// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V6XEF1n4QkF+dCiGjNdK3OvR6h+lBGdyXyOSNqrtc4xBc7gyAH7wLNKcIhbM
yoQcVaQaJ2ojadgB05CxKD/RDEqV7HmxUUObRleXk+xOizgYvOhBHFn++I5j
7R7pKEIdsHFGxtuG2/z7JnrC28/aqnTqSSb7LI09VpeBR3i5qQTUU00Sgbpn
tgdY01FvrNqU0mtFPyO/lM2u/BNgOlRfXjGsJIPAQoXYUG/Y0n9fYFzWZxS2
TX7H3qrltbMGhtMuQ+nWHN9bQ7qHb8KPtlE51nbAMeEzQDy/7opEqMdl/PZC
ljj8xarorQILdRFy2/NzmezSLyl5lUxfiHZaUJWbdg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JkIRgQmHsmZvinbh6f/JeSabqA33opeR2SIpcyZh6X76yTehGyBFMHjRvJUt
qMMXq2Mu0ZLvVF69UfVlwBw9z5BbI/2z5dbCp0tBQ0GHOnco7VVzq70q0guO
vIUyj2LK68FtGZeT+PQr7CpuyNIYK5eiH++oPoWVmz+LzXvxvPMy9shTfcod
Utx6sQnOpOAK6w3oXKbxmCGOM2kwX2hLZBWuE54z4xYRgragW93si0bOaEVY
Q9dClR8xR8B9XDQ4i7PNKHWzNepcSlbzkYLz/UDv11QM37gpPEe1RmHdZ3Wp
fkTxoFRoI2fOKRdetZNy6RAzCeNW+L+X824wLxqtmQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CGpr3b7NZWSXCrl+dVj0QZvA6vD6+JwAO34GxKoTfdMqcQ5tC9WsRfFpSL3l
S6I7V/f0R0469JFFUbK/CiydVLuziOo4hCay9QeTSj+lvCouO+uCPZGe/mYC
mBj8uzZ465zYjeRq+1I6rgln3oSWfQeU6zq/wg02VTpzsSC/4U+2xvbOXwMC
nBq88OF4IG4tq7TR/Wm+W9w5qWY6ayEom49wx9xH6u09m//ha+1vdZycNyzC
AiSCbTemAeuYEFgscIVykv//q5CG6j0UNwupRMs87tg8EHyAuylGX9N+kto6
E6VN8tGFWK4GE2Gz6tNzcHrZb/uEczogx1p9ZJ5rqQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pdqr7mjh0I3EiQeD+0VY9lRmR/xHwB95WPNkoSID0ijqC1RuD7LtbxXTv+dQ
Yp+kfS1egk8hLnm3088fwrj8p3kY+szYEiZKSf5fHxYntSkJ58tmdLYWloB7
G6sDYDKf4pvEODZBZIzYUAGYGsEDxUqA8BrOw4h1Be+3dE3d3tkhgXEpQ0Vv
u9bl5gI8bzk/tCmYNvjH++7ZKvDhQL86HsJDcZXtEHBHotj6yh0aW/7fFx1I
MBVgy1wojS9fZ9bPkijnDegzNBCwmJ1a+7t8Wf8IvpWrChDkPLcfypCjJJA+
7jAfmEQVoMXsLJNeXbczKluPU/CnA3SI7X6FATR3Hw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IywW2hAOTJj1Q9JSkuDZmECyVqOXT5JvrcwVU1TsJPkT2SgRWqd4SVVPsLuo
bZeJcx+KYVNM9I2CJnjlyNfCPbesFhB78K4pTlYgitacJAi90Oo+cMsVHboH
SrdJdRQYkLw7Zbq8q2TlOeodNr/PEFdytoC2T2YWBdrKaGs4m5Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Oj6X4dRc2FBMIhyEBwGjXLrAPRgZ0R39cFXkRceJwRn5td5XDEX1oAk7hKuE
LCuC2NSb9H0dE+8jd8aupttuQOmCNRKRWbh61R7yZNniMUgg1qf1aGirdHl4
44dBZ30H9q4nK3//hm3dNG9EjuOx8ttG7ye0zbpocnPayXyBLhrBYNcNdIzV
2zO/gH6s39H6WONkp3cwvODRwCTFhzLnwE44ykwxpokxiIE6EnW9WcDXdDsN
KhAvJmHcqdjOMJe5d2KTqV7ie9+lczTdpBiZD41cr/1/fNL6RfOoNS/1Valz
Q0iL0xmYCE754hQM2zLMEGN0lXdL7Ab/YRt6OaUrxknNBinwGJlXEqCh8yCC
zSCKOhfL8DMZV4PySGkjB17qxJWCS3FqrppZdjIHUkcV2xVXf/FdqsJn4+eR
oNq2dcdjSEUwpvfgKwMTW/2bXZFXe+mFHq4XZ8GM96F684pZAA47t020USRE
WMGRd/e+vTQIWQ5RBN9U4jFuxR8k7bUF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KDFqoM+qeGguJro+hOA9m8HP2r0cmVPyiFlGYGkMVmusgJ5vV0sElBWAeGPR
nsnRb4vP7zreZMScJprc7ctrz2Ksap8pB6GdvOd35e7wo7sovM5jw5JHIyUM
vv2jjoGjkdX0MbINRgMxKY1nf8mxhv5wW0FPN4aAP5BOtqTwK58=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uL4+yi/CId9igG1ooqpGIopa0D+jbqiMLQR64XX/vcmn3pjvyfI82rhRTEXT
Bmf4ND8ksbahMb6w2hpReEzXJhkk3kvg0+hEyFGp32B/hy57HKzq2NLw5Plu
szimjO6NQSXs5hJVcOrBrMRkQeXpJ/zygKlS52hZPg1jUII4QE8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 253856)
`pragma protect data_block
dNhvM13XFepXWCNh2YJuqJBCe0M5+rqtekRyKOWqzdEej8tWWjTg6qsFxRUD
1+Vqk+tYbf/Y8nrv8n1pVEeG4jXWQGuNNr795Wze4Yq0ZNZJnY2TlOE9N+Wy
4o3QftBRp7k6ZkP9zTGB3RkPa1yISfw392n0C/pA8QzAevJ1juJagLs1YeLW
ocJDs2G/Ku/bSVd9ZEFEhtsdABamUoQlre79j67P4W8bIh1SgEzk8+2gKfQ9
MQK8lewcShfYAUf8+b+6RWgviTI6GfS+4o+YW9XKudbB94jYDQpBDU1kYrbC
pL9p+n+i6W56tf8+IYtp2YhOkjfQ66Z93OYoJfp3NP4Ww8WzcwTFFTNth0Fv
fwib2OzPk8hjffxiynGAOemrbb8Oupt7hiPQaeLyMtHEwlMhxlndypCJwgdK
AWOxbVw/Wo4m2MO39F0m3XaKjW+tvBHAiOgaO37dF4o86eiimqOXTDfx2zoc
WKyFnnqMHR/2+eQEo2BPbMkHe6qnsJydx2043Wl8JgQhqsyj6CzWfhXw5+12
9BOg+KRUKTz4tfGCq6gvfgg6C532MGpHb7OfUFNpoG3wsBEJ2wexFeHXTEJ7
cknrgvjiENuL0UhN8qeysJ4fB8iB+vaFeNr5cZ7EBNhJezCnG3VGu409Znn4
0FmEM2Eku0zCpUwkcCvSvKEAS5jUi9xwk+/O4Cgo7AW9rdRpGp00OGWNA3ml
vqp9Ee9q7PD/WSubfLw+7uDfjEl0GeADvmc2ckGLVKqdlwnb4wwrtbBIwCqW
JrGQtOi0eJXybPra6sbvhmxa+gxw7qupzkcU2ZT5q178lfipgul1b+fORGRh
IMaf1FeQuvpEuoRNBS77PsYDndCkaiPBYIJbkB8h/lPj6cXC8Qo7Fzcq1UBU
3fQcaST0zPQMuLtoRNua3XKcLJO2uD/PIsfVSuHamDs33i/i6AJP88qWaWqk
5gujgElGjGMugHtItcszZgETfdyjFtxE5qA8PB9KrEAdUOsFUuWTua4C5LCw
/KyHcoQkbNGrgGQOhxp1/W9RXDjYdVBUZV8R/FzA9kgg/EoqG4npcQSUye+E
ejs15rhiOngaMS9w89qd+WclNEg6OcDDMdyvM0t9k3NHQkOBqGNh3TIafOWw
Kd8+ieOM1fv3zXdGpbGLy2mdKvXOZyye9dT4lGR0SRs6VXOaA5XU91SxJPnw
bAIEyc7AP8HRNbC+IcNK2TyHFJ+cWTfCRBoSMSKo/uyuHfFh64jfcDvor+6l
SDuoR22rlWPpfROrdWkU8/cLgLQoqlW5aofkmIMpEHI5njtBWt1qwqa4sxhv
6Z5+GXDAbbfgsiGjQwwuB2RaYA093/905Um3PuJRHyYMNEc+TrjWc7gva9B3
B6GzBps/clBVLxqVQzTc5SdV0e3SUAn1H3MyD/py6zhR1dx0UT/86Q5LV845
Ac2KRWvPjrHtX0Wqh6eTNBxgOSqwsYaHdJ91aE8sYvmihfDvCXjUa+XpMhqZ
vMFVasQFttFz7t0xYVBlh1Qy3O/kGqXoxg8Zr3ubtIAskDylYhHlmKhMASVu
czASc2klnP1RCNh90BJUKI8pe182fGZT5cssvizAfxThmTSBBkIagmPBPgHX
3xmQYz2IvA+O/kTTtFtmz4KH/kMWcdc4Malfobdyyu7p/mWeLCjx8rVM7/y7
twwpyB8ftaVFHl/sUomHbawxlaO8KixIL/mbLe5iWVEjtAgb3e9lvSYrTpgC
SFksLMCDIjvBEyKseSNdYGtJ1GrE+g7G8Fws+RNNzpDqvbpd6tK+sG1yCy7z
bM3XL0naOzJ8Q0XHOpPuohzYUO6nElgHq1t/+g1TbCwvQUxS+tMHE2LT9vhh
derjsZjq1lzxpyiIerx6y60RcWzPIRTWH0Sk+jZSoDYKoZQ71RAVXfGi1ZQt
/nHjY4V65x80Te6DZGiC5/JgucjMvPiMHIngfsit2J5Ngd0BrDZl8M6ePaVX
C243xv+AT4gn0BhMfXoMCFVxhTSDwReTmczGguY/ogGqrrx+NVnWE47bYGqz
Ak+GDxSCUf/pOd1/qqKAuTf7YvL6T3m7YpwPiOVqiTgm0Sgk8scV2rr1jiRp
gvxp6aJ1bO7cktU4Ria2BVrvbjnBjpZ+Yj2kuUlMl0h5X6HvhYn78T3lkxih
iKA9Dcm0L7lblXpMal4g9YoPWy9zNxGCAi+tJ1oQTmJ3LcCQo9CzCPPQ6J9/
6hbnOCH1zzOoFrIOlyg8s3gUxfAESsGgPAbhDzwoJExeOQVTxdkEwT5y/bjC
QLfGHPKMmVSyTqpenchvH5WmmRflF39MdpLFbWLSosUMF6kTaJ5JXddZDLvA
0XxXKhWq+aBRUlCGdjPjkO3EHjKgJPcv2zWnLkRJt5Xz/430/JUFTsFE5Jdw
MzJ7xC5cQiuK8K+5ONwh0+Yj+YL+qDvbH5X176kzIMYvaFbSsG5ISGLewjXQ
FR4/YEBkZW7z7JF19e6GFyHbonChJqCYn0FHDHIhKxUfik0mA4hoLAFHl5I0
PaCGu4RxcT5+mA3HM+9ZQ9ziMqX2q63n/qYM8AWALALg5gw95pmeQLW36SEB
gNt9uy+X0izFCJgp0+FWZjZnnb6JH5eR52F2+UXmtQj5lrDCm6Vhdza7fbFv
FXzaPsAYl3FVPjPOwQ+jjedVTffLMOZZyvrVmCJ9H89h0vuCK3HvWZtCI5Lu
R4dA7UUWwQwzXoz1nw+9hnbsTDyjmuRablupw1APkY0qMQK1WnB/EznWGQyS
Sf9uA0bqtLWhZdpACazRNxe2uqSLSWSIqNyEkVJNHGvooRqKLirBAO34aHXA
bxbKq0z9npr4dfSvG46fjmEl3Wp4JBGjw7ablRAEVkd/PZBrIjcPSXjm4ajt
FVj2KXAEHVhGo7Y4ISb8ZRM0x3WLCdn5OrlBxDyRUmhoJmMxycYAH3B0wJT1
Vkb36+8Tw8TXU18icm4COd5tZrTx/mCjZPLueRPsucSLKZ8V3wnLrg6g+HJM
cudbMm7r/gCCkJObg/Kn/E/0sAESnDx3byy1HtbSoSg3kkGwSCdOV1/e8IO5
tD9EgeuiG3Z9R3tiFS6BBhoqds48yjUJP/IG0iUYZ0mSixwIX8MwKZBOynIC
0l50Sj2cE8sTAbVwQVlThJtM5diCo7n8Un7wyXvwzR7vgGCYj4hn96dcedwe
Osth7mIteyuPvhXWxr3gU5FQgrqC2Cx7x+v8tGFo0OVldPMxsi+N5LRrp6/L
B5OI1YF1zx1F3oA0r7JHHQadWYBVpiHAXv8dOPqcJXNEb2MnK/1FlAxZ6bjL
t6RymKDwTDEB1cgmp7DMkBLo+AQn7zWrKp4q+Cdggu4HfjpSUwI/qduYUP9z
I7UKJVVz9u+xODa5SPPsIjfy4rGQqfA1hc6/48ANlhc3gKldXhfw4Z7LBxhh
X1PM8XUnzOxAufYcxdYHKon6qCnAb4mLq141UlaRkq8H30OzucAsUczfm45o
Re0BkdCaZ2NYURPr3m5Nj7L17ddMqxqZekPqW/cOkMTMRGLHx2RVyAZmIj2y
io2oCyagcGIctIa8rbR7S5COD7PJRLSyOxhxm8jNFPgmS9UkgvPmLnly/A84
6LwtZQsXWmREtVzbJ1VbQ4dnuPv0GSISta+WAega1euA0RYPpUQswHvWcqYZ
wY+vtqgfM8oHc4teu7+RRwXy+DF7YBbmoUvbDhRvz3MedGMA+1/I2GIyJ/HG
bdIh11HenmEDv7fqa35FrmetFy3LwxyHhv+8OH5/fNb1SOfN60tPGIxQaZzx
JBnoe3WG7QSGLKrjcAZPMUqor0i/Gy6+5N3XcT4R9IBzr/8sgiE6BhLZO14S
1ZD81vjlN0vGUpUV7z4xTIetr6k89eXXWa0K/Vzj36P1Es8p1twU2yrW0GhM
q+ecIlKQC98JQ6WgDLF90iPehb5YKY9kTUHM2yrMKHsniWpf/xoIXyk0q6QR
aVh/DCBSnHVXBEkdgR4TsoSSP5QVoPFlC/tNqbH71KBtCk3KrV6meKSBlM/F
LSy7VrHEI85OibLLAzDlkAmY8zB1tetRxb6YlyJa8m1RiI7YYMT80AHwBddM
zi3STUUmh2cYOIF/I2NrBKvQ6Ji5xaZAwWLoSs7rlmJDI4xSW4kVlHYtk78z
KPNsON4myRrQuPpvirkzXB3NgHf2DMemo189KzqkPNjiLfEpNX82DcFwWwXM
dOeRfAWyo7lStd0hMVWUz9/hooXdjSTBbAF4B+4eFN5owUtf6oI/mfhUyn7j
/A61wZ4anp1Rt7MVcdGY0dB6bq53+XYrAILjCKYZ3gJ2iDqdsodEobsKwfkJ
mfNFi/65XBNqSfqh1rgLxObbSQO6yx2cB71eOyvNLT7dUpTQVCeAU7YDx9dg
ucT7XL4fXmhNj0ikKJrZTEYKindcneRUhVDIZgMog98un9lQFmcVFGvWHt6b
v/iGP9ApcGbf+Z8cjTwhY6lJYtm/axB2FSgOKoEsfYnzClu3s2ehQNZhtlL7
B7b3yPx0k3O6ovFh+Wz3dH5weHNUE89dVQBGs2XsdfnJIfocQhvk+BFPDrX8
i9TSQF1DL2esUZNrOQow5/X3L/+1Kdg34Lax4XRrYj5YLpgm9rScaid+zlvj
ZIkSYv3cDoLh25yBWVS+577qdoCEmyo18revS4t93HZvaPNHqP7LnvJPInHR
H4YF72Ksdem4Oy9KYHqEsUx8mjA3L7r9cKdTXdbNUce+kQ7y1EYTvEvp4L81
7irVBlFZkRwDsHMAZHPe6s4p/BsTGFyWFneOrybTd8qR2pQY5KoKEHKskfZx
uU7dbJHYnsWlr5lQoeoUTT4HKSCEg1ATtjIbqIEaQ9mq0fKx+7b5r5hB8bsh
KdGaY7LVBokJ7xZcQol04wSYlYazJdJtVAnCZQZx2hPxhgXaMTP0A5hosQNA
IG3X4T8U4jAgeq9p0Dx1sKNYmTJiZPtqSRd5Kx67vD9/x6nHw1/fIOSv6Az2
mf9T+/YL6/iOHWCFXCSGUxB13AKPI/gLKfmzlmTmfl3FYc1b1FkLDT/1VX1G
Rf2i5KrGeRt2j4axvABsx6+sjbkLDjrLNuHqwYKqpBoTrGYNg2TtJEujMaF2
F92wTwehW6EfcHS27oV1XxDNZpXoo4BTpueI73YT+9RUe38VDhwoVatDRKyj
vMv0IwjVCtZn6sKxBqiavbOFnTUSb2vqB9aByC0/VU7XkAEFGUmYToBO2KoD
qID1GQgDYT72m3l/OQFVrW8lcQhvmCCBNhhnwTV5LXxGRlPT32qteuYS8rS8
zeRnIp+cA9kBOmNMV5Qf5jhY/lxthxsarO0Fk2b6xe+WLL1XHeLORFMYDevU
MdW5vKYGSxezgH1zTkAlq3am+/KVS5gY+bWvA2bHn0kOP6y5UmLcBMnAA/ab
HwrKQOBAUP76LiF8RxTOL/034EoDAvtzTtV0R+M+LyhnrGr6bKlbAT3zD6AN
TEbmiXIR8t+Ri2fr/kfSDF5mM483Zi6us+q+2/34OoQIJ9dFhDpB4Irg1k+e
Q4e8WOP2SsTR9HQqpBruYE4gMKCCEzVCuJVVEsL9HpnRRbhylRuu8jZA+14A
IlVCfxIksLhK2ya1ZDLcSeHFa24dAw2f3ZE9EuCEUIzr/uPsCS4QoitVXY+n
VXvjjJCLltJ8etX1uqWRvXDemZ5h2hIINhLnYuI2XQ7/UYaN9aKhyQqI9a97
Tl858iRZjxKHh6jXSazr9YDa02/pgrF8VyEdurmqyHZR9JWOnlW4PVihOkz7
ViUE9nKTfzp4vR09dVGWCiHuqe7c1910wBbl1CCeIlDlPgWa+59ILlgmAzVm
zi3LfEkknf80gGDHt32YUygiY+b87BPyVb8JaueKCaR9iVUxR/omBh7qoNP/
7ywp1/6Kg1ppLVxt/YTJ35ZCXm06vxtnynUZipg1o7oZIJKrTevpzoYwpxyR
5BjXGoxJIcEU/qrmr7GQziWrT748XUtxv3eDGZkNznSuGgKF80zyhyfhiEin
SoEiA9SIsHkNprn/4KbsJWcO9Up6e1B0PBxUcWtBYVe7UJAZvTPpfGio5KRX
uE3FwFpdeYEotI/k+a6oZvSwhnhqVW4omNu4/W2y4npQ4/Z2Fbj74voxpMla
fTyPyXlRXZ5stBB/IuawsRQG7NxmqGbe0/RgKUaH+CBznhkdpINzokxV0CHK
o4E7zYMXub21Mn/39JTg4PC1SFlqsMYZH/zMUJKyX+EUom3utcZH11Y9PvcT
j8if8oKmFOXUqgIQTEECajybnl+N49Zo2fooP4zrzv8RJEVmKt/pWPUTo0ex
ug7JjgpSD8YndgB+FPJ1et7A4GdJHJGd2LybLaJb043d8gj8celeJSsWDDXK
gtcFSTpW5OgRqm60hMPlAt8YriVjlucIu1fHMcwJDwtr70Q9cuzH0Fu3/eVz
NNE+vojMHn0jQ40CC7As3XoPFv0PTrXoqQalOOMgiQdQz56aDimW8pq4ajxE
bv1NH0OxMxIgqXPkp9AFDtPElpKMyiiF4IFo/baGHUdCHlxeuYTV5y2eWr1z
NFW2i8x5lUPV+DKb7isYea6KkySOV8AzfaWwYnwldgQSk2Jx6b8LiXWbjsKM
i7N7PN6tKg3vrXNOiZv/8tHQlL5h25ObI1aJzD0RIjWis8XL9VHLH7jemnKS
BO86g59HjFnsxzPOu/bBpkVNj68J6LD8SHFHeaXwXZlcHn4NYxj9UGzTiqUD
VHVfu3ObuivOipFtiKPpBrh54xCrGbrQQ0OpgrBOUDp2z96JV4fjQ/Bf8NAu
/x3HN8DMfciLOFEvrnHx3rkU+mGH0xl5QicBFGmvEycVgtVcWEILTXKLaZJU
UzOhTqwCEdlfokhYnykbPUs+991euqtkXx8/ZBrhrXOLVstVFPwxh6i/A6kB
VBXtzLHe2aKtC1Sm6P6dOWin4rrglLlDmQjcnsn+VICBJT/LDoAMs/Dkw61s
bAWPsetI+gwI5pJB06G/7tw1Vgyy+I32bPY+07wsyK+78mgK4PpeI/MZGtAn
a7N/rJ1EnVcKcMBME409O91caOfm5S6JFE0kVWw6RlALCls1L/Dwzmgaz4J5
iXoCS6Pf2eWFs6C1+Q95pnoTVVBwipv785/XGn8qLUe8eb6uB10K59zVfutL
08XEdO1N7y9JGtp5QdgYePQ091wNoJEgVKj4gz9ufE58oi7NPSUATejgCIw3
PhsEKIpX2nizduZ7ULHT/2SZUZkNoccMXpzZQA9JoKqzZOjWpe5CNcyKLGDb
jZjyLN0o/3TXH8B3op8Qo9Ncz0phtqwh4fih2aTIAA06CbdmGtJS8tCAHj87
LhkOIBii2uVyK9BRLocF1ddkPB29eVcglhlAAG75Bw9Tx3rLpflr2/HW4MzH
nrfLf28dFhWg8PbG9UM8S3PLEf5E5fzBiVbDUtPfHDj0VFVQRBSDX9UML07v
DibyQuX568CJZnk5YQGDtwUhGblXxYFX5i60evga5wxzXMmWX2ZgLm5I2NrC
vqT25yI1+rF5u3cjCj23zeE7XzWiP4rktBlQywWxragod21GbmjIHtGVahwW
rbwQXeFY951BMtEns9d5Y6+6l7Q0Qi8ntJr11QK1JYuJsG7oT+fdoCJED16Z
uW+V+m2gTwPlhQ+R+iSYv5GYx/UROYuRRyjo42WbwMpS9f7C326KeuO+rjR3
rd8WARW2Ka11wZ65X6rCWT5A7Y7Gh1Ib6MRztZRqhlCl+37nCHu4PlHa17zo
aycEu1+Rqoypckag9+xkjy8MnWSeV9cor3hdc2TG3gX5XY0Kb/ZeOLHnUG+2
dGXjfP1oSFz/chaOukzk1iddpzU9Ozgabpm4FEwBFaAQDFEL7aUt4MN2gftp
ajcytpXTXs3WiuceHigwee+loEv2eJOBoeTz0bQ0XrC+3GCobvPINd/oJZBE
ewhC9usdJYlNrD3WRzBLilAImmd73TZzHFu8lSAMc7QtSYR85VDw+J0MngRo
ZdIBmZDuVoMPWdeLdNUMc3u0/7dE6W83Y/yRk031czKtW7ERGN1+hxgwrWE+
LLYQgTJfbbOFf2McYtJtW7Sq+e2nB+CiOGNhG4Jx+SxvHHKamcFJQ11Io21s
RRuoEDKznjmAO9q4wP+SpRs+Fy//HMI2v8ulPa2Znt4GcC+ynuFsienlhrGp
F6EAnyPYvejpdvv6Z8hYPKuH/vPvyi2ktQhnopFdtSXmaR6GlZ8W90VJIyf1
/4cPHa357Gz4lic7qAFJzTgqG5vZdvWtm/awv5dwAR1CJBIojtdHX9usdl6y
77dVHus/xxrdVGd38R865S7HX3S2BU1tpPUAg4Bev+qTPN6E+kiJTDsHfN/i
7MLCiY+vWO+0mV0n1esWz1eKfrva7vxtbBQSrn912TTzQC061FAsJE0WRPSU
UjQT4HPFPR/sk0dl7y6Q2u4uj2Q752gLhNKx6WIPJhXzdENLQhuyaxX2Q3ze
Dr83spZCEfHASWe4jjxe1OdJFvtcYX5XDnAnafeEjpL8eQnpMv/MGbJhYXZK
pMu41auNFfiEdlW+wdEp0RrGggosOcGKTNFK3MaYjUEA78cA4kIjUjfO3ZK4
ZzE0raKIV6LXWwsKcfpWzBCHuxTB8trEx1YOJ8FwIpVFWYkairszI238ry/Z
Y3nCfnm6sMfMTCggpmCqwiWJAFYfjvf2ICqtFjt0ebiUvqoSS1kpw8/aaETb
leTN/B3JXL0Ydz1os/t4fOKihaXbxxtDFvl8W/ObSwywdKKhlHbm4zaXcRpq
gUXXOEpvR55Yy/VKFM4PyMydOuNk0hCM21+NGPqhLJ/t47nB13F/0TIxnBAS
L8deXt9zMXN5AvDSEPJxZSjdqjfqSG3M+ZM/ucBttLuZ/FJY/aphwiTUKdf7
3Qw5sfesiPH81NHiLsJgOQL0ZdmsQ2DBzOa0AO05+DfQzDLJrCZ5jKJ1kMIU
Ne84SvkQREAyj1yEwodsWAGK+01S/hykR1WEVpuB6+w4Pmn6fCqGEk3FOzVJ
b9Q8STQ5oxLtKj0IKkZKODJnv/svxd4epl1DPAjobnx6DP9zRSE5wFiXruV0
9gXRyjZ3pT7EjZ8mSH/u8bIIR+kjcL7LHclDmsZvLy7nLCA7gEN1Cy6Fbx8k
I4F9rHKklalY4LR1j/jBJp5stTTUGsUdF4CpbCOMgK/j/SHFhNsVmwqRAPsj
Cx533QlWXoASVio+Lhr8MtoknQYgDn0LUe3BWQXGfbU+IqzI0RLOMd6+zDUz
+8FnRpEx2MVg8JTDgRssv1p5wr26HI5R9FhhmYaCx3qvEwXIjP570p3Cg/tQ
YTl7Z9IjZXbh0pbInRjttW5/34ZUvGHHgk3qwqF22AezwW9qZbSKMy+9bxpT
BRiLSNDsQ6dQBlyESVaWKrhsQFJOIgfyp5rzXnPL4BIN1vPiWER5t9T9ELXa
hzE2QgbhPLZ99fpDT1jqvrw3s4ckkksH1kvJqWTEpOcwDdc5aECAMSOpX8kO
nYc4hzT9fQt68NgwHVA1MpugYbj1pdS9W0/+9hCWogFbtTmFFxkF53af3poo
Bq4MwV+RvDumftp2hxlqenismZL+pQgx9w2bBKJcE5UH/Vyui6saFmuOPFHo
zDAw2whv7daWq5nJpR4m73W7PAZGaoZgss/H0dbD3TCha1Nc2IbhsOFT5Kty
/pRAQpksV2Sbi/ZDETfg9sDAculU1YEhv7roPvdO3fV1HqN8eshigPNoe4bj
AaCsEVo89xxVh6SzOfer5fzgPBBul44Elfdr2WgW9ExDDI+BHDLj3xdS8rZu
f/QYo14QVpIvA8HQN4YhOjz5ZcU2Ve8k8SfYJ7Cckb2Ku+zgSo/1tm3PP4OD
XoZlRR6QNgyO/V6gHByguCeLpJjh1NlD2bqNoCdM7J+UgTJqrgNmbCW35h2+
1Wjc4HbVx+N7ssHldfmPwIj0ByLnZ0iHnY67fNvbimEpQRobotNjH8uTr4bx
wIIOwo7rynhJxvIDl4D966Drmrh4YO+XCpSpC1IPj1zkwFiMpUdKMTNz0Col
3D138EX+CEtNYXnFKuKBqX+Hp+xRHUXE/KvRHp5SG7/s3qStbTLkTWPaCRpI
tL3e9WJpzZzWWLzw5Fxz4zGtLuqIX5HVxROjHNMNSKJQrHho6G+CbNgl5S1E
ZB0ly/Xu9GHvl5VoJIFBJGYC9p20S1dEx+iNHP2jsib/64yy+ytHN5R4RVKp
TVCqPIhOlKZ/k6Qlxl96O/IaUUTJrodpNDqNriy6tzbv4Xm1LB/lTrtOe9If
qBU65WvUinvn6oclR4PnyK2i1ClWMVR1q4YE2q1ASFfMzMIoMh5s8xoAgZDh
jNVhPLaw+XoCQNjOMyN44UIpvZubQsXEvj7IZ+mNXCuO56cHb8sl1wbeMan1
oEFDaoea4mrxnAY1Jdrv6Hjn0lk7fbeHg2WGCOmBc6iDzktH0ekE6QLwlLFB
TOcRiyb5WAfqAUMTTqdM8nWajLUAp6Daw81wSJZVNhUBwb/FD/Y15Ua+9k4q
fdh04OLJuBgqUHgfyw9uUwWCYOaM1DH4H1l+VmNktRb8DJdHUSROO3VGY63D
WkYfgQ00VuX5ZmlhEedJHS+/lndUNr65lYKVWK8ksCdxN6H7U32l6lrGj6BE
v0qMB+uadjju7z89OKSGiKP5dVu5h1Hbwc1OuS1JlLfAvtpuX7jZXmWnO2b2
OzgauEwjiMlVcBX2tYMcMmMifWxWaNNxreQGnPn8eZhbDj4sjPEV0FQFsXlj
+Cw8pp3F0NFylOqJ/GBp+dN8frfEeEzYxyyZJ66Lz0pO08yX9+F9S8cidlLL
0J61/B0qODTzYJhCvXcXo666QQX8hm/dCQWUBRMpTZCPQM92kNZ2ZycglX6r
Dcd3zg7nlVIe5kH60sJ0NGoArzjHpHsA/7joO30hAwbKUkcMRpUn3rMKc6pb
fWO8P1MWjY9gtaFARyqZl4lTdLMNcn79TDnr78Zk5Gu4560nuLS7MfZYJ3eH
ZFQiePapY/POMDADnfeGFz39FLVQnuUt6KOqohXJesBL6t5+Z+ySafIEV7Ip
x9qkG3v8emFHyzeXemgt8ut74tarml6u2OvDQ+bSzfhKkm3/O7z4/yYTQFoA
cWUAwkPzavql0Yp1UosQ/mHGn5EawFvdMEWinQYKcPWflzIumgc9epJPFPW/
9M246573Gwld5MN0J9rJppcqF2Pd9Lo+F5d71fIYAViXABovMdXqN04DcLHa
Opw9bGF5LqRHH4sJagU9CeoGuUSy4y7P4VqSopLceE1SIA6+ybsFx3NCI3i8
u05at0FBv+fUAlY1M6pKF0ZPBmn5tETdgndVFMNUkWt0JPP0OCw8A1aZ3cIg
1azzbkaZCTrf5LMAo7ifnEA6xKAPEhntvxraxHexJEdrjdPXiXdWhaLCQzN8
I6dXOjc3AB2pN+cceIhTnE0Rgcgu0R7/6ROHnmgDrN9n4IZ0k7Ydhn8c2YsZ
OGRs+B/P2jTQdU731fHzsfK/3vAYDGu2VD+wWXUEf9ROnTE019Rv/99/AQeH
82hUjo9hqShzrIgtV7V8ogx83UyYGHeu5f1r25bkWo7vmrmpYjsw0j4kxW6n
lQFyIFEWKtGGMWOo0QpmwNMm9NoTAA6DR4+RF3sSytNZToF/arqL+EbNY4Wc
vgyppajtcM3X0IVjJ7u55TNr8ZDU6nZbhXYsiUyae4ugmuT2At7jx02UBG9p
KlPCeI0Il9WRKgOcNCmIupcRWTmxQvdTxp3rrtWEHthI4iwClg1+ZoMKte39
gySeYe4OZq2VF2QSq6J2vuVCjzqyqHF8RfMwEAdXH9215IWr02SNlbYdGbQF
NDIXkdAfM5v7sfgp4bSWnB56Y9ZoI+XbYdHbbAK/aw20VkO6AZdKiVP2VxNc
7U07zhtkyJcN0dvyZYRhaAjjjDi8xZgZ48iV67RAUKD1Eddz7Xujk0mCy4zh
8uyI62WCN9ZtLc/ToZgeRCYjI6NFq2iqnPO7jTY02vN1IxE+K4tcgyCW8r7b
AjB62Y4Q9KoQCf1YpSSJCEu2E1NgwDODNQcV9PSi0RVff7p6U9HibiuSA90S
Q8AVYMl//EgTOmYkIJwL2qBbp57WY6MUX/ogg+OWJzCe+XFC3SX5vBFzjHob
zNq60L1X8Eq5kLXJU7AEJHC4DA4RUa9po6bgxDbLBfyv0+OO0CDwK/Pc2qJg
Qezal4J8GRvBfJCD+ATaLFvOOHNInkwRECOcIrQeyOf0FLWjwd/DxHQqXQ/Y
3FMfE+vWG9Ljia38SRLqwcNoyRTVnrOqtJDIVc2sqrMG1ae8Cu6aRhsIij5H
FoIWJphVbQm/wPpCxyWGgPSCBe19dPQMnE0au/qwgElFA2vfgh4c6xpiZyd7
wYsxIgi9vXjo4Nv48ofD+PsfHelhpPJ8/paaTKqtp74fNfJO/eMcNkbNnl2w
ap3qGJoXHlAWiGwCAWTXeqKJ/bzCYXEwACAbxuIIRZjB/2obJsssntnVdeE9
VIzSqzAOpCrRE+qQ7OpdOJ0rh/uXfO6sJ8lbcVNnDzShBZp7aew3CX2RAjet
79E3in8i6C4N/o+lDYR4B/nU04qz8s0DhWD10YHBqAkNOxp2aihESJ99fdxA
iS0Fptzy2zZ7at/JIptf+Zr21M70R9ZNQdIoG7v6F14nOrhQ4IInUeMBF2ue
42IvYAEojsrlTNG7lV4QI3YKWlcCkyBRoeQfUKwdC3yFfnZ06ZtGbawVXCHW
MRwzomJoOWWTyx9Z4BJkwcK/4gX8wSpB9p7xNbAKqijcN8wmTvj0BWmwlgJL
BoHUISTKR8G5cH2JJ5g5hBNMNgxVeyQGmGwSMNpRizIcpXLoBziR1Sn3Dgp9
CEXf9FT3u+ojLzDnvuDbxhXT++n0f5zgyPCtghoVfWno/6ZOqqPSuwOw0/uB
0onJhmEG2ErxHeGL75jWDHt4OSROzCS1Gj7DBwB6LVLgHvCRaqG6wvmV82Ws
AgiwsmIvhcMWHNo58fsbezK/F5A2drRYT6zZ8Qcc7iTknAP/ID5vQEqOltY0
mO9xqP6CIJmai2LCJy1Hgg1464GERRQgTZN+CH1OGXUl4PxNfmPhtYMiGDF0
4Yl4RHNel6gww5jCdbt47rc3iD6Oh9ucolGo72FnAlBl4l0II6gxn6Is5UAl
wtUe6s3y4gl8dNEe4lRhuKRLwWULT8zKLLAKO8ok/4HfynmrDpOGkjmBBOdO
WBGw87TchacP9uhgMhtmrh7atL0cY5Lb5wOzAri/muv3Tw9ZANTwlrM3vwoO
MTbbaoNipbIn0xBS3V4+oO13t1kiOP/mWbjAmn0Bgm6udOCRFvG4J3p9hprF
2QSIBGLYLBduIBtT06qcGz3P1TqDeY+iCfti9mLpIPGYGuAOOuvZMqAhVEKC
+0MYGgPbGPbqgmUkS9SW6ASYh2bqO7NWFVt0WojLakdihbJJDYNIZ8YCoNab
tM8OiBYniqBLc6UDTwfwW7VT9UHFgPKEl/IkYcF9OfNcmKP4INQVNdtKdYFt
O6HjgcsKMnr0QMPORMHbE9f9BaffOynA1P+27V30zJ/EyXGXdV2NnfdxR4Yo
Yc7u1jNMSnGQZnY9Dd15usMXIFHH6TZKI0sJnLfYxwwN7VzvAAZWAVK+EyMc
6R+/MxE0bIfzOkWnu0VESjbDTZMJKs19eDV/pxfKCCeRu1sckMriey9W8HBM
hbiQBfjLitu12kVG3vVCe7hTZkenx59QiRDO8wOhxPderLeB5QIM79u17ypq
wIYB/h3QEKzw8c7dikhrZ/3vmVZHS4wM0lTDT7Oj1JxlaFl20EjyjYRWgn4y
wfoe3snMFBj5JRxQ+a9cdNH80W433lykTqSpYYovsP/I88eslIjju6befhC8
LP1BNOrq7PvC5wHIN3XLDy0F1ieJ/92nSlR/Bkb+LOXsMpm2H1fsGgsLk50R
Qc942uQzVDgCXwot2hDXqwOzmsPqr3XEVj0iOA4K+fa2/wmgR29eJeQLDq2o
0igPmTrWxh4OCdv2MPGxJmSP3ox05sBC8a9gqgmaLZW0V73Mnbtzv4u83MPA
acKHY0rMqNjrloJlGPu2NHp0uXXZcZNUNnanCK4HocVEDiqLCnMSZsJXnd+n
rSnx8Zyg8B+6gz4EDuU1mFqTelpkH0ZWI8WdukuO942NM657ceNEDt4GucVm
tUKKlQH36891VgFBqBLQgXGC2h+36+XArU/bgZw4OqVtn8BD1zw+VwUF8zVX
0qmYqZW1h0s6XwlWLfOt7u5aJRIBK9mISsu45GXidozG74AMksByJFCgMxAD
ANdEPcKlRfWaAFgaVplX0VcE+BjrRDHeZZq9PV7gSLkj+II232IihBmePRIu
VzqwqpKObZcE6dGnojdmN93JjyEyGV19z4WxI55/aQPZwMjhM00ZyzWy3jmf
vP7DRK9Jr9airfIc7pPoXLE1Bmjt2o2P5C6H+0lXOwm+nT+4lS1hUIOfbsoP
7gMgKcsEUOH5HQaew1AgUedPS36lJEVHHwHDiQ6OqZAXrXPozLgguzBu44uN
DppeSB2ztpAWk2GN2Vy1IszaPShIj11IugVNyBD3p6olru/UDMmCvv0zwyO7
ksvL8lk0vrYUCniH+MT+lLnHsUV/5swBXRLGfHrxbTZW4zbGoi/DeF8VduJG
5oiiad/zhJtFzU9MP2K4dia3MCaW+dqMey74eJ/pzmllOJfPWLcWDeJV4SKl
NkSR/vQrycxDj381eyvoU/3qdplJSWXTufdEH+f/jqQEJcDcQLcxbsCQIWPH
+h/Q1y2rexu4+CKmhpbVnzUe3j1ceT6K7Sd7+f71OnGCUKCg1FcUDdYPT/6S
wrbCvQ38QHPH1QtbeIAaMQtFTPNzZVJEnCUlBz7F25kBzG0WERdDpr8Ogbr5
5mLZs3ZhI9XrTNdugzZ1g57yERh9QCYIqSxg/KWZrI2S0Bw1iShhvTVggmM2
KbTjljS/YFUAr3vzDKT4+vZVyTavDzbd3TqMYrv4q1WVGV7i4McL97TqzGkL
xEBjNpspuMuSi6Lh82nX83pelu8XyopJvEGX0qsBpAoxL2xo9pJmpA1H6gWX
alvK0pqLa4rmsPgEEquntHyGqb4UQLMKV0h1tUOStIEFHq/Vh3NnFp7svSmh
qhWN6pgYkyUwrzQ1lF72IqA5JiqoEUt8mpURCiWk2lkiCMQmZVdm+R+HYWhi
S6R9OUDjvUSQyZf+KisRS3R4SGu4cZYuRZFucwmJiouXzmaMxFbsrHkgTwlu
jZwccMajWSrR41j2IP3BURugM7kxS5B1OzrZEuz4XtjERJHjrfX9A4fW/wXW
yEqVdydu4D/Clvy3r4rotJN8Rds97ddnSBZjGnH9N7FBvrsL/VkHib85iM1F
DEpmhXSZDRCmL9zzVOtBbbk+tSLqAuKHu+MV5ughQnjOE7GSEH31UwGZNcjY
QhWcYy900MfA5WZWaa39r6VnsGnEssk38GajXKPte1w8FaRlrXO7UPqFYdg8
KAs+f+wiQ/Rnkxh8D1jLWCJuobL2Ubz6RTOZodxR7JzTeY6o37ofQpBst1L/
4rVegt7bz975JC7I2kmpoMy6E2h/fSIJQY6C/Qc3ATelTDvDTh2Bh5w5A3YH
F/BHyUHr3yQfjNx/RcGzx+zSu8jTj2illdUsVhN9QJ6HlEPVGskg6kFo/5oe
zFw1XMrCb3zrVdgR7zdrf/hj5Cml2fikTn/J4rHjj6ixJj9gs3kQwBHQbpxx
UPvEBMB1eRSWchXGkd6O5n3Fo+y2EDwh4Q3AnUjV0jhAJ2D+pd3sw0d4U6ku
km7zoY4lIKRgvjb4lL8IuwMwbi/bmZTKaucdUKy8C43FhvdzJb0KSaIuq5hz
1m0jXJxIxhLRcZylIXIQXA/4O/XeZqvmywlTvrjSznAwJzw8e+z972y5CdF8
5FwPB5io1gpsI7XZ3jGOdlJlXJvgrrC/11kUVDbvs0yp5nLpiPMfTIWaGLqm
UmBLu4RnkhfR9f9lGfsLUpht4gMV9m2j7PBSHr1BSWGeGI2eWLR5Kq7bUrsP
CIminxKwJfRIllh2grUg0vl8rpWPCZB7p9rT2aW6tTMrKKHCoGEm56TMKaRy
yvnXaLkl8RHl1f/KIRARfiJSZcfLnIrIJro2KeP3huXb4/Cg1LaZduQrSiwh
Ecl9+T9sWIyyTjXVrCIvyqTQmPef+YBJsd5RiptZoX9mhH5rJPkUjIALkK00
xLRbsPaqQyd5n5imZ1Q1b9yjL73psF2zEfWbTsc03uf5oI4wc67C8XkXOp1E
LD701Xb/J0yfUc9DngEJs5zZNlKCTtLd8OYZs0JXaEoNMCFrV0If0x8DLE30
nkLLrU8o3eU3aGDu05mDEduosjpUGzaCZS8B2x2+zPTG2GU8hzPBOAB6+m97
Aod+VSr1YHr7g3JKeKJVmCTHisobPW9W3ImWTzBlrH/RDTYaOKvp+kTUudR0
0FN2m1USEQt5QhGURcAmGGw929Il+WW3P1Af0CCE4877BDpPxLeU+lUZAgN/
rgjv5aMRKzlym4KebEysBx2Ynoi0GH0Lk5RyjOqBrzJxPZ6JPp6LfZf9JpIJ
YcXUBpGkl2aZlArgSe9A5AUYmVFFcqChX8fCahdMMO6j8kACBNA8GufVG+xy
RmQShkD1hCbicRGmgWXU1X+Br+5/gMsUfNmozwkEwpnotjkuXAFZwqeWx0Mh
FyQfI8AcOU9faB3ELteveQeP85OLbdQIsJdYghHDSMbTwK/0DF1knORxio1K
OeOOs7CTayVUE5zNo2zPu6kmK2pjblOj6kjZcDZyY5vY1XOIWwrtxAdCagxN
UcA5htOvcXZjUZogvARRviMW53zE9BRFqi4OeyucGhUfsWrs13TnDdiAn6Br
HGxXEiQGqJQnv8P0u+M4T3pj7GjTj46zIqAdySbzd+b2C1W/SKDkFfDkxjJ6
oY7iHwX+h0adVmDl+f/nuIHxdE8WpaQGUs2tPzo8vVmha1hoJ2HmEgg16jzK
qfuIIQPwfqxXqLUtnZOutNxsJcRPwa5FKfF6Z+3CTApyF/VPailIfkqjYUiN
EmPnbzRx4W72TPXeTKFhBY7qF3CAE0oblh+midwO0VnbG3tzdQeCaYNB2ncS
Hhe980jsGtn0Kxero32sXp0I+XpPl0vO1ggO/oZTUkM/8UgOko+BFvx5WxFm
jQ7S1JkeqyTkYT8tmrS95hchsK25KP/U+aHkMpvz494/TvbkCRqUq9hyr36L
RMHeBNL3hAlSksxnv4bD3FEv9/qvAOw4mJRaukyOWYdwTAvQ7BOo5tExj+tC
l7xmVNy6ZkRCUSupSkxVyjadmDDwJ8o/nbnqyj/X3gq35LNs/OOXoq/cWoDT
xjUoIGVOplqThbFVAOt3Hggz+GpVmswO8OEyrtnbiS8nQfgombr8ZoiP5gDu
s3OeAvkNz8pM/WWhLcQ5obJtQXPEPC9a5aO61BU7tyGvBgLwYqrcAci7Awds
+xWuItVQKvF+y8ZNpgjp/aQVEJdNL4bnk/5btTjlvvx4+K+HluoN3fb4reUb
nTaiTN05dL9UraqCtSDaPDWvKZZIRtACJa1r0bNaft74vrqv/mXCVirk2wHL
YmujnoL0N18RepW390pFsmYIMU9zxTSBSoGMoDePjQ8z0Sj0jgPEjfiIclLH
ziiSLe40XNwC+wyk9uJCyu3tEJLOFqEwvBHkf6nmHU4TLZgi6mnTFN/VwWTH
3b4+k0rnJUEWdQueMTFR82rT9F0GH4rs9PWBHWkjtq8FLnvI5t/2Au7L5c9A
nUPngV59qk0fQFxvZLK8O9Rc0SxLlrIsPjbLIWZNVHJQ7X59wdAPdek+6Sdc
1qKXt36XYnhgzCO9ROWyYLrxz1Ay7g9WaFrIGLyhh232ZVkyOg0pF7niglHP
hKss1xIBd+DtbL9r33nXpU1vRm0bncSfy05fnKnIGDb/3bZiYN1XbhknOaxJ
nQrceurnMI8bVVZooihLUCQ/2pqwPJY4J8OhyItNaFdhjAMS8NRxbd2/QRdT
0Xjd34dBu3Qi9RC/bWhPbcG0aN+9OTWnFnsaE+yruF2+FgSYBprNmO8o8sTo
uqQOj7lvSA2UuUqFKumIwEiVitBvx7kO8+nL6bA4hbglACZljmpJ2Rrasl+B
0/e8k03wYw2z6i8WjHXWdyrwunTPetF91WyGjeboqP85hQoDso2FzdImeZDv
GtuhqKUaM/jpznizj4BJfXQ+2bK0IAKVH5bRy/pgtOFqzht0huGEwrXrhIhm
nreHl+q4y0XSh65X4I7UIuxZaBS9SHWJmCVsMV1XLwowWpoMR83kj08A0t79
jg4x7is021+1EAl7YEvnHjn0AdzHIo6Nxg1Ux11yj1dBr67DOr5P7Y5kmHxn
HneSEUb1GCo/FrsbN21/hfSdmgeh2IVW8q2DavzscyxM7sCPdoYL+K6zjoQ4
zB+J0K/z/z97VtAOa5S99QBPrzuqDGB2jEW+R43VUg3Jv2/W+4q0K7CenZsY
0XApq8ub/T3DeYmCgK5VRe1l3xCo5E4TQAbqDGpEq6G6lsm65TkjHDx8QX7j
5GatVKr7haHMZZtyCyhreIkY2nirlHIqzw5iZ4xWo4KHMk9WlSDX+JJFNlH+
YCpcHGBxvdyKxpMoVWHZ1iI1HGB+wA+kUrsHkQuzfxAs8SNX9A0IzX1F5cDY
A31XmN9YqoUQDXIcfcZO5mMZQK9bmGpknd/PyHJ2Od3N71GWtCyEXho0dGL6
5bDjztqBnuxGxF+ccTvGCFJwlRnySAiCtMRZ6MNkFq4zUB7jSZ25qJ1cQTMx
RVQk4hcxXFFwqj1xmtPnlQ+hv13jzynrmloizAzfYGkuAfjwnl3jfz7W423s
WDRkMG7pn9cTqwHoHTteyybwGFV4kYnxXag0TBBN8Lz/CC/Vqn9H3UuyxvP3
QceOZLum2ruB52i0X5ryqO81TTaTlBLMb9D6tu5WCjes8+HqQ7TYkc58pces
DY5V+sW05pSGTwV9TOhM2+VjyqFDUoS2zKJCxRxO9dcCYneomaKQW4UatTSm
QZs5ZUzbrFqtzzW+6OHn+93qrh+wnrjEip3Z7kq4IcPkAIlJihvdDR4iXQRL
GvnUGnecSkcOOUAvzprpd/7RTvaveGGQKWL8y4qaYtALx0UcCr4yy8CSBCXc
iQur1fhX/a1uZ5crfPi8y4qaR/582v+JpTNnZ58JB/Cy1hoFA1dNof3ZPBQ4
hKzeAXZ3kkj7B7+7sBgt4XqEInxRuv9Na4AhrfpQS3+s0pEjhU2IXrGxg+Pq
xI2ppMGwYd9X4IBqjMlYdVEzj76HVA6sVuLjNbwa9gS5YN43lmzRf52U0ttP
PKvpmbT35cqAbR2hyMPYBHgBmIhT2xauXaFrH1oH3L7rhw3y8zcBywnjJyi/
dC5fXTERwDnaFuAVKncVlEAvJNIqIQwzSxhalhcJBt7g6bgfEqe96MmC6lOC
RNtczUfQRVYMSfK+d/vFwTygRVd8S0bV+/sMCx4/2jzYAJ6VR8J+qKi5XOjo
sXuuZkrtlPDyZ8Yms+pHKM1dbQsw1kXVWYsbJTq8lDqQiuwAautMg3ezd2JU
FRETir0K++VmXq6/zNyxoXsItXRrmB/cPLILx1AKNCDxMH4TrhQ0jWiQ0qKw
HW58lI9ky7Ai86LAFuZKQy7GjzA6WH9jbhwHbiWCSC3+CuBcg/ZGsaNXLTRE
Qzx60R/PSCuRlJpedMl0aWeru/4TiRgoZ+8BI5ZsS1tDClp0fiVwCI89dnHb
WtfWXxtGnchX/zVXDSKyKYs3yuWv7LojKEoQaxP1QeHdvGnmTNEMkOIkIUji
1LCGSqLdQyfzqI3TceAupKm0nKutnj5vViETwmm+6wR8+3f5Tw6QNfv94ZjC
HeE2roi0CO/OTNi2jJcnsFWyUjdSIdmj3kbI9Yx/LNiybFemrejY8qj5iqk3
AqsU0G3tnts6jphdXQVBrlBz1k+7MqLgAg8E1tlBk1m84MmjFHKsXJLJB/JV
fZtCyQb52kiDrpnXqD/IwAmNdB29fRHuElGkPOPyAIByvY3WaHYI3kgCuNbD
CvN4je4eY8noTrJLWRg8GofN0n5bURcnWAZUjQjOYiyoRtaC+fli9YOKiJWC
oNCPAqv1Ah7SONYH23HuPpY7ehNIosT2hdha2uOBSoX8FJfBt7Ze83YMej97
l06IuuldyL6DlvdFpB9gVyLjlWfjQv3PJC9SaevKEuF3pvVqPh+F7Jy5QCCn
Utl2mTa8dPOk7tUZcKORlCQmCd3MT9pD+Cdtjbi0rGqtG8WXhYyP8v1PXLQB
firRh/gThYYEv+gHFHOo7M1sfCoLSyPisCeBxmvzkopKQW2y3y/irLn+E9eK
cZ3AGkjgROi+jYQf7zDd15DkvIFwEYM/+S2MYhmnE/5Tanz9WDN3NMkApq7r
cDTfE/ixvXrTFDvBBDEGH2JVuS7I4jVYjPLlNgVzMdjoxAtYWzWqGgoRa3Eu
+Plrf/EdF4XQBB/9UDFy2OE8/BA/E0AkSvsXQWwrkxSZMbPpZQ7PpIezJLLx
OBtBb6t/DlpVfDkI8MLrhALilHujI7nmZjscMNqG3AjOt199f+ECFBNhFpQ5
TZ5qfVDuPrlPQcJ/SbgpiguUKfQriztA8qtsiH4fRNtXZna/c4+201okMkDm
wGEpTTZB/uFEse/yZ8I/fOcnx/IweXLjSMxy4Qvs8+5a9p3AB3wc1IO6lPWK
ivECH/Ad+p2j8ciXi3g36RHtR44bn8YmC5ke0AmCjwgO1KFVt9u3cptCsIbQ
uCOUTvNNhudHjxZ3aJ6DywITJ1Zzu1Qf7MHeK534JHHzpUHDQoT1vsGdtXs7
CE/70+QSYKWk8VXQsCap9l0CfSwDVM9p1G5tW2k6Eoqf7MSuorqoI6gH0FZc
loC5PdM9CP5C5aPryrMTvZ0K/hekps3OLAA+nOTMQnz9lHtOpBHbJIP7lr+M
/67SZRwjjVixDl+Ka+T06Noq8g6ddOKrgVeDB/CM0Jv7rO28z3TSo1E1sjU/
yzodnOikM78MXiI7zPG38t4MaiYzgSyDMErfPkIUPX8gmcldpxWNMRISnkxa
gSBiNC8z6CfEwxYEsh6ei/SdHGNDQLedK10nXH0NwsZaLe8uMNR4P5axfhp/
mgi4Pj11CF9tn/nN31r68RG44VPg2r1TAcDFljl1AfRpZOFii7q5Vp4pMRRl
tiDjGIRQNC0Rhu0T6E4ebIpAOy+usZbtSMV4FoZPpVb6FjPyAL5UKvJf/tSX
Nb9iol7KgQiWExmXpPRM6CTCYG+xc9H8krESWTg3Bm4Mr+5bKFPHFvVzRUFE
UkBNcaNgO6BJmZVgcbHgFfKpOZXBleX4xVKtG/gVCUgqYnrcZX+yTLhVntYo
TPOYOW5eptcnZEH8EvMKTBu2NgnuCoalGK1AyT/QKgNjagxrepaL2i/tjKiH
+Iq4E/QByA9p2d7whvV5L2sTRoykWZIVMsutFtnyGr8kaGbHisTK9eoPMXaT
Lw89o7c4qKd1t3/LflRUL9wqqloeSxkLMLb9aElKTrMRyKjrOfvi3l0jzoq+
sdDIo7sxpI0wLsFWthrRFF3c7NcuearltQ8r43UY0BP4CeEOTRssLj9VP3Hg
26RVf1iApyLaPReOiKiU352w+kyMfB4nQ4T9qW4ClTV7Z9ytckZ/zaQIVo1v
iyZAjVfKmyKpS+EazDXtbB1dEna0Sphqo2FCBF76pEoAqYP/ax5dVqj2Pz9P
5K1/Xu4+3DOnzGHUrVnPNS8XhT6GUjxeGQ2vPO/stH2649VgMBSPL4Eo0BeY
s5NS0dy2XjdPJrukFZVhVdbh4J7wbrwxWbD7k2EBeH0D6HfsXPMAyYP3qBsJ
HfkJlB3IcwrRKXq1V2Rpd6PqipjVxgBRCZ+ba7GO7tzOfiUd33AL5+WXBQDj
e4cF7w3cxchbUcoQyeLm1wWnAXdMFno75hwEWEJ0kGUuscExAuPbiXeSAQi+
XEZBiBbWLUsMw07mlNls+zeC+4lLmxLQyVBzT1A7wATv9PPs/bmM+c/zHCGI
TPb+DB5guyPzguURTxz9I3Px988NqxafMLV39FShEHKaJDDj4unf4+KuP9ka
Y9YezgCzFeJhU+diG4f2DxA0lYSB6q3okE9Nb3l8BkTOzu8LsW9HKgOJnsPs
23Xvogms2sz3jbdCk2ITWe6x8lamYJixXFqY6mTzs+7ZEBteUHij039T3ovk
l40+PBspymaTKvIgQrAtUB95jez7dgZ/7xdkvb8cRl3MFfrliSRhV1Pk8wTP
XT8Wz/HhjTXIyJpdwTFGjOtNEZ7DxJtO4xsfINMRMoyd/tZ+xrQeB20U8lro
1Jv59t4atD4rFGpZNjYkNkU3EoI/OvUFy79G5LNtOOfuMz6QPGmeoKDNNLQt
xaJDxEWQuyW8k0ftp9w2zNLR5+MEt/S6IfhCfFe0WOLRSIU3S1qIEgmYByj5
2PR6Er8j/X+TeMpLBT4VEpiQu2i+jTR5LWZ5t1FQOrVvt4vcPcfIraVjfeSQ
LyB5dqhfdn4r0omflQCR9aYufNYHKHkFYjm/XVpqUqC5lW5FTsiCdTjVfzzM
vxCHrO5OzmoEm+m/tV3+svUVyg+TAfVW+5IzjtdJSj4WBM2zELRz1wmUOIAI
DrWEG89SvHOKmEA5hW39/Cgf0cVOLnBhCIgV1kz84UOl+yVRj5FsY870VKbQ
rPKQj9fg5278r5mXnWmA5LafCW0K3BJaP7PWcNPxvKIlrU7aWjn/T8ExjK7n
q3kwh7Rb4k8+LKpChOFwXFrrk6QYu3hj6DHAfamYbvlQFfFrBRGXsf9EoKUk
a+UYiVmw2FY2Ykxcb/SJOGm2wkfIip6ZNWCfahG25bCPbUkeuIz7YuC12wBx
eVSaYVPYJEu2S2XVT/R1ye5Q541znGLI50Jy6hO7HbroUt7+TX3GR+MXxFhk
w5SOzZl3pI5KXomfPTo8s57IPu2PM+agJFrvzIgBFNh4DRjhFckdFW94AlDl
vhpEyH2VZFmj1EIAu001uVZicoaz8+L2sLtJs3wG9kUfO9ZofTEOU7+hjsHs
OstXy7VGh2+xFHzYzpWLFmdRJTGFCYNmWDAqbTVog/rqkDTU/IDOixzMAHIB
4ucj/lwijVgvWI+KI5N1qAYdIwkghP29BSfqTAmx1+wbfv2A+fUszwhOoZ3z
SU0QofOMeT0bit4kPgVTI98AUWqM6y8D7ylzFPT2XEW+rjblKXcVDEkMat+i
WHe2WePbFpvGAcriWeaJxbICelSyBkSkcM5dGJU1xUNNo+NUwEs+HIuXZjWp
MafmgrmcY2IjjGF5l475/k+IsBSztQ3w3tBH1yAxSzcdMuGxFrzFUQiwrEFq
ePUqOt8W9k8LejfYOSRFkNzmJhK6wato4qj4RTlbJ3R7ued+BvsEi4NqTOCq
jvwk0XNyeg3T9WOv4I0IRbYVgzau9xIWjk43RZBOCLdOoO1xCqBsKlRNoJLy
DycOONrhlSqKO512m4UWRdpNvcKJPD03iunE9C/k6JnXh4e1K/N61WjxJYnh
iA6Sg/RY5exALOGNZ47Fy+7EXRaNSQlgnuEvKb5z83+9BMFoToMalV/XgvK+
k+zpnFfA0nrBTFZww3Iv2pZf1yYScSLDfLSc9qj8y0lPCVxDhBkCgqGOkEdb
mknJyh8I0EG/ID1/GyV2Rx+PFfxTfPeLYRt5My0qE6+ZxMesC4WheClk/vLj
tyOdhlXoe4epwcUYbG1CGYOHl4uUubCkXpXsXByS40H7YCR/vQ0Ys8DiIk7J
hd690QrH4mT/pAMDK7BpVHcby+QOxbDTkfPThyC/oPZXN7MIb3isuSgDATa/
x4I+E/jwgGDDFkQkl6SJ9bO2GULqFeVutmrJQMagx7jmO7OSxthUegkB+hWA
RSQxzqmp+kLouPZzHRbrEMcjqxNxvGmUsQbTUH45WETzkycDcjYwb+hUM6Sw
xToeIUOB73ozPB6R+tCYEpKbBBCgu7Zr9j2oZKkLEV/Q8pxvUJfkeat8Qjsw
trcTApbNKQfw3/DQeS7e6xtnXYfHtl9jq3s64EEkMS6Wly7D+nO5u2LoBJsG
SqwGIqduuALramBVLBYj3uDMI4y4K6cTY2J6P/PJGua2DJXobPzdkdrpiFXd
zGsrTG5TJnpKzRZ9kp+GE3b2dSuLW+O5oHf91Y38nz/cNHZJgw9JrlFwOJ29
ht7uyqEq1C19Mocn68yrqCHbDOXtouXH3BmA1wNnYB/HZuHhrUjJa5+9yeHS
d9vhg/ivk/xB/QYkkAie04KFjYbtlx01WGnl9maFqcaFtm2G1Y6vkxqP5HMz
9pdmNY0dSh4B3M+OpNEmz0qKRuBUZVqnFvJB6+Kjt3HBr3oGVumg7XtWQjJb
8cE6V6NPqrPfORPe7ztI4ARqtLb5SerTixfDFz5z8CL5nccW9rekEz6zeStX
INPUywXrJG7L8G7ZLtTFTMkNkbu9uw5vZE4PHikeOYPJj2yB2nRjDxBDdpdW
pGXV31XH6w1MaLNFmIgZRMtKsst30eck3f0gH7yYctI12do8W4OAsY1fvjFc
L4tgFVd5d30kD2EDijqt54x3qYxeYyl50H1VAee2f5WNZ2L3+nTxu5lXLWIj
Dlz/QRA1bYzpREudwB0VU0xM02qyiFyYFQq2ToLeUVIb+XePd1+J6lnTfEPE
Ewx/zXVcZjl9YxM30k0xKnD/lUFTPUKVavAQAX9lEBAbvGVxYiW6ySwp8PA+
o25fZdnroxtT6GV/qVqEruQfMfAqwyN6SQMbRPrcGfTVMeSt7q03gPvR3Ytr
GvKUzl9sTLLO9kxR2kcBoBeJ3yFmPF+yf5Xg43Ih4LLCuc9SgZItMBPN5pnn
sxCZRIry8ecGqqKo8yaHAXZ9NfSIQKHPMTYW3R/J5Z2W+LBDGo2PsekcqXHs
laoSmdhKHz6n5tMzgLkbNQPDhrIJLcbHeq9y+wC3vG0p6Eb7oZj1fDoqDJ1I
DrU+fgScsFC+XCVA5DXAp8ZPB+7hV1tInDbwr/SNEGJ92G1gHXUX2bUz80jV
Rrio8LvNv0fO+FjfUvGwxDPkAGCsLJz0UNpV7fBe4JmidcH0IbMFWWIIaHRk
M2lzrqjiCr87stIjbe0Fo/Eif2F4TdkBQM1EptzWM6qeEOYzdU2UtflvyC65
aFJI0f+OPdomHVKcN4j61PbtWy1s+l1zJMnu7throqeYaFB6CYxxlL6wb0Gd
6yLAeVGPIraQKUi+GWVCHl499n6/FXqFNE2/c/R/xrrGwwPD/2P7gmA5TlQ6
F6ViZwtAoWwTN1gNLCUlxSENR04yOObzaWaIedpmOL/B1pYgoxSzbrDuSwU6
vgFx9YslTPjNhBUVSSd8Z827cR1YKfMHzodMt86/jewHXdiztXO0Tm+pua1v
iKFrhPzUL8pvJRBI3Aqdsyx4mvaDqfnkwFngFz9cLfJHtA9/haR9VefDBfR5
UQw43j3TzpGLQ7LrR2aYZC7hWbW7kSsfUAaOadFXIQ8R7+WEfz8RhAFJcFUF
T1BLf6fX4e3bU9nsZc4uOSl1Uw1MigO93BjJfz0ctA/vcpt1bc3SD47qu7Xi
BERFPpoMugqd6/UzNyiTH3DhFI/8kCl1bLCWzWly13Z3WCUxRuTZeF+iR6ym
lxtNc0J7U2nXq+DKa3p7AiOVAiTaZQ3F+4i/LdYr0W5HQPIv1NcsjyOQNZZ0
x6aSaGIbtCy4mQuXKg7h5CIo9h8KoZwKrWK5BJkmPZoO7dG+rgIty4ngIRB0
hixtNjvjBz56tiMrpUDedEWdsuIbv1peqD486vktBA/+gHu6qpKjUJpRP8cX
2b1DQKqOxMLJFitu9ugMurcYPP+jJKEARJn4VEyNL1PW0cqZyKIagibXBSHd
H6GuhV8lVuLB6SpFOCSkAyj9hbSUGVpay3ovgLggwm1PB65ecD4w9cCukeFz
yzRzdcK88khkeYxQMVuMOhtflBG/S7DWAK1eDPSuFaKfKyeup3kIS6HLE5Ko
AOA06WC6b+67vbjjNbwasrQSVfoOP7oD3iOB7wRCPmcM1f0vrEqPdBHvM9Sr
MMce2cFO+a7c92B6oCNarMugC7ESdjpbIE8O6B2Ke9VKsht4zHYosMT3RRkv
4Y0BdX4Du8vGPKvyow0NPn0gt1uMJCazGVbuMe1qBpKGxfZPrWFDTzJFblIJ
PEFDd96U+Af6jN4bJMee0L42uPCQxqmSwupa1qvR0ea0C3I7v2XqGq8jbX/z
NLvG3ZgJQXiJ0k6Lo00Rmo4GU/73nnp8s6GeuhjohirqjdKOhSkpG7Q7tqbt
Cm4KgLRiiwOCA9GelRdzTWbPxrORP++0NB2UQCksAAAO1JnS5qb5+rPkTSHY
3X5b8WsPg8SrdJ3wgxBNy1aUtxipFkiYPnSfqQKQUaukS4019pW7QFmGENTK
aAZA9deNeNxFfa77GxPAzN6B5Z+MjXsmsjmXhHHVtNsKRvWofG7DW0XpE1y8
fChaDIhJG609HSVLCOHa/WyM1t5dlQnMr2jHSwd3wtMznXhnCLRjmNCyb5HW
X2LbueyL5jdpn6xr/mtSLeAwCl/9tIdCIbPAkIIgZNFrdkF0nkyQapethTaB
5fn81c8rzIeZ3GWsLO4FTVSsMmiiNFw98kS45Hgs8c8UyttQj7TYyiE7mbA4
UK0APdLb08fIIeVVK6LopMIEcVA1xQKRDmWrRIKsuafI4TVwYbpBIA99x02o
xduFvL4yXVXteneQBf8Y8CeiMgRbiWJ471fdnDBwNZgRrlpGcSZ3TiLS2X3c
AF2PvdfLSq2MIXxrOx/U1/H3O4zX7xhuhldzBAId7FE7BKDSXMlPO6rr0BO3
k2Czqxn6bVlLUbWiRlMpEfoTbh/xG6nbnAGfSJucYigoML0fUeiwN3CN2o0Q
Qlsc77/hmTw/elGbnPqLfhwIoYOb6U3fVhJxDk/+rj2oDmAbsZMJ9neqCx45
zTUyslTJrTHJzuM0DLws4ZOr7OMLa6X+7r/jlMZrBSJj42ycTKXNCW+zacCs
2Q2ryPY60+2RGP68rT8Z//Eg5tzAqEuT8tt/YMijVSQa6i1xsc04+D2hnrGr
2AW4I29XtqKM1PLy0alc1ONykZsfj7i0GFyu9AOHf/B8jeaeJhBnMnry+nHv
1SCTbL9ybu+Ko4mUie8HwN0q4BOpJ0ysoS0SJgGi7P9q5I0XIrXcHtW4j3FE
4KNTsOUf5o9F+VYACOrFphUf39UWpO0E/M8ybxQ8S8pNzaJOBndzp5u2OOrD
Ffk3/O3daCm3T+i5qNb9fi/0DtPasKD5txT8U+MyCE1Yhe8JoNMk8ymtOQHc
WsYP3be4OB+tiJCV0Tc0BWdCMiBPN3BEmNasRDsRxNMiCEk8gViQdUIBBhnh
cirH9b9jgxgjZ0G9N5Vaf9IQHmYnLkrRvCjXYeZK2RRhHAbji8QGgP7gF1RV
4mYkZJTeEeVyphboX46gIOrwTa/PwuyWdtZbkWvv58/mVikTLrhzbfzK2n8f
JCt5kMod3KPUzblrrFN4jYAWxNQKCM54klOeAIOvzIWFpOsyafYiebGyrMlC
I9N+X6ZcLvaOpXv+9e8xwhJubnLkN0ooXpDdqyW2v3h/kKdRxHOv+LUbhDe1
S4OFdcIJq62QqFpX1ousgYd7Z7fOHNBLraBbwxoYMrsSfehOq/k6dw/Cm3y5
RGiKt3IaB88EgQda/H0UtwMT9uNIf3AA7XzciOxunLVbN8aX1z+/cOIvTvwI
dDMf244WLS29gGUR3hb9/NU/fBT0m5m+YgngBQAenPTdk/ZIAyE6bDdBAduW
vTC/CR3v/zxc+c0O55QQXbxVSDWe4Ljp9wY7Ijv8i0uloIG03fuLIx7xnE0S
4UcGxoNP24aBzWfV4sWgVlLWDlTNfd1Tc+UMmO3emjTFi0wlAQbqw1SlKBE6
ml59C7vYWLqUmqojYYLuF/OC43cp+SHWjhwGYWO2sFI14QajIwwanc58+2rb
oul1TUe/umrOMheWv66S8e2bzea6PhtlccuAk5NW24GQnGogNWLHyUNIEwG3
i1/jOpiou+PDFMYKocGv3YiLSmt523UGwMDsBIpOh6CH20zIzz0qRF5ZZRGV
UBJxIGRCk7KPfDC9bYY4QDwSfYnccMOuwlJ4hzq6xkobPhUcElzAzJzk5KrH
0zPRxUEfLApR1T+nTr+mSkuMEMINkkde1z2n3oEccEdVsIaBVMoe5TiNulpL
BqRzjdaKackMvkk6Kr7HfIZ0ECegChBKI8FfUYw+/YdYbIL5VIduDJC0dRYy
G3+2CksDULssqK1JHcmXL/xFFXLPG3JGuRQAMFRfUQtp3q+msaq04U5GMDMm
JGUOgVdrOaPhxpzeq575ivALQzB0M4MNuTkWxI8x1Sxq7Ld5B8CP+9bZ+xtV
MovGncOpG5cQBQD/J6EGLVdf7wlcXRaZGop4o/nNQnfNLDOTNTl7VBlhPcYO
EMjyj+WEvR70N9lXAtjNLK0/x0/PpfSNhTWnbrVktKLy8A1vsnwg30fCtN+B
240RO0huwflGQ/+Ya/beSjeUUTylW7jY1kWLdDDvBRTk2IHD59R/DjfQkvZ6
UlZIN+zRFINu/OEh3evPs871Z++AMERTY9I5mv5f4MMtGwPFUk9WJ17qmPgi
xSHIkxhsHjNdP3wUl+hHoHwlDQzvoMomE9VCv8iJFSpJH3bCsYENBjUxC5Or
RhOpRvDXKMZ32x/qKsO4lq3b+supf3xuGm2eJS1aF81glP41TeaRNJTyn7D+
GgSSb7Qgx/w0aXHbKY3xrvskRU9bmzgONQfBLR6mBrEVKcbmxHv7xDYSkRE8
kWqxYxlIWicQt9WHzRgso2ApOZBIwuyXOsfk93olc6d+mL45bavMIP2+x6lO
29madUVhm/mGni/ZyWzGazoTqcLTMLiQ9U9VibKrPSOHoOW+NhMzmqnl+O/G
Nu57SGZ6TLAyGxLBwPMUnJrn2Okdp6RE4+OuzmQyVpt1bCPohCb9hecFkNzL
XM8vN0po9DYm/QnrholOG11gW3Z72Q/d3uKByU/G8XR2TBbvZ6k1Zr6bLNhI
Arz2RQuGAeU5ob06BQ5ADVkZ4zECxD2IPSEiy5/xFEQ+VlVFojkRyiKgNv4C
XToQ66dO6qxPZz9zG8DII8RZw604ThUulpeNkb6JLIQfV1o6YlYjr0Wahcis
V8i+ksviOROcbwjCybdeQj8XO7B+nLat6NE6gVeHuLvf6qEjatHuJ9KgdDSe
HGJOT8rV11OsMg3xISfZxKKMc5JD+d4A1D8Ggwc17OpZUDMpQ0xRzoWO1eJp
wn7t6qQpGLYVdW9Ht7cUTD4XZ6+1+XINJgxHOlWHbW5x6pJt9qCohpHUIRS9
MuOeITNncxZ1LO7yD368qHv2lHL2TwGgc2y64KXAXOnp0UZzOHhcNutFPNMX
fpfKGsw6PTkargp9FDCWCphEml5Xnr2A1wqZmp0lVKvkEGtaw5YP28CfEiWp
PycYl0NZuA2JDohErG17O+wxhYy8FsN3EHBmSMFaM23hF3DxMW2eSmPuGO+y
Tsq+Fsyf+aZIffU8fm0iL0emu+mL12WJewsQNXdsLMBoYApwba30YErpdTVH
MG4ufz8S45ibt8AZ5FicPScXD2aRApPtu2CYHUhmWCgHR9CvdKDeZiAIHIl7
E8UdtW6g6pre9IN5UEyOnawGcuMn7b6ACiWbyPZgWnMjNhqW9o27PU1spUk8
uD1cLhRfDKSLHr+BzA09fA0u4/xD4JrWCuOVst9wmbaz/dS2o5wyeWF8+pfT
BWgs5qrbNQGPLSKs/Sji2F83IPLakPoTKaeYrftOmtzBBlUFzFCP2eLFUg9Z
wOMm5bl/i+lzDNTsAX+JiqQxEZiPpbPd/rfzGaLYafgNXZ0bhpogigXmQFMF
lggrv3fKVm7jeToAGm6yPnsson6wcU5pHhdmVv0h7+7g4nrmhuzjVu9rRrTh
9ivR0uN1KoBMl0PzKz1oHNbeuCioL/M8WKo+7h3Re/AgXzJXl9Hu4y70oB5j
7FChUmD/505aeS9iTI672FBLW/CRGi3X9Mhub+QqQVHTmBQ3exHDZZSErTlx
roVWyerqzRoIsA07Ge4mGmBK0iPsm9c38FNoR4rd0FithbsTkPs6FuHQaLUp
kj3mt6NaYLwlMxgKHxjVdn2iCLJqqsW9FWO0Jv05/Tid59UFgPrGXP8fCkxE
XPZQ/CS1UpBbk2WaSdi1KshAO5WJL5p5TWhIfZeIeXgzhnz0LWlvfaAdCs2A
dJkFVhncYGYm/HZAbYywYi/Nx5Z9DzddFMB0+bgN7gufH078N1OShfIXGbTP
OpcYzzihT1YK4CvJrkKbm8Y2nY7ZzRd/J2V0go0bcXPr7WhCWsEHwl/OZpO8
13fzp1AWJjLXZ7SLrzvf/tFu9hViqgu4dLmEvEombyf9sfKoTYSoxRNKslgO
7kDrgJ6+L+2B/4V88RPWrprsVbsfda9Bzgd1Zt7pqpM4+sVRViaOfLGsA1wV
xwJLBf4s73u4n3etDroj9D+Y4WltJg3E3guaw6XfUxi+hgfUjRJybBS7pZ+f
N5KP+l2JAm4US8dG92u0IaR8OZ2izmz2ZML3IBGVXm/vPxBhgz1/PoS3s6hv
H6Tqyxa8UQHMaV6DiVstRhOcr62s+h0v2pLj+/EsZKOKx6eYT4N5ygYMn3am
p+arX5aLBXKckbRNUyPPc1DhtIdL1Olo8xKu/PKJfsMxaUWaMC4xipZqwQYY
/eWKulcElnVbxvRD/4uE0J0bcfFoRdaSXOAnEPOvyBoXZbfudgv4CtkEjwt0
FRGXURGFlR1sKf+5BGB0Wp9Fra0raCaso7WoTjTN1kOdP6rWPhlXFP1pzhnk
fjLHPnmDYuxq/v8NWi2LWI0qzs74f0x6lbP0Po5upUHZCTJQ5KDm2BGUt12i
8nab2fn2AZG7QzhUc5tghxmvTQTBneaNl7D8eV+CsqpnJeDPJenRpA6FPA4N
3lK2jPlZ0OfbWHxYEXVebXEWVq0wtd2hcGniv4XkiyhlzeNuNeqq+XK3iiy9
ERczFo3gNf7SC/SnWcck4i0k472QoKgzCjPMxv6pHMOWM+0VOooEKVhY3L5r
HhYjwyDJzZGwP3EfabIJUmU2SLncB2fwvJ8It2DrsP6fDzWWqda3yYSD0SSv
SVZEWT11eRdwn4MIN5FnhduwGjF2VC0dmcA1XeSa0oQ9P7LU0pOFvqA61ApM
asDr3zjHAESNRq8jGOIEFHPHsr9nXSGKFAIKZj2g9vZEahjlSaD5y37Kea1J
1D1WU7YmTDeSFKrma2ng+3lrbhnyXgyVqgzfMFq47/0hf0C6z32dB4y9Y66K
fN6wr5azWA28QyWcX5m8JVfmpna0lCLAI+bn1ZbOezXfCIynokuLW69Y7C6b
MvKTw30ncBqdLJzDGFGKpKdO1P0uc76HQB3pi/YGYvVqdSV3vIuI1Kk78r7w
oKpfrBcEu4Ocmu0O8CbpI0I8AiMukGWQ//qYCac+YLEQDP+x+M5BdCMJUTRd
w/a5M7mEVk+9ZBimA7JLCVAFc4eXIBqMGGaC0iS7arXAahH6pZ6oIk95Y0/k
K6Upx7B2B4gQ1BjIS3FVzoViSedNyf43fnL6+IvSCo7xTL2qam+sr8heQZTP
aPSPSekps+SncewEPzbuEaij33dya9E7ycprGxL5dmxkDdVrLMSXRZKJAoxb
fZNWf2wZjs7aniswczinMPyIwwwNqqi/fwDaYWapWbaZ0BwQVmKbiumHykNi
J+hXJ5lkzaknzTULcGAgrTp2C/NjSJERvFyuKgW3jsGZyoRtda2WGhUQ8LiM
mUG0/XfN+nuAYNfGkp2+G1kx/thiB9gA2RN3bSgsGowjZj70enEuyU6w3pMF
+cUbOEyGWRxCbioHkSUOXLRWWWSdfDOpfK+XsgNafMqb7OCqMLH8lmEV01aN
VmuxRSML/Ng/AOTl54XeUc39NgjFQdqBqpoPl5lM0YAefuDjxIUMOGyjnnvD
zM37DOhrVQyQ8SdKbKWSQPqhILZ9JUWWNNMWbY8sfgA1WsvU+iymYHcnu0bj
cZ8s8+yLWOuYzt7HVTMKh52UqdjymNLw8ZAnbAZ79xzISyZ/P3BFT1JKuZKB
9r0VlYgdiUnL2WnvAMbNy07Dx28dexTKCKSD4nSft3zZreBm89o0QAoNVsjf
yQwm/9lSIFFeJTF5mctRKQEqckmvTO/NuzHK3XH31DfoBqxIJgJWxxY4l+lA
YFyYrvBXpnShg/98XbUm8InqMAJbyZRedDvy05JVa/sQtsEHXz6qyTAIMeE0
dk6RbH/sEmFDQ0xvH/O7r5ZQnCHfSq9PdxAE6vOldyPn1zYB87OxgOUoHGT3
s5z1LvyIIP4eB7DRcKwXP0CEFJvXbFe0jdkzVr1uTdsGiNdIyX9tnPb6WdTT
qkYXDJhuPveeCrVvrQO/b7kF8R+y/a2Vn95c0DckyCZ8gfg+s7UGB3KXGNKj
V8vtJoIx9y+xLP6KkmoyQqMG/W/uc/c/Rz4TCd8hioSJ9/kyIyGaId3wCs1r
JNh6WYjBMAsj/Zdy5saxdcXMl+yaD1098kNw2/c30YtfB/hXMcNu27fecjLW
/+jhGxThrMV4aEdr0sxct7MPo/NmYOv82/lP+XhWFn4Guha2uOOEN+G0Yq94
GWaZYkLsvNRLOB/cf4beayUYaiuCeVOp8dbh9w3yaDz56DeVD9l9ioAxajRz
aXkgwOyzntZV2sy+lndlp2A4Ig0bWEbhI6Z/PdekTlbPO8bblzkAntXGJn37
T5vuDUFzSqfIabkrwMJEje5cOyWBoCvSR0Hn9GzKachSRx8+s6Yve6soKNTt
o1ef54ykCGiFFhrCS5SmCKHw0/y6fIYUbL3R7082k1UKNS0735pM4Xp/nowS
86Rja8ztHcXVY82mISZ5boeHDyfObuCdHs+TQu/0kaTrwkCt/DhzxXlXhJiL
+QfIsOmeNqy9Do8cpiorZ3ZfvEANLWneTKADrgdBa6cyc7vWYwchOMtATb0P
z316QM4gsb0WTHWpfdnXdvBxdts37sK10/mSE+vEJ38eRRJpo9jNa8urRobS
cm1bC9KlnIzTN1bQXFMTnbMCjSdtHWsre7c/sjtouaCOtsE3pIaxIsAzcZ+/
EIhAX8O/r7vvfjO4uuYpaljts03VYwPXJLVwDvlZeiVjqt6F+xb4BNiOMQKc
CUacRWKJOvb3Ea/2QUxEXXdmL/ZDflMyMktvZnNZwXy0iyJ6BWvSzALX5TuW
eKuxNqNJDFoXCtq6N0Ii55HngTXtd47rl3iJhTpJuf9zGgRbOAzRdQN55wiK
bCojlho2aj5E12W3DcRpJNWSunOmr4B4MhTqXrpD1ZeUo/P+KFQnxN+6LcVF
LPnNYwUC73VnefCo6rbQwlsGywI2DNqxobdomltppor2Htf/iGlVgFWw6IBV
ZDIVSrBpzauSLTz1czltZppc6JZ/rIK4a94wm3WOFRWDGXjjIbvMecCs/vnz
zMIZs3M7uxp3pq4oQHvXIRAh8GQ4Jg9pc/gEpJfuxFxgERzr6D49oY4OOYVz
fWtOLzGV/9ZETxPYoTkAmFFWSNk0fs/PAq4A05n2lsIc+aV9GvnR+bTj9TRr
WV4kdVyJU7rB/a3NuffBsVDYuv+G2qKeulUiUuZ2NWPFfqBuqipf3AEufBEq
bx6+l8RIjtfdzgFjQcvAyPQPQG7hwRndcxcfxazAv2maFZPwnv1e1GMXW3v1
145LYZTqO9tt4Uvcn1SGs5NcOCqHAZ+NHOx143CnvvWTMG4TXg7pO5F3r9SA
YdMTQ2cUpQfZh/avW5zYyNIY3TOGqDEbrfyI4Y2tw28J/4Su00w0LJZ7dt0s
SX4GPYOzJXV2dsVcW/tOrNocILWYDYZ6qwHnp5UV4mr7jHXoCfy9CG/64VC2
simVgwlYEeB5QK8kbnQI8HErP789ylQDFFBz4juLUrYn1cMi+eHPDEvAeivA
bpPjlAUSUY0PKN4FzfnFFftbGqAyEX2CrTb0IO1rCrUKU/TGETJwkKWHPMLq
T5wl/Zk8S9eqEfL6lRDxNOEk4uALhPUmoDLknId1+Zp+lSsSQPpgh9199Cu4
dy0ZDf/h3s96CWcMkEuG2mVj3i0IU1OkWV6egJDMNEn6N4dpR+piX6/yZz4K
bf7Xj8oFBQPzLMkqPkM3wKpwIZb5A3T5OhWkxq0/JNe9AEk2OkVLgIUTM0/Y
vak5y78Aln1NxZCasEQlVsEf4vE3P+GsdkOVqUe+ne7BToxYDc88PX+gS8gW
5gT/eDjOxK655HpADRAIYsy8+Bmmd1MnzDDkkPPKHA4dzGoKcOrXZ117TUvv
fppq4VRY45f8IFr3Yu7VGmu5VGm/7+/E+sRcXDwOot5Z7PM/qxqgutWvawxH
tT2ttmjZSoree/lhHeI2UGWXiCKE98Z9OCfuI8cdVNlawEvwkDGqzZYbbE+X
ZKCXImrrdk5Tec5ZtU1EdzKYHn7x65axtfJisrBRNnF/l42tMHUPJrdO3d1A
1cG+ER2ZWvwlpgsAqRNeWjyPS6N2yase7b2lYq9OgnMjt/42vdUsVLdK7rdq
YRxukX6d0+q+jqCiFhaTntGURY66QgatFH08YgkStzq8a0znizBysgIQkNYP
sDS/lPSQZye+/EhfELB6C/AYfRKj6tyw+E5M664Xzbh3y9golGjQZWqyTcRJ
AfdT+5vmR/F87HU2EkX81410xZgll7TUyQLW669qeJ0uaq7oLq8EhNp95UsS
+t1AukMgMlMbJaeuKFoFogXCnBpl12OA6TQdt+T3D/S1+Gx15ikOVO+TnGu/
akeKmnWRIGry8vW+E39hDH8RmidiUnxdJJ6Y7Ps/jQ70CkBkCHTfDWHgeGcS
I2mhMeXcfTTL1L0iZJ25p82Eu8IL6wbI6r9foPRUknkKMrDtZhq63LmmwjZO
ulGK5PaxezUSBCxXTQxUo43aIPOpjVtpdycXIDqKXlAn4eeQvg7dE0QeOzqc
4sqtHtI63yVT/RKZze/5l/wkdxAbEG7MHsmt1Vk2bEB/vStaPyV876hTiy0O
JHcwoNkJkcEjvSLIgZMQOSt0bS4hN0q8M5P8bHsxJsobEuim4VMN4XdC3tnf
sTCcuPKFI1pwc9O3WLtNdQ+F55KOl7EmqwtZl0cGYOC7jkoya86SEyeWfi3k
f7wsliHa7AnkdIRBcsDW/FBOtir74Y05jqmkFpmV/No/EPmONUMK35VkaWXO
x6QAKlhXwnpTdg8pGg3heKSoBs2dhWkKJNzAnijKywtJ4ljBgMbAoN9wStRh
eRFhs7LjtdH1edi9ieezswErElAliTbXiKSLe3/jxOKGsm01pl0J8CrauKpp
pXnhdMw+cv6Ecmx/DrmfW0aiWj8hEsasfdvw7bVQFXDQVqN/Bt4jW4MQFU0q
zofCJwAuJkq5ZVH3WO3tPUaS4S3YMQRBA/91VC2+wguboWnB6XchMt3UB+ES
6rTA5ovloA/hE69BkB9AukrhgL9LLgtmtoOFH3Zzvb5yA2jzYiNnISNNSNsy
DEnBjejw1bfyW48/kTOXMh0GI/FsS1FhAUs0FVycRkJau/hZ/hVi0E8fnM6B
AENLE4whV4aFTJ5tqO7bfTmSL/Bf1OHc2b7cTOaau5G8W9JRlVGwTaAjLrR/
f30swCRm1TuZkTDcwlYaefKe/aGh6UguO/G3/P8YhbQmy6fmEYUA3A7HXMCs
84EvMW8jyx1Yte2yAsV2S/80puTUQO/G3FsY2CwR/P7E/p/0RHbKFh4EJtxq
+Zoc/mY1TT7RTCNhtVc7xUPL2x0XVsfaTo2qwQyjEwZ57CaBT43SOX5Wb456
Bp5Jt0jfzf7dj2utAgOzeTzjgchg6F8bGPH/NWfA+Lm7InmboNbVXmkVbNY5
zy8u+A6IYChuQ2mVp5nTHkrjr8UvVyD1wJ76+QOSXvGdZu+FB3OB+E131vhq
KXhm2FaJIzLDRpPOddYR7DaZBLxhpWVyQuhuYkwpATiVU84E+/Cv8itN+ruE
9+RBejo1h3qol4eXQIUYkPY+/HsSNMYQNt76ZWfCB3fBtwzIXNPjGiOluJNI
T1j4/fiVxRLhyLYOrAxp6RzgCaibMIkKmyKYtkkXlsYYZipkdq/RJdtQcsUu
KNpSGMkFJimRUz2uvHta6VSLclBKdqCjDIeDer3OuKB1rQtr1Fp580m35aY8
FPmJV/6isN1P3Kx8swbMH90cAhKllHMgfxY1IUX8NbWEg3cpQ5XTfHZiNsYw
k04uOuIR20u0QnkHblJKxN0+CBMuWH59pW0O1k2z68rlD1u6bpw+BKje2zpc
uPVQgmZlQVVsc+5SuCV0mgXl9Xbxxt0LoHznbJrDt8o6GVUgNa17h25MNY4w
OsSm31Tgqk3wkSS774qlZy2uloDoKARnsxaKELdYe5exTXxXBTadINET8DKa
gbqTFa/8BfaOt7uf8Y4klgEemyZPPiAxP9lJOqWTJXFeNIzQcf8PqG+4ETzZ
f+wqyO+r6f1Nj5WqVKpNC+H9warSyjlgdvx7yyWPTAsYERys8llc8AytD0BB
pHhPQ8T4tjQvi4v3JvErBBth2uJwxHpDIMncGtpQIkrJck59kp7oMENKBY5W
tv4c09DUljSfA2OXhp3gfmgSrWE+lm7LFAn2fyv22qo40jFAQiMKEJYKAUkt
ETaNWDiRRzv9TZJPIZLyPcKtx1Q330zdibcsb/BdCkd/LQReov7k3X6SBSA+
s8cO8VQvmS2hWFW0FAR5CzxQMqMEPrEqSKJ59BLV9rElSrobexfe0s2otUmJ
sakwifJvurs++cgDuP/5kIUPWOQFWtI6wwjlVXvpKUCKr1oUikxSr+UALHIV
ZF7aLBwKt38VyBzuGRId4fn0QuBoYMtpz8Grtv4l21kQYVaFHOBm+PK+NCDv
/RC1fxHkL31PiyezLMBKDM8Lqm0RiXO2yhLc84eEv4mPji7n2L8G3Ss/hFhE
F12Gj4yb6sBJJfzzAikeLPrDbmCBlchQ1yRC3FS/UsVnOYj6FQEGUn/FEIHP
CQTsVYcMU2H9QwtNLtEkyt9rc8j/0IivAWUdyw74N94x/NxPaAF+sfvYzbGq
qU65jyoX1qVUE4KkR+2MLbeg5n5rczhHBz/oNsXS0dnkxtzp2iInpT5YNWMD
9WerVo+HQ8m8B3BSCS6myLwPh4F1AZ3BRuSzKrYu3R7bH65fUmIl4LhyI5q3
xD6Ak6ksY2tSbivq9unW5CwQAGY7/3r2+Y4Ox1qT/qT8zA3BS0rd7Hnm+wTr
SnZ/Hmr+WNQZbt2tw6JGLEsuZjCB8CbVR6T10ATgpybpz0EQexZXb7Lv1XBa
ak3rEuYsfNAwryqO5RDq08B6Mz0sYh0xM+h6Dk7tS6r59SveV5GkdjrjhNak
NJ+v4cpd80/5r+rByOPDpA1WZZIgObBIt0ietL6GMJFLiOjtgEVj6RUwNPMj
EISHJuNiEwWMuxkkrlNL35ouc8sl7hRsedn+v6B5aJsvoQ5kH+h+pBcW+hq9
+NEOFT2tqTgPEDpXtN+iY+zG/XFExECtbk2S/zFx3R768buBo/eaflqz1BQ7
LbGO5IoiXjeYFywKZPW2tMz7/YcAgoLbECMeL367C2fNiaVD8namNPV29FbI
ZlXWfzDIfcCPbXbMpEJM4YqGjdUccwENG/fD6BO6DMM+RCiqhEPyD3Lx0LZA
UjPfJLvvpMs5v1iCbHDre2nXivZmfpLyQTovmHCszU1uvk+JJDZl/dYHjDt2
0fngeebgN7uGPnrHlBh1CQ8krPrTMJpIYAOPvgsYawYGBIAyF8bh8j3ovnOi
ijgiTaGxxjX8WKQYGPSkYZgWS94g+24l1yRd3DA0VGRNtWMSqi6uDrfeJ/HW
mSx7U7386WgOCRpl9gX7oEtAGBiqlGrDEkbuL4toiFQ54syD8A6A5HGY99xu
6xOjdDWRyCLMtANGBcDg/U3DdtajbY6hqMuLKmIJHECtee8gi4TqMuXbcOZJ
SAUJ7iqWam4s1qzw7zH1RieghVUKAv8nTcbqGFT4MFUVeTWmMbV8JoREJxf4
D4Cg5SsTBOhsG3ekqutS/p8ycw3RlzqEHVrvkMVQQ3/riinacHY+z9IhjrWp
WuRkALW2OOH9+hMO6HQdRTOnwr8TcYWuqmS5+MbTuQ6vatKQA+XeFt3Od7VU
7x/HhssMziLwGEGaVYsqZ8kZuKqcrrU5oVwhUqNvtXNiZwKa8yPWVYasksOU
629cgOMUl1egMSpQl81t4MQeMVoaj0bIkYXbs/MKBQR9hwBaC9r8VGVMiM87
zcattaSyZux9P77Zvfs5fzwBTzOyC7hfYaN9VX/7DGmR1XGvtPaG9zGbOrpZ
cRE3n8M2RSusteZ9adMkeozt1/7gRHq3ypjVEow4NP3WYOb7u2LyVQTXwLog
I0BKYblAj0TI5z0LgYX7XBsJlkB8XmUaxTMFnUSeUcQll7g3ojc+FICaNFxg
TJeZ8gmp2/rs6jYyETwFqcphIQQu7Zk1GsH+pdsSEby3Zq2rFUpoOtv/Ts8i
ideiyr4wxxEhvh8gAarc9rxH1g5HtXP4ATQSEs3eWXusvCDNZdiewYQdnZ3D
PdM65KYCMLnMqmZPYjfT6OXNUAdNR4s7Xny0ZvHBQrEJI4HBkibKlPAfk2gQ
G8yE5VALU+4lP3U2pywXp/fToGnv2QtCxQwAZFVLLAEq4ZXJVuMxaWFwyfRU
OzcFpDqJVfgTbR+3wYHE5kHvnk/uiEiKxxT8nBc/5GaWJsMFHb6n5rLi73pF
xV7TP9FCCjiwqkhsOB9H0d5T8l7fzM4Gd32oA0+rPVwMw8EjeexdsSzEO/y+
0kXYWFwc+ypYMrH84cRSugcJcIwh5PoDEP0h3IdTrTVwwugZlEUh/6BlEG5F
gXvakw+hnE+eCUZwiv5mMjp2+I+nnBUP/LrRM5N4AZ8g+Le9TXfhxs0j4Azo
Pkg4WncbTLxo4HziWIK2i02rdj8PnIKBEQK/kN2o1SgQGP4D59cEQgH3Njwz
U4kp1gsxOaDMv9WQJIUiBgh4wwb2JAiEzJMvNhDmqMzifK7XJJVNP/TmBjNr
SEH2jqQUbOnwPIBpVs0AgvYjYE46E8mzQuk14xTMRnbgziu208gDWPzowMys
XNe5cfPSEFed4dU4l63J8PSjWtZvSeBlZvpbvNC9Du5YarAXlXF9fzn/yndb
Wa+bqYXOH/0Ubcw8H7gwJI8oHaW0n3ed3+iO6jFxnOUvqz2CiiXzLkYAc2zH
LxvAjZPhFUHhGAgFgUecldDip362o0nSJ64Q8VtxS6jAqJKwdu+zRoQ6BCus
cNRUbH8JEYfOfuOdqDHE5bHYXgtoT1PEZUeQItnQiYkE3wQyA9uKwiInA344
UPGjGZH1XGoxnJuYT6T/ZVvIHJhYvgh8oDZv84w/EV1O2y8yGsP8ev2YBEMX
HAd0marHNtg4AS0/aTQsawNtTvyjCxHZ+KitxxAtlXU/U1d7OBxH2zztPOY0
74lLxFS/6GNJu3OM8pgHimmoYBqt+4U4yTGkui2oX44z5GcYGQJdNqS/5QGK
2iPsRo4SBLfGgwCV7eLm82cDHBYv/eo6epacLsW0YWKiBxagR+8gdXTqI++x
ZeMj+hUMainPZRbEu0KNpHIljM+1mwbRO5g/0F3x+Jgmksz50qvBZf92cDgr
iMERjqMNDajs5jwx3dGdcH5Ef6fMS1kHdKAY726Z481UA84iY6UgUzxAeuzG
NFMQebl0185//zrVMXmcOUrlg3w/fPVUUJjahcEr1b5BivdCczPGMN7xj2rA
MVO4ty70AdYxEPTcga41TOE6VdC1sx2m8asPasa9rMD0HDNdf/h6I7JbKIGb
P2FvgHzrc3QuBCZeYcqj7kwPeKFsWHqfRCwJ6FQDVr5ZKfWs8pUj07EncRYX
gSQ2qF9m3TLnlObv+FoA7tJnpikX+y0fJeUsofHviSwttWIJRWB4GRiq7eOu
Z1cnPvMNDzg9PlEI0CkJ6ZGPVHLpRZl52WAzh+aVXkpcDzXNoPpDrnwshBtl
v5LV4q4tR4RsBy18EJxGDHgx7ENbfkFuYS0Kl70HDu+Y4shWv2bBNjncCcm6
JFkfDlQ4uS4WKGFmbxqxCwbyWyOk2Vd67KRsso2mbY1IXjwLhNWQyWx0XlAX
AnzyHNnAPbBLgtrEs5jJrjQr6K1/wwqf8zPuhUmE6Qpthy2m9NaFRFuIRU8F
tLkWPEOOdbG8j7a1tO/hV5w/WUG+5O9r+kn7PgvZwYYWqQKJamqTjGQSZ/hY
Olwgd/x6Udf3DZ2b5ie+iLzDg/aE+Arx0V+/jVuVJoU/+tihwFTUv0bJWV27
lorF0iRQBi+QC2mZuCciYSyFD5OIuzKC5gW4irQ2pUZ1TBN+LuK7qcfi332G
N7aZjNWAy3vwKji9KzJTFQ4Z1++Bp99JhnVYjEncilMlj23NRVaMl6ftmFrs
B6It+wBb98OOyzXh9plGyc3hmsuNkH/Np2x0zRblobytUXYIhmCyfRMJnfjO
DTNITT00nv5hOmXh4L2+H/4cf72McZIojYs0UyKBfOo/bSc3t6LTys/vWJCO
iFKYoVpyjkQhOs9AWWbBj11Br9iX89XobCkA8MGtbN21SO+jiU3BegrJCVTV
UzPPVp32ZrGaA1rv0auV3L1gMvRUxuXdWDJLsRcq8TEvHpEwCBG7xqQ1YtWg
f4q9szL0NsRg1wGWGxpYWpTB7qSPlPNRA7xkrCQteV1P0UR57OGvyLCzwOCn
8TuwYdy6qA8Z+mdCdOcdN5+Qvne++2bT5PDb+9p2dhRRjtlR9T7rJ8IFfvZo
lLqhtnVaypCGscp4kb/B+GT0Yu9Bpyb7NU8gL3FffPUXCkoOMT58JikrUu7H
jXMmK+n2YYe7sTIi4fmJMiyxa9mU7kJTXrxQ24rTHdMY9mi3zUXrqy17yBAB
v75lJWqstvKliaOQ8G9EwLxP0iN5dJfnrxIWc7Y7xstFzfRtnol4tZ1+N9Qk
92r8cpheNyugJTONmw/HEXubj/MUl7n8OAXlCMh5LEC163X40eXHEN7ay/Pc
nbbD2aLLf/27hB8BdAwW7sh9+TMOX1ucc8jbKRN5KMF5PkvXfnU6o+Lb0G+u
laMkXkHU0MpmIAE5Yv110qfUtJYHmb1kC0OFhrm1klFWkm6+4EX/ghfOEBCU
n8S1eUXSaFQ3OsUE6vg5lCpfsNRS7aLUHsH41sgKLlvT83UeejLRTwhmyKwd
sEahgjosuM8MZ3WTxCgjgi+MKdYJvcvXy7dfOlQqcKjQcFb+fqrjxAO1vAuY
EllHh81QO1SMRCGPBMtDMqcjDQ9Lby5Yf2vbS3BDqfRjwpMB4ZHGGl37+7WI
kSuYeeNoAkV55cRyJ2Gp1cxujiEM3QEHmdeYG/3pOzGB364I+GEaR4gT70uN
kUGcMwHYTSPYpEP9vZEq3IRaSZT4xbzpELorYxk0l8Ww5+Ja/lxXQH5YTT/j
UCPvs5twjIaR42lWVUsuFFh/iMHPW5lzQqm3vCVcyAaUzQI+31uRp3DT40QY
3p1T8Wh9E8CRad3F6g2DTf6b69F0KDXBUxlAC8EDbw2CnNKTQ1zPBfdHYlar
WTunYfJ4YggymeerVusCK/wd+dGYtf/iAFzwd6tM7ph4Ns5fh5rhrYezAiHc
DnrO6DUyUH5tGvlM+Dhklhx6G9UR7681FPHfsOcvNPcuC+AiTzY8uZyuEYib
N/Bh40GLvEq2SBBGErJezrRFL5FDhNBUWHbTwudTjxTuDnxHaSAfNQkLXXRl
V4kcMuy+C8FdS1ea7uNvjH5iREjW/sLn+Q+OFXYlmuYtmth2mTxxm8JKvKUe
B6XQ7AhqdzWSTtIeq0FvG7TLPSgE6SLYZ057FTprWJkA1Db//JpUmb4KH0pP
6WN2G5/5XojoWCBp+B/Nq0sTXsjWCCREmc3ethcLkWL0tXHxMAbzFLtormqO
wy5vv02OppSpDujmL8lm4JZJs0aCQgdOGTlWZ8IQLl8bRj2vTiQY+6xAaBOI
Mxk16GZ5UmZp8A+ew/ejXnGEIMHSTBYqIpZTHVH4+y54iJJn/41DbdwjrUU5
JASoAI4Oa6oAU6RxbdrYDnDffox0ojkmawEINPiK1SR+z7cbmJBoxJLeliZv
EB+lV7zoPrcKkPdSV2zMQgomhwOZBaN6JWVfX8WXwj1OAvh02HRwUeKqSjCw
HsJLkflX41whcmHQCM8BgbV20y6dxw+QbD96jJ6NjrL2INJemL1/ySyJ+VdK
Rmgz/1rVR5tIwv1zJhpCv2UiLu0rlCTi4LsZoLPbOwlibVVwKaMHQFkFpTXg
0oWGJmLSIyQFCwmZAvJ6AbasQs3QBS+uUuhuk30Ws5Y8zdw1dgmZVeu3KWJv
iOYol52/h71DLDH3NJof35WlqcxphE2rvP7E0wDBHz/Q3cCT9viRGnd+cmPz
sWYrzxcQFOk9HyhbdA65nJqlhHPuV5AUWWBCHH8gv5s8/6XRqOjTFGU0gJ46
KiNV8vm+xRURCDbE3/iLEAhXHVcH3CNlnfC31bWXlHf0NviH9gDL+q540urz
XOX4CLx27h4sdkFZu2y70riDHmXdDKTv0VBvSIV8rk4ztyqg9OsiKETamuBh
o4AZgwWnSQKIKX2j41DP34aGq4LlIhN6/MlpU/ma6N8W6/H0jL2As+lFV4ET
W1ysEc7IKSeBKrtTT0Q5OanqyQRXDarsPXIvWzAWOgRqlvCkSMaZlCTzBXns
ZH9+4cw/eU3HKomHNcyuyUde7cPQyqG2tHaTEBAieDYvwHvCgZ7qzY4N+2CS
kUeNzBkf77Lsf1xzuHBOnFjZWpV+4Z1H0o8mwaaEzTAOXlqVpbo697Pxaox/
/15qCR7oyBkLF/Y49qrj/zYVmOHl8CyQgeGYTZwg8D/SGnBGN6SQjWF7+Z/c
UAkXF/qfMGNH0pFhwpfTYCMcabApXyog3VlNdxvO4hZaCNPy6peaC1kynbvF
B2CcQKcBWRfrDetxZ7aw/p4DBJZ6XFwGfhQdgtbT6iNnFwNKPlj9BGx99dl9
gRUScD799GScoQaZ3dp/ItVB1if8JUxo9NHyRaWdPWclm1PCkYb8eMBBddFk
mjRHQ0BZbfP21iMWn+ltu1CnDxSOYgsdudeuBcBHPjZ/9mdZRVqOD0sRYRb0
PuZ3+i22YEHb5czSonEn5f8FHeea/sD9Fww0NKDDrpB8HVAwTi9uGxx1fdTZ
FoxDUI/5o12myzxtHCBnpVV6CR/NINlPc03RY6Bp/g+jfyPvXFm7wpja5+Lk
uQgbhOhPPcTbnvexER3ilm1AIXJl9O93+hKvr21RPFGn4KUOl65bCJY/qEPt
A01B/AhIrrqUIBTBo5ynw0ISBLL1bnzjYHE47otA3jct7EankkLhp4zikFTj
59qPuKpEBFSkIv+mVGLnznsi5tLrpoHxGQ3By9yiL2UGZnBMghbq7B9cWsEE
KEGnu6HPOuSJ+nmycRNkLbYdlpL93V0Oay7QK5HV63vPhGv5xGltg2LStgdm
+66trAf/dv4fIv71IUU3lJ6UYaIiqBYdqRKxVjsVH2f/ZbW1TI298UlB9H0P
rqAjOssMTvt8KixEzsExr5Nz3v1+GgrMOj3dLftMShOFw595QUfV0Fioc0Sd
i3ogrtfVUj25xU6ibAhXlxlHEjWICbfejCdgKxhmWk02rqoPTgZFNVWqodko
5T4FvVQU2gsMnjBDejOmtP1qXjjisinu3sAyEAPwG8M42QFSuA2/5Y5PVLNR
NOV8uJKjOE3jQ8OEonIZM2RYuGkPpJp93jMTqgBmpvx6+Z4wkFrloCB2bKwx
7aqmJOxNMT/SoNNSzGrBHG/aFqS5mtsCqWSIwHr5JFBoyAu0x30IdlDfecMO
G38l6PGug9j9ONvkuogLcDszAAx6f79AQi9xRVy6We0xJ+K+SrtnvH/v0MQO
UzU7rZw/MkkWwvuD1fIsHtqA1IfNEkYK44aN+9CCezkoiQ/7SZLm93qfCUjk
IV7PJ85R8D+ITuH73ryeGvDOCO6EENjNySk0m9qdU5Q95SWVEAMOjjsqlBwQ
QuC1dtHrs4QkmOcVqG023vp9qidbpmnJK4atJDrWnpf0BYCYJeEszgaOBOAy
UAfHrmCByr90tdV4Rq7nw7vd3zGWIjBp/eNlpfG/TGNc/+pZHNumX6yQCzwa
EcVxyLIasMmZPOuxQlGERRpeCM5Zg4770QGqYdbH0+gdF/RPc+sjV7dm/EQO
78G44DkgcINm1Jd4k3yZFFBVAgt9/biWbZpXmKjaozZEgL7Y+NxxrVFH9v9m
qtUrznEBZq2aKFKkuvOLdoOnibzcHObHdY19blUHn+xsqdDC7jau2JKn5uS6
IIaH3ZbbQdaazKenu7brImRaKCdDyAUs0YVkqmB+WKEX2biAJ41WtLdozx1e
weORxRR5FBVgvDdne6+pZSzyub1OLCmG3ZFk/1lgNNjXrpw1HIS9MWG7BJc+
7sA3Nj6KDz+X883sUeMechhciWq/9+aSyGvkQWw5LEEh2NhJhuvfvf4IEuMM
BWRBNabRSr2yfLYeYZKsN1KejkG1hlr+uEbdqI4dnGAVFLbqfihah5AWVN0r
odFcqk0mHX3FO7/ZqjU/ZGMS3ciYZ3JPyGwkhSbLRxxBd2t7+LsCp9A8b77u
pUeAq/jZBvd917kk6taxp72H3VJ1czh24OA/hvhEHRn6UOY4dT3o1yZZuPy3
QwC/lnbkQBzYzH1TZlfLibBT29BaDzm2NZSP/1nxcOGXzJBQIp0T6R4S0doH
yOCmaZsM6fOGcSyjUGsov8JinIJmnyYEA0k8mjCaVUHHhOTeh8WLB6fC02Ve
7cjJcze5p4unvRXTwZVxgON6UVtza70fYvu0wsIud8vbb7GF8eOYrbu1Qnbw
j63+F66ARWQBxiT0kq180d9b2nO07ni+9h82evAybjOqymk/+jC0rTD8qW2N
1f6Y9w7gLT6pvIcevBCQT/zuYFxM4fHaSSFia+jKgkdyIx3ROqf4Ei9FkOul
EC5Ll+un8aSNc4QJxTJdo/NwCpOYe2XOMm5BXTblO3ZsswaJK+cWFU/JZ4Lr
afiHAmW7EvLpPf+zyVfcPAjFluDZtGgKXYDLesu3N/2KKUeGopcjgsGyDRYk
EO09zs0+XFs+D3DTXvEC/W2ByK2FT2cEesqkQdUIJAuuiBYcz0x/cagjvf/z
TDjjnaQLLbh37ufcQzB900BB59hZgtzd/taGUMtbomSU4MqLoiBuJXmm5E5c
F9I9Rnbj0X2fjaQDFfdKR2+X+PK8029PfSTiI/6zMtYwpemgcnFynvudeE6o
daaG21bAM4dHduMj8GE7b0j2DiF0vJg1ujKdtAJhM0AAFA6qU2ff8+1ku579
598XoEHVB0JIMtNoJPJ8CiMDFQjHE9ISKejBEwogCCNmqVOzug+23bcGQdp3
GU/qu5O1bKqjuvHWknLksaPcN/kCx3EaVYw4sro4nZr4/03aQ/f1kDDYHCsq
mxvBz71pf9wZQBTAATMPBB/aEFF7CM2lVOyEKtsJbygta/l8ngMoqTE+qrtQ
vFHhU8P+lrUD4xZPWSq6/HZVyuXRTGxGjauwPxtmepyE53uYYEX1TdesqFN5
PjZDsNU+3IplCZVfilNElqFN3vcFEG3mDyX9k7vevaVoLoSp/pV/dN/DriR5
pF+W2Rt9IJLsf6XlQiml6I3vRKzDOD/YH1J2L5FFxunMQfJcAscDcjgsAS1z
wYEd9HE6RyQmDchXG3Ifv9ia+rGJTRk1kt2rWIZJFs4Wg2Tvi9eSTPPX3nh4
fQr8w8YH5TIlCsjHFP33Qzn/6DQSpP53dCueVZZjiui/UKWQ5MjM8p1aD1wm
ZNFcjNzV8JOJmanyjOMTpRZi/4bsRSYzGpS5JzGdMt4ShNNH8lVTvCCmp3lZ
bT5jEyNu48gKjMsMJoyFu9qXvJhRA5b2bnElP1ghDH/irY92q0oCzlLF1RBM
kbyMDe2dYRlCCP5yNkiuMwe7/WZp/C9E5XLeFtbtNyfrxku/GVSjQHnRyyBJ
S56JZgWFow0zl3+Ip1Pyd05sX3HZjL5LcygEHwKaphX+UE7eydtaAv+JPP4Q
C2ejwnehjabxa9AQxt+0oezO2o5hoaaM6TJ9y47mzAX5kdbCve6pcZEsnLjz
l2wDWFjat0CxlbeS/fCepUdbl14QaTglmgYFP3hFevz6Ut1XeihGyKW6oYib
+frMXPNJBzxzyeD0KCHu2Tljiaxg6w0dt88ctZyMBIB/FNDtAkZeoU+aiMVz
ggph2WCUNm/2Q3kVIaY9f0eF7WC9r7dUaE4B+VVncv2UEBlYi1fnaH6SxDLp
/hHqATHzJsFcUn33Wj7A7dIyv650eb5heNzCQGDe7EFjTaa/Ow5DdI56eisU
dc27/5iE5kWbxG5bAjtXy0lgOApuC28G+/KFWaMQsUp0Oqi5sJOuZnycT9wg
Wow1KvczX/CU7j9fB6jJaZvra57wa9TdkCibcWlAUEM6U2GiaxIu8yIfFhXg
p5tFrZDYtpR/xcj2MD4YduPUs7zy/U6X/xe5g+bYTTA2FlJCIS+Zyq+Vfva6
NbPqW+TDYA7uSG/SJ0QXhHSXgxdryGACZljhqJnE871FL29RmUD7xcUpMADW
feOXWy9LEQ5j4hYHrpJCNmQdagcto8eJ8U2nQmHOgIIZ2Rui85K5bkO4GL4U
+PO56jkq9hfIesqi2GrktuT8vssMILeumrh2yMzalYJCyt5Vo+IBfTMXNGUa
FfD7neUmxnWgDqAqq+QWkcqMQqNk24uN6eZFViErvc808SUMUIomfcpVbbdw
QNa7RgRaAbmFx0iPnspDdgkeyeGnh9qH4zIZQOCYUCYg4jlmfCpNkIrbMfoB
w0Zt37Z6L1u+ifnJ+Nwj2u+m6HtCr/Q17A02oCvkO/O1raTLtMZ0Fw5nYXDK
4A3hcqYg+KUBDidgI39+Phem0Ay0mxH8kxXWiF4W3epZtZtqO7ZrdWHH9IhA
pD/yHLhzhJlGaDD2Zc3ilhfKX1tEkplXsXYoqOY2BePtUK+CGPKJkYtQkB2d
l6ZQmkqeVYupSnJoU3OiyNCx8lZBxEWyYVR/0yEoAktODERJOOM/ik9W6nkC
Bwn4NxhkkUfhfZv8bvMb80t/RVMlzGMAUuMTXd4sGcbriq/Y4kwM7xTdISi0
9BnBkCD1TpZZclqge8tfRI5c1YbnaNx8jvg06KXHj5uGe6AHYsWXRb2fUy/R
3eNu4+8BrAqW7sTjSIGjMPvQWGiCFQ+p2Hh5O8Fg7HMJDdJXc6qW5krD5Q3w
DE9ee6AcTZz1qxKeNXy3w4qTIcYuy+5TVuGfh6asEfYygqcMIVJZgw6BFHXL
pgU0DnGqvyoqoVeLlOkm/Jkucf5NzJwlNkAHYNu1+kmouGMq5u+/QdQtX7PD
1xBKnh8lfef+iPJ09MeCjRrp+zzKzt+tdQMmoIhmXr7tj/MZD/YVV8P2xWwi
XlGMx0asycmqpEz+3xDsey/HKdhkBJwXsz7MP6Fk5QgPGwoXsDPT2M/DKNCP
8JwFtrRIUWxeotoxwzcg5PoOJ4xEIphFdLEJYJSlKs3JvOO6VooWjQtQ6m1X
3Gh8dSbYScN9tWHbvR4L5kvwbwFNgXctN/Tf/9jgFBAF/uMGe5irJCa0UwZe
DoHy0jq3ZP9MvfqNoqO53DCznj51As7MkOu9NOXJHC+pZUOIxuSJ09iCB8J5
eLV/sdizKDml8n12WfZly/KHsDNe728QjvttBwgHzdOFFODhkO/oE8uBay8H
hPduC7RuB7JpRw9yCoe78kkUWjzC87DsB8XU1kK3MWAAa6uGk1QqLREQAhc4
nIlEI3MJbITnyLesqYiSORA0NleRnZKLHtPLBSyQzhn4EZneOetjG/QVKpoj
LpibZ+kt2LvbwUXKkyAh7amj/aoHeNiP7yDne/ghkHvp+omR9ykGNlIuG+y8
KSz4JToG9iyFBTb5QBxjrARzgMSYeAqYqNkZTZ2wqE30BDTh1NDFlPsNOdfu
hy3bq3djQEF8tUlHWCq3qJGMqlgI1F0S0c2JGsS0zGhwTFInfP5nE8lDds5w
2UUInd57Zmp5jKD7LPzUQ+6P5FP7b+3YDrzI/PHD8vKC22fcjU6EPH+DMHoD
Gn6KBMWLkiybR0fYN8cR/ZGW/BLHBkJX5u1LEM7/XsJ4mueWBZ4sJcOYckqR
54sXtSp3x0354XQ58d9T/02teEmiABQCad3JUD/OMrLM1nwgwxUWElywzFNN
AUxi8lCdWT9xORWD9tkGKHVrrBsksNLy3Qz8eMclqSJRnvpAV8j7nr8VwtVz
88+tE528oiSwRb9z2qEO9/fLvjAQX/0NP0g+ZtRuwonPUWVZcoBvyKY9ueRG
s6NBdyqyMlq2hlY4Rsw7x1priVwoRoO+NGe9BDZ7PD1l195DhA/GUP6iyFZE
g21SmQeBSlQrJUzZs3F0MMtTbBpy6LvgGhoAHITQ7VD1VCB77rMgpIeD5AwH
/g4RqvmmzlMyRTyF+g7FlGBkNgUsGzsZvYs1iFX5lyQQNYcm5Jo0G4Luz6ii
x/cgFZffCILUUz+17FkWLVjhtMoY6d3w3nqUh7STcktHCqBQAKPk+40xaAzl
cywmFIzA/IXaynfw99iLuaJdyisrfVZQjbfiK50/iCnlI/dnQ+g6Br7fYSeU
o5dourkbvBN8uVSfRHd3oNrHT+55e4P6sY7m13r5TF16U3w0f/g2NgBRG9dt
hDlOskD8aNVVBxL1b1SQ3LUnGWS6lRA1C5WaN0C0Mcb2B6TIASe/8rhFfasX
5veLD1KeBGaKpRRt28zrCHHFN0huiHtU8YK0HEWwlr++dub3MiayMQOwMwBn
SGTA1afx5qisHfWpyTZ/PNymAOpXJNaljk7DgChkTZivp8JWdbGwV3buRleO
hblgKpkelv4GGu3glMbGljVjRwj9Y3tNpmVZ5S3r0/JEsSV66dcQgCAjo4xB
yN+Uxcjo4Fv7+iQFDTw1vtqKaEMtpwOWHoHbVeOzut/Wf0LMFA6N+t9H/rLm
nUmoQM85cHD7Ns/4WBqHmLQVjnmbu6EbLe2NDRwXm5jh+diaYQSWuaFYaJF3
o5EkiV5Rt0FC/sIqGvBWugBV1N8Yq0Ghk7beJops3TIPEyqBLkJC+Jc2jRDD
c20pXFk3UqhVIj9OGQItyxH/SQQ/IjhiDYhMl2gdMfLHnU/rxL6/rqloG5jF
7q4f/gxtA9uHT0Y876Ewz5uHuDQSw+SXmTM8uFmwioyHLbiQjXlU9OuyajHc
ew7AVqYSpu0OU0vm4BauNw8Mhf96Km8ERuOf0uNlTJPqE1D9SnozHbfV0n2k
OAdNRwG7W6cphmzSyYnN9+5+254u7hl1Sff589rL5DHgfqP0SRNip/e+1nkv
/vecUSs1kfjJz3K0dI60n5nJgUuWSGbC4SYIuFx9mO3XZ9ytycyplPxsouwe
aodlSNO7l+abeLbD/e1VWpH9ryg62iKSvwCwo8bm6LmUChJmAk/doqv3R5ha
vmeHDgVhtnYvAsQ/PVb55Z/Q9Ec0pTx5c9lDw3NImovihxiB2R+Jp25gcneT
uEuEkc2VzZjsiAM2PNH+lAYwR2AJEi6YEtAoXbic02UfQUXqju45GiAnaAN9
LbhIrKM4pFwuljzzZdl03/VHqByf9Com38zssvl2/joH+sPPic4tmuHBRpB4
xI/OWIF6AoecOHuzXK6ik/Gid4uGeLHHs/ydxJXVvE9q8/tv7IsQY4AXcT5q
q6tzIvTZDO5DBNr+kREG2E3MheVZA2PA51tVcg2A7moYwkM+yOvfRwU1F+Y7
8jNvC6Xf81QuSXLMVgTSmkBifCujlSpJkqAHpPnTpFDqaZSLQsybBmPb8RE4
QSV6TAjTzf6obFc/wsl5AJKgWMLRIyHoijWKafQP2GR5RYajU9IWODEwuFXn
7cdjfZ32d5ezHcO9BjfKja2qOx+mbvpQ4iM87PjWo69C1bW0pjD8XNnLl46P
xI2N5csEpGu6UTFAMqNDFswZiA5xmdLOgAnll2Y4RM5R/77YkeywCknwnrkz
9kFbBqu2wJhx9jI+032hyUZVu+FU0aoYx22NH8A/rXMFJNqf/9n3cYsdH0dK
oXCbmMYSSZ284j8+9FoHJvyJcKG961ejKUZ6jFeXTIgxMzNZnyd1xFJxgcLO
8vaMi+eGvrxoqWSDCcDk/+Uo4Zum1te6qH3LUnZdkZUvwl4jC4SR+Cqs/6Qw
vra8OxFpH3hJsoSSrWTDV55knUa+LjdD3esaPEWVFfg6dVmnFSOnuQhoAHBw
AvK5Ms9Pf1F+Znq/+0h8EhvjfSnFEiixlKCNhjNfv4cZL1xNAwn+x9E4/5im
s30dK4D+TQ8akR87AKqQs0Q90sw/gWawf3/Alw0+cLVb8HPs94KN3Oi+x7LG
9fsZAb5Q9NXmpLyowu2bcI+13eGs+Mgn1Pf8pRYeE4wzgUl4mqmonLMDgspj
R3CA0FHdubYEL+GgLMqM1P+aLRGCGwdZGuvjnsiWYyaw1IJuDt0l3aoJCieJ
qN0YpWdEvf0aAZuwbQv3Uww3fh9qglp/MSlJHb+YVEGOy2UB8Sawla97rCXY
wLSep2jwOMx6pKoTx3pic4667rQCt8g+6dp4ElHtzw5/FEPH/Sx6U51ibX6n
EnrqvCWmQPLvTh/yd6XJezcVWcjXEzwsDohGgFHvJKVsA5c6B+Yl8nny2D7t
A/fJFLLSxD8f0vApRT2LK++WE2CtvyugT0iqk5meMoGC1V/ii6e/f3R0OfNv
iNguEQ8vr8rcW/xU9WFar6TmjbFqLALnxQL02xyZAHdml3xQehebrM7ECeN5
defvBFKhJsEsU9NjZlZg1nGqGM4FMnA+neDRL59L+T3azOvg+2Ab46Q5OE0u
96Ppzb28YgysP+sraEif+oAupvfqHztXcmnK+JpIWQB7/7m5J+gPh4m56gWO
lLHkFW9zUd8GIPQg3fQQGZnFAVzSOwTUsyH1ztB2u7wCqbyMquh3GUeNiNJc
wd49iNL8UJTal8UUJKUMnqo26fkRfJJLh9bJU0b9+5aKBvD5Lboq+TCUIo7T
1D0ZduwuYiCQXHV4mXiwe5Z7JHp6LeNi/bKbQn9+fyvc9Wd+YPdHZeQbYRKT
HTjCXdY4YMh/ZzhSzjQKw8uPQjButMsgx0BcnydUZxfMUjM2gpvzXf561UEv
q+5Cvfj2V93UyKzcSKh8IIiRD/iIrce63lwF1xiHUKPy/x5/9/oZuJux/0my
pff4Bs3y2/aMMv9/5i94lOAxsOx+5fC7h3OhQAAoFY6PS0t+Ie+bjWuyfkxO
wQufQFrfNWZrgx+CacfrARwgEltsxCnOnB1ZIjyWROF21ES8EKaoj9TXXMeM
45cv0BYGUS0Y44TSiMBKUbJiIKOzdazYJxNW5v9qvE6m7KRDBFgm29ib4lpa
aywNoAAyqpwY8KBNL/lzt93tb/7rupry2RxH9Vw9QwBHOmtplCwPImM5geEN
mynRhMQqQPMTKImaGd29YCPkp4ikJa+yLGv5C97+TzeW2fIxDEhrf4/O5c5a
EEjrkY7VWRhH1fSZ6fs4CA/evzldyIcYHMTsiRLtWqyuF/FlQtIEm26taVDh
sZaPVqdmFDXXvV9uJmdefSjpEBsJA+YiggZ4xp95j8xVp8CYSrG7h5oRCqwm
FsruQpr53LM7+vN+kwiyAUyKBtiev5sOIRR9o9ljO79lWOyFjNGyhuf8uo3F
N+5tbvivbK5jkKJGTFDg5DXJZXlKcoN55S8+c3bZczPjqSigMKGy0/vNgtr7
bCja7cDDfz+GuY4cY7OBqU0K6KdyD7c9gnyqDOUZTHsYyBJ/Qpeilg5v3tUc
ChowXt1qwOZMtkS644OszgxlHzhNBRCoq7cMplLz43S38A6BGvpEzZQqwIxD
curopzAeRuMxZfLmW2TaD8+bIy5LIYWvXSNLeH05Hc/K39iNzRPg2PGmhMW1
kryJFmkVsBiSm0lrNQmxzLN7sf2PiFXxI2lDDBQ8Ga2bt8iu/NWoClPcxQem
Z5EajZ7geuMBjOsoVQo8922by3g3+jOe5NDT8Jmg+YaIie5flV75xCtGvsjd
RqoSmKBzQc+gRQ65Zibyp6+Bz7Ye6nIxMrCWG1Q44rK1l5MFWNUamiAs90VB
haSB30hwQKWX3HNnq8FyocX5dYluwk7t821optMKzkh0dJRHa6MPDiM+/Ved
8/O6FAiQ/t/Dx3gcbmRuAeYpXcIFermlycaT2NWn3NS8V68rMUo4Ngv5fpa8
EFmHHYrgDZtTEqqAkXHMtsPa3yPdDMjItoyOWRbHp1egEXeR37MY/Ot3Okkj
fstPnfpTDWMzAe0H5PPxyzY6S1lWK8DWRuO63M5b/l/pxeyFivhheC1XmsIX
fywI98p3Dz7BMc9dca0QxyMTMz63rnfdtUuNJDxTFECTTqe9ZVqoW4drzoYY
UtEGuz8ZqacgKUOrV93csr3foh++C6GpRlLYGxf4Zz46sezjJMGFFA9a1oIa
QbrdBveJcql6ws/lgrqVIwWP2ZBRnZtxhrdzZI4Tr0Fv8qO+Gr9GLNkFxqcX
FBix4FGqQchBtiaesXfTHfCHpbV4iKHoQTjk21hEGk/pB9Hmf1865rWmTKnH
6NsQrax5PwDHpO2ahDZCVu4dFIagBXBW6YlRqJsDR8s8tGPBIeO0lt/NlAE4
ZcxKSxRUVT8S+e4xOyJd9mWOrPdg/UjUVEZ6R/wFNcBe2hxwd6kaAvQEGCwb
MXJn5nZaB6sMYv4Rkl8K6tisIBpkJ2K2hYNqaU5hFaT2R+uIE6fb/mc6Sn0p
pA7vKB6Ymoxzhgs7Hhs0LlRNhdgG0MOoVk6/imvrq6p7t9FCOi5rDERy/STH
bXGqFr8sJCu1ZlT56wi5FYLHKdq5sgpaBGhWrnRH36zvZ1Zd6C/gBYnoEcoa
ZYO67JkVLzRiWpd4Gic676xjmFHc9yiJxGFAkD2UDWT9w6BxuuoLXQgRQKyC
4jqelxqaRGQoL+vw4JvMDE3LTzXAc6QL4FhmKvGNdRlesQVdZdRZttaONF0P
AGxnLOMgAe31Z5M3JnQFytqEL5dvuai7mYZIOcLbWWKdFCFx15wkUHQbZqk1
PZ5hyCqjgZ6VVZKdVoUsDzxb5yXiRXZ2CAvG2nfJgdynBn2n9V0H5LFhNZsJ
kSRwOsl6V0ufFUBIBNHfN03mpGHtZKx4XPQ8xBpqjg+JaeNyFVyuQ61kobMg
2FSVLXqzWKnL0HdC+35LfnUSNKNErwSGewXblEqx0GMFtTkzk9h4lObY+gM6
y2oov8c/6/S0SoYpVx3Zd0WIG2uXiKusCEINR7Oc4wDdpl/2AqnzK8cHimyI
+mERO7V7l2XhJ7AWdygjsxlmJrGZILoe9Fm4PudZaCD7AIIuTV8s8kEdO2Wy
rtbsfCMrIDMUoCen70oBRPbiPZs76FzefGAaQGH7ZP9avBj12nqCOGQyGmxP
RDGIhjzZZWT/+4B1kbQ6BbwlfiwF0KICRBkEIeQBp5eEBDZtQcQNSpvbgOgO
VGuj17r2KIxH5jov/jU9tF6bq9ucwFZXh4Sy6F3IJWPoF/SVB1OQIjmw/swW
KlNz/zNQdYdqSB+rPRUqeZi54WIfqjiu5rBaDhYeIWT3dIoo26uIOG81stiY
7+XLhGHEr9fSdsujIUekvg9bHir0UQIkfNVJFh1iSYmoxkMSWNR8YlOR5fXe
Tyz1xtMyyTGPmcqAB67GtKg3YtBVeF92YcemtW3WhFvAJoNmbp9LUTCd/5tz
T2t5Vj5CiYs/q9D+bcdggbetcdn7ZhF4qyoDh979vIH7P/dqOxfl2mVmzF6m
hqVcoryoketo0wDw8UuM2gAopdyGO3cwAzSU02C+TLyPwpAKosCv9/2cxc2D
/jOdA+QKBG7JJB059wIgLNHLJxxdHNejlyLb7lsqsbxwD05GUMNt5IM1yrmI
dr9m6ZZFuF3lTS7TcSoZodRkm9nVo48C2UKZRUyLvGppFoJuGFV17PlEnume
2Fldfm0p0pgFIGkxUd+MI4+QeoGCRH+ZiQ+HDmd4MnfzUouRFMRz3rKElkhX
7rj7+L4Tc/ub2dpkajjPbzQVyqrMztydaI5ZnMbbDhZeDejAbaWOZ+ICIGZ2
bUOodFCxjb2kgHP7u8UkU7YN74dHvMx0smxq1gZD6JgKIYnQmC5SrjEGLavY
JoHwR7w6I/Sb+CjhWOzTzYSiOZnYA/ViZJXJo27th+zZc+BpgGoiIxQtKuOg
1sCKXi0963ArdIb8HtD35aWttAa7WXgCaBGLDp5jENuLHQLQ7QoirJZMzY5W
dV29AMoq73X39CKTHDFurLvyZa8JLtzr24aATsTm1nbd5w/ed4vqJYSBQfzT
RTwiPCgZOTS/XTEvRN376cG1lpQoSzmRLgh6mzqf+FjtjlwrrVxUcAs20933
rmqsmNj/qxNb7v0BiFXUl8nP4+JbM0l1sSa+ziwJfUQGUWtoRt1ZxwTCqZ7G
q+9wOKBrjArllj3kmTV4rdMr6eoWweL66g2pj7RGGlorvtvisrZMdQt3p2qJ
YRKsUSXoyk06eNKpOUPxl7JPjpMsOedc0B9Edmz3gmFuFIHDUdPHG2TC7Gw4
YGo+2Go6cxTjumVypydRsVSPVTmHPRZ0JDHgpdv+oZIOBZjMexUIMBFYemvx
blKFj7KgQSuWSi8EZb93w1AGCNA0RSJ5dAc+dm3rQfC0O53ITSmBx7WBB3zM
it7SD6yTLZsmBVa+ncTYWplSGsGhOwTjLCgNeZMFx8LRBEnhm2MFdTTAxKJs
NejGaMsgG6DPFuspacFbGrw0fJD0mjeXIWFYfUpsbOH0ZwDHNvO+wlGPvpVt
MpYUwhCUFeorol6Bz9pT3rDhCBAPk2iSAnSeMszS0otcbWCVthf7Lm3umOXl
uAP7TQ9Yme7LICcsF8QtBfmT+ab5FQThFPuZBz+Xa8vKU9XiTYQkyzJyM6n4
k+Uoecq3VUFNu9MXLHYt7tWgsbL6qHkMAThxy19P0fA8UzHDEyD6VXxNgrKX
rtUXSI48wSlNaz52xeFgZi7Lvw2PHNBK4FK1DUAxqv0WkS8NdWvOpUKpE/ia
Ud3gKXjDerN1CD78hvyTyrrcguBFZOT3oTTJLEe3jWXNjyfGFiSYxpfQUmHJ
yXeFDtXgDPtsjPhxQlFuQ1d7wSibobNYgFerzpRVX0musrtxDGi359KXLowx
9qI+6KNwDzEPQrV6OFUA3Z4OPRTUQhnGgJQ91DnIBYOLKEs/fqv14xANtkmt
DfvlHnVZufMkwB3yj7LlIHGVKfNPSBvpu66Fpd+TxKOhl+onghAQdzOAPqNc
qh1/rPod2BOsmlZ/9Dp6RIlGGcO6U7OcjAAqLgUf/xEfQVl8P5zRD/gGWLVc
YyBNDhyUvXh7d7pQhM/eEi2j7EYGc+K8HpHqO9s9WtXSBve9AGB1sVbNY9A8
Q6sQIoZy7KyDK+UsUpPnzvjOmBttRmoTOJtGiG7fMccnEGF1sQ6JTMnY3Qj8
I5hTOZgz0s/b5b63DcS9No1w0kkaeagJ1OfC0PapIvaLJ1ywih+35WO6Mf9F
mDtYKEmAXK3zjTiyPOeQvUfKaCsQY4CZBYdLJo75uTxsQpQBkNR0HlFvH1+d
7qa9R4fk20Lf4VMJJtiwIeJr61q2rAqn/n+BiaxRx1pvZetKp92THgxklkvI
oV17pyLBZhnRy50sW7kbrry7pURGrRRGI8hx3bmw/HYiC7cptHgwmFO/djrk
YL1FIDXtAfCpe30f+9BtdDmuiQg9nj58/n4aDcqW4eIDKepaQguEWrIOCPW/
mEwog5q43QHoxcrkIe6gNYWPSONvvNoSFdEY/diK9qceeT/VzT3KAtQeGjuv
r9AQc+9PCAJZRD5b6Ux1o85Bq1mt+oom6RzPOaRR4+Ldb8xpP49NC+fvS5ez
oCGGMoZeWIewQ5AVrt1Xv1ppBZxWR97jR9lEzwswxQzNBZ+ZsSMmFeEBXG69
i/XJVxDPvD7ANLFj3rCXLkCaelcKJb9P22spvmkjPBV9j9w5dwX8l6Jv+YIg
ofEfGSPFlb9+RxyN7rf1upBvbZBPJg8L+AusED42yMwBjCHnLnLkFYOa/rWo
9bIX9uYumRw7634njDpfZtOeB4beqTWsbY9p+aUuiALI4Oznpsz7H6A2bMJA
BIve0Jw+fQ9ra0ui9bwZp+sjYUqogoXEZ5c0PdlBGfKgTqxp2vrTcRKwD3Qr
k5XQ8yTQ6Fp4Ym0kVplJ2HjQEjgCjpiJ8xZq9G+z/QuC0KPzht1rNGjYSndE
Kv/dteIxDgqLt2RYygIIOu98A6iGu0GUF9krKQwSTkYN7wCVeH5sbkXF2kz8
7IiLYC8VNHfep0xVom5sIxbSnCAvxbNsGwLbB5n9Sokx1VUfip0DGxWum8uE
QsKpYe6xA6gj9vyL1EHgQyk8t/iWsPexKg/v+5ngQzorn8Tq+FuMNY6jQCTP
LPsZMIwjB3+FVIvTcWaYhypr6GIprFS93zAnpZSobeRA79DZGxH96N9z1rva
g4r/osl7UtRJtA4FeDzn5vEPXLBQcfMAfx5bRhzLr4fm8USHpE/8SdNPoXOo
g7kKPvkS8NDVV+bh1XFEqfxG3qhoUak8OdlKVB0/ByM8TDH3IvXOnaWVLulk
vaVA5PnzYqN4T1XJg3Uk7nLjZolPuFNRjU6gJPKoFVHztrUVAFsdQZHGLHqZ
uWIVXKny5GMnV11TXUNc2hiQwuG0XNdQj95r0Yhjg6xT7fgTO6INpmndPSnI
gUQ5yGHZmIuP3V3DDzdf40PwOzbhmVJCpN5ZNeS7sKXqmsTCz5mstUXBKuWn
H27cMqc1gEFlpKH3hzsiwCSccks47LAh6+f+3egebF8SyI0bHI9h7gaWuu3n
5I11PyXA7LXWXcNJoiR3NeEEbtco5ufyr87MPmBctTU0PVuLKBgE5zqCZ08J
io8robUZJ5v+vHAbXhLrn1IHA7bnfUvcBcXFDdehc6NfsSpChabT25mnhfLg
+Nje/bcaPQiZcYwevqRwXrZjBW49XDnwIFw1wfUYKypbcL+AUgnxNpmS16kZ
myAdq02oThXjWIuLthBKVGGpDxeFll0j7opZVmyEDfRmhuVmV9zg00z5siSP
7Sc+Z5ZYq03QAFjl9cwxEWP3VS+hwKmx8zn3XE6S5eTteang79SGk4eloayU
EXrx4eBg9elDqJwPTs0Bvaar9dXs3AS1KRTohsBZmQyqaaDNSX9Kk46iASKW
lg2zVJXsAjnzj7LmwlOsKNq9cbV2+fcyeHOwE3EP7DirVALOvNF7NGCEhHAS
TVTHsNLQUmCfc5556yvxYYgmEyPXqNW2jIC0JAE2vjRc09Q5Qo573rK5H15L
afHLTv6R48GxBBnUm2IupceR8HiNhexLvbFfYBGBnuVZuNESIGlVBsDtIZ/I
ZErmGnB6zV0Tq1oOCzf1y1X585VTwvd8rIlbgvw0oi1doa28LjlbOpT32mDG
GkCMyk8peteQWSJT7nNBQM3Mlh3+FGcujr/gZPaTVVGzEq4D5RLcgrBpL+z3
5InrFVtmqPq8HiQJgh5Tk1H+SETaHsr5/zXJrTDu6J9Ujko0/ETngC3bDc2b
DPNOK+1mhjdF+DU5x0yTBjTpMZ7H/nySMOG7XgJPSqdHfM65dGOBjJsSO+vN
5epqd2WQN3vNnSNw/MmPeAd0w4M4R0bcy5rFimd3WRUGbykqNkABS2kXOuSH
TVuIC6ltCbSspGnYvGradlTtzmHPAvQOipy83jx3h997BV3krYxToNKDvOOi
j8KO8mgRznoIkBLMC/xBlXAGuj1rMBOHKVLDrWD/z2vnm8oNs87A/2n5z3ck
zksw4XDmN4pmgVg3jXVuTJAuJQKYz2BiMynCesY+LUtPxjyRkoYCZn9pZDXU
0zT+M7u85PSqBb91/OJ1+fFzZCkxmgcl+TUyCSNg2A8+EucSdpYQHyj8rRLc
yj8j+VHP9XJqYJyJE4quVO4kP2zklcQGYK/ty7zcGaXCzUFKXBlXMPtld8dA
twkLW6ZMyr6ye+NCy6EDHOO5b1jkbv65Ym7jr5Tik8+B9vZxhirdedtYYCGG
mrsfl6V68CE7/cED918QVUz8vq7vf0t+vxYaEFeUFynVnp28gUrrwg1HlIXY
tCGw91ya6A9BBbIx8MWKohPDJjqeeWSzXrqzRCZvdqN3GteFTd2TtQDB52RD
x4WrfRAwJL/c26nt6HpfgGGNhL9+/BP5/PMcODEfOoFVb/Cqu4M7EuDpnglp
lEznagu/yTbtQP3Em2yQu3i20BYyVSyIj9q5Sr3tgtFhWT6b6bz8iQI8HGa5
PJofSx3PFLcU63kTBZc60YRoktivz5unYRGGk3fcR2RrDXVo+FH3hvuN/ELg
LyE+HnGSTM/PxAi63cZ6uwb9R4FMo0TuxObPtjOe1Pu9UaYzu0Jn5vCVlKXj
wFP6N2005642wC81zhICRYP8WgnGmpC/z4OyVoxJ4/N4EfYVeElCOHgxaw85
n4xWQObxFcUNXS/G7e22oZJiPKptnrEObqZgtwlx6TkoVmGQjXRF1c4bzg1S
8+9ngCwMwMOSunClYTXodbIUQBZcv0lRclAJTvukaY45xsuQlXR+ztHtxpl/
MegTuVg68gzLo5sd1rXxXHiK2UXBtE2VsedgNAbBaKdPOzbHB048wcOsNtOi
Vp4giinWlGpFYhuIFkNVZxKv1XZeDWCF8uF5GVD/4SCsfEfAoyAfveL4+nJl
6eU7ZcOTqyWQinDLjsTn7xGGWgWGAv9UatcAhNecbG7CtQgjIVb6YZeRhZ7N
N2+n3dLYK302rO1DLRIaYiYTFNYrbr4Y87erqYyxu8/boiEezuo3ETwD0Vf8
+eiN9PxSyB7bWtLzLWPZ6An9waxqXZigN06JVH1EVPlD95KMS8J55bALuN3s
6Tp/nzu/L0gbnbMXRLeMqtlYtEIWHotw85FkPHaW0oX/u3Ta208dGMluCE9x
fHQZ13j14b0iE5e228dufh0Um5Tkk28ouwpwUaCjCiBco3Di6oingdJ1XSDK
XKGoiMzZsQYwjRW6U3STQvOrRF8cUEfvA6iGcTV6tMYOJ3b64WsCafysxhtR
2RRunzBF253JNdznZumvemOdkvNvMTyNPaFVTRgS6W6vXHcoi+qm87Fxn1n3
tfx9Fkza2j/uGDqschWS7F3qvqD10jy0q1koIdQhZF4IispVLxHF9tgnDYnt
gRP9myRIzeCHHmMU2tt+YZ3rnslu9U8UxMc+ENeh5MqwD2sAHmfHbCA/s2h3
+PW1W4vEHtLjAsn1vw2JIs2qqD8hUBWt850BmamKnRwgpHx5GvNp9Qjl91qa
DvWImU/NaW15NyF8i5zLDL293U2Kxc3lTPBuvfMia5XsrVaBrKdxEpjF9fOR
0Zh04iVqP1jEZGwLBE3aAqvneERaddwlQOZFwnrzquGqN3qvpu/P6o79i+2O
ZvxHyNeWkOwknG/nJQWQI5SPZBVoRGYkOhO5yfanLZYPAeh0QnFUTLGOJ68Z
eLK2KV25FoUIrfU1dmkL0WuCFBrU2tDN3gosE7d3woqleBYZ7/T4ot4xiGph
R7yRHwlFClKCdow2OgjWPwy82Twlj/D7Vz6nSM9QrMuGRhxEldn3YtLtUncN
4g42clcBSS5XueaDD0T3T5lIafKj6++NU+YWp3C7mR+BfmtiSaNXKfvGc5J2
X4ahxYh/MscWB9eB73vBVoWAIznXOxftnjBP3SbHPrCxH+jUhj1O1prs4ZRt
qeGcw5oX5KWSbDfdJdefzeItvjKiOYj+WLV6kh1VkUB2V69o83i5kdkNhxIJ
zsQbJuMdrt0PJb/MjwGAI/UEPiqwEAzGv8DFu1ghN+Npn/toCoMWGCoActpK
wGXVBcx0E9yyH4O3B5D67kne1cBj3IzWDjUJn/VmKPpUTcSfEefl5Wcjlr47
Rscg1Y0mUnOLkdmcd3U26jfYpCv/YRlse3CRc5BRWKV8CbbNZTkRi0y6Ud+w
PPKHvrqieExFmVjwZRiSPuI+/EIOQxVXERrX4unnx0VdKsNyko+zOyNt0DPo
CKmYuNg9VTTBLr0Rfg2jwc8PozPw9J+klSrt3SJT9KzVvZg949aPuP4SVFdb
GxlzX8+rL2rwt5GQnJgPj0qEz8yfDVSgjIKjBZYdJrRoLsyITzuCo/RDiQFT
XSuXwwHHjP62be2ylUumyvnYbOSp5goRAuB6WPnpphehNIJtSC+HW4HM6Kxq
AATTLrfs9y+W1f6ym5xchhPinULLp28bO7rG2yuDjVQz984Fr/837YFGjT2J
z5sLZoG/W0WlU2eL2dtYRybFIMb6nlh+pI4AhATjCbtAqpBGTVh50KBv3rec
JqT+xHz4Wy7eePX6uUh8G6hTJ1hb+M7TPyeLsLxfVFuvQnotHePSq0h3zWQr
XecyHn974Os2l5mzX2IpREIHM48SZms8XCqNP2R1RSP7jQ9M4H4LejEZ3AT3
08U1JwTMJIFBLbvv58kESmHH1b/RRBkK8OYAUUu3SrwQ3VhXNGDpvZNmhxaA
V0BE2vwZtJYbwqyQPNjvOlKOvQHBHnuBxpzi/TJSXNrXwhTF0nvdF1u6gRFu
dtrLawzjrp/j9NYdZsdcZnsy4cCd+UaR7UdHRRXRPlEkf8KS4pxcGtwOBJNM
V8gP7Olmv+7MCHAmpHbHUSx/VtrGK5dyhyYN6wJuH1yaRyBb/J7jMWQpXSzT
G2TPvKC0qUH8K79hd5pWBuFVcDETRNl3ZVIfsnXfcoCTyDbOTt8JI4HXQrpy
TI0LfjM2H4P//OmS/RtXVSVqDmvSTAqXUp6ydzMB3DhPjwpEzXdBZ2IVRoAr
IPkYlDTVmzKuk1Q3v/AiDjLIuysKYi8s+XuWiZjmIprGhsi5O4bZsx3d1Lwb
J1Nu9oC7F7+oXz3O2HRpg/jQOdT65xO0TIlrcQgXgl0m4c/Y9GmJN85s+DaA
muwU2vdMuSAISS6awXWs3UUeAr+xW6XxeN7oVI258NevxmlT0h0MEQ5zgVcw
rbsU+hu8s7X4pIeM4Ih4S0xmS+GJn/yeJXe61XMB3ZgfRO+KvhOXgSPD6fxI
vzJv7+WdNJwxOEhnzU8grcd8qgwUcQbxEh2ICJrU63nQJ0lrEfbm/iasRkbd
QvyYgl+FzJyag74jUESsVOcLPuEapb4NC8D2F+zusltLJX5yOvkS/MXJjux0
SwO8eDmOcADufmFZ/HjgoFhHfpkArSh9z8nzUw+hgSHo+5oKpY6lCH0dkTeF
Sbj/Bibl0t2duzsZK4P9K5lwO2s5R9whV3LNOaD/bsDU2SvsHhiz8DlJft0X
kn9bDNsiECqIMDcYMvDUgTYejiB7h3QgiZfj+zhBNnbbn+HheWjI4fWhUnVu
v59FWnVzCiHTfxwrdmpLZC3P3YKUZmVC98Qb48ZnJnDJ7zvrtV+VTLX0XeUI
DjCuI1nH2n69fo5e6S172b3ldG4ltVpFkj1sG58r+tZfQfUa1Q0+oZAloDHy
Uv8fuTeODFK0pQtWjn3Fe/54XnG6kpeUNgaXcfC+gBOJbij98pVikkpprOq/
roTrRWSpCzdRDdegtmBYxw0fAIsGIHIvFv3B1ThVX95Ljh9UcLhBm5PbubBd
aVxZFV/bAWq1Zr4X1q4wflvWUn016VPpkp4Km1X67mecIuDwwwmLLDkOeLTR
Fm1OXtHmdsuk7zXsmVRtQKYxlI2tIPZ0v2huN/wdxEqKoSSr00w+Ezl/d6X/
c3pew0MTppiXlU9KBV268DQ2kTsZNP0J+u0XxcOWaGry1ydrspvDlJlG3Q5I
FJThn4WrjdGxCd4p62G7EZtf9F8vLPdYg1VmiMy4rCjDysx69GchfCjQ73DK
t//UeS7YUgtZZYfs+eHjFJwTbnaZ8XEuKK36FJVm1ZOEreFy9DxaqB1o1P0N
rajZzJrC9p/zycUrcSccZT3kW5oV/djaEu8/K2ybmQXqPbs2lpB7/osZ5quZ
C/E9SMw/QCTR5mYPJSS139wpisI3dbPDzyAZvaeb8usspdsjTiafUDQ1eZt/
YcjJn2kGcQJT0wBoepUvwtTgNZpMblox42RWyqe6a+YQQatwGv8kmhrCwsMf
InPWwGhuXuSV1fv4Wapcl2V5hdwCBkIltemuSozrzcQesQYN0qQwJt8AifYJ
MaXrJnZnQ7MKdUUSfSft7WtxoaQ+2aOYHfdW1iY/2E40rtciHDpZfkpRY7g8
vKjgG//9AsQgyc+h9HHRwewZNR2FzDbE2h0DPGXqzzZMEw8m49sC+fNzua9U
EXqDqxvKY3wd9A4Kcv7mfJQovhxfmwa0j119re0IXxCUjIzVjPrPEYNCTaPz
gHqIXkvW8Jv/s+fQk/OeaNPxe/PdJfes0zdodVTl6CcR9qfvADqplAXXumvj
l0ZdgPu6FQH9hU3pOVezHw6SKw9I9NZFVm5Nj1QU48mYfHAn2LQRmWIQBOFv
n5cDWjVeqU2J68uYjKQ4witw5/m1j4MXHYTgf6TyZYVXNfGfUTvS1vY0AWeX
c0GGRebinQEpGOCVd7EaXC+JKGLZ7/1EvWmO4FSqu6x9ST2frkh/Q9QhQP6X
dUc8jjzSnaTQ7okL/CVi9kW3hDDNttNF4lERzTQjZ1w6wxpspTdTk6wI5tbv
u1ExTtzKriASmsABXrQFPjJc1MYHE2b8qcaNzNHs86wBEjszj9hl3qfPDwq4
KBkGMsh4cqfu4xYxpTLiCnoPU1BGpN+v+M1VzlQVxSiuTZF15l7fQUmWnGG8
GsOdPvYzPuuj3k+KWbFZeUHqRlyIfrJgEoJSo0t/I8it4qynTRfAOum9W4Wk
vyIaQFh+BwzGnNGs3TnKydTQgJSGaL0QE0w159CJJA/QR9UyRoR/hgFPamsd
NEIToqVqdwX05UsDLyJHg3WOh6KpfdTBQVN3KdO8B1Yf1bG8rcVwh/o5Bq7M
rgW0+Dw92zQ3cQI43j/ndx/5B3WTNtTZeJIoxcfHOvM2EY72Dk1BjU7oNC5t
mWNSzpZonHY2xJm/jwnoTolnTNDVKhYKXJALKo2dl71/wbS1fQ/j0C+wPRxB
inExSJWPj3/YWdYzcIlYzLTzQVVQ9lxS+3GCTzlvFpMdtIrQcuLJLHWOeBky
w87C4TnlNB1mlPS7f0uSM4Vs17C2z/tEmraVoqRmAV3suwNHAEQYAO8ijiL+
scc1hBT+tpGX+1pUIPG40J1axF+Aze8vF2gNFjsj/5kQZVaVd12KDD2OOxEz
8EtBxx0gf8R+tZ1nYqOpiYX0covA4WpxLYuZ4LSPLLQSJEEY4IFsgWUc1nQ6
NBas94zQXZE06MLvj52agG+wRTvvKgMMWTQ4SLH75VHJfb4ANcBZPm4mcgvH
INIXDE+D5EeHub2Ma+/Xm5fHpU/CZzrLqOji+OB1JA8/sA9h2bcl9sHW8/WG
TKtcAyLZxHI2sc0JO1q5tjiQYZydHD/IAdBmm18wYx7hmuV3YTOX/aliO4yX
FZG3zsUlsUxt2T3RiSoWFoHthygLWRGe1UcSPCDc/LCdDvvssrwuisL2I/cZ
XUWM1PvItmsLHELWvkOEUR2sNweBXVuUnodMoJ5IQgF76brdK9eWeO5/bssY
bjmYNfBaB1BMPtCRVovm7lTVI8GR03xavwFCB+vJpVGotVmdyy6ekPxSLzMR
N5oL/7a0HqPFJU73SIj92y9xnHauuApb5IbO4SZeddjmJJLfLt1joSRdt9d8
SniJ1Os/7E500nKEkqM93qDKlVdsvUVUqrYzcnTyI5m7IRnhTGlfjuHvzGgZ
Pi6hmi41Yvr/R43/W51hVsH75KcjzRdlOLI8+i26NY5uoZmFYStPPE73AlQl
gETC6ZuzzbJelgB9q5qkvO5asI5ad/wesByvrccYCtJwwBkraGGDmRHub3v2
TNd1Pb0CjAtc3Pir13BmENNIwOXX22z0BPDdQy+yD4XEFu4w0EVXhizdNksy
CutRkguumwUNsQ+oNkDVok4njviRa3odNyNELAk2zTH77aZ5+EqVKqnPgFKL
8PFEtombc9wv62oq8alyt1hXfab3/9X7Tprxm0szei+YQPkxBpeVjjj2svsv
Fp0nHvvQxZt+adHuu5JbdIOy7hv+LEpzBSEbWnm51hUZu+YYqcs7H2i9IvKx
/NjbQnjG+tRx+m6/nSGEfxVmgbV83nqdQmlpvm1YydNR0sr9IJt7E5PD8M+5
U2UIkt8hytC82zVs3WUOih//FtoVNyZuDrnvApH44Y1uTJH6ruPsTDyR9CaY
zMnoXdvRMD7vwrL77SCDVXCjcxx27HRAiYYkevC05OKKchTC+tzm275HjlHg
JIHlA32MAhgN7ShGkegWDz3C9WaxkFLy2jYfnZFGWYjlmpNUfSbvertQuIV4
/DeLCW8zCJ4niXkWcoc/5vBH/GEPV8jrM7JSV6Ij+cFOKjreloW0ZTw41SJR
LdFiHWDPr22beBdHMX1yBoqgLyaG+bGRZgS+9GQfu5qgHfz7wgLdVyQotS+Q
1dsj45s/OY+HldYKsb6O2ZojEmCq5RBbc+6RDWUWTNdnaL48TY8k3WCemk5Z
lMaRFtiVDoJ7OYt3Enfpqe5hlfKzcVT4Bg+cU+aLkS37nEtrGKttFmlJbBbn
5lMT6sYugERR2uQPGXAEprwoxbHt97/cIqRIDwhJN+yQggEuBpQVqLOS24Nc
uFniG9XPuQ+dutrBok7oxGdEJv6HuN5MAWd1eMz9Qbr6LO8x/p0UEkVUH+El
vEY+b7sl0oxUlHAl6zFrg2Rmh05+d68a+AEhxaAh1srfanh4Tj0if4Y3JEkb
PcECEpeXGVnukl53LDoOuWHW7Qwqb6M9/zxoisCfyFy6eils8TW9mnfRg66q
2ONZwJtGeucZYIdUuiBA5581vMXDKZdWD3UdqqjdUFNk14/3t7iX7jGPMAub
WwRbTmCKCxcwmu5Hkl+WqO0EE2k2yH7dnw/Ttdx65zbZrdMSpjf9MC+ZdLXv
2t/v/1WCYczvzwzWsV9aMMuIQA6f/f3JQfL983y9z2yAAkxstzpZfxP6nlVQ
Ao1ZMLc2g3HmvGXgZ/4Y2O2jc2jsTUDQSSLi0/k5GefVsU1yPuZ3+toayveF
k7SqOzdzLcIw0cIJhkJbsx+UdvHIIFc3UfdCpE32YLjTC5tKl6ThOsXKpsxC
IV+QSmqcPI74zdT2oZI6Fn6xVtWrB5mjVlzjYHsrPQj73zBB5BiwmZrVDExW
vgbZYwGn76zGgtVmAFp8bV7I5OHX7Yfyqs8TsBk+2HmQ6Y1sbpam2nPo0b9G
z6RrMqRVc7HfNXces0DOqAG8LE8jAv8MZMjW8GOE6U0Kw2uFD/ZuGpbkEKIy
kUJgMdoJOSABC2XwxIOe9rHOz6ShUkvNOiarbLZnAhyfYoQEC1TF3I7wY4xn
JM3tjgyrVLaHOj3YDpeeuSEMhTgc2U72w150zaGuysX8Dmw0DktVaBjOEFwy
fhFYAW5tthi9rFckQSraopvk8sjr3KOztTLl+dZaUONb0ItifzCct+q6bGtA
a7Yoi0OZK/Q0YZv4dEx9et8T8GXfw1HVFYAfFkYKp5ZK3U24Cv0STi0F6Zf6
luC0W/5PT2fl7NGOyQmw2v0MgLA6ttNYclKdDLbJaAmOTQ/uFkXTu7QyRl91
feyhduzyoafGhdgbtd71tbJiP6ZL0PSIT4ti4WVGwmr+Cbrni+acYOU1dROK
+ihfupWojADgoCTa7q26JDhEvpEG3t8PpnB2pEFtsjsJ1bOM4EFWQqKjdTaR
LiyjS2f+Rh3DHC34YCvxErKjcNvBvphGah6Dw5t7cn7IW/GLrQtrJIpcLOIn
nvnHcEbCx0WiLKtqyJxOwcBMZWBk34kOAkTLUhkN44whz8S9u72tu9SVa4SP
Y1F2DI5BCplYjYiSuQFfHsO9lSVnFUIUPU+0bahdxSA0HwgXMULQYLpnDd8c
1Eos8+wqhKQyqf019TEu7re/2sFvj13vp0nxWLyXKehMYDt5hzWVIYVESNv7
KO0dRpIOkaLrgbZjhPOHh9MD8GxgotStYcL/BsFMUzpX8rl6O19QI7LB2MYr
CWhC+TRUN5LCw9a5LWA2p+ZgpMsJDrmZ4N/wmuy+4bjO5tkn1/Gt5n6gUu3S
fEprT9TfKrAylD9oXlnc8/RxBfC0KBCNBWDtUz1bm6E/AvhgVcu8Igi6ytLx
PPlzs/qdoAV+cIzZe3FomCqOP4FKVZAjtzl0Q4PYnnLrkMBqHgYbjJs/5ZkU
zUSg9J/XzsKKBuR11VJ+IAzo5m4bAA5do6dCamF9XZ5XpPT3dZND/h5nyc51
HoS5NNkQPkB7SUt14egY69YQ3NlNL5AqV6fGGjdsIjBy8Aw59BVxyN+D3VSO
7eCRabzwY5LiAWsAIq7eS3gyaWIZUbtvj0lrRO7hU83tglSpXuwKnMyYpRgv
j2sqsfGlIHS9jqAFGJo3EaMD1j4TyTD/fCjmNgG1I8slWuU6BwLadq/OcTRI
tMRHUwFPOnHLpjWuvGQKQyoHEDphoWyMY68MMynkotPhHaBso2xy95+yfBlG
xTeLJ90StOb63dBmqmzLS1ugq3NR6qr98nQjNRI3hhlYm1iHKqmndAyM87Aq
xeznhtThtZzRPE+NZdybe12JwhXbWiLVQw5wh2CVNoqavOM72fUg6cng3Dck
uL1rFeR66sJVV6NalvutqkNH9NDld4x3IFnOJGBxGhOg4GbyEeBvKwCwgTVU
yeIEf+avKCTJZfVS7h73f+2vvJ/iF/JDZphexI9qV0fYH1gBLpLCZ6FZf9J+
aRfHhWz7536/OZ4P03/vFCG23WZqIIEmWIDr5nzOUK6FhNF6a+xHs4q99+/B
Aamk+hMwKd0LgZLSPEBTKCklNn8GH3CqIrTcwpfLyIQYSsZpL/D7NkP3kzje
S2aPitwl0YAI5OBJwqo6N/izpe24910kVKjyfH6NxOTnPNZ2CU52PMpc6Ffq
dittgzcXz2ZI2LMfaQlFP22for89vYxUkDTqaHX3kU14YdX8nIefM3O9kuGb
zqCPgUeWbyjb3iR+FJ8JmX/gPnqaTnDwxOGlJaMzOAC2V44aRUv64R7FpttT
qnKXGx3f9oJj9iyC0d28joW/OuPj8rXz9EHAPAHHzaZRszSzn5Ml30QI1tVr
nJDmuVFfJi3thJlWUvMEK7/sshcUvXsmAJp69CPH6hRfk2f2PC9ySd2+5Bwe
esqkKc4R/LG3q13lxZziAk8Babb0IDvcWMFrkwWIANF5rLMsjuCJ7PWoS3YL
SzqSq9AMmOV/jtfV9sFD+ml85EzIVPSizBr45uy3tcRiGZcFSOEBWJE1yxjk
Ou1BaJc4KE/0LTrH1xy9F8PjkCpH8S9y7B1/h5FzYu5DHMZZJcm89z3xszF1
ypEAkqOLymAUXyggHQ0unUmtDTgJdCPERLB3ZyzZ4HEqd4Y6Dhctnj6tJEyh
fqcrhtYlHQavDk0Z4P6OhdTm+PhbY7zUhtNvVaWBA1GRLBozKXq1aMLnuP6p
pi6xp7FTSTa1qwGYwjbSyGdGC1LR0RJdy9Db01KUS1ENbWwyVclaMubLsQkW
0v4brXY2KpbUlba3zCx/zdEwp2z3ulpl2lsPTlEYB73jpyaxSdKbaT1w/Vye
Fic2uzfFvvZwgSY/nmuZWyP01ZEYhVyjLs/HiG0zjNUH4CUGrC8JzbS5nx5M
g1Uia2UcG1VCvqFtxim2OFw4Bce9Zg53GGgJIVn1k6nw1QJvd+hTAZ9I4Idc
w/BRs6MLUgiE4Rg+u0naKaeb3ra+rt5o6lgi4hEyivf4qcS45qccAQYeUE56
iP05yWDKiX/gZjgB9gmXQxSRlTaqdrtTAKUi4R+ATzHqEBx+4V/YxFjxbD8t
M3wNw403TfwKGXERh5vPEvyNW7dC2z9vGBLxbcc8/NwRqX4UWXATodiELMex
2DXgohEqFM1a4xhkp9SLIyUan/7a8WvzLcMvW4JL8xDh4V0u6YroygdAA3b1
q1xlqZGyDvqotmQ22jkmzJ+ssMFVQDBPspVDFzCUX6OZyIaPTsjBx9rUPpMY
44w7pEJO7dvlFkd72+ZltnFcXq33fOrR1OkwQkbPR4uOqu/kEuBeB6uhRkf6
HRFJkIHt4qJqkcpalqWDmBKtBD1/VwOjFhMEtByYVghwMPNNTTmscqh1Rg0W
P+ZnFgGv7cvHklv3fOrWbwSYXMVBrFCqq9uNE1mwJQpLxeaByEKctv0Zyai5
PGER8fSuw/JjX+EN+5Q4YiTOiNMc6TpF8FiPoYQF2Duj4zNgVZ0EoqHf6FGn
EHEzfq/rgnWv2jtfMF4jp2vcFga8fziCYLYNy8SylAPRFZGuZVw/qCEnFKj+
fQAFtiRSrt6EwH26fSvCvBPaf/fNo+t3yVVgyA99Vh+YRlAMKI8h1WbwWeux
YeR/BsPZH+bFjEWRFIqnufaMSov2a1DSFMYW3aBPejP8urUS52umc9zhW+cY
tcShlVMExmRaXL+7ZyZNmsMAS9Ew5vVddhhmQrTVGCQnHLFQWU1Ct6JIdqUr
wuBGMpvLLMVbf4HwBUjgWdj3dY4LWm7Pd7uf6ib04sgMEQSHRQM3FUiBjRIO
9INx8WR03pXgFbHV6M3JQSGVgWEnl+wVCCYwhFbNruP2Lc9doDyKk4fgh3w3
y5hMMHOr19Xx6tN5vPKgHrnzegzELMViL4lG+rYoxzJ+oc65OxSSwGdps+Nk
JjL3Zgnfl7jw2qymGr6FR7bKzn/w8C7xGZnK3Ls31QbPlLt1ns5nmmZyWaUt
5HsXbmEGmEC7I7YdkMhrCc2VOQhM/CMWS4WZ0SZY9GPXogl6PVT4cCod6CUf
TNhYhGVgSTMUyLX1D4ybbuHMnlTCH3uAljfHMA14AH0yo08XB2khTrMpPBu8
4BscuO7jRE0lPYvUsE/0cTUZaiDhRpWHiUNirf0aAjvimco+czBrcBpWQvj8
1DfObKU0ghWXryewwak5X9wA0QzmiHIjRBO5KyfhaQPWzOVRUfO5IoBhfeqq
x0ansUGIq129OvUHJIkA/kAIVJOwvYT3/SemoAXXaUepElpxAFLgZjzMFmOa
VrL0XOt86VGC9+GUyQa4JBLt4cLR1CrMU47gnNTnbMRyfMPeEuRbDTQDxAJl
LMFrWLPws7Y/qVs+mUA6d6WGd3UUI6MuyWoNTGOiKI1qFhbul3YXmlgrvDIB
/fBYMZYePerLJXY5ifdGfvfg55+mE3rNXNzexGi/G7NBgS1xbu1kXXgLBM0U
j+dCE9JhomAi6ilWAOAWarDHA8Y9PrVYKhdUU8Qe2e4TXAd8fQQXfYiGS2h9
5Z6rzZWucJaa+sYeM/iduWxTwWeNW4NmT40jfhAaAQzj3mR5Ty1dQFgTvJgW
PMsb1Nw45OmM+BM2h7D19dU7m43tkhsTU+2qTLb4+rQdKkOSNDAuWujvFW9L
6DXnwvZ/CDkekqW6nEZ6JaQvzYpe8Mv6FQNTnA5uYGVnkndVnyE5JbJibM99
2nRJBtq9NwsQSOIclV4VfnUofoQB4fOSSnjfijqNWIu6MwbVx+MEK3sPV1qU
xgUpRfefPMUcbofszhVb7ed4O57+YkwG5n8ry9bP7QyJH4U43sqmkCM5kyg6
cDNjsxEKiEUSf14l9qLR9V19Ssuho6s/LcAJ65IGoxzU4czTACzftgC99kEv
XhF6EDo6kUJ/8cnNSA+1UuVMCqn3pW+kRzrP6B4dbPyZ2fjhG5CjHUJfEcdj
0eV/JZsGo0NmTcPV7Ss4HtWWFRt08dgdmMBtuAE9N745LPlaEzWJjTjjXzF2
dgpPUxcbDJIRqY1nqpYiHJVkvgOabSb/hw1XK7tOmZsw1t30TIJNFgd9wej3
xRQZeRAyNqrJb3dU9gMvuDKS2BkqC7mmu6jMwX7/CTyB820P/Ggo62Ij+5Gg
T5lw5qlijFLhqvs35033OeXsrRlUpIEi05+e57k6I9EVp0sbV00/chf5YVLI
05vW/lfQ1dorNKelv0tVrEOzBTLFtoN2vYYnnraDkLuHsXkWHznh19o+z/xJ
6hvU5bUAiECWugehRVG+QtfdIjqL9JO4mkzepcjdjbT9lfpUI5Q22aIAA7E8
tNiCXSG/EoPMu3CKvszwu6TR80ZKrjWuraLj4f59DChx8nHvIID0VkYBDt6P
pxW3AHtJa7DH0jhHxudRJz459IWCFD+aEXy2hcomeljNpoF5IPnKjNWrAyDB
MF5JPxJyhzHIdXGcTmD/QccfH6yX2kLATW0AWgw5pLcKOMxmPF9o1fG7ygMs
dlnmXXN2+slPa3iIiuArF8vCc0blyhTLFpDNWsCQpsFUKTg/YOghpE49xkHb
syEGKsAOqGaxH1wAWeDjakvvZEhvKMfemXQtdroTNuYIh5b+yCnYg2QQ1cos
I5/506CYLyQt1ubqVJunCzNBucCmBmEM39FIkEtXeB7bgryYHUXl7R5aMAp+
wtxaNgAp7wcI+80tJIGdgcXrcxHrU9f7chDdfp6cIXPaXorSY57AjbJknDV/
uWTMDxYzLlimp6GTOBG//R9/rrl1Bpi++PG08RJtr90QpJ4E5k9wy/sSSEZZ
gzNEDwZGw/aIJkvGSh2fI0qehveqvBvAPu/p5ZbG1jMwg611zez9H8DTrYXi
BTqEl3hw3/CGPi2RmPa4fceAZl0f5fmNdMeFjljPs/ptvf9FCAxQdiDXQdXZ
mzJf4mLSWwnMphAdnOYY6+FKenubdTElp/5TsQd0b9RwdTti0i2KN/WKqmsC
qcom5JZzT85+VHaEP1FoAeXtW54tlWcLuEkvXwtqDZuISQaR7snITNdovYQh
7M0a62nw9dozF965wLQ4SsiKgUYFKmIrfZ/HwQSz6+ieGX2JK9axTI9WFAvy
qRyXMMExCcj0aVJylAh/F9bSGEz7RHM6ccl9KNXy2AVe+h4ejg05jlItWD+5
EjF4gx7vbOip3QVxISnhYehwLA+MHkXCnAaucStuhs+vx0xNG3pbZhiZzNke
c9lW8NwbWUw8pibtbQMzL/ElGKDWti0JzRXGiFz07e+mzdlPvEtHADv+A0bU
1i4nWolwZFD92Ree3a6T6lpeKi1R4qX88Pi2b03ITMy/DrAI5jycLJsrJGQK
7TbZBJ0+btnikyaUfbzMFo6qW+4BmPdwb1eAvTN/ryUnW4p7hZfk6fz5LWdK
uY0YZfd92/NeOR/wV4MN2WojKTEL8sUV5Bsta00DcOLfWJxiNJwrOo7qliwA
IRuh8Fa3z+Px146aFAxes0lZDpeTvvXMJn5F2eTEbyxtN0NCarz4k52WS7HY
Uz1B8SwVYLhY1q0daSExZ4o4QIE58P7C+YAwp/87pOKSbnt/3Z2+OozHuQs7
u93LXn8orSGAyBDny8/lqwGG0R6T3XTIVpsLL/zuRKrNyOVyWSMwXiZh9AwH
z58pJ5icwNKDCjbA7mch9Oe5V9jcY8hTTOVje+qWlMo8kfThLapkkgYgIK5K
fgtRfuz1EWFFYr6OBUOCrVApPLHHJQ1DQ2RFpZz6rbVgotdK0rF7rusHeCTo
tExPFgNFBtCaI+OSssbryP9aszkMz118JCSPvSXzoSyaRK/OdmbjNrrYhvTn
oNtta4myvKI8zJjDVb8RletxYGobMAoGRuCy6Y5rCgJGCc5n2VT9TaG+h6h4
hYsgiP1VRv6AN5UOcxV81s4y14jH7qKtkqGHp3MhDfFHbTUjo8FxaRXptjLe
u/u3drNXWJCoiPqrUimSYt30aLKtTcsSvMQgR3mHFxPkRXACg9X50/BfDusG
Squr70eRkJyw7kPQiek7bVNNGs+pUum85oGRZU6HQYweSxOI8ZQXggvQzw6T
Pr2mdMEHj8WwUiBRw8gaeUNCqLBl1mgdZn6bLGJHS/WuDnmEnIBegZ0tVD0s
Erk89G9wfwYgFwKMliLBCGZ/+fMjpYMhCYE0Ke6PEOt0HOXsAzvWBs+dAgIo
tm0Axpem+rH+71m3EjKrWhitpqFvw/2NNyp5+PwZB7jPQ9gkkOeo/1MHkNO1
/PnozoLCxW+eCa+Zd1q+RAs0jOnvO+gC/KleKIu3M1lPnOWx7c4gmW8Q7Bo1
XI559g4xZgrLojiV+ucaaJXCWaPLG0hEtt30k1ukb9RlO6cIKMnIruGM5Hnl
ai7/ahAcsRwG4SNd9fjbPzZpocpkEeqGvrC7DaDHj8HP+05DsHm2OFIhL6Ul
r4FqZPlf7aJ1y97EdWDW7Nr9oRVxXglWtAROevGEog/wIBlNi0ZkOlLMIxJ7
MJsPwv44az4E8Ng5AHyqqq6np1sc9uKJM2e62xpcSB93HxS0+6lXAIm+arH7
CWTyft8WtBBHx0dJg37y/QYYRitEXpsuYV+IpBgTqmJZ7/3BPAWkwjhHOoj0
sRHrgubPN2T3LOyXX8GNUJnV4z8CNceX05iu3jxjCU7mzZ1svo09+fYefoYE
2MJEbJ7Jwv+lMx3BLkiH0oiTtHS7zRY/ct+nfELMlqh+8AchkZj0GfqA9KRn
zLJLxpLZlADzAWjAr6vMv0NxbpKqBnXIfJEf2FM2QOOExP+2vTqeNovlNNPb
WZQP4FzBpKxuoppzGiiAeIDybBlwu40fGrRdaX1tgqyEs1KmDfing15R1sbE
qXPMriaqq3ASALnZ5WYse8Cqf44cR+HI1QwlpYNv3LLCEtqwMKQO9vDk5Nyy
8aBP9yffe772OxqBeNChJEPGchR0skbS8DgdC0YalrxFjt8ivE5xFD1zMMuE
phiZdqR5NjOLkzuIzGfCTW+B/Eq4bf4qyFdElYIoJ1h+OXmgT7hyvcL6ZgcC
qdahsZDVkBvcgy9JgRzFa1VggiFznxd250k9Ox+2HNKDmAL7ltszqJ/EZFB+
F5jlpxLZfBjrkPLOC8pW+Ff/4r9q0CLPaMmAd1C23oxYuD/RMEHpX2oqPwei
nAdxXx9d6Fv/TICLI6ftMdhBo8RRVn9VO9jIm9TkDw9Z/4pStCfCv2nby2Ca
rAPCoBPeFowu7VGBzmf39N46kqBv8rMELe803SbdK1/i1xMk6gbpOgVrv1Q2
ulCP+8e9PwSSwGFE4HWSBPcn50m3lc5zWrxCZCAzwkSN/9zjlYarvgpkJE8V
dW5veiO1nNWu1nG8HRLREWvL8r1lgQsHbVZ2dYeVfBDfMuCTIAaZbwM6gyds
mJWoStpDsEudG7A2HtICLm+Oe0f3E/A/w+Xv/mIHRUQ6vCYxoPfMhaolmGjE
SU++9gXf2fH47dPNRLIi7Un5jq+vaiGq/VC9o+gjTd9374H2Xj+ZGErXU+WH
s78S5gC7qmqQ7LvkK851jW4Hsrr5baJ0/a8sxlIBaA2D3zA0x9nVvrGUgYHP
kjR8PkhjLlHImcveYF9Jd4DLGyhYv9hf6Ee0Isbl+0mYqd/QEj4Svm32lR2Z
Uv+zdFIEQPoQlFqe0Q51qQ9NiJFev1Nd6VZ8fKXUesIHFbBmX2I6IX8vsvSH
T+TziNn4x7Pmf8CTj9U0H0NEHky3WhfbHHypSaApB4x4dZ+R5LDzzZEjukkj
Nw4kpn6lLJMtjw2PDOVLzZqXWZD/N8uzGQGcabjdAtUEYr8Qm+A7FXhm0JXt
h/cbmXb/M28cSuGcLCu70EXSDC9HxI2nCAfCKKo5AgmoBIclZVminiqGu+OK
C6JoCKdr8+HexVa2mAzjNXUHwTuIsOMlStJV5N7DuhiOdpb4XlV5ve6eyONW
LSliOnG+lj/ZJ10LIZGpVoBrW8P4/SNqu0yotifXmqE4IoyYoaVaeaSzbb0h
cIXPB89gvHvy5gONyMIF/55lWKlqv+wAL1GnGTiewBvJV3GmYcWN+hgH9vH4
vPJ3XDciC0ncF+o6T7CORUqbOoxqmS07eLTh3u58cevk6MeQHjkDOII+qqrW
1lz2AFQVtTLvrtybXV4/+z1tqw+IjhzqFssLpIRq8TGgVaDaCZ8ujzzyJBcL
GzG4x4+WYhdUGWg9nPV7JB10EQuv73/1QNeOb90YCgCCMfpsl5w73I7smcGs
zh9Oh/f//I1sAAo1Wc5y71YUUsD4bykLuFbEXMbhrfXI4mD+X7A+ehMVIKSx
7QLYlqRXf1iuyWZUVYB8LzLINY9U0Wm6i7SSpCedS4efcUWGqozpgS1mRo+o
VnCWvq7b18Gi0LnNhjv8bcNcrKLC//4S+68dF0iAVVnFrMTS6yodsZBoTeRe
umHdNVfqi/utAs0vjQ2fXMJsZai+sHCQhhyo0ImIIx7gNF96lCb8vFpMGZcc
MQVgmy9dVBeljXzZQY6MuRbZ+naTCbIETlcD5wkWKICgRd1JJ6gNi0EMInGk
kn0w702tqqKfdtC7cdUHuZ0lLHeLnrxVSFvkCN7ptK2Xuxc1R0tzEPbELW8i
uB+/tP4Iw+pOJ8LIT3pOUZS/dle6ubUybbYitW3L8l1F3om5JZRBauyvEJVq
4hja49efDaEj0J5OywO0/s9wfLXqHXs23qbz+uKM6X/ZrRVElw8C4z1JIvc2
gKAOMbdrrQSaQBWPw/T+tFViTZWjkKfKE6hrl0yLn2Q9nzGUHnyJF8QOpflw
i4pumj9SMcdCON26VRRC5UVLLeqLfjUigsLV8V/LE9LzGWYGm0EsQwkaGsxv
+TIULLNLx5S4tad5rw0VV3jLHm+cKN5gyIghQtt8b8pWtYVnXeoqTtQFvF8r
5F1oF7rOtgGpvLm5jQqTAJFkxxRdvqXBO2EAI1/8UpoFnSnrKwjPvxvoF3IG
QGQi2RcwSAu5CcJVHj4LKYtJ+/Y/aHESVLHOvyDvupvMFsGupdDa2ZhhRMe0
t9qPNMF8V7/w7VTDeZRSwUUEZ6txdWt6uGUJFeAmtHHpi9PgczwMf9q+BCqP
U4jlhnyZcFH1dM2UithpMiYbp9bgIeEGFVJGtJVKRWqL5mmwPVC29sWFvrHw
8k3TyPwJk484R6CRCKyAEqN6W1m4Snx8dg6fiIctzle8bsaal2VlSHUSxIFw
HBFCHlUob5+ePk7CmMOzuuxz6xUZ6ysHjCe6Sy477TODidfdpSikgYJsgO4n
39JweHMOoecvDm4m0vSK0Eb0rRF997uXtBRG1t4x18TB6UMCUkWg06Jc+hoA
sEAkVYFbMsBNIV/cEMO4vyiFNma9DWqXsE7WBeWIk8Zdk6mfApXCfFkWu+uR
m1Z7dEzP9mYkxen8yov86SVg3Y0V2bilDkl8nzChy+uUd52v67wdZ2WOl6g8
qvth2HlvTmAi1kcEhLGq63bu5WORg5StdS8mdFKVLbkufbyexeMoRA8L9MsW
YYnWeHyT12SnqnDP0aC6tkY3wELn1WfbWgnH/PEqpd/xp4ER7g8sqti4MhaA
4upJRMP/tJgsoxy2qmBldrhmetIRc9t13MyMwDbO/W7OUGY1mCGHnxFmo9jW
T8Nh5SiKKMnJlCFHMHG0JiUPWd6uBlemBpcUpB+AlzEs3e3XieOdMPE8SBTG
LHmEhWA8NkKq8fUUAc6nm6aNsFOSRXJa7KVDKo/xXOlOFIriZA/kgYT7onBx
KsOd5hl+NgWHlFDxSCKFskc+EKQZLG6joRyNBWoHzolTsFn9KOQWJbF/7z3v
IJsEngQW4YMpxl7cwOkDMhTrNd/0O4EWfBOWyfXy0TmjEX21s6sha+A2hv6M
r3ozvkN4g/KIsTkrflTiVopNdLia4XkmPThnfDRqc0/A9STYSHnkC3armlIM
BP0TALT4XBoXlg+W1uKKtJsKV3l1ld2KL10xCdALurYBFk88Al+99IlZyV61
1WboLAx2ZHgcDrPIDk++PUqy1vlszteHE/UVVXDJW0fnLqs8CPtDAzYO3B5C
82pKFxM0ELIszr5qKVambMjPoU+KUJkxcLxXC/0VMO8Gep6XOMrcLpmWS0+b
5Zk7xrL1Nr31oHOhCtrE2hoYKcH9e+T962noJV+str7wHNm9Ph2iCawccxK7
buj4EW2mLaWLSSloJekv+6nWwcNQPMDquNBlAzd+LusvOLRG2b7QcCTI9sag
n13eKZeYrsnSvpsLEUcW3O2KN6GoWvzekBZmoQ50Wqb1PyEtiaY9plmX75EZ
AbQocViJQK10oqKJ+oxBG6lROujyNkDYl3ClPE4KM3DJAfZvfY2fsAASDKHv
6qcWIkl6n4uM29Fp14g4TMTzef/Y43DC0yvn9ZgfTx/b8vEOpqRdF3pOQguR
Lop/vJ+M5ZqSfvd+bksGR4RJ06e0tLHtaDBWGq2OCNQBhsPelsQn/bi78OJY
VDeNGRuoi/43jYBojdU/1mWhqhp8E6PqjxnZbcxCyyi9KyZ3ABE3u3Ji0fY3
i0rsuyFtoWjY7jQalA6rCEEiuLyvvLysTYSby6HujZG9Ux9ZvrsM2sRr7Stw
xhx20fIhabGORbO8J5osjMbogvfTGjBco/foEvODc2uuva/BpnrN0X1g/kxo
sOyu9poxkHjYnHyaEFsz3u9Zyky78bfv6VlujiJwv/28INsvOiqWKmvviZX4
n04DT02lplloUOOBQlpUt8KvrMSEedv9KeUF37Pn2m/QHmrQe4uHb7Luou7a
/WHeYsu3hLLbaeoESV41ze+0rNSlGiQycTzsI9ThUk8kIF42GSaeO3PJTb+D
gMepsQsEFaBBLszdenPO4gdOW7gXEc2SO3rX1vq1SSAnpP376etJZcxHXTz1
yC4b/EWDYPZyhKIo1gyDwRv9WIyF0AURjIknyBTKmQkELr+KxoFiHiOq4ZGc
5M2AAs1iw4enMPqtRNb7SakcwPs819rvTLHGKI5CDp5T/zgsC7Ba84MVrGWF
pPZV+G0YH6BRKfL2UmnKs+QmoNjmzoQst5uDwUBKGj/aqF7akZNIcFIe5kup
rmgDfhdIIq2yQIZUwraqqcbS2EPibOTbsFQp0yxv+JrK5somxc4V5MRiLr/8
2yNu01wZem2Akfmd5iWt9V3R4Q9b+kCf/AZ/qX/t1W/UpSY4c3qASf7aVXnl
ZqJjrG1XMzjg70zuX1zzTk5EsnCKvY46jAQcIx6u52/rM2XaViVy70rApYVV
GRRcZ6J7iIEjM8CIvAz/WMJjhhHk5AeCWSqPj4xCuAMdym7+OKpPMFsuS1vU
pcErc/016q1SAXYLCSs0vnisKQFLfjgsdGkKobTdtLfx/2xfMnKqOXq9FlVb
1IoHrLqYObq1U4NdSF+15xpPhxg2BjkeUWHddvSixIrg7CK4okiMyBvcMffM
aZV7vmjn3aED+8fRKeSd0Dfxy7eHtC+jUb/IFnkeDzUPHQiKQ98I1x+EMwLu
nADc8JiIvYmhA+O3jLZozUu1DXsNnKJ0BBlFA/vPtI2xNS0v1QzpvYja4siX
zKhvBQ/Ov0WBryAjZ9rvAMzHgLRXQ8tHKGk3shJBARv2Iqan0LCmyMQYjZpH
NfokbYGVhgMq4ncNP1C31scOeSXAdhFVL8PQBOeop6pn9HITWVC+Kvua8bCX
rNVsUPeLbOfyBqkoZKhgsyjlI8CitdcwsJO3DMuTYhp/FqD7gWE5tpSKuQWX
mt/T9FsPSFxZpmyBpM84Rm3PU8Vm2nr5z/Yx2IudI1fRoYQwW8ntAMe4p5T4
pk9Pc6xkoKXVLZoqQb0iZWzfVQmLEc/64zwPBqkOfbu3L9YTlygKlZpyKY4K
qMZWhP1uc2PEVHYqo9tAp0Z7BmH8/0j32dfxJUtCnToSBLPVjN3yBc7v5Hsm
uG0tglEv/BUS3aYK0NMGeCPy62Mx7/tkZCq8mEDTrkoT5wc7AjtxkiS+CG9h
WSaRmCaJZCwhTRBY4NYAiwv+y8O53TNpFWh0SU/0b+G7rWzZ9E8PV+fyjhMk
yl5YRU/RMiZkxk9bI6zPbHZ6xu/L1gCMjIZUoE76hOv556B3cyEVU4yCsiQJ
EDCm7sUp+NPNuWoJTqUTds7Dx/tS7YDyMcD3Us8UGxH4oJSIeHAxpvVxkVrb
r0Vq2g+6Ji0HZhZV244u+LOrVt+01dNyFyE9Ls2t6oDGP4DO+lTWQ6Bnj77P
PcsqpjoikhsvuCvh1bwyftZcDnNHZQhkD787/QcuX5ucwFksVHFoNnSoCAbJ
IRhxhic7LTHL0msogZp/HJ0qOpUSPT8lCIjgv/WBK56s2j9DskMTst/QqvKS
xp1NMeUaClBW/g97o9IJQ8JZEarZZW89oH31Vi13KMkhFVm0NEgPzpEnw1Dj
QPFoMRWsasTbADie/RpxMV9Yojo+WFeMU2AhdB3PQ+XXQIgymKdLwm49Z4Bl
K6+M8JlYo7MiHA8ZARIVQ730m3StPEdVoeGZtRRi1h1K3ov8uiLNqJNJHlR4
CXtD/jOwgnhrL0zfxSKAmYj2IrO5exgSh23CbgdYRujVX8NfCCryvPsI8GiW
AQX4Sb+vA/2LlcpNmkkLpWcTX5i0CfwOXZjKAALSpSqrj//qgOeTnUxoazOf
R8+oieyN3cs9GilfAcLQNh7Wb0umpsnAwKkKdANPXOJ9YpzVhTsANhVWTTL1
YbJfTsJFKPgmm+FLd2As0+bVR/FOlQE4hzIYkCzS8cjxVniuQvz2k5IBNJpl
PCBRTsbeNuu4waUiTXdv+jtR1EnXv66ut9rMpWr8m/9CDmGJlFtsts330fbw
y9lASE/RBDhyt5fgnw3QIG9wcudWnrFmnJVYNjLU/F139oYoyacFS3poKnWl
QjKk3Ubt0iWiNfoU9GdkKc+SklqlkXgaJ2rPOq/63CqhZIMdjZ0/u0iHLIL0
2vWw+6t4Zn7HUaGy0PPFCCslLk8+fZDHRT9o9hesCtAopxIveyEw5+11AFuf
rD2h2ZNRoAGXrDBnVnVXqonQAOYiaYajduy3urBhJDHNOpxn87Qp3mZnFnnQ
aWmeYx8A61GO4M/LYxnNlO/IndwnNC+6tCjwjU4gtXqxy3rsm0UXfslgC8du
MeolR7o6oiMBvQ2lU0Ale4ebXXDpjsQqaLLw6cmrrssTq6oA4ufNrGcz1yof
Et6x1QIL3XTep4OWcDYnDeCF+Xi1/toSb1wu5tgVtFZwPW1t/qkNmeMuuAgF
Gq3L1uNsbAQ1+xe899X9TbauWdjiwlxlTMRS6pWT+ecwJ5FqQO8pyKe5RIMj
OQICKFFIy5KcHpoqqo00rhDCDp8jw+2mK/hhbsyjvCfrvivNJs1eBIK/KLEz
88f+qO+hW1RmEfsFFM1lsvaS0SY2L/vpuLj/TWen4X6UzUSYQ8qeDcv3Vo4E
/GsxTq8/ylhl8lElKvIXWuw44+L5jLKjp2vUFQD2SjI7GAjgm5X3dHDKxipa
/POJFwN4iGulnFGaZkB0UsGM47QkS0VDLkxZ+9daevIKjPXG1w19XIMb/w1R
Gx6J8fza8B9gllhp+IbRsmykKFeCq6APeIBG/M1YNinDPIubO+9DduJ3kOlv
HxATc/AIErjp3ey8YR1lOVvsYfg2s+02lAqUGQJrfEjADRDiOaT7A6Eh0sW+
FDlx4C9R9tMSrBU7badj543EX2hnNG0yj477FtSEx1STOD3p1IMnPxxVIQEV
ejrkYE12ogN2TQm4PHXU/7YLqpSOr+As9JV7Kt1q7cPeU9WnSn8hgyq6Ocqz
5XXh8mC33uLH3z3rhOeL+jTqG43gGgLRi2PKktzdgO+Gv7k5xDw+uQPcGYDy
ERQYUOzAfRpcU60lUbJxU6MzQ3AlpxvNhCBrQTPzZYqX3k/K3hifCciYpnho
hyUtbAtKAeIS0TYu9XwCOMmj93e7kmY8sfbS9OvbAawgrlPS5NWqZQeeu7i+
/jMMbO6CM5kvOn9nFB6conlqqfWxh43jOy/QJNKlA3KtE3x7PL17nknLq/mC
ob3DzaOtpvRVO7lApu97OPRCH1PoK3EPGoHSSaddY5Ir21nlDhbgkPeP2o07
7XiN+eNNoxO4rlXSf5sxENCf6Uc//8yNfb+tEfeHOWTauUSA48erqVFBEPq7
AfsSWKRZlN0PveY5y1mW0g6Gy81Ibslmg186GZVsTO2pKhuaw3FKI1G+iObF
Z7uyObP7HQCysp8ZXJvcgfLAHIO6hRsTyVYJTXSZ1fnxALB4fKi4Ai0t1b5J
Mb5AIjd7csQ+2gVomjhaq7SiUodmhgEgS125pOnCP4en+T0NWEDwI/+XuMsb
PVSeQuNzPAEIpiP4jWwJlsg2cx7cZZcDGPGLggtCOx4rUNsjsz4NHj5sMQR7
f3iOPgAcmkSKoEksX/YwscToudT/aAjSq+D8BtBfrSzPnNgvCrVv665fAZK2
y2xX5iJj958uqRSVSiVPfTDM008Jls0SlryXSzX6LDe6zirkywVu+c1kqxt/
vrD1WHg6lrhnX9WutsNEz0Z9BYzmFhqbQAKCUnn6sl54TlvfzInm6yl0M4k6
qOfwHSx02F80I59Sh5MEHmz0ISiHbm6AnDhpf1CeW6EJtSkPw0swII8/2c0k
gz5PjScvnU+bpc9jkX7VbCtgnaDehb+qJHqE5/wqplGc9rUIsQUMeIGy/HHG
U5f13+ENvR/PA7p3UfpaBXbZ/cZKZI89tHrIX3jVCrTQ49BMHqk2Ev7p9XfH
feqO1kvZQBWrLQm21h92IkhiJ44CatguczVWM++NNJXBhv3viWi2WKsyezH1
Ujhv6Lzba/K4LkfoYoOKyFQU5Iy06BTUCUUuUS1z7H6JQysg999+OwUWaAZw
+gB/0Nigf/Evi3AJUyuN6yPfufqDjpCjNLJJhbcgOKeh7krKaSwZfptR4fZ/
s2F9iSOZlyYxg6C16KGebnSDn+LzOXKZ02e0/HBJQlfC1ePximj2GW+Aj0iL
mCo8lKEAAIp9mkGC2DbcSboUx2gqh0h7dyD8I+KlmG9iCfg1Ycq9qMnHeYF9
xafZlZFKA6nfD7Q2p75t5WRdk/ixMAEkrfdC/kqqbwfHh29evJchJZhYuh93
AeO7Mu6pNFrJvC6nm8xPJewyhc0hFifNsLyP1qOmas5wCe4Au0hTbC5zII4f
BcJg6Q+GSfE2auxBYdqbgC+5Ymp5U+mV8iUXS04Yb9DroGLNjmg2v2LnZGR+
JxDuLujxnMYs5Oi5sfRqmLtnD9dckC4MiUgHaenYWz9QzumP5doww2YmfcMm
swRJaCoZu0NUNLrMOP0BEsf995o1ZRQ5t4riRsdcpW7eTYcND6cXkTrP1jGt
TnMSpt4wUr9qeAAN7L7i/ofPKqAriy5b1G3Xsyqql8qTUl7J1eA22KvW0S6L
Ir0z6nQRDg2dGGXB/b1ZwfZiK05cJN0i5+9zOYC6SPAXRLFiJpZ+T5gBEfkx
0C/wZxU2Qm+JoGASluilbdz0okU7d2HrAYOy67EKvZeUYR4cJL2zPw/F2/8H
ROv4fWC0du+aY2ZDt3H6z4Su2FeWL8PwvmgcISnq0pEk9BlZhZJsxxb8Rsu0
n7MqIw1m9mYLL6E9Z6ZjuHvwmh6U1eA6sE83a09cL2Rz9SB8NM3BQcnpMFDP
ioeKYjN/nMVq0087uJXHV1yEBJlH4ilzmOyBp11LCEgt+/SLlVvG/ei0tduG
HnTHtZ0OumKJS/rakyD7S+VUJ1NmEXDkOuB5ylgEp2bKRdROCqN1WbxW7Qfa
OzWjhsGijrGddSc045eSi7ThxClcvLpFLvPv6Wmjg+0SMSsqU2V+iZiACnWw
Q4yI2SA9tF/IB1jhYFGTnqf1f4seWBxg1Wx44F4qSA8FtRhuB47h4YZ4xXiQ
B/HdwTDQIaZ1yq8DkryyAvnJi77EmsXEZl9lYF7/1i/HeB4eCgaGE1nPJwuP
R2/CGbgthRhA6sAtzhx52ZwuCj60CxoE0ixkT2r4YCL2InLJubST0Q47wE/i
g96XisMDmk/njUgkTLaZqiLG2iB9uF6oOhh/bq3MTPX0c20XxW/mfKguNJp0
GsUEA5UGFpGF8MAgS43gSc1V8NlxzD2ezm5ptMmTY3iYFaMuIId2hdy+1app
vl5nuSk+Naz0wcUWO26JlMYGdqeBm8BL85Yl87ubPu2kA/1u2+wZtCEJ/VPb
iTvckWhtO3jzb7QDgTfjBLrW/QMPFoMToA4d/cNlEVHChZGENV1B93aC8B1+
jM62nAoOdtWzsMI6W2/+YOnA/bgxESdeQq0d0VK1Fhuhj3vEeavR2oSQjdsi
tcHVHr5YY1JuDjkPB04Lm/IJ+4J0DjgMeX1WH9P67d57FUxoVzaF5ZjhZJ7x
4ynVxeu0BVdtwCaqA4mJAoWPtfE7nYUwuMSJgXScmiKKDcBQHQPvFI3rAPKp
qNPehRiN30YuFbAxDLYx72vWx8g+oNMoN2ddIYwLkG6SP5w1xCoROWgnD5wf
Vhrg8H8sD1i+COPcQnQ1MdxsmYRmEF4D7xuVmgiSz5xeqxUmeK4aL2yILMIT
DWhg3VCFPRN95WPeqk3ZX+4I0F3ohAUZYiV7zr3UoDFMoxRf5mUnOReBDRjt
3p+IGM0t2/70LqvX9RlPSKX7HK3aTPSq0KUONQpTZg48nSXlrEgnMhjS4YYl
uEJjTdTpvaSU16su0n2XhcufB7rTEAsX2TgNWkXICRrushLOrdjv26blzqME
E7Y6aMet9EQg+hkYwTpgH4s67XUuNucEBcxv9j56LI4irDCLpUnddWtStFJn
0A6HzisT+BBDBdXG4CscWkFqrTxN+zra6wI6grQJx3csRCjVOt6OK67kQJHt
+UjOIJLGWwxzEKEbJRZ5IdkPgClXvyRHHo6vr0eA3Vpb0rpL+bd6oLWLIi5j
TL+shanaTNQuY0b5X5eVBl2aVLUgjHKxynO85E2NyoMcDh8A3lBIVg2Nec1E
RibYiyM3AR5WDmsbZ8ip9DtgBkj7rXcB+u790RjWppSWy8TQuN488de9RA1m
d5z2LBbu2juJ/xhNS4bgwPiM8UirKHNmeGggWkPj3N66BL96BsM6miEXUGwz
X73L2EvD9KCDB2Uzusr+lPw6hs2bYy0HpdMTpgm8c9Pcq1prO43Q0rS+8qZ8
eOPTPNFd+DMkl6+i2uZ+Tq4exeZYwhqR1YeF2qAHLLNKFosaIo8iN675YW3C
uoSgBvnH3IlEgbq4ZReFwyCJwfnVBjL16oShmitwN++MqdlC37kJ5t6sa6dY
2HDbdRWHyx4YAc4/hQsgEy/lLOVhG9xqsIgVfpjIZLUDv7ra1h26D+dk73ss
8HpuSz1e7Roju3Ct+dvkpGk7fk0gMJRLlvx41A99Te69iJe7bU8UwbN3iYPz
Fy0sX0a0v+JiHHEPNyNuGLvy3IA7s4c2tlDZtlLnEBCVem9+tT6AzSyiE1bj
J9Nw5RDaC8tUkT8XDGCHfV92H785LkHq7WmsA6bLoB7tqXuDSrf2nDIqJFl1
SaR0bpLXHdfIQWKW31pUl3dXVjko+LkjERceVCsb+UDnkov1eoQmt2Yd/Nfv
KdMpqhcMlFmHwU+LL/DLkS7+WKKyVda947unQrEH+9lKOF+NZoM8RdEclAx+
3PeoboC8QcYC85ELGalU3Jucl4M2r1TXYb28zRCCBsACchtXY3TRJKz1/XJ9
QYqcY5o0ObvBMVD4wZAe5rjbrob8DARsqfgDEaW5qlWREzYZ8uf82axYKkt9
AhCWlWVO2iAlAuecDDiTN8rkxdi322zI5fKyJI+pR4XIt6h6yrvOOcf0BpLg
7Uxgl88yw1ZDqpUkxL9rE4C0nqhMpp/Q/Dqi5bEVtm5jE0R4F387GBDblFNP
wUPYoEXfFJZY6S6bI9Xlm1zeElDMewTu848kyVPpvX4X5tGe2Sp7EtBxZVmG
lsUcKtdQLBxr8/LRvcPlyvImSGlbc6qBTbyz7bjNvk0ZZa0tLLDScnyP58n/
VwNpXASDjornnzr7zSBNWizNULxv+DTWqUsWBnoH+DSbIwGEk+GrXWs+YBsJ
seTlwMmKkS+lbtNCT7wKOdxSPA8ieTH1FqWv07F4gIVVowBlAQ9hOkPNse40
N0hlYIa+U9GBS/5sJq2CsrUWmb9WDTVmWwvm73YMpXmkG+Pjnr9+ckZpumk6
SO5cd7SVkfrFeed1iTb88nehlmIIxhIUBhWnr8vaaaqJ/tVPEm2eSIN6Ol1w
h8ybpCg/P2fDedEk+7qUb/UTayKp7EoYAavkr744/cHlksado8pHpjNl9Oxp
4rxxjBl1Bqqt8m/YsOrJfI7Ju0bI9RW1szWbhV95aImqCi7/sf7N0CKb3rM8
omKyNmNstLpImj3f4Vx1zFJuLjOj9qM6CkGv+RsHiVXWMY25iCaU/U7VxgQR
DxHDIspLBfIuf33u6NAA3bwnvyUWw/0q927I8MkwMYqmcnHXRt6Hdcu2YEeQ
wQzI5kFritV5bSVEfG0DCQMC0s0hNrM3nup76g2p/65aE8P/aJS/HOaAZ74C
bBo3Mn4ujElPOdwfEKc+7c/kag0JziKJl0IAwK7AU0diqRKtlSTF2xh3Pav5
28rI3qnvqKS5f3eWK+BSLhjTePHJV5vqD2pVcGoJeGGgXIwQw/iZwhE8ANNS
NFNjhrKZdoEwKNNPA7wKQACDrVGdKKVWpkn+qo3A8HkaiIrCcgeRclLYeoCr
hw1NSDOb7wyXEHjXUVyegsUxXuSJo2DJwwUi7doL/aP0Y0b95esUpzVfntcu
V0C7FG7wpt+6IHX+PlbLSyNfhm6XrY3SQf7p8hWeQxn2GuBrk9mP9qOLeNaX
vXZWn+aMY4qNzoUnRa+wfaeUHPVw2rM+3zCJDVhzav0DHevgkr48JtI/fCvo
0ngw9Osg/4uIOCHnBw9Z198iBjykcNVoqmRBfaS7O9WLLdEhVro87K/S/TsJ
raciWVxr8eewCsPuYFjNzjzYM37hDzcbiLQ8vQ0iksooVzuQWWKAVQo/KLn8
t9E07StEPnztPrvjEPJiep+g5HszkAjYduBxFXsNddn9CYWk+zq8zvyDRITp
tuz1FrarhdMs/6YxFV9MqPDu1/8zCS1sYZ5SlsV+RQXNnX5Oe/7mT0343CKM
BIxNeNI2SnBYPg8KKS6PfB2Rk1x5oKy+ynTvoYLUY76FVKK3HHBNwaqx+qr6
6YA6/b4sMp+EwkbM9NoPWzHKEQh7M4iaC4QTXJxgaoXA9V9Wp/lLE/3kIT2e
laFzkGMuHDI533nQXiz1V9ynMbq1RNSoDEeSB2Z3/jq8tFq/WZ662LmERiY8
+db97oL7Dxx2YoO7oKT4DahM2DRMdDhqW3FGuX0X+wRjR4Q9LmkLqJ9Dd2k8
H6VuroFOcoY61ELaw9P5hwgpwTU9rf0J/WAD+wfakGbISWudAL1XaZkpHVUP
Gb4ym2XIoyFO+yOY+sGgOZ/xdfJQSQHknhwWri48PhLMC4AUiPXiGmrF9qhO
ZE5JT8bJVbMjw/Vm68tCmFPdmn+xAcpVWyoAYTvuaCtAaYinDFVCcm+NAPjW
t13DDvmYc0KNIfAJuDjCmJ/lKem20nu5tnOIHV8qlKuFFvCmlI3BNBUWLIhQ
t9JcKuGFx8rIdfpC8SHLXZ5yoANDTZGJJ/ZCzcgYBC1bAXHUq/g18BFZC/Xd
Zp5p0dhBZkwsd7T2Gtr6BQpxqGjCuoold7lnbZ4mwW/0LxLvSEcW6pa69Z3g
vRYUiE8xYVrnT8ppFSyZjGJ/zWgiDrgEf/Copl1i6b3zlSRGvWnkWejxzqom
+BCtY3X32YD/68q3dpipESRry1JbpmPbmxJK6JR8DnHSZwks70FnyHOKaIQP
3l+4MCsuJRkenWV1mtgO1xvLQ2IXuMLbQOJdG4R/MwZ0yGtFjgYQ01tzPJFj
205ypGyhvChdKYir6mJw2lpYDa29jYTHRSG3m5WOTxxRWRyXTjU/LQQCuess
2sssBbwhSYiWy34lpVH9TC2zeygDs5omrwKlQ4V71wxr49uzJaYkq1XYGEX+
gxCZqHrsNY2iUNJuoeEhOkrd8Nnib0unnODDOJbLklNGSmwY7ddkPZK4QCrR
tuKP50EfQh2mRuG/kKk/1rhVFApBHUwhkQhp+cmzSSRnWBo0qR6gskUuZqHA
598XLCMLnNKuxvInuf0ssLWALMwoZCfHn4rHKRDowZotMXBDmSJ5YCiolR50
CNNp3De5ghWEVKhS+0DZgY9wLz+R4UYJpJIhlKNDm8iFBV6zDgSfsHvIGxMZ
a30XjvuY2tQ9NQTmE6IY6WoVDiwtOGhzvFu3XE8EXJLRu7bb6UGyRDZm2RdU
Qrn1paGYuByDKLJ8xm5Wem5CRzlBCJj7bkdNp+I8Pk9j4TUFEfVbhqMGB65w
MDGf3mGjcNIHCksiQDHAVFqj5rWtkzv7GhLOBO8ixAaqcE1cILg/5e1LZ4Wb
w27tjNLwWiiZvHIriY8+TvSXzpcm2Zq/PLu714n35eW/sFlLmM76DEFmcIYj
VMa3Os8dqmSKf2tegoxxwqK3OuV/IA3/Obu3ogXnYhXwJa1p6n/8QRDOlOEL
OyBC7+vnVIsJ18cQgI+1WfvZ3+s2bi+20EsctqKOlSa6Z37s4CLSBPAs96vj
fgpCjo79pM2howKpReSs+nCwEQIpJqW+CRSuBqb01usGJpBL8KulcpkhiObV
g2lSIj+1+k3db+xB4NuuyL2xaC63jfRBZRKAzoxweBSQz57SUiPtc0ktL7DS
CjZ5/23pdOiR7ggzJexhQySyX7xRU5uRLdigSW0covipdaTPHhWlU6ijG66j
SJ/xkGA1jj4vI9Xt4KZsvfVu04ylQleUvuZf6uJHnW7mxkYdbSFLuxSuKaXv
up9NOupQc9DahaUS8OWEEKUIb8hPS0rgO6MOsqskdcYNXDXkwNMgEl3zaOrH
uZYk4SPuVMClaobJSdma+fmk51t33UQAr1BdXtuTUGUJLJFH8LxJBib86qmN
FrYv+t5qh0XcDscW+VqMUm2eVuiUos9jcNsxkjrw3X7JwO67xeDHpKDt+p04
QiaA7rsZ8VhxFudvAzEPeD+Sej3oqbwga2xqB6DvDbdjy3ug2IZ/PQbmWkEz
nQAkWs8nflcCdu5f+Cotaq/o0+g3M9J7iUF2kDMgPOw+4GIirT8b1aFAj2De
bXZKeyUSOjDJRLXTsA/b9dmjzAydRIbDckm7XDx2Dg90AcgsV0Hfb5KaPXBf
YvKgUwvkDwmFlY9+ipLe7UcjZ7JsMMN+didicU6dBns946YLW64beJT0uqVB
rdFVQDYh1RxuPRaYIvT3uVHSTvd8xCI7jXGp6XbGR1hKgU6SHrygJT9NfMs6
+SOBO556xoUUpr1Up83OLe4dnHvAk/58kLHTpBJ6bkg6W+lzLgi4VNkyE+UO
0MxxiBPTr3UrVD3TMHi3G2jbjpshKDxwVQrOzgdMVMC1RL98xEMUXIekGABQ
NyPWZ31FvtNJTdviTq5ewWt+xssY/sO31J+aSoSfDNo6kOWCxPPSiCGhFbzk
zARaTt9TD2o6MKI/hkprnH7NA+6zNOb0h1wbgO+kQPbnQPScnL60Hdv7lfje
sCcbYrIrJ5A3cLkzyX2Z9E6hEF4XxFlhyvGExn8+jG7UU8mMAoGcbGJl9FrT
vVbJpXYtYTlpHGDCNx1/CnhvR+wd8VMzMhPelqCIK+pbyDNNcS7keGLT67b9
uw9N0qt8rwdf3Ld4HTPPDzerXkiyohjPWS9AWJXxRze3mz++lP2pDPZfKHNs
7/dsIHKixwpJaBLbvvtBkum7Xw30vjOGaf1/Msa3pMvHMlAgSJV90duzJuLA
Tjs/mpF3bYyy7wDFwddbVUF7PutDo8trUscBXDKIMZK+mk8rHKhrO6r4NdcX
IamlZXBuQe5dkrGEn80xilj6Yimaph9mb2kovedEWpWl5CUvI/nd9k9Wg+eZ
xND3JpHQdq9Ra7diV04v1utsyrO6jL2iiJBzBhHQZymiO+ZIImiJn5aIaASg
csHFDNfzDzzv/ILdsNSIMfyMYQRY2y8efK532SC3DY1dwplx61EITIKWIZx6
eOAD9ZswfYHniT22CZYNm7JH/0mqxYR2sNQHKOqTKAnIxDxIuUhLZj0Sv/n3
kETi5rbpBXc7rcg3i+alLSnClTtwwIhRi0izjNN4PBQBwLThaBvp9A5OaaII
0nS0QvJTkToC6p24ufV0ghO8L5QkL0N9KRkoKVZYhqBGY5tqtKZP2sLKeraH
WasstJObQ4vlbaKHmWrgZstK+eJvJxPOT+riIJl+wpcXXearvcEJMswbhXA4
GDGNg21gSs3HR2f12YfCYmFc77rzsoNtWbNF6LyI6Fltsu3YqlFX6+ANbSXW
gmueW3Jmpxpl2Jb6LianjUbzcP4pwqA8LZvMMJR9ZYypO88/fFH2JVjQJyi3
k0ZTpENACj8uzBUpEoRaex/gRH7GePKq1yulsKdRYLx2V6cqX7L5NHb/psSn
xeuyOZammXkfHUt812U0LqrgTTR4heZCdWcaO1TmHNvUAjAKauBFbJxqE54J
G3xqkRJXsF/y3oNSCuNYQG61Fk0L5FTVqn/InzicuAC8pMfhknVVAaa0TFVe
CWokbkSQRECOAh2RB8peH+D9ELk1FVT9mWYucEiHD/daf6LvISUlDiX149Ve
YG08MjJyLcPFa/X5uJlUSqtICn42ULEAitiHBAxI5zsGduoYOzjVhwYa7vnt
yt/N6KCt/Y9XBl1jLqcu2HSSHaUVdGqiyRuLLwJ2VMXuDtpdOuXN6j89XM6L
2EhFeLpQK/INfTbpGk12vWhM6VjbSzmwcGAzTiGHoAauE6YadK7YdVOm0E2r
ICis8dRK3If34emli3RzdrM4hPG6oO7SQsCYRYg+Td9PZAbbp8lNJ83EScRr
Iwkz6K+JoQIFORNUwx9uiG7uGk+oxVSXPV/RaYNXCtA2VbwTEuJUUExcx5Vg
rlGe7iiQUwCokU3xm+P84Llupcju9vuwrfJQTv8h0z+mPxpzYERovZHOaSq3
RZTuVf60acd/oPwIAqXAFYHrL4AaQYznCiETjOEpbEO5DlXQwQednHeKHY/C
5I7zoSvPZv6MACMt7gRh1jPZpIeQQs2pWwOZT8c+dnyWfIWawLrQ2lZDt6OM
aL3ZwdL3P50ylTr25JtSbIpqBP2gSB0FlYKYuhzPsWTFWXvN6ad4JaZKrC2/
cB2n0ka5O1lvw+Xb+JjYvAZWsx4aQwTPj6ccE7itP8VfbQXXxnU40n9slmvY
u0w6S+erCx9+K8aPyemyY0rCwRCvv9PsYf8DOVn7X22wqqieq2YfUoledxme
O75r5nJwizoIMolZW4KEzXQ30D9q1R+aFvRcyvc6iYpYpNMonNTUUOcguHc0
bi7aRfzI/lt+iLO2/2DcpskICLhDgW4DZ4cx5h1Z5kYKjvm+Z4Rfkg6FPj7z
86itb+4WyOzJnSZ/WfA/83BiND4RtIot03tvT4x1JiOkmFa5pP7Mm2JDXfOL
P7s4oCIJyzA+KLhx1snZsuHqBdebGZfDDBERbtrmLzwWeMrfCAqysDSuRjc4
Kxanvxs9YjkEDMXJDquRGQBD6qEZMzn+GrCdZlaT5qYx0eI3/Io28WDtRuZU
ejFTDhvc+lq3Z3lJgU0ceBG6rp3SLuSFLCS2M1Qi53ww81+qyvZh1umH2xm8
aHyHnTpF4ijwJsgFenZ1yvJVr71outkJTRpfus3tO5kctNH/tVUBp71OQz1c
TnAUgk6cylWZ+kjinvqZiip0PbVGkVzab0Jj1uiJtzJK8U7bAqMNQpbncGtQ
551X3rAtYpqYc8p4C7k3/+/u2g7rJPwqyvYfXqLdE1G+Jfqvv/zlGiubqZi6
PB83gmu5oERvMGjLMs+ClYymIvXC4qIr8UupdSheWbrqsjZ0gnrX3Rwsxjnf
t6mJNqTO4YCSgPx+e1Lh7lV1pogPazguC7r2Tt2mwh7TdKWJi8mPkaqKz8BY
uLd6KYOSyxIBufxY39LfvWIzx4EztiK95oQqQTMSpNrHccQV9TeZN+vRM52u
0xrfJA+tknfBGYZQCVjMUi7GPlrYS6TI/RDsgZDrf+5o3A1t/BY7nL71JP5J
r5NhIdG//uhGen8pBZddCbNdkn2O1lO3D9yGbUZu0ZPlIVxjsWRExGcsEDUI
lBVrpwSwdx7RkN1GgbQkJIl1IGkBtY4FBevezZNSbiLOk/6g2IIB1Um6EODY
JcA6M90UpagASsO6nLZHGPRdrzAtMhFboKWKxbn6L/PUbLr/zy3JBNTQlzL5
o7f8CnaWq9LoUE+yNTSoGnt3umS7sFkDWteJFAYq0VwV+LIYavNsj1vWEW3T
+cfgKK+WjvfMVdXyzATXLT7UU75z9+2oZNzicDop3zxTWzfKAvT7xPzytsaP
6JU+bVYTyP60smj+XR/BNFKveiG3c4vvD43SDtBC7gUuQ91tgtpnJmG7u9nA
Elxvf1COSHeIPGghEhNcAEvUD9b6u8u4QHnYGYsboI0S4u+/R94/4qK2xFKV
2wOGcQXl8RBmox8ef1orJwp4SxND6msQJfumKelRPiJoAop/M1GLPuC6Qnck
Sw5iDbCgze5Ub5xmL7zcBuNxCoT8t+RCVPHi9aQxys9WvgaPv/ktzDWR5UeR
mLWVqJ9CLdwbi/18cIjKHE1ZUYROJwSSgRkkTEgKeSg7dRliZ3mxNkq6PLu2
BREYsHZhQ8O9XTVN7ZHiYiqwrMfHTLp92iolfWe0DEPDOMTYYyw6S/aKh3KJ
hOaTbdcuo/DJz9q34kKRXgQlJ4k7MBVf9bFgPRzSt1hgltUitvQoxXRtBdjt
NzgfJ0Yy35FhLiGAumq6Ya243jlEWC3B3kfeCp6XkT88MnXAbeRfaMTYwvTy
NKPzKfmcpJ+EAR6O0jwYRTacdXNJJZ0XlCDaFayO9eprevueA4xlV46L1Mip
z/Ti/Yyk1KahoqwbM0rGHQM6Z3dlxxAadtUSmERVTE1xSCiHdgHF2PfY0zV/
/89Q0lJV8JWNVV3A4AZED2deV2S0yT535LlvkdfaekO7aYReY1eCYk/w5D1p
1v4LH73u2XRxgqLdnSRmQ6DfXcagYHs6DDPdNlxluOvQgj9B5/9wJyO3gSak
d+E6SD5fOSRcfDGQeOdqKrJQPq1NNfl8GSBoo/f4th/X5gzdS8+1YIe+ppoe
p3zWLZvn8zOowP1AjcOvfUEn1XasNTLOjp8O4oqSh2w1dPm1awCttjBC9WBF
sZEhdTWeWBfHqsrNyDE2tZZtn/2qjUCO1/7t/JDB1P4ZlFG+QrHSSSO2Lecg
Yd6+FJl0Q2V+6x+CR5xPKnv2ml9ELIMSMajERkgF/8cSV+JiqD0x/AJKhajd
bIuPHcJ2w+BZOfE7sJbSz2yZXgLJJnzCEFkR8uVi/WoLmzOSaRgMxHL8W/fU
KvGUf/XSn/sJOgRbB1RthX+m3cag9yuzmzTMIOakKFEqGzOyjZuXvEf7jv/o
RbXtFtNnvJbR64Zq8tHZdgQHOgGSHAXrYIXLFx3TQ5PqXQBrVHDILTqVcBOP
WzHGXRW6YLR7OUjPADVLuMuULqOGi1bGKVwqsPNaOoxSfX4DiQAuBkFK4nSs
c7FODa3A4gKSPRIMeGVNIp71Yi3M9OQtK7ExOm9GdbjZ/X+3rXp+7xDCok8x
K0B+YpVXXrJaAQ3KjGNdNugNJeZGMowkatdsaDfXClqMfdT/HMqStn2zDyjv
MN/kBbjXF2ZNZPg6emosRZQftIZtNrUn29TdXWFWMKzxuSMcJWfgNTA2WsFd
4sTIRO5CQj+RJnocoFnwUrAJo1KKzqZ0T7Mt7B0G4bIyZRXGAP2yz7nxgmzX
wZx9XJZ6tGEYEyJG7odHTURNHPc6HJmFItZhaLVa5TrP2dk5NfFgOFkeMcRD
V7FHi5ZP3ldfQDdE5Ur5bFzHWA2tymx37sfoM2bMMUBFVoqodanrfqziNA7s
E9QKQ9XitljyVnUIa/MgGbi7DTC+MKsrAuy8beMJLEiMDFheZLArRoUHBmcI
f5A/BWMPPsFK3z9KVpSFtriJM6q4iFGgDDYKhCZgobrywxGq0sfcJi4hHrv2
Yj85l/1bvFh6RRyV3Wks6AI5XHv1Q8IksaoAtdRPumKPQ51zsMVWq8L6nYBp
FZWjVHyu9btSqj5rFNntmZb7RRlvQrRrYM8RQLDy7gIh4qOW5724JGzU3ZIB
jtRePZHGnw//Rt0onKsaCCygJ85v+l/Mg3SXNFriEM5DgW2VnFlTNtUJQgZ0
CDF7iRRGwa75SCKvh8ufnXatT3zpRw0B3HHuByGb+dcR1N2M/63V512OmV/9
O1fkBjtUnZP4z9pnf/8tMgT9AyH80CNWctWzxc3g7NmxzxVKuenFXw6B+yuP
uWlV6NYU0VmeT86ZHmjkvgjYDnkjIO2ts9wltPUgr5RQZXVwJ7olXw6Bzd9X
RnTHukrFTAPZTmdGCJL4XnAFw0OR1XZv6eaIHc1lzHpH2BBEHP433iCTDOI/
8SmsMFy5NqisBqj3w6nvzkZ6Fsl6GD8HXlgcWTLpy60amtnZEy17Le4pR61+
/bYCVJaCRnZ+WejnHZf1LxFkoTtWRjkz/Y/50gsarnei1y2YafuSn80iXuhw
qQl/KbAJH0r36LSasRuTtpqLbHsY56vKGCycrUOl1mHL1xi2r1GOdYfOYN+t
KukeCujDXWKrR69GiIpIjAu0Dl3ATrjhC9/7cpJFVn8ZhO+Q/3ZQQe5Etaqx
QVc+icvJpMWDDPg/EOE0XS23qB/KTP2wimApuyBf4j5WStqD8cjc/ebDONxt
GUvGQoVGQmxP0a//ajgNUAbLl/9Ark0r17s2jt7QM+pplLWaqyMY91ueZNj+
q7+TV9j2+GYmIxsO5+PuQIdcb/dX120B4+5kObrd2LnVtlm1lSH7/KvtFBho
uppLMN1ou8b5+xC6TKipMXhl2J9Ymtn9+Etk1u80VOxhOO2ncIHIVQDocw3Y
HqHGg3/KENehlGhRH9ChBqcmxTrsxKmi8PMxg4JUHpe/Viviap+iLBeIa/to
PX5DyyFYckNCyh33Gr7D4x9lT+w5ML9fhs5qKZDxXv80chg9fQ4mUI/gAtmV
yuCJqZiixG/sfuHY+8ZkEG1bP16+PNLnHRhVnma0zSQnsUaohGWgqlh3YxlY
uOBe+1N+omybbX0nqIJETAM76oQxuKsyCDZcEPQlopncQLFcf73l/LI5lzol
6KAKtCt7SOol6vs58ENM/7pcNMquaAR58H+QshDqBJG3pCF5+oeEniC0C6HE
HxPVIHLWPXObbHfCoFQ2svWemYpYhrSJ0EmbZ3VTgDrFZ1HZI2v++VA990bZ
aU7OnKv1o5Mwb4V0cfDlE3PxK2HLL7qukk225fRaCIibcD7yCptZe1ijZDRQ
7TI/QvDKLXJc7eY6oGA071wGd6lDtguNddNYiNqyExTga1jaNtYf3NF4ZBr3
DpAxDIdg+J8Mevlkmkj9cDVes0iYMs35ilpdAeWqfRZKbOGee/nu6bAxr4Ch
RhOkKrvtcfpAme+cSWhXI6O1WL1O85rJFCTpjhSyB+HQbLILUspzsitMqs4e
THYocFkwWHxYz+axZ5dNCuGDsRaDkzaWA5w+PAl/sBedgFeudhkGdUXU8vFX
WFfeFndFnMMjWGdUXC3Gn2RojmR9W8biB+4LS36DDRwI8sRoklz8qssZK1WV
sNKb6HV0agy2mXXmrd4I/jzPVI+6acXu1JdKJUaF9IaTNYLTt6P8+HZXhJEZ
cfJv8hl/Z3mU3Cwg25T2nyGTPlzOtmAeWqZqSeOWTMBKLKPdRIWDS5U54UjL
XJMbhIkvBCl4liaEuHDJEtYxZouzwSod1k1dh5gdma15GEWE/8KTxmg5auKM
N7pIPFEwMZB0O0gl69rUv6ybtjJyq+9DWLvtU4Ah1RH/mFmnqNgiuyFY+2/i
VcOoe6MUUem3KRKQn/pGFNBN2p1LtldYR65Iqe15h9RwGRz+YabhI99Gdn4q
jD2O4NwUAoPtMUUamQ2blpnmkU0giP0SxB3yHfesoLvYRw6Bjn+tam3ERE3p
8v8OjGNE1UvVPpODaJCO7X+gCxLzwBVR96/gnIPoTi7U55FC7BJwtvErTugP
629Id+Yz/BNHqMlnTemniXuE1ocxfKCrwgP8ezh2WqJKZeCUWesyMOJM8fTW
StNoTHaXmECW1k4oCE8tZKDmslOvgXSOWaw6dxDfHgksC5z5jVZ0Y9MT+UQy
ouns1nbSedvXcmdoQqnsUgHFkbWXT++uzesvtXTDVqAG98ohD7MtBswHxSNn
kTaZSoOYv5bIQo9sxgncXn6yWd4WDNunE4at5IsQ/eloY0wDn0UKrp8zPuI7
CLsdBjPjP7k2+IcLHJL/0u1FW8gBZMu39kx685hfWswsj1S7U0FKJ+ugFEgO
oqqGdnt3I0yXTsPjXIPN4Q/NzbOPRagC9Oam210RC8nHU5MudIke88qOBIUz
MCSBmH/Nf78/qT+yrr/E+PzaiKelvsUw/KcvnvgpvF4C/nqyoX6J0RxViUGx
h+ofqOf3y9pmvjyj9z/wbo9YpOpqA+bCxrGumA5O6tyaX6jDmmo7vfifAtBX
PEqKSSy5HRzn4kToWHTIPxG00nniU0OcRFvj1F1q/oNDIiX5ONj1JtovQbLx
p5C4l6JPN5xGzJVkLqNxayS2PWXJ+6uJAsrubhk/3xzU3NE3voKGkxvf6+Iz
OOr5SPwu2ODV5DUe+mfwlkkIFP0naX7Ch/bp3GxuwSoyPBh7QIQ1QJ32xdNO
oT7pgWxs3QI9rL+Rn0ttA+9sA0lbgCRi2fA3PRPY7+P5FPo8bja89/KCkMUk
fj4WD1SF7aJ+rcss07mKsfmnHGFb0Ekwn0iyn5XynimKVrnfwglwplpPR6WA
zzhCx/JC4oSqtlw3summhTw5xJLa4agYSsSx5hiewwlS107A+YvqmV9Lbwe7
IFVStkdsiQQmL6TbWkLZfqD2JrfXbRAHvWNR/aXFkBp09mFNvUlW4cjW7atH
cybw9Pd791sLXRi06k+LZ5BqSJTNS56Hx70WZDLMxMNNPT5oHUL2hjIsaWlQ
tQ+KAUN5q9FTU/m0n7gaUJQDw3xQ2yKfWKrVjaTvEBMJawWuzhboOZaUBwdf
xwbeglKgyXkQOO2sqnz5iGa2i99ij7GNSLZa+oPW0vhlJvUliSkNq0+8UKo3
GDFSoLVn2Jdqyuyv6cw2CrvgWkWkP1TSAeiJHf3T63UxQPIQNYEJYaGTwCaP
3xN2JVj7jyfXCgJzx9UYkZ1UNNE7ZX5vEc7EfwIBDNQmHSkeEwRwVLRJ5WAJ
42weQk0pjVGsZj6Sqh7nSeBKMPsZ5ofTy3CTRsOj9hNCPsl1ZAr9zVaX7ZOn
WTQe9rKF9i0tZ/Yl9sypmU7ScjH0HqHaVFk5Ip23evHm+3nc2iVD5QSxZ/84
YTJW7v8zJliIXydvCjysEiQY1h24+4f70eemq3siGuExjVb8gvt46dyaSMMV
lLRYOUzWcOFWf17OsUk7OLEy2t+oJuD8lZfTlAdLWG/Jhagqt8fEgwlUcJiq
1V/adFxT2fEmS4A8LxL7Us1+x+c8eqfkbZajIKe5yLllMs+TMjt07zASKi2/
SZclAjtXVctnW4NMHxI5oeJ9UXfSsYNeqnaNZLgdZgXtJXJrN5rKukaARMZE
N8fF6fX83X85yDohHIvvmXwwi8TZdTzX5rrT9glRhl/lalSWs46+cdvP2dHc
JcKO22DMwwEKTefgt2gZCAEz5HY+ZjiYMask6OCRYws0ouoW7M/2mTxj2SkQ
zb4DEnIycdiMKw4OnsNzbiCUMIaupoqi+TqsuwsCCOhSI5d0Q1zouT36deyq
y/CmfLIt9nsFhro/gqHvk2+biPp1XoSzucSI8ocXShLzgZUopp5R8rP0AjXV
BmRz8ZS/jtwks8oK8YJ5QH1fY1aXCHblpZ995vMl1RolPfHAEd1HM98PzHqs
WU2pppnXgyqNkLsplXkxqZ7HuUJH/vg59YTBqw8HICMWEn0Xf23mlOk8NRpe
+DkPJ/9CeF3DdBt1yGDNBi8WXP0aqfvhr5nTgG6sKvHHc7IJI8ReF6JxCvvL
m/aXuSqOjpCh1AAcfxNYSbURbpRj9VcT6ZDKw5X466kBKbaZb5tCRReokasp
NRDdMsAj8R6ZcxDzFFbFgMJKttMP92VetH3CWpxhA73MTIfvqIKA6UjW8x9L
doJEu0r0+hz42qDx17Ltk7igoaH5T00cfFks8CMAj+8UGACSat4M1lfM1HYQ
nckXmc0+V6Fdeo9wTrac+uU36d/hlMpBulKHdqXbX2du2bU3bRzUwlY48BrP
ii53XatZSd5PSZ2G3a9kbIaEN8drb5g74MPYhmg1zNtwtR5KBOq1yx055R77
uXIPzlKn64OFRQCVDSwU9w5/YuN1PJq0x4JqbqlGy3x5zFOZapWYQHm6BYYE
GiupzJbYcO3HSw2Js6bRY2n6eTIxvuNeV6xU6RNztsjM4CLNS3pa6YIm3e5t
QQKArng0FGP9jWvwmz/wxsG83A+XFuwAxXSh9fg3mY1hBKMWDSwkc14TXNFv
T7TySdoiY4239/G8ZrFhx6NWI+XwVuV839w1UbMWTpqP/FBxReipdRbAe4lu
LtuR3UjuV97U4ZUHZj034d5FUEpPvVJj+c1QiMn9SNg/IzKbPEtVOMmOH12T
SKzilJuXa84YLpF2d+DO6mrSMbJw4fG6YMKl+L3IIhSULezTgc92eZi3SUIa
Iva1sxLF0kk4ez51piVNGuQwUSZfWSj6Pgw4YRmT8xr04bBJcScJ8FpW3tt5
XtY7kYAEafWAnjWBzAmX/xd3DK3BqPG12c8GsAbGNkYHmRwcRnOuNdqrTKQX
9WFmg77+bH7SIbkUFlaZTfE0fQx9ZHh0feb8CKOTYVYDKbdCV3MWKq3OABET
1Clqdimc4YXITRy/t03eDHFXwwm+u/5YzPQYPEGBbXD7ElJQrcXmnnpRYjKO
cZBxkbc+uaJbavNm1vCUA9aReAZqK6Lu0vlYGcW/uDKh237t2vq5vqB+mU5g
osLZgVUATnlpDMZG7gVj4Jf/n0a6ZkI+mvRYIiFsmvDayrtOZ/I+U/+WSv6O
7yTh8UUvIcfCasJr3ksTXJK8Bmau2tIlMd/pBpY69LwEwY41WpAFx4BlgNYj
vFKN188P+aIuRGAqilbAYxGmw2p3WRYkc128Al7T1MQCzguKKVBCaHbsgu6j
g5AtXdG5tb88kQbuBFkKYaAqEDULOeJk1K2LdojR8edKHr69a5Ck+rDEMSah
0G/HGVvK/b80X3ePar68eCcu9T+pJjx5wwhYp0NIHYsH6ji69iteJLMvOnhT
qx2BwAkWIjV7T+aUbSN0a3YzkbcH/xNhCrdMc4exCuOUYjLKP5SIJ5A1Oq2e
hj+80833NtgxmNpFS8gJskTNxDAQTroPPMYf7ug1WMLJzwQEU5San8DH7b0j
Hgs7xx8+jXipaDVn4YLrQCDYr3myE7qPgcOhnaIgulKXUFLTSvXAKyasIOgZ
8u3SgE4eaQeCHI/OF67VRt9erYePblwB0BjQIMfT6kOc7TH+7sXX5B0yJWci
IH1fqOPO3YBrKLmj3weFG2/yXSkbXRfI6OeAEY8oy7Iw5wQCyU9SSLIAxgDL
9Lywp/bDHiXNHo4alr/5iqTZpo8R1qDx03R6ls69BrXzE1V1Fdzku2wItR8D
dD5srjKc4a2qbka7DvEIWdDB6+k49N1bmT8wKmowM6FDvHEftrBKOPU8LNGO
KszTM/JUwRKi+WMm9hUGcQ0eKSTQKEafPQVZnRkoYPUPzD1XGgtY38ObBQDS
LhXzrJ/bQzk4h2o9H2Z8QEXllRWYCtHwy4X7jII6OS4x79231sBKtGBmJNH1
caV79YXIYXUVGNws+/BYGc3uzhmJ5eaoetM0yq0TWVuI0gFSyIKQEjYQ6PGg
lXYi+NvdIfwSTRqf+W0GU62UqYgTS+KzexnBmbaTX7w4R+9T+a2YWonHRadq
KD6YRgymimF2mkJVjWFptkBgW6YZhTA+muT/NB/cvWtg0kUBNwZynSapBoJc
Oqk9i4Kxh/Za3hxK0GloAvpDRBKLg5qpF+GUv+8tAjqGxL7ztTeb4CAzac41
JhFVylpu0OYuo+fSpTGS4y+7kWeuvRr4sdamtBysBX1RIKOusqyDSjJAlbHB
3iCKbCS8KddCb09Ew5zBcUV+oSgviAgMLfcviLRs1xxXC4GDMDu0mIP1ZCb3
2xDlCVRSkiK4OnE3Nnztzj3z2AfB/6PAVGGRAn0/eEj58nvB5slUDXzu1+0o
1V5WXme5SwlwCf38Rc/YnbJHaIqGb5TEa8t7FViYqhfT43fhT2MOvko/0ipU
lvsRuQVl1dt1Vuk5lSBQHDWOt1pSWCCsotcygcaalKL0OgxIb7gNFr9+cCLV
MIVJ6NMWNnKzZ/kEIWZg9QubdiDE6v+u+i6FKcSsNo3zh3KXnLOKVQYmRsfl
XPrZAlw14oNJ0Jc6GotHnGRoAO1LtLFyttljprlHI4mhd8cRQ+QpDlZJ3ZMT
Aww/jC2R4SQ7vBD6m9ZYn6kL8gGQjgHACJhXxjUq14g2DTWyiuAn6u2GBegC
Pop0U7ySfEGbOqtHXa/6gbsh+8F2HCwl7QMdMbCWCHTy++quU3JttsFFfXnQ
BXEB0rcvl9hISaWw7nTelG+OkImptinBOj+NOELhuN1E0Nr00NwWnaRLv2jV
PrZeaMnhsfV5zlM3eCtxHPsVMNZ8wd2excRiBb4X+LsxpuOtLcwXWVhwPji7
QTiRtMmKz1Q5XGCbI4gydUKmh9oMO5P3AneVdnNVdsFynoUgM4yK73be+9b9
H+e6kXniVw7jbC+HYNu9gfQ1FLpEMchEbk9rqXWShbUCe6hSGRdnGFaKX3G1
HBrFBaOPnLN0KKlNdtYPI/UC6vU+HEqSAxJtFBubvfTtiFiyyDjdBYZxlTIl
5k9hDeTLRYBbAq00DOI529bFKjyU3RoRbW9DlRX1MrbmtdiBhZnGj7pbydfP
pGH9FRlxqH5MI6/hpqBIoYZ9WRfVd+Ti5SOW9tTult8aVfGh1y6Fyv2HMSNv
XK5G4M3IXTZyvVJuSGCpMTH5dVud2bNf64LE7c9W3lgyeolHlyT/mrK1Bdv0
uall/QW//RdwH8PgJ/JzFxMqmV3GdrKwfElX9WpXj4uvImL4Q4BDdacZN1ki
nBlVZhuoZOsWiq2cullPwzRyDzRUPEXmIaep3y15RGWsTwpoLuVj+9wEPDZe
qMED4ZpJNR6eZp+8crnJVtDbVBrAsyVHMbSVtuosPKPX4GNaQmVrfW2EECKI
ICCNY3sKt28cLyGfgDMQB8jm1NF6ME1YjIBR9cBuiYMPrZ9gOfCBeGq2IPlp
Qcsg74MKJlefNbtMdnaw3qMD9nyN9kexRcmGBV0nRmTIjfEHXbrizbsI85f+
NuzAxWC+oHk1dr0htvOCyeoXjutP73vEI5WEge8zF8GHZYtqF0e7Z/SBOPJF
J06iTUEAc+bL1rd+j+rZUMwFn1Qq7B+z7zAQWbVClu5ZZDOxcU1PE209hpWD
32m/ddKcXa4ifbyLhl2VKbCdOx0/uOYKU/k6cxK2AipEBQLoBpOJbol9FbOE
x/56sH5qXo1ap+h2zfG5f2bblRYYG1Dq9X7ktdfa70KsZAs0yf8nA8GDYABZ
HuTmmuW+3Z37PP+jY7jSuDmzS2zuVuMNg4RWS9c6z4k2EoSTxfqdY95Yrn2g
u6+FRH2HWnNFslif1O0f3Akb8uP36b22ivzqwGt4cGeqnMwhIfRBC6wKfXAl
fdcIM/KJef+6r0BHiw9TsBqPdQnhEoHgVwMZz6OILCfDySHFQt9RU2URA2su
6jINcTdKUisaPmMaTrZlt9yFkj8/N4VzNqD49cBcFMYph+iEi6jByTKuukht
f34RT1awi2DxPSFmY4CxjV6p+puYCBEDX8QC30ZVrjv3jWCRcImcijsXgXQX
BLkYloKtCOV5yc/QIs6pQyCj0ChBGC3lzXDiHZdJ1HPny/kO5Ka/P19FZV7A
h4ksQ+U2loDXRAqXVKJq/MY3GKpE9V9ShW9gBwDgRiUGiqhEMv38UX0uXC0j
/CXyPNVTF58+IRKu3TgizFwxmjGt/8slw/uY7ADm1enFZI415xKZs6mgW3X2
hGRYbEjV8KxxUAlZplLgS/6QU/JVendsqEMQn7YbM1lMEYbE4MvRDMXlhUun
ooFaEes96bki9078SeLCrJ2xjV8qZnQHhkwT8S0fpT2tTyElvPRPI0nXo0uT
StMnZXLe1hPy3ohEdXh8P5GVxJp7eIsSLNNFNCt/HVTPI7EaxFbxvWIUpS3y
7wyeSFNApgiIabRw6zKc8yB+nrT/nXc61a1VQtL2JooPcaTrKLxwwvi/TAIZ
6cNhZa9Yp0Q5LV+sLwIEsPc/4u4Qqsldl6ne37Z2YaDyq9p5Vc7PB8BCdawU
6dOuDuBjZ0vO4JBihQ7lEaa73KJIHBPjphMyv+EukeIcCD60KxNNwUx3fwW3
jpyQ/egG2n8m2APH3KMGjyH3KJBsMxBdzDq8gGtPniQLFjrF8EpGrRHKZ83P
aABSxTRPW+HNqD5OVV7BIF0s516z5VD1nIF4OR43FbiL2AIzMpszR9bcfWym
qtu5uig8sLN3IBhJ+lr+jOsgR0Byb4o+yLS+QCqlL5NRwiLY7b/kxK7lipV/
xCrjDEBB2j8rA1Ix+W8wuPSU+kIccefR51UiTc3YjZNWna7xcBiro9x9aJ3S
HnDPirKRcCjFaplWB6AEUi0DHlHRxQ1Gz7BwRK3sC1iQ0F6g7Wq1tDqV0XO7
Lyw+099FDxV0tqPoO/wkacD/pTZF+Zn6HphvVkMnX/VCq7+qdN5AQom9DKvd
gVW89TAIwclsHEuv5umdK+sT/peFBj98TClVU++oANL836JFv3cGE8ErFtLL
4KFbFykjcQC/mEx8d3QmJEhlZk/+p9VDjLQZU4vd4fGHnqXq/qJiactmYId7
WlEe4THhtGqH1JI6vnJNtl6HO6D0S+2MA5jlAsxei8xLwOZ3ZZxs2+HtoRnn
BUcKoWAO9gG/43eNWWU4rjYxlKN2XvVW+ATAFsgVrgMTA+ckKeRymtttUHgK
iipKFlu8iniMDxNuW1wG1y32pndnRdvefn5ibRIb1T/AaD9/KtQa0PVheyM7
01Yx9ZVUT0cFo8M50IGIC1dkMLMupzfH+rS/cmA/MNYMCXG3E08YbW4OT4le
c68mvmiKA+Se39fetg5kxlzFTfHyCaAupu/4mBTeJrKS04HI02dZBakiIYoG
iMLsgYE2vGpNyDyLoZd4Uta4g1LfLrfau2DGwmzNg6F4s2QxYICAtIo+R8Wx
dhm3TVwbsaboEa7IKYsdlcwXWRhWrM8seY9nEBE4zE4gKWbS94mwTe5WVFxu
f9pIo7nQJ8s+3l4v9NdZTAY+/bMbxBDO2TwiwUsgxDym0jdFS8BjfHqR6Mhw
KaN9h/56hMo9Knb0pyUhkKov0N6PwmyGH0L5x123K3R++jJPlcktGDGmRjix
haURDErcUygM4QmzXrNqYu+pD/MSr969+EPMOx01BgLOIT+f/zlBozutJE5z
ipsVvLYMlzrmjaSWNfYCfN2XV0/G6JbLcpKM9JpyUFYbQte0DLlsC3lrDDdN
UvTFYUokwkXM6+xU+m+w8CeHtSiAIEb68Zz4b44HBZHoTEqu0pDPy7NtJeJa
ZDVGRaZYAnZAWjq8oQocxW6lycT0CD3s3xr+jW04egSWA09ojxmD+hxXszDH
V0GpwJU5ap/AxKiUL5MpzZonQ6kPZDuloGdzDJR17WNHBwCM3tJwOl13VWPw
zT7l0GVFvC7D/VXPHkN1ubRUcj232OzceIvsxFREuL0hKkhaaGTsgtmAna9e
dFUfTLq8Sj56qQtXaYesdV0pMTF04xw7ZoITGYmefTae4At4VtNAV9G0e7R2
VIl9R81oI7mAvIaoyAF1j8XiCkUiVHxkstC1IHYIBI5EBjzXN+kBmrYhdU+w
ANMvUf73OZAdtYSOz6fQcesR1J1xmospnH5jn0HevYImCT7OaL5smzohKrlI
T6yXaE3gq0n1IZprdRGsTYw7qATTvuCpxk2QXXN1tyJcoUkEKmxDiQHYGxrQ
8ZzODl2vpx+XXE51jcxGitMsBl8WEGAS7sG/pFgprfBRQiAAKe2y3NFXS9wg
QWq+2bHs0MYlJz9ox8favsnNc9r35NjStHM8uA04e6Lhv+vLuwbG9N4Zb54T
QL+a8CLclZrpJ55kEnrckY4Gq6jdHZ18D1gtP8YEo5/bMYLaTDPmz1TTkQjc
W9MlalpUD/KsILkcT6+jc0TXl1ZcCF5AXNH5if+3vfZFQz+4sDiv5ElJ14QQ
2jphxndGO772t7QveOt04St0exrvAISuDkkNVeq/lE/ukKisxpdL6eXYzT7g
+bW0cr9dd47sQdPBmrjK4fDC3UY0CyQwmgUZDmr3g7Emfn+xj8OPvellmkr6
gPpZewmsTvPVYyLs82YERV/3ZGi9llK7V1wtQlXPbPztHt9CbYVSm4czLw7M
SpcuqReoXKrzYUWSA0yeQ6yGVY4bq45f2E2hLe8z1HyjkfGlOUVV9JrnIXLd
pW6d2c1cCzdoimO45b4kQJXRC/FmBCG+maruA84PxHd5sV092GP5Kn7QlhUY
CXUZjg3HkF7yPi2Rx6uTZAOguKt7wdOkEdAv5bVdpHIoE/wdfzn/Pwtb8dl2
YBDqaVoa6wHMgrent2l+ISbzRPNBvWOlli7q15NU0tz5Alg0NRCkSK3f+XNJ
y17TNFs9YkHVnr8+kW4yInmimmKn6tgICfuiNK5wVWEyzVoUjBhgRmkgUiy6
sdPgJ8FKeCzCdo5ygzETWj5aGjdDwUSlo1wokJEG1F6DPYA0B0rdBY4vqU4G
FhFfhtRu+nyG8P0wcOuUuHp4yJcCCyxyhg+RX+jG2KzN8nIemAjuGMqcYbIK
xhX+K+B+LIbNXoGQvzDDIh1Ex0EOjweUrJW2gr+5RmPQYNHw5mmEsjWNxUo5
nYgfJVcVRNIqUS3bP6Ifc39mTXTHfTCzFztNRuBK5AR+FRFsdNiVubUr5pTq
dsB9LuGNeYlg72AawsXkGflAOO4SUZsWl02YHsq4D2/El51C+mQLJCiE7pWa
pzDwNG1EZ8mSUj4MWtAm+N2etavTAB8YeHXLy213nF5Ky2rPGqkcXPFwuc3I
QwF+/VNG2mJYTZeL0Vch7cw8vwBA+NbW2z10ca/UZleb2hQhyQZAnZmImXRR
vJThQAPngcKIxd/OGkf0+2dFffV6cd3FrNPCS5W4A2TDPTqwi9HhVkHypewE
y5+zMRPNrvcNGrkPKWalHCiB5TUr/PCzA1ZIgHfIhONuZYpysBC9XyzUfAxC
y7DLZvytY+RVZTmHqEwdxw2/hbBYdw+odM+ozmY9pyR4moaZCOUHdh0XHM8R
KoDKSupNpz3jcbAvVzGulKxRu9D37DV1V/+EUMX/yG4dlr8XHv4QDdMJCN3q
qmdHX90LeCwZWo9J9+1TdYkI5R7x+RhWzVnejvFzS9BHhIWN33SGbYXrdXa0
aKZMrcyGy27h0vsswO1dobKUqADPilPvYFJduLqJHo5Bl/zRwbeFHaccAczy
EmES3aupElqFU+rx/Y9bsqSrxyN4K779+jl7uW4SdZ+O9L8W5bkuyOpRaYQM
QwewQAEP4YBINi/sfwiFaf4HZmBu0Le42r7Kc+ZDi83pWZsIT4z7Mvp00UGO
7wPX/ZOSRNBK+a2HA0FYrW7EB+B3dX5avVnI/YnUeQWASIfv/lTMrpEwIcxr
sYj95HPLoKfoSirW26u12SfIvolOhd07L5jXBXZ73epbznwO/O3sMCVqFuVz
QtOBenupL2rSxnC7atnDmwTg1rlzu1/uDxz6y6UJvft/1Iwp2OzbxN1OPDaX
9SItrXHVsAbgVxt9qRRsFFSKJyYjZeaPDzTOQmO+r3KJ7Rf67RwSnc9ZAc6a
k4PxNKbDQfxXVYXqRMGrQf5KmIAwGPPVCDf2HTwUt/A0jX3izUDToQEhMNQK
uJLHSt1G+1/XxgQYPDDl2P6R99icBoIhcJHspCcwXitU+e5FgQ8c0Sj4f/cJ
3JjbkyqltB47lGXK0zKwRmEJz2l74NEYoKJO7/jrC9RZb0yip3zNELw4VuLD
MLTaujZJKQnyfp8/NdKfAF3DnHe9bI+RFIGHg2hVdq9xzzlektFRDK2CzRK0
5Q17qU13TvXGroyGd/bjYacts1Pa3H2zYXdAEwaOSH9rqZl0beopF1fHgSq1
CHrdBkCUmH4Nv3ppP4H7ENMPlbnXm40nNdgxrrDijj7ec/CXsDgwRsprfsm2
LExa/7Ctn7UYFeWBzylDs+6URKJXvGaJLakcJiNW/scOjstM52njZd6L3z0f
PDi4+Pg5T9XYpE03JcopKjoX4fsTxxuce42ALpROHHfgms8pk/F2JywemWr+
Iho9RB0eXFY9LXbI0dHbXlHqEi6LLPmkccdIOrqz2uDOKncA+LhAlJSAea7R
8d+DBm8lLoM58VKgLgohmR9f9UsyObu2pBW7eqXJf5YtlQkc1n+sw28fI033
AnYCuGi734Z/Qz7hhIKGIuKVDQMOJOR+JzQr/0vkhehoU4Mnkzf3wxESK6dd
h7Wp69UvpNK8lrexlRnp3fFi2TiTOV24Kfg4SWFAgzO9/xYA6NyqBydhWO3s
XEbNWYAWxBdzXpcSatqOK8PGHlHcMwyrOc41k2L/F7NaH9TKAMJ8HxfP78vu
Oo1EmLTPUH5meg0DAn+fSacwA6DjCy6wJSk3ftPUGsmnov1xEs3LUsMkh862
G3LNC5Su3vrlAm0he0ezpvHi133UGp2K0bDTcmCU9mfLfi0vqeOnZHY4pKmV
ahNAhO04QzUFnmp5TtGJAP+nCVh4PLFBhv+SpWKmyLYaDcfBbS/vSEOEx6uZ
cLCkhbX+II2gdB3FjwtafFWq8+xTrpefAJfAh5EweVeGaLyOQnkuR5r8rSzH
OkteBpzqStRn3oj0N2YwW/oczH1C3ZJaHfsGknvHpab+PGkODjtrKMeMSsKb
98PNO4cefGo/V8gl1MkAHczeXD1JWKfF0FSwNaB45O0Y7HIabwB7NxooAX2l
HW0+tIRyUuXmPycuekCEIQU7FB4DBLURxKdRoRqHLZrGy+hoN3PA1Qgtx6wj
UNIpUnfOxKcv6BsIayx5KCJwA513/vilyibrQi3zz76STdLrRDPdV9H6osEx
vSRAR67YGsptbLCvdg4+o79MDlPNvrbD3tnSlpSvJs7qiqWmm77RP5zu1kwr
MNHYL2RphfpYkvA2Jy6B6uG8VJCZJcKhhUSBTQWKwK33uXUgxyKSZkzpTkFa
dws62C4xBtgxSUJL+Q95pXwX3xMc9SNDKah2JzFn7bF6eYwHmL8R8h5bo7vJ
3MHpTEj2YwyKoYwPbqMc3x7cn+4LPgJ0giUjXJpjSHB+NV9wZtgFJ5bNwviM
EKuwMVL6L35SkgO6R9aigyYxdBFxpIfEE2007OZ8mRsNBVr+lTPNK+HsFPaF
GtvN6zNqdn0cSrnMWMa/Vkh48Fe7AltvFjBSywHIrQTkaf7fp5IPpBxj5b7Y
F+P2Y2QIkBscXhOrlvZUouX6Tkrn3F9xVcJ7yvhaUyoT/UkpAAVUPCWeiPZO
atiUXUilM5pF1fJ2xKBBWH5n0Xeu+G/pV9trqFkgoITQMFDzJUrYmrcviY0y
lNbSQOy4dwOjCfVfofFFsX5USDbBybzDG3P6cXSdxaCGrrOpGQb68QjQHzSz
mThRdYJvfmdHuGRqK5crfugYZZ4PYuuxmjQH6bXer1tPKzftAPfibDvRuCII
VcD1IbsEbSfjCBzbH+ZHEO8+y/Xuy3m8yUP4t0eW2e78wbHY4hgKbVk9Ygr+
SIFtgUPFbpZHOIAMr0GTGkULYSLFF5FPxEhVHLK+lfXnH//hQUABXhLHkme8
5N2Q0unWZQIqaQ82JbrpwdApEDPOZXMkDZPkDWYsrJ+1sDIUzhPdEvX4kSCj
QyZNj+mGToXUSluV1/3g39uvU7jQd1TR27qX6GBMu/Mq8Dxv6h/jv15wPkO3
jBius6MrHGRioB5hjU6NxuLAqBdOM3PCRwG2oi97xcjs0GegqTkUd/rNouwe
to+KNvXf91LFhjEL/n0/LrxG3mtCdaE+toQYwaGFNRkNNvUp97NmV24sqy0r
acxy4Wqh0e+npP+Y17/sqoVloJxHAI5pCiJNMa9+y2SNjYRspxCGCUgnQgRf
A8xYRIZDBudIkg6fJ/uxd7rYJdmdhgGhensrKZCvdgAuj+Ad3jtK2bzcQqxs
qzEFxgOdRkyj8fNVwboCSYQ7YnF0jPXJlwBkHwOHtgSox8nZNLm6v0Gb2Sv2
Qb5V094kIQ3ryLdWAITBjLwaVTlCREi4JuxMjj3vTprRgoztk7EmXmeZoD0l
7sTR9q77NDjEEud29Gm0PakjLST9IZcObchJrtmlAgoPS0qBju3e0e5/DcMi
gGljm25WkNBQ/b6E0hse1ZM4NyOwXu84F9uMrrXPCrI2QFXAKuY52LuYscpW
3qJXSoRZLlpbLPSUJZEUn9vT/EFsWiiGsnwWwlVFJ/WArstwxGnO/b7C4CQn
udPHqRupkDPkeekC11jI3zhtr3WmQOzOF/NhxEq9RgusObRVD5qOwyc4lCVU
eyi1Gg0ZgisDVFY73ce2p0laeBPT0RwvglTdwAFchIpv4nR8wzCdPqVZiJu5
dkniYW2sO7FDuxZSGFYVhJxS2mlTqUFgJuHRDVjvV1x4k80ypFOW1MK/2IT3
M0GcagrBuUd1hsZcwhxDdaqPQBDqiB+ftICQ8cmRN8CdcXErlmL2Oja3S9bF
UwIZ7ee8miG1fOsns+w48uK6sX64yuE16f61Gy/jAa5xUPRA3Wcq+xwdcrtf
s+cV5bTjLW6Fu1gETEwuem94MeeCRIQOkpg4j8UbEVfew9EKuhbmyJFR72Co
cb9UZdOj+/dqwpwXF62uxI5yZHCYzKANWhQPsOZy3ujEJuI9ZIWiu7obMy2T
ix+xh8A88kwE5jXAjQ85Fe/5YeTZRRrflzuIbds/XelkUshgNWOglJ6tWek+
Rwn1hXVT1JVj5x0brdx+8DmntMbmJSlz/ypHLdRwdo22wyh0AoWGmZqREI/+
uTmiKXjIeWO80KIxY+69zmrULhMbhtugP7lVu+kpX7Gxg9JPhitYX93i0ITe
8CNFIbDhV2HrFdmJapEIMBr09EiNQUKhHWq6mvsPLxPGyW1dtZtc0jlFyUyt
J6vK7khydBrLo49stugpHMbDohf2M1wbCqL61+vbtYe7YMdYVk/dU3aSxOoM
4iE8CP9QGMSCBvRGhGSrlQqY67NEWn9/YpprkDSwvceFtqMpUI6VYzon6FeR
fntzNPfqIP1BlOFqk6ZqF+ghK3slrSP2Bv2dPyJJ0WAIPBMpuCGlZvB0pwF6
bPf5aJFf5KLAUXUm1WmGZuSnFW7U7Se49lL+e6Z7QRqPePMqgWnhOrlTBjw1
hGpGRoMN0HbQt9/dFS5+dE1iREvbmStxHqxC6RtizCutkhd/9l86ipZe9l1g
V3CgVsALr/eiC+fQKAEZ1zJA0cTXSHJnKEXlV1/pbCbZxNMr328S8+YvqwJU
jhHM6h0LAOX4Un1YWJtbrA7x0rw4t2GgvLRfemNuDNIA5jeZfGsCr4kHfJ0p
4049BGM7h8FMu2wooq3PHhHgc6z76aSENPgbCBXTrGURdWQPgI59u5wD3DWs
ng7xCxKs6k1E2cxtfJ8aRhNGniHmbbnSWU7JBBVgJ5PJqR51iO7oeIhKPBYl
Qv835ijBU9pcFORPxC6L9pxHfxGvrtHUExhaA2phB1ym99RF7z6vTbMHLCvB
1BnoF1qu9YnIXUMj6OdFQb02kHLQjvyTNjUJla4LMg5dGDZ0p6y+750Od8Jx
cyRsdUuy76LH2eVfoy49TCkiGEV9Jfj0c8Grzw2+j3B47SEOcKGb5sPxZcW5
sW9FIu0TzhalNEOdESeZR7spo3+XbDdq9cF10I5zcGE5GWA0iYlDvUbNC/c0
7gIgpq+EHMQ4gfHvDdOX9t0Je0bapTds3GHvc1FVVcVgOdWI3p/PWs8dDb+U
3qpVqyOp2KS5GFAx3MbrG70bLUjAYpYuOIeQivQ1Rc/cCQv87JXyLrxz/EM/
/zCw8saxNTUZjiZby9yH2lmlAGdoYKX8+RsE1+c1kjaTh01s81zNcgMX6eqb
mG5SU7PGVBf0FrfgQnhlIU1Lcg+cZYhswiFUpTnKeUA/LdzOL4rHRG9acZho
hWFHwQ2qxsvMM4cH0J7Ol4owa1cJuprxNIS3SN15qyg9fBgFHHwa1uYUBieB
tvYW7fbssu0SmZj8CFd2BaVLd6r63wz1ixprj2+fsHXTc+4TIaRrAuFB34ej
0mNkMGsaLwxjBgC0YOsMgvpGKDWmf4GvZzeNeKcF8x/ZhvYHg7fJ/WOLcBzr
5wHY1ceLzrX044GWmixf9Pm5wkVGNNWDXqk4c2uucjfCs8p9ItHKdiqqKBYM
imMe0jv3vavWjW7a5GFyxeki9sfgiCXbwY46VV2PMdlp4UZbmUzsoAzseciJ
GThFTQLn7nCiYaijjQ/s/Ac1Ckw3qiEQmA69fSDt7hVNdgsQ6dTOfNQ/onWI
6m4ACqNKXu+QkXTkVSje3RPrr/ZDPcXU6LhWIuFTY5bpj2QQiAOD4Npua5EB
QaaZs9Fe2yGA2CBhuEuMJTPj54ds5SZiFEH5I5dI307jr9cW0ROMt9/TrJTA
K669j+O/3Qw347Jkfle8JQj/b3KOxKAkjviSdEVky8RJa+8z6eEPEv44Tbmf
EWkmqghT1EOsw6RIWQcg4uPKfPThIF9foNMVKsyBmFiblekD1Nh92GKj6w39
Z2H/rSPYdUpV8Io+oV/8SdRZ1QUJ+c/rrUaOx+Rv/TviN8PjqU6vkIM2e1Iw
rRhNfz/MuPJFQ7qPrIWQ5E0Pfbc6m6vKVyrkM4vAAZXcpMvF6dGQ1zvNv5hY
aed2noa3FGGYoEPjFlxEFQ2BOzB8seadB6AhYes9cgSshvJOfKbR72HIZ/Pd
X9X0HakmYDqabXLNgcKI/GGQ3m3ofVvjnwvWOoSaNi+0XN2OlqhjLha7AO4n
1su9Hkiy8zPoYwQQ0yY46m42lD/jyOEIJFYxN3n0+GXCcxyj9Nj+fNOC2INE
68dkwJLVgE3B0Kf5DXCYyK6rxqcrflmRM9PC/Ur29KQb9n06kLbE6POXkiUR
0EzfGIQ5cjV6T7N/e15hKYMqB7viB5mbAO2U8vK7HOqgwx/OoS9GDbXK7eYZ
WObkAqEdln4FuSLYSSLuEV/ha1ZmFd9u/xpPgQpgfnCgIknyKySBf0ZNo34o
LJn6SRVETT7c4dRujaVrL+2KuAVr1ZaGjnCNJhudw/7P/ByVczuj0TuR2ifb
lMNUfJVFLuRCjhXbpSBZ+OFo3OGkHib6+HuNDi5ppPmlcKjoZyPv/kAzbdQk
KwMjNxIeMXh1QQeZcPV/jcYLmV8SOnzUsmEpn+te418zB4du0dwHRfDgfv4k
5btqyiG402CqswyoeOiU5rAlEmF7D+X0/yJi/9aIh2+1vMiUQFf1cGTxbQ57
++Zx7im8KknbB8YuDuxcYmPJCsER/GchBofX0hKoQJ3xkVaCKTHmPxnlAikI
fI0tb137zKaNB5b34av/Qz/0ohohMzZajLVRvjELyBeXAiBNAYmXVuGpf5hw
Kzbd18RdIvIem6MGdEfSGbeYcIzAjDDd6bBWmuI423g4ccbHb3ZEhJ29oOmB
J8Wa/01M7e1FBEpVlLOh72cpnkLMIKr8DsQGQ6O4QsSjwCwWvN3bBnKijYAc
4GfkavKuiI5JB9QC13ws28qpHsPmSypsPtdHELUVfeX5Z93NUugyuHrf+Mhv
oWv5I3w8jnX2jK6CIRzr+H4bFWVqJrFRjV74/S4rCCELG5Vi7wvNRnN/pgmV
EKTNrrNqrH6PcM6ObEOsWaVlIiAIJg53CfkYeTK3l4xGmLFS4anTiAbdlHjf
HObBck5jL3RFviq06+CoAj/5IhseLkYM/EG6PUYScPfR6LBXzT/1hEOQZkA+
d0n1rOtv4tryPQDBZBXwN/rzbLhqEG235WzHjR+SIO1YN99ikiP6/xD6zYAM
oJpQNYAYJ/e5dBppAxVATAkAaqI9pWVbTusIgruC9+QWkBPIckpMM/VwwbjS
anvqwSUNjil3nESwIKtFzOmMtcRJJn7dYyJ2QoqYRAhYGZ23sBXMS3WKLfH7
lzT0bmsMLNDW5lqUKTkMawxf+xkzAMjItF9jocNCVW0uM5Z6YRBhINaJdg5t
XS0l/Gm/Xyzv/ykBJmgQ/3Yc54sK0/zcZw5OFfWKpbrmCb6WVmP0H+ZRBPb5
+c+OLiTe5yrZ0VmD6kjIsBOHbAOvyQVs4StHHcKEtya+Mv3xD5n2ZvEoN1eU
+eWdMP+Jyo7btBCo3o5CS7Sy42lhNC5zcW9fXQc8KzcvgVINZcBbRjpMscPC
bzR6uJ5fX550fz468WtdMfoLEXfec5xWn8hRGZEQsWcfAnuO2KVxSd0516Zm
hWRqhNWpxkwq8QMkj+qX6h7q4KNfrM/xyNeN0NqsLBRIe9FhEDkkE/brfUaW
upZ825IkPvL4LY7rdh8uDUwwS/eptfLQ+SOBYYr4HF0mPtZumF/tag4yDv8T
lN5nffQomvUkT/pKs4nEMBSquD5XI+GwBiGCPEM3RByj9VFaLEq3ZPPK4MvT
bvjHcQKgNGsIsJuK0L47zeYwXygXS4p2N6reUuI8See/zuNu0MVRQvMKs16S
eZN+KcEX+UQ3FqaXJmJMbTzq9017Idvj1Qul4z1a43IRQN0XFpdIa9P57dS5
PgEGYoow+ZfQD9W0DXJryVTE7miJG7cxUGPFFJ06y7euWDHcTD7PgfFxwnjF
uYBYVGDuhYrS0DCAQEVW94Gpq/h3Prjrke01497qJhuqGX41g0Kz/4zYZSHv
WaqZk9yZP9Z5vSttM4M88yFMpyEKegMR5RK28Zm/Zq7JjMGBy64jXQtSfurw
7/j796YHGgaxSP9SBSfViaFbsGYEHTT1kCRg/3HZPf9wS9S4zXLZZ4NloemY
o7K5UXA4jMzS/W13dQwc+IY5ic6sa2vqsCxS4HWYRMuLFRQ4uNoi+HZm1I8y
d2kTlUkyRxNgbp6N80j6kGE7nC7YyofTM0mgcvKDEUIiyMjw7e8kX6/X298m
DGSBj3oEt64F4xNyJXEg5jtCIBVFwaqT+4LjRMoU4QmqYXS/lAE9xxJXOc5q
ddhmJJ2x8Azp/a2gWT4e5JL387Cx2up6Qy0OFPfrPPgxsgw9y10dlOxzBqrF
r1NNNW4P43MnZja8v/p7U+etr6b1yqQNaoMkiD8nALIduXkMwrSFa8g9TqII
3Bs2CefrCHvNjIgjhoD+pPWlG0RG00F1Wddd6bsdD+R9D6qxMVgQoMCJApZx
7628kIhg9Db2KLOL3KQg5L0Uytzq4iGtS/th+PRcrDpm6SeHEU4pGCECYbIt
C+5miUwyogU2s40QzJT9WUHzAS7x/Y+EEsmHanueXm/RfPSLyJJmdZULav9F
0r89arl2E0B+MVoulu0irqnmNp3kOX3L3rPACCMhwts8XLvjPdr0lQu//K29
rmm3hxpIbDVCZ+ZFK7X7OWJC1r2zBUye5r4nuvbvFpwUHa2jr59T8zqAFiX3
QYPaUNxqc/VPl8dXnFY9zDA/aPrz/VDwN5VMpfZrSTC3V4ebJJWYDLAnoDjo
DnfYnywYu8YfXOKgzDCQzpcBuZDTbVGWE9AhljRm8Q++SCRxOKE6Ysxt+h9G
cpaaEc79VBCsy7HWadA4OlHNF+fVewp6SNI5gz5L3K2iDofUWb5IU8XBrtCK
Dlw/FLu5HfDFLkGJEQgbnnJncaxp+MD3WismOg6qROBOvaevgMtvwVc+umtU
8rnE8CK2DqCL0IqIgLjW59Jgq9uZU/fPum2MyBHDCWUhd1SD4DcgUElPbi78
YL+EbRjPd51DKJByJhWZEjsmhRsfO4l1JF0h8u5hwqjmAPClwFetIIEoE34x
rW16wwqeUR+pr9A0mPJH65X1zjybrks1fQi1I4HXh2EGJmvVQfy5aOrA2kwA
M+KMZTqnAi7H8W57urJEWdAq6U6isDkAYJ9ka3ivguR2KlpX6qmZDqY5+QBw
7UFfJYY1rjgwl6HZV4xaHGw4W4fy+c6kVx3kAMw+RNRQbDOPyjKEHYwltWy0
X6+h5ZuFjGv7+rfKyvRQbH5kzFLZUcOOOB64lFfLrARo3IvCln0KFL4bjcmm
4a6NoqqadZC2T0xuz1PFPlg14WJzBm05/5Jk+Z6oyp4lzY1VEso7sjcxJ7BW
vpNU6A4nsPzJhLBZTdAZEQKpzfGzyZZVXMggPngrWRUHBrFNnpoYqOekWrLj
Q5b8rxRd+M9dxfKFvaKh4SX2gwaO+E65x/qQcc3vYJlgy/10f1ziKlM8aF/I
BqTWGYWA7H1ceT1Flm+L2XgVHKtUUYu4FMNDLluoAkemzYNhYa+o0z3AdhXW
8w/iEBYt5KntGiKZyvBKHsE1zlmqw17TY6q3tsWGgNmEi2aYt7jRxmF8Somz
3KPD8YRzboojLG4msCWEQTPkZcDLg4yf8bO2nUsNjx8Gn3U9m9JotieRuQTS
A0Qgbg71p3Pw+VQENa/drkR2BTO5SviVG0EMDLnIs9frHTO51NKtl3wZCiU7
mBcMdUY0JZiz+nCu3SfzbJwhVWsDLmo7+R3zjFaCiP2jU31WXKs8WkUrZFy8
WphfEAQi3ZXe+IgNdJ6PfFk95IEr9N6dIGxxhiW7GxjkfwfbxeRsmAuPwH0U
4AWA5ZhmOQ8QSSmgaCY8p/ptOn9qS4TbTBVhJnjDllB1DZ27QPatNqogr7U9
JIbMArxa8TGGwQDmyk49tO7BHD2Tr2nY6ZunvopFHjr69h6PKQxPSncjwZVf
JlZ3ypXoRAJxfN6pBnmJcVJ+1r8LmgUT5p+8GiN9lGv/gajnI4pelbuv91qs
Bnxff82y2g3yBw9kWrYwX2x2uzP6nrGCN8d3EzzF7t3AvrjDCPIqFeM5Y3nd
JB7qPqGgLUF0fdnhfbESSbBUCgCkmLuOLPaDrI8aA2QXGt4wFUkl9hip6OhA
kGKzy2+rneizi5pkhDTPkq6BGRaTHf01E3MenSjosSaIT4lLQyC5K6ibaBcD
jFWx+uzwB5vMOnd0vyNuZfeKrEZ3WvspxyZ+Stn0eQyzWu+K/DsDAhCoXi7h
wOwVOee6K1hY+xEE22lQgmPGklFoU4XicdIFkhVQJzR/7oW0W3/3O3vZvBod
lNKWqq8jMjx5c8npKRysUUYlX9KZfyZPzxMlVpjh3ZDRDJxKIG94kzsecrgA
CnUXET27L00/DT/IRHG7EedV97Mv3x4HXD7Td1j/H/sRnub5Bi2/O1ZOm73n
UCQ2d21S87fvwO5hao7meUXZt0cUsf/PY5pV7ft1d3ZcTFPBi+ggK60mKzs6
AuxRg6ovRX+LG0svgEF63FaH1HhVS+m7qyIxpXNytgjZfyLJLzZcFUKlBzh/
83hI9tkMhuuVXACS+VoVVbP5PgpqAVAGxfz1tII61XX9wPCDFqKmTzI5QW5R
x7SdCM1EucXZ/gkmpJx8wbVZGhv499Lw9+u/Hsq/7FBLeueqs/xtLt2nHdVy
H1ByFFMzUYOdmhgxBE/GpUaedu0LNlEF8ZKqIQe4tKpHP0Le4z2Rntpn2LWr
uwX784D5xolwF0yybyWTNKFjvk0wCuoC2rzhIGXWnb+bwTbdjf4hO0WKWZlg
EE+SltPkeMjHXWqWrrniTrAkvD8JniJj2Q/DcGPa+x3zORkrwCw84+L3n3vG
J3mGwScBggqnFrUs1cPu18IQRMNchdDrNqlGN0aYj8MxoWgq59JrNH3OpSnC
QhuJoicvYC0y+12oB57GjZpQimPafhL1ApHpmHMSV6QufaPjGSIUHZBLgflY
6efp5caoLIN89fCUGPFXUbk9FemSuxaN6BoITF1h7qojb3vtViHwcuVENHFP
fqnB/KIlN4il68tl7+Y+AMjyTQ2psEyC26mxuU1mMHVX2qKC822FU+nCd2yp
Z4yzQn+pBSXvIppTBJKPtv/kPb09u4SVJrkijhHabHyeB1t2OAzSvxHKWCK6
ZKQXAdCou6pkrS8XmgMKO6RsfVGTHTJhJvpQyQ5dGTjIehAUHLeFlhx79exs
Udhoo7py8n9tmIY2x8DVQYDDbGvQ+hJRj+i3Ibz09VN1MtTPP8Vn0deDMxG1
h780IDxBROphIEW/xLI58Ztd7ooaWneuLkwc3JfU3VMtWM+i27BtVD4ciGhA
KcBZkBio55zNQbEf6K45TzNO9nqptvnua+23NIQ7ALXvUTdC0VU09qvBtkSF
PCPAUd9DeT59wCUTUDUDtXzy2NAAkhBOAYw2+YNs6a9dqA6sPtldMHjLuDJS
a3lE+qdUZaP2+oc6PtRn5pYpqk5xgOdtHh1f6aLW9xtnop+3nQnOqLnE7ExM
hM8Z52z5gPVe6XojVgNMy9Y99ogrg3cWCZ6a2ZByuQNfsnyr2G5Ok36yeLGb
uVrIWFc/wNPvM1xssY0x7ccTnci07ldK7yBSqETHk/9S2Vk9d+CJjYBsXhNs
zcsIG0YIwSoeXLI03f0DC1xT7RNLX8Enrk9dv65mLk1SkTyksbanPwEDeXF5
Fr6+WEYXa6IMLNOQQhTNE6hj6OnQsgChNsUruwKh4NMEeAFKDJzBwHs2PPrS
uHmxAn1LOXtr7OsqrVQa0uwo6bIVMgP3o8DU6pDBsucCweWfkRUkvhfWqb47
RK70rtina2mZvPnkdVqmIoLcvAES3h2C6em01x+FgQqFwkDg1E8BytUiPHNi
LtQ+m38K7zYegAIrNXrXbLMg4oAjNJKlik0zb6laICfyJHfuY0Igbhm36xDT
0jNX9DaW6Kl1SuLiV46NCNBnb2L9/Ho3o/0pdu4FjWHy6Z7MlPuC+8if2dr4
1qczEB34F5uuKawEoITHR0euc0CzNTPDv1x8qysNPXUqw+uwpayd1o7WZ0ZQ
gRbR+dshLMJW+QYFYyABcbm147h7ZnaNK6Pftqw8f0Kmz9R77zLF1ifJO0yU
PDhmjS/5uFNqK6sR/efgMXXzQZQwixAudEf5+kk7vff8ZqqXSWKwCMB2ayEV
3K2FO34oi3Bc1v1vDsbAjspPFBVsyaBGIetsjKuo067FnAm0ZzKhMoH5loQj
6wTQELHdhHkfI2sHciNKI8yilfS9RabC8zouImxtnSuyMFkwjKrgtIiJKAM8
0ye+250R3Y02AUsj+XTAMQz0Xq+UoYm1FbFBIaECaUTqYRertoLzAK447lsQ
7mPuoKpaDeEdsSAEgrGq1uJsPeWgBg9pLAINgcjGbRKMIjDe7cSL4go2l33F
G1UHX8vvcGAli/cZmJeMygNW9bqvJ6uNysp2eayf7DrxjHS6VXoLD+Et7POv
tsHUDa1duBoEOCLZc0xI9fwa2xd1aw0scO7cJvB8cPvquXKEQocDAlUAS98D
7GZXEHioopf9bQSTjc0bGMGIS88LvTE71RqI2hZxxxdFD/lXkZIrnxn3PyTj
9DrrcTZIiA0yfYSMDm8GDZ7n4cSL4ST9GfEMi8yRgPCsw688blq/ndnj7ECU
cPXXjYsSxkukfN4limEs/YuHf8fSthwQd4Xra36QGf5JxNm1TjVvwByBgkMJ
4olhFCRTMAx9mjXbc4pr6oDHMFFgDRO7PlvZYqd1C7rDbTrVYiy5NWx96mRt
jm2wvK52vtLWE8+IEfZyr5YOBlE4VFxs/AMEIgSbKW34i2cZGPZk/NnIlcHn
PVxriiZlJ5dW+3DXZEsT3SBqDU+IF1qaW8nW4KIIz4Y0ug1m/CesnR2VbGm/
rctEn+F8nvdOOT4MLSurNJu/rGhO4mbVwb9FsoBzcOzxX5JoHb9iWteq916a
ddEvmnmWvehdX7yZMegXYWJ1V5JZ6W4V5jfk3M2qLy5SMbd3NGLa5kpQEPPf
i6iSZK680L4ISbZoWaX4A73SU4dk1jdKnLe8bCqgN9RZGLwxozODn7rVVVgZ
2McccufLcTxh+vR3aPzHQUr+XkjnuB8v+jm7bEr1Wba88reCQ8UxcAG4RivM
jJ6RRBfX7RFQrpbobzN+FwXNcmyq7ONUaDmDfNXQFsnfRqWrfOOqASDPoea+
1MnEg0unkIfp+0qtWHlpML+wyFzfKzXnUo+8SCX9MQggX5wxb2RD9KU2fMEj
b55fuGWUDVptnzvMgv/jEPG+jPKv+eOuDejxWmkyeRFbWED4u24YXcezIa/s
fXEZl5pFtDbJvbWeLAgasPsN68FAYfJSzCgEq4m6WrUfRB9vEzmCI8pkZcLS
KO4k1o7eta1/ySVNicslsHm/sNTdwTGHGeR4TKAku0B3aGcIcBWL2mCo1nBD
hPpZxjCaREqbRzeBCGvw/F183J+Jh4H//zaQM/flsHxjQ/zixi4ogMQC8YcH
ffurWHVKJH2wl6I3rqqA2FHLHhkD+4qlpI6Tw1oWOq/Wvg/Yoxirb28CX42S
nK98BYE0hqtJYjX8LM5kiqGm+9KHUk12LMXV+yfSUVNyJYBqENwOjG48cbaw
9+dItWe2a0yt3W3+cXsuPdTiJiqAz89kPbJ06DBJjMEWKz+k+Wn584NbgKXr
9jgSxXaqQlRZ7rG2gVa5TMi3CKmU00qqdwLxkCOqZSlNW78by0MTnqueoovR
II/KH66VPQq6ZOaosE90ANx3tMOchmDhvvifzqKXPudlhxzbomAR5pmQshbv
L0wdfqNQtprlulUPy4n+vL13Tnr5OxnMDU1iEcKfOdUSh+u3jlGUB9l2jZeQ
gJOV2weefGzJSTMbEjY0DOEh1cAdMV2KfJjF/G4MNYTMeagDpx4SnyCHVS8T
yEW/cG0Rh6P4j/CNzI2hXzEt/I5jwV56HGTdromAw8xMv/V1RI4hEkSfDhgr
J7yTau+o/mtGLb+0uY4kcMkKthX4RExRXP62cdLkg5hYFG/sR77gZrtJDUF+
opy11IDDNwdjih9B7WusrXN4ZvoU6n+q0S5Sa0+HZ3Irr3nccRsWs10MWj6A
RJDJnhhbZ7Hge8Qzw9mzFhCYuDp3AkEiuKEI1zUhZGB3V9qViY8MP8LlDZWe
ORmol9OK+cN8EGHGGF25miYp6ItynWi9uny/mHOdZVybk+d8TtwT8oudh0Ww
c04KNC3hdVeHw6grpZdu3ZwvJG3FQIoLabu1feGkSQfWaYasCWB4GiBXgla0
Moz5m7Q6gB7yFJunjvou00veVD7cQAAeiEWY9+q6XELyjoXmg6gAUJeI1Zek
oFvUfnGzY/KlzTHscW8swIcMNH8SJRk+Lo8wJdol6ifDn5zkjty9Kdva68DD
GnW1Ue7bEyFvzHeoJlTdhgaHuAJyRQhnJ8s+PsAnMXtuSbB9mjCW2TTAe7Qy
ejuq26kwdd5ys4YiPn4ozY87qPBqnaDnrn/UMxBaMOpby0W4GUpntTYyblKj
MbkBc0uNUkApFQZDGc45/hke6u/43o90vgJHYlks60tUmouPNTu1W68ui2Wz
yceW3LC/sw7XIbxTZkrCFnqUlJvw6SC8kxq8i2y3yECuTiwYkDVT1lIkR6jJ
SRacy+rvFyNxw49BHzxBDNv9QaiORiTI2IolkgWQX6/K2vI8PprBEvi2VYbr
iQHwm6XPUKrvD+M2q5RuG7QNOQ/0jsoZOXxLRdYfEChfhyy+YiW2QwL0BmtN
WA3i0L1zoaATrUNBEyw+PmWPSI6d7slHc7C4CEoSe20O5DHkHC2an+TYBtHk
FufxkWlYeo06+BQ67j2XzgzjcYBY81hjphFN4uVnbpWosvXM6tP6I5n3q+zE
2KHv8XaROvHfiz7VeB+8qxbwmME12DKILGPgU0BVYPwgxNCIlnDEKZI7hEXT
k0eu6LSprxdr5bOVjlkHLdhLXiOdMUrZxIQZu3Qqr5U67t0tCSACNU0zVVit
b3sMvFsu/F47tbTtXoze7cXYPIK5IKS0QNvEQfoSq3ZBNk/BuxQJ/z1zJa/A
FlgZE5lLwp9dW1m4zglqi0mdI3CfdrrJV4yVwwKtM0P39dq1UccLtak5epve
APayEfnQIPbH4q82uxQ9GWn6ELv4RYZxj9DA447bzPY7ZpDd+xw3Up6/JLW2
Om8NtvQoTCLdoePv0MvqapeZytiUuQnUOmmPw4l3ijaY0QBqIPQpWTIWHbV5
OfS+xz5T2DIMCbYzHe+bljYDjDrYXMSEkMa9kq4htShKqKsyzZePDBg/919V
YAMvs0rRYCn3nyNyOkt5iQ40LJ32zy5+WDEFGYVP1Uehnhhqk1ZNHB6K2vx0
H/GNKgtoFNupRvv01WQtuVx2Xh4zPah2OxmUyfeI3kLgzS3HS8swyDRFrfXL
zqDCxxEZu0tYrcqA7U5gKmTHCYnhAr72au80eLvuhLQzL0RYQlXugtyb+LUF
ygF8i6J44EdUfDXgzINGTxNYkAf1YqK9V8Noy1uDlRKCDwWcBO/rjPQqlSzK
hxO/s5HDlfsX5vUFmReAUxgvhrJGa2yCaB0xmeTUNjFJZuaffnn3oA8ZhfwJ
7oSeCUfk6d2PO1t6fArcnzVXs4rwdJKe4oTYkUcOZv7+9M4ei6QYILl+Z9xK
ushBd0AUQC93qSkz1NWpLFxQ/mNcxPPseRfW38mqAs3qAr2b9X5hNUeEZnLu
TGqbhd4KzyeJ4iLodZ0Oo4EjO4bVg/hFNzsEXVLXTZVgumU8akh4mC8AVTkg
8mBiiMn3Zv3KDIV6ZKjfzpMdnyHQ2KdF7ayGT1DZ9JxqOj3WqgU3ipBkdV3u
d14GH0PbC9NtDfZxpylZDKRNaulTiH1ATzi+hAK42HApAIh4QxCEJvvCcbxd
DdnnqRH2tro8e+Ea/CeDu11UgrGU1GWvJfPwTEoUkTWJNNJ47YjFskxVJfPs
uT6xBmDoBtTKaKzOGGVTb5o6dnNK8gw9vW5+07IxaTW0i3vJkrhAyHTIDosg
VPoqvhhW3Z06mRE8xni8KATCoRvN7kiVCA71U3dGVZ/fgvyfv6qN5loEn1fF
atng2Chb594E3LOalTRJGY5gyR/hc6jxHekHdmmDSEp23NTt0FnkoJ+o4Vuj
lP8WbMFtlwi3pvdrJPg/rl3VS+zBh87fQt2gpH7GgUmi4i0e/0QzabhUEHrk
g00xretFCNQMaUJkNFUamR3s2tDlXyVeSkgPTLwutONWukQP6QvLZ0RTydUr
wSzuCSYOgw79z9KgVK5fXJwDP48UcSZyejo/WMVZG1zUe0B6n8gk0dXcDzbF
i2XWuIF7nubsk1gTIHyn6wrKTPXdygxBQ56wMNjG7vI9VqRgNv5sflU9aSXK
+Z9x7HujT14YlYyx7sVJYLIhWdqW3KQc5ZF5RdoQDr5DJf7YEKnFfQuFXe0B
Refw1xImRPJG5dkd7j8sHVZNElzRVuj/0Bv/lf6y3eNKLbB59kqKFxy9mrQV
Z0tcZSgjAJlloHznRJygvVzg2jMI8JWIeoPEIhoj6xuLgzB1RJRx1q95JyVA
sVPvZVuUzrQKdb7EM/rXb2ToNRFfW7FGJd8reE/Zr73QO1fH/FFtR9nejpq3
snyj1GrssXw4YnKtpmHlWQb5k9IQXZoy3Mp3wmDpg6L/iB+Oxlyb+340D9CY
SIn64AOmSqJLVQ0aIoM25adYtYVzFdbVlSAm8evKqrS0Oj0q8AmFohcpBBDZ
v0aw6xzIoZsfevGe+Sq9tb/jWM/ig0/1DAI+wTvnrUnCC8y6FLwe7ONbSQrC
KD+o/667vDmMM/x3bL3o3HJfeGa8lUPpj3YySUZlgxvXQ+32NGIxgulLyejf
nBV6pTdDpABcQs/rmfGvfPyldIIYpUzlcEtCVE9k/f+Ub9CwHXVtOkIUkdXW
Pq31GiCY64GM7RGJBb88HBKBQJO4Q4Jagj0iUP+dA7+nrBWxk1jsGAFbxgtv
NPHHPIhXlJjjOk1W/C2bvPD/PAX/4UdH0piRQBfZLMeQ97c2ZnCzozJDs3Tf
Sj4PxfXNYsewd6G7J+nalU9ScP8U/m+FKlnMwptNzsYbu0/sgcMaQ+Lb9oej
0yFt4oAmdEsdTeztEFGUrfYqSa8DeXo1gf9cZGZls3AVL5kQIn70VBRVosZ5
p7a+Gc0YYdtyJGuWQK/LcNSwu1YTSucf0nqUCC2YnrwNm6Ir5osa0bXqhanu
bR7YqhrlvJhWC/LPvUm2rhXSkfxwQQkO82sP6aCMj0sslJpuvTtoD3y+lRyt
QPrnSSw5Z1jcPIho1R065eB58wpTTnLhAza7NxZeLRkuNs0JB+csSPHPMPWA
tfbH7U3WYn78a0w/KTgsYy/pDPzEGSDrLij+HxoYw9A00Mc9ZcLoRbp6Dj+y
dJritbGQ2uin9FvK3bJu7z6rQKJrb9Tj5QPJgOYYwuwhf/9pLNIisHm/BRw/
IYJ2EfM2TZLjesJXfA5SOaVfUKdRf0TZlnFsRXKaMZme8N8Da4bPJAU5TQPk
2PsHJMV4l+iYOrD/A6brmuL6o8dyZGTtoVY01nAM8jVgRSArNyfv0x6ezUc8
vhZai+c1uFphIH/YLjB/tMrB67JqfsYvvDf0dxg5Qtoce80LnFwELB06C1aG
BgDCv4zTVJpyMkrL9RM+ry+ZlsAjt50KpGFQ8suGUK4BJ0QtDXarkHvm8Zgu
o5TF6L3L2EkwiNUDbrTQ18tXTi2BK+Zq9xk5/8Oj1XKa2JuJ/NZxc66j4RIP
i1PiBnkZSK6PuxQ7SZJngtmkctFmqaR8Ilfq+6eJIPs42izRrHXssQ56ehLD
JLM9I3G/+5/EHoyD5h/zZpYQybATS5s6psoSGj3H2iYieFK0DkR9DHnn1CCc
d69Lpu2w37VDVuwyyeSif/SShsotgCNXW+69wbu6wWEiI6rtARPc6OTVeMaj
2/VhcWLWirluCPl+iTwe0NBXQSrdChkGC3x1JunH8BCboaXc50BmvuvmG5nt
+upbAQwmI8okcoG2yjVbzHyXRgd1DpPLfwao7BVXDoqdcmNkNkO8AwiHa+sF
Sgye2A8Ld73PREXRQr9TCXt01go2fKIynXe90XwEJzm4q+/ahtJJZ3+folw0
OVXwtFxESjQpeGC0L0u1z1kSF9WVskHv4QBiJrEQdD6nYR+k0HH+yiMq9nQr
79IASfGfFrlhT9YRBYqhLL4Z/7VdJnlFZB9M0YfK2QUWcFwWkcFSLSqRNdxq
EV6ycQwcsAEzsd+Gu1BAo4RTRMv33WpRIQ+O4kBIy5kElX8WganJF3mQfbaQ
eB3CCJVLeqT5t8d8c0erWiPZr+pe9K95wgesHReMl92sl9IUXaQXy1n9AO0t
HaUuxnvXyLt+GfwMA9+KLnrkwAO3GBSR5YbxoIRIObE27la82UWVZrf92Uo1
V6aSWmVX+gAgAVTtGh7QknDE5/5JHo7X4sKZQUGHLGHe1/dhA5vOSAkM+Q3p
h4ECExL5Qbt8b+y1IPQJwf6tLpVnozvWIgZpp4mJJ7bS1VrcslTUCs40Jr0n
bcUUzcnGC2crjvSkGx3/Q+8i7ZU+5OTgJQd0XHJKG7V21UwLsPkY9MK9JXes
9ojQLsqj/T3NFDTOcmVXIgpL3QS5WUWiK2+Xx8GQzujzedcZRluGTQpbNkAx
Oq8ENUz4aj/LEDBMYrEGG3nkaXTbjwR24JjHloWwXLRTdPQLDU0LtMnISTnf
h5CEG6qNl9a2k/iFVJGp4EbavuDiPDpFgWUspSNwIl5xvE16NT6TC3MzxRzY
1GYY8LGSAAVjBo7svgsLM0aRAxpz7DQI1HnKxI/lpSypsLiF0wm/rEQeSzBJ
BC6meqtKkz63dWjNq7g/jX9o6NG4qWNbpZBnsPjebUghvtiXD21y91l9kamA
gOj+w93IqF+bZwbEVoROykZ6wgvZOqpbqIkAHevJqMj8bhO4SUvbf2Csw8KI
NBQKHpK+eeOA67hzCuYrf4woOH38P2dW1ODTl5wtNVXPhiPyF6RGVYuRvQF/
Mb90QS9bJVkLX2a3gCWoIWK94zrctFLWVHA6YdogMpcXrrHt8DqhVfqcgNek
baUTh3ifDlEd9RiKCQhdaCpYI/yxIfqtImH19RBC1OFYZQ/9gW7C7FXj2hpQ
P2asnzc6SI/22oXWLjZYq9UB24w0iVgvAM6p1PCTNhM6L8f9fzQ10OrxaXMl
CDHakz5+wsmB+p4/Oe3EE8W2iC0G3fVUpFBGWrTkf+y3Q/oCVg5L1IytksIl
NaPzEgsO88Q5DpvpA/uIhN9VkiTKxCjZQDTALrXIwhSzLTzL2hW5HNfelXbw
naSUyM+JGg0LJF6POKzNNqJqj+2MMo1ns1TsboB/yDCIZhrIlqHgxb4KzSVH
AR3decXLsBHwQEnhT9HsI798l8LvWBeebFkVOq2rTsrbA0BP3duLjkufA6kr
hEz7y2t1KtsVD34L99SmP7txXaXiGdENBEffGMSLbCffl+C23vQz9E8rIQtN
alw91jjfBU7uvypCbmIcZ/WJsuwbmfSI2yT84yVmO3s4FiD5X7Dfw7Y0khgT
/vUI7R+8wI0zhjzreFexKOfBUl7Qq3lk8Xu/YwUEjSN379yv+lMED8PjjY2j
qZtu/b0790L5nLWtq/ctAdEsSXUaV7UM/bSY+6CtIHj+UHz/tU1k/yANdfXl
eZMD55LiEP8DmfUH7MuZxktk8M2SwO7R59slskx89KYROE4pMWcQe0nfD2xR
61deDtnwiLwCEHt3sUXaU8PcD+qSZBYMVS5bLiFJCbnLRYjVxO7/2s6fdYWH
i5/kQNV23dn6zQOdYvYo+B0/pXECHcAc1EWxxl+fKV4ex7G/s0VwiBDWuImB
kYKMVPRaUmP5CIrLxCV79N27HcIh8BMxxOvEQyzY/1oSsfe8BNWUTCkAnfLW
B+n6wu+3zwPQK6UozkJvABM6fiaYYoaM1RKf9pIllfh88slH/ySDjPqhd/0Z
6VDTPiC6L4SsWWXB5rqa8Xfh+E8ZRxkAtJZNHKLiFebe2qPzaqtKoJpOom52
s7L5Q8SV86Q2yqefFb4jKi/38yIXPlCUHpDUW1J0WmOSO2M6Ha2TMrjosh0K
+AtjffqZ+XeD7ntYcQN5uhuBQGIx90j8K2G6tp4M4AKoCNuoPNGWDg1iI4a7
O0ZdQJXy4zQyLLT/dDKYTXJ6P92o+JCBf5ZHDjMujUQjSAEt69VjoZgoRilt
z1UUdEmD4sP+NePPQUK9aV/GxednOTBRf2/jfFf4NZdTFMSI6U7C2caqJbof
7VGI60hGZmeTgHIhrNqhZuEbQwV+uakbhWJBz0RNit5iTHfBV26QNCF2+qYv
1bXpNaR2jRlH+Fqkv2C1rBnCQp+TY93tzkMVsfM2/R1D5Xpz+eAu4FDR5pqe
4Cz72ZsJoADTimpbrEFVwhl+fCxwJRKHJQwRMeVtaocX1Jx3a2yGayOcZsre
rALJItIXNrVfaMkEzqBJuxEpjEDhLnpZ1Li/Kg/7Wi3sr4cWqTl/aoF3na9J
43iwOZdrvz8hyPVFwPCaPk/ONuc5NwZcKyKaoiwUhfiBDK1d0FzH2BYs/y2F
wnsSFBd7mqz6B0ToAEtC1+uF3deAyFwfe65Y5GYtvgHpMgrrWwVJjTnlbgOl
j44KsXoTntYIZDVmHpLNtbgJDceUfYt4Kn1BfM2QQwqCY7wAvhExtR5gmUJo
HSpGTfRzCT7cCTBPUTJCSKJEo+Rz+k5RiNQ1CGoc1ULAiLdSDLRozjlNlPA1
AFQQ7cEVZKS/3WVH/7OBKPfgkqSVQ1MIXOG9CDdGimfLauu72q/3Q3DsOR5F
BtINoGZMXwYXtyFJljLjqXVFnHA0P+cdKFhVCcx0XooRuS8p75sZAZtCUwd0
CAy6OC5Oq5VbG4Mdq4NwqByrNuCkwNy6z4Fsrwxlqj5xq9+aEgRY+xtCmY/4
D+GzMjMnLeDh6j2VGNltJMN7+0dwCF0LENvqVPizez9kkxY7bKH+Q9uqbv9s
xt6861+jtgIFwPJ1cmswJ2rVVlYENZf9UBi+mmzvOtu6Pmh30vcCbOSaFLqy
z1fp/FzJD+zDi6awVAfxunTOUhFw4me8YZr4C3GSRksOPx4QnfhG+BEkkkmR
nAPK5dWMmsY6mBmhOzOGbutL3UqkksmXS82oBPi2W1A42IhkDJiLbaWH0qAB
i4punP0Ko9qYjzngpnfZfBv0+swuwXkblyAm3C0R6MXjRc4YV35pZ8P2E8NJ
KLHtGjjxasLtkkt9MpBJvjFNIEHRS7TreCy/6DhttMsIfgsMJ/ysQOf0pUNA
KNdpapt74SkpIgUOTdYWW6MLNBwVNwg38uJn12s+0LrvcIk7xnvcgGS+YrMP
90lhP/c44t770xYumixE/lu0vrmNCK/SUt0A/H47/ZQJWHB0EQNe/qAEPGjS
ePI19nZTaxKa5ZgpkRChgpHEjX+HSaTUWM677gXNX5CjDmb3QKkbFLSf9/V6
L9xdeeJxSpOIOf3KhMW4GotRmFLGmHOdrSpkMqGQA+EYNclopUMn/hDe1jlt
vTdLA6Rri1tbUBTHoqxIxzkNcx9kQU2HMXUOspwvKrzAYHyMlU3V4ioA8spo
cdpmNW4IpYY8O87NiB44cMs6EHCvmsxZEwCjMFAcYRD736Um3J2DEXJtAKTS
v0JVyQDK9TeaD9HvEPfePnTeb15L+h6mNt47E5AzWU8G067wbbbauN2CN9qb
nSbH3gBI04jOlvX8umaiNZd80pV6aUa4Rxe+UzKOvCIpFZHyHmWhebGZWZrN
xQ7ob9rTs4GZQLR54oCmtz+7qkT1cBHZn6IAe0/DOE7zk0TrNjCkhtGyO2tl
fNTuO9FV6QypbS3G7RTOL3aJHg7Y4uUuN1CfwHeqftke/JQWrMSg+cKZwfdg
fVUQS/Xb7/SbFe1cx/C9V9AB9MCLkN41zDBuqmmruHAKiRqd+A3l6k3zmJQv
Cq2FS5ciq6ue2qxbMTy/YeHb0G9SS8xYNotNJ0yYuIhDNCVERvhZd7ye7ExV
Ol5gakNsJLKltxb7STIg9UwaQXSs75BaCHY7mdAF+T02bvkOqj0Pet2apqb8
o4u8DvyowFzG6LiAfwzfV6V560Fe4znmjBBGUYVJOsIH5KaY1kKlp+2BcKQr
1VxqqXHzZVDC434p0i88/MbEyoyFKhrbR/1sS8/tkX43a9agAYHvt9jpzRHZ
lQ2G4Z0Tlx0/glpQb4wIWm56NT73tP/rLUytgWZueEKz7CAIrPLfFdYkMUKb
V39MBSJc8s8RzxeoqhldVT8u6pgAY5sO/7Du7ZDnBC8sXhv9xDIe2d14gnb4
2K0R5EWO9gt6+ekppcG8GUhoZdSLtOMHd1qo6Z/g9N2yiCCwT+es27KFgbGv
kegB6gN/4txrxwAc6DkJnQSL78H23Wb5QBSnGe7j1fuWi4S6PgfGEPQHKbZS
OBVL/IL80MxjI5LWtCPtAgOyTCWDItCUPfJewhAiEQc39IJ8HmAQ2E3t0KD4
p9nU+Wch4ROqDEhLR+Fr4qHdTHRpCAhL56ZF+8QS78yoxIQ1OoNJJ2xBhUp5
S4qf1U6ckRHtMHCYDlEX6cPTA8wlA9MTDA4I9kUJtpk2jmXwVDp9EI06IxjB
sipwnEn52N2x3ktKd+vHmKHUim5FYDkrxgme6fRQFeaKGl/RodC6pVFKJQA3
o8Ff8mBB9LLAbsrRgIASclImsE73frS2yJwjHwmfgvtLAfxqAtg+XwBYd6zu
vsnqKbL1380PUIOoEaaes8zKWHTfaG2PPNrPQItrLWZz/IialisfQ63l1sbp
nzplXICpKVzg7JiuHBQudAWpkzaHljgXlQ1B7r8LtQTEzhfb2GzFHU/9ljiL
Bsn9sP9RvxdfrPc20vaRi0f6YIbTUMcTDDU6kVRfbAQ0SNPjFC+Xdta1BUiV
3cjvfzPGhjz2wQLUVpdIl8rqpy4/hwJkIKMlsjgSGsznjx1GyBR83SWbL0lH
FmYlg4xEFWHuztJn7/JgdhrwVFRsFXsZQ2dpwtjuLQuZABU5Fz8ZkbraCtYH
kWhESJUbow7pu2hR/wmReZNqAFPHeQJIZH33uprU8UHv6KYvfM5vBzpR5Z5X
rZTpRaK8HSYNqDxz5pR+JAN0/h02ESKc2B9HmKZ2G58ktuVfDvCS1jSkvkdF
GqOibdDhFnBhcQpaS6ZkSoXm/ZVJz/M9b62oBRDEiBhiLnrISpeWBRS72F+B
LBGpadNP9usQ234TwT2FEKuf4f4AhA7+nNIjkXjo4znAaBjFBeICNd8B2swV
wU0vWddt6R5v/6bi4YNU2pul6WlXs1i5qBFQUee+IUDfiVE2h2+DpD28Ne7D
QD1FJDVi2P0LiPT/Hr/cWOZrnHOIUICNNMfdNrJXV7nsL7QQF4lq8xSlTUjz
5pZ7Bif1OyB8IA/YMfObD1O6Rb1gIINrAbyeW4LwO+WF27BhVg0t79pgA+HW
6US3dpnHgPq4vFXLAIc4aDJXa9LlrZDwwSc2Ni/6XPTYUN2Ny3lJqziudqft
ruIWipd3Vl3WSrA+MLVOV1VE+Z/BaY2sl0RYPl0qehfd+y9y6dqIye8KIJQU
tGcFmtoWYM4CIlbYwC7+cODEYVn24sKlfvmmDKVrsLnEuYm1iXCMk1CNIf9o
nYsElwGYw1fRGYpdBM9O02ay3uLKJOVuYj4iTaorVaeZOJjTMJFXtrG8s1wL
U9S8FPfRMTTlE8SmHVWkehXV0hs2GkwW5IYSoy8ECcu0lE8h3qyEd8YpnYY5
vp6zi6yMag4iSjNkeN5/mWS+zbqf1EY2SlmfKN+2pb+BzlgQlzZRJo5wC+Pc
DOzI+rSBa64xuxXNEIbQLNWkZLbojNQgm2xZYwiu5qllOkuNX6Uv0QziRnZv
2sbwDGJ6pmpETEOEXkc7qbGE5dj9hMkM6IQd/XMRn6BcewV6G/rdLxEroKcF
eeIJ9d4fLpCHzBda4jk7tLmLDriSBILa/DTg0MSa9SO6+GYX7isuCyzoNnmH
AO2FJQtKpGZU2wZdBmDCfkDiNZarVTFL2hGnNf85UADHDPw94sR3KLvbwgq1
AMQoJCHTDf6itPICqvVirhhE8J9XyFKNYtMkhe+tHIxIyJhNWPZ10zKTXJ9F
d5gmVWLTUiNe0W6u5RpqM45W/QT/lXhlJWvSFqNKvLfswzR3ej+DM82ANlLZ
rJUG0mze0KiIn535OFaIhPkVsz+5wrNQ14q3uyCuWTHyssTWO422Wy6zi3ce
0r0920+ytszA5aZ/SDfEcS05zL4GmFuuz8I6/yw1Jo5AmMiLyuQy1/B2/ZPb
A95bWVtdGvix0fGU97SgZlezpi5tNi7QeS57zMSwCuH8kD6y4g8N2xkAe1Wm
5Z1mkRhOQOu938AqnEcJuQnMzTyQaPzVb62+rM3BlmctKRBfNbA/6/FQpyfP
UO2gCHkmuubMBQ37R/y0Tq7b4m3XeCDHrj+29XhOj8U7zN/6dJqeWvOFnmng
KwUg8QqPPJUzIHlndXd2TYsjkvLMumhDX7umZ3s26R7Z/54HPlULjR54ojqj
OrNJwowonLVjPFGS/9tNSHJh2NpxzNDEpm7eaYPiBANmXnFYNLUKCDH/eo7F
HYDdh+33n675Wr2pnbjcoTbMrNGNGoeZmO9dfFGjWbeqYWvVJdbGW/BdTxx5
sCApqd2hVbcHzt+VrRDbGJM2NqKnb0XOql2rcvnz1SWlJVQmJtUvZpU3eR4g
3tjeosmlWucEpPPU6G/BkQWcHos5Iwnth1nQ2kpHDi7Ra5F4h+5YH2KHApKx
mhN9FY02/YwMK/17FzKe+HEFt1ll6pcAQ4hpT67OavGinyOjVgpDeNCSvSBs
19Nwn9GesylNIrZRP5xQTKhDEJfAxjTe8a4uYkmTwnZgdZ3K727TpC8OuXbz
YXLFkxco5z3Jg8XTWhdIUXylDnOPJV4GsoIctN/Ukpm2C5SUk+RLPn21+s2e
FBsb3j7U2b0umCwAWgbugy4ycEhbcnAHdhL5/Ln2BvBqVU5UcHutp3hBE1eO
H5UpWyfxKM/yED9LCNA6yEPNkBaTmJ5ZlkI0NdW1SmnSY230nhyGoMhxPCdL
sXwZWhS3YGIJEpMF2jTWe61lpa1Fb9RM1Z27RdmfN3czAeOQwvNuFk0ccsNk
AoMd+nE/UGQhv1UeuaIzO+InkLR7QDWdmrwhPnnJJ9hmpMz3NQDKukEH1JEq
mGM2XDde2vX0xzS18VpVWAfgs8QYBzTXVOit/fy018NfjYOuT7A67dRlpTQs
48OGksN79JmwaTFQu+gZtiDcTyf++GClMFcgqg+h3rzsQkPGxSWz7Z0ochyw
bYsbb7Lqa1skHFWzPagYoMQsC6sK/tlHc5T65K1IHuebiIV2Bo35V3iqJT7w
xZESJJ0GKtLTvI3snLNpEymlKJyergqlePgDM/NaiIeyCAZURlQ4KxCl0o48
z7eLpYvEwVQtXFS0bp/Yp4MKAzdxd5CFIdyFH7ZT2jMUNCKftKCPjXWI/ync
QKLRQoAGw/WhUWdI3nWvFMtlI9FG3xmdOGo+AL5Q1H4kJ6Sg5+kSV3Oy5UKO
IbujX/VMSJYJaPFR28rZXa7Gx0uOtEQwiJDE37lb758vF4sCKxYcZbNcbosn
izriwAuQp2B50YolHbnacfNGLSTIyQuCBLEmcFFl9rRzzmc/4fd7I6x9B0RE
5cpBXbSveqIIuikdVsPZEaSnUD+9T1LhqYTyKz7xUgl2mMXvTGKP1jEjoEJe
9TnAxpTaFxCyHGtZNTtuJmGxvDhB5UsORWaKwqap2umoFbGGiHgk6+tFuUrp
vCUQ63ni2ERpPkkCt37UMjWcQNPb9Bp+6+5AnnekkYbrbm0UwHniP7zeDQRw
qXsXPD0+xk7Y614wh0Ay/b/lFCospkHuwfB3bjpdVlK+etj/SOvkdhl4XZ2T
pxx2nBvgE4kcigt0/C6wBXxl6McSbfxnL0hY6FQcwPXfCDKpD3fKqDuaYJ8c
lUIXTI+qCniUBcmOfjyo8oIB5++uWbJpTE8i4raU9w53Ge9XkI5Y2scNVG1+
vZl2f9oJwlw4VE8qzVZUBiOLdRJJnYhChmD1rTAmcoLcxnjInfF32DBuhhJY
wP6CfrSAiljUGAcdVp9CytHS8LVt1GnWL26zl1doos5qnmyCqzbqg3AdwZyI
PqPa8wrmLsZu4OwTIyVkKkfAqU3lVV5BLayVCL1pA2lmf1PpgpgW/Oo9VAe7
xopYpcVb/8XS+WLqmOl3Eo9a1jFQDHXufGRPifomkmWbTGupEEzsL+ys0lFP
Fo7efSQwr+i4lzTZi5u87EB2hnSQoEPIJMg7H/QYUNtmhOqzf4t5z7KEdGEB
wj62Hyqsx/gUeGKzh9xgUjWiZiAKE7hPMXPUGGjRpHJ+Za6DGrayAOj85EqF
5c9kydMQXT3ecdZjw8YRJaDaj+T3QbKilbpykqe6CMGL+pwGu17wP87PhSe4
5wbIdsV1QY6V6e1ECC0d1s41RIfxh3ZL38Kb3RiAD3X+iM0eWabHPXYCrgo9
U3n2TgrQbCayE+EepXzv4deSDaEeAKzRdUohJO9cEPcTKz/nrM3fCEgQAzfu
txMlKdB1Qn6VryhYxr5KD5/6/HDKKqweOYphdSWo/ZPAPk5GUmI0x9U1Avj/
MaPr7SaBbNWDXlRq/BxQd37sCqRR/8wBMEntJvyM/0L5M8nxns6Ouve64ffj
4l6Bm7hNArAzVcenNgkvaDN1E5tSYS4NrUIlS54guiC7Tr61XksZrv+oZjKJ
EgHvTKOaAXRGfWtAgv4ewENuiUdGZxGY5MliOmksJT+nBOBdKKlTiqeo7mSm
8GgLqvdJLv9QEs4nybQCxnoyXljk8sqm1/7mEpFHhaj+TWQUyU/N+ggLgvSP
IsLqmgvfmjcCjqSLGxDNAG4R/8c9TTztGyQ7DXt5zwBTuUSnLeIK0MsYgRcP
MGeHXVSuvCP0NoUmT1oxW1CaP6OHUkldwtJ3UWQpVqAorkq4eqVgACDIwFCa
V9TyL5oni2Eg1KbcGPitJsllUPlLQNMgPYgXmLOfttuhs8hjpG0/TSEZiTDh
xKfZ7AzLOrD/9qymlYm4+FRYqLRhvK5iTPR00StZhXp68/Zf7DxAbCXQKZsZ
R90Q7gNNYvbPe0Z7UdXurDKLsGnL1CMLs5iz/qC80A4qaFeMJklGJrBwgpCs
nR3kVF/d6ajkLQNVy4FuiD5TjPW6aZjkwqBlIAl8OftglCsN24ANslOB8qPX
O+Lmf7+BQ5uzV0JW1G+vKjYT0si0Z56/A3rTjaaXEXeBGib7Na8FHUFi6VQK
RnPwA+1+HxiIlLht8S5KXA3KBYg0D4C0UpB/fjvOaD0qt6oW4Vov2nX8Wx3D
PMeNl2EgkYzSRZxHNcfrB+qln21YMfc1sBty7xOesaH9cBDSnFf0bHPlmJLM
XqDx+bX8LNn+TKKhdQl2GMIeqbRdDlq+SQH99fsg6r5qm18eMjt4OCybsRTS
WNFadqIzSirGlpFsA+1peOuOXmPTFuOpzKxG4BneZ0JAYsCwZcaXoyzvrC5U
G80PqjlZ+u66uBD9D3Zl219/CmCf+GfeRehmo9Jd8FiNyX8bx/4AuXGAx68f
zQcWCHnSzrVYw1BLvji3Hm4Awh70Io0G5d1R2YQz5XT5N8zjN8PAiGAyNZ2m
3ODQbS31qjM54UKbVjgryVKufVlgZ1/wDi7yvPzK3tu25eerZU7OzfxYBxPD
hK3dxPsI8w4v95PNvxavivEk8vAZNmyBrYgEUyGy7t+Pa6Ip2G3dl8ATZRZg
aVXdvP/lTwFadpfBHeaoao9JlvHEs0PyuHvw66gnQi5ZGJY50b0It9DWU2Zl
QPiO+EYyPCMjanw22EcyD8OAJHEaRVMQ/nOjzSC+GJHeQcxr1QF6+WANEC+b
ssCYqhtVOpcOoW2Xgy9FuIn6NPtKAgWEENGDZujJduqNarrSVp1zeBgV28TO
svbGaBvb4NP+peEpMVish/UqCyIj2IiSe2b00VxmORhg3Z97oD3aUmsEsdMX
aGC0OoMUpoEpJuval75tYdg3TV2kCZfJZD+OBn7FxgaCM9cULtmWteyCY95b
WVqOqVGr6YyLacCEdESPQELzzlJylhiSQ/2yg3jUOFEqfBbdRl0CSsBh8BoW
0MMz8163uI9CnIUbBaF7m02khDVkv6GmPRUv4u+1iHNHnsElxoGoPGrCGqkm
Cm3e0m5s30yrVSwk6Kh9x0O4NQeo6tW8JDnqLr0EayeKQss657YUhqw2RSda
UYJ1anp3eApwL+R1ZwTxj1ML6egaj2nLd1KQMlDbySe31/2hGNIivSr71pgU
FdNhvClUl08GGagbgcEpKx5bPAYsTjkD2kF+k3uPQXNqSp4bv3x0NW7rX9Kt
kFRXn7B8r/EFLLzJPnv81yIznX5v4Pn0exIfTW20jVCogFH2CGECIUwc8API
WtxqOPVuHdSfWqvDNHucH5z7SO3hFpM7XE4FVJeqUSd3Eim0HPmrnztA2e1H
Z9zzyrOkgpmQ60Cyu/P+gAuTICQKT/P8IV4UXoTowgJqeaTyfZWNGLFxp75r
FwvbpyLnWoetLZwW9W7wU5NljOfhPWz6zEkxk2+vSz1fOQWnBCWvJYiM7iWn
RvyHyYe2HxpMNF9kL+wLjol9ZOiipb+NjgjWXZA6EoEdStMS8VnbrP+I/NhD
9GGiMuDBTfhQeZSkjHOdh0rehk/BmzNtS2OOZ6Xcx4PbKjy/iN0pqGQbBIct
LMV1QmQhUvUbN9HzYSZ4oJwachkz+yA5KsxjcAATDW8u8kwPSEoyid4dvAq2
H5BYlU2hdYbMgmXrrlR72NtEmDYQXxY847A8xywqE+FqpRSAr160+Onf0J8K
tZOuIJMwYgwFQim1Z0YaFRNmaifmAuS19gM8ezVVihkw2NtCVHWRC9NAN9Be
dVi3ud+GjWNEhl4PVxtLMUyaVXwe+6CMrEUWvB37TJMN6N7nDQhHBiDdam9i
rLkqyxghgut50qzlsWlm4v52iHJ4jLwYp2owyQgRRXmaMqXR7PbUUA8XZ64j
KnuudW1qoz7cC51Uo3y6O5rqlxB4bZo2B415ePBvkV+VbhVuD8Avykx6Jf1w
KfmBDxpwoJcdrSTKZdFO+XtufVs4U3Pb2v6iTDA+PUYCNO6neC79Z61ntqsQ
Envr+TVmyKoDpPwi6YVB9B1+pWZ9ZEW7V7dbr4Mlbf038561gM3kQBfSFqDQ
ZtfawRgAbjPnMUHLYmAOqWcx5Yu0PjMfLjzCNWUUkTcTzDiiL/T1ZapF74pu
DFUHrkp030afndUQMLqCF8YS8F3cp/e7hVVeX7NGOUDppYUNzrhAPjffhNgw
M24d51IqQ6YD+eG0NUjb1CuAwxFPBR2QFRyuPZUu06VH0udgaIUcQndAH3bn
MD3xxKZqe066NXEVCm/xTpmaJ+XndhSPYtIyQixZmeftQmpjKrB7nHdMxS6O
Bzq301RjGLd6HXxr2J2KACspFVzhOp7tEBdt7qC8krZXeuiL+CV2TFAXYSaU
ypxjG6yNcY6A0JWMpPpITorF0L0JiWdUme85ERd8DxxfhYW3kJ5zXO1d32wx
fXbZMO7nYQ6v6u2qjYhPRg9FX/U8oJhrX4jcApg91Erm5j/4+41RpcANW49b
CFGeh7upAPo2A47UtFjCGbqW8oh9cynW6EaAgaT7KSE5kUlm4R55ieogFy+9
LsS3rMiRGLhjIDTjLh8JC7tGDJzvov61/p3fpDZX7Bn9RWV5SIYorzMzc/vo
GGCPXJROHML6Fhrit5TWRrqeoJM9pZJZFz8Q5WPk7TfGt3mQ3DRvuoGCtFAh
0SLdleQoI/+X+s8YriwX1QH9ZCxodnm0ahyYtFw+2W04qYCo7LeNB5kk3mX4
DGU2Gg0EWGdsaQTDHgdrc5HoPn5B+/q06JPaLZoUGNixiNUlFGENGO9bkBM7
Chz6KpbIz57PVqu9x0mziM5JulZhbDD9/YLFV3+Y9HgcGM4SPnMbXtWZHPfk
0qNxqRx87xA4SLSFtSB9zbkWCZJEQ60Ci2ivcj6AtDeO9HEgo35r9nzmCxP/
rs+ogbEAnOESjlp95fGItpn6xPpWE2S8m4xXerNlDwBd2e9kVNIcnDwSaI+K
ZP9aWLqGUCwidXVhyp3c20AxSrxR0bRb6JvgHkWM6WDSGleuh2iXngF3U2EG
K9N3YjQjGrA8Fm+8NIc4ASuPfydsbzDXjEZ+ZE/xEiXU/ap7XrgVVk3cdW1M
h3A3odYCodc0nZimNkZfJHuonswJ6J7rfsGkk9tEA2mzi4JcKpgy2Khps075
49Aky8+kRPO95nzOW+aQIYDe0uxSUJ0tOQdaavRqUnOl3shgCK+2A/C1XI1C
CE3kqvV5v2oSovIFQDBebTuZmC8jX0Cl3Db0BN5CeX7M+AuZXuXon+cr1BYS
TLd1w/b6pQrCe/8qxjbPA70mCcFvOj2ko47wgcEDFNxIenctiTdHHhVdyN8z
MU/2+iiMYdvR9fjDypPA2pQlSt/VFB6/KnHwBZx/7MXRuAkvu9cQROKChK/+
gmEW1ZRORG/35cPwwxdhIMvcrG9gmzBgM7U/d68W+Anm3UlYjzLcpP6/aVoT
dvCSJdpUPk0QyWfcvDYTc9fgN0A96LHsT+TRzJA00mlylFRTVFoYV7ALg4RB
5E7ugvvf5Og3Yf0LoMIPiRxPDwbwiVtEdRAZPeF2bP8gnIQ+kLry+WeBcX5E
c9HG757WpIx0XujYS/J7nne1ESylkahIoDvF1UFvxhrYWqqnMswuPIrJ2MN2
dJMR4AejaQisXeGT/QNQ11qD3cPn7m2EmHA6cHs957RROYZHZzCFWhImK5Z9
+Gfh5KlpuwZocWnm8xloTeZfr7T8FC7FmTHjeT+hqJW3m1aFW6zI2nS+WuyD
UPMivo3WZYBzAp59x5kB/o5B8wg1sZjc2r6YUpcm0d0papooP47mh7fwtMba
ljvBWe0uilQ+Yepv1kd7byOfStdb5W2e3JrDoLc0uRXTZB8/MnuDz5VXiMle
Oi2DYp9nWRj0YeuizpB6ihxuhbo4L85HjqK/MJfBP7ftQiOsXZxtHCPKGD4z
MJFJ8NLqJ965aDw7Vq65+TeGK8fb5nWqrw04YDBa6LiMsODJMlOsrHO8Roa8
Skvpkye//Kg8HThurDLoeoo589SPcR0rkVDnbqNAA+dJxnQ0cNd/F5b4XLL3
GEUJ5Wd9jAY5CVqXxSpSxEK+fVl8PXQ/OOl7fyAr0frh4QvpZFsi+o1G0TN9
/30qlDqx2bppDttNcummZyITzavK1W+qn/WiCHsPkng1XnJYcx8ESAF9D7x5
59tiLHY/42mcvsFkt3k/x3IxO0A6coPBzAG3Bbr1DTr8RjxiGH0nC09hris0
shYhLBeQFV5/9di5zaDHeop2+0PPBWbDuLvTUryfOQ1aYxYzw/c8lfJRm/Nl
v05zQIRbKd3MZlq1pJc9K7lGaAJNeIpFc5zj+T0R+8O71cRibH+ffQtTaaZi
wWSInyxEAok2dQxBNUNclfhIFgw/EAI/VbLcKZb+KlDT3fBmzFZYRNeQ7Rqr
JV03eqyTzztFnsBFjm8H/p9IT4Eqc2is0QGv4Azrq07EuNW1QVuv++lYvL66
0MHBY1/HwH6OhMhQwSwB0RIx0flvdf7ibTe9Dpc6ZRhESuJ47XBDeduBR4Ro
c10PU9ChGSZhGy5C6uCJcUhnWEjgn9Bqxu+9VlXDcl3LTAL1jr7OfGH2EeU2
IdWyuyDoZC56QIAn7HzmI0wwi37wsZlQ5PXa6xkaqN4+/dgcJrwiH3zdf4yn
WjUoHPxjIQad1opARCEGcRAl9LUJms9rpqc3Gqz1YW2k3kOhL9h1RGWGynwD
/4/SPmxH+R/xLdTXAEACpsPwOyRbpp59qHBMSQEo+MPOVlrEbIMoDPh26ah4
eFBIGdm3e+NlqXw12qpc321KwJPOEv+UEgI2HCnbOsAhOgUd5oUnBwVYxJP2
kgtB8noDkVPtBpdlnRJ71aKfwt5pSVJz5jWJWORX9u8JfaNua6d4npZHnidi
VkLDsiuAc96UJgfrkMYWSIXQn0rqALbHjc8ebx6vXbdjuGCKzjnPYzn8wgy0
3IGrX0h9f/aYCSLuE8SSHu3cWbW4sBB/NFKO6Jo3iMPHkytE1zuKJ7t9StHB
91WSiU4KGXFdbZLCfrwYqUYvmTH5giVOvl4+mOrNf+Jwd5EWEo2MXuq30lfd
17OEt//PrWLBAcMQ+VPE4L8YFYqHJ7HFwI6ejavtcB9Lqd3EX5iZe5K9Jswx
fSvaXgAQT8M0UNZyjBIPQTPq232zPBdPvZRqtooC63T38uIgkvH2rht3SJpB
Oiwn3PWZiyGNKObKj+zWIJu5DXz0A/D2NtfT9SjILPPe7zk/iOqplq+UyNl3
gSE8s85zLSqoh9AGQpXs2I6iSfFAYvMgwNihKgVtDmGqkWcZ6tYwbb/JVlIl
KjP4QO6VixQDF6WsYO1RI/rr4w4eABs9y+DrT5wh/Zr55hBoRXdT1U486/cJ
3QHEtYTxEBIKWKmtrKJEYvm+enkslpnF6Dj59JJ6QI71ymgne91b1WdF6X1b
UxnGNFwJLzhg4bXERUmrxrIkp57s5CyL5+derJFbG/PN3th5+ttfTPJpsJGZ
WcJmFJP93UO6I0TmvqZDEZqQvVETWvK0+gIZcdLjR5GOBpQIdarHOxNOaJUy
5eAMtARoX6iTrCKvUO3aQplvE0C8dYml+PDlQVtJ9nU+DiDoaLy5+G+S1ZcW
C2mQLYYUAQ51XZBLNyt19hsacQXFHWOgOd8wDXy3WhsiMeu53D4514ZgkRVK
f2Cpl8oJJ3+c5/Cae9R+EKtlrLXOrVtjRkVk/BqzuxThr64JpvPYWMCfGr/6
VR9ELTvZQ1M0d7dkjE97GSA/6qNILHJ2CzW9ie/y367TkO7fPE9nddJDSGxT
CaFuPtaWYhOIxH5icn/GJH1QwCPl3HrtxCdoZdcvb3H91TPPJDfqwSOMz6JF
ROrFPRNEPkA/APMw9dIglFnhEkpwNEzxpW+FtKlNHHRlNyuIOpJCxvwrvM69
Fchl2REcPjBqlA5ln6ZUv/tht+nHzjdPmbo5VWz4EnS1tMtp7ntYnv+vmotQ
fN7YmsxnpTifoAHnk82+CH/ST1n6OONJ8in6oLB9SoEcMeyJTdt5OBke635Y
LHDRN0JfgBFCEIBccKJJCz+ilz67ILKc5tu+R6e7OmiSbWDaonjF9NITAUoz
kyoYrDfVxi80kiz7QPwLFgkoGPVPEOBcQmKaogI1y6Et4iTcXpGts3lfSAwH
h5BhvDWZpgyYTD53ratubbl7xbDeCLTkEMwvFPLq3qIBqbBld+l4u3N1UMAh
G2WuKa7LUgEV5E68a23f/eNnJU5AfYalTy9HFUw2e51foahDJAOEwZofKTEx
PRlIj+tUJWoJYEIUI9yHTDF2KndRdR35N0sA998eyYZcNsnD1KXPzFqQA38I
rlAl8X6CQ25llpJLQ4C9rwUMrg7KCwGRrds1QUrphIXGkANFTwspznY/FjS6
27UBXp6/PwAl4k1vuspFAQEofeu/34/zGISQ9yLITlEbSiavjE4Nm7QA/JAn
IYEMaYlXHEIvTX/UafqoY+32escpzKictmYVIEvehKopa8gql+yh/IXoVdm5
hEZan8MHOsaQyQIvN9eQUtVHMyDWUjmmlZJpwV5R6vlZsBUD0VZAAQhqPHMc
5UbRfTwZKn5Iv5pjca/TwcIotuf4VBNXMSeEDLhRONPDD0Vz8GL6rGE7qrIV
vaodr+0f3/myXGc3UBgq02cYeRm6Qg73yg1iZ8KR+IfNoa23ZlEBC3eFYjip
ccrbhdRO5PIQQnbdNT0XR5ZK2/E5OGv6POYu1qgDXg5uvwdVPf6jxYl5urMC
NsMJQ2+54fzZEv/6p1Ry2qtH9d5msSB6S/LSVBAv9626AyQEt2kFp27vewWE
3tzCZZt5HvI7D5cUyBZl1z3bed1H0nlslC731BozLZDsEL76RkfIGmaoqHyi
DVP8rJ9TUV590NvATImb+khAcDAS0RuM2gF9efJgCCW+TbvpnArSglK9fnlp
rvZfwmgmIziBmkVVzGxbFpmBboQJgvRZLGlaDaba1Q4u15CjqNoGwSEMTQim
3v7h0F/aTWaVaGog1sT+ELFsFVTM0RSKbD6XblzjBOubFywv96i9+nxH6Pgm
iEgZcD7ub2ScwFbOMDu7UQnarxPHqsO1C7r2jCzdcM2+2pkSv68P9etYiw+X
m9a1xTZBUhlWUNOYBE34RAYPHMA/W7KOHudPcsUYzrSlHNLX0CyAFLcIVbOP
HH5ka0SqMDRjogj8UkvvdwSStjhnDGK884oDzbcNgKCIeXz7uQRaXNUY0RO3
fPsWSbOstOLSH5eXkLBYY6TOhN9nCAD8Hk3q5iQPS3nRED9Lv9E9d2FpVR1y
809ck58dL9fVjuf3hL+ewD4q+bnKzG1f2tYc9Rz5XSHeAVHtw2WgWPzxxdEQ
BuFmDODUUY5m56Phm4YNvCzwEMVJM8GQUlgqQOjhQejPF9OGNBFe3GkMhAIV
2E6N+tl5uQZf9YL09UJXrW5rN0vDfAeBOlyl2RYv+Z+Y/NOyFWfTYpV/l2JU
kT0VOwlDdWKGBtpSpEEV591AtzK7Aui46J/ULqNJgZyq/HX39f5BlKB7pTUS
EcLdSuL4uZNw0lpbvOuNCJUkvpZ0occMmuz9pwWNP6cd6A2uQPi1ntQMifq7
B/6y2diWORvgTmzYz26/u4+kvcAgFnV0c0ntihSPenYQEoo9/vX+Gq4Na5KB
yrx7NbDU6XUJ3hCYatQ8/af+IpuLwOOWk5sTtaVeNya193ChxFouZxGR5JhY
ANrNL63NXwV673dQWbBCmKve8CxBGkcmdwuuAHKefo3htFdH3z/EnXTzO88D
ObisS2S35n1Q3pi1W7xnrOoFk0Av6aaF/93gfc88L26ZTT2cFhNWgarWa8Vy
KvsasxU7EWSJW2fnGe7lovvaEuh4kUOrx6lk1z/Gw+5HHsVHptKDXW8yLJq2
5RB4cPQWzBO8cdcEem4lT5b7z0IB9TliL+1s+5DRXjK2ia5rwV0s1IgBWPcY
p+eD+qwyr2QQT+zyizpDx8MMGFvxEB/cPsnM/A6RB6674A26xyosmGLCLJq1
eXBIbcElUr8O9Ai/MVEvSBW+jLWFadO8fzU7+iBm3DVvfW0z/8kBhsjZCas7
gGwy7dblttFQ8qtfHz8L/cb6oY/NBTkaUPHpiKAKRgWwIKDtyiUx6tMWGH5W
ETU5w31IYlPPAqwQWHsmgvzuuv3+X4YitZ6TBc6NZYZ/drEfYTzREQSNwbww
iXz4wcU0xatAvuRlPs5/pZdrX+OKW0Y+XCPb5NYT6G6/0QSOdQac/a8y6lyW
9Ioyrh1P5ysKRNeIo7ue4Xcz/4gd+blqsxsm/7sEwkCC1nMOxIOKVhlcL2Na
++bse4kuD9zXP+bE0E7WepEKyoUAZ3vhBGOUO/ftM85XplWpXMP9Uch/O6r8
SCDt/q86qyKYnKpKwFQBJiF9VGhNfCHhl4ofsBELFabTw2FNrMYxGr6KfiFK
MesQbbEHr3pQVPvv2v4nS0fcXOGsMtNPKmPcwDnTAO23nrsuM/Xoygkovknk
yyn44uDvuBtHJtTONqaHqpVGBPT6a69x2jLI013Q2hkhgbcG/4Ke80tRG/Re
0WahndzVTcJRMdPR8u379JQ6bHswHdRc5AHDe+JnoXsrBx0sIAb3DbQee+Uw
uPI1RV6j21Tj2zfDYEIFVpwds0Df/Fq3zClyWdczQ/arVzUYfvGb1c18pChq
rg8wyNFzu6WmJJuI/CyEBl9IbhL4FuCgE/ij+s1kp70MsV9s7DUlGSnRC3yT
pQJ7XoOaoWAistkH1mn3a87xWQiEkuIXOdsnYMZHKNSKOpACRew+iYjum6Tp
DIkaHpMlZe0nlD6zWN5sH7XUJtY7o26npeuX/+YRqE7jkIK02r+TwOMpotMd
EblDrzrjiCPMQpLoiI3ExhT5qCjMNnR35P/8h+ga0veifaKxxQu6fDVBjB/T
mP7Gjq7ksysX26Ip+M8HrrnSHMgGzVZl+YTdcWOF+VYKPS8Ycyy7SCAf1cZp
ZxkPQZSiX8KloK/O8lYcG/l/YWvg6AwYhYk7lKoq4yweptwsLkS/YvoyqG5l
dXj81I4Qi1yZV5IeMYBmENyHNYhJ+qGhbSbwf65aLj/8nVlTbiBCiZx8LIHw
HNv3AqSc3z8qhBQqnBmYY5jVDBtn4iwQWqbczm45Epi0RxUbpfTqD4zyEFud
Pac1e3vfe1ZjxydUsEh8ICmdQj9WBP87ogmoJO9JFu8xR302J8p+ROxxPM3b
xpFD0K4liHYC+Nc+SicAZQSgiuqks+GPm6dXb3rtoSpBhVGjmom2Ni3aYdqU
zGPd1RTOXou1irfmIMwRVpVrr+LtzRb5eN/cmjEZ5XubOWK9em47adZwmgA8
+dcRGt44eLVBhLKRBCNfD6C8ih1XgLQCa2ywR0vPOwc8Oy5nNVKsSf1pR3pR
p3XyCsQGR6KYYWq8u8kuw/0liVlqMZ6mRXIf3zrey6YoBQGJqB0O8esqcrmo
m6I0BLGFc4+W/R5xkvJqNOvwKY+eVp3op/JHoE1Lt5xptHFQM5/fUqd8ISJC
SXqpjyHGC9zKAVxk2OP6CE6NqzpgrIGGGVH9CN8UqHxRRrEhMMSgMYUUHh/d
qSxp3BZJnvLEPoE1IF6cYojtm7vu9MXi01Tt2iahQ881psWoCmhgs9JClkt/
9SXk9kU8WiKtCcEXPxJTSezq4T3Ouh42XsniCksVq7oVXPyeRz7JiTA/1nHK
PAc52KYN9zw5zbeTCW67Xk3BC+6avk54kNUdtV/lFdK8/T31y3Jj8L6xz/HF
hRRvU+yZnUivBaC35M32WHBAfIIwoD2zWxa7KHsyOGn3KQuOOBSTG26LOynC
iOVnO6dlnFgFbifjyiwbmUqzEHCffFyVDSfty+N2EnrdsKY5Ns/fQNfYzBie
TNMf6vSrLT1KdQv90HWQW23T63sam3qeAJn/7rui0GzEvRf6x434hS1lIjPi
+Tg74GrDpPp8BQ7gtq1G2VGyhRb5CC21ecPvHd3n1DTTMSn+ZGZAEG+W1TEZ
XREHwcti6STp3157XRH6pCGmaKvaqt9uNN+D7DKSleKpaxGrqLKh/2G4uUhc
T28C90EUpAQYQaVzzlEIohO0mBlguUuGoPNAB9YYnKOqkA2BvHhDSQBZ0p7G
ynC/Uz+WTxgcXCtBqTSVJO4V6sCUT80xYKdQPMjm2pvZ2jtDabJZSt5NAJUJ
9tlSxFdebIAXD3Ysw73hsXW6ZuFr/CWTQXKmDn4ORauFeWZv/+Iix0WIV2Oq
2t3n5YCJDXK2QJjBLAUvjSMI9+zH4E+KFzZG6AnCvZn1jjY1QHLG1Zs+nwGO
mu99MUbvQDqJsANMgmapkngyiM3y8XQQnzx49ytv2T0sLDL6j0aVRPlUfs13
1eFqZ2ELOxVugbR5DBQpbr7zrRrAj0k+gidnrauisbQVVFafyk9NPKRadQrO
U+3a/VqdQrvdPT/kVmwMM1v4RdNrE51UQc/ChRSM9BfuKbUsTJldbA6BTAN6
fcvpxTWwq1ziFbxln3Yf+WrpwNJW4qhC0cdYUlZyI1rGEp17wsoEl8RcEzIA
+5pVdTPRnEBJ6dxvcB8HlPBTUDdZKQ+ccAS7W9QPGnzLbixiwAmVAsFAVvon
ORDQHvYrOQTy+Nqo8rF1f0AUszB6QnzQw2EWsA1vVfWXm+JDjyk3GD/l/CZI
6VASl++kVW7fM8am9i7SSwrqbnWmM/zeHeA+qCt3vvKNVwkhry6iFwninng+
flgmkqawUhI+dEvuNuas5bRnbVY9DFQQAUDyFK4vgAt1xT+XpvBtA+kXUFbC
zOJwvrbIEeNGBT2fXgu398luTnZw9FgcvRkmtl/pZ/lITjsN9wM8Re+SLAig
AaZXR86DWUw/WllMHmAt0q4IXVgj/OYxov7cy8Ev3eCb1JGt5Bgms1a13F5L
I5P+lIpI4sEfe+GyZ0FhORB9saQYC+FbbW1aec0iY+mZfAOsJ5/Vg9ERKWa6
9HKB1DfQnEe8s87EdgGShuNFrtcJALzKiwPaVlGxlCE8pvMV5LvhLkNZFALv
MHX7xcOz6uKq7N4n35p5mOpJzpiaM1mC06Vk7ZdzIrSgHPBlaSR3a7PiZdN/
jiDi/esnM8EyqcWLXh5LwQwH5XdF/xNs00aF2EPESmc/J/H7i16S+tcWALGh
NRnN6AivFfq29BAeJ6XWJ3rWRS+vT4hEVIfPSoVbpWoxLq7Xnvk3qFPK2liF
HUDWU/kAN9Xu7/IPNqY8MHDUB8UKVpVAtEHsSL8OUKqV74SJkLy0JemeyOx5
UGJr/lBYk685XwQWVliiKoQOmLs7xs6xlaFkC6TAgF/4p/KodgrLQGgzwgj8
hUqBwJiWMwtKYKSMyh2k1SukcBA0TRQ+8CUKeUQ2cWoNGkqQlDQHNvPYIrDu
FoX4a0QZPgErX9EPFck4dGyNPHI9kZRtShAHdL6NocSgkPvSZuhh+UCH4gDA
9iY6aVunT5/crLKBQzYvuOnRskZ9D854SgzTPQSBjeOIQDptnCcowLLxiNCm
m5XzlWn6w0W3wPzcIppCeFjT1cGE0ugGxY95eWuHrshO8zuebQEfd1pdnm27
6SVnA8jTbnB1/yFOGc+DxzSwz4QTK2eb05njUD6Jp3tIa45lfvXWEUMI4zlV
howm7UsJgmrzRJB+qTSvey+O5vyZ5TmJp5a6eTMG3Buyz5vhNuNrAXqgqZAb
+QTzQpQoTiTyUEYrzSFm5qebdMkg82hNt0VPtNL55K6gzvrMpmoqMqQ2AgYk
Uy2Q95QsA/mK9Z/k0z9H/slEXS/S7noq9Xi0W52IjEOKcIzfuJrJsnkD6TyY
zOBfwdz8XvnBefWVduayOLkALlLj40CnOlZ0QH9QTXywfIXPIC6Omh7RxS/i
2HNSSboHyzsuhzOm+jFoPAVMfy3Zbfajnv4nc3Urftdaol+3owV48JTRarhW
S8bZODux+48q9/dYDgagFnQVptkcHhSwdH6FFjxtFAUb8SMq/xGM/qBdtmSh
SFSMM86bj39+u+nO+i+PbXWFYdzyKLJcFUv2JuR3dbQZcUp694Gq9CXG4p4w
c+4gYOUlab7l+hCJOekx4aLnnhv2UX9f8yz87VQyzlY/holuSJJwiUybhX2B
GQ4v/MFtC0USnaYq7tgbuyh9p5D9JmcNTiY4glcn6iCmAaRqkQOswDckB5Jj
iTTrJ8Y5kIeuoZQ/WtUVJL7Wihc/QbovK2T/j94mc9v/+YRDOF/mkBCdObtP
CYIM5jFSLtp3XAxEyijWPRHq1HCqC10PipwYIATZV0/HJ2P9cF/VJuojPYn6
WSKp1VTudLybU1NIvkSt5FTvV7qMSI39wkxZHsTPQLhLq1s2vfB69cn49reh
0SBPFcauw897em3UObzPncgf3TGC9qofxNSqHus5SheGcBG+dAXlXEXFV+G7
ulA4SO7RbRG8QDJ3Uiw2nWAh0EIgIsV5px7YW6kd+9LjCDj44lfCPHPOBVxu
MRY/SvBddqHjgIeeHoS4/UUbHdf2cbw9y09STEd6cIPRvK6NgcqjU4QL5l37
NNpJZ2eQ7iE+uOzmy9P7RzAt0BM9hisP8+Z/mgI4O0gNvBxT5o4/SLkmGXNG
QdLx/twTkB73KFT7QsTxbLdoTFp9YYeUJJ6o/n2TiasZMJSbXeYz+tpUdAwf
BRTn2qH/6cc628ZWSHay59nRYh2CzQg5ywHquTwAswWaOCGvBcrx5PBN+KzN
/vvODCRINeFGjb0CekN7qJE14qVDUmP180MhRPiMzJV9aeY9RC9AYhzt37va
Y3350AhQrYcOftDPfzd28ix6wXaxyUZn5CproLT2azQmpN159WB5a+alAt4z
8frlSnaIii/g4Hid/0HMHCWGb24ryPkRiYKjH6wkngZHh9QlnQKlIH5bcQlH
FXqZ6JBTZ66gS3mIAHzcCzF4KJyRikbjOVwQIOqT6SD1wg/lFwGOl5HyraNV
GWTWC46Y5ZclnScU1kAjexn+JSoqYjm8Or7QMFZZJ7Mt5BSQ3oTei3YM4Hde
ZsX/2PjxsFJPePKajBi9IiDmnGAv84vSYrJpWDRutB4gFSuMC3d28EmlDOuI
atnzTREwobDil+cO/wQFxHD3QhNkwGtsNzLlkk+8gms7MLu4EyADBZLKOMI0
HjXhqolg09hW8achYUg9oT5xhSaeZvhlznycDJR0Xot3GAhQK50vCDf7Ynmr
i7ZbHGGVjRUnuHxqt4+fqd/1M17tZbXUf1v/bcU4/7fuG9WWRxETT0EwdL/k
6/UQQ+72C36fjcNcYrGsSKXOM31z5nDhwn0QNwufdQawxs91gN/eebHgaydw
8GzdLgy/hCHaCI6DQWYGqLbYr/D38lf2K3Nk/8TzrCKHC+bv8savurVesYTh
C+fBP+0cZymVWkcur7o1WZh12dXPVCptsY2GrfWSG26eBSIDDulOpirYKGbE
YNTGmHjzxbJyXfTKxuvZbRDbhaV4m2wQGs91yVPCWnZjptFaOsGJF8gWXwLv
FIgffM17LlLbsyV14tK87Vl0cA7WsWxvcJ7ClpfjkMsNFpWWOtPglW8Ru2zX
EnfL8dSYAXVuKBTNXYBBAcUfntVF4QqaV8cEGgL3gSx0Ltkc2DbYAaY9joWv
Ak9lR3iybXCxw873Frf3SPkP/T8r/8VG8ZLZU5g5RuuZUg/LDgYFHPsz9E5+
zVzli5sCMgSkB7rZaPGqIviyQxo2hqcIoWc75HrWnp8LcLcgwcmFF9lPJSw8
vNYHyYd9NauNgdRo9SJ6NLJd45qs8dDvwm5np1y3+qBjqmZQdpq+CTC3wsyx
i6mzCZCi4f33L+sQel/fP/EhTa84oltpD7upRZOHAfYA6sp3qlkV+emBbwyX
87Dl6gqtzfbBLLIM2xHj7kM6MNjZTGlduB4Ylae3IvyGx7hZRQ9ZuVUtJWaG
M9GYQLlj5P56RaGeJyLHGFxn2prXPaF2i0RKIQIWtzS/N96eA6EEGQM8WmHR
AUy2Udtk8DKDkhtJfJud+H5slq+S3GaLWtUASK1h4NXFGsyPd9B07KB3JH59
Iiiw7Eq5ZSbCN7d83UqpEjKb51SVcmNx8IpsUY04pMNTlZyXe1dBdX1DaMre
QXp851oHWkxIiGjCLqpLLXu33wNr4124c6QdGGVcCQsHkz2taoeRKOOtBE5O
MNwC1D0mUzBkvdtsq5vohzX1Uj7bIDHEE7bqams3WvrXoXzMtQIzM0seMXFL
5BnxquWkly0Ki0QLr85rO4tIuD64hNRusvbszWJkVPucOoGyX60PR3+2i2VS
4jBiESCdV7TvqgcMfHez30J5mArahep8shG3/1banhsAIbHVYq4mja0W33LW
5KLUsP/eVmzXT3QWj2iOIgroQWRVwUjYcKYsDPtdljNRUG61yjXsPVdA/9Eg
cca9OvjCSkBy6hgXoN5ShOmw6cQ9TYYEbhLBeAuIiJRmJJj+LiRqtRHWhw7U
26VK0RkUaJ/oi/wziAvHKaNN1E1u08hLEKcnEbYZTT8DETQfw1bP2O5ekkMt
VOry4KbvGyr4XRJBGo92MheiMQyynhrSRPMsqKowZurkyCo1m+6YAiKjq8yh
5Wm8N4NCmTMCS35kSbbTI8MxXv4+aw+Y3oETFG3Mz3WpHJqyVRxY5NCXpEEK
1rwzlJRT5vPP2ysq9x2WUIoAfPfRs3DxILvI2dso+iZ1b/Uda0Rn8cvzJ5mc
6+8sd3oJr6fxD2RB5a2hy4axAqc0PxOaT5TKIgKIpRNAmwrZjf4nMCusGCoh
R4kDqtz2WRWaA+wl5QNwWkjvecV3WRHz9yxHY9RrMA9ABLV3SqxRVShfXi/3
CXPZbNE4czjJS1yD9YHyvuMwmlNVRSDcDdNQ6MDVPEsnbEFV9d0CJR9fBs34
yLm2+lvOv6RKwiOlbTesB4sbi7PvaEwhe8SHdjUEZ3Jvn0poThqlATltOe7G
Hn18PdP6PQR8fovVPlgvnxULUDnT2WNCeGJzZwKTZ8v8LVZehVMxkF/t13La
7eoQrZyI7gG8nCl9NMDqcs0gvzxkdepO1jL25D+Y40hC07X8s/Ep4WzdwOaK
odbrj4W9VHaLx4rBogd+X96ca4v+LwnJbKApyD5oKRg7BJLhyIvTUU9puSsV
//4XO5v6ExAFkuvfGZ2OvcZ8zOlXJvjMiRlWNrDZKMWOtyJkyw40okmRRxfC
8Wp4IqQ6uuhjlPxpa8IGED6J9s7RZ1uSupgOOg30OQYjTyIY9ZLCE6mDn8u6
Scq/QpL7U6zNcrGUHsqtfpf54N87tXa30D28nKWgwZFqWBbExyO2TMobRiPl
EbxUo6G5jCjTih4fxtKzHnpTHXlPh9AP7nXq24kW3weLuxDcFBAeGpcLToXr
WYtBmJRhZ6GD1VObft5hrvEVXty33+yR2fVfSDM0KJE5MWQS+JGvbs1u24Qv
A1SowQFPqB464AeHx+E07kY/ri0qglDzyNke9Y4LSGfltLijIpU+zqVgKmDT
vguWNKZM6T6npy47NRbQWFLqzBYflefB7/OFOo8PTB6ktHY/cBYplwhEoNrX
9ZTDpFOLQSvLuP6TqIoknXL7a8MRw1N59j68786CaZYnaNJ5SZVzZc3AIiqS
PTMEFvZ3VdIIGYuzamWN/0UFSS9yaH7Gk5hxx/fkFyAvmA43WoL7Lq2+ehsm
tutNFbIn6gALX/S74cEWVTgU7aETu7kUrAy4mByzdWOjC0rgtzbFfp+9ElvS
tHeGgX2Gdw/Vv51hVRxvGUNsF5rLc2gf+hJqvkK31O2B6wGwWP1t0Xt7HWIl
MbHHgdoQsVKaW11vT5zGl1j0tHPDBtixpAmjT7aXznRzSbSNo2Z968PGoiHK
7EAZXjIOzYD1lzFiQUeJDZkjzWfAuZizsoYVdUMYj0FUL20RMttonjESKS/e
TWLtdWrx6CjrQx83hEU92iVf0bVCBR4fpQVLAyhNzVtKm4Hnm6ajOGe7zEoS
RY2iuAdMnsILjVXNgCQmKmN0VnUOBcyVsJOYrWTI7aZ+tuMtzGo2BCUgRpqy
wUZ/hrWhZOvILLZTlIUuEqoaXFM74cWMK2Ncu08RxxtPiAkEr+oaAqF7RyLZ
/O0aYzcq2v7vh57yArg41L0nTwuZUC0XI7XV82QUEfjJje21NW2y1hB3TRRw
FUNQ53KF9hwL4HjOHmY/D5tsN6lJ955rOuVA878tSpQRVhdvGIC+Nx9bOxpS
PCZ+37jj2sdHWfRon3jXuSGEWyWy1sqNL5UAsU6aert2fl5wTtc0wL/NcsaO
IPIxfRq4yONvo5m0eOujrn+hfL9QJrZOyoX791JGVX7Yob52gMls1mSrA/Sk
0D9CwhymZl+VSvYSaDCYlilb9ROpUxqDWzRBCeWMWrlj501JM1ET9xOf3rWW
GC/RDjG6J6+BceXiyrKtoCW169eKBvJMghPFBQ7sQImzBsHywVJGnyZWeh4V
Ab6riHR7qAgn6FKjTIIIkbH24mnevxh8ldGKgDl+eVc7rhTuCZZEB4nNMEoP
3d9EG638xbX0AMNuod78VEYJdt9luVkv4Xtz2K90AA/85xlX3Q/xpQ6rkjft
8b/5r5I8bWYALC9IcruJeJJW7QG7kcIBIxq/3hLk9dheF0FfXLJEfU/aJnhi
XbO3Kl1MxBecoLcdcpu8LoHrSaVHhkKbNpGKC498r0uzPZn8UukYd+gYyF6c
KOGgTXXPNo3vkR2h0DOYB7La7FCM+pc1GuGDhRv810hNuaN/P+wf4wUIVeVx
WzOeNKnvu5k9hS1cuXqq+RhKOmYQnSqWP7k6MXlrk3SnDMR/KuiQMwaw6Z71
ILnBwPDYEgkBskZL7DF4geIAOlGsBpWFSNAtec5l9vC840YGJQqMGX9PgeRi
yFJIMLohnlnz0JJH4uJQn5eLi6ZLn4PDK0Fbtw9nxPJGTwsQGM/ebNs872PF
BmjQkD5SCwmrifCVOh4+sLFRfdk6wG7fwN94KglOGG4XZ8dUKz9U/2Q1TaEX
sR+HFTR2lVpvNAweS7LJHxvU8kUWec5hmFrejIR//tWJLY5fUCw4ehkRdPxK
gbSOipYZVbH/nClkJviziKdoeZQ6RDDgzae9tLvQ29hdCWi4B81Xef7bqisC
OeTqDrBeuz8G/2fetFBVrywSADLcnwkwDBqSxgMMjD8VW/7Mtrt0WvVZWoVh
aHSgsYsGyqLBMjjNYXs52/sP7QESdFs4HmOHh8GMeOqj8GAtYP4hSWfXiv4d
K7hZbHwT0d7PjTS6ybFzgemgjBlXlUB+U26bELHbBb5/66UEGBj+y2zLPQCv
anMhKBTt+5KxcVBJKZlvlSBlrfQlhkdrw+3Rc023mX5Yqsz/zJAYlVBT5ze3
DcMzmYrhNyGYS4eoT9eDDFDCG4B5KP9TkgbvuYf27JF3UZ+JonZWA/X7F+AJ
LDB1zaRzOFRbhYfRRF/AIs22u62zff/6bvw3F/8kU4UWkY3ahRoJjBNBvn2a
kjKZaUMc4HgrTh571x67NrrDXdG6UvSDfE6rE6/bwBMJ+ykGAxNT4Ga61Mug
tic71WDzRHrSoCyKLOpet9eiGxmMcbUKY+EMQqasgHEAzNVkJU7MUcdSWAR+
NHFScIIiMHqrWu+JluhUxiJ6yJtCppSki1j+xDEy9oBkDJ2MfBobnobFlb2Q
4Tf8Fu8RFKaQMgKBrwPGLZ6RDLyLtGBqJ3GeA0W64bEJ3675RQwdfViWja2O
LHbRiJp8XxiKIu14FhWaAGjiSYvgVWn1J+lV3HHqMsE6xGT7DLK0ElZdQeTJ
Dc6+jBsXsDzUcMolaKip+gOf+kkArsDRatjBXHTk8+NLmNZGdroxmmddvtaV
EmfsnN+BEMJhP0tHONn8KF3IZSKJEwkZb/pd3yq8Jcr+vVb/tgp1/B8DOA3d
3rT/dABuayok43PFCjGdRTuXpR67CPU/kB1hlUQcX9aBReZ29wiXJ6J6MVWn
dntcUNxYGno0z7mBycl66q8YxDEidbhLe4jg1F/Rz09y+wpQS6ZIdmrsNc5V
fNxki5W3jrXprdKC2hjFLc6M0uQuYYP+DPyFtH3j6JUjn0PvDZqKPxVyNC9C
kXZvlgFiEUAGx2J7y8+hfrbNTsSTByj3IuYY9B6eaveQCzzuDQ4LfK6l58W0
VTGgRz7F6mtLWxnNlCiy1bCRNpI3UstNbwP+M8ZuUNWwjfxZ7K2AVWAYMD0y
wrzbkg2NEe5NJC4vs+UkuDf88y8Q/201lNhqJdYF5wv0W4hWN7BgI3IVFYt6
m2UCfXzXb4iB9xQkPSW84k+D5SzvyeaSIlYO2OfiRxitevIMEucNYL4tE5SB
r14NuyEt0wXp/ZBpTlQ0L5X0Yq2yR0zIrWJx8jxcLtMU7ykuka+jNB37zYvk
64dNMZH/x0o6kq7k3NQrYPlfjRt+HG+IowXYA62qcncXX0TUe9v4RVvkFvH5
9NNgj8QzjOb3p6oBoFUm9mpjqhRBXnFrjeX95ACg0Q4OtauCxaaoewHxJX7H
alDaU5U9UZUqe6co5um6heZMQyeJyKOzdqRd85t19qqSu6K8IbaffGPf1XEb
YaiZ6AdEVOCA+FK5G2HzcYCakGK+YecZSXpyKcVphJ2MVaCo2uBBGTKx+qFD
M27/dn8GeIGDRJiDe5M9xPMD4xSyrkDkpI0t4UvHCaAxNTB6cD2tEiqzO2Vb
1Rr2lmIF8ZxpHdoT865mkxy+GsKO9hTxocoIb5ivv13l/M6Ddvz7uGHTfA/n
jZblrzgRnHgfjOblVRpaQIN1Ab2lcv84ynbsTy+WmpjbIZIYvS5bkqYfq+FV
ttGdV6x/JtXEoS43955OiP0VYOL2GWD1OzX0lEwKg5TXeah4BDvYWVS+sj9V
uvVGJtq3KKfB3w6+SaBlyFB0Boz14C0eMo214FXfrHALCOTh0lRUax+nPX80
/Edhgn8AToEzh+WxZJDau9VlUAYCHBDQBaQwIwzzGkQ83ijiYqJCuexGlJGH
8KSXAsIHJvFq4Vi5BJyyPkU/uR1faU4kurawTucNVPTJ78wtMJiu4yphz0pB
c/ThvBO7z7n8nqR7q78Gvv1E6NHDLcE5vR47G4ZxyvinR6vqaj/Pg2r97hiQ
1Na6/12w9upHQaIiTVbDpLVnJBWYp1ksiIbl6nNHKwkS7zE8f6c3OJwkCvuj
8e5K9y8arCrgK9XE+psyaIwHhHPorueB+GQYaOA/EUnvO7SA8dEwzv53sCHw
98eDHcaQ8gXyqKXBsY/VRuY3oIrPoQFbFnvDODnoCVnHnJUmD29v/9BODAQU
J2xIAAb+WT0vQaV1pkXsxKgDXAZgT53vKh5meypAaq839/v/X7W8FnDoOxk7
/M3sLuGdRtldN8u7P5V3SZezweEAiSdoH+somm3/6yNFCY4JBS3xj3uiCMJI
VFA4cjckHGd18WUDytwjagRlkM74ydtbEHQILGANER2QgK9ETxDnEDYp8UPj
Xn2/qDOuAfypTdTHJyGlT2h5pQneKDNvTa5pNWCgS7v1g3GVliVElZ3dX+lq
/n9uuarmwe8dA0XJKj8kV3jwb0BOV+w+6qNO01u8GmX/P5uREuyCjnnAwq8R
tsEh8wkSogciqhu7mMvIuZFB//c6nh4dwKezbNXrv5MAaAR/j/kyYEsvfdAs
oQfUUYgLR4XAN8szrmJMSn5wV+3jFHCjPZI4Tei5x2pKbX472As5/az0hfK5
cwSx58V2olqagakj4gxOtkh7sPl7FuC2PsABn+Vs3cZJOueeTKlUmyk0mtQU
k8mJF3MTXwOqMb8q/wtY+m8eNJ9ymVuLQAPVfxPE/iI6OrasBL9CP0Q46/jU
LBhTbtW3Zfun9fJmCIdN9HusazDXK8j2pKKBdiKwbayQD6G1ZH/5sF6t7SZY
tL3mGbjmH+W8dZ41BPsrMB+KdubA8CzQbbxI046beNwxEynhcQ8r4Jq1p57L
Q/tc3Jee8+XO91fdbmnXvPFZLoZmzyeEyy3VR+qgEs2ndFKGAYXU31jOOq0L
t1X4yJRSRAeOqFwjKgQUwX0chyrPLeR5Hd0zdy40fEOuT9LfrEB6PQV52QiM
7/yBI1RabtmOBquTXjfYE5AyzB4olRDleAXs2txmVdhUxyEBoiU6jluRjRS4
4JqDaJEAs1FNabERASFHeGP0bsWI9H98KwF2QCVuyfyn0YtdzyUtpC1yf+A2
bBtoCAe+CK8a3tiAwNGXMnU4IsERudikowgnXuMHQgL+HghEwQCbiJ8vy4/f
IYC5TaXdP5EVZtzIJZCne4Itvd/8wFsDWJTwbTWBdQJnRAEtMUKcuC6dwGTj
FF6NC3/7FI/nNsEqTe3rAsU7QdVjck4M+0cCrmh3peEpnC2YXYuPhXUX39HA
tqu6SMXTlwUkQg/z3F2n6V1iLi+AboFv3cIe5RSUrdMBSzAfuiWV5Uxcm9a8
eHu7yBLJWcdARhZ/LsS2T+DfbPkTyZzfNtceC8UwiOXYa+DSwnGu44C6WSAA
Wf1XF5CaM5hqilt/xczugKOCMka7EOWwcrzIcgL2/JKK0ZTAdDZGD3Wee5zK
P6S/hXAg3dwO+idKdT6plYlqmvw3R1sBjHxuSEgiB+4XaZmGFImPvIjHkFDa
fxvk2Y05Z2ij3a7aSrpd3ucfPPJ5G/8M+O3eKjHQJhLkiw37GBIuf/7YRzl2
+I1FV47WUtODN+vZ2yMMOjmtnWGz1NWC6GUOn6AquudQIqtF2VDR07fWvEdL
B5p99eYWlYwgL7p5VHZFPfIv8rPB7V33vjpiOIqXpLZ8+8a3joilCTfcFaso
gvD6uQRjyYEJSqX8ghaba1NMTkca8fYfx+CGwmty1ODnCOLnzJb6gC0kPSWR
hamHxtfVGPVCXuy89Zj15OGT6QfOa9jcF/CVa9WQ3O8tOJ7vfl87ebNgAYD7
3k4+O/y93j65VqKRO7UAoppvtbjDiJ87YF5WfWIZJbq2bSnV4iwI1Ll+CCn9
z47fRJHdPHHUNUx/b1KooXMakdVPiE3tz+pHr66Xuq/Gy2Fu/BatXa5YXypo
wkX0HWL9SfvrGGnZq3wrI+ncmmKdRDXBQ2aoiMNrfw7whEWAePRsw4FBdzZE
4tIluFmAqP5q2+3fhwvhH+Aop4yQJ2f1QWZxxKkPBIQc0Wu7O7KDPWzp2aAb
NOQYoVyqQYu8lvT22JHha486HUVp1RlIBu9BTMHjCg68yMnuURxCxfaK6YWM
tVQIgGRE0BzakhyAR3rLqkTCRUkTcjc4B3CYDkmlL8bv3g9odqvOtS7/2bd6
RHg8IwfIbyBAR1dr0YMTPpNFQOBjThCERE1R7wyGH/CvhCUrMjSd4LPbyIgx
taR/bc6ma+42lGJli+RPFwJNnoItfAA5lGOqWMnZWKB53XfbrKAzkAvXDwaj
H5b32Y/sPcVhXfk1FaZEyiLgCPRPJvBt7V+xOIlFpuzuYy8DQUzHNA9+eJfD
UVfGZruf8cp7nsUa4GOgXhTOGwcOaDONJAwurGTSET9TGc4IbTr2+5CVFHOq
8FLKcdPQvg98mJFaxqa3dLRO31XA/ljj8B5T/a9m5wDJi73qTQQado1ZXIsJ
X0K0qtAS24Ui8Z57B/A5mfvQ1UopPG24+8WwJqSg3Nq9tF/aSRvoBh1P2HVv
hsO/I0pBnu2PqHPGJJ6oadEHsxwhy/EwoQlG3SeLIlcw+tAWS/llN7RDsBvf
RyIWCVHwpjbop/rYwzhK6rn2+IoS6UOLaEvB0TLFCM/gJrX81H/R/pfpElzP
goJ0LfRFS5PEkqbWKLmEETHy0zaAg6yMECv/UEjJnXu6g7TtDNnN1xnpvKOu
BvkXWI6x/frkb+8HEaYJhDWg+ygPqMChEdtA7WIjQX0fBCfgULbvpUbBQvg2
NNkG9H+RR2lJFxjOBKWQtIU1tcbF5VSiCgJIN1im4ymCvTX/Ny/dvjoAmaBb
+zUMXTbCsiiPB/1goe+KT+OLbYaRHmzIDDJXYVIQMO+t/6rP4fn4dIdAeqk1
5uqwaiAiq4lXnC8itKaldrKpAvZJ8k33ri8/Yo9h8HEm8cQdAFMJsw9fGIVH
5goORhzapirrb9n2252TekTxZHkG9+ZUzw/GFK3CcSh1aNgg3Gn+ZY1PTyW9
9Amn1ILn+WupgU3VulQLRyBTf961L6t4Tzm0iYCizh2lXtv4TD4EQA0DokuE
ZZODiRGCx3rISlDzOH+g4ompqfYPOM2ThSUTeZ1XfG94lqAeIjoo4RHx/AUK
EkwKlz1y9nQSk4r3NvpQLQK8TRs8CYITk1AxZn2UvzmbjpK8Y8LP3BSV3kPb
KE/wAMha642841CLxPcbSv3275xsPhjdzvk2JGrIxMQkm/+50TKbjlOcbPBh
m1rV0jnmcIrTvcuDb7u7aKHJJAi6F28tnRbl3CTNpS19Y1KTRMMjlobiYQm5
NpWm9IZGK+4GARpjI6Mh/HEBU2zyVJCY3fKJPHy5QH+763pfH9PUQMDdH+1S
xw9yNzDENx5TdOhVd+hhck35dV6JBskswCqxL1HEjh5WqOdGzVh97SKLk5UP
MvEA1etJkkVWeGPCduQMLSXvFukMdb/DsF/9ncYwFcRK5PMelbHSseJ/NbB/
X+A2KzKq3X3rC6Y1F/IdHmRNroBFbsDEj7wdMQ3mooFeVWa9kaARlWIx6jcN
+Rf0H/3LVcaCBa2GQYa0VHpDSApnroBNCjTTvcUsEnShWY+Z4SdydWJkIXI4
ytVwZ8v/GGxpQu57mAeC4AscEDaHDWCct8ZsYeG9AmqpuD9nXIelkHSWaiyt
6mS11iB75/OuGpw4+KvqCOAP1yw6J2TsXJnlYg3JVGimUMyYir0Pateiq/2w
/uW8Dt+1/+fpu2D4i5l3UPy32kY8kp5dtyDrtiDJ3U63ysH5qCMRscr9FMmC
Q4R2h9RVPyRobz92TQWkS7CJYsUNKL0F3NNzM7GnFcEt9zUMVSN5hETR4I5O
TOlBQ42MS+lXQZyHskHCJDvJJM+jXJTaXWdyk/pjfKoubdnEDtYv+lembkFU
sL9uooPBsHmX7GvseurMPfRIN1uEfxyB2O9V8rZb0feXFFEEqhwwFCxaia5h
zjdXvBneLSJtliw4XyrrJE0x1P4EB56j1moYCPQ7SeF17M4N8TiBGBlueFnz
CLnvl1Gs1p3GAKq2DqMIR+Rw1AFwM623Ep5ysShCXOWseqsKIL+nQV0WROvU
T93yhzTFgMitvfLyNpIhAsy+XDqYcP4ALqSOj9MsreLhsvGzH7b1a7OL7PPe
BO/ctNGRTHlv1+b3mULIged6h38VuNWR5ygm8j1WzxPggnt3BoWABUIprXBz
nsLmPXm9rh1eJzBTxetRak4uRLUEUxaf4eTKUXia4qmMxVrI8k2IpRdkLVGc
iqEGyeqB7djhCjdJ/HLwMYrfPUtDbH5BaVqf8WwekMFKyiBqd53TTdAWOEoj
7dkeDNDPy1mrhf98o7n3RHmEeiMTA7xL28psdtoupQ0xQxYcjNbuDdYfleDI
NktU/3nHxayNUc9ojuLKLlylT+fUv/oQtUJzUP/DS+I+fFUu0C+ib0ZvrDMp
zTNaZR0nzLkrYhwTS7vEkkgA8ewlt3f8/N2nfJTC2wHUP5zOpeyLR2HQbq9B
wqOZqpNYJZIIZEHHA/wbJ9j/vvqLMjY1CmoKqZsc0MYholLMATLHChop0hx3
ov8b3QPFAQQIKW7XJC21k0yBGyWQGyda/k8ELKAgr+mfjtPuANuvEIjXvFFe
x9HIvDFAHWdVJtndpj2UDxsbjf6QkqH/yQM+LuVAY3LwNip4/p40XubdTJc5
ITGDz2jFC9Mk+YIpAcCVYqn9n7xDDsyq8dytIQ/b1shKojABjuIfMNFD0XN/
gVpaIS60ByneJzTLZrjMybDtWcolqxEwE1VISYRwv9VY6fC7IiFrRsQP4n3X
099N5Qsj7suFXIPBiGYISa/igy5niRY8mX16S7XsFRr8Jfu50GWUbH8vmXHB
UiY3xk9idQUAxckUBCdWZU4wJZFXezr+DcC+SUzDCFOq7yU4RVhsL8J7tUdC
bhnImhmxTIe1VSR9MFqdngPaOxczhfasL06PFfzUtlR8E+fpYcRKTMPzFrxv
tplGpdNQnP7KchSFIgPpkdXAQ5RSRNMl1ZAkjiI/1FQiOiIGoMYa0M0nSt7w
JC0ciOaA9473uUl9OUBbUqGl3K5+DGDfO9zAYL72WYK2RtXRptI42Q9fiXUn
MEtCTXVRcKWYXw2Yo5SrxBGWgjW03Uy77xq5G1GUjMMwmkMjCOhZj5ieuTg1
EVGNPpytB/GHvirvv97iYv9EzC8FAjiFH1E80+Lhxd9XTVYu0u/ZdAQCD/uX
7+OeOETvfYXY9rXSQfQloRB1u0MYrbP0lykXsm0A7ZokiJTQLBGIuF/+f2AO
rEx7sT/JNcPdVXCn1E3Kn2MX7eueztPnIJeu9nmq7YF0YGzr9/uaHU/hcAjh
a4DN11vltw9XnwiXOPZTpR/M9Iyt/wHrfdzZuL+1vl0ZDtIJq3kNUlaV9cER
rvhqLSOwjCgQVeuk2wn8pU5S2DCmKEh8oskGytzDC4GDn3XQnoGjNktiZtpn
S6I9yAeNoxeoJ+jbBYlgrHz0c7Kjl1zp9W6PFqnAGJIPWpZ6kJABBztJEL2K
gFJd5y0+b9Vi+x7S+qi+OFhk4ILQ6lqMspcwgsZuENOmLD8qyT5teVFvryqf
EnBP1VigNhGBiYP0NTP8h5ehL2lH/gmJfSPM3C6RPGEUi7kDw/91yG3EpQ6o
PxSL+kgq1mW0qltNpTrBT8gYvCFg7o3L9Qm6meJyIf4nFwXwmYqYU5zKLznu
mllEiG4xpd1Qf4gB458xc3yFcKIsmTDJlgiD+Y5Glov3AEoV3/F6D3nTRS2O
QQyDZ8YXmEwjZ23bQNFtRDq1HFo3AcEtz+wsqZRRZa4t4Bs8szNllD68OzwA
GfH7ZNYivau6znUEuS5LJzGUHboLmcAOo0QQJq2F0NVj8m8V73jfcvSrHxay
0x4IglmSkmQUOrgQmRjeTWwL7S4sLzF0qoL157CwRd5tH1MNWWXVJJCCRCl3
y375MGNN1CYRw/+yyZ1YbP1bVYOfEzSPa8sspWLO6rWyVl1XoJvso9KWdBKb
gkncQVWlhvOBOsKrXBw0aOzjglIzJA2MITdqtOF53AEAV/AtwqtGl6wYLu39
Yz4T1W4tzYfaGfkUNg3C2osPPiEz72FRVbeBlIch5wtnSTgUAFO/YVI+C1iY
IKeIWIZzEy7kiXAv8JokUbrOf/1n6RrJz9G0IT5Iayn87M/xd7aC2Sg7ORhS
e3hzpViyCwa9MQsIv0U4s1mTby68h8VNDqyJjJhLLPSuJE3Lbcnh/fUwhpIA
RobQqJC5GItYaHOpgQqcxyucyHPKqqF4cSlnOqhaww8opJevMt2jOgwl8ziX
vMdC3YaBk/uVVk0pihO0dv9DU6Q90L6Pdhjo8eRfFkVOavAufIIUVtvRUWg7
Q3ifIV5go7Bkh0sqOjNjweEnnifc10HpAWKk0+NSKMCRMVlt4aoEQzFADXvk
4OBsCLpMppJp9SPvPUAVrwf9tuqTTpe1PhOh81Ge+RfBDPw2JGRBouDM0SPE
Dlu3QzL16Lpq4P5x23z9RUrPEv1a+Uj+fQazX9kziOo5/adcDpk2tJHkuMvq
rJZZQv/zHPJij89OKEPtCXgPHkQsjWtOYxDBBFT6iZqejzxZ1sa4f1HcKv7M
wpAJtcgBoUisq1QOy74apADmuGK61Y5XxCSOkrZVpNU8MiFuCcsGOVgPnBT5
cjChQF30rAWd1h6ni+KVaB0c6/agPhtWYxL8nXCBSXoshr93Ov97TfWhfeBq
pCSjYZfVOZkhah8ouwjfZLQ9CmIJ/4Gj5eMaPgGzYI71tUaCLyYNwn9SsUgU
XJD5Ze02d0C7uFzdbPQ7lZ/lLEcBZLtv4hD+2sLOVwV5eWmQ0DNtdj6FDlGa
ceC+7sEKTHOca+SdgRb9MfgmFOFWfdi/54A1s4lbB0WJpHHqkmJLw89CGSuJ
6aj+CCqpVZtmtFfIuXhnlaTL+ECCUyD6/UlpsAAQS5lm4dhUy23NbpTLb5T+
nULFcn0ZIIUqWFRrfmJumISqxj2loCEZGkjIbWJw5tEiNkiS0MApU70IV8AF
mu3kLvabXdBenjJh7l2xSR0bsroEv2IOpiMTwLWwTPP5Z29K7dmTmOLeznEW
8gUmPUQlaxMUTyD6bgrydLtgX5/HOdDA0MB1l1dNIkMdXafcBO6NOXz0yvf4
1LXnHmcCLvBrzSYQwfRWknfPQS/h6J2d0iFOKFK4FPuVXOMJvzXtAkQAjXTg
zsjn7ndiAbq/JlTNyegj7xOQkyJV+q+MuMIq26wk6IPvqNI5eZEIVCCr7mZ4
Xuai95kXSaQk9Dx/fGICN3zxVkNYbmiObdDEHv7m25Ub1/c66MyNmHAq15f3
pBpCK4dWfH+CR7K7NvJqKgaNhUrlRmMma1UF+ZA0/f49djYpruFpGs9vsUZH
xvwqsjxj3naO7I7K1xBlOzsybkhnsRa1w+dLASgMA1JcQ6/BgJtaw2Ic1k6+
YQ6MP1TT3OPuVsgbKfJx/E3jwXgNz7NU+9asvfsbiE0jCASwNzNv3hQbucnl
OD7Nz+M2kGd1v4Kh/9XimZBkk2Gev2jHkKCtlSlZnUjOBBMSePyJlJgIsgVe
QWC4QU0teOqrn+OIOCS21PQmVL+ij8t/4He3WiKmOxAB358X/UEIEPEaCv2S
8nWd4iJQX7023h02oXMTTE08KnZA6Z/77uL0/A+cFsHNE5x+JPRzoUPT4J8F
8UAmAOKN7MIRDOQzMTn7+7V3sdoIWEPD7h8+UQxiAj74hCgernrJnLOr7Hrw
kSk6LhzqEgbpKwoaw1fKRfbnazSHzrTQKRP2iSv8FDa4FdJ5GDFE4JdFWx3C
3CkBF0GKWnBdwGcyN7GSYn4inYU4Sc9qFRzineOX9n//I3UcmpSv7k2xwZu2
mUe1JX7P8G6n1GWrJTVl66oeUbYZZvciG8EqrX81lrj1b8x1RuaqQvsaiyLw
/94H7h3O+QWZl0ysZ2Gx5xKWfdZk3jodmvnnlWwEfKIfdaJ8eswZj3Tj/UmJ
MDaOebGUO25M2vjXgtImjPwUCOmmzOBzLvKIODtxQcaHG+ErT3eNBSMV3Hne
oVTRRItx3KebrZCR6ak7aV5ES+Tc+zCeRr71IDUa/gANFTpn4B1pdaG7Dw81
6eS3XJA/ZSiED5rfXZviFEG3rk8c0U4ySS3AvykrwWEYZHUbQu2YLXCVZm3Y
0aLfRmUWVJSaZal5HhvSCi05Wd7ChQ63jsvB3xvkybXXLIGR1pfLB9YabPAG
GLPwF14Oa9KUN+atqDa6bG6a+8U5QIqBA3l0dVhX5xdR4Y5xxR7wsjdANVV/
6y7DkuEeY/rGKaU99nOpz/AeRDoCAcL/hQvwkRtx0Xe8yCR1KwEnPGRZoBkL
6hY5TSEI1qIsBk5P2aKxO/u07Vufm4+L2lbYYygLU0WgY/VDLc62gqx1NyeL
MgffQNPfbH+77tSAeixzs5w+10HYH865Rw+mwQ1DFLEZUXkFPNKAZB0KJtrt
ZoKJz8UkzJR9hv2j6z0xy11jvDLcSDNcZc8Tv9kteolyf92+pQpunzRfvyEq
2VBeaTGRbzUlOe1/sAHBCWNfPv9fFdRmEosspAJhaKhwD6PDQfLY/n06p3kh
yWndlOBhJwvfm22rGEPMnAZQx9u+vkFfzfgO2OxY2dpgSzieHE+jydzWCBB4
114hkVj4sJiMCCvUDo4CM67sNpTJw5CXzORZu+nHTJ1jRLllQrMPnn3N/5q9
YHTZGDzisYfhi2apDLjQ2A7P3obza3wVLnf4DtdjrDuP8j4Oqe1i2aITcpuX
uA2dSOgcHdpY3kz7livIvNRzOYsbYfSAQgW26Ugw30xT2ptSXkeGl0W+WtBg
4Z+Ehu/Q9mQP2S6cjWKwB6XVDt5lZQJae7N8v41kbM5mBtfEMs/S9/eX6/eQ
JqKKu5reg6MPn25xdaZOiH5FFmHxmb1CSvlVeX6bANwQoiOlev3531LAZfOU
xE5n/ZWgrGf7I68x7OmGvrw5gTmlHXMXVsorQTZv61xlzD2/ktEzODJVCMm8
LDECi8bCrUM0V78KCYQToyaqWhQvTNz03jinIqqTKZB+T0S4N7CmF8Flicm9
/BEt5vILm6A+tAWxcyyE2G3hfyatQXae7xCCAIhLM9I+bMkHctN7G6EwZkGX
1VLTMuk8sM0Rl2ol5hhGfuDKmaKPj1aYOEr2OlWwgMl8Kil9NDprxzA4vLuX
DVslpJYDQLOSPLBfcRLD0SmO43MeIyrHvMhsjwIApFHCfz6v6BOcDgDaVZj6
o2vMNOXYMPTe9dsIDj8e+VGvcO6IR74sBZI/vWZ83xaEy5gGoD/sZwe0vXdK
nAcWnYYG9Nc883iIRdjHRZYuhGh5mRgT5NhnVfzs95qCKlcNwCUMrgTybJpW
VZk4pkrJi2IXOYko3tONlCxfgfG+5q5LOQeDkxyAr3mzEqK5bQmBw8p7jiQd
I/ZEPPuybfW04G6kqdez6z6T1fMHv0cL6E2aN0/AskfJZI53gZlyQqPSZNxE
eaac0K7Ol3/GsJBUm3DkUSnJW963QhtNcsKjIV7wkeUDumHcMOEzXaT0dcD6
YQu1e8bmSoOOUTvdh90YjsnmDYDMOOMscjCn46iuLYt14MWIMNxaPbdoNGZy
UV1tBJ+EtPTFrlQikG2ocZQADAnhjBsv6w+JzMrAh5aS87/BxWwD+sl4nWFO
z0ByLSxxLaZ7Gnvy3yG0dccNTgkdDx2erFGX0T+izOvZXeFVoCiw99S2X4Us
jH9bmO/hbTsPIrTjCvA4oYVpNefZ2e1WPDK7IVgKAIBKxtIfjeK2hvzaDkaI
HyLVkaQcgBz6r3eDdysWGvX1DndCONAvF7P3V3VXu2cRYqUK+naMt2/CRQ9q
otHfhMVCkJOHT9vUxDoXN4zHYQPTjnTz+tbvQPrc19yZBjT2xCOPKgTjT/TF
BeCuhaVkromhu3n9SDNBcAX4yRiUPRVtuvT0HDsFAxkuhctdo8Ru50IT5jgE
+O2gF7iiMbQvAubLAaJCVbq97/iW2+LcJvdZplT9L7LRgZ31n06ZBBB+UcOP
g7sFfy7ud0UTrugHk39FXbSXwRuPZhs8SWl4pOnP/f4sAfv118x95kG6W3bs
Azv0v+mAOzuia5q1Pg9ZGkd2DayCyKEqUNbZDAf3fWSKYwl8qQCXyyqSi4AZ
rIuzeJ+ehKkYuh++BHKTWkNz1Xt7kQm5R76jGFFzgO98nql1F8Ltgsv7sFi/
ljA8e6a9qUWOZIUEJQItms4cIlAs608i/h+JSTfW+6u2MydOKi5P0k6zTNXa
/CcmpTJAsimOW5YM1LeK+L0HQQPio6yAD41KMdIkAFFqZHQIN8C5xdGLsCZj
eb0JHwndf/zPfk6XpE8O2U1tG+y7b/JJNgl8yaBmOUi2B3TMrB9M8GteHGxQ
g2biB0vghmKMtxBBGk8v5IQFxUBLstsBvnY+9t8y31fXy3oIValBFKNDPYcC
HBF5WU0O6AdaxvJYy8VzbvGKW0BhhK1APEnyQrTXE2uRVKmIpLLu7i5us78Q
Tl0tv0WhAobifoqyp4I1EdpgPW1pIs/3k0LjvIc8DToX0rvOKmSWrF8ASUsV
3wLzkqGE6PtxUYwM+HurM9x+lL3Kq6KLV1TOA+tpb/ZFQ0jAoM4Oy0eOzyvm
zh7klbtOkgGumm9/Byk3DD3NVPl0Plj5ZiPW9/+W0EFD8W1LuQyy5820SW5s
WIOqeT0uRmJ7mt+vXv4Nm8LBm8ZV+cYeUdrSam6A4socbE18tO/jzyvYwGEB
SeQrts7Vf/sHiyzgb6rDlV6hTjYGAsDzs8kyzMYo8rwmCV5yn0bIL2ZI0bxX
HLhDE05HseomJd3ctBCsfqeEl7E2JKDGoo4JRPkQUfO4tBxxWrhWlJ+6wopX
V6T5XhpbZ6R17FV2D2tqaRZh0whRZWA1XPotWMbxgayNB3WoodxGqf/IOksv
tpmsjI+ZZeS1/TBP9wTP9MHTqe2TsYqsYtncsnusYhhcKWpR9DCH57snB0yO
D9hxEF5DMFN17JcfvNsJOPmuDxCbczSZNI7rPkIXdL0UzXeBtwHFEuOs+kUO
8MgcJAHCVMwAbcMjyoD/bQiVINcOqwuKrUSt8TtdZbdyolqcJ2VVPT2Mi9lZ
3v3gCwqib1jzPghxOBtkSX3pFV4T0VJBTWamY6TBlpkdP7B6irLO75icrFzP
U6YaFg5qMLcSvlUC5DGQWHaDudlRqXoDIjKMO1uCrgH2CTuFjuVPx+jV/5xG
XuhPJVj2AEqg88eWvxzgzVncOp4Pym8dfedpJTKbXe40Jw0PzylsdVx6x9oA
mCxzMfn9kRUw/1jcrwBIVa/9NYNaMt4yABXR2HCPiq4rNUshrQABIwcdkaNF
pLSC5PaxWaulGCXR8zWoXaTseRLGD+3b57R1Ea7BhEHipDWst/Mni+O8qUXY
6APAsxc3Rktmba7Z7xwhWDgxQQpd2a0duvwmmc6hPiXp9VeXhNTrNNGh/UPO
9LfYgP4JgediIr/40FEAo4w881mcFOCE+CP6KeA51JlUfeLOCaq+R/BZbT25
vQuKe6If6Xk5bYBMjhkdA4TIo/fjnTye5kRdJMBlQaVA8NY3HNXx6Ang/j21
Ax+ArQT+rug9unt6I/71Eh9EaGOsp8m2N+KkpR8ggUoXgpntQICUBNgr55P1
iJDFl+O5UbhShNg7kHWPyBM72vZSDHYT85QV142YYOZiT4yQ6uC5/83F+cO4
wjwGjp+LHAFHVQFq0+e4toZW2MlyKk8j3G4WKmE/0c87idw4iuJbgoaCVugv
K7o38Jna0QgiK734zRND5Z1KrikHdB1luH/fgWjqdLiO+6cr5BVN2m5BF53D
Y4o6gyzjqWv3RzVn5lwsFZQGLv2JlR7jqqNSoeOaaxZsl4NgQKxJ9b/5E9Zc
q+D8GuqAqkArbYi/UcNtOAzOrHcaMdsI3HpU8ZrnsbPfkBySgeTBLR3JD23K
AfJfWuUg8zCJNB85V+y+4kCLH5epz08XNYCiewDLOg9pCl8uXWUCfOooB3x6
gKox4ttEyjlYw4U4XcMnQOhEEAJUYEEAplc86a6cCVCeIJZg23lp4m8Tq7wS
gvEy9Wq8+WuM+s0Ylkeem7Z0qSAtzWgEotS8JRpu63kyKt89oQm39Y9v+inA
YeZmhD2RRH1C902o/GgX5hZADcnx2M7/ZhW/mC1Eb3+WtLihqbIPDYEOikZf
8BQATruJt1TZfBpeLWBxiLnIITU1526E7H9lslSE4oMINguV5KLMKzhUc/Da
nvknSEQf402RMqSMlukHZ/ganCtu1zkE5OmduGuYh+dhK5xOw3L2K2jYbvWK
xEs/E4Q97tR6IKrdSPhml3weToNCrw+K6S+zHMRDNZ3Q02XFZkHY6ImQVJ63
66YkRt1DD8Wl/5fuW+hn37mYnL2OGjQs5MnMDXpzG8gVdkK9Ei4vjKLonIuB
xBdpBDMNELm+irQd1f0kYnrNpyEdEud6b9esOQQOQYLV7HX6t89tn/H6CxXK
J9o9UXWwibVeTHe9eAGnxVxqfwHCQFcG0OPZUIbIHckJWygijW5/PLlsRgAC
suOHf+zjtS6kh/X2bVL4Enr9OfSRXRZcYDRcJnlBbGSRI3PqiZfqTzBe8JUZ
qjWhcq8F3Sg/2t0/isLQkfJdy8JiL9rYmWOg79yeijVJ/0rmhqGd8WJwjCkF
URip0UQ9qMKdUQz2HZqWS6VGGXH7/i3uvNKno5TbZ9XEUVolqFM5orf+YMMM
NQNJN/KZe0v9LHnnoA7jGXxDwgwylNJhnzIq+DvWQF8vIVSoK+fzezbQ1fq+
3e9qEK8OhVVGr8Ue2v5Tll4xDZn0c2IRUgraSfnRY8Aa7MY6k/QkfAuGpOlN
FtpYO/z4ukcUO1LFgObzqvHUloIOfIjGqJLvVek1s4HFVBj1mCQQeqAPINvG
AiQI3tJlKDCUrlAkdrhpxuTZZJjTOW3tU0Rzkdj2HEfx3pkv9xvtkP6F35FD
Ax/Iv88uYl2A1F6Xb+Ev+6N3Z8Alm/GaWxkXV6iHqESwySE+m8TKe4rCJOOB
yImxDHpjXMzmrGX8QH/z8Aq3jRTxR3EpdAXSfkq+pn7Yu3n4FsC0++i5JnkM
kqc3V4Yvet3u2Vz5oTHFalT7AAyEWZGVrfKErho9cyEDQyXJwUYJ8pQLkNLp
4DZKrXbLnDWSNlJLy5eRubOq0ebypIJurLJw9lPKfgJzGXwP5LtyuzWoLErb
SjdebBMGnltYfg/0H96wTr6vAgMVk7qa07/+X80ckwkLiCR4sxHOWpVRciDX
4qXX4kcH1emEmZmAdCEFChBU/EfQhZ6xid+329HFE/bhoE6yM9b7pT/zqtm0
5oc1wIWLSm7S32UyRcIUnhMwabXppewej5gYQrnlyLvBf/zy0t6fbMUj20lB
fg2ZkwRWMyyUNtVGI4cG/0FsJDe85xQyOBTYG6NcP0LvPqrVpIwhyFLlhH2T
UnyLxuhnjXAcVRyezsK9PmTkLaqOwGZM9nfmM7eceNGl2t+sFK15vAsmqRNT
aoNExHZSWxSWciGkclaQw4pHiJNdINgKHy1vnUnIIYCPAtJYNs9dC9cMFdS5
dCw00/MICoezuyqezwROAMEtEthT053j2Wb+uIBdAezpPGJvkSs6bAMulxO1
G9fFinP56VVKh2eiyN1rwCyHoXSMroWD9zngTBAOGQ4+2dSNFFnvzHi9J0Yl
C/rz+vhdwEhLkLur9IgWgvQjlIx82xiDuULMK0Bz0/++qb/YT/zn8afojOf4
pNPN7V8w77ekMyYjA7YCtdMtymopLLDqMUz1PHFbhpxlACRLdLYcLtK4miKD
sXeBWMf6CUjjkmpCMt2CdCOB715PW7BArl3RbETNHxRyD3sPPj6bZf4FLmLx
mg7ZpXdmJHRvqsCi61P7rrTKbezfLtfiDDLTNM9Wx8ff7ROEhkfziEtT8/Na
OpqPIse6hx6NtjxF0nkTSSziFHktYFYVewFldk7ar3XSxYK4xnJlmjAWYiaK
0QvBSqzD07Vsnzieap8AnWaV/5ETtmkSmQTtMz3gXXPRaonc8aCm95ofdy2E
wpdAA8gCqeoGGHaDGiAvA0IYqJ3m+R3Wo78YGBbm0/Bq3tkNIdU7QhDlSTnt
ynrMbHv86zjYmjqbuCfyyd2jbYOgf+Kqvb8qQafGU7MC9MqsUbY/TPKu2BpI
oZm8Dnjwi49lSpFDRf3AzA1ZSQEvDEibDi5yjnuUdQWlTarq5WKevMHrAfb9
maK1LkDhKXx/+HDxZNuOtPYyJlGjqGkt8mUipgN49+a7c0IC6xNbkgPKc1U8
VaA7+b0L2+s0m93WVqmjT9wEYhkfRZl7iGf6XDuljv7H2uMKyvavPhEWLNDY
esxpU3ofVyuCv8nFcoGSMzPhfom1IViNiV3+5KU3pTZ1P5A8pVjXigLxbiMg
1fC0gwgS/N3lLhi4pkWBiOjFqSGcencFJw+GZN6hfbYAGfrzpir+et2bSKVe
PbAJiP3/LbHRMtSrKnibUFu4S/sX8i9R+GzFKKvTD9/LqD6NJn7Anq95NJYA
THtP6Po/SIizTmDe1boyUm5Gszfx9KsSJ3XJJIwkTWEu2Yys8QbfiCV1G2oD
s//Fu83GJpnjGvH8kIeN2m5dBp8Ii3CzMdJIKXrysBAwxLHQQbuIpS0YMsi9
DMmI/mV7cOUJwzO31d4/no6jNMhitJ/RHQAd5V+MieOAoqPIVl8cBCIZTKBg
vxsCpkNk4ESl0v6s6k8FA4tLEj/eLXyv3wUx2TdjE/L9S9Po2sMyq1SEdc3f
ruNxgDWtLWxyYCHGzudzrUuSp3z93Ab20nXTuEZI4EDnVpSUHWYtIQ89EMzX
vH9U3Kck2ZX1KChyy9aPW6y4tVjU2R7mNhrOsBva8DSoC2pyKnugcM5HAa6d
eo78uKjSOTosPdtlwlvrD45jcSAz0QZDORoDXW3/jthyxTE0/fj3UeVIBpOj
h25T+3jbrs5iaSTzPD9coB5KnfM+J9KvNKBMtWg8Wp80ePl/sypqm4UVC2+U
hjcmjWIrnuoh23AsVuusVC8yrLFMe8FfyGWdqwzc0637T4fJeE2ZnKOAF8ro
ZnkiOEH2GZu2z3ct5RqMCa0i+i37AMBOEqx7DJNHl8VecivkrXKwGJULtiJU
nyp8pLu3o2ocZGUdcjzVSScfNxmhyp/yFU5Br9Ta12OWKx7UNa0TNUn0hGMz
5+LI3W2z4hNFOOfmXd/55g6wGyn24HPHaog+10dOcoXkclzapHsgqAjUwDcp
7Ix6GrTEI4wbUrxilt0CsknQ7W2Vt1Qf/zAORu6ynqKlfA+mgUXQQcr4C0N0
eDiWUuA9v2+DmC9QnOYilhoUjyEa5fQrP+ER1MGZWpDGRH1j+ccrUtXY1y+J
CjCqQa3Zm3MTPoDweLa6/bhtuzth/t+3Y+VDuFMRp7T4O273tyPH95xxBg2v
J2m0Z1aao8OgMo8Au+RPS9582X598q7tjopyMVjJoVRWK9uWlubUqp6r61Cy
3rVIOfmA/ji3tZWC29ik945dIhGva24/0hG/hBUIRXBXfw0S82xSfiCtLAKY
8kpQNv5ub9fggdsUU9lfyFLcUb8Sqht47KMxxHjqJ77IFGwGxhSR67tpLOOM
OQ91wqyKzUT/oAE15seXePxSr0XxZWUEjWsF4025DTRAfHYOVsRa0fleHEQ8
p9lfhXWQD4vLJ6X71sqQ7jvUMJB9sGvL1zSMkoKZ/oIjmpWZ3uYJa3t82TjP
mkqSkezkIObRIiPEaxDUxQ173vQrvs9JKlI5844tqEO/gjyAHKs/Qu9mFTYE
i8VkhYU1IHQ4coTVTSs8jOBzhwtGhksCollh2c6zq3bCf3rzW8ZYlTbKCIXB
O8UlIuA49PYz+3gfpa5XoCnW7UK2FHGN3G+kEfT9mNenDvEhLeghZAFhBeoW
8ajNghpAW8KnM9+b6OVpstxmf/aeBn43YdX1M4SMKDaD4vIOSltX/swkM5H4
VrxCntYOcOd8KpGEuQjHIKFCFMbBkCXfhtlVlxSssiYP9hCyPU4ytHvWpfeX
I/vR+/CfmpGJjXNSJ76AzkiMD3ExThUdXDMRbOjd1O6urlqlefGZiWpdr2oe
czkRo1c1UN4htAaDYWsq/s8c1hPfZhkg0dPDHCXRkU8zaCFygZ1/NJW2R1bU
MYQuX/fiUstQDVLNsj6d5L38ioIVbSNpmMaCnuwJpT4s/9XpGJvImK1aRKs5
aBCAyzZY7QtkXMaF0bJxQ6xcrsKWDlTe3IDpkK9JD8Tpc/tQ4SJOB5sKp421
ANfvS21O5jjByGw2kZXTvGOdVKQ9uLn3x9bN4/K4TYzh+K+kSyDyIGlg8Vnl
kK4Xf361w8+YF32OGRyXovxT/wy4yWfRNNWQpxhICIkzyufrJUloZoAJSG/s
OMJf2Klz9GKkP+Ee3ikC9Yv8r0hq+VQjs9hfAVomwYbJgEh3WfEbvKkvGKBx
Ql+kLB7x1fHf4/TYv5JqLvuG+S5Zmyp5zU8HVaK9qqgrn5TII2tXevJjeju4
Dd1LIDDI5VOTLuPVGe5NDiIP08l6s6BJKL4/wg8US1+Xgu28h9By0/+50KPZ
Llu0gNVoyY0Y2BaQHmMw/OF+Guynj8mE81rfO3ImoNqicRNZ9x6dnCDTeji+
mN97o4SKMVInQNE7zFg8FvVkJBElrYLPsirPb9O66xjXxQu395J8Kpyxgik3
dLOhLOjcuCJko+yhQavGURZkvD8hf9pYbU3EOgnTSqFngD3HGoiYuCaqkms0
tq610COWMs/6QRgJsJQYwx0+/XojWyC4z6Da/opoa1xJYhpQCDDeu/SZoNeh
y8Yv/N+BGWJYCKKk9iu6Itk2oGnPZFJ13hZ7K54Y/0FDGkbDLnANHknz9qYg
z7iuGH82wiKCj68WljXoqv8b4bDLsMMW1wdgp+KH4atzFmtcptSNy4XOj1T4
f51iZFMtAgWTCQaJYfhKgsOmBqcQsFNvfWnA82vgqWJFCVtTdvXzXVK51v1z
gUBkxasPW3xb5dK8Q8bHX17haPozum8vFV1HEvkBFo9zeTzGgq9jnv6fcgj5
4dgsaQfCB81ky9IYUFhU45xiZM/wpMTyOqk7nIT0l8Ko5wi4zLXI7lu30VhT
H9orq7lDN8bbNIIuPx5x/3Y0YJw/iu20iCEBQwT+UDeIVIeWkw++39EFtEx7
I89Cm2QD5zQDZJfvuX+/LS+/c6UzKGWWHvpB7GuyePdhm51dPM0qN05JQWEN
tp08yNq0l2VXk37tgFsb8EBkeIrCtkzLjE+mdjUdou/51TxJsR6qCjNQMpp8
dBPToyk8lo01DVkASnhGEqTP8TM72UxXYpGKEguzYa9irmmRyva5Ed+BySG1
XlBmxLLHNKokhgvb708cLosZCPp636HGQ1ErrSb+pvbwBlN7sRDsB7DMygwk
4IOi5ZM0Y2bpJvLdZhYnBW3V2jLgcnPNKr9ogDGT60KL25ZRQ/K4ov5rmT55
4Scsij30QmSuFBGaATCvXyqseN9C5OqTjQNO/lSplU2Al1gOh2SNAS5KlPgO
pqMry4jqttmPue8K5lxRZF5CpWnLK86AljOYV70n9hpW9HsnfWqrPz136wrk
CG+IlRE/BB6duz/0IG6I7eI1h2UN/D17rQ94JSCqFIYwkmnI+6s0oUrO1lZc
sXj/JTwYLtCPgf4kA+AAR+R3OFMFF1V74fCtIX1S4yv4vIbyTZz2TB/f6CBT
8JwhO4LnshKMxxhKjJLCPAe9h89KbCBy39khGRV6h/EYLLLnyjH6qoSpU+Is
4COWzYLq3MWh4VCHzI0vYBtCaLx0fHEwMkUZM7iIVZQ9wu/InkCgBATt52S2
KiaHoRG8IJreM1cZ2ZKPyBJF3Ng8kPXNjLyZRV/KXay9g0S+4+A5AlIgitKE
Oji8ZdNMs2f/U1/Xfh7o4EF1LtwVdNPVKfoD2zFcoCHqmnW98ryRFPYeJ18G
WcZ+hjtErLOPWHuIIVrwC3Z3HCuVBbEeLU/w6lOf+P3Lq/cPbYrFsMLbUoh5
UQi047JNMrpZU6oMYNdmfZKjn5Zx7w3SVFsk+Vp1wSMX+R5HFG9EQlI03uzL
R2eBChBio6fxdnyY0fwAxLaK9gf3CdHVtsjOGyne1uhQqyD6VeppcFwKg+gt
SQWGtPZx1fALTqXeQwsdh3immZdsEOaX9E75mDmIntQ2hdXL9Ymj+M7eXxAl
wVfkQ82+XliEf50kGuGbB6gJ3Stu/JouCwC3CpM78B8nnYysz3WY8kGQix0a
b3KiDsqTP/DghhW60qVCRhsfwtf6NhKAta1NovPdRcz1murHJe0p/MB28aeJ
8cPF/zKjjcJKY6fC2RU5MNxBSOJls17bnxNII4KcY/S00DWxGi7LT43wwV6d
zRGKPFxKr8cqMhZX0peyMPx+IZ2tG2/JrctKeTqaL+At+9F+eRcIoBvGNk0G
WSTK7350ZSQlIK9pQdfiUijB1fpF2UJfGElrlcjbhFb587hVHQEFtMB+i0sR
SjH+Y7p/4pb26pUgeESZjsuGO9SKLwQE6At4Q1heo9BhRZY4m6g/8uA0pgBL
mG7kEMZmrlTwAGA7GpIu+jLUOHovJN+1NUZ/yBuiGtYd4PRNhEZlMiskNdxw
PBzo329XwAQ51ILmt3BUT94kUblc69TvRnzKaX9B86goXuhi3dMC525HWAT+
BzULQN8SzxoAhoHt2TyBJ4ajSiBqZHpjihs2AbWDl9eibrqtp0Gfdc5jGkzu
VAy0iDhEtngYjrMWqbUdzPclVyjF1dJFLLfkGLLUwAJBY0vFIwFiTu775Jtd
I+M87whcPbhQzIqq4Vva4R7ESrDV1gChdCslPSz1VkFRlPcYnBRCyAM8ttZc
udM1bTOh+g630RkRH3gW7j5ka6Mwk3Q5raY2xK5/FoO1UksFfmtev88E4z6i
QbjqBjNjkTiQkbvrmpI2Rk25qDqjQFVmwgLLOJyr6y0oziK270v6MyOmHd49
st77Pvbom711lXobavBlZunBsf1B3p3q+rR+Nbja3sL6sh4VmQrj390uljY5
1ysMzOT/GBodKEg1kZlAJRk7Jz6QwQqpGDCocMLH+xy387XREs4YXPjYjwXS
mCHfOuHF/SLoHnpY8FLf1CMo8Rg1S+tYztSHnONlzNJoXyCQWApFZm0ido4p
TcTP6afmRE3Wdpqf4WBNd9b8n1pBnhg33e36qVEAP3/FL9120VoA/4YqcrxE
H/zUt3jW2+1ypMSWkebR9Kf0Rb5HMF8tzLFgWrs5amsM7kKOKje6WgTWPZSP
zlrAPXucHj2WquSdxBGhhUu6WzI7xKOZR9y7ay7NsqoezlEqTMZPDSEYHInd
uTF1+BkUk+Mwqi1cynU5x2Z6sKkXnPz9iIrkj4vYHHhOQ+680wSRiS3oqUMn
4Duz+t+icVLhaz9V7coOAlstcmeZYIV7Qz24Gu775WwGEbaSOg6tdz5pN2B0
5iAeE/n0CFhe5Y1MFjfCBzZ2sKgjzi0gZWWqmPR7XYfeQwAa2NC4H9kqlMOS
WSc/60mtSXsY4fUm2uzemeMqZDaSQseTQwWobJnW4kOL/rFTmj6QRXYuypKt
4H6Ts9F6eo52tPWWeAZGp3jG2qrFFsClBORY1xYZwInvisaVWUE3/y6IwIi+
SkX85ikB8n35TQ3sMvqJubie+H1fUFwhb7jCdzfWY3AA92pv1uPZmZOVE3GD
zyINM1KXxF8NblGMFCRzXVryAY81AuIGqlhT1InMLuVrIA6d+xtFLdsTYvAS
N92q9g2SCYCVs3oawnCExO3V6/6VU6cT1JheOGkvk1LXvdGxul4OOzLcF9EJ
OynZc3FUPxLkEHhu6PQWDHnuLtfqce448RQb3u8/HlglV20ONbyhcxz8hlR1
OcDSkMMwYiKA+iOlUICOYgvdtZo0Y/EjAogUPQG1cOiY0kjixf2g2NrlaU6v
mJNiLhpHLn9HiEQxe1PajwivXw/5FJXkFuHo+UI6nnzNLDiri9IKVFoYRsmy
F3lAOuwePJRDzvb6720Xwkp+gG7djiaWMaSVejxc+H71EVNK/6oz3q1SCCQ2
WY0y1eviiz/5zPGWq/8hgsbw4mu+ZjFemWntU1wDTd5tGQ72vp+/mq8RQ6Jt
fhLa9UPLQkf4J4ziaDRHIp/itDd9S98oNJGOA+J/32mWkUiSb9uc7CTbvUCB
OsWcFRl+DBGxbCscckNUoqWXd0lYIJdXpCGTzFHKY64wvGIpl4K0ll+aPChJ
4UsFGccYQiHX2o5/v1OQiokoXWniFbN4wCoZPkHFCYmqjza8zn7mFgyjL6h9
nZhKmmx6zi6V5A/R7hqNlzmoDpDdPKE6LiLu6Gn4RO0g6RfckaIhu0+gdCdd
FjNWAhFDfE06Ha9j93srtbjkrTsmhLwiYsWP52iUd+tgKdaMUUuQMCDvJeX5
P3BxE0vJ96E1oPBNIBwHvGHWfXN1BINF+nsBd5ehrb539CnqqdRfqjX7Fxb/
5uA64+gZDGRWAVWwrX+HAo0xMq8AqJRDhnSMUfrVs7DY2X5l7vSBAL99jQMY
u5zLcv7Qz//+u/QO/WB6XoE3M2ZYNsRwwF6yKAXLxhB7DcZDepw7J2GrQQtx
nG4wjT3kOPlxCGWJBKhT7LTNwCy9Wn5vAzOy7P5INZiq57BgHpoaFVifHo+a
K03oq6uQycmy7rjV3b/pV+IKXILZRriiQeAmnW0o0hsVdvMq72um9nwbUwes
+tRK/tqfj5BCIdBv+9RqNuKuAFWvD6Xcm5tkAWcXfXI5i79T4KX0lQ2LXL0I
XLA+mNqB6UcY1nxr05JSeONBA/6OkBYedZ7ZoLQ8I03NNJ6F1/yJQjP+WHy+
2zzb/fMR5N13eiHQL2E3WEwKKVE2qnORF6jGlJCKlHDjtCh6sITERJ7TbVVY
TPluaUjaea2wPny0A7LQ23mhgC03iItaV4wgcv1b8tVHYdM9Lrz7aqzKuEFV
FI4nzkRjAgiQ92LoMD+75efDN1CjQJEDEPDsH3AX0yT6n+uSmje3kJcXptw4
FV4rr2kR8ijSwV4IOg2wAwTlvzPvcmo3bjnBCbxmx3phVeGoxl5WUqG7HqB2
VJ9crJxxFu9rGcVuTXqRaGpSgThMv0zwfCBaTJNMWLawyqucy2yumTitTJx8
jeqPxUDHNvoGGsrkl7Zs63/o7BxwfISgN2qn9OeZqeXndH6FVz+7VXbohiRG
pAYEjjzAGpMzTQOZPgRHquLUpon6BJE2fbBT8Gi4MfQeC211wovYo+EJPczB
B3jM++KLKH+MlQ8v2IlOyEgkZEwkyhOsdZ2wNLcUIGIsjJJwr6ioNS4yglZ3
sok6bo5G1J+Pnath1//xn5FgaQ7Sag1Ca3gx3XFj6Dwj+bdEpIreBAFT+WbO
DfKKqxKIg8+CM2XceAyfdcBc0rg4xA1a5XSaOSFZgqLHX6hHuXyOaj0haL1n
+uXoQKfL7c1nDLyMHlk4HcADvoj218EHPop+rk5ALqMwTkwio8u8RJayEvx3
OKzk/dQBwbtmGPtXM6VY1ywC42d+do6HcLXfIUwyEXv4nNxHR6OOOaWwSFbm
MnrO7f9JVhmDryfWm4nG8i1ZJUUr7GOHchz4cl7ZTMGW7zUR5Bgc1MnDJJMH
suD9EkQkhnM7DzcrP3xU4Yue54BCKe3NKPA4KHM6scS0IZyMgjnUUbmnmlsT
aEJQFvfeSpK3P3gX6wm3Op4KDBi2MeBy8WkzbZ3b1+18JzJ5LJH4qU8HV0Ll
yWcLh8Ov2eUb9UYbBmbNJxeGQ/mhnWhFwQjsQasv2yZPQx8cCVM1HrfZIOQv
I1w+AWrdl7JtOOkS6aks1kB/6Kp2dlEkh8PFQZG4Jx4Zj/s5BePSMNz89yRo
0OOe/AhpTA6Klte8V3DqHEI0Hbs1RksaOHlwAw4aeJTLRoB8OhaxLh+AKXyC
9MfCfOdx5zo7etpN/V2m9aeg90ulJc5RFpYPlYHzp9eMmswIDoktM2hU3Yjs
XpB3ms8irsNb4hiny3SVsx107fx5cj3TARdPu+CR87vaHp+lyIS7w93cDPkI
bx/Ge4OMO1Zj460Vv7d72mPBmtggB6nh8QiYizZlrvbC332eB7lFKxemkjqK
LDHK4YPcQF1/A3l8b2WXmsDKkjrHs59uA7E7hLkB3BAiQOQDMjYM3dEMjzFY
yf8zNJmhU5penm3204H7po3nDNLqpZ6z/AL9d2aR9Nrc/M3XxMeUCPUSu0ui
SqaTDhPLNdeUJlo3ds6r823YTgY2U7aLXFjZpmQGozjTitjARsW8/7vqh5Wm
tfHQT1VODi/faDXMPv7ujyPk9BDCDYqk+lWMvx8zF83BLTEZKzdBvPmv7BnA
IWc+87mMcEUNltqavqWOiyELWzkQtau1+RCoCmHCf/Ux/fzJSeMSNpxT9MBO
ATMltL+htQ7UToOAkZUcCZF7dQiVT9gauDRr2qD//DIIytPK0wCWwPXXQ6gS
mrBhNBQLJVtAiNCi1TSfoXIfsPfUnTRtpFVI5TpC9JIUhxBmYYCRo4+9ni/3
uqYenzbTarmnSrNsgPrbDvqW6wD0bJ7TRKJMfqeBMsCe2wMjx5LhJEkmsLcL
RGv4wBctoFDcwXNO02kZMQZz5uVxIIktvXt2kvAtvScpV62Lmnu7RndfYCFf
aTopNhWTCEOf/0DdkPqp/QjGsKl5vUhM2NYdawfnaBaOYljrSA+rrb+4jsJW
ZZEuxlPcPRentOnh5uCcO538ZBOY9QM4hbPoXXqhx6bRI+NMnFiAWGOb4KIf
SSWZtnitBY0OTB2FMaEzzL4+EF4JpZIVelJLfCR+otlPYa+dfxvz9xWoawhB
006/TfgtjbvQOemcS2OzmXhWqcL0Cnh3aUCdgE7SPjNQAdW5JH+vTQ7mT41G
UVUmC8LXePqeuU9Fo64LU2Va8qsxP8BUmMl0NFHylSXMnQ0zfWSlSIJhHckt
0Cqmvu5qUJkimtlzm/YoJDa/1pw6DqUFJusML+FoolVny1XrGxZNXji98DcC
uJcK/BaOIMCdxAPDYD69dueuByk/ac4rAUZ7ESKpWpVxBaqESONMoa8Dn5De
Dg7ccr9Q7NgnmtwzbObEWElGRIhheQkOLkdusYdazdbzwnyZ3gXU681k/inG
TCMsO/nSpVXdESivok5UkpCAONOXut5PISZ6sqiO+NEnWfN0irEh/cJ8eTh8
S5RFUbR2ku2sUjej1Yr4MFAWqVLqQ/rCO0HHwnQnfLADyhVDT27csSTk6QD7
iD030DXXKi/kVsHbvocMQu4RqVsvRQka5Z8Y0dEFAALDP2RyQtSkTVjS0x27
N/ZVHCrOvv48AL5pxQ/o4iYC1etdJJ9BJeGSIXDvncWmmoOegqE5IFlNUbnV
aAQcKxUgbtVHbZXCbB34a4QINZ1L4lOJE6o3EocGyIWD4zw66AcfchZyp44V
osyQZ89D62I8DPtD+53bJrb8vDu8ZoOXGqUnc2GvdtXpaiGMFZE7kgVmB95H
3aagVmIwGHavduA7a9d6/bD7TUAvm1BTr90zmMzDJeXSW+cZ1BK+TgkeHrIW
3vKcssn0xnCzG8M99GtQqFenHT3rM1tlAEE0SRjunT+if5bwcaUyOdveeY/L
krnHubyOU7nMENn6GTUbceCDxNOAqgL239+vLpqNBsUBu3JpYA6DPNA+1SP/
x8Ja6CIYyrTnWesCYMeB1fudcLhTib0crY/6kciYHZ2zisXSIhBGnfwkX0G0
mZemMalWFcbHU8YDyZt0iJlP15ZH417sGt2Bzgamd7n9diUbQqJOVqEJ6DU/
3b2v4VZ7M1t7j86Mqo5I3CCARftEazFCAQB7b6NJUmbfWa7Wh9OSpyBsS2ev
46Qr4kpLOCg4pQRQK9f6eg//VWg5hlvdLjvHYARSz5uKTn3BC0OpT2jEQwSc
85rLtzd3p1mUCwCRXle9rx/PStWmwyGnddlt1tOzY+qLKQXZab8NSPUZuQ9J
CZlf2IA69FJFMkFvOosmADddB6XlNqk2TpT1dvn2KYe3rgFHQt+ChifuQliY
hzADYrPek+ncNnIiX8ys/70CeUtge7Tp7x3ohvRVZyfHB5Q2P1dQLZIROiPY
G6UMUV8gYIZOdjXFxzjjyLfO02lb7IVInbG619JE9XRJaI7RcHkjg4JFgd9+
xuNgAoBV40u/EV8rHTpPbH+7OW71FPOyQy4/YZYv6uIeQlGdADJ5FLFUvh9H
uJ0uAtolr/D9fe8oV7lTPwOweDjj4vcE9EIa+0tydtRGhBbUiC1Wy7xy6zg5
Gy3GNk1ER6UPzuH7EaZBW8hsBwbaN9WDZ38yF+JEMCYLyqjcF9iRngy0hDnp
Iyh/BCoNDtv4k1uTAtFwGkWg9YSipsqXyH0ePpXGhO7tmy0p5GvLTKxSMRW8
NYlEHCFrhP67vSihQW0Gn8YNtx+93ATsbkEULkS7TOn1GwgSczT+8qdMfXZX
zTP6fKM/ZejPXlvqZbP3m/VVfE9N7EJHdO05yyPNY4DxEf5JQVTRfugql72e
Uz+QnCKsF3qoZy9kpecS3JAJk5VIftreN8u55Lgd6PqCDbs8kj5m3PqP++tI
Fml4HROZ7p41QvDW46GFDfmIWnOOb+ndebvy8vn95vWxPCYdU9GGv3pwrQ55
S1HPJYWnRcMql739P+C82JiRTQbsARsCl4lxfIDl3Fm1gvK/LN7oOO5BYLw9
vjB+hvuawfWqMbGoq3//mfVqAN688fszkmWl4xeHle8PVZgCH/U/m1vvriMx
obVwgNlGdCaahgGjXb7YWMd+AV6EJeNdMRpK6k+M/OlSH8HjLLYIG3wSykmA
fgDytxhn2oZuKM1SOR/nfdCn5qWO0/ltk7PlRnmrpCLwxa1prQN/SUN3Rrwd
yyVc+O26zSGnFEeDaQm73kmgAiOBw1qtDRaXr8I6cy3dZZFN1hy09rZWd9Tn
b5seI3PQYZLv3tk9l+qYhMpZ33iNoZ0osfMFtAxM5IzYIiNd9uv+k6cvOf5J
pM/qgHVBHYIASJtupmLjVrFbx629deX0VxUeaZwMMOwB6SYOOr0IUxP8EM5u
nOKGtmHhnxdyocY5S95qqDB8mkascW0AT0ehiIib6NmmP56P7CEVIxdEzpLB
gmlhNLmNf2iOIs/rIQqb/kpFjvvI5mDgR1D8/KVnBbZWI9gHvvSfpcqCXayR
zwcJtz87woxgVro6gbYZj+mNBrPv01pMfYi6TFcCJB+eC1fEbVsc6WMwvtEh
tZU9Rb0P9EoSHDWxkgEUBIBuw4N5jBYgVTer7ha96EapD9HZuSrSQsRMO+oG
0MK6fQo187Yr+P02RRjJFeII0na+jTkcRgC4l42zDpgWsYELz/oimEsGe5gj
jK16h8eTtdjM7NT5bM7jsnf5Wo8tBHZfyqz5TjB/z0aOx+HqhCiC7uXWCZ91
gJaG0BiuYCPcKg0u+QjYRdDI1/iBP9Ofe5L5yvPJ3tJ+zSDWg4Zw0BDkKnGm
ipIaF7gQ66bURCKHCCkO2vChKovCo1h8hvLvymXJkfwlwEjP5fppgKfdilF+
ELX60HbIFwnjyDd8REZiYJRU2jKpk6mndswg97zU0uP5BDBUrUbvMw12/yau
K/bIqC2f0JZFf2Nb1dSdJoz8hiJSjjA72JiDryfeuJ7l692IjFrXJLBiW3nB
sm2UW1N40TV7W3Xzh14db5v9iCVBQgSNvVFg9y/mobNyXEfKUyg2XSYBSHuG
Jx7B/oeEx/hsqzmHKNYnNiERa3VJbJwOEwqfP1lxssJcV9VyU8y/VEr3KuCR
fwF7SMxTqldWge8osoPV2UYItJ+5bfVGeKP1qkq02u8Jxk7+UvEgjcb5UBqZ
IDapYUKKku2jKKkSWAVKRXP+oSAi2pqWv837xXk4zWkoWYWxkIpKDlhbgAGM
e1r34XhGWEN6Ga2PtDJtTIpZwyFUgXTHRLaNZbsHxIMFbcEMWtdL9eNgvJOX
rjnrun3TBHuIfj6vVMBaZgeVqM0BhtG4+HXOxj48funbFxwmMTlpNJtU/wxQ
Y62WX0nqv+naISHBHW1/xqlKgEHkMl89TTu3KUsldkHi7ocuarJ7dvHdx2Y5
L4gf6ADfSYhF84xx3xJWl53oBzotLJV6ezKGIftLM1yBl40w3Ofpg/EmEgt+
xSFU1FgV4Zs+oLpjnidm3qAUSjC22sVSI/zfWXYEz9UNVdtz34L2Obu4FvkZ
UmEOjhb3eo3L3c/yErD8zrM4FAlpnUrwalOkmyU5U7zqgoQ7+Aff4WJuO5UB
oYZM4UoIMVEGgKxCOu97jnZVlhiGjNceV+AhTm1SiUos5pXIsSe/JzGYpJPt
TpVQnP17P1k3VS7i8p5W/6ECnvXksbtbcNB8GqAXyXqpwV8jyy8GfX2ggKnh
2D8MPs4I5+4mt28rIoyiUtpjnPzI1iMkx2rCgQmgIUKZ8wS8ZFHrKGBagYQi
/qz9YMEItDfEEpeDYhjpqcDkfmesfH6cB2DwAo7P7Swbl5X74M1daPn3PCfL
ED4RBMe6qaEtiWeg+SFsNfxH1OGq/Y0xVhd5o+m5VbjEVCwHaY9orD6T9eUm
xtjUpuKYl6B09w66LAvx6uFQkcJGLDy+pERs3frvfZr39CJfrtC9H8nM2zcg
rGGMlKfigxxyJG6N4wkx1/WaPbmdv2HUVY93WvDy3va66VbYn3xRrdJM8oHA
ylBSOx0SddlJzUQeHZ4vGcQqYAm8wIqiwmYci2quPoeVTL4eR/idnz+oVree
WMDRJ/7yWYVfOWkeOfXcerUVqG/Z8IkssmI26YcdrOljnTkwlanEWHjBVLPa
UdW0FBZjRXzXBplXkQuRvAG5AY6Buu/rn5fU9BpMf4/oszxhXIlikiBDuYgI
hjRMROwqEyuwAo/OY7vle6Km3UpqyyU+WGOyw0JFhZZv4L4JWZUxjB6fVLTb
fbdy+gKcEti49XMb+7mFQAtRsRcGKTlHAGmXxG2gcbBylTYTddGleQx2LmdW
7S7LAz5Ni4hggCHKKLexBuniJKWILf/G3DwRME4MeJVnA2rhnrIzHeAJHc8+
F7dd6jpL187lvgjdilUXIZ+SOFVnMSCTDdwYtY0uLGb6sjmhXb7e67MP321b
p13ZuBq9e4kiSez9WvEw+dktHHmMRuYt+SKIJEXnk18It6TSzyasIMWXVu5y
+MmVxpy9HxDKyx9nHpUwhamf4xmIzvLo6YjsidzJfEGVrKgtcCQReBAWlCt/
E4iXwRT/NR2sOOYiHMsj2fD5BvwhENOfFAP/ZJnu51GNxp8Yfuktbmhr7Cnd
MJPMgj52BSALxJUeiCl7poV0RHhGS9fZlBrFTqpj7va6sQ/5YjRaCo05izn0
zqCA8kNcUz1z5A1PJZS1O6aLTX6CnScAPJf29nw54ahNrO4AsUZb1ZiY0JiE
8G4KAThDd6+I5SxRhQDD6h9+U9KtzM10qN4a7s++NSxmtD3I4x+x5vcZuJ17
NohFX0DJqQJQsvqFaXQKkJJQMuhVcHczGIL18OEaIXHjU3WvzagCsgXHENzv
EPF98Gp5EnqvaxF5Yi5g9W44UNr6fdwUh6I9YEjcZt4gA7fB+qy8hAmJVjzf
DLgQocOu9gqEQXh3PcnLITozUtNSFDk2jkQzQhump4hJpdT/7YrfAuyYJHWR
qBy+pKEBOCBKX5duyhMqcJmoUFSTZuas1wxMvsAylU7XYMRYJa+2vJfJAqDD
VwCaQ6/Hk4y0uRkHy3ZUCdLBitmCt3d9Jj4BIkfNQ5l1zBzSJiD24lRav0L9
NVFmX6g8208peOtOkaB8xB+/7FeAfWtnea0XXWTRYSL9+1cwVfYMTHIGlIbb
hKvUJDHnS8ctsibwpBjc3HvTJGDvL40BNn1m0ewIqf2dt4pGWavYHgId4NTn
GPhRIAYPkqNdNDhFmuVo1EKotN1TGfoG6JE7w6DmHEUwLSwl6HBo1MvjDVh9
AaqJkIQyzwPu7Gi7NdhRT7+l9MTxEta3k5PZzuGYD/6MdMy5HmqPoZ5tdNO5
3Ds9B90AFf2Vef9Qgc5ofEGSE0r9+1lOuY9irbQuu3ZRdfRTqKNZCuFqHPat
1p0ND+8Kao6GuxPICB0KNrXW3Q6af2evKv42VpGaQXY7ycTz/9OWnwmsncL5
bsKKm4G9UzTPANX+h2Y+U6KzlIYZ8eRCd2T5MmWPyXVRgmtqeKlIJ4O9PGtI
p+CYa+MlD5/frTywNVrHs0qIkuWDQSj/Ggp/JKNIKgmgT9vdfgynaGKGPp1F
APPQMKoxrjT2Q9XZv/gR1KdW3BofkGvmcLvkVOir6ARyVTp8ns9ExY6v1zvk
QqrzRvY9UoUOPywR6GJwFgpikFLxO+RU6gyOGAuEieK42B7vRS+Cl6Tlpi9a
Dyb2kbJ1rqyfEoZnCMicZclxtMsenjV1Yk5Ps6La8WHLgCsllFaVqaJoiu5g
9ZMwULaiSn5vEbNsX6tyJhmw1UiK7pNM/fLv8v7JAmb+pr1Pf6UD/FHKfrI9
Dqb5AsSZR2rdS5So47ih6uP/s44bKDd1QG+L4XT00uBMA4SlUfGzgjccnBPs
0qcbfr3N7GUpDKgPgrAaeOdrqjAPVLpvRQZ38DVt2eMNtGV+i7FnGBaWh6FQ
FJSnCwfATZGcFAAbmJAZvrgYSEc5cLuoNZRNOpFxUVYmR7wgWYrLj0S69vdH
rUmqvZQUT9ljaBZD+E2GU2NsWSZP2WPuom15pI5tzA+3gA84waVSVN8bX/fM
t3FfchSBPJ9ivxu6Dz84hHshDv5G+Qr+cBnjMOAmgCn3ysoefjZpNivUQFrR
kzQtjZxVoNG52UbBvWUq3lZNbpAm6zaOBr5Tleys75o6L3wBwEFoqOeO+TG3
F7Zq0SoMgF4nZgNPAsjofaSdZkQn4nR47wgCoRAj9QDAwSuf+ThvLfIvSLfB
flfTZEo2VrLFjZ7cQfu0RytKKjHm20ZTilUyFlKzoWKq6FmCirxbmBPZWv6K
XEZWxHZ0c9vR5UPzatC/B/yS8e9v2c1I8ZsEi/ytMCWKEBvqug4Eyxxpe6xD
9JpiFezn6S6HTn1Udoa7MsBmcOsOUUip+hKWxXyNqZ1CzrXmtUDinDpj2XGa
rjZmZOfbAqp4CG+PKAYE3t5Qzli6eU7CjmmqiHSy35ypazfIYy8cDFH2Svj1
XkqYY+SwDKQff8Z95qWdp6XrGrK/3TCbTIRfB0qJt54+r67ilMNwFkeHUf5L
wH07ohiGiErVw6xQD+QzTXpaqjWW6LhTeM2thpBBV3vhzII+hmR2RjlcDXri
vEtY5ZDQi3PsAOfV6PSz2LFkTecCTNxKQUzY/9f8oslh66FbduUSOPFinCkz
MhbLX9Yem6PKj5LyV99ZW68fvf5q+5m8VLNSSNsy2jbck+bzfx30Ezp+Oqqo
/5vWb4QKSuE8f5aJYb61ttIcYJvegYqZKRzHgLU/OZ/EGU3Mn1UYUFzy91iy
po5Sc45S7JqHVBWbQErA9XsVM98oqmLa/re9IMgNIdZgLqooEX6/E2wpYtRQ
lKGjO0BfbRpmy3c8ghA32l5nuYOU1mavjXeFyVIfmHVc+0NcbFvs8bKBwB6Q
NwTUB+L99Cdy1o3cFE9YjP8cxHCLTnemlJK4BZPe9US2SP3ZwvSciYEGKoOR
LQ5VliaogTDnr+q438LPwcc9ZQw2AONg6mI55KcJz7IocS/XCivUeq/PIb99
geqol816BIr0ED0msC+qkz1OpYtiUOfYK4/B6mH/J+U23a+Gd0oeLQTBdmhf
NMEY9YK2F31DRcJKU/IajC8s2ZKB701PEeIiQkaUA17Tl0LhTL4Gh9QrLTOx
ZMhIkl4XZ+2OosWZXz2ePvNjpvAWydk/xI+EYwSVWge6lyssMbnuZOX/zO+N
ruJBosrtQseRJW1wUskxodbOzYwb2wmVy36Adcg/B4CrH0/uiL9XF2zata26
PP7TOUypLbqr4EWEB2XeCQaGfUeOoZ91zS62l+35CVGRW9JNr2Z/zFeLHbGx
5h0NkbrRAtAu8qm+8JeTqLB59+O1ShdjdkrHQpZg0R50mjqKEgHsalLVlvEp
fG17ReciZLloVuitDeAgLeGHwqOGu/3aSoPeHphi/6U+bGG5IMUHgWFhAiRo
dRbggD//XtFV2h6GhyBUxoYnjlQsQTZa0Y8b2g4BMIfQ5K9kWye1sLbNMqEd
EDUe00vsv+AbTxe0jyIQimjnVNRvpS4KtDNNBqPHU/jSmDAonX+0jR1vcJHe
4QEOmKp9kL3n37GWPdICgkIG06aFs2FrSgYNyI1RgnT0fhabqZDrYQMrooqq
dXvVqSGXjPNcs6kCvUpnHRywBC+BWnsJj99FNrrQhp5nRIB8QOUE3c67tO/y
+hwThR+c0uU9JL0erygJ1Nnag0Dj38dxnB5x8bnAHnA8fanwx4PdBgBkOV1B
4zxZz3/77TjXP7NvJCl1K4KpIsSca3YxWQiZYP4LdjKkD1MlhaH+8t2Tm1jl
RmKPF6kIDhnUILQ5YRYfqrUwRwbou1pUAJuDJYEc6TJ6gdtc/2ysKnV8rWmN
jR1sB2fYtreY+APLCQTsAUAuZcTpNn2hlNuF2/Jio4yueytRaO2kuEMjHrAf
nnqR8O8ktXMz0NcF0B9EhbKPSjrUBA1RbJlr32nPLom7/pOi2HLW59gnuJRn
b8QuvHG+o3XbEifUHOmRBtfK/fk7DMBoht16MLpGUSilWHO4v2Lmtl9zWJ6x
z1p2JwIEyE4b/OBVlRoFxocU28SWqibvlD5koZioum2rAO0hNsVJeHcFEl/j
xSQwHmDTLll6EmIN0cjd85lrBQ8ibvEOe+5MNKzpoxuYtg7mZzvJZOPu3Xpn
IK90bGZgvgKl+1iyEAGcYOBwlfP0EwLPlaWJ5dRtZ27qpbKHIBMQwHySbGAP
44aaryDcO8HFsQ0u5zmFySvdrWgyJrHBm1L9MlbW2Io7w3ttGpnIi1+q/ure
DE6Rq+pWNiKjCZ8ZfM9lbhYtST1C2wUEftQlHcLp/+E5Gerjfvekgco4TLbX
e9raoeruRqB85Hf9Herg6B8o9JanGDta1Dg5rkR0N8HZGjM8MlHsjGLcklng
WrkASe3N5JzzKxPHa3ILrn11TvitTyHjQiSfoINBnjy9n/Z4MORrTmpTIJC+
fjVDtRKrOgrgYIonKgHPCCTnzUbVPJ1d47CMPshv+1gJsTG6Du5hScOksUOV
Jw04S1xk+YFeYRUqx4iNnMci1l9IJ2tZ11Tmd0Gmb72tRPWrOhpYY6Abfgbz
J/BqtPM/4ora3lj3ANXkd2Xc/TXFZ/WZLiw76RtkQZKaYZjPhK1uM1TtNnCS
BV7TFOD5jyZX/sezpgKejW7adYo2NpEg05U2Bn2VMKmAfHES/C4NequmDicy
hdf+x1Pr1aE7E3sAJ9IrKIoKIbHszxO0zuqF2TWTuZBi/5c7zgPYDDmVIcM1
KflL94CTNCXN03xMo+6FpIjG8qSlC3GX+NDVMynY3pgIzWvSA3xO9OlNTgEe
vZQfwn1gdT6x08p5b6QpsDLMz4ojWviOoD5U9080CczWEwOA7QGGyjrf2DkD
RPd3urMVl0cOqvpqNJGD1WAIN6DHrQ5K8l/vDNrCdNBTMb5009ZyfOWQPdjA
WAVE8gp31ApqcYDV0MnZBJ9C6E5ZxSzCKPr4r5ELyS2ZaVn1q5sVG3q3Y09X
x2h47wiYmU56ZOAzJSIjWUZQS+e4iuD9FJnc47+n1QClqUfkY7/MBxixM3HC
bK0r+JFrQQNNHXStikYDhoZlnumAaWBEAxWX2r8tHUAmQUimN8BtUFoWPpyB
gTj8yzRB8xFdWTvkaULY+SlwlecCjQPj+eq6FTzmXk9wva/mGwCmU8BpFp4U
Bq+pUq01iMAza8DITeQiwHjsrknZPsjUhdjnQHFg3TJg3nZ779jC0ENeIsxl
eCNbDCb4RLF6rbDxifZ+JXHCZSWcFUAYQYWp3/RIgvwH0yjbkcHakqjuBIjd
B4ovit2DH4ry4oWzmAWt8IgrgYt2FlO0ezNulHfvoWko023qRQPsDrUD7CdA
gsKUASj7h8uQv74IlP6sCKBbxlvuEi8HoNhe/Jk+NGf8oydsw5ZhHgjoDfiy
jcSl5Q9jUYm73jaJdF5qaWeL5KjsvhI+MBG66vsyqKqQuVGGNH3cs0vsKr51
fGSVlEiH6ZyW2yVoco7j0MmFUuWXKhHCP4twhpRYZZwDy1oPIwVpiO7lJhQZ
2ZfiDlFzkXdBcZkEKY6k54kuxQ0BBMI1agDxM382e2qlvkXwQkcvVJpfuUll
CohiGjZyNrlMPHugK0+u3DH0usnSakrsLDHGd7zyZBklIMr+4jl+rbyGk2VV
IcqsPYsEImYD8RSEhGFdOeiXyk3NL9KKx3mrskn3qR/gexnUJ6maGSO4z8dJ
svYPh+ruNtstc/0fHgUz1lF+IlwXV7g2XekAXuNfH0l8NyIZP68ihqu7FzMa
lZfP8n8+fYmJc8Nko+a7d7rdLcCj9cd3sixCz5gNULJ8Fy89GxIKwn+hDdQn
t/SHIWdimV2N0lS3g17h29ArgRU0ChAuGNI5BFPNaU034eNZbyZGuODEt1EU
Zh5p0O9LNAaPih0X+to/WMvjK6Kzz2y1sTA32gdfffOV6Yif6QMIN45yCkWX
UtNhsSSONjZS7rE7bOQFAzueUBLi4ohVJFQU2iNPyipa5ykPoWWgJLLtcs90
LjDJ37/BOVpSvPsQTFLhLSCGcEiEONb82wZs8J9RNQqbblFfo02UD8scMbCi
Jg9M8yCpFXz7mAD8T0uxeHxpSHDVK57iuwe1I6oR73I6wvpQp28igefjFpZF
jil4U786Uv3hpU4TFb416OwIjPo9M2fc36yHvrpC/93NLH7SDkEUh7/4gFHe
UeX0bz0ZuQQqEaeFXWbAfc4WOUsKD6XDuc0pjhKfzls9narLa03y9bHPmpe4
uxPuVbdN2nf7vPL6o2gVh6NgprO1qAodxowNwURtjclGoUnnm/QdGHEh3yYW
aqkDMaVsIDNaB4FIQen3ShEZ2IYJU5akSpjSyU/XXkwW+LJk4uE1+XDdXzbH
9w6rXIAOlGf7EuNyKypFZNrqqrrdgMA42el6hX3yd1dEOxzc7QIVTQq6SQiT
ioyGWSfq1JvAJdrXiFc16K+fg9/lU2zgWAyWDOFIrnCSLl//dI6/ru6q30oh
kScSDmPdHPcK5QJOL+/Djl2uImAuwqzPWbeSVRPWhhvsQGCGQt8MGyj5hCks
saVKYE7RFyNTL1QiJpc4c24mWce3nIP1J02ix14CRelW5QmELw5usVwcQ2Xs
qbThm7j3XacxVmMCjRGM7NigE8ZlfdvmB2qmAjRJvJamIFjTzgYvgl/Iwm8a
JxP07jFhF5eJ87XZkUOnhdS+qMKz9ldu2/dzvRLEFGZ9s4YOhg+uVbIgx/yw
lBmH3XodezdWV+NbLPJoqk3n5JPN/4Qbuk8EQOLdF7tA9Yx8jaLFBG8IAkiO
UdmA6FT1rz3F+GQbJP3lvX+pGGdn0gCAIo5Pi4GDUV+YscEF5TYxIJFzRMPG
MHx5LyVSOT9AvQ+mhJNK/NIF4qOOQuQxBzgXCqYqVxPH053Ifk1Ee/v3VvtD
eHjGcHDKTwWTEZODQlDIChdq+OkVcyHb4iTkjXgJQ/eplfl7ENbjFVoxkehl
fMxyhTOoqslzqGA/YB9kfUxGkEKg4r0KaqQhujjDt4hW0cOvClQOPLoflP4c
DKLDKhOBru2biE3l6ye3jDSCzxwKjBDIJu8oJ/l4Rp38KAASe2lufct10izl
T4O5NtRZYIcvs79vyRXOzl4ZW5AMQKs0ggLidTezZsNk5DGXeyL28E5UcA6+
sPyPKRT+05cvEESl9J5+IvStMVl2uNiy3sgGIcqJZhPzTpOZFAKJ7yv2uKhU
W5Nz3YfMET3/ij4PNUXqsGZ6VHcaMIOfJrxcuRq7gXXoNzoDfwrWTptonh1i
PfnppC6CK1L6HSBnecWvBAvsq15f+2qYdvzdlfpIJAyfhLwQX/wi7CoJLXfb
wSt4Cy0hx9p7GMC1py3qXGW9F0ai90s8E604NSFBkR49Pdh5MD7Joi53FMFC
TefAbwM5aIu/WQANUA2/fAmnwO1Eqgjal6FPjQSx3U49ducOYysx35fNabrS
QE+humfbopTqjFQkp9pHz7PZXgD7V2xTx9dTBHrt6snYJ/q+1+/PhHksEtzm
Zflb2TExfditMmQKsEgqpiwlwpYe/S8RoAhZfbLEiEFfPnR2+F61SrufZsPr
R9acOwZp9yNcIgrCeaubMVdixyFFQ3ZfsjXLIjcqMu9k8ppri8QZxeEUhvye
UGO5gHBDyomlDQerJGe+DgL7Uk900bcuaNOCwi0umHSs2+pqjTnmMquzPHcC
smZAHqfwfEJTFbylpZL2cW8PDjSgnLceQq/nNRHgGxIbKsfEvAemdDGE1tqI
wJkP3N8dv3fUXBQTwDLLtxi0J9bziUi3Le/nPzbh2I+1geJAt/sN5GEmZNcR
Pl6lNxKNgSvSKjZb/FqNcsFvn+ephlqCPmMw+bC13s0MecyH7S/a05lwlyUB
56knP7VIiD3+F4wj/D6gbrt/JIKdw3q0APtdldPUaX2LmNPylfKI7GHhbNWC
32rw2Nl/ADCDAOHhzACUGBBjE+ylq1RZDfONeC3h75/7GKXmBkPBJBCK42zh
eo0bLIaylQEavVfA7s8z9AgKgasOzmsE5gcZ4/Q/rnonQvEDrOU/Nn0do3xs
ff4aVsoqvAtTkjat+rdOde2QBfCqTcWI+NZ036WSbfMLmXgXhR6vfb1DYXPq
JFP7ompFfPUFtRZTko4MZ8rErlwqwXA3P4O+EPjxWjWReDqUFgYfWc18da3P
FjdPWxFdymaF3RUUmZKmNsastAIS8V6HCaCIhRspPnwgaifIchWJvl5Wr452
DnoqBgphZNSgph/UH59b0LYqVcz7WILBO05lP+WiuK88ivH5/98OXl7shCN/
C8mHb6zzNsiJ8SdntM9ilVb8sK7lS9bEbVoEMAI72NgZG8tMcn5T3727CTDD
uBr7jZNqB++VtnKpDompCtjor89lScZqUFfhU2jzB0Sb7RclfoYXwX5F/zQk
Dj50WhKSEnJUCf26ntUsOxXzwWJq/MAL6g8X6gAk/HEDnYMtHPSDYbk4Hpaa
rXRZgGEBm6R5zsU0IxC7Uza+wmk7Wz0ZQGS13XUZ6TFmAljlUMXMiQSgWChK
WouQha+MYbSxNIEPyt/XkOAdUbcN9o5/PaRST/Tz8vHveDYbpOerIoC0DdvO
lRRYgPPS98kK5dPm4XAURdCEV+K0SPD33Ewj6JSvojdgPINNpxjWBJupS9Zi
AVbXrq5wFoEAd/wNczXcuCGOOzALI3g0fRDPMfd8zr8+o6gQW1HU48Df0paj
sY8br/7s5dO8D7xogXwcIZhnx8kgOyWsICdY9phSFVt0+KAd7SESyD3OjjgC
/kEGkPI8P073LlBe3tmC4haOd0XUSBdsi7k+5BqsFBJqwoP5soV58CfaO1+b
bMlSCI6YQY10orBQ6ti2XQc9vLmvzfJorflbBb6VgN2XHcPU97SUGQsAUZsx
sXjJPMjbXETb4X7Xejax3fTOmEHBQ0XfKoLXgeojjXu0jnRm1prQn0Sakn53
eR2c/S8l5NKkxCJNwOR/zqyY9LUfejczwAyz0262GUBjCPHCqe1zh7VYbSI9
pofx0F462NLMNYXiBSfhRinp82p1k++d22Pfk7LRz4CoVhYn3K5VUcaoVvO5
urJxtENMGL/qWjOB0+xzQTo/pyBCF09g07fwB8rkOvu8fp1FKdDNwmLSMCpM
mc6P+C1CWLYLUvm3q4g0oohCvaKarDeerHyRhql6HrEZQSAkxYTBIMDQTALg
zSlbbx7Y6qqlAkaNkhiUhbsSfPmdFNGrTZGl3QQDVhlXDdPdGmlCTqsmNlim
Gwd1nNCsmlpKbS1GqkHPtIO5nhqBmzFrkhIHfhyVgCtjlsDuOOHl+23J5HzA
jQlOBzo7kOdvcuEpbGeazAz+916tljoBAET0wzioxmMgRSaJR/hYyvvAHl2P
96ZhS/mHbAjEeaQ1yTNzpHhAPlKwgfg6tsEBK96iRfgraT9MiwbgWOndff6J
ankrRFU6PtVoJQpTQM8Qvlh4IbB60Ht7WLpSI7ZJQmPyhPrqOaHYlcyckQW1
4tqlzrvftoJMUIJeLwpMbGCiBbcMBtMNpNB2hPVGOfW4WwJwGYtqz06XefcM
7rcPCwM9l+m9vqLWjK0bf1z3D1XC0gYnnL7PUjl98JPYxrzIckzmGiBPQvh0
s2HW3RDoGL8TKIrNeyCqxIkFcyOapzqIvvq1G0Vc1j65ZPDZqWxs5jEW/MX7
IRW/85bAV90tMy187SXc0kjqJKctmogj6kJu4aZd3PjMhMwI//Pd3ry2nz+r
ncsTgJ1EOmrHZOIQaLip+rk++zrowhYaKGqSC0ZB/LqCJCe+DjytRGC8vZq8
Ddg06bc7/6GTN3Bhb6o2t5yPFAL8N/C13J4Kgi+LxXFWdZ9fmN9FnJLBrBu3
8XMxuiLlZlw3+LUUnMnl22pHBE5o+agxOK7auKjHYnK056xM46DMiMsAoQsU
dPgbMM8DUNT+6rI0KoYSeC7h6WDZ0GS5jTjwF5rY01HMGQLisORLCSGBcfyb
wrY2rEjt4VqVoGG8qI24lp4X8q9PPHID9ey+kJYq5symTGIFX0y6C3rgY3dx
72nrPb//IjwQfekl/BKSxI1O+tII8Nll3WAps7sUTtqNvgJ8rDmmP9RgMA/1
7ocuvO3IzUvIU8fxWR/QpE+COdUTVFSJxH0umVjMNWc74bgwt57Y8TJ7q0z9
ukFfWwPESAoX8cnXeOFMmcI8efv0mV93Owrm2xEf0iYOWaAfIkEgXL310Ies
ZjziVl45y6UEUajq4bqzZ84b/SZ5eBybJ/x/plErkCqCeXxNAC5Kx+oSVk6e
A7D7SRS3rpUpirbd0WurlNh/qFZHypV5CY1aY6MvFv+00xXye1Q0rFqhwxbA
hoBytMOaA/Lo/zA3FjlOismEiusKRBJvdz2rKOf2vLnJdXi97IV2gXIkJDbT
gAWLC03dWv9TZyuojXGOAASQ0t1c1dOuvorGa7ttNSthu6XZLBIkv5VCUNld
RNHyiU7go7bS45GWaG9EWwF8B5tYE5cL5Nj4VlDCN2+SIpmI+9AiykrvXFEv
VM9n7hLHa2tc90+u0Uu12+bol72bR4c4Gkm5ku9ErzIYajppiu5CsHmzKG/h
EPPwYZGjUV1u74KbqzBma22v0mgj4CF3rqYhaSbwhvRxCjzRxdcsi5wLoP19
GYhOCHBij/HM/XBMZscIkK/+eUWP7g8/xjHKDQvR65z9M78NCNe57rAIkCS4
LpNxNm6yB/AJBhRmX67bc6oMT8Y66L6ypcMf2UwZ4AOoh9eAs7SD+1qwuvrY
ZhJKrmiwwhjYzVUIzNAeaWM/IDjxQ+65XiYYW5YAU1oxuO42Zazx6VPa/BDS
YbUGGjG7+9Ood4p7Su4TAJmWHqTlu1OOJpZnYqllODeIJtYVzNUROf9/exMw
/FlAQojiyMc+utF9xtABj5p75l5gptQnZkn2ppeIINcV0Sb2g/iWmeTkVjRM
XRnFcA8QGZ3+4uWB6FZntaWWZzZg/SlpZ6qoAtxQiAbb2Ct9Ok7880x8iSGK
Ky3k220iLfV6jh0yIvIwgE4tSHpBa9slfNed+Sspa2l1xAinhffRyjWCstt2
NaIv77jPVzKOtBbV5z+3dX/eh7p00H4nT/sEIeHL35F1uF5GrHwzqx79fqEl
HkbpPngTpXUHtEwkzo0KPVPBU+ITQVVZE0pubRHNpG7PO/Pe6yFcRghqZ+Jg
AY2VuyHLCDDNn1rhT1vibJ1LuLYE1A3lkG5FdXqAwCQ3GfRpEO+eTy/2ktyp
9x1hH3sasuKMsIEDvIXDE/mlmmRaoT+V2eLxmI8Q5i+VS3XN+HvTks/g3MRL
+zDVG+8Nhw360SIwv7bqgC6yzuVwoR6CD6gk1/EsWInrglvGrTBGp9JMkTBa
sJwPVYSOQrRdIUyQL0ps0s8oF1LpCK15fvFmDU9z5BTB2TXBf+SmSk+HSDDK
ev+6NZz2p4BcnRFfyquf7mdDGX+ZlxEbpIc0SmT5jBgZNFnfDpbeWJY5sTYc
WNh3aadIDX+PTETZveOto3myH3BR9/FRjMdNobO+tz1PtYr8YcnY8bMmsPgp
hFsiE0q2LB3e5dmsLZdhUWtHehyqmkVWyjCUgWKeKxiPcMTb/8qkze8NZJVx
e9AeGw8DGZV3LH+oPaM07lxm6lpelkHfvc+duiZrhIQUWAb7isAMWXVOv8BX
l3ScCDF0rZZUzJU7JdKUnBOd7Efxa4Ib7i2qbybzX/CK/E6wUY1aJLtl4QDS
vudxjEyHWrwerymt0zHB6LXtj2p75aBucbTMaWik8E9fNka1F2+DNGce14Lo
Dc4ggrnwW+gopiFzRrCmd6C69fMqjisFOkUrgGIlJxItM2rhqYQb4osqJ2pE
T2J03A+j5BiQtRSi9IIRmStkQH0xs9fi5JiOKkqgGc1j6v4dJsOOGQanFa8h
uG1snzm6KG608ntpTM4xEEsgWC2FmI2mHhlQ4paVOkMWTi8Frv66CePTyM+I
OOXsbHVwD8hPxd0UaNW2DlvcrjkfRCFKtpPo5DN63+4Q64azbu72aJ5dLTSJ
rrUHzZ3SqMuKRPyFi+yCXqLX3lwcfRHWeYcSAAgbowpSEGmzcG6dKpojJp9B
kzJYpZoBogcOaAs1Gb+YazX/zSYqobPFJjUP+gryZzDWIzpz1/dY9YAGdgKT
S8NCysgytsWtDGzn88g9wZS3XPqKf+q+ke3qPZXLD1H8EcVw1UFAQym1gnKt
nSMLhJY9jdpi8yV8xRkfwD4ISTqkaEV1hja6FNRxePt6Ef5P68hvb3o0UVRL
Gr4594Tunnfn3w7n93Lryyqem0yfIQx2TIOt8MtB1jBvUuI5pTXp84ljvGr+
J54fkI+xPrnmdFAHJ0+/RSDiBS75JWFMmRPaTBkzFvan7aEm8mxdsZG4qvD0
kUD4ug5ByjUsqNDtTTIH8PyDhu8CzGeDptQbRz6evVq2JODEkSFAabUzdLpF
T1WW4IctCfR9arb/5UpUEdg8Uxs8tbcp+nBbnsDX9TgaLLPhDeUYZysnNhk/
bQY/yKn8S4t59G2Z7Lp/t06MN4TTnKzgCdI8KU/DH0LfaCABMcwUtiV9frFt
JcdNzidd+wtsqWve2jNJJeabfGcW9S8TG4DMnjTb2ewUyCpNR41nyPGIdFcB
qJzFqJxEJyLjQypO+i4KXwVHZ0J+NovfIlOpW6c2eAqXKeett2KlqRAKtYGn
yEQFT7lmyGPnsXvX4MU+z+L6e0endKdDdBuqJRq/eGemZjbEXx43crUEhTZ3
UhJ1Ia8A5BceLQVGp7rKfK6m1JhailGfCVe24a+CaGUM/LNOU2Ku7QHxec7D
TesAb7y5qxKyBEdji0B9PWjowaVoEeComdvv09rKQlGdSbcQxWqiYEYAuMbb
nb8uTUspNHGKXY9WwoN93kg/87NLMyhFMNtWzWiPXEaSDlTHrY6sJQc/Bdyz
OISS/xT0UnN15Gb4Ui2tKZcOWYNkGMBxdqRJ/JBWIiafW4+ywSslCqAWiPpj
l6K0tTPlfncofVA0bbWAKNKs9HWDRRHGWmJH7g9mduwAVUbDRfFrLk7XQZNl
ZCb1MR7kxYoNSfUY6mNOn5cjLPkOpypM5Nu74/lDvJqFZ4M883pU9+qV7iCm
V1QLS3npO2+fIIJ70lSivAiKkYt3Woi8+MidMdAR4mGpGrUvdlKZ/1zUusbn
jg6uU1TDwJmhiGb9rsCQsPXuXufuoTk97dMsDfm5Etyd6x+hO7jdxJrAFRPu
F9clJodBCiAJ+GFlWi+hTeYS/2tx0gsWvrbqR3ZqTFojbe5vpPKvGT3N8oFf
6u/jk+hbqcuR8g/VuAXvnfTBgsgTBpbO99f6Bp1mWBANoqyr7gtAaVTpPSUP
a7+RdqiLpWHzkrNJ9mEKKmhU5E8Pk4pP3lSjj9Eaw2dSm/LpTsq3N0TZTtVa
T75JqjT63Yz7j8jwc6WCo4sY4G3A2RsVw9f35UTcuMk4mrnyU117KfdIa2DT
dtxltn0GzufJXKPNj2fppXKg6BiX3BS9JBNXONSLaP3pg2rJ0K7bqgKh7HwJ
nYtaQ5m2y1hoo8glvSjn3pSeFNRwDD/SsctP6gszv5sLagct1E23lEu3MzXe
x17/AI5ZcEQinDKq27/Tnbm800YoNEgqrMKg+sKOwgZNlx0Ys1838A3mqYAe
I+rRskONprc814E53XJWTkWPuTr7IM8Sh8JT7AV8mPo/iATBJ6a4ybZXgmLA
lT4dAGVoRSVP/MBigpal3D5lQDCUcyWd7KLV4BRSts61ZHIXOF2f2HxSgdLN
1uLyhm+cQ8RSsdu7fdXGyYTyYD9e2FRYKN+eh4NAxTslqwSXTlGMr/wWzK/i
L9wdfe2TJK/rmq7zSORV5DKr+xSYlcHJa/a2IJ4QSPcFEDX8tWuDtInGcfAf
1EqJUVEskZdWE3jO7I270ZdNch7gb/c+tv/yHLzRyW9IJ1UmRESCtdBVD0lQ
hEnylSTcuqmgyKlw6w2QFjIWXYAxcnhPGvQbiXpguyeMPPjQDPqmr6IOqSAE
SbQnH4ROMk3fGYR+w2Z5P9cIypc0RruVnaWfzn9YwtHI6aMNIPTyqA+fzL8q
TDdQ35LG2IVFa2XKCi2GUG2bN0jJuXkuUOLU1VCttkvzOlMgxu3S9SqXLd7Y
mfGyOLgJdTI3C3RT88irGrFRpfM/kdBx83EtUgEhPLvy3Y3z8cQSr77MGxUH
EP79B7IIA8/q2knq2pvFLQpbrDOCvzcucbV0Xix8YCBjKfvPFuKxhgJSDZ+n
wUaZshcERfjkqLbUSSyfl6cMXfp526WpXtbtO8QnhR/UDuvyWB8fdb02gG9k
Pyw0Eev+SZq/33P+AkBKYnMakwUX6liQPHIF3ehCQTeG6BBPUjZ34pV+Cnp/
NFRkIqE43LcUV8v0uhp73hesB3x1C3ORTZdEg6qOrD1d4SBfvex9OpJ/6iEU
DCcEJqelhH5MuMttO2ayKoOeYtSOp8rOst+/gLR2aNzVibsck047BtAatpdR
2BXhtl5OBuTQuePJGceaMBcH9xCQPodFSgncFJVpS9dY6QhHaRr7i796Hw9M
2DIEqdXVvTQW1UJAT4YZebHFdLSQotRSYTW0jKicyfOhRDfgBcW2hl0dJEFN
PDEbai51JI8DcgawxX877ln7fDCxCW7NUCdJ8laxDqSUL6AyrPa70905c+3e
AZjgIvsfGZ9FMFnhdxKIECByqI5BH88pOOFUkGhwQyTP/gbVkC8JNF6Kl/mQ
IQ4e5WDCIqcpge73xx2AOa+9EhMc34DKkuCk+smnCg1Uf4lIbdrG2yXqePkR
YGW6n+QAGQ7RKxhvnSZmSrEKlNS8YgUHD2wUd7ALQGlkY2JZqKAMRaN6KTie
qIid8hqF1CJMD7sJhhL/7dE4CEwxapEM/J+2CxqD3IF/vyUqQwQxIdDk9OJ9
AhaVUpBRxg1G9QDEbnl27F2dA/aHQnmlmDkcn7/v5XyC9xO6hCGfG9ds6wHL
G5cN6do7uTy6AioLVHATRjI9C0pfMkSQIemaNmXlO7/KQDskz+wYUyMmpHtm
9DVRC+XaAa376yUxtOoFRp7MD+logQb+IjVo1+yKFpclJB8z06jTo9+shKoL
qQQaAsolsdsIPY8UWNksZPUKoMn55de8vpZAtTN5zanXcpg0h6Gk3KbyD0bD
x6h1qW1BKoZH72ODGvOk2rPYElF71I83e1AisFFpRzuZPf8CBr/DzKw7elP/
jGQ+f3M2G8kXEv70bv+3AQL75T1IT6KJ66o55tIp0AB7GZJcWCvVF9LTY+vD
og9BZIdne8CZBVeTgW38rd4cCQuV4gZyjkcYK2BYYRq8jvR3jk7uuu+x1UXm
ge2OoYQ9QhZmYHraWJYZC3V5SVmiRruE54D+PhFu7+N3BvedpKFXEbGVEyxj
C99GGcLJr+J2fjMEXOLhPUd5+DSfHxKaMTd1gGLkCXGjDApKKiSHkNrH3tVA
U7tqsa6MeUUJmhy4+K+ECGxvA2k4UDMdKX8YcYIGWBrjEXi57o9aosoKM8e9
g/vJKQ43E1T/SeUKzC0hymdYIG+H9OMO1jXu44JpTe7Kz2uThS1gayFMZghg
+U+0WpF34FBhk+MSWBsznPowT674cyR1GKhosAgN+Bxoke5QSI9jpzsMrfzr
eqt+juGjHApc6eG272IG/HN3sx8Tm7tRpEJSa+ZvaaW2TybeEJvJXKVtxfV6
kMFv44VWB+hB4BOseJTvwpbW2ynAtevj6K/sFLRCmLcQ88b0eolPq1kEUvyw
ZYbPU5VlmZDnQvaOwRCjO2qlf2DMS0N8ZVGIY+0+svMbUwqcxlAaGHMmZ52l
vVIeMcuB3U/8HGeVdU+4Js94ngS88/anIVQB2EYX6qVho/81+Y+LAZPLKnQ2
RbOIftEngcCavbZJaGfBvAhRLP3dG7m9RAf4YcUaTiPRvDpOPWL0qIZpdCI7
h44NxjRgJhWAcuYfO4Jv4aEtXs/utlPXUwj9NF0njrniX3aA9qX6QM//s9Am
5b+rfnhCwsooaqTkeHvdugdlewFFKlA8VU5gLDlxpJGhzfcilrnsqmUGN2NZ
wbScfe4HgrtB0Xqdpl0V7LOb32M5VGpyTBlUIO4c6GmMDgMyO5wJBbaelxxG
35Hk1l6fGLqAPiMolLV64VRYb7utXV34epYWMvByVbkuMM3fMvw/Vq0daQno
dx8CQTtuQMA3pGhod9hpEdTs3hH4FSQiaVXg6dbl9qzoz1LXI4WexHgFGUBF
sErRKhOOTbVEdfYVKnLR5KIjPoFgwipyM8rBc57u46F29e27wYgBIXOvJX7Z
FdopivS6CHgsU3LbHIUGNZVASEIT3TUlTevjfAdnt3WKah031fwDMI9QMguT
azfBESA6eLtg5DWBtg6DoGeeFAXkrc2IBlzQlVJ4+mrAdDRZ0FKUUzc97lU1
wKgkHiF3c03EJ0fX4tlelB54AUNNjy4KHlSo1dRZa6s65/X63p1k3sd+WleT
WM8TY8pvf5Xdb4Vst4+dZoh+U/qFzM0eVgrvXx5sDcyc0u+82qUSdRotZhT0
QzbYOKS2t+VVJaoIjuiy/cLSIjlnK72G8WvZJ/ctn9YYrwGE7a5U96zyRN+M
jt73oWqomMUGN6gmpLiVIqhdnTJwYyfS7TwONSpp1o6L1iK39VjxyH0KJrnR
c74OfRqwmJLZpJUwtkrbhseLd6B2Fby1EEFrBeVnEoHtKO29MmBo+P5whoc2
AyCbSBlGrPodb00vTMJPjrLIFqTG1/ivGIU00GkQ6OzIginnOrqniBrtiKX2
woV7G+HOB1rnxckrp0pcRn0tG8ecCyw6tg0XKo6E8pE+YMSH1sOrUMyp0Cou
tSBANOXzpOps31QKaNsegYsZPXYHhk4iiKya668mGM5S8gjgGc7wHfzi8CHN
W58QonWhVw23q6nKwGD+guFLTyDt4dBM62GbMCU+sx8+2PEZNVENUSUnN4hP
TBMx098fwubUeyBKrBj+6bsKwEkjuVyYuTZvbjUHhox9aOsJt3MEhFFrnU9u
C27+7Ws6fL/i7g6i67fClYt/AIOdIkbKXbulF3gX/DzwMl8TXzxfLYxXg6OD
4aWUBqofzisCxdqa6yRUDZJc5IjLuVhDQk8f/L8xXklynTbLzlwZDZQClDAG
QnL0AYUBDewOvCUeEkcPICgsXqm0PENvoWWqfmDVvvMo8c06iGCGJ+KvfbLo
nUwBgQLrM+9hMnf1LeSPYAnr4lCDj6cWoP+W6TU9psFGsftsMrXMowHJqJ4+
qxZFY4lEVjapaNktgA4b+fjJ+c4HWJVVcmdxP5+oA01RV/viNqbKpycX1vJL
E+AYZ9Ia6lF/P7zWx3aQSzy29Me/61H9syv/Yl2YccrDbm1NhqoCIopca82E
6PgqNvbFzFewnxXE0tyngeT0t8K8t5rWYBPZ9Xaov59HVmLE99PGQvHnJwB9
wo7mXU26SXsz/k9RM2d19FxKvXyPJHndRREcWu6AfOS5z/CH9gmMzlFWIrny
woiWQZZOtjMEiLyMpnJV8YGmlJ0DRKUyIq0GVuk4B1af66pXl0UpshMUslUK
eh6qME4EWXn60arJ5vEjz6fcZjh+0mAX9Yo13U9ixfbZ85EkWq999avJjMiF
Y+A3MUCsBGBnm9s6OZxonBnKL03cmYogx3WbNdFC9xyFldv+nCtMXxG8WyO6
gdJF3s1owHZDhOZDCp3NQ8n0AXEeM7HIfKYmw9G+6qZ1OeIeIKJHuoMrt4Us
v4dTz1Abf5Zz9H/0mxLzh74k7Dpka2hIPjF8YId8/jkKmTJInJdhgvS68Lfm
oFtaSiTQz+TRLwYYvIojJe2wYtFq8U+dNx3whpEqZz2cHmm2T9mFwidPjO4y
YF9O1SFRUn8nMZuMPfXghupPm4gYYowmFV1Em1aOIldQe3OPFIyaodfgIp9T
AzNOIS+Ojn9iTuttGLLO5nxxoPqEob0Pe1vFl15UCYofdDYPofPsQJ/H6pYc
iiEnmFAlOIl4kR7ZPS9PW70dCRLUdSBCrxRg/TDUJm7a8YJnIzAxYwRQJi3v
BydaG3htEvUUDddoSniq0yorMYSmQcYNvf+k6QaN54vO8HhuBt9tkk/110L0
CE7w0q46w8ZtOaB/COadcAnu9JKfuijM9gJYLCOuK8/KePAEpjKXhpNTIPGI
1DJcRgbjzQfhz8zsZcy2wu2AmtdMLhYqs18IjM8pLXauc/XqhRVra0zPAvsW
VOuGyZ6zxXui+3O2+MvRNQe/S87+tENR06gXI2p+VXpEPNwnFtTgrLC2ADsn
156W6bOYyaE7CXZ9qdN+A8wO7NjgnKAXF5mU5wm0D5CWlyyP9hXIqq2QHA/i
MtIi3nav593IvIBKMSXnRDM9fI9T7g0VWoRwO1D6iW6o9ng4OhRbA3IReEI9
2Q4XyfkTssEu57xssjhmA4yHUbgvL0YlEr9gDcIyzhhwfz3kzYJhX2fuUcj2
aVARFacsy/7obppFQv+XeZr+51bfSNor9JuO+KdDMKudF+Z6NhAZHHJVUlBy
tsBUMb8MGhRb61r7KbqumgU6PqaHsZmvKHjUnIbfoahyON2okKLykisR7aQY
G8t2nEQfQvdNBXov3lXk2Xd1hFehcwT74lWbTue7vsO4UpuibV3ruCuJ1TOi
7KpWYt5iMHez/Bx48oFc9SdJfy09kY/JtfvvZEtTOGg7NFLP1gwD+hBNKkQq
vE7EiircEoRO7lkUNS0uIPemAoR0jHQa2aCemYs5vm1yq6xjc4FN5rRLIe1o
Rzf0J4v755+lcxa90GYD28tWZxBeXJpct/spoPNKjCY9SmPTg89g0kdOjFgc
vBfQRxSEe43B2B9ZPfFB4H2NMq+HWSTLDXgVfwXOTdzjwZg/OzoSffDsj5ri
LCmA8waWboraXfM/Ma2NefdVK391YGV0MRaWp4ghKW7C2R0vtHxxXNxnw6H7
8TXCWbwDg3fK9g0fUDPNEWi30pFPOg5toiqic3us9+yS+SMtcAu5Q/xURWH0
bTTFHaxlRegMil+sW4LcF6+9V/rltyS8rhk8Ed/LHLujs+Aroi74nJskKe2e
v+D4vlnMDRz6UYiz3efSDwEAZiqphf/y3IK99IOMOjtG5n+Im1pErSeKoVre
/eOI+VSmrD+KTsFqZfdVwlc1DwOdQYUwxR0ryeaavLtytP6L19t05cRi1rL3
2vyrTdEY0YyMQSf4elpDLBsACcdJK1i40sVsFqjIqdU4QzjwFt4POPmRGE5w
OqAWDIkWC4WP3H9e+DQMs7YE141sFflBl7oKg1N9jqbHeuetUsGlzQ8wcF3G
gLemEs6+pZ/bAr96iGcMBmJHvUfjjVZIMlmIJ+Bwy67MFoNYPJM4q/idL7Ka
DbPbsJVMENkm+g303Zoxb8t2PdcusAQ8ir0Fl3HsYIOJS79A+Ormr6BeUZIB
R4DNrEqnaqm45WFl2YtPqyIaZNI7I5PDtYF7RBoAScqOhSuPaDSHRewBu5wv
dOeAMJfVb8I/8uHH6fzjYfsXGU1V+w+0AcD5+WaqljYHlyDGsky6h1EEUdoF
AsIFOGU1YF4RMuhJymjLj7qvUuhVXEWKqiNG3OxQI63cXzK8lxYpcL5iwPzU
68MXaVE+sh+IDJ6KVphMKRF1bA45bmesOEkqtX9SCckSrXNIYL9s3/1zwnNP
pS2uozQvPSMTETd2zi+7bJRsm4SGGMjZjJ7TxInGwl0s4fI4KJL/2R803CFG
PiYD2hH9UZZEiIPOgCfJoIuwP7mZccl6AlOm+W/Td8PDr5uBhHseoic/xFw/
SVETtj34cvOg6tqpJzyB6qZAGBGli83mzuKoRcQ6n5OQapHrXSoOa2yriH9L
ayOQlWiIdGiSQTQuzbOJUjWhSUqZyM77CtH2eIBUg8sUqqzoRV5nmNG2nemZ
/mKkxUyOY3cCBeWKMDG5VL4cTaXAADCMOmSO7zMS5+l9yYAYKKMhro0vwNix
U1m/NYqvHTvJGjdEe/bAqKp+CbUfSZKVgimNnpKFD4+47mUt6swUB0AYDkiO
HUG9vLVZGJYi+BTNHaO2ntv5xjsaea/Pf5Oxr8XStvJ5LY3oUbUvwakRdSTM
kpSKZubYoCtblMHL3/jSmSCKovWBrZt/hwyTCChFqUSRm+wJAKv/+0pdD4ne
0+vKQETxHJzOrXW7cWu+De2wwg/fghjFIXworU/P4mI/PcIZeWGeBtJ8xYV4
K/OfGESb8IxUnqXU8aM+magiLONQcJoD2yPhABx3e1iN5/I3YzA101TWJmeo
KqNMqz5Myk27R6S6LvgvFQISpBrVfOJoIkZRoyJqsU0qNieAN6g3S/n1PkKK
F/CvBV6Z6Hms0ued/nTzsVtWItE9DME7V2ec8wQ4pT1FV9VRepNne6PxBr12
x3tenm8Pq/wxxVJ6ZGWbxlL01fKgsTT0kewkIx3uRPbOg1nJZE+aOaSjwFWH
R5k0Q8IrywaBFcfm0xHZuCOKDJ5/7/pBYhUXRDP/vyM4mosHq80LwTNf1q/p
MlKbTmie/nrc/gOhd1wzaMi1sNezY7T9HdxNh3xsnOiRcIagXrPd3BooeNLp
o2H9JQnyK5KEDowk1O1ly062WfXWISXPD4RzzS9wGPsLeFxqcbup4xbF7xAM
neBJpS5P4UhqiUbfjFCuglBObpeQXXXX+Aw1MQgkafU3Now7OgMBP+/SckhD
YPsT6cPogQkrRGrE1Se2H2jLQLmNN8Wyfm3QHHgZxa7zgvlRKBDFSX/nan5K
wJhxVVds5Pt+62nbj8NV4oGQJnFHgkWFBbcccdwVdHfBaGOEST/bJA7V9Xi6
e/jGYvmKSALSmmjKZtb0tqpPbY02PjE7VZ3t6v5mxRN5CajVc8KMYgaZ1p6e
efwmliSwXcXz7/sidCqVyDRitMC3V9/g2V1S9bTwR5MvToisn0eLb1Pe0X1/
Uy0F97gFPIXjUdQ2W+sdXdShW21Nfd+UV3BTd8nrfckjSV94Zaf6H7TCpiEO
wOik9avVFp2pqb37XHWLLPsYSkX0XlJk+n6dwFpGRHYowBcFTxQBn33zKfUF
FP5H0mw6kYzwg9k45t27PWdzkCUygPuOeB3KgjwKY2SbYpB6HbdY2ZwoNtMs
egD0e7dpfZ9+8p4aaz/qLs2IT2fGQYeKZ7f+uteK/r9z/Op/RedVEC0extRJ
VO9eNZnWXt0UNrM1G500IB0X3wuNO4FeM3aJkqMOGyoiF2LOWasQhmFx+ywq
1z0inPhX4etAO6e9zg7nI74zAFMsD4dxpurHpNBTLNDWp1Cqkd9ljDddiuq5
Pcgzl5Qru3/Yb8nDazeDfOF4q5YL0r2pBKHU6ZEvrrDBnHCtDSqofZmdNfun
33f8JgstZcDJ2XFsfJJPycrk4T3fHGcfOwy8DdFcs/Hb7E0x+hIFtcTlFYlC
GAMOZK+dyEjV79HwcnzTWAVknpu6Pofv/8jw8Zy1JHI7xEahaE/I9HnJlkHc
wFVaRbipr1frbYhbR9yYr6r3I6zQXlw5ywUkrOR0LEL85ZfDjZT5C6cYWMvd
Bm7iVYtNYYybKh6kSjp6AeB2l2BuFzzZlwc9JgQPlnLcszJmpXt3KRBtNXdQ
o/a8E0MQJrBHo6M1G5CbECy9USnk336PXR6LW5s28DZPhPhehEK1+7URm1t9
Q1FIBxlutIQL7IdfZ39D93MDq97L4ub1iclK5RDXXAr4sIsAv1zW8fblCNcg
86UrlCP9kuwCCjs9311HzJIFrU11c0Ev5oifCQSC3vJAwBCI0eJayVR9V0v3
VQWlvufsZZHvCheXpjMzLbjfvjFCjeIwk+3hv/g3i0XUF/INTRvfC5X1ZMrc
tLO1UnRu+Q5qm/RvXCk64/ZqYIl1h6hAACrRwn3QYAUkaUECkrKajPX5HrI6
be0u+qOCPv6zPPTsQ/kD8hykgj+RnHcRtXLGger7LhLEivC0EKI0doPnpiH5
hjp79cU++t+AE1iAeuhcogq4jBMsZASJ7O/ott8Z4/Yy1zGHXv8mCLKQbImm
YxdRckAy55kX8TeGQ6IIkCs/C9zuXJligz+b+/f35qr+e21/uVoofFFpds+R
KWFRIOCHDefFSQW1Dv/OPkDmXLhzQbUmVVoaWFIZz0C6s0iVslHT4vUQYeio
gSrrKj02LoCJjfF/4+5Qo/r3HCudZaaOOmFlQT1eZ9WQZitrOq844hOG8r3A
Z4QgfBU03cyygsKewWkobwyuqm4NQYm1hNiNMFXZlpW8128j3gubIuIKidQV
WCtmqtlbsbXPp/7GzaMO84mSAxyQ63nLhT/tlI96VHlJAEyC9FnYDVc7a7HM
DnyRTuQn6bOLB1vo0ULjFS8GC60svnfdfEHEBV43N83uC3x0xzX5X36w1wuk
AJ+p8+rrWSw6/rIo7OuQgvWePcsXkljVDSC0jz1mqzD5RsgpAh3we33JaMXT
Nx+wteUm0u2WAffKEGha7mFBalcLlQEtZCzZFGfUbB1dI0RXy7pjRQKjvHu0
wTh68fYYIlLUbJjC1yeQIjzqrEVcqEKh5SEd6qhj8UM+eA/WyBkh3+ZHcuX8
/aqsPAgLZBBoXBlwN63nkya/w+ClHDjNHkuXfxJzx11a9HddsUI0UXoX3kRH
DtuToM/uy048I+s5UdXfqgRaCWihC9CZqsWdJpZt2E809gybOaD4pDfoy3B4
dH7EonzBojk+ex2AO1Xut8hvh/ar/ZUByih0K1qYzpII3/C/eVGDkLsKajk7
acdRFMccHl7+6wFN2aFUysf8N3ajl/sfoLaeF9JtmO2yjIbFDtEJky5mlKVf
LQ98PMSuSEmxp/u0O7oXGOA2BPDOJ7UQo98+dBTg31O4g8NKmRG/gifi/AoD
LihCAcPx0xEU7DO94ykAKi33IlnxUipU/ASryzHhVwXElAcBr55yPnFPkcjK
ERVCcaFIctTUOLV/J+uqxSxN7dOL1YoFLw+VOssVFZIRst502XIlBXcQzm29
qIyEc9EOYXAQMEJHCjvf/n+xrUe7waVdX83kxnbqwtVlbd0ZFhg9+3vvEQco
Zim3Ioyurw161A8G4fEl3++38RZTCj0inuIGwGJkmE5UApp4WtZUrwVJLY42
Otlc344ARXlRCpIk2i+yDUo3sfItPVbLT07ZnMXGCHOrg4l11gpYv7sN70GZ
7J/ylVKb9fvvLsCmK3FWOkrc6njMrqywh5mpoo2swubi4xs9cNz180wzfp3W
vwyDLhUnVbHdfqBUU4wG17swjpl5nDoN8gmu8OI7oWBQxI2heSoROCg34aZG
yU0D3xBHzt5hBY1NFxkq3nyLBWDWz4e7iMwKcHGQaeRhY2CgPtINALwkR6le
3btMZAmEwZ6t/lmRWjBqIeW9BjsXc4pHV4jYA3D4E5SIfchodGuwMXlbo9uJ
mL8zfvyFYSNMrrM9VuU1fLh87SFeYRc/NYwWB70+rM/mwMF9QFZ2cFCwdiIt
cjgQDZ+0NdM+xMgCcs7i19D9N6aROG3H3Fz0Mp/cziHxSHx2/SXRycn+osvN
wdHJJT7JseRgU7B0MxgRbf45ZK2NxZaDVAHxh9EdpQyx1uAkY6aLzArUfZ4a
aTCdOCfBSwM72dGgLCuSvLm90tzR8MrHz2YUA5Ch3qUG8U78T7C7q1DSFXAV
FiFUZ1l22sgp/DK9faYfXgr3nYNj5RM0rRgyJkEesbn/nUXHXYC75uqV68CS
I8FFvn+yBwaOTd9s9mD/eq+lDyzmgjaLxuZ9RFFxcKKiYXLygj19hHhx8rJf
x3YcSGPNy+LzUeRgPfBbTush+oxk2yFS9ixPFtj3lTQEnuCLVC3ztS8UVy+w
H0kj+87Qw2Dq7Od1QJCTa/ox8H3HLFQQ+CMq+kVDFCFPVG89fm/YSOU4ftiA
HsyVJ2XGwWCA/q1ombE89py9cIb54yoiVwE9QlvMyWefqmXb2snk1PhBaJf+
fb88RPLMFr8Hdy197nEIekaK/RGrt7xXVzauPmjsqa04RR2QqyWoSUGEBG19
sbqHshodcV3HlOx4NS4QTbfSLL+kCVIp/f98k4/0DOHpEeJnFPAbuGAht4j1
qki8N1mSv3ncNeyvXLAZuYY39NgqwhedGprWw/AtfeMRq6EykZPxtg1q9LFe
Ibhi3NmUoInFatJYp8IoEFuatFxfyUtT8r1VNNtRUz2spPeeCseqj9q8vbQt
sGGss/3xrKB2eC1BBPHmL+JG8btNbjbCiFLx14uIQNSa79bgk1Y5wimB5Pr+
LX0EM/Jn9FkVdzaBMEyjA3Z75r9rX2rWVz5Z/9VinkNhyjVDpAAf9fJwcNTY
MvmYx233aV41MEBfeUEHp9fQxHVd9+ZApTR5F/9bjrnHaDD9GUQ3vNsDxkEl
XkVijaE7WpVuqeQkV5G1zX7cbIREt9r8PMQ2a8g0jVCBttY/DxH3TLqrujKa
Unc+4Rwk8/dIRdaiJykg5IS6+2CDA6FNHUmhwO9lZvyIbJ28gdSmqvcdx8N4
tmsUxuDKV4oiRsToWoMlzbDSGXI0pAcyys5i/IrThfgNQjELFcGgq5EvLCS3
UZWwhCzqsyEA7z0o2kAOtIw9967JcqeqnayTeTtJ1bXTto9TbNdKDjVZpuLt
PgumtNjZoamEfTc9nmTwJyHVt5mKfTP10vGUbAgc1HuVvrdBwid9THTKlxMe
hy+J8My/ppg8Nt4R4Z7vKg1jkXRJJoIdGDROgqkCDLAUCRe+o7sEzVINQVZF
HkLzO5Omw0lzQNIUCqfFPsI8SxpxPBE9up8qBXrujlO9x/wnBNuI5BoL6lzz
dLMJ5AimgwFuVaI3P8IkEIDAeppg15U4SOo3sDskGiQJPlQEC0qyPlOzGQxV
xJso6S/IFpG3kMNwyU9FrpJzBhh9ywuo+77+Nle823sv2AQSyEfjPJcltW7K
f0gYF5RIYC6YfQf7dQKlnyo0YYEgOvlC3tYdZUc8/5sAX/oXV1xQc3P5N92F
AP+d6vyqkBQ/h/DuBFui/lRJE8XpTET6VDFtoLBjI0227+PR9S3ZhAlbukL5
PFJNP5KlJ+aiEtjgni1p8RKsb3x+CVLFV5+uy3KvAYidHXu0ypoDmQF0aooE
h2yu3v+knn7++N6N7p69d4lN3kNZIOp7ciBa0ysLDVnbv5vD8vkUdbtikrvg
PGZ83A8b1MMb/S98GKPMEAa3G2btaXYZB0C7q+zhagRbwOsYit8XEAE5c7KB
gzujZL5bFrnavIKVNlhhoHG939tSZaawi6nxTi6yZI39mspAutOYBAT3GDXI
SWaF0hLcpxjIRKn/cLvSdmfWBYrHZ5tZD3Ckjcun9YH9AyOynE5otq/bCkiT
hdEGBThm3qpmhdnhXsY2NJxuAF/WDHkRItdKNKrJ68k/GnH0qc23TJsBUTYO
x2YnUIx19qYRhGgNZAd6z1Q1UbwW3pPItZVr232cZl/Ml48HSrix4Kb+s9FQ
F08pX/jV1LNZpJtMjAxHE8vR4XIcWqSr9SILvIzXpA1Nb4syyrW5RVb6TDtm
PgEflj1oxOPZPusGU2jubAtYbI/rZ8U/LRZwJ6DvvUgIIthE+bkTZo4mswtW
ZUEIP6GEoFxje7G+GQpbgZrv2MXkWp6n6IbeAa6q/sMPXp12gXO5XRI11Ppz
hIyapdGw2+uTt4szSdByt048B9zsWa+wQoxhnfUJwz3B94KH7G6dSlx+nMzT
2Wc7TJZ1Pt0EIO/dDJa9oaDFBaANtrBM8kcgs5EvJHGskwlML7+5i3H5f1vb
EvSNQW4gl/e4Al1abVfuUntHl/NcD4hlDh+vCnushxkJyapMGW/6LyzxF1FB
MQgcf7ZGEPFMAsmCnRH8qJ9xxA120Z7S4d+wBU5eVyX5lA2YNdsFLa5fLfmA
ipEpwrJc16aSXH0B70RPpR9JVlNMGdwR8ZWX98jdU9o4ftDRVGbgBvozDlkd
iS0trFrBD3/2jFc9kkGVvubDO4Dqy6kUwcOoGcn6DA5XPFAoGvHMpD4KsWMp
rtgrsEK0A1FH5/p3s4T6dKWrOhIe9ew16yaZMTKa9iEkMjMoYzw9qxUqaOX8
3m5TInhcjVUErYtvEs5PU6XhzgzTMw4lFc4aKBLwbNHf9QRd72Tjv5Z0wLqt
8ofKXkAyZSV/gCNb3S1rU0JPiezUV9nSjACLPRH0OZT9z2mDgpJrIjctegRs
4zNoa/qSGlI3u8Y3j9cX1NwgfmzTRTKyOaAYRLmKlKQ6LIjcRpL8QuAJcQr8
SFPu4KB4aK93grAahhYHn1fYStXD7wQ5a0o5GrIbnmDat5VbT9QMaqZVPMmB
yv2vaDOJzvPOP/hOOv9jPLy6STwl9573W/70lO4KFnMAbx4lY4wY/Goo0PWY
WEPbCkgBswY3e2YU8ttG1GWOH7eRtXSWRFAFWlZ5qveKnoQ5VcYwoHfA/MJd
0eHt8LkjTFmroe1pF9XAebte2EqgWtwBnTbDbqd8HJ2hZVTIQvYp+rQZ6ieg
RTQAs1XyPjnOd5oBVRwKe0FWxvx2g0IGVsjyUjnRo8G2uLU6k20Jvg5fZwQq
CB0+5EDTN619ESCUEtwix1CzY3q0tSoSHRuEqmGSiENnTd8jltKZPeeyCO2x
PLTcXR1HO9uxW11JNtJE+8Xq1kWpYXUq+7WM/NPGkFdlW11cYzDj442ZzzYb
ncQOyKjrH6AvVrhzpJNyRpiC0RxdcSxDLp8fiv6BsuzsppXfdozprZ3CsusG
j2xQpwJgSNyWpvqC+3L77nk8ra2jR0qatwntKQ04TVG3LNrT7LCrsclr9Muq
n4/XjwxA4whTRNj1Yjbkd0jkLrD+Hm0n6INiwe0FoQ8VHs95G0zj8YN9h0bN
noPqBrNcqyZwahXRuiB1dU6ZEqthlDlQsR5c+q+9QTeBk3xxQp1Xb9Qw9Rd7
Ya/Bn1rnkEtUi+PrjP+DQjMjY+XFPMX+tx56KHqBcTXyKo4IllujXDI0gbNh
4Sju0l4fz8ZtXWuoUA1ObSMuZ6pVM5adhNcoKvoHxg8LNOmhrqBffO93qgjV
dJmsloGRyXcWuigr9Jygr3LrN+zkR6iMDeuAG5+1FD9d/xXgdiFY3FyihuFA
YKShzQdh0W4ofcwcLNlI2ZbM4ZIHsRUsXoefQCZGF1lFbJs9rAkl29NQdxtA
ZevgysI34DCre8h6QTNwRr9RLn1Yi5k+8Fd2TgbYZYB/jBC82/ayTuOYy4R2
o/5iuiicmyCE6KjiBS8MThBymZsW8seWZXGx/ZeluEmOjsY6MZ1/hoUuEp/V
niYImGiJ+2iZWhgQvakESpY98JawAvOagBj4dwqNjyaUegLoCQ6TF8KMl2Jx
5WBDEvwrhk0S2YTnNl+EQagLpcJLAElCCj2XFV57dlLBrU8lM0PZQa0VJeSy
mIFPanmQMzoq+Uf42CHAURbfNpsQHm4JElb3mK2tlKXcbsECKdn0nh+dGHN6
uI6FeQW5B8uIvuOr03i987CZ+DA9DsF1tT4LdGy7KM8o//SbAFNzSbAkdCiT
SRgqJ0OCPWZ8mfPcj4/v2xSjoqDv7i+PmQTdAOtNvo5UInvK3HN2vGpuSjnW
NZz8OjpIlZmDftVEZJ7OKzDIXZhex2fNFyizsj9cIXZmbUF0AbVeCGg1IDyf
luTaaV0BnN/de12deOAjLNqbIleKO8c3ur1Q7tHIA1+ArxxzRUrZN+uMa79o
LpQU1RENjbVunOyag1ZkSwtCOJ7QKn8ArrgcMFCqZRhfJjP0qIYdJFWfiRwh
ZMoOpi2ZAZa1c4e6QpJX3J9DmgL6v8sczXFLFnHqymoj+6eJw1H8YZ3u4tvf
i67lXMgs3GJVL8Nbx/dih8AhNAvsKfXY1cIX+d5wBICvcrFQ1dvb7ugPOxPC
a/PonMlH94+4vPBU0pXYfxcfYGnW82rmpBcmVRpagnVhSyPkKbptEiBOa+VN
jYk7frVD2gCFAhyUk4rHou3cjbddbQ7Nq9PdLnyXzz3W1XKfRTJmvOXDkoT/
gBtABDuV5zzNAEAcujXGozzuzm0aiZ3HpvoM5He5FLoDiPUtp0nq4yqn7gWK
jysC1jhF8x23gltF9hJ4WfZcrNB5zrXEhkZtMSafoScI3rZYCafkuauHAOcB
wy901KU+kKauNh1+5a/pGx798Y8WuGPoOuUaSV8bk/vC1FXVTKHYiQdHS/y3
o5EjM30iTYVS452jyvWuNF4QkrQvoGkRfZ5ixlraMpQ2sC65lAfZi2fQQf7b
0a4AG9GUUx+y9vTjilhnb8vqzaIXejm0ghjijlC0qwmYuH3mJG028NL0EkfE
OO/7mKGwK8Omj3Dvuw5W8Qwn2eSenE6vObm9PKnLZnV6IIs9kFWKDM9MNgut
RffM3xOJFZo78ZYXL6QBw2vKmhzxOgcA+yR//6XAepaZi3Emw3/0W7Upu5n7
LU4J84gcX2pbEhYMuTgNzFzlldHkO+B44BvHbBvyOdABSTSyikcI7nzJJ+dh
32wjSPadZoTGNKYBJbquiGrB9xkUWjOG5P61XLntLKA0vV+9ZHYW/hFFCorm
45y8yNu6Fmab+Uy2UvmvEZiYKDbjrqOLZzkfPyEsdWUhVaUfadOUR8mNgQDr
V8ODz3qqeQnztbwAcG/u9VF6DuTKJzlhBha3R6lI1TDPr243pL4Qtkcrb0+A
QBlPMOwCXYSymDyOktITsXmf36U8tyHsQIDqyRMKSijoOc/YNdmrxGalSfEG
H0XkzBnKl6Kv1dr0Ex4sUxrMoFv89mwcFldfS2H7kOHcgqJZEF6w5cmJ3Fxi
BGVATPg2BuRn9cFFEWysATRQIT9hffYsNrzocPzbTG38ym+sA6sthUV8DNdA
qPfC/thE48n1TzorKh9L+1VAjq6DSammz335poCcAKCKbz1ijQz3Lr0BRXUv
s9YWmsZVnuyRPGMXxBmjnP/UqEaKPn/9RVXJlt8XB0knH7JOyaj4J1TwnJoB
aoOQDoZRfuhOSDaVAF1aYUOgsWlICxz5GISfW3tmc/LHYc0jtWjB0w3AYlL1
J54NJurRECKXFz3DAB/QWM1r6UoMqclT/VrYmFn/KsEom6vWqnlZX82dQ8hN
42eame3adI8tq0BPmNNhAp/7EcPkpxpOEcsFr12JcCkaDeeikYezj+5CFRqy
CUfI2KJ6BRLSUJ69+83b6VbK7chFEkiS9DPKn2kYhH1vnCIsjv0pHVRnQgz7
c1ZkjQhCEJCdLneak4YvG0jdqTU5yhlZ9hsT5NsOFsswtqx1xtGOYEGzw0rl
XNhtQaOZOdOJEe0+vEQWzSlTIa4Ijl8kiB5wL/WY9b9Yr5ZZWvra6Z4bDNNl
6BjbCOHjAnvMpcIzR/iL+zdTEirkwsDWfYXzMkC0RaJXgZGcrKwHVIAUf0ZX
efBrdalotmqKzq26ZChq0g3gD7PpdDBgg/UCNbjDc16gfEKHjGUj5hrdKcRq
ihCI7anW8Mo0jibWoP4BUWXGGamTJc3ycMY53Pa7QYXYVDtLPUMjYA8/7Iuf
N/0DJBUwXbbRYxfVAJTLnTvCAhh6dp+3geW7oV+eljy3sgWmctK7PqIx2vHZ
kCNiWOjjzc+8iR8yrES4GOhSA16tRO7SsUCowMdnV2lQuuIaVe9ZgXTnqdfY
QnzFw2LW/0IrW/CxQIAhQAOtg5k2EVI/sn/HZtLfzHhPGfMepHI5pd5ZC43d
nNuli7A32I1EsK56bIB4ESwwyGvva+ct8UxEyQo5aZLdi98wJ0v2Zs9T5tLF
DQ/wRGC31iRXFO8Jl4PFMkkxaLEBn/vJISETaPPYMD7V7l0YHQG6JDowfc51
2wJNtlkZvhVvK9mr3YZbft9/y4k+7lMKKsXAHCHHrKaHdgcwkus7DZuojJ50
xC2i5VfDyHnGNDpCwov6uC/Hkf42TMKIiVFvwm+22d/CZJ69HZAunFiWcw4d
Fv0zull/1dpAbEgeGttBeMf4lzuIUuuKSR6n/0mF9r7voGiOFNfXaJ+nJBx4
beA+Pvw8VI2R/Y/I536HgVYFHvE12LKYg74I8rlXVcgBavxUk2opN4R2DELF
FPWPoA/58iwkc1rU8e2vmYzzVflQPQGPF0EVtIuKoGINb5L/h5skc8mZMSbr
QYaD3JymLSndvA3oW/U4bGgMJDYC8He+ioDLvobyGfK2fP46fe2KPjl+jRbv
oYfgt1HNoi/zQMia+mmpxxfPYkfX+LPM0EAQb3YIs/I2NrEIxbpX8YPNzWxX
cTLJ5WfvI0/aPGoLHfjbh1BfQ8bVSxcy1xSerP/Gv3yOvWo6hO1WZaPB/9lA
8HZgFgsWUWw+ySwLkm3N9rhtZNUbwbeVCKNK3AN/vowcTT5m4+lVjIG1JfoD
0PnYRpQe8yHHjabxGB25/aU5QTeb+/psxjvYfQvm34a4lLUqKkQx+DyP4xyh
ZPSZ7HJ3qovP3b6hMlw6kppbu8tDEjxkI/w+roOSQtgCqI9FWWz/asyu3cZp
P/03o7/e21iQX+dVT+KBTjCfliwffK36zfKwP3xwxqJjfRUba50TAkEbCmO+
FYl38yNJIHgbib8y9Nn0GSI9IeH1L2TX8MJrDalky7CmGZMm6kZzqW0dPSHM
cv02tC62NBaUWDX9d85ILJUKRYMgFd3A2c2HSSdKBzeumyreuzxkUw0wUFwA
mhlTGqQQytcGmE7W8TYOQ2ZwHT/4BnEIg7Rn8lijkl6zvexnUFT3dBkUPuoy
vHw5z1PcOIOIFJ5/yofxxWbsW9fiuHSm62b4DGiKy5UIW2D0mDyY787PQ4m/
W6ubccXO3EZ8BrzBmcyKWbPWonlJA+j9cY+M/g0hMX2GQuucutPAkUczZwVl
Xnj4ijBeJAWaWR1GwdEVI4kKoL5bhy6Yt1TiGmpwMZ6ZSOc2Y0ySov/t0afW
+KRZMULFDXYLmtCmiNRcVUtR00PLDRFR8/I5AUKfDvwvUnI6HepuLkprmA5x
tJ31ty1xdRVZVTZMHPIy93wIzA6IH3NeS3G6qVsFFuAEtFJH9sUKLVkJi+gI
G5uVGfUPCrTkKdZ4SBe68UH64lJ3AuzeIbDltHdZnCsIFdkEHoPjUrOUkHQ5
++Jsmks+pzhdz+v3Z8SZyzW0ZeKyOGmsiAMi4r5ihcabaJ+3zAKqqgO7FSRq
fcX/rz8paSGRxAitBH/rYPDKtcfgE+Jive2XmftAVeRM4lP7iBSUkSqkZfCU
bCemQLyvmgVgL2VpGfNYPZ2Agc3wN12QfkiQvvx66aguJdJysIyWHzBvbtH3
gUoJRkhgAeK39sbBVZGL26xPPZ/iX6C685q8IIGo9GsRaNSEb3V51ISdpwiw
tASO1cOjqBlRiYXoLbqd/qGGt0K0flMfXqEkUwqZMlKquX2GasJ975kc9nBG
4luXwHQon5D4Rrc/M6gtSdJFi799ltEsegiGc6NSWBtRbd8SKpxb/Yv2iobX
Wvl9Zq7y/Cwh9HAu8pfLE09JEnWrZiFDeik02/hNBX+48bC2ovAiLut9egT4
lzrDN72J3TyaPIEnkZhcMtxYJpPS3xNJvv/3XfbkJDj8ubXN5NZWhQIwWmUC
bz8IV/xlvo9EY4d/B7dv5xi2N88ZEr2lkJRIbVWGLuSxyEDhTGmueoB4ZLWu
2LYXKyRFO+l/OS1ObK8DnlBAtYb+z6yAzlltKXZrbqKX30FA2jOG8Ir27xaC
yF1aj2fL7BIlB4wtikiJAlE1Mw98D6XEPVtsUMpbjj4B6m3U4cg96FBWq5ZD
MWo12DVkv+E1p+Rx8GNIOVHaysHj9a6K3dlXYlP+lPdUPiePv1OZADSAu8Ed
2Fd8kpbCzNVJxT34YifLIiPVYbwkpYPh0+grlLeWNJrbhGWihtvIlIb1On0D
pS1CZSyhvhQm1h/YoKDg+hWnnkn1KN9TTMVqrrAMOZ7s9XJ9BjQlm2Pisn0Z
xy0UMBF070MnkqS/8/rJ59uDUf5j26YWVYDE/721zJTB6vCzKW+CkvK8v6x0
Qi2A93q/xoiW+BCsb5veZcfnejKXOkGyA6SplaTGQCV60uKJ0v0V0wl9z7cB
jaV/JUEkPHEzryf4liTszxrzWq05x2iBaddfnJ1QTxJEsKzwyvVVqd/L6+B8
B+hmx+47j/EaqiX1FJ79hffgQEtBnZS4eSfCgJhDbhri7CaG4kLJ0O52zrlt
59wYk82Crw0AIMr75iOLMyoeclkcG9gyBSFUR/8aDy8qKTgq9GYFMdXMxFW6
+r44pAnXy/++hfHq3l4n/uEQzd9/1xleVp4lxz/HrXsV+7GsRc0xWEWPEN1d
k1muK/ZX+TS/WxJIkffqh6by4tQmn3r1BcQCZALmf7CIMFA+6FdducYdJg1T
IxrK49RYapzdjGBUl7G8OPi70gWiu8fKLzloMiYu5tXqspPza8x7sFXZezmk
shcT0fI8lVAILHliHsxEnseZpuuKPmS/0scLsWXC8OQ5fSJcBnh2BAJlkQWO
fWTDGscehMT3VKV73Ec51bNbSMokJxbe++BFB7v/h5wB8ZOKKdmbWBy1nf8v
6KewJmhsIIzFLG0vs7oX2ZIJkGvoBIau1ij7CLuXf/NaXreW+r72f8GSb93X
h+Z+JmDAXIGxE8ZcPX4vXGpEJQ61dCe2imAIV7cr0eK25KTNSAEZ1oGmbUQ/
ypvXmlBrgW9LnZFnMT58Fjyo/MvyeOGLdXkqREFUFjOSlDGqm/I0H3QjGhG1
pjxtbwuWb9mqbFe+dxjAGAouijBbmvQM547YvJtTCt90VbsZ+MR4OycTYcjr
jbvIVzj91HsnVsbhBm4c/uFXTNrh0xbE9R7QMe+9IBb7jdbfTgr/xo1KYP33
NHCXan/7K8tofk4WLWIN3kgQdfr8jo9D2VhKxzSNYaAmbfl4mcy13VE0QQtx
zioHwMEmZrf5o1rXiuE9WeWfhJWHpTaubOK1YYde1LnYD5e1zAZ4DwAYG9E5
n0HcodWuz3AzZzvmYUUTM+KbmZg6McsmoU/xJKlyqcQmj1z6RAFwIuBE6PLC
WkVIw1L8pJOtKOnkxmpEwC4FvnLxohezBVs/tjfLjUlRaoXNQAM1xgvECm/I
F5ouQG5k4QnnvQ1Hpoqpedsq0B2/Q1boxezk9firRrYMFqvwVPUvrnlUMV8x
ImGpKwc4tm0zCKv7jyWE03bcBvTj8BwkJV7rLo2czYmp1RzmONxr/mvr3ZvI
OzVIuZfgCEWnARkxkaOn6fpYav7OWmblonHJJRDMXfOE1MP1d7iLgpvRwDBp
G5/XqPqRPQZpbOjKPXxwOEL3UU2NHWhqDT649vf1dDIilbQzV9/6rUFaWKlg
J5Yuad9/SrUrH7zwcHH6ftL/EbY1jrtw/LVVgb8ucO9QkhQsK316ksvYke/3
3wWNFw1Ji2Wxwl3ov5AHl3dae9S75OSlCSwWMgmhyZgCJSZCvybmaKDd50vT
HkUPjxQWYc4ydjorPzrx03Au4QZh2r2rwzJnbtOSfD5PYWmDOtj+ALMCxIl0
rptdu3oMvXHouAVlpAhl8hLGKHeDKimBtec8ljNy0oKP0f6/6A9uWgzEca6E
SgoB2doIUnIdcsq24UEWBEa5/FALtNblXij0BZR6WnF13IaoGsXOTpBEKDPR
HSSbBeNriejLSWRQGlqWTa/H3h5sJS6ylHR0CjOYPIV8tczH4QmJDhTsEtFv
a89osAI/Uu2B/pEJKI/g+hfeyN2xul7htkALQmvpkBzKSLV7uTX9ADZsRgBX
gcuD4fr5qsSpf+e/dO9t//B/EFcGiI4sX0pEr42L4VqIPgTzjxtQirMsOiiY
CQYgfz00hCkjiSim16J3cQQIRR6vDk3tvBGrj7/Hgg+CmFnMWHsOmjqrDxbZ
gqurQzANw5WG5MNedmJbHpkA8Fh8O49JQC6tkj3634rHGNA+MSnO//Ff1sUA
N5B033eUr77jYZxBDlN3IOH1Q4VX8v2pLKKdJeZR2dy9sbrl8eLBy0tUrLtU
spFhVc+FhOWQmFTlgfjGohfBJC3AVDteOzM2NPlBuG8mZQ5e/TZqSaHBeA7/
SeaS8h4KZCQzvhWBzpDMOD3q0wO3veq3y1JrKVCYyyRSBCnl1aa+RxDQaIPf
lagrNbAFnuB6lP5aG0h5nbSbJDfaSSmnjeeazGFwx5AUw4xv8cVA8EMIGhAc
y9bH+6K5YD5hsaJQsux4TXZ8mhXOqQakMgs7ECNdTM10sPWrGQaw29kwA0QD
7HJ9B+I/fVgwuImriLINysYdpnlZcr7iD3PB/i9RpHrgNaSaumyaj9qPod6i
qZIBLgQ/PMmyVaNIDLqfgNwLPHF//BElD1L6t5nHSg/ILxpxdm1Jb+kaRmKA
BYQXyb8zUycW389TC48Z15wlPQf4u90JVGmldAL/TpRJahu3hP+0ZQnGfhA5
1Zmh7zAqRdNECoCGJlD1q/eoAY2x6vrcLXO4TjXaxRVVhBJ6l83PWJm7kHg1
BEDk9zRU+VPLifHQ7f3GnpVCNM3Giipo1+UAOGXjBYUKZRXsQagPZq1doxV+
FtiZwLHWKANqrEq8PKHqz9aEGs4nL0m2/vUNRJxJxm3v7KT0maApkmlFAnf1
AJatZZoIrxYH5JGiXDUMU80YrAQkClyIjrhE/J8csc66j2Lini5aatfS+o/3
wDgs+7VR9zGvO5yz9xHCg7GphHWNbAsBjJsPapeFWVfBasAmkH6Y34g1kI8B
XUq+0YhYhY3LAzaUJSCv2sScNfoIMEI5/rV3+bsJRY0IJWa4Qf0IrZyjqDdX
60wbuE+cMzbqnYyFf8jD810gcisSmqS8SaJntt8HJD2bnehNme7DmVI2K6Kf
z74FEMIfJobk6jcDEgw/utpgD6BnFLxMawSuux0gRqs4PbVKWNbf7XAHN+3b
jrMJ5rl97E1Tq/vHUxdjTBnFO+DYT9HoPBgSwHHg7iv5oqm5gr7dqzY1LXRM
ti+wuMJj1lzjEHZlQh/brnICU9Yxry8Y2ZtOYsnsBAkovzO2qc3RAW5QuQfN
SNaH5zUyEp6wJPmyRqpk9+wnwqPLxI6oA7Ax/PpwwOVPv9zxwXI72vDy3sLF
eiBt2dws4Uj2yu516Jq2lHw3cIcENhnzR4dwjZGj6sXvvSdocicRiGu602je
G00xsy2gRxKPjYJd0/DsAE35yck1bhbB8QaYbwhipV3JZWEw6Cezst7KlHuw
Yv8x1kooG5zU3F0ksCKWLrL55fLwhRSAN3B0chUvlaUScWSAPciX6cz9DVlH
qJU6IZYBreOcMsSC5rr/xOzzAWPnuFtr3LEGHxoAMr9D3IGikFFrf2/Hj3Ow
DSQqEDfr73PtgL9G+XGbN+hcWoQSjbyYBmZYxP6ePg5CUs0eMzDk3L8VyY2j
HBGnGFJ52X4LU1A4Bd+zWtSlAXR78nsQzV91CAvajoQe41A1Sa8m86Xc4fQO
ueNxmp3X595pS50NWW8Bynx9SuY4jlFc1JLMkSRLRugOUot+yGymEWSrKmlF
Zvu8BbNAjSRb/j+nRQ8Q5nvohVDB2kdF1gKtfNgHoaKeGE/NEg9rNa9XOTya
KDqJOoFGcWnTClMKmBGRjmk0LyztDZvtgMl5o4TR8bnr6vtrfZtEJCyjFr/T
aBG+/Lo9jCLSYqn6CoINa7Q+KHcoLzxKipURBaYz4zDKLZumuM0SUPfKp9LH
BhPRpMHWAdkjdy9FlE3DhoFy9nBysthnZxDJuqenv8lW0+eJSohbMaL6bzef
wlBb12GOgf5MF0u+Yod4HBnLsHvnoVjs2r26ES/2Ro5qhaXOpw6yIKL1Eb5a
XBrT4Di6DVyAijoK0NXNZAmD7SqLVGfPoVcczdQ2FcYLwBORCSs3IZ0Uek5u
CoBG/R7uI1KNGp0SdSPxLzqqhJyzON7UhN6ee+mHWBuj8aRQYaGCWi+LZrtG
U686lk62SS3wrfOmFgGR0bHGmkHk/a3ad3s/cgcQwNqU2OdrWzblOGTlX/bS
rWwu5XyzeRM/pKs1CnfygHmu3lluFf4DxVTcJgV4ThmxlKNyiMtugesIZoTV
gW1D7lzso+f1qmQeR+RHgsLDd8x0u5gpGyTZnLI648CURT7zHgLX/Z3o30cL
6PLDRcJgOU3T+W+8OP/GHliE8A3Ywc0Y+uv/0lB7afiFNpYwz9490/2hfOZO
46zMQuzZ4vQJ5uCDoV4e8knCUKYhNN2rf8KLHNWW00CBkrGKRA5xJvpE2Yic
13yNlGpVuzNd3lkUMu8LniV2qIaVFkkuxmTaW5vqSi1KHD2qlHNkGHqwkb7x
w51quRc7Hcae9rwnxG+smNWoO9yStLva/u8Ylw/NyZKhdkMPl6fT0NWiN9Jj
PiKBCldC99s+DXf3WphA1pn5vif87dxkTZoNiLURt8eDdGGUfmEGznZxApei
dG8vQoT1rIQaTgCVAdcVNUrG+M/XQEAPJjaP90xy3WX8KLyzDZXN0Ze62aaG
vVPi2pFSHnugYUaJ95QzX4hw8DEBp9OeB8gXe3PnVB18/MoOzYXuqoE74YOr
ThV7mPDPVQnTytx+UYuWRmuB5hhlvAnMt1Zq3KFSW2kIzJ/Ii+aBP0QAAkiB
oq36EA07fzucVmaW3p+cl0Mn9fxfgRU4UHOpBFFZqe8J7FnHNDjh071zXklI
payUTu/JWwxSdKarCFr9saClR9Jevp2YisVREObDJdGOdBKFG+yRGaxvGEa7
eNAXcp7KulGtW4UcNnwpbKCL533H0G0dJzTtMt49JI4vFSM4SY3WsBq4TQDO
m9hhlntBzQ4e4R150znK9pMhpDL/nR051Rz1sgs4UwYhKI8CQS/FYf0BDd0C
HNj2+ZgsaR55wcaj4eYzCvoUcgOm1WrPCjb30VCwUcFm5IVonQE294FDfWeX
O65sBw1abmOgdiOstpSdj59Sz7w39Bh53pMwZ4yL0vrEiGyr4GVWWm6vAghF
UI7v9sndeWEe77rr6hAixvCKrs0jmTaBLCI7whaL7oaFTnyYcTdHGOWwP3sZ
imr6av5j3NDAmaDZqctWe8HXgkwNmYwPs7+uodTvE1jr3Be6ug5JS1wcWQQD
oWCfEMfwXbd7G0D+nvtODTcfLqMB/Zf5OSgzAxyIGN9ifaQwMx5mGkwxYw/+
Q9gFAQY+KXT7gv0x1jB+knfg4bXwz52s90SqSu2UyaambYOkjVfeGxCWbQTb
TmlIvMweKNSQfDAPmFaVYOJHxfGOLiVa7S6AcJjWsHjb7zc081N8clDekC6W
gEIdVjUl/bDT+JVB8SOkXfWoXRTf9WT85Kl4rf/A6wky+plVeFhBArF3SYS2
Um4RJmI2jRZLiCQzj0RfR3FUk1QCtITJ5mYBAq4e1DSciTFqiXW31mH6TdDG
M4qD5KmMwPlOvcvafCrRSJuWtgC+Pb2KhxmedJDJhMUhEQZD3OM3CPC2//1U
3U9+l8YEmzkZhvIUfCtaiS73t6r3K7weLuBJdz3zor3Ic8Rekd0ihdaCvdPR
+Xn4TyevvWvaH8tfMNETBYhFGzvE+/Xoa1bFAXJ7QRlTleOtysf0T1qzLSzN
2nF32cl/mw2Qi4LVGITYiZO1BjEmFBKlnGEot0gKkOSaNj+KcMgOXu8mT76Z
n2758rmlK1ddDpCzejeLBPKILU9CjVtT2cvIP7d2HR3pX7CqTA1KE72yCv8I
F/8sul7zFunO4bGPNd1vsfNDt9LsKiqMbVimLTD59RcNxS7vlNNRsDMzvvcS
/x7reQZuLZ5fiufZHSYr5n0PNYu7WFlmFNOgSU1ws1tGDKep9C1UQuxoumFb
F1F3L6pxDyCBO/T2nijXXmn6G3q7bCxjXkN7OjBydvsB0LBNjwusx1n1Xmtf
s+Q+bimf3tHX2X9r1sM2T2niJwagBYHWVBvKHQ8Pm6M1G91azhyTjKd8GpxW
N4R6z+Dqhw21btJG21c18iCsK2T+xiJ9e3ppZJOAPLN81I8oShDQ3ie/l5BW
58Z21bokAHy3ZFqmWkT2ZxTFpFmiI93ui4d0eTr+mrpfjIwcZLmtByshOh59
dhmpdBzlZpeTsASgWpk3WUPhMS8Mt/ygQYzK99Bxorirj9teAnHnCWW82r1y
OufO0PYw1XK3yFipJt2Gko/rsGYnntN8lBIbgTK0Y0aKoUo+gfkmb5j1aQ0y
VqlptK7DN0Vd3e9WRNAAXdA+28yb/bTSmRNIvb6nuSY8pawftqxADqKjN14C
pdO1nezwZGEki7ek2pV1L0dlnYA6yIDyDfMvAUynGm8OPuFBmYxRO+FgXRg8
0yPNfgotaTU6Z+PF3VL51t3aje2rRNdyRBJ34CoxD/JiV0dQLfiBZ8trXTEx
n6iTjOSNHSFtJwASNF4lqk6Tf08Yby1D/Ge17zXXmFLDViVFObZ6qLBYforz
CbKk6aSAyK2f2YIQQGF30dCp+3SlmuBfrW5QfNT3wkDiA65wjaJEVHJ3DRk2
ZmKihy4tVtuFKS6KGyZnVf63GfWeEimo7QFFvPMvGdQVnAJPS5byUuQ3pQML
5oJMLqkrWe7wjM/B+eNm7c3OW3XNHQDUUbZ++a1kUqRacVgdmGEKB2rgsGHQ
hTLW8KK/IH9L4mdh37TY+qxdzR/iuvvAmDi7Xna4ZQm27VxEGahVMNlO/mPC
x+KC5uBQojfo6mjb/StKoMImIXO0DenXtKdILfpSNjwt/uH4vcJw0VoNQbGO
L/WUKN74j99rOZpi0fIqjJ60XUXuq2EBm2IhGZQkO7NqmbC704tQ1pfBIsH3
RVpx0Uce9YZ3W84ZcZjVgwF5ro49rlytXaz+rg4Ql3Rgjf0RLOWFQeuyxOPy
iZrNhFNsOrXbC6rgycg5s+ihlTz80QB9g2odjRDGpnX02WtFUkmRYwvH8ukg
YPT8/08LG4ZZAi+0TPihrmvY8Fl11yVfi9b6RYpTMCjP+0PdJUZaLVgUlbqk
d2ZODWF6j8mv838DJRRqhHP/eOSTKQ+h8OAkbsbjJa8yLGG3LwUTvKiEqwGA
jxbM1Bptyyg7bJwGrczaqxhnTZcRWH/iyYQ9bLt3UvsdrDtsSe7r1FvmbBzq
d9SWoa4cOwq9Zy95e5IRoYPZUhDyPQbxgWknz5yWHo/q026HuWgerjYHe3oh
0aIsLOuoV79ypepU2UNZVp5/FYaYDsZx5AD9/9M+J88Ea+NsttdEzMfoU3lV
GrI/2cHLbTl3ZCC/G59Fsshmq3UqWVZQKr+kpKwX6tdbz8X25CA8AC5jhHy3
NfhDZcZnAXLgEFlYDgZLjRCfeMelYibrt4CV7G/JY8v/StQHidAUiRnV3cZ2
q1mmUsxHkmuxVuC2Z7QVIHpBO8bukaGcn+XXnL3WNEDh0OgGFQkObvACC2uI
/DJ6pOGMt0exkR+Tgr3yStg8oQvjAtPRsEvAqn7FTRQ/K4iFeIyUAdQflrQR
3hQV46+LZXIgpmHct3DyxBFcGSpoktPOQkn1Ds8t0hAG+N2w+nwUIs5MNdAP
kO0T0c8VzOcQV0AecDt29+MrM1pOlBENfaw+JWwZCDwW3bjlCxTxAj5bmlJm
t9VnjEyjG5ndKB87poLRsDN7qdKcftPv22uV3g3frB8BDoPMoo5a/lkvvH4P
duTfkhqG4QaVZCHuONFFOQphD4OToDZm4Kyg3mLT6nYTxb0hnzLwBd/fhd+v
RbX1IIuMBNnC1VmEY27fNSNV4PJ/ZugUwQ5qtuw8e1zuwDPJCYdquuRBhkiH
9e71Ql9fWMkjyxkDhsl5UkiL6YC2LZM3+6piqKVv9hWn18g1FKm0MQz/7LuQ
9YNR/wFbT3imuFS4iXGmEntjUYlS5Z2i2F15lR25iUES+tGBVCY7Kk4JbVhw
kTx+VC/L+q6oKGvPu3kd6anPElMnpIbhYCHGNxDCc++A62YxYrZ6TSgNr3Gp
EXigzxGHbXb2Ujq6osWN/t/AH3Z1+YFeF6/Dzc2b5HDKVtME9T5kw4aV+Tw/
Ni03qg1mn8FAXB04ky5AKlH1hmGT1P3ahhmXWVSmeIMPUnhZaoKrVo1bAFlm
ysj2IUzg4XY3rm2tUAmAIzTm8HnxWANCGIyCo9sjHhaDvxfUA6sm0T5kNIrP
qUqqbVqKD2de47V99UHFpNpL0RcD4xU24BSwrDB7/fWyz8ejb9H323C9Hhii
kPgw9GNivG0A5HetdtQVa8I294Dj+EsFMLWWL2nixJ2qXlxF40TGTkdT39jF
/LwPwXGyLzhrudprKk66+lIzRSnZCGPB3PM/gLa8+WRQ9bMmFUctle0vcGG8
Zn+N8uON6h5UVNaUD0aHTQmCV6BUJO02B2auLvWTS93K3KscRvPXOzAZL59k
hZwk7Xj+gQs/k+FPEw03FjQCCeEd7hkwPZPLNcejYN4GO6rDnEsIy4I3Ethq
Ow375siR21S8z1gXuDj3uUD/zZ863AypthtkxZT/DAQgCyheHqYblD/MgMAX
/40SHQbddoW05DKUArlQIas9RlA58ymPEyTcNHymt7BfYef+eU8WdDiciSoy
Vj8MIJq/8hKgUKoPCIGvuMdLClagEkh3MGKIbEVH6meSaGgZg8e3jcVCpqoC
srFOhjGUSf3gF5nYdaKYos+EqFoEFeNbOsT11stxLK5tWqArENT+OfCyHJ1V
N/v2qYWTuJv77wJCHQHfEPEC8AZB8qupOFtOLNk1AXtsbMbku1bt9wgrkdBJ
+ddef4vbL+/soSSD4/T2wwkkEdqusf4+t32yVJ5m1zaVFIMFQsf1xJD+gVm3
VJSsfxkHNj6ana6h4W8ZuiaHRdWPHsDwTra0FiG4vrBabra+r2IyW5rwonjY
n0QQ3JThYApax8gYvOcYfeQH3X4e/VymICtsrqMuSqPK/Cf66GpEXoxtRRba
fQ6HTNc2xky5ZoIThX7fiUgD2fPPXQumeGFsCiXT5PQeBK6bqCI/i3Q1jBzt
TmtSl9Vql71XuY2/8Sj68wxQMNmaCoqe6RAMF0e9Cmysf4TR0UIpRTJQ5QyM
mGljrccz9Be0oj71bklK2GaofhbUELS/kbT5SZVs95v9BKz/seNT0GulLP56
0awr3tpsxH9JyvO3uJnVdXiAyfKk568+VvojXTQG1hMNx5HbeoMaeZ7Swl0u
hS/B/Yy+qAI+v5szVfXzlaCvClT2FccgBMc0c3cesgZm2J4W/npRb+EfUUIC
ALm3Mb67YTED9C/XhLAzdb8Abw/SBe3vq1HXnv1qBbt/VsAknxnkZQjpYUTO
nrVuFA+D9uMyfMlEzVTcwA/phz4GpTKMAkcdfIm2Gq2p3qiP8WrnevCt35ry
0roMja3YLXZfMXd2v3XmuDJDInj35rfJ7apjudh1roWTEfLjegT/C4UgT5ot
mYksDSZQEmajx5XnIk6XFAxEzKMFsNeUk/ulrZCfVoGZRma0Sz5uhKgPeIe2
ps1uWN5h6vioGRbPMrXhgX4Zyn3PCcgoWw5FECR4vGuWQdL0/k8m5eIhrHcD
B8+dH/ii300+vYVZLxcOFazrzb7PrGkCDBZVTJ/dNrB/aN98+FzZJLuZXcXU
d0/VuaP2E89+1CBpuixWQ0DGfHBtmK+UqE+v+YZak9LiFHsA2XBXxPNKmXAN
MJqVJG+QOssEg+tFUt3SwqELBbIE2sPVnViQupNReqYVf7Crss5CfkEPb5eW
katHtPysbyl7v7Hk+rfetRncEaJeoYhSjjF7Aa4/Z9wSfO/87p6PlEAnxC9h
dKfwNBt9l6jib4wktpa5JapbV71HmgkxFNIVtBPlw6uLnldJbrZEoB12xH2J
0FCeOgAcp65J3sOVaq53sLRbHyj4pS/39hJPU81SlUcsIhwNhrXmat9TP3aw
1zyDuY1+Exzxzd08Y5b9rLPdqY5nWog6bTE0ARzRJHvcPpxkOHmS5n9Sj9Lr
kMur6QeN8yk4CqYvzmoWByKq+IjIdz+HWc87g+4Fl0LAuzSlZEyQa5c/2PI3
rkrxMYoeIWYWXD4Q//srN9abGmOUQ4aVcFq90DCSUsFb0easKq42cvTqnK2Y
rS/sCNAQTt18J/YehwQRYj0UTMWOi6oiY3U2nqa/J0TvyJrPzNt4V4aaR7jF
uw70Q1mndOo1C4sJ6Q5vZfEveuNLLD4w3AIwy8xX3Iip/3cvzrBylMFQMl1Y
Wup3IYaKCzahxj6hPmQddXSN+lQPwvftU6sY0+RwwgGBdl6fcSGKqaOKpVOa
eoMdp0XySWpFhvagyochJOhOraherLTO3XHm+3m0Izq5PSigMIo0dt6T3bWk
ca2sBQ9ezwYzjNFW3zvfVSkYI8oGHRwH08zhDsV7/hYEoJ4vEJUjwnyJzJlA
WE6A6Fl/jF3S5rgddGWaStJNtQhS0RosfPgBkplyp5D215n0UyBHsIp5DFdv
hOtuyGXRu5kUlEwbDJbuKMVoeJQqp/+MjILpUsvy9L56uHkNSpAZ0Vm5iNzw
TYNsvC61jdFTZLTg7HSOjntwWb3z1ta/Zmbo+DFFKr7jRSTUKaQAzK0UaSCS
N15AezYVPlyd2zHm0bry6AMR34h2oGF1nL34XjC6qycC1jktBV3qGuEb8z85
gN6CLEoUjXVX0N59pKnQ/+aG8Y6lm9JE5m2+cBrpg1SNaIMR91TrTyNTlzIn
/pYqiYmWSv2wmdPfKyeDZLLnfV7mL0mJ4+Cs2kaO1btL1gJO7Nwc/QRdsIUt
uLMoWd5YD4u807lC4yGX9H7vAbUsUaVvUGUXdRdl6YXz9tv4oGaJAphzIYOQ
cZ6URbqzD82NDMhv6IZHhvTBofe7GhS/nUJz70s7rhb1zEn6MHLThyYZVnnj
6LQ7mQQt08atSYMU6UdZGEbtcWVhuQo47WHqcdsSd6uh/XZBd8/rneA8z3TO
GjRAiSvjmQ1nc2mtkxtgb81GhfdpfiyIilF37ifibKf4RIsRlm0/GFJcPo6Q
IsPbDMtEhet30Z0XKEZPbdTjguQt30pt4dBMzoGhXqVCePk0fXkdtWHbUdFl
Zrr3EGOCm3TJVDAC0FIQEQi+tv5H+sMuRSQn+FTeSbvAkZhyZsHz5IKIn2TJ
+lVGjfQel61N7aYTO9KInslEGajalb6ncTM5H1NZFyHw+4AsIj8ocjb3mKmO
jra7hPsy+/n1s8/uA3dapVz9eXAVgFtFly1BCR5i9tOta7n43FLaOWVZQFm4
8ELVVWFQ4To/kaFasIEEeZ7UuPelp6gL9X9UPJhhL9EyqhYANNh3h2btCctG
+rb3mN2tUfRyfrMf67nkRFeScMnP2DKb1//5jmrlgLI+NyZa3WbqkEVxcsQZ
1Nv3m2VqYE4vesx8wtZ9cx4u8GHw7M/AxXNrf1Md8x3Tt65BaSycOQfUqzjf
hwKPEDdY7aO1FhGsq4eT06xNbMPLHUemm09Wi33CoO32JGZC04y76k9Olrq1
ZwsiZwNbz9lkHtmYOBqPw5i4t9WSlUcFnGtqQJxEozmDnibGkeuiVjXLygbW
8Q1Sw76ZGO2gsxhbcBtYBmWpketA2zTSw4eK0lXNrPSJtIThhsvQxXVBQVw8
RJqEp83zIdT4hpJhaJ1yHGBUw4WvXCAf4VfLBYM4pkg/wbsICggDIH6K3Hhi
whNEal2e3aNhe6elfrTMfGXQGc+uIemGSeY0YF5gLmmZekq9DAwrAZsXqIJT
vn2yFnYpcfGmzrhEueB8lPGFPGWC0wDg4yCGjJ4GHM2azz13xe4e/moBz5VJ
7t0aAkSTCyEOOvaYxpXcleRWjvilKcqBoEFCdWluCUNS/6fzoD9vF1lMAkCo
OcvVVrRCBbSdwlCw2boPkLbNSPLadWbRkn30r0u9D1mxaPLGKb/699YUkDZD
dPuM2BdyWgZt7mAXjb9FJEJ3ps49T3xNmmlBZNS4sinm+sh+Kb2/HiKTIDx0
g1kFhUI/Iw5EpP9sO+sPqCUjvNt+9LwpN+7drEUZvJP90xV6v3B0P6iB/0aN
pXCbjpT150EPCitdej33E0QgDOguzx9yYaBO+1XvfTmzFodOdG1ywFgyF35e
2+JybTSBbtp1CdzWVO2HPmoeQj0Uu6IJbPopQLEMDThSNnuoXRmVJhgxjGaT
TDybG6DwntXW+YbR4+GZvKIq6dP6PvdPcRk8zoSOB4jQLy3+8BCst9ADVEd5
1YJEwv7PvavxDd44cHwHupJ8jcShCWvfMr+GCmC9guWFL7K6GCHnBYwe/E4r
AjTxuyKnVvJqphOj9p14UeelMWN/4Ef2Aw3dor3y7tt6L7nl+2pVMGw/T6ly
dRtnXsyykoHH5GtY9tiokJM3PDx51yhy5dJU/DQctcZGG2pAJlYYyALzjuxZ
Rvt6zk/ha1IdkR//7Qf6HNzOUkTIMqlobV0HTCdvQ05YuT++7TIOqLFxRYrW
bsd9U9Q3exDvjlypuFo65wdf1VcFV02X8k6YbYVcLC3afiQKa4wKGMgZxe0P
KGAdfTbVFwmQGh3ZL0FeNyDZj8v1Z2oy1nB+gHBIGc/CIDAWTY6O8zuq0fer
nAiX5QXnQfMox368qczGd9JOTfSOCpIlsSc4NrsNf0DaMx6lwpURfeIopp/t
bg3X83/U54JDRfztp0iCDs7EisIsZm2I9pSVh+TyfL7T1mFuGDggJB0NdUn/
UYpHgR0wHQPG52cWi5FmU5L9g7r89Xs+6TJt+rruoLSiH7u3J4GEKVjqaAW6
eWlZbJklbGZyfmunyWd4gaSyW3RmOaJofTf+bdRTCaPLLu6qDFYRkQk/rj+n
NylAIEtGw88wgSzDNTMvG/NPXbSEZNwkvWUHIkiLpr1qNoKefr21Hv2Vrh1q
6GhbLNt/yzmYMW75CvQ+Ah6vZ6JwBWpkeQZaULBLwzFnncRr/TUf1CleNP39
BYsA8CJUyAsJljpsBOvnr4VOG1sy2NjuNVPGQlXOk4q+Wsh24O88FlkVGIt7
Ba3RvNzQe8/ZBvlLWzgS8PAFIP4NPUErJvf9W0bilODgq6PmHrjo1XLdiXdp
ypGVyK1dAKMX31cDiRCgTxHCuXCit8QRWxxqJGNTwX5RPqLH26nQjjPRc2DF
sF2Qedu8gCIWLyRLLabahfKxlRKbHcvdccbYA+tIezFLqUqty8N3jwKNPlL3
ogArw53yI+EEtpeVkHOoRYw6iQo0VxNLX6HKBpgWCibfkbKYzcudcW3PsMY+
HS1QlhxGcswpT/xQHs70CWwCLPqvUI86auwsUM3OpnVn6D6x4I7ayx94uH/6
IzOdsf4HA8/qKlLzwiQe44RfCWaVFsv/O4ixyAgnWUQj8QxY6NRDlhYzOs20
AuPkkD/VqvA84qNy2bvPSe+t3JhdIq6p3hD5MFuD8Vmizl7YT0SnSA1r2R7l
7THAYmYJTDaYcrsqNMzBBOWuuT55GnZOvOkvmnV1hEhEkMW5xInt3XBBmtLu
errNE3K0Kr7EsbEPxHw68eqv8hkJGn3yS6er018xQiL7rLFqy/SGvODVPZJk
csyP//jaocaXh4gRp04DOMbznXdhi2uOCx7oxG5fBvTXhMpAz+VrlexG8+eM
dXGmYmAODgSolmcQ/b3d8e7UVdVTwAOY65/CUGumh9mYTEVqLwPCHfzeJOzT
e1Yc4XFCYSF0wN81GI4O1Sk9AMEhUtXieZcODfgk1/gAnOlWyo3LthRoaJDX
G8kT5NheImjwhcQiwN2gBcwOIj96rW3qRTtYMuW0P1YpSd2PvIbuE8mXu2xC
sgo04YXyNeXJIcGM1xkVnQ8Kt9njI0/ucMWPRye6ZUMGmhu7wKtiCTmnC7ig
K766prtsADBBmZ82ccQGnDrpW8lJd6X49IbF0oTitpNgHO+gVNYRyKwkDw13
MhLKrnWO9iaxGmkLXifvGAt5pUR7hxPsv0nL6QpfqEauiwHo2Ji2hmfOCt2f
LLMMlB7ei7Ww61r9TEumsXcPTcbPF71lwrp0WimzbY91Fd1aOwFKGiqDcmUX
6fqTsYIKP722U4ZkmN5FQeuvu/ZeUb7S0IxCj0BPYQCmRj3tyUFoA0ta74qP
ec3TRYtqw+3JdiFqzZfoQgmznHpkG4a+L5gOM6a9Zj3cpEgTei4J28S0nxWa
A5smqPxOl0irqfvisG+b+CPy7D8SJAJjLLjwzpJZihViP+HsRRSTU1w5JSVX
XkChrJyOGswRBvmywOti/tkm4IhocQGti1wUKmuixP7vMjosvB/LV1v+ZkNB
hn2CzLK8vEdAEfatFbQeRhTsvOW+uQSJnyRJAuiOCI9DLQKX4vNf+Gn4W/Qv
uI/SaAysaQj+4s9XLxrSF2RQrTUoZ0y93bSJw17KSGAHwv4gKLbSDlPzxCaT
1ZLYCsZhg9erSxBMA1vFgOLke5D1a0WwxUqpdnaswVNge7o7m5JfCGLOyYH5
bgk9JZ98YZJJOT/MoQBtJ5vWMli8SX8+byk9mXNTLUNjdN85HF+HQdBQt6np
NAVc7XZquTuVYp2YeWY8cUNT0QJ7ow7B/orgQ2ipUPde406d2YOWrhn8cJkk
vsZsc8zuPpZ5Q7biuU4szY1ygGKlTRzpaPyIp6j5eRyYeeRqOKpWy/qYE1p6
XNOsIP6xhpMsfz8HYhp6IMBRGNfYi+e4FXWdtcPPeNHa3DFLCpfTOA/o/XRG
7P2e7FgVIWQDDufzGEDb0fmpaF+dD98rFfzbAKCPAGXe4PyuQ6YG0aKe6KFR
X98SG1HLs0Z3bLuRNwGkS62oddjpEvTZiLX9DPQL4qmVmJtQF7kvMPouejAw
8PzdYoHupICL7GeBJ06gohCbK6Hlwleq6ugKi2AGwdW9g5HfIhugb+WQsCLY
W4g3km65cXC1D2caxgoUAN0QWSrP+m1D5cJWGlInhQnglbwF9z5mlLj1dMRJ
iWBME/1jXCS/M1PnC/Ie0VP2bIwmOon6TnRJM6G62l8OkieWqa/NiDDX8lYa
TLLjveK96r9KI0dpdGqzxgoIlT9OTb/SqGAZeOQe7QWmcvFJ331FnoWGds0t
cDzBrPTLUHJr9mY4/48zrvTfoO2hUxtmgDePVFiviVRDKoDFDRYXM2u82UMd
vYfxJ0cEvawxrDthHRxoyOHfHhpHl5D0ei7iNCu69i1CzIGyHgfFshr8pfb4
w6gYD/VK6czyGCM7ES0zblcIDm6NVFha2P7ESI+ec/48NOGzNpmEPPPDLxAO
TVt8N6LLA531aMwLESUbvTQP//TisJ5ji80z+jniEeuvFYx9Bljx1ECuYcqz
9R+tDsEd+59NLQk4V58SI50DSn0OTAnbwnzF1XnUXaUknJ2E8DHp0LoBjkt3
OVTufZwh3H5HHzZDIwd4+hbTzFVDyDRZYIaI79LVHtXPdJWZTTSSMm2eVpj4
NZYvkbseOLJZxtKNFnd9+WiDN3HvvKRjwxs5MdO7etBiacYHdLJRK3HjoeUd
DQyaRJzT0LwML8p6iLW38CtHgRB646pIvJEEO60UcEb3/4cix5DhvwoXelUP
qhcIexC5G32IFQdoeNfdphdpWlullXlSZDGw/UsfqzYdqQFULelqsSXx1wiE
a8Bwui2CPykuewkHnJuXY+km6oGdOiSoAm5tI8YixRwiKuGCVKkG8feU68g4
DQkX5L6/Wy/hUCx7deUk42CSSBWUUd7aUz7W5HovBqeMlm7P8HbSk9QfY6xB
bSe8MuJf2Jbq9KpmPaHbIFPd0D2fHAv+V0ITQ5HxvNAzd+OSz1uEfdpjBN6I
MI1LGp9HM4aGqP05O0vo6M3MKN8ZmytfsRVcIILpw5zDui7I5jFlpoGWIegg
WZtftBzZ6rrPxa8pirOfas0Ih3xGhyRax2TSvPs9gUGi278rHw6d4h99oinP
CFsiOu0+FaziNdw3z0+8ax1+tx1xLcafyxID76tkj2fx5DObkt5FvJPOQnKW
nMwCG8/eJxGznUX5uCi9i4ZUqVKCoKilmtxNkqo6hH6dP9YplY1OtFlXSTK9
Jmi6i1e6HIXVSsn9DPP8sJfkcFaQbXF7vwH+G9ftsS2T20XYuSH4skeMxCA+
gtyJogSQcs/dc27yOJuBYfyh+scHMrb4hn5aClYELb475iQF9jVC5dScrpOL
EVm0c0aTMisyNkI02HQtPAg3YIlOtq4uoDHbkqy3O03Cgv2EaoAiqcjoYs2X
6kGoXzwtmeeKesJr/qe17Gsa2Q4678LNRa5DGG/GRxqya/4WsxhsyAf6mw/W
tSIi+8O3B8lqglSCaKi2Dlo1Ra9WZdNGtjZJOIPpzSkpBFndntONQgY4Kyd4
NGXKB4lnARny9wIymlhzoGyN+jvgqpL6UO4G4oSJHlt2tQFaRzbo/8WgrjnF
sP22nYesnyOA98hx6EUxlzW1f8YRgyn4OSbp5gO8mConU4QaQJnYXvZKHjwF
pP862HvzYJANLqmEL59kXhCTaqn0+c/cHn1aPh1zicGGfugJBe98dtvNytIX
5wr844mRqhHWABcTtPbdp5w311pwSkWeNFXKw8VqoHu4wwf4Em3NPSFpVA3L
0CLp5jkgJjk297f6u/vrJPuN3ZZMcJofsIJbBD+GrWA2DWspasB6gCufmJtz
RzzbOFiysR1fu/MdnxPBSPgJdpb5SiLjVamFkQRRKHl25X7gEU3Jt1VmCGAC
tU1GGtkpLqGZdrbP6Iab4gV/ekZ94w2IpQOWxTtLZ3j9HA7E21Q52qPkWGAg
KXFnBTKMDw8DqbvuF1usIWcBTfGCAvWBlFwP0/lUM4MBkAVhVvVZaoyCiRty
gj072Y71EI0RQTM6HOoJfJqU7wTmcit+IOEMSR4Fv1o+iyPtQctCrh3Y3wfe
2Ow0BeZfdGL2UiiiomLz6o2zOhRx6+WHPcyOdgZCzY4ogzc0f4Nwh5g4vS0Q
N2qr89m+Hvl6mEOnbidkaewaOWf3Ny+XaNDMuD/2JXIScnxTB+zWzwkERQ+M
4f8+W4pK7NZ5ote2NT7JNtHD/+vWhlJgRAZztZ3QIwfrn68Ftpu5H1Fx1vXG
ZpldBMaFu9Z23CO/BJFBBDYqHm4DXdoCkE1+LA7+c9kA6Tw0jk231JmpzBW5
MfHaTauLjRlIwBcRrQKsMgrHzhEFPStbaGPfhryZmB35SmbkIS5R9usLPIN8
gTQesy7vMk8ZqIu6rQcqOy3R+/Ig09IOuOKYoxEu0+MSIjKokkQWNOO2broY
JCbsV6r8sutRuBGKN7Gx3A5HJ4vLAooDxPKg8LcEo38XHg3ghGIXY3V8t5FD
0BPh1wOOgut9xo0+wmr0/HAYOqwYXHVOprDHjRqNG4bv3rNXUkIkwj2e4mx5
OOfPcFrPNNrJq0ONX28KrKjKmQlbnT74shSWzBBf+3wavk1U/Siv4J4NtsiY
zsJPqxdHs8eahN1RuzYkd546MtPerogblBBh5URUpBPpoZpbIFXvviU0KMfZ
Ok0yfy6eFENi1AX9IBwAW6pbh4IJj9uGwMjizSS9Nakh1H333lToPImdvm4T
Rf/6AeN2aSANtkEU88V/fbjRTXSuU1ejQSIe2fGk1QJxdBvmL2folB8erPd8
BKuxz3T8pwt6MCYKzz2rGfNfWzeZm8I7Ue82AzWNLkgSnf3IYQbc9mcisYne
sKy/YBrme9TB0ZPHYmBR6PbOb/6K5LCaBaiU5PCF2KNf9A99MQW1UQXPpnr6
TJLZU7ANRUI5Naqg1aSgYdh+oAlXhaiHF+W36AubdXfr7HC3cg9xM1KoLpIp
uBiwoqxAY4hHNHUDXGJdP+A9poZc8MMs4Br5nSpQ/7/B6XZ8Z5nfroVg7pc4
eKCx1KpjpXoes9pXlQtBQFEml1YBR0yfTQpyzNAuXijxoqevlvU4HBb1VF/6
0p1deOs9mUQMltJkWMfKeBPlz/XigB7BIKD9fK6+d/caegtIU1BRLje890OO
pkDPg8o0xqBKPeRZC+7myBJBC0jMJudSL8ZWNmoq9vlKFT2WVV/rdkMusIAe
kzKAjca/KF3Elc5mJbgJzQI8sfpJDVtW1dpgJr5pl1+A1m7Pj9DoD+KGjglK
w0Onw76OClHTmIaNxgPOLTQRQ/lElOxKXpkpJsAKoINIpHXEeqroVTE/Zp9X
j6s93ruKkAXp31UPSKfjB4zS1xPVybVyLoxz6mcMsA5hqvfODwTb87tY6Jzu
MSmmrJwbapypFyP4kHekSihsW5BghU24jkxt4EsgTFffuopAE0ssDs/BEsv6
jlgcFGN9miDnE7OF93UBclZahn6goOiUmwqrZBE/r6pepm7sJ+HEptZkeOTd
md7CGyoOTszkTKchc1hRdA9jdq96+pd4SB4Ucaz480dNrwWSzvvRWLi5UnDq
1XeBcChJ+Wlfkg2FcbOexXxzSMohdxVHhQlyril7Dgc1kp1wcBWJwRLY6c+R
jym4seyHt516YA3x1AmBSqBgNEBRTEWSsvO3Ih1HtXNqEWMg6WnCrR5tpiyy
hd3LjJR2fGcW3YEiopiz2flJibZmVD3Kf9UiU1JD7F+nu/YqjVk4hc0ZZyv2
sJoe/Kz46pBwmJH91zElc5jfywLzGwjFStI5tryGFikTU7RpumAkUx39UjeF
FB87sqtyAa7VHBQCjn3VPnJrbUzSs9GJrCuUUX2//n6SUklKv7OEPF2WmBeM
+WARODHzGiEavWyuD22Ul9uJWdUGajc34KEWGS1FAPQAHYTt62mJo9pzANc0
Qq9214MvdcXdgdwgwfjsWPRggOTQmcB59fyYh1Ad5ZfcdKL2fdHnewtE0YGc
gaRFrl4jCN7oQ1q6Z3q9Xolc6+fmGynRXBqsw6TrEsM1vGpY0qcI5+lAn0it
VaMGbZraetmM/Y14IcMMQaFCHSWWVPWr+Hb3cNuT9BM/hJcisgrpOTJKvARO
8SXUacTYEbdSYnDgS0VaRUfBoJDI9aKdNgTmQNwNQmCEVGZb5ohAngfqxZGm
lFhmze13RUzginaQSjpRSyeDqfFhOGZnmuBE0q2ZFHI3jN1YXi2hbilTX/TB
RRA13HrDbrnfPY57bn/16hSdP9tp4EANgNni37+qvPUx0Yn19HfExdxOAGw8
oBfAlXpsfyS7jbfqIuNNOj5i2WRI2np/9/07gUHjYiHcpdgNNkFC4DaZPUTe
VBXLqHmRciRCO1Rm6HSuVYNxz7mzjP2SezFwFU+MoaLTgZoB3DaO/M+GRL3b
bn4heV6nTqIOmg4dYInV1N5mB3VGWlJSmJ4COCgOym8+cwv5pitZobqHAKhe
7lT+eFZs9S8jKUAQIV3QXET1OZsb3wWOxGbPiVLnhiVVXSBPjivFIK1s8LIK
kdFkyZtqm50kbEQKzMZKH1l91iDZHBvRKYNwxvHI8zlYOesI50hntrK5pmUn
ynyHn0cih2MrSB4F2sw66apd46KDPEKcU+sQdIC9Z+qTeavUaWbvkz5Qbj5x
T7T3W5NwEcwAC+d0YH3ICAc1lNStFJ4ci/0BhkqzMpTvODevwwTrF87RIR3w
JkXEdWV6JkOStd24ZFBznzoWDoTiz1QrTm1Nn4dXJ5HN64iI9zdfrEKO7l/3
vuxE4FAvET7ejT+kqwMjw9fZaOZH8RG8VTsP8pA7sOVCK+R5A0ijjuToq6p0
R2xeCGz9+iKqASFh2VaL66yS/v3L5klVaUin2KL7TdzHi7YM+9mmkhpgjFge
UDcVprM1Ev+Td/W4cNJcCN8Mkrhjc3m8GLdh77z1aqlRohmaQh6Aa6U14ail
4mmEfH/g444x2OYDuorPVPlL3cJWXetVSDJKy7SqVpdKTyu1y0ErfjwZHeSf
Z+w5Wrqy57HoEq/u3xT7qV9ElCBmd9jf2y8liYgoRc6KEbBZiVf+feZy5jtJ
nHiE+tpitW73IzzyceLIzBIFzddI2nd6alN+Fzmy885lz03gbn0yGVoJQ7NN
GS2WDNEhgdlad/jrmGvi/s/Ksz9kZjMgvDmcgwKteqVJrZDZx87MUVaMHJrF
fuudyjRDyhaj32rzNjaz2NW8/5w9fxkMpqj5PTRdER9Op1MFDG9JbSykmeZb
PVfDLTkFFUe4vxdqR76zd92jHmOe6lNIlZplAFEjfVNkxgQOwbyGkBNXi3d0
HtYE7DHluCL9UVPZuU9ap7HdanfE3a4uV7RGP+6iw6xghmjzuR2b5vbYQ0/m
pIloUqG2JwN9x3yXZMWu1uHh+wpEhhHQ31XJV9u8SWk2xih76BgZBW4aJ1H6
xmMNQSVxGMsjjKU8RNZIYeDNQfCM98e5cqa6d88dNyJUTb1yC0W3XHAVZesF
EC7D1DLZVsQQ40dKXFO4SV8yVA0Mqx+qB3167z80h+b7rbiHqZZW3daxercB
B3zAI1ELPoj5szYAXbw4WwgvKbaX3GjpBjx8XGqJWlp/3VFo6gMY9K+f8hrM
NEqBBgX4cQ+Y527B+sDjNkqR3f8PsYukVNUdZpX/WI2OSO+09VyfagpBOvDj
+vUuJOUOUT1bIp0mATbVP3Y+ifjBwsymIO/RM5suRUFMzGmPDa/jhzGNEg1M
YbgSuR+x9j0ENxcY7c/QQ3RJ75kSEOxZd7etd1o0JmEqRu+UxPDlmwTkH9nv
e4u44OOfeShz2M7WsBhibS8BexeEi9B0i0Grnp35alufx957JO6Wx72vC5sU
fHX/zJ4sz8ssokb+akZ+46A/iNYUyFT2ctedN+MdI/0Ux5xkplwK7lzPOkKo
dpi+QNLfsyJ/Zc5Ud9DD53in4NlNBOlVpqSwwe+DfyYWeZUuF+gCAKy9QlWQ
y05ZW2PzKh+sTNWczHA9pqTIcFCKtjCQ9vrBwn1qvDtBfqNYa5/3plifvm6D
S5nSQDwLkN4tWX5AgPtlioLEyi5gne18dm3u/n7ocbjO86iwfD90xpLCezXv
ch0rdy+z51IkA5Dlzz6rsTcRm5fztCYhdCQz2Fy2gd4fhTNrAboLDVPHCB+J
nyz6GibaLj+VRIdeV5IHS7HzmQzZKZBq12jUnKYhVN81ePrIvgudXNz1YhiF
DzkqRDWI+yMQq1jc9tQRjG6HKIraAdTinKAInHKqNStLID7/iUMQHLF+S1g7
z7oekiBOetYnbrAiaOYWzeNj5CCVhso+ia5R3ikITEU8js0gXzT2xCJN0tCn
j+STqqCqd6yh9CEA5CCN53//XbvvnIsEO5HGU5ehhz4wh2q2z0eZ9oEakzA1
wNiLQcF/ktc0IAUBC3rPQhtoQK1wkOrEjKfsIuE96yKqrtwxmJIR9F43ti0M
UK6j4kF3S8Q0iLkG0BZwWH7Vba0Jtm7ApvXjyhipU9ZCpaAXJy/KoYphUAiv
KBK/Lo68Y+cmqTZgFF48DDq7jmYcttatQdF0nwuHDr+0pfVtjiXyMh+0/SlL
rtgjcha9yjPnLaz+hQ76RHuL2PjmN94+wgOmWs+vpLkhwIEkc1sPSXvHIRtW
C0V/fc/RiG1CaUn4aIxGhAZe9ic77FgzXzd4w8yWVu9zbFd0Oc4DABfxw7ok
tnGrksacxzQZLYyhmT/glsGp+PVpudqWpRqz+8ky3YramkRxQfVIJ0UnelBB
5FaOqiQAzqURUUOl7dUmEAIZIKeHEg7+T9/P3itAS2yioWVEZjnos9tCZD1A
jinsgnBirsEbSv70PaugfbAGgfof6zrmMlIGcpwJX7lXrMVSh0oxdLOjolcW
bRO3x80wK4dxNqS4BAJE5RZ45Y4+Y26+EEoZPYoGpTX/EM5/5tX12c+UsH6z
Q+NAQP+qoZIsBU3Pt1T3om0748yMWp4ZIRT6+cIHZbDvxMpDabq1WRY2TRXU
mziPfjlxNi8jLvH2OaT8tS+gMim0GhgMUiIamNEbOyuviKUqd9XSEhK9xilA
WI7TiFQHO8hbMMG3x6biI8yZaKW3Gn6UCGL1ssfbsNW+Su2tFYdrt4G25TJH
qEtr5lmbbay/HldgaPPYzRxgq9RgNMDjgI8U4ct3BcX2T7wm8C2i0V42EgX8
g9w+6/Qbb8RntPhgXUE5SdMNMiBhFUZCAa0yr9ioXfTcQ/lE3Shb6+iU1tAN
d4ShXvs9wAKMT5p4uaxVNT/hGGjrSBqevD5PNFBU3gBd5S3Du9I+erqVYIOj
QDO3J0KKXeYU/y2l3GRDIWCdEE5a7FwpR3yv5ysnwb/EA/Ckj/YV41zjavBd
BdFdDyo2apHYRHoLl+t01aKMxqhNpEz00DwBUtXDomtW3ufVBGtyaJ6oX4ZU
pWrNmhsQccWIQwNGJVG3LIC20StQYpAgBPJLWqQWY7V5owoLDiHTekLZDB3d
y06NW3STZ9cHp/LUQw4flEK9HsbUlb1Bs0X1LHnAQXArnb0wQQKQi7oJTsqC
NjgoGZ/hxW3/WDqVwcysHmqwrPBSsH17v4UOfPaJQHRyQIqr4B5En4Xbwb11
+2dOt7Y0z7Hg75UATS+c/Wkitas/U850eymmYx+M06CngOpzxm7QruMum/LL
eGGMMPfqs2En53iPbUwtbuoNqEQ6aLHeqt99iwOWmfyMzPTEgc90fgqXDsgm
uc+ub59dsDgFkNhlOYYbHfXBXvth9Mq5xbY5alqnL42kM82gbZI+Vf/PTdym
xZLbURaqOx0dhIJsEl/nYeWBHsC/B0gMz7lzyTaEndVSDqx9iFchJnUTVgRM
v4Gn8vdTmI9iyoYuWCMMWCKjCRV3m99sAyxadS7Qw3v1rtJa5yeZtMa8fHKH
t2Y2135tSmVnsMKwMlkK0Le2V5DRy+AElr2fh1EL+2KAcQy7imGKaMGso1xH
ySrVrYV3lPBr02dyykqFCGQvmty2Z0vmOQJ0AuJ3QeCdovfNxafAHCYluAJI
eoYvq1B4Mbngy2gjCnov7sZjAI9VF7o3xREAUeQuZz6EmPOD0DxtNc3CxS33
wADYs1qG5lTjoqfsX4a03pKSkY/0eDM87dpQNbAPNHm07xlIAUO1EX4KD0Eh
NNEqqGaPcJBkD/xKSqpspxJHlhm75BGTjxCFoQtMjbeuB0rlYOI0+G3KboK4
XjdjgPUEqhRvKdUwKw68b9iF6s6iH9KJgZLWbpkCpmJlKnN2QfPVe417PQ75
GXjIp58e9ZDIGVN+o/a+xXVaZ3QUb5QdBcQdwZApSc2xqzGArqDZSiTLz1aI
tptFF/Giq4s/V/ZkSF7UvIjLoRzrDR3vcdfMJgGeaj9YT7kKurMUXrhEiQH2
TFbTA72FzM5C+Ydt64YXICZCNoks01P5I+Ua021YirqqLyISh+jHmdQESy1Y
PSeCOPVrQ0juASgceU33cq4ZovIE3tv3nn11YUcnYVtckVRu3s2Ufw59FYYg
tJ6c8i0s3CyBq5xf2UOxdvG3Sjgz3LAyXqgGYvdYVMtTTnUghClqRdpkpoui
Nj0isQOpn+Nrao5OotPRqHyfnx7EwLc+jYHfSXCz/+Es1TGfhgS4WpwcAswv
AapobeA7cnBNQTAnDFmcZ97i3UA/rp1ngkP9pjl3Ru9X2J+BAMdh5YW3TOcK
tQFH1FEp+CKZBqfAg2I64Qp65DBaD34MzE3qGrb8vJQkxl4gcilTdirvksmQ
Wo/KWmSJ5Wy+cKG6OoJI7Qvwaz7P0b9JmDh+uxKTgLXlAByFvGGwv/l2fLHp
cuLgUyw9bXjEzuTl7wd3tqOFvzzzjLEyu1ZUmfzqxlxEFeiJ7DfgtbsqO32Q
sKQtwzqwMKR23tXpq0LyWqfQvqpBl/sf4a5iE4ucMpNPR6bfM/TGPNeFEztY
QiQZ9IRNZOjpsSC1e5NAHhwH8yDjDQlYn4kJm/xpxRaJgp1U9VnSIT+qYrxl
A1PPV2OOlzxddhg6Y38JasxNosYJdWbdo3zmDkHG2xKPNfm9wmL7aHtd+WGZ
n2aXqVbHAgq+vmLCE4Dt/j46p0Z3jg4iAomPnIkJIVmBJ/ZLcWV4Y2qWpa0T
L6CYaDdmxXQpLKwj2J418nbALlXly2jKQwjRCtnOhAEfvQTaLVq6oOtvGa1S
qo45rFc2tp3VspSAMrY9nurvuoIAn19l978qs3EnhIDIDmDKtLbQU6kMuKwj
m18FBI/vo7M0XC5Tg5qF5py0nheYiIKtcxZOxTnP7muKgDPzHv1xS0D1KT+K
LriPfEvZQUFocNvT1O7xXkEGBYD37LYnhRzI23OAw3mYtO/m81NNcTOFssbp
ugyKbaYEMs0MC+5hUNyKvpN0jEfCzmM3wXrdDAuzN9vi33Cg5mdT7w+iVf8f
96YV/D0Qy2KQShihNx2Iya6c827kWuxBiDZG2Pb3PkaTBNTFz+2WIG69rvnD
763C8cYraocNLGObDxh3pRr5EDQIaq24KIzPjgSe1D5vTELlc8eiXpkUJF+Y
B+QP23P867ntESZZRJADmwDNbb9m+S3iOZdycYOh6dy2AHcmK3gvD4AK5qpG
HPHH+nWqjxFab/PQ+FttThAB+xvYllBV+MB3J6iO4ReoRweQ7/hZI2Gm8kmH
V6Of3G8CZto5vBrnyCDtzoigURj5+hKsN30jy4CVyEj2iAAFPCEqABGOmw7+
uURCwIB0cO8a4jMlHebg+VIYmdJE9p5uLxH+9pPFhmXNf936ggK2V/NalQYF
WPUDLD7M638z3xnKGijrvB2eGYK3BA0Q+M7Fd6aVeF8szsc9VWNIKy737YKS
mwjl45MML6lR9iMIKUpErofYTXSdbDPMSgT9tjQ3XtUmCT+FRVJXmfufUTsc
Y4gKSUn1T4SgBrFy6f0hMzIAut67//fICdd3AG0d6pi8NHURKeciPtpm3+xK
y6EKIelqZvvKI0aQSJCqvQQ+rxFaSuWUjL4Ql/PmQNdGk4e3UrJMIUmcb8ub
ZAGjWq6YTgOxcZVTyQrrL5mhI6pJX+TxwJmU1aosTlSFRIrz2A1XyavvksQm
Nn8UkevH0Zor0Zm5/0m8PjElxr49ub37vrWxUIZalkwmf5AQzxtatoBt2Z5n
jN+FAkkfV25+leb/hS+fYgK0UiOz7Apb7hwpieFy9iZaSdRBHXGw4NRcStjj
Bezg1iughPC7mj7EWJkWP5BOuZZrZ4GaCbt/2Opj99j/Xi8/9HZZ9BllTEYO
pgYxo6mkWVHnInBhFsZVWbg5OKKBfurMH4cuk8Qh0g+T0Zk35bX7MYEQT12M
5jAT1ndiIGvBaDlq0AS+YILoqUUmxPOBKcrwi7cFBVq4O1vC4V7HmzcOKJON
ALSzrpvtGyKqSuZXYgEYqn7jZAOhxnCWTXM3TttV8AYsF7+nH/ItBPeOon/x
+yqmSR4HGrue8Dy0Eya/Rh4VgXRBbWZ2SS8Eclpy8Q4hN0dXGBuhxfDuvSdc
axpL+4XobIyviOH+IXaobTmvumQ3ARhNSZYJi0eB9fCpvKS6W0F2kPurTS1E
D0YkfNv42qIzYrFkSrtDKZs23sDj9pNJ4PFDEDSykfrcpq4JnIGc0LgVOa4K
BUIzCjbgN3HpF3weBXbifqtUhz9XM8ZkuJcApcuFIB718IkuF8z7K7jGFY60
Ph7Yy7TmOeqodFaOyM61OvI7iAboyoUIKgCcS9UTHmoUnJ/uGMZKh3mxv6jJ
Lvs1dlOlXuyC2I5WG5qGie3SfmhqIU1Q8wd/NuxGBmO5pffTvESfo2CFgp/1
5ZfK8iCSBTriuXa3JJ2gsjSXKO75Ogf/hNekUuiLa4DdemtuoDghVqvmNbv/
IH6Q8OAvOIaBpBcHDgQAmZ8x2mNNPdCKc40PHX9xuhyXQC+sCbbDvrOqVDEm
AD0IAhtTSP3RJM7B2mELYhICfw5HqY+wLqWjZzmN3A2Z7ThnRr3+/+ewVZxE
0djw9gfE50h/dcpSOwvXgHMD+4R3I3wuExVXldE41DP7uKE0D0gEBKT2GqxZ
YQU/D+ebtKPD/KAG2fGCvjlEUib0c9E6Zd6IWVVhWZKRisz8vSHDgnEhHz7G
YqdpEoZrHRsoPUAK9Slc6JV25jTgK0oSM4gDq+8EjJB+C89wEUvmTVt1yIbB
ZHxedomVU0SR/0r428J+YVe+znNq71XKF4MV+t0/NYNoHXwbYHIBq47Tj8mb
vM9e4K+uLHQSQnHspLvcwRjS2heUDBLZnRKtX34m/YYRVrktMpArD5Xqr2jT
aI8F9qsLrLINbMy0QE2foGeWz9S/7wCzpkZC2U3rHetMiUaz+nVhb1eVM0E1
9s2TP1+WvPLbgvyb4yCyU1GAVCmfQ8vhGbD46u+wyyr9hqVVXCUgFyVN1OCy
ijlD6vMVUyvZ+ngGrhdSBB8RFjSX8YxI+waHmyig0JngkQuUiGTG2zBPBnYN
PUEd2w2ETAB+p52UjwryvNBMRHctyc0lUT9f4OmmnUzvwPhiKnCqcnJugshD
Wmh/KpdnOgXd0RZYp8lgGZQk+y+7CzqOQp87GLLezm4FmWyNtAKNV3sSs0x3
AgyZClddriMK2JA3Ym0yccyh08t3Kwhg5ZG4fAZA0LJTJZfSy5jqSve1/hjN
GHcQ4KUy3GEFC0fhNTxzxSBE1u+etfW8irlFMw+5WUdgWJksgy1f3tt0OD30
d735Ddptbgi53uYW+M7xgrZCl3wHfMZ5gdsGWhX+ZDm0PAW9zsv6x0XWuMaO
Ebi5FFV1Tt9basvyfoK6m1LQX0/mUeIN3BnNo8wP/0KYiCYpU9XKqkJSQGku
wdq24hXHIEfHYfZ8bSMHAOevSVF+palDObj8KF9l1LYWSFBxcy6Xeb1Ivsuu
desIzcoAdJew12lBoYWGIcMaU+3ph40P3mvkFMxG7+nEElV6agvyyY1oLXWo
pYaJGam1VYozoXIUR5Zi5DouoChHLjgiIBfrAYCUi4ubnUkss7nsRjL9MR4a
/a543VA+haEFJ0WXhautUa9paitUe3g4VG5x6uXDcUnhG3iNbqWbZ6t4ulFV
h78PtV1g48R2i6Z9L6lMRlQxO/ncC5/9dn47nP+NRZalM5pBVPIYOt2N115y
RKie8JQPJyATY1GwqszIflMzI9r32QqMhwJLEXJ7AE8DuXioKcSBMhePU8sh
MnJ37sTAQbEcAA+3KL465GH6lPAvhF3JpQpwrGjVkbXWqC3ts/uLLx861xPa
EtVLp57K5jheFCeZQqVGpbiE87j+v5TZmx6RfRJRbJm0FuC6jWkFAyKl+nuK
NEadpTOFzP2gQKQjB+2VBfeF0LTFXGniZeZV9itMw9JU0yBt5YT+Bf1HA3H/
nOKtdyzUl5pwoMIkYD7rgXxW2+6XOXIpyDqPgHfr310/MvVGxzVSFvj0W7uI
jAdEn4IuFCdE2aDqsBRuTQtKYmwztv0lh6tWh6p9xqvUzplQJr36rM8H87je
/7z7xSpCLcI9+K3Ge1HvQKu88M1wjxY4f0BXuzxf3T9tCprL9TrEXr15J90n
ulD09CVlUFg8wzRROn/JDJRcEYnoxkkWZM7hqynOj0yR5lXkqOAV2q9g+2zN
gvsAc8dvBRSq2XgYnbpld0EHTqQJ1RUeX4uBxJNijglO1y19NCkOlVaBT0z9
ks/09yVAkYABJkRD2ilhtBH14jKLe/jpOvOWeAphCBNvI79YZ3lEdjicLdif
E1cDDLnDmBfjJf6BC1cHVbb7uJ5UquUcKQIww7UijbutZrdmStIhK3yrsBDG
cdusoIMpy1WO2Ugeobn0yk1QBBZZDnbj1hb1MOhStOiU1N75gu35XkxhWrRN
GmXVo/CqlXMJZHfazV9ruP+kmpozxWkL3sUsF1+bFmThB3VdM9ZA6P7WecBS
8m2emPG37KI4D42lcEC360/KEhWKJkyuNhvtuWl1xtour6hIUX3uiMxTj89W
hlDoF0aE9zA7yyjQCFucDXmmchZ5JTYbTae134C0bJbOfgVWugUybHA7ePPe
eV/8tAFV16YbfDw3lqhpi93vm5LpFjTkaeYpuFogvqo141rn/BR5Ym+8EjoG
fM+Ec99mL6dRVYCYTPV1AuTBgcgrM8czqlJjcPrGuRvSAYvRnCLsqgYBBueW
b8rAkS4bLDWfXRdE9QoWwaBwPdXN4ztFu9sk3qqZ/ymjmJFkbATZrL7FJQU6
lGwrxR1Ar702dxp+cNZhh5cjDoDyQWttyzV7bG10O4uPgCJW/VAT7WAJo6RC
x3NQ7TtgbOdT0hnxeFdXDesWF+ElpG0L4VXZ2dxIMQrNWTYscZ949YF+GO1X
cTofoIEqYDYF+wNwQi2qZSNvA03x2wazZEj/XiuR8gSN7tHXoEPd+3/3bgTn
1K9t2NEU1iz99ajI93q5mq3s9hIr3lM2/Bws7R+aMvRCfO39vWthDz5k8CYc
Qkd+A7j9ZMsYN6kgcExF4zHyROTfgKInudSVhz6LCTnteXjc8uvioFaKoBMM
lukMzXWZM13L/KT6Vm0VZU6w4KgmEkFz8R1i57BCUr3AvkvZjutof022wPW7
Mh6mgzC8B9gvLedfy5Mhl+CT3TlZFgt5wCGDUxRYumMXOFebExGHPW1wJmPd
LlyetDjS3jOc/D6ie4NTI8cBK33HCjT/85QeF2XodTmYBbisS+HR/g/psDp3
TYt4hAe9UhLqdEapidPUAxVy2eYg/AWFOUu6pvou6KbPL1wPCcHQ6co36ls8
LFkO2v6mv4tOOA0IABkiqUGBLU+bkaQQbV+mDT5FrNk4+zx9wSM8NP93BaKO
Z5rxYsuCRlioo632WijhyEu7xkCgnz9CFdGnHbbCk/4ogcYWhKf4zcUtuV4u
2+JDGbuzTrShFslTWZn+gmQPherq2SoD1UBrEHWy4GjzVEZgTtE3RkKPSE4F
2HfhYGTTBt87mLJ6ik+6gTnCGBYm0dX6gvgB3KV31EE/MJ6xRIb4atwfhm+y
czT0bzknqnSVevkf3VIJaeCtHZM02spjym+wRkem6XDB9MQiuwpf59mIQQjr
ZPosEmBQ7g/ifaE49oFiX8tGM02SPjUIU3/2LKQ6aJrzxsAGE6AiUcbVIfxI
6P9lE+jVc7O2HV7dmUSV39QYFvJs+1o1PLi5Y0ZYSSlf1MqZdxziXAeLVtnJ
a1DyOCX4kyEFXbWUD+jwkUJFwc116Q8FftKyAy8sIIwpLLJRUshzlHmP2fSr
V4i5s9G5j47rg6j5CLrI6hPHmh92yC5dPgrXdzpR4Jv7grHAvJBO742srv/O
8PWG+xtqKOvcdyWE/uIQ2wU8VOXX1tItrw2L7RIj34rN6TgkCBmwwwTnVJUp
q8W/ofZsuYzceK07FygtPBoAnHBFwDz2evdckmvm1PjXNx7/TuFJixcwT3ln
gP8pnoFnQKgajbcUTXWpw4GSaElaLvd2/O3hpCO51IUZ4NiVpkW1NlxtmPSX
x2SuebF0E1XAGm62hqPbR39nZiqgf7hmESuJvphqMgpKMnsWWho0ILBARb9U
A3hdtqJ/LIRsSLQgyqfQl/9wVuP888tEjmwscIBzTdRRS5AlrqPPSBFSip95
qS5p3r4hZwZInHwmAAjeadzkfy+H6dt1+xuCjujyR8p6VaKqHA/jTwMJJoY6
kIYhW+rZ495Nbh4Ic9zAi9y7UeYEMdJ5hMvXSr4oogpe/VJCv6rdLIHt+U+v
OrbUwghR58kQqqhQdR/j+jMTyzNGhKMMyFa6VfHDKOSdN4b0gHzQaJcJIZGf
ds6X0gRAMwkePs0RicTuY9DjeFKF3SVbVbuZqOdOU56f79lWJHpzDM9rrebe
+uT2ThPbXnuztLqOkJFlsZvRSx9luqM9yittFwh1gW5Yb6gdI6TF0zKaJqVK
AbWE238cLjDwgzT2fLiVEzxw6mU8j8t+zoVXso9+Y+lYlq+4nQhEO5ixqKCs
fwOwGMIcbs1sNM7fqI16DuBG8b0Pa/Yohjph2HY5fsg94WHKha9i5G7tpK+F
h4SSiKidmjD+pKcBcPOL4+7i7ELSEreOeWGtG3COCHuDHVBb0H4nHWgkWAFp
BBLBwgf9O8bfTRAdQpzn+BDIG/sYUDpD0gQh5ek/1qq1Unn1ZGYPbfbN8Yx5
8AmnmplbOICKhCczc5nuFMtg36V3mkHDmiXzmKTX/P57R/SiiKfa/E1bg/3i
YhQC+Xt+Wba+pYREkg3radNqWL94TLPuAw86Yv7fpxOGDPg+wq5bU8jq0Gco
rrqKZPjB8b5bSYqlEyk7bJHofQH5Kw2g3pkRmk0fNgHedeX6NW49MES/LNsf
uTUMdPkBwe90dLyLINrNNSuFR6uqGEUzc45dYOqYrW398VlQA1mnlFZ/jLDx
ZWHNe7cX2c5U+KX/OwlrpaknvShuJDM7/gAxQErmOJemUPiNElHnC7ppk5iu
3JBPuFNPCwJdn7OgZCTOCcUOmjBasNb8ZdFYgqXFaWS1bTijCSdAiW9Xn0a2
RAw+E8L/ArU+YuP2Y1NAGhepqxxeq1zr2WL2tEbvr+JVcRSWIi5QWYIDeuSI
qGSJUvn5RUoqnObPwNcDeHDHmso9PFA5R3yTm9EAsaHOurwcDaxhIzOB/LgF
9iNfYdZErWG/2HxyXA9p4EWoXi2wpSAjrSK179liSYYKAmGfvAyifZm3Pl9b
S0UMNoBAYx5FZTo9iCizUs/316s2X5WkAU2eyPez5bQ+QlEk0Vv/5r488GGn
jbSTxKeIuJXguncTrJ275wy8YcASv79Tj6tdEiS6h0O6y9SRkoyh7PVE5j/h
nDgEmBhF8jwiKcHFJzvQK/NrevowV8+u7eCPa1u5SQ3GZHI0cffvDaBqwLiu
5svx87qA5+YarmZhzrrK54N5paZd33V5QYJdQrrsXJxw7021yVFpDb56vzXz
0k73X4zVd3QEXvpuxdr+qFvWymqE4YELW0M9vVbAZ5NqFsl93EhXc2k8QE1m
3/csVn8gKKZQNZ/qbBzZCwkMOxVr2zX1vdY2PpSnACoP94bXpF1ONZkAYIgN
jA03b8w7BNtSoImGDMaFCj1KwZy7u1bKOj9pEBveJAoDfJMBxGcWA9Ec3X8N
HB8BMBeIYuF8WNJPP3PhT2nhaJeb8VCHq/dbHvWWlrY15RIV1yv239JpgqOi
clA89mt7LBI/62VH37hCDFZcrrZj6LU4ExbnIRIGPBn5mmaCeY9Q3WKVIytC
Txpw97UIt7VnYhP3Xfu90bbn2veDL48sZAvMEQVORtIL8JYmELhNbgJqiyTS
7vOk7gNWCDTobJgJ/luCPYoAamqCfiTD+4BfnHFgR2I53Zg6lQ2miietYUvC
KNt/rxJwkPscz2Z6tYo6/bpYdS72SAfLpzXyPBd1i553ZUaie5zlZMrbO5/B
Y+FAKlGWd20tvT7Tp72v6ukG2jEmExzh/tiynZgUm0tuSChMwLyKYUl9hKEX
x9AvkNA17ehQR3jbFZb+t44kra9dtfR7xY2jhIuKq9LBdXSmVQCI0E2csplp
N0raXKYT5RwuK+6AOxMvmQq/KBCmN21ayxAVIT3D0jRDTUKTMmK19JY2JEWb
p02Mktiz6xQnoKfuBGonoC9pmu7LShCsJX7WSnDgLYLHHnL1Vck2c9Fg9Ndo
9EceNLaCf4Ko7T7qtvbJv8eKizqDr+Kh0uf7Cj9QGlJOHXGDz4+iywv84X0A
dpwqr1UyJTW7ok29VPzyNM9g5rIKckbcZlbczHbjjhNC27hsVlhE7AXcjhzK
dQ7k94caQqFi1PRkXLeggvkd9DtBJXzAWdNEHi4956hyU5xO0I6dC338GXzV
OaFuIi69LaC6k7RgR1EhdUubLyjCtcMbnovcWogLOxL0cBXAtgESvnUqdi/o
QiC2y7HHIGLVIMqdJw1LQuhtfvNDnVbkiQnJvv7bxYie4aPR6KoKZfAQqY6F
L2YZy1pcy+YyyyCg3kqydqmLQ8lXXG19BMS+PfDlS+j8w+yNvAExdo8f/3Qu
5lWqve8MVgAzItPI6vdceGjm7BTMkc/fqBxekw22XfQdDsJrr+Kq1SgiNAiR
F+Xginj1wQDZz7+WIlHrdM5LlxZVi0azzQcsuuKrd/5yNY7hHeAWg+JL+za2
bTmUqRsaPxi5F4x4xs3ZiRCEurV66iTvQy1j7olSzcAWHB2lQzzxA+nm9z+5
S8CryK+0efUTpHHZ/qj9xrSv/PG8LStyUkPsC/5TBdQGBscJ9Ap6r8LsQRB4
1oL/4So4RTqXh6SwxlGZw7k/t4xKa84US+ZF2NKtCklRyzdkJ5Ih2wwLxulX
txfOGZVBZ/eiyhGjQTWyWJgkQ+ybUlr9FzioNkkb3P/bLFVtL9YXwennCXo3
mNV+UtwONeY9vOUfZnLbFCr+myqPSP1MfJl5/cQiIIkI2CEdEI2i5lRpDTF5
YCjpE8VqqHwMeTGHhhURhakHcTnDbdEDitKDjf9/qLHsissVGsWJwIioxDFM
RYNeiSRZsCDSqw6EpkXc+lj38QhzxKyv/wLqaVpNhD35w512WXpJLf6wyPdY
4mWrmPKt29uL5X9zmoiISKawVxVw6co3ndx4zhwvQ+J0gVLU+DRo0pZ6Aupz
69x5siYJedP0UP75YhGDZv2x3MteNt5V6kettoqWweu8CzHkAIHpBR4Iiel8
ucn/7b3NVgD6C2aBuhKTKVc1gcEsoawE6zPoytPVVHhgSMJEdYsbdj1mP9qa
WUjG09Q+Rbu7djYtXs9OHT8lXVwFwKajXTY250V3xcoHmszR6Q3BfnrZiMsi
rclqzFk81qHuvg+Fhpx+wizM9lacm/4hRD9CTXUpVEL2w5mn2IfgekPk7lDi
B1BSHQ5IPtuLe2Gimc8Q5iZ/TJG1dShMMSMttWRJ6S9a0c3+XDgZodt1sQ56
ONYIcgMfYkVWjUkY86W2rF4ziURl1jP+lZciypGIibGt0UKBjgvuWodtHrPF
6pf677bfVRoAWSpXEDBxY7yjYZ3rcq6D9to30qo6hsGdMBD13BOu91d/apMs
mf9JylZTcKZjOKMgOixzD/VeFSasfilyM7DTDLNPMeMEVtlilx1gVFaK9+Pu
lRb1vflaqvuMvqo5jw7XDjHb1oGe2ggz5ZBFrW/TXcGzP0n4s1YJcQoCA3tg
mQTHWP6/3dgyQxAew8OQ7RAhR5W2PwKUE0WJjiOY5HuFPSIW5z5oL6iyje8K
9j6wGKOwqvHKpNcRbpjeyYChiP766Q7vgmm+CkIzDJFLXTWWLKqvgzdUP4wo
totW2P0fkCevltRd9aEg6dl9d5KlpHPSGfFBdKCp+kvYEG1WU0ZhCoCPlK9U
KI3o65GQDPBPhnaNlzQJqfvs1cehp2eyIxnHIMI4tc7IFzPwKwunmpNCUYBn
fiFmYQcaZkWTMgdmJFsKfZWFFLZ+9B1+c7BITJm9zhKzFkb3PoyXUZXFlGwP
K80d8nPtUoSswiqu6hwF//TEOfER+DLAXy8wDqhL3LKkucAVeGyPKgnJKQf+
W/tIWtHnHkKrP8QdIyru2aXPfc/visIc60MHtLTVAz14VLwPMulFou90HCAz
55gLQ/BZYkqsaBDn6cjx88ZIVIIWUB2Hi3bpZUih7AwW2JmAHpUKukRVELGt
I7B6SaNnjshjwuXNnIcZ5BBuJOFQNd3cUY9l+a5bWNhoSo7MwFRuDCA84T+M
vzGINj2NGHXTjEFa156cS0dZJlcQTBPxWalBYRWxC20XHLwg3PUjibroi45j
DjQt0d2vd/p8yWF3b/4MgtGODhSNcsaz+O8T6SscJW7/VZQCcC2j2bYli+j4
4NfNiWtYoyT2p5069IIV7eP86xLU3m+AV30jqFtnAoM7Z3z4swdGAOUM1OhR
A80zT8zz4knB4fpFUKPPHICgNX3wq/G9TjJfr4mhSPDAmqQCxVdHft2AmvR8
RBQLaBt56d0YZHhD4T7TkMshzP8ANATByVyFAGkYNSfSCazjur5lrzjCfZ9y
Om+yIWsgnr1X0AHKdvhqtla187m8QkBY8Yo1HYgGC0vnI+P2pGIne4gOSR0w
nI3vg/cmG13h7wAf8kx1SA1THL0FSFnh0e04eaqIcbCd8n8uU/7b4+D37toA
E9eFK8LthgT1jpOL+0JUU5WiYE+gCorfqE6njqepUwCwpoiAvLtidiiIcFoY
1Fxc9xg+/GPVlYhmtQEzvoJoPBIZff4gEaEVk32Pb+89yRFAqYGT6QnQ6Zub
RaTDdwzKgWOiJwzGzR6HYJS3K68l4XWvw28PGboQIasSpFhlwn3GhjJEndne
AGdlbkjISDvXsOl/amNrq3Wm6/ok7v1tQIS7feSYMJd4j0UbLgNIrVrW6wVq
HApvxT84PA1fdXOkx8uGbww18ncOJ2dsm515pwp9uuS/suKh+GMgaY9sZ64x
VPRlWlDXQpxN8LogrLLDUnmTIJgCACaPK596jR7k1O6HmHUQonpB1Zkxssir
UpbhDdGDgSE7r0/a8+NjPvGf78sk2wLg1Z/hCw9jmPGk0VZfBwtI9Rw62jiD
gF5E2jCmhBzoojMYbPB11pUdJ7omcaeuZCUoa0Nmrozni9aZbZgpwx9sTuAN
Wt9UrZEjBGmgBpskgTg5mNOjSsHZob5Y3fuZMkXrBexdfi59laVZPhcF7SPn
3w1n1lXlNQ9nO3F/Yj5o1GXoqqyc04vRvd5L9DsXBxTjkmPKUD1K85AzE8hZ
WnvLa5y9zd5iOV81G6z+olC//boOiJn2xGXo5vSLHoJY8tgLMb1YTFCGmOKd
jV23ed1afioy40b6YAW0UPNyZKhK4ENnLZRLAy1N6AsQ3gEZV2hC4h9BhWUQ
/CEy7k5AyCnu7E5nztBrFwk3QCvYCdkrj+RwrR+xWI1pdkKMNEhUJ1TaNAn8
W0PCTChrrwl/0JjT9tmLx+3JIhsduxruv4gm5+L2RtLgedNiIq7UO09k0aop
7kWNfTKv5wEF/guT4lxCOM/7Zw7t/QrIrVKMjAGMrHLp0hja86pZwAXmhyri
qsioZKIyNo/9ypKY/7DylIyQyzzteZk/WMu6VwQjODdJt5pWjunm7K8NZXpz
qjJGj3P3FxY/rO1jaa8ryVi5JSl+UbLRI3LkWCtNSo1tqR+yQXEdsUo1xlLO
MjG3+F/GytJJeBAI9IrKxVp+JyVmxoPtiz69XhAIW/vzFPSUgXypvblUzVRe
dDiLowI6ENliaBJaPusVNoA+yjk7SDukZNQLFuybLZISFb2OJYV7A5wvMxV2
MrWlbMH/k/eD1Jp6ZQsA4ClzBM2O7qnhkYTTkTnSaKc3tmuruTgqxBFqX1O4
ZDb5D1KAKMKrA5FYbN4by5stu/3o83sFhsxjbOalwojKYvk3eHGQqDCI6XVa
/gOxrTQOFEM3vXcbyogVCQxPrp+4+wOyrnA0EkJKYvrYdRatmrcvK8NBAr/E
UBJ4lzcgE8UiffnQI8IUtaSpklvu+ckHLLzf1ZKgUPjAIMOP0U4r5bwCibvw
JDMmwg5kkwJnkQwJYX+rI90bfdO6RoEa0PEPslaNNvf40BECpDuAidRIRp5T
CTHvBW+mBCI/5u3PuxMW0tui48nNn84LDxDQQU/lftHGtQfLz9Ms/XSGU5Fo
9lK0MP3jyqGiRgv9qnUldwAjXUBS6eXqSsDlbFAKk5a96OxACpbNXQQvXMBg
D0fQOcTl6fqR7GoZPECjJe71EJN5QuYs59BJnZrMNoJxZzVjST5RRjjz0AZ1
mOW77+GvoWml0l/j0BCgNO8mLZo3IAnm1PhbaPLcslTLj1RD4FGybCIZJNus
TyylK2S/wZ2DfQeKn5N+6t98wLh7fJ3TfU4gBrK/uu0+4GLaWIbmvmy7IC7R
AF/ORUf75jyFDn6VuEFAuJ/SW3NEIgop+aulBShezHO8OQDPsnjuN7DyV8Zu
doiJ8P006+CrHdfoxq0TG2Qn8hTTRiUztIq1DhBlhotfqmM9s2fznAvwwC+q
7nJSielk/7a2MpBHipkLDeIpgQxTitn/deKMr3v/XonRnpm2bn3uUtb0G1L4
PXPucIYP+YOSumlJ7YXQ462ytxc3XryYy2xQDgbYcMPZk2XwQXXSLPscuEWE
6Nw6M/WFaWtezgOoTWv1YtesVcG+jRI5+EfOKhu1gSghHf4yeOYutnGYtjyZ
oCmKcF8hZB+Qkgymze9YCLk+Tvx1tzLXb/CcCDbQo1XFdi+knh1e0uFeESk7
wERMa/NkfBAmCmQHdT8rcIaop8p4lyVK25JZWzA+10Ha9m/hCtcSr5m00RSz
+xOLnYWCDvnqh6F5FpAY4ZitwJLZiYjsKouMszIx6R+r99ocQAmfsEb/xm0D
nlOBTqE8mPb4tftk8o59ueUTCg/DO9JhIoQ6FfdkmZA4SxuWJevmHdCBRagh
eSQKzvf02o4d3fyict1vpodE8hYH9pkqh/Sic8ZVd88fEkSgtgcunIDjUiX1
vRz3BxqqKCaggSeXiXSUFBSQsG5eMkCl7bdg6jiy8T2LVf/Z7TS3m/GnhyOD
MvD+0JUa/1Wykk/8WdUH0aybAq4wzrNL9i3J8dESN0/L15La35p59rNSajFg
3TCNlS3QysSIBrrDJ1NWEFcc/mE0g0duOgg8JtYS1DJTgDkLBcM0EOCd/5qz
vWt2rhgNf4Zm4W4NiZocHRID3boFEUjqWv+NTLesv52MWgiFgKeB+en8KwXn
j2lXHymsvH+qz3y3La8ZTyWXfMnC7YFxB1FAVVTCkIQMqocjbbJoZ4rpcaIz
/F5uAhqNjF7XuxzI+YFc0Z7pD+RF/WQYTLQh952Z5umlvZEepC7rJU09aCRS
H6yXpNOvSWPg8nlwCI8mBdveFm9wFwoxdqMsn1BJOLO9ykb93FYwnvqw8dGp
WuEa2snMEmtxIrsZSvQQgOsz6FV/Thv9yq9PihDitPvVb6X6bM40o4ba+CPQ
zJBkwqY1KoVHa5OZ35ir2VBULvD684RRhCqy8ZMpRaLkASViyGGyUEcTA6lt
usgaErsqbiZuGI6UDLyTP8f7vbcKlbRxDk3Dj1fLStDmaS0A5YuZSDm+Om8G
CXTOXu4WJMe5HPac/qODhtH+w/Ook5l5ofk2jeysSlUCeSElAa2DtKL/BLiq
gCP/dCtfbWjxl1YJYVXtDmHmwArOf+t50awxgSoT7DpWGgRFASXJIvgbu2o/
3nGVkAeI/R7C1TwHWimBRMBQdaoLsef+idRLrliLeeuMgV3/MEfm1D7/yA5O
wnA2XTKgw5gHbewt2NJaIkHhGNvnCnOawqfWD/Vl9V2RrcF+6bOCaBui3Kbs
0tADCK43uNxlDGx4uUP1mHsZtyBu2xByyrrz/K8De8114/tpYqj9dvUYE3Hb
nvECACkvRA8DwgrsLTcks4/jrjqwqLzahDmMvVhgiu0ZwqM4zOS5K+UTZqZG
yOXKLMh3omAlduLpQnhsmU6hRfgdXxRq4AxP9Qn6QYJqWPprbwAkKJQBWN9P
2MfRWWArfQUO7xmximoZalCqkR1/0gpd+YS3BDm7DxY/2VDHj8wY1hwlzmDu
2uAfuwHI0AA9rzn7fNUoo96UEgWv1FQN3DNADlPZG9osJT9XNJt5vp+u6M35
BOXqWvDmiY53rW1O/EJQKQhy6D6+J96zWGIY4IzT5tOVEde8LZghIGcr2yq9
dKtC4kHGyWrhBgy8waMpwNqnnb934XpldYlsI+p90AseoVnLUdhdM2l7+ETV
3LSqUOESjgfirakW/NRoOUW1xY2r4nSMzh8IprHo+sK0w0Ehal4Hkrr2zn8R
wFAVeGYKV4bIPe+WZUxxUaZtNxASgS9lCc9uxgq2SuCjUGO/dWK0VnryoSbz
BfTx/B3nYMad1qNYFozDz1MRlhulkHDwOxJd5pXsBgmbLKlVpL/ljEwbV1jo
KpS2T0z/lcPk4iZT6C9015mydxbO6WCZRtEGyRp0bOVFJkgZAQcmflqvWpet
twrX2qAS8szfluxUQMUyWiHA3rBDcr5Vvuy4mU35eFvxz048K0dNUOrJVUsz
L1595WvN1ZPe4xr3tIXkpnhgCfwO41DOMSTNOI0m8Mo+TWnblJOHM7EL19JZ
Cd3LFiQR1skDuzfc/oU6tO9xjjEpgOyvIcgO/bpArWFtJ52C4shxoFUSHWHG
GKnmhLJkgVlK8qR7orqGofy/uGyuhKYWXzJMvM71NM366dWFq3Gq0fAW6V0i
P5OQoGSydzfVPFfB3jnALwPI/sqVbISP/bi3xfuvlfMbSY6ULSp1bIpv67Yv
Pjl2jpLWNqx7gdA2m/9BC9Cn0TpTtlDlmctwDr7/dIGN1Cz1NlwDctxi1pwO
Kb0ii/pZe3RHhXu5ECVjyzTCaGN8mY/2HMu9gTTsa9PRSS8ciy8UBlow0h3k
KZd1Sx5lP9jrHOnMevvcfvikyQldfsu8VyWpiAZuti6ce28prPFXspawSZUq
zIvzqYhQUyzn42K+sknL4hhtuN5cUFO/UyyOfn+kYauIpGJ8PAV2k5akUzs6
1R0esWaJtVm54C6lsjRicjDHeOHoA1S1or20ZmUstYT8izFHUfFz/Lf+6/jN
G/uTgMogevOtGk9hAO3Qc3IJET1CfPP/5gguOg6nbnbRnss39KWByOaun+SX
QSalYLbc34cuSTnnK6/4MojvwDXoVYmFXNHG0Pqn8Le8bAxhll9SfjrAeVNm
m4R82q4hi56x4HXA5GXmE67iJ4nL3Zo58zzts5FrkFHRDcmS6l9tFy4AsDe0
iY3DUM/pdnYmlh9viGJUpkMf0jiVKc111ulr3PDmKOnANuvCcDH3VG1pFQYV
rQPpqBcoFCNvnKLIXYmSKlk1cKZ0MDaySm1Uwlv+oNGG3fP9twRzvFfbN1Z5
f4muTmeekmy56Y9DXxizrBIdtsnJwJo/Vb3SAR4WM4hwoJzBLu+uLtO+xuIL
nSXUtIHSxBtvNycQLhs/I1s/jI6I1Xe/9Bb3ONGa3E5pz+QsAx8iMknDqaFf
zxEXFu3ylPzkNB1/3b6JtcHIfA0FOF2aH2OG8TTgZNkH5Mu5isXS1K1MiiLv
4l9eLLB4xXh3e4/FDzVOEDAFt4V9R1UMqBnlA4mlMhk9KDvWVHU/NSCiByHM
dIO1EbDv9Z9K20287ZU9mKRo3b60zmIaL0iez9sSIIH1+c6ZnIK62ISTWJMh
ZA3Q2S3ZfeA2cdgorQQojEHgtPaRVBS9dr0iDS+UM5yjQcKbBlS2s0fjO4/f
w6XJaBaPrx4Tsez5Q1dZvloJ6eI0tE7mqR7PlBDwQQlYuzs9irI4m5x7DpJW
FJnmOBBbQRwXa4elC1kZloREreumYI1dMA9n0UR/8Mo7z0KIw8uJcQuZLMQC
CAq8wIJn8vMDsg03D9nafAQ4ZAoweGxrYn9hh4yB8DKB2XBRzaP0ud4QQ7nL
0ukBotq8GN8y++ryY5Pk3lseYLECHRUCnvPEUsQlYqJzVNUamR0VG7TYYTNN
vzMcKgn5nZDsSIhok/FvpT8TR2I+i5rzoLTz9VIUq+kFSNRvKR3t/5wco2s6
UhrjMwBE7cLuoAhdhcy5bJWcD/oaQOJffuf22uaF8dw4gtnaTAgmbTOjkgw8
DG9F8ovAsajyjSp9MSkQy2Jh5Y/88N2RmHBkkDNRAgl7Cjo5OUTEjviohr/k
mWzrDZsOmReLP5aAPiJ8f3qqoTf5ZXWOzjbrS0H8nm1Cx2tokSSw+ruotv0O
2U1pMN+NRATWxyU2UOsktfQj4AYB93EE0CWoe8JDuLc62qzSVpMRvJL+aT0W
m7+825i9zRgidjnDPKAV8coSC3QtqSTb90M5l2DV/cXxOJY/bCWuebR0hrB+
7KBHYzL9JFkWLHr5q70eeNNxushDCTVWeDAIPnoFsl9BPwCgwf/pMsSQtKIW
6Y568vKYUstjOnLwlxacjC63YSI4rUQNfcsIz//Um0/zgPPPo/ycmyhn/0U6
NALzcBtyrX6mBtyVzlo5nzBJTK4v2DvU0JemmQ9rFi5CzagZZq1XRlsFejm9
KzQVJC41VotEB8C8XOzdV/ZS2o4JH/E/tBDG9HexYrxuelPI5TrfhA60cqws
F/amgVV8SQ4xH8Ci+W2NjPB5/BcMf+kDu2iUYC5K2Ch2ft2RgptLAmGkoQkc
ioOzfl7hKqq1s9Uz1yFYkUwJoxrWyAUD1JJVuYHc7rgjvs41hR+Xpoi28hB0
4GbG4Bx33h6rhSv6hdWQuhrxZOAxQ1j+PiEYng9q4Ao97G3Tg7XwgKOAmQ4M
t/FHNGtQ70UlXaIxIxbPwopglImSMIm+kyFH1lStPydISX4W4cWyI3m8OyVG
aJ8Q6PPLzG+CCq61bXkrpTTsXmL/haJM6MUvVbCCq2IRGpJVT4Vc96u5UqcU
pxfHBqtbONvC92Ahw3x5PphuayjQlxQrYbdURfaHorrcOJvW+pn2T6FavLzN
H9rMMSgNjZ/C4kb5gGyn8VnbLh5gcl1/EdlA6vLoqStwyl6gU8nSa8KkgLfT
NCXrHQEXYsPh3c4srMqwzDd0LdccEUCbytOHDhxqkSPl7wt4PFYTvploV9If
BB8/r8wlq1Ekafid1MUXgMzKsdMWja5TysVjw7v1kKNnoCKvC6RCadh4n67a
j1SX2N0MdCNMXNXmjkx84ro+/J9Mdiad2o7CZ3QWYr3ykQTikCvzCgLatkIn
iXanBC7CCIrgXJhEly+WZ6YijBlntY0JQQPC85m0clffP+mXAGZESKgw3wss
kf3oeht8kj5EbnUxNWX+1q9qTgDml7WjslkKeQwvtA28hU5pGnXg6AuyE7Lz
RNV2Sg+dCrWZOc6cen8A0RGcV6q/null+dW7PAIlXSSfAq/LfRbGIExepxSY
1macWiBXvmAlOAfVJK1II7/ijBm4v3R0zBUzhFy9mpy71V8VcrSsnLK1JL9c
4hb6KmNS/lrEBhDG6iYEd2uv3l3dpZY/jpPP9WeCQgd8w3eiQBIPHLLe6fFe
qj2HYM3BiIjeWbzQgYGY7TeeDeaVIY0ovOBfW679iDtTcrsx4QC5NlbTYlrB
2/27uTG3JkVuDrKz4+vnMSVwtl6TBSjpua6V2OYm7UsuZyuVB+bKXXivhufA
UdPmSMOl3yZT5KacShtZIiLtMRDmeC62yNdKu4Jzo2L2VEpVS2+Ievi8VQne
1XoG2YNq1gPZ0WHiBZd7Ji0jXmPtgmRXEPacvmjjsVPXWrd9qzDaOBHu5hOi
hYT6BCprRkOFcH+b2JZL++Ek2JSrXsukw9Ei4k9WVpK55OlCU/lr1cqk9YCn
OMY2Ybzg0Ng5HrLTMghlgh3FFQzGSTmVf9dnmCqxEL39IRmxCA8pf6wI3m6N
3jCkd0ZAmMHzZ1e1roQvR0tbuyH9/wOBDCsiqF05fUUtiIx9o3ZjNAy8FIH7
erRshiaw5paymQQwlJ8H1GgRhaDNb9UVJk5drzxTBtlhMVfVPk/l0JxfeIJ+
y3r2BkEw1rwYm8N9wGuZ6pXN5vQQtjJwcdQOzCXU0c9JH9Lbw31NiBlj1soj
t+fY1FiNEgyPAImRfwyC4nkJpj7boHYBpAraOYKF0jKiB81WY0nd6Is3nUgV
N0uvwjvKQEj1SLuLeHVO2x/cA9MelT24h2fkIMeMk8ke08jRFOkjO0KKNjCR
gRcYGa9EtezHEPBEd0uzJ3utcKd+712+cahYE7VR2na5miTi0ygr8oJdGWoY
m3Ld7wSPmBEMoK/9Ggp3JDDldMJd6fUfHC4kfYxtlPlIyNH1QLe/u9IycZAC
ld++t7KTG32BRmnjlt+1z4KZrAm5m+XlvYhzIl3GmHxzUgxcm7XvC7bS0q6v
FkBECYRmZJWBHOGUhgQlqajghz5BmId3AeSdNovLvdAdcdlRQtKDcfPgX5E3
5YhujK5YTFvKt4/jyRaWhqDxg+MwSYKs/GLVFsTv9Rqwclme3tsNSw3uEYna
4kHuagYv+1WnlTIkyf4SnQ5eUkXFjBma9CWqZxQk0/v+kXPgUwKdgoqCgrGV
edMdYfaYaayhJnnqvhCy0+6OcbLDciDE7GGMVxGDhZiZA5VU40i5JH+Ny+Jh
5R4rfiDyWvoX62qBNLpCKovtFPZZR+ChVzOSLo4lA+h9iIyhYR8W4pYP83uC
6UVrCiB/SqPl/OProbjTnXVpjNTcgBFy7H+MXniAyXu46qhLU2zaqRqxpffZ
9U/h3WMetTnq09KmX7AtUxPzqf/U9eJV2cUNYapDlA33ZNUz7vM6U3scewi9
p0apGYdcI8+IqKkEoXZRHX/nUJNeopGULSTOImAS6mrEViiiTfxhPKIA0+sS
O+f2y7navTPVaiUVD7AyS5rwX6//wrnXAa65GWR5CQIy8s7FjtdtY4la5XSl
n78u4lJixqfssCPh3t3HY0ZWgA5qUPDVKPj6c+afMZ+mFQOUNb/seqQSPtLi
pmFYvZ+sajU75dZB4G1Tpc9Zo8IoR3rogb4rWtmaVkX88Z0ZNinQaiUrjFU2
wIr9WF3s9H805nqFpPWhBGN77KHRPrEsDrueRb0aquLmYQpRdGJQmPiCyfXV
jyP5ClezEeYwjBT0r19i7URI5OvpZVgKQQfyMiQ2ykgnMPYFHbi2Iufo5Kwo
+6ZSLuIAqk4Y/bJXnOVV7DczSMssoFMrG+twhWpQbAL4uSrgJ/YBbKnSWGnJ
ZxZ9VqZBP3AFkWHoaDnImPPxA7fOTYSRxkT8f6MFOVdf4tX94GEVhcRdvCgU
Lj5O81sr4cs8fK68kB7r0a6mfHRJ87zpD53iI/Xo8AIgmc4zmD4vxRYOpCcW
XaXM4l00SlddK6dRKg+hR/cymHVEujnJAdsLgAB2orZUIaJhyEqabHmiUa0O
2MpIzU1p8hk01mPYmEtrA4Y5EDrSQDBSdZKBLxkutdssq6AOl+X0C991d8S+
9Haxs69M7yd73LsgBNZ3xGqh84teFgqkKtJcpmKyF6qIgvq6VHMJZbFEkWb5
bjhc6tH9bWc1JJrbBrax1ZNl0+N2UK9bpuRh0yhPo33MinRQKQn79cR//KSu
sktcPgFzM9QzB7TeOgxjjH9Qy1n/5Dc/NwoaTKlXZOhPm2RXz3n/tuhaYqy6
hqgyQx932gD5aLi2ukDOapxMwJ6X1/LWfctXFBmgvi51q+hKiqK2APm+Sn7G
xuk2Uc2mxU09+O3JWV7B/gAminf+yrnK6B5N2K7hya7Uzq9IaFLqbaa/Aorn
/stEJqXJhYNYTv5gu/HXfUuQUKPUS01M0EYu3Rw5IrUVSKLVN/NYbvcSFU2X
g2eWmlb3XHyGRuw9EyQzWpCwDn/mdBfDR5046AWTet+/nJlvz6NwBPiUkoCu
rhYPTI9euZp+8Fp8+l4BEOK5ZHmV6dutyN8mXnhlykrlnsJlrT2WWhml+xqs
Hy4tRIAzw6jqOtkfeLl9T83tHApsVW8ROUcs+5ZyIy0HRf8W51o+EFN5PMI6
NCmPCmPpC0M6SIv6LCJbrNLYx337N5OUkqQlC8fhIeBWxGOdg+RWJM/hq3pe
o0pw1PsZfR6yLbJooI5heusWFQvP+sZMm3+ELabmzRFhv39R/kkUJoBpD9iE
bqmHJwzinp0OUDpGOfRdxDdxnb+oGBS+9nXatOMYYnwjTg+lwSjzL70KL+90
5HeqZYBO03rGWBSFQqURK4GHdvW5WOT4Kz1cCTgnT2P6jEulMyJP+ySNAZif
iOVdyuXffS7jp/YUswpEVrCCtKZcp7UI8uv4Vdh6CzYDtj55FVaG94Z9xK5H
uQf9Xc/nQxyYLwtFgcjF+rYfweREg2NetFgeLolXLvKqYHmZ6m8yLVC1I+MH
rIn+cHpGZrWJPNHMyNkWTd/F72W1VfmWFu1TRI93u8ixpbsG7sR5Mwb3Ys25
etlMyEOvK00fcj4rKcVB3dBDyc6lhCGxZto7e0sY9sg5EzLlH6zmCouvUEVL
NSFiAIkwsTOvCS8TNmqx4hCth8kK/+FeF11I4zydkEE0ZyUwzO1U2yprTWqt
RrWIkNzUBsHTZXYxDgLybK2VjWtuHZJlIEuIUOyqXrrpjKERwg/w7jYRPS+F
ve0BpVaX/kKFpd+I75Md8owhagbFZLFAbqYzkF3jG9d513E/r0sT+8i91hFO
D1+L6hHhlp0eqoqbufv9umAWKXHhiGAd0yxcE5BGx9bRvNJRH6X1RDCq2rPS
YlNIA2gB4qJIMqew98joAVj2X50qdm+zN3R8hhh9mTz6DYOWwNFPY9b55kH8
hMBoE8vyBAqzWe7aoqRPj2gNhFk2AvlfY0vi7WJOtWFORAGZmttNxajs7FeQ
YcE00HkS/w0I2ZxcS9Ome7LMw1dwD2WElvwXOT6khsl8wphn9vjzfO4D6clI
4yFKUMMgFOM8Xvlu1Kq6XqET/LPSUiBVO4brYI4HOcbhxYLO1Phi4o1wvEbB
TIv+kRgcAXvAoBnfOV6V8u4rT+u/WjTl/F41PPR7zp825DbiTAi6LUu48cix
OCf7fZOkHaBgjyTSIYjjuHs6NyyqPdr9JCopMrBjqKFy/nQBdI8GhugOgW0f
yCKwHvGTS4Zm92O4hbpV6fE0EOQ6Z2g0z2/lioo7HdUS410eaccAoJO9jrGC
NSYpMMjftXUguGqXs29dEyay3xERm65NYm2EacS+ZhKOrNCw29xjpOO2CfPx
tDNNg/kuw9fKscnmH4Qjv7FIkpNGjHpX81VSerGjawpqCz98XYIoeR0deUva
8fHCqVLxsviX0LCKhfmb4AQoihvtbMdN3OIX5IvUWPGrbfuhCkIXF9Us/kGg
eutUxMpu73i+3fktOKRsK75nlJFpLFImycHUnc40eMIBk7LuTRNBc8KT5LJc
3rh8aCBU1eqgLVl7eA5G3qxKoBIlU8gDNunVSniulKtg4bPS1KASH0eNKoLt
7yszwpL6DJLZEmGpBINAnixtWOgYOQZhmq/z0JoRUX8SUZ8Jb/6S6MUN8TCQ
eRmCKas068mUiw4x+B8rBSgbV/Wba0kuYsrv0+MU5AQUy+9Hb7rAVwgdFcBQ
o7M64TO89yxh1OFgSMoLChSXf077cqBVUIZu6hRL8Z2U4zhC9aDEx6D/p57h
uy8NJt2DxF+gkQYbft4yikMIZqXZi38blVWRrgmMeU4ELtE5VAze/nuyWLNs
ZSXg8rRZtJ9nDwfwKiahwgn6iNnmNTueUomZdGX/xJ+BzDOlGZQGWT2aM4qK
8r07whV2dVSjO1jV0Z+N7IZAQksCDBYg0N0wSK3yRjLHchf3YnrhqNGtI+ie
+ukCR2MN4BVe4psqacF2BZUjvzy5HtunXdwQuS+RJLg6yho3UIudzjkbRewt
gn4yp+l3/wz3YGVX3XWGGJiog9aKDroafPw1ibWNrM9ste8BW3qEHpX65o2b
W2yALdrSd57VX3k1LHZ1PVxCHAq9BRryIKXTtRpB2VnxTL8zQ/g3JLUVmQ/x
oEyRz9rjSAUNLWqdgPxylRKRQXd5WQxrh74sipLkX37eqRog9C0hxOkF998S
SNdGWFfAjUZrVFPgchRRbKoF2jDkE3ddVpjvk6QkxwocAyJxb3TZVc+Y546D
mKHxa3eoqA9ZUEmesOke0aHspNS8bJBrIFxIDxFb/fu0aeHC22fYl5NJq0VT
MGuR2MhyfBD8jYNaNg0wEo25XdFXKiaAEtgPIqqpfGeaHXDHc1PK/sNAkphp
6UYYxnRGLn7CxmSNEjJcgkqtxeZosgzgcK0+3E7NnB82yYY5aAIZ4Ja9n7cb
y300XqOui4hkDJHeXzQloXb9fZi+7pNNt6tDrPImezBjEFadrx00lG7XyaIB
VlzXMqluc7FhaAVTQlJ2/scClyiM/vGfgJnDPDGZZnNlL+5lDPcCRYctg9vw
8loeumX/WfPI1V3OB6yIHp87O96Z34Jylk1kPZfLLSXIlQRgSnwtmRtBVGVV
561HfJJrU6pi0rRR8LHylqogtcVq6OgHy09ZaRZh+Mpujpaw5aVJ14DmntVk
abHgnEhQrtLJ21XSF5x73f/2b3EQ/JCdJoyGzthqu8aYdnjsKSxB98lmUuJ2
ikzh+5weDlFFq/NQ1BhMXho4/rjq8mEmKZ2LEItKvT2f5sPPN/dEJkEEXNdQ
2ELsY3o9T98QvGHiawz73oM2Echfh/wdkZT6IkR29AipKQPgeEAU4dO5YHox
IbuXnt5S12ipMCjR1T4F/oOzRVxybkFpnmEdbNZ2bEtFmA3W6D1TfZDKKROH
a9Bf6rdj6XmMEzZiR8pQKTzmr+gxuoMu0eCZsBMrbSnJ9OWAHdAwgRKt2QB3
1Eb2O01eRR6ZN+iYMwoX+ACezjihEJSNVg2jaOmqytcKHIVhL2CceP44kBTA
RlyYkd8XzVeEhNZQ3z0J4iFFXEed4s/ql5dYxN3uUpCi1EmBR6tLVs4Z+uUz
5faNstwyhhFjMv4r0L9ug1P/elkwKMDfpTGjNt1jLxWfgza8i7711EBg9sCw
wldjYSbYQxzTMDaBFIkFSc/kLvBoggaEovSkGhQTJSG+dnpPufXnbDXtQMf/
RbqYFBh9zhuORpyEJNwuvbq1rXGXL/SBaqE4/ET5w/AI2Z+HbqdX9GTHVHM7
RtYnqMseKCNlTi2MS4MyRgX1TkOxcG/0npmoZGZuU/LXTOyJ0zlyfYoDYqX+
VihcolzS/5/TJP926Moxh21o30alaz6KhATV/m6bl/6/86p4KNnZ1lttF+j8
CKnxBOEAsCHjHjusrL8bNJ55vDHEo0Jn9yiBq7Y4rquzKQZB4jeIR4dFH6bf
/xfOxiHPviTRx+WV1zQfXdMa1HvRXZg/6gcM5YtHh1M2//QxasQJ66T3iE8U
BRrWCZRfZeVtSBiC2fSaGjMZZLJ3gBLCuEZzsGJLNcaS2MHz86hiR/+tIb+C
Qf0HFQaQKtyuNqlw+hNjAJGC2zvEtASHf4mQ7xQcjz0F4Rkrv8X7DxU3iFS1
ZQBZWaqwARqz6QT11Ex+qZtGH3GReHengNGUejxzJyIrJot+KVjjImbusFK3
nedrUa33pSa6M6jzDlfwx316BJSe2JVSqg8m1WYA/pE0ELlHOK6j6IdDydq1
Wr1hLa/d9qZKyfQ5PlUyAERoQaOSy/RbNgAbfBn2ytdupyimG8p2CoUWjgBh
GDhJSfOWGMQJ/1Fp5uXYlAcoHq+zpIDJf7rEZvvUVdorr7m8MiEIz/ZVinBo
dYkov7MTTnKGCW7/Em08s3A9ToGD9+ed4eEZhPZhmxpVZ+GF4PAp/c2yNVeU
pRX01UpxkSjbnofXftgm0jGnivrLvYtE66Jf7aPBVnTnlw2q3P8P+RWDZ+m4
Lmg8viCtMj+lO0xzMvIMK6BQuj9MxFBW6JDLyLXRBwTl2FMtzu3bRUHITkVq
2oWou0Qlv5TMza3MhlzCuDRPHa6U2jparWbZymZNfNECaapI8fA99vcsHYhd
fMf5wF4Y0XrD7AMuB2uJoe9/6ELdjJGrpp7Zzx4wa06toJ/L5refs2gaJFsm
xiNUM+jpw5/cCNPO2krFsdGB3zQf7c1tQCLynrXcrLvl/y7vw3X3X+6WJg6g
vvEXweWpkNww1VHLfaCKYO3AYlOhjXzbkHPccG4+d4um1S+VJTNy3dM80b+T
IYUHJGrMXTOeScS2+R3ffMdQi93/qWPKTyII7HYeJ4IfW5NlZtiisRebwzgQ
w+XHUznPLYBPeiqrWPX+o4/Ef8IrDzgeaIxH0ziP2lnwmGM64AmGc9b6FJaa
ksMeGVa1sVdr+jLAEn7kgzMU1DcZ8/s1vdXEXEPhv9LKiRcHOrxaBzMVxrZj
vgmyPqmoxw5Koz10Num5O2pG0rkNTpjFVwFaIvSo9s6mEutigau04otWb18+
FW2p1K6DhWX/PoFYwEhPsfuNBxXHQW0lrGIXSNRiX9w4prwMFlKljsyOMlUL
QOlV1r/wUVm9gj/PMsefmTN3Fw24UpvFTwlgReTPUO6H2jo39xzMWdSxJH7c
2jRkDjqS014OWtvdaI+UrrmDBOoyiDLr2KqUc9TVaZo5EQmzcBnKVLxWFzoZ
O0bfdhFswXKtb4gAiPvPpCYti4YbBb+Ylv9x/jovyRA5aZac69vgrFi8aeJT
B6fHeZEK/nr7boeAbnJ+WTyL0FXG2jBuz1qfzvqnDWoqE0AHwILE/qIWthK3
0XVaDWLdUV5zUwuCjdqDYmoju4zsOdJ9nEzgoH5SB92Kdl/PyrfUIGE5MaSo
HmISORzfaSKFxgccYL2cdg+Xaq2Px/psG481+f+KXKCzzxNenSkN6C0OBFMS
mHvXc59vbLgTNosY63CEeP+JOdyd2UJEYgygHna6QfGAzo967Ml+NAK7jcMX
ZlCb0jruXqqd/FzL5fZ3gTeuR7Zajc66fcbhIox38pV0JfTghABjK5FyVfGy
o+tsvadZEtYffJnngHGCziLWgzkeSXu/XhqrUXMTTh+DNqgQ1IFZyFKYXg45
xglMYVy6tP2nxUtkgo3gvtQ8enM+AJ1mHrW/wIxfthMkbSwt4GEx8+nldr6z
Xej9ybn1eypPmNrqIIDPxQuf/DTss2yPBptnn+Bb+AhaKfXEiBGlWVnvyySS
lXVReT9WlDp9+mtiysAGdYOtvjl/WtLz5Z71whQTvPDviW8c60roQAiEkG9m
7k5oeUC/SlUmqydeQhCoJQD2LaUEeH1ftvAC8nL9b1OTdL9EN55LNIl75Ly5
+Sr9NHMITYVC2xLxNkf5iPEPB2rTTYR7DtN51FhDssi8lrCSjgd7hYu5m71S
ZPgdCf9ZqOjPJFV16oXXgbhL0nrBHRRRSk5LTAw/xdyppo9Ntz0hPO1zbB1F
Mn/XYOQQnSzbjHspnLOdwnbPOvEw6QIafK1gkRd170MkDdcnEu30tKEHz47G
3AgdDATfobjYA3XSld8z1S7L8l5yogFAI662qyA2hE45dAsdLzV1aKeruvcf
1cFPJcvuCu+3ok8h8kI6A6EA1qjAak4icmF/KYhx/sX1cfCDEJz02SmLM/Nt
DjgIiHQXjbbZ69GcWJl1ZS7M1cacCwEIzwZ/hpRMkFv5rnHYZGrTEUqyoEys
9cBSo3AE3ainlGZTBzoGvEE9EBYEq7Msf62lmOBqDzjH1RHhJiOsDXVOF+/A
V8WV21kCcOYg4toptHZPcnyFoHxSd9PMf0djK4yfc4cG/3kyU7CgYPIT2Mpo
6dAC2i5/HBWH37RNcGEeVYsMa8kwasGO3Jz7E4L4XCjHvsWktSdctcj6qRLd
CZ/KnZLYEmcC3z4UPlxaWrM/DB9OiSXC+DWwWnwXoHRZxKbVl7zkHawO6YhU
/jItGs46SJmE03X36JDyt2IOa5Mw1Z1LwbY285w+MuL47NJmXe/5cECjUKiM
WPAOUFDgmyyx8vQss5PLUckk9K12xqoYSz51RX8rPQykHgEjswianhT28tyg
AqGOJ+Blb1F0xIqHGDw6S+VHm1xIAx5S+EOZEwyHZNmnbI6Xk90QZMQvoypn
/vzabtGRHoH0rOAcwkfBC25aMfoneHKyl+/XuJJgeq4mXk9q74OhlZJUXhi5
4LVxSRr+e7ulgDVetvhLhGYX33K5G/PeRX612RHSRGJjgLPzqCIs5+IOqlj+
MQnXwJDqqvzrFAOrv/UxFCM7QobnXf6LQZpOeaKExtESiOAUaczoaNZtPyfa
lQMAEvccfAs1wTKcNTvDlEwZS6N6ousPdWoOkbznBZ8YLpv0sX5QLLtysfJS
C+V055WzIG78ch36ZgrmOSRGtArCNeucXGNSNnRzmNEPFDakuqH+Tv7Ndnc/
h2C18jEUBl47cozuvLVkiFBgOgiEa23myfZctF6zpvfVP5WLxVkOnyYmUFjn
aCuDGSzg2+6CcwuoFEO5vYXuV5ewUVSxU4/IjkgOXkMIYKwJMsZKFc1KLOpf
0hDU8NyXNGbEbJkn03LAEbXpqprFojcgFAKO37Py/hay/QSQfepqChYcb1Sr
JBB+MIk7kX4EucfdgRc1BWGJ8M0B1DtPqyMM2iRee9Kj9EKyY3iim77FwotQ
SG403g/bWsaJ2sSTa64ADfCaUD+Xl20u6tVuzaGZtXpN5/54HjxqVXxz/5yz
+B9nnb7STBPR3EI+D2qxGq+ioyPqwMTfqzNbjAevsl2xnLKmIGxpYpWwv//n
p5thw58AWOZCuiA0IJQoMvThcaakAaPkuWJYrsFWsgsl6s5CRhWeMQKyLJFa
6bw2T7kITjUxFhc0yU9woM66yTymYHWIdk/IR57fvDTsznUeyRjVW9glZtNI
2xk8hXKHXKeyG2gHU+vWgDzMxR9rq2M23odiCmBGsLwPWjM+6bZZZOhQ0/7s
2d48CADqq5FjnqbxLDt7jxk+D8E0P/5kryAFYi9d3Qsi6CbwbGIo3kfB5cUE
1PWPTqLGl02JFjWCSewQwx8IqGBh9nnSmFyaa+o423UNvahRb+pv6kJYN925
VdADbJu71WbTXfuRMgkUdayxic1xzJdgELgJwlA5WaLCcI0GOGKok39k0SM/
O6AqGHXc74//qqg8GfCKT94NAjlVv6OY8DtSMtBk992tBn6fjZAKcNudTBJ6
ty5PjwblTbYPq6DvVT40SgtSnsnIESMZv4x5SnOx4nevuI1+buSQoiwXUGta
R+pLowYjEWg6+W++HabYbfc5xi9Co9SQ4tJ52ec/QrR3SA2EQlUhRyRcgWx2
O1G1qyLTS7W7D997B2QOHIJ4sl0HB9/zQYXd3qT2tpCDMVgiQnWmqCBc4QD0
RSxbmTpJxOKg+UbV+CURkuEUbVg8UrLANrNjxAoT+2aIHuMr5TRXfaHQGBu6
2InBJv7B8Pwy3dZtMNHtK2MdBODzYyOfG0zIJTiT46ZZmqUUMo4MXysdTEIM
s6jIX9+UFvQRn63BrCQ0X1jvuqzmVxgRMqSl8TkT5snI/vSI2GjXHkR9+IFC
M4Zgp88dDvGvgQBA+2HqEgDKY5fZwsqtXCGTGBOreDT4Hpm4dSDfQHpiu4pf
3UVuxjfosTuVWs2hxKn1ZcdeW/h34AS84r5SZEH60IQVZTW3bOnDgHroof/5
AzoBxBDBg2tZNn+WsjJeLixfTOYDGCeP0RYuNO3bJ5XsymAURcqBKzHnaMPf
cFJKXwZgL/gLoijL8W7XGbwDzojHanT1e5FZ6qgxxkkXude5wMV9S7qfwON1
fpwFpTEPwZc88zSitsbs+62sp04cqK2JdjrT+HwfR7VFLyLsQLV/COSPPf9O
qBFzf2Yj7rHOsWY9gx25451Y1vdDfjijKsz8oDYjqZ2CvYQstZBdhmpxuMzz
WYwoFEMXNONCQZeFy1tSXSr4NPEmwcBbPQqzux1CZ/9d0O493CxojhJ4B4ym
3GSq9EGnI0O6hKBEfFKI81AMty+hVC3kX070R06prfIBOPac7XRWYjHx82iE
NHqfFnCww4dc1GKYAd3n7q7HX/wOIIQGqVyvlkJS3LLNpZyTicVNQki5MN78
TISorzy38TxBeNhB2hpByjjsE4fz7iDfyCOp/nMGVXRz4EZYwblkz4zxHzii
kCWnF8RrZEr2QXMD+owy/M9fdVEBEHAW0ipcUlOvrOjmphKbOTMJ+p0Agubf
o7JXUua3uZFCIzRKlrtsATBBGzMHhUuftvkmaO8PlPub/netDmSDevcuIba3
EqdMHCtfALOt4JH/nWcuSX4sgfc221wkiRabKhCbpQsGZtxzHAOmWsz5KR/z
icqsX5wX4Cmd5BJpscPP/gYDdQkj8o33tyhJRV5ejtwqP881qxTmcZgQndxc
hKRluSlq7dJqxxPccSh2WAnjIA4f/pirkqq2DcFzIhX0MRllzuHRkaUE41ug
hWZcUtMLrmj+M4HDz0R0u0qLHmSK+BbYNhQLhsrSQc6RcxO6ckmnF81NE431
OAz0Zru3O5m6mqEl63AAThWunDsiEeGX0PLnrOBTleiBrrx0m+zShw/oBCz9
EHZKFrnw5HyzxUhR/JpyteVZobLhqRKKp7+0azFstt8WA3Pkb6AHZGeWDOfT
f8XFPTZqRvz8FNg0XiUUWLn9EOPB3y1ivZ5uweBmBHJd/Rt9gr/dDmDRVFc3
YuhJVGANQzQgqHybyNfVLdOFXmeHpiRzqvBos/msW5ZKsLdUoZKG1uCS/tvN
TLNYQSft3R8dMudfR6vhl1Etri1VyVvXweegP8tlSXfpoQ5wXVMbJYGpGVmi
dVXzQyQrpS49SsJJqFvPeKL0JUFAOuu9HHdygvoSzmc1a/zn36UDlASf15xa
Vo+ZC09cB52J6Zg8fwOAuIVAIVP84BE6rGgf1VeUen/LGrIohC9aff10XSj+
U8NYofJAdiV26Z/oZeSJs8gdHWT04WNsGm8sqsOVw7SbzNJrrSmEOKQJV/O8
IEnwyCQUylmRhXjIeWCnLbNtC61ZpCS75huI3xhtbJcnzEYN3Vl27AdpoPsx
C552yDvNbbAbohUV3PhJ+J4+kShTskebzdndJp1o6AkZm2PdrsqyKaThkeRr
g5E2bJTjF6VPORTWobz08ECC14y9ftfrulAlaqGcsi4VYoEsKg62h3UjI1+S
RiCjQP1wNwRYX0X+70ZIbxK6Sc/PEHWiixlRczOiltTcBndoZRwRKi15s8Yl
fv7o8XeQ+gDrDrFLw/geDuJDM2x2Fm3KM42PptvKoufqwZjAWJAmAtolEEEu
W3e9g3gwESh66G0qocLTIIMohKf6tL/5x67SIcq5D67RvaXrOnB/I2v56/bC
uwpaj0GZZeAq+/r95JW+dzlQ05yc9+3668QLok/fGMlg/OrW83fQkbzrPgZQ
Q9SaXlnw8eTjRmdC3ytfoytqX5ozwW6BgtOCJBIP/Z4tXD2YTpoNSCdqQYRv
ouW3g5uAqVTsouX8/WPKmc35iGLZZ4O6ePMjJyRnaLmW2LZLRzwjhWGxAa3K
zC0ulPtznSsXg5Hp7j7LDUjRo8Bo9ItvutcRBvuQKouHOA3BtYmH/wcaf14y
Ex3xa8oWoWS6kKNv4xB7p7vhl/JTPQETGEVxA+7z5kk5KglLtz6mD96EU7te
kgjZvvXZnR7N6oJBqXZEm2UZiat+BVoe3gXI03sDrJMRQSLb/rEPZlTJIVO8
EMV8FS2YzKuah0cTSlpu1CHtLHN/8NLKgsruLZ2VwiYbH0b4um4CO0j9DTCr
nQtG7yW7hRpjHi8W+pk9+G5SsxQmq0AA3pBF02Mlqb9vfBKiUf4rdiY9LpfH
2mQeEnT9RHEQHJJkX02DdCusUDM1Ixy4mU1G0pM55wINt50vwoTdAg4hks9N
ipcL7YuTYPdutnB4WPn3u/XNxy6DUmh2nfL7ufhUNA0k3JI6uElUOa5nqJVC
q+qMc8ejDqanfopIP4cplNPh3foRp09MCAziTSR2fTNBnQzi6NsyBf/TC2Q3
AV+DwvoFKKhWTe9Z/UporN2pNs62xngpgbAvhvhpFrS++LdtcRQZniXeyyGI
TFqL/I3+JZgeU+fog7K0jRq2xpmunMkfrYLsluzbhjdOa46QjCbv/Y5Gdhx8
DYFUqbFybSNBTNgR7ueuv5bnFncut1lOZrA5ELEjx1d8WHYWDSFStpgxJnYf
BC4zblBwkB3pvLcqb4WvQna8nnG4lsXYkzdYeSWUxc0bTMwlKvPT6FktwK54
pfK44Xu0KI5/ml55Iv73G0QnXJOvtL1ZEy2XRvkV5v/KSKEYUeaivyLNp0Kx
q0wXSepu7hl/bFa8Q0Id0tTgzVMvjvPYLw1pDTUjcpxC9osBcomd8PkLBHMJ
cn+HzAr9SLdI6xIZP233Y/TcegsvPPuHmV32Y32vuhQJQHpJVDM2WbrSq48s
VaDUVIJjKnv47rWynWURAxxESPZAS+/KWl+Edo5nFyar9EshBmOb2Z+aWbQU
TGKx61JqUT5Xux8Byw+tNF2bjvjKilGVL+GD3JsA2etWiQvGiX+YVLJiChTF
5MCRA8IGj/fwp3opbClR9F4ZWMtluh33RiRbMi+NNDVJDUFWNRJa1DcqoLb3
Aniy5g7CHyY5lKxcCt9UHTbyBU0OgHpz8G9VICEsCCbw8EKp9mFjAa8Mf08v
wWLIAAdJUjVhyHXNXyH9sk4ZrKAX2XvR+VJwf5akeNQGh++1RwOEQXm4U0vA
XumRCAUKVWIUCRCmlqjq7B7nrq4FPCs3XX0YRgKKdPiyD7halnw2ncfhkZ3z
YthxWTG3RSiEAnjn+hHef7XjCvS3DWZuAq46Ve02U3lyacxsmgnorFET4ykF
inObGhPH7ahwsAAnfWR2XhZx4I6peRyknDuqEL3dtcmRR4gazGaAPOq0QfHH
g+Ute0VTAaNfg2yXIg6ZWT01RBzlCVbEAz6h0hfPgB8ZPWsiTqFM6DyBpqx5
Wb6Q67lzbZIKWGpEDwsnmFJiYGJcfWNvULtOGmbtecHc1gABMsoETuAV3zlr
OJlK1quCUc7Mg0EJwYkRqSMpPAd5Bgp/n/etaPLW/S5tznUVgdB4XVG2sYoj
TMBlR5Zbv9dKuZQcwDekKZRX+J46/P3CM780971wrCLL+VtdUuhXKKn62/GB
A+KrTNfE6gz7UrXXDtBVMLF7SWR9rq8EZ491Hy66FDTq8OryqxWXiK7P1pX4
v4rlzybT+NAYqSnLTbBdpj7z9R4iK1VNP/t6JJNb3g58iCQGxDR000XsLoXL
ZoiTYhnrGZpiWcgMsSux/NtWsT1fN25M8Pih1H53TjFjDZFAD+IEAzg4OrLv
Gnp0mduw6udzXjhbn5dav6WJAkOl/hpCdf1Vd48B9vUtLyXpAtMlvo+fUR/S
Sdu7sYoimGwFKX6iLUogH8LKPWG8zXa8IQVBZojnc4g+et1Q9bp5a5gfczKF
1ioaJL7+qe3+JNmfbUZxkAqLw2xkGnBQ6MjqdW+0AEf+dAp7cjr9y+lQ21Qq
YKgxlzDPwBGW6JmAcfMdAbc0WRkcxU6k037XW1pYP5eYjSuLG43x1YgFUV3t
3zk3keGfg7/8fKbfeXMNsvthbp1jZN6oedAjfcHKKinU0eKGHdhEqt/iOqip
e9mHosJGikxDWDj9bbnSaODIMPuc9CQlxGZ7F3gzUXWRPdpMUs38T8kxMkzl
w8Qs/1/8/aVgCS9t3WPfVY3PS54xfLTVNEWw2sogsf8ylT6eB2JA4EW/JL2L
ki/kcpuJU97J1r7nUNjQcBPI9xiBtuJ+AHJutJj1xdbxw8n712cosoJS6DfK
0O6Wb43iyubUQXyfqT9lMCRfCkJj42NLr5Z6PoZG7RpV3w/uxr4PEyIp1jyC
QcIEr/wUwSnl7KjvshD3ZLn8nEVLInubtxnDAQd5zjtKTzOgohSP95NduWnc
KETjqSMvuEDLG6PKlkBvlDc1sSov24q8fPr5zbbx5LyuCQpuNRnAwkukAVQM
x83N+olysu1VpTfJNrAZE/qgUnI01yPPjZIcPSgUiTzR4WbS0WzpdSIrFF1E
T5zw0LgTjMDyPEVtUF+fZ0ZC2ki4/a7wxW1z0lV9i64MTG5c2o57bKi3m45G
4+eRx0sVceTvCNKb1fTdpJLLKqFFfLNszOqCkOEQfsnZr84SaVmfRZ0UzQnS
yvnVUEXXEHvt5RqnOjlW6qJWban63pjfSr4jpUGmd2fnJOLDTZGTfPdK+tl3
KvxfUzTl7M6IzcF5Fhfw0xOXkXy8PIwpAZ6a52mFwY5VUkuVIoaDhCHsYLsj
JuXWkpPbKKMDRUBmsdW6lkOdzkjym6hJz8t0CrvkGbhs8X3R6Iis2HommfBi
AWpYhoxXSpqBxvV5atHc7L1NPEaSgPT2ZCRAaTIDWIVMW8o91iSGlGo8thYg
NZVSOB4oMpYE87ortPOy4HncO6r2Pect+45s97N1kv4DEvy/Ds8Qyw7pp7R0
VOEmRXCjbBc3VBdqOlLYr02M7XnA7Mn5xRjpp//cijGxtIq6IL3gVOeROCtN
NxCDlOK26EL5MMcoP1e21KlgSwJwP4t49ZjNlRpe2unKSIWeJjk/H9pLmiTO
JsNt2NGCojGwdw5BxToKIg7z0XXb6BNW5AEYvQSItzZGP9M4dyEcbrmLpIpG
4d8IJgfvXTQg9DOIDl/AGtPT4Boq2biq6jfETCvL21/YNpzTEskupArhQkyP
S2iF5PfZO6ZWZtjQe+6CSgv/nB2bs4ljqNPSrEYsRYTpLUkp0qv79uWfh1Sd
GeThSZ460zGraywek66XyASbjBhg8EPEeZnsBqenQXtIXgBQtmKX4HMbyzbG
6ybsRchuWDnq1nVTzYqmpqCluVeEq/gRuQq+LrgGtBILlheejYHtnWL5QjHH
TJuLqol3gnAPiFLira5FdyTZ9nARXK8dGiv8yeW4ZdQPItKmmsZOsZN7nOEr
L/2C8Jv+OwWEHVubicz89f/AES7wyBmnaD9SkwWkwOd4PmWdruhZIi4Fkn1V
LcJd9Jntx1INr6ctCPVvqudt9UXGkCqocNUUj/y38PiulN0Tup7VbKtQFAyF
sBV8Ug0yF9i0phToGZ9V4I+zWk/gmuZNLvXwQ8mKDD1pQDl3K0eXzNIK+N2b
3xtO8hEAmEqHlNe8MBktEhP5KbRBqlqE03/ziXfeXwfPCRXAwRr2hpVKe+FB
MMOZrOWdkFKlMvJRQ634ejnQslCkmLwJlhqPyhDthbseORNxW3AbwW/9WhzZ
alzL8E+yzCwckxlMAfpo1YxmwcX2XmbP2zr06UFN4WU+fxKbYbecPbO1QmsS
5/avOmcBpYDteCeyxsnFV6I6RobntSqgSfTrNpQIFZZUdRpBV8OIooHVstvX
6KQWH4TCN3f0zYZ9rT2sMXD0ejYTAKdIx0G26jn/wgSRoa1L7Ilnt9c0QvAJ
tbj0UQ42pVjlXOrmwEeM67FcTRdLfsbLdGOO0aHD6oAZzqNXtoYhgzhuBA6w
aLqNWei00Ur1tb3LrYoX9jW74MPMG1rNfsXzCNI6kcc/CyMDvy5BctJzBJkM
d+ogNwWUUSKRNfYTd/+obGlKpJOBS2WQ2RT2hpg6mV08+BBsoy3eucnvc/00
J8MEgNAd3kDae/2yS39Q/B719c58LT1x7xguMckIjeP4vI9lvENJudqNOTDE
Yt786dSzAMV6Hk82f31bN0XTPKzahaAyY5y6HYblMTvlSb/c5ncggkc0EwW2
CrbG/aa5C7NK7x3HB8s1PCApZiRXcOCMsat0qFcb2BNXUBAVPKcU/squu8WP
mEZLMTSrO3aD57zJDKOEFc0FhjdmLgjfCBuCihX/wrJB/L0jGhidM084n1db
2+Opz/fG66kcIsoy0/P5/t0beNDgcBuBs3AO/MXwMmxVdc40moJ2lgv2/e1F
Co/X2TNwa368jmLSG1v5EU/bfOwaBwelFfvjwYDyrG1yxc3AaCtYydpeVM41
XLvn0yQ1niR8oxcIvdGRPMIaq2iROmFgb7OGrj8FIltRiFA+DDCGRu9vMYi1
nSiZXdc0ACGvElWkZqNEiEW7vQj2EveZdaFdhjNvvWzUb1J1THOLe1jRSIWN
FcFGHbn8vwPccR9ta0WmSqt6pxVnkQdoP/ZrtTwbDEIuDkCIbDjCBFhfw2TX
PhEuqn+kSP2S9bI3cPzVolTEXh0N0/lVJQJYKjlEik2m8T8TSRFXzP+Z/QFE
2eYErFjozMvzuo4WXBl9B0DxApPOJnBsaojSrjvTSSGmN94f0zwNI1aFWqfs
9nOXhZyvoL2y8P5u2eUoakNxLopLoQLxtmRt6cP+jKKlmfTUY0sOmDWNhvKc
iV8sTglmREFZ91SZ3CgDovhfrCDmrEHcw1sDFOvhbZAlV9bZVpVMmlIf4J7A
H8CoIG1jtsv1WFHaYvybf7wHT1sWbm6f77ZxIB4eMM5p2NF9Rf+T4OG6aC4X
cVSATyMeUjtUEEOduBUjwh2priELy8bnwu53KPb65bwxT3w3yGibYlAzFwfQ
bzWBxgjVbd3UkPUT0r3cE0iA58RLkkla09tW/OlZvH2F6ErQzmwqxTtg4gwD
/YYsuHqAtrA3nutii7etwE2+WYtSYFPeCaUCouXL1FMYOFgqiJz0Km54LV7Q
ZJ/ge0v3QyDDa2ByupOzUcrYDL/F/3QyQpP+wHezANbF/BR6APH5kOqhRfU1
9dEC9geUnNRSBzZvG2I+mPqIRC7+OnTHrLc5zYYEquVENMz8uSND4JtiX592
UZiIfr8imocEqRJ6D5jdsZF08uVLVvM1/b0ASZMZi/2ohdTG9suUVTZLvw0I
XPuSc1vhyyLCanujutxI6SYZXtPe5OEns87UPBE58jNmVpRX2b/l+Jx7+7r7
X9jvKDsTJ1+hffariUeKWlkP5hA9a/CW1PSX7kQ90O6FfKQ1458vu2K2Bt1/
ueP+A4ZtEJeu/sL2+eTi67DvWydXIwZBtT+TCcTZZV2UnpMk7roAC3R9u8El
qwOyxpgELevdFdCGRROuqMwBVwtP11rK9QsT1diCp0X8sBMQ0oQC6mhVIkaK
mizCAGDUb8GzxW2+iOjGUN4tNN8xkmKlCINUb45LKNEgT5WgvvmJBqk8Clmt
wH0aRFkzsBFQXpjrxvb+YGq42JNX4UBf3QyByJJ1v8pvx77mzJVjvYzwoUw1
hzdCyiFu88FO5AmIR1MFG4cUNL4CZrmRbZTxbavBXTfmlbWeQk0wZf1Mq7kd
y3VBR5K2Qa74BhL2vaqk2dje6ITJIEt4C7N1WYuuBuLsGPRfwDi9FnOZMV/8
SYxvzHtg8KZEAWrxRAvpn/+sjyKvAYmQ6OLpXbxmjmTXwcvvVSQ5Rkhc6uCe
WDac400zwfUzx3LnNnVBhMgWsgsGOvaQrxoevaMNBRF+TCnTbH89rb0IQBHI
TGOIXXPjHWzoqIRLoV6lcwoasqjHZ8AQ1SHG7irLY62mkkfZVKhlBkG1L18G
902zfpcg/7HZogt4VIwd9InBrcdCecC2eHuPRpQ2iC/YbwQKfxH8PQWqkxIE
MYIVPiZieKmxDIIN9VkQePZK5gcGpXELh6NbsQw0peTKuz6yWerl+kHaDyh4
c1cTi/1AfjW+cLPlCEmk0hCTgh4G6c9HVC655JZmhlWTywOdZeGAqsH5G52l
yU9/BM/edIEIuq6cxqklkrZwbZ/a3pDEgCAz3iAg6QtrNlXy1kzvoZHk0T0L
f3/mS1qa+M3l5lnAhxHRqGeKwvl14wzHEQL1oyGn5qIey97iKovinLaKCCVZ
AWmd8q35ssO3sJ3eIZ/uEbGa90Jj1HRNaX9HvvOBjnZYgZVb3JLjOTNxfceY
lPxCyEV9bMpSIss2uHPbS8ireKidF9sWqfG3Gg+QrY81YVcGDuQXxO1DHKtt
W0MuvH6kayCEp+UuprrCMXl46ZzuQeVbXlB8m1gu90ipZs/o3HdBmzSpIPSE
CZkONjEsKMeKktlCojs9ZJ+ip4Sd/0S45WWFk5HbrbehuXEVgn2KXMYVLzhn
a0KaguYKnF1ZSQxOMOs6j/LpZFk8Xda7NEfKi6guDPhL5QHOxMRTZDTzy4Dl
sJz25ATGv9MFt8zzyBy+5LGW1kwaQSjTYLMFwSR8YrXJj3oMPx54WlRZSgts
GycWQPh/XH5qN6KB9FEb/Y0On5YYcIRIjP2dDD+CNvhtyOk49KkrIgirU3iE
snkfniVSvm33s2j5ntKfgm7mZRR8/oZesYzrI2DtP6ELOPvIH+ZrdhI4ydk5
VNnG4kZGWkK0ZyMBovmuvVbhdf6iDnAo6jSz+4utly9drLCXXNYGtLaGwrFn
5VEYt4LlAE6tbs1o0VUZVCtL6HePz6/9t8Ks1vyJNVIsvhWsBQkZ51wDfYR/
8NdRhi5/iyu8D6SLlVEmpnXeoOgN6EEhoqAePYOAqFd4qFB/vHwlyvJxmiHw
XuwU+WImJVPFkKjPKTWvC6KgPT8byz6MxkLp3QSkaPG3IBzb/JtDnTVr8V0+
eDLuG8e7oXhgsaxVdS4cPG5i4DnFLInjhv+lAcCjuf3aoAfEYTMUf3Sqv2ky
mscTz88NqvRFoidSYX3YlbRBxpLg+Iw80+XNo40ZxtiG6rJimTnzCqj6eNfC
tWbq+3Sbl5gl9XzBxH4SQ1FbNHLpkSYln8LmBWdvzRXpmCztbqkm55kmq6z1
eoVb7kHJiTLnic6z9Ml6pgCiJvUNJbNPJnXBbcSji/i06qg4fBXDysy/gRoY
TBwfyUUZp4JXzz/9cVSRxRy/gf8LgUrNdJb/HpfXHuZjKmFX0AIeposxkZVI
YdmOocO6KtlSgMYljL+7OhTl2ooinOB8Cvo8PgMB88Irwahtfli47WXVDV1R
JZiSyuYhjA9TmPkCdLlpXqOoUNGRSg+C+rf8p81qxIj5Znihte9SPzc128lp
0Js9fUR7lk9XGqugPvt/BDzsQbkWwRNMjIICCtKXSK2Y51q0Rdbgt4pS7khI
Sg3dPv+zXQkax93eV5mng3Wf1BMzrX54Wvu7/rq6e2659qoPx4LDrRcRQods
Mo09O2mHjG7GhAIOls0pg4eaHUWnkWqn2Dl3HiGtP5g/FirLi6VCdnKXR112
Qbb3ONRqA7SqmM/mYI8BaRLoMjbC/e9OG9QpBAV6khg2x5zNm3406A3ZjvsB
3GxKL0pqFadwwyDQbaMvaTYdVuEIwGuZPxkMC8zlrUsg2Qytv28eR24WIXdq
cEIihW94MlZ/DCWoZSIVn7/eKvMDnPKgbkUTPsyCiqjV95//nZk5hK2KsIhm
PLOvtnDjf89R3sTKsf4F05dmQCuSbMiEG9ixaZ/oVEsBvrCkD7NRthnZ2SrA
dqlowIw/M6izOk5CKQTa0oF2QQL51kOc7hg+r5WMBaOlD+sEIpRN/O1pYUiJ
el0Nc1xXnrTrd3VV7j5HT8HqbxTNEwUQrdP2L/e76cqU+y3Bcm/a+z2ky58m
nOsa9O7KsoUx+W5T+6PszavuZHh3pMht/GqcZVjAn37wlD85TaCuFsyrxGMc
QLBxELMmpH66NPftoEJA8kvFLorR/m2dCAfoy8dRDKbA8I1QehT0mwLz/4od
6m4Z8fdFY0F9OoI/LoGjbDrhDRjqruN6pTaihXCtPSW7eHc+Q1FWGNfqcjfP
tHDvav4rMcb3z+7ztpVAnacQCVuGUlgBv7+4XNoFh7a33bdzE3VyWo876mdD
+E6re6aBo1z+wn7DNsp98M6EebU5R2P9zPB6ECkiVPGl5luqEG/kDcClfmfh
zC0GddOj1Qg6F03u6GkLQVFCOjAdlxe2oypnT6Yt307xmo0mGq9OZmomYvdT
1eb262zvTqHpMcysB13ZEgeTn2Wrnf+D6loTOJkvUesWv9msHCjJ+Mrsj+4g
25hmYVKs14+WL9ISaHL6PPsl4wBzRMrphN2fbsX7PxrA9hCAAOQdlIVTb9Sj
VwmhdNS99m7EpBO1gZaU++NWVQytfQviBlH1Gy3RqvbwpE6iFDdXeVvjw5VP
msQSB6t0fyvPSVLwzTwb1PCKuHnJwpy/br+xkYNm0HpLi17/TxYx7xuyNvFg
lvNMeiIKW/uCyIsLjAUg3vh128roShYX7TSb2eO8rbz6ny5aQn2mH3Ekz2ie
IyqE7P2t00pQxdskjLBuPfTRlM/XmvvIsjwmmBigKbnkBp3cHmDSKxlnqEqq
y2yFdByynRiy4HAr19nZHGwnT71bvLdHsIOSF2Xn79fS1hgH4nHvPCi8MVdf
L4Hka62cAKcEQC6jIU7jBE+Ww2Nixut1XRx9rieBbeWviXy7jiGuOMN/tRc0
0bNMKQWcFXUEa1QUHSAzcbry2csTcYMzWhK9+L1mgRtALMpDeViJ6N66SYMr
0HeT0W6gEkAgFzfEzzTzr5HYrcxpFPKMAJzLhQOLlD6tPVAmu+A4AJ2eVQY3
o+ZI1QH6NCtlHeG4Os1Sb4AGrBVJI4uBe8oyqNXdOtWY72tDZ/3557pKWPQ0
n4qYS1CAIhksGRmtyRDyrfKvdtuPv0mqhBYq72a9gaN2jWDh0dZRoZZzMDL3
KXKmPUKzVYt2GyGaV+17u+tDdnaQLk1RM2lwSSFE7bNO7w9aTUtjOb0S3JXc
KkYyhgLqdR5cQMz7+aTpHAibEnun5mHM/slLbzswD87DxtYguu84Wv5EWY6M
Cz3dXEEmpMq681fimjYfgd33y4YTDMVN8HHp4VYP4osbplgo+1YTEwIuejOR
xhUc0WmtdfTe59VclrkyFxhD+ynOi6xNN9/8i4vnD8C/qSgfm9E0Dsf84pzA
2kUwKfVmjV+4AAT0E0yIsiasiVER9b7w1GJVeZWArMPYuWF+mDzcPrAXY2fP
XTW0v08FJ8K21YqvseRKuUBOg6ef78fm0AtQGCuVZ5DQp/HRsNbjM55d+S83
2e7zt9Yjdfjq0gkwVd8r6x4ZDYL2JGjmxcXE0AekKwet//YN1dNKl9EpbSv2
pVB2aM10D99ybIToQ7NZqFOchQyF4rPUbZW64S6dpL7FHcNpkH2aE4+ds3Fe
IsfrxMlfbovFdX9SnHoynhuQrGXVSffs/VddkAdq056jOK7CZmPZwx/HNtF6
An8NujvxsrC2GbL9PB0wPJKKrHnqeBJu0YZvGRTJoCrBIHJNdr5MYUweA60L
H9FxnXlqV3q/lMNoUlHUpOAvxr5VQTdGlBeGIwQlhUgbDUh0MqPKiRJ0Kpis
n3MRPoxvtF4mCwGbwEebbldmsAsYvlAjp/boINiUuuCaq96Y098Y8ZJtUXpC
qr8dBnJreFKmttN0B2YAAILQLhba0aHZvQBMi6z7dsZu3+Vo/hVLK7/mPWiy
8QsyBLb3oTdrQ7zGNXJGQHALxaSkd7xR7g1P/dvBxRqAnQUCZvaHehWcl1xh
91aw7fYT0ahv6y03J1+zWw8xRu3DpDLfM4YMuxr5cdURlc53xLrDW6c1agzv
DmCRIJ7kgYVHV3LhVJphcYYebJra74RwZ+wa0AcZJkVPusotmcz/ziXkxuwy
RGo7WYHKVTI24Tl/SILu31Poc0FudK2sQAqhUuCMhyn2iBdFgwV8AHGYoe+q
oHJZUh7kNRyi6xosbZ3o1DE6Z4bSCIXE2zC5AjhN9dfIvYxgy4ydHjkTqjbp
0RMlqj8ky1aDbfMROicaRSlImGfE/M2niVMpBInUbVYLJFehNRxRLmJ5KKkz
pouyryshtMFfEo4fEKQ1TrHmrsYF/qNP3PmGcTBentHYiXunZt8549lF+meU
6Ej3CTvgXmaRtPEyOaT3Zw4zX32MsyG2udLXmCn/5mZ4IrKjz8UVTE58jLcV
NhHx+tCRUZzrzyqiSKzhg/+NiYr6XGewdenQTStaxduOvXAyEd9ajpobXqwA
Jd5pBwmNumIMveSUUJZPLVUi0TB/NAq7u2afsTYElNFe3NpSTOWa7Viv4x0y
5Af2lVv4mecw0SqnVLvip5gQiodlemAUiJ1BBLMBJP/s3u5vOT9lIOGY2yX2
+AWsZ9kkY90dYA/gEun2bBly+zisVL9ld03M8xQ/ugY/hk2jUU+9k8YSSRtO
w4b7P+VIJr4DMsTaePROTnBdBYFoYy00ZESVy8tXJ2k/3us9uysJlARUWFw5
IuuYchhbo/71KPYnNYeGbZ9HDuGL0XIl3sLZl5JRsbmq2RGeEzf6ML85lwpf
P/3ko6FQvpm7ebYKPYKm8lK3FGnBUutp6R1ap82iaMe0bcdJxgrp2QnM4OrT
hN7ZecZSMZ1nW6l6mVwAlWsri3bqnb1FjAZDfI9uO9PmLURnNOvHPngsQw6q
mRiqpR8zzMAxNdZJIeupG0P+ivNYoT0T9rk0ASvdYlAzw7REeI1vPIB6GAco
YsuyemfsCKeki9iCkSjDqPrgjTK+q8Qjtnjlp9h9nnliUFe68/hsaFkFxXQJ
v+/XjXTbVHAuXiN6FzUm4sDxUYigN9vNmgutq6jw6xVlIjIcx0AUPE3dCXsz
362SxBXNLh4ZCF7ueP7BZiKqjkihJHzuDeIDUGhVaNFT2kOW3uU0BG9sNPBw
E90loSL5FuXFAxy7qz5GXoJnKrrNT7GF6Ps9/3gb7z/JC1bCTmZnrJ+1b0Qn
/N1AR95LWkv7VehNfU0mgJDDj63rVOw0FNoIn8xJPNg+zgvAtduaTC25nFjP
jECByosp9GdDpxgc+JYBK7i9WCZpuh/U//q9/NIOmmzRaFvXVbxgHfAOe4UP
8Uq0Gz5E4W0L+TQyj3t94m/lmug28+XLr+yM0uQCEZK4fZETkmidsOJTeNdE
uQ29ugf8kguDEvBrdwuYLmkAfIn4oMZY7BR6eak5ZJSodcBPBg7DAqi6MWv9
pLmQ2BEhxqEigne09PhZVJVqkWBHE781quHr+gQnC6bFsIwuZm8COFeBTAFn
x80kDkZSh8O0lOG/MONnixMtTKKUQcqIfnFN0ZuZleNhwlBv3AkRsDPGCise
JKo9/jwoGUV+P6+L1ROUJi89O5YLfIUM9q/TmLV3Y3UfMDHI41VSuNwXX5P9
d5NawP3PSJ78V32XeVFupfJNkUK7VJMXxEWTqo32JM6NZk6UdNKR2aA94P2l
OhChJKbpW1OKz+t508w/Qx1kvElHFCUz2/pqLdHYsFSDUciWFArda9DT4dD2
zC55KlXHGTpXQ6qVJ1UD0v14/5yZUAjNao1cnqRcZ+qbqquNjBoZcPPIkAMw
6LeK2n5FsxjQ7tDqJbrYJRI9NLcz02SK7NxQHl8atuLCohahqAi4FZ4encJY
QrG0cUNr2M5nGLYbA2/GxmMQQuRXMTBC/Ayht63Ywa6792enB69bNozrgAt2
puh2gpKzl1PMP/3oH/5DqihxvDw1IguiIATuOs1Z0Ut2y+fpcl71EyQ7DWhR
DoDjfMVK+e6Tzx9CTs7J5596rHT8wfaqzjydhvSHr9AJlksQcQt+XgSp7SMe
cDrgFaFMQMjqCeO7gpvQmuYjQ4/3HjSZLoxqRP5R5cZQJMQe1LpPugwuI+Uz
yyQ03qQovTDTs4hDIYztZZqbhV+UeQ8V1UIxptOqsNLkSLNfDmVaWHgigeSM
KKQI/s23qKvG4Ui0iTsFYGOiECrL9UsEAxwlnDfgwcDH23ZcyUE+30+xf3Lk
u2+b4N8tTc/mCJEbFWo0vBOxzuvL8JbYVdW8NyS67doSB1wFYT6JgZMTWaVn
geYHMIhHHeFfp+QCUxtlPNN80BtMDvVYAC01UdAvwWS549FL66ZgRfqJRS8w
oAHarmjDP6IF+YSU0TpHMEorNdZrVQ8L7tiMYWdstqwrdHVI9rjRQxz4sIPK
KHkrdcTzR4EtaLfS/n3Dze9tladu39oN4bDlDQ7bDYW7QKa48mIhKL+BIkcX
xURvoSZr6NvACUIZFDwmHuwBSLOx5L2bl8N5/uL6JSQnjAbKTM8XJG6DIFb9
MAT3ADCChoCx4ApN/lnwgZMM1NsvazcDGMQxOmcKuZ4fjm/xaR3FPi779u9d
TSphsCE9FsabejZsItyITN1SOxE77eGgJBIsmSornEjPrquLPKfg87Gm1qs4
VTB1z8e2jD18agg1IGq/HG9nuMxagHGGPwxlqftZVJJ3J3wBCGhZKMqKZJA1
mmhYTXeZipIRYJp0JGLJkNzOMdy8+aNkiwqvvR5W1PxB4WnqA+EYSxZa9+vN
eg5LC6y2GB+qB7o046emMjufvYT3M+ivJxXoquWYGXcMPvnH1XnjX3C421TK
MuSUvlU/yhUgQ+WAf/zmgSd3xeLrXfg/FpyX25sMCJ9XQU2jMAUPG6dFInma
ToShSomFqZ6DojQli9CcImlU6nxGEg9z6aMnTd3jQTwjL5+jnilbnYcqXTfF
P6pVytou9fcOLccvnjtOh0500Wnh3QFXWL72uFcDStlrF/PwBZrtJK+3AW2g
IBYIA5phKjK7RhCT5b0Zwh60l0hY75kbUFkKr2dfm27q1ngmPvQfNXTRD1Z1
sotyHdUeulyZNyyIHVFKmDDyztAsot3W1Zh4udf/ReIuq+Hp5IizjLlYTypA
pwc1u/eOobPcZHPywY12oydn1mEPGeZAWFoyCBPVtH4ncYqb1x461QiKxsi8
eogiwqCC+Nlle1MFHkgJ4sgqigRMWcgibwPlfx/XBfZvNi3tifVU+lJoVe1L
B2I89SL/NJGEmFgAgvRbfKgQuB5Ujm+EJpFfP1GXRYJpkbrEaIdzDolO+3u6
UtWCF30v1KXdd6U0BegyrCkNg0MaKQBDwbotkETsDkGNhfiEt0vyQg/poXxj
RRjP1OJN/9+lctBxR0ElFkMTvfZk+oM60vKi0/VlGsS6/GE9kbZrEomkpZOk
43Z+2SOtB8oytPb+m7PDEyj8tt+XZI1c4k7ipngimNWE/pPxbYUa+I+cPTfi
98bGiwd7XH5It4rn/7lwpkFDBR+35zcLpn3O+0oYVoerWGy1ETUY06TEl9U5
bcqxO2JCiSvm6/YIed49cIvsG0BTvfRhGp+L7zRmGA6jRdAxbGiyKFWcdYew
CKBzcOITw6yXU0vymzbdDog+81u+kuZhq+N00oYoh+tAnck5yC3jc4PTU4pO
jl/XhTN+LcrDpB2f1POKH2w6py+5cvY8wxxyhtPe4I6nlj9epjFDx33S3qRs
z/yslBVziX3Ny88+Pe4T21A/IrUyhZb0sQ4q3b3/6zrdnEZKNA2YuMiINQza
pg+8Uw9b7J/YVa24DkUOdU03IDuaccawSnbgVrNi6PFpzwRlJjizf0tOr74z
4jspVHWnC3bDP8GLz1RAnBc8ZPYFG4X167rARrYuTMF3cK5R1Vzf/P+W9kZW
IBrgPr5jUlayRuynLDBKYaczAsuMawKP6FkYeXllNTo9TIFa742No6kWyOUy
Wh27FRTmct0Hu6LVUqJ6QeX5i96TuQngYJRW2c73n0+6gpKVOD0d8uooj+tH
y3jxtRXvaEZNjBrKok6+vFv4f04N0B9fggjdRllmv6uDPL8TsNSMQpelcua+
pzwQ62jcutN7DHNyETWDBiAMr/6LZ/2UlJ0QNim+SpR03TNxIvcgiy6Z+/mo
VH0Z2Y9v9o5lwHRoz0W1avVXY6g3/ZX7Zk+J7DR6TKRTjKRxktWg0pwd0G3e
4cFOQxKSxlOs/sAMrBrlFVaWT7THOAwmlBZALWUmHVnQB0f6wrmyCBFTfGeX
IgiUAI2X+FbTghEi8VVBN0tAcneHiooMnFQmhsmNr0RVbz1MSshNWyKFR/6l
sh1ll2X5FLmxURl+yokop5Awo0Fsq4bCDUs4MG2M7HvGJPd3t4uYjj5SZH06
uI9q4+zNdCD75WLtDP77uwTGOiEBVd3tuWgPNq4zi4xj1pgzSvYrVmvKWmXo
Gg+Rr/kQbLuei9AVkjdE33REceSag1171QjJNTbK+hqQn1s/TakTTB+Z+wMU
L1M/ckAdWeOGGlbelxNSuINL9RRZ3KU8qI8c36/lK6hiZmVmt42sR7OwQ5SD
7wGn0PnOVBbXX4XMAvdY5yTrurWCulTUEEtKJpGLqgGkjZsZlp2GeoIWQv4q
u7aZyrYVqHaMOAq3CR/RvwOvDCu+zecXg4fL4i5D8U9IZt0DoCDBeT3dxjh2
ZL6PMnaB3L+sIv9J7XgA96iJrByeSX/Aqqf95R5WbrLVT2cpgHM2REpWFlvF
UwXUTcKQ1MA+jotU4rzIXTgFwdpMj6JguSalKjFagfd/Ik8os97kHGDRTGWL
gbyJzVYJ/Cn0qJUFJ5cB5D4kaeP+6r6rPXuYUlprMuIwDbpnlNVv02yo6i4D
9jbbXrKfAyWOTuTeyRKD1tcKAsI/1LvBGKQQZEnIxqp2X6D6F3w49Tp2t+P/
fHr61LjC/4nFNJxj/m3VHJ02xpxjl+5dF0M6L973NAvX0EYg6iVKX7/RpfQX
J2qIw0k8r5D8e0roYM6z7Ro1yxUz5hsEyDZiGwaM/xHqHHOMwI1rPJ/m6o2W
xCzWRsYn3ewvn8DSrP3nwBxFs1pyB5FaAthsW0fMlxzFPNP9Z2klBjW5SaB5
dglmw+rVo2lpaLsG3lvNk3JHKAafMAkXKUC1Ep4417Oz4alsh3fMsvIFYUVd
vOpB/yxJ2i1xWNTcXxYrBZaQUBVbA4myf3uUkCS5n0vwjPhHhkUgGs7CDUqK
BfvAhvIAuvmlHB7wLnf89ohJSWKiSWirrlYDdAFGsrA6Cak8HRh1j8f9jZpR
QiyccMsdx+Rsr5rJhcdwrFeq+SD0And6Teo7ms9SvFqGVFnlSoWUhE6+gEaF
ZrmhcQ9iyG9hNc6zbygpU34qEjQt1vpC81WnYZQTKljuDIRGFHSpnn6+hFQT
EaeY6BV0HtPPzAlHruovf3Hl0IPiGG3ycMjDtuEUqUHuC5tl0YXeyG7oQ4BG
z4oCVJZYe+1eNqE/K4jRf4upqC67GSdg0DLvZRrvpLqj706ew83mnj6THJr7
ohG1xZBhm5RnouPqBOpB3LdmjfXJ9d5Lr2oo44nJy5bXjbuzcgw128NlcM44
stY3s8cwHcD6tnT8zwz1DNsMwPv/5tZOTvk+HbinGjtm6sH2YUmKVwTttWoK
deEttHaVfsILGiMA+9xXQle9uH4/mcv8u45xHvOFnmY11VCSzuecmwpp/UgB
1S2FBVIUIdNZl1xzasEi3vYnvm93BQvBpRMxhHB+kvI/aD+XjlpelLcPOpR1
usdlRTAzg6+7/+taTo3XlJOA1gm76ijQRJOxQ7uYVA3X9Yya7i4clkVPUJ8N
CPsyAa2xlyse7ukKhldwNpvZEDTAmPTfI80qRwPIh0n3d9+whCFgfsiQb5cz
sTO3R+2Ez9IWYFLCanFWG7d0EhcRfvhs3xnvfex0dx6gDpG7zufbAcQnhK2G
zWN9a3yY6mRXha39CzMMynO7xL8LsUxC+l4D4QHKrAC6DX/n51hW3tgHHDyo
UMW/0ZNQiS3KGK3SnOf3GFqmikfEIwlDAWcuiCpEP+vweE8sRxuabLF0QyNL
75e2+y3METTT02yFr6vNFsmaFDt2sM8DAAe04CPB3/ECXGnWVkH6u/uOhkf7
ZJL0HqPljCtHh1gkgHACOYHy8f1W+P/TohGnmHkb5mMuG98a69QGRA7Y8RZW
MuMCHqL49PEicJ5yRm7wEZuQtQtanGCLhF3rMikMB4XiyReHGEc4rqCJ5sEr
yY3MdxjcK89aH2TfovS2/PEo38SzUrYf+CJfwHh295JvzBvVOU6iTmmRYE6e
fK19TwCXMu+eqaHavhsnvkNP33Q79JbtnydeLyA9u8863LAsk4lQ0ujjbb8k
FzNlBYxcN5MQi0Rw7olh8Dt11I1odBy09qPMVrzGV+58KMsx7b3qIVvqfXVo
4oOCjFS/1cKnXFXgGy8p+WSysJopaxOuL37tHQXJzxhSrRKtryWTtvpjA8C7
T14cVnZ0piwJZPqQLuCvlJTobfRd0OlPrr3MyxEqT5j04kvrxAldrppS+iAD
6B4iPbC6N8CgF9RKq6gkztIBcvML28JyaP3CFIUucRJ/rgBHP/p9ZvzTWYoQ
7P+JQkj7S2g8shCAcBuO3FuS9cTg+mklJ83Fz5shnf2tXJ0VqF3ulDfYi66i
bCyoevgjerUEDNQ5sN2EfFIdtlCG+fSDA3tD+n/hY+4svjIkspOK7omlG/64
j/yJ9TPJvye5Sy3tHpkI93AT1jC6rKEtczYxLw4hel25AJ8vY6+V71jpskWB
EzG7wM2bkElcs6xieaXhvM61zyTi2AE8Ega3WUpmBVp9opUYjlXcJBGFO4f8
y6VILyUTBeCeXlNFwrW1nVhYuKZZyzkW5UHTxgIeWaA3xck5vbFENNzPJxqD
NYue6Rp/UrKuH9b45n8FwrYFw8DQNj3gkF5ILl6bsQ7aZQaWS7NA3UgcrO+I
tlIsmxBOXNOg7VA7FPOwTzdWQs/xNrGEbTt2A90W17P/r4VvkP63aI5jG0Tt
oa45In1jKwJ60WzChCIJK+1sjmFlcZml5NE5rBxEc03q6HDLlrDtBAbjm3Po
SosmKz84/UmL5TlXjYAECDhJkC6qc3LLJmlZYiiKhUOna/2vWV2n5Ns9cHRS
45+kQmsCxoI4Ch0dVsAUVAiRKa8GDvwHyfPE55URS7/1B/A/DkIH7oJtPQJp
4D/iu6CgUqYWbdkXwe+cg/jjT/y2rkVRppMuy4jyegjIl1NoVJS3ru8PXlz9
yRjO3a6ZRj4q5dNloupzZf1yGGFLoyv+Ti/EPiNBQHIw4WMDmVbx+KJBsPCH
3DaVK2kjQivO9I8XpRR7SYwO5BnN8mWE8YTb+xoPLrVFvQOnsIi81dRF7OLA
0tlsAzezjSRkdf+qlDn9VPFAS5wV+eIGQkcOl3U1zGMmp/YKIWvAxVNqB1Zh
FJFGOO9Ll81plCet/40YwfzbsfipIBx9E8WyOt4arPCeQfakkCRWjGRqV3RD
IQOI/3fISVNlhpipwdlrpBAPxAQ3i8vQ02Xf9nMQdB1el5WleDY8asyOWp9G
iuvns8feiYbBCrtTpt4/kknuvvdL5eT24gZWd76It3zfm/Z7FoE8OAlLNU5k
s8EnLqlT1b7tQUQJoQdGvzLA8pKTJI8ZS5/gcvhxcVuLeoEu0JDs06XZVOFG
SU/KLJnY+YpXPCM6dRsUL9WepuyyNm0/dmZUfFItVS71xFN94MLbhKVnhqcv
G3fvee16K4u/tJ40y/NFEopFcpgvDxayUmdM30hCTFulkqcadnR9ZiyPYe+b
Eb1gbzuNjQDQQ94i4pqZQw57DOX4iS5jn8m1Dz+e8fJjSQOjI1nHt9kxL9P+
stf0j+HX6nRVE0s8IPuKo7xTi5VH9tf0K2j1q8ryLxPnI3tXkO9x3zloumRd
eJwt63pnUszTWsguGp+oUpOq/1XZmlpbUixrjQNhmZYBxD5E+6wN0IPEh3Q1
paXWLDMbayROK/KLiWVtlI0zxGj6gFvro5JtlEj6siQMw/cnNCFl01+IIEkf
cz7DihVMwOb0ZxsFk5VzLR3JFgkOSahKnP5QgZLEjlqllpTEUJo0burhtvRz
lbs0Ay0bCL+UNeP+lRtp6czRE/gKUd/JUU6hN3H7u3XKAMvSYN76fg2Q1bIV
SmuMXsvIEAoOYpxP0DgVqvdXhhk+KEO2HENz0fbRLrtbF0pn3TI2vTznkfqh
Gu4MZjo++shMLKDWH2DPihRVHOlOKYlsq3Hmr3qT4t/VVf/ykBrmYsDhsD1n
U80QH9qR7H/zkAh1cetx3TRRTDlK4dXPNY2H8egejMvFtXAAPcnLx2K+/cfr
/XG6xT7g11KYKsHPVPcUHrmWhWv8H7NQjL5jE5sZfqWx+Mw8EGvvqbEQPKN8
mYWuHn+jIb1igd26qlcwMYFxOsP12ZKYc+Or8VZ9w8RAeB8fIbQqfAjlO/jO
ohyUUW2gLoJ1Cgw/mjcIg/zo4/TRxX562O0gfT9wdR4NYZ+vrOtC3UBq8Z06
9TNmKJgVS3KunA0KumJHvFRX0kLjP5feJySQ0JyT2H0P3M100PWN0/SynCKF
DWMn3aV4esWLlHpk4/TWeAcgnCE3iVbbNpqu9u/poysE6ctra6wY6Y1HT1yD
beXBAEhox5M/OFEhME5bntcZKA9+t8Y1DnSEbd/7ejMY5ocf8HexTt+7ydub
lrzxyEl0spHYD25+duEam23NxEjUDVVDEKTQWSg0QKFtqsNNbAsDu1U+DZzX
UfXzS60TbfdsUaEyhTfAM9GUKf35FQdH1p639SS1IrATC/dYJSsnvda4PffI
c80w4gHlPklXwlt+XR6fOmq+8r+dO31surEU+0SaUIH1ceCMr2zOAorJhM8b
oW+ytdazY6W77L+4pKo/tlK7jaB9ebZVclld1+fSQEMVprdiNQvDA+CW5Pav
L1ym4SQDue67xyWBOR+nnRZ+0MJh/nijDVXOsUVH008gmm/I1bAlDGM3nkPX
7cp2MC7G9mLjZqmMPlxv+fRBEXj5aLbmn0PYMHFyNW7i1MVLy/Ps3IH/ElpC
hBoHIZpIlcNgSy+ZvZqzpR5gyA6IM5ZoH4RhG9EWj3jkdl0F2figEfuVboR5
QNwJWhOZA8h/OLKE74/XjQ8E5qanIbsA1zcA1O7WlYmLrImVSCOuu607R9Pt
yThpWWOxjXJx7yvTkzCJcfJELQo0Ri2loqiMUnJoW2kFW+bhptZE7pAEnY27
5cqaoGQE7p+OxJ8cyjJ0IGX4uCqG+zwz2yo6BmED5udP+Xs6RZ3Vd9Xv0iTk
BxLFpptiNNX5omSXXKsIBuXYULPKxdQ1QKwTeaKQUjOO0hHMFgZ2SbbVdrtg
JQDJtKJT7U7tNz7VblMkOj80ayM5gCE8Kym3KhPQ8wmjlf+IwPB7/hcv+NQ4
HKsigtkVDWW3ZxBfjJM12I0h6pBqAKzvxzxX80KEsfNIu1gIQcuIGinDknbc
1/At8PI2l9cMHIqzqBL83q/onA/VzI5vcwlM3ziDR4agBPvn6pqOJArWh8+T
YoQ7VWiQ7Qn6XIIm5nddBBmmsNNYcPspws225jw264+eVLBZu49eMl+YdfEb
hq4u+YrjtJs2DS9iKJgRu1F9KDJ9d6rgW/NIulm/I8AxS4hhcqUsHthcUZid
/bY5Drgzmvo75Y+WovrZchGHjPGfHd/kK6970m3GgfC9R3mJBnN0aaHoa7R7
bmuQst5w8sD7ZFr5L1gt2J4UHfqg9RCdIPZ9lkbmDotBq2vOAsiR5EKdUgvG
3RMIxwgOSjOgxzjqbwiWlXjWAJAvxGwUSMTN0Shfzkl5hbHxGwlGHAL52deg
zR8tWjStEaiRsuopYR88zuLBQAtLkqqBZIcYNpxbbX9p2+DKwcidGL86PXVI
IEfTb9KxtbuSQpI3KQMW8qnf0FLQtgpKexYhOC5sdFN9AnrHdm9haeS+Ey2t
GeyqI1gZThCCdVa01z0NNo1Nq6Oitg/4dXYIbkihuymPcEnwYh6A53K1zukq
CAimxEP+HKIcAT4bIuDJuCRiKmk4nJk413Q+ssWK5tb54zez3diixQIhVnYE
NAUxHwr6bWI18eM1XCooGsYJ8YVcIjBhWGBwxM41yUwpY7J1tfUwdVCPGwEI
YKH36m3OOvxOPwYShXh4W5PXHB5Vyn/hvM1JbHolIf874BLOjXp78a/TSsWF
43Hk5Sw1DQ3zPsu3u8HleFY1R/W+/kdReQw0RhBGi6HB/AZEj8LRWV5pHbIv
mmcUwM4q+C5yJ8VgOZeD7BcTuH0tG6ROcg/DipiY7KNvxYWsdKyhsvFUnGrw
MN1/KBGPkyn/I1NmbORsQZWhXXeNIXvDP/Rc4UloW6RiMthWfWzNLgtRicaO
1azGDzJR09xM/OfkYo9UF9MhdB4q45yZKLL/0KCQQ5yoY5W8Jgml7hwKwxoX
OLfPxSc1KJdGdVHKf8/jaOOE2+t7i9rIxC7fe9j6vrX1YzFFOxlGj37T/SZH
VbfanizOAEd/0ZiDqgVfNSw478F8Y951J/4heklATtAMQLUW4HTzOL8eYXnU
6dYQOWleTQI0Ps24cBHa0f/l6YIEPfkbRxS66rBG9XKat9x9/96DDWtgGOWl
D+QDZD6sOwwn7Vx9AG3Pd6kIqzAqg6RQri4MBmyTtbwrBkbLfLO/trEonj0B
cAHvP7ir5AISC3MRAMsfl0giPEcJ2mwtS5lmMZqEnJJOs7UZxGBuYjAiMwWq
KJOugED+femEBr5O1yieG/2P7/eE1ylCe0HvbLeWuBH2vu43uEB8nnHhvqC1
K9VyU5wYjr1TRCFSTgajw6Gn07Rph8mihEmiu2LHnD4Put+gEHU7xUZ0fO90
5NnGrNQFQN0dAqcFirVowDXWByCgN75tE6MjkJ9bcyjfSnvWe4Nzr7FkALwL
jBMdRdnm35HMUREj4Hvb++EFpw8Bt+jSP71zyE5d+qHtWQx2GOtM77f7Ms+V
XuQweOB93p+teFUqRnjQ3tpYarFFYsgqsRkHYTQndaBpFGuWEW3yw1UBzB1U
9+Q2AE1ys7O9CTnl/kpqb35/v2ODj4aTq2HFuQjncmx6H84HsjX85c95sOLU
V6GLJgLP3tI271EyotvdCsOyTglAt8HmxDXimjIGDsrLnzqWUZYhC7FUX3fO
p2zK0VTzZDTYvprqm3zJlZfLlQRnmTmOPtQmRpehmyoDpv/0GcSmbxTurZ3Y
2nEGA3jC3MpJ8jz2Gmv4yCQx3B/sdzSwp6bcHaPKKCoK1+RscJL7nwHpAuyr
sIJqVLV9lfl7r4OcCPDNX7F7zilcjZbm3QVXoXNC4MP/5slY/ZUhSdxW1Hfa
DLZ8CSc6p5Vw3l3goahRNa7eZDmi+xqfSq/dOGfRnCBtMUy8LTYOThzEW0M6
kPSxLXJJYsLDd7QNtYV/O90V2mcQiaKRAApM5uCrSJwIJLXRXesBPRTx96B1
cV1omp89maB8PW1DGAICU27U7xNndGIiE2j8sVL393+a/ZEDD4NsePS2Xl9T
2b/lIfCd8rAvgaAiMhv4h0URsGzhcGylPvr+tr4R68E6kLw6UBAEnm1qOAnB
b6FbitpvfvMpbhD4IhyrjQNgDAG2J90KNXMnrCUqgTqCs/ZlBemBxbXxTTcp
DBIwhMvKWTRPXfU+6KimmC8JpE7nYopxfnktoclwrx1H88i/+/5LfDj1V6sP
yN/Uxpr54h1j77DtrIfmkxMyQ+7DrWeKXMyqvnBUbAewKfh++HfzurYsZhjn
9fkmeZeOzRvh+ybcYz+BDSvL7maNF8tFPvULVtZeQBhxaGho3eBvSiwY9Rnu
GGOl/TlIPVGf4RZLb78n1e4HbRPBz3qQc0l3H3qhCE8iYoFZrBVeNbsDrjtp
/BbanrNwJBLcq44hfwBwsp0DMC7wS9G6u67s9k4IQt18gPh9UIMX1zgsbesT
W3aVU8EwukOPUBffNgUGHQFkc9pysUSvoI9nTC2+E+Vf/uYYyZxErbxG4NXy
YZVfl0OH4Lii55pquzU7z1G0qNBiHMn9RvRrEky2AWiCVQdnaqD16JAM9Fat
3eFRx1/r8DP/G6zPDJq8uQ6ujlfzUEpiMBKlBJka68lz7pVd+zKxJwPQCm4i
8qoTmpUB/ItAP3CHHCiBz72WSsqrs+q3BIhLHqEqXpPP42p7K4AWYG/B88Nf
2qqcbuilsgPj98qn9JOi0gCZlSHaIAkS9VQA13LDbOYAxN2joDCHIdg3k0oW
f62uP+u3Xk+HGhLd6wxPIj+xLQnwpsnRgm4WHEIAAJJL+mMMlmmUNGWm5ZIV
RYmbSbOXqn3H4kzgwBjzdwvvI2eGas+xqYLoQntPOXsCCEtDFQ8XTXKLZjmn
qzzyrQErMYS/SBgrwEoHU67YESrnuNf+hRR5PEa/z+Mr6lzgw0QkfvNIJSrE
yp9qJUcXcQF1w6x3pBf8SJqcWPb/5on6H+O+rnXwW4RcN1cIs7ZhfipzAvmy
MnKOWY1Zjd7c+lwEGbIm5FkM1lvsQNff1qaTWC9/BuCfNnUTzBbCcuZlK4OL
wGyRk30yKe2Z4TzHMjWQS9KiT51WwBO2sQyY0+oWnMgHw1pWU+aimWb2pmnW
8J8tFnBZSNAuVoOfdKDmd18KfSsqJ/FyzRGW26ha3gp7ILdCqW+pFOl0wbBh
hzJvvOxuLmeE/ixsLLUeO0qCPUJTOKj6lJ+GmwvLTU3jodGpiUu16sUbFAea
hZX2yxsn6SEIRY1sYbY/FAEUn+Tht9sA+Z6a1E+5vuYAeJFbpaeN8mB1FULs
dX1yYwTJVX39PxAwe9AvnKN5/sNaB/mNuv/X/v+gt3IpXpJvIJhwNr7nqBYg
JqN+Mb/btnhS0dBeuu2hPCqt01r8m33FmgDHtNaAok67IqRcHcdotwGCtho9
Oz9AhJacOJKTyGhWL8SFrMkuNnmsXgg0Kowt0wFt2QZlCLTjKsJw0x0pQO9E
QkvFIpnucFiWbXmT2PlwbXChkJV1fcVMkVj3w0jjKEgoZ02cBftC1EsvGc/M
iGnI2G0U6Z4LI8e1zW7S7n+9+aVh04e2DTsGUv8+Yx0IC4Ep3kTJnsuNa7fn
4lTY+CJrCliT+AKopS9dQ8pyLAIQSPzsj0HqnbfPwgX8izoFbQoqsYOW0qOR
/CzcGUWSoZfZxsmZiRIPuWRKtL2btbnXR5dhy8g5O5XhAc2GalzO5/DTLgLH
t7lr0VSV5fUWHBit/lfWntoYtl0Hrm7E1v9Xaq+Q66vJhi6CYm50M4KLU+ln
D8loo2z/K1twEYwiYnJa8aE1JDoB61LtYbLzJzWWhXhWdt+4XFyOywTjfJsX
g7awIQkDRqJMOk4hFpO8e4fg60bs/rI8T4yuFI8D6SyyfUdENS3rbroR7UaU
hJD3VmHZOxQHpxjoBeta9+IBRWEfGto5DzlSZijj69ft0OnhjWwS5YkKYR5u
E9XEiXh+hH2SfvujbRo3Y46qRJPthfKxGCuIUsUBRlaYaFqs5aVJdfk6sqTz
vkN6TL5VAzbfWKoOLkhptG5MTN20QSVWG+aBwHGLXNyqgoU2/SkVo1Rs8+KD
KNOu5Uxo7PTqxqjmUGxfBe478h7UT1y8JJ+ZEYPHXVYtE7ccRlHapJkVi5ea
GaSKx0DzCn46ecXOyZm8DQfa641dPqXuq/WC5SjYI6FlwRu27Q9ZWYURbbIq
B2j5g9c4NmaWINPv+wwlk+Kf/fmk5XLHLTmrK/HSbg+L8hx6OqLlU5PdhOX2
+7YzONG63pdHDMQRQw5Q/dBbQtrtjBdNTSJtYSssRkzwxB9xppXNu6XehdQJ
/7uwY06bIcCOB+nRkOJN8nPy91Qgyn8hUC9ZtlMgE+IJ42AoyF2Hda2B5qrK
jo8esGutUt+FG3N75UI+COhnXWgSyW6qZ8Xs/SN/uh3LztN15mrPqcphF3qJ
9vVYukQ1++n965VHuy5s+XAB9CJfRNpi9ltcQ+GBA8q0Uu1XeA2cobe/BRsr
wORN/7D0aP9GLlOR1r54jOWDt4CoNcFq9WGImL9rBsdPlKM6oOnf4BA23i89
3TDLsXQbDgG8EmyxsdTqZrhS8qHBoeDjNexWKeYVOmHYePvO1Xpm3mKOYi5X
qlmo5Puf7jhof11H+x/uNWpG/sB0BCGa4LxO2PNRFnDItj9TAbtpVnXttGUQ
IEbpqfXuI1gbSR3+4Jcp9cVWXU8XY6RgrxMlHGuBaI4t4MyFuDZK4ufMVRBQ
TInjpgIVFTje9xi0rPIWCTKC45zXqs+B+PTJISZLFc62xybfliPiYk7o7tfO
DbXZ+hX0S4Hkr2nTFygArAKIC7VGDCeSr+FlrT1ejeimefvQ5785Z3KPSlye
abKAhaAAq2Nx9ao0vBu9KGnHDD59R4XaQTwyzzFFtLbocOHKxo/fHaQYgczn
5+uRbSAKRu5BKlW8pQ8aM0pVMV+9roXfxa5S+SZkVvbMHmEcJPZYJzvTd3Rr
XuVIGnGbjAjrTTOleOq5ovicBxPQjkOF6w73sSXeWrbrZfG/j9d1LlllNSN+
8Hv6CEMk2GUTy48YHSjhfZnFIGefeFx2TeogIJAscTxkRqIc5O5jft++z5WG
gAAP/qZ7AY2L/jEn/jRDcNNe1eqPk4Y+UGkU2kXDyQIKzc7r+29w3fW72CXS
dqjsUYcaybjl+jAFJflbrO0hbE+4MG98w1K1+wOgLjM3V/SxmP+SYdD+y7Ve
TIDHpgSeWurPhjEAIqV1xTtSsbh9G0hUUV3gUpfOv7Yhr6c7G6GEU89lSqIn
CMqHurxSQZClakOeVv7E/+8DWiDVHQWxoUZYzn21zHU4H+jObBO3IInJo3nv
NKHdDGd8JtM8e+DPpp6Uk3rV+ujS6/1Dtgz2njBWHYHxotl+vMqpcaggiuYB
ZfwHc6L8p42ysd5NTch8bRx1BuhAiCqTEKQPTj4Ts0NuQlqznYmIGjdyrsFD
XyBzw90dZ7EY29LLvf54L5sEug4k4ckhq2tY5gJDhL+ttkYjKjuhT/yNb2H5
NRkA1CVq8zog+BFchO2QqYfMZntK531g38yCChpW44jb7VrR3dhoisd+DsBt
LEBFpYk3TmejhkqVxJcZZjWxEVb4p9iOoyzz5WAIVrjJG094y0TX6xLxcD5A
kkck6XuGWtQYzERMEEuNFHgj+DMLYxXvnJ/jIH6nYoXllSHpNZjEQwRpRU5o
PoooEjkPQzVaMDLVDllB747wlcndfwTOFw6ZqR+jyPss7edvomwFaQVhnHgy
81JADOpZDpdLckjWcLO9XkjOqnn3lt2kzUMdsTYHQt7AYfjhLSwJjmmPmR9z
sr71vchsw5S8YJeokP4xRnpFWFusX03e3S7K7nkKnjiYyEm62HfiYXvnr+kZ
bbeEz4ub9++E7EJtlmJLPw2b7Kojhc0oB8mmvo8qmAskwi7l3rhkC0kC8o8R
0LB8bQ6XSLW2Fpj3r3tTb9VXjFaqhDQxLJ1Mr/rdeGCMGdDGvKckMV1sE6uT
YER7LickDPP4p46Wl9/j/GSEXYb5YGZnX/iillLf6lgq60Cxb9arp52X11mj
FYTMuQu8bMU3z1rpgBJC12XnU7UlyKYZeJQhlSnG5ibDx8OvtGdKyhu/2P72
OV5stgH/JTaTMu3k/xevzI69w6MIWh+jcJe4qOACOaKU399wAuSObmpFEJfi
gPtll2UkmGl3eQ6j1SXW/ide7rMQ5rM/H6DEBZum1cQWFD/a2G44oxa3C40x
tzNk8hNv1XIjvuH5qoNulshNfnWeyjRwN40PpTjh7y/yD/jZkUnD248juQIJ
7mZFLHDE5CqHq3G8Yo6+tVt5vM/hHbB/76JoV8OMAU64T2rPmtMkX/7G0w8/
EZyH0IziaTJW6oFWOUO/HqYJV/515NHGsa8xmbUlkdODnCr0ehlz/2pNhPeh
QfqgK+ywIPxOS30S/hjzHKfA2kQxNuflr4rTXQXlEfOLIXkbkR44p8Yg/YHe
w76h0nHS310u2nVqtCKMzLr8sCHfw76lscKIso/Jt33tX9HKzTxu3uy+egbL
s4TyAbxVsjoZYk6Rd7Uw7Rg7RC2D6TD3PfoC23zY0Et4GOaTwacLevwl9Ztu
Zby/TjBiD+LTpwaiYJpQCL+oFvofQUZxAnIS3uE8zkHb285kE2Qk8IaJzCxF
4VEFWNJ4GYaTLRFPVU3/lvJIMzb9K7qfhtSnTD5ZWmB1LwtRMFsC4YDCL89J
sp4FnO+uprshs/bmudC7WN80C9uA0F1huBfmBv95eJVsBQBkVFCdjvxaxG8F
t8Vy5VcJ0Uny+EjiT/YbMCtM4D3d7UQ2m2T9ZcuaJoeFLHnT9xrY8dIYmC1U
nblAeCRbPvrHyOkYWIEJub+pw79szUjh2FV3EQZgEx1pb9ohqrxScgWPLqr8
n+dR2mHLyxI58FVbdH5Y+0pjb2SEHH6/bOuN+CngNhQOtChBZ6U0Rs2VeG9Y
4g4LmBOszaS0v15Nq8K9Y625HFj2+6sAs2cX36/6Kra3ZAJdk9nZSfCRvZdQ
Ivw2jXAXeyCgxeOG+Saci6+Jp8PaW11qMh3WBD2XnqKMZnijR+lE96X05giK
LL5mNIJsotImilfebjdDNfVlP2oVXn3/g9c1Qz6Devde6LWKu1Pnztecb+xr
dMH4rdjijfFOa61YaprHa51z+xJquEdAXt5XuwnCg7oS9SIYf7JIn/UZc3Ov
/QkCcU2p6iITa6YIBmi6zRVnQXd+Eaiz12Xcsk0rKPW4Mzo4FeTZqEHepHol
EpxgpUVr/M0EfQ9cRVZJzsbB+NMARB9TCKyJ+1f9/vvmNI5bxXaLeyHPBhFx
BAtLqaBjBbYTomyggkDyrPqCS7XYui4DtN/ipFhBaXY1gWjEDXm4U2vkMvUV
ZpvIJu5Uz2cEwG2QpYgcVsxrSM3BXnGCwEyVRh0wv6cwh00wbFsYlNcPQOEN
v8fNnnxOuZ6dFs82rM6mT8HC8cXSw7mZSDlFE6DT1EI1nBynGHfe1afhofE5
FSmVIXhEArDYAe34lOZ/FYMpztL1af2sZKHTJPkFJKuMarQAmXqK4AYdQhXV
ifORjc2q1iy5IrONm9HP86MyUXozEqMilfuddguZ7csfZHye8Ic0EI4ZHaxE
VwPZ/mJpead1pBDTF8Yxe0nHFrBqP9aLAmOwiKjti5hwnMaTqh3lTkk2p6Pw
njkRo2cJMliIxkSjmT8EPsORgknD+L1s9eQ5Coha7ACBx891E+j6uR88YkGE
Mvg1vT4FVWH+txdrvtb7sNZBqeJsAu8+vGZI0e03zPUDBjzf8z3D4W2ALy9Q
w2iwSL4FrHCTcft18vLgDkjaXVrQYbIHHxiY8SSsu90Duwy17wlaemM9b1tl
0sacpBTPSQcDE/haerK6a7JRw+iYecigir/NW3Bs9m/BsL8x/qygL5UqLW9m
MvIsfMFQQ+Y3SXzIc4+Mfs7xTn4Kdx6OZwdmJcgfmtHmPutEyuSXLtT3FXoJ
qK/SZ70XzgUbB/mflSgxhtDTaG+tBx+CWVPOo1/z5OtE6JP2RPUPL7YjQ+lz
/q6J6GfQqrN/5MpXoHSwv8hQq/dG4bCa5OIOJph2v/MbZmLzc2+ENnMkVzl6
PGNoinxoolQidohmTpXcqIV3VPw3R0ljlJALmzjNiQMDoCK+M2+RPTmdB4xR
Hh+e4p4O6PjcSzdHN69dz+W/3Jou0B/OIb4Ha6juOh7EHzSo0oC+ACQt8SD3
7Ke+4TXIFYzJ9/AQAIWVtZHOpOQH0VopmLxToy4tfF5GqTiiWOWcUgypbWcc
vz6OYplLk5z5ypilefpetl+fAV0iuGWezIMLr7Fqdm7fbkCYPzLFiEEVvbum
ee0AsYy9UUssD05rWMXmM41A0TND1/L93aRJhqw/GDDJb+TKcPSNzBFto9g/
FVQScv6BF1jdGFsKjax84V2dMgvEkeA//jlH9e0gwyz0aGgTtgnyquc052Lu
ByHJXIFz3/sIXoQVUxbE+lxy95NgSvfuXsOFpcGYPgwc9vffgu89zAjZC0ZX
Hx1nd4swxjlmXXWOa0GjKmcDUmvs/EmQmOwGujK7ZjGo+pcZE9oO+wanwTE1
3OM+tLX1K2by931KR0HfwbSCkK4LBOZpxsfdfbSN49UT6kUVqYKl0RLCnwpV
dO/LJQ/GAeg0TOxjn+jb2mz860lDk4h+SU0fHKj0up7fv/7HzfVnqoXzFtxN
DMgMHsDpLrWtP2yvHxXsVGQDpYKTMWcc/oLbI7OJZU95fL07ZAlI9IOJ8rIb
UN6b0VtNg0BpTOQVKnEyUGKT0toDnQ0D1WB5m7SONIsm3cGfR9TPxs3TQ4rs
QhQGaAdA6fBqlFJAyAK2sQHmS+fUj5+DXvti8k2QSDH/l3Go0jyArg8Rn+sy
pnnteqP53Mg2PRWJnBxTQPAa3t/k0vky8BG3t3+ZU9HxUJCfpCW0BG6vlm+O
49oUzi4SEPmkQZn4EQxDJJhzAK3cQFpQg5udIZSJCUJqU97akMdDblOc+iE3
myEugXeDMwqCPe/I4RKdIFGxfA3ryBfv4g0aA4W3Qi+5NBfBnrE/ZnCjKBoH
VXcmmZh+F0mEWJGrhw6S+W0Nrs4B2VMS5jk6AfcbayLR7MULZigmqD9UX/+E
M8sadREwwosBkhKY3JUAbXOhPCuxvIhdesL+9ebGTeDvBvMivGz6OJJr2ouH
U0+kVss9YcuJat0zwjHXaNCD9koxmuUxjcQabj2JTJuhbRTObyKQyXOihX6G
YHrZ7IYKxgqOFnFpH1VNRMf+Yqa1mEXWCME4tSsgk4OD++n/HjKlObii46A+
spIlHhI89s+d2NXQHNEkd3cdILBblamXkWUyFnw6q2HPFASmOZmdiMYnNNcf
onfNMWbZhcM0/xpPtIOmvwK25GPQWvXoJt8ZIynp/1W1h5k0ebq1eWvdRMiq
H7xtgK76ZddpnhJCrqiqcWZQi9oIOw5xRL1LB02I37mC/Ai7/8fS4z14QAKv
BNtIiv4nvUTKtMwGAAaHKOHLyjJu7g132TQVzuitb46RXCPbuka+9sEskzNZ
6/DjbUu7OpjFnGMasuEmddAlkH2ZcTbqqApkwaQrzwmevk3QdJhDm116y2LN
jjOSsYZY18MqP7UuRGs2gcCs7EzQIB8ousH3vrx8EdRLdMdgvIlWo0k1UKcu
lSDYBGoCLU/eWwssTpx/6NxYDl8w2zS6H0EzQWTNXXazNXGxl8NfaQBp/6nE
KJ+G3/qwHVoJkNkeXNkK+cwYnl/EAlw4HdWm+LW+vkHBPne+T2cv+DfYbJLe
VrhAxBfH3G+b2Za+9cVE3zcrjVgcGgNNcX2WZG8UCRbh4Yjnuiy7sre5YGm7
3X9shaJ4KLaq+lAiSvKLWhy/Be7yCcbt3DaO0ElNKCNEC1dRIIAwBo0B/9kW
RxmexTItYTT0nR8tTX9YFrsfZO/nWb/VOhXgCDclgcpvOsxQr3MRz2xJIhHo
Pc/XnQ86G3HgtNYffslrEre4H1TMVZcdcq6GRYk9Wm5CzEkkLNqy4/VkMgnP
v8YLXX+QBIKpW+PTjvp6/pm0WPPpfWIJ2Ch4dEBTB2LHnQ9BvGcSdyJCu3sq
76FRBviMFqJAIBxyX3ujhuXX4L3jXdRdoKEEFxHpJqHkT7i6YahAebeYBGV6
9QP3nBgEEeZZNTrlGptsMP3NF1p3RhBrOMc7K16uaqDaXiH8salsWKS9gffj
ctdHhQ5kzIwKD/ljXfM/l4G0EA/H0FGKFgn7Zp9KRuZKtCJcBgruyNiaE8Gs
ApHSthX+JtnhGt4oppw20uTTERyLDqYEatwp1hqRElnrGd6JkVqD0FyE8fHR
CMkX5LqBFeCryTGfPlOevft5uOppq0TZq/HJC4BMIxamLNyv9MyszWbMyozP
SHpnHkUhrJ5FR+HHpd+j/3Rr2zMcSE5RBSi+U4zcQVBGAtV7mVfFqR4glg86
jshfRBMmYk5h/pLn7Csv6ipQe6Kg7DUczGeG6aEvMV33QwyCKHhHAi44S573
t6+R65qehyWhjQw8m0bv/wYSZnW7nQmFi7LqSVJl52ItiVEJQQx4uVoSt7Zc
IqZsoYiO/qmmHbJeyEhC/G8u3ouaQo5Okh6Ds5d6rmf4ZxreRjxJZE2MpJ19
fwYno4pR1BSzcYu2d9wzPDLDKR5LH9JHBqOn3lZ9TENxdzxA+X8Bs+IZmHEC
Bt30R9Qa+dZyhD3Vnx9S0cLpUXgMZBx06WErJJDRVVvZE6Au+2U3/IL7c/0s
WJcmj9aQmAtkVVyQlISj0QdOoCDnnnPV+UgSJBfoWvTRn9fgoMJiB8m5hP7P
DJ4f1+VKqQpW5eKkDeZ+jmWkkffX7NYQnRO57ToaoNWx92kecV72R8fV/LIW
5EH3j0SFTYtlFWA9sLXZNuyNkIA+1PXHSOWkwczBiw1j1a3SUqbODHbqTTM+
nD4OOVrNv56lhDFuyL3HIiAzn3hqHIIvP7O7MAZr6XLcwBRzDYoF1Elrx5qM
gxsen9mwJzX5W0UBHtIc+wrm1aSfSPXOu/gXxBKX0EBwW9RB+mayStoZ77dt
2mTAKBVFKPX5Vocmb1fX+5LUmm2rl18/F0rWX4y/Gbsn6s6nbrhG+Y2EDj3H
fA0yLZp2KFV+exvm554W19/N7MSYoANlK/zo5D1XvO6BiT3ezW/ivNtQGadx
EYg+6nmL959bNah2+SSizehPLuSipk2FZ7Eu+XBBrDBrwLaggDcbA3Zhw/Fq
6ZDKb04qvqozRW2bMK+9EuKNtTgnZAbHx+GPYst8wqugeLdmVNkqc53shvx9
SZAzG43xGXsdNDtogVqG14t5+lUDx/lQLARUxVVMgWx4DgwVZL5Na78IUuuf
DBzrLW9UVXgczDV26REga3N6mU/vOkb+vG/s8e75k7Fm5IBC0CVgRva6i678
Z3O4CFGTQuR/OmfCGn7ahCaeDODWFcQYUZ0OY915+1OwddQnLDi/cRRVyDPG
yAtzoqpRYQ4fxJFJka/EHcSgTRcDi6uAzWNiO9jk5rGFAJXwBQ+unuodzYwA
JVOD+/OXG+gj9E03KXqo1Bi517eP7X6tT20lAXFKxdeGihrWqAeozrHUpCap
2YrU6t+CDwvSTc6a6+qQdxnYIZ7XiVnjR8l398fSIpkl7DSQTpwYLdEcibZu
xP9GE9tYaR/r/ZVWrjcq7ABwdxJR5sSuHFMXO7/S/F9XVjUf3WM5CS3v/AnP
EBPnbOb/AP/ZF2kz7W8+1F9bQbN+4mkeXESQLyIGuH3KaWiLFIM4Q+LrQ9VP
FGFqZhX0JPA1Oxlxd/Br7+vZYxY+O1dsPopTywCJX4EQ45cOz4NVaR+ZxSh/
CfKp/s08r8jzXWRzlg/bnfwfPYG5T4o/7zCN/X9FzpPT46xoOxzdIeIcs0rn
x1NtRAOyKvGB3zR0mwBLAidJPr2wJ962xNHHAjM0tnkR2++5x/7lql4L7aYW
fQZlsHIj+FxjOXA5R1E7BeHcjh8EKT5ZV3OdtNVNNa6gyiOcs6/gMU16opH/
FS3m0KQtI90JqnzZsEcOtJZEDKblIqTreQhZk7NsiYQC5Xtv7FeO0/+cGApI
LWK+jTSwPYmnZe/6qYenDBjq6gsloK+xhwJOuIICxLSkJwRJoM/nJRGmpxCx
otIHqzAfVKQm0irLvgSpAjIXUPU5v82daopx5i4UFiiFo+IzrcWT/8++Lwzf
BDFw7GkyOUAqSew6SkbWVh8ihMGP+PlaZ+p6X1Gaxnrscom9ld8YCpsXoXCE
dOc5avcKcfo+GU5e3Xx5cD9oGBJQEDnZlG7gQsKWRpGWJ6x9eRqOLGrgddBs
NuRWFw0ewJXKv6p1m7IcYPJ/Gcj1AIzjhqPuJQdhFzPUAWkQpNdBxQPKMFyZ
BpTLNCU65LozbTgEjrIpvnBoG4eQVGsuduQIhqkMrOcP8cAkm8NMvwaP/tzn
xoQDOWR0vZkmv9RheKZTN8GPTJ3dexlTGWCS6b1FEk85E61TGNJiB0ZpKR8o
dee14queCFBvgICWbvG4gawfeJ1h/vVwEJhOLBgjm+9ruLnlfafV/6ZsobdK
Kr/kdF0i/PK56eutewuq2wSW38RnUklmTpTcfYQ2qEhaEgJTgxdqAmJJeoRt
wWRO8UKkgSP441U19nbrZOFD3SBTKWPUeddBkhvzBbwYan1+S9dNONrDOuCv
XvZpn0/fsGv9erhtfvQ1WiL/PHUf1OdThC3BvNl1kL4vNB9FhE8L7aWN+2qs
pT9Gbf4kHl5ny//eYNuFJvkMIhNaWwGIYH12MNJTUwiTHMauRJG9zRvOMz9S
faoZVk3liw8rN9vfl261vsTvFrYdmDs/Y2UeLSMCld3L7jN9bol/ASQR31mj
AY/kxsLdDDeCN25DBFzg4k+3UZDnl2hz7lnOYORKScdNN/npaI34vpjLFl6Q
KI6k/PjoAizurijpcdSrRAI7UMlxImRbt2IsQmQQ1P3rZJL46/gOY8AiM0X2
13ziHadmNegMQHpEIHQA52P+3z0UG0lC1mMRtE2igcJqxL8cpmBCUTz0WjWk
9kH8rdnol/lJ5TBUbKMbOAUM/j2ubGYHUkXlau6Hj1+x+HlmKk8LaLe0cCW/
4QRa34/NbkA5nWxjwjSbAZGV2yboaMgKFXgIBRkz3Qzamg/bz63G41XsUFVF
TBkOzOR5W6CtoN5C4muzmWB2Mo192Aio/rxu0RA4L74Yjs7AKxrDDSuZh+KI
MrlIx0Cup9dUArvkYXc0i9IJZLt0TCPK9E3PlYKnJzsk0YaiRCsvLFoxAZlB
eAjUcAJOHWAzvse4yMqfi0EEkphaUshs8Q2MPsZhxXZZymQCGDniP8iR/q0y
scv8AecYF/8gomQlnZXKxQop5PslOfy/AFmrpBQQcfjHgQj0HaiPVFCg555P
k/ZVORayO4LIERyl8Q054KBBRwgVw/mEcUKQoS/wlbwliizFs7zrDYshBnXE
LBlHtMCwg78n1SEBNZwvCk6tHNn5y6v8F5dRFxP//ecN5VoXUET+bSve9rG4
nu3SNdQIeIFXsQwrlKmLH7/OcXK64iOnvfu01BveEOh03CC5nNr2x0oT9EfW
+jJAMYBAaNnihMInDKWRnX3bEmyy+CbMmetdpRqzYu71O6uhAT55vJspcA3l
Pd12Ar9jRzF/pkbTdTqwRmDRXmrt95TkAkKzwP1x3BlVA/6aF17QuHfzWFFG
AD9pUsu/mpBBUtDeQxBmOaACfcuL6WwqCdiC8aL17abX3+TW2qfvhsfjk5PZ
fbndAfcHLOS6d+UffcJm1IlxpD1pp9b5mw+o06g8/EO+cxIGjcWxTGz18Z0S
plb7n7gY2HJUOa0XGN36rx7VIYxbSBV/NKGyZwC9Si4oEliZ4SKBj1/KBelf
6ifqnpAD6ZVrPvdNDHmMX6+Qcu9xkivyxH1uJosB2KMBblaQXgIUm6oJjIcO
2b9EKthwN/KF3g1SizpyI929jSMtuBXmvu9O7rJ56aThEPkZCmBh57S34hiO
xVY49Jbzp2x05CuMnwPxKMZjUYiQtSqlFdYyYcYjU3BwzEqk7lg5kyRHI1Kc
YllzoD3NJYahXsh65DO8tpgSZnoPujT4YgV+9jJ/DRuSEFxN2f0nYm6sEcbF
Mf/Jg6nY8UhoYV2Az/8Noax30eaoulXklFPNbF+LJ5jBvVsjDSIiGVYPDAZ/
eGkMvb2XbbFat2q5T7zVna3qTppnNGCP8p5l4ADtHBMevOIXKz51Pioa5HI4
PttGLNCcvv7F14tE95guVux2cVkHC4n28xRtXcPIPeSKyL/cE+voCgxN3wlF
sGKWk6c0PPjXBUsIxaEZyL8rXMu/Awz94H7jFlag0jNuhcNjkFkIfGt9eBOK
nCg4YkPFY+dWRiMaYfiY3oKia8agpfO6oPm9ajQiaEuJCDg+FyguaZpdS0CZ
bUWQhEhkG1Zi9DAbUA7pW2dYL0AP/k5zwAWqRjzUE85x3fK4Uy/Gg4p9xlGN
v+MfWbyjLQ9gVIlGi/Qy7Q5Rc3sGqiMxrJSKclwRvqJHw4VNiX5kIvqEwZ00
zkm6o2HZjQzvRceS3MDJXLsLd9HwnQxsxitP+2XHx9HqnU+0A8ccN9uOjYZ6
zCipAD2UYhZaz4gxHhooNTEaPc+dZkfu3x6ac35h5bc4KviFUMbbUqzcEBWL
hY+6CYbZeyrLAUy+7Y7DwJPqEDex4CHvVrrR2VCyZGASTVD1d3ns2DxWTG4j
wfDp9DoaqdPlq5laagHc9Ja6uDOcIQ9JIcLAVLT8qaRZse6RI6Ki7//XltuC
zyioR6uIEDBHD1bAi0SeWDvqj7U2U/h5h+IMIlOg11hXN0ZuPUlLrRYDmID4
VSE31vEfMxrcFuFjNtcM7bs2Elyc5zPlc6S9GD15QBuxAIm/9PKkiVsjT2Qv
ew0P1z86FNDM63g+7XnqVT2jAZ1kb0ylzQP5oWZU5o/MGkUELHvp96tc1Ua+
/fB19mO06QwCTFTQ2FUBgjk4i3dUqMTtxUuuZbE54S5ip8fa5wHMBrOG8cQx
10EMONLyQ3agFBNhN3AEWegPoNuRU/QszSCrpidGuRh29Q+ZGlzngBkxyRct
XCJin/nUcwM7agAUp6bkHwT90qL5LVkxqkE+kVkaDMD2fB/gWpCeO4DnKf/z
gU2dz4dMnoAtWaMx07JOnD70MxeiAcMNQY9zp/4MM6Ad72PZddUjg3kNAXRF
aixZg8+7rSV8+mfozGUz2Xpc4nJtTgvbTITKT8q+raRhsKUQKpL4naCd6JzH
9xHoxZeC2MfbFZPsYAA4tIysZshSx7kO/rFtM80ABgjQOWU5etsh/d9iPOhW
xDjelXrJ+a8nm1WjjCwXtoufNugTiQpznDodtrXekE9qZSn6bH/8aUARe52C
ODu2i8/aCJaZr29se8jVaKNFR3vqwiQjx4mLgBvz0gTMF82ChQI/jrJz3w5l
nD57KNspLPykys0rW/mszTWFAMsHzfMeiz+B2vkQQ0DausHV3BQMIAmtnKGt
Zl9Mt3go0E/CGrpES5MiYlPZHfJSKi+NtsWxjc/UDFhKS3fOL9obvmZ1cUI/
CHDFR+oo5kjlDkxMDntXh0EMJJUW6JafkQpt7k1FNit6ZfWOFEXSFR/3ls4+
sdVDrNEUvi9fJCY5mun1bIxnyzIV4PzvyOHtZhmpYZ3C1cPcP4qGLhTIlHbA
R+nfu+fUxgKImLuVH0SrCBHwyzN+o71Lua7G9QnwW5n4TSLRY9lR1uyu7xY8
Sr4T05dYNT14Sr62xmmHx3UUkQbyKFZMius3baL+bpicYibZ9M40A8lX9C/6
GNQxvi6hLHTSqgs6Or/jcsqUVWeND/EH8qBF9s2HmOQPLSQdahmDu/T6DsXK
dFG+PRe+kanTsY5jQBQco21BsBJkUaH/LfKEEjonTY6R59769Bpbq6s251Dn
O70n1euYIvgzYXTs87R1uv1CH7NkxfzObRVEzJdaVpccoKVX6E1+cUQn3Hs6
veIYedHTzAXfZegYmp+JSDgNO5C8dCvvio/PBU3nJAQxou42NUQHKM7dSNkq
dhiX29OyrT5YydmVQIVJL+YIGr05/UUYTvEtpZC0lHHdPQ8lVVEdhYj19Byx
dYdEDwac0BpL8/5GKUPMM4csBHLLMRxSlooHGyCA3C05z0AzdbFj7q84LUJU
uX49PMY57w6AlQouO/4nElC1PsrqYDJdeLKlxbzlNgVjnMkI/q4+RcMVxILU
uFJ4RelKW872thQ8drWhCSMw7z5U1ZnoqADvrYDEB2TIFTPCiH6giLo+Wgkt
JfmBTRYxcT8Rl+SCJO4EaD9P3ikiqhbnAXXNXSCq+tv3DrT6EwXiov+VHWT1
layQxnawvzUi7sMJFNwsqxwq9edLY7la/TEJX9MuCrcdF9QsM5mxgXnBY4ck
UUkmdTubd5LsrzmN7XunLfjV4t+Nxe2NJtrhpQxEu7Sb/jrOM+9OBu5kVzN/
OyCqvnczk6zV8GPsXpPIcYA1fJrO0r77kS1VMviZ2olTNw8alR0j4ceumoHL
9M6hdflwOdeP4rbClMMDYqDyHtaq2safUwyEC3HTK5WkY7OFCixMH3oP4CGb
s5MGxfQ74+sES5TTjSYwX/mClQw+HMKGcqNNgWmOgRMzw580gwdlhEQaRJ97
JJBW511L5MM22Ut621cqYKoh0mT8kyRwMxX3IpEtyxwfr4Kb2wKyJw5q8Z1p
TTQe4XbwnRNIaGJlTaXCwxSYgh2RVzZ7yAQ4kwTn5RpxXk/+1ahdGaAPtGCg
mj2lt6Z9xENwdnCCFz2mNszVp1fVVmpU5xrwFgcqQYegPqQWhenFp3693Ulo
82SD55OWAv/BPP8pSCJr9ltcdRunYnLjUZY3gFvqlzefbKV8IiooglBezC6p
gm6Whrz/dN/bkzjqvbo2CeosI8DqD2LNpiJ9sn/3TZKAtpEZnM2Vn43GNPtn
TQfIZRtSRMRBR+5cbox67rmJzQUKlEYVQ0Vel9OsyF8DjcZIw+GZ8WMPD3Pg
1v05m2mQK3QYBhJ44fXQGlEmlIHBMi49fUfAh7rrMXFXSV1eB+e+LD6Eb4pv
z2siSPti+7LLAHIzSZMj1pqvMa7YAixDIaPeRRmNgx5kngTHrqD50Ni94L+0
h5vzyibNRdqpfAmzOHkKaCefuDL6sptEOuXSE7VrZilBDB/WyyV65VRZqLWB
OsawK6fOW+KYUOjuaksBfKp1cAVCnXvwygQkGe5aoUqsMu6A4uS4dRIE04IT
cXv3vO0ZTERJqn+wLh4TU7e/uOGX9uo0yHjHxU+OLeMRC37AOeZi833eco0T
v4LzJkcQNb/EaLRvZ5pmF2jzwiTG/72evKJ/A6Y8zt6ii0Y6oG9GQ/PFvw7+
aB7ShT39ja2bUcu0lb795oGAsVHs2FNEy48qBuk5ItFDjO7yDc1eyG/3VDmC
QeKd0tvXfgLb/oGgg2kWjf8jDg+6MXKpZDFjEXuRe0YPobIA+ZYX6jdTmW7x
poTQX2hLrImjITTa/MTI6ZMypJRs7lHDvlz4vkSPJjjMk0p68F9G4pJim35H
zkMjuv11UENlI352eMlypOp+SRh/m4uqxSoBn+VUQu3qSBG6RJ1qr4+eGCAo
AC/jfw+PbxFl6ahe+xYiOrJaLIY7wtPhKkiouIfREb5D+yzGxUPZOSpV3CfW
VWjTRfdhnpv4ub9nHTxFs4wiyFK03rbnvJy1d1+91eZvNyebmzH9vlVWL8On
gyfYcdGZwGv+D10L/tGealz6JpjX1n21WztYrGQSqw0XfobBSDWvVUIw+qdA
hFdZlVZE8qCR5G90rL3rO8ogJvc7P+SRIGDvKp/k6A9U7DKzn/IuymyySkvo
VdT80hFRA0UQBWI1XrupqXZnxqboX7H3ZHYHohRHrPkrxfHDKlWI78yuO5e8
9s9qFI8PvKsrNSV5VmBbXCuePRSERML1YEIyWGxIFjsN27WMPrqAudiebdCG
BxzwToWdmYQiM9p+797XVMdzkRrUi1WCHUv9HU50iuiksNd1ykRBqGtOAn4K
v21U44AB36whcJ5u7vvsFuoE4icC11Np0nh9vunPD6x3egd2ZkC6OKDaKnLS
SzrnoXlWH5hlaJIsNY/xrt5X6IL66M1LC7BW8ET4p1RMV68RFC7I/+Yy3mBx
A0TQ8AQkDJHC7ys9vKuQa4XQTP0D7p3htflZmGPqdAfbpnVlis+e4VfOSx2h
F2DrFZDVzDw0e+8D7Cl4rpetdOJ9wa2FfMskKGq+b3m2eGjpsiFAz3QHZD9K
BLd/qa5+bC8qKhmApn+J7XlE1pXjQZDuvADzkIlkDHwAPQAEXpYf7xv0XQ7w
mH+IMyViYhVM7OOkVuKu8mMORdp9M+VgemiWCP0zHDKijjXJAEtHb/q7lErv
7lC606bPB7LBXZB96GcGtCtPdOg8Qm3ln+t+PZ3DO05bpCBnIuR6H+v58sCC
TwfLgw8cCl9eHl0XBXxcoHdLB9OqQzxuHIEmSjOkYVWKHqinbDno4UtlJux4
s6+MY9g40zEYk82sy+cZXKRIYOGgQrOu/GyMOCnvpF8I1oOM24uAuyDJr90L
Jxz65QP3BPxZOk7V5zJ0y44YV6noKsHqrVCjDNUPQ1VE/dcHzXSulqvIkKY9
SGudBvpfwFsiFjukfxZFTRansPh+TwKC4baM6hrIVHMGQpt+8gNs+1B0qS5i
68wlJBv3UMal4pC4aJ/LhrFpK+oZlPiMJhssMiVHLGHzGQ73Lay/UPW/lbgb
G58sLhsO1SiosHcE8VgNZaDc/1OzlOfrT6XK2Gbnjcn26ExiPpgsJCs2jNSv
kGhEc7obQiknHZZFe3RSVz4u3bkSuE63dvmuTur8uh28O3RvGNruYN4r5JwN
WFIl/05OvFsyFYPfj4xr+gPWFsYDSBHMzZBkcUqiS+br2nUap+jrQ0JVu9Do
oT06k9Buk59kxICqJGZFeY0xfUqmFex3LvGJzKi2t0KRMFgbNE1RKWNTPLBa
VPduYZx2cy0sfD/2DBgY5cXUkLvPE41ZfhlAkW7MvwMOlcKX9lHrSZXhkDC8
Px3biQ09FKYYBXcN8UxlebDnBR+MTupYjxdqQudjIIA1QtVlynRIe+vdZdRo
2givInl7q0xEJQTgurC9MsBNHYENOHwhlDT7AEsyhOjv/emaHDcSoyHJcGIS
kxIVr0NPB7FouEMifFsoIWEmT2s2ozUPTHCLOFs5iI+20gZiBiTUoEiDlScW
MaiVo0ihtASl09COKvALVG7fsJrtt5yI7XRSC07mQ9wWJQGmolvGx7VFUePt
Scyee0v/2oNv1Qyvsw2LdwpzdptUAW63vRY5Mq0Rv0gDI9ov0pedwsic7sOD
7E3Iv4pelg/RQdSjxPqcR761MnprRcbQADSjtErPmzDiyJFwa1p7Ita6MSmX
pRJsIIjlK0sJnXuaBZwPJJAr9pV6lwsTBkWstbe0qOkUIjgHVQ+aSiDvZ31/
+Eo+UHBUPt8DEO/f1nQ5pKvFP4WBB2mGEjKdC1uwz94hBHjCnSUDXbEpZXzt
3lq+d4/nd8JPjofzTx9q2OVElTfva0Is2TnjtlGjiH5TE6gLFFxm7SaQ2wFV
/DntMQWi/LOFmZDvdFB1VjAKCx74Y0bAHPEVe19ixQWZsH91t2gGe1b41A6t
mVyt5jA1/LM7kgdXpqgqe3cKgOFaMHFHEYPWsd+i+THmlRy7XgoHH+Sl9wf5
tl70ggFQ9ploNB+l2vY22qyGmF18X4UosKVfuXY51XiU5+EYiONqvNTp2YIK
yhSBVaaxJkZMUJVQAeCEHuo/MYAU1LZD8N2iPmhRD0G3dH8/CgvW309Onwcf
KBXAPqJaAilzcwbKre5FztEaxOMxS0yS+krBLEJHqSzUoINvSCwBKYUu9MiX
uxPqa32YtvhUYDG/XLK+JONGFQjqyUXfwl3ms8VnYMjKSyR0RAirBc+MPRan
NOrSmZU67pnQC2GPTw1Ig8OFBFM/GROKIV9Ln0YyKiUq+P7otXsnB/+ImATk
CvXvPve1+MedWnEu9+fUenJ4IjCE8EcAikiihPfKA8A4HBwgnucORE7W3V9k
2qF9NSw5PmNLu5zxQ5DMxm9D1PyMWw2WnOeW3aD9bmZxMYK1fQsvs0GMxADr
Z28xTnn1ql+1rkEU4mMYoqOtmvWFotqjUxVQH/GszLW0lUfYnIy/nX68/E2E
IZ1bfjEv0ztScjFJtij9pEiMN968FQYGrKgOdhRNkOS43GmQbcXre18B3qg5
BgUEngl+MthFDgMca5KJUW7uE8h1Sxe0jz57Ev0SgIC5alex9AlEDLVy5E9h
qnO4SQVmIXRCMVatjGF252KwRqJYZ8hc3jf3wp/9FBJdGTS0BYdAv37vVWOF
c9qcvsKCUaLPHesuM3aPH2/4lh7gUba4f5TT6HJEx1yXuLf0zRsRqQP7cz3+
/zg8LOszDBiUsho1d9lU4E/n77Drmsc3KLcS4xQc6fa35S6MRwb7xx9xk0vO
vmS7KL18Hg4XS/lVU8wuFb+DQN+vYxZW6FH4AL16BeomvTpAgDPoP6Oe4lyp
ECFhd8+PATsnz22WqGU37YwEYBDSkB10wQ57fLULa2jtrgXf8qClASkcp0Zj
kHxT5xJkZQFXn3reQtc7oSgzjjxo7bG3+oaC5q+Nejta5tAMwoDkqR47pZFY
cdPUDuC5XODOMTiS/5ETxc+HxG12u28rHZxA6BRlcr2t7i3zgr3jGoIMq425
0mwpf2o+FQXOfiUGl/BBZYTllePMzjWp65Vw0mbQBXVxige6co+vG5edi66o
BnZBiwfCq2L8unU2ThrDLj1PWF8cWaFjUwfgsetbGvT8u1mePKzbic2XCTx4
88eDw1PNP8Ea/eq6nyD+BJKVtH54nLfjLp+bez6hnn4Ngwl+d8vNuEbU/jvZ
xCWrx25C9npRwIKxHq9C925lUToOJGFKkTChXxfFlEPpeP3JAhBsyDaf2csc
42gua0JQpTCUZWPTWjprxxilu0B461Ldao8ec+Om59GunbS9vHfDR3jaOX0a
HyYI8amyAdbqWNdrj98i94LOFttsZ7KkbH1gyK2K6GiSTgvEMtp9JvpFRn45
ulWG2PKNBav/WzAfuUU+Tp3hBM2ODqzz6pFwOnZZzS6faKyA2yOmcJMB9AE0
nICKXvAuBh6lafKsgKxDOTqVURlkVm0XxY1bK1wJbIevlGvWJ7yDYRkov0ZK
IZIsEcFbwT5O64XuFijIw1hNlA0uIiDXIFecBVHgfXUT26cUW2aX4zW9w8OS
6HnNzjhipOjF8IQFMpPa5Few2Ogy1B6E/RLNzygN5wYUAD+m2VQz7ruVrfwi
Klv7lqdTbxkiLJJqAAEu1K/Wwsdl88ln1xa0HSCSnCIK/YfeUWG+ABaXzitW
tZRvSXvNGSArT6CV4ndZmHSMBrsSY1yyIz+bS9UMHZgppfl2uk8JcEI6ATYz
EgmEXiNL7rz5au3+FPfJI8MEBaRZpSA3OREmkHwSj6c7NiilWR3/tLmapGhH
/hiDEdSaQU4rfG4WGR2SQIYbDBIbpZyh96DY3xOusBzNcGUdvDbDzQhY0Ua/
B4/PMYAXSJ9uxy6PznZT574zZIhmXOsvPUPozl3FEtr2nUDsNSgfso997i1I
5cSMmlLxhLhZHLJmmuOG6UBtRZL92kUAB5eeYzSzlFNHav+LMDDC8noVtRjM
qdNj1lab3H64mc+Y2hj6/+HxUUlTRLFtowZcit/5WuSu37/IJVG+ZW+xAeOy
OiVdqToynghSkQQn0w/JkhQ+IpggtC5I4/kqbN6Dxsyk1OI8fE7sIhRhuNPA
vXPUzoD3jh44+KEkzPqrUUWYhL6LXP8sRQU6mkEs9Nm4a/Hwse6jXm5BO87n
PLWafiOWdaCYDtMypu8QlSfeWIHcXRodRgWyWOnpZ+6J0k0GRh318NM1QAcV
dSziut7+s5l6lwPX0SxZqqFKjcKIf15/LW7I/8kCIJYFiCMnUK7rwnuGg4Ub
SSSPuFDmpVq/J9437zuwxGYw1c/9fpUVrsyQszEA3p5FF06ZmHWNdUJT9scg
eczKUAGitMY/3460MCmhAB36D+mHqGkRzQkDnLRTJ/QJyzVli/wWeQnWeNdQ
dIVpFIcujw/ebENxFDd4IRAWMUNYLCsx2/ICZ5B+5YhUkUB1SO1++tPcCGLi
3Ky2vY7yvR1XdTj7247A3ihuDfIYmsiqzJSxzS2Qgm55P8XVUXzr/VyDh7jJ
PTuENoDnVk8tRhgKNcmYCZu8ZTFuFkGN+l5i4BCnBrUGrzDxIcrVoCfstMvM
Rfyhm/dzAK8z3Y7SRoECBV+ZVsjk/xejM+PxHdaS8m/Fh/SjxwrLl4eGmDkD
Yc2lzgW1UjUazQ99CUqh6kajHyVF9fmjnC07gHVMwhV9SBRNcgze1Pp3unxn
GNmszqxlS0a7a8zCh9UVGFkCcF5lj915ZfG28KqHsWQYoYBTlv1W32MDsTa7
Eqm8gAE/FMSu4F4w8c9bIWs1BLzUHOqNZgjItkutyqhaPfb3xmNb98iwSftx
Fb4wtRg3Xqvm6kE/REY7mi3BtJ+CSBsIXzSIlzCj+zRFPVd3AnbPGgeW2SA2
6aJWknpUQ1zbXZXNqzS39XYElTlBbVhUWrgZog4mvu/cZP+pFRmS/gH3SWgj
i/xrPiCM2XQ8kNKDn9uA5In75wSnSABZLvSSJawPL/91zUzcX5g21El/3jkb
vvorLLFHy5uJ7+L131iyEMzxJKBj9GRAr98T5Kpynz8Bwmt+BG8AkJtUfX1/
pim0yCH+ivnH/xsj7N8itMRfuYLqvMklA21Gvs+OVWMofZIj9HXhOBP/9vvR
9ykhjjzNyjx4E2BeViT8A3TV/SlybI8vFSlXBMsqf2iAzKHlokTWs3b486hu
537+wPME4dv4zUlYb1VIiQ9I67PmOw6b/IQDyKGGrdVU62PHuDQk1VZSvynq
OHBqJE4owQTZ7Ugl5Hp/SYcv/1zeRUSqBI0AIi603Yu/6CQffyGlCN85obHM
41urAWoeMOR+RsxcFWB8Wo1+vuOjNO4odiUA5z0a1t7A6NYddQ0tIzMNtLw1
Y8IwcCd4qMAX68E7HMDNsaqt5gaygTYkxvrT5OkeB9ZDTrEz/mT44ANDzRqj
Q8loqN4EdF7gfa6r/vxiuYUEsLdAi039Ug7nAMuKNUvBrKXASOl4hvbkMNdM
Ku/kkqPId7aJZdWuTtLh2/5hZ7EPaAJw6MpeoxrV40RO2O1tkygZxNTNHEDX
sdPSj6iXvnlDtHbcTRtM17oTSZow+X21oE2Dt77+UfHJURlkOi0iIcjIfzyo
eeJBmlkUNsgvYtemRw/zCN9uKyymWm5DoOxeJ6BWH3OAGJeCwxm2RmzT4uw9
A2jMQJWyYfN4KtdDgOrDLvJQx9Cv5su4Oj0mZtHik2tdrsWSvD4qDMKy5mKz
LG570bGoimvsOSYwvHH5tPtQdYIAEKyY/zRi9D2G6hznOZ+IBunpNl633K4W
Kqo8v5z4yv7TvXwRAak2x1SP+xd1LrW9TCEqCcPJ2L+U7HQYsuxbNtZ5jr37
wXi7FBl1hMweK1lkyqJIEb8elxv1y+J4zpuEf7QBoPT+MsXjp03t6TFkaJqw
2Dn8FhM3X6HV2Y7DLZDRI8CMQdpE5Qwj5JS+LP3GWkJ/7ynXWohFb5JfvogP
Q8GKnqH0BKMowUFIdNUrA5GZopAZQwj9Feg/ts5AwL0OLpZ8vVJofA7DXLb/
x7IrykpHPghAGQQpTDGJGFhtVNH2Oz2zI0XRyKKFVE7Q/783su81fXedaSsJ
gQ7cMYhqJ4k+eYiztc0WU4j/SXp1h8mU83w39FOzlXuq1Epxph+6k/nTR8y3
NMQWd8zgrs7BnFAzlaiSpw9VtFN5uzEwAzZqtUdTmzeiEaj931z3o8B5LirL
HkFuvBrrkiFROj3lmezxB0BvyY8nNYXi1cBkOdW4iKBqbEHeomyH+8lAOXgx
9uXWgZ3UJCz9cFPh0+J12RbfJXvufXLk/P7H89Aht/tLmPmkBWPBa8B7ax9b
zlu1X5oELHywrSklqPey29XCIJSEJqFe+btIqMzOw41mjD3ENqdrjwdj00S8
vj3pEsLb3FEouceSJbGGQOhx0Wtb+Ndg1vKIdcIUgTYH0cNnbDMDTXflTCEZ
H1hFACwfeYbiuUPT8TtGhla+zfTUKPYpAkgYMWeG+fyrOqHrtmQ38k2NX1vT
m5BJUdoaoqAZg43qIxO6KtjgqOOMPyUuG1aIMBBFqxJvNyGUKYc6URchhmrr
N91nceFk26nZoy8o+Njug80NlsQkPPkspMc/kcUfhPdW5eiyIQCvOXIzAk6g
y/8rcZ0d0zNcq6D9NmksF4Xmf99m4KSQ1nW2NE0zDboTfyrYYvZ84o/1EFLO
8DMfl00haD/bfXm/oiCI9QzmKF50VhYpn4Fs6vr7Qz11jmygAcS1ZPktLXvy
UOphMx1lLanFxvJrL7X8lqphFKmES922iPHmNPWWsZdu312lX587O3ZaLB0v
DNGTF9bg6NwojxGcq+Uh5txrhJLoth/vkdQv3qBxMGwcUS1pOTSoHCc7DDPx
ObsNiTwcGHyqZ8EVimC9hce51U4IdF22n9KJ+IVwlUhB3VueU2cCQIyfgYoV
x3wwNxj3SrSerMKyNgjvzZdMUb/+1CVuyXLl/UJC2jomL3XPsLJy/uDuMER8
H0WMAqU36kcRFItFz2vqnlrkq58USsaGLBbP4XOiL193z6lFUKejp7daspsD
vvmFfq9TMJqpAWHCl986hy4yuKUmFy71zYbmEApCxkEov9LnyPqaL6ygXm05
e2uq+66i9Plie46W9nl5rg11r5Dxjrs3nUkO2nn1MdxGdaZOn73YMiTYUInf
hrNmV7EoeIB0GlGPMrMPsKpvCrMx8PkzynZC4I1sr6uvCQ5cBvm6ok07VKp1
BIcnuc3UKrrixUO3mb1ClfgpvjIFjm7xYX12fAynA/drLt5g77g3wBGH49gW
Th2c1JdAVm9fnqbfPZuOqZyw1NalM+LmErCEXjGQAzUoHOWhaxKeYfGUwnez
I7gZACph7WEs7N2AAFil5hys2b82aMaVSN1PtjxGJGwPH7gTs/tX3xLMxAvV
/IrjckdHKq2/npIGRgMYILIdYAhLvbYYwLM9oE8PIlA0GvKCU3psbTP0b6oH
DThvfw4bjDjklRgwvnojTr7wEBgsnXoH8Q8a24HtYn5xgbhAWQfMVEvs6SZf
Qondpuri44HNLPNeHZDut4Ff5WkgQm1aHjjJ1yJ7UICrBvbLW0AsEHQKeFO4
Hlvk+InVZVp/+5W3HpLjKO3mok/gFTVt0TeKHwUrVEO9SEyGVES2BxZtTwt7
EJCwwsEo4k8ellQKGKs/jIiDwzpwvqQnUX2h5/KskqoHqC8/yhk2pZLBZZMr
keHLvMLhmAvl+H+6oAMqWRTa9bYreC8B5EqOpTzENdEZGZ0l6szRSMNl+kX5
6897HZHJLR+XT1+oeeBYhmr4ryjbJMDzj0kVqnpBeGIkBag65laJtEz8SeDb
nmDwJ0ySe3PdSyo9Y/3ohjTIThbbfEbuNpfd193Y3ABMb80cUsRVOJ0ZOJjs
8CAlE3WfV2fZ0lmG1+n7OpTKIRTCosn/lMG+fbsPGDIBpGODWAdgWtY9SHhe
/pV5EY7PM73tWKh4VazkGfuNJBbOZIiAGu1rzMqTLDYC4JIR6vS9O39beatm
5YqSAb8V8IbBcAK9eAdjD+Uog8lf/3BK3FZrQKhtof1cHxI0KdPwr5bqxJ8u
oVtVoCJQcuPeJJqRyZQFQx1nCuuCpB0ylasuEPIxhIgasFX7uELr4lIaCJwQ
KWNLNRl6bPtYH6swQfnSSsxF/8tUo3BcUhbM2HW3veBcGRGeshC4lWoXkFRD
J2MMXdX0SMEn2cp/u6xc95pSgBrOcaVXUs62C5QeOqilM5u0+hWp30Cxc+ao
hqrDt6SfqoiILQhlq4R3VKGiHIqzOayaJieuQTY1DtDxarTctIzBQSlSXWPg
IOvrQbuHN2OnvUXVDJ24eHOYWDyXEeVDWMr7LzphZ0cKK3p6kQ0UdpKYnf1y
Z0O/kVSu/+x/mF4AdgDi7G5n0I/lVmj3LugcK5ZhZPGukx6jfNSB24ZfgXLl
YELajWPYNsn6/Z385pKmV9UBu2jtj1yONO0rCUz7izhxkqE2IfJYdl3UQAj0
su8p5rnHFbKDN0jSMhHc9WwvYW7bz+qpfXv+9sUnG/na9PuFm1iLMYW7UbRe
9625yi1+4ElZ+8Hl43myoQmFFZmXTmrzmS8iSOxjjFsP0kqwyxAfP4mdwh//
oEVWweP838qYthRsqfoW0gSgbDpqy0tyRL0WAoD5FEmma97Mcs+oOkO07AN7
pvnPI6QezGN++SXQFvghwfRqkgizHJGH4tQRe80zNieZ2xaIbAJzctylEIcB
tE7g4tNkkE6XkNTd5dOYHO5y2f0yIGxJBJnQpclQsPj/uzhHegwUgO2nZ0sS
apGGTXR0K517oFsoXplIsjcq1yIDY4BfaRe+3/69QQc/fT7VYVjrI9IIMwbB
Mx6p1adOMh2wFACKNJHubyb4GgHCDgFZH0rNJYY+u4iP2i5/viB2ZOOCJa2i
yxmsOftY3DvlDYf5D6pr2l0od5TzokRw51uTyQjbBSgu1MTEUCgXaqraIc+H
BKLCK1gXgsgKJ8z3yKiJXb5AQFt68k0TX7F5W517XCLMpwoiUTN3/6MpsguJ
yOzjK9RdLStzkDkGw95xEz7jJ0/YR10DY3TR87VIYWrjzOVOunditZClFvl+
R4pzk6kgFIctHUHjlp3iOruBqjSR0XL8hghWwwCH5aNwy+wJi2VnLsvNdwQr
M9CwzLU+71VYbzpOLvJBL76XTTfuevlUNXaRRnu4kyYvbhMOjO/fSuxdAoYS
/5wdiFCXMV18mHfEYAbtDX1QcsD5P+jLwPUIIW7MqR8w3BZ0lRxbQO2o7o3O
nytIB6CWzmfhloMFVGvjzjaeg4Vfp3XgXvdUtIZMOWiShYktIHu4mfpNN0xE
NNHmBhx8JoppvYz7uqPzz+X9P1XRBI3jnlw+boDpKTDzeKDVLNi6HxHE67tn
2ShnJ1UYO9Htw6SpvmP6288hj/0ZawqNx9H4FWy02Qej7WWkdX1fERTbm104
kDjb5LX236G5LAfjTe7y4qa4fa0G7Tt2VJQe78bOtr4eGdszunq2Skmvq49w
lV07r6mVETHO3sbtl3IJxO0SezOcjuVzaQgiFGX7nX2/qQ5LUVcfafazzO//
IPJk7FL8S7XRBvmaG6qG8fbufiHwFTpxwsSscLVblwWrsEsS/FSP3qH58RYc
YIOmwoByT8MoAwyJSMFTu0tDpohKTWPrh7x8PPnuOq4g/2+LiloB9ZKcnXLr
oCIukh2zk56vSPFOQuUrFY5RTn+j2C1k1FHuJnubNbkgYJE7T5HX08BKax79
PRAb2jD5HYNX71lBdgnEaGUoEk6ZPyBsZamNw7ZqP1NvSo7F3sDKtW8mnMn4
x6cQbQVNL2mAFYpBTOZTtvfYW2ZJ4Xbo/QvQmWBux8SUqePN54jg+QsR0xEf
W4ZjU4kaTDwUx3s/AkevNIj24iI6zYRf+LJMbAONPzq2JaVstqaPx+YY7ZXs
PubWrw3RlQMd28AuM+TbPk61Wac90ytCpnoiX+PPHeRViSTG0SAGpzIA6pJt
6GEGiFYg71ubgPH2RKlAEs+eG0NtAC8UL8DsNgDhQ3cgVaDbbnvBj/KFykbH
y3Nr8nfDXrGzGtGJV5rDISdx90GnV3zrXO+V/lQaaMmX0KCEz9u5RA1wHDQy
lgYhHqBM5RfpiNEETmlppZB0Y+v2gC1Yi9Q9cBIBcEVBicZUGmqrl7VV10cA
zQ+nJSt5ibP6KsB2p0b2Pay22o9jLhgag09Z8uYdlhyCqv+c1x/fHLrmsfQq
aPX37bmvblxjf5Yng6xz+jVO5j3MjB6ve98LVXyec2UR4o8jfEALL25OjrKT
zsnnUxrw4Zn+WHHRZHqBBL8gs0Si9kYhcCkgpTW4dBOv/vBmk+0lk0ZeDX/o
aCCxlVDmnsqZYA8KH6Khcvs2/wHZyWKGzy/k//6vuEpCfRGpSlZJNryGjm9z
RsgSyTKwP147XuyijjsWy3jNK4Q0OvSo+9n3xP9t7Srf4wZ3fLf2e94r7BQ9
84MvGSRyo8oBJP7sQpM2v669qj/Bj5odtN0jNGVOURTi2PU4uAUfZ1KSRMew
/EkWnZacOQrdF91OUnszdAivoxieC5pWloNpjiHCqmMGrThGJDz+cH9Xmjez
tqhHNtmKlYofOSfsUfmgeGY8s+uQ7Z2Ew5b7ncOYne2uRIZ8eUXI+ZbNSTIs
o2zAGCp3BKm5AAdfn9UEPfFulYW9BsJgbVOU7XL9V/jWMaZplwuLFZwAt5qF
zVh2QMgAAaOwjgeZz/fuIRrnMDtgJtYCYkbyUpySSRpLhmgBmLiBDmnJ71pc
38nMdAumqfS7Oaig+zvjjbb2phAWzXIpN+cw7CmtDMQrxMF1LIW4nAMZz8dk
J8XevdXN3BW8C51tZZcNllPy+q+/kXLCfG8GTJyt/exERJzZ0P6q8onzW+8r
qhhHmoYjtPiLHb0MZIVukUWAHnRTNrq8cCiDW31fB53O71PN9CM3Fqv+xaQm
Zmj11POywJoo1HgI8axnvKvj8e+75lARGPWzDTvOFvjqNSUqq0PYWtbuE1AG
1D23JOhxeRJuvrSQ8b3IxWjN613D6Q1+e7Fsl9K+ltPETfHYH60qDyase4Xo
8vbbec/6Owgv2r0HwQtOc6/Kn2Sk9d8GDaFnjVGMjUzegpyOuVztTj96ZjLR
EOqJYz0mW4kOg9RqjlcoK66TbsVvpEenqA3G5CjGbRMfx41gZcNypa1DALSq
lycC3gLyQF3cBP68KgZ6+S6MwygraAW74jB2AQhKzt2Zayj1yGX/xrLDdIn9
axuXRynPeR4i7vIyEKQ/VeItI8WOmqPWM1hjay7lekA20GNEOr9WnfgVxWZx
pz7SDyzLA1VyBUAI0Pr1FGpLx8kmWDIdbnCoomvtaG4BMGXBjJy8SUQre83U
FkWU8MyASLZ29F2N76QhJolc/R+kj9Apb7sA9o6bxWpbDJ7ADJSXQURC04Ud
y8nuYKyrIx1m+t6kl7kv697jEBI2llrpSzndlmnB22cxo3rf6BQV9KBzSrxk
qrLcj1uRfSvH5udcwPPbngxBH15Tu1C/w1i/VOvCDnhoDYlgjWnxfrhuco+3
eePcnps4ou+vGwHdmoCVaUwWyA4SXP9+eN9YeqYpQD9KlQmtzyN3MigoQtKA
jsWy6e7fv/08PgAX4434zREi0k6qEcYdYODRdipKY+j4J10UdhjvMNZFp1Sa
fG6RqQgEGdVaTi4P+ZLFM5+Jar+AED/3tj+k3mKlBvoEZ+8S17cBpcldVHGj
+dKLqa8IiVUQUYIIfj6WLJVa+sxwkgJXAi2AnqqLXX8EprNeLUZNrN1jKbCF
eGwtX7Boj4mbfzBTBA69s3gbWgxjHq4dUmUKGIOl8FtmDvN+BS4dFs46mmwy
u1MhzorodBWbjDtcAWGnjn9vEmoV82bAsWAZe/lF4agJxd46JbtUqKMsPC53
+MUyPdhdoPoZc6InN/xFn9DfVoH7jNaKE1LuQrFWOHHLnvyI6J3FVAnnw8m4
u5u5OQdAqHoGHA8uPPnda1OTLHpJ1iTpH076jRCU0MkExlCrBUKatf+iHVuF
84m5fELh6LBQrsNFjkNNGfeI9MVOn0tVq1j9HIxIaxF0WBdlwJtt6oB9njPl
UlVXpDGpGDT3nFu1VyZnT0qXnL5zNhGPQFKVEas/vXvvHq9hlViXZWt56WlM
LvdRQGNG3xCqiAnRe15Oqmr/9c57Yg+u4q3r8cVdvuXcJhc9NcV2507H7xpF
3frPlCqLkzSoSKFl+k5Q+qBMVgEyj1jni4tqXdeEyKK0aZp3aNLp/K0c2mf3
6jgSkkB5tOzEOKIV3PGOqcZxN2ARqVE7HbgbnkoRDrILiQcxumf0RxlwfWGv
2jnLOic+NtwTOWKQueNiuAHuVDPn/GJWDnuI+qzvWqyyRJk+Rjmem0u0bbVv
ME8l945iGr+1YzvR3eVFs2fTLTzyalHaSBVGmndmbJpNRkB5bAioBsuHJSsV
vKQZZyvgR5liR1HmjlWcgTiZ9m9CSHg53FLYaS9MBJav4yMim//xaYG8/vUc
hDp3NwNSJy97Wke5bj3N7QnhFjlcj+ccDs6O7zsGteTb863BRaO4tCQM+JiS
a7Gjt02LKF7BT3HWvwN5gTs9l5JfmJRazo1tXutoCDjD785YxPOlpXCpDdif
uTZr+MadYIq6R8S91ca7sZIOglVpZpy8Y7FBv+azvfIfzNoz7skWOEcc4djK
HTbvTWfcvQyGevOPbG9OV7ibsc0Nm7hJd4oSNR464bPF98ljDVBUHuvN9PJW
fi8oqZ8xUIUaIyWuhUGpFZrLBZScWJE7kjcncRe2iFWxH2xgwXIiFgcucMVz
uXg2q5ZzC5f6naMgRvAl9CTy28ycErNI8zMZTJht3wSdbxYFPCw4MVaiuV6f
DvsWUKQGR7uYq/jhIJGDIx1jGjNFw+4hPTQ9MjTgfbKGJ4fFRE9DnNKf9GPT
TaExYXlyhNasTXIVBwugAJC973CnJg0R4Yq5F5t5O4RiCsjgaVee4QloJ3wi
nP3LbWT2N7ZEPAsxXFI9+GVO1RypuX6hamIFDOfyBZd8lWQDaWlUigUFj3YV
qMUjcy8bN5vPs44cZ8M7tFrBvgTDQ3P+b13XpLi3yug7gBUQAYtUf2DZ9XC2
/QsxNwwCSsZ8mn56i8n5MhNUD6Aw3QBJW/D3YKVapo/PCx93aauS2/wjbaO+
M7zBOnApLZqERaMpLR2mE8037O6Ny+lNoVJcVYO+3oH8+scMUoJjTA5WDxx7
UN+eUG6XgIrksbDuYiYuXvjGySGblRwS0+/gD5Y77m1QScVeioXPCwiyWuSj
Z7MIbAdrVj7MBnraAXn8SX2xw5dbIxbpcCOHPmL1t38OODFNnCXzXEeczWfn
TjFj2FtJ8k9in51LR1ZxAZKlSfls73oRrMEHgV8K/RdyfJOUF7NisntKDkEH
C8Ee6/a6iEUgctig2cklYuL65SVvQE3f9iIrkVrCGe/AhdtuV22LKNTONn/d
l3K/DqAU4nti7RF+l5mocweKMEJ1DIlF+qo2d5kQIWw6cbkoqTlKwcgVc4/9
YFjQP9/mUaotRE9IJRS8pO0sE5Vkejo41ZWOSzTMikDO3DlxEg4w5gbCDAn3
L1JqSoY5dSlNaQRstDzdyRtyTScdjXG2prsOtHJub4mcRYCYOcqZWsyWdIE8
B35MzwuU9AAP4M3TBssk8LaCkMfUFF1yauNmDlsOr2P2sR/TP/w11vSu+vQL
UFg+FRhBLCCglQ5gqEHuiDAQVCa/R28C4WeepMFaP0/j3K9hVhgwuwPE36Y3
9YCFedfojgD4CUtmu08hDsgnsyWPJ7NFglSVYhJtUzAnApIgg3UQLoOTWgVd
boCMpZSd6qBiKzwididjG58WHoK13hPOkv656pOqhb/qiinb3JPJITFRHuPJ
I9yADrzVVjHmJlYE3LeIqieMWrt4KfSISAYmg5qo/lV9UpzatZhXaY7E5lGR
lcgRkZged2El0q31WoF7I1VwnGteb4WbPWgbVFajrSxq5VqEbfsEwd+87UeX
lhgG+UxIiJ6vVJriIcP+Lc+Ty9o/MHcS5jQ72JzLfy9/avFTINfjFRXIg7Ny
KnV4g3NEZMRMy7Os+2un4qVVvWlP6XPF0j4ypkWTnvO6w+o1H9UZq92x0HYs
8YGSQiHilME2rsn0FX+iHIP9FUlIZYtUtMXve/AW/f4TOpKBx1tyCA8g2hFH
w9z4V0EL/Nyek/PcF9NCnq257O+PPi1FD7pFinRM53mDfLvTwX0AEb5Vc16O
InCtEuy0ggxaunoJAaTm7eFobEYmhOKO25E/V0itsGLlXsfOhhiBkEb9i346
4NTXclO1rcK5w35bAgdaxoCrDTENQMPf+9282h6kckM5Z0oUQpG5Cc6B1OB9
n5EUET0Qqxf93TvkZQ4wXYq519o7rRanV5AQutGQz5kubeUX9e+e074zz7IQ
Nk25jVl+XWQQXgfN144MZW63PvkuM7Z6PhieeoDuZyNcRMEOjiPezyi3rE0v
ucG4tde4m9s3NqWQN2EDz8rlkbg4VyHwNixLbRw8zd/ddCYdxENwK1iw+Kr5
Zjgsuhp7Y9KfA3zxErFSK5BMl855ik5b4GquGW+BOH5YLrXqnUzgRipkkC/9
OiwuVe2qRZ2MCnHpHyqRy2dBB60V1+cf6Qwp20LzXIJKmnHRYIazd4WZWJIc
2oLiMdTKH+4jxNdotLIvZ4SewNnW5JLCuOthIXIhQWFHmDxYMOAjziTg17B9
r9P12hVrSt21bYkmKH2IMhOLpGSyYiRn6J7J1JL40Dc/x2VCSIrwX6btEXXN
jbHtCqGRfkn59fck1DciECFkljdafm5vqL1yvKHgme6YLvQ8thzNSsTVkD+8
OdBvJLEQ4bruQYktgfrklPEPBAMerzXlS5pLAjX2DtGVDnhlNg1uqFTRtV+I
uidfUKGnTxZwuprxVxRaImTj1lXd6e3sUmZV9Wgjtmhy9GfLZriPP0HqiGRX
v2xuWBjLnHYCAbE2L0vhi4CtLRvUt7sraX0Jbpah3YoYXAFeePYbaiK+vgje
MnCHutQewKIOBVOCyPtXm3CVmWkN6Pun/x3cGVUYb+v0Pe7PEoMLxN816Cl6
DlnZ/esPWAKeFHmBV90euBEwal7qUizTKJKoH7pM3Ve8T61vMeoftefrzcFh
pxOlJJC4n+/AoIZ4uH3oLjkCGc75qPe/VeiOAvyiga9Y3JjUMsZeYijCTr8q
H4Zq5pDx+c37BPLeEbpJ+rFnCLnzr7sZ83D3pLDZzwDdZlnnkp54Q3PgL/++
CJZamAB1HZhNEd/wKkgxcdmXhmNV6YxqSuJMQaQGoPCA9vC90Hk9qXrjdwGD
6F4bHvFMp3hT05AhnHtA2jryTmY3Pfz46/E9vyl5oJZZ4sdJv159HyR2Rys1
iR4qNk44H6epu5C/KmqjqYQndYWb2ThC81rGzZWNZXBXSBuiudvXmTxGEGDI
qOhZScNCG9Lo3P5+sMbWeiVUjbz33AkeXcuE3ZEf+yADsNwPIYuOJO7J15vk
JuKyz7z4LMj13St6C4dj066K+ZRaW8pHDyDxz9rx2tHh4vAKpE30c7jQaGi+
gXx/2dkXnAiXvcbwapIxQFTuVCix9Ve+I3x7ayykLHf6HYnrWdOdF4lx2dLT
fRGjfD7ha/3DlYYwicwvHVsdizgRX/S7q3HMKYJeHCvYWMMWgJw6AY6aiT/R
IkEs5Egl1YM005zVFhp+oxZnosRbeBJofTmnwYJweU8fhMAylvRXAsncJH52
cypQgcLpzoMpADMz+IJtcd9ZLAKgswDDXmwNeKiC5wWyH4fHZQLdpTwCm1Ip
8yYqSqUEwdxzulHM1vf+EawgjDDe2eDYYcmDBXUA0vnoSksewARSjpkzgVUg
aqWgYyhIdtV1yNhYzYwChX/TenifKQSQeU36mTYa/QsYLQTgDOcmDFgGV4cZ
BHHqEgv6+LsJWpwNjpgOyLClDJy9B/J5NuEERNtkv0wQHJ1DpySBm2+AbZES
OGOxA8++RaRrJu6iHKtvXMbyP0FhMAl8vWlDpluuGxUNyGNaGQqUlBGjXjlk
AU85PeKyWe1cHcybA7CMg8dWk47cM9GsqUkaxMYpjGZhe07VNd5Ci/jAZIGI
Ajskn7hZfAt1kHWf2lxm2XrYj6bVLnntpSL7ssDtItFN0PDKGg865KUZrJdv
gruN8R9H+8bOtE8CGvcKhvxmKrpOUdxKSoIQ3pEHJodoOaY04uScACN65Ngr
ktTSS36cDNqbTV6VArRUV/sB8/Kp0wPpkaM/nvV2gt6hx4ro2cIgSB768+KW
2m7eXfD2zop/OHM1itCD32aS96rWv0zWlG8pj1k09XBHck6wfkNdqTPDkRQV
daVzLd3JKGm3kM8h/3Eh+lRal5ND4eW9++M1BKM69NIXRHQblOg579kA7bN2
Ip4/+mE1U5GgcQEC/7r4IMv0cdJq/a4e1iDfbFDYAPfHQ5ITnxNQU5dZRILQ
ZvuZT41K9ylRZUqKGCgf6u97Y4A4gpqlEZMcECy/F9zRRKNETHVVOzmzs+4B
8f2SY+8/LbJkQjXBvc/VQ4McI86nCpPPcLILRWdqi/iv9UI/X+5FQv2LKTPh
v9xjmx83oNkvGj86mS2SrINnb7V5eOQUHwb5ysYnKGMDUQ6fVZ52LogcrPdO
T+pvBHE8+8a6FrKcEF44ZQcv0WYEGmMmALoxCtMLaxYxWZnEngQ5tJVbLL/2
xGkjSVszjojRpticIg3duvIulBABDwSHPud7127obCJFVD34yNpXUwrOGCqD
hgFTVr7gfS7h9U/AtwKcjbMoj4LdDjPV5gy3xC7eIk1bmLxdKe4YcaEscibb
0UQlC0bY1xRHpVociJx2qH/oaDl6rlOptyHdE17Y0mUTEMmw8uQusaQ79Mj8
ld0FNa8sWcQ8QaGxv4GK7pcQfIJyQDJH/XtsYVhy/Uhiu+Tlz10DR5zzYFXN
Al24EIEB92GPx5bioipf2XDg5hsTj5mWaULNRF1/kJ8huymoezvCQpUqdyqH
Xfj5ekRGAhjhzlTSlEQrmjBlFgn2SeIH6Gj7I7yJq9/tV3nYzoN5kXWQPaCn
rzhPFRGQO8dNGslb1O6U0f2l1yWdfKS9j5iOLxYXyJBBeOm4OYhfa6veIZJG
sA88eXxRNVYEZREzLrR7vk6ZasSoCTajBX6JJ1e9y7NPrSyQc06GzrtHaIW+
nZQDl2AKDWdo19iqevN0iEQ5wFQM0KMB4I0IKRm8bi67ZfIKvqUXslfs2pdJ
0PKDLbl41QgrwOdLKZFE0dmianGkKTQ2IAFgW3I6z6WwNlrmZoDo2+ig8LAA
JgGu9JBxsQXwHcRx2lL7536DT5og8gmn5n6+4ma527PT5DXoZMoEGS8WLsfF
VMyFCiDM46gAXq7yOsx+MoWmz/pOA7tayZ4f9pVP639jn2BupA327Yu7mbkC
zGLolaoF1sX2jEoBhcEJw9+g5giD9FLK54PNJzBsZlpqBk9Ag+LhnkcUjj7j
DruP+84hFDVg2Xub2HpXr6QnRuUVOcIRg2RZ9t0xc77olAapcWyPkaXxJ1xE
etmOMD3Lc//fvxUfF5CRnmnlltog7Bapspkm7oJGVkudOojMpXy6ncbXbT4x
r75BV2sz3e0yx8wLiliEphqvAEOJPIJdYESKKtov6A2oZVbGkabSyclUUx0e
XQ4bPhn3KRHC2IKIbUlWCmAq9sSezFmhFI57hGC6gx4S6qVEA/HJ3m0Ie5ZY
s9iF6mSWCNu8MsByn/MMT1M9R7sua8wD4T4wHxEwN2x625REchXHaFId6RkM
AhVao4ni5SHGmM5TtpJr/OoQLXGLWBdkVavYy6WXknlIZ5j+8h1ltNVbnLTI
QAOidIP7ahD/8eoMFmkpHyzJWQu4WZFcVqh2yciDgIQBAPiq5Uf4xwhHsABl
zH9gl7x7gDZUb1PunFZ7SKYvR8qiCEMGScVGbIQJXC43BgvnY0tWEzU67lBw
WFcgwQW8bdyqe4jug7F+W9kdA+KOUg+S5TUlIyIKZtfefjFf2Qttp32F6Uag
UxF+p7GnPEaUuApUlOztsedQ86h8TmIkgrgJxlfg14F8CfdRr8p+chyYRzNf
2+f5o3fObZ0AB8C6XGohoBXwN4ZejCLo38mZ2vCS9y59QmwSb1gWwc/o+RoK
WDIvGDIvH1VyJ64cIsXjKrErrvxejJFvRez2ObBr1y5G/rD4uyFpglUHz5n2
6EqyStOOQya2pku0qwKLSudWJqlTBXz/QvugrYsoCMMpz5IzAR9UaERN/UuQ
WK7TE2zWtoAEp7/Mldu+tzRWhJcafhoI9nribz3vWLoZnuVPbk5nu1gzN5pn
xZZAw3LLgmQqiHJTaLfPo+KHL2bIi5V+alKRe4lFiNfZdGPtZDhY5j/3t1bj
w8Z7rgzRf2mueXxHMXBDSio7R0b9HVCgIjncQ4fstHYJh0XcoMAa0ZF2m6Jt
hXhEBNbrqKm4On4edhAZqlKpByZtzKMAVVtM5PhzgBp+4zQuEZ1tAtInHpRw
8OiFsy0AmNI6pix5TFjdbj9BMaBA5QeUSCwVdB3FN6wpc+yxwBIcUDwxQ8QL
0SzEjDzLXXXhNwm39NODHCecAsMCi+UI4iMBA7cfOGL+jYaMK70TE9E+kkiZ
frSooUhm2CpZc9Lz6lvgWPp905yJPEnxeJzRX6rLVxTO9457AbgdDmjMCax7
5jCNPzzNJg6P4JP4vGBLNwJHpmF2IzTuloyF8r2AeHpBsrV6YhnKs9HLIC53
zwGk4x0Ld8RLHhukxuqdWFA9+jU988oxxa8UTVb9AYC44GTrYlw3A+WyqjDh
I9nMRZPxvDeZY4nWS0SLA7V1FR1LK6uR4XyYeoO4cquCJ6crj9zBaOzXmQMd
joEiFP9m2fJ2fF6hc5HC/N7/wGyGCZSwhrjaYvv/T//sTEsX/gnseh76eQqp
Fae00hwyb005rRWRtzXV9bn2FWnQL82yKRam2EmNeeZnxq3JAf5oW3x0H1lg
F4mPqG2B3xmELaGG+X+yPBbV8EBqSvUvyg4Hmkj2d4WdiBcCtBl1xGmYxVEl
EidicLoxO3E6bxX7pNYmjCP1bNj8yt4Ha3G7uFmjzmemtthLu6TpuN4NxNnp
1hi493fX0njF8uZHQOoBe7z2yuEBU6USmr0eonmJqpOMF717tjVgAFmPGa1b
VTjOnepHbaV1I1KIOr9rt3c5CdaDNP6g2ZlEe2jNH05QO5d+cKAX7oD2iDyP
cZVr4lymRkqKS0/AhE08LIpE+gafxzFT9+JTyvJNztnCWdogTn2H3BdYNA6y
8r8wDcONi9zWbI3wfA5uqLIrKODqePOm0K0XogCJ70p+JwKQIurj4qnvnd7c
PBc1xC6raaibeRTYXxJ3q2BPV2QnhaxPv8KT6kXb2P/USRCS9pFtgz/vYdL3
olR5ToaDCuqhJYbiCCkqQNUo6V9FhTImN9yXbjRrxJrsJQo1KgrgvKVzHu8y
g+ZxWd4hLeJGoXu17uJ8djOrMggOSPlqMLornzp6zeSOP+PgW25zqF/aoMAm
/l/lrzY+QTB2TudRUyb+leOO1NeGNgwqnPXXZps+M5by/877nynwtbcvFA5x
bnz/p6MDIRvLXXIeqC2GGp5nZVb3+fz315qQJaI732j9kmmhY0npxkdInd1d
5LGhlyUQwPxTQtS4UrRGBuvUXVPd3rVHYz/aHE7X8HUyBCuUO/ek1pCep55R
8INybwIcg2kLSlsujNamdFXBRsCTq7XbdLqKKIUD6pgosZeACBomfac5hyx1
9vaPNBx3HfRUrcZ7VaAYclQqJ0N9L4bzR+Ts7Li4q6j+ImEwtt7JJcWrFHIG
WY28Lep45XVwlMBgjcV3y2Q84lHv1BGbE8rMvl+CRDHPnJtbEMxFSLooFZrP
R7SU1VNpy1lRnVKNT07d7BxwwzR7ugGNVaTShCCf+8gE3wSYROzSrPhIg6JA
tG+F8CVMUblnhN6ZwNpHbg8akiGOREO/uopaK01KR81Hdj98HdoUrhV6I1r0
qyeXRWJxfY/JJ3Fi2ArTufzkNsRUi2ym1oJ+0WHrgE513H6/NrvKWEQJjaRG
Igk9lPA5DGJan2nWls6a5//pgoKs5bZZSuVGi7eGUb6ZcqW+ul3pFqqDzLVF
oD717svuTWfUqjmveKTHhgz6n6j4Lhqo/O2h2oF1OCC3oWAgamR1lbkYqgF4
fEe8ROdGxy7IOVoTUUAUaky5T26excKtBRYWjgNxpO/mQuFoEkylX4zdtY72
n+73F/l+5ScmK9mrqtYW6a1EjmxX9tc/g21b+lFTk6by43IGyjEBHWN3MSCd
fCwR9lRheFeWiX7kRjlADL9qefGLCwkqi+GOkFMtQU4Es3tSgSgT0PEDRAb7
aVhBvilnUueHVuG9i/EABJykYQFXL4dfs+SNwpKiMewKtwYdDfyyQrNIXBFf
FQT66MZ4pCJFC1qrCDVGy8CgQWGcXojCKjoHiA8EhY6Y8W8syNLbZdby/IrM
oCM+JAGMMl4AR8ddGq+m7tOpgRkhcFmfUzJxAOPBWTR4/YlKxEJ+ahwmTzRY
j+4WwOfetn4DkiLfUzHceQrAWzAtEFhgI8u2FdZUl1fw0Wgy7gFofvmmfLWC
KDdt/qiGsq7PSFs80wc6ulchuM4LHK55ntV+6x1gSdmLs+N4nEtt/miVuEy0
ICo38v0YayuZ49BmKISMIvYoU4Hzkmaotd/1iiTW+mb3QKKCHGsfWJoHGxtc
zf96j/uF05FiDDBao8NyO44j3ZL43CKN/qaE/1xBZSQHMXerOBEcFG1cRuKb
Kj9fUx4vxEDn7QKSFMtb+t5IrfJiYHzRt5UocRNMdcmnJ783hpfUFz0bigBe
iBRw5E4z3uLjOGTWpm0tU0UExMMpMYGgFOPRCCR7tE3Rbd4hsBd1iKnlLWMv
ypzYZM9G8SkeZ9xACeK16bAPonwS8K1q3wUVaVH/mRAEOlmGl/7YjOEABIdL
wkOQ6kdqQX50R3o1KeKCavz/AcuGuvgpXsXiHiMtqd2YpkzqTqRpQtFEG3j4
EFz1Wbmky1EKOdwcOi5nvWsBMTw+ulZB9Knv1GVwwlhuZYKiiNHYnsU7HkoU
8DCGaLLUBSEbJw4APC7ztMlQTrMtC7fzbxCPu9C62wJS+/kCc00eRBaXtgoM
Lnfgkb/KjFMzPDVPMfV1lvL3mE/p+CcCxT+rB7d2H37luOaCL9UzlKmx6GO1
6HTadF3TphMOX7fkGCXD2VX9PaL3nchbe8nqFkfkNXAdrkxAHO1/vqeCmo60
0bhHNIchYK4+kA38gKe9YATUEyHuMQIiycfWJYov7gw9OZZnMH543tHdqdDL
lDSS3ENrrTjRrkOElAGNLd50xXSnODMq0/rNBnDZEjlGlEwfa+17Ais9WQYy
ze4r5ry4GuzFYYfJK2shfF/lZWF6yZDJKEwwTsU1gJu5UQ+l4NK9mbL9SfeE
Hqb4sLdVtkiyyOZJTv6A+kwXLg1nZdGHX0JTcN4J8ffUtESsSjDeoYJ8bMHR
Tw6kUFx4tNj5chGpQBdcRLt7/3gU2GY50CLuQRSnzu7swwd5p0zZCcosLkUp
3CPQFwtF3c1vmnk2qHYOJr36NmSY0GeFBfK8HwQbOD3MLs7ckja9D1lGV+Yq
fChwpehC9Ew59Waw+QapRZPkeGSiSDDLHuq/0Oj43J2DcsAeFQHCF1jLFaAr
0k9JgqCprDEd50ISJ+Yoqgt88Jx4xfWbSeO0WIEGcXZgHiIQdcs7hQa68M67
OZ099xHsjSc2Dsl38yILYvrgQ0Vm1fKiOU4bHzWMMmO2kMkn9TZUW6GVUdOJ
klwBdGsf36r+p6eK7B4Pw6he41u37eIZP88kMpYORJOwn3xeTFCQhKV2fvDF
iz2//F9jNt4jpOfPt9iBawTJOwIuBk6CcBow54Jopoi7nYxAK/16jU3r/AcU
h7LqTSwxrp7joZFNWijXDH77qt8bgs45ZNMVycqhFi1i5ftiVBa/lSUkGOOa
8VJuXnII0WHIDb+p4REQlsNKduAwM6jPrQKixXVW4HgWLCjl/lTSyvlUqTFd
vrzpyvvgJVr90+/SmySlC3dXvtbYIAbqKxN5UCFfmOHOI0MyWw8qRHJI8ymg
y9gxMhmHbb4QTVBvh9I01OMWF3TOviurmD6fZiNISOgLh1IVA7lN+AYX4oW2
ha8UMLUG83yNlG7SPdV5PRCQHpt0/9EWbCkRVfR4AasF8xw+CD/y3htwO+VB
L/H7JLAfH0yHzgd49TThnofd8EwyFWWKobnQRpzoVlKnW/Nx/Hc6usp3DPTj
lhKSK44Qbm2kA4Qe3C+5wv2tlMd91dWdDisSWVB2/qwOSWR1LtIPQmMU5uYj
v8x7TsqeTV90Vm5mKIJzOjegI0YvWozpsWRx8Y9hsGxJikuFaqvjDPlgJUb0
Qy/v+FWE708Lurn1p1pIdsKvPV8P8puAsugRjI27o1uqb/UijrhIPktE1P6S
fiY6iwj60GLPe97sRCdkwZgzp8n53QZ6O+jMtpALthkm77gAZMBHonxomOPz
pn/DelHxGcP+aCdS1MwkK4ypjRyvtIh6TiONXDAxltLbojONb+dHdBi0etqB
icmO8nIx1/UZPS/tH7s6hYF4s1XpIPHGhFVkaQ1pZRm4wlKCsCzIrXeEQ6TQ
5wYr65FvvDM7EZizCuIElsGMHWBwpf0OZo79zVk1/YqtJRRrg3ch5QNHaISs
d/FfE2JcXHOHOYd1UlMwhN7CjQcB2uZPDm6mudTeu1XYWUr2WIfM0tiyJtGR
xrYf7DpNOpJO/JyIR8ihcZYrGfmcmqXI0Pl7LF8yKCIGB4rkKLhQk6jK+nsB
uTQkitmh0Giduw45K2pNlc/QIRy9t/MIAvq7W3t7MGWiMPRcIVn70LG3UpVe
Y/edh2LhTgV9EVDuJZF2uNNfmgX1Kg9v/soItHSzPcbYt4XZN53pdxviaD/e
HZ0SWonWeYEW8HKDWJrKzIVhiLLCDl0qLr/+2HC6MDqFayFT5yaJxUsql4pQ
rnTa7jZqL7yRbUzD6bDA2mkrciUZ+40EeTqc6VO0VRhy6gJvW5taM7QkAaAL
0s/mVkqc4cmbQPzu25iFmndfBp8d0/JmSb4uaYOqzWRjx3jmhStoFQ1FaSAL
eWbpRzU0aqpWney9qkMT7Rwg8s6qsYWRBfoEMCuDm3TTQq0AvzfMsLZCm+FQ
MH/2En+ob5BDSpAg1qunfPswlvL1dJoJJErEwYAKmkvYitwYmjvG58g4zsU7
1LkTxr+o5FCSYyn1YnX695UN/bwgqm/1TAD1SNniYR8NzBpcke+VBPhZS7hd
uJaEUbQqeNyTO5VCm6yiTvNtGrLWvHhentaSBR0dOFQbaxH13Sd7UCffNyAm
lLSXvCd3hivo3vhIcP/I4deNqYuwepqCuRj7yDIlkRRS6Ix7S1Nbicuqc/o0
LD7oEeQcq3s3hs0tzywzwV82BjStmRUbLsi3cOUgHKLwbBrR430MOjZR02yJ
GwZfEtV3d6y2892Aw2mzRDtMlXekdFHE6GereexfLejGr06+a/zIvPNipu+h
HmrRb6y/5Bu/YBakSRX9A/9ArAUAec8wAupO0d0LLVkzvb56GbFEntY1YQUp
2/ouAoe1zJme8NAX56QQuZSEqp2VaQ7FMEVB3r19Wcr0JtxkTnlKegEEGrwW
alQXbBfl8nBaomU6WEIoP3R6rdfja7wonB4X1X+xzs5R/3CIOzzHi8PTfY1N
YpyPri5XcRKclN2C0UDTuElaZW+Z5/wH9SZaLbdNbkgVu8h43xdXwomgN9m2
Vb4b3Ef+i6VXRMbiHihTXxq978daKbWRnxi+EEfLZBzTHdCWeQMHPX2eUIy7
hn6oBjcOQvMDCUXRbOl7H2+8IaMY2F2c/p+vkFfIXyKU9rcfLVXhL+IbmMvz
oPbWybxyPT2C2zxze+RiW8ABdktKEBYu6kq2sl3RZXj0MWIl+HGXeL5rd0+1
7TIp7gNSZOPm0PjskVv4u0Gu9W8XKGRd6fezrgrk3Ud3h9kUA/7D8zujtZqP
bxQig7zKX8Dy7PA0ShVZXFRe/vl+ZVD0LUCgTPjKz8a7uuFUL5Npogk0cw4A
TzeIdrtMLXEUQQO/7Jj6Xqt46/0nQwgXGz0BVnOaniq6cFK9oUYnAuysHXnk
bVlEu5x8ZVwihd/uoyGt89IXvLNrreZLM/2zPAbxnDrL/bHirBhfi8doEk+R
v7VsR0vIg/2vH6NkiNz6LKIA5GKmjTEINilq9Pe4gL/xOANqH0QnbAHPjk9z
8T9+WyvMsqgoDyCuAyU44E1FnJ4nohi620nVjC8l22nyIPt3nFPGHc2q7IsQ
VGKSsn49dOM85bmomNSaqJyxCtXFxRt1DF2mn97ZScsbq5uiTWtBwNSSoUdo
mei14aZTgIyaCk26Nkkt8iMPkRCJtdJxxnTbNbie9e16jb6Me2dxuyxvGWOo
08ansOGoYZWegOb/Jc6Ubj+j70w7Re4OWfOX7qAEnKo6IESCks+O6G/m7ZIm
MazHPZqocpZ4YI1/p70k5R3dzqdNGB1CjV9/rozktBGIwLn4le1m3pAxv/yC
Y72hTLF7FDvaQ+h3HrD6XSlDSjrzkGzQtughjQTwoVuIRxopyZSO/tomQkv3
Wu265YnzaNz+tG+6y66BHwB07smezx2pvSX3vI4OIa16RolgS7LLLzSfxown
DilrfN/+WrmJYHdkMOA4gzaoW5bUkgsZydmDElS5tIPuAtxETuk3mDfqiBBD
N6kH8hDvpEZ36jXhU4ftysu1cWh+CuWGOhgveIpQoTEFcVXaEuLxCIEd1Kw3
HxgW2CWFbgB/UCP1O5n56noX9XJMbTLJls1aAsk1FsGqmkhrO8JRN7ZMCcPG
xIz5AlhN/X/qu14Dc/x6kN39y2GD+WS/++uKfe0gPsP0mIT+qtdGTF0sABWm
8RNAYf44o5SMdamjGy6Sf608WI1con+K37CpbkZuVJ3DZDH1iefhcW5B8gcE
vWnkUKLb8z15/RsoJ91oAbYEHizwt/3wXpYNLbGH6cjyqmFwojruz9Zqmblz
LmOtMFlBV6zCEjFX3P4Om6lDaLokafEAGGEI0NT45yfbp4mRfKhZ9jicS7Ol
cbYqakSVvHis1/oS/C4p5NTOW0P2oC+9cDl8hvfBNANBqHPVG9v6GyjSR/ty
6yuG7LFytv8ONYMqPMQgME7yatG+bs+jnPzJQ4qYUZzBUrV17a35/ta8znqj
Zgh+GTm6QHVnN9Qn0Q3OaJE1rmFZsXPGibxHE542Nt0d8LEfn2m+FOx3K3PP
hEE2V+7L6402CKuBZLSrIwsjusBIn0ZxMndGccDkgDp1i9dCX4DKZwUC2RLE
9ualESr10cRyzEQWyuPD1lAynzbeyQRQyi6L8gUbeY+OCAt5z4PlxBgz9Wv5
W7Tly9JHAHJkzdKNE7pHBoQZoW638pO8KSPsjueUx5B0YpLTs2Oq+Paq2E8k
i6qr50KqLlgKLqmdDZ8xHET524FOZ4nhQnk9Tz8yJuGEiBl6lWo98MdjAlmj
eRjmVwse+B42a0YXlqvXGikJEsvKNzT/Mw4brLrxK8shbBPoWqzSgHtvy6Px
1OHgjD7KaqqOYwcKKslYdfTJ1Q61ocfR0sEA2/lTIsPagHIBBNyrv/Cuq25X
5jqPLBkOdJPz+4+Hku/gH4/CTgRX0ID5T3YfQuI/amZeuC/iIpi/DYQ+eYbR
I1LYSRMS5qt+eRaX2P2QviDy73Z07O4rdqZl9OsBmbd5kipPJdR1ID/GiQLJ
Wpdxoyi2V4kSDSWqgnhVhspgwrEFPYQRknD2IUfFAF0qLAtXry9fK2KZc79S
ezwQ1Zfr/o0edCcI7KBRI8kmMZLxVg0sBMMb+oMwwXIOtOJGrDAqEyNNZPaq
GQPddfihGiYA1EEqmaM5ng5yEFEoVr06S5z4Vacc5K8rfRFAtNGorq7nIl5G
xzP0dcXMsS7oxif7eJV85pFXXgNYeoQmdr9UYmEzlkJ7Qw2ah5EqCzGZXyR0
pJiBC0JuqPhpyewWcGpoIOU78v+mOc9lQGzdp9R7lxnBhGtGWr+gv95UGP5v
/CXYo+LTSi8WhXhVqwIhDdmd0e3B8StcyvDQMR9bHZk3sJC36Wjth5X/gtzg
g9xfvEp8F4X2Kjqu2mFPisSunOi2DMkQM+YyJ/42f9qDwsnWobibtI1wOUue
En3Lk134RU/HfaCgcOzwc99wTclsnbTtDCtrP6S2zJZZgO5IARc7jt/LzJjU
woJosca5m+ozj1whj0uAsUfUUHnNPwqMs6OncGBRb1iLh/R9ZaHvr8nvJMu+
n5gwdnhq0keaH0c0mFYym91jxprTAIciBdANcO3w8nJy39703Mfm7N7HBuJY
LcMRlUYC2RgFwzpRHh1fytRBE+akpSOvzMZufkrtFSgXMftxZuaZsL+dU/Hz
3lutI7IIX0TISMmIdrfnFEAgDaPWpx41AJleACmmkmd++94KzQXG3K0p4Spc
n+WXVzDs5FEEYHERRC2HZma8S4GMxk5HHs6EOEi2PVTm5+Ij5Z2TmH065bx0
AGQ6QfH/vDMwtViTJPiK7g87heq3K/B8rbr7+psDuRQRP2DaqU/4mg55Cz7K
NElCJfOUu81Nc6BfIL9TIDzVcRVOcvbYz4Er4LZYZYJtWyVw835QL+2IjFwR
9r9KNCkguwzyFb+FEl4C9i+6XREHDjFD2zZ6yRJUCpPAis/l985Vc6EomOk+
Avwn/Tz2ABGFIs50XzT1TlNVSQiItNxELxkp139/+M63FqfczRnmk3CgHmAV
EjWOXKKyZoBt4ZQXJQgQ9x8+jHebG0z47aQuOLCc4bz1PZ6x0DxTvtwieGId
TsbXjlv9hPCWDLpmvrJtt/SotsNN8X3PhNDkYpC6Oz0gJBIou7NvwVVSJPVW
Ipnq5XNfS8XeUXw6Ufkl3c166Wo+XdTLVplHquLPeJwKsHX++38gxj2cTMvJ
lr+H5XqrCCTcgAl+BDkIi5Hy2j0rvHTXV+ErZ8xArfOO6SMPSgnH1r+XsWkd
Xza3/fDR8nEm26TsBsRuo/c60uwY/4hH7lZN8UOKbrvJddp780sVnNObzwSm
XUWrpu3/elF9Mp7p7pqICQPnQCV2+RrlW5bhz5rsOt+pVvXvi0pbWR1jNYGi
npvveQD0M4i8iwyDffZa4Jb2LepOy0PjfyRTL4/Mj1h9R9fLiopxqRM/y/7t
njwT6OUs6LtUi6PHL4igRi2ZxH27Mh7e5nzHnik/2KPi5mmvJCHTxj1KfuoQ
Feigc1iWBX8eaJKtEk2Vurnr8uQnVFMUlcgusfad0lmyaAllR6cWEDPb7o17
kqXA3MXYJ0TZgaerLIBKKvnKCrTj2abYiSdIyWBSscp6RpjAmWjbC7IhHQ3k
TZQR9/E3bIFKrtP1kaOLAPDEsMazU0/4Uzh9+ONvC/Qv1aUhFPu1FK60L/4M
OVoL0bgswhRBEkGeLLQSNeU9tqRtiFo4CW63zZ9/gz04+ZHi+jM3+ge16sKM
iPXRqOXnnzqBSFYipLmy5LEdTjEpAb2nc/CbkSdW/rBYwiYpPp1ISzi/52l6
W6C5X2ApU4uOX9NziXP0Lgxj+pFWGxbAwJopVu9lKwQfR3rByy8kF+T+65wb
haZG+v+04dTvIZhG6asoDZcr6s8UwfUdxamoDMlj28s7iymyqloSIXAgEYPG
xfF1bQYBHwLmZ2g64Up65S1tnXS9nYUCgPe5RTA9uUPbe+8mDqCTT7atTZo6
pUKui1llaOeLzM7U842Vuy8dBLg3T6zZYo3jUdwYl5zuZm/aezjGZisFbz2b
gMsuqfMo2lAE6Q+FSSWIAYIP4Ev3Ym4BOGSoBBPFsiN/FD9HnkdkNH+/ChiC
Q7XiVtGzmNMF+IQlPn4owX1QqjJ7FgALIDIVDImC6iC1PWdq8XGPA4fcB4ZT
dlpun2U3qsRJJMIqtH8iw1IrYa6fSVvfZ7118WT5GvwpvMQgHVvn1f3A6mRq
PQq99Tl4xxRaVvfCRhNZR5hCWCBTV70HKHbxvq8RnezpbeiSSJAGbY9bkNwB
8QwU+WlwP5NntlmDQRSZQ0dg0nidg3hi3sl1wKM4G50oCtWE0ZKGP6ki7E+G
IN2i6MaVWsXYyZTPRBb9p0GZp8oyHzlqXL1tV4zKhwav2K7iU4kcT4jSnj23
n9TKdl88frKJi/XdqtwLTuUABTvOBSN0i8Io2089D2fTfS2IBUHAGrhYt+zX
/Q2a2qDwuI5lZs+ce2iq3bzZtLtOlAtwWf/X4GKYi8MuLQbghxJeItcCPzLo
/+Qb3CWO2A7d28N7s0pYhPL+41pFP5tLu/T6BU5ImOCZUpFEkgyD0iByn9nz
5StatALY989ZkIxE/SVLXVy+Qv0GMD2lkGwpxs5dCZ/Z8Cy5+AnFo5ipCWbd
pPoWVSsncCx6rtrUMOAM1QrbGYNgC4PQ9BgjW0iAXsM+Id3TpOvgz/Xrjqzs
1R5E/lZf7mawlZpHkLebdYfHNF3bgBiq0SdxXtNFm+iUlweWCB3FtJ3tED4c
W2oHSSMrhLubwS6THTbnDJYux0lb5LI/LDZXkCRuOMf4UgmlQkf2W+jJO7Z7
0QrSOxL4TBy3IzkLTduOEdw0xTTX0jMazMHGjk9Jbr6kYeRMlsF48b07BGwR
M4oBR5Ef8L/3LIrFXYLjZdc9WQOc8BIjpH5upfrC4/QfqDfD8vOl2Igz9LAT
A73PZZ4brWQGltzgnW7ScNOM/LcLFGD/2YtiwbI3Ru9ZSJCDv7zUc35pKB9h
XbbzHJWY7gbJsAneIYDbhUDZbfYitBsbk5XkSPQ8bBon2yA4kIyV4VY1Tihm
DNhiP4cXRP0iN620IKNdx6W/Q0vnfHO9a2YLqpkhGMIpaKeNx1KJLyUj/TsC
f8t37/J8PyXD6BhHc0vodirBUv5D9TAx60ZIx57r1jhwd1XTYEqseAMwhbeJ
5LjJVBSz0e9OkezpeTQYcU/XLpjzYyQR3F1auil5dbGONOEcEj4xP/8ocxI8
ikIezyOZg7GzOKSX8268i5TpMqFke+E7P2NDsg8+tzKQ2Z9/6KpDZ64zlLep
9Eqoc6VHkU+UwS0FBoMZKIF7aCPFOsHjRPjDEs6J/2xhZEsHC6JWPlWglJbp
B+Eys8nWGDtmC/saBBPRbnfr7ZmkxMyC/ytt0HL2St4qU74WW9JB2tFAthV9
qRSCOZf0PqDv86xlcH6E4QtGMsecilO9sRmiAQ6ZS0McixH00G73gIK4KHBZ
Tay3u0HpQC0NGzdqdarbwWvIBDDHk1PTcSaRDe4Zz2Nl13dYrCbJMdz0nMYd
3xTiHh88OCKgknunFnRUg1CsKJOzl4ubgbKmfkY+ZHTlBZAgSQ3vYei3bUgj
mHjOSQwiX2f4zbB63smKqWRDN3OadbKgbaWNOn8Dty8pIwGRQcB+WathUyi/
N7/PpPqvIsNolnmGqUpKq+nFjGxYXgenfsZ4UJVhDk3QzXemenEXAzljCVfU
3OEIKHrEXuiyeb5ozavlxESy5w5y2Sawn6K1tJIOZH3SMNta1VzZ7MdhopX6
S9aM+XN5YA9R+rnUfk8ASAgMBCky5nzNpflPK80I+THzOmzTCxap67pHOdpH
xYL+vx/JP0ABX6dEESGr7RE7pI2qtSKUrvHYoCFa0tBByCc127GYZw1LzZg+
07hYat9agdFEUzRgTcrdpsYjgVWFcW6sFNoLglG9Wz1PaczqXBA2B50jsfTk
vjCGRnJXWuWJtlrIFG/dzVde/QtXHXsW3xgc2uu9dAMY2viebCHflKZDYWaX
j3j/oz314DPkMD0vd3gURjSof5MqGvBnvzzKQwOp5fe2Yw89VJpsq1lMkTzC
2UKeWm8ST/RgjrINeuVGaErw0Ch0zKl5Yeq/zouccRp/tWAoZIKXTI+IxZUN
KSKkKnx3X403vzmD87PDVVYqop6so/uRaKLWCWBV6gJzINAQhXDZ8HA+uWjd
UDTX+2l3LeCWlQ8JQK+n8rU03kAoUW64dFBOeMcPMUwBUA5u9iFWMhuSepTb
ypTGdcbhQWMtvTkDgJDDQvQU1VsDGcHbEhjXcSnLHhzFVrbdFGzyrPg9Pk/y
XxyW/SG4KU/j54EbbOmcHAuCD9V2NFzloQZDOy+sbd9j6iFKCJqOIEUjeI34
xFNCfouVwAfTgwGa3bviDdTmEezstaAGCarxth2wi6SDAEEfa1SBys48Cm1i
y9hL3C5SI70GJaHy77E4ApaRpjPzyDImPE9DvJiLrNWExOmPMGyi5BG3TZ0Y
pjhL7FJljMEraCsBZ3CKtkdskZAlxesjHHul5c1npSGkFlWr0B55CLZebm/7
LL2Gy5Z73Wdg+1Yb2H4XAbRBjEgztzoGBljae0NhEys5uiKmiTN9yiFUUF0N
XwV2Q8LRZA6WiVrRl8hyNxzi6ivTDjHHU06J8Y0lq5j/BiOUX3NG4h77f1FG
TFicHlxZ0ydMmJSBVK90zmzNrNazpzN09g6DI2WiXdtZF4+e+MVj/mJ6PPKE
VCLJQpCbDJMdalV3sqrmrRKJN4IN1lyslESOnWQVlZvrv3OaRjT1efFW98Cy
jnhMLGFIaoDjQc5Wo8L8LYJYCHQ99k80gHupIonCYnA0nfRTjqoM7DSKWVv9
d4dsg5cgLWhZDvFAuyro/WOCuJleGyy4TYEMO0tNVfoStZCtKTYj6m9j4teb
w6x6O56SOd4oPtAW9iLSws9D/uDqOC496RnZfEB0h1wVvzOiTYtv09DlpNuG
Fh76nANitetN4mPyXlp5VqTRTwynslln4IQrMijgF2ZVb3Yrg48M5+EOcrOF
J28YZhWEMJIcBmYhnBVecyhY0K0Cciek9z9ADBx91nPexykyB5o5H12eaqfF
6Ln4si4qvrjrhQPkFLPYZRMO4dOQKQ15xsXWFLo9qKMV4IA3AuD0YRUmL3IR
543XoNO4toSOqySuEWcNzUs1KJ9kl1YfEfj4orE6StPzydzLuIj9D318p5FJ
fvH1CHyNP/9NdSf2WfjbtzQF+UkXmPvkLOcCxwJx6WD4IY18NM4Cvd1iW7gx
DV+MfVUws+BQOOjO40GGc0nlBS/i6uXW1tOYKIuM4wAlfJXPxpJsBJwj+Lv8
0X6JGP0CCVBTfjlnJlTadXkyyXXMPlqcg34Rg6NjqrM3b+XcpgEqOuZfUm4C
VWyH254cEUjAt1dO5lxCRKQXNgPg9MVs47gO9hJ3gyIyFgKpZHGN2q6STMxm
f5lAlvVv4XzccY/uw8PadWmIXZ/LyKoRnc7LVFkCrm0B3ruD3l2VUuYX8MOj
7hunqrSL2WjmhV+7/Z2CTl4HWUeHWPd6QpKrabgPjja6cr5VcTdJJqM4fO6v
5ImhiSRSXUmHYJj1ZvTW5jL55IJQGZbQnc16ddd+HF0U4vQgrAuBvfYC6fWz
6YrMGhYzrjit+jkji0UQVQrOslWSQ54CFk7eFFKC4451W5zkj5Mlty5uYUcb
PTZx/TdRRNCoTmJrUd8YW2JmXILjqH2nlqDRzW1gVlLYWNo/V3RxWTaFx0ts
vx6teFV3fumRh7x/DZPzxAkp7sj1L4F0of+MDHaL3zmKkV+HYSrx2gM9DYFx
LAOQjxyZVJB2vAAXexIrnDQPhvr5emRLrCK4qyuMFofvrYyE3Fc63MRk/Eyw
PokIBGbQdEdxdNbfIrRoIi0/gxrrmKgrT9d4w0J8n4qvtcAP54QU/qcGK+VO
diIGuw8iywkHqQy9Nee6V1XNz3Mr5xl4xz1jS52rW8xzKkUgvoDuZr0hl84F
FfLP2MIx4DPpdggQWAtf8a6/Bh/YHKECHNv+zNHJ4sINOt0VtF5o7jsV9R7i
N6IM3IcsQfa827OxJNFkreoLby0ApqvKYtBZmNcN5U6Zqsn2KFfUbcZrysH2
l78hy2dGL92bQ2dixLgYE2neVwFy9hg6H4WFoLjMqGEA6ih9ZIAqD7hJiatu
zByzF0c0dc2duYTrwvkJOeNv5vcQ0VTj4pm1QnuGdHUh8YWiycqwEhG846ym
T5nIbd0nRZqBaOAoZ7qKlyV/hunuQUpaoLg41Qh5GmLrXRsOXoH/ZJXQM85r
pQWSpLPBBeLVzykIYLicrIiXcUUrP5PjQTuRiEIeJpwXrKvUtuHZhnBPHgkt
Q41sETEQZtTiVvEVcv3Moz1QTo7ex/LIRO0AS/gAfwMdSaNvprlFzyf5bS42
gteSri03/vH1NfMqp+VHMBPqRs3yCAF11sXa9tSnv/O0yeLOlkst0OQKmbFB
ptHnUVDLqDzROUg9PVmtBGJRk8nIn+fbQvunnSRJ2PkncrqAHVjoTEWTpso7
AzDrP1NVmszl6Ug/kfknvLJe2eVUUMZT4O5usX1Mv+aA7hr95P/wLUkjV6+z
hRm1eirAiTlnFIvkZ1zDsOekvdpy9mAj+Mf1iL9F3bHBcSVcXenUMvkerjSP
T86KqnM4wA+7r2QpAb69kcD1T0H1SKcPiS5aocQymilYx0poxR54BUNViCZy
TyttNWD9NrIm60DeV4t/ouQ0NSQzmSXyoNiEZTJtZYLSsCdd1QNi08uVr9kH
H1yqtPLXod653stXD+FkVZeSkpGRohLaRomPHWcfLN5S14wHS9TMb3ZTBxpb
KkpTJoWzXywLPp9gaDLNtVNjH7eniL+drmKXNmbsNNeQ0RTkT91OaPT1bskT
r1Ww/Cs15XyIXmX2oBjuKA45vBisDurxqb+I7zJbS/kXIf7DmAYEPKcjaGxQ
F0qw0NdDWummetER7PsvU0D1Nti0OzQpYIRA7yuaCTACsq0kzt2fUpoW/7LT
8WCWv1/dEOR0bwe5/zxCxE6CVHfpX23UT8T9nrEgwHUR+OOHGEu7+2fYgyEw
odrwY9HIgQdEmxAE9z6/7kB6gPU6YLd8sMMDYXknN53iNr9Qck44ii1TCTKD
i4KXeRM343jDk5M/s52D5WrB7B0L+BqgHcIAcHAtVWqoJGkCA+EiG1LymS+s
cDQnNqoyLV8EBSk4bAo5hpPddrobkUEqr5DDKVzlPraz+4dn/18lNWWCm6OL
ionWvpjqH8n4jivJGIvLcmuu9KmmimtqxfxtkEPQSEfzq8f2XePrHyVZ+OSZ
gyPeA0h11k1ylNRl3TIvo/+HWmJ44I9qmfFIa9DEfgm0ofZ1xpNG+lX90RgA
PM6TnXrZpAH197K7zLu0wfTJ+S7DbXnMIv/7O6bdM816HHv5RHN4P4xYRopB
NkZH74BlPgsqpJk0JBuxq4HYZtL0DGFOEP87WJRcGObt18P0LL4m9vziQCSb
MoERiAlMukWXSXE2rrlG4LfjkDcYXRx9nJLQ0c4y4yuZXn0GE5zj7aCwvvNc
EkUczFnotVxLCQ9lYIOQ0wHnqNQJIS4zvPn+b+nY3W9OUaOifP5GdDMof4sW
/T33cm+9Csx+ERfVJar/iQ4phbKlt8n7qhGk+CR80EdgfoxdWhSX8BBTfGEa
c0RAPzu6DQPxdntQ41hp14E10gL7lmJtsoO5bWoxg9/IJdxT1uQ1jBKk+bkx
PP9wHs+3w132ZGI9wbCM78ikU1nNbYuAlVVttAaEJsRBOQCipO6E0prF02OB
zkbld+/UJ5UedM/r1X+km0oLi2F3PcRaPb1NMlYlci4OMmRt5+tzjTEPohZp
5T4ZZpfqudjqLQYGTQDQPaGbHGEg2pNOQWeZxKZ9TbauzpxgsOuYID+qnmtf
mk/UDztYltVSzG6vFwYJorW0W5JykNdGKLWyBNR1Qy31lCq4udOICw47cuLl
/DgyDgQSvzldhRJQITSjM/tnBr6XADRZDjrLOmyW3k7d/9OKxqUeRzfgji9X
HAILTz6NG+Tc9nK/cFQzghIcSMSyGEWJnoLQBbIj/ixqy+OEensogu/IeA95
Kp80mgheo+JgcBvIuBzjXM9jbVwWWyfnidlu8nDz2CmsKRf640xvHF8n+G0A
HssVpjYGq+0SKFw4Q6zT3QFwZIbqTDZgGNTyDwG/cmI8TYZCYPVJ9uWpcNjX
6agnNQqdKj8YyIGskjm57gOgx12sYBSvNG1yBoXtE6cY5R4Q3/DKv819mD4s
cWjBuukOxgeWPss5EUe3G1mfA6pB3E7C/iQ9Om3B5JMsLDMVqc0C2/D1NQpC
xZR039zWqNYKzEgIM15C8dU/K/94eTCDHJ1kMZe5p235s52/MH/nnPxWhoGF
t9kl+Hx1F8OlSmbHALG/jZC7dQSy0Ek/d6pO/b19T7I9IzaAKzeZR0UHGZhm
/S3PGQVP1B6JDRBiwOGhaznMPiB9qDnfIZ6XpSZ0Y+kE8GfCUg3Ct4oxpqHM
Yr+t1P9JJN96z0yaUb0HTCeAlYyQ2UCqLmNBLHzx7MIbdz+/O+ibg+A/mk0W
LX+c/UkIYq13ZwSZ93lKo78sNFzHBt2c0kR6iLXSOiH9stoXGlIL7M1ghd+b
loU5glo6q5MAPtJ4CaOAs+ZN7XkDU24cYIjoBresqwgQ42MylVwKDA05ewUd
ngyfUGQFDZHAtsPW8D4uh0FE2hSybxDKn+318YeSZ6UM9kYb+YCssXJFMa0n
CWaHPF9D7fWYdLs3ULw3dej/GizpWh7EYrCPVCTBj/idT+ktNT88NH6CXjGP
l60EbUQT1klENhBsj9z+aaxY5/P5U+mP4+2g4/EkbsP+STUWWnLKKy8BqIFQ
j8Gi+/HNECbpHDEzoy1m1kKI4JCTqXTtjP6PNqdvUHS6+DvvVnizHj9s4h2P
VhryUI2nuu6mv5MIX8Mqm8Bz3i4O4/WklIG8HS4wnnlgmrK84ghLmpRDZEq4
cjkg2KYQ/GY4OGg/M+Hx8o8T5nEzO83MkLfc3Nw2mui3GdD2KcCcVhsKQqtk
joZzaJoXWSjt98VZKR14AuXp5qW7RNg9ySgevjMeVjFxxXUzJ2HCjS81zqba
AZVz7PXP5O7N9ep59Z2pPU9B8Wgw63Lg4U28Yu3/jadFICwQLq9lsy2uJg3X
B85ju98POANbTF+p3hnO0M7FdwhJ2pq4L6llXfLA/U1Z4p09svFJpKq6/NNb
aMN8YsgXgyaVo5n4RCK3Z+6B1AAJPyKiWuX/awiXllWNYtG0xIWQcGvmdfgk
WZhus6xV1hWNEcVogGlzheVRdbaC1dHzjxMLI5wLLlTejJmMdserJpiD3mCG
z1RsDiXQuIpzncH6OFrRkTUGcpYLE4eY1aIf/LoIh2jW4/nLwgsT6IXGpT6w
mX/Xx3/tM0t+tPS52MTmD0OLtOb87OkLDlz9m/vu/OMiXmFaDU0vBYfYN7x8
edrxXhOeNzmPx0HXODB/o/veEpVc4Dd+1GIySI/0mxk5SBBBmYZi17ieJN0b
mWG9bc4DkEyh30lvrdaTRYGFFrc0quinbx6Na90OVKfIX3reF9GmjdSQHkjT
KRVT1lv69JlBkQwCqj6pU+IX/2PmE5a97H7PTMiQQD6YlIM/Pn2MojikIsZn
hpAppJXkF5ft2CfnGAm29NdlCPXAHFnWjYRbnMyRWlJ4LgJkjJkF66vGL0OC
W50EQ1J6mDDCCqZHxqp0jpc/VKqqGbaDc2ARSCsO/zSWOTVPqts66bDOcefe
AaV62AIKoVRZ3E5D6QjN6hW5KiniuYaCDNI0GsfBQbODNDoGA3rwK0/KAdDz
m/Grh0i0Kkq3i7gKShUAoRfkX6aHAanb+etQV4LeCQ4aAszfjHSKrjDllwus
DLEohVLpYLlChkpgkIN81m9EVnGTrMseN3rUR8VSuPpztFo38SYx07jsD45Q
oHN9KpHzUKYNRf4V7Naq4Zlo3B+KG3Kz+AaFZ7YDr3r6IoqBptN6Oh1vDi+V
xeWVJW0Qg3/8bFxiDs0mSsRATcDOyCUXHxd/0p+stmgrLYOeF/0M21m2Edzt
6D2PS+beJ1oCtzie4+J1MVJa7tGNJq6BG8lWmDnOx/0sjJjKzCnwekY+2Um2
sN6h2EF6jRH7DwVFuqfJKYd6ssRc42Bi9rCq+enHl2taj41V0CFj1ydMmGRA
89F8KYPH+5dzYKfawxrUgFI/sZwCQsvJAwcKaYjvu3smK54sdyyHhgny/lpv
xLciO/4cDn8/BRsiM2MBZiFphJKhiCbEdzWvVJ9Ewk1PzvVCFJ2RTEP61+/A
A6m+615tO5RnG0SGIpmD/i2dnIu64HyLOQXqWJ67fN5z7IEVWSUYWLxdgqtt
LbUlnK0yoHBN5cM3WFtJKtnlq24pfCBeRjS0Eo5HXISF/jzxfmF5JMcvYV5a
ToE+QlHshe5W9Hb9pi5ZCfSqesDh0Fkj6uSMb5kvP9MnPEG4D6mB7OxvYnZX
FIeL288e/EIYrOR6ikDSoARC4jfuih85yHUk7FTOgtxKq7RuHK84W84fLEPu
dInlMCgwLqJzAq+p5c1y/No4Yj2cwkDhTqJmGyC/a2vHT3Ql8XbS1+F3luu6
BYf/969w5KDqIXAed7NYQpdD3XXewHgNMTiPaVR0llTnsXSQidYpSCdn5XFx
PYYM6b4JmsbLdIcL81SwzAsR80JT6wzH086sBao4LctYS6ke0HgTh5BrRl/j
qUtIzy+ehsyNtzGAHvPiOJPINtpw1+eepC2PZpC5ln3ovBwk06e61LVUns1o
FygzvK7LrUvd3O5EzjpN6or+WYuM6P17tcjOznY1qP8xog0B1a0UJXRq+OAI
bO7GXDz1/uG8wvTJabvakXNGP8eF0GdAI1oaIuqwq1ENKdt0M9jpwbTDO+BR
1geDen8PApFeSy+ZSQqfYJtwl0fYMttpycIB1NcBXWneK2cS70FJ8AMmwGeZ
AxWFiaAD7M9G9+zNoT1jInC9HmCQI+qTL3JxMx0Vbk6Q+7aTLZweB5FgGwSj
Nuz74leq9J6d8gzUlMJRpuY3gjFz1hY+8hz11WVUWICIPT//vrbtZULxjpqN
ynGlYWBYJOPQRGPwvvIttE2sMyOMZLOFRh2rTrnTyfqfALAG3gv98rYO+HuZ
ZK9BNAf8Ge1k6ZHvwpcIFuULBKpCuqo6jJRD5CKqTb0EaZFctYqt/irD/e8f
Aifs8Al+shq2ooNXcUTXc1GHMQTCvUD04CzfFhZhyKpg5kGAWpJQw13yxEAH
wVpy+0yAdFGRJNlsOTVk5Rq48/ociGXJ/VqREjpuRLNFyd7M3BNfXngXcE60
7N3y15SLbxopQQ5gCYX8mW1oA9TuRf7pkS9xmUKYkOHVWIP5vg5auW1ymezc
yQCf4TBHAEnrI461iIvQj/FiGXC+qpauZz9/jhrckilpON4IGe1czlfZGBB3
1eUu6IlVErBhLeZqJQzXGnOFyysBQQygbOENI0r+atsugKMilCEKoWXhXuKG
b9yREy33+oZ42DlK/4L3x/cY17fNxXKfXGDX+H9NKeoPIeOIxRqZiUvTjc0b
eDNv/AT5LjCFYEv4EGD6R02nY3L1+U+xTVw9ztfAopX5T+GUbkdQm9kRCciN
g6+sIn1V8Ezbe6X0mqKcuFF4fW7yhsYQTyo1QUu0VM4HyRfs/UFW+zvyOafY
fCuaz7b58GfcLcEDIhOjd/Ye10fTIEMD3HSlDga/KdxbbcZIq223ECoZ1GwB
wVB+bJ/QcZmte7lHPBSWBaNLU6FX6MuwQPKU1+6aCjurdeSlVowTubHPBHY3
xaNbAl9Mx4acCKI9f0LRXO+x4suu5vUheCfq5SA+8VqJfBzUnRQP9vaVynKA
OW0iejKED+UXT19WyhKRX7pXlQGyfmsAoCTTA39QO+wUZZH+PhEVwX7asxGB
643rRmXdTpZU/Cl1P1Ip0VDkhYM5Q2GG6ribjrQAh9OhGLpBK2f3XWCvoUP5
Zk+vKIKjEKPHqqZdAmLVAnh5I6gJEGngfnd5r0EkpVjHuWz9wmpF6FISvxe9
r7NqcXoi3iYmLk0A2f2p5VvHlSZW0nqxARIp/PDs7a10BriBEmMGaXL90Lnh
VpjNRQfNcLyxZG2Rs9zmHSLL9UpBFGzR/QbVck1nH/05vs8EWd7LGFkZXn80
jW6FPMWf4l7BZNOY8R7RN70JgmlFZzPIsWHoSXEMyefWNay/BpHfi0NDxXFM
eUbV482zCCjWoxCfhPaLla3XX9YY8jZGYnuuynrBRU3v3BDIMRLpJ5fkU7ta
ShdrNJrPpT5Xm1hRp+0J9zhZJJ40cQOhHCrJgrY5PiTvHwjM5nZ24vgpsfxP
aKwY3CdiM7YXsP0F14bJVEYv3jDQpkYzGAIBUCbvEUeg/sxa14Dzkaxu+YCy
2zRa9II6EMFk6NjFzNBvXvLf+sR2bG+09MxxGoA8mU3qgvF2eHiEfBuRY1wS
mR34Dhszwj0RpZpGKXRMbW4OhEBI3ViiIo3QaTK9vwd/LuRrytZLDOlQ/AEL
mNjTJWL6sGMu4bAHN3jlF9uAuJnFXVbEDMxCBPsnTPlJnj5cGXLan7wgiMt2
+aphl2Z5lmGxBpcAhGjkmm46M742Bn6/khKoi3WCJeSf+2S3cxJAIIkj+Xj1
retYc7wAjoVDQyLvaUsWBCa5QOjS7XsbIT/GJ4GjHSXY8YXft3PsmxEMOYww
i8CXdO78frNmA4qUzE61Nie1simwQYA+BxO+ITSacjvbJMdUS5GGpHUZIWUw
09CCMiAjhkDo/V13z20z2oetS2h+RIIYH6x+hWXoMxOUe7kee8jzn2ONKx4s
1lWTstD0qLjcat4OV+NdjfwlpN79+57yE5RfHCg78+dJP+Jw1Vpn1C4qFlui
9dBoNHfu3UxEl65VdBmdjpQUr6TWVXi2PscZ8aJrvMdZrHDGb0n2UN2gJtPu
CmVvR7xRgaT85qI+MPVIfn9bHxLtAaKOp46VUVn9UjSkZw12SAW7eYYX7Y5g
uPkFAZRqodUiTgjU+zSD8ISKDAZw/LuchMa6esQg0VJaVYLPTWCZYclfSwO/
ioDi25zQcJSfFURvvcKMkHi8BNPJUhjvnr3UPSYqU+2U5f3ghesGyAhrKE8Y
Zol6AZamx7L+myOSA0aLtzHNtpM/LehamyL4IqqUvyhpXuHH29cMYktkI4FC
PvUAVwlJN4uV18qeMrYirfm6TXT/T4aM74BeOy8AFrLHlbpUDD1XGDuv0m3O
3o6VN3817f2Ctu+Sq3nb2fihycZdMr/3vYwD7rWeW5m0XP+qvHKpzsVhqa2g
4p3jiQ5+0d3iiYY5+r3hvLXqJzPCyDH5I9+6zEx+f/9H6Klf2MNMT8Ot3TTk
ChtBfZKIciW8KbuxzkR9XiYhJSpRY0I+96+CGahP9QeRoOMoA7fCpZXWyOXT
UIC+v7MocAKTcfzD2yWImiZ4nDwlKJJ/3EosvJWwAthP/ljOn1NM5aTzuKDW
qk3bM3k6x8H/KjfHcR5f+uk6dbijjlwfKsrvC2utkUYNJ9fBgYKZrSRq2z7o
XKyo2B8bEyyyOJxHNm6QRp3SIPtVUY5V/ndewRkImTN3M8rfZZsQaZz49bfv
XHJ9phkSrjoHymIWUtwIr3qcNDI1Q4d56C3XD2ee1MjatsrgvgrFeQbw7C+3
UYqiCaYPoL7Vx/yJxWT7Dd0jIAYq9dPI/SWoCmM28NbjQL3Y7kSUcx9Yeomm
3JTjYYdTSSiBCkvL36Zx+oz0DRK+M4ZCksTDRIX7e2TPngU6mMD87CZ68jE6
Ei7SJ7+hEOiKawF/syhWvrGN0s4TLmtebvE0B2FZ92U/6tRw/RtOledWjpGo
HGYHZ7wZdDh2v8R4fqinZtPP8thG/AYM3nQL2j3Z9hiC49ZNwO+rxyFf/ErB
7dj7Xf+JXK86Iol2DF0H3QZ6FOqbY1GtPv3zPQTHKe4BKOr2rFYQwcuoZT7z
QESOTnmURl6YzhcXNPXYVP+n2tFMz8CrcCIiq46bNTem+18Y2/EDDlYP/Z4G
GItO1lgvhNQlmlUeIMl3OJWXEKCrUS04lF20ywlDqPzqapUDWuUiN8tKV3iD
bAIqhdRVtRObE3+9BCk2G8eMLCKCCnO2IYD1yU6zyccgtBY/vY2WXoFJqqSr
q/QGB9dCh8zuYKp5ONjuKTJRFhVa98ydB35a34X87ZwRTWVHFXcBD0euymfs
ZVWG/2Aet1g5KoVAIcG4mFdLuFMSLIPuJvB/5y+khGVkYB/iYm9I0ppp41Zv
nsNv7g4/L5i/tv+YZ/nvO2ZUpbPu0ktYtB8jYwmWJjWGmaevkd6CekjHhAqA
NyIfwOA6fEJ4NTRRdd2UiyTSkR31C9Hp/GXkUFH2Gmfp7BK63z8jOpfXDVvD
U8XY/CQcRVkxew/RuhW/wfstzyNuenK5GySFmFIGhUUArnpnec2p5ZsVXVP9
uRi3R2O8JHD42iqWVLma2IZJM9fMd9aq5eRN4RDvEzF2FhNf+rqbdONeTVZ9
yvky+RhI8cLGI30IuLyhfSpSRC7Jkc7WVJ+eExmgj7BOujuj3lOCrsX3vu1s
rDsR1p23grgGSpQkQ8z06uPMzyP3lWdt3WI0xmpo0NNkITBWw66mLoV2hn3a
zB8PdxT5iZA1EHM4d6eECCR9PgzrQZrMUkN3rMEsrGAiXEGu5l3Uf4OEjiZ+
r1gYjj0dFcWQQI8ETK54lCi6NIDQb3vk4uRZMEbKc9fzGupx1yAkASvBRt20
vpCQ7W+UC8U8M065HNqrram3Pn/gFyRKMYh6ewjoZtt/SqdKCLYh3bMYiqdl
ktksHDLMWfbA4NgBTmviGEVMMeWaY5YJLACyjBpmYbFlIuYAjKFnhvpHHHLp
q8WgDYMd+gNFZLIgvXJwd0EvLjDPOMOfBCTMpLupYvJ1eW1U1Ya2+ydDwj8L
oPuH0ul/Odv+n1naAQfbFolo97g4R4tzxSH0dIuEbq0HKsXYamrT3L1KHEe1
7zwyOj3ufLsChw97AK4a3BDnSUsqZM2Ga5b+pn+uDsTkqSkxgA+RRSRv9N5E
DzCgf86KWiyVmqPB0swzDBh+QBNkahJ6v6AeWCviiqSkJeSDu3Zgco9HZF4N
XlITW2ILYPnMpl1MoJ4Fy4lYU33wbl2Vzv7I5E1JjOhoyaOSzWrtVEaiRBvt
XS+uKHAhwtyc+jN97OrQZT/K+viht8KbXlSJqpp37P+mRrLymRcgGo8i2kT0
ojOb45J7VCedX8GtvdonGFVX33VhTLkimNtkc9dgj1R+y2ipAjXOpQdk+baX
M8OpIz8ziq6iaTHDxibCQxLQBOrP/FjobrHLWXUox80D8udM6yKg1j/GdnIZ
VKHzGiX9b5b/FpvVuQk4IIutnGI4S8YMStzIwGoRoMeABFlUVOq8l/B7UvCE
PzYW3IWyJ+zrKMmqmUFNJzKQHbQH4ZexQplvVND/CXBljTwK9h+fG8waw43i
I2hZVCRyUfBVbqyKUESvDNpudRKBkwjH+SqXorHQh/b7PlanUX/ECBiysaV6
ecLurG9pEFgxU585Kiq48/DLxpSjkCOfvFLAOhznt///arpyBeqZGqKTb4s+
OQ4jCA9kjc2yOaXyoT5QG4In1cB/skPJMK9WrjfLo8AoYPZ5PU5yAv7KY4eb
kTAqE29cwElyAAS6SlZKWVGtrrXTarRT1ZowggPDoHrUx/VKCKyAwOPa0v8d
UlW0y3HD5axOC8hSJ9TA4pPhqzQXMSFztd6DKm5JEnpYwVwQArDSQYJ/vAfw
KIeQrTiAaTuGAoyJg3YsmHnOt87/Rkx5Zbs8iBbk1djpCAqSBzHHVLkZJR+O
OnJ0tKA8RbcObkI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGOZVjEvF4rQT/lL9cF0n4yHtosgrJ2T9n384t5zzRNRmTKLu5pzoiBiTYEg+w2LXp1DcPGkxnZQKkZFp3DeXUWSv3ULTKzN9SJVmEyVXOLEEYTV5IrmMjVyEJqagWeKAZPfHYhZKnmThwGFUkXS4BgiZWS0UlS4rZhdcFb/SsPCYCQTmZiHeJGPzZ/2ubpUuHhea8TacS1R1d7C1g+r5oOIxB28V95ly+H3VhK3Cx0A3trB3nYUe07cq+H2SOqnjssobO75YoEOofS4SSvfVIET4KsKFyUHwlKF7b1e0M2pBVFhaMYtMSawxXyjLQxQGtnOpVmrlIiG82d8sDOpk2q+bzVcTyWp4xZXajPUSCbMs0VKohEMGgsChroYZ0dMlQYE0ZP3dNwqCZdpHRC2f1QbMJy5r6fvZsGLTJ85bJFSSmftECOTVHQtrmIUi++5V6OkrqOTc1Tcalxh25COTsc0p2aKbUzIbFlH/TfJ6Ar3o8g5Ti5MzyCVnKUtYyogQUl1VVdCmojoWOqFUDD3j8QRs0ubgZKkyJq0r4iYRex6DxNqgtxQdo0i1SopMf4S/Dnb5xui708sbF4Ht3XYTONvPzTUdo8oEQjWmu9NScELA5RiGBSw4JZaGYB5DCjI8lPxPCw0Nc4Ic8vFIbGuLI2vgi3tsF3imcwM1yxgTJiU5lgNrZtrYIx6723FValMHpGamhSsyCkNw3b5jLKTy2dmhDJ96901HNF4duFn1H6Vk07HwqWN30qiNCJvYB11U05ddOBgwvxifsw+SqksnWOY"
`endif