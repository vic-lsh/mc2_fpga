// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fcfwdxTgc0t0bGgoAhm96sOOVRHjTRZu38a12lAV3M7QThSCiKWwUSQYEQ3t
fJnjB8iTsnNCIepkLeSRdNN10GAJnQRA1ljsKU9d+azngfXcjLvC7hfSndVg
hzM4MsT9c4gpwkJ3T/egvyVzBw+wSZUUObQyc3v1JxFw8sSB383aUsjc6t1+
MbtD3lk3xgalEDXOIye6BMI7pc0CmDdhN2qfi8v7VogRlIRvnoV+XrV5ynqG
lauatAjs/J+WFBl86vLaY+tFPMD9ujYjGjf7JCo7XjifFPAvKKAGRhv6tWFJ
m28PHBYT4AHDDnyVqO20gwBFDbXU+keLIUdRbwnFPA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JcOkc4VZ7Rw3lzttuKgLUPNlj6aYjgQiT0wNQMIt4TvWiblcj/HJno85PpRi
3rG5VloLF+pmkMae4pGuE7YRole0ub2YszZQoHQCMSLshnlNmnuI0sdf0whL
jNul6vBej4fa+opz4a9uTLtfUwsvrqYdd77jShCuEw13gfxo6O2pPlZoVubl
yxcOBnTYVxx4ZimLKZndSSbYjEg3H05FlFnn9wr4neVXv8+wvAfCcv9/0k3R
mc2zEwuxITh0KTLVLk8P4jwD9c9tZIbxgZI+AxtRSG6FHmy6jw99HFmFzDax
JbpbtM0wZPAQRF7R9yGG4qdlbFhv5WBniO+04h4Jyg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ut6qwDctaaWTu8HT72wEJC5Vxol5vlLmuR+ruK+GjEKL2HM55Xeb836L3BAy
V1XFoQ5mHOAdzW71IQGcfVF4/dFdzXU7hdvTZMnLF3JcbBYj9MJPZzUUYM3n
Mfjil97Pyr3HdPHc4baRydOnqUYOaxjohM6WzSl93SMXk9XlxkzXX5KaLnSd
QRwZCXjb2x48xSLgbixY0WPe2mex2EQCXrJNXA7RISPF9ADcQ3Xb2LV85xfB
/9bb4FL3ozpyAcuUgicWTLwddl211kvTpWLPQg4zaNJVJ+bl4pWaoynlaKSI
3tZTYwpIoVYPsRua6r8Ix+CNaHgPqscRiKB8vYGipA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V+Dj8kFfiFecYNwpNJUeB++uCr3tpTPGiIGjxfAVGQBFHFIO+P56vdvAG5fL
C73m9CJdAs/inTcPfX13H60EDI8dLQD4UPTAPWuntnqtVdMjfCNh15tdbR5F
a40Avq/OwLq2WajwA+HmiUAuGWHVie10eq5ctTKSh+YH4AWAS9TX/fYJ0b85
wQYcc/rldlTF/Cd1iO/qMVjdYR3voBwdT9+cKVwYIUhCXp3wUjZ6FZEC8QIE
U7VWCTiYVzThJg3kPlSh138J51lLf4hJFWBSUgk0BppalzbXMVFMazW03khw
vPpbZqu+lNIuxfc0Ijfj+0K8CNqnSC5yc1KkPbuFBQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YuzqloqDh6GdM7XZdqS1JPVmDGXYdX21WhS5b00OEgmbYSci30k9J1qIOTSu
vaGQnk9bm/npKpKilw1AHShleYGEkvavF288vx5MWlgZDpoc8a5u2+3Em25V
5Xg8C8ovcHqOpsVPcrV/kwvNDtMtU9U7ZpqR3xdhY0oYKZp8/R4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pYPXRpEvFuxHnRnKabfbhJVpn8xEosO4fnE7eRmnhLcVU+HMDedYd5OK2KMm
jDmNPqJXBIKuPU+iBQZa66VTnFdX2gWcSqNvdFmtuGAso0mFNUvYthgQmlGI
Y3Vv53Ob9kcbgEgDvHWsTFjqP7J9N/FHMsS74VKS0jMpJFtQnFuSNjthBMPb
WQgJNMy5imqisOAK3TNPAflNHRe0sheSLlcj1hK5SUSQDAqKJd2m8vprvH6+
zNVhW2ER/SLCblI5nESbYHhZOlJ0WDv4Z888+QN8IGVMyOQFQGCu1eXqVvZP
Sb2q7gQ2MR/ssoYFoazoWxqCIyB+AoStVZs43uGI/dS6K2XPA0gZfVSMT3qb
5gHNzv2lABF8ZdsSyK0n1MN9MEuH9GdWrXdrt+XcsAjDqQZ5sE+8OJRahgFw
lYiPbT62SRSa6EgNGflGVZM3XFaMiWWaA8JbazG2onRMbdC8yQoDUmW34DrK
HMRgOZW8Zpwc5WEP7waerGww+SCMg+s8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pTG3HzfKEZMkw1dMnvWHA+oC32VW0gInSW55/wYywWVYLKcthjb40fi8ErvA
1QtmG8Hkc2zKAAG9EvBan/8zIWN1l9HzP91WIWq2cjy8rYs80odd88su7Kjx
U+c5fPTjTguRwY77i6wVAdkaSRpl2GyLRiuIYPrnho2vvSp39Io=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q8lbAJYw1VVeZfzDWiEVebmq/izvIr2WASoZXSdofLJQyYGbDo3zEqvXWgH7
v8Wp0CW/iYs4x1P/wrXi0C2dYZn4h/GvmZwV9Cm/aeFgx1qVsS9/A3+B1O6p
KkbjCm/hsZiHUUwv4nyrLmlO9MgQCIlVJ3weqL0UHhEpLblx+zE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16064)
`pragma protect data_block
mHV09If6dcD8oS4/SuRQIb536FNLaKM4Or/U06b27KwYfQxeLXyR4VFhzq08
u10JxC+iHO2/siCAu4E6kBCSwDMFOAJmjgcszg4tg45votPln5C+V9p7w3Hd
u+MymuUABOqJgOrfOA2Lj9O2K9XHgy3kPN2PwlF0bQ8l2TjkeFvy7Ua1HDom
uMVsL5fvQz6Jqtgtw03u5ToKDavdY988Gfa7WBQl3QjTK26kdooba1C0u1tB
VE6WnvsNPkzu1J26PB59d4MJkceYhUeok3IqRA5TcYo87wb3kvS6pLkkJp2c
hxB5DbRx9Fzlg0afW/GZNPn+B8MyJgtRUYa2NcljRq4yqnTK4Js49BN1Sd4o
50IsWJ9hpgoSbGJxsDSOeQyU/MhKGwSpMMxrVuFI/TdR2zK9Bxbq2C3316U+
FdVbgbmyNV+RSQWdsTQuKmXsvqdcOhfdfeg7fdHs2x9sWz8ibWt4l6yCEFb2
+Yo6POxDzOucA11utb3/vxj5penMV0asxKzpLnxojDXyH0vxWtRMHvw+VMPT
Skh0ygrLOo8vVbgBhGC3A11+fdOO6sICF1X7lEPOBHmHtdOYw2N4EdmErDOK
ueNduwUH2GWIbVwQHwa5PHG6EFxBjGx55UHPbdXm0vL95GQDnUUbhpLC7Ysk
SWIEZx2NirB1GJiIU0m8VWDB0e+xPfMgDI9d5uJcRAxh1rjq8oeTkxNy7WJj
t0Adwqewq/+9cMiyIOrymjoe97G/vOHfrYJE0J9GAXoQNZpTcJG6diL6AX5j
s86QuB9kWUXKoCI10g64sPVWb3YOXkR03WrHYctltnx4w8gw9ePB6AHPd/z3
WMWVNs64worXDL85AtAv2C3YikFYLCowYVjHG5ms3nOMHMhnoZM8NGwUT9eS
MKERRnDdzNVfRITh/9EZ9ZgRiH8E1ybP6ScGJdBDwvPmFFX1T9O2ozREba0H
i6bEfF8kIpXMnK6V5VG3NSaJLb1tHNfRzK27fyqrQWP9RpPh6ucMecNueV2S
WqcJvW2mFeLZ0Naom7BMnHTrajbIX1oHQRrIJ1AESWNEEjgAFuCpzupouUJQ
rvhj788EGEchkiyLVHAFKmVjgENuM5KB7CLwFScxbg/8mI26k52AsiWE8+3T
2e14Jbpnl3bSkEKSstWzhnFeQex7a1P3Uocw8GQhgsNrEvZB3fN8fBEgsXFF
ON5FPzFbeaZW6/lU2nQc+k1Axp3LTb2hWnmZgVKGYZ4Lu5YhUXoPgxGvZ/Rc
NJLjSV+QDBarypr3M65NZuaCaISOQ6C5n5EFg24g8QeLR/U8a2ff3CNDEGmX
9/fHJOIlT92QBE4StYFKfVWikD8VcrktWLNry2dNsnaptzWITalxJZfEgh6F
wv/OYV0S/iTZ/PQ3cpWc67Wcw/cRcDcM+AxPVEbfN5q4LLAPlc+MhZB+HfZU
S9aslHej5FAyCG2/rrG3lBm8tuqJ13fLakh0MAMN+O8eYLGxNK77WQqtgOew
xoPTfnMw64tNRhjSeiUYks2/rP5oPtYUsIOjR52TWjbVAG6WRasK7TiprQWR
a7Lr10Q93bHSZviZqZSCk/BTB9AJ1ZUfdYAAEKqezd4PzjBIVEmk8dy5cxuE
5aXHYRAo2xxRToZLU1rVd1PoX1QzYyzJ8QFDZjvAVz1eX8GZy8D6vRpeMebF
cRaCrPHrmlu5CiRZo97FuuaTLl2e4RNdpUdsCk53CMzrRM6Hs0iT657oqaKT
4xQ93dBag6DWpmRYdkzQ8DGoGP5tRtIkPB/6h19riLQ/PtFmC/LEoEYy8u1H
F7R2TeVpBJ/3hpeI76hDCRTYViuYUBnAVSP+4tSuKoOn43kYb7NZIvWg4nNx
0nXhORT0eRZEahSp9Gp03F0Ddi2JmmnuPKUFVQVXuDRx+SdpdHbi3wlvRa7P
yxP6YDsV4HbYUbp2jbDRCz/Xx0A9BTa3F29Lg/rIL8/AEAYHc4SjU0/t59wO
BV1stwE7Dj7qKB9wUWiXxAzCOaphXNcqOblKR3cZ9QFsedLPTf8RwqcIhy8C
K2fh/7dR4OHJ019dqx4E3FiQlsAKjEt0GUIJ8VtAiSbRnHhl7SJq+yz8jtMt
GER6EsZKdM39r/LbREGtH2PkeIHA12FBhcBcPsyRAIbTh8+kyxJ8MKf7hSMB
PZVvzjoGpyWNaK/NM4FpV3yeahbzFGBrgjRRawcK2P8OAJyW+JqtlibxUOXW
JO/W3SGItjyAHaRjcfU/+z80kREawFSVuGLtAQAwpKmYB/nkKD7gV0fy+km7
yviREKK0mCep9FOo1YWYAH2W2nmk1PEufQjWNOZSNSJeEy/ZJIZHKYEZz8JN
vRGiecYnf2PcLnOjzlKBC3xxia7JyaYwDhaoK7AjZ+4aRLHQ6PSz9cwZYvZ4
TEtj4ErtyXa0MlUNEpzEufkKXQ8Qc3UCWzSorTZTvpWa6zKTSFAzuKbMSG9b
axvb7f5hSZUGWk2UHu3D0mMD9xYRmWizCo2ozAFrn+0wteliSr3oV05bIICc
S7kLVOJl1k581Aj7nKrzASPhuDDoeL+fHbcycEH+/zY8sbZUWak8BYMtSaG4
SxjV3WvBal51t5pnkRTxQwq8+ss+5baswggP9EPym1sIYdW6C0ZYIcaCwFco
w3wVoDIbpNX1ZocbBGfBvUwK8aJsFIP3E0sO08eq0MMdeN/HHQhO3xJLjtf4
3tgc97iNBF2C9/6LiAGmu5yMR7OtDViQs4DZKSV50x+najXKSHil8dITI9+3
/DuP8t6kTmiqw0ztDml4+KxviTEEUPhM/6ntQCdn+pQLp8yOt14NKplX7fQi
chR/g5SpxuFfjSaIF+vv0Mn0uU256TnSXs3DFp9W5jfywXbfVwjhpD5RLXst
J0eUr5m06ZJiB+4Dq/1e2M76hH/hHEtL62vdkV1qV3Fa34xWTzqf7VpKaL3T
J34xukkvCZKxTqN9TqMSG0Sx+MogmOe/G0PpW+vpmPOZ7nFZ8fbGXiBNzYDo
O7KnEhn5d/lZnSZg6zORHDhCYz9aMXBN6nFb9DrZiz9NQ+I2/Utz/8zkMY8O
omufPmjUcqfVAGcfKXRslX1iP0YHKJ7FZ6T+ii4jaAl6LW89U6+7PNmOn2XC
PnT0fuzbRzYwmeSZp+EzEYsX/DAe2S8zJKZdacfhq3fZRr2gcyJ+6gfWJ4b6
Ev2K9EiqXBzX768hdJSjG77HdUsnYDQlG4MM4bJhGftv0nGslpl6bImYTzdM
t7T/6nvAlkdNRbjz8ZGAj1yY9/vMQ/LgRrX4/9V1VjMvtISJeL93UvsSGiIm
Ov0pAZ3l+JefzAs8uPVR4bbnYDHx6cOmyz0vyr1jJ+CBfsnoHVj80RKUkb8w
/mbfGOsXrmWADjaYpbAI0sFR0Xog4qO5wpqGpsrj1RqnzkpaHgyCv5rFLuva
ggr27UyUuQjAR51C6pvxNaR5ovjmKPze5sFCWs5Lei8fX2RcqRHuSbURUeAB
H8AshPjnRWXervXnWI1HsueYemHNjbEZEjYo4Wc9bnZwAtOpuOvSqlhOxiRc
OnuHoMwHo5uACk0UFM5KQs3GHw23/EQ2mN5/hmz6nmJj64pqOXcYUqDoHolU
khNTed7VaKjV4/HWRtrkdOmccRcLCYZkLrAXu7aI1+JexUxOr3xSn2TA+IeM
S1j+ymhO0e5jw521BMLckugO77Ixps6lvMaIPIb0JoRy7sBydE1jj7niMwHV
nGFM6rH8u+wt5plT0F5BnBlJKuZY+e1XqxflVmjW931kMfI+uaOB7Eryrht2
xK0Lpwxk+A1r7wz09tDkUkBlFIXgTtoILKOEE3CYNR1M3VmIBJJkO6PjZ4AV
45VCijhHJmNhGQNZ/p+qRZ6XRURYMGzi+yN1MWL7Kvo2JX9x4KD90mZ6OwmW
flRxKYtdadelCU9vhXN7CZ6GyClPqjVqUjaYX78pC+MCrB4Mj8Vt5HiKkFRq
Nk5EfGP6hko8LQM5bMy4IeBpvnbMbPjcIRA2YsvvvXwjcnkgsTh0/+MaZDih
zQgDwIkaRiISHwFaet21+e3SRNWljzoFWVBZVgDIja5BPmNSN0IFuiovhjeS
upVpQLZ9/3GJnw6fi2F3Q0Y9TLfsE08hxPzNOa4Juyg6mlwLVjb+FvRwsuve
vdDfiV/ukjRqYffIofqJzH6cv9S6hIHP1xm8dgAJHYaRuLRBXXjN85tTQH4L
5XrrvcYncTQnTPxMSKVJGkkBarMBEGK77DJ9JWxTLMHQhfJg6nScGP/GyFyy
2sztbS0yLY6hFN3zeeXCkKQWcRA9INDc9mFONsStDnJ2yE+SnHdAV0hxfOIb
JO0mG1darRBf+GIU7+Aj3dWb8QvryEhW6m0qFQupHf38POTOF+4ZKJ3dM5ze
VxLn1tt9zDnSpbQc5gBqiJIsFXKtpDVytcuje3E83y90lXzE1zQcmT/iietn
cEsVFHan5HsrqKDwU+jODgiVX2BX8Jyy73082Et1FdQwEQnoimjuMwsfkMYv
M4NFOAfoXDlETjCK2nVMoDo0oQ3aqybp7U8qlhZu8O8Xqlzg5S2D2kMPZ3g+
KsQT7o0d3FzsI+u+qWF6NZj5fxpDIph7bSGJY62Bb9YpCYlWvLMDTmB4UC6H
GgdNtQVF0V7y/gTbDetk7SkcAfxc8yRFQw3h/Ca85YrIxsINFizfqGiciYrY
drLMQbtoM5XeMiJdL3LAkLsFqwqzGcNlDYncmxztPMVXGEbNHKJj5mq9ntMZ
375jgI0j58u1l5lSolRZGjbco96cVVNwCFaNIk/fsyxmfJu4jLJ33HiCgEfx
vJhymX7/IYrl5tm6t1C9vUyvtTkangtQS9QT1WMgOToPosa+ryY6IOZZdxb4
U2pCYWqoKKOXHb5/QF2D4oAtoaK+QWK+yIxK1U9qn7tTEOcF13SG+7baA0Te
+6C17WcFJLeZkt7AJzPGKf67Pof7OXP8C1qzhquTFNOeJxnku0sm7a36C29h
zNwuKgpGVIZpik2kli8bvYyRNM3RGueaqWRq5kE1Jl3FrMgfxeCTpbe1J+vo
mnX8PQq+hcMQ4uD67UTXUWvMH5uT5GizPXO3Vb6CbKEq18jpWaaGGtTCTXhX
aUIwzL9Bty08vVhA+aBqmDf99aMUUmJqW5KhojOQO1UA1I3WG1yKS0aBpfNv
4ZYRvikV5ZU+cdNo/n0GcEOPdTT7r4zNFTHdyOiUPrULyogY/pu05J72e+ln
Fnb1iGGcNlfKkDNeSCBBvef4iTNLVJveqdWwTVUhNt5N7/AXbyladKPmL08S
pTiQq+jXtoao7zr73Cc2S1+mRRyX+JGNKnkTeG9GzQR31iFKQJSl6mMIZ1WJ
hmXsG7QKfVGMLXXEXsmVidO+qJbifLDUIC8vf7PvdLd7yOwpQ99K0YQdUJ/e
oLG3eH2fhe+kchBGjv0ooCndCOSIQdCMVem2xEvyjHJcycFVrGPjdPFcwFm8
Op13r0z3bEUmOonQvZnjnHuBUS8E18FnYfvOCMLM0LsI2G1qdM6YTf5kgbvq
xhXyPyzJATlpwOar4+qFZ5LOKDBWNbmr7TFDrLK2dX6giRKv0kH4qWHmaTuD
201J4ZbJF9VEYQTD39cXVUDzF+EY1dAs9U0NDFWpYaf97HO/lQvRGJOHtWEl
j1GcY5KVV+LFTLKZo8YFBZgub3nDCct59BT+40kWsRcHXJj6RPpKz1SfHzlr
300jOE6aYfNxZsFa5+S44F3a7Yx0HMSKDFIgJ/a+smfQD2xbmGFLme93jXdV
Vu8fp4cZ8zWTOBzRnkxo1RuVRXEEqiuFleWVfW/AzOq//ge5K2Kz62GlmQmf
FdeDuk7IdZWmJpqRcZU177pmMkr/fI+E/caPuVM+pFB2oVN3lGg3rw15vQ6p
QMC3F5BHq7ws3+qGcwwlQtNyJB+JXvLvZbPHehMi/ewYM4ESJxnLkEOm3F+W
MdJKSJ9MrxgpcE/lDBvdb7IeucW4oJVkSlrMpbq2inLy60WLj+mGpUkcT69V
psnrCQXfMjtfovbAJOc5e5OTQVaw8ijbQ44D8/t4OzHpMLw1KYUAlxhmxdAo
or9KanpUm+PfFvgDAKh/UJLr6VHY61fMmVVFDOJL9e5RH0Cf0m/SSlgsMVuI
IKCFf2gp0pmBlc7TroqDnjVZW1KKPUE8P7uJVjM1HXMNtg0r+R9mv62PoOY/
So+JskQ2soZW0EzsJKs6Rz1+PqL+fh5nMrmkXylddW37sTMNtW6GoRylTkfB
vj4zFvvLhx+aDlegWXs6Mw3GI25QMyUEVkRsMBKV4Fg/ItgMbPtoIhnEYe7E
bnV+z7nezAe3cXJihCCQ7pG06vJOQgjSlWXAatpbq2z2aLFzEb7aMDYx7Dzl
YjSBXKTg7rVNQd2uLCVO8iqmfo7CMBnVVF0uwNh6QfpLWa+C4jXlxCdLgnIc
wxX1Pea2DxoNFfhEYu6k9gAZuK6nyBdjAr+NOYIc6uR5F7rYIptTxfLRG8kj
ocPX+dazqmhQylMgMV48xB/ZBe/aPOgR1RyA3SPwtAd/xvGvFDK1HYzlA4iy
2W87UovbJXAOgMgOFYJ/fiyK88xL11QOoH0kpTec45HN9Kfcs1wxyELQnsQU
kblEoaHypJrT4zWlsZNme97nwjXwWpkduSadarYw70+DDNL2AU7eV3aXNTUl
Py/0FeoPX8lo2CXTeMQ1Bl75kAZxWNMCj0vMAGiUVXjTFkekChuLDkmMKFrU
AC1eMZkgbdKTO7EAJEhpkRCIlwLJl+jASx7rXGKkW4WOOiRP8u7P9Dudcq2b
jRtwBcp423YiuAJMFUDRzZLVIkeCxrWFJv4sVlSFomiDs8Dwja7eTO+nB7DJ
6QvRrCUVLklIDmTqpuo7LrA7K9zbaYVn1yFkHgfSu9C6Rn9N18nCrEeNpRsI
l2mBo/ZGBN4aEoNRJTsFXhLTGT9H3S29YUA+WNRPQXtuRI4wIZmm/jryfuhf
Qkkwpw5k7PSqHm4cgF0+jteTptqE3Tzc/yK4jLf4q84Yw2l74xBRyp0Bsq6a
8a1y3Wu04TEJOtcAyhbP6k8Pk71yjFovQg9y03ue3KaS70NUnO6EGA0yk5gP
Fmv1PA/A/EzyJK94i4UN3vxh3DoF88ZAgVutkBgh0OxwS0+Z9TtJh22qi/mP
q+8MMtddkp/ZSAZmE76rrPulkS4tSo/dztqvZDGrC6SBnmyXwUy7FmaB06Q7
3ZQf5xNi6aa8LXxyCqWdKBroCIttDj3WCBK2+lAAttwuKEfdEmk7W5ljXo03
ipLQgWtDN805GhW0FFu934FrO6evXKu2x7K+e77uPOAn8faGxuScEGbx+w+f
dTgj8z2ByviyPndj8mtJlr6iy1UdRkdSOztK0YvDUFHGs/KzwxtbDsJdXmTg
Q8hStL0WaAc8DI/bpzcpmxZuos6zsD4UuqA35krHme/S4HK4thEHxC/YJfnJ
z6rNEjV0ScxU3wo5sln67lEXlZsCcJjjM3ER/2gEpkVWmEAnXhNlW5SbRP4g
ucsVey2rZk58jWMUzvnyTurIFBpgzC7Cu92Pf5KC2++hw/qr+N1t4QrMLV2J
XAA9ItN8tSbYe8BMozwFKRXLs08iRKmohaMJ7N5DBV3RMLcCUymwnLwylm/X
cbZowSro5Qh9r9X/Hr9MKO97vjQ/r7vk7hSMVEMyPcyK+DJggGWuQyxyuamB
USuASQsQDFDtMJ2Rw76ckfPuZlQvslUpFGqqiw5KWljDC89Fb7TbWvA8dgQm
jiFbJQxH/DpaqTmfUUjue8lgUzNlEvKT4Mb/fOwDSWm+Ma3q9k5JE34+ck+b
fwbDGKsJV4r4+C2lojaxdm9qcdQODi27JG5U0kvfUx3QhpyheZX+1gkHnqEv
Ds53LNpbd69lkOpX36k9srTFXeaczAwcYPnQcEqjjp5t/ju8kOQU4pXog5HE
aRF8w09227LX9os6BW3QLfJ7scfFDzOaImMThK/EJO0rsnWTr8BDXHYSIwRt
0yxAl37sz2hGWT4Lo+qwLHmyhvj3vCtIzpV4erOoM1Nnw9RZ/7Lu916/0Yxr
fR5oeerM3W55I1qQOwWXc7k5Cor+aOR7nxCb2GMtnhNZxHXJXC5cRLaqOP3s
zqUm7WzRO1faRH4wSwnta+Tw3XwIkT0cLsE29vorN3snzd75fRXlV0OvsUOX
OuA1C1WO+3JIcs47pT2CjGXhyEXDvGNIM8LZFA4l7vUkHIut9JD8d88cHuqQ
Q7KGojMATqr9YRHkOS/fD/EBtEmyaezpoJ+5tKVnmeaazILjRvOIExHdUUZj
7PSslNfQ06x5qvoQZQGtm6VjCpDgFo6+v3UjK3siyD7qQ5PGm0Yv11mIwq0M
r7dvknkJv6VdtYtKn8uYr8ZNYmIU2t0IUq2zJkdN8btLL5rCr8qcd8C3Jr6X
OF9Iu0braS7YkiRql5UczqGAEvsie8WVoYR3QzSF9jYhg0Eow8JZ3vlJMgeX
uUp0yM6l9v0axsu/+F8UpavBbIz08k30QTVGG7gbWXsO6ABnztLkMXisWLoC
4wc5NLzwy2LhZIqv3HPEMA1pHqIrV5lR0I+yJGrjVOrRtqMdMNS1rh87kQ0T
Uf5BFHtECXb/hVptNs+Meoo981dI7+/V4spClG2bBCtrzf3hFTrhI5a3f/ff
cTzR6RIAo1S0jV1YvCx2yCFdhQ+EI6d1Lpl5cLxdm87O5cUL1MCgA8qezIAM
XY08HhKa8vFPC9Crr3WOH6+H9HAsxYwFI/0bjvlsZ6DlV2ow0oLMH3J+jHXA
1Ht4ZHLqKqFSEFt7gXyI+iVp77e/PfG7K+cwkbXAnHTvaF1Z4ecycP4j1clP
8YE0vM6dPTMJ7hScMISJ1X31LA/N+7gtOwhGdufLxNGjRinad7ukCwKrRvQ7
CUMRbCZSCA2atEcwC40g79r7DZ+UYMItZJGg0g5FpBKxBkXx6wr9a6OHuj8y
r+SgOcPLY45Y7L4jgGxOoVU8LfjxhMvXCDmFee9+HIdmUq28IrnFWRDs5qCp
FqWCJiOvMOPRwXauq5zSbEFoHL4HMpX8jrkirkrwNA3+2oDiFqZU8V2s8A84
SnH9aExLCJuE9NvTiGH6KMX08vdi/Bqvsuh51TtBFxUEqbWn/lfUnnbcBGKM
XiAufJBRxLpLoJcZ5Ma0Htr3Y0FbkDqHEO1hwRabHh2WW8kY+xoM3sbY4VDS
qrjaUyLqN0w3xfbS+BbdmVXWfvwm8f3NAlzQZHvYCZ9AxjBYYwpMjbuBDl9r
5LTriphnUnfzikDHAboaiYr9vww/RwuoJc+HTk5dVc4sdEe3qK7fTQ6UWBC9
bcn7sCak6LwZ8To6roBU+zqes2YHo6m+NBhGZNCi6mTOTTA/tL7IWL9vFG5U
1MxN1/Slf2qNZkziDMXGxnoeEc8m6+mg8wjUItB8kZcMQIDU02V1reCncqbu
PWtYtHtRxKypnd0/46MpJWDZX+od94kQHMy8obQLCA5rvyOjQEP2amDh+qfz
DDFWfCZRYjnvtf+MqKFhJ24cL898fG5CqXpbvMIX/MqwITDgS3I+2UnoTjb8
YflYQxWCWX/fZsriWP0EHS03xj+CXNKeovavZ7g6OmK320kV0l6LkeXmk/Ul
PzvijN09PREn91SMwrO8qK0AXb1KQNTyhBMBiyLQULGVbe9LlIw/IxR8WM0K
JNav9Uwae7WFwHCkI2GDHYyP+88wP5fAw2L+/QN5WZ4udH4csiYXxEaThSrC
kJLDLbPHyr3RYmctdl4XIjGTFF3ti3cokzddl6Wdmwu5pqDkHKMFB6R4ZiYZ
v+WBojmf7MapFIDXGVKEOspiRkF+t6eq7o1nMkHXpf+1UtF2hlOeP4t+DuPT
jMYz6J/tAsf+xnGmCtlu5Tk4FKeQr1nM+p6A2pUSYoBwoE1w1gdP+HHIiBKl
uK2yhb8EbzRHpO8gICiYN8Qa2TMFQRdhTM/IYVWB6+G/Dk7SEz5M/ZUMsCTs
xOcXsZ/651anQ8QEE8OUZWUxQIWq68TyqHGON4HGSlp3UoHI1fnplrWrmbbN
TM89541szkZczH9XlitUvXS6/JrIyiuCRq0IxzpD9wVN3me89jJN6D8zC3zI
9gL0oSXZC0Npg2l9R4JF7WMqmXjB7887IuLxFeR8FgZvHTUgTuf2YzCGpQ5O
7OjuhyrxGXWqt+K65IX2m3DIlzL5A4Mas/HYrkwFS+yrVr1sYf37ll6WLBpt
2RB4zTFM6Yt3bcuPZhA4enK5jJITOmzavrDS63gTOphL8oRyMSlDtiZAsNkz
BF1y+OnLfUYQsXigbgEzOQuYL9/Bd0RSxQlgHp8RXqp3DZeLYnYf+Xs4PGVT
NO7Hw45m/f2PkpqZBvXPFBBpcsNEVOu9dCfBYZqUgli2Gk28/MePQyQHUoLW
Fm85p59S7VyE3AL4WMk+WbRdtK+gpZYsJuZqyQlMYXvzB1sB6lPY2nuSWKDA
+NUYg5MLJpaCQLjQibaseiFS77cT3+2vxI5f1eCkNwhoDn4Yo//Txcp7q5ms
5YkOS0dtVIkH87zLWY0xOGmrPDI0ZJDOw+23LVeZjoFsI9a2R2v3WKe/9W4h
LyZX5dp/t2n20WNKw4/I0RZW+FV7//w5CxrpQIxIuLWkCbZytH9UxQq0MML9
PsZa3vp5SZFKuPQLdilWOTzcZ92A8+czsmM1Kx0/cpJPzwVcPxRsI+/s+oXb
3bEQSkDBVkO38QgX9aJk6MIeUCPkzcorz2AfdX56m5BcLrmh/pqZT0p4tFqq
oOw9g7FCg5V7cvYJkDbzyzwWGpbLkBzPgX2Z/w3NHHQv0ueDevJ5GreOMHBZ
/eobaTqVaSgZ3Su1Nou4Q+bMN1HmqcTy0WsbvDzHZiDojLJNImCF3MtueIvG
7UVbQHraYZgYPlKnDmMULJaLxY55xzendZcWAczR1AzR721BS7P3GlvIZkQ7
sb7vmj1diXDxoNKS4zFh/FBbelonEUFjl84FzqEwkUbsAOxojY2OsnOJGgKR
VwK21TXYQ9pcEfCnwnru8MHE5X9jJ+LwD3UHDC1/caILdNU8yvYtnihHHZfL
vTtBv+5patmpsgwKpmNWJ7wKIUwbPUpxAmznBS2WKqrpwGmCcqJ7kRiXfQEo
1R/1TliuM8npDNXyXLb77yLEzf1ufD4hwIJIU90pLgzPl/pwgsdTm92FX4AU
ADxhRPHUm1Ehn/S6LAb43QS32kJqc/3uA34gQYs2jVPdsZBM/8ZyEdarEhCk
dH4YjELJZBQaxX6OKgNUMBng7/oijxvkRR6aolER/cvRVwYNmejHQzkjw/Ob
vai05CViVjizDh3cHUmS0HqS1Ff7gCnKzjSL47L0ccvszPm0lrZv828VALDT
T7uS7va+BT4xDJsJPSN6V4gY4bTInhMqMXyMrkXAo1VsEp0OPV8KzQQa+wff
kYd8zd0bM0KHfo+JICerFbwHgiaUXjfxcNKqbTjCa3ArxKjhsonrC9A4nAPy
hTp7KMEyt5YM/rrXqtAzCav86X86FwjHbEM6m+j8SRc4aL9qHqyPO/miA7Bq
y8zGBLkFy9YmcSfeMxqeR3oQmW4RinSoDcNYUlJForc8GQQAP5Ge5OfW3B0c
EhlR4k0ncVf9Cm4Rh5ajawG8Y0nbEq4Q0Sq1CKmjm3U4DbtD2cAgWdwisLQx
mcsjbRlS6MZIC2M3u4BKL9APdaUTg194GXKaICmW/yWEIpSSWTSh2Z5rcI5W
ua13A/Rq4c1lZFrw6ox7KAw8Nb8NCojow6r2G6eUpBW89Yo+XdRPmEFnngUk
ewWHaLjyxr0/Cu/fmTmcHx7ztzjJc3lupeRYPcx8eDih3SGqs9dNPgBP97I6
iF9jH+3Ok2iyURDTk/Gif+TOxKwGAHKndaeRVp7p4F+iev+AD8bD7YxOcqod
1g8adXy/rwJIBzHXkWKic1fk/fAquvV6pK858HmqwZUtbQUm+XXbDp0MsMQt
jylq/GOTl9NhlWAB5nDBUqrABSxi3tGcuwYjLn94Ilp/z3lAxVmDGrbIyiSc
2tZWQ4bd2jBLYSrTXJ6ZL64cyO6lYSZWhsfDx0Slk2Ff4rWwp4dklW53Mtw2
FEF1h8i9Bl8mewLIW73BATbt1Y6JTeoQEP5RgrjMQVklA2Yn9CqCXZlOfhVk
o6C1F1dggaqCxFTbxM95uQI5mGZiw894fzolskBEbiC83A3ndmsy65Xybvvd
6RItCJlsgaCPtY8koCajWGD3gRvzeTIv1G87OPDJacjNsSruuEZrBpPWBdku
7+bSiZ2SE0sS9kW0/hSwmcoBc3YViW4B3vlwhIpzyVkOr0UR8kjt4+OLK+mk
ce2l8kd9xArx3rxM/zcsIO2tckE02F1ugdC/VMX/taOXBAj8rmT1oLULTYcp
MaPMitcuzr19zybQBUCkKAk0d2Kto2ExrkzVxg+3EhByPPVgIcwtY2v+obW7
I9eQSG9XQ3UTegr79yUIs8gO7+jSPJoVKoqvMv1MEon7WqKJMPY0USceWF4u
2eHlgZDUUQKEKJaZnoolvbJOrDYJhUz7/PKRn7ID/k674fvoVl9pG13/kdvc
ocLOt58KO/jGey5AeAF/lyBaZLax8x3/N45lcBlN+oJbgiOL/z4bwPin2Rgq
LITzbs3nv5cvl5CNxKpCUE3SkhhfC2VCN04LOzWEDpUoefdrRvk/2Yx8G1bi
dUilTryaybjs55sSEdhaceuUW1Suzu15tW5zDVhisA0yD2C6w5cYOWpDxKw4
tSbzq32dfWnbYOqukGkgKQaPXsLtLy5Kc0EELV39ljkTuAwhysf6ZA5jAYhT
eDDcfW7hb+ko8Gcom0kwHkfogPlHNGXx221SIBDVkhUvzSqGrMSlGvsm0VLq
Rb8IBMWjAs1hOesYEH3Edoo3anai+3LWB2HMQ15QWLznibcSe6rrIGYipifP
iPiRltB9jAbsJ62L7FU06nfwb0Hx9+Mzlg6/un22xXPsFPWR+Swwrti0KsqO
hUmlybAkOZafo9CzRo8VffybqMc54/eP9D76MzS6UJKKfQ9FN3GPcNXw9Yd1
FnBMD+aADyS0Rq0ar5bVaAoGWiyUeJSpETb0SJJKVLWIvbmd8iP+P6HNZnnf
eRRvtPcJp8C9G4/Hp9Yg0NF4yjpBknanJHPQKIiVBC2n6IGKrxDBf2SLcqHY
FLL7AAHxMxI1Q9lucCPT68wlJwmrE+46R2gwY0OnxQ5oudyLOweQtrMOysqD
JcS4G82YgaXRAYGKt3YLYa/nFU+Mf/+wg7UMXbtv5szJRCYEBb9uA5kqdLos
VzAN4sjy2M8ESVvh/2VVLgFfO32lCK+uT4INh8d1M8jxjCxSGdsEN8e5SiGc
ooeb0FYGRQbhvQ2l2etgF+Ho9whZ54J5fBBrt3Es2p1fkPgm51KTwXblGeeA
uZgzVPqiEaTdVyL8G10Q090P1K7YXevFYFBHUAKc3C6HBCHrDbpy5h9E8Bco
CI1ICxka9fDfUvOV+vATmp4It/s3+Q/gHpWg9UjM0nB0CCqEC+1bWCwu/fmr
AO+9ZgFiIr8pREzmnla/32t2URavWAgm5hAbtX2u05TWVHZX/VZE25ueaX6K
cn4qDoUVlL7Ewpo+4S49bzSxW9C3MnM3KGxbpBt4vngOUPbjKMOYDP+wv2YV
81vR6CZe+5+X1WO2e7Y8WhjZ8BlnYvzcHadKdjti0JamrRseBzV2lpmHHPQd
VdEXHbGb2VyPOfbaAPUNEBsrBfcaHJUhnFgXO5tVskVFcWW/jByeW5YsaUKH
siLP2SlBHxJlqrQi3/wvlOPJdrDTZn03TMCA1QtXMGlyWvbqOxNmkSNrTT4T
Dhlo9XgRUNPY/+hA0CbqAcok7/iD8ySFCiDbjTgRjCEHVsIr8zvdIEWumg+p
tJmeGeQJ4Ca1XKXNpOSUagKp+o24FzuMBcQbFEvGDakLNvnz1ratCUDjI8PO
WkfRHpYlV+pZTxxKmM/s5FtirfZgTjwFFJhLoZxpOnkN+EQAu+7lDMbqj1wk
uGZ8JG63zhWisyFOnIIyaS6YvYae8kCVQSWc2gao+6JSuKI1wM8hgzMIMT4/
AhkZ3m7X0+0aZ8WyundDcIM3xB4Q+kDX11dU5MvOY1Nu2sWwF/Rg8WUnChFW
bg8vObYo41nwF5Y+E4mvJMjPnFcnr1UP6fufyGGctLbt2dKmpNI7EeclRaLs
LZCJLvnbE95TNAjixxPQFDwwXfRNzmPp1NXWiXFxwljRgrCd/DClARuXtNX3
r7MRNRnY4CCY9MWh8wWByx7q5o3dZSPg7LIjU9qA3ldyZHbHLF7lddPCpbLy
tvFFtMSZI4zf10gq32iAEWYeRhMS2YfJADkVZ0guPQGsNywrQkeL7ytSiFqp
Y4a9/sjU2rDIoPZSoJmzui/Jq4/8jacJhU75zgTkvCOLOdUnIE6BVzF5abd0
PBXOC+lNGgn7olxVmtrmjcW6f8h1Dgy/S2QChKl7QQ+bRj9AQHKMO1MLM7+E
57jmRXsrOce4DcZUSUZL6vpSdmLPO3cVNaQ6slK+Om1xuVcbzh9kPoN2cpYT
ybrsDdR0HaTVVHDDr+NgxQMtzyGM0rP7ueNupeAz4ubSlnWEjBvmuiuIBV51
yWmpKFPdks8yS+M9m+LUVxDYtYCoGcgRAz/Dzc+eyirw6MZgq+TLbcUnVMxh
amro0FUHqt4Kb9XThvANPTXQHG1nWTUImrsQq5d3MOOQIoPvhhQEC8RMVjLr
OIFtSZ7iQCv++2iUSfcIJes/L6tY6FMJFcHuuP08cdMFQW0lfBt98Z2ATcok
nzo41UoDeI1xWU8i/8grUtfHuWvxRR/aw9OF4XLVgt/y6dvGr+AcccGE8CK6
PmCG/r1/j0aINvb4lKYoFy88Vh7Bj9/C2bnyC279TqmCFrNXQ2VgJ2Oyvc1i
Qj0e/CFmBtg8SfUeVQr8qeOVGXZALzGvA8SAVgDMQcr6IXAeuHaw1oGwImGh
M5ZymnueaZHygYo//2g2e51HWtNUS0kqr0vh/tFN/OxLLoWWuCG/WyUoqQvi
bROsUdbqDVHHVF0Wi3fuUttBunPupYFuOtJjiRXyw+FNzRcoc6+GDBX5RpyE
/5/JnQ8LXux679McfvHxqNHcOB6GBAbHjNdvN+OprqAtJe6mdPAcmspLfxNg
q/VZDPaXzLX4+byqyaCQwyaS0lRm4NwDNX8cXheUrJlBtE3xAEt8BxiWcQvT
g+o/Y7AR8mQIdZYqM7GGboDePwiIH3XRE7Az6MFP2cciNxFTe1j5zmdCuFnL
DJCsqxleFq45jsds0d5pdS3BZSG8A6HP75KCCwMWWHha8Fo7uKUcZl6njGnQ
vUn4ZLcUJpm4L2jgqJBoA2fHemT2B2ht5kOUPfyK0tQWZxz2VJchd2PeDyz0
gG/1mJZEr2VP6fEt5xNmd1vvhZTW7I0tfHMsorcqZYFTWIpDguwwmrv/v7kT
voSDngNHUXrorxNt1w66p53mvyJERAPM4QebrDtsvSA+0Ibrpwy1bZbgBJzB
ltjZEeidVg7pNw9/uLzospnjnkiCuE6azgcwRqr2PLh3F81PzGwUsUKk4Lae
EAVre6gKgfibNoPI6DZ1KSPGPvJ4s+qnMDk0MbIfH7OlQmwKF3aHnAKxeH1s
uG4B4zvURzHcQou7YLN9vZnozJVu1b8piv5xjAt6M1N5sDVJPlVcILi2VRCd
ExzApzc8L8Ed5HM/cGg1GGxkvIk6FvUCkWVwfdVZgvIUJciRf90icxFI0iFQ
Qs9u9RIgDgwXp/bAqbbj2P4oSR9Z07+/01DOsXbPGyaVoXd8LbyiOQ4qDUf6
U4eMrTiALVVUY7YpCSjj7QcANppe2Rv1uxSxVMpThXbJGebRMdlU4vDoYUl4
9CT5QIhRcRGME0sFp4E2pftK4d7kwJh+RNnE/+Yvnsw9/c3G7nnD3pKRGs6Q
aqfshlgUP2hz2U/XHeqfVaQ9Y5KQ0d4pm/+JEY8o53XAD6VJ2IBtVrDSLuW5
dw7NR9axQE38Hnwo9uCBjpJnjiM0OqUEbE99d09s1zOIaVJrlE12xDGj6HdI
NDZ2qSli27bR2twCtTG+qV3lE+vW/uCQk8/a+G61tcVTrBUVRh1j94xoCoiJ
56HclNpaePK+v1FxZDzc3EwCfrssqaOk+a+fPsywP+b2vZN8V2PMJbE2xFqV
51zAfl0ruvWQ0fEJkZymyWdsQXVH7uIHcvsFMqHCKdKfHtr0njA+Dljy1LbQ
DUG6RfVDft9Od2YOL2hPgpIpTKXYSdyVGvvTGBKKOWNIN6w7KG4qVsXbr4my
MvnKf6dTlzRB8FVcm5aiDrCkr+cIlZb7WyyLKYYXwDyFNhkey4kUQ6y3olKA
uffKUe+tWwkPwaPnyAsMSbnB6ZF7vi2iofhq+AodjpQORH9mJO2ML4qtcsdM
4nkpoZzfjKg7FQfD9HfQ//GU7ktvI9W2mrw2sTQ5ZeZw1jF0dRcHXFAB06d6
ZiaCcCiwHA6y5aE2e7HJbySZFOEfNj6l2hVkKeHSYOatyuEE9YBAuLEApu3e
3BzKUvVrzo5CqhsjqvdbG/EIqfRH1BqoI+eCRIqIKukXRyldfMjEHld/2+TO
daadgDFhI6oTVBu7Yb0CqHIXnyXJYyhhEBu6CCRL9XWQ94NfoL1P1v1ewDgE
eFVfzbzWwf6/iLyJZ7tQvYGBwhAaQHqNrB26KO+Wkb88jiB2oOw53merFFol
BbvutgopO1kW1HtyGAZeUw/xyMTqaO9t1wLBuqsAJ7I57kBbcCUz81UQFHyX
MbEj/p7ZTtEtRaaYQlPDpHzT5kaii1tSJQ1EeV+VlSMkfCXr5HJJaFpcXvoM
Gc3vPO2OXjfHpr2a88lLxaMu0dg5Pa+mNGTuCh74YQ5drgbunA+mlrDdo5Bv
SA1fVr6Z8uUSeuF1xAKJIwWrUC3hzoJ/6aki8lT8ANkBUDW8ruRh4MHz2gBL
ZALWzGH8cVwPZzBWpBfz3/H6U3JInIvxru9dyro8gmFgEjUOlvwZ/3S93eMe
drSMLSCPcKWlMFsFbHSKji6sQtT9bW/T63opmwHe+XdnxT+grwMGVVem/N2D
WQYC6CllLw/fOrb5T9Zg4HkZjHeFU/pyYqrCSK28wXPk3348uLHSOE7hHjZ/
eYmc4KRtNF6UtnqOe6gCAU/h4NyByIlaZOMQZmj6TMgyVTShsCqz1IUBqsQL
hzgsqgyQboA//puBS4uYS3QxRUVs2Rx1xZQ7DNO2Xk5EKrmqKBvBX7ko0f4e
woz3bKHJPKvimytE4CC5PPOdz3PCgpAjnZutzGCGsfcpoOxkx3QdWknVKX5q
bFpuoWOAmmJNGZWRR43DMYFs3xigv3T5tIYxaaLYfZ6tfV4zQJ7bozcKHFIA
pyhJJCfSYtE0xQnEyda2RkDDz+9v/LpPcaKdgkER2CDQ+6b0miM+gIy86NTC
GmBB+Ji3cLvLQNyPBSsPNozSe7C/nF5hjOXfr/AhbYCYPDool06hmsbCBAH5
GEcouTO+qzprxE9fSBLUeFUiTCxqhxgqyN2CZcGRF94g9q1j82kRccmdSI12
bB9cf1DdWQwOFS56LXtcg7ZL1XH4CjC89Ewe6NewriWRiR7uDweFJjz4mvse
jA5lT2j6EsPmnhrIlZxMgZvm9N7TPE3agfWTEL/L+BfMingHvpikiCQA81EU
9lTQcmr7CIzcj8hen4CB5E6lWQL+R1abTdE3E4+obBpBo1zrLtBcxW8tynh6
LTHprHlZvn2Kg6+3EbXiP1WWiE/nuuxrt7P+eNjYsnran2HfuLlnXjJlh0wU
7BKnHqYJa7Tys5GHvi1TMpzDrkZO8+HLtPWvjvm4qMHN7L9PM6HdjGjxP29b
OnlkrvnbET/s8CjwKHJZU85ymldE+loNBLHPwJMBgQbr27hCMQNSk/m9nrCy
Mnqoq/y6yrbvKvO+Z1d1wgLBCxg8EAs58ScWotWPFV/MmS3SY8HPxfUX5h11
ZBCJn1peyR+ljSZZUoJrjMmXltUUmtZlDFW68Hl5bk20FcMSHJcOrp0xVtrA
TyikYV9TfiuFtSixxQ8CnMxIrchpfbuTLAfNL8KizHRdLJ3WiDVbgF5bX5TM
e8Au9Th05L4qfKFC78b5NhKUZTcdrcIo4pOULMn+pI68kzh8S8Ti7yGoSP9A
JyOoz88lnoGfAh7LYOBRZZiR8V8hY+sWWBrixir6aM2IZf8F2Z4YkBT5+IVE
meb/yMEDJTiGJxPr7cZl4kusazu119REfq7ETX/lJV0baIJ85EBhf4YZ5LP6
F1GwXX68zswweG7SrbWmM29dxl8ttI93ikUysGaisJs5JhPquGiNREdEUd69
Ur67KnoJIQSsNxkRo2H9d24M+DT1IeE7R2t54yZwzXy5jZU+f1PX5aQE4fzo
h/ohc/OD6ophg3AcqrW3agM4e2OcrfwzQAtY7aq4AEnlwz1sYBJY5FkPRr54
zuRwfTmDDw0ts6y4NN+xEQkyW4AEQ0rZ97OtKW3yOVqCmOm5Gi5w6WyPuSlx
zYFn2pqFeRDfDsKQy9rBFKDv4nC8BdwKqogS05gdhN4vJHGLvaR6H2l6+x99
epSXo08VTA3qtB0e1ZL3R4E9PAkktc3qpcT230fLq7vmYDQGpbfFXZnJCVpe
iUX2EwDJfIp0E7uHwtkkOrKb1kK2xtyLojBdufpIvm8+Pz93Lxkoa6qeaU5R
0W0IU7uowGnrkA5wNtbRNSAHtYEq/YieIYM3x9+Xo5KEzOg2rMktwIK/u4cA
ezTi9GmT5dcoGuawo/+O36FJgH97MFNR8sg5bkila1w4no6Htb1kZ5tATeQp
u5wOq7RV0ihnHW8UddVqN+Uw6y3u/bNvHOmi6ewNXn1HeZkzPUuT/QKIlbiF
kAanczZ4xWCcLIV9QYRE3VkppY+DsfCtuAD8rqbxuV0iXu8xXNa8bQDOJ0jW
/2F196GSSRzcyxM3sLHTYMiI6Uxl7Ec6DEFZ0ywCzw4obIH04wsBWCDAp4wW
aQIw2Kn9k3qvgVikVEBjsY+SoL9lp30Gilah3woI/PcwsYK0pvshWhC66BM2
60GQkLSAMyj7ka4PL6a7BzqqhvHS0lZTQ5V5U/dmrqwr+Qecp+BV7ntFZRZ3
gkYt92Xlmd9Oh8nQ64KQ7lSd64M/E564zITqAPt1ySClAvYqFh+cP1304CBn
kRqlebWp0Bip021gOPry1PmY6W6V1KlUtnUsj5yzgrr2WnjrIDsAFgtMQdQT
FVLntIKm12d/rJRaJDAp+8K2LOciDcurOh8TQjuf04Vv638RMZ1VbaklOtQs
BlOPAvlw6PRL8kcKfgsW+p19+pewUxHte58q2voM0UG1wuRZBpeKXuFxA8x3
So7+Epg6w7twIEaul76r3c+qa49vQAlGXcRyjYSncJLIojOPno9SFRU+/01I
8AWImsX7VcI9lEuX3Nt1q3pv6VDRdPPjkqEgBbN6gouyOlzds83nM1h2nF++
VA8jNAKcIlNlODWY35P7C5wDG3ZTtSdZj+ZmhliWjDBzw9Rw9fNWBvB+aU8D
hGJRFJ75xRnIZPt6GHg5RU9YaC5tlpoTV/f/LkLnb8kplpVRAPgdL/+X3Pj4
JVV3bpSBWQJHdZi/YAFOlOMyMRgyuvPZ7D7bCqEm6dYCok75luIZeDTTjMH+
ZFa9DX96/Ne8NKXqYst61epQfl69qpH63dcz+CUYaOGIP/l0tpns29QejRpa
YJ2RkyujDZfw1WJ93eqyd767R8HjF5iEJ4DIXRBkzG7E60EwEX8UlNqc+GDK
L+l7jTqc3Fb6fed8SPXO6WAoGFpZlz7p+czsWuCkJVA3A/KrYYbRETj6EGSL
xZB2cCoQfRbLix3frStHQUVFJjF2zf7P7C9icZVYQRNjEWvH4H6QMH1CewyT
MnMTlB/nQC/C5xpz3Lk3m2R7W66SQ1ioieYEZovHhB+qDfM1L6XCIpO1C7wg
mnenAfweJ+7qCFW82zdcms4smOZyWnL8K+UnH7gFY1uodAerP3U4+zgp3maF
mMjceBkuR7HilUpBD9owoxqXpk5G5YpG52n6WJ8TjLPpujnDAlrvucRpoOZn
w4WSAf/OezC85tleoETs51aaHnU/zd7dfhbxkEdqy7vAAem9yieOXw59Grhd
NRsF9y08y+II9OBJIRUzgJxPc/EV2s9Zjb5aA8nS7PEaabjpv1gnhOprgkO0
rSaA3Qd6o1yklTSr3oBUHFJoZVPXk+bJ/DKxFjdxKeb7Ja4bk9raj68dGt9O
NJJzjRD4VERz4M7YAuoTG7LEdS1vp7K7SyMRMnj9qE9P1U8KjH7KHFhanZuw
E1NhNX8vNl3Z4yYwPibzA24Unq6VIw0Vtu4bn5IZCIyM3Dl/XYxKR4TrCQF3
vXrymRw4VAI6FEsAwL33RvbViRxBdomGxYL7nfWVBVY4q5zltxzLqtypUs4D
/CX3a4Kxty71Xl4qH8x3V+EHx+Bjl9sAZphq1p+ULO3npVy380B4zMmeJCBx
GtDyYBHnYpW8ARESnp6lTU3IlQdNW0GcX/xZQeUdRHh5SdtuUsOtLX88AYF8
TH19dUQt8EElBFn4eaOIusvC5dkqxOHtIBbe7g1An8xY8cSrfDfMd/RcoG/6
pb6Pk0ThmgcKtM2xylg+8iB3e/dGwepmPorv7122JCCoZNM9XjR2GqsQ/Rff
853vK+yEC2S4dpqgDIIOlIQ6CB9/SnckVmHuoIB1JckMNNhNX+wpBdC/72Iz
0dm5SjD94z1WCkxLiN+yADUdn85AKJWxTt11Ngc98IN//WYAqlMnH6PzK9kg
H7eUnWlw58XrdaGsBygbRuMyMEEzTywJ4HqehNdEFfv6NzPPybm+Y65d1ZPx
siq6eOKruns/v/VcUbIQcjyNyJBIVI/bOfK18zBOewwgPVAgvqeyE9H3Ue0m
Fc9ztr2MpTxR1yjASZRo7Opujtu1jbVm341DkFgY1qQ+SR1zDo85eBcJk6ad
Xdx/AB9nJ0n6Uaa09GD0m07qsGCmMwVJPkiE9B/QR6r+GYHC3+qXk1bvPuIa
rxZGG1gABF8AxUapqK8rwO8HuiNvQ606o/YSOP0WdJP4Njbnk4s5TL5Z2wNq
wocGZ9QzU2oxEIp3sgYyY97xQdux5KObP5OvT3NEI3xHCd06PPdWPw+7+Rrs
lzerbiaM74AbFpn/eAt3BL/vljQ/t7Ep5dJLf2Jcf+nkk3jjxmAkYu5BTLCu
t478RXssG7bBOgdf0mvnvQdie0CEhFCAtL5+ALmrYJxRLZAibj1H5u50r7s8
+l2koJAQdy2tDydWatpCZfvoN9M42SbCra0wtOWTDoVwNdMJqkyD+Q2eFsi7
GE8fPz1G1NZo8rarBnbjJV7JOa91Y6gjXP4/4ux4FrOIME95moZawsM7ZOHv
e6G47h3rCOuQhv/rlwnI+u9vq6wiuA7zNbdylKUztV1MV7Cgqi+lmDK1tyU=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1L6l5otvbStvUYK9pzh4LETXYnCbyTJZ6n4J+XQWs/eobg3l2gkV8OXGE8EaL7yQZFt4xdyoK1M4KEy3OLFZAigsnnNh5DDGE6P7+Qig9GW5K7hF9hx3WZzQiA378MF+Qs4Llng7GjvNzzTFdSF8l05If13kYU3uyEAyJDspFVEkpSs0QRdl9t0DufnDfYpDxDbUWWvCqrEjJSbA6H94+rDBhZx9Jcty0x6QfTAvN5AMVga1fXovU8QCOjbz52y4ypTDYfHUSPqOCIxzAg1ad56rDGMjDrH8grORDrYUtuKG5h5Uc8ftGaGuWaWf4IjKEdMtuq8W7Tx1mEbWDAkeUM+JzrkpfHHR7Y/vEvOzVZ6XSXhPHHHSQd///eG45aCoQqt2fE8lMI2VroDO1/qG57iRe7Zvu7qtIZ1wUkwXEftC6whf80kRo7FpneAEloFq2kJdeovtIN8qoORIq8fh4t5DeZR4RjUiinWLk5y/FRB3NTkCHLOemhELpKvTFW1kjgU4c1+cAVRFN6WY07bpi4EEeCRwmVwQCEe6RL+tX4BzivyrmYOEst+PRLi0aJGzDyu9LIoygMKT0Pid9NKBLGrksfTl6hJ9k47d30quzvwMAJX+8a2KbVxSqs+nQB81dx8QFdsjmrmRGkwFTxaHkmQUmOVfkMpyT2lcDRWujIE5vna63gE2CLxTCinF+Wp6JUjtkyPOPM8MHJDFLDafGLVt6CKzgww+JdInfPE2YjwT7JcmMcsboaxtOdIXQQo856Bl3MIHN25RkHB22qmyCJd"
`endif