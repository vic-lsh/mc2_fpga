// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B3y9XfQIKQ4vR/SmW60A0+SM8akM3oN9X6Pd40moyVuWy9su/7cR86qPABgE
qSvwX6vBskrvz7ROvJM5TpSuZApLLbRIYzLSmsMGAWdtmmWKu78sq5aztuxc
Xed0V4sgKeCCYgpiW55ga+w14wMM2sO6n0fFmQhkbYSGIW9ZsmsrJ44o0p9P
ZPSoOfqlA8uue2TQbJJZqnt37oP2+sBkuBJvOjItwOc2DNuxxdVFNM0jPvf9
O4Ua91ZiP3t3UPoXrg0TjQhfLN4veuIF8HH5TXGsqsgB40rlm3T5GQ1iEkBB
qWhflhljrq0pqDnM4HbYTDjWqIXRsJfvX/9jd6R2HA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cI5qa6teIEAh77BL+NXaGrKmvlKiiI6RoFRMg+KU+Al88FS9MXDgi8zRkguZ
w0ghCCtfwQoSWvcv5Tvu5S0C9z316o9RqCq14mGBIK6DoW7BLqqaUkwsMVff
jM5F9quDaK6NmsgxI4GG9iC3NaT9jOP4/z63Vwileek89J6QdqTwxbB8Pwmi
B/2bGhkktzAL/OucFLVjoEC5szGCSzBB9Ycvg6UuEH4GSrSJ4Pd8zkT0tbjM
9BKCgSyI9ewyefC4m7bmFhbsxwwOxwoFExpiomVUmpBVk8psKhvz6c2xOVjt
pipBurwH0uxOjN07Cu9MQvOeiujBCIX4su3T+EUTew==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ifx5sxJOz8lGuleXUpauugRUNRuHWBlzcGLml8bvtDF/IqcPigMX+f2p8401
bv70xdrXjNvOuzSpbLQB44JCxxB6AwlQozZefH4zp8rOaxNaja65seASTThQ
n0h/kvIAV8WaQEkScD9nvBfHM3s66ZI3iYuvSA+Y5YOYsOz3LdeZTL9KBvxS
iCqjyXGeMKCrU3wxyhKWLT+dh2KKfiI9/wl6DBvDKiy6pp3Yzob+stj0CzAW
C/4YBYp/5EYk/YENPhVhh0Ku0RDQW7PZenZPqtQJnm1dI8+wnj9zWqA6IqvA
t+UXJ7Dy1QIYJoJ29DKRcvVGnxscC6rNnfpHq0c+KA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IT3OyVLvsLrCP1wntlRTYfKsjxGbXuqNqG4i62pUNbH48eO+/7tpdbvgyC6d
7/rsMzcL5aQtLAaq9KsnKGyMKvJJAm0byFfrjIytZJYJamhwu7jYVNAP+g0F
5fWsGGA/BwELDqmi5MpyZpilHXGKahcugq6aRpm2D/gXPBIFzeTYUOqGdiOd
K5RA2bblzqWM9oKJCIp05slNwTnJymBViwt7+OsoZh3nx0GYLUnmJj9N5tX9
4b9/GUA0rf9n6mSuaUn4T6WKX+OKPhEcp/cLx8BU2nFKr2Q6DP2il8Dj5Rx+
hS9JzWL0qYxo0Q3MtuJhuW3QRzIhTWXo/lSy85TRSA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
abef0rVG8OlkztOsp9NKGvbuXSvUE+kwFw+KGsxvUjMew9AqpQ2NCz9ijuV3
7dkrnVnPMGM0dV3lF9QTVr8alLKWV5DcDZBwYWQGSaeftcg40cf4z/pm6Msu
DRJANsxAyZ1Aj2SZMYLfDTIEiosbXTrSTyVUnMb8TnXPplVjxTo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UweHRODFNk08QYVzUwczrUWF9DuXqi5DS05wxDVhPt1wc4a26q3AtZqGvQr8
oyt/NizV4ZYcAdZNTV3/8/ryAM/wnLMBr6DHSq2zKa4XbAwwTLfVP2VmrI96
/K2tDvz6WH9ogq+Xl5/wifTblAcYYTVz2be29HbP2iwWJq4AtwcEI2m+XuDW
xni4bmJeSyGpKs0y9dJnyb5sZJb34xkKGtVZVE9y8+QQWs7mwix/TVqvp9WA
hNe8KWiAA5sOCs/axQCsENjWAiAwzhVmyq6WK8p8gzRVaVilqp7+z9EN2qRe
n4HQvImOB618fvc/m0w5MoWMUM7dPDNbSZvs+vsbT25ML05QfJkARlvka76J
1rqSoR5xJ6THO5j9weXi3oQqA3vnt1KNFNst2PbG4S34L/MpzE0XsXWdfH+u
iK/pNC9Y83tABpKQUSob4pQAUpAzBKBq+vy469Q+ofqYVmRko08VHvT5/JQ5
p1a2iuLL0CMnaV74bJ1EvWC7uHSqKVpF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bkn5JUBhW11Ehlhdbi//1DREciIcLYZHjVYhE4H29nJSQZjbMfrsw8Z+Kq1S
kLQn49aWqcukee77SfQNAJ75X/bJHfG6M4kA4M2j0C0pcI5r8VCQjuqaqKrD
yO4pnabw6Efhaib0JVGwv6SuZV6CZkeuKLvxkmFmSHnAG2YVw8k=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d3pCWn7VdpPT2/4Cw3IMcZsu5k8Xl56omQ4Qsiv4Lqm4No3SyVlougz+Tlmx
xtJ/FOr2SR+IIpun7GT8JkW23SsluAly9kobGiri2TwkkqP4gtc6Torcw0hw
UX6UN19+u//YH/uZOC7F/ZuAiFOp2ICXoS/bdGP9YGqDxHzy1UU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13008)
`pragma protect data_block
qnbq/NbCIIWrrTSeIePTnJJW4erw4HzvDm4sc/BkK/0A+Z33DSNBwMtupvWa
UCrfjnfrK8Ag4ZLO3DQQWPnM8LkUF17ynT+6iwC/lckDJr+xDJ6s8zvJrXh0
KXo4rsh0OByodtTmmwafrIc6FErCTa1Es+H4LQggFQKQD7iVU62qy1QZzfn9
d/IAWiO1GswJXLzOC5L7GA1uK6Xcvih+MpNhkmbBbmh3d+JGm1m8gb2ULkrC
NZaQZ7WYRoFKO4hJj6G+VDLTIHjb1fHTGdmb777ZRLSvIYvlRLRLNT+E6kud
3BSsEiwWpoVRtu5m5U0BsGB0tHYxx0DKC/TbTzzLZDfg84l1BnfaD4CULAHF
37FkPr4i+2PXWneWkPvuWh26WXKer7CTNWiGXXxKEt9WnJTQvyY9YcoT399y
eLjrFXTXotBsc+ttqJ3bBUOM/Kqfc3OQYhjklSCrFR7SKwaF9543OKf7dq1B
s0BML6etb3lzDhnc3RE79UknT73QTyNMsQFLk7ffKdcoeJ5wuJPJWZdlV3sf
dWDB+KKFNTY1lKN/KYvascdzSoVL68H7t+qHoZsMA2+2boHI2vgqHoG1OwgS
wBmIDQvP/tEFQCLWmWkzEFIj+KeVkylJMBZnLct3PEqaPqaw5AgEwvQLFK62
cZvihHPlILa9wm86WNqsd1+gwdCHDym6IZP+LuzfpcfE5tKoUEuL68ey/K4W
Dh5pZk3Ef3rVO5eGiHtDIDXzjjwIBQUBJzvDQsmcC1DAGlcVGyxI4tKEY5ap
10PGO2yJmfafM3bIoXLx8UiD95k/3CRoM+m638hKThjeD+VZGus8bcWHqb4e
3bTXkO72RetAf6zfaZABuwAqIgQNcZXGeA/i9e6HYxbxhUx5r0169girU8Qr
uqgsimQAw6JQ4d17cOpW7dQcetFoavnvU2U/lswgUKJn0JQm+dvq8ml6o6CR
7fKvUjHMe/Srsxz2NbPxABj4Dtc9tBxFejzuOoa0ejlmNbgcAOU7x0ozUSfQ
NJmGPj7deWaOhu6S8pBkz04ts4OBSUnvY1eIA6HVluyto9KnQXuDHkQdD1h7
KT4C4PzdcYsPcngLXuQuS0ONf7UI0x82p/QwcyA3iHtbWj/VZVLyaqRYY/DW
YfKULmLSF56oq+4lU+rKTYtcgK01azIHHTJ9B+Wizh4EVE5qYO/r07A/nPX1
YyPrlerICgTWYMf51/Qc/SVBa25oa9Wc1QeL+lF+Pwbq0R63UZCtPnKDCckb
Bc6MnbuO7sCknaHWDyb0+ZemQCzCYBKhB61ZbJldhAvNVHz7zK36FwiQU/e6
dLZoz21ZGY9Cb3AXMVA17tiUGRcwphT92k8D/TYBDpZxFKSsTdIZWf/fgC8P
+et6OFlyruktbOXpEP7dlzkR75HEEYJ9E+MJGKVszgPaptKR6OJ9yX9fFsZz
0O2IOpcYcj0drYm0uO3j9Fx2/aSfxmORHOain1Q2R7p3/EaaSlu+ijzqPx53
Jt8Ys4kG6iHK7DokzSQBhGoF1xH7In5Z0B5XU25BbTGXJDzDFu/kdE8+RUtY
k43OKlI2f0rHHwWEyZr/AC0BEPy7R53wgzROxVCxYDYEX+Ku75sv168r97TU
19Q6HY5fgBkMbQUBRQMmJrP4NGLeYVYYT+rQGU+JKkBAnF+6keU1+c4uJ+35
KEie8N/sH8FyLP0VWcQHoUXBhIEurCf/LOxxW04WPR3qlMNcwTNob/f39NXi
7iyRuzzzpA5qjjZqE6l6T6oTDEBVgshVFJ4Wl55Ru6v4Xu1c/SJGfWK6kInS
lnv6d2/K9ZYwKoDouGjr79/8rpZUCCPJKHJUX4rtsUw7/kZ9AELm90RCTwLS
lesSL0D5OoZ12mViFLXrnLIHHb2eTy8SeZtznf9JyPkeAlxx+ueCTo68JO+2
/01aVAUDwle4WWLaaiEGmSf9vocOIy0EZDTbGmAEaFzPe9I33coqnoTEQ+mn
+tJV2dyavOE5JaDdclXWerctLuxCyd5irV6Pe1PKwu1aTbLlfBmOO31j7neI
23KXC+8kKI/0SrxNx/+HrkHlrjFRBUndkn6VKasgmdX9BI6s0ds3LS86hcEt
F5zUsWfFjhuvSEFoAcbdQkzAlHRxbLVHsCoELlzVypU8FrMl1Fv+pEYUZQ6f
mBo3d7dU2cVvKPdqXU594AB7ZMe85EieaL7cZ6k80Reqagwxo09GfCdggyVB
tDx3ywFvNG0DJn4o4tPSnR+2vW+Qb6mM8fs423OnjpkNDNhbTD68i7P46ToJ
OfFH+QAJcbOkcblpEnVqusrJIF2EYYxjr2TeROx2shwWlt6Q1YtHFiDuaZ6e
tWPMwURi4OkSys3os5zNu8Xpy++itZokFaAjlxzyiYhQQ6r1Jbp2G1I76V/u
ffbx7J5GIr4DgVnR5jUYcAeoyQAFaeZurv5YKXs+2qUEqmBskmwaecJhq84M
R9REFhYD1JAiEqSFzjI/P6sAQgMmYqkWqsSStepWBWGj+dwT497Dg4FkPtf0
RjKKtaOO27nmLcXiW5/V/NtNVpxsYrQ7j/AefiI87/OTUTzWHBmkFDJCh9sy
0IDsPR53f2tlzEHz6b6cTPpipBKd0qUXdXrQg49FCFzu2EEClJky0LSiFPzM
9vPdCrDtdlGIQOW49fz07xx+IPxTFNUGcKlkMIfV5+q7gK4BioxqUPf9NFLQ
uZfbwN3hKQdC1czK9F8rsAVCfW008B6Dxj0+tjL1/s1Yjsp04ZZlFzf3PxfF
6CrXlaC4uJsFCIlZCYj0fPOuzi0k+VcZ1ESWSYv9L8LIdCsvgwvzu07jk4+v
/aMV/64zFRsJxv95Z5cp4aJM6WlV/dRjHUidCJM2u6VoyBlvs+VwkwLbLxK8
JHUpIvs4OWpvAkh2FbNrS8AKlj9nDDBvYcn2wqm/yunElm6VHsXON3m1ILSO
u53J0kz0A1IY/08m13A2dvTgSNwvbqnG1ciDbQ1v7jIOpUGaKYx5vInBluK/
TjWx5E3TydLFJ9HFW6Mh4nuNfmFKYOmc8Vg5rr/SDAm1P0QQ8PRe3UmtXWCF
8DFN5vUH2JAIK1QknIYswQzs+xpb1T0y6DjV0gKSqrqFBGghghfsvQ4ZGapl
YK0uHEkoOqivFUSQmnDcboBGoPyR/TFgNRe8+rjEtqw9GCHDGvL3vVVHWVAt
8Hfg8T2Luwd4NGyN6ytjd4UlC/56rrKxL89qnjFmjoXkqHj06mExFaff6MIg
wqeaQFAXAX/j3qbfEF2hfARhKKkanmCI522eKngei6yHIpyTUet705AjxaUe
uUbSYFpFd6eYLNQIbgEJjEz6J3JcWAhYxIX+9MXnI/QM7v0jcgIMBTM2MOrk
RwM45f/gKG1u4CzrAhAm6eVUgiXPbXezv9DcTIrVfFKRjJsKyr5Sxh5FORXh
31q2Svsj7yTagAb5IBy71K48rxKeGqj+5q34b6aY5mWo0YFHcbRJeWHHGzbd
LzYbeJ+tme3NaoDxplfepriMoiVizNOK89dFyez+eo2PNxIyq55KU3Sm4hoM
JIduv03FEnWN2j+Gx2P54GfDknXd1vVoyVSgpxU85UXuiEBXoTGVWeMcg9N7
TXw/4ZZKaCl5/1YFkcX2c9I8F6lyQdf73/6DEVGHMXkksZlJBLGElhU1NqDc
BCPMzbetNx+AaiJKTII5tI1Kz3ROLaFmZKRjOmHlKsy0R31Ec4kSrvtjrArJ
rIzM7BRpsL8KFZzcScPb0lVlttpZXRB/18m8hvMJK1VDkof66HvKnSBe4zxg
N3memkz2xb77fHDXm7GGerQV6xIPse18cnYfZXIMcrLuMuCv7aIYM6hdhgXw
TCG+bw2Ap/7VD5UlMSgM2ceWmS9RCe9UhsSVR+FgM2NIyIGAzPbiLyBwIN25
TtgGaQfzehMZ3yF5m08h8d0JsH+FJFkcy1U3kN8BydDOuU6V3/Y7P2g/qagW
8tD/4x5IWlGJcSorabQxImSRxKO6H9l0+qmlmHkYehpiaJLFrEPHazRdi2W0
VioWpP9T43wKhL59CVsy9BtzuQALO6h/+JSHiTQei8XVjbrKuxNiGYPS+2RA
XlvjEkzfRVx89f2g0C3w3rpJuPRXo72H56O5qz/RQ8OnWUxnCB8gUysKhevj
G/HtuQGxl+MaJcBUbwEFZIU/187Bk6N/k6kwTYwZMGU940Z6RaTjA8uAg2aH
F0rtv8uZHVOWL8B0Fn5Ywzx+UFT/Hyk45DhwlpwfogZF37SCjzMVgJZXNfp6
Q5qQ7uwfqvd12M5A2tWveYbDTq7E1sI/preLFrs1zqvfGpuFzRxvWwoNyNSx
d4qt2p2Rkl9JJlQxTdfuDzg1m/Q6biDd0GSP77+/dBcAAJpIoHsZCZ1bzlvH
rPT0guMh2tCERXdQGM6OTPnTOxYvhOBXZEHfUe0y4ZVWaDxutiQhOH8Bk4Km
j4f7XxDrH4T9x23hz2TKzuH3WmbyNpkX2WaRKV95WmstQnBN7qMcx0v506pG
Oxsz7QZRsK3eOFfw1yK9+V7hyUAxKU72FcFkJQLVLT+C/KJEcOdmRnQKQUIG
K96lM3n0sGrYw3XLSOAyoMwr+joesuymD1QaMirBUh/NXCmotrsxbCL4knK1
dNsiwSqP5Nr3uoPWpXOY5CvSFR8IUXNAlIuJBmn3FCHlQAQ7ir+DN4KjgXNr
O5lDe6PnO2bg8z7O+lYGp9Hx7E1AvJcLMehQ8Nk9/ppGk9AvUlU1+Gjc2R07
25cgz41VTd7nkkl1n8KiUPcLeFTj7kWgN/tEbkfZFpfuAcARLo4hOr49E5VP
YcltGb+MUvAisOvpyIU+oLACaUAbuXdxtHCmqMh/DB7IzrmITN/0wLANgcm9
NrQVeqoJvnPofw+NIsxqdo3ois3l6omASP8Q5yreRmr9qWHbD9YBRxXAy3aO
lf6eTPa86X/DVL+Mr+HI66DznAagaoyEqtV3cplULM84B6rTm1xi7Z/Sn7sr
lf+BRaTFs2u7a64FE+ZpChPM51VkqiziM4z8LW2wj4Ybdf3CmZiMN+7K4OZr
c8ltLOrYGN3n/65GSg8LxzlgD1kWIxKaKIlgScefFm0TEywOObpJ/a2RIZ6x
rkbDsadkbjnoQ6UfWpEm16AEgeU1umQkn2ZdeQhxZMocdSZKCZsLtAJ2Ak2B
ZTugPQk+AKlzG4h/9YoolQO2zpSmdNYmN7QIomno2c1udzNwbZNXLTZQ+bLE
aTE6udiqGrns7TH+hG7QG+Dt+542FDBzlNXIwaGra3lDIV+912O9pQvvrVyJ
CUCQC/v8eA2rS26nIYzLOp92X6MwxkpGWz+E6L2PEIHqUAMIdz0dRctkRgc2
a/06X+BNIH+KzOKvrEGdOFQN/vVbbp+4AUOGleVrz9+RJBPvFZxnzDYOa0Jn
TgA+nZ+PghjvmAXUIoMqbUDB3LlsoOpVlnZWj+3VsXHi6/tc3Ulck8ej0EVz
nH9kUrnkmLQHKRHNvKCN4TwRu7IUCNAVPCneGAJHhhX4DOqdiVQhplA23/MI
H1qZRuXkpucBCuoNyXBbSx86kdc0Fo6tifUBq0b093jxEoBkRX+uklSVVUun
4quAUbhDAs4lbSNIF/BFD/6VeAFgbrhIypJy6ce1wHQAqhrQp7FAHfk1iP1P
fFHhJNpTa/YHHcJKDEFnzlTjego6y416E4BikAI/lqnA7Z0cs8EFDIwNjuYM
spNP2dX0zVtdp63xf4d/GKwHj2um8J6aThzZgmN9XvAGWqiNa6piXpVWoU5h
o4XYaAlUt785d8KDldMiadGmAcz55nxzoQqhjxYRMRrQIcF4KbFr+lu4Rkgo
rEdwYgGxHGirBFLXxQc7flecm5+PVm6uBp7V/4G6FkB/95TZoaoSzaRjwgSv
UUjrrFxUhtK3jfYUCWZLr0y7XKx3xgsj4y3qYGF3xmGMUZjuCSfJlsjgZPGk
z9A9RvPhjIUyRORmOtGqPi0xavGpCRg4ljJsVCfQ5Pd5PDXUuLNyBLaw7uhi
SoLIPWEMDsMdQsWxL3UUaUmwS9Mq33KURHI92aSdb4n3YSScRFuTYkBiyBop
kskY9WwJifkoh0E/+bEUhdFCqBlQBqhvU4n5FwUvDRHwuQxHHqqbYM79S1fB
0KttzxenPzfLrAV/Fb5g1p1uMOE1T366m5q8rvBiDHN2Zq3mGH47FnaqQPy3
eJHsVr/4v5mNu/Cd5vnZR4R+NPLzED1b3Z66lQB07ZWCi5n2RC6IZHLdtqBT
EXlZaLhyGQRi3TJqEMI2nmaexh6296AW8WqNMmPTZ8j9YjX/NdbUq386R/Wc
PkcNa5RYCgUal2+lEA87/7RS9bRP+zIcu5srw7vgIpgKh/mhJ3JPnb3w79Sl
ibpbxw+BoMMKB+h/Lg5SfMhsg6VFeMx7F2HaDNQnAdUwOD0/dcDIWrx7nZFd
k60AUSBKwFZcISiZ8l9GpeEs/oGDzJyw/x49D2dwxysRbqUzt3XiOIbRbycw
oDfzta4PyuBsgGk5zysFiKeCbSzK2M2+JHyqkgNHLbLSfGe8unmM2wzjqpK4
lQ1qJ9gBKbboR6iQjXgGwdJzhG1GT6NP4RtJdMCC1aOYCo3IAtN3Fc7zuX3n
IUfTpvfOW3783AneITaAB0EQQK3UPylEXiasWu16aBc94ELq2EIdjaFYDHRk
XCxeGvVeRyKijlYqzbHcYBKCVpaHSTFIiqd8UGROmwJmdIOFDhQ+A4BYx1ph
+TzNXVxwRUr/5Scok3uVQLAfjZeq+LxpEb3iHtYxmZPOXYDxs8jVPKQaPbHm
Tv/fkdEbEMr0pRw98IVPIjyyP6GDjJRT4roAQojw/CnpXy1J368TqS/49noy
bNyHZqf9cXzq+k+asN8x/gJRbg7pv4gobaPThjVMuij/9B5SzUEhCx04Juq3
2T5U5dkay/cr4mPOiacduxN3JPhsBoNzh+FWpPIWofUd/ARGF1ELXE+0g/jl
3aExxKFLqU1GLllEVe0gTiJthIAPds1s/shBSxlNDnAmdxdVGewsjPWItI19
ccjjnbYu0/ztCPXqPOr+l/bRN322dVJqjywZizIWfFv8UV1e8DGtLUr+9/hN
DxOWLYJR6QSide3p4jXtlfGZ6zbZbBhSY2w4A4bMEIYwMw+9N89f13DUhEya
13v9qX6K29QSk84b9CzKCfVtkHV+/bu2Jk77148q5a/X3w4tjtYMJh9g4GBQ
N28L0QaiCihzWAsYYsgQxhKu0dQHF5Fhf1bxU+wUXrHypbgjx+8+K8sGcnhS
UMSkVyw+4QSLkQA36ckDei0DNBFesotZYVWrcsWLKqKjVAs6CC6cXQVA27HB
v60ZuFtqel5QkXtVGH0K+ag+y+vfB+d7ApBkaMRFv5LROnn29SPzm+KSD4Mr
72YDwhMpIX3DA8LSPwtmEi2wp9sRJpbWP/5RyLpKHsBRma4dxFq5l8VS+LXq
m/bKsPk19IbsxeAOXy/84YS4NuC/fl/pxDX7CnYU0fvMROsv/OasOiI2/BeP
DRlh1uMtoPoqnuI3lJv0Yh0SNJTyqVNrblMMsFnQk975nh9KLgJidqSNX25j
SXRGo/n8OUo2cX6/+aW26isOcZAIReXKzDh9GPoiekK3ux3bBLCET+2DUMih
En2wzKP/EoxcGty/zWE89RHK60NUCdpXQicLCCACcZDM4cqUa2j+jhrZlZ5d
vL0SWm2Mt1kPRqtj0JFTVfwl7YTKDKu3R17edErVrhqR5lUUkmuPyMhj+09U
2AN4QcIl2hGsTJ2571E35KnWomWUPYbBUbLYrLa26h0ZWwe48QcBSf94P/fw
hV8hGK7RdfSIZL+3chq5ABFFY5x376FOY1w1O4tfCmMnTCFzizKbRcUmNhP4
vDwmAUQOLlYdih3GEvQc4aH+FwCUlIwuaQ751utGg88OruTjUvWsuDXJqdb+
Kf0yRSfrZX0Wm6V/ttQHC1oUPj8ABWOiqBgjDYm1ml2080nI/UznAMvxvnwE
B4v4AlOBXTyMoiyRlA7hGwYNN+xXnHoLORlZoJqid2F385ziDkMxhE3A5twe
DANp0TB6djxzhe17lXaXP0qT5NZdFgS3ErRScqUJgHzBM7GE/NCend2SMb7O
7L/bBMsNoVnfpN/Uge3PzhVAPEPvIXnatxzDyLfa5HJScIbD8+5gINxrT7P5
H3keCBa/RN5zJlmmkncod+9UCMuTmT122DOA4+EkXbo7jk/iyiDQpGF1KA6u
gR8ISb0JMWKMhhPBp5XpAJK/ashyv7+I9kAtv/sXlJTX8z7/PzR4Ylv4LXzu
hi+L7JwM4JfnnCq4G41qgI46TfQTJ9qpxtR1FGeFulBhaFUxtq5oV5vjwzT3
fV2RHRWHwGMXaa/JY1/Ch8obChHfn7iWuxZGlH3/Pb3ErWmmIdjyIafdTwdB
6ncpgC3TwxWJ46tgDYiW74bzIRiAgRN7Rl2jFRwdSFgkP3ML/YcwHdbVTp+Z
plax+4hLORqWi9OpSUs13crbWUoIKtEuhPFIUje1LmXtCsDrnImwFcGdIMa1
8wSDxEUWMznQ9onU0lM3zZ2Wy+32rXv0fUT1KpARkNo9eUq0+7lvPBLtUIU9
CPoI0fTq4oD9/r3TOLKCWlszLefuZ6XtJY+CLfCbLwmQVD/b3RGfmLrLbhlI
2Q4QlL9dkP3vqrcujPyiZMS3aztvMb3tWFc89wdE+Ho1GTrEjmorv1oz/T+J
XBtedlOTOyHx4AXHYcIAFoZEVNSlW3D3I8t+btKi6oQtrEzhE3A8jUdaeGv0
oAIlLEm/4lEgePfIfpsnZw1g0JHvJbKWs7LCFYoUCz5ANBMG9mIGP1Lb9O6T
druIwP+fUjoBVU66nrwcLgGzidyOzOV2ASyYbkfQmp3YuH3tnG8s4tlilKGi
P8TVMLMhUh/xtIDBuaI0IHk+t5I5tBjnOwsPhXfjshXxKSTyb3vzPZmf/IMk
fBXGACNGuBMn0OKeLV5ZzVe36tB6SmYeqEHMXiuL+aVFL1P7HH2lawFnpsQG
kOLSljtIZ2jXVvDnKwOpkqNn4vcxvt8ZpGoc1mnV2q0g3Cp5y/sJ7rfoabJW
YeL0Tnb6Nk1uU9sNBODgGp+0bIYil8u+VOP/15b8q3zEp0ptE1/6Z9Mkv2zz
aciXSAyTmts4LVHRLOiq3WE9FvUsA2h0ZWpxwa7v+3JwoC5XisYMcc85kb0E
44IX4ZjHfx5wnrdBJ1sHp5cvySQ1Isn/4IQwvSJV6g8isNZkrV/Hm+cDqzX7
41cJNifRB4Za9ZLiLvrOU2j06U/kpe9rdsVwYlC8ZPAsM9MqBFtXgiLqahTj
jnkI2X4HjaGOxhY/CVMKYthMRMnVELCWFd4I75WxcklBsvc76x+xC9mhUOqF
Jx15znZ9d/Hjbb+R1B/Iuq7EpKl0NjfRQdzNLLWyugx3NrqV7y79RRMS3R+f
H3Y3xboB8pWAjjs/JZmcoDmTMXNpzxsjitUSUasY81xyoo6infiwnz0AktEK
hJM8wI3ZiVJrcHqlNkWMop4imLOk5CRKIeOi91rX183AZnJkRbaSdyPXF4FH
c0USno9vUy9YH1XmTuQsNF2vjVH0EfVrZXr8TaRFw1vYFVOM6ALfCgtBmS6r
8glmoaWcEWXRzbFcVx+77Gy2A9oHFSn4uxQzbvNjg2XYBazRfOJhd/p5ZI+B
r6wMG73neAMLZ2GXMbxPo1yVXLUdP6gGuWDzPSiopfVmWRxf5bB1vks4Xh8G
opdgsf0E0LtjSi6LnS3v6x5BDYxi/0Wn/j91yciWARMBeGNLEw2q6BSyPrGZ
TSFFoZ1pfumKVNdMkcU1hJ1Tof9FGxfwWwV+tOzi7vkfpaLeMLBZOV8zvMss
ZK5HNjarP0YI/iX/RqmlAdJNLtVm99MNmZenR88CH3AYZrppViNZ2Y5Y8FhJ
el+Vf3XQXCLkUZX1GkyTvAHEGEVJdGoPOoaV6VK6WeghxwkuhDAE5+hsWI1C
4c0orjaWeUbRDwx311I0KSPQ6wbOT+qtVIpniICNe/Y6dMRUiW+0rwPhWF0j
oLElrbsJHApt8lEQwqeplx8vgfqXYKBy6cG/zelLrzejam3pVYMd2YO3SKGZ
XvrKBs68mtVBQi9Z0FRzoxMJlLuyDq3TtlZNHVy96ivnVwKbOvSwXSyeEDpm
GLubWCCrwPE5ER7fZBb1II9RWTbwMItnXmu6QpqRr3izYeyyyQS4TwHspKIj
BQzbXEnzkTWFZ9VHwIj6lMQeB4FenBoUPWfkAiJt5cSTyTo9NyvQ+kpbWRoq
M+81Px9+ObxIx2805dz2EmuvBe1Y5geXmx1DrAGXMRsrQ1JrWJ6JaW7O06hy
SULj9z8A+dDIZ2wTUu8ROvzY3GZ5oLPqa4u7KQ5Vl+R0rFon/I81UpK7I7ZT
IWTDZMtdI0+QDSDECl0TeWfszybRLzwGt8inVsx7ZDRWa2qquhIgDenVF2Np
pUEivjF4BSRjc+CSklcvo2VVOLslx2bQ34sxegPJHajfr2pTD2EPXOKo4zfu
JOzob3r059uJn3WiXh2cFZmFTR7bB9zL1tRue/xFnzKUmiNlQRxMZqB0nysc
vW/677j9lG1FXELld0F494+K5YbQGvN538IX+C3LKLp8kGlthITxW9SCW8az
bXsXtzLVEHQ0kqBuGQZibEcgHE1jpu45XPT2vEhhvi5W9k9+0ojC2Ioh6pnj
7yGhI9oAYhacdNWepPE+YtSH+AYtDPmCBRB4QA6e8LZ7LTtpe99vcWQO0wZw
p4b4vdyHzfOeM1Nl5iVbV9tmsXOKtR/PErHxcv97h5mbFy/4VOGXIDGzqyE0
NIgMfXh9fkUpcbOqq2va1UCSr1w/yWukOs0tWDtfyzJW4I8Qb8qnQlevmi71
cyDkaDVTyro2VVokdjwciApgpif1JWupwgVTgiAUzjFyDbgl8APl0Utgl6+6
kAApQ/LHBg8YY2LAows5GJT0jwLj8saN3vbClqAjHZ137yGLI4tHNnUSBWtN
04Ue7df2cbGxLu8ttJDvZQT+H6lmsm3wTewe798SGaYK77nqeGtWsEjelGNE
ppVf4WrKoAzswzJS1AXJEZwuSnwY0kpYOsR5KLhlJDAi21KfwkjJoGnYnyKP
wBN38rrKifQ7buwhsxCQY3nNUgX1Oqbd7olIxADetzy+++L4mmvFasGMzOCA
BDyns0+cDxsPdN/SRLtgkpbg0AdtY24qHJPiz+i9W0V3PTGeEHpfsB45Uaw+
Mrd7c0eZnejDlpXA1WtzJPhuJYWEebG4aVFOglv8PZTnlzW/ew4bPoE9fuY5
OpIGueqHZ/b2krphoEeST93VxsoYOxT1+a8DC7TxDpQmJ+XUCifK4lu9wXNF
hGW7V3Ek5tyl4jhYHn8dqB6/w/KR1Y5Wn1/WNgCV8l2YSFFlr1x9/Iqa0Fhj
E4B2cdzL5N3zMNg4QASp1sxRl8C2u+v8vtysjlrlw9NYcYTJFHlkw3LoN7zd
vzR3OTM1k3YCpbIQzttj+dsLG1LYTwEAzMAxAuCKSiWvgwnN/xQ/b9KwyQF6
rkmNlOjRyct6s+1debjU0P73iENAtMjNUc/kgbHZKd/1hTo4HG6OJcGrDsf2
1YunJNcgGBPmgGdII8sV2djQjwDKOZzDja8iXTJ8qVAweaC843IFlaZdlKZj
5r3aydeW21esUA2hSFzxTPAcodNEzxv2tGfa16UDwd08A4q9xQv/Ixtttjod
hIrz1VUW2AGtoVE5yQOeZSKJtqPE1d8NJTdfMszydI+hytSBaNOibcgHj0WF
Zzhw2PcAjqBuTlaNx3U0vx6e/vGOM7MgiMNgyh1uIkHqjj0dZAJvMzgWm61m
JV7bCtM+a66XQOsc7OK+GErojXvkTd/7TSBXBV8HC2fqUhNOWQHA5AgvhZng
zIYm3HBT226M/6nBKBosxWZkK96Wp0oyWO3uYMVQM3lx6l1eGS463AoYYqtJ
6yXqyWy7UNbW8k8iHD0kpQdOk2XsTqR+CRxoczPf6kdkv07Edd72ytmPLZT2
8LarLSApPDaKrGHwo/uTnob1EjlMPYnyNqBaO7YHnv9+jBaab7Yyoi/AD3tm
NM+nzjkn4oo98KN24TCqYh1GeaEv/mPjlLplDtxHmXLg4+Of9HnxjoHeti5o
S2vjHvUZ1+605PDnoIh3pJnl7YxtctAIUy22/7NinoNNMxIae6jJdS4ZHSwb
iPXbZMQMiPb2ib+ALkDv1cCPz6MQ5V14HD9TANbGhjtm0vU58IbBVnOgmPXH
F2afA98pWm7YlD3CohjYNUWdtRPAMLQskygFSpH4vCQEPXt5dYNcFvIAu0gd
pas6SIxsm2R360otN6oQfAjb+Jy4jf1X4yped7hlsrsgGALNsVoT/zoOB7yr
84dCH1ObXB2IbxKZciWFH7PrBCqYBJ/kp8V3yVWTX2p1fOlxbWL1pVUwmxWX
4YilLS9Tp6EzznWhheInr8O3kDkN2NzJgZTOfIKU0iJVZtno/AuCVhJQinyD
4kxQwoaCYjzp2X06tys2TXhtbaN0YxKQT6PXqMrONUgkjdL3t7y+N60l85/N
cEdu+Ndy8sKuoN/q8d9ul/4UTMwEh4kL0rljXVABdYuELu3J3nBR+FcuOc/g
IfAakyKN9Jvg5+8Jp48UaJAFeJjTVBy+zWVE/QNDsdVLJ0nwuRHrI6Asl9m2
DibPk2TyDUuuq1YJnnRxjFpvqOjUnihaLkRJ6wWRpHRcu7UsTwjGTklNJCDR
Eb9yYZ9KXbgbYmjrZIeMKJvoRYeWQWhpYpLFiLwRquofoS8d0Nb/UoERR4sA
Izvu5xDKmk1ca4qDM1RQEMv/FnXb03jxiz9eghX0qufaLMWioZfWOTVDkH7p
zHu2gwOGpgjyoLCyqkhJACp32ZbikU6MMPj9ONI10COUNi6Srgu0tBmbf2WP
16sn5YgXfKomUWLKHBgEaicEgd9ZQk4p4qq8+LOGXIfufE9KJUzVA0ju/QfV
F3SeT9o+nzfbPBL/i0BrDKgPOdvwTqO3/oL2g6meG/tRyRqCiz3BqYKXNXvj
NybnHBonEp7yrac2VkXu/6BEEWoWFyo+2Sa608teu169ZtYvdLQgNd0AL00t
77e2oXH+037xtYpjT3gT/hVbJLPO0N1VnISwotMAfd/vdiwtR0KH4vh8g/cz
RuWoLzvL3XJyTCG9bGXUX7w0bjTBrFJN7fGTHC6qysYYzah8MsqhnUpcbHaJ
SzmGMk042lnL21pU8D2FcMOpL8JWLP5kIC8e8HV+3z09IFOGAEPkzZkEtSMt
3qZIBUQE4KKNMJnIv2/aCrH76j0TjHJLzNRMF2s9CstFbm+RvZDkB8xdziDJ
glk8xNhxMGGBURVHHZG3+0OUW9e5cUSKy9e98EtIib1+ipvAUUWFuljLenoJ
tQVBwGQf1HaPMBZPY/iDkqlbmYECgDsH+6UXX4+TlrBdIy1u+UTlRbdnR4F+
X//P0RoXZUt0GMhC2OzGKa0Ko4NqOUaSHUaAPzVpdYmKnFuY5mPSwWP6eGQK
6jU+JpV1DTe189W5L6reqOzLv22Yk34IjYPpTS0QPg/SnTGMd3otntprE+Ka
2dW9HLkjYWNYfDf001GSHMI8Zj1tEMxcw5l07Ss2sVlD+Bkw4OvPpXnC8hyF
B2lX8sUTyW2cF/b1jVYcyCvy8Gs5d4tQsr0Kkd/B6AKGiU0ypjhjC+GG3hzQ
PrHyhZ9R02h3K2ps9Tp13nXxyAMe1Zqotc0+ZpJ6vt5A977L5lkadN7Wr88y
ogZr0bjJZ+4eL3lUmok81DY/O0qmongGVuNEFbQjUFDBstaOs4HNtX3s66V7
mLMMDpA7G0bDXNmUgWVwBS4YXJJISJmYEIFiMZ8tdFyYZY5nW4bHJe3NUTId
Kn8EoOgCZxuW5P0A9JEyznkJo33HVqcD427ISa839RfemUyNzcALcQTDQj03
c69peOo7ujDPx3Ljv0nMjHq2wIe/IWLxpRaMUa1Km2sSvQi7e9lgMw+KSX8V
MzwEPGhng9k8RJx0gDY+JegkM+5HmNQJbFhgq9dCPRucHJGg5ZWbeegFMD5N
lPhMnXuecqeN5OHf9mIs8AiNs7/5xDHBUXnPhb12E3Feg3xQmbMD9H9ABVFJ
JZYIGjLDvXSDMZVRmSHrlD6nFDYpT2hYW/XAxDeBnAvJTWx2ixoGRKL2n6Bh
pMjULl+/qXw8iDbKuHmxxbYf6DOsR6OkgHErKxjmVQG3ielZnKqw67vbvdVl
Icg3qH/a8gBa9xdEdKgLMlfJhhp3bbVPrxotowjI9Rn83tNDcNCGmWf0hwok
zWwQPGMNaJIIkSu00FDrUZ+rVVogOhTWdg3IVAFm+omc6x7f/hx2uCj5sqJg
to78TIug/KbaRSAKKGTy8gYN9vGi3EQuOCGf8NJWmLN01i667JR3Ndi2fVbr
GKhHLwUQHCgv4l8Z5Fkfz/INI5HjQ4G/yW7vCefoq337J7QUSXYJruPHA946
KWwk/aHGl3jsJDigHpBTYufvNk5/Kt3oaGHpBR4HyQpc1nryyj6LIg0k7pp4
tkpFtmEefCq6JJaGPugi83tQQb0cK4hwcheRwd5ImgLvNJWyO35dOz9MDPrg
bGwN1HDtxshMhK2HOAAN+VJcaTXapHtB0bEUC6WHjZoPs9b+uG7Fj7iGpVcK
vXDYN+6sh6dkbKvB+/1YT1PKzr7KdBg3lYezQFOUWJsgp5DbTawwi4tNHHLw
EeJvsz24ISItlRQ/2JVKZ9NlupYJKPYS7GLhUUXSDngkJMQRjG729Q25/I0v
Fb6uOFyhZEudt4zeevZuUnF3d+azzJVxvVuvCW0c5bC/2DGkvh4dUKMqjXv2
xtGn2xtnSKlyzEMMjz/YjlDxryx8R/H0Kf09WQNneIUn9usFZPk9vIEv6inP
xLuudyZ2fXJuOmP/JjWn2Y2D0+Quy7PiWEUI4vnAhI2qHl5AWu615RbztaoL
3qVM9gMdgEFUla0QuHoP+P54HCfKdk/z1B2OvcACPKTHwPrYtQdOQcRq6g+1
hBikVzFRGYGJPpLMAl1EC/0mdODw4KaHYrc3xEQNcYUirE6yY+9Wemxw5v8l
BpdVN5Cvw3j768WkoaeEqnb5nao+5iM/rsyUThbMRfMLTtlXWnmrNnm+eNbs
AI4tucBihFMFW1PSju7NT3v8Ug5DOSwC4ZZsDUkt9J76t3cCoXyKb3YnrF5k
XH0tx2/xU/wJK7Jyhqh/CJHzppFTkR+5Du8ckVuQpGA74UsAh4fcCb+UkYeI
HiO15lDlucsibXmVJWq3OmfMbsqu3Qxw/dEcoMJwO4V6BpdUVeXVa/jq3Xc6
PN9hIz79tzJxWT4pFLkLO4SN7fe5C5IivzAQvCD5FEAa3ZHUPdXxKtGi/suR
KBOBoBGhzmsWoDO9BZ7sVoM89qxEptxhFB9wq0Gpm4KtdXul8xQsGe9++eir
ZUXt1JLEXFYYIq3niLhX5HAXvRAsJyZsgxP6UlgF2QiZsKDsL9H4VI3fMYf0
F4wylJdPa3lmM2xUfat+bjqBcR+qgX+Sr4KtEJBv7wbRxl8H58sW3vcxv5uq
VrfiTW5mntQq4zwPjNMIfNLcQAo7gG+iZCPM68AwqcxS/Qm78lo6FxQVABY5
tu3Xz3eUlZVpPtkCgMWlwEsLrrrqo7pw51Eaxp3iB8VxcT6gapvMfm54Xjfb
jcLfWzwCPB7LBIGw8EhcsE27YDjzzg3bPwO62+YmbERS8ue/WORfw5mo7Oa+
OQrW3vmiChjAgA3mCNblr7hv+GfvNkaqXjUZFTCD4WeRx9UgQPLA9pIBtpmp
36cU7TIViIfrV+uskYn0Nf1lRu6CQGcKnmQhnMNEBzo4tptgxww+yqeSNEzQ
lYc/QI2lzZVyk2JX6uqvK4aNt/bONlGJi/GbyR5RSV2p3PPyCO8ZqwNYh4Ny
a3Hkpp9PVyytgoqtZBhU0tlMNlt1229j6GVnRR53auvFcebU/lVsuzKIYg3p
7L/TeKT6eZHRNmZGfmpov1Tr6tKdEQyGWX/TyVnN+WwkyPpvjhE3Xl2ttM88
iTnETNTIyx4RWlC84Th4rATQzBzz6r0JtaLqWkrc05RIIzQ0hBDO4IErxSth
cJMNli6Rsw8ouCFfaOoPoP8Xvf7B+Z4TdK1YhP/jrjBkJHgKlCVywsfmKk89
qWniCDRWfE/ILEiF2UqCp0l4sNnc1ijdPnosb8O9nyxyhVrglN3cVF0zFAJb
adAV2Vg965npBwdcM7VZlrrIKyC9L2zjA2oR/ESYxl6kfW3kAOLn4gXWFBeV
5zYBnGAZo8u8VOP+2V2lGc0+ETeW1P+aMG0MUfyxyBYupwdDiHmVZfZTBVBc
11wfsd4NQgEfvpE5YlPIdDcAVmerWiiaZ+HZJsapsTOJkfd4Pt+Y+CjCIaSl
4AN7J1IeEGa658A6TeEfvziref8kDJZfD8rG9xNHcNe4f/x3kw+zLGkn7iiF
jprKYQ5kyFJ6XDrWDWocoDGHhwedCbOmum8NsZk37Eb/7HRIh5o+F4YnNsce
XOQiN1zUnSvTC9Z/nzazWIrbfIs/Pyg1Gm07fAZTAPXyiFkJ+Usjb9XNGx6t
9g5/0RBzXGW0S7GILeejMdpW28zhj2guztvM11sdVBvyx00MThA3laaZd6b3
R/AWBA5cE2zQSgQAtzpqQYDdwURO1V6lMT3tjzaMm90atNhUrdm7KojyJ6cA
QzMrdjlDxEas8fW3TvNjy4lMnUHF0CxZI/8A8Gce0IG18MHbqEv8MaB0IHDX
j2+tLtggJypwZ7fnDnMSuhWJh5SFdM/SAPmxcp5/caDM0/UAmZAXy6GzHADy
lKxBR50cL51vXZ4wdYyP9jnz+GjQiE0bj3Zvu/JXrzWwFbgBIkswSdLFJLq+
ppiHeRycePRCulnrAnIZo8zmeEath1nnXARQwoqJZnyq++LD4PJ58rj5hDWO
mQnJcNUSKFsDxK6OnOv4R09NvZsUhFcjjwU2znNoVX46coArBwZj2daAR0vo
gE8ztz8eZ8Z4Imdw8LiQweypW3ovaRNBG/7i8QuGRdjTISf4sFLNK04Koigd
ptv8UoOHnFTZ6sXt+aUgloasghmDy/qiPdlLAggH0ggqS5v0gkxMxjvznMAm
br9VrCm0JZiCruxaglUI8TqcALUr8zXaWXRStAOgvI4xL80yoEGiPOXqevHv
Hg8sszpTOGkcUeDjOZLiFSqWjpOguYL48txHz8WyDIt9jDdruVzdBgnyAFzR
JJtsaDfxcUB1Q0Jhm0Z10z+TN5IH1InFL1qt33WngL7VTfwAVlWQ+EE4oKkm
cD2ECUzAtbqPwFolhFNo39xm3X3VM75zUhajKjIxWMs3satrZjbXUK8BjqcF
2bfg

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzf50UjfySUDSJmQloo6NQ9/USpGnRcFAt94AzAA7ubxx+gYOFsjR8YJQmUXFIR/sK+RfM8LWx9VCrimidvmO0gLliQmDhbcbzIfaiN1kqFNK9aFv4dVqsQyhTtYnIPSDoTr/aTe5h9HKYgr8Pli7X9c3Ux38EsUrYrvW1TYOraN25MYUUrNypZjihUMfYpKlJfe458eiCMh3tFbGcsG/U7qcWfRNpPatCnwuD1bHryqMMHMG5B79TGV+aKSMbO0kLUdAcI1vmKoTUiZuM4igFNV7cIg7YAhy2bejEV9tDS3RUvWthi7sQk6FvEfNNZ2uDWzgUvpxPpvZsenkXiN188l4Jl7yXMHwHSJGM0RYlRw4jD1n2N3us5yZ37k7sEUMBn8DmYv7SXOrK451oRD9RFHCbQmhV/Psauqy9nxHW159YZAxpL7KK8gr+r1Nr+Cyg047Gcc65qzooQM96kPOK+ihqFionYTcFK4U5EFvO3cSckP6w2+l07clmEmJGBqqRE/AwEPFjK67l1X58tigvdrNh21qfAYb1MiFZL+UwPd9cUPtSRDhaUY+aZMgDQ1eG/fNDfGfyzDc+vC4gCTBtINl/1qYR/OLpNBEkbys04+iIcuQGdONVzgny8R+X9EGHjSH9UgdmQ1t8ocqgl3CtddnbSLRi1tbqa08HQ0vSWY8rgIUIA3oVqp1CPi2IzKw1VP75HNN3xQ/mt/VFvMsTSuvuing73c4OH3yniDMsawbDP6BXIXsfJYcSYr129d5nmOiaiCt9yL7e4IWjFALvm4"
`endif