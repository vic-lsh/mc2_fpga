// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fkLklBhsOjRGqL0EDuohDljmb2BXKVFVwUFA0LiVn22KJhPzwfhsQiyvfQuh
tYuzDkyEFUo5OGbmikt7m5qTJnG7+ZMOJZHH559/0dmhnpxOjlykNfq2vI1R
FpqKkjD3PsTIhM8Oy3ktntkao/fX3qz3pVoinAoTKfg5kp6xbOy2EK6FPED+
KM+KPdF+bheyvNS4ZMnc/gjf1XJvqKvMGA/PsiAkUIdAS3AGcBhxbUa1JTN3
kGe+YTjCt3m+PEN70cAzScAIjdezt8e53BZn0xwZWS2YR5IIM8HQzBV8YFNv
kG+kd25XeE2i9qj0OzxzTxx2z/KrKWpfoRMCn8KdMw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gsR2epVbZTsMlE+Jmkqw7mesmGA86+nbyQQ5rZ9uU5kdDCjQuRiw8u7SzQfE
3rAyquf3Q6COLuitnEIVxfXyTjWTUcPzjZ3GeCgiE5InaeOYOgmyLpUuRN4X
rpRgt5QLxGFSY/tt8izAZ9kWeCZqhzpU6+PH6iWEiSosTz0bOFS5jYdp0POl
FTcL7iZ6T6WL8ZjR+u6nbwQB/D/5YVCocKN+TDxE0rk7kMXNK380WVk1FrVS
/ytqNcNZ6vCh+fQCeCisUi9yMYKAN6WxVGRdEvClI7DpfRpHZhiyqSqcrJIv
hDfqod9zr6YF1kg1eXw+GCB0i5pzhrOpvqtlEK0mlA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
M8AyaClfDG5JVtckokZDpaoDCML7b5zij6rqypnhUH95I90gcH0BWG76QzBG
vPrdhEj0QAMsFEMkiGVKN+yEECxldNZ7bxHAQ4xAPAnprBHlQmAyF6yxk/6v
vHDZDACtJEVn5kUX4WOD5518Zxj0EYVJeGnbdhHNfQkzxi6Cm+0oxnSCgcp9
ve3HvszuHuwMMSq52gpgyBVWEuhb/5u3DmdvaIBODZRRswt8VF/xdYHQUt15
I7Np41rmim/6F8SXfQzr7u/P45E7lmnFD/VwWWJRlLi+zA4qEnb1oV6vwzsr
xeewd/5S8Nv2JeWLh9rZ3LQulf+e+tj17GIYjuRgzg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kAaMC8xe1QMNT9Uu0i+CcZO2MVhzDl0NTLo69agP5eig9Ib75iU+uar4jHmS
cTQNHvbmMOIKPiU+JweXwij/MpHfBfIBwga0saQLBamzUnlbWYvEJc562Xi2
Awd/J87L3DwtSleoTNUe2pQteejwoq41XP7fa0MAQphsVBKqDtBs+KszdWX6
ZTIXii255I4Ejkre6+h6GBuvNcixsI0NUe7DDOE3RKtZrfKUYQpSRFecIsLG
3hGdzTGKdpeZXZk2liqxsJPMq2mBztyNTRORXYw6+VqIIWaSTW6cr93NUo/7
RNIFdR8ZF5Y3Xe3C0Ri3/TQZ1zO9u7lnb+Xg3UyeGQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YFzcw6J9hj2u+2xwgrPaurGVJMpOvF5ZthlVR5QaiGjHoUqhaMwwi0ng6V3T
w627yHcHnCfGYBiQtJ5zhrGLC5Ur5R47ttdx2rdn8SPhKTuStuj9vQMgW3TI
JgtwH/j4L4zh146JKWUgtHatVQ0UuDtWWYuXGkogiqzogTixTT4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bI9qB0USUvBIJK12LpUMl7843jqo7HCyKy90RwFGny8CKGSj4YNFHBjVBErF
ez5wqiWwdmSX1LtbfoEj2000Vw1M03KCOksHi4M+tht17ka3+vK3htggjtrz
pUdzkQavqr5UeaVMTcpNW1TxkxfIhFqBoM6Oo/a1/DpSFgSWYwRW9gm4J8qy
lj1gaWWt8vq0c6A9iVYw5zuOm3xejNlIKV7AyxuaXUV2yISizL3bZH6BOZyU
Ca6MFsYgjEbYuT2es57/OUJFhsX1ygM55Y1q3+YVLZsrm5wibLxi0U3V2aLr
U23g+rQS1guYc+Vxl4m4rOdB5VfBrKNJ4XpufAEMHfObk4r/jbp9kAL5eiaU
ew917vJQvPFfHVyyZnS2feGkh/nCn5zbhfmUaDBWM+EErMw8iQapGNsWChgB
3rSxzuTq4PhCVffIDMLYdNMCLcYgJ6B66h1OuC2A5i/WrOifxFy7gtEpRi/B
GeRDGF3RNjSjaZSsNvU2Acdd7red9LKh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K+DubFol1uCYjZZgtSCGJ0s5OVaU0sk8PoYwOCoQZna8JgmnyxAQVmaQHhWJ
HfiKtJO9sHWczaDGwr+dpfGuhcPR/UB5YV0uJ9TueUWO58bbdGtYP4WH0c0j
zRhhXOLg6DyNgl/3k6uG+LVKdHn0BRJjbve7j6F+A4D8pSEELVM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eD2bWNMHkqeLXsoqHbk2t4VrmlSitQT1o/YEEeooKpP8CGSO49CjYw+u1Ksf
iamzNjrmCIYq9VvdUYj2saxWvyThyB8nnb2SjzH6irlEJ2OSVW6ekxGjVeQR
i0zqkTjm15QwmKmbrj1jJ3N/t2t2jYO0Q2+NPCMKc7Wb64vCkxo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 35184)
`pragma protect data_block
yJ8nIxfk5LR9GZ2K3PB31Bj9acmF5GwqvXsNh232sPoB94krGTiXr8z8VwR2
LjEpC6Vht+yEXwBdnQWPB1Had7wAtPYpwmei7HTHjTn+gCw+a7M6FQ394SGJ
e8jHu69sh34WtztRV4/E8oNnE4Nw648E8maRqsuSMHBynJQLI/Suy/AZmgm8
VfqzyacViPgZQXvKOsr/8W9WjHr9MshESrRNByYFEXXUTspkVoRRNsZxPGns
6znQWFz7yW7Zz/rdWKAMdNRMpkNXfLjPF43o8wbAMC9P2Xgm/V3u8kjF5Emg
42uF+9472RSKDhbOQ87B6foxghjd4fZCLDKSrNamlAGbmadmc0GcCzyGnWMr
7vXg6MYWdSii/bygpmvjmDdbhySK02Vg1H+h5Z5HFN132IkraDRtQQ2PrMtE
37MuM0dG622MrI9UExPFtcJUeINEcj13YA3o8eSl5zT9VO6YxSP2lDgectrV
1sTg6YoCgvgkv8y3DyAnxN4iw7DbV70v2oFF6wb7t3/3+CIgPtY8cVPiMHlN
0isF1WbMvbSQVzd6YonXUYHNRfVcXP0SugqzADKtsMPbngwx63zADOTcHmB9
ZmafVM4hoZn0dVys3Lc9z0ZCiWqYyaUSMO7UDs90XMu+Imxxj2HFNSbl3SD0
tI3eSTZRAA1QXCyWCfaIiclTrDyBCc00OxFXHAgwkF9u+pMv85PKCX96pwkv
H09LS1WNusaDH52HVPRnCV5RJyOAsKcn08BUjLDiOeMhEGtZYIOxlT1mxHbW
5qt6nejKoGrDT5BZfi12f66dI1gEnuNSQU4+v4/4B5iR/SmV1cCzhGHFAqF2
2mXUIveobnwFkyNWpwxmKxyYQW/Z3qCl6ps7V/nlTXd+xcFTu0F7woYMEIFH
+Ks4TAcWM+tgPbnt6OYjCZqWbHn1Kv8kMM8bunlLiy++ePqHDkB7Kq8pnzDE
CQeadaXKEaJNxcfRwOesx+BFQD+8QvuSX95vBeCiaPn3dP9fGg+QGS+pK5Zw
RmPjE+99PR8rinVwJJBKHRbtMduHTB2YZ8D/zIflf+nZHVStMNS04toc8RJw
1N0RudDZP0eePr/p4QwjIaO4b2Fgztb58XO+kg0SwLpK0bQFQEpgBl9hsT7g
2kT+QGaCIVQJSjv6A9gS1twEDtnAhDDJ9jLA7M6vO7vK8H5XMFPXVZbFDXDv
EACuOnwkxl7+/fcO79rPmk+fJRZLcJvT2fnR+r0pnIUrg9Hj0vAHIVb8zv96
9SKTIDaw/24J1z7s0bWXkTC72gAU2yBKslsUiQ9bUHykiA6wXXwjLjKxyedK
aS+hnSKVQdeSAkkCGzWSRoQxbBz00HzdfNgomgrrfHiC4hptssAlKRije447
UCP/04mRwZiZjQPz96TI2p4sl08pifXzf1Mv60UgSF0TU0P68JWxkgugMWht
g3tL74cEyIsX/Xybi5nyLj2Tj9FfZQm3WjL7FvHRoA2ETkHAAHZWICRg/Mho
O6TdX5Zyy2Am8/6k2ih3UgQLjjxVkGIBIQLuxjEycfX2IF8FuMDXYw6W/azo
7RNar+3V9PLXZjTCxd8JWAx2e/cjK/QW70nl9frxiWqgzNBax4oIHrzxAN0M
A83FJKwxcyp4+3wBJWHWJu4XJ7/vShrVyHmQmgNCH6VBjilJGS8nhF+TW1ux
34qvBVXzruPXsPVvLgV3No6SqyeqHKMcRw6SX1Blga7T7Jt1t7cpSA4N/JLh
pDcdhNaRXjh0wENbGIrN4dlQY2d6tkIrOS2ksdUOBRa9SAfhkbuV6eRbuvh9
5H3EJTJ6Y0uKmd+Gtyc5M2a581hH/Ahom3tCfvRaGilPohdJjw3H6TFIoFST
CRSW/ABdRvdtKDJ0VzBpn/xH19nc1TKQa6oFYnEH1thpsIvuxbtEjw7yrzzN
4n8JnuT1uSwM4sbmLZ5cGWnTQGjThmsGRmskkSy4SqbM+8N14dHUTpnau85c
T0WufkXan+Naw4vD1R4uU4Zoonb2awXxAm6qZ5J+WRSYt0kWUeAMOkOclcBN
sJFzqyVH24j1d+F12XVtKGgEX11arwtt/xjgGrMQlkHkeguhQrYv5x1yAGNX
Z83rLNcUvdBmwdxuAZBMz4DDyStvbNA1odZBoqiDf8J2Xyc2bBOKfn7pW3Ff
VBM6dHS3mPrJpDAkEAjd1uEVPv7Tc2/0syIW0Q7DhvYDkD0OwRRowMcDrSVH
Lo23pgCoMmVM5DMmOjy5GFfDJWvZYM9EinNDJJ8XJtAtbakoyN0TdBfLluP0
OxAzXwCTtWY0C3kx0ZQTlTx6Ljak+KtBH9bKwwjF1zjBNx2oND53CxM7N4jD
T6yNM0XB23T/jnq1u3e4x+CGTAG25T6RhGUlwh3O5iL7bwFYQX1JBvOfZdAz
Wr1JNB0S1r0kvif2dU0cmHasbdh+3hceRRjAfDZPfeargUAooQ5JWzcfGrMq
MSX59x3GgujryZp5Pf4vCQeip/sSixxz9bWljwpg/Oh1GtdsfGMlRF4vMfdC
b3Ra98kJDJesFq86EfXEcDPp+hNvlkmWAyIIxmkhKCrGB5sgIjl7VI58Qkoa
jI+gcnkPzHKATVbBNf1dkKEz3MZSYL0NuYZIa4SLC2H7hM2/usFTT7EeljDW
wsiJjwJeiHvEshicPaLlruykFbe+7LCqBW5dd0TMFIbOy/hj4Re/OY2OddGW
doGVll6FYn/Dnow7p4Z8HU+j0c8lpazsbPL5GthrS2oeMstUk/Ab8MhqGqyU
WAnFQWZZeztgRkW8vN/ZHXj4kgNjrWmWV8sIGRjA6I5f6JMIAS9N+gEH5iKd
g3g1w9Yf9LCR0edlN/VApPyItU1y0gVyi3jFuh7TSCPEImCj23DvsivEytTh
JsQdHRN1a8Ktt9vqrJKI69Hf5lXikWM4X6UYTzodvJYQuAowP9Zofq6vhW5h
HThkB22IyFd2upOBOhgLgpVh77aaDWZW4Rt90hoE6aoZRIIGANoNZBu2SBM6
kFHkZ00SakN+MprdZm5zoR+byF99i73YGfSpOgN8sNyUJw6gp2Ayu+dlhin2
fZxw/+LnRLz8yu/4CQFmB+qGBKbzr27/vNlvkalOB4XXFWo0Jz0u+/jhAUs6
W9QDpkF5ww27cFs5s5GCLobqGzkubfClVYOSedBLgeogtmERLqKpk/gY5oYk
VY477vFkG83jRmFCRTErOrrlt9+yamd2CDa0iDSdcoYq4SwcZhZq1T/ZOs3A
BVgVH7dwH/vqZ0NEkATXYSifk0vPbC2wF6JD+0ZgVlmhU5Xr1TScWH6qQLS5
pE401c5flKuGkrPpA/tevJU9RULKPN5B2q2HSWz9zP7adwOydKkicYCgqtDW
zzVko1y2U2JxhR/2YF9PpRZ0XJzgDazi3CojIjzPzwfK58C+2DHZ0AOxrUpx
Du/QBN2Z3VRIA+J+z+ZTfdMs6IIFQOVSqWEjA6eQvmZlXfOe9scU5PSdw2Ri
DLbDEo8HvL8/6Uk8w2FCj6U+GicTapq0voXfDoHbH9Zklmpk7SAUVcI9n9nM
Ry5OwfeO70uDiCPxgM0TFMzT+jZ1RHgbgphNWqu6QvpTfWUYHlERuxqiExtG
IFCHI/IgxRFh/zdy1r6WPu9Zwoo5pgXfM4/RnHUd2MB32DcaCbsxiOK3VWGC
IAxEfj7Es7CTSpreuBsq5PBTY8nJeQIhn9rB6qIlcwMQcyw8qNv6+Sk47IXH
6XKIflbveZtsPfmy2larZMviK//5WHAF1m2yPLtZsqnOHTSIv+CZDFQauXxs
cT9mYWj7Fb7hMtwzlQu6SozdAMJhDmniK7618Q2aQZ26oT/XBWyj3V6gi1+p
mOoc3kp219CmCAfUkK944nim2HekuzhcaomZi5e/r5Ro4DVXrpPnlnPJ7Zl9
lJ/e3tl5B7nVv+ekjrKRpKqnXBvg6f+3kIEw7W3/GnKhRfbMWI96ievTGrfb
tsE+9AL0km39FZVQqftzIN/CUwQYA90sVROHa0T5inpkwqnU3xNEwKm2sNjh
xDW7UM9YHQmH3R8Jjn9r3+FtZttmB+Ta78qyTjm+ZS9PfhPeqKuNZKvuAt6J
xJ0jcYotSh9mUj3zKaF699KXF//TbMz9XeQI2K7eGwPXWy4ehZp2MZoBn1ce
YBadXtZIsL1ZRcM3ueUZP2NCs+PsleGta30kmf4CLn9PxkPnnBJhnDWvyMlm
rlMvRK7wLWaWyKLNwL5OI2bfRZsW71QrlB0dpBOhpBUTDRKR/zVi6YoK9enJ
QQQx75NUIFkSbza+2erzMwxXeZ+ilv5uj5sGxo4QnWDUJbDgFHd7lK+Y2O07
1MuTB+OuP0oogaZtulpWh2rhqSLEF4Ey9Yc6aKcmxH6aHSRXxblWqBMaVSt6
wh4+xW6RiWEXYWTSR5R0lZVVYU+iQQLGDZUruH5bPpNpEaiU5KyZp3d2OD8f
x3wZZsbKovExJLe/ZDXvoOBkZWR51Eq4R79BCzANSEKIe573V+C/LoMNjdTj
BJG1JzSe0jh1t9wOzhOj5tHQvI5OeoZTOnVS5GOWXq3kB0lAHKabOqW/IaP4
YPVABi5JXlvaiOAoWqS7IvixyNmB3S8xQz2omZsMVTW2ceq0xKDFIDL6FoCE
N+i5ovKjdHlbr/f4/UfRBy9v5VnhK2An0n+YuIK5UpzeeKpConrjhd3NZG2W
vTZSj/d3j61OqrAr6RLWZK+g4Hs+abvGKHpQawJi2pSQb6f3ahQHOJ3YHG3Q
u2KBWzLvJPRM8YyhAnwwvgL2mWI3nef07rXw/TT/EByeJtYQMJMiKlu9uC8C
36j5Hl0Js29IjctfEMfgR0VVr1UZ/ZIXzolhSKs35AvEI7dXHMF8TeYReqAN
wI29+o/DGy6/oWwr5aUxPs+yw2WBrCNL93EB9WZtRyzXUc37RZxp/Q5jG0A7
H4+4O+6B7NVJ8Izdm43k0vS/GmRGyON69hv4TkycHYiWz+8ADgOVMo/ge55i
XlQAiECwo1YY2I17ykLC0W6RO4zI7dzFwYIXFlO9ySfUBUWdxRhFl9YNp4G5
t0yhVhLS7uvWbvq3TV1FymiJhpcnOuF8W6gTLNzwrqfHDrE43mu7w7AFQorG
B4GH0qklOS66p3ZsSbMhxr/spUa9xTM3pdxhEX4aNwY2epPkHUoDP/aJHbxn
wr/dYEjFqAzQUqtvXXXFU12LukaWORRiL5L4zETmAdIFU2m8xkRfBGK0loW/
aSJaRS0h98BogMzH9vn5+aCs1sdkxutWLgWtz7Nfg43PhvVshq7xHKx6tmFl
yZeAyL5+cbu/nqRsSUEa4xIYi+gU1/DemUoUWjxN43yO4fm0kIk0TvUqRO+E
Q9q/qpuvFOitWq0iiWuocebj3xPUfD23TjBROmwejOLb+SV8WX8TS3rsVc6R
Tovs4tD24WR+lrWVHMGYk5+ye3ZZYyHx8chTVlvhVXZ4pNlXqayZgwBsOkcj
ddJ4QyWJycOOY4JQVYDOLuO+qTCeBE3KEgB0N+OHGb8KyY2ZK0XAYocsPvJd
3ANMQoOkH67y8txzxikIcFLwiYzWHfEvY9oRa8Mj6a3g4mUfWjYjXEO3Y+y8
tl4UvcOr7hDoKQNyiEi9zLSCOnzpoEkDPH6HTMzjtZ6AIBxvTnAvlJPtwNnK
ZW6+z5ITi/1Nfkz0AZWFPxHq6fFRcAxIthDKokAC/98iqhq/IUOLq6SmIn47
lxkYir6fzf1nkuwToN4I6B34aLQEmmR0lmJR/TQoKNK/PGli4WSCV4ZGkQaW
f8ctbAkxERBnu86fLK1EjCCsKQ7psiKT4QcOcec6UAYzKHZj3c7CmFcDeFUZ
wh8BpwacL3nWM8vF8PoKkidl6uwlsAoqOZmr9quahBRiZhEyvPmfO6BP+Kkh
IzP6lTHdgV3qumdwBF7qFNjzSpksqImEPJoy49yAmVLN0tPQAKT9qaNSYxvu
Osd6q+YslKGJAKs2qT0hJPV+w+JxV15oslLXvIE8QBmzeqcWLccRxTEWLe7u
uxdCMjaSqb9ooCoD5DCa4q0A/SwihZrduOQPdywVkQ8xF5q5u8LcuhJEuVvP
YYMnip/aS3VVPWa3a2+yxFJGJf48HTCHNiv1FpXrQhU0is88e9B8EeSBuprR
Bw2cn3TGXp4kUUSJsDimXzWkNZVwQPv44IM/9Syw+TEXVXV28Qip5C1Y+o0q
7Yu1D6kzvhhhmkdzyTfyADSgQnLP91Ef9J7pyGM3yAkNnVz9qsrPWyt8fFSY
lmSv+gVcvlLLFs7qlDIMgALxN/2s+7ZLcSOqTq6+HDtSPj95TC+wNNypfoLK
j3eag1WKN58Cpifl7Q7drgrAV4ykH1zqMkpdhLmMTTb7RA9q9M1V6mUPdgPQ
HbdLNdW/R7g9LP2ttYiKrh8PUZ+lH9qK8BflH1eKJrkp/5FUxvIoZ28tvq4u
MY9JSvoH9zulXJHLebXm3O9OEHlDsqBaa12t1G0MmNXLfvHbvwM44KdjOWpA
ZB2pgQVapgbKEFmwkrh2KLd6zd8ra3fZYu49xVsnTAKjayVIpMQjjTl6SXEr
XuW43lGJgdH5RThf35kPISEhHo+0Ts172l5BbucwjSH/G1EzJbXTMX2kduRJ
bdsn0QIYQXW9BbKZuuthtysLmpdUaSBJ6o8J+czxCxMYhm4Ba6i3lhjus6V7
LNiIgd3v2nui5hazu6MxgqArO7WcLqoXOabHOjaf+HZyN/tqoikSJ4MOwuXn
7ncsv96ZUtQodw8hWez2b4NtgENbUQowq7/Civ3nPHRUCk1wCN78yjE5iBs8
S08o/7FgOE2gh7R+Hr7OMJPtS7jFQAzTQFj2azsRyPKqQeBS7kZtwVcXobjZ
s1JxOyNZ8oPEObTn89JDxpYZXnkvqQuJv6cgS+ok1UkskaT6agXzjI+KjVKe
TIzRuRkpMfN8rYPGDV2ZEGiZ9/KYtlVuSmXUDdKczjIvWDDr+33b1b+i0LVv
Z/YVdT0MYKrYe6qdeg2hWziF16NnITNOmTeCFTjKEFVeikqfKBSGB7y1A9Yp
JZxBtNathSMUg322KoOCDpDpe5h9JUegTsoRHsm1Jqi3/EresQ3tPtgmnVE2
A+oivQwGP3ls8UJZu0EM8U1mf5FqeCM98z4gQ8M4Ew/Feh3/oaVYSqXXFNwW
5G+qh2EKL7bMLUm5D1xGJgQP9VnwtjPDQJLAkKTyxjPMuUQTzFjc54USI1QL
rrD2xgcersq39yAJLMssBWZUQvBMVMauMP/Eu91bWo8r7Iv2i7CMeREZC7zC
+RgKfL9UljmExFYeA53T1U0IR1XkBz171RELB9j0p0g5llZ4+J01JGYlNSnw
iDMbIxPEIuE+10oZVURCBel3+owL898qzjjMzjqq51m6kpbzEEVrRzkPRIhY
TxpZAf4yU4QOVrD1BXPDazucM/N3tHyNtzOpJmlK5sKUBjvszbzn6qnxXeIH
E3K7DrTQuQpQbUZbRSwS7YUMUYN7lwQ290T55jGHES+aefNyLDd9svtm5DAM
D38n1xQBiy4xY/BHC24Ruoyiau9o8Vn4jz/Sw9EbHOLa6H1/1P0Vt7dwNsnF
DqSVdTcn62LhXDgSn6s2vwbI4nfv9O5mz8WLYS5MTfPuFhiDwKWLO22OXdwR
TE87aOi9m0sR2qJOVWrP8vLjlGmadSKYOzTlP4Qu3YwPlo4ThRhvrh0CFq2I
YESy638kQTVW5ghOBvDhyQDJprmKa/Tn6LMadOLpqbEpOqUQJs0oBQznQSPO
fBWcGC0lzcoUfe9nHRRLFF/zEe8KnqzW+dWsndEEGOa5suHYyotFHXZ6eVH1
0OfyRqPQUXaeAKUMcwDvMbLD0ieWWCx18Qz/k6rYcyK7xPimMyGT97nj773A
8IshHaNUoYiRTlkg0kWoFuzonN/RggBfKlvZQv8ajcKLHQFBl2iqtJEVNFYR
XsoaENbkgZVo3dDsvnkhdRQx9M3nwp001Se2pC+1lpNu2CTVe5jRQWnf7shH
PukAsvUcqUxcMfMI6ngNq58G4Vr/v2Syw2nrjWPJSzZd30ydYzlWXckPcerp
l84CcWvITY41tjHiHGi01BJuWTi41+LxWSDSqgqFc9UhzFiFMMdH2yFLSxVh
zoNOVEXNyTxN/MLnBug2RqK2taFhNHq4FFSHGEuHTDIcP+/8GgovBmI/Luse
m+r7CtqcWFzw9KGDJ3u5Xpo6UOQfq/+7gob99nL2+RLZg4y1DOPbtgn/xXHd
Soyc1CRrV1r0X8WU1EfeqUlD9UjIlce7NkcytwpA5AzymLqKo0gmkeQvcTVO
NH/vn1Dh8aBdUnqWStfVWHaglK6AVQmzPVn33pKy3TGpUd2K54+wWe4PNX1m
L4x83pQn6uKlynHRdj8sfoBIrARt63AjQWU9Ezqy/Kor0gLkV4bhgTfxQC/F
ON8DNk44Tq2dW82ODO594nGyVHBQLFrJypBFeoNTW0FpoXsRzmAufDtdqhwo
cXVUCwrvEWvPn9Q1JzPQM8BJ/9tBkVPzKST8YxGz1kid9Jx0EszaGkaYvYPJ
f9umr5jsBfrq1HiNi8AVyOzjp8TIFz6zWrppR0+SoA7JX8NWkz4mVzZmlOli
PtqPQj4tsQqNEqwAXnMfNAQDD50uFmhCADl3JPJR33UF1Jz/C7aBRKswkHd9
ffJ2YtkRQ7eOGgMakhZWt7a1s3t4t162APmLoPa2CiZtkFsJW52WMe4CwW/r
0eL9dCxzINaASSVzvdycyhwDMNN3+Hp+WuVBLaoUJ0j8dloiZxjpfE6wfdbq
PuC1ZTM2eIuU9u/ewqFeIbJfYA3g/0u0I8NyJT6gNVG7fmrFuR6zLqpz51e0
djTxomga9KSWDRnTG2HY7jkrxv3SlBZc3xRwgBnelSTQYJToOsR/ZdbrYiqO
/yHH5h5IsNJ3t25Km5DKqUFgktKVbd2Twz2w6+aqc7Eum4OF5hiVfcJDWtYA
HQML3jKv1bpZf2SHFk5yTWjas4lnpF4+pcs63nZTushLmyydeenAsIqilhce
ARO/hcyHZN8aow/47TE3zUQDiPGSPxTWVv3AEIhFagwNP7bRuqbDrzmvQocE
sNF5OG3lmHaRul3o/+9fWiAh9dnEU5VMFZ1Prr6oWLmO0/kdIRcbkjt/25t/
+KVRIBNOMdbFv5xb0lHnRoZY73Um4zAQ1O53xXLE4QWk99dZ2avbf31lPX1h
BkOFwX41zLsR76Gt5+oJzGu4Cf+O1Pv2HYquaipUqOtzxef7MUTJzqQCnyTT
7TWgV1nZIOhdfeGehlnSfkCjVlFs3biMMNbfuWlitMuoFC0iHHrpzne9+Rv8
rN/UdXjCI4VVcDk75dVJCOarYuVSHHuOCJUxQVxE2V0YqNNbxxjq8UcpNKnv
N3OwYTJW/7Wb/AtwnnIASgDBN5Gx8jM2lXpv2CrWZv4p18lq7I7rCYXq7pG0
vTSq0bz+H8LYEozP8hd5+k6LUu3eUC2ZT6K944PPM7rYc6qsm5kSvh1XKuP6
IlNYenMaknrni8am3EodCzLOnnMAjUp3iGvT2zwU100UsWs2RaMV/Xva2YCy
0QKdTLP/qgQLmSGFjSbjLrNi+KYsCKwFsJrhbsdo+65MvYaHydqCcDIPTsz8
YYq2bnv9UOqQPS2GeG1nNsYCpteMUTD/U4AcZeIMqTxQsFBjvTStPxWOs719
XKJm+UDLqJoSxr79LJCDr0GA7ZZLs60Gx8u2BfbZLy8nvT5MVO4KmdCtM5uk
R0vaRHsg3gJFXnXfOA5HAvFYOwg1tsY1McgcJAvRA4VrbZFLb0e30qbvhhwD
5g/+2/HuDBjWavEJA+hDFSWUqlE4HBGgPpCf9VtkdyblwH0WV3R3MO9Mrw2d
vhuKUI8fABjFJ5Mr2Di4W4zwtzl0D1vWfz+hQpl1nxW+Iv8Zit9KnK195QCG
xWViQ0fe1IVwwnUHrjM0EDCyTzooJ3EqwAiuwoktMsOK4ACx4zFN+OXs+7dh
NmfBBPMRFncAGrTYdIwLtQ3AU/z3qV8T8evQjAHdTtogDT+pEYfy+/6eBBLl
moGnDSQMYqDKvDzquCKIztXNB9ORyXDXw7Xq3NFQLD93ojFPNbRgGAgboMf3
Hdy3ynXGii50v4p5FVy/pEengA7t2a06iTNItjxfeVMhmErbpEHWLbCvXea6
iYfHMczsBMr5B37KfPFKvY3JNdBhXsjrkF9BcGk+duQRnS4Uw4g7nyFHpvBv
r5zjLE3uEbGPrAl6Wdiltftvei+OeSsnvT+qtgV1C0SPXHwqS4nDsmBvZdEe
qJ1u9jnJKdxSFjXiZl97cGxg9nJOQJRNhjS+aY3FD26D0VhA4B0Xt18OR/db
wjh+R2jOeMbc/RUXlw63Zi3LKHCAYa8f41hoMDuJ1AacmGE5NJ9sBCH3yzdQ
VZ7aGBsa/5RKfc3l3eN9yQ2+z1XcqEa7jeBURgGjAbXESir5WkTAlHFrWvdW
+YUjgr+/8/jJDnarXTKSCJa/IMPXNqBdpEc5/Xj3l7bcJV4+qyttLctcEyw4
qr95OCkAYFGXtfbk8G0aCmgXB8539GDk04PrKnrcnBJq8v9uo5FunVMp7w2h
6d7kq6sqmz2+ej7O7Ra/Y1FVfumVFNV2/JCRBWTNHVikT2/1fjotcXS36cuk
d0+HDO9osmCD6FI5tlOnKqw6KlSYNVmpZD4b0JaEiA8xhfbzyTvyaeMy26ai
LHjnUjZvHBXjJbHCdWWnt7j+LjBKGiqgPg+BaEF8bu9FX0G1AzLWdVMnnwYe
RUhlfFrMqdRE9LxgxOVVZayZPbgPMFAB1/SQmRx+m3/xfBC0GpvIixs5ZI6D
c1yDsQbsn1PgfOX2gi+DN8fYbY7OErya1/deokgo5GSE1Zc3QQNYm9pzOR0y
9Muyg5WizXViicaLdrmj2f0uqEf7zhpkGZLy5JX9DBIr8f0qvpILeBIQH7vy
IxcPygd8bHPZXECp/hXS+pj+63SfNLE4pp2/158SrsJXG0wYWptM0MbsLKBh
NUbq82UtxTxTmdQHw5Zj2djx4OaBRSszfpa1fJGpTafTWRNRNaoH4QB/pLUr
siqva/zP56mPTQaKSJL5Piv8M8tiKhPM+XEFXT2DLJdixuOCNJl0RZ+lbaZH
8fe7bu27xt3QTsDpayCwzK9GIdoK0RK8L9ho/KH8pypxinJQdgyOaVsuKXJx
uABQBYnVeuzBcE9g0nWjyc6DVDIS3InLChE76fz1DtU87xwBKZIOX6yovGme
6+Cv5KD5QBQzurR2nFsYtb6cKDZODDqH0hKEQuKmMrlE4Cf8VxxDRsXYNf3x
RnKMpAypR3UpXkGf6ARcEwjzGqIBk8ItFywZ7/lScwRZkIerLkbNLkkH0T5n
y/0beUjmgSgI0eJY93j5NEQlP0x9z8Wmk8FZL71JfiyL+S7Y1ZWakc97LW5q
kM+AvzlvTFIkWviQrdUYfLF8RebdpxcMYrz8LTrCVOEyu9mkAY8i8hIOV2tL
qdm4KrE6zCnS21Z7IN9sQ4XngQPiYAMClif6lGHLkPpwtUOhmFQpS8l37FIM
PcZqIqopBeFuV9s0jHQsD2GG9LeR++9WwvuiWwp9mwsfavFeMj2X4kE4uExY
ZR0LtgwVw5USqRuc1lwCS+gjCrZsJrH73l5ViPKODCGUhfXChrsmkjlIzv1F
xcmWyEBi1Ax6DOpgYJPWG2xdOCY+qHnARShpBJ3YfVOlEHztcuyaRnpvLjft
h8iXYZrqmHNc9GegbfdqpbNnFLpQO7+RoITgm+XAPUGHjP2YeCLprkN3oW70
M7F0cKLQ+5pqL/+Dfp9KU3xEharnVm7PEXGPHwYhrjvA2k3Ep9BDiU1uGsnx
LHwbCWfS9tTzSe4SxxBGkxOLzX4ZWS1SEMK4mIx4+mWkyKepdKigBYvBh5kQ
udM651HOCS4beRnT9T3UbyIHDVokNM0W6cOJK4+COg7qmfmVPvn2WoC913xr
OVmLxkImN7GFxJ1PZR1kl7lCNIuto/CVyHZzhclqirc/WtLFrtJUhUZBVd55
pF/B9wYSmLJnA7OijgGi1ST+kT/cz3/MGLyaJ73UteGMO4FlCwh2fYWXoI3K
Kg7BwTBixywOemfTemKdGSDDg766or96tF0tJvK8k9KWsAw2oD5HiChHpUi0
+py+r0uqHMfQoCjAWGUczb3e7G+y5OBZneesGkqJosfQL3yRa9PTymZPyG3u
a880QG02N3bhsqszS0iQzeQn8sSb7SQe/PX055Gqxf9vz3zQ6LzhaNEMRMsc
1gi7Rmr4LqZMFWvKRbYNynq7xVYuUvzSw7b036ZX1tEqKeXCfXNy82A5OYBN
hKgzFLBMvJaXOGQlAqVoNyVhVNlMEcZ4i0hTOM3B51LqvVmUypZ+IJ1tngNq
OgRXxempRckVFBJhZpYZ5m/xaMPrsS6GxulmqCQZxyuluB/VMO9BqqWDWCc0
FwVOU59r/3RcrSca62QJOx6wfHv5/wNPDAd3CJf/y14/Prvko5repY75lcU0
27pmQVZawJlN+IB1OPter9PC9JsbjehahbIv24flRyQXHXJsN7xVl0RiJUSA
5T5oPGdJz5svCFy2EfDNDV7of6RLMHFhRO9Gjc5IBnyIRUKUMNbgMTRcgV+D
WVaQjXL+4RLr2j8bL73xnK+SLeYpQMVfukEzYECG/S1rHH+7XyLEaEdQW33n
SUiH06RcdCgyRqLz6DWgR+99yARDTRY5COPRiDBPmuaUjpmG38fpdg8C0sTN
eHbsV27bFLpH7qlMeoZoAAIJJEy4RIPPjJBwc8d7hOK7J2IPk3Hm/eXOKLX1
42O/4SU+AZk/QPSfY6X5XSLq5i8DlaJ65YUlWlU+vNk4Es1vgYNIePkifmLU
7CdUkBzAuPcE3jrjBTzt3jYQW+/CvidWpMiO8IBEJPo4Mmz884G+qEAUwYfh
gfOUhPBiqMo8QW7yFKSHfnMDAVyXc0iL2G6HQrZJOsBV1U96kdCi1Uvpd3j9
wJ1mSk6PlrjclQssM3tvl8sAsS0PcJP9o5sy9YalmlXBuWXxKcBjkNGDA6y7
QSqhD1xllKKuntkRGWZZrko+pjJuUndHq0IfVChaI55MAxIRbtpt1n81ZZHk
dMrOki/4qTozQbBKbRjBhTO1dSNZt2rPxetKSX0T/S/64hQ81SdA2EmcCCMU
iaNW973AdwHHHNmG00wcjSMqRx8MNQzy8aOX5tZ4TjyJgbrCa5Zizu3oGALd
rCaHgPDUlxWkR5LZId4x9bmixrORL2BGfAQo35U4tVACjOA7qJAraFU5sxwn
ZDpi5z2vBF8GlIZjqDNlh8NO73XADyq5fJzY9c5Ly2z8WyypqdDyH1Vv1gj4
SXdK3uTih67MgKkIGRbsanK8mYtG1M37u1Q6N3bh5rovRYxpT56UfYZLDl6b
prUe7GVR2qUVJdP/GRBzSjCsd18aCGPVJQHtx6UWJEuB5IbA9Id4D+rdgbeP
NNkvGYyI4Jb66jvZGzLTU/6y7t5Qh7rtNc1iAuqt/SOGimKruFuVwMBFnHLb
ujySpS0nuQTs4N5q9NXuBbcD2Y7GDTg6iye/0d2jaq0Yhp2NwuSUrtPEgGP3
9joGieXmpQM2652BD822F7mFcccbDQc6ZWaRP61bg7+p5Xz4IJ8R6q3HK6Kv
G1orXizoFsfdysK3hTF59le+0M0SA/cE4SME7zKOTTk/qUrRQRAtqNWNWy5L
oHce156XmAMpK5u7jtKDNz/wim2tfmkrh28G5bD5WxWt/HWtGKwmlbjY5ypM
P4Z4e7+zMPVGVz5e/FAAVGiFSLcaIVtX8KWoB8MF7oMhr4v0HqPljYoxobmk
cg/G1ehm5tu1BSOf7BicW6Cue3XfAZ2nj9bYtgAnk5xExZyrp20rhD4yeIZY
E6RMk4sjFw66VVDT5mYGI96AbArahElhJka2Gokp+f9nyiW390ZD6U/VMU2G
ymS1Ra5Mj+jTi5Ga+RLdrh8aHW6aFnbFOnSJ1LgT8c0RoBF1xZGgpHHxNd1o
8Oods5WEyCf80FVwdzwfVAF3y5gOZrnb9uwfqMot5GeXX7L1gIfwG8uAlAYm
ILe4j/8Zpq1e8OXuGDCxD/hQd5OUl+HY9dtZZU5noxM0BTmd6jI9rgULXdWq
umLzAeMULqn4hlOm63WDpWoHqB/uAwRa4ouuCJdyV4sMQyY9tuNgFe20Vl/S
bIXTRzBPf6WHRfXWULgigTtSDlCJKiWTbe4uva+uDwEJg05/nDxSy86AtCBO
s8JWrWXhLv667YTkxy3NeW7Dy4ILiZiDNkgU4oSpH9rl5fFN3HPcANit7c+1
yxl3SDnKHCkrzeo0bV+55oFNoDpvegk0wH8S48mWn/YS4uwr/e4PNPUbbkXA
ShGIQ5K7Bf2AyJZtqS49BRfrvJx7KDTUpz6oBu8zQwF8O6VAMubrDKTtmE6E
a9QWmL8bW/XOrnscEJEuFSLqbyB06eE08iESMj+05sJRKYF0MCPnyA7u+Zd9
+ZrHF9nna82u44AsZSlm/PuUWBmWm9VKi8BHp2CsQVCMlOA6aKiIWZfgJL2S
08YJPvX8MJX/b7PBJeFtT91FWysvyLOROtB5up9uOqeXyEDcuU9WQ+YEgUK1
ac42OIyAtA6012xa1ak0iBggWo9yIEibxOjlVHZhgmNhTcYhcqc+4rr0IGGL
LSLmjo9Tzag4vxoemzCR3VRnJUhM6/0wONPEzouL2ImOYTMNff4+n1F5Y2Bg
cTEYuv1J2vLFtpx3b5UWh6tpNtpjsMFqao6DdBWYGGlccRkZCm/9PAeWjydi
x/QLYb+DSORXQXM4e8gmREWSeGlQLav2x5aSD+hfkHI650Cw9nphrozIz0wF
qPjyLspKJ5MhY4m25H8LNEsEfCLNAhgTiw4lP5TjC/BsVLcDTOZQmaZw1mgr
B/YNIrWdqcljjKbGP+G7D4v8IBt11GfIaYM4ojGoSn98AdR2e/oX1FUxkKq7
eeUrk8UhHSHudMwL+R3QkId+EstDECKLVm5qs9+yJjxuKkFFp84ONr07YQf/
VaZIZB/WGackfsU6d3CfzrEr51ceJVW+DY7qWiz3+bmvmSGom2sk6DOGu7fg
rI7SrBL/q72RzlZ76ZtwHIFLeCf/hE6z/Ah5VmwsMbLiL5exlFmBCY0Y8kOq
ebgJnnzNDX9dgKp2y8pDjqV7MtXi+9zVfYpy3YV6hf0WiSKNfGm1zhaWu6fz
RIKdqzsLZCE+xZUg6C9JFsQaaVks7sihSTfVMwnXnirzLlGdM8k6hPLczSUh
O/1ApJtrH06ROGY/itnwoetNiZwoMZPdpChVnFUfVPgiJFtzOwZxQIWnYPUu
KaiuZYgqy5k84SlAmco8ZNejEZ55uvAAMYwQ5Ev9x2UKlk4gtWsL3kLaLBdK
7yDOFi3+58gxkYKdIPI7gpbLVmRXmA2cwqHn/kVAQkaSgt3GzzniQPWeoEsf
xu6UBxRd0OWypCCAZz//k8iugudiIK1PCCsnQwrSgd0ufwfoCbP/0n/Gh2Q6
6anbqmJZ9lcCmGA0U1JgSi15yLbiB+nlu2AkjIqsYGK3bARRjQlfQWYWN9CI
VkoMs0w8cjobxTYmn5JOaxqHsb8OfdeCpyy1oA6UIPFtxY/yem7DbRg1f7TK
2skKQKE6ZA9yHM3NE6WJ/R65BadwjA8YP0ChGHAJFg1q9PUx467FaD+mlmd+
GDtrX4R96+9o0yxa8YPgWoliXvuVCU16ngU3UoF/CVl8TSvaT1zqoVBdb8Li
XIPQ71EVmthiwNCtMU6Y7DLcPouQyO0IFWL5skP9/bpKPHdBTEl4h5Ebnfcf
etX20T89lBNVoeO/FqYveEoRrwddmlYPWsWkU+gcJhq380tzxUETEyAIeW1L
Btve+uu0VQIr0FbHzZ4T5xTt8rRgRpyCv59b9y9LlGlfBzSFxBuQEbJLBbKa
9jf+cwuQ/RoWW2RNrdYj16smcCCYD31haPp7ukI1vJkMmxMX3X8N/3nRwOYi
mT5Al+RogwypOwsLJ24+NXhHeJEyOq0YOKIBoN+KV/qWKqMhqJtyNJbH031H
8sg3kbmXHbe9ontolIogcwdoHJFe5tp6b86QRBrMkHQg4sUx1w1YQ5Dxovs8
xEbzbiCops5MhLBD66+LpRTkv621+JcXRiP0h0qaM+CxCaFrW/iFyIMe6go4
YJ/tItdBfr3GRuiMl2NPyufhHZe99qn4RUSUHxY3PFDMNBwMdz0boKuDNn9Z
UZ963aMNDn7zBlBL7tsaxqeWoIYaKxMeIlhGk/Kih3+d8z0cqdIAeKH5k7mU
WqqNI/uvDsQGl4+nlxOUgDgWkmdbge/wZqUNvmGIpcuX1rItRSdAAnQdEhdI
gGKJf3tj67hFHbCa7bF/2JBcY3IE8f2aTdxYon5MJ7xAOD+iIvdTKBQBAGjl
DeaPLtRHBgEpvF0+KpTZHIg8ilRdsqDBty5lFbPolzWs/Gvl7MrLLd6XkEHM
7V7SithxABoUZ8f6HjnatD5sMu4cdBqTj/Jr5fyokiUgG545yQ0XL7D6ciYn
vSihoB/j2y8EO4/J91D2MPeK1x3WwnaXRPg9rnXfef9rffhKjfSTqXDa6M/9
337lHUQjpoMbbBG3m/ozQhySzlFn4I1nQOIpNv1/TWvt+M8fQ4qsjOvdV4gB
04J06UGi+uj83wmUZZAs7gUV5YJRz+Ee7TIEiVXr1V4k4yrxinunHEC34i8G
dC1DioVw9EqRvoQNMlVYuqTCJejWTj4qSCylZhrx1/Py0nz79V4Q3srHg57Q
cF+5CvCisnYJFJTMxhkB/zUbexFhDf06nTcr9q3r8QgyoVLgZdRMGu1UkJqY
Px6HmGymriDbSPd/eEBJw5glwJiFHdmwS43XKKEyssHJ9XmAEht7Q/rEyJf7
azj30U2GGLS1c3be5r3oQxIinD4llRCUCj787slH47yuOh0eXormfKlyr3MY
YXt2rdvW540NUEIdixqyMnxLOlb2CoVbFlyihfU84Oi/BXJuvvDrrPqHiwEC
eVJYiCvDcmBNA8XCIABv/Qp4YiNZskZ6Xw/tKhQvbXnxsVtX37UmgIInbdv7
OdyTNLXsfghAubEpU4Qs6iUJRS7Zs92LYP4dbt4K4fDnwopDR1yoztnLQmtF
rqekFtfiJARUL1X8fyIZeBOplIvT0UG4Sd11NPoPHpJUIFd+UiMqT9h3EA9h
k18U62dgzwop6dXxM6WwI7kAWaLfNLG7Ut7QHVZP6y4M047ziDoT5xOJ8qO5
kGDGQcnBSvhwjIY+0LeWtRB7y/NBEcevRmzwhWRnug4oGt5gaWWZNO7+00MJ
TmKUePmQlOfagetK9KFkiacHbGkrrq61xULiUlQTUlFUnencs7+wrVuXyHTd
Ts94HKVZeMza4xq2x8fFSVxzjSNwj5IlWg+rsgv9JVhQ1QGQbEb24HnWYyY4
MMysRfH6k2hAj8CFpZmMp+MqUW2LvgzlxOBJHvznXpQd3Oelxxtc+wz+p+ey
AWgcuRLjAF4fRMUnOnN6yxIaag1Z90Nb46sCrgRWLn0xIhy0350ngYglHNS7
1YK4Nlw4C88WszNEwJ9Am7+X2OW8z1ShPX8zyBmZLnsR1noYxSDmEMyCKSxp
TlmHIuACUzNBXfAkH8fMziT9JTBXF84TrTIAo9hEPmcjgKyBVR/Y5z4s9DfZ
ZhjbhqwmVqLe16Q5OYtj1pWYcF+/VVAJPiGQHE8iJMSsEChTsqx1kP9WrfGb
n5lp+C+KLaGILG/doDrdx9hA50J0TWk9ZMUpDlKrKd+ggAC4WoH3qX/eFTw1
s3Y+zFeabwfyE4RGDMMczJnzNBRxkFaT4E4V1Sa6PSFVl4xZ8GXxRzSgNmta
2hgApWGDrpOUN5bQb96potrdTEly4spJAClN3zo+u58xc605FpuEoFaM1tp8
VndfAfOmWWT9oWiuP8uLFx1win6CxU1WwqxcfLLGq8GEDMxN1Fpd8d+wXa4+
yTFAWEVpI4YNMqpFY+JhWyg1TxgOF1SqQJrlqOvXm5lweQvfiAYhVvzQ6Z5Q
AbaSo5etMygYOpax9nYaTpaXSa3FihFjPEjQv7VplEOJEs4qGx0IuNxjIqBu
cO1CrGNulqcUGEqMHMcN4qi7ZVGhvWK+ABNOvXYgpKk4Fn6MoMIxlfQEEJK0
jTWLAid6Pr3svpiIqFfh5hC7RJK6BLZ4D7DJPtYNygvXVpSzag0LTHrCRv9C
GR82EVs2IsuozeS7VYZHv0t6Jtx67b8gmwMoU5v2D9mF8MFVb0zmdVb3bWel
Dx5hy2l2+FQSnKznIxSjxHrYPMSJJIUqmuDSDMGuqN58hr0qzVd60ft2C3lf
OlCPWfOGMVv+Yw4AZuTKusL7JrVb4p1JRKDwX0IpY5GDrV6Pl3Mv6nEkASsq
nof/X4IkrQKWlOlOFUuUvUHvcESQPd5pNBzE4S1M7pYnmGDQs91vI5kuTgWH
q4Df7NzLFfXWmQH+t/fxE7mInt0+NS2Za8aKdCY5vbZh82jgAHTUO6G6w4aN
boamJN23IUzPQ0ED3Wi6NqspSyxDbcfvtM9aM2YPlOkhRquowLEzR7JsFmmX
ZIFBX+27jLeKmnwOcSIBlZ66YtGQLT/d/vzU0t474oIJiKlkvpTQMoBWcINJ
Usa2zGWF2Hhp+9krDX6pqKOBckSm7quqbRCwZ+0N58Yc0+47O7Um7KBoctpJ
U1LVs05fMgAwj20lOyev73dlkmcroIpiI7rpnIZ/E7MpbvH4pWsyK7fAFj7E
6TBvSIAkmTg7x4tsdeXbgJVCY3RiaLA4o2Ras/lgEZS1PFv3lvbjFhQjHDv5
fSYK5Eo5xM68GikfE5RnFCUNFFqfTYq89KOtfn5FYUWEdSWkLNlEinSGlrBy
rkx8lCXM+QSRNADr1JzKYBZuwmNBxAX61BXvHSSgXxH0R8mI2hSzCGzpWYiD
yso9OZrudYDxqRk1kiCI1K9ASymN0+KM7XJkaHotCOXiMlDPdDl+8ySywrRH
tsWxu14ouVx9A9O6vvBNsWx7FoVSCUT3HgbzL/VHvTFgNo4Dn/nfCzHXFQu0
q+DYhQzUxeR3gKiqnFXqcl1Hu6vl0dwW15GxWEM1si7HaOu1z9jmJKLJEQ7L
3Kfx07tva5Ay8arxekyMbYZgBTDLaidsTcUtWQG6A8FUJjCHXEwGgENJSHa+
+mZu2aD9rhxBGYp0hdDGYDEWz0PDppCHVuq9pxJhFOtU/HICwOgEk3ZUqzz1
qgb4xe2a7eJKVl+ztmbAfmljiOWkL8DTcmgb749iinPnp1vvI+YNFmIgsqEo
6OR4vAB7xCSkCuiDMA78FTvpzUQVKax6nhkDUgAYCaGzryTX6OvL5mUAzfb/
7pH0QsdRnZNwN/NNUM2CY3/bdW7+4Ld0b1XMmkwOetq10SxqeyOvn+sdqysU
xVbcxHKEIaLNHGQgGfZRGO/Pj52Rs2NCEbLe8MqA9sCwkbYN8PKz3Mu5s+hf
c8x0kP+sRxqb5uYI5o6wcZFKD7km/l4XFkHX0sLIC2fczV3r24T8ctV27Lxo
9tzARO32PbtB5d7RSEkqLlGgi94NHwhTLjPrtjeXUKkJlimjZplLk7Tm5YhW
RGNeW5UwmU+XmyXJTTpMkMMYMCDZ9AIuD+XpaJfVWYCfWW8Hbuo9iSDAdi1w
IRq+Di5HAKqY6++ciLcpQWmUnG1ScIWOFfTm3MoVXPU+C/BUyxLenHlnF7Cr
0DZ0jmIHxdJ/L3BvbFmxSbTJpdklFE7Li+Pikc6ht3+xAeLQzJFd+ncwbEtF
W8j8/3xSViTbMOxG5TZrFpHKi6TZ0k3t2pNCOi42zyAWDAPxHs9FWHEk8cAY
OJ3of5YjPA/zU3lXJg6JO1ydOsx4ID23MpGtHC3UyGAV3yTVAYMlda0V7nDL
WOZ0XO4yMSGr2JWTyp64wnuNj9qETURyou81+HNj4wiw7g0ptdVleVeXuGST
dkF8and/kLdZInVE9+aWfidIkJFSl9j8Jk9mcPmeR3kG4r1R2k2LnpAaonaL
hQOFOa7ghe3ot8x5KDx8B4BNuBnzHHNnqMvu9BYELptH4gy+UQanW4SqGbZf
SjzaSE0hq5mT5v7JtoNI4ORdYPVZAAkSlwgqgIhKgkVRLp5cS6H623O6ds61
A20pZPdU7t6/0yBh819xdNa+GD1RJwQk2jWuP4hNm9kc4zL4Tsa3w3dhTgbu
nU4AAQXkKe+V8Y5TxGAdVSkzOgZoAERGm40u8faFLlkbpAPeR9PJlVzXi29g
PLnsjzQKO5cxJJ+LdddMSyCTVii38HvJq/0I4y5hjMEJih6c+05ylJDgWu2Q
Yih3wiWi+vPZEYh4xMLLav5PMJbmetnN9DQEi8AxpHBiThjeX6HUshskNkZ/
OQ6NbnY4B75j8JRQR9SKzI0sM85vPRxRnx7hclQmsr7Z0B/hSGeDni+9eiFl
4I+xCq5K9wp19lr5TkiWlr8oggQJ/Ixq3jHZqbQo5KWGLqXs0tKDgNY91kxW
rc5Z3wXTFKKcpgXfOn6/rsnM49PbiujqzgMIzuURBq1NuMmTF9k0oCz0bgJF
MyuiVGlttFqlZULJoZ6cDsk6UdXTU3nAltYfEL3dCw4YSJOEPrsAhUK1j6VP
2mQJsv5C3wYEus64M8v4YrTif8iEMZjH96GDgwpdoWJLhlWhjKIdx46IhyQQ
SpII7kyJJJk6hDwsQKyvJkK2UpO9UZ0HaTsng/ugjBUaNtvsCYeY3gRBS2+X
QwK2084lR7HH6Xxq2nmIIuOb4hN40itAfJ1Q4xThNaO/ABVVauDeaBOv8piM
naEbRlzbMG3/K0uVwIkpzkQlt0/OaajsQYVNQq7Y5HAKFEmCU5ObVFjQ3RQg
7fogf4wbeqVB8cmn+ozJmJLY30bGbaMD5fSV5vHGOi8q2qRvTmw46jyC7FMu
T37IZLrU1XHX8nZCpkjxsTiiw5/8VRaJyu4Drl6GZaY1Lmh92jhe64o0mZnL
c82fEidBNhpCXxSaD7iiKGbayBklYR2b5T9ZnLHX7aKHuaFuz49XZtSWZycv
sxufcL0FFzvBwAbXzM+KfVZzz8RR04uOrt+qMoQwJMK32xGaPnEQAIYM78oE
OGKvjzunGGcuaI+LWd9N7X0QS4FZv66fyf+pOWP0O6sGEB9APY9/56AlgQTN
qs29g2kceqENxHzjA2Yrh+tDW72+aizBlWtUF5iKsWGHq6h75zKHUcWdu68l
WF64ICGkp/GJd4CT56ia2SCzN3DeAuWLh1HgX/Nl/ckGPAcIkIEAQcZ+Ef+q
OWabtjPv55eBiqUwRXr3nGUVQNrA+9Z/TIrun1/zjwTDGJNDdfoKbQuBTbDt
F6ou1LRGjFirkhMEor6Pm7qwAcd+CZ2yo2lBzaCZRxDCJZhVd3t8MotdSY/F
WnFtA8E31hW4OHApDevIFt8tv8JbzND7OEkF0VxiCIWgDuyNf/z4wXlrTJnd
Bx12X94JP30nXHViI5dTH6/n4VxZIkI6p0U992lWSb/R9Ih+nDvtIAWtj2Vp
wJheRMYTsg6Pdmctrw27aGjc/vG904Jxab2cyzo13XGVXd06MATbo6w71Mig
NMoK4LsTLMFa5TqmaIurSsYbz+3uOyhhWyCKITln2D0IITpcRBwEuHT6mET2
L/D0dcHEe1EqHWNn+82CQ2hOz4NrKvIFdpLWhS/KbHe3Nk+TDf/x0KdPK38J
K04X3jMC5j6+JOt2x1ZB9ON5Lteqe1ShsipV7O2AWF4h4fRYM58rPa7q9hMA
tFB7AAxZEEbzZsDgm9VmcvrjgyDtbI/uF/4jPY6iMN8HANWS4DjUf8YlYtwV
lVZEzPyCp8XD0N4njfoCtsnTRRNTUbTZyIV0SvtVZU4axkmM+7OSHkaXNEBj
u+VDWJrfgBr3S/n5ZmgVi1Wlbe4zsMEDRnsWXpnnroQaNO1s3wEkUtD0kg62
H7NTb6U9bzoMtU/mIx8tpAGXVlhTDyWeL2Iu0yfZ4d7ol+HxHrtvlQ+KHvvC
ncjX40oOVccO0z2pR79d5mXy5BuriYD6Xzvk0KaTV/r2Tvt40BQNSuXMQ4bp
/kgwO74fcJDE/+DCmfyi0tJofWJw900p9PIC24WpjQppkkY27LVHObU2q39+
BDDOr1xi+NWtcIG3xgnoB2WcGzUCEsDX6a5kZu7sliT1kDj/XJ3UeLz0ZGm1
uIrD9oWMrZ6+V+jvdCGRHtEsUPQGNTPTPSJOiZOqMb0YpWMJLb56V0/6mq7l
/IOG0Fq1UZ91cFxaylHkNsYzrWgu5lLqzqkbnSfKLn8h8x+4lRYQt1V/RMjW
jrQxEiXdo7fZ3xNeZNf3JSoLbtAE3dfO2BAdv9BmOM8KndhzOyDkUPzVFuJt
mPP6/to5O/GhuDk8UnON7a3OD0Ekyxtw1Trk02AGyuIWuxuMyhTwGdVqp8vJ
VsTFY7lEMsaWfgCGt0gPbEn39BDpQlgVNnDZsZI2i8KczbZ5sPuOocavR4r3
V1AVgBXoUX4JBNB53Hw+PwJkPIoV0gwI16GI20gLJUX6kECY6epESY1cVLs9
yXjHcKJMdxc/Xaqv0UlxCUfXSo0nyxxdy5879EeKlqx43zT6ZORQ4jg+dnbb
I/MvUznpvqlryDNgwO5O24iOS9GNjrgz+B8q2uCPh3ppNcrcrJ60g2UtpeST
n7vppMG0m0gqxFejRZdGVR4w0OaaQYZdeuAq5CUB7iB2POUA5AKiTtQklZXV
OnCbWnzToMbo7GlFApQwsY7CbfvY2BmBvP1e03zdOZnBAotccijVSfh4siuL
9QJHv+FEZGIHhdf7e3uW4VEmttPwGVGlAQ0YtPbIHRHy7d9wLAai1YSODKBQ
NZF3Q2m9322Be+ySHQ4wwmbS/MJAfdHKDgw+DFFetqRgawy3S+t7upz9wgAH
uGrBcn2NrWKC7ATyQQ/gIGh/HH2LxFX/Vq0v4KVcTrNjrh8zwvGdBKeivqhc
ro4lVOC7YVZd3ILyvMav7tbEXWp85hcS26auDpG1mJBgAqYezYGximKVR0ep
8rf6LJ/IjlqulaoZTc0bBgb0U64rquwD1n+ygHXYieO3x+KY+cx1R2BQ2aut
6oeamVrUpGiQD/uEPugq02MZsSiBnIs6TnsSq6CMUmpPSCfibVKPFZc2+s6k
oeTVVz8eYlbB/wE7k4ufhFGKsI86qZ/wYdihB8aQHIOfpfJL9XRsvWKhd3jS
E4A91XnZS8dWUnwyi25/VE6gQLXTGp2k+ufZxf+MY0Ozcbi4stYhaNNIJEWe
7KSeSWxJdYV7dFLz9Mm64VVyqcN7E3L/dahSBserJ+0SSpwMh9hU0eNFij61
+qydujF/S1052XIImk6Fc4CJ/SYkQ+L3bPNA3ChRlLqzw44erD6OKfjlhEsS
9l+Z+uaobjYUxyny7KT9QuT5kX/B+FtdcveA2RVYE7Yg2H46YCPB612/Wk6k
4KUkYDe9n8nPO+FlT3R2MqDggl2+gavY76sE00VMngin3Gf+7zbFRawN+mPH
HVR0C7VNUwrw36yD21GPCnrQZVDq+Jm2HgFtXDbRryuhbvQVm8ObZylTzmzl
NEcndaTbi1LQ4os0fz8QZRMG1hnwyqJud/y2JOpnohxq4qqdVy94TMlSKQ2K
FG38IEIrmcfw8WVhZNefRkT7pRfHb62sTTHowzNz11ew8Gj7m9nTIdobpnYy
NIPF6SapZMmBaxyWOB861RFLBwqZIKRli1FxzLSo+6zk2WhQk1Ju7tI8KcY/
ArKmHF/ILqbvQUdH1BkMRjlRGC1o3HPot5E9ufM1uLouYmYtMevu8TDIHKUv
JIMNCezgzdojeFr6DPtfgpnKI6ZmQcIy74LqSa26/LMT656yoXW6jZ5gyX72
UPxcs/NaPQgkmK6DbhIlnwQGvLo0xW1+zJEJC+zbt/oXy1NafCjkOt0a5jkO
VJy2wYr7lOaFkpmjfBS/pP72noJgButmg+WEmNgO1Qp61pL49lSq7QYONOSw
xu3yNLnOgvELS9UerqBg6ORA4DMT2OKorXcxf/yFDtjUJq+IgzA1o22A9Ztj
wHJvBrS1Wq75cT5vMucIYIPYsTrCun+H5gW1SZwluxj0VMPjWgTuzsKyrvTB
H1FUM28lirefk6BQ1bhojTKIo7phmbNN67LEGu/dTcXkCydroX1Czg4o7XRG
E6cNuZ0TRZxP7NSQUDSHudL/L4nM8B2ArG80o/HIuMiore3K3YpXZOUL6495
9qjnqgztoQuSyswqQi76hghxQfCQTpsTGw84EKNAVMedYnAWjFiULBUvO6Da
eeIJUNoni9BeiTwKDKv1zd4IDeBpOw47hJUjoZ0OQjpL60H4JMFrt8NYtGMA
bOFW5LYnNhzSMRQqcEmn1bqnBFUhMEiCzdL0SCS5jtO2ANCJcqWjeZCP9jNr
yObiQBzOy4TUXG7CZzeKYtRFHJvzeUNx1/eEG+mJmEdJqCK89z6HKnl4IgJ2
jqqvcHi9Ng2cg3yYjFKckO84EGNY6e1zp09wc3jV5py1YDx1+bWIbXCx01nP
vlvcRmbVVYVLtiGg7w45qjyia8ZLDDXB1Wf39o8T45CGouSWlqtzoVQ9ZcOU
jx0iV3vtheZ6S+aBg9fMkMWhzlG/eGQsGXJsf/xYBOKJy5DKa1rrZRglpuhf
JAGyrCyoczdRyrsz8WJxSbNwgP5er3fQeRqHWHPkPape+w863Vd3Rb+GedUm
Ivj0IPXtx9oAyxCbSD43A5Fyk+GaM/nkc6602SrM52OQeeucxfEYZEseCb3O
50e/kNIjcNbfu+d1RKwKwFmAiNU0htC71YbaOhnM3EKK8zcz5FUk9/TUAS7N
cWszQvCYyV0rmPVs9zeeh/rcwOmx8GssRJRh0i1FnCzUPGbvqheqKmjd9osq
Kde6PnQzlmyK4IUPP9bJM6JOYTaRU2R2WVEjYsbURa6d1RvSzQ/PaEQFL942
BsnKGWdXpHoYl5Qu9cSe/iaQdPgYKB8qci3qNvoyY5VhWnWRXFAbBQzt9hpn
OCBoZe40zLePovQ6tcHCKQSiV0ZRg4IODzWnvyf4dyqIw2O1Ot/5rMhybRaA
WjW2d1sDzoIgx4UASqyr0+k8orY1ATPhtx0X5/ocH5HpxGtxBqSfX9j9BfZg
ULz1+K6riJFvgJ571FCCppDbRrkcrO0DHyEO9Kxy9CC+QyDaIPSUoqRtYdLp
up3rYJTCbqnToczn6EiiGcOnXvptyyszCXRt2O6g811zo8uEj8OEX+JFe3XO
PW0IcHYk0XiGOXduaNCct2xlkAdRLZQD4FWKsCj1jKzxoBkBS3RpAk8j40k8
cFXkBpdg0sVGSNs+OYoWzfr+lxgjQp9FaVpgXrmvzDOloVuEFblK8xOHvtD1
79qasr16UdsGGAkp+GY9RRQTAL7hmhunfhYyuPzcXWWi3UFFCHBl3FnDWj2G
0kwR/FWLDVpKxmUIL3UV2IC+SUG3eNhs003igC1Ivsdoid6Y1V39TtCrE5/k
33xazxmXmBXVrPbKuG3qNOvNkg9HIcrft2om9C1aEhphR+sYAdQbeFqOirMP
HECmn+fq5Pc9ye/J39HHWwkSIo2gqNq1omFikH+ac/FdoOnDAAyfZ5trN9dA
02fwx1QRlGD0bUR7LgKxirNWW5szsl6JQqIS8hQ+6fw5qeieD/B8qBAUsFp4
s07WqjXFP9e+z7Tqbwl7SgemWzeH0eZ8f+IsLV8iy41Km54UwwkRQZBDojUX
CFZpTE9vl92KHZwsL3Z+XH4SZQhwBvGDftQGlhWpBUEf9M++NVnMGBZAjUNp
I/A48s59I9XuF2cDTaJiU6aW9ZXmjpzv0h6ZtG8W4rnbSp+8Gp/9xzoew8xb
r97O7sjlV42nrDOOMnO/FatA5X49/5/DRnT6g9yTXbUfPsmEin92qfJjheL9
/KdAfYQe0403Nu5m2pwisOQs8cEImzl+VhBmFkaYkq27sHIrFop2KXMPT71n
z/d7M5TjLahg+9qV6z82elwpY3AREfGnzfF71Ttqz0+QuBm10i0prOTGnfEU
j+znN59KlsK5yGcwVzQECqUIiRRPjg5AD+25uhkCAkNjZBV+dHNrXlt3Q/JI
UL3dyZSjJL1BBeyU8SCcOFIVMBWeGxEHtM8MVbN06eSwKFcd11nVqOqwldqY
MF2XFEmPTksYwkVsnpMjo6ITpsnjD+5QnUebarETf80gfZsZaHX6y1sG/rIm
IyMCRdJIAuGTTZbut7XLhLZLKKbf77NlLS4UuooR0fkPCIbyQ9u9S55uGy8w
9ySIKNS58S1f7DW9nR/K3IxKrP9DO+I1IAqDhj+SoBjN8KZQ/6p+5xYcE8hx
Fa1oZ0bDMVSo24RhOkyybjo8xg1UJ7lej4wEpupQPUDIgKM/bwXG7/eA7sNa
a9WBJuns6E7zni/2U4ZwZXIwYvs/tdqQAI2N9muM6EciqUfJyF1H7YxfvakM
I7VSYJxVbsTfCdVzRRnisJNxoBchlqrQA5DkSXQavQS1HCoFW15N6cyHfKOO
UiiG9Hbt96vS9vbTeVHeyPeZ0xev33dm1WLVLYaggpEGuPCBc7vexnCG2JCI
8m51HUd6Xf04r3clm4Z0P42q26RcFoIqTZjS6ar+Pqeo3TddZt03sNKtFnfy
avWX4V5duOEEiwLxBAOx7K+lTiErpEkHQgdUpwTxBKYGD4/ikjlTOIMKx0xb
to8m3UjsaBPEyJlM0xkJAomnn0b5v7okyny/laKmdgMCKE5Bj8RxAGNKBi7c
GD9kHjY0WIgBv1JCLPeITEs+SD0nHw4mQZiLfFbAHoR8HDrthgXCLLShm7MQ
qQarlLtDRSh1YDElaEZTekFNWPzVMe6nXrXaNPaIpHFv9ed5/pEnMoYKhCLc
QAGLshHNlL+AEO2FyGYy75RThPeXqU5AYzYsSVUwsyh9Vhxrt+ks8m0c7YVN
HfAzegIOKEd2KAVzvMNE6WFMPSM8200leD6+fOYbfKyq03jI679u2oQ2WRFA
YJobswCk1XHhlU8/b9sKI9mTJjVnTC+5i5Kkf7JCpikpTzMP+9uyfLIGVSxw
mMTws2HZFjGUjHkK+wwhugHlmRc8bpqykCtUrdyU5lHXGy3dw8fKq2DhhTnP
leCDOfVuse0sPug0/BgiABlcaqb6ulOQgVHjZwVm8UsLX8wdjTpaRecqjn+8
gMrB+dStuegQxEWpAygi9vGElOvfjmDizZWNP2RF+292A8fimF/6fkeBeh1X
ALJCz/YH1PJR0uyhBLZvOfgpAh+EoAA1AgUpG4kQ1tfz/s9ftT3M4bGbQMbf
UMXFVIYmBo60f4XiCHJ9MQs3dgAPo0nTHBXGCZuR8k8vaux4AGROkWnvtd51
WmyFO5f+AdHQ6ke6d/UGmKV47vRoeacieyvPa4GS5/rO+/MKhvww/f6KWrKz
nku3SSdb5Q3oieUmSCYx8QVIODHelioO/GJawC0YYBrGvy9N+xPEUigR4ajJ
MfREFiQrbCEwQ3UM+zswhttZkBw0v1ZMNtHweZzjl1AW7v1QfFC+CQu+9gEH
CJ3dUzNncMMqWls7ViwHh3ws1N8L4SeMBM6QmIynTmJMPETf5yB7gfMUssrk
/qAJvaZ50AqP6tXPeXtx4FkVJGG6S8UcRFeryianztvTUQ7bE5ijgg96ZQOz
KI1CmP6nUNt7VlnM6wHUIJFCwIxf6JsJMQKY9gG1c61xiXepXy41PZkxtN2Y
bvY1BD/rX7cvtAQnMboh5CJBeQcTNjngGElRIfHe3f/DAZGSqlmLdeXenUyg
b1XjCK5w2FRMrgxJja1xAypOgt1JjtceCn/7YuDp73d4lVcPz8jck+0DPMML
EdLnc896N17OpJjPDUnmKMMEMdPN3Oq51SC/dGDqML/LbuWyKv37YahHaTJh
Gmmdhbpho/uBfhw/jcLVoQmbdQoj99KEfHSPoKgczq5gJl6GIcByqRHChDnr
oRapxh+UoFJugnpJc3ciI91dpSbiNL/y9q2CPovKgXRBpjgIgAma73tLGKaD
Kyl6NsOMrEXSLjAsEZnFVmgUTF/FeOuI4VC7vnlYypVjyU5T4S5esW/zIW4h
ilv+/rUBC2KkJt7Hy0DGV+GPfa7LMQo90CxzMOyacEnUFX5Hm65x8iQ4JIES
yNQg0kH51Xw2cSjPEIaCiFOS0nhJoio/fr75+lv6WByBeXfgkalWmoxDxM84
zmX2SpgygO4nhsqKdLm7yzKGVCwX5/dOeF0Xa5CWg+YlLEFA+hMKbP6zH5vD
NP+YlhTWqwSf5wPu0a0w2GhRHGwhBzqU6BcNA9l5o+skaMWF6e9rdRzTfZf+
BvxtlfTo6sBQIZnXIVBxQnadaXoQSlpYLIt/wAb12f629yvlWKUDlCklYwfo
ZYpNMv1CrrWxkXf4Imnlduo8DhRDKzxZVnGRFVj69CBaFJCqp6GuRXYDZVtY
PGT1lAZy7TZ2EcuOQooa9w8Li7DUn87/1bdhAvRlzooV/Dr+Qrn8kiv1DVNn
/bW3X0NXx2Q07Gd15JlM/4JKUhD5SNfRuJwvdZcfsIuxJD0LiyKGqJY2+R3c
ouex+uhnGt1x+qwn+phox8cuuBCZYZJHkK19TLmqLg+GLxrPSrP4GdFA0eoq
KpsL0qNl0kuXSjU4MoMgVAw2oal3+e/atigh4YEL4MebE2xC/qGrIH8AhcDl
UxeBLCUNR4eHMj6zpdcJr1K7aB4+iN/Of0yyn1AwBMGA4Aqq5TFXpi6cx90Z
RUp054Pnlceyl5Xma8WknGpN29UzxG3aXI0ocEeb73/5afFb7W9YWkObLl5D
gcCYaHbTqigCrMpWRg81gO4V2d+0WQMCnyrZB8yF75HADqwBVjlwu2un2RhX
LsbrhEzYysJh2FiFF2eFm/E/rI81VmhQVtxEIi7NGXquNTTqgBQA1wt7axPN
SU1/QC3GPXhGjEvZE96rd2P6lVYHAgD9VUbM8SACWfOatbVEhFS49ErhH4C2
4w7jAzY23SXZzMQqw7iexvFTiiiSV2/3178wT37IRUqLheR2s5wcDQE/T8I6
HIXBQeYDuprBrsAMdKeGuiNrjkFYt5cZu36OVyoZPlY0i4vllqOdv8wNUMW3
e19nVjlOJnFQD0MHqCKE3w1GJxtUdu7ye0FFLk0DX4dkNwjtGSkq0qC7aTDm
2opcoSI4qBI/lFR4WUwyALHY/lgeRYhUjVst0LeZCpjIvxNJh7EjyGWMTZ7l
oiaaq9Y9zZD9I8eLBHowXGWIGj9oVeo2bL7ZMV4c3SzI744d5Xr7dTBcWoub
llw8yv0zmJSW4QlujlwW3iCEUs5qISRMaAH1hZunEudr3zl1IvReMj5bKZQW
CdSJypW8dXoyENX3O3LtOEnpTLNgraBQm6SLHaraGEWP+vfGInfg63SK3Hro
oODeV/wK2jMam5sNL1jIdZxpqkfJvjxvO7yIc0JchL/3MyBrZ5aVSO/UKcmN
Dvl97kcSykgd7QdKKNIRigEk1uqXGMGmJtGI1X8GEnjnh/LnqoyweUzNNjIj
kBa9enWaPI/PP3ovXgooz34Jd3EeUd+q4xQnb30mVXIKVg6koCzWcu4tYFt3
NjtmZjtPfJDjAjAVhiJ1O2SPO2rYL2eTYQiQLKALcF6sxiYvacUzlUtkdp7w
vVe4bH8yj9+LvPkHVYzFmWY+xiM5eQBw7VtGr1xrOGVKp7xqtWsVMa1foL3+
vhftbpBe08kl0HBVvu3Gkn8yGW9fTK/b65sb93SoCK1F4SqXvMGPmPZZo8xL
a7akMm7Z93EEtq4Y9aeNE9amXt9DMaFrwyuGZDXzEZNtnsNzcS1e+oQ4ok1K
A0l5MoVFPSb7LpAdDTKJ3vwmWuxQW7VO+OzyUfSvEgN3AvZ9zOIQLSIUfB6l
LQxErmn2TLb1Zr0kcPNYgP//wQSjGM6pL9r54T/tXMMt1yKlXeUE31rWRmi8
Rf06vRaxweAqP10K1G4wIYRnl8vphTKsm2tVNPOTB7xUo3Abx2YMgpBR4ltJ
2pw7lkWdiL8eEZ+DQ5Rjrz/wTlUeVW1DqK8oqI+EOzBj7DTSWNi/VEL6jYu7
N2yqzGUvPkEW8MBEs/CgZubm8qT2G4b85LxozLowHyVcous0grral+87nsTK
JUoQagg8vQMLfAr2JLiswy0IKmL6rJSJ24lNRf6QfW5oz5UxGrERp3mpK+pw
gffR/2qGt7avfNd2Dr3iHVCrBrY1ESJUUZM0H0gyBmqb2CxInK35QXEewQ70
EFkF495NHSCOKLayx6VX3VCza4fYpFddMsyjT0g0SFFERPhw1dD9YAmkJzG2
jVpyTFS+dLPiz9AJByD5DHmdaJofECNM0F3ohh8hBrZTGU7RTdohSLtHAvem
uKbGpbORO3YF2mqjOKPaoyxaUUk1ei1TxcaKO7T/QV780HeOAdXds9Au3j9w
uLCw+cIQ20QN98FgZrXG6jdy+jY+6Z3LS1ufehRm7WJQm0WX5ncbikxmT5kb
lXeklEh8sXlWmd668MBmSsMCkV4tYo915TIX1512Y0/4agZ0qh2JN4WMVhpJ
vgyesu9HjmFgxFoxj0mP0kV8u162BgYDvsMPsIsdf7l60iaCCt0saO8P3fd+
H/FHrVXnbq+D6Y2jPVB23Ui2z3KPMt42iuwAeOmkm2K2K4owG4KHwBoWK0LN
0O0++ana/R4VyDjwyu/ZwsOmHvAvDP0I+R7gV9r0O0yGqXr/uhWDyX2HFrKS
VkWRenjTLJRusYlw+yRae9tYNRiSM+VBtOK4g4R+AVOBjOcxUEuJw36hEUqk
zTbKhOqn5VVIbgYdMv1ZlylSuCfY+3WL3md/7a9teIrjIsqIMM/IHDvDRJYK
4ew7bEyf3iY1n3ONWqnlmo1yMnQdsszRv622TUk4a0wQMA+w6tps43vARY8k
rRdyL6WCnymzxGsuV+/v4VQ9xZVH/JNcG+D+62KjzUR/GgVcHL7bP+XvSuQz
RO3LGIPuMvAV+Lg4aguGF8BNE3UdMPLyZ/+OudCEJ97OeBKAw9JHPpCbRhqv
yCXoJR4N7prRubRgm9xLLwPfcSQm/ASmZpNy0JpI8o7WbEbJwI/dHJbsrEB1
UBk+eM8aj5Z6TnXBQt9o29eLK8lFnyDVV0cnDc0lehNxoaTaq9z8bQcLr8vT
LBAKPFA4BPL05qdj+TyVrSMvdlafhIQnHx2V597t8Oa6xd+pgkTsSRTV+Yvu
4J7uHjpSwqGMnTAp1f2MI1SPgVbIdD/0mPSOYit9zRzLZJT3g+s6h8QrB6G7
fkYeItA7HN5hYT40j9AOwO2akKYoG1at/j0EVx2MLgCF8CCAX1evbaOiQxRa
l5+WXzxOyS9MblwtDhJMcYCHXLxDfCWg7nfho6JYSmXADRcmb2D4qzzVmorH
q2ce+mu/+lVnDAWQZODhzhwmaOcfwAvbEiN1HCWzoOeFcewRCRMP+MVnTXGL
qVm06/zUOyNtYpHVlGfntwrsTsSG18r8qi+0putvVh5SBgbTRyBZB3c51nFo
DpCyH69SdM9MJlwJL52u94moa5dHWMyCsMncndRO71aXjYR/F9YOY9hW/3xI
EbhBJutC3G6ZPK6STXO12rn7TZ3ZAVpcKvMiHkOlHQlBEE1pLqRPywmWBx2D
c3eKF3NOlWVHBYwxOZYyDxShtd9Bq+CJiZAXogplM1flGDvYdsBuBEnSY1xA
p1htSpjFKnPbkAfAufuL05tskPzhEDNWce1LQS8O8gQ+6st/E+oc7KWcvpQy
ytVHnEFotRSIWEfVWs8E5Jg3romDRV8Oc6mpG2dAPA+LvC/WuC45E5DMvLL4
+1IFyaXpRhU8UY6Rb9PLVMIfC4gdTrS0Is4o06EN5ODsLF/ffbp/EtcOYZyD
Q1cTKAHK0KxxQ0nj3L4MbErI4ERQAkElOiLvtL4QUE+pAfywGmMvS6blp1yj
6gF8DpVWipJefVjztGS4Mqt6gwWVDa4CSLEojx0btz+NVFdsrIIcdiWXyk2k
HoRT/BVJsvWX7KM5UgVZieIfSuqHPMt2rS2O/pWwNKhIXTudd647Y7E22hak
XTLvQ/N/9563Ruk4bJo4Y2DH1tZpE5Kfu+p3saSdBEVm7DbX8O5E5vZYKFKP
qbCvW0pKCCHHri4ES14xvZ1NBAO9osPUxb/AB3YajHQGw74iDqxZXmZ2onED
BrOWT+Gx+R6NPHkyJJ4u5GxApBgKvc3Vevr2yhmzQclw/3a39Bb+5ovQ1yN9
dYY2cjfX4MVG3LD7G7OWg1oqH/6pXq3/0Oy6ul3b2Mnb9XWcEmgu/5O8Q5g/
3cVqB3c8KpiEFP32ybZ7VX31a/PhnopRLXNxP02ff/ZIbBvQtqItLofRmOws
JSaZBNq5Srdab+8OC1smb8leT7/WqptEKnRxX2thp2VLaNpyG7OAgdBaJOPn
/OjlRB5eZ9HiJ/8dQqSjVM7JZF6o4Z/IYhWN5QDklxBIVsHfzQaCO4j4jJ70
2TG6CDZBUmY7d7aJrmSAlhq/pP64uNKCBqWyB5T+coQH6crmQoXru/bizeWc
6WNN42eeM+uB4YFtOSYpjzaaSvctjtrl9+D3/RiF8VYdqgRX/MqtZmvZVTiA
jhyl4m0MzpbDNrZifVCmXKbcxKj1WuN3u5rja8m31Iwx8WxaVctw/UVYDA3s
V1Pq7HKa8u9xhLbMqX1YAQubR/QXa+/1OMVJX4gG2d46Q9ENTtOg8lIOGKom
55xA/9ntDi6Us9vv5+bx9RPsYBAHoJ/Z9bLUNBtmKy0KFFp6GzMO80uCFnNT
WpwvWZ0aJfsqVdJTfCZNHmashXRDpQoreg4sbLuZVXghU16ppxfyQ3zwGFLf
hhsVhEABFBFxtLxRmO0erUzTJbH/XwibyCXlqlJX1Y9xNA+Kv44qpTMRUeLW
fdwNpNhA9A7EymEBoZRPaio3zStRJiUsVDOK+g4eJKs1U4uLRChY3eP2FIvV
Fx6a1Iz1HHnt1djcVuWJb/wVpIckWq1b5B4zd/2fs4rbFqHWTBKbG63e+YYO
WPrG0jcFyH6sUm3DMSrQEQOGyTeUcNnzpJyi/dr0NOY1G0+ai3ZD0QIw4BHh
3Q1sWC4JCSmta2YbxTFJO7GSKpv9lvGhM0hT6YwBFHWzEoDXw+CFnHS2WA6g
zFKEOudey+IyrEfqLaYDuqm0VxN1C72GD1ASbZ3I5FM3DmR2C2gNgz120PXI
fvQ7jUqQ+X6wYckWG1lV7GgqRic3mj0lqScNI8vMOyllSlRT9SwD0NhooXUB
GsbGLHPeuWdj+SX+Ilz8zmSRy8iecJ4mJImw0Bx1/IKxnUlToy9dO9ccy8sn
t4mODpbOxnsYTtarCqvZzYSCqsksr2Q5RERHSkhAE1hUl11ytlpnu41UJOnP
U0Czui3Ut9/qBiGcaBvyc78D4NASjYNSpgreJNLsNzC2IQkerH+LscVR3M71
HRXE/0PLTc0un0HqNQ/Ttpt0eADv/Uvy0rtxXhrQGoTcT5fAWq5n61NyDFue
6YFAN/Lp4ajpSi4W0CSU3g3JwfGdqnBtyOyE4CxqEk8E6E53RfGpWDr0Xcdn
aCQEVcyu2odMB27DoEcB0cXq6mVsqLOaG0rrstq7GWX1bHjnjxLpSnXHVego
wcnPleMTrw0I6m7x84SfVakXClDfmXmJ43ivEVRP5ugE6M1/cmp4nW7w2vWB
RVHkrR72mNAOiK3FaodGRqTsX6Seseq5y6iKNVvPdmKNXOzsLJnewbA19Svi
Tpmb0n5I334BMfSxvGk2UFGrRn/I+o9PP8h0hTttX4A9qXK2blpiDykL5eVI
XPXJ7NoaxCr/KQ7Uejl9cCPftErCt2YPdkCBrEbSCmkeOoDxZPj8K5JeRFz/
FnYRg7zQJt7smaKVm9F8bp85BFThEgxmPx/votRtP5pcPa1zPnpJb5rJEwb2
ssTq8n7Sll5D5Ouq8q0AKCC1uQ6wXZbwt2rxUiFteYxki+oAEDIsw+11Ufp4
axErX6BNlgPiRrLlUPmFXjiL0QAdxDAdtLzftvrqbI6zGmS2+NDKyMaCywUT
qRhhPEhDXT0bGD3eRpIxv1zG7XLocYbrO0am7llp4q7uT1HxLHI/6YcTyf1Q
aqUmG2GTmSKKKn+TW22CdIvj/cLRY+RHcMXhY5sWoQD0lY9qMSq9zrMjMql9
DCVsFkdRQxuHjrjsWcjOrHW5P/gxE1gORJAvb+lYYFaxcj1A0ibuYTPvSdGF
xNYlvm4ySw+x06Z6iZyFERKVHa04QC7OHFPXfV0AbX+J39CGMzo7007L7Sgq
6I3OCcSkVTow3rw7zebzfXSwOYHEuhS15+G6Ha+lVbiY8/ELPNH6xnr4yzdS
oITICwNdWVw6U4ygV2vIToSc1PNIUdVQsh3lMtsqL3QFvYoZcnuynSAVXLrY
XfYwlbABZiqzgOCh/ZtN0+YCNe0YiBdzJkxpEJs5mGZyqF4p5W73+GnFGouf
ba8tZH9QTQrMQC92pMxEq47uZtK1FXRQAXW2UpojPfKIwj/SjRKiO5huFMTo
1EsLxwEOBijt/Z5oXsWyeEcmTQ5CbSrz9XTzh+TN0RJjWg5h4ROP4j97xA+e
p3WiNOrmNcwT3s+PpgDC0kGlfcBgb9SYYsshLb1GNOszLsLE9Jb2+ayqKpWq
li1ac5z0WCRLHRW7KrehKWU677VHhjFh9ztltn/uFkkd3zLmuEteFp0rpJAw
IcSbLc39/4Qck+KO58zxLpg+5Evp7TYem3LwKHn0h+4y76MerZ5Y57A6Vsui
koACxPh2K7WIJgEO1P57nG/TzaXVu+mSHM02gRb12gBHhfDkrZnyfx7tGzZW
SLrr/fl7+8Yw1zg2z4b+BMYnstWju0P3lre1HnuhrwPHV47aU/+EFj6+341T
+LOyrR5JQERt6zIATg6xTPBf9DH3fgJdhCiMdwIjo4hk+K4XfcTgLz3XmffJ
oBFRCHr6aRIRZ3EpFfb5gFXZhfuu14uochyocFO3LVbgsJ4ooWIjn1DIBjRs
UI1O55zRXG8UJiZjas4cCmCoC8t3QhyfNr6wfkCzxgXylobAbjoGUWY80QQK
kgYJrG3deiYf4qZhCoBU97jZD2ldXR2BsW4WhaAaTyrNd1djhRVDKMVaymjL
UM0J8N0icvrNlxyqLi+5sQ9e/PJIzRXeYZd0d1qeonuHt9iM+FXycaTXVAcW
3euPIyz6KlX06jy2H14ZQgZyhYXU0PkH3/FZPYmgZ6Dio2X7Nb3MamIYso7Z
vG4a6KgwzmNH66I2CwILcXTcaEiq2l1fGOUnRkz3aXEmWQZIyCH4TXdZrqwT
G6LCI68XfjNj3rzSevnIAF3+Lhc95KYqKJTr/Qbm5bK7g2F0nW4gIjmaS9el
D+GSxsUGZmLkavlbZV178ik5jpXRF5mMDy2kacIPXymACFYAweIj7WMGHetN
eH8qhhQxGu+YlfMXKGiypu8JPx7PMBLcEiY1S/ZmaUehwhZz4fwNqc/bfRl7
XvnWblsnj7eij+WUohIP1Zj+fokp3a0reAoMWC+VCKecBU144VR6Liyykpo8
30U6BQ9ujpb7Lc6n0AAv23MvJPkLI4hCsUlOLx4mWVtlbCmyLQ98WIj7a/ZZ
0VC+QrqdKAyU+jkNyd0Hdi1y9aNwEhkE5o9Tdy3e5lxRbb9FsGF780mDzS0F
QZfPJNqZcAh0elhNVk6PobYQDJUnYXOgXqCVqqCR2yYelAP5MlKcscB49dAZ
yszlUkC24dFND+yYj9KOF1WOz/ZJI+v7tJYDAc7HP2e77RSTkWkMikErp+fT
ydxO04kMRl92hjJ6vQoiTCePRyghSTGFKio1Djkj7a0puyvj7nuCturVm6Yh
P6+ahwrafJGFRSdDWhyDxWdbMazqAyKP3glakd6g2kPBSoh27uXyiccQFxLL
SJM7EXbXAYJRgMd8NER/0iVur/z7TqqwINuhGllxgyVkGLROQq+fWIzTfZ2U
PGEXRYLURzM+T7RU+OVDeEEmZyrBm43UptQPwRlgaUhP+ORQMlsT3FrdeLBq
BGCAaTjBarSNz8LzjXU+JyDD8Pz563ITLmjlrPgVLQsYRz+mu1Z8gFtL1gXw
op0cmvdH6GDKBUsJE5hWcuYOAtIbaYr21WWznmRGFCielqKMgmBTwvci0fSn
V5qNRz5Nju2KdtUAbaJPWrqp9P41a7j+XcK4e1A/6kzNt5f/2XS+BWcs+hj5
0132cK5REdnSKb6jDot4X8IboWZQK2Sfagy3Jq4xHuwn17dOcMA3Ev9ckxfP
8hs9V8IyticVS/XXztgqBKqjRqzzn1SR9wAgpJKYMmYeem1Zs13nxUR3B+MN
52/+AYYFuBeBQYW5chRIN9QhGTp0nIjs6PJpYqlYKxTXfUfLYAoLLpHJM3Le
KOhTgOrRg2gj0aJj76t3Px683CmKcOYENL2qbJO1gakUU3bW3XNHZqoV7EGC
OX6jbcdd/LM8Y+BaOUMp03ZpGdZmCHcVG+BWqROgjLq0duNikAGftQ08VoT7
hbzTzGCoeGeuXSB7dAGCRO0z+y0NzkQ5uhVkqEPPNi/ZVjWFhqm8SXOX1EcE
i9NoxbPphG6wt3dRvI3btKOLz84QLX1yJdzzoTQN9vPEMPCLvEB9suy1VbQ4
mEMaAMDLIlI6S+cDk/hskk34uLUiYIKlVGJF/nXfqQg+3FJ9H8Na0jPu4JMK
bnfvfIz3s9trXr5xN7cb3LAnW2kJX48QYq/3AIhq6bzrNnjXswPAplEWPRrt
bzoM+cRnwJivyHI/ewHmpSmofy0ONPtw6FkwrrqKW3iQp+Apnriz3VSTs5Cx
jWlgDe6hUXT1g5Uqtt2r5uLUaeqkrInTId77bbqH/orEIvdC8CsdmGRKc/xH
cOPTlSIGDd/kpLmGpLSKKlZI01YNnt1DUSk0/Sg7DHh46Iqlg0mPvjWRm9ii
ld4syKUMaJjuqkyzsYs22YdY1PcTWpdHvyNaEdyRmyHhd4RM5+YE6V+JNfFv
jmQFSSTQOaMKocjLw5o0h+drzET6qCLcvKzEAYAnFSEo25cgF7m/t81ecD1Z
Z5HrPw7WMGMm6ss+SdpFK9U8C9cbM6J1COx1UexW/5GmnDYSSARxc49qCWpr
UB2nEzG0PwD0UdWKMI6jnHO5Za65ytwdWUTJnrj5Jyrl2HHjoTkxBtzS5J8I
cscyeJ1OW5MztMA7TRkYc7dNg9XRUmJ2LYQ7ka8YtfNtp/ynkc3xTayctHdN
cGX2Pmt34UmH1elec4Fyjrp8DxkhikJ8R5Szs6McIxFBBxbIIfMJXIitqEuJ
HvSIYYiZ4YVaaZ3XhOLnJ4VPLqCdRxbDdV9t0C3etbhJrrMWl1EjA3DU4K51
/WVZPyvtiyEnSn4caYwniYw9CZYJeX7FcSw4S/8YcRsIC6pDvNMFfqPfn1jL
AqNEuKP2igqKQNmEbHD4TtmrqT1aqePValSpQYxQ8XcxI9gcsKomMpffMALK
9HLrkXr5cfuNxDn6YK7T90D3Y5IYm4EAQBuhIKuLp4mOmF9dOSGpYKtV3Qwi
WRj3Vg/V78b882RLCzel1SqiyYpOwhnIy+2Np0K4rI0C0CvB3fL1Ny2HlGWu
Rc1Tgd6YuDB1abO2wtZ1rMF4yt2xNVvwRmdJTSfXscMc7n5XQeoF/32Aoveg
gziAOL/V43acQ00JatG7UOxZkCLUHF6JyUamhfAKyPj1qaU4coRjLyvkg0uJ
bdLHhIQQ6oliBbF/N3110mLLGJeUtxUIXo6ElkgwfLK7hueoqkFu5r5WrIaj
06zZ09PAQhohiN0sae5HhdM3sDRHKZOyHU5GKbrHb22uwKnq1sr2CTiyQhro
ycSS6R/9FNst+WAg9MXesJ0FKy5d1oXtE4AbfNXt3Jod/Httk6Bnu2xkkm4c
G3ACLo7yvKt5OaZ3Uf4hSd7tsLQdM9DVgE6TusC7G/0Mu2Cd5tPpgkJ67TBw
IX0CDYoqpJae/l3TSMTgB0D2/wPeQw/NtY6FQ8bq4IfieXsGaIEh1h+nY/Ka
HRyHLUobtS1jIzcsmh5L44vuCvxrZMqvpreyLjU06h5QO4v/6irLv/wN0tmX
4a0ZxINCuYXhSvrgYW+h+O8hBEos1kVIXqLrXpamMcBla4xPlNLgJhG4sKfr
A6EJ2U/+T/ozdKkok+kxN73v2Lgy3d+HsoFeKyisixnA1gFSgaHgWt5jjAMZ
bp1wWUbWfySbW2a/HB0QrA3hSY6O7yH/QDvx3mTG4BbywGCiYWvVLIHMM0aF
vALgaaQRfebt3FjfXY3+75Vkpgifa1jYZM7p/AxI6LodoHrGnojDoFizPO8f
yEccRfPoi9PdkI/JbbTv8eVtDVkrUgASgGAXGOOxnP9O6gpxotNufkvpnBCi
CbRgIwHddu5/bjtSBoQlONlHIpBaYxeJxAH2EWaMg24BJ+YllYBdXvTl2Jzi
CECmdKtj59gvWOuROThDYgbvpB4z8KUhn8/UY4vgmBZODBc66MII8/0liNEI
prmzrx8yEBG1/pyZ6Qm0gUphPqJ4SFy73sMW31HvRQEdtJm7L7X1wrOlF0YN
dHP8isiNltxPyZSegT/y4c0jm70FdYrgq+VFC//UXDjifc1ddNAQZ9EIEfCg
AEVydph0uMxBn1K0feztFrQo4roPtwUCR9/gSyg6oe7b6eABDG+J4ArpkNiU
tk5kJDzfHJbKvkoTpj0WyWLzwxQUARmrTj4OOZTxtqf4MOkbQ9UzYyAepD1q
adN1fdE7CtECe/tXSwgNUqA8OaRFaWkEI/vnmPOn1g9m7eNC7eUIJrsHqzSz
LIKNqXCj9lVvLtpPLbk2VjsOaA062a0wnWNScik59TATfNxbG3Pv680yuGdq
t3MHkNvmvSfK4AOFcBGA+vSXoS05pCiyr4ymjHdsKbHQ39gU4SI9wCgXvhhV
h+FZgdgFwmRtdzx06YhGjyvxSJNHFzy+fyIl/MqOIg0I1kBYdEEwWIFVTkUP
MeyP8ePd23E3PUHYbmScBsicc8jP/cmqhhbJcbzVSrKKSs4lCfQUP0F8ec60
0bsQgQtKNImcJNFEiDmOZHWGrR59ex1lbKMA7GD4P6V+TWYyzn7ejEsAQ8jZ
nc65CZFyxtRIDPEn3Pv1nbYPmOKAqWSMgu23Di58ikyYY9wrXCQflQ9SBL/m
YkoD6iXSiR8vhWwf9GJfof3LjTBvJ2dnVQWA5wkKBqxdOlm4JhifHNFlXEJi
EDQrGzHYYKxDtSzfdfTD4y0sNFM5EEdYvwCnzr9O3J3U/8DJxnHBe6gL4b77
DX8TlyAqBPKCNSp/+MvS1M4eRRK+Qr9tzR3qUEwcfePsVPFUP/1gkf1F59kG
7tO8amt3ntakCRUa8THZoMcTeKdmZqbl/51MWJzspsJ7BHML6nyMhlFpEov9
gyfI1pmLuHbxaqqvE0Kci+ILUBnfoWT7o/0gDOcerh1pBiryaEGHjmhu12pl
FAz9NNvzpGynjpL1IKSRxepnAgZUdkLw2MU08NcjbwV0gfP9rPW2QMIRzhk6
pkSZ4nXXUIF6VVVNSnp34Yqd/mBxTEs42PEvct63nC1OPrY7fqWfwJQCiv+p
J4XoDi32UFCYbUfqYhDklSDwQEi6TuxoNUQwnU4XRWkF31OpIufaeiqj6xMF
lEb8jqI8Xq4ck7xi2o6wL2Z40HNrP77Fs5Kc8T9aWn4K8H15Uf1qm59ElhLN
SY9447b/Wdw0LAgXQyEd5cAMsY4waT2aEaOoquAAYbtTzDaTwQ5KcmwDfp3+
BKZFfh8Kw/bW1cSVV2wNGRUG+FVBWwrtarj8ntWV+rbdzbPWPF/WiHpaXREu
8KbAP1l3ZSULdcOgVnZ6LqJpJUa7SwKsHvhKfssPD6vrheCjbvrM+6iwVZDa
Jxhy3NAHdl5uhyQAh+Ftg0RympqrhhejtEsRZOivJyFg63tS9Z6ihrBdjfeh
Un6nMlNTe9UGJmRUt/tKOZXXuvRoKVkzBm/9YdvWJSaO+1YceKmSpfgVQDmR
KmLYvoiU3M3bFs9yNJqBGCBaWNkxur6DO+kDA7RLR0ElAfSDF2qydsXnEYSX
AabTWYK5476J+DRZAnRW9EmYCs+Uho+2ehzb77ez+Q4Y4/YMdCqs0IKh3Q2G
SRxBz9mA2cGgGb3l2Keh3xa9IU+3VqFIzLx+bXRXODgnmYfSdA4IPzF4G/SJ
tHgMrw3IhKcVAHISqjEh27NboS7qXx6lMLwXmAdgCqAzMXIXtungG3ttJiCh
BA49+wbbBajTrlahTStQNyzBqhjKLJgfqiDAV6UogVFsKrHyyvrTv8gHGSxi
3JibzzpEQ0dVtutESbiarLua2/ei+uBOeFq0qemOySYGF3FThpbQ8KYPOJhe
G/l0TnHEDSgjpBQTS5SCjU56B4UD/Bbkk8GDdkIsquX+04+3EzwTxRn/Pv6Q
i+jZgmOu8cEKoZLMycZZRxrjqnaiZgCHViiWqdANdJHl9hK/jLDQLI5ME86w
00aH0MyGxd5PcPKSH1EnN4zKPj53i3QOaRTIBul3pADOIDg5NmhdzsA56MSv
fc07bEuxNxQ6Rca/YTqKHKZzuXPJi/9p6Nar3G5D7rXyoCPsMMVsEBMdXAqM
skGgB3VtPvluX/jwvBFm21nxXouR5SETENGDfiavIm/o6h+3YJR4ckubg8V0
yh3SC8Dtk/Y2Mq48K/Fx/DVRNXIrXtSkRFZ+jhWCQu4TRqISKf//C8phahP1
htMM9OSEapcsp/BrqwQBCUdooXrgvMCZcIPy4+5bqHr++p6OrmCV2PDaFuXX
KrarlBx9u3dxDxSzZRL6nqhzGIILiQwbCM7K/ZIDW6auGpvWdXOo3WdyeLJX
BXLciqAO/T9N69t4KXZjO4BeW9b4b2XGMOrUsUhAyyh/3OM2UabDsNOJYFVb
Sz4/YUHT0Y1Js8DKPYdgmaPDduvFEHY7U8cxB/yUhyZqKQYAcBirfaYA9VbW
j/DjKMc7NpFuvGkQ3upUAq/jaBm9SujTN4NFlJPHjuq+c/Ra9raXHTZEIC8s
TKNOvYRt/kArhU0v19+LY6dtbeKfW8NWxPF225R0JwCPtteo1n8TWFP1wrlT
YjMvgnTkCgeVzLvNYxLM6FaylQg64XL/z0z5Jf68040p35Vd4HliMJqScASg
bQ0sWWe8P9Tm/PmtRIv2lhzKeP6H0AvzMh68lXx3fmjG2h4OppBBeDoOB4PR
t0/LATLLSd5L9Ps2w34xj7fqS40Qq6AazU1CkOLbXk15NdNq5td6QQFxE3Bz
Afs+0cp6JZrBLz0A6kOn5II8a12j5I4ApX1c3EcLQrPs+RJTa0WIVIt+GeAZ
AXMkTjKx5jLVdnEke3vhI8uj8uaX8zAOuckniOQBzGSyPP+VJTN191UjxZ8i
EYbnAxxrWQHtu02RL8KYAiOPQpxK1+OWsy5KdhgkN9F2S3n0weXscz6UQqZ1
HMSV5sdMrCujNuBnSVnlrRuTcva8LTLws2afjcDOilSDgV2uEpF4rqFXT602
NIXOGbXxbFXeNydDqjZLoF0XdzVugXS0/Zq97iXCPoyKRcAkEkJ80q6IdvUT
5INZ5wSGupROD6YOFZoi20hIv3w/GWhpGFlF9IaExnWQUlT/pwqtql3R9huq
TpqiesN3wOs4XoLwWZMmFQrlGUOyIHL4Nr20VrIW21daEnZRvCoDbkmYf/54
z6nJZCydyXgJ5MMZ+P5thz5nqb5e+f/MA5vTx4TsadmrawTU1zmf4BmxciZw
swIPCZtJaScc64Vq5wP+Ig7ck1BunpMpsoXpypf6bRydrREldti8EruRM6x+
R1MugpJvyjruvKHwL1DoFkKfdNa1Kpiew3OnPKPwPEtvjQwBdl17JWPfLV0e
mFMgxsyhsurPnOJvX3NWIbwUwzEK6zFXxt2bDlbCNTrqPhKq8lwYLUyAJkbS
ZA5lq0/J0vE9guahOiRzIld+8yd/1exdYAKBOxx66abEwQ3Y2BOOI+7ubMOY
5xkBZZyKuopi69Rgf4PyGmmbLvGPxdDGQXNfF28maaF71EYEE6pfuC1Y2zT6
b3f6k65ZkzzNfnK7bBSV45gOz+krRNhN9emjiV23iAjFP5CLZmtpHKwDUnuY
yCKve6cCqhGSkEHI581l8cBia5epUPKPJL9X+tSvq0HLJOAlGinab82sGmJu
1XIEMwk6o8MUQihj3hpa3sntq0pJXoADagWl0XXiHPZdUvlQwACNVvOMcoLX
QDd6aAzBZeIdpytT7Ux0D3AEEhf5AmZJdshpfbLZGG8LaepfvDtsx9L0ieGI
8HJxEVW8puGk0WHzFFCFpwZl4QFDUDuvfLhGhYEHPcPmDDmJNw4uQFxYm7tw
ZFFxqlN8BPCP9KifZYZ0uzgHv1WBJ5xrmrHRo5bEogvDZ1QLkqCeNZ786soY
aVthP/HR3U8qOzMoRiKL0jfVZ3P2MzOCBDKxVLydylkwOxE4KVj/zE7kRsCQ
/UG4meTNF7EVaFcrIicJ1jdSl9fMkOkGclZiPdpLfuTjSaIscrXd9NXuYcys
/xa+DLwyifWeHhuCP1VjHZKWq10nfOhRrss+qX2coEdwcUmMDvsyqh9V9q/J
vbE/BxJBK0MDi61JlLg2EqmCdcDey7MSE9VDyzdKSTwHQjAbjFHlBMWW0FP9
UDA1zMQ1efjqs0uZHdsjyQynt6jI+lsMfT5mDU4O7TcrHtdZfJaOG2y7KqWO
jAj/HvOH1BDFATvLJs4xbG3bxMpR8tWUkWe0KzhDZBHJdyhw5/mJ2JqJBRs2
aoeXrEISNqTV7T+nHobUq0LPtxFeptvirqS0ZhDEZEkV10hqoBfVvG658iWS
FBDJvm32bjo6ShYQ6fT6cuxaknSbyuHhXNfCGCYHJcR20vDG/HnK/Ss28tCZ
gxjmvLTJtGubb8e39bjpd8OOBkrVS19T3hnnrqZydfuLgn9dhCUTkkzMZALq
07jNrkLn8K605SGwDhfQCYeNqyO8uY/bbGb82a6GlSgA1n9Ldop1tmBEFoPC
TOJPnQDuDCDFDR/uX0nZH3KO9HRilLamff4RiS77ZezYFldOgvnj9cXcMlF6
AdND18BCHa2hzYSYraTsZ4RFCInBqIh80sUAIb8Af0hpFq7Of9ykgpWfSGeM
PjmvWkQmvL9DDOa6sDFAvUQ36NP3gd5ZLuABfZKHPnOtKOGvPaBSo76qO10S
qx0tOP/OzOcmGg2U/K2qJvGf2mDsa9yfGHv03qAIAsFFIleK79+w0/tCHrOG
nDsrEoqnU3rdLXv1N6JO5qs4CrP6BaivozIfaD4SlqC36uFiDmg5EA2l0vFv
7scL6GVNAyXGPlmqHXtN2P0S8iaEq508ToNV15plW22Jg9z4t4xn7bM0hMGU
Ug29h84I4QWju+A5MCpLCVpBW4fhUAr6WUL/JValnT9TCSpJB+U+vxIoisQf
TU93MJIgaj/EjwSZRRwetYFfxCpVR0ackJCm18dmUZ2AGrPymZcydJzqbixC
nAgWnWqLYz5RVGmr+5yAbwzxqTzNg8zeMcp2FKWUDbc7rNeQGUb2NnMFvTXN
JwpTyQ9dfzHYueLsufi8Tt+RB1KRThUy1eFChBZSpVjNoDJ9O7iucEUaC6Vx
fw1q3AEyf/G/o4dRm1KmsyIG2NQyGXp9WSaSuNf6P7A+Mm2otKWUgBV3dy6H
8IAqJS4U4mT1RAb4h/EoU0IRMZokPM9u1L3e/FdzRp6oLcjLPmKo+gHKNGMK
f3IOi4KNYxLU0En6O2v50nWMvw/OczBQTdSIKOvBTGsBHBQyO3k9TsSl+DUU
1bChHsT6H8qwgA+Kaal6euDHv9SxrDjPirjmysD79sm07BfaFLyugg92QQ+5
INNEoOpnCfCwy4l89YR0m1sm8Gug7y9pLbcP0KlrnhGrU5zJSwusY7L1T9ut
SmWZAf9iUiDX1R2xm9SWVrLWihBQ6SC4rRPIcgx2pVy7owQ9n3IZJlXZmoCA
bsTyVmpCN2HHCvozUhZCUBDDTJ2umcFLE5wOlzPul+q5U2vJYa901QVh4x7F
a9LQbrnHDmE4XhmP+mt0m7/xDr6qh/JF3aDOARKqCxntH063qsic3r7Ff+dt
0QIhJ+Z36nHTmeNDdrsr7XWm/B7eCigf+w5BAvsobmVGMUI6ylbjA6AGyX1S
Xg3WGj5XXSBeSjq8i5J6lX3ubA5t9xnuOE95X7f5O0TbrbXMVGhpasxmBSmw
ttLo92ozxtovjGvk36Ia4ZGXKylHhI8suJ0GF4kR7rz6VQkX5NdcuT+ZS5tf
gbWkezEaWq1D0WcP63ttR5gnGbGI81hrBsxj7lOCh819YMnPR9tzv8F3sVGW
xdpGZBvqJDkTAkNErS4qwko+nUleW6RZXKUJtxdudhWESLD64ozOcCoeUdHu
4BIGqjB2zj+/iXoDw66yGbTqIzKwvFcf6pJJDnl6FLPRnw4H1s3/hvcwdpMo
LlOI/F6gcqZ9St0o6zFiGb94EAJQy6Z5jjh8baOuZN0qAETcSxvOfNcj6s5b
7FlUoUNsFUgjTn9ZhzFK6AVkLWGs430Dkap1e9YMaUeP4Idfrg7QftkuMt5V
ALENDHCCaAv+/UTXI9hTZ8SweCh0qK4v6R1sW3I+6MChfChfnMLeVG1Qfnk3
5OoCdJVchBA3z6SKrVdETjXhNpBsNUXVDwaN5SZd8YHhqKtnhqHjATb4UwZE
09OGJc8GWmIoWEO1rROR50OgVZdIOFUM1BtsPqmbHNuzDTJTHtiz/3mVUC/W
r/1SXPtP68/yy+eG3bYvav8B35HCGVzu/7sVKQDcZlFlvWu3rRNJ8Md4ZxYk
7CeRyx7ThvBTnzRnEtssIFRCZXgZJyjEMPbvSw1rvwpGz81QsIVWgSp98epf
aFg6OLfDpGrQFnKa1S5BJH5zAxJakjdZoPidO0MQaUa5Do0Z0NOK3ha04gZi
sfY3vKz6pq8Rp4U/zbUrahZ61nthAnezEaySdZtx5JMV7B+mf+/EbSJ6mRGW
dSGQp2LINmEZauFnrOQ7ydewDVk0P6EzrWSJDweSik63RS4grhsup5MlnE2x
oMciplSzYpvvo9F8ScCXRSz7yZjmSs4vaWwca3aWcz7k/D1IPdS+o5SD4Vo2
vZT3FibBKLjenN94NbIoY58CC2v/C1cZ34qd/apJdKqISwGKmDKKjtbJE+26
2ZfoYwKry3KRCrP+Bx5YcrmUt0FgghQjJ/n1H1rD0SD7ExDZHCamJDlENB+0
vOr8xTjqHJ4vF1rtrTJu4gUOkSMPDhaY95cnDWqCIZAeNqi7jnGe10D4RHND
YK67ShR0ihYyo36W8vIdta4xZtABEh3Az+yChW01C9iZ5W9E4wkBwkVFtBc0
mpt+NzTmIr2c8ttTMSRuHCsRXbNh6PVXRoP3K7RLV3N6dk27Y+WEY8XVL1bf
Y22iMi91TYBMS8n3K2c5E5Bdxpu48m7W783/Y7GM+PBlsERMLbcBaCYnRXu4
VtSi3xGRxMJUI5FhLFFY+kIMOlC4Q+hkXW3naB1UciFPNKohIoW+EefTPIMX
z/UuyX18zgxnao1rFKVKiK3gkirm+x5TMELogfUR0xK3kA9oSuOKUd687hez
ina+LD1H/VP0FkaKukwky5cBtUoHwvcVK6vptfKOaVBkiDSrVWzlLk8mJM3G
M7wzQo+ylzXCo+y2xelw2fm77FFZjjkIm5aGAd0uB7r7gNi8FyYMgpbTcTYG
OWjm8UbJRN5juOoS82EjGVZ2XafORTeQfyPHhAnFhNOksVVCLlYg/uMWCWCE
sRRhzTE0AuXfNo5wSVwyZcCSGpeguVgVRsK/0ilCKvyKwrfllUHxJZ2grP5x
C1QSQrXedbkrC96nx1c0meKLgzKsaHk1mkKVlUMj+NlPh8JcLZluA54dB+sO
MW3CL15EBzu4C+3yD9kJ0tf0iKtxz4rJND+CFoiU7JaFh6wWqdsIQh70TxHS
WN1gasUgAbdBrzxdrro7MbzvEP8jLQUmUEAXeJ5tSWnhjYGxNAJpA3IbMBz5
3C93hXsI5SvjZ1jwUQo9LcCO7MN33SpcXWAFjBLSY4Fct4SeDVsXJ5nRUyxM
x8BKDO4ICidSlNKrJno5EObXDcJhtwMGTsdXSL8SCaOqRDbNJy9RBGSy+a/0
ycX4cw4YpdcAMhlWW87Xbzsv+3Eqm0BRF1d1Eeb7/8Pk12h+8+6DDNIOteXI
ihfuXt/MCfXp9db/TQFuqyAZ2Zpbn5QIyq99qrtLhZqev830YbM4hphalM1C
6gvh2uRwcnPxI/pmlP1hjT2aVsbAIGvjcnnQdpYputfM//gUr6sq65a/vM2/
WmsApa/3EypQho3O7GJMXNZdlUnqGz5mEKcw8xfqrdsg8hDBGxyZqgATQjJx
clYu2Y/NkXJOMpW+dA6JmBgzep7l6dgcuIsf7NXXcM7ME3lYBeF2labFeH9N
eY+N/Tw9KECIpjzchQmpSxfr8ngJg/DMyUk038mqIEolwvKR5WFhvXSLkakD
5RQ9eZyRU22uxO2fKYwUAJLREMMxQzVn+unDvHapiKJ3INOV8PCzzujSSqIe
W8jWoooq0nPlQGaEAbdr8oPT+NGNzNyM8PfuqyvVioTfWdMDV/nqYTR7shBu
gYEdHgqoDkf2+F071jNAK9/rijgzW00I8qLqhxN+IDAG+AYtVmn/kzrCGhgo
0HF7TK5jSvMq0uasKKY88zd1MPT2VJqHw7sZr5uB9dX+6hTvjJx7nvdRMtAa
KCQjOc4sewSF2xK7OP54dgpPHHDqvx1ki+wYLLGVbTTA5beae6HnQCJ4HCcJ
032uOhdD8bHKKvtaGhaj31RsVriY1mg+V8sefkXiT8dBjf8HAwmlV2nxbHmq
SN512EkWhDm4VMYD2yyHNmmRaKcO7qrQQCnx2lYi4cslYMR567oOVlTUWFIq
gEerEHSrD4Guf30JRGH9FHhSNcf1jV5D+GI+eA1tsPyXTeYWRRJizCZZVzKh
8tf0HWWWyayNH/OIfORvO8bSVFkDcgqKeN9meaG9cjNGgYOZLfaf

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1I/On3jslA9pqSLUSDie+mX1GQxJ6K/5cg7i9WzPmEM5HFi8a6TMwWTf9qfjHASgC5HeKPNPzPhemRzbxeD1JqlDe9DjfYhNXnQLfZZ42KhU5ORfFkIFnkIRJOruZdstwxH/ncVZly7+PtelYUb+SgE3rZLd9Ur1vThv9fazhfLEIOTYt1Nw3vkrHH9cKfzwlWQ5qa34AZQK7AdjvC+Y7tZoRUCI08TO3LLSo0qOvpOn5fabx7/ZC8q8NvW/kzKS8nkQBvPY9D6GOo3tESwVViC3aBss4sFPhAM5TI2Ye6dYozuaKGPaLSErf2T/F5HmLdw2G1nT6ZwbYZCwE0+Cql3mxwBd296CQg0ehHvF0dQdJDCcqE76xrhXduE77YthjqZaDHQ7Fj8+XoQmEMIruP5hGsc1FDe5LQ1T+7nEcsym8Q/EVwEuUMV92F7TX7votSRjdzdahcdwueQ1ccXCVwY4295oBgehFz+ZzAFso3rzdkfhRKzwZtB6Ao2PWRnMdWL1XihiJGsODZJX092VkKnrSEGOTDCwjL+6PC4kFWdjzN7zQytwhqa0vQScXPzqKU+PPHVPhy4Id5liaOQsURCWG2QAJD/m4SbGLSRY7O90KdYK9I5oYEOlmmMSfZogVWsYxGLy8S9Kj9SPGkG8dDnuTfMG+Hi4OxEPZdLjn9ea7dnfRn/a8duGm4pQPhwEYelozXzbqQqoD/Ai5OLV2kTqMh0TMXXyppfbnQoEbdPVlxBnWHID4XL8UlFqYEghcDqMzoDEeAspe1WPcw49kxw"
`endif