// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vpEWzQn77A1KwrvGPfFRRV2cIKHtqg1J6H3bgF5UitOZMux8qJsi9HW8Il26
ZBwYnH/DgUt3Pq8pJz5f7xnqn0LoOrdMxtWhQpezRqICmgM1e8wrOHCC3jrl
CR7jukl6IchGbhukqyZnWoLdm1i9P9SjTJoKmEKbdfbpUrIEYs1xZTl6I8qm
8A8lHly+HvZD2evBXR+DgPyRHOPCxSm+pgoCLEhAwAiJ5eT9iwvGrKNvBHV5
wUbFv12OOgRppmFL7aKxH5W1dzi8JymvgsT3ZAbVYObRpVr1uJJYWlpOBVcp
+M9lmdwnHcWU2iud7O1xzZvTVYtViCgXrPLYT9JPEw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CwVpc6jTV5RoyLHO8FVxJQgmZf++dS3oEcXnHRSfVlHGc/IqdEujVk0bORBm
jbqXzE3WT8De6yxmTBpqBkpPy2nVTCNN7x+0mHTzIGmkzYZWAqtslDeZ2Q05
hMGYoRcpY7H0aeOWOhbzp1Z3FtbTBeMOdxM0Kxdknh8eZUK/Ew1DItV07+RJ
eATPzsTr/zYGzQbAS7mTgr4jZvPY4u64q3Ar7ydSoGA+2VFUBFx3HzTgWTcK
BwtEbZkWLSV16q0VHk9QyNIiswxRFxzL7psDX4rPkPHpipsY9CPFEAatSDNc
I/geqyNu/AhYnfuiqoSm+zLRu1A38XTSzagQH32/5A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S8WBYLuwf+G8Bchrl3zEJNk63rpw9FxkihOiS2OcJ38XDW2XIf9ox7gW0ilm
N9v2WJB3L6PUntUs6pwQTIsi0dbUGVjFhoL7r0OrnSIcbxyVUtToV+bvqk/d
disdYnAaIWdeJfolt1zvC1f4ekxFVZ7WC8dvarShlVw+fchfl/TdKlIBq7/G
Xhi53weHtPwCCs7NDxwKXwGZe/a5oBeHCTb4yoHoQ19djd/0LZtLWG7K3XS4
GoYG5OtXJJGPlw7Tr3xFQyB4zJooV4Hb2Iu7cHSMSR/EN0T7J3rz/sYoUaO1
IqLxtguuUgNSVIV8yJxClytXsudRKWNNG17ydg4zmg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JXKbW3dKjJ8xjXlfymFmskpUU3iWGpVRxDe+WROGo3aONKle666/HM0A5/r3
ZyxqvojEepyrbCem2TL2AlwrZH148KY/ZBSP39YtKuDz1xLKUUbpFklxTS8j
fiXxUz6D3suYIOX64hJ7kdUVqXVUTf36IKfgIkcq8WTjKQnVNETd46rJXTwL
6rwDj0/ZKYIWhFZu3QYINoEqzFMKoSSz6b6DIZr5irEpql9BzgfQdRAPUaac
NeYNaMsk7bydqD1NwsojKJKO61KpdnFHLVC+98uBQjMj7CbELnSk9SwvgtEo
RDARxazTNW7+jl0tamiIDiem2oHxilxbyj8yeDk4Vg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ea9w8tjNshfC4eXweXMlbssse/plBAk5UoZbJaSom56DxbE7Ut+hSDtAIhXV
25CYLZJ31GeYaraF3BBuhQJaVBl905aWzcsim1IGN2wW1ssApOO03qH0j8Mv
8csLtqvbBwAammOvIz7QNo9dIWyfBSyvE7zQWrHjmtmgUK2TeyA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aGxrbTIFUZA5Cqkly/+iE/fuky89hWVDaUW0ylj2pFbv0fiZi3uaYBlyhU+g
m8iseOc6uv3CPhzXaVS42b5SqLjhjF1HqZbGihljmgiOrKxRF/PTZ/dOxivq
bbsNKEr+ref4PP8p6jq/QsfgAnrHXnxJAAz1MOnMsSwnLO/0QMB0lRgI5A3/
oD2VN/i5BDD+YVfaJ5Xayt3usAClMHN4qLuxo6lAEAHNPAIscBQ9N97iHcf2
F1JW0OoAfHkQrDYAUzqj0UXGxVlrnhhO/t/JqfBkPDFMTuqNWrLsZNL/YdRw
OwM58XCQmd5UKaX+Oj71bsqTyCdl8tWkfesjUC0Le7ZGrGrQve+ulGLodV1z
DSXvaKUP5ZGWRr/JsnA8RZfy0yLQQzHLmur2BdiTUuPL+cGSTpGg1mufnmpt
LN0ozU9qIu28kaTJzXFyQtJbVFpjV8E7L/hNE1VgKyycNzPy9z0Ms22ZuXZI
03yVEKnfCRAs8OdriRBeblo85aug/UF+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NFWWlyN0O2hnqGvb88xAHRreg2MusUtSG8JAmpSJxjns76dZ1WzoaBOjS0an
ybUoqGtDXp4swN/5mAoSIKHLwrwHLBfS/bHW8GZmuewWmAngpPjh9XGOjh5G
FFAaFEtcK16SC1q4d9CCGT2fLoTnEINKElQ+HPJz/EwTVsvUpSg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KMy6K3OgRPTyrw6BNEt5LXN1D1ujt6UxbcA7TdnR63yyIU08OvuCdDM0B77h
gZ4621rSWPgz5gP18wGjEPmMYuk7KJmZFceOFpebZHaFDZoxCMhc50hxdhF5
sbPK42F3F7qGXTJxBLhsD2a4u3z+ZGRu7euz9KiiJEePJx5TROc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 38784)
`pragma protect data_block
T7YrXE7TM7/dqzp3mGh+wiXqbYiwapZZEQeZ0iypeJIkZCiVWPYZCJHm14gQ
dROY0yna4SyvBD9WNMI49dXVQNLJpV6KYCyofWZGyGiBMQSXWUNZSQeoakhT
TlbexPj12GLpkXiLHfuPDvdnr7L6wi7NV1ZMRgOUcbdKu29bTqSY/4IKxuRz
NLMOs2S2fsEU9dmiSp4aD0UW2gFpomP6l7dylzB8ryf9riT0/zkgnX+aESwY
dD16xoHB7cO8brKF80t8M5V6Yw9cdBSawADGcfDpsE/1BS1Nu0ue+Jlp/IZx
/45edSqbDjzdJwqd0A6mf9puUgODfZAChUc8TnEdt7Gtg2lBlqllWYL+KZ0Q
fIV+W3v1i41Aqh/caYjo2nHAxI3lQhvxvFHg07XqcvbomfBGy5+i60ddg6ov
f3Yaq3Hqy29kU+T/qjw+mGdlgw9sPpSwJEaxrLPwrwPxQwNa5Nx4sZMnM19a
EhyVZL8e439+fbOv/flZID8V/HsYjorO9PQgGon17FHix/QbnPNEiiv01nYM
twbpBtgIyCCxUndW2XFz4w/ZXTEk3QCtre+Av6f9Dp3b8kwO7QTD8YRwRapi
h6fWrb4o2uNZU7+EuC1f7ouz+bmmgNSvEHQyuEsdU9YycVnegZQ8zL9Quzeb
KVZ7oedxx2KTte7kHz26+vBmr6VT07sXyAJRNMafGlAa2MSiZudfMyq2J3Of
B0r9M7UxNxSSwK9IorFozxWtq68J0YQxuYAdjVWLDvIzMZPRNa+pVOLXDSSs
0BVhNoXp4TXceQda1UG5mLD/p71w99lipdqRsQtriYX6pEAVKxW1HKBuv1PD
5TC69Teno/uQgdVhMRVhzu6tBlQoi30+++nPdHJv5B2LehQuSsCAlMVA584/
vcvnv5bQl2enZU0FbWS3cAA6v1Y2ZYMGk/AOVZVVkPHIq6DUNCCnyTqZinQ0
9H+5KQmYdLZ+HboLgVRAr9rLbjGXRB3WUtuZl2xZA5jM0/4NctVE3GwpYh2x
N5mGVgZLVG7mmEWqoc2VQhy99j3h1Gl1Ni79vwO9x5uJGNeix4KtjLMcEqOQ
vf4Vh7L240u3BM6kO709669llG1fj+84Vh6HItj2Joh/yoABqCoO4IQ4SBTA
9hZLfHitzlYFzTN5okCNkTY3TTg2mMLFyzMBdkqWXaaojjkfYkyn/l5fJrqL
NVY9ntwtOMVu0VgBgkJLXSf+hOde4zK6DzZoVxd1mx+ESjJHjMTgvjfsHmCs
4JZf7JciXTzyy18CWnvV32ALXuUTdOWKbuhFeIq3m5dCo3X3GVlKY9Q5lGsw
TcvVHLsgBXQ/u+3I47E573c9TIvYnuQ0LJpL/oXxmIqAP92xXbw8KRYb601U
9nfhxV+YZ2irB67EJhNTYv1851QjnqaCmUUsebPahPJQ67PBMvAbVZmThq6G
NU+xYJvVYOnP2j3DgEsm1k3jloVmivNqfWy+6jK9asqw/ndmmyq17u9vGBtm
RPmJs8kyI+s7HCLLHl4U9RyyEVCd8p/+igleu4q8YkQVcu30FlfeI6MBx9VC
zA+jJdFz/cVnTTt8TaqrnW4V/X3KXIdOkxMmbKHvoMpFJdtFPF/650E+uMob
BkEOdNpBNryvYdmn6hBum33pMJS+aDFiqcYnCqSWcQPr0PHa04P0n2PjTYQr
pRNyH7w3uphuPLfOywM2z39JFteF1YQwK6ubltTj0J02VpRQyZznng+QQrst
I5NXhjdcFEohbS6yWoPafP/zNQGJVOfAr+EKY0Tm2AcsQZtPDA7/bxx7vc5w
dnYor+ym83acKpKe0JU0Qr+ptiLgK+eye6bZOHjeqV3uKEIOEmXc0xwO31RM
CIhqgJLQHrap1+/jdXgwu0PlYj9AsN/rziojvoAg865XEQveFLMVXNhhFKAF
JJPK0zAUnBOt3+6uCnw4knXIm4o7EJmdx4Mjs88hru9WNtMXOz8o5EdHsGqZ
XGQhWZQ9t0Zo+L9QzA5N+/r6LBpO/Y7mkzOb5G+9b77F7I0Z/sPhgVQVHcyv
oLesvsWtsDxjtTl3Zjjbu8zFaDBqQ9sp7UywPQeZvHWxe27P4ZIQ9A5fs9g7
Xsd0C0a5uvlDxX4j/an2qlkj0rujJ4hOU3Bfc/bBxgS5p1zliIOOvEZCjl+a
qD4EaFPuzwmRwC9O/tY5jPfKQSJ46s5ez243gXPXz5nBtdTmicqF/4aPaumD
olW/zx2Ydbw5NmCxcvR3CbmTAJWQstjjFaCqWEv8RFTlZPhdldgISP3WGrba
BhYEWCMw4Or604h/r043v/pulS/lIGYOWrHAkiPvSFUD+ywJY8dJxELBt8xW
oC97hYTS6VsVgmxlnrBDzepPVeOWlJMRdvwyjrfD7Kdn+f3eWc5y0bMnZ7jz
HxBuAp6TexueXpI7tAEjYQ/sRcfGGtumRWv+X6wuVCm5odyUYClLNWCEwqSW
8jXMjb44sgBreMNoiE3MQkhbF51zQyXS1+fSoHTueZJJbl45dSWYK8LUJjUM
KulvwUi4Wi9gaPUdLL9jEwqSFL6H1kkeHw6CaNvVVU/Bth/EOFvzxVSY922g
4p9BkLkiYgCqRsQGwy3+gduIvGd6E3jG1fQCDO7mLKlrpfX5BBsqR6FAFQC5
iTklJaMX5R/ALJ3LyA7jaOWvdm0unGCjT90NnJKI5WYDfyQR5sJluVT08IAa
rHrqbwduFU/3SQvq5lsjHoZT059kEg7hO1zkwcJj8t+cOImgj3t7aFmnVLwu
QahB0y9uOxwNOqxYmiNz+6RVCl4a+VT7jJmz9VY5oQt7La//usjCEHtY7Ywv
vLWrdrd3NgXGvEOOG09ogGGKN7+XCYF5jz0+BiKlTfNPH11EdCY/hMGdU4oz
tPv8M29qU+CkSGcGAO4u0bE/8a9XQieZYEath8UPBF0vp/+VTyqL/1I1BoV5
igc4XAkB1RdcVsjX5DR5bOSdet3Pnyieu7Xtt3ucD0/F9MZv33L+vnG6QiFT
QjQUTM1nCb0H8ECQ1Nkz37YukoVu+mJRhrea90wNK5kypEvKUFsncNfwPWmV
SxBXR7h2hnm9P3s9LJDe2GTI/t6DQhF1NjId1INw1/nNBxgHmQGAsy63ULtY
Mhu5Bj4CdDlDut30lRA4y4tBK36MB0dRpNtbcbrUXYsjWwroiD8qz8ZX1jjJ
BVbMPBKNAHVEtf1rzD631q328McRgylhLLv1mKG1L37Tab9PcgHCeLoE/hsq
NSSGQh1Fkh2ASSKtRABdI1Vn/ZaeaVMVTToC8H+Yj0IJNfR9G3868/Dpr/md
v2EsJy2bGZJvcUqW5PbfT9YXQYBRoGTmQIzM2LV3F51AbfqJBxhDr6jfuWyA
AHOW0Kgd8e6FjUhZ/BFmVF1nRIbtHNrM/XhkuyqbAkYUr0epkLap7Cm7hYz3
sB2yv9rWvmStTSTjgmi2dv3cE6Hlj2OmceUv7POIBnEwFQkbl4ODaxlp0DYG
bWQTNJWFooESYOzof6MVi6Xl0jghJl5f6aCVs8/QylMzTPx69Wrshow8i5py
PI1z81dyZ1EVciG7idtNyaRKmkk6y0GBXaNnAoN0cmGiXQ0GEqdj8Ru7ndXx
8Ek2R7mniheZ8sW5sWp1LJKKR9Hy26LTMHeeGSXXLl86HzBDjcjIlOJLeJgA
mhWst9etqLBNVrISqTfdqBnnPkLNgfPIl4oBKGstgbqwmIh/QKe911D8EbuY
5XocY6ZRQ/yPypPovS1Y7JC08hpyok4EfSr7DooUKWA4csYZBz6s8o/JrOVE
j5Z0XoTb4H5qVXpj65smJTF/n4BE/UwvwztRzCR99L402Jq3A/KzdK9m5cvW
1+yZ7AaLbuTxOSAD8yslJ+FVoqdaCk2oJMbCS1dpC4p+fKKOFZC/kf8LjQZ/
UfdEV3kmcNrGPFf6VtwPuJ7UEvwiLbNzuRRLHZAGCGWOSkj/rdnmq3XhM0t0
FDdOp4VGWz1k9R1JevcF33uHHF5rGp4UdC36CU5uWcUstn2oqkX7Dgv0tYN0
/JyhQwKtD9+UlNodj/jnY5sO5V3usOMjrnDJilg5MgVRpJDDL5AWjh9Rn5Tu
AtdfS9Z7WOaOQcydEo0B7vSoiQIrWz+PA7vZNUyYGNVD/+BfLVRr4LsS2/Di
z8bYUam3TrN0mLRrI4admmBbr28/H48Caqm2EFsSpknNm8zWFQoRQuXZWga6
RT0tNXOR2N7qmB2vRu0rjU2rQ7yQuOJUPNboAeKhGJf8R9iUo/T8C93p/erI
FRDHzFxIdniAmMhhdJzL2vs9C4qX62fsk6Asl+ViMVfk0/H/ce5zmDPkXJZ/
zdtu3Wraz7ULbJ9rhfkfI9BYG6L8KmpuNv7lWl00OLtiu3WiOqDZZYLpR5H5
pxg7sfCrLWxogZ3dfd0mUKe32IOilQ5gKYWvURYo5Dj7P6UrCWScX7ICjdZM
Gukc/McLE9DvKt/4sCLMUW4lIxeSAT18NTsvNsFMzkuUk3wnfGEIsSH4CIcG
XCUIjzAtg07syUm4cf7UjBnI0VyyQ2hvE1A7mmVllIfxWSGPBDEUQDUE0CTw
EXxuKdIeYFFRSlwtyOwhMzbN7errwcmXbogxpI8uismKW4AhcwJpsqY1AFNQ
MjkZDB08at7PEAMv/MOSF0tl8Muv8xMg7kS/qfbL3z+gGgaLazG9ACrJ0cAK
XuY8IK27i6Ly364h9I8Luou/RxbVn37l9JZ+Oo3XORc6M4I/b+DjocaGdFVQ
5rAIUBHMy1IvpPKH15tZaS7vkyM7HRqaPdu1jVIiFyZdDR+DTToNROG0l8TF
2TAKiYfHZMHv0uqqrLJzt8rnjm7iYBkBqf2XdsrxyBqC1CJT7VtehD2/TSGm
4w6b0bMTH9DspEn5y9F/AcaUU/dcdDL547LbaktdTWefB9LCzVPSfAQMVRJK
DhuZ06AAECNUlISBc2ZC0heaEHmimyMG9XEdjL4pLuZlLZlT7/RamFn07PCe
w4N6K4+a7OuWg1gI23+LrTxjxqt0pmUpE0JV2gnvnh3OekKlHBJ5Z36fUVbm
zsv6mplspchALQw5BxVUvye6lPj64bBz82I8q7U/bMtiNCTUNKy0I0XmFKE3
NC42RC/hmMuQITsZJ1o67Adf+7KOgCKU6SrncyT1AC0v1EODSHwQQeW76OK4
fhpePCuj3l9PB/WgrpBQD+Syw8e69Z+bdVj9M/vnXuGGGOuIoOubVfxo/cjg
LYUtH82nK//aFgijgEQUEytXm2cUr1pSVeZtwVApBnZK9m4PLwVJluyDcCy8
7WqfM2D+nKFEmxno2R2mAYfzZQ60JScRJtttFaJi7omI+hukDCKRWj6dnx0m
fPd2tK0fulWU6LVV8bbn8uJJGR2fVP4dwkWsNtY75qElCHjozC+8CNK1pdB6
/cBle3I+gTzSiP9deCeN19o+TUKMapkW+mZWhZDEy7KL5N2dvEQdIOESp2uP
0/z/aU90zKO5pMOA3kT0ufqlHCr4CEfI5qR+lWVQnOxicv+tAl2mcuq2pFaX
YG0y2C8zJ3CsWfJOy6qoaKd2cj0GOyM4VJ8+cPq9z/Vxi3rl3bwUkwk5PIVU
/pB1Z8LDvqfJE0vCRJrUAGz0sF1F2r32XM9Tl8nlM/B1FblM8FC8RXdxh/93
ejUwXuleBcO3LKPA5IDEtRJRKOeYWHHenSuLRgmmYr7jRjK6ZyHNaQfMBqlH
cLEbK6zUVnnkWth9TqVZmRANaSxinGY+jL/V8BIUWEmHGPKALmrScWj4Glpk
hPKKb94sb7w/eRUDdnzqpx47ZlPP5B+3BEZc4dTx2MNTlJLIqWJoBjHokX5y
eAgCF+AycdELXuwt+9P0P/2eEO/rQGLeQDNlHktxI4nJRyxnZSbjO3EfmIzC
nw6Es9+bwvjMPlvxKKrMHaKk/C3CRsFKsAOB91YJ9q1zOqOp6tLKRZb1eP6C
0oliKM9DxY3EA/eeKZyQClvD3A5BjMp3jsZKMLAaeE9iBph14fB8x0R7IzQb
ga1J5Dx1iW815TugpcQaWbkdAINcK2DYzpyxVSDVU6jxeIy+XuD1EtKTwm9Q
QORwyPJT9aSF8BXD9bpti325NgXLUlaeZpTDUs1XKxMA3WTXeOgNO+98dByL
6/TROkZ0drBUJQH/niMZO8VM2P2IKyQNuEEviLFz63cwzIPl1fljT8P8cVuQ
SrpPpzs1KuwIf203RU7CGD0vWy8YNyWlzxf6jNLJT7Fr1cGb6qfSIuTYxo0J
XFzgBUFdlW6NunKz70ux4SFBkbWUs5Zjzb/8OeqLNNevrkxFVDpnvYcOxcww
FoqRvz0LDBSDUqkYoo+2c86f0lAjQacKALo+YIAS4aFRXt0+jIwIVwr2b2S1
9yNj3CdHH3Utkv7QA/2ob5XzaoSTC7DPRsbQGzcN0/s2nPlPyUN2gh71I9nG
CUCQTQYEOImeDv3E0B7skeNsA0jlH+FT7xX6EKjICJYBZeYQS4ouMKgGMHqn
eBC3DMEeMI6RnuS24fGDdglvx25s3ggHncE48/Rc3Z8+D4RE9jgbL6nGB5cV
gYbsDp3STz/ni4SeXMYnIGpZ01ypMgje0OhjT8Hog7DYuX9Ad1/HWVfbQ+D4
UEI8TtRmD0pbSNMYXxfbFXHt96my0g+NqnjKu+p4lssP03FNRXJ7zbDZ7yhM
+CVQAimqedtpC/K4logNXyPFEQ4ORdVJQZIxsGeTSaDnR/sVf7mo3nzGn6BR
cHAQyxn4RvXOUbYKtpYCVSMbB6qEt1i3E9prtGIGT0pVQ3AZjobLdGRMNPRl
RqUBwI2CmlOQyqakB6ZMTzqziRg+hm/hBPY5Z2Iq4zUJPK5XQt1PLrs+npUG
zH+ZzSO2hDgdOLNpJhE3am01RX9eg12nuo6Cv2i0m//jAk2FRAerapVmk5Fb
OrpvXCC+cnHXZ0xy2C+rZ+/PZDXtN0I7L14HyfHZEDPJESihBb3XuFZXvZsA
BBcY02lF8TiVbPhakQ4zG8+JrstjExz4WkXLn+3hy3GECt1ixietYwrFQkuK
eF2ogT8BmtxHgNvFRRcOuAkoin7Oq0ovK+RvuuObvoJf38usz7SIzzMyNNdl
ZnbSPj+wa1GTUA0NP0mKdmwY2bHo6r5ckdnxGOMmBh7v1RckN9mhW74491fN
oAl1KKg/L9R6+eoY/3XWyAG3flMT+5mgYIwG0GeMWZuGT5Ux3q6fFMx3tXKS
3pMgyaoza/2ySkdvCrEINTaQ+J1/drd98lU2vC1zFe9DeGFphbe/V3ct04yb
L00Py2/wkZlFp2BZIbc5mld1HdRNgIz8aoYnGY8AU8Ekk5aGUNkzH/Eg9dXo
0wjXjyA0stDtclTwMKXiYGH2md6lE0Ys/mQMPAooCNWuFUi8O2saiboU8+70
Hr3sCKPd9zy1vXW33p5/a0tcOMznCIBM4kG0UtqcvQ3tlMezcKJgDXBHHBrb
qgzfmjN7UoTu0uaIW7OxppJNhso6bAOPurw0nenLkIVuFdnZNku/WOlU4a3s
I+WVEsyJ2o2YxnEA6fVoInNUROuaXdX3Hio5cQlTspIMvXOTl38AnN6Y88BN
/wCjC0j2CbYBCoFuiYLChrV5DTCVX3N+PHS0jjcwyvaKxjlobKq1OFzjBGT6
1SGDW3KxV1z+kcJZQ9PZsX4CL8oTrvwcR4YB9+KMTiSMxO7/zrzzsZZiw5/7
RwdYFNIBfG110bT5eZYPuUkVbA24+Ve65AuFVgpec49GMWjOlxsdxgfPkA7p
UoVcadJIcu7TqdIHo0jpQNzQv+wFY2iGIcHlfC+6rv0sarGRQa4K0svvUlgD
57eFxWr96odG/UHLSs2F8QtwIO8LWWIN7TEkMqvXDybkSYI38kRvQaqLcfhP
IyoTwLJAEKS7uw28HHjqHKxBseliSfLRU9oLHpyGpGbcMQpW4l6OLd78WWe5
LtJ6F8DMVhTKYyf6iZefxQvUX/mQ3Okg5aOAaaIwdHZCNeY99mkOkt2nmlWh
/8aKtU7nQ6xPk79nerg0nTCuHDXH02pultX9irc94OZkcJd+vIITgHTl9lZD
Sxo5Tl6YXFUwn6XXHJxockPVFqANfRKIUK7/jCPo565iHoPVYasFCIWmyxVp
EyZ1WC1Sxj9WEyVCZZQ/7QKvGbhB/H8GdcB94UeQ/XbV3AM3CP1B/Y0Riyh9
V5Oz3HUgAsH2YTlHGyfOSuxO/oTMQGmI8M+4xSAQLUl62LSgnFq62BUU1WgF
/DkhS8Af2x2wF4Fz4J+nWnO+9SRUqOrDKBxcnyXncquUG73gtRWKCpeoxhe9
C89f9zU2rCBqsfFTlkDA3zIypVS5ZD0JRxP9GspmsDZTDZnWeEEDWk373/HN
dpEXQDO+T1xsd+2eQVeb33/15RmjpeSh3gcpdmGfJDtjtquPAMU0RcshnDgj
t1q+zETOwBr7C91I8l5xg2Bnt9aPvWNgcF3HecpG9bh7owDwnhuwB7U2tXlN
QpgSs4T4XIXd4KDow/i5nd56pjqPQ4+miyv27Qiwf9b0OtHXUMQrS4TlxvHR
dRb3E3PohUTvyrTuAUCYQgGBc+bUp2bUpab9/sgf4TohOat3LSg2HQ+ONv4/
9GhLLBClR6ryzqxjuwKUq5rspodYnSTRO5cGqd2/9vdCLHWAdNXNhkn28Z69
4bPKY5TLElbR8T7Ox4jg6YkH2nDolTIenAO9d+DZyZpNjTqPnXTX0uLYeYd7
10puRV6JaUvlO13c1mTi9bo3KtP/d+BlWblWdSKfRv0Bj/Re64BBJ17GFLXu
ud44+BJ/gtP/IoIPzS3RckxUFOta/SXyrMEmhxLfuNWV80fL2z0VFS8goLiW
bUhO85oI31dQk3/y0CsdjmiH1h/LcqvHlvv8mJXKO86fqtLUMRDxKHHQUPN/
3Zoat7Md7MSPzPsNo5qqy0hcBGPiHY4BXRbRGPoq9moQXtE56v4+ytzkSNCU
7c5MaLwbbVJVZNBXMeZNDI3UxEL1+c12vW5dWv2WdB3cCrpi40A7rc9oN8yU
KW16kqgAiZz91iasqEV3Tsd3A+fDzmakeJrtRx7Xqc/I5Pf+dhIPUrl5Qr0g
sMDz/avYfAoBcbeXh8ugbpfPWoEiU7a9jeMehrAXBXn1ns7mfj7mCHiIAKvn
mUrCQU48p/iH2L3/jL8GmFvIqN0kJs+v9TmMn/mijtsBGA7wCXYc/P/Z1Q3a
rrThJwg/2R1xC8qCJjyLkSRLPh9J/cnuqjbXFZxM0fSHeuYkOoTM4FdZf4qu
Ptb1mrgyCEMpWjSz2ozcoEEOV9ocXt/Z6kMJfRqbCOHuFrB+72khYBLJY5Zq
oRdRcc1nakNgso76iZ2ZiUSJgH63REBepKeOe/qB2GSFf0M7c04MiNsaP0ev
7Oa4WMp33fXRgABqQ7O22YE+KF3dF7l9ZpOMzigt6p878r8XgkNzS0GWogJo
9vfiq4i1eoPTnV71cU9BV/zZ73OOdZc3V6XWAJ9o5IdWonanVwfCZIC31dRX
EKFV4LYGMzuNnbcjHMszgm29sBtJ3LuMKbOQI1bd6RXFm93d5kCnmA97oOFy
kW2hNuiVQC5a//msoze++56iWkxmdXnjnhBmG1mNp86t2rsjH5+ouIa35LTU
DBehOZcxQHvwcNqZZOI4R9j/Jmr8Kgw61RC6Tp3wf3VAZc/Of8GuSCqx4O7b
LmUJr4hFUy+H4Z6VYu6Ca2nFbBVt2mMaC6YiaupY8UzFJ5vjgwo3jRwMvd2E
RjIZe/JMF4IAwqnZFG4l2H6MZ85C9kZrkRwL441bLT2YY0Sl4q75JORU6ies
0Mo7qtTVMwezmXvajnHhykwxO6T3hf/pC3v+k/BFddlW8Aa1BhFxZIh9ZQm4
hvTfQpiCR3QZb8HXdfnP0ECkm2jqmMNpn6rAARbKqVovG4ynn2MF6mQ/LNmU
SvlkXr9k1e2L/xyqN6BfPnzCg3Z7un+fVKgBtKAvzCtNFvEnda4ctIwGEouY
gtgVy6oKJ7GImzIgONxwxlwCk673JpJ2Ic9ubO5oKJwJNntx4A9dWHiF2RF3
+3hmJWIWUFYm9MozRidgq4OfgDhImUqDl8zHGcP3y1AXwlr5KA2ULVuMD0Q4
3VQWPo176w/qJMgfFraLUdT68KPw3w7BVriVW3C4+34RnxcK+mbAfSxC3V60
Nlq9e217Jwxibr10cbONIFKUzf+Ie6BKwICm0bK5lrswIFDkFpvelKXo5t4g
CIhnqWtrcCg3HULYt5691QF+0IDMVv8BAMdj8k5Pig7P1oYedUpJxo9KCEfr
BQeamAv4NGX0Yx3b1ajr91ZIDSF0sUrzLgGsT9rqI3lLBoXc1axzT0nyVGWm
o4K/wxElYyaJHwiWHeCPeOzgaR2zyizFDVEXd5q62bVaKNvFVnp38qu/AeLs
xFXWdO0ZK3wrWaRt60T/xeOJiVvpO0rgH64FZYfDE/gca0+QuJ/v3eearsXi
NIswDjg2w9LYne/d8xna/zAJFudlzAtmv/d1+MvCiM5M6g2hRDh1qAHjoeNZ
85vY5Cl+IHCMLD6v80T1IJr9UqSVP9P9cMAOFvbVA1y66VJQlsuGeBM+7oAl
hNy19u1epYPbqN3u5469AjFhF2AOCh3ts357t9RouHSsWq23N5xmJvOY21ql
QZSON3NUOBcT/0MgUsFJqeMVvSCbQyrYlEQRbL3T3fAUz5KFeEXej6YteXnZ
d+OE3S+rEl9BuXnxXfyZr9AKcmeLk7L+zFV/dJB9lgM7KxsxohHaJyV/X1qO
ZxF6RnkJAjwrVyDcF7HmLfTqewtH6r0SOaLHTmvdPDaU433d4UG2HQOaVtAh
MUoqCWfGJgLQTfWiaCN73uF04Lq7fcnDKYXqi6keAxJsytui72uZczN1R5uu
8GcxpwqNPBYYSyNUlEA/90ddYIWdvskB6QoHEXFZCZFev3qTyI75RzmQj/xj
EO4ssIOu70xCNJN1atpDxIcwVENNbO4+Pn+4e41yay4z9rLW0sNLDpzPTKZ8
0/DZmJa18I/PragVo4b/I5pP/sQYuQRlroZBrr5teH5gNb8Ut8G/e2vnFmm/
cxrF5w2Q1kDNSelaI4frIY2WIYLYwWmjFPRRTQxPpRoaSQLZ9ZKb3QnbEFbi
v+HWICbUgehye0+fezbKg/ueguiE3ALjeCnum8KmrETKUmpTDXCP9DgkN6Q8
Hskt2RWjx0TnwMbA9dK6RePGjzl/Kvu3VApx/Ft9mbccWzRA+a0TXDzVFANp
j+UscsTI2baq/voTJGeZc9J5eiC4XQPMMfyD1JH5MGLIx8SCXWyNVNbDmZBX
tA8CAy6W1qpHkWiDAPUR++fzYLNAwjrWsqB2d4KIXHbFH8lpeEewMzEzc9Kq
2As+R5PJLEh7ZyJo+ABnATFdppoBqzxWRIRNchHboMg3ax7IMlyJSm+bC7Ss
yl9PF2XPnROjZZGjZ5PYzoEEWj2JbrMkdn+j2Hz/Y8KaYHeWX+aHjTJIkHw5
oK5FmEUTR63IJOTiuDP926s1A048BPlRxZr8nWONmCpucKjvISxwCFLnh7zK
HhvLTkfDW5Zij0xuzoRkCZNDYcYnBNVIxNhC090EsVKG79IzG2UeYAXKKpPa
zt1q7eyxXWwpN1FktPuXJ9Z3WiRYEeBfvOSi8Zu+X+xfG4oe4N4yU3Sz7sR3
tmYT0yqps7rgRyLqyo+kwh+zWT9NUJpnS/2ATBMoIGGhSfdnb0V0IhyLwQ4T
EunydfrVLDBmnZaTyr6el36IIpv7rn3lRc84qojLGsvfNoATR+MJzetIA70k
szStTSgFU7sswcrdes0BTY1m8Xy3IcwAlrFM5FU7E+zX0d8gdGPcbMqljHOw
DH8qrrddoPXEald2ann9MAk9//TUlSPEobTIqc1/ZNgtVmD2zoUjtTLiDhQl
8wFrMtn7K8hy5vHm0ArqB0i+gtBq6xRWKHy4avzKsDYpbhDQdwJNgpuMfSqD
unwlaciqpybqnDnGTjr5aykY3NGUYE/fZDwmbXigDjZP2sSXKrsNR7VUuJ1H
frBK5bj7uD7P02rEVPhsD0fEzlv9EQRiP2TMqqc4P+CR9dT8YQo79gSCqXlx
akRF4zH4X35IUXw1GhiiY5xqSKZe6H4Bs4Jmzxs79LcWC2VpadjU+3ZiSFMG
fte5mmDlaqILWE8kFcidjbHXyySRl7VI0UyLMZ/58/Kcy3YY6FvCTR8l068X
udM+tMfofBVgRsxeceRo1seoJkrt6LcK2YizzIjirmXmTe2YX0KDJxrHlhvW
9f5WLBufBZ+mB4ypi71b3KHVnDncf4doKbpXZvHhBloL4IfsJXsiqaCQym1x
l1x8NwuquAh5P/X6gO4nCzB7nIViBnyiY02q0tfliELwjsIYJXOw97K5C5Pt
/SQZouVnPTdZlAC7Vr0NIyAJss15MvNRsE5fWi0uU3pZsiomyBqRaGAC8Tjc
CJwQ+zKCA0E6phlu2oj6aaVIBI//y/3eA5zu/lB/V/jw+IPaasD60I80EorZ
DIz/1xdLlEpDcSESZ3KkgmnvqmdQIT4vYRVPPPhBXavUugesyo3q8Wejubgn
vt6rjcr1QdaLxT/9sRiCnnojTho8aiK3AUFXCSaMQGPeUmy0WNY6WHeIt2Qs
lg1TNQlyw1GeJpEh59xjghogVUs8pjxkTzQZr0+zD7cFcnFUJvMNkxx0m8oD
5JhOsEMXhgqLc6XyO2Trw3ucenO4x/8e1Pvf2qagw7vC8MQQ79v5Qogm7W45
aX8GuRXeUHiDu/DQQixWVK/cGIEM9O8P3sQNaMBMLe8jz9OSRDVCBUuk3yGM
+BsCjGOSg/9NtqOyYz+J42nO+39hsrZfV10NUTHXIfz4j56A0V0nQXZfK4W0
kCkGVWtzerQwWO9s0BJioeoUxAeL8RugYUPdYt1YXbizM9VoIHmz9jJBTh2c
ge0nJtMk/BCGOmzMcXyodYpJfI+c3cTITUgcSooBlxibmmO1mgSHMyjj1WVB
3tIszuETxxepT2eT6JY1PAPHeaVbahW7eAZi/tgdp/fEOQcrmwAdu7QFUHTb
xrrSZewWXDYCS0EuiiQbYzL21c+Yf7qzzP5JVlGBHBPo3F2EYRx5mzfelsMV
98j9DOyEtu3ChUsOuLpmmCBtYaINCQJnMe4aEOmtK8xCcFo1JKtYNkoe60vV
QuEqCee7zdWmKepyg1SiTngDxnDlD2nbEL/Dm41b8qVzTgTqI9sDHSk/gn0N
Qz6Q/FA8FUaLh02OoZ5J009nbnoYKoMrVx9GocrTdRElJI6vR3qcZSzKSTbU
3IemB2j+/xs0Eid/ia+iPNmxgLaA19cZgDlBWkM4LdUica8IQrO6umm1+iNk
WR55oaehwzN/kSKwDG2OKC0pjuQC66fk+Yk2WceFyreu8cV+z+j858KfuY0w
Ldy9EP4zUrifREaBOO3LxopYKQUL5PvFxd42cdfBrrf8qbDwAAb6/qPmAvPM
NFFMvI3VOcjwaqn0MacBnwkjUjuelGCvrQcnaJvKFVglARDRA3jndf2c3mcT
imjZv2VbNWS/BX+VM55BVN1Ba4TUojpbFMHgcQcIPP9FO+S8UT1wr0bSdk5l
gNhktyPIsth0niOSzoprnwWr+vTMUb/9vmLvI4+WIpDcG1ilTfzk2yr5Lrx9
7a5jXbitlfBVoqEHS27gl3SLbJxz2GLvGt3sQIr7l6mmxztBz0pru/qdBBMR
7u+hVoXqriCpy40H648TTfZ4x5BuPbMf8QdYH6nmlb4kSL/BZAsAY7BZ/kpY
yzmHhJOwAa0ht/fGekKEi8Ec7Gif+Jzky8hERUR4igyrfGIHGgoTOv3ojDhN
pspVM+ZfeZ8oJUve8M3bMRURLuiqmcANoFwOrXS2VB5yyrdVzdwDOUteWOCx
6c328b5Qf2E1CHhop3XQelZFbYH08I3zvUd1lPtk+kbaDla/u6ueMNQ1Z0DJ
BxLmR4kZ4g8hStR7/dBzxjtpyg4NapCJPiLQwOtC/akC3yZrAV7N0LSrgjaJ
EaJeB6+W6mhQq4emduxwYiBanTZd95cZcVR1SPaGIGLiEXb/s8B8ANqet2aS
Ik5eMX5ee/IxmcctHTW0vaZ76tMTcj2VPQszE8OZDbYSU85UXqfREITKAiK+
2QiDO51jQxUatMOg/80+Iac9B985laAL3Cy88BpUrkde+TCvyTwkGx+TWGLE
NSEAvSQGTJnTeYpd2VA9GbxE/7lUpbSO7CWUpkmh7X4peyzK/0Gr/HJhRFvE
VvWa4Mw1c98/CMTLZdwwmC54MsNN3ljgFKfX2TAup8FkXmZ8/CK8FvqUW4f4
c6af4p3TNNQN+WFNYoVqZ9vjU34FPaF/QOzCvsNbttpTR3jGoLpl6hdsmHCT
0PnxtuyRUYYSJab/gIAwH3AFD56QXYA+HF5OwMZOQt30F2L7tgetR99AMXVL
+Odd+oYcqbyalOqHbF61vSFrgsBtdyjg5GWvgLu+Yyi10znDXIUMTWK2EfOs
hHiuf7K9ionJT4qHGaZMFjzT365Y0cbcQ20eOjtsR5ITWYEA0tQekO+ksFdm
Smq3XqCKh4szgtCrbrp+wF3XU1m+C64Ssom9X2oXRuXWNQdB7+RbPXXC3hwB
hC5lUWTYVHmXP0OpDBkhsOdPnsb21y8TSo3YY5IjsKlrPzLRkS/k+46h1Qkf
EitBETfI6rznnEMxeIii7mwY9zY2beNXyNhhVDAu8nuD6Zn/fvw7p5oRLPtu
af3W0uoADITVVbyB9WFgkLcVuO6ShMr08HgutBS/yw+bFtPmOrDESBO5BBGJ
HGFqnci8cInXPOeQcMj66avI0anWClhfjGHpJC3o7SIq0OILMnz3F9rcBZwq
J+rO1p/4EbpzE8piwew1E1Cv5mYxQgeirfcDiFIHRhkw9caKiMLMc9ZxbPjC
B4lyegx0Mvk1DtoaYd8IyAKW/RllgUFi3of+SaRgs4ztAmr37i/OXlv4an2/
Kz2lUP/tsEqp0FBTVbnl0LRGHomCc8MM3jtf5y4O5zaI9zSfU1YEmCIjaxK8
5H5+omWAxM79C3GKue3nVlAktUp6CFsD3z2BDWOstyMCpSIwhhe8VUVC+grj
bJ1ASASuDGKGEiLYKfAAztW68voSn+ogbJXRNN+/eMpHATrD6a7g+afy/xXH
UUzM5Xno+/wwqHxlGGPqulw3VkFzEHSo9zCDWiHRIK0D5XNww/lRC738pu6q
C1ayXV5dPpYGuDx6kxuMqjvfNDlVpJbRfPj8Xpa0ygsgijW5xHiXEBlzPcbB
uFu1M2zZA82tQ/uR7Z/1EaTC8Zsag3hQFEWpfnKoFaMv8nDQ75SKpXqJogGX
JLT1eqMgsWdkTcuj41zJo9jbQAdR4io1U5BmcdREk7d2qLmnHfQXUjCUz5CR
C1kN1P3zc1qCNPM1W5eZ3wAlYO7JSuU15ZqFh3ZVyDWT5GVr7duY6V3OMmb3
1FO0xVBYH/4q2+vI2W8FGlfmjny7DMtjGqG/8xgaOAyYgpFOskKU5ER3PzMC
vyl4oPNCWXyaQqSrS9qkVgHBl/FqlTHnUGmXsUt8UVyr4YdBwPF9TuZ4zzYv
PGRpNkpTz/ChAiUxG3Wl/9hkzQDeke2dE4sdaayWAE5aRW0FCqkSfvNIMOjO
+pmB2TOKxf66/lsHEK048n0Pb2RBQg6SyrY8hLKa6vyZSbYBGBsWsqKAGZi7
52aHDPAr/7CWSLo7t3RDfQx8h+jeHrEK1tyEx9ULDtW2UgB0U4UyO6iKdwtx
59fwTxsyMa7Ub3UgEqIBu+ZYx+C+9DQx1WXBWNu20LIbLkFszmLHqsICSjF4
K38Ekvv5IM7hb/g4hkbg4JpMqiPgl5FBh1gsaIeLzbnieMVElW8fUS76vnlX
a61yIvKZ5Exo9ZHt37sdcqUepka79GvrnRYk5fPHvVkhOYc7nPMohrAj+JYT
swYW92lACYuO+hXeRQaOkn4Wq0HswkgOoyhHVykQlTCORB/fY+5efssZEEW5
9Xi0z51H7y+yOwuE03QUMWHJqicxO8wPUYK1pBPSJuTWLNwiUSqyJfVlgn7Z
hYi0djz6GX92VCkyKVLWYXXxLFDiU6aMf96mbV/fM7C38DcmYQDx7/GzbjuC
J3bSwBs64mpA4jboimJijw4Z4mI39AF+4LpLTEP6upGyXpR4gHsbD0Fz4ZoP
XexH7FdGnS726T3gTJnB3RzbzpY/I+dpUsF15quy7ZXrclYz4wK8+CrxDK6a
SQeswtdJjBLftGdYe2ZVD2KH5o9OJtgeae/XZN1ExH/qHb+xjITt2OYGQ/8q
CKNMqpgDFv7Mtqru+sl3svFS6VSIfHcnFW2TzzGCzgnvOzlNjBaZZ79NQemu
hrgTYO6rd6/eqCTqF359tfv6Cj9wkw9XzkZf/dErzNGU7S24YSEXIP0Uezuv
BKr4ZPeYvQKBgtYIYOQ6/4SmzDKegk451yfl0jR9r8gzKSw/ISYpUCYSSrTw
TGgLzqZ4Y0xKlFp56bgTbk6SVrpoIhb7jWtck46lnr66HpMIAac3We38n8p2
6w7GCYoBO87nbXKflg/Mq5lNPbyz6dFE4LRpci60FJpytOsgGZ5JUvCsiLJt
Y8SQJ/h2nfTHWmOXcf/w3ZSq0+fxLHSBQATw2s/7MgCD33kdpylk0ul/jF/a
K7WvX2ocNYxbJc3FUESRYgiNt5gQkpLQ5AltSEbDFygsvZ4R2gstoUY2oakD
R76MYydwLy/pBfADJ32JLuHhi6oW02JySCxK32mz/cNBa/JbXa55hrBlg5gC
NqfszGO/GX1Ug3Ae6WzwBY2hX7/sia0Bo5Kir2r3+7ka/00kUUNPgbuXRSmf
qfeeG+aGBkN2myTrNjvCQRr2Gf5WIYVYQf1C9oUPFOJrC0e7K9+wspT0TyRN
7mhpFpujixjHZT9rp4aT1MbHqTWvg2XVAzklbUCuOMxR+woJh+R7E9IXjGja
rzB/4IlTo9LWHxcuuup0vyruHsEqSlyDk+HVchoRg8k32mgwUPmPIFooefHP
j+FGoweNTZSZTTG6Z5dVaosSL8/u/nUjchSDGvSwg4m67+DQqi89gbakJKIo
fepaKpJvJ+vPNIYEKzsBF6jHNeR0BQ77Dgzz9h0LBeePyClXbiGItqKH1D5E
bFaU0juFrVtLXN6iJwT9o9LEM0om3PqZJLzvYRIuPAfeY/wt4BZvJoOFqHel
P2gGQN+9C5F39U8zl/WFg/ctIqhL5YjTxYoX6uE/923Ayum/C3Lx1Vn5IARv
g5lRqlRC/96cK0m6VH2QhR0c7aDxPcQ7vhLpbaiiRuX5l9c3SSB1sJ6Xbm1C
AtQz7ZAKcbR3k8Y3ChZ8EY3C/aDRHp3EahvJqG6bCru7vCWLKLTUwWVAxvX5
uckxvJyCb7FPYw5UV99y8SMrME0PgTK+rNTG9gYXNvBT3WdqI37olBbzeuAY
01QfKJZ2wEaPuQg9jO3aLY4z3ro+K7NNVBT5xSPhR0yMh8OoFBpque3IXeDs
2kbnGlH6srijnpF8OHmQD3chcyzsO+DMbkf8b1c0Gq4tmyACw9Spdo1eXExd
VFQ1Amgp9+zPhDXMdKMzUTxB50QQmKceylohEAuqGFShvejtFSQDtw9Pz2Zb
N6e9oGWwszhdccoTAR6TmLuWTFaxOIldMNocWiv/Mdh/mxN4D9XQhfH/wxzU
TO8N+EA25Ja7DIq3yp7GE5FiIvbaZYFUfWLYzRNash938vwOII+UpWS97ZKF
YAklaCzIJDyFJ/z3D4uAiMU/JAv94jGaYRhBLzzRkasOGHC42Qv/zjB2jlk1
GpjanS1hT12v2e4lewaPV/gk5tFM9J1j9CmnYnYqtvsZdei5xpW4ke+YOdCF
uI4Zzmi+8EWZhObnm7gNt/9h95kKHkUVUjs0mqLuBtQ0RZjBVsfaKLZIv/oG
cVBXaEj2rcjtlSvCz4hkQwDBjIz3s0RWnQhZ5BWYek8EpJMqCgcWPignWDab
4CjJO7iUXOrXC+xofdBSlVSGXRW2xzlbZS9NUHt4u7Q7CfjPVp21IYWFEY6z
4aaql6BCM7wRcNkNlehvh4cuI44WGrYeXOwGsXjPRbfU0+WyqOiDvFEaAVHL
t6M47QpAo729geo2KaAclAT4HRJ4VSSa18mL8LNf8x/PmN3YYHEb4GSD1i1H
UvdeafIlJNsG9TBztIvoE+ziaXAh4/oPzYscztxzYtIH6Y6741a/7kGpVsqB
saJ1zdO804x8gRaGDRHi471K7b1vlJ5wXK6KOI11+dJnYJN96mONga2xJ73d
38ODtWW/Hvzm12cxjkGpJyIlGmjEHXHAPH7dvt2ZSjI62Ud/wFxrkDS5IRqq
8GcYAnAERyAKI+l80vXyvXoo998s6XVer/ipLQS5khXixLlhQX5dhrJd4ZmI
iIf0FktbnkIRM7er+VhbPWTUi1p8xoW96RbhVo2k9PP4cFB4nnySs4zHp96t
0G8KoIu/gXFUrJHOv6farIH7LbXAWrHhikzU+Np0z8zxnYMuPdKCnyornSEQ
MaB13MzyJ+S1xckXgOiDtSHcGf4NQaoKxCIkPg48co3yeItVefwhQ89K54JB
CDvQHg7kcekzo3Y4bAgJQjjNXjR52Exy6jDN7ROMqR7YTKLrTIEYYOF4wgIM
FApSFpNjR2BpcN+E0P0q592Y4cJRjHLPyIfA3NXoSetyhUV90FegIi9nMba3
y7ZFuheqdszv9lXq3jiiGcrRqptW23NgHOm/E+uTKKwViMdpXUG/FP1PYZsf
ABwkepp7o/LQ4ry5gEiwj9z5aiARctg2tRbOAWjtjq3M0fWenstygG1k4QVM
ftSypciKDsNQhTPbfqdFiy2uy9+LGbyqYNpYZw8MRjVhoj/dm3+TnXWaMngD
/vd8Vq+sqJGihjeHdLqMi+KIqW9N37bH/2UaFtsBpn5IuOi447b6g487PyVe
SuHlP+fT1Kao6nZEZDAmRK30cdGFaN3oiWyiuKrw4M1oQlyCcCDWBNWTIcsU
NslZAkowUaWlaSG74EIkSmQCmPWruZmLYx7OP++HHbw4MjeyV8RDBdvT6o85
JR+J3WPsdLjf1nZY4xXbWwUFKvxSioFRFp1OoqwcCtAAV7B54m1wQDt5HEDu
oVxBc03jsmKr5j5yGAwswFpj6ZNJyQPNKjaZK1g7Yan3fl+DK/6YtNHI9d0x
/be6VMLSE8TSOejHrEggfeW6fLmuio3CCRHZX0GGIWa+EtSMw65KTNpqc1ut
QhrE0WSlwBIQK15Bj8sEEGkxnxD1t4rMUIFm5690r5ct7nBpc+eYD9T3ibW6
mayIWcmdB85yFD+XZEi4xwuigDkUbB90gUDsbhtJH4dv5HKWjjdLiX+zMrY1
/b/t8yzdKvn49JO5MT5ZGN4/As11IRD/iJNNsdDyroOcLxBjrR7oPO1DMpDe
CIR9+OEl0UUHh+UAIS3Hw1LAfQEwNm8Dzc8G42MkOXMxeWItRPRhOI8zsf6r
bU4D92hZM866ugHAZsF3J+vvllqQW8cMj2q8IwiV3dIscrQgM4gCS+irYiMg
vSGFHS+DZKWRyoSkMy1WhSVgKJ9IcXQ8+eNJSgk3/KTCHxog3SHehQp29tec
iSUEKInOhyFrmlgQPUw9psJxmaQA2BCyKWCtGRNq2jjUBSB+bYEJFnPXOJNk
AKbw1mt2wIAF6JLlXxzs0KR+X2YxtLR3LUOy/XqtiTS8Sx0dJlLgVkPQNIlx
kncCF9K3rcwfbleMRkA2mnWaDF/5XFVL3m1mfzLhfG4lG4B3vzpa3NgnKdmd
WZksosDmkzonVeb2iYSmft7KKK+MR656IEctUHxUifRlH83r2XRs2jnggXuE
RhakoCZ08e4zHI26z0qCopVLCc2SJxgT3xXspbvwSb6242PCBU4gOU4ZLTIg
5M7bjzhthLqPhdknAAvVVDNx594rBH7WFhxIC2gDMkcwg2ofl3bdGgtPLLVh
Q34q5L8SLY8WBM5GdRKed2Ik9Mf0NP+pjh2YkZthXFCpvCgw+bDAgecj9sLZ
kJ4/fmPvCfpKpOGjJQSfXCBdVjiED/nW//Tsbl7wLrSJxx5ANcXoLC1wiLfz
s4bbnWv4oumCRE1Hti9k4Ss8y4CUaUXbIm8bQLTO+zeDDeEUwnvd7LZmOwVr
P71dE6w2ywnmuLW62eWNif3PZeHuT0bn0o7LUQjw6z+0ygLe2iWyx0GD+lms
E2IpDT44XVs0dB+DZnYZxzTje8JEjv05vFYD/ElzR7hlq6WQBfd0H6nNfyZ8
vD/5HMt0we1+3zKK11h/Hsf5QoVeLLdpaR/JDJXBwqLeEwBWZEEADi/Pr9By
HrqmvK6Gp6trkhVleEK9yCZdWD96j+m57pG5fE6y3Gk/BsZ6dXIJR62nfRCl
MzS/U3PMllc6nltsOAi/K1gJydiOSKfdEX0Hn7KImSbRwLxEwakG/GRN5G4o
F0c4J+Kizgb+45c95aY1Q/kMOJ/DX8leIl8lluhxfUEbdsptN12BfSjczr3z
Vtn5QyyZXlHi4iHzREnOtJokLQdzgOqHJyMIrIOeOXJQEzF0g3cN9PS+Sj9c
swbmTv+WvLtVTI6eRiUVCP69ONrD2pOYeueWI3Fo7/QWimmRPKJDk0VY/si+
6BMP6fdjkoa68s9d3bnzoKBjgjquwAjxMdmft9cRC/hauo+sKcp5JJ1fq6mt
vgXD3EC/tu/HmsIrBn0J3lT0vVdA81JCVEM1EQan0fWibUQmfkjG8nTLxkbV
mtCeck0ZrKJzXLU2kl9cTg/ykBr9LEPsA2njbQOeNcxmDLHhEed4ptXHAHFA
3a8hrOwJvcAOsDsJPTbVQzC9L+73n4qo+0R7XS5NeRHI8G9iVsBdfdWi/wH2
yQ1a+NKM1hVRDbBXzOOGRmmNrTfBm+qjJETJneMFoJuM1nEolAKMS/nnVbJq
Ia0U4A11njiS9u0h5SKpBrytqkiXSICIAKGd7ndsrImEZ2w/5Aqhr/IMj1tF
852Vqi0CeRXIGKWuf6BL6d7P5+sHsUYHdT48SqrIS4HuiE69J9xX4EHBgVpw
GLmVuW1ZMabwM4X9o2NzxE5/Yg+adUOJRA9RZ3nv5Vgo6wS9joEmybPcC0kV
TqsMByjZpGCrE+p64ZL6CcJdEXG/BRQUxpt0h4whW/TTp6OxOCw73qpmL/E8
BJ3z5NoTU9rPCJ7AcZ354/1PQNaTxLDiZlU9B9NiaqXET9QiWHLZ/kxNr/mA
IITwjkh8N0QZH9pb0iI6spvOYTXPzKLb72n2FVEEy/gX+PHM5FNmqnaVfbq3
K97ERGm+Plk2+pa+pMJW4lrn4efLj9IfCXo/LjDH3ba3Aa1V4tISPa/2sjj1
OWI5QcySfwhhzn67qPkAbEV07tLEVcPeY25yAvnJ+AVlTLZmE7hNWGq741p3
zepb+gDVcad8Djpn9iO2mQ2Ekrt5mEd8u/SzC0B5Bux5FJ0+5LF+z/8PiO2U
XiejFHpugIi547yuzJMngHHHkJWaEXlf0BcXEbHAanoE3lj8rGhcfYyPaoG+
LZ1g5LbZcdjG0wtDY+MvGdh0du7eRWRJa3Q39LRThxJPNpQwJCBArr67ZKse
2xb8JAEXFWlXJ7F5awc3bPZ23MUhNlJbajbYwVFn1euwRG4nT7FsP70APKgs
J/Urgchz4ACjkphwdcgbICDdej2NTPa76dVcysVeqkBcPRNVTsFseEX2icsu
4gnCCH0BHzYDrFDSKUWclpCiiJPvVSRFgABSsBiUu8xQ+SqCllVSauyociVV
6hgJ8dku3GqcmKGKJFSA2SSO5yb2fY1n9v0GeONuAeBhpDlrH8jxzGkJKr7E
a8tkhrqynDZpBPdvwufdEzMo+2Z0TFo+ETJqRvx8VM3Wp0Aa62I2d3hv5PkN
oX152pCdNz8IJiHbPBizGfWsG+FQBJ4uWzdmjalhYpUM9qBOsQPI3O3eO/UI
LooUdAhAGNKBVUC8MfQ0KjCl1EsQ+9LeULNnwYNuK0CVqXbqpy2fhSecCPbY
u3VV0LrsdVz8CNqDrO5i9NDO49MOkn6AwBr2LqPWKKhGxgAYcOsQiyhXDMgs
N1yK49wTzXX9B6H+IlTs+lmfA5s7bX4idnuIsXMl28lglLdCEcpMXSqXanqy
Ih2QHwS7E2Lj9Qe39OD9/3TFbg+n0w1Szxpt1WzzwG9mMVVnN3eJKoSWHYpq
FCo+tG5TVT6CmAumtOBkEfBasVwwjAYmb0mCNkk/tiaSyl8kJQ4XqphsKpqE
A3zfBt8dUm/cTTdsruJ5fjqmsxuz3dX6w3wYAhTXHHb9k3i/yrv9LAy6WuY1
Q6bJ5i+Sf72x8BJpcCyx7Gynm6IZg6M02BIhST1aPUTp8Yom4wUHAOs6kRAq
Q9yCVd6fsIf8B4RimmXBN7nuyDzNXPO18Lq8nxNsuP3kXdsDa7THR4p02jXP
ay1eU3c+S+oRwpnDJNGwGLFGlI+y6WsNylMWkYsEQBWOa3awaJiPWwgwr0Jf
64A5pv7/xd4ZK1q7zimWmq4PTEuVKyT+g9OVa+CfwB+NkL+dWyazgDFp6tDQ
GChddndemEGwlY29ALiV6LL6uCoPzIGx/z7QOr2diF2uyKd6f+6WFtoC9qfG
nObkcwX8ldVvUi+V08WldL1lXtPGQuCPCWkCik9/WfJ1XsmWvg9HBvrB71SX
l5sFnJf/9lIbEYOQLp8ErGxptVz0kHuL2iI2KuaPOSZKpziZjhxflhRgwMe9
rZagAdzd+X5gusWSG2Mmh5gOG2C70slbpCZTLy9H+VGd16FNTvbBStCAq0Dx
475SUhPZPOdtMMyx2PszB/5HtpH7OhNBsIZveQzfW+CBTz3lh51sONM3BduW
MIDwPNgahbDcUdB21S5L8X+tqruyqyFLTY2X6CH5WuSVrqlXtFcM8O098sKo
U7zT/r0ZJZbGBdrQawwnCf7juxZU1715/VT+/cecAXWMX/MKWVaQQxfuSYNy
gjdtOAUYImconewZZ0qG1x9kKr1oVmzeGYfi/vzvRV+g+Q5N+RPx5Ucygn8b
VP6pkW1wf24Ya8nPoQS9CGygkm43VM90hyqhBsig0V0PNWvpulf4gbr4hcA2
TLCBwc+86mLESx8waPgXiHDeVqbQQ/Ky/o7e9VBHxhp46BXFYIgXEZwAOGN5
TzWv2Dz9mETYkmWNepDYX0VwvFOti5x354HVk5HSHWbbgPU7O/aen4Plz11v
x3r196anFNiJ03c1Yjc6RZWt+PsQdFxuKJJrAqoDz971QhFiC7ILmOt13N8/
i7Ebq5ol/6olW61b6gqpzmnpuHwXwusc8HYzzdBSrFLbatcPCk9xp8OSJD8r
icB6tF092BYQbsP/li+bH9JtGWmX8w49rdOYWyccadNKpegWfjJ5uD7JSk4G
iU+u/aR0HLjfzFUbYDVznfdtsqlzV2j5vpQkKkxldzlLWNR7/mUW/EreLaRy
2JEL57cei5ttrxwZXwezrtunbOTNa0axG+7CGXcxtTsy1P1YnC3dgx2qnVt9
8GcqLGWRqrzluS/ULWLRN2p1tGpsr2NQoXZGK+lFWhPWcHqo3OGICLZLAp6i
Q4spA59r77cwG+7PUZcPzLYHtbWIXYsjXYS5LMhbZWHQcu+sBNBP9Jx284Jp
AxdjoUS+n8bIxR8Ue2m5CpZ7UV7L3zQjcvuLkgnUkjZzr6XHHCj2zLMg+aXr
DywKpsrkHjC2DhBClkDBBXT6MMcWiBK//Sgh1hR7yfIZoXzr1Bj3ZAojWo5P
FZkMFFuWOFJXoI7BNE3IRAu+qO+T/gF3Kgnyt1uFkCj62932sq+a6jExLEf5
Z1U8+D6n205oDpzRLUPoA9siG81x3nfDVunRLw98VwEslFMeyNpOFx8sL43d
cgA8Ngqq01vxz95SlYZJ9uNY9OIwe7Srp71JPYiRozTzhIPQFRE7koXLXt6s
23jFtliSJDu9sIvHJUKB+gOuEssO5/6UH4saYJVg6JY4S8YCRyb8NeSUStRZ
yrpycFb7tVucKdZghFf2VmrotEN1V8srJ5rjvsqu130g4j6YHKiZUO7E4Abx
IaYy26cxNj3YlloVmLIyTFwl56WOlizAYqtzVAjIGdVVPk4fjsi4V7UtwJjW
+brJwoCD5DPLJPRm5waKjYaiTJ5suoIAetSQ2567V2uMQrsY3oxqMzqMG5Ji
Y6sBgfeop0pKC1sMSNcQZZ+YO1QFwM9LSXU/qNnFXbqj2fj43pUX6tOM/nZT
Kt5hSC59NrjICHrINjjtBtClO0QHE/5nndF+VVDp8AsuMFx9jtHmeuQqGBa+
cBz2JlBUtyZdr+8LHXP1/IQVYDmifgEg87oqPDwW8rRliTk6D+vWfXHsGt9X
wzWpP5cd0p89sj5UhfQzSx+XDHCPrd7QO+7XYstlT14DM1p2vKZn8ui9DkXg
LN6mrtI6MNxrnEmk1UKH9R81uzADS152WZZM4WbmWnh3XYLIJMrpzrw8WlD7
Hm/yN8UQXHgT+XE+oVazZLoRK0Gw+P4Ke9b/C5+vZDoJRbRP1Ay0tOgj1Hri
RPblKX3VuxjmxV6rosMODA5JqlI1eBLRgONsveouHeNMZVN3TrEdXFM46SV8
tQ+a8oyXCfwksZogrONU966ZHUnC9M4J3nhepCBYtjm0d73XyLZ9QWBaC+2m
tVw76MA8SXQnQLJhze0AmKNWxpKWpR1ZimB/2BvukMd/9Qr1OaAdfTXvD7fD
KW6XJLyopRS7ZQLZ7OOQ3+V83SZ43NU2sVpx0yPUFAGx1TvKFTyfTS3oKZil
VWA3IAACPhF9eLWCQgqzgEWgUAR3QIVVAYhQN/2PRDTrL6WqV3vzy6MvjRds
g2JGUetgVSINRYmLcZL//yMyVFOQY+NGaI9nVdpmXvLCbcN7WoBfmxN2qvUm
GoRXmr4euNe8xI9O5rq3zjydXFVpdrTHzAqpXXlbocEhTO/EC5yuddKEnFIc
6XTPUru78eywT+iDkP7ac15Tuy4QJQJ5QQ+JR+Kyj9xIzU7l+/j5XTEztxmU
kz75l/dUzSf/lCnxkkdmhuE57qNjQ6gmn1DfIF0UcGGU7WG6EHEA2rcz1+Ak
A4hAVSMGV1M7ZX7GFwiLEGe3OzmA97uiqIvCte56nFHs9dkx4dkY6LCo8b8x
d2sY9XefNLChuYBqh3D/zS7fQ1ZLTRd661P9UJCCKdsxRz22DIFAAADi30WS
Ocpazx7f1j9eXoflHtneFv4eDBYs4AkARKmKrZ01DVpaPbd6UowbgSVINI6e
FRfY1zO/dPiPt0vYiin1Aqu5lyzSxltniD+f7RSPRJQWbC42tshNxSm4e7Mz
rlIW4gtkMq0ATOgIelhwtpqPJebD2quPA7dXpXxlEsx9fV7BWQFT/14EfCAG
To1n0/lM8wZcRSU0RCKD4BVc+G4sijhzV8WnCHyw6BfrSTe3tN1Q32D5jvpm
F1bM+wKLuAzWliYGmxFwnWnPK4meMYEfm3qYbx9aPt04q1VvHBwEBcXimE/B
dGjzTpEgJpCHGmkwCRw4zglpkA6u6Z7CAldoQp2CXleU7IGOEUzAm3CTGkAZ
5/dX3aHczOfH/Xa+DTFXP/9/ppuOioY4DFV1Xul0zKSV05KUeD6qMMHIMTQt
Jdmd6aVHChn+PgNzZfMk5bDatjGIkilbzjbIgzyHQfajU5n1XNUuRFOP60TV
au2SAnnPJQR/2SErzcR+2rA02xivjzssgSo1bF7bOq+plTAeOMcSyUN7Zask
ccy2omSZKAQ/oqp8uU5RJqnZz+CAidZ+7pQyuMvXnEWcMEnmVyjHfyVxh9gq
XsphTGd9q6lnnlb3EwRfkPGLx71Og8taKUfEvP0rPNems0iwPligTetHBz6r
jzclOluyR43ow53h9vBkc5ebSsnzU4SHE1jAJGo3fTbj4tTTu7Gn5JZbJHGJ
XSond2RwA9G7hj7HDCiNft4u2GKKbKBYgYACOdsdfnEoZyRSCvLYI/MOFEcz
k5YP7ZctgUUP1f+UJ/9+tBjLWXSZvnu15bWa4kyMrZ0szCC7RQNZ+jko5w9l
2NcbEuHQ3CcS++ENBfAT1ml1zz/MzmHhCKBVI/lh863ULiZPWF6D4idur9Rq
Oz2Lx8NpxC5Ac7pIum+T4lMEdMBIbJv3YxCTQJOV+VMU86WNqqGP6pUDnSVs
a3eErB6ay8KVT336ikjrGm87BTIZDk7vtJYW/XSQDwtoMpV7khDedR1C11WY
0gFQp6zee4ZmrDr9Yfp/VbvE48uikhY0zUN04nttD0f4PeS02hOUtoPOoPCB
lt6k13u7SlQXmIOI75ZP82o+ktW6WkKQRBF1mq/ZlMorZthEEz8UNAdP01Ic
JgaErTTWj+2vNerfOu6f5+uafFQjp5ZecWdlblZia/Lf33iq4N9OXKl1iOFF
mcqv4AiXS533dT5l1+UIdeCh3TQaKBMDtLbZrtDo6AlROfXjBa8/qcTLHCtc
5thZNYfIj1IMOnEQdimsnZkTcmCI0PBbBpoL2Q0PmI9IKjMLPTb35515qzE6
kXE+TY6vCXO8twI/qiyNH9NWeOV5ETcs5Ito2mOG46hMTC2xd7eSFoBNdqxi
7/9CVfpVm3SZYkPxn0U1vuw+OxcuqJM6T/uZ9/7XxiF8zFskJP7m+itAeHAN
555HjmBBAbrK1Bm3NhSVuUdRHZwzfZ1pzoFH7cFP64CPeJTtCUvwpTgy4I+6
ly/1LfxysfdvRM9kO38k9qOKia/b7h1IVYNMq9wOEaHw3D/06i9sCgk19DOm
qvPzPYt4zAKn9Z3v7gPKMpwmH+p/j2cjZ872sfGiNm3AHbbYO9BfzdyN1e6g
ggYwY6tKCbPhfq9ad9/BG89kBuFqnuEle2jUrGqAm0kbNSMLqaNYxoG8fxyZ
SO9mIf9+1IdyHF1o4dEHgOoNwMJJxPbxXMcTD7zdfbMX0K9+FxmbxKsDUlsE
LiyP/u1iP1uhO7e8Nu9X+ZVUryA26NfzoMtGVIvhJ0OuztZ0C1UChqzx+bOG
0K6UdAYm3H//q7jD1vrgZZe5J2M2AOs8wXYjU2z431ps9tO/Y5k9w1Exr/CE
vyPLIPEgdaIob6f+reRhOK2hlssTBOYKuqdMggFuUzuIIMeouFVRr12srwnt
9BrcE5FpZ04cP2uGEMAXSvsY1kjL2eTWou6soS6CaqVd504wQfCfMUgaJJxY
OecavBFma64kGgX4Z7KbeD5iC+mYUpr+NWY5L9pEw9hq/1wMSdsuFJNBiBkL
Cs1OuAt8tGzgVurTEZNZ3k0P6tT6UzqIzEftQrAiYQHQrw8aht9VhA43f94p
5XYQFNokLMlvjTT0q2Itm8YR5HCYs8Nl4jAcnZxpVqBkwj4Jd37xDe5WBJqT
egL6Jgx3EcQw7JTD8FS9cf/aJz+P+tJ+wCzoK++xP/txhGjpVJOyS9zGdSO4
XMzI/rth7xzqvelGQwbjwEKCkw7tVB+609wgRD40kaMQVcrzAvSBCcBaTJZ1
3NxqNasKLKwFvczPlUoZZfXtHvj9KHNwt41AKN9Ky0Vy9VSb6RefFTmKZehG
m3+CN9XgS+qMjCBXl7Dh+IjNSHRpj1y3SCLv0H7I0afTqE4X8+JW78SaNC/5
9A/4YLZZ4bK2+Blbt6ve6yJ8l4cCIrp4J3Rha81X7T3ClTOkJEysZMS0QSTr
Pls3W8QmDai2o6cKOoEw6ML6dWnWpSPdNd23CIke92KN4QhpPAthc2sRfdMo
0jBcxf+38E5mS1vADSvrg7sFY4Pzrq4pwgccOHdvxGH3aSNO7qBKGe3XQ59n
JbDnTmCVmf6R5AveIRDr+2P5VM31kP7s5qqR+FCWtBLMSAt720f1uIlnWgLd
tYgImOG95gMgRczlW6cTlv6+ET+BWjZ5ShClc2PAOWCtAP20qDM9uPttxqMz
AmD7JoLvcvQMQT+pC5Uq+d4kBDmF+TfD0iNqe8ldMXEB8RQ0UIyGXcGR2ul7
L1dzQmlboAsxK4zjAw8CeEY3J31BeBKoK4bSJqdPZb8jL+PBPP2kH0lPxf74
9+T2FNMrfzcDJ8lze1Z+FTaeOf5GfFIL/hLUpecOq61dsH27XL0FElGSKb8h
TIFn/j8oPgkijtGIcYkEAVGAkCb24a3eI5y/rYB9nosefdEoNB5eKeoCG1GH
sNsKidRvTuOyfFm9Jonmk2f1Cr9q/AdB+KJR5BuWRjTuACXyf3uDwPmsgjIc
CHyACOADu9s9EiRy5ucbt8fIKUxpVFgCLP6c0cd/C0rF7mMyL/IzdXQmflKr
kuGfY5cO/IU7PFupUKiAI1l7azPFfWBLkq3SHA6BDbgTNm+g0wDBGms5XVS3
M9cnMPIx6yWfOnd4f+1AhN1QtcSTXAZWB8bivd6y9tTuQ5qqt/BxoSZtbAk8
+v2qNvTMWiMLu0cWIBEqyLaO2+pULzRR7kQyyWUhlno9RND/Ewy3v5DI/hXA
UGFHFmd1u1fODMBvAAM08JqMoK9xUtxJEGvBkMONZwbl6l76WD/n6l2Ra8c/
/jvmKR74+5A130mNoRKQgX+J2tFHfb2Wa1JFQnlKEGm1Bax1eIbQVH1U0OKt
SJn0KgW2aQ5DQV7q0TQsP4bYzl2Hk37sg3zi8/bJ8x2kQsJ9FcNKdZ4ZWN9p
Hju9NMy2uYWmpAtzBBDVekjaibOfGwbb2vy9a0xuAFAhT4sgNSdamWm6A3GI
Af6HY094BWGIKzOpIGGnzeo1rOR37lZk1x3U4UN2zmngo+GwNgNUFgafsQn8
KnEWRKpQv9pbLlz4HPeTFvDnQPUyUDvCxZA4BK2gt/Q4g0o32VzjINZlwfyY
DQBNbGN13OsvYjS61fLOC2W+JxeDeuWCTJka+xy377O4oEvFe+CWlW3ZF2FA
3SiFcpWC8NrSa7GLvzxslKQlAqn8JB74oBKeKNlW6xizAiAgK2Ddxyt5ixdP
RaYUE4hWoalkatVYKyYE25KHJVK+vgnMj0QUvtlcnC6bCVwcjz3bRniC4imP
XXag9Smgiyq3wBA8tsx8yBYha5pIJoyEk7R2xkJalQTxkTUaycb+wA52gIhJ
fdVL/jyIDsomfyXRdWEK1I5TCPCKvn5WTu2xdv9csbtk+TSUMU7T1mUOBkL5
Yp2ZQKXf0laf/a3pWdd7gUQ+Y2G92OhzsCVH6A0XA4nRQq3MefjKIuNP/7FF
h0WBXMZMXVAXXrGt01CfAwKqVue+pL7m9b0xbwxth25j4leJOs+cv5T+Dd+q
kXvQ7KZROT/YBxgwNRcQc2X5EtOclWKd7Gg3ZYx/0ruHI0jjy9rg/TrmaQaD
xxsRKVaWl/ENuRKWYzYZ0FQ6sUwcu2uFTJtaZCw+mhBkprbLiqFsDF83qq9K
facs0tmNnjw1WgAAnBbvKT8zVeskse5EWv1lhDkjbWbWtlNbSmKIjVwQiQBO
fL7DuqdDZIrIlH9uOuEscWmSloN+9IR4dMiFmJNUlOt9In1xgyJyrro/iYdG
VAq1Z4nNb38bimfupbbSy6wvy6o9zJM9bIAZALUbKdGmbAv0FD4wLRuwmVpb
W3MgTRWz+gfzf49HeEBX/wvAet5qOhZ2d9QlqbgVlUjwxgxlZ78bDAdW/gir
4iXOVVBt/Ytq2Qcsd30bCIGo13aQ3UQBNY3nEX1DysHiBce41bgc4mwsXdS7
wTbgA2MwzshhOK67fCzq5F5hvbQ2EAPQSrJe1JTmk/ILMel4pjgQ95PTACBs
5MsIhe6c3LjrvNHVlahVlS1OTcX0posp8PUyUMZDPxvpp/eQJv3WT+LB3A0G
+5SVmBEu0HJ/bA7G+UP19RY423Ngu+IKq0G8ToL2mAXyYBtHfeqkIvxqu1sc
/MYwEXfC3xQMb7xHrqPsFdrf/RLWsyFdLc3R90tMcwHVijkSEkfle509J8JO
82OcGYZO6wDWJ0/yx3pBVJGzXIHSyqdSolnmrH5Y0d760Ln71f09CycUZc6f
7tX6i2rDJJVH4rFk4DfwtQxf4PARwr4Gt34+ax6sUCPDLrRHhPVk9toeyIa9
14HEZv+G9mpIBCPw9WasUIpkiO9zeqtvhXWEVaqhx0Lc+W6sl1kXYnlcxK1H
8BdT7hdeGX6oUf8YOU65XGjqcJUBza4ypxeLntszpbOriepyMJU1rz8hl6ut
KpwRMluoGb3FGKxCPngUXEakB/qojLYp2F+Dw6ZBVqFJKa2VUC0K687Qw5jV
tnJUR05sOIpf7dAtVppIItf0rAiGcLlQe22PxSb+HzgdgONHWxeBGFWez3R4
hmYtGGEJn08OhBXzPZYQEbZ3kgpIDiihS0zri+Pb2YKCDjeXCxqfs4h46E7+
gt51BWg16CJAqfAodAGM4xsR3W6n7E2J9ZElorGPkUOVSvYTrHENh5XwJIaF
f/fyyujZy9pjpiDsEdoPZs4RGJXTnXbzKqmE1S1pNT6hmPQyFldXYzQQCClW
jI8HuKbg49TirGQv1hOtsif6dbvgKj9+ZVxoqbK6iOEW6+s2PMbVgOK8nOA9
YZrPFMESNrlRKvg5OGA+v6MvqgbocsE/2enS9emxJ4hYIsbXleITrLgMjf2B
0UbA7X7P+pEhJ8ueAsaoxzhgKh/VChqvCwUvHIvLpq85JsQ6UNEydU9dQBlJ
yJlIOiaQpJDrw4p/OXHi/bmY1SpdxC2gpjjix+7Tvef89efjqWE6CZ42tbLa
ANxVaTcQfoopFmJVbKKnrcSN514sF/1gFyPBxbG08U8KT2awgOezFW0t8Tn/
PVjvdeuAehepwGK6tvDK+baIxQJi6q99T1jYJj6j3Yecze42yLg8lIvNFLyF
aPdmZsX2eeTpzbLheuAjNWdskGA0eoCtw7VY8LK7ekdWBvNkBz6xWbHaROsL
0j2bAC2JzN8OVD8+eZWQ8fkXdwDMHOM4SyoasEOIT+ojB41CWw6gV/mN2eVu
uEDU0JnmhrinzE+qVSQgbvngOXp6VbM477+eYaXLattjxTU+5SY+iskUm2h4
b/g9ZLxw7dpl8QEV1KhP62Ty8zr3Gdtyq/Z9WkkrybhY0IqF03ztXCtMUkcy
4Nw4coz3zwx26+rAYFh4nr6YhNtJOXriu4VND46SpONkMffHyV7p+aGpwAMv
qximZO0C2Anj2SJJzqp7PjiF7RjHYuTikKsJNb+XqQuU69wV5h7cSHpUBTpx
nnyTpE7UlLRBAVBW9XBn4BKgMwyPI/PEh5YAkqS7aOZS8cmLaYcmfrpguSZ2
RVcKBgm/ygP6YO1FvvW5wfD1tGboAZcAbEnAh9EJDkq1teCcQ8zV2jBwLZZ3
vX76meLm7LXDSBNMkCypPY48r6ZTojiB5h1HQWuMdPQdszMXmnXqLpwh620T
ze4LUPIengbV6y8XE3smcNERjWdOuZ5HU2rarqtPevdGsrwVAKRcZisvi3uu
0ACrriIVtDV7qKLdCBj0PZGWbn/kNt912HHHvmNik4TjP64+QWWMfxWK5cvB
Iw5cSBsjsKiPpLhU4l5AeKEILCd++jyAtC0lBp60mcZu1CSmvt/tkqDdFjF7
tiK/sy0cDSXEdRlCptq6e5PGlJYCJ3SGtrMIUTit2ekoUePjb6NCsZbPzGIc
JHK348js60LkziBCi9bez0dE8Y6M1gd5pAQ/dYq0wT7VxER6kjDacs3lsCkV
m4ky2ePNOZvQZKxLN8diJYtTY/1iLYeqLY2dFyY8MpJCti/58nd9DZz92i+l
GRolm30OrK00wSsGGOFJqv78lOHvXks5bBDy0dzA8xMqanXK83WxcwWzG/Ks
2zfsxvozi+Z23LhBMi4U8LC2nsFs+z4I6gYW/0RP0M9zXRiBxr2I/3jTmkGd
yjYLSMJjZv9oaQ7aZKr6auCWg2IA88rIWm9oA0FHtWsq9s2v8aAyTy+0WklR
dRTs86pgqcKdkFE9LAB+bwcc/dKCaCQ5bOOqLZF/d4vkd+yDoF6Mr/SyK2B8
Yh19ySFx5GmaGm4s7VszBdY/eT9luWnA67OR+Hdxb5FyxFn/L6MwuTowwBH/
wcB4SB33e7QkUBqnQ52CykqiC19MFla76oxEmARw73mbiigzHOioswgMehG0
5v1pZZp6VostYptoemn3PPTWsyzhlqBLqIxW95ObZi+TrXxAQJRrlZ9QndKP
aUugyX3dU9wrqdc6f9DmVvJkYJvqBYbUJmspF9IA51E7HNWTIje3v4EClnDA
SJr+ziryC9j4lVnU0iImgjr2S+LNB2kdOc3QjkdbEPx7TbwO6ZDNrDRcAxrr
zhlLp3OAY9bP4zDMNdhjTXeXmjiAVUQHb7zbb7WxRCWlPetEEmZG9L9G9Wfv
MZrpDakV9DN7KHOc9cra5OWaNrQMNjAQzH9K8pnhyWUms3rdzosGRzpFTT2Q
p3OKeQl4Cq03xLsL0o8fNG8+T6CDoSCm252K3sdXZb8XHJye+wyC6VbCNY1U
8V8RseyZAjbLKE3LXS3/Q6Mwy6U18hLa+BjH+9fwdI4V1OSUBB4lWHHQqjjz
WZNeDGPxKHmeGotvcqRPvbzREFygYHuVPFnFSdiVCJO22NHWnhMNtAJZwUsi
qiA5aW+l/wPw4rzYr0KjfWGzP+B9hctkneifBDIMyzwZMIo5TiyUR9vmKNUU
fngT/CyEUE33dBA62NjddToHcJv5/OaQ0xkleNnNu/ijTOVelXlMGyl8mVwI
64H8qyue4jHbxSQXumSaB08Czvqxnzd1feMOazGHquPPmzPFKL2EcVcdQ1+U
n5ePVayuCtIBJ03WR8aHh6iE8q0hCkA6lhdSfsyhfjqmDVYBZGFqz4jGGtDt
bxWTfIO/o1UUfVyE//cKVgI42s1Rhha0qYN5KUIl6HpMopf1Ez6Wv+NEQt7N
DHCKtPoFqbKkIOcYp6eaI9C7oJlPU+AMJCphf9ItC89VrSIpWFpUWJE487aY
nJ1nRH9OqqZq6ygtKDLXkariuSxS0XnbDchdHxJuQueBl9lbmuW2aFGUwz29
J5dMTqCs10F52VVsTAZKmRDZIknSPOjb5S2N4z+gzC//t3F7WjLiVAVgfVyo
atUQ+WpDP6ymRaOwTGsO1EuAd//uk7JPhhAmQuOGC0xUiYdg/IyFNmNjFYB5
if6pJBL4YgKrYz1n2+sLEAe8TjbBOuoLYFrTpOnpjNONwnhVjtOHIMu+kglQ
RhlY8OXu6OMgyb5Wo2TfDBNJHgkMzcXRZlphulI7sawjhUnkyQX1fMjQFhu8
P69NJBb34WUbI814qSZvyn9G34x1boLtCNAROmwwPdCMaYmRzyV53jzI8+Zk
Sv7CQLcqbb1reFGAclRXS3pfN8LE4cdJFDksOgNG0iK24In1BlvlBWmiCsim
upgs1Mb5ogrGmbRfSguT2mhLAgDTdm64sZYe8dqU6wfNW6fg6yrICnHOlVVv
gPo+Ro8gvHVhTKOobR40TVA/rnwuHZHyRfM2qZjQdGEdze5KgxJw24E172C9
U85Cz3HONDo7xuLHHL9PmrjaQ1VKBtZqWGK3UkaHWNsRMM+JS80DFlzfXl6p
h8aFicvChILTmLdSUF3Bi/iIVz43vpfBtLTxpG9Xcr7pJ/2M4auP17Qtv7wl
Njt6gmKl9943Q+b6O5JTRXbJAe+VVVsM6WtJtiQ+m9ZmQIqSm2wmUVZ1ncFZ
Nun7dnD7DBsAqq719zaHnJfdVosrnsXiUNYdtJIcyf77TgLsFDJJCCFZgoMf
F3brQitq30wR7wmE/3s8qqdPmJvcmKOP5g9zsZyyfXd/g6O5zFgzKq1IIjiQ
fs+gxgutea7R1rvgpwDAGivXhwGACW8IMxhcPgRrPNRIIcN+0LmUNaEutHlH
CPogqBPahM0OOlkT3r7Z5mgUPrIc/vht1tUfJeDeJ0CTJNhpHEPKDhxwADtg
6au1vE2yFSh0o044PAKt/7v1olP3R4XLGkH7ldpwIiGiM2q/w844ZeAFrRAk
dgR6ejk1B31xauxguyk2xqVwpf1eOmQZpJ7WacOawfZNnX+cDHq/U4diluWZ
7LJsGhWhAxyy7ZgFmsM/wTdiGbEer0FS9ORMyAYB+pO7cB8UssKW6x1k6HqG
U9B2zg3UmSDoa1jnMgnb4PS1jeMuXVRybW3g5TnovNS37s1KIOl4KLb5W+0x
uSzK/rNNAH2NborE+bF8OngkhYJU2SXj5+/2jCvJcPwBNTrasP6A2oaWZFDJ
p1Rpra0XDYntqh8oZfgTrab1ACMu1o7nxTndVVjKCQkOzorVmDBwzDaL4pAl
Ad3rwzy1VGtpADN2wIRBdgMnkWNQ3VtIWWANOlPXYo13stBN/w7XrqxzWGZg
QjjpvG+54He+jdLVi1WgDQd2JVRyVdWFn7xw+tF8vpod4I/AEqq+XMg65dST
Y7wrXISKyYwRxdh0p0ApJKMYTywk1xG5Q6WfUn1/8CIg7ME2D4vrtuoJHxfF
UlwAS+UJ5uSpBBcfhCNE1Hi/pUpRpRgU2dxiroCeNhG6+bKt34NkorN/+GZG
0wTpKgZ/yzcHu5DhugoRoShuv7mnb4Yn0CUw3ibtF5hxRrGzHNIB0gNNPXgx
OGVX498bZSijSv2PYiiX/B/G9Ko+jBRQwocUEYISr3UsR2DiAKjp67zLaDhB
0vi3Roq8GULVUtxJszjrDiF9qAbTscUR8Lmi2LzkSILgOgMjSPL3BelF2cWe
Bb47H9TpSlYstpHzJOXLdetIc5+PS8ezl/bIsz/OLhbnVvQfwtU7nXHPnJb6
GX8w4w2gaWbOhnsctow1ThWNA9ggl9ADxsfUJwCTgfx+7ce8oYJMOSClOLdP
MJVI4X3vQMgrqOCvjnuR2wn2Bzc34PXwkfDAeFJeu4YcKLb3h27UNh5nzqO7
neogSSzvlSqyiUZBhP+J7reXvsvZv0qz2GW2I7WxbI6UPM7L03ixa4qCx3mD
LJk+XAVl5hMj8LX5gR7V5+zTSTK4PBQF75SQ7R+t6K/IR8v+vsXKbmExw9W3
cLp79t82DEGUJQdcO7vgUo3GOStUOD2Tnpq8FBz/W2W3KVhCl3avfuX/70bv
WjAmxA+SZ9LvUaWg+YixY0/lUPq9HLT8ciGZJuahjuxTNcfNs0s8tb+BtANV
8xQ+Ce8UNCTiIBCqkzYaiajI4EqLIV3SSlWhSUDGbypoviJtpiAw5ffbVsqs
UIicPMTSqCrcYpzbVSf4LaEbXm6sx4M/C99AYC389i5fhrnO3pTd4sTig5N5
gA8O6+glztW5nwjayJivX9EscitdDgE9ZPsO/KyFWAO/xgR0OBZqSsAO9JcA
FCDBOCdlvanpBSg4En4oHSFMP8RklyaX3PIjublKcBfS8vjGoy/FAgAatjlX
ndIRzjHul+0F5A1JqdEotAwVkXP94fQcsBOd0Xjn77HL/td4wkyPCzxPCG8/
Nc8dh42f13FNiYgIz5u5+u4NiN4wU0aMuTAKmm/I7oLyxYw7t9PhilmdB8YI
04OvZQwPrvMXG7jkpibgZCL0zSl6iu4APqjvSkbEQSS+RydJ8MkYiAWRugMu
KA/WhAYY+rdm3pWva6Dpi46i22EoajvnSewlemlu7bPtezQVvpFrikdnIgqZ
do7nBkcnEWUlWHlU2AdWOLLsp+2jBHWuFoLKSouURhEna04rrEhJZWiNf34+
qiySN2Lzono+xpkNHNZ9M6l0dQAUbaIwpyeSX+hQTYFKrdwZh5iRcqFArBBG
nqRb2BIjcxaefgqXEQzLh/8C+cXyuJaPODWbc57LFRTmr7IYvlTfkYqMAWAi
4eLM8gx59r5wTjkcFx/2F/ZoF71VR1LI28vTQP7C3WXI5S3ekMJnWj6Ep12b
PsEPi/kgpAv3ATuEaMoe8wABkhyuQr8vYcGXEP3AXyg3Itc7iEkXP6xmN314
TSHJQnkF7ohsVwXbZ/GDiKSSrcEnzZGnSMhKBP0QoWap+8qag4S9qz5fPFJr
F1Kk8ts/y4LiVXmGp7txdWdeRFlPlTuUHdpCqpurBtQ9zX7hx4qBYpzDkRDt
332olP/zeLy4RPINaorOQL9qUplTrVRUFUghgmgEAyCZKDMvboQt5gifhs0m
5iqCQMpsJzhobhbBXTv1pDBXrnIj+AlWxP8DzpsdIWSqC//PxdzfZlKQTMLw
LtPgwnDe+H1ASduHqfFUgTu7TsXPFQOHnkXwglcaOW8g2efVS8ul5w9Ldtcy
YQUHc8l14sgnlLSbU7NtmpjWaa7Bw+b/0fNIx/OCzI8M02wjbykRNiRt7UsG
Oyc7Dd4uVRRgUrILIEA74W511O8r2SmatYfOy9SOzYRjFBSHokdAswX0cFym
hBP8siPO6MZ14fy5h1v1rTCk9MbrNSRo/sHjbObokStBnb88VYXocl8m8Q/c
b54MhY6P4TARmKBDJzAHNndljaIKPyWWZoC6XwW9234tci4KWnot1eC7bcKw
KtkDV3oZrxl4IHsLJd88Gr2wf8Ja9mEaHaXp9Jbp9fBNtVRRCzH6MuvjtzbW
yzdYtJXADC49TY3iSUo49DX0/gEeIQSO+Ozesv9xWf9yiczrVHGvpt7jyy3k
6j/sxDEy/RoZvX7AazhlQMTMp6G8UIWG7E5J0yX4gS3DSAmUGckVIwLnQdRa
nfDHG/H4RDkG64gfZDBD4cA/D8Xgt2w1JZ7rp34zk/FD9QMZ3JEHLrpejYxQ
cOu5zpSSVHvYE81ExfSSq2xC7etH6WkXLtb6re94IdchEvg2ieRUl3z0wQeb
0fyflvnJLLhVVEzXW//sCrMOWY67O3qpzmDYbtzWW7sugO+L59VGNf1cp22C
ygLOBH2mRVdZsBgMBGim0sm8ZhWaluEkkbNnqxIEWrRyHTVlUwil+31sNCoy
pGynuRgMOPwbQPS7JLrS78QhJJxQFXt+M7K4pQ7SqyuDpAfspp8ahhcTcHlr
mybh4BaUkE+QTSzRXreLd37FdFp4eyP9KjW1Zjv4XNP41T8HXU4z9HhCmfni
O1b7yllttnVYjNWQNP2FzUOG/tsVwkgI8QviZLQPrp5tTPQxTCaDu1MvO98O
QOjksM3WEIfPuutjjet8yCxxMjsuQr1zpRSHGH5jb+NLnhQa/+LpL1Cqqsuj
lwU07dr3e03NQaDEz1Oxzh4pofcfMuf0U25IMsAnlWRyhIgf3rZmV5GOY0Qp
cBcO1y52YAd6aEPnvwLXUfuCE2ZA2iM9//c0pCuntow0SlE4ZID3EcU8O1Je
ibal/FzvQZKq4AHNMtwH0lFp2Ns0ERbpoPtvutDW0wJaVFHOvFFUex0a7j0w
8UC8DPx/Bu6c6CHIg+HXFY6R1H/4x2HqaN4+cCmRHomIzPDcDQc7VObnds8n
u6UWKjBj5AokqC63gfU4SQpAMn65Bog5x9L303FANmb4AKGg4cja3SKv8kPE
I5zjwTEX3Jpzpnroh8mOx+FqSpk3FxtKOgVf4nEe41m8Hca2FYDzYrij4PyI
V4LzZAUe/pv1eI+TtozHvkVQiQTW81vl4MwOzwVVq3Untgxsgo9qimHwYZ7o
5L+7UqteMc0eJ7fJUtbqhyTJhzLVK9mSBEMvAK+h3lZ4fPUdgtCWg1iUOizK
lPpu95d182VzhsZ1Uv4LxoBFMALgi+ApbHv9AoTq3Rn0q7s2D7jUOXhGjpXJ
sJ2aCW8okfoW9RKgkfnWff2Jhbk77DE8rAzPY5aUf3IjksFBhO0wVYflw/cT
YsY+7zJXdjDec4stFQuhUp7stKIUqFesxM6MQYaA0GSmlE5IE5eI4T9Bmdx2
OrVKfAXbwgSDH6gkQiYynxLDmKMLiuhxCZdX3sYZBNLJhMijNrh670kxvuAc
55v400k/V25tlxFe8YpDPKLx5H22slCwoJeuamn7GBJcf2Tjdi3mzY+ITQfu
CLJNvPxEyYs02b/hjqQEr9FrDr43KRE71BR7sr4b5sgusnQVfDjg8LuRfdn+
5r/kIS2PNG04DNcRIZtp/MBmQaFS2oriGn3qghQWapONCvKEPv5Ai6botnoH
c3Zvp0x1NvKVVubgkfgCKyTSP5k19tzPiyDtJfBFYSEuEHRbM1k2zfMF6AX2
Iqm4FHkuckm90OTTFTYMcZ3n1nZUea3kEFwEFgSTkc+gsP94jegx2BdH+BU6
1tgDATCYY2ruGJmxo/aW6zsQDdNnac2vopbtm0Xlx9n6bfhWO7fZ3qYwF1JM
5IqhXtCqdpe84ltE2ADzkFdx5v9XG+P0EqNiGpxhls5Ppo/IHfISOjcocruO
wsl7lNJ9LJteY1B0VPdJvGlgtkuLi4y9cyVBCn03yFYwvDaS+Rdx4xRavleC
2KxeXVcmKE0yl1YLLEs3AtfaweGiBL5f9zyCbJi4nab1ULF97s84vDZ0xciY
lRyQCSFkQEeH/mglDX3V5Fa63PkB3iueAUjeiALzapKJkyPMCFc+nziLA5OV
lt5apRQB6mLeT4ZH21Q5LcO+N5+z0xiqBxS1eSPT5Jea4uE9Tc5ldZi0G5Y7
KHgdJWNn7UYL4bJvFJYI78uYs0K8l7m6ptqpD2dUkzK7LXTpP7qT4KKh4HM+
hPQjjUPpOH+GpUkRvnygqMION5Y8TiKOfWF5z8j/XHFqvymS4p+UIzbSwSLJ
JduPB9ENYE3hNDPuPPcdL8n7AQ40gQsMWbXvx/EwwT9+jL8hMoGHAM484bt/
CK52XjTbGzR+Y6Z9Q0N3GqRoXNo8uUDnd5cczApUYOzcYbcui4hXOTltyFhl
9d7t31GLjWJxluVbge480SbcLbjdLTAE51GdRSjTAvZcE6Yd2IAhPz2Hgbzz
NuCyY2iWlpMNup3frpV45vbRzCuYkHPqXQwng2UwRIVUUBPKdfb4Y756svqM
gqXx1qF27GOrXzbA/eIkElmQLAuls9XvUcuODafnueFw4QCTmCjiiVEy500m
7ru7t5Jc2QBE6dSKLr4I38glJpz2HJr6Nku2qPcCFDLe5jhWSs65UOArkihx
Jus6azQOM/4DWos/NyYJ1ur0hZtgfze5OA66oW0f/dzfv7yPNKeVWZQbBGgg
LKboIUZWFo2YzfFB9DfYeGuMwszHQF2/LPZ1Rt447+ApGsi3HyDEA+ta6RYz
MlUDBOp0ycr0nr84drIg4RCQdBetm0MFcFMypc5So87JBKrS3wBOLPRJqQT9
2Rf9Z7l6mwvqcSdmGRQk6QBwj2nljuWefjCrInJFYqQS2+QDvaVH5rKzEpvd
WTFpQmHNDDExETVhlDyNLdzUfqtZFifS7ZcVPtZ4XafwoC+0a8eXrGR9LWJb
QNaFJHQke/rTfsSHAD9k+lqxfu+nMbhQ7ZB2Hn4rRj6aZ1BO/XiBo0bVoF/D
8aGEPOb3T2h1LNmW/6++hNPoS6BiNslDqfNsfvgRzBOHOEvgNxOrU43+fFcd
pi579+rjN3ysltVloP8lb04OTGbAPhL62sA0X+y7AjjSL+0HTrpHjVoPxdgx
Um38xLVd6wgzJi/3mNYGZLq6Icgfjou9XrZclC8f5PAJXeSwPbMqUvX3Ztpn
AmgKZHr3KFC1PQrGD8TkvpM1GzDyR/TMY/e5i20LN6fMnN+NYREWRWZ+CA5E
3RB+2n+MUOiGoLPfuk9oF6uKEJkLR7xitMfdCUX+v718IWaIP6Ry0VPnP50j
UgQ38EP2w9Ajcjmo98Dj8Kalqe6JpCfG5jnYzp8M+LmlS+rsR0TUIG9kOoDu
Bj48poX6EDHMXHq7KjRGbWFPNHfgtlPljLFKGO0Fn/5A5sxiDZTisg96ja+w
xbFwjL5PXC+PMdb0TZG599wIx47Ri/JasXqBrd2A2KzcRB6qtcZ8//ELRr6H
qslQBqqRghUYjGvdnmeRoUf08xGsQWdillazd9dxZZy3Qyy2TwhtwihG+/v5
6wMGG8mS8tvXnCGrFPLF2NUhGa8O42wqy8BOV/IKv+dSzSjFz2o/azbZp8Ty
2jN2ikJcpYr9hu8+RClYpbm8vriB+Mj6xf+zlCGXWx4atwEke15Vy1JpsFBj
TV/rcj+4d+imIkoB65zREYYuYYfFEFoFPAC1wZB1chjocE41dxSLSSST/s5f
AAoVquCPHu527PeKQxsf3SM4LTDRKWPrbK1yqTd9PLwBILhz8O/oClpWFI74
BCAmO4s/VeSCtAQeY8xz14Zl8thmcBNQWWdf+vPZbZB3L9221hrNxcGUdzVC
QiDWY9phYQpLwQN4UtHJmfeitsdZqBYB5ROQum7bIQreuSQSlCHyTrhcMFlG
2sDJgNVGfzSx0VZicTnsV4jUUcBbiSSETMfZjHuabpHhG6c/2xkrMFjdffvj
CoMbtuPKi+d1XJgnLc6rIVWhUUe/ISVOCLtKMWmlnM4CmP/tjOARQoB2wD6q
ZYChFBWe7oqq3aLVT4Yhki7aCzDEr6hTRiRHlHqFfhLrIVogD/acmdm3yb5X
HVidSMu16xe8QmolbEFCiilbTi9YdWGsKVC3NIt2e/krpAGATdODEhD4Kg2e
/nVcjIISWOw/CkA3Crwpa6obIR5TE7ytGRwwH5rKL7vgkEVreTkJmUogZdo4
uX+K2hYFujdlM/OlJ/Kb2mikapUbT0UjQmJhMuh4KjKT1fKsSrcFD3We12vr
wa1tDJ+E98prXaXs03nhqTAsRNVNP+QrZ6+6vZfxQBnXQyUo5vtROXyAU9zh
CrL+IwJ6c047kU1ngxknhOUiVBs4F+XKedMRdXhj//T7OawrdsuIrGrj/m0+
y+Eloe+jkomESy0fUVM1YZBlLhPVOU3jKTUIUI1odHAHpYOKCVRQZvM24+UN
qP7elivgpeSGZNIPjx447/5sav3OtBIuQhJZiTe5qAa/em3TMyL15CSselaM
1YEMWwXmaULXZpOX1spITuon4MX6+w1t96as8jvjXYTNE4Z2d88n+d64L1J1
Ln7ysrDTMDX7Z1hEU7ZR5cZH8IDjsqpPB7WH4Vd5GTIlSnWa1UuSemklhkJN
B+tqgBDaEdH9ma3B1j9Ox2DRKqrR8ZXCgscMiwyzpaH0bBCSSrOSenMOs4S2
d6b4c1CGEhvJcDNxHaYrty3rfwf2xEJN2O4+MmxMIht51hfpQWnfSlRQTo9G
pbOzm0qO1fUlx31B+jhRCfknUfJ1BXMSecjP5rg3zkW4tse8h2WBDPGraCTu
wdG/lt9UlKX46wN87IN/EcsI7jtJ1nj3L/tIsq4IrhpHZdd2QxrZV+ikr+VJ
5edl+IthhxuDvRpzQr5s1gpxd8/hCe2G+4Gx1orASxVC4EhUoRsGv57BwvsT
dw9pgRsIO4TzD+r3nOhdiok4tyS+0ghJx0261cyPjj8fG44Qzs/h/EUg3XQr
bxtb0UQ3awsdgctfQz8RcROWN9Zk4OGGJjhnhSsFCixOk5/pIAwYPb9qcl0R
EITHk+QG43pL7V/doBB+BS3EiovZPyxFVwwCBnuWwDioZr6JW73PV6+dWPB4
Bu9pXyYydit85SEDgbXjw+HQNPygkg38IlamfjaDcoA7TQIftSPcAx4D54Mi
7biJWumUvyOLySzwDe/3RH6gdudxDdp0fuXQ1Ff4qWDxIdCDx/8+Vsk/z4rC
eovUUkmCqNvpUjtaRara2jh2hKpaABBcymwDtvKBRJG+EG2Gy8kfqM341AOa
sCnQNOCOVmE6pGZqutbxXbDmNpQF+rVUmqFNx2P0wISHzj/6aG+GQsbF/GHd
rXQffDKY17aU1+1MO8QvcCn97rh+qloVx7gGQld3Oup7jVE01qhIYmQCGRHN
XNA5m60JUS8UpztiIuGSHx0t1LwdTVKDdVrZZKE5ShBm+DAQGCSTa4l0n9Qf
VPnpcOhUCnpVX2+gN2RkHqfUiKHSmSqrTFu1kM9SBD5IwSS1YdwHHJ4VvdPw
rjMMM3BFp8nFcn3M/aR7PFGo7+2gQ6EEz03IvTNQx0ZpUENVuCsIkrFd2yWJ
3cnSl5w4jKD1dVm5dJA1ZjcOaSJfyhCMrSvACBYVCCrD7+2bg/f7w1DXn3Gn
/152ZOM43kcTMwNgTZdpf04tNLmYTfMKZfmw1Jn5f2hgiB55XIlXOCIggzsn
C4QikQmnotp+IdyvEYxBaO/wnYLn8cIHlxDWeRyTgQKWVt1KsCVoFDC/MPyg
uBHapL55t+WLfPJCjSwFYMP4i1aZZn2HGnNG9cRbif574Bu9661PznZEIG0r
Gaa2BegOgP/RL1VC/t9NNZgY1uazeYPc5u+or0tIffayYbov4sAVIXJWFGp4
vIYRQe1A4Qi6mWZ63phLgCkBxPr5C2fbU6w2MHv2YrlPuWFo32rLckrTJD5Z
c9bud96/ls9dDBKiOxlYwSCT4hQXIO0zByjf5VIzEUfckOC8OcVXVzK/l7my
Fg/vR/+fG126q2ucoqMzXHzXVvga5jYOt2WwIDWTWvbnrJ6Bsr1s4esuh8wW
LDhMWJ/3vPFpdU3hC4f4sRt5IJHrfFBy1+Bwxyio8EmrJ4oI945l3wLfbM9F
KciaMFRjQ2eRA0BrMTK0G6YiIQU2hNb+pE6lpz75Lr9prxmasgdfLEAYYRza
ZH/LV6Q7oMgVrkt6FYSHoXQbIXgNeZaHLIx/NOVM35cB40FopY1WoJZR0emL
IKwYxKJTab6whmZ1VU8sIBhdv1aa/7y6Un+sdN2tbYzb2Np5tzl1DyENKAFx
+GebgmXXkbHE/IMYVZpwgZqlBrMWfLVWa6CqDQt0RlaszRhb4VZV5i1ymqF9
sZ8Ao3UJd92gM9SEHqfDpL+4wxlyVtAc93FhjxlmJ+NVqV0+zJ485Vm3lVu/
qkA5VtxvH64ptj1pEDlDLD5QNA5lQAvBbwDL5eaNnv1dU9mfU33clsosUNE2
SzjvxloTV2CrcGHyh+Xut2H3TokzLzYjBVM8fL1YYZdkvweEqkIVh+DmDAgU
s+PSaXtFXESjaMusneq5xkzQMBYcGVQ5sbQDneCXicCFBi/voM1/fZNydeIg
dNLCKjMRr8yaYEItgqj/PxSu1pQneKa9IJ8FHWStsFYjrK4ccIftUKVX7i9t
fKgRFeIx3EWNduYEbfxso51kWgLFovV1muXljuZ61Az/48S4U1rkpMCpiIvk
iPbTV7GrhJcLYiVryDWBKPDZlDBkuH9vtSBUUBTijc6Ct5nAE2WP2cMgDrzc
f4qhmCt+aw7RqT+gH/gXsuT9285635vDM7HCO5zJU9STbvOZ8qwpxGkgejwR
bj5DhXyyIY1KON7RB34GpzQq7CyR4cPzHEGH+5255vpa4b5EP8xmfeZA23Iz
CY3dGz+1L9ASrKqE4Ez323viSnYwhmMNO2PKQV3eUzYcVCpvGfSkVnlT79GI
WBwj9OdijY79JrDmEJEysFRkW4DAXNvwV8ezVHq8/IAUUcKAf6xqPDmM0o+U
zC1r+lGXIMi5zu+9PravEZAgFJz5OUMS9eqjXDst8l7isVbdGkSisBzocmZW
4KnTZqDhQDsDiWsBg3fUyDyrk0uKLHzQEmvXOzFiOMT4KqLGFDXwOVHpcZMg
9vSi8VxFO57UxTOpDIE0CVpL9fTU/nrzS1GV2+g9H0kVeCivRl8q12VxcIJm
7zB3B4J7CEjoyHNXNq3tw9b5eTQoEX3bUZX+zCqHDWfpJxwWYZ5ow5MjQKFe
9oOXs2cZ7UVBR+vTS8IF1cpdHnFUN/IBW3+ay1T7vS876TaxeuIUTJXRyZZr
6KTos37dt4XbBm6WTXfUEGGy0jh2yDLTB/JML37iOdImXQFM1cYjbmjsw4lr
ahkxtHA7SEPQrTmTrA0VdxAMLGCIOdMbsMyZroBCZCsOr8NlLn+DGnIDopfd
pMRCADC8PSSugKJvLG1pbaLYMWxHCHFpkTH4Hiu4zWDm4vo38u6vcQVQuq76
HxFUcJK7EDYOw6Gtc0R/f/0a4XyCiUyTP7cIWI7wn1J8Rq3Z6+X6MkOUW55C
HdGYToWJ3ZK4bPP5EqkKb82oLjdMPZjdmmb8pslRzRfSk17izjlzPd7Fc7TC
mwK7uG4PUpvfcDfbHxpDHZ78M9n0hhshTPxcppneLl5j1/yN4Iy7RIuht+fR
upWsg3rz7aQ9UK/5KrIQkW4c6SuLuKevogLnubMT0gYoR7d/7UpM/htObPIf
LHEu5MHD0OP6cxItYc0QkkCw4/P8DtA2W5liiCLSOZIxc8kdzayLnd06b4BJ
aEdufH+CpVrB5n5mGDfO7CXYQ9sGTqrxfbQncHsCJ5R6l515uqH5oJuAallZ
4lQsnD6BH0Wrn/Lt5DECmV8eUgp1G6BedmV3VldaJNZGYmY3JRZLfoOlDzbh
bE65940Cfm78vxrUdgjn2GxjkcoSUb89hFF0l9B+isAzsbkyZrh7Bl+OVfJh
goSu0CZIXFqx9vN0oJNwNNLg2fUwg6kpJ4smRFjFz4+IgxZCO0S25k4D1YA3
TSOGq9kBw/Qw0zAeiEtxrLcRZDmW+ZUuDwmv8UyzF5qurpBCjuauLr+cJMoo
QYE208HOEdtf+xPL0t6Kvv3/hsEF66/wf29z5/aWZ4yZkCz8WwF1Kya4RWrJ
+TU6u2Ga8/BvtJ+CO0gxizN1d62mmrayOveQWR0H/esgOiY0UgS5PZV/wCoW
Ek3BwU5wIKWO0fAE4Xnc2bs31CXxjAtuxcEMiv5WRJjNkpUd/QQryd89pJW5
yyWJnsEoh9YlQfgCE6CjlU2rvig2cDj8yP/mnNwx3ADbGADJQQIkCNzMxDDb
c7evmb6VhNoocIJy5Z8QSBJQerJO4I2kA8ubzd5TBe99rbxXKf12l1WOnKnh
0Jfcz4uJcNVd+tfF9Lzt33v+dP0/b7ImEnQF1DDCNwD1vUGoxrm78HlnoxBx
z+IFIDapCJoFTwcU2YCj4Tsi+rUxMmpVvpOsMpu0wg4rjjzjG1hRHqdIBlsr
nR070dTwOAcgM8fLiZiGL6QfhkQTdVSzSpOt1hH804zJ08Kc/q0hbrsWlrp8
sz+dO4VQmt4oX2Jr31dBpEpP7wCuYeynGbZ+RUX4jpRDTr+NG6NiCuivA0lx
X8N55cb7XJqxu1EaFuC9UhHbZfd7RIbr6niUvW5vdnzMbTZ95UnNAbr/GJPq
F3UUWeOYFNXN329vsWWUMcMzp/DdjAisaqk19XxKRvdJnpsZqYqX+YWdOK37
EyPE8H2WEYkiURPEHttoPUmjLEFFJqrtvxrOvppzHqX2o+kA0XmkQLq3d+Ng
1uaVPdqrDqjYhZD858/Te+u79RIMp/hakX+PKC4pnd/N9mAxbFRVFIlwAiVp
OoSTEZbgHmNpz6vStk1GhbEoWAsXZE8z8ad4kvCXEUGVSkPaznF+IrgySwDe
qVmvrjJ7UlW3jTMc/i0m5DvM4lfvW0x7ZANJqjE/p8+W0UanwW13ZXMg045L
ci+BSR/Vism/5R5QHl/dzPxQbaGJbODr54js9I2rejX1Q26jL6E7h//JBuRo
nIOc5E3+G+22+xem0nscDhKVm4xmg8k1sWn7FnndNMIULpGIGDQoacqDf7qV
GZdCW79eLWR0133S7CVA7KrUIBsHNeEBMKbIEwP6V7b+FATNvc3HlciKU3LZ
7llLFUUOpebjE4TS4kpM78ESdPazfTT+LLk4h9NaT9ge9By15rAKtTJqiZ0D
cG60hXU4ecvJ5iyJKatD8dWjQ4EMII4DpPwc9KFMJV7/kc6c4CEjnJSfoaLk
45to6ccy6zJ3ra7VJxEj1zh4XYScvPhjLXsF9S7a9SN5J4Aip++/Mdnd10lN
Dw9JIMabzkfpcV9tht9VOCols6greif7zzWHzIfMcN5FXm4Z+XBaXeWdMCji
DwMGSPVBRWV6kVOAO52SG8iEK8hXZ90JKc1Y1nokiZB87iC8GQ1hXydy2veh
LcDuNisx440PqOv7eqPhMvfW7vtf1DROPEx2CXp/AnGUXmTUc3JsWNyfTnA3
pgeANgToCQ8kh6ZVdMCFI8rxxPDOqU0u5atJdEoM2CsLUcfsbXAnMDPtHbnA
c0p+zngD3djgr7DbuuT1rsVWWIBBm702x7Z5md52GKKN5K6Ttzjli745WE9q
K1M/AEsQevLvK5HeDWzCVrekhln5OJpHhgL0SQxRALxZSdYccUFMyWCZkW9D
JqTLSFN/WB9rwkW335zKpTNUCL1Xe8yYbQl8JYElxw3eq7ETdG/OT54h/Mwj
PGcCnGJOtM3oFBZIGuyP0Z1Oumv9yOpi0v/SVwcymjRLhB1B4zDx9k6T3R+N
VvKbTwxTCBlUnMRgt+Dbe2lEOnrZziogJGzXYcZaxM5FNju4o4yw+3oTpZe3
yt05BZjpmlaQWrGAldHsLUXdairCA0lYCx/WRJOazjNkjBQ0lIAwxOODn1Zn
hPWgsiKZkAZfqbPg1+ChU+tGY2SsVZ+5Z7Q9phQLtf6Qe4ybSvH3nGBlZ7b2
w6xc4oPjt73DsknS91/LoY29o+nHzLs9VcoYlBXZfBa0d2jklTYJyJSm7eSO
KshaORy3jQhtD3YMBooDmcUQDN/tqxFgtSHNpn4U7uXAhLNLktPREuG/HFr0
6Z+xVYyRxdmd4/0VUHgsjASmSoE54q4PYuT/+Aot1KtEm9X10Ol2zhGOoD/T
5BBJ5QvNZZtkwcnUY5jEEp26r7xxyzTp4NmFBUNwRCIs+m4n8aHk8F89oaS0
HXI4Diz2mFqorVWoIU573JLpRR31bELrHromStGl4hrMcHQVKNysngam+myG
jUt6nzfJ35mIZnTXfi3Ug3Lf4jt+4+tjjlr0Hyf3e3wK+D9ROgPJw2TRDZJe
MFZFibvfZU/B7NcUS7kXoEBppDqITHC8P9tGkRnzpQ1EjB7jEF17Mvt28Gkj
9b9PtqqOBseZVxr38c/gN2mmLOJjly4mdq4h3ha9Byuq58MWnn0RAKguqb6N
iUgAn1NDqSagikYeUO8nHrqSIFBBqHtxzBvVN/ZoFYk/UuUBbqZWYrrDmduc
1dBbFeTUvj9S+yuculQgrfh0pSWtN67aZacr1Po6ruuJjq79+LaJ0q5vCnaS
+U39q/ooi6gM2oC3pgwMCRs9Dq9zdcHl0cXcsGTRde7BjYJhWcKWqTbvtS70
jYZ0A5/qzIq8u3HB/xlApdThbMufVIVSKRUJ6sWU6bQ/Q+fIstH8ZXPQ/IS+
7MXi/0ZTVO2tsjVpBRR3Bei+fy0bisQxhk+SWadw6fQrn7wULSf/az9mJn2b
kUYufJ4JAOmNDiuAa/1nmwFcrVNz/7jMGsUj+kby6gC5GE71ukyI+zX+nU4i
+qYBXGF+6EtUDShFxXP48vAxCu2xKVJt6ImDpQdf+45ACh+JDsNnWHKmOnzJ
CAuC33qcLH5JEALYdA51S/FlL0/L6h0160RNBCwNHrBPfcABbupK86iCpc+J
wMg9uhDbDTir84p4Ifc1IepW7+zuFL0OGGNgwr9sf4eKkIeKI/naSwOlgYkN
+l88VkOWXpEOFHSaDCukSEcZakI0dmT5n3A5oI7j6w8XCbwcI0PmP8PE7S1h
CsJT6NWDuGHfLGvEIHKu9MpM7YDDxu827JBkzLMyEfcrtWqDTGAEWbnFbstI
x/Sv1hXfpYtgSrKibgIrpgcUmmbiA8UnHWB7tnO2oUCp5Cd0IpJNa+n76WKV
9n6LBMjp3xE4niKcybG88tScHG4fMHhq/yHygkJhOhFETj68Z/xDsmbUV2WM
fp8lWepCwj5zGotFiB1MLseQ0k5zTAXI11WraL3uUmYW6DkWUPNC/GhgKBkk
qAUCpCPVhiFug4y9b93cPYA6aL2qfNxwSIEMPADDjlymjjlmSAYclUjtwkSc
7NL1Kme8S13dUQ09/elLI3kpw9KOQkRBwSpxishwnl+v1qjjg3WnXTmmcnrK
uONthUtZYoP3tNpLAw3ss6Yf/Y6ffaoiv5vSkquCeBz7F1rym/FhfqflNobs
2sv3Dzsof/nWqgL/PotVkDrNGTMkUYtkU5GN23tUnNTyGpC3W4BNkRUOQ+CW
VUse9VpXVpejCSKHJq99GCty7bufzL0sPRFY1mHFgVrM3OC67taJoDmAnmlw
pUZ5HIVtnj8Q11J/w6xbILriyK7T+cJMdMuixZxaAcDndF2GzLdYeW10gKu4
LyVyisBGmPx92Uw04szDpsW+YLN9T1y30WjuxI0ymAqIwDHyWxUphKvHzMCi
4OK0AS9bszjdIn2cX1Tcd7lF6HcIYEzMa3M92lhdbKThHL+l+h7iMNe5B2Fd
WTawkdsUdwI7yvMgjPJG7Wn7+ZlKlSTpLp/mMipwvCu5jiYZ9udwfr2WdOAi
VbWUB9Beqi5KgigwrosvogSaEs0+j77jTlDjqJeQcI75BLtFN/F33Tkpe5N/
/isEN/csp3eEk7UXyNoYye+b1srffSCaj1TwoxT1OCrLfNa800Gc5K7cw0y/
L9c0zWSjj1TDOqR9aLXcoxJC+P5Ydpe95W9Mk630XII/DW2PntWrqhu4o9dB
Yv69uoMym96QbgJaU/fwEn6XZ3WTojgFuWNPzdFTlI/Fd2WzjXTzfMb3l9hm
2+QcXGJpvFH/0rS+gFdRmPks4hMFbA+ms4tdWjYQdNx6kGXq4IUWmNlCY5/m
/V8muo7im4XAkJWJM3OiDqPScWQ68d9Yp1Xh8yXeOWWGyPvLf/JYYJtT4/8V
86A+QnITtaDVRve3b/3ZBa3yTkjXdlSoo8QkTRv/6x85FTM6a/vx9p5/qtkN
58NMQyDvddiPozp3Rg/3wf4AzZFW4x4KDIMGRZTo10yt48kv08CEYeXonpuC
4fdFUrJKqjJab/Y9zKELtJvF5Cn5vaOZwhEWy49AcEkoVma/WdH7yD9P+fnW
GPBgQEJad1J3DgfUswH76u2uHTBWxE8gVV5tScqj5LJGbhDRrmBUBKPg+bvg
fS08JAdw880oIyH1WLAUHETrptAS4Ret5sIOf1q5068Kpxeg8xP5CzTPivUo
UYeKz43ctm23dN/V/D3vdMdoSonPEZtCVLLi34GaceTuxLw+GypCEC4mblEm
lrEnIsSjHSU6WkiPXjiK5eCKExke9IKipFyduPfH1+171LOC9vGafOrmfI1z
NoAMcdfHUVHYA27QYEEgBokxK+dHs80hhkJ31X0ifHKjMljqkc6iGisvdAla
BPRjGX9hSa8oqu38t9cxiuMviwmE0U94gCOH0/JOab/9BxTSYIwCwAMykLD6
pYVs1iOxY/NqodSuoJGh74BerOHrUCNgHbBlpw6gMXEbim9I4qu7v+4oiShD
ltovML9QOcYru4/bV+NFYUAEPC6unB0YmO1gvIYdLKYWo8y921Eh5BZyFeCd
WIXaapKOp4C1ZJfx1SalYS1QTSRf727niB5KG/XzbrTDhszfulXjjbG7kNmb
jnkjv4ky5py/IyuhL+aPLTgVp4LKkg9P4u5Zx7wGLMhUTEdL9Fm0TrIbFOoj
1jJt++b7l/y9ou/nBPsWegyoHuBIrSk9ogTFWCd/FSNJqGQsSl+KWSdxedSa
UdV1h9h+QRq2cuv0BHAQ5ILx1vai8P6QCSIofaUY7vE2sSuZqjshhEZwdrlU
n5RmZiT+EpezBs61ABvv0F1eZOi8mvyPjQ23INy5SWcfOWG+McUCeKx+j8KG
JorQtbhM63s02hzXviPRIq4wyEYI1th/7OaXL9twwAx3wia+S8PgcQCPhBiE
bxfkX4tbFmRNi6R/ZBX1h0cgEw7Mpb1piOlmgtsoqeOEUUM+H3cRalW4gmK8
X9b9ga2PK5xU4202BtH3p9IwortSy1HOiQZX8mCVHKBXlfyW5+BxWzA3F/5X
0+7B0lqJQpbwd8lctKUqu+ZgoKhLSGSkdrA90r92Uhjozsl+ZergRsL8SHzG
YEvsrTf3RR/FLwTgnPQ61EqLFAW5KCY13/hjXguodkwqwPgTW+dFsRaw4OJt
DgVGXu9cyThrdjPCQFAEeo5i5ircbAlOFRjhOKIchLHXQZxqgHmbfPOmwKKf
QGyVnwRXzmGJgKfKI9ruHBfoAyT2/U9m19b36l0+OmfTWTOxDOPcAxjUD3jB
7WvvdleKrIBQgLDtAUpZBVNX1L4sBtmS3gLGW4Fwyx6Cud5L0+5yH7n0ew8+
iBhvSqLYSuVtvPont7/bMNEqNrboGW1NY5BZIUwAQfiuV8khGR38aqRXVyfs
qH2P6zFaXvOzKXkKw8M80s2fz+5y9u/lPjUQOdEkV9UFBB2oi6xiwjmzpwiK
u1D4ve448/r9Z+FUUg1pUPIYDkem+8L9AUwIJH3PqoIrTEDARMn1jgHKeJrk
09UBGJQLlW5ZYtrj5aSClS5AfxWOaB6+M2OLzwIV2LmsUj2D1QdS3n3LSyI4
onRxwkS1s3tYL+NhzCLl0kxEkK762g8Du8m1hdlwrJSTG9zuAeGbzZSK/yiA
cPIaU3l7bqctxMN8Axgcy67AaX3BxqSdQkkfFCT+zKrOz/x/0D+INM7Jq3Bi
+1H0sCHfSCdp/ubopM5TShnnMeSZ11df2ts6DQn+ZbkGyTRy+vdn8Sef58VD
BAsPregTdORTtdL2rjwdw7oa7x+mXyCUQ95miF+ZsxDDuDq3sndwMkLVmaeU
AQdYp09HjfH2kWAuh5ITzEY0DJxaqhhxL7rkrBxJhFO65yVf0xmTdQtA9Vkc
YtYMmuy0bvqhEQa6+UbPHEYJjwc6f0ChfaDTNQJ2mVy2vuZ2vi495qZEj/0v
eaZkfg8IVPg1kHqKvZBCZcjVq4mp6bcU8dndQXwrCW1drpFHSNmeQvAKRmmB
zTRV9TV8Gnmtf3psvdBe3ydbpoSaqLMDED//nGqcG6PNvYd/RyoZh+BkXLuK
jLF68xLdXKRW7mn54nV9BZjIxo4+MVqTFyTTaegw8wS/YgcYbVP7XZ1fTthu
MoaDWdMfrgQ0YUcRVWUtVlGi+oLetzFHesycTrTxLrMtn9EFISxE6AQaMVAL
Dk5mTCvqrVXINLMk0qLZ3fP/Sxtx0MDTKpyb6e7i1OdoxKNAyJMaDo7Z11nP
0v91zinBn2T6zt5dludKVuvjZV8iSwwx0RBkfSzUYaZQI0C6NjxGxeKNjN/f
1lu3ZOTaFH/BFRfth6FYtnGCDS8uymC/zD2Tw2TO+Cl9OtPbcRpCOgIzHg65
1qw4SEF258oMetlgHm6BATwGBacAybTw7OrumvvGNq/MFler4/r3uEHyDFpN
a8aVdBXL9empGWW5oIYWvWJV9LiJUWvxMRpWc3bP9vHnhU/ZRPpwOOTJEs2a
9l3D88Cc41J4gaZ/O6gAnZSAXJd/saeEXrPCLJyuSgkdgaCJwVF1+De8tYJ7
B16rQRDMG5dmfMKy5kSiY0plzF+l+P7O71iB2j99ypXhmtbHdHH7W2bOI7Ts
RPjTSciq7iH0LlS/b5s/nbclM30v+iwqDJJMDhCuqYeYSs4ZlrKQFaxOB7w5
0IAbtx0fyepsOWfbkKhSSjl6Gx7gqvJKlaBEYDfdSavFJLGtmZGjmNTM6SZ3
l0GFlT7B0SKJyGm26r/9/6CZCB6ITHCjLnRWbF1Z5h49ibb4t5T+noeYjiNo
eewsGbd+mg3T2PIznurEoQKAfdWg9SA5wP5q4ewbMCty4iDv+DpSzULGlEGJ
iX+2wZkb7dDFExRrXXJoHY2hy1B7BczJNQb7JFWSuNnVGe674IGF1qRMyIRj
kKAIinySsT5htBV+1/VgImsX73AFE3KDrPUe4L19i5uWFCKJkIQQ7UyrbOzn
xzMyXH7pJX5z8u3Jh5zVf5FSlyZiw/Xc+ZBamp+K7dqmly8CXfAw+nCi396F
4LNz7H2T5Vd95QGmDvARYE6aS9bBB9BIEs3VwvOajR18r+xw1roJD6U64AmH
YfyHJLyyPAarzY263D3t947FrjO+xLkpm9fR8dPLi2Ox8k/mGPFwlnW63z08
5IVcJfCPdyQhcS/Ugz1wG/wGpmbvlvx7zlb23/hwf55j9cGiuwv9

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiSLraD+qEb03/szXXd47zuphepuJVkXHNE8nbFeELNikSUsvaigkMGZlpJLSMg9Q0WFbkDZJNjj+PGHvTmCF8jL6XXGtMI2uVBWJPpOtrDTTA0XmOrkPJ/F4tz/l9YuZG02gCzKip2xOW/o+IJXro72kYMUD9u0dWr4KuFSe0IQs5VeU0K+LwZNlJkroAebvVmCmnWVFzsY2VHUQdYQCAldkahWfXbXbq7VW5c4he7udhlay07FhQPyoyFTfc2O4brWTYQyfZPrPWj3THYDdHQhPKObXqHYdGDOP3tqNdd/395UaagtGUU+kxTFWFz7OZzfbKWtSjHMmgE2eEx7a00gSV59Yc4X0UW2StM0qrP3+mSmwRbpGyb5g+zACOMCk8KbftigcD5lrIiJy9dDn2I09CS9sg6sJ4X34jN0DEBP238dy+Pc+DN+x/iVWfSiUdhK+2B7aghYMnbeg3E1enrSky0RIzE9hiIHk0K1d+qfNMBMQZiWyTfvuztG6aiUpfQhr8nwhnOAXUTB3laQHqkx3wIcGpDPWathb0iVsYGoX490RlX+jwLVwLzUNgYeAZ/TWlmOeicuc6xuVbq5muKup0FgiyUKwuxYGtB/LgjgWRYrmBF7lcuHsBPWMj1WXNR2xPwqytwzwSfCTDsvCD8dQxuLTMRQu5H6MBEavm+IG0qCag7zJpEj3FasCLJBQIRPMvo5fzLMQhz4bxFt57/crsiisW4Cn/t0erlo7j5jlJZtM25x/JqKBBMWro7zAg9sNXlG4k6hqnVrQiNwcRy"
`endif