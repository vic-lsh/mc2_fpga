// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I9C3HfWBPsAqkf23Yv5/zzd8IODg3kk2NpPJHClXVYxfozIfyOqOH5XCquB7
yuR8czmyJH8peiKcqzZh7bbFJqLx8kaUl+qtH/O6PmOLM0+09ZQSCL3GoudI
WMfHIdjzpkh3voYTIn8pgeNg7C+bshVgZpJF7+jW9ivY0zCt1O7tkSXTdHd1
IHM4lygsbK5JglEQuYNpWP5iQX7x3fB4F05AlmYyOZ1Si1VBd9kaQIEvMM1n
omygttaSVNfNQVv2GTD55b3Dho4SI+U7vzO6srVY+HutkgJuw4j9JwSKZ8Mp
y6eCsclHWU0HK4DXbsx7vkHPzVrugUxZRP+WHXjoyg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hXj45oitwxYKmgLArF4+/KhBktPtnljufY4/TTUiX2vgwRYlRI1+rcWrget/
7lTCUj6YoEZ25HfgkXMOlT9ukgcs9HEZi2P/tX5zZxQN+ljjoDBW6H0TM+z9
Jt0zGrGl4Wn4W1VuPFxKPbbXiDl4B+uZukhh9orV6GsUfL+FgblRCerXTkk+
3U3vFs15+8XTRsVtp0+OeAKtS9eONp3JNGk3dEVQcSMCQy/mQ440f8LMAmnA
T3dIFk+JGQ/YaYis5UekdLVhf7j0ETbfxVbwdgC7Bgv76ZXxMID82xQTi11b
LGL1eLeDS1/ckSLsJDdpaX4VtCokbVztwqmlSNlI6g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JTW0IkwvAb/h7oj7TvU4nxrgbDiw86UpDEsBexcIfqfy8VLLchibjCwaK67a
iqMOUeWDa7lxKIwAMQ6e4aZx2RGijMDY8lxogGPHtpVW3gKu4N8eUaz9gSnQ
v9aoFSJcJf+IZ/3MMorQDOpPWOSushwHkGtRnS1SyMeHVhilSVAu4G/w6ImA
to5thw/C/g28f4r5XT9E4vrgHqe+ecImtfX9Dio6d4B3nZdM6dZFIdXHGf//
h/JShJu0d9TDmpc808Auo4+jTxpO43coRdUeO+ZMCGaHZwXtHs57dmmHR3ZF
ZfHs+peB0ddZZjpAbuJIaUf7dJUKbB8RolrFQ70hvQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f2cZVNCHflrvHVqxheELcxrm2MWATaNO+n9/MO6Qd6r7YYCCcx0y4YOepEs2
oYTm+AHMjyNxp1YvvZ0XeUtSTPsZCSqzUz/sIED/ICGqfhTacBxGduePd4Fv
urJoR+e6vFVV1cupkDRF2SJDsg09PaAYFNHiIW1vTzxcNhs0r0OfLrKGiMqz
0vhHU5tLxD6jp6PG0TM/o+xBuK+EyPMjsvjFXboNeVjQiQ0fqFIj81Z77dBI
oDtHd70sNR9bFKSuWMHbVDE4oEZ/pRgP3wWqMBb1+0Y26ja5mjy42qWgwK5P
B7+dD72+x/9bOwN9gF3adeAyvgZz05tIr3gq6ju4VA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Xcka86k19Q8jQCLr4JF0fZd2jqsLB1idbISrHQMtH+40HHL91r4i0yyBYCT8
5jmPNPyHkJReyrLuc8dTlFTKQflMU/vQNHiKjz126fGhJyBlGPIdlqYaaqPf
eOKsERgKvPOsI8gfCnIKVbLJBjqZTBRnoy3wqXF6B4W2v6Nkr2E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p4gq2/RosCOdDpwP4zRq8OEmSOuPz7nu1MfcuJMI5dju7R6i/HG+jnfI+mhX
vCvpO5ENXK6ygIjJ9ERgH9Woofw/UjdKxbGR1ovR5V0hrAEViO00m6NTskeH
B6wmLZY8tTL9SfegEOg3G1IrRLQIajSVT4xBJsmLq40vh8DOazZRI/5So6xl
CSJdmlI5unAcBx3wMEFcjC+sOqmFiezsxg1NVmd48wSmVAxiTG76n+zLShsm
qLT19IDQ8i8DJo7opG3D9QWoC/dW1XQZrXqFz6ZOuBngyRBBICbSoqQiw3iE
AXL6YW1qUFVCDZ2YpOy6pByHfALSW3iU/NFiD5sxOQXMLh5EZgUth2+2ptoW
Kt+HQvbkSjSFhOOG1BenKdQ277HJjTkvvqUy7IOYRaPk5dYY5I/cSHc1oRLQ
+3n991tYZhCPTVvWULK8xGGZRbadLfCMHlCL68YMkKL1m7NR8hVBiY3AHJlC
+Fwb64e647HVPJWUpOvsbSbUDUXp+ffK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QQw85Ob6lQCpXqXE1PyXMTjCy3qZASODTFR8oIR1KSstTviCf2pwmO4wTyN6
8dQvJfFgYv8c2GbW7NwD+nH4wN/Ti+E5fQHvTuIdZnwGTz6iA1jvyF7uCZUv
uVZrEcAuKyXuFi/ShUvLly/ZMt22NS8i7uudBVxQlPSaZ7VuAos=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hYIoQAwb6Pg8uirT7ZkrFLqf9MN4HZKbpP2pH+oAGPGucIy9S/qtDw8+IEp4
+zF3tR8gaaK2uj1oEKeUt7cf00PkTC1r8IEUKg2Fuu+pJeIcGIlykGLQ0qtY
Khh5oFtEBgHqVDxJP9dsYGaHa1jM39GvrYV/D3FMYHiu8ga8LLo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 992)
`pragma protect data_block
CkqfIDwTxGZAC/3mpOOJPZ1I9idaN67PcHkThv49qecOXJyN26cA8IWjv6Ar
LsQpPC8Y3pA/ZnRuwowLxMsfr+B3L0WdL83+c4GuZCC4017rX7Z9sDveMtEl
y0IMVkqOBcUrD6riaHO5o1u9HM9BHO1FcxcF6BJhG7ke1fbhvhhaPCYhByRt
uRjVjyWbMWzBcmDY4N9Q98mqdXXoMG/om1oBkjqIhCyL17A/0SFA/nclDT0u
krt5qXJH7vuGCqWnvx6h4ymr52G9jL+D3eWRLxS2OFwPVdBPEHD+d3fTnQtf
2zZKV46D0KbtRumTVYKZ1U6pAN96lJkD82hjkxHhMoUOw5inpXvfplhdk9ZD
C1q1WT62oWk1sQfSCCqJ/eUXYJYYTCcJsnAePOWnmMVlXN4tNh0AbSD72zyK
ldbtRwUKhaf4sWS6j1XVaguIFApmXWKStPgZYa7lLZbF3vLy0UF/kKPTzRuj
6fSKIP0CInXYRMdIcaq6ftQponBINc8nXiFaJ6gKmS+zELaZ5fQipQyWA4Mo
hBfALvorSGhvOrtuWluTqwamSqOpPzP9bQxa2OeJbVPX1apYg9bgg9LziuIS
i+tahn6pUhXhr2ci9Ba490OQ6IeAKFT6LeuTYxqTfFhzUcWbl9fml9JTw+0G
qkFz+FmpEWAMTuDuZ5X2Wqu1tyUQe3PwPkTyamSZ5HAsozP5wr0YOcdvqBmd
NltNvQ9HMtxnTVeuEsO/AsqslCQlIcQTFk4EOCbVtKhSlYjmIWQqdX3zTUTh
sYZQnOxqLmm+axFrPg2Zh5RWOZAOSYjaCjU2I0qtBhsNROEFXedEHmSR7BxJ
ReBbFsCHp3nBecNj17oyXzUfH99zSE1LeWh2PxX/E6a/EgzcBx3hbw3E2AwC
EPY+97j/VdvO1kqJWeMx8F4AGja6EOaSE5mZEwYdh09zRr07rJaqJ6AxzCL+
rsZ4So0p5QBfkLCSEttF2pHUd207k8d8iZXjC2H3fbS9blOqSH5qzWFIpzWX
tGrhlAH+jLcHEVNfp+nwh8ORLMP+3jtPE5whKW84gA9zEyO57uwaVhLcfj41
S+MQP3nDMufykmNjEovWfOXg+A7V4su3uI/ij8jINu8x6ZVHs7Q3XM42onMf
X2w+QYIa4YmrmoQEW0zln+Kc8RiRWACLAEbo3FajbQtL4Lp1778AV8ZGrevO
saoH6eTtb94EIQfdAnWEMcXxHeg/Ada2ueeUjc89hdmMqEr9K8IFPfUeg53+
xYTeE7T70zyckqK2snZBFk2Ak1ygz9QLYSa2dzVM8JYzg4pK5wLTDookGkZR
Qls=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoz60MTi42sAEGm4h5QG79M+uVMAp2/2L/KDuZCW34BU5rcC1AGrNxSdAXD2Pg+xjj1RgzK2o4CHw9DWmQQpr70KMP+pmHqxkUSNd41C9LGDCGrSI2TVReaH+kXx3L9+IJPvT8wAa+TsTtbB1fBdJgP7FdQron3gwMBod/u6dGvCjVck51r0zD/KsxoY05jP/QdElkkgBNovTNC8TmYAUzgVyKMnUAAeef2AKpPWbP45FodRZSMG2j2rweTuv8IoRiRiWVovSVALjLLZJQYVd2TqWt/Kab8moSnuLpkgzd10Rx0DstwOl64enUS7k1BrsZsEzJp0jf3hPzk3I5Gj/6ROWkqERkiecFCaUxwIXTYn3TNBZZwS2e/ukUFsYXBx02Py2dL/P7neFY1mMRQJKNadPlFwjprdjOi8O3hbQgycSWAGHmWSQ6qpo+mzkEG0JV36pKZDgVZWPKlauyFaR6qeWPDmT3RGBz8FOu6AbciN/L8kFG9oAGl70/JV+DKPhCyEEbZ4XiUIWIQQDo/XAXu4DphNyQAltaG6o0KAqixcWuE5z+NhcrK1QP66iD8JeGuKuOTOjP26C/LNQ8HLm2rG064e+i0VPB60b/T0kFyNwyscOOSb3+si9cPnwSmUFUZvng1F78fJQ/fZSMTb6fgM7MX22h+b/TRwP85gTad6Y69fwoRrQgPVSGqhZJQ4IWnE0tf1hBYfbKA16XSLvWChNyC/8Rn9jnR/hl46qMq74pN0pbgozms4oKW5S34RiJKuHb5hWcMI52EY2z+vJK6S"
`endif