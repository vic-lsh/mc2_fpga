// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ot3jw7JwdDteFAD3DxepZR7vivpeYzKPUjTaVupIF2OezPe5QglVnYdUL+TU
t/st3Ot4BHkjovKaMTxuSF/Q4EIJUBk+3VRZSfoKH/Me4xZ4aRDRr/uzY55k
wGYSvbFwAu9CZ6JGU8q5044ny5kt2e7fCzFvIU2d8M396BR3IzQLdAYt2IRO
IVF+CRbK7uFMWfPloAmrUp1foCUgO8dEc5FIF7alEE532qejQSxKZrqGCyBy
mf2J8gSbBUFyDUEt5Pf0Ua6Wkqzh7uLrCLJjSU9mbbx6JorkIkaFjWozJI4I
Ld95a5BmEfgLmxPtIhcmNHCAKM5y0DtFYbuIBu9Tpw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W1l3tb3c2XRz999+5FeXN5ZqVEF2rh7ST/SuF5DPwSvb3QuTUQss+zDAV8FI
ZSjR9L8Vcjrs73wkdbbcaUmqqlhpKe491CfdLNjSuBZzBi4ffeod9UAabwjS
EaoMBfhHaBZrxpky26oqkODOdD+GwlLiQ6VW0E7uWZcazNxjbXBYCUtfRJ+M
f4qAYGCQU18s37rgF9VBQ43ifWKez0Wq/xjpZ7YB6vDghaAzyb7dKXHQsLfZ
4EB5pmdjbv6bx/Ld5vbeLqDyCqqjnuGn3KhKeWuWDhFI6pCBbffvgbg0QS0v
cOXFMj5wqexPNHwJ+qSYi8SpkTwa1CmOwsw36b0BTQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cb4Ur69iKoQESasnxb8mvd0mX61p6/EcvxauJpo4ewa2wjCRJSo0JLLP79db
RYQM6Nxhrb9uNO15EjK2dApFu2VEnstacx+JQSZjOezXjkwuGVoqNAU1aOUV
RpkEI8IerqEbVvjBaCOcClzloVxUObynzFWmW2HnOIKRNEYf1KTQmtaH/Oaz
wQ8gwRSc1Kub4Epmoap+H1H+ICKiU2fIHI+KI7AVgNdrkSKS+wWZMFpWv9oK
opFYhwiPNoNwLP2c1n3Obii00ov2QOiHxGq6yEoRWxCM+TPqxX8aEFWjx282
utBNP2M4ldBbvvUwG5GR6kxPQXKpME0fxukEvzh/aw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hBNm0ejOPeKkLGcL3atsxu754I1/87PCd5/ykPic0R+m+IyGZ+nnMNsXSwKT
DhL+Y3htGIYmQXfsHNiKpHA9WGIkt0v+U8rFguQyF1dNxLR2RsDfkzjevFlo
HH2+ewiATaj1pQO/rrQYpgC+e2HX1VORb4FzhVPMQqBdFtaweH0Rft87ZuXl
tXHV4ZqNWRCNVM2lR+ZWihdF1wzQb0e6BlMU1mLHTa02VwgpKvHgNWEkfHUu
08zJygBYyPFs28llQi3zyY2G5Lq7purD4/Zrprn+i7B71h74q7cACG7QGrJt
Q2+izSuCljzKCs3dJViJWWvm4C1zWkHh9Eo+3EMxjQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J8O8C16tPGKBmhheI5kr4VyEVEoHp3d/oqFiJamBGXKAkboPrCeFFMA/7Ss6
m6v8rUbVoWvKyZukt9i+FgQhBOJsZII96plPtdGzpYa9lthe8PfTVsyDbXej
0Oe69FWy/s8a4AihurMAuucXzTleNb6c3RbKZjFTN6kRxEilnOE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Za/oLauUh/k99JoK/Wx416HMXquFBLI5xtepWia9vCAjbPlP5We6dsycQSHA
lrBQgIcIfqTNBR1aqYOlPFx31YF4W1ULDjnWSI2uDjNSed9MElu+6+saBKFj
o6/Kxvd7T0wftV1CXKVwFB5w2+52ellDH52HUlaTzRoI9vqpzUDPiwAaibuJ
pvPFYq9kCXK3zMtVu/JdhzTCQL3ItkgNH5PIfu7dHCoLVoMIAhpsBGnmZTWL
qoQ06dP2Xp7/Wx68GAY1+JtpNto8qf7gglVMyLeyy3UNZPkGE4GDYXS7l89L
1Jfz2YNOiUxwWyHRV5qoUtcXpVLZn7qSwke0co7QoujIIx4C+dGXTff3/m7m
/PWmFxVqXUwR192l7uELkLflQ5KbhyXjzNpZMF+iOkHaQJSzEmrxnCp49N+x
ch8x7WC8LuzGQeVuyT8bRhLXI60VN87+GhvUnAOPOhLhab52m0TaRjO4kSBs
Kio7KsV4bci5NdwZe4RPmRJmr8jqXmJU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
na/MdNGHXNT4Lj/IRTNgMGDqybIcHLVjwvyGpkXIiJMlUgmn+LrH0ud58HFc
nNCDuZtsEeFShzno7zn4zj/N0W9zF3Pbfd67/d/ppaRa8itI3kLkx68zibJm
gH0v04gEG0Pb8sOwRdTUfOobRkPGMsiDs4p58hVbeWufE2bu6kU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L/gWIB3WekIXgvm02FsJKojE8YyL4OAUYiyHKUAl7HOU712xTFAgIuHTIrdc
xUn37Zb93kyAL8+9qJ4y+DczmzTHPyC73xF4UZNnrImljlPuOWc6LQtotEYN
9QSCYpM2y/0Iu0WBJ2jNGv0kuJkXbCyy3oI+RJF79wz4q4puxEA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8000)
`pragma protect data_block
V8KcmBxZA2pKAUVuFvAgDGsxvtkACoGU5gg8S19cpp0cHvkQcTCB5rWqp7gY
cgQUKXENMzE+tUSeEpTfM4QCyXPiz+h6LTr6WGbt+f/u4ly2INfki58aZL3f
SIjdBJJzNLWzYnqkp+Legsd9L22x+EOY85fFYRRQGTCOG+AySvMdIw9Qbb2u
aKJb+zgubj8uzT2i0Os1ohed1B1zD+hWfYkVptfpifEDrJaLOnbHEm97uozt
JrcAVrWTIcWEzJK1pp7uXP6SpUE6WxQ03WaQh1K3kekkwBItdWAnIaFrgchf
/Qzcp/iDR1eInxsjCa4Zdkn2t/EccIKKEcujcbvnAh2lmokKZ42NjA2ERbML
7AKy3l9VcXH7pxfhqCRFdijVvyCIJrzm6ji7GT5XczmU3Y5TJdjSqNpgZ6hz
VaFc66dvmOlvrSzw7FmIcyAc8dkAGNyPJ6L8xMehL5PsCBwIMydDwrT5BhQy
FrBMZBWio9YJLedNOOOxTmzT2Z9u1xbhNxWs1QdR5Jb5e6IQPGPczKTKgRQ4
vFAH228UMX0Hbd6hsipOChoUjBROwMo6ERAzD52PBOhUzT/vLNCX9oqU7f4a
LfmdfxsL4LjD9qP5FkbOkOGGRGeYFOCCbVrs38fjMcaCsllE/t2Ulf+He9nq
4/ccN3OqAcnQErlBFCTMfOCxws25G+ct8IoMhG3Jkg14jYk4fGKmxdwXDg2V
/wQ135WjSy/doPaGklnSxKEXzjptdGWKVov1HO++OwLCMpgYI3l96hX+rgr/
MhqJsJIvL36+15Hq+mInWStrl1FhhY/d4dlAsYtIA2sDEiZ4vegebZrEjd+X
5pAY6TyO4ovsMVpikCfzrDPET6y1EL5RZPSMC0nbZuTXExA073RVDugw70vY
1XOvdxo9dlXFl8JY+v4q+76SPfCySoitv+tF/EAfDJIAHh0ngPDFI3lWWAKP
iWlqZB0EEkdE6SDRUqwBALqtSp3kFr89L6+g2oxOJGBjL8y1tRg2nfZ22RXX
OzZM0SQtWskQOGG6ocs7TuITgXTUHOtH3EDdcS4uAx1FJ6iLNqXTeAyMfszK
Rhg59/dvxspeX5+W/4/bQvApubZizB70ZXf1+aI3LtuY0RfYa79zYWweH5qF
RQ+HGx0vPqOrsRGQQqI/f7pyCVDmQsV1UXkAfyhnoXZUE/20r7iXDv7shEI4
2caCQ4Xfma4/C5S/OEhPQK5zsoD7GOWnfljlBR5ccBPgWO+8z+KKT4QCSwPE
iCXkvgdZ154uht1C/qAcAP/UFkZJX5PF0CNIJlhuodAfqg9NjjXmE9CQjA8/
UdmkXaIXYiFIYcmqAbcv+cco9nnpJEwu26hKgmLsN8Z7bjGUPjz/0jmj0Poo
vVkDiiaKb7cuU3ddH7sIU4f9YAJLliJYKWUGmOs9FT6Eu727XUE00YOH4vay
7bDcYSMX0LO0ogUsn59zcKEOlgJqDN2CYT89U8Me4I4NVtDwOJJYgYn88OU+
IW7sZK5cbMw7Zb15wubXEyTfW/PXsaPaOYQuzipYeW+7vOOdLiopLWzFiLKE
jdhCVmMgam7LjBoz3WOc+ixAomdFSuaKEuuRgdVmaGHDKoiJ6nbXxlZZb7tH
AgaisauP7CNjiyBRmb5mjwFrHllHr7rp/oj+MC+eJ9/Xqbx+u/rPeQ5ocBA4
36rHsnKEth8NGpqWq/TVj028raB3gFxohGegDPQnFIWpSyJ/4m5/i+qoWZmA
Iis4JnjjTrjfCPFNOVpCRB3unDXl7mMNboUmnAIwmUEI2L0IRumX9+2qpxSS
NJHYmwKOdTjFuOZTuDcRdJZ8ICA/aCg0TGSI9kKuQ7+DLC5BIFK4mdHAmKbT
mgOP0p0QOt80SfMtkUN6hsqXcwRDIt8QqoNVqOIYGRejlA5CqC7p1mdURLOM
heeFMDEi5XL5oi2m5QlXVKJnHlkSf2zeMz8MyPYkf3w0CyHgTPj3/SIN/+6H
ppZW43wmc+c8jL4fJMFHVvOJRdw8ECBKaxd6pYnnIrvXDcBlbD3VB44gGiuw
N+Xd63F1csKifcE+YYRRl0MiAtyzk/W75+Dl8iZNP1c1JsQiagchsT9V3JkC
xwVj9O0sFNZIDNk1nZAGf9vnGa4//DzYO1vvbxA6E7AE5BvA6lLg76exMgjp
Hu2h3zD+kv/U93SOBIpJHHfx8jfQWEi+hSrSILfwlnfAeqcdlotv9/NiaN97
Rlv9J+6QQV12TFAds1odT3rHMIXw02jJFV3cQxEPXb0ENB4zIoz4g8K+QbvS
qpWP0gJhRblpk5+ZL5+oVDy5Fp6JlgR8rx/uzCHej9xEMcOlqKIW0wB9dGZP
DIRqB33Y3utjCnuq7PhVNF2KKIPoJ38A8xtIKrffh3luEfz9M66IDLK7vmwM
OCy7RJQHWjsDbZ7su9YKZly+XO+3rA/3rc5lpwWhIgziBKJvVm5Ab3n7i20w
2BAEcMImug9HY/lDKYnb9MrcAvzc/2epzotAmVytu/osqC7BEHJyG7pJIvL5
U/IV3fcV/ckJladuLLEJdEE7oVE9aTz3RWVuu/TsAeLdVFZuEPN2U7kRVOVH
ta0MUwEnxYDFeAXN2+CNAPv3Sw6ORacRwF78R6GZzls3N4RRqh3LmPt3hmKF
SrYTOTDxucvTe8Xle33i/eYO1JdLpG7b36AWwIZVGn5MXqS2qjST8bWy3zxG
/ShCN7zZ4hQZeVrEoOzJ2Rl2+OufswAod7knaDrOrre1McHfr0BQ43tlo05q
en7e7S4ZUI+0EeL4AnAagpagr3QF8yhrKpe7rnHjzKa/xYVVJmgS5ZEMXOfv
f1uVp/ZVSv+UGaU3XYjLblWTRs3htJM4hx1at6CMvP4pT4tTTgfGP9/Rwcdz
12qalnnspfZ8ZLfwgxKIPS2USExwmMcIfixVYjPPgLBjPM9fsxN6QpPGjAUT
jL5WtQ4/MuOAoU84js7WQC41b8Yym3tHM8jyGKEoCXzSeql/80QrAHncGK55
mlnGk7nj3j0yb9bWVz4x45tdxV9Jmz98cKfeHtp6Xofh/NcTfbB6y84/DdAo
VTb6xbAGmGMrxiZ15vXocFVt5DltaQyOzZgW0SYwSrlBijM7wMuiubsfFzST
FSpwfgZbW9//PBr8I8T+eCRBIUBYbpJjf1jNhFee4D4YL/vOw7zjYHPN0p/l
K4mq3tgpXX7yQOx7s3qS2KK/ugN4VZDR79DJKMZYig64GNLIDVcW85X6xZ56
pYWyrkCqWf7I6F9Fjuh5Tp2gAunBTOFP5oNFek1CQQODJX8AGD1wX4sD7yKE
YhdwmJY7xnxqeKhHzPeKhNdLCibOqPJOQBCeHhb0dl5PpomB6p9KR+JUtypI
WLslOT7V9Sbic1jKwSc0q/3urPxJRtRIzG3eqPj3jBGDp5l8Ek5pVw8owQWq
90G8QxF2vbaa4x0u8IpGXu0lfU5Gz9QEbA3brD6pSDQechLo9ikkMlWDcXKo
2yuTAThBMs3PhImaA8jcMy39HfmSuFrQ/XMajF381gopJ++xwz5jxPgZgs0B
lTyfcw7w6ZJLtzlrlBGnZklkIMLSca63YSS9A2W1oJzMQtU8MpauD0eQg0eO
WFQOPmkFPuj/wYbQQRofsGNzfUWGYxLme5mtOAJy3fhRatREzGnkZd7Ljx+G
y9kTgVNPBXIPmwMqi0WiH+bvecwRO4He0wGqh/+9uz6weqJgGsx7XNpG8Xwh
oneo0Jbb51VhcbkkStxSXJoPj/3mvS8wVRR5oNW0CRIzQCSlZUlMezhqZ9Wq
CuDIgb8b06DdA0ADNtNz4gZR1YbOjFdZcffSG/eofKu397Ci0fx19197JvQI
TIMV7Z1AAAkAUEXejN5l2aPdIpxfmC45lMVAAWcBjcdlFdbAKug5n5WtZHPW
FNPams/NPeMfsvtzEJ1yA4kzKlbjwyOWH5U7yDSBbhDi6PfXbbWN8GWZhH1I
8v5YIsgyZuIdKeqqoN2/pQD201aKb9NLjOsOzwzDNnlcsLwTEFwjhuj8uCZT
+B/g6p7a4tbC4sUN1DDNc9VqN4fP58VA8FFL13KB9WbwsoGcLJaHKqWKHoyh
yAADlWwtlZe0mJ5Nj00wYJzDkKr+NSvPEvKjUYY/Sa87h9pdNgJ1IujDW5jN
AbCG6XyOS4W3JxtT5OubSGkXcBm5t1p0hvJFmpYafRb8QKtGpt7fZncdMmJ7
u6F9AeCGXAlKpdNE3AYI+1eRNUvldMeC71MFmBgXZidF3g6LkT60+/woL07A
sytfdv4KXJ3qZQxJlWX3Ul+tP2QTHZICR4NJTyR4S9MeB6toFywENI/7rWEd
oQoxCjaO1Bh/xmGDUnklVw98mlaZtENhLPIXtaPNbdVoeev5VklWVttBzlIy
sQREDYR2rmNLTF81yjMUDtp8UDP7QhBbpl66f2py7TdBYD39BSM+rhh3IM+x
wqnxroRaZ+rz7ycnY6x0+V+MYU4KCVUYh7tC2bB7B4b+1KvoWvVRH04kIlZp
A9TCo2DoQ+8vp02363uDCOHaON1B6VX64wUNtpbzLmu7j5rzHZcZOvL2wdCr
nqHZJ4vwwMYW4H+PxtOrhv0tFRxmwvgkqL55U93LixIxbZxTrk4j+mR/I/PH
0xyFGSwfARasd9mV4SwMnUWOg1E9UwiLWX867blJFVIIg6iIFyG0bRCSnHh7
g8sDQZPpYz/yOEs4Zt7C+Z4DTSiqqtiY35sf9pZvsdcII0qZOfpjGcD/Ywmd
22ROhGmidftMsLKp3H9o/8pEsoBXnWThvuGup5hZZbA2e0qYOQlq55Frn54+
VVm56hf0PRdy3ZMbbYxganCGH+8QxlWOvIQ/RtNfZ7Dz3TjbCTxdJrWHiMON
VKBX7UXZoCdwmot8vsT73jIflg6ujYU5vJvt+r33ytJSc44GhwQIJFZN7C0A
cCle/Rfw9DsBzcEQxFK2sZ1U42I3rQ14dPdV7dxippATt2AaYqhtLao9EBRK
aT+1RQdfG6MM0iqIsH9OrUlIjjRra0Vdlf7X5ZTIpk0/jtghEKYmoXstChqy
aKhfH1H0rwR/8Mu2haNth5hGznjdqGnyBmwiP+LL4B5Xly6zd0+LRE/9GRFR
FMMMhMQqOPuC7TTFxeb5iLvm2UMTlgAVwU87GDGE1l4OJfWskH3yX2rwvXnQ
4Miw95oFc2dSKcTPdlUAPROgsQ5myYsOqwJztG1XVFtO6C9QkJK4s0e2C+CH
n9l6Dw953uCYmrdCChj/X5rcMbpMScxbUeeOD7eIxor+LWdiYhhvZOXwmZFN
nktk7yX9/bqStoCWH4aBe8eFIw/6Io70fP9zhL3jQPceX0z+HVB4IxuOLosK
fEj9Wkdg1uMTO9Go7IemufiwfCW92MqaPhk6TbX8IBMXSzPeFg89sc5WMvpQ
ZQ3/GzaUulH2fLcc5YJ3K1WJPpuQcT4KKpOcLRxVd1VpXinBGaEB56pYVmkA
xvceA7ssd4TqqQVn902k1Pmx8klovPemRvnqKk2kBdMogQLzvhhaVN0c7y6b
fZumeLpO3+kUBOfbY+H2hmwRtH/+F0sj4r8QJf3GPZcr9Nxi52ClRt/oFJwx
54BVoQySzesQt3uSWhER/hq1u9dBjcXDLBaXyW2wmM2fmKUVFuFvsj//vDvR
C/DJ5o12keXZ5IYfhHomBcso9zSirp4i0zCNkZOPxenmzKADN7KcVhDtd87J
YSwyXOOWqHWsgDzTJQZww6smHZq7OohGkT5B/LrWA8krklPPICFHEK3o2qG0
KETNJd+urjtERT7+s9lOOnwX9D95dCqpAa0Y8W1r4JLEzSlndxjz0c4DSTLN
e/pRIwerpTqfngsY+kwk08+uu2w065C/FvIVew0TgUzCKKKMmUTbhevqkuf+
RlmQgnYrddF86doGLknzrzr/KGjM1Ic9O3z67xzBUdTyLxUQOkR1RGLfCFHe
WULJ/b81lclS+eKcr43GH4ZsHwB8rbcSd/m5CbRZUT+926Pp0zfICPgtXnWR
QxubirjhK+YHZGiAQf+7IT7txkn1auGiuTQTjDbqXk/3yDkNE909bj5FWNjd
pQ9/4Rp8ay4OFI8yZmGz++1KPZ3p1o6fRWsORwayssucXWc9G2kVSNoxRTjk
uIrIMRb9xw2SEgk8rr8uROCx3kITQesoDDjifTxjB8UGA83GYxFGjGk+ibfJ
KuIbAc3wQxD2Tz8P/WCaDfpRUjSDlF8ehyZYoAw5yMSgl4im333HZVn40cnD
kEcPFJSSYyZ3ElcJ/6opTaQ4ss/HdrrZQYfXBKA6nzmama78SABnzz/u/U3P
c6j0GDaTKvMSqLGnBfpYq9NPrxZYiZDFAssdGldgtDIWPaBX2YvzAZS5ddVF
+AVsIA92Z0DzQOQbpPzJuWy6F/4fUKX1bI4QElBcHOLXwlOI1NLY9RgPd2XZ
3WWzeU+xf8MdqoYmHgzoeyh1+wXjlfEw6WolFBcpDPxXsx6KmXKK/OSExOWp
YvY/WvT4BopGfMKit77eIcwhEcFkB3WyfYNgCyCkiOJadoqqo4A7Q11SCQx2
Q4cIV4/JbZQlqq1+O2s6NcCrZjbnbHMzti4FD3okmSYaDnj46HYZHftoP6T8
COb0X7i0sD7ROp4zJd5sWKN5DkiQQreWGBsxNR7OeqeOW+hY77A3W9TtR9Ut
bcnYtJbPaKNKwTvNnLmIt75Y1SYmAuBVxE9+gitLUIAVzbN8UuVJfanise/R
eZaIehrD5dlWjH4wZUKRcs1wmX2q3ahVJTQ++qPTSdtbfxgl7oRAxibWPzph
nfowcuR7vH4CRAAmtpCz5TyZKBEaYk7Q9pDTnbLlQOnS1cUe411pMiv9sX3O
s7g644S22q+5PwtjFS4H3G/cwO+UQLB9HarryJZ1m2itvWbgaQVZyaLizJeW
DaITBNV8KgLCOl//b4mWYnzX+VV65HZukasCcQ+fENmI9wELGoRum3VdR+wJ
Ltz7xRD3z2kq9bFBGDHrLokjWYNfNuWkXCMhK9j5+D7nDu2xwvUkf/rCB2oP
ux+pUSyHsZK+iVY04R3dyF0iV7jjc+pbepnaEzZTzv2QYBeJgw1XQ/a2D/Sr
5682/tPG5kMJD6j/m6DtTjYGQWBl1IBYufWjtUk1n+rpRyjxszHp391/Jp1v
WqBvWZnR9oojHVYtIo/n57ix0at6k+5ofXKNOxV+fjwn2QkYxaGgk6QeZycC
TAWlTScefwf3m3E7cPZmKCtETX8kg/N9kr23TmRrCtfeh8ujCUUADRnnTNia
dSyDD8Yjo6Nq/hEALO44sDpWm0lbkdIVoOT4gPnCl6rPFW/vQNoZ+ImPjAsZ
UgbWUgGuyrzc7LROtPhzriXjCnsNbQ/OzGVo01UAvmkkXOdtYqzwsCSLEJHQ
dKoqJFL5yx7BKwdwnZxXm28kwmCDQEumoMEm8F2dUKLM7XaUP1IbmImgCNi1
mxVs1aKh0pNzFSm9i/eXyonB3C/rSdXmJIZ599NVtdUMS7A0GeeBBmjwxqeP
khP/dmtw8pQ/oSgtT8zpbAcjenLVlofp50u8N2KWG8+jKwPupEWhh7dOS8l1
PicvNwicXs1MSrL59LUGQAr6CqnDhnbYOLLBSb1Qubs77o0sjVcQdRwZVw7m
ZxFSawZdKA/6G4ssl11U+fgsNb45d41MyvMeCNLa7PTTC6tiCmVw8w3TMA/H
YDsXNZv9DUt8qtW5otj7r+tnHwruCyNeK8YI0RzAUB51XVHLtttRE4B7Y4TC
bMLi8BryG2z+N+xOK+7VuaSlQZA0PAlDvLuDKn/KnaZau6aSqtOdbZRZ8l+L
UK9MrjfZlFKuGH2GogMilfsX7gLyk9OtTdW+0rzPS+SSXa7QXuCjkOdq+8xU
1gNwTvx2Mr7RH9gP1D/cIuSG8n/69hIV8xU1YEsj1+GuBS07RLrlTSUN8MWW
wLFooLO/Sr5vXH0T0vjAptCysEC3k+xDbHhZmzjj+ml8xkYFTStsyvqfd3n5
ZYq4Rvd5TZCX1/9AohpWmzJRwYiEhzr84hmp08X0rn36K1KY9W6yK7C23l4o
ZDg7wrTc8gH3g8mnyEBaKouXEplm0l8yvjz7eYRnw5saa1WfbXW6iLXfsm50
6xa3OYoJ6PgOnQf0HMmqnDnR0FEhmpX7Vr004sRTBDkemJtWJlBxZII/bNSC
lpJkIhff3dcrfT9qlq9W1v3TfS/ClR/U8sWXDhjaX2s2znAdMbb63TKvNR/i
0lG/6NCJ/n7rff9pYMrmQfWwoRIEUugcwuHithTChz3cWlpkLnMKeke0W0w1
ckvkzcYfxOJOIPMtMd/gow3rO6nZgMUOUGchTKOpQsdtyk9Yy2tfWJDean1v
iTTZnrY1qv6kZBEOaxA0VcCAEXrbvCuj9pm8pUZsKa5DDx/qYPHPYm02+4Mq
Q3I+PYyxZYUEv2FWcT67CVs0w/feXcKmU4+QkCY5W7lxtAlWZjtwVE4cgd+l
FTPWop/SPV0yPJmLOkYAJt61B0/o80MRO+unyOOjpdUqeNvyustUPlX/PCKu
81JywsC68oUpML/BjFyHDKlq5YOdBWhvyETegEF77GsfGDv5NbEIC8JOM/cl
Yz2OrN9LZu3uDXfUYc1zGPaf4KAYH6YL+ny5Eykmq5EWAIZrljij2jYUUf9p
/kP47D2CjMmBMjivch6w0zC67880uSA1qR8INTZ9c9UH4ZISjyZZs5ye1Vwl
UoP2hYyqceJ43XEWWgJAfyYHI9/E/uDwFHPA6GTgoPFloq0kQ8OvifmRb4h3
flG5DkTr7X7UpqaZjs4JJ3wokyIf5vvzvVTl+rZOMzOVTdjESfiJKUSunY12
mGUM4w4uV2lSXuYTKeerYLrhQJcNgvy0al+qVrKbYGvVJoJi/px91Hi9TZQy
07mT8FCSd1/+DS5gDuBcSRgw2kIbrUaDtW36HnYTFVtRQor8aTXETous/Bxi
dfYG7dBNnRE0E0fBt5fi+dEgvrinMfilcG3cXuPNV621VL6CHaslI2xQIz14
BWqrEmqflLYne0iLIWUINe/qfQC4LL8OZaModP6KbW/9FSFCBt9XMvUnLC+0
frx4TpqGUNCXgdcOyGJUZpD03LLZiZnNEf9mvFM4AxhzlChqpeZky8HohfxC
lYZZf9R+5ZNcm14OtZxCNiKO575c510ibFDHJZ/nWklSbV9NXdWIsprNTldY
sY+5PMR69SnZYMeharKNsD0zroStU84ASxsPKNY0HOGOD1rQgbPFoKzfMXX8
7uZYHT1ElIxrfmTosqQYg+2G3OlM1vrWIuDlp68bXC6+Wm5xZ/pIXGRsvYmW
aaTykhqaD4kqlYL+lCbZRnC3DwO99KSTerCwEgk9QGepBO7YxadZsrR72AWB
GL8C663n1vpMOsHSH/KTY46ecJEfLy/zO34qHkISnaD48SUleStd7P4H1JI7
i20ns7UdYULsHQzSaxz/CqMnjXIu1zFFeqS/yqDKfhzTzRy+xkNqQWhQd+Lw
3H/R4vx5JlTgEblYYnSC+M9EjS9LjdOdXyBlCgZrHaNt++WYrTrJANQMq+Le
mxYwEnA4NxIR0J/nRrzf8bIezmJH5BSAie0L8ePJosPEo5XvlCp9kHBGL9vW
/a/ea7nCyhakmfPcExhNlQOlroSrU8IwIhtoDpQbXFqLDZZ06JRQ0/1fSkcA
NZKZ1j8B7vQUVaJYwuaFDj+/mI5iMIeJbZcOYF7LrmIiniDwSENbVwER5Xyo
8SP/bDkYjk/YN9yutoVmzgBDMShzK4//WVWIqMrYHuDLi3G9mBM9QFvAqM1g
9oSN/EZuSlb7efJSJarGo32YjQ/rWHkBQdaZ4ObB2AlAwytU6wzWz5L7Wk3r
TDs/lm9PjnNo3yJEEQ8tKxQGaoJXxreeHHVXD7WlwNUWffWcHcm9SVlxC1wd
8eZZ+7HR5x1i2cNs/MhTEih/3vUSyN0y50hMbttVxaLcEnJQ5BdajM4zepWz
rhbaYXY/7RmUB8vi5R5eOXx/YIosbdG21ZQ9YqgmzYImXbtFgEUZba4WtsW3
kkeyPEAbl+YoTJk0afC/+k7GVh8/n4B843BWD4uqtviNOPJPrboDfzqMbj4E
jQa/uQWJBx0//u8AqjP8uHZ2PagLghi5DYaVcEPmZWVj6C8iyb2BO7U6BM94
egj3yz17isMdCN1bWZll+XMLYuFybEgpyFAFhDG4+K5ogdSxj1dyRxnLe/fM
tsdFi+AwzJQapxSO+K7hGhrCk1H9eIlMpcnG6cpEIVZY+jXynZwwNJF7ilnL
ItV3sb6S/bDd9/iLXspHpHUiNhMwJs9plqmi5TnnqNLOYe6w2h76aAjnJYnm
2HpFR2xP8UK7/jWo3C/qHLCpkCssTd+CAMov6pgmDXRiABsS46eM6lOWjZHJ
qiaeS491P7MwPSU8YBtljm4/G/GEhnULy4Gr3tHCHZoLq5wzvgZm23LTPbMa
Et6JMmx4YT16XN1ixy2rFhYuL7H2jZGJyv8Z3Z77YxT3aKHj3nX52fCI+0dr
tfIKgF7kT0Cw1UXTTuZz6rA6K8Py0j59R68E6d2lpo8ynA9w6BLUAVmOmITY
6o/aGUnpURpmyFeCAXI5gsu0ES3fXu6pgXmac2MSzMHTSh8W5OTYRU+GiVg8
HfyrGVPYCv6Ic4/abcHgLCInDaTb9I5dX9uykjpOhuuNKlQ=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KzvAUcj2vvlD9u+ql4k0fsCoIrGjqFGSpFpg2w2yig2bzze4nxIkqF8L1fJwmznptH+wnR0Twz7uyTG0QXdIivyIF771nWKHp7RFKBfevdZyCObEa9yvCsxi57oRa182VVWHyJqsOBW3zE3x8+CqrVr5WE6Zb1nItm/rCvX/l4MHMeYwuvRn32O/jdm1TeLqRgOBwkv/M8U00G+9nYt13ADYw+gj1Zpn6m4jA9mwVUka9Z115zEXal2Hyz9flA2LBZ6Czmo/OylXAEiJSljW3Me82oji5QqaUIjARf6QU4pnKze3BZmu+sItTZrsILXsxP7h5CGwqH/+r2oR1yw3NLvej7md68Y9cwoZsBjoSAq8oyN1fO7PmX8Bij/P6YZ81ZiamxthkTUqWXW+45OVxLUmTfdy2eByKOiqXukY9G9ptkLAsxregN7xMnC4GuGbLZkrKKq4/NnZM6+uX2yCfGYOTyGCqbV9DVEWhCK66FLzZ8sqr8tE+vsNjVSAhduPXIUvbiG5pE6vkpEX8Pupxu0iVTJ0D89gFaiG+W1eXkXSFnZz9GP1Qwa67tC2SP2hapoIs2757/grW8OVtePCYwA0uhrJgyW19plaoCtkxeqSnwr5WVnbf2gWYKF5MuEmKNZMCPXxYd0L8TU3sckw9XPDEjvwkJQzGrUVcuImuc8VBCDrpE0fFvzW4DhXjIbGWZrjEBFodRhDhft3vsTp/+TcoQUFwovfMGIwZgCRaJ3zRbaB6ObLC0oH6pJah+LjWBXQ6jHc1rQmNjzm1/ZOlJ"
`endif