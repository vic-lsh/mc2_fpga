// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RxIb6hOTHGc+cmmBHgTexgwDQcXbohwWwATLLw/CN6ekpqoZmhR5HdjvLNjD
dBRwQQEtksLSDSnMU0Xo0WLXm+/ZqniUwF5vdQ+6RxnH+ssg+zUi/o2McY7I
0SpR74N0l1rnNCx/LK4BimuTaeMseS4rrNZ+BbMntEI28qqSSrBjf0fLT9D2
Bu2HD8p+jdEYzhPKKdks/g2M+4de9pEvQMxGQpbgXfxOV5o/AQ4vIRhTFb5L
IvhqUTNvLlvcFiLitFkqVajlI1e9fQjOeW90mWiNdKL9RVqNy3GNkHGV8EUU
0ihWXl0ca6nT+4n1zxzXMg+XUOMDGrGxeywMLbBalQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pVJlJXqW2lIzcpOdUfT5gBtW+lV2BBIDkMlMJW0FhC0/Qyxtg+6MJumSpYw7
52NtOY4tfbTW4FeyBdVK/1KwVxUygvrpCIzMDLq54K7uCdcR/YNoneCs1NdI
dL6Uxl8p0lcuD48+8xyLPTQgcU6myO24+YfGSpKLojuZCebiQJkoitIR7ABX
4A/iO3WL5LZH9vsXU3AZFj+FlCmWwJMWlfeIkpaOFPhrhwi1KxdEVcDwSom0
XBY0SaSgV68u3wZZflh6S4Jxjtp89TbFFXKrlitczbvVTxz5sStCd5N54ANb
C/Pg508IbDjVlGq7ObN6UFlc0p6p3rJ+Fwa2iVJ8GA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UtAakgqdVT/5WPjz6Lhd1vKD9vRiTLTtFM+BiM6aRWYPNDM6jHXuqfDuXW6+
UTE92fS5NjreZOOanSOQ5ntd1oumZFDWQrafVDijC9etEOpT/sIw/rNCjERo
M0+NLA86YZ0TV3XZL7lQLDhKV99fzmjOK5kDD5bRh5MQvFGrchCOnIaDACBq
i1kVIvU+ES2p506kWHFYFrO/IkzI01K0z/FHU8eX/jg7qFuy8lruy7P/IIsW
jPBD8WzUtsosVYAMSIFDE+a8a1P+PwN+s06OLLqdYFXWMqEGSmFKDKJwSYip
+exsiGtFS1tLZaD4Z9YdeOcJo6eBhsKvRWF7aLWfwQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IeHOyHZQ66sQuvt6z/kxpT2IWKhJaacHTGHGf6gxVHzPyeILysUrQ6dH2NgA
d5VkV6f1lBTn7prbxTJTkuuOzSCq3bC1xRI96cDaDrpz0KZVogEFd8JtH6w+
OWgrgZC777kGtv4YTSViS7xRPGjzVQtb+862dDaBxGgrcNiwOC070+jJ8YBE
cwE6KhlVHV5KfGNM9V/QXorvZ5UXOQycLnETPPVhISlUBfZUK66oLBVXdpcM
IyaplZsqJb60luOnav0NDFO+XDo75Wu9Pe+iXIBBi/42oDVF9h7q1yKBS2x8
XJi1ZFk4oIVTTl3GixheRNsH2jQ1kgL139AyXyRzQA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f1TsFNIKqm9+5Qv1H0fZe6YAJ8iVpMd2MpsDmy3jiVMRO/OVpRUIN+AGVGhF
29coAn0svYJxRcWRCamZUi5EzBEho3Ks1GJ7DjPR2WRXutlLUx9T+q+rW+/N
fPCZflLS51hc/dpuIN2HQeDa29gM42rRr3/YtbxwYpn2n6e+Kls=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uMy9a4VNsbpTCEU/WmBHX45MADbrj+pwfC/5qTn1wnYsSAPOxW7QkIBIT33U
WZCbsvQYsYcVsC2yFVgOLG4vm6wnW2iEcO7xVhjWW91y7qtkM1raS60FQ5wz
AtRI4vrs0XcKgIG0/oRgF3owVYUkN4e2cBt0tTY5TL+TCd3gOTkUqPguOc2Y
4Kdg/u4vM+IDiH1AwEJiHgRHpQB7HsPMPmbDHaZEG4IAZPb9bnSDrsBG+Lht
L7zwO6vzgezssBf/olVtSRDzwToKmS4YAxxh4/4DbNVv4xPFku4usfvbd83E
kIZP3kA5mkiJrihkjgBX+SxwZ4J0zjTQUSLSxyYJUXUieuoXEYjdC6ytNSnd
LiByNw0FrYnSHWHX7/RCnJuw5vEsvMFHkPuYwo4YdyF3P4qDozaegD1j5hDF
sJRIqKgbqLqo/Ta840rXgnbj+bYfCucSVxOCIZtqXgjxMX6ShxLVu3hjJZxz
6BU5MKoxiMMSZPE3COhwIBow8S7HJr5j


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fRwU1fMzZ4OY6TUfxxlg5/FPI19j0zxqg67aG9B26w214xdRYZde948lJfpz
FPVFdByVBqdA182PyYztr/NT72reRa5FdsHtQz5tgyv76mB5sJnxEN/SKS0c
vKvnRU/am6pabufZo2P5x6EqOhsYqksBW1PMl44n8Vfv8xsmFCk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PLxU0oFnKZVbvD7Ajf99Ni3tResT7S2sMpoIMqNPk7r8/S/ekghFrcs84gsO
FxK4Akv/KqhcAKLthdOBUBQpFOQcAS5nK/ucK+B1c3V5yc96fKdZ9NTkoPco
gNWSItZELvavnltTRlv+Hk/syHhr6hf9IdqYSB3NviZy6HVCFWA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 64560)
`pragma protect data_block
l/dB/cWRi+KjG06EMBy1iJeHDQRjgowMQxxS90w4+R55mbtezyZdWLI+xdrk
bmarnVZ8ioxOfAAa5gTFW1XUmlfxaSPqLFDdhPLQEzPVROgaJCxkUaEPn2Ig
o7y839cWSxPVQhWI4LLEpSkRVQFDi8xbZURZwk0ZPvykn0vKTEY7w4hY932M
sjOjZc6B+tIIK8/iDLzcdD+8hsRKdNSKjFsO44yoXXFCrV52evxPNki4M+BF
q9HSsWSuUdxFz4piYziztib+n8bdxyWVqyNDtVwWMpr5c6zS3L4phv9hcgcK
SDpUFdhYYdXFa9rjwguuYoV9FXwjVncYkXeJ0bbsS19B6CO3C3WThMcZkVbZ
/RXCL7JAm7+0QOHvOwXAB/ehYHUXenjBsTvut6UCv+P48AirOyI0eBzLFWUS
5QI9pr+lOvYalWeM+3bCcA+33FvRrXgtqHL/01aVG+AteE1fioIWG5SJXB/z
jBy2Q3Jct7QMWkuru3pd8oolEs7k2RkRumIWDsaLO3mKdDLy2JLaXA0veVZ/
XK+f/227RNvY9HMLBo9bTkLkH0WgeheLi8ovsZ//6Kx5GyW6ioYbOitM4Ws6
T8xThVGm0Exl5D6EDa0HnRPYHPnyBASM+vJpfMKmGjYgqRFADTmZDEFDa4oz
EdLKiRRwzqQCnG1qzjG8Rxlthi0XmJGdZAv5MK64+HMY8dNx7nplPZnZr2L/
vhnp4PIDCsPRiUAixJEgFeRztJCbcQs1tiqJKNur6tworqvH3U8BfTq6FmIH
LWBrrP6Wzbt6rzcKxidKDRX31SYLuI9zE+mjVzEJHJbWvsJ2xDgjiP+7bULi
dH/EmKR293C1SKzImihc5KRb5zQry50D//gpQNC3cJflYJy9jVqHy06O7OXj
VRqD3ZxpFscUkCUQGF0oTCfShRdTUashhAg7PEBIKvrQQvPIGYmGpaGwgRZR
l8Kat+ecHab1HOjTz9RMKGdB9M3hvSQ6kB6Ak3Z9RbL8FvTa7cndyq5pVp0v
gZdudIqzdcYRS5g04Kx72RhSbT2oJmaXRUAZtofo89uRR6LvDZiLjDdkn8yT
lNKTR7WUZeBgT7+LtgG3uxfNCNpXPQQQtiOYDygDKQpnEWLugwJMXWr2bPGF
o90VjrymfpXDKU7DhfhwLde8o2VQxNF2KD7VFJudfhyF4ijzh5YBbnrEfP33
N3F8GL1t2tckncQpHVOH1usdBG6Ma518qBouANBwEEIpc5EWApwykfqtjo1j
ObxsowwHQMwup05xLmEVhxYP7WjTfdUtHqzRLtsSKOxGluu/mpW12YCphZZe
4wm1CgqBIuf7ya5fNGrNsGIHG0ia2WwzzCk6mjph+F0Imog7gG1gyvFmFXS1
2Mp/v7noja/QG0oNFZz+PJlwiySu0l+UKcbdRlyCcwymzcha4V0+eBsezaef
/6Aolp9BJBl2CXcPabR1JB3oE/lCjnR7RNClwOwvdlMUB7zLHxmm9/eXl2da
tKfhBBqgtBtPwHX+EqvLd7F5m11ls1AKRwwOnImwguwmij45HinfIrqNX3v5
++oXNv/eDIZxmI5RhpwJ/pAwyqqf1708fBELPK/OVAQpRfBpEfwOAXK3J8tU
eHzMT1XvhQfq0+UjzftmSxvtsSHpPhewnyjynPVfuXmG+d+H7DCBXoy/MSt9
RqdtPpRsr+9ZjSOL8wbTwyOyQweaIPknZdnARUKauMB09fpm6uWBiN+6Pwbu
AJEmlkZgYXAxD186tsp2wVNSTzvl7q29Ly3pk2KtPBbOhctPledvYAat5whI
9aLSxfEpuzlMNICEiK6y30LCIANMYX/CJ5eZX8BUTPP2KTMeuvx3sglbDk+q
QLDt8yw39ICQUE1YE/qncMAikzdtX9uQqYxfE9AuAwZ5YwNTCCntAEEcwo9u
gxmLR772MQIEomYgdgZX0bRZEsrycOmCJh1Vfiy/0OaZw/c+HmF8uCBQ254N
KJyn/uRl8QW0u0NpMqUfj0hldqTXmJA+zCd69C6y43vWI7MVBNROSzU7I1jL
kNUhJiloVQvFoAFGwWgu2LYuIOk0SnaFyMKwRrHokEyWX0wXgJDWfbf7bjyB
3jrvt/GSptIbV7V59UaXB3JdU1ruYJmhvSErWEi0QnL1R8cJJHYBc3R//54t
/eGgWv13JxcRkd0bf0bs/BMZsiToroFi9m78uxGD6BiVABYhSkc+ff86JE7f
ByTWaJo+BroQwA36dBkccHCQu9KjM+cZuvR8qR37QL9OZ6VXCcnAUTVPL7FW
/iTaDo9guz2uVP5FNa49ONfwgYFcnkcXYCL8elaOHpgvf+4KtxhTA5JtKVLV
1vyA/QCCulY/bNggeviSby3VGxG7keEcIlJ9FqktrrnGBo9mBI4DicBUX0PU
DJzXRGW4UcwtixyVMrni+xN8zENQDOQ+YIXAHGupmn8Ve/NfwUR6EO4Dt/13
aqZumWvLGrt4mjK+b698LkrTXaWONBfxT8/k900k+QqxHWBAAlapWSg402Jq
7Wn0T6bZvlO3gOV1ZsbXyWLObVAA+wJvwmnINf0xF4S/axpwND9sO1TKNkUo
LUTOsCGwO2Zus8tfxlsgLqwtLtyvgHP++ZUSUYto1gjwFlBn4+K3dv6+mUwG
EtKgqF/jjkUobjGcoWvZjYbI5GamZ4xukoxG+7K3ObVIYrLs7Hs1eRIgdWhK
2S6GeyHkeKMW5xspOBNPZO1+GMW72bzpGEU9eiGRa6SS7EXG2LGOPK6uqfR+
TramIp1EdqPq+hGRPulmxJwq/gIgbdXMHkpUIfa9OEks74rj+bwZeT00FPo6
o9c5QPij7TL/1LxVmHPupLYVhVUbgyf0slEVMVHqkbdrWS51ROBOxj1s4ADd
wce2SDiAnKKvQlIo3H+vo+DqUDG/8p9LVOEoxJuriHavH5NfaKMzmqHT1siK
gbsPy0nIfI1Beh9vadb00fithTrsblAoKT+O40fWuvgy9dx8tM+qmtQsW9si
PRyx7PcGm7MuwPRiWpil51oPqvAvrdPP3ElTm+0k97RK/9Enp00eODCdNdoF
H+C7XoLisBXbiUtjhIe4tvCptv1IkSfMuMKggTeT+pm7Ym2EtnTusQXOWiEm
tSuztQ4AZohhRUhS6dkwuTx7SCZOnDE1hcr9PVe8WVrefRtZgCKCl+U4Ogbq
+zwyRd/U00k3iaIezN8XeeMrPj0k2+AQ6CftezbeN4IS1U9UA0hwIbDjTkcR
Rwsmm6y3wiANXtHRC6ExvkRkKuuPgeWR7k9VLSRGJY2UaVVzjVyjVzEOXYDI
Bd79O3TKLrB4uoBOlE54pb/CyRflirWExPpCtR2THCAf7kTM9W+QQQdmNfP1
ODD9+2yHZLYwb8puLvuDPeQmcmYObuWgxrwjh87fXLJuw2QmzNrDTtMW9Pc1
3RkI7Oc2gLHXuJzXMnL9wWCGiRCzXzfFMFdph4RTo+kGjHJdESQXwfexevnW
NpixYAFeW+sQcvEvT+E6Kl2foFHxzT8A5cweSqmFK+Iu4b/dxUACjBtUjZKh
aGMsFz5BCWRbJZEpt8LxntSlvWftp612ubwAfxt8Zfs+C7f9TcAVBf1px8Hl
6rnWuKIOnHVlbbKuPfZVFIjt0ra6n0+Q08pa9TLsTVTGwp/Y9KW0mrrZiUi/
084+4vTmW83K9+GkBte8jTBe/Yb/U7Rls3xJft4nyFySfwqfy7TjDFpR2Khy
BzvXGj4Zo1WQ4C/cZm/LUx0X6A5KVrldmVojgXhiJbcLQ+R01MAqdJA7FvCs
AECYaLiUO9+4XG2Ah9JEHp/j2O2R9qTsrM+b+qOQI2QkC7gV0z2mS6R016xw
m6Qdo3bfmMMieGNzW+lPSk9cpdj4Q0Xhfc7Z6eF9RjWZsi5Cm7OyjxVgFZwb
Yo8L/uP5SGFCkXBeQcPzJ76Qr/B9BEYQU2C4tgFX/HNjm7FKgE+Zyfv4Z3YW
G2xIsg3aNhzFSnrzv1SoMuDY6FBVcjYVvld4BrVi0hsZYludWO9Q3NPXSlBd
pSjyl6t0ROA3CVJeQQDwUW8rI9pyUoKLHjnRRTy9Umx7gB4qldTbhS607wwI
ZP1eQ3S9kL/PMBc1EabU9cSgyNfIlXvUqzqkzEj+eDocW6HXuMRIgz6y3TOG
21kikrAx0hutj06CdaGRVR2uhLmHsLB+fqhFoagI1UeOtyLt2wMPFHBGpjZ7
kcEnCLGYPzFnrDc+KeuYPk2iLVcx5WsrGlwada6HEHQ+ETezPksu98fEB741
azyLeHRN0l25BTg8B68kbIuCL66GDyeuzf5IIIaJxyFqV6WkMMgOY10RnLcB
awNyxNxmMClcKpukLL8gSeg6tEENkg6i1bTe8GmimqbV/x0NGjlFIgmR65gf
R+nL0iyFamHUVxtoEdA6dnhEg4NkV0CU/7F3myaNqQn+ygojHtYurFONuitj
Mjt4/Gr52+585ivOY0VE3qNHikMPhSNMsGUNkkn0pNNnNwX3f5hk54VbDIMv
w17JwPIX34Ne39LNUGv9gZ7K07I+zjyWcq/Hg9psaLM6DcShdp0VYzBPOlD2
2yrheyEWB+ZV6OWLzCpAGxEScvCOZJfBHuWG1pYlipcFMy4U2Ul3rSRAdamc
JYAWE0/4nvNsUDPS7fFaGQE++Sa4bmtalDOzvZrmbpXsvmGEZJdoCxUIrcpE
jYrJ+QBDw8lR0pwAlgzxLYvl/Bt0iIh+Bv67CxGpwroaZBo4RKwMyUr8L9lK
iYCWklGULtnVFec6AOUD3KKEW7kzADxj0tcdBmt+foFw6V2hKR8OR/DppSBV
d4nvrlOXuziwIEpHUGiFMQCW/j8nzByLa7y+LRobg50wPZSDfX7EYqPKp3UG
VvtSAkg8xxxaRPXv5TGbMVM4dlistwuu5nmvz/WKSswWxdUvJxCuGFVPRT2Q
U5c+ZfBJGi63C1vonQ8OlZToMJOvupAVeBORBbBS7pL/f8REJE4SGLUYUoOO
DzT9ZLr+LZ9Fm7c868PDXRlxLOwfV8dqSKXjP6JF3Xil/EeLMxHra+ZVM5uG
gab3B8u6mHQEEphKlQwhBN5sZjnczxMquMItb9P5OS/+FkXb7H0olqZnjItM
bGXPr15c+v6z+LDKPu6GlEZydn/VRMkDvgLm3HGXEDmV38R4QtJUUqIphVne
4TwBotpykNy+cr12OQFSqU4QriQDPkE+xYMYvB2ojnSlj1xeWhXB+VHC82Pa
18rJkdXTlwUFL4MdoTWpNtzo6lnofFGxthL08i60cCmkVj6wdIzdM3ngGTDC
RaL11ycYCxDSGyStmCeLztfsA3UMeoln4p+8ZPHnhWZMZK+bxfwZMdCbKMTN
2hNvjfgKOXwXea4vBFd6PAcMC6sG4eXHrU3p6oEqNsjbX3HyA4lr1K8bjUpI
B/D8lhreKKGnLBTv5p7fwUYSqdyE8OUNfkOjSMJAPh3QJOpcdqVH1a7ENIoe
dJVb0nhun9Rpke35f/kVygDYyBz3SS76hBTqIl8Ci2FEougVzJ5ygB4jrk0X
ucuN6QuP0yRl5QrAsA65pgSTTXE0wqcttUea94s/K8FRWMaflYj5hiaUqqr/
EtR0gpXbCZbjUJgiLYFXfhSB8BIAijc6FW4MN6VUhQ3iR8sxuKJQoKDCFv1v
d4P8iAFGehIS1NF4/sVJ+dvNrys/8hMKvh6bvLW8/GqfhiZlXxwfQqr6J/ha
SHvwOHynhJWeZN67EAFsJKw0hxzyudKULQJTU5ELCN1yIFRu93FxD/jV34AC
u+rYVuOFYePl9e5TU8iCBMmU+zPcBK+xhx9p75t2uEo6o611QsZs1GStP7xF
QhwU3e6PZGrOYDaPtUiE8daEQ3XG+zRTA0fYoeDdZWABA4559BcXpCpBRrF8
1y1IVzmFtEmGHuRK4lUpLyITN1eh5ZQj7mFFp9CatbHCAP+ms1ubFWYKlJgF
DXqaeKAwwQtxFz3ZCtNt64IXnEX4WAay364lSDoQoEbVXr1isA8oUozrndGV
l6Aor6g30WVueQzFNznPh3eV/iMi6qKLFhvtG3MU3gaI2Dt4WMznQcF+KQBg
6ZD8Ty9dS+Z5xCi7JFIAYrtQyXQq1AaUKoPq36fV99W6O1FbBTC7ESI+5M2C
0MCv6aBbpulJgcd+74X63XD93DNSaSLXoel93MNI3DL3h0Olr5nG2y7zvipV
qMp7pm9gvaYtGwSHB4HsLsxmWwFOOEAXgfktGPTcEtf2QSDkcIzHS4Udc1Jy
ySzwuf5934EmzR5KPP8AX6RYVG30cttsKsM6JAYN7upWCH0HmVdjh3YCZL75
Bh7KrfEU9dCWMIxgCdoJDt6nU2QcajCKUoWUZUI1pBwttzxcCx5z1ErsYOmp
kovZwSKuH7KENVt0kRUznE7zLR+ZwjGJlYP83wa/rxjpo1B759oYv06aq0Wn
U4ReZ24QS0YgdTzUf+qWYZXMIfyEt1AthTZz4sTauyE7orF+9N/HXkc5eA4L
lcD0z9ULto5j3SbmWc5GBz0RY+3ttoA1E8yqNq0xoIZj96SEQRSB/He9SW/l
Ilqf45kfgGVB3v3dSgyKJT3UBJOT68AQUN6UyIxavc0DTKmveRdXS7v/cVTe
J9P1nmKfdIljHOQNt2br2gplvgCdTwPjhx75x1d8b+3zTf1K/bk0BFka7Sf4
x/At/KB/8Ea9BQYnbrzVSJeX+esBy/jDKW65IBKpKPGaf6C29PhKJlXhZ3Bv
tbh7K79Ac7HnAsm20r1KAA6SH1KAH0fkzjSlXvMVTdJajWAaRqmFthOPUEHA
eYSdY+xtSDMs/ONAPiKWdssXJN2ymZPids5360CwKeuMvw411Xwr0nUnx+m4
I1Tgci2TIL595iJF6jntOTxAE7C+KgQBQpG0Ft8EeHM4PNK0+Spv6PQ7hNEW
gQqd/NDua7D/exVcJNxvE+5ayaZSIsGGg+L1RsvrCBTIjStJs55x7gEImD2p
qkITAqJ0a24xKj25Gh+GgZfFqbo3pVwEtCBzHgKsqkRa9jjRdB8OAJQ7WHgv
v8t51R6jWlfGjXIe408wI/5akhQUHAK+ki0ppFHduF3LxW1Z000q4iNKCWtH
Xqj05CGadKGl7xORUdJn9n6D/trZqmZdHVdhDdwFWAuwOJbdeckMsIoyAQXG
bgbOgvXNaouvjkHUlW5QAInHjQGDguNVaqDzcx4/zwkNAxKdHY9nTZ9Pqt9w
PCAQueRcx0Xtuk7FGPfbyNW965sEOGlf2r2E5coOLdWTPrpO2PQsALF/vesD
sKMVpfyPh0SYUKbTs2L6YPuTUmsJBfQN/pSVdcGAr+0gZrwlUIB5aXugmgYH
G7BKnfDTPGoac36pSo8pYP5QsyoEQfo28NNPuvxcUcHK+gc1Y4KdAgKrxcI8
ueL72Vw+H20jeUdFxR3hWI+LvMlce1czRnsPa5O2Fov4R3/EDyZpMuA/WRYN
zFxzkE5nsvpVdLzhzHuZczS4wumdZc+rfT8+5NWheymPMoZ32bhVaqeeQigR
JDQy31nmPm2KkbTIYc4EKDNANzKinKcesonPYSTzrRDunFYRFUT24kN1Z/3O
TZwxPfPjkp9RI/FpPDaoZhkLpCdEti/KhrpJWDOxBJoCDOqfU9wa/PKqE+CX
MkG3kgzkVTEywowDjzJ/mEotivLdQ3PdgLMBXQ8vaTV4bc4amMgdKYZasHhp
TE0h7tQD8oiT6K4au0dvS9jPSjIRuwgKZVjo5MGfsp2mbTnIgp1pkYmmGk4X
E2kY7jLE2U04fKeHZpna59MtIILPA4lmckYofrvB9HCFKJvtixNkKNbwJDNM
dUhBrurzZ3yWSJGrAvhBl2UtOY8UxSps+2y2+40RS876wxCD4hbLMEPiuGtC
SFpSnhll4Tr4SVQE16XR+McOdFR2ORWSaJIwQm1NS/TN+UavdgxcEXIUp5lM
yKjDLbuRkTJFBJyYeG5UPzJz+bnoOk+yOjqX+ovbq4XxpEMRlbWSjJ9V3wip
tg6saYzgG99HdCEJzTH1YT3MWR6jh4+JmehOn6ihbn3+skwrC/a46ckyandG
Rv/f7fujTTCsT/kkyq9H6VT9q2NXq2DKoIYoXEIhqaK3g5CBBrhFnKTPzkYV
BzUtwHGodQvaq/k55bAz/tPUT2noRqJrbzlwF8ZIsID46KEJPT8fXeQLk/2B
ON8vL/bg+NJmqpcEvrrloXqxAHVAUVM37qHXDn/xshB3by78vGfxfvrusns4
sLnTQ7meeZRg4gHtE9w0CbYUQf9Di5DMligJg/Hp+j6BTMWwm79hlb156b1/
6ZLZwv2BE158ZFNvyUvGSI/Kli30rjuUWyaue7n8fz4cTrxF+MJ4ggCkULqk
hoxe+aXiKYVm0SZDwHQJQSNrpnbsyjMqPxLx3KdBzYoPoMW6mzVSUtepJElV
O04NkL/Zrfdrfz9YvNO84GcVlJNt1nphnOHFqwNFujZyWWU62mhGwUUWCy2z
AvcKTFGFOPvcsIjIPa/LIqPNVYGI2nKiYlbpdW5SZkVkeewSKT5GSiUkH6uH
XlNJlXcBdsW9gw63IoBitHqLi+M90m9topCrg63ZZWjdxXocZtZXcQ3tOGCV
SADz3aog1g+DVzDP8Uvn0OmaYjA1XV7kMdsyq/DzGRreG3TYw7sKQlRs9U1E
qZ4sFXMYUXPu2ve0I2WSjFEa5XlWpGHjozclHE5uTAqQq/D551xMcSjg7PaK
AO+2Dlm4yQoB/0OycCkZawq4950yKSUz4YNDKLsvocCPhNQocsQYNSLwnnfg
NmCz0/aENCZmprxtda5tq2rIq+QmOnjz1ln9HMvm8o/jGLJSMd5pud2HY6kt
MM/G/NGeR5En8zss/a/EA1V6UkeURFwa3T1QBAg2q79nCYkcANOaIjnQjloe
veCp7bEVmIRQpfWUpjPmq137K/CsyS2FOBN/9oq87yLRo8heQmuJtx/bUIQ+
QfhWlOF82hZbWwtY/FMxDAgvZ0wSe5R7TRKyLbmYUXTCQLJrmfW6AW1j+ZyM
zBH8cCHhnWEhAwgf+t0P8vDRdZeagcYhvUEHagZ2/nwQ97mKtJr1oPkUydqA
huhto5mS6hRnArw2dbHMAkIhFP5DfY532i45ePE5CTtzMUb8BqLrArhUulNG
jj12GeMxaY6GYEt1FeOrqLSzFWuSTWkDyl1VUihdEzIVPNQ6WR8WMyVJOCyq
euiOnEzNHT0hLKIGDqYktAjrAZh272UMu6eLhqohfWkmD2QRKQFq172fSU/u
eEVHQW4wYOWZopOg1a7f5KrlJLW68HBypIuDL86Ij48c5GrEJsnrcHeeIPb/
xfsYs+wOpv1ZcXokmik5dXrt0ASq1fe0ojrc/Q4OKcYH/7j90sHm69zdKIUh
sRYoc7E+G/RNrSoac7iu/HdJQSqL7toivz6CZEB6HUqsNDJmUF+n5mbr3vwz
75rlR7sZjax+5pEjK7coPMvmINckNn/kJ8cUnkFgF4BaFDR0mpfrC9Xw8Z3C
Md+xp3x+jSjzRrb9PgtuPf/Iw3xGJdPfzO5u7GwZXPudvvEwvdLrH9D8xfqs
8/QjUV7A/UMQIQm3+jl2ZWzRswUfshe/clM8HoV4OR8vG9cbG4Pv0B03t7B5
i7swBTtw4l/uHklS0aaSxD25u1DhUCyWbbOKLWeQv/zkesqaPxFeKvo25ocK
A+59r3kLpck79DePsnS9sZIlFZmxx/t/LmXdbpF5ImgdjQ3stWpfdXB5nJ4r
UigRdc9vx1p9f9YwH/3wZVlZVJq4EMRndjxArS6acXK3eqHfKi0XUGr4itYC
FdsUxVFYRt2+3cMVy1oXYnv25end5WzBSsCF1NPlWV9kSOnY99/l+Q6oATXe
mv6M3vT21zFpqSZ4IpnURM0ikhPMfANlnKXgPjPbBru1XajnHszYuX3DIyfK
YaNKVT4NrUPH3EmTuTn4lV3SmcivESklAeKCbW2ipmLG74wBydcMtqp9Vqxm
1TyOogIJet1WCIuXBSNTmRSQyvRwPfAaNxgBzClZT6+tP8P1LVtRvtxdS1l5
N8PD7EHCKD5SLTTfjPfEZ8ZJP+FcJAD37AZaiW4ViL2T3F+GnP0Bk6HvrhUb
PHO9OCIByzkd3bsPhTAYyEbupGosZG0vC4nWHM9qId8dqgvgGHhgHBMnhJzX
nmUatLuGbilv2UxEicdSB/Ri6q+QW7Pzt/VO8D305W14w6k+WlU9ZwtCqKEc
2juVAjQt/7nAWWBO+zSndMUvV/W/3wyP0tqx5lUBXrv+s69UKtwdUZxaa3wR
6e0KJpOVQPHaXXU12VLJ/x4CZ2T2PikyKlBeIhNpWTqIUl943pBf/hwiLI0F
wwiCSmcyjH2jLxFU6klZCjMc2hFTMnCg/pskPL1S0SR2EmfFeSkJ58I9BiMQ
zJNEY6TnaforWl/Ta19E8yuz1XfnSzrw6jx2k0FBCqKUHr+ksbc/ioW0hgoD
g2ATrqtzjjdTztd0v36MoYplqOLW5czVXOgQ3s7LivdQ7lWMmSWS1cFVanPI
9QCxwSwHmAj1mnjY0xbAAltGJEaupVkiIYStmNf4cq8q2dcXY9zk581iDyAS
JE1sLLq/WjCIoe0EmuZMBx1tG+i/5aLFECfoIcF+WPHM2Y4NBkAZDduGBKR6
w/tVaOZ/ivuScLm8d83kb3CUn+9kymzkoWJhT7bsxzUkDrxTfbfOaEt4Uqlf
bS1ain07udVwWyk8E0eLtntbuXmh/bDDIVRzJOeVu/5g4U5mt+WK0oXasCKH
krJyV9LackG3HBXHOG9iw4i/xa/K9C5Lb5ygRsgtpA5OEvHuV/jqfUhoVINT
whpYM/pVJCK6OrOjZMH2qsEIRORuHldiF3iZJWaD30jKNa8v5XgEB+ROIxs/
AHmspxjp3enXPqIjyr0RRBvTWFx+aUe8IJmIjfQGg3ouV7qiznF//f8SyNAr
YOM7ZI9TetmMoli4YdBsAaobMshlLnLi7WEq9VJkgzVVjrgZjLJ4LaQX0Pgr
KHAUpWyvkKNBnrSpFpYjm4t+6MulKwq3ihjsouofud4WMDEZf2WNCsCcnZiT
3RGKmn2EfiTZjzYoW7mxLYbAS3sogq2G8bRy3AQ+jcfStC+RdmxPd9cecY1n
PAeizQqvNdXHZUZGOZjVCAv/6f0MR2OrDDVMfIZ1ePFX/CnvLPH4HtA/glct
v6fzBLVZQJKp2off3GlFzggZL0GROU2FlZBV5QWGWwPWAdWq5oadaT4G00Wu
/Cwobx/7M7IiwMbTRxSUkbluEJnMHmaatkIxACKO2Vm2PaFr/yv2tzZ7Y0TQ
ED6iFlWEdkXXz44Xf4oLv6jXuokYNqw5ODuuIgOk2r/uOxZrDawGXPn8s4KQ
5EYjyEXUx8doZZMwdCkrExCNf84RoWiMolyVLZlo84fG3E2g4ApOrGG0n4zG
Wuw+b3i2dKHfS0vMbnMm8UUY3Wf8tyGHCJbyFglZEcRGENjYPmovc5VULa15
QhbI8crqsq1D2nJ6MKyaUYwl56VSGVJ3AWu//7f+mP2zFbLkTWLmHYBsPmg2
2A+4Kd+8erGRV3LrE3XNi3IlTyqT4mSjFPAmics26T4QskGW/Wg/KP421duZ
pBcJh/B6j8VEiFzKhHekvfc4q52YJIO4WZPC1bV4dheBx4X9rQIpXVmQPJd0
zyypHWuPHjOtn5tIq6HhpIFtfemQgbzersfq0ufp0TvACo/+5RKjoh1fm3/S
iIaWZfBo7onpOchohrf75GmJYabsvx1G4A/oUNKR93CS0ukNUpk665ksppGA
mCdbm55DcoGiDDZdl0K2oDRxiSJ0QkTm7IpyVwnHy6pRUjXWx1uj/y+ipPM2
Kv/AuUT1M4oPtUJl89TQlNr7KlBNpCIqX3mR06+ssNgYloztXnKSDhp918h4
tMVXIGgIeXDW+BkPWijJGJw6Dp90u7Mx1L+WTnKLqGPvfhXd6FXBndKJHJBo
zt/9uNGk+3m6E2f41ohM686agIyhRjbXYqtij8nOI56pWI8JDcmKJC31rsvF
7XYF0ruA7DTPQ42jAbzz4apZ5cX2wfAhy5AQ5QeOFmbqNs+dTeynuAxi6F3/
PvcTZYcikeezvRrj5sCdJzgn6iEThf6fuNnB+DnLL4jQxQ2eLwPBB9nYwtNT
8UMJvRUUMUIr4RTskzQf2QHJwyYvG7xFrjrfUpeH53shyFf1dVDa7ghAU8he
m73TMseyuJpMY/U35FDqRqBiOMeNKSAz8LlXSF6W9QdHzcxSsWGnrd2joTPh
X2V5ss2jfpplNeuPyK/4nJSWm8zvo9rISpcAl0pbBY+iHFNyvYAa86C+UoIt
btw2JZ6Q7OddC0d8VxMhl57XxfNVGpaCLK1wIifneZfRVeueW3hnCquFodDe
5+HWHK2rKwEO5w9/Qne0XeS29GDwZ33i+AuA09aJM3qNOOQaNvotaX4ktDMY
37AUPCi6sKdM+auTtsycdISXQPPasvg5yz0kLWsJGuPApaY29Gp1JUFAowl/
nn9gYHfiQXtJGmQ86WwhsHEUDP8II+x6nu3rf6Tlee0Jnu0sPvlGwko7iWDO
8d+2sREX8eDNAUhEVtnKz0alWaUM+eFbqXhldkav3Hw9KpOlsYqk+mL88jBQ
/gxv8u4RIx9YRbBUbDYLeLiX+U3uA6kEmbK970z6UnWNpclukbQQqktqjWNn
xcD1EQTBwzhiqD6lJ8AOnZoh4Sjb5jzzjm39K+j8OkT9ux8GsknT7iyhGM+f
VaRdTlDLfZX5k5AKvTQZXinjLzqsdmNnpyiWD3KJ1WicHtYBB+Wulz2JmdUD
f7652HLWMnClix3djAcI00bDq/4pSU1VwyK6YtaK7Gy5N8bhm2S4TVMYBppi
xT0kyJeFQl4rLV0e4XPYuS6ujy7Gjt9J/DX9ANEyg48Uk9dwk3kh5CcojdGI
+LIwWEXb9xMbI1rF5JWDlcsia0b2DYWVgOoUbuvxwjwD2oTMFvztaIhLyn4C
WAq1DCuaJEwkZrI5doq2Qt1ut0wyYjsYVQgAPH1PMJAoIQKDSeI4Iu4rEYV1
cIOKhpIWpdnS0hZkLu0RkV1kvqAH6YU4IZ9+gJ/Ezn4THe03tR/FUXc/iLvt
tJTHHMm1ARxqCFd5BZuVHAmnD+dXCYyRnC0Py0wBEexEC++E7gdpfWd7HaKQ
vtzBDvYP5WHC8konW0CIkjc9OV1cDePRwyeN60he5tK+AUGHr4g3LNHBSorw
HeoXhTBXDsTVDTBNQdsJX01wwfQx3xnBR5ijQ0sdloTALvEbiUBG1c/3u59X
ssDJ/pkH1BaZM5QEvnzK5sYAyHnJR2aIiaIe+y/XUvlY1+1vkEGeyVPZk70S
wA7raynz562M+1UoY68f0HB0FfAIypgREYLVKMhs+PcUS/9JBUx/ER6ddEtV
bS9HFkhdrXF6H208PT07QZ1eKpr/m3Z2gzRX97E9WwV0j2GHTuBUYL32TLQB
HA2ndcWZcseBI/Au4nKedum+rMkmtKuVV+xBCAvp7ai4yk5wDGNnM1WOA1iW
EZaSf0MHDFj4pWwlut5lU1Y5WTNICoFeFAjx1ub//GqGcNBDed7Hwpd4nibL
hLWPF75siQHJAtbvWCn025svVYAbmkC0MbrezxY4aaqsq3NT6miBg9sDD2Tn
Gm7KYdTMLRvENKwJAgnLAf69TFt9QN5qipWMH23X/KOEa0P1a/uIzshp8NFx
2zOrGAcfSPwMf0p5Zv72WHOjrlztBITyVlxvWnUJ5vJGexYtlh8xS7RzJQh2
7m+QKi1bEXrf9274m/Y4EgG3dCEgEpwIWycOVKaU+deAMclRwNFeVL6Ha2Tl
vGRHnNU3gAJX6iIq/htE1g9LbE33ZsNd/9vg6vjr8lVzoHQKA92ECS3dpsrj
jTkgCthGYDkChycGi+SfdadLyodhqeV/BJE6guyHAO9yrdOt8ZHhga2qAwhF
5mrP4SdcgLiUgxrchguostu9cn1Zi7yHwW1YFNjsiSgjldY2KgQPv609N6gl
t2gvr93WLIQHEPUgmca1vGBQU+JRLIJiOj4e8393dlQme8lWd9Krx9Z8PHij
P9pqE7iBlrvkX98AUojznEAYFeE3pmeFCKSoGc3vattt+nS8LOTcCEf59I9t
X9C7x6KXpEOBXkYOXKW41v49HuX7KM3tfExY65jgJ9gthZ7Neo9lCcwbYQDi
qXIW5EoO+XI7oTml1GfTugh+7e0NzKZubhiEnaqoOAaUEkLl0ZonECx3kM3f
Td9PEIlpEkLr+XzrNS75RcbbL1oKgDQkPrOe6SYU/Ldvy1thz3tXUfdI4/A4
1ZMykxOy2wHPDcO1hrznXCGd6e07KhOi3xz41l6qkOOULsLq5/WbvPfebKpk
OkrBDtT9Ycq1yy6DkAMpgt7+lm+4qzV6dGW/5ExrZkLeLvajawUG0AlPMlIq
rrz1gFZzrdxMcqHc8GUD0n/r2VEfG0TKygOoswXIc5KcYeOurBFzu53KiV2S
K8lxq7KdkYLPkeDiDzlfagjXWHJZHq2ztw7Tj/PHqxx+gF9a0ETQIMrsgGnG
YXuoXLG4Ulj2Zvn2V6y7WSbpQwclcZaZQaS2FKE0ffsZ2ZOoZ565HfVVsqxG
PyIyiMYB6uQwE3ZGcsemt6mg+RMQndpl7zpJiTwGWjBhbL7oB+pRwGxd349q
PQfUNALHY4cDyd5TSuzGz6tZEoRJNsuwbpGWfcRSLf9cCHcLcLvGbVCMYtYB
pnie4CwhulvYC7buuHdTBWMsXtV0OMkWSGnaDLFU8LWxM3vcHoaOh9wgbNkY
g9PAax/ykxc92WE0oVrlpL86BLYmOIVbONuNNGa9uGigYGO40GEhJ2TSFtK3
ctiLMXTXG4vgDxh0T9pxIqlOdDMANlsUl7mwrdlmgHutv9hZ/Y8OyNzYJB4O
EQztlm8X7HyCKRh3OARkLxPsqxkE4hZgKRkqwM8cKYX12eHnYLIefDppdNXU
DoGFew5afEM2QqxdppO7wtVeuO/k3Qu0YWT9bSP1uAeQNFzFMnCbH1OwK2Nx
UrRhkr+FikE8K8ZaBUMHGH8reLIyxWUEbTf9P2P9gU6RIPvRJRQmHeoWCWuu
Y19lmdCe+35nfiWfvsHBlTumvgcoCCk/g1SFgS6jiebojsboNL1RbbhOPhlw
CGFt6QnRb4V7nlm1wCKbgT+GieUpx7SykT7cR6gR2kkMfMOXQ2acvMXwDmDr
82rAh24Q1Ubqg6+LYdB9qnJoIg+gC+1T8jWF0Wmo1YWM8rxrN5Rgr5N1RNr/
Rg+I/ltkl4skjuoFUYdUVCRJ4R6pR2anluEb/hhD1DtoVpEbkmNvGMS0SI6j
XvKIeWOEHhSNrBfY9ItYsUz0/hfh46rFvaaNSIyi5vC/TB9qrjxWupV6oFMJ
LZlAOlnLQaMHAcLeoxqaVtb3pK1AsYZTQHi6C+VTwsTZXuxgf1ueJJZEDVNa
gknW7COxVH8E1Sy5hBm+YxyqxcMYAJ73XrboI33wzWhoQ5qFX8cyzlIaV+s6
6HRFC5Y0lavDxmI+kFuBx0E2LO5NdMMJSPadBXthGRucebWBnsOZklkS+wuU
EO9BpVXJIjnvW593iJ6H4imvs7hgihhYe0Cl/wRatseW5eUQy0RlYFY1UGB/
iDEcmFus8qNX8xTI2CLGccT1cH1eJsPYwiWx9Rrm2RMTUjAWE6umX/Nsr1p7
/P8oceRWEG/90ueGVKB8YQ7fmwtJ6sR2rDX6sPAYjqz8YntgRNRDCaM+1jVk
xlmhKL8Tjx9/vDra++JBpWjkX2IJjnyOFyslIu8E3gU7Im8OEJWu6sil2/Dd
Q8Q30bi3zOLIfkiVZDOxmM5ReJ+g3i96zB8ZqmksPujAkYKE5EnLzcsntfB8
tW68HUW6ZKi1uP82q/NLGchtsNO+32WwK9H3ZNnG5X+f2Gf7rfuMDupHKBec
0Sq9DRlL6LQxM5gKPnOaL7BNcY4vktRz7+307oOa01gSI24iHGIx4T92kjU9
Q7nQIkZX0zkW8JJTEA+p78Qoa1d9J1ezbWQHzmcywOikZKCXUtqnfIL0RrUV
s7HhszT/qYs94YSbD0S+falIfIHHPiUnA7R3Sapnu9f1Ntqfgc++frfqGzom
KwqFA6nIXRxv+j1cMjksgxj/y8E53zNt87t/oLC9JQgYIvfP5y/CBJgHGMcf
8hfBQk1NJWHXeFVuHs1CiNVtS2GeBgVxq4Z9sLnXQ4lp6uWwvLoMikd0658S
dlVVouabD+qHMFu1u/ptrTrCl6MhSYVX19Lcj1+3Ewfxv7XbV0ZHVRBVcit7
5oHhuCUu/B9TpPLszsgofMoN6JhN45SQ7sgwnPzzEFwaN6CHDQP6dgCRcwd/
BybG7RI33n3lHSAMmpwdWXRhgtmx44p06RhVcecW+vp0IYVDl8sGvemj7/uf
M+SDt9wV7+/X8CTbr7dcCQzZ7e9ZCtnb6pNr8qsxcBytjiiA0+OEfZ5Snk4z
rq7Q/c492FJ0BJvZ6SDaUQG3DNdeM3e+Sp7UZtDMlHMMbImBrlq8x1tFIgRW
75iaqHFEcPbHXbLmRbywtZNp7sB082Bv1MQNKunU/UnxKarTsoRLCCEaloTT
3P3KC9aycKUOI2xRs+96AChCCTt3Pj8BZjaZRRdyXOgsa8k0uOhR9emIy9V+
GlgEJxQCDS+dXEIqXUec5mwvRzMmg9UgzsJsZOvHvZtl4lPcpf4pI5toI0PP
NG/eOdrNOMAe7D8HU5vdyB51V4B7mYTuI5WAvfuQ9U+ZEpSdUUn0C+tWwfVe
3NvJz+oaXuFXUfxflQsGw5oRqBFMWOtMBY+UPPD++MuNQu35eXoq7X7754Fx
PjpU6wvAky+EZC+FUsEgrvfWV95WjzwirX9rVh7wcgP23S4f2Z2jwx8XgZ1Z
6DpCaXSg/Vwdl+Sv7Q9G02UZtAWTYSdlq2unOamusOolfB+rpLkUfiocHkBP
hWBZSx5wgUXuUDict2LzZOObYxXAlqhJ/SMWLX7Rqy/JAnbHu3erKxwopNCh
+IHiwgHp+qgm4MrOQ74FjaMqrTiI0xR/C64dOoKo/FBDrF46+lf7JDaQ9Sk/
ZOWCv/WXnUCRIh0yMDpJmROT6O5d3+yyvy6mnGUm4DqzGMWHvqhP6yb8MZK4
sE4r/SJoPCZp4+qOM3WpkYdlr+Uja2GSMCvlZR8cju3rA7l4gjzETRHrRODh
jynVXBK0Ue0+JQNhashF8YBGhGrDRmWPLb3UAtHEXWM0ifOx1jE6PLEmhCUB
l3XR5U7IaA46GL3v7i1cH8VIXS0umZhKUxgBGWvrhV0VzMCTDzmuLhRs6GcO
zDqGDSodVza1iiKqs7QBn/PEre9TZ5aRfBdTJvh7i8zQmiLAkxZBHpRYuo50
G3FojjPV8iJXwBUs7f6xAIpcFIMD2utkHHeCXNjUoS8ZjMiDkLluHk6mHoPY
NngDyprjd1hWK3cEDYI2cOysoouP/8wfgb2DuWpNDXDXDEoCSkSf3LqyS0cH
gntHqvjMg1kEx72BYkKJ25a7uPk/hgNpuzNcC3TBaip1/fZ3vlmCxSZ6qhFI
zmN7P0+zgzfQA4dMrYHTiOD2rv6sP9QMQJoIhDLD1RphqxOq4A7CK1Mc8JCA
nlZTl1FyXItio7sUmUiFudc8OBaUdPq7RzpBiEilZcFXWE16iCAk4TfNB2XY
iKp7E/KNuBOBXOb2XePphi8SAXewL+Mx+VrfHaH5Tk11vOClREEr/asADEas
GRXAWxrF3YJFOlj0IP3lDLdk1crm8PBe2x7O6NDPYLCEJKVU6Ew5KXVpzvix
a96xpuFt+0xUHCfGFb80MNMe4hPGrtDSLLaayB+k9ymUo4lLh/agqf27zcc8
KUQ+W+net+EAijtuX6ZsyPMctKljGZfZPwSgmuPDCCA/vJ8yzdaDlIGx0aCk
r/z4emM+jL0Mwkl0XevSxCB8Oi9r+KAsaAC+LbOB7HuVAyliAmX2PjnIa8Ge
4gFmmkiVrRzVxMcLu9aUQNw5srth4HasxtAA0WUONE/coeorNjAeeIapBVsv
eGU8oE654CexrGDTuf3r2HFqAbW5e8+jFTSGQlaIc/LaAz9C0wd+T204OGvL
tcaNI+bhD4xhTDaXmJRO8Xlq3GDgUzzIsk7+SfwNY7yRf+wlFsD8cz5lcur4
mZMEAPzCoz4KyT5E13hMeNwYDjHEf/GpkfVU0bXzMBM6VLu0//3zICwUV4+k
/YRkjS8mM4r0gRXwuaf7k6PmNnZ6iBRRL4fVrYttAK9kCJ+wdx0xE6klc5Pp
ksLzpzGuB2cjq3pISuwzbTWev9GIACV1O8bY7s6M2ifwh6VnWjOz6H0UNQ7I
MlpfUOu5dgM4axr8ETYryWTbhtK1zRvcOwPZQMa9u/f5dGRRF/+/6PzqSvLe
sXV3FiH167B4DdR8wuezxFqc+dMbOOW6INZNjEs2c9T/x+pUUVW2XP2T1bBR
VTtixZmK6gZsw/LG31pZdDrUtCdOSeGIi67OVb5nJeu882T+8y3b8nnOV1Ya
2wMh7tUrKJthywGPgLSWMpSImxKjwPA7F3lCIBaqtS2uKD4M7dLJTgbiHnpt
kArjfk78uE6vewAph2y6VCfqfmSqK+QWwiJzUEifsu7JMYd4YfX6XNGjT30z
Fvj3/JyVHIsXTkNjI5jJSyVzK8G/C7r2OaMFYv+VoTAKV943MAbX+BLokOUM
JD6oBgrQwFETS3cjRkOhpMauFQNKkDwMDkWsMT6yGj7otqyvHvqBMGykWTae
tAc/jSs96J8ftbz/Kent5TVXlNG6bBbeowMkNWj9meHPaPJ93l2vmYa+PWYn
LMPZ01mCBHpCGxKej0KnX+hDitsYfvgwficL37GxifqqCrZ3aC7wtJyJ41Zj
Go7m578oh5R7cpay94Ofqn+3oBeDRVno9v4A2LXefCF1WCj0vxM9PVSDNy23
Xp06N7Q/WGpsW1ynErM9Dx9OFYYv7FK4OtBCYWVZGVd12PJyTcNAzp8tI/OQ
Yy1VWSdogD73PARfllw2y1H4pwZStKIYTHeAEYWquCXvM3qxkR3tThRw24mI
fsmUBYpE+fYgbJyVX8XecGBJW294KRRZIFLx8ZehemJuqSs9K56z/r1FIV97
8W9rZxt2oIxbhq3CgjzZ8dMgRxb15BohZmW0RH4cYvBWV9JlWjnp6rW1KuET
3PonIT/AI1vQYcR9VDZw3+mV+/5JEybfMPO2IUpDl+l5JMNX9DHl8kNeRa0h
vYMDk7DBfJlpiWdrPcMB5hJzS6vNVW/GGGiZ9H1Lqt7eDdpwtAMkdq5jUkbD
66eW18LiPxUMwAuHVheVdIvTJ5pB93+V9KW28EGcSoO01kS6y2yJbxRdHw0I
t47ZRTxXlJX1tgs9UZgBCzZd+s2BjHHflbnhqQzbvgf2Jkfut/uB+rfYAc73
ctmbZmXgWla0gBlIwYoN58yDZ1xLeJrpmL1yvAcmhVE6uNJ6u8XN7aHtcc61
dv/r7cfNirSYgghLe8BHjAs5aL3S3LWdZoHXCiMlQ+EjVIe08XYRQXIkUtAv
jccFSuhlSqOQ2FdDozw4cbk9huFlNw+GCsdJAmiVB54FHgUyUvIRBJJG4OgW
nyYGhovDomUDhjPecbJHq/oe3YEnOe0t/vbrduKMbTM3FsOiBlusNJbGQF36
Udw+j2zEX7Jc3xp9zWJzhAFQt5um7937t7NGuIJZx0w/yGBXEqQ2A69BkX54
n4FOmYpV44Nu6wOzdKY3gjNQSatOxBN0mtefoqcnd1U1bAB6fqKCzbloQeAp
0bBFFWEmIs+go9oVE3HTwkOsaC8HNILqSwF4jLmfKuOAOR7ko7WyIwKIA7gA
ofhT8skHLxXEw/UK+LvFi+eWUbVv9ug4r004VibiGOw6r9/0+7q70FiIpXUd
eshIX6i+6DO0mGX7CZHDNkTFma8R7LFLSZCH7v3ZwaHzDuMATmFh+ZXWN7wz
iRpp4BJExYtyH0NVLqmv0LG9pU4FlZgoN/EkMSUL1t8NTHrwVKiFWhN1ZbdK
1i7NjqBndqQWBPTqQbpE71OLwGUTpEjJO3aUFeBLlLSgW0Vm4Il8iwVX3KGE
3xfWSmc2IuHeJ6jRWTYPiVV/oieJ+pdy4gsDlpSKsfOb4XeIqR2MP+zYoEyx
QjTaBAVGd5SpU2jx5YLtvnQlkU9kDEG0Tc/MKyNAN7m6146pOg1kCpkXc8ik
ArwknJRDjddhmI8kZ/8ZchlW9IsPrzMG8VQcBFr/Lzf9jQFA0BxRRT5J4hUM
olr9CG60NUZbaBqjogR/XBgLYQHNDjJSkBoTOkt7YMV4tCKfbostzfnJRx+v
umWfUVT/wnbMd8+a7mqnApUgtAqHAYHG51unvFRezaacMCT/pUfNxCrIE35E
NiyVEf65OCS9HKoCeVrKnJd2l98+UJ202ZrHSmuaPxrPQNTwxOIE9FaNPP90
Oeiik2IqvQ9ZS7aghKtUF1nJI/IccHX7Aml6yFsQe7C/eFYmKz+KZN7s/hc5
rwdv6EB3rkxxNpw0tdrXi+iQdnULxjHrJ/K1PBxYwcL5c0la7kX2hyAXE3o7
aYWE1hSFfVXsqGJ90h/UK3JbFh45vTq5HWnHKQx2SJTkl9UKnT8RqgLW2++S
0lPOK2Ps914X5tBJiyoackzCYn/mAfsxlYDLeYOJ6Z9+ri+cXjDoSm6dP7vu
ngiAHe+Wq6gnBZ3QLNjQ4etHG3pi/5m+dG/xx3mZ3JaFqPwmYGJdbrFTKzvB
ugXIUD2qCU7JvuTWlGXJGVMWLiEzkUfmL4Fh7Jnxd5FKC1FQqi/3sUpL+tKI
b6JzZsjYS1Io7BqzvSECI37wP9Inamr0vk3dH8X7Y5HBnOVdxdn3oQkKtcod
qJ1hp/iK+dtt6SR4whb74yVgMi7B492oGdkco9bK8yd8NlDjBi2AQJks+YAv
OHycQOVgApSaeVxDQubnPdJpfNweATfar2xb9Tphsz6nhJeYmgJDkOBFrYVU
aCJyORqMac5+QUUsvxs6BkDK5G2FkbqkEd5ss1HVNFW7KhyLaqcNaTIvvzTI
sq42QnzIZBDSRC11vDwk42gOjhFSKWnXwPjYQ+aFTJhwIt265ujekv2cIlCK
A8duR415XcRkoNNnPlcjXPWxq/Zfwy9u8ho3wPZqom8RpYdKvrGu2HGbE9w0
cKdfsNOnFYgSC0fGhTfI0fgDmVgl+5+DRQ7DprD5bKx/60h6RHfvq51pY1Fh
TcHiVej407Mzg7ajUxga58CpuA+U/xRk6p0l5rURBReRTrxxvCWo4bmIxhmF
+TZfCwrMebEUFczs1mqgfGkwICzQ8a6aHIly97Z9IH/MFfzzFBHGlUTeX1oG
0WDTxxAY056YAsnrmfsZoTzp0q5xdOv1AN/3KeKY5uZqJ8q/TWpy1tnxIDIm
jfgsa4cAxPu4X4gm/TVTgXzq2CuGSVkdwa1Oc3bRGAgVw8Byr53Y/e10m+XG
NrzJQkJFv57URRIZCIiRe8usZu2IDYxWVilb0oQ4L3ndK9dH1PZB4B6Leb7J
ynmzSL+R2kiy5XRtaUPGs9n3uZ2XjS0sU4WY3oXr+hgrcuo9k+l6VZgu6Qri
y4zAjesLxyNQ9tzaDZvsmekDbWxcBWt79WEpi0mWjz7Rm9jOWi3nGYNbZOWh
b1y3O4dcesQWzDkZv0tFASSKR0Ipdj4vYL8SEBoj85PWTWdKU2PaEfTyZ4Hl
ZIhQ8K3i2ljEztmmTHymvkS/bl6alW9qZEQij3FFQImV1ZlkO8mHBKNvAQrn
bcjhaG+U1SwhR+J5LqO7iR6kD59fZoE9xc6Yd2kF6WnizMOrWx0u56/SUPR2
UCgop6uRqMe+WWdQs3m8K7B68zV8AZ2S97O7ZD1r1v7kMvYr8GS0qVDRg2Kl
ykFMFd6Iqj0kTcAXQRodR7bMmndcn8NG6/JC3CooBhJP43vO8S7Pb3oXEQo6
gDc/vcpQw2jjZ3habG/icb94xm0yb2s17FlTznZZiFv3D5ycw71XuZFTcFbD
BlN3noFLO+BMQAB4cCQHT2aZFYsM5i0AJ2ddtsqY2MNkPUt//2ctHILUcJ02
copD+KCFB9/wHknKuHDMQwrcdD5s0AxQBjofsNLZNjROUUrnzQtIsGSPTXKz
MG6UwxnB4xA3cbPEJFkiKce6YB8jZZ6tlsONdLs4yDVUQWYCC865BozUiFLz
AYi8GUQV/PBynvCpvTU9IAdasRd3eDX2XpW6EQPjJKwvwwheSe6FqAgVEzq+
y2lyURSAYQFSg2yZ8t0gvoacRtLWQ8nmzLqYBtckC6ekHjv4evhS5ozxebde
Zj33JfzmuYvjtmbHCiDRRjzz3JnadmziICxl+5TKVhUmAPuzohfHKpNAW5V0
VMJ5m3VfNDALT9o6cIvB96/vaklQ7H8APsUzBtXiadoNcOYl63JcKblY8+ZF
NP13k7a5t+kOBF4X4ANchg8AaGQyGgGpDBXL7Eau8ZVp0eyilZrpz6BCwjox
c/osXWm2NewqilFdr04lTZqzpQzYeyajVS1ybf7g07DhlGNllI/oA8TSq6zh
a3kk65Ik/VBPYFIioRd4TjMapgghgxRk4tt8MYZtB+reOewXAzxPscBLgVTk
oJ4Harv8kMBnbiphGHeOilzvTVgBEmtBnrOIEn0sXcotEkBT+ceGJK6ZuwPe
4RiEpeMVPBk9owRyDTSOBRWd3yjGRwya4NrLwAKEh5wbsSwb/FNNjnhAGVmU
k0+fjC7VscmBGi+yD5H2xdrA+7LTCY1f+7VavKZQ7XTWMtL5QMIeWxMYUBik
TvzuRjceNB3WljizlK5Cyk7ER1pDCw3cWbVa3goIzxITP3Yn/Vdg7QtKw74c
RBO9YHYHKOvaZY3nH4VMjIcnjR6VgtyWPhw0GfXU0Q0Pv8wP3lCkV+LOIlQc
lsBPROB49lOu8bMoOjhsQ18A+Qln7NIR8wKsT6R/82c1/VFM476vzhkr7tk3
dUt55mXeBuHlxNk2XuS9N8L6J415VlmKiBQs3EAR0QQibAy9e2N31jvBj8VQ
B/GU0RRblrCWh6tL0VgN0hcJbVXRZPpN8ZRBsQX3sdCPDzYUheayeXzpaEWZ
JLo2cGqSwsQMiMKGg8h5TtHTPqNBAMNEZXoUVoWKkvKFGzdppVrIRBX2IpYU
0goLLgsYHl5zmWKLd2MXg2VaEjOkdo0CqME8/9g2WGHT3aw2GRIdfJQGpp76
WrbzuzAzB5KIIYsgUpp9dxBPcN4bPiwVSn1AnduwtliIyS8ui30oyjeSDZvW
udSaJGm4+/A//BrD2P/9mNtX676oVsrHNar2t+sgX0UK/4bbldQSct4gzVA3
bq74G86O/l+TKvB5ecMRM/miXYPsxvtiWrmQ+1zlhqDgBS0GQGbpqIxH9uJw
zPkjMTryHKdkL4dN3aBy0UgIkzbnooGZiLForu7MOgfBtQLZoEY1kToVXggz
miswdYYcMahn73/G72JDP7wc5ne6jKvK3COrEeUAm8PImHuk5NykAnDW2cTs
4BJm9H0VQH2ovCjkxv5eF5hoJKV6aKExyydwJaZsR3RR0++3LRsGlj5mEpiR
vlHGSIOQorX5GpS7Mwg2bHJlgpaRMVGjarhlArBBqL/JCKxSdb0rfmUnOdKK
M3RqdB/rM0kf3L937KV3GI4a4yxg7DeKIHkPnnyezn9HoLqDo3D+jUCREXrH
HFUszlCchLlwL1RSFqfOtktGXJgjPl7TsHLNAI+eAeGxZhcw3Y+NG7mTWdCr
6t3fUFRFPPWYHV9IrMQfQwV5M7UFfZXi/8RnV1OKWpABW4YckaRreT9NjGAD
BQGXztwXkKNTrK4KBIYoUlXMbY8OUyxXYd1B1xBbUdIA29eQMTidLNdb4rpR
cxEuZqeFR1pXZgZZaE9XxoXMpCSj3EpKaz7ksyDRVc+SeY0ax0mk4RvsRvgv
WBWu40urvERA3tVSseK/wuCuaX4lJJKfi6TyOjjTF+bUPprRpjRsN0HHKEww
qwo8xrcm8Z2BrlD1/tjF9M7oCHvLc82gXtSEFz8zXxNjdwH9g8nABH/KeFcw
7RmGjjg2yBDUASSIGHsIQx8lICysmks34+GtuJ9b2Vo5rraVHNCAyDrR/0I9
XSqUCNkLW7S9hglnilWGw0oLdbJCNEX5BJ8WGTWPf61/EBUviTVlPaha9wW5
9jUDax4l+iWT/rO57jSfsD7YZGTK7GncP7kHdl3rPB/uETiXq71B5ernK1Pg
eSH4GBOvB9WrG8SeMmNeX/LRNbT0U6V2fHu5G5fiEQphTpMxlQeUsC9uLBSA
U1J8YNJW3vbsRAFYjwJ6pPVaXVI8mInWBA7I1p43BZzK+EC4utxPZ6oR5tH4
M0W9oXLJinoEpuN5v9AbKjq2b4Q1M1mC4Aty7x/qCo8yh74zyYHvrivQmvGg
VQfhNz3h/I21QDVo1pGjT2T42TAO2ntHJKWf7rj0D85E70tat2GFICLbkpoq
MHjvc7B0jikp4JSPx8RsJdi/SkxCZu5SUwk/Bup9EOpIoQ+u2SvgxRcoYZuO
sAxUeLPPT+tlLEyt7tHv/UTE5SlrEVt5WntVRq53LQZl4ro4mFJ6e/fw8EmM
i6KeWVvexo33BqFtrNHAPMSbTowNvgpBEjsQHsHsgCINM2c6c50ymrnPKXk6
260/edygRJt8tV/BTfcOphx6ZyKcpQb8c8llEMFTNMTh0mcsHxV+t56cTbVk
o4yTOAszacpuk9nA5aaxYvXCex4Udq/TAw/xWVRHTXb9+G3A1RdfGu8/7nOO
nr2H9m8Yi0+pz/Y5pFfSMnP28QMbicPFyL+0eyWaI6C9mLQ1j36trFe1Z6Y8
6r3e/VBAvzOJGnHBONz+Z4p7uAqKmw+jIC8xNbEzJbRfAnkOhFaZUFf7ItTx
O9TUA5J3uq7esKLzyS2RePXLPYD3q4FB2p2HinKdOdcivZu1TfgbF1xtHO5O
ICufqwnf8kviAbHrCROGHaY/txTzG+v3uLlg1Qe1UfLn0cramDY6N0pjnrh0
XiDJwYGYqqAuTVmgM9y59vlTeYvawJS0+kT9NJLMQCOBrmimdVyifRAeDij5
dmXfCgKKju31hElee2AbbfIZR/T6+/thc9o4mP6hRuBPIgwTF/vMwSonMGNW
UnnemAAQYegsAY5B1F/CtGSvYMY748peU7gzRNDIFl0SdVvHeNvwHxJEVHCr
FvggA4VBA0xls9FVctsDrXSMFv1ULyLK0cJvdzpuaJrxguVewVI3Up1cxWPa
ZobsMRsEF9SrXMZMyjj1wHjGRfcLjh9msx5WCM25bEnvxPQ57TfpjjOLlbZl
fYtsVq45MjsvWGjjuKhMGoWi3lnjm9lSGAw9Ao0WBaFlBwhNtKl8D5Ls4jlb
zJrtTKSiiJk1l9YeYWlyxmOUBz5TL+Ej+gqibyYI9TaKZP+4HmdDZY+OP+SQ
6h4HW0nn4/9xJ7Ygwwc5t1czJHml+uI5W5SqznQN59Osl2Nw9gyyRxYdrawi
sSHhrduxdaMUBbjOhrjb+n6wQaQBShBChYQRL0goNY4SbnNrY9/x7vF1WAX7
tZdRV8oyuUdjZo5oH846Kpwpxf0JzsbsHXKRwPPa010x4fX5KI91h7catRGt
W2bYBh7IuV56FbLQ3aSWfQCbk8f+tAWUHWmSgKD6WJYgYpp8NNyeJSNvpvzp
P8XuJSkKF4/u+XYyrjWdLenoi9rQ9/8wY1E2v1fhdu8phy5pB2j7mdZWdbmM
34XOMtXapAtAfcpW9bKI6sqYY0aO3VqBaV4vxUP467vdjertHTbui4HF9f0D
dJPobXptklFhnHAW9xq8ugDJaKS526fe3RP5HZk0S8el58b893xL/CBXpi4L
GI8YlpsVXoCqeiTP5w5cKqLLWcnZy8CWBQ7EtPMVoqgaZozK8xRD3oKqKNn/
ttR4ez+iGRX7KHRH8+/lz8ysGNXdKiY4MJgR2pCd3UAGHucS2oQutUsjAjvr
8a1RhPkXYqlGzJ+a2/TOfvuhF3K4jX41mqrioTY+6ivzRiFPIe8XeEN1dbeL
KPc0E3dcW2Xdaxoqd70i3DSX1t5kh8om86H8v0O0SMW2ww3mN8Bx/rAMinJu
W+lz7mxLgwyTbcNcbOA/Z6rijgSpZbmJsQmut35Xw0Nn6STEV1vT70cZMVmS
fp9GacSxYMnjAI36Xo9Ffgqausv62bjm+1Jz+wDXfUm9Dz375QSjh4VIdAAF
RS8TxBxRQUal8tWyFjyVYWw5Ury4G3Li45ygWFLTPp2reBGqIH36pQDoMHDk
/548nmlV0wOzCIBAuo47A5898X6saM14AFqDFONW0DaC5lWScTUmTke/v1ei
bF3dkC6zd0G3sLbvjvNMQmTGIu9DTAL6ZYBqnG3QqWSANGyuNt9YJ00o7Rer
k91sZfJKlXLWxPOoa88XrGLPnIZnO6Ejn9icMHUL2ffjyGH1dnMCfngkLIRX
ZlwEaVXyZsFTdkWzEMukuqcFykjd82ruMm4xKf5On+S3aW+djDEC2M4Isyt2
qjroCmMnhsK6oP7vDlXNpFmJjDBDdSlWU+CO4bi1mvgotk+nGvL6G0R4Gd5+
YrGx8pyARwxvM8K/IYNMGM2f26iixN8MoGM9R0Nsm6OTFQkCXFuFzqm6L2zT
uqGwuW8Rekp2zjgFWHqAYtf7OQJnofBs3LsstJma5LKrkt/J4p1ccgKO1zBx
jkq3ew9cAZldvshUkbnfJ7kIfRxeFnKz5hz6kZ7EgfX6wgK/Y5ePsjIsSIQW
p/pjpwPsJoBzTMd79hvAa6I/YrwxJqY9056y1r53IkKPUhxOXCX9k1HNLJzW
8yOn67D1yv3jxcHrjU1guMg37/j0x7fbTdxRs51aXRLenkB3UAm3XNsXd+ju
D155dOThBFMChr36rxwjRYjPQ476FQxUDuXMSn3uHUwCF7ieDjVAr84No6gV
2qspcizifBpLIlai2N9uI4/RPrsz5cMCDWatkeZ2ArxJ1Skh7mPArdiwx/RB
VnI3g2/fGfrjtg+6irnfkIvHyY87JHDDzYXa0sHZa2m4BA3DvUjUItUrR1jF
L5QB/TkwqcVTBLWW2WudOt+xMHH71bZ2LAWCv6akBNoejnptU2Xl+M3a0o/M
7mm5FinVP/FmGRFfWYOXZfr5y0GvaE8Ogf+7omvGAcJDFak38FqPD8NeUzH2
wxAe8Db9ZCDqKrKB0m6x8hUn71R1w71O8kOn6WZTG6jUiPWkaFLMy1BeOjzS
nLxSGqEgCBMHKvFdGNW++gVQgv+cWqowtZDYBrow7hkmNXOgTYNR87ha2bMK
duib/pESYEK7OF4f3Y1hJileOlNPNbEW/+lCEk8lJU/KLA3DNEE60sBLQSlU
vvh9P6uxy86taVMzBEWOgutKiC61/xWUqrijoASnu1290SzJa0QvYYx3E82D
TF1qVZaig1+b1iwkwXa81MyJIgmson1d0UAvSuNQxFMd556xVMC2dzfJAp/Q
CiYsTt2g30nZ74lqMrlvXPXJ++q6TqrIdZ9wXiQ7stywGx2mSgu2GmX7BOs/
hy/vkjdeayo2b6YevEbMqT4lRohrMjM5XuGAMAPePA5RNS6CFLJpcfFiTv/1
ssRm3uIuxldiAugZD6kmZy7/rnba0JKHUH4aBKhHEZGImReNuF9kdBclzsFO
VBdKsrlkfr5e2KCyC7gh3W+1r5ajOeQ4DMM0j8lIc2PFGHHPKpJUgpT77wvH
tUK8CXlgofOP7kPaFq80ZVgi3NvFGPCz4VnDJNt6X+Oaqz3uziht3zHrhyWu
iuZLZl0ufOIghBkqZ6a9w8fscj20dHtVAbP8E0FO43IDv3qs90V8vZq4Lzl3
uBkDGtjB18WymfbbrPWskqFrx49yn5HgFvsMcc3fvz5t2MBeB1JAQmZd1Sy5
ojtthsQI3UgEGrNFplls2cbmAWHQNqCuTeQKwp8x33punr/lIxsHoKNu7kcU
n9xG3qyHtEpCITMGz+8ucm+GsFHcG6deZy8/fT/CAkkTzzlwPLiYoNOwva+A
ZtAnLVytJXE/b7gyZq/gMWmOySOuvWN+ifnLaF4gsGsiWsAiaVHTTt9vzBlJ
OlbA+Z5Miygi4ys74UQR1iNTyIADICSw1/Dh7uiuwiBlU+VOJ6nihBQFbR+A
ZFQhd3vXJGywZmI1+LM1g98vOFq4ZaVNk5wdVMjQFyRhqYOa42QSsAmmDY/+
Q9KVq/vc3SWjWrxPKd+tnXPaQ9imi/19uGazkrtJ9y9dk48NRwO9EGeV3XQn
doX7oQNiYlzhsMLQ4kfwMvJ2kNp325dedD7AI5mlSlcxXWlxVFDVEwMUSIil
rV0o6EBuxG9ip9JvUShRsEABkefRiAUq6atBAwDNgzEGw3oe7JKEZdj1+1/c
7RWrX8uvlQ0MVGofntJTFRhmonOcSD1eFFLEa6EvvHBAJCwjF+x4Qo1lq0q7
JfgriDvSRdQ3wXH9mUKhhfQgxYIud+1ol0PxCxFDMTeuVzYw1Jf1cJoPAgT7
1ZIdjNtpXhv6TkA1zf98anU1DgMb3Js+xnCxS0bfX67thCTAqHI+Za4c0CGC
PoKMXxWyoYw9aA4QB2Z8VCwtOHAGtJY6LPSFuYoP3NinUnqMKFub399SI7ri
+iCjeVon3M9kbN7Gf+ZcU6fTbjQgoVDjmrm2k7BWKOplpfPytYPQ/boM5Ub+
UzKU4PdnFP/WmikhbS4qBfmkS6m8Zn1dfOXg2hSFhSuW9p+ENEzO/KKHgS5F
4VaRUbioBJY2nks0rIWOSnaUHMVAPFNCxDJ96bGRnb8GDWbLGV72sDg0VSs4
2AAzee+3DTowF9v0MkFire/GbB76QNEqkiRJzjTMABRwZrQ4Wy+vW1mFa0PM
2M8rxKs8fJZV2Wey1wwUoAMqYYhpnr9spC1qefqnikXGmfPgA3ljf5Rn1Sx5
w7hENGyGMX1GPzwQf9XZQQjx/rLL5LgOrH9GFlyC0Z6uJU+aSO+ErZHnV6JU
ZAzRSQ88fui8fjBr2dmjC6AbN1RSSEmfP/t26fv2uj+l8vTRbV/VjR/U0HRg
HeRIiQ85t1nKWoOd77pHv2KythGyIrthPBWmzS49sN27EmQGLpQsjPcmy2Cm
JnyIcn1SX2BMCfdOBbQYyP9sqCqrUGo7efhsHdnnqylEFUcefcqWLZSmseFe
LUL3yojLCapRvGCw+b7cZXAF0zsWozgYtA0Tiv5CU287FFV+DlAi1q6UX34o
pFrS06xQNsxcQdEvQIfPnIhglP4SqyN0rnA5REm3zo+MUbpTAGu5i/deZdAL
KuRQb5IA5hcJ9M2A4Ljjh55wdMFeQPYd+vs0B9sf01fdaT6wuhPSwQDE4oOj
UnQM23Ebcy4mHjjl9uJHlsiXoPljVLY2pUccnBKmKnYTz+6RjGWLK+1XTcXG
lGRp/QrHphHXAtfjqlWVq7tUJKrZD4gQPD4KpZkYvIu9QiXP3FDU0HSnUjGN
HiqMpTaQePvRNrrKg5zTsYRI/Ep6s8lN2Tlmso+3i5CHqOfJEbnNV0McOYH1
IUPYm25IKPvjhfbq8EoCzGELLICKMsdR5nVtX5fPOp4xASwOLXtX84qrDhhf
dOixA3i85Jvapjo6OmPjGXbON3bX77RuTz4byYFuhOBKAtW9xoGYSdUXRN2g
HfRgfx0AtJTcRSQgLBHYzgu3ucGtCNWnK8h3tJNbL5evBKyHh+CA8FPTpZS0
xPSJUbMMALIvaUMUvYEtaFT0wtbKhwBB7iDDqmlqJOkINVv2eZAEWv5C3/2f
FzmhF03t33duHhxelvem9tsVZk4IQGKRetXFfvRXdBaN7kZyWFodwis5wHJE
4ykKqDk2xIJjGC8dtt71l65YgfaEdtSP3TmlzwwE3vFIQmS36RLgzX7tzkh+
HpfBkXbAMoU5JJwlRVNrFfjxZX6SPaJYtKs6ffYcPcXqwrJkL5zUyedGlGPI
esBSkrfDyVqFD0zTCtSuTG30LnzNiZhiWK7KoI6G3WgyltSQMFJaWTkoawUK
gUvl8hjRtXcczQs+lzC36rnW6SLXaOCJq21AfyS27/tKLL20vftLJbOX9kot
roAXBA5Q57h7JqAS+F6QHXtVE4utULhgn/vmOV/ooYNH0AJKzktiDjzJdLg6
lVWHi/EOeFHlKz2zpX8nzMY5IMYX+zVuoEitIk+U1inG3vcP0kagUCHFarx/
r6U6yTEIJuEIUeCzNUXlIpoR+jTBbEBc4jNlWe2NfSkTdog0xRzeKG6qRMl7
e3CzAfUl6xWoOryUCbX20MNNB1sDoYp+ZScg64ApQIh6lP38S2vGxVvp4C0+
wbCYlXkfcyYxbz2GBpHF08VLqFvs/PzE4S/MVdenbNFUc0gj7LsjKDielgxH
F4CcOoEeYZH6T8FFfQkqCoyg4MZpMmr4NKPvlCHqqyO8ladqFMopxCfUSMsZ
kv468PlsXdq5324cCAkaJP9Y68siyWyapOaOtEqQZRBcr05BdpoFNKsAHXYV
VCUlgd+pxC9obWH+MqzU2va8xl9Pmung9Y2GTM+K7EdDd9jX8O0ieKjj6N5M
17vPpVbqiWgyETqwEqC6WD0EYiLJl42TXuu6ZG/9phJRZzF9SXprsXaouyg6
PjZl1vsSKlGECM1jO+8YEkHpNomDCztaJgETXcYKu8o6Y3+G/0jcNuId+lZ3
aZEbPuvFgoy6xQuCPPwHf6ZdqotwonCFs9siZgaFzRdD8QwnqHICVng13BX/
Nyh+nXsLeIQ0lUl73ph21vkynBEWAi11M8/7Vnz9HtV7r4d/isyVt/PgcRh9
nkhJanq1b22wk4drq3rh2oKhJPgGDnC2azHanWuFZqYh3wV+fEl6YwbkgZWR
ab1qho4cDbah3Hn7y+qP54TXus3sb62BPt5J+TT00ZGo+J+mes3PPovY8IYY
00tOM/Z2rQcc5hvHQQqI93QOHWsjErbuGDMn8UMX9hOBZCTFd7ITUMIzpCkK
gbyHQUmI+XKCs3NRcp96HrjCRbd9bKPqADK6gw0SYoB3OebbRc5V6I9SU7hJ
uZUXVCPAcSVE4UhWBgInZ3V/kEpJgYYFS5SmBZJJI3IiQJIqeztt1NLWgwwZ
RMd9JKvLzKMcSMhUwliv+Qw12TWmFH25cLP/mYioh1+MyvqQZVM4L/TG1YRE
hAvcd44oXDq3ZTDjqu7YXthA69VaxUa7a1BPzuZAbi8HTDmeLF7WqEX5FWLn
3h+rCqCeaLzksX6y/ZE64vfD5oyKW6si1dnY2olxdR9jeD/liSCe6yccA7cv
Szd8s60UManQt8NABO0pl3bW88IzpNE4aY7ETXoBlvZvCZ6X6QkCf7zEojMq
OlBxAGXpdW2I3yfWPUhPRgoSHXn06EIS7tksoUbAbGGzctq6BMIJnS5LwWtR
9YrMRNyBOH7RY2oI9OA6l4Nx7fpPCeNzYgRpOWY4ZLdvgl84NhT5M89FHe8c
NtYc3N0TAENkw/B72+s7NnCGx5UyS5c3lO1x7j86hEabcaoKXILML+S3+a+T
Xq2yGMVx+/YJiMthKBFfBNGAnZy98CHRjyq2cjUi2uXQ2m9TWbR73+GXJsYo
MSuA7Sn0/cvRxbZcGS0uCdLLSpdwMv9NiOmaMjmt/+yQesDks78L7rSbAmek
SylS96wF2ACiYhQg70U2Uj7GQxgwEPPRVGjPMIIXUCfs5DqVQ/aozccyGq9i
vjrCsn7gk1ghid4VlJjvYDTuUzS6gZZrAjRiyAwVmYhwIL8lWLsd/QklWyT0
QO+j0ddnPbjqqzwFIeGQSb+7H54p4FZW3Fhe/vUEj5Z4f1bkgIVGwCic/ksV
1p9Nb2YZiW3USZqizIIh8ZQkBUCTWVkFBW/bBEK8mJNVjKACfGAp34a1wD8e
7GMjmLtZZxPoPaJZjQ+7An00Pr8jXYHC8tPrlYddaW/1lz4aw/Giy5Dzdd2e
hrO0bo2cwbW6qFR16A4zGSbdIjWz1vGHX1nJlbPe3/lUfCL6/6G+gK48PLRx
pUAXfyvpr8QpmjwJ0VocrWwwSwKlwcOQ8Q3Ps1hMrAarSD71STD3xYUupz0q
fTPgX5xnrVNUykzb/0QiqMr64CMyfCMRVeKwBB1kuYSi8Kfk1eGyhoC/Xy0O
FRwzA1Nd/GXU5CfglJIlTCr1Kmy3079PkPTR7w1jjT0CBQkuWSgbyjj60oBB
/v+gMinzoFXx+ozRacGjikMd8ckViFwPmh9LNeVQoNEdq6LiNinXBR8MHNEa
MDsBQNzALs3JBfDAr/dviBagWuIXc3K0NkrPoQrrsRSftSdccn0AXYt1P2Cz
U5hxjc6br/e4rJMbPVdtrGo7xgEVrSFH14j/bBzuqvyEvkrdhAhIZLURdWdT
bRJxRPpO+qyHbyBty0MuyXgyny9aLtfMLm6NIF70bcsXyMaoRBFxgqqIbWrW
fZfIFj4PIgf9xnMvWBakljDTXXg0p5+QPSWGx+k1xuOno3oqlO/JHxCgMHWe
bh2F2/b8doC/UkzJwS3SXs1VLOuxuxzaSivbWIv/Fvp0CPACvfMSIJa7+k/9
j1nEaL4uhstgoM2iSrJh8OUG9mmN2+ebgBPoD2jTMm8fOt6kreHXkGKIJ8W6
VI4a/1yB3BxMrfko5ow1UX10B7csZlZMPQaVmTD2rVB0m9tNmdwGx7cb6Fcl
KOxH+E2PygkVJixoL1blyGwoca3JyHfTN4dIhJVBAj4we9xzPONIK7J5FBVH
+IA570m4G6KMwFXRnp9CZFnBibH/mLdpWSuzy+w+H8hJWxc6Yb/yboQASik1
bKFPKgc287srMUkpr4/DQngDlRDeFeabFkbgrUJgM0kf7JwF6hJXUWLK2vk1
MkK9O0vBD7zbjKz8WEXkI72SsUH8J/H9LnUEag0oVNVMI9NB084pCF6POcom
zM1dT+iwdbeHQNO1U2boC5gkyy3PEV8HiJLpkzekEgCxePWdEpk+V1izU2IC
XOflHVcYPiY0S3ZxMZTDhN2xobXlSbWGSUPLDm+AzJz7sPbHoEPr3Jb6/rSz
zzp4CkaCUCvW0lgFdKwBa9jErNrqoeJ0hcFlxW08Qg+ZtUiT23OPdNr6HOzg
XLp9YLjIMx68tPLjGYv5cZpFxjVXT8EpVOLXFaMqinsX7VSSnVBCUTsgAlPo
toVbrHcJBgxFn72FI0ydKNfM6pH9g+QiLrCsE1V/hKh5YVOJn2O3EL+fZJnF
RcD1Qh8P2EJSW8wvle5toliAcjcxBrfAK9d+AVtuawuDZvwEVIalaN7fZogg
kusz4DVmAF6MI/M8PbrnvgSC3rq8VxUxQF9NVa8fkI28jhavyqthBISADHOg
jDMyZzmrrJRYwMNwU1u5y6VXW8RcaorDLbr+QzHTSjEw0XwwoPr4DCg4xHCE
QERemvKdxL+iwGFZswq9SfiygDxDkK51K39dzukkURPnGb48dORNES37LtN6
Hr+/aJCO+f3dSXDqqGXmy0OAO5OHAVEuaA2JKizNkSDYLZJI0rAmVEYUxt/g
xc19hnnNJbiWm0tgPThpvbBhbjxDW51pOPMOx66yTYnfbLyQv/fEtEIZEnn+
K9oDGLfyBOP/xKqAH13Ygdft1GHYqv/7gjtcchL5OOK8+rMtsVfXPjZe7Fh9
1Aq72AN44VWIQUaxmOdBiorqSnvfsiCgi2vL+ustkw9qM34cST+hJ2EkHIGD
vKoP3PGajLVNIfG4wk9a5xlRmCrhG6JUPbmipJc2UtF6H3cc+rOyUj5s9JX4
sWFJNlEYyQWJtXppLM6dYlAhg6aHxq5dI76vsx09bhpevVuuVlqNuzAUWTyw
TbnFYURqjTETxEAFAxUvZo7AAuxCzVhHnVrkDl6VnpBl8E3cjgTTgZ6C0gp/
wsWKk4X1AHqEWCSwEvuTq9ZDMXQILJRcy3jcX0TPMo8i7eg0fGZEqQjh7iUm
HlHrkPIpwUw6GbFqxpqWWU3w/Wp9zS6lNE4eohKYGMQPLj3gNC960N90Q50g
qdbvb7sQ7y2L9YlzQ6eUFsxKY/WUK+HZ3DwpyBOjOtU2Haq5fsnzpAK4ix3n
XvpRaHrOQfJRoVCnwtBUvC0iTnerbVla+I0kxetWxcTGDnIA3golCKYpi+dK
onnw65xRTxBtCaTn1JJPXoLvq8DUvi0r3BTmuZhHlOc3Mz5KIFaQpOLkPQ1S
dXoOXDzhG5PIwkWLaFFNlGKasesnriCJrmhtVMmqWRTnMdkTwHbb7EtjNEvR
8S6Fu6NxQf3MA7GMc0H4yCisfwkLNBxQsb4rAVWOwSX0Y62lbOJHIQNgXBup
/1rvSWZ9WxeR4y08nYWlCOE3CWmsQ6DKW3PgQKWpPFIJ0IOJnGh08t7/Pv0Q
B4qMsj9/5f2QkFohQ4SjglPKZ3k01BXYSz4j52MUuNpsYEV/pZ3pE+ESFXXV
ldRtVfbQDav9OwLt5NL+U/rArUfx+/oOqpFP3/RpcThHc5c/2wkKBl9JpBG/
26eABB+lYxUth4n5t00KhfYKq2abHlKL+1eKi+DOVE4G79f/I0rR1ydwyRBC
XwW2qMFiKURt8ub73nOaI7/d3CtKjLS/e6QL8OXEsoVlrOocunRTzLTP/1Bx
SWQYix3fh27WglwJNIM2wbUbcY5awGJ0OpEIUYvsMjpFSPTccpDtWmeTMWam
JrwaBS91DOhNHEhodyP6rGBxzUL+SEm0OsWEGZy1E1YmTUR8yYv397cimToi
W9XsciQ9z90FX1klmgVf+6pE6NqWFn/QBmDqX2Re9gPaZB7dHA5xT8wPDKlC
7I+6YdPvW+LoQM+iP9auZt9lcL4libhgH57c+WDjcDjG68gPot23F41EAN3a
UlOebVK9A4TDZhcK2WG1zm/EXBAnxXBJX9AY/CxeWG9eJ8OAkv0ouOd3t5oL
sX63Y5oD2DDdPASod2eNL6jGPFTbezNRYJ4bFwCWDBG5KdxNvVpuXoKnNhxH
JiE+p1KnD0k/96jT22MMl2tHznwToVGG3p4iHol1WTRf8VVhiC4WbemmDV48
QbrXBq7OYaeoP+SjtArxczXvAbZGu3DH6mrPlcKW4qhILwDwU8f9umLADnND
pZn25+UKeFpjELlkjFeoM83ECb1D5V0gmYr7ZlJUHWiDCaunoumwYDcAUND+
CdLCjsARjpwTmcv7WdqoPputdjKcULsRKuiiQcSj2oBW40K21cu3xAff6aSM
5OJPAFWwCnHwqf3ue1HOaWLcoGMar72208nyDF7Jip6+4VHCkXjw3dopJzY9
tTqd3sasRhJxUVVWOEoTo5a9ia8137fjdaRgRVxAArO9zjiaWSs68M++cvS8
/O61ooW34jXmq5ENSXrBj7WKr3/NNrAAlfg5ZZLLLp+XnyhWd8cwDXPKrlfO
XamDz+PtjrZgWW++wjOiRs0q5KEiwGVLoTMmmugepfav1YOiPgtu0CRyZWj6
/TCsHoCdv0XdSimSNLQ5nyjBW/XapCneELk2Rez/9E9Z31bh/IfXmjcr+vz/
tqFO9vwF/v0x/rX17FVGNk2S8h9WtBKNcpHHKQRPqx91faUWo/BxkFGA28Uz
4YuS4FZyMchIzE1HvKKPggu25cAyP+Q+IxcrcrR8NutH/kN+jLRRP/i228AE
ynPyHKUx9qoV4YjqCDXmdktvwN1qtkOIm49D41DiMd7vQMqu3A5KCDPg3+6Z
1dpxcOI7l3dEb2GOysQaQg8IQcjfDMEPl0h9ZJQMIxkZdhLCwX+QuQsABDcT
QstdUAlZovjjT/qhzP0C63KI5d+PiY2NqVzw0DDiEDHSSWOzIrqn5viarxlg
UMLuL/2EeV/9AY3zFCL4keQqsqhSgsHQ00w1yo30NejbMenYy3n+n6sJBxZr
yrCWUofXO2qXPM+dBduk+ro82CGoZMoxfpXLFjER/FM/3BLt/4Wr7ay/etrK
qQMzCY+5FQi2fthEPq8IOA3wzgBXcsHCVFkkPhIkaA2KxaPfL2i51lSdknOh
nXXKKOk2c3HE2lKLBztfi2TMByi816rM0N1WR4vEan9lQqHzwr8+Mx5yMiRz
1zjD7Nd4wv8Y9JOAAVkNEqlvl9x0cEpkA3LeAl5naojFDtQXoxN70N6g0s2A
aDj0Kt33P0eCD2B38ZZq5LAVzuKNHdhHWc+xFHHNcCEduIW2iUpD1JFDNF20
FMkmTnXTyl7gepBADSTLRFnTHPFgjxWLMNSNOgp2mY0uzuqW1n0pHQdnnbGu
I/n6xaWFhFGu5fdD99AuxE08C/uPRAArt3ZVq6wlKBvf2Ylue4U2PjpkxF1g
TG+bRcRIkozPBHa7GdEncTUqZjFYm5tjtjnFoj+3nTPcjusdMRhNGWr4CL9K
Oushw+E0YDVd+dIIcbWN/w9NpHM09/Dx9IDqqBeSWOyeFABdLtjcpoMBzbHL
CMH7KU6CLrqaY1++Y7fMosV6bbllBY7Do1aczTEYO59GsVuC4TODRw/6aa1g
lx9vdWO5i5jldk/Tqf3ihebLOAXVA/GTYmO+gndJjOSACYpmJZwXmi2WDuOI
lUWT2Cd9NH77ADpCTis2eVs8pvX63YrdfOPC8V5pCbU0NMqBuK02f65Bbf9b
mGBvy9gbVf2nciZWXpi55YcduSmzMUa9C37y3eugHlK/X6spxOLkqeatRLWM
7J3cteFo33WHvYjfENw3sJFdIV3RebLUzSNxO+dzW1JdKOdndG2hefDBJ5v8
CeKr3I/xYH2FwZXHsg6BZE7ji+MfRXGXp/YNTu655LY63Fsk825jSkR+PJCy
er28YyBm6a1yRnRt9JZ9+gquKAY+drottQxIviac3Uotaai4gIQg11Nb0/wl
bfKeyj/pIyGeE3EjELZG0etCGFiH5xLzeH+W4VthMWpVSlweOBQifwGjn0sk
vDeiHlLFTiMfcruUddQvgQB/tvXlUXDLlMWh6OXJ4iAS03/nby2CCk++H7yW
as0WK6zbkAoTeml7aiWGVzymC0H3OLx4l9kH0a954URjE+AQeBNfajSjzI3R
/k1swaZ07xuZFTccodB2Dvta8zYRxjqGxUFZ9BZl+0MGoK+Z/33xTf5kkmpH
Ctqh9b9dozgMpHZ0fVLjOL2K1AjdVIatvsXH2QJ4VpMZO9rwueP0QGWfZ4og
/zbZDPW4Bu44mtkCk8ZCaXVlZox03ay6NEKdRJuE/RIfPAxmKxVfxOdmuOu0
yEiK5V1s3r103IOc5D4V8T/h3mH0bwZ8vAhYmFL0a6yHFO4Fs+QBhZcYAGn1
nKtIYOaJjDbVZhygFX6hHOtx0Th0/jSo9F3yZOz9DajYCEljRnxRuxJQUckx
0lMrl7hZq9tPGKBjiN0JO8EaGwNHYJ3m9SJh7ziRmcVnPJLgi+U6JASg3gDk
TF1Vp4R1cmTkzMPBT2airfunV+3DAR2RvVWos3rJrZK1BmNqAuqAafg5QsRy
PPLbK4t694kpNT+xjGTF8YS8xLz+eHjE7IgTLF9AWeudxT+Hi4rvScPbPtKb
tFJXYgHGt8NMCrY23gOy0TR32lHVBkE7ny18WkJc35cOHek1ItO5NL0iB5wS
mzAR11U0fWqok+O4cnvuGzHRmovdZmH8i98KH1l7iZW6/7R/YghHVMGCL6+o
n131EhtuDAg9DauY4bv6WCBM2bmv+x6YOtCpPRFU6fA4+TYzY68gsA+4cCvC
no4M44GZSewdV7DrhZDYj+sEgli9+ckt4fn2cV66cK6wVHdSLXz0dpxFPXYX
Dq74O+V7FafesFY8aTGinUxz8R4qbMDIqwvGk0+o1FAzUteCbMvjHYD2mPxe
hfwdEGRLaWkJpmDQ6+qD1aig4GgnW8CV7EGkXur2nJLSwS1tarQboXPpC4wt
HuuZPGBWfck+QCBM2P5VwVyH1neuIHx18Fjifaw8jK1FOS8gpVz22U6ZutFc
INwHllQee6sflqHcWqknfBlmVXyHe69Fb0v8cmYQMGqBoayP8O2gKRFRl2SO
/QOggx8BYdOkwKtLKYZz5Y2maZM4NNghm6Y6q87pxf5hbUuV/JG9zExdBaEa
GDtk+NL1QVEdmkd2diufypDpnSs3Evd1mkcamZ0U734aS6HadE5ZAIna01Fl
KwPe8k6XQTKUPpPFPqwOeR51Zy7WA4dqw6hhtOacoea1QiugnUyqlsuFnE9d
rYmKkR+gj9ARqKq6jRltAbWPqATkdEBXT9KU2hT6aILm/R+uou/hW9M8jzBa
D4tn8eEwPaHop0LojoBiQzOLYr4nP1AZcapdkA1+T7u3K2BHrXu7nmqmAtpJ
V1BMSz5I/28CqQ6vhPKwfmCIcFLVcNikF2pPFdcNeA+O+E1JHaJp4MC0jd5J
aqxLsrkEQ/DsahfsJfG+YtfQ5gGlUbbvLfQot39VP+CFZtBoE9r24VQQH/Ec
++8CN3f2SyNTuKF2GJXX9PiFvg1X+xXnmvZ10wq+rB/cokJZM7pjMw3AfFau
Lptuijh94Dxl6W4XWPmA5Uu4TX0Rj9D8WzrmFZG+LyaSq7jmA4sVJGYkswj8
Gh1QtWBUYB/ItUzJ0+VDEYMeRd9A+8mZzHorTQPJPX8r43Fg5owm7n/ZR3OY
qrfKKgRYrQ+b8yTvi2SpMNGOQkD8NB2nB7xOwe1+ZQgDV9zwUI1t9NV85AsJ
FwzomCKJpvSAnam1YngN2i5B/4c6bp/spELVwW3md7fyn4QFChn5wxQKJr5F
x8acMwvCCeEgxivC80gBzLPYhEHlLHYIvxerQw673zZTM8UQ0MwHKVShL2JE
IC+agwm8otfWNR48HWI5FK9sSO3k52neq4E28tbIfg+jT7jrGmiyNbSz3o5h
x54HLvL7tKMSdoXAjLWeHlERblxL1syV6y0bhNNc80DiZQ8e5KTJDw4Eed0r
FfPT/vxkhngoxGoppDL0H6C0oFRseCrdiqrLRpJeJDa4OmbeeB7Y2YvutKlQ
0MPPeziXr0Jwx7H6Bv/fcHu/Lctn88sjXBiYJ44RPOBU7x4rd/TOb1lLHORR
xkdlvUUODubr1fSoBPKcwelNYRJjTNunjC08w8mbyq44aVICpXAC7LRhXxRZ
hXgZowxL58FnxTINZQAwiB8UCJU+IdgHerh5zGNHvvlVM5eH0x5gg1Rwbowv
QtUuziZk1YfSY/TUd+0ks3kxHD4VkbpCXBsHtwuLMqlOYhakVFErjFCAHVY7
aabYIWnAaF3HHcPLru/Tb7pNTp93v4qgBgb7PaIvcANZlTN93te/TrrQ5ZiU
C1AnNeRlfJFyXt5xB9BKOLSL86cbqjr1yelXqUpkNo0N2gwoTTb0hfxaUca6
yVhR1+i0ByHfj5OxHQvptjfOlC82wStKBjAkrWX5o8HdlrS/9PwEwOGsXUoY
Yggcl8TIBlxTyRaOlw9SQNOZ64/fTLVeTYKuGCrZ4zk8YS25EhPBRB8Z5+wk
CwlmUAj2y1BGmcd3xkhqywpJyG+8Hrkg6CVYgD0t5xCQkGY6zBFULNrRdYjt
ojnoz+IRHA/ANhwNaBjTnwI1f0l7J1PpcWMrKdEmDgNSap6RSDlCOcSzYtBu
sCIvP6YCAFj7b2WOWrGqi+/eJwLWFHvtZQwyb4CEOX+R/DPjHszcUU0Laksl
5pQs4XlOXiXdxzB0ZMhe5a9rdbOwXtyQUCM3iCbrmg+xaWDthd9U0GNFoMuw
lUJosbSzRTd6TIiJR2vczj3+g+RRAo7a3yb9dacx3UmAXGT0cA+nJYSMGEEj
eKbT42CEx5YGVkqpI1k3LB99LTHOifhRYVoRgf35V7X81U/Vq62CGL13p02+
eaMft6PfHwM/Qk3ExC+3rFYEqu5FtlTW1LpZuYd6rP3og3AOWe8qUWZ0v4ai
3KpIFXpakLIhVHRxRnq5DPq0ylDzFdCxS22Te4pr9/qb/LV3XdHzTb37Zp3c
4r1JmRjkDe6RRKyfBWdiFogz+pdEhJ5yqzjyr4+R2zaINf+TGeCoHQV1bPk5
V3mOpjYi9ioxFzp8+inaJvFgeZPsV0kTMeufiK9G4DuGekGbds9zHtfnKeQN
/dFJiITsHPA2J4VQKQNbcND+jzhP5S7fN6BurJE6ji/n+60Clo2kAAhKOGI+
vUUo9Zo8GCl9L0YKI2lvb0LP5AICJS27eqJHtTJDoTUGILascV8cfSVh1O5/
M59fdHCWlz+dAYb7ps9uCMKQkJZogeVqhpF6uSN/QjA8Fs9MIz3A2ZRaK+9b
t08+2FEm4m9kht7VNgklUhV6k3fQQgWBgnM5yKv5q1FsH0pTDpe/E3WFHlo6
Z9rkk8MZ9dUm5fwTcrq4yj6we12ooXnu2DzQXosUj3g8JKdFbls9dQZg6xDB
OHbnMuTTwe9wSH7ZiDxr8lB0o4FbEWFI/ukgNriArA3k4Rf5QzaLkWhFhkvU
V3TmOhTaKBhDFTRr4EVSJVhczFv42owQIFpOEOGxYQxxrOs0udhv0Y3+2lDr
TWq8VSi1RuWrBZvZhFQciU13ST4AKwsk6X2DhcUj+uw0cyE4SL7Lom87gvU/
8E0szGwBaY1YaYaPMPDEwOiQ2TD8Sut32RSc0WR12pZ37F8uIRqv+Qk7gc6I
b+NvS8SV90hcq6qO9c9kVKqQzOL7gJ80L6MgGdSFQQkE27b36amo1Y6FDkGc
qGNidlDwkVK1OWD1/f4ozHcZiaBhyuC6yWXKBYbsVtp1Nh+azpTjAjxhNpYc
yz8uVdkBt57C8XLAYFMYWLbUQR2G8aqu/kX02ySVVtCx2L4e1HTXyGuItfuB
JpFSb5X2s0aEBOPWGiVX+Bg74s3/V/nP4c252h60TOLM25bJbgHSakIg+4gJ
VGRmqsAgSlkh9y0E1OPUj+M/dS1bGSo5FidkrkZC8ZxuxfAStdcaIo+f4gOT
0tclFOmTHb9zIwlTN+XjMezcWqSo7fHrgqVrvCZltruv8gWdnT97rHAOp5aa
1g2C8IcbG1GT86+dPguOpGZ+WmT1e4+8IKM3xKpfWgAR0T/EBsDfbrqbMaAq
9ngEozcVuBIY/3qR92iYt0/aFGTCN3CNAbHGcz2/d2GmQDOhXrHPSKhifP5h
QhI3s6+m+2YzHnnX/ne34MQ0Nrg/4UQKowVik9Jf4o8SpJ90d3rRIGCFEfiK
MWDpbC6OqoeY9AMcdbol31X24Gwpq2SV7ABXodpF4wE1MALBstlKPkuBoMIG
ZeOpUhUqkT8AWy5Le447tbrM4EZe0Yb+V6qSa9er2iMFG+Th9ft0xI894223
LsQxvIkJHcQmItFvnrxSjnIXD40XykC93s9Coqw6lvz2g4yc6ajiCFT2l+GM
L32G7j8C0QG6AbJAHLriwf+ShlqzJtmQdtvnjrsNAErjtb0q9hUYvNiEyJvY
uX0MqJjcyCkYc3WJkb/+3hAn2xL/OtS2ttuFUl7WbpC8P9q5PptZnfzUnZkL
AO7wye9hS3iPNQWPKDs1y/ttNrGeWhIku5ZWSIrmKUf1vibJTd6GieBVdgNo
LtfRSw2pBbreXkHDFJ9/hEWFxEzmH+8+miL0+6rARfOjjHIjqHHKMD8WNA52
044i4vcCFld64Qzmgn51BIRbX1VceoVlrr3gjjunwepmc7y8dq9Y2ycJuY8t
NxpRdAjfxs1dw6tTobMhCU8M9GbB7Wt+A9l9lnohoIzSMKxV24RxWbPh+Tdu
iRuj0Pnv/Lw27TnOmKefceqkYSpy4iSWNNye2KnIggm3PMxReXwwhDxyX4qy
Z1/6Ax+AK3pDRpHMJoZcEOFiunSWi1o7OnsMHx6iAI6wKsC7PwZ7kTPnLiTi
Bbr/ncJcJEXtFmaBOzZPcLWnarZ5/Sv10GxqwpboOhWPOwvQVH8Lyp5eXIqm
J5gunqlX5AlDF82ay9tAaHrafZL213gr3+Cew/o16cFdcOXxp/BNEpi95oJE
cYuAj3d4HWHMzCCXavL7Vu5w3ToS/XD8/29HLTTMBkx8rQVUYZ3vzJGNKAIU
CJx9jCVqfMh04tUyN2Q6HhBtNnATCgKnh44moS7IE5PqKp6NogVLNYgmww1X
CCb6vjCPQBw0Xcm3SJi4TZB3ioLOQSihM9dsEFKDay/aPpiI8R3JL7L2G1ay
Ny0hAKPjj+Jt2uFNsxrDlCd8DKkJmexYIi0hfDxSWFOnJLym1+8je9ogKo/5
H4NKCXY/lG/erwsB/VIf8ZUQBOZLCyyCb0jhXkZP2A+OmN9lOjoIZ29t4jBY
euUXu15g+rmyJg0dnbDnzm8N4hR6cUZhyTF9gEoEH6bEgNOwuQ3W9DzcYc/n
5ERIykLaqPCuF0AbAI6FH1UjI6oUTCqdolPYXA9TegGDhGv+giEkhII09Cqt
jQfJiDJTFzMH1PxIujcor2nu7jGrWN88H7NpeLegWJvEAYRJOPCclnz3vSIC
UOlbzM3fBYwTGufM4efZee0TEptzQsgGB8Tdv5KBkH7jHYPI7zIV/aUaLAiX
kFgiv7LZB88CSk74Rq5Xxj/PwEQUn78k2SQ2QZg4pB1SSq+2EwQ9YYqtRY18
QmXVNY/edIHpZSvEivIL3JJfoipr/1at0hljbEflrD8AMHBgE/3D6al5J7QS
KVMfxVSyboQoL00ldsvrbHxmxglviVsP79nb8TLxyageuB/Ykka8LjqBGUsB
9gEXS/8QFKY1SsDJxxYD0R+AyApMdDExExHCEdCbQIArzjUMLL3C5y1PelqG
cNaS6nvLb5lbeMCmRJsSI6aAaoV+gk8PrTXVsYiORAER3PuzlgtEMmRwVe16
Vs8H38N775H4/yiVCEliQIaBoFT7A2k85rUeLN1xOzNLdlnSch99wq1GCgAP
Kg2SAcdVm+pqYCMv0txMFauSXu+rH3s12dt7ybWDVoGHysJZe2uKDX6lBDmq
31ACO3IKJSUajsjrcNEwoiYb5fyQwqf/6FTh/cF6y6bKVyZ1DwBzNhog/kQb
3c6Y9ZbuxtgVL7xLY+FgggwftQRUVykzzA52BRqareQlqg0gg08+1nuhEvQ0
sHOvRiT+MM2Jar5eaApWcdwT8QYl5d3do8AkHuMQjZiSvVfSZB40gNhfGMtI
Q/1zeS9ZvW5T+Rm8ZS8MXC4qxv8PG4gmhpv/DIBCJUCto2wq7CJ+tkEnuUOM
x+Esrkj05JRfcqCM/tYtm8uYm+czp96acdeoxzAPF6upABnS2C2WKnXeBxf+
/aX+AM8uwDATYK6yYXQeOwYPpYkTj5HAHvU/pw6z49EANWDxbRpwr6ZEPibO
la02TmjJMWHHFjp0EAe1iEahtYakWQYt5fPmNNc5/4FOiXtkHhPrvHgB7D2D
G0eDuzxxylb8pnqy8hzKVN77ixdIxwY2Hne/EIb/JDDA037BpDr8A7fkDVdN
Br/ZsYeZL0zusavnmKbcV+kE9DDeCa8u6md7XH9ycM+YZu1c+qEYxohDTzFm
5ClIUtJPmON7+Np8+7npare688jEZPyi8QEOV8H9REPHKZi6FYu3B4XG6mXU
g3SMKye9cXHVHOnChHWdSp4dmgU7Wubfy0Zfy79Yikgo4ya/dMNG/05QeO7D
EVp3mE2de9BN65P6CGiL6QY4tqR3cmxymZkU2kTbdwEeHbG/slKQFmW1n6Q/
827IN27qRxoEuF29YujBdoG6je+L1MTgUdILADosu9nsWAHPbB5ZwfEY11ta
Sgu3IAMnVYu+e3mHF1HRWqgtVqWmMJUh3YbiPaKJObwjuD1mwslqa1lpf2m6
VbqSdI9DAxplODgHRZdvyvExk7h1RF4IctLerHaNOk5gg+IYI6+z4iWmajXK
hGN6Vl4lD8k9CnL1xfIrBfST8aioNGSRsyg+xqdGHFkyKWEnEyW68Yl03Xw4
r6IQEERpz1gcEhdt6dRBG1Dz+4sP6hsOjD1HsoaQ/V3jMw0oFuZktL5rggJ+
ifpljVCtVr+f2ZLcSMoiGD4SkVgzuwDPrvZqaB5ctySVurSNp2+EiSqMCDfb
a9w6xigwSl3E/2Gk6DR9ifGsytEvqvYyK9SDkxOeIm8R8PhRGGh9mFo1NMCa
6YFw46S3aouqsOH1YjMwPg8MYWk8/aGfrD8KIbjqpKlkby0B5s6xB2VzgsSx
VLXoEHThnOCwtKYWAq+lQ/aRQW1JuN6TJRinUCPZeCkQnX+pEMod77xHmVwT
5bBR/q8qtC7QVZbj6Y+QCHDLci6FwhVD3r9pVbf2nu0stDbx/FCWYrk5jVtN
w0WSDcwG5cumUvf9j8fEiczNvE09beXcKvpvc8t7SLQTnk4+4Lua18y7e0Ke
VyBvRn15QQTqcsvx/02IQ+xO3fgKa0hOEUbAmVdmw0oVSmf50Dw/5cXq1VUM
HhmjYRSGnGu7uztIqVa5kSDUkmD+36XWg7U9TN8/uH2uODPrU5JJKWSxFhX4
mnnHs8uJR3rijCM7andHZ2nyC0NmSSQ6RceBUd0ke2MRnFq90GmwAKYi6jV1
YSlwbYhEgLj/sfsyuTLPBOkybTVZN1EeBMcsswgTc68Fm/aKIZHR99Q2dMpu
a6ej3dFgD+ewG72AbsLFkOknxzZOOMCRUAJYG5yMqJKLCzmF7t+/O7niZdb5
vNhaHaBs+JbdZ3zVNi9BMYq79FCpWlhu+BAglXIJSGJpT+Knsc+4YoDUUy7z
ea+TxG4LXUZSwgsFqPqHErWm/T30swZFETlDFyEVnjNYCDTlVDqM1f3aPT1J
Mm3vkTcbV5nLeey48niWvYW7u2mG1MxgASkzgpuVxxOB7qDJg2fLEg449yja
kjYlt3uIbIsr8QnvIWtgGCYNc6HnbcmexKEMY9M0Vjd4HACWyAR+UgxRYFRc
jztTOqqmiQ8ORy7wj8oZLZEpi5KbwyGB6EaJSYorf+wjWH8eiSYcFey5Wbu0
TIincfT9eZr6wse2P54YiHQ7AmEe0IErkZXds8IxdR/kwHn7plOdutq0N6O4
XmTKAQ+9CFwuYK5QVIzxvdYu3N9x1tIB5X1/x58WyZcHhwfkLbhCQL/SUmqn
X3ZgK8TN4wLFQZX+KM9+Ef3dSDe9RWoFH+7D/1QGNCvKSS9VgEP/8JA2BXXA
8OxeQoZte6uRdocY9bjWQ8xLh3vvZbH/jh8R4XDGLNOGqMstIO2JoWaNWc/2
DHwHfnheK8aMV5dTm1r+Xh6zRIuUW8c/+1WGpsThy7AYCBZp9rt7DMIri8kg
IcNSsSY9VjhAd8vbgrh2PrlinRrB92hn8YbiavYRw1TJ6NG/lKp5vSYmTZGP
LHTxVJcTfJarmuQAyxwI2mUSIE8l4QyBGIH3jHMbobfdscQklvUoG+YyurzW
hWjYrQRg4fNqkaTCLDuJHO92huns0xl7itVuBkhpEaLagEGal+yli1tlYqj2
D6DHQxWeyIjiPwx3pQI9rIBXCupgUgvbXMrIGlAghqZRbY6ZkztJOGn/yaY5
VaiJ9Q+TRAKe4jTLedDBBAneNyZS8qj1nC4mXR2wmCkFe8XAsQDmGHbQ8mC0
oPlLafL+ayVMWfl3MetRNyibNoFZqx9zT/gv+e56ENLA+WZ1jByi2mikN6IM
s+SQ7v+w8cjLT3yKBqxKgWPmLj2K1aE54Etkz+woo/5Dv0pEjRuHCfgC5yLb
Dck8wY6bP5dpU6X+dGl1ZxbQU5KKfyPfsAi54h5lwJqtRXvlrRSvxP2y8bC8
C2iX+5g4DNfyTdOYUzfLkbtBovl5QenSP7GgcwoN7qG6EMral9qIDVOkn0kn
CkS9ipXyGFAeluiKWghX36CzowpQHqUNae84FKdM30o0uNqyiOs+zlo5LXv/
UvdfMzOB6ywNGsO1e0qpaZtdpev7Rr+iRRLHRNiNcAC+4Zld+HkiEaDxydwD
ReL+yJ6rHDQX7ryxV48WRTX0QDcgUbdQV7d8/sSr6LBzV7O1krt81iF61fIv
Qe71ts92XbgivjCdh3U8m/ip6zKW2CAI2NioK2xquUWkKww19kQJLP8n4wtr
FDhSnNFXMd6PU++ZmEUbtMqkLcdr3ST8sePSNzMSt8xTa5ZlZP8CoUa4C5qV
has2v7jkQAkQsKlw8vhukouamtt6XgHApnqMU2I+uIjMs13RzG0okAxz3hPc
5KsGv6fNF3bpZVR9XQxA+w2gIrDqJ2NN2o01HCFe/gIzxwABPa/EHRcn8GtP
xDhAilNcqJnnaJy8PcvYLzvFJHJmbkbqYkl+CO0C0g2r6jBlij5ENhK0SuHp
Dt6UEAzXYblEcOGVMyeOjnJenHh1nDx3MCODNoVmHs/RaTawD414ozunTZRL
iCzEtHWs1uXRazkfiL06imyrG8t2+6PwDW4OUjWLxZEhKeiUzBhGpfOXuGdd
A7/CaEl0+nsjnikSnIgDYA7YX+/WKTPMOHAi3N2oquOxSuk3N5oT3auWE2XB
Ch1rf/1SZtzmc1gZEjwyZ4oZnJpg+9dbOaTEBPc8wBEU6xwGNIOOaW3QGsU4
03vngiYwqfWdgbf9IeAQln806A4fVTxBxZjErle21weR/39pI81UpLpQ/qBE
28Drhs0kplCPEXL007TMphn8RHiDRCGbkTFUmfNQBbVZomK1egZirAMVXRui
fgM4G3ryoS2pdIdRkDR7s22p9wVcPjGVu8pEnJgR8JsGauJy/jie33CJzINA
z0zxdWgNlbHxy9A/O+NdXYA274qPjyUx7EsfN07i2TrqafZaml8FFj4QQOO+
SBHIkwxAyG8Qi4YeuEqSAULPR1Za09u3/VjC660ZB76at6UOFjH80CgH8l0q
01Do+QoUhB+YydyA5XLNgKT0H/hT+e+2cI5IVGJK3c4MueyRlHHU46mcDHZ6
GMEMYzIa9eHegFcYuNBLLZZJSzN8HKDoiiVPEB6tGJIoExdHzF8zD5vbol4a
Vg3UAfc9OW/Z4Ci488TGq77AxRMeAzS/zg6slyezC+VPNFobh87krRO696Of
qYK721X61biMvSW0UPy+P7u1YxPGiqXA13SeEUJ0ouTMI/0XWMWf9AHRljoK
yw3ZMsEJGM8KKPfM+b5mp2zLQeft49DA3Hn9v/VIgOsh+vOHS+6ybVC0rT7g
r+Dw8Ce7Kjz2GV4R+3rEgzBr9vK0GmQs17w9EVklnHFgdcwmS3Oen5N4n2gw
xR0XB4n5bnAxpL2J0ckbYdYPgt1k1l/QtyY4kNmn0NUMY85XCapXnyuSTbJO
/gtQi68bzbudqPEU8wS+FBb3vac9YIohCAUbrii3kldbOEKnSWB9NBqe1oNx
Aiz4izYWglise5eO0urMY/LpX6xdj0Uf+smqfF/47rl8d2XORd+Im21/m2c6
6LEIRXjR7TKWeezX1TNpF076YFkv1NvUgVhrhGuUKcx+KXYVQ/2VWMfNVB67
GhA9SSskMuItFoF208Zcl4VzDiTbjT0AQzN+5G0sR4xQUQEM3fx7vOUftOQj
MxbdfuDkzLzP+WCw/gV1axsXLBunrWx909qakk3ll0SVCddzrGGGIO0EDYGu
OBWs0BVVPDi29YaphVGNcvVuqAIwi33TBXez1O6EZ2QF83D5Ag6IVOEvARM+
aOIJ8B82UfQ7wotx9b5C3EKXaudXK3o/v/TnX0Aa1BNjwQyzYDAmUKibc0pF
N0iGH7OiMHm+9Hsy6Sm6ELo7zNpzfgnR8QCT45Q5cusnF56Qh3sYZ8OPOcxS
qJNbiw58QPiTraEg0crVNIXzmFLrQESWpSM/VRLHW0THDFg8b78aFYt4Xqxf
di2FOqyJxuDasNrTcyioFa8gl1JA2cQpcRKWyCkUn8XaqRx9cINiT385BZUq
aW5XZ3Wr0WoOIiM6EUfs7ZkBSmvqymxJRqRV0M3zknTvHBS3sIkuWHGbXWzY
3uZd/Mbnqy9N7nj+XHrbNgH4lZHbg04N+k1g1DKnwOP1zGyBEFKBY/CFt/HX
JBvq1Tv1E01QuMPM8HXmBCnLkJIEcOKJMLmQWh7q6FRCEXYzxUUkPu2v03kH
KiOvttMsfReWkQDr/OHRV5HxeeNZwDflJ96mA9uGmbjDtFBMfRtXA+cJ6nA0
HwMLpi96p6wuzSEF0WtpVcpoQ7KFhA+BPORKcbVV/Sv4ZbEIX5eHWJVwYwca
vzRUhrg6AINSNwnlykC5jK2LW+8E6+Z8idiXkvdfA/93lQlOYwsqnvzFH8qR
xE8XAx4MFoHHn62DdaUO/ZnwFIjT2DG0APfd6K/sgfia30P+Bkzdz3tAYZZ6
UA9oN253LyP7JpqARj+pVMm3ap7ArKt6pgMQEOwnR0bKzra0lhTgYIaUpIkr
PS4mTKZkI3M4yvFXXZqFFjcTcn9ah+eGNBv0nEeK5/SBTRDe6rFKZZZXjzAM
SoHi6sh0RVU687yCXDV4SeKahVErzLwM6DeiKNbI/+I7SWL7zm/DtgYzlGEC
bh5FPCU4W/7Sw+9xhTDJ4SH6MULvdAQ1w1At4M5d1qH40VGhFAdDd4yMI6IK
zvZrHOwCOqbezUF2FgvGhs3vCqxc/oEteDTU7ldQFnUNx6hyHVvz8xsdYQki
6TyfS0V/Vt4iUo+G32RV2E5Wk5DUMUKZuM+0X0p4ntxdQ0SqX4GGIJ46iRxc
EfX+anF/aeqfEJOUDq94KhgWhkKdj1AnDRQZaad7vSz6CVDQnT52okT33sWR
uC682thWOQ2KWyLy/RZR9DNRUJSUwGzt4SU0WqAb/S+ZsHblHISoka0hoeEj
LPUOlYvc1BY6494bLu1S7e9I5RuQH80kkEdn7Hidl1tOyl0u+osOwrl/QM7K
i7ieN2cEM3zqB+Lk1JJGjLmScXHnCDbTQ9pRysaI6ZUz9bbztRMe/NfETACX
7ZDLPWKP4gJt1733oM1PCLNrcoGV3Jj87KzMsSajsvrZQC9rjDs/AZtDYXAM
7psqzTguaQ6EHvfgJwB3FMJsldbvCOc6oJTAV73kpS1pm8qKhCquA5yp3J64
AhcUJkvpmi1pwhjb+huCndYe0rvJj42HwD3FkftmbQlrpDGYvvBVU5oCP4S+
KMkzZ/EC0+gFRD2BQ2S6fcMUIZs2J6hsFJLX/GlBNJwiIcosjVAFeoI0vjD/
eDl+xh+NvF6Jg3GVLJp2MpuGpkSVQ3xyDLtoANGU1hbKBVy1kTrTZair1sKH
TOK7kezsaETG/8msodKdMlL8z035FyFoqeIRMUnyYyGSJGl6GNNIwKcLAXHv
v0MlRfLgwyFJwFpZf46fbig92srtY2VZkH1eH/9zjr6CBfszSYc6bFM62dEf
NLvvdY6gU5nPs3VlW1sONJh9FFJk5HGQm+9OaCzl7fcdCMohAu/vma8lOdaf
LK60gwIdvpqiJyUOLebQ6fCSCqPLs8Yw1YL5gl6+rS1fmD/qmq5BZNKarWzI
bHRaGpGRzAwsQYReMSnDTXQ5D+5Xsfzxa/YIUyduPUZ+tFdgX/SyQ7GX3CHA
yNZAxIVJHa11HaCFwOhzj2JEe2bUoxiJTpSQ+yY5WuKrBOOBViwNHtSfV1jR
VaZTL5n/VV/RJdu5R0a7JuvG5MGORIZoCC4FJ1t9QQiXur47DXWAXieZuycF
AqAWbSqwYh+cBF6Fs33e8wgPmPG4e+4wfGP8/LLWIJoj+UQDqojNWBdL+bwH
+UfSCqbZz8gsL9oqbGnQeIkqtUUizEsUwGXuQ6CoI0CmXPuuf96brHkaJ/Cd
QwyPNZVWHLmMPiu7HAM1iGj3ARxhYCDuSp9SP65hnqvFdMmASjNyDF41uHly
pELEEnDCk+XhLd5abqOncFAykFNme9xQ4qlKY6PU/UzW9aixZBYDfYdyLXer
aFDZazMjEw8zX4AHVl7j9h+cdvymHgnFCKhy1ZAIFQWozIh9DK6gZGUiMpM+
QqSyJAA5Ts7S7ooxLH+i1rBnAOZ6jltkpS1NYqlcm1gwMhp1svYzc+Y6QKg2
w84jKFs5vF3vsvz/ZxDTNfJwiUQWzTii+9tSKePkl86BkrFI09kF/Q6qByah
53WutRY2e615sHnsOxNYgOo9kHKP1Aod140CAvjhpExPD4KOvf5qrEVCJR6h
mN4t0yUC0ZzjJE7RwDq18CgEuZ5rWIWz0xSfUAjg3FKbmdI3NN8vUf6qx+oZ
5t14P0s6j3wZuQ48hMAMNwuW1oSk95HjVcqWN8g913HoOs5DeSZWZMLOaPgR
qGL4LCjmT9TESTu9DSmTqgx7wh+lkS0+yr/VEUc+zveQPiQ3TKeJDAFaPhAJ
9GjX3Kdliw9OkSr5+O8WapMX1OA0Xwfck/epQqL6cnNaOFYLWgzUt6ELoIap
FYig9tZ6h3+RmQqqLa7Bxb/LHm2Q8GEDpw1cdG2dqUYIbiFw2GQ6SAxdVl8J
Wg626nZHSdWxcChqre1wEOuyI7QiMDGUGsbzop29jzANjYF3aU7s66+wAJrD
ZHOp8AwKwZ9v6oF8FQpAQqBf2g++bUQ38JUCyvp48Y2kjEQNgIBDWwFP7zyT
HkXu0lZtZR6pWaVek3QObsK19JjFlYaTg9wOCbUDhB7EpeVnVbMaviTEC14q
xcnDFom6J0HZ+g7LJ6eFje6QORvfoLyXn7qCoOZvscpa6rCZSNvD/d+B5hIc
8cl0AHTtKEZTALRC1Ry3LUduF2R9/+jduJZ4aw81/P0ztK6ODHcmerI9Cujl
ynK/TEBAqq2UUwiGf7pHlPSYofv7VPqEOWUfUgKR6yIRNOcj7YsOanG4UNpu
bLpyFyCLL/cd/OZ+Z6fylZ89P86uZSngfrnlRMnVmRfr62wndcxsVHqZSYFP
3Vi+uZ8CeMFvLxPBFj4+ETw3KixqRqnnIRuFlMYBQXqlotZ6MnVC21zVaYtw
NprDcF5+SO3CJ6kpdsrW6R1QDqcVlh1x+0/AlTdbeHQL/U89UwwC7BrIAnjx
gwuB+8iU/ewmzaE24/1wkcs+EkzasmOY37A0N40f1phpVkeeH2Xd9PoDR9PR
3nv1pspWTMGS9RLr7bpP9Br262eQ1r1ELCXL6jmx3kpC7yrGc/tE8phSDJAQ
XLGkV02QXLSEXHdeXiDoKR0cgBIJn/Uge17LF23fK4kLMT0veF50pd9B1nbv
h81cy+YHU4qkSBEjGXWOIZHBeGLG+WPqBTiO8h35mxZJF54fAym3vAafY1eh
1jw77rF5M2szBAw0QcNlLP4RoYRPFKnNVkM29w3dcr9NCm8xK4pg5itIPUnK
ixOQ3eWYCmRsuOwJtCszNIOwObQYQ12JyQQ0maIv7WWILw2BG2/tOm0WTeW5
sGl8r/lWpsOZDPULP+lH+T2yB5MAso9gMvD7aJ715Br8TWWJmGjX9dxw3oFu
Rz7yKlT0V8sm8YuB56BCb52sl/e146z/qWrAiF4gIOgQo7QO+XSXJHziHnQG
bYlSS5dLlXoPkqxFe3qUrehGhIGLVvjXPEP4kCi4r13dtKiuVp10HMmfS+Jd
0okNWMCTEv8eSGq2eUcCg7BAMHi5PhacehB1iPea6GwVuaMxIU7igoyb9Ov3
5Tlwy+ZfUgydBslliVrRvZHMhoJ4zFWwPl+t5eRLOOntDHG42X/Os8cb2INo
ZJYX6oG65UnwEHXfCktENxmYQ5YpPPZk52Bsnm3DpGxCyi4zxpl6Q0m/detE
Nsb6wAJ+GMatd9HUpoEv01xHARJDb3bke7JOTfTYbcGZdpPKFHBzXhmJv+aK
lKkgnimEEd+LtVAE593ZNnxIndIq4ti1GyMOzykGEAEwX4n7foeFmPxn8GYo
SIy4rWhZJdNP1pYWseMrJmURqlswVT/2bo/tkh7s7WzC3R1NPEliDPs46nj+
YNnkvzEtkMZ/8I4ymHY+tIhsOVgDcuNZ4j1ozBx1Neuxw+xGlWMFt2l9ESEk
aagxsRGJT4k3UAqketM0Oyj9fdMvSGXWC5ian0tvs/zvb6LsRhot1JbBnXtH
GuD9iLaq3A38o0va2FCbAWCd6bubPnTAV80gHYujUHfmbBs816JC6BuKP+fT
oNHbC0K/qteRpDf7t42Gef2zXNozgxebR/u/ec13gtWACRaiTOl8uo43amMc
6WjdM/M97P+toyUteY61Vnmou4BOcfH2U4TPZ26OEa4ZWqKK3rx27rIsOQEM
utZV5dkCSrCqHFckXirYsX1SnDHV+LHW9vILhx2bIwL8SxaLFQi7lWu/gUKb
QzsO2Kl+6sD6wpCVkkNKbi/VAezwJFjp5chlJSoquBt2gWV08q2YRIT3cz+R
CDKrbC+6i0j8np569MH2xFAlHm4x2XAYx6VdJinJG3hidBuoHI0t/jTUqaXa
vATHmBWO5CKb0JNN8BpltRqDactVW8nc4cQ8bKQJ5XB53BSRSublZhG7un3x
M+bMvt2zOFsLQDwxIApZEy40wv6xrvB6fKWauHMPshxNz3SDIbug/WzHSM9c
1CSfxppls1cGZSBsKl1Ik37eqVHzxNNspmvK2zaTX9X+lSJfYUnuxTq+cVsE
rhsrj8qkYX1PnPkrztM98wCl8AYZVVj9rYww+G8XAEerk30lczrqdDmcWamU
OJwxTnC9MW5hb5DB0PCG1IdiP3Gbux6ff8E2+IGpym74HC4b9rB0rLWX4IFo
1gp6H4ecY7tXYDzjbgfozORBxtiXjR9i5tiqLq63MxkuNAI/bjU+G+Yx/hii
T52Anl2FpgM51yEFZQIOaXOZg6NPIQa9WaBfGpn2C63RgboCrBCZm9OSf6iu
YpscT8D9hy3jf1R+pnSnrsCHWIwkMo8Q+zeler3/TMv/wsmRBH24wT2xVmpP
C5h9XscYw72pqQ6xtYyAdRFDhUXG9O12/+B0RGf5Fpizb5HR3jJbaEqdZ3QU
TSl/hpVR/niA77VC63UWQDAL7rRvCzOHj08cVXRT3D/izsVyL3QSHY8MqAP0
lWfxq0PBrPzIPPQcbx5zJ/dKZN6WYuO5UjbX8hfNRvSecBoxbVw2ieNVNx3J
AkBxNpzkAs9k6RhYP/9BwJXOrdBVCMaSgbBQmKmA81mg5oVlOnsYOaAD0NWn
N3wKSLdExByjDxZTdlw15G//AKIKj3evg/iGQ0t2WVNvcLGzraEx/kcpL4X+
/oUzQ+prepX34Vs4MnFE1ktMgVaemKNNLNg5/D3cm+rSnlts/HOuV3nI/ccj
AUeYyrqfK9j7rXphTbHwqQSUjFnHoYgwD+zzziqHBZSCxN+9Ec30OxK/M85o
WSbV0c7++FP5Zx4M+CeKhLuA1nMs61Pekqz2MnetIaA01faMQXZ6uJELrpGE
suBKkAqCaRl683yZlAPoKLMWvtv1IrSYojUpRBuNIwuKgMOkPX97xf0wD3fL
x0jZ+F5/nQiacD3h305jmrIrkZ6C5bE4kjtb7Ler1HH8OaXABjVPtEl4Zfxh
R7xOUIi/7jdXrs7nbpD0uMpnG9w4HrDS++9uTu3gWCiBfewNlUb2dSiRp5mv
zNZnfjcoIBTA5n+LwdhnQf3cQMxEYfOdLcMOGbgyx4ssHW0KTNCr7hNXXKmc
fc0uQxv4yKnhSbvWkQKvyHz/qweBCBtqN50Pn5wxK6AVrC1/fUOyAhwUIr0u
g8D7Da9pjrYPzHFf1dTn6bm6lW9VNwnyADGtOhm/up5ZNsNtyqjUd70fb0ew
Z/WYzGqP2+Ow+BCzC75XRJ5k+WHGl/o23Z4ecUH3J2vTZhDWu5tW7HhLyhOZ
bGNqZymPfLmWIo47kGm8rhMOpD1ZHgpueJNN9tjX1m4vtvfHoniyzhF+GIbM
C8BENsO2bAqd6TeqRTstiOA3daueuul5Bl22OtW1U9kwftUVBKuZ0w5jWGa1
sT0csxiDpR2TWOVPckowi+I1Qdd/uzUp4ZG5B83rWPdF2nRYj7/E320Ulmkz
J3bZ/QBnYmBTcYIbeGeQYF/t0sASpcdFXdCh92dalE0srWCH23SqbciZ6LcO
THwit7XsfvmS6khVzBPd3nuyIedUATasXJVD/DfPhS4MdemggHbHNO7y/boM
wv+Wj4iCK7IP4pCO9dMvQz2Z76dT/qF0gDbKy2XR6wb/Gnq9nZOyRihNQ7mu
bqzBTQ8QNGpftB9pzsN9lvK4tmsCaBgogplFSXiH1l2eWHeiMNrjXzcK+psD
Il9j6w7RBqvT7GST4Y70+yY/QyQOCRvZVtU3QRijDG3CSz1X6p6m7xtd1Vhm
zNsKo9MHEzlq4wSAPC1wfHnbkqZp6868T9wrCvj+SLUFzxfc3+EcUsaBGQV9
tfPpw7e2eKywjeHtWNNKd1UrdzoiPszgw9IERWUWyjb9l09QUWIPJCaUOtqP
zcuvbHfv4VtTcR9Bq02ptUzv5tlhQf0Lkew6Bw/7Bj9Fjwfg0+MXgUFogTk3
9LOl+Zree0K28DDUv7CRxD6VL9JOZd0+6Y+DIKEFiNQR+X1HbXt/fTaORbh2
HBJJYCOCn3q/srazclp15yRAyF0XfncsyQpC589aaYDG+rAwhhN+FnE5Y2bE
cNKY7uupRYWuTv4az/Kisb+m45qDQRoMrPk8SReoy0xaijUf4paqgY8Dtpqn
k7mknexOgZW4yuAE/UnCvD8ap1FvOda//EUS4CdVrQC0b563rZ1+ivlC/X52
dUM0sK6yVFFwptTQGUz2Ki7G9YfLjet6RqtyMwyY/pXK3biKoW/OT8ApcxvI
FaVk4v0GNc2j2+800ueeWkZoUpz6b7XluW4l5Cq6SleaPatazrmcIa26vyw4
ppcMIWiO5nItigQFRCIUo2UazGSgfAhO1V4dQE0mbH97xcQByum8lYRYUdzT
qDWZAb7VHXwNgPqcPbUuQQISjVjy7EDe5MS39XeEYTIwygK9TQX05x81K7MP
rsqpGQPvD8ScPij9W5TJKPx2E6+y0c3ArLTLLhHGO+OOa5KFDAyVMgzIWKsZ
iKMGLizs1CHobrRdNeYt82mfUq+kUTrVW/WyEqlIIe2SHacjnaO4cINN1BjW
W67EekW+PyX+PcDcUfPaRXyjRZOzmG1b2FjwIbQbotFGd3RfIW/U+U6jMaJG
72LzDle53+FznDknATAexQAU2QE/SJR208JTdRXutK8Lxh1C9r3V123Qo8vn
Ex53+KDQJ+tES84pghtqu/8IHIo6fSGJSPvjEdhAaD6RMyhTlkGS9Okvk63D
oLbGI+bTAjMJURo2lUdbIgI3sOcSrVFoZuv490UbWaxELfwuFQ2Vt5VxWrdW
ZccpJuqK+D3pvMl4A26ldxIjwVCmCbJhNMjQOFvuBMb+c3UO08V8ShYssDNa
TOG2UkTDwkorYjZux4cmfngaHjGF2DJOhxR3qgjp9mQRsNeJHBSEh6wIaL54
r39MRkLb/BA76vZj80mHCJsRpr6x1+idyobTMT9dd89NIOu0jpr7jkSwx0PH
RJz/OSDIXwYCCd5aV9abKH3loNe+EMBHs2WpmsMT3HJdnmnlfJs+3zAtZasD
WCk5TsckCMnzZh2jkrA+Bl/sE/uWPJr4fTtN43HRG69yB3n9ZIW2NcJgSZ/a
MA/vRWMf16FERwYTBXUhwjye87eDfJ4LLZ3FBrCl8REk06n2h3ubPv7mgLSC
jcyxU7r6+VF0FYROAVv4K09pdlJg1l+GcWIdItIKmJdqem2vZEDq1exFBezg
gZFmjYC1RH4wIsOcFnWVqXfvGKOMMk8jhfMm4XRiKZSlFrzmCkIso2ZsaEaz
FM+XvDX0a8g62xn1OBoLESUAKUSKM6O0DkwQEMXKRD2u0KYmxnHXeQdqtR7D
uWKGtIEAQ4nySCPVttOnU9WAy+UxkEpflOVDlBv25MGdXiEHGY/4gGgqafgS
9E2noXRSME8WY97n4Cnj8DBN1jnt3eg8DRJHr6Oq5ccjlQI9nGsi0rkFToWh
gPa9O96mxrl9lj4yF9cz7mURiKb5PPLH/qWSg3BGdfmIbXi+Sa+iV8BQy0p9
cvzNjD5gMf5hd7wpXl6sN7y/4cAYY72GXEvmzBPEmNOYLFe+x47+4iQT36NX
3cuAhf/IoQhV/8DBZPeT6B0jt4zU4hYKuREj2perMDwNvYt7TBqWUMRhWefY
sOfVijo2avJq5ST2hWPpQJGseIMq2XoP5g10hj2d9Nzt1e2N2iYTc9JHnSdO
w2nMnXFFfxtSSm1nFOr+9TcRzyo+tCA9wLVAZOlHRS01mlPLUf7MlRytoTg0
9vp0r4gqTfmk4w+AmGcwkA4dkF1NpGwwUK5ohKomw52y1Lc5ZKTJGuJZ6nZf
Zl+2ZKGmPBG0tPZ5++bSMJ9WQ3QU0U+NeMCSgqZj4YOUd4kNE2tOtG+mjlXL
ZX7MePw1M7T7T7tgSJyLBADGXILM1Pd4JK38dn3mUeQs5hNPjEid5Fxx0j6m
35HbPmWGI8TIOcEndktiQxz4il1DZBHFUz+ZoRzfLXKp8GUKZwcU8DpYZ+9I
/z9pI2KvAyjdUJ/0DMtodd6oNXnFf4KNEFwiWRDhSgEOxgIHPllp4EHe1gim
1wxb6DpnlRiGrC1CYvXqQfyAXFRN5tgHDQ1SVv7vy8OSSh4RlBBS6M7QEOhZ
/j2NICefT5L5l7Lo8ptqlQlXsdD8kwxH0hHFy3J3LRtRPPT7mez9Cik7Nj2H
nZK2KoktGQfNa22cYtZ8iifFzogKZiQ1ZjCF6yXSeTsdbM+AfCR0+mlSByDv
FazCPlwMg60Qh+/WQ6KGSyDHJQSXV/CrJe2YAaLWwdQImjHi7O7ySQbNtOt4
cMkIR7k94nvuISaN6nA+UPGv73W0hztE8pxfz++rSEBeMug0k/rJrMYnWGkM
wbFEBBxT4uuyGgef0OUDOrLaio5/w65NeI22vVvN/28VFuFvDMADrgXArHXn
OSMOGX1230hn724xQR/9RAYkod0bh2Kkw3joaNbHOuzXwYsLylZppwJCaM4Z
YeOoKKEmRgqH2Eu5EDKwM3YuuzGhKhYn2tDkfFlPRmjr7YzF70iN6/kzwVYN
wn3x0kgy/Mg6GYena2y8oNPD2v3wFBDF+RrwLeNunT9Yti+OJbQIaM43+fNE
GkKCxXKoxd7j+yNBK2bN44GTTmxA/J0ogyn3Jn34eEvcj2dtCSHyZ4/g2tbh
Uvm5/krbNhPBEHR4olGTtDpcBWSX/vTd1SI9GIW+p6jhO3ULyNo3ZvaGNIdt
9NWDv1s0yxuhaBxQN1JXB8C+Wgk42ak3aZWj+mxDCR1QNYZw8U9xrA3hpZGV
T/zM42CbtdYLMoNHry1J/Umrwz304ZzLfbpFWR5RbvU9XZPChwhXROc/yAGj
IXjAmhn7oLY84ZiH3iyyoNljF8QT+qGJVuuXZZk9tIqKKMHHh44B+JHsSwa/
hX6LBq5mTEvNoAEzMzHxU57GqYU0RFluAf6RWwwQ9nxfwioFLAsaVl3rdArr
Q7jCi5qNCgQY/fqbMnNaq7Zrv1MVP4YKahv7YMLovAtWdxXwm0VOfbIDBoWP
GO/hcPoZ87u+wf5UypM+ls/b3yzbFK6ocOC8hGVOOBgga5DRyXYr8Oe7cZ96
q3jOfIkq/J7ZzIUWUIeHSaDvxpyq2W+hXyKqvY2JK7frK+7eOSTt2neQTazx
hLtU7puRKOBWf3y/G0zHj7ermUS7GOcwtpp6+Bt4HANNR8Zi3xvVDR3g8Wpm
z7owMxJWOJfVTqK1AnGcaBzF/hiyPSatwWEby1hY2/F0kKYtkA+7wLoGY3ox
w7hIkpsFMBsAO6raInozNcYLvd723vO7zu0UfJCxwwCMVwWDLhQeEadn08sM
uWo3e/cp6z9DdOHhwNtfg1n5Y6acnqJRrJ+oOiAobcAm+/lI/aVv6sbjFORa
43LrBorD3bXIpGIeiUq2muUVA6KlpxFfoUAuy3dVmPdmxs9RUS2/TxVxxfWr
Qytbp4RAnDbfMseUk1o1snubMp4n4nnRUHS8X22ASlGWS+pEgtAs2GLGhQS7
hRs7s0zCPFS8kcUUvryJFaOXE3davmyFYuKWT1Gi3fAlWDw5wY/d66yqaTGW
7UX0Oz1j9VUysbh4uLkUkfVrWyVpNx8xyuZSuxp77Hdj0YyiX4JgJl5mNVK4
yHI3n2MwBLZdRniLc6L03Uc7eYujxzgt9KgoTLjmwjdzg4E+f4eGAXqF4XUM
9BBRAJ/4tBfFHh1ViQ5C/HojzgtVyRG78huzhe3AUEDq1AVtajdXWqeCqfjM
nFEKOmOeC+Jd3q45j7Cy3I9kJWAwzBMMeLCpkmE4ufArIUXdVmd5klVWdBba
Osnek9UaxFgmlLtSzgovYVS1272VNKV4js2VzIui5VY97UIslUQr6Kar7cpD
DMpfoQs/0EHFK7Y8K1EMgFbVTzhXCA3aGyAALkoTJFOAG6sNyKVa3SCm1mBm
UTkhPf8nn9geL2B5vYuTEUwpVCYfNbNnPF9S8Eh78A/BsG68HiJb3a3p4Fxs
Hg6wBV5Tvjy1baBJuHYFv8xBEG6VdDpi+WIMI7BLcaja1kGMdCxWwAUzgrjL
TJlZ/iLaoLUG6df6HUs/R2ntiosY1SyBEtZT7DYM0+YQUM03pWiy+YWzEF9d
uN80Hww4vteIOtHxZiZNL+x8x1wtm26lTIM/yBiygf7WLl9LXD3iBkWluDMN
exat0HpnyOUP1jytfvXj0Tr+7Ewftb5jO3MNBdmRlZ5uOI6w6j+gLPL8EMOx
Yd4ehbrgTCXZHXGs8oRLa6RAUxUZbrqf6lDeerDq6Hirk+Y2OFDhX2vJWddn
JChERD3izp0G9FKRxptH/1JsPuqpg9lglwFCOh6s3Oh9kbuA2bbZufXJUshu
r+brITvyEW+zFSFimHzakImlIOr5zTWWmLte+O1bvGAZd6jeD0GTzzIVmqym
/6BQkCdoXzlyE5SS6OyQ+51a+3CLdd4COMFJcgMX4Y2v7DkKoF9ok9b409tB
4UotM1nJ0uzEXnwTlVmmtG67zw3YrxkHl2vn7K7XR1xKlSXYmR0xLv4rQqkl
TNnKCauP5VuerB6OKzruuVcotyCN6wnqJImS/by5XQwHR0OChN3DFgNgt3jA
qm74kUt5khKc/5VyQ8/JXK48iQ/GIBQB8+g56WZDm4bmGk9XfAasXEzdoQ1a
9rJA78VGObjhRlNtTWx2BbDPB4QYvuyrbN7Fm1nh0IA3X2qD1Kqu3Ew0qck0
n1ysNtKwUZAqaBVmXwPbgyJ8jrZN2dRMSjMehDj074S70OGVAof4Tj6Ribob
yUTLAo+dVkpCWuPRj0TRJ1spDtipHc2JXEJp3QMIZGAKJegiKe6BdpIohQ16
/CXipRE/ldrqcfz/KGvi76TbZ2kb9WyrHXeBPhvh7TUmlpsEOGhb7zpuasPW
ZkROn2jOmM//aFwElVy+Ip+MHdIJtszOo6COVUR3UEelV6ep6HS3Sw5ur/IS
Ipo/s/IeFT3+Cz/YnIZYnSDXJCMLM3HTb2U9KMavwPEkmZkp/XjmDXt3fddG
keVDqN6E+7ApaMESWUbthkn/DQnFtdDxwonRreDbYGlUhS8yksxvFGL73F49
cy6InTw7heFzbNvsy1SKnkXdWvBNMyTDScoWZWWEc/vsD0RllOb5nvEob+Df
vxbS2p+LsAj29/fILSYTy61WwEXroEHOe9zZ+xl376LAWal+xs5BrGcGq1su
QFIBbN4BKm8/RzboQTn8LT3RnAS2NsVRN49gUIaky9ErOC2KvQD+BdUIOJMp
9BfUmzeTkcg15H6SpFjsUXwFORXMo/fg6CqomsmPDmt86onQC+E58ZHKeteT
WreGKEi+Sf1EwalYZBbMCXzExKTshURp+bTLCZ3GPcVBOPJWBmVIYI1cO6fV
tULhJf/cVxpmWQlCp95fuDxB9pRem3GSDys3KX+NbWgAAZN6+PE5bDtdlwmA
o7EmkxXoywi2rZVmpKPs9XHeNl3DHDS+ZIIc1AusJR2B9wLaYJe2rd0Wqc4s
Vnwi1ITfHDXjusPxT9qujihD8Nr+xK/W4sbUG5Nbf5AYVbcTNpsTPdR8ZI0L
m1GmP9wzuxXjc8jqFHtbVzmb9Nb110Lrzo1KckQzjhyeho90hHG3A0NeMRc/
wJ1D20lerkuI8JzEm2DgfhkVj2xOWFKcLZ7RMX45+6QmPNSfpsv4AsTHjchE
vlnKSrDDluicbt0ok91AMpFG6eCtLZhErmUDBxN9/U8EeakOXTeMzdH1idjp
NcZ0x/n2Hltqwt69VA9EvJNvvG5H2NGNHT5V2chwGeR216C2TS1KgkzgSUCP
dx95/GE0A8WeTlqs/iGjPlLZ3VYjwxUk7pqzV5A94yxona5VHSR/DdMUthuK
MdL3nFRjCDzOWuLS5L99RzTqdiIL13niRbAKZ6uiKmEKyclwA3nLek9B55Wl
QvCvsjqPnDjzzM5TrBKEdpzmve6RPQvTqNYo5mNouBtoYzANkbon5k05X/8v
zDRNAF/09fbgURt/8qNPMUw8CI0kfumL3x+eG7KBwmdMVySaU4Bt3ti7fS5u
eNRbcEAc4LsuRPk51PM5LT3+p3B/LHFicBCfOnzbnMDjN2dOI2i9cgMJ5per
+jZlk9oLVEFW0cDVbAq9OA9BhAyuaSFvj+uLElwFwg4DHQfZ1J9zw9hecCRQ
2Ekzolb5sZhsOjFSzpC65XKqM7yusaiVyqOFXBUnkNH/WMuJizKumK++0e9t
GLdP1yzOuFVQWlIhgS6rjxZ2Yc1d/RIuULg4cXmLsOYov7b45XkjtpO5MTEO
VCd95pYe4rT+T4y7KwZ6GvqHcmPd5V8IVJ2xthAzrtxBWCMmU1Dv7tp2oB8E
aUXZYt/sxWKnyavNPbXXlBvyjApPl9L/dNfbEPJhI0oL4EQdo8cq+wFKjibl
Ts5sYsb3h2Ni8vAjsq43Jn8k0EWblQRV+HgCOWWCUudBs5UzJj38Nsfh/KGH
WA3hfLkhL+Q21IPsAGkfmBv9SS1qnqFVlREgE+enPQq2/sfAomIsrLg8Y1Fw
65p/6xyPLjGw6Qd1Gpn7gji+Pcou2C+Vaec9zCv33n+ilPqCR77BU3N75C7i
4IfNGrY0UJl9U9BHadbB3U8SxXcuzXh35ZimWjbS12wJcFomMr6xm+8syZ/9
B4vqNv9Iw89FonjnWath4j34naY2B3jAR8uOrUzCcq9OV9gkrZkl496gRFyU
msh5ZHJOhu88Zdut+dpe1wUKOLgqlekGQtiHe03xT90NfPpaYYV2RziX04IJ
+Cvdz/GdJaMPnAQdUUgLlIEMK2/bsTx2aI0C+WA08JshvOgFhBsj/L/Dfr0M
g0ear1S6Ul4mViLEGz/q4vZT3l012LFsyRL/IKKGS1HaMlgJGCg+rSqzIc5n
+CBHL3GXA2VlbK9ZjnOKLnQM5VEcSL/yfJlh8tMf5uohlGaz4YXkY8t8693f
EeXsdXPloOEiHN2iZujjHXm0iLFzyOc92scp3/6STtEi80wJQjephly1xfXA
V7WDTPrqNJPYuzYfWYT4EAAGLZMo62KMgusFGL++N9t7Sdb3Qsqjn+8Pfs6U
+l+Ys+r/Ci0oCBavR7mmNuZhM33wSDDY1eewyPHNdC7RPmRyTkmDZ2JAutkn
K9TJdSs+jSsfafx1IXArJ/tmVg74G3cL2TE7NYelijTB60AfHDPCIYyxXSQj
Lq895I9Lt/WJRBIwAX0iQCRy1knKpb8JzM9SSEwKLGPCaO94px4ij0IjYnjK
mAHL8mnJgmyUiTFnwJYQDWIxiwjwkhOrdG1Eq7T8eMYA++PNLr4c5vP6G7Yc
3mi9ZMFHG4JaOXj/dTmHmAaN0tRUCLznBHZWo5GG32gXmGHZ87xaHeybZnnj
Hv951YzA7AMmRYJpL1JVmGYHTVeOfrXC/fxYWfx85y0EfT7lJH4dlOcBroPW
tJ/dcy/KV0668hivcYhyoBBdxK3XouRI3yA62YB9q1C997B7pAYTsWPY/uaK
WWixkvN7Vnf5w5eOoCQ4Ds+jVV9PdFTzcWwlD4qlfS+6XvZh5erJ1E2blI9u
Zy4Nq4/LC+CZhau3Lb0oW//g+0Kx72NDGq9LaYyFNAP7lu6+abibNyFdGivK
k1q/tQpUyZE/NSB0MNr/mTBGJhhB8tGwB5m/dBKoAHShnfZMiDFyIcod/FC5
IXiTBTwr0TYua5E6QxQqYoip6F66mNcHCkEcO46NPUtCS3uRXNZnwD9G1YV7
lv2w+QLYZcl3K0sIVKfA2P79pMcGbRlqMORsJQ52Q2XP+tBnwPvcq308NI/v
ELdH7kfvW0HiC/NPJT1gKnFkemTYdVanmOmXqo+k0cOJAPF7t1o5e9qVW77T
cfcGQbGGAx3/ckWddAs779Tz3l3dJ2jCpPkpOr/um5EosY386LoJvPG1Cdj4
E32OCPHCsfgeMHLatvTkizhMoyx+rSE7ky2KvqgdL5kC2/Quu8Z/S++RrrCI
gcYeRuJ2AtpvrzbnOtjz6J8/nLSmdVoW/yOCivoM4h0qsHAsAPqDq0aZ9gXB
x2y2fJjVpX1pPJ+MeT0c1jZBMS/QOQUwPceqoWtKC2mtPXOkgp3bwH9vJTOm
pv+t+dEqfsx/WFCrmD2sPwVWhUiM6tSRDEF1QXIX8bMDVdxZiBaASn4SL/jK
vxt3WXuMcG/JzzgUOTn4n7P4Y5uOemqnhvmOfRqzWakTfP2Duz0Um1alBylm
9Gp0EMdVLxg3X7e0XC8+Ti+qmxVBwGW8Q+jmyBnB63M0Nw7CW+KTzz3sVXG9
JU7AsC2Duu8R7OrwqJz/4YAMcuHbYNOc2OzYhY0UEksRB60ZpMEjUAHOzgDU
k5MsWT/SXSXhfFqx/sZ/trYo6pA9lDgP2XBdBRjyGSJs5AfqCI/S3h8SaBXY
pcTeKEUhxo1lKgVxYiZ2LyRuAGm2VMzF4pSYeDttDJ12nPEAc2qlGQlzBStg
KXZps2/OAqE8+2DVKXqSmWSNHEQKURDOnXCAH53IMUEfXgcfHV5Fs73xF4KW
EkBooEZpORzSNQKIwDLiurj8qsft/Z5dKZg8tiji5IopAONJKagbsvrrHyfk
UR5c6IGxEn1e8DQnMQnbAgDaJFee7VlPOd6FV0qZyE0gNh/iQ0C38DPoxb8T
oytowzv1aLbnF1J51XDlBXM5uFAy2yICCgFVERayRIJ0e5NSq15cLlDS8HSS
PHW1IjhldJaIiCCitxbDvArwWmn5RI6bWtCZN6s14qKrjZn4SozRYXdJRiv3
UnH7sKd1bRC9ThSoomXFkO3F8snQMz2zaEzWqTv6Tt2KFa6x4K9yHpQ+IpED
GfNLjBiKdcRx1LYPDcLnCEDdUlRafv22cHlxedtKWIPQhtjQ5vaCFpugeSxb
hoWSJA6iPWDHV8X0ejnJdkt1sT3sLxVoBbfwaWoVcbDTReBH/K9ufJq3J9rn
nbDRLMqtJr94z2sm8SN5kThrKwgf0mxNcD9SCQhFTb2r8jAD37Zldz2E5bgd
gj4lPOpRRrK+aZy8AuuwdhCGC/ejntyTNhnUwt09QjOd75wq+LnsaiMONuNz
G35IlDziNcMYZxcl0ZCabK/7kPi7np1qN6DDQiHRClCcim3+ing2Y5sWumNt
BjKeE4+M4t8Sfckp2Ci7i7OC5KtN1HYojdIc68ie9fWy53jO6C8AGzfab31k
ybP8W6FZISDyw+2wMhvhXQzJVJzmIwLd+etxUmqVHkshNph3SAEpvV7i0e1a
PlrKolUyTeSeu7RjCRLKCAkKu5Tpobgo2KZxv6s4pTRkQfIGErDbKC6gQ7wX
63/P6+VHi04P/gDStDJwDOgJdwpNrHMaORS6CkHG9exFscXgIEfGVPhvnidW
SVTnjpqAvKMThaGh9MMPQApLVVrAjFx7dSeNoOoXR+AkQ+XOSdOLcFxDRjSY
HW6hhgub+z6gbMV5o1JbCQ8pJZR1HLfjuqDL7WMVy9VzoOVAuHzTC8eJIjUt
kHwpeNf5gkyEgSxD1Im6sSin4MvyiHXPyvMJKV0Br0lxGOwNMqLlx77uDTEi
6WhuLeeWtdzDn2qRZ6mbUBPrrfVq0EBLEslqahPG8yHWX04A9M7WLf2EZtWs
rmPnyfbQpvEdkd8uWIcA4FTqP2/pjcFpo4h8p+A/AMDVcqbxKUKBm17NSAUG
rYZxlxGnSNdja/G0k+hjsJIDm3AUVk5vHE0JfaK8KsBgQJOmTfd5RQOnjv2Q
WOqY2eE3686zrSKGj4SpIVbnhbQ7iyJ3eZhoVayU6ATSBwbLdwEqUv3klVip
HLUaA4jUMCx88/KIRpb6k5/5nXRbn1ByQyD0F6V7zybQ2RIeBna9Q2wxgUV2
M0IjwRGAijjjLvEnsifslXiBs6Vhdf7YCPDxDE6fHwvBQRtQvAXfXapUo+c0
gHpjQf33qiUxr3UdzIJPcdYbatKpgDppOQXgz5jXAwL1aMS/sUG2u46KhxGe
6MozT2Cj2fZCXbIqpxBfrM3VE/AfE/zaXy9DT0gm7Qeash/ByJ7RxzHyd8ZU
h3I27+S9K0+FUR/wAekhRdY0OOoHcD3Bdq0r4tuHtycoVHBSkUX1css21aiy
IhStF0S4HEfUgrG4oZLLM2ywb7ctFimWNMaYSXNW7Vgzum0xy7NO6V0BiZb0
3YtsOUCRRvHzRjGIe2UFUFer2BDMUpb69J//XUASRaJNaCPubh7qC9r3oKUe
jEvgiCwVzYQ62qZFYx0cLjvOIJ5rOhFb4Gz+7JJvXs238YFjbDshy9uYj8EP
yhGkO/zsN4Zcsn7IYUdbl6CcF+cGB2QUqQ9j+Ay/KU3WLUXoqpYwWTpgun6Q
X9chb8azkFTYT18C3EEU+rYQpLlgMx3fCK2nqNW6nqDDYz0dRfWjZY4vEza0
DAQ2blYjc3PdB8u8RooObn1dph1CAI6gC1OH1VEQ8UU7zgQfqMIAD+56XOMB
9PKn1Q2h94Rgf55p5gc0GQXdRniHDI7ZrHv7MLR8RS6+hk4t4yTd/X+WKAq5
xR1TgWqWbpZY2VZCkisVU/1JuafdC51Gu5b5YDX48f1GyE5TDbOCZ1TSTCC0
wcgmD9Ch7Q6rwVhZz7ZphYMFWPhz2Ud1gX4tyWfF+CR7ORSG2cD9k481PlPR
9svSyJ/ZsSJNklITY9+TbcEP5AMybUzW2aKNmBKpws1yNb3eClkmhGy0aAjd
z78rslsSJ+tZGxzBfqE3B4xJPrhHv2NAjZSJJMl7ztk/YWkgLa9o5ZDu2zV/
idGy7+Q3DDXzA7elRBo64lJKp3Sd6/0c53UKNC8Jo81LLWXgsCnl/WDQf4l1
nPAcznPotni6T5Fx9s5i5qbfwQZeIClJ3pMmrEeZ+6WQ8HtUggTYjWbcpLQ3
rX+sxc9C79AXKWhER/5w9RnGhHVfdf35u4v8g1YVUTeiFn2bWCeLjaXL2mQO
ent7UFrYVXFGIQS0El1v3GnZYd8ZisY3litQinr2DarCtjWP6vJwfTx6trZz
9f/Sqy9iI6dHWJ+HpAovhXUy/i0KQEa6SZ7iV6zYYT8TP4wjgmhSh58Oeiy8
jtj2aCyKTCPbNDTHfocQHYeUYGNu8QVj9tC5tjkuY9QUQ5Ee+bzMQfl/nfip
SjzhapX9ZfZb7f/W1CGTAdGfcBS6/PYVLIuBYpRLq5MFfV7AKZiQog+/58NU
ox7d/8+gHxgsd8Ng2qY23Ne2ApYISQuMiBRcQFkLTYPLF16kUiAkMtEvVPKK
SL+QCY8zQNtA6ZP7BUkP/EJYxRilGU7zJEDkS+iXEy0EYiptrI/r7Zlu7K06
LsWOEbmu2c/TNtNm9wX+Q13eGbseH0ItDCu0/jfaFcgY3DwbfSwfrm0G3pzY
FIhPijQi8zuIBAFJhZMG3yPCo9A7z7zgAl6eWJYbQnsMJMowcVB2Fr8aU0h0
F++8YDBw0vNKUBvzSML7zqnim/ACZrdYzeMHmeZZ2/O6ljViBCsIrYCu2aR1
2Xo7PAfCoD3sSabfa/rxAoaqHWEMKDVG4C8yqxGo0/BMlXbpNgdV+e81bUjV
01p/YSALpgiM+Wh3byQnl4vnAUpntwYtFmyLq4reTTTYO+njcPNllYKi6Ojj
9QIRcusqL9gp3C2iROQ+CDu07jk7+yr443YmsPG0v2s3lobMseRyGlUbSscG
Y+dLMJPFSMzCI905LbRzE8PBLIzxGUz7dBxbBOZzZC/et+Z+1L8A7b7XXUo7
whS75tfEyi8Pa8/uWczcVx+6chAjhblgS1bJcsPP6xhH2SzSMFNXE81vTC3C
HKqnSKGlIsgRg27pnrroVxp8071x5W7ziMzKsWebt2xEqOpPcKYwowdURq0W
oDNkHWbif1rZ2pH25OCtbts8snmf3U+aZ05Zh+5z9/ENbK+jmaQmX1SoHVAs
q5y5B/q6UI0du8bduNsQ7ukc+0aUHbbJMVJJUT2DaW0FWDBufhGpLJXyqhMH
DxjUleNRbWec1kuKnS2MOVm9V4SLdGKKMLFq/JuYThNzB5/9dTFKe2mCLq3Z
eTo98svb4kbpKqA63YdieSmI0Mg9wGm7Kwma1MarM/OueuNmfL2IKSe+mhPG
hWRc7fONJOL1wq3tq+yQM1ndMBuZ68MzeqgBPHjqZBqAmGbnGo32fAymbXlK
21ySjkK8JUT/PKI4qe0oSJPfEaRdAwfTNPJ0xB+5LhL+SMQhK9qhi0+0Fh24
nsA0sUXWdZDGMJoTfqy6Dz6J+Q21ua1MgKHnHt7D3D3Vks/fc106jReMvkav
Hc4qoavfgtEPQtcxNvL/Y81m498CY1kC63EKG1FANeYmVXcSFbmDjvDTdDr+
zf1uIqQ1wtg54V7Odh52MYgwKoLMO3pROkaQtwMiNZNrpwA8uGY5Tqkujrmx
3h9Fb9hy6YCSn0TZyZK0l2XNxu6/2QYB+v9M7GRAqxP1HL2fBaTpZ5Qw5S07
BzVta7lMjDQmBRdUUAO55HaIp7GRlvIrs37GusxlCu9fVzNh+VdU/B65ai8h
zpAUg8nNd3RXTE1UJ+l59MQh3ikgklFo4tdOFYmE5G8kfZymeK/8AGbh4rPx
GmzKouj77tovoQrcUZmjrnSW1E9YejnplRy3/dnHpkLDBTW1SIRY5Y+idpQY
QRnWVPd9SlQ6uT5nx/isrlzjK0tUxO8ccxSGbDyQfnADti4sNeFd3+6O4eZS
cXCfmU/ru/I4sR2ASnJa0tIthFO68zsDPqS/P6Eifbfh4Gx4PONIyO0TRXY3
vAvbzpOAFgStBAayM4yiIiHNnPF3DogXrBQn6FEoU3n56EvCSaQcqIqZdyVy
+6l+iWFEH7m3bbuFWRjNuDeSANG8ygslB2rKLHGWBRWmXTGoLsJfJegMuq3m
HMUVaIWJu4WCDqXWpuiUGycnu5AcxcYvhyLcB/m9ItVYxqurlK9PYqYNKtyu
pBQdfMQ51RN9YE/jt7p0h4FEkKztETp6Y/TFfmM0LKt++o1ghciDBsbUR/ys
xqTaEVxVq9zfEjaqDpdVl879bXPi4rGnlVshnbNdD70OME4LkPhBmN9Wvllh
GPUPP87qChhnkfWyYezrm0WmHviA3E8LgqM2RKYcJrVDk1iNEqawJfplRoNV
ZEQs8EhFhLwR9XCV6QyZVNnc4AHCRfSZj0YGjxGWBu4O17wCUYCkrL5b1SAe
AYhx/Hqmjik0O7WX7QdEppMR5AfZcQ7U5bMGo2OJKBrrsWuEvAvpBu+FpAqo
3eVlsgdfu/2+wre3CiDRpKZEkAdmK3xk/VpjbdFdajc4lSQmpkIcxMZlpQk6
en7iXP7NL5wkSiVbHF86gSMGl9PVJjzDfBmAPXu3UqO0EowjMOvxMgBm5iNb
W1HpYaoVBzNPVrEdeunTNfsoS3ycfOLZgLemlQMYtHl27vQZHDaqGJ+Nj+KW
Ng/hIaZfbDwNo5I6igxrd45BhIrlwz7PQNYmz0nV5TGzM5MOAjU6ygwQM4L/
kgMoRpa6DueGaPESJDej2yFmgTjdaqXwPr8tmOJWFEs2GUyLh53u73ugUWmz
zXI9APeiWs1CpYB1FmJUsFKVL4YogcnORvMWXxs85i4wP01SVq5px/DLj1b/
aHHoJXzK2GWKzY+5dMWEz0hMZOtinrG+iUIbUCQKpLDwYwaiAk9lAl/nRktT
VTs8FXB6xyzTET/51UyQNL8ERTK8ifpBec4Ql3h/aJ6MbmNP1hCkoxLO5FXX
g1jNvvXx4WpAUXY4FWa/kcTVJTF+ANYwDAwjzryXgt65a5Ei7Jw8D94vx15s
pWLVplxhdZBkkly1sq/idqI0Aq6Eer2IrZSX12onJe+IIhCxkZCrUrK8pO3u
69BhozKAm3D10V5EUbCnKQdE5LFziMDDna2vmBMprj8KFz6m+PwPWK982asZ
EzNTxHQRh9egWT6aSdUSQUTexorqvbrnhzBs8lcaqqeEc0ffNiuXuZUmrIbJ
qGLq9f6++haVLnCgNpZqAvKaTIXjExh0iGpC9FQGE3AKqM3Wfx4ZRUQU1MkU
FLsr1i3loFmJYRiVv7jU42QmebGWxIOYlv+HpxaF+t0geS4LNKkiDVNuqtRu
zwjHPszX8FnQDutHASUx3N/ve15IYUsaRc57Mn+fLWsoTyae0WJbaNo7Ys4Y
IOnHhY5Za46hB1fbhssVoYkIx+0HZzvaQtEgbkh+N4UqEt8JxDMSOhS+82OP
h0qig1LOiploBl1Q+mFg1DIUsr9glkgAjg/Dry/NHiP6AoiFpuJcf31WHAZv
zSPngOfMrZkdWsU+iNwFWazGGOusBuPqpoOnqsu16rBpx9iJgjDs3RpMY60c
CFZcnD7++neu7uVuxXx/ui+6cSDe8KXrKmEjs2CEF6/4mKgQ8N4hExvNiOoU
BSN+wpsAXxSL0nXBMC5eU4gReYxdfhQrzsC4XPVjVIPOOOU/IRLpQN+TX5DO
22sFZa4IXOB0t8xB6P0NHZpDHi3kjzR5A8wzOewcyiNtXxk3iVTu0UeiXC7Z
ZdK6KRQ1oTIUTmF+kw0IBycRbcbt2fbfh9ug1qGHoL2bxhIBvfkbIKrEq4DS
WNjAuadgAZPvgBJf8o5x5bFFrbqCdyfpeWl6U+IiNaKGf4ZY3x0ut+jv6Ds1
vLSF3ZRomEaADc7F38FknB8Phmep6Sx/sAOrW0k0BqfFhoQQMwIiLKBOGsjx
iJ5Q+Q8vCTrTJg6hsofbw2DakeH9E887SMo/K3znpTPJXkIRB9DPnmrMdSA+
Ps6etdepCZj0nBESKZJ+gCVyxE/buKyvcG89F7TMm5G1IjzB0SyYC7i5zkj0
LpbJfjI35dvwEotg/6yKR7Ce1czUnoQYrBc9MGcOoA4pL/f92dUt4Up/pWPL
2sgr0FXBhy6SP5GQ1PbYI8ZC9+8eKR1IZgUe+GVAf+cA6TIdklo/TYKKRWn/
V0GTwYi6P7JYHnCwjcIn/YjWsc3EKM2DJDy+guUk8DEgeGsGuNysDn7RDvJ6
xyAN3snCMZ1JvW4XGeR1J+XiBweznKybXxu8VuYucohiUgYXAXOuwTK2hfBf
tGSceSJVVR3zVeHvQ9ADSNBB48b/yQHx2UiCJtwofNQlOZFgGJujIM+sz+9L
eYp7h96Y9rnL7/Y0kQbM3XsEbOIqHdgK4bkc9Cl6JJOWYwHI1HVLzVuLvNk+
txBBYUsOZrHuCGrLVJgTVbzg4WL9KdwbiEzmJ3bpnyyaYrC7pM4qm0KbvXRf
cPriW+GiLO5nCZjBFhIvQ7qIFmxnGAJvUPAy5qQizwOtS4Cg9jVt3xxbQRQZ
RWyGcg5+a16UWPLsFsoDHFfSTjdKP98T/rN9tZyLAj4aLRQZOcJfZpLEHvhF
OY18IyfNCPLm1QYJ7MrSsABIgJHlQrk1aevNxfCWHROVoDHtFTRDyMUwwFnn
Fz31evPqAOaN1y4yd6Aj2ZZQ39AuifRQYQ74Klh6x1DbMdQwUIawx46j7dQK
SgvtLG6AcWp9Q1p6+ceIRwvkjCesZQcxBvCG5AcRxiaZL0llBH5QgAT18BmS
NStXOqEOpSPA7Ws5iKywAER1zFEQYi2spF9VC2tsLvRp3NY7VaqrBa6X50Hz
zjzaVN+UjezUuLPlnLQvtMmvk2iVYX8wnyU4ga4tbZZmtQQEsq++CfbQMR0O
Pq2Hl5YV88nHjSadJ8hmI6xZi72Rb3yygCbH45bjAH1aHRGwS/xJb9j2yqzX
SmpBa1cXIQ15L1/Zjyx38C9RDhDYC3fy35HyZrN4wkCiAEY2XNY3VFPE3H+4
SvN1BjLkeR4HFV7pJQ0lCnM+BkuJ240R3e+sRYOo0S8bc7ZuhT1yys71CbXP
xs5ko8fqANll2PSSZ8fb91iasW6F1isMniOMCJXKCw5zTcs2J8wTj5b4+8fO
J6WFuJq/usyI4FKN7hQYhoxkAZTWBobuYRzgW2B7+NDBtwJeqwZUwBpSwVWB
HMe4YbEXHWYJA+fFNZoa/PxLIOwSR8UbHxkm5UoSgkewzhi/57K4TobHi3DF
3sAA/KkX1iYP+Eni+xH3Epqn6Pt3BtxorE3Q1PA72zjYRq08gsO8ds5QyE/e
z2f4ZC4QQkWVN0TMqu251Ujm5fL3qW/kpR9F81nBY2C1cVVgZ31kMV+BIttS
sL1K4vycXqAApeTLU/c9WEPAzAq2opr39XGqaNoAyXTomKV0bSnsEkSX67cC
HvWYbDG4Ht3fqDUUzPkmy75zPfGfeu2BISPetAJopNtf+BiM9tOlmSodNBip
a2658RIEvmn2Cac0OuqrL2+MfpJdDRLsZjZmVYMlBH13cOPdjAIpFzGRJfp+
GEe/DCb+MqguUhEeFezDxlv21SEGZneBbw1yIbe0oAx5pu7e4Ghhtgt6Xl9u
LzISpzJ+3LXeJAXFoTHrDS6+ibvyoTxheAYdIhb6aFbB/iTMz4INr6ZiLsZg
0cSJLarYFGeuXO0sQLtCpPaADDuVdOx5KTiH0/NC/Bki/OissdO1x2sPGDSU
hRqU+FVUY3NL3CRII0cYK6Ni7x95JJCHzujOoTMstXf9h1aqh+Fh+ofdRckD
iWwLMnjTGdBeQgjTbk24APT6co8h7vRKgPzFVDFurYgOeK3r3a0r1MBCUbBa
R7gdFYknCxg3VPGJPx2kGCZQayTzeMkGUQ1OswqrewsLCn7biRM0lEEJAWri
r0Di4EmG8gdnjgjDAQAbrfJOqumB33+0VZh/gJzsN6sA5bhAyBUNd88i/9n+
pUr2zJGNzi+Lv6OJoR2uvWAEZr0lLqWgo/3DUK0eiZTwM+E0qseSp+COX/Dx
sHP3Dn/iTyL+iL7K72JVQHkgrYitpgMrKt8EDoEH9R7QGETgcd2T7JD+eX6C
0KZ7y6JsNwdCHygKgnx1IAn+/64RIn41uNXU6sqZ43sXxMLbGzITw0Tt7zaG
WNpeNgKcSQ5hj75ooZXGZnCAX/RtxgdJutpHMDOtrKVygO1I0uYyorwoNZqS
kBj5VPsygYhSwRQIeCGuniHkcDmj6w4swkoyw0arbaOqVWg6LN8ROlxHG4Qf
+GTJ1hn+Ha5g0Th+bc9yhFbFmsM/jmhzV+UojusIpMSesqmz3lzqBYrt4Pii
5kmur6U4fLMJeZ7vxXMAiTEe3wF+57nXHXs05tZGxQZcfgkssv43XNaUBbIm
sPp11v3v+4BIBILBHXKQejibo2qSgA4Xi1UZU97wNAupPxpO6dCoFqmMnw2A
N1X8OqO+/z3Q30gy+MQBAyyVJrkh4hQPiwMoD7JKGQIAGqLcpDM/4MJGgqh+
j/0/R9IdOPqiu/31xVuzqixfHwq+rhDF1fXaEMBQcuGMsVxUzuL50nrTKCC/
19D7nvDH167Y1tt/45JXfMw0qltM4OgqjQt9OKEDadfPTU9WFQPvX+Uv1GUh
3tz+coZKjeRFBWwvnumJhlQ/7AmKPvLrI3uoQdu9qYSUFD756ikLjZ6kNKZB
ankIfXOHlvWRftZiY2WiGT43EgOFvVCd/2mzUV3Y59f9QBlBoD3CbKLYAq26
mLY2bYGNJ+RzAqNW7dmRqr5oq08zf2Qb3INhxDinFEOqn/IKV5cYt41T5fAw
6KjnrI86070Njp+pLfcS2eJjfHsY7Vh/1YJiyJF8ok+kWzx4MEjqPNofLVf9
I8soX+p+g3hhzdjtYRTB+p4s2z/nXT2ofwxYo5BdL+cBj3+a2V2g7iRpwf/f
RYYGVqcrvz2XvZh7gq37TrM4NddVnLL1k6cjz5N3zUfLokLp5BC/st7hSkqQ
mqTsz2W5lF73SvEiANKUxWVYS0DfkJzPB4DOhh2NFDZ518VlVFKwv25WeFry
AiIWiGxhK9IhK2xC9RihxWQ/RJtH0ZPa60yRttFPYSIGmAOa+Enhtoa3J8Pg
UwWaGWk1YvJcZnj6+TmIa+nAkn/bMb9utKkkQhNuC2yrPaohgSKJuLAQ/xbS
EXM6jLRHy0ALRMwIyl44LSGu/5ofrsco+S4CGEvFpRe0wkG6xE+VOByu+5u6
Hc/8XRIpRUxh71YmQg9HK/L2K5MLhaPehw9cfshrdwJTVSfaTmc0WfxBCvPE
e61NSISXu3U0Aqs2jBh76UQrcfiC5vqIxCuOL6B/nd/CdbESRjxAF+e3Ck9p
10yrbAfdZfGXT9N6XFqL6SpJl7Ax9wm1AMdUNnkULR/V443UoMBg5tNaLe0j
Qii6hxn4swU9Eaf6/5DLv8Fb1vS3xvE01/Ow+VA9alU1wy/dKJZKb6xuu53l
4PmY252vlOVJiVB8Fqv02kazEWjgWHMhDcgCgkkAUioMS4JKqERpsrV5Qoev
yIAb90rT4q/48b+t3Fh+gsLO77VANbjJ0RlTq+SdfGxhjgu6i1qXp4vAr8pJ
sXAHQms5gXp9gY3zNYkZlvTX7PuO/Vh0KvGE7ZZgZ0hmMTNRUuJrixlMBJZe
/PQ7/lDRpId/grabOVNmWvGnfr+9vPe0GugU54UrxfuEV/q8tBWXmKojsGKa
pflvsARyFA8bcgjc2QF+y69FgGW7c4QRQKsbipB41oFbFCtMouBNt2mgbuGJ
PgCR34zAZOK3dwQCYsUpWxuDvtOmF9uPfRVdlslSiQkkGgBilWuAHXHUAsyN
hbDwiNIgiNLR867NMPIr0sGcCbd+cgu/kk61F+kcMxLeYhKorkAcsSBEOdKl
BLNyZJ3gFd67JeDmSHgJZ274bwwPMud+9FstGbCGSO3yqfLMueyTtssmhMBn
4W3hwSqVIxYPWVKk4MC3J6rvz8AdP3G8i5KSSjfGGMVcLGbcgDrEJy3n20z1
/a1XFqj7/TLOXt1PXppXL9xX4w9Y7SSZ+UgKISFpWobGF8GdYhNmM92cEK4X
jRTk8YZBeGONTDGc3qohrxrviE7eVfOlQ7AIgLPivrtql1n4Nu4vo82J3ecR
gOQjgA4N7hBMPbg/t23SM5E+VrO744GKbxHMWEZqNtkVsrFFC0I8xcB5PN3b
T88tfOebLHNuNpKZgwx9DPUOA2h94XhWFjLYzFtxq7JHA3RXBZFx+MXq8npB
b4tCHtV/ytZKHQCHUyO8BEjtBIn9HjxkoFl140jPop2Vkz3T8gTGLkt3I3HJ
8cfcG6gJ9GrhJZRFwsVCKw6LXv0BlUq7PTild9Ti337RbpuilxMtKSscSIXO
Ai8A3uYHxQvsZG/6tnF/rmShM+7AKZkIDZaB7AIHWqAM4LrM0YwolYKSd4h7
6Oc9qS1zrd9ZwBS6HlSTZ49C+DuSA3QKA3dPnEtz2zt/+jC2l+o7hmrlyYsi
KDu6udzofq8yaKhL4ZobYjO8LPuSZWpyUBszbU/ZGucw7SO5Vr58ymSK1vby
VFX+0EcJ2kdJGW2SYhs3vLulzUaKS0ogdfGiN9u2aIi2Bo47YRKvnq+xGwBw
XRHibQ7PRkeH863/MJ2S++xyq2cP3I+9QwRQcDm7nquKQwp5jV6T13VbOebI
B4THaolqsFHQSsBUcdzFM+uAXW2kyG6VIGpccltAntfKdsqDBlk7FD5l/mLw
8t0B7zfnj0/+LTX78JsY+c2iEAYGkV75GjVKvy6jtwUGiLHgbTjLlFx4u779
ESc30X+gEAT2OO45rssmlGL451tSMK6BdcCnQThT2Fjt3tik7hHLQ66tYuz6
+wgDT85BqpQLiCEiZshF1e/hscbUD+5ClC5BZvrOFPvE9wBnC2gDRb/9o4iM
yekZtMrlk6MIp6tNJ3frzI7O+hDW2o832B8Tuy5oLHUoR4FE2DF1cVnLViCU
0rA5qMlJ3Gg3rmhlnLykVINJbXW1LLHm2AQb6sniML1AROGk9zKqTkIEhqWp
LdJdTnlyyR/5PASaP2wx4KydFzWmU7QDsxuPyniUzJUDTWWDVHSvGWk/qpTJ
shZmjn4445u6OGHQBW0i67go/vJEMT0j1BdaCtRoJsp948uPE4UC9uiQbXAM
nnr5MVAxnjY5piDBvO/vxJbLVUxIbJI1ZNnOoce0x1Er1UVQ9CoGyyU4enES
DMs0AUYbz3gShirKwa8toivQYPs/E/Mv2ehohBgywO6M5+qQnAYIfsX2x6EB
Siu64axeDz3YyY9YXMqVNuSFMNtF0iQlq9bJvv0SMDDb+f6WLQIY3/zNDkjg
2Zemme9psKSH2x5HOZlRdKfjuYsxEA+A5P0KM8E9hY5ZiI1hbg6zsTgljxGO
q8KjXW7Tx2IMPSHHOVmkBX1IY9EHX4k3UaS2iXoYEkZjJd1E+niO1odth3au
RFg4qN1fFwNUVodSmKQEkZzbw9KBNLj0Kj9hTsmbY3QT3y6TIQUmvU21CXs+
+lseLoljwjsEDIxLCcJZlZTQQTL8k0pptXfY1gYqqWpR6kvcgrSHJ4NP/o19
t7RXm3V5BwW9TQ9cXIeA5Jgo6wJBjSyKs2pSjPg9SdljK5tIVx2+ydLXTNNr
HCEfwiPR12j82Tf93QSp25/GRhYnrhgyXYdvJdrq4DPil0NG99mjmNN1Cy5B
AYMbJ3rOxVzvOmlzH1i29nNKI+LEgsJOQL1tPo99s9H/DOMoPeix8ZLrSNJ/
Gc70Cm7E3jox9Vk2dsz9Z3GzzIk2SfbKM1JtWPcp11mIgdr5detDBCqWdm+q
p6c7znefCk4dug6Hb5Vj2RaCfCux3xMA68VjZbNCWcXSsNx/nFTWHYa1mdzy
Ei/WadVIVNoIYwd2UQJ2G+p5CueLcqjesbiQ6zXieH+EeHeDSkp10zAT0Dii
iEPJYww9E/kZPPP0s3HqzcXKDMQKxNyjmTn1WQ1mLje77NoJfT4LEUV/AGl1
ckt4DtuHZ0WaLXYq58NeKFD1I+DBvF3HfKsCTDJKeJyaSs6eLNuL2U5DCP3L
8EYanmd5J6+2fEv34DAHzPDjAgVmTcI72vKw9P1yxsysxjPgP8q5CNiP/5AG
Dk2duc88mRC8sdvEE0gm2e4L99se337XjAFR4giInWLFnu6RFT29qY+gtasu
K7wcLtDbx2BX262cH1Islo3B4DGdx9QLCB35Fo73e8pNU+RK83Aan737Idkd
aWnsPPLI/E42hPC8hpxAibOyAR8Zs5F4YUKJHYLqhGbmx30LEuhGGugXHzyk
YPDiFw8a4hMgCgEPQB9JS4kwKz42HbAge+jeC+8Js0cOBtI81Ls6Hizpz4wY
ARaj3wvwO5FPai9DVd4iNxuwfwe1CkteX33/pzEPUcZytU1m7oMB5UfV0K84
wP460KVkDdWsJ2HxfgDkL2l8ZhQubK9Vd31r2OlCsFphucK8/usWYHEP3ryw
LFgyM4BlyncyRSvl7ZfO8/77u0Or8xiWZhJd+wGsRN17VvXsDY7+2Mw89yHO
UusUQlh0Idg0mz1qsxy3RLAbjuEiby1TIYCTsxBxGozJ/XvzsynolhPT3igq
CoxRdmeQq3/eoVxTwjwekplFlltIoLDB2wHiOnXonLok7EDabwcIZwOW0aIj
tCbiQHVPKUKp9xMaWhSa6J5OMmqgBUgbVpXSpom9jmCCik46qDXMkBaC0awe
edMx9O3+o4QnEb1YxibMkFJAI7gWY7HyfDqmh9PvmedreS8A3pGMDLYeYK59
hb27gnKpCUVlkZr1/KX5SOJLTv86mmrgVFI+z9gP1nO56dlOFxkcChZrlqdo
DLmpEVt92Bk07Mx2UY4kfL4PGAZh/ASssIlDoqZnX5je8fxDDEFNTHXxkdEh
WI8ZVlv/fi7Hfk8XhdqmbsskRgehW99wvIBGpJSUrJu7/S9TzO/wM6uJ4F80
HZ5kPH33N/5uHNnx+60jRN/w2yXRlyOTemNeBnelvgGeiV4YPLwt5RiGQBTA
sRh2UE0AGpAcRpxN6ZouR3Lq9IDCrRptDJJPR5wnC27H3m6pg65WFuUsxWOs
FTIbDoS1f9+n2g2WfPIepT/H7f154frL6U2m8xQsWI+HB6CsHvNqsjZxX5+V
vuvtbmPKhE/pUTcmxQc5tX3zCKRtFSPfA0Ck/3lvQ0XLddeeNr0wPknHypiD
Ad97nOxsyiKLH4Y7CeMcc3obimstXm1S4waw/O979UxQUztM/jKM4qiL+Nt0
fV+nIh3feSGeb3dspBHG7E1HNjsK/g7nSNGhUeFkoLiG18pjlF2ucw3zPgZC
SwqfHnSi6K2G9LAsF7dJSXVhTkFvMekJvPOuQ5PpnOgMHGKcNwrp4NfokCVg
cVA6xgM1ug2hHZChOtWch+yWPl5DeOBi+U1jsLz67ZhvWwL1r5+iH4mU9aMe
BZbVjnSzwVPKal0CYwgDIy9AEoGlWLE+bZuufLeRJHwM1zUHP7P/7HrBFXPt
NmQubh19HntrM4eqU1TrUCm84aw1UpyMfRGxDRTlfXGADomp4kIml0iwBXjB
ir5shRcNBCd4CLApnRzLewDb8rHqrxmBdBiz+N4jsIL1ZHP745AHaRl3zVqH
jdi/CZe0cdIr+AWzz794I7TKS3yBafdub+u5vy1mG3T6AE7KoKlNeRawjVId
kDjCwV2d3021EzDaDb1udrBRJcTwXjjf5oERa/cHXSSwhJ7x4jKHwiUCxUPP
gmj6SsKF66wAJExYCBhQb/KSrbBluZmBU/rA4fdvwE6lHYZWOORK+aoJwsfO
euuDhr+agAME+Qo80wc1ICnUqf0h8DdMNWrNW1cdq38gVmRmb7/D/Gd5XGY9
Tq92kgstVMIAcKtU+EZK14i2wJIeau96rYFiO2he6E3Tt1LKrjSlr7V5iJsX
ZshwAKmb2n0f+wTq2tffaElhpAX1pEWButLzVxa1qTVN6WvWUCNpSCdRfDCz
Cna1er4wjVLUl7+BJuwoSwIwP2x5bx7OuP8sP2ogCN3xbAvfcsgt3co3u/eC
v8+njPzWPXmfb78xoo3qQZbIePedcLzlaPlyqLjCByTPHLojT+WMZv9UYVTW
4Z+BeJGwT5OSRhXe1+IcfbsRx51LH/pZlB8gtWAp9mWSmVv4+4OpCUFWK18I
fscAL953QK5xbIzz5smYIPeK1vaXQYW2eAQMUCLv+ROsgfkbFYmI/47uVtnC
4IuiGYYlVZok3cWs68rBMScbkym1mYqlmmjt4RfgBtYZPQ+jXHXHoEtPID0p
bu9w+i1diVBf2gz6AQvHU5TCW0LoG5pi8SnF75GX6hL+fNVrJaMJj1afwd+L
Xb8ULBnf2OpqRuNLmmTXndA8LqN2r4MUuX768EO3d4zOhw0YpvUwWWpf+vCX
ZFzxPh/XLfvXx76+fvWhcWE9su0qmDhRbaSz+Kk+XjnrYbRW8iyn5Oz42+KX
UQzlVzITO+vP/jJW7hGIMZ8MjP1JQ18GdnptAMBXqSUn0D+9vl8jYj948TQS
gN5MYZ6xJREZJVV8XEASMmfBq4EY1W5ZXjC1GEIUHmw/hbkV1KffhtEvxj2t
wZ1ssrRHsLkjgM0kih3zJLzhmkN3WIMvWcuxoaEDToDRsoAA8wFdG3nFKJPB
Ntp+H7a+OqALqhLbSDUPUu2BKH/S7xRjg+9+yN7DmbG4Rm/Oab4Zc2XQi4fF
fWej7kqfdLQ8XyABdYqgWPQ6N5swpfkfqRmWdsjwQ9OHDX1TAwW6nXOscNLm
ECFoM7mUrqn/BmpDuFXE4ltqD4DTSdb3nmVdMJ00z95ONxYI6dOyu+rU31yB
pb+Pm/7W0JD6XfRGrfuVPL/Nk9RE2bsKFwglweaGVaqU2TKRxf5JgkC0+uGg
3lKM4Mq9D/WYRlyd3aD+91aPGS68g12Sid46NkbJwybAr0hRTFyHmcOu6Bmp
I4lcapm4rLNR7pPq90XNT/NqeQrMnTWQidwbDXYBlLDw22cDFaObU+1rCIfT
Z9xe1GL+tQyiJ8gYSI4UO4t0wtBycA1FlkXxnQkLa6I/amDS/bm//6PO5V6l
r6yIcIg4SrlMo7fWVGPrW+dnM9pBb4BJnEiclLEGiTRoi9XeFFYhWTns6Y/1
qzYkirEJ+X2aklextwzy3JmFpwUJSiOcSm67Pd/AcfjzqPtXVNC1fLA8a5to
eZM9cyZqWj7c7k+YOkfshfGZglgusFBKvTIIlki3zWUpmMK0A/q9CvOE2vNh
gcwcd1y5zIcshRbV5YTYxSnye9xdosc2Xe8MRSJMHDCOgA1hkP1qa4gLLb84
CZuP7BA6fpwDx8jj6eb+ZRycfI8+aftQ64m5CciUYmMZQjXlif1c8u51G4ff
Yj5Z1tsRpKniZRjRVOOkCG3RqWDOmvpEp2/uFR8cF6+H7CA1q8lPpVsvN9Ls
MPrsbrtg/AJSJUdRInFLicbQ6j5F7izqQvfbxXp4eu1JJVjGPPrqa0PgPUiO
S3O7XTzfNo5MbmrbTZ3YC0sTHfLbQD8KVVwPEfgw44F2UWg9WU1jsA4yRqLF
LGrUdr08dNf5Qb14wLHMeyiy2GNEUTC4g+eTFcUF2FCUM+S8I4V1AJBV8nSu
RNWshPCskBJNTY/Z4fj48b+4BR7w4ag85DmnzdLgRJYhHDAyvWDOezbFDQ63
cJoP4tk86DFEn+VoEV6jfsCjr+2KFptUOoOLi9IG5h21tX7XGzTgRLNvAkyD
a2ft0d5WBvsqa0AvgseOY3YiKxx230aWoNCrY0GXXKuR6SGriQckBv5ZK0tj
QyALdtR3eIsxDwIqQVjei1EQKjq+Z+dcu2MpXxkDZMWNrxI6QGs7l01KWQyb
TvkgeisPyJ4GH0tEGb+rJSjmM1NzxGrz+ob5MOD8Ha4hEbV/O1A3NHcsj6pr
AciaeQLp/eZsGhSA4ltFG24BcQwg00efWT+1onHe6z1S8SsyFYJy2g+eBZ63
2w3AmXHIx3mOKWLsuWKVhE5OObhrPVNOjf+bRqM3TUq+326ANtx5kpxP/5XN
m6zl1XVuGRqUetFO7ZLwuWsaaCxDzoBV6mL3VP63uKE4mmptSpG9sGNfGWjJ
BtRBDLSODr1B08K2so20CSU1lv0GqC6TVCmQL7z36m5h9nB8nZhcUPGJFs18
TyuCLxCpQBVZMINminaicaHd4mRryQyhfdYatzi2TTkYRLVhGZNN2uIGfrJJ
DY2id8iDafNjgTGTEVVX78H3xjZHRBGtHVWQ0MK4PuAgmKNx3eORAIBo+Trj
rZNW3vXJWPzmT6Zn0tb9a8ybDTz59cG6OejFTW+uSOU1CqnFz9+lI0bjoUFE
tnlBPmLu+rIhT6ATmRwKqgcBx7GYIGOyBalsoBg2OPbt1eEXZ9R/7nvT+rr/
0JTAqsbchCw9wf602j4uC3Ybv8az+R3gk1pNl2IPy3S8LcOyq6KsycPBousC
EMNMooLc/hj8aaA7nmoNpLHk1HKlcl6aN6rUTIGETlIgxBfSrW7krzxbjB1I
U6b3O2spb+pEC/4xCB4I6cf5pYWIWi2FFQc1+her1n2QNrr7PdPq7ADOHDfe
sR42IDPKu08+3ENkjyRzqxAce29GRGNivFJa7y1rEnLIwMRbP39eb68W/2mP
+094+3rjHTChiU4X14+HQJR+4zq7TKJMto4eo459tnnd2dIIIoXmZZEgb3kC
5JcUbX9Nfb1PKXdhd+z5XpSOMsjxvFl0O1b4ltmin6QALgBAZYpoPsscBSXg
/xgvGbFP7Xql5Oa5C98QdsZopATbZpSI/UomAu3BJy9PPY5Y2d9Gt8H4Lifm
E5CKCRAbFcEZedMCiW6kMFOv9dylio334uCAXF0Qg6mcedaJ3FTCQBpe0Q/j
/NF7SvrBYxCb/6NaD8dHEeWxqX9I/HB4hY0qetcpAAa0MwA8U8nZar6mIeKs
/taAxpfh6Jn/0nk4ehv8BdFBcbUQq0KrmfFAyFp9a9SssZeNxUpT3XRZ4aX2
V8j49MEETjo7TDDpZtn9gHxBUcbvqbuNPZYICOJ3HiO86Ot8hkjlxvkfTHsE
GuP1NIOIvs/8sZZdm+dGYi23W+g9SQssJiCdxiJGq6UtjHOkmKM4tgx+esSm
iCYOJub/khTXJA+2ZsQ5yKgjfdrrpac4WrqJ1IO6UqCpxBUsiaulJRyLUu7B
hyNi/sXnSrfyma2IekgP9Xyk/cN83IldPhWeYjaDWqDwzdh4WB4W6Cs8Sc40
/L9m6q+IKmOc0jola/vUJ/GckNNWWjWU4P6sYKCYiixGCVqbn0Zo12XUjHAa
SFXVC4XvZBofG2Abo7S0B4DYENmKwJBVkAvznIVdVHiydQH+ajrgvLvYyBjw
J3u0fIi1wHl4p/7RGz97NSCpOQOyH9WVKzBgsbFm599VtuenNMrgrt8Wuls8
99HcS29B4UaG7JdXWQNLNg/kI1utB8U4ISSBhDM5S2jaEWEyaLZWo071PH2X
8WjmCDVVFvvPS9QzytfPlnptrgpTzZcWqjCm5Z6KvUi47M8zhO/oNovilr7J
EKW7N57/zWuCOLOpB5+HmlJOCI7chbdEySV5WtsMXZppjJ/lWikj2rqLcw9W
L9mKWK4CV3WBJyMe//nWQ2rKEoNy8guLmsJwkgdwpVUkOOE65Ogd/v4eqWYM
A4U3ipbGM7xiIbbvsi/LkkIEmgBgvWljskWIdaIVAI56HpHzui2e7UVSR2XB
eTD9ZtjaFufVCSK3SX7/yJmdpe/fJ293VsdHk0jiSkIBkEl+YLeRRnyGm9uk
fl2tUHgLYhPTSXITLcYWEAAZoMLRflVMimCsrh6KinvJDgrHwk20A5K7BheO
qhGhWFps8NGu7EFtzXPAFPR/pFtA0GxeO4ZAnczjMs9DCjPVJnAUKlgEGK5u
GejEIA+PQAwnGwdS3/DRrPdRJw1GhOd2okVj3xUGzt7lSNy8erc0G0imi/jA
Uu2TfmQ9KUld7VcVtlbmBYUXDnaXFglTZP1LcBCm/mrw4yvvU/cABddRmvJE
nn3UPIbhGwDoP3P2/k3sGQSaql4ef7Kf0FRryuFf+8o+AcCtG4b08g5rejZs
P1EAdeKbDCQEfeSq6R9S1/qii4Gus/ZOHFgLYhVPgEoJcjxvi5pvodeISzN/
2IWpoFK4QiucKhP3aGbWTL4VO1xASyIunBbBIRAlK6gX8075RgyScuknIN5r
kqzrP/hLrrgQlEnQ71VYZlGnE2lzZNrrefjTnARWxzB0okO1Y4tRFdNoUkG2
fsz6WRQiK/eSSem+mzsi66ImlYSU8m3HA4WwqRoSCw/UcI3MV+MoPwl8BqAb
oA+liihbnEXSVH8UnXGD9sBJHSOZq7Xd9GRzGTC7/KT9BPuIXG31oJsraJ4v
hoGndSeHjvaEgz+uq3Z0BpwCY4e0HCZdkH+PzkmDNTb9dvpOEZZVkMhGVajy
ydMkiFfIDKVqPXbC4RgfRGBZzunSkaw+v95FUP/R2KDkShRxBaDyFLLh+uOE
z2BjxCHbp+ayckfffeVDbxga7xFJH8YemDsIccW9we1NiSrie/QWv+v711AF
QLy/1obXeMZUmEQOGWxNEARaUNYD6XpJzWtXa9iL6K5rRa/WSn4ta+dlsPr6
Z1HdVDuMrSs4I6lvOzhkxpB+/L6xK+6gM2rznqF5rg4AgwCGpehPdEFayT7t
xo89RKP3Qu9xQ8rfGYpp4rbQhYdG9m33++/bzBgWmse6rFno0tvKkiULHV4e
lnz1UkL+DEvpLTGtO3JoJmuYW7Ir5x+4wPflAHafl7GpuWMuhkBuyjmEHC/U
VkaIG5Er1D9SYtSs8zj6IXn94IQl04/q+Yg2XQmSLppfuMcTCZKykPlmHek4
HeBc/AvlfS4d/0e6lp47xq8fWiKxXJYF1j9ipfNrY7ZFZhqN1ytu469OLMN1
eDeT21f4S2fooMLgqJje1dGUjSRLI/EQ0xcHxCGgX5oGEPG3nRDEMW50Z/1h
BLLovZbWsHKDz6u7yCkpz1t7XyjfKCkg7Fuflac8bC64+1LBiblYPXoJMd1C
ZF6mgoRkrWf04Meh8OpU/1gyYQ+VZjiWNO+y+N49a+cNqBL8MXHIJzrGdRA5
tdqsWCl9B54KoQkd2XHwlNhRagW5jirs2Pf0w74HWFRoq3ng8wJ+FIV6uMml
8Vu+6bdq6jJK4T3YHKqkO+pqA8C7Bb+bKUFCm1ZAoSdUV1aZs34ikLgumVe8
RyvbdrgOjFaiQ/YvCWeYpY5vGHQrhwdvvnHizjAG20IEdu8YtzLzVFAx+0xD
Kfby4VFAc7fgPpd1nUCLnJgB2GMXDUoOKjEDIJlspko52Mdc4Iz2Iy54dPJa
wbEihX0SfxUgwiuAOh/NbgsfCwUy+I3cPd69W/41DHSsCODfpK/hALohDsY5
FaAl5KRrLBoVGwlLTKgiGC1v6HRS0+DT63v4nqwyJFXBjGDw/t04kOPoBWet
GvN/LvhL+71RJ4iAcucNpAM3YBCa6iAR8pJy63ndW/W8p4jSxCcIM+8B97fl
cvekj2N6cAJS0zYqq1xYl/AF5lIHdYQL17exn96B/KPWEjYwNRx/9KpryIe6
mdD31a1V3KBkziQT3FfRU2rAlXatadxHG3V5de8etBzxxVMIo/oYbBaMo87O
c68jLmJ8LSQdmNE0qYSAChdmRpMK1OUyswyeEKGr1bibsdK1I3L8f5KTq5io
n1JbD9mL6PYqfY5vOW0lFFmPpm/gfT2Gg5uUGOxt0rgbTY0Gl5Pj6ge/XRXj
ZVohOBX1TmdedPx7e7ObJVZCWBxGw4BUwhVSNkAKIm/5Q/LFNZXN6OAUX6Ix
Toi/q/3BS6E13atjFM48gQZB38+vTVPy6iPwcVZVqmazSRhYknwKrKZ+kEvL
XFbliGsqoSGHwL95qwXCw5eTeBuVM+6YCatJ4IRdoYn+lnTUKuoMilWPrYyz
YTvJlux0JsjpD4xKB1DjmUbMD1BTAKb3YSkEdA7VVjrrpbGrcu7gnXYk4H5Z
YIrwPQH9eojIntDbN/1X/aciN+tdS4BosBTjPdBPNwlKHEPfx8n2ruaG9fG8
VhFCQZk75p9bF68o7gIzn5O9GrmfxLqzbmevSmMsh/lgwLfeVF1jDDOQEuPb
ZY2xdbOyfzwXLO2mRm+g52sIC95r9+z5AvVA+4Gpws4meDK+gsfzJd43z0xy
bdc4HezZwj4fZGUPZfylnazspjaPaexl+ZaFVt4jkUJ9iAn62yZhs0e/rm0c
b6O1eTZ8Sd37BMxA8pgwV8kCVzc8w/u/uj/U5skczR4TD0X6j9bDBCTg1jrn
FpB4if8Q47K4F/TgzWIreKmj3amnI3Mb2KzBJrD/vcO3CjDxTli5Sjtedqns
Uxd/z4X86KCblY6T1D+jyDzBBQDy0Msl2uvwBbB+EYjnGR8N21Hu7tWfuf5N
6+mM5wZnb2owU4jsUoyYB4C6XAivcrWWZFlP6IeUSELklBL3IqFYbfv4rkrl
gQp2nYd7J2BTuJV4Yk8DCV7rol9/3ZbJMpWV70/pqp0mTr7JeYGWWJNIk9Ub
5zO79vmN357ZsxAw67dz8p6la2hY+qZ5uMkbPoOuOkrZyiL43tIbvsxDCPwD
njJjTV8uC+PvPJQBhlSDJVDim4xQj28xRZhuZJXhk30gXGE1Z2RB04GbycmE
olFok3SRgIy72QfUz6MDVW0YEjY+SIw/DTRim+DxUpr4EqZsnX51K/K1Sd/e
P2VTy34t3M/vKUfAtS2nviCRm4cc+i2SQxKdOHZtNM4ygipbj0g9WudaqsN8
s6kAa6W+2BCjIvv070ayuhrse28Y3R8DKYJFSlZdaR+p/McKj+RB9x5uLmvS
XC3RcgTQpcJ6nCAc5h6i9iUMa5R/CEj2pZ85KU8uJPMuqFk/D/x9tyrQi0k7
3kkGjjbAKapV8g1/KTNROYtqRXtbVvUYKLmvVZLyujiNLrFQte+uU/qn9Hgl
5qY8FlD/tqgmCD9CtQ0nkDPSa7OSo4Z8LE6pikYTPfKGrnciXVe7J8BSOga2
MLdQZhkYmYKq38mMX9SxgKRsJ7NKerF+BJ82Vott8FFoXjG8QJsvlUOWkXB/
z4J2bLzeeqtE/RDLWUBHjjHC4P4sSVPN3koIcQGDrkqyRW0XXVhO6+LmrlGW
iZ+i++JBLO/XarcMv9jZQ0qvBDr75MC3uuUVZASmDWv8efa+T0so8P1odOyD
vrESPW5XJmNpfO9LMR2DoHuRxWfcLxjSX2RRF3eoOo2bfV0OMBEnwd+h4aeL
/xqYWG7uonvv8eddlf9uQfgJHZcWisFPtzENQjcXM/ckbGRD5jZnNYd8DUID
wsxl22rkGwrMSDVx5MxgphgAlneRdFSEfZE3imLdXfS5M+PeCCqYiQiWx0rm
tpvwi7S8JxrQAJjos7HqsdRMcUCPFtzjyETMrIV4onbeT3LFP45jN7CR3LQ4
PFg+poPMdnPb1hkmxHY+Axcl2dl4LAcPUoChdoo+l/OCT4z2wEZdCwVfcN72
QycslUefqwfDl9MzhtvFlULRnj4Z3e8cQCuSbIgIdwNIvmO7dGvQOjb5SZjt
w1PG30dQrG+17jhxBhLKbMgYil9oghxLF7D4pvQOKnOCKaDKkJXbLdVL9cLf
xguLBMvIEAvsqKzyVBugLPyDx5CWKyNFSQ6BqbeQY0yHQWjbvhnNVWKJgaDa
VjHVwdrzqtzOvILzcU8Fj9/4w6S0lzCorB3t74DxdezL1XwbM9AAnIHsgAqR
oo5dbBSIZPcYg2LIstdrEsFnH4Bue8OefbwBdxWZ5E984Tb0Z9xJ0+huOebm
Qa8MZ0chzTO/VF4k1mEt8GNvBI/1fCHYJ6JFRFiJIwq47RdwsfVoHhPwsvly
6qHXkLnHwMrmESEEDRcVH14nAoGVEpFyPWR/0TfJJdy1UdfU/8nE0eaX0KPC
Ey/OF7S0ACKn3Swx6wAV60ukd4cxie8CvSwRtERqvvnOSw7ylz1K+iTXhAp4
Yt7U4zLwBubibkkL6Q04ndeBRnl+6u5OEznsTH+rGSnZ+RLeuPobXKcqQpKh
tfUIbbfwDfUZdDurJKyyy9+5k3fKjO5oy1ris5CZBaImqEOFLx6OSkuG0B3F
Pi3CNhGdwaTC61B/ZQAt2eZPrY2FOvjDg3z+1jlghe4kvx3ZSo5jb+Hm1mbc
PNxbrrO4yqibUOL9PQL4QpQ6k47n2wczOJlQT+oEA86rxAAE9p6AaHplyN67
973EJ7UnFpR0wGI9HCq1pf86yUtbhhK6fnrLrvCCg/9ysHouswn0yhdnchJ4
fubBIz1eCzhyG7nCC1ClxqxL4kaj0EN6I8LbSiYevpsJumdmOCYlp5BQwGUt
tJjhLNZSoExXYx3DpicwzMYeWU6pfOiP9cE5mbGCSLTPrY3yR3TYN5WZdhPP
xGy/rdoBw5iESCtyNCbU+JrI175xIngB3s874IEb/o5eqhsHV3jnvJD0DCpC
Osc9KoiQ8ZkAoVwojNFUklfEBB0PCBwICSSZr6KrdBTNJtPhZUSe+AFnNQQo
cBuDr2fPP8SShhuypWO1tlGWthLiZFgXf2btU13a8qRg/gJML7AIFLc6T+Y7
beY737S6YgU4T6idoIyru9q/poLwoVRNfpubmKv5IC5Kr/m0+moT/XUx7e0A
iPbfnXyOAviwYB9gLTlqD/yqPMtq10DgFYXTmqbC3pmzXsHRNM13/g2kKbbR
utXhgX3boNPQeQ75FGomYC87FXWL7CtnJgtUM9ri/tvOG6MyzgNMg1QRv5tz
OYmFqBtNeFmVRAWYL8SY2CPim2U+Gr+p4iZ4Uxb3WZ7BjLeU6E2GAd5A3/1S
WQSzgsXCjsNZSLUcyGBr0k3G7nv0WzWK5OfKO5stFeZvIrpKFBd/SI2elaUQ
/fW7vZQH3pgdLWmcBFuovyngm8M90ICN8HoJTo4qABxwFxwMdkYRJi8R7eic
1xjQpEo/56XYxUR1TUMyK54pDKMHjhe9i02ID5G2sUZ0bJgwNOhJcucH4UYV
mpskrkrEgKD+cI92ZmjBzKSseji49tdYnI7Z7lJlvV6kVPGoCkIH42y3bxFx
HLBTG+u+tlZwfJaZFiBEt8VIJmC+P2va0Qd7v3Te+gC7R6k2GYewEbKoonOX
Sz63gSwPsfd/5h8XsYCAnCHp4UIywh3k3yKAEY1Alm8l+RqYermSSVwYToDE
dzmTZ+TLCRVyS19CO4+9qUyG9f7g03E8MuTC+wVcWbt6CNjNLDGs75i3yS9F
tg5xw5z6fm4atXl2euX9HpNBk+xSw84mS8llm8dYKtQPyCt2zcWlijFr7e1g
LBshW0LLup/RxumNT9XU5ZNyO4BEStd0chnZlsxU

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGOsr8kMFYOekjNQnBEhs9lyR21GYiOhF3vXFqT+oNI36NoQuwDrIKknOekZARuB0KGnXsx6ULpQR+iPvShG1Nw5sM+YgVPtubAz9+VRE624pfIQUwGSGgJK9rVX8MTz1/RMTs/9IoZ4tDZo/RYzUSzoGs41Xecckgwbk0IGySJBQoqJNZPXEAKk9V21upd2ttNOCV8QdIZtQPeVzXDRcxmH/7L6q1J3HxvB/RQeringNUuSa0XMTYLykYswR3CKaap0aI0TO4dG08qU1gGWGrxchRIbZJ0aZZKk8IwzJhU3fFAHW6Q3m2EjFa+0xptLARPdI+geKnIMkgeJJaXffw6qiEOT80upMSetgYLzl7KXeXoV95tY0t42+2AK8fUwhrC/66Mmr3bhWR3W6Mndi1V693oDTFlYpuqYTcxQ9kAmV69AwUEEtsiq6o/WjM6TL0FAOm172iHRq6/AJKpBEKvoAHY4WuPHDFDtC/3/odPVqrZIF5IqZkyJzxMFhbjszFHqDD2Y85NsyVnlHOgmGo/Qf/tlJinJcmynDyCXR0DUwafDEIDyNS00l2ssqH8YwswSIy8yLyVkYi992hQCZlrqZ8J7J/W8k2dLhJFN2mvX9ZL5JG8Xf7IDTcjBrFmHdwfEbPtDKWz9+2U0i1vXKczOFse07Amo55tqr74dIMpYb6o5dWiDc9Glrkm6wgVsUPxmqxxoAGxZYfVaXs4FtX6Q4T2y9i81a40Q/Yn2ITr7n0OOpK8QYPGfRtcgMHN+Tu717yUd3b3xMy/QvBTM4sFF"
`endif