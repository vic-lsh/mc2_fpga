// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0UA+guQTKaXQU83F+Yd1tg9asdOu/GKnA1IrT2d07wqQ4+bK9xm/u5YRcN3x
UswcUwugY0AKsQzhfF5G8XTgLYI2pqgFPIdyHLoZA30pKl8rd4kZuwoZAk3L
ZJ5YwyGbWZZX7uYV2WafmbR76f1RM/DUGTd6Koqg9G9cOi5k8gA8E4sotGDE
5/mJHXmcQ1MpOvIrEh7Swgy0nRPKmFiIZGw2+34Q1VFH+ckwS0EFAMh+bIUY
pckxLp/XSxOB5q+dEEyg0YAxIRYoE025oVCc8Eq16zE/6/dXGhebgrPBO4eB
fArhLV52ILy2lbhrotCL4XOPrOvzxbkcgFK52jAGLA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mWjKKChuKa8OCpXvuRSFsMHde3/joQhEltonmJToD1gaZva9Rbd+mk0N6owf
RvYwCNMu2FE0T5FVVzvpvad+AYDhzUYkpLGSD8nwIxO81Z+Vow94qo4eDviu
YcW29ESYm+D2iyqJzKkVuh7YFbw7EJgJhEkqXBHHo3QwvwyMJDUBRzQ3bJDj
+QdKjavoDY/gsNE6ImMW7QpjSrKCLMDexHQSCstch+wI5oEoieR2IIGF6oJt
DVQ1nKthiZ9JomeXI/TnJQh+VaVhMAhRc8GeJwFviMgikRa31YHc/cO7i0Qd
01egbTddJoO5ost9uzs4vEGZK18aZksS0ltJZvGcbg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qCeorZn726oGNMsDdbkekVkHpiWA1FUsOVttmkYdyNaYBkRreburkJCQ1ll6
WmzrCn3FkW2dmkGTVV44hy1VugzU4Vb/LhAoZwdlwoQZi85tZrqD43UjBmDj
GB11JHYOPwO98nKtLdoEbXUyRcH4frZUC/fnghSLuAVf3z2lSmfGS0/Qx0gp
KiAq3C+kY/avQ+wB1CNRgtWqN/8FSJ0x66Jx/0Jf2eg4B52y974XruzIAN2n
957nw693VWCBcQuY+mr9mFH4YEq+f0TXgrpJiR6uEH8CI7UcNMjQa2+b8fly
KBl77M/zuid7MRul7+RB9lasN1XqYr14LRoWYjUoXg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C6EdfbUAYjn5PVaBPw/Rh71/Aumf7p3Jw7LgGX7FuncqXiW43wbLRX1K/3rr
iUNbpOngqndKVso0YkGPCWbTgkotQwPn/WpHl6WAanynqafqlxxLWXPV2X1q
35sJshNG35aM81jjX/eYZx+O7193DExsfLlbXO2cba5BwCrR1bim5tBI8VsP
OG6flRRk+pVWJsFvY0g5HDkBEqIHKknoCCoMiuJuOYU+gnlZS0PuBjqmGfcd
X+hXTu6KnBVyvhlLcpFghh3OOJ1cxsqOiTsAPRcdLf9knAHF+RZjyzJxUqDv
o/B3a8khvO7yOCjaZOrCkJLwtuwACyVUYWYZcwO8gw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PFIPxzqW/xcd4ja7JuK+zl2MsReT2DtpgZGqmb3t8z8irD83egF2tHnCYoj0
OhpvjtUjrsb8MH3VZ/ZPgTq1w51okMdb4w1UUGrr5xn+y7ah/ykgmmilue+z
DJQ2tHtyjH4EqKLZuxCn0G3AZXlHaJqCjJuQJ0I7qF3DN4vaYrs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
S1RYzkASqzTd3EA51qGYdfy7o7cejmsvqZPg0I83KRF6CI+jA4BL8u0KE74j
B60QKpVFAb+TPTz0sH6cMz4Igtu2ZVA7JHsBsNCjW0CZB/RQryfXmY8vAqE4
XPcBfTXydu4gULQM0vxcYjbxqL6I2pjZMXy28Cx2QBGhKpKZC1drIXPU/86g
ERNhDiXw+sKPaoToFt0q/iGdgBrXFSL0qQaFOEP7Xcwy1uLBaWhhud4XM5JE
QcNi5A9w6ZdiYU7i9XzwQzO8pTr5szJM463raX4KbVln7lNtK9u72Ewije80
pg/9/XGfJvMzuj2ZCO64gEtZvslTwkQMYJtcKPKQp7hXd/FNxuSwX/dlnct/
dGMxGqCfcEuxEWXvUNJEWRmQwWlR2oa83cJz0Xw2BSXNi+GyjXJctEdRaL3W
z5e/03XDQcgJYF6BowcBmqb4+PEhLUKxwcUdpJu8jfchj7ZfdvLLrGo4jMx4
E3SSe9z0U+pb7nFvikFg2m81ZQ6qgX+K


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bRvFlaiiRg8Dh3zIOzw+H7NuUemwCHhIcDDGdCdMqIW0fmK1QoBsN9ejzt2o
vUczdEUOxpitXMW5/ZT5V+E2AE4nswbwDEXQOkjNC4cp2hNVaWNexB8SzU+R
u6ReA4eo9SJl0zrpc8ZnO1vQVJ6QrlSMcSHgkm2UqVFWvUPnxAE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AKSVetlDzEKxCtuHK2UCI+Lle7sxijTxNrrVoLSv8+M65VR9oSgqaNiInNkb
nk2ArAZ8j/f11RGVcRyLXG+Q2S69ojejJQUAWHBnKOdeKvdD2he4qtwa6LHI
if+84+cwLrJuEy2cSJx/OZyVHDousOkdVP2O9zWbP2MdfNu45Wg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9536)
`pragma protect data_block
sNW+rGvL7tq5RsPsSIdpmWsse5g3zL/Xioxi7ao1atNOdkWnVbF2yiS3ru8f
BgnXeiCJFQaz0RIarcdvLDRUFWKBlsIZUsK3j3xTcGxQ/2bstSq4RWYRoxpy
6cgh9cuaVkgj/qswemjOE8lpPOGF8hTru8kxbvEXwH5XiRI9E16S0GUkhzF2
TGZiSArgK193H3Nf7xTetB3wSQI/sZ1Yn0utMoh80k2JPpp2+VyjtqEiXLiq
R0s/yE9jffzmlt32u/ziwbCDnzYhG0oZ6DhNO6n9TWnxi0mmUlEQh7kh8MU2
Tq7c7R25P516CFor2voSrdS+dobH/g8bj0zW2RDYP6g1semOoSF6lGBe3IRt
S98zN/mKU4FUEkiIRFkRYOlTKwimIu4Dqkcw5wzqrsRp4lPF6fHCfFH3CziE
CdxHme23frY1dz6WA/uwXMVZv2t81atZls78/y9kyp50LEIAdOjZ7pB6Amu4
4oBNVZY9Agezpp5QRkhsq1zqpal22QXJCdwpUR5jwQNepqcC+46zJD3TkwGB
lZRFCXrcahVhERi7pCQ5ARFjhDMV8LGxp9gXYJUu8q65e69ExTFDbee5aU2H
T5o4ACvAeRqzZeAkNkg3ludTySHKk7EYD2SWpzUyemcYoaHzukW7Z6+vSaB1
CetBnYxrvd/2iJ4dSJ7ymQqiPC2S693oam4aSTKtUhhZ3gC9xGH2E2+95Mas
npr96lpiR9LDvJSljB5QWDLTztGKL3XT4KofZ0e58NhjFBfKozzUAKJRHTmh
YSBzDBgA+4Ic+3PlLEIPuaijFfbCclhtqqdRhzCA7on9iGYTElMX3ehsxF95
qgr7b1OIVcXPLICKgN/nx7f4fOkKZksux1d+jdRd6QmyzPqB1oQYC1PiJAww
Uk+Vf2Xv8/KYYJP3Uf1UwTNvdNTTYSTXb9d0pdnhgrKR0BHUcGIjoTj2JWrv
blB24TfKrcW0DHVcA0elBYE8H4yPgTGWvT2m5TusMBb1rCQL5DclXkH72MGU
FYGBv3h3hQSL4gEZVEERy458xznnujvo5DYs6pXLLnqSiZse0aaKuYfvuTCL
A1YWQeie2U1JqU0sVR1At+ERlfu3meVaHbB3q42ZYbGgXkrHFhiP/cUwOvfb
P3Vys0jckMuspBIZeN29xROS7rb4Tbq2wmt82xPFKLOrrH0ALB8a5ulT0hNm
/O/LUyTv5Mra0OEG4c8Bjcsx2CsxTLeQL+3tvhYzdBQeNj7uzRVXFmyxkjgq
3ZRy0ij5dnlB1zE5gcqwrcyrR3Hh9PdGSuYiFE3P8teSt8fXVg3pY7HtCvc0
w68gBkAx7Z7E6vjOBJcpHVSORSgPcujxqsCCGbqW2QkLU/6BjacVkqo28JdX
XsTn8oSvlwJa0uJiWrhBWs3azKqxnhOKl9w36djqWUinI/Pt0dYs5WY7TUpa
XxwdAtZBBncr/1LGgMIDZ8UAbSmiiN7KigVAHAu+GX3Mm1bewRsf+iGhqkWf
i0KLoQaLaz4tHkLshVMTjSwzhu5eiJd6wVe9CPSRcjxr/sYDJxGPTTIs07Rf
39P0rXtXaJ8XiTuXfmuokmpiM1JcCS6VXKvONiy4N6j1RqFtRtEF7dL5UGkg
HsTfThpC2eWlmyMvQ4s5hpTbXn08m7yGGfZWv7zfQ3FMKvjwIfqu8o+FeLf+
avKWysGNaHedG4MoG5WL6sg2kZw3UcoQijd7GzmKyUgkQQb2S5vWVdAPfk67
iA1LHa3L9ZHb7sQfYlB0ON7kZ0328Z0LWgO4hktLbqsGx0JezBALVGjCJnym
4LLwzT5Oqr5Wbxq5e4/3mldpkECQ8pWn5Rfb9MvPfRGS193ztmJ58m+U1plr
aTlEpppyuyz9wDeY6puj8vOz3DPo6DOnTfcWKDp1+AY70SeolJqXdekvl7Ph
wMlc5o32aLExmg9fWgD/A5X6AXft9459FV0oVqO6fFOs3BrT4vjwbjYkb5BU
vkv6ZbN8O7rFbRV7MSIlUoDCKyTtctnSf134/C18F/6Uebatm9tdd0o5g9Zr
fshBxAe9/cZ2MOYYMaONyRv+9ZPJ6DLposndbMM8jOuASWZm5UH9JampZqXg
NxeC1hwIRBGJRyFuYT7KS5BoEIBbJPeWPQbRXXknpd99T2moOGEdeK6JNhtf
pyCYgA67OEA+Abvt/bM85MkAp0hG8pPakgQCeAkTy7bBpoGZ3UlTEho+zdoe
alneDbONfr31zKJYai7oXTugxMYD2D1rRbbQ9Phtwk40MM5KNpJCNeqSnTTu
MkyIdo6pjCA7PsBQmrkVdlJ+AVEBBh33lzvEiDInXiwttFDtOeJumYfiA7Md
R38bcijzP5QZzy5itvDiSp5H7HVeGzRUqhxaQn4wksGz/oANtSg6hsjWgnXG
woaQWDszL9bf6+XvPUEXrBunm96BzUfu1TX2yea9o4RNfXu7f1CzY0ew5hz9
MEDEhXw6Kr3Iex8gwIAwiH47zsy7SAX9EO9x2t1JhqewTRFGzNAY1YajCnuk
SpLKs5FhdPkSiQ+G8rLdeLZ/hnnvs/nInNZTP+IwxyFArQQs2GkLEVx/s5oo
mNbIHXygbVu10qHOf34Zgv5uBM6bbkhe8ZAxc/v7sE9b3KJcoGCxqYsXWc7A
dQUQkWBqhtyjqhC/uYcYLx0k3RgkFOfj6wt2CqeMCpU2+CPbp+dcjAcJNboW
vHl60daejrW2yZSUGJ/QE3Lvr7+7BT1Q46fPOk+OrXuwSczJsp1MpjK53DW2
NNYNJcnfHGPH2NcuNkCzKrxP1cD0uFiFd1C+ineNtVAqBrOBIand1KrkkanR
x2m3jDOhFcBJwwzmI7VYtxbF4z2L8tMG7c59F2kf4wACkvSoyIjSMZpnfeyB
eLk9SZHDqGmYz9NxIDiT2wyhI1gV2SsPDy+Vea97duKZ8YM+MLfLc164w6Z0
uEK6vTfJbKHpLglHqY6IFfUaDatrDvoM1sW+PAWSR8E0kp04wgtQueAgNrA/
QxFTGdja8kyijSSqUekW3UhnKc3wojESK1VaL4frxmMgKgoz+dHmBVY4m0xg
T7mFbGo+v6lTkWMEsLg3WAZgy7k15kYEPJKHT+Wbd8DtCUU9vAIuzksuMG3d
NAexP6a0y+gpl3XG1M6XufAGAYAyNChG/+S7RdUHkNO51iq9O7a/YSRh0xPN
8aVzYQoA2Lkrvf/3j96DErC/opwncq4v6CWo4r+Xc/gx9zGcfh1ykMs0fwFg
u8CFIHykj8cp5w3POOdd1EjrKt5KQOIssTTgn73C3wmASSPnbov1PepU8LoB
hbCLqmFskv+6enrrv0DxM05S0e/FuXacGeQyty9CjEnFKem5erWZrxFsrL0m
7G03m+LYn0AwxJXq0A9QmwwzEQ90bmvyBg4sRVqJpqLRxVcIYGJrPOYpqwYf
qvta3y/auimda086zrNCRbDW6mEMTgQrRriNCnMcpUCkdHYS+Af799RcoAiy
w/T+XDw58Bf+jQnH2In4PIip5lQhQBmaPoof4yVspU7ZCwZ66HJ1XOo7k/h7
XUqd5rSr4YS/66PjvslufQmdIB2wlELT6zUfI/mCDdGv2vocPnmrSaBnD4Og
q0jJe5C34GHbmiT7mOcrAKVllTmjA2ZdteTRWwXiDWiIdZsTlLM/mM7fUl3/
pKWZgVHjxooZ7oDZrCEMizTb4AmqcOV9iseBQtMlVoGJBRJzgcsvyy9r9UIz
F0vvKuqChvrqy8WZLTFSycI38kjoh/heyu9NbccaQu7I/9/kEF5BYOjiVDys
A1tXjivFtCDmu2F9kiQdtx8Z9th22pA8kJpnYD6wZ786ED/hg3JNWjxBPlFG
inrHWQObEzdTALL39uGUIF49R89HvWAg8lWqy0CV2Pu6/noE8dZHQebzWSOY
RncX/hZw1iaJzzdQ0WkM+7m3DAQCv/uMeTXQA67UGrtJYr4VMdaPwfOMsr8h
qJWxGZalMMqR6FghMXeesb8EWDKs/FxakvJHYhmADvn3jArAbzBQgMvsG0pg
QIBH66vIRPiN4jb8LWtti60JXCAkSqgbZ/nIiftRQIxnszfoIqvkZMSMnNTo
FAV7/egJJQW49WS9s08zl/yTHbn+I9jLtzDIqNrPVidSRmfllDtBtQM61p2x
zJb+yQ6g9MBXxsJxsn1yhDTx5IemcXnJgB7FjFfPBfn2Tak5T7xT1GQaV+WX
7DkFGWpdY1VnAZ3S71beaBTcLEFGqa709gQ0qcmLYnZxF6wykyuGyqZrdqyB
bS+CJzokxvgScTl8oQiXOs4daZVfCEmdNF6OHuNnJdU9KzypSGKPMt/KWCFK
tTC2/bfMBTu7eBGqVHn/YOWY5jhEeldVwGa/CbJrgaNOutt8aUGRMWp7Hw2H
Nqo+I9kheyPqspDeknG8QzcuPN1hyGzkh34onTT8Jy3urT4oR2lF6QKWug/G
Mbb3Ask9UrB8VMSR8i7TPV0hvEjXIMwaCJmQL4RCgm5Y1Hn9LgrbMx2JBTdk
DgXn2Ea4LN8lV7KeZFJEplxcUL7Ehd1aHOayD+Y82yBRzLmxtHMVOFErCnwh
4vus0X3QK4ffS9lricw8OV3jVqoq5EejWb29QTI00Won7GBlAot3muVFLg9e
k8+sLkrj/7EKBn84L2FztkfjBfFUHjDGWjiDW2CUEn+gkpehKjPqCUj/oNZq
6c6u5xrY7HVEYmIE5iGDKC3QnR6jrPkL8fnUg8hr05fUQjclR9tIr06VQoMW
ocDTjTtun/Qppv0IEWNPzfbvgTNWyVDhIcW57x/DvavWYFIISVcsWnvqlKv/
kFyX7JccMkeJsTC9YhfWClk+qDJplur2kVNHpe/DLYZ1jJ/v71W0Ebnq2gmF
IbrJuVV2+w1622kEp8E9rUykw4W5ylNnX3OjB3cHwXOjy6AZHVS029s7RQG1
Kqpj2IUAn+rGFPcGhEkVQZEkjNmV8YM+F3Ef+ArtoD6/g0Z4Gk2PcRXsZMyC
ai9DGglPCBUGwba1IaBQ6cdef424nuXb/Y5SUqTUyNPqSjD+RMPTVbj0b5lp
iN0YnPkq9SjNnTU0ytk2e7Qa8ahbN39cYYP6PLWXxZiOm4znh56UcxcoGDi9
6dmEqgnYLvT4hByRf8BHje5WRATlYNMFa/93aTEydBA2GeOiGfX7iMebhwXB
H4/1xGg2PwMOXKHJPYMSMo8icCnwFAah9oEPoot39+5sK8mfzmj3DHPC1VZB
rAL/jGi5YvJkskxeLVPZWxcsprQObRwVDGahxGlYySQRPC19BFUx4qDZb6m0
aWx0XTKSNaG7UXSvvTc9BcTz2V0BDWtVcB4Z+ym6VSGQ30n5xLrkQyVqJlgm
/VSv5Bo7Dsb3RF6I7gl04NHDHtBftXvZQO/ZrX4hpC194gBoZFYOhJA4sMSP
V5zf+eA3/HWPC+PX272YVG40KIaggo8TKYL79A7AqPRSv8pCYLjkwoVKV+KG
Odg7x4SwyKkbUDT3nOM04dwsYgZDVUnbc7mtcNTM6kMkBKHPOrqyIolC3uBl
wm+MvznyWt5o/7RLjm9J7TIqYBfhgNKQSUggk2v+2JL26Do0v6xtCjaN0Zf9
ILqssHsTlC1FPKV5WL02nwSFMK/8Z17SDcnhWAI833pH+QnYl63KXBon4eRx
OttvKaQbd6S1RN0SXiGrD+Yop0a8krI71Q30qQCCfpYHx/bFVzgR0vPvcgS6
LJ0nCqgaE0HzctVm5FXPXhA4UiC4RKb91xgiOH852ffQyrkkOKpcZpk5/N33
8riLeTdPYrogALoLaZNN/VPEuEGHumkyE/+566icxANtnhmyoM4108AOSdzV
Q5GS1cLS9YhR8khAY/ROjT8tkDyzop3SVw0d/GDX9Uwbx70As5hgqhu6h8Nh
05RjOls61thGbJAMpu6ttIuoPbIizy6QA6JVVq7n0dXz4lOFJTZxe/mJPGCa
uohVw7xYtQ4i8eVzXHS/wl+CZUnRwn+3/nWf9JHn5TtL2+iPurJdPVU/EMJh
tzAGFpqtRYW+PlLpeptUYWFdVyP2btH5hoUi8ZSk1JZLDZvQzoHWeTde0SVu
sZD7EQ60NlUURR6SnVMMR8cBH8LzN+7P4p2ki445DOZLNXO2S3c23jbVOBXp
nyTibzmexyhHsgruXm+PsLRg5OWBwSZ3jZAgQ53jVC1yHqJcuCULEQFs+QZN
84S9hXMBVOW//vXyc6pInsTkAk9sBi/yyuI6G5kOT/t651BbBzv1qxnnuqGA
GPHZC/A+G/2pax67HyowFEPbszy28BKXzc8ffTjyX/Gm3eA64COW38DuWUwF
O5uxS0uHqtVGsqbTHRmomviScqcMMj2ButaXk2gNoRfUT3jCnPvmFkd7FPkV
3kbIcU7/Bx9vxIZjDHXbOgc5rUYAd82GLQkx/soPbJ/l8S7pg8Eonc9OZHhj
pCJP90o3LmABaeDuNfQNLAVjnch0X1kpOmYxxaWU4FtGw2Eio3WjkkWnC5Cx
0gofLuTNidOQCuff8T864+KhRdUIYw2yn1U2y9xHMeqKXqx3sUp2ykkzbHeK
boPIfmjIoSdJNPkMSpkHU/85vH0fq3znZ1DnBGMe+yOap7uHn7pCIYuwQCTe
KZKn0PDdveE5a+2wOwWg0xpZln32JLxqvaYrhY319CVJkjlIcATmrNPWsKFG
eN4hCHVUFbcDwA4mRRMXLNdkAgKPzHFDNyXe9SaspCUJr6l6cjFRWPdbNQ2O
t9vuiBIOnqkYm4AyKSfe+5L2fz+YkjdTTtAiBNZIEw69lNy+0m1TzE6g5Qux
2lUipZK0GSijhuhibnrkjIl5xVDyIj3iVyQiMSl40B6kChxtTM/PRTtlcNov
DDB7P6TF0IJ0xTRCcn1Y6SfTY2+kuqvKfAhB8to0WGrDJsDbvFHef2sr8Ddp
OhiIwPbtOGLsZgKlgymsWoo7JS7ffWgagka3wHxIt9lZEoJRvr4778RozG61
EUEOZknxCXLdrlvIIdLdCJnChwIVv8ouPQw3eSXpoNq4zurTD7eb590EW45F
O6UI/CU6WqlwrBCdKiuone83NBhxrAT9G81iZlrMTmVr9ZdtIhDtsTQAw3uu
a4qhbVaIMWsJnXhZVMKSir4XfwT//GWOH7ix0e902Ko/Yt25oQKphwAFZcaR
K0qgsUVH25P0ABoVwFM3LEf42hVW8OTrzbe9Wzf1OeoCD7+WiPPRb27+i5ox
QLHFMGRMv0FA3wXdBk04Y8mLDI3/7uQ6NAgkOpuHCsS6JZXwetNyr18gMj68
PKVa6l5F9vOwSv8gble1w6fhrjn7ItbpCjcFoiBNd6B9s2Qw2wOdEjOxN8FK
cXSNol3AB5VaM/4PXKcffaR6bFKx+fga1O9yuKZnzfZHEjEkBSDXhuFf7D4C
2oVkpc0HVsGshacLrL4rtliiQhqgqLi54GHV18bU8HTPNLFAji0Q8iIXhmyS
5I9hSRtWIKoVtdzcpyReOfXQQn8dm9Ir7BcJjn1+XDNCTTPJQBtcf3OB9yCc
OLsdALSxDoX37H35pCUVY4vSL8/6daux+GIP/hYF2HRbREJmCj/jxTFRkjOv
WuVu3PGkxi93lqy6zXTKH7Bie3jNQN0kz17Pm0ecLwVDgGgp3VR90s70S3dT
LqOJVgJmNAx2nwMW3O1mrovsTXt0/c6tWGMX+84ctoN0gOEo6bQIrtnHDMn6
1LmgfNj9y7/CL8BgOO2Ij9PqRYPpzwzBTFVCVFSvkdCXHUMNzvV6v6TUu7O8
bnU4DtFU2vTcUlATGbwj/uT7jOHI/Kh6TRHPnGg/R3Go592v5eEU5SfJOb3v
CPmZZ6dTLqyywPQzahH2ivghru/HEmSAP4XEwCv+Oy8hPstxOlsVNjBzjsLg
EgpjsojhWwo57u6BZwMpR+Ap6B1mY4ZGcQ1SW89P7SMliNRuyj7cLcOGAdif
F+aN2P7XYHL7fx95kMCC1OHu2aYgwhgPNnxEAaBOv/yK8vQrcVVHpvOxJ/t7
MLhp/H9qqSunFfT0ApFfEvwG/2npLZ1lM/HskA4WCFNjvagB2gwH+lX9KpbZ
7IKXDQ7wNwvUSxgyjj4GcV0d8X6gCamdovep9Liv/GS0SqZ3gpUYWPA6ewGX
S48MS1SEBBTr96NmUybLXEGwJuvvGmwAy2uhqoxt9FtTjO6/o7Z1+JVDpaL9
406Ubno6QDlEgdKXLNZIGnVdeRkbkRjo+928of9hH7o+N6GBpveubtVUr9Px
f4hcDf+Vwik33cGFIUThgH+1YJo/cKxBwI0oRGWB0JT72Js0AHPFRmnguhcb
Re/lvWB0P9eV42StnZoQnJOPzaq4IaRqWfTQntBgc9tPtpbXbnuFpkt+DwND
kImDYeXOzg1iUpzGL7YIaLer2zjyamSlbrNhnN9D83X8QchQbQj+K03MCVPd
WRKWgC24esp/RHOGSwFcocBsyp+axCnf79EySh3QALJZHV95QP3gfrm633n8
FaIj/51olaHPTsm+0m8PrebgZr2k0hMf9ZW3KD6TroKKO/FSjnVeS3E6xhoj
1iN33bYMLmQW31+37/XC2c0mYhkSZ/SgdLjNVdMUocLuyne4ntybhUT5qibv
reTZCBoExtWI9MdAZeACMrlJM2ILKkGNMN5yQ/6aFlVskCZsQGVv15ukKIeb
0fE/s6KQumx6buxPVdUblxwIqAhgU+ABZc5Q0Q3ZBiEy89QfOf82lE7R1Elh
I6ku3g7CFmf7cEleuE7uTaa8Er2qRsCoSu+9WdfG6J5CcM2Zimd5K7mp1lzD
h+AAsaTwKFDgS5dRllrSbdgCm3lNkV436iS3qn3TvM33o7rp0G0JYQ1RNcbF
bYprJPmCrhs0Uwo6Fy39nHWGI+l8zMGB3EZ5RqdR0WANwvV3Swg0gTfT6wZ9
qHRQc3gHMOGBnYXfgi1RTybf6Dtto1cKdzMUSOo3eJ368ZVgtML9T5Eh6QWl
oGByM3JxeWRq0pcMrk7nax07gU6bOR9WIjgb42p8vGN09zYeEXE2kNkA2rQh
F1v+z6i7CxWK/lpXecDElrfkCrhzuycTvcrsiGB5LwFKtQzy94n2GUqZRvAi
O8SsNnp9ZPnKLD+TVYz9DnyUtDLd4+xab829w1Me9b80H6Hyins1GKrJ60uQ
J8yZcSbnZAh0bv7L1+Bu6XCdoxzvnN5HVzoJqmIEGZOKibjgx7xUsbRMHEc9
rtG5HPIsQCr/zPxITihFiIScvbA8FSh2+nNU+e1V9BBQ2m4OdJUY18cpZDBJ
gmD+x6nnByDpc+AsEA/QppulungTylH9Hem0ojfQw9giz/Iy7LK+LRaCXnvC
/k29yO4Q1TVxf7tVJGZOA7teVr/SQ57Ya6VrpaQmV3txWkGEVWbugK8HLKxy
25CAA1UXlXt+LvPA13z/HIukAxy8si3WSJihRRsdyWGREnfEczrzwjrsFxFl
1J0gcw6VH6Np3NeV52biBzPHOe1emfBd1pM6dYn04/kTALPtPKje0oZirJrk
ka+k8SiPy/0E7YepBQ2Ku7hdU4qKIy3dOFZAt7lyzXHbF2eHhT6iyRFijL5r
NrLxDPZoygRLBqeaTgr059VLRzY4iu/RR7tCEk9Vk9mLsPuL/VxCYifWM0ID
/K7dKTn/IkVZ3GORGmvkeG3NOZsf48jOrUwpqb04VBDB70y0m1RzRhPkdupQ
gr/bXIvp2UuNPUO9oB7UuA+KuM95L5X1BELK3TprbseuSKn5PMiNIxmg0sSc
XuXGcMaYzeRtengd/TVT248KQP9S1o0Cz0DYeUegLfavqDdiVWzf3NZycq7m
IqpjvHllJqnIYWOxoW5WJ75K4RcbI2v+6MzL8TWW7eNM9aWAfQawKdXO2Ath
lSl8vG4vFAy5KLSAlQaG8AB0J/Cc5I7E/eK37F+zqsXew3rvzvHZIC1fChBi
PVoYeYi72vZ7V/o80D+R7fVUV7VI6zB0yO+EBsEvXf0NyF47J4KCQWGx2H0K
bKQVMlbpUFJANLKUZ2cY/bvc4aLmh36bYC6DJggvwyqAeS61npfo5vrpddIt
+Z75WimV/EqrzWwhQxyEPbwDL1b8UblyMLQI4RarmB1St9FiYdEZJVUJ+64Z
uPTTeR7z5q0jw8b2a39zNKcn23arFwU82jzYHBu2zpkYGEKY7v/QyKUX/STE
h9JI9NNq1zObv9d5DpVyrgwQktoyyIIks57jq0Z90UNGZ0BrJspiR5Z+sRLF
wkwvVqcfS2mlCNY0ttZ1H3eyaVlIdI1QRXODrLWJKcy0xHbW2BTMmSb7mGyU
wr6sYpy0/5+OylhdGakho7wCurUYWnu4DCJapIYr2WhozNTk2hAjugmp83ah
358atF7gF1j3RPZBcFEHlx8zZZRV79eB5yF9U/+gyJ2y4ExWx6bgpa6QZpd9
UYc39I6MqOwCrvciUSGURHBLXM5ZqLBlzM62zcdHblZAUdRCJnUtvACl0lQ+
T4bhR508QWGaHGKp36dVUZRu9JXM4ghQS8z9shIZFBZvOwurafmJ7EFjyAqi
SoVVd2PAE5WEzC5yXbB+hTMbiFtls37ZMtK5l3f6XWsfIF4BcYv9F4WxTSiE
cE9IELB7J5CD3puHwUSJ7zZ8efr1EZO3kpuhYhOVqcTrh9OCUo+Apn1AIjIO
7daxWNxHrdW+x0qbGuPiFT5EZgC4K5eKHMT2YO3jlzG7ItQAywgIjzx9sH9u
eyeWfLcCu2KZ4ajhfQ60wjyxhBa9/NWOILII3sW8314oG/kJyYChpixy/3zU
OgrZBqCCVvmMd/XdUoaqBL7JmdvOptueojmcQVzt1xXDwfMdpg+z5xC7iP9F
7RGNpQOjsKx9sOlJW1A9aWetDuuIjis044syzFAtrU34YBNRBWCZTuBcRkGR
XsFIxA1e0lRsWUM1ubG8okAJ+ANF6k47h+A+dNdpG20qccnK9ZXGt3uZbxZH
eaHGYaRA+M3ByH6cFoY4s8/cBNKFPRYndejlryxH6PMVifBBitqThksvAqtE
kXcvwDQ+yE6Jf/E47jpUurTFNl2TYTjX2H9m2heM5ydhbfVUBt3zp0dGxqZE
+WhwuVSeDpLQ604rZM/bCGkNvfUH86ZvwHnHikowpuQ68jm3uA6vg2ibXMav
GXU3VqEv+E2InGSYWZBsOCyhp2AES/XJiCaMSZEHhM7Co2vl2NGmPSXqNC6B
mB7wi2mAFbNA/s0lJPs6UOpACmsx8EWhTT2UqbirT0kJlLNidToL0DRz2LgG
0W/xiGVSnGI0J0NAkaVJs+tF3j9iArb/kvsa/YVR3iAZRhuMdJeEX27ZCQsY
4Y6NRYbxLvqwJIEmHT584OAnliBRkhAND0lMiTU3PjBod69RO5zBpZgJgJwR
XPbnpA7OsNDfqpgzK1ngU+Phn5eHhP1SfDSg/1d8UmdJgqrr9wYCWpYIrU/V
GG7MFs9m00l0K9UZmYP4ebAAQOWrslpi6OigpAXoVbkq72k/eA5XLsFQUAL+
TJJRHBKj8P++YX8pMt/G4AhZrLbZPmZ/rWJWpod/JN95qdVQB+bBXCeE7nDI
coxVHeWwSD9lAAnuce0yV3CVd2OtJRkck2qUfH4OiH2JhaKkEr9Rbe4OZzAk
2DB6aH2aEGakGEdO+2nutlLc3+YaV+Zcc8PYmr2EzDiUlSj6n21ooykApru3
ceqlwS+GkThBXJDj1dSvpymQZaen3Ky1H2nbb7dNOC8HS65q4YO4cjXTpwBp
Fj8JMGmvySBTqnob4YxZpeXup85cbBz1IfBbNEbn6Um1oAwpcIqD+/pd4x7H
lV+UxblJx7mYIg+GMDeMCM9w98/+tKch4nnjZ3TD4vmnpVwVHc9z8udDLQRL
n8XU3zIP8tmSFZDVZ4VorDSiEQR92fnPaN1DcNCJ5l4UzSnOv0CKUIpp+KFV
rXIXpapMNlr9yu/aQJZ+lCNVU5cFUY6EJgsEBub/Zp6jm/w8qtp5mESO27u3
9Cz9TLElbw1p70ugav0ci09pRXG4CABmc6tYzTS2TQTiXuyAUQRVuBw3ds9B
bOhQsk0sOK2E7xf6cPmySQ8NRwsdZANh5GK1yG3nDsryyH1Gzee1Z+F+sza4
pKtvCNGawWYz7wM5Jw9fpc0zMl4jPmEyI8wnp7AZp22WSr5vb8/UzvcQ79ny
TKXg5MeAA1AIQGW/Ati5Lgi9fGcZSz296/+ZRmk9wM3S74yWJwOEh6Ksl7lM
gZBja8iPiRdckw0xktfCEW3O3HKVUTAh/2KAXJDw0gdCQkWvYKLeM8dUV4B4
G4uvCVwiP3ixoAk8y4ufj9eatyGV2xhjRLjStS1KNx++Z30UsrbVkr5sehVM
U5xQdZkq/iS+0la5pHW9ypu4U3UxcWLWmT/Gx3mXIHSvsfkGaAeKISGkzGM7
GgWhaENA5qT/pcR6Up8PJT14Uc+DDi/6680XYptpMuxsV6c3cz/LfDmnJgpo
sChtnNsNM4D3C0kVp85iknSs+I4I/Rex/Jx1/E63KwEhB9U6uxqfjYKY3uER
7TOErJjZlet0+Wwxq7j1N+gS0j3JQdbFXn2DcxAfo/AAq/jwa+JZkRsp2sO2
NYBXxoLS7/t9uXCQOg2JJwuUvNOiIGUbcYXqWw3TTXPbNmkn1kK8VZhw18E6
xe65Kz7Ll16V07wUMuE7pV5vGBcUzYZaGvZ3h46GLxuEihQJBC0AMY80moEV
iZL4KaoDE2P51Luvgdw4FzVWFfSVhyKsCWzBmGSQE6rASCRg5I8YZgA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfLNS0rQG0Iz48Kx38OFyeRW6L9lHRWMbucJT4NosYdoBP3MOA0qFI34Wou2KX0PAwRL/Z9pW70AD35dIfDMe+YtmyVD6zA7K42fsQqcDspbZq1vN5E1iIu8ewwxbf8nKIiNy2DNYJmvMSFaR1g72ED2FXC5FKWgfvDDUAhQeaOtGK1OyGC/pJG6hQxU+shFI6++h6U3zwYbjRDQR80A03dudJ6OT0DJ3SIIdqspGaoqvXjC39z4f9SWxuSaQTtfsnM1m0NV8IjEnqraLGFTDgXhPAnH96oRQRfzTZo/g0QM0BMP16SiUNWvsofBIL/bC22adJLpwq1IrwZEgl6Aak5Kr47G0BVbnL779id1fTL8/KsCDJ6ilpLySJVXtLPps7VdVzY9xgDnUHb6OCR0w+Owc5cE9GK6PY3N51Gf5NKF+cbgm4KdWqBEDy80wqa30xFuvopd1ni5YHlvk6O9sYCajSWJx4if7Fcu20rMWkkAayLvsxR1IcOFMFYyzJjOsRRRCvRnzvkWNrjW7Pm5EzwdI0yVlHJjwkslJPn5U1Ll7s7Q2hIyY4exLLI1k/Xq6oH05kQAEhRRritw0FJSUXQcAlcO5kNoYBZHjB/ML+YmWXtPddbwZ0hs3KiwrscbIW0yqWnAnBSfCCO56ALHpckmggxkMJxm4Vzlwa0bjMwOZC+yfBERUqN7y2qEQpHJ+d/ZSAjYUwnDi4UdRpI3JEjNnSXGW6ME7EvwswCq0IJXHkJNHV8sJmSfutNhqDygW6nLgdV+uOaId4lXxzoQBTK"
`endif