// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fp6qZZJE8h0zkA+z+9GNu5fSHnNjVM0bNIYOIwTYSKmIi01lEs+MwkDZEqjO
nv0vCneuVRChjNJ5EkGT+RAqmcuTfN5r7h/QmOdBKBdkkOCJRp1DcBAWMtw3
9fMyAOCdn8iZNaYNRKToHTlYnyaWhLQl5i5JQJSe7si1TCfa6vP3L9QAYo2V
hpDhm6AKQ/yD9ZZV7yxulleeQn/rOaxtiwavDeChTYx6M1c7o+gHThUUp4MV
GzPrn5YY9rikjiPDbJsRaxW3iSG1inN437iKyAOgr0lAaKeqiz+Fj6WSFzSs
1ktVf3c58zPpWjWOUEuowZ+D9xoS/cWdt28hgERsow==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K5IGr1ovjDatQDVhaPsNjwtNF9mcL/uFrt7sJWgflX7yIldNhMbmH6E6YME/
ngUXPZJuasaw0zcRwe7FkjdSLCeqscVv6gxiusfgh+mAGkmJFeFrFktiRixV
grhlTWc+qXqnK5QSEsyFS9F2etLvAh7e57KvUJPpQ7ItZ+hGbZtsHNVWWTDP
fi1cxeppV4grplgyLDlpfRTRk+ILd8rzl9jUCF/hM+dtNtt28KTvP6cNlRO3
TEQ5xlxmUi3joYufURniJFiGtOve/kPNOut/HUnumdWmrhsWu6FfUaoCGlB8
7ALWXX8hjwkQl+DrDH7YTqyxamkaXWefO5jb6oz7eg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hyv66ohCKHt6Df4l8TaJ2NN9/l6ZI69+Zqasu/T6NhC05Ftmba9IKSOoFLXP
VxoHQkxmZ1Xcxj2isjaT0AN+/R/VjMCuUkfaeBessoCcMFal4edA5RL91Vxo
A4ipdkGGrH9KtKAnCWQ0qH3reGAacegGecUTpqsnyrFH4K3OmZu8KFP+kdgT
eMGbyNrJzdaoc0I+tOcYyv5w/wDrqboD3ztw4OeETcbHESANfY8XTWgmxKFC
46SDw4sOCgs7bjDoJRAm+2NT+/m5dLBOq0FpO8Pdl6tcCADmlTMxa/K+QMhh
5faNFdiT+7wG8jghBOtdPOK1R8SFsxRqROVIX/WVBQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MNxGjktMa2lxEaeDIRUAgjqI4obJ3l2Bb5BO+i+sA4mN7+r+/iNMKLeBGtNS
lqrZfhR8EwEr4bc29GtP5k8lRpaB3AjAN4z/5a8eWzCcvFpoPYUJBUTL1oXc
bccf1rlSqRglHh2P2dFiRCTYshWcs3/cBItQnz/Z8m1AAGqAJyHPHy8E5S0Y
yz9lF4RZlS5q5JoYGbxoosNWAe2vY/52cbLe6p19iYiWl5gk0uq6Jafp4sG5
1nAwTkzr2gu9aK7Lxg07nYa+SAQtLynm+R0QKRrxusOynZBvuNIdKVEEvewz
TFh0XImzsrvRGSs+ovy02pwnA6CCl3kIF7qRgO5Ffg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n/get6tjnoR7v7wvRx2z7ojpG7bF+tVX1qBd7DIxr1zQGLUydIyCP2ezMibe
fB6ewEfhVPno8b1erNyOClPH97owuOC9gcNiIOhs3t+mkePSSc1vB6pLtqHV
ESc033mgnkxWEPqSj9Kt7Nzzm6bxfmt/c1OBve9i3Ziv0R0U7SE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DM71kDpEmSwvwLXYCoghnx7ecCieUG9+XLq9njcxD0jylVcwL0BzHJX1QHsr
Dp76gZp7bEZLoOVNJbUFdZ4lr3Zfi53m1Buf/HlrpY3c8dqhwwdlKid9VYwU
8ofHPJM6SssLNVNsgLpZAweuAKPc4PGhKLdF7i9b5WUZuey2rUxhqPCpNNhw
oPTJk2B3XEu2sR+QoMryfNA2zV7kPRI1f7pyOtz5mwYDL6WByM5VLpgbwkM0
wtv7pyuXseDedZq7V5rfUpuM51VNtU/KXOO/Ig31Jh28+vqXFtw9sNMGovnb
wcm8ab3DCQm+E5ytYoJKS353cv28zN4w+/J1EPKH8aggupu2U7m4GfBZSmDb
5gvTNh9ZTMglrMYrKL3f9tySli+9P8ZEVbqb85IoAdH3mII385VtcDl9b6KP
YVQ+xqnQf1JQPYpnXWt973OwGUD9tp9Nj36gSxLcyN2GHEz+wTGRNIPJ3cL1
u0m1A5edx4FhPeEU+3cL1j99Cvnh0iBC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VQ0WyHTFf4asNKZduFE84WcRzZCPJV/AkiRK6E8Fbs2lwSEORZUAHuBdtuLS
vsEhaAj28//EFyYZdPRWIOVdnRwa4O6cjH49t5ZwVM9LRjaf+/PYshJaQXmj
oCZEm5/nPAgbO16VVTaoFw3xSk9VyO6LmCLUEPXX/JT7Xkr9H8Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mxY0D6T8eKCHexITyHkgH9saPf3Fhx9UMVYfGtEJgX9PklzEHq/fm7m6u2VF
KPirVc+twAV+PranWfduNV35wy7yVdmnTU+NPji09PVFlquErgJBH/I+f4vh
AizEFIYpV5MfwWNZ6lb/XPjnB3KM6NamN0mK2QSfRXs+IfMvYmI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26896)
`pragma protect data_block
kd2W4+DxhzRuFdlpLj4OrnJJL7iaw2VlAIK4cJjP51OtNQRBpQ7zPnX7C+zH
rHKC1NYPMoqRHo9a0YXhF4aD1BtnSpXsoOs1PL4WS/UD7457evI5iJdaFo7j
ZDyH2ybu4e2YWyMvthddqvdnI1ZcWlDkpYfYlQpk+iSOFIRmNJhGeAwtp/YS
TsFuJSoBXJd9iPhn9euhuLZpc9PrtEhczrskAfu19w2q+kuLRPA6ptqlheBn
/rgOd4l3hj5ibOr1pA6SrwrTe//4jP8Di/JVt0VQxXY6dz0CknD1w9wVCwF9
DxYbKgyj7d7G3lrpguLZlmwgYzYtrq3eUkbszZr8WoCK3/kPPuVz6FX8xT+C
QwB8iPy0hfYm/qEAogrTZ2yncklZGgxwK1qCCDVMG059qUOkCkW7KLh5gG5E
6wXC+fr8VeK2p/EeR4sGFpONwe9KXtc1G1yIB7UOlCPJ4njISnWL0bHZ9PB0
QR7LrfLxgkoGeZK9HGp7tz/8/0aBUFdgnZaTb+f1reZnzNo0zU3yrDeClU4u
dJSarntzixQ/rzqYOXLxYy0YRlny05WmEdVaeIV+Py9RJSBzoDVzfk/Uz4rx
4tnjNIbGqurB0WgGa5qVVZwLNywNaCDnuI4P+tAgL4GU0KfDzsCq5DxJtbq4
X77eE9XWWIm4cSMAmGIQ3L1Bv7NprXKzks5J5WQiLZ2pqHbumgwBT+QY8IxK
aL9Gv1R5MPtRRAaCtcV+U4LECWx7We65eNHhNpqTCtSIFlXg8TkPhSOTpqWy
i9zBPTHlKNQSWkOXhHa/CovVz44SY8b3a1WG9aWJ1XjMXmRDNvBpTMJygDd1
UN9GkhGEWf+0ScgQTsxK3RyPElOKqcDdcC/lDguA1kOnnQXBrphELe6nXFee
0tJzp4BwHV8ygpYOc9ydBcVZSmcQ82COm+rfL3FXtmJ2BsvLeXykdOfw85yp
IOasREGRYxTrhVNgGUaDJpwNjp9cLYuBZFUvuslPRqovewAEk3FF6WC6JNX5
ERJN/vLNeEBLXR5acdAj9pGS3Lpztt6Zki4Vip9jHYL3ynIAYsRdnaSorR5V
Zt9mV0M2H9IA9Uatq8hnQKWfepkhn2QrPfRdSR7nuoByzvPj7clta1NRIhpQ
67NQcJ61oONHKYnw61a6EqJ4Eo9+jLSpGP36YShiIXcCcy4uVrXTUJaUCbTT
JSeauRtYtrJWjmSJsVepMzzB8NfEFeTvDYP2yld8ZdyBBAJy4CxJbtyaS3nK
CkP1eubHTTrKX0T2de8AgoVFBLwouYUay9KX5/r6MhnvgtcoJ1y0g35N/Z9m
mUWlZrPTq6lBh3NC+ghuClrwGWIs5+4ZZlmJZyJEGsWa2tiJQL90TXFF59YU
CnyXfWL40DjyJwktxVmCO7FDx6o12jbplmOGDHcgCUnmHIcByTvbUVtxb6Xm
7H/WRR+9xp11a90YDx0RiTNSc2e9mb7ChNxLmCpW1h8xGtVR3S+rQ6MvpB85
sqPTgYkCuKSlRhasR3orY/q4K2zmiH7SfOWfihuaH8drzhaCrscTfyzncnen
Mc/cBmmbVUCXzMPc94khpouU5HtG7ry/ipoW/EQez8gPfkLbxb9tgsROe0eB
oK4kvzx7pOeVCgv9gbqOkdm00JoEYf+U2nJFd5Fs6ccBsXE48PtLdK2b79zC
LPMaiFwzUtDbfut1ttpu9bK0drZJ/DUfUpL0Ff/3puaZULagxMJSB19its3V
KJZHS5QiAOHThC+ojWCzGbHXsODmBZyBkC8AFdzNcUy0yXSCz+eDLtXRdsw1
xhNMYtdzwLMMVw8xbnlyhqpea5Gh4flK1Jpz2vpxiAcuypKnSS4gPrOkBhNq
vV83Jn3ma8ul9/hNI3m75JHRzQIdJTTp0kAqiSCszBxMKH5lg6t+1XOj9Vpo
hqpGltrESAzYxnmnrvNF9Krv9cfAeMnSQuaOtVTX9iG4BEbNND9gUSF1abmp
sziPHW1cyGAOfQHmdfiKbuH953zv4Npi5IMBOjjxqVOyhUndX7NijWTVhcCG
3KSckgbMIT2N0XYfZOcZE1REmKe8lJdQ8BiEghl2V2pQfEmmEzb6cryEdvUg
c3aJvm90/qR3ONEzT9xekFbR0Gs9A1kSyfezHIyCQU5TQg4G6VTB1ierme9+
ubMF6umO7/HAgFu62yCLcc49DfXZc2MhgEwENAykatPnCjHsO21w75FZ0RV8
LumLmGTSsgVMscLRLSbtbl0tvZHBhy10l/1p35xhV+iTWuWH9T/vP4+RKxUY
gX3nt3qA1f51NW7Yyw5RYkp8szYUUQr4ztviApwLdMI0sMt+LayPxsOWJZ7R
nGdkuXaBpG1gn0V9P2R5r02JxSxvJL4uRkcVbJZSGuQK1VfW9kzQqCFcsO2O
5N3CSUpGrSVa8OBo7Uq+uwH2oDIldgz1tVRHccYns6cFOBKL9drxPKoCDuUV
QX5OjENGbTo82irinAdb6MEncKa48/PWFm4u3tbxWqpbLBqEPFjRg+N2NqnB
vnj85PM+Ta3AkfejbW+KZmwXtHOyvhzW5aspWjbuw2o+NHIKlHYfTJotkUJ7
1r9HEBY3GJio5IzScNuW9MCAZuF78Hxp07j6UcYz/N9dR0tyMJae6tZATAMy
G23QkzgVK7gbCKsn/MIn58VREbypFpowd5P1bV+lGTiOvFrpdukE8ZY3MW2U
G+hTGYrLmsuW0wIBrErich2zElgUDeKvooQxAxmdmX57xWrc4FLCB/k38fyk
8+slsxdQa7ZynTopBKtBUxC45bhSAQKxVCKm6RUXuewnPIQmEltjM46TXC8u
89FXckJCQ8fmWx+HNDExmSt2qfPrjHzb7/hm61o74tNPYObKyh5uo0k80jRY
30tqkZ4TgOh+VG/lf2cTNvZ8tawQ02+Xy8mBr7CvVQCF731Gw/rmD6sQIaNR
AlMPs9jn50CPRubINFwWVCZ1rn1PLzyk4pzrDxUusARqsvWMCOktO4gtj6+G
XcIFhDJ3RoXgnSnhcvXAviagHpUkF2uaevVRWL2b+ndCP70x86YubmAbmQb/
0yVFBIDn5ie8/o/2ztxe1xo6dSl1DtBaH+6nsWqX0U5nSNBmhBU1O7A8i0F+
dVy/Qbx2i3RDVsenLo1sRav+VvY5CuJoLSFOxZnNsajhfNGhognoDckhEU/U
PSfoZM2KSdKSOI2GXeeAyakO4S2pW/JGrgWmsO+qBWhsA6tCMg3zPiYndNxi
fdnOHCU0WhvQwRdt2V0yixAaAKQYjmrpYm/ZWerDhDg9TxJ600kFAt13LNgF
0Gk04PMXsjStoKczSTtwHINdbSLZm7Dkk/38q6iBy8hqYFeiXCY2DLhoW4S+
ca5D+0I3vzrELO5J/Y6AMNMarXtG7sdEsIqxzITwwzxdH8KyYOcPBeq+4geL
JxP5R3y9C72ONStFayjFX6KR9e/MYYi6m3ZC34eOZav6toJHEJprNq5j9wm2
NyIFxuz6FlpTqSl1k1a6f6vZ6PG4m1J2OExOKub2wKHJ/UdL1TrPJKipmRqb
/nCwBzZK4JRotchKApiHb/X7FhnvKGZy4/OOuWO1v15pAimUlOGLJNsZHm0n
L8RsAJw4dc1bddpCX3T9n7xGfnldxds1bJsUXcr5fFVwE4Dx6zQi02imTYPr
TBBq2UGKls+3IorocSfTkGiDMXXkQXfTx/YZJhM3Z8NSqtHdPY+QonOu3tYX
VT4bbSNmg4ZW8ycjh6LL7mITTTCx3jtMxzl6iv/w0DTQu60nOh/GDxMW0iiF
s61L6aucYjxTM+Uk0HCTE4fcpgturS1SsO/OpP7LEudUlkhFpZRSCrNxnbuA
72MzSgjwzFlyyuV6dNLuUBngXTpDWdrDJ4R8ICElIRu5O+vv3q4pgKSWFV3y
bJAxHeSG3FBbhXtdB5IGExtlPe5y5whaWDDfsXNTpXpm8QCCnEGZ8cNZkaEh
VFXRp/mzFl+ZDE32kwNprMMf3YMgFUJGP/2dyExjLiVOxB3UJdQTRtESldHS
jYDewsXIE7kCZveivzhIPtUNAeCMyA3ntfU5wBiXDetOHY/+Kj30A37e0dI+
jiEIPhUuqnqS7WZLXwl+JVKEy/vBImk7b0Cwj4vg3Wms6aMl///XbLBtv5e4
qXcsQgDzaaU/xqTFTNdKHVKC8YJ1o/74E6KMBqBVG4hMPjhEWK/QrwrVi8GI
dM8FzQ5SRFXTEJ2QMw6Liw35YWJCswccMxxBJMuHtwXWsD34j4hw+B2dueQK
g94Eo7YnId8ODcNJD8VGiOV/IgnEk4+RVjRPHEbfRTZtBGLUNe+ZRCG9F2bt
8rEXezhsB76QAtkbifZGtqttiirIW6qtF1pgZR/+dD9/7c6ESJntJZsf6U3L
0bQs9bRYll8tFfKaniY7q7/tebzY5UwSL6zrnRX9IwUmOFhTvlPkRm4DIJEv
1LSNQhj6SSDSXDUu5IUhDnH3BPIcxs6BsW8EtzhKYDha3zvJ8O4lty7dzb06
dfFz+jth/2tfVP9ZZqidiU3oFiTL5+SFK2GrqWRsJelsMphT7Ikdl1s/Kq3e
HUD1O8OXSLcfjsP/PJFSA/Eb34p1kb+ZSRpn/8kdwnFZ2yHtIrYEt9alPFYo
nHyMSZ/URJDtNPWAbUqMJ+F8mW8/Nts3dqSNLn+aIB3FjIAg9ls4XE7EF3/c
gsuV+pidbmpRjdw7jjl4VQbw02exwgeXu3wkPNDiNRFJBwI/00h/zwEaukOi
m1IV53nnQjJTFpTLft7lbVtoH7PSfq+DuN0t/BmKAWjj9nZatmyH+HED41L8
2aeKGkWCvuXlJ4/qJ8jO9Ts4neUX/k3g49UIwGeBKoKlfKox3vjR6016nYoA
0dnyRnLLfolZz66zx6+dJ1izSZDIUXBa7djN0w0CMoUXoeTow0FpxDXXFUfj
nMguV1hhlc8hrt9EzQPzGRBwnnc2ypWbr5PwNeZlWwIixanGyMG+Fc7YwusH
ld9ZHFQUH6Olq39qcezJUBzPyD7fMvOjOax7aAmAy3lPdrZPe+2l5on4Hnlt
ZZGGO9TZ+kslotlsh9AjswAfbxHhelhBVwsZIJ7ID3x+CoDKZOQlUi/EfZ1/
17U+wl1/ZgwriVSERUCh6zuWQS1DoTRjnBbOF78Ju7El/sGdocob9iYPY/Un
ivd/gECd1giDKUcMDyySjzZB8suECyFsWdBy3EhYKPPeJGDauUyEiAqEqKur
sYdO1yUs0ukZcIPbfRTTjs5gaG0VbcPaENIB23Yf/9Xa4+uqro4sRS7mhqo/
re8kYTVz7s+7DAeyeiHpfYkyN6sZdtJ7mLs+qQmWoB9c2spMzHPMp803psXf
wfwTr5/gSH+UYoCi7MqvGvmiRpeoAqowhPBn1jy+1mQcjFeK4xVmiYsbvpA0
4tMohOVEdWbQMVbWJtVSpTndt0gUH6zm/Bikgf7sG8BfcmkKFrP3MctruUOW
im0j68WhBOs038n/V63TQoajE9PeTXlZkuLyt8iDQwPh7rdkCGEBLc5HDpoJ
hh9T6KCCoVuvjNWPgyqNGsS+fw0WmzGEXLuczh7Luyduk6ssuwMYmqVs1dpZ
dYsJAcpTB98Ff1JqCyds4zGkSqYNm7AfAhtfPuGkBQL30gF64Nd8oLta2faO
BZwk6v9vCBoCmKZbCy8iCMiGxHodANkRreQ4XfOizisghdoRZvCV2HtP4hKB
MTAF3jjDMQd5lJDKDtiaZJk+r+FzQk4z3sYgc4nCHkQAGii890xOSscquIIa
T03GtIFff5vHhXz389l0SgWfnYMASpqSyRSJkd4Am94R/bDcxPUtkuSDO3UU
8CWwwbmwqEihhVDX0rDhoD8mUMMKDhkxMsXv0ubuIssz1uvsDWLKtNAt0Xwn
0kBDBq/AOrh3Zzb/f6uVyjQLjImfhdwV/HOal3WI0QdHixuJxisMKwp70VJb
N3vDQtu813ap828b9spqbjx7k7aY7/+Qi90dp7mQ9w75lejgaIES4LVclcqa
1f12fC+c6x+7EEkmtG5vYcgocQTZn3ksYp6sCfP5+XeO5eRyVzKTe9OWa4DL
It9CCjYL8l07DJ0RHSLpgirkuh6uIdCtd3d4bbJzSgorK/fdm+EMvVgVJOBY
UDy2WEEQrwaBBRqjS3+sy4WDjsmhdO0ubDACI+wfVCMFpgZiUSNeEn5rI7k5
W+ghCZmx2XoFvSsIkeXKP/TPPuIgK4NxX6NNNpEmAGCjGE3Vi1QyOZ6DSq9U
u2w04jNemfEmEWLF2IDZqNcjIkeTM1JqptQ+XW8o43yOcoA77b8EeIbGn8Jf
CI12NQdQj9m8e14ISntMW0ot3yx0jcfOU3s9eQcbDLqRY2F/g27xOpIsGmq1
euEAVbvgygNAsoBfPBD3HDikosWz5uAxeKBSV2aUByT6PIRe2YwgF/+OVLME
rQbuJkInMc+kJ6Hgw3mFARqOf131htoYFDbnirqZGzbxc/uY32cM2CQ1HqBF
PO07m9guRw5jTUKfiW0FMlap/ddvh9ZAUMzwrS7NQaJhzLPp+tHLOna3B/F4
Pzs+DMLS/4fugN7XkFE6teVfPNoHMquHx0uzxCngGgp0eAsGyX04wVGSVSkP
4iO2X8+E+r37CdxpEszMn+d0S+d6SOTBJNckbokZJKjtcGU4ACcl7oxjzi+t
ePfQAt9jkUGhvRCCQjsNAge9UM000xO9BliqQ9EKuWRReX+1RZ0i9og9cykT
21kMucJupKRQFbi9wqTYZnwiCe9/Vf6fhEQEyrg/p3leONqZjffEPlgJsnYt
Bs0Aenz6RStUuALpNaPaRjCsKlAj2iCRDKeAmafbLy+pQE+WrDmr1xB1t6Nw
LQdeBvjOAsPQ5C2kpk6phzijeoYBx8ftsK+3K+2EGYEY2expM8g76pp0tV6y
fPy0C4hvW//3fWZUD9+m8LYeR7YcRGJqB/AW11RcaqVWmjSSJTEMud+daPVp
XirhQIrEk/9C9Ke8J1PzmqzaonRcCcjdYxn2O9h/GBjmLBUKTAbM3gyHUEOF
IIT56gZK8tSnX/0jCwHjugcFOx5QOCC0FIEdTLl8r5+RsQ6/qj0gtgWsD/7c
/Vmr90k4fG2rdVfJp2HXoQdnCrU5YW+ehRI3iLgXZ30UUpQ3OnedryqLbJ52
jEIRk07LLRSlJJaFM/FGSRFDMXF0uHGUE/17ZvKZgFRLTVA0814jhxLEX8ZO
Gf32CtSUqZlzHwQK1cQbbEr9nNsYuFRRkHxUWFQ095/5HZ/hw/sQFHT0H5OS
8Zo7skwBFrCD/gSu4od1fZwNVxlPJ9uZa/DosuJ0iWZBFLrMdhurJfEPtMbx
6S+JeLBtRhV39yYFRs6qcssJYt7eQPEdV08ExYfN56URqppN5/OX8IeHX6HX
Hpyb1s1XsQxhHFl15NgKvJ7cVqC9zKLQbUO5wsfllcVGM5kB2af711n3RCvE
nHXbmSUKA3esVcrEE2uJjVLm5PtU64nqvrBnyl94ADwthICxsIOL1PqCC9Ag
Ds9yRc62uKciusp6eG6qSE4nNHibrvPkdUCfFVCUv8P0o9E8o/OqGmDBSLmi
Z/BoYWR9Ov0EOcVgzHJQhbpM8+daT1fQ49pTETQW3hTDjPz8Gls9IN+RhIk3
iFwA2vlniEYR3u0o8TAhTF+xv7A9rCv9BW1xEf3UvQ4Tm3NoqInFJQjIe7ou
U1zHNOf7GGBonObnYUjjmPSh/6wKJC6vpvY7pXK9WrnuRAFc/u/XPpo6IrEq
wCKMRKWc1mBasoYwunh8QyFppQ3s89EH0xNS6NbeV/65+XnGfR6K2luvefMU
XY2ZnR4J1pmnrRGvEynZ7c59+JMeZTd5IrSHuG1fpHVzrvbFv0rCQnvRO30T
QIJa7h6Csa1KDuy1CvaEBphopRNp7iO1z1SvjEKj3L/nMd/AK3massUzqQ4d
VfVRlcHPmP59TTY88eXvIeG5fgMcVTs1dH67QDYY8e+8bVfqthrMftntAafK
QFkkVgt+BO4ru1HgATcUnozZn+tbNabVueGjn8RlQFjq13inVa4tI6kHgtI5
3lUSV93ndce0SJ2bPe9EMPpWb9PmiRj1zujitG2kr1hMfjn7u/DZKj12maPk
XujIghTZwA7vtxx/t5v4B+JlwtQGxl0TR9dftEa/BgixqHO/ctU2pJgCa3tt
vnQpuJNtUiY3EjosaBOEsHhWaC+Z0BYxOpCwB2yktPUcHUzjqccv0jsv37yp
SAmZ4nV7aBhc7p8d5Yt2PA/kJdQFarAD6RrxiYcewOTCB9Mqfw6q13wG/YZs
tcoKrnjEDJd//fsTc5MiPUrlL+cLmwpcicWVmNVgNnm8iWZj8nER5MOg4EbH
gqCOiIte7wWqS+xJU++2nvJz8nb7jpByX+2bAsYWR4geNmY5cbj+HZdndQ6h
rkuzd86nCVefWLoqcyWFyGExWEInFO3/KVfxWGP2yK09EY3jrcSWGUuMuZ6s
izL1NzrmP1ew6k365mRRC9vNfO2P8r3Wq8mwh0bj8JgOVBGvIn8RZczA1zW2
R/nIY7ye0KrMsDhq9HHLsC4m8fGY9FEmtMR1B+n3aiWc6fmFR98o0P/gqnkW
qxCSCzP6gsn9gToc82fPJxZQB0WNgtAIyPODW+vi2Hdnr7hEnogAe58LA7n+
Utfz3BLa+kIIVMjTegDf4FnEHGP6Vn2GsMmADDAtcdxG47pIh36T/IgYXukd
rbjb06vdoU1lVoHfFAd9fkCKhJUaeLf9oqSvvv13f4nH+hj8xVeaHOZgBo1b
5D7oxB5foir9kq3c37nOz0y5tNpxOg0EWelxTir/ipC1Irvhb101hHQfXDGr
WDJuV5HYNtcNMCRaKeSR3DWU+TcBPYzfHgnHBUyCcVt+QogXNXTLDaTu3fsA
tSN2hqFJgWWMqa3YCI/oODtzk7Tm/vwte+wvHulFqxWX+oTvgXQNfqTMWZaS
bzBLVeYgbd6L2UtwE1PY4+6K5SiHJN1TsO8RNY4J4y72SXefq1ZBofEHklIc
V6Ag4VSinaNcm7Dvc2MhO5B5bznWgqrbJqhlMLNfg8g6B8jJB3VQBIpB17g8
0X7VDPUU+uvQiJ1pfamuAe4V0RuermUexuFgZzyiHyff6V3OsbYYhq66JDdU
YHZrIFBBzQ0+tOnqfk93ktwOkzIKmzOzE//AkmLcP9ofita6j4YK/tSXVcc6
aEVYVkelZZTu3v23aYNqq5nfRoTON6qrnXit03VwU1aYbyyJT47kA436XVwq
hQ3VbTVc4jV7Wp8E1UY/YvIOhhVzQvjEBNpnEUgoTkT+HIDvvcuLyXRNCEZ3
dRMaOX7Z+0Ujpt13Pscxd5W1Vh0wesjF55BkjnaY0VWGBsAc6EfAk/RNipU/
fQIoVsZ+7hEiTGd4z5U2wA0zQEOVyLHxFzLJnUErWEZZt9xyo/h4P9Pce3g+
srY+BxjApjrCGTs7PTNmxuZ7Ks7iLQs7XU4XHbPDWzwd5s+h39xUJoapoCMB
vRDgzi0a/+zwLf6WzwO46xExBzrsLm7aJUijOUmWQO+ZZbJWKeYvhM/Qd8Cr
IJDmHQqpVXZoURcAgao5XiMJvwKN7V5lP9OsXZ+KY83j3bv+n4TY8ZXdyIXh
SX67Vnw2oRQ4umGLJDCqFerWCMTjVy91i7VTCvpuGKXh5S+tvO8tvflDd+7j
fChClfW7uckxdbGGr5QjW0r00v64vOQiIATXvQexkIaew0QfSN4+PDTQF8B+
238AMynuIG0j721Qh4601uIvl87Bz/pPz1HGvFdbZva3iWXPO+W60MN8R3XY
9l2YrvRSH8KolxpCuTTmAPer7wWu/r08irRId7WavtdPMgOn2+16BvLdCNFI
3VJLazNonoeKSVIcSxhjWSpHYEknAQip7mjAOYvhrVsnlG+FXROuJvp51Aes
Dfk4lAfzliZ8QXA6y5bBEXeJC0h+OdzywfCIYmww43/jUZqDQLjA8/4uGIj2
5YA49VkxjAmmNPTgVrg8xhg1jcheyrMB4g0DV9+q3qZEmfM5LYu3fCUcjz/P
Xd0J0ziiH8AJGVCWSNe3ArZbKrsxIFY3Br9GzL+9hZ8UlxSvTgmkViFvrQvn
dvePG2tC/bUQFU6KvJCA873ubYZIPeCBPce1jEW58zwZZtMr5J5E1+zTNRBB
0TuONGHfXAnpV5sxZMUCDjLDUtY+nxFqRKIs6bCm7GDWF91jU9avxHrQtnZj
vO1f10ZhrbzW90JdOg3o/R/FMji2YwTtDIuxGRtpkXZ7BsHPf73uSjH2Fccx
2hlBDoThIAHNvl9rARaVH0R3D85zRY1chg88uXg6WEHDpejyEDTXi4GixiYk
Dt1ysFp1icRzcbKERCaB6vsqSe6WImswO5owCpixDFc6gHF5Dof7q9lOcZLT
gyFPK58VOtCYg8+0MjzIIZ8gwpTxGcK0tQ5B8kpuWzVzXCHsRKCUGgPgiM13
Yjwk5EFUHujltJbnyO6XqMNkh5DjTg4yOvmIuzMf+j6Quiwi8G1z+LS70CnR
CAOpbzb9sldwfzgf9kS6N/ShOUht5zNOlBVKQmCD7N3OhSskWo834Ipev56q
9CfQu+pJtIfBIFVX45DjiHxuY1bAGct2/dlSCjGAljClDab3H0beuzUro4RR
wFbkaCdiDpqdRkROTJgzK728mWmR4TSgaovo2ARzcWZgfV6APAw/KBR4bkie
PQgMmhy+jxvaStcgoLaamFYzBQb5ErFSvx1KEIaqSLs8H1jeQujHERvPzobX
O9FocSADO8gqD2RtsueCM+5PiTSnjoyKtRsOXtpeMT3hvLGwb7OZzdfKlCPF
NZGv7HWD5qvXR/uzQsWx4Kj06PJN6l3S7El1KNxVP6kQ8AFBbz96FyVhtsZi
Ggg/ZjJNrsnTCqUa2aDac9ep8UCaRtxcLs+/7N66qJzIRrxetiwteAzMiBsg
KeVIokngiaXXsaL4FOOfKROAZ/uLPcNRoRtTfs9KkvZM5rL09SwwKvWlQUSh
jhpeyvz/MjsGzTvKCD5xaG6Da1RIjG+1c+HKa66/OetP1FT1VU3/FCJCQzY2
d7v2yv7EK9DKId51MxNWKxEdo5HBG2ks7mTPAEVX+0pa7o1A2o+OdQxD7keb
IH/mUDFGDChZzJao++3p0DJaYw8FO70gZun+5hP89ju0V11KUNUU4K0mvFn4
9FJHxXrf62DVEyT2IzYe1Ys3xZnz7k/Jc+LX9C0483pdesOwj1XrewupNhzQ
BQv+GvI3/CQ7FUlKUTzWFu4gvn8jBDCBS6rmj3NGvKy6xm3aQ4kQpcXO7W9T
1/LUTXLHpcH6rBSjza66IW7q1wrUTUp8TiM49y9NLhivCrw5g4+J5augBJnD
Zt3eJ6H4+zHi72OirQKmrz/Lpy2R4AOqRnMfGmUu2DwrYYoKkdTzUIGr/f5o
FdmCucKwx4vlM2FrlFG9bjAT7k16lfqPYmORb9vUb3g7mX+K688btvU/kq6U
FV5XwIvrIHe9QaLAZcg52vzpUwxMxcVJsugqXsqnuGB6IITmuKGDGFcjbH2S
177tW2MR4GtQlHRc/KJ28eYfPbIpLhzJX+AsqTgznJrBq47AbUuctehuzj8S
o3WJ/HtLtaNpOA6JnIMmx5EG5ilOFSZYFiBZiVAgTJm81bQRwf9zxDH+g1H4
K035QDTqteAulvIkY3Il1aw6DCuKa5DV0v1yA9XSNjBvX9Ow0HVHagKFTvWp
LqDqb64hywq+jYsIu5snj8usv31S/laUglw4V9MTzE2uLTn3IaZoUj+GzPwy
1lROtL+m/mdfDC4JHTg0Brl/JxawU5DGZwsJ5F0sBRw7cSEzgv+q644/1x5P
9qF4fSBs2nTkOTPbobu6UWYMxXV9jMugSfJ0y2Vyy3mXQNcA1Y09vIJSDMvd
9vQmuNZGmK85RtsCAtvIgNHQ+jEghRave4w/19YRPSSfyI9DEt4HDRC+3JVs
I1kLKRwgh9DO2194kjrTwnhF09fHXn/u1E5xnXZViy1LYdbOOINjRWk4evkb
+i5f6mHYZCNEH4iI4o+fEE31+piFK35xbsvIlMbjyVu5ueKqUiFgJlnT2ztF
YbKtl89qMQkjI5fRXR24oNuNOGRZQnpg6ML+o8k4/uuSSzrsonTSv7r63rws
dcR/GGlL4Sd4BZE07cUo7DwAtQfoVPWT+gIe5vnibkVPuRD+KpSNGnxc4NKV
VtdFZUgH0dwnrlD+ZZoGafksA6UByP1dB6q0Sy/SbDt1rNkQLqqf537ycUYt
cY9w9OhQ2oRMTKwaU1QesV6xKcg2SAFSHEaKmYIBWawkrQ210g6SgeTmQ3WS
8VhPikbMfhVVtOApiAnu1OakGSWoed6+2LGLtrlFyPGE9edtwFFoF3fXzC3n
T99h6mHnIb0XQ+tBbqXC0u+z4MOvX+8N3w0IUywMD8Z9NkKzLva4TJys/gmD
elj0GhQsbTItzGDg5q7qw1mOi61E/dGZ0YsRC/4+H/l/Sj+IEs705JSnvCnS
9rovggPGd4Vpb5h3dqWjHaj3P2zdxk1r8ubHsnuEh070+xcBY6H7iEBVMBfm
a1dO5p0SGodUY2swmJB1PJX4TF2pWPWAr6N1I+wd0xk+Hs97H5ih/ZFqSY8o
njbwA0DWM3o+YlxCFPwd18Lfwz2rG7SDrm4fgdKcpsEp/3v2kMOXuLg6QJQG
rWzSRHL3lSbLOLM0By0OuqfxfCX1Fs8kMeFikE2qlAp/veZXbibFlSjUYOx3
MpA3GHwQdr67r8qHmd1SuFLFtu284NCvF3Fi6i7r8OchmSUJBiLvk5GDy6cJ
Q7Y2zyHwf41xDJvb9YNzIbFWFOgax1tYI3eMXZseb9HV1E/9G0uMupEKEohH
Uh81OJPoMDDVdIHzhIjyQ6ySLEM0XAVXH3qCgW1f1OXw8cNzFzgPLqWgFy9o
Eu92TODAeLOQf66NFIgef0o1K2lRyqGAOlb1imVFaeYVpYurhaKCackzw4FS
SPx/79Qivz4/9csBnirBxbJ3hkusPS5F6Hfm4ldKwpPIPGMEdqV0ACZvRGmy
n+/PSBNpaVA6u+NcXQOAX+41IrqmBRZkXbmAFebooTsam9veg6tQHQrMKcSE
Whu4sFytsU4ztlWs0ugbENDDHtHhrD6nMVGx3C94MmiT70FsgMhbOqOCAoJ3
RtD3dL9iSTMoOOpEQmw+Qepj355XqH8Wo/EHGokVbyJV863mK1kVjzxsGcxy
x8DhH3I7Amr2CTmtt9s0/CuvHzwBrY27psv5ZZAy9Ne0QWgfGw/7rykNnrjw
I/Xlk7REotNooj5yH2L7DGM8QKsesC7y23nCycr8VUENkhD8vfDjw0rkjUZg
XtT0EsycDb6IiF/v0L8Fqk9tzM6VbhfA3U5DKK8FfqKKmkkQ156M2vezqVwp
UKdQHRk7stJ3MaAQj1FVdNvirR31WqMqpDs1xUfeiWGU/4G+OzEKToAYOlIM
vOutsAc6o8RIWzQwx3biS4EGcHTelyEA8sK7JWoNgZSjsPeNUQqoIJ+IC59V
hcCTw+IAoHQVNz2YGaYhJ8MJwuoUyRdoGZDeii8q1GX9SCqiniksVRChMk9O
bJwn0YjkAmH+RjOzX4e05KF4eyOxmBeVltgtvqBn2/5FckSWfRAdl/qFc10A
wdPRpvEyLe4f+SlBf7Gsz2PCbnxWUvDaNr1laQy8TnMU5SFpY1PEOsHLVbAf
4r8boaDqZ1IDiXiqpVBeB8DvAelMJrQc+WfbtLIon95U1pXit2FM3UpC2Pko
K2F5RBzFT6xq86GinKtoz7O7Sq8+UeJQuhc4yOqxeFfYzbdKwr+HKADLJIWZ
o5sWFRad03aNAWExuY4ODWPaDactUh1amPMs2UQoxKFa3NII6Eb2iSy1KDvW
zze1oKS6yyprSbxnikcvtlc7FC+qo3r8RIvyE1jRCc8oozFx7nxyxGOxlXba
sKQYnu8HQ2tWxJFCQeZO6XX7zNP6nwmj1GNvZfRW3V3Ig/P/C+DmlJPNR410
Eg2/SvO5trqxYRoQ8AceXZ/a+uxrxP6D7ZQvR0+5HWluSL2CjXEUos3stcqY
MpCRuWRm1JIcHXqlUVrPWp0XodF3vyCTcwn1DVsDxxdTaRFHi8JoQDn/iAz0
oKz8PbUqaJD1XAM7ORSS0b+wE0Yr4Rk+B2YHoaXCQPmZhfzVPGpDu9zL+Pm6
ZOTvK8bQKDUrzT7D2i1WWKtcmBE9xm6kv8oIsNqusyi5EXgvTDv53QFuY7Sy
p/A0t0gyh49d4/rJUllItQfpE+TPCgHjf9JiX2ZwO8yvPDLEDUhL3oKe+Hrk
ZDJ2KTWL3R/7gzW2MwqzgwM06Hp8Vvwckms2Hak99g6Y8pvfo72cQaikXo+6
Lt8cqXu0k8g1D2akxwIxnkt0xX7Yhp4UENWL9L9ILTXIjytXEdft34CoIvxL
IyXqBhjQOuULcOZFa7SzCSG2I6gZtWhe4X4L1Qn7JIpKdSy9KdCum8CqQsDi
ay4vqAU1LAbm2xYycmvjqF2g+AAYg2CDLHuCvuPIMarlxiOym5JTKVay1qLL
RBsseRsBhAnlIFATFe6xjHs9qqMMeBgiEjXQiClCZnCwI7tlZH3wV1g9JQIF
nb4o9Tc40WZiprgptqj1qm7XotV4IjF51IRmc0xtqCr2H0Ksze8iQ7mswF35
BeVB741CUr9kekc3J9s716uNL2tgn1y+Ao8n9fUkNqL/GIEx7k+axpDxlgRU
2KbkIebkmbHY6hLCjRC5e5vPYKWvuI60+3a8xHDDo4bqPU1RMW9ZuUZWFUD9
i6KBYrReR+zlYwvrVjecNp321Qohx0EI/OZM08/BjnqFEnD0VqrOqPZvMqkb
DFA/Duzm/RfHssbbCGhre/h7ncIZB0FclwFrJQnwF0yDErSb/ueQLTo3GVpL
ohDK0KiAo9kxxQdmVfPoByRPpZoU5UDdPMZXqOmZZovp6772kmJfzP1Yckue
dLUZ06VthjIiy09EfDgnZQxmC43K8XcqY6LYMnRnkqNUru1QEWtCAQpfGBbb
EbFuVHfN4EHl502nhuR1P5dy8vUPfS4Th0jodWYoEoDBYrsKJxRjRsvFEzcM
kK6K0oqDi+m0n8uqKQoSbl8BKvzkXFGCg1NzmV97ZzE+T1leGuViU0OBLYHg
c/wNYY/x9TnCwtzxKDRrRFd8tAdGr8I3CKefrSVP56H1qWR4en84DI2BGJ8Q
HmOeofXWeZGlaClhBsK8T5rx1L4aX4Dc679wetBOHQnmEywEjykTg7bn8ayY
tBEjA7c9Vo/mOpC7OjoREXzTx5IkXg/MAGW+qr1x//NV0Adu8+/D5evKR8j8
bpYk2nNdGaJxJ9zZHGeLG1NDP/1b8+aMXfwRQT2sXISA3PPanOJUJM9XdGfn
h19KaSjAGK3/UrgWGf1vM9rMnA3E1sa0tfRt77EN+UR4dU0of8sGg3Tc5euJ
d70Nu/CLNjMOI2Ag0x6+vU1/W2WT3JETrX3V+Rrm+EikWD03cggHfhqtOcIC
Uf3U7ZM6umB8AHPE/Msl4DfwT3wH7PfTtDJu2AcsCamaRaF2w7Y3yNHrIWMj
YoLqRVFhzv77wwJA8iKR89bcJJgut+rVdDsw8aCN/pIYWLs/dFrODnTSe6Oy
fP4dvWbybiUzEJW+GZ3yIbbYjb4gB+C7WJR57fDgOP5P8AtkleWX4UIxbtOi
EzUeDlAfH+UV4SjeYUkmrNMt8Ebjt9H43nd9ED7VnUDUG/bzJZG0DTSk/I72
yCTsydHhQr8hKj5A8TvulUcvpydefvXBBHXfJxIrBFoQPa9WewBogdgXkfLY
5+xys7KNKkpSNGjFABoHcSjAXpFfY4nHsl9AtQaGrdeDX5sXdwommNweuVyj
dPYaOQoznaUyMK9IN0sY+Zt7eKfr0szsNK58RHSghz96tmAYhysEKcZNmUhz
x/3oUyDLtXju2Q0NLE7f2CxHVtOyBLdmWR1yYvjjJMn4TyixSeREoRuYvBPn
Gc3BuH6G+RA1aMjFtCQvpCVoYBSX9U9MNP0G/wn9zL6BJk22oGEqcqd4wt1T
JcePekaocnVEcbIKBg1RhW6PqU8prMi+hmvOk7dBoNsMmd1wJjZmfY5U/X6y
o2YG8ueNX/aMfzOmaQxzBImqDNmNFxBwCnR0eHfdIhnw/Iu92SipS+96xL3I
ItjHpVtWcL50YVVOx/3YyEHfpjees4j38feIixqfg3eLWxje2ap6vhQ9IgPx
tG8WfvjHgDj2Vs5jOh8pkxvJlWg+2XagOVFpgDSPCUOiX0NnENE/xkWPGIji
gUwvMToHQ/Sq0TLGdDkV1izEalDz1d6cNKvpY06AQlkw7dRWDHnQWyGrobzE
eYtoTzfbyiWLoYIVKV+y2dr9gGAqVqi8k9u+Of/I9KhsEi/LPgCKihTY0yck
DYN/uWSb5W5Zu7eZ2tvw6+iYcul5st/rmROCUoOfrXDKsa24/n/Fb67t0KZm
xJLFHvqxMkJVsCxiPlPg7FBAsTr001KTp2m0lht5weDmInsGFUvXPFBK3Pdf
BDdfVJuP+3fAeCP/JaqsGmR0ihWzRIrux192lP214v8hr0PrNHplbGXWxffT
CQlj5SC92ESHvue6oHhqlRl/3SD2NkWnKEQwDL+bJLPnZL87uhnOW9ekLXYl
cCm971I3b5lIzHz6uKxccu+TnIpisb35yVX9873qddL44CB0oe4Xor+YAVVW
e/qX0I1oyQbUEb3Q2gmce/N65W6BTJDgJnEeX6xz1Ue0IP17ifC+1Q5GeQmg
tdkxMQRMheBpxm00ft+6jgcLrhLT1fKc4eZ2JP/oweoWoIOyHvon2GHZGgYr
IYHDaM8ofSS+k8RzKK8S+jGgdr3yTZQL2N/VwUTv0NCv6z2Am7AgxLJfXo5j
N7gJjPEwJJR1dFchNwQwPKved2Elsdbu2u2gk8qr7Jvwx+Kr56eWgdsUAmgG
nsRwNMwb6JMg7fgo0etCC7EP9+YtKjxang3ADJiNpb0MzRFqwKit40VnFA93
jKJk1Qg6L6Ba8aFde8BDsznD0vJvto4byHpwHv4unhs2QQE8OsAZojCtkh9G
2wsbLETx1+Kp2FWRH7/OdguTD962HQYsZhZBk1SGF+n0KrfLbsE4EVifefwf
uls4tjNypPJXzZB9+qEdU5Pz/alX/BDS9h0JpAgBdRPH/IVR1ld2kiWqa1EP
/Y0gplE6mfC9gFnufZ2J8mLHkV/qxn6zAA4vcPZaW3FCU4eMMNlZufGCSUxU
XP5BRkDm3k/M7vwzxNOylmuzXxV5jDe9wd2iv7u0rh0cpTI7vhOUcXEzoU/t
w/ArUyuz51KWz27hQIBe22UkBJmn94evokSQds82+sjIfYSr8qTodTYI93J7
UpgVi1UBrppj6f3wvKITYavPmUc5QydoVmBmQtj1BN0FgkILyZa04q+dqwuT
caxhNuvNQtyjQJ+D6mk+k3KtLbwlFkWixNWzJbojRbqeAtXRBQs5bXGg97SR
OufnPf62PvCWH8BADDpUMqKhQkn8HHqIoaDKjoNfxPL150op6/QABI/x9RUF
zG7yx5ktq9FWkM0iIdtBYjoWyp1WeUoSNyAsb8DyPjCcK9QKChnUoc+5894v
pvJhStONEhCwx3vhrOpJb9X/0Q/njeF7ps5c2rI7h8bIb/LbKQkV1V3U5vuz
e/4vOELfDpndsum4I9FSF02HFkRV4TZjLETBIFnJGpjSjUxoHniRE+RR/IxB
PcEpq8xCx7IEVqWw6U+sCh7X2h8V9VdPr+WTT7k0YXjkoKpDRiZZBmET3ya5
55LeRaLWemZ9wZsm2/bB6dOxY2lL1OJIhCglfpOSJUIVEpxFOkhT4a7ldaXz
+m3O4SRjakSV1KBwm27rhDv+o1dFTU4+0jngEIDyEX7zVZZMJ1pQ6iYnKxrD
ku8SotT6ck3iM0jnl34NauSpYs7woF3UQ18CRfA/bv+tSQ8oHzRvMmwwYFpf
WtK8DTNPdAM+xVV684qOFFtkkqcKSh9cksOUqKMFRKgAPR7moWityIz7t9zU
PaQBLbXhBpKzedmqGmtpTl3Jj5ogYPp5r7cvl8pspJsKv+FrtXHdbT/73Ok5
USOaakFpB57TrFnXNfGVzjkvkapsoWwxAHTFTy7BaLEfVyQY+48509p7wnB3
AwMy/FbodHGebn7odVhx0DT1nQqJKCuhEe3/MNdwnrDe1B6OiAlF5XkW9fEg
ldq0Cp7zVvHstB8AhfRaFdck1pfv+HgveghmwbhWqWmmyyF/fdL/BAHB5pHV
WMqqoWTJg+NQnm/6CEfvtWj8XOkoBsQWgnmLa8fXgrcVesU8mQ1lp0t6UW30
N0Da4ykscoHGHbej3r1ema9BoLmWn2QfV57Kue9w5rrYCjvXHSGwn09G6rTy
xxqmwFRFC1HkmCk5FyhP6IpF66ug8N4/4esozhe7IpGfQPQ5vihtrvjDWwXs
+VhRTB/PFaRepUlUkI5/H7xgmPsx06SQBQeFo2Hk8h8cYqtMJLQm31eDjjZr
CtJoCBvGTMRZnFP6MoiRfv3zua9lQWBuNlJCnP3xOqOzslCOrOOy5zaw/WVn
AwXpgkfWHxCtUXbK+S7fnFVl98sObWnsncJBXIo3cHhHFLllFFu57hrGbfVH
mG/8angTq23OI6DWNkA238CI56eGCWN5zMDWNqIoI3JntDpy8Ip+ldnUhFC7
wsJNW8CidArXthw6vaoY4P5ym/gjG2wbYoOhAZGDdJ4/qCdC0DPB4yP72Wqy
5iHf9saG3j2PxT4TDrGq7YlQuArzN/YxGUEd9CB9vVHC9AYIMccqbN1QLmYL
9a7JbWEk2Qlgpyb3EeXXVo54rT/gfl64L6e0Y5VgkjmzR2FannsYXS0iZUti
jTUTXTC30CLjN2TCvQob7X8fkV+IrAgcQOn+KUtCfRPM+Ab842FjKqYD17Fz
JHBiGx7SUCCkemfl2UI7rPFc/7V/78EXMbv3zBttgt/zkqP/9zl5nii44163
qvVTtAOUM+PYRY/gKBiZ3TBUvFidUOsmV/aGUOI7jMoIWNdjyizPcDaN5R6X
qY+EAXxiJTuP7nGXc5AdPhhrbAuOLVkhiLWROLyFCpRbCiS1nKD2ye/dvxHS
y/eMlaFjAobtzLlZpmSnDjZ/kCEpOFuJMvl5YNXsdiS9SlOm4AXEDzi6AoSI
Ny1V+9e71/RAeNKYHYvDchPr3fSGz9pLBr1ClmW7hm0RV0bWeNE3ZpKqb6Lp
llIULio1OdOFzbVZJoMSOFGLOlgvxi20Jh2bS6QOsYWg1fAKIn2pqDXgIBRG
JV7e60/fXZyGCdR1UTKmkYEYGwFuTuj4pxNIz4NrHKdCvEhhOSbNMRfr7rr4
LsqGUC2eZZFK6Orew+WFEz+q0S+orjA4Nj8wfl5UesEtGXU8IZw4/Bc7uknl
Km/lkDAsy4xHeRwzdcctBszABw0N5Hh3SvlIKJh6Yv85s4DnbpuYn7bc/nn0
VYh5sNjN+KjcsntBISXYOVypHIlk/ZtMoGTkV2umpcxZLv5c1I8qNbLqK5nE
XOx7XTuZ2uU76kOVslkDNBDkeGTjVlEJnVYIWf8Xi0PxkzUjCHk0bD00dW++
OdaIplvQVLMuPtxD/rHoJyreBOsjIxFlwjSy1hZTWWKamgAlIW2KzMvFr6Wp
+3O+c3gfYr+uxp6u0qe/TdS5W4PnLWWJ249JcaeLLCoPv7YiAPdao/Nxul+4
3pLFUplnaMReyKLpdywJDPN/qHEvx4SPu+xquFeTjXWDcbTjk2UirnyaLj2C
iJMUG7t8vHdnkCMO7nhoG+FLr/gtYxRGRlfYZbz1QAf3/SnXn7L0HO5fNH22
xAJvNfWLAtDdurCTbnBc2nqcza6HIAbS6xfHccCE6EDg2x+NYqv/19Ptm/l4
jsfG/dxsorkH1qlren4vsobV7QpIoCij7pdUI2rpQyaUvjyBj4fhxpb4Xtfu
uvjhri0s04RhnKyV80UrziVDOL3YbUhaBJSAZziq8sknxmehsxsVc6DqclpG
Tw21aKLp55UxqDQZRgfACHfT+G8d/XdbfTsJhUdXkwxOxCWeAoRUmmvtn6Ju
cS4NUtk6qsRFF8SKLJ1umS2Vjd4GDojlEKOkcYUTXGR3lylebZGK6/f8ge7i
j504YX6b4yRtEUM9Gx6mvvdaaTjfds2FIn1jc/OLOGb3rC4uRpCOX3lgmTk1
FBWNsFUPS+y9mByqP0Tmby7LxBOJm7MaYZFiYzg9YFgk89lknYc9Yqas9yl7
emOrY4ORNNn/h4dYKXEj3frlSO8HefTGkWyY4soCXThG6CPnMxdixA5Qgbuf
UamN224xFYWrREI0ASkYOxqwS+fu4PK9ab8TmajMvj5217/88qXWeK88QSpO
loeOJOTHssaGKD/qMFtfT+tfyvfjaov1FLXlI8dmkHw92SzLNk8+ToVRviMF
VHCcYcHMaHn/XXmAPJkYEiE4YYA4j/LtjijAekgnIHC1QY1SfQbdCAsp55K2
kBxSI/D6LCEJ1KbjPEJ0b0z4KLxSC1okstmnnK6oG4YAzki1wkiGPu3A0/t0
ZhLFDkmPjY1qWP//gfzJhdUQHVa0Fe4Xakk9N/+3JPLTQDxXx2YjKODRbkYk
BXJUW+j/hW3jhkZHgs2roKMnwTVTwW3YJOEBKsLxx7iYggyahhWoCdIO0IGi
X8gQ5LuAPzhGu7OtRzCEb9yxdTF4TFqWScRlIk72eUQbBMx2+csnC4P4KAmQ
Rg0zTSouCabgRt7ShZT9n4HmDR7JLc0qtjBuZTxg8iG0hhpWhtA4mPLAwAa5
naPSlopDJ95nB6mNZ0LP0y4aUZ2dl1DYuVImUnkuv7ukSyY5i9HqsFcO8fCr
BDqrh0xbvFMinPVLIN3GwEiY0s6ygJKJydxNLPV8HaeUeAjOLOCkb8qQh42l
3CdFv4dydoftRQk7/v+w2i9M40F5PqYEn6C9h6+8pMKA+rBIJwZ7iqZOf12m
gysXWIdJgx82M28xunsE6WSLop0tvQkD1NcH4G2IUGTM6vqcZ392wGNTekyI
Ggam5aa8is4dqLYHO2e+YnCEH7PruqkIoJuotBQNA4GhkfFpkzj4rWYu7Sae
1YWNhuLT16UFweRgR+pJkZIoh293iWNSQ+oSElAKUIUu/D2yin6oi9hThk2N
jEKPVcAgaHEkrMGMcWeafVWMjWSRjj0jB2Y5PW3gSpUgW8eGUo9IGhCywhZ3
/ICNUKT+BqoNeB7ESy7jAy8/oDkO/16UnxZywqGyY3PVS24YTzcX9O/lysjh
XQ6ff/ZWs/0c0FknEoMMSSCLciuumlP3hgUDCC5VSTmesJKNq3JJW+nTz3jQ
TNsHDY94Lm6lCASVUUmus08u4V4nDX32rBB8BflFlXVB+fQ2QN5KDJ2Lsc6w
CeOsKB9eMDhxmzGMvkWaYT5kqmDyQdJiH+lwdSMn5mrTYdUrCyUMIImwWNHg
xX70rG0L8smtTh26pIHWwlxA4FQ1qyc6P+t7lsk4euUWZxe+Z31pHhxQTQs4
yyGWfUPTXmYsYHIrtRCSgPUrE6LCLWHJ2CW1eigvatQXaL/fhTDqwDGq1V5p
nzZWKZJ/mHHKQWkWrl9876ELmvG0qEjllqyiWvwOIlYa7qVUIcddKcmNvD5Z
UlMguZaaVQFOqhFlF9kHjWMKkNBCmnTP3qtiKkSMTpr6ULjcjugiSAo6sS0/
7EwxhEehwNnVM54ixZQpihee5vO0HJBDgaLjheC/haSsw8wdBTmzee0/I8Kg
1zm1iFAU60q5M5Ejhby43EXhD07g7CRmaMNngAwwvnSATmvxxDii+kbv3M9k
MMPoKxilhcXmyHRTxCvjZkpgSZrAQpGuP9wbHl9JW6MLg4GdahRXUcZN3/yK
/BHETC8X7cEqt+QDr5cVxiRp0eCDnDAUGBl/7nzACLm5YbJZ7LU5XMHhv5NS
IpjrcEFWSwL/izk2Pui0JsPs+5TNJWD379KQkK1k6FWk19WCwGO7Ay2VNJzY
GR3qXcYCjsqkHMdGr7VmpEnA1ZZ7hXpIYnqK/cKgp2w3pCg1RqPTcDq2yGKq
8t0DPFAX8sVxIReLY83q5j1WY25iPCUYTQfXFoAruBHRnzSy8c7SIxr5hJ4l
Hi2d17mLpiEoCA8+sZNJmQnIihmf4qx6eNZDbGBgMH2OoyIcInRXGrIPIVZF
779n1m7aUR8ZuaqR/p/5ZB0wChitVijjL6Phf5nQdDPl4dQ9RvOkrvuppJ/+
n0eQbgsp1Dkp9Ix/mySwXq5c4vAg+bC9BeodCuPR36Q7B0M4r8NohWFS/VwB
UwTQbQWpuWeP9eTwaEHZn8J1F9qhmHO9R5xjPCbKKVJdrXeo4YUhtVxakR81
rEocpcjQDnOP3hp/NZ2QLmN4FC2b9zdpqDROkh+xk0uYFWYL/+6edkDFFOHj
bIyXv/lvtkx2yQXb8R7ivbOAOpugptlwAsdzGDF4zqP00x48juhOe3oYPUix
WXgbLHqzBlTqmxvWkdTRrYhn19nQB99QCJat/qD5+xhydIoL40EzkKdheSGm
pGuX4igOYetjWs40ohUN/jK3WkEXmSekM9iDL1cx1vk7RksrXZ0siOAK4YtN
INcm0+1LJ0nsIJLLpfsbeKnE1v127SXIl74IM8LBncZ1A3/xHoA+o1bYzPEP
4/7UUi00JQbNp8ReNt2MTx28v4dEoDvLEVO7XnvFT7d4/vUuSbB4TMx/wXNQ
8+MouzsptBFTJ1VTJdEaDC3tRAIAEruZeY6ebxNBXvhJTArAoUQx+5x6cNPv
LN+QFcSGjncIWNCSadbWxqFmJU7XLUq9+9pEnnhxjLPFB4r39OlwP408KMfk
FKZQQXhgHzKqZqQVnErs0VFbY7lJdfz3l46ELSQNK4YWhHkSsZ4Rh7lzRtUj
zItqEgWJUu7RglcgxxUGgoZP6133GcCxh76EKuflDXWib59Z2LJjVITq3G+N
OJE3jRtTmFR5Xs9Hgyy0E/PV2OCGzmSgf7YKVIEU68MFTzPHeRwK60cvPKIK
tWrq+m0R2uOlSmlvIv72i7fMGDbUQEJ+4kHtYSZueysc+nWOwKbGKXzPdofb
NpYPjP2x8B/Q+Wfe8dx8bDiAA0BKuHtcUuioqwIc4RUpp3kmsR3t8ETlCFTe
5/PolKiihxwhS5WpjzrGh3CEsiLNAxCA9hJ42Gy2iKweGRGEPQU+Y40efsk1
hTaISXM0J+38sm017+QG9iZgy4e7ud/7kLuatrWlTVwwYXqHs5Tmkv2/+4da
+wi6ZdNWOaEPpvWmkTtPZvPE0dPZURmBy+l1kHlic0eoJMDc/NHA93Ha33AG
tTbqPBuI9OLUd8kh4046hxfyNwM1cVFlTdlH+cF1wcpcE8038m+sdeXX0/+Y
UncpSqrHSkHJXNDdtc05qXdyKMgfhjrEt77kZ/sGnXTmZRCmtqfixN8zhULU
74Wv69N+2IqdjsvE4WE8ntyWV+3TGPdlnFEpLjrVZiLFmtY8fdZ2VuTHEUuL
87YQs3nivY7jAWu7Y8EM1XbGGiR0vIsfDnx7oHlI3EwcoHYrdR1WiiTNRkje
Alx4/halPr7UIJCS3GcbzLHOTVfOtCV7rJDl57Yw9O/ygcg0zR8lA1FVqjON
zs/x/oauer5mIOmhC5q8QTHa6I6ezVE7np02mdCt3Fsh3qq8AZDZslWCiVld
8PtSAN0eftgCX8Swt2xUlARtxseokmU/Zl+bj+wHQOVtpeFF/wwBliYsPATf
ShnnQoP+qP9U8tPJubCviX6POidGSbDIbr+2N9o/Wb+5K9a5+fWg2pTuP+XW
GL5ZNi5YfeMb+4Pa0HR3l+WLWUyBJD7dTDRw0b/RIA+wIEpcnovXwTDeCR2Z
gA2P0iVPteBcJP0HNAL3krX1eCwX0QPkNTlvoFY405HSqomfbRdsPzRRVAZ/
Cyl9R/qqpDEM/IwDDR2XPVmcMyBeJBX0lrnhZj2crDJCJNkzRRQ9g4p94Rri
HV7uggifNg4CIsQtnYk51fFFnoZdCjCndHrpK/8fMNb4IpV8Aw9UpRHMEL26
2BYpWFfhdaKdRWVf0S2vlkn+o9zH3lgB9+UbG8s5tfba5lGERtQHgHQ58Oq/
bbmAtQy5iSCATZSDgYUCvjbjUFH8rJ8/IHyGKis/G5h/53jH5P3W4cN/Q3W1
Q0a53B1PUT1Sv1LlK9kKd2s+CPIyWfVtgBpi9joNfUYfbNgQlnZkBmntqZ3y
sJUhFb/FDJsUA4Hogs66s6oySRNvke7OcpkotmmNjM3PziGLVKOJYFxpYUxv
YVWbTYfGKnwhBRn8172V0f1otu+ANJgbCG4f6+nhxbzOzO1iUK36xRleA+Xy
7kjaqF5TS3nCt03+WKyoowOwoUrdEZve1FszxiaB1GjL/u9WK4tJ6FE+tCrr
fl1TBvS/+rO/5Q8EDef92sqRbXBCvbfGR139nd1w82PyBlZIfC0ps9DaTeGY
uw8A5jzStsETr39GsZO26wRUfgUWZSTq1HIDHUbV9ixefgonAjQ5LfHWIIO6
apKTm7blnjnqwK5uPZADHHPpeuxG/uNNH8uzUTcrQ3XYw4FDCBH26JndtQNh
nuzlrm2sz7+JkJ5wzMypGp2aPP7tpe0iBGM0GL/N2AwnwzdE1HoXK1an/dvZ
SPEdbMT7Pq5rcsT4v5h6LtjRRJgJyLoGLbvoI0TlAY9vVjEyZqXV8/UL7x48
+uj42m5pe4WRatbrmLKFZKJrybc9XxsGW5RObIHx0okQpPaTlOISCGZRc+jl
HAnXtqEtsDMSsKWB/EodR1Pw9Rq/g9D5PRj72MJkB8WB4d629IcmWZj/+xNU
GYwh0Z+yzKXqI/DwYWPVX7bCTN54eGFwU8v1eq/4KtTFc4CtfOT69HnnVxFZ
h0+PQZ5q9vCFyuggadQdYsqJWsvktsaUcx4PRRFbS1HTOQWgLhG3rpFdghOM
jvZsbSVckbHz82BYukk4DC116vh65xWByRErAcGddhpu988iAxWk07USakol
c2tyjyDqe4F10vQ3qME0cSKl3BrJZn1ewekOALD3v+iF85HxbqsmifsZxxPl
0boJFZdSLDPGxIR1OT3o9kijb2PRau81nfN2MI/DkWrDyicqa8gqThZ5yZVx
fmcW7emY7xpMz/5sA1AT/55mQryKaFLuElVoCgg0/gTxzW4/ef4tCsGOdFeu
rJGYN8BobImu3q/P5eF59R1Rzqh4l0WrStk/krCumZ5q1vk4ezLZQ+e7ylNg
+yz00T42MxPYxDhT4rz2ewDyiVHOiqUK/qIwDvEAYU0lCAntCfJ9WmbMEobr
WhkiFB4WImQIWP1TFh2hgcqMQQOPMk6srwQktEJmPMzkRPvTgE6Gb8j/pnkf
UVxwYybAXjux/rpMyPTXes2MqoCkpPcC7rE5SuiHeQjW3aWIsKLdUC3Zu1B1
grzTfLlVwH9BtPef54xl16EWy9Mimrw1ZxTQ9OXjfOJu7eIq05GH2At9mI4d
MYY6bB16Ds4pqoaSMhHSmptAaj75o0aZdv8zz7563a8ONaXfhh51562lYCKT
KzJeBleAfObOghDKBGurWRzPMLCBmTQQ9R1FxlMKhkPoIhOGP3XvHuCx5YHS
CGNe6X3JsArVmzSFy7FmQ0nNUXok9oSCrWt9jjDA72m1nGw2ayPHsQURRo0e
49N7bF7B+R5uAhLAyTrq3zaZOJMUdkMcunrwixajyY0VRMvSHyMnMaiJSRo6
/Yd765ofMKvgqN2RBYPzM3Y5DTtPF0HNPr/iSJdMUWjB9YoeKf0bkZP4WmAm
z3+pRgsgQ/albCbvhN71+6SMwcxRVw2SVkeaAM1p8s4WcEYnk77TXdhMECk8
YKUHBJQg2K2CWI7692ftZ8fIvFSGJnMvd9P2e+zesI4a3gVwKMnmzt0j6X+s
7IZuEXuEqjG1aZTStIMm7JsIKjKVgPXg5PVd88FuKTEm04lq5G/r9tWklV6Z
UY1UgGxPND8Jt2rCwdXADEcxWW/+crDVnnaZSIt2lvnxHr8o/u0oZTSSngUX
cvKrlsOwdkSqPhC2rBnBkmOKWoSoLVrktErtR/X1R3ed+xISlmp6W6RcRal7
ggzlzQGru1dXaj27e45XzMsb56dYL+2+5dgG4Vz891HoTA8tIfaLw50FEIIV
L8//1zdh8xo0oOH1JxPGJyM0Hq9KcBSwQkM/ketF8F3ZBc3p71yDDcfCqeTq
g7YSwrXP6Uus92dny25llNcxYy28hiSZyj3eqrx0NeAGewyxFlOHKqP75z+J
ZgTkF0gjqwaCrVmFuxc6vnl82i7Fn3eSO+sw464QI4z9XhwUs5w9Ln0ZcRAT
OmwANLwUV6e0XsP0Lndd03M30qCtkscGjNo3lm7eFU73MZuu/opJg/Z9a2M+
FUU8+o8hIgPZDUaRcHDyWKTcgPZP+iskyWcTPDfru5iZKYn8b0H09t9TEnLC
6trA3OpiBlLGjz/YWbo7rgCuyFoV+hkexpW6GBRe4OCTZ1V1uGtWyBsPncE2
1f0s3XYMhcq2C79INLxV3fHf9yuiF1eiyRUGBOakkZSYkP1Au2/BBW4cNPl7
gcvT0QRxU6qzejliWiWQQAlkYm+BfnGIQWURPWXENQolNtlf5rBdyevsteA3
ECui7kM5dzaoU++c91g9tMyd4gADYdg4dAuROrKI/+jWssHcTe5oBRihBapg
frNPJE48CXc5K/kZHOCn7OeifZkclNqajyeAgd3mYqrJkSkeTCCmz6H8mCxd
Waf9l8fUBSFwp0AQVMYp+u2vHQls+Y7ficTs7RpqeeLTGZzGe6UYfwRJpH1l
Y42U8LmLC6J7qMJDDB7SOvuj5od9j5vyXs55oKojggcE5pFjUMBthvjmZosu
5v/jSSBN+5XDBnAJ1ZvLVdlQI9Yzj/JHKUtIAShDidarGzVZ1lX28hdZLnzr
nCbiEsoUupHVTaaMrLIYHRaCc6p2oz2KmsHHjYGnflEExLciWYD7K7lo1GlN
zHegzHbLY4beM12q642Sp0UwUZ+QR8ANPds/PKvEcjLZo0rEZfF14OmJ5C6x
FODp3hTBiN9z3NOAVZGASE0n69+iDZOBTuOOLYL5yiEqvEInRPKphKXdgsUK
WGDaG8M5IXo7ZvzipBWMEsHnIg24//74PM6jl4M4opunJwy6eQ+bgGQFZKpE
Yde+iFR7rNnLZoln4TUL688sZRU1dvlEmA0T+3Ju1anTw0afOuYLiJW7pIMU
S1QUtGQVSF3QAVz4lIowsBfu6D3MhrKEhh3wkjPii40/nwnVEskdEVaYrXEr
MFUqStYvKin2lYIVipsL276shPB9oOIWnq2VCewlDRSnmNmBBMAOeflrJB16
IS9JI+GJWS78+oNPIadj2awmSCg63m0jcm8xv4zc0b6fmkv6CN5sfnFDwvkf
qmdR1OrFIF5Mrh+kJ6YMO6MFnSVLAIab6WuZ2vvZcHFogjwWeQyTssi41txx
ANe4aAY70v0osVCpYqnMs3OeiYIWH77q+ANc05nXJhi9J2veTcM7Hj7cPXGj
McGHEbvxayQXF0Dz0i7bi1Gj9oJY5z8SLZjTr7OsMHcsdE7s2BucuQMsqf3M
448m3mL/rGu41oAjMK8BPlzYY2OQ38X8FTlneXjMDZd8KOizMehObArtDlpl
91r/eVnZ999RCfhRVIyFINJ3d8GrrJGFEl+ghZOCd6brgQJs2b8ZH0XEqvuW
PiLotADR31o6tgNhL33zZWIPajhA4ZFdMfyO59pmwsVnDREqgM0cJtnDx1Iv
pu+EERbxiFUuG600BuilL3BpXuzjfor8EsZwFGnEDIOcTWlquWRC0xIiyock
9f8KAWG9px6TBhC8UjspQ6wlmncYuy6JHjeJiw0wxoZD23V5sJdr/rzPnnii
FAPxm8oLPVDXdQ68XTDql22BuYOTrvrHvdcIbq9VDD8gmKUfZDhr656MNZyJ
2BpJhVwn+uiNzJECKUqelG4YWesqLacZiv6NQCSgQhPXd6ReiXIo89P2aHbV
5hizGDj3OYgrKuz03230Zkwwpu54fUc0HXscPChx22X1IJE/JlJUGLgP+oIN
5cl7iXSXpJwxsb/TzJht5FYKt4H1G2OhA3us6k63Ak/N9Dqk+6QRfSYi+oZY
eK9/Kx6J24CVJNMwXB7k95CNm31PSvexKHU7+ZkGeREdQZyuhQiQe7JR8bBk
JQfFR3c9hgCc3fA21c5z0UjT2Od1o1SMGUEmndZosMoD2DP/fXJ8zMJMi1kl
/oyIHLT1ZFx2NjU9TAeqYBBAw+A3/pvFeo6YiCulV6HyPpbUquuRmEDhiPcD
v03HeDmfdjpGnr4MUMhs9xqdSqo0VAy/NjhtdH5NEg0uPAAN3/fE6mltpPab
os7pXdeupiufXT2PJFyTNAihajca1Cayn7SSKxpV1obCehJb8pUfwYSQ9Bp4
b9z+FUJEWGNileBcXF2XVIoKydilm+WwiRd9JQsR33/Ej1Cr5j0dhNhBK4nm
WLLtiJhw31pudCjIXBV3ZczEm1NxmYti3oDFEWSNr5p/sKAshrqWKigycGRL
j/v35CgJ8zxkYsegvQkiJF+UdVHZS34zH/temOVM3jb5rWFD/U5oPtTWYFSR
XlrJzgFyRJCMR3lLv1WSOkX4u2PMij+PG048j3qales/S3d+7ZCh/A3zEUQ5
H91cZfhgsIWhWgOFAaW5mojNKoy96eS79oEttCwjezGsd7XtMLYyVPAMyRGR
tVsX8yZHH4sOAshx8aIeZh9uZm4B0C6RNub9306sOZxYD0dzxaIHqwULhIVL
/DwQ61wrtIcGi93QneFvva2wDQzlPvtI+DeUdeZQVYLszsSguBnSZVJuoLPe
vte6x4siqD1DLG7FayPwJmj7/LM8K+T6l2F5qyvj0RE63X1SdmR3CzOzPUuD
cD56djvFhJxUIggJ9kpV2BLevaidLL7NKW6JJVMZyxwFa22AeIwnVa3EV5No
VGokCN23jEiGykVsy+mHDmmE6FeDwCn2x/aOag0CQXbrUDhTw69UeJbHpd0o
/reLDS2f32BjWOVZ3akWMZXRuLLR27q4MPiC5b1pCtM38asZO4Sz/P5lLYX9
a3DwZJI2ecJVEMFGyjq8pjCtBUFUPD5OTZvJI/X33Vxt6WrV/iri9RnUBaGz
7/fjQL2c25gk1FtdwxaCJw7ojMOim87jQrsZ9S3Tdt7QgxyXxqMuO9VsXFVc
PzJ7rRvBVu00dl5g4Hlt4VOsTMvTBsaijxnnWLUSiRSPobt5a943FpVy6G28
4oR2zqMvjObHmhK7L8R6tqT6sRX7x+f1aUo0HHSIEzzZsl3UFnAa2iX8HZBo
t0xmIp4zj1HYDox3QC22K+Ty/eLa/785pulJ+S7z5Ivj2rvpaE1A1HKccW6B
TY4arJdRCPlos8ymev+Xm681HTu4kgHaUUtBaK+5C3riUl7vqHb6N4s1bWi+
wGQQ0NGilQhFWkWtYooUpzQTkShtBO+9UEgmlqufxgJDdwFSYRjru8C3gbgb
n+5b4e+VPiiD2HPHhryY+lJLL2yE3ltpw5rI+EGVPq0HQps8jm2M/uTSBGfq
FstiRKig63R0eUXZ6gjHKDAJ/ihmjTKB0Pk1d+H5D0MiWX+x3vygozhNA1xk
4qU9LkLm8uUhwWosY+ivt0Ln0wBx0FR0oP0QuWgZjTcRCcmpevCf5nt0XpKO
GIEbKWufcxd1EVZERq0xPCIU3WMoSr6KW6n7hVSbG0Rq6I+4h6qvjXtGcD3v
tjMKHiIkUQOVYnbZ0IanbZqfXupOfHug8iGaFDiIhOvzPYMJRGye9ktABm4f
opD/beTl4hkhbDSftEaKLQPJGNah5A5bn1d8H2NUZJel8cs+t/VBTvmrP+yX
9fyzsTXAQCat5AwjXx4AWp6vyCsz5ofYisZbk4QylybaPqkRzGzDozYVnb/S
RTXLoIQx0f7A+T6EbNbdE62AxpswUmrK5mFsF08wveEjgk9zgsAfbQCroyxF
UTdMZ8jnQEFiyn1Yme0pniN8HkyUzMDgfo9ukAVkrfdxxjzGK1dS+Vkc4UDB
92ppX0DsxCDT2w27TGXL7eo2nhDKJxT6sud3qLtHCcgzTRPkzTPT5SWJKghX
ypGF44OqXYkTr2KQcN/Rre6QQagKnjKyeWZT2lhqMKcuuI/NC0GX6u9Ia9Ci
o4XIbWlV9ckycfoSkloxc8wf2525OIolLLTNfOKW8o3Z7brZoXEytiAwzYqO
sxCHDye2KPk6qoJU1Q7AT1cdpS6EJ63W1OnTbqMN8oxIewfU1rmwlvONtrzz
bFMTYafsIKaoAG3MlJ02K8p64sFN8cD3Pna+/W8AYVv+xcEm42NBUCwgyEiH
qzpnEj6ucCoTONk9f+D9R3JlZIpMj06mkzKDUlvE88PRxeA5eL0p53D2JOjl
Mh4DbkMlAFViF4P8GAdHt7xMFp+0UecwycPCKJZ1ZacAkzrUCqv3YLCHmW+5
1GS6HOWRizSSURJKb53zstKPps5wG/nl3JDYiOVxUd0AuxOvpZwWkolZBgNe
S0BrO0JuYSkOreXTkJ6z9QvHZomYG6vPXKOgLlRalQLkJuhEXzgz52qDMNgs
j5KPUfc0Z/LDxXumPWYtHYpN5GGyQWPsSPUQigD0UNg/z24idSLYUMFaTdn4
6tB3fev1uH0gvhBfAIDepMmp90tpkka7+uBQaybHolZvl8JoLmOkuT0jBdQb
5HnpvSFizQYOXq0WUrALGTd5YrmwbuPdisA7u6Xm7e7RZ3iASo9ogoXq+uZT
bwXp/IGgPmEFBOOkj9VE711BZl6aWMfg8hGF6msWTDbrvlLur1QPnc6c55TJ
rMDaMuw6X1XLiqNhq7gmTf1GkLTv4Pm9+zXDwdXo5hpinLEiCYMWwA8y9l8k
KD4s5OXhwcX90r1Yl57nfLvopaiWuSbcEHwDHE1x7lj4/T3lXo+oHH1pQvEw
wvvs+cb5yVDTTzXdkcO4qj1LszYBXsqBXp0tbHnQNnAnv84Urmbwo3mQ2C/c
7ajNy3Y0g23/PvK7yXr1RSIJlmgBshjm4wNkXTb7gKj6iOOS7vRk4xrpGaIc
bFj6EkttoIItOIxO5ITadZ44GG5lfRmU0IATUSw0OBzob7CfSZ1fXIcF7aJG
vEUy8W/Z18nDEikwMQ2z0GIWNSPAZpHCtHi8seNSvmQJFfK0qVaDCl82TrFI
7TCkogdDR+7IBQMhHAyrLI1iKjLFObLSmq7scQOs+6VjeF0ugqaRKRYh0x19
Nyy9JX0PaeI4HoxUvyKFtOJ37uGGPPfXzF6+OyjpxjW1/IcdWHr86ulVq/mu
EcrUJpn8fvnzNtHkABe+pD8kOmPA0ksMNdqbK9RIBLs6jizYL0IiSqJIq0FL
rxCFxwWNIo2tlAMnKxkgJU6eaj+AG5IRGH8XWf0GJR6MsVfStTFZ/KgKo36G
a20j17/BvseJN8+xDKWVXz6rypS6sHwP0DKvggyGt2ODJ+25X3iqgOy380Uo
Cx+kcJ9Ox90jTrTh4Ex40A4XZYgfdwLoRhqAIEonRI6mzSnixvYm0qcBaz4D
GMBQE184wwhwgi/U5X3JRhWoNZ54iPaVP1tAQnJx6kTy6sf0qxNJ6ogtC45D
UpShLWtdUUgEgk7AdqOAdvmxbxMsKDP4Q29/zzRSn03ckZkFz2k2DuAkX/5w
nVUQ8ypELT38CO8m1Omb8ZtoXOZBidq35z7TeS9y0WeLKno23IRk9nE7Pg+c
YJkUjTwakhNZ3E3fZKUiNSAbV0wwwwNR3jnLdg+MdFlUkCDHobwI4+gOzEek
WURCVizZR9oVK7Htj4O5JFF5ZxxnnDQgFIkgrqmipBS+S7Igs6D5O3lG6e9y
HREiZ7DF7r8LJ1BI5QhCraDFo0NRorbgxwfhylRHpXvmJxr1EXFyP/FKSGVl
+U+wEOH/L1lo0jCWndKNBcD3fDTfO6N/Dt5W3rmlm7Iu4yl5nLj1pZ1S1Xs7
B9geJwbtViE3ZRpmxrxDm6Bips5SrSeD1TKu4UZ5n1gPhKmKt299yPBu1epj
Bg21qnTgAYF/1lFBQhpZJVNnlktqAZVZ8kUUDrKxcq24xWQNLH8pDxvALloL
lvNWN6T4t9wh+i/aSVYZzBrE/RQDaaC/04Hig2fCMZQ6a7alwZXyz6LaXeth
SvYiigV6D6WX5jIfZuPjZdbkSPdug1gSGZNW8k4XLLzvvnjpZ0mrT3/heWHu
U4VBV+UI3rTdwhvaJQzU7att3yRm5YBQZU2HyBptmFPt7MZ5fmggdIDf2iYr
uJtui6J6CWke66bO6Gtnd7NCsTsdKQXzTTsFo2HML1FGM6Picf2jxw9KLfh+
QgXZZyBNyaz2SB6jt8IyTlvFLQhYH6MpEmzUN3OPIUDdrmvquV0EpKDnPupN
6VfroXkCPSwfOcUsVYa81Xwb4RuDjxD5PuB7OTmFOf3MHNh3+Yj0xV+H4cQZ
dVUoybT8DuHdOTqbIYm4zC4vMbcUqI0DIjmQ66Th3UnqcaID83EFMgFwMjB0
dc9213KrjjeNBi8NlfS9Mc6ZF19rZalcHVTbAxlpIV+vvIjpNDNIOXRSQADr
q+SPxU18vZeoCZJKNjDgdYLGcojIq/kNYnBG+2c1MWjr0KdIt/eHPMKCaSQV
UG8mIMHaImubQ4NKTcuWZXjJypEU8U+RltkYV9KjyUIbwc6ysGxMmizioWM9
WYzHtTLngWlYhcVqlbx5mKY/0Esh/Nkm04E2EGWtfhk/eUXF7/1eZm4kRzx+
NIZKvy0t1NIz42Jw2K3ABtAp9F2vnoAld0RtiQH2WEKOSkAUvzZjhJc/nYqI
w1WvQXM8DtHKzR5j6iU3KMTtJuRpAl8Cm2+wQfdSakJnynHCkaGh8VfQxufp
rbqAed3lDPLqmbv/PRSQjSBPj3Zu53mxufniqDQyMhFnCUyjh6s4c5mBiop+
ptjcq0NJi1cbpjSE7QBkA/eN4Y0wz3EmalopoiY4q4GfB9fKrr+KW427Dp5w
rRj8q6rjYtpn+W1F+KyJ5jNrioTKRp/MdZUtmKTLWJkNfhiqgKw9464mJEGN
Ve0bLbSls43cQeV6C7B3zbR/foIwckmPEzmkcFNsElZbil4ooPbhBg5m7e4w
gjt0I1SsN+tvEjvke/H2Zimw5vcMLmpfA7hxi7otEQ1cO3O4jqUSp2oa9yt7
bS5hz2Lp5U0lw89/hpFRjW1FCRWVoMd54sn/6TJeYHRNJBCD9gNrfl/o0IEX
ING259E2MoFiejaSfLz1Mqp/rGvPAMbkvTdSn/rFHq/3KvN17OZn68rpDo9b
hrEzLLMCNXoh9M+BLey1vxk72Un+/8Qv8toWlEL8xzk3rV1FuO99YckN7dhy
1I8F3OGnAh1DmKB520TD8gNXPuU3GIo0OU+QeYBC1JyfnqVTnEEZmqj6Gx6e
UiJGVvHwTaJw4zgj8YmB63jMsy4UKX7mrtktwr49b1zTZHFLNf+Fsc6EgmXG
0IsrSJHKulp9r90hqSaElKnS8D+XXcBS5ZRoPtmne7yK/nVL2XUHDZoOHC9t
LmCiEMV3l7zoS8FwZXjZA87Hq4fUpGPC1pZemA6GW7JFvZm3bC+wMh/bau5Y
VmHNCCsVnTVmGunlhE9Qb8Qx5ZRGy9dpkolOF4KxpVWvh52J9q3UVWplttjC
hzKZeQ1t5eBEgGYmR51/YpcllKCbkxEjeAfkMrIzs5h89NJCjySmLPBXOX5M
54xMxbFHwnw5WuGYHFBp+5t2L7qhqZPN9wWlp9aQnGPlfeMd2XjXzD34WqYf
1vK/fmtVZJdYuxgXAwFhAp18BsFtqvXCk5/CpMFMjIe9FgSfPEI2kbQdQd63
ycr7uZOO94QDO8Yk0JGEekhTTcNdUesOgEF7Okbvab+ccndiCMgb1pWrxaAI
l9E8RHEkaHQw3zVv2/rEFx5ELehfRd6lM3hnl3wA9SagZEFOFUkg4FWbG2oS
0YNDdXM4lo2V5ZbVUTvS1z0ZfmhN4IahozzgMqS8699aR92OqbM2b19N1u0V
FB726LfdhhXvl0nT8Uq0EQuOkjsWlMJPQEqugTZmWC0Ml5MUyzcISkhKXfDl
UJAzYee9dmJviNOTyEWejtCQaxkwTrjH3YK3K68P39G7jRahsRT0Xl/hakw2
acDRLdM0qSXmrLJ+oVUlF4d48So/9RM6KkkJVrW0hvd8gaLy2B5D3yB9HzU3
NUrgHEowL1fSRy/H6cYKkjBDVVIddFB9f3pcqjTqbMXzPLWHs1QzeolNbWhz
tSQQ4OMQEJQ7r5iQEIBLZ+BBiseFqdJk8Fj63PX1EMaRMbwQmqnJazWPnMNg
uo4AiF1RvuXL4Uzmri/gCDOX0Z0HxMIsrTWzibn4ppz0l+BaP55WnQvVy5Ta
cbN17r/nadrknQ+nP3WcPAlOYjUsaMm2bM15vKGLsyPmE4ynd9QOsK5+u/54
HzuMS6iN0Ps6xSiJlGHMuMsYwSy+EGh69g4AobUL0sBBJNkJB1X21+tqMLdy
bt6xDPdAc9ry/BDJgKXDaXhxjWdxMcCW5UIrD4pYnpflj7UiTlZl0EURHC9E
CAgOZJ9p3towIOHnyufXERI+K5FjCkQTcw7Uaz7UwqtGJ2tgDRNWDlg/V7Lz
whCunT05jQfVkKSrI2bt5hvXW4LKVuffvlw1o6E6WcRTFfJTq8GK5RF/AY27
JIEvmzvKxRHChkP1J+lwvauwm7aB0aeAmidwMGjXUjde1+IKrXU4m8gJoTDv
CjiIgnf6gnP50+lEtsDYHaqYXu9p0cfGjczzoYujJ8POK7s4ZVY4NrjZNkdA
9tfMODOHrhMz4DbLW3SuivANRtnZxfv82c3gXZLGloAzATP7djMpLs5HiDEk
MCpBOwEb4vglDvXLey9sCx4IiMJPmqLa31AcEYGRZNdr7GSPQawi7c3dCUar
GsWS2ygTdMUl6Mz/87O6IG0rrlhd1ljlYuD1HxToKkdJhsnUpFXOfbvFgW0p
4LNQXbnHbCB6ZyhFCTUpIrHScfkbr7NmW0s8WmHvF8j8GSCb3SmwJyA31uZL
J23PoycMRY3obZSB01nX9Lk4obGkeGC3HqfykR2uF5O782M9FqTxkJ6ldr/V
9VWvYParH+hevqVNFS3p3uN07rpGg86unLLKBVyZJfA93vTQ4Xq6qMTlCAov
YzrDUtNp3a5/7p9sfTvCUY+B7XglZziSAf43Vkj/8ikQM7YglIIDqGgGtHVP
w7MOLqAT9ERXsd/woa2vKnbW6ta8VgGPZbxP2jmPN4bVw2ncWBbW+rTgkC1X
cEC7FYLavainSC/IdKEqRmU8/lYpmVBF7h02c5592i1wlA6a2UAAkeKiKWBS
bdLFKjAYrnLHcsV6eGK/JDWDwS1EQP4w/UYgO1Gmqq860Z/wg+CGYlGlJj3U
euPNWAk37p2mUrSbhviUcFp1HwhkeJ1OjnB1PR/WOqsIwF24d/9OPGl0UcYq
23P14ond1PRQCQLFLjErXBV8CSlQ2oqmxDcjWC6uXye8rYg4T7iMkH9hRiB/
ZXClpSnqN2LklKXudEH9rqasIVptJuHg5OFwB1fm0q+HgIRtH5w/E77+haTw
2A1fiFtglTbxuioba+GevRAjS46VtKUcUyhMpa4VEk0fgcD6cBv7pS14zhgO
bVIKWZF28+6SwvRTfV+zVoNqolbjghJk/0g8shHlJpUHniz//W+ZuM89t/xS
mbpwpxHmrw9rbs2GUfWmJzvowQG46dGNT8zaX45cA0tRv5YSiHBlp4Hoa+lD
YNBid6kAC/pKxPGD0DdiVks325V4QcXEzLVT71x68MR2hGCXKettEmcdP0uF
fqE1TaP1FDXhe0mZOUlr+/wYr0z+1N2sBstp4Nv2bgrP16qZZJaQMJnLTB7C
aC3IQsCZGq+1z7/wUcf5z6i9ZlyGgg/ZhxaeTJk/0A==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGMX1T/xxPltATdG4ve4HuJxxyQuWbC80WQLrEFHIC0BqiQBeJTRV3Rq/8kAKfh5YbzgFo5gIZ5bq42LdbYorxyIa4sjUgsf3xcPy9T6uBljl4oj4qj6JVmTh6nNTU5s3FqVh9/E2b4nnVYsL6sWNQe3nrTzSN/gXJET+ghF2LuTvfZbS8sifuyT/cU5XNkiRPscoYX6/MwbbBRivS2T3l3SjTXxtA6l9rBKfBa4t3D9im1ZEe018laBcxlCuBN9e9AIf/jECx5YNOPF47NcC502eh0CW7e/jmchr/XWjj8ftBAHrzBz3FYod6nnQw4NFxaipJxKFPFVuxwb+WEQhhUSKazI9jvu+GzaXGc9gGo0SyA4xqJ5FQTeT1wMtqbkVStOZNI0L3uYmgySeF+qLL3WFhig3R9l0qGGMTuZ8IXdN1sd+TqUKbnZDya1ruLs86U/pBSet7tbbSr0nS4WkeM1xhmsm8zb9MbPCZGd62J5+nXOG6O7Doc9l+NuQayDo7FjgFga1ahQzQdadKQqRSwOy2bT3+eB1llMhzWkoQOT8LuPY/SelXOCrjespgccI2WE/SBIIYmgBqpeXAv2jyKxae2kesPTrn574J4P1F7zipuWuGoQTGYzaKEQr2Osw7XuOB80xTr07ceh2qPg2ttdHk02WdF/Tx4KLbk0MLuqXuVO+KndKg3X/+7VYMzGesG0gRw9CFgf+68Ro/tlc6SBRS+as0sD/7JLafIh7f7UD2gxi61+wfO+f3difdk4UettKx8nUBhTwKhyDlgwTkCA"
`endif