// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YyotivqAZyCltIRZFoJmtPrE3IZUzgr5rhejNLv4uhGY9nF9IV2w9KgaSAOA
l7GYoxn5KmJ9EPrAciOUG2tqFCLV2GN+J3ATwPg3LxXAkMBqf2dqasIGkUoY
QjElTtu4+kUuNCk1EBoZN1nqXvt2Gz6py680stPtS16I64hgE2Z4JI47sSUE
uLOrfD56HE7WuPfX0+6sLrYEEXAok/DnpfP5xx6zw+vIHteRnLfzjfog/6Wm
f2sBtqiP7QZf6fS24lpqnTcyRcNVV+wvvaz0MLb938KJ+UNAg8lOqtgxBR05
HmD2XHRYNdLbKAgk1RY2D2vHbHc4rm4WnY586BDLYQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZCGpZEBGQJsN6HX0wDv7pHjkp16bzJSejgqq+h421EHdTlJ06uJDM/OA0PEV
uLL2vjLGId4UoSIYG7XRy41TrbaCTXN2Dr4YqCFPL1O1dk3/MQ83whqw4uon
H+Oyxqruw1ykC6rU7FFOFRZLzoWPI7vvDQ0SrnMEl+KHCXLqqCxQrl0VOOWY
xXSf7OwLJaakA1oJjDcQb3osvvv1tu+9YxmcTzExBwgfaopTpWvAvkdOmRT2
ZxpPysnaTpgGAaIDD1reoFU6QjnJxeiHoZ+3HvFFCB/UW7pls8fjqHVIAFsu
2U1RTHiWW83BR8YQED0vtbH4ZregootiIwibvsPn8w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gunmNOR8limd9riXExO8mOkcjLAlBEYIBADtqDYH/z3PfkcStRLi1nnbHsWm
+IvguTqz1ByGzzfHZ6/FInHJ6f+52oKb+8O15O9yCv4Hy6A+kXTgU94yftFm
qrl6B19nRhyYRDiycaK5mX9RvJPdb5iOHrGp4UVEH4DzIAB+F1MeseaPMFQ1
LfIAwyPYt+FFSe1Tha87dpbBHWwQpdJdS0tl9dwdca1AB2MQrXEpKcPU1FrQ
5I1xCP8sj3Phrkt0RxCTvz/4W79bccB/X2XI1Y1FhHurIh19Pex4TEoiVHzA
/VDaFAuKOnVpW9/rgQEFnR7tTtLLivDQgv+r479tmQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TwbujmOBKMazzYXMOuWThcB8MwN72XV6yYOPq7zmk7NWfMep5mx8q3FcAwcP
AnwhLIHGoF+GOwzR9RRSmrWm17hhdf2b7GlVo/bqkv0250FBWJf1uBrMswC4
ZvzwfClfWKj/Gmp0rw8dC0Mc0wtc+PNLrmYiNKXeG7DQ43bFryXfXFJT8GKo
8ub3hA32kAuGwOlsWe2cZ3S0TmZ7XGv/9tRoe8RDmoHXUUuqFaAFk8L6wAx0
ZMsCj/ObjALkEniI9lwRjk5L1rTr/OkoHYMQlmq7z8fkUrq6HWyUNj35gnTF
UxMvpPwb6ONcFQ8eEgLMcwwq2AiMFH5GibGOkAtg7g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mXYEScpaTHuAIyKzRWEuuhl/dA5efZPmbaL4fDTWLWUI6JCKOP1Xba6flSSC
dGlCYiV4HYt7/PEMP9xIYYSPv85C8NBRvzYfP9WRCLz6mLbahExMadDVG4Eh
zKj647WYvGkKEl3ThL/NHPU0F41ixsfeEdCsL/djGm3oNiU+WPQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Z6lQc18ly9Rmo3Rb6GENMYHefx/d0WSIMncg+vt9jSkkWbDhAhrYegan560x
b8k2l1wLE4pmVF6SumjRLtKcvAfDfecvObUx2Pacg+Blc8XdcynGjGXod/pG
E0O7DbZnbmLybA0Mzl8kRYrOctIuHNvbDwhmBrnuCpYC+tSm/cqTdWHZGVSE
fZAHKzXbsZ1WzcksJAJULUvUOTNlC6m6/2WvY0pr6lPb5+S1LmoXMVou9YL9
SDn+NiDcvZ6qMnrKCFf+zcaFCuYjgmk6y0BxTYmFM3SN5Brva5waA9re9lNN
0wDel064XhZbyCvhnhJFWbWBmXtIpNyKkNCUJI4KiNUArEBBa9ZkNWk1TjM3
D3OYh5Y00tFQXsektoWzO5FEbssUlvEvJy7xnAow1LggDkGw3gqhrBArbw3d
8NNBxxMM/qmAcUyJ6AysSmZyJ1HNzDq4XAdHMDMVE1cvpM6s5s5kjSEvaNxp
JZDkRXjonHRQPXxcL7T3yym0QOIfH1PG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T9Tdglo4VyflUNzVvsFzwNUoI5hJMLbOUlbAo58BBhE/nh3qDVercE7dgk1R
X+zmXuWg+adg8vhZ6VRR5yshN6sLdF4yJrcN96i/nzzMdF+Cd3e9ATo1u1DG
z+F4zaBPOIm+LXKqPvMKqxsY23ZyVOilrivk7ABWMnYboYlFfsM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uT98O7tLlfqHBxK763dUxfSp9ob95BZxwFUVRpNO6zdn9wfxtfT7Hf/A6cIS
Em5WVtFvgcPYX0tO2kcZq23YuNv4uchNEaubv/TP5SypaFHUmjgQRCIqtipj
qI3f9KgFaqkUT8bwkCAFgodCjNdX2dXS6fqwCLJVU6OlLg+H+zg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4624)
`pragma protect data_block
TvTlluj/k5wCHMBnIVf9N+dfWlK7CHUji7hYQp24XPA/zUQ6e4SrLXwpBLyb
jABGqfy9ubhQoz//5dDImLoz849b80gPSyW+yK4lrSu9A3TMDvn6TX0GFLpL
6aBwCkyLzUI91uRvLcibivDRlE4fe1+c2Omstwm0Ck6u2dj3p+4UbkyLZtqI
n0L5btEFx8i8SVSz88G7F8qmOA0ICttxL32LN/nE5HmrqQUCULg14cvUyYB5
cpp+dOC4RyuRVsYVekjcFjBtDqON1fsnHqJU8S6y7QYnevB9tMZjrFyIhXJe
NivO8ZUMOi4/36kSrJK/zWSae016D10Updyj1FE9QPDGHVcD8pgFH6caa15f
dVqwIq/Op8tI9XP37T0Xu/JqUHyn/hlRTMT6+kLe7G/3z/9luQVlfbVyrDxJ
/BVJLf6Sf+pW5eazbTVDDXK10Nr2CzP0iHYgtfYTmjrP97ghnj4k9RlaYhk5
5IdSpknCuS9o2KiVJpIRUTR3w/46x+DntvkOPELBX1s+cHptOEYS5BZ6T48q
xJMlIeJeYWzaYoDgrh9ZbmFTkndy4hIv3ebCIGGMaUO/LQbGZL3tR8wGzjZ9
3tnGPEOANlAXwTKUXOWYtMJsZVy0heqJc0myLheeLQalYdwaocMor01zvKVK
Gwx5x2FqYnNkvSDFmVtJU7ohNVXO1+bkULDKwp6ecvNpOBS5PTzMOEqwa6cl
eXfGIHuQJLMs72OFtDCPeebQF+FdfdoJ/EOsRiEvDuAQnu2C6SxzJAfh8TPf
Sdsr9z9qIzxhT/QBjLLnOZuy3gVifrAjih+OM68pD5x0ps03eADmRE7f+Zw4
nRu7NLYxQUeHRp8ERhOFgJ+qwZdjAQBocN171FSn0/s4w2xDXVOxXfSQk2Bf
Az8EtSgTgCFwD1d0LK6/ZVyR7jSE+iOoGPeA8v/2b00ddXPkLGku0YF9d/C1
T5fGo0Uv97h3/eZkMBdlg5rwDgqEf0RK3hHxyc4KPnR1Ee8heiksZbJU8GE9
GZ53sSm7SNtHOc1veePSrKRvsiQ3j1Mu4bfLqNIr/4XHc2Gvax2JTooFuFbq
8b8u1PT1F6DerEW4e82huecwpG54Sc8BVxSgytm9Q/xFb4SDH7dAzvGoEMlv
13f71VpalTPD8p+Otxmk7wIvHWASIyLr97ZVkL2koGMV5aTroBdz6bP4zmBg
zFAQaG4JpAek4TwaRQYIJOAMdxmtq5Ldwlrr30yTAthF9m3c1t5FjUNu9560
1G/ammBbp+jQwSVSAx7K1km6rSBDHGvkowN4KGV1PL+jCMgPxxI6Xand4f9J
KRUW9e90+r4qxzXzIA9SmFdO8l5xdRejkzwpFFIUiU8eEz3vH1lGQZuW3iaZ
T3TDUrmkd27sDGimHD6X8Vbezes3cl/cfuX9SFCz+dBe38SFyJCTP/u2hoZH
RqZ7RKa68PGDox/kocoTkrYfThyc4dyZVJfs6v0SEiILhGtuv/PFdV7T0dbS
URBkLjmr5eCLoizeAM+QTpjOKo7dCsl7/3f4ors5bkDFPRdHaPl/EUfxS0tN
z36fq6HHz9rgG88Hgyy0BJoN0qUJ7ayQYX3uT4ayymV81xDxqVDwvolGDLke
xyacN9u33hwsAJBJ6vHbBlIMlm4pwpBC3WXsoRwzdnGjlCxY/rqbfKD/cmmB
zAi0tRboOhKhWnK73x/vdfSR1EafEQ5bB7Y2XDaD1ULgsGjnVCRJ+rPIChp+
wMxkjNSnYZMaNKSdktjTryhRkOsjWjIhT0K+9qnVBRrkQ3+LK7rEZgJ+UfL3
GOMxhHx/bwl9ZvXsUT7h3ffKgQFN8ZTwH2oARLMTdmcLGJ208ctQdgsVvC/z
u8Gso+kECdhlsFZGnqAtYDR1tnE0AtgmmhwJp9skHWsKgcTPFZFi2IWgDf3f
8kMT3I9k1uLVqGoj2aWC5ZAirpjPK4y6EkU3tAqgsZGJw4SVZzZPX1sWPjbZ
YGBmDKT1xEk5mBjG6EtSGE1PPQYOAZ9x+doL5Zi63t4QBje6d2MxcuAtmE3n
v9q5vdwNvYGw22JfkoiAyF2FKWZhioT0y3LHyCrH9BYB5ZpIHx0LghNi2jvS
vFLn///Tsb0B0qFQvwnGL9GnUap36mnxoV4MjXA3veXDDFTDF+NAOzV1KAfr
TL72iJAPKUHkB0oU057SltPWlCPpOqU4PCjCvZn6lyqwoR/jMAEdqtrYFHSt
M1iBaUokEntaNzUdwoU9uLC0KGuFZUH8sUJxZATy72rM3ANIvUquf8jGf6+V
lf8oJeQebIC9qgV3bdPmYcTpmRgEINWjgkDNxP8Uzg+P47WZQ1Fu/KzsCUxl
tNQvjKYzPt/G7dG60ITloztAKn83pXYwHvhhRTsUgh/EvEu6vyLsDe0k1OdJ
QNpKCQvnHENT27bEdzK+IONg/dfeKpKLGSJ6MVvDXoWDLCVIEES/h+X1F8fI
07ANG72WSqv0sUYKME5HcIO5lE3kZvJ3/RFVqEkeFpa46UWuIRqV19E0LF39
mFlc4bIgtLee6eycnJl6bJvPuF+80BcTV5vEZtyZMxOHhnOgPYSAP8YzRuo2
s+yT+HN51ywI7WjR06c0tfIVwUkp+a24soP/bUEVnG7uway9PrepeL1aIONj
Mrsb8hy91aIuQr7AaKRKKBSzMYErHN1NSZyCP87mJgAt2IxlDInMJf0pQ8Qv
yi8k4JxCM8oUejP+LdiTi/jtTzRZDTPmUPVt9bnpt4qTNbZPYzoFJFK6ifc7
S4JK8+bCjxrOuw7uexQKxWgxW3HOSMUGh2rCUFF8n62Whnkd5GUYSi5bM40T
X80ekqZ1SIWgtk5/n4iKrRgP8RR9hIr2OM3GK1dntYYPk3f+0BJ15GBnns5q
Br/U7AcrM679eRUHikyNOQvy5CzsHLrhonCshwLjLCbaYKwLRtasiOBVX4Fo
5IN88QUyFJ3IgsGoox7jk60/rbBIshRpx4W5bbOsbfnV6swEGFgXFWDpgbvM
/+C/jcQK461/CpHXBLagKSxTMYEfrjZ26SoW9ffJqpOixneyfpVzL8vZWX7o
mvxgpmWTQ9WMjJwmPyCyeNbF+Asj8vLeY4LpzOzqG5wKuuxg1cndBsndap0/
LNEoPQA7wQ7bY+nk/4hWhGkMUtjPJrho0Mo+5TOxnx1cbdXLbWgWVKBrjRl7
yIwUJJfYjuPOQ54SQBE7g6h7gin9jc8n1TdEqEdk8fqI6qW5JYIHC1rl5nBG
wEI3XXnXYx2k9lJ6yS/d4SxK4rEr9295Y372LsxP9mLqc6346AUhB+0B7Yj5
IkPontEWHXiusXOpfOQN9/q+No//15Cm2IjAOI9OuY8o99uFCxXVLL9AWqmZ
aU88W65lJhx8lu+RSFMgSFRkqk+Bz8MoB6IJQyuf4WCcVRD831EZIsg67wsH
sNTN6Z1Ino8Jd6idTkmeTV/bvvMzBxsbtsMpKKo0TtilXO4vPLt04tcPxzu/
hpxF2chOCTsnE8FvWio1W76DOjZPYMu+KPfNbLMBH2UPufH4ah5Q3nwTKP3/
ttx6JB4xDa36uM7KVtbla96+lbm0KA8984RWkE4ITbvzE1rFLRZkSTqh9Q1G
0mB8/LR8AOt7oCF2Y9+MO01Xdkf0USSR8m///JrxAPiOwsXrCOTSYnvt9+0F
wJ830aPQc0DJCGk9mZIVmtnlyz+jEOVr1fwB1fWmLuqVD1Jg8RDTF096G2Y+
IZCZDWdvHQcJz9kJ7H8I7rzCQgvuoiWZzCuGTMw0qCV/z4BhZU+FaCEnmT+W
yrvZTKj4BRcXuPiocPrQMqSEwzUGyqh6pwk6sD6OUMU/goL58wLQOswmeaEq
g+vlaSdA3toSOOa4HTBnqxDB3rMjAVe81GPJlrYENO9OPewG7qseyZ0r8qjS
Hodh6XEOEz8TRCipqQLo+mIDfJ3uV3RpsGiEMGGb0Dh7h12rUi8uHj8BGRsv
eJZ0li9hgczzCz+6HXpHtbfJWpRwxSKKNRQbbmaz2ogsafvd30feGbUU3e2S
THYSJnnxZ88GlfhHFIWsURG304sihRHZ6Z9x2nCn57zCAO/HfXcO4WN6n7Dp
2NWFoKasTV1XMFyMwfE+/XryHM5jTb0R5/d5J4Hle2qcl2up0uzTGFHHXYCm
qaMwWNEYWgdxl6nHNBmnzwoaEnaGBW2zWcUxUmzfJR04KGNiKjJ6SZZoBVok
z+5bVA4clOp/3fUiseJgechzQLTPd7Qsem8UO6kpCCfMbcIY2rJHNeotlqn7
PvVB9z5hs3fnTepjeS3eU9eB/RM4Ecmh6714cUdPchxEMU72C/k0cleq85e3
Y0BtTf5dA8YI9MiyXf+GS+bDhfUP10EtDbgMJLzco4CqJP6tkW9q3lh/Wp5k
reM7KvxmKnTWbX2i9dxlY+dTnYF356rP2ahzm8b1q7aGlxNBurefOVdtxgcj
qsBQa+b80j6PyOpbXv7cmsmglleUEaAGS+2aoJ+CwLgHcM+xEq7euw95zbXH
eIPVXAUZOxMv+6z6rfwv9A65VLT4HQ1tHXCjo4HHHrvvYR8k3FnpuFIMDm7Y
r59yIuUD1SRS8ltHmB0rCH2kJUATDAMlWIwJBUxVJ4wH+r20HWgH5GxBeVD6
U8f7Lp4dq5MrsHOrv/LZbB9d3w5rPyx1gzvAoZvCSfY6JPG2JMJuYtSe9kHW
HhKgIvQBSXEgvm0tZ7uAgjpvYgNyCV3n1xcbDj0yjWjtYccHEuzh5uAlgc8B
VL/eIU/ZL58r05PNl1Zt/kO6DVLMhHS4aLrwolGvFswgHDdqK0l8oow+uw6u
o7HUe7oiJs63ymsiJk1nv8NQBJxSPXGCQ7MrHDryqBIqQctNcpp7pusRUs9K
fqigNa6/BQlJbWK8xvlv9MIybDHR8XgOZ+cKIvzskG3Rm86GgzphvNW24q/v
q0lE8e7gCJpeR8/UW/DCJisnvXWNzM/v252drpptLrgWIBpgrKeZRze8YfnH
IxrGDjIySU9B4fkS9wh32mcZQ80VzRqQpv5YmcP5a4/90v357AXh1vdK47qC
3ewP93TscKq/oY1Mr6COvQ7E/Y4IitZ8DjyeQHtyy5M42HHXP66WPa66YDoZ
SSBBUWnJozok/eTVL0AjG2BLQ1h+alv086eNf+pBvZF5OPDKKEUb412zwEDi
pfO8LdX4jOJpwggiWyFpQa4OgxiRk3FHcPQunZxqmKMRkKRleQ7cwyUHrWzB
vLyOgRfs4z6AAFSm/MFRzyF2ONJA/wlbS7F/808fmNYn7d4qHU0cbm6Hwrkq
ZEUTcmQ7CpoksPj6arBpuZU+2YKIK0aks9dlbHPaqm0/UDx4k2DlGEbfAzS9
8EuSUD5gokbQDdkN6OeJ7kMnbR2YBGkse6yTwNtsjiRwPSVwSPx+Xx+AC0lr
Skue9Yf5V0UxETJ7or+MDkaluBV5Y2WrG5UhRv5CPX9M4F3iCvzSLDTINu65
rBKuFTEkT+zAdhO9AD4JZJJm5KSOxws00+6HXm41ihddd/VFKVuno+bqDG6h
atKpJcqI3qqTD5TLit2TSou7d+8mFyI23cQCGI0J/0oig2NBa998N+8zQ/V9
hyPSZf3k4Spf8854wz/xUY1fyYnKnxKbnPJfx2vzebHRamhrxumNC09qGYJM
tYypKg/RN6QeOYaoV+CpCAkhdcGZU2sfj9c2RbjScki2Tk1SrZohvQPmlPr0
pyJRG04ne63xeBoZhxkEjGDy0TCE884+i7sOaR/CfY4RT5MQanx9bEEbg4jn
OLpDv7+qnFKFxxgcxVV5sWiF0gUlRBpHqmkysdl73VwzyUZUYYOGkhBPmFVY
Fp9pUC4Egds0kK+5nhj7NeTz3b4G60nmeJHLgHGvh14a+c+NxTTKpG9AyPxN
OzsHunA8Mc7pmtI+8SG/eJMs5Pp/OVcqkZU4NhrkqRZTF6jHutRmH2LLHtk/
cBmmcGGWU1D/UcpSH9PY1cRinny6EydNpZf6LoiMpflSMnDI9TG65H0i/rxa
NQLYqLs8DlZ/gDoaug4267t8K1eVDZUYVld20tdn9srssOVSvZYDuqb/Jqti
4Y79NOnDjhfLjFZwDcZg+YthNCqI27ZzVjTyRQ/+bh62QlWDNXJC1GxXyns/
uxnBxVaOg5t5tl90Pg6ugjPJLDyV4mUt9bYTRtM5e3KoXA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyIekqrE8Qw80EMyhSwP6w0ehvnyisLmrs2Q6RAJkL+mB3qKDuC+Gm6Y/1PeMuOLcyG1t8uPw8IQvn6Gj1+g1wjd2JyRDLXSc5eCYGtTabAxgdKBil9moww9vjuRYn/vtq7opcLTILXEgM7ugsFy0uDwLprxRtZLCM+yr7+qJh+8bH/30d03ABy6VJg55KdOhTDe1sCxMhr0a71utmewwU8OK7uyXQsFhqrqCZ/KsYvvf0tE0rcj9ens8Sf+gCQFIxvFvvBNlZQlbocgl27YvB71RSEk3OH32CvZiM+mjV3SwIumtD1jGqv4fiIjTICBEX72gSgUo6SnAU3iiksumNDRMYlIkVQ8/SUiuHLaTwaTxM33JvhUDdkLtO7ykTSH4t3JsRrtHZNo/C4GVnxGhHV7QK+S5Y6H8O/StvPyaeUfgAX7bdZGTl4LF29teSdhoSrCaAhVXIiQhxBlNbnNb5xu2qxpBQO/f5nYNw87leVkpqfCzUq8gYFXr8cX/hqPDx26ToknhaP2eVPzeFhZSkb2H+P531QhuoA/LR6lDX8kygpQKzFpO6cH18Rhg5aiaO0sbuDNAgfpF4kcbiacIw4Dp881T5jwQGR/iRTC8+QFtd0TGkFHdNCUcNu7kEH3FuLutmhQQ09+UdQ5AE57lN3PsbdSemf2UNkw6l2O8HGGlizM01VhmIgh30ooBRGiIY0u1T8YEOSfTt9hc65u1IDjhVesVR06ob3GpAlOk/07r4+r6D8Isj99mheWQUImwvmEvlIm2HILMLt+yqybgFHc"
`endif