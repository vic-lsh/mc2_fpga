// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UNrJqA/iM6cFIMPsER+ZfzngCzMepzKuUNs4dB6qg9x4Rrvsj1V9xsWI0YGL
S5ZrinLuoaE8cLkYsSVZGphrfexE6MicWwexUT7qR00m3+ULhonXg+FiQWHE
mb8oxCaNuOPhm8Ggr1sTLEoAg+bgNUGmyGDFR8J6bBM5Qp+qTcdzefX47tFv
5mb0vt75SOH46HpuzbVvpt9qWLj2CYUB1ejFABrUVNO0nWUhe/9OQmQR5RUA
7ymT5Ydcn5vBnfW5e6+D3lGQcECcm+lywNli/9xLh7uyz9/AhzSHBidC3YzA
UFSrxOyichiI9VkFHnt7R0zJL5+BBfgdIqqLjmq0Hg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FwKZ8mG75RFYuZEGtw4Iz0InlEe6yYRT1SQBqoT6mA+tIlgnPVDa22CQUxR5
IMoXWnyZQRL34v8/nqAbpNVlrqoRsgNebTdrpmVeD+v88w23VS/hXrmurOKp
IT64Muedpq7msfvBOntyaJBUQu/uerf10R0OYV7uV6QbHVsQICFFLAhWjgKm
ERzTKV39PB137Sxq+BLXQZwLl/0VZ96Zcz+ocWIFy95J5qksJ94SxYTMxDjt
YEh96Y8fVnEeRxG2PPgHaEu4xDf7bZroHl2UnP6Vg5W/IFDW+KbHoOEp2VwZ
l4soq1mlXsfWwD+igr1UfK+dXqKeE1iqBMSShPZrCA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jcs1ryv0pB45xtFliYhuVEtM9Lc8i3kzW/xzR36DbjErLLMw0Is50aB/blF7
yJWNAlI+QO4FqfNo4p+vU6fZSFovgIDefLCP4ueYrML2CJzJfYok4C1kNsXq
5fLg0b0NfWXQeh6epW3P/BUcm2tyDRLQLp2at7MOQBcQQSuq163gjKs6Twq0
DqC28oRnXJSm9it/+5b5RLXcb3OeHDe8dnPb+BpezptSiBKM8Kfaldi894BC
ddvSXUfPYb5u9eI5ZIWRDKEGQyyYYcyhHZOHmOf/Bw4YG9w0nck6o/Gj8QSF
7H0c0ej7l43I3nq2Ql8y9KLoFXgdBEfBssBxVk1Dtg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GsoenAOFBVtqyWvQW5ma4m8avwE5Dqm/d2qEEA9Th0se11nvUzDSG/HxIcoZ
WXE8/ycw5KnNREvby4KEjKCkG2+ou9HBujACobYAh6IdQjOk4h0po/5/hPHH
/6xhs76B5qVSoImZoRdy00rcIUnQCOLUjloaEPEmYVbPg5xHiLYJYa0HZ5Y3
FEBXnPxHptKi6TsZHE+NqLVkXGYcQahtLjttaqB12O4aVlsla7jK31yQXFjY
c9LpIHfTitjESN28PuiyzziwxHnXuj4KBuGtpUvqon7onksTIfK+ub22OAvu
7URANJ3QW1SwjUuD6337o27nDo6hcXnDTcVe+qE8xQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L6YSYhycwiBKDD75PfOzCM4AkY6GNaTSLk/aQBdENT1M3A+VYSg072mAHmxM
14yLE2AxI04vhhWsy7pDMR/Q8lqGyq54XSp3dJcvLKsHDeVqbH3qbZK9wx0r
pgCj44at1TFBvSTxZSUA7dY4l2pSdPKaqQ8O4u/jsDJp7qMXR/Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MnEp0Dg5yEOCgJkwg0Pi+PyjW6JOQag1pn288zWBgfBVuzx2sfbQK82fEiyO
scT0oPm7FWjaZq6AnjyBLDVolNKTrS9V3a42cKDZrLFQX+asnLCRBHiyEyTA
m96vfsRkBXYSKDpd4L8VUc4IgOuTvDhtfnaSjFr6dtA+d0rh6VU05sLmdCP2
wVafdJr6xrEm0EF6BBGGuuTY25u4xdhc2nOu0nR/tjLpsNQEWt+4rAIVH7sY
WaqLQqPSckDLEVzxlErYsM3nqVn7Ck7+xCl6Kpay7aiRJq+ODDAKovOALQJC
rriz5QQ2m5s4eEFKrlSJv8CIzDCP4fgcOz0fWrXuUHw8DtP03qFQ8rnZRSvB
Dli3bwD8EioGC93NNdeeETjAvfiUAUnlPP6fJNkvcIxFZD4NzB4+u/aUd8BX
IsCqQO9cQv8O6OIV9FB90KE58BxN5k8GG6c5lcuZxGptIZKaokgaodxikpgr
MZLTa6UfBiT55Ay9OYgU93mLGHd4DIA4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aSjXvQXPSc+XqlwL1ZC6hbLpCIq/KLPoJtK4PAEHHPjEDmxnJI8raMbl1kaI
5b8dGW1IEwt8jCqN+ELZ2MS6BCqYbjG5ITrMpnOmo9hDuDUDAKzRSL/6in/7
GdqkoPIqi41zlZmSMlpjIX8Su6XaTrQ94wgJRCxAB+61x/Hhb+8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kjCPaqid0PpbeXqfCJZqm614yEHQ6xRg+IYY61P/AHuHfZLQb7dBKjHcauvy
UGxzHT23a/d6FkNb3aMOH0+9nJY8C26uhoueDOHPsfnmzCsUYMCbMskDr3a9
OjYgf9b0OsvVsKdukAzhqZKdqGzkL7E6c0+F7tXEon2eEd6kLmw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1248)
`pragma protect data_block
vk9cBphMEk2bv2bUNm+UWcA/TGDvHmFrMPxwG9FewD/2G9AGNbSPjUSHn95q
YJTUdNyTJ2iBaLHFgfE39nLgCAkGKjFx/jy/3rYQyvxr3jCcDmK7RhhtJ8Qq
0JgGZi3GNbh5au6Eq0g7EcixnwX+hkT8emPc+6pPdVDDzjGekhs+vqZf5ydp
tCrAEtBVisiJCB2oANErqkI/XxvI3/mUHbW2u4aWs5hLjLhlyJfdARMdagmi
J6pra9q+fwO+Gr5UB0oIJpAO2hUzl+g/+5F/3wkaURGmxtELF+XLNhiwkLvM
qZtr43tXDgaNwTPy7qfVk1aOgXJxB3DEg04ipZLhqUvuhojDY8nBMsDxDO69
lVyeNCc8i2imy89JSscrlXdCpDCFkb/euI0UHZEr098W8mvHqycBysO7wxsB
S1fvtxSZ/FV5u9kVaNqI+fYDJ8OTRKh/7cvL3C7Oe21aF1d04OCz0ex1OdDE
4eRXlTsX/ojMyKw3c2temXnBiSA/XjFrc0bW68Qsfrn3A3e2xpHFGx1LyokS
vLXdKVt+iOeaOAt9BBMUNgcf4O/gFuSU+3+NOOo9kl5JHs6NReP/1p61NnQ9
PNjC5YFc3du7HqbwNCbWJJhNnZ4/IRzk/Sw4mTB2heE/ccup2GZLEtuuYMoH
DqX/2lmpTvYYvIX5KEKRm+HTEIMmfHm6BjIPUjNyt0d6e4SUQBvS08DAqilc
l/RkVgW8p/iUdjSKjTb+OLcgSTLT86LAKbD9ZhlUu0+c5AQBUgJK4FoEP13V
6vlHldHLBHd9XJ6aJuMWI3eXcPmP47So6eDce2hgyC/i0fFSyz9EhckRnre3
NZJJFXeZSpNDHeLnAP+rhEIgKXPgHlLfDrom4DVnRpFUkgc8ogRAP8pzIclE
EyKA9tXHM96qr2d07EPDjNHbuJMdj2TLusTWg2El/L/rN5hvCYKh2NzzNKWY
attmi3dh16lnmltWkj0ZQa+1ks7M+tG2TNvtKZphxUXEVNlrmVAPWK7Fqz/N
NqPMGgH0OisQVOXCfYNrcREVGs1nJ/IbZyNbbsek3iZKlnnAeh1B+V4JB631
OvGB6Hs/nu5i9jotX4regNJeqejbFdHtv2kH+7YxVJbnpV2mjNunTye8Ql1W
UNWcj36SnM1Va0g9V+kbBgEdzHgY+nGVNR52eJu5My245asHILhZfUfZRFWW
JPvHDDGIEUsGg+doS0nq3sbRJR5c3ZQBRN5LPOEwJcyabZwnB1P3mvxn/SXv
kMMPHYLVruLJq88ikIKIMYpSfuoj2lpNQYhD2FqvoHAgzr9Z25MzXkdfgpIR
A81Wh6f79GrIUQeSZNn4xeA/yUtVgDv6OfmSy0jNQwBRJIo8dRv5NWQNn30c
aQNuBPRScJ25CUxzx7zaR0SxI+Xy74+d5AOPnMh9auAwpokzusxysGMMKsP2
IwBgGThxcK/zGu623Hxs5r/cZffOxTjaOeMBPLYYwVAZkPr3G+Km4Ui3jsOC
KqJnx9W0NIHTE88lPqWKSkNUhc9za1pToP06QjVJFRHdFAs3wum152KIKZCF
LtMZvb83QB9Gj7DqdfM9FgPCoTucG7/vwVS/CgLfq0atPS+mkPwRO9hhq+kJ
UG0ZHZTMbqzOnuFJ4Dyj3/otY+A2eWqC8ynG7QT3Wqxv

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdttA2J+T9ekTkPySoSvhHoeC2wN3YhiyDbKrky9RS5Cl4EPQ+5/sc5sjqEGMl+ata5YzXfvnB7UxC4OqDRKXRtu3HMHURTNifoP9p7h1SKquQUsX4kulsa48Cig9VXq6vg/tWHlFOOMJPk9Krvg1zdnbWmO+S21eMtI3tbG8+AkRXrMzUTvDLnJ4avCzMVe8f4VqHe1HupnIrr8KANm3QXZRMkGe2Pr6oeNrp+BpBXJwetCGSYT5CPl8A2x/Q3i2szVPIs07w/I8B6jLwF0ZtJn7ucd5Yie57icPWH3zMNp3aC8H+M7PHTH8TcrxuOeXCPOz6mR8gdVNGj4R9QpB/h3frKkb/7sRomMvvh6eAusk6fD3Eoc4wD+uHAxUNE0zUQfMoPU4Kf2bsy3td3bAAQ+cid4UAgkpxkGTtD1v0ltahEt7Nn1G3TdwpkPon9Yo0soxXTB6Y4CYv8iWWOQQvdYQifapac4We6DaJ0PciQv1bA8oBpkwR7z3OqUGFpHM/hXrCyZZmjRp5EunvQkZxBLVamBgB7jZWV078OrnfIBDKQxlV0mS89GS5893QjIXsl5wIUtYmFwJTErk7q56B54jXVPIU/Rfccsu4SP7BkPYCy6va7fvJ4u7J8aE5aJvkLA7fecV6CKL+LcAinn7+5261zXULNKWldj42bhfP3vw+3lRXpiAJ+C+pwan5MMy3y6Uc6cyX7xlQvU21OkBK1/jP9nwm3gdMdA7Z+qdGKxTsuWnnxCJqg2lkWJptDM3OSTNiEyCWnq0bKdEZODrNj"
`endif