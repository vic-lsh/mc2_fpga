// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C9h0Ecmbrj3uFrZZu1hakRekf9/HDJw70i7wNOS0bzvtcgF1oW86Tzx012KV
3pclXORw+418D3ztB33frcidIRjGkN3Dkhzv4Fuvo6UbS6BOQTkbA2Z2QE1r
dGXtkwG3DxaLKBUL5d95MjEPMX6wumlptY8uwviPceZzAHQFSgqOnNs6Dono
dW3nOMMtADI2GFkTSbSYNxsLFTEm5o+328d/3q98Mr2vVX30vJSIMs5VWVin
RhV9bxfTkRrAiidWRqcOo2XDccC5DI+ThTRSfeCXJJyWZ2nnt6NFhJiqX4OL
HW11fYW8nbY6+2O+ZFX9tTDGrprFgzVUQkDSZsp47A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EYRp0BrKWiw8OLt0eRcrgAc9xwzhNv52/yS8EGCkSZvVVopjn3aiPYEJzCWH
fXeurv0pWqFBXrW6lWlAGItrPdcKQwhFO4fs3okr3wpAX0C/gJDfKUs+uQyJ
msXnOp4HXOvr/SCxn7Kv7rMM9FAbOuZ76N4eAyfLVwtxclL2c2bb4ktAiqN/
J2tMF5KuF1Y391F3n8+BAxsPrOPz0LK8CVpDraaaXrLvSu/t7WfckrNl6vxG
J77JX3qEhm8l0mOB+v+Tzo/+wk8XGk4PIAaiVmZ+q8ImslKvEgNJA9tl/Arw
WQliJJyjm2GvC5Fr/2wvLHeSItoYeJFlQc7PgmecnA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f7ns1hRwf8006L4YLPIw6OYxR8lHNSQdVgSMpm9xwfhCK9IO1lRmbOkL67ss
nm9sNqxBg16KdS6jC9mMFl3uJskBTqL88HOZap9N+//QxigVIXEQ56J9aHMK
GqIjikVPxO+lLu2PliTc+R7QUdSDY0D2Cebi86XJEXTPMW8dEslMNsiMTbyY
gvE4NWP6UgxBZk1tlM7atVEKgGEyd9qiMl9sryM14o0jr/+N+Um4nHaJOYxB
9uTjPrwYz+RvrjHInbZUoKUScKGDWLpr7ghKz2o+YSiWEEtd1nf63EQFAQzs
S1ZSHibuPHPNlwginPS7DcFzl7MqrsyoRpZqzqvedQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NMMvIyFZl3qfU1KkvX4GEb8OHbha3QFMo9cCTtUK49DWpY6v5orAym5rb1Ag
elb7uRihpUj5qcHw4c1FrYQOT7JyPZrDWkVDjO+DgN8lMtLL2eOwT9rZJsj2
QmU2Gp1gM6Fd9SYqT8c5p4hcxeA2SVf9R1YK8ob6nFIA+UGiwqPopRdsXaR+
FjpKZEqHMJ43ODhfuALYb9Qi4ICGa6FM5CHhaan4m1lXX3eHTZttC28wweE1
r0Iumo/4ADDJ+fD5rdW0/D3pDKkJzdHATcjIISOTon0y49nmbVQ/gGbas0Vn
df0h5ghVP1RvxcGsprBTwFgVd+w9ywxJJ0IZaaTkyg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n4yrrZ3kxqnG3m9PVOpGLg7ihwq+JUoJ0jAHIkp5Dc6dR3/M0dJTwbOmBMId
MonXLG3rDgdv71JAHhOUZBI6AT84ojAm71O/wNJmM1PWroOSwc7M5v1yisM8
Cdp9ZLf4fzSWOfW/WLIJ7y/4MCwyAqRgD5FCk/2+Di5Ch9MJw+Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HGbCx1eStHNnl0q1oWmuH4rNJbQkc3zZCUXbGR0+Nc2e/xfb0irboYLIgXz4
b8sXmdh8fc/OvkE/svGlaNCzMLp1tEfReT7gTYsLIQWasyBG2EnG1XDFLRa6
CUxMnPCH2kYrXcxcG8UMB5MxqNewL4xUNWNSIlNeMxHHpY79hnZMAercKOVQ
xEW1vWGcRBZwzPYaua3tSSPJFlbBEkSXDqCTXAYFsxRKEXJlhTOBaUqsJrk3
qI2eo9jwpS3zHwtYuzgd6H9bmIMk9ZSvBD39eNYD1eA/ywWvu/QpF0WMI+UA
YdEYilitxcpXgMIoUZXzVQEnzJz4b0ADAKRVewKO33uI3kOL3kQRcWg7MclW
9GmRt0k7hzIW5inyZ0IoglrU9Av4HY2lFFxPIg+FK1qZMw/ugH/An36ks3co
urVlUj2/W+mpVRGaBCnFDTbS6H4ffif9U2pslywYTpsEnR1xQT5QUBQ88FF3
fapSagG9wSAjHmzR5sCZPs1eOJAd3dRK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tLTMmGMxbqOvnuqs9r+zgejrO6+1VYqHpzrLOhxH1XBoJtz2bHZ8zlHIQjhg
ynbCT8BXFLo1B3FYSltcFvgRwhb0qvymoeR4Vv1IG35OQXVE5B1+K7/uxosY
lly35J98ebl8xkUwbYwiWM7zqtZITyj4I62svvgZn8YzC0IKNek=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gVW+3+wxDrz7HBK/eZb6FRKsJcOHRXo4Pf9honxHtnVpMmT1Pv42OGkHwFSA
BjV/Ey+RlFBaXaPU8Q+CpjCRQQeoSL120rn2/gN8MhJEGXuuOmcv7h8oYE2m
/t+xxgRVNJN2Pq/OYPHdxV3uz8vgiLf+XR5En4akZFESCUlRj/M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9856)
`pragma protect data_block
1hAQO3IRS/hfhIv3hnyE6FL4rz78PkP4RfVDdBbT5TxB1cy5G0ffTvBrWn9K
CdSdg5B3XRfSRC4hid6+WQzuU7zfWE6Hfja/FMsBuQGv5fn2/GN19Fc65Sjk
GbKSIygpryPZpw8hdfWBFLvDGA3fMfdg7Uw7JK9/VpK04phPlEprYDYK9V4C
3gvJmdtH1c7rNic/2g7CYbETQoXEEK/6DDTSgKU+eJJYE7dk28Z0eVxard8D
z9ncRUo5uje2tSGR2OFdIKk8KipKylId7+0OiKbtqw+HeTjD/G9AdZjzSmJ+
CQmXY7YOaQoeTmVnaM6M+iOQKdYhpQYf39yQEguzvGcg9HJOtqdTFLAh07Qb
aRVxndYzQ4gUi9I0mjlzuzJKwHoSr4TOaaF9KHMVfB0ZVrOIT8KnGb7MjEsO
/WD8C1bpC+w+ZFE5W3PSpvTKwVAUiuZnv9+0zgeUJAidPf4QFrqMVzoCBZoz
+OW73VY+XX5+81gB0AwaMpE8dQaG/6zFzqadA5NJakgsxWyBaQtEsOWe/Fl6
UxKYrBxqepVac44KeEd2SwlMX4pCVXt5ffv4XWIvT87v7H0FmlKQqAf8H5Hm
kmCwi9pTfJUJKI0zAzg7eVD9ie7FXAyQADf7IFXAv4/apa8pHVabfvhLlcMi
J/dsFxuDATE3e96F54O6xif4j/kVzY8UrKQ9fTO3XTOv92G9mChrSKf5Zwyv
lQsCx5vbWQIRjNZr9JrEyYc2mwn0Eg9n6oYGnl23TPMpepoY+EScqwV2XO76
aIUH5Ef++ORBz39K/EB5RQ+VJ+Hi6T0kr0R80D8tHHRP1qiHTB3KlfSuoJse
671il72ts7Zr2fr3YJByzZw/FySUOStSA3ZOBYcqBxxnxh6oiesxrsCaJviC
9U8vsBR/P30/9gOTsbzuDW6+W0T3uijDY6UfDUtFe6hpEpoAJpZovI6ryUoE
yjTqDo0yNMiZvK6xOHUluILwJKCIjn5wS2u+5cXUNWNURXr63oTu2riU82ix
eQmSvaAcPsCrs62WI7vnJPzKGLZl8JgwWwDchglgY0dxr7f8lt5bzR8SzoXo
Q6tXcS1tsxXI+bcQkhG9mShg+/qK9NVewcIXTfofd1mk5lvoWsizX++S9yfb
OC17cpXBrPVFo5jEnUqYLnviWSIPn6YDx34gtYsNV/+nvatSa2Egd1GwiGpS
dKyVvBY8Y9k7PtKw6FFovM6Kc+GA/n9WtiR2QcYLLvCeIbxJHL7FZE8CVpYw
KR3KDSPOY1qNMllw0yrdhKNMEcPdGLzcDHI54B72pZOzUcDnUTb1yjXzi8n5
msDj7eIrkLzgPXq3yr20+ZVBRPYCKbfFzyqBSODywwBKxAvydub1DeoI/tCX
TNjbjmbviG27wDmBald14Njb5P4GGrG5VxSb68s1FfTcvNVMrqRis41GgPX5
H/bUZYvim50q1TeZc0u3u0gKMZj327nmHzZxXOwTI1Rj8sLyMS+nFh0uoy6r
TGxeYagF1Y5mWvxJ+5y+zP+8GDx1O/flYyloVhnUbCGK966whoqTxu+ZJJNV
auO67Mnv6Yf7Z9rJ7XtVBNlswOKi2cm0S9vfBeLUaL/g+O0X3/T5uwFKOxl2
/YItLeDAfbC6iKKgjlt5mayzeZ+LmDc0MN60eu+sRbwbrO5r1/OT1weBVBoO
ym2DiT0vUBt45H+HYZ9xtxHJGvvM22NdQeLNMgDFQJhxIIaEcoLSK9P/n7PB
XO+OjTs/zLNYBRQngHs9nvgc1k0rAjtv6qnIEdelli+U5FoKrR+J8NgzzYQW
3JYtlJ4WfTgDSjsk1x9w5o+V3O2bEqVe7uYtBzgT5wB8xpRmh9HHhi3ATq7D
y/EQ7eU76s4+WwsCLvXxZ1RU0Gslljg1jITkSu5hZ+VSxU+gRYRtdaX3Zfw+
8WxX8TDX5Xt6n+ONsioHZs5wQ8x8gehFq6zAjUATKtPkBqybJeq3pbwaGLTJ
hHiMDPQN7/m3fX/DkhK3t+fTpLM/jyvkYV2aFKowyrMOPsGq/1ek5FJVCaPh
p5p5yoK06ctM+mLRmxpLDW7EO6z7oq8G6ceWBHrfSPiapmN6hg1+vHoV6STL
VuVe53pMEZJxwcSQ/uSAp8k374u31nHn2tTKyHEtJKPPLTgc3PnlJEIMHTcS
FeoKM7oRm6OsClw766ZaFZ4RV+kYFuSzYwSD6d3eIkI1qLDbI9CTQv43CKmR
X3MN2BkIg/fRAFqu6vrBtX1FcPpK8WjdTtnqdwqif9kMvnwyvbCnG1LFKR+f
CLHHGe9BT2fOof83kVMujbqzrKBeUh/n2p+zjjVwK8TSi6C7HN8eokWEP4X9
6zdJFiYdNs6n2m7nKPFj5GIaej4ip8raHLxlTzMSxlhZcqre8rCDyV31zN9F
mpAZs7FylXcjwMztaA6sd5mwbwubbQAfnTwBzcbkPGYzNBcPxgH0Nh6BZgMl
Mfhrxet0xEoK+eXv5Bxn2fBgSrwssyh6lBp9gIYQDjDSblXmIo/thF0Y3pyU
7NI2lVqpZhJJAfgrekMRRS5GIhIed0iyp/qPpuzYi+OKW+WdtR5NkcN4Sg9P
JQoXSOQH3FTjOW64MJggDMtQQf4G0LP8BCWfDqHz2xsZnrAqqLPLbHyDkOn0
nMu7f9UjuoTVKjWUCqV8iT2F83O3HpDWSqCDlhzfqwlvf4fvUeQQ7sxKcJ/I
41/KaIExYIRQlELyczus3lJ/50U0Ce5Krx413pQQz4Dm9ODZ3PwaXQv0s1we
jVWp/BODTGeCvMNUGK/lnC7AQJ7fL/o8UfhPXbBfxcwWUljYQFn9rN4xHFNb
b8bmCwL0ar2/q2xKydbRk49MUtnK66ak+bV+88HHKOhgxkPrrDUiMTqR4ugf
anU6q7Mlj1vt+VEiM7tJNiKWlSoWLjs8AzCIrdB8/KDW6lAFU2zXu/3BcUF3
FyuSYRnvbnrRkLbMPFpiRYUA1kyfXP6hJ2KpT7X3rlRZs+rwYZRHUlv3yAYR
aixjTxfnO18ESRPbd7jyIMBn0L36FNC3Bnv+8KLZHdcnfiLv2IstUGEKHtbr
RZWOb0JWD5c/gAwaTjzzEfSPLSrrKm23nU3aAup/S8h8YwbpLtf2IxmiAg79
WFkca1VlbJln0lCW6GXxYlTWV66Y7QpfCkwZQVwaRSBZfumxdvurjApAXYnb
ao6G6zuGEN3aRiroUFAr0YgoJjcVozzAyPt4yME8QYBU50RowakLBMaTVo6p
0a7Udlda3VljX8MYnYQWeSDL97BLIBiDzQzjk4ES3ag+wlCuqH+AYnRq83pS
C6jyYc4XRduqHBWr2yaKjwy51+Oes1zI3Q2/7FbDRBGlTiB6B75cmggL0SNb
jmC7GmSFGfXkmfWHypfmN1D5nEDAmySkZlpwX82BYxWN7zLmoIXhJbNn6v0y
A1C0Yk31j4lKmlQGJz7nHivnL+uIRvdXCGu6JEHTwTU8x0G00vT61IDuVA+9
2+70rDZ0wO4wfIHldJvxUgwcz11gVooyuQ7U0SbcL8e9gpNqq4Y8pVO2eM9W
TV3SuX59bhk3evu1H9nrCcVKPumDpqqY3fNB9eJV62TVP/6VhR2/uc28jaxE
1MvCJ8OcX+dFEYkKatIxmZuTvYOAc2vq5ohqGgcTCRytcls1J1gXWj82LPtF
Ii5By6/q0Yx4UEHdIYqCbSuexY7xZF1I+lQUDpI4YOUd0/LN/o4f9LVraAfe
uExo/0y5ThD7bkEijSJOvLvmOCYqOZRg1EG5Xv3QLHyLnY5ZhSDT3qhfcH4p
3afwqTOpU4mWCGbgDtMT/7dbuis3zwfAS2KrwJnhhCWYlIGm2E88gOBkZUhq
XdFzgOPZxhTWrRm0q7ntZqbVgInyx0pBaII4W1VdiuHjmu1rOjEeZgtGpBzM
1wNX38X2pkLyLmHwNRzBPeD0y0/h8PtD+BIl2H4CEkBMuS9aXK4wYx8YpqQa
XielEy+82GWD0dG6IegwuGeTUVgeXCM8SFSjfbtLsw42mh59Gbmj0idiYBUk
152ToxXTUcxtaOc9TbyPZMG0SLaPRm/Dwm48ks8nmX248VmWQ/HQjiARh/oj
PTxiToTWonZdlsMUdbaHYpz6pID+hIY2siFP6EJJn7KYLriaI4w6/mIeU4tc
HW9bvKHGaiuZ7VZh7AEuYo/xRMmpF/jjdPALvtgds8JvZgoatN4xc//JvNyH
g6YavonCjE1gSe78yGPt+6dLd9UCSV+UgPiLMSBCHqRgQbDOM2YAHqFnQ5od
BlryJ7My+ODKpLNVPmk8yc6Wt0Za7UrdLL2Y2337YVtmBv1AUjJQXgfPJBYu
nWgMz73ztqPiGBXT7ySN6Ztlm5TBNmAHOfK3Ycl7ugdhcKyY1jq3g5GkHo7I
LOVqMKkAJoIOpW7jNF6PB/1auXVCYKBdJ5a8B6D5DyrE66pjq7NRK9eUrH2X
/f+CmypzrNCdCS6ATMlCZ6GEdZpEIOPicJ30Wt89mxx+kxKcCc3k88WelXqo
bv8HnDudG9eeGF9YqgM9URWORHUq37s+KcxSz0INRVK0DVnlVe1yj0Hc/H1n
2vMzrEZkDBf0qScBdEwKnk8MFFISSyNeZ3FF6aB36HhMJwdqU84aqk6Z+pcW
Ks8DfoPmA9gk3wlZAZRKJQ61o3YUG6y6fhZDzesCPLHHMdO8mtOr30xEi+ST
MfUyqjCfWRdSikxyo8bsO9tg6PhwElmxVjW8+/KlLmrP01NCTcpiNf1Lk1Cb
mxWtRoye1+pMOt8rT6oPSxxm8QEX3f1Pbqc94yHLxRHjDgGX7XrvEUa6M2tx
23gdExDxTwBzUljsTwAKwlaXh/vt0XzmE/DyNlvoJdRCRV6c0pSiRF9EQrkb
pP8gSw/HBJph6NpBkmCAsBkO20RVAxEH5HxwEfjaDwjf1oGUgPP9RRYR02OO
9We9Ki1Yx9Yxm4z7w9LKc5lNf322B8wEkxWCLIqStVXfzQ4i5B5oFrN9Dyl3
rt/+kf3kO+z+Se1SidvHBmfbYF/mXzZB1ohOJkK3ZLTNyyLDZUxlzCfNz9oi
3uJamzAg+Hzu+0f2LtFGHZ7axPrqbPcnEhX2fvTwnLHTL1xve5JmO7fx2/ZH
ZfX1tY4bbha9umWmt5Ihk3zL2SyGSERo37NFIrzAZqPEHNcoIkTaBJEbae+f
41vd8jnp6l1H22nZ26m9YeaGBGSE9OD0LXDfyYB4Ck2BdVBn4x2tviikqtFs
3O08Ap++3GntffASdkQGg/s5GsiFtQuZV8zhQY0iCIyADFWFghNh0QbOl8/6
bVHrOA696dcqiMI8IxDC6p8TZ2UNCX4r/EIxbjPamklqFlUgjJYbibJFNcVr
1W6OXZcQXiZxSffIzEIZUsd5xcOmd3xAwc5s/suswzYhe3N/xNyHy8C5l/T3
zO84pdXL8EHwLYg+I9MM68Xn7/+QE+cpTYjxPBMpINt6aMdCiVP4I+x73pos
WlFL85QSCveMGzuvBheFpXgJrFtDIA5N99zw0jitKpTEs1N96dmH5a9ZAXjn
tyhZEd+AAp66j53jlQZ30713WaSnsoB25fpVvmn45u1CFvITW+S+DPM1hFQy
zRIjbxz4u8mbUKCo1RCB83lmMOokZ7ujeihF5GALxswFqQlgP7i/nrfVgX2o
zihGKA/+lBX2mSORhyUWbdoUBDsLwFzbSUb8HquGdYTPehMJxJYmwIjtOwp1
winXzdhZfGOefbPXGosqLBqQjl9a9G8LAEtymgoCmDh0/Yy4bW99pTb4ap7A
H5GcqrTY+jLStVbQqcFFxujhCUPz4bhkMYRyWpnhQ5TWxrUlZj8v7wVLnrGc
VDOvSJCHtjfovm2s8lJ4qIDsrydzX9khTjTFNYfsDR6cH2FraPzvd25yWyAx
sDEnpwIxfYXaeoki2qW0eKW8HJDFaNRHugA74TACDI8fyP0g+jzMwh39bNFB
KQAnySz+wxcg/VLAENfSk1anTOsE5GdV/gjuerih0UNmQEUov6O/A/p6kWOJ
jTVIwnDbzI48XKNE82tbe6jM6B5pGF6Oh0s320rre1la42kYE3czHMpjllyw
R9QjR2iMzaWWe6PHyi8qSQdm1Dq9gOE0Jy+D27q+Ls8yL0yaPtnhrUEUxWeL
st6gdKJFgCTbxFvUBpi616LySWSHub0+9eD8tef+4GMSmHNLBLUzIFCvPInK
MkWNQ6AcBHFNZubf4tUFSuLUQjc54KLaWxitR7XVTUl2jO1D12gdleSDjDNG
xrrxDdeuna8+/sBjkc930iuxjNk/SvSmKjXYDI+SMW0H8U3WoBF2TtlV9nxr
s7DfJedDec50PIbKStIM96mH0tahoNfYx6xi4yW1KadQtXriiPGRL9uiSFrc
xc1Ov/RkJrXsGbK5AEPc6BB8oXzLyfXjbuwrMmXcrRRtQzSDaPq6tO9F1Poc
FygGwti/ZqHd/aK8qTliotBDj+xvalex8k88cERjOqTFy6WcZwNYprwIoqoo
AvMetaQiDKTNZhjHoAHnB6fBfYoDYr9nt3lVvZowY1Bp2MRQo6y3GuGYbfhg
g/R2WYLrQuLWnuR0ml6Bhz2NAVhz3ni0R+Kpz9X/BsG7oV/UTiipVW6ZDJIV
VxAZaqixlVSC7zdLTf7Qj75WztJSWQMvtS9BQmDQyOGKQi+zzYrXHaLdJD+X
grtCYz5sqifJil1rJIj5Ww4ff08ZRwpCEDbeRIzYtre4RvlWLH3fq6LM5B45
gtgOvUNO+FtgApg5a/iOhSvqSEX5FyoeesjdAuOw9UZI7Lhj+PrhEt8jq0jm
r7/oQYHjlkF7K+ysOS7gBS7ucgatzm+K4DN4pEmV/akir3TZUJXoLah+36Il
uwpe7LnThYs+U1Mw6Jpks+pqqSv6CPfCMADIfFyFoGofA5ACTpetwPp857p0
xNcPjzLcU2SHxtveludiCNIjLeJffVmZ9coS7acEChIFXkSQEBBwcuI0y9Oq
otMe8crk44QfOgu5pU2AzhcZO107hH8f8bY+nxc+Oozh3Jt9o/LtI5GPez7Y
HUk0EISPZzrKfIQ1Q3NQVMhXeUGGf/yE25TpxNM4DkOvLHusndOZ9IT1BNwB
OpGlFKiiNH2XOWx52Qtm0AWNMimnQc5M6l5cWj9m/Q9H1QWMI7Pz4pAcjLG2
0EQVTkF3PMzAh8NZmQVSFZJynfXUFXEfdIzQY/ihtoLmV7Mz+UfebBZGawEX
OSPf+PGcmPpUTFQeu5rHJwJA1shFB9RA/oKHAElOH36/WHWQRcbh/IwRf1kH
/SrsDduGYiA1vZZfo66uYWw9wKxzhjiA18YoibiVyuI/jD9rCHAiEmucUTLl
hYnFzdR7t2nTyd6M0JHFPq6ic4VmnE++JfVoTlDLnisT1l0hD6VlVAvYmm13
0MGipk7E03BU1SRbNJKF61fLtrfuBnS0aEzhAnYzGdL/5mzljKaPNLA/Hf/t
ZM7IH6ky95xMi2Y6hGbc1oWBrdCHbeuXYwpQK7ZcTi71fAC/7jaWpHYD6gAm
cFPINPNKHnUj/KlBp7fZfe8/gS9JZpEKe9d1u4yMUX9+6eexZybJBrZ7Cj/W
naI4wuZyHPPjweM5Hr/47Y8Uyl2MGxg0xaph+LVWiLQEnuTxK4wXRo6WQCIj
qElOAmk1q1xMtN79fsWOxAEMvsed5iJcLqmfNpMnILS1q5Qz3mJISHXXZAtA
atJIhtEs/bmUOP2Haf+X0nJAifrLzFUQS0fh76PcAwHIcX9OsUYifI35joWr
HL5cf/z4ZKyw9BMXSnt1tfjE+dlBjmKdKiz3MaeHZveywA0YUvgB9Uxqq9qs
MlUypULJ6+Z9ojZ27MH08aCNtCS7yMMQqccBh8TOLR5NNi9ZZZhROKUdd7Zi
kuEmgubrc0xdABL14bG6lO7HxI6qcQfBnpIqmSP/kixYtFy8IwEYEyB3UTvM
WdoSOLovyubTyv0h5GlzYgSyQzPh/3cyxZoPsIYbt0AcN3qkHj577dS0MoDz
1qIERbtAHPqqKiDWnr+I/LoPyu8zGRCYIuV6s5HbAo+VO+hCNkWphEYxJ0eD
v3OuVTg353lCZ0lOQX+NWtWW6X8bzxsPRhOA+ynaP7/GTl5yMczbOejqXUtb
q8ktdKaqBOfVZqyoBJVXqsrP41D2kAYB4S9E01FuykgiY06o/RGFLp2sJbQc
oVLqkpnoBXTTD78Hog6pPjm7tyzPiZJ3v1yancIpl6lqeMGbsQDSGlwZ26TN
OnPQFj7x4xnghUd9YBhPEg92ThFwFvS8u0SrWjQW8+YFdyWckCBjY3uYQzrC
w5PqqsA+c2vB0H+7GMF0biv4ZqSpnuHUadlFyTuUWC+auc3dTpWitobb9yoA
Hj4W2yJNh3IDdbKBYSukof4s5Ip6jZzQnEHwe+n4w38srbQ0hrm1GM3ruxAO
voSyOyLo5O0ohz5iRr64TOiCqNuKuGTxhZy+NGV2pYq6mSnurJ8H0HiyNoTv
NAhYR+qy+haG3f/92MzGxnc02emlX9Z3PYRicu+0e2BuaW5A/NCGE539Sza+
da+rrLRYrT7ys0Gtbor1IouEwnHEX8i5lV2umHof0UNoB5AhldpC5PJykqWM
mYvy4dbDYOJSOx93JW3qNQbY+HmcgLxoXykkPEwbbOhJ0cN0ZFUazdwz+kw4
nA41o/wjIHIc1cO6LBCsCdwO/EIPWJzEt7N5Taeq1YNKtDfVun6+kdMPRuXE
yKWcyXGBQjdiOH9rJj4PTZFMEQ828XEhEJkGbismAcd9sN4bPwqrRMeJXT7t
rHTR0VzwMTF8QuAFKTKuw2w1b2Z99F+IgXUQIUC2vqvNE7CmEMAaDp03ltdb
xBb1V895+fc60EaAMawMVRQMrVF6jXUM4GUbHrVcus6ajeicmbXnosF41z7q
9NujGGfOuwgxjM7TGNYW7Xy91qcfoYmIo0E+VtNchn1IHbYkYOrjMOlb6jNB
yS5p5tNJH7R+dUqcwaTb2DvhCQc9ANOxM5f0N7GcFpQoURaidiGIHk5P8JGu
y1rtQ+Y/MUb2kUA3aLFBURYRg9D80utTrJZdaPxDU01PayxFqsKxWfD3KoKK
AlkkTE1ksWWog2SIcKIubSNwHTxg3OcDoI25eeXjwuCGd7iDiFPQVCpZawm4
w7PU0YEkXJ1kXR1lFySkGipWEvXFm5n+efKHYtacURS2Nf/kL8nYD00QQGJH
XYUPRV7LP4s+1ced4VO+bjnSCoer3Olu6DWUAaph8IH/L6FFLyu6U+CFl2Jy
fkcDXW/Ty+Ify+2pbtubbGVjZKRv5sUroPTOj3E8O8baZEKBfDa13DP8dl+h
lYfwJ7vihweWkKbunA+s+9nZvx20VbxgqECdz1kUh9lQBGfAGg0+fZdRObrR
nnE0FH80iKglZ9vo70/i7O5ghpS0jaNR6iun1iIkjOlrifZNu3t8eD1E+m/p
A6EaAqTa9fUjpegNSQzSp0TuVs3AO0ewF7ablrQPRp/PZR6nxp2dG2MeYi6w
DgS7ZD+9132pxsA/XJSpQO7jPbMBZiHgmxPy14INbzIN6XoS6hFTmoXmCbvD
mMmdTAQkAHzzH8r/0OnA+bTHCq+7ekBDulNWmyBzJQutg0q3xgn5a6+sA/kj
84n7eQhs/maQ35S5ewx535ot2KDyLW59Elvzix87PCSjlRxqLzCwgVo9Cljm
9F25Tla9sfjlRu/OwVQeJLHLk69e7iNMVtznbEfTsO0eprEY6s2dQ+eoD6RQ
70RFz2505L9eVvraGbOp7yaCDbZEgtRNslG7P7/cqjVRVrqRhU/+ZXKbV5cm
bl+bELewckTqCV01nU2afWbkYdxWqGh5PJrzNS38O8GE+mtUejk2SmHNS31q
0+QkkTwLP34ULloIxR+4U7uVwp4LJsF7IpJwHfi70nlZrGWY6cKaXiwk2Pwj
EZjbvRbFMl2PevaSsfIQBA1riqZQ9HWJtTCEHYJskKLyEGiO2O2cqQPKuVpP
8z1w++qn/nmkr1GPeEQf1QhgD+iCetejjhkvxycf/WRq+fQW0A6NxbT2bg2g
VCdvBDQpPBThdHDGJeIjYgzNmVDIaaVwAlzXpvwsIkrjpET5zurJGVS8I1vH
Ar430A27wM5M568zlImen7t/dAyW8GQ83r5vnjp7VW8O/99+C/XVJ+EoVAkF
WckBwf+4q7kFS5JL3EJvaPEQ4KwTdfvxz5C8a1qhSWJDQMTdCMy1kKknpA4Z
T8SwS9u96HW+dUGCF4Y+jYH1MVRDhIt0XY2GAOtDbSefqsff/PiE+8J6Gg3b
7pX8kgR2JIEHtBMWysDIHFDaudhy2XPFY6cXkaX9muCuQaihVjzKmD6gibvl
WhLzl/USTkoU8dt1xTbDv65CPsBQ5cgW4Th3vkmaKoRvxE/uKvmMmryN06DT
UHkpAkISPY/AmPw3Th05aK5PSu4CVupeeycsC4MUgfF14vVs3LA8mU4sp1ev
b4MVaeYT/UKVImzaLVOPndWCdJs2CRYdTOlJ8UZD25VmspQTwcyb4BwwCJ7m
4ihY3Q5szVhtrHA2zaSJpp8oAOFhlZ0oKYNTbZhHk4RGIuxRwbqK5e8P2E/z
2iAOauJd583NhFZOL15Mcne8MLgQdOZYH6B9xgPDHiQF6+Tgf7RV+bAA+vYd
Uv2X3UBbI7Q2aBf0w8TC0Ng1IZ4XqYnufkDzaPxNk5ZFWtyNAX7D165TWnaP
8xGDbAuW38GdwGKeuxeTome4nD6KddiPeElSVeXmOor7gKQ5yFDSqLZfpPWP
U1YC+qFX0//ixwQCZrh1HSvLxrBC7zve+Gu3WR3XhjzHekSlxVxa8VNtV/hq
3bDL6Bjrsa6LtvbeQxd4SlZF/rbzkhaxRsaFWultT9XNpx4aCP81dRGoYUuW
/TuqKPBjw9hOX6wN0AyRO7893nQMkHG5Z3fK2osK2o+XV/q/KtujWfgDKs9C
WyHqzjjOpEf1ClzG0DP/IEPSnzs1rhCXtsCrHpjNEid5naSDxTQMXvUaGakZ
rGb4aE3HnYYFk9axy/t9icfDN9lQJmSMN2VuaO39aUIiJRi7Los6ihQmt2Ay
8yYTyaGEFs9C06eOYMJ2Vlc2+yykAJAiWVS+UDb9ua6IgMkkIHTBjKmUFN+5
YOYx7bK3HEzZpA649oJjvjJI8RePqosLCaLTFzl7BySmlX7aW15gQv9n4Ll/
VZmfjHO5Lw7B9gLvWD1gab7n4dFP6WNB7DcgWSOUneYOXxIJF+VpI/QCpUgO
hA2xF1N7M6cQdkZMC+1Vwemjkr8tU18Gzx5OZWyLhSSx1O3Cwy0QzAcW39kP
O+7ds3pH19V+kUONQmsNGUXXizleXCKwPMhqUTpTXxP9HAVq/Z4mnjWvBn+m
ifVO8QCyiQS3rcEC6e2bJQu5BVq6PCvoIH3t5W9AjCwqgx7GRwtW+MF8Q1dk
lC55e3ia4GuXaUOr/g7SZnBobW+l5XdO2Mz4lDqJVoGgaCvQQHp+v1lXRzw3
mArlw/wR6zgC1pcTSUZ4PTI2+T6yzpiNCDAwVY4JENLucoB+3O1mks/HUTJq
9F00HaRQTK2HsZ12xo+l7IV9luMB1b4EaN/YWFmHIr7fy1UqR3aW4xKnqvBG
336Hl1UTMyC/2Ztg4jnm/8lYt4QM3NZwbMiuWDkStwqz2XMOBoi0HAyv89OF
7gL6YCOb+GjdwvkhdiknAbL4IMx3l7bEV3bIvHxu0FmFcjzE9CoXn+rTs9o2
s/x7hG1w3ctbHONthNFMw8BuWQ9jXhbnCv8JuLekSgHR7n9JBTuw/WX7rv5y
ZOm5om4GDsFYld4Pc8EpKL4ZY8xwxD8mez3hZ7B9m7EuCipZziWUlx9OrzLQ
3FNHly9kikt1ksMj+VC/O+ZruucIRQuNUVyRvCDqztOYGcCiAGBoP2/zHE8B
2adGK4kZhGbUoiATHneuM3sXGxfS1K4pMFeKGn98OnJGHRpUWatCDKSVyi0S
Es4zlnsloCd/qG+S900F8mH9+z7H3YetLqsgE9EGb635eXXm8HpC5hK8vhQv
FTwtvh7/qKiulaFOYVF528L3XvC7Raq6ggE0FRWNE2u9vIvaSWiQT41/yqS4
GZsFnRX3KM+60l8jccmyWz2kRSW2RDVNoxrXdpA4Sw+KT0htW+7h3PZwiuq8
zWo2TvnU8WMp08MZI+ggiVnJ6uurYjQN0m0TjjX4+ZXTz+N73wib4ecg7WNZ
RqIx1Nk6JzX5svseKITtUXEXLuESBEuW3mrV9p33ijq9JccOHhVxklxvBLO9
DwgoV0ntLtDmCYHF0D9sFgtYeQfwFOky8Mi/aSN5ODAzY5OQPux+X1/W0VLK
9N1mfttRogTdVWpUVAE2IFXaANVJoLiP6yFAnGIs9orVQmyxlqtA1rpJbMc9
uWPCnTB946MmZdum4tcxRzroW2jJZowAA8zu2v1zdReap2bPZRG0QcXpKaG2
lHBwvuWeZ6FVaje5Wan3X9+IK+/5SIXD2UYyJ9hj3ZeU2G0oT0U+vd3qOWrA
DysdEcTq782bH4V6GgSG5QSvBtet5wMHzvMeXYjlxiYadaq6rAgVWZlbcyVm
AZ95ICJw2ueUK9QIWc+dAfTigzuGGzpgJ6DlvTMcXeA5pltf+ioTl6s43YS8
TqJ3hj1tKlWmOL+FKXhUutyiPQOPUSlTsKDbeVrixDYEQ/enoSHkqn8rmgtH
fXWPdmhn8YJxCvdbpCGnD7qqfZraLAo0ds2Bwu/agT6p2b6f5/RYR0XTf2Vw
1av9DAqoJ7OjvRVLIsIuAuAbmF1jkIsJSGOY1RtbHM4QIVfFO87jfaYay44j
UmzMW7XCt/z/xtpVD6T1/4l0qXyexFFww7Lb93AOFZSano8a6unFu1Fk/8hG
7ud72ivrKC723cdU1vd2WKL4B2r2X9bVPZ/rMfRpsP9+hFp+Agld/3pONFH+
tOEmqAUjPVbHxhLskDhJYmf8SBgsUxAuKtC6BRYNMkb5zXHByIMVlQYqkFjd
l56TqAk2o8dPDVdNqHkNGH+9ZASinNd3uIgvVJgGB/UgAM2YsDMJAoi3G+Iw
fgUeMDy2klqavdXk44GxJVhqgq1XEJLiIRbZ6m0ja0KhuLYXkS4DxKvb7t3o
ejU6X9fJDc1Rpfly8nXZfHnR++h/9/wWlZkOGM6aV+Badiu6lFAHSpFzbQKn
3w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMMdjtXOQ4SvnupfWiGA4RIWevIPtETZwmV6OLXCg/7b0uLNk3ofTRqIY+fmuBacxWVgQYUPoCR9BkM9mKMJWVEcVwhCm5WSQ4V4Y2UprK95x35GDgeqEa1TuWETVKzKpMTcyOptk1/zEDm8cjSravOaoVjJ2Dy7YSOSTRsPHhXUtvpV5WBqvMoIq5ULzz23WihZSpJ8xlng1XfDlkiu4OzdIK5DtxIz7aT7ab5VUxeCi73a5nz2tYgYsIf5sFj64TmU9ax4WoFAJyCq2UlfSAMsncBjk71WT03uVfIXpTP5AXr9QAotG1yb0LMHDNK7E4MBY864FvKK2Y3hUKNGC8EGDyJmVpMuy+LSiZejPBnEG/s4rf3OaPIDEM3WjCe0f8Jxex8Qth8lJ9c0xSl+DtswaY2DI9q2Yv4fxksTDiXR8xBAjzPq6WYcQbsApJNLyrnvpnvzwl90WGG0oCdF5cbJX5Tb0yNZuXN1T7tPkfridqZG08SUIAx0XFdRvA/P8e1Hsch4hDS8ekru3Vl0Bac0cO7vqB8hZS+ZUs9NFuT8NOKp+2kAZ95INp76eekaXSOakepb3ntjru269vZEKpQbIG8Wh+ynI/3c5GxSB2SMpf3YBlALIhF+jI5FQ5XvDajm/1vYBJRSv6c/yfA1EmOz0NxB1eAgBBQunoh/1FuUs7Nc+dqfWqR1RKJbH/+k3FjRYiYaNhvV1N/xDMpq3xNE7KugSVF7ZNrvz4G0YEw7QxuvJ4CGdxzj9RfRbJCWSTPOd6RBNDdG28kn5GDwYDKJ"
`endif