// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L2e8b2gAmcpT2IpbZsXbxT7yJWqsqO6enb799jXXD8Vte7M0edYO6rAVkheF
SHHvvf1Lt5IyZNGG4EtGTmky5UiV5eRLCoRpILXxkCwI9Zq6yd2i7g8hSMLu
KMX94tDGdreMWJE1XhjXo627eSZVtboT1/BCDjyblehTcB49zgukLXHhIq06
73UZuc1nohPhCDlMYZoXtZT0I1FWt5xL5c5gSoAnimW1NB1Ujxoyj7EqBDSo
GUorRvu2UfE/CA7VFgrRfOiGVcoq3E4Ku3tMZNPL/ZNDJKgBBDrV/ALVn9Mk
MqXCeTVPhoORJVYxTg2kAlpcvsPy6m0CRIIp+JyWtw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZU/D5cU09MdrDiEKfFV1UyQdaqDmM1XXJecehpF/CClwX2/j1oDRlfZzZJts
O05o7LqzBJkcfcqyq1pposTM8DboA4XgM0FwPD0b7lwDuHYox9d//hyIHLbN
m6wlk5pkAR+tcBFdUI07r78HZKp4BhJD2zbx+quc3LyKiaMVmupU31snolMO
BHOXZxqc3rXW5bhXikbElZcIe4avNxUBsZFgvgMORr447yX4T0MjoJiFny0U
8/Zzl3BWilZWLSIDPOZH32QfW9WixqUd9hnOjNPxXZfakqb0uWCGuns+iQhO
ht/3QFoJ1jdTO8kb0T5bv02rbSowhl7ez/X1uufIDg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hh0K5upIoJI6Dx5DsAvPBEcmad9avntNZG2uAGj9mPbfIDcXL4x6ecbThXTm
tFuhat+79/Xd85PPrSMAE5U4CHpi4GnEJj+nvlMbeg/8SwwM47Xn/iqusXtb
siR4crMbPpemRhqx4PDqriQtqSrbHGXzYgWCvKTtKqMmfkJ8veJgLSjmTsCJ
l6YRgpzasbzZaAl4gxl6plc/yrNLBSo8L3jdghRk9+4uqJOzVeYab+VWi/uJ
qJ7S/n7i6n3dPdCORepkbtRrG/KxV0Sk8eBBCJl8VBvRaZNbZbRavugZ84JF
SEF8YrWBBrtSuftb1aRNCRQDZj2kBiIOMG+gBQ9zaw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pZbWxKE4tFFQ4WGgldsWb38PvjeGzTg4SajVrNbsyCEAEgG1Np4YQoAlVW8R
fYgrN1bDrBx3J0UUIVF3Qe83RrW+1Txch46IgKNVU1two+I7/VCOlsS/xfP1
eP1sMnEnazabLwAFxr/r1Uyf7EB/669a1czKTCO65m+r9FL38QEnOvAVYiR+
s4fUHSOTugRJ2NQ2fkVpZs9IPmnXcxDQDA6HQkoV6gYkXv0sBxsI8o0yTm2U
H6UdxiPZkLI2TjQ/De0X6obccsHIzqQIs//+wRsG8somFBijQzvdlNV5Jaip
3bKTfFqOiCqcOBWmmWyew+f/H4KjYGkgcnfPIBfmlA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kqErxvCFem/vg39t8CnS7zGtg7Y+iibXcGYgl12yBhVUxxXW/ZQh4tzSoP3G
IMYGSd0x/K1yBtjpNqqBQwe3VQQYgHaNSOlB0ODpifZs5v61Z7Ajh1/RH7Jv
b2nwksQHnBhIFKeHulp1Z8RAcNCf1sMqo6DwO6coOMAeN2nmfMc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nIDQZrCdzvLfOzLWnK49+AXZTKUfPCZMSf+Jt3g2G1bJu6JxLw6NIWx+GnSX
P/ABWDNLzP9h2KaL7DvSJovvryZb+7MMD4zGePeyUDVC6icF0wN8yKg09JTo
gNyzTFCKbqOxCrrly7X+nQzwDy02mDxQ/OHzJPsd8/iDQ91Dba65wy3lT+J7
nqSbK26sy5tKNxmiSCyLMzrq1wgpi33MmerA9l7+6PkTEBciT+Re0lW8vANA
9i1sw2zbtbeDHhkg0ENHD1jzj6IPCGikg6cwJG6DTf4CqxSaxooW/AkiayRK
bTh7vLnITTyH0pjpXUwgFfwa16GbPaYcdwqhzNQwmgCcmY9zEcrzoJZ9DCiH
D7YuU7ZtD73cBlhyzLpq7HuKvoKxFAJ6AuEZtg+tVLsvMB2dn5JpfloxvgEE
Jdmqwf2hNrKFrDMVRQzEoGne3KVOUipO+bhpJ1tpazW6JCcDw+QAwxdjyA/7
cJCbC8AZhd1VsFRP6T2ICvoyPb0GAJtH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SkIMN1r4FyJ0eonZ8uIzfR5mfHrPIZLcRyXEsSrczpZGnX15/Oiq8Y7xVkqU
zlaupe+j0U7dM+u10WyqOnIBCN6hFLqi1jrzNIyuWkY1smYGYPoxP5DeMKyu
YFKDF+eCELhpfQzRxPbyTrJ2wy6pTOx1aesLPisAqHMwaJz/pxA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NI/bwitxeyj1ozDF8p4tpricxNKGpGXajzkauidxZj1WFWKmCaxpjW5G6KLr
l9b82KZLt3PqSB1jDZ7sirlgCR74JqeW3qjzz4F7f/0FqigK8wpMnxTTpfFH
39MrEUXweF0S6ZvYer+fFnBvfUKtLvapOql8ttNBbqVQXuKjHgA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10128)
`pragma protect data_block
vRAgO7Y4edi59y/xYa+jWWCXW6+w2qZ/69fLcTDTU9ToUkQ4KkggNVJcAu9F
+ladvLVGWaSVR7dePduMKTJZLmMJP8CFmt2cZteSM4NF+cKg48v4YMzkd5km
+osgUu+d5eSKdfT0d1R3I4K/sUynmMrwhpYyutfWSsf/MuRwbivMNHUzV7d5
jo7ErAJ84JFXN0ewpUHxSpEzStFHQfvPtTh5+ZWPjBL1C50U7nJKmJQZAGhv
biUf/SevN+wX5d7sLqtUs6a5jew7qS5q9A3XltzsKg68XjA5pzkDGfxmNVer
Uj3Jx9xtc0se72oSf8UIW6z8C3I/KXrHQXxRRFpSrMhN4y36n5vi+TJJjYxC
JzpkTSJFlOjeQc070cDFC1cvgkvnrTIGIpAVS8blZ3O90CNdf8yV+/Fu4i/4
hlTFvE5e9nfr4KS1170TAX/Yy84oUTWZ8AWuBmn86nxbqeU7Z0Zg/xOGqh+e
nbV7KRtQUPacHCZQ+S9uFdwgpnpZl9rT0/w4daDnA1PGslMWlFU/7J9vHVpo
JhLtUjlUBKlvLOsx85nZxP70NvlyLfN1IGxJlFv0mFFBZUKPDVTOrpIN1TPH
Z+MxTg68WX074iNYEaOjUXij/bRHZ04x9jUr8jnadAluILc/JSdZeNh+rK2k
aRYvJHvJW3Hmv6d+Gh9SP+FhsCUM222LoCwoBxqItVp3SfUnI7N5X5uYReiO
KuwTO/Dww9z5H7jEgavdtssXu1W00rOkSBuPnV1RpW/NjbUYvyakFYubvVWM
jLw4hXeoYz72BSxR2RF+EEQS+IaDt3bTakjluRmcUJpfAf6gaRn4ZnRmd8VB
DVcqzsf2MM5PTXciSR6gnurpULkQMtYIEDETUwABD7402NZDzYmZtKJIzvTe
6+ybzKD7rzgvY96mROWl9LLnNt/PIIk7EOVEqJmmBpiQvWW22BiAJfZAB90u
vg201tnBP8dFSo2NL7lpxZRmtU3DOpGkIZKnwn+xTo55rB9XFD/5S2CsTtPc
j/rjoyPmQZFRT9RrkmJcJ5m7RQMY5az2ftHI9Y0f/Q791n494XNuxl+F1wgG
+RegDZNVCQu5MekpqeZNXFtoCQPbMMMessD9i/1VWlT10gtF4lJO6dw/Gev+
C+bughwhXJTwl2UbultxhroDVJyhXDYH8u7OuaT24bQLPih/RGlThpHiA1Pj
/VGYoE7V+HHUDzlh6YMLs1YV5LOe2y4Ss8AHfehWeEF5ufqtGAfmVEhzALvw
CXcJ5qV8FsVaG1fb+nCQLAtqQ6dHaHOFqmVBtdjYhsg1wcwUScBTw4w/uZXF
fWdqz4PmS+8qLn7P6BSc52Zb/BYyt7qZPj+CL2zhC/TNGO6gMU1YWi1/+Uh3
oFnKOt72bCR6z6BwBioBVgNjn3PDNeBIlWuHqPiMQfVoHqDTdvTLekMlO3WX
tHajpEyL3KBjcaSomr9Og+MGbtjZdR7mpQ1f6RJu/qptWufo/zWUf6+7LsDt
HlDU3bxxTCO7D4h/5Bj1UaX5Zlyyg7fLjkuZ/n1KxcNwv+IQtKT+vZCFxKQt
bBDbLP1SLkW7t8VX9Q1tUF+p9gxVkS0Nf6tBFPw1DEy52IMsEn2439aZSIVb
bhQdp0UlexUxvx4/NRx4ZSePbO0CmxbOFrvP76aZLjGAJD5nKPRtFVNOzPwS
avNkJYeSWp245ZQTJClBTzFP+tQciOt0jlUkrnLdBiUBtE+KmWD/VEd/08Mo
pc0YkKQsJxaAB6uigIzeZbRe/CgB6WbhW+U50812jcn5mNQNnEZg8RHRs8Kg
ORW3HQiwI8Pk2TAo9DzbsNW5+w9VLWTun06qzjoCKMPwR3cMSN4Z72AhbJHC
+0WLCo0BxgghoOHAd3nZyuuyUbS7Ic01TshKJIBMr578tdieOBCvkWVkVdiT
KlIkshgDpwGimoCsdBgXmuY0WN4p/0kX1L4EhJau2evWW9WFIhUQy/unhGaY
GwDzLASJbxHgHeg0C3Bx4A1k6dKcl3JdkDIz+A8kGTx6cSDu45zts0EmbnIW
dgQf86wKh1GZ7SJR+X4chwafPj/2owQNPZ4+WQrXhHvBfAKx8KF9pov0a+Rr
NvoSnBoKc76r2GcNHXXNnTh/EJYYLFwIFChfMBhbnPVV1sM0IhXfeZawo8X6
N3ibjMtzRItbS+GGLWXxIdMBO531HI/X0+XeGHiDX2sMKswlxlUppx2MsHff
72oBcbc4ezH3Lr/XG68u0dX5/KEp/06F6J22U5H9//Ow0QscBXGY9k7V+LTg
A4ntNGnze4XRhRYuPw40do7a6OfPREJqx2KeT19R3igk8qODGCdzMzUSml3w
kFniDtCf3ZKtR/zyMxEv91/SBNsGNM3IF/12gee3+86yXyXlVbA/9RWoBdPv
MglHyAfqeWPMFq4DXb3blA3bzHbRqBCekV3yYrc9xwdrJYBr56QFMJuNj7SU
8zHuUeWVqPjGmTmemcv0NVPywnURc7HXQu4aVsFV7Q/GnqKeQJGoAAWwD5od
YHRfBO+7Z25W4JSD94zbTZE0dGFBLc2PPnKPt7bNzzw+2qHOjyUKxsQsJxLS
7qYxPb3y4qbhHp0X2gq2zcNBsIm4ZrzTzR3Zxn81Vy2MB+6m+ENWpL3hLPyy
gRMH4rWhDBlb8P423roBDnbvUmSIABte5h9yKIYz9dVS8R9VAgf7OeO8aRCG
EGNTm5cSmnm+BkJuQZJexMdH/vRffU1HQV7S8bUkeb12/PeimXKQaeIvsllr
tbMB8444EjB+hSGNpN7dnp8jz9P9TQW9e6s2lcp8HH3S+np85Wpr4mV9eDah
nELOgw5vcIGHLQsHcJ0gQUpFnzHM+K25T83UU4hbPKofENATnjC2QMA9JfpA
haynAoCdxpKUoqqFXlCaeqAyPd5t5brAAvP+y/4UWTNZarsxhuLzV3ZHLLfu
5UazQEh/8s0DmgNfxCtDSwSzZr/4ob51mVB6nfIpyhusadpoqxrObgcwRO5h
zj5+5F7F+mTLERoEIv3+KwYhJILIVW1epDiC0u29zMtXBaaBpr5yzj+o9nO+
HDJyZ6FFGoW5HsORqN17+sNvdymlwekJtPzrV9vgGMGP0i4oNrd7AZujPVKd
GdkuXnQVaTVNuncNGNQYVl+sd04PKbp9aKBiAqFgqDOVYeNd++XkUZrgQdHz
6vosu2GMBvkWjHtSRi287xFBhFs5BoL6/4hCIWySOIsNMhTQvxb14qBKpSLL
yhdjlqQ8IYhEE0uCSSxBHHAXbRMr9qFxsfULeGjdDwJ5rskbAelLO7D/o+OC
4PPk4vx77BetTbitRaOntkUG5i1ZgtXqIm7H6WAI/tNoJ1C9R0AmWMneJXfg
PPQ2u/ra9K80rd+XcFDQrl6H5Q5hsTRvXzO67i8+VHHStDXOoaaS3sermDyc
md30REoBvgqc/ge8BCwFgsh/PkcjudtX/fLahM1F67KXw5DSCCZNBCLTnkWF
FkncGGyO3Su00/5H8zMpE2/8WCvgvbZg0P9m1OYmpb6PI1s8z4R57dtCztkY
/2Hn5d/oOAWDyFxekx77d/kgojOTFyUegJ6pqXlZ5PE6XjgnUwwsxXFvSu46
dEZKa4Xa0DvjNyo37BykoWagHs9g2ZyBTaHGVKt8FqbpEYhqlvdmCzVJwYXS
+nd7XivJ29kj3cWOFX1bKyqqIbFxYYTZZzanbkNCfYwUCVPCap21IE2h1knx
s1h50rjCtdgjmFiA6nHexDclVDKB2mQEtixEHcNASY/AQPHtK+GAeCVdLb8m
EjGzyUROsyFqXd3ptiJ2X9XLxCaGH2FWnyP3TKwCJSa6ec9nCNrct2DT3RiT
+G/ILveesrCXRZ10t2ywNJ1QxSaTG2w94zozYINaEowPj8+49U4uACs/7gEp
23rYweGr0whTJ8fKGu1nXaWjaqloutC4R01YZqWcukEhl1U0QeGuXctcaG8S
hpOgbcMQ3C6vNiexikQ4mNdzS5qBhRXTPu4tDVEAIr1LpuRI2KMURXpnj5N1
X3EmwFJKj22tEfe8SgVZ3n44WbaWAZDb/ZyCq6n2c6BWHxbq8UhxVfH6tpt5
Wlw06xAocgBWjzRbH4AIhQnMbYlXTauGtTceQc75kM98iC17QCTVFxibAKor
/BVF7D94enNTnXAXQLZkWhz6iFVkmmibG5ZB1Gmoe0vs6gZr40w/cVoO47//
Bzw+e4b58Ftka2B+Sl841+deBNy9qdLGfE0SiqAaCV5kXXU93soUbloKIPpB
ytQgSUIe/uOu2jUYRzDkOkSmBF4Gc+AT2nQlen1Ug1R0HnqTzndsYOplraXa
IcOh4u6e2PKfKuh5yVDOr/dK7RjV2OC9MZyZV13Q5XVhY/d3O6OFVKa1eUKL
XIsyIvhqjwitF+Zdby4H061+GU55cIVYOm1K7ah210MIwYGKe76446AfDCki
d6un+1WtK3XOvXJJtfGfnV38d4z9wtx4wQy3cQ8Lq0G9GGRl/vEhNK0iEZ5s
zuyyod4rlssHvgLyrOq9iN1RiNz7PDB9cDPG7LqkeqeGoWS1mbchjg+c264e
Chq0rlvUUWj00eZmKc9jEiSJsK0v2Yraee7TLOrznvkj9GRPZS8mvsFGVWYU
w57cvGnGqzgmCdqF8I/0WpQL3qXehRdcGkciZCagMyevlHtu7w7CsW3lP1F1
B0DhRe3IJ59J1jrAKU3YXSOD/uRTSCiD5jWHcQNJDaAi6EW8kAKEKg8XetqC
nW1pGrfBNspdB4+BUKSF9H4xu6pWqeDgrVJvw2129gzSpPSTgnchjvLoLcUr
fKvVDQuRhTEo8+0m561fkUcplv9xxrNVa2jsIkI94C7s75yct4zCHezG8Xuy
V6dQwDXnrJEua9T6/2nXAXRZhK85fDiyHhxvli4Ezf/906ZRHGescPZuXbTZ
YdsjQJ3ryzahPZMNQEAoZfaTeMkRlRqNleEFeQukdllH8qNshF95EQjLIHAv
bZg/178E/L4OjLm/1yf35+Mvfhp62jz/2VLFgV+0bEgAKEbrALqKhYY+tjCK
81VfFkmNDpNX4xLglupGVhrPnbep/9ToBYYG6FGd2WjgRq5EWnYPluRCetEv
abrlb/mF8dHj8wkAO9Q091aYv0fpydzWO0kqMkqqMNSX78iHH8ceFyx3QySl
BCBMmZ/3z9AhGAtWyXER9fG7crHOQW4QVvW9V/0W9EU6jdeQ+dDCSOwvuyz/
N1kq5F0KR9pER8tiPhIgwhZ+PHiCCoXP8elENzorKuR5K4TaFbqArR+gJlfH
rFNjqsbwnK0a1LXl9HA4ypIJAvMuxa5egbTLlhX0xNwCcMs3hpKTT8HRLR4P
HY8yxaNtVo7Nt+kllBQKR/cd2zqcppgYE397P4F4LFTM7JdzUTIT/MH/gVL3
4+nppuzfD3XGt0jKoo4Lam8lFQ/tvVoFSR0B4BbrBgMp3sSRb3zqljEoFdFD
5hu9RX9jeoLLV9maKCBtV+GM95ziir/z7Y/hd/pCVNhFtyiIKSwZhXJlWSWX
ro8Bn2wVJuoT9stcSXKgRGhuXremuVvnazshttxHXMtVSZgLUCwggjFJZ5yX
w9TQwE7gNfrCWttPglcp13hMKcZlgAALldcOMlFgBva3d5/CKfUIm9MHgPm+
46MTtD6ipAGYQfrv1yHsEZyYKSLRT80LL27P1rdDybOomXqIW9O29Ukr0aHr
BfwHaTSKy7q8nazZT14Z2NJ6PdXyQ1hGVQZm4XHKoYT3VtFZJ+NFMKor/ovA
o74ReHjrWyt3drVPa2FskZxG0YTT13Wo+wxfLEKwS1KGJjltjmro3GMTo9Av
KSnqjVe6H3fmfyRvCTIrD0wcVvyLWdRz+m3XOVMIJsXtLpGYsApFX36XrPsr
o4zF/LneMhVs0hHr3tr3GtHxXGQhU+sdPdVgsJPlzHKXwJcHHVZ8Q6mXXUAO
p+YfqlIogrNJ3rgmnF+i+vJyWhjBSk135Zpbul2Z1xPD2rC+pGWQoY/PY2Xi
5Lsq49asaX/yXcKDYac6dnwzOOE3IgVkhbLwG3dFuoAHTmvCfgvPwdDqtSx7
9l1ZXperu7RewxWHfIoSBlT4SZMbgem6VvjY/MDEm6wYxC9GCUNuMHbkviBH
ZOjyOlVESaNF6jywl68qhe4jbyj+ubmI0u5FBnLsWGInDCs2giv5qTAAP9o0
GQovKSFGIYygSefEnXomyheQxLOeR/6NpIaIEoXGC/h4h3GnXEU7BMVO4B/C
iHCwPFOKexX23rP5TQ2YCHd30G05k2yzXsCEq/i7QbEla57wCHvdM1oHCBtl
1TpnMAYi2BvDHKBpZadpO8PXnOYqC166Qlz/icsXXHT1acGyqfcvk484AdXm
oIse9mJC0jlgyCcecI5KQOdKtWd/ABBl2nPJBGb1mOMQEBkXqliXxv5CVI/x
37+DRe+ninpbO1gt07SY8aazKQnvEkibyLJ76LClP/C56u3CLumhiwterJ3p
eXno+RMZCJPERveHlTYXmB+oCOu/RbrMSjkoJOtSyZLk1wumyChZOgn/BsJJ
e+hWLHDapsbz1/7L02lF04VWAe3zmUDk9dzdsBEf0jblRe1Wr95BShV+Y1Z9
WGL7TzBSmlYlN3bJnKLHHgS8SZ3bazbdFM6jp6NRIUYGPlznpwEerz9mE1Y0
tP1UNuumOmkljrhZR51Ph/Pl4IwCigg8lsdP0e/xlvHFT92TzDik9tG1TpmR
aOzgRp5jSE6hSYyfGzvuyJSZBhFXPWg+2Fvts0oxoMMgrQnLNSOXzPNOCPfH
x/YGw5xMxN9AOBKkxDZBfkzfqduBZSBSIzLN4CWFNW7HfrWhuFR7aGJjbLQg
N/FSULVYNh49ExxeVwVOin3EUsfik7yAi77Xr36MAQWUgPaASquREUUExmpQ
mde4GpUcPfKRdPwvZ9YseeYoaEg8b5UnsbELO2F+H/nGb8KxyDD/lWvWg+zW
WdBMHB3q23YU6z6tFM43V6O3FIlTdUpgK8u240QcSuZfuPartkiHRETBLF59
ru8dDdOmi9CuCcJ0gJLTTton0CxL48ygZefzDsGuMuwnfAA/1vkHjjrcrjlu
GM6WLcHiGiaOsr21NFqxKU2uTKS7EkmFQTbt3BCyGS5sspiaIKMWDTGRr2z/
0wNrvf6hHXBpT4RMaUYVfaQ6ehHPgn/ZwgDOxmtnmsyyjXpVnLuozEZzoZxX
ZVu304PzrGuYJ1/M49gR66tP4Ai7yxa1e+v+marhWFgpCmsSPipP/Uu3JUOA
In6JYP1dHZ9ngYM1uXjTJwetjlG8B/gvbNu7wBJXs4fzJ1WoJK8Drx5QlpqR
Leys6m03+FORbDBuqOHxwA6bspolqYwjz6jZxJeGWAym3P1AK4FfxAJd7+lM
WqrLM3obSO53+HJ9kvN2wB5hdoZZnyHELD5D/sMwChBWL4q5Z84S3F+gK5K1
qHOGoVKSPwoIDlIHwTpQtKNTKcDpmh4C4O0G/LDYgYuQlasuR57GWCRZbPKW
NpoRpDlLD6wMas74Rng14u4B1QEy+sYkOr+VtNnh62F1W49qyUKrkUWKjVRU
zU7zjQQ5ULvscnOv/HzipxUJtkjOVG6r8HPZp3dqiHP26xlmJIFg8b/fCcoP
tJRqRO2Z6sM9h1sCwsKLmomz16ce3zKxE75v9QubHoZPYxFfxYP7ieezXEnE
xua6mV/mdLMoBglYsQ8Ii/vlmdHbcrfQZUlO8QojbU1tjTWrwnWphGy8EwY9
RfW/5pAJjMlt9i9lPKCJW358qErNPBc+dEqx1P/vK7SWDZAlpHS+33GJfY+T
P9AzcPYb9ZTPDjVxLVULaL7YKefbgCXvnGLqTam6AmO4haAWErSp7zKEwltr
uMeTg+R/6NfmOfgD/VRVxMp/pzUTacOkHC0ZXy4ue6bsRa+aYZrR9cHHOrA+
RV2fyl245XWtO++KLBc/KzSy+XCyn0wH/uG+q2XfGZ2PGAsWE3cn2I1AvBtc
vHMBVZPJ8Az20JAdg1xOGyquBKwQr3qrHmWoeyJnRktLfaG1UCK+y0smTWqJ
JaB6IULcTsk/nu91bLOCwuL75XwT+XEi++LAvCgIUKsq76Re10Ow7ldclObw
LVAjjat8fZcAMhUsP63fP0onINwpzSNb9fg4OnO70pkiEjtHwbiiDeIJxyoq
Pw9py2NYaLX6d8Uwpzkaq7CYewy5YRHdbkuA8M7+5zE7dAslh5unlJtZRV9X
if8xtclAb+x7J+N8IkfoY536ElrV+UEwBR9T8a6+mu0+Y6pg8Id7QvVCiezt
YfelFpTg3nU51pX3J0Ej41KCj2q75BWwH2BuI2Ln8p0k7EeNqk/PJlalFxPU
PFS86N8mlduScyKJTeNZw/3qTtiSaPIo5A6zCzNnyo2Bpz3Gix3dNuKXN/W6
7EQZaBupZIAevTWmpdJP/mvYP/ib5P1RfPmCRyX7WqfJGVMbfs2BiYyDXIe/
TbWO+enTkfbK5xGFB+e02JnG/sjbsq0OqPndy22dCEBx2qqDV73+ayx0Qv3Y
flAhdE6DMV1kOLjtkBxdkfE5aKOiISz0/33Mf/XdZpauHIgv3ei0cGr9MTXx
Fmo9/u5EdUTrXW8+D0OGGFdjxF0YCMOJq0o22v30Wkc691zz9916/nOoe6Yx
e5+SE/rrmXeQwZlt/8gyg+psNcsEEVPaNo5gphmi8a1UUyfIOsR1NP1vItkw
taM8eucRwykA54NfjftiOJI/Y45ceY2pWdEGNs/V5iec7YwQUNpUsDRoO/BM
TPRVXiJJN36oNXP1WsoQNExyFyaORenRWVXFGH6/jWdPEklld4egZv/cQStB
TfR1WFoZeIEdSZygSkBBYust5uRURXzVOsLtLtBDZ4pq9G1BhzJ5vCnduHdm
JqqHkQWDx+Ymobztz3LqaLJzMBQMc5XRoh/nNSqt2yj56/LTZCC5QN8Le6/L
wgvGxInrtJdpaZzI0qpqKEvGW0MmihJw52oeIkfFaego8Fzj4oDjjAD3ySUX
lXRUxWFx5o4uBAicuVhEeOB7D4Z91rhxluQnLh78wL3PTltOVhSncSAr/cFs
kPd4b3EwlP2IjkBRHGoLxQfYn23nxywx5roUDqs40Z8fhpqnVx2Qg6GqKYVU
D0U8MoIKFFi0idlzNQntOKS8ZQrKW6ZBvGSgGCYyQx3bx7EQjOLmBWISQchI
1aZwBzKJ9eyKZtwVNzOEmCzJhMGxFu07z2z5IFaFzJ5JLYxiuprBDkapRiSU
4WTNJkDcbNGaVaUOMI9+7a9c49r9Nt+iRiHBu1TF4yoPt3HzePiicSBaCGtN
dUU/KmhA5+7xqWOPXWVcQRt/l4LvhvQNIJp40G07xBYYwyde73puxKuEKuwR
YrG0pnfVqphlwxW9128mSB5Cc+5EE4qCSNftWn6C5D5ACxLs8Xy/o8Rrdwl2
iL0Qc2au8VY3XccshHXK8fHGP9r8ryKKjte6ysnFHrrKvfSqK+5TNMHWM5/4
CwNU9pV3IPorVVlN0WmPlh11cyzEZV3URMYA/OxDcXgz/p9T6fd2BQWwF/8A
mYf4K0m4bCBI2160t8b4wxVOcqphFRJmtszSgAUhd/Lb88vHdfa6qrz3YsLi
al7Y/8fpdNzamVDKqmZyDiLG/TK9mgDKAmQT1nyHbOPW2RSrTWnpn71RNi+g
ZgI2VIOeHsAIwqXY1eawR9vvbGJmfYwLc5ZlHUcJzmfmRg1jdJ0KR2Xf4wbQ
/x84PVc8WUADIs++HHQ/WQVJPNUoJMr+tcgfavJ7ZvGCiHzqBaGQ+4wHmhRI
hlWJF8QjmMyKWlIgWXQRg9ROIKLV8UI7hhNZhTpJc0fHcJFZaANyVBptdGcM
J2RPaEGWHwmMOq7e/b5YrggJ3UqPSnOwz1kncAeDcYVJDe8Qd4paVkFc7oz2
IGAD01hBAry+htdfLWEXT0zDRTKpOtKKybDRB4lDEu/ZOXzrbAW7SQwOv4/1
D13r6ZJM+mckZj8SIpK1F3V6+KVJLJ9vmXIDvAug3pHXLcgWBle4Q8HkLSLV
3AF0MCDO3FulU1sufsH3ii/cNbmVWkaGo97oo90Tbr8yoUqdxcaGTHdxkLEd
iCoTNYywtKWeUrOdc7idVCYjkKsBIbfNEpE4HDG3t1YT3H8eOJyYWWr1Uc6J
QbJ1iOKOZKPGtTijRqH6D1kVJIfuCcdLfYYFKTqEp6CdzZopDrTWMlG7IkNR
drVovXJQ+tdrKM/GjMHPNL0lNNPW7W5bfVyGvpz9rFsyqVexZqvregjnDS6J
/jiFGPrqcNlQ3K6JV5B7vcYztFW8L8Xk6y6VtSGWApoAfaSjf5IUvWA1sCnK
8jLLKXIj6az3gMijg+X0spIfDjoAfqXVo6nmQgbXKLtprnR5D+badO+VBU34
Z6IbNPgC2ggJFp3JHjr6deU/bwXSUuiiwGIB5OYSMpQ/11AcgDO6eSZpcmd4
F3UrGEvim1SvmsmDu9QLdI2wrKD34XRrrcCFFRN2TLGckHnBzTf4IqbrZ2Bv
anSwutLvCFcJWHRi3Svgx98CZMrhp8CZJ74urIeFiVg/YbITdhoJSOfACGxD
GVE+hy1/47MAMHlOJDEeV8tUH9NfNwz0UNKZ5g7xQT27ckSckxoMYWHHFlma
tDvDpQJnQhj2P6A8BXKJe94KPMv/ZJcdrYIPSs5p+YMgGaxmAeTckdIO+GL+
2rDGyZ4W/S/vt4z/xnJSGPi4XacJygp1xiu9G0gUnXny7qn7L3qF/GZ2b7Q+
McgExttbsR7r3vrZ7d9BYCcPUSLgYL9lf3Fyh0qEh41ekbIjQAybiWTh+dQv
x6AWDE99HIenZzojA/V9OCYSHQYe1RV01tMFfsXqRQwu23YvpKlZQ8QZGEq2
ULWJYC/w6xl9c6goqfiQIF+J9+VNkakrVFr1s2A4kEdwTyp5hKlBPQ/ugwoy
aerRvn41BNTI99F3ysl5CRzgl6viYqj4z7+CJ3GMGA/IOOxwV1VM+LOf7aE+
PGzeUuyP3pLWZcNBrsggY+g6W9uafGhU7lwmlLSuKcfNM0vvk88JrRr/5rEx
bCBUYZTrhSpgkjXD2voscBcyQSFrt9plXf5UeNqfC021dy0zHC5/Xr5PHo3v
ZqOOSueq7tRJLGbVYwU/neo4PpJkfT2b77GZ9jM7aFCBo0ZzLKVE4WJf+u4h
FB8Ckq4KFo/DkE7ZBZvnOrOOxhjRAC8Q9OiHGYpunjPW1o4m46vbvT+4lJ2B
jLHjX/OjB9OZQgAva2/8waO0/0lL/SdnAYggFy/xc+r4XtSzVMJv/wMlj77R
Fst5sVncJ7dSdtH94HDNowKi5WoqcUz0lAhlazk+YaSxCuLQ0MscohLQqmvD
YQO/mSaYs2c+9fHfTg1XaKfq7bFrZMtH5IqQhOLS+KBd/nQC98ypJlFfiA40
HEAcG1uirsvspmTzigQNqV2KRk6ZeNpf41fWFM63L8jrJmMM97esMuOw7GmE
9jtBJMQtq8Lx9X8A6g4oPupngMaPDJl2Q4Q1LqH47u6jRCstS5Y0UiA/OuCZ
s//Cn+NFOLLCUKw7KbyGHew1hpR1nu4gdIhU6QeGpP4bAuP4OcXHg8+E7sU3
/BQiXClsEYs7Ukr4yiRr3YS2QoxzACnOdj/3GZmIylBLqS9lnNeY3rdjKpPG
vpnsusMROD1jl/opL6tzyyv+9fUqZXWnZ+fUKhDaC4BYmeB29BiIYxakEHkz
DXRT5kZ3IQnhvMEj1VoUK9NcHtJFfUWO3XFgI7CfPlXN86FKi4mhd5XZlH9Q
3tjeFSDY3KNS5gWYJNv4HV7crf0zfI/qN9UCVKGBSkooOmEWT1YQQQG1Z7lt
qQyWH1TmnAdf5r0JOyg3Lmz55hk/1rGHkH/Cg7R3lbGcVhisxwkKyiSnKiZP
SbFRWapgiUXrAwsqWdiJU+3BLkHLaIXmAdZj5Dk8rlnNlphmbN4iLpPnuQ8J
i9/3j32+C6yfnqweeGof4+wOJWtVCmY8EFBuJlAzqIhrDpxHHVFcvGuzginj
lQjJAYvd0MWu6z7QsoZ5VdaylySSM1gB2ebYCJIYI7kLEJuZiUJLHn0e+bYN
4J0EsJDzio5kzEfUDoxnmLDyJJe1riBUEaDbEWwLDo6g3PTf9h1smIlV8wSE
AmMITjwRerHsB/nzANsRe94jqXMVlu9BFP49XQZ8GVvF/TEopZU3J8i9QFFv
2mW4FfoBz/56lsX+ShdcroL8vRMLj8sJA27Hnvjh+5fl3QoNVclmMcUozv19
H4JHFy7wNSp5AKomFkadZyVkTeFzKmPTI47ddppUDaYYe72FV1lrdh5AdaNj
Z0dshcWZ1U8pzoQ4/ecjjwaOLg6BAfbHVn+W2XAZpADlQJ5X09r4pIs/TjoN
CJBA045HFnJrMJxnv96zJIS8glObo5UJS3JUvJ+U5esbNgXHoIwdLhWoRFNg
mRu3KmprBeKI9LHAsJNwDrgNdVm89zOC0t4FBQd0ytMtuVfdmLuaQZ/HuwI6
6Dp+8rwGU73FHwzPjGGSYsDgGe3Bamm5X7xOsLCaAuuyDdtIp8D8uPdrs2cX
jtf+t5+4HZBAFhxAJFi0U5fvHqQTkBsD3bHA1oNBOkMICrEgcPJ6JhTu2d0N
zzw+krDEyQVXsAYP1XH+Kl6f/NPQDDcLwrFeAj9gqDSdUvI0L594MLboRowe
doAGNOqIqWwrNdpw7XTyjPY8xQ13LRNePuDax15SO3QHcuUq8Lo6f6ilp8OR
qmr9aWAGNuQeE4JrV1KyaRhcY4T/aNk3C/VN5bs4JU/MmD+nLUuXnpFwt9s8
96CGYKs60/2TAGq+O1DaPTXxvv51Bs6FjypIK+A1WZjSeGx9jh94YIMQxGfq
pD2QN9u/Z1sBJ/kDqJrM/kt/AhIfwhRPq4rFgTOzZHmKMPDzaLat2xLfYAFD
p07lkpZJC46qNUekcX8qZl0pKJ42f403koUeSNgEoF0fwopd2TZwDsKNe6Ey
/Hzm/o8u1T+fk7CW0To6lK7HSmrlZo5YSN/kkznY/xWj8CO9vjWQ5z1l9Gjx
oI3PUreoYPYtdXkT2kVmXRTitM3WIVrUsOPZJcVYWddONJZTNiY2Gt35iKsd
EXvGjiD8diqBshUoJoMB6mUSbUJNU0fpSQF88N0j2K+IHyb+i+G/NttaHcgH
2Et0sg7siPGMlISoSSzmEqwRs3pLNSzU+SHWPESFyZVVIKSogSDOKCO9reME
BWaG+m6KvJ5cZ2dPh6jcPaKlgR1DQsigP6y5ffbAZKEIfzeG558Rma2j4HEZ
hZOEuYk0IL/eqLpjO6EpZvp9heOdAaNrxc0kI5s20TeG5zfyUWYxJSTFu3a9
82AEb7aHfwpA3WiRa8MGbns1CgTaUQWPb4AgWfp54vCi6f5nSRD+xpqQIeib
Vr9hB6nBFuXKzJsW+uLELyuxvhGegvf+CWd683/3/mrjlZL7A9CqcyU4u1ie
HVJsOhDYe4xhspifS9AM2AzVM3j1oKIhctFwyIEunRWkBuVtEn5q6IiIZRR3
c1ls

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeizFB+pCXlGjrA2QzK+//v4xHhEZZOKyIm3Cyv/G5IvI38DrfoOB7oQCzclCZM9qLvU88jtDnmjje2uBkbuLjFVAena+ISamo8b5EjfaQzyPhc+uB2sOpTAXIEVYoyGw0dzMc39URn7+oCmX4muy2mMdgf6ZOhEMdfcTjURREUjfkmpRAEJodB71vPhzo2VLZNTUk1+rLWRDWo5AaBF9nN9IcvxiSSgR29uyQgfQzGqmDvnJPfilK0CfM6b9E1Q9D+I0OsjWiS0XxUWpTKfcdRD1QZYghAbdD0Ak9lm4nxjD58D5qNiCQRVMOuSEZw8k2sKBzvSoDDlZ5NGyerETbS+4KBaMeRSvydnjqS3ZMNclD5Iv8Tn2nJZ+a9NIyKUfx1hmyDhdshwlw3RjrVL638GrBaGRaIj6FUNnpTzaDP0TOdSI5ETTyMs2DocoDK/Mz3O+dOpLzAUDQU8bfJ4dINnSy6wos51Di/IgDumTbTdima3y92zzl2RNBIVG5hFCbkFp3wpKIYbg1CNLYwVVddtgS3pBaBvYOX12zG2iF1CCn2nZcfNsR31kT2AxRCrHxY7XpjWEUQlemNiIt8ZPhIARgHS2hTxLBkW+eaEABsoQxCKDN+VpJguM8ZL/lMQXhxNP84856H0gXuuZhd9crtbJCpnzMLT4NJitw7Sxysl8jUMUagRV+dGZk8lYr6gDxFNZ/j7cUq6sIfIEsoJ/+u1tUv1lvapUqh7Yo5AixECDxY87E6MlV38W3maIPtRaM/7pXEhBR7Hcl9SZPYy934N"
`endif