// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pt0EXY2sugWy4k0yD2Ep1t1506aLjTot9y7m9Xspi6G2T0Aqpl0A5n+Ia58J
tt6k6aI2fQRh70BMDhlECviGQOG0QYYwNNQCyz0lkX2SBlB+P/21kRu/gbkx
WrXurcy66a4MP4Y7gAr4ldp5T3h3mm5C/lZsvQXVrIYroSof0EThbMjMEJH6
Z2mOhan66mv5lHvNlwRZbvXtCDTjsPEHqUKwRebAx0oaJzfmwSgFePY7JtW2
IQz7WvH78iZt7tZ9cea/v7zmhferYnqMTKtvQcZwb82/v0sySchMfOvnrtin
55VQzx625JHIbIDQYJ+tnTqcb7ew4AYP5JNIohL51w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qkJxbv6xKM0Pm8ko49nV55/xEbJHXDWKRimeq5H35PntcPvrr8I+orGnX7gW
gVACQ5BElThWsH8GMrSxD1nx4bsrtPs2YPGiWDPJPra5O/uEqK41j18Q1uW5
IDv7iginurc70Em1DjDXthmV36rAaoRQdpSuhTuNEj+Legx1P1c6O5xseKeo
cZtQy/ZOS4oCIJH/1RtNCOQ1u0mLPNuJ6X3psrWmIQSHUkQqqROldxtrH7Ki
c4LyiMQHPBV+nD7E2WlMWRHG6v5oXv0HXvq+GvmuGZQj7Qo7YgDw2XfV99vw
sPn/jlJAssAEt0c55Ogyoh0qNvcrCTGRAYoiC3XM7A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ku5QobRMPxhV941+ZSoMhGdx6a5Qw11D/3ozmzwuY1u2wbhVHSA6EAaW182m
Dr4fBK/zAa4yp8Z5WaskD0PVl55hdwBmMwurPqxuAV96x9WJGN50mnRhvvAm
uPiW7+pteXSc24eID6QNCpieOhijHi7wNoE+17i7YwE7eeo6J5kjMe+1TjBV
5cnTG6+zjyowkgmmt+c/RVnebBI8FsFR/m1KmMG5bdD+a+TJSgIWL2g0h3oA
H+vMqJRSTSlL89Sjtb0+YlyrssJlhdq56VWAj6qLi6CpyLZyZQBYBLkYmqxP
bp9ODL0qmbTGOQRP454byCrOMoclAv1F25xHhfDVfg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TwdL4Fpj8tmQPIJWtgtsblakIyQ7wESTaplmbn0HRlYkORW6yYBn+exEbDk5
Tn63gUEVcXJcroI8XojOxT4FD0JKw1xQnCEl/WLhYVczcWK0aplPIbThZDjs
IgpczqERsw2ZuGSHrL5USOpjKL8uUbYK8b44HqZjCcCH1CLVxNHpPY0fT7JB
VOx6bzOSW794rrHS1nfjXoL3bxHqlze2waKYiwTRgS2nDjt9Gm6PmCJUlFRK
3ECtx2uVqbd+XTqpRsFBqtRG7zmYwG3K2dLIwmZFJjDeXtu7i9pYhzKptDDy
qZla1BOQMPTFEDLCSjAQw84rswJDsdDia6AdjVMDFg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qb540xR/r3L8y2pDWbAamz2lqDuTmLPSYNgwioJ7KcyPrKvsBQerjeoePou8
itlpnwOOcMq7mHUNi6SnnyaYsDDlp7foIPDCDwI3B41U4eTdJE35rNSqHu7T
+XP2Giib2Zw4wYsINusjnH0fYcd7UtHKXWZz7GXUTGZIDl4E/3M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kZMyyjMD3pweY/OhkvmP2sogAS9VcFUD8tSFTaUujA4N7OVHKs8ENIACyEiO
ZlceD7sb0RmGiinCq3y5Fjcezmk17ddYQd7/tphMNwpu2YK21q25gn0xcu/R
ePlzWUi0fJHLMJ7jFbhjSZo95vSCKgf5jPvi6iyvRxMclrJCSvfIx3L6bN17
C499gRlgrjLKC4QBbfYfTJZqhsnOFOy5eLw+RFcsJMmebCRj+hACTjvj6yTL
4FhApJKb9HF5AoWj6JKjTOZFdyVLZKrrYkGJo8hGR7TS7tER4oWzXcLOpfSo
Kz1RPd8kiKdzdQzYGOf7Wx8A4IZLt8P+s1b0L/9iVFB+929v66j+Z+bYWFPn
LcghxJVDfShOrspJW/8ibGvHjlXwKqsOFOapIcl4JrfwLDyBDahPK1QS4FwO
iylil1k670xG22DShAxHDqfCMY87UDLMJeWiXYqUb85XEq8xQ7axf+Vff+Kw
/n3iT4M2nxtJQ5EPRNbF4x1muc4GrTht


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TSbTShEtHE6w7WzwZ/A7FVbVP2Foa4aRdO9ImOIZIlmM575B/ss5JMN/Ldc7
OviJKh5h+SzgHTRRLSZpv/GcbVRQPQ46uQVy5LFxUdp8ZePkmnrmDQJT0mjm
bHJDA5+x6mkAOoDMk60FVwXjO7hj68zWOXUTyvWV93SKvv3TrQA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cCkDDWkDwN7bG6N2fHFxgl6zOLmRgj/vkvzC5tztIe36homKX2pbrupa0V85
3hnEgSAZL1+snN30Uq9w4vx30ins7jdVbLGxMNEZCTJ73zavkESQveRmvRzc
cbTCe6e4pCgdAalFqzRKVVAl6Dsg4BZABAi5vYkVZIHW+FW74wM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
CViW6GmeTy3Xm78eVLAB9WtfWy3gDdjUGNK8Mdk4F2P48dtyfRo1EEYLl+UL
RJzgkjmVu5FfInqK1Kz2A8j4DE92P76j05h8X/iyd+dIjHXzj7eRnuNejO/n
uPkNwXnkRESiYzHFIHJ/jDy1OTOzueCfeUfeD/3SZfr3Q3eYe5Vnh9KdDNi6
WO6IXFol1lsFOEei35rlFW6RchojNjSxW4qvkIkNg/CjUjc4SQDzHBmDRsXx
BHrbMtrszGH+vY/EZNoIAmUTx/O9RzI6Je0jrXeDwhhpottTG8QJTlsIzZFo
9QeuWpUDPsIEPinKK2wGDNQ5TYoxSW6s+j/JSPIBy0vjGOn6S2xGIKQyV+jz
OnOeXjpOW5aQfOf0sNDBgwxav/5aUPA5n3sMPh7mswjwzuH6lDB1vRdBnsGf
35aSNXqOlUaz/xNKDqcnZylREJY5ejtxiPLWtCP439cpLUXS7rRnTg1r4iti
oX7CgJRbiakJ2u1YjFZ91/iGDlm69PgwDxrXbtuVqMFeyDY/gOnEZhNjiBqu
TjEhcWxGnU8KhEgWe3MxnmToQ3HQp6f5WZbFJMe1YARfLGavKFN85bY4sBSM
wud/rDUp9AEocSOaGJH0INRlDP0ZTdMbMmd7ZgHH4qSLmU7yTJJcC/KlZHZw
ym9m6G/3hW84TAZqWDbB9Ak9ebONyZM5bldKucAtDPJQ2Ru6bD5pjI3OoGTC
BRgV7paGsPn4/YoEoiPJdLG/bnRxvrq2vQBIQT1XIHUyjrE3oo4jnnhT61Hs
7pX4w1DZgfi/OEh6UlFLB3Ln/E2RaU1pGxaaUQSCbNrC1nzOKFhN47puvOMn
o4GmTNxnOKAhjfQmzQrU0OpGARXgNkVAcNdkx0g00m8BhycgAwVlQ4VMAs87
Wd5GIA+L+z7HaeSiy022x309dMCcAvcm9Srdbg3impcy6bYGnomVwYApMaD6
Fg0EQgfDZKPKaaiUXj7FWiX0Z3QUv9L33MFBIxK+Xdj8qu/p6Y8FDTIR+ucw
+sY1DuJEnl9FNgYnCHVrTADT43SIEm/HecTaLa8rVGMcSVz/A+Bd8JH6fgcU
hWR4Tf2EcJKqB2cvVZ24HtUFNsemccmg5GEJtRIC3R81/Weavs6ZUWbR4V89
FuPaHiqySUZjG+s6RWIn8s6Kn8fRZ2JguqOceMufX5QKXtR7RmrhyrWSR6ac
Lf2KsHjwLlBPW45uuoOMxjnondtyiXmbOrDY6ZE2xKNGXqdqyeZZhM0lCU6w
yrOq4Shj2YYiM+PROwL1n6uNEmJ2JrPjJZ98KjZTGVJg7AzgTfF5zoNkdeYd
a9s8wyY6ExDrqGowSlFW+FD82w9cheS3+fTLn5UenGOJBAdlaz+Gwg0RMQIR
Id4t8Lc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqcCHPdMM4ruFCIUs5QiadC04xYpCZDTWPxUnQ3CCjwypaCvXjmhBv7212VEHc/xY0U3hwk7Vh48fk+ViPfrfc7G61kjuXZxy3RK1aFXR7UjgW4lWpDw/cqsCa+LucF1lPOn9v0HR/uklVHoBLIrzUYjJyDFsUhyssJfukE3zwmWp6MgyttFKkqGVi+HBxSjnp7fkdd3yQamB1GTY7mt6RTGTvJKiPrB3yMbWp4JXwQVpuP9bsouFYxpjb4vtakd0GPsoqgPh0l+0k0QLknQ++tDn18KNjL/saZFemk2oMrAXMuNzMoD1nGW/dkRjmMxxTHrxElj5d9+EotnEkS/mx7BBDbZLxnweNPjO0eqFCEdhA71I6tDRIhNWCF2uMXrDEZnsw01bIg7/2TW1fwkIh/S4E35unA5mtbd3+hOZ6p+cfJg5xMMLWV22k4VmF1SD95RZP83WzuYWWWOL3s4OdXydx8H/5Ymqd3RB+tOuO72U22FHBOkmfqoVwAOyEkG8Oz20EVQJWuyf/P95ZiVezwa91FV2txFyn8qUWwIPFM3zTvBgQgvro4tno45vyEoG+pq6ztbqazQkKJjd1HaGtXxzxUahN3SxtLgUT6VdE36UfqOn/2QgSZyObX2r7iaPENJKYZ8BBLHy9851UFl8aqac+uuikwczElR586uFTo6L8D5aTQtnFg5g8+FyfKhdWCzYnGaIu9qzhJ5tT0RzBfuw6HK0MAACI/PTukNM3gfvUFE2SAM8CsdpvAUZ7HVzOB6uFlpd2ORT1Gl39ISKynm"
`endif