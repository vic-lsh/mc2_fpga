// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bkYBdZlj3k+n75d1sTIxKvZNUbAr0wfZ4S0Y0QZeosLJ6NO+W7pMEuVhTsNE
hvio8+f0YPit7GcTisTC5HcQe/nNWMDwaKgxeZxC71F57O6Bundh2a2ANuYO
5is3V6ovOVaZoFMuxGjzEJeJechdmL/9kvKRWtr5nBZLUgwzO80hl9LjcD53
GQRwQT6inFXcVKn9RJwKjODuKexr384SjWTnRrK0ZKd4j0DUieGi5i+kaHid
5av2kGmo19auM69OdYic+Mj4ZT6FP22twepUMatPVoneDqA5mvPdLMAh9c2d
QcDNMPUYNE/nbZm+4GqieiluJLFo7ljqsJMcC1b4eQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ig/kZsQ62qC3srYArCT4HvT/uWEhJwk/jT79doKW5G4dYwni9SM82uYQZ3C6
k0BUB8ELonpwNCOqCZWyUv7Bd/qvM77N2kJ0qNSgurU8nPhyEgI7jW6Wxyzj
U9HylgIko0g6C6n/cMqPSM0/8/FSZ6A98pya4FZ02ADncntkUkB+WmA6Rc/7
GWvZ28YFseS2wbDd1z+UMjcxmTPcTN8qdcxt2wVTkNc/3o9xAlroDmG+2+Ks
ArcCccVbAVb0Bpyu1GYNNGRzdaK7dZsNh13hVMId+A7buvt/PeEZ+2T0JvwB
UU9Bk7OeGiq219BDisakcdcC+8cbjgaNlXmE1pzqqQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WsgkvgfC7Bke0urgwHmgkR8XOYZPVVffuVX8AYG8dSWiEGMeIhgPIcWyGYaw
bBGnzvvnnelRAzOjhUon/1iR+esUQRikURmpuMt7dqxLuz6E1jm8+dDjfl+G
HpR5DGyfgRMhUst2i1CBBbBm1JZrJr9jGKQVL29Fe74Q1c5oRhlZwx9pbWfh
BVHYCZ1XzEpg6cntWfOl1mUDu+2BksXBuSVd6LgqAODjiuVv4YhpA+Yv7Hg2
wuWdA2bqDf3lZi4w7YxR9ioAjDEAeEpXNOLlSADzpj/pYa631IHAp4rU1+ed
HzZmXS9jx5WodITf6Ml9bjjGmXfdzVfzW10xBuLq/g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TDeHmRBO+T6NFDghpKMQ7mfFLe0bjMr6vnE7dxiLe0mPIjy/s+8yVw8JSubn
rPS+pmbcVlPqJig2bbvrVKQHbgaTLUtlbxe53Zw804w8gmEYuTXYW9lQGZzJ
TThxHNNVgBF6HFcUg/MG4rfs/9KNQNyNRW2220Td/MimQuTdfIyEfH0bGi26
Im1wQF8goSnJ7VHZdBh59l+aZmdS2vFcaWo0LU4P537BY3W6nfMyg9pFMl2t
AKf5L0iLg/pUlu8yOkD3GwngaFr9y331wghPTSdYUMATSEQBX0069MUbF3ku
U1wn0Itbl54mzR+kMG6Tssh4wRf9QjFCSSts/CjPhg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sbhPxMT/Fs7eCOeAD5onrWbEJfmqRk5/nYHyDH1Z7MpJ1U/qKJ3LBhckRFX8
Mc4IX0jwjb7w3cMp8Yi8we7JqjPlncA0qcjLLEwpUMYTNjg7L4x/MFWNbME2
v42XL1zz1d+Bqzo72A+4P77PyW+woFbfGyq35bhgORWYEpPzh8M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QHxwC7jU2GxoI3FywUVFhZP9bd/g0QCo32yvn55Jg62Fss9ELVx534ZRf0s9
ZjS8QHXLdHv8uJVSJ8aahgMeNBRyx70Dn6DAXwVazeV1SY4B7ncnOI61W4wU
0QkULuxNRg68mat+VrVQBBDMUDseGNPyiEcSwys2bqEdRomIKT5Ll7lbFyra
F8ho0d7dUzFVuz5yfIciWgIbqOaq2+hiZFuFlwHGHJBG/igBkQDiMc0fswB1
btIUY7PzODKaKl8CcHxiWCZ3DrF6qLw5ZX1oU8lCfySQ1Vmd7neHapv7vK1m
KubRB5VKmjUFUH/tTEPEnUqrpfCa8girVFB+LQKDoGS1TThXq+1awC42mqhN
wLbPxBdrx842ode0vah3XGpi+AC2uNj1djKXAPHKYbmUQ82je19Z7WIYZ9hj
qpQ+/Dxrc644h9uh5Sc2hA1hKoa5EvrB97c8e4cefvYkHwX89cIjeB5XVSXH
/FHiTZLHHJQxht/56ADrhXxuSkE90Alg


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mJOIQ975Q/esUkyMwvCGrEPmZ2d3wbhTi69TwlNhoucqMHgjaR/JJSUeY9Bj
XNlskNTe+HA4Bu6l9uvDJHWY2TOJXQiaGhbOfJOz8blYEEltwekDpO01T0N7
JLEX1KZT+9swvM/xvhLhBloSkPt5pBSF0zgVxp/Ui/Gvh896emg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JYCO9t1AU1AoYOOLKjdmxcFgB1OiADjC4wLltNcaNuA6zzXyCAmeQOoSMtjG
yuow60o/ZgTyU51UmU1WqvjK/yJmzOjfuatvBGIYhkLr6ynIkAHhCpBYo2PX
GM+ecGXORQMwjGWTbdbKHSDnxzUcapVb5OJADs06TZwxe3Nlr/0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 29856)
`pragma protect data_block
MozUgHFwhlX+5kdCP3e70HYdvfzuoJ3QeF8wRfCQkwTLtV9PNme8NmP7j6qs
GO+qMr2+3PUzYbMhJtegexNOhxtfomDDJmkAliL/aVgvfgK7NuX3u9sSOWxL
ffDdJx3xn4eeq9nvR8MBcz4gBunWuMeg31s+WKZgjRyMYVnmHWg4I55HXEeT
T8bIvdK9Akkg3wlTc9zIo65+FqBaGl2T6zIFC6D35EMiN2xDzJgU9UgzKIe5
JaAINydKFHJ4jJlz4mz03LUPrO3bnu1I1hOFsj0Z421DXulIy/IpI5pcUi8O
LPmt0nvkG0nSJ65R5T8QFzUIOuM4Q7iJkTXeQ/IJ+69hvtiEhjq1ih3rYBUD
xxAgw2wTh+Bz6UX8/LO2LruYbXPXVfBoFQTDW8/LhsmvD/OiiCOvVBjX22q9
2C7dw22u0I5RaxGoB5JqWLYaDGEMwwF+VaUMiLe6CSXnk+Bjh6eZyQ21MFRE
qqPBMiAfCr+h5ACjQ3VR7rhVwOO5RsZ3WFSEnYOlxtkS1XP79Vg3R99zcWxb
olwkRtHZQ75FOsrvxBaCE3wq4dT4QihYmScYrWIr+/POpMwBi4noXnQI7wNq
+8Z5DDcmR6Qs1lMhzw4Cgf5GXvK7wl+XkDIFb/vLSuGehCLGDfMX3ecEIhAh
j1nNVGiewyo+DwxaOCLqoOOZnLHodaU86zmaIXfCpUocvoq4LgZqv/h3lRDW
yos0gN8T5HfC0pcqo091Vwf1ueSMiQGND71IxHAbBRykKyhxpjBQ9CuiNDw8
/Dmk1zLNPGrNqtwal54NcMwxNRcXR99c26TARlP2CU28v4DpYxQey3OHriJJ
qMaxMypwbNzitHRg1D5yoYI3brB6Ba1i0p+3AjkkFiM4YGMAgwrS8PZS+7On
I5EwQP5/Un3aq3O5v7bs7K6qUIbBBOT2crSRAF6sjZURKwAo1zNqDAh6IGhp
bi12LfRiMU8iU4tVVuEkDFneCJIzknGSBB+szJiHkZCiT+QIfKzl2kxi+wIX
k7DKodJBId2tcdTsbVTmRao2N3xGdDlv3F6jkgISPFK2VFANxUvav9f6FAvh
xcF5qbamWDrbQ6RvTezkCeyuj9ztyegKPZWQka8cM4+3KexdumxeQ7ICjlA9
QFWdi2tmg6VYthbveRootyAoI2NXrCCAC4tYp5kjakR7ffjULWngNJBwdgul
04vDFWIySnO+dKpOduYZnfnnoz/xUkPz9fee9E6Q/hw1l7/dRG+aESv5mvKp
mrGoc2kZ91YAcG0Zb3eXbFbyrpgoawBwG7Fn92ZLnpWuqQ488FRlVjZgxef9
+YWB5HKz7SQhQh1lpPKvlm4SKYYfmCES2Oy2PJ6tAYXJ9jgZ5RxmSJr5elcH
UoAYiEOMIeEdC4TP2eXzsG2vuj1X6I1glUzVO8amxYVta2hqdXUrqOcQmEBl
loFnnGZuEu8M6Wzr5Fiblq8bX/eZ7Ngy1PV4BH3WITEVteHobGFi0xwLij21
xL9xqxWrdEuuwFOAC2uAnNsV93sgW4HkuIVBMsrsMatUA7CnrkNV0tWafKYS
mUiTiditVC8jKf+9VIN6At40MHsvOlQpLKKa/jm4MNy+WzDbjqZ+yFu3X3iK
FYmLwt78zCjPUVdtsEd0XKqqHZ8L4bfj0D81TYzuRuvwtXEc5qDaUNJZdu7F
GmhEkaLgJPQZYJ66wQo4WPlYM/NE5wNCT1m+SiFKYuJQfsQJ6W87n/aLCgKd
yRAF4fAJH8fC+ntoJTluepTxP5q+MEY4197MmMBYDx3V8wpW1b9exEpYLlyU
+rv14hJFyYYz6kCr2/JdoYpMActX87fs2rzp9SFwguQN+HyeU17PlHelDMex
3X1aJN7oe/hjGF1k7fyVxa03onEH7YWyOOGBoyPJq6zrN/qQ4J/9OWa3VEis
4aoCb/y6Eraq71Znhf6b39JuSqIKozaS3WnBJithaWeTN5pvOuW4wQH95R6i
1QfvLHoe0iwzDtHfrfcC8Umarkh+qWxhKDIwrpPbTpJsk3/Tstl9U8dp1BDn
o/XXE2hbtXG+yh6MDmcuwGFH5kJUuMM/mZzX6Sfm20Dj2jHbtQ4IqWiiE6wI
ViGnoNU7SB/5UjmJ1VjyRAKNg60IXOhVbLoLfVe/Z3O6e0JP9fI1Gv7+hMSC
VVNiEnbqGU4DXMWzZ8hke7yS6gI0ziyvjJzkqkronRT2ERL/mTOWIbSNRIKl
xCM1YuT8CWn2MbzSE+Mm+AKmi/lxeiMvNcRKQCLjRFbPHcnJuiS/RWXEzQ6m
MLkpfezBMUPev1rp/D4RbnMDjWLnxy4s16YeeG/Z5378Xwi+UsAVHcbKb6V9
8lwv8OfLgIaOLA9DiyMa+eugtLyB/4x0qpgXgTorMpoocDZU9LE0Zg5KmeW9
MFHgHiv03DIu3GMTCf3Rv1CX6Zjev1bihwZTGVGXHz8yUoRUFVAFSzgBEwb+
qFdBdNZR9q5bJB/y3ENIeqzammf1GGZvhzCd3RaKAUyvRI+Blnt/I7xiYRfk
GVkS1cM9xqA2xFN63dWDcBTMVzwC6VWwzmaogmNwXsrnDxLeq9cnMazKMa0h
zBn49VX/xNiCre11Ps26YnXVaT24el9MfLZDkK1x1X+MB+KbcJLmdmSox3Ht
uvcj2hC9A0zbjkD6OrlHGYhr/yIvDNHKc4f9Wjua37R6dx8DhLI2EWTfF22x
THL4XQyqZ7+b2W9ebBTZXGXhQq9VZHZKNZgPyxCIDBRuGATG7W5QiOU+9qEB
ICs/bg6AuBAwPSvhdxhtVD1PPGfJefi5EwG8NjlbzgP7PGZFoN0S2hxF0c1A
bHyRWNwNrHxbsJzKJNw/2S+abM4Ya5pCoLEfSpcl9BwdN0kDs1bEUS+QHFp5
3McpUfntWhRFiTqw6bAcFsy/75SdDsWl8G0H6cm8dHOTs3GWXrm4NK1RqiqO
gF9gXoLOQENQztR/u32zb2rMhfVkqZZ6TRB1Behi+5mpExzYCr4KiN6920O4
OM5/oTeOx10wX0SfiA8e2q4pux32Ga9d8vEayKb6/1S1URWYW/KYEf1xvh+p
RAyqDxNefstM0pb12ExDqzsbapwYoOBWQnTaOwG1nBwAZ0k3oxRQgOxQwX54
5ahwEjFNxYCbA6oG1nDuy6Ufo7++bAeJOQx/ERNukEkJpLgSXgmXXgkDRv2i
A30FiQOtGiw5MJ+RxlzLRO7pQM4UxCDExGZRkJjnmttd/HBq8CIp1tS7S8O5
TYL8Vd3xHBAVdO4ch7YChF7yHQJc48POmoq41jWDxHLm6osf1iibiFM1o4lK
Dr/cjjJlb5B58wFXlkVPZSGMx5KHHuPEOnL1Urm4vh3QYFDPDsRZ1pnTOPlY
WuGv0s7Sqi8R3CdIH6vbx0peRK4ejsgK/CGrWgfN/TcpmuXyHxmiY+JhnF+x
aNKtr+TN+KbMbnWFaYgzJpC2ONwa4vF5jbmmjM1gJDXdXHsaCwuxHaebCuV5
GPIhvlkK7iMA296ODr1BLpSndfVE4HV7isgpnROrerqiElz3Z7TxNh3UaKsz
S7zkEb8Fz64Ith3lAzG6tIaKnfyADBu/4AdBhRpTNl2krDeCfBW/8NRSZSOA
RP2mR+nuneEEfqrJWk5+QGC7S801nKJJmzrdDSHd0wV1q7AnqeH9YrmL+iu2
icT5+fGpVfX/MVq8czCH16ER+FwORm2tsApshEvX4wt5IfUSYwReVseAAfmr
qxKJC056LSOuW5tx+wjicdz0DVFj84qntoRiUcuEJgvoG7izc/+8IJqZRXZT
61m2DNLtWd8xAUQ+bBtKAMGf2l56n4NkwRUlDw/Qn1qW8y2NknUNEibdXfWq
lG7HPDpnaJOSs9OFwMUoSnuSEwal+fOc6NCIu2lae7znrFrVdrZsD+ipyCxm
nmp3WHpJPZqhYkYa7gPQgoL9ERDllRmM6UGYnRsKQhr6Sryuhq6TA9e1/qEg
yKcQvvY6iGrMSTazOfirjQU5XTj6wCgrWq0dgFg0lhJKAqJ76KtoBt/6VJ+Z
NACZXc+KWeM4qPpA+HHbTGl/QB7mnJGkmKHKBzLwAXbg09yAwQ+DAqP4ibo6
b+sb7rwxaKIKx0pSbiqq8DvWC6W3CbrPtxMndmyfcplindyjyx0bMZISDgmb
96mRawmxTWOjsO0SdPr1m/nVnWeIqCL8vkYDJr6SYVap/oRxaMnH0nUeJmSY
UtYx7TLSvkgKQ8GiYQBmtaHpMR2v/O9odc9z0VnkhyvYFX9LrLax2NO3l6Wb
43AxTKR8hm/tPTlv88gXg2cQPIdkKfxsjKM/noBdDSxjgqr0qVsHg7hvzIev
MVBzC2aXcz8f3JwPKMabma7gGglz+6AJrm/EMNDBjjQiNbnEM0hEOpNpTQUr
rE/3/+Oyjb9k3lriEmJHlaXkOfKVPYsZta3T2ZNqImw8XCMCBbJ+VoBtgKRv
9rc2c5bGiu3WRp6ISkaDh4RRFZSjd0afvOAll2LJzm5KkJIQG5sObUlXkhsE
G3AQZDa2KHIs56lBJhxVqUVPcOV/eFoKUk9DWTGl2Q6/ubxtTcW7Wq0PGNNj
Wd1tw3TFewcN1KGhv7jsW/SZ1jEXw5CKVNQ5Z3FKmIxohQU0TlQJoEHU8yIH
I1cHo79OzqMINCHT+EUKFBEsJARP/BhHl/ECGEoxZjMI2X/NKBRtSsTl7LV7
+V44IOQIenPDy3M8P71tujQLXr2zuw3EjhiEWMq22VJL4cCp+6BE4y+7c++Q
TrioIlI8HMJDTp3hFE5rgpRdXfNaEqarfRo116N/71r/zWeJbdcSLyT0J8P7
QIzGvctzUdCI3ctIW8AjHS+iZzUqOvSWzyaY7DieLlUGiPSZ63Yx33lmQEaR
KRwDKiZlYozsDugoxPQ3T8PYDP5LcA183USGqn70UxChet1Vh3HnLdDihx4m
sBiBkNKs9Y0v9hLQPAu6V6NHu1xdwr3E3PP9w1Wu3oRGXioZ8T81GZ+Rz7JQ
r9nzdVKLDi4Pd2sMsKdSr1LaMElD9qOPma9yvLgWMu9KFnnADMUcuOXiuDuD
/E2Bkm8EEfg8huNw9xgxDfIkfBf7G3x2lUwXf4zstIGTLojig088Yv4P07mf
Y/oxub990r8sT0LgJzpjIewGFj8I3z58EoVbUplBT35OvGprTId6TKSE65cC
aj4dKQlR96YfzvTwAVyc9LT3HCus9ZHCINLR/2Ie+n28ksnaTr33nN0R8Gnw
l98RjFQCfUVBA4SYm0WcWT9N+l6hOWm/NsDQH4Yo70NVZ131Sw1Wy0lDXog9
dZAY1gSxGFZiNJhz0AMs/gwLmZTLy36s8VucXrZxpMOHNnylnP7zee52N3mJ
98fOHzLYWcN9SST0sNViMv6Y4a2hmChjWst/CFpVkH0qzG0+1mLAcmFEkn8Q
rEaOj9Xj43ZXtK9+rowF/dC4uYy1iiGCwnOqeTALr+qgc26D3tSthDZqt09e
fqauNP79O8EjlfocXKMqB3wfqzhwTpzJ5XXMcIycocbYI6mMfPdY2KlIsOp6
huKZOL9rkrxIsmXY+0A+wBDHx8rlUbrH9atscebh5EycFEY7eIFTxUkzbBJG
qk3Hn2hitokI4cclKh5MSUuv18JiiGjQTmQpWoZtPUwpEwFB72S3IrvHfG2o
A+gaV4iKmIm+LsxNxSFhOTFVf2sB2g426ESoKhux8VigBJnVZ4GMv7L5Tem1
DF3rsPR2rD9WTvpyWpN7Z5D3F7llbqky0DbO12qYPP2iHwoIoAAPwWzBC2dV
FxoGRX4bQy0Ub2ZGgJOScKeY3pKZhhB15Z8mx8umHHfP3o4+AN/8QDNUHgfV
OA8eMhUZH/qeQKj8plLRg3rc50DLNdJwH0VHTZLXfUV3Afw64v53IpYNKXjG
Xm4JU94mJFjnqEWcNDIE/AndTiKDQfrTLWA7lgDCb6RKRrC+6n1GPLXSf4ZZ
P156fvQYzny+lVlxzVghSSm3l4XxAljsEKrQ9YrC1vuFU2JwF1/rHVFk+biW
Oi0KcSvP/cVtDXIqrke5oAO87CXdgRpiDZtxO4IPJzZh8fP1SCSE8WtSUGnn
8HagKEKj23uLw3vbTV4g4Znox3/R11t13NwrasFCBTaXBRczpWk7NC15KzpG
OZcZGfrTQsbINYtE829XD35lO4m1oPMa8aaOagZ682h2Q9uwNvZ5gZM7w9Vo
78mqPQ44wAs1e9Sy5UnTRP3GmJnLqj5pjOCYDz2zHyKRBpzO9Ynm1T3JxwjI
XVy2Q5AnUT4VFmeUiKNmqF9oRMP8c2ceDgCLSv4el1FAKLTV523JWj2c8CSY
KhDYQ+Os567f2Aw9PzJdoXJTxPoJve0378OaRwkvZbiyCAqMmgqfBXIYdVuv
yCRUVzWsNdxbsFaSs5P0IX7IBKcbBYHZcCzROOq5JImb9KfUQFawTOWKNYeq
VrrGS8vy/ZHqeW/oJTgXJdwCkv2POgKhVkzMO+9o7VDpzd3E/AYqcSMGR8+8
pq0G/dS64Eo7EIZwml+xeD2BzPUAx8lSX2ImMT+IHpmcH9iqeErCkPGrut2T
qhJrtpQU/Q89ag9nXxl2GHteU1t2GCG76xRCJ8nlWF7lwHEPdL6dIhDqloZR
WQFg2nySl7yoFsSEvb7vsqBYTX9PER3K+O2gApRoqIyjZXnmZWsYirSQRM7j
yDasJ7nWdWmUCegwnVkp21ednLUQncinN4O5ajxLH9rYJA+8DZe5TV0njCX2
26o8XfrnzW44kZMI0Uxh3h0OVsv68SrsWlXpIjxv9z+v36Of2ry4t1a858WM
t9k2ybr9dgB/ChGMwWQW+YTtCvIet5HeohYs7T5OExN9FLz8mLG+ICc03NBE
7Q6oKeLxXRZAn4sRMjREF4rDD4Tld8ZJxGkB22Ioclgn9S2NAoasliOfXSgL
Nkzy1Zdkj9+A1UGXp2GMGMYU1Jrq3BPk0vAiiF7Mxna+LStE9nFtkhN8vTBD
lHzlko/z+IXEe8cXmN4RNKQQqscWClpkzDyw5HLSQXcNm+UZ1HKU/kSctD1Q
UYohiciebThc6cEMmb7hxOMDcEjB6sIFaLpTZ+m66CHBA3gebdRBgGgwNQpC
erVgyobh08kPjwqy1Y1g/dnpjwFEdJOFL+CF0N/IEfMc4qKA2zXwQnkYXRZu
qwRb1nZJVdKMPeldDtG06Yaak8b6QbFYvirOZ0iGAo3BflD5h31DEuy9o+aj
bhQlBzgFx+NvDCwoFGa47pRLFutjBPnmlu4SNEEmSLrkKyulwsgPrCh2TXFq
Zy4x53S5Btp+otYcxmkMOzDHxKsyICDaDrj6O/tDwXq7g0NHXfP6CU/rV+90
QDa21o4Y4xshltF66L4AJFPjsGjT6nvG9P8HhmdNu0v+O8mdliA54WnP/Kc/
cGBOdU3YVkyr1qIdgF0rYXfoZMRx34UbJz7T4yMIPQRBjPok9vxm+Cx+xXeI
rXo/xeU3PUP++wCLGBRhcd++034yV5iFbgzDmPNrP3MFR5QHb30tjSUeRrio
tPRrkfngpsaucFuGSPHoOuIZHGSP1T0OlEU/YSg69AdX0glz5VFHsKVK28Si
0XNykIJ3ECGusDmA2l3A1F6HHQnBgOShFhCgPd58rqC5PnkPH8oPmo6MpU0L
9TMn/gkOJTa5hmqRiRUkwocoH/ZeFa/qo4n92t5N960hu9PmZPghm/M3lukj
M9LA7r1s3vqJYADLgT4LwWqN7t6hVQL0dGrCunWAxeCV4XdrHtUseTDgqkKr
tWUOzF42gq/LutinYDuEKlYJenAXLjGvz06Lrx/rAxo7QiEgy61zyuuQJvd2
put/HSNTsrMIoBXcR8yzIsbAihCCzlNDDYBNY515WwkxGbJCSvCiL7PcaiN3
2iYVs4ONcjljNPO+bWMqWGF6r0sOQaO/wl+vaJ3mWbOQqk3rLG9kDFWMuwvN
fsdaXnW3DavhFE3PYt7f67XVEbMTuSV4VaGdpXm4cNUPTv3mWGWAT79PtaTL
q9MqVUC2wk28hbE0Bcb4bYoiTB+q/ul3KVFUQj5n9t2zaZm37T7TxkHzK2oF
et9UR3xO0LVsqt6eyC3pANYh1YKntRM2N1N56xSHgFhR70gaqHdtoN/OK/CS
ZBfRS7H0GVbn90AkY3Xrp2ijKqSlgI3gcTiq9pJ96ffgFOF/SciejxPOPcgZ
tOm2B9bTmXqNbRZG2aO95AisuCXz47uCnLbyYYantIoXhAx5K/PM8KW8t809
BW6BLX1j78P7D0STyNxks0E2qVq0GjLbOECALZTtWLDadAMtJl08lfBYC4HO
UNWC39UA/rcE4dzFKQFY2iewO9x/slHAvtMEUgu3WCR6pYWF8tPJabBhB6+2
eaDS4zUaKh8RbapNFn0elGi6JlJDaArAiU7HUjwsRyj7KDjNZI6m2chILubJ
a1yclV48Mavk5xDHJg7s8V2bVoY2oAcg/urDeQ3EqFfUpBStEYVo6gC9PWQi
AvytM3FDwH85/vjv/APhCEGMCZ/iFzcJ/LjZi/fvfE2DVvcW8iNXqIUP0VdU
vB0lSTwgoVBQQxhOWEUay8hMhQdP9fz+wPUievS17oGPEfz/fRYHW02FZlZS
n2EbElbDK8yrxeHZs0vl4ATyYcxoexm5BG/NQWQze9PdbdScAOMExjJ4wSNY
N7IRkFgwNfu8TvmWRmAvIBkbpWTftJfgdWMI00yriYMOKyAPwIheyjTl2MzG
REW4zPWJPKAip0mVjmVt6sq66q4YnTVPbevLrTczw9FazHS7zdu6+JSO3A2N
767X/iXGJZ+7RJhD0SXRJBEvOEP5vPpExRaNi0i1lFZcNXyJ1Psixv0Gt0fE
Wtv/ywgOoD6Qmbl9Qbpg/R2cZF8rLDDyb7veNSAtPExH3cFkIGddFz4QWBIx
03cE6sfTSov4q5Y0OP3WjdR0caSm76ZaQtejOKhzvuhlNrJdL6TIgcG2DXb4
6A40CBy2vlbBdUs64q8tk3MLxNU9dzBZUgJDTqJQJwx0H/o69HmdNKoGpw73
sjW5IS3yzE8VN16M38AjXJ0bSHyY2H9kS9wqCGkMpqoFRoHRNqM9+weD8wJG
P4I/5NAWqTDvacC3rnVaeEbZsjD9e8k+E8yKIuAomIHQDht8yuJx3eNMJvqY
XtK/RfNDsKGyb9w2+viXxqvs6eEEMtWC2ADqA7lNwpx4Zs65aPiKBXv2SGEh
J0INR2mR8prjYNXe0NSIGejgHX+pqrLwG6NK3xYBWt4r5mkyoR/IX0FJTY++
y/pEN645GmK/5r7m2hVou2PL/PVD9I4qt9y30A9nCGowvIIJB6O72T9qJeC9
h5XVuox4jV4sc6mGTOEIS53B79QJiPnySwQrx5/aTiPhUuHB2Qu+v7KxMB8f
kl6BnQ82j8G48ulV67tAjQwrh6Rg3yEP2gPee090Tw3dPFm0Clf7PMLtGus4
u1sPXzeccrX2UYM1W1rCl004+Kxibi79yqwWrxOA6o1sxfQh7Rgyx3PZEGL9
5kUvTMdHkb5XGbWTBkCoM+I0BZkqsuwB2ZlUL4S9rkNBl/OdPE96BhmBOZpG
vZBoWvBXWMqOVsISHDR7HDsPrIbgX7A939Fw7ktfFTxIvuuodzMFHovLHKjq
92zM4e2hnV87JSVR/BRY6jPy+CE8hp0Sak9rYD/SyYlswhGlz869ULlx27xN
BhGh41XLISH69IlYDskvIYUN0tUaq3SgVSIiG6RCJaX4YpNkhdDCUbSBBW2j
e35iL6O/QZgW8Zf+E4BAFrCJTo1moJVR8mveKA1Ma5LHZxj1l+oscTxg8xTP
XrPLxRildcXcIcdmRCBrIW4W36DkbsqlO0j1kPcqYlbsf86Jjgpu/7BmVeax
dn4ixS/AN1B7HdWpNNtqgHy2F7b/i/P+jtR6k+ziSpBzZ4KSBK6/wD7MYY6O
HCt4SpuTKaIcYkumFhUATuUIE+M3zjgQwY1Fn3OvdOGH3NfPkU1UJjyvRdm9
iu/uiNKeQoFA98lAseRPg/EIPtzcPyfcCkXc1Ime6SvERucXay71JBVeX093
oqiIEThU/8OR6PZWFQF7vNjeQLSJ9/lm59RZDfy0oFkCr/7nTo3LN3Us28pO
iXSNITYvliWuX8YQCNNcltiRmTMrGjhVF9/i9Ru2sM6X4rks/pv55re8niIA
0sYa6gW0Ag1DB6tRd/TlLSjqUEXktfRjHtcUB75j6qD66FDp4NM2APmD5dDG
OX0sYQD24WwQi/EWA4sDVRA6O+sphtogZ6/o/RFvtwYDfaPFveVvpgtyAhyk
GdiH5/rrDVwXR20cBhMpCn/N0Z2aMVXUD/ipILYtI5hvY8kgIo/Zzkf51HCt
zfdPMdHkpVLd3Ym2fCPlOO/970iHwuYKmr3x3s/gRgQIKVF3nyTzlX7F4dqs
gpf2k5QnYppwtqQAc/yIwbBQCKO1er/mBX6TA3sBHNP/BHN/6WzeK5U/+hny
Srtm2zbsrpbWZ/aVJ5hvoBr4f7dVULYg/3B++s+Xj6YNOMo3AT1QBHrmVXzf
csfWRIddVM8GXv1fnJUZvoTVC/7icR+t51crCWeP8v+KWMa17CHyZ4t5AbQY
PPJ5rJBm85MlagyDTmOq/016BYEBMy5J6SnJsmBoM1K8aFL4UJ2YMmYBP70I
eeVw16fqth8eMalGWDlFbPqjOqgN+OL9Eu7n0kebnIx+qamrZM87IgbfFOd/
jOH+VCQOXJv+ZlECiTrXWQhuPKPaDggNmv3R93VsDCDYzdPd0LS2f2fzqOtG
DN+v2N9xEadcTnvqYR14MmSzB+4ljmGigz1sBvfymGTqTa/v1zmRiYqwGSS5
hoVX4JfdLbEdUeZ+X+Lmyc7ya95m8DpbyaHhlPYUMwl8dU8OmAGzitqD1NdN
DSu3rAil0GjNjn/D9KzkYaBw056/pXzRJLGgx56vRaG9O9blmgDNNrJJs71A
jZBL7J3eMhnsBg55abmTdHbpGCbRYCOvDFnCP0N2hWq2YmvYIk5CkCObzpck
WwAITmCQPspsCcfMlrxm9SFAK8b91GfwAsxslOoi0khyjM+l2Rf3eYiCrTLg
+SNutwM6ISCVgGxiHWw9CY/HNGTpVL9jbAuggXGGYqWVycTj8Bf4iDu2qTpZ
hCguB0dsd9JW3v/Sc6L+IzNZ5npcXjQ9jjczTRuvgpNjBmrQ8mXteBNFiG6m
Tmb8HEPS3MSDuKk+/72gysHpR4QBQh9jo0XH8hHwf7PP74ek7PX9STJki3ST
ccq4gmt6XAdyK5lLfHjvRHweaeVOaoPlIgrKiQqd/ZppghYsAdcZmfZZDuLT
JsZ++pqc2+ENpRP2cNKESyjRjRN7Sf8O+bHQaTI2K9sBsv5X0GOD761ekCPr
QOTbM4oxRNPy9+nz8bnqtxXNymzCRKjSVbun73QeyT7aY6biI5LC29wgtHoR
lGbCZ8qyt7vlskOZG8F72ooBvy6JGvCTpw7Fs7twjPevCCUJ9+GYl1iCHBXE
E+V8TWmp4o1QbbNJBkPKMdlJTgsQ65UtKYmwmk4I7P1b6HEGmtK0Mkzj/P/K
hTK06iZhs3E//Ry1V61aRT59xYNSCMnZ8GDioY1Z0n89W5kEe7SLtMODIGIO
tuncBjfQfZvqakiN7lZqG7keirFmWxR43LVHYWvyD6mjc2kEIntkYmOgxj8r
D7eF3Vlx28Ytfn4yRqDGcq5Xon4uapcoSokAVc31tE2y9uUGt+GtLkgpTTsx
TXCIlDPJJ0VK62p06IARDvvOuUv5faMeQRJIau07JlepDW+gxc8RHS/FAPQb
PLGK2acv4FF5DeMDgxE6YfrBO5DKwGVPoZArV6Qzo/t/hj1GRU7T1c/I8iyi
Vvv6LcEECEGX3/lMWG9wOMXbQMZVRtsGU/LMMLsG8gDplFZ8e1RKuvpD28eJ
1C65XokMlwrX2QU6+cTFHgPOa30kVLlkb1lA48wiwaeWeCfPhNmMTm4k98JQ
0yooKxknTUBnm8rWb1yGyo2ENW4N0B6eB+Fk99t9BtUqM2cSyE1Enspd7g9e
q3nW8f6XMzx5flhw7EulCzcEwRngISFqHhwuxNf9byR1e3OoFhS251gk292z
2N9G9VpYtKLTRkZE3SMjnbYZBSIJdQBuEsCRZKzy3ZYn4frhAw4IoycTeMEO
GPnxz0FLtSPkvjZnxcUtBPpEH31j16CXWwXy16s9BbF4LL2cBJ0O3HO9LmVp
fU8jyswEqBsDwrxrVINQr0QgP41+7eUzH1yeQZSCFQ3T6aGa4yHc6U7HXUCN
XSA6FIidZeZI9y9H611W4zLj9tMbVGfJXv9ZUx/ZNVtsnarEbvtpogSVrsnk
k6I2Zt7SheNg42XA9h9vPvaDJPpgPlaMuR6kLDhheCiDwVzbMQ1RXkX9ZeRf
wUN3RIffLYSAuqbxZ4xMXPf+MGwun/TS1X7HK5higqQzE1+AcUjnjstPacsT
X0fGxNvtnJIjIa82il90lotP+gZgjlaVYyF04NLspO+T1qGg1jRMEWsv8FUL
GS1EwmNPwrjnZHbm+lgchKNO1xgcaAANx7S4X8xgDIzqZjwWrHhwRWcRSbEX
xMBuKQjOEevNvdURVr3rfj3hA56S9V3nNzndnvu346dTQGdxauR89iKewgi6
6SajtyyoFzA3HerEO0KSMRNpE9hI0Czd2n960Jrwyp2jQ2RBke/ohFaNXWBi
49k7SNkaleeEMnwaeR8dxOkGwaGMQ+26RBurHyWUA4K+ZwZcdN+iw7uxMjgh
rprv5zUIStWkUBw4TE1ekuKCSzZAvMrmM3ghuUNUVMXXUYWShYpffmHsERlj
T0ioGAXvVSX5wmleDnbFz4uSTjh1lMflRw6t4ihOPm8zMBoS+mrwn/KsaWpQ
UhHr2aYMrtyw56r4SxzIUQHzfat77Olmdn7b8ucEhPgwBzrrRMLKUeZB5I2A
FNAi9X49DfUippoQf3elh7Ma1VGXNOTHYDPsGEZCRE0oqbOfpb8rAxEmgIkG
lpCdGTBhXEorxBf87ale4xB7OLOU+Mv2np8Fi16Gcvx303nUOmKzRmtIZIzT
HtYK1D8vQ9GFuoE0Er6A6mwEw7fIdrESIZ9mmwmVs1H0G6g+364lXv/6QiJu
mlLdY72B5ujMmKiY9NpevNSBgUPjyDmgk1wJYzHTUDqXST7XkEykYCLrzKxA
0a2VuhGjeKgSRnuzWqgokq3c6VH4NNpWy/rVxZkfNd0UjeSMHD7zJIPYscji
E3bn2OsyxaBhDdvlUyLA7oZmixtNe8Hy+5XFOu1AiNJiXkJr1QNtNzZ6Nk3O
fzypd4k340KAUizm1Q0jfX6aiAIpT1bk0F420Vorz9oEAyxFFDaq5ky1k1hV
L1KkahpH2sBhGH7stlIhYF5dvlO1YRfw8QX29n8Cse3NKh7PzP3VXEDB10RZ
QHdgf+fmhHY6or98eSn9vDbrRuSPqkv2WmMoF4PyI5EzHL0s0KkeQzgdKPVM
VsnsBX95WWiComLYZ3FZUdELeq6jEluZTyi5TrQ5MdMDb89rLe0NGg6haJ7p
wIdU+Cpb+S0vxMCjs+GQ2bA3mYZ3GVgh1L6p9JikDEJv5nGjfdHWwnHLorrc
clv/HY/QIb9dujf80StPaRu1Nccp1eP63ggRUa/RCCxpeNIGxy62K36UT2HM
/FY3fdmFSctkVB1ehBqjtW7rSKebGB3ZxsTJFz/DU0sHfRDe/PlCNhgo1dDw
I1BMtwlKQSt104wmiU0ooMLzPdhqXKOe4P7dpAfTa2D14oEfWRZDwBNjZnD1
uTGA6dXIO8kkJIS48BaCD8JKRuXiPePK+u1dTeUuCrKCR6utlV/sj22ZsCvC
oCNpDqVXtdeoiBldksneI8MdQz8tpyqjYZcUbvnC5riV1mM4lyv9YRtV+d1v
SvF8VSOhfFY3YslGsAqIrp2de6qyomVWU+4qfQ8kR3UixU7uQfIFDtxUHshe
MwMsplEEfjs+DsZwgijHgPR9iHm2zqF26e0ZGuo9FaCJU3okvw9PfH24P74f
tqZ7oozqpY+NeSi6vCwPV3VQ6bxhPflG0NqClfEJJNKFIcAFEFNW+SDQmLsV
AuOVgggnXAOmigSrtLn/fOP3PRR0UACWtVIpzGYW5b5WYmgHo+jQVtUjh0T1
CCMFCYAXvbif+op+L2rihIVwvhnIStMLM+/SHsEqmeV+PtZmrqLEBK4ORY4C
ZMTRvK/9lQ/1/CSXrITokWJS9BqCzO7JS4sAxPfWAcwSw1Z5VFK2Cm8t18Eh
5lzt5cuIj0Df8wrzfEwZvrn6/nUpJcDxuht1yQBjkTiqCAIaKMIsI6IyqJAY
O2/ZQPa6f1L+h1tLsYJ6iC0Xlp6EOWgTjQxl1ApZGm7g6sGbkyOQb/r+qG0v
yE4w2FfhAt8AUaGgY8/vHR8bmWfiNrGwcL8/nd/QLDimORtcaOb62f2Lltop
03N3M7Id+y0qcWm6pk03cJynqGABDIuM+jkQ65CKy+yHCarrYxC2NjvFbDOm
fPUZ9hUTNKtiffjJgf1gvoMIKdIpFeS1M9k1rq1sSJs3IO/fskPSC8vhl9og
IJoKcaoIpxUNyATJ+1XACmN5xf6E0HoZiTXYH0r5NkHPKk66tu1bFA7hkLV8
1PnddP3B0h4384TOUzGyBe6yDbbg8EGby12unMkHC4TWNhkUuA4BwTpF/ecp
bB9h0Ax0WtH3hUDmnN/z2tkA7j2/y2Ac7/BpjFZyiq+aXCarBSlSHwmzCG4Z
9WBgfuxmFB5WU6RO39Lt/7aXdODc8xfoyvs15i9Wbnq9eBEK0afwbMLWw1NP
8ljzzvHee8k73Xya2C5sECdGcv5qDjbUfqGX2X1mdsqIeKEiYF9JM0UsiPEa
WJ7hjpX3kTGse8XeDOIv/CcipRSVfNJSVz6ymKLZeSvkBIIGEUTd4Gvt9IuZ
8mI7ZLAFQgDJoovW090yeddMgmv/fBCWO00CKHZt0uwwp/Vx0TaAU/Mrs3hw
S34F3qREUfa+OHfedXYX9LV+Kn8fQzXND+g2Gnf/dIx3IGV8PppiwzaQRsPS
5GGLDCpwh3+gOSwkKjzn3LH1giDm8K+RWFtw5E31Ty+5OBfVpeE3DC+TeSBd
n60fWYmZvd0w+MZMYsJWGBeB/FxsNmWn/750hBF7nf9CFlJnwCDz+NFAwahL
PyqUnO/e22DIrJZj6oAim44/UHm/DX7HRf3cUkjlpFasvXrIKN0oq4XiUPRl
eh8x6Wl+ameRiglSAYsoQsztN24XdZZiPuK8bwtR0TgJd+KgKTdBBEz2n7bz
nrS+jbwWpmVxbegXRzP6b6NKNjvBW5EXno7ZLBXTTiOkya/yyy7fJOB2qa8w
Z+l59wGOp3O//eCmFwzR7b1hKqXIOGPoJq27ehuml05LLldqHq3xBRIrv+KK
Qes65EynK5MZ8so4N2WLma7Kz25/x8q9SOUJYMPSVo7ZfHoo3hlXbJEd8lVK
BqbPsAWwpczqfKl7T5FZ/p1/TRvGYOSCuUHRQzR72kfr2I20/S1HU/jRwAHg
IeBdPQEIUDz0WFMfFGuhhfuLfcYIEUdi6hXtftD/55fWoCGvGgwA1mc6V27m
idnqNN0vEAigNFd/rdFfJwKciqQf4styGPV9huYSChETSAdWXqDT2YNmfbZ5
F9fFv5TajQKXrybQ9y263esYlILZdLIvD8FEe7wseQvUxvc/iJiwDrsI2iPv
q6djgbHFvmGJftVB4GMeddpk4PoB77pI342bq+mQxKkkEeKCXaZew2+SLU3p
rDKoWEh+nxxGjXhTHzBXYddqVMz+G2MnegHk2RK3vKAqAWdNhEC4iSTuSOgF
+dyo4RnYsRSt/Rk6o34D5uz/WxH9TD7V/uMx2VFJc2f0Ow6ltm0sMKGP91GR
FZy1uJkmAy4Q6TedKJQ6PwB3+soR5Sb2YV7v/kojJaQxve0VCmb9bxVCVDcD
aRM4yyXZI1zzF2oUMHf7dAmX4rmKcqn4H4kj3Ab2+g/dRpBOiBDuNSt0KN31
l1D7kpllxTu2x40nbRQP3ljZBcJxF9dIo4PBOZpYJ6XAVzU6aSogFcLSs27D
QfQZzPjL5uO9tKLDRWKSzXOrAb/vlIHryH36ZuTmglfGfUg5ZsqkyeYAW3a/
5uwBabhKxVrCcofERlAd7JqVtqU/JlprPiDH59A3BOTte1OnWGgiS7sf0oso
DcDCyzTdl+lQe4ZeAD6Bg/qj9rgBbp8Yt25G7Nhbxh/1QtBqz5kCcSN+M1rG
5/4j1ksWWJatHd8NLN6MqVahFl9Bsq/A/5tofpB5raocsF5Rfni238RT+uD9
fKaskebvsOJtaqxzknFBTbtBPAfw1NaKffZVzLu6xULkdqvVPDTo7jKy4w2y
MTAeoj7TLZlxxdvkqouKswHDZJsDf4ReG6TtC+lHzyrJBuTg/pT5MijwAsxR
a8UXWXUYLPW8iV1nJhnVbjcBrggTv3TVijtZrpjbZfcusc4WvHSPqUzEpJSo
uD5VMx7/DniaoDN5ZjWo1L0N5FNuQQk1H1I1jeaqs6e1kLjl0C2KtB23Twtg
rou5M2KoxEYCUshaZgSL/L/u1A8yhv/lnX+lV8rE+F9yZj8xBkb1QBxfEQ1f
UOS4e1BxkTMOXTqvZqxJpHtb5G42TkCEkzg+QqVOh6WidL8yvGo1FjAZt+Vz
r1peK0dKIKA78m3m//46/wpj2mmqU/amJua+fzJNtX5KufOj3brNFQzaTwcF
3HA/qKkoeC+PHtdV+CTY9kUCDGcDC5B9cgxt9k7bRj3Vkvg9ysWJitsYzWxM
k1xKpOyyKdTN0nlEnVG20GWIg1JZMiyWuCtss+4ImOEa6WyT4x4mLHAuink7
nBeahLDhXhSZwUPNC5L/VrDTVWU/HJkpNA/2v3MEgT7vtQ9qThhrxEygRthF
2M17rdZRxtlGcxJl4E4bsGaYtj4rfhHvDwqdapZUc/nVkPEJm7uLXj3uR5tJ
gvN36yMErwfGxWpMdN02rrceRqv8ttl1gFD05BqGv8HTyNRxX6CTN8gcAsAe
tMW5LSkzwl+0ByI0t3gRH0zyvkRM2pzkmWVkwKZh1OrWK7AYgzKSuOaHPChA
pqXDHeMjckISTyNUyP7bzExE7A+fl7M28ONTTf45R3bx2QrROBbuGT8QTp14
Uix20xQbCWrMmycZ22b84+HPVgaXcouVLK8GyV1MpOMdKNKGHAze8Vw1ssk6
XVDApkCn98rgpP15UliUIgTdWFe9DGSnBM1/aOHvGDWyRPWfkvOsHhF7Is32
+JGR823ora2wIw9wfK/UoEwgRWIe6SQ3bI3mruYnxPyhD1WQVeUdoT/o4TGy
07aOjojCwyMS2WFTMwinsE1lQ20Shi/1vHgernGnfyw+ubkH7qj1JsncwQmm
8P76gv6LqH/cAxFpz0fkGgVHWVVMGE6GZUAEmoCe5Oyfj/QdU7QI1aYhy0Fg
rM/++plHB/PMbmRBxfv8Cq9s1mkMc1NC5XNKJRuT9oBgJWSpHni1T8+DbHiu
vchfjUsRfdLeuB1ZKHVE4LLHZa1OFHDLcUPfFKIjhFSku1MYYET8ad3glwLe
Pp9tnf+jW8tscRVDRr04u4Nt2t3rvYaFS9tjJZrlso9DiiTskAtaHjIe5p+Z
+5h2o1+LhVCXmunGpU4h5ddg5u6gH3BbyUD6UInFIz4NBQYwGNxpXkk3cO1n
xcPOHGrpAzWJX7LNlP+f0Eyp+Q+IC9ma7zHzVMkmse/qy7d5gtDPRpzB7vR3
xZ4d98+8g2Cy7si27lwQNvOdX7baI+ZYCmDHwzJFV0sEsvfR3SyJa/1vN5Jf
LNSFlL2AptP2kiSzFtBjKyMF/IeeAKhkAbYJJMRMKv663dn8pJqbzgEGUeM9
tLX/UOjgwxZ0JsBoNRfdCiPHmloWV346nzmnoMumpBtZ1WWQq9hDw91a83q+
+YnWZQJAE5VxJ4e2/bVNhYwGRlUwiTb8Lgn8yCN3vRivypQr510eQHmBinKD
oE6phgZcVnFkf4imdP4KaU6v5iWL1SYG2DddSSRkCOECWrElLN4pZcmRVDbm
POP7Q7zVBg501J/sPjAjueengq3wFsTMxDj/cXRSS+1QxI+o2XOio2VRavgk
10AuzdjCoZjrGT+YFeL+2Bha329NW1Po3HtsC6Wms1R9O6XErhwbcyW+r91T
uYfYwpcIWvaf6vXwqKfH+aIy+V8Ll9ry4jHAVRvfZznAYGiPA11dubN5lAym
EPi79qwqSrQlzKBxcqnxMOpl04GI891Z9PE0QjbLQJNKWVGIpkqJCntBzmAL
n6YmUwiIx4TxLtgUiZj77xAGPYegWxNrOjIh1CROleRCkmA+txgPXy1Ss/gr
jngpIuN8v1poRMtNGmTU9NsXe2e+TyRWUEcXesHftGSUB7Isp95xySTTIhLx
nytShaOEotzum4A/KNovmxSSkI2HI4FlB2/56y/H+bnQqbLypfpXfv1EJU4D
lrNIBmWT0v8D+LarcU3mITNMbR25boZI1IM+6ELKQBSX5Kd0ZM4xdQppt7mk
t0iPEaf3JYUgjjRWu7N8No0d3ERc0TUYDWOBmYf5BoEW9qG1FNVFemBo1R6o
WKa02+dqIEU/uCoi3woOnKgauqN3oSrD34/KdTKOxsQ833hoUOmVcF8ImL46
lKePRuTZ9/ycHOhl69+juuJBqMj1JQbFkQbuuwcVn4bxVe+F3N9+vKR1UhU5
gAuMAi0OnexRR0F+SIFlq3CV92cTiVz6eRrQDfsO+IxrI2EjZn4Ptm85VxZ/
sky1nVuCskCLFs89Jn3BtnSMA0tnnJ6WMu/Sfpwulgb2ELsaf3b5TZCsJMLH
WI294qEhgO8mo1z/dt5b2fH2/EvZjaMqKMVUKjZm3skYIwtI50ROvt0FHa8j
DPlXBnSkdj96FJXVJxpMfCcXLFDnu7z9wjmwosP8m5lG8kj7YNMWQHOVkzT6
HaiBOjYdolBqr+EvKiNRhZ+gQbD0XosszyEPWsfhMG4QYzouPiHWm8eba4WY
VM/3pU9zE+lPzLh27ydI0BHPeOyKjTJu6J5ZbpesXaSGw0wojI/LR2HU18p6
693jbv8XnTG4P21I8jWdrO5JsJV94cUdnWOjtJGhrJRXt7dtqqmGXZIoXQlZ
zk35quSXZmYs4zrLCT78AbivSXRh6v2pWUCLfQmkprmaCsH0W3ixuU32uVgz
EmrgR1m55W2jiP8rRgI4C4RcHxIePXDDLOCvQ50jFnrwt98wqn0TeRGc0pX6
3lu43bdiRua0RMfNI8sDO0TSQkzoVbN3zRnw0pO5UR1eG7CH0kbKwEwHUGp0
MXQ3WZTfR5K//IbHowFbDzDJxU5JEE/iBZ5SJinWEHL4BkcklQcvG1hBqnyM
/nlRVsUWHCy5UubiXawXWH4fj8gmTOk7ZVHRQXznr0ZFaRa0NKIHNKCHGIL6
Y6iSeJ8+mnWijZcqXQIKeYElBF88VJyJpd5CWA1GW2mV055hUK/z06jLErKE
oCEsvCghTJQJkEFJUc0GqMa4UHxB8iAnajTdmS1rL9U1dElTF07m63ZnxK+a
Q5fTRo/BQAX/NCTcvW1Ea3uFLOp0OxzcPaUl94RBZf9axPxSpEZCi0390BG/
UP3ykmepQpjRwt0r3ve1igoUh4woLDafir5rN1H/+9dDvzK6vyVAyqTtbJYq
4JtmFyicLC8WpWqlA94/hi3Q4VTIkv9MjcPX9vS+lEtxPT3jFbRTnyqWQKf7
VBGVcKRjxW/YuDIZNPM2hS7A1JM2tP8f50LngMAwRGz44AJoXsJCiavKfUqQ
ZsMgDU+gbxPc0Uv7ePEYM2xIFQocXbfTRowd0eGgYvVKh4RkNbhBRyRJ/EbN
+BmBVfLwG7+tMJRYaWqk0tk8DveienWZpsQPZOm7eSbrT0aqZFBPhHFZA3xC
BA73GzpuDIF9RHdRn1QFbhbPgofwY0AfWvjP18H9YLU0md2sK3rZCeHdAQI5
37niXtArvafecyQEUJz73t5I8XZBdehsXBgIiJV1B5S/4jbTCcG4d6JIdwBW
TZi0Kd0+jx1JmIvGGXOzQYu/KgcBNjbbaHQ0qViQZYLn40JMhGPNrq3pHXJA
YOuJTDDYxFRHm/wdzUDIX62JV+ISnUhsJbbPeF04yXhxfO/pONoNHmwPpnfo
aTfUlp+EpsKwcU09lZnyX+oFr6P+QWx8oKzuh/5lxSxTwmNZm2ZIYvWZtcyn
iRzplwDinPWJRoNc8Pa2x4KWDu7PB5IyHaaXKxjlTrbK4dhEOoIaX5mMJGGc
4a9qFNWF3eBWk7MiIYKqhuiHixIzEfeknNkVWl1ZmnoRwoeVhEP4kqUdTx9E
+BUZmY+gofE3wCiMXr6DkyXvoKFXbN0jwBSz1bcLNITko41RL6DTIKrzAIHr
pOYfARWkAxzWANt9abAzUkUub3zwY78fifgRKwn3HhISeOolFV+RtXsbT5qd
wKTPkvsqdQRbX1uD+pWTyCQuqZFuDfqMZxQ9k15zgU0yGYz86AvmAmza0sGe
dHbwdVujr9CLvk9dIRg4dxj+4K6xeAPGLKLE9+Ow+pE/aTIRsErPuW7513fx
tJVWhsbwLRDhMCkr1v2eNpm3X/95KXkhI+iokqA65QwLoZg7yIk9D0etzShn
BCcg8nWksMN0BRL9JUpil1iLVPdILN1wekp5QO+KtJB6D4YPIc+Y4tzraIKT
p5uYFufun3Q2SWsggsbGwm5IWTIzmpbjisnLBnRofOSs46sGfSi5w7yD7q9U
NviGwoZqVlLUvVZ3xSfYFgAnLslR2DZprEPyjbW6rzH5EvP/T8SpiFppug+V
GXWZKsH+wrEElYk8aMyTxUX8DbypXwBxrdtucHAhuTVbSdc05eQZX6vo4kkV
FaDKZL5eiGk6XsQvssFiagadSZU6noqwineQ0A+umn5sahHlr8BBxFk1KR3d
9Zvbqml7lK5NnEoZgd5qcqA1+aRruVulc6CUBJYJDFCysPHt1eadWFt6ujKp
EyiK/M5AkfQiwrb7oRmdc4ICkmkncK4oFq82xe3YY+fLOnXPhyLKQnraaWyQ
YZnDTajP+maYh3jkTroAoTgZ439F5rUNW/Ox6RqF+z6tQIQQE463Rf+jsHse
fjWdC1CDLxoR0khxscQlCefyR7QjE0EN4jaacHoMF2enj9cKYMn+Qp/LQT84
2cEMPUKRFxS0ihEePXKaY0hgaaJ8fLRkD0N53zGgewpiL2ms6oLzHGOgwatz
GUELG6j3KoAVEEuNRYRkMRlUOuJJF9DBZQo9CtoMIvYRt1vc1/uDE+B+q9id
bplk9W5pkaoqAhHyber3kV+0QHmx1DcwMpVBBowyYVhk1jGCcNNicfedMO98
KHbIZ/mwFGJFmvITSEk95jND2hMcfe8ADXzk904jjwnokQiEEQvj5IngjuOX
GOHfGOKDKILVtPMfEfmNwWsinZKbY34qpwJu+SU7li2OhxHWWQQc2cVPqNlD
ys8E1DD1rRQA3UF0NqrumQlV6z0l4RoMrs79TQwppp/UcP8NLuul6N8Mpt0a
RyXzrWU6GNI2QtIoUxVXLCGmpkILejBuGpxQiYzqX4ye3+jOQau38FpHnk7z
bUOxxthDsT6+Ya5M7cKBM3FCMwCRVI4mpLxIvaqeOck4XT/8USbS4chP/SKB
hz+qP5x2BvUvfGVD4SbNwq5RueGzowRy6SMfJ89Zx9V+Ca6hrZqf0MWS/lWi
9eCmYJ8WmQw9H1Z0RS0gdX+2vT9IhaODwdkqi1oXDHgGANhiwADbmhG+YvRI
V5DDaJ4q9qcopZpY2jjlnlJIc6YWa7ytH7HFFQ394T10ZL0vb6daL2qR55vi
C0qugfgsN0uCy2L4Hn2Vh9hsNmVBSkshCC/B9+BiQ2FEufNDjCPmlkyRCUTU
nQHUUDe7usSUujGn8ckEMYMvRY1eW7nxdx2cSBz0k4HWTwX04ps6mX5pwzN1
6EzOih9MBa1u7jSqYLjoyzNV3WtZdfFo2s/Epk2pIy4zQQNpHyjON2LH1cdF
n5KtvW+FcxWjqAzGzkxRcQXRC2760Wix9prH+uxvyxlu4Uj1e9SoPqp6O6VR
9E3gm6vh47ULjgrWBjWG41tsg+B1+1LSntyDCf8af7aF2a4NWYpoSkCfnP0g
oPVE+rgVkVdJOPjkEOy6kVG+OIErx3aB7XHWWhwzshsnr0f7hxntK3lmwcQf
96YXDj041wo0yBHGc2DMmogpTJNOzxkLhbLxWYcQi3R55sPuNtWccAGeTgAB
PbGXugaSTnxuz6zRXtyQAV8X3CJG3HKh3WN4rHR9PZKt4snXNOkxBcM8+lty
ivdJLF1sEdO34lNZus1w5xbQelXIO91k/L8H+HE2BxW4GDBjMdN3YND41cmA
pY4fuphw+JRnYD/hpN4LiyRGv+hQPL5XyzGsyrSG4VnM4e7FS6wT65YrCyuQ
UvxpIWvW93xi/jrRNUYGrfm2SWTJkbdMTh8eCrF03MUpTBzx3KzmRqXxYh/e
05pexX7dm/ABB02Lg8c4JgridjyeNzxQlQiOQpwQQ3O4St+xM+6AHh3iSJFx
cMyWAoiSwwWZ4Qxa0Rc3muvbKF2qEihmU8NQYSWRFn5XOmbTPA/n9GWuMrK5
ygNX7+AHjayFSniA9a/UjfYtMU02fQ079Bafh8hyFpCrR2hix+KFOWaxDC+i
zo3PyNquN/XalUnGpYyrogTX/taSWOz+8lQnWuY2VwGY/6g7OkTqlhVHK4c2
vM3k8NwnvdDf52xQcKkFhKX8NPX74XuhEaKg24vnXRfF84D1Cgwat8T40nNN
Jf0s7FlGKMnL7Hef6zi0wGS1Tzmfioqvo2ujS6pJ7q/q2Jdwdg5R1gYt2CwJ
YBr+KLWoC11x+3Nl1mQSAcGW0cHwx26rNulF9g+Wg3+sdwAHzKLvJ935wrlj
WuMoC5vk0oL7T8sBnQPoS0FpVnbwZTGhA5Cj3QVPWe4wsx8STaLzYDwRHfEK
JknPWTBaviUEqCniqv0FN0MiAjmGwoX9miPHHz9/Zp67tmbgWOBRKUTnc+Xz
IoR8FV4dPYFxQ+bnlwmIlnv0yfkk7HgK+tvxfdDfkAiyoKnJodC/ThSTBpvf
tPrMYAk9JX1SqOHdAJ0HSXPOon7oxLGLv4vb22IhlX5QZ8l1QKc1AgUlppbJ
QSjbx2PtaIDb+gaxgWjA5XjthF2CZKzGcBUtlU3sYB27yLExFCKisBD5c+xD
9tm48csr5bIRdoLzSAObc6k1ka55vCpEmYgg5omqwuXNCflWwzqFwgT/rYi6
4SuPTUM9HhJCFOgu9NfgrDiN9s6viMbjabaW4DrbQdUNMT7uZDFsSze5nIQj
TpY4faucinVyeYlhdZJl/wuePxudL/9hLPlP2NSonNoCgRrTpU3tx0nWOnxw
kPQCXshPbfKXf05+RQ991ii3Ii0RtPRYzKLc+3NVm6wRRq1LDRY6aFc/Rpzw
gtHHqn8xyFFz3XSI+9m/QN8Q7zmITbjacSyaWmww02OFC8Ojm8IfQnkxwLvG
6rHZM0NsfeL+NyjHUMc9GwWobvycj8F9NoRAkvpAn2cJBTm7+4xFoIX4NaNz
8y7vKF0Y41XpjA4XN68Gzv8qEm6++X+zpzrr3IjsRP4r49IlLNrx6ncHGP8d
tVUcFWEhNOrC+kpzuDur2K0KhwUFktjRVlSi9unvyyHiUtTd+c1Sltj2Kchy
S8zIKBUGMwADIBg61EXxL9YmBJpXja5IXcbLuaoapI+cEv6AezPQHpb9Yp4W
1Vmrwz74YAiX1BeSGTUEGqnRvVf+b/prId2gq/i9IUlBOJi968Nc91i14LpC
fs6eQ9kJQ59DtUBpht8YeshcHP5MihKGun9/rZVdC+cjKeOeh1MUycxDdcKa
4YlyR+GZUsirtXg+kQYLzD2cC8YBILKykV9VKIXGE2i+br6h1gMIeTd+lVE4
452xBVgW70wvKhidL2vorCwjq22y338xphu9b4yTQ6ynZ8jcSBZ8S3/jr/CC
dxm6CipUCLO6BvFNIu3i2IBlVRgHYjqG3x5/IzL619g65MSbduKitFJwJmwc
x8xxB36IJldiJ9oRww7jPxsTd7N/udURxJv4ltyz8GFvsogcqAz4yIHvtG3k
FDex/YzyOiD6o0ms0MvYcMuLqe8OkF+Iaa8DIFfrWSP3xJOPpiUgn0QvlY3r
MG1PS//8EaM4jXKUGc1cXEdAYbIzSwrdburCuyxiee6yh0et92r499g1zQkL
ZMO3yCHTfF9cCbYUnjFQKVea1zvBqfBACAaDgzvdp7BEpYhGtXojuC3DJMJB
qxYpGkGCKcbEORa4hmAto/46Ew4VZEjGkcn4jIXCoHVVSINqUkEhHkXWx6tI
y8QUPRIMnQkStwi2KPgAw6B9AOPO51EJkJt6z7sT8/qq76C2n0zTH8XQ3rmO
xPBu9q/ZcyifvhNDIfX+4ZxRMQmoSW6l2JxJQnLXAUzLDawuB/d+I/57DQ+S
jP4/lcMg/2miAGasO9UdCyQCuvhDNg6So0kRH9aBf6AVYQhTZ7jAvGb7jWC8
r/13ey9MwNyX9yRlSzGkiup8YlAOxzmFKwClOaf7FH/3cj7WJua6cLLoBJXv
tDU++K/wJlW2tews20pgwkN7V4HBs6esCaceHolgEowaq5vNQUaiJHBmw0Zk
q25zfWS86gVWqt+Soh2khTfv2cvLTEDklPE+PA/8Ha/qzUmUXzqS6TkOJ2S7
zapdkR3pFIi+AydFzECaWBsMUuLPvMWIfiX7NRPYeMmyZXYsMRpcXVeAH1Eo
OJCQdISvvnK6vUL24bVs1x10wSkDTI1zFzEHxpCCxlLtkBjXciCcisAe8Y+p
re3V004YjKUlRM2+AcxVC9RT0rdc+NvAj4mFfhj6OO413gDAd/iDZ23+TunF
mEo3le8vyDxYqyzG0WBcVunDQlem8idoIqpVV0zzv2uzvSfizsKrXIvktVd4
JWujBk/gc+KfsIiwNjeF6EKqQk/BIVYAb3/StL5d375+BmnpsvCL4jchO0EW
MsSHxuOvM4FvsBDk3WTWN+G80jfmfhdsehlPsqeg3pIYNtpPDVXoIdz/sxlu
/adXKGnsvymYw0oW7oJv6VoLp+RQ+QlnadjxpxNb8k4RKTEGeiXnVt+RO+fG
xA3/ubKO6sDbTtk/p1IFTIJiSmKA25IefNwel070hkYK3s3k9Zq08qi9M7qh
Y9Ub4RrgP6Ijcme0eLEcnKjgVfxweG0dYcRoar8hlJLA2GXrokt28Mb+NNPE
n5Q7LRXxWPX7aPXPRucA9ZC18p8ROETOEcELiETEeA/VMtNpNFTsl4BYLiwB
9z/Fi4bcOFkAaLrR2boLDfbGGs6iG5OC/SXhwCR9AJ5Eub37EKc5rS6wemDy
KWO2j95g1BJBp0cRBBbc02qlzO2CF6+0yfXybp7ihNS67iiRqumLv8pkqia8
UmMqBeDSeHqkEJEKunwhlJHc3OmC5k7uCYkn8itLHEofJYa4GOMIL3F7v7E/
23CpylBoVanVAZlz128BFgcoStKST5JACviE5FxPJpcowGD255AzEg2CqBPe
xBaKeGXazL41DHNlq5Cc77Y8rl9r9CiLBYsblhpaCFkJmghUxhwi1JyyzusZ
YtaqFEX4sOcTSx/TiJRZsJQnZcq9k6I29UmpOLiBrDDhYzAKOsQ6YyEghWdK
TQLhrd0BGEJO2y6jUmzbCNX6VPir5f12XeC3EShVcDhMoeqvsrU65p/0M3Ta
REs0yTEjBUkpRVPkI/DENYHmjbJLmwdbhXNJK4U9HvIdRYcilt/5zWZ3/7ts
dsODZBjspD285cqimAxm86G+lNGyGfGna+fiqNZEV3BycdzrXLKeDTLx/wb/
jaDu9kNX2Zqh/bDlY8XJAtgwWloBkw2m+zHkGfEbRyJ7dxnp5WR5iXDDKSpJ
wtsotteFBN4RLmZZo2EwmLJGH4GRaQVu6hUCo8U2gQTlapqOTQZim47xmIlu
/lUGtObCF0xo/JqVLldJklPcJYiddlm3ksBpYsn1l3Qnzv3PebRsp3CQE/l8
QIfaspHtB45l473htm+zU76o8BpOdk4p7KizTNCfr1J/6CWBuxoKWAEcCLQT
ZUqcWpgTelFN0Ne7WflDJXsbM2VI3c6xq1TEbgYaQYXZzBXqpA5r0IwpfxCg
yfUuQv4iHlhpETJ8ajDiMsPPTGtkt6KDRVZxNDQ4yJGzevQR9/ehlC34OiK1
klEHRO0Qy0QgjMGBrZl8lUuoX/iClld1o35js30/aNGkDhc5SDZO50aWYEGx
lapR3dBB96BqQd7Id3uZev+Bq/adZvQHrms+qmFiNoqZEPzaIFv0FYOTZQZx
M1WUKScvdl6ts7UQqdJXMMdr4PPdJ0VMKd2m7AO/y+rLazyLzDKkyGCcamhL
N15myyebwE/3fbTxijA4JqGvHnYRi/qRHzlRGr3ADcN2zlD0Ib/zUHekazKN
ot3aVM8Mu2BSEGDjlqpqL8OTytBjmPm1t/8tBfAUwyLKa3zaXTtATv0Gm48R
1LOvUJW54mlez8GAlScNAPTG+g57kmGY+m4EBvrDvK3hm6ERQj4b5JasYvGf
RejBKr/XjRgqRFviPWEqB8VubEIXep+wHbIX6tf4VEald5vMnmSJUeVWG9e/
HeJ5XWzRnh0sktCXAbBmbt6jhzDTXsJCZkT0z/y8bQbMuf8ha8X9EPKAHvY4
bhKlJXv/lWzhS1z0ivTXQmJro0oQ1f0jsJQ2uey6ANpQbbX1i6R/Htry/A4S
4CloSvpaacpj439A64kx9Gn2pdsHQIpTY1vpeJsm5u0qNvu8SF7SgCS/NVW+
Ak3GUu0uKWcwu5xibiDbAsPSE3wUbw20ToQPnmi2S0JAUegQHd3zsU2drC/I
qq2TznGrwsZ33FfVRYtfmlDmnbguWVc/tiWKaTSI32/LRRSSZODkpcmA5DU5
mlf8fFbqyskpIuZArvK/xmCPBHjfDDv4VojGfEWRdhRFTC6/Wy17zNO7XaDf
GfYz1roj24lf9NTLvx1fNhJUyGJ9EIbAHIb6SfWekO3pmKVHQXhcaVX+3ZSa
h6Pz3MUNmyzxijGQc0yYHCDOD7CTyDvkOWN7frNxZVnZ7xVJNXH0N0cxu8gD
4PZiDhykcPORO44GazeNxG9Pn2sLhtD+x79WQEL+qDwZndZFcV6betuFDDzW
c8GXFdDqlTwPrT44QCFtjZD9HkzMvpk4jxCtyk0Ynv1POlXp2/1bMhl3guQJ
Vh5n3e5H6PPwjXAUcz3w7TmtGWWKVQm3ve+fqOIdqd8YATHC5DmUf1xm1A0v
DAtC813MWUURt3NwzqvRxe4UMwPq41tC+YVFCj9IORVHMNWNB6STOy72/5uo
y8xd9ia+1hyHTQMyb/oxifHK9WI2UGEwFpsS3Mq2spvpcJ6G8JYml7a7ozs8
+2aSantamY1edCqw4AknoTGi4APM8UDbi93HrMZJejVlDfjnzMmvsrmWEtni
AdTwdDrxCLKEC0JCcZ5giqq3SiYp3BsZwvYmNcHMxdYC+ACSdffhcMDxfPDm
TDiF1CSnAcZ6fcozwYm03Lbf94BMjrKH21p3ugzOaQnQwXG3m9BvFqCJzVEf
xAFgNS3l9rS9Qeu0KHgqhym1L8XKP9v38jUZTVnIlPEHz/9Vn1KogjCY5VuL
/OSNzIyBCpcA51zxroJAOkSMmkQItEh7Y8Y5spa2UiMNuxvfNCthobxKttxS
gWDbz6J54poLf9tS6IHk+ngQPTO5CKwSqjoELsWhofqjzap5eu4SzDfNIgGt
0X1K0dJ00JQAyfixM//tMdilN+725wdFWT2JaWN4NUOXt9mbaT+QGfZxrcfl
2SuzAmg4upKFRBf/qvGGNr3gSzNkLI+UdnCcqKnUZXpn3sJUGqHjUMsnsJcl
83qUvo7Ia98zHCaRvzmdHqe9uXwr/OJu5/DOUdiF12d+f4HDQmhwoBDp+E/C
yLIKiSPzpFzJh1i+i/0GrlGCzSf7T7n/anU3K3DICdjEAZPxTxvTfOmZj8Af
Ue1ei1aRZrynvUkugjAFKo0k3QmbKeOIx8w3RBtV3TJmEvwiPCM4jt3i0Ppt
MqTamh6qktbyEQFsj5h9tT9Z/D7pcBMzRI0Yugv8KShUSAce/wvDH0SiUDc/
Dp+MYiZ5U1JhrLtt6FpyjRw5OdoNXaCPr6sIFJFX/1FINHyUBi769tv3Ycfs
cHQrLMkJp2qeL839tDk78/AbLmUlvAHdzGWikQ64E2sFOaDELl9zfXmdopJ3
dqbtUgc93/nBOu+NN22hjG4TbUFWLgJ4M+Wwj9bCjDxfA8KD+1LXqbRpl9Gn
07hRJoo8o9hsQJgG+3zXVbEzhur9b1GfrzXbiGhleg7+W8AIPNnfylgz2Y2B
qM9IQ+qL+rnKqm2imr63XLstUrDURiYpHjce8gau/2Kidhn6ynRc7DGJEQ4L
18u47M2P3cQX9/W+lp/ruxv8NYug7Pz6egMHLWyw4Tuv3LsvxMNIvvjpJL5j
G/lDGPXM5Hj+c5pv4LzaIck5gtPxmCqSNEMwjxtAAM2vy8Io1DVpV5MC86le
vVPRdXj7OyzpV9y7d1z+jOwE0bZCfyx6Kcq0pHD17G2+v6eriSz9WhvtHscv
03JZ7PXeC6VpUnS/JDNtEdOr9IbRb49k9Ir+BWje1tf9G78CBhbTbEGdJu8p
nY9B3sLqnhUyEMYHHP45Aeenh3KXKm6iIsnNq7cbY70k9uWXl2DlLbyhJpwV
rCr+sjJDq1yxiiwUdAPoULM2Yy4s8b5zxT4y94lZ6BAHcXoemphpUD03tT+n
2a2ZqsDzUmticTM275mBn5m8D/G++kZ/RoPtmRvzoWKkG3IzzeAY2YF9McSL
CiBnUBxFaFQ4rsStDNSlTg8UqZbHW37te+GduaYkk74gp/YvA3ij66iA2kDe
yqbfLQ4rtWk2Gd3fxOLM1fQFbI01bryi13DjjYhB3ZvzPeCr1nXR/IpzQedl
vW8a3mTxvH9eWJHCw819Mh1FuOtg0tzQtBBPtMB86Fd4fniilwxy6Le4JJAF
kkJYne797BuZO9Q8JLz3eF7CGMym2VTfvnx45+inffRErR3fgM14TQtJBQiH
/QpkWl3RRP1op+cynGcPIhNhObR7OkvvBtCAM6Q2/wtToDl2EGtcNM4GQFst
j2vBitxgxsG5J0xyH+ZE3/5uDXr4KF8zdQ014rjI6GxpZZLcszIBfh1ybTNH
g88U6BL+JR1e/mZ3YI4YoiOdXIOPGGmbxNKHRxBgKojIw/C4k0GK8nYAJUJe
pZ3VWFmjEE9NLVKI/d8zj3SGZz3TsAZI4R7yBmB9NHtIJrrlFvoz7VobDeLO
9gW0IHZS1Tsqh9upwaikFBWdnhv+a/6i3zbvnmZGGfyog4XqhNPnJyAzhO4l
YMtvKXRfzSZMCiK1BuUUu0VUhU7DMhX8/ZqKTlAWTchUCn7eiBPNX/IHJwnK
vAF4EVEEdvM1m/6UdNaRGQJrQRo2mkWtYLvBU4y0w+lvM96sKGbJLKOsgdLy
AiveTvhLtuuT6QqCUpwHZ3J5pce3jKSLCNX3mfyUFV8bR0BAwXtv249oIAgU
tgAkoK9Xs0pqxcZb1AyjsrujaRvYITs6VI592mpNObVWB7qxGphM1g9G/Jvc
DC1Y0qMqakAG8o2orwDeqZZxxkjITzpJzhwJWtbyZCebWpddF9/knOeHxTZI
KdlQEJTCA5lYKf3lnnp0fNjvIBOMfh1lE5rrOcJ2qqui2pg395C0rOr0t/9B
pLIpdnc4yyd8O7jvhwkfTYlH7lfua7rL49seb9VMxdpQDC0TAhF9XOWbGxrR
kOxRPMpbfz/qEPAr1JwapytgDTLinfhBTHB66GpXVaPwrNHZ5YGTKQJAe7gh
zt7KBAttm6NrJBZyHr/Sm6DJT6JTS1fOgzMWRmPiO//kBbp+Lw5ZWKfyb+qq
Aywog6KJlrwD+V+Dy8JBPKippNBuWc/zCYdBfdqtjznMar1nETwV//rqCaz3
BouvNs2zp0/hPH6UnflJjGjtxAoPhr1KL5sXxoOpNSM75U3KsnpojFMbTLsU
2wa4oMihOnGY9HAOgHFvZubZdEDVLhkOoNA3R3acb7stQLchwyzcjTUGrMgN
sUQD9Yc4A8KVwi0RKPkrEd8lH+uUhTPqWmTumHZBGoozqydhx/DgrxxKQdjC
LNTpjQI6xMsaSwjNuSjGOwmpDvWfab4+trk7IRvScyRd0GVfoeRD3STjddFB
cdJXBs3HeB+XTPAvFmPSlV+/qmi5NrwWJQc1UmpXRVRvYtSdjlcONcZFUv5y
NS1uF1j1rQewKBF+cL8MdfgWRZtjRXv/tikEr/cFBffH0wyAWSJ+LLRQaWo6
JHsLvo4XbcIqaLCZKk0WqN+wq8CvaFMk6HyhhsAVN+xHwwuFL4sWRvc6C9pJ
748kWuEUM7Bmx6qR3IN2QBvcnAKGskqg3mqv6GVa8EK/kRabB9W/I+AQgee4
U6TGH9Owqf8hRSQwHm7GXR9latgb9/kXH9sRgRHkmZsRyH1Z1sp5b/+s/VOX
tcGapAfHOcFTjYsxYfAP2DyGEroecno6zy1P2FD6cNtSh/13lej9dxyz9mhO
YAit7Ws0SLT7LUJ7UjeCcNhcyydcQcajRgy/f5TxT0YPT6t2vYLJB4240tk4
176PnhFGc1HLOmyqCCOl/IqNFJQJDHjmj/n2gdfo7hmVSSgwvizeH4A65vQp
G0Z5W3/MY1Mxirn5T+UaAGa6Eriw08yqMe4uNh++9j6tLvt8Jp3rPaV/kS2Z
tzWs84FarUWzEdjbVPTeSLLGdkPJcK4IMG8L2FeGHBKijfQLHSUfh6R/N672
iUv8k/oNTH/U7iUaaItEvYiIvQw/CFuAKEhidg3YRBjdkWR2cxPgNVx42Huj
QJYpXis4zIYEcN5CYR6WlTGuvMaeHbU3omhHECqQDPnGbkuEPApImXre3+AA
Fkg7C80qSuoMVPlJf9r2KmbDIfLSUvyM0B/woFu1Gqo+6UA1lK1At8oFjb//
sZDVcIIts3jJQI7epjlyHuRpAO8rmx0lJmfUKfwbYvOO2bOW/2Tc/EZJJXJZ
6+rUfE2LxswH3M19EYEgon/T0vy+2bRoAs6J5HbzjQaF+50/ph1+C7mOFQNG
ZXl716zoIEZJIt8eHZEl3/S22c8f/uskFmKLCKc8325M3nXPLkw9WTChMcA9
wA4cjc3398IIRf0Wwh8yK1i6fSJDLbUGCyvnxODXA2saoNSaXb127Z8E7/AV
Ye1FC8c86muvCOAgTO8UEG2A6d/CNepWkz1o/XHdzo/xZs7ElTygIneoR2eZ
VcT+/nB9KkH65wcmXwjmGytFoIQbv108rGKpjGM+vWHHypmK1pdHHVxfN+7I
VmbxhW6y+mtJTgYbTJDC8tUOq6G4RC0PR9alfOaAPHgyK7vD96hc0z4W/1Ks
yK+0EMU+BHTX+AF4umOo69J3/KuFjGQBJdGQsoZjLDQjBt3WkvGvAWTluwtb
yM5CdscK2eLHMLYQggXbT7WJQZ5PbyPyNVDVNHRX/WzwQJMn8ub9Onghbm/R
NAj1S5mbUUp+Y0n8JdBES5Dkx2zvNywKM/N8FQ2swpFv3iBe1tfCuwENslTh
JJ08UOjp9QR0l99MxYRr1uvU6/FGHwsdpIKUyodb7zLUczegPF2YfukQMSRs
qNzxI4zLo+Sd2Y9L52x59rN3ldxoGRtlqfhxy/SscoLjSTwugx1FxdzT5HiH
RpLfyfQlgK6S75Czg/V/jpXgQPoCHGB8TDN58JFP/spvSrzIMYLQLGxOjDhr
BsX8d3WSDRlnn9IcR7uqv9fZ3+B0qdq3QehfkBCam31+Cf3cx4h5l6etvuo6
zjddhpeUm84IofSSKk6U9za2zL7v5c+Vy7sezhYV8/RRJeUilGBBKlITrAMp
1XvUyYr58eNQT3LdgLowcWwj4Djlu+hU+6CGoz6U4idOAz5LXUKjq0Fp4ThN
leE7Vg29ynPx+HlU2cW+IyiOadxOJ4+NeLGdWQ2ZqelnTucns2TZCoiSfChY
gi0t3v3VaOLyVnB5pOVJEXHnLt5ygOm7npdhGAaytJI+9xowzG9pPkY09c5f
jWdEx37UxZJ2lsgC8xS6g2dBPc4coj91LG+TWjh+MJROjIGQL2pDlPRZkAKU
C0M6KK9I8Fpt/1h287qf0ukxnqUje5pS2o/wYfzOa8drbJMP7bmz29nLGxuM
J10WxcH7Z5ahnz0o/xO/FSAVq4iUDl7OnoFxGxBACGWZjuAuHew1g77BgX4v
AOD+MY/2OzHi2i+UtPxyglVWpKqPnIx1nsTfHoMiVugqcPISYZXf/6zwMzcc
dWq0+F1xplnAnTYUP1LLODaaIFylR+72dSsShHpauwCXR3bNjmdYEUm3MiQt
oIC2ok4wRDZ5FsJSvdm3XHqtoIgwL9QlMwjgzSXzsCpRwpfgCqAEEnL13tCg
Nk17OFs7ZwEl+/FzdeUP51Ltgir9xWqZhhVMFy26VBd486nwlSjmVwDDviTU
oToopHiJRN4ub6DlzpZXeexJseTqa5F/KU1L2K557Xpopm4Sl9WW2reMJkxO
nR8Zcez8PRa/rAgh04uPsNWkxJczPARcXflCMCDXkwJjEPuf8T3XcQWYmKZv
TymzyL9UlzyY+8gxIbaKN1VBPy71tbav6gOVXqgJOnwXmBpIx+aURYL22VQF
xN2qPnPtfvYfVBWQFQge848tlhCJT6r1XAhg/fvN0l9RDTc+r8FJ6xjXtpA5
EzG9AP7P9OGKvUcQn3ckTaIjJv2rsKMGFnBODl/+V/4NJDAYLVt3R/QOl3vI
/4mkgCg7+2Iy5FovdqVrWc7F7OhgXc2R2nqmv99w31dIEX4O7Yy30QM6lsF5
yRyoSMW7584fTDMN9oxMk37HJr5NSXUU7d6hKLN3vPM/ENTtX4nn/3nmC08O
mVfssSE+5S0HAGSsBAu65+stmfvZ8JIADfN6zPnbG/hkS5CSZK7PG88PwdIE
YErMzFAu+auEog2dviTubpZu9jqkkNErd8pQO73udMmptQsB9faRhjL6LwVz
47ZawNE5P5FZijteTAFL+f2WPcJoh4eZFbOcAznNB3fatSZW7ctwULY0MY7M
KMFfebu1i187Ekei00C8kkBcNiw+wb3d7cFlrMAnPxcBe6SBnhTy5NDuKoU+
84nFcxz7rpPYiM6AJyGygE4erH0fVyWjWpdB8/icIYMK4dJV7z6K5McGnDfh
HEL+WGD7DV2XWayVMEIK32L4NBf8g7icJpB3KarZ8N8AkVlb08aI8FAs0htK
syRY/OFL9qJ1WzPMc0pLsR2p+dD3M816GOVhxFMX9q5c5OkUhAQtZuTyxqAg
3l6dsW5fPEJSPN7ZyeM3O0ZvqBNtZKPVoWZRUTbGNEl9FnAElWHIg96F2Kbm
ByZqOp1l53PSw2mdntuHLm+lBc34k5uGHLOQNdc92A+z4bPoajYGHxX1i4s/
oDFMwDkmlTVgooaopWhJEoXjzj8T5WfkhkAiEFYLu9UeqpzUPdhJGQZj0Lte
sJ3kkbXM3nFR/2feJBpAu62EJy7Gq/5f1z0Hw76REdUmt4d8+70aYjjQq+W1
JIvchQscl0YFKPQ6ICTytUSkRxbvaXmPU5v165szRVwqb9bRgXpJQhAJ5P6f
j83UA65ELZfQXiJERqUafUYFKZqM2cnYF7rKz2DYMSW8hiWbP6w3BEp95RTH
F24Mp8502Hiwecq59cCV6YjP+xUqEl2/qGqlZFgrJb372Up5cKbIjKOpQjYk
C9WJYZefXRCWtEoglFtzfZYHmy5hfPfbwXeYigrTQZyWyc1nJQ4Namr39Tc9
injlE3AuNy2y9uWLK3fbubPynpTYNMlVXdR7p0ea4B8nSFHTNgslPsZAII/Y
6ELUWO+sZ8YJ1BaGazrW0aNNrQBNw/tp1HniIyOHPhKJBripkoUSCBfso4Ae
IMUXm687CYvwCncxgESZM2LZCmDvGEbqDHN0oyifWjONoxQPt0Ongh7Xg6jb
HX2wQ7MYFAW04j5/vwdXgdecJn6qyyLrmxy7cgaiSOgPPyFQFYZ5NBVqX/Rm
Qlhd/B5nzAa+6pcPk1GSnaG+Csxfk5cxTGHCFtlI0h/bBRdV9gADUSOMNDUA
XhXKSEM44HX6AX3l+vezSijqHsSVWgY6el5MRmL/tBv3fvCrOlX2/Z42ow03
5AdBwrDNxP9LqVeM1FljoclfBjv6fcCI6FOBy7VkoqmNwkqB5kfBUhBrj+qe
9060rXncamSyCIASfXv9lB9BbJqb1iMAugstjlor5oLujC6Tj0h4LffpyLtA
cWoOG/NzpmYQYQ8f6L+r/QgzQbCd08SiBdo2YlxV+AKla9S3+paFEepzytPe
1fh2BdJh9mAlEJrRllknY7r75i8fFSEjo6RtTy9NtIXdpuPJzC0oHNRgwtHO
S9rtqmgcROvC9tdn0n7mMrXwiRgaoFkW8rbfratTE45a10NeyfGpOxyfZ4Cg
Q5/+CAo1o0pOV58EzMLql5SqoSlqScnBHjjhGxPJL5F8wpvY1OeIaHyljmVt
ZipYrbGV4pUrUVQkCiut8bd/b/OB+PA2dz6r9pgH0FMFHFhxk8bJ0d6u+9cI
W5j9DKK/ycPCYF3LdR5PvaPAJneh48Hud7trjFf2IG0WT6Wo+BtdQPf146dr
RU6Sqc8t8d89MiYGbIfC0OA1EiAigg7PSklvKL3wImzwvVd7F7yeNP1Cz/hP
GN4VpZvLe5b90n3wg3LUfgdv+Mb4qe+yEUd3Dlm9t6r+fLxXyjAaVBJmJGhm
BWXgD5vLs0U9phODHszFfhA4TBSDXq06SEmiHrG/8rxl50g3pvQZvrZDeYO4
BfJ+kQ9GXJip8K1n1+VRBHuCZqbMI/VXsPGI4tnRkBRhvX5BGVpu6K/yoOWK
AAWCzppaq5FCvXPFRKQYz30ToQMavjn5RQ7SlxtMhvZsxHmUQOyNaY5YzOAM
8OGJuQd3+2NRBpacumIk9Fge7sduzS8oOa8dCXWHBA8LkXxEKtoN69Ei9xvk
C6hzLRTyPi0SW+7v7vSC2ZHgbYU5p5psH7aUDyqCWRlIp6D6qNe2RQRMFLq9
grzzvTHwhdw6JYNjDgifVxtGaR60S3vTWZMx/Y3p+S5u/0HGsuaX35Shq7EB
gaP4aBrj8VwL1vY9d76dOOBCLJOynb6WStZZxD7jZtHIirHh08Hg9ou9sJ4V
lJbW1Lbx4KQ81Tyu+zDQN3b2HuiW2jI4QLYwUZvzgmveUl8wwCGGcK4u5C/P
4RmiJEe8xVfW0pMhd8Jp/ut9Vnwh0dEb245nAXMdby4i7onmhdintaKy4XJq
02YNbGn5f56NDiLbNQlycH4p5VZacjoyymfU/LPxoClNGapSeHP1gPBudbAX
KmWbDpXpwrZXh94Ynl+PL0w4IVWHME8I63gNXJv/kzC7DPfpm/w3iRmJaSbD
xpTE1Np/+Uq2TqccpqaU9zU3KfCqxvvTtuKX0N4tGKTWCTiVd0PWpPEZYhOO
1z647X2R4JtJ7qJKXpjCx5pLIRAlWAgVvffTM/GeTl3wNSFGGEyMNnAwUcHZ
DlfEq0t4JxcD9FtPbEjsnz4qm3jlV4cyd8r/oEN5TQgYjyYUW/8ntM8QEWgs
oxAyjuVn6FAUq6QIqW0E7BESGRZClXeG451wnKNcg0grfpq7BXT6pQAAhCVt
AU0iiFqa+m1WRlkbirfIpGnWdCeRqfwOKdsPG1WmLy8jeCG7M1luF/FNHhHS
d4ICVoPps4t+lzWqUJ40pR79nNdQi+maN0mkOn7jisMZmsuVa+VDIDxQmG7F
ASzdni6djYcgKrUO3o9Q+K9dOCSPnCpQetLUB1ho3ULqIywiXvZFFfpc+OeL
qnJ0t1LHGQNRn1V6VEpknUYU0jUnXCtyucj/LojlD7T1SqKkrT001S7LQcHf
QE2W3WdKuEy8TqsXBZr+nhkuHWoiap3L+NWxzRHCXYdLvOFsSR+NEKJW+GBe
/mC+IxxKF5oHq5su1gfCH9jV+Jqf85wsxGADu9liLGT4ym+xnAfxkEVmOjeS
tCZQlmZEzVOahOBOW+53tk/FbD2yAWYid+oCC50MxMZuSNNQrG0Ifx2vUryV
/Uek+7Em4BO7celi1139SHeKJKypCxETcfnEzyVuEIV/GVBdG4GolielwjE4
hvB4cbLVxfumdIyVfUyKAmXB1DzsYCuavuNPPepV2sHOl/xbUTYzxfwGbWnc
5CDiKZep3HUyYma9aNkW2euZLUUHkgKmSH+/0pM0Y3xkHBxzoo05ZfQN2KSf
1OCjrNMOHqxwNIR6rywnCAOnWyW4Ut5f1nGF0a/qRj16gMAHVt8dYpLLpOy1
GKVFz4e5LNYbeICwsKyyosUc9XXDEMuxfkIfF6xAhO36dfwFE9LAgncDF9XH
Mg6qwpCAhALfxD9T054hZpfZa7+YF+GX3eHQKlgS9LxCAHnfbJu+TtyO/0kz
JxnR2ERzvFyNBOhteKHWdaUeutGt1aEIv2dv5lMM4qZ20zm6usz6M6iLdxG3
mU7VlwhQ17pVqJZVARuCbDgh9gvu+fz+lDBjL+e7HSGDGaT72sctS7BcplE8
HJqg93OPoqQv1iLA2lg9qAMwiEQ/6jTYnAEJFfxis6x+rlFlReTpnx0O7sWl
fypDVPI4TtUECMKlpy5RFe0W53Gkaz4/PHUjoA16UK5XjVdI9NW8JR/0p8Di
fO+AqgEdVlvOJFmITjcGSKgUm87Dr7TMy22bpxeTgGkCasMR2TYbJ2KVZUSM
IHltlYv7nDyAtIHCcCcuLjQ8Qz1k9qMUbx/NGoenxWls7TwJzRjGYREdB3JR
oQWCG+iWTn66iq0x9xNqSNG4YScfxicPfaFvKqW1Bt3nmSrFz0ONNR5sJsld
FG8Sk+ZL24aq7dwzvVcW1vRx4ue8GWMc5nSuRxO4+QHGKZaZbeInCBcwHrca
RptniTINCbAglbRQrAI/8J1TWaTJARg/uHoSRTyMckXMLMS5ss6i+3/T6UKX
oosrXF6ndd20LLPAaoIAUKgMZRSU//uM7J4f+nj7WhFw6Gzg+PJ1ThbitNME
zHNoPsNBuMDmDvOQBdseP3cq8s36hmiGFBDzrBzl8uCeb0xfHNSPih6GZAQB
QEYV2Icgrq28y7xYELFHdzvCaY71UUt0Zc0ELwmWCz50eTo+CKk0OyDKdLd/
Kg67LcWW+RPCfxqorfAaszOY/4KSqgK/wY/aeGc7SagkN9ZJtchoSw0RS3Iq
oTQd/U+2v5nRBYgSlVqQHvQNRzZZaTfKaw4pxFbbxrwKg4gk18p4depmQ3e8
gOQBkKXWfwgh5cqP1oKNkKYfWbhfOvtRdc0ii+zcuvnSTCoAfz/Lckum0zZr
RODMGfooTi1Mcvw4sXiDx7qKJj9Ww/dKO9Wxef/hULuJNedfe7MxIf98ekgR
N8whBPQ1vHBvpSeyJl5QEr8SszkjtPSS2d5oQI3GtHdksMlDyydeg4dMZFMJ
UM4epdgUCaFKBYvvpjDN8OzGDDtZMYJpuMPoxRi8W3UOsNGZ8S5pwN/yT200
XLhDEbZYrjTvXMdP0rGdNfA/MrbutXTjodqpFNax75B7TtNVekYNmaa8CPzK
B2Oh20yNMGFywIzoz1zNCga7uoQ+o3qhJ71jMmfoOj+iq9nzn77EQT8yPtH+
YRlheOb0CHdG6yNB0Zarw50u/NkVGGPys3XDECldkZFLrAogVv5PUbgiWkjR
aMCEdJomWiB6PsWqhMHDJL95NnDG5BIPjAODQAg/dUtyCC8CC+x8qg+uuWZ9
LguIywObtrlKg3jvYeVnRKWrxantfvXChJb11jVkaJvmvEMTxmbyI2IFaahv
bVKu4dGO2Z059HCzqotUX5IDmk0klEZ8mLvvURqTyQt+Sj9MPHKMVjxGrKgp
R/xbcgOL7XdbZ3JcRltKPcI8Ij5ILNmnsZCmSHBL7Uwb6r6ZhOASqD+CxAl2
hTBRi6L5KzxRHNhMrDZVbX5yft3yMT6W0lz34cOiSVx1f9Kd6vRdguJRL38+
lFZ/bDzz+yCUHcEfqKcffK/Q9OMWrheOR8xU4ODKiH+T6ec+/XYQf2cM+41c
3/Xslu3MVZw+mFsJgw6v8eHc3cmPHcYT3FahYBxp2LIOd+maTrdyph8is6/6
q6YeX3EGb7dpbifm77K1ciNRJpvgY5KYqYEfK15Nh3w5H0fz2x93skPBniuU
MfAV+IFBoorjm+1I3z3gl6veifRE85209WX1jc+UgrfM1rrnII5CrpjJxVPE
T6AWzYsnROslJyZcFnLHQF3KHEx+K5G6k6PCnEKrVW4S3STwWp53L7NlncnE
CCdQ+C1rXmSCEHnuUi/31Ay1obsWQP7wJgU49QVe4zsOkdLRrbe2WrUb4rLf
TCv4Y45ZE0kgoYioWdVoxLYf27sGzWU1uNYG8/vvJA+8XeN8LSExW+BP3ImU
Zf1aPCPoUxSP7tqdwep9zP4wUaeg6b4nOS9Y5j70FSssLQAaDYf6Fbn8VTAq
EvfWsKnRa0O533AD5cxPeyLKAjTSMas6TXEuLYZtNwGpDDLY4/L4Au9jKJ/W
3rYdD5KO+xmoUW+6TU2lybiGoh8GSFi0yYFKbq4hkyUvYOhpZ6v84449w8Ay
CoZ9TjoiUDd9Y6MTk0BcnpZIk8iQGzpopJm2G2qSmv8Ex9qoZRHZdzJwhxRL
I/4lejeapOUsdOdXs6+Cxmh60vajS0Ct1rGU0B7Oq2vRrE3FwkCaFEI0rSS0
k5XtUnSJ5EHg8E2FoNJoqXVGKxZq4DfOxumxeuzqclVIFDrP4bAkWoFCVE51
vWMnPNqeX3OUab1G/ys5q8tTMvkW17xTTiWMAVjTlwNeXtlAQ2R5tKLc+VxD
W0uiCb6yCfTsUW6P8IcwzcBMzbDfHK8zNnPwVAqsWvxmHIkHneIs+6/ue5fw
h+HgTEmvteZquauQcJo/FzKdvZymcGjugpoltzwxKjd6+0je9/UrIDNF7iqy
RUBuxvGFphJWdsl7QrvrU7+z23shk/R/91E0Fu2jl2HmmFaHA6Zu0rAdkWaW
wkEQjX1dnDfVK9JXqmXOAhvlZsDjMc+4wCb7Osw/gs1n49cVg6C1ESpEOQLY
SxvaxDlCP7/y8z6Zn4nfoJEzqFqL+75m6sa5KB9ydLYFuU7XPQuX+TRvqXQP
tgYdh4V+PTMTfUGriZO+oeQI/LdlIRpXfXIxIRMa+/hOCThHATdzqWoS/WoO
iTwtSuSU7bqTWis2uQ6JF1cMCVRWz/TQNTaNwLiP5+p7pNI8ISST0zA73SX8
3OczTWXhOPYvPCjiQN0SIsNqEY5h61yTSfrLJW0n9ZPFfYbwl7cToMQIT+8O
NEGZ6V+tSdTFxHFZXaCOI9vlYOinxtP5Q+uLXUiaCJCbUIrR+1hVZF7Rdazm
bxmTlpQphbt9OU3MMpi5Puhietyg5TBtzsWHb+WO2c9jgCCLioCKcK8DV2E2
e3Ma4YXIqn7r+tr8TEnYGWi/KGMNI5Ty+nDT/oMxWQ9ypb1QtVqt//9nOZwt
w27yHpNvFNeagkwXlE3aCA91QM3lwMWZOfiBIy/Zf/YJrft6L87LHXRMlLek
Fw6Hs2lFi915w3xrWMjN/5UFp4Rqdyvj7JsZ5lWMW1LMqmgbxLLkLI+hpU9u
UKS+RwgdaMmJsxW8gAZB9Tw67DX9sTXvj6v6qOFEbzkVthOttQr83ydbbTEj
XANX1eNbYr+W6YdmO1EdTPtjKmESXhVv7AXgFUdY+G5iAds0IChd53yEQXX+
dUG+QTdTl8o5nxYoW96m22zSfccCTq9CZqC57gA/j5hwCC8q/ASU61vzBL+G
bCopTwWn9NQSfVlhhquYZK0ayePn

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTzhVU9rYlzgrhAZpcJTCL9snUTQNuOJGAuIS2sPpf3wCQy3VHJ6R+Jg6weu8kbWUUW493BShCVAbg7gezywU0nR8EWCIRQC75Uwe+KCvoDIa/4f+MmoIQ24w9dVKVVYj0d0rEh05iNcIuj4iBhMw0IuENqBz+0oRml1eiSQt7egifn8CrDdxEtl/qeUlH4TJZ9P7Y1dr5hm8267feIZ2Xs0V90O/SdCs8A732rLiwvNxobr1l3sCKtyjk6wnAGThsDf5xwRHwwnyUPyv/ISeHslQQLLE4eNa0902CFbUAJQHEklkCbGtwzh8iaZcypS10O4hfVjnbuFFYBTFAHYttC9tZC3O9PaP8oYw+MUb+jkET9mXvnOs3nQ7hf2UT7+J/h1+GU3JzvXcpZgyg64P1qK+l4eyT12w0o7GKiaQJeBJwYLA4Prd06nI9kY5is0nA45I9VCYRzHTufTs4YTSodk+sy9ll6tEYNfTQ3u30xBVddMdnJWP/btIBcOr6nrYm46tznVQ46oxuaeH102AVDY/PMj8Hc8dg1BlkB2TCECOA8D2TuNmdAq4NTF1QNaAJ8jscOTUs9YILL5Yxpzq5ufOr/w0NaW9l1GFu+3HR4BQQNSDTa+j86XPa6itb4uEA5KpYjfG//n9mYvdvOpiCAhIwdb7fEjJ3CTdncPlHasXQ0bOkznoGt4lCB+WtKggXaRwEq726rWRkIpMxxdSObwP6RuOkKRbW+uLMdYZtmjY78+Kn1H6EyjFnXK6xnGQsYEAoo5PoiM+uVeRErV4Ka"
`endif