// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PYFNLx3z1o5mig80to/VkKLraBhwFdt/l8SlWEF02QgqlnHdKGob9XCVVSsd
mxm+9ltj4cfdGh3PW5slfpR8wMfl9r7+sWk4tOvjX45flAel5YFMkge7AwlM
+BJN96KXOYl6ZMbkU97HinfmSmTFo48SPezzQanDM+yd1lAIYiBZtPN4q8mz
dUvQvPPgGGGOHLorZXAVk7Bw4e+ofXwNtx4kF1dlshJDVjC00EMK+Xp6Jg1I
4hjEsSKw/3UDmsxp/8vbhqJedYfkKOgwNizhykuxBUMwYQbuMjohagEtCf8l
BBdC/HFBupEOJs93iNSYbX0TNXnbW5t2wBe4hmuDVA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UGR8YDSO9gMm6FMpZYmckHW+6TDsOKekaKWUnADHYK9OYvZ3UMLs2HYuwpjP
4qhII+HtmEbMPxvdvzera2xTWp8hzIbFwaYyAmjY5UQMvFo2BsfHOD4bsjUp
aNRru+HwdLUGqBra5p7/jZ7bIIMymcz94d5FxdEuoYFgDINTeB3IQdRfh+WN
9bN+CkYbY8cr/AVdhQd97W3L72XBno40qHteylV55MTBD0trJOotnFVjhski
aL/TbyulUuOm448AZcpKmP77h6Goygv2KhYA7fGeAENBodtmQsbfqPP9kKQK
uHYQKT9IU4d3o+e/qCZ0Dbo+Rtb2QTAfelwYTHL0XQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Erj6/MAbLSEUbNyiBg7TKd7yIJQC2LF3TSCzJ107ysMNyfi/cMl34CTWyL2W
o0Nu2nT2mO5iygegqeLeQMS0x7n1UAkGD0QtTatP19vvKDehEh58ljb3jiY5
0fggtVQVUIUuKxRARSWXJUSzztQ18imkTTRs+MZYVD5L3Vf93Tb0IJbTgnM3
LiRzmuj/MZLLWN5fPDBK58z4piB3WJkjC44YrG5eA+cjw725PTxvoo9gX8XC
wq1409V52RvvKbSiEJrvMX6LCpcpWZJG9HEAfckRRR247dG8ZALf6Ua87cwR
Wzxnee+H+X2q+It5UeYaMt1g4Tr/P5HRLbxVnvjUIw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EtYvmz7iEdY3B1jdR8obBYm9OS224tDgjyxyXO/kP3aO//FgtRUOcw5MpJi+
lVG1m3NrWM89uwDmgITGPEIAyKoL15AIVcBniKuz5iOvaotsJ+9pXS+G82vW
B34d6hrlxB+/U7MRmTa85lA/Q7O9mxplROPSjriacrwR3zc7UR/0GShkNfIm
nbpmkBU11+XyXqvOPdTp67q+YKZLz7D0LxqoU3lVTd2UefWBcV2GEs/08Osh
52VMEu3fQm81Z9odxrQUhnl0SSl8ORaz9pvRa4P0+YhpxUNqG2bb0zFbWpsh
gZ0fl1UbnrGT046yNAhGFdFqe2cYdYSeDZG9nAOZGA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KgRdGuWrn4lGxMyOQYg8D19aTvBJpcMmOfLM+gfAUZyV6oWOgP25JWJ+InPN
Gm1WaguiThVVuJkk27jlhgA14Ml79GeSqYMCyeOfo74Fx1mb7VDSGnwaGqDG
WZLoBWsGe4+ScELYeU9oFHevSy9/A0sh4EHpdeBflnvCXqMer0A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hemEqhnnSzlwDfLquqbd1DhXvfG8nUAmyErfr5CbfKfZ315iaGFFHdr3swpH
fyAiis5KgvrhJDwDE84gHabvs3DWafDXOpbRTXsOjEv1Fp+t8nCdN6jT3DiR
tBtYG/Es62QdydzRj1XuEa6qoIq2hl2q3MCzdnUbCKYUmuy6f7ZaSkE0lqAU
dgmRgNxNddK5eEuCi2kpy50uzNGiNvnRFVertZVG6Lw5vetWib4NOgnfUdnk
JhH3n9v/hBuFH+1IdQc0FhHe5H8zTAm1GmVhOme+SDIbganCSQgMP3hCQ0FX
y9BGHwyp1rYBWsC4pSULg2dc8Vgc+vr4yJiTtdovrl6BGp6eJY1L9b32cANR
bMgYnfufTK8jWgGzjNXbomuKuYkX3GCiq51ZeEi0IUuuLhTJXUhuVw5MVqar
YEwGbznnyY0PGJrWDWwJ3JPFvTTaJj+uyggChzIoU7npo8L1PDFREW7WvqB+
39Du06mecFcyk6V8OAKSqigwhnhdJ43z


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O9vUhzJg6OgyhOkSD6MCys+DZppRADF7mtLGiMsP1YOf+y5021ibuxWyQHLO
Knk6xbJnQM1HGHc21T5sstuYb7YPiD8rD/myPTczFusg/AMJ5lqyTmKZOdHU
TxY3+b895csJKmMD7kklnOEpZN8F+WUTJ+PdLWL9Lyglc+4oO58=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CwiDZEKc1q8F39WJF//y6UMNYZm3uPt010780YnWN5lryAP5WfV1U2N+qTP7
LfCQwK0arfhjyOTe9kbX5DMp1crKxXTsdtohgLWo0DAr8YYwg94+f50z+COW
bSGBzjy5lMh/I1N/LmHZc6gHrVT6IFaC4LbPLjRbB+EVOkHwQfU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1008)
`pragma protect data_block
GD4otqeq2QrmBPXA+OMWYQrBvMKRJmHHbhQIaYDkYtgQdFVn1IvKHW4v9lI5
7+sY7ZtkGYUuL1Mts0UpsxkDOQl2/TMaXjo6/NjYv34Cfj2TXg70aKONKL1B
0szZjSPrM2Rib3UtSxe/BgsTrzLVZenKCLYQjbfzU1UpX5UCk70Y+xwbJk0H
3clwlY2uMX29F6oLjBfDV3SuhN9gB04le1JbTCzv7jEBiLWyn8sM/r4v4W4+
TnZYOb2Pr+eOjqqTS9gkyZjTROD/KzFzcHzMhoqwIDdc/yN52/555rHJFvfq
L7C7PMRDgWn9qXupVmYnY4OVbeS7PegXny6n5fay1p9iEXczimZBYSJJlQiJ
rg2H+LGM0tcNeSMbCusTzUPdeLdjHioSUrsCUV8H6ULzF1qU/fre0+GbR2m7
5YQpSduRxvV1a2LqW9ss9AP91aBrrdRQt2UW6OL/tzhOmsaYkFSCch4pcaUq
TTE3Amo+1mkMz0mSS1KojeRMDmjOG7zIVArmv39iSb/F9gAxp7zYSobhbBbT
Po02TKyWv3fixNcGeLYeJOo+hpy48s0qKcmfRXAErs/1odsCWkBh4VjygtCm
PYmOMpQeZiW/scHIST4PcWO2LYzgjrRaA1baSlJRJikMV1iBc8VkFimBaafO
+YKt23Z6iAhD0mH6JzjxbZGeOdDcvARv7pfaA4TV6BbTzKWh4Rapdg2kNsEy
XuApJJgswzoF9eHtg3P/nU4cJ225yWxgYBNzwJVr80EHb7V7nfkLOs1/mm48
Hl5UcqNnUzhzEeYCO9hBaP3vD2+HellTx778/05yV8HGtnXW476poJFW89P2
+vcnWDL8e4hwHrG4XU4LNS50m2CYoGe6PjtBT/Wh1tYh5McqAzONMnrhqAw1
sIY2W1cQv1UFTXimmDmi+qjiAwcq7RxGfToCq6Zi9YpyOfGRXOW3BY2qDK+5
Vj8A3oK/9f+SgDkuE3DTJZQN55oTphGar6E0Qr2/G3Hgj7+CFSYaAYQtZf9b
eE5jdvgJhYYKmF/4z7TPAAzw6pctjHzWPQCCoKAhDFdKVyrA92Bc1gPMlM8v
chg5ztCuOGOkh1rv1J1BloeTl5TOYWcQmxjvdKfAfji6tYJV5I7USixVPOj6
oalDSo9Xt3slHRvBojeXvjeHlrQ/a5GEabAl3wJrKetbxZWoaujlZjC1UT3Y
nzKoqqcEMSgA88pfLxI2IR+WS5XoQSgGOxzjk+2ClJn/2F0EMjCPBsdelO53
sc3u1+9aY0r71NuOTa81sUfZz29jM5UVwE27uxCyUmHxIOlG7SgaYKajuX55
joGDrGQ1KwrsRQAGzel80Dx2

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfaOIM5x6N6R4ckEuyI1Fm4rYyVQoPpmXorWP6Z416Aps7NiLeFuUGHJC8mCvW/xX8o3oGPezj+Hxu0bo7vOl5v3p4cd4payFR730Dn/B0vY7CEPof8mPc3TCg2XlZu9C5ZA4Lzx8PrHuZoTu17vElauqplozGvcLwWg3b83KeRYqPOO3YfD9PXYXQ/BYW54pJqmOW98IpkzbSnXV1LPDogiuKfHcCWy65Tss5skNHRt1mK8sBAmrc349+jSSnvHBiqzliwnrS8X8ttRU1zAHhcR9M/ltQKn0kurCw2vxv6iSsFjSlho+KfMULbXkkYH3KiU8sNcgXRWwWRnV8gybdabKkmrfLH0AhoN1Dx+7BexPwH5gJUokGeKRuFPC3FTqtlffk+vkVlO8Je8rAl/ikl7QicVqfMqjfY/cN94Qwceb/Hhd9fNCj7HRtLALbMVaQWeNjBoXqqZ+r0U8kcRE30ChzdDDSyfhy18dRRZdVBS7NfxGcoaGtd43y3L6qq+EL0vb8TbHhAj6hLzhQs4l6U7Bg+fZkC3vMVMr4vjPdHGh4W2j8qr9Ct3QcqQeoSLPouWLPNSawrHOgO567Fay+rqp76Frd1/WxlYMmYSpWYz4a7+uakbyH8guiORp6vQPel29cs5h0tpe2dsXxL8/ymAjOYLprbEhZyG3xGLEFN/EMGSC59rcmu/YttYWQUd1PaRz8t2LV+JcNLHoVxfctKwk1FaHEbaoIsiL9KIWtb4yuAUrE0O4XPYNSiv529ayEqUfjwjVz0qvG2HmITfBbi"
`endif