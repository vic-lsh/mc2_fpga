// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jPVemM1D3PWt7UStvDb0CTDUOaB9IPfleAzBwma7fNAv3Lz+Uf5SXK6DlQHo
/iU0cS/lya9rglBgVAGRkttjTzYxkgwWD93mVz86jXS7IUCqBx7MZLgk4QGr
m0wwQxS0RbbIhBvIHN1r+5munbfx6qGGu/Hf9FIrNHUTP+SnlckbubdriCHy
9iJjRqJIL8z9UUOggcmnCCQp0nQt0xqQuAiIgiSDQgtS2GyczhxRFcC6lfta
9ZY8ibJUQwLI4kYtAqHUZ8mhUix+gwXmbrixrg52en6s6IMUIaMFygTDTNrJ
Rgc4gs+Vh7q7bbJG/DlCNMd4dlJe4H24pr1qG5qgEA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dNCKV4cZoLwVfBh/6Y8ebqJ3bKar4uj/pId6eJ3nwNKm8UMUS5Brvoi8f7g+
oPXaNPMkuqgwW813kdiNstoCNMFQBHxySvlKJMWqVDdTQr5JwoGJwlib8dGD
qPnxYc9mOQhFn7oNBF9biHNJHCZFs1QuiKngFXBjrGBELe5YYp15E1IwOaXu
HuuAomsYxWpmaqQyTwIkHzq/Qc+se+EOm85AjDbWp2bnDBSItcmaERlcckEh
9gA6d9GB1nGqpWmsUjlK6Th/U4SPoJg+GW2hX+8bPYuV6aBi1kHIgvMYS3/6
jADpd4FETc09LB3yfP1NX2ohn8a0pgxKL58VJ3r5JA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
idG8lxMPov9V/HKmEg1MhiMnvqO2mLv737d8wQhT6R2KoBaDbwLtZLiy6YHl
X/p7f0nf3m2OdbBtJRcBb6tEiiqOa+Khp/jEOaMk0zi9Zc5c98QcvQCGzDR9
rVeE8S0IRxMeZ5P+yyc9IUVKsMH8+o7/Rhnd8XvuheCTeOQw56b936O0Ofu5
font+r5BySoOOq/04m73fRHxttH4H9QZS5pNl2lwKV02W4kX+YF0BBR9FvOt
20zFibM7hu7JIkqpiwtAGpfBjqpARFbiywScZkjCujcoHRJlsEyhp/e1+GDM
AmneQLhg0HZuJA3jfwzv0ySXOUPeXizi7TPfu3Qbfg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jQRuQ8yuJ3FU4cQIfRQHEuIjPd2qm3TfLZx/iuugc+a1Y8e9ic1kXMxPzCZd
wopRAHGiB7bsfWmMPnCOAIQ4vmiUEoHOUOjYZ/V5KP+HPdxBnrQrRk9PBG1j
fV/mHGssVOE9flbWdhRDkV8Z5HjNfws01x7sWoZUZVPn+ZlNh7+J+8XxhEwO
2R+QV/eMJCfQD2OoYbBQ27ml/oESVNaFesj9YzJHw4NU8sL/l0smXJwolfNm
9ihXVQz4Q5cye6C0pVClUiwqxtzQz8TMXQ/qW2Cjm/7ia/uy25u3zVOLVpjv
Qrf9tFBjc28ROnfjLn9UBJ0w7hLahN9DQXGAq7zRfA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LzXLpV+IooxmuuGr4cUUCy/yOeJUXoKpgiYsB6rBAIrbhNa69oZPmz4pZgxw
2FSeLV4EHgfqHdNXeFlpDPjXRYOa7HJegW7phhrH1dPHHWq5E8CvLG/g6lry
QvaDAb6buT6i+/4RLa0UF30XqYe72/mm9zOC9BGH8B8O5rtRifU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
No5lyOk0fLo/ym2CHrh5OHIiKcFlrn1RoUEsKHiJuQzTCD2bByhIjZ/4VLU7
fVVxlM0LnkK9VVFA3HhtDEnETNcOYOc62kKwXpL83DcmTvChCSIcVs1BXOr0
TglEO8/ozl9NumVcIU8tc+cDjG3kDM4Phv9EGqEzttSQ/rOr/I21fTqRtoMu
qAiFcDeALvFrFrSl+CF2VpXaDoUQA8wu8ZZnuuCq+FQCl0mV0UP2ghH86k7n
Tsk+qTT0+m3vgcWLi//MprW36NZN6Y0k+Ip7ke+UG8ImqU4KYHKyZCsR/lvU
FWbSqJSqtdVH/a06/Cnp1tVKpdsZD+v2QlaYezBK+185zsTMN0follJO0xPh
PE7RcyZWsF4HUPWlfsD14lDRq2RAoQRjmvPEl3NXidUMy/GgKcKQX/bSAa5m
on+HlmWWGEIcwxBEdCHgrC2Bjzuie8U2RPc9kj0CkbVKnp3l4jwhHtJqAjeG
sx2udLpLRPOLLfAGoWxAp6TZesq0w/So


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MQTHS6hwyiD3tMhikqPnkKxmmtgLFhcMKhoGYShz5B2kExO9TmagBaFH6j9c
2OFmlf+DT73D92rKlblM7VDYXUV7GRXuThlvTDdyFjmjYGquXb9Q4YGCLw7e
ElrivsaLesTNZW2mphFHGK8IVd5w9fHJhw8XSOI0sHZisXxZDak=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ryE0rtWiZ6X85X18qi2zuohdhSAZve08pgdcObOY23YJ4eqOFBbz2IhpqMpW
MCejixFUPXDTq/nUWjD93ntullss6PpCk08q8FORGqa+m3JSEJYfdhdAS4VO
ScDfbNqDU5DO+M88qwoc0uHUDXgmwTSsHBHIA+wUc/2AwgwVtk8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 79472)
`pragma protect data_block
ZfXYBargEiyu6b5UJ6phFt+xwT6DPDhk6Nc/PUbyyDV0roOr4DxRx51sV7Zo
q9jyl7ZA1tvZm4BP8YgWSyXSX4Alnbg7r0GJutnyhw/1pVdV4g2G2xYBjsWH
YLdFhgDFCRqNL4XXPOSKo0APzhgeitvEKYJaq7rToy6kM3Jh8A0MUsJiusCx
e0qqVPDwF2oonIGGGWj0NAz4pHJIgFNIdEP/C4elRyxvcQZTVdT3iQu3xfdc
zSX2ZFdrsQ9YHL6/ZA1YVCE8vveJ4iQGQfM7EjT0Vh6R07og+2d6dtU3vdVL
aXBy+G9pEK4zZq5Cg572eP7540uT2r3H4tZFJubJNRCjtGW59iiAsRL2VqbM
4Jpiwb16VZx0+Iwi90ogd6XrupDwGZEjU43vFQYwqO5IV8a+iandAImiE18m
sKpXflWxyhU/toguG6bfDif7hdHmfLa8oTabO1t2D4zI/xd6MwaduqsAyJ6a
gPNbhR+9pIJjGYv9qBypsCIJq3mpC4ATsBWICK/4DeA+sODPpK/KLZ/RjBjr
y3/Bj6FUGAjaFkR8+wqUBBuj661PM8ZIU2CqIrJtX+fAsEUZ08sT3XgU/M2U
oW24yMynjtGLL7q/1O388SrXOi2wuymNX+cZSqoSIgRxjgBm+kfFQtCdXPcV
K5cr8HsujWgL+h0W1QecsLQ+u30yfODjB/OBb8lrr37Ckw1r81+nBTORS7U1
2jzHheiYvj85PS1szkyv6XlzB5bTFWqeQEWSahFbPJj1omb9r/baYlFwg0Fp
KSziMXTVl/yHOsB6y2WCjDSbyQaIJuS0Z355QXmHHtuzQ8h+hA3lmpmoGO60
1wT7TrY6P0d4RBSqeclK2LN8rFYVaaoOtf7wkWV7KsG3yd0vWdCKim/tP20y
dlJIRPl35PcKiQAWzrYm2p4Ka7hPAp7mZR9qSUpjtlNjDBrzEIyRFXrzKec3
fiQRE9indvIj06X85kF59+F6XiA4UJNXSfMMpCcj23A0o4tohWonkXvhT5Ll
uj6oIdzk51KLtk8/z4xN/W04+arZcLB0Hy5NNoF0htHlYI0upOz/K88fOKda
WKk9f7F75PXm0m0Glb4ivQiMTkVocLu7TNknrhyUGANZXyMmdYEWr9Cl07RK
mf7+/06ulSU4NK/yMlp1ZsnE8+0C5860HxvUJCpLW00u680c2o4q7VreRNHT
IQ/n+M++BkKzPN4qBFU0LYvlQL1l0SQEbYS6WC0R4xkotNMMp9t9/+1UjKmf
c+rUBlxKeXL9ESLE9601uWrqHXYypza2CZW3+cxdFmgz5SnAKJeycXaIDvXQ
1oMmLW3Iga3odqIN4khUwd8g09A5/0qdEGArGQIp0XI5165zGWDFdzGw0mO1
s+DV5gyHeGQr3ZCCnMZVUR+onq5BMfN44xcwLy6ZQ8iTlI0mDGiPi/kEq6g9
e2WGCf1O02DXImTr1M0mvWJgl4PhYQ1KNbdqGb18uGAFMenS2o4s4GmJZrnP
XvwA8oP/owDXjfBgitt7FgTI+eMQ09P7/jJNcIxMWttn85Aqc76SOg31jLD/
wD8i77WW+nkQaHs6Vk4crgWASoX+IJ0THCGNgT+9XS4051PeXNfoVINk59Bk
Sr60g2rclt5cKY/ZOEO3qdl2qprodS50xfbCE5h5YPpDD6I+i17Rq0t8FU8g
S7qhY9Hxw5iwn91NdUIak2XlG6VoJundwujgYoC5EkRVcbba7ndm3QDO4NKf
60jbRKqHQ8CNYF9ZNPYhr9WyUsK/jEgt2KxKJH5tbk+UC93tKbwv3FcWadWi
jt/0lrlpuW/td+vWID2GcCvm5YUOCXsJJ7jZCXUcFJW34k802U9ZhJk+0zF3
+eKiCy1panm9wC+I39Du/W4Q1BqVPsxG7H6vBTmbe0DJeXAZcpqQjjrrYDH2
lxMaNaDJ7Hi4/75PD5yC0OzP5YdeibQ0n/iVd4Icz0jxdfAQaNN/qKNp63v0
WX+ipm9QRHACxkNPitB9Nz8mE4+MgpJCi+Fyp5GTbbecHoDWrExcIuE490O7
oqEg2XlKvuesUD+hTi+lTediznW/6fTIoCJZqYy2HBPuVHuLQKzO6jFWlx4a
mmW8FLn3JVT9RD9ZX4vGJORcjsQ6R43/EsR9nnrFi0yWFY+R819y3WszFIlz
p7mNWIPW4SOO4rPY/zWLnByYSmVywkgLyy8bpTv3dGRLcEIuGyHE9IdcvDm9
6jWRFyRZcWAwQtdvDVv80DeEs7aCzbXD3mszfkdiJgssrCAQdcTW83QNGxZ1
8F8iAIelXh5ASkHO8nJb9Nv9D81C2RpOQLvuCXnmyrBEzKdRvQgupMVtyyMa
EAWHqHisANOi/kNDmX19Onl3jHeUIzlragPn8wSms7k3nqtbQ4YECqmodG+U
fivIOc8Y6LEWeBzLO3Ca9RS2OOZVQVp5QC9rWEygRMuILbXaGRc4+/DGap18
UqcP1PZir99r5O5QaYlydJdUy0ePWNuAFKoSQgbrgT1ZpfPXScAcJJ1ca1ER
HmypG1YesdM/Lyn9zwJh3Gx3zQVlfL5V4XnkZwC+Gc9BSlQwm4jHaiH3Zdhl
kit6weed/YNJE2GEX1JOaRWqizOFdW9T9tefKY3VwGBAzV4dN7GXiM+Fjwlc
KL1rkgKB5OuR9Qu9e0hKAxzGcKvnvRL2UAnYAZD2GC6Wid1hzo+jw/RhkRyJ
GGtfOoDpp7rzoYiSXf+8MrxO0bVhZec1B0SbPrpXw4MTrUp14C8rKAuirVON
afnoMNetchRHkKrfFXodAfjigKTnxDTuorZ+onLlGPKjgiOq8hjkJ/oe+0Tb
wM0cYWixDCTfYrl3TTnvx4vADIvkoxR89cP6AWh1hm41DojYXISsw/qzumvr
GqRnl6SQnINVFEUw6FFZ7CKPKKNVnZ9+bA2SIZKVgdn3oN0k9C4zzBNCTugL
m3cTjDX9EKzW2woRZphpJuddN4aOdHvQEro9Hn5O5qO1osW73cKVUPII4mmn
oC98aQm0D1TtMDwWGDoXbZWz3YBirNx7t8fBoVCHCGHAQIM7CqAaLnvo8nEy
0HU4UPCPyVtNCqVhAiviBVCXqJl0EUReH89IPo1rNrdZ7xr5Rjfe3GD4qkey
DE2Np0fqIWP/jKw1031drk5RBYkeE1ziESp/YFpB3C6LCWVAqYebbsSZlgfb
/Rt3JFUBDlMtxPGjX20Mq9CNAJWJK4EELPuvKv2Cg0oZ2Q3QmfSd0/2eUQl8
o14JFNYp81416TnXnCzsjwDaBQ95lWUNfh9XOaUYiEddRasFTIFINf+pc0P3
EwiPbcUiOtZ/Dc0gjd4vDT+kw9OEN0EadxI7mQG8j/mJjpsNYbFYVMIPNv/Q
Yj8n44RzdQXegeSz++rHaWw9X3cFNWpx35VYh7rgWKj9qM89JN1Ha9La1mqh
SvKNVW6irkknPNakEfg0wW6Z6arlFeuXmzC8XdlMme/IVzgXiWJN5pCo4vD8
wCOlFNmeL++ofIuJxj8+KSyoGDrNReU9BnmXHBOIj2BCfgBdE09evnpjWqkL
9aZmGaXp9yFGYgHamyWN1IsDAW9raLXq7nJQHFPZloVjKESsMQ1CFxk0evta
0DgP3szwBSQSfF7E20RD1jaadYn+0DzV0kWsmE0vMbN7OBZtYa68URKP0CgJ
e2K3z3XmKuFv9E1DOSYA9BUAuHC8cdIVCpyoYfF51quqH/UsLXTtEcM3/gTf
nXKkImFalL8/vBKYgTDCinMM/O9mvL7pUpmsFHlMcESugCl7qWffCykWKe0u
Acj1n7xRnS/kfHZMGDj7H72GMyjOtoFHQNTU9IXDvPGqjMN6CqEV9S9ojZr3
RucAM+StCsufTUY35ConX0g61WT9KPFcexWAPGqkkvnYZMaC0NwdW9yDgkkl
/ZBuuQvorKENWIAPrX/LLuwfbzrqrXMxnDP6wb/pnhpU0QXmMya8ZXBMEkoV
MoQu7yMvtEziJQdsaixfpb28GBfuj5OlDnurkq2FaKT/bFewAxwV+hWdYf5q
X5ikIekp3kseqAEOJahIi7TON0QR0794AkhL2LbZL6gWkwC0Qft7fc7QlW0d
GI2jki0MLMjs0g5DpJdsbyqWgdgtKWcrr/oegzSsavR4TRr40hVwQSgjccPQ
3s9koQ1NRgdLLH0XYFER89DVxFEPjhdo1TvBohcW2K7S4PF4YTeQLVPnKCyh
GfIefgXdYOnhCiyKaoN6W3zmx1N/TeVH6Ilx+TVsS/TxaiawB2vtLp96RWze
LmDK+M+dhzukcRb7B0HUMT9T6FPIbKwengwokY9V2a+G/1MKL/9skPfjsVA0
YButtk+DsXiuE2e8VdgHwmFQtZ2dYIorWZtmMOYEBOVk5avuamgBB/iLPC35
Ox/q44+20Vb41Q9hmmEKzNREdg+sB9zTkTxWqCyjvA2zQIpJkVAcckqxNg3b
nJLuPQlKQgxq6BnQLLf8fFFvsRCo9QNajmLbHKXBwXURBFz42OOzdSyh3WYV
UVzoYozjs7YT1ONY60d1Tep565OLMe/z4H01B7YkMwlGXlHslABYdklvGHdp
tuXVAnyTSjfFiAaQae8/mSb75dwG/pTblvtUZPxkLnp36WgMFIrjnLKtMNZS
33JG/wNFrqACuf134OayEb838fFrGJ40T2tyJx3Am2Z1pcl726PYUywgRUob
N32GJJTkC7sC6LeRr2zRMUlZVMXUaNdXT+hq4i5RrxSkXwvErrL4sbN2kQcV
IoQ6hOTg0aqNabTv8VBRAslsEjD/qktSNrrYyg6CmX9+Gr1sZ387YlXrQ/zg
Cxui+y5kbYNnG6MqCFYddFOJYEXArrGnXW6bRw2CaiFI1/BBu+qf/CVt2yqs
Y5bm38SXxIlNiaMC3tt6k7VOlVKwQzWa/whN3PvpldwnAZOohRH09TBLCovq
UMLg3gBk0jOZsWXn3AlzP9KieZrqkAs5Hbdk+yMQSc6Kzq8cos1haXR5KCQB
gSEd7MPEAiDDjewrb1+YfmqUyfsXgTZQdTsWQdpcC9zDWndyYleQ4pAG3J6c
uLmrp/lCkzXUuWa7SWYtvzmfzdbhlq4EWq3hDRTCYe/Whn37FKjsTrqzgFGf
dTH/ZUnN80pHiay3hGy5QcuJBD9eaJ17ySiKEmY0d70NdFgdLOYZTDc9IFvL
Ps/jvwFwteQTt6eoeZfvp4vnGpT4SF7pAsGs2LMqPSDBtwDQXHt/RFYoXj8J
CEI9Pq5orAbSw8nmT4lMSOpb+pLwzT6PmxWkmec94z0Q3RNg0rbQQG7yuI0Y
XS2DP7UpYJ0QF8uWJ1D6QfNwOMtM7hHFo94vTqJpQLiSJqW8tG3I0m7K+ers
e3Z7SfwHeuNz/LshP1As5veiKYufkXuXKdCYZr5A1wIBEzzR6AG2ByMeO9PU
GY1YIzqPTICa/mB9S6lFj6FSjfxLAnkeHaeHHUMrn5HiwzssLln+O3lTmnuT
xFQROiXKDn97LeXr+OhXeOUyViBOEqqf/HsFZtSdnlvc7xrLe/KuAsEosAM9
hTIFRz5DVJA8eqkBrt3KRaGA7e5Q9k+Qht5V1vJK2Qhvs3QcZziOHo5+9+u1
zXZTsF4GHfBjROL0ATvpW0dSKGRHXOe7DHyndomwzefiBuD0w891p7j2Yv9w
+XaY4+1I+pUUks7lBHt+c9MRc4im/5DMvjLaVLdjA8XP+rDOais7FhfzVpeU
k/4Wc6atZ4xNkRgflL4t2Bkv7sPJhXUF08HK7Z9po66z1jzhoKuJNHCnwWOx
70CDfLKj/KZx6dW+J+7j9N2rASNtX3KnBY9pWMUNj0ar4s9HY0kZVqV6Bz8L
u8H4m5thBv3njdSwflpyoLAyaU/N/bzW2q86hSeHhi79Ut1pKWLzFOk9srTD
srf9/IP+Ds3Yh4f4+y+fVsPzFNrhSa0PVRZeWVVmEJqL2mHfQP1MoVV0GB2G
hAfwHkOw6gBvBoQzC+yro0NQ62jRbiZ4xH4GVXwWrMdxw/RmR0/23IsR+qU+
bn5Q6cM1nkRYTFm8wCcRY8VIKmZCc+Qb73YIhAEe546M9cYO6bqva9P1OsP6
2P0NQSx3jD04N7vG9Q9jDD+6BMIuR1bUXQwkbiP6x4YyV+prHKhpJBdxVQa1
CLsnwR1V1gVSzkPZN0mh2b3/oIq12sE4cMk9o5Z36buoIsJZQ9ZkDIfdu+Bx
qUS7Xd6aPfQa7M+K8oEk/V7JaPGNi+bjwhLDYHZAaoPKNmAggo8w8rnG7Z5O
yDVG+1fM3W7ByIt74P5NCmy1gYD5oI0mGOB/uNxncoXeofIFSWZphwCr/CMV
QQP3/s5p+/duzvGsKplX1Q3VZY3Xtj3zMk0NuFQ0pmGZaYJD4EhsTMpmnQ1v
/jE4P0AMkxj6vhecvDUrd+DemHf1VPnIdgiMyZdLWXnofUME8HJHI3NTjoKJ
hFw9ujPcL34T61WAVaZIGPv/jgqcbnWimG2PFE4nvXB5SxdxY1hW4eYWII5/
mSjfUOeSsY1YHz+V5zG060zkPV4QWbtAEyS9oR+1jotb/ONfaRhqcXZyFil0
Tab7mYnhMVsQbTWzjaeYShA8GDqbXV+nmvJ3FcwtYdEGEgQ+3Q+jpQvPx6ot
vEsV9t19AqkU6hnqLf96a8iL9rS/euRf0kFgZDnW7lqoTfpiKRpEJeMytsqZ
xqaF3TjqZHynLtL69Jf48awZXETBV1HXHLYpAobxGJrlLeCasrIHDCb6jc0S
ygzHKptbz8dS9rwamgITRsBemHSDVCF/yF4QM0diDcc1k4N2cm6Z88gFQofL
a6LT0ATrhz3uVzZWE0+n6WK6qWvrLGsjY/yr6ZuC40HAyEGTqF9I9NbKx3fS
uVfCcqPZV1KHQN0jhbABPVq8RyAq2r1zpd9WrtciYzJmFINb4QD4ZbTDG35I
zG0Ru2Ezyy3m7T9e2rCiY7c4+0BrIIkgkJeEuna+i2zkH0T/0wInf+KfNpSn
2EGVU8GGq5J+wlTHDJ03e69ias5KjY6JodR19mROWaGBPE69eUfIQ3SxnaKU
oEMzXlBgQ7EcBWecfTSU7wT3znrFvt6fFxbQAR8fhty9wTFBIS/0ImEv6TCh
8HrqNaJFOKhesjmzrXgLqr8mTic5gwLE0hliPU/dpxiWNgfGDPL6XsdTB0FJ
sgSY6fB84WXk94tcRw1l8W/JobRY5UpPHl7HLd5OySHPo2O7PO9LwUZ8H9pl
m1qeLdgGoFyC72YnHcS26wdUFR3nPbC98XOVe0E4TX9cOGxwZLtP2Z6rHjoK
03YLlUFopQ2OXtB0g0mnfw9yO5x45ratCCkNqwqeNU9HI1aTCf6x0VlD30mp
ptQIWzOoL6ewksigj/JP0T7ZSVXKmRV+URxGzyzuYVmwyU3/O6Rh25ifgEnc
+x5hZkAuZTGAR7fuuXV5dtyhIw5L6L3bnmENqYfUNXZxvxuaXsw19Kstw+Nx
qIEaD+3bSWokDpO1kAZEeG4SgnL9tf3JJdz2RzxqZJc7BvLA3clEMjyV9Z8U
bGihzzMCXv8J//SdKIXDWOgaCDXwK9LztDULjivw+JrP10dwojbObnWdcYaz
metoDeiTpuuvKobtk2aKKSWKN+n1jIKAQarjWox+0vP9p3yoOwSbtLw8vThh
WpSPNrHmCE1/BLMSKtAIzUL6mN5wYbGVzjdDdMJ4VTZRk2YQ0gs5hVKQfi0e
4bGYX8bn3okvwFRFEc1Frp2f83ACQLp2HOXMa1gLeWFuokwZmJjPK/0k2M0v
FUdjZFngNGYsA9r1a9m65WaHpgxVCe1j2ZMCGdBBQOcB9rVOdGs0Ow/dC/RJ
ZzR5/t/NAQlOgxCadXk9iak9akzhZWvDb9ZX4Yx1+C8EM90zS12arVznMoVF
OfoRpXGWXmQoOPEve/6alVR9QTUsZjYtXScj6ROhjs6Md3STvwI5RWr/fjeo
6vlaEqGTL8vmtx33JncQqvfDlU0Swpnx1lStbL7tsKqc//Owalhc3yVmpmUl
D4xpJa6oRs9z9fkatgXxNqPbB9g3JnG6POw8qH0o3Md63IpiV5lPXo9P2opw
wZLekVOeod6DN7ZWSrhU5lq4/NCnp5IvffeF7oaFpsN+qAA08O6TNll6wyjo
Uoey56JQ4jejzkhxP2jw4ieem6quMl0Y8yPKm5cs3RhHoCx3dk7wEVrZEXkA
xLwoY5Evwth7Iz5soL8lWIQBTF10NMIxuxeL7TVraBaxJNojP9XiNB9l3a2V
UQGbMzEJkDrvkcTeF7b22vrsowCHzIHEYHRJ09tc8+o4iuzbBDcQjvfwCuaG
rBdbj7fKmwGrYOvxBrsC/PUqtJ5U9x0PMpEOAKaK9uGdpdZbHT0Y9Vjxc2Ed
QQisg/ABpOxzJqWxdtV2i6WZ6tuZ2gOZuWl1q/n8AJdhe+u1uVWbtFRDxuWP
dkSpziNG+IEcxuXj2cA7sOFmfu6WBi9/CucyWwYS6tecLXGBKvZbfiqjo9kS
y3yDTsc3WmfnL3PxgIlBJJzlxk71fLRLPmD9BP6aPBinty+TolSAzs1yzAxk
K1TOBFvpvUnUCRfDm6eOz9WzN46HJxDkWWPuqgavhioFsJJNyIE2RJhsJNHy
tgtuRlqgyHTs+QZIo01wPkuJc6pk8FkBEqh5mwXy0RwwKrdRPfjG1Si2tV0X
NNL5RjEOcmRyWSuBCkopERuDXdlKIIK1w00kBmWXolR4Coj12gYSr9GQNP5l
riB9qiN3vB9jQXNNppRB36IZrgA4LEBiDCpPZYUaAMhyt4OSC0wi0tu/rsdB
TGk10jt52y72kj27rSYeylT09i/3c5LAJ29Sh83Pcz+hV8dfLmV/ewcELS9X
BEW5JM51T01DntaO5SHEYV2EJ80SF31kZCkFFNZ3NoGvJfdMkOaPEuMJ6DXv
ocpkkoTjLr6KcpeUW+PKG0AX7fpzK4ijhVrZuiqTSgrL+M1hVLh4HdpIHpwL
bsmN6ZznvR9s5FK6YzLPJ5SmJu/hj8mL6GDJyD9OwU+3us1NLJqYDxsDOtB2
05RSSVfz8XXpCZmrfYD9ubQdkmnSVV+dC01lzxhVA89f1XiqrCWxxkGuMdhM
xfYrTegitAPJMyp0im5+kZK1Q45uNC32f9NKrKdlxNPh3cvbL2Y7dQ+ftVfJ
0AvR9K89EFEhm4Oocp2iYKDz4vVOorU5ZQ8fwT3ObmTooB8cX879IH6kYroe
3/eae58rrGUjvamjuCZfTflkt40msPtOXaeT2FMHyEsRrJWBUU91VdegceR3
KExMxXaFiAMcbUsyI1qv7TvKBoLn8tvuAPI3pK4jSAp0i0hTaRgaWDf35wkw
6WFxYmpJTIUw3nSb5bLvgGA17HPkdSr1m9AlZ3EDRMi/cpdo/AYiy/JwRCIa
CWHFrI63Yx5HwS5RT2E3XyWNetnAEJRmcmsekBf5j8HSmWNCJ6g4t79Po9vE
SkatVgxZg2Qnm6TJwt/bqikEhmBZhyqIqN0hZWBOJxsfZq6C6CuBbdhlqz9r
NOIkbJR8XsH6BisD9ONirktLJely4YZlywVaezGbkhIx/xp72gkWrilNRz2G
6YwB8T/Wz/6ffz96s6D5aH0Let86HkLP1Efe1kuaWwerDXQpv78gUv+LB1wr
wNoMB03RZ+c16AaZPIv+ODFKMQgWjsbWZEaPTRhnNT/JFpXxMziE8LrtKAIV
rjQ7o8AtNWuGsJddJTiUpu/Jg+N5FJpzgAQx8aM5XqXbNAGfxOCrzDRFbFA7
OHG4g3j4/Au3cDHay2VFeGu/txn7ahLbL8km7snONoI3M/7dOfBYuRtPb/oH
WpQl+l/PPlBdBjJgCITT88fZripSHarV9P2KfRxLLtiGRc5fjoMRoZfPlwUj
nsen0d9A9fa5zRuOG0KxcMbiCC/b9xI56h7ftKLJ1TKO4ff61gcF+24R1jFM
Cadoeq772/Xsxz1Bi0+E9Krvnfaw0EEoHRrkHrUqqTPDaWr4M4ooo1XiWz4A
0S3tObn2XNjL5XawN/OADLjstRDb7ffaqH9LRHw+nZlFOrFHrAo+I2wq8yEM
sxHO3Cc4NyCgnyV2xKoz07wVNq2m1cRU+hjObkAFhV8GEAee6xNewV+OGNHX
s58v9vZ07QfPpDrtc6LD30wQ6UTw8NtMnubqruwcG3HgtLGT8QR0GINxZkv+
CupXhYFJABpT7EKjdpo2SyF0TtDuQ47TPDj9ierGWPa+1yyus5sNb9xJO0PL
/9D0IRMX9nPEmKaT5twPFgWPnBsQ+bNvbGXdIqTr02zk6bITiI5zsAw8Wnh1
77Kvuzk0pCCKienQKADlL4svEeFOvQ44IyHg8aCfuoN7F9oMHMm5fHpCMs3t
D9bl09/pgH6MMR0Gka+o1FLDHbdtjTCT6E0g0g4SOVfngN32lKZDVXS8h/21
lSBVyBB13Jyfbg2oaGlqsATUkVTYf4xY3WuiVOHb5qrlWRWsVeq5HlmFPlrf
rAt88MSF7kjGi2pa4WGns0SOt+iFNz6CRqS2H+B7FEvqHKX9xypKlPfJ6OMK
61qVrTsiFMf7/GKuRGrFYGSL6wmHHbongp4xtEOo8r5rhJFKNfmDT5m7agk8
557XVeiqiq1exQCKYowAPKxYOwfNPamQ5njUWOMLlHEplkK+812p6jPsK38L
SJw67cs5ZVJA7/1IcgaMMMz6eEnKNU4BXp+1IFq+LjRoNyGLaKGA1u6k9lD8
w31/2+eCV/mgjl6M94a+MCcpZikLAf6+k/GD9x+GBpkB06tLasZca8+bfD8s
LiWUoqp6ZZaBL8qXlyGCgo8WzPiyRr+bxsBkv5U75zHcgPkHVA9m9fBwsdYi
uAZLOfm1P1x3BHMjoOkXwRAcWPVeYtO9K09d9DzZCbC/J+KDbOuuKxM1/oEr
hKxXGe+cPXDsvtl9kZkf6edmh9IGSSKiCJt7cNDchgD1ob4dxyrok2vfNY2w
OsekOrPridIASgjsoBKwP1dZudL768hYe3txZU4GgtQ00AKN1MMAzcAwYxei
BzJ56sqnk6y20Oeyzfa41Hek/hkKD91xdgPHCb6M4l85ky3OmxNaJaW5mdip
oFovlMNqmH14p3fvhmN+XNf3VrPXAv+S3g8u3n3mUB9tpxIZEehzGVifp29a
vpNaYTvQKOC2yyGtoi26FT8zEu4gtZuclYU3UiKlX0IHMFcI9v53JJ2pmoCc
eKTjX45W80v9S8HMRLJOHOnVxd9DbN9u6j3Do52zm/Gpss8RbAgx9+hsyE6q
OGZ3QaH484elpNGsPiUvQawJA2fZ4PYARYMvz9/mms4qzgSStAVpLfGI/1jq
yWn14CXMg+dGMAeQl3he+xi1AkT/4blo3u2vD8DxDyRCRgoXVYnvygyUu25V
7VkhO9411Vpe8QceYIzUPn6F2HiRyUYLpVJ6oDz/XnLBN1HDUfaGkTWJujuG
ffatoSh6r/RpDve5wQJEGYHrq64yAlznD19+GRX07ozIK6adxh5Oh/gq8igF
ExOQQW0VFPtHoUqfRs4DlT3588x5JdIMcQqTzPgEawuOE4BX8DpLJkiNGM1B
7MyeLk3N57OyvAsVyXI2TV43Z1+o51kEdT+MJ68mLX06i4PF0XHRNLtuX7wu
r/pxRVBwUTjkQ91Slk84mOSgnXM65zs7V1xaPWgHdZvSXqciab0fdZqM3twG
rC8ozad7wdkJg7mrYkUfvApsiQi0/iWk1iPx3gAPR2QqOgZgLhIio+e8Key5
9XMhZXJ235lq6JPgRySHQC1o01qgM9iuwT6sacO4y5lcLgmCjsv8CUn6Q2Zn
csXKybJvKxcAgsFExVSJBOqsJgkzmkPoOlsKzvxJnE4oKLM/6cHpFZ+R6dwW
bUOx7oDcD2d471GzTCvh2jDvBBBsfX01Z4RjNxB9azfdlbRgNcdST1yUTblr
bbfzmvtyKUFjzoxTzUzcO2hgHPmRbMr6uhshMyETkMVBeiORn758ZRmJkhEQ
Y6GF2xJIbH6lwB+U3PTjcFw1/wJu7NX2Hr2J3MS5hhnHHgdCq02saXG2J18m
bix4ttTuThgawkBlwnIr1FDuG2epfIxltPW4fUbVQL8ObWfRTIeu8loY5o9b
VvIhEOpcfTLKoAV+99X91d6/6oeQlOBpCDOTzh3kfiCv0ibJf89AHp6KkXA1
7H15Q+3ajIodYush6MBIiG0m6B/Tn2mNrWvzApM/JPls5G4W9StV4MvjksrJ
ZVmw3VAT9MhWiKy5lyeiuxh01i9loZinQ9YNiIdjjSvrq4szBJd7gDpjwCmn
RPr+HoTEzqM/ETp21Si9txw0RczNb0ECYI2LgSDhCbL63TyDxAVgvNuouLnp
GiXGuD/m7Heu5l10wOdpp4ETNPxvKerkZ5GwbH0wmw4hZMBU2bAa9wCpy/NO
qBMA2LFOcthsbNSDWzxcP5EyHZ3PlhXeZCvY6QZVl9lkChngJfgE7QkOe45O
XalpbIc1oQX/IG9vZi4d9jIOGNktjrjXeeVnBM6TN1TS2Yl6pZAH0e/D5KRQ
vJO4I498DDH504VtJLTTQO5xPXmJlZMB2EV+MGu9+ZENGYaIopCWX8JUUZU8
HQ7XAqcjR/jEtO+mfLE0GrrmHpjzwFnAPWcfEiAXM6ftZiV3MfEAxdBPwMMK
n3JkiIEPfU/w8TcwYhK4eqoUow/RwcDnadYDVAaGsQafh1FjEfAtfeROS7GI
GaY2yiRfbh9r2NX07xx0bcx3gIHSxv6MbLb0vNs7CLlKO6guA1FD3uvYRf7c
OTjxN8sRSo7pWgCrjSdYmh7UFxpuaeg8h2o1cMDGG2xA1x5/nZgIBj2kI5NE
VQI8Y8ieqB+NrR8INl2wd7n4zmK8+YE3RGikVKbardTF88a1TabtX8nDiK7F
sT6QfLdBQx5N5Jn6LZUzMETqHSk9lW/KFb3DtYeTJTf/6Qve/s7wR3kHioCa
wj+9jSMftytLWxZr/2fpW633+z5qzYCpQb1yqzJ+0+gERYygENgbbOgfwtbY
OQsFmCRtM9j9Xuzs8DYmf0/mduM2PYaRotqY65k1JAXiF2dlC5vj+Du6B18+
0tOA17fZhZHVo4faopjz3M0CsHXUXfAL0UpaS9OQpP5hZ9uDk2EYi7rfIJCU
2Bek1JxEXehC6P/JzqBMXIxAAJxSHrBfLslB5ASS5d85StS/q4sqLi11mqen
tqJfgIZt1zTh7LtC5cl++4kxaBslBJVJDsKgFljWTKM1aqKV/c9QC5Zoyzs4
1syM72DMsawv9iFVVXh1671JtOXb9G+ZO3YpUJMnhwiT0fgIq+n1MSpSP6HI
WOCrRE/761MdcLIYAXVsdkrSwXnLVfGgUv0P53EXGeTEHBULVClGcUrxC/q6
5cu42yBu2xkvvCPbbJUtk/yEFdFd4zCgdoKT5DJAzZ7XDWY1lJJD5kGB6uuv
+5XvHdox2tr9j5pwWlhbZzCTjvS6n7MqE1/y9fhtBBUV7Ko1IxM1qKpc0aVA
zBPa4Z8lgqsBHLyX7mYSjnHtMTPCjy8NsInRf6SHBhZyuM65ID8k7N/sD/o0
BzpqTtjs/iXtv7FcurSx8YzxwZrMz8wFoFQDOfG88Ns5tPr2Cfy8geHFe/k4
VwPZke+sQigbHF6ndl4oKYxCCCmeIdzv/lAJNytlajBza4TOEqgQJm1JVECq
3lJBqhqt+93dZX5ObS3v6WAl+BDcVHllvSX0xtyir3pY956LqHYosJKjIZNo
fcfDd7EcT3oaohyZRAWTo+Yj/8/8aLOX4GV4cwf2HG1XrAvWYq/WRxz6SRl2
y0iD9FTz6TRDW9xJQ0AaiurP1yRgiMMPhWTJ0FnOXa8RC4WjM7jJV+FFBJ79
fOIT2+QEgyeMhkvprskg3MfLcdz1hb0ttg7Uo0rDli964/mDAsz8a8LmQU21
rQT8honTg9ys5tSTbACTHHZ9EAWWNESgGGEg9MMf1siD6K57FquUJcRv9oJe
b0IWqB+5mytHJw/PWj0Z6S7noZsE3BeBOPXbzkxrTG/wFiZkpc9cxHgxcOZ0
pDKwRn0F4fgqpuykVUHhwQq9kbXWxhHwQ5DnUI693O4nzPFcw9GQWmJVM5u5
VZMepWjzsX+LX0BT/deqIxbJwg1KXDJVYVIn8i0eaUeex8jlOszdTJ9+ZfgI
bf0T52PdQwTg74VDKd+ZuWWnM1sXY2mxfYVkadpJwnMNvXexMu1Wy4GEwtoK
1dy5YqQonHke6XEPrHhaJbkYU1dLE9KtHoLv9AcSKaRZAXXOcCqr5bRlZ+7o
9p0VVazmx/h7EjKjbfA4zhgKMF/TYsEdh9DD+kFqQutQfNVH8SbpgvTjH/jc
IqJftCvJEr8tW4Y6tHkWbVYMwy1W8how/FMLHWN356lsB8OXfSS/Tv5CerjC
WU3z34VYxlaFmZxEdp0VddJzLwIDn7CL0kezegDTfgqrxGXrQEi3DKZz9NAk
Nu4EB8AAWl1bQw9rSnhk+0TzvuKoXg0hVro18KTOFkn02WvF1e5s+4e41+5Z
Rd3vwcPtleHkjEC3Z2XHzZqcA2pkCxvoba96ssTsD4P6UpnW9BlUQRxGoTxA
pBH3REtRLfCVTE8OPM6d1WOregJbkMJSX3/hhjh2NENe/0wl6nzStLAlVpB/
fu4VAQkxgHXrMIGhZSjlyO6AVN62pRbwU+9YKIZDlJfuOf0hqno7WE4KHUCk
718lIfQ9ExAjORUDCV5WrSD/BRa+41HBzxXuWAs6qU838YKn4Jan3iSBXeK3
ukzwT9o9uHJ4udBuKk2A06Xtb2b7TNot7e+Mmd0/MVxi5dnuDlyW0MocDScl
CMkQ9+pDgDNysG3OyLInrqLDvPCurvvSSKmdB4pe06amAKKjDusa2eLMKZSF
Qzy9Pi3mzIoRLvNI+/MMHd1xMuyyFszsQUvZLx9Tmh+NrHEyBEBOxCEiTooH
2vhkCO7r1oVJMaN9FBLnbxwB5QULw7WBydr2/feem6ltOTXAbenRMvDthZZK
U44xFPmyeswW6cHcstA7/jSyah9fvKeaVU2z8vF8XnQMXIiGcRxH58GnzE+y
/CqWLJbUgNUQ7TzlMBoxp9Bc7S6nE8mwxocgBzYjKq8D4SmDJriUSmjssACb
ARE3i2A4jz5t3XYvfbC8geTq7JkrAYZPksNwSRjuoxwhD7FXC3YSTioSTLKO
qyY+WUCSY+ijoJ5pwX+UJPhQwujRLQIrxIyFoGjAIGCdmCik173ddJmDsuTI
rOQ7YDUNB1uJ9dmrdW07iIXnjWz+zUIFaDFnbfuGurEIIVguvQmaHCpGgyy6
JjZhxu3ufU+zS7zOqFKtMCZRyouZmEf09dL5sxvOJrPA/P+2Db2EoBkbD/f3
OKlAwzCD0N27STO/WCDNo0SNp2p4gyotaIBLk/wEhxt9uVAPnfiheiMN6Qjr
tYqMCXd/qhH0CqQ6YO5A8CGevIrlUcufAvhwNwncRvfODOhC2FVLMrQuJenV
8IenG6YCwdptSEqIyRVzd0PCfi+I3iuuP8R/DQe+o0D0OPUwkw3rawkEcv0/
TwgUYvoL0zKW9aP+ioz/fvFULgck3q2QX+6Q7yzrgIIunuxy/q5krBXulHTn
w9cd4mqwq9A1t1ngp3pKrTs4vd8wsxVNKEYvY4AU+6Su1EVe9jKT1hwoWT6H
cXMnJ2/sGFQ3IpvZoVIkpO8UIL7ChpzNGI9B7bWTT06xkJ/QQ52+aFxokVO3
JfySoExZ5rR33tgD6sJRY2Es5zZXG5cptTMh41HTRYD1uDx8IBIl2nl/tIlp
Q/YaoI5f1Ab+WQVqaRC7YAZE4MrEtjud7jP4bJE2RzNR3cOJd8faOuigYBNg
ZJyEkoUwdURu2fn2sO+iNNV0p7ZmuvKPG6+RaG9SlM/P/PJKyakvJ0ThLMRp
Ys98AoBHK1bSRzgTDRw+XQBThTHl+TLl4pHVkSfe0vMEha/jIB1rblS+PPXB
rLjbl85azrZbY90ci2khlOjgJHT47Tywtffn9BHyQCdEQFPJiUHxh5fTzk3i
5vPbeoiX6HvNtkC2GvUdAulFHr3j6qpNDV8fXgSJvv8+ft/+A7uaSiXmR8KG
aWcJnEo+pHF1T4i0UaKtX8hhvPa3C+MUH8LUmgKxsRWo76lOzNR7ZqXQu1wg
/nkZOZ4AZzY8BCNitK+fihLPskYTtri+GK1XdKh7W2J85/1D9YTwB7F/s051
3CcCURBZ9NYM0K9dqSh/mpd52QE9lBj77Er4Iix/tjETWYO8YChk5fbhtEL7
DSn2llvl3ykcZPuvXSU/127q+lKNsr5f62m9CSmpb9zlzyHDAI7Ao90rYT9T
HG8ZnAZBJ4krCpVhdowvOE9d2lYvqTWa+l0zAEAGvACxp1J65a/ogrV1rTSY
2aVeKiaIgnpB6y9ab3grdSBXPdwEUdIt98c/xTObA7p1o9SJ0h9arrLEHubF
geGh+a7+1zvWRCnvVqtBafHo7Lf9LqM72I9mG1Ce+ynapaIQkmSySTHjXwvk
bT4Nly1IWZrriAwxu6fPYY16ENnDYxIdw4slRAp/GsEGlNI9aOqJ6KZ1SfwJ
pjA8psZZ7XFseHkVdUCapE4/ROyzlm4LOY6J5+ux4+Ui128qeUUGfyxfnUbF
abgq6VDqpuuzaWBdrnyjcmaHQDuKCkiJ7F5lrbGMJSPwi/dTVeKQzGlpTcna
2B8jtFsoR7dybNfbBW0mL/trz1gBnaZo4KzcUkOoHvIaCeBmm0Os1RTHvLVk
DQsPpRG68NDVl2fl5uzHykNy9rKgPlE0NB2ePLqPvB8eCNqLqEfRj21xqMsA
4Jf4O2L1k/UB0+aZKfcRFWEAQZ2ZKEK4rxglfr1MmVBNBshJldpV5uZcepDy
+T4jcFDcd++eUCkKPjis9qNUqTPBBlOhQnNlXxzhgWx/QNm70A7uXC6IDld/
hifNeiDvAyH6H6NEfyrKBj5o30T8Zwpum6W61LXBmG0l+1hJHixR4074QoFq
gYWJA8dLxnOMJ108QaHkEKVMFkpC9wqSwO1clkS3ZwB1+t4s74K9pZoi3Azq
dIotWH0SZ1fuHC5kPjs0U8FltbnT91a7xLs9uqZIRLFF/yjFFEo13jJSDSue
O4KrgXaVqzXj52Ignrnlq2cism3TGVsyvFRONn11vI3w65N9bW7D89In5V1N
a+Dd9dEsehEaVw9xMLC42Ia7Lk7rbCyq3o3VXo/Cv6C+p8yHTkPlCJYypAT6
bBIdNQmxvWKxzi3Eu+vzVVjQRheL2hIAOE9c9hzshK/4a1Y2L8EvS3vutJDp
O5hOBGaA+d31e71VsLQKbD5KJc0lWvVrnI/oeagkbm8lc/FjINRXyPVvPoLz
qbUE6zZ04Y3qTTriTFfIigmMoSHiIgfruaY28b+maDrl1o+ng4MTaCyrtlDU
jZjM3VTdZ/tTz/mjbxQFaE0x0pT3Hh+ShVNDFahYr1oOerRdRmJxZAi8MjCZ
tTiuopwrsO+nXynxvf5Y15f2fkMq7n01tHjAWV1J/Q9XW1t9grZZjHZVKeko
kjXEeZOVqyjX1sss56qIS1mfwhgBaZPhKlmQHZIFfhZUAK7qb50YAF/Sq5jf
hkX8euN6ulFsWO72RLzCREuVsx2W0AsN3siqqQA5KlIxdMfwP7CtzV6wARvy
L6T1VDsz8OgD+drbbKfipQF2rMy70keZVpNkCj88Fa9xX/jiwrAAAljqxYnX
zUUoZRUJIt4972JDp4pIlmDVP7PH+7U8nXyG1J7cw3+op/fUdXED1WtRfQA8
IV9VaCshmaHhT9qZctaIZ1H55rDep723wOXINumHeN6H1zGBOCPOmx68RmiM
aGIJCfgWAD/HnAN1QVxbvmONZmTHdx9VrVXys90CYyPJXvNTxu8W8LsNAY/q
2zw+jvueZA01VbqxKX2sRUqemjb1S1aBVvBRAC7vxmsmNUDAR6eFDcFEFBPK
T37mS7dn9WQRsr4LqKxkBGv/SlhkdC3V7ZBnb/7AbwfUpKQ6IbfHKngYAEk0
yKRJ/2MpP/9sBPls+0cAQjufGiLPeSzWWP8zAMb5AQ6mzUzp2x03uB7IkQsX
E5ivpzmtp2pvlLOkMdUW0AX5hDH7cOYbz21i8Hxn1EA50/uBTDvwEAuRVEoF
vfoXuRKLLJ4NfD/NzGIpPpeEVVY6K0X+Bu4WyvAkvcfJsaD/JZMAJUqYSv0C
DtO9FHR2Hqziqikt0EWkWGfALuZg0LiCJuJZfeG4n5m0UXA0SNeLuqGFK4sE
iZR7vi9R4Zx7NljEo0aseXp3xvXggRvpYVGw2zqyE3A/YK214wwYwycURE8I
Iit+1ZmLrJzxoI7TNClRBHId7DH7BRxgKC+AxVPmJinlXgTBC1EDRJjNNxMV
/DQr9km1N14o+rSId2487IlmPb4kaTtClp45PV0q8qE/NnKfdhICgBYKVY8B
xQ4Cn2ALC/XNY65Hmzw8/wWGyv7WO2z+t/WXVkQna4qNqTT9A0nVuh6XaJdU
O/poVIYUxe13wiFJrdb/mjFbmQnegdwuS7I9qaxzPpwXiELM9n6ZqF+57Vji
jV7O2K1B7aGxsbqOGpOIJAFPvp41eoE9mSwNuEHAMXorV6sfne1NsyAcuwZn
LnmZTuwVd4WEwl6pdwDP16ytLSvlRyZ5TJaLrz21XD6v86kL/HEsoPqblW+h
9ldWsEiI3/yrbufE24PXUb0G6xr3T3SsHA3+YvpIOTzaY6+c6l/2xJhSnpF6
O022fAL55woFQNO4s6a8Tjr2vg01Japawh3CETKuzhCXpPlRG2Y3zXXfe4Xg
/ECr57r+ZVhhSNgWWnjtyq6oFJarxQgHAr5FrbJzJz60T4BLAWlY9Si88fnl
pUvOE4WbGBCtik/VC5g5mSqThOno1HP31oiqEXcBtflH6efPAE96MS1cYiCg
TubYUBL8Hnm8p9vhxJjiW5ojrWiMRENTQ+f1vYVnsjE2c90DfxJSY6iGTXxS
EPwew9Q5K9MVGnyV8ZiuNn9AQyTUkFxaCg34Z6xsjfHuSJUuN/ojKHEBalof
bWJOK7RHXuKDpyHhNz5qYYi8PvMlQPWja4TUH8Fz71+PCzDZCxdMJMbzaERq
YxODas6XYpYKD8/hxE0AKGe/fgO19fDdBuLQmHqKhUoeHF8KllQsnY1Ezb2u
dU14FiS7wEh8xnSJ9NYVvOu20aodKOWeylrGwfyzuGaWClhJSvYRvoD0NLFe
+ZyEfQdUbRAykRp6oCbM0vnCArnzdQziok0k8KzpLaq/dcMCKip0e9w/vvTG
nBKjoRSDFczMJG8wUcGUc6zD5Af86h02tZL4rvNYmCq/u9BT+wXnHg34KMU7
R+PuLx+XMv+fi9DHKuKlQKV02QDHWr0LYo8nzzF3Ya49s5lJcUxWyW2frdxh
fgInXyW31nKTXMVED2f0VLg386lGKgDi1OhLnFO1fJgWFtJqF5jKBnYKRuhp
Q/K2j9p2cLRGn5CnbIptRhM6IpOzb6JIqbmnk+R+8IDz+gdIipyRsmFYLj2g
t/Lr0+TKty2K51m3cpJRHxkYrt4xBxPyOCz8SkI7OzjfcBfKD1I8j0qAadKK
h3XOcRBYxdguI1qnzjSNjQadPrK290x/bY66vcLYaxs0xPe7C5y2IV5F5iVF
L3x3/itgpH0yMsNmsw9M5iHpimGwp4ZlDGMTnBYZdd0t21v5l7UCLjoddxly
OgW+Bb3Pi9KbdohtOFW4TJoDlWmzwNHWmn5C3nUIqVU7ApHy/OIUkhkxeCe9
R2CVV0Ktt4qW3T7xhDWMRA0g6XIU/fyY4KbAL0shzrliSTco3L07z9xVkghd
a1nA7fwZ5mtj+RhAPgwdNeLrG0wJBzu01lKGYDB+TjgDqUZRCYh3WMqeQV/M
02HhkwtRTcGtn5q8UCf0905Cf4VYetvuGm3yozfrLnu96d+jNK3jB+gKQsnU
9XjEuBy/JGUJvU2TTX1dAs1S9lLcMLwUCKasCrDdgLaNxh3CkWc7BGS0wmZg
eor9+T4m8DJrbB5echYrm2PTLcbmGDIql3UMsbJviZXKBCIGGznya+KWu5c+
jYBGz07vml5yQcFLVT9Xk3lNNJj/VsQjI3zeNudjsl00NALO1Trxg+51atfQ
qF8T0qAdjoz2oV7BKO+igRBQgzi7w1vfaOya0dc2hDehfDC+sMRFJJULluda
n4LC/0s35449A/DFS8XEJSmZONmWpUsflnj/c6OfD7Q350+9TS6P8qA8PZJv
RkpYRFY6wy5WptfMmkiNA++Xb2RggZGxKWAlz6GSExMbzEpurdLWmTBBZ3HH
DdJl2h3I242OYcICl5wtrpddxc1DV3gUghQuBRUTK0bNRICHbpl44jVU4Oqc
zbW5W0XdeMPLyiufjIqi2VDwcLpRJBU/nalluQdFX8oBcOLMHjBSv9SHJgHa
GteVLK+Xy9HXCCikHnRLdoBcJjQ6NIBZgiXs9/c8sRdQetx64ks3ETKT5WAf
SaP//Yn7Y+1w6NH1OyqKHfht+IFBrzdIU7DzshQH4KSO7LjTKfANJopjVm6q
vBBqz4VROi2OZKmUPJOWyW0xNyR7ed6YK1i9lhhhb9Yo4mfVD5eN9z2dMGvO
jRie85bnj0Cls9rCDUmY0TnWrCTjvfHGubre5JSz1NPUsM7Iw+MfHGfIsxrU
RQTXbaocuHCgHAeu4hda/m85wA3fu0G839HfgTMOh7mQjN+ca3B5nQcvjTOC
MJ4EGtrBgF8LpFZoU0Cedvri5aHaJoOpKkjq8vNEbq6ey3jGtZcXnpdTG4W+
UOEqoSMdXbnk1+K4SZygloNJe8WV1uxOrgpaoq6wrCmNvACMVtWWjKvQgCJr
AL2fCW7z9sc0/+ZfpXk7g7o1zW77WRajmcRosmQ3rZY7lZyz0/F81/tUs8nA
165CKnw3x0jnxoeMTCLqFoXFKq+7qwWOyy8Coely7kkPdoguqS8zLldes0xF
61Hb8b3k5fNWTAqfNlitTyYUaMsMxgpX/xrX7+wE97lxq/+WJ26cUkS90E10
NXJ3cd2ENvbtACDN17mpdS1GXsstnxBqAmKtpDwDGHLVijZnrqnzXuBCp4uU
Y9UQav9pwE9iYGE8aznRg0K66bTrAjcv0G0v2dEuGAAbsl6d3MGNPS5/0iCG
2s6XopksKDYqex1NtS3cAlU7lxVRRAbHuCdp6t4BiBSCwiT2MAsXOu6IN/jK
L6kMKwpBqKeG1cSJZ+PZhHN9fK27iBWv+k8eUoaJvLXwkyeGhKK03r/SRZOt
sBQj1aoY6fK+ABGxx+OSm7geMrvAP+Tuyup0KhatSQQEcmlJxHFDmLz3hDgx
naqEAUcUfoKZ1u4z80fp6pPJ77dqS+kAocvbbY+FRXlhQmZqiyydxxc7SNlv
vY4Ezq2wUGGDRufNIVedu2MVLAS2UytWl8z26td6OMANZwsX/e+PFv4XHv+E
hVkObu8wG6ePrhmIS2f4Q7VS7WhI+5GHNx6GqPBukp0oCzASw6zYSNR9X980
X13pQ2qnJGA6qGQmNasyaGyFrdvWkJ47OdIkFHfhyvtY7FMgbMki1M5qA3WD
yopoy+7FBK9SXICcC/Tx0XssAyUDfL4NQDoVNE6+DkJfmQXfqbqpN9QuX6q0
AxECPilxY8z5CRY8kgZMgbXyh6uCBa6AQexuEWdCSGRoVQrr8QyWiszMC72O
IhiEpjHB85jbrNJaYBBL9p733rnCDDD52d0PIJvisR1QQopQ3KDnwwaychaN
UtQaYZNNF9+65YeSrFe9KcoFj3jzXnaoFfLCRNV5CGBcyOunZATIbvXT755Q
ZixqStWJIEef72xvFkla83zt9ym1NFaPvFYTfY+7v0nTZPtH4+lTEc1BC0Y7
px4gPgvWsFLmbOaZ8/STVdidmwdv8P/zEJhuG/c00p82/dD8r3d61oClsa2S
468akMbtiKKs2j/xkDsX5zsEYHaMTHTxSQDjXQk6+g7jXIcu1mPUETf8avXx
nhGzgdraex7Sgrjpbg+Y1FSeN1Wk68vbA855MrK0QTiw1e0d1ybzH96FTz7a
H0yOJO1zxaClf9sXqOdHAdrVRnUOdCH3aIUvnE6vIHdZ7cq/nTr47f+Ql5gW
vEnj6thimCnOqMp3s5oK6VHIZokg1kAubRikM1ReYPwzKJk3jWYG4/bnIxWa
ZhmtMZjTVYajZdN9HcLs0jhtxcSDp6ksx8n5ZLm2iWOtCjASN+WbyYP/RsnQ
BrcXYEukGYd64VxJUqscOPVtTbvwIP9VYerbgQb9VfHj4AjAEPaI9RxiI4Iw
uQsvbf40PSL2Rpu0CFt142dmHMCvB6j766tXE9gwY2uxwNOP41S4cpR0xykn
B/GvplFR+LmsijmT24EfXRSrmrCJpo8YTzSQm0HeuPqu4OIhV25+wNbmSYV/
QWKNRrNvDZi3izw3J5A41Q1VN5fokZGLvhqP5CESPgF9jx+2Sshab4EemEIF
Ju+mdA5C+dN+d39o9WyhXBkqP6YvUBFUTHzGh+OH2GBfvOga2vA6GiiY3ST9
5G9t6Zfmfz2o6AfPJiGQJJ0JWWxFm2YUTsz0aGcXN6FlLVxzvShZYreBERRP
UVhvPvU4ytvH6xuCie5+COs0IB4p32fkWvWL6/LD47T2J9lI2NW7V88Yd1Rw
PTK1TJS+YTOpKh/sAwwQxaNja2mtCpS/n6muZMfzfxecNIIV90WyyTSn599H
dzGjn23tFFWI7M6OobPlJKYSDlENY4thZaL1wGcRzI/RcbDf9pOSZlR7ELu1
NjxlQU0bRVxbBe/0Xb2xKG3x7Siu2BwwtFJxsf3wBFjHLHdw/NgWI+OQKiaX
DqyNLgvu+Y3soSZXPUw7Vy8rfoOdyfYZqKjV3zZ7uL7FJkKcie7cIfAZDTVG
g9leahuoUekKYh5PyH/lEUy1xKYj2UFFIearLX7KkqZi09oDl8ZEWrHziE3L
iEiKqwufAjyu4ypVDxbrzTbych9CkOUuPhGXzNZ/a56n0IUDLTG28BB883fl
4uWZSe9uSrkufw6q88G9AYWvE80l1NGqHPJvtaOyz6MuvnM/aiJdFYhm6V8u
P+A91WNiD/IETZfrMN/L/PVGdLugUYsthxxFCNcjYZqq0MDIKnkyKvHm6NQ3
RkzLocf3qj0oCxE9tdk8FuO393hZ1DE4v/2XupCo1j55xQmHUYuahRlU1PRD
RibzQEY4KArFgl4pe/VGyH6JC1GDnjuGHyzbuajWOcplP18j7hvITJsrI2c8
75IxGVldusMaNl2TLjOae2nP/RWOeEBlZkANE9EweLV6zHxLD8SM18162fTa
IF9kIyek/Nwa1PeiXhqOq7uEoT2/P0jNVv6unVcPPtAWekNFG2uIZYKInfnt
SWJ9YQF4guE55etjryO0pkYXqH7noQQT9kQ6MCZN3Vne2gwsDi9NC6ZdsUl5
fWPbLLf8qJnQPaOHuqwmE1w5JqbJs0GxfSLg5psazN6VP+cpCeJX9lLC6+kN
ToRwtPUBxznVJTW3FjBMNBv5SxSu6mIOxmmpd2/5sRSBDFxaHY+7gkAN3rQI
x8EZkBSVYMtXke582vj5cMVVYRrrZga2/owtJjG/HD1SSBiwYzMS/K+YeIJ/
5ommjg0+jGhbE2mQ/XwLYqrcIOLwln/LavymQ/u/rLEgfZgaXvSe01VXY76u
zHVd/viSi2YVwwKPAYJuPVt/e3Ya/sAxHHx6p0MSnX4q22yJcvxqUxxxSu4g
oPlXQSIQ36mkxT5CNDA1YwQO7E0HMRxhoyE/43ZfzeZRlUNUr0sbUgQs5tLx
x0E+0YWMmHazbaDSFEzufoavnS54ELWNcwQHqiXosIgvKzFtdNK12zdGIyFw
gQBG2zGEYesAMYyILdfbdNFpXYL36e105+7SHAgvy+O6oA9BzvJybhW3Q84x
h3eE6qb/8Ob+GDJJivtjU+EZdZlGBe2M5xNF14dOEapJ0k0zvt8dpM1NuO85
2Digt+KMW0lbicd8RtoKbjsWKG3jdafHkpTQWIg807Z+RVB4t/gel9+Nns6e
kLhOo7AzG8UahR/QddUTcR2Qg3ZKM6s/UvURoRHe45nIA1kxt67YTJUJ7hHP
yTagzEXkc/aFgNv6P0R+w9AuXB/R35hJXgHzMo4lYaoAlH/HiUniO9oFb6bG
uxdOZmq1VFwPT96H2DkHE+TBWRpxh7ZL+asn8RH6jVS8gFSXZGeL1lhIg7dq
IZaXVrdm/IEG3p6TDE9K/2xm7F0EHN02p/RAqpcoL4jhQzFfwmXj2x7hUvwn
lYAmd5deh4DOhWuAJhrKm4IqEiwKmM/7QJbsvX/IwL/MxPrs7ize0u3uqURl
6TJg/G3NYuE9YaOq1EsGDvCVoMhWAUbGioOji5q05G6BAeMjoepKLpCKjefj
0LD5mC/mvPmeov5OUQIgsObAlEsFvt4oUwgQ9C60uH48soF/+qMMyKJYVr54
w2PAq8fZlpfcg7QtAaG2Co119yJMAERgyKv0OBkl5+ncb9jvWQ+GQ9QH/1pF
j2ejS51bJyQlSuVgVKmVyfCEaUHT55yt3Vgt8kp2ftBPIBcTrO67J/yInJnU
fCcqcOibQ2iyMIttaTSsD+5HE4ihmtoS59o5gSaXh5uBbjQGHJzvb279WwLW
3YYhwpxUKwDQ3w1+RLEADS5y3q6y/VsHLuCxd2SFcmUGQhM0JmOAag7KEXTT
O+F8axr+0kJhy/Nzv5T3qm4vJKAsqzQHHWzcWx+BDrkeaB+4KF8Dvdb5A8AS
1MSbytI90M2Xtxd8OTPW3raSTVkLc3cZcJZ0vJVODuKYPRdM9J0F1XCvMWl/
cgKCTpprHQv4ub48csT+g8zuiqszDI4YE50rIxyOBAT6zb3vNT3dNU//bx35
rSt/lwt8A8p5+bAW3hwHgtBXAIeOXf+c+hbN641egbsFJA/PORyrsLIUS/6X
Njcd5F0spGLM0MPkrAAx1BPl7UngFK4dMQHjNZr7t+z8/zyMtrTdcwEDba6h
wJqOAaDmaXdugklfJlNhTgXY8/qyR/rgIj2dL7Ce0TKQD0FtkM2ZFqEsRMi4
kOnHm/o+uwvm+g4QXVN59W85KcmpPfFQ7El6Bl4NtGKFbQ8qWEHBw+PTuNKQ
w0cfuo03D5EioVFHVX5cuKlEnp7u/q8zFfxZoAPGoKWCidEG3C1tRu9g9hXn
vmnjEj7BPRLhTcklA/UnSHXHK9hNnroMToW7SL8KuGlKMH138hW8e4ohyhTj
GSSyvU2BcomI84TGwURHcHp1PuOIfUuJn8EQRpWcmGfqkDwGw4RnGmDF8z2a
ST9UxCAgv/ajFaDJ3lKtAkoryEcF6e9pfxz0mL7aCA0O/FDqXCycdoIthI8g
imhSptSvRr1kFLrvuWOCO0LB7jMrwh/q8YmY0nI+8UtEXwS3xp4JPYZRI2cf
Vvm0+07mq/C/RzaXEQovNHp6FTGp5wroHtGn0h5l+B1ti2FRfWAIHQAiBVoE
Ww2V/v8ZByBd5pc475CecTqC14r8msjHdgNSkl1Ji3C3sPugvDO9FYvkjdSL
Q1qZ9HvLNjciYh8x/KVHpfNmvuBNmwJHsPMqmKQb+2FLi5MiaTHyuFSby1R5
M15rYhVAk578j7c2zhEaUVWnTFlq23WvkRiFXtZtewBx0EXaQBQ73e5RLliX
H0HkNWyNk1DUrmBhhOLaH1ErwYm57k/j2fKBV1yN99hFINVxp/0nD5tNVK1S
08s7UUThisxeeT5vQ1mCfU8hRk/rYIzV6HG7MrOkQ6BkVEgOsz0rmAaygweO
Zs/tlLUej98FjWK1X0HwI3/NST5KD2m6/Bfoln0i2uSI4OyScXp/KF4Y2Aip
YJE7OuEpesFIiir2mailo81RXRNx+Yt9+OoWimOx7jWH+j9TptJghm75DEkI
FHq9W4noc6q0aHmpcVtJQsELPB8SxLL50LC6BijKscxlsaxq0yAmiyqdm2Eo
WIusmvrublsJWo+3xKa6rRwkIK/yj6gxkIllL3Boyp1VusOnzwQDeVR2wzj4
6UDaW7PrL/EGmsh2yHk8teFWSAI9VG9VcbW6PC23T3y3j9S4vla9QmGqKIKP
97Ytroq7d9pv0WF4/4SBxnZfOH2IIpGZAUsRcfBd5FNR60NQadEtmg55h47w
xEKMO9j8dWd8oOcrVjxB2U9FlmRpG1ZiqymZiqdJHuFE/6BX1Ytlrt8jz3zL
CotkBh76uLhpHZbbyJp75buzaHbPVrK6MAIYRhRsY95vn9f7Sk6sQkkO2lrc
Qn8IW5WFDdOZMtXDHPW8q75AuGboelo3E6P9GpqAsclJcZq+6DHZ1SJbhJM3
DY/YR0zKcoqUM5nzGp/YABzRoPle/byGU8t3D2VikAeCC6e/Y9590yRb1DbY
RQg5JPhglxxDQe3C+aPCASaeLy01YyoUN9YcJ8F3ZGVHHpkBjot9E7uJD3lc
KRFpmmMY+X/SGVXeSAwgLhaQV4tRl2WY4xcD3zIwaOzrFdBmX+gqq5rQpODh
Yaaj/P7LvIfK/iO/t2WIOui09b+ZwEbyvGe98rKWbVPpvUIkZP2ggAsYta0w
DTn+dmqCWT78L3LvSDJxEqOMgSbUs6w2NZsBk6e8B1GD1CJ3eTGfbhNM06pt
Xxz3FLgsOZvmNQB44Qccc+iWJ8M5jC6vlxHhriwLaV5+P7JcyR9IXAcFbN2y
42KV4f1fdc74/zL8f3d0C+WP7UtjURkBqH4Jg08GNqmU16NKga127Iy5qhaf
BGafDHh4YLH2aJs9dv3KAjZGshbdlBXf/RBbVYVpSgs3vY4u1Q2xWOrp81Pw
Rel2SyH4N8wLTc1dayfv/aIkVhc97SfhbDXmR00jqB9RkVgDkHQxyK5jIAnY
37pGHO8xvic92ZcSHL5Dh6vKn0CYxuvEei2v4HqMyfj90Pzkz0IQzqZmf+Ys
i9bVeX8X80DqT0pZPZv1jACus0O+RBOIv0XJzdWw+5vrkNbhK5Aiuf7AwHUk
KO84C515P3cMKX3Kr+hns/6XBS9ugqYlpXnCfuFoCJ6VBdpKZI2X5omXG8Vc
Gb4dvzlD36I0oFbIMfUjPnzADUfu1w6IoCZMaKA8nYpAA1RNlLGWFUuNr0iV
ozZ2ErJHArLItO4ofZE8KGfrJta/Bh8weUU4CYCMSSM+K9floPi0DronhmP8
fttAVgU1dgZjaJT3GMEI1SIYOPXqpuK/KafrVMo7jK5rO5t3d6KK0q2dKZN1
kW5LNyh292DSpFM+K/PwIU+n8HZEy2ob75e5drIWJ81LIX3inNxGnDDEri60
UY8BHU3gupKmVsFAirMdVURCXjoTTIESfgBCc+5CY1/41upnqjW6+0LCwgCa
1Oik7u4BFIFzw2sa3W6IHlqICPcf2U5w+PE3oOsd2/CzMghRegCui4I2gybS
QAn0QAOiksR7L0stbkZ36miSBNq2Ph/QAFxUqOAsyTsLqbKgW8vnNtF91FGt
5j4WkzEnmyvIdgSRQ3VdIJUkrAzfrOrCnDdF0hpL8vig70qXn3ellmVXBDzy
g5BF1kbepMeFTKEYNQs3Rq4DHJkEmsrbnYRGfJXQWQHCSmMZfBXTwCLv1CE/
vQu2REa6xMd5LL2Kc72BGHQ7NviAALecxZQQ2Ri3ltK3Vp75oIssLOAoa89d
se2IfFATs0kUJP7eeS4rSUN3jIcPD5CN2qY2ybDtbRVsuj06nwAeCD1GaBHH
/KvA60IMWPQdKQ2mqYhzSnNaxOnRZM2NZn0h6uDCQ32LOqs73VmbhovkBCUd
JjFYfF15xGWJ4RWRM5q0PeHO+znFwr2SDHTJ8CyqjEBNB653gKErTCzuyel3
ORAa5rCpIC1nMcW1aAUnlIKpstPukygdqnUHtTbuCYb2vkMyqQ6RzJO4jM2g
rpp5ktjHq8aMqfTOs2mF2Xx0LitDmk27CpHZi18mHw0V+gpyr8UJg3eYabn8
4xoiXPs14QlVzkgxUTNOIcTKBsazMR5Q+33xknN0U/K0XCe8xEmYWQnzU+1N
CohYRNI8uNbIrzo0eQmn9MrcQNC39pyCbDV4JqqwhqCffbpwjiK4lNW+C07N
HWiIpu6DqCK1EywiSHrbCzvtXdspTf1VRRy6a9xl0Dew/cgmmi31t86kCkRL
MQl9j7kzmyOL5GYog2Wz7y1TR5zMkMlGhDeTv14Tdhv4mehq6jJo8e+DC2kX
AkyPPePphCsEuWcmamP5Ep71avYfrV9H5i5BQAr6H0OUTtwp/OWHvBi1+hT8
aTlX8QrG0JWqb9oftfjudAXU2KCO6QtGSkq0jNKSVX8sBdycdIJQ+y786/Hx
BjV7K6yFojUVAA+50cjqcaBrwmdEh5uHxB07pQQWfXV65PXjdd7HUmwXewCE
Eifbuot3GDp/AJzQycziuc+xlpE2mtaipiCpdfJ6n57gcg7y7iVyIl3Mpkj6
i+BbsP+TD/XAoXJfNGiskry88YgVHWIAir9gewAy009ivfFBU8sIn6YxGsaN
JOnzUVAY6vsx+BpZ+UQPW1RFLIeM5gBKCfG/uvkWYPxQPpN17ekvBhBE7Gam
/MYvxoyLzMtWL6lwiAZ6EcT09ia7vuqisIUWBiM6FO0yg22g7WX2FoghVM2D
4HZPZJ1UazxqiWku9awaBWZ2hj+Er8mwrJvuU07qzxbqLoo4/AX6FNEU8ahm
OrVHUNXRIg0wcN261f6toFflE2leII7X1wKGf7N03UuatdE0DPSw9segPndU
hRTxUbn8GwOrUfOXbax3MSYgy/YO5DNdsRpwKhK7LC9D6+GxT7bBQPShK7vk
GJm0BoKpjAlZ2fI8VbRL2lvIuVPEnZ0OBUwQeEoO9vxBk6ctYDk46hLYdIRM
Rvv2PShtQBBr/JNtnWG+6JpUPF/yjtkFlXJlRz82yFzcNACjaqJMk9hurnVP
/oQJvmwz0l6a1hwt5XKCrnRB7YyCpQn/0S5LahWwMd5dW52PZW7DL+5l5j28
i/KmtCKRtdkBtH0PhpzcpV9JuCjTpJwd5PqZy5L+7dtL/AcXPyi1WCdRKtYJ
42zZILwYIj88kswtwdZczNxqXFapp5Ytb/j7Wt6pLXfWQcDySB3AylO/DGrL
+heM8fwyIp7BqTySvRbhGQDCWFgyNR+V92edhHOvKMQDehiltQYr2KNOkb+J
AdmrX06eNSt5QD51iBYafZB0YUntz8GS2F0oynn0L67UnL1ryvLAy5GiOPlK
JYj5b8yux/73BRHUduDRrWDSSJuHJLq5aZSGCe1ZzckKX8TsIr+ImthMyNbT
5TAVXr81h9jtH79i4e8QjbQITVLkfjXosTGsdEtL3UmqG4SNGNPF4CENPIKN
3jyuXQLGvq6tH5oHF/KsNHlb1lGfovHTXuJ3zUyflMzowJXVZqpFRZG91EfK
rAM30OdgdPr3mM52lW8qJX+J8FEM/FyiPh80BfGEp2HMbxkZzvrEJRSfFaNs
WdlvPsVpnuisuzO7/k4h19/6pOzr3A6XbnaTeAGgvY12LDuN3M0K8/i9nFtJ
USFrVNa/H0iuUVX3dkW5ktQrnu6fG9tz7mhVuJ4IuZnKbSUoOLchNCpogcHR
hNVaBUkPN1n0+uRQiiz3vzjnGRXocKjYMpwD9OQXv0veIcprFeFBP+qGrTle
XS9qLW8+7199QoeqEihhq0C3p1p1jc8DjPyJm89Rs3lRStLmNZbUdXVKHcWQ
goJhHoYcwLxLvfK+GvAQrjmrzmSPsJS9SE6SVfgMqODEtIE95QaKDyDTAVGg
qozLz9fs2cGytRiev8LsWHfBl44/NpSZzBFI508tCdymoTatPWiLQpAha5Jz
IENofiNsjFurP+/ARdjAZTMjMYrJY8H1zpEDe/Aa0iBo1k4wj72EC95G0TrV
7CdTVHnfgIbgQ8UqTDifUPZHRu2HQdd3Nq97qIjLxUTJ5AqBK7M78vHQmhUd
A5fWsCEA+JxsH6w+5fvMEGaiOu47uiEDABSZ7QQ1z3UMVHsrkVuDP36+tokX
DgBhGbqRWg0k4WPPSdxr/PqOSCscJrgkFh12J97y24MHbT9/nSHvCtij1X6B
w5Faxoa/ce0KcfjbuydKvcGe1m4fdeLxXvoUQmvXRBccAVJ3I5/12reRhJJm
6HRS0ix1pOau8+f9AAXS4347xeekqInHkjnjExWvFuEBA2u/On3lrxG4RYag
sWfmh3Unj6HIxz5weHcqg0e+Z1D++3Ht2Q29pOpGAGnLKR0nHvDxsvUPh0dx
/EE1gJhLpBAGzBgrLokVV18Yr4raIRjUsoRyPaB6EaOTEJLfOT/2CTjtB3o/
rVbRKgtCrKhXW9Q3j5zi1NSKBznyNWa+OtD563zWik/mRrbbyUYa2Mbo84CJ
D5BvWqUjWn73o2JDJPvM3FOYSDW5hQNsVnKSJDTStgu16ib2inm7CpibkLvP
lL89nqAM4LwiHEiEdRo12IfjNWp4BCtrYUvUChpJNGnjRO8OxF71rd07yZ2g
Q5JS7dwbi/nJwL9MANJhhZo3wjanoza7eBraNqIYl6aXpHcWqwrKiGhtt4on
XdjORXdOkb7aLx2FRmtd5AICA2E49ntRBC46DL3DLZNregCldb/QYA/q+7sQ
RUr0Ht1TTLXXzAyWFeKKroXaIKoEgNyQu8xDiCX7o343EnYhhGHiz2saTeBN
LUNEpMXQNoPrIdQOQNkhuApjoa/09yKh1Sk/srS8qadc2LYjgkTks8rkT+68
2ydUefgJ8gwU8/xOSUquTR1C/7OjRhH8vsQuDg+awq9kIy8IdWIXWWvwSSbm
QLxiR2xXoqxzx9ExyX/jJKdU3zzs87Wi3Qv1+YpXT4Au7KicNSjce8ESF0D9
jjCzW5y2CxUibs0r5QE2G94SRCYkXPStqlrE1Q9vFGF42pZhPBHVdxnyTJXL
nhUAzkQbqGAExGYgakAs/kn5odh5TMaDcA57rDkRELfNHPKnW+hH1I05cTEB
C9CI1W+6BPmYXEMyPJ8i2lU2RGUklweBR44IYghdUmjuJYBFiVB2CyscKb7B
dZ8TV48KqD8GZc1yfjU6UvErXetXgRJ/QDDG5k9IzVZyHIXVeGrqupgI0K99
Hw4tmTpmELsaAkpJS10y4DYAwG92gdD5I2ySgCO6ZTRdAtbtIRT9bkrFFWgm
yk21Ybjq8oq715EMM0ZhdpfVTF3kfayN1jWo5W3NsA1Fp5K42j3vQrPhn1Tv
ZOqHRUWKUGGkjV/+9Bu2vfGQAzjZp1m0yDiVwjHWbbUA36ceGvHLVQ/lV6j9
f9UVbqMaP/koj1CrOQp/xWjNTqemilyh3cmlc63Xmt/FTtn34aQnu7oybpPd
xJYI8xqq087CRrFUFMHsXQfmYDIUWMFZZWH11dSnO1uSz3+A4SLPEsX0Cz1o
nG28ErRn8W8nVs/X2n3iH9+WelWMvzWZyLyZ1IbULd0jZWPZXDTRD9QtjYEt
pdNsGbbp6pkMOCHOesbWZcRIWZU6mp8uLaW7nBPWoAXhHay7IXG0iMvdtXNY
Pnqx3VmjRtu2N8bIekEbdg/AjNVSp3bOTNtSBrClFM3EOfpYEKCoC3WdQymQ
FFezOaiecABPzSnkeDHoXrYeXXSpzlt5D+db4W6wcR4FlnkNz3oSzQrVBgA2
49qxlxEO1qke4k0RP2ORvWpmQkZBpPYr89oJYFCcgQsLNCz1kmfai7wXiXK1
1kV3dGR5dcdl1BUueBs22VQqLR+Lb50iDPgMLndfFXV71LoHzmjWX7tbXkh5
/MisYgNzgUDPvYd780wyRdcMpi35nh8shEfelbgsxsD/iOWs3JnNpR/av3Ff
Jo3RpltfwjKYOXPfKVSKg0uE/AeP66fpfHlBLkDhnQwkGlxNd8uPIrD8ihvb
+LkF+4cdk4v4UhaDv5hYdd8ZISuxaZ5jj+pN/IpBOHUkJc4N6B/LsgqEwKL4
DL4KUgYmt+jK/NKem2stYwUnITj07Xnu/fwH/1Ydp+aH4z4tk3dBQoj/0Dr5
pb2H6uaNsY2H3qUlpOiEOtS0HMvUHDQVxRwG5IMFteL2WOamiX+s63oODwFr
wSRxQG+aeEZBj+NjJogxwtigOh0r7SPyi4QrtDbxCHyuxnFXthl4siiS7xOX
bj7RnyJjE5nf+vOhTDiZVvqv0XpKaDQOrB/PyQU3cXoG3zh+eDzT7iWVpaDy
I3szIZ4XdhkVwpQFzvYqDMOP02VT9dwnWASkrFPrTXx+pPmcY3CqJC5/PV2O
D4G4w1uOFThvqsx8BglKCnZoikcmsFO1M1JyOVlk1iGztkTc3bUAVo6CWf40
FSqM7aYueOOC9TAz4yD7fMpOpZHg7PloQStyan7GODOYOoB5zRxDZkxzNYhh
STNfLe6HXvFYaaecMsN324KtmtUW+til5svYkvDNnvLiYU8apqQlH7tDn9T8
W0yjwx8xFYGf0HswmSkvF9l3mxxhHjJss5zr3pleLwdHHnRP/dcJlpX1NrM9
UqMx2q54pjYrfruW6Skz2zkj/ELyK7UMoSFHYAl8f1KLFZHbz0T44CdlqyFi
BjjMLx3YNzOmwmiV17lL77fUcmIYFmIZ6LeVxgcHpllvT3uyF11nz9PJPH1r
ckbIlxhKco82xtxSKWX8bUzBrNcbhl7ndk8OdmYllSNepEE6/UTkZmiikz60
rRVQA9sFwEZEVOrj6OM6iXGrGBqsC4r+MkiuvWfsv6Q4jTXTPnRDg2BB1cWP
hvEQXjyqz2kG719BelRbEek34BDhZyIRf7Wg3Sq5XyCfTQQUUo+DXWPn3dol
37IlR0bpTpWOPXwwN1CRANx9tyci08LavJVgHS5UPvsnk+xpGVe/GwgM7H2z
oDeTTxUZpjEOP6tjXysj+QjPpYn5dhq7iDM//TOvzKrfIzSqj9EKg7lltIwB
1vZUIR4bTPk0Lo04OehX+dxvrVEkRC7pGvV0UJWjMZhJ9WXZc7RAtdfand0X
QZIAUNidAHMf3U45o+lFyxsQ6W+F2it+wB6N7ktPFo4qh/ZeM/nu2zvPOOqH
0E6ncW/i1yRNzVBfBVW19OY+M69OVc5J2XA0+IGRPhxnKMAga00rfcLsb3PV
wXKI4OkhZmYfu4he+G+vXjpn8+Pjb1Z2H/F52jWI1yDUQqSIQRDVxvFwPLX6
+RQvG1Fwph0+pEmYX+nK8i6xG/TcVEVwIUZaT1HV955+8ijlFMj3ygLTIYG9
gL8wsS6cF6eKtTbo96umwskVATOU0g3wBJhXT7fpJDPz9FYMRXIJTLuo308m
FBM/NZy6z72kd3Lc8n9KzdDtztwPW1Tmafi90lTIgoM4xl0v3GIkKMF06kfY
Cr/v1dz3/NdkaQ6bwyi+Pt6ZeX4XYbN9Mcp9clN2WAtxcYvA058g96cS7fmN
HJR412CNbvKELDaZH9CxzTnqEsib841wEn56WJmPl8At3O8HyuGgLShzPyIz
2HgZKDKjedQ+1nuH+n3Y9GFIgRIgMiCTt6y2ixc2Jd4HhUhZZdkilNdFyf6H
XkdTS2O/XjvNzlubHKF0hCh3YPJBP/Z9XME0WG8MP1TwbjSzFBK3IukoouNq
bjBgQYnNbaIEgjF2gL2Ajn6HN+Ioo9869SwtF7IBlrtaLMvDX7H/gDnzZywC
rs4vBYv2URTEtSUduxZpwf9pAEWwoliMLCyycdyWcwCiKknoG8AnQyBt3XII
3AtJNQWpZhiNZbEABg9UmNJ4ByNqW7qOXvMVohObIzZoNtnuzHcNoQFK81b/
YVgH8dSu41b7G8sp5r26Avz06XzXobBCCKiZmJ6gJAYwYU9k3/5mDGJGdhgr
FMW6gInOyZOCF9DmZmjT9olSNx6ZraSm+X2qk0ncUUl+SRrH3/IaTqBWzfd0
iJAUIwr1dWkvQqIeyFg1WsPznCQfhDjPFYdsc/YnftiFl8aHYLRnURzaw98I
9TyZKJk055NG4hUkgtKi8zeJI1okvsRVzrejdq2SD3Zl1l+qgshA/nGyN9Ae
p0HBJJcP+hJ0E8rvylvyaLmWlgwdehvdYtCAEyg1oNT5jkbSp/3vbQQ/Tg0y
GO5y/cK4B2Tz53Xwv8BPKGNk9UplJ/5gwIx3wrXTkSPaMgu/6bjfLYTY/iQe
d1GB+crV8snoCAnepcVRxd9PZG2MdevOgq/QHORXlpoHrePvtL+fRGPitGH7
gilqPNe7DdFP9XfV27Z78QUTnmptVX5Me4blKvYEednZDLPvoiuWKR+DckZc
oPGOVXs0m8mg8svv2taUJPYz8Om5bu+z3u+kYUHV2/E8qn9UIYlTVzd2H06P
Ls9skNGY+sZCupOmLk9k2vP7AyazzBH+bRQk3R69XYzEWIsUXxfIPoTn12sr
p7nCRtcZbliHU+F/p5vv45PF+RcT+fgoc4X8tLSa+GJnqxQntdABLX/RzlHf
wF8ymPrEhePniaOEoKX/SuW2snmzrPKLi+Oqh6o4xyNpypu0HBnIFKiaYAZr
IA66JI0XBgvALcuzN6CarFp788E9hcC8QNGVFMTev90CzpufpWBID2prLdyq
2coAMV+LT0XlaVABhFHahFjFe2iLsIe6GdCLlSI3YGbbZ9SHER/5MG0CyZ/n
Kawm1xd7749qXr227t0kvy72lrScWRVd3PMYosBzHk2/n2gw2PDgIwJWbu6h
ZchHNwFV7SoA4HluEU4dRwjyvss4dTSIzrcP6f6cSypnNAQ1c9nOK9v2+d7W
bRURmqTQwjAxBwzppwbLn9xnc8jK007pkb63He//WMuidpFGngyJlkmqthy2
8o63jN6GHVlrvJI8+PzQRDVVunRBYF8Sz1SMTHtOrRb5/IK0U6xEbxqEP/gh
M6pe8HGE3fuj+FAQzk3gDlyQcRnSpaHfHDmA2bEyMv/48YOoctStwb667m6l
CRoUieXX047CnNI0xztrtNTRGEOFPuWl4rSkV91WHM1pAh2H4JlX71FSN4ak
0g3C3lsEyKRwrtWJlCGEPrQm3GvkWKCj8QaczH3Wmfng7qTqVJwFdmL3im2t
PLghZwro06IlxfgCk5ciknxbgZOLVhdtW5kVPcXM3GyijBCHVRiFVVD6pO3G
iHBFynT+oWrFRPd02gu050zIgOsNlrJ7xdJ2/QumNFDGdvbs4ndSbb0k39D0
CDj7oaCN/07pdXOj/vxjNa4qQ48xL5Gx6H01y07nP7bsiIqwvinEUWJxb2E4
hiezIFKOSxAkQCfNpKrkVYTM99MQiGua1d1lqunCq3fHi5lamXE+aTWDhqLi
sPSj4TUaE5n5FWKypKjO5RCYF997S4fPg/3AM+bjZ4TqAj7j884d3BBCcOxV
yNHYpDV/Kd9l8g1QucfAez/D3442GkOws3BI4NYDnN87x+dNX3D3P4TO9OSR
prToVT/WxFxswCqXSpqUCA3sROSU7jBZ0Kn2TD3Ugtklu0eCciriSOt2laiN
xK7qfTn60vBHNSP+P4v0Pq7PzbNrxsq1olN+XoZVxpDs5GZFoXv2pYBJ3sDz
Xxv/sGgnM6QD5xqXc15KSiyy34W4fOivnxfc9p0okaOxPRd3Yu7NKoc7NcmJ
cv5My5eStrsdGq1XFhpCagFe+83J0CAgjMrx/hHXwGWIfG93UM+KwNIWiMvL
64M0um0P9aCcIMBb8jyaJc3Y3+Otgjkl9m5tusOWv9iNRhEfOl5IUcfycQUf
lyIivG/FzrVy0dZP2csSKqNhxkMgov79ZuKnY3UFLDWLTMuwY7/pTThiOhcR
LXBq7+Ehyl6L2pc+rYDx1v8MNauygTzJ9da/YfpwqzlLmeaMxLEekRwRVW9B
Wsv7XNuch+rqRph+wSdy9zy5TVuwXp7EiRiMIx7ZN+bDQalnhQFaOxZuO0DQ
iai0TKLLJPgLZwefQuV3udynpgtXGVgxkGkhQPVHLKFmgQi++bikooG/HaiF
3NGYjx1Jq5UUV+58CaVnWR0UfCJJ79xrrTGuTMNQUCl3wr7eA4FaeIGb4m05
oFtfU8yOrL6D+U76HvGHwJPUNb+voM/V+UFOwU3pzCrgtjTK2HKx9B9Cw3/N
H6HyBsP9Buidzokaie64d7k3KaRMWftiRfL6R1GxYxivkv8r+Fh/xsvTHeU/
VxLtuvX3B6IBtoHuBA/kPI5BtXias+OEpXdJQnjPAZnIQLyaSF3fbEpvVju4
1nBPyV6qPGwSaTaOHrbR1hG0Py6ePT/2xoBKcs2ZgSfj3p4KYzzzfUDxfqXv
d5zrDXZPEzb584MWBe8tCntdtXeEnRgZn8/9Zx5O73v9tbMOBuSOyc3H+EjP
ySeYGkjRDpFEOHm3DNAVhSfjmxnCoZinzxZvfhPnvt2H4NkA2p5Adfl5Drbv
035+zTCX5q/Mr2x5UG15mS6bebhDX0XFP6HcZ6h9NMq/986DMooFmMvuIb0c
0Mzcq18IUFZRFFXC5kDpCF1NqsE9oFr2hYt0qpF/8M+/E4jxMbm6l/HXW0tD
gcNPn2ntCSB3Hi6TxPG6Vo+2jMy8QWgAZ54tbxfT0h5bMgS0LQvJsa0dKowX
1yGWN791bLFKfulYwgnCRcqHt2DpfrWQSubX+00EbcxpvFfHg9DvowD6XQN1
key23Zky62CwUnzNEa0EWnlrQD//gqP5hsrp38dVZ2hPxvHY/zmu3i9rbYj3
bydC0AucrH35D2uudYPWL/wwvW+MzTanwx7qLpvFrx0+rDcGG5MDaQ2c5yrN
2GRLtmxPWR6WDLVgKytWx+CzcOC/CVHBWmSM1VpN954Gzh//4qSdgbGXtG0O
UNrm0mgaS1EM9xPkauylcuHqFT3ao2sUV187J6JnCo3wxa+J0uP8EikQz+2j
J2hUg4cLmk/62FyVeYcDT7iHQIuW2YpwlQ94L9ba8sHua+xwqx5bXaN5tqhZ
kfUQ4U2/SxRVti0Yb884JCG8bqN7v6eyeqGrMqsmgDCaGat3ad3XccWCSQ/B
BhEoSLm6bQdx/XBQW2SXPjKyNYBIp7U0+eSpTjp38W10Vh+DuSM01HbMwvVK
Qm26moZnfTeb8OQPraCNSh3bIMrM0PtNNAudID/qB5UrN52Z7IlUC0ekmnDZ
hRv2MdhRROQHa5s+Tb5Du7EIvtCBz4Pq2G+1DndXa9maPXnnhThA1NCvLWPY
lCWjUtRfWvCG4ZHw+5jw3/Y+ZXTMD6mQUK64NnlXNCz+4jeHjnyYWihCU7sH
H4vlxBWSVOvizRBdyaZ66JWbTPBObQFm0mu/8an+EmW/qtHXHJIE/0EFSypF
5Q52I+b8bF1cWyA4CoK7aV8F2hoHqQOM9tMXWaS5wmm2kc623R1LGF/sdJZ+
dKHvmt8hmCMnw+/XNmXesUZpf3GnSJdYtkRY/riYombVRM/ePct6R/Gud6QM
iVaQcsKIqytGxH6DSWEYuEyI3fqK1aWeikR6CV3G1xdiXkmQT7WscyUdGaMU
cBV7QizP76IpbWvy+TiHn+qUVAOOSOylkiBSmVw0jGuc3qeOgNeUZ+2OH0mF
w9Z4/8CqwNCCceo0RkWNllvrBz5l3mLNRSm1KwdPYbculE9IQ46jMm5EswYZ
046XWCNrnt2qOiF2/jn7XNIemlHUb9JLgxAGJUg76rOyURTMYxyavEmUvjvB
VIS65wi9NMzQpvJH2O7cBGwi60tnaf1XTtlDQI+WCcHn6lU+jTIxHpdnhx2+
kuSmgJUKjyklvPLjGVLikS0TSrXvNRkHIRr6eU2HDlFiWXKSCR8y8+azmLG7
P+l6hJrsFOAqp2cFXCQWjk0a1kE9/G9D9MyvPiHa2XcDIFrXKCGE65pTfcNo
HJfJ9Nf8DT+vwPwt/PuTcZhspJURFhnouA/2blfQMGhZDHd4DsnCDygVleCF
Hs66DTYxkCAsTQU0AmA6A+t6VHME+jwwS5RF0Ub++mq8ZEsDj1z9WpXQNSPZ
S+q0dNpR2Zqms8DASkg7OB5s8ElQ9wRojQmUlxTmFfaV9B5mIJqUASo8ZWYL
2oUltKTOjtR4Ai7+m6Fj5J/cJO29q3uIHELhP/4AhiKjk1d2GKhS+Ywot78D
VpuaLXGywHoXDM8baEVlPk2ZlPSQ1g9oTgm7T6ztgag11UT/UlF14a7X2pPj
DGelDKARB+OocqAF0dfDUmFF2DWesCAAKyd+niLPODQYeOQ3kw8Q25DwqCS3
nenFH78ziJqtUiwH6iq2SkbEmVfX6whvmA9MRMHsq+anorQBWoBaljXJiM/e
oghdzNsylyHzkI8DbhZRp/rOkBXx0ASwVrvPdOkhmi6DJc3ECzm+fob0DUT6
NUmO2JvIyYrJaD1sNdrL0LGIKOMka2b4XisuD9BT5Z29a0ttz7E+S/DxpKCG
YEeenDtDpOAwixCrJB1AqtxfxrQyuEq8D/zqZrAPBhv0HEx9taeLSuB7qoh7
B+jLFlRnuGn3c66ha0eko0EW9WUzfWyR6JA1fV6IwsXHAswkkIkhl4QuZhdK
5SviNMejsHlPjY0FFk3wcEzVs8KyVJZG06j2oJ1M1Uh9DRDxgTNBxEpPe8uW
v7tr2PkB5Mgdqs4c5X+Eh6Ypiy1DFCPAuMFUvEOD3hL2Jz/ygVrXu0iYaLuD
1lMHyspyA4LSqN5dOhMVqyS9ZJvep2DRYnV/SY2mPAcPQ0/bDm29xP2AwssQ
YGoByl77xmPih+ZDNSDDz2Y8kxwGYWks/9+7wlzE9oMhVbExDR114qne6By1
tcUg84O1BrROFc1/cDzOiiRoFjNLMcNVECc4u13oDEQJO25/n0JJerHHDNeI
YonfXjGuv23+b5rlhTKIrzP1kEfwo9Ul0AUCqv1EZUqGaAfpr/6II+Do49oo
os1tiVA1m8CKVh4N6U2HG+8pDx0/k4mGggaBNdicfbrLuotJxINAF4eUijUb
q3Yaf0yjpyTA12oqMGZP6PVC1UA8aMu64Ej62h8n4ZQyo5bi/fxHzpoGzkdI
SGw+fHQCPkUbZ8Jx+FxurNx/b8znlFOVs8yR1KaKvG0rn5xgDbAx7sOo/I79
nTyQtpmHkcZsKv0EfmOVZoew/CLaLE+2CzKTf9dU6EG5omEKl7+CxGUTRoeF
cUXxUkQIz7+hSYlCZa0+ZIwlcgcKZJ/IV8dWA4s6dY4oTuX0elJD5DOdr9Ux
XGzivT0lOuZhHRS/drWLX/pU4Ir9P8PsCclCQ6OdlvlUOCAhd0Y8lWBAFcFX
SwKn4VkUtVVpexQ4Mmz6aQHt43PqAYfwDYNqo1lp2zRhhwfeHTHYjm8OjX3w
90AgHi4dfjxGkBeG1Yrl9gwdzvbsCO2IrJqojRnwyvipoQB7Qm8CI69pW9pO
9UZi65Y4EHsxbNTyF4450LS9WNWPrRxEIfZERGFs5pzHRAUBMoMk8d9PZa/q
YUSNHBx3S9w8ApqDMPSzmFSjsdwPPQTV/btJhJnSbnxnJmNXaeuGvjDHIGYd
pwQPW6pHQOAVE68qAiGfMvszJ7X1xw4227r4LIodFYXe0x5+5/Kuafw7+M7c
DDsWrxR++CVxoDN6/Uk/JD9VjJIwnlRMNDzVv90QX49LekXuqoc8Q/4cN/ES
bMlK98N1U46X393/SXnPd/9Y+Arb2hleZS6yFvDl/VltSpvuextG+Ry5047w
+MTjx5Ts6Ze0S1UyPqGVkcX+VMXzaFF9EH/SqUm1Bj5zLY04PQJHomPe3io9
BRGtFdbAD0of+9iudB4zf5bGwLWfZ9DeCmBeL5ZdOmd4d9dSieU8gElyrsME
GPb41Yh4+RQJCv+roZrldyrUTh1SM+BO0DZfTk/aIODUxclbDUjewUQVdYsy
+9Gfj9Yupz5p0J3L/q8E8mJk6AnnjDOItLRXntjjXBim82BbtrEJXZdMWVL9
34lG9jGIl56S+lhFRPzqmO3Dsf2EfdLTLmbck4fqcQImF2zoMYhnvAN8cqt6
VAIfyNqE55jkZ4qaLl0gXSnEed7dIBN7RrXfKMLJ2AgkAEWb7/dVmn5EpuJy
+zWt7o1zImXqf3t9Le70rQO6KZVqYLDZf1A5C0rPYFJk8hIVXk49fIVY4+RC
Aucq+0hFz4oPQj0zS2VhCwEJs27AvQQuUkma0rt9gfirjhRBqKdn6L+0MnzY
0HScvsiNFL+9fLqo/KB8Mo1nDf0/HrMtUXO3C24DkcsXao3/oDvjYbsXILLl
kE5dO4oxkQKaGfQeI/obYRxzbd031Zpe+xdDrLwEFLtoP1xThgxPXS2RPNSz
JbvUV34SyYYlWcFHlIzJFqfBKmlA7M78g9hvL3Li7U8SUG3gCF9iIOSdOn+X
uimK30VygWlvfER70NEfDgYQXwerv95fhgLZv1jVXCOitxXDIO8p3WOhIWeq
fS4dLNC+qq94bljYJTfvXPHWfv2Y+/y9/Ewgi6ynliQiOmXnYDv/FgcsUUCF
ssI6u/ATjtdAOaa9wWS4zlGIdui9y6jL+kldKuHcx64+o74uMvhGSULzZJ4y
5qjRTPxcdGrwo0ROIRxlXSZPRMZPheCUdXqbn9CutYPbyCQhdseMCbPXl37j
V0Apj6tblaNBookU1ZeUvDWN1UdcpcY4yyOFfM5/bc5cAk0vPKWVIvJRcy9e
+UFUo11QcvDWu49CkDFpFKjFqop8qjruQcU2L4dL/Fw0gUUM1TXwP3ztsenT
dXK7rsWtdBpbPLP1x7VcUb6P2KAwUUVZdNsCx2avDzolMAaOaDQibUAecXJ6
ac37c8R/oQs5aU6K+8q9SWj+RfFmvBKd7I9y7RM7wuWLn8X0Ur8zRAW+uQh9
JAoN54ha7rhrWrytZQE9XoI+Vwm2FptjwrFdddGLKZd69g/+sfRCZu0UFrak
/IlXFcljAoht2g2pGpQFNWsW1KmSc7N/g74xPm5ZUdXESMaBDeseURHftesm
vrVKVJiJKIfZcYYPr+AoJGu33h9ihZWH454JvH6s/eNV/mr6U3ijr/JOJGZp
XtwjpfqjGs1D2ds9Tl0Z7LK/eJudWZP1wxlLodZ2ZaUNoCXbemWS50aVkUNj
ko+q94jEwAsXEWZ1TDKE0WpYjj3JBcerQfaM3AUHF8Y0kkhCMOkgkzu0sDhy
fFtqZyOKA1iKTiNZXH3jr+un35e6pNIwOmEqyN5bYXCUEuBMCsFzmtiMVCy3
a3J3Vo6kQYYVrED27vaFXj1Gv72JcMnsm60ipeKU7s35W8ODWNWXoKvivJ3l
nUSdeJ5qWz+VJM63euzPIog8UdQmRkVBIT2vrkgYAhr6Ik2ufrEMJfBvPA9p
MeV3iVozgeO/VLzt4QxR+eAyytjyrfdCefDlJYWXw5LZnkvDuJ9xt3bS8tQg
ZuDdOtAQNEBGQZKTcMJojRZ7GPXduOooRH6TsGdDUKKeZdvyRM1oeNNkiIs5
ykOWxfdSjhAeQ8he0a312bSE0j897b3QTUHWiSPRILkcUPFTx8QVuPelQIJh
09qm8eI7VKf8zNdA6uIxJJTU3iQImJSnTzieAg8TTQNkrQyVQduJlDPn43sa
7dLYwzsumX/CZH8N9dsWG5FVkeI1UZQfhyL+dMgZ9Q6/cy7JBn7a0+6Sky+b
RHaB+giHF1Z6cjko3OFIJB7dJ7vsQoKTYwsD+1On2cmND7f4eXZ1H6bXJWc+
5d/0LsZccq8xVfQFrNrmCCyIpwbxsUS2iTEn3QNbahQ7k7aX9EZPvJ9FuzPr
kTw6ApUbxo49Ilb5wfS0YPmsvZgrxQR/PSHz/xEnwVfX6KgZA8uIIa41IwmW
TtC4NgjlEgP8x2DOlcHejHoMRSA/Oc1YXOPlDxLWSzACdo3ncrYTzPNKgifl
l36YnHTt9CNACVzddgQVoi8f6qSBebuKqmPG8yh/yP1t4Ow4XX9ndT9NnLN5
iYw6m/yLxs+6Y01O+ZYvcvthEI1MX5mF66YcYE/Z+0REG2Hwan5Mu6mVQVmH
U9HXguC6sWkvnYdkpMwdsMX34ulIchp6ZC1RMANXlcW+/Djgux/hiAD1nrVt
c7eSrWfV3xOwgS5nPJ2meoGLCx1z+OdQWfMHLhvV7k9+GJrGakQxTiTrgcZS
bopDCZSGnMHLyHdU76yy+nRyi78C7DVwC7BVpMe6Y0DdP78BPYJ9bQjjKXni
WbVLRFAvtzCFLl72cPUuSZaw4Kh5AJqRVbAZvtPIdUrSxBc2e3bMCHCmdoRI
+PCBjQ1G3Xyo7/NzLhH6kicYzHFA1ce14MlX8fL71DCUupKngx3jtb49yuCH
0ym6KUQjkp6kKltPQ7+wy3MrlfcaWSHApCfUGL+e8qYa/S1vBoZ5D0fILfhh
ZIS3ILGYBmlyqRT9Pe7aR6KzVLcfAMyGrMG0rBXef21QnBaM1+jI5s8udBA9
AJKgYHJMBptIFb6OPDkU4kYNT29NzUBMQmv8JWv0C4d4NDdoCqii+PTM56bj
2R69ypQivbzXc9bM/4NW/fmzk6PS6puUNgw+s8z+vFhdHIVMXNTjMV+vAgtb
QkT3S+23DiRnPb/zidrx/HlH+F5V1LpsUU0vdjwRQh8uuoCDcmERKlQs6hCX
Yf6haZt1DIqlpc6qrTnercTSop+KaUWgJyTmpbt8gbni50N5sBKyPXcdeawG
T27ZayL9CIejs06P45DQ/JL/xlu7GTpJlnBq+QLbPMx3t0Ah2usL1aJ3VyCB
V7nVw/iXcVBYlk3+AA6EyK0wToaXhJqrnl454+iY43UotyIlp2ndVPd/BMzu
guLNY9RPlRPJeIBq+ZpzA+Fsb90cEbN31zhuz8r6jrof2qPlFCrT063zN8f3
fJPNd40jbJZVr1UuyPuf53guZMEsFctCIHCIeAxBFCpzQEwS2vj+vWIiugT1
Xwud2sSc8kiufflR+qhFUQINwD/61WtEfrEdY1nQkLYeS0LKOAmHUCAxuoZQ
jcxkuY/+NxyXQx8vsVJbJX6YFPNJcuoyLJ5oSLgMEDYlMJNCjXSDcmVE2SLz
djti+LVbocDaWP2452weLvnJJgS4flq23ke8C7pgbGTFOFL/jhAC+Cgd2/nO
vudiQEQf4Swpzx3hGMIzzxFEGdSNzxccPjkJoKlzD4JzXRuxl4HnKzdKqauD
shnGKIicGv5Pcgp/uyqFtYSdfynvIETLBmDDGItHmE4pU7bJTZ98JZQAMcZr
4BNZQ+2HRpRBS0JjJ890I2G4347LHO1iAnjx+kFw52bic+QBTe1xrVSs+rMD
imMoNhUdwsnqXeclZ6PQcMxDR0fgdwwl9zmt9iGYiDltwy4SboAIbc+4uVKa
/9YEiRoxG5rk5tzMGua4V2UE15QtBbdww9jQ1I/LrK0Uo6AaHo0w0vW9bVCq
DloBIbbv8UPTFvWGZIZsB+DHbxENQD0TH4bwbVMxU8zg3HsYst3AyfCguBOt
mLPEfDJwXNkPOrbp+e99XVQqbkZ8p0k5C2CeVWm+yLYWd8EjFFawBxhXW8z1
mNq1IzTsUbtFQetpJ5Lrdau10/P1k3ceK2BdTSqe4CQnB0mvtTpaLYkXwbZr
K7Mx7d2gZiuKsAD3XUhhsvWbOz4jdXRlKtxXtjLEoyzKgZvcD9sJSkHXr/d/
eh1+k1v3Xk+MRT9dANyEQjpKBIx4m1LFRneR0whdWjo4wzPNSK7iv3uyOtft
HVnK/2uph/8z8EpdvR+yv0NBgHAZZ8/S4VBtaA0RdLFy5Ttq+UA4ZlLfELlO
6mOq1VveoHWravht2Kzd9Qwco+nTQcqthw8mUGSIDSc4ELBXNo4i/cQooQ7o
Gf0bWU0135ch4BJnB7y63l9NK5rk6tjV7akb1hwk/P7tXFOKEXuPno7wrNBo
1XKvluqoEx1DbXP3asuC+CLd7rJwp5dP4qsq7pd5PyBxX2OIKUYuAku5dBMK
ld8ehzp7rm7GC21X7aoFYg7RGQNMDFjvt/pPEVvUpvU1GsrrVAE6a9dOdYWc
Y4J/vB08TfnvcCWek0OgJsqvSStUl5iz2ko5l52l1QQyTOnVhS4SDOGiVX+w
x6e+Oc3eoEvJEmXN0FTi7T2PPE44bkPqSjluC2pLMdxk1ChYr5ANIKj/4ZZN
kJizJvjYaywhI1bZAEWPMLj21tiKrMFPduaCafBY4E1vqq/5ekzZkF2Ye6pk
5G0U/VDhPTQnqWmFczSZnkRQS9+bGw4D5hFLHc47QeyZc7CStg0khXAfQ/EM
Abyok1rwP4L0nKaB0UfAzlsLSyKhAZQK9HII968Vwp7Hxvqz2ibnDWHZtaE3
uiJ698SUZ+XHo2JTT8SijAnPoZgVmVPyTw2mqdDQNFg3eVARwsdIYkoeMP4A
wcYQhhsh8eUN3LkzvgX+1b+/OEkbUIx/OgnseYq0FzQDHap3KyCAz1sHkFa5
jrl6UsMD31zjK6PwQISQtTMSHlIfpeBmPYlxb/SEV3W3/fefDjnk1z4qoQw4
HyLuKn7HJFmkppUBDLxxZkEAa7L7jnxSL5KYkgS12pr6kihZrEefVYix6sty
YTWGRO+MvEklNj+V5im7O0T++StZFjAAKizA1qxFDVEHPcPXEPinxHpa8gPR
a3n2JMuGVa6a2NB9UEr+L+Qqew7wX0Jzuv9I2+btikbqnYqbAbeJ0oKO9c1c
bh7uzSyQZhL9/9DnsDPTJERflpv30jb7XIhYLZVQl7c46xtFMAprOvsD1pLK
ln6SgITY5oevDnvVBKdwxwD5YeqHddIY5sHW7s93qtManxWILFuXvxwd8Qve
t54QEqbtOknmpXGaVBcJrfnPyq8DaISOO7707xCbTcxDgHIlOgjzxQMkBzaw
rqeP8ybIkWu50AvJDgo4XszvQ2GD6xmuLwgQTjVLCWYX1CpR//n0wgKeqI93
EG/2UwSMjEvqbPI34Wbnob06vmcBA/IhAzFcXriEHIKpz6AkefWxfObeUuy4
q7ZPtKQS6FCUEQtsST989A+MVUXQLlDPyfyx7Rovn6ssbTpskN+CRY6poTtB
IUQFeSraL0CULEk5f3oNLZmLrTydL8ge29L2LSF+cBmB5J/778nlvUbcJL/J
zCbd8dJm9R8biniuLFVaSVCafh6tyPcCHmj7haMqRQ9BoEvqxM04SraKNvW+
9mpZB0wMSdHly5lQ9L1CGOwtsqvKs6sceFIN1xLG9l3YwhPlRx8ApSpNDQoi
CPfw/WpNtGk4bFdD0W8l/RCLJfFpZ7ajfTp08X4svV47yzUiQ9AaPzEEtdR0
Nd1OFnPrW9DGqDB7iX64zHv/6rl2noVD318iHsSVhHjtAIQCkNwcAq0HrsLe
eLCF2l0oclFFwLm+5fHjZF6POJtD7tuGMitOGwprfhxLQVZioo0+NEF/s6As
7ByExvT2C9t/7b9LeHuqdKL0JqXHAE9GB79HSK1huousLAVMdvJ3sCR7cEz9
a9OiWJ826c8i9yhC/195CFQK+HFXbRz3vlbC+SZKZnTjSy+1GDVyseCIVSn4
pBHUg3vWuwwcrK+u3XqpyVzVqzavf8DRMGc3n9LEPNnScpoU8j4gS5LYWFGW
Apj/3poTC8txHn/3Mfy9YT0t4tuW0l5wJxETx7GBbk67YAEQ0oEUAUIbOuiP
CfFxln/hBa75XDbIZtz3ciXnJwUCBdXhZXBvk+9qQdEoFtOml6HsnX4mORuW
FjsUKsE+FgG4o7iYxzXxUzd++2PiVC6utA3qaj0R7Uv/rpL06FgusCoAX0Kt
3AjPrYPYOjwxOMHZYYa9nd/fQJ68i2I2/QR53RaoJAyz8rCZC9SQcKKBoMaC
45vjiOiCcfEelTskNMep7gVr71vzBZCy9vvv7QyGRNIAV5/7jmuVl9369uda
iDC3YesnOFitxWvX/mQ/dD9Fw7FpAWgKjceEZ9FJB8F6lFx+S5j6lfbdGQ0U
0WG+zR8JbY2JcNqr1ZUZTibx8+qRWXuV1u6vnZj8DCCvGb2Uu4IhL0k/qauS
HCOU8euyzCb0TOxhHlmikBcOjjCCEDpl9ymU73dMgBfDI3TcyFK1rARGS71k
BtryNrnveKZtc/SCPQSAl4siJisfTQlgScM7SAxdIJQt+AXrdeSq9aK8bXy2
x42v3/rVOZ50CXSi6KakFLKvl0gTIHkX4PcgnlWWMPRtM/Qnd4QTUSJkM+o1
NY4HzghfikRdu5AWANwJKkfr1RLj9jXqi6v2r1hDOk124svgkhT+VsiMwTpK
149MD1OJeuCg4ITb0os1UVpGJJFMWBfApG0XOOQPL96e1vRd4s+mJvEP6xi2
qr/pasAsEBgR6R/mbVba+pYhxlBQ7Un9PYlCFU6JV9hUby3j6fO/uXWoDULT
B6PJ9FGr/76w10hO517K2voD1BCqf4j5jh/JoJbX9Ufh7h+uVMErrq8dgeE/
+Rc9yA6s5ByVpamgTxUoRP/Mz5sdaj/cC2q6IYvMai8BxlKezGIAkdLnj85e
B3lWYJuLWj60nhxg3sdCUZJaNs6B1zpCUn+KvAQiOmUNxP35eFCbYGFX1dkp
DvrFv8j5F9vZLfsiIeOrvfFRbUHg3+Hk0itjNDYHgaBT3VJuoy7hZH4dD8/V
Qs8cXG0hK2W5VT2WqScVyREGZg6raG4oMit7xi/zJl9TtISE556b0IQC1ujz
Ou/SJTg1A6tfPSHGP8Ao13qiPufN7te9Q2QDJ4Gkd6gUEYoBzeFIfcS+7J5I
Lkfe8HLmfG8Zd9hJKVtcRijUEaJTY4aW2t1eSrm5sCyFrFp9wemplho/nP3h
cBFnc03hIrEZ591b0fVgse+mzvbfZo8zLfOdnaL9J69CNZM0rZkNx21lAWn4
WIh+Xqd8IPPPWNSZgL0eZmcYx5Krr57zqRcpVnvZfI/A3UrXFQOYpb3Nngwu
3eCvic040+wQjZ0ZIvwCTHqr2dWh2Rqd/h54y1JJCgpk0rynuf8tMqymiBNv
QzPXi0SC27G5pIlcXgoyvmhRvV47cAh+GRZbbnkTzGqjgF7/O4HMNNLE4RCv
Gv/OsZf7edYmu+Tbuz1+HXvS0B4QIRmtohis0gz4ub8KXOm5hwFsB2dDNxv1
XKp7upWOlPxeBYV8HEBZkueRI0QPkdGXGa+jYG5QogobtL1Igz8rUIJ3dQRv
a6wYIPrYyBRBDEzRZfr52TIg9TyQclOnIiKGbqaPTuTyf7JzT5yLmeSSjfoV
0RF2L+I3uNOqCMjBEshLH/JBnD7nK1ariELQP3n8mRHjj1wKPGGeqVxIqpLM
dROfQ7V1rhb84bHR/QJ3elni7Urq4N308EMnnWVH1Ax9CXvIDIYW6ZU9NHad
Yd0AZ3rIG4PNaTDM75G5YJuoxT/xrXOw0XCzOXBcV/Han7ADCYZqP8FQE/Mn
jDxiuMiUJeM1lTx+NL21ExzJQp/wdFGrL9rNmHLSN+aAsBZ3DtNbExKqTQJW
OlKqFZ9h2R0ZmKdaDCs8VHUT6rZ7P3MIIdy8waTpAiGL+21uhtppvBRva+JD
hn4++gLivqrZR9ouiUtNbeAwVOHT26gZrSIm+IdYpNe20UHuJkvLuVHbcUIp
Otz2S7jc023aTP3FcKp3OsBj26xoqRLymHkfpgT5VzYS9K1qM3drTeaLaqsM
O7yCxDtBJncPk/cY5f7Ew5s6GJz9aHWMW9/Zp2O1gZFBGBMnF+QcjooAa3lo
opf3wQ8a2xOmdC7g4erGQbFb9qI1WyMRGtwxC3q+j1be9MDNjPSSuqhht7k0
P5rcdPukWPd3OGpuMxtz4TJo4m4WVX1Nfkl9ipqLl696py6St2hn+CQt0ryA
ZdNqF/rzdO3V9qMet/cWkPyBfTtRjSh5k8njjxlmv9yZLxgqDjQRerRiVKiE
Z8YLypvRKgpjyKFEt9Y6sLfqVaviCzI3Cl+b0S1xQ8iFy1zQAYEIfpLYpDeJ
p4EQqfwX9/BOqctus2VPBzmBuYSW4Lr2WXxwK+VQUcPnXqwjLCXcjoXXhund
+RPISLL2pIBhtkVt2Nl587dxe4gjiuJzwgipLQ6+1qz1pHrqK6X2DaTiaDD0
QTP2Fe0k6+f1yzL+nHRov39v+BtDNV4dSp61yZfdTffa3365Cmi5L6wIH3O7
lhebbfVb9YE2C+AW0iRJkRUrrCq0a8kwiFR09dUHiZol7mpIxUqa01WT7RW2
huhOy9ILPQqFJSp1NBwet2uFKsOonQlLvvxHa5c3vOx1g4zsrUHomsvb1sN5
RIt58WdbYWebvyF2YqhjYfEfIvAvLW/0MT5s6vpF3nPF/9sMcPVP50uDwDj4
BJfhTtIsR6FlN+9i49ESautAnXF/en45govCwKnmkr41aVQy8hLKMNZNUGUg
d/qZ2a12bKMJ3N1sbYrReAR7cVW0+ZATItXkXTZCcCHlpLfwwiWVIG/zmmBL
n80//assI6ounfKF00FtqKUlPRvwqDamU6VyGTxTb3/4TitXiqCwQFn+Yfld
nlOACbLfmANjnNoiMtbJxrqb9o0BvGQ6fosbpyOf38aNYBtttCGYF1vm1BXJ
zkOOKsVuijaotgV9XiJrRRl0dfgwv794th4OtSgqY9I32fegWJL4//WuukUR
CxGfTViw2HutjCtj97DaHT3A3s2MAEkfn1OhEiA5uIdN8cUF9K17Q8cjhzhf
7BOF+EdpABitbdUFWUfqUZAUmo62abXt0hyZ+SYoET+YpUV8t4nlyN40ewYZ
qypYtgbIo5XUjgE4NfsEWtw0hDHysfJS1YpLGgm0Q9886Qg2mKeeQARtbsH5
dkU5Okl7elroIjX9btGvbsqJ+JeuTSKeeOXIWbNUXqAxFUsge4qroL15HqgJ
BU+QLX37eDi3ZZ+vyird1sWNSoatRjc8R20GiNRBXNTzrWuO4nG5E7qvVsJl
l/8sd7wsXlMm0mIRxOHuxvKqAZ3Z5kRyi2tSOyxeePtgF6aNxr5OXT0Dogta
JD2xxBG1/xxLsLiTfv5hugdKvANKtmzmOoOqsfWj59Lg8myudZiVDbWw3pRI
dGVJ7AMMp9Oo0XZqARGLKY1odAyBMcwNFNKpkiWH75ZCsr1A8A6xGV7rR/xm
zX+Ra6zxZ0TNjrs49Pc3v31mM2YJKqVH+ZQowF4DrP/FsIVt3s5jXHJNyz6I
JFh0qfohkTsEvY4vYHAmshHx1QAhz8YZT3TcUX+rpfsPlYG+9Gi2Xdmbj9JD
VfzkqjZKogTG8FhVmQcFcXDo3tPS9UnUhQs4ImuQyPWdVxw9gFY/wR4VRkr4
tY9kBo/WGb18CGEBzSrIoEvfoI4A2c5wYHIQdI0C/FsKjSDrgRvRJ6ghy/tN
MKj+eMD1hbQR+8nOyXuE093Q1tw/GKgIBBVZwUu/S+o/KHMm85xCLxitISrS
CErZ3ikm3VR2JMPgbG9VWUfP6/k2NPpdmdLZSytuS4G+w43Pjrc3ywD7yKnK
TYp/xr9eis2P0Tj4IB0XOmy2KIk8HsphqrrmF49jWIu1m4wfOKaR0m0QkHot
ILYML5Knb92jMfS8Qk4tv6YEgkaRlwkWT6/sqt0LrQjLihihb5R+oAtTrbWq
ozAOoLwr8Fo99WDh+cJrRNh5uM1GmRvGyfQBgY7FOx3Ic1hI8OBN/sFF+6Gw
gerSQ2G6Ey2zISMRwI5BimwhRooCdhe03U3JoV3piI7Cu+/F4vjs+GliNAjD
yWe4/Ph9TcJAUgZFqvXcHcGErMmp+wetweIYBw76r9k4QpRU6F5Jjo9vT4is
ydyNBWWbp/7XOZwelmQVq+YyB7CDbGoCz85j6N0GxRkSjB/xhCV9TnvNFZLH
jcYm7VtdMFwgesoRblezVL44bZ33GUbznB9ihVd1sOma+vKgayFixMBhSH6R
H9E1ZpDyzhF0W/Wod7B8nntPjEDM8EP6X3ZIqb4GE3i7n8J+Ra2Gr/8EQdd+
gIHhahwF5kUle3m4lEzDmVun0FKL82KTj/milK3OGyWowmP1Ampls12HHfr3
AdokiBGGIFgLir9nijK7jRDhU7TaSyon6xErOI0a1fsHMq5QBVFEEfX+vzjv
fzbSL1DT/5ChMP9Q2hScVd48tKLLc/6KSXHLOUx2kGTEVlEl8CFFlpKUb9vd
z800pr4YzXjUir3uAHv318ueVUwP7ha8W0Qd9EsnMUJASbvxumEx957fog+2
YPGcTlGexsVfGa3LHuq8U6mGee/76pOIjYzc7B+h9XTLfOaiKT8BGzn0XxeM
WyHyOCiPzSgR0N5DVKuafvFKTPk9X8HP8ra+/OHV1Xaou5Z0n7ACWBj1KhN/
MbXBleinVpcdjECeiVFnNXdaTUMCBTC68heTbKNTgQsHWPwrysIYR0+TYptA
v3WSurvVP71ZctkxQDGfoU3Sldmg8ZXe9fXenKp4PV8az43l7jRbwPpoec0E
0/0pmkl0tc9TRElZdU+kRSpvPQ789eFcOcv16W+S1U/JrtMGTx8/i8Ykvp7E
v570TGCpq5a67Cx4tYtnZkuSWW1QtYysloYCS3O/sq4tkH5aTwS3w1t+Q6ZO
e/X17elBoAA67hEd8YfMonyDrRp4Nl5w7/zDxiKarCrDQj8gNFGgdfYRyugq
pBJT3then4d6w030xGoR3sIuGcdHyWV5Z2UBpiD34/vNLN5GB5E2wm7V/Gqa
3iVbdFneuKsGJeQxZVfjb8JLVC6U981e8zAAcCgV7DQPexLInmXVAeZvxZvc
wPHw05Jxu2L56WnEPoWlei+53k3GMW0a6dcic3yLozwfCCewxy1mJmizMkbr
xbMBVZfdci+p5tp4OoSGWEVDO1EZdYWEwUh8q5WYuHt2hZDK7GnLYYos8fwC
BxYQgQFZ1iVYVrgQh82ziOmxrCvsMivsNSBzbHaw2yF6/gzTmsQhWQvArKTN
CFb6mKbJwamMgmZvuabqE6OCzyle7tLILx+VnxmkiYoC4FADtvnd7y665n8v
Z8TsqZlaQYFQirHh0/YO/igBwwlmA52qtJCph7bvRXsJwWLtorWAnokWwZoG
I8hBPi94kO25EWuCeH9ybICeoQkA6/IX6Z1+ODoTsjAzFEmm2xWUvcLrev22
p1Lsx7U1jUu7CEAcOIq1PAdb49R/FNZrIo/Z/ZzFMh7SM2iMARW+XRAKxv5x
ZfOp+2rZiEZ74GjUOkqSdL9dXkepQ+vvKp58KKVKiqrfPNJW4Wd1OL3uk+EU
AR2YN3NnnmVRNQ568eMsX4OMiHlJm0iNDpn6hB+es3gPz8/m1+oQ1AeznS61
5Hu44Rrr42MSfsNXn7yaw2m68/WNcYO3GPXZRNR3xIAa0RYCO5vWFhU5NykP
18kPFVlHE33cK4+AgsfMrCzdMtwGd7ikLQEpKRJBnU5IWJJ9+CsnPaGT2p+a
paVK1NrYDqs2zHOVjqBm6by+0vfJEDlZjmLGY3llER8NBu94+Plj37vIXouz
O8bX94vVJ8F35gPjzM6my416ynqn6QPvHfnOg9qQmk5u/vCK0lVRQ6+SjeT4
vBH6RJh8oTzpM+sTDXZ3cAPmEjGfeKxhKuONvLLudfewgFhvp/oJRI4jnzIC
Ik4BXfAkm80x+H/811KfdN4KDZVbatBoxnwlOGVEP6OVEWmIO/8jmhhbr0go
LV5ZiAnimIoF/4ycaT4kzgNBT6xe4DdHZ31rsFFKCnPnEEonrpyTYu20ukYx
OLbBPy8UTeJ2CkHAWgf8Cy9MdNpaFQuPI0KVfIK/8Ozjq8JpabMivcoYjitO
Wmcw8ERJjm7g3KBMF5Ky+KGmKnPUPCvHhXQcxuHkZh7BtTSaiA37BIlqtbfn
MqhiRteMVB1GI8vjHVdcMkwJ2uGUbTLJTmgCZCp0LAei61XBloygvGrhw3HX
hvyRGvWPBjW87OKGdT7e6J6hf/RQG81B70THYO6PN0UmBFAnDaQHNESa1Ne/
Eo8cR697Guck5yFt6i8Z08KLWN/WkYAfqsTloqGTx3dh2AHx8YK8AlUeb9Oh
sSdTqpksCuDfZN/iRg+LeqNPPU5QGGYit4xe+hpmrmqGafey9JRs+xGUDtTv
REMT7RB5QkzNaGP2Q4qHWOTxyL0Zr9lx5n4TFMyn8s6bBH31diq8UBI1/k4z
OdlEAm0S1p4GAuuIT/iumdoyiBBKnTIliOT7fUiYYcVGqpHZIfrQPR+N0HqS
D0sXclh9Xqhf6C2YUpzG2HK9C8+yF+ACi16+CUvS7bDzafQEywFSDi8IzDQm
7tlFBABtUCS4KGqMITt7PpiuzKwOj28SiLvluDGq24T0blQxDp3g3HVJs/03
ILWbcjA90FBqs+rjIuXeJZ+JH3hcCC+yn7fnCnDmCQzRPoMWZSgqo/zu3tz+
3QNF8KXuCQodsYzCTjlu82MKgD6aleRWzhaE8ekFnvjzFv6Nhy1C2otdacf7
cFhi47OUTW6meOpeeuvnVQKjyutZHHKXlOSM1voEeCvPJrcOlspEyRcZODzt
gKQoTV7WkTzrnmxJWWub2CB90Ol5gsoIABf2dyHbBnJOUsMVBgHt0u9/S4PE
tfcvtBGjb2FEJDZqv/Ir4oUTXKPfCKJgwp//DS1G8DIqWV49x3QO7IWnkB+G
v18HhEuH0BdDd6c5nZbJXc04vy/QwIWYcG+kf5cdFleW4oEeSAcCcWv+U+7E
aSIyQPSGWqGY+novIVMTI1CNlqy0wLd4IdovjcusJ26U4bM/TuFvXuca2XGa
qgQ6rnHZ9gsLohn1MX4fostzW7CN7ZIXZyZM4Cn47qiAe9MkFy+diMYAiu9A
44C/Xg8yIrFeFsB3NfD9QVob2bVJmL6weWQtJM9vBtcEkY+8zGhMd/6ikRHv
hRWPFXbC5P7s0vxJBlclL2jiTvzN6ZM8wIj9rDVglLb86QHpL9VHbOUBsdQo
DUiMKF21oOY0a+Gg5Ni3zlHHEu7giXigleORS6hJ023avvnsrFn++YCnbK7p
jpME1pLxsY+ZWfF1fwlbKJ9vWvw/5EtmDCF0o5d+FBQZhRALnlPkagoc18JI
EPmyxdeA7Xr0Kt3KYcqtw/wSaJYBHWI+MgcNIKH0VUu6nBuVy9lyj5EdtaKr
CtYSOIQiBMDrs3FZXYGP49Ps+UnaciICZy7FHslIo7yHfb+oYWEWdjKAAOIw
QbkTn/+Jzv7wLoqFPqoRd7paZE/zChWOtKoBk2LTaMrzmuBIIgvdbbZszZye
JpB8k2cJdycBPj/L+r/JysmpiE2UubJOhQgio21DWC1dj8AgdFHWwM/sPvBR
obTl/YF/pg/v5PS5b4XJGN6QznQYtcdgcuBvEhWcefKcWIPl/1kd3rx3Jibf
EuyU8Z1kw8NylPlkkvuelRKQj2Qn8hCAbMaZcDo4elNBE+Ha58CmmGK1/GKa
RppLVBtOuVCGn0AUeMrxUPnVx+oaZj2Xfi7lbuc6l/ofvY07peVTR1KTuvl8
mFGrrHugzGfBCY4QZvfor0gaCYeegPOl9O7izVDHeznDZPpAscgg88V+Hc7m
il0NCVMNRCC5gshQi14hn/wburxeBTn7RX2l/Efm/MrYKpCrLdeE/fjK/gCd
hTLxwWVL3WnDPRMvW8ZYlB01RAKQfP1F/qwBD59T2fMA8qxeJy3/pdgHpfO4
VlXrfOvKyK9YPvX5khWt4L0X4ufQD4kNNkh/PkaVc/HkJJwEsazKBV7wZ0Mn
6Fx6kDfy9L4S0rT5SRHOhLzoVT5oW5icv1DKLbZZ32nWXlXMKTkPYL6rQXPk
4+vIuOClsJl+YB9s9Arn8opT1cpSSkQvMvhK5E2hyB14LmlmEFjY65TrEuHJ
0Is7m5YKzcIfQKCofZSqhrDY/mYkr9QqujE1HXFWF63YxEZi4YZwfEixOodn
0T4g8BKyAIR17A8dqMXf5q6QSD6paMPKKOlPMxnWHM6j3q+rqMa0AKtksWCI
pT91NihPPcKp1b51NdPuykGzS8288sggnoAKhqMWt+YBW47bxcsEyCkwnxIQ
cvDECGJzB+2nZyF3J8+UKmvHEFXX7GFTr78pqKyHWzdIQq1i4ZN2a6rI2s+O
Ca+saRdAMYDuwoOl5Yis+JjTheNRdkf3VFLIcEZ/vPT9ehqa9GzP6asmYQ+Y
xCzxm7deJSYnEukERgwwbggyAT4us1xzdqKxe8dpI3b3otw8UiN/rLdupaJJ
fGhYpEu2SqrgvoOVQKXXnDOh8E2qUhnFhh+ao5C0TGdUSQM9uVY9sBYWarJp
ApUz1qwkpL8I/bup1Nt3L5AbiC2bSF7UC0HBoSi4jCR9xR7jznouMzUvGQwg
0cAclFYPGPlOdXlPBLn7tQrLXOwyetNGt7nNDi0UgeYsY5Ie3/z0xd1D06rc
ukkKb2P/WzUdkilHTHechocYrHO7tkMgJpq/Jj0fJMW/J5c9qs+nmv4NLT+t
R/6XJEni+bwaP/QS5p+ATbicTs6c8BPIj/TA+JUaQocH8VHeBu78nn+/5GPB
LTnQ2tGKaPFPrCtr1VuOSFaTZXGowVRRepB2ZdzZW2yaqvOY/LkaBCSePBZ/
4x4Xby+vdQ1ThIKL0A56Q07oP1Ab5+gUgOYjDt3sPgTMtQfgR82fdc1IzHxA
SMaYJAs3/1/km2NUo8b42gzUvFsiAm9O57P9a2ryCD+8uaSSPqj9M7a3z8qU
tZmBpfVbLCShhQuYuegVvFAL2w5XyACVzlzdnCnwsXRp4ufjcObgu19s8/87
RGFZy4QlNhz8qnx7py2Nz4Xd9MCdTHWXvsq/8n4INWmOtv2JakKtvUQJdRCQ
rPUBESRXRSfdy3cUUf2DazFxx056eJG6+CuVxwAhF7ubLv1celKhRU4OrEQq
8V9CXmfPSLa0L90iX47huxu+yjTAQ65oR+wHH3buNt0ik8nk5Ynu3JSGmVGg
I64vX196iv32LAPqX/pzhwLvaA92+afHRV5KWrkNQooIHa3/NkrpfuU4QczQ
tonrtb+plOfoPYy6h92SNlKI5CiL7CkeO/9epr44MRAw3h9JeOWaSuzXpsXe
8pcaLB3vUFheWHTG5/MGt9FC+7HP+FZxW7sEGXeel97vdpGyvrIf5ZuVwQeh
0jkaHrG03v5nOgcipFVlaYhXMrrnQA1pz116ReSdE90tjaEbnxBC/2skGMbU
Fjvbs1MtpFC87aN779pG3d7uLRdUtAuzTaL9P9SA+4eJJ1AC4+2ljpTcmM4t
yLKWWvyVJO902rKZCjtsWJFX89RyhbHpSG7kyIdVDxWyeGtLXAcyjQhNxtuS
jgRAsst0lt5aP+5UNvZOYDX43NDKSrnVZ0P8evBG3UmOeNvjD48xopIPI5Xd
0YQ4kaowXrjbBPgEv+qWw2k6B7XVisnTsQmpyJfbs5iLH3dyBlVQrg1OUkjC
qIr72s4BfXeoqJvHqUrqlgNylOdNnfd3X9G5B8/tL3qT4bmhxPAc3pUhWCAa
V2K6HEJg1OgKgHRzRBD8lJkhJTNnRVi/G4v16swZyme415YutXN1qCDfDUkQ
C2U/QUEZBkja8j9DneQrhdHxVaA9vAmfrE9CWsAyADGlvLODHgM5kxX93A2j
8WEo/X6PUho2BJ0ck7EnZBct51D0XyVLfDdyXA31PKqZMESQC6r8JF5IN/FK
0z4KAUrEPX9MZqnJhUYwV9lIwKd4IEqXt/LHHPkhj6GKzIzg0BfgUTxhmOxH
mOu0iiMSfAhI/km2/v2UpHkw1d8g09xkzXG+IzAGN8RbzxO9CDqV37Z786gX
h/brKzKQUZEBlmPAzWnP3nipU2o3OR/2GXa9sivTo1iAg/DeNkzZTnMIJaym
I3hEF9kcXsNXKya8aKiwBba0cUFKhYZq1VqCSRAysta9brfWPWxvpN3Ky2aA
rc28u6VFUpV3u56uBzHCN2oi7r0nr8sCWMkJqsQkK7QXteIvF/MJyDjpq367
JRTRjIWnRSweq9Y1XzmPcTfoDdRvlTdB3rGkeB6kvtP6x0YceDnOzwM/yFQv
9HxlOO+GDkmD/tlyVLs4gIU/iXyDzuZr7Fa8fNo9dbjrIuy/wyroJfNiH8/S
Yrm5bbzz7U+zTQX2/LrlAkrfz3LT3el3CIh/07BWPe0BWa+cBqxNeMRRdmkp
J7TPx0ps+ERqbEcm+n5hFJegbN01fZ0IocFyGkvP7HLK1g7uQW5c42m7pSYx
FRk5bLJ3Y8rZX7hHd8kZFBcq+c9TgN0GVl7qvKoNlZhPO2weSLxGKcZcT9q1
QDiyXH7I9Ps//90YjYul35MZEcDOVdHA/0GwsCSuxc5tigwi9A7vwv39CYtG
LGLk3MXXjG5IRiNmtGY4wzkU4+nk5ULelM+tH3ZBqsHjK7Rfu8SQJlfWNCHX
5h/L9yWRqf8toxRKjiI4uzpMMuy/8RMPM7JPeVaty3B6q5EA2ko55s385KGM
lmCTPynwdAWmObbocVo1U4Ti4+f7rpj3zOj5ngYGfLE9FMZ2f6VXGfKFaMfe
EGI+JyE+Hv1jOoUh42gzUMjVr88PSNqs2kz+9b0Qg7jK+20oJEeH1O1T43ID
1Iq3WOLZmYne6kYsI//OGcHol5QuW1HtWMOSIxjOh7lZcKzBzQrQC+YD3hlA
P6T3WeYqHXQpF0j00renY3Wnn0CTD8uYuBrf/mJB7Q8uv/CWX5AHZE4c3vC3
DOkRv09qBy+45PLx9Lt1KIWiWH3kWVlPowyNwR1zKOevZTCOTextdii73I0A
DgraLTrVdJXiW/HLzjFpr+kZMXUzVmTplrEN9GPIdX7qk7A3yNpMP74iBO6/
xfbck2fhIL/CtwBmLth7GshTcV5Jp3jXAU7cKvobx+ukTfEAtJI1KTWrb3FZ
XOHHZ6WNXFmKAPTl9oP8PbjbKekH9YX1+/6kXTxaf0c9+aV6F1oxLwSTBQdZ
Ww2eNbnFOtqxGqgaxNBVrgm5q0vVFQrmVhYXIPZ/46QT+UZGmArd1k+Oix7J
xPI1s/9eTIBJW75CyHwY+0QpX7PnS1dDCQbDQFhFItjLPZ3lyjQu0uVqslKk
B52j3fGoa/vVWfvJre1JqoEVPwGIUe4NnUSdO0RblEQK2zUJFMCBPYtpGGba
cYd3P6oHIfRcbH6eTfdl9NbV5UQ4ns1FxD0QiN97h+kbqWo9Nd8JYWtbUaBQ
W25xJ94KgHSMRVHCYFd3qhh3VEnVhHBNv8IHyUgRIXQdfZTchUNwFjQK3Gjj
O5jXvcEHPbKid1/VqwSdmDNs5scuN/98JnRHk4VgZ+uo0mm3TvIijypZV62e
yQLIVTiLsQaQ44+IuppC0kr7+Y4ifOzbJuC2TI9U6VOg60eEp8XO8Vtg3FRc
6H2J0PdUvkH6REZztZgfdKjG+6+ITRUtjYnENnyLkmqv/wBLT6UaTs/5J2wQ
uValiALFt6qwRWTSYZQgmLYGmyUTDpfWURcnyRWxY1KKph1OnziKEgNra4Ok
ljREDcewqZPQ/SdvQISA86tE6xil7Va6ORtB1WmGwTN2o1kspAm/NQiVMLob
sg5ZTQHzWxxTmiaE/M/kGlAafBkFpYxOvSGNdvGqBSlyFP+bZmpvl73TMsxk
D4ec9rrYkAOH+rlWidAbaqn92KIFx60ipjuCuv5ME+V7r4CkJ1eZDTDySaVi
m5bI+OasAaiI2Xdy3FXtGC4Ts3F9/uSYA/WqXZ/VB/UlHvnWpT3ocHrkjBTq
TVqxAvo9FoLbYsyEDCgAPvrXFXUNc4TNg2p/BhkXQCaao8ev1luIety7WFrg
oFem4YGBYiQFOdr8Do/1kwFHDgkwOMcM8OHagsxi0/7bpH7MtptqrllzKF0w
vMkzPCFuVsNlF4ggJbjh/UWH9Fr8FD1xGPHeeRLYvGJsnSAoaf4tSNKixjCM
pi62dzDHrlC7zU0f7GgNVp2dnG73TeMX5miGklfH0lD/58k+ta/A9+HefpAl
VpZa2eVbOUfE7Sdm4nJUx9A34L2IUUC3yf1vbhhffKEOmQoYM3tcoljMlL+g
qIuSPzaHP/fV8b7eAC0iygDL8enEmB7dNLWNHA0MUTkUsSNacLHn9e7b91tc
iO+ExuTP5w1UiOfVw3HdvCUUymvl3PoXue4hIBRuIb1CtlNrUQH9nCwRWEkJ
Zbf9h96W75uY6Xj06dOqTPVcWWoepfbAXX6IJw4MwnSCgd/3su4AS9GNy4wj
oFr0miX74oFpVx5H9Y3YnvpDK0fcPX5uUDbbCAKF1mxMBl2zrtVpJlmASGFL
e2X4qpoNd7U+Po0oZIMzZxjswcXXrGRQ1u4prlx0La6Q+pSfsC8VP3Hnm6Gy
7SmpTFP4nf4zFfRi4XhiZispOpuz1S/92rZ3WmROzg6/cFjh6A30Tmd95XKg
5fIvKTrsUO0TrCcNiEX/EAX9IecHohDIovvD0hun/iMBxG26PGJyRflpaqvU
/za4uJN7I7QStx5a0jkleDvQ7NXqjqeRD/yOiBuhJFlDkw+Z1BkFIVj+WDwE
cQjaSbIHWkZ7WZQjbxG1fB2uC1UDPR3B+jBXL0+ZAaDaojsfswVF6h1JqJwp
nsg+ENnY2GTXG15fPo2YLM/op4SMXgfhRZTG+UwPU09OxfLpch+A5HXpGOQG
mHC6ijTfLVxzylhDhcIetRgi1TEKddKWsPMm0QYbPfVNpZx5X3c/bQGSJpDA
fLP1bLaLGPQC9Jhp8AWGtRecVGTmZQ76iditDzg4QzRSzZSfIURpREnisgI3
2wxaA1wQXV7rSilpNjxiausplh0RjlthWfZcIPtD6f9oYlO75M1VfjaztW0R
sj1SJTUucxRGt7xEmxf97/CRgsF7yXQ4xQvy7WvFx2LMCfCIoppUdhyNaHdd
xBJ5sdvOqOTZb0+Rdkzz1s6dDGrtdXGWIfI25YWqEwVZ/rUItTQtCWG4PdMr
bGe6NWySytxHyqURHbUo6n48Mm3z/K6tTHsuTXH25IF7VWCwZCzDAxWVyBEi
pUaaXVQk9HKdAmHGLFotVqabEeZ8FeNKALnt1NhDRwsvSyMVYScaVH8T0Q13
rXj4KMpM1Zwf2dNLDsPOJTXqO+Nnf8vrkyWx3Ujv+Ogs55KRORHPPptbiK57
Axu5jNhcbQBdJDN2YdO/bXiZNvmO9Hj0ErvfBoAinB08l2gI+CoGkRrkIqA8
AoFliNE6SbwokDDaG0oVjiwjPdxMpmQi0/mUdqEu1NHqYYwf31rS2Wm3epiI
qxueskgYlmColRfkLrYky8Esm6MKk3h/KXZlfqHMXD+2k4nCvqXHgk7Z/TlU
eAP2il3ZxDF8H5PR4kQKAt9LTkkSMXKnYlxQA0DU8xYBwtYklb25kvquO89k
EEvPRy8z+2SEhmptHb47WAccgCDMmR+iuiOqkHZIom7cF4YYcnGX7maoH+EF
Pv4p3QIAhNL8St1sOLblFCbOVVx9JQIQUNwvfxLS5PAM4TyI0MhMh2onxXm1
rRCr/q7sKpozpo7FJkyu1i20DDDuXFsIyxn5QDGjdXChzuMN479KUChsqi8M
pfcSWUN6URrXQFRFJcZgqcAKEJonVUv8bZjRv7MXFQn+QIoJoZWVpZz2L2p0
SzrTbIYB5svdqcWqc8FC2xqwrGVnEDOyR6QB/wrl6q8uHf2x8yt1V6+HVQAk
8rsALvzeOf7HYj8Bo8gXfZprDkXpP2J6vFIidVJZKywY01cc6EWkyfnu2NsD
Y+z9OSCsVODoae0V2gx94U26Xd/SpEWw2XWR4UHmgteS1EN5rkXbM7ZOZdMn
GxdjzUmunEnWHlV1xqofzx51x/a/+GFjNRG8aXDu4yXPDW37lHiErnylf2kz
ey23HKKOpQA2G/xKiQ2kHEd2vRZY2g0MfR4o9IkGvRohd3XdhKMa0g0+dv3V
FA6nTU/Vq0uQEdovgsi0ZfMrPbNrZoIubCVMtXFSfmHyRz61dM9hZf+6EclA
+6wlNdOUYP38QlpQE2ruYMBeEQ9+bbaGSai9N7L8IXGncMcSAfaAkTRknREG
wB1t9DNyDSso9HDsmX0Fd4wctixcpbWoDiCG2GRRphuq6syDxaOnqxbZ6p5u
7aVz7wGg06IyDbEJK8Ss5FnwZhbnlEoW/IBfu2ylsq6iD9Nx4JKryd/7CJxL
+iOgL7Oh64oOBO7rP23FEgSxI9Wxgjlv4IjYA7b1R5cSzwFhEkKpi/hHQ7aQ
lDBGvyCb3oaqN9mcEuNaJDZqi5gxP1GPbrF0QQslacp5hKmmogM7VoMqA3Uh
2eMLWrkz+NHvnLJRMlnCe3/DbWClPyKQFZE0E8VXyYMq9/IXhyL4/mqUEdwz
WXgi8H07TY1ctATsOPhSTswhfVDoreIAMoSJZk7oxdqrdsddwHqRgo4zNmLD
IY3Sg8BJhOozjTp/omRZNBosgLsNuS1aUxGrNdp2wUI1ad8cohOxbxCD1Zhk
sErKYCCTNdpzyTqCfXyWBJYVTZ5Ro0e8Qv0NvVN4tPQsltySDzzgqTvXn2V6
hdORwqO8NY/1ZoyJbHCNhv+CXkW1jn+h1STIeyq3uoEDqnFvc/grgZa9k0Zu
Shr9wtlmyebn9JLDv95M0az2wETcgE3ActyvKfYxjxg681VCWMjzAzlEpW2p
jXmQ0LAhYpC5OjgWqYAeiM1MaGSvbZecxkXLVrouDGVnZRfwq+LaTKKn/WHe
MujVtRjHjIxyYSMAZHH6Se+0XZVwSXQeTK2kwX5Y7PnvfaQH1G6V3IrXZa7v
IPBzOhgEKJ42nRDYQ8g9b+T/YFRsVuMJfmG1C7I9EL0TytLyMLCavMTuUAGu
K4aB0FBc14FtZ2j3LwfNouDW5tNFmFk6smBXJknuGG4NPTSjTLqm+mDktKFL
vBzXMQP5I7NjrvJvXbJqLmtSNfpAcyTNitDo2EnjiZ1kRcqeAhRGC2DpTmcI
5tAS+TxT0fF4GeozzGCLPHV034rDBnFndFM3Qe1iPHBVXfP8NZo1fI6qhjsl
+feg3zIMlxhHq6A9q3Y798PqCW25LE03mWsF7/2javKjmI+VpNs31SiGCAks
aJefuH9ePEb/o9YmIGBRYnBmLep77Yyejwr3g69uQrKBkISrfe56NWjtkHXi
If1Tr0o6b+263cJrtODtf7KTeYXh6bopg2jot+D8Tj0GZKLmrfi+Shjs0Ecx
1wA8/Yb9hX+szWry8w9kszyAgnyhTipI2Qpg+qjaVth5tLQ1UL6/NU2CkILc
bh1bsm+hx1q4TPNMDkIGybChBkw33epG+q7SmhEmgLLP2Lkhe6+Ci4RuaCmv
K+In4rdlZCWN7gDjhPVVrdZPZjgT/zABr67IxYDOm+9Lex2mlHWotTweXYYI
KcNMWrAItsYn7iL3hd53oYW11GlorIcS1E8nAMYfirjGhBRoEY93A96twhEq
ebZWzrNbaEcOyMauvaOXHKsA9C79n7Lxyu4osvmHl9kzWTbnJRU9MOe1DPBC
s7V1Wvf1kz7EplqekGu+V4svsTAD7qpU14+53HJwo+s6Spek7QjR8yhtKQ/I
YrJbkAkGeFeLTGYUsS8ebfLZMYiDDWVn8zIaIjZlI1NONa6zpbuCoH4M4Opg
grLnTDulXp2+MOgKi3FoojMi3m1TFjdbDiYhIdROllFkSMfuXvU6OJax/EIj
NwSPOFJ3WQjvrpwhCeu54zTfJZygl86N2mfIpLrOJ1npb0ddfc7SBm6opUND
nmzJ8P1Gn3yyLzRbsd6lWSLe8s5IFirIozjrEbaQUO70jDV7+X7DwS+3V8iF
KpZ7EpPiFZrdWsb/+sv6BkY+7mAvAIQZkpjwYD7DdlpDCfPSvw+pH2JiJn6J
+jGIdhxGtz4si6iueEsJnOsPWM6eU4DCSiz93NTiyL7sFYf82TEDxAwTZUeh
11hFShpkYBCAuVcDbYc4F7lN6ZOeOXaTrcj3gbQbG4pOETMcrOilxBk3lOMA
Pkehgg7BE/P/tQ3X2UgvtRdRVZJo5FXwMXKcD/e9JVaGf+pdCtiEr9l0aBfp
Y1ESWJ+x4Fn0zd5J2JbkghP7OOrYcGZoh6nFeSdFyu/gjBOCysmRBSZIKeHC
92D3nacnwBpmQTSMhlIMHi8d8wRLcuIryrouk3WLI107YlZri4MWEhcqcp0M
867W8NwVQrwCZELMnySYBSM2VOi7yk4hKEUh6Q53YjGpVEMgpxo+FDJiZ9ix
P3C7ZO8S3gRKyQrJZCG4MnvcjN9YtnNC35a6fLb+vRnWMhn+8COBRSzYw0sm
LUsz7hkAzULee+kNQqEwPlH2EOpG6AQrmzaaQiFD0sMgQCDv5KudlxCZyZiG
e27WWaATIVfTDeHLW5CrG9YetYgKI6CYCwZ0/YTUerXQsdJatz6efDPucfR5
SDf1BPfl7VzLh8SCIVME+pa0cF49eqrYOqqY+gZv+ovG1Nyo60d2sKtjz8L/
ewSby9EgBfUi/rxsREQVxbnMXc3yJU6zJUM0p2me9a/DmT0W9ygTi3syYdTm
3cTP3CEFfVcEOMpSwvp5/Z0EXXMiV3juqLLzPNASNVLz3ytWKMi+groxIBwJ
GWbfwomIXqhAZG4h5wGkrxzsN9wdt6c3wEkBr+0KUR66I53DJgOIR3JKYYVg
NYxUKDn/D2unjrq7uXiAOgpXW6q/xkTQpTI6f+K6sq7I/jviC4+KXc9B6qX0
isqHK/Dp5wmfCk+3rRkVOyaT4aC9YdLld0xoKpBD0pzz0mEZdBfkVDyNghnk
4i1IcN/4nsVEe72wGQguiEsNvdRtolpplKu1VAq06bqV6oJeLxyhwWTER3Fe
5q+GHlwXkzqfL0Ixwy3v8QqbM7+2a9Z9zwP3qeK4NNAGnpX0+ZBp4Bl3xfMX
2bEdi15bQySH59rcyN/QZHYPlobKB543kxpd/6mFK5aVZGHXcwbmRpnLHJ8g
E2Ale2QGNcc9zWtfKPDo0/xpP3GAefb0AGqBel4P9sgvQc3KeK+ealsqqV1U
02wKdlOqysA+efyLrdoLy4u7LPZqxwkB55DkySKOpSqc08r/OqzSVNx4NrBc
RCip9IUcy01Fg+VVTdCsJoiA7zUj03cM0hvjvbo9PH7TFAJGkcB2P3Qc1ldN
ABlRjqIVSKHxLK1G5qYxjCOjUs8ze+OfHWBMt6zJUm9zwOsrhqYys97AnteS
gd5HOhem/iyMwqhmWktXAdOhRxR7qqntksOsCp4fipYRrYvrJZv8crCG1V5Q
XynGUYPyeWqeHOR6wvKbgpSoyKi7PEgvMSTTzewAxwPXbclWV2zahVyzFVZu
P6GBz6ZbLZ/yFu0fK+vwZFE4FB/O7x4cQKoaucInzi5nkuouZJ2x5f19r/dz
u6c9TmvNSpwvWYweYHvGHJkKudmrGu9aq6BdSR2P1I76nYRPlGSm3pB7ywSe
/VSLhE9LyucCip3V5p8WNdUjqIIpWw+grtFJU4ExZYTJy13V30wSeHkW+0sR
+0qmWXVLCMfVHAf9MYZCWZb9uluBuxuplrqZCXjb/HKbi2D7MTjLmCPkUB+t
PdrzrklQSqKOtkprpQj2cCMxms5y9XIBtlsogO6ua5uY1rX5mPjBqNcGiKXj
/Fm21zdC+ZvX5qwIbOC7GRjyO8sNuUyISzHLlh0GF6y91924q3sIR63K2RSY
OCtQn7eY12S6rDSA+ZzsH307Sczsn+Yoycptt4cwlXb9jZfOBgIRHsvW+aYL
STSObAs4o63lC/AMkCwmcTucTjRfZC6SEQqdpl1TJ04VlgUyWkD/VFejjLEs
8BHATlLzU0C0zIw4QHkH/vfwfmjjPTujQjWFFJs2sSg/InhRTlDD3c6mDd9V
vlnBH20b4AZzjAD8O+P5apY2Ix1NKOrbmXR8iiJzaV2Gwfth9xf0sAO4M7Q/
xLbFmiULdN0tfi7PqTmjZPREOXbLR68NhbTWEqXGN6liasxMIjXHaoaIMoha
oL4YMOMcpXAW9RWVRO83AR66VffJ4kBpejtyDc1QgrsL6Rr3C/vBBX0Ocf00
pkTjRb9+f5OZGqhdjU/THeoSnlzx7l9n5E9h0I7lnzBzpqvOaqAJy4zt+Fli
TZ2L2vSsUmYlcbYpNAVAoqohWhIr6MBaKz1sdOwRfnwcQuLnQnVNc4xKnb9a
uPR5lkMl/9dFHyXI4/zKMoK8ZJB4CJnjdXsIlDTS74F/qptnM3rWT5+WzSlC
BrdFSud/bT2JN8yNXHTfYJqkyoVOX3HcSvtFEUla6moM+iQpGvQxKsCQ5yhI
fBdejt3lzkgl+wnAII1UcnKC4fpr6v4Ca1yR3hs/JmAvgCqsuX47vQwtf5si
Amb+oJa14XZvoKgtN+/K0GI95ZjcDc4s9/8eAT6mLwXuxuJK0PU4/zac0kCE
HgjffztiMGyXBR3/B4/Fwh/HIE7XZa5rlDBzv1utPuLaKWSJg1kT5CpwovjI
0c6PwtaHYdrEcWOXvgs8DLid7Z21374q/aIAVTdXdTooe1BXmC+IzicDmhp9
Fj7Q3T6f6aqRmmgP1JT3g3/QjWq36amA8cJe4Sbk8G0lrRrkt6jWPa02K6CM
SaAdIs8g7D1DIIEFuvsd4d9djTMInRWCOGGrFVtmyeo9hI7N2EHyHqb8w56k
ffXpN2R9xhp36x99lmUQkkYKnVutxWIxhm00S3cSvWmMAA8jSEmrpwKOcUub
1nP2NAEPgpfraVQ8N853pFVqUI0vO7AI3wxYkpLmq03CXxTb2/jETuj3iRG+
xcosrqqhfEysXfAUJsKsHKFUE/5Sirlapz/rD2j3KJxRHLyLu7wBm8QHExgm
hAkNcv3QVJnPd7JMk0v8q9m9iOwn3NzJza0WgdA9GSwXEXxpW3e5eIIoWEu0
ZLFwGaH7SLE2nxEqooMFXcI7S/sFWLSAsUKOFI7K4uvoGjKV7N3K6tImm4sR
9VsiOguys8WOKKsEVsQmeELnMrPeniFqRZ0lI/ASjhAbDNSW/0DDc5815aA3
WFtEym0eSXWvhaD/H7Q04/J1OwvbAEy3/3yhKB8VEQPE/c/R4qlFjsBjsCT8
PzFwOBDv0W9TKJt6gIYf8D4olkYfurTjwqWUMt9hjMD3x/CANscCi8itfYW6
Az/IFHbbnZmIXl2+V0TD3E9A+0xo1XlzpeZFnr+//HnwR4e6RTJAFtkXYSSY
cp6ct1IlTySq7d3F+bsvLKHTuXSHEZRZl77nz3A39+TDonUVVyrBGba0PNDC
LJcnIbYfEk3b6jIv4TTjhTc8M7I/qKAjrgkg0e4OatmS7l2aWWyu/ANWIDTP
SguW6eSo1Faof62sXDgiVqK9RkrPOz5TRX+7VKTH8kjunuV5qMuHcjO0vBmy
J3/JLywbxYhHFVTgOO5XcHd3g/s/DnyGS+wbXlhl9M4sqsaLFS7MwpK1FtIv
mnUfSRxgs6YS8aJqThIUE1Xna0S6UkI3lE+6IhKrbwjbf7sC6HPwY0eRCNhn
GVyWaJozmNOmh5fIR05hXYQpKLCjZrAk5LakJdat3v3SmyWjCr/v0eyR8K8n
fYuxa3aM8InWDJgkELK9dutUhY+cC04etoJCBiQPslBO1JmnhLnemL4kyEfw
HK4447c8zyysa5fgNjYH8TyucMe+pT5sdTxa+b0iATgKTRhVXgKGpFqAVAUn
wS3aZpsBer6ougTJz83e3FOVXLnBxkSuv/JROcrDELX+QFMuDej75+rq+gru
ORJnn8pjPLU8vByawBUowutbQwNVzykgj0zZqAN1P8ul38uDzFjk5wly0Wun
rKospxyc+IiGV4Gep4Mw1Qm2NUDHy57KAEDTtuEV+B8ipQTda53FepttxTyN
SNWkZgsXB2qXAdAwmybJuav7u+08gfBeS7g7BIm2yXwKyEWWYiG4xcE5w+Rv
E4iwFydb+OU2fwIdrFaJF/Z17Ox1pOxPIW7mNPp6Eodp4SNPXKBRxxFqHTCA
XqI1Ss11+6xunnkNvk4JZfeNRF1O9vgMgyl3TBKOXPDO/BSNfGy8N1U9ytIV
B41xLR31tpM3kpYHUlMkX9yoEwgK8JFfP/XvyJ+WpRYp+t0wgv2ybELBYhM8
/i+tAZgigPZASEiR+WvFMR0g0QLprelSIH47V0gXHv3+P3LTMMuW8Mbcctat
N0Dtnxax+OL+sPvPA/Gd6goutsQSBb/w8K6IxQ7U2rdyEfUCeJXZZgx8mFAq
xTtBjpqvLz0n3FEv1XozaHKk4K+GNyfPOuB4bPVg+MUPoOLvK9a7vsITIAE/
wwlv8+/85Tjojfsm1YdmfQevCwnE7bDQKWgZ6/O2HW3dmKGWk8C5gTAGd8sI
FwLwsaz6trMIrT9DJZc2tYYIgtzFX9soHNBMcEqHX8k2YYGYq+ECbQC0JRSL
talielv8xK9DMXFA8JuJxOQL/xKixS9HcCgqK0D+JjmBNHjtsdtNRFiGMu+L
iWFHbcRz860BegV0ikztDbCgwTqI+zNH34Dz3jgQ2FGJhRS/AROvf8crKn4J
e9RzlZKOKlxE1gcg6+RIYrWeYyBHgBZ4POwh1uv9Frb4wiFwRGM7VL/qUE0x
95WFUnDLus6SJybh25Ppyi67WYeVMCfErjPPbXdT01vp7dBXutKfRnKqRF4h
tW+dx/yn7zjz82N3JPPi6AnjUlxgnORbn5zUAoQMbXiJ5VXtJDfqbsb6pyfY
xNz7939DUx3FnB9QFoh1ObL17jdLoQfw191Daf20wlCRpBggFync4mksv/vw
pX7aIKU2Mi/0JnKjzslb101xNhLs4r0NLLu3Q6KyPU1mmv7il2RgwIy1XIVq
AqF3UOXODLzKwqsjegcMs/eoVNJ3QG7fL1YaEbpSzXxgBmm9JVxHqFTTOimt
TrC9P2CKUI/8ld1eAqrLqn8915HI37a4CECAB96SEondJjyooVYim9dAX0VD
6jkLORoRdKd4S1nvHDtGWUzzK581Y6poAYyRczKSHbcl5Qw4MQw+fz6TolEy
O9cXqhjWuRqGZGcWuFxxxRXBxJIOlv1Z5/5h4OmPWAseHoKW5d2qDrT63zfX
pbVhrQukHhTeP+wpnHbJGXUxaXxOZsTLgI/ybsLK6KoUPNu50RAkLKpGDAHP
qOqYbjHZVmma7HQuP3Y8N7nFXv2J8QRm6uj40YUmJkqrdukDbyt8MWigEIRb
VKrLjj6+Gx+p/40m02P05dybkECbe+nVtPj+tPjWFVAgYGRg7LzyUV+v8h5P
tgZDZqI2LeLHWTbC/BX5+hV4yz3R7Dw74zjifqtw2ItBDiqI9uFPGpgqtksT
FEqOAogJYD3FyLDXjzQz1AqF+PKDxUMbrLxtxH/sRBLPJsQvUrxaTGAtLr7o
XZoZjsdV7dOm0pJgkyRYExS/qmaMmlcWnVjHnOYGTqGJdn+TA8XIsWCmN6dB
rw+Hs2P7AmhBQ2Np7HR7GEgmSctgQLTH0sXJovcMj71gU6Ym2SiovsovrjTn
cpBvHk8svNHmQvJZ3hJDhS/81cN/chjgj4XCeNpT74wDXMSmeDxvkrB0Z7j8
WER/NqfvaCcP8mwGRObcGiXJdtuz+gleAa+eTPkvKzag9AdjzXvN8hLdjGjP
cTlJueBtGUgvRvF4x/ClY4Gr6Kde3KDf693XD46t2skO7x6hYp4X3jiWb8lL
x6X48PSxHLb54xew/n4FCu4KyIXKjdUhUqQ+lKUZpNIN6U6C/+0ElZQebz+D
WEAd/bKDLQ+euOOXbSqb4E89Rk93kmLvIABnrmL6RgxWcAF+DAzU+fSA/GKO
RWfTfiWrzW3wcLxPZHlfCi2Verc1EweSrehdgMM+B8dXjsXxnKd4OiRcjBJr
c4vad4XVQGx5PVrn4qCmqlKttRiAEPsvKlnVy1rGzKmuRw3gvMocgBeIho6Z
y2KSC4Ed51/tzHEWNV1fArzCjjT13nO12K9jEjtXMq+W2xkkB0IHfgB8W5Z8
PjhVSQ1QgqBx4ro5e/ElK1xxNoxh1JoUmZEWtwJ66x8QHeDNV4fUT/+1Olm6
00ZazFt3Stowr1xt7GhcRbHqft909O70rk71lDJEA4ZEvbhJBRGpLSVZouwz
x4x/LtAKFeP9GYdXsJb9W+B+BV7nLhVlhpWARYjNr51ltGFmutRDgm7xO2Yz
NyR6l1/LPztm3xcHNB4pp6maD4aqNKdv6rtTG9IAZ6nON72nFM1RpoADzBhP
kStwHhQHqtJ/fm9xbVP17II+BxKuDdjD4mKXEHwtcUKEbrfIyce2K2EsL/Y/
dtg7m5B9bkGoA+xMgXRSlJyQ8JRVrw8hDNtg2i5qQlAz0gFMvViqWk/NlIOq
bo+heL3o87zsTuOqqt/bx34+fQrysD9p5Af95rCguaULDXYNgyvBdLIBlvlr
ORo9RL3h9yR0B4Ode6pSsr4mKG0lYwOU00PXcuN2wuOTS03m15r0B2dsNJqV
Tvbf0EVJvFM1yWCU+sL+jpPIrZo4gMoIuK9aitTDBSEJfx/kOC3aaThdkBl4
ZZYUjJIdlTAZRo9glkMAUYDdR0B+aT34WV2xXUN5njJWoB4JFfaitD63csBe
Hm2h7XfrY5mMANS8B1Nm0QhqvFukN2BMayhttd9hgHJN80TeQE/QQME0ke0R
ZF2+La2irilXyNLkNk4UBewmdKUjACMAY2E1wVo6t6CnEl6+fy1K8oVgT5Gd
VSxYwKybZPgDc5lzlCU2zUJ1FaUK8HcyM2CvbQgqZC9eo9kAkhQZ6RxT3/ez
oGE5GZb3Zb0nRSTpr/wJy71udS4Q8hxwQTpK+88tdwAOzUGMkUNBkqjhHi5J
Ks1uhNMsOuYrShUa+9i8llBTO09TnboAYwasdiKCLOvVEdBW+xPLnhPoHbO6
WAKkajkNtj1OqWXJ+yMInJ1PNGvbvkDedeWl3LG05x5IV4Madsl/H3oitjvE
Ur1qZ2+zvmmPaBdq0OQkc8AQ6Eq+Avf9HfxCutwAhrrsjLxKwuwsBiV7mmQu
yTBz54e7cV+BmVb3572Xm+wYPFY3UhJsjMNmSPLwBec90BW0P+tDSIl3zszC
+3ZkmDVXCnoDInvzV3fLi58BqTzwTelEwLKYDWQXDuqp0UYQkpq/zr6hlkE4
xZ+tIlL3xOFXziO/W6nYvOJjEw6524fgywJeMNjUmNL2bn0fyshJipmezGOH
oF8qs+e+/GGphsYiduuwIKI9HEdy9AT3uJCvlJ9KMSKJAOd44jv27q+iHZsf
P3x1UA4y6tjGuWlzI3cmPjBg87uItgPl41HqrpwpSITdSYIjxQGSzvxxUc5s
NR1SN433yqPRe/RSU3lXyuMlgsSrVzSjgs1grUoGbbORebNX4wwFT8TCaOFr
FAmXEwj6G203SFXUHNG/Nrr2UQKf8tqFgCmEQg6H6tQaAMZRB3a98Z3dCHL+
U/Ni93xW4uFmk9I6LfJ+sE7jAPv7aLLFARBOzUlmMajgy6F07J6Lv7h30dJF
XYOyBMBkSh6gTzr1bd57D2VB37orZslGyY9mZQVFLSTO+eOBNyvS3hKwBHxZ
wdmvZUTteGVZzngKxXucZzivj+g9VgKrXNp15FwU0aoqlkRDG8phnZXN5DDC
uUbsWO/4dtvQkXn0TvqT4ifwLNWmtFCv0anAN5nBfLlvAAwU5ZvH2xWXj/9m
rKpOhr2l9/saGtpAJ085DZdLxJXT2DOVpNUZvGduv7Vt6WiyMkcr4g6ckEh5
eLkTmWDRjIl9OCNoq82w9qIWuGMZTI7ZBAaiaAP6lq41wBbtbQT+gFq99Cgw
y2H7nc5gKR23k7x7KxVt8g+1vRjs01+CLQ8sWDXXhBVHIAsrjl5KzQ7lmWqq
54ONbfcP5M1rZd0ZNaa35IT1dA7ejhHC7/9iX6ZmrtbQQmm+58c4YkUnDsil
lL85uelruILzYrSMgZsolxaUhsw5EUIihpMPzcO5qxqHzS73RCVBvDlXCMPS
jgkC07R/mmgRgXTjNqClirER1Abo0innxLoMwf5Gq/Rka5ilJiQhJI5Hydj7
ecXnE3OiTh9okFXT0zXzY3Jn8QQEwrjM5W9ofU+aA8Re2FpBsTGsfe60pkLp
lOKfQHeYJd8XGZ6qHXD5jGrI6nzj4zrWPNK90traMJVp8jviQEKclJbyd+me
hLYsAdbUfUYbqoy7tOsRzrHYy0XaFgpfQqZUTZTvkKTByVPl4SFObbLMzXS8
hMk/Gpw4ggxRU/UD49Unnh6V5DDxspPKMqIrpc7kkZ62PauCRDh6FFa9iQPl
/5shvvCoYI9ipXpl9HcF8rM1xF/9jQ5N5K4dSjlH+TbmxY8lC+s0/QXU4Vjl
V3Ss10Sqg+y/MStv5Q2lax27PjCQQ/Ys/DirFN1JCv+ZZLxsr+KXidNZovLr
xG1OL1/m5ilJlK7E1VZ3agd7MG59GAukHZhIdHuyH26DUlj9Gv1bWdgPkZBo
txEBHr+gIHBpkORuWlRXYu22IixA/6A+WZm9P4rb5ALZCtK7gYtKg/PRgqD5
n3JGVY7ExgLI0fuFYv6s6vrYKX3VE+lX5aU/kH3t3XxzjSUOcc8a5uDqa3l+
fVLLZmjJC8mnYAwaYcmzXeozIvtvoSFFWGYf8TIrKMPZZP+HEd/zrdU+j9RJ
g+FDiyRn17qWdD5b7cicVuG+bn1rv7pJsmbZTuZ7JcB7IqM5cQwgEJeWPIVm
dUV+YZQFNlO1rKETsrqAuiAp0YvLAfB8D5B0gI1Wa66/4SYD30ALX1pQVEV2
pACWdevhqOFXhtTd1exOBq860Oro/MF/9WCJAIAjd8dBG23F3UMMzuexB8lI
/rCnJJgbZKuDNHvthh9PdHLr+weclhVQX3w74AahKybYVTW72wU5AMphq2ay
HpiT9gWX1nt9yaAhG3RdQqgLLU+8fvM7jK4rVeaBxMijl6DlDAjFvc4G16fQ
IIJsMuA0nOzW1fhU0Pn7Vmg/dx3ZNV2i0eM07KiP3xb/jvUiPH8TgINVu5WQ
lxTjs+0KW8kpK/cNrbj3EqW279IRtkF/srM0IyuxFhH4vtsICzI5/AURr+13
CDptcYJdQzsvWJOjC9eoLQVKw0kCHStBbUigd87aHwvJ2MEV0YGROhYLQskW
7/QPcNKyanvSwknouMeEc1QDzB5bvwswBcYOodXX7asDaqJGXGw/LvMEHgZv
NNEYS/iKlo2wv9NUa9F4FZeZhZHCI1YyBsjs9lAmBD8amiDPqNnIQFNXEmX+
B9uuKmg2UYgL3YnsJjcoMS+gmzMabDP/p8fZ0pbJkrFxfba6zpgYVwrcxS3E
mQxnKl4EAP8Uif9hwB1dwlZO0Evjggg8PfNrthRvMWOXek3LEInvIMKW2ABR
FJZFxhHC/9gN5ZhwGaF7I9Ccc+tnUnbKr6epVxvv9WI1pDq2+Ir3xRZbfQfB
Nk/Czm8EPv40tuWi0e8WApl4FMnLaIwgky6t745VkBH9397w+3a1A+U/RSkx
SQfDq6nrSqi3GOAvysjofq6VTxQ4jhR3Bl1aksRuqIOJ4j4RzdJqWIO5zDDi
5EIzqc1T5GVe0TskSFoQSWJVs5JURCuGImd/fxM3lqsp5LrtYWoBXI0PVhmZ
4mUUWdv5dPDSW8aaCUfZzw/QnxJbW4h0hO/nRQ9L8J4HuS4KG7zOo3YzC3Ql
kdH6+5ONPRPE4BLq0r4Ydd0mliFvYjJRW900iXPQIIeI8f5bSujkCysaeDTn
pweLfYT/5DU9+ukNWilmaIoihPAKCdtFJEWUSKDOP6xD0QGIgjWMV98HwKBg
xllDE+e/+fOIdhriaJzXL0k4rLlUKIuPhfmMQU9GdZ39YbjmHZNly27bNM3P
oW5Uqj1vuM4uWP0PyN36Sy09w06YSXlF30BctXSfRTrR2/C4tMOWkA1vC810
DX3bVISc15MVWKgHQ3ymjDbxqLTPwK/gITDBamr4onrIEQs4HMRoSy6Aih57
ai9hFmSsGuaPMXTQ8XUTK+QpAr0pG4T5gAsjw5MYnGVDPXEeofOeh0QTYq6y
AzM2r4niNIm1OIJF/UE6ml073toMWBbRkSB14bhkOjT3CBUhohZhzKTJ6a2I
zw46cU2ayyYol0Zwd7kCktWvFwB2w4F4F4yzk2Q1kgV3trp7eQsDYT7wu74N
LKNmxNjc8Kyp6hhmlYpI4voHhacLS17PNfuJiI4EzJ38RP5xyKI6JjRbS4bw
3Hye68Cgy0naQh9uiyr3FA6VHyBlt74kISsJks3qgQi/or/eFBnsJ/HGOlqf
25jEpzFBwZadPKPSSqv5KPKyOnJjc8ztEDZhkekgYAG409RQ5Izzu/Hf7SBg
UsKjTrv05TUE5NqtnLrDDHCPwBQ+yxkZN05S2R94WLcjxb+pU7qu1JvVdthS
6iWPyG8Wi/TvAHOFYm4GmwQ9GIHTJOS+cJHhIqb+TNtTWPGFIV9zYOgXWjMZ
xRBZ6kvPm2s2rvr7NZUE7Y10+5boEGxDD33Mm0+C+Zty3KAMKPg0dObifxUw
tDQvTk7+vMzVpuqkL5e9j6fA/E0/oqDaxmVuSwMaOn5koLWyeJu4+h7EKUWH
2n2XO6bLvoa1oJdON5o6rJgiFogGIJaMOiG/vpYgTMpqZ8R2oetxx1qmVUtu
q3gwrLJ9SwExjn5pHclJzH9UJ7LVyIzC/ZGYuYlub/vgBOazuTj+YxI0ORO+
7fsjUvHNwuMYf0NYV0IMBASPYwjy/eX1WienrprRSvzEY69ks8HbUyY7o6S8
u3Mwz6IH5lRqwJ/+hRNZspenkQ5qxKOgc46DJ+GX2YN8Z3FT2FOGShu3DQ4c
23ioeR8hmlXKsJ/QQeBSSaagj3N9jHHbxByeRwfhVTvmQPcZPSqLDbJWLLPl
cw92tYng9gqkkfz/XA7WBOBo67pvkGrrcBmCJxjU4Qak7Zk0UbHsv+bY5QSP
ExAKQtK9EpN1eIytzFSrOeP3SUkBYif3r1yy4UhHW8HatkjsrNQD1uT+2zS5
AqQR9cupn8YK4IRQNrnrTHv+EWhqopVKm83OS5AsvgZpx4+qpIB4q3f7548m
RRNYpduShOukFWsImiSLBMceJxq8dL0gkQmUyqe/ZeCKoS++srdvq6V+DPfJ
79dCjqbKXIiiLOVx5uIyGpqwMTg0cgPPo2/RWYeWEVBcr0BMFQzHnwl/GdEC
akDaeuO+bBMJGP3BHRgm24ADJpEOq1WXhTN3WqqvzERlywuXC6ibzea6CRun
Hdfxj+/7dE6dWneMS4TbSyglGtQUHaYdnjiROs0nJHIA9U5ET0NtQhDQaxew
f0m5YQFhBV+3Z+xf8qw2eKeLo6Gi8otrdxoPZrvnj1rRqQOL55gaqxH67AoD
Yio9zq93uhHUms/I4fmkjro7mGaJ5jMB7XSEULHBgBeEJx65W2feAWMV7bcx
Pv8PxgAmO/31e7L57Q+L/R15HDyZ9OIlVI50r1zC79cl/FZ8Rv3wGFLxCyNL
WEQhI/F5wapRrcijQiWLIZhVrVI+CrR/uqKmbhslbJuK+/wVRfmTlSVTUBeW
QVm1NrqqC92o5v56t/2OLQNU//UIsKV7ad/FPmb7JeS8FJQu/CgL+ATdSiIX
+Rci+cY6ZcXTUlBeYna6bBqVxDetl17camK/nrxnxzR+ijwrIe+Lpr5aCYnW
OYfeYYPNol6xSkY65ayDmjxKFgsCxC9beGhg+GAsfdsuURNKOUviUJS2vu08
izNnMXcXfJbaQ7ANHTzB76yjK8owbYD4ViFDkGvpibsTyLNpsocolgo6/WOp
rAPcEMICAN5m77UdAOJs8xVG7NWfoxRn9dnsRvM2JNqPjKG3USTHB0cJLOQR
W4I2oS434bzU+HDTyGp5z/6FCYvN/j/U3FSPZ2CxDjQGhEqAXPWOkLoYhNzo
Fryqz/8W49ptyjvyWn0PAculxPqwJmUGd8Uc3i46kzzsyvO4JBjTAEvDYOw3
/pbtnPduKYJzjRrSGrzff90Bva5KsTb4rD+zIcGWkNJGxK4gdrRgB0biD/qw
HQKODlEdPvPktD09Md06lqlDOyW0Pq0X7us3FAClax8R2fzEaJG+uDoLU1FC
F6BhWr86Uyu0MTdtRvKla5aeQBTCgVpc/zi7+Bb3i6QQ4c28m4XsbwadVuB1
FuEvmI1L42wyfSar9biwiz/g4lsM63DiVj8Mv1laKsIRRs4YW/fUifQ4IJ0C
93FhXNaGUKN3ve8MKKH6g0jfYpa/uHNAEzCeXzWJmGObZ/7fmQMPSc0+H1Jg
EsOWoQjV+xZ18vGt3SVlx4gJIgAi3PysKdpfd8IIjbAwp+05b9LgTQELaV0e
QpHjlw2VIwO1Ny6a8LRvIu3pPU3VgDtrrkO10JfeO/aPwNg16sjLQsEZ1zjj
+0rvRokpItQIfA4vYZzUA7orEcxHN/+RKNnhS0PMr6TBymhyZCDVzZA4qEID
EXrTdK2/xMaI74JZVUWh/ZSTf2cEdUCjsd1wrbmgWZHnM1Sr5BuX4FP4mR4a
P+5KYZiC+46H7Q8JmviBAEU3gm5yIvJt2aKe8rPJ3e0VqoEi5tytDqwEsNWZ
axxKGwLzosOaoHddQc45zXL4m7ynWJeNUo5/S21NLeZaxcZQH+4Hg0Ygl6eJ
83nuFvHnPFSCcV+iiogAdQfcx/TEGPry+OOpVnXSCJZLW10lOuRhgoP061Je
u69J4cMJDOAQg3pDxy9czk/jQYcUUSunJN1sFHFyI9q7zLyIpY2uX0BJaxTk
/GndnrcIrRHkWy8LaSibW/vAuGXCy/mychim6R97CGhDDax6vtMuL6lFaQpY
jEFQ1KZblJgqCqnfYcPueQQGDicRN9ocDf2688AnyPQmnwa2clX684QmSh0m
qzOlyhYKMGaUUMbREnfjyPGMAkaSp2pnfUkuoeLcoBC//8VNoCaL3voaCZOI
FhKNgt2E/RJzjNrLIFjlthBCApcQ4iCZESGT2lPheS6EggdPeJoEY7xrfGv8
Uzpc5msirqpOzdVga10t9afNEo60hGYTloDdxm1yjJ3y2Rqn45z9BuTS2a8R
q4HQ65P28Rzbjm5FV9wSgqLypAGBcSzH6UIQlH8EoBA29Q5n/1XihyUvpGhx
hAYx5mTx1tSUNumrpu5hyC5eN9PK5OoOIN7tZd8iP5VnTvJ0sZWu14lezrzj
DskAPX0SXt03aOjJ+cHM9lvbDbWiPvO4cC5fYwRXgkwMg13HcJ2LoRr72G2G
E09FdQNeH7HbyISDKUa4GyEHNk2xCEvNOx53ibT9Ij8/krCxsRrHekVkN4aW
TIvJordTYlTtXXGgrdyPTdFKElqkXsk+ieDpN0PMfJSHBJbB8qqbUE/17XP9
JeGOyERelBk4YSEeW8uzy8zRtjiRz/s9JzFoioQHefaonk3nI9zhK2Y+nkD6
yfYdjI1o5Au+4Nb7TstYc0h3ZmstpfM1J5EiB5vFlUO7tDLL0i8lCDqBu3fw
/rYx0Bs2qxcBeNjcDrtgaLYoO4xBZWNyxQaZEp6jyoL6OdvwNr6m13doDljE
7O/xRp6c5rSnwQ+6SPdF5hmQtXxUJK1rFRekzOQOiHXpsaox6cikt1oY/h2d
9dtgQSPynMJhJYrARYnq9ZqFQUPTj1kQOfSVS95HJph27UlElDKc04QtzduW
sz5MtWQ0TxEaju1K+Hz61nR0/pmYurdUr9bOhNg3qo5Vcal71zCQ1oA0N3Rj
ZqysJQn8spDh2MbkGHlo20X59ePnkMPXJabIv0MebnGt8/Yh000tpPgjgxG8
dxGCH2t9FQ+yL61BIxr7SqWeVMcl0UnuWXmKrhkns4q18ePNEBXgeX8v06jO
B7mxFXDjfAmZ+sXpPNJdCUoe4SQP7ESgCgPXz4lq8TsqVL8TgCPXBtEpcBC7
wrLZ9HOCrbMRZVdFhhQH6Pqgofn1j25o46hb20t+Vts3YagMLVwWjbKtG5F4
ps2zc5do4Ny+1pSwav2A+bEqk/vngkK9oeVjTVOlVcCbmOoCoGZhiUxCCQdK
1/epnOZqU3cnAS/V7zRUvUkS/voNSMq2dWtvx5Rcvjmivrb0Bd+De+q/Q2KZ
sb1Wj+dF5m1ehvOguE6VhXqv2dTmkPKggtNU5TjWoDo25ENzqmRz+doq8zmS
JL4gfqHCe6wHvpATXNqrtvgEovDGrBuKwKghE4JDEWbVpp5dIZJBfCOinq1W
zI0vpzv8zlsgGYdMriFhwdkHoeCW0Q+mkEqIhaOQxBg3HHPwl62vinERQGCn
2ju7UHFgZO44Ev+JTRE/pXon7m3Gv4w5FMUO7KSW3Po60iXC+OBiPBseT8Sp
Oj5u6bUtEOWpA089zNmsnyiZ7kRNw9c4XD7pdQfx1bVxb3xHrTYPLPot3yHr
ccjCXiN0mzk/3YMIWesIHmqmzZfpLCL8DFBCVGCHKSTzay1dfeQe6WkOyK8R
up2zISqKbIqHYAPDT65qhnAx2juKkeRQAwqbNcKGdFi6Zq6BeAzj6LknCy06
toqiSJfrI0SY1jCoAJwhu4qju3wE7GLwtYn9t1Bj06ue2hqzfEolJzoUevsr
vjoQUu3oKw5Xl+U00x9OiM+En9rWs8MKMVe7N6aaCuYI5iX+gkY/0pRE/D6f
BXm/2UFQ3Y9hUAVjpoYZ+wpNyslsw98yU0tMVNFnbRQha7LoceHzfoA4z2z5
XipJJYg2a8L0JFXWIvjGWtt669BkuZg+2GjhuMgKG8+zKXrDhvTCAX1ZOmWL
oWcUX7ZM3SuO6nzj3P3KzVGsDVOBYa8ds/OXyMMgu6ldGA2pp6lHfpxOlLm/
h4lwaGKnQcR1N8/r8veVD0saAL6VdOq/CMapdAtmT25/7wGGvlX8fBLjY1Mt
qQn5uVd8wZsXvK6ODdy2b3YRg6YEs9hANAHHHs8DTQpHloKVsBwcYeZc4C6v
H8BW464439YtvLghaXid2Ny+++mrBGwC6AoDGjID9mKj9mk+cTVUxxfweh6f
S/Rj2R90AHeAPSv+2Jgl6OgvUfb8+yeJflt8nV9KUU34qx+9l7ujRxq1rMK5
mq6l98bsPWhPpR9z7i2L9HVPX8M4V+uw0tGrEgoIjEbNBELPRviw4uDVNTeF
UyHR/md7BeZYRZY778QTf+HegZQWo6SE3oM0unGTT/8tKjnr82j6Yh/Xh/6m
HQbpHGeiRgYHLwvJ8zbmIKTAuvWrJZiksJrbLrmxlwyh7sPiMdUKrl9QIyBu
3Lm+VVEO2jFsJl8sorWAZNSsSizX4r9zg8SDYgucNsbS3QZdrTodtXHME90M
twiWx9D2vzndvOIufbwA0GVJARjCLk6YNNAxSwxl/T8hosRimCXvwnKbVNgJ
ughRHl9QQ81dpkx/YKj7jraPtdysXkjpQ3ZvNFb3/0w9fn7aO8GfNjuheHqK
JgsC6x0m51U7/mWDFFtPqsvdQg5v4MrLrqG2B461qHRm86Rt4wphPTErHM5E
mmRDigVvmMJak2Mn52wNcVGfZ55OIVPqbvMvSYu4qR4pCZMgjoICRqDBMN3S
ZIivODQuDY9wsLXdbaXdmvZQs7l6z1VvIc6yz3K7kHUEqx+nznomX8ffwGpQ
NYGi9BaSjNO1Eb0qA1gSGjtfsypYrhs3HoRqbQ7qQ18PFPDmHE9DRNroesDS
I2yK45zDiLxu2rcXfy2XdxLXPfa3M2TVhCAd/Rh6VEbCDGuAeUAP0Lwx+dJz
9c8DIpl78utnZgO6GW6zy/hl6ZbNOLacNWEv1reOdqdVFUJJ2gB8NHMws+Gl
qMjPLNXhjF436s4NruMeYXMmtH7sJndrHGBapBW4p+Ptc18ElxfPxNkqij2J
L+05+P0pIHK8neke9jR43xxPYqrfEY1eCFZqEzs2DE5RqZvPnRJo1Q/MUT0C
D8YsdFc7eQH9cBrpsgHpDRnVckEMhZUlkaLYDKHWGWE2rRQuevYC52jL5AEJ
ZQHerHodFJOqw6HCo8SZpeLwqIWmb1vh8eG9Sca1JDG6IolzFtIIX/PeCsc/
wM4fpTr4Z6GQSkmGsGGkpgrzQq0hVa80G06LH/Gf4MpEzoq2M73EEX2JkQ9j
vUqEzW+exV+Uo7tR0RXq3w/q6RtbFek+tJqeJf+9fUmPx9Cvp0l8oh6apEk1
GFrWjIT8r2cn15DVg1RUZT9mf6XW4o+U+f8CS2eVedwVj1/cNsHQtziNorlR
RAI/oTmVf27AvCewT4xd3lEiUUXx2+IO4NrBOE7Kl1Ot+M0AVPKhcsIkmQkM
nLntx0BzQCcnCH3afPI7B7sL9qrgsatPVxaHqCU6+ggxP1DWRgPUaMxwbLcf
ExM+HHDo8/k8332LyPaevWwQXSyV9l1xJKm9cupwMvBCEzygp64ujChAP3gp
0aiGo+knWTHuCd+932me02US7SVms1P9zqLf+aQ7XPJ8z382+J3kUYCkEmSJ
kPA6L4wSxu4rpiniMGEGPQTa3EbSnqfPo5Io+SXFOZ+xlVCdSaUVCQKA1yqg
wRvGPVmrRSyCghLoIIVglITU/KIE1VwkKc85jguE/W0x9uhR3IbQzEGRNmGb
bDA63DymaPYrpcfPWsiWAEJ2dqVBkxBNsdRKzaB34jThzYUrFrCh9XIAntId
sh8QQCI15CjiF4A2ZofztiBgoVMt7W6SrxQXul7GKbyaGx5Fz4Op9mnQybKi
jS54wu1SU5S7WkUTikQjM9y8S2tY3hgwpmhnZYDCfjyUSxh7fvL1OjVUnLn6
Fo/4+CE5CX1klYe5p/6Abm8mRJaSsdc96c/iHwX9nboKCyAaV9ESNEHMaF6n
z/8yd++fN9udzybZIY7N62D1MrA+zjVlK0f8yQH900iocpAqDCTqDfuYLbCh
DsLn4/BAVH+KP5zqFMa3ssXDjYJDi+9NJFYUZzRwrCkf16LCt+wjFv30MceX
clAz14tf3cmks1h7yyUXuDDvpITyiwSO1UzOorP/J/lHKEPerK3zexRyiKUj
WZGgvs/+x0+9/2B5/vPk+I9P63yQJW3YA5HAgj2oZKOLCyjQfqVVy0q4yHu3
s3FSRqwWkNIm9YZPxsqgLPEiOuO1aTsSdGvflfTAoBrZp36stWsVNfc6Uiw4
DFr+nsPnD2b3LU8WSrm4NImlnUHlND7ehUEFnJRx5lHlGh2ON4wMYrVL2C3t
GkQv609qx8lZ/x/u1NNjHnkAr9OJqMuiW/6tApAADVFbyE9p8iNNNHMBdwGH
3zp42Z3PpXIy7+7O0gBzqjGAyTUQAJlhca55ywpV2GwQ5/KdaPJJg693Cueu
0Ufjv5rJWOPiGCUf/8+zg1ze28F6TG/rG2ZB2JIudIwGRoK7HhNZElRVYTEE
UjX+rKbcaF46vlkZ4BHheHg9z5BoJaQbtklIWAcoLff/fd+L24MuHRkHlfT6
3VA0iETB+87aOix0t5TZGz13RCwvtk+ajoMllud5uezJkJi1RGbtEVMeGlSW
WCneYcueBRDRaJK+hhfDy7XVf9uuVl3PvTRMaieJ038lLcmBQFWqCWsPqeyw
JJusXvGhE/9ndBFKmfPXAOr0uz0tFWhIv4Pl5Pzw707U2ANuq1tXWSgz9rv2
6edebgE886c0R0V7gXsJCjBYk66oywtOa4AA41vpLYV8Bi7hacx6aU1fYd2y
FiEi/L2eSnAu5AYefsb33vTGhdXnJe7zxo0w8oX01P3MyerUqbKYp/kEsHD2
HMil9Tiyby9CLsA+TcXPhjWdwTQXZrTymqR3Beyd4AjyDR6HnJak5nGGMlgg
p0ETOP5eFyZ3xs8G8NXBZimo9XQccDgsMsg/T5BjUbbU8zA/QauoDGKizz0x
HzfzxdYNkU5/TUOBqItVoexUJm3MT++CYFpC4mysCx/9TCX8cOp37v6GqzVK
7jbtNIFZr7m5gIctVKnsftPxT5swx+qBi9B1lMcWOAm0ezfIRGnFqjfC6YKJ
4aC7TW5NxvxeIeHSTzncEvgWlCEg4d/8E2xKgi5X10z0X1p4cnFXOjpgoy4c
v1QIx1zrb1SDlJQEjFRIVrZVr6AqeJuL7KgST/6LlHxu8YoJLrzKrz3lYnbu
9xmdAOvJ/SMvLcZUvCPVuU1ys3ADmHkMwjsU40l8/wiIhDan5XybV1aGVomN
gtBS0ggxHyDtQDAVtpWRuNAsKlmcL1JBte15CYUt2C7eChsJIZlJnjoif6z8
lei5fEvZkbF1aoNqO8NP0RvXEnkw0oXA3JwZQ4L621Shojhsnrm4K0LJmxn8
pV/6v2kWqTlAIp1pEE8kzGJScG9hbS1lHo/9RGw3+xoX6lzc/uB9tpMy5sMz
kVUO8KY2anhgzdLRtqeNynmAUe1bzWZLgHNxHdbnRJ/fGKqZJaLBzFSeEFjw
4oo5lwHSEVC/49V2z1pDmHoB6e5o9IU7iZnuf6EBYWcKEAd7P7wQuPfNtcOu
dl8zi+bjpltTp7wxoCO3uc5T7XxgPxihElhPqP/neqz9Wa0da6YFVhun8zYS
EIc3Oix7aeyBXxUxC5HAtK30VCUKdDwQnZ2hrQICbbRaWU4WPenw0lWrZ6xo
DgMGxywGIsSbV1TOZedsL70ruprTFQVbCJUTM0yOrZ4+pYegPc8v+yynV/DJ
JJScBPP6w2Dlzk/mshw8oGZw8Z2WXj8YW3RSJh5uqntUoiB0Dp81fo3Zuqam
AgT+MwXplzs2JsG4wGUgs9sJGUKJfr3nxmwBtQAppiAD1GipN+iAcllHv3GS
5kw/fXxZhBfE6Z9MHjV8Q2UVHnVbrc7iwVhGp54xIse8LM9/NLJWHq34XpcL
z9l5MNM0eUC3bKHl+O/H9YJq/sWB1l3llRkMBoeXBphWU2lqRN2Q01q27Rpm
Qmv3ygNJd2Ru42U1GNnPZ6/4+ronQMvFG/TmQmOaUxyuPzRRsP8vikIPnRJe
eCieCX2Due5Z2bZEHZXO+h+zsmZgSGDQKr5wKvP4I+trYztkQlgatXJNkyvQ
SmgNW168C6XDk1GhDFBb6qxFekXcivTuwkfX9CYiSVBKwFpFZnHHdWF1dAkJ
9kTTJzDBhwP+uqDL/oVlOuOz0YDErgIX9y+8fqOKEEwEnncl6PM4cUzWZLDi
lwyWjTYKZbhGZnK3NvEP3zWvotPoabZoK8gfuoc98deqBcdPcAoEErUaIUAV
Fcby9hi3Ey1+rj4rISY6x/VOiNzyM84iNGV91kvHXUHbcajjjUAjB/v3ANqg
cjE55w7l+AtD4VU90ueNQrwYLo56QBy3llDltISx/1+NpJmWhGVi/ffJO34n
iYQedr9+YmWg5Yqe/VYUV97SbeqN3xlSSD6yLNGCb5Whca9+QWvYvcyHJ6fA
OQAOxIEEYny9hebOsr8zRvCb42hVzfQp85TFTIQUWOiqd031Su4ICpBgyUrF
eZtn9Pas60YHOHqbgKZAFBD3jBZAGi9euo2DhGcJvEnnajBCnlQndeFo0wJV
YWDot5+JDh8jl3yOa7VVdsjf0fQHLLtqsrtnNZB6v49seDMQ5nmu163+lRO4
6KWiLpoN/QSMad4pbzAuBQc/JVzFQ8VOTDYOZoCZp3/hDFQgkIX7XDiMkhFr
I6SMkQcMf5Q8jRipBR496KxtxfhVUuXne1Yizz/JafNfAOxlj+2dr5bH6AAB
s4VlC+UzGR5nuGmynNPHONOgXnAceWOZquajOw7UR2ZsDbqko7Iq/Nd86f/N
yS/o02BOhsjLO7lU+PIa4q5q9aCRbLJ8iFFSe+AwceF3flUVPZBUa2lRLvh3
AvvbkVnbMQzj0oPkkC4GWQksghW4gEWe1MbrDdeghYsaHXs2f/YvixMg2Cnt
iQRezZTLilWjF5tYEgDPaZ2Nk6OBdfyoWbECTy+ShzBLyDD8AbZnWI7YTK8z
yZGwzdnG4Ali6UqkKJ11JHKObHKnd0zYpuynGyf9NEmaL3WGB2YXf2fIitLy
KEnwseLBeB1365zpSljXGdR80I0jMyKkLoyJ3VyMmeE7Dzgl9ke19bLaq8+L
JKB9zuuEGj1qg20EjUeOLMYR14R/wo5MfdxtzVdUC+GKAEoJn4WWphWd03oN
l+yT69OXLfj15ONOWzyKgx1xJ0SKA2tPA3Loziw7HvIgYOSLR+Oyl2gloIqy
5ABEry/xkckNkOY3QZwssoqn9aCIgWqN1x1GdI/1Ve4ZmdwsNOdNeXUisChc
jEX4wqoIKXDiza+qSeDWNB9PPuaFzxi1WbXpYqi2WzlRJliMPdNhqs4JRQVq
1yXMUupa+6yKD/JWyzPGvp4wJnuopg3aPjFz6RdrbUFLGuZ0rmJ5KyD9QBSo
BjKH6BMg2f6a89Gi3mpvGTMblwjDPBKzgy1LtZUS0jK3zwKjEE2ygvjaYNPs
QjmhzwqfVnyadDf6IiD6ZZO5NDiYBVwJOWu8kOk3Pr9TbgaO0ssFvpe2E8wD
rh6lXRk3/cTorvjmVeTpoJPkkYI2JyITWPi4iH5fvaGLIRjuXqUijS5aSfQR
9zEg0fbo/tM2ZuepbQUKZqSqm/fSCYHSq5v7PUSOA4PuyCEJPyWrOPi7X9Cu
mjCB5dEmij8wYRFR50zGL1J8fzhmxmScdV6MUncGCPNeC9p37cY/S9SG+Xjf
XTEDsPf6pzePpOBuvrMUqaNcoJcRQaXcLavWLNbOrBxQNTfDVMGdgQvWrfl7
2ziYp7NPAl2G5Jq8+UDGCYB31sKrP51FOMYJMsQBkkXM9yj0fRzBCqs6L5Cy
DJ6yAqmBdOiGndvlERCfrUnzbptdnKaMMwXTkJdPSUFtSM8NZOcM07wyixVV
33SjCpOWc1hULysiaIKDLLCzhy0jU1IsEf19cp+w1JLifpeO6Zibc91MrT/N
ffbxyNJ2i9DFpXpyr3zy4YWSF7l2cEvsoLoztOGMtRrEjQUfD4sOEymSG+Ls
G4mKvVczYHhQn/gJA4W18XNpzY3hhk8WnggelnFWb3QD5wznkFHiHzQ16EqC
R5j1kR2s1WZ8aSS695cjv9XzXTomxFIwytu7y6nyMmEb5WnyhnwGb9sGDwQF
zv1KvRXpPG+RfLFxxVti/rzpOj/0H1q0Q1IpVQUCg9uVVWhlZPT6SeuHcxSW
pSCVPcgbFS0eGf41MRMK3hvtm8GPISLXhkdEjkarVLDU5FNsHXqzhpkzJEav
cc2cXjpqlawLBILTZ4uRQqkbVlpVbtUUaZ+M95ufnInDVv+i2UfSEaXlEA0T
q+N/T0EMI9SP4mQ2XL2zzO1f9MYPpGesrvX7QRk2x4ia5J7/HP0G7Oy+tP4k
YqZhyhMUd/6tFfeDtUDJQNvga/bS5856JXUpY56t5e1kKST4kmtegSkR4Dke
5z6dqZKdKMmRqdPimRfJh4iCEMUz67ARKBRZt91TUmx83iKW1AEhMPXte8+Q
vZ3O3hrxRpzLxCk2PhzXljK1nWND2OKLihmh47X5Q3aOVhSA6gEVm8NK6ln4
AvvDTlh7OKjC/I4qRlre4EcUJg00CxsKKqNDXsXF2QLbJR37gT3IpGHNBWsx
tkOWnprewEnKxZBdvazSTayp3fUfPKi7vclCfQzeaYPETxhwJ60If8An43X1
KHR4OH9vP/mGLqmj5G8WTnpZposfKKsZo8LNhwjiS4aGKu7kpO+Uc7pjzeeo
1hSYGKCX0UitBao0CSAJYXbnDHW9TwC9fJXEvj4mcrnyy0W8mI58+NZCct8I
+IaNaF9sM15I8x6nV91pLvWAM08GC3ZUhbQPcYAAonUn834R1xv8XGa8Ni9l
FY+0zeYFc2P1F+XQH/ORo6SB/uwbBWinna6v6tuzV+Ii6WnHu9B999zExbHb
nPAJLCymQHmBnk3rffyDTAGmPKWiIEGFrbCqd4EEnmoIXLDA1o3zCGw0zE9q
UInsjgtIieoWiE0A176GKDEUpC1dX2+pG3K/1LUw8zpmIU6MImBX6ptXH8tn
BZsuvVqxejEDXW7KTYBgSKaKLG3s3hz6pED/N9rMQewsAN84wdv5ChFdj+D1
35p+kR2cDOvOWz71YnhNh5TfnO29nea9Wvgm+YORXKz/A3r9pwr8hqsdjRJh
8rc2a/kidJpmbQOz+x+rCZlNRWPhfmaaDz1aLLvjsIGJhYFzVCVftdtwk6QF
NrVq2BHQhIK5+HMNLergmpmaTHiYmxCXV2+THS8CpSeOpwNFPKmqvMslzdgU
HMHx0zq1/YutZzmJVEXPRABqHQU0jynUhxw/hO4rDrb3F46qhdRHG+d4MGCZ
QzTJwQ5Iq20Y4rEVK6hFl2ZOS8a/22y31xgqdybmhtJ9/94KWiGJxxhKK3Hd
17QyRp/yc4ZF/TmK6uE1O21aIWzVYRlBO7PmRbqSbTlwb6dH47aC5wQftDdF
VLVyg+ot4OPXvjLus2PtabbCip1EC9CkNz3Qql7LrCtTpEZwqo+8ljFttGfX
c0jxE42bJCDuBXPhpHjav4Zw4uHzS+SpdLAwFknqOS1+249/74Xrj290xu4O
SGjao0ZWpushNES+vJehIxImTHPSHvnYNuONlrTZzg2wD2BMEHoMolSxZi+K
K3Kf3ovOKE9RoqZqyGgEIfI7Utgzi2SvpTwKHnUg4dmdXO9+fz6CU0V5Grss
DDhq2/B4mjOOb1Mfnh6NRHyZa+HSB3K/JVeALf91KGJr9vp2iDzP3RCLJeFI
j4AwhyNzYgHmW5WINszRawZv5pSRJpVLaaGLveSiD1ZQV5qmfLDTmUaFzZyx
kftJWw/HLD54FV6Mt3QCYfygzOWFCjV/HcnyhMGUIlSRb8nlPckQecBZEMFU
87rNof9huO6vEGz3UYgxS/QFGA8E796KzA6iyTwrVgz5qUHTkUzjXX+EYKiy
Sz3js2oqNARQgdte7kwXFRB6YVdarZ99ovHNVQpgZd+qTypqzEefU3V/11tr
TZytV1Oj/A9zT2xLHfLlVVDy3oNi7JZpHK+9kX1rzMzGtW6GVYuyzwaSi50C
x8NzbXnmx3M+117R5hDSKtLtW6CxHO7FOVV22NE9HwFHUlvgJQX/w2FC9o2r
OFA6cP4PZWtcLkadkneg8fv0ilT/KWY3O58OBA6bBeWkvz7JkjvSUj6ZWTld
bUHOI19TVNlFc0P+0GgppaHTIv/Yf1QBdPARuUm1EaYsX8mMX4kf50xTOnVj
kFsdsOTbn8mFZ/NtMW/+7nhLxiWuGqRKXXNhWYWw0RHx/Ji0OCt/u416so8h
DpjzywCaBJ9Z99fwhg4aoQgImhIFk/whniKy7librWPLCFsTLGDchhea7Ezs
1G+3tEyO6s/K+/HoLrPiET/VHiqJ+NY11m4lbu9IZDOvhKZeyhUofa6xGgP2
kxOiYbinlM6EyJwZgy0ofm0lO6OXsBGGgBgtAS9oeXfB+7aTnIMnofX1h2Wy
XSNnIjhawIj+Q76GIBLjnhLE9CN8OIWL8jzXpy/nmrNk4NCe6mXBwb9SMXcd
kWMRB8GugdUGXGgNx7jrY2FwPjG6AVvH5RAK5FMrVSV2YB4QR6PM1iv74Fmg
aqlUPK6ddSXQ9Vg+0ugXia1sqN2AURT+hsazEUAC+h0PwF2E17cIgOOl5N6Z
Uu8nSANpxucVY1uGmhoFAb1Vmf/hDInALnwsxigLmwF+eDJ+xg8VyqxZg0Em
mLFyosfDBDrTw4p64osuB9KEvoh4eiPXNrbE0IgK/Bxbg2Xdx2z72xWja08v
w6MQFnN+GNSdjYb+xVuz3G4XkIK4TSWBRkSRSvDJW3DM1FaTZpl4Lo59x5Fw
hsu3GFcmhd7y5zpL2dIalT+2gyh3MIzi5DjzOpGatO7WhtvJfUwQAXB/FKIC
XFO4J9CsmLDJPZESdCH7STGQafVacfQG0qW21LB+D/v2JJZlzYLIwwg/yKl0
vNlebfDrOQR++vYwjd/0EPZdOHVBxZXfoRkZFsCGXvMWDYVdO2pRAr+6aUgT
Nb3dXJNUcI1lObNoOS30KszBK7CFs5aTnRQ9MTYNKwnxvFEoqL6ljpEiT/4n
GyGjKFDOdgKgiuZ0ezYeT6cgUCxb0WWc6ic6QASEQC7U2/ksGR8zOFABac7B
D8hy8WLb3YqY356W3548DEb+5G3agkEyZdqdVD7agX7filZDF4X28j2hFwl8
HJm/MfPRzys6h94AwoRJcNWVANh03Wy2MpXC3aQsqRzMxLWs2iAdbbg43gtI
gSNtisUvNavlP9ZP9Pmoygi+ppY6gpw+DWYtcRvyhEb4fAdyZ9Bv3GltyOdO
VEbIkVdosEfBIr5BIX1qp1i4je1wcxYelHO0RtfCoNj5mLs3sOtr+5ez7Aek
YUnyTlFQXqUKe89z7ZqGDRo2LMCkLUhcsiK83aUnZQ1GXfQUboBgV6J1WFxi
+Zazb89nr95cicooV48wxjDQCtgmw3/UlRl3DvByHvez34euM2/n8mCshRMr
cPWCs7xWQ08u2t5naxMLTHGzUf3DIFDXtBvyLo7FXYzzkgQ8pzg68QZ2/B7z
amMReLXZiLFfkQ+z/VbZm1w9W8hblbJpVeGKGuGQAiqZ1QZM0NUoEv2vV5nV
cCN4OHdSsy7Z6fCv2GGGHjvzUb1OHB9VZFDqOlXtXarICyyyvx/MC6kNj6tp
wZ9I4zgU7KYqUBOgHVqP9iayTjgQsV89zAqUns36mH+kdTI03lLHZYgxIT2c
PBC59SQxteoHOgcfJwfNJco3OPXGhtnvfNp4DZNUJnHkSjafVaBVRV5fYAHP
mrqP3GEuFuNiMjiB/+UK+sr1dGIyqcDrIcTNj8HKf2fM0wzcmeVvbSn9Rl2X
h+DqLxe07XDbSSJwaZCewXyZbxb6tij3CXPpTo43Dj4B2LtzBNpsJW4eqSiT
4gVn45y6vhQuA4CnjebauQnGFJpI4sZSDuafuydzCN58ac1t8OWoXOb5tnNs
LWW9m5PHOyeltmZeabk93FEHyaXtc2c+rq2o/bq30KbDBKQR4m0E92lsfw7O
rC/7z269Q2y61mdrfOaIeEDfIom/jgGVA5sbyjRt3f2VQKe/oxy/OjhmPdtD
EaZwwGKAHbHsuDAnqD0V+oNIL1+42s3Qhf04MYqj76LP3iK0QZrs9Iuocfu+
s7q+wneZy8rL5F9yehwPPyzmh5aNi1AHLHHYdSg0fBevTXKtRdmpZ5dDC6/w
N2eRYivaqlDkwS4hcazyBGi1aPoAieUHriITbf9EFuw23jxntaUi/xBiLG4O
5DoQ6LOMs2X6fSqxmXLd+HKMh3DJAd32WZBna91GPeuG/11KCCTXgHIQFo4U
4FVPifciL0CBSl8Gj6Q9LDmZXhJ1xYkwwZu9f6D+TIQPCTwfZc+YuVzfWBo3
go7Z0D1i/B35HAwtqm/173UWXW0v1RWCo3tlHybH7nvEJfx45mH93RQH6KL1
VWLUO3ROaAEfaXyKlqCIepAV+w+J7KX1D13qlm/nN5YeI9PaVEqWgONhkUBL
Mk3Zut2LIuvqy3W3yCOG9ptckchEHZDPqVy093w6sFRAxmjBWrz0dA646Fwr
v2LGUZ3TawANGHOB9FKmFoCaKtnlR+8cUAt/S6FhCA20qTkfC25w0i7ZCLZg
siplrW5Pzx6pXynkNZwXAJerx/MORxPgnrgoBW0rdF5CtpCGin84Y+3BPrNN
gg3SX3BQ/e76PHitpuDNziIAVkjcx1ezGU1ks/UWMvziGKT019gAOmqjWOIT
jsmxlWB7YZukgb7o6cB5H04ryMsdF3eqtBRD/G7GQwh2ipEs8kt39cMpEFm0
tiuj+4m07nqcAaJoTwyt4bLCj5wY20jHpVQIeJQrMi4oHSXWC4CKUHIvyEGq
U3ltL9wi+I2oVB1zHWQwDjveUhRHS4qPUlr5C5a80O4xie5SqFtqV5B+xf8Q
oaMZn9kQAzkScn8cP+O2j5uxD6OVr1ncLyyCJM+de3wBESH+sbcORwA5e5+5
oJJKrVhgt2qUOqQ0jHUpyyEoBYuf4SZmTpk6m7KtjNCMPY3gTotnsZQLh7s3
8rmyl9t7sE3cFC75AWpm+Y9lv++vSogTt/ebhD1/w5lEk4yoeltWNHplmNq/
jOJZNxMMmD6LEw/pZWLnfkSDfrw6QXHWRNJ399GpMewJe/kytdQYyXvLC849
eVJj8IgNxWrcRzu08j/Fig1v72zCwX88cspgpxsFylPVgBypPo6ED9b4u9SD
ouj1Y87m8IvZyOstCL4Jz402TvZbizYpUsDEX6uf3/MJ8rS2+CV0lUBvCcBG
S9nTlv4cjpokgU53iORS03LsF1j+pvuPn+T3gAt+75snNy6cSlG6jB47YS/F
TA68hI6J9YQiquyA3Rl7GPd6VW/YTW2qa4UldyYbEA8WZMMj8wqjJ/Lq1zWn
WYZe0oh1WI/aiZMoIo4x838R+3tUSC6IomQCYuTcVcC07qMLTq1OX2c1xesM
HgQKnn6L2NPkw8Q6qG0gDSNdWKUdxtbib6+tz5Ge5klVOXSuoItYaQet9c4Q
PRxy3K61lSEdflMmtGal3iD6jdh2sAhl3Ro0jx5z81ZnGejxmYZsH/OMKTGK
rRfVpu37At259r2s1N+R+5o3hyAfLpZg0XUbtmIINfPeX5KTNPRl0UgrW50Z
Ro0asplRqvBIs1HPQPtwrBlLQvIHk2sWzTUPhhbYPme6UMwNX2k/znxuSndE
2oxc5W69GGoQHrWrjsr4O48sBk6RZPfAHP098jWZn0W5SbPjPOTAQ/6m+qfB
YZTJLsUi1Nb9krGjzfkkKvOTb37F5bXmA6vaKFUfikGukfHqT+PfQ7LfI+j6
/fM61E4mPW9M6hdQ1XLvYtv2QEqXFKSSG9HOW/CuU+7IReaa2WYE8wqJckEB
W3tOdzIoC1q/jVF0FhZ7YC7IQBw/UqeIS4RbChAlSU5HyAoCeVQInggCjgE6
Y+ph21hcv306sDwOknylYTCZ1//X7qGLhSOk8eeyCL7w9tTIL0N9zTydGqFJ
CMenSodwFEwjciTaFlEjKzKDjk5PMlQ9uPPIAMkQZgnN03dhgMA7RC3fBY2z
3LD7AAHGa5ZPKdipSL17ScXe4GfKoyO+zdUwIimXt6j29gjbcgJbbxkB3zFX
yQzIaN8wkKsNnCknPe3QafdcCYIJXpkEKvHsuxi83ROM2u1AvrZU7Q52rEhE
HI3//z4GszHElae6n5BsvmQh2MUUALgJjCUQuDjgVAn31R2as02XNuc4fBqF
5EnDXOfgl0atUNbrLeKWxM5YsglbcI3+Zx8saWb3kDNfdv9CZ4sJQ2eEQN7q
te93+iEphEmeCRKbkIby8D22vFIn2M8FQDz2Ar5LsB5tHs+6TxY5E4r7TziI
qZMPs5SwSSUTREXeOz82zwu9SVEOn583zwrlWF3/B56vnkfjNJrZtQZK15U5
xyUay8mOQyl529P6BV+FiLhb0K11F3HoBozp0xk50naJw3P3VTTnexZdgXkO
pl/1eHVwdB+3OM49ECKBYExJyEB7t3xg/GJ9c3HDh56H6QIZAPjzsZx7dv4L
en+e+HRySRV7T3nvAR1g8RRZ+mD0CekFT/ylDgz6wYXZigB3+N4Z9UphWqJj
HmQlLAaHNq/dd//5N76JCGvkJ4E4oDRRgKYOwbDeJJXMbg6ULTJoeMRUI8KT
gygBQamFq8N7ti3uMOZaaKUVB1BbTJTNlsTEO83hbrRy73vIzaXBC2sCPzdI
w2qwnMldhnlnQIDEwNI+8C+f/LnNF5vKhjkClGvyAkrb5cufiyrFLFBMsIUI
EOYuIIGNS1rXPxuavGAeSqjqcL7AOfUZSJ7kU799m+uIfUUfBbtNzX9qfpa7
wvEkF/qLPRCJgmF82wqvFlateLRAQK9SPBc5NfAHFVPjRDd0jfcSFboF46tW
YRJZ4YUoPwr+hTRNqZznpThmpvyC1i5AyM8jsPPr93h11HD4dFbPHnSwmdzG
mrsrmKZTPlgVvqnxQzAqS0maSVWFv4wZOUAgOB+RNYpmeHdaKUjk2lFhupLR
MBn5vRiNK9QOxEbdgVlZwzXJFKdh0u4dZc8XFVF20VMpKLnkHbc7mhDBczzg
qZLkQkPlyoNqnh1FxH2RM3Dv/zAwuTDhgANh2LVUNB4K2JzcO/Pvst49GvrJ
LXpOxfe68u3PpwGSVmIiGwxEQPe0oRUH3xdLuL+mMwq9Yx7W6CYzdtPgvb0r
P00NDcyOug4v7amhTPiSlXYfuP2gofcNUljwtfFLAjS/hxBw5n7KD5BKRfmY
RKjHuRkLNumwQwU75VQKyoWOxRO2n+tyCgr00lfcTxypi1DLt6pWCezHf3GM
Gh09o5auYfcxkQA2mp+8CgMv1klUyK4KXljsrIaJgEdK3MTKS63Hhn6rG30E
tDPl8SLtV3MixRxiwKOKDgfJxmqAP2NRLHugjX0G2MdkJ8W51YBy4jKtnGQR
+Yarjt1j/W5Nn2sAG8cQlfUqWh5+KZM6tlx5+pA8u6eQZMeIS/KUL7GFGVhE
5cGFypqyF2x3vfyfJIEMfni6Yud/yOMLigAFaVOSDBtGGM5mtKYcEh3XJJ5L
bZ6GsVrRu9vxv8cM81oZl2DjChKljseIeBmmRaFEdNOvf0qurMYqsQ6T5ctx
cxiobwacDLGnDgDfhDzflALoOXBKxGj2PYgKsKksCiRxA8dep9HtfrZ/h2iA
ypxf6PgGHG5nH8mI56wdVDw9+JXZOYzUXaERa4JjgHutZfkBqKV8am9AfEv9
wG2IUlJZI6rxgStCZEgshEOcA7wS0YgIKNyIonZEKpQJiu801uvN+h85UZ5F
1YLVNFDren+TAzgn2APQ7Au3T4l/R9fhD9WeMlPl7NFWMcMU/QBWWyAI14df
akUnXp1chpvioa19oVpaKakkmTLfC9rlXpF2yfQ+ClHDmeVbRL1szMasvnLD
UqvcftCF5Qm6xmmj5+w5Z0cd/Gzn15xBrX5N1Fsj5ni3ITRdDGyRnYhPaNwb
hT3s+iegut7QdkmMG/TF8Mh9MfZCyU3kMPjjdICQQoqqGsRWHglZT+NHffbI
XbSqYCBJ5aftgKmnceSetHQGomUTQlX15w/CZdc3RYwcSxmplFIO799QtKX0
EBpz5fMQK7k54NtJPd0tgoYMJqI7wCZXaAWlh6t1O0DBViNHbfXnalx50JHh
XZc0QhwsuMyCI5jtRz3DlXyslLca1p6dZ/W6AksPvMHX5VL9m1pJNgiWpsA1
AxGqfT9Rlo/qrB80CvxLpHbHsloMiqQhrlgNc7k/tc/y7lS4U6ruWhFsiSgN
A7zrDbVObScEZYGSbrF+e+IbqZA0ss220pBQd7zDUxvfoZyO+t4Q5mcCC8XG
ptPpZ/QZze76lpjprRxJFdRyttpd9SPXJX4ZufCgP6pn++E21XQFMl4gIYi5
d4GWnhbNBsC4Zv0OyZcSdXVP5OjFbw1TELdmSogBMIOsAW5AQWbABJXgpr88
PSATARQRvInHq/wUc9uj9rOvCyQxIywFuAh+gG555Fmbgg+FZv5M+RbMIoxq
KDx0HozP0TsCYKmiAlK6TW8yzin09ISl8wlOsVrsTmIOpDaLC/sJtUVQQ8rE
yb2VLiZjh4TjERRzCKNvOHDPClzNOVxoYqCL4Ow4RSE220we16En79mYeYRZ
NMGzKI9O1z24a6jJboxgljhzAhwDZuPf6FD9xxUGYvYMne+lp82tfzpNq9fn
ok/nnZlyZf2tkZPQFNjjJ3ycCVV2jLaXhK5KCKA5yW12yAuf8pnDNE9Yd3e8
9jhXycWUG5aUGonP8vEGDXhD6fbIyxJdptrB+f1o/5CFr5WsoSpMuGJ7R00n
sSu2SUpJd+0pz2kCkRT3elku8JpNnX52U19IuyQMiUuI6YP8DKAfKfCbLijJ
DXpWGI6znv4Eoiy+Ke1UxQTUgrJzfHlCRXCFdbVhTVSd8wFYMXhU6I325tjx
uGT+7fZPIVZotRzjMm1RM/H/mbYEgeyXCYoWDxXd3nIx6wLKlKUgn9adQmbu
hCVcdw17XT5v1DUKCL7g0qkU7hY6iFnzNcuQAFgC/kuTYlHG6fAz78razCxG
e9pvLXJGtdofTlXAWievW5EjjnVyPrwmZskyIeyMjuzkdiq41r3mo/IvSGLN
o3HEeDduCXKj4Y7TDs3tBpUo7/yyC2zmb4sW3t6WUAm2ea2/po+UYQUkxgXp
QMVCx+cCWduOLU2SIrNHWUHIaIKB5ZJ76TNC42kKN0UaH3AzqApKgjFvszJs
elGISj4uWOjdyJjiazS8hZhuXWme4bRcCpbRFlLcuAMnXIr2fy3xwhzrhTGi
c8q2ZCdEA8wPZiJKPiDZTZXxrd65PkRqjPYvlTpE0yGhbj6UACK8WwLT4KL3
oYFclWVsh+TgSUz8bj4ypgD4Z8ewheZ5oQ9whfXkKgouJt/Of/WjWE0ll3re
zCiaeDqt7DS3WKiSzbPVaNFQdAMyxmEfn7v3UF/QN7o2jlvEigvA5jBQIuis
wcEusXJcqHJ9OVCOa/DxKkiD6RTVqzjPONT9sK42dEydtJHnodBaLnQyvax/
U/fFMQ5oBd+4AScbedjNinhfpJkBdAqcJcnOpUyBIFYf1qJRZC08Q0PxGpYm
/d2tIF1Zgrg8rjOFtXJf1CBtXmAfgvDl7OBX6jTq21LJId1PSRsmtXAo3rdP
2VIralU7FUfZMQjBr6plNtwXAOTEoNiX5qUpngF5fkLdsTZZkT7pTPbf+A6u
3khlut1dh/xS6hQ4gUSWe/ywTKkiyp+snh0mEWoP4D8sdJSVcBC7NEVE/3pw
qGrrINoNLOUH4wWD0YS5pWL82+b0aruKcFa4Pyif8YRzqTeB/nyIHSVsnl36
XZPVF1sArA/4G201V81WLWiPph4G7n/T3/How9KTxGvTFcs0TfQ+VPfb7GW9
dD5C7YzHpDYkKjcT4Sen0SP32c0tDyaJJPijNMJ0tVY3pRRc25jc/T+3mTIC
Tk0sC4b+qHOcaf6VXrIXdG2BL+K9rARqhMTw0bywPnJ//6gQHskCMq1oReIO
IemHjanMNeNsBgDyCKmnHsppefQE2bzqyS+ys60n06y8TFfvL41d0jPbfoHQ
x2GQ/mDpiC2nA8pC0xBDx494MMPQCrjlJFpe1U8BAD7yv8Bx+TNBMBEDkVxU
l2gT0jfOGrKpIiKRsrL4hMDRLGH5URLIgWndPml0i6Hz08Eq5bWGNPlLLIwd
hdew8TIo8/GHHguuxDud4R6qCoTcyESjQ04ZJRwMrWOf9Zf2+OS9fMw5N7ED
oYiQZqBKmzkE07AXY7pONoy8jQJylp6NhtSwb23GyoPVnvQJv4IcTmHYzcR3
Z1A3et/E4gBiGgnU1cA4V/JPlGGsCK/MxbKEWLOlx/Qb+wu2nMWRHhzp0Hty
j6AbVdmPo9WGaDQl8BnBCP++qLxWHfpfW8vfGUElmEnGD7gsZissxuMAAsrq
fgiYxT6PZctMDxXwxrEixrAUOlcei10ZqdWICBzTy7Y0hj9+XdpjnQZI36Bm
rDPXsjzkSVv6YZHjfA0Upr/jdS62zYHwqpdtPxwSLvS5wMrNIy8hOkmc4Odt
AT23NVlBE0X/EQpVQtrqui9Bb8TBoXTIfQSqyyTUqHxPsxV7t5vqkSPFCwVl
BGM9pczQg2JYRWMIR1Qv8iUlNni1CN+SYJMCfvpVxRyVQl03xsbfXK4o4tbv
AhsCC6N88BOV9jU+bPxEA1KZcYVk8wUHO0hxqZ2p/iZoS6Zkf7kMXfoAUEg8
CVfZZrItJoy/OYGZA19MvKj4RvViObYvGBcPjYTf+gI0D61RkZ+TBtP468KP
uvJmPEheFpmha6HQTvO3yEWc82VKw0qUkUzaEJ/nZ1pHjLolOY94U2PYqS9W
yTpG5RVPg413obCrhtrAhgtJdbzjWqLb9YoinwqntNjHOj3Ry+qE62bxs182
H0mgI5WfIGgDJmy9Qs6gWPHnpCH2mDZwY/HhpDCRnVfWIXGXzy08CL4g7eGU
xL1WLzHZ693mRPyg3lCuBzaqodOik+cgZGH6SEqlAXu71D+UJ22tM4BNVeaU
zWnJjylOlwO0UTWbI7S8evOBjxDH0tNEJKQY4OUewMHBEqxlhJGNMPDhtjO7
gnjk/Hf+5g3Ny7GJoBDUreXWlekMAMokQZdDL+Bb8SXWTz9zgvhPLOkpT522
wkEfFqDswPiJbM5svyNITidh9oJNw1D/+xNNyVWR28ekNWBKVhwarDLitM6v
M1yxJNg6Rkm92+uJJNX9ZFA9lSj8l0ZiQj/74bbQ85wLPy1UVijtfzvO4+wL
pe2AXQ5AOO8isqzznjUXhuawP/HdeZH3mXXB7XyrQc4B4Wov2xlZO8XsZNb2
QIBBT7TXOQIS90YYKFZQxWY/EpzYcmer0RawG1krsDYyidVffMPHc/NRlGvI
sl+kucevgtEENyfXGvqmNObSCEW2BwlBo7sC+Tz4wVaugZ6n4bia2TTX4973
7zQYYFIoEJaEj2yUJQSUdpwHGFJHLA9n9rRRoTLyxjCDMuf2y7VQUUepEO7f
P+jtWWL/4vGfjTDeAoae8NtjYe347yvsDc/k3nUPf3zIS1SlI6Zy3LiI2VUa
SHh3yWy4SnBlBVKvfFZyE1YtFAleq6CZ0NyKdqz5lgw38/jqRQHEk5C/2h1C
ZRsQaKbD7wuVNLa0qYqOUVXcyd/azb9bDIQbhV6MrP6uUq92FlMGmcHFC/j5
SDzIsH95pOOPpetcT0IputJJOQykoXi8z6kE3PXht5JWkXAFmsyJSNJHfHFj
bXiDfRKwDvODZWX6MAiLP04WEiX00Egequ5P9GGuxrrUBYKLgY7VvOaz5iE+
wDFyjyOnbBdWzdDTnmiK3RMWTkrhEaImamaMitsK0LXR4D7RzZ6yvq6DKrQI
qpPaNZm1L6nPGl7/sGXT5/8akC7C8GHYVjee4/qToifKaOd2i+GnOt+iGPHl
esjr8dVyHNycJtTwNy99yAqwNO70scYVJJZT1DkRksti7+FxwYAOdSq0s4nN
OkI7AtqK+DC4o5qkSZCD6z6jQbNDN4w3LBJXlcmWpcV7Qv/ibq/uTKMlMeuH
KHPsOZNYLElQ9JEOaArWjElGHpWLHXLlFwPyADlftt2OCuKfYOvlGGAFam/U
2ULAfO8auiTFc9wT2SrUYOkOjQHWSRBh5CVjGgvzloXe/Q4++eYSO7xCP4Pt
eXtOo9kSE2JXaRx0Id5Kr9hd6UCoKdYSaFIYck6cEhke0Os1bwEmrLBYx1IH
ZiiniycLWuZtgU9uRu38jzBvPnezceCLVaaVwfuj2Isd2QQLHxySgL1WwCR6
4A+uu9o3umqC9rSZHryIRH6TGSu+Nr1QhnDv0A1cWrswlwnkqcCjBELcATLo
gaUKLF4fVYm0HrsSobreYrJFYv5YPhqQp7flypXdEsWUwe2HcqEM0bXm57tn
sPwowjS02/SCoDLUJEJvGctBiHGA4sdZ2tXMPPTcKBYLonu6B/lkEi6TFnlw
LLqj4dmOwpAhti9DMkGInaby4/8O5CbaUCyiDJUGp/KiVvhTBNkm1OuGkSlF
e5sXO39zyEozFtHJK9OnormWuum0gPbPeK0f7peElRwD6d1zOzR+Xsldpfaf
zRJLDowbcYZDen5oimPKYVL1JcXujrbbWWstfPORX4NTbbTadL1T0xxfNtaL
WV8NXqfEW3j8yyA+iBh8VYiYh/6h3HtEHsdYsSATFhTwjZS3JEuN28Wb12dF
gOMHri7I/EOktHKLYgWuvWpZdXrzpBbLJTqgtehbdKvERo1+JDbCABHb12h3
CcVzvi4Njmo/v6uEBU5XW7I+mk61dSuWwTAJBzDvr1kiCdmfI1JBNweoBi6d
Qir+kpnS6xdfpQnt2KazqSVW0lfLicKRpzGRHQ2R04OT722m9LtRkyz3Hpqu
lTdfHLBrlnNLeTCgoh2kS4SQPwFaHJNvxZRmjzK6YK3K77G11mWaGsx7qLEb
9RXnimnlZKfc5mci86Yjj10f60vwUClZ59cXHdbE90y3p99902pVv2EJmQ24
f4MnXMcsgP+JDMN4vDuyGoHGjnl/WJXKPGofno0r7va6fny/uIa/NQoyx4pz
79b1W+lr2uzJ4BzHPjy6POqe3gwKzb+41TyPrUwNsRo5ADOX9m6NP/4cRXpN
TR1CieK3UXykBxAMWySPZeRjKFDya6ZbYws53rnnbDMUabc8Fh4YvAb5Aztv
3SfjqNMwI3dgmVDbM1aAOkuTGm8nG/iCGq2fWJoOJwc/IeuB5oLE/0edXq9P
Fhq3FmKD7QY0ogkjZkfbIfyaH23WFQaj2HdPTMh51Hx7K02oZF7iAkeswvmL
n6n4n5WEu2OJME2n8/SOgCuYTVPR/upZa7GwU2C/C6fOT8RCVL42x0Qc/CDH
udu9AnzUIJPUx6EadBS/eXt34qU2uE46vpMc8ZWuQuFJNHJUagXcUDLfUXRc
I75+eretWSBD5sl02DtY/bHbQuATXyPsSmIO/kUYjBshmfZgHzAQRi+dZWJX
cmBdyYbyTPw/DvUTGH4+d7Vlmz4aow94xTaEl/KJD8HITcqRZabWCOh8ysXZ
7Qd5z6DbjYaxPLF2aWBH3r/grJ6flwfwVydkQhV/ifArtQjcQgDPcc1KTLWL
GuCaUsRkHhSeIT/xIE/R2IK+LfrLlan5jJnSw8DmOQGDzfAUQ8fmrON9HHNf
DhS4eMNN4hWqT7FOry5/xQUX06f3bj03Ws4XDOj6Le2zGGDFyHqVBi2Uwjf7
ZyhKLwdU20hmG7g155Gkbuf8xMtpNyPp5tfsaBAvPZ85tP8h2UItNx9l+pqK
7CvFItNkMFG+8zl/2vSjcRLPqwUJrRj2/HDEMl+akjv7mhmDN8ObMuYERWXJ
dgT1jaPgcUlFLKHi0rMk6QXWm3gfu8AKtLNX3MTIaEzAyWI93ywd9KqFeKwn
lmMI/gQrja25dViBQ0oJ/96CfutDs12x+DpIW+DWlu5x0txMv/7RJ9DopBkP
Avh8uUGLUWCZVnkkGSpdV1cRw62SIMZGr3u/C2GTn91x0NkyO/uGzM3Js/Jt
2A5O8kqxd/YFmIBXjjo2j4y9lBllAmVoeyZejDdGciH5cT0cfc8IfSAJqGuy
1L6zgG49fjJf7Oc7WJcYhMYN0ve/EVK4vHnlj4wXrNHHNRzLXpVzz9SCXDip
+VXWZu8cnSO9StixOUo9crff2xrMmplz9VwxyqtmnShn7N9fNDUdYBKW+49d
yFjaXdBVZfg2ALN63a3sNWJ0SYc6/wGZY5yAOqbT+6z36JohQLDhFeF4e76S
rW/odppOgKcCpJg59g9AMBq9CNNDN3E7o4GFro1qhQJIhFa0ue7KQipHSoRU
zcuRnQ8Ir5bMGkoqp5Jvq0QjuPKQQ7MnE8NAIkPb2qy6BVdDG0BD9BuJDqSQ
GYnTaygmyvowqLRgyoOiDZuRQh3V+dy4aVwIybq5VDM1PPyxFVfdeW+60JGW
g6CwMCunsUtfXhjV8P7jIcoPVYtXO4nBTtWEqq/CWGikXWMM80iOetVi+6ep
gRDueP3UkzWwVInWkd8+TJ89TuN5BsKWSAMmIey131AmP5G29aNr3P0ToTS+
sw+iFs3efYiuD7w/Rqn31VazgEZxDxb68fjeziMkzH2YyAL92D9IC2WHDq5j
Ldf48xX/fBcLDmHQnqUQLgFnlpsAIph1CcUI4V5ObVbmrT7fFSDwv8bTLCGn
t7lfnHJ9fvCVnV9+Qhqt8bGXgx1TwpNNRgpniFN8U+awGN+Qa4yfra5HSIfh
cQLoG/knlQaUKvyCtMaY5mT4zfKr2qdq7zb+lC7hB7bSAkV+aDcUR0NhJ8wV
jxRrYlxzU4muiaH/cFLVPCZSnGrMKt0AS9pGShjlviZrpdQ5taBzqCFFT/hL
IIFrYsqqcT0XSJtNAxMhNMtVh2r+PFJgGtEsn9Utb/D8t9YaW4yvKWzI3ms6
3K9cVl7GXDsv0QnrLFDonYMlbI/Khyx4etCazSY+e2WhhPMTik1+d04mFAsw
ds/DFNTmLioJCZRE1jb9tnBN7RRfld9u4frncYkDX6exAs46F+27xUJcQR5u
RM6aCmF6Z1lUBbFrjWQqwvAPWx2mawuxfa5SXekHO5qOo9Zr3NkWpDvAIUZf
ZtYGuzaToERcFwalKIEFP9mSi+qksTKpq8kKE4yrzkII6HRcfud/ItqjrChh
pkizGGgqg4tWylkafDxvYq9uTmhUENnDF4AZWyKC6SvANFxWq2sY2NaJkLcK
O4TXCK8ahQ1BjIzPI6HmKY7cvc0aEUwW865YlMOjixXZWjuivLWJ9U0IFIpO
9qiQ8KUC5fuoCsAtC96j2oJmrpVHqJt4Oy4PeFtDCT9cHUb/AoTwYURGtLbr
SJBFkp+RlLh3/MsRXLh7TbLXznHA+5iEUB2QDfMEr5ceY/38LFcsqq9ykCYv
eDgA+tNNCVUAcsfHpxUtukW8KwN2lO2N8yJu1CsU5qN0v9QrcWkQq//Q0B2k
RGkei0N5vvl7YK8xxqjpzZQdSE6Y1nc8wdG6QbO2XigeDudD1leH7RBlKSDr
bqIRUVAwBMxX8Ooha2SOFpKaQvSI84Au2ItwOs4Tbgl83TMGHX+AO8iqXdiJ
46Qh+vJLEoMacbw5X6adLVbzXGCaiMAaVTHIww25xgpQvQpG/HekA6g3iUJQ
ihKmOki9lQR1DIu+qhEM6XZCqPi3Jv2gTObM9WqiObbLORQdyZ/EoyjeT9ew
5kOlO/fUf0fd4ZHB9QoT9jT5xfRf3/s7Qc7nqVI9rVuzsD4tvlajdJBfcdk2
WN7q+CWja0UcygErmh/Tg2xC6PVT4rd7XfC+070wbYE6gY/r5UEQt8AY8diL
ATWwGVyDzO68HduQwq4FWE3qe9OsnFvgkwIUbGI6DCCxI3L1e2Ycu7VQ/Ky8
T4Pszp8y2vDCzbnJrD+aR7PVdofjrpVuU41NAGxUjd0iMsGtbB9XkhHgQMql
S5o5043DsYzGLQpol7ifCcHXRc/Dk4q3eiidcbh9DZQ+HXL95ng1RQ9bbevM
VYkEnpBnuP2j4FVuzIEi2PDIAofAGOx90JYHbUvPW8i2fHuWNnc8hTPxCePq
fKEwazNGgMe8SA2GGqUgMdJDTWG6Ga0H+A6srZucaJajUjqDvif84MlQTiAp
kQFKO69hfAxiS7Rl8bCHsCqtrdrRDbCUqp/4jLYEXfeiACQdZd8l4lESW0jc
aKeKpgXfWDNTdHyFT17DYDc7w90iivcCxhINFSgN6RGCE8dyOL5yK9ori1YI
6Ki6p7sj1wgD3YQtzWf5ugOcGJ9z2FUfFMRxmqyV4lp6RpqzrMgxBV+pWXex
z5BnVYQSnWgFu9OxQ7PxCbVGqPChWkXDCXMnGlL7etyFHQrgEIN/N/tosZPU
tQ4e3tHn9QqWDb/yURdfXJJ5W5bGXByI2IjwUNlwJjBEi6pwNar/dQxwGf+S
ygrRrI3XueFSPYIYvBMzjOnUTW40mYcTTXRzD6v9Wd+jLg+xn0n9QD67n0Cc
S+UYetMtflbcvX/jRAJ0kHvlq/iQRTzggqxa8VmaN718FbHBFjBMF6b7rw9n
F2AG6BcNNAXtJF65JqR/IsGU7qEiz6hUpovDtoAt/XqF5A1IRqp2yUv8zMeJ
ItA1TeYnJkSJUJ0XC7nfYntJPJViFyNcQ69avAuz9JnwNAKPqFB9XgA//iDy
jauBb9RpO+YN+n1rQqar/NkluwYpomoGS7D5u9qhtAYMS30Kw23llvw4OVPv
XtqsXIu83BNjE0QZBLxuyG0+zn/bDii8kXMQRrYodXxXLzxD/8m8Rjfo5XJE
o/c125WfBto9gy3U074zQ6FmKCj/m/mz6Rq3+fPy/aBW1yaCoP7ngY8aEYDN
rlgYhpR0O3D9EALg57Bk2R6H0knLYmNdG37mL//WYSbuCtrqxSTvaf6IhuNm
xM2x+zv8IF4dM2swlWeCap7yNpC3I/imVqSajc2KYppEzZWUfbm0RgORpWFm
I1byRKP4wU/+Rg413vwIdZmFY5oQHCtUxCnS66rEu+QzKUEHjHEZ0erR3UL4
m+ZlAFJY8SifNBBXH1y6SVn3SL1KNySmFqe81YGFejUuG7wI9Hqqj4ZOFH1M
+xmFOfiuIW5ac+QMOTL8e+oHOo+l1t4uretPxicw7HGTIhVAeCvM4tPVG1am
FT/dGq5ugs5vwPJNVtxp+vrH7Zk+pN/c4rMJCCUAD3rDC1ka7D+wVF7o9+wn
s1NPDnN4u4nLQg0AzW309XBoqNIjCbENdHt/yMIv5fcQG85KnL/6ZSu1ehNw
dT6FTbX/4z/cIkUVlsUH+YPaY4SAYx5RsEK+7zpoYDZc2aKSM8wsrpVzQ+mI
95AztHGLL/nk8ZbsKJMved3TElG1iJgJHEIOpqRhO0iTjUwZN02b7EoLy5lt
LeySshtXoqrh0k+H2Zk0DeUYzx6Bf+CkZjhczOe7bSb+ULsacsMcRswvDg9G
LyjMNc36BNL4dTp0ejqd4v7kdLjv5yEGwH/pabkBF2JMZmMhzNowjSJITNBb
f7/xmyCDLJqBkY8wpcFieVAtb5DYLc0wXQmQ6aoXnfzE3BuVxgL99/cFFXJY
RoBAqv9L26/nWI8LUBT6XkTKVysCLgIbTRkiIYgvuoenVffx2Wf/W/QOiksg
SMHFX8TAFknttfA/Qm7wlmOFtoHOoxb9MDMIMooe7qja2u25j/NcsgFWDj/F
xTwTTlRYHjzwi6RWE3ZaiP6xI0NpClM+wjQiN0FESrhPx3GfqNipMw80UHBz
kHQe+VJoSgxMardcZ8Th2/YDlVGKdqFcHFFeJaAleBBmZKpT5dJjnjBA2OUf
IIgUAkvOSYXMIlgVDK1uTZRpcUnh39vl21cfZUGZcmFqegW1Xw1Vw7jqwWs5
PxtMd2aFlGaSSE5TkCdzTNkxrdItdDiZwCd5pYOJJiUewRoS8BvG/wpz2bEa
jWt6+xrrjHSJfPKdWcyy4KXrlWSNIcyDPEiKPZLKTcJ9CM6DZIs2Dz3Q5yQS
p0Oa9rdxUC/kuE9FDK7Z5S2rpaRadHTJu2829SaTmPoj4MrTl2vwQ4fVRPPu
BYEjgaXmGQut+AKafWT9hwYd7h7s3wmJcN1OxvbuBnie2eKPkqtSlFkIQpQg
8A9RJokEtHWTZS38Iw0NxBE0CaC643q+9xDNv5+8VqbhritXbpyqydvA7soc
ZJCu0A0wvTZcAZXrqDh5CublraIAVJIMqz9YQHSqstX6GT6QrEa86jdMNe89
CgiQksD5C1jTgsqESQrSL/RU9E11D3zs1omiyDV80IDF/kLUay90D+147c6L
zQGSlyp+hte8mUl3w+sMtXZqG3yG2NtKYmHvDeDkn9VAXNwXrg1MqRw4SEpE
qnP1UBKzMjMkgFvTohJHQbNZS97ZE9+EwqI0jYOtbOu+vzmcWhtFf68F40/a
X004j4OicokfENSGYnr/tAPf3Z4jpvkske6m5vUrg+//mhYCBkEKUqRu/IgJ
1MI2jmAu/pioq7ioLgX8XRxbvDZik2MsiK4XpFb7wPwj6Af1hBlFCmuriIup
2UeqdFiGhHX6O+xSFL+HqAKEm7QeZVMIed5ZMttQHkrayYXQ5AR+QodEhD46
wBUBfjppvKf2M07asnuN4o4wR2oSsI2P5JXhC0/SXUpc1KCsSw1ADvol7sEA
OzaR+QRsneSzYVKFZmOVE64U58H+o7lXD1cR0IyUHx2wxquFGYRUKz2umoXe
S6NIIQPKBb1JRf002Fc3QlDzCmNSv5RGLVIs62l8NYML8itG6U0+NMfqg3hS
acVgXAGcM3BfHcg28n3n478B6eUwE8KpCaZPEb31fGr4mohn3QAk4jreBYyb
opotVi1h1l+O3Cq1+fuzXIzIG8OK6LnF4zR8VEvxi6SwdT/62zK3fLWH/1II
cepI80RF0H2JTNiwCmS+qBPnMA1HzKUrXcr81Y5lE01QJjxlmMy1odiprsdH
6yX0gGAPe/Mh3ZYh6F9va0Mh6yqf+YE2+dDqUBPiVAqXsMWkBqOtBmm9GzhG
sgJhRfyt3GYo0jHxu+7rsgKvIaOOMeP/v+ev/DmnSt/ZPDblGKdQqv+hEbqo
3W70mXB07x/AVhLIIcN0b3TxOUsi4L3ndx7lLxHglwajlJOH/R/6XyqM130i
TCY11pkxdNwqXtdlj3EL8F9hcm0j3wLh1mo5Qqzd5bTKI9DLMkeR+1OsDo+4
nkNGv59MDFv1htNGIlw5U3M01pchIV4ckMLV0dmYk1M3Gb2WMko79xcNW73l
wmT0CIoOwFWpxCnu9vtni9rAlHcR3NZrFPvDOhK7doMAn+WfpNokaHlq7YUw
N0caWTyXpsjWdLV7VR3r+AcYxqzhFbY7syAxg3JmPBsYqPbOg0UlYfNdk/bS
OSvZa9StObtqkuiUjtBPwK5gHOF9+NvlKQ6NiEpDg0Kaxc4XgeNOxGSnSieR
L2TlN5+h+gbM0jVqt7/RhtvooVh8Rezmu4GCCGLS/VzoL6/w6+AtMn9KbUiM
NILcgo1OQEv6ugsmkUdgBNydnLvCCOohpMBv2fvmBmYAc2EDSQqK0BxEqEAr
P5AHgADFLTnA6mn/x8Wpzpwit8aL9a1axnXrFrkmxjre9aWKuPcXVrSoFuwX
EUlGzcZ9LV3u+58dh1XnjwvmjFpwveCk9Zdfwkh950Iq/op3FickARrc7KHl
3EQwtoTcSWgfSWhy3J4b5EUel6GpPyt9YxmgHlToNDcKms3q/1MHqNFjnqY6
xKu1rkAT46ZFCMt0+tztggyEcUc3q3hRJ7kGgqd4XovklOCQOP+D9413uHzG
GJVXbSFHtdprfgCgDT/Vr1wMLcMHYRnLLhSXFVlbZgM0YUrDZ1jsXuwqu0sX
r5CWqUcTpyEs7jcTWv74HvLwioVQRjBb3HVA8xJTWofqd0cfaJ8wP+SzAYH0
fhXclPuzxl7LQ4qeCjrrjT5fRkDqLGfDjFKlFexCAdt+qC9xJYzdRa4AmLrl
yNoxXSBuB6NVKOdONgo2JmfHC3AusbTTRidKwing9+QHNoB8sKMREEOMSCTi
7QTAIFAFH9jEOOt5VWAgy+MI/KzTSIJ2Eun8/lUbRtR6l+LVVsakj0dcjGfX
EWRnkzh3xNEo87VaIitQYttAheyABSwzhlcVP/5kAQXW/SKMTHs50Am9BQkT
2UsMtLaL52sYGQWMx3G7TX0XMALAu7AE2Gi3EZryKmAW+bqQl0ot4R+D1KYG
szoAGtxP5XqzaBkN/nTUuazi3dkNBJs+ifANsytAPaJVGwb9rvAVj2NEZe8/
qnMTF2iXq/TnKphKhpacrZh3SWZGL55dpnwEni5Xy3KldXZHIOiZSGVyhc3w
RcO94rTcWotFrqpUmHiqkAkHdE25CVoLB2TN6N4gX6qKsCEJ2cEFE4h0GvJU
wgiZy5XIK8I/KdhgwOKybIyFdLv5THHbja3cIbpdO6y2k97kotedNtYQ5GVh
5/fMM59SNtoberMaopuluK+HmDb8hiejlgv4raX+KuaNMIXMKPakfzQjC02I
5iLhUgzJwkFFGJ1yvW++XqxJGLFgBfdo0HxU3BgxPyqJI1ZdeZnPeRZiR9W2
hmsUQbhcgIwFKd30Fc07xWnFoopnaRkXcaaCz80PJ6TOkdJUIJr5hYVJkGmt
kEadIEoWaqKOUPmyyxci6CTDd0xhIbk2vve+yzuU8SnrwysFw7aV2xSXq/EZ
H/KdaZZmuk8KDzS8/VTB7ilnc2wtJFxshT/sb2tDPULm4mTULTkLP8HcSChJ
r7hGHL72oacE93od/u74ZgoX74pGQUGGkGk3KkjOkCLb9j8P1i7dwxhjZyhH
DcEEmmL/j0UiS7FFEh1To6IChwFJ4HoYUpLtPSh+dug5Eoy4xK5RYBpWplHZ
dHyGC2GvDsMmbgBYZwtMcawouVzNWkFv/tfXfDiGm9AUw+CzOp+qbarGo7fN
RCtcIrCYN7Sofw23oIss/e9wVkmhOEvrrkS/Zb4x9yGL5YsOMbuDMJARU6ih
QB04JlnGAdR3BekQMEV83Rn2ufVIvhy+Ft6tVXpKsZZFJez5S7Iei6JTrHIe
zMpR8ulOW70/jLOqYJ23S95t2dXFEMR4lU2xmAAh//HkNAdHvtWDnW5DMBGF
ZL2llCLf/G7i5EJPs35FqRTP9PFZUIcgM6cqjMZWtNuKsuBWvSGSeM7HhVk/
Ml86/Ak92sTsWxeBPfyqaEh5pbMBZGjG/KRiXSk9x9aMO50jx3TGZOXifUEx
uuMgXos7WDYCzZOjqnB/Cc2DilrRvZ2rZwEIEd+lz2o7iGe9UZGGqtBcvyh+
ON+ShJTpU+eSE2SccR7f7TQxf2XBctcieGo5wHcDgcC20XdO2OQvwav/jV0o
PZkYiKSWEz8iAvTa/5FRfXwk6jPww6Go3pnkzzv+2JadpPtMIW1WrH+n/eCN
9zH7UpC/EuZJZJK05jlqK4cfecLPi27z4bDA7E1grx2HobhP5m/z8El56oL4
sSLR+xqg5fT1u1OIfMEMfqYg89gi38blHwQmbUPBrYOLnGT9Iq3UtpLQp0GV
UheDqpLa5yxdqV3FPRnIbjHHXKMeKhVl6sEYfYEiOp69vpjex2tW/JBS/o6V
ni5OUdFWo6IoSWYTnDzm664899GEhGUbTExeCvxvMHvul2p8k1ZmkzIPVojF
uRgODAO9fHcEbhd5aKJxCz8BFbiBRU0t9ZlZfjMzvRLaW3BnuFYC3oo1ne13
37Hcsy/fWN3wmlYEJYYuuLDBlrzRx95l8K46uzJZ+58fM6HGG3msly9sm2j2
YrM/AwqunjHpesRpY6VWCUJzA4cW3JzYdjsuXuC1b4vbJdOPCqjeFAB0qgTy
XckobDMyk/cpGTom6DewzjSx2/84xFNkI42R2gfzk1r0WFzpWx2Osm8iAHW3
Vm23YLFPDlp+Z5tJzqkZSX/14aje8VNl23Ts+WEXiBiCQYwokUDAz8OnNbqR
OEMq8Unin17TP4Y22qMNSfTGWfXPmK03a6LWZ1jPOGHWYeokgpQ2cHBUaPSB
vW+RiRW9v3hxCnFrgKmvjWrcYqG09KQPu6HqxeSxH39GBN74vU3bqQ17DuPJ
1x33R0lSpSUuuWFcc+exM7T/dXqazZH54P11xm3EmIa1TQ5RPN3qzK7AwERK
Qvy0QsTVwLv+ELYF/8phEhi/PN/CLUOsq2B/xljmviysCf4YIs1uHzIz0Uk9
yyf+pB74/ktoecbULT4afGOUm3kSlCU5/q8ekGRgS8pQAr8HHtvOTBk9Au+3
892KdLeD12Ke5l1WqQUGWr8Q7bYGux4E38m8AMaqw2rx3fs5QNHXhkITOrG9
fE9goUzCI/NMOhPIjI61HSDdWJSWhfnnkPHuoolds1k3RJfLNFCD4Di6NICw
9rkRF3SfVPq+FkQDQKo3P43A3qZn/IunWUQ0pyNLHHikAVWPfTydEZxlDd+P
6IIKfxYAt+04AvwTCIiB/RWJutfVj3saDJVwMXyo1Wj8xx3u/bultMhqVhTO
lTyn60cvndj6Bd7KmBzrrSmytGZHwF3o5+eJ2HaT5b7H9F19TCfsNDnJqLyc
Hm5Rs4zDHObV8vvyYfcHBY/eBp//Z4YK/dMid1uujb2iiRAiPif0NqrXbvB3
sZbQvB/ERPGx7iKDeYrcDjSwl6G3RnGkh5pJwyg8O3ZqogEH/qIASl/sY3gB
/yHiCf8DXPntnGT0Ba8p7jpvYJMsjRyA/6b4He9P0cG4DpYzhM7vcWBQ+kk5
tint1acHEAh0YAPLSWumVy0/TPTg6ibic5wm+CEVJDfvHNeiIcoFl2cQBGnV
ujfPjyhSV2NBYlFw5MzPNnCJAJHiCFbXPbpboLUdeK9SOIZ/MDbZsqvk31Zb
DAhX/TvsPfJIuE7X5HB2sgeQx7hvxCt+m2YWEU/zq1gjT+Dm9Ecisa8cetmX
oSwD728371xJrQN+kgExCw7rYWlNrEjwybLbSAw8qUkBwMCCC80MSQf9Qw8H
k2XLhREaBqF0xMcafh6ZtTuMPqY58CDYqRb4ekP+Eoc8uYib5g0dnyyokf8P
O+K0gVJOoAHa2FkfvULCeBB7IK1YwwpqR7DIpmNsHbJ23MkkVguTnHwvT1kJ
n/myZCZNP2C4noExCSaHo0szv9HW+wks8QRnK6Ww5VjPdExsx5PQXqoJ2w8u
o6Oy0LAwSmE3anO6BWQN/YYQ9DsY0iwBIH4Hze/aTdJTRNYsSrDgg9rnWXWV
aOEBgvjcZOcn/JvpiigPPoAaxPro6R+TCBe3CJRo8UM417a59rBW1ODykoxP
tSfehRLpLOwSz7qh882QObCK4auaZaRtEu2sILzvlyN7zivK7GDy1POb+jxV
mTuyipgGdzWbYCGJNT3exH/PwS59zG+ejY7EAW5r0cwz3IPeVKW+QaIAIiej
Rzr+UgBW1GSFwRFhC1Dw4575Mwm7iNq/mSu/oo8e4wbD1eiQbn/iQh4b7Lqk
CX1OyZ/A6vSwHSkqUTtzUSdUAFnb9o12Ifn36Gz1i0lSuTJi4B21b2VGzJtp
BwUnzb7CAuokAbDwHH6tdFLA1Xderf8hujcw6kNyjdDV3qUpPvLrHqCtI+Ar
h+TmOW14tqAhJ2aKb0MhEpjjSlB9HsbuGpnMaXIjD1Nl+K3VQw8oAmIL/EB9
DQT+p8nLlln0CAppc79IB7jzIc8SO1/gw/itkRwF8ckgKMjEUkTlN5oVwsIh
N0ddsmiv0Ah+tXJVcRms7wZwOxWRDlVKOG7TTzYucdDDtbOF4iKgHWkJvX/0
Rlg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpeg27jjeVdZzqbjln0cl6c2nO3cwbFXBaz+q/OT9RgQKS2i+J8J9uRwqM24bvOrnnC9oiVIekdYdVLk/1TV2TAoAH4RxkSQoYYjvOyFgpmu2i+4gcC6t8l4SR3ExWnyAZ2htKLNJWepPLgE1zMiKbDGi8I4Whul7nMvAE0XjwgrzGaUlXaPes7EvZhGkIOJfviKKvZ4UWzle3MtuStqyLrey36DzKaROW6mHzoYkwhuXYczipM0VcOvEH/Ggg4zid42Tv8r/HJ2UXoiAalKJ8aIZAJR0Yo2+2ntS1cyG4nyvQV1R/9tMqHhvPzsKe8pvOV7i702rvBMCdN1mM1BUUwHPA/EvZwl0woBT2ef2DKMxLnEUTYgaXAjeNe4GHQkkEg8pZSqPC4RakQH6+Qb7BUjmKQiGXVS8fc3Z4jTb/u3xgnWWxWSZS8rYGZPhz1JzN995DdjDm6mMMyiZpuTw/jZj9eAtq9vVIOV0/yZFgppcUvhlH9vS8agzkvqk1AC2jTmvVHBH7gC77Wiaiw9T3NbkHHum7TZrIP3mrwnqTbqjAC1Dc43Ov1JlYwksVyIHqoFDOKLkJyVJci+QDdMs8Af1XvbPUXkxacWhjNaQZ45whrxNclgd5e92cfg2THjzo1YdY8Z0u7rOWU2eBfhkl43/JIuyp6jbQ9vtpsVDjvpb/HtxOgGZbssVx5grtFHOyLa7P0N7TC+7UVAXtY+uRqACMiHcsmYIRE6ZB0tiXLgR2dqFk5B96jWKiTa1Y0yZeOeYko2SbtCoX+F3LlXCDCjX"
`endif