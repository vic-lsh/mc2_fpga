// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kpqcpn7NUJytP+4PuHZewL9+2X/lYL3lsgnb/6mVKe6eFlGnf73KBP31OkWC
NxZ0UhDJAzrnNhykyDmUixhEELN+o3P0GCTLbjxI1plU9INH4M42ecHm9ogk
NTJyDxLCFipLiWyztmo25m5RQdTIo9Rc7t1PtxOYpqqECLSHDv0MS0i1QAd3
IrrK6aqG0QwDlRi8O974Ko3q7qBrYY49H3UYUT+CkOmHNBrALoZiDDQ9dHwk
SH3VvW78B7/YFUKzn7E3nu5dNCen1BqKJTPIJxkAzRk7ePPz9/gPiWe0zKs6
zXu4HwwUZALqAE/BA0NgGg7phI6bEzXhHO13ou7lzg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Rk9lHZIM7mm1p0ciuQRRAzAT+Gw1hP3ZH+WOKxqmBcMVe+l83mAeXiVhTUMB
q3kMkyRvvZQBvFFNIMwTkS8aUUmQmkxHo3bqwnf0zbcqkZWSYJDenZzeunmA
fGrfDZCSaaeTfcgqBZm0Bvgn77vYcXVXc0W/U9ydtiqPFeyPdotEJn0EHQhs
0yifRUeeaOh0V7d6VfMk0YMIOGrJNvvdc6EcVChvfxtaecprKut+DGYkfYz5
9Yfsat5cQecYGEJW9L2PjFrqY2iqoZsaTbtx+qfFYB7/9cvQl8CpPWkgC7yP
0ELP7ouJNAqRifbFwCfGb8+LfIIRS1AM5Qx8YtqdoA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DIpccT/UV52lpc659a2I5wLI/LJJfckzKRRPoCOnp9kVylApbSlqF99Lsmxo
oHi74VPy+t+VI35HRr8/nNuNV6YwMyQBna0lScesoElGYp/WZ7qI1Pv27OI2
wFN6+Il8j4h9cDabf33IWeAmGdJeD8+XOZTmhy9zeFk907vwgIgMVnYVRbH0
a5vVeNYdO2bxZEGcmdbTUqi5VGoi0OGVGPkt1O3D4d/cebGeXhZ46nHC2cg/
0peGGUezLm2u1kW76UjC/t3e2tsJ/yOI+PZxmCkKLKlLt3K+3L9ziqjUAekd
coO7iFHGYJje/vMfHxkRd2sMzZuTirn6YZwVlxpzxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d6DRB34VvPGcLCQ7nnJXzkNsoZpXSpL7JohZxtK26okhyQWPNEjiCFDj1ryz
08BQ/KhRSVYOL/+z2fYxRZim5DzEJwpF163WOXnVbuwyW1F3Vtvmke2yPPpc
4c3f+oAMSbEl5URdHaIvbI2jXpUQW2OOUmVxAmEwxOY4yQG7hK98MzO20pIz
h0m932rR4k2p7UbtlW/Et6kYf7iah/nqD5DM1pEnZd0CPYW5sjhRs0fiN4ZJ
/TCjTUVWg/1MhhwfexwEAwAPMrSJ5sAu5P4/LvCQuUIgCmjH+fWU84dBcnLP
d515msjxM+YYlM8Mvkw0+emlOG/rbeSkaDxUVN8k+w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q23GoY8GF3LhXI/OreP3LVt43i9iivvtw+yG9mlO6mRExDG5i8twsm7kW/Xc
LmkhteMMuVi3kZr3Kty8hmrVxIfoyDLlroGikmQJ2vpEVYpMxItkVMqAaSC/
fg8vzTjec28rFPV9qXpOL1pnd+mooZTmm/S/LOhsfOGDpLj3utQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XBzO8nKtHv4W9W2xEDBUSGV4Ayt6bLkPHMWxtQJK09OTl9M3tkMqFJKBxtj8
5M7Qnmd5C+wbL8Y1+Chjf7TCUvwUWkoIwik3Btx1npSpJg8mDsskSGXK5iDe
OwJbcxFfEmiXsHN7cmfJZ2VQTLUlf70LOjiA0FBSOP+4KQxkdqBzq7uY1MMH
hqRce9YRpA0kSeYZXwplLuVX2eIQrRxG8f8Vdwd29U5WDlah/RdAtY3RhSFT
KRQov5gknM5d/MErpjUAuPTSukGqii1SLrXCeISOFEekVkA06VW6+gJd23qW
7zTAX7cdtDx3C+CASvxZOwjBaEATWMbib1lVVkAqsVjX0ze98BhMGtMosXCg
OeIRhLHoI9gwmrUKyHtleapGj8+7WkMCfSIcllBz0KPlmTsqVyzFz9VDabLb
AFBfTq+FcnqNVDVmxJ1j/C1hNh8N57OpJ0h3QduuHa0dRaMxZbLeyIlqKDtV
CPcBZyXW4E/3RlqVR2n6nknzlU5v1Hek


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m2EK0YudZPEUH9MmohxGxO8TU8C3KKE1YfSPBz8W1RaGfgBuC28GNYJZ5YFz
Unsiv/86hxG+lFdUtjOEgxpwJtM40KLkZVMNECGFAmHtHQCiwoIzAmF/6rY6
DA/c6IhwesHr/VK26fHnPLGgFMkilTDqq1wE8G5UczU6srbaJMA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OMQZjYcK1X2aO5n3JC6n8N4ZqKpAgTws6lTHK8yFwclL58yD4mMbNm27NbqF
7nCwy9AhQm9cFUYWtaIsbnJNncB1BYsp7oesxUIqyVtnyu5+xj26eoaK8pdc
MHFdIe/sGQyugReb2aLwA5SNeWtp1VuGFZl+McrV0tv1VxeIkR8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 623920)
`pragma protect data_block
a2E8uXu+9tPi0ER+HAIAyTMfKxLxQLqzwimJw48l7CcV75HnZLjR+xv/0trJ
hcaY7ZzFcEDVZhhrbo5Lq3qI22hJ8Gn3XLv8R8IqpBobx5oZKjLeUzmBQdiK
KZHPrKqr2kEegK1VuUiLHvN8x3N1cCGgQm4/ajcuKIyvaMPKSa10rtjyzTel
7imJcfK3Qxk3BRqdD9yn18LRwjlJAAPtskECD1GVMyOwyfw3d/Ew+4G5GL2p
XfJ/upkFGOYzPb1oGv4QwXSr0OfjnDAzt+vLIAdi8VFebOOYfF1tt+mA+KhK
vxicPOF4liBtzmeunmPXr8ZGDItCkPKJqN56qcv/cK7Ue0qYkY36RuTSgB+T
SggEAzldXJq8/tOFChyVh6RFzxWP2bxHa/YCvdPoAHLzeMm34dmujUChMCY9
GQZFWAn9ALO5LUal5vlzbt6QxfFQtVzUHbkZE8oboHm/eU/uju9VqAB67X1A
xy6sm8cXY3n1CNPaQwAAa+0FUijQ/0hbZrEtZGtxyjzBgOJoDKxB0+i30Xb4
9rsLWiPguD5yJLFptj6D09ZYYNhktx3LDyV15zmz3Qfh0V9NnTNOk5qBcH+W
B7TKc/ek4Y9ZnpuGIs8zg99sacUYwq9e+EgI0+QDVtIgP2OqrLA54Uez9d6Z
Ov68DYshmpVSeogiV3mQTBlwGB4Eo8I10PWZr8Paj+AsziADYP9Lyqfg09ck
gH/eYDqiLYFiQqbfQt91T7WnXafwIhIxm7wtobMVZWKE1g5NZu6NUsHwF9Ux
0dyW8Qp8MOOqnNPcmx9qwinYmX7CpG7JLpyZowjKEq/gbk+iHGuT2oyb3x2c
O5H5PzMhV0GDtNG0hWZRUvet8VptLcibYVGwahkY9lWqwEVQaZvtlbM+pdIB
mbYSP8XJ7AkpxdPaQ+BaJGnHzdm8Iig5pn5LmlCsOYaA0/32WHCTaWiMNwnV
o6tcpXvZnHEWdXc9aV3gFj4S3ZpTT7abUoWfXss3ePKQ0LgjB2SBay3JGgSv
gEEdAoHfyGTUxQaa2j+Cn9+JnbYHPxqLe9iRZfwaeG9nGfzicv56GZFZmxOh
C/EbpA0hiG9xmape4xEPN++zXJa+Bz2KfDVxwbDurkeOSNT18fvZHgwUuT8r
qlBDTQTgddtGC8/exrUilBYc2g8Q6WJ4qaSeTvBFhPSfP99K0/LKVXwLoOos
JSnQfKcYyiZDR5dp75a6ecUs+5YMuGmHvlD09whA6h6FfQ+VSMG181ScI5L6
e4L+nwoBPrVa4yBUG/lYCPJqU5ObqiqaTeFGEOmG8FkboTzx7Ho+GBVcm5ix
A1XQEs0OyEAXrqZKC5ZVB45UMkZr8Z1LsgInXfPaSQ0ImTmj2Uw9uU6cagL6
yKpVGO9tQMzmqDf4vDBY5pHTC3adPB8/cY3y2VGMC1BWHSbXppn2MXkbCONX
Pe6NDOTpt0ShcqZXFn1DYJ9C2igD/vd8g3tAnxRVxGUZEUSXRoH2UuWPMAFl
nWcSMGwAjYMo6iTO604fO6ghnQrwAs23dF8lLIxi5Lnvdjp21iN+bVO9+v8n
ACZ+c7atmO7HrieOAe1VFdyNAN1JCV7SAOFWgutwb3mgto9i66Qqe/Sm9mzf
M/BdkBiEH5dth6lmu4w89e+bW4AYiFcRnR7AYc8yiC170VzR24HjT0MA4gjr
5xX+8fvgl/hLpXJqvKrnPzmGgQOvztuh+Li7fLAMJ8un8kwKKAy/2iVeasYm
Do2MGTbuEPR3dzJEtvhRTH0vToHqFcomyFAuIqT8EMTc/1ejOUJrsvxJBvHC
h7oMSs8VU/CZgmqA4MeU5B5yAY0BmEBCIYPFCrjWWVG+LFjH7DES0m5pdGRJ
QXXTtZFxZRDGgWk8l34lH9fb5VTvvcW0X/Ir3uU0zUujIKM2oB8dYMbysvxa
e3QuAMSGrEybPo1e5z4GZyN0b+/C2LHJ0/jl7ujpUdyAUMbawdmHn7E/FcrL
k1YH+keBrBas3N/CW7gmgyx5W8Ncd+MBN1WiKFpm+PQIsBzgahHk2Kk91kwF
Yg87lbkNh9HlJ6YKX6pTKsepLP8qoIt67xf4QzibKHydHwJ4Lr8rMKmrfGgZ
BIgHeB2d8uRJvQ+TuhKXCpCmm1RlSTJ/lUOaugXI/MzLRvHdXuR95hSW2aQZ
vjPvzNQGKC2FyEfH/oBdSp+WC7YPegKzwRnEHvkyDrxaP1/cLmBF/V6jFMUp
WX/HIrNaPedfLDK60J7XETKOdZ3NZ3yrfXn7zbxAntWwsyWseYD/rLDbwkhl
a5IPV85BAgJfIVH83YeuWKCf+mgJRmTcKu+3Un7ZqjjNtjzerDhslMPY6xsz
M5kt9pRxEZ2MJseTYqwag+TNXREOOVFccoF7XeN/47c9lphz3NVoaBJ1Xaki
PnoliTQfMKIbRgevr44tqOSbScugqC7sbMOM6hn0dQX64fsfL2B+p3I03HEj
IHSZrgKbvuTqOu/cI8Btjkc7VNPmo2jOK+hHI6VWOaoYOeKQJmcY2Zh+MyU8
cYT3f7onPAZGdPH/XXseGMnjpaDLP5Xi9SMG/c3eK2Ng87X6VTBXs1veAxr9
s7lG0BHCm7gjrI9atJyB3bmvF3CyNaQQDmIODKJxK3jG5IxhGjTN0b/BjKOz
erg6qXIiirv1rwbYENHltzvDD3WjdPQC09mJ5Jh8flhQYVDrc2BLOM+jK6rD
/h+XQytgl27bh8ywnm1Br5a1tZaYVc2qNV0oDy54LTrjViQwQNqcuBhTzDFt
/MHMgjNfsAmiCZevkgsJKs0lkb8iy95Z/09JQVz1y67LHS0kDtB+oWg4lACy
oAGMAtRiPPIRtO4yU11a81xLdzp9D7S2rpTLDrPBu0JUuCO514IvdleJTcDV
+oX1Mdk5NwW5vHdqnh+GeZAGvvjLJt1IA1XqM4qAjDGIl00T/z/PmiJekuhI
KxYU++HU9A6o5Z/vNFdFJTgDn825Tz1Ikxpig2hHUjtVZcUIW+XvARyAfUdy
hZn+XpxClshvbu9A1SMDkxESUrBWxPS6lDmE4blghGhWYCCMUrLx7e0yDiAS
qvhARvRerLqpuo5WcvfcbyocX3cPDGAhWCcgQazk0C/bhEixPtjNu2vc3bC1
i+Y8Eo4RE7t10ZUJs6NBNQcFxFzvnvL7qIAUOLw5jVbLUJzyy/6zvXxNnA+U
1fhCc9mb+vBsJTaLz3VyADYpb9OqmARepUdS/AQPwZ2ndlPzgfhs5MA1Qwhi
Gi2NL1HH7FAEJ/Yd/6S6cGi5kRBenjwtQjKh23txegmGbqBukg3UWgsDt2YQ
e5bXd3ulUYG6IKUT6tBKIFCnrPHT/pGzi4O9F/u4Di8XqIqcIjkB+yrsT/6V
qz8F70eNPvr7FqYeKRm1GWCTQjk//IltlPHLZIcyPHmPddCBKhD2BFPuomAh
nNyZqoUrgZqJBhChZVya/JY7zKfo3fS8kfY1fLZZu0ztUaBqyovolqNJNUgz
gaAizB4/HQt8PF7F0PabmfCX+js2zR8GnKkTVgHVm32+K1ITGGD3fkPQtknh
+VWtqgEljIDyTTOCUWM93LZZ5nnDrs1mzQDm8wtm882lWVvrOktDY8VkAMtt
6lH3xlTu24oRII3VWvUdFu/xbe7dM/r0eQZOuOrRTeduxCOZdJEGV3viIimz
7VkchhBSmNIafatfpCqjXXKAFNN0tQghOcbhAVOyrWa02L7Tmpwv8zY9/dlm
VRwHsebGCH3vuMOvXjGFHR/1Uq/7+16Zqd5mhMitDCY9+zHBNgPKtWpSPhNU
leRSx+/MnHsdrtJAourlxQgu4ZDM04rkbtzvxIBUXd1MmNVftuLX2bh/rjBy
hEEmnfgxuMWwtqt7DJGbiRzfxusrdZhuvXXIlDr6u+XigB041Cvqtvcw/AAf
hIqzRUcxJe9kFMRpLXItJ9G4t3LpfeCFZfUZFPw8H8FHm9DLL4nJLos1LsxH
kHtnJWtU/faZ8XDmC6TSxRCzg/+Gkl1AmKR6qF+ZxkW5qyn8qTKUHYqGfj6B
uFI69WCIxSfiJLCSiTM1mkXGUclebPsGZVV/La+9vFpYVH7Su0QtdOmcR+JE
7XUuUIqHr4yLjh040LzWjDfxepgdxMj2MJAJTuBmN1nPymlzJGTzC2GqDbWK
F/YrLXAy61iC2i+P2Aq8ZZnncLPT/YEeO7+J6kY83Vk4gWx5JM4VhiImBhlb
68UrvodCO9YEfOBBDbX/HbRspESeFhMePFRj/YuZ4StoLrApjUxohvMP/Fdh
1E7M7eSZroGGYSl0XUloadRfjdOji6jx8q3knvjrxp8tL1J3l9Q4h9q6fcku
DP66y7zNcRmDl0HpaVZrk9BI0pmQV4tKmWGLC7iNjbNsf/E8OgkmIzw1Z5nh
RnmuwI+LxrI6VWtE1gV5EIYi3ePc8QXJNzbMFZ4AgrQBg80+P5ZyL8wwqRsV
y6BcmQZ64D7I9WS7zF3pcfiRq3eyVI2lKGime1Xs/g26dRBipFKWdSt+gWKP
cu3B5Gus0Czv/3dYM2WoScVXixTK004LBmIgVjOkUt1Ns7ZwoA5oz4AYENzd
jtSt+bsTjTAMWeLe5ECSeY1ehoD3m8+Mk3CTVqGm6OeOBhE7S4XSg5lN4bg1
39mfv7gNoQKdsVqccJDDsrCe44ZTnqTXNp9dUTvWzVxsWFG3RirF1NTEeZsD
iisE+XJwy30/acoGcT31oewcnokyLdeGTvHNiYPEcR5e4qrj8cda/wDg8ZJX
pRODKPbtgLR10yq06jX3jJOMQ/EK/xRln+kizR87xlXV0ozK3Tkwa1v2cyKx
kh8iOSDr1ZEoSjjw6AxgR+8iBWcQh7EFUVzX18xLCTOmdH5FgjyQklelozJH
PXo7WBC6RXUzr317vWykatXAzOJrSvk+PvAITabaHG+TE72XQPFpZUnA9a01
m5KAl82s+pdwzuZ33fQI9HaffKc0iRaFdrV0AA1bKQNKsHkQwfFtYQREzqB6
l6NzasgYCymgr5QvrrsaPWvkAuVHI51hluo6QoLJa8BvH4+KP2tas/BOaNp2
x3qaRJFxFzEpcBdI6VVUHT6LDtUowj2BQVVoLibEAhIW5aSOSdzgedynakfW
da4czd3GE4Kqg/JmElIIxX//RbzjnPjYHVQ/KUqcA8DpvvCGb+cuJxtOphDC
OypAxP2wVTyJhXIr6K03VyFoJx3KZIUnUc6fTzKqz9N+5WSybqgRVim4mAyS
h/AzEq76G7liL9AZyTqtGj+FufnJkF9r5fGGtbx4pO0vDLXPNmTPXYepXBaL
a1XmIxoISt1UD3eRwjel0xsx7b6yI3SiO56HthbpKRNLE+c/x9l1ohOYPE4D
Dbev6yOuMXewVbaq6cDg0JE8mab8/VyO++yVm3CsjDscM4cF1jjrEfRcxtQw
xcUy+d+kcGrRs8yc75vkK6EKbLkLMGjytBAwX8ja5bI6xrg4EXti2seRXCi4
IIzR8s/bJVnpOSqaQD2hBl2nbOEAM4YUFMNvuHrXpjPzQwxOKhY3v3+EQvP7
EEd8HlNQZynSJbTkpMuRu8qDRBqxQdofMvdTL4S75Ib5Z1V2EjRAUvPezkNt
C+zUXPdfjf/5Cbsb10nOUkI4Y5RRalRPclpd8ESARwCPUBNCDXoZnKOsyYv+
lnmvpZvGeWz+NOn2kX8tg8ih37VTgur99yKdiO9twMXRWd+NjLVEUN+x4Ik6
CAkPRibNqT2qbEna0y6l15yGM02dYNNgFMR1/GOgI3j52qyw3M4pcbzuXWhT
LgNI5h3ykGFY3KDY8IoIIeqFln8QqtpfOkicI8tsy+9OFhNb/LvoUraLSGDx
+ocMDBhv84iRBduPHojeAHA6wSqebDEBbwnZt4KKAm8RlmcegFd+mE0R+O4d
k+fgeomFi88gsQEzlxw2elRXakIqslgvgOpWBbnBhD7/hvixd/KdgOh1U3Gv
hFa6hc11gUjHxrlE217VBjXPNagn6RshMtH0z2X86Hv83Vd0oWCHDhMJZ9fc
6NBKJGe3ylxvfyfcsEOC/hOA+0kBjfErhrWntTLLUWA4828SnFAz3Cu2fpGE
zKHsG4PqMdq87YdkDVRk7EBR4tUMYb6cwBrzvsWlC71PQmwNSV6wbAn0BSFt
Z0wvWLJOduKvGgvmWd5MshBnZLZ3hCKDZzMf0YfnURDvCKINhSh2CJMiJV2s
ngKkU3lM3PSiVb6fvzr9mBtzqgHN1k0UtVtgp2rlH/L5d2a51BScFpadMi9/
+Gpz8vqeBM+7M/8Z50/3qs4HrGiDs9d1mdfKWGZWZvqFJH9ffxeTD4BHK9LQ
gRj1iC1RqFDK3ip6o7PWBe6CicY4r7e8KEwrTozr9wrHK1amLFq2x9S47xKf
tUCKQNK4UXWUpLtPITSu894bMg3mIq0AFI1fkRmis3zUREevd9FuXdNwVoiC
hHq9Dw+66rFwu2WFK5jGXGIx/dz0ZoLBu6Sus7aVKVN1TziSPoya+RwjJsTv
DJaosXVGDTR8+jf4yTxCnjv1qqeRN4O3buubq+Vuj7ql5VvODrxwSlzSVt1+
THSLiRwfPlmYqd8kVcvfh730JwRs/IYVWinPnb01OlKNX+LXBUbNvXpxQQCy
2iSRW4AaU4WWlTdyRivLnkf1DkyjHotOmensQfitnLx//0Jyv6uNcxx7SMfm
fqz89KP4NmCX7Gtodu8BVbTLahvNaZ8g1S0jCGBBKg6xMm5j1b19GCPWe+7M
ix1oAy3fuRUFjPPCAADWdaCk/hEQH+1ei/Kz+XOzjKCs8p0+dqZeKWNlyopA
gwl9Qs8bIM3TS3bBTYqbDQUxmP734IKKt+4vI7ptgh/KwZykmV0Q87ISwGBI
+vE3Z6+BywSTawtmlu3H42etGbbyHsFLHp4MiKdLAWmh/DR1z2LPkGaaY7TQ
YXu1ypgV648/X/rgSQMC4+n7ZRX4uo5aRJEmyuzQMOe29KYA8aVgpVuojl0V
4aYNDJGP/qpcgVSogY/gQOaQF6JeKZrGD+2h2whZDmdezY5rCHSep2EbxnJl
szase4AOhHssBuwhAooAvnaSX8xdnWUi+SFpw4pqOO3xahOymS4U3rPiN62o
kZSE637EBr0i3jC7fbSy4owD4u9v9e6OUX347ZE5JBc9m9nxE1ekVFog9J4E
KwHQVs4SRlL/234BOMV2axCKWuHiWw0VGlsuyYIE8Lyox4WLiXdPFkjSXstA
Dd9HXXA1KmGfobz6gyg0+0jpy0FD/FXbWN/qQC5Rlwugsv/h+N9SLaGIuGCy
cBgRFGvnRTDmj04c8aoL1x9hdxcLpd3n2H4mXvO8OkXiEE6eY4S+m7OQsEQr
BK/t0rwoFuwrjcbvz9tvEvfyEZplCiSenkLBd+IOtoG6RCxQhxmKmlxBi20Z
aVt+u945hRVltS4JqCzsNZF8i68O6Kh7IGH52DxkdIZg99MIn9RET9BqHu1u
BuXh98g0xePZB1FkDpzehJ8LYrBqP1Xoi+HZv4romMnnlZJFH3koyOojaGfx
gz43O/WNSP5KHprSRDzyaslVj8Zkupo5hebKagLctDOpGe0ImhyqIj+wnByU
ZECc5avkwBWGqNCqgZ6moCs4n23lhxMavsWtt4YbiJCl4ZV6/Yv4jgmK0elu
qQ6XHXRT+4PxDW3BJTqnFOOX4mEUi7IrapetzNapMXDbL6/MdgebgWznNoJm
99e2lJeQFDzboUFswxWZ2+7jyuFoFD+dLFpfT9ewe9rZCRjbSRMhb7gxRSTk
p3BUtea/hES6Zxk1BfqDggGdil953eoMycZqFd3+StybMlxzeTPIBl+UR6/d
aiT+EMLoljeNf4ak1dkGBsg+DIZTSxOe4Yce9kRR1abzWq90n5W7RULPKnj6
IgX5325poULVcIkWmBnDP4OIhuYZZFDlx9CoWpbuv6n04Fp14Bhauu9yU24B
z6YkS2BQQ5flXHbOXBn428L7o7pO3+6pPZl2SK8ZMXoTdca9X5QdBnvT1Iq4
rEJZIs+unxOLZJPeXvpS4RCrLBtTPkg1Qp0sHhq9HjCfWO9dNVmeU9eQ25D2
wlt3SsdfDER927All3Aryf6/Z0VZGMwv+0pKdvj1wOQ3U6/e7EFBBtvPvwMR
lpMchQnpeJ5LNShpSqwGYUkOHzrpE+QE9+CwwGIs4wIj7AVFE0PtIJNoFaUq
zuSv2qZMQGJftNmpPs1pDiV//QDY9qO5nyH7jRvMdRTnvtvk7h57XynWfUU9
SbmKQCW2XEU2wXQgffW19+1w1EKbrK/Z9QC34hCcUidu+3Lup/il0v5acHSl
gmr3VdfDYXaBIn7m7X2iVdrkBv9QYYyYJMyMqUpShTxKhsyaY7for/SkqjvI
qMZm1sDsEoKmBh1a9hyYapbRYWYcK+I7BwYF2Bz5a0/GMBZQdWdQmkiNxmWe
UR7pOy0gHRFjZ2v7ylOK57k0zWi4zkY4I3EMwm15r84crkBfb+mf/Ke15oTo
rAo5D8W0KVskTBMptHfcdWCynw5pAlmAGv3dY8nCJL1TgTEQ/s5SIXuwxBYO
19j/rymxGkPZYeX2kNtlNJUqHLgxc5BREfvuMUZ+NQdyEaoaimrE055gWbX7
kCKWeHZcZeONgDpEbswN5kZpFM64u+vMGlPeWFLt3KtNG/99JSkiZwWHWY0W
tzRgu1La8hcRbD87xFnE4uW66WLoOElF1bCos7hVoCjjYKMk8g1gCykVU1S+
nNEA8vKBzs8G4j5pFDTMYePW4FvDV5/3J6dVSfCb2+N/4XU8rylpuUgW74bQ
9j6gHN5GhKtmgT+E50HWGFlL80Rg5z/sxwb8eJ6HMCa4p8ncwLaKMQx9RzrQ
yxFMtWiLAZNfcrUhrUMGzbaFkyOff9A1XyRqGqX6Gz2hrgunJWWgyATgDOWF
4YAfqD2B7vHD1ND4EGzYC5I8k/CScx9PM60rj9da+Q1ISmarhorHe/zbZpX8
HmV+1FdzqT2+JjR2PXXykvAUUmy7L4iLbyfuWJKwYdSHgDYaXMgv9j9AhOWh
/XIdGF70OLs6rrhpjq3z9oQanhpLTwjJtQ6jmWvsqBpjAXf5S+4WzW0FfgBd
OmkDHQGfUdy9sPECbqbAnruIhQEDekJ2Ar8/JIiacsuvgOyKY0py2yV7/yp1
hSUBQlNKYqWwqfswEruQR5Pru20Q5XbAIb0TOKuPStd4MHyN1+r2cUACaPLp
93mIUgzmzZehoDPBSSo9lMSi3wnR/7++kB4Y0VM57CR0AUUpIU4jhVQeBAcs
LH3NduML49hyXkdfSmwffUE1wHFgvmUh8Xzh2t6mBwngPACz4Hk8gbcEjkLt
7xLtG/O1UY3+8XKn/eqFkl23zMtyERJyd80EtAW+Cw9++4ThfSoa3uzOk9xP
evfoH9DexEk0mYtbq06Ovk7M6B6aUQf1zc4U9w11iEjBI7qrmDYrXvp9aYdv
A6FJejQGCRgxbbwDDF2NmcZwdP4yRCCzuQXgGjWL9xuJbn7bJamZB8OYpgPm
NVG/0LrR+jER+51Bu41yvIixrG+4tqG/zFCi2XgZQzRkdPV+ZOmcSLZf8PUZ
pp6RxQlFLjL+zh2hWWlBh99SqGSt1ixLPQbQwWZJ9btP+xeDLo9Xs8QUII4L
telMQdhiPK4DYl1toT9Stlu2L5OSsYneqRaLA0YxCeCQdG8PlTnLpVeEXhpW
DbYLZqQUVeAaRA9VML+MwTyY6KrbwButWPLs6wDN1rXO9cjLxlmkbMEiLWjx
UecJYmvMopfHGqHZC38cCxdOFxQ2Ivce6RYLicVwjdQpucPrjGoXLvrvEvRM
3xatU4KVTPGSl7ni72fbIJT3J0nw7fRJQomS+Fjj9d/zI7dAKzsNU09Xi7b1
QRC+FlxBoLHMhrcdLhC1U+IHM9uV4r3V/TFXXDX16RCZuyMQlDH7JRx1T5fa
yMT2SLcBsfNuZc9JRQ29KlLWQ/IEsTyftTKAhTELOOyuQn1HBQ1tCjtwXSU9
Fm+4ctUU+Efv/tfgAbMFqw7c6aty08BcFNpmODXGHMuAfliW8dSa6il+D5tz
gJ5oKZigmVkwateQjhZVQ2Z/jMeOyKWpAgAZOS5FeTXQmE7RPi+z8BsVadfm
K+YREulBahbV+AkGPSxoWS+YgNRti/wqIVqz6vu1haW3s9HALMC0toDS7upr
sTHPu8tOChSUsS6q7YStppZ9pQuwnSABA9jClDl6PRL1MPj6YdjefR146p9l
qUodX7PUrLKaXfiZw309QG4bnuUvaEgnSO6SuqgqZLGKvobtTh6ag444c8N1
/gdgAoN9FrOL9f7lMc6+dU6MZmmyvE9S0ZONN/guV5OwyBumQF8Penu1rSWA
dI43A0kWMZLLD3c0xQL+mopBLQFOA0DKF/eC47dQ1Cx+sx17GP5IQxDOy775
fy51BCIp3wLt5yRcogLjXo0iy6ex/0idL3INqIgVOOO/fC0tbqhcZv5UIfL8
eZsvYvCftauBY0KpJL6JuB0D/+o7fHsyBX3XTGpGMLO+r2nUWpCZDNdoYsPG
mG9q0oOCkW9Z07qMxLlXhHeiD43qaH0eSZKyhoJ9AivX7oOLX9rGoFucCm/t
47AkZrpCveX2JNtwAqjDq+IKv+XQK4WX52X/fhf6jXedS8m7xSYijKRza95h
XFqHPtkPsEr7VF8a5T3lWdzUZTahaAoz+mW2DO0szX+7lBaFlJG4txC2cJX1
smCSLUXvGHslezUx6TOSsL1A4Wp3NZDsKXJTPiagyYm3rxps1gJfILMe0DX+
VwKaXm0G3c094YsoFuml0hp84f6bg3f83PAiZw3uEkfQ0hS5J2pnvOlaoqgC
sO1Lsr/zB2OJ/y551hAljwRso46+hIzFyDn5dP6LecGoiB5PCcYqAFxKVdGi
H1nngAwb9eBaoJHfAyMf868i8PmzxRdFIOtiCCiWZ9Pm6Mx8rM+jZaFFOwTE
DTGE5ft4IbiPFUQH+xhoGw4WG1hysGoEvBvyN0O09Xtw5SwCFmt+B7seMEw4
mfXA7QeRrzsJ+vheuhx29TjGvK70jVmOABqgGodbGNWG20tG2Y0UEI26kHfT
DbZHE8j6e7JhW3KNhal/JlcVUB2VTDjBUO046qqsKIZiaHDBRt2h0DluvXQN
Qkyx8PPl6JfmgSeRsfQb7VtjIyI4jTjBPlxxN0HO801p/QFnJOiS3wisbTBF
TG2olVBFc02AbpRUdLWBCTQHgCst9+4LNr2dJYW17PK/22dLSB8zpM3ir4W1
2IcKVKSLdDoZce+LchCzUQ/PBiDMGpelNtYCcl+/AZz04Sic6woJtGOXjbOk
5+tqxjQValPHe+QBTZg6+FsG2CtidgnHsJ9FmWiptMpqCNIHVXr8Mekayjgf
ixytlCKVhOpzDhoqICS6X0Bd3tx8kPqskpnBloVRqkw84npXUIhJHWsUUQrt
t+HZa/Wsrbl0ZWo4sOxrZhflVaPEOfgwT00kaXjv/6iZ7hrS6d9IRajYt4ox
XprmnK6hJMs+UeWwn2l44fZAxhc7CdDbQTtQeH3kZm5oNKsCD8kU+EwRUf+j
emnNq/icyAgvkKflFgCK5xxsUDVQfUhDRquHkdJHPokWiMWuRFYxzvmMi4Kn
C1d9lgvFSQcsNSDnYK4E0vY4SDPlp21xf6itbouFQL0ld4ddnDjJ8pyHOxrD
yvxa7on8OOehTDdTF6sIh3gTRi5MLNaXF1p9Sss5PtVV16FkeCFyx41+3xCl
Tx3hzKrU6sBFswo3oddNvwFkQOFY2UmL6eK5CGzIHQWmQv+skJp5DMSiTW0l
CPxo7w48qjNl2mLVAq2EFKkT6KMFV9xTBoOxTOJKDc8Hb5SuiXO3EjlEBMxs
u3G1/LMUGpbMO/yuvsoMGGlvAVglOHArHo2EP3GnW5izW4nJs++HqcxKy/8Y
TLs84b3bUyDjNXxM4V/DtgB5SH/cephhYyWtuOEwn8eLB9MJGVuf+0+HACqJ
NE19X/2e/F9D+knvHALvPmXQaKlUcc7Xw8+ZHgBu0XzGUU222GpkSE+NjPtk
Z1uV9XhvtHuq1rqmNlW0CyeYmgivF6xgScU9BV05jdktnz75WzFoMJomayzL
FCplFfYsw1vkdDlRouaXqfzT6PEn+aT3AIQ4DCdVu+tOM4vaBaGWN+JmKr+P
ywQa7psCTOvL/nSGcpBoupTR/J97D+cgrACPeR4lKXmtotm6fRDiGJFe5YnY
waCzXMQo7YgY03aVNNsZnsP+WyA7/shlnm/Yf5YjI3B5NtWApQunyhhU/VLd
Jl7dnbA1TW1avRPIwwQlyosnff3lRse8PdL9P4fzuRxFFFS/eHgQ+tQyumQJ
Z4DHDReLTm0D5l45yScOcvmgVWfoEQf/K3yEWZwJX2o9HQMVrTZ2u9ewcBSE
yCsalhdPt9D0NF/PajrObfA7GDeCzJi2hf8KIq7teOvap9CfHE9pFytkaJhA
JrL7uim1ixZUemfgrcXIiUIcxJG2siU4++2x4CrEwmvN+nWMXPLKBiOmv8eW
pD5q3t28cLpu0N0ApDAo1+mhBorYrA/S4a7+jWLBeDVXih7E6uot18GYB9Uz
Wc4692+Cf/4+OUiTJKo9rcofyF0/JWZxaOxJwxn+X3di72gpZZ+F7wNLd/w6
UvRCbMLo2tuX3QaY0VnzbHAhrIIBGYMR5ha+r+B7MUDJIXjf5o9qf4Os4vKt
I/nPuMOktWVIWIPmnOgABPV1ebNUjzpsRNWdSUzsF2RttbOqWeeYTPhfvS6f
ISWtjVSHOrTuist5ShnYUh0L8r8GFEfI+mMnp0hW8NlQeypS4NilpReO43iN
grI4AfPFosD4P/L44XvLbgORBZwUJ5xYgrQMvO0119QUijJ0LMw0Fe5EtRSw
JIBTLLeDeLyOSWz6vXRl3M0yO6Dmao+5D2mbU+EhKNRmBHXl8HD83I+UNr21
ITdgBNk9Hh5KxPSbVQDOxP3KqhjGFnkXuuZ4saJklCQTXwm1VBH9btvddpyb
AGJkKvEWnt5vh24yDzLCJKZG+Czz0+vYGDjP5YqlN/x2nZgSsrnmPib4mkWs
HUloddVnjBtI1JUI6aUuQoctfdVUpilvhLMssd4iLypa62X6PSIuddNZMH41
z4af49L2Nt9T49wSdDiQrn7YFOO3rzSmAipj7I0cWX3LgBKXLJFGMg3mh12m
vh8GLLNxclv3l+bZ5wFM55/70rVqqX11A9GkR579zF3pleJmrZ+nBLoBJHi/
K1jiJnVzQKIYHTShwjiZKchbqVu3UQxS0Uad2Rmc9X2RIlkZJLtMqCPTsuhd
VlJztgn7s4jtbMXT+pWe9/vuGis6IPkWdpyTklvVTf15PPeAaCF1BbdVnK04
4aZ6lWyxYXBrKMaazQAqwIqH1g5kXrNfiPIqSWNE37WDtHn+6i74jA8U3PLz
gYdutMCrdtEZGcckzY099nRZnlKFak07pobwQMpOeNGi1e8xv7RWWmJFUHad
VKZfaH4QfgznB8c6SLR6/Bur5e17RFrijP5O33vi26ZHvlFEbZbh+9PdZXfo
UrYFbwwm7ZZRtNaJEsmM5kgFW2Ab2trXPZBUECpsFSf0gZ8xnRUo0LIhOjmU
K36CBmhR7FSLMN90CJqbrkQCQYBV4DUATSR3yN/beMpMK9TBn4CUY8wtdmV0
4frGL/1yjl5JE0CuHhbMJzHXvcA/0JjI1J4Qo5wDg2YRFCxqr+sFIMZ1wut8
cSSslaeu+DCPNH+SBfUK+mBIwZy3ZoQPjPun+0i/MMl3uU6pvPTnGQap5/su
ZxHCbdA6HV5FyHJ8j/+93S+X63BVVuzQ0RDQ0F+GU4mn2OZiwAALg/4K7SBI
z7ygTn4HdzFn0GWjs6wcHVZfVBvt1jH4IA1IaS9xI+D148e+5Ep7PYuqIwMD
dCSoCUWgGbfDlSAiUf7BiCaDEYdUCRbw2WUN9G0KgTCWhmnFpZhfgHHiDyGu
30SuBfdBLodK9nO37HZomxeOeydWRkX9rYUfKtievKs6Ufiq5cLuBb/4WqJe
FozzRyXWIMf+fKFg5PX8t5WqzRUndI+Mu3r/1nbgP0wVj3umlfQt74jfdc2/
Nd+1EfP2W94hDLzLZunV+Dgdb3jevtNlrfLzKrIdNFeX5UxPQFnwjxvpVi94
pb07vMrVJr0fPUZW6BPYt98SbJ1mGk9SUYKML3OnxE+BsQrrmT+LnnO+2fsS
deGC1DkFniPXsaofnoR9PRooXgrBsAQwHgdOMme5hqShh9kwV2+7KsWsV4X9
Yg8uOhBR3E4nnKJ2OMaDfFU04B0U/tVFKtFgPRQA/6+s+F6H/Jgz1WgykTyO
803RYo46MRWFWmS8EQc39DoTlxJ1R1cs0BjInPQ3TGZhlAOgR+EVdy3R2Wjd
hnYZo0q2AS/DsjITC163Hn0Zc02PsEPBIYKB0wFMTZf7RncM08HLFY/QNLE0
M+6BoWP88E0OgEuIxzgw7k0lyfDw6cQgIwJDOyGiDg5pzqOQUek8Kl73CISE
+qBuWLZAX0Lm6fYsSG4d1CsQ2UkT6xBiIDHarU6h4/VZtR7TRqvRtd4qNLjU
CJdYHCRwAQf9ovfKBLSqOCBtzfMYDfUlnyPqiVgGGrOpofbuYmUkVILoeqGY
UGHdPo/+uXFaBPwTZfZBDH7zwKsZHwmdsvSTiPeJ4+BmWb7ZcAeUFpYook8P
80IiBTfXGuAKInOpAvdFJ/OUPjW/c8B0ycf2kXZWtpOAIn3tTU8E/mgJk4bm
x/L77nduZcZSNQhQiwdR296FULMz+fIAZKacHpFFabxl9b7ygsAATUTAv0Lz
2O4iZBPXbU2iyHOkWjTO1BKFwTWcPenl5OX3KqJDJK22kZHXeuq3aANjshI9
ylmItxuhIul9bkAjd0WsWhZ2Cjowe5MmxeTVpTN9UKQysy6MMEgPweu/l5/f
WFxHo56q13fQHCM1Lay+hd0IiGBh7w6OtsCT7eDcy93ycO9lAplEcISDLbL6
9IXHoecYk/9z5ZwUbIFiJ+qdCXwP+xux6uJHpd7/ZyXquW8v2DQ1jIE/bNIP
th6u0xxhcy/4q5f04sAMDmabOEWB+1sHJC/yK8bR4yNd7nhYPsMpy+sMOS+H
t54E/X5e07t8muMSVi067+Y6VFuSD8VUlL0H0GlqwXt+2yCYKM/fu+ZTUggg
IrC8I5/0gaCmnIbBJ9LimfhDvm64LHWGjo5PycaEdK00ho1wl76px9ucw0On
0ivT0q/+ZE5hIBSCE6XhYXagOI1ZVd67agqyXvLFk3v6tMouLgmPxPRH5SMO
ieAvyGh0zfILxGo3pr2HADyiZWsh5pUpX8oP6eyDqpcMZN9RQvDyB6oaHqRa
eAeERtT9cJkJVis23zwNQZG9t6e4yPXh7YwVAI0OUjL0tnsuxgxLZ5bxM5nb
wsKyc8zhbB73gdwBjfCoO3GtD+bT8aADxcqMbPB2gMtrknA4mA435tllZwh6
NA6orqbyhII+JwUCPNNDM1k8F9Uh1tRA0VYPHdWx8XprlGh3l55tf1UBaHtj
TKYzGsq5KJkI3NdJuN5jmvGCcui8i7Ey1EZNNYe/L3FXcD+g/TLDEUXm+DmZ
eVQI0ODT0rVahfK0rMfhlGJQgkC4862fe0wkt1ctillxwTczfqneUO5G0MNY
wirvjAm/45xSUhLmfc93kmzAaPbg3taRLq6ywB5WUTVNFUxSHVhs3y2FIbcm
TGK0Rc+tivF/0FPP1vcHx9E0+cmsBREvzi2LAuoKHQ7CBNv7g4HQoCG47sIQ
Zg5X14GZTXBxMKCFVP2yH/TgAWf0r6OEc8M1OM08Rybf63z5tnUIQHZ+cs1B
7Dl/0xPhgqwLFoDkp758NJjoW5tlpIp0/PzmbiHjfRxeMtF2sGRTIW3MDxR8
O3FwN6SlhxIhwiUKl3ovHRM0s6wTt6QtjrFUm/GT+qxedZvewa/+sP/56oiX
Z2ASz8fkhLO55tuEC+fVLgS6qe7Q3fcPc2trluB4oYSF7oYucHK0vFTf8TI1
l7CqxUc3ZnYwCIiTi+iE69BhpQdZcthzcY08/piCVHbhtvVVdOEnqrIwv9r+
hZaTBRqRVfczVbLJaXnBkcfunXASkjRY2tabo6p7VznR2VekVLcmUAZORSd0
xRLeMjlROrCDI6kDXUOgZ0jJCJVYWzDVOPAoC5XA3xJo92KOBO+Z+8HAXRKK
X2hB+i98JV5zjM4SNUq+SwEiIxTQpW3hN3UJgEFA7rvT0iqZ5FjWS7/BUz/s
3j4MmXomqaliyF69UAT5UA9J7KViFAIdrh/n1qnFSwhHw5fu37p2r8Cmbous
JA7YW0DwOe4BEfj0RtzKZcqaufPfYlK47QpEagIfqhrt1mCkQt+MG9FlYxQs
9yp8n6qWKgaLdOgzJrdfxiP6HSoW0lfNcFzOGfoFpQgQsIN92gLw9HALvR4f
zd1CzHIAtcRP3d10OOTnFvXxYrVj/fVpf58SwYVS/DC1WqudNTZKuyh7z681
h/awTvzFBaEh7XkO58JBlQ11Ftlpgbta0u47BngeKW9TUnPWYZnB8la8nH9E
QKIVsYtDM2U62InT40L9t4sZEr98T/zJAp8H0rhVxYxWZCr6v9vx183yp7Nd
/rBL2F4RAM4w+Fy41coFZHDIgIAjD3rUhUg1vkDzxw4n4xOaNJhdgYZGoicS
5A7gFWoHnvwUBvBjMlYpfX2VUMpgSToJEFdGoOYpvwoAOkCoF+V3zC2DyWYv
8/mk1kDoQYPMR7IyhpAv/uqZTBEnPMM/mdySQEvTIJKuHwpvuZLLW1R1SWKh
Ohn+z4wU4GIeM8j/8XGhXlIub8k3uODGwht1N10OfRPCmFEfhEt0Xwo82xRo
hMwcP/3NrsWGW+Rtkm+7km9nx3P+Z6qLEmqcwOk3r5gi0z2fgR2XPCbd1Gv0
rM6ocm/wVVPrYf7nX4hQpct9MdkCeBQ5qtwfwZaKF+4klk9qG0Gq3GWP1+96
A4HxfMwAKEpogxa6p2i4z3M+z9FcrvFtK4KgUjIGxfeSdYuHTIx/wuZyKfkg
ruovRTfm3vp5wYaZ0SaAB3GwZ8ju51uzlmo3RjFqcoz2Owb8WeeWy9MzIrJt
mJd66g1LQG7wXEYSKUIp/pL04+hnhJP7Z8e3cKaXGRgZEix7ShfV2zvXVoUL
097skD6ggFmNVuh2cSWVlsPW9i7vC3+I08ZLt0RTNsUbi7OYrxvx4xAZ1yV6
nAIgbhLV+mQRMReHXIgufIw9y3VMHq8P8fqegAe1GdD9J9KQfnLwClskz8ro
R6rKg10pEwbtc23aravJuhpWPGGgPLKcdXL3oBtu8fT8W6x+6twLj2VX8VUs
/lv4qZtQM7fMWn20uBWgi7elkcYJXaIDJe/7re/8fBw7sWoCrtcWzwjZui//
wrG6LSi/kNbSp2cr8jI4Ek9biNlyP7OJJLWcjAuHXfFNvxUSkmFL50kw+igq
5+y67TlusrreXOQZVQ4JH7bkJi9P4Q7hoS+/LNUX0fRqXFNbLaU+lLhxjamL
rHRS3jQZyecpRBACf0vn9NQPkLULxiTbNIQLYDDw63g4Ksy5ao5pAyufXRvG
7fcSPdNgEeYc4U9KHvOVLxEiLgusIzpoTqhU6fFFoJwI2SFXJUoWpbS1mmxW
SzLBY2e2xe/LOz5AD0P8QAY+jpRpFXDqUZlNrog5ujGAuHEJA/3tkis+1288
7HtWXEgxnSyXWxZc5zQzKCGs4lvjesGGoet0yHIwFNIlqb/9njnopPINf+4t
MBbor75l/oa1fHLnb9eoMcBm4bUeejeAlylpj2AwWxwZIG6o5y8oGfI7pWPl
w8/4bbXPDyZPueYDeWUbKZ2x7zcLT80PzWS1AzF9Y9THIeyq0aUnXrfdNpfx
UAzRimD6cUkVNVBNt/1RAu4Cto/uE7It9y+iAaHyULmnwXj2n441UbLSmdA0
w7fVYLneZc7U7t1/e2GWzpao0yOGNWP6vav3aPeKAc4xwO8ZidppYcoRJ8F5
NlSWOcPfyllN5SZIdgSfcHsniWj6BxFQG0Uw6h2XAn/X4/Zqzj6l2/yNLE2q
UQmzvJJ13Xt5eeKc0iFGy8Zt25p9BM7EPdIVO2bsaFky6tP63bASZ3dlNW7+
4UdTLu/dscOx8e21Hc31VaZk99TeWbH474ZBqsl0mlXm402MhMp5gyzCOuxB
DWd9XYoR8yL2ZpKnPCkpU257DM1rDaFw8DWotS7O2RVbvJeScW7nXmrqqVcH
Bw3fxSS1TC9cvwtSd37PJZBNhj7wNxH4n0Hq9/sRZ6QnarZUzHp1ShrO98Zq
TNVkyyCl5YxTIyYPJStkj9ElMEi3NnXN8pshtCC+NcN/+nVTCLx7yVhovGk5
GmAqEAGCBJcpL0LnQCFCVx1WyJsOweqQ3hBCV7s6NStXm5bkCYXjqdBan0vy
KlRAzZARQE+3sEpR02p7ueEqwlzE7Gv/CcHp7nnZYnp9XLKIaAVyP4OImNS6
tWhAHT7UkHF75uvHlsIVCckY0690jY9LrJRFgtWhTnhuoeAEWOiGKB1x3Cw3
mdxO1khYdhruZ+k6eUSScMbawcZKQYo2TH2vj8/BaOSQ9XsVpZ8nOGR+fNbL
0DmXyNBxPCtvo+7+EUKZx2neseEdSXNc36lKWDMTXeZWU3ELLWdDRZ3oNPyp
YS7hQWil1XNcwF/TKmFgs/3EL3l2WreJwUoF5Dzno2/MXATeKBlleyOfz85M
j9A/g94ux+k/5r/ygZImHGy6p/znxGWUEoMeJnLzV2ra1b2S7Kzalo8vbaii
Ryf769Nb9Uq5V/pcWbITZkyfPoPOdl2+ntjI5v3fbyNfVP/QJ9hd+KigV8vp
vdEPxl7/2/nkIGP2HTl+CYvFNsPoiNwRyuZ2C51jjKbObvx4mqqYOMN5XgDJ
Hi8kq5Y+jnt4Xxc0wXdGdBuwXLdbrbEAJe11Utdm9xrSFP4ZtLWa6esPWHOP
qM7mRE6R8U6hXwQ/3anYVCJDlfSo/o7S51ykKVcq088N/4IplLL5FnYx9h6o
IJ0PSCdnjQmedNZp+A88CQmJp/0iuFeRmkz4bHTiGPtIBHjLWH1xw8tL1njC
+RplqrNahL1DtmzfSaVXgu9QbtM+065QW3NHRAOlm+8W8yNNi/wjiLAn3neO
OPOMEJjv2pfbyjajBzuHzwMNoP14pk/krRP4KoyZxEzD3uiSeHqjHJ4Njobr
vYgCqV7qHQKDiO7Zty4AeRXSSsFWWz9we93icTx89/21vPaXWZwQ9QHmQlG2
AWUK1fp4H9eiPmJhRzP9KA7KI7ttvLyqXGXSnDaVQ0RJytmOq794/a3fa+vc
zziZe3sB/IZPvivRSPoAoMZnOxld0MQ8kbrK/+lvppxmoWMcfX3Xjtvdlv0z
c5CmPuxPo/6MbZ0DA11hJhUW+sK18Al1xZYAINE8SyCad0t6Je5P8F6mTrPh
C/YPUcibY3w/Rrz67keNdDxtH3ZfpxPQ6yQNwPcY/ApOy0gd1m+I4NymenRX
Q93pJlpHwWa+uuq7dTirZjuDxFkwi/yqNYJ7HxHmSfRBvfAW2uxlg1bScWTA
sGKDW5UaJQjy/gJth9jnJPplLKEwRHZ7aDjCMncx6hEGBzKXH1hQZXa3ajKn
mqBPC4/fQolt1Qh8p+yifuHakirtie5wRvWythauE6AYIZ2eA0T+gUAPx6NI
i+elSd3JiXSJTLjyt7nUq4ppjmSAaA/wTWUwo0CoFzCUdGES+NPhmSeyvUvn
i48pegtaWyVPqswmVRcsz5x25RpAQ6ITcYw6hAJta9z9gBRqsreMpaiTp/Zk
ut0vniP5V0uiVvn5OnqB6oTVulG+Jikoj3KhPYZdswr2+eCJGZzyTk9qQiFg
PRPc9/0zKc+8+FYGzRDi9FjTxvOqmPaCHLylkXhLDiZLaLVbq4xlwEh+/W2C
NIUvlPksEVs5w6/ADiYz6ga3lS5ypGaGob0rREptYHa0uFHCzrTcipy8oQ23
3x6ti+3oIbyeDsnp5Curh3wDXhARBaanjYvmhYv6c0TOatRyWWIi9MRX7CLP
eK4JF5pspZ5V0CH3w40ISpTcDE2Zq2UYTMBL2y/mRojdPLwTfdI7ghNNE4Yc
xX+L9fk+Xxh3JiKmftlgTDL7H+SzeW0BjOfH43Nyjo9zus5jdyvFlJ4VON9l
BrhsxYUpeTmsHzBINSO+KTaBt7ddbzdC5wptwVXsaMuOud+X+69YarmWuh8X
zIKeq5Z3+hQ5K38C6yTbFETaN3xvDzNkkdKJ1tQKuDBDQk/ENFZH+Tk3xaZf
S31bwb+5KaAJOuTxAwBLjH7iX2kn84/PD6oT6TE6S8a6vEw9WJ6EJyXjckmZ
l+nhap+SZabsswEJlV7CSZR9fQ4h2/RjhCNJWuLhMFUyGmbS2oeab83jr9L6
FjN9ZSyVuQpJYde4mVA7GrLwhP0J+CKA+AyVfcVg5iz9SX6L0KUcvo9kjzyc
FkWIKPsU1aqOxEdSJ5xJFG9ylMnRjqlHDULiXd4t2gOjCyYeE3SVmkqno170
SRT6EPuHHFyWWGCOrtaeehccfL2i7iNJ1lG7nKeZT0kGOZExDAVEe1PXll/n
8t7GtO027hb1HpkO0qPhSKM7/oWGDMJJiSYQyCx3eCj4nz7yZD6jOlObUcav
rcUKc7SH8ZxMMwi110igZMAFeAAVt7YWeB9ikPxcbShC0iWBvIip9NV1zBa+
OyTXXUovWhCrUXlZ/e00XUTc7OeJNb9d+6cdkB1CUxOYqDnLH7TEvDiHPmFk
MB+WW4UN3DB9ddSAYmNavXma+mFerV+ozTNfMME7lOKZYkQDe6Wh2XDcJ+kv
PBINr3L1bfAEpKIqe5CX7cleRojaK/tz37UBWjgzH2VRNOZfKvulmfjgTmES
oHnGS6HgjP4xKh8vyWnqLTUsoCmhkbr01z6RAedbGlUvfl49U5jHPCNZ3psn
2EwY5gcBZD9pLkJO2OIRBh1kglCOycPCbLfsc1sSVkX1Wru8k9on4guwo2XX
ZJj3VrUzOdiw70rG6D5gs3WZUs5u45u0/XVTfKOEq8N0uCYQS8mpkY4IOuGF
aunJlTUtiMet2XjHYvrlkLUeESNYvHE7k5ytftCxYAhvfYapn533SC84MwhL
1pd+0Yrp6zU/SVk5UzrCreUUwA13qYS63LLGBTwo4fHB5pqy1oAg+OTtBmO0
T6YXm4ShHyiHri2M0m71kKj5U0ShEOjpg1J9yrMG0WTVo1sRctxnSBcPC8i0
S01j3No9we4RzytmB4D6PXiYILeEkdTGgucp98mj6pLTjHLye2W0L507vFEP
7oSgR81dPkxoXJoq9QHY1CoMDIj1mirIfpNpaAzu2/Pto70ibGFzCeCKRUVH
+38jJRKE/BSmwHdg0bHVNyDwW9V6LkuJDn3iO1jiDRnUFJegmxNXDx7rPLUX
3tLvMs+k40TXu0hRhrpfyEI4qGK/fEIa3VaeuH3jn94QODMvj6uF9Mah6cxT
YCfWfqf2BeZ1mLH2zs03P7OV02RNWCrap91fBVTzHbnbjYXlnM+8ERrQJkgY
F2NoS1ilT++aleDXcw8oPx0GJjIg9LJ81o7NeQ5ag2rlPxyAyDwnYeObGpl3
0bleqB+3LwzUA2nWceqp527rokI54Zr7QSTDuwkRq9NQ4eXJJ5YpHxiyJ3IE
qwZgu402i5Elv4aUQiHk4gONypvoI1oPyHQF1/JR9bPETnWbe0+5l2rsW40k
Vq5R37W7SJrPzfweQvq29YCjtotSXBgnrs+ADbDO8ygkHhcJY77U3Ac1xry4
t8F2ZMjlkEvHYEpjREaoFR0OD2khBxwiMIQ34XyfKs0Yhq8AQOJ0xVUZLiMa
QmJhvJjS2vLQHHCzo2f07E2UrTc5g2OPXQSH974uxpsVWqlOkBuAZKTwGedk
GJXLmAUpynOSQt8RECutod/N+fPRzsG+7u+VxbsREWYdDDx1RBKloJ76N103
FuaOmD5g4tfW/81GkIPvD1bKzPGLPMZ+ZvVdcjLuKdaCwk8KGemDKti5sxX3
a32jxGf3eOiTyadRljMDFsKe1MqD57o5F8fwyR+6RAHFImfpnTnxMmwriC9a
sx4owtvpg4YgZngj/4XOxhOqZ9wbCd6cqmwc9FGAVzEyaOEf7avuQk7qpHjl
rh1VyYiTvQLfytXyo903YamdQ1D2DEpViGDgz1GjfA777+xaJmuilIr+2XUL
EjrhgJBV6/obU809fXdahNM3K5iPwnplPn6EVqKpuANQ0Io1QQ/eyw84l9NN
0Dq9Cf9BBu7q269sJH1Bw0sx3V1OOsZBnkJhRMBKRWaVglzsK9I3cV8xvJ8d
NSDa2ivb3rJabj0W3Z7Garj2LerEqhlSyrYzR7XUinK1R++q44fNi0/b+Tn5
RsTu5sNuLdjTMC1CEkQhqzpmP8JC6MnW00oKqZyfdJp2KnqxgO9+TmGSKGvk
wTZQV+liyuIpQw7TcOSX/ZUHL3gwjCxipdY7Pm12Qum8wGhRt/sNpoZQGBDK
dJa2GVIz1zTB9DEh6KDsOGd5qjIH4hXjHoG/BDwWLUqY0kL29zf2mv8un11S
9ZHRoDOQKainacgcDyi987wq0g8/uZ4g1TTND/BE+Y+Hv/661/+ZHzgff++n
uVqpAPjoZhlDdXZ1hkB+RlImbnI3et6kFFfObtVNObLZvojGl75SuoWa3Iez
Hby7JBIs8bVfYnoqxs+SC7+r6gIZ1iIQjpwjt/Q196umRg1m1Q8Zi20RN06O
zxlmGY/tLXtZJzO6rV/UdGVJL1t7U0fAjlk+VHacn65Ph0+giupoBEP44OOx
WoK4SyzZDK1Lj5oyJw9KmDeBl/o6mnVxyh7ovolW3HiOJMXikjeI88cE+Bgb
ZFylzFuBA9dRYOpBzNdHWY8nKW4saCyVlneBltNW7ZTTfa+RTkJz7N4fVd4p
yKqzncuB36s7orDybtHpUyMinpB7pUovOOIwXogYv8sefkvZjQU7px8NvS3Q
AvnNHFN5T0A7AGfU0bidyU3N2mD/h7GmvNhy0zPaFS4PGb26GhagDMOP1j19
RwEsHh0flRbJ/YQo0adEfIGkO93J64vYZ0uzUvOM5c2Sp7oJM6d0CFTEQaG3
A8MgfykHENll/WLrrqJ+buanFm5fM3kAb70S1L24qopSSy8UG0YTLXS3y0Qg
a7fVAoJFDJZydtlbrTXUolCZoyMFZuwBj1i0+nBIGFccfi4ASBdFg6UUgM0t
nDgtnrv4/JYnRSrOeM3LQa0g2O7lbVFUEmemxys6wAVoEzEh+xS0D60VPwC4
RMslsznPNeWtddQXRZVUHvu9wQGrRF3hZ4/4WcHmik7UUNEid0JRZ2w9wa1R
Ki0pWdgYfs2s4hkS06961zcSsE2yULqBiZW3QpZs6kUkCgchEqqFssSY92ta
mPN2m1KSRc1kxG1pum91QaxXjzSsHaVIc5HKn9MJQfAxDsivw5u/j0GAN0wJ
hDk7x17RRaCavAY3XAHcn4aUYBjOl2DDqqDDe+k0otqhT1WuNdASYldpXz+O
AErpfJZ8NxO61eMDjApg8R/8oNgG/4fD9F/QRSfZXryYuse/FAmqPWefP7Sm
oOrFLA9ZyR/ZDvO8WKZ8Nj1K1L0WppODa8Od32J3jhTuEUEzhT8nM0GrZTgL
//sYlqHBePWoVtGOQYIYK9ens8n2p5BOvjQixd5vEoCVNLduGyt0lEBGV//t
l8zrHcuw/2r3avUqgFV9sx7DYORcZHPiYRVbTDUhkvJ6T3Io0uMH71WI7jjy
lWkgpW/EORchPUmttDxsrMB5jw1fxifoPno05bQCr5C40lIO7depF3iUuX/l
u9hZ1N9tPLUbfp6GG0L7vkI5Lej8U1CiKrABjTqhuHaRkF+IgwDqaGu1pP8i
RdwBQKm1bi4G2FDKM0zD3rgynLCrac2ae/TUvmkt8Wlh678h4FZ9A/kth4ks
inQaK2s83yQVLRHjVs/sVQSkhEGgNY8y/sQFFlW9ZfyPISMWwtKJ0wJM/SwP
C6Ifzpzzq9CR7P91vpTqFaAo5w796U3oT5f2IDsQ73pCzYLDO786DZyENHXA
ELiqzzwBF4pDBymBOvfU9m/MzJPol9meudnY4C4X2HapWGRFUoQdyl3Kb+zr
8IQj3YGioL9zo6I5cPJLtRVNwT2XpuBb1B9oYFvjnTcxVRbklvRyu0KSRwX/
lRNluqF6eF/Qb+I3yIy/ZxXLcjxkibTOibqjlE6wSSBuPcq3guyuYwZFb+IG
3ojii5PaMgIWULmi+0ZYQ0xwwM1ESgeuJu+6LtfEEL4shIA0vNYjSDDebG5K
skXEmdBJjMcla044baJ4cQCKacFrxgP438YQzWFQgdoG6YYI6z6ry+FXSaWv
FdDyqNKENO4tvlsbITPQemQR/9DcgVZAgsqCaA0ZEHvUNytu9LgTQZhmZDjU
lQaypQt1sTerec9D6Ud14ip8ltU71gGHkpoVuQkk8HLo4yENDddziFIJWPMh
57PGHMEprmCBYP2nkrvSXzCF8cMrMhhuv4dRvzpa7uT+3WRn6Vxfyv+K5JG7
yXaLcrlvzVTPOGq3Txhra9CQKaIaqdRtpdN5KlbBMOY6oON/Az4EOh37vFDq
FMRfu5bKemZZHbP5BU1l7GqvJHDVEwmv9n+xnxOHrhNdl56JPdIMK8wjmaY/
DA/yw4NU0rlI/zTp7YVdpNkjecmmwTntQkw0kxUo7hvPWaHyAF3RbJCKnwvk
Af+vb+Sv84zZqVFL7BUttS41C6fHEgAaasDevjr9wJaZOJzVyyPXUyMoTCrG
aFeF5Qbn0udMmt+BtlGCDG83q4ET+jTe0sYd67z5mKA4yknIb8c1s/PosDGo
QM/R3BZyfSCQHxdwG9eQoXJbROAblK7zE5wAdA2MAyAycAp0aM8jim4y/aYD
LLhRrmdqziCagin5ix+vOAUmezRnprN+vc8HYVpUMQnjSaSAn2ZW7p7FxH2s
xccPfBShu4mB8Z2GLB9YPmwhqJH+LWUYp4PCDp9R9jcwiF8XiqoNIZBza8wJ
XTAjTPe6J8qs+CFT33oRiD07x3TG4r7HJnDbrdC385tWIkC4qlIDEDL560iB
gHzTI+3ZV1BTV0AGcE6I/Q4hqtEF3MYsOSHCW4FDniSikIj/n9XQmOPgLb+1
tR3XoYpV7R0LkC6vNjKHWjxI7b5Z9q6QP6kY1iLNo5qYfHI5ZliOqDskhNdK
nyL9iBHViR4U/hcyGlPWDvQKsk9HvF40PWb8xyJ+BKHzz8HeXrzYjl94Xr/N
mhcLtW9I/J56jL3RpeylQ/tsUhBA5jWRC8/8er8H0D4no3gb/6lVfNM0XMyS
L5HEVIlq3iItKwm20FWuh52Zma7pH4IgelC8hvw0tKPD0TFN9btprP4knZHR
perbaEQAupXzFx6L7CTwf6O9EBcR9leP8omRgqdUxwTG8oyciIf7jenyJVnt
OaW1OVwiEgkGfG9WtsT3JurT0FMxBvKasDJDcr5TVmjGxc+Td3W8FSC0kjzY
Blb5M8kPvi8jimugKbpf/eQTDI28wu73TtqMIf0Q9uHHiwR8lMJUCXMqfXKH
xLAkzZgR/AQ36wqu52k7ruEmeXGO0uq5j2S3NrCBv9GanfpHzZ5d+k5FJ++j
KzofJX1Tic9/37qMXyUWO6b85ExifyS0N3/ulZd4L/IpcjYC+6Kzta/8rjgo
S91BO6rf/AshP01CsYyks+YJGucgooAV9wEAFIEcxLUkxjIdzarVPsGFpdz3
xi2fj2C9+CkmYXUywUJlBdVAhLE25eYSlhVc6rKUrpY5kdzfeCFylSBAZfkP
192e9PVbqdfs1papv4LSmkJ0gbDRGB6WMhY4p0a8qNr8Gj+Ky0FNTKKkhIfE
KIEskE88DjnKKGihzFfGef3Q3tCTA2Kdu06+ezL7lTb8k9AkX9zWInSlgrJJ
JToBKKddt1RUYHP/GqhrEaqnCJIVKiqecqtSfwLw6kaM0BRlJ2j3LFC5QYpb
D7gNMnJqIal+cPzODtrSEmzM8kcFdrGClrbg2na+P6XyZaNpum2zwNbU9nDJ
i2BxlTADfVH0+ZZd9jUaqFwVwR3e7zWS3sot9mt6goyyjj5imDF0qqo86CgT
OVRxxzxeoemz1fNn0dTbjIzW3VtTihG1yXqdjoRwxxa67luv2edOtZGzFjK6
15tCICzyjmT2WxfZmK1xq79Q4KRvHhi15KU08qBk9sC7htNgfmDNI+VnbETL
/OppFlhocdquLvicVeF8t15u+6aT9PdxV2XddVoHSx+VB8RMwXhojdjNpnbM
hKHpsSLy4ZOOFhs/+Rc3/20E+7wEkn7uCaeyGIw+Pvdq3ITaCQKcyuiENj6L
jJjG9UdIHfbUqwV+DI2hFbcIRaoSIKDB+hQzvCdKqyUXe0D9BYt4/3kBOUVx
2vqEaF2VwZ6r1faNFoGdegfu2edEE45QhJ+Mgb9/Nxe8v5PsrOEiyzLiDYzQ
0SbkBFFqafPspFa4T+Qbmn+k/hjOIQJGfe6BecV4FulL2QaYTY7RX5rG4l0W
I+pjroOmwCJAlerdMNYbBvn7tlarjxxMzX1678Aql49NlAxmHezm6n5aO+Cr
i+ZEVpNkVdY8JY4runzixhrqtfMTz0tDfNP27lwxjItmt6MsdzTjFpOB8hSW
9b2PUJcRggbR+kWbI0/jHPGTlNgE5iLisBXcd4LR+v4lHJEsD6mC5rDkYMJJ
RTjhpoWTWspjdoM6Sql6wCQxVQ8ICHxYvJe43CAfQmjePmR01GZw2vCekatQ
JHkmxUNBChuDFE+mtOf5jF+fqxwtnOLdPTcy0WRSwc8u7zA44dPXJKz+KSkK
RPMtH59WvaE8gPLZdCz+0zIMwtso3X5EfFAqeTB0i99qf9phMVtG/1DDPWK2
cJJZJ6EPRDZfDE6RvLRl9B7oe3Z67HlfcDmX0sa/960PflU29uORfA+hLS+8
dT22tyBQQoSDgJWak9XvX4K7Cx4ZAlDu4lQ6AJaPvtDibjmV/VcEW4kUUrLg
j6gMN9NBJ0oJiwRIXS5qnlfIAUdUyqvSwpJMkzAHy8bIOKwJvYbAY0fOWR1K
x4iuRAsduLLwbCapUk2KqhD3x7dtEGrJaWnCyg7L9tCgZI5p4KmTAWeuTE8b
Sc6RYIBLcdSOeGOcb9m2orHzgGOuLWdxfm6T7a8Z0LKccB6v5zqoHNKOb1sM
TwZCP2HM/nNmT7X0xQdz3nyAPJu/Ek3O5QDeHAzeNUF6J4XT7jxoXI72jINJ
jMDtKSGPYEJJdJQ1bGx1H4ixovkmQi2RH+Dnxe6rmkBoH0sV6/Ex+xJtKRR2
FlidX9o9xZjBFcwt938TQ8/H9wufB4HrsUZOKNJBahiapJExhPFnJfmLvU0T
B27k2SaEoiHjV1gEmHV8HTwLRnC3VD+pDFxY9GZ22QTqCoP4jhgzzFXGZDRV
RBhiQ94FQafnA7/+QXj4F8aic5RHIyDW4rP9ksSdWtx5xjVcvngo58t1tfSw
nPn32eTHVBhpKOCd4/33ZxOO0RM/vj1rgx0lKqSqNwIsUbnxpb+aCOEaEJns
AkvK4JKuK1+Od6FjDjaRR1L6wA48NXuMW8HiOVSaeljJuBNhwfVdQbo1zgBK
oes5SXVTjhFzz3SNW5yeX70sYYHP1dlE8U7EWUuXFIKAMJ3iciqYcncXJQd3
CQReC+8Gf5atO2ws4jOLrBspLMpNtKI3FXw/iNmoYLAZUUK6EgHHaISW/Zqx
6qu53ym+SVFvXILVEyOErChegAqe2b33ppsieKqZyfn2dkYNSJrxrJ6KJiFV
RjFQnNHUCOhSCyU8nVkWGlhIwWQaBzYa8/JU5v7e30HhhxlfD8cfsKKLmb8h
58kURiSA8v9XFINZ4N4mV1gQUvqbP2dVo6eOqRRlQY1SOV6C09iFBxs9Yclq
EAh+yAocOdwNjkMHD72MmjXQPFYoWPEo8KDmtR9XPDBRYJFrY09t+8d35bdO
UZRjcJm1q4vhGjGbxnUjIzqsFNuRdN7B0msFYXe7hx6uwkVzBuDvgCyv8cIW
qGDXuy6OnjfTbnzJQPYZmpXvdWhOULNM2feRRFdTxjDhSd+tvOO05vIR3Gra
HHBXJvV/Kg7S2LsJnub40q/jewH0WoZzcExnNLlvQBxSIGik+Y4F7Bn2klSJ
Uss0SYd8SYRZSTUcKQaMxbB2VBam+POrT+R+V+l0uV4v655GEtVUlJLrhb81
ss8Rp3w5avppZGFQFQPIvLdQ6tjSsxqkDeAfgjd3yAnBaEG1amwJf+zjTNsa
ODOWw5YMThyEwj6Vrk2icHvd532rZSbGEEuZJi+rZddAxOL1Nw39r+sbKGEb
w5bsCKe91OypKQDmD/wXBn711eFzzW2jJ6gJyrs/ireul7WwDiotHliFMNBQ
hvZcOy4CMNtI5gXgy5VeilKYsekAAXnICt9DrhCR3UZxu1fV+u0BtjK0/Hyl
8r8BibGCbOayr3PU40CJeVhhtJX9qRIyJVnNURQIKtGxkIhZ25L2g0nOW5yW
wP5Or7FfjvejzpsKdE9a8qTPCAg5Oq1i9AyDwBw7xFvmrqAuAbuWCEXLdZ48
F3P2UngEGUur9ZoI/sHlWxbOjINV0QAVZOmPVHo1nDoYSurVbomJXaeeN9D4
gPWEOSueQTZkXBncdo6X7j/k96EPTy8X94usTjHMjAltrjouUzPSfU2jnMkh
mF/0xonXHnQKqptqk0nxItDEFl749TjKlNQY5q1QRI3pkC8WwC1M5+ejuOWz
ib0B8pI0htJpvTcqDrNw8rBXGtjDVymkTepjWchV0/HophMRMUCjzHpA/S2K
ttQCO3HPbYpvgXGKe+QY/C3gszpDsQfR20t9C0G6YeC8lBHVOwVefcFaFxuT
YHQp3zBWfV6ZAxBj9+2gkYvcNn90nBubjHTnqhUw5ZK9+TQa7eDQ+gh7p2qJ
u4o+N5usK562BpzJrYZMsEASr0yi92nE15+sr3rLH3PRYyyBxgRSx39lzvvd
6pR2qKlnMto9/d28PR+pDcGYvxDlL4RCcig34BUaDy4MRitUcraNXsP+2mhJ
SY6aAS447feYF8Q4qzLnMzbsXU2hHonbf0IFB0IDAc7kZgnhL1rfwTNqsyXw
bMM6Q6V1SyEMsrJkxwtKRA95ckkVFm7aEZZQ60rACQO/zztFzxgNhSEMmwoE
iHCB9Di9hv/7ME4RN6Kqxm39Uxx/SDTJCRatnpBr/HYa5wJoUlV2CB00XJw2
SbG/3TqpN5jBucVARUKrsDz01OyVUgkXfRUwANCd+vVEOD5HMuZ169M98rb6
xEVG8UhvEMYSPDwi3yLha6itDsWHVvAWZSKq7DdrNHui/KhI9zom3J6K+mV0
MDtq6r3BSlaxuckEskLSE7/MGo458fcDMtSPF2dFY+j18aqTPBtcFP57d37n
CzhsUgKAttehLkEQd5+eTyW1GamxQcsXQtR43qhQFNmrWaLNZxy1fdVFYWUj
9+kTbVHVO1Tn+CwUIyLLVYVUK4/CRgB/rHl7tHvTI1QSJ5qJyyG0yzt5ImZ7
shp650CzpRv47e1U8tQQfhr+2gM+m/KS6EABFW38jenxWNbPa0VpinW9WR4P
z4M9ozYwRIZawbeawXPHJJeP3y8Mm21B4N0VCMFJUbRCNswLuISpaGi1Taeq
28WFWXXYjTmxuLyh6BYAoN3SGCjkXf40wKdUURBvCWS3t+cwKRkVi3BjaxY7
PMBGsL7afZ1o2M/rG2niDtETkzcPjG0yn2svr7BvJ8NCNRu3mvoi3ymA+qkI
zIDAEQY/0nYHIBYVtARV9C49VVX4OzTZi3X4gXhDxY40xKQjyGWa1zQb48Pn
gt1u+El+R/NxBwlpNiNY5WGJ0mm9p5AuxNwvmySHgY12lTFb5OwkwnTELyRK
Y1FBP8tvBM2dPh2ZMRhAKeos8eciWgbrwe3oCKmKo14V8dSHT4tNuW00ne/W
XvfVgjq0haycFQwG/KvdrQSAgHxEx8LdlSfhEvK3h9Cylsregxqq3gV5bC0S
KMnjttTOoZm348DHFs3CD3jq5VkoEZneyfaLW04FdowrPkyFa1TGU/h7Xtv5
sQEg5fV0A3j3FfWibjaqsZbln/5N+OyWIXIO8Ouf4cbQYWwws5aFldkPE/8X
6QDDqhBf6jSWr4+lBgIiAJ1Daw/88v7MCpRsnBRUhsj6+Y25khNrJD2K1fr7
kNG/vfUMa69tsulgYMLapvrdP+qIE+PsEpBwGtuU/bMKkbukxBV5cDNmuZux
1J02vuJYqM9lVYGsRtv7Iz4zYl73euwxvQ31jTEGIrKJ1HDok+IflqDAuwYt
DwSsDt2YTlwE6jxAnBRPPYJ4f2+KlGhGZmn0CoZ04hrXJ+tf1YWdLddBzhKO
3ir0JHdM6bwhCWThUQ9DeHpSpck3DpKp5uRkkpFOEHeilsd1tv+UaYp+NnV+
Lz9BhIVvkn3sN4uXS6Bj54T16BPZ5CVTyqTH4tEPhts4uBqQ6lNFgLYc+jMR
+9QFIIaaewKFaxf2QXUU0GJWuLS2O45qZm1kSewSpflvI3Hpk+upljGkVojc
vLBSo88xuTciYubIZsiZP9JYvyyK/kMQ/DnqLX6uuc4EX9fjGTJHOx0Wzk7A
xdCTel6KCKGBPzbnFCuYqxDxN/Eun8seJmRTayA0n/HQXgZw2b785NnnXaa6
HtTmq+a4gfRmJa3CM7MUztpSy3FefF2Kpd6IHo0gvmrOCHCpn4MznDpccWYP
gNyQq1z2Yw/43Abfgr0rbU4DXDvC+cV2OsV86CWqpqKms6mXe7YyXu65Po4+
4qDDk004aRkqq9IoNYtJemVBqNC2U46cYwFWIUxySDHgho1pJcLHoJUySJSD
fYk1FhImps72JsmNQcTKti+VBWgiIfA710rPon4ifjfpmreyO4liDwTMdhga
qe51hyucMSe5eudpWfdHERYhNrQ8p/wSRv35SNz/STlR8qH/szUNxFTxcFbq
XyjxVRTGVwbqf5J/6D7Yk6GarHbuf6Imw0HOjWAEMqYUWHzRzVdXQWNnzyXP
XGh8zvfvvIiSjML84w1Q+8zKLaeGbZ0fZORPa9yeOZQ9k3fHRNeP98q0yHq8
hZccLTtuNZqbbxzBBiX2v64FO6RP92y/9KMvYb1M+5f8jKk4hUWDxIz88rZ0
ccVZRXK5j8vHwkLG+vsBGaxX1KTRVNMHZTDqHBPZWufKJkhaqY1ys5BdeIja
Cew4uJHt4IhO65twLFn5sFWTMM42quVibBVUmdT+Xhc46TkupuNTZilTvCko
gEcNOUwTlh/Ss8sit2EHissQfWzAF+emlh6R/Yn8OU26rLShQD0IgvCVycLl
mtmDPTzp/lyLFBcaViMRl6DUKFp4Ggf6NoId/vqJjhGRmMBr6Kn4bzpNFE++
+t7v7oUIRS1HSQzc+QJsX2g+XDQebiBLswUiJbf3DZqHKBWL8J7xro1HCH4Q
guLlinYt261H0MXDcu1L3XTg0Zif8t6ZmYtKv1oO798g4VqdNJgCb7d6AkDO
h71dr6PGCApdphAdW5ol8ff6ICKfhJdYwj9JEr3wvf+z/icmXSqdEQEFIRCK
0GLgpzgXE5uW0oWpsEyI6sbfQmUF99976ivd/oP1LgRT7tF9gnHc1rjHuVUg
cs9RmpsU+lRiKnMCNux09r6s7TCjWwP7W/IjhNc1ULW8TsYMCIfdGdaCCYc8
KENE2VIiYhWJ3CxmmwwX/a8Y+B4glZzYLt2MKwCbbuWUYvk6VM4Z8ux5i3wD
hhKxpicu/ZtvYodQhTBkZzHLUXuHq0RQ17Tvel3jtUkKcP1jsJcsI+8I+N7d
REc31j+nr4th7PC/uKR9JSQ6TT2LbvAe2sahrOSC/evn5HRrE2db8ZMMtJNk
RKNa0iYoR6VIV1Xhcp/xD8+uXSXq7JkpG7+pfgbEsDUZhXnyEZtVN/Sh8axF
C7vlPbxnZlwr4chke2OBWJ1qmAXfPaXpv/5BU2HXX7IEQ5uTy3KS5bmN8XpG
WpCexwNCCFHvnr+e12p1TPzXLjTq+dnY71KMic319pPMMAriRy3kkHFvvWXC
zWl5faUS1z8d7LPjvG9krmA84HIDdCrcV2A2Yr0xn8VQHBzMpdgnx8S/VzaP
Z/alDu24IRscXsVMtD8Qzzkyv0p2HeR11jMhkd/SEPzYZXxIgGfJgkZSCVDb
U9edBPACfHEa8QsKElwljfhteEVwG8it57wFk0/iv4//9FfEoU6mPLKWCNaf
ta6yLOBBE3UWgAJ5QMocUIZhCi0kAVSviBlPAmOt2K9x/A8Y8oT8KjwrnM12
DPBrNArayz71oQ4Kl4RJjtuCxQEvCANle+cVfBz6TN4juosdXVYuMX43XgEe
pxRiyqZ1leZ9R3rSmcLvDiWrwx2geipzbRfFnesQqmjfA7rEBhmGCad014PX
zOVst+QuQZqIID9a0GkuHkG0nLO0UAHCFyole6B2f9l/Gq0pK1YnJDkzNQuT
dd2wmpNCEYLkK0okn76FCLbivP1hid+3+5t4B0HIGao4WnwASmyzyipgYfYO
lJuFNWP6x6alaPUlGJteR9VsHaumIt4jQ5dFibpQILc3761TgQU8xHkFNLrj
WjRsjeurIa7DjhVeQxLQ+1GwkooQZvmJiqlC91GdLzx5c2h8dZ9epRomIVzQ
sc3xhd3FidTTHxl+N26bL+hl/pmnAuYdd02jx1CUskJA8O0BoTgCXenJkbuj
MIdtAuSIHhVUm7+UPAvU5C9Prpvg/oJsHVH136+6wJOf3+aZNAk8Jfzf2iGK
e5+rFrWJAoHWK0XEKdtmhW4nC8DQcDMZNP9u15v3XOOF76qDjSNraUZCiexb
sJkoSxCtrkiAZCYM14eQMC6/4AFjRWEUWlmAYRnBWEf4hMj6yTuv+XReB/s7
J+IoJN/0YKKxr3ZlwZM9wnG2/zaFZpK6YGGQNNclZw3hIN91+nuKx3F4Enkd
hgwph1ftKzNPFbmaiikDcPQqQadK/YW0TWI+dlGKBXt0apB7JF7C1KfFjEVV
5jPtTkXw1usNSfH2p1uWII0nA7diKkzBZOMLK4/t+O2hSBZEEKfSlCNHUb9u
Ivz/79ptQHmYJmeJnvXh0E3Lwp3ylhGfciY2TaMwu5WS2RhqdM8Oxv5Vw35G
v/Mp7ubrm4rh+TQIXvVxJu2YyDEZ8Sxr5dHSgoc7U2XGmC69rpa+U+liTSsL
f2IULRqPul/HW1izjHaJNyhRfhfMZHd9b2e/BhWo7xZ+1JPun3aWyW1QQDxo
wrEAf3C2MTgugVjxb/uS/r4JnMbvBuGHuf/HLD8z/G6PSAgI3gJtviQptoW9
gDcOE8K2s5jWxG+xBjaux3CRM5J5xFilkjTauZ4pNGKaJacNNMUn3mZYfl4m
+aqM9wIGQ5Yfxb3paad8dbmVRM2WTAG8pB6/l0XXkCbKiy9wMTQjzIf86+cl
CZpfqcCF+j9kiAmQitcudpTWnYLoqbDIetX1jh1LatchVkV2qv/m8HHuMuqT
Oz2mCp5p1ISdTsJzTqdf5PE1chb1VDuGzYHs91DLQzhoj/puWe3avjI3A88H
hIIW7LHWaXYDPG4bB3d+5T0p2jPEZSKaeShC/sdXtWoLaRKFMYnqzdZ94O4E
qDBcU0tj4KNYmbCTEHX5Ka3Dw+v6N9y+hU3uK3C7mpsnHaoIzdUlnSaj014f
NCqWyTubxOzU/P1n+z1CHgxzOJG2i0lqp3vez485nWVjrztkyRnX237PRyzs
cmLH9YcmqQO+Ce1oBAZrm6trbCAZTt1nFBweWRyT6qNLnBLen6lsVpFh6xCP
cGqbgu6EJLnYsOILOv8YClSqchOwLUeM+zkI5oX+6qG7bfveaf7VgDN8TWnO
kHOYCmnr6FNM1v+OYNP+Uz9mQV6lgC4tbyCN7oT9Vk3Aim/asJF/Kk8U0DXW
Ia51oTQ8rA6EN2Wfn1MkHshGoiibOmoCDUarkIE9MoVgNSMueFdf/H16ddxN
4KT2QDNK2HcWo7Z6nBQ42PGaO8LEVS/s7uoLjz/9s9nsdWNCHHqSwiU+/Lrs
UyTFVRcrL3S5DK2Om0J4x6Ib2SPZIAd31JgFowT0kU5YsrXghtjw4gTBzc88
6EfUqzBa+4xbWAC/FcOQnSFSP2MDmA0itoE4ZJ1/jZ5Kjcjg1N7vwQu0w0z2
bV0XsIhk8EJMEghSTCLOSio9BK7eOxG5TyKmq/b4oZPWkl2DyYZrIWCLSCtm
sb50bjuXAgVh55kFWsUeYrVTlSHM5UOCpoA68FmWsVvKXkcMXwjixRIo0fFt
Is0G3mvnSIhhu82x6RrNali3N01LrIiwBDdAsttdYMzGcLlM/CHT1J/yS/ZW
5eEV0t8rj8KAmHu8oYTr8e7JqJUkY8D4sZH8TAc7Huu5qbc7mDuDXBv4OUQ5
XptyrdGHWebAL4FKZsw1dVzuBmuBn5mesqkYYWUGV+b4zCxWLHQEX7gitiZo
DAS16TxcO8Y/XhZGjhEALKTaqSZECXkk6I2VsexjfxfSZ7h/CLpYaNfs6Jup
fYWu8uf0qZnBSnAo8dlcMZ7bEH4BdW52gnKn+bdxP0ggt1vFAOvrg13ke63q
PeKc8ogDigP4/r6VCDQl6Kkb6Y4immE7GHH+g3vHt3PTQ+m+9rFhAOVHKAop
J8JO6t4c5ctphQkH7dn2XxIFZJw6UazTH3ialFyyKv/QEXqXzF3rMfc22wbZ
fmIRrsj5D+0EGSWKmRebOQdvV8Y09wwsYyOBtvvbTVPGyr7bSMyNxHrfWiRr
RoiMUaruFO1HJyG8472R/6LlJiT76cVBtVfY7FsjsizsPSFwwyE/5Ec1ABUC
qY2QjpGU7pqiI2GxB72MmqqEAt4slhPccf9d9l7KcZu5Hr9XIzBKrps9FSTf
SibKTLtaPU8NKkoKQ0AJezX2PLx04g1TYR88Tvn0YCZc0i4mgxN4Xa+v92qG
Xd0dd/ek9R/FCagiNMrwhVO/kj3WNuXKebtl/MdTYW+NfOqm+79mVWKf2ZxQ
92/f2/3OzcghuVtY8AUGDDVyVMO55u36+tYnamwJfAazpus8cdCKA9fWCpgs
+Sjorg1XQ/a6CX6C0F6FRJxtLmI//bDXSRJKnOtysCat3ORdCW9lsWVQyYeC
tOhSus7MLl/lo42DbO66fdZpWFfIjPVh904SqQWkgutgab434clafycTnsqL
NDbbILZLZoAoHPkYQYRAltl6aFHr/eObfVD5IgTuH0vHGjQ2y8/LhZj3WIOe
af69Iw/JKQFSikiNtgPSA9CXstiugN+5batlQv7MD9hW2fd90tJ4gWYw0c/s
U1MGkNGNq/s9j/j0NUWgueAqT/k/m919bP44pzg6DmbkG3IbhD1WDvWCgDLT
P1i4ZOsomVr/Dl3hA+hRzcUd4I4W1jWzO4dqc/WL7qiETqpQM0qiZnlN1x0b
2Vg6xN81WmdSlRH1/OZUmXrhRsRqR5W6CPXmw/2E9qRKSCZBHYx3wLca7MVK
42Yto33NmUgFlecNOPJ0GscZlDqV99r+s+w1Z9Jtf5MP9+w8/jkYERStXY91
q+ixyxU9eL4rcH4SE5tF9KG3b63ALZah/VhlhPK9I29fC+wY5veOPlcR22+5
MyI8otgL26yYkvlv6Mq2/AlVgFcckggn6BwTCzfC+cObMz3zGffpLu5vjFTS
t+xeUdFw3kTypyhq1VlFrEzoFTsd31CjKOvpxGUXtlJ98ZoHwMovGQLuizhd
LhTeMGcCH7u+dqHwiv/7D6MlXPecHrXcNiAmw5o1A7R22XtRpbRrpV/b3KAD
mpSffb3pfQauIuma941EZGjwfLNQOzvjgPkjBClNpFk7wvQw26UeJMCkXjlK
jPCOY8C/2ZK8IkcDVib0PkeZNnahnUu+Ib/Vnxv/syvnYgmV3FlaY02lC17W
gOrty2SwEU36o83JikZxUSIjogs9wfR5lOKx7x03pyJjNaLz2f26nsuwfpJ0
xGNiiMSA7fI4qdqJ5XFPJRtzDKN2bEMGUfKEIgaRa9Vp8i10GAiTENx6pkO9
RGidea4g7cmwsiyuG/YiQIw0TNRzqhcmAs+i5gIzxqdoO/h7swd0wIz4//ac
bzPMbpaoLADTZja93IGjIIvkZvkrkeUgaK6XSa9iAsC9edp9EByEqsn/2GMX
+TJOvxLU98ipMB4tdVwhvIa9rUmohuHiq0dmGPkMh4L9sSmyEh8Mx2+63bo3
LGSG/1BGkI97O2iv0N23OWuOXO5NyIG61zZUNio23ykGSZBqFc8gyDuGEwD0
mUR9JP9uLjzukGM6/D0zSTRoIaCbY4buTroEnGXZesX8KIu6X67E+6T7/1iL
OOoV3tTVYasNubSfI0ZJ8eiTDTHFPd3FT0iGfeFb6MQSaNaEWSmHtE19iYVM
LRo8ks6Wis+oemdt+MpOdf72UvcuPjNEDkc7+YoSpv6uAa1Bi4TzScV4e+4z
FlmZKIy+xheESLuHSxowQ15Y79FZB3RD0oPJcLp+yN3DONRSt2rgdUJKb/wR
zPKdNqv/mKw4fLiJEuCsUh8TuBz3oMZZ399TxrvNsVLL9IX360Q3uhSIeG4L
KJmv561JzRkHXhRabmB7eNuJBUQQaK0YI7mKLGOb8zzgDx21hkj655ugrDyZ
SFzJvwLhmg5HFWkV0xS016hGkDSg8j3Op3uV1vLSw/kgjAAReNhyIDX/PO7k
Zd7e7SNxxdpLhIyhX74pgriKjo9PdSuhBEvtxb/32cIa363bgAjk7/rfSkwV
ht0PobmXrWGl34YFTcUb5bUwni6JESlYLRLbfbanKxCbJmMOAx4Lx0d4IS/2
Q1cKOCmb3sBUS6kxQRtzEzDg74OTvW2DzkGQIiilKC1wbRhu/7+TwEQ3l/pX
zIM89TX6qmpEZTbVsFnIgk1C1Q1NO77/5hfqs/IQU2WxwEBxsaWFirrFkK3E
KHN3V5PHegiIn8VFh2dJK+zcuOFNAdTQzhOJ0wRvujsPcBMog6ZFwYZN6hKH
U7/pAbRNv0wgFhFk9oqDvW/zN3ZrAkCUnRDI/EmQk2EZ8h4Q64897QiG773X
Fw/Bt8U67Vcrj8DAaLj0cW0CDU5IfnFOJc8oolPdz7mqR3gFZAvOoaHdu1eH
YXwUGcF4mlfR34qi8bqj3SsVkQvfOx9hkucyEhLwAjMjFOzm5seC8hrK2jGY
1S6afgP4gfAku0a7bGAYvDRqHUQPCW4qcOzmha27pBsEvmlzPHm6MBur7d5d
PD2XdzrXNLOPq2Dok1Frm9eIAlgZe9zfHv9IMkgN10QyfTKvkbtBBdq9Ry/1
kA7EWGisSI//cq1Tihet4njGccvrgZgtdid1wxm/krDZ+ayI7xFXtTPGulXR
68qMlFmSXWbBGCP3dgCMgwwkWrotjmT3U0rwH21lNGou3P+5jt62/dQejPRb
OvsKbENl6HJ7qoviVF8ZlZh0fQgnfFKEZ3lhVkvodG2XJbOWuJG+jCM5dj/4
NuhptvchnpvE5miOKeA2mw+LNEC9eL7mFgd/CM3j6toB8VNevIEX9cQY5pk6
iUmzaWwLSMghrZVIovxiTMkeltgN57nf9236+xO/3CKMvUmce5XHm5KQJSn7
vRO2yzlCWFitqrAfwB02f2YvN/EICWyBUuhXJtuFQ07fj0rI4PZjCH3uvQjt
aXlRppSGGIcsQV9guiGujSpYq7y2g5MFdSMAg1912k4LO7kNmPLCoJk00HTO
n0UkgJfKd562eXqZAii9CC/pgMrG5hHlX13EATNYZoof70PkeJBbKtDdonRZ
tan+k1Vd3qw8bz/f+yfZ58G7Y3QrVqzy8iDa9yY3FhtXjvDgJVZtL2M+fe9j
tniaH7t7MeyFkGNqoUDLO2M9xUbBTeOup2z0nzdGNT/14ChLUiaXK89SD+Ie
izJE761/NtOIwd6yMmYP4HUSvwAlGhnvqlpRUc7g9HWLbw8TOzBlj31hbOZh
HJto7KrXAWLjX4dfbE2JN2q6DBkj7reCP+H5mXA+usptEzq2zj03CtnEN1+E
76hGoH7T+X71sF0CSTvw+u7dGQa89wmq9BtCl5dD2C7l+C4W+txClsjIdzwF
dyAgnxpYjyE67fuuDYx3TM7Jud6B+TZ1Nxd8+t4DhCUDpAvGW8QsOZ+a9VzB
5hgKvDSi4Kp3hEryiQlmdiRAIQeskFE9sI7k0IuW1f7ZPrpmsO5pVaWYayRH
I9VRcDV522WHuBgGp3COBy/0Sd2op4YIDU6mn1LuKLWus9GXU67xK57NFQCU
qZyuBn6jDbE2nL4/HEQuSgxzpjCsKine8HUhGw6sp3v8/iaptdE8kFIGKoz4
rbCs7YDGupvbYDmB97zTTVwYfn7NYyq8bPeQxETcthZf1ePQpwfig1qIEDqj
07QHKNXPA97yXq/2RA+l75XGQ45akWDYQNdxG3Lu2AoRL3Wd2D//Eijlwbhm
RhjJA3xG/Yh7t49KeqZ8FqiKdv+y+5M9KwSyEwk1z/I9uLDG5Vu9Vh7tD2SF
0DODDk4EZBOv+u58jGINqOi1jUwFyuQm7mzl8o8vNltUE9ghqE8ZW0yiUiNt
LP/wR5ETb3eta64OYmkLAkgh06SMlx7SKNXgm21w3VWrbjCP/ShYP52kZ8R/
qetQAV1wT3RC7Wy4Poudfsa81RQeGpGLmXDzP9Exbh6ob3GMN3WI/2y6wALn
uQztjGPKV9n2bfsKeUAXGmUWLRxowSkgD6KOQj/nQ8pUITLKKvKlCuTdwrDv
qWbwJOoIlUz3Rah9yn4BNnPM15GVSYBwi0e1Sl3ztK4gwQAI15U1okx9B/gu
uXr/Ffhkv8a/KWtf9Ppyhte2dk5rcblFc+y1iPFEqUT6gATRx9sGqAKPLXVQ
72EzDQxoPea7oVemYarhaePrGu6LRpAMoIj/08Bqd/4VxZp8byJBcY5ICLZu
6ZHdHs+2CFWd5/G3vHzrumqN8wy6/u2tjaVmh4bVRIR9Qn7q4KR9nLehygfq
/pAhMm9g+R6di6CU6Z6M6CHzan9YxoEqpGiibu20+X+Ji6ejOvmQpr8reSLP
2EuP44wi3V7/KtJ4QAoZ4AEstfekew0S3LJJA1PR0etcDe+wq78LdTNAEKxu
wJCXpMrWJArhfnw5x9rkpRdS6ChEcmGYDnK4Fl2nq/WgIGxDsEcQPCNPyG/i
JbqR2uSXCCGLA1K7cIcUBrCpSI1zLXwN+Zag/6yAt62eFNr+/VcWm0y9OlHj
MkC3Z6QmROg5nKU3CvH/DGU8em2ZCqHUYPVDApvt6DSaB0o87kJ2O3IZ79kA
Kbuxj8NodAoZj2I9UbkOTrHG+UXMH36nHpVpliXJ1hb9qMe04f74wIYQdHyO
0QfTb+bCC57++OcSnnq41dWJSOyb4jcVZECzLmzwUJtJ4DKoAzUT3tG6J6IC
mSNG8g860Y3RXNvi+Z2Sf/D+T9QcParE0ZnlorS9HsYlVG8YnPvxshIQDcbB
8vyHwc0oLXuyt6OMYddNITnDyA7/+SRjkXibOGYAgIVD+HmTET0nrRE8nBK/
VDtqkCOnIgPw0E0uEc5KvvxyrviwO25mbqI8TAl3LwMETa1ATYco8lLSUwZK
HPl4Aa8vBnIv5Lc6bRF9JW1wyy0oNLgKq4UAuajn3marZ5IBVYXI4SG1YSdk
Psr9AqoEt6DJWlnyVP8czemLN/5Kf7CJz8GV/IWamP7FP0jYJmU7SiPI51kW
p+paafKMPJyKoKvTcV4A2nOfx6p8I7sVghSn3V2/Zst/eM2y4dwWQBU3KQ/P
W9K1Z3spIOW50Jkti2Ko3iMfuP2Nuydqug7NB9CiyDgNsONOPm9omHYI4Cnh
9i+lcaw7OpwdXmQRd/RYaFyj7MLbV9Ake9KQKOcHNeNha77GUDeG9tr3D1qG
RPtB18Ur107S8bnjdi2QPE94dlY+uEr514wEtDBE+MznoW99ROzEf7kmWM8R
MSvckYzJkmGE4TEBFNal9y4yJcMcbR5LDsRSpuMN3BkKK/I8dUliySgWqy9g
xodwHtmj96nf0lLU/Lk+YtNcoVbH5CTSQe2abshW75NxeoY4dQFfqwOvmBrx
dCieWJXEtPIfH27VbGvBSE5cwDJTzLF2XbAxxtqwdp2Fk0kQApMf1rE7VFng
Yr6xMi5pBBJbgEgqf2JA8Slw2L8Sg80YFc1xvPh8HDB2Evt3kdigK5QTPCNQ
mgkUM/+/0dvBqDxsT1Ci3hY8QJFTk33C4okn9lOKSmhr+FbWqs9gxV+v1LYD
2kcDZWzLN/3ipMJWFqb3boQnuU7Mjydbs0yKXXmVOi1Id6pcPoTnxtKW33Gu
QJF+UBQdMaWFOvyovF9599RYB1CZE8J+b7xxIbq2/6uJ5c+/n9+IHHMtBbYz
3lueXu220mnghbYDZ+HqKvSS3L7r6Lfl2qYHtN0syijeFo0WWDfnsC/AUY8u
9MVewIh4uUXwMv0QWgYDRbWQia1xZpvEH2D2FQOd2XovuLqyJDtV4diLbMy7
AYPJWtQW8PNAE51/fmhCpwB/DyKlKVwuPLnIVbrHvotoMvnmY1oO+l5kv4PG
zwUymTtjILNTm/XjRTr45LHVJnHtb41LrRiHUsoz3F1q+FnZmqrnJGcEzv6y
BqHSt63J4RHTrXN3zgc16NnmtlpzBEJRGeRBB8jhdr9e5I58OMja/D7gqkmq
VwFv+YPcdBqcqScqBLPukkRloh3ny1skMeZhI9tbL59HkTU/xe/CPNnqdP5Y
mzoxcI1lLWmYbilqJr6diVtpES3772TQe95G1bcRNNGIXVQeg/IzHFilGIwk
LRqW+RVJz08Mwxgn0UQWSGXZZqHurb4Gp8rrmuG1UQWMf6J4rRq9zHY+t4W3
9pUY1TcF1kq6ZDYJeNvC585MlejPTOjnHDKyAALvspIF2dv1ovg5xflnKXgq
5ej2x+eTtl+fvcx71q/qMgk88lVJr73UN0dx/UAjePdro6bXUf587DPNjISS
5W7P2jXtnPCdWdUoUdsLrbmGJGxcMfZS8nbdx96pnOAaoccTcO23JvLeTfWI
7y3r0GR9BP0Y9p+W6Lvgyp30vBhaxmptYM7lzVCcy71IXOYuBbhdylp7itVp
oI2ixKwyRWiU2HoQtw9jSVj4gRx7eCFpM1NVJbiY63zwZSPC9QgEO2idDBxK
H5wRCVdQaBOBncfLNqdAkjPHZ601sDVMFUs4QXn108OyiJKBwKi0N2zKS23v
uWa/pRSj76jQihAZ6Wm++lpeRIZP/JPfWLyzRffLv4KdMBIG/4AQJziCF4mw
50hP3D/XjafYiKNDrtXH7a5BBp75uUBAiikJLYzF9q7nFP+1pJHmhbwJwq+S
V4GFSv9A+6/s2VeWdJIRaLIvp8O7jccZ5P5ZEkh7L0XPu1PrZ5eTpYqyF1h9
cxaoIVanjq4MwK6PUNUXTttEm1a+BFI8lB8GNdBWNQBxpG3W7/7WDzh13NbV
SNteyO9dVx4AplJ79BHh7dDTzLUIxohtWbQ/YTkMaykC04c9c7Xryn0SCVCi
qEbLAIg2gxiV1LZugTnn96tLojzuEdBzjlTLPqIe18S5Ebantw542FByj2nb
g83eJoAqGNuBuN6z4NeLcn1j0zHTPo+YFTYEEzaxA4+CaXAi+Uf8Aqiwpyp+
g0EV98V6t0BjWfzb+oZ6X51ILEKe93csjKmad4/+Zq7goArDUXW5FyIH0nBt
R0CyMbi+41bUGTlfLzovfzRRfeTagKrkRNVZFKimu1Si8z/nXeF9ysABb/z7
lb9JKeP5qN0VApPSKOqSN+P6f73H94ZMglGpB7u3zjDbcjq+qMc3rvP8vPvq
/PpUdoTrUjWIm0FnWMZwATGKJ86x5TOTDEKsn1KGidwEGbtaIJrrqno9dopp
W6beMGWO5f/a88uA2pSVTcBJxs5xjWwo8DJ14wEO/pvG0RQaraDgCWA/qXDd
jL2gnlH+qQrg/AkueeTUKCw+XLFOM6gL6m5ul5nxkH5wMtN6rhvpYIFhuk7I
OxYfVtupQXynw/MISbQObRvLnWCFT/KZGM+8Rn5QWLaLiSIOEnkC+0oPg/p9
avVfYhWnrvvJIpT/JBgjxC/4CA9ln1Sh73990alBPs47vAFNKvGgyirnRaXa
//uurQMTwzZen1IRsh0Q6fOhVREgoqKELTkKV59BPHVwDCwVKokU1xNtU4Vw
SFKSEVPcoc/keBWTdmRv6mgeNro1qMvvdCij0UpqJpZQCNnzqxQ59vfyfS06
zYLJEeWSJCSLhWRaRSEcGpPUXq8V10QfTgK+G4xVBOHQyNpHJ2BcScMguZJN
upB2Gwyl/kR4Yfrc1WYGN2JwaSjFiaCGKbi+Z3fNHJISKg5bFe8NqVv7TOtA
1CZhT0M600RsHc4BLudG6ma3M45fN1mxeTsz6L0/nJqVqtNpab45W9J4SE/M
TutAWVuNXSdLoWvYovasXeQbx/U8n1qOPj/dFYg/7+JnXzdJgAGt+WDWT84n
2k8GTUWQ9yHoa2F5D7IlSLyjUIWfSEWxkjqf+9NNMj5NyzSmDu2o/JBHAvB9
ysmEk/8DNI2l9BKKBAmqBT1ZPQR/0+awZyiEervaccXym4rUt4vWObOsmoMF
kvUQkXINmM03ivl0AcLKwKYbWbCG5GQSNdXm9q089ulw4/ThazCwbEH4MG1P
3ifZRYy7SPNpks/vJflm1ik4ofV0HWKjmCjPBhpnNhx+0tZWEuSe5OJQ+N4t
VPvP0tjVSmsKhp/NczZHhyaFksjMIJS8MLTWLe2/LjM6s3D+ejmk15adi5Bx
cWgNvHiGsgKqpRCsPhDej723iK3PxPvozSloXX9ftT4UdSR4qPQRqYDlc3Qk
IVoLduxnZpIVyF59spVOadP1RdkYf4Dl8I0AJ+VyYqaxBpSh3gHxqroeggyj
cK3wVmYfATPgpeOTqU2a1p2Y5cXZyw5egts2XHQYF4v2D3Nf/rHmw9CPE4Rq
JjewlirpRxSpN2b5Wi/TFTbpv8DMGO9mP8/vzPTHZ6tLipp3LuVJgwDY86sR
q/dKsqDf6MXt8YhsvrqaSapgN50DcGQLKhSDo8z/3lUYkx6CHOvWpViVuCpl
/LdCZbr4m3kEJe9J0yqZpHb33C5ME7L5lwbjq33dc3UkmM+/YIOdc0jIORJv
1yoUtQS6Um1WOX8ZkCVp58kGWfZD4bV5unKtlOnMvA6IbsP6HOyxVXA4Yqsf
dCTtm/D8wktFZE3jYhEx7WTjdxHNrclkpA7jH3w/68E8k7IlRpJtu953SKo3
KplhGpLHGokRgQvIK5tJVMhqZgup64E3d8rpm8HKPCd4mvsFkCB6NJJYrFN1
eDJ2L24SLDrjl3DBORVmm9FRoHIgTdwJXO3c/LuoSTZUyhIngeU3v3eyGLtP
iC0Gsdv2qEXa8DWRh4lEPise/02kHuqVxF5/ik3QsgxI3e9YAE6kAywgl/eB
WT+ngtnDlZkjzZjoiK0rDC4y64ozfjL8cC1jKvogemLT5QSAJJC7W/FU76ic
Gl6AwtSfcokDSb8zfbN32vvBX+at5jVLapJgq0a/YZ6hch6C+YpzslHP+QP8
FQGl8ZGn6s5w6S3rB63cdwASuvVFtmydsBKPSsNE7wUFfvUkAjdoMu5hgVQf
fOQJXfxQaxkhqOCI8UNJPLevJfvAKpDrmB76otfWtAI2EtYFGGrm00uGjqrY
MdKLLJdIvORJSll94nCVDWg4SVW7MAzZ58lPj4s4WSZWeK9hxo/opXRu9G7S
dleGOzOqbOcquCyHWp5DeubMKLHBrqUwdJ51vDgN7CbJ6G/NyEmKiPYnXJrC
hfQPj66VCbB1N9mKAxrryq2QhGWmOAk9Kf5FhlVAE1W1aZdeQ5+yP8FNMehQ
dOEvDrvQmUlNKkRCNL6rqmez6WkcQIqmSaWvnFxXoKTjDrA7cI5y4IvQHJ16
3uxcLmYq/HyUZiO5b/yULbAAIqpAj7C5z+C//W2w4CnMeWCSGXgiHmM6VX9A
hoIQjm9gBaaYTSSgZVw5bJte+ZrK1MRsvt3fvaBy/n64OS7vdsKIIN+mafgO
jiDqScptuWQqqe8+ULa83ENiwcaaQ39tbWybNK4dkB+pnVTunnwB8f8Qt87x
wItgF2tDqYvZEwOgAaPxgAOTObcH0AUFkxVFMGmMHQaHMwH1qWVntp71go24
aE3DHaS4EYenyZRyANcCG1xgg/tsMxftygbx+kgvY4OCma+uBInWV7j5mX5I
nTj3O12FAysEBXAoDQwpn24jhCkP4G4O4g7Def/2YiVtDHZZScLbh4rdYArf
UNfNYguunRe5my83JcIpaE9kCpLNM3zCNlQbedPibLLXbML3Z8W9tH/KHyls
RG7e78YJjDd7fMs5YECd2yJdV5b7oZRP6a+nKZjJ4eLMHqMjBO654dlJ+kHo
SFerLpX7B1GfjuUfD8hl9/u5bJZmVsepw06wTS1E3mKVgt/Ri1wyuJh+IXn9
/baZBTAFzhFoUv1adLo87eHnrBHRK8bnkGldnA0GH9PKhyl7yKS19NUWyLMg
u/wHGdr/CL0bCYZAu+BPpZX2zO+ljIey5UHCDB3WZ4BoU8xp4hyTdDLRYwx3
tiQ3g81TCuEULhPqV/jRZKHoE4vRlRt1XYqLFpnbS4kerccOhwE9CK9ERXD7
oo8u+Lu2JsIcXBT+I1OZMb/azSOkkGg1o9tvDUG0t744yXlhtQKqkb+55Y+N
Jl7WjC9H8FT2tniolM3nxkluSq5OyYDkqkCO3wM5tG92e8Uc2t9lbXHxI9oe
hAw6ulh6LTAhdBNuBKe7C71IGrSzYScGHCZehig2Xjsa5l3TKnN/oyMimFe6
OfwxFOUuy6XOsYc7SfI/b6ykknSaccWI7ZYdmgZHNR+59ZHVaMYWeDtnFrSw
g0fYvBiQFJmZM22g758GXtqA9dj5gRsuhR6Kou7gtLkqYeTKZPpm2qlDpjAn
q9ur92EN6dWRD/nf1UPwxgwx7hwQirX7BC0i9Z83cV9J7Wnl7GtTk/Wrs7kz
WttkDNSpxWSQKMohyXohp7cI1RwtEMHUXDFlNLpX3Y4zf/3xVgL3LKdNSxZw
A7rSQFR5tEiWUgr3nSI70u1e7oC1nVJMlXQIwg9/a/HX3W6kB+NYEnakcMWW
llDZ6JY7lgfcL9w+RR5u7D40IF7k0bbXsFETbw7+Am8QhsvTikdEuy8h2WXF
TeQYLx283Uk6i+0G7J7bOFXwj3U2kG/XI9r2ZkpOUGz40EI+zM/vn1z9Y2AO
745QIhFuL9lL4U7TBWhml0ZgNDi9OVXKyZz+eL+hUuUmHY9EZ+0i38T/HgQs
Vn04PFDH4WFyad8kw4vyDUO2Y1DejLuOqkFxGjc6u1dyxrPN1ZdpAxzPnndQ
m1ZkL4k6Pjw7EsLUWT5oobyll4j5F/BC7i24rUE1+JNvfodjBNhWV7gS5MvI
01mgD6qP7zD0m0NJmLjUssp3XqLKur/n3dxcWv5cvKzRpxGc0MujTcClpA/2
o/Ac2+kigZUVCOz90ziHQ7bWgvfvo70x+p7qno0QPfJ2AA5HXgYGOD5cC8gG
0YyXMxX3wwhA2tN8zj9Z4f+JxUZW+3ptj1iSIi1G2EgvhTmfQbAAOOd2azBu
YmBBR9GYcMUmx6rEDBbDwmTcJqjkBqla7a+r95cY3+bvrdfr8KIb7FomBg45
gyjjfDKgnzqWVeRs0TTA/SDVuchQn6VhB15ACht5t5bueGJ9KXFBOgKVZzT1
ve3l6UcJkjp8141C+q3Y5tjx5sQ4xiSZcmyOjZPU8cKw/n+k94hkf1ygPqkI
u6oWyEjv+0Dfdhk/GuV2U7aqwxLkEu1pguXA3JKH2UNWpZA4pmX5Mfd4Q8iQ
sZar6DpJKGBg/IbG+PGurZO4lDCzuUzmQUiqBPp1CGrcdKNJdtzNQkWsewaj
0vleA/6VtDxI+Ws4vwJXpOdno2TEhlHeQUTwB3gxuy0satCwj6ZaomLOtcwQ
FqGHx3vwRdOfLgdpZHDEuYdM8zdEE+aWvrS9ZX73+C05zG0xVHyC0EEIZNS2
um+i3SDXfTQrR85Uwese5YqaWTlpBkyFkiHF/bVIpnPs3gNsIxRp6XDBU6+P
DZxNm0qjdqEHXieJRyoU7Jn7UY9y7zM4IyRpS9q4ukGvL+tMfoiwPSyVXJIZ
EXWPj4O6AZFJYXxH62iDdruaLIq4YczazkgJQC5iJ90zOJKG1ICilo2cLcwD
mlZyPeLboS5a6ytjLcCLoeBhAv8L/1Zk2bflxMCw+NAznii5OgMoOFS/abTk
59O2QiOgpweOGrPzYTl+lt76GvqZchm0gBP4WuhUM9VRcIP/Y89Xw0hCXFdD
FLL3G6pzQIykk5yLSW+7Ra8MRWk/qsd1Mn5y8g/rphO2LtkP2u+QHPOcNFcP
eGrsb4vJNf/cBUeqEpf9OIv6F7w8m35BYP8TQGxgD++MdJPW761phEy5+Lj9
zMWahKnOlbVB5p6B6TTD1q/p1rZ84UB5kd6gZNevjRsl7qNMcT1BGJSjkwSv
n6KXTADJIFuCWqLhZ62huTy0KP86WGfNhs+3dUK3gxUO0w4jCRUnCK3FL6Ug
oSx9I7wKwdg/JRiQj4LOwAsRXQbreW9IABahNhN7HTOOo2M61CnjQJEm5tZu
DaI+Tb14Q34rT57EPi1qemGUsm2RO4rYQfH/iI00CW4d2DZEJ+rWb5zYmOkT
tNMBwjoJA6tFjPa9lk/Tg1kuJJjeFvBlwvfA1c6rq5J6JLKV0A9UyfW/9nPD
/VAvnNsgvJqW0XSYZKHo81D01w72S4wOYZZ6h5cKARTXKRay6Hcw9MP6m7LM
ugRsAJJVLxk0jjKWeu+4wnemm4W/GL+8HcI87xbmn5YpWn+S/ZRF5bO94tJh
OSJTYYY7190Xs0uqRnUO3lMAHG3CIYCzrlGmnCxpFdFani33NA+oVYOYgyKo
Czg0NPTGTaYw8GfuGKJob87gHftZNXOipBjxYkQ0EcKfKEejdNq/KadnRd6i
56hNL4kx/9YkiU1HXGsOhdWCVEKNlEp+bgSGL07pg3M7c7NQ+nqgX2XhCbCL
fp+deLClf31rHq2BDNrFkZRGVc9Q1Ipb5hGdGMQ0xA3brXtoU5jxewGafL80
is4knUl1boPyULN92PN6v2Y0AayCN25Sa8kwL8AzowtC51oRp/ebrTXpxL4T
vCQQ8A8gwwfHmXFbizstXIIgt0vA6fcTf99kic004l6K1J/X3qsx8vqDPELs
UTruMyi1TXp2vIzlEUvqhm9rCsxaxCOBvSHVgeAnWVhqmxcr+bihXJtvG43S
9kKVml317sZSCKYKgYKT3XC1byuL/XNCJQ4MARhitzNaKbQntNKrOwzgV8vH
GxyAjbnMWVJ84q52vhv0F0Iv+xkin5cs5o923mAtz0g7oe8oEdCVuGIko8Wc
MqDyud0iiscUBnyoSPg0AwnyJ4aSVnt1f2OYtzJdgmcbHq9WpeXD7AQUZtx6
Z4pi4z6Yl1xEkysna6BzlkPdd0HVvPm5XYsvVlM54I4/FbxQqrMxqXVuJYXr
gjVX+8T8hEsFg0In6oDLkQi9BA7zVunbbJXHfvajT7jXRKEHekFMB321K9bA
jGpNwYxnkzy/oQaJASqkXdJ8jyr46WtQ+CZHderMX7n+idTsmx+dfoMNDjRB
5UTHrwlkrKhGQ3nEffhbiyO2H1Bt6Uw8WiXuC2rbR2tjoXdn9g6NKNRb6qon
1R8VVXhSvTfEbfj+Er4sOog+4l75Rw0n7t3Ilw62cev27YtaG/CY+pAQ6Yvl
UV5PtF3my9Sg+SdL0xV0P2CC+ZT94iq5jcrBqeNZZAn/MDSNCr+OkZkHBmUb
Z2tvs/EJ3iXwtEyN13Ih5Ht6oA+OQEd42DA8x7u15Ta2IGWikSszv9YQhb4z
7HJaf+Zmjt0A4yivWLq7J2QjrrQrW9lWiJybE8JExVDqcuJ8+r6ffHxNDHFo
e0QVXw3nNxR0fwMcpOiRJ8WhP8+nTrADZDktEbFAL1Z2YxzeMaUQuT+nrpay
YI8lpY7mvSo3xmyAwoi+XRc4ZlwGgXRjF5QbOXen8xZ2ci4d3t1vP0CGErJM
Zh6qZBMuuE0o8BhMu7PS2UWMh/SA9WCBFntZgEWTU2WEcM/jHnoVOCgTn+XL
78kIduQp1Oq1gh5NbdH+IgsJwADKt4EEk0bVE1vsFH0DZeB/6wzxaxJrQzq5
V/0Z8VbOyAERxK1N6s83LID82BpgXzgSSrWHjHSWR0or7DzM56g3kc08RoxY
NaJWLC1Ybi9AWTM0HeH1g/FISJ1JjaQsaLd0z+kxnQ6hzlvqsywLk4E7kQ6v
7fsRWhCIQEVwS76ads+nyVAc3Ml/C4YWaEhco7sZD8pRGEdrFiLbYPaEkfUH
WVD+w+4KNmVh/OaMJZVL7lnCpn9+5Fib5p0raaopcnsNqf1Aydwn5/NYnmx2
PqmXWhvZvOOGNx9cbtkGY9zYgApLFDhEFH9vjwAAgUsM3GmHgq2z6s8F2IAI
NZUaC65I3KNss5yU6JkV/RdAjnXg6pxl3Om61s10W+00IbmYPbjh4LKah4Fl
khb+l+/HCilgIJNt23M8LaeCK0MasDYSuKoN91A8CbETM5iVSKYgg8QRpkWM
EZprlIpR+GQB2ZoGVG5swXPdF62vIgFh1uKdLhiK53S3l77BPUQjurXf8T/n
RIg9ER12h6z7/FZik03kfBLs2rXKd+pCBJRwkFLlbZ0EMVYzyszvIVgOM6//
0KnOFvRI2s+ooW89hMdzqojGoe0H2PcupMQ5ZEh4OyD11PzitQ+Cj5sIse30
5bMgteWVkPpf9DKPhv/1Y+cOwkrBNOMBtfOHEsM1Pa+nDG27Fwuo5vtuyGWT
RISenwGe5nZ8ddbcp+GpVDJDLcOqNehSjWSZjrKvnCKDPZoR605WABSx9c4X
1ZpU91tUTas3BolYurrP+SjNbxzR4ilPYZeTMbzdY4wygjcrx2dIaXHAPxfW
Lk6McH5tYEdVrqMgW5uiGMUAq7XK5K1bbpIiq6EorNaabP0p5D6L+qvEK8E2
M3GJrCt4Z6HGFc05VznaQ2zipbBW4psbWcGSSftHYuMFgrstM2vXFeUq7C5i
HW4+NcIPZi5O/k5z6LsUOjmd0Qi4erMScYDCCK7StTZTzTknYjDadA3GcP16
coymcbYkSFHh/6jTs52RYJhWgNFujpunnhjpY4EAaeZm5CptE9WkNpuVQMuD
meB+v1L8A+GeBy06GVchDC4vwWvOzeG44zixme52q8He4bS5vX0I3pK/imN/
7VLoAY5OO29gsz7sc3R3/cZ2zX9vGMt3LR6la/kl/jnSW4tVxJB/MCz/bfUx
MIW/ddnqpeKgs84+ArwbPJVdmlYUsUJ/o+67fewLCatHuVwvf5hEUfGNoHaE
9sgvX2iyiVdlBtAEQjQLQCgUJMYZ1Av7LRhjae00nLnx/3DQ4pizOUWVuNJf
Pqh20wY1XnA/8iP8GNTFhZQGdFayqSs4/h9GUSbmiBBAfWtm3n5FoESm/fkN
PDErcrmeDHaBKvWlibP+s+iDIRblOaaKXCmkpYxNvN4DCCGMPkuDTEw806B1
I1nHRxDLkJcz+7dCD0G1jcLB55ly/tL10GV728OacqpxuZzi14v70Jf+ijak
zoE6cwvRgXPmPKCkz0bemg7miT6/ikSNFAxttnFDqLJzDKtfXWuJgzSRz95d
GvmhWXARJGZqhqvgfJWnH/kqRK/WyieYkqHfkHrzz84w3omJ9iTE7W3XIuSF
SP/B5MJ5cpOo31sN2s7jgdKlhmnG22DkfXxnqkImKpAGf5A58hUuMiHGib/i
15XHKoz7ZCkgKQl4Av72PfBzFC5iESnZyQcOS10GqhAaLijyhY489Vy3pITn
j/XQtn2gAnlBs4685j5ULpqvmM21D+rbo4BwnZl4109IZ4QSBYnGXgxu1EPX
G9beyrGc90z3NLLQhedkN5sJAZw1RLmBPl5infstgPW7poHKlAOdWxL/XP/D
l7cYoFab7s5i6HHon6rV655h71ICUSCWSgSWbYTH/R5bnrYSr+I/s6+W+o7T
OlujptA8plgdRKxon9/NUUC5fK2L1MZcz9Q+AD0AfWyodGfnRU/Z+NPRFbAb
eW5iV69lNCFreANJskePh7+Fq9RNWr7VvtmPp0iQflV1ilgrKkE3xZm/P5pu
5ym8GPMhYx76aTJb8antFLi49yRXQjDQuTMBqglht0xQ1J/GMRm8U2Wqm3i2
IV/CO7Gr9TNz9DqUdi7JznXyoyFlQgct8TbTT5pH6+uksVxnu8gO1TDJh9Ro
FrwMMPZkU5W0jAUtvcL/+rPo6arFxZpID3rTXZNAtXn4zgp6/AWXc/cvIEC5
o0d0UbwEETOB0mENiZp5I8CQ3AuLS3bbE74l0FUiebCCXAGqT5f852/t6gvU
U5GRVrrf3Rpjjqn8sddopMepnyw1Axe2OBwGNhMQm6T1Qp8FJNKR6J78qwlM
TU8VExAogttlNK4YYTA3hs2iE1wDMKt+iJF6VO21+08b8KjGzWo4xaxgQSKg
kwm6QoZEKuQQg1JDxobj95ES8LdFJHqL70ysQiSYMKZwcPhG6NUHrOfdJGTe
2DIyasUhvlZXtMJYymcTahsaYAyxJ0/9SoQLQ+tWvtKhXzyGLrFA3BABuyLV
MuKYdmGODSgHmko9Qf7B54FFlSUCRsPZYIubGrYrUVHdcYHMkpa2yQbfDt7N
FMTyQAs/spEcW8t7t42zJoVlPWy97ZD65efncACYyFFOlHzc9+2GtdXWQhNm
Kh2PrCz4gYkAbMmEWLjQxJMZsmmmZSqwhbLN67E5U0EiIwcAl9ldAC5FMTtF
t9F7r3eQcHoB63BxeLxrIeAT+H6hoqLQInFJ2N5AfMW0wG7xzOjQeNv0iX5v
/+2LJ2ZdXM/Ab6EQbJgQEDLz7j9cyZjE9oQHwun8XLa7/rmhMr2vl4Mfj3bD
DYKaJb4y+B5BtNbufMnUcgDy/wy4uSRtt/UXgeULBwqUBHY2hX3knpjZnXcS
3L1P6OfQYTcst5PtjDAO4MgZ9gKCmtuCg1kuW7mNFq6qCRvUU30tIRWH/y/0
rXXlW31Zpo0fGDDUxE+TdS8TlmwFL+8tzbQDlgPFreUx6H49/astyeGZh/D9
DIReFnYnUhj6W3WKFaVsJOHzm/cLztadWsIiCligWWJh+8ErE8VlWEneLRr0
QwXHyK1N2ZOW++L3EjmNpMO6I0U1Njc/0BmvO5bukc7N6YHMkncxzCTa696a
NO3poGrvDE5o1723Akho+B7IGycdoyuECV/8HpemKZ2X8rHbp0FW/8ILFvlg
Y01iM0NUIPB3Bg2LwEgS8zd4P8bvXa9KxrOTQKZDcXh3/ApypPDRy9fCCrIi
rVd15F9iIP5mD/7CFx/JvV4URiZQ/vah1lBwdOgdKVxdwC+zonjAtRJUBZPv
9WfqhQM40Z1oYFfVAbckhIcOgOtef2+qkl7seN+FkZ4U9QXsdbEz+LfnoTQX
P3fpCTxbBLKmeXwQXCg7B5uN0crVsa9VWFFDvrhib45x3hTs7EaM55d30Iit
Qcxd4mnXRV6VdtSQfCsHQihkKXXjLj9r+sPWhRAsSbMKyYUieMOr4b9AXiAT
aJlhgS7pueJwKh63MSSOnv5Q5G7SyYbrIx5c+WNBIdeGKLkQAGOA5mm0792w
LnEEZG5sLNSB6lmv7Aat5WVDmNmETNdoz/sM9vBX2YOxcdDXirfhDv93SP9C
5AT+zAE4tuOCEa5dCQtBXaWqbboTEky80Tr1jeaXvp4rqcrWQuGGWDmL4G5r
amDJdLRH37TJbUA1IGbgIXy2oR+ej69AiKyAgovI8SeHZCh6DHEiriKyrSBv
A3OaTRjZtY56R750dTUUXbbMYGJoIKx5ZXbHWPUgqb6UbWiV+CNfUdYHD7Oe
18db8TsB12kkEnhnZuxZkf7UxCYU6b99UHFJ/DvT/jyvjohrZY4qV2u8Kc41
UkO+5C0M3VfjhD6LGjgJVjPTGcv0nOb9pMY8Pn4bolJ7hqE3deAzWwqR/z1D
tpclBztcina3HWekXc62m/rrYZlBZL8ZVvO0VQCuyXXzlvCDzPfC/vazeWTH
Dju/8KN7Z/a74Cq7u5piv1U4hn3UEKnyYqz6cUkhFFsU1d4zB+Y0/cAu4R8X
BzgYwOeGVJNBG554PViQPgUwQDCsGkCqph7Vf6AzGAT4bbFzZn5emjym6OLC
4K9cTmKArTwsPn9qCgcA4b6uHgUgMoO+UMpwDSDCxe1zaDZN/BJOpkO9Ewl8
ylTTRPHqI3WzGyBpW7XoFRdCMGDXHzk0/Mpthnaz2YK7lFKLrpY9Z2m8oC6D
tcSQdPTvufThg2P3ndTWx9W3Mhhwr5rbX3vXUz5UHm32FjoL/iRQd+k9Z/bq
4HyNcjdMnNW90c591CYjKDBTNKhTmVYm+OrV+N1FXvFro37AVcLTYyAXQ6UE
sw29FoGywSzf1A/AqCm8N7IxJLIRmQC5I8LCD+MzOVBbvSi96xkyHKZp5E8f
I0gbPSvZhDR/zxaBETHzEpeUw7/z5rXQAQaPnmdvgvPis9pcwUmw771HQnVa
3GdclspE+lGJGTlYJF07ruByuuXMQCG8XM2s3HHEMkIY/PeiaDOr2U/1gQ2c
sxyuRFXz+Trdjv1tUyfGYnPLKVBG9duvnurqi3IS2sf/0Aw5Ahd0agu8uY6j
evSQjgiETPobWZ79/d6U2flz+mOCguy5QwAiFM6iCL3+pCmvLI3hrwM9xy3G
bPaGfFMdFK+XWoYU5W8ub+YEvAjLshFrSinmMdXyTCo4ABsI5uI+QqY+TE29
1bg/cBaEWntBA3z2bVglSgXlGf6YAi51zhH43mDykDY+xNhjOkMYReXV0THW
UqiznHzkh60w/72E+vzFWGyVxsmtkpz5NsUjKu/ZolNqJ2EorgugLnDHYG+4
5/rYyv+CAp/EYD1SakLNwQ3n+tmfGsoGRubzdtQP7dE3lkSw/2ZYzb3BscS4
tMstHKeMyRt/sR9wtGsblSGutcFNWgnlxaf2XoT0k3QEh8CDBBZA/9R+D+p9
kzMK0gqI1uaIZz6xFEEqafT73Fy92cBoClcA8oEf3HIEoYlmKRgHHXH8hFQK
XvkJhocYEwchOVNiIlSuqCH8lE5cK/GYCd0DahDkDe07iTMouyXIsQaSTmfz
CHzZCypr5qQmDAgq0lh7eUZaCOKyUVPipomd83nDyX+yDnCI6iWOqG3dG1/a
MS7KbFtxi+x8R2aB4qXihXdsN83w6aJZTeaKe/FMGnTNdMZgDXvg7CCNC6KT
e6bFXyXXbfacrhQM7ABiwx3cvvS65sqBv38EWodWimGUmMP/xjf94D8a4JxI
NJCRsS7/O/0AvXAHMlY2daXznLhdlpWgl2uVoOGDytgZrKc9ynEU8mbCJER8
EoYIm9/Eb7UAiLKqPnq/Z1OkSObajm0xeNZL5wBwzm11xMhODGjv5R5RxZ3E
Ni1ooO7xrqFBdxswKpRteV0YPv1fLG8cvgMFmKY0S0ZMWVldYuYZHTAyYVPg
mRH/l3auVODb2CrZwTc4m6PzRQe435N1WRbz0FMM6bVMdqXDxEtf9g7FLxot
/DYfA3psPqGb660aQFcCPludnJcPh1FzYoLW2SbNVeSsS+l7njpvTdso/tZ6
gDBUs0EmqVeeAAnxllCAzw3sUiHxeMmiD9yppoHgYP90lycIcx8FWVHuTyei
z0/RyxSkwjWGQZJfethQBizzSjRG+NzL5XOOPTJQ7rBNvgnUE5zjPkVIjIIK
y+KSX5EzjB31wxbd3NttG+5q0i8bsgN6Qnr/NbyVHn8FkbUndmDnC4atfrvw
gIhuG4WXnjaOD1/x/gbvRCv3YJXsSAz13pcfJRTVtZJeo0hKYWTDJz4/ceEv
hl2z2ijN3ZeTgn3a61gcFfa6y6OBX+TtPh5NOx2RaO2BILRxfjuvtZpceYwJ
ITSUypNnOxZbavv94SP+wlh3V6S12+fCYeKyFsekg24N8gBQVnVWqLH5jUZF
nA4ZW9l9gqfTHPV8jiyucX24gztIIDkPXc2T1eX2krT0K32zwpgjMGLU+xv/
9Q/L/QZVw7CyiZlpo+SAIhOJXcp4QUQxBO9vFIupbVPU6luG1EGhAmnagIk7
Nq+Voo3S3FJ+AMjWvIFmU8tBoS4XxP/Ebfk+rMpNfv9FRw8AV0JKmDgb12bK
9ABXKUP+tAhC/xFUt7cey4Ve1VqTvNOQ7vUU5ksxMeDhLgPPDIEp/r7kGjEV
kNrcgGfeWJu6zLQh8MQKmyzRMQs8g5b2xHklddgaIwvqfSP3Q0qo7S6dlVQh
gPmVDhQHqgTwFDNl4xWiRFQYiN+vKXz8wb4R8alRcpQHnNQODSA7inxMPk4B
ubMC+K6QlZneR/WxDLnyim3x7J5udJtMFltC2//9mb5RvkH4XXpnV+brbsb6
PW1F23nM6yVzLlYMlZm6uMTxsEiJyL5iV1t7A/cFwDg+Spm5YnxCRQKxe9/B
Pq7bIFZFsavzfL8ZnjxyOLumU9z/yOczNZU6W+sAzE1SxoyRn6KxRdPn2a4W
5xnkv4WVSSVMMc3NvCQRyJG8AEcvf2CYz93LHrfpXw9WEq0g5qmu/SV6pM3d
r24BRBNsT5Ju8RHaUGwHOhpvNbm6tR9xRoACK4IKNi/WG7XegwbjAJq5hcV+
1gDDz/0ncZfgZcnt1BtJKkcMc+K6HuhKrBQtLOcXLzaZ5htjhhMkMZzgHM7I
D2/6/W8RO90Gx8D8xb7ggURoWP8IpIHrQicOF730OBev7hdQYPfFmzAd4rmB
0QUsvamJQZefcuw1zUlY2Vr2yFZqP4kxQdwh7EdgDEUSpskMbmIO4cEveMil
DxrqVqwxhZAm7/VVAczm0nce1nJIoYJqQHN8+sxJskLswZqEFmTNIfRcKmEK
jeGoSCaIdzYHZK3N06yM9eUW9Bhpsq3g16eiJ7qHwQSxgyT1MRJ/Ix/A2i2m
R1sSy+q+V0lX5ioc8UFdl2sNu+iUxv0Lr6If8EvfRruH+8b2D/PgjhZGPRU9
Bhqdwoezb0pcLZXL/WNBrXEv04PZLh9xzIM5+/P4smOALAvnTlLOfA3UbQLd
Flmh3M+WcZrEMT4mY3mAwI1q8oMF7VGf1dQdcKmcjxE1aRMUbs5cA4m+iJ+b
ysRuqJDik7uqE3CZuUT9Y4/CO7r6VpEHITfMOp3GR5iEDSSzuv3CTV3z47pU
STiwS7f+k8emUAm/OzKRHhUJSaCOtt6mi+xL1nBQX6MuhmgMP++eTuwel952
wsY4UPC4Cp6NaudoJAVUJaCS6yXop0bgULD4tIVQjJbK2LylDboJ1vbCjtA5
M2BhjuB6bd7TPw96uacVzYZ+KZCNaZ2+hKjG5j+hM3H2AxM+UDMGokOgHpSD
mHghZ+PQ9HF3Tb9NIgQ+IwNoH3oSEIac2rbCAXNcavt+Jc7ghMbxxTrr8T7o
lly/lmDNQtt/cw+Vs7WXoZUQQ/iNftyUztVNkvSfOdbDiRtwl5iJpZcscIHv
YN9qXVF3Ott8CqgcnbzxsfJu+qZHflelbNgahGQhpvQrK9ODoKhX7u+9maTy
35aekKlgMVLkTDyoJvzgPPE/GBr6zzxoP7KRtw69OGAZXZ+rR2x0A97opApN
lkFJr5b4dBgJsW/RKA+w9qU2FF0XZJyX6dZC8JFQuFmQTGctcuB6ovG8cF9w
Ou2p52XKfOATEZ0Ly26fVXDc9o86pNpTTI4KIjMRcPTkaf5EzwCcqySNTcQs
Nu2qasvwJolKUmE6tgubofKG6zaGVYTKlThTkJWuECTFAZy5qQgIjujAe4lo
tf85uyn/d5J9WyBfIlHkjWvF/T3dvYMdIf8iPgrdv0AUSsNQ6aWzsVVU3wGE
5RLTnBlvV6dG9k6WU9d6WPvo9YeRuBwHpd0KH/jK29gokoISZPPouFefvo2W
sg72LUgB+BCwVRpxKWZXeYSxLM/OmyDNzyg0/MnNNLlTZPf9L3QmlWkLAuNA
YMib0mOCWbF59OgdH5tadScT9IUdUF+o36ll0vTFLab8AUQDSnko1fz6B3Oa
JNuweACSa9L4CT9rKlyBZgZz1GdKyJLDs8SAyfYZmV+YYJd8I45r8B7XMQey
XWrCMnhr2nBwmOkjxpXtppVlrm5+1iBgJP5mC29C/G7AdDZDGIFZI6WHkDRl
lOJZLuidCe7g5SksLFvqISl2/Q+hOX8ARYulhTvYluMI7R2O3SmXAjeBkea4
2IKSePb/dNxKVLaKjB0dcX7w9Tllu4eVHYzzWkS2wvH3Ho+GTnVJQd3CHjg0
dVMi8i/JlKDZf6b+bxzj9L5SjLdeQ2R56IMqmkDqKi6oxZXQT4N0pYrCb3aZ
liPJmLaM1YDRNwrzmA9HfLooVuqEm+sUwfVKwUuBUb11NAmhGXjhfFQ1Xxs6
asbgIduHybLWxBtdDq4U/Dxlx9a7MWMzrjemPI1rsW46rP6CI8uC7GMMSGpp
urAWJeUsYI8cLKPKvibVVvxwrJNYLz8JWYVioMhQEckkGYGiod7AY65RpptS
7MnRf6U8uwMuFEBZYgGeYUVJtW5uJ8+jNUN777v+zll67RKN5ffUWOmElE3C
rk+fiag+Vb31oQoOy/J6h2L+uirqwcdU7HeC792iKKD8auz5pCGOYfuhsENH
1tqbCTlvH42kJk6oDprLPBsVdnhoSNQiJlRxV7dyEx9OALprvqEG66ih8l+V
ciHHf/vhnbXQKryjvqqjMVgtFMgPTdrhBsPONrhsZd0BdUfR8Kf8Y3G1RY6J
ee3edENrW1HZkU18I37duLT71ZC2gembTadmQSCLjZhbdl/YeQ6PQ3T1ISOK
LI6Z/GgUcf7lnDKS4BUWV5xj+Xv4ZclBQDz9WRHVREgJoZmJ+0OZV+AhOFtL
rxfpiRRgp3Qj+ng3mANrWCBgJsLNVxbQMqlDoXFYTvcVFz5E7+tjWYhmaeDM
WPBjVlCZL6mfz5ccuQIdxs19NoMuoH0/YQTUfNt2j4fIfdk0fClWNn0KQ3ih
DCN0v4wBHiE3KHcmFsz+fN+Rc19/8Fup8dKfRuiKkG5BTL/fnFrDJXy0KayL
DFHFenn1mRIAZer1jOGKYeynOYQGKjaqm9AEVK+ia0RCqVQ9bHGI60NwXelb
X6pcdiRT8lXOYQPAOpk58+zKrtUPXvnG8lp4FNuM7jvJhmwgRPkldTS3Qyjf
GN3f4dcIuKXR6ut0UQoMzvYRnVvHg6HdsUvuji8LvInvoKKcVETQVHgifOcp
W8u6XyhUNTIK6HsvWxg5gKTr/AYG1r4iAsk113ltanfTQkU40oCe1FsJpgE5
a5csoCD25tp4r3TZP/UQAvG+/qBZ6Q2olWIMX3zlTUrzhwMB4eRxkm1DnA5c
C8ixiIO3zw6RkCbQo1rTJW7tlCfUdrP/Yzzm3y63pAnexTPHgSrtfkSFRH4y
rFkqlZSTu9Ix0M1X1DqpeKf4/aND/YrtdAHDNTs81AhYolshWmXTrZ2R8H6/
URr6KW+d6oh+HCzZsKJD5zf/Qh61/6QWCRipDGaSbVeBedwKs0RQ5A8zsNS3
Dt7TaczTkHfstzsu5zYpeh56ztXnWux5LCA4pi0Eh3gLO2JuqBdmzMNv4Cvo
wyxz7TtW+glMIQORaALIDiVEO7coAFSmj3UMSQQBq3tInKalo/bXuUWDKTBQ
aOl6qWqlf9HBY0D6A9FwswfnFvPGtJOrrb2l+82j846Eq7tlvogLOIxX21Y0
xasFGbtbD06AYZy2HhZVCv9JdJAZTpX1mp2hgp7xGWptkz6WulfdGVDC3p/6
EYl4XEZx+2H4diahHDoWiKwCE1DUR5S1+06RAayIDOPcrQU7qWFFBVI1fEIa
gFhTESRlsTvHt3oK8/eRrmMzuxLMxi0ZjIKUkLvH4XA0AENQUIu++ZH/CBZN
kScFok/zfQOCPFBgS5mEMYr7wiytDaXNnLe9JbokZkjZnoLy2H0eIvfoUKmA
9sD9a8tYrwT9NV4UkKMyTEhTSJDHI+9AQ5GG07UP2Gj2vNOe9LCv9kYabkZ2
F2xoE9oV3mYa30F0Rhm3M0dxLlC3sX+4QVPczu1acJHQjfkVyChJQF4Re/7M
LDOWbJF0nABMvRVM8rx4Hy2j+Vv/S8GG3R3287NU57QoRCTXUWT/N18uyraf
nWhrcrii/QFWZA3aDeu+/So3oHYWtCKJhcgT6rda3yauU9CRefbqsiMolwk0
nRIYyTApX/JqVHDtWiBFphkG6xsqe5+UHr/CcEzeFNyDkIukPc4tA7FaQCvq
tE4+LAnn4WKTWuOhDq1jE0fWgcRd/z1VEq7jDFqDYIJy6xk6xURMJVslG5A8
qTCoMP9GxhL06+YRVDqNu1+gXuUceNk+Tx2OEQGRAX3UNL1l20oGV3OVpJUn
TOVeISc6q/KnIz9lJlBLVLOml/j046RQ7vAaq8fGBY8JNGL3x5dnSgzhZol3
ib6PUGvGvUfln9wAAYHEELF1F61xjEQBP0hAK+p62vSLwH+DiFYvfSBc8gGr
Bw7/vUdkIUD97WngI2VuLJj/mtcEO5HBQif2k/9QXNmn9m9bWaXe+ZJjoEuu
E1lmZqlQcJjffdD62R5OJ68vp3zMGnzSXOIjbMX7dTDR1YVveDfLLkr8M6TW
aSS9xoicVawk2lTd3R9f/isUM2WrXwGtiiws4DgMQPjN3MQg2OUi0vInLO2y
kK9gHt0rRKhQbgFsylUB9ZlI3zBTr0DVCbd23YsJU/Q0PiNVF9f/Wjt0f/7a
TVK2TfQsfLKcfyLjkCw+ai6C/SHZXUdvObQ2RVK60UHjc/MWdkErqmOIgC+c
S2N7jqRayd2YD5XM2Aft2/zFs6a8d4Cp4XJJ7OHqricPlD9dmwR4N+ymxjCx
Wt88DcvC+NfFK10P8XW0PZdDrbqWciqP/zZe+zgYTomQFbxOsWKM7vWMiYMM
q4FLekuD+BjFzHs0nOadv5nAgs2Y59oJ3knsTpwdHG+LYWzsT96EWAZXYK0Q
J2CqjXb4PhyWCL5yNSm0OulayuD2QG+dTFnSgMWtlhfGbV2lcUDexePRPlii
MTf0klBB8QV2NMVyxhHlRYBc/FceGV1GWx+qzxVG03cSEYziSVKVk0cYReYU
N+sPDPYg6sbnPDUOdecBA2cDuOy0FWcNsVvRGJKJBHwfGVqGQx+EdvWqWm+Y
RquATVSaECy3dw3yW0aAlvhTiEKSYdMEaHFzJcXhC63zkteUDujLIzyUB9ae
gj7l/MPSxqFGIee+nS8BcqY/D9b3F3vWBEsOAFsu3iIYJZ/P8uep/zovCogz
w1EMvOOvyRK5pA7gTqhT+/oR0AKSv9+hBbMZ0Oa3yrWCm35FF8cWdsI/eINU
07o0uT8mSUHdRZZR4Lf8G/FfRRe0wjopjq23z+NBUZQ7vqaV5DsICQ1Fll2y
u11WD16+o0caenDdbnWB/hdcyrHjjZ853hPujL8U1WTPND9eKmtIU1GjRgIF
TATWuxGZG37uB/bHh9VNcOUhr9s1OxT/qE/+q1hjgPGYvar6kxVlnuhBdXIw
W1nILA9y61ZvOQYV+9GVhgzrYxFUoii4/CQwP9nj7OFDYjlukTVjoWgGz2N9
XwDeZ6PNSZU3Q3R0D/7IiXQ/PYXmp08IhsmzaDDWkBh0XkYwpIS5rh4F6ZGT
LO8iHAp9p4FjZ3feq10QGJNPTJJwkkDjF4c2GCKoqsg/ADLeB+R3btH3bGf3
PnmL1j3Q1DSyHPvprLqYvZc6qGCigFY2mXLJXByRrkqmRipU97cNFL2fbLz3
NnRjIblPMJ0I3gkpLOC5Ez/LIv/eDPYZ8U0tsxOCtuUuYVAuaqsJolLVjbgO
Bm5oZlbXXheTOi8YIjUC7oS5a9S+xxsXYl/UCEC88a5DyCc8m16Vv6gbvqfo
d+OT0i15/h8TbN87V1KyHk5pZMPM2WDaONisHugZphH9vFZFKzgT6WiB+uBk
CNzYojmT/+3GOREyzauarvcBCig+uhZf3VVHZEqrXbrEi87qTD1CogEPsUx4
Ua65nc6iuZPRx5Tw2CmDFw4bP7SG5M8q5FZsLvdunN+sFcQhasPJi2yc4JFv
pgl25szqYrFgbkpJMYTN8Ts63ikLw1oM/GGgZJMTsZxkcvLrCp5hBEn7gxNm
vKmsLM/kehxw3H/wWNWq0rCXM7cTLPeW3S3gaRVxtCHCgzJN3ZTLPBmcNeze
pLGdMJPng1CPuJebcSm65wYaEs8bvJzog6bQOAFQl9a+7uABfgHL6A6LshAl
v72+jR+05SFfvI8NfGExTztSwjOZmAMmNxOZf9z3uM93IKkhCUlpfatxojnm
uZ2+xMU4QtV5wlk4hxgJzQPBplwQflA2gecN3GwwKrkibxVn6XgTbzOkYDjl
icNhW2PIn4N6tAwM4OlIyN108JwH4j85hlAcmEleLn75j6fY2Iu1WOph/iJQ
AIuvWZCPIWrp2k9VhgPUVUcJokJhAg4zWnPnGCBxaqm0rduB5bNTu5KxruTE
nAHNqn/qnCKSxvZAiXApIsycjpcWKiICRaN7Jcrx5cR+4s9LfYo41LNnzxSl
i+U1m7qO6tXrvl3JgKhgPcWPMmhxRXHtZ1f3y9C8aOprhWU5CLANVXnj5Pdc
krWl+Hd+jeqVOhKnheWTzhitcqEseIcdFb/RbvcKWiwBLVrQa0GtNGdZvD0P
IZU+3FOR4hWZ/4nrGOanTqJ3iv4QO9ZcmR5HgusAZaaZ6mEETYYKG4TthROR
HnnhgXxvdLCYk02+QpBPzI3v05iPgkUUSXiCuL3in5YtXzqqUphTjSHMbOTu
eTQoLel0SoA1Qm25Qlq6b7LI3hVbci6O8czqEHlId6IcjGvXRUfp/5Gq+Kad
3LavaY0FmPppXUqLtWhr8EX5r0X0D3MwIfVpdQGtU2W6fLMNfZ20sCJ0D85c
jzdibSV7/NQQFtGN+Fzma89G5OxJbnKTFORE9whSwG3+7TjFmtiS2IWdS2ae
8brfjGBhIgnuwhNk1xzGaT7HLD+P+qzz9dU7UY8czeAGEUFV6/6GjsbEcq/S
hU0BZUqLOZtrvPf/r4rCU8+WqvIICbaNc+fMlZVtUEpCz5FhhI974q836uGf
GrUQS2mf2HI6d0c1JI2Lqy6/2mmSi0GMhBMTN6vjk0scpqfn9ES+8uUMyOq5
rQ6gsKncOEm5thsnPk+vKWWpytU14fcJI4Jls9vCls3iDZ8/vu3vQJAMJto4
31tY57B3OwdaP9955bhy4ehqp0Ex5XUDkNcc6sYPkLIT4nHPt8PUpMSkw37c
KrBNVSKKq0aNUZCutNVtNsVxZDcGLxtXj+WsG1bZDzHAkbvms/PfSipw3HCr
o2N1r0LBcrkHfVsWDrOovm+TWip403nPHUBJ+xwKQTUR49B6ImUITuK60sfv
Cx/Sp3G64bELUozKASPp9QKTugUUTqaZZEcCAxL92i7JUIuJDx/TIvDa+BTa
+cWB08WZGkMDMa43k4Ae92+7ttD1p7XAcsoEss/Wu4cicRSx2fog7eF8k0HC
kWjA7gXnGYh8mdGfZTkUMnLe89WFwFPRKwix/ehw4ZUf0TeSae5kXXvA8QEv
bmrfgM2PItb82du0c+wIuTCGea65lsie+JNbzzhPZc2qvbjqPA7Sz1QAzg/7
bqvb86ms85OZa+t4nh/5Yd2zZ1+lng6JAVbRyO9ScsRPMd/4S7ZeYbyu8bo0
aA8lptx8PvDE6qYYnKYZZMoG/nq8rWVtJualmy1GaURVJMkGwz+9cky/21Bn
+PIo5fW0beCFn3zOAmB5dvkUqikjm1cnZ/uHyuAut0sG0UJwuncmf0rRLlyE
xgdTUOyM7HDNqmOhnOzjCCndvJPOFGTyTUe7uvrVMzztHqVG64fdU15p618t
DrCRyNHmL8U24xBrCh22wkcc2eRrXdpOz8slKWZlj0DGrm/QwC3uHxejdxmc
nhtODYT98gNkaxZkMKtBIGCYgLCO9dCb8PR8VCic1fHdNAVnYMK3arqrTBEw
7rfJyeZQXXQzaxcEwH2/bxTymk0NZPiJX9Rwsp1+Jl8q7bH4YKCROuap1ay+
HNy4X8XyA+AYrlZyiPD91mr39BUd03CRgVHuyr9ve5gqucmGJFVZDqYdpKzx
9cGaIbpYDaO6FwzUsWTzu9IVL3Fqje85LVlA9m/K7f6XeiPxEe3f35vPiURq
s99CnK322g4OYL+vadXQjG+npsnEG3eECnH6kRHKUe4dpPdoFIeN5oJD0eoT
/1r8sI4srAVUrQKY4ELBjoToQfWeSotQ2dPQbaasRU6Tw9B0aGIh1PkardBS
kmms5E3S935Yj1LzNLj2y+UcYVkOcOXc4lt4Nt3p0KvR+ZZglyd2r0l+j/K0
7lCkq5OUBvv7067gNRnNDIU1yZ8+QRVjCE6xHfKkIz+QAayCfseZEXCw+MAT
6Hf5TYG4VxMUv55jU7wBupouIu5wUrTKR94mSto5HhWxN2u7s90/hhsEwKfP
ia5qjKLjJ5Y+BS+16QikzNV731Nh4VgPvfrO0XG+H7PpUyxwkL0srEN9i5Re
wZGYJkMqw4alvadJSfB0PVo0FaIzw6CWdF5G4vZnLWsHtUXwV1yrkJGOuyfj
P2PRoUn/Dw9y+2wbZ9dvTgfX05ORNn6MR5VZgoErdDmmZqKMmAHJiS9Zkw8t
MobTfmBixvxF1DXBVn7+Z0lfYh4kLUpXT2cIoWnA2sdo2PqyUElqzUQQ7EGD
Id0vZSja90yakz7+C0l9p3nYsFqCw4clLTZtH0QNUp3CatgaUdf/pHw4Xely
Q5ssCxZS8miIEM0HTEPGlNALsxFUj/LOLkLs2kuqdimYEemdBW7ensdAOYgz
xLfdZz4RHIRC2tttbjB+HqapqFTb6oWAZ+K1mQiaMGgVQb3osLco8daEM40v
6lDRPHsy4Rb8tqMZtn9ZKWdJvBJbbcePVtyzPznoJTw3A6dn0aSmA6BpHtCe
hYR/6orOPSY4AiDLKlzwwK0bHq4gu/mbeonO1VVUajhJEjWSWJ8Gk6EYOuGg
csKDuno34OK76dqN5VXYxbFivrS8Ng5F1Q47UtcZEeBxWcxqP9Oc+7DXJyii
GZY7+fBUwXgTUNIc+ehKRIFqEHqpkyLGxeZDLWKs3qwWFMXyU47s4q+JraGJ
MmhNmzwPEX6Z58Jz8eAxrNNveHpiht/2weQe7TShkbbs2/NME8I8ekD4NTbR
cu4KCbxd4L7MQ3iG2hz8sPuKrRIvzcpNzn0toFP0dODAYwbW39FVBPunMlMl
KvMHkZFgd8cbikw9pMhL7HE27FXYNlBv9TtEUfzUYCntdhg7qvhqSMNTeBhs
j9JL1li5usNhAXj605bI0ZmbbAsKi1qjRXdeLpQ20apQYrloqtPBGSPtw4Sd
gFkVt5tkRTqlpADPCceGwyR0iRfEtPiEAtj8LK2gy2MrOEy84clIutEynXgf
JvkWY/9OMXmrIrggWJbWzpwPGnAbF/MvOhP/SpSctQZOotPv0ffgDRWbn5RZ
NJx8yq5isoIFn1PtqmUmFAXwmI8U6/LYvjmdDFJHGviCeZmq8c/haJXMZwqK
N/iGrvZmjeNTNmkOslPfR8e8DkGXur7/t5XsInrC7xKqvd7Lvk3lcSR/FSOo
/PDG9dQ0eYBfeg+Ln2p4P6jhlbhs7aSQYkt/4+fx5BW0E+p6FBvAkJcjsLpC
iiiaLQXCNL76dtldlu6TDlNXULqqav4DHOhdmKnqEMCwWAbHMutPirhtrkrF
OKUFj9LO016c+EgLZcGiSs4iC0K2utMq+qlz46JWnKf6j7VJoCWh3F11W+yS
MCyv/h3dT4XLjdNqjQKUBYUheuRh8sIUD5WQYJMY7DM8pXn8zMci2UWiDMf5
6NKLE/5sAAT6pDE7Um/n1Ah59e4zQfXZZdwwkXo+/lxl1+c+zZU25byTJ07o
+k9dtNRGdH8PqHBI97DfaCnFD5pC3gbOjfaQ8+rC2AHrum3tBsQ2JQPWtIt2
qjkky3TJkThW3etY4Qs8ODV5MBP1ucG806Q3zBxmrYPyl2U+UmYSj9suYJ1+
XEIHGhHf2pYNxXJTuQrnjxoci4sDVLLb2Ob5FJpYURNLYJ7H/3FDMbuQXqQI
xkG/nM0MflWznc9J7lS/e43nrLqISFtf7LTwPSRATv6pQQ369c5WOHDcxub7
Y54hm5fEuGLB5yWNAnctbow4iFAgvyhcXX3iaTtlfjFaToHZ3zHtzuhp05At
leg+D3HVtHFHrI3yQBZgHmuwQpQowWZFtDFPckMw0OJ2M9QQYa89+dxh5ESw
RiEWPS/iriJElMsz2JQ2MkiRt4L366bQ+DhRqv/7IjiP3vYXkf0xloIemlaA
t6oSgelZIeAVrzrau3kz/3RgKJFdVsob0D2WqDNaOBvxbuXfri5J85M5aFDP
j4aMa615/yewJNhnN8atO0WFeqHtp4filplD5CAV6RbJqYJra73psRvDCHIX
qTrkpNvrbNSytZ/yGqZ5CxRrrfqsbbk37RY0g0dbgQwzjMDBPNHcudKT5oxH
zSJkSdEOHeUJV9ePwOup+NSlVrS0bbGkm2CHBuoHkBykDO4Txwc9wooSe+Ey
Q5SVX5jgoWlRe6kGQB0v77sJInTn4a1OAh8fvYH/oRTlAsECp1hic7HybD01
v8ZWR9K61Fw05p7ZvwUfcUxRmB/encRad9Z+ls5RWm8Hcx6ehopu3LT/rEIH
s4XedHzlgOVhRP5BaoOGHGetAe1x9R7JMCRXP2pG2KRvY22ZDIzz8t6WuV1M
TrvG5yHH9niSFD6n2+58gEC0jtGIgUQk6yIpeWTNw5HX20bu4OmBz0H2Kyfm
DtB7W/qhQgEzfZOmJQa8cDJD9XJ4/CpUX32FDiduVPp/7g1a+2VqaBUmeY1w
n5aSeGWuIvUxwbYwNTCm2/NLAMqabDqaPiaMGJqLAJh6LFmqSsjch/B6IZEs
Ut6jLFCN3RKnUHJvVIS42JC86+xpdtCrOvEwDZ+MEbo/qdLRIeWwRDdtt2d9
lrnlLxnc154rrC480ilNSDQ6SqeLZ/rQAMLCHoHX3wCKboPcOGBaGsWFkHno
ZzAqO2TCoQAGpEnIC+GGVonku23Gd7tZmPN3SCABcUhEan3IbVKLz72Djf0B
Q3VKo6S9dx67GeGJR1oJRKeEf2BTzQq+svHhStyaOSMxC7IeGq1lMShZ1uXV
D+Djl3sy+xMRg9hMZ9I2cPJ7xjwymFOLgep9yV3d8q0fbmt3lhwmtqP3hy+5
VZHRIjp/4orf61LJP82n4wtjETLXT9h/fNOpjEaxPUjnAuXekUaym1prfDWg
32kzfwT7k+vUC0mMPQ+WVtgW4z4wkLlhjJenH41l3ihcWlRVLJaqN4cM3vVM
5p+cNq5svZqLQv21ea6o41DChrM+EHyjLFxOYAhLdMKpsZ8qW21qI6wIOe5H
XacWcjjOeBjxsk2jsK89lAXiaKnJUM8hMOAt8HahDWec91FwiY9fRYb8p8gs
gOkoUPUc0HD8AHo5HRHXaxXzvErCq29IA/1/+BPAE8VXBzuDCYL2Fhne1vsv
p7hOSZ3Dzdnw+sLleWFyrST1VYTSGEX7878y8lHZlJvaRmaERWlvl4RaGfMj
vRD/VBfwUv4AnE5dTZeOwRiyd8Bi5QgzOnTeChZThJICWKKlLsWwTw9995SP
pR0JeMeN2gUSgpgYrrbXKpAxAopMUbzdIkMThpE7hPuReCQufS4imP3Omc9i
D26RBO8F9CqfMHJK0EqR5Bq285+HIP2FF/PNKlanwMGTtD/+wtgwc1RXDAXd
tl8Wy0bujqyKdhm01C3dSn5cIWEftW+opuYYOMxiB6+n9ss+mdkg84wBARjA
/w1rxuxPuDbLw3mus211WUxqGORpCXKSfk4oKD0eMrtjnLq+S/onZIaExTMY
UI0aAKPvEjgTNGp2uJq1fGOn4mPGXG4Gm4UN7g4RkJH/HEqx/BYQLcTNwDmq
mm0TxPZm0Fq8AAwhpFihwhQyhaZ5qwflZyVfNq8GGBXmoiTw7g9J9k3g2DJ0
Bjhffbx4fCSYLd3G0TRcIeg5Zv3edQSqouISSM6uXHwIOUa6WqhSiyvMWGj/
MINoDnSGWjJM+XtmC498pYbbfs9d6BXQ1GxsR/K9FO3WWb/+PbLfhA+6Dma5
ggCBnKzrFxbTR2X7h+7e5DM7vpB76/njW01/RpTJUdCaUEvE8ZdKBA5OGOfJ
6XXtMiVCiNDmQbaJD3+BzOGSfOSRnagI4XEbaJI6YnjIs8DuV3KGJgXdmQp6
TESKtWWFQpyT0SdXp5q+M4XcB4Mturf/8ywHcD8o8wHCfVF57I6cOs8ShxF6
CprYRNF98mrtmqSsTX+fiNsU5lMO4uRI1fmsK76iD++r+e63yGHQxiGDnd+D
QGxANA6jvHEcAK/bRiTAd+3roRpJgFxNiNIHosCHCdIqE9cW49gD8/f/0Ztg
4OOhQpwk0YttXg8sYC0cnD/tRbR6LtFg8eqOKFZaUO+dTuzKYYctS8tykzGS
F5Kit2iRFrPXdB3O6shavuPs7HJIexLIUkEOwG310kjTymv0aivuVNHI5v+j
zjRSl0vb44as+H5KYHRYsOQGEScXzTg8q/Lz9m+R3O7Y7pOKQGY650KXK+lO
RnXB9xL5GoRCxh0izSd+bahWsfmYcz9UShsxvuAiCw5AalD+MpJ4yRafKvqW
Qqty+2OLeBqQk65AngSdX9taui0a4qmRY05y4LFuwECaDW7BUEddSpFsJs81
qxkrdqnyVRVJUR1AfMTbbGYHbrLiNtsk9n+ixo71Lze4iB70/TLE81s0zZos
P4I01dlEfBxLtN913+F4/lWUzGt0cwgJYktJ5XP2zbwKH11ItNBTcN2iY4j3
MmqJsoud/5V74Mm5+TGZEQJceH//Mq2DZk9jgLhGvnPPacgywa9vVirLckif
/hs0w0N+7RW5IKgVXakB7nkqRMQurMB6TRKsoLx2+XxHvFdDKqiewTJ4fqyx
CMSenExlFK0Oo6sB1oH76eM8jCXoY0bk6l3golDFOgcBWngxptG5KzSGgkNo
Kk8Koy0cKlOz5mV/ue9xaSBEVKGKmA+oQPL8+OsN8IFEWmqMeLmoGtVpRlTf
E2U8sH+bbC8I2xM8lqeYFWhBcx6o9XrDQ8D8KqPflHwKIkdvMAQzsA96qcFt
EWJTo3SIdC/qjIQIK3HHCtPc0zz9vBtjEO5MIqjTQORjbzKgr8rW/6NRtoUW
iCvsJUvTeOoyolpxbnLiptrUH+HVQd8d1JJaqvjBidV4Jsc7Rp/WFqP7StVx
AlFBtD02KgslEuMLMWYrbVkpu/TlJsDHGZMma6l59f4NcCNTJywQqkO/n4pz
dgXEW3+HW4ndTIaKbepahLmBvSgf1pPWraSDHkPySwr9O4WYoZQwYgQIOMO2
LS3ZEop8CVuHGH6maS4w6FThUFK9+8dp+n3S+f/Aj0E5ZRNuaPUvcLAHkoAS
IMrnGEVEJACdkNjlWmr2xLAbjn8t0O1SA7UgRDhiDdcTRrEtd9V7n2mvFRwq
IisyskJsJq4sf6JiwCNgGBZ+J8xNwCb8d4JJUZi0ofhVtILs/RiEFOPCtYBd
L+OmPj2qfvRHb1p6dCmCwNvPNX44EuXyysOkHOBZeGHqS5SbU2ApRgn4yZ22
GSoQMHyaCvuqhDdI8v8N4upDxtTXxgqUqHT8A1imB4/93hIOT/iU1GyyMZ1y
h1S1z/cawUuNJOYGdjoUhqujkbmtm5Dk2WZbXoeR0P2xviSy/SyVC/4zZ1L5
ENOFSqW98S35BCj+u8WsmP0Jt+7/iGbZSDohhzjpsVgCvKBCnh2HM7TPMKf4
JiKP5s9xbPyRDlXDW0Prok/q1qfXbMUc4XX8SkwR7uv7tBfFwJ/B2c130O/+
2RWocdgT8xRBPtDB0p2YvLZpzcX9XzbyYJ9jBvusuJEFRfJFFbxTEVLFngz8
wk1I32iot+UuPB7AeYxObufUaPFgi8drpyzzZ2qHqluEk1W6OEDJkavvMZ32
1GZDyZZFGWBel/QjwNDoE2RGUe1RGlMr1wjyW2FhXMLtuExJvKhxXdtCYMOm
revu+TDeV6JC4YFJOdh4Qbaly2eolWklV62bQESZtJpMxXo8XBiS8XSlQerR
yTiGN/9zV2FCGQxQp+9HL+s6d4QAUXQPfEdoRA67FVG4mcGP8RQKpEyiP5Jj
A9LixS2P5S2eSWMUr2VuW0AVirBy59QHKPiTAGDM/ZmXcohjOOa4qFoPMI54
BcxPgG6oKuyr+9ElFPVi6g5lXvGbQZY2ELPj8t2RcCbJoyacrJKEPj0aPCa6
pUW7qdP/qfaoyWafF63rT87dgtFzKKiXbJm3Ev6P/lObRgKkjj4YDJkd4pVk
fHH5oFzhAR/WETtNLbWIU8GNpa7UXUroipEVZugDZs/YdPcm30Uy9PZrf5UT
6tCBQPqEOJtRCSA84s3areI1bluO7+K9vBmIiTqjYsO7p1ER2DKY8GRlgPoV
FfaSOCqMwbXMY9Bza+ogV4Y6onbXkr48WJZU2+n66aDvsopjdzCJJHreezbK
yllrJrkSO10ruImWBbZwNaxASEN+rUvbktZYxfGEB/kxkx9prJ9cLSzqI82y
k4JDoDn2iQ+0njtyON1g3UYM/5JmWaI1fRIfpE6YdEvyMbdZ4EyD1m92mf04
o4etCBiIZilVP7Z23Zw00K0N9+7qSeR+chLgmhNIz9N5n/4vEJbDgtMKoiZB
4+3hrL1NdDLn1lWbaiEgCM0DzBZ5zYlKVuVbbioLejsme/8zR/+mAFacmjz2
zFMDwDtxqGyLv9jLgwk6Ev12fFnAjTA02VgOa5HyYG7QdzesOxW2QyY2Ye5H
tUHC3E/5ctG2Ab4M8SOnZJBQLE/JCozHG6ion0eLoje1vmS3xbmqt4cnEOPk
sYcsf+tCMweoPDOSpkhUR7hLMtdfCK45ZMJ+oDH7Ogq4Y44bbHAKNMeIR1o3
ptub9o+D9KRQD4c81twMSZsf0LV/gqRNRma2h8jgKKVMEQhOZozrUESCUoAB
B4DWuWkIs5tW14Kf18hPtCfh1ZUzxBdfbFT2VPzI9WFvsWVG1paIa3gZXm5Q
FjqoyfztlzTKhi9FS/GJaZxEXbE2Ie0TB5MdZqnBAWNtgVBekQ5nFr4Tm1Du
GS4s3aPgibp9BQDtu87ENDFxAtVeaiOLt8cBwTMMHp0hbhjd7Vof8LrUq/B/
MEjno0MIBPW7vHX36/e44gVPJoZoOEDej/LZfok12DKI3sNcdUpZZpZwLDWy
Ib5Lb/fhquf/TgPUO8KDbuHiPGRxu/xUgSxLn84VOoonOTr1XAM3/xUl1/la
KkOPkPeK28Na60LLGmwlMK1NdkUG5D3IOw9J49tfSt9u/KP4KhnGTQJxwOba
9cizpYgX2iBkbZFamioFM9bp4vmmm3wvbdV0+w5N1yAmQZOOC5XlzgbJXkeU
k0CNYHu4Yni/z6Og1n7rnhH9yFpoLqRU1/cdpyvXpLFKe3U5HysLD/TsH+ux
P/BPjC3ZVixjumAEGhwiGrIxrYqSkMrKugT8BPS7iuOkgBqXIK2x8NHdQe5f
TPFOXzlRktGGLESM5d3zgTGwbXfHmtyeWGjvpMayiMQppZEUIOtdEVxFJhwE
lKP+i7ed4YmwUrVVL673LVVTjoQgyuVgwUwzJVC2nuhsAUQBA35yBfWBBudk
tft6lWwtTiks1grdCSMmlJnVpdUC7rIQRGmdnCc2XUzMjLq9yYq7kdx2u6RP
3VreXVOdF33CltBIAaWyfB7T5U9E6NuFXRzk4z4tPWccMmBotQrncJnY30rf
L/SGGRMFk0uquewPGORz2c4Glkx0aOAjbvGTxQdPCpgMUJEI6HI7UXL2f3XT
nd0t2m0Rq0xChPRYM5xLWs6P7B4musUyxW56lt6iQb9RtRDWmO+V0LDE0xi7
p5mUMwZrPZzTNZgzO7MIsxEt064UpVnTVQfkdJ+szKY4aZufw4YyeIoKUbKD
XD+Yl3X0akpnSx91Bb+xcU0ZYI/cpXdTNdwjN/051aQHlCs6yTsEaMEfLC68
Ebl4PSniZKNMXYpIYNJCtB6GqhkADPWCN04YpAWlDNslVv5ALsu+qWlzVl/J
PJzfyBb2dKIEnv1FWRQeTdlhhcWnCmk+YmMDu/uS0LsBicHAsOMoykwvErf+
cWvlwj1OqJLJo8hSCMnAeo7KrWgRAPko6a9wC3xB3htQtJMSrgZlI85v1uqf
9FiQzYXu+p8HBouHy/CAnsMtNAo+IcgxR4X68mL5D0lOG+v9hMtOkGjKQfGm
lGeZnPSI4/SNwQw47ptlV9R0AP+x3B+c8MIu0e+yGqhGbtTJ9Ql0W4DzNoek
m6vZa+7Q4jeny153/UO7++sgLICsPUxkLEY86dxf4gP85pOXaCNCcdDr2kxS
kDdHbZVFldlqcSondd9ZCru++uLvhL/JTEP5kzZcsY0dsJAMAgtepX3h0xn+
7Un7ocJNBAtFTBQg6mHU2RXSByGYMu/zUe7cv6AENuQF+fiL2grwr9XHW7Xj
9AAZ9i5WYAX317WK6WHkeGJSSq2rSR0qmQVuD3E+J2NcrzBL+Dvu7BsOJ2Sm
GLf1/gJhqROBTT1WkibY2oqxfz/3jgchPblGKLkZv7L645lQRUx1iYrv1LdK
uSip1eaGGcruhWddANY87Og2pjbEQqDx9DQndgETw9hXEbWvZJO13CqCZXHI
MQ5Y6sQWLKV4RgxWcUhiOe2Cd47cTE4H43FGHiu0F8hT4wvchUvTeeMm9O4W
XRMINa9KJlHPUSzZ4b5lpbwqZzLRuZkWT1jeFuEm1SJr4ZIgQhbELOe9edwY
nvMfMUtUs7KEZ9m+BJDP1tzEXnKwSPVCEiwsB5HY3bntbeI78SWcYc5B9aHL
M4YQXSQH7fv0nhyZh+ebOFJnK56HUY+QYdEmn+OVW9HOhw5+hOC9ofG8uEHu
RsSn0JRHnKSjWFQlUo/ZT6XlfiGpwmEvJrxLqM1Bt/c5ipuCzKASvigZl4AJ
4w14DpDRNVVw/rLQwbiq/iWkCB4CnbArx1IFTtjzI/LWw6hKmrLuOEZ9bjWX
VZxT5sXutXeZKT36GvqOTuCQDahg/YOQh6wQXFGppUUfzxvDofbSKBFrMrAl
TJWIMNZeyzxWgA4ubVxy+TLvwyBotDNZRxP993+zzmuuJFpXS9Q66+gzeYsc
8l1Vmpfp3oApvQT17ZoJ7exnusm60/Scw+23smYNVt1vaDljhXSy1G0Dtc0H
omuHRQ4yDFzOBSHP430mg538B1tVMcZ8WsQ89KGqkXcTDi/dpUilIvlsqet7
WbiOGSOXXzXEunQziUYU7cfzN/NAUUlMvEvfDm9u2nxHLzJDbGeSdeLyY3yY
Y1v59PR0CbQy4RE2ZLu7owK42erZXvTVmjIrD0fh8EZ1L9eo3A/53r7beC6+
P/5avc6o6GFRN/CcV0yUvKVwxvUVi8w2jvdM6QTU7BSpqBgRYCBIj1pmEqgC
/O/nY5zHLswdjzh2d9Md0p3bWwODnyTgHNPT0QXgDTAazPtfKM5H6V62Ladb
+uJh4AD+mIbXQc9wDz3rBsOIOS3G7paNfcBt68qoxIvxwjzMSIpokis0qUs5
ZJyltA0tdUfFQVgtypD+XO07VXPxE6n5vMl0/8huGLZBAoOoUhm4Yd+5hIQq
B53jnwcGDWLkcvXPR6gbJwkuB310xeLxYLmsYI3LdkHmzqeObvSdr/QT1p8k
y8oAYQpXaoe+jVU4ty7QaurDtTjcUrDc8S2s5HSTV/l+Fd6V17sS/8vLVT1P
H51AntU/mIUsSt5eAcvS8c+y3fs6Rc1yRfIWeqVoyQ+vdn0aBH5zWelhjqk+
srVp9HN5fU3QxAkGZrRilz/0p/VVUOWaFqeSVBIZqb5DxURhbsn4tj3CA2/O
T1Bpknn6Jw3JbDjMJ9969WjWnsYBcL0AZQhfwYzRQ1Z66DKWyYExwssD8e8w
gfQv6iF3kQZf62HJ/9iO4OBxm5FI2fMv6iBUYBp3ftKgUosGLazlXWvFD0Qq
1Up+DhU/9+wssZKIyNfo1m6NhTl79vrtVIy49BFO/RWs01jCy+4ZuTgDnB/O
uO39bihnsfm94pmxNk5lg4fExTUITEn48YPhJszHUtcGNZBgaoypEqGTt5oI
bwM8Zj76In9e+OmV6IQ616tXD82mxdhh235nim3nbYyYrKcmW/Fspf06jS7U
254/P5EpsYTWn8vkUBdyjXs3sm+c26ekONCiPbMDtmSvAtapr47TaW+OKXA0
Hce6VsPc64Hgyk4T33gwtWdZjhsTi5FsV5agizDvGml1z4If7a28ZGmAgS4b
tZcnVF2B72ChISPllG/O3lXwab2snpyYKMJJVxlu8AKxEUlbmWgC2GEbgdi2
AkkO2iw4MKQtYhnR3SMG3UjPJO5UJwsfKFmHQ5NFciDaAh9RwDcOYEEN5U8m
e1/t4x/3VWFz28n6v/8iTOTojgzvgFJqepxYOBAvni9PsDfVCa+nlzcWLfOv
0yfoPUWnheeJQv14vxojw1hqVCMsekGkgMKNRmLkmbHUOG4VPEVKsfLp/GZP
1DGL+GPjAEBa99K/wwBxfPXY3V4dfSU7D4zUB61f7KivyJsCISyMOrFccqoU
nZksT9+Bm3CjrAq/SaugkkuF9rOniVKJwlu/7M061/nidLXJeBw8sOXTuye/
stezkNoEEza4Z7Lu5yrJRBz4Y8FRiNo+xVZvsFSz5rfLN6wd+QODr8vJFOHm
mTMfVL3kJxO7izr0CRa7iAzERo9zoiN/rYrixvb6dMh2dyJ3krMe/8ZgSZhn
sX1nrB14NhRVnC8PCFqzkbtT4eGy2LE2Z9C6RzT2P/EMq2JUnyl8plLcccTi
lS0nuXAnzj3P7HgG8z78qRSOxJTmCGu2FDtDf5yBF1jfLZBwebTuPDPGFJkX
erMT/6RNRIMtL3yc9ch5i85yCfQmQGyErbiafZ7BBcqgq3y4xGqYzMfY1D7b
QkuLf5siHfcOoluoEqKBSUWWVRwZVDXCvQ9jqZ7Ag1AWjPQR1MzOQJuJ7Yl6
HtjfJA8SOxn+ft3ADCdSxa2p90q9C0Q/oEyqtjUZ5RKcXnoQmpdIIOUeg3al
u/QI+JfuLfsJydVvhUXA/dmMGVh5QBr1wh/kahJqsS8bsf4N76Jera3OvySL
tDNqpoDqthS0T/61+f4XxbVTVTw9Rq6PMTKXSZLmST3kcySP8nlFYtnSQpdq
M8ez7+juM3Cr8v9JYy4CHMu+vuWVqKit3NRcmUGxLnggIdnCk6U5iJ9Y1ezb
5he7ESLaiksNxEKK5EhbRx7JxtLrOrOuVcme9IVXa/LpaobRPXAPR0SfRahr
O2iVLty/owenkcFv3xxSzcyNNcEn3REsQ0kbPgDFRUwJaqKsqj8j7adUYJjA
6HOJVK/ZZUAdS/+e0Co+wDM7gyVZHDo007A+u5EL5f/Ha5H4E8bEcMpS4qCt
IEbI/FZras6uiJkCFVpyMuKH6fVuTUCzuHaJ0md3JKEc0mEJGRQzkg5mqk2j
WupNkQh9ir/p43uQTkHJZ5Npkf3tPkXQZLT2HvFHwyYBhp34preG78TXWyh1
DTQ6p71jx3uUqYfMwqItSBkIWi2m3MJZ+eryRc37yugjB81CIrgiOA7Ce6Xt
tEZmdRvhdW1zkWvuCQILYIyB5LM1+8EvxwreB/8jTWqGHZtsZsYlznwnDUXl
WjGcnO5C7kJT8aMDqc6zJZ3/W46jHgHInQj5PLZNICn1NHhlx4bLaP0M5XcE
28HDFyWz7FW6qJwN6GfdKECTh0zG43UhfT8+z6yBpf3rshXxX7uKR0riGdeQ
WnBvj1CK5RpUaghzqn4X4av7N7qIH5LfLYn0k4qd3CmiJ1GAXDcA8grx6Bo1
/GSxC8CAqmAlOQxnT+FDOhqgK8C4BnQacIbIVrEg1iKWzdY2wQut5Kp6IlgC
m5vNgJchrkeD4wjyKx6FoGlNjzhLC6D8w3NWakTVXbFEGP8WFk0KpJuBS55C
F0C2uilsoKkCv1FLOpWVuHOI4adVIV2euxUZTt5gBqbAaFBkJ81OmbywFf20
66LNGmlBbTYtRlocvYz+TagvbvzdneFZo5tjaykqGm3bE570sa/Tk+Z5NUon
N+D2FASxv3QFkmcQ3QHfxiDsJ8idq6zoE8wPjA0r6R7UOWiHfsSuLfIwRkB1
hilLtK0CzRCeOGKa0RpObEA9laueEJ0D1RcwVnIC7tk028JW3TVJ1oN6nGOa
4Xj3vxmCBI8LvshXDhnBNcPnMh/RcEGjZ4OT8Zv2XZ9j5qLCN74+U8D6W9Hh
6MdhQsPosuyUSvwCn4lYaeA29nEyHsrWS0kCQHDRj36oDC+nN58vwJAcef3F
SNd0W3J/oVFbJ2NBAKfv7sgzbx8LsR8PQ0L77jd5AHrN8qqyLgD+hib6FjHL
qwjlALtwc2/7aZZqqtuSrIRZPJhW3l7Q/k6lfrH9J4DLcTQJQoCGBW45ieM5
R0l/d/h9T84IQIkQQoKFgfqPqojoRIygapy+rjWgB6JlArl1Q+w2UCMNQfjK
JsFh+h9PvZqp1WfBA26coII/suol5tzHm+Z4+DTXvnB7vQdNQgOtKz3DH7CU
Q/3cH+u9sJ3oZdfqRhtrPX232y8hgiB5khM0VLrMMVj1M1TRp7Bzf36TSpY5
tu2FWmM76J/BA6460pe8q/qLo2TlqLUR75QTZUGNoDe+MuealCOTA5Mg3RwR
jINybLiIdx/kSEAdyDLl5Urgywb3Jll/CF8mPvgoe8D4I2LAo+UD+l7Zb4Bi
eI1JmNHLPaKljlT+m1Hj4NrvaHlF0bywILvaXeS2jdpq0xvfMwHisLc3mqnC
MhWgSflrJOrMSVf4vdrzHURp2QVNTVAsQhdSpdJkr82yPb9KRgErUZFMPGoZ
93Xx0SfCM0f5SqdU+7qEzzZYs3c0JEOiKZZxDYs07yroZsVaQY5SKRQTD9qk
NlGF/1A/XyY9t59tUJ0vH9aQdeAspehDrexLdj3yuHZ6ik+/ZK7QT+Ukgsnt
KglftWdFmsyLZ28w54ocYov972HL/8uV+ACXxFyM3NoxBeXz98TWwj6aCnbN
dcHuiMz99DEkzbWbxAAYQ+PRgZ+7zfio/4fFTo97SyJKzXmjf459TOs/uE0n
DmWv+kN6lWgL54NxvOStkdOeS2LNeyzodkn8SV3HDG0kgEJ7ZtijLpeR8mAd
enGN5rdgcH8qzFoQHpii2vMDhpG85A8zlGNW/dj5y5Lh4I5ZkLF/8VGx8utZ
j6hKOoTG3FPMbkaTOtN7XChLDHq3FG//OmFQdJzEUMDU4wI5WgfTHKBxoVVF
HnEO4C6u+JagMK+Lo58DytfhcZQE1Bln6tomRBjri+M9q8F6/HcvZQFCKHXw
EJnPLYiinu7L0m2eWyvqzPDMHGIZIMjJizBf4u1yYTII5DMdH/L7I3U5Pm9g
IuUX7Ul5Z8vOgyj/rhsWkUmHv9m/2JhC4kh4mKuODI3ctMEVaFO1VlgN2yF2
Cv+XYYT7yja6vEsyLQqdcBER6Ge/F/yDxgfxgXv53WQ3UHOtLSXkbYsRP756
roZad0F1+bAFADfVub18X4wHvZ8UuA/6j/pED1vaP/xmHyHfvDZrS6MIWaML
B5d8xQBQ+VrOIjk4i9rzAXrX2iN0CfIfdw4IvnTfMW202ScOJZoEsdW4SZxv
fAtV09LGfT4RvfNyNnbZdyGq1W3gt6NVjV3naKvoQ53Vxm4hWj23hvg0rybf
POHdPVdpvpIiiVAyepak84fI0CoOgWTGuShrcuG7h04YhvXpC3I/ESnYIcKq
yfHyNZWDCx0ipg8qccenllNzlk7wBkgvSh8ZbUjHIGk8OGoWRkziBgsX4N5H
/I4TFRqwIrQhh3yeiIBY9XpDYtcvvGC8ocp4QmlS/skczMFGh83uhoAQHsxE
B0YjpJNXGb60RRkU8OlHpR017oyVU2mNSLok0rBCIjT2U5O/7WSJ94yy3QiC
/7fhyCbzUu0IbmfdNGRIJ/uTItcincTj6KXJPdrOnafXr75Jd6KnOR/YCpQO
D0/7WW3FagnNylyZFXuWcT4i3k2dklA7hXRwuqUWsd7PLqoH0npxFAOpXKvx
ZhSPzofCX9paZaJlM4d2OjhpqdQCNvU+eTMihQ9XSjd+cEv8a/B5p7SYaP5i
LDEHyzLdwgGrteCiK09VI1mdJWWtG7JGBDq/+zphxZz/M4mWd2Jcb3QtnSpX
PHLjCphvvSyU711Os10wLMJDVrtQJth4J9+zboM6wVDpfBHE51vh1TGKS6rZ
7fbG5T6fqi78w6I2pBmasixDOmnHh5gpYrNnfc4//pMxI25cT8kSCx750wO+
lrV6hhSpJlBmuAUigt/ORHR25Ldbqanc91bROAyL7EK2FAfZZjB7YL5U8VvM
Fx1kO2b1l64oVt42DIz9e/6XS2a711nXBX4WD/glwR7Foq99WpaUEOpdJvHp
zmJGiGVElPtve1TXIi0sg52yLHJ4RiLO7DH9NP2y8qYYhFDN8pHysg7PBwfH
VEClEmfZXnhKkPzZ9mrNZTt8FY0t8k239TZZD01h7cHfVMBU1c/EjlrH/QKT
+sFpkQBHNTEdII57NXZuj1eYlau3DhyM1yjWc8C4Q6a4rrJ0oxWyywC6jjtv
NURWbp6J2PzMUeASUL4CAktB9NW6KXoAL3niWInHthAUws9Bu1qQnm2ML/0T
0DDgUt9Ku5F5I8fQkMEBW9cLLRyogka5KeIZxHr+dVe0uisYp/AREQE2ktSq
O2iuAOt6kE3JkxfAyTDJpSkqAh++Z72qeTAlkxnqoYKn8PwmKtIiSH2A2a7X
XEbIdMqqVXZtw0+oXMTpmzPqr3PUDBicfOIU6TaQrGjMBoYt5/BXioSguf3b
b7sQL2ykXMLkT806Lkq6PqDEAUuspQb6RoipI6SxuqHGnFVHS4V0Ct4vmENS
zaQRRkOvkYxrdrpa1AUAHL4Q6o2Ylp658Yt1FjyyXpQZmuAy0EOm8NNoClKU
/+teTyUwZn6pLadT/UZSZ7UwxvYwDArHAlzfRm5sEstbvocE1lQqeUDG8haA
gKKHaBNvjSUTuLXmByBnjIRMjRMoOCbH0kzge8dvuzrkI1b4TGLjSAZjgreU
S67gS9UijEryBfdnzGCbxbf78LDf3FFdnWESSFnUFiqxW5B35mhWPWdwqf5D
WvcM3Z9WU8ULFInJMUImDhELAN7vmxOp7KcCjVV2NC9koLtK4wRMywWpuakO
IlOSrAd62+UiNTuHPv4IxdRlrlMx9rpa7LUUlWgf/ABKf/m8evZ39swQbh2F
7mReoPf3KzRTnu+qIY7aDIake4wsfz/L3tLSOWMXlQlFkldVieYGRC/zdspc
+gl3se0CSA9T3uEbZQwASaZdwFIh157KHfBnZ77zGy9us+lkD0a9ZIxxpNZN
855aAKZq73teG+ewpve4m3qKdBE0/GJ2bRHKsu4+r9JeEiPDAsyTwtqg83Xl
chw3ddri3K8G1TJCb5kqOLkIWbPzarGsnRYg1sL84J32wunOpV4/3CUO94S/
ZJowfnBlIJw6lEXjxXhTOc2yiDjfs4OCpskW8v+0LlTboxp8b2//cDpTOzYC
Ry80t0gNM4Gfr4ZgjbiTrwBbaCSS9l5EkWXt2Jy4OZYMHSCvniB/gIpVKQ5E
17OjYp/UUvIU6K5jUpFzqNeP+wTqdRsGI3L4hirnijR5iH59b7+arHuweuDn
1Usy7Fobmly0IM2Yfe/FepQst3G9Sm9/s6j3Za7MY5DvUxlfy2gSFVTyDlFF
KUjvLr2JywR0xRnQEcExAYh8hQnieOxXXUVX8To5g/q4Fef1FrHsuEbvtNc9
cNp6VD3N0QMbj1TTu48Ap/hfyIHNsEUjK4Z6E3tKqr2DAZ0LtlVdFIzGsIlG
8rXgGuIsYC9BLVHpixX0CFpMbhzqKyu2NAV/U/7kEMyg/E6WsLoY/qQQfAQ6
rrOg00KhiwLaR4mIvx6UMvG3z8ml6lq6uwsXjzXmw0y1kQWCjbsek1jOq6b0
2oE/lwclii8xZDPpGR0Ixzj0mGQTRkABOgTeIlDh5xVQQs+H+SJ1YCiO15Dj
HRCMQ0MVjOa4ZpqSm+EK2/eraQxWLEgekGf5rjmTZAfyRCfNYQCWoRXe96kw
fbpRP3LKAClWRbiFhYS2N0H5SBrWAqDtR1nFKkXmtBnxV2PPrGHvpBpRjO6H
LVhCRnmNq7wC+pgg52WbYkwA16Quhm5jPht7bJTHfKbanzPCAp29WBIpE0mb
WwadymlJc8RJCed1P+bUXXPp9VZbB8JrFle3Ut6I7JHXb9aokv9cVf4N4Amq
+CkcuHjzj6Cc635y6vChg3miAiTI8PVooK/3VUT9fJEtQDCrJtnevofAT2R+
0dHshNiovfznijv3+0B8oIVcFR4A1882VzHJEUblVij+MK+ybyeNYBBFU4WQ
xORShHRb0G48wmDLNlq+ktv6ZncYz8pxiixO/qvxXKHXn7yp1baGHmZ361oy
UoYBY5z8JAw5l0pTLMlYc8DFmdS46KmNWM6CObXEDj0v3vY7hhTkdYHxbUQF
1eUiGOvyCh7+MgxkM0NT40Q/VvxeZKcWm/p6wrw2/yuZwlY6jb6zl0B/Gudw
JTp+rNTkSTCsa0Heoiov1O70KD4AZ221eG5Utou/M0KfPlaQ4VcGRUvkj/Xd
pgseJ6mkvSeDHXUjSFvt3vZ0qsLGfmoyS2VNXKehNOWcheXYohPOVQd/xSiF
ALEHgIKnkq5SmwvMPOrFMi9nflEXQl+88muhxmEd0DRH/I1O3JiZk6fTwWJg
+kwxCpnEV335Y/uzIxBMeWHDyQutZBJXiFRBJNrT72Oh9Qr3oPnRVlbVuJfn
ZvdUpTmy67mzUqX5IgFKwq5WYEqftPR1JlnJj4RxeoAEWNevRmLOucEBTQmh
2OinKZMpM5+ZRpLo03J3y2Q0BSeH/wEDyYrwVKtlDOs3+ARIl3Bqm3l/RBFn
Q64iwRxFbdwovGDlEBy2LXEwRBFHEgwVcRRnppXPwxUWsR2ncuoLHQISZE2a
MRCHlS2uF+Ht97m6G3pKzZ56x6a7qfLzNbRwj6SifAgQn2t9D/KMHHQ1NY0p
609HtBj5xjRz4KDnMWVYRoMun42d7oDbdOtx1V1HO9GvtPzH+LqMKzw8aIZw
xRuXPlC60ujTj/EQzKfSOtK43Huq9QWNnq3g1iV+Icr7JjuqVY6XcJ4K4OcF
lvZu9Lk8mqf9KLwDAOwbl0u6BlLrVCG1xg5Eh21MKz2agI/PefQltNO1WdYp
wdsUTQh5PzpYUlnX/Ud58TTUMQRvhpLnJJEsSfaHuvcSI0mRIN/v5us9wHVJ
tWkKNCd2eIlgMJlY8Wyzg3i1SG8+xkgAW1z3Uz7ztFvMq20CcVMx/gb4Hm/T
F3qU/Aa7yCxG4OCFZ1VsC8F8Jroyp00tg7YZo1sANf8zc+JM1ZonxN/29gyf
NqowkGHLOKbndU/wSPC50gKJLq2qBiTOAGPRqhOLXbkLd78IaKNe/YAZT9+A
UKLUjjSOL8vM+h1ES184SEI2CY70Ebh/T+4Wuuz6VoP6tjcy7eXtErU+H9bJ
+5sj4UJdBwESx9ym6aarywjiDopuvm56GpoOxh/7UmBL+APfue0H4ls832lu
Wv34R74fNy56g6msjfys4VwLUqd5UUCoDUvKqLLfQ1Slp2NgeN0f/HCo2QFi
olAxBI9NtpwonJqgfGH2ZX1ZqMcG6Kh9Rb2E31WZEuBHBvWOFjSbkPVG7bEa
bLkO163ekVpDMRoP6wvHIA2VqJLSmtK7s72hj+bvGTIJh0uFgfaGJFORrqTM
OgDe3hs6ADpOkeONhLVydLI50NeS4oV191FjIY9cdLBHVJFFI4apdDxQbHTQ
qDNjOEsULvp2OEqw4uxNk/sVKzYlgEirKZvxumeiRlcOZ7ChlzMaA6jp1pL7
BtSffwRmub6FS7y6/FlqW+j73LD1eD9a/zgmv1Yls28JP6DX733/7GfInhHJ
4wmrq8ZWxSjt39M7jrUTaj+XQSDHRNFTq4mF/ZRiA2ZX3axwQeGregVIP2qp
jh6zqvIAOHr5tS3CwfMmWNZynjvUn5qj49g833WjS5kayqvLzPtK3j0fpI+s
y7fXbAwVw1PrzkI4W6I8A+jf+Jlrg0ktd6aDn6xA6D5A5WN+VILmCzP7jPsB
jaypdEHXBLJ6d/cBi/pX74/V9nOQOlXNanbzD0sJsjrcFc1zeIDIDJeQgAqD
wZzeLep5uqnweBjQr6fycAnkrCPy89Go6vehqTF8X0PooQavtavFRpKdtrbY
DRbNXiwTeJi4LQa67XZA0BoY1MijhNjjX8SUpm910Y+woN/U/OjfxWZrJeOZ
2MYh46nsMgwd3Ky4CGhpp6TIGZLvMYYdiGiC7Y/72VO9kJHRKZqLnvrsfgpH
5cXdPP+HzZ5EMcvjN1KUmeTZ3cilrlwvCNeZ6H69bmPSTlDVqlIguaRfzfIb
zJY5mN5IAYDHV1kXE4/OCM2aqd9XlcSBW3QCY0KduKIsPfpXBMzX1R8dgqZq
MrQ+n2CDpo+/XHBHcjiUuw07/T/mfLYjLAhCR0ELpXsfgJxTz0AZCS4bMBZI
OddX+vylIqW4rwZi9ti/0FgZ8uasB2g6NR6ySqLoh0DNHszyrVRclMCDkKqt
2GJw8FdXaPAVZPTvXwNjof2Rpv3uyQGD+HBixGgfsV9j1szlQS34L3o43m2J
q9GYPR+uYeJnAwLQe6rbinBVgz9RVVD2hLKeI97QjL7vHwt3ZzNf9fx4zwUs
SA/QJEKYKqMF/uFJhJ9y/233pNuzlcrcckUYeb3X8E5SzR3OWkXBZN6lBqfm
CKzOSZ4hQpWh8YZAyDKaXZz3+egGf25/smsuhcYjiLaiMN2vcxMMU5g7I9M2
9hdSA4vbHc1Rwj9szupxtNcYiigIZsNL9lFTSvpidarpGzDbQbYyW2dj/xLg
82F7aQurbcG5At/eCq9rEUJBtS/ltsVkL13jKAIoMCtfUx/daGlKwJ8jyJM1
JkhmTC1w6pKqwortgsshp6gS3SiWm02nBel9icGlj5q4eosA+RNVFiaMhwdB
R/xCVHoHJFMkHrpas0Qh9Cvj4vbRnGQcnaA6wo14iN5o4Zs05OK6HrbVDN9s
eugLVh6Zl8AhOkfGEGFLX2mKDy2Or632O+DlPn34kwQuNh9YyH6Dsx10369l
/0agCpgQaiek+5j2zdM3eHhRsq5Q9jLk8lf78rhDCJM4uoQW1qMIwwJcKZMO
vIgPWBV948zPIemcVrC64Qp3qucS8wbVW9bHkyRGP/pgBZybi633F7z2TnFC
PpyVJZHBViW5f3BqTDLth6YP4eUEBHG9F6APPY9FUDWjOrH0HOJXNNpCTunh
b5XiSl/bkABvknFD644Zqi3dw/XDXy6aPipOsys4LJ02k+oFAEgdoKV37LS/
R9MrsRJcFSptPBU6KgyftE7J7KHKaHNuk2V5keQzkj21vkxixfNb6gijW+aF
rr7scdCxNlCkoEbH9fMOcmBL3iPO8oARecKK6Gn3Z17WD1y5BCjQZqfDTgpV
Rh1mjV45toOeX3yeTdwDy90Az/N/18gg3WlcMuXqHe2cAiWloaQnWAo8Ojsz
7YsQfPsc8A/WJ97H9HJujCKiO6jGVtkChB4ux1USLJDFcHefxA5Nm0ngeqb4
oFVQGD5/ZU6Ak6olif2IcOqfuJES02DTcRt37beTbO4xgBSfDn8nugdZZw3P
SnoeOnyaoqEVPWgUTcfFI5nGj9G2NGZYUkLWH9WytKkA6cmLsuqsneR++Y9A
nVV7sOhIJjuM/Agdp0KJPEKWF8UVf/owJhoWyqKLYA6IApPZSQQv0bIhgwdm
Wrq69rcrzVj8RKom9kylFN5jcSNvJ0LXNffINxJEguvTwpPy1shweYY3QJcL
M7M/yQr5BteUi7CDSllA7hPw8pe9uKSQDUogZBgdW5m9c7X/rOAVADBudT9W
ze54O3wamnMnMgZNPJNWp6Or5BW/eYszyLW6iJ65QhT2XPAxuaOGtpWE/T9j
q8OXd7ZNSKh1sj40Af5PQSGy1EKXpXnbE5iBGX+cW0cbXBkAe/YXEJoxuJmA
xqfVivyu76Gto9K89NloKLE7RHhCopaJ6DcS+bh6j2BztQxsXyYC2qXifAdb
BbfZTy8Bco2PUDuYhfg2PY2omWWg9bzS1ar44b2fwotq/nDGveM1r1vemDfs
RmdLErAcqS4OcIhESJ7y8Yrk+vR8r1FXRVhNRJGWNwas/56hERb4pzFFFRws
DvkgOAdcEFg7s1Zv0Tp8FlrhHdNRHZl7NuWq+dSDAd2BJQ7/dgYadzte5SmN
o0LjBYmJjoSEkK5BtvL010qFRcGoGAqvzFZrwWDHVKgSinX4GyJ3KbZReZ5g
my3ieDqKJsJXqa5ZmlctN9llHq7NJvyQfK3gbPOnDCMM9c4utKgdI0G75Qn8
VOW2bAf7XlzmfLOzyj63QVyPEz3/INx9YZqmgqd/nhNbfoKubtK9DCN1dXMi
0UG+pRLMQXUFeJWjI7nfvmAjvt5jvyhcXqbpQBSv2UvnE+bkOTDizqePj3ok
MK47Ajz52VL0kXANq9usMma+jsBOvAOQU1HrFdWP5erl/kuzg9bhHVhPf3VQ
zD5NSnPffmlacFAd6MplqMQyOmjSzwhazQmeO5qzXnOitzXss3AKejHCSVqQ
gUtIFczXpxSafsq8VccZeD8QZgelc3ApWOn8zFPOGtf+9LFNjyRv8oGrcC1y
BQ9GIM6LB/UHnCVpqUWjMU6NUuAlL515tameiUXXOQnkFK/haIqJ2zrOHDnq
5LV6NKygsIB8slqdY5ZWzwtbLl7Nh6x1i0ZPz1c5D0g2xMzy0DYF0yN6WQDq
cVXvlwoYOOq7PTKwaFbUTJBO9CNMr29ddEstpyzKBPf4YfUmcb/B7zQv1GWG
C0RKmzhgqxTPH5LK39dNhczq+5AstuCzpWPg+IUGU41fiiCIafXV1eI2fV45
Eg7X//oGdvYWuD00YYzpxFByjv1Gry40fV3nJRff9xFht+rlqBEkYzwA8bwa
nP95OuxrI5g54wgb+vOXwEIUN3bTapdeqi7kst8iorn1gIw0KLQG+HYb+7Nt
jXQD5pfPzazw1+3myb8btSgPbi92fcX7juqYqXqdPd8Yp9s2G1bTlj/y9svo
yZ5hp3AZq+KqbyA/v+ibEyBWhwxL1hQ1EPRfByARSQRCVTExK2iucWSdZFgh
TKmSFcoUDaJP07pPZNByhdFJoWz4C4DEPTszcaeOXx5pNDSSMHAtHSat2Kiy
i0Z8SfgiiUAn09HPoFnD8GVryJn3M1AhSHZIAyxaK0OQJXE07LrfWLW30mGG
zhro9xdxlisVO4Rn4a0DMgMiDevGGKk+rnuUOwK307zCixVMORXX4AVYMVxZ
WhwZwqmcCv0bXWXj7PHhZDbHNcI5Xa3CeNCwUS3icql0/rChoReJseRGyrMO
Vs8cgKZvwVko5n8ElMOdHKTE4BjbuCJzBq7owSJ5ZICDJVJPksVtrW50F7Ra
jrdpEx/9MhJMCcc5O8W6tH3QbBPePuj36qGcjYvhf+aAB1kGfvkOcf+dr4Jh
TY+rGAlDuyDLQvP3+NGUdqc0r8eLgcMhFtptxX4+PTgI6Drs3lSWlLBqqUhg
m6VsKOZtfUonNGEC3QVBTekkAV8fVRcOI47eQ+HI2yGaeuYpEB7yMvuqOjAa
2lYf9iJoyEtEcfKFc65adQuxZRyGivYPiSZtvLO/vsYnC/K1dkRx3c9bEu4N
5kkb6qyJmU7TfLc/Qza8iZQDQec3aALw9lyS8MgFsAG5zjyhYgbylWQBP3eb
zne84ak/wZR7kq23AFEPcxITKn5akL99zq2iNYNVfwfovQi1WcWxbZmfw6Fq
6Jr9+Bw7tlge2CSCrvaDsQupZtPgBsBnpL8FXYU1V8ZMHPrtLinmnhnfq1hc
DToQ26QlujRqS7V6xp0rcETHApuAfVJaJK7UBa4sfUzmnJ31/cNRKciXhjzA
RiBvW2ueTsi576Xi4zJ0rriE9sQwrVmzZwzRf3TiBiPdIE00Ig/fhJxIeYfO
u7C8zHeT2GGlFAr5Iu0b0IkiiTvGc0oq7K8srfYkeUJsys4s93np4XdlEnrO
h+w1XyoAwssnXYs7jre1Ha5aLUe+EfDCqZd2oWcU0OU8B560GSV76lQY57B9
8odZfTHQWDDMqa1X9SX9mxCF+nhVZ9sfxBSFinj5yhV+vZbJfTC9Q6u/zIim
NUMHv8ggD8IUPBphyXB2WusJ3NtSvcidZMg8Ar9IXaN0J8bV6Ry+robEhiV3
qTBhJmVGd6typfIziWYNAViGXKpv34v24bMwvnAGaeT9ICujwK221l8JiFYq
JrSjPafv15FvhWpc+CtEoPi7QX8zqFDTURJC70bCPZ2+mlE8Ey0dcIAGBV7l
Sz/6hY3cb3qQOKxltdJlzEXLg90LtljscI80SP9Cvt0m3yqVl4xe6XVcMDxr
EH+1S9a9dLVTPaQvR7RtFm6PlpqEqBAxQOp6/XvaqVje7poy1N5NqldbqwV0
rRnPvORPadrqjDa5zpW2fd5wi/QH7pyg4gq7EXylbRW8NjRmRlbcMB2YDEkK
ye/urZb334VXx5wZVn0HAnmPZDGbpmkwfppJELI+bGt11RzzhehG1Aov+VLs
ptRqyaJifGJj1M8eYNrErWjMJIHoop2AjwLAIp8GDuLWshbovDPzL2XcUTx2
saqO3v7saZTmeuF8PN3XOaZg+yCJgeLYkvPQRDsmDlsj/vUO8or/8G8xCTeW
s7f0ZiyR8zCa94OAc+b5dQOH+aQM0Ixf9qUzeTUOYk+o+9KBKUbKuFfYJFS/
t5yfkGvnj536qfrjSUae/TsDIadl+p5JuGiayucn2apGQbDfNzid7KcdhDHT
HNDqf12aaloBU7TPy0BWcr9NpgK07fzwoJKX/IpsoPD7FoqRFuktc8xvh3+Q
3ugSVBWO6E3SlkSHoRvUSvlP7PnQda9MOLQpaMf1E5JYPsyUXU32t6Ud+I27
LbwGzdGSd8WRJqdz9CEPENGUsYBYWMHn/Mk1TPpNjKAbm7pse5pr6olLIg66
htqC4CHzFhx6y+IuKgzddCOEkyeR+QUYbQTO6LCFocfkN9NWvyjwf3HdbZ7a
0m66wygo16NdeA+l0VK9eo0jXhFPWJMVLZm/dnO4etwKauxkBNrFWI8rGzEY
R+FJJ9FTOx5B2f5mlpBU0F5SUKdNqU0fmotBzzKqn4eRRE512rK0iDZgulRz
OYOfmIIQMtiRM79uH5MCJHulrUOjvuywjS5jYxqhKHpICxk6kEA12BQzFdM7
6M5kVIh3b3JfrsjyWuO7K/Nl2Kj4reyMzE+FrHVb43QDDJrf3CZhcl+BQFMg
6u9PcqhTYqepIPDKodRrm/ePNetlCnEAp4rl0x5mgHW+sUniBwoXWuF3WmLq
7fV1ZGjTD286ocvJ/LviLou8bQoqP0n1gcBmjQYzX9/g0Ca8ZCkw4JRYdzsQ
3gGuL+L8jS1ZdREKU8vKrIAvbHOlE5z0ZMZMqW8yGLRlRyB1X5IoW/EKGJoE
cIyB6UnXaRNfeTYfVuLjHjpTfT3ZUTOx2N6vzukgfhWcPTc5CNGc0x7gg+OA
KP3qQxRdXoYXG4Ao2IIGk//KV1g9uOpEkMSnH8U1lWDyIuZDibpqpLKEPHpg
vXlXVKp9Za1GDRVRVt201TQiXzrUC8WezUAfr6tNsBisZUKnnL78oAKbDSpo
PVfzAMxwO6EnhdNUswTXB/DidRIZrhiWQeo0Wkp5gJVMkQXMgpKLaRwq26T5
7ErycC+Nd+51H0OTmaHGf9Wd5OdZfbctarla0c9O0Rz0xMvAYU3wF9to7UyN
a5EO53NWtDcDuCygDggN6q4E7+OCEOmv+oXw8ZHPSFiadiBIxHmL6nhX6dDn
hfssp5ykt3nlFYxpJShuiBXk0MbDqEQbeFG9lLjrQov5f1GpHTPKtZ91dM9M
lubudEiZ8ZN0gfr4pPJ+5aB8G8/y3F9bkWJ2p3x0IHEt19wr5t1R0h3lqI38
UZT6wvIMCALUomP6z05GpH/kT8+SDuBz72+AeiIZag0auW2j7mqrSTXlgUWk
tQ6IyTrws+kA6PDztVe0SFu5ZIeKHHtHmD8oBAef5EmDrTSnyH5IHRZi+dmX
1fQVmGOwdm8+JovKg4YPxJlN58YtPZ/fNGfMeZdq20II/lCa90c95U/BlMXR
FK3nHyjPErTy3XmEzaSLUqjXeOJgp4zSGmbGw1/4OMs1YkFufk5wxFytMWsm
REYJ3vp/SJzeWVBTtPEWX2/3EH2C52Q/ZDb2biwM5L3e7pOEiO03uZf91Bf6
michFlcyrf8u1+8zkcFdRw1nJW5ipR7XnlwyBX45fjyCbM+iiC9J9jj51VLM
HY5PpyBOBOHkBJ3XogDeVXHFR2B2pHCCPSd+2vcx83X9ZmbfVgAv7M3HELNL
lZQ9rWtNkrdaX2c4nn2/gsPbGCNve4tsWj7KL3OpBPtS0eJvzt2eVYKWFppC
bqX7psHfOtMp8wTTT6N//EblobdMm1Xsvgq8pNTMmAP6wy10GveWKqXKKbFI
h9qq2iv4XcYTP+jxyrqFkZl5WWegdTQDFOsf7wQZQ8D+sUUDbiM6sPFBXhW/
hMe12f7q4lEuO4uSZdycf3iITfNjB37h2MXNvUuE4VRsIXmBWNMjr9YnyMzU
9ZBEojwM19LFuTu6g7UEenb+Fxzukr1nID4Hj5/j2QizgrCY0lVvzLNPoPct
KZZ8qw0z9VgKe6OxywDihv40DIl53BTVA34iYS0iubmjZogjvJ3S4Vzpk09H
59dYyfk59MZ/AS+rn6u6EGA7hMaB5IhGv78KQICNm8RnqmrRytSiPJyumyDY
iIcENnp94tdXYTrDCDsOhoEGDnOLKI9aWGSCMjSUxlPEAXLbZEXBkNCX3Zx+
imr0oI1yobeMARY3MtnHQzC4YQeHAUvCxcaUoGNukoIrM4ZErC94/PvI7xIm
COpOCLg6dN22TM3slkGsVwF7qPkl+LHFmNqgGBlfvR7qr9spFBbPU+5ZrdkM
RI9DhJnAWGWlwn5oueh+HvZJbeWCm2sE3kLtKWb91KsouUfZklZZW8osML9Y
8MeQG6WRqSDmP50kZM3Q41HDHwjni3eANpVian3MmmFkChuPYJ74QPFqBe2X
6+wAfv0xsK01Yl0ic67QghmYG7rVgh+N61rfJPKHipeq8oTFepV4ifWXyBts
E8fY0jykEAi5kqFUQit+cNopfbdBiGv74WdCNjZ0heKHIcII6w/E8KI3J5fc
4SKmVfaoWnjnnTVvogcA7XdXeimEfxbRKpqb2mr8ViJxUe9OjM3+AfCnfy3Y
uqTT7V66ni2CK57ElmwOzrOiEpcyILSxIBEciKtLwNtFQnDejSq2Ld2Ei8t6
xtShJiTfCyrmfZzOn432oZOdygwtQe53CxTvlQOy0jF1Zc1nQYpZfMBLu08+
PZX8ORTzQ+MnJxpqUU2lcwk80XnMksYqdw2M2BtAr8A/JyXZu5hX/bvu3pXg
HF/lvRzPFrd9fBaSDaJQ8McCPWeDG7OnaebhrS+vCsqUxCjR1cfIkCgODkb7
iCjJlPBdL0kf5hODC+XoeheOm1O2VWLhP/A/pPonyAiS4900mpo5kmmxNfIA
Sv9ft+01h5uUuGhtWQJ1cYd+ARnY3q+2UKzEWOjmwE8BDPkREyXXdF6eO/Cn
US9DII124om7bIKgh1nYNWdSdHVR2hwNezpur3EMiJ8sAzeLZgD01Hb+1IpN
ZMx3WmvuedYOEiY3GjlZgro19XUAEU56nEpMuYycco/VudMUFN6Ybq8w/oCn
VP7letiWv2kofu9OyInPBMD+RQZjMpg+NCYdwZqjUg81EzqRI917UiqRjyoI
VZ8VEw+0esKtNS/hSFdZDTg7u961b+zTwwaxTstKxj0lf4Sz0VcKqGZOW5hj
nMoAmYfTDjLjw4JscR7Dy3VTE8nTcQEHctaQMUtvMiJ0b/MMjzVQVC33Kq9s
+gvoKTllj/flmtT5icRBNbExYdflzKxLLDFMcOdomfK9OLrB5zpd0akZuuuF
DQCbx3rueVIDLV1lT4esr0heUB0LU8TeIcrc99gXzSCHdO8i+OCO5hg9zj66
KAsqD5yBlDka6SFHAi6ZECuqXERMFw9s6A1QteH9OLlJm3AZWKboZfNBltkQ
riPV4/yyrq179SEAcJUhmvxeyz0okB7AVzD9jAQuEuWrwdJuzUvG8dICxzh8
zsghuszeS2dzSXxt7i/yueZ30TtZw1k1yON+2YUE4/zqnEnd1XevbHx6vEJY
B0IujrLwkNP4dE2mDkFmnTi+qIOJ1N4HlWd7MbttCRAdVzhbr0uSEVjRAlqI
YrDFRTLPIGVvvLrsqAIogT6N2lnKxBRWp85crLuG444c1jm0AU3JFL8iVkjC
cTjEt6lsKigo9nB/iHH4rb/up9QJDRhF694NTML57xhklwCNQ3FthiZSEKlm
d5R7CTp7TOUkwXCvyvQQYF7ONVKgEzoAUzO8cVbnS6z55XYW/oLENVKbT3Ro
I/rFy6KVih09TrH70Da6u2pWbyzDOX8HNMPFKLh+A/PPUtMNC09OPK70Lsxl
MVL0SD1JkSnj13N7J//fiVhwHwFbDb79RuWsWrPokpZB2WC+XETJR7f1S+nw
Eoa5Mstg5I+4Ooj3EIJ6N7guWH56KjSi8rxuQoKrtVtfUGWZKBbkJ0Ck74Sz
1iVHysem175nvCQKCDroawNbdWbo0SYeVYa6CH5s1XHwuriOw/zJ8m8bhFxc
HzU3u/036GMFjP8JkU+UyotztQyhV4qoJTUPqg0DczBmN7DGCCj+Wicf5SzO
DIo2Jlcjrz8VS+4cwpGOgdFF5609F4MyYLmbnyfNRJZMBdS/yiy5Gbus6rnB
KOzdOGy83Mb4up3T/sPUGGpb4NgrRwkZ7ZlFvew4JQQcNQZMrRm211yZlKGA
2N5EdI2JJ2R8iOEBfZkunvuq40urac4BW6MOTTNzS8LJN2uVd9IrG1H0L4s9
+uUH53UjKZY2lOeCAFVwdTqc7gXms94TJFu2zRXJ6dNnbvv2tVsSnFssrRmq
Sj9OIJ3OJ7uPJz15SpZQUwMyx2/eXhy2tAcbBRpf2ccNnxxKzPvU6/XhDHJl
YosVZep3M+HAkEptdjMNH3WFQKb2dO16JxDx+ixEJOu0/3D0kdQuUIny4q3b
FNJqumI1s4oN6CkERsxFijkFeTyWXNtDLrOoBan6KEnl7uAzNqDTAceLWPsx
NChGJ9DmUByGF19cZEe8WbIFoVshlZK+TII3TvmaEf8YLXrabW9nCLE6gncx
7eHpxhIy2gk1Ytwyq0vrqOO4DCZ9yFQAPnkS1Pg9QnKLqmepo7mxEc1VYkdv
/RMHNLfiBdHI/Wfehla+eKgVe8JaaOLgZU1Qrmsi0VgP0wj9jKDCtdRMxxST
NLeA0lxsOXvGinXyBqrEJpkBrajrNaCkOUVi9oTnDiJ5UhpApzKDwNhQCEdz
DrjyiWdd9NNSjLm7B/8957S+EeDMJ8gRXiNm5GTDGlHpHlj4aQxY7/F+rjlj
5GmhbEb82A2nWNknyqxkv/o8UMJ3PDGRgDTYzmKLEAlYZGe7ne90/ZAD/Mni
rESHcYfmA40haC9fX+jBE6LXWtBWHLQIfdtZQoYG9GdfmhZQLHN8NRb15lHh
BKTr7taswUZbIJ3w2ryIWfpa82t79B5HmpX72pxXbdsB+FdndT12JIYZ667a
Kyeqd9BmVrUntoHvCb0q9aU86cYhyLmOP3rqDhSGTzfRy30nvI1rWw0cu/+B
3AsCO4CznqgtF2+8t/W4E3rbSv6sqFsNpMvYRsX75DEL+O4nO/T8WJTfJwnc
aT82nNU7C/NklB3HnUxVbJxMjt3h17jTHibi00PIR8MqHRgGeClYV/oj2QtR
fYt8G2QihzuZ8cyPoREb9XJSL8NyrcTkroLqpddghPR/GFhnTdb9k8FflUzA
nBW9F8e9/k8tYFj6sOuU72AFVyIcVjxWQWzyzQ6q0CIzRRxsjCAw8wYM6B3b
oDqpLzadwDiFJzOuCW4r98cuGUqa9PkhavhgEVRjkbIubxltbhllcW5hxKXq
cBMg7JMNlw1XILc82c1bKZFeTqp/zHCMPgqQkgy537OLptk0y8Wh5gaJ0JCm
8/fF2Ioq+Xm+5corO/NQoMe7SY4VqBipRzHJOXCM3E2UchzvIM25q/nwo60A
FAPCS/6yBYqGru0iz7qtUkx0+tZvu4ZWel/v1D1Mb1QOifdaoOeP84FCdBGp
W1mf+41XP4686/tUk0M+CPj9DSh4n2HYERXPPPZ8Iu4DskyqApsj5vJop+4v
NUKEeircgYo2icblAqF6O8cHg8bRgz2MJG/LsPDSI2hmQcc+oCotbdYr8V1p
NUTCZbWIPhnPPgJzeA3kDHOe4pfkBsVlt8OYC1URik+KSvzOOqd5Q4G+oz63
SKJ4VV/hM8wH4l5fY5+FzAYtPcAgAxJbNLsdmidM9JFuo3jWuFKT2zhDQruq
1Wq5WpVMZZN9u1cwJj7PWlCh5/WNBMxxNXZ7Qrc+KVKvPiU7dpxfonzx3Hpv
g4NXgdjYu79wiV+npHGOskLdT9xFabfNjFGd2J2/TqxxoJAw+Pykf8aIweMV
HFApb8Zgquj6m7yRwcjKALR+XhhFaumjiJCOGGczAAonMJ6E+eKk5gIF7OQ+
OioVX1Db+FNiKmwlupB2mbl7FKeJaG0ryn2ezXaLP5s4bMZ2IuSf6PJ3vro3
QpQSxPjd42caXiia4HhMHfLXTx0CqrQb7789Va7mx73jp2DiL6zfJnQyUqlY
vbDCorSSp4/VkU/NRfsBDlN3o7sSzgzRjZbhH2lC/MJtcXUa1+jJe+s7QR4F
d3ufroWXzP6mTTBA4/4V4TyRSJZYNUMIEIv+0gEyOYPt5w3uvIywa+50Vrcd
PwLJjo1EQBnbn5e3AT6vQ64zlYJ36g5K0S8s3urw//CxPv+FEICGlQWZltZb
/nNvoBl2k0CZL+9+SuW48uwRbZDGerWmmW4N2VppG7NbIjsJnt2PEQpwP8+n
pjETSIXGf1THCJEbU3sx7/HDJLnoQVQM8dnlFEXWhFeCStNFiF/VCblF7SH3
Rh23ow3lVH+EhQi31LIVrzL88+hBfZTwH/HmtVHb3Z8U74IewBCxLArMFSI1
6YDY/px/q3lCs/enqXdhpI2/67J6l1z/I7ZzhE4MXeXLFqJ70webFmrV/FbK
P/0L/4itLXc83u2GcQ/6Qush/EylIxRI8iQ4Sv4MnCnj/tmSBnEaqt7wIxqB
d+HwIu91ANbEGfukYXzTupPrZNnJN9GlznllmUne08v2RLfeYAjo+Qo7wCLq
N2dgUpGO6GSNBUUtPM5ANhsN3AqpmhDW17AH8J/fMKahBXlik/mxWcHII2tB
vdYgjzx5OsS1/Co0s4Vvgsq5oBDP0Q3S6tUA1tS7ecHi4usccVf+hOIStrOE
PctY4GeAglgW1U5cuVyq62TRSrlSxXCRKpFskoLTQGeh0fyejmZ5CY/M0zps
qD8vZdV6lHhUPym3fshpIuZHRH2Fy62XsnmOe3TrrD/iPyua+RHKZsfQYFxU
IKpbkW99EwAH92ob3vL7bWZEqAans1qcvMd8CQUgRS1yAoFXG7swQXcUQo1+
OdGcxIndb9MEP/4b9XCBTxwSf4FDwP/5clyZL5XCxWr4GvNIRw8/G9ANjDzx
wyluwWkWmN5bkx7+mhMZUo87bzWSh7mmJ9iGr9chtqD1KEE6ZuZJLuGTgiv9
ScZslRLYVm0flghxoJVv6bnw9fe8tLn7h+5nT6bt7XNyRj5ajtiDRJ1bmjQa
dUzEBEJ7piWNvJmdUQI4Qcj7PvODk3kj5rx0mNLzD7vKRVynB1DyVGPKFNRv
S/6Q6U6GZqFFOEGiM0EcE7+gi9TpToXBt0rsC3QJ1RB8nQ8V3RLD/cB5K9iU
ys8/0EpCuf8KUsodlMQk+SDpZ3ZJ6g4i6LqVQI7DFCBcRxaZbldLqlz7uF4w
TB5A4mkZsteAjxHncb7anw0T5rjr05NpfdQGNzDt96+SMs0WGe/NP3cSXqxO
0NmucgaH71/JnGFxg5GkDy72nnGNj2LcK2TZhM/j6PZLGz4imeIqADkIc4mq
EBuj4YgehYXkIwblDd3boZLBjmcK6XBZ8wQHjVYdrvj1N8Ov+ReP+Yb5aBpQ
TF31KE23LM1XGEkHBNghKgvzY5kBc/86VE1bRtMAslELEJ1JqOZDGXRMn94O
s4Zfjs6Bi6fVCzQGvXxeyRdxCaDscLqHIeed2tiHp8QwWAhJE3/ZzALmPifc
mlyZ8fh2N6yz3O+EWUQEqrrUpkuXjw+9es241SPWEm71Iyagw+WXKXx2DLZd
kyjM+OcbUvEZKM28oVBwi25bAoAf5J5j3okcT3L6q5pWYhrTHH+rakuCjdgl
B9iyJJEdgBrbW+eUUcFH2z8LxYUX8IVs58c8GYgkNdLlfGpr7SdutYWtOa5B
zoH6RiNrwmVGOR5NIEXLRhEgDW1JU27CXW2NvMPxB4ZBhrVVKBTeRNRvU/dH
HwhNdmEeeNXG9TFGuhGHcjKb4bmoPmUpQ8w6067YqmX3c7+dVSL+R4Fm/mpw
sz0HauN35l+QI+dS+4IPCnWVXDN/aRT516v5b2OtgJzAhHl6oqY18yibbjom
dU3OFfuu0u3SDUeCkGtfiSRJqtGAlB+wkgs/6LoephtlNHkD3nIhjQAXr7zS
/MJfiqKyAH7vC7Idci5n0T1E0j4v+T8833rTzs5hqhB2l9wTkv123ELeq92W
UDsI43agPCwrGzua08+sVVlnyMrDClnw4eAtyF7xyy7ieubpQYhr5F1asIjA
R+KOf3AxYzWGTUqCaI4WuZszUM55v6K5HAPysx+F/EcFuLaqEgFChN0K2D7q
veGLxDJ1dvcoKJ8wm3XcdeuCz/pCYpi2bF9vMFCzhd9mruydAtdXK2JoL1QE
MQemM4hLukTq3GqT85hINj/hCYPI1rOPPPU2yJPUu7SOBRYS1ejCMzF2Ewdq
PB70NZpi6qPn8FyN0Cg9xcf8pkZr05u9kMmEMKLOuUJ1U9Kt1yHiPkXT2lL9
0CVpI5Wf9QcCY+8H8Gg8JuOb7qdJRmq4+frQFhz3Md9/ReGWZRLdOxds6TKG
fswGMFVB5CtIMeiZdF1up0Zz5DbmPFavGWfu7Cfb+67HB9ew0bvXox4XA1iF
mJQDh7zXPhZR1QslfDyZXpgdOmpTmH7JMt/tSjKlo5+Yoli1fIbUX58PvOYj
Fo+DftQajraDOzrXPpr2ko9dzOPngIR0kl6w68m5FWHPDilfugV6s+O8CxUI
T9yvxxE8QT727fl8s6WV13t7FFOjfzcZkLwBbtN1oUbloVQTyB+DC3TrUlwt
9nv6GAkIYCj7aLXyPV2RIsW9noDgW4zUbihkSx5iN8aaiHyeRtb9WhoD760y
qxmiGW6nriifpqn1ivOK29brs/3MuFfq4+Fb3zD+e4gXcWVqrA4Ls0DHDBzB
/jGWB1IDESjrb8RJpeg9eTaCfRxzDCaEUvMA6iuzU0ExXZorhQ2sTuZ0mP8i
L0pp6gG7AEhiPE2CmUZ2Y6rIQzQYNGZDGDczNw/fPkzTTdCbwIn5tCqnJMVN
0KYRGzJIU1r1cDOUmkszMSpOuf4U5uzSlgnBhhMFVwC/jhbDq6ZQxVlFziBR
oPCeZVVnLQ5yrOqe/VgczIRCF9Nc3bx3+O1m8anuDJXT/LogrrgupNaUaHuy
vyAEfqmkABAfIxiT0CyChgUe9YFTGY39qPbFq9DduToTIrLDsTKStfTBo4IX
/x3xfbE/ALcZO/2eHOVECDsBIbD03HlQDJHL1SJVkGD5gMUQjAnpj+yyDald
v/5VVGfTZWeE3BXuQsrH7qcSf9PgvJ/Z8I3eZGj1KBqhd+2LmrG2Rx5e26xM
5SBhICFSS9Hu0PBOyeelpDjbEpnBIO3KJo7LiI+rCT4+NYWRuGxyuSxU5Ktq
J9cNosBzUxyYPGIYff2SfYckc6gn9rSPpnHWu+mkT9/LA7YyzsGKuA9TVMR9
1+GIkGBQmhH3HO32/kAv9XJkMo+B6mRxjSvakZyOPAb0GxqDI58EE45oTUWc
aSbB7SlqJKt8bHfxPkhrgWU+E/El6KN8gtGDHZHPVD6egXJfnA23pfbd88nc
2FejFYzIImhuRWnU/kTYVRVjrbg5x+llRjvDwF7eaDRW4IevfhDvQUdHVxaf
uXMDyuna5bxAAkZPkfaqfKWWxThTBsnKE2uKqYMAoJwTzgNBNSffba4UtZwR
680CeYU01kImaLaBz+g2FAyYJ/WPF8cX61HONrg5ouGh1TQ+fsxIMjuMmJaC
xE5Q3jp+q/ulZOPz1a2r/RL9hzCZANley7NJx7HseKBlnfYvpeBOQkjsy4f5
dNefAhZ9Z0ccTIxL0c0uqE6uPh6zSYoWXYwG9Z2xOhLnwraaXY0a3D1KAjlT
dDAkZmdiXorgfDP4yYOvEoKo7XCBptM1pJ4NSmOs2PvyE7kGPX2vBIMyS4Pn
e0UG0LaBp+VYao1Ge72gjuJgEDNSPVsKhJ0tDYGluRSMjzIxzcGrG4wReEOt
EltVmv0/8D1UOFp8xOFOoSeaBMC4AtcuY3thXimPgP+B4sVoJalgZjt23oYn
Xmyhi7pd614pf2maWvdCBJCDw3bp2mKV59jWa/fyH9J3vT/CpggJhHTNWD3R
SoLDIGfjCQW3PzpCzp5tdDuxqogXiKPfO7C+pEbKbbV2B0PGsn8rYvAV5iox
59d3aP9pVLyl9o8RBNMO9zHBUxx/jVpuwiOgaapJEKSthYH/p8Q7BGuwd/Zy
oSnnttXqRJKJX72QGY3QlMaU2ZTtIqOr/99MKgtDuA4f/Qod2mdBtsk/6anT
avvr4iWePsoTBMGaxx+pLdbaXiApKkg8hBmE1zRsSth5YwDjJFA4x5svtCdf
fH75QX8/QVbFaTA2lIo8uRvC0Zf2Y78h6LPxtucLXVnGUtfKcaSXKlQ01wIp
kVQpQI65AcaxGcgheIqRscVYPGGac+mafkYXuQzTQOV3WZZwLTVaUp1FqzAv
FnTwsbooIVFfvEc9+Z3foADMDePtSJNKP029dektanXtuqzAmURZnGpcybsL
KLlwsfE2+17w7/F1ciPsgwspMHS7tWPHmLcZsmAgVEnSK1ivTNaaEXmWZDXE
ydx2Av/nZ5y2/UtrgaaH5A1Yu6dnFF9IgYMIatBIH+lQX+AVDO4WtIZp0UMo
+PIVyeaPRpAkwB/tK7J4dY/jL3v71j4ZHFJHuWGED2FvvQ/xttHHmd9EFFX1
aW46xNxbQd6tqETClaerkBUUcFv09I5nDPdQTW1fW3jHDAoC4d1NyETXNsJh
+aYnNdK8gsXeVX6Pi8qKKtNBYuWS9yNQMCdkJQRpFSlHRC2LwcCvjuddQBQh
r3sG7jhzgDj+WqI70itv/xJpQCb88THGlWZdtLpyhDKmo5PD/EmVe31P3WxT
Eam9ElT9+uDjqaiR70iVhcPeFvEOURswIlAuzS3qBKt4ZD1yyQSy3CoLbztU
DncucBT1KLDBVRTogwYofIg2MnTLpPCzjO0zRFuTmsGZF/u4/RHpQgRYLo6W
kDsnZdAvn6gCjp8ud8dPZdEBCccJgq4DnqFVLXn0UXTvVDyUsfL0c1UvlDor
v4dibdA1pHqycdvlslrOqNhue81TdyfmibxW5Th1nMH05HKwHj/iJo++c7Ym
A0Csgdm7DognFkfhYSlfI774P2sd7c4RAaTx6mTKF1jtDpWvv3mEvNuE39X3
k3eVLKWKFpc5ErqFjfBFzwCH1HipHrowRauIhGsVtk686ifbMf0P2kF6BtGr
ogLms2TD9fQ/cExVcHIQcZIA6s58FdSaStrQVcqiCS+UB6ajMDsMqVJTZ/Ae
YoB5n5pV4VTTrMwYE+4AcGL2iugBrnG2ikfPcVMY5P1iSUNRxQDRG1pJ7FUB
bqWNkDenPF2lI4iDHWeHLxpubOBbrcoo05jqAFwCAD7A+2oxHM6h2JSVkqKc
5PRhTECOUmYPZUlpJuOwAWVNM4+xQtr2v8I1+CbhTU0TiQjpg96ylSLqcz+h
NymOEcgEo3CjoLkZWPfFGyd9D6w1UchJ51qV3a0c20pvgazWKVd0lh/zKWnY
1DHnUQgDaEVF//F1RBTuMRKwQeipqGynd7q4N9DTpEJL7MiZxtGR7hAm7wr8
+y7c79tzVHT5hKZxyIoL9ofnvmhK0VW10ia3/14UvNlaJygJloSUTCdjAYU6
9FnHh0IZ3qJTW0fUZpUM+Ytmx+eW9/JrrCh1ufKtYv2IOxpbR89DW0jrU2dX
tadGbySYEOmMiOrZYt80FdSSkUEBhrQDduEGfl/2tsoGn8Dz1q5OSRFx6fP7
XP2a5ZjjQl/QPDG9Z1JFVlDjfOkCdB9QqnlQwHtTjuB4vJUSWnZ4U0a5zcg+
Of1cLnPqfZhSlM2IJr4xPrxwPg54WeOnsDGX7N+QJio9XFQNAjjKUT3YJkMU
9osRmIolv6FCWdWH94ge2gSVePF8XTqJANRRMBsm8pkncaChY1XVONUNyThA
NeV5ASID5J5qhYR9/91xUqAgQlLuYg9FshUXI4Em8yUWgVH26aH1y1b40ciJ
555eod9oLgvoNtYraQnpfjfS3PWuYhkBHXZpITrfwkE/AjtVmNBq5jN7Ia2P
uolfCNzNndSn63oBT/r7c220KZfET+162qPo1V7mU/FAw2YIa5SjsbxgP/UL
7R0ufsNLj2aQnZp6BMlZKdvqq5aNcgrSv1AnXsrouL0eqGKnZ50zxTHTH7yc
R5yLrkGmpnVkZUoZEnKwmmGhHzIlUxfBwlo79vHtP2+X2XV4pHa55SmZPqMx
nJ/7uHp4qTnl++Y+9wXmYtbhh6rQP78/iYT2c+vV6YXoZGK3KU6S28XC2w+m
pCHCLMrktKbhkdWVglne/NOXk7uXTVhoSgkly9Ws/+Tkm0yiVXszBw28E+Y0
oD6tse5EwUzDZd7MRRr1aDQ4jqblOVOk71bOqqPJjjRrv2SpYrsuV5s6LsnL
1yLSXby7QEs2+8ypHEqBFhvc43sMHQDoRmSnxmLSAlBIBc82jSmTANNEnjwu
u9vvZVVSXu3xDQAe/d4MHV8evoi9paDYx/qOHMFLR0NxKZDHEVChymQ/U+QR
hfZGY5oVkefqvKFbPCt1JTyIxJByeJ0Gh/P8xfC3UJ2Pw831/6UCEspEP7cF
pOhb/TNDepm5Gdn1BdtRIzlDEgUCUxlVjeX6mNkNlStg2jABVNYOzzK0H1Cs
NIMwAC+lU3RH+bquTHjQjwK01w9sUypm9hmMhEJZnwLwjU632HodO73PYqS2
p8qmyDBvzoYg9bL8q5RZDGzh84LVr3qnKbThuUI7hMLHnDukDSxf88HFXRvw
hhWM4uaWt59Gt+NqGSIGIC72xyrDjgNXX9peqDSL3wKpcJSmPvQ4wpCgZoGi
CM1Pn7kjyabXg4xp7QtDS/7nhH85OEnUu8XGDeON5hDvMSq4RNsuexji/s7r
th4q4lUF/tcptGsR7CjLhotIQRiU94X03vEHjCKJqQia3l/vIK8TkzFhVkbe
sG0WIhn5qaEHsVor9Lzlq2u8FuVd4yKd+d0LpdML0aOVzNFGXVuIN3ddNT45
tWg3LzFhrGm/TYurdNmwnuIy9Ljuh+9+Uj8xh4zd328y+aMbSEqzvGMB0eyJ
Tdzlcp9py3ZuuBV089iHEHpaWULyNh4w019pqIBSeRW+vWDPYP0CPO1KRm+8
DX8l5vF98z/xK/l73Hk5JFB7ujJOZdXvfJKzO692HvXbHXo5QULQEwJ2HwWT
hyFkUHi6Xoqc4rDAAsYPVFbf/078n6ALUyUfCv1JVsMncmyZ16NYvBF7AK3v
UX52ad+zjipUYM+WQ0nvVjlzkQ+RXyLPyR21LD5rjuE/PMcRDJ9RXAu/RrNQ
JpPsoLzYlF8f/B0dXY0ERojYnz04VhYa+PUmEEiujUkSdZk6G9OUZVTXkSzn
Io6U76AZnH0ct42TrfkfuHR8JCCj5dfszBGcfV/oHcvFyQsqyIaK9BaF6By+
ZJQcgYJ/WQOLflb79dk7+Uyicrim9EHOH8DzcH5y6mS5IWvilrMorLRCT/qE
8LCDT7Oc/ur3rXKfIeFKCr3YRIFkzA+BNces2LVAhCIQY8McrdvtC+KabrER
Mo6d7Fwtlgf03CCKW3wh/7F79TCQN9GzkgSDpCzy0tIcmhFcWSgDa2Rbpi4u
8N3yypYKTpUgXedK4Y81nIjSSHmVPVn1LzFw/Qhk3foTgv3hb3KjVUpo/85z
zitZLcF3X8Bd4Cn8bgplmS4KAg3HVs3iZjHfcsTaVnPJmrsYW2zRNYChWoyj
GFRFSwUoDpkHCsqL7N8aCz3DHRQaIbWKecYLtYd8qsxp2Jg2qwziZYlMICLx
00ogQqRTJ72YGwwzCjDkSB3y9hvp25OlMnYGKj642YO1jxG+dC57LZ5O8pGi
TKaI2xlAuqR1KHt/XNReiofQONnrxwo3lxXXM7tzQQTD6X3tsOxQ8GPkT9wt
sMBGzPc1RTWAJOHp7PSpyYiTwEvzVwt/OTtX7/932rrkHXKf7e//DOBv1Zal
+XLEeyi9JlbKcqXQcqI0Cvy6/DJ2hadu/dYrmElmnbVxrTGZ0E08j35++b3U
GV6+APV9U8RPj7zqtGnsbMEFMe7ZpNpf2vkwuEmvCoD3wQMTKorTXcmUqu45
t4XAtHA6GVEdbC2MQCfU4r7ZNgRvcKbqFoCZ/4G6wYQNK0Im4g+Pvt+52SsM
pnbrCmtboRyeD07RQXksvVnCI9SrsjRVqyoApbe8zE702eeKcLiKBoF/TY0n
QOrqyCdr19zlx1xql+LBlsAvCdukwmJlzNOsTg6hYQiWef0u8VdzB+0PgGKv
jqkuBOqyUU/b2ASFUu/AVKUtvu7Qcguz4iAle7QmuxPPocBHQYb6PW6TxOr/
aAk58b8WuOTH1LDuWWgiCSt8Fn0uQ/aiwg1YvAA2dcr4QEGMaiuuSgGjdOGs
BlNpsSRlv5CxKoKhsj4zWH/DQ8ajhq3XtFVM+vDgULlrbJ1Fm3RoMerE4Dps
fY3qvE1pPcd8DzTyTsb8+VOBAg9xUjEcEk+aD+5QDSO2lZlWx8mAJvKl5O3F
Yr7k5K0/N4HqRertjmI9aLEMjME/zKAfEcS6Rvo896rQHhkTH3q738QJ6a2R
dSfXN4lbHWsbudxSIDFvaAyRqLBIb7yaWGjqwWxk2cYO7Mv03OzG0Xgp6Qn3
6/mCH2MybGP2k2AAMO196TseLJoFZgJpHFQyJG7CCfkTzdcvJUS+sJG0DrxY
VrBXpBNDHvRMF12RiFiCiDMIiaYLWZdw45BmJ1tZCxdK/oMLVr1s9F+NwiAJ
qqp/DIi4MHUuFn+t3x/yKNXQlJ3w8uLiMFWnAVrSGN4oUqPxJvO/J8ZXFH3O
C8UqruiQcI5/pmK6f3AV6nsdhs9dGbTnnz/ry8cRod4OXu22Jitdj8xJLut2
BJ2QQ0JcESeTPAkyIan3DEYqZg9wuxcOZUwzrIHAKgPQn7WHq0I+lpgpPY9h
HT5k9HiQDpsO1azibXnhXu4tN6oPPS5gqqSyFDrf0kXMjCjjLu/vcIxzoeVt
FLBnGdCVnMygCAFQugBOy6bJX7P1oHgm5VAJkivPVtgCsKpMwmnUvm0fWFU/
eM4dNA2WArlhwn9kQzlpNZmUBJYraYHSfDnVU5EXPVne5/B+WglVCk3knJj5
w+PjYGHD6PSswuXIwrPK8eTw0v80xZZqBs2O1XVqgegu5z/ogbJhqYBMPwNL
CcMjnRmcLt4nCHiHgZxtP9wCXypy085c7V6e7lmnyoBbrOfcbBbtrZqBQmI6
I4KVrz5D3bHdJGlLCzHAfpBuydJT4s6C7lWS3X0frbKSNtx/9oYsxtiv/kyw
r4XolBqfHTXkNNae6h2BGvhryZVukjTqUwvL0DiX1xy3qMhrsnlI2ZXcmLnm
mAc9sUPetKtRW3sbDWdJTbuPwHX+JVMKLMU21wH6Jys5WThvNSlwhxxPoEJa
cKgLQ3xCnf8/7KTIG+DclmCKdcGswFhulqBVpRc4iL5B9d593NSgZMQmreab
NwnnaMUqQxb/QkUrhvPbxxNi6YgRpdaPxNk35DZ3nVH2eHX/mnicjiy3WS7Q
xPNS4krxC5vnOCpIPpxEmUy+DwcHgq0KD5+BOCbQG3TyY1/5PCxz+Q/PjpmY
z+wJiFbjqaaee3UJdZ+fnXI77XACZi6VkuC9Ij3huzCI+QqihczV3ali9NXc
T3m5T6V0SsoVXkxhLs9aQp4zc5UxPJR6hxcVoa4ahunmEglO9uYMEn4XkKNT
+0Ee48c0kGp2si/IEDgX7S6F3PYm5Er0D0jGNLkrYQnDbc5mWDcelfeFwPP3
3v19Whge4q3XdgGyWgye890otw+eMkKy/XPwOfM5589jl089YX6xVJZEDa9D
fwYqYL8HPCEXSEuz5afFGfTSDVSEKOZBiKOXWcAi7/vLXsknu4fN/ormMBPN
fIZ6yrNC2GWbVUa8TVDuXQH6IWvtwKTvoXiBJfQHcCEB4/ymc0JpH2DdnpCM
rhd9XfDMFJgNtOPAlTpVfiUq5sSL5cytIwVQYH/kJ0fjP7++HEtdOaEgeWsb
14kkGfdQdjg9VOEm2GuDR1tPpCYODhAruf6zXVbnI2Ra0NEi81k5XzQGq54R
l7ZhBxoO1F7C9xwXzoxuxifbzUMnWokgY1zOmAP1SPdR0rcIfE5KPIFO+KU3
8c1ri7q8klBipBfVimDBr7TrOYwknd86MC911YDZqOqC/UQ93rjhyPVvN5ZT
oUpWo5/37tuGcC35PnVFGgT+c1xuUDIAwoWZzuvedSHezB4JCJhjWAJ0eXVY
dW3ADzFAmE2E9kLvHtpHM4p7Au0UxgmSWRnPs+tHItgt6HfErHQqNJ/X+DgD
+9VVCdTflcRAKsdIUjKrpGWMZmjCe2kn+zJ8ft7AmHRj+MuxgzNzuCaxdAaC
LezW2gMFEqvtYvh8JXsiRtvDHWxVZHMkMi/TkEmy+V/qz3EROrNHxqi2JqB4
vO4zWWXjtBI5M6sS1ueYZwmr4T2e92f1r+6864KOdDm/NlWQzpE8gWXM6y+i
0OBuGAZmJC4GzHZ5LnWeACXrNY0yLTaSuNrINHU7DQ2u1Z0MqIGFpFSoob7W
uakZQxOj5vU0GvO2UH+w0lPoWJ/7A8jL9sHkjADnLf7zLqaC9eZb5++O/1Ab
vmp2Xl+QSpXh+3wff35OmkQoaH/b9jJ1J8tKy8fjvTFqXU/fkFmSWD86HYcY
QeqlO3v1ZsS20qCLodjUBri+aloagDVGk1x5BjzPwANpCOVn1yIRHza+0NQE
QtIeQRvBdZwJ7slDnD4NZg0QhH0ddEuVBqAqGH4HOJFWRTtRZKUokN4yIDX4
A+GFNgBAs5LxL/x4sVSxMgyDj5GWIDRjsYNN00RlGEKh/P6blMLJMT8o1I3N
IgFN5qleUeWNNnuxQ5ZKRujH21M6X3pHv8xRrhlzHKUML4AzWInDLYb337Bk
2fk2JF1FW8SMC619TMa0EEXeYIBWh27T6rmxOcQe5wBcAsp2H0Fd0ilTDvhG
OiEcejQHju4nf2OVeGgP23QXCBQqr9NtPjnvI7QZb/Z5VooxKD8Wqlb8E9Ul
wqpSbNW0PkODZyRi5SVuy3vbTr+cesj2I6X9IHri4UGkDlqf3R9Q/x8wMV7M
rrMV/OKs58s23VLY83WYKtBGOM8h7ESS1THv/tvMQ2bJC7b9st+iR329WmJI
gZe20VbLQXUgTuNQWa8n30ew5AgKd6zgaBLXf30KgBc16w9MOiYFoGqOnYfe
8VGPCUz1FHzwUsXw5vEIQ4WnCZZuYDED3xnRwb6J7LKEqr/dXi3EKZdgLpUQ
Naodc6lzL5dJOMjnJXz7t8cT0lVC/eCR5Qgy/XRWHqFwFpwlqT93hFHNIlZO
nGjnj+El1s/X/hfAcu1mJAfqB/XA6lnwkfLsRBLUJobn3NkgoqBJjwBCdpOt
DG4SI0hrRo2dDb6LTrqJUXwAu/lgBslnIffBsoKEEZFrqif8xaS9Ciswkxsf
+tLL4c5IvBHZ7kU8Rk1f22YbyHlw13j4TXdghfNYgtkwVjD9XxV1/rvraZwp
TtKqWxVNcCAy1Ic3ihSfCHb4xsszciNFpt2RZczNdq6QTUg2wyv7SgFfygnQ
2jnWBvcXv7cCAXGHI6Snafiir0uv1r4bMzYOH1JVF/e8ZUy4L1Wts0mtyRkE
22VHBE0oKHQZ7D2M6NQkRRsU134uVCsJoDa8nwX4tMA7WEafsjzjP/xthTx4
eVawKpTSYGSsu4jl2/EQiO1oK34eDk25NC+xRwtRjtCgd3+q4MkUAxKm45u0
vfo3+4powHNvATQFE7k5CoRNcuN4i5/dziONePO7DNPe9qUBIwcgCmnSRC44
EviX4klOX5BzETiAE7804a0Qq1xzRlhKjMo5lqb9NUbgNare/N7yfVAJvBzP
MiC9f/gZC5hmgSXNth1h4dnSfTASH9Cv7TTU23S6SHYcf5cCqBweAaeik2/1
IXq0G1pJqK7c3e+77WBgE5TRW2N/3ibSOKF82XSDgKl1fAS6HL+CsgPI22uK
KGuzUeeH8QanFYG5fxMbqG5I4DiFDzLh96Jwhfd6NJjkRXW0Z0uUHdPzUGGN
TeKBUI5xaGWZfSPdH5VoX7eml+1FfllFT0wAxIc4gtlzqCtrho4bUSuezdrN
gIRaQYHeDyNn1fI0xePly4WRtYXXDO7VJ5SErgOk5nAvV6bWQdCVzAoeA2/T
RxpPWePuhMoDOVaD20dhOD1Eog8FaJbyG5mjVpYNFvt3kzrHU80CbdGSKoz4
EmRQMmDyQdIuOJ4NkehXLn1eLhXQSAonooYar75czy8zif3TWFcjKLoFA4Ku
oikFqnPsH2ggzp/+bcPnXjVuFCAwZBHz+PwL3s8OW8F1OXuzLy2MymfPcxiV
tmc3I5qiwFhwPO2F7ahFLLweXqNAN5nAcVeLckFfv18uMYHFBAQrfliesBh9
ScPlkiDP35pHX/2fVUPk5fkhJqcjKi1fXRyCCirtstGtT53xWUvcbTi+kM60
QE2zo3fzuEOjY2ICU4etOIXGjfZYsmFBhzI2peWf5YcKWW4MAO0r043kEnKV
m+o65YzEV2/XT73edJh29ocgUEhEEIDa7ryHYyWV2PYqg6DewD6KumZBaThk
tLHC+KIJ/A/mmcTnki8ZHRYq4tOtHQjEO7phGiMeqL6stT+Ohl/d/ItNtnv4
HvUYtTjgqKtVs1YTweyuwFu6oXib5mCOWqwzPglHAivcOMI/HXXzr5AU8LwB
yXgYCTz3m1mxdlgTLuaRdTqGcJLrTG6YE9z9ChcW8Gt+FTQx2CM+7HOpytGr
/gFWLVdKmzRX6Jwv/33sTKqjZ/tDaVWqrSkl11jUfhxTPDDoK+64D3463l8x
8X+OKssAMlB8pdQ5lPocrrfp7WibezS/ik1gQCtT7fUK0TVNU7ls4tmYgHUS
qcZDOGGjq3lvvvcpJ+FvtDI274r+OXu7gmHwlfyqPujNy3NE3UXY4uwZGXfF
WhZ9ikB+JnU3BpgAOwHikTJMCI/vQNwfkvOxlUfmypm+HDwNik61J635AgBN
vBK6ahg6JkFzgYjhXYT2tVuPoseyCPVbshwRl7JvqBvvuccY6E1/iIMfK/xh
476lOcZPbuz5tfMTmAvqOCkzvhWUr2+FmJNHqQEY79qZcygk0Azy2xcFnGcs
wEDAaZ1kSJz+pbKTnXW+iEB3MhHTGKolLAcQfB4hhy7KzU+tP5mvqfiyOPNh
/CrnZYo+MuzIyV6KVQnHO1MRrPMClPQ0lEf+Q31TiXZ4XCU1TH1rVLgjF8ST
Oe4xzeK7/lGnaTsuniXSSoobBtdqECt5T4po/s56Z9/H81pyuonktFi0TY7i
in/MbpqI32xzLV3LlZQMRdpCyfV1m3kgTPG6iXuJpBa4r1yDvWa+RB4nCzi7
g+SyjD2ErUZB8MMCUL09wQ/p9K3HBHLQgusT1sr8f+GykVWT1+FGiq6wXR7r
t1sN/4wjKmW6jN00ziQS5oCg3OrN0xXhNGiFNGdZJwLqIk8d254ahBranVcR
OHHLHidDA15cr353YuEHABNTOAYTJeYSDVv3rbJ+zD6snP9aXzLExNhr8ZCG
vmrq2j4c7WyyOURLdpmKZ6VXJtMqjAJixnlRBl8OV21775ETZRs61KHZogoQ
AO/iR3jDWuDKhiMmY13dz4KDp8jOdZp1dsNFiUNfvfCr8aHeZFGjyH3ijMdG
zunwSS7D5B/XSSluwNhYPszAuEAWervaKmJLy1CR/GXHpET0FAMHRJKI9j8G
K1RX208Z/hgmx8qIR1mxgC2qMoL6gG/0STgKpjCobb8e3EW2ChQ1Auud+CKX
ruoHSQhE7qpMJn4et87OZ7LzPA20X9CKUHr/Bq2/r07AeEIr/Spp+83X/SoN
wEgmwH0pzAsnk/b9IbO4Ov8sejZY2MQCB0jgBMDQAVafg3IO5PSj1fqQaS8T
PaTx7DSEq2ML6eTFEOEoucqg1LQynogDUiEVD+nOtzVejuhlso0x1ERJ7q24
sI7FBLJym69FDo6vcqGDV8kdZCft47dJpfqyB/aLH/jN4Ldr59pHbXHocuet
zy+q1B762BLtPm1qfY0bN0mfubheylGRlur+4JcB+Q+RnHk/zFiAoVO/mJtO
athxMDqtvwuKG+xcwrNX2q5+so5v0invAA69XfoSKqd20j5SSALt0X0k+p9L
l2grd8CfWJ4sS2TWOGCAhJmHc5/YlfWSPpYznYHwdPK104IoqtZEGVAdYQey
RrSIr4IzNJpXHxaS+loKKOu3/deEHg013GMf1oyUA2xz7RinnlL/SLTZ66uY
QqAJQadRi881LLcIXYdZz9jzF1uqhkVNvN5fNE6BfmQZLgse65rbLUFqeAeQ
Gg7UqpCQRX/7CkZ2Lhv4R0P5PBrpEh8pZbq6nyi+pB86V/n++cdQTprbk3Mt
SrPmcTZWQL2hLASXkgiaJw84mLjnECnyeNhMw/3vBvlgUIOlRlJzTWr28dYk
V/4YOEd9VdDI8JaNeD9tVogIUSVV3SB0miOwQ8XN+U82b6GDNYnGo2HeNGFQ
FdxQB1h7GgIAO7a0Ai0yjkRvYpTzF8XwlSyUMrBVnHGgsoWRY4qhcWwtA1cf
IQvYujGDVB+8HM4eI1BF8vMKGp3lPrzkVzvx4xVM+C4c1pqAVAys+n7IbHW+
3/2rNgmzUbFAeiAMXGDhGz6NpmnaEQMZZfUYXZY4x6En6RdiJRdcTJ1XOPEJ
0i+s4DWzlepuBDH80nuvSQtFrtRBjOVv5tzDPi55qVuqfoHE4ld/KOIEq0QS
vc/TSbF+1GmvxuJmedP6/662qcynASHc4A1aAwTGEM+j+lNXQlvsCnWbPBNo
vTOG0lUc5DbWJn3haxLh2+mlc33yHXX8ccfK62WR6ygPSFdJwIJG2aveXRkP
8VFqM5yDlEbfFqaphuVbREs5Rlvlnd+MMM2PPgJZX1JuT3ZxpK2iAP6Av8HG
s2jIdqN4jQB1OdDYj4dE2coQK25EP5CkDyCFbWkMlz+yXvs1VcfYrYr/Next
1y+am76i/BVm6C97xV/TG+xRV920NrDmJAPXgiEdGRgEmXCidk5Pv3uhsz6B
zHYYMM4ZXJdxR/13IolQKSgULV0RGmBepkAymctwMfqf6j8RSeUzcB7Jn/1U
o5ltQQQOvYlezacyNbFKNuufhxqSTykxQ/KsfQkI35dLHGXl1oHb5ZjFxwn0
X5IpYcE+Ee2kizmqGjW7SaWSSk0W039O0HHjpR5dlCXTLvo+HSIcUy4LM5/o
/K2XdGCINZTN9HUYxN/khYH7I+lnd/3+v5s+95CHelYdv8wCBuY4sY41cQbp
ustgrNKnr8sKvgmZ8AfrGtuVmocm7pDMcv/XS3wXVJypjJmt0K7dhfRzjuv6
tRcjJJeIJML9gQ/gKMmxRPrl4RaLoz0yq1Zosfy/n35XFPwjzYzW+a3XuZMD
JpHS7KJTvF82rBaIpfGhww2zXoRiT9h4t/lqqhTprRLKd82sDQ4i31+FsCrL
Fb56fUxyGPm7I4OBeDAGjSL36gu36Ks6qbwBwbzEtWScO+th54QfAljgAN1C
SDhc5mIzUmi4b6NEgxASiKx9ItA5fi6z7LtHPdv8+tMXKQqoAP3Edx0kiWwK
Eh6ysNmxPgLuo3o1+6/jQ9sc1lPjcD/g+A+tUpVgcJHm8GdV96+Y9LwYJGCJ
T90RPtoK3ZBiHA16O9JcsHl57E/qPBgp//L9sBcIBveq1wtkGKc/f/jdzeFi
wdztk+r3SQFf71Eg5l9IsxjgiwtI23WYVIETD94nzRkY3Znf7Sy1oRoU2atj
pfdgmL3knpU7kqhmMgrsRFTTKDfNVfTKR9QR4VqaTZjgFzD4TyvsKw6qNCgD
JzucgrHnM2JbFG+dLq6uOdt1Xb2Iz84OyUzDomto4yTLN7vOs+/SArXtmaTR
QNpSJnjkBEDfGumOIDEF8JFy/3p68OJwheSKjV2zR7xQsD4Ac+QppjYHUa5t
w8k0FJqqHayicHS/qh8sz/KkeQ0IJjpS8XIUXsk526ixGKL+RWyUify1UTNA
yGFdUn63JXusmPOjUQLIjVWVPaUOf15A1gsdAOdkfg3zys7Pj41xBR7bbwTo
z5Cg0HyGWRBozikupy6aytk2KZwKB1FHgLle+QbZLY9geL5ZqnlU/+Cxe6uq
3ehCO5D++DOv4IN2fvJ2vuOi6EPHp95i75E0WnnQsXCIuxV9TZXSiMaABUYH
GAodlH56JtAllEOMbx+jlA/7K5YUQAePx+p49LfQk6Gwc9qIyxCt1BdnaHV4
w1UZJVRj9Og42YmfOQitZQfttct9JnWnkXj8TEpwG9zp6NFx0paN60insZqu
VuBOHSZXye/1wLlFPKsUR8TAg29lhjUepW69mxGN2zDrluKOBq3OqiZqeXS0
NFW5sXkfHaOfXfeQ1eQf2k+hZm747g5KFASHJmZZEYHHIgICh7oPRM5GZWHP
bbGPgEhCTjkRYCt/5APWG4F0TCik8k1siDex7vlVKOodH6d8PsszYLSv0Ghl
8AxnDdj/qnRNR2HZPY2ghx42r+mbmq0VMtvZ0Di1QfveK5BPGHmwCmwtuITK
RTPPQ9Kb20oFsAjB5P4sZETxaSnYK+spfDguUFRe5QKGAvANSokoBDqWPc2p
paF6ha1l/w8gaF8sEsbtJXXibohY/K5ip3YbYQ0+ZEi1uTKD7vdaLibBuWYU
w53pDgio8FZ+NJJCkvV+bohbtLGGWZllxDat5KQDCRP/K2uWCPx+NMpy9akV
ZJiUz2lENsWMFLspE4YtxM7FCvliasN8266u5uoXDkLisotfRJ07F6PYxjiP
6XRPydyp8TpsVnWZq6HCSq5+1wAKOpelJmgijhXKmcz6PWTOL2o4d4z8IyAS
6MKETQNmboEKlDFTdMOxESb5A/v+vntFqRqm5pF7a7AEiwi8pS5PT+fMHlH9
8LL2Qz3FWtD6b0AyAtp5ayKAm4whcAMJHSI743qaCKj+t5RYJu5PL1cstCbO
Ka3ODd/ScXIvbWV8rKDfN8rFiGjXsqs6aLx4eEshbf2hrWRPVcDLqHTYOE/m
qOdKo/JyyBYUZKP8jVvpQOCartUCBFGWkJvG+pJVzWzPhHjKTH81L1N7gbK/
IWbQ2EJc+R4Xm9WYu7euxeOMxtKJNmHliUbqLiBcXfdEbQiyj0uY02locZyx
UDrOG5hzK5xfA204YgvqGp9+I99gOI9uQzsDwSRVNakCvx2c3U43xnqJt8Mx
6oo1NE22EpYzI7ZFp2HrGt4hZyNSu3mU3LMfsaHTuY5jMrEkkakhtY6UlkAD
B4HFN1WaKfge4dlMupBZtE1HjK4HssBoxEjLto0ESKkrJH8RXK64g6OqxMXV
TEOIKmXV7BtFhHxyrfKOWyeiK/pwpGv6SqMDzhWPLHxZRNdodlryHPhuNuAd
I9oar9wekpD9rUgWWVsyl/mX8Ai+Hw3CPENCviV3m0iHGvBo3OkM3Jdy8esw
k0u06dJDN4DYjfenwQ0w5at9tU0MwtTALBZ7Yap9claJ8H+HZTuM4aFgdfXv
2rHJBn2fUws//aH/kfU/2UEMSatzEdlCIHVAlNUYfpvKfT9vf5GcgugEm7Sg
1smYdecFrmGZm+mSVBlQxBHIcYQKzau/fOZU9I9Th8dEAzroYj4wQ413QoyZ
qB7UR9oeBRVYOD1LEGsK/hLSxR7XT4jgdyyZBfQC5YiNqTMQkHoaLku6jEc4
LFpDEfax+drDkAplDCIQXbtl/4AC+iBUpO5Z5HG608zCWmMHukX/u699r2Xy
YYyoF9pOdzL0IMY+W7WvJR7OE0irViQ74KZ/Umeo9ljZE2/Er2lIRov8d7JA
UXPG2WCkeKyhlfp2yxVhalqFyzxb/12w509uryS8F7zJ+wkjHjW5KGbfsUfR
BzS2urxfzyTRrqScp2EMTGC67TchAEIsFu+t+m28GIyZtFIdbpv89DzbIibs
asu+AT24mjeah6ek/fi6rw5xLqcFlj1Q9VcSwGUYy8K/YQ1S29KjJu8mpe7j
Rq6cc3qM33JAFHl0CWIk3mMPF6FTI/zZ1brKnMh/sDlYO85UwRlUyezQMJx5
kME/HAJs6NkvS+dgw7b25DF1nVwdDOuhXuPVzvrEJjd8alQrx+e8L6+18Nqz
BL3kT6pezwlMEe+g/KmyJkYqV2BGBzqL2SVqLQuUneziT0OJnUtNGWtOYSL7
dPW9mBBjSZWY93Sf0nux+HmBqkQNRqWoqfOhABc1dYHuN+3cRlW6xlw6lQBg
mER+OHrKc4hreSvX9Ph47cRpN8eLAUqIzzr0i1sfmNTQTtloM3LWkq/5W+bU
GhtQMcf2FIYg8kaAiAACPh0P2YnX98R0ZRxcPohDe2gQ5fN6E+E9+FCGH+ZI
T2FI17EuHGaCINBT2Wix5rVfJreE6nlU86QOB3ze3wXroKJHaYOThEve0z4c
aIfVTiD5H4HOvvH7hNMANklfLRIS09D575WfNTJ5MGeQiF1kordGUnZtWi8Z
SielQ7V4AguqRh7Rt3NMVrc/d+JPfPuhhGLKx56T7+4e9/Jp2hiGBx0k8K8P
fN5hSVB16fSPogiRRcPiRirzK8OcH4cjZdha8I5N0yIsrP1/ntKSZ4OAcKfx
VktK76fkdrAwRCSzTzjSBC2lVHw+6KKFhOvIpY1oz/PIILa5Miw1gbkAlhEA
i/pdoGVruxZDacC2psFDiczhMkVPnmHESEq9gPPRSCFSyD9BencgHKprMpKY
xG+qmyqxtdt1jM4IDSDB4e9XJ/sl0YT5bxOd1xIbA6knaE8nKSJDUZ1VXgnv
3GvhVTralCkiQdh6rqvlcvvwSVJgQ5i1Kv8UK8O3QJ9LmBq54LQs3VYE0Zr+
uOciVabfUJbaOJwhv8A6iu7XKZUp/ZCVBLBj74zWuTt9obHNDwTNOyrvIKle
Njb1D/0zeTo90/1NP/iScFscSzQHfphkoANRFOda9DB0iZ+sDucAITFxIg19
YH2iCqHOlxuEqX2gZxs2foBg/aFsIgUdDADOk2+tUzrzeJnWVHdnGnj7UdqO
n6JIYhHC7DXzx4ptHPD1uROYZ0FhhR0Vy4b6h/F8n7zgeE9O5iPF1gRCwSrG
acfW/meH3MSylnuVClXtfvgWn6IQPziJKbkqCMcErR+s2O2QbM3x4Cd0y/L1
fdv+AYgTveuy1Dma964V/P00SeJXDPueuPWkip3RuVyeQpoJz3v5Ysbt0AgH
HG/IGVLFy0C9OsgWDeo6QU+dPaj8+kl7v6//NaagzZEwKOF9oJGskpipfv9l
/E9hy5ANLbTAlx9vOKuDdXTqKPFmzq+7JNldzqw5TZm+zGpyZ6Kc/wUm2i8E
rF3U/q7PNvBUpznsPTLs+9RyFZ+DgmPBURY6vuQALsnmFUwaedAKDdGwa+W6
a53KNtnIrIRRipnd231tRwYR1tetLxwBmEWT3Lmhte4HststtFcqt9RqlRXl
UJsDeQzl8kIGXK6XrcoOs6GbFzPCcKGMEgGj9Kxg7gBW0CZKtXpnA7iovFnG
sQoXw0WHAKdgxA4twUHktKMxmMaCJZGl+xn46FUdZ8AF6B1PorKu0tzkrMxK
71OtGoWdUJan11h0NQ29K4VI3RYOpJGnZUjXBfRr+5bKJB3uBQlJ5LUtUVcl
psvMoGcNmXoMeP9/Po6Rkv98cywOW+s2fZEjZ/OfhXhHkEPSts2VWbwkyyr8
STTwCQCs9/ldiJB+9Ru11Y9e9KR/iQl9ohFUc8JpsG6klvfPaanj+XwNmDLj
uBhNlXthCUmrczcCJoQUlc259fQ/QBgAJjJvjRdg9kpKquR3qQl/RMvItrqi
gpRihH57TF+R9aIXVO+gIr5k310iCIXiwhvYzBv8o24dI8iNXnT4v/lZMxAi
7CBrbIkHptDRrDvjGIDfmbBOp5H7w96YyMomvcelANI/B6MKteUyzP8Q3SgW
zORDvH1bDKeJQQ6aTnkgS+yP1dIWN0uKPyIpOIIFpF4rTLs7ekqqw3VYJA09
vj4QyuLac91yiiO55CHD/5rOexI8tLxEJPcsWGYibTwc80RCuiDlHrhWT59N
LMFC8EHGxjHhJHruE5rJ0bIb9n1Sl3BAjUnocP24XLpY0dqFCt3J+quomOMB
Sy1lTJHIwkWOeYSDsCmTiTmMP+0fq9BnjzOSkBWLqI0BZ4ZPWbazxCHBA9qq
qveszlo2+N1ySVPHygvH6EDA5kB75O4bD8EMdFJiKWL8w9KGyDbB1NhohFX1
4dU3tfrvvde/QhCBDUJ1uYVTTKweK+yCCmchVTCRLuL5cFdo7amF+LNO5Ap1
YBonNlj33uDb0ASyaDH70N8tjKTGZ911nv39solkTjpcpgT1E3ufqkTtCrVf
S8LdcR9xWNPAghGmjTJ8ISyWQYHorp3x3iCOOvDsbAK1ouqmYEbukXtVA0tN
0Gy0iIWzLuDc7Mo/3QnVtPsHmptnPNQBPa0Cr/tQycScrpqe1cosAJCWgmZK
Wsaljh2qj9UaKjX8RXb8/W4AMLlaCeBvLJZnGnmi+aW1Y9LobKYs44ZzK4q6
annlrPpCbEnxjeaOaeeqmpmaDuVu03b+Y7sGiRJKmjMwmPLKz51JDVOZfZG0
uecRdVleubA9pv0t+bGXL0slSUAfr56027qEjA4EN5QJr+txghjIC33+GTDS
td9edHp/vbwXhSn+AHiJsTA9tVOxfQ6GhdPal3Gmr2lzldosufoaGF0a1ki5
Iqez2LvDHioadZOCU7Zsw2gCCGQYCSz0cCO6fhIT1drlepHCRt8tWYjuQHyl
R6AefqT9JsG/2WAl9im3dNeoTp+UjqCjX2MYvDp+LZH1l56yfeNHgnN40xQ0
9lfNYuZKrx9Rtm4q6iTseKZu4kHVaZ2bUa2Ns9xv4icEKMK7++JMJ8vcMQta
1mD22lzBPsi9qiYiiABrtBkUeESrjD7y1jAUdAjLU9W4YvdWIcDZXm4fxblb
UFTZCuQW74ZHjWzErW1aSALVtnEFV3RUd7s0ClGUjQgHukLP6gY8yjvghiJW
mjyKfgZRH2fCDklVTJzs/KPY0DlXNyDLwJBSu4Fkowg1TElTPggZrIuti/o7
ZNfF9dSq3WR5ep22hk07zH2HaWafC997g1U3WdR4VmXakeZyhQBttHFSipGZ
yghbP+TiUrDvlayBRtNKElrEbDfRLcQGDKYeDendYzwTOW3SfB5DKOS6GmfY
A9vd9JtEJsfGekTgR+Od8nSIjsFo5+36DmatxPmCu2eh0OeamMHRJrCdKwLb
fY84wT/G/PRMOEr6VrpfyTK34P2cJjyrslSmrRputV7Uu/LP+I+/cRg/Cwps
8eWMK14LPEcHGC3lRgYqlTBuPPawHyZSwVqpu5796OxiA8YkMy1Au8GUxPVk
Iz5peXFQp5vTokEi0ckwUUA3ijmaycCSW535r09084W5ghJYvTRjz+6Cib1V
jfRtJEm98PxtlqEF+GjMxaFj3W8ugVarh3owFcEPjv6ES3/D/Cis5zBBEDnG
Ce5VCQ4rwsVEnM31bbE4/KQJ2ngesAuYp+ywuJIVmhQQbRZsPhXE0wH1Wu/Q
zcgaL13v/5Bn8Xb6/YBynLCoab3Utiwlg7hWyVxglOakbHNgbJBk+BSMgfsn
FXko6RzXidypY1Fu3pJvwvQfyMbfXuZKTI4osUyWOKkXocEFihpNVmCzk2m8
FXpgWxKCyOrYDtn51FP3aFb/cYKmDhTAAajGc9OooN3CNUQIjKevbZRYfTFb
BBiyJoZ4/Lunf/wcI4epwNOG6pFxtYPmzSagpnAlQ6JLfatbkxuU/4KrpLN9
U55R4Ftcg/EZByRYmJr9ltBOwIMfOFkFk2d57kRgBGnH37Hpah354FbBZovd
n91zL6D0zLC7UyaMHDfnw8+0ObTzL3MH2n3jHadvBUPUcyrpY1dJDhGAWcSK
BIyMQiGnhsh0/tnHlx7KkYHAoo5BQ31BCMBtrWhg2U5n2n9I5Rek4NGhO8Vm
BtnOl339uGs/xM7a82C5JkhtlXXNozN4NjRLZ4U3hhufaTgKYS5xOdFVt1HV
GWkShekFfLOaaNSeVZ+/+OXYNv6MDwCiStuvnDAT5hnr+OLc/pvkG5ijn2Pt
y8sULklLNBCjYkOsp+TDifH5o3yoBHoNWFk9BKF/KyaeaI08InASLOic3YX7
rV1a+tiVmhL7DpT5Lsfv/lMNr/7WkRfRlPxrdb82iLXaSwIt19uYKgCN4lDA
JVJTtXyBOrW1Xh0OZuMJ7G0pZOvsKZB7GM5RYk3Zb8tfqobJbjSiOuEp3Rf/
jPstrxYgXR3egXHRGJcgADAGMAN9YrXR+9BHI7tHRLKRiILU1q1Q8Ct91QOa
/zFGGB9tFDhZLEi9E/2m/oj9CgtZyDmVescxsqanECEUegXN0FxPMyWFfAqa
4LqYWOUDxlJ/uDJVkw9/YJDAICloZE85y+G+D07sTmcYrrLDFq6lb1wPBpl3
L4ThiUf+1UKBqt1i0V/uuCFWiNfgIFoaEzlfT9RPmlLjDRiMdBfROiovL5q6
UZkGmWoMUgYFKkUQApSvFsbRhGx/APxUKS3EXuAV5Zl+QAeU9FbIM0pk76yG
zw2gWoctZNhH19hHO7BWmwY9GyIy+KDx3k800Hzx4emVt+GGntVn2eYF0oEl
r7+6E5lii33m6cmMt+Jzo3Z2gCX5iQuji/ANezklLXuI4BPICq1Do/3eS4I1
YAsRPvQdSEmKi+BRdn813w7qfR2g5kEKOpb18usTSAxLnMdUPoZN+30QktZO
uSnvmuPA9qYFpjzRSkYuGatc07goCNkZkn5NZL4jKiwXE0M6+WR7KLPp6aZB
FhBiDA7bdz7TkND+66HSv6ZgwiyA+j4UaYZUhZcZPOBcoyesqUNWlkMrG9Mj
iAwdwCnGLGHpQJmCoyZoekA64Bw/7oi0g0fICJRQNrmUAEB/0C+qfsoHoTKG
iQQxtujHR76aA3WsUdQ46mLcLLiS1bFO+JyQeHcXMMdYzIuYRwARqnOEbd5h
E9JJuGlc5lcixn8SkLTL0/gvLL5Ca2aD4api/DUFNsNWmHz86WdEiTOs4lhH
P6k9IzeHzQalPDyqbZ/ogbJXkXWpsvulRW1/eEfA76Ot7OaHOf+BM0VeJZRh
fz9uthRdwpt7D7fD+Ds5527Vp0AaLGQsCWEQO2xOzuOxt0z69sL8atYE+CEn
7yC08AHgfl7JbC3kYWleKXcX/l4LKpX3z2XQ94lD6J6r7um4pE87kgfxtj1Y
GcPsro+9LyF87qTVr9agAwptRa6R7ct4yLN6xGDCHuvi2jZ4Am27mMT3vD4f
K5y/tfs71LIOB0TEy+q+Sr7uRsWMfG0RIqPx3kHKHXRNw2vqZGyZkMiNUOuL
pm67K9tadJTI9Xj/ooeU1w8SbLAP/oToP8YmO3Fho75U+yoDSVpWADj2IlPT
0VIe9hWKE50KDrZCzC7BVIIl8hd4FP98G9i0HcY8Gw/dc5IQS0RB9vuKQqEZ
5rEFtWVfAjQH4tYPZ+r14sipVVODhyFbLN/tLglwNmp/s4yQDJ7CDkccLXHS
FRFgdpfgy5sOy8oGPXybtZOzjSRJHJiPeOUcRptFTWdnSq5maBfGJtpJhPs4
BgzIcV1Wn6At4GzgsSl1g4NEuOq643t0qVLgVfqNkx6x1kQcwKEiOE0h0Gqq
mHcUK6ZBwRExrbKKVnZIP/nTTIWi6M75Zuhn1D7TxTS+f8kdg2a9PFpbKM1r
t73OwmL3x6tglAlu9ZplPK9I5T3tYRebiJ/JNqDMO+mG/11c/TdGpfvGkb0F
LeAlwbs1UBLdEoFMHvcaUQBJe169CWU3Hj8fV5OTdAtIlE9B1W6fevS3Ihpz
8llSeAhJVqVyZ7HQ1iLulrHSRAoPXua+WiPn0EsILsl1pr06TLv3n2RNBPJa
Zf3pDOudi7xUGqHsYO3EBjT1lz0xxVZfIIAYeu15FbcfEgSUyvFQVSYhtACv
ypLzYV0JKMvhCgpliTf+f2YiE8f/3r/kmi4mdSUfmJ8sWdcGbXQyWZuh3UMG
x+p6Nk9HJn5eg/03YRt9n3ED9j3kX2bZAvG95p/6OdqebpwxDm2BUZNeyqmt
lkAGnfpu1nMzBJJEy4ebeOffG1oD9aYqet7g0QJj6eWMsrlZ0CcBuQWjbj9E
hBUGd3rwWBbY7iN+jmlYML/SO62O8833JVwCeQEIgQH4WRVHnbfUbCA5ZYLo
Ttqh8uI7neZwqzy51rlPkkCQiUtnWGFpTsHxsMbqCbuLYvVwiN+/hGWp84ag
MUjonOMRtJcz7nwhda01U6vCDR0NOrowy2Bu1U0LQplXwq9jAd9Ak2ajRAln
p/jsmGa2mpUnM7ryooeNtQ+JXeJAwv8QWAWuhhfsztiiNNmWB6UBd0sfXv0B
R1dztabbFIABGM9H3+nwkjk7YsEBTnjG5JugQf5UJzE7UGvP6dHThBVrAtm6
jEREKEr8dZvL5P6wqazpuvHY7UPuWf/7AP13MxL5uvi2JpzOugcSLcayuaEk
eogmAVyjxVlUWy230jVFkNSJ+zn5E0MS2zrcD2cXb2BA2h7QdIB6rZGVx0CM
L/so8Q906jiGt0V0LTe+0bLgxCzVyA0Fdnk1qcqK0izvp8At+jk5lGvJCDPM
0J77FFl44m0o/p6SsnUKkohUU843TiF8PhNN2h703rKxkMxo05awqW1OU3tE
3pd/6Fri4nnfBXdMuOiX6uWcnLRLYVWkXINIFIaIST8TJcH30A7zjSJZYN7I
+9qTblqPyVz9iaq/9ILrEUY74VEzChNLZBrec2l5rIxVq1UrduIMv09C8cYK
hev5BiAX1VFIR2HY2ID8NJgHxzs46RRWAncoqUjGR5q0hOc2agdInksfPMxp
0eyEs08rzmGgyRGcPOf9TZvtzP1zCumt4mZl9dfAsTHsVvK/2EIba16sviL0
97c2UKZx9N/AZLMGHEcfOmphxlEd17gVvM1MpR+J5XwQ81SBiWjiltlPRypY
wY4WvqNNtsjODjED1rexf0zIYT3eBnlGG3HPM+CwUf+nbXGvr/zrdVnQL6W8
/KdV4HI6bYkjNWc233NLNE8HDNmUvi4o5xpGJj3SAnE6LdImfgVYPhndNqcr
IDyumMCkgwRzTrXfUY3itYSMo5qA8ND5ZZJRCTFK4/2CUjuhMxW5khIc4vv4
D81y1s/yr6vrokr10sI3MNztLpQ1tlWyTIMXGKaStvnMCNP4IBUfAvamTBlA
8mlPoIfrKqPnzaNH1sBipBREedQ3qyTGf/H2CALrSDy+nB90qfZDIYz3QlMA
/QqpYiIdQQM9ReGGmg9DOAQulpn9uMtIg7JvDOy+HsbzGM8I8+IwpHyDF3LO
OpeJdcneZ1Yj7U1lbBIe4wqItDvjVod4/I4BpRDon6CWAJjYtXiNOjexkaf3
ABZFixtXdnmTER0KlLcwcE0NrM+a7jwwskH+xJYU80N9PQO57Cf8/f54c92U
q1ewXnVEU37lxiP6QcbCyXhe4bMCNKKUDSmjhWNHr1SdCxgOuxWOG8SoEJ+X
dqO8dEIXsd/1W59RRtfCbrjwT1KQVKvo4HW2U9oKZehNhghpAcILpDRc/4Ft
MBlr0kdz8ZxdX10/UlhDiVN23Q9o5XzNfajfZAEZjmFZGVSaPM3dtWkUiSNH
aM4940wqgwPzX+kWBr2yERtMCpYv+FtIfxKrMnMnpWTSTYByifSTYgYAgjO5
J9m6jIFJbv46eA16Qylv/S/RwGlVcIxXRtnPoquakWRX7xfAYpEOoq5u7hkh
p+7RTO+Kmc1dHU0IDhQMgsQuEhEnH8+F6/uK6vDEiAwDkQPCTqg7f71iEz7p
DcTePfRh/2cQz7PMpf18keELiOHDL057FG3LL/chQ4cepio7XtA7sLQkN9Kc
9NyoZQPvmPGchxZQKJcUF7d2SN66T5rfic/QsO6DZFAzuFeelRWJSIliEDR9
vysLljqwuytIhXdvWxOJOVCsTzibQbprAlGWr0hIrEH2kR6lghcLxz+UUpnK
wdexGCf3exjo0Z4HORSJKURMaA4dcOZ+2+5kN84rCmHSdOFrPM/HA0XNMrzD
DMtmbTThPtyAsCe7ojuRE3MJ6K/rTD8HRqtG0b+mUeF5Mc6zUuJpLd3Esnis
k7YXE4h90I87GC6tXEtS1Lt+e1k+I3WyZEFgst1H2d6qU2u7DPtrc2F0p4Zq
bsDSFYRtLHA/UnTQAX+KWUO3Jt9Qk9LF5JDiEkZCUhVUmxVe/6AglFSsSEU3
zj0rRFql9WweKSG2+kKMnkxSvD/Zeekz88yp7WBaLSGEz2qsByxextERt9SR
et/oM3Byzr4l9/KNlfmE2kslRBYTrVZLrPuRdXUBgqk5wRRuPYce9ZplLY8/
kRlRHoPtX3Iv03Qy+cYAKxRnf/rXIUmTDedQEnm2r36XAeIzrNzlXjysFroJ
rbj5YoNXhlJsGi+QCwJpgPxAmTPTAG9om12HrCfJ9qGb8FrdSELkydSZPKTS
9ekB/P5Z8+6/+8j4zr2GSYVFdtqzJnzP5diKUiMi/YUJps4jIhFdPTR8KKPq
35+HObFXxQ4QiWz/CJvJMcTGz5/EccUIsXuZPUdU9K3N82IRo8MTo4VFcQEZ
p0V8hCLzakQuTS1Q/tkkL0exzSXqdE+0GOfTTzgLB1OMoJQdqhWqIkGX4NXH
dLOkqTOew6La/FhnEhd/gCwT/DLP55gF/teZSc9YU6CqtODOhebx3AUuEorE
XKbjvuQkIXeipcikj42A3adYcO7Xelnwhp23Cv0kFQmAFpTqAUGFy5Dlq9/C
KuRRjz+5MJXDD0t6uclkyihacvEWjTvoIQcLp29YAZC3QvdyVGWZgP419fFC
C8G+5/YPeDD/1h6vzzJPiC5kUH+C6Asla6dv/DJ3gt1FBmqRlOTQ2X7u7+UE
4AkrogOOQGIxFNTIMLTmCA8qhRbqphS7L0VlhivqfgPup588b46Rq/HWxpJk
JMZPFIJlzrOfwTmf+UtywnW/s5f6Y9fFHhvAHUoD2GpPsny1N1oGaA+OmJbV
InnxZTQyxKMvCvoHzsJxmfoTdLfP0tkO5NDKRftE3hHdggRwvkf+PWqle2iD
ZJuqTdZyWHE/L2bvdNJMdhtvy1HJ31+7LYD63W1LuIKWyyLAmZnOtbI2igpF
QsbggYtHWUdP2Pb53E2ocAyKeBwnfIC4FvTKrc9MBPcx/I4VF3wlvVmT8LFh
xbH61cPrt9UEOR/mNO0WrL6YJ4ACvfE+k+NnaE06Gauk2gEDuBHYUPNWYc/I
ICbHCVplhRtFteHyTmlf1xq8Nf9nHZqd9M/zxS4xJxsbigWZb4KN3MEenIVy
14Fnhfd1Lz3BKvompzelql9ke83NFNtaTGdIwImmJ7jYEfhn4dCJzsZqoDLn
QWJ0jHk2yor2Y37lEA3Esg1ob4mtoHXoCXNxbI8/90paydt98ySndiExEIkA
xprchnINObk/keXN3FZERrxiqcOvDnXx8BRL+a3trEKcSEr1mmlpxFrVN6VN
VPnqpnwZnrk1b7ZGQSzMCSDexpMGgvgcCXvX+l03cSMgeGTPYO1pL7U8LUeq
kUaitPER1dejzEWh4pGOaHNX0+OCOUAvo6ttVpbK3drOl4da2PlsTIsrFmBm
HYXPTHZPIp+CmPjXwP5Hw3LM5j4e+qi0D65s1zBfGvfnb/XsW+F0H5dVC528
pv1+/gqL7Ek1owfbxZJXS2tiY7EVUzZMcFEftqxYLmCV3lnbJ1eREikmXseN
nhNZtXrP2aCBW9Ox8vW81LUhaw34o/PbOg2c74ji5xWSiGJlmvFJM9eIsPkj
6ySkZ3Qba+xmwn9JaYM9KeFEOL0GBxHP9UfGAUqXVAxKXbSqgl2TNsYCd5as
2Y2I56xgEquIxk9s5MeYRoacroiiWE9b7CCWmWf3cDEhqbzzE9gM8moYcnin
mZf/S3is9guE6UxU038ABdG4XMuUaeTOTQ7geCLCa36WdZxItrZ+8TLRFBs5
iEwxpsIcvFtIvrEeL/o5ikGQMTkPfIKdJKpXZrf7mh3Xlsys1pXVRg9V7pnn
d+Y7/8XtMPNRuCDb4DYk3BpKIS82HIfF78jRc64Twt8vRnL4dwRJiHklxAI2
t5WD05EzyjbvsrIIZT0UHKtb8WX2JOyM0yfckBPtMq7WVvfEdgf6ci9DaZZ5
/D5uC+KIW60ReLFwEygvbhkFmkN2V73FBZkhzuChO6rM/zFkG7iTQOsgdhye
XqABtiC64ng1VQUK6BsrbuONJTTmMtnD/3GUKTO4O0a1lgkpaAM39kWZLxFH
uH2rw0w+egab+qN429UeN7JhqlNts/nhhUmIiTLkGfrg1paln4hIn3TbO86B
XB9NhVux/s4V4t/ov1RzZKg8ACscmC6mMEhuczlUVBdG+TUeCj0nVoXkOFoR
J85RYaQuAC4Y4CRfZBOex/o9fk43fHOB6xojeIIL03M6WCS5sikFvdT2dWzq
gbzcH58GSwvDy/RIBTx3dBp/bD7Og9TC5r7fN81/kos5TBqqJ7vmpSic+DzH
H6XevUGYbOxWzLHxoOG64EIxjv6wOruFDPZxporSAEjFMzhgWSTi4YghgLhg
uDS7UdpMkzDq+xxZ5QjNHzvZN7J9eJBr2gRnazWXy/AbyfspBNq4awgEDq7z
qayGQr1ry6KMJ38eI1xM9Dva5NvTi9n7Pqu3bMm2NrS4tFoCb8YWOIA9/BIK
ZT+syNzgQjSo+UQrmlZM/JPFKcoEDeQHCWZ27pMOeQyb0L55ZzBb9F9MIiho
1FDjp2l93SEofj3MGKmCYGd9OPzO5rRrYtkdOCruLiC+Bv0P+l40KG5d+wcX
PG3H5+PQD7Ca9jgS/cbnoWBuwBXfvWy34ASAoIdEma6TEyqlKhoN39MwROL4
Abl1UHk5k+1CXMDgwZmzOdpThH0dPlX89Kb5eDjr4W87WACllSONnl1+aMeF
rRke1fUMK1eX0SAjQQm9HS+zNY3OS7WV2+lCg/oZ3vA8N8NLQuCx1nemOQH7
sHj58Pqv0Q23sJKgD33g94Xm8TwSMF9XqFFQqfuBFSUGsKSmc4h7VKkRR/qt
5pbgDXG838/HYA0sH9lJJpgd4JwqFmuuAnygK/fJB2aj4qTKR3jzDKmNcjE3
TxvP7ZCyZW4BPWg+q+jIBtvCj0CDAEZn+CXSJg6EuHQcl6wNfhIuHcWZEs6H
hHrea8NXn+kAgEgGbPLblEPbQ3vDDPfwjqqhhSpyLaHJHjZuqUPrY4DZrN+F
bZAIqjlBGZJKh8IwrXQYFmLifANiA4fS0llMdiEqFA9kVPV8/1O/VEl6Rot8
717PahylV0OmvX5QfkLoUJtVc2Rv9DY3ly5eg7dJnH+bG2nH6Y8gVFxgwVz1
JsIgnZN7VfAY33tHMynqQHFfTSJXWfQHMAHsyBtkRQEmbzPvE9rWrTg4rltk
QQeYIfRTCFxSJwQ0cJSeRNX2up7aQElo5XgIMTrfDHvwNDeTcsr4OL0S2pSX
OBAShM0q05YOMTOFoTv91aznN7fNcXpy3UDanZhBAyng9gVWPAE91xwBkc43
wiiHVn/8K/APg9AhSq93OM7fcZKSVB0dBs8/2AJH7TidKsRAnu/gD6JhJ6eH
F10x97KT9EmY0GSztjexqpR+JDJzs/MYJDOq5rkMx2GkI12dpinSruzyz257
oUiqE3a0Yz9JFyNYZwmwbHm/1Isln9d4wX0Mt14we5z5voJGy91ZtTPScZd4
mJpCHieeb+28AhVbG4CupAyqPk0JMH8fBt0qngPrC9rfgLmmVI2FOU8RVc7O
+08z+sMzOBxmdwPZoi4YekSoR2p1Z05A/zomL9Eoh+N6z+1nme0mA2caRpL7
tuOzceEYYDSzb7KoSloos1YJMnUTYcuTtVa7xYhzuh0xNHvJSsxyFMa9IF3A
5sYjttpanAgivV5pdC6fo+luBtM78RhAb7Ve+bXZoTNjNKYOlPny4AXk/zlr
fWnwYOweEEqJiC67RorlOwgqolZ9TiAENK13SPkQSh1jPdiXW6Z0mW5AWZ/F
FTpBOLDHcXKuRDUwsYEtiSZrZaa2d4Qh1QC+yKvl9nv6Gs7m0BcrHgaA5xWg
fZmZqir0PIHRUY4LM9KtmvP77JVaE1hVUx/TLKDRxx4L1HzWbs4AyhP4DGn1
Z+tI8ZPz31MSRI42P7BbAottC3a+x8lwOJN8QKs1RBDtNzpwl7TK9oex2bvg
yTYlSLKaCPAOznSMx81ajhzHkt7dDsIYIx+f+aeiCkoxbmW4LoEDcxccjCKF
yb7K9YzvFYAp5dkI7Yp40CSaIO12uoOUXxetR4y3OF8SHSWaoRcEQ6c4N4n8
iIH81o/6dBDiwEA6F7guIBY9RWcBKqjl43nNxzbuBSdFfSoI2qAb/dHg6btg
gJJ4fTooMQutNI1Lbotp+B8Z9fRVn7JivzwcUUV1ZIgJvHxTtlm/rUhwSpOH
rusnVP5hhkEQBByk76bmoJyHzYQhv1Z/1n5mhI1dSIXjFbax+66bGTVbm/yT
Q1ApOpek4UB2m3V7LQQrSbL1sUMCLZsrjA4fXeBcorGflBN788/ps59P20Kt
Jxn3NgDZVR0a0oASAu7WHemD9RwbzLpJ1jsIPA8JHqVxUjYZQX82WUX3zVIM
ZbTpZNOMRQW3uNuXz9oMBZPffAVIovay4GUcUNK4TCUd3ru/xiFARjcnqxOV
+UseEIt8SGnppvj72CN1u2/VjJH3JGpNrD8VKZUuA0Gab80di7tiLmuBtJy2
8DntYv/PL74d4r6vSi8LHJQlTuW098OvyZhnDFmO27VYYzb++XnW3II/zjUj
aifuKrC9i9+CRNhwDmb2GIRxpEiRZcSC61LyjeYRzFGSaS4fDgZO8aoVrqNu
tXoaeaUs0IL0uFVMZDS8uSF7B0JtdEM1384wYwaeYsoMsby+PM4rSqz89i/d
RiYdfyj8RqRyWWXlEfjp7NcUMgUeybfeqDtg6NrZcIClkPx3vHvewOT/dAwi
ex8nKAGPG3EDQPv78nqSZf3YQ8UNZdWZGKMbrpKzQf4NOA76dYW/vTj9Tccp
ocARFnMuXByrgBx9L3eOahPcbjYDE5PB7XmKfSev6VNALVWzBuqcQ1e0Ej+6
u8BUyfVbyksiSIF4ayIYUsFMZIU7N5/oQZ0vUXp0/atmlds4W++B+k3auERe
Fehl7BDuVeUt3DGPL4Niar21T0F9QGYzUGiADc4uxb1RW6DqxiK/V04F4DSZ
152eoEbkS7KtMYUfcuLAMU0p4ireFyCWuOfJQTrKT0joKpBDjyAWScl1VUTu
6GmRW772nzZqAajWcrF2+kRK1eBlII1tFMpMYwbvua9v01M4Zi63CevDfsF8
0iFxOk5JldJIAB1Lkbtn1IugPSWTHLXKl6jZML9/sY1j72G55i1rXTRLNoFH
ORXQzvA8k2qPoPTuiBopVW7j21qVptyR811QQ/bjSz63M6uIO83uNgL35qaP
LuHF7CvZpk13nuniUI3kfglQukGHFF9kKITCgOUzpGarFG0cOVdyhJiqkSx+
u8KchCwQxrOczIjMiGvoo21OtM9VK/NTKuBvb8x1ApfUZO7CqW12qydzpHHF
MpI7aDswjoNlFf3cjw0VZXz4zOaG1UHDwDQMBWlaka77MWIXZSptDhncwVW1
SlFZWT5ICAXxeD/wdBN/V2ltSpbL+LkP+QrS9CLWKSNselsSXvnBGaSYHc2T
aR/FR5pW/Is6npM+B6s6TnTCXi2k/FZ65DjJRYKijHR3H4GfL1arHwa7CCBI
n+rLf6PGpio/4B5z67nrfFOoPXSg/s+9OXFnZkeq9EcWvfsz3RJVYjdmTU03
s/KvG3qWBWXu/O/5hg93629cf5OUeUJnwF3st6x1g3b7/0BpmZ3ofe2nET80
ee47ni043rRUyWr3folMqSl/SjgyVQbv6trCmGK3ODIGkOlvg5deZ0HxmmBf
93S3WoJvLZlKBe+jrBVG7XTfawWMTSN3tLqwC5kiVhCRSYO134q2YRiyqFKx
L9owBSzCaAI1pTvBJTiT/245b9S+20AU1P9uu1LjGjAr8EvxVnZxuvc5DhzB
k6nhg8hf8NZ0nBQ8aOHUaW1jUiGY5EEBhWNvop+vnLsH6rs0NggzlkA/fvLJ
ohOhlToSZya8qEpw5HU/4jcaWnxBIgUQfjdHbfcUvF8aer5bdZIq6p+JXPm2
GILa0SI6xCb4CM/cYiqUc42LvYW+tmiboF7BiJtp8A2xuJ/h/ygMyXsFJ+9G
Pb9pTg884fTW/bjsBs4ZeNdxMdcoc21uXxA1dstb5OURhMeciDRtTD+NE02Y
QZkuhYD1zHvWxCnhw2Vcvbw08DwahnSL4OaAoj+47gC56bp2dhPoh6gR7H/t
9LShpqsbsSKIkmvkoj0ZuJAm7RszPkiKupL4K1iASvgM944vif6aqjx91QW3
HJtzZnPTDntEpSigj3FSTO/MqXC7mWOqdXsPHw0xNNC74RlKxJ5x8rYgfgKk
JjupCfMMiGhuS2YjO/DaWqiUqEwZgOo1ouedyd9ghB57XOeXaJp0/ye6Uct9
Y+X+eK8rHlwWjtnlPWV/mmw9mzZLlQPw+Lynz+XeR42I+pex9uarJiD/fdeB
Q992qKYcpaxlKlrLVC6M3tdOuypzBrOYD3eT1SPQBt3SZADniwtsCWbbRrty
OpBMxPxP7SmRTRS+EdKXl7fc6ZLGSZQdg+l84XQ7gGL0DDioLEUr1/ujlsIp
75mc583x2dcxre9m7FHe0+gRZq3AMrJAhKSeAApxMY3KtklhTLzpdXTE4Wvt
eQmDIxzCdC0PkzOombIqkH8h2kS2vAb8B9tRiwDKXb877YjCz9mZjTsEDt0r
wo8LyV4+vienI/Vv9CfvYAExw2lBhe4Te0wMwaGWtIQjaxQmKIbHyhPNqskt
2KmlTXUMX9hYwwaGh07laO+Ra3Aie2p05ik2TCHUo7c0FuKvisVA1mO6V5VP
3O0njJD/ElmddbssCgg6g5c6dQFoPFZBEUretXzJyAZuazNfyyaWd/bdUA3s
1CudGyis07qxKzug0BYL20tYR/irX4mmBw43XVR9inuZeEtx6JzDEujo3ZE4
Glk+NEp8YNF5nL4ZAHCL5JVZ3HAa2/TL2GGYWjUtLp5Zkr7jTAzyTK6+eT1g
WmBoErn5lQNipxggbra7oW9uMlLDC7qUtSp+wePXjPEFKyvzVwohXlKCUO3v
F+UUu6mDoe56o4v3lxOTWhgGxCHv/4WfBCUFhQTJ4FJ4LbNv5wcxITNjxhZV
ha3s1ZauW9JN5j6Mx709XVpJRgykaLYuKC+nLI/aqwtC2DI4fBjUWFdoXqF/
00wfA/6IwaxEtArdUOAwCMDznKAd0G5waLIeDObgVXNT+Fax0TBlPK9KknT1
niiCUsF9WfIgtKyJ+XJvXw7FdCG4kzIIUwBGw+0x0/zopjXDO/SLNWMD+Ukv
wGM11yU2hFslWDi/rEKet6kVFEZAOn2uCD+tC8Lv0xlusntj2OzJgfDG8EVw
QBZuFDXwKi4EDT2lPF8Uyi1/CYcyuld7YeAdUOtZmdkY8XsFmiZSFxrRfd1+
ddptLlavHgAHnZXDx1m3h3D4Yw9ZtlXoCQsZ/k1F31HDKGXLiEzM2+ap9Qbx
yY1f8LCXQwW/kUIp5WLHVqfFvGVtGj7x2OHK3CJVp8xCdG8R0ksBiOD+wEPg
0psv4hg19W/Jjv3HOsO7Jo//zYiO6mn+7xv0RnpYzwg+2EvSoDpspBMMgS9a
edtXCLs5osJzGVdCaW28xl+k/KIsewc5MB7fXBkOxRIMPkU/UPe/a4UPu28U
/rGZvseXW0VJfuDc+cfc3CV/JPaGqGltseK3zPLF2iCDlzq6PAYq/a237xVc
cGYlwZmn5Hudd05g7qSkeHxhIUicU2O0mFJNRZbyKIe3+0axOrDhitirgvH8
ygyI8yFZRhL88Frz3vc0cOvAix9X30sE+V++IstSdQf27iKMmZqXyvkcMV/P
Y8HvDcxpxkHcSSzABkz/dGGM3oRU9oXLRapKTNeYBI1XpLIEg8gYFUesqfbO
L5SqYBE+hWozzdepmwLyVGlP+bf9MtBgh0JC0DGz7ClIg10xmj2Vx286n3g3
2wMWGiVP2s2cSx8M60wLHJMhH348DVGVMJkJ2unzpZ1gTwRi/X81liGa2c3d
K6uyEXIye5EJPrQPB3SzFhuyPXbKHH+lRFsbEGTUhtQe3KBfyOLrjDF16eQ3
TDjNUgBlvN44PuaG7S9egR9ovQYsh/a412Pv59aTMujrQPQ1aoxo20qktVrt
WEJMBx0D/ToqJskiFo0it8hUurbtQZfEbD+KgmByMPsb0PvWE66RUDHCarFM
niQCeDdl6SJ/x7KCxv10yL27fSI7rA4itu+MMtGlbrr8bbRLD1XBdC0QdS3z
jL+adsbZrTRJDJHbM/+Ut8wziJKiNizMr1wFxwLNXbobyvGEt6WjUdonSQek
W2wpJWN2xU6ScURqOcBgryxk3sWLM0p2xCwl7cmYcj7k6Gg7+QY9VRD3tUIa
oAmsB38HUyehuC12yLTo9W+2xqsRtlTXzij8C1RmzLDQrrzKAJ2RARxfI9PB
b9kW5onHNd7uYmTiuqU6L656KcPdhmnHb6nQyyVUdn1Ru5ZWfFuMJ68gD0L1
jjuXVZQuZVyF6rTCu7F9snud8tdcA/klLT7Bd2SBM1G5pw0GIpT5K3VqMnDE
7gL/7o1y5jvbMUeEXZzLMuN+uDHwoRsuE4tuHCytMo43G/NVYU9BnceS7Fa3
tHMcj+Im8XSaQf+02lK76nJxGqO0IN1LKsy9mzWcCYVo09UsYHI4O944i/MS
CTMUeT+19UV50LI+3/P7JgLQQai7nfUBN33X+8E7wdheUVQ50B1viEF519NW
7NKNSJag4YxRu2h4o4Ahpsm1Ndd8xDKTvWZ+ETRRwYCgJyc7byVJW9iL42fM
8qQp+tpkEupNa6M+nkyDMRh+N12HeLzLft8xxEItZ8fcY36KRDnTTHCtBgQB
ke8kT8IBQp1weViPvKdtqrx0KIA+Td1MylHgm9/XHM8qq91C6l1SPGogLhn+
YTCXW5cmtkvXeU5x5Lpqnz6pDnj/72TXX0zot95oF4JkpQurBigg5hNM/LFk
8MRzv0Rekmfl44KfNe3rF3BvR32Ms6ebYMTmV0ZP6CtNZgz+UfySoAKZcJ1P
r3VUvkRIAc1Y2d3c9CY9RzLobpk9O5mboStIwQuz6Gbf1yjKonBuZC28q8/H
Jfb/KRhCeiMA2DAfglBMGxK9kBEwC/l/rRcF5nRfw67YGVe8XuC8puFNUnTD
vYt8WHcikNdkPocsgig3CZBdO6DXXXZwiwaD6ZXJEQ6UppOvmUQ1BFLvovJd
3g9MTpm3IoOBGvrgL+O1ppCnO09hZQYWFC7sD/g9T/mnk70LYPSb9OGSoD8z
sPT66tgKonTCpAzz6AOXuMtW+B562AgfaNuz/OxWxLV1yqQJjB18RWAZWXDR
nwQpFUQon1OgY7pAwr4K+i1ISlwKHrjmSI871JQcxUlVfVMZRGg5Lu+FEcAY
vDbz5eRXxzl9+OF77/Bi67GDXVbXJoi0j8ClDwpuThlJGERnt+jDhKK6AOqn
Q68/NGmYwuGFYM4viLU91dwsgTRNqqBpxDngwT19IrYQpwy9eU9bbhkn8Zqd
J+A/t/KDya1jlyLDZY3DgdJH0ZgkzfIf1ngH1uJm70PTerNy0wqinn8l6Vz7
CRVA2Q37+qpdWvBFPS5uVuqoi0ONX4YDbsav5GUlshCgBNbuQoqolG/BeTCn
bFPSStNNMlf1UeA3jaPfHuYirHQuocE43a8Fl5PdThCi7afxynLwJqsX0doJ
BQCtI8wwA8GGaq+ByVfDdFnzPQHn8mFTX5Ce3UfdbphXqx4FSMGdA8v5jXAG
b7cMIwbr7CoEUag/EPaK/fw5RtEHqAk4G4KpIRy8WIxQB36bG1ieYJenbxjD
flg4i1PtwuvyIYXW2tCvZ9BS7f0grdk2FS2NIRWzUl21mT1TmHaywjq3hAB/
pgRWCGR3FT0GoU2JrVyAzcZg6Yrru7tsXIpK8OBhkTDRmAYyu8MgL9zbQVUd
+iwsr9awve6PVtZ+erePlK4zW1A4PlAwdQoulWO0t1kMa8XR/VDzhOPGyzOR
jiiXCQxxxBETa8Sx9m7QG+AurxsSFy/RP3yi0oomN1N3GsHcjMHjy+7tk504
sgUWjIsUe2Mb3Xm9SpCIwL23zcEsHbbOHcTzeJzjp+nLAKqdQwMEmvUPQIVB
7l29bTCkspxPZHumfiQt7Wo4MqZSqYHGY2GDpq5RnVBTywRLindceq39RyUO
t9JVpaT8SiebD1TDH6fm798STGEeMSZUUBPiIhzrB1L5lsoS6sqNweFMA1A8
EMvbipoVMyf+hy/j4uHEfEL3+AELIAiwj5RxB57L8XvsCphMjHGCcnGiCOVy
J6ikciklaxTLPETR0DUbMz1ZToglF5Lbdk3sIp6MJcFxp5nnnOcaoQ7eSXHW
cChzRif0uxlaX/hYBoM7a4pnCs6cXnrdkPvpe88extbg00N1YrLCuDJ14Nxl
CAcMzXm0C5ILg1YPF6A6eXCZ9hzCh6o03BNfQVbEfiS7wNWVzfLiSijsoIkw
aV/FydTjjjRO7VVkHtpbetNMLD5BH+a/JtHStA+w4kO0aw5SFmPOsLRpJIQt
3Uq67GX1+LcVcSR+Vh0FaANdnWxiHWCezyxAObOwqQiJRQ+iaWsIX+btv3A+
3Bw7wMcPgzt4lL5oKxauSlSSVsy97SXnEAyhLfh4hlM1KS1wy/tUf8jmoknq
oXcxKK0Vq/fRjB7cMeAzDhvv6GrPIPzwaVAjjGDuV6E4X7vUBIHFPD6bQtmi
EhxcHAvGLsUcE6rPG8p5OZl2xmXnYYYpsXTp3OfCg6mPo3Omzk9XyqthxZ/y
CB/L+/suWwIRSV8i1vtwQrI6G9BHyWpPAnBbvj7YZpBhI6eEvGxpIVNAnd00
bddt058FIYJuvLeN3SOkSsaJmaxdrHlORR3BkwqGNoW1hNHh0cuYDbz/wNIM
xQNCOgvVy5kWvdtIPYosrcaFDvltPS7C/+QG3w71Ie1Hrkywgc7Z4Xe7b11A
uD1TceDhngsGQ9nd8ZAR+HnmSDmm7NuD4IlHlMQLv8dytaSi7FUZRENg1ALE
UPPjFoYTLWVDVaZX9bdUn6+1PUR09RVmGnG46hE4Sk3UujJj8u9c8dCVFxn4
IhNFJKkZnlcA0v0dQXIiwTCZiWralR3BCq/vzDLEVL4OjjOINzXkq2Fquid/
8guZ+ukzzK2RIPTJDmEtIayMpYHUFCziLD8/WNPldPSgUtY941+ZUjlUYOzr
LZWNtRVVPvdz4IWUvnEWgWg48UNbIdU8/sSHhINICCgQv+z7EhWDI2E71USM
BcGwa1v4hNdiIiKqOlj7iHbUHdxu58m/Bgm8aTNRjJb8UrXz/xaXEt/ZdAmP
FY5FLIGspG4BJhmhgvEvz9glF5ejmFWZo8zLG/KFnQsVy8Z2wOlTcjytzkU5
rkgcr1hyC1eaxCVC+pc4suCT0mZMHuGT/OxSWmps8dnaGdxFOTptQw8YuKGb
kNskxeShScF3/ubR8Oxx84hszpJyU6B30Extp07MLVICTkLq38hJ9vrGW7L9
l64d3aIed3hH3aM9eMCk76tnGesTd14yfJ7AUAp1exD2UrlbkqG/ljg+3UZL
bQJSi4QbkrLA57QUYUNeH6ikFF9YBUwvksC0Pmm8umlkD2wDCbTys1ORauXu
9G2HozxzQyU3M1bSy5s/SVnlIQXjKWuXRRqdvr5bhi+z3ocjhqaKVSzyXNdt
0vxcRY4aOjZnoEVGdGxwm7jJX8kp+aA3i3GAD41HEuOWp2/b0oThsuGkB9dz
wMcHX9XcqY+48JCc/I6DXmBYdCDba7WtTlG2EJ8KZ8cGCjOAOSI1QGdiI+nI
tGuW515KT8/E4JOOG0/NTWEvZKunGiRfrlE3Kjf6ZchK4tNGro3rxT07Jnck
ZT/3/kq2IuHkseUFzcnWSF9S7cTTyAzqtvYIECeC6HP0NkwH4lowzisbPtqO
YoVaXY8IWrW1KykGAbtnhCwXOgFxXKp+xwTpdHG++dRgmbePpITYcsct7T/l
ixJibuWSkkH5ngOJexEB+GqGbd3vwF7M/6VMMNfB4DMkVo4lFaaVSe+RzArq
f74tWtPFH4LN4KmDWLFoOeUZFCjv+vml1Ulu4JOYGpPv7/2eMxPleBvuSn14
4MDMkKCc8bpvgTDWjjA1b2PFyJUlOnnYhj9Vm2Q5USzFKrfK7k0qMjyZohcM
nizN1zBKTBT6OhoBUUhWm7HYEeS16NUURqUoMmKuIiEJ95lnHkYGJzsuduM1
sNtUeQuafOphjDaRnATfkqQd39qujZTSlKZkBHpWtk/9uyHQ3u+T4xn8iPL2
X99wjm7Fm5B3+B8WGHWfCy0K+dTTmfj06ziqMWgIG/qmAZl/kp/OU7LsLyhl
CMuDc1rX9XBIJRtbaCs5+aY/AxWiMa3Vt7maBpwexi4u97EIa/XOR7e+ZePx
v1nPHjKEk1U7txnyRcEqnRUn84tisyTqHfmfAJ/XSSDnAtqPgoYKKxOPUqeY
XiyOVV/0PpwZUy4X/Pvt8SgVMU6+Id00GQ4pLyUU1R7x9vx8KCrfAyNa4V9K
i7gkLvBDLs39uf/+DjkaEzm8PDn7lgYPX3nSYqGnywu0+1i6HXdTzzV+wcKh
O+9fNUD8fIl/x3/ZF7ISwBkkqF3KEVFB3VeIxIneXAxQ9k4da4I7a9r+/FRN
EhMNuw0TxIyCXQtv1x0ni2mDeCe4wCtB+Z+RHyN9r/JuLlvwmwOEXZqy7A6G
8SipTtBSoiz9HQWMoeyXw1xws+qFRftdvMLVTJtzG5CyAo6QEylOvZsAu2KX
WMvB87shEuHU6ZluFFNYbIwnHeo8xkvk8DH1fSAz//M2Jok6YwtnL/PNeG98
D5/noA9nqOJYo1Ldiab1FzRnWDGI4DCdz1fBE/HzbnCHW7tGSyTiFUa5xh/q
d7hRuAcDV8ZXm7Nz2QhkvLy3+DHSW94IaNYQTblur37Ju16e+LOiCwqFCezQ
EC5d+ExpipgDFWpZRSBZV1mqv8Q+9UeJn/0o5lb2QXr8RfFkfTzt4bLiW3de
LgQLkkIx6vCyO+gxFkfawZGFK7faT2QY6srYCAjSP7+CS5loP3uXjvZ/nRI4
zcEbjK1w/UZlXU/+eBURLgugKIfCqIrPXrLr+YU7y9IvJ2hCp5F3ub/1Kx+x
nlDoqPY8tUC9tRqxgoNmHgafaqpB3CgabSmh/F9YJ0Ser/bVL98lACdXxs0Y
xeT+k2LsXToCKhUCtPoFCDSmrNhzJsECbfOJ39uMQRDra/sG9dMI1zjh6Gzd
cHh+sQbtMN3qqLBqsj5Ykj3ThstQAcrrXy9wCWLKKLBovTxPYkPTLdIlhrnZ
NVjSxa6yu9WrVvjuVsDniurLQR5TvgjmtnJU9OXB8SZ8I5djFReE821NzJlx
+DkU0RUarhZgSLVn9dYxQdXvpGvBVv4HVtzhSdpeayCrPBrnEM5wk4lBlM9p
atRBv7JuNgLxd0wy5Bh4GqAaGonnCW/OdMvUpWeHSHb2X7EDMqR/+6LxO5fq
e0ORLd+2SVRkXMGduOrU4JUEs9lilxidl0ui1T4QyLRMRO5urf+JY91oFU0H
zUQJQUa91rkGULSl3JDto3fT4dUOG3xERF/VqfSLJXRda5uP/pvwYRfjirAM
pQl6bWXEE5iacdFh+KEFET6bC0yaQg3CXptqmSN8MEQTe9sEshakN0m+uUoz
eCLolsu+BCpZyomOZumd+o/Lo23xdOogfXEAXU8OTMlOqeUncTZmm+JRVxx4
0Yh5/gQqBfKYYgMAqS8H1oFwNE/nl86PuaaytyKaPSx9hwN/eaLvlnCgWCnP
cozSNyKmfcITojkdz8s1yqhtkU6Uqttt4QlD/EjiMdSV4B9CPNb9V0+HKQGY
yaWDubkp7aIGmoIvapxn2AG4SwCK4dyrp/AlqOSGMcbWO9iRcFwUX79FQcu/
Og8TuKO6zUiAuo+knUEfjUhvTtGTvP/NFTrgJmpLurCH2Sdofe/zEi8SohI8
l3bMH+vl+4RP3cSSiZySlh6buugvGTJzsT6GOfTTuFzgxO39T/EEyKFOUDlU
H2ICAnwZZcg2B6lr7/QI4H5M/9XEb9igrEdmSzyjrD6AisKq+iYNLHM113CC
4r7llAgbqCkyq4uuPm9ynfFd8jbtQpvGe2jSCVUqsNqF9I8x7lwKC+lGSsQp
Iv/y92qcSQJVECIlwTgKtnOWH6t3LGN3xEZs50IucSDlUc2GADtp6d/7UMeM
ETqoDGNW1WnAaDEXD3HOHMT9995i0ESiqC7BWOvZguiymr3xhnw6pV+YTWGt
OZI5Xbo8oxts0RGDjEn+4NLnPzufh/9ow4uOsLEUwizCJ7lMW+7GzhW71+G7
rD9cSPMzjEXhXaVxHfygVwR+atKGyIf/wBXpX21w25CHTdPUjWwXgqmBzZil
F5MlcYgC9SP6TIwUSmZ5K7sDWEembRsqXU+uItJdiAxvvmlzg+elavLJJmg5
c3LEcfavGVi+wr0M6cpbURZn2HuTC/t4smn44inXVjX9O/leKVXY4/++ugJ+
J+wWBVmOQSBqv8JXecfCFuC6UJ6TIOIpqgLW2MHSkQjSrjAk2kVjTZGFIP8W
HaYqd/Mg/YPHgoZpwalJPYpAbQTBD+GTMRb/YcJ017Ts/o81r29kGtA3F19i
BzQYa3DY2tLt7/vslSX+9Le3N26NdNsYf3yu6XdCqBcScH/4gejaunrFe6gN
DDuAW1C1L44bd/vDxYXxXoK9RkVRTUT3paw/Xj0u/mTvVwfFYhLx2XzSKnEn
ikqJRIlH+Sy3LFDbl3P5ydrflxjrleN4vqs6F8TJ99suG7gLKtMhaU0v4WNl
z/6dEsHWiks3Q7sKOZsyOu9zJ/RZpKdANLwbVjNTQEeQq1hdfujG0MhnyRtL
R0iI2TXh7KxsXmYwjFZpNgFWrV/P6p8nKBBYhe5uDO8tgIXkhK19QW4QG23Y
0OHMhnjJqROhhkwRL7ctKkYD/6FnBOABJVBf52DfbHQpo1VeVAdV0b5DvfDW
TsZ5cdSDmjOT6rxuHN/HE6ehKR58tADW01snLAOa0GZJVAQ7aPrJmwuPpNHq
SGRuRL9xJKHjce4+ZUr3BNEj/t8+oIwhkWJHbU2QhT3aflaeJU6s9oCtWKYX
ZpNfBrf048dMOo95h1fQtVbZNaH1+9wTVsJHkxUyEuzPsT0Y2sB/TAuujZfB
Aa2QrIhQH1aJTVStzVNsKpiqRNg259989/RCOUfWTjDlvTRoHW7IdPBhqqlm
4fsDi23FrKy8efpTZ6Z8mPWUFeaOkbmCgoyKKnToAB82IBls3ZVGokQbP/PA
OTnID5mgV1CdPUheX4Cij0x4q2IIhFwBZjGp6He8V3y5aVcuWi+FkSyJJhF1
9KUMghQ8r7Vn1z0kV0V0Fb6JsxaPrU0Fw4ZzimJXtdSNjb0TcvwYC78iuZ1u
U1ynPBSsU4p6Tyc8xTEakR8jPvJqUHlw8DP7CtB9graZ/J2D037kDXuV1hjz
bCvTcImoPKcM1na268kMfs+YmUFzyOekpoQ1dXoW3LA7kpx86m7C1dTmjLNG
q8ipg9aZ9Gxw2XUaOL8hrZaS+u97j1QUJTDr+HvjSmd/WYp16dtLSaQVoYL6
mm9Wwbz2VyFNUXQXL+0xy/yz+F8/MMwaWfNLcnvZfiiTMJAU7OdIppy/B5bc
MouYjMiMDkMIjA2ACP7Roj7TWWfEloMmxJhu+6y2am4oJYyNNk0Hg2ffmai8
iYVXVd12bUvhHfJYrvYFyrJXAbO4eKMneiWkjGL0prEZ8/bg/35jB4jKL5aT
jiAwyLjWgaSyoKkGamdguw9f8vSZkm8h8pSg3750P8netKhmBt+xwTTcRuUK
MEICFyve0Np1yfNrXvovB1pyrxWivpmPIXAqQSWeRWni2Y4PgBEFA+AxQSwa
mRFV/vFq+qPaaKzZhCxzbgJXvXQ42biLQrbKBS9ZwyBF8bqIklP9jKWtf38h
X/uvwXG8wxUqnAbnqyZNn94/roD8V2IvKLhNPdcKqazl3azJuc4fCofeyL2J
Vy/wHdW7N3tldwM9AUULERwwb0BdhtXw1jtA3gJyUcaSE4qiIvfjEPCL6D6l
1gx47ppq6NNwYumUZgBihe/zxMSpYDkanLHrYbPT5D7hq2rRJbqs7gSTZN+7
V8O2ILlb1OcBj6fMO5F3WiC3On6wd+5naNMmaYqNLel1pdYDvXXHI5TUatLz
pmIqfLTkLOgwFQMBKJJHbWZWXT142P6mWonr24vbznGwVnyGBelvCAvwyna3
QQh0YjxP6Sml+h1BjY/xxfKlSlndHBA9FwybUwKOIJmkibMRJAJG5l2AoDvf
VM0AdBOiOlcbXWyaPCN1Ne/e7+4o5RPQTLd4akb/IUqbP539xIzwPFwK0/42
xhEwIubGABbYyNv8z2qNYAirBSQpBZhcE6HaxtBbhdrh2xJY8naGd6w8fjhj
3cNaA0at5UKZA0BLdF+ca9MA6502jCwzX5RDBDueQ8w8n+vLLReggCCo2nPs
1Ms8uS8Do4VzFhhPgvFSggT1qk0um93Ls1fMA3IsizRXZ6F/EEyOQbvkilrS
Z5vpX0LDTLEmiIKXtrdI3gv4vxluoxfyw0ARlIlzuKdGXEL25qtSgZKkuGa1
2ocBas3nc8g0OnPe4UsfRglfewOdYEWPJ6lpyZvM9PKPVnHcSFvWWoPu7YDK
rL5Z6B5jIR0D7e4aPnNqRBl4MgEzeURmFDlW/WQgWNhAn8K5Difjt/N7qLtd
Re0wo58Ia4DjPJKkFYhZFhjB8fpADBJbtVG9FhMlzBtTO6xjl0whCctICfnT
g9FOciG4ytougsE6zx6juYQnLuG08ciFPIYHZtF3n/fCJrXB7PI6se3yyw94
zUaq2kVYnvLd7/Np1YxxZnHYgfkaLgdyOcPQyaBzaIrQf4PmVk3y0AsHFaFN
87YNGuvkKxZiuX1SNx+3F8L1YmfYQrT8VFSiNbFmPtSUYQtUhf6Gw+I9t6eF
iw/Il3ffVW0VxhD91IafuWelKC7jVYV3D5xtLJBhBYpsHqotMRWGFz/drMLW
sLhZVYNPsp8IjIDOebGxJ7HjE+3Mb78PBid0DRjJ6o9ZiTXl0LmSq2N6xOJC
buQpNpjKXhfd0BP/rYXRTPwnABRShR3omSIUiL3ar2V/izl3Ipk4Exzk/Z0g
PcoZvwFQzMx37SRGAnCwc0w2YfpEi88nyCWYh89EhMwc7M4UmjzGRPQAy45U
2QSt24D8kHbEbWMmzvzkeTneA6qNxCIru/ZEw9ZxnZUJ3t//5rQqR1NP/3ci
IVJOje1vF5yxSxdScgvMMGJ/5Ty0N1r3aQTx/16eG7w5L5U47Co7v6WtVVrH
G6Kdc7HU8yEVKcCzUkBpRCjjKB7QOZbEjWFdLmDDg/qp/ks02OxhM5K1ameE
LfQqukO/ctQbLhROQZXhfMUrDOu4OBgSgkKkZdoPjhquPtG3GDfELxapJSzY
bjQ+BeP3UrEHaTczYRe+zewW1u6LJfXg5OfHuxZ0u/dwBr0Mw9JSFfIHIrIy
wNVgFNRQHxTmn2mQ4n1pYphPTBeL4Wqq4txlcUXU49EfK8wPZUi+2lDRdm8V
S4zRZIVBG/iHeARV29F+Fz3Gw+Op6GiaOuQaHscVliJPWPFQSE1O9cVCAs8l
IJRCbBJNGOQjLpdi5eRmth46WajWhVqDlQZjPgF7DMZRjzt8o6FgAo3zS4IR
ahbsmNiNqIysGFUkfWK7syjYuADTX4e54p0cUPTA30Uwlfv0dHjThXZ+MWe9
v13y9GXz7SjnwthGYgbURe9cl0mmuJpOMCiX8J15g2YWASY9y0uEhzBsnCpk
yZPHcOiQZNk5mSjjYS3aPMDcobAMt4GRc/ertkMq2Kl6TNZDoiRFtZ1JHm63
BWarcwya8+PGlwDp/mX4MFqYvzk2LAkXvm5U+Chsju55KCVko8VmEkAT6l9m
KNkHtTu4ALR+IXRx4MZNuHAhFFGk1B0XuCC+UpXhm9DKbIATlavajpkKNUJL
mr5mdhDZXY+cjCpfu1BydsnCYliarvHnRDgJ0dxoCmIuM9WE3lKUHAuEANke
uMhNp3aQN1mcKx7YGvsqq03WSarhyanvrZ8NlHDA1H7txAH7wyyNeii37uhH
QMswwRusyVdnIvn+fhBaSgWVUwu0jyJZCLreBd1AdnO2uRWuKAqJah33hlu/
SpeaPKC7XO3y5hqgs2q5A4ncAMxhArEv/xEr6REI1Jlb5Te3neKFISlgumNU
cp1izv7M7js8ywPwE2KMuIQrC3eBJTFIkkK8c4lqyu+El3qTXkNKcMzqprXu
yPmT5fmrU2noB7/Vvqgl5ljZlHZNIgXIBtvmIJ98b9eRCgYd0XENcbQJf8SW
+q2ue4d/1hcP2eP4syx9ehDT56kMy1C6D1SuyL2BqknrkPUjtFOthFo5ZtCf
Z1rBDEklQroXgSHXBxcB8+9U689n88YtHakOcZOU58BywNuKxROJYkuTYJvG
tn1z3m30XUIuctKF7cLsjtR0tjeFyAYAfefF5NQt7kfVOona/PsfY4NtOE5d
DmIdQgJI8hLg/GEKTHwu3afHIIlNovXsXQgS0Y/W7cbgyPD3rFktEfjn8DB6
F/a/YNQbPJ3e2gOMwBXjTBAooDR9oPWUEBajrvycETnIrisnuFYT0Y/GCEYU
LTFSP+/Z4pE6/9OJxAEWovgAM2s+VDn96RfmTZY1G9yPhN4uWJvU/igh7aoV
wW3g48UX99yBtJBFiGep9HW4tGE/EK7lfOazDyQqDxJaped5nLfnWz+lrT6B
q2g5oAJbctaNM9ozktl1TqOz0CAw+BdoovqNWBJYSqzJUmZ7u3qukkxyqBnz
QFPIp31caqg5dR31O92canzClMHd8xxgVYO/ZuxIsW5PlhVvldWNYcmlAvlw
ZfT231SPBN+RsWQoHN3csSHJmEHNPSFwu1/dCWwmo2k908V6hf82ypvW5zvE
VtGaq3jrkb4XyxRSbssMkGQqumGjEFL7k8URV4ohfLYQ7Bd56qrUAMlQGDuU
GSKC3cKTVhgGOGIWNxjYLgvJG3zqE6QFUkL3BvIm2pbwtgYySBnaY9VZGUad
O0pXD3vpZgoB3v3ug+PcOLVDVl5LC0k0uuIMT0HsxE9BwrmBbSu57bnDfiRp
KuxaP1ADnzD/Olwn7sjM0QsCNQUVYdkykCa6OWuDS992gYmspDbonMbZaeYR
LBxF40mympG4P0gCiS6DNu4nTLLYVu05eduRnbhZNDiY9Jhe2Hg7Gr0+R0NB
uabMqRA00fnGN53yQYPDJIpcNBGOjDLp6R6FE1dGvQ+A336TE3Dt7L4RchE5
xbilpSth13BpuCDfxScqufLyETP7eEX/i9zeAMRbLzFN3Df8MWzBfB81wcOc
912eI2EBnTwnsXAiJ9mKcUkfNruqZqsX4EJD14FtaSeQAsX2QAcOoEWu8PeK
tl4d58lYZUYvrDT4413AMVvn2xKuQSKzDQO0bKhhT43Ph1wlOJFf/JsbC+Qq
km2XTr8a2H+FFiVu5lydXnQUCHNBITTwS78f6JCK4q59HHhl8Rr7UmSlXqIJ
UTCuCBpJnpQM5ugwU3E46oq4SyQbYYjEY/tnBwbV7XSuFYfcIQoHfUtegbwI
znLeyGSxACuZqCtY7OgCXdzoOVyLE2DdkpCNPFdTwIEndPU4yH5kHCYsrtKE
s6Rn0n6magh5OeF4ErZgvyhN2D38nOwUJ3InfRV0TuAnCbtCzlxrJw/lJL5Q
RATsAog50VHxSKqzzzTNSmAr2bX8jg5Z0x8CcOPLrKJBmJslnpOmYTej02tr
KWxsEaiWFWOX+vFeRiTRjOugV5yUdJ/BFIb+LpRQUGYFOj5l8+qtW2Dkqyq+
155nOg9FTU6nO8lSJ3SstouY7/vbQj66Lt43WTHsSC/EIgowWIrw/Sk2qHyl
09/oxj1V5wBnqg2e2xO3kcYNIMLqVOdjHKcDBsm/DGSoE0XnFvEwyyEM+NeL
5f5JbXJNYhxxhUhe1BioLaE8W5DpUqHay3zpetcCHrZlE371GwOLRMZRtsiP
aL6X5uO5stME0S2TicW+FJb+SoWA8ZEqffAHOGH5VQx8x0zqNAHZs3i69tP9
N2K79bpo1vqActqJPfCuViV/+kUGtKF4tabX3Txe4VLiGfIEZ3Wp56v49Dp8
k4Nm9BC5Pwrk632+oZFWLWh9QhB0OKtt+fxOV6fA9s+GhR+dr3ZPuYQQhmqP
fxpxqkLXOYBg2a90m4n/jcRXteGZuADlRcGBYCkNYsTjw1dFbEjkXhMv5/W7
yIzm7l75py7tcEkLgBvIIY0b75WtXYWyo94NHhHC3dirhsiZT+tyhXvtCsyD
noLWb/s7lIV0w5JzxTl4sbSA6zkBjTUF0F5Anb6qvrXJeqrlyu7pWVWQCkCL
ohUwDOzpAGjdeR2Bm/S5RHQc7A1JTGYdYQtzOoDZidxN7+urs+6tAKl7Tyr9
4B/0Cr6r/AMddLCN8MoRzof+V5Nd99YFh9VuGmYqK7urPErFy/ms/hXzdnT3
mnhCKvJOHvlN3lzv0ukEP3bg83gzWFycPZESfHUDnHQLJOrz7mqkVy+XWf6A
00Z2RA/qXRfXt9K789asQCRCYeY8ZWVmg3Aem2IrEUhtnk4ccr8+xerI9MLl
uepWTi8L7SmvPnWk54wxZv/uOYS+Wr10plYtkuaOUsZ7It5ChaeCxp79KI4J
tAdS5GV8L4v2zk9+72DQQsRFMpxTN5Hn+jgXCJzQ7aOlpGLe7pjE/yIGdbKU
kS//KyWjrx1Knx20BE7xfngHjMLufuBo38Qg1eOwRQWo4cUk18KCEvLGAYGa
L+dEe+jRIl7QUbsNyqvBOSFMNHOmxH0HizHbsIkqWKYlgDcZXAUvHhrRMex6
5r7th9cubjNVIhoMiUyD9Jcixb7Qw73fnGfwGU9KHWOfKdTMSUKrUXusLxvN
UBnrpRsrzmoKU3hhPgRcpHEk3PXij+wzrsEzxT6Idu1vInPKZqYPDvdgeLBe
JKrIOpatThrh8BKVTcBsKrRrba9lP7qjTjxXfnoqNTGb1nrYz92jRLNDrLzo
HsLC9wWYmLIufLfgUHXpNY5hU/g6BoNE49lI/0dr0F3kzxYNomfJwFBGn4Ua
aNo/YNzGK6pSuCXdPQ/lKc/daZ0aUyp/jhebpQZkcV9gEPqbFtLaiuOEcp5m
izIUzJbj2p7A7gLRUlZLyBIi52oVcZm0ycX8uNTPNkoezVNiATzzIcU9pQZN
vuckfyVfuwzbv+oxKqOoQhT/j4SalNYRV6bnzhdqjEHbDfG7dY0IwLypsNXl
BaobRhw/E5RQowKqAgfx27gzc9L5KbqkOPxkDe0UyYiGd6oobowfsHz3hfF8
OvIVnXDtxqe/o30RsynlrIMOoIjGcjAsIN/wKxIzIfQmsbFEqJDBiZdcThNl
IlN5c3B77JiOIb1/W11igAwCAvqRTw1M72P7pu0XBw/g1+OTgilKVVm4viHG
rOIuOuZvMoLUb0zMyAWLFXuClGKq32F5xEtASHLFqxiKdAyUGitgK840JWo+
2LCHO3cWNF8l7BHvqBfEfppBtTseAhcB7M4D/xuO7tgAx2uDl22W0LT11o7C
WdyOYtSg9J0162XX6tYe/Q+D1zZbNiUiQ1BWHM4WytVGhiPw9Ayup9AOf5J1
I6ZYci75v0l10lPpn0ejUO80RKFZ5L4VbizVkL8ltDWof5UZlm2dxKAPHtl9
RVl2LxdMRD8apkZar2hLyEsMOZ753Ig/TPKKTcd7wqQQKitq0LPI4AYSdi6e
egZgd1T8hkitjZwVEQ2y7mkWv0DmWC93PtTNMxx1UswER8o/yyxqmETzCtcL
x/u7L5B5Irne37u+zyj2b8gtOJfbBcBlktyN0tXUwUkXJBtN8o9F799BuEjE
I0j4yvxODWJb98RiRzos4O/XuGfqh6aijFwNfh+Jl7byHRS5Aicxi16fp+eN
QG8ZpbekUgpVzKYfJLgJzitQjMdIinun6FQIAhk+EhJOd9hAQTj/HjTzaQ+P
EM84ZQL3mfuiLuO/fwIyLBnYE5GP09EuZYnQQvQp8YjDWd1iWC2II4qIIOPS
9gkYkZZA6yN7CSJ86FGpQ9xfjVrZ0GKjwMtI5/2SKqavTLxIetQ0tnSNlQyE
b8oOE3XpNE0Mac3S0oIPrvasL3cxZm66URkeGaClXuavzhNzcS6Lj5ZkerWf
nUs7DPqfeP7gAKaoiP77YWgypq3XOeTXE6sbJxh1OvBZNmmpiO3ZQVfhd0h0
Zlw49EY6YEozN0GMC4du0NXePfpmu6LY2YMxF14rRc/Qwxx67JYmzjQglNyH
Q+B/w7JiSrJTvbvS9+O4gMZ9/arx1AMLjq/HSEVn74V7Qk7oM/7kHKRsWEOL
hzOpM/pKJ5rGbfUANsNZzKrWz9mlaF8uQ7dd3V6cxj/TXU2ELlznjO3+QbAr
Img/Cd6UH+5Oo7PmCF1iek5d/YiQeWsmhT04CAtUWXw0Zq6mra1aPp4JYeJP
IVIzQpvsPFZm5FKbi1zkiXt62NKiZt13RCz0Lp84vvtxcg9XXkd64eIZHLSH
H1WKwj+r628l7K41nD8k0qxoM/xI5ZBgc5dtqOLLXrsPJf6lwkFzlvl09nb1
3/dNa+j3pnZYbtZAIQFc8JKS65BmQctOI3YWfC5D5Y9vHkPffdbVqELWOv4d
og43h6un8mUDQIKOLrSp0hU4iPobY92pdX1R6xO0m+Vi1qi0+BlhNdUbdoW5
4HUTCvMbpQyrn2RSUAh85aYyMcmza6RuovYgKOVCOk4EaSvR52mB3kQsbo0r
DyRaitow0EiP2t2DepQNeBu45JnLPy07pXZjsb8Og2IE4SOI7+dFf9pdEN1R
GbvFbovc6WdsaTzOSedAca0o4n9gRz8V2sfBeBxzreA3vRPUC+ekfS6l+jm8
97sYn84+43pRSfOnhpl+bhXk6j28cu8Opm9mdDmZu/8RMGyIaLgxXdM8BCva
8OYrlKdv6ro4LXFYNwtLh6cnhIpo98zEe7Spr2amAFb8RHuFQ/YmJA3BjSpC
M8m76qAsWMm6IoCHKlv/jB8reX7fIm6QwFvU5Gc75ux2huM2NwVRD2bc3pnR
lDdlPq02Y6wRA38CFdUG4VmHHtU7gIUt2Dp2VLX8vf5FM3q3vdJlIFJPRILM
sOsJxzHmuTcPaxsYYGemZ3Qjom8xIRZhnGPMJSmkgth2ipl2q33NORhAq7oS
N8r24cQZSkJdoq36sXkxPB2AE/VulgZ1u7o0HhWz0Yd1FE6+49PhmCXmCrlY
1l4Pv26P9tl3qxE5ttpgbXi0gpL3JkdlMWmwHxG8wX2Ibkw3ovujMgkmq3ZC
lqXUzgNVSqWaR1NZYTI3rF0Z0hT7k+T4ecYrO1T9wHrBK9PgqIg5KrZLS65Z
h/NIb0RktoM7pQC8V19JqjqUB65SqAnjjm1PUt+A2yG3OVj2bqF+7Ijey87P
E/O7vhLssOqcKUU+5nghkVnI3jP4FfCkow/lApGG8cdH/w2hemjI3yFbUO4y
6rWSn8opj8y+0Mu8G1MSOyHKY+S+6DMmYKghUS0oC/JVWgXvKXa7bELiUvcS
ak7Yp/qShEAFMH9A2OQDfvnL7QDL7/9UqtbSUx+XoSXG8ZWtc0oE1HyFCByt
b3ZF+o2bsfXCebAehU7qeH4DF2yhZOSB6j2fXqJWn5u6UEtY1wQQADk+BC9N
gqR6xJBifzqUnykWvb58kX4LIHQk1FN2vf3DsDpAL1sLPh0gK/QZP81bTmjz
P6CkGVbJnsrDNYEfN5atcd1qlpEGBJ/UIPLwq0Buz6CAP4+fnu4KiVLWw3lv
oKLKIy57OKJ6cNEpPlIOP/+9EXkyWRRbpkosmCqyjJogci0o0kkTSvTBKoMj
ZbwWC7SKT0T8hFBvR2zbkcO5aanUc9JZXH39Dl2quicUU+EtK5//F3gGXCCC
KtlPD3FMuJqW8lkqSYwr666jXqbnacPhA95GceXJXbrstEcwcvNyMIsaRrDL
K5GuUaPWmo61I0N7DYr+EmdDQ//Ra8cHmy4WGdtFCrr54qeUXUvVaykSm/I7
gr8u6Hj61mZoGqSi7FML57oaHYHtMOXvXLvryVP43x7yamSM9HZXmv/hm7gj
+ayj7kLJpqO/GR4PLEvv+arhkeI+KWee1znCjuTruqjL8SSQSJSV7sDZ7sCW
8MF2cQHwOfx5lKWS6+OKBDH3AcsGwOzj7nMQi8GoVyw03Z2QzinLSxnrSZrv
9GxXp9HXnwIpiBq4Zyku3x2SNKHa71rCwvKu/psxQtlh/3cnePrO1Vqjh1C5
N2dX9vYWQkYilIV5Y3dc71qJi6ilNqIsA6YYcJtFWPWsF9tRyCAQiS83bfaX
+0ZTn2JuLoVg5Q7dJxClqnnTuMOnoz/yqFIDHQE3+7vq3vhBdp2c2nTyLLM7
eyGbZBZXrUVeE+qrWqZ6gtJZ1nqRK2l3EEG6/rdD3JROgAyr+xBuKfd7fWdz
4xnwM2xkWmlFy64h2lupFl/muRs+0BjVFoBILJn4yH+jjk8fxtzzj5yg1evW
mFDgKUDAHnmsuCmqQZuakqR4kVEMPJqelZslnuDEj7hbO9510vkT39jggRnW
GqESCcr0oD992bBQ9AbA+ASnW9iCHsNbrLyJBdaQS86IaFyrUDMI4c9YPCXP
QTwtafiGqV4mAqxehTB/j/q6bhgI7AzF5HJeXKo6K71Hb8MnZZtLjxM/uMTV
vt+ymJLDtmzsF8fHwq3CiaFTCPJ06hDEqVSmoZNdPxzhA+2ZY4cXE/UzxBOU
ozVbtgagBSAJloUfgiupxNwhi3jIqZ0ayzuHu0fH/nnGbx14ndfKDR/+doEB
QMrioVYRZwYr5K1j4nlrih5RpyLxHpiCYRvx2Z4dDx2d1MMLhjt0njmVOeAh
db8QVU74MakLmM/uCTzzAWcynV6Eye8TTteW3gaxffjSOV/y8MfyB7sQ5+Aq
NmYhYgPghHejn9qiA/GPAMxyf1ztHWz9ZoyPEfm0QLOPyAfWxF9Bwo/GY4F7
2veNfmbTbi0pO8GXwSSWOgnKV0cnweuKhUwlMuji6QeyDGeq6TJOp1T4klT0
A3dnl/SRqZGwNdH7CnGR445yjd2uFsEc3CarcWqZo2j68EKmPRHIeaM4Ga1j
vlIOQyQFC0hzurM+EXiRlwDNCQhCgiYrdt5cp3Gt+XSGP7e3sx8luGGWDx8j
GeS5a1o1Pc8FkcwklCUqKjGyVedxFchlz7sBJozMbmQpo5ojpXj3LhLZrxFY
4gmROEnygkdGcQoIHYtrfr7y8mIgSQ7e31py9RhBuF5q6kgyOHFdbo1YPPPK
r0EGw1j8HvRh1rKv/Zl9BbzfrqaXSdHeiyDjEyHDWz8svNovM2RBveinDeVe
e1n8GUNvrtneGzLnJ+UpoRVb/fCfPvFzn18Di641tlyYl1MoD58oNSOQzHqB
iy05fRRvQaZIGExTZdx6tburz6OZL80Dp9VxJ+3/AtcGiS0daMlYCwYs49/X
P16YUv0XbXVvCRWgWYVV3k8Kh334eNGv36zjRRJKaAd8d2B1JMiHssKKP514
SrzTE3HLgMb+SqQJ5CSQmEIpdeHavIiHAtQtxvIkBbz7eqM0upG3U1pVfzlo
NgGQCLQMt06SDgghNzVG9e+LBiy85zBVXtl/6LvaBrwNkqpLSmeYE05dhHNf
8jTfllYVOjEt4itzIpKow0V01GjUWT+URf73KtJm4QiQ8kX4pJqPhubonCPW
R0o/U5jd05X9lphPedErI1LMHq0btXR0WefMs8EbZj//K3GGF3ctgDlUs5Kf
5RF/2835+zDhh73mXg78Pfdp9abrdCmPWTkpFON3GjBFKbnPGXLmUdBiPJm0
PY85rWDw63hWrK2CyZEzbEBigY1IZ8BS8wxN5R995Ja2B3RfUFK1Sgz3r/JX
65L2pss6kgKpq8onIfBwQBvohd74hGWY8j0+j1TX7IH6dqTRWyrIHHosizNv
JGeH1BsfEVl7E02X/bTxn+OJYuj/1OBFB6VuFy7gqMq6iSOPPtYbFRdnhRzq
+EgfSh+c8XSv9i8CjKUYsPH5soPPLwv9m+DoCOj6FAV9053/ssB7Q5Ajsq8G
ZLrt2O83qcc2D4Jk0wb4/mvfisLm2JoOkft2uwUGQKS35+VaEb1m4ucGW63r
Pa1TJjw0RZVpWoZVzL+fubCCnZ14pgKbYgxELED1qHkFip13dud/gitq6RX+
QSLfVTiqiZQmP9VmI5TTcPIGuZt0bH/OpJHROBTl5ruoCjCdvywTwCD2eNbQ
9Z+2h+CtkjBiwkyp+gt7F6hbDmeDS2tBcWjH2ajLgbFCkyblK9kSbg9TAW20
o1hfBbmyP1tPyrL6P302qn/QhAGExdno6zqaNapVvknQ5GaDDbg5Y95Oa/Ii
WlFi8feMV4fuAlc7VpIAQYalf7XKVZzUk5ftPy7If3tKDUQj/6tXR0yUPzUS
DRWl+18zr8N7TOqWRFD2ht2pNqkziECYiW1HLhVplLrlZQQBv4hXWt+MXzOR
j7glMTq0ajHbIxzFSM/YsVANXljINRKTWNxesqOz3JWdiNPAGqmyzNIDh6IW
XUIYBnyfn8ZFYxvnqbAs9zn9bcIFNOc4BM6ctw+CwxKSJb8DGuVMKjJBoxfo
rldOzwkOIZ9zZLyL4seNyqgvmgJzO+4m03mRBMNcdeI67M/YbUfjGadOo9Lz
0UD7+a8XvTLbLkfqyFHq2HQbOxYyo0saEgEMkAycq4+17Aan5etY92hKbYPl
qwi5j08ysLnShWiRXAfUCKdWBIXo7sSOaA9I1GErg601zmrmX+fw0fhbuLTP
OzdH81kZ+YeOCM5bDlpVQ3HEo3XJZ2Crvm1UVt0DZ+ph3lIa3Ns/zmL8frD1
wehNFJ2uOY2eVvJoGM1dWFShCa4e6JJ5iM6LNLmv9NeyqyFcqw1XhVmMzBan
uN1QjHqiUCkMNbRl3rtONdkXlB1Do4ML18jYO/yvAAcLqjTxuEwNRGAUAsq3
mh/5k2U4pmpjupamAI+4mgK1bIDUM427ZXStJ5NM7W7YtiWtAMytxp10Hv7j
WeoGGnv/cmMFkkUCmx18qF9VhHKcPXsrHsIx0964ffBssPgISRKYnQcMnAm1
LuuGbAvMqq7tZR5jfHhtSJUBY5pvwOA8vaRAvf1QpwXreNlwD6DtwlyHDGq3
CS9u8ZTV8O0E1sMQf8bkJD/s+h8+XlJuy5dwwRKLDe7zg6diz/jsySW21Gei
aktkuALMTfhLMk0asJeGDjvtdAkkwobkIfXlSEcd5j3NZb3oT398iDpsBHPV
QDZy9Nd2U1uV3I8kwVKRNxNFaaney/ra/n/KXs6f7UB2ebKwNU85dcQbBIcO
p67Dwr7++JiaFaFF3pIMxm+ir2D+kjlhVBQJinSVODZIz6OawAMkMXh7sQwb
vOAcOGQTLH8HnoUvfK2UCjpaZufVM1AOLZ10hSgG0uWksQPngztSKcbXAUNc
DUqwK1+AGiROIhY3ONa7Edd4w4GyB9hXr3XEGp14aVT9vr5fPBFanqH/hm8x
OjqLN78fplHY5qBapV92zlUkOta/zWDsaWaUXgQqrsRQzurKPof7ZwByWuiE
U/pLg2ho7ZM/piQgWuW3CrdvsDl/14p2CHvf7ck2FEl35uVV9iIZFLRDhwv5
4s7g8dldlbie3QF9W/fwn/qcqFhv5wXwBjXJKpMVkaw2ZctSXdTD8gxhJysk
foVlXtj+Iai7cunu1Iyj6/rFqJrTfBBMRngNx8lpy4HMktxxHX9WY47LXUh+
1oAQZGesYfO+fhnPOdXXz9SxCz/HSHDNono5/flTsB5C281VcSsBr0FHtxgC
8k5uIWcZE4Cqsd+nJEWMQ2kp4KRwdQhtP3IL3kjwXqfTC2UU1s+/KM36nYel
n7ve6kuhF7p705TNh3bvZSNls88bzydJ702vLa6Xoz7ZYdCitxPSp3JsPTy0
P04ihsPWqCStqIiV7ChZvleAgmEbp1kKcT4BvFkwWN7WjUSpMi9/cYL2eFEP
GakJDG8f5stKvp+KxMnHfp3v295fdLiSxO4wngKqF9Y8I5AsYvXGp6224sUa
HIYiH3dyokEMUIr0F5NElRADYI9H4PdUZkqV0ryr4DWZLLaLD71v2SQ7hDlC
67ZLxs2bA+aYvIs6YIOCsNXHRD8Do/k2k7DW4IWKhCmwFB+2dV1mYhvec5Ne
jSrnZCR0t5sya2qupXPaKu0zXeT0ViJKE0WLL8EhOvLNHShIZgO8klZ4JS4G
C8Uwn+lVw+ITrAZaC2pe7Li5WwotYQUMFhBF0vwHuH+/Olbxh4D0IEcy5aU5
cnHMvvBSyT6xMdDCP2HyjFFgkaa+8SGov2jRQvLJX9XuHf7+kFbRLPzOZaEe
fPMaYgk4CxYCWOo1NRKqk612XyMmK9Sl1fbkbHMfbIrSwP0OylWVhVx/oyQJ
mWzQQ/UwGjw0xZYNBhPmYlFkmyahoYtMGjFmiajQN2+ewF3MgZOb1aDvdhG4
WRcz6GcZCzHy2uf9n7u0mjhbsvaBeOdwiJAoiUy5jNW3XNl1Cwf4Z4urWuJ4
8wXZO4G+lmBymBy4NkeuksowaGQD/R57O7H5UtVKAapJrt0dKgJXEI8lgiSJ
v3/uei/rBkFo3fWcCBg96+POsCjxzjvLaWrLcS8dxsAn7UPRKuAMdIGz0rdF
4j1ZgvUMsTUNPrn1yIcl1Jp21/L7B+BniPLnlW9znj5+ctRRrRyObaAiskrx
u44jVx27QwS62O2DMlDP/Fj2xb2WDIEeq5hOEAlc+lavyOn1OmxB5QusOGoN
k8n4U/U0Cnbd8HknMEKlgNQFLoPCcQRn4KuKKHdBe0PJvGW1GDr6Gt7fYil4
sevpZQZyjZ3iFry8tHNG3sqTCXF6NovYVF1vD6cqUChcFr9VmX5bcM0PIw8Z
NJS/elYPnWfAcVRVIhQQF2WlUrMea+TYLxk48OV4+fV3RfFhslTyw3wzfUIP
ATBx0w5jKOqMHT5H0fAooyr3NyudXGJf4V5e+r59PdYIwCUP+93I6gRDQcHL
QflTKrgSGEQkK9BByFnoK9Xqwk3t21TyAQo4f0R2A3djHHVlxxpFfRs5FaKa
CZ+F+r15rEgn+bcqEeVue1LFTP0sWYSzAOPYaQ+Bm5l0GyEqTvGoWfwgxxP8
5Sg3vWKwkBwS41yK+qWD7c7ok2P6+DqVyhkpwOvPCndueo/ptyUtWoa0hqDz
aeuqWOtnOWtYTNP3tvsXR68XZmgaduwafACgwvBgilHlcP+0x+pxPcL4wEH7
a0rNYZvlUJyV6hAUDJvobXFiHyX//fE0WhAW1+KI+e4f5OCIYIH6fi6YU4w0
PztFpWvtXzrdWLDpIdrhb3ULY3wvc9YBgNKJUXULqOZvC5zSg1n1vx8ifUQs
QrkP6jC9G0/FJP/v2HoMZp38nv7mEA4o9IN3s5Ouww64nRyWxTNRadJC4VNt
q3/SJxQ/uzyCcOkTdFjYO8YgzPbW4h0cTotr827JQYFtFzzKr9NSfsBbLq3U
uTrpB3L8tEflxgVIVxd04SLvYFNLYFtNpPmFIzCiy+O4wQGhkC88lgPqBVlc
vVNqypMLe9pyxH6hQkj5eJbNBmj22YaeKjL44BtM7XlMsyT3TZYoICFmUmVE
kSa3shXlzJTUXSWYe4QA+fJbmnIXjozQMoIGglPRlkFcTHNprF98/5Ab88Ei
SrfOfnFmBVwxfqs71i3tteV6NoDiU48GQd0DD5QbquoJ5uwh474WwMCr5Sx1
yxyVxzLdv/+mcGEIX89I1fNH7ECqYse51fioNkh9E1kGCG7HW9H8DS2dTbgZ
INM7n4ZjjsmP0YxI7WbMVayZcOaJuRtrhrz3jWtXm7HoF+p4+cZ6dDLHYYv+
JkC3AW8QG4VyFf9c4aZT/rKKBA90ZE9e6I0QywPp3QUWS3HbRcb0gz+SrR+c
qNzZxrt5aMrJ3rD/9AuCtOo9Tm8EeVwjqu//7/wndz/2bztrFJi0JY1d0ds1
dwXrdo4opYQFSXQLSFxJ2s4qxS3urti18YziBe/tat5I70mlYsRbiOGAMCIc
m8pAtfVBkj5OO2aAMmi0ims3I4rqIK4rOru9uxLdNtsIJY1402ShJPGv2Sif
5QI3W3pB4jjSfMTBG4kKH8cG91bVUo/STVCg7jdfFj9fooPL6ifzKESmM0Yz
8OrNKrtSMfEbq974NmHeeg5pIGmPeiwWLtdTb4nhbYrzFbK9VDzKsSLb8CuK
RkxRxD2b6hdGj8zZ5zgqUe4a5Tk/MkfwiK1nmNfMOM1bqPQkpoVj7UfXej1a
URUfSMGEJPZwSKKngtvIE0vkSBXJQjnz5CH1ZJEyqHfmkS3q3BycThF4vUKI
w7/+rNbd84rSq6Eex5SHAPT2ZluGAUw6DDnVum1nkcH+eMZYm1XQOJ/09VFo
oRCUDpD3WGUyBQgFgkLNM3f2ecAZfaEc8IYZLElA9SC4Y638ReQJXXt/N0y8
E0zGylgu7t+QEsL6zNLZhUKPd3k3+CrZ7sKZfCmF29S6hiNCGhw5aJ8jrZCz
W7HCQ0px5B5C6sIamKLZVCjAuIG7MRKAVrfwuKIewLflV8c2c5Sv8eOQ/q0O
W7q5vZClg0B3+KPTfMCjH39v2ek2FLGaHj1ZfTPjYS/fatJGGZjC7yVJXFn1
wBACtgg/I6JhEI/iYbkEqQfndnZcaUAlVYBIRQfh6hs4Njrsevn8EjXsZdtX
di78jXnlV8RGDd6gky9gj8fs+c7LKUz+x4Fx+1/jTNetZJNlrlOIlZFOwGJj
UVgGxgtr1BUtEtLSOIrXiXTD3L4KPIEypqC0OhpLnZL0hStuCftSZK0Esgtj
OIsz7Iyc6mFjTY1lXUJgXQHeKU1+QNkAty7OllAzH6jCC+iRSFChByQkLEAa
IgGc8jH0w91PclysFhr724+snst4V5CjTS64PQqT4rs3Zv6RpfTHXKTx7FhS
SQfSNVhPKll5q+52crcis4ZaKIVvmpfpiQzAC9fdgAOM47jh+7QP7Vs85Spj
gM2gd7dusL06CE0Bnd9gkxfyyIXJSpRAPgiT/jIm4NlK8GsGO7Kew2pY4AQz
u0929typZ9D1p05qMn41RZxdPLjAbyzVQWld2r/WvrBFQpH6rMkX3GjnqhI0
q7SA9/Z+ET2Kl/mkANWurj6nO9KI1X5HIH/VnVUgpnLa0/5tp/d7aUSm+CyY
ReYQHqHSBaf3BlPqw9xGM7yteEW6L8ovPa+mE9dC6xnVwP9v4XjapvKukPdi
hWabmM4+4fGc3ZiA/sPd0Z/XLQgiEKEAC1FNaxDin+zkOBETnEPH0atev6IJ
yzaWXMA9lwiv6ehimHkmfUXl4lRvHsXLWlBhVSOf/Yo4VWOsS5ssbpLcTgmz
lrnV9FVbim+jaKFAH7N0CCjQB2sn22MaYYpdr4+VVWCzG5dUvyqTUOQV42kR
XgYGS8N4i0Ywrf/GG9QcID8Nb75P9I/nE/ML6uP9YNgPCv35xnKwIERi1RH3
xiJa5ucN1OOhp9jfC10+rZw54Z0Ey9HaNTB2TpF4y4j1D91gf8AK5cz/O3h1
vkpAa4tC0DKbYxW7PJmWdcdMoGPh4UuE3vjTYlmeZ1DpP/xBzovu+YAS42HV
OWztbtnUtU+BU0klt72ql/HM11DHoPNUhE+BKqpVqzfuTkMTU4E7tp+qdc0g
0qL1fF2WOtPIYXzbS3mOAhwBz+Mz5StMt8ULvF1ayzjOW+aCIRZOh8JxAJce
24lKn8p3tG+gmzNP2z835SAypJs/xgpNtCHDj2m0kN7a8l3/tnlxPzMkj/wM
lMmljm5RfoFhaKfn5lg4S15w+KsuPBHSGGIhm82OobB7BOYTnSZ8Z8tnP8nN
XZTYHx62zXEiqgz8E+e9LKlIr5kX0sj1NHiUgSLiPxoJO6L7pAskQBCAopRo
4tsm230Rs6EAnqrssynoFjMLePwDHMRWUk/ywJQ6stIAahlNLhDZaEZO8jpV
t/kVyg5oCykH+yWmLeHsEXFXKXbP9c5k4Fis/juwTy1Ki67R2XXrHuwPBeNE
82L3zX1WFK8FELWjz5sbBw/7fQ4K83Ei5f2TFc1iur0kP883hb7xhJlLmuyo
w6h6Ynwc1gPsf0xYbz1E8jIz7V9EkbvVOqx0g+c6J6OiEx6qBrgHx1ftCv+4
Fb9ClFPgfEWNIH+19+tgL07phKZPODQVIoC/u1ZV9JSDPHo5hi0gN0sgWRLl
LPck7tgZZVrPU4aPJA11pkwDXsvpQZwnziN+enWgibmqiEFFeZ2MfjnjTM48
9nakZc3SxMfraKuA+FqtOZ+MUOwbO251W/AV3+AzfcuaMeEcmUOMG607d7sZ
DvpYJTCKJFoyXHjny7Yp9erp+13abAv0WZd/iVh074oCYt1OgXPHNvp5u1dh
C80qNNnH5HEmLSCyoS+C1X8CIEH4XVeF+KK5Z1PdBROLXdcEyzFDB8so/ChM
W55/haT3N3OAPeFwBM/Nsx+ZfT684XGrjgn5AcYR7Ns0SaiSIARmHn5m6d44
5Dewofa7HPaLW38IS7+GV2te0/jdSg59GEnGVrXxlvqoe72REY39xxCo6eIf
qTYMeVGZXS6Q/BDRRKsXH3zXGu2fBR57Te0xp0LflyRNGKUMgSpFMxtMWFS5
3KHLE2uZp6zaCerwkPdgvNyID24b33Ho8Ydu6rkXaTFaAQR6LJ0c+pKhnHJd
0KRe9bgNc6/LQj5j7Jl4AJuzq0o8UiIostonEDfQQWh+5k1eCcQLRYDfxm/0
hAOlEOTbgLgKq5qCjtIhRNPYIUmEfukQpr/2HvyAK+TNqgbG9G7IpH+BCihK
uTpVRVchiPA7tJvUwuVQqLdR0zjIQsNRPRjVxl8zLqXnyz86KtMik/gJjmie
KeZCQlUH7NfOgDDIpSUqZPuEllcI3cvjv2rHAcxN2xAVqQgOjHKxDSh1nvBk
0DJG8SZnMsqB+IvcPzi3QJXPycmrsXA4naXBJUUJLL1kGUn6f0ngN+N1P8fP
VPXgPsX/e61g+ScxHwwvMyA167/C/RmvLvqUDQTzt0EdEmYw0ElNRLif/FYT
kaylLZ5roq++b2kKpjf4W/T+rlvdoFhCnEncuwYY0ErNb+LTvIr6O00MhF/G
n/9HPlh91AN6q6mFTUw3x0shjCv10qVFo3kbwf9jiCTrqd7Wl8jKAi+pMufh
zaWzoWVkM5Dtaj5nsb0E0L02+S5QMc+LOsp9KtUjNvEjnH94hW8FyzBD9+yr
4RHBnRYue2W/2IFXvY/ou3tslLQY6n/NzUbKZ6dS40rz3LqbqNiESLFpopdM
kYwIjNhwcAIsqSTJwWNTiX4ohR8wLyGQYkRU51a2RdRky8EXqlCKSaL/8R4O
NeXJ0hZ4b8RDvLsHtRMga/hx6PqIycj/3OAfnlkuynZo+T6wu2T6dmY3ei9b
hzStAeLd5nPeoNFEoDcJTXxQ3QlCMp0KRfdnOb2Un1aW6L7DAXb+5GQ7bx9b
kZu8t9cNXuXc18e8UBLDqJhU3YumrrUmgESlJVPQoO0IuMphf4WxNDr6vtob
/cjYRxoOkiZQDol3qMcANnIn5GPcTI9IOnqQXEJCI8zWALgjxXpRxQQGAr3A
KuBRsNAHkCEnDhu+ijZkLj5YowtBywU3sy7KTIUnczihrSbBLR/jxHsWFOwT
N0NLztRrqLF9ZlV6yJQSsXgWE34unmoIKX3k6Vw9VA1hOSVu9VtadljGZ/gM
Oo9AGq6d0qtl0r3jpZ7aXsuODrngM26tHclbO4IDaCfazKmM9JFY/eh8M8wc
Oe7BpnrJQ1vKSP3Iu99h3stBRgm9uaNhlox3RUVVYI5pI7o8qJip3yHvh03o
gB64AA3k4HTjMDyzF/X3cFamazFF9EOMGav7sFnWSh069SdeEnVLRqd8XdyF
PSDoee+pf/NX/PPJnGlxlaxekostxYx9CWVN3JBUVe1rvobChBFEPt9pQez8
PqZ6YBxStwaWgmT7LT7sZHc4mnnl5BeUJONKv0akmbckPecSSDiQkbrznq4w
BiZz+vfllfkI5KpVvO7idXq1uHpqDkhCEZmToPP7ZTqv5G3AZ40ax3R5x+8M
rQI4oHMgj33QJhewKF8CBm1jhUIHQOLBcl2jAPnN8d4GcColeYvPFk2bHqvQ
+AtpHDeoju9r6BeEoc/BrRpk0C+Mqo3Z0MLB4pNaeHgBr7AmDpS2UpxbawNB
is5cLOUSrZ/3CDxslal2M0XaL8s0qQQObmcqJwynE8qFCPFGKOVugwiP4M0R
YtdeCR8gLm5vpJH7+32r4n2Gc7VA2GbE0hIBsern0CkRQscKElhyuVD/gh+b
Sf2LwUPUS/7vbFPL7nwfWu6QUGrdL5E1EihD2dtSec1wLylZtj9r6OF6qc2w
Hb38vKZKisFVjXJLjtlVrRwGtNFRr7cvqlvaqRcp8dFfp8dj+EM+ZM7cXs6/
tmgssQLiv2ZYyFrK/unGojQtScdV63SiZpdKsb4c3mGBeSWWdoKGEcI3w0gL
abo0QDFtPqe0qAnITb+VJj1SUBp7G0026PVRqihXj5fNTnKSJFHFcJnzosV2
jNPDX428Cre8o3pRn3MW+a/+UmdnmkQgU/iS9Qdx6EoIuQ5SV80uY0pUHtQI
Gnkkt0TNozi6V3XIh07ZwmQQvgzbFcmRBUvfCwC3m1PYQyYHtUU340TANr/c
a/uRU3eZE20LCddnHoJRn1FM/1jXeSuv8DfHpRPlAugimDgqBhEsbKJ/kKGE
HbUVfxJ9XRwC+LIxHgeDra4+UtenY0yd1NCx/+KQFF9l16nYWVECRqPnHGml
vQhVoGS+YYag5knAXluFNc8ISxO6nVLdKGMEsdKmvBoe8/manJJ8WHrKKAHE
l7Fmv0gSwaPgOCrBjUCr222rsYKKh6rUidFBCfeWFTcKyUjeyPzeQq+il/ko
0rSgiVYQ04NsSRh3XYltDyxVo4HiRfZRyE7+TESjXGiNWuqm+PBlO7FaD5mF
TM/njzhFRxX2GEcIcp6TJG4usX1IKN3NHErHAInMsnkN3QK1paFoS1/R+FOf
jZJdf1txiNTP6da2gPwlJ5k/rFTz6SjNlkCVHeBmGp38r2AMG2KNGgn5gwhB
zhK+dJpJl9GQ/xOj6+c4VdGwfv1WlFiabgLvCSefQMIVmMBL1OKrnkR/J3oV
QJvnyBKlS2td0+niCD2CA7XHeOpsb6Kg/XWpiWK7g8PV4sprv+IRcedkDfNM
JMbMbO8NzVXs77KVn6OBPr9kezrlZdgG280r2Yio5L6USf3ptw5Feou1xAU9
CKzf1X8on1+HLmd7PScf5nCSy8t/Bk/jIs/yWSXj8snDVeZgA3PieOiAv1z7
Eq2YDALDSMdSzxuiwXaUNnUUaL3HVeAsx1jSl/s6/ezOPtwqABlnyvvd7xue
WiHWZ3dDBoIIdOZLr+3fXe7zH/+MMLrv4qMprC128ZzRRSsfG5WzNKt3K7TS
XXxBZA+xiMg4px+Apuj1dCfjrOT9mxv25gHJ3qumQy1W/38U49DJx/UJW9Ew
4KqmeUf7EeW/dYgZH+kh2LsujH/vlZvCIBNYoocOnTQAtjCjGzhj1CtL27OZ
nWuc3BgB8roW6zBZS5v+KPwMwawiKoTdNHwyzx4I4de09y12oLM3+FOvtHle
rLX9kdy4R/KAhK6icErDcsF7VkVAqCy+r/1Yp2Yulk2/C5zXu+39xZUtp+OT
VTGR/DnNlB0puMlBEc1aA+CYUXrxas5j1ekGeAerJuQ19QPJImUqUS2R3V5Y
5HuSviXAyle1IFOXTGv/pDrZw5vfWBwTly1vwNsJ7TeaRnKzOFIp9tOd5Kou
Tcso8bQGcDfh2tWKmxDHdM79WeFISb6Sukc/xdh3d76ayvxIT8aP9B4eFFcA
NyJ/YUzjSVHtMXnEZZyZ74YYqBym+5IP+GF57s3Z/CjECtGQBiiOjYEpNuj7
jvpeqH76b68O4nAR8LDM7LVFDchMlaiufvD0rp5UgKW9MaRM8/3a5G3U31Ig
uNgbA13/nXI31xD5cnBLo8WBrlF+dql+A8yug6X6pYp1x4+6mAZUNAbovavZ
GM4ANCsJH1MaEhpWpia5PRLnsvsR1HayZPXvEOryMevB7IVroOkaihMeGl6M
VaaM0r55Sgd/fU/P7dPcRJ3thhKvyBnIhsL3d8hUbfNKKjEgwZ8aihnD88lR
h40UCxStheYEWsq3EokxFZurr/8c6NDHvtPB1SDYR78wW4n9ao1WzBFzM3Yv
u59+6feOv9B4blG0BdM8e39KMb6aI1SecLCfy5qYZzzPYGQ3B6au3fiAuatC
137La9ozU8OCuMp/SHMKVLS+D5Sw0C6PVOAPq2IBO8PEI0Owdnadtboskti7
sBbNWyre47TG2u5quZQBk0UlK5KB+GBAFlDOpjlLvQ0hsSs0h8jmRbKIr5N4
DwB7Mmgfq9i1Azh8+NACCbrQoBf9cgktM+3DzLM/ivHw8vUKsyR2s1XGB6TI
Sp1usMW05uzMXSl4pwgTunDbTGxpHtT0ySGsoANyVGvmXF6CkLLF8NG4yN9c
BIppQzjSGvkttwQg0S7lwIbhTgBFRqX8CR9cGEo5M+KRkK5CeRtJ50iuPppS
3I7Y6ssO3Uj7In0w+ljK33U9ILzgW3nZH2OjlO5t0zWo7JhUYQCuwMLvWrcS
f1JsgQvnGRhruOrV0WJ6Wfla5Xnz2MHlzy0rNJro8LboyqDBMNeKDpLnPogw
MEzctedE6bxyvfdnxAmELng9Gk/JHbsOiObzHBGEccTf0Zn+ZddQSakMwXlI
y2YK5ey9DFHvuUQaPPJLBQIIZK6MvhokKurRS47bQ2fJU9eQ49LvEsX+4YkO
4pf1i8zVN+ntA2BA754JJjRxoUfo4uLBX+A0E4brTSQSH4qAQSrVYB9ISVQ8
OnbsPbONU9lBOuf7YiPH+eyMqnX4SYeZc3uG9/5q8+xv4jsVIdgvTXGGk6Cp
y7w9Abe4/xh2wvxNSA9B6Ucz48Q724uy2BhwFZypj43l1VHyQYs7X6IOmUAB
ymDPMyQOmIYbkHUEGTC4LBMsEIwsU/S4/anTRshK3Zs1XWqPkG2YTfRVW5GQ
liu+ucB1KvcZZmJcdV2uEzBhvAqPWITF+Aj2bcDhFlbFqMo3w3jEkT7PtlrG
hT/IRDVd7GpeXd8ZO2bHAke+bNu+RY+9G21nCJd9TMjB5uvLZyuPV7zSBoWO
5X+WalGu4Mdlcf2zs7bY5PLYdBcQRkrOBmihObfPMeF0155YoN9swjId0ZNz
ToLB/n4AJaQHgpDJj5GZN85KA2YsdbUTTP2lFR1b4mtVUiDXnoaxMa/ViiH2
KQ951EdTSBJBmQU+HHmj4ySYeLOpK2BxldvjqEWaHRObp07OZzkBVXc7tHci
/IRYBuMyWuh3+yEO0Vhpf1J7ZsfXnoHlr1jTw+06wGoQLt7i5Bpgaks0wVY1
4Yi0TnaxnstJUqn9ttZAD+gR4sqY39z4WsMuSN1Qw37Y7OisabmOTYs5ln4W
4NVjDuX3NHhBZfFkxH0LqzKdGwxA50C1FuOwwKd5nCUpgCc0rBLKKgAcQBTt
J8LYKh9vBX0dGf78DAZYISkysDPXJx105t1WejHaigbU84paPEri9s7niWAa
BjS/Q6yj8ESE8JoJmJYskmSWJPHbHY5wzJy6MqMuroZHYTaS7y+jS/jfUDeB
Tg3u2idInRU0MG0jhM3AgBbjLOxumk5bHnfbGuhwhZ7TSdHVFc3NSywBW3U1
A4jPuHWPTK/aRw0pAcStm5/E+vSzI4jiISlXvmFZ3czqYOr1j6+krPCoOB4x
lnmScRDkO69HVU381a3IElYAbOYhj4vBorGlq9lpqfnU+rXmONTBpnrpRZOi
Qp1rEpbUTnrXO33PJ/L9kBCveqPDD0OiEF8eYwY0Hv1Lukmj2vq7KNqHCqVu
A2lf9tilmg83wGBEC5myLVPX1GvaB2J4R2EU3qhN+0QBS9qYqqRSbR/x7j23
0SPgmAb5/Is71CvHiXDTi6hAC2wjgw2tiK6SPDiq+e27JTly25Z3E8q4BI6A
vpKPoBFb9tmiSO84j/XXl/OhhKDVArzw8+NwXdJTKBdg6dNnXBWjTshqmCAi
cXJ1OkNlPLtL5S8GX63GFAzQLnqFWi2DwO8N3uZpjOC06UxDhcdhoibxOht8
GlK+jm20QWW7QalFW0aaq30XGfxXuJSw4O2QuifqhqFFkMfTw+H4Ap2OwTOr
fQ2x8MfInag+fy4X10EzCfv8d4puVFphMCM8SbaS46JDErfO9rMAkyxTz+ws
UA4w6yPY3beHdE9NE4aP5ni+qypp4gPYBZ5Iz+e7PWlnlCJzbIeDvPop7iWp
zqOUvFzaSCbtnGRH6z+pdQM8PIhx1cavLE1hxV1MfQUta8DfdxYdj+s2g5WM
UHOAfPwLgx2QXvpeDt58SAi5jc/EN4qmFb72tSB0PXyC/GGlVUn4ZOAUu2iv
4XTHSM5OJ3K+dpZvlR6DMPbKZOH3eniivAfUxOdx9nGL3SppoSReeUhMIGvp
IU8DRb7Upkn4XlK9zraxHbdSqc98XJDSXYRL/9Yv1EDcBbwPBHPimci7g0IS
lAefXxcUgL5mOp1F5TxAODk/NwF8DBHU7CrDHO6U5N87lLD93Iry1rzSpB+J
lcJ+VEloEzvGyklw9nNcevyVDdevOsHvdzt0ipkS9/OIe3LKTop8dJJ858ks
CzYk3MWubQ4x3b8gq08u1fAyH7bSflWFkC7Y2nvdk82ClMA5QYn6Xf829GRT
udtkqyDdUZAnSR2NHKUdaHO0uxm1aiDrkhvWUiW9c4x/GjTjmHV1WTl7iIQQ
fKE35uN6Zf7MSEQ6ln4A7dz7MEfLawQ+Za2g2ZEZFDRCjotYKPCEsDRP0Y5N
2bc8B+i+apiIddXTV9sX/mwEYVWJJ8npRvuIUOuE7YqPqBnqPGOwwvQkXzKy
dWp18Z5OVhfS4fW+N8dv5aSnxkP1H6aF4gUUdwMjl27FLZ6do6fEweXah5cY
wGzXByQlVjhAcHLldXnhkshFEjiBsIRr8BGgAc8HgohEtGoxY3J0Te6s+LJ9
FhRNwrnAG4tgn7xk2mZZGZE/SNviPCSFEhFYVPQmiAyqp/MTtKvKMAD/BTss
N6mlWUg8/FsY1UJWXv5avuI7v087zGqqXRY8ady/11FDi2qYtuAGAkkrCaW6
z8UAzbZIiQkTJnaVftIWEIKQvHCkFt6mwZpbJDQWtc1/LBd8nyjzE0TMbHqY
07i7SFWXqX5+KC5n2g7SdEOKqoYyE077vzb5BWaaO9cvUF9AzlOCppAgwRL/
XWPD4psLOQKMIHIxCubi9adGYaAdXiLVCzH1ttKSDmpP2/HdnezOZJ0bPBvF
ZUCMdkWBKi37IRC6dy7ZYZMxiXKkLexh3rFBigHGMTjF6Ug2GCFM8ErMqUTs
9Z0zYP2tB+xgs+yH8JKr9zaoKiUELs8VPJdRe/iK6ERQ36W6CCZrLJJ6HQ6Z
Zo8i5zuh6u0bPNmZlPujcRk3jvsy2em0mwbUU9qCvEqWJjsTDqyJGPLdEmG8
kbbYYcZB+rNKYmwGS0qcQI3+dnKMoSjik9h21yJA+s4qV8he6IXxKvowmp65
VrNW6xZuPkv66CFlCyDNGry2VLxTQ9r7WxqZjURa67X6Zffh6o1qc3pndS3J
6CO0OWslf/L00QTNjBRaiob2nFO4Yr21N+XoSMqWmDAwD6JInNpp5tVci6XU
B2xFulZGwzeuPS9qUGR71faDKh2M/xLKEhvzXUpZEysE2AyR3QR3xy9Y0LbY
0K4r1+xBFS83bNV0MEDOvDRvJdxVTY/XMJDhRCrIsVCChN3H7HyvAp+a7sof
1ErjbSDL4WywUkzpaiyhi+cYUBWbIYto7vgi5a/cZZg7PwdTRF8m0Tetpw0c
OuWzq3kXBqKL082YET6zvzHfgpd8N+FzeYea/c+7Ugpx7lM8FmJXNC/lyBAE
2BlBvRme7harCJJMNNbBGGc4w0wzxsCNQRE/RTuhGH8eX0OFeMwNgVt2T1vd
SyYRBdY0i3AXPq2WMX9e15e7dnByP0RA1vUEK9SI0DOKuCj8GahmwWAkvqfV
PPSj4i0pJ5xHFoDIFNZwkSEsIyjZpHmecR4nSzMIlxv6mYWsy1O7gYxBxPsh
auEbPkE0jAlXGBFRdbaymQuyhgK7Bc8ch834FYc5w0TcZLtaSap5sFDcmrXu
NR4YTowzAFBvpyMk12SXZ+pXfdgs4LwmbWZ5X7jMWJIuUdM8YNBOPAW3SUcN
/jt8ww0sBcx3o8gL0BrEoyQpXjHcoYfMORJxX2h1bexB8/obKTUKHnIkP0JK
MnOq6XlZkFbqPqKvdQJcZ49MjGHZMrTBXROeHo9evGEQk96aaO7BbNHRbohH
W10tS2cyHYfcg7/OBm/rlTh9VkwlL1wivavlV+eAvC5nXJXOA8lHflr/26+J
agTnp04r5/yPKz5RDAPYZ8C4PjFDhAeXxzaApsgldCRxoyN3UYPgdoRddOJl
b3WTajWH0ye78v73tcTXTtDAfJKhLZgEpuu9t02HnygpSPmgJDqBnbekwqa9
H/SDOGipFi8bFw4bP4PfILCBvFrlSWBeJ5e95CAw/Zcyx/p6+8+JTCcJrAQ0
YlFDulQDimryYAuW/p5SHpNLt1TvnZlNyu3jOZ/0u4cgrHquTF5t59srs7qM
UkCh9UiIWR6rfZ0LxE5Nc77m7BB/+WmXoFFSxlYU3YlyIAuEQqqToeBXwLXq
zWS8pCSOyhqwP2j17JOOTEYivV5vfEl2+r5jf/ytibBDC2RqOZeyXxz3SfRh
7/sX63ToUga1RKAcPA0vL/ypY3dZeBXOLudlj8imfPVYCepeWoUau2Bnj74U
aVUIC+/jyt7QhDgqGviDpmflP6TnbfCXSy1pSymCVo5nD6WlQmP6kuS96lQX
6n0bXkwjLq6DKg+nV63pnaVcLPOA/Yj05XcLiamCQ0OoIOfE0cQ749TmKwCH
/xCt76Gt1c6Ruc6DzG1VBlP6XLhI41Zg16Dm1LTI2jdA1OImM+BV0EItMazP
mfOdy4Qkm36uH9Duoln/0Z250GqplHKUa+sN9IVkU2Pq1fpRak6wB875MDKO
ksrJZrTg925IYF3otr3M1IAyquuzPcx6rHXKQo1H1Uw4kLVdOBzbNktZlaHv
kVEolfeBdowUpDXjU9XD1FI9dQ7sOaNyXTDOshHBFuZXthw+wSR8kGR+FJFc
ApE5x9opRvqQisxIUhCU4Tqc7TIdn0T3sbZYaP3oQYJ13cff7rGHeJeP8dn3
/51cGLJqbUJbknhg433ho8P6wFhqy3OAZZw74bqxxuj3sQaWb6/+MZZyqugN
zVBAx5nXXXB4Z9+g6SkxvGB8YTjgYY2AvPVmTebQ4CFpDT1vWWUVhlf8OQLw
7C91GZxogb/VJGlPEVNYT00NaXaY2LEkORPLxGsY0Atq88vdZx1ykF2vv6zl
/9PhUR1Z92Au41tYr92OevNBtSr/SQpcxHjA2XqOR7KxB578eRb6aZTLgRsl
SvU58my3ngg5D/aqINDKkdMzbWm6wNEmK55zlBU+zL4E9AoxiOWxqNQIZG+l
GpEd42EPfM694AHGIWtEdQU6DEB3n21F6BqUVKj3VD9wroZKKZGgunlKhJsB
ys5X2lyAcAgHhnZGc7zxGKvxdrkY9WKNYsCHCZpzFlTsCqLXbIMdfITwHIIL
KJUUWWj4J9NviIb1yYxU3EJdYZp9WbL31cstBsgm+5VC7jY90aukR/6b3LAD
gnzRBxpXKf/Zsrgw7mdl4sDEwpQPP1Gcw1vVpDdePHDjoc8a33cdpgscn4sO
Pz2XeovTsjHYNucN1AFD/55/aApHg8MSRtv0e+2cQw8iXAIh5+Dl7X1hxRA0
tT6jUHkax2Ckm2iMkssD9sd1tcJt+rnjQ0zCS2VGHZfkBnPEFXQH3oh/JF5a
3j0EHs9i3tAafXK0eW+6AYuKV9ok06ec7EDwxQ7LjFwVPgsZCgSwo9jFwkF8
Z1VMwfDADUSEw064MHSbFcu+KgFS4UTL4GATsSDzBb31uk8kTjRGl3SHUb8h
GSnuZAeZy7PPfe6TTmvDJIjr03z3Q4lGXoz+K0f7Dtax9Xtxv42VufOoLLG1
/U4kDZfvm1jzGN7/meLeysPW32n/xgEgloq9qFidDHk+7GVMUQL8qvFCU7eH
6M8esRH0L5ptYXnhckhsStK9JY6j3rK6inemCl2VwpuhF+noAsBsCzkyF0pQ
Xw3XieVhomtGzu+51VoKcshbA5ebGYASCxolWWHsf79CTtYb4DW1ztJQ7aSU
Dky4+0TYSj7H48Xlc/jkoq9dDdma20YiujS7fqvQHp2+L4zHTalYNsTyW+Qe
9oq+UkEY3Uy5Aw7/tpmx7QNRKPOnrKnqvZg/1H3k9XlwOZ/VKSh89xoEV5af
Er4dkL10I57TKpzHhs2S15+5/0+uiGbmazG5fgDMhl81O/tuF6F7CHXzm3yy
YKVelrhZlFFuPSKRjGbzung+i156mC2DSuvMv3fm+B1c49Ro6vy9OLp3Dl63
3+B/XRkpegskSxF2t6xVPTKCJKkoktwia3eDB9i/KHdo3up4gWUUROhmb3EG
gsMouHMULEsjIO8lZ0bSye7RMGziVcqSmsGQ4bfJJNHrUa2h32kmST9TZD2W
MNy2q0RfH4HL5VZVAnTWiJduTiceHG4ImGhrwmHPhw1c5I3IVI6GbitEypzQ
m7MrbWysNVeMmp60Az8GUQ7xOp9QHko0Qb2ArUdQ4KBPHosUD9B7+hqCk7gp
zN7dkJH38irUEBSfpQrkm+uuOOFNpirhegyLgiEosTsoc4rQem1npk2ldGA4
PxPNGBSQk3uNKdXZ1hvDfbq1gAYNHnInew26iGlmsgfBCvRf5ZuxJY+45GSE
vK+af/U8c7EDxo3zY8DQwFj2s5Vtd2bRzd453EmEvzg2N//RjjybDo+PwQuU
9B3JZnF9+t7OYYJqZmQMlQqWiz3S0mRGINq/IFSfJNg8cjUT7j8vxlh6+Eah
SFxeuwX996X+VEVQ4LvLnFeRwEmhXmjMHzAVA9ZwKBLiEqWdy2UJ/RmsgoZ6
XiWlLDCRZkIr+a6Nzdcn2gLvcsbZOtGyuwFxbmS0Z8oAMBIr+NyVwswEp2pa
nWavv6UXUze4W58Xxv1F40aSXs4flchJ7XhS5wU7Y8mSL6Nd7oHR/TY3kMjs
6GOzydD55hzmAwKJISgxVdlAPtuU3Uhya+1wkyj3fnFTiQtB7rKZ0re01JtG
at91l9CnMDnjgManCNTewwCMiVFQnRx9krxidw2E/ii4xbjQBHR3P6N+5Ihl
Bnl68grOAZymnYl4pfaPF3iss1svlVcDxaqwEMfuEwx9wMX6BfLb4f5XSBzG
qq0KaaNsNMauJ8aTrBgA/mBJWVyABt3WUwx0lUVQFRnpmWMf/+QXPUnYDld2
Dy/x6jMKZRpYiAlfBLsoT2teSsUSbEgSheNvgUsSxD2sGqRkgWtq7pw8aKJo
m7ysNadI8EDsi4X2N0BIVQGjwQMUQGr0QIv82vAeNR2FPc7Mm+BtDJmGOa4I
O94wYYuyxFqDCPdUT1vQ8EZEi8c3SBPLvOUmRE5xySDDqGAVRzowopumcMIc
tlHYu3buEf5IrT0Rh3u1ekRdEWobnzUWt/t47SGq1yImcqQsCflmwMw2vMH3
5NNhNtsHMqABzHpQJKemS2S5mWyczw9xeJ074p4HddzxEqansKWf4hVPA+hD
Ead11rt/NabHoAyFA9I3nCZztHmZhLg1QKGWPonSy9V1uLYBgJHJ6b0JymYD
iKo9qa0ZrOjD7y9RtrvpRFcd9kTjYxSEtvwbkqUzgJS6ek6wSDcOd1cLPvI6
9uAAySZliAywIPaSvwtHrjW7P30KY/bWnXDWnMpvALVQYPvC9lYzWJB5/qLz
LRX6vK6PffGqJ5Acn7eJQzXltbB8CJMrxcbNqRo128RF9E34B2uUyrt1bhNq
FLChIf8l6MbBgBmrbd6pRH86DlnYsrS3yj/n+BWcRqS+guXl3awFZ8jONyik
KopYrhPmBFHLJTDs2uK86TEpf4yGW7T3XZXOMcfv/EhMIZr3tCDxQB9GVadh
FyE83JerL54r+wUNekDBN04W2SXIaKxle1stegJwuMMvKNTkYweBOF5vUjke
AHPnKkMNGg2UYffbBmWigXV8D9WAcyWuT6t2up9a6deAOVxkkEHlt32FCdSn
fnsF6P0PqKHMkOMQG9IFy39Xnm/gO0QzABhgkq2L1DyXwdblS2Yrk7U1a9qz
PaSW7BvWKU9pM7yFVqlupjZ94ZN0rZUYx/cvpGlesHXgHilRFKBmy2OkHl7F
ZZ4bOtqMNBESVnhLotb2Oyhtx1fYbeMIEInLaX4KzghLj3rRlp/LUfYdvDu3
tPMGhC/wM55n6OTOQRnuQ2QdAJH13+ls9eP1fYSSh2PUtGbUpib8L2wG044r
joj9raqCl/2c0CflxT0n0cGsmnkIq2XfFrkHWME+yzXOQIJKfYCOdYg3rQb0
7iivMItV6iezJymOUcH+5p1+7/9ERlekPBJY5SovOnjZX8Fz3TybvneMnNnU
g2Q+pYmgWjg/RzxPSOSVb987Or+sOT+2wlyxBnjvPDNm/WjXkfsItZIwZjff
as5+61fGtYPJ2sLbSN1Qqy6I9fci871nk+qap0NNSJkzMTilhaIIuE3YctcP
k8Eud2JsbJT1sEmLZ2qvLCOgBQJKkLgXdf5xbCkLnjL2knZ3j0ebgsK2bZhC
LQnVzNQUe0RXmO7MmFz5VgWqyfJRW2QbVCUU4W0d3zXRnqU/0qtKi8lReeva
0JoRjDP6Af8hT8DDH+bVmP+TwkJVR5w1BgcFK/NZlZ7oD6pe0vb/YnmJPSwg
BzjpsRBORwXBDb79Bz007H58YfVPya82Sr6VKzWo3L7Z96drdaBY1LeFmCpe
q4liJHKnfD3yyJ2k2lf+W1Oa3PKyT9sKh2JOSj8QG11Fvwn4tmrmojnvvTgx
F7C1weapkr3Sfdu06Fv/lwJbI74orNfCPZgAknf8OTRqHYNS1TPHqH4lgOdC
CxLsa4nzl1xgNCUf59LCoUDy4RMMXmg1Fm0261YH6cjHYe2eN0eUhsTNB2x4
EbA1mKVtf8uJT1uKQimPf9Lp5Eot3f+/3E9Jp6pTvjfh9v44oSaQ8PwymZeX
cx4rPE6fG9oCAp4X3ER5pu4lUBThXD+j2vNJKcT9gxfpXVtxJsJZFda3Cdri
cml1PUKY7Y0eb+X+rE4UfQ0fH/SqDASRpWNRnDGz4Sp9h9Z61ok3hTmdGJ5U
UFeBJ2O9aNjn7PTEAydBxmXEO0Xp3iYGcWngC3X9QM0rA/4R46sjVHebobP5
4cJ6e91Uas7CkfbVFKX8Qp/4G/S/vvN8diIE6eTJPmNmudnC6QyBI/2LyljA
ieEVUp1eeq4YsJvKb3lEhMRVG7olzTp9zUa2seVQaxAlfdw+Tt+McBrXwW3V
0jVlFr9q3FC5sR0nvkVIRWpBJpHmwEGMCH8uX2aGEDfYmY9uMRhAQ5sSJzWz
h0lEQvTDFwAhSJcfTCWDoTErrYN25drUOQ3z4GhWKVn+1reGrqn5K8G8k5RM
k9Vos/JftQV6hhwAKUi0KKdCo1QAjMsfP8LTu5l1rv7ZOa271weSStQVXGA0
XPjcXaBapvKN4Cut/nDFsoLPW7UIeOggxaRl8rvN2m5VihuS9FhiBoBATnhD
22MhA8E0j6FiH1enVhfwF47gQBXuKXOoVtCJhswRTEVkJe+G+IqL3wSBmj4I
pclpy/oyhK/PAsi04UHam3mH0UEHVBGXiMdaCfnPq7yYHEHpjQZ+xaCteC+x
tkNzVVyKI1PrAl3sMnK7vwmrt3llmrEuXLXJj1OFAxtYw6XM3q2OKg9EnsIk
/y9Vs/hUm82fWHyvXBaXaFa+nAU4sDk8zWq8rqrCIhyJmNL0TuFYqLWMPnfj
qrzg2xYGodsuHlPE1nxtNkFBQ6DWuG19oJtF3ByLd6juu2kz4S4bwu93a+fo
zK4K2JZdl3TMYKlNQWpzOhiikNiOErze3zXmA93K0YaallhoS6M9KommKwvA
U5s7roEXTPqWJI90TKMnaBK5NTVVCD6GSyqeZdwkVqAL9hxwWSgvDg4VuGV4
bYA6MItarOl6wnPOcch4DoqpXVQY34r4SyITdoQcNl7QpYZGlS0ti7dJow37
zi1XIBlEWOIBeg0hNorYqEpojEUR0+aAxUTW93y9U6/84Dl26OSUFXKm22XU
TJzRtb/bVFeRuU1qTkLvZqr5f9ggg9sBaMPa9Pw9SJj0ojujzn7aLkj4+x5m
oIyzheGYfAM/pxYh7w1yG6ZlyPxMVroDstJF9iDkzjl2dmGyY2U841S1//Oc
7JdA21e+A1s3rAao9X0n26uo9LMtFR1OHTojzSA1SDXUdkTVIjSCKQoRib8l
yVIiGKwPFsE3g6W4JqRiuhd/f6d7y0Mfw4TZWjPaWdPpgzyLEITf3h462VXh
/k+xT5A5OoheSfsvW70Dth3JYSR7VW8R7C+hdR0cD21wZZSRLUkXGEQCxmO9
JEP+tDCuiDL16kYo3zGr1AAlJWm9dNnEC1lvKTIrq4YreCFnY7phSSEDZXZG
eFRPaM4d8sRrUQRULwgMH3S8ZTBzsmNOZeIS3virirk95IzWtgisvSQ+Nhc5
A2H3NtG06EMqOczp+qknA68tHMPfEjRz/ROCI+MxxlcoWlit0MCIV6tQ2JVV
g3VS34TiZaQ6sK0RWCEjh+TZ2DdCbfQE2F7IMa60LE5F38EHygKvI3837pYw
WsKWQOLQZEuIGZSSogOisp7xNuEVPIT5cG2S8WVQQmaDHx89TI06TgKnreGv
uZCEaNDNWc5uwKJyCtnDQ/iKGVOO783ranOnHfBloreDvAmWkzLRdYQpWYKL
4Rz/jkDS5Ttv1muLJanquYef7um7vQpYIE/iqBRywHV43g0dcOsIj5nV0OhQ
EKlHN6wluj8F5Y36s2V4Sjh07vMY54MDHThd1Jj5trpskWaA8sI6T9QvmJCn
aB/KXbeiHCmQGfxMHAoP0xA2OuNAoqqzZiNjtfks6OF9r3+BXqVVTHkjpL3Q
wJ3cjwTyJx2uy/62BaOZT109ZmJ2sz9kADejimamK70Muudvb/jP1+FvDj1o
mRjq4RYq0gw3neBd5E5djjR/C5RLom4VCrEceJIhwfpfDwf2Xm+ic29w9CAL
gYsXlY6J5mn3z01W+aM018UupjPTK7FacfAJWvcKbw3VHBBSRsqFVQoaDJDc
OKpWPZ1JXOEmTyIkwshfPBgRXnO8L0EiZ97tk8FhgvzQwzfyOaZM2twntYxS
DwEDbmWiUcPlmu0seXtgcOyGtr/BgKyUYak+JKdhqtU7YqhuujYbf3iUlawj
N22Qtqu8wzpKuEoc0AEnMU/FOO1ssOA3djP+zh4ZBTGhDlATSJhBH0a2GY+/
uoxfi3mK0SJj/YfmwWXtxRgK0RW3B2sFK93rIzWTXiqNme9pffxKEWz7CX1N
UdyjziEOTy3BuEcJdcLYNrtr42Qa01wI3tmEESk0HREmeiGOj20Fwt752HqT
TmpTE/cPvYKNvYVtw0dU4xmduU3AomNug3s+2GYm18dyVdmbnbIPSLjgLL4j
LZHY9AdGthaB49LlAZYwyPtcVFeTXkHbDUQSUfFr6WZ0eowKFf97uhvfrNcH
FetBTJASsSxi0yZXcz7D3TRcFKFdVi6USdTioyl1hEse9VkEv/OLydOG+obt
KIR1KoTkMDOwE+kkM8nFXO0oLKiZlvo1XalsjE8+sk5zLDmTgD4VxppvwDRL
kryc2eMGGsuRIZopO/IYlo3jFKh06ASXTyjfS9WJ730tgPSnGmTZ7qtR9Ex7
OY2VxDq9kJGpkl566s3gGDTg2v8gAaSf3+GgOZns3r9g7woEim1N+GG6JVSW
yOlT9ghtYtN6itUIjmH2IhV9N9AH4/uz55f14QLf5SCL3hwFodLmtnfdu1rv
kjI6pxo2oInE6KuleJVYPFTtaUEgv21j97v4q+FZnqiWKwQahhy7EfZWsKSS
xQF0aRkt8H/inVKZyyDRYnav3Rgx9vvFQtdpm57V1Ir0BiqUw130NbSdbOxh
A/Rl8sbKoZpHo9FH9n9JUTJhdd8owGHqYpk3QUl3DOgj7bKAOM8rZDHiMU52
UCpM19XnLXlpB2LLtB34eE/t2dwpYysYS0VwcfZFBSDyfe//qS3rGe2MB5BC
noLOJ4eO0rGxQolmbNCHtjYcTtq8sLDlp4Ldqe2KzkC4mYfI4OzuBhHEjd4A
jfoIrEYTuetQn6p59aZOs3AHZue1gdzR+tfzd5BxHnTR8/w98UHcvpUegmLI
0Ikfb/OPeTZSBZNBnS9mK0wN460liRYK/pqSu3qKdtEoAYO1Xjhus1M6x27B
O4fq7iYbLeQc78Mn+JD1AATbXVXUYvv8n9GNFyDasKYFWFt2ITuR7u2xnk0z
7QVDo7Pu1ndg56mFY5P0l/xmBO5fAphCUUh64BnDi/SwzwufUEQr2H28zAIQ
QJBYg72Xqc5+6CwcuZVfX/ZqIGLBWaqct6YktUdFPIznj8gw6GzgLf0W6PFQ
QWtxQdH4WKtDwwJKAlfgreTS9nfscBSHUMGDA62t7Kv5cH8CxOqVj03TKwX7
okrx2MNvIBn36mlXRskgFnKeqTmZc/EXU2/ltXJQuUh9zOouWw3E0jaCY++H
0zDDWlhGVtbVka1J9ov4ouvdH2/x0uxBbFtik8tCo8DozGy40iYbIcSgNMoJ
qpGGJhP1T2Dz/JOSTEfz4Q62iilPCVBK0oOVdp+OL78Q5e8hXlqfnZ4B22Zx
wfAvnwWhVl6C3baz8OrdVQ4YiJHE3OeNFCRjD5ExYZN0g6KOaZKb7sF/ikKr
2H2x+OsoZruAkZzLH+FtBbSmppWtggwj1fZrepzWeUXBA/ZzUc8FsQNDD6Tl
tCZAnvKmaBKQ3rSVIXt0PONF7PPN28aqMo2TdqfBZVfL2+w72Zv0TGfuVvW5
LmymMn+ezRLoog9YXSxReEkYJsOF1mz0cllkOvqC220AmzP3dmjR9xemI94G
g4sGf5rerTneIkteVBvPrJVZ6Gag/klEhMfiQE6Hs3PI2aWjBJKJXt66QZzT
c31CZg3/zXMyg8PzgxC/EKQElQBl3yqx4q2CQI+rLg/rKuPckgKm/xXzZZmd
TDVsEE1/aLFTvl7Xfsav4F/CEtC+J9K6CuhH6LTYHyi0QDqoBY+xWYXHDa86
/1Eh3i7CYw3H2NMdKJjNnltNq17MTfUHn14sJMdWIPqsP1uiNxwAsrweAdRh
HNOQSnJvFJcnYmznEK2sO5ZYdHkm7oBLavzCLbbQunag8gLLvZ6aS+kNmKdT
1RFChaQcAhUkQG07b+VyZUjyRLXIauTghkxVsNqXA+h2hagB6tK/24SrLUQ4
Emfhg+NYwV6o5CH3Jv9YhEDMRJIqLbsfHyvJWkaorByTFYgSKmEPfaHEaoZs
CxMD9UiMKgXBNO/2+FGc1AE3vo50iD6CfbjoGlsFoZ+f4Qa4hSKshryfY0HJ
wX6sqJpV9eitHP9C15bvlSnu09pgRVSESrpVBeYzTiS9++ohN9Ti2XCJD5+7
4sjqPheXdw8RyZmMUkYzOUbFO5hdJTkWqnySk2iJLiG+1H5DtoxUzbd/O672
48TJhfupkVqhDmn/F177DRu92U/83GFLB5wI4c4x1afjtSM7h033enXAcr1M
HtdqFBCbI2xlk/b+NjBicqXeL5gtR6WSmhG/5oVTN2wlKJATJT6S8d8vf61D
M8TBiBPc0MDxAaNFSQWnq/HLJJHFMY047THcMS5dnfed8pBP1VkgeuBZycrL
INb0meaSfCxNfBaPZz4LiHbTEFdyLyB8jskwgCLlW2doK4KCcCnKhxVMEt8Y
ga20ZThj9QbQPMYENiobE0U9Hw5CFbGNyuIQ2t47GzCPf0+2rsK0tSCEqa+p
rKd148G+4BKjW41RPTWDb+bbYoNWY5CZVAuEyYLJYnuZy40Jz/z5U/f+XjFW
cvocqhgtJ6Hy7/MzV+fkprwNU1XQVp9G26ypi6iw7OptAwdylU1h40uzb7RK
Tlwrodlt0mYF9ReirQ+E0JcJnsbx/3bdOeGrdqbnA+nxS73lUst2jlaikqJh
dzMYw0/K3o0lsNJQeV+pKKjw/mMkpS6sYAWA+XsZKpq8WCGBf+P89JiodZW6
G1fDTQeFdgtaXolEhTlF9xEiMCc0S0SK/Ju9wDtI2D/nQdt6ey8s2/c+qFFv
bxXKqEJQBsdIdQawxZU3j5yGOtgUgczujXJU8lnXKY2RpEJbbyUsEIFauMhA
N9nxNfMWOEbOv6VdsUeFPLp2f6eTY0tVRbRdp2VMnLlxiwykKDGl/KzJgv/0
XWMj9ngCCehv3Tq1HnJA2kZD2cTVl8dN4YEHskbzvCuR6YkoaJDXOUxiyB5R
SWcHOM7n7o36sO2tMhJcLsq15ik+U1x+k9scFY+CU4/YvVaKwhcgJp826QWo
nJvXQwBXPAQLs45Z0VeGKSFrtD37KKv9QVuGAnBtbgOxTS6DT4K4wOh3GP4Z
nRpa7iQK//R1tQ+BlWtalPOVSsXeahP5So+R/z4QJOCUUuU8xCz7g8ilXOf6
oVuS3nFFFs/KDjuubg6jG211QhGlyV+c65AZ7cvkuPE/Bx9Zwuy8Zngc1qz0
bDr+H+0f06h4tjMkpi0FK+c38pilnQJTc8N1yyK5MaVdtd9UpDhvS+gwsn9b
zWMI5TmKT9SHNLhGyUQEKxaz5r8JPKcqlEgo+FHVoMqlG7dTMXVOgKIUh3KI
ijqTEX2gvdozt960LZzcVzAkag/fNr9PLLjvv0fz1mm4T8mfkzxGMPj+Qc/0
mYXmwTQXDY0ip6AVtWFanO2g04+VFPBAQe4ByQSYLbIbvtx/Yr/x7JYaHvFv
YX5PlwcruaOVfnw9Z3TOSi4XIgI0eWk7/UR4F7TEju4EFCG3FbWtDh5iXaCA
vvyNzzDIij2cmCJ0QNGAQIfi8w146afwWx4bBIuPPWu87kOkBwwbklDPegup
YCJrDfKr9KNbLs4OfNlenveQFOZ92M8klcjJVFbIoZziQ9feD05p09RBQ2ov
5eH1E/EvYe/go23s0hK/tWnWS6oxKjxHyVzCjK2Km5pA0/Bp4Qxmtvn4AvmI
iA8r+6I5309tTR1dDarUyhuXajafAKD8ISA/FOK4bCDz244KhtcSLORjV6ep
ADEa6q+hYM3oyqqvG/A/EvsG7ePNq3V7/SL96Lyz8X/8OrHvTuGyBKTejcNV
oiaX1E/f6gjc3LuDUSMRbDffCZJYKfT3jcRW9qqxzVmmEokcMmTCCK73p/5m
AG6/5susFT7woHiYmAUglnEsVP99oClVBD4lKtUKmrPT74/7IrlNg+VOdhr2
Zco5ufFlAbFDN4bbuZApWxwzzpnHsJS1G5UUSpcvE1drJLSZnJByON08mAiI
SHaolFTzgD+glbDcsJG22q3xVFHXNggIava2vybTzaLs3QvFbc7RU2NL/YbI
eZJKk6vrdXHwhMXa0LGkNe9SfGF0toXfSnZGvZSm4RHuUk8t4ASVWUEjhKWe
Kj39viSFFW8WC/KwoQDdixAXUGo+nk1f4vb8VY2dKBRLm9J3vah8U3igcVO9
qeo4Q/DvFPdKTU3qyfuBwyyG1p9vsdckRD67FxrB7+tSiA93liTRdMxTTFrB
3q1z4LwUDZX0jKM9qXEtG1ai0NQQRdipixSd1ScJ2zvlTRvH0qO4iILJvZnv
q3l19sfd5assFEsil5mO8RN255iUhhJxZJossNQaMi2PVH86I6MU56FyPtHS
PoVvGv7P23EiFyxEoP5vR1Xjb7O9RDbZYMG9SuUiqYFYaieGx2cOJ+mo+zcV
IjjaRAEoyUTKDeQzNUrh5VLEz0j4JGpPgWplf7r/j11hSMB9qr1XVZ8RSjgN
9JKJEg/2Tkn3p611bszJezkAVNTtpAsOVjNgR9r06pq1DrdkSCxwgEUzPobP
4eKkHIokFejYEcKP/zfzASJ+sUaFRv3qjiETkhRMR16NPO4VRfQBjVJuHMeT
7+mbGB8WGfIFlbAUQk6mlXYTJgfk/rDr75yBctIB5X0k2noZKA3hiSxLKLsi
FxW0f9URVzAOdQLVxVu9SQiq8uw6mLJB/yJSZfzuxuz53O4mPK1Ed6xdpm0x
T2k1wXgrbZq25CcJMrGkbATQBG4WRwUuV45R/Keeaj4IKv7DC9+4wVOdNJXN
V2xtEZVS+K28QK6LzZZS5yTkOycvKYRZj4sQYrd3jotDZnuynHq24NgIbcSI
17W00a6Vk0gZ8xFsgxKjNkt0L0x80iP15Bj+xUQ8MvRUoGWEcKTgfRvTz+rP
C9ikwp8SvsT56xOh5TAzuzIJG7B/heN4zfJ1iRFHB/TQ3CFvMUOjySXC8Ijm
rN3wdaHYvv4cHVg/IXriMn9brkdlokz9nlEV99Am20IjRQ5eiCAGJhPI6w2m
8hH+rP/+Tdt2AnPPBymLPehgPXa7fg/BbANPx09GljExxkLkDrTxTnXtF9LZ
LLouXNr313dEdbufEBmGbKsXn6VpsnewZVaLyFZE04PK0oBjOiaaYs9CQkJ9
IXyLqtUyc9h0R63ts+xwN0hzzRnNbbLB8E8OdLEg4fFMOUNBc0DHh3RIjkEU
sNAmUC7GocjwW1C9g9Usk/PQ2td/NNU6tHmk75oZjvs/B3QOiVQxzBwn0bhj
h/qnxDDLmP/NbWoYtxOf37ESQoynrwkYnVdQ0uwfgKqZgHFylak1f+s8kAzu
s18PTq/1Dyq2/Kxd6HakNRtsF+5e4fTm9bbCdHaWiylWR49YT1FlPtLEwnZf
6JqN8L4i3qEJj8Q/pFhxCRUnMdYN6VBNatLezC1aJ6sXTmIODjn0tg8Cq91e
bSgtPaZ2IppmR1KCZFRtwROVbEMuixXs1xuD5/j+KNSJBjbQQiYPTwKJF7mc
SkqDJ/hR3SYDMLoX393XJ2X3k3PTS1supZnlv45k9ZYXSvM8alO5lNauzDP+
0PKuMYeHfxCyLgtCX9iO4ERXrrB44dNLaE9Kd04R2fE6CIcMLF7X9iad9sjE
iQX159CD95cTEDgX9zMxB/Uizpj7lxJgGuEb0H+pGysv0hnmNX0lxvvKexnW
19c0ReBFDZuPNKlRKALyoKy3TrLLfih4UX03lX88PoM0h2WIi4Xq5/h89hjv
Hq8XisNdyoAvY/G/NaVpQmLGCqSg+EqgI9m3UFyvbMHvXjPOwxDk7E/dJhtA
BSwojjCoSdGFdn9gnumkgV+O7jH3+AAC1CQ8X9hLm+FZxZ1VYF2FbnB47epk
aMUE0FgnTWvwnbQlYg7Ieh2zYmSGGZALwg6Qb4oZb0fth+gwekW4mwPY4V4p
EKXGxmYUYVErXugYCtn53IzkwnX1NpAJNqJQQeGyjBHk74aZzfitNliCrGvO
kn9+bV/TzHmZyj6+4phY+PwmcBHjeSJ6IDuDF5xAlh+gkRgFOFYqr8AsIisc
WZfQeaCJ+VUzS11qFskuoWZVLF+fyKX6nDsyImQwwCqdnfOJC8DTH3bT1qhq
mzOUIDF92n/biar/mCX78e87SN34xWZeUpFrD966pxLKBtbreU8OlAtwYK20
/Y4HWJJWqsSSzpFBhdyzsieqRY/hR/IQ/AgF/afkRnBOL8a5CZ0LHgMfYSSl
Ff11QwT3V7remvTHMJKlhuTsZJ+yUVeykJmIvOXPQJP+YNg8F0wzrBGFF4tU
y9S9He62/33vk90L/3ILSvhIkxZ8zUgNlBhIbTNoI6qT/WpZGkoZXt7ortj4
2aVMn6+EWbeDoNegLgqP69TpxlrfA1vu2j2+JCpgyu456W2B5hjurJHizdvZ
h9eFpPnkcli6FSXzm8hw4JD/zmgzXeFNy5hmzASIagoEpLs3R9oZanaZNbAV
708suI/4GWqhFZCEjIs2oWxPFupo7kETYvbnk3D27a6QhQZry0EMjtw98q5e
5NdxLXbymEe9nw7KhgDbHhc0n5VWstjqSLvrG3mzsLImG6PlikBl3+8MPMYU
1M3tDit5u1oFlTrf3x+YzW+qfw/pgp3LKJsSR2Jq3kumGdlVC4WnxHoYinE5
3r2kVkJG0XV7MarZaqXUM0+hzRNt2INOtDGJggxI9oq6xsbYc8qyyisBcnPO
R2qkMuUVqFNuuf4lPCAL7ZDbGMcYR9EpNkfhp9ybnIdkNfHxMzgpmDYv9F9E
tSyVBsj+ceCqi9/4VnhRN56ZUeqJLKq9QMk8IjF1GJVCYgEa/Ed/Ds2Lz6cf
7vojZGS/3TVLt7/8j8HZugfMVhNnDrApIHoA1Zvf8WnLEbbXjVRufXdAEW8n
tTboltUB3VvuETJ5PjxUduO43vnwk3B79BWfhcZvgaCEPEYxB1MOVGv/gydT
peEKWazGAMGQIHN803J4w5Si1RLBKwEmhAIKjiUEZuAqCSoWDzHVFVr1FK5Y
h75sC1Jq8uLQL3valPNhoy2fssYcRcL3Ymwcua4/mjsS8V9NoGm7cLo3iuN9
nN6IrXoGI3y7FdmuKqlImZbJp+Um4D0g5fZ0vwF9msaVUfJUnKLHJt7Sm29J
iMxS78bjZtmBYfVpB7Euwo3JSkQuqpWNBZ4NYF9h6Ob05PGbyR1i29T2yXHU
lxKqvlRFI93HlxwghCg1cMGoRqFjreunYNNS3uTQP6ALjEqKPkZnU/MFpCZj
Xtib4RZILh2WEDRjB7I/uySpIyj30vv3uaK1ygr4JHDZ0hjqJVoWTwP62mQX
iPapal6LwhFwdeJiDSzuFSCzVC/SrhBTar68Ns1h7aQDcdva1isWobUTcnWW
ReIZsA8L9nVXhJVP5uvl/nEcFzZ0LSehdCr5X71C2bBQeX/U0Ss4zfP4zQug
KpMXHmcl8DXdmqN/dwe6IJrHlOFDSExLt9pU4RO8RKRtDy29pn32t2rdIcmL
Hju108BTIX3sREGWr+0NBzwLKKN7RCy4AljCDX1HYeqStK3c2m3LNHQdySLk
uxUWWb+ALks9PUmupKCjQ2gd1uTOvYuTq31gFcXNY+AE6AKgSkfsa6g27jpA
ED7wwUBPxP7FRdv8JOv8B+ue87VgA52JDE1Ok4IaafGeIZuJ4VfKn54fQrhP
9D36yXUQjrhaQdpvSBZu+3gKB2DTADVW+Mg+VnVoh3obuZQvhWtRCRoxA65G
WC6bKRN122jp6x5bKfjEUKuuapTQSb3tZXVUCxKDmgRppFIExmfQoEG1UdrH
dB6iuwWFOiB557aE1a1fLnEQ68fYKuECNAplpHH9173oX8yxYrzojLMezsBC
9wsvrcl6jMpS5o5BXBTAs+Hd2u4VrzOAV11pY9xs/AMK1OpEZkzjteiSPH/K
j+rXOkfXb13VS9J4KraUygkA9AjlLr2NTy0rZxTi2JyoQsqnezXRVa0U1EUp
/myy8pdCerf4tr11K6trwUJ+coQjKNX86Oof6/oF0GgmnT53F4McTiUwY1qr
wCCGc7IMV5w6J3BAOFQwfm8CsYk+4kLRiVUml/xiLo6VywwvYzE9Br0Uj6ic
j2mZdJwjFIh5xC4v2/b2o2g9Jqd9Dr94X96X66/pQbwsJAzTzJ28r+d+njaq
j+akdE1IQCmFMB3Bn74dwlFZKLO4Dd5YVPsDp+bO0fSGKyqc3YT8ehWA20L8
XiDPvx4YZlX7d7oDkCt6BfZM8IEF/LaT1dUClxog/cFPxzZ9tMzy6QbZSmL4
94HNKY++8dSGnzetDbB6Quuz6qUtHLokD2F6JGz49v9PFkBB/X/dQk/YL7p+
Au5vDglkAocg2sLFgg2hbXe2bICqu4hbWkXuP+P/6Ugu6VoOm+HKe4lqUmyV
ByN+c92VdCnEIma571tf+duKbG7lQpZPLB3hpzcVyMTTvCALdwMI6umZ/hcH
r6CRBfUXzKgLwIMx4Akj444RbM5NZUfbaAuKt7JTGgxfNgp7ov6s1IHzJ4TP
Z89WGvTS3scypQO+5s1DF4dGuKldgNkfHViFuM29lo+FOJ0Q3VDmGi96tB13
164ytrgvRaJtpty3RagnVyk6jUQXCnWOZvrSR8jI2Myp7qsJw+5UAMfJ1DJW
fStEI/62+z5YQH5+x/9lu3KPsmxEjWGkQjLh5prIoYr1gXSWQfIZHMxWnTyo
/fd0K/xo5nDmrRhdz6tuOEYuCV+vPwl8k4OtKGoCrtMQ0k9hw1HTkxgLLKUz
7ArfV9pNpd4NBQQprBEH0Aue1N9XBTvtugIXhWdjzv8GxiqFvfmaW5SYhcjT
nzxiG4yIlRL5EV/dZwD3MahjRr0HPqIkAV4E+NwO6dF2pH3fsqSampCS9xM5
ktfeQDQqXKch/grUDDeEUelQVK+uwHNnbd0/T6eYvkfK4UaIEXA76LW0lPyl
TJ1AHBwqqxarsgyJ+C1Gg+5QH3Ba0amExlcZ1eCNvQZ4dx1REkgNTuszrffn
3qkDw1JqmVg4dcKbGUJBYq0OmcHqjyCMyg9jxkrIdfZLERIRJRUgy9wd1gg1
21ZN5ApDMn6XAmk9BZl7hPZqP6ZGtplgWlvG5yWYlD9fgXiEE32+jNsePW4N
0CBdbyK6uJGvlqirC8Qs8MGrWOwZ7tfoxhJ6Ttwe7LptJAGBItp0hnC817yC
gWXjMCeybulXRwjYQInDSdisrBAYdKgKTWJ3FQmwbDSeUd92jmPKAs3BWjPk
GkhW4yv2vv3TtTrDgszpzW63mmGhmtAN1hcxLDhFnhgNsgoorPXTkHfXDN2A
Waf5ni6Kl2NcAEt8opLFNsEAOxGTixwIILbthoxbIrnJ8423c8nJnkHygS9L
85gXkU3OOxzU+H35jI9hZeoQqTe4ktfyJ0NV05U8ekazqEb6v+27kaehA3vw
dVKXzczd6gS1QI5VALiukaUCFQuNl4r581DzOSd5nf502hsNfmzQoiZell2N
8RJZvKIx8sljr13AyaEXxI6xs+BoMzYXTsOl36EHdvnA+s/0KdUUaRU+LLYT
tM0mGCW8UetdYd77thA9MvXBoEXEJgStkkeCbgJ8e/aLrhyzh+Mllt2iADZw
huBxBaSlT1lNbynpn09g039wwYQKMUThZB7MrRu74eJnpyQgqoQbQWCocbUx
hnDPW3t0e1OIsVHMtLoCOGUDAheMkF52MmnpcMOQMXBW48jqh06i3RImDgJT
55AfxI6t7nAExSXEUTSM3+AaXfQkiDq8E6QU3c1xQYmqeHGsIPEGKbuMNHDe
SCeBe8Px6pGRD/TYF4vfWSllFvfhGcmeINuRm70ec0EuQXcRlDF6AnL1az7T
vW4qIOEb9X1Mqfg3viyeWzOQj1du0Klgm1PBgeMLS19SE0MaSsz8Lcr5NW5+
nv/03m/pSPUS2oXGQxCCRnhzSDI88ppwiPAgBIasjWb4UqU3JJc+f3P7To5d
0fRJhwYv4oeRixl8dXi46TLVL5OEBjx0s5aKCSIfqhYfnPNpybzGf1LdBzaN
RNegv9Ql8O6M/jwBz+CsZLlY7+26Dl0AqZ1A5Nv1y1QBOH89RFwMD81CHDLp
VnZlwDVMsczK6rbin9d/jvQIWseWpJ9GLoC0+2hhqEDh8qUjb8e61335aH4t
Nd7s3xW6ICmghVCZHHFHNxa8YAw+HvYJ8b3TvDaiIrqrfI4Vlzk4WixoH//z
WzAKRmp8lkHdC3n4We4QfeDfOZCubm050X/SOFDGWPIIcWDjevRMDHuJ6ZQk
hViqm85MR20CznEWXwzhjDZLnz4L9MOQk38kVNkO/I2Jz99mju2XTlu2R/E9
HBNuV5SMemHHFVjc//5w/XhgZGfwU47MX050iM+slRIBmw79XNgzdaBtDu2e
9VJyGRATdiQp5BZZUZuGHY1jhItqiJ5ukqs5pMtcuvdmRZgUTPDjJd9s+sNR
5mUNuj7wR3r6aWa9lpebqefk8qjHhWq6OF9CN3th+s+jtb027P6rWcnOg8q7
M0Ev9/NAfcHrxpcoZF9miCxY8Cj4XtJlMt1ERWiTnYpZCHRCvG6vdBPo9Fbf
uI2yu8WXg1kQKqe3pcOc92XOQWgy9Ut4+aVli+RybWPLio3MAYvp3upTqEP7
mPZdTXESXQyxVMqAUrg3th8bCYPl3kdCTpon3WyTW0N/k7ScbsQYKAsIU2EA
SHHzg6+35mrIGI16TfLsYBrkeYZYaVgapZisECmvwqbGD3T73iy8IcUeDBrt
G21nLOdUK22g5v6bQ4yrrpz1AygwSiTNuafd3Ru/tFNkL+zxg12YezN3TN5l
UNA+zh8dryIt07ha0x5SUG6NZjt9/XmFPHYa+lrD4y6fkfd9/hB/DtIQIh1q
j5aVUhVVT6Jk+RLfMuuW/V+QyJ01Cc8VFNlwpq0xVm1zs2132J009ePgxOI/
RsfXP1NvHWXJ4Y9XFs6uTdlRjzgNhvMGx79FkG6swC4AVPf9PrTVaOj5+gl+
OHFgstiSbeTNDKZFus25qbsopZrzRSOiTEd4KsoOOGQe1ucbAerWD28V2d7/
/KgaexPfkG1hvnMAfwZpaz526oCEjiSXohKEpxeLbDoZZqI5Shvjy0otwzoU
8MCec/VTc6V4AvUxARf9gG1UtY5InyJBhS/44MqWYPsbZHw456UTAeTsLhPI
6qjwvFT4QJaX821DEd4EQWPefDbs7YN9njBkZFSozXNsDW+Ha26zCfontpjL
PlxOOo/vpSf3VcBOFC/adL62GoeigW9Ja2qYJ+t9WDUmJepUnzEHfo7/2CUk
JW9OktYPU6GcLTUJQDrKLSL6WP4p4jRG74vJzxTBFt19jfjnXnmj+WJXpitt
nhrmPTVS0O46hd2KPQkpGRuY1MLjlNQ3qY/q49SQn6yS8tSpF/5bUvfQ/mPS
XXtOcAzbBw2ZX2/Bf1CFEjgO2qt8iSUjZXZoj05aseDB2JJSY5ytnVEZlCWR
aqOpcA5flseM0hNtUKNk51UjTDQJ/YFMMD1hafw+h4Ow8O9YR+uF3g1iBYuw
rWXMqV/jg/RmAOL/gYCNVEvtLExw5ACivHJMxFv4AJgUCLOYqwLAXR1bH1Rs
uwDBf5ntINQPMIfjgra9SGAUV0q7FD05heo2cotaf+QL6A45zAYHZpyfCc3k
AjsutmxHJM7B5J9+ilQ1yNWpFF+WYqjbXcBztiSuzvNRqX8Bn4/3UV61Nv84
9THmv/wFwXq3ErNpNWT6L2nz/4NVyRt5teObz6ob5z2Y+QiKk7T+4ZUDlOqY
k/IP2711ps81TOJlC8lQyIJTIEOIXuaVVICS2NNpOhyf+m4VppT1P3CeKuaR
HHWOyTtCqw8TuKt1uqBTvidxGWFXr5Iks3fQ396erSy/39jWS+l4DoKWTLYo
cNxKr654+esCy6q51pxcSDhk2OdwQLvMyqFWd7zgSZRbhBz10YPUrIpDQq59
8J+CpcmZLAJ2L3J0ulSqfblE9IilBCIZ5Q7zQGi9UY+yg8Urp8VE40J3d7fC
SNMLeBwT4TmfeyS30UvzcVVzzgi1mgu7f6+pDir4v2Lu6gWfRNsjvO1/aMhK
vqHBOC50J4A7LnfU3WyQbri7slXuoYIVFsk1xseOdok0LnI9yvgVUMfNE7wX
UBc+EobsHC5zoAgEbn7jYQrJJbxX5LJL4DB5P4omNhWXJvY2vfkTIq6F3jpx
7FC+smCQF7rXrySCtpxKZ3SFK9xUs642cfSklLQJ71JGfmtWmeqyfH1wSONI
xQZGVTuRJFLytxFla90MW+nkV0HA6T6ACk+0UVuX+WSPC20rL9M4ZeYtUe2S
H+07RZ923GfItqtlp5hBjk2AFBO0LuJYuBZqQaqeDzTuTL6cUOjzOB3T59n7
OKd6G8ZJFt6nHbraz+BuWEGkiivYnfcqkgeTyZxOlPJt3ND4+lr3jmm/6+kP
6vcsA+Jny1mHlDzxVYvLR3fu0Au2Ln3huzT/yX8EM9iJkmwHretmXekTbtzL
8cVO/u8jHwHjzqFrOJcsOcwr15kYekmiPfTKKZeW5+czW2B1TYiqBSsfZJJZ
eTBbozna+QdEir+DhgI2ciiVDauloPMrpUDjbii17f2BLuSqdmzG4uzXwYpx
/xtYWwNSya8a7ScO3zjVNulm48OuS6cj/gogOM4Gt2+fbrqudYr0sK3OPiKA
NYTw6071ccI5yWdUI9kmI+ezCijnmxnYQqTlWWsYZDO1qhzx2XOEl8Tkee8F
7WHACY4HzW79rMPjmVsHbp7rzfTuUBvhz5Vnl9tTIRdx1GZ3yJsU60mmytz9
LfkqYhnjtb8IRsLTKgbUrEki9JQW8ulX1RUI9wgNGqhQQ9K4vwvpXEtjoaRI
vLD8q4l9Ef0/fSjL2YuiU3ge2j4tQoTF7i8ak68Z8NmiQ7hmFnld67kw2kP5
BudSzQr4XfG80yp8t7xuZRirSS/5Bg7g5LnYoKLpPN4i1PNAjfntdFQtPi5B
cq+0oyqnIinwR98Bk+LO3j/L68mIeF8ZequPzFWUGJ8HUPgcnKniIpMvpRDK
E/6FoXAu4syc/rz10iDMywfYjFkQx+eTuvszLJeHSyPVYhg166ZIYl103KNB
7cBD4ODzSSR9J1iqR1/JnIG68QL4/RtFL6KRDLYBd7seSCNNAGwHQzh5FBHw
qJEBIalGKAPhnwpE0UoprxDsxplx2DAXHsPNuU630Ieed9iiEuJ7xI9bk+wM
/Pz7DVg3wEh8tdQ/fnBsufTNqnpvTCrJ/Yi8ANNlyRKFrfDBENY/qwdt52fa
vYrX8kOkVg2LgxLkVcxeO/Y5slt7eyjXJewfZXX3h54I/Rkutvsv2MFBbC87
CRpNe9bHLcTUs+2Rt/tYy/NsEWpB9k/Mq8JW1rpbYp4ulMOcklSMv3RDBxGY
QWozrB10y4/3qXIc6Yq0qjZLGIrCp+llXj/fiXIvVxIKnsKHDzRyWN4rtAfu
ksWGukJavmL16y6Y/Gp5aiwJVBmBDzNpwb7i7na3oGDN36Jv2xKyhFzfuHsW
k7yCd03Cz9IyP+SANKMKtKE5o5lB62xRyuq6G5zerr55WG3K8ZhT3YMBHH5w
mrabHTbIdT27klruEIJK/i0rsj604ZZU0vsW9EW4IDVg0jYqUUkWMu9FfZkz
Rr3u/RY/EMGFEObfmcZxn3SaNGbpJNlYW/yx+QcMdqHkU0CppeF/R3RwBJDv
tXT6LySHKlp5UQnCcmXUzvGViRz9hbDfLkAmv8a9E0ibymffE4w6arUrTQSl
CYFV84lTFAtTsmQJMmnWSjklaZe+5136Ia5Rki7UwerVu9C2kIin+N31MUMW
yAiw+KKO6UbQMLoI/USo5e+1AZZuKiL3R+sauiZ1nh82vIcyGRXy290ISmLG
JGGYSnodYefTQBlVtS4VSqTHjNmCL/CvYOghRPOUzYE269QVCEpt+gdcn8wq
xgYMi6Cx+XsJ9BBjoWgVG5uJGNrK6sJij2vGp0j78msDYFvnLIakLynZXdul
OdDxBTH6ydFomP3BU6+HqtdQwZ4A9aK1cmW/GSl1uGBq6JHaTocaqgHE4snU
FgmtwjRunIxgdyiMGLwQFuQisv8RgRlIe47iTAHTchDjKeXIKjt4Mttpgd3k
wVmaE8MwHMaYKLfYwvPXAy6iUC3FZBuu+2gB+7rJXcE4ZipaVxC9KQuXPZOn
11q2TMtybGvIM3e3wmczZlPcJ0PMqMT1Rjuf2sKJZfYf059fvxukpTqkjb3f
+tByqQcdOtuO8QwHVSs4LOGrqGcBjd1DEENq8lUW6cbTQzRHD+T9LBizdwYq
M2RA1L0jOKqWbiGctaY2ZOOVFrwV8n3Ae+kyypZDopLKmPRQjb7emWpRkCZ7
+sEEMvV5lP0vDuGsjAfuqzxsb9FB5tNfl5eEE2w7RSwEluQrxhx3wOb4RKsZ
aW66iYEBwpq0HLFkjiRhslS2yUe5Z8nJERrX83PEHsr5a47cn+3yeve1qOsT
SLZq+vS9iUP9IQz/HUXClDr9qAkp7NlbuDR5mVJQhH8o0by6nlSDNUwNDtX1
4TcM26vt+FIUabat13C3jMpfvreybgJcln/9+dxJN6xxEhJUslO/07I0730n
ubMbM4C8nWhI3zmYFS5kauYh8Xa5mHHcLupPzREhgcFX/is7/gvwqFUPxgIz
uj1cLwj6eY5dvSnnVcwnvtLdFM2//ozVYhVv9s6Bl4akn8waLwO5Up/pgpE9
fjza1Ox8aOx/4jS4b0HhLtpL+3MPcBOj5WqFScwEBLhcP3hDRj5vM58bzlBx
Z55B/MiMyuw26OXzUc1i5MpNT5aL6Ip1o6UjkvJeHdEVyImTVxlKjoqeQv6J
O4hsKMezJ9BsyFyNnsNVgmTjzmmJbPaL7/msl+Os0Bt72O7oTG6+Y39je355
e1H6X7bAJTbbfjY8v8/E8jss+7uXlxk4E1SFBT31JuHnuWNMpvRr++CBE409
o4UR4Zols4cM02E/ufnMV+kgbm2D8uUIo7aWAppq0/dJIrZnhUc2rLwHM3K9
SoWhrx4Um2sMGQ7RPAUezIpf3O2PbIV9ZhbvZps4IzkguJ3ckElkx1uSBs1m
uGQseMXsDsnIa9WdPhfX8TCj4UZc6+QgMNnXCtUPDx7Z1yFi90qGIiXY11jV
NRYNzmBrq4dpY+MnoRndK2UqpRwoYDJEyA7CQYg+uBLysiObxpIZKzfvmSH9
TV/9Au+kTI+/WK61phyiQRVPAA8Ezy94dYk89Uv1tkQq1GR0zxirj/3JAQWv
JBWIyYAiKja11lzxu2NdT4f/bU1Yy0VQzdc8ztv1a8E0P4IqO0G1QK6FEOwG
YSiGdg7X5o28rVCq+VLuC/0ndhtqEcsC+U7Zrn1Vt2RFsJXdgc58Jjc+XRjo
/YltUt7f0ACJfckucd+/e2BQeljBWnV21UDj2sjRAXDSIbQiQ3aBy3uqCpF/
2rfG7Y849zK2kNZfpdpfr3lJvSWak7ANF5gI990qIh+S2w7iz2cgzPgLlQFK
p7MwhfIwic1zmwx3S6Hq2FyqcZqOm0iD8L1/Jzjg41kxLkKOeWXqGNLyzfnJ
F/US9bHWDgmSVk2qOI9bCEcsiXvwg1TUgshMwmFscqZ8LCfgrA0AfAYscPpO
+Qq9tq9apO8olwEgILLa2SfZl9zPLJlxvgEAAR/606B9O+Ga0TJP6z5y4can
nJCcyWloMVxzH/o0WpZUxnyxjQxaw+H70JZ5JiNBsyf3mVzTOrO+y4AvSygv
BXQhihwq9AZd62XjobTc1Ux45jr/+TlUZhLRhRvefr+uWRASYoFcXN7Try5A
4d1AMBkeEK7Rlioe0xbN748Wm7ghWfazvdezDaWYulY35sE4GOqml5tKcz3+
VEtSJBo0gtDMC/zqgBSrJtPZTsoXKN64C7Ul992s7Cwl1OP5YvdQid/AU7mL
wINDuh6b8kTkNH9HQnJ/l2oX6wjBRqHX/DC3HMc5FUAplKLvSzBcvGtsUU9A
OwdAayVNCTSfdK0lOK8bokV4H0Pz7AK8AAJpHE/ANasMUNssi7MqC/cckBvl
126LKBdRZU/MPsK/BodZKuMFheQFLSbSV5iDCRP/Ja1Lo2xy9l26RFcuC5KI
kUAE4fJBvQAlu3xSqhRw14RkRBRSzP36QdsBmUiQKiT6rORrCMW25WymVqAb
jKpnWc9NV/sECSOgemYVhpiquZUbJIfKl3p/B9p11JbjDhSuM3nG2Uz7baPh
resTYGrhhr3u4ASvMNGKfzkbf6Dw0AbfxRtsOLlp6OCx1iBwDL/JsLIFg2Y5
wa5I/zkI4gqjIH37m5geM2cnYhWCLV5wuphLEkxirUUJ9nDmDrM7g349noK7
UfM5Rqj91WeldrOcL8fyzYGofgHNAImyC5FNlxnt0OBWsoY7+5UY1DkWMa/i
2YYTRG26wNqXf6qgcYy8V6Q/xD2xIceUa4fkyhDDrbRh9kk6SFtngM55OQK6
JuRslNhg4Jdw8k5Euy84kZaQeIhAcdZanGyFzWLisKs8aje0IfbUfQrk4Ofm
9YMr5+YPufnAdWP+jV72AOu5RVstCRMJBPKNlaj+mN9/+Jfx7241T/3MLb9k
Gn6/pSDvBnPK1rdj37DgN76sZvp3dg2O5Pa1oXYO9s+i4CoZz1muPjL1FtQC
QzPILlSpnTWgrCbZlbntk8zZtUbBa9mb0ee9kME/SHOJWPFcghKvJpD1hZds
4c3/6T9P2t8FlNVy5fTyFpCd8rOPUGOfMbuA8unX8GI/BhTUHGb6UHHVnK/B
BDxWdYUeRyqC80Iy5peQMnKFrvTx+CE0boiodNsrUq0pTSuJG4lnTKqfoooT
OjFU5px4MPPD/y8vFijY7rQoifjMMp+29xbbdS/Z1Gg/tti2AWZSf5bTJljI
KiuT19gh55PI88qx2yFcTfmgkFAJbTRaebOh3z9ItT6VXAs4BmxuXtrjW0wp
3LBiu6azIFVzf1seyL/o30BEDA+Zba2KEFklK28Dz9NES3T6rEduJ2sPV/ac
JPECq/kDjeH+n2zZdF2xJG0pV9u+MuZimeZAiC41WymIH63xZ6U+xKEexAM2
CBUxRmGg/1/EpW4SXTsLmuEngV6KA+FuYm/KsFOcC6/HjvcMUTpU6TpmzsVs
4JKZ6RHR4AhKIlK3KKmBL/d3J2EbPLBWDEgue6a0Ncl7+rWFzVWCIeQ88qbV
BflgNxKdpX/Tjb6QbGbcYRgXBZpW86FZ5DBY9+n0s4f9ciAxr4aYe6nRm4px
hBHAStvi8L/o/O7UFI/BX97fMmrVB7Kg7TXv3aAO/mKLBj4/CWVHfTCS0LKI
JAto6mMeyMxPgnE/wo32Y42MWf9t1vlfi2IqEH23HuYgs6IcLYzAVIBlM0cO
YHBweC5vyyiYpMQ19G0qvIHEmnqLv5Jyu8EJZmbVNvjk4W1lrm80UV6wdTWG
nmd1T4GELIdiLlHtbonDJovwKSrLjv8RguYZ/q+nSlwf1LZL+I/s+4kiatcF
fVbvXuprHkkiXtqhELUQy14yCPwSu8cm8RTQ2CPiWBvzPzxLEoRV3CREOzNY
wHFswxpAveHYyd6j/Op6ZojtonnxcQGL0uLrFASA1qwzpb1bDJmZo/Gl8E6J
ZIGYMQ8ty9lKjFx6H5CO1e/pT8WY9NTfg0W2NeHRSi7oZdukOfhgidy+wvv4
f1pTCa5KLQbcvcGt7XKWLi4CJLc/GnpLPe/Txz3VsmrpILjWNmk9Zq3VD0LO
3+UJyQ73tyrWZwhX3wMh61Ja5o44o11+Oo+kUn9FGntPHqs7joVLR2jhuQeP
5kV/m5GWOO+AgOIGUl4SLRN2gx8u17trD0LtwH8LhOG1y993+AQlZKbzPvKm
m6yeKgaxyI54pEhhChBW8dmj4fajTISOaa5ad6TTF+2pO6pMSsZWm6Sx9sJl
ESmKVGkKrmm+L4KKsOgIo/SQ9i7xx2QBiuIMU7BvfmbmMEXQdGYhzSD5Dv3O
nmoT1Ht/suZIcmdJQ6sH+R4TxA0e4rQKWOJZ6SPXV3N6JJs/sPFyetORdc1J
finnmVwnYyJd944VhekRDMRXK0LNqGt4gWE4ohkt3dd/1VMMcuyKyMmUCPhW
9PQOubL8kMMljo/ArSy7G5DDrIjvr788hNy6YKYE5A14Ewgr2LlK1Jp8jXgo
DfkSa/EWGRVSU0jvzg1pyH6u23jnpxCSrrmvoGQOXhximKTTt0+Jios1gztv
tGhv8ch5T4TiUrI1z/oyk7STPdNbd8uwg3sGGreWGeL/yesYnqCqCyNAXI8H
ykwMHDeFGHMgv70v0Af06yOVgdqa1x9FeFuPd5HwoQLlhHKRK95FCIqNXD8f
4prUsyD4Y9IuU20gtmLVxtKABANY5i4c4n9Zw3WyG2uYYn8Gi9jB84kZUP/T
d8Aq3FqYA64LfxBoI3ouxgZESNM4IRa/leTZrSylShkr5rb+w9w0bTpllo4m
98PuFxn7bRKO35FiET5EON4fH+S+Ve5+D3umKwyLgVhXOThf9laysb8M33Mp
8OSs8D9FZmGqQtbra0z/ZPaU+n7NVV+freD/sJq8PIexkuUjUxa5VIG7lEEz
lhsL2Di1U4Au5tE2wFUHUWKZJOE5LkzUPAtpr8HaGMuXh9IHgSNR70ocI1aU
XxWnNzzEzPWkdClBXF2o4CNoUelLuWAza797m7tYL5yvy/zDxHnOiU/DeiEB
yxOqrxjGOY/0NdI62Y73saFFvgEKBAhFuC/DIn6EHAtfAYuhu2JP8gV0Kh2N
DKEvh5E0OhH8SKtyYBlM09rMX1VvXWCDKeLJek1ftk7lVAdMVS16hpCG6KtM
5J8Klniow/TH8srUVkPnNmSSc7uozoldqIeO12UyIMELbrHgkvPtwOLUlnKf
dEO+djGuztjX0XtnHxs+kdBtan3FpSHfdN7JI1mSlapMdn1biT0IrpPyQUXa
xmOG49ydaGBldaNqWUoDqSoZh/+sErQ87j59nwx7EMgjZPpuqmKNCNU9QAKh
6yi+1DDqAom/Q9vm78hIWKmSH0GL2XsDBcJu3KBGnBM+OvdnJCGIuFl9Gl8o
tP+8qaIqnpgOQxIz+8r2hqT7LdekQGkbC6esDdfQ0N4fT/tm8MFopBu+eTWx
vMfrRVuZq0OGhimrADWsqamwExe0QtQPvwJmR7jrM5RArV8K7VI1Yqb+BIJZ
yguFDBdL8yRbcyqueP/QQiJjs04RmUD2UkpjdLBKOKxQSPHMoBQHwDKUXyjI
XnSyNlXhatU9qSCYzO4jSiVBIWVJv70D0iyaCwbbYBSsjuckZUstlobiPvSg
rCas4jL2VryYi3ZnvpGRhDn8d3aes1DYaxuba44dtRsvAV/Pw14LhQQx0hXs
BsYbmtP8R6SJvfoef44vYXMpgtlVfChxgc0cm7sjvCO6BWTfvHC5rWw6tksk
ro/1jMRu1RXMXpN5/RH4m5oYq0wqYX9QfF+V2rhYGCU0ipE/H4oRk6MSqa7F
l0g44RE30wJNKsSy7pbAOqWUvQGLbXPRejMO8ItA6p0Dv8Mq1XW5kj7Ez2OV
zatpDEBpUieG9QI+ROa4HWLBZMr4Ce7K/NYhrDu8vCE6sh5q222/8pCPYLpC
hdO0wbtLsnDdCkqNwBW1CIYqCxzQBggwiiO4UCnasVbGu8oLsxj0H09KYu2B
wqHLjtJlOSbRxW5gVwGxu/Qu2qaMwSfqKcYwBtcq/KIgXwN4sNBsfA7p1QqN
H58JiPA2EEY35YtFEVJ5p5hpaCAwfCVdO80sX+YliqkP6EZbVNLNJKz2k+c4
kMCkKt6bSCYRt2Y1LuX5/JDPLlZmFVlltvLi/ErICawdwlpy7blqHXOqjzFJ
rxx7TwUZ5DwWN4inXWn8MhVWHgy/JMweR/VEB0mv04YirkTyUE6sUanV7pig
IyUo/8NRVcnw8vmIAL2heFJFf/z6smpGKpVeAzAXU63YZFzojBCG5UBygvJk
pN+GjNj990hMp0d1bcuF5/0QD1MPzninw2ZfuxWP+YdAqdZH2NBuYgIpToeo
kQ9ijeUtQ+YtNpPdf5m4zlXCC+93yp4c8Rxm/cZodtUdMQG6dGqQ6C+A23z5
vRwBVQJM7Wj43ZZLMIxuNcqDzS0674J8WbO6Ev6bIqVRhEdUE+yFb7lD9hcs
4Tm3LOwXwfPPXMYY2Gzefhzu+hbsV6RkinSWMm23euugw2NnO1BrGDCtynr2
HpUoaKIT8usbhbcEAGN+OpRTrCEkw+0I56FWtoxhYNcGHEKf7E8stU57sAmM
9EUcBRbhNyVTbMFlyDQwUEV+rqSIDSKAg2h5dbbf/7X40TryqeMzAAJczz5e
BTNYbs4tSrQpu4ZXT4KbVZHWiASCPMsWOrU10q9t7WyVGxp1uvmst2qHbjHV
bLuzaKCMXRtctr5jYKsERo3qMO8Xpio1Cx3Qvl2PDJGdmyRljW6ukgoBj7Wq
G/4ewoi3YEgjHTTAXP4qdIkPV9GLM3dZs1eNpPwJTjRrpmnpDsotAX99gR9a
lDQY+HJ3cXdu0S35jzdhl1g6eVRG0gvQZtqP3ga/BqhYRtAumJh87AbxDB8s
6gGXFOoh3HZe6Cyvv+SjPtQsTF7gmkgfwGWtlHw6UEPzDIg9cBhbVAHUqQRb
uKl0aG1LSS45BEa8L7wTor808NSdQHOB1Krfte5Wra/vz1gfEvF+I9JTjnuO
kZCU2Oj2XSt4oP4NwLDwaEEoiFK7rPxRXpC988CphVulh0dW52Q5w8oKonSv
2v6HMWLVy6CbbuxlKGe7ou45dGjdx/BqG3JpBXPNPa+U37m2tCIYb2UD3+n8
+5loucFSwMuD7NJQaHXOa6PFDXq3tvy2n0AHhFByGz7aathIZVXRKYBkjzM3
nt2k3bcBs59Du/qVkETsUyIxA7JgzX952xZhdMc511ewqWrY/fsUNd9Bbvyq
MgAv34VPFtHz9XxmxaWYMzeCMAP9LsMEQwArizqzaDM1IZl+g3FOSO5CLiqw
7dvrQnPonBmTkGLSR7v8TP5d3S3fh2sK/ofJpTENZj50gpXGdDc7nYx/c7Gn
VB86VVj8cVzs4/fo7V2DQiM9F1cnXDKflf3WALjFob3s9AG4qm/NoQq2yf2O
pJjCK8lz1a5k0Ot2TlIEJ7KzUAxLTjl6VHCS35jhSBzqvfiG1Y41RVo+Om8S
4oMFQwuh6Fkay+LbBPBlYo6jHn7yPsQL3BNq+ahV2ZCgBivlMnL5TBt3s9Xa
NN+P+jcH8Or4w0WbZayET51Zr8fCrc3BR5/rRZT2c1Zwj0w3GQTNHzHDlqPb
0QM8UEJMRLXBUkjF/qky9cHpBQCM3QdfYYKRkUOQKWMOojkVdGwbvYcVLSrU
5DvZgKnQV97REmdRnI0vrZIjE3WAUf8REfQY/flrsphI2uD//LTlov3IZGyE
kc+z02FluD4J56igP13tDPdG6HAk+amSXskxInk2G32Y72iFu7xX6qg18/X6
7F2dZhKouPKlIXVIsrINY3y3/nwE/CB+TMVTrbOVc7m8iQg4GYztl97kAmum
EYYKFzzJrjCYXYpwnAQ2DPCrGzrdLcksIGIgXjsUaNY6I8rZfFcptdEWkk0g
Mjp74g5NJV/YAGHQ3IWSZGV/jRD1HoSnSFZ9y6Hywd7K6CD+SImwEJhc04Lm
iQbPalb+F6cqTG3tDrIY+i7JL+i9YoXeKPmiUbYOcW9WcvmEedgOJddKk7Cq
qkFFcal9bxIk2vdLU3OrLfdXIFg4MYK5Dfq6C/iEt6sRPHVl5qVVUidSJ9fJ
TzLj3qfUr7VVNMjDfYKeO9tnzOwlIF1ZGWTW2bDFIdWJfdafJHg+kMZafHHZ
Gtf3bk0ybOUDZxugsWEBpnuIqhE8vE/TKCeME0wVp317OkRqQx6Gd5eDvabD
2Lh5BDhyqHNFWeDg7YJufsBHdJG/4sJSS/iDOBkHDKdlpa+F5j3eKx1zkm4Y
YA2QEiBZp0NNn+FiA/HPW9vWGyONrIDKWkzmj+yZVWjaS1NifZPuwnYP0HAj
3jPkigRsrpXrlkORCQq9kVmngZM3/yZwz8yZvdsjOdfGCTOufYYkZz+FD1us
bpu24Y2K+HotArbE8xrm897DJsPq8TJph5FoGds2Zsqh/7rIq+DpJCkHGLkq
2lN2v8lx3ywU0W+WT9+Ib/55mE8F85k4p7zYmd+eFlNpKfdzXCaGeNDwtfVF
71vp3Zsud8BUezjbc92guzW7+QLki5KjfGORq7h9rkFcKWfK/1Q6epby1OCA
5fH1HeE7GmtVlziUltWaR7XcncltsPm7tYvJRs3HeuxjhBoug9Xa6at9DVPx
lAvbYc6LY9//p1K8hx+N/lGu5Cj7t5RL8pv+7ZcUKKCqIBa9LiUcN+eWV+P0
IypeaYTHng60MLlK112OxNCWuiUcPnxToY1CDiNcmSdTIzW7Bzv+rE9CWidA
wGY274vBQ8AgDOtqm7pO1MXvhj2aWNL2zBcQU1n28CcsgzTT/JEVXWZ4ewGK
mB2zqwRS0Usfxqrw4Inv6+2d38ZolZ5V1NgxPG6WAUrZa+wQyMFwRcr7LTZ5
YQRViBZQAmWdDDfaYldq47ouj6vgzmB3jPC8/rh7tODun2ETufUw3ubvNaTh
xcBr7rgzZ+bDs/Ql1Oec+9oXdYChUUA3uEpGvLr388zk0Qqje0zJBgWM6OJy
oVCSWKk6cO32gWhQwAKA24n6t24KbbiW1DXNg/fEJwGSPHeuFQ0a/2D0XF0+
ivy18UJUU/o+OP2Ju3n2LguJJpZK/rnUqsh1L83DAJk1I6tDd+1Y29Tpsj+U
X4XX1GDyZQeBYALVxbpGbUdjXmO/ewDvYtwz7rlQEQIIndQzQKdZZz6NqoIv
AOEAUWnwz9tii0InonZHwujId0XSqLamCCpDaxDSxw63Qykw32avk1SYxs5T
+jRETNjI45vRRBjo6SqHdg4L84lJ5WPguUADwrL3PQxnouzDUzpHxG7xzFgn
buxbL9PXW1oN3282BIxOw4vb3T28J/ELXKWDfKGfcSzrD9WCHZ3odyNnnaxk
yde7hrUPnt/1LcK30Sn6JZ5aVwNDnYjpBZD4qSSYWLif2jFrSrmLGglb6GUw
PHsE/gvz6z5Fkl8ztHroeg6ZHG/ig1mz618osv80YTHl0DrdezD/XmrgGuz6
UFkTHIXpoqKfdL2LhO1YHWTKejp5glemfiSjt2PyBQzb3/rHOQBzaU1tU8ye
wSCem+dc+uRozwfVY4h+i6GI3t4gMEI+d0bFL1PPWzMWZPx5S9N9m/0roI0e
G1J0Clwr/u2w5qgVXDX7WeAZlZYYFOD/S+IZnyHDS2BILBr6wCrJ64s8VyHD
fo/eMcJeOqBUNeAXQ1sTVCzvOYJPiYKE2ESGDpXNAxWMhfvhWgGdNQ+azUyZ
cJqmlmAyfSBVTf1S2SogI/2iStGioxP2Ac2Nby7kyd26lLvmOuEpqOo6l0fw
j6CDlrvktW5TVJOWCCMFbSYQWnthqYdqb53Q/FzbkbCq8IfFHc6DpraNLfME
8fCEt8VIzSkSPouaf2wJ748xFG/SRLP/AQJU0bQOX6ionBebQH54oBH22MC7
X79EKv6ZomH9bZDYY/h5LNiftrHEuohpYZNgAkq9JnUN3q/eeKYFf/McrG0g
9kO6iY9+YauyZL4nMlXShmF2Q+Bw3VN2Dcjyda1t0xYbpMYqst3ZOostgpw0
w+bNZmRP4oFSMbnkXDkOK6wkZCB/r8+BrP6baOcl2tYTZyrPvvGPfIJ0RK14
5fOTNsEviIPEMqck/MVYUqR6xF7SmSf+EH4MilDMeMWynIgozY64uMra1zLe
RebHJTAgKfKwBHfY9IcEQafBE2uS6BohCB6HJn8feu9qWWFwPzISkpGh4w9b
oRDETSrOq1/rCsLq21GdnVy2R7HnZF2E9Gc1W5d89yrSEHI2JRpcuI36Gfgy
MG85ZtQIwa5P22jAZ42wUgc0K7jc6CHIT3UXNQ+EHEmw3abGzTZMC0uA0F83
cJVRK83EoCMS4xWGlvX0c8PX4Xn4h+O7xjw5YRe6lQI+Ko2Hl2IlJ2A82GOE
vdwaAJ4cdyAmmOx3bal75jt9QS5vvW470jjVT1mj/G7CDg8pEqtjLCYrvw+l
8cSH/N+V4unNuyefyCueqxmf8t28AiqNcuyEHrhAcjNUNh8bDLlWSVA5ewnX
7YPVQrBl/AhZ0Wvrn8f/pje6CU5gG4mr249fhf3e8RcvKAFUFMeitcyK2EtI
q/g7vR11jbs/fXJkjfKnncfVpYlIldruCt9CcvPPBaMfROgm31s0JKMYmnTA
mVHw2psS9YX6ujWmiNOpRnNElUZ86VkDxlTFAc9SzHM/Oi4CdqmEE6RDKwJh
4uk7Ae8tJ9+CnoV7loVDBKsRnI/rwWoqJliYY+qR+KJeRct0PFC1X27seslY
PwRtAO6p2xLVc415+12Y0Ev259PLm9eWMnAqJ9Q2fmQh4InQyt68nUKQgqHN
4X6VSGs2iUBjM3ptCLt4aqrLR/69xyyyuIQtrGq2k4qfg7jY+9OJ9e0fQ6i9
mTLdZLeWLVjcsihBv/iqUg+7vfQf1cta79mv+6kXDah1UJVVyE9Dw7cth7/K
o0YQDH93WtC/xcxkB8XKkw7cYuH8PIxmSOW6f8TDq5AZiqfoKFxQYrwQLMA6
zMUJPEUZK0L/cGD4nC72dQ5ebiNcYufUpYlZzpJ1Gwoce1vGZl8NGrtiqZGN
pssXOBKW0p1avEKI59fQiq+hUgyns5DO7ansWBK9pI+8CHNm+QUY52htFbTU
Oylv5YpNyTFwMyLBXgdBPKbDMoPKfNKkI73zgtkPaHhWEmdOzncc0iZZrP+L
Ntl7b8lNAkgj2pj/bmuVi0hwTZIHHjx7qL53VeeVeyNyv72rq1+ESudEXdyP
y1jKw4/deiTdWag4HvkoNItFp8FVwpRF/ZlyBHV6MulppFz2ceqe1QZRFwBJ
xJ2FtfeJmQwFfZmgaBJ/b3S3hyOlA+D0wB99kvlzTbFts/CDvkZmpwLsSZ0W
Ko/NPzSfnszgsy7xUxBo0w4WswW+ggpMDUwVev0T/TxXQz9kwaHmWvRwzZ5r
sXsEi6jO1iai1pjqoAmHLlxNItAUaNoFnVtO1SaAZP+YjX3vcbmhR98etLYO
SYeXn9zEHYu8xO31rQk8e1yYEBEs1OmuGU+c5wsnUjH6MqFC+29zjk8zPQQP
2TKI3FKQrBVnqiRG7e0/YnLLycjsBr++6KXreZBlhlD9tIaqea4/oNtWAXyB
1jRIfyAHCBeCwA916EGdabvZHdkz1dhZkseI25W9Txl+OKjJE8VyRJBI2GWR
5y6QdeOXnd0PVUAmtasJOHJIszZG2PvpSsiJdhJflVAm7pADVSaDKyUV02ma
YmFoCYrUVG+2x03InWGHdDDHsHquomZkw5m+X+ihSngvQ7vrwbI6kw+R1RXS
hsfczznkR0KkkaSQRBMQPSSZo0x0oTUkWzC35lHA+xqBmGZnSEYNYklksd79
f5ruV109soHVXJuzbd7eMxmPbOInWaVOt11I4durqo/GaHbbXs2o55Smd7Sb
yh6KNPY4HhGWd8rJV2I9Q8Em0Vn/lCPIcnpooV3PCHITZMHT6zGpZesLvgby
QDV5XaAXnTS8e66p0oM760MQriOjIpz9Fyr0oC0DLDzATrQDNXg52UXC50Vc
VfIhSYjRMUnq1nKhM0xlyHXH4E9rvabimSF3zUuYGth3TpcxeTS4kEe4AtVB
B65/Tv7+BcFgAzFF+lYhbQzxGC4kHpw3EhQhL4G7seNGB0L6BzH8hvwMkyRJ
5DLgir5TVUDRYMdEU7fg7BaCnd3gnE/35wTKfC/QAEk3qgs1K2OO5mY5Ij9t
FQum9P2xNkx+D4JjYbzHBgx/RVDIlVoz7VzEikujomrjm5BYHEmcWUKn5hD1
+1E+rnWwAIRoN2EMbya69UbN++kApEZV9OTKTud2nUhVu9O07JFb1DEAdKhx
4atmVKOjh1GCGwHmieQIzn1reFMpa7VnotgQlt/r2wSRfuiPMFMiEMEYs90U
7ozqMZB02N3PCM1aCf1F9t8StJcJqCxT8DKcKtFQ5rBjdkcAYON1wsHAdX+Y
ufvMtG9bADLIoRhtEVBQ7Z/K3sOiQ/A0i1ZipzznVEcg/bnK/8iUiHe5ZS7H
SOhTwnUk8W+p2lqwzlz9lcQQ/JT6RguhkSGPsKahYEcFC5wmb3hhkhP8XUH8
3Jx4E4BwAo1fGt4hydxNYcn/wlqSwn2i9xLyOb+P4/+o8/bhxQPIe2AAa+oL
Mx6hNeAfzbtWi0UTR75pDD6DZlOE3lp+ttZ2zb46gtQKYlDCen+g4byNQGLe
J/NhJpNIOEFR4xeZgfJQnzWSEhqbqhJYQ1obd+fm29C+OuU7cag/7oUolLmy
08tqAQYTzmq0WpphYpJWL2bqUgoTao7fTaxxlxhhe1R2rHkEvAd+x9kSJPt8
6AEhKCbkWDoYadWE1JCd7yGJ/v5C52x63+ZtkTa9sOAP2QMM4vy5OizPYL/L
BGtome9iO7gozlCK6ztOTVi4br95KwK91LGlFTFzuVpMBEQHKuc7m64DwSJe
NZYomhdjNHMx2X6Ylll+9L0o++qw5h+5f90foU0kZAqwA7gUNq8qUabtQw5Y
nYD8YydM0RWHNQE5r3YliJpJyx808ETtOImWw0N/ToLOxWVbHa6oQ+V0ew4v
XfXEA8FsMEEL4OlAp/jdscogEdgEO8oYs/RA5eAW5olSuiclzwwxupyOZM71
Y+DR1ufTI5JLWM/nR5ZgNcWv5W8JjI3nsFLMwJ8QbDieQw66oR2v+0MBkhlv
346oihIJkCW8CmMgglG0vOPopE3QgMqiaYRCdWTMLMB4bAfFQVcCUmumCDpT
Q2AXolA8hRvYV6yMaZf+MccbkJ7lcI4+81NQhNSwvj4R/THI5w8AFdk3trQh
svOdUmdJBA+nViKqbNZGn0/GNSFr5x1YyInj/w84F1yogB58VmD7ZmA6xJJj
oVFBCzBB+I4ivCrdnc9FfTVkIXT2i9LAPMgNGyqejTwJo8S95o4MH9zlMVqP
AxeqacI+/f+XW1mq4h+O0vmaiXDeEmNWU4inHCyQ8aPGXgaY459ZeLGzb458
tk1RUovuihz2JCJI4VnwIwG+HT0PwtC4C6M7r6tNBgMqCMF7kOzjpWYVrmyg
TEsKiXL8Z36jEmYQOEgqMvmBILTsqoSadXIe9P1r3kRXMewzXuIdyVyu7afX
Sxt93J6TA3+wFcUYfPYBPZGwSuhnZ3yCnUL7LeYrxRiK2epegaYA3w1ez6fp
+cE+uqledtDDr9pCgGzdJm1JKk5N2BbV8fAIQm+OBNDhpoQRUp6ZG2ulHAUj
mMIFjny06JtJ2GN5dZnN+R09E9m64HkwlGxGE+Co/U078RY1PRNxlT3/gGcu
wbdMZipTppWZ9+IPxgsYaeMPq6ArKS5YbJnDO6amJklL6tgJWE1SMBG1yxRe
tF9hygADatg0LRfb9ZbkpD12xpBLXiuXLL0CuJX24KTh5F7oyCQcdS8lFDKA
NeAN1jTEVkqYiWYVWYbtoYRifCUxUNz9hmrjExyO71eSiDlpZ7clQcODu4dI
tecU0ya9Qekhpq2MurTpBiNUAxLB6mhi+19qBBk18TEJH/m1GuWkFaqHpx75
IzKA10ylGfLuR9Scf6UszCgAuAb9n3lWTZngTKbM0q/roK2YcQ4QwrJMUVBu
0EF2A0/81GsYfMlqh5yI9eIfHACk65D3+/jPB74TEtZ08k4vPP5Hc7jEZTEW
iNGKp71mC/woe8lklUWnE5hUq5UjOZMPJmrSyZMoGyAzxnHb0y8wYSt0x6Vt
HsPf0e4sZ3flTae5pPqUzyZiv/XCsip5Wyp8q42YuSq/2KjfpEkI46IbU6N+
PCdwaadVO1i+eGdbCTBwyHgqmuCO2ZHcunSTdGgCTBlO15skZzvH7qoU3u/C
UR07+2alHAQoRin5/Br0zMs6ijqojiQKjgITruQsws78e636mC5DAHdvRavC
ycFgJeroeq9ZR/XLLcATRGCW8H2tRpum96/Vqe/+BZXpVTBgmXxQBvIbAkqo
RyrxQmvxcz+COnweikhLh82OLClUpnFxOZKL09m7Ac88mtF/6YTlyodrIPiA
65Rw3iENAYMO1TjGwaO9kTGptT17BV5QCh1+lagZfrwWXpbK7VYGBXvY6nOA
vashED7GqXazdqP+7qaVKsEtaED6+CqVyRiWBs7G47E+U6ZCz3woQZ28yA++
bm2JSwJvCC3SEtP8jSQYPSzWAAFn6Jlu6t6uaB3fF7O0ogvMn5Ex/vYO9zjo
zbWoK1FJqJeIDv8NzXxLVs2dbEu2KBShUqJpiFFe5GznR80ddR6pvceQUc41
+DOdIgbcyAdoYZQqB/dX/qMThapdJog/kf7a0alcW+t9/yA9yIVFBYHQIv4u
pQWnAdMMIHeSsV8RRnS75/I6TD1hu4vq/RYDI6oEasqz90j4F+dlDajUHS33
GciK1vYl+xYMmBxq6mHDFKdknIOQ8qriKJuFZ36/fFRBY3IoJgg1AVLTEA/g
Hwv7pn/6sj1wOp3qUtx4+J7vRLke4K1hDOaOQiIsWnGkL16PY95IVaQ5ofMi
3V2sUVKMrYwTsSXa8w/nDau43pIToWsCuTC0D8rXUNRpYfJ3to4MhO6Gv5RN
g96jgKroXoUseNWZIx6jY26BFbuzOxA0RqL+Jgnk/iAGnu8vg6bBwikq8BqW
1esX5O+THG95bNpedaYFG4BwWHXvuQauQHVIa9c8N1HU+3HQURP2M1lWAiH2
dyjaQ2TtfN2J5XJ5G7d27ib+9IXV/4/tkUqRW4kiGLyYJFIYTsXobk8KJYjV
d2GW5sm8K6FBuaizfOyGtXKr7X7bSZqWOp98wNZVtWLKVkPmw4xTup7tIc/X
v+3oCfrml6tXgHNtf0ekKVkJhKga3jDczmTGgEM8pJ3uo7HbCuagGQFwFizB
xmJNzTbm56rYxsZUPYiN4CnEuxjLQpgdVcnZM85GA+cJfaLDsyuQwXTNvY6b
og83fMK3DCbjD8Zy4Dzw96NdVTFnCqaUVdRghllLmYkuiJTOMu4r09N2YveH
GfnxjRXGXvJuO7ZZazpUGkcehnGxTx8CP1kXtz1XzC2K882JLcHnID3IRJK0
ZF90ubi5CHdeQDbf1ozf1CO0+7W/2Jk3ajjkiU2v+q9LJfIoyvAjtWcupklh
jF+Ervp7NrS+839lojTirPqbAyhx6m4NyIKcNHIsG6WAgXKO2hEkAL6HelNX
NCwH1M/8rNx9j2GQTED0OY5t36xs2pEXPQKp/6lsNlKxvTB7NjOqwom60Fd6
HlfXaEln2AqusNPDcvQMzBWP2MW/sqicv0opdWVW/Rzjime2Uyc6aLvqfaWB
1XDakd1Tb0ZEoVcDCYPmwk6DLN/EddoSTHeQXM+H4pWXoZGJqJacXmrBFUGS
AssfIObH4oBUA1PofMw6CyHCXw5WB0FfjoL4g/peJl1YOnKVLi63Ddwh8WXE
oAvvqT0ad+Ud+olDz9oJwUA5uhaqVLvLULYrTcTTscbAwiZRu6iC29tcvdTz
nBVLfbmwhOs7MyZ8Kfig4HaLH/s3qAPXb1nMeqsepmX7u223FhP1Hs1ttf8h
6RvjKD29ud7gGuptXmdH8NgAQ9AnxWS+mdr5J9KhMufmxdfunqB+xjRaNV1O
lUTR18lXERLUX65QfXsgSHv78X4MET0k7Ra+Hio/9rGE8mhnqrRuc9IIrJ67
2IJ/20v34TGQuu8fbhoSw/t7NtmCJpOIzhazmm82UqiAkTodlNrDqH6Td57G
cE7mp/9pJvgdyeCo+RC797eQN96+ZUHwm2fRtbctJS8i6FQ22uOp3HzgZ0OS
KeMujLqFaNB8SLvPWRDo0PzP45at99x/v3BqK1gK1A4tT2Q6mvT7xAGWD0hn
y1iqMrbIXVWaZyulIbXjoBsIrzNvwuUdNHN3ouaXeGfaw9Op7KmYIrT0cntN
osNBIyGD5q2jSaslsRL1aSXhX7vjaVpRRrBF7unFqXqWvSolJBVHUM6hcDB4
0zsxf3Ycgr/FHr9CFdqjUuEhLqKpp4RPZqnB0r6B5aD6dxmEiU7Of39Hfp0M
9VwuvJOzr0G6u/4PMbzCWVAkjfFqvuJRhOZb7L5gqrFKvLq39tgteoGKwJ8X
7vUTSgiqabmUey1YRHP6l5wledP60uRXzzfOdNFCbixwUzERi43CFAfoAEhv
g8yX/64Z5HTVkMkI74kRQcI11PDA1P1V0Z17TF/JnJpBzbTFFn+psFMyRTbO
i/xSK67z36Vo9gMP71mKrb/k7AdISgORCtzqMZb2tk0vY0nbaoku5oG7ZpIX
keVF6HOejFRMDvBHNT4LEUH7Ox9QcEkBG06zKWndy/8XMpvpVCH+ELQmPjvO
Ynt8h6Hclj1vcenPxqEUAOSSjEHTEqA/9PXnqZWsdfKMfrQQ2lXn+hsvVGtl
Mgd/d2dDDjHazCakbRKH3iaNBvUfbH72HeJvMYmUglDr0l9bZa9SmqUHPrhF
gOdKEsq9vMs+0MB0rnj1PB4ucSPbMS3ylrA1qspaGej8QTJnLg48c4h5Eoyg
fJJ7Cu9s5qeFXAXgH8qcXGdgc4tHJE2mHXfHW8zSGOElD6OZMD57XCMfUy3z
h05qGM4qcWYgY+nGKtzkbXqTYv+qMlgiKcATvabTgc7fMpJp5b7UsZHqBx/l
5XsSeescdTiUoVa86Wg+HSbaTXILxf7XNNK9IOu2pBxGRPbOqa46+3LDu9iO
er9TUVtFJr+1qNlUATV8//EArv8YyMp/tTWOdeTeoBRMHboUp3k2cvUKvcNO
0hxgEJcJNKbJXX0BHXmgmr6Ibtzg69B+n2Nz/NWPuSjWmtYUuZdzAoGF/TVY
1LL3mYc/Am8xB9ljI82U5DstgW0jTjzrGLRBJ5vEQtugrr/fJHUfTmbHyitY
s8wQWhgw6Rda2gXuacF7BggRLg+s+2DIOzLryZ2bLEdbZGQ0wgPSfPQErw7E
0xEwJ0MNokeMRC8Ogzr22aKf9ZDlOyfYAWHudhsg5ZpSRKZReqopMiOd76iW
E0S+fWsyBhNDuMTvSeo6UccStJzTVVREG06R7UCg1AkikoI7yAMYMeat50wY
gcQZVHISAS1ozuUl2cIkjS0gDn30i8GJ8S2Xut//PlaXGZ6gGuROquXnxgz9
+Cl9hjAiHxuYpRsgeq/cfzXNG4hy1u+hAzSH45WgHp4IqsnRfXLpj+gNpj+z
GIGoeQWOeeK+ntSRQmmlZy8NYZolIxSquClFXHqcncfMqzjxQJeGJSmGrCj3
pntaTLu818NPYUSFYQCo4na0cP8rl/npNy4mU6q0qxFPqhCsxQsUJLqmTWYa
mV2NX7DQfNK6YWBifRB6lgoXLbPtwzwSup+qmvBigsWf0ifviLzvR7G1+Tyl
OG1Bmg5s3qugiH03Mpc48eMoKgeNvw0jLyT+X/dp28/qaFqqII/pbqRohB5O
JNKoj/alX4UI+3S1tXDUuX1jAjuKPwtylyieHnIRj14g2JdDR/VsHyYpf+4O
/0XjFFQW08Kx8MEuQSRMvQa+/FYQU1lsS5vgeAd2fQuuiTIaLgofZ0u0U9t8
ln+kLTmJUTIn6g4rx7owrrslCY9Bxnop8EtwFCAlB4VD+UiLT3CqDp1tjPBr
/7M216qd0TKAaR+CGsMF/WpTTwLDBeM1clBmD47FhutF/WARyZMq6z3E7Qcn
K7P8sNGw5sb9aT2Lt/csHNz/alssweMReYHaV1fflzGxE/aPqVW6WqQE7xto
1PYG45z5PNU7Aubvx/1WOoeRfjL6nkIatSSXtDJmzGJBgHkJnig1KMzqeb6h
jrXpfhz9/EMnmWzfQWDRN1S1VmY024Nfd4wKAsr+3qitC3htJglN7onhZE/K
PUoOPPDJeL63tniWP29jBlbmpbMvx2GM8MyxfAIi7oU1frwfvXrvN+5ASmUa
y0Dy0mDm8Ou7wDCvfSQsaiqCb+It4HAfczxKfbpcYAvP59d/VQCxvoESOmnb
Pne5ohTKr0gF0F9jQU6PYBrfmNR8qGv3MJmJPpkUzgDXJ+A28V4qQoFXnrLg
tm6YGY6nExdQyNQNHWw9tIi5tREu45MH1BJEK9hg4jJ1rqqagrTK4X2ys3mb
CclJuer7uT1yrViv1gI+p0b+DpGSKb5UIpxqawX/dDRTxy+a+c0mLjExrX7t
A9MUkTjqTa1yVBOqT9yXI1EKfwWhCEIx7HAU3uM8QOdPSVuCc6M+6TmS65gc
MVqgaB3jcEpPFFb1Wd9lMErnQXLho6T1yjvAaPJtPRXeoIzuhgrbs+63Ggdn
6nbTZdUwsT7XXMCnZupffdGeRYTqrOrZp14o/3mC7//zYsa0chGN9wBfQRCH
DJP0dYT56Rw5AiA4jl9tv6R85LEDvJgkkyOulNRSrBUc8v8a+K0tmaoMV0oy
qIwpjQYWfHsVcVlu2bfyDAUYxqscQqr+0QiJDA0XQR2ZQ5AduojF5h+sIqd2
xlHxboWIxY7qiV192EyNFkpfOQ2p1nwSkyxdXU28cfK7uOKkHOg59DICJx4m
yIpP1UKDykJuFTKd1wDG7KnDPzbY5AE03yINGXBTDC9vJP9CSkpcobh+xYtg
TPJePM6kTmHgmeqZJ/kp+zKHyhtpGzd+nHNkmtwmSq49HM52ylbx8fmR8r6A
BkW18yqxR9ogvlwtNwikXeCC6lB40grjfQ/qH7srFixpRkMTHHaRWEz1hr+t
WJjv+9Pg71POtIpZmmYCOnrDgaC5PTEK+L4XWoJvtk8kdvd+TEU5g+y5bWf1
64qKtMaJhdqIt7JlL7m5HdQ8AXYz+2oqYo/pT1C07rRqiChM6QXlmXMnQnX1
ScrnWAfPrdLvTI3m5nCvNhsNVz/FXvUVsQtBVW3P0gxmcSwlLzuJHuhDJlwQ
gaSUDZUU8+QTn9kdKvONWGOBmZt6CJcDK5/0Bta3WDkUqaV/iljRZxOG36+C
pxDpbXAA8mRcxyWZTVKY8ec77+hfAA5ZDI7RdImwrgjVgPl//D6+NciXFngU
PKSsD5WLfhzR5tm0DTq2sZCPNFBXaEISPjBeL0AYs37Rbonk52ky3uDCNlQG
3Kpcmks+AbFCmVPCcTXUcGx4Ma8aOBVhn6CcZ5bqIVQvLmOpeO6DtLez25RJ
7i4zjjIsG/QDAx+j3q/1nBKGS3Uh9uxxpGHlbeXUtpfBDJnl4MtPwu7DIUt9
5T+bfJeTuFIRrroGOTEYbWG1r2ziNp6xa3sQpmvfBXeCUpleuAA0fFSMcUxz
KXytiNWsflPGkKR4CbvIYWN0orhwg9RrrZcS4fBFDvfe/8PBU+UcjJPtc1XA
lz5rC+mp9mwxTnoNN6Y+Zl1X9KhWunyGKMnJ0uSx6vT9jRK58WCz207HNloY
mJj7C1aoM3ch8aekugQAHLfn4ERQ3TIilrRBtOW5pbdwj0lvlppi2cwDgeTq
dB0SeK4lwrU9q52kVOox3jtSRuFCup/YOqlAIMRDl9iKUHNGi8zhm1PlZVjl
ahptSNNKW0XcX5dJ8RPcFztvAHvTEFatwJEAzs98R5R2cBOsDYr5X9JI2E7m
QY8zggazJsFeg+vM1kbRSbJvYynO4UaFR4G5WDEpY5pMIaRmuybA/OGkz+7i
rMfzHi1cS/9KMY2+hjYCKSwzc0H16IRLNsfCsifcR9gqsDbhvQO3iIfrsM4f
DIq+nKykTIHLEMPUdq7bNG7YoQ10kWO52seudz3B49lzJdV7alQ/je5OPHBA
5xSCHNtTJ7aLwhqDiCR7k2wXKeMfhdyEqTw+YxtB8k284+05MsvfnRqvuFt7
gLEQC651cKQs7SaEMGT+vhNr2VfnLZXHAawC81fG+Bto/DmI1rQEwwqTa3gd
RiITRZN2xnRWkc/Qrfsc8gW4KoobYoLxcng5/vxdI62kxmeQSGataJEzMv1C
W7PRpaAU8kiBC6fG0Jy/dEMma+SVAXL/J+lptSAQxRfVzJBZW5UBTHjhrJ3Q
XtJf22+9NfWqhaX+GWIKypQmhQ0jLu6mBFEfS3IDCqKtgiHA3FjWE6F5DW6v
i44ud4AO0bIDsD9pYhcAxqZKIme1e6rk0Gd5dtfl+Y+CsC2HjCLxclSP0QpZ
RcIO6XisTCtCY49uui3iKZb9oMqWPFWzZ6CtATzZKTAOTY5mKQDwXcL3dn4Z
3ig+7UnUdYAxnVTcAjphhKO4us3dUfbJYAIAtEHhnzeOlWP3VWm1W9+4GnRj
e2bm+2O9Wy4mHJdAksToJU8xvZQU6Rv9Sl5hS1Rr8QlyxSRG8ad9MSmsrg5S
M4t3UyP3QKY62pkoewrvjh6/7PBe0oyUiPCmQL45ZiM0cA0zBNVT4ucwn5Bd
P0p5JfAQQKrzOR/+xBmjisuTtneITl+TLulpC3BJtEL06iHTTBFtUl7fJaBe
wHAj0+B1upjL9Lu4RUXdy+3uRDHmdRC4RlpxJUQcWOGn05MGYt+Jj0I/OlXd
PBNzgkhRFlMvjZQ7ZotvAWeTDxREekWCx4cMNZhVfMbUexG+QcvndAl+8ne3
0BOhK7XKT3qpvSmKsNJ6waVKaXjugFpztvdoLPy1UEkdvHdvHuEv7VJ3AuRM
6B5of4W0B8/Jg3EEadSSIQOwl685LH6PNyvoWimPURQUpesu+VTca2qkb0vk
HENb2bwvJI0vjYoXzgti5DrRyqf0BLkDsd0ouUiN76RN8bY553EqGEVroq4+
g9f0MMoEsUB9oAAQ1x4g/lhUyWZPgu5oEtRY6UoL1Es+4lVlaR3ehXdAjXqL
6mi2FlnADBPfD4BPGLNe6cVJI5UDOblo0dPmIHtS4YiOCNxZB15CU1WGwWfx
kj2FnjOWtNG6alDzSLlVTWx4m8KH4JQ6MI9EXEBMZB/0WWM8xpmq+a1qnBC3
wDHK0MqDyZWLBE6D7+LFpDruCf8qDsSAxG/I2cCaXWff06DuH1njL0rkcbLE
HkmKsjpTkNREgKI9xBSORkms6C7Pd+US8iN07ael8joLghRD4RrMNmH5tDIz
jab3WWsj+NvP/h6Vkp4JTFGaeboAzfpEfQNXhhs8mabRvFEpLDCUR4DMd4/8
/Bv8hnQ7MuRHhZlFqD7OAkbyfYbk6IgTXMZ3okuIflWk3Gp6ByZ4QbedRzkk
NUnmrgybD9q73LOtCoqYHnuw149+gLRHruEeKzzE6v3WFGCcyLnQNrxLm3HI
qi8TWq5iI/QKh+jkEF0dm5U1LplvWlTAwZljHuWxQFni+456LYHDL1m7vhVq
pkPuba9ocVWzvV0K/5NdMnhqfwFnu6JmKa6kr/21CsEy/Oq6eabTQvJy34Zd
Dak6naBulezFB1vtN/ON+tuP/6VZrMqVhMiu/NIkALPoCf2iH+3CT8yMDlYD
t4BwQpV33Si3PqCzoTZ8iuuzph9bkGMdeoKpP1nVO8b/aMWr1WcoD3TW5ZxZ
VDiFQ5t7VmAO+eAha2JqRJLJ1BI4bec3FZOBeHygXp4p39VdZKhWtOsnZAPe
5+6q7pA4xZdBPpBZOyclWZjuasnROGoXn4ywPSWduZW4/aB/9zb32kP3MDqs
9MF1wxdYvA7dJccazbPyPhDapVVkEpQrTcEvtClVTKjwsQvdg/yyCpXq9xbp
y21r6o4vVUDK4ntRbXhaPIlQk6F9YkGramep0o1lWy6/TfA0mauwD2uDGkTQ
dffwGYqDJyM4F0RoGwOQe/dwsHpZx1hHpY7TNS6FfxO6gwCadhlN4faETmhF
ggIYmccvXOuSSqTslnufjNGuoRF7doM4gAqueAjHdJuYag13r3omR6cmobaO
YjgskDxmCcvZAfYZ5JuBo5xZqZyN87aeBNukYpXY7atITdHgbHV7low3PiW7
OYk1jDHHb06sPrJj+juK8zHbrdS7uE1wWbfdQZ9hwGJsydPrFUIPFGlf1VJd
K0TDr651wQdJLjcvagImE6vENxj8tqekx37DVWTDc0vRBwWVlUBopKTZ76yE
Kk2DOmRGfkEhF0UIpT+tIBd1mHOTpL2/u2RXPPVYynDAOncqRCqOF+eRtky/
4mT03dtId5kp/UZT16UfpDElWotlbgC2+8ylaiCte3ea+zmd7l6z1/+LmvlT
GQOhPpkfS2mPHggQqNcwDeSZH5Zg0ac83Wq7ggpL6WGYL5yDgUfgklRTx09C
eMzY+/YabS6CGr9Svr/ZG+gylZ/xvqXzLDEquHxkReNGxeNbJZR2WoYq6wHz
MQ2JHDFz2FQDavFhGbUeiAC4ibgy6bb/xsI6eqycGJ/Qf6avPGjEat3VJfjl
ZVYQBRZXsONxG5oJLnSJ4fM2coLVtJs/Zto6+V6hI38FodhlAj6Nr+fLU1dh
R6Bfdy6DxRCprcvX0kLWiPZR0f+rW3uVeT7FPeVMSBhmqhJ1Uv6WxfxOIxLR
Vituj4TRDXWGwELmkRlH+hBH4Q2ORcG79rUu3am3pSI6exDycy/e3P6X5Kop
vWoy45O8McYHaYdsTQL94ewmyFhKESzJz8xSPRmjbNdSSv+O8bk1ur1sSlwq
thJyQ8NiUJwWfxFXayI3PHLjVfaWtoxFQs6AtdtnP0l50j++RXuRHmTLSdRU
KshKsmPDNXx81i1XtRdBEB7bsTCiuWhAssdvWTfQ1f5GdTmEu9uCyk1NEba5
//+jK2c8LTSeiY3cl465PZIOJEHi2SoXak4SOUgIQSkL59xhX5cDr+D3Zw7P
dEwnjCF/TQEYwgn+aqRER31l/UVX2c5pL8ygVMfQt+mH86/V81kqZIkk6KZx
qWUXyIuLNU1lT/SeDuwGoVWrQ17s3H29Fv9uP+qbejbmjNm7Ya93pLRKDWS4
zQ5bMrTchVqDxVWoVZJcvGB3cMHccS9sdkT9O1HBdA4Hz8r9Y6dn+03vXKnW
jAPHnlTZ7jjGaqbLOsGb+8IpCGqqGwrKS4UpXNOS1VNQMHyYzyZTNoGz4kRu
lRGSkxBNWT/k3WBFqkT9jjApOADMUeGeML8RT93pMxREHnksONlRr/Ekt3AP
wRr9jL/jHoOI83/0ijx/2KaGJodnnBjqZAoanOCa276l0G48XGIK0GyIvO5D
cK0eyzUCIbwK4WcBZaLpQ7qb4mo8Xb9M4em2VkFP2lh7cnHbZHhYL6YbyMzt
kxBfDf+2Vxu9z0LIS9WcqeqvkIBmtqEzqwhJQynUoEttJixZYBDa7CUpho7m
cHCSvWTydEhIFvo1BRxTYelkBYWEljsDJACxycFoXjlI8qQ2DgQJVm00K4CY
7zUs+WkW36LFEW0iQJAc47VKfaaa3ABOwiHXebW0TxvhdPurj/Oa0dFtd9qn
mxpunb/jkuQMR/ZOuawlANlYwqgHdtaNlAtkTWQIKoBeFrqWV340G+IMIPLB
ECd0GHlABrRdZBHwEfmofdtvQKE+pbTAEvbSvlPBGeiJ8W1Wpdk91Aq+rGXf
dU04/N6fJsP8UoUekAvqf+Kzbz5eMkSs71DM2s8GgEyNUpjH4XRKzvo5pU5W
DhVkRjdtx9wsgv3AS88LqGb/2cXLKZD0YqNjZH8wnDpPm51t16p6elgfYm90
79czaFxiNlu41I6kQ6NGtxB+4VNaWc5bopwCdetd+btermb46hafC9gOz9ho
Ij28fiHOHKrdER6TBlu77iFAsCuEcLQodhKyJ6HsCFDwBLVMlobR9Jxi+Qlw
R2LmZ+rbPcuKRH0miYGujHUBsiRf/UhDIYUQqM4KmYBsZtWaaIJeWi2H222D
pDAfY4P2aSf9WL3JnaWNCmu4CjxWZUaopLec53R8iLMuHePDZTpLOGDjv1B6
i04Yj0Q9D5C6faDBfo2S2fST+ELThHWuD3dEGapSXFuZgybk5cXF9Ks+STKf
RlWBIk7aZ+PCVBmpzHK6x+Q5Da0pAMQT9CMheDdIH+TkB2s38E3DFjfNqbzV
0XjZLh4E1UwmgRKu69M6QjI98QwomycRgceUz1mQ4EuUMXQaGVMKlnxgGumL
pHR0/bdcJRnNJZ71pLrSagB7Jw+tCW6FUtFt7RysOjVURxKsgAMQeI4Rq/Yu
4dFtwoNUubl4MXg+4Smo4Fm8tqlqW5w72QvAd92QL6yF+KVqEjwfbO1BYxoJ
MQP7ZmQLgl+JQyWdc2O9JfipLg4kvGEVIa1rfXSJXiUKX7tBnRlsJbejctVc
BnCX/fL/Bb7XRBUxaM4LtYTdty9zI/wS8jgEzvrG+JX8+NsYhlBVALHZt++B
v1Gm8o8s3PMx2nUS9BcK3WhQq+DqAZ3cu+CyeV4/11Pi7X+r1nprKw64gCIN
G7jjmWs0Oiw4yFtRhkhU9J34A0JUZXGABS2kwg4uA+g0Q/1e99Zagvl0S7Xv
t8yMMnUVJuly83WLsvbTXGqJu2i1XhsO22JWVzMs9Si+GwX9R72PhvLuYZhT
bRu1+DDPl7U5KPbXhZc6aCrR3imomfK7Nc82z+8a315ep2ASgS/JPmOU2LbX
alrh3d2Xq37BpGulAE2cAzpZ7iuj3tGcauJoP6YRsgfQKhK9m+z6ew7rDZzW
OELIXU7HebZyZj8RN9qZ/x/TZqJU7WrjIGvFZ0maQO/HHrW9+bn3wWzLADKF
3+JCnxDunDLYCbbsFv68aaQm4JGNG/SyCHw3c3Br2HElvJEwW7LFm2ZdsrDD
NWTzVoSjvyRr3NTcS4p3fZBhmgBqMElGnvKI3icvXr+eOEwtf1jD7CD08xXj
nbv/Be2y82pJuMCVxyOjCeNT4hho7asQYwx3yle7B3l5CTQMdprdOEoJPg+Q
xQztLGysY+mtWUOj/hDsrm6jJ6XTwsuDKSOrua8+rFfdOdVcdFXA6sUfgN4m
vATU4cAp9hpjxvHID2NSZ5wEAhwHmpFkss/YLVJOSubzTlFMRGB4rhj2Ippk
VMiSWHj+L5Annmty5httWiGHFxwT/xUOwnKUARkbNWeXtpzueAOvnRwyFPhT
o0JaenylhMvTOufkLjGYgodtp0Szvk83OMn7NlgsSyqHL8cUYOoAsWjdxamx
Kl3QuaIEPcouoKu4j6awzNllHrumRkPdcXCOMtLqPErdbudvRZzlrdcFCFyx
plSXOoz9Aw+aarVrBLmoZ1O+cuL4iKSQxh4WLhRnufs+9X+SwwrkOYLzC1so
AuYn1vEN5XJXaRWZTQPEhg8177s7EFGVtm8KPdQ2bRM4dTTSlR7PQggBAYP5
7nOzmtj7AWY1mc4BqA33MAv5DGjtX7e5qBoPWfgOf85G+GzuK2TFI6DMoQKM
sSJa8/GOk+1vVKNftw1AnVHAZ0355LGFHZm8OH06ZFa4Rx00Fmg3fW8TSJLJ
5OtRyNBKXIPTu5uPwCAzcgjsdCo5Kv4aYV3zr6gX5ZTGJEKiz4BaiGvi0ksl
2qmd8HezTT1wicwD/3uceyip+1aDZfaoi5Ospen8l2cF0n9i2MFO1l9d64/v
miiNShUzj9F+81NlxkJsNmZQUchmjAjIfxEJpuofL8SFNp2HtKI5JHhde6Vy
S2FtkuWWq8DW5be4fB6Gy6XKhAREKA8TK+ux+ot3mRbucB/casbxv1xJmuS4
AUUf4iNVNuliW4AdX3dBMg1ET5wLsF7+QyMjg+caP88d0DT9tHgLE38DZTTC
mT+JYOwnwPbVSz7jH3FVcC6tfiRpw2lhc5S+Iamb6t+WK9RYfZH4pku7qo+O
AGb/OcpBqjOUBKy3XQvdOJnDkVLZHVtdZSdlqJycOcZQrCm+GoeECdqDoIPw
ZYb0iU2B3YoiJ1j7qi9F+L+KebW6d7Hf5q5VB+s+zHIrZBTypFA8seJpBqNo
3Pb46Wp4RPgQ0sNr5VJQP9jp14ZMXYltuybeTR6FQzXNCIC37cqTmdq2jIL7
y5CD34P9tpGOFRV7iq0S3lwhq5G6GYEtk6d7KrFDJuGI0DxbtHEo9vMHAkcE
yj5tVhlwc1g4miPyvkgKBvwogIPiW+t/GZ4uNM4q0LJhEnpksa/nADgd51Qr
Qe0zSw9DckYHn+nVXiX7mFIJWznKLRBoWzBQ/2fb3AnUTIfmRHTT8g+J8yyn
rKokU4CsDHTM451WSwaKMOfxdIdO8rwRyUKwQ3+9D9HIDO5z7PkPFXQEtvJX
6awXqIuOFRCKHc+Ltc4ZJ1xitSx4hQYQS+tFE6u7KK/2hLS5FN0I5+GpHcFD
7mbDzIoC1j0L0WJmNLxwDlXD36iaWwthpvtGWvPl8l1OgW2339Zu9AJkB8iB
PU9C3YKWp1nEHjSR2e9R8ZeTYpDR+7x6kSBYxOZ2qoACJftRJEx90tf6rq7B
ID3Kur3SxEG4JekppVFuFry+m/mfZ7JfUI+anioArvcth9ZN3OWgKc6NJJ3N
ei7KNoH7kEQQVQsb0z9DpPaA37loP1TKFTNu28+1tsD+nTs5xYWKedCh0Nqp
5g4IM7uY9PkRRiQ4Y8tXyAu4+wMJ/iNRd+RhZ60vno6UKwXxjYBIdAWIrg3w
MPDXulmPqcjmRCFjlGQU3myFwtNTyrNru281Pe+kZMg3j9y+p+kMo4FZMttp
LQUnc6a4evtRZpfoBU2O1T/Kn3212X6dJ9bXCjLyHKXxz25zodBqiheTsXzy
kq9HywQ182pQcMBds9Mkci5UJIsZjs9pG03Nx+5PeO/0lIY8Hjs9/B3OuriT
/GVFIjU2e1rCq64qk6vqd6o1pE8Nk7LaKmPcrVNgwyxaxJXA7F2Q2fKH1jUK
IWlRSWaTStcn1N4utB2lQb8/AcXuD9C0bxLCPYMMmX76cahptCm6kfPLaFJ2
NnzXgMYZD5d+HkuiaULf332BryBI7RJQYB1qvhGMcU+Q/RscDjUD1aV7AggY
aLGFxPIFt5OKvMVuD+8hIlGNrIqHzvO3yP2KJOkSf65XCNN8GzvGW4OgallM
AUjnQC0BLFEXL+XsRV2vLWNW8+kcu5VXUcwSZOrrC3AlnHcHltN48rp26848
ZVTG35n8txBYCpH0HWQjJhCqmXw3bM76tHSzWzr8dqej/5HJ7qLkFDzwcmZ1
a1aOmLqhq0Jq56MIw3vglj9TiO4Uvf+yV29SaStmql/yPuBIgBQvCTJfBYTD
aCRbj3Z7Pvg5fu8zNoalG16uA+gN0xbdHgnrNewLlJFYVMnMN+V2jq3lXlAX
Wxxt+SKarvdOOqQPu6zsPpON+PiRu8sW8RhMzY/7916O6EJDkODwWbf28QYa
rwy6lJIHprlRVU7dIXH3T/Aq5UxLxbe41cbXxlv2VwTQkos/s4suJ3gUphYa
LwAuMnK38aQ+V/OvBuuu41U3/9BVKsxpLhaI70MT7Uq63Yx9pIFATpfAXPMN
+guRErqLOVoXlx1BYReyBS0bAa5kC0gh3t/SWfF3gFGkw5fJKE1Khoo3bA4t
9DMKurCS9WmZqFXtqC5oyoDgFl7aUa48x/FMIIO07iDvzOu5a8SzPrjDvuqW
z+eBWVqxBSeKcCV/+9/pVgU0TPjJJrpql9tW86JnYevw42jtFqOqTPuBYEiE
1n6v5d1DbmcNwFSWtNVPQExlGc5m/I8AMfhwYoEx3H8jttljwXIZl47oKuwa
dDTgpDCjxr9YkNhEx/v3WplLjcEDxKcD+0q40TXf+nbrvCA1eY3h3VYlLcJS
VyNikzPUbS1Kd1SDTJnlTXFZ5I0cl72h/XrDulaoIpUxjWOaZTpJxfKCDz5j
b8XEWNQH2ObCVj+V9bx/ksYMgbuYCX652EtNRCSg+8Dzv/geRMU21PlBiSv7
xYoyEuqRzjzhz/T7Kb5yEgOm0wuX28t3/fvs8yQRZO8H8xHkX9SaJk/UeoMy
Uw8lseXGJvTnGFvZCWHpz9Xvel6hlfkDjrkEt3IL/vxYdK5AbCZ+FhPnmuFv
CIJJz8W3Eh5atrJxJhVxaY4lwJLpksApVbZPVh9R8krKS+Lhl9ulTCHVVa4B
MWpkvAFdQzJhdWEUGV2Mz2AvJPL5bLWxbQ0TZcpv7L0pls/GPGiC0VrPvqxU
nYXlf08zdpYEmK2wsy5us68DEVxgWSeT3Z7qowX44PovLkzAlfBoRCLWPWZ4
feR4dqhu9xnlVucbDMHM331JBJRUimnl57TvarJR+dGCnAzCvf2o7W97Z+h1
UJhxqKBfiGc4urT2ojhiLs+pprtVOPCO7fr0bKxt1uAsnoemoZnleCYeFN/k
iNnKqLo2TPAcbFZH4ngNbFvBltcWytaMLIOhDwqpVuQBP2Mr+LIUW2cK7oIQ
wZlpLM1+dDhiudS8qclSY2AWN/VMan991Q/D9scT8K8b5TMs7QAquTvC9v4u
FKNczeXXUzuHelRCbwpAhyMTgHs1k4ybkymxYlvbZHYhLUOngOatq+Lppqs7
JRZ9M0Vrw7sXA6eTmjvzCqJtiFIgfsqpvly0T7LjmFaOBWdb6lMPsuhChPa8
/g+UI+qI5xYfcm55vHojbWcalrt47YstIn7qiWJml4D019G+n3okDxElX+wo
pxI3XKphHxhblN60RxC5azYvtyjEmqLe66p2prmHlCQ0TF9S5KU0M+thNbQ6
sJLS8Nn8ZFp7TZQSL3FY5G2142t73eUlw5tfFXuspZwK4rexzcuWJ/2sTbrC
x9jLUA+pHBJ34dv9cBVQArUJtL/vQWI7ukcw7QzZhA/SSr3hhjx59MxpdSGA
EOz4Tt1qk4pQlhpDYB/pXymiJH/aOpQ3mYFC0yjlb+at5c1Uth36ABP0GcK8
RAFwi269nDbZtL6VEJsgYhOqUcUtsadFXQa0jH9VSzwvwxBDgq84bLrNVA0e
SUbJ6f+I3Ohd2H7NtGC5MAoP/QOZP/fJ88+cn0Spwktgmh5N7b8hCzg77UWS
czTAknM4/Z+tB6/OFhDK2x93dqcTt4TrzCdFP+jAv941jQNj9XfVeLmvsMI7
dhIggjxDYdMHAar6jIG7h6WdlxgY//ePDHhCPTXHD0+Ass2aBDWoBuXGVLDz
l61QXBBadJzvNfL2ILZzLYuBDYyUKX9fd/a5wg9n7qkB36jIpwgVhBDwph7L
SZDTrjnIk92GzCC6KROtWDmAlV0Bj/lgSo37G0BVf4UIiO1NJ3P/dPNicB7r
Djemc/jUujVXz6FAO/FUctuewv0ryh5KoFT1OahOpc09AeDktn4e1zWbry4O
CahxrwvL3QI/E1LMzLWKptJyRbmEkyvwbmOUkkEHwlvv/8hfaQIrUXoez+rT
6jATjiTMCX7Pgmpr0X6E11DiPjGTdQAJqvi9o+bdn6WbDx41oIgAgJo8f3lT
FpLeuYzfkYyADBxui+CpTU2GLDoxmtnfBOIiGLz6l44nQ0t4HBAJqfew7PnS
7wdF1hQCXkPz6rx4noEdYSW3epogDuVo6tDzwiaBHVQjwLxd9gQ6L+bamD8D
T7CzdEr6eF0BFAYHs5Cqtm783WMgWHs2sn7bp2AdkKBMeFx18xat8PFoBgW3
mF3kn/e/rgaXP6DqgREyk0uOCfSappgo3UUUJm517DJ9B1q+duCa0dmLWT/W
+577X9erIaSPThyyzt3bfa4Gc8bCY9N1YNXBiUj2zrwvU4mcN2hKFOa2cPBw
shmDvfT6gbBe5G2DPCp4JiTGAxpUaWpXcuWO/E2CT9I41RBTqY/08zWp/Seu
eIHGy5JgTDo6yeRAHdu6pf7soj58t1U+b7CTIWP13222GNSwGx9ThTAymuHg
70HRUnXdhtiMxF/AIJaUBCc8J6cG4YC5SkY8gacurBzn97pVi+pia2OLZ1u3
wMluQVNWoIVZYnE1LxxKyyBrklRaWlYzcgy7dXq1laELvaHSaAbNQHMI3lGp
EnfW2nrpsDF88O/BlUScCMQK1c0X82RPcAEzNHLqQgmEY7gIvhvuNxydFonk
KgHI/4RnN7MHxyiBt1R6f2mppG4OENeBBiBXy5jYL/rJXphzUYoKW9nXH9T1
FRRDJGulSMK+Zh6LUxDfixzRlEd/Ny1QW5pm2jq87o5driutTA6YzWdX2GpQ
Djsjh8S2xmrVPDyDOMt3PicqJfJsMfm+X07cSiRI8hqlsrUjJ45H7EdaqXbN
mSrTESAecYO0la7GIDlkCJl7pNO7+6iqnOEEzRL/W8xnQBmZSuPHwJR88/wd
cGjR4uLAYy6exzbkmPp7n7FBr95qnUNPhfPNWKVeOCY8eH97NbeWJDZJEGus
1LnlpXKX05BMsnHgmnzReU+gqAqCGuApwXQrBRLYOadz79VStZOkQZnPomMz
09PM33eLumiJwaNEI0J2bLZqXYAe/k1Mb7nvUy7yPcon2p59OG+Br3sC5tem
rByd5s3d9a0XCkBAOVeiawDsZfYOWv0zxVrD8JiM9PIr7Pg5ogbBB5oqRd1D
kvsZ9IXrRiCVlu3UHbS/FzArEyd9AUlVBZFdR5BhHRvufFQOHwggkogrRsnq
+lxKJzRSXQLX/hUWmx52fmY0sifawAZkHzOdrCTAJnuGHyycfwVC/YS/MPa/
/XkBlwNA0mUNgJMOeEonuxQCwTrvZSqvV3MAVi0xk+Ws9olbLvyoHs3VP6i7
19a3UrA6ZsTTC4228euC2P8nXcwhmgU12fPpbdgy4/gCZdtaTvvRTICKaDAu
IoONAbZE/WxNzWj65B2UpBlqvL2A7mOM9ml4dQw8UqBPmsMWH7I8sxWlu45Z
ejhEzV0Xnv1xe6X1jxdVXntR9gB9eXEw9G8SQpquWANtepuI5BhtkLZXB+v2
r+AfU2jZjqNnvVlsKV5Y9orrZtdp6c1I3siZXgNDxUxRFwX5XqMbB2D2JVJf
FOv4/lM3AbIZpjltvlbs1JDi9t06X9uERdk9b2YjfNjFQ1yKvebKRFapzG2/
sXvm47dCLRMAmxoLEKs3iYt8yqm7ltFS3WVz2yC5qPPmZ9AAxz4QXlGHDt3D
+bmkMp4ACpD87ZGT9sUemwe/0TrFBk8Kc4zZO2dP6dgHjjvkFwr06K8BptXl
OqY849JKJGc6C/2oTsESaysOReuJccMgcnhcEbdhB4Ts+hLmmOmtg9SqykKT
WUPwJfUwTwFg29KaNz3ReqY9LSwH8C0MDyl8SAtYESekxWu2+kbhuQw3BFVR
GhQy7pANdr6Ba3NwS3eA6fdi2UgBl02amAvu51KvJhjm7V7JKHa8xsgq4vqe
iqIX/JWaD3muWJpe1fv8YppsVvGZ1yFH4B31pM/JXHUDIwBd35oYpHg7ptjR
c3Mtye/5ZUU2MgFikQRddinZfVN7nCMn7rOsOJRtx4LLwI5sVtJ7yyuo/oeJ
SolEy9B0yGKISpZVtArW+bSf+cwlhyZ6PlAphN1+NnzJpnZHTv5WfNWOmdsg
I+R/rMxZ+bwmkg3LWX+rph7PaKAxVGXbL4s5qvewevY38/DfVSoWfSdf0Dpj
Pq6nCTl+YF81jHxKuLtWYg4esSsqDclLcR0YQbmCfxvTaPUd27PfjPQql2RM
eKCH8UYleoufLCUIyWAbNC55WMbcY5Dw92xpuTd2JWscr68gt7MchFucwNWy
GHwqh8nnY85MWPuVX6J4t9nBV26UKzx71mkHtQ3IDd38T7zs844zQU9rhbjZ
iGbstwOkGsz+uiiHl1vEZ/cpWTC8ndTUvJxxjQKt65FNym/+qFw920EgzwCQ
DnSeBF7cHQC6ndGzrKapjSrPuGIySE1RTOktMk6DaFYKku/SoL4vZyJb6i5/
VCs+9s9o0GX7KGZNITapsjO85xBnQ5qrYYalHxLzGGLXc7/PQN8G2AzN15zC
1Wr1ss6pWJ+qoVYEaX6xXG71jDMFAIshHsOthHONTku5PC50yiVwGlYlwcpi
J+IIlrCEAteOdbQ247ehT3lY+NBkv416c/mAwk1Sh4xHVvokPfdeHxH3Zfdo
X+MLP/RTidyO5ro+5DO1/2VeEiZ/pk8UsWFH5uFOxvhfIlj5PYgeee5buHl9
TBKnsqKU9B01y3CzqCUcjyHyZgYqK9qeIV+gDqySZ/gOfosv/o1ZXJe42Zpb
c0xlB4cCPjjbqz0UXSBC0knG86A7Kfv69ROxKkgIAkJaBRy/tRfDPXDXxvqK
IpkvpD1KmFgnQAckimptiWHNNszmSfIFA0bMBkgc7gxGRKA7JCO5YdcR+umT
ZDEpA9FyH/DQpL76N5gdvrFT4BCo16sO3EoaUuRhYVtZqxPcwO6hrnNZoPBz
U74WCtFbp1CN6mHE4QBG32Nbi9EbrhaRjXJo7xsFbF66jTRh1dpobtrA9A9n
VOd3ix7b1dVA2ql0f6ih48xAgK5MkVt7UqLYTtrGXEOkJRmUVfNdOjaw7ygM
wUkLWE5M9Vya6GBYm8r1c0Ko093bVg4PaYT8cx2Wnvx3ns0+x74KiRSmTSYv
9Goo943AiWERbRyYvLGvIaQz8biYX67wQ+XUj6qd8liOOB3LI79TzMRzvZ1a
KGq+DbVV/tTzeiKGOPtA0wvuShMywDXsjYxi5qvYrhr4DiW61x1t2oITwJLQ
oNtGy+JDkt5HaMZd3CqXJz98xrEvFWMx+surARjYb3XP/fxjvaDPD23yCbkm
xuh55RBaU24HjbOl7j7TjJy4qP5ajujN2sRzlOzsdojPfJEdn8E6vxPMWiOn
8weCALeiFp+jUOPAMQvlPKONSek3FEMYFu2fwp0jFyRqU+bC4nN+7eFP1SSn
0yBSPLo1McjnqC0upQMvQgOGyaqx4Fko0peVsROqESMSSosRyqoiSQx2WXt5
dInchNtY+V+nheanzMwlKU8aKFlCVpT6pkLHfESADGHnYEsVXaUJ4v3kXYBZ
U1w2kOLMCMo8TGf5cK7qaAsLDBax2nqNh3VfFCRFwMuK+phZm6h2FIr50b+A
yOFTuEhjo15H/d0d55dKV6cS5QSNsdfunt7Nj/MLYZa7TsCKA55eeIzhtROz
/g26+D3LixCkwCzFPvuYf6qNmv0PQqEwxIAVEAkrfrglnUSqR1XNNjbB95c3
9MJL+ew5s5yeok3AKO5qtaFh093j09Njel2C+6zQCMbMEqYDb08ue7lf1RPF
dGrxApzX/AuGIDyzk1MqIiPJxhEyz1h2e7+Z3vGMFhd2i23kVD7jHphqNRwY
aNDVdvH/Z5pcnv22Cg0cs2RreG2+hqJvpx8lqW+dMbMm0QML8iK91UD8bFYt
3q+H+/PtJxZ1KNv/M4t06hQfuSTUNk4Hx85vWKIkAnV31reUAyqT9OGq2KIQ
p5xIBlwR2uiEDR8mHCHegA8JBXgyzCePNvIaCIMp8gisHR86ExwzX1jE8R8f
3EbDfDc6U5YMq5AsEZ3wCDzqvJerHyqA73qux9m+fzOMns/xFXZ9HbE5/T80
ohQ+2wXwhszBxh7PSBzm7wcrC+rPKwTsZ1QOFg9Tl0goi3QJkcrDDmR78mhr
771EaVU/y60Qfwj2d3mh0I+OgdkAcbSKbPNClqxcZZs1scNFv60iofKygqyC
HgFVpBcRb8+MgV20Da9gv0KrrAPMzyea2Ugg3eY7CAZbcOYfxZAjyGsWZDGk
OA+GapiIOkEsw7TId4iKAUoZs2jK61XCExBjr442MUliLPbGRBtvk0cU6xIy
+BKQMpvft72GEbI82jX09bz40WnZA6FSZ+Y2Nghj7ZlNX70phQMdVjF/Xkc8
rHybe6djWyckvZVw7HmFZHeCgWYKGy7r/ZSXkEdP7d+qjqic9LA75bkcJCB9
heg8xyyWgmPLCLOpSZrYK0avFDqQAlnrClT+XGYfAuwsz+9NByR4ynxELy3l
NDc1Lq8bEvIefk3+HHTRQVVd+W8pF3LWBdTS61T2Q91J4Sh/1cgue1j/k983
YjJiFxcRKaZCI31JBw3Se8JxxyQaZVOEd8FIxbLhQb0NsOIwBCefrCte2oiP
fWFM7oA+d+gOmonSw7AoFPh1I/310FYmkUFQTTKawjPNz4cTK/JH1qL/IsXf
wWLDlfk9lQxeYFxIyJfCPguW8jRw1T/uPWEYdqAHhg4vI8XICpjYUwjTKO/0
NZvmkYNr9Tj/am9VphkplD8tWWWRvyiKchZNRgUtCE0iEHFZ0tOy4P98HhYI
18nqyeNM0/Q3PVlonGYihl3uNrDnWkeIplx73VsjbLGuziLPaQKQ+FpS6SwE
Tsap+vw56wM3uYsia8Sk/b1sgpgaKvnJ8STrxbJ582YY3+kNLwpspnd4+2Jb
kxDjq0hQzWdTAFeN+OpqGeP+jbMouuzZ0aYHvMZnmLxwqRmKhlT90NG1DN7n
oG9HntO57o3uz/6cYV5td1Fm88qGenWcHHn6k0rmCeEbO2q/0SVRtIz5EBmR
5Rtt483sj+083z56tLUWBH2aI2n2ik7MRPuwA25KYuoj5yL1hTrjRIl0GAYk
Pb3DnMj5SEe0AyBKhseOtZek77I3SDgWRkYuGkS8y8luRGFeeLF4eJe0Y57o
JMv1TZe1Pj034evDvs4ukqIPFItt8rA+DroFeZk0VU8r5iUSVTKZ279gGekV
vV9gNshmBfgdDoA+N6VvEyUfm/8MlDJdO04kVSOKaTFJDu48/FKg7cKG/VHT
xkt4KjekJNwrz2+Vdynd6tksJJQP2YATK0j4rylfYC/wbryE+iSZQkDDQEpg
aQFWng/Z9ZnEUC+LUV3Wam2CDKAaV4/kfmUMUx+Vf7qMdxbQKSe1I7Te+YGI
pMwKbXTZLFRDrISS/7JsImaO0v0D9gboDm5/4gtAceVrCUUlwOyuJPKVMA5m
LwwEp/ycTiOdbe1Dptk7Qj32MHTy2rdUoXd5WjJqZT7N8mg08aII6AmpvzrG
jxuo8xDVXq3iWw8U3rjg1ZPeaGc1F68MYZaxN7v6E0IykmkiNAUJG5vCED9d
z9W+HMmUMMH9a+YdtbGK1qI7ukESo2LiEkSd2+SEI3yiA1wiYyHjI48BcS7n
Stie5j8QdiwU+a6x5G0kzbhbTX/tzU0DRWofSsjhFijzhthxbV42/btp3U/0
hvxUThF+bRhjx4PCDlxStPEpLKGriXq/pyNkthhCYmdAslIqVMRcmdU/CNDh
eFN94TMqXHZQqzFf/IEqNV4BaDR/LyJxGW/b0RciH9G/gXJD+idjRT06G+Uy
lUYKc7ZxYq9UtJTfqwRKlPXdqlpVISoX4YPKk5pShOLHfnUKSYxgkJbYH5SS
ZQaABomeHKLDva2ihWXTnc93rr3D8inULtJOtHcqFhEDnHwSfOqWPIUWVYrf
rYJ1xCFIsl2di0T+DR9oOK3uxQCrPA0j3uhDrxUwopsrhyXgJyw5V+MPX5F9
VAzMYk/ahn9XMlhOFtJ5FZlozYyQFvGt7FgVHjt6OLBCTTUnwCabVE5nuT9B
aDwL25Mq9eiF1iFVMY/WUZn2+k5OBFpoPvmcbAVJ9hkwV1FBigy1xQdR5ssF
w012APLUKXtK3cKUUwkWKEpf3ID5+45EIlF4ZGNR/xsgZpVcaN4MAnr4Byn7
N48aI4qLf2KjDltu6pduoNcWnQc6DtcL9Z+QbgWw3gjm/u+VKVgf/E6BlT5s
dE30K+iz7lBSe/v7qDTzwKI0E9sd3kNSE5tdNSf4Cmvkm5xSfARWupSLcFuq
v9xFEeQgnCupIhmUfp/SPbg95gsDMpj2QuNkhS6gjmfOJ86W4NC1m1N6tYJJ
jNAMP/o8vh8/5J2xR8EgApHBeFYZhzxKRY45idr9GcaemDU9GGrbtcymX2nL
fuXv/PbSXmA+RgLv+KbIIq0pEIyTvVFpb0jgEYR0k1SuOFu3TxORMjR3hx+a
mfFtHcwCNaX5xTU/XjqWyhPGI47IL/D7OdfPbJelCqMaPAu62QYgjlj0s+Vw
0/vjJghfLLUf1N2MpEBlKKV3PQC+OV2bwf/AQ92EdBE+EQwMZPrpJhT+jZQS
+4xoyHj5/bYPtQ9bl5HFSUqTW+6E0ITjWCP8Jk/MfH2BkkLphRmXGqsxvXw1
UrWV+gpqi8R2mDkDiX7TAWQZJF5M5bkL5HaidL+KudIGBqLw1lVPh155+pzH
bbY7BtHR9odP6xdeiQ8ToYzTqj3HedD9wkM29gbMqL0lpD0zKomW85k5lP8k
ate9CAZPeCF3J5hSv1j9AmeCfetCjXxP+lebRviZuPjWasfOcPHG1YVHRDZb
mQcu5wigiCc/8mrNhYRxKWGrZMFxGvEJRLZ441sVxj0y3/RZmuF9tycPQaB5
MR5JfQudT5l9MZ293eIRqbsGxXx8VYZICQbK6Na2sgWxVgp1kAflNvcgIRVW
YjXv8FKyMHBPkqQokTZHMiY+4LXOBvLF1eCrqoaYG68gav8XQQ9o5hPnM5Lw
E81A2CaVnuknoa/6O9ap6BqU8hZiqUJseS381FU695b7xgGS3ujvZTokIGiv
Ca0WhYd/bH4aspfcGxCBxATHamEyIUY743lGNoCS1U0lSYwZGAHqiAVyxkgL
42mB90Q4oywf7YckVvHLg9WnBBhRXF72d5NdB2FC/ooJZ4R6pMKYhDX3A/QL
uTKeWBKJwNUFExOlgYbH6fS5ZqJTKksnPlUnRaQHsoFS63PFBsjmrVPzZRqR
b4kSq9uco9s8oJCnobwl/vHOReyKy3PSSlzv2s3KNdZAlvwz/5M/XVxumwzx
0ph0Uc90wji9miZZmH0JtDru/3TWkVpOOg0Ual0wbJ9H+yPvthAr70Q9r960
TJeuBLZDz2FuAPw7xSJq4J4ekM0nIiVM3GS2n12jKqUsEo4y1KbnrqEUxeua
djwFVSEkhzJc5/YlzEkscnWcWARTtDICnDmOXD3XlxfWoAR0913nqfvBtkK5
cQYQR9owmf78rfg9hIgOLe5vxGXs2t7IcR6nPCLBMMrB4mViSExTIQiOwOpb
/g5walRsOTkywyX0RCbwCiJSfFPZDI+xzvTLxWBzAMNqCQ5VeUb0e6Xt9Za3
617aVABbAG3FxCYAbOIq0hlH18rlGb2EfmEu/cer5mxWI7JDMK7SXB1zlA9S
+qQINFJxQdOAdQQ176mRgdYoy/hZhyQBy3ojrEymhvZPW1oGq8iuCIcJCivM
k9X8ZmwZKGlKks/Hi8i3L8rkGjkLNokH43TYQeYTaIxPmFIVctQnptUkNm0Z
LLz0D4hWq0dTVu2d0WLFRvS6Zps9VCDXHR4ImFokipMljnYRG2MtWaaY2bu5
VTOApiwRtEYUFUebQzamWbxeWJwmivDVqNwcedSfN4ZX+lvxSsdota37q64q
CQduFiBAg85oywYX2LsS9i1KGVlNyJRGPVI0o9LMPDSyudNPWo4BXix9nRAO
O3gx2sxJQtf+OqQP9bvGp4N8BqhwnscHmaBPyuAkT3lWOmnAsnoMdJDQQbgN
wTgAFgJUsNANu0cpI3Hv1sAeAqklTk3DhsvN+Yr3Fj8+XBGZJMxrnnLF3hPv
85NgxHkrQynGi7wiBijb18mBE9S9dgBRFDhRNY85RLm818af3atwtIsFoP8k
Dw9iaarCRCG5n8pZAPI3f5nkjYdmUog/v2B6jt9Kp6We4E6Vhpnau1ITNvZX
We4UO3b9Rad+ZVZMxUp9JYvYblvojnLrH51TW14QLiBYlMmABsHjGXqwDuwX
WQTtTLDNysg6mkeyFAQl5vkcTrBgWr2EPaZvx1MQEP2YaETcPKLIgME+uJUp
FqlwlXD/1qsKJTTIbmsIEjaP1GibjMAbxj8e+y5CR6xIy3/Td0KYVTIdKtr/
WDklL1xqNQZlPiUcnS2UQdPw5kNCAfZBSurQeFzdUvYuNZEx5K80vSN4fy8e
O0xlHtkZqjtCY/o6YQIMwQRuCQ+hR+ddpqKrw0PFZOFAkubjMkQpamena7yx
lERicpJvlOTJHVLiIoHDCRwtY8OcB6wThIEJqpUWWsvMTGq98EsZfqHZT/r7
QFMOBpOLVTS0SGFn4lROKUr0kHk8520iAKF0HyC4tazwnS8b9ufqW1WfUkqn
IpujSPlQISuktlFKYbvMG7nPoXFXC0dMaz09cGOnnNUhnQbBA5DtSZah17Ql
0FuKWyDLyZcMpMD3fpLe/6+nwu0p00CVh1DCBgstP5ctOLYYbq4/YkksrLaC
ixnC7eN8mXroJhReKo24Ly3gBNk0JR/Wvga+tyQgrR76LVbmCG630tdJI/sg
JKx6DEH+FSvVw1onxBA2b2a0iNZLtEtX8lXDsU1OkS0zBNT4BfEi2Yc9lHm6
qEvEikjA3APsjivGepfiffvgn4yl5OHRJ/UJ1xqR71UyMRLEN5SFN97VSktI
VNV5ZknJ6H9kD7lpT4GFn64Wx2BcJT2k+NAbr3KF7Z4AyZIbG/XbBzsY7AEp
Q0VnFXFmlNTW3WDBWokLjc+D6Cuv105yMG8rNUdcK5iysD/M5MKHnbHxutJb
g8QU2lILxLT4rSKdxWEWYAbQCLl0ERHnmty6LMmQLOePoKz4otSSej6dQAlT
BdenBPVEpL1YK/pW8UF8syRWsaLoEj6pD/E3Eh0eibqN6f3zTuIVMt9EawJn
6K8h6oQDuXgZdseKobHLD1GuO65JwvTUiPv3QnyR4JzD263g/c6h4yDeCKA3
x6XxFqSKkUGT+Ds0T4eWbDM95NsSlMkZmZa9HD2hvNMwpO2Jo0D+9CQ0gg1z
qdGAbhc2k9fqP/dPz3rnXCcJwTCsgqOM3LA37vduL0TeGy6WemjY1F35coCj
uIIr/eX3cn0XAEgzmQiSh7/2L49iGaxos4cy8jDHTBPmuBOkXAnYgtHQ5VeZ
5WTfU0I4FWq7BREQzYKJdZ2VMeiYm9BE/zgdYoLom8Y3a4QiP1/XapaOcDkK
qX++mSSoLwIgv7sgA8QBPqR5p/C4sg3fO4oKAiLS7rJvgxB3ENS/555Q/w0b
KycziayJW4JVF63DUwwyjQ5vpKRI27DEaiiu/JkXC4sTR/BVIhBwkpY+lG2Y
7C7DjHNcInZ6XNniMRPkahgSS8sxNc0X1xvhhyMIgzFpVSC+/homOU0WzFuj
SJrpK1BChJsWZZGJJ4G/fnpA1VT5rIzDxd7WdVtubZGhckLaMoK78qVJAF21
brOan7xkIA8Ns/FFvezt/44OoMIKGh42N+4l9pUr9OkfJOU5H8slg8r5F8X7
qm9Cmd/qzq2Dx5lqHL3fSXS2XUGQGg0og0z+wkwyrKhRbRHFcf/jijqFSjwc
aVRxRlZfZVLrNZdI2TrLXxiFd/z5b9YVbh58WV2t1Odh62RP+54N9nTYNpxA
SAHONbfH22nXUa7sfn91Ln+l+4SkrlDFV8L+K7ld8a5kgGn6OKBRhjmpF+Dx
9gQ6GNqTWYccu1GLyd8njvSK+22C0gFB24s3Ow51AJ0RCMiC35AU+cpC3dke
6+a+T+ua57L22At+fzkSQbia8nrqg3dyXuSUCYzvzJvVYYG3xlUJKunzXxwH
RwDcIplihOj473dWbzuIiNAiDbMLPuAYznNpyzketPqf3bktduFVh4BTYgbl
96UBnRz7Xo/yi7/65uvf7xpq0K0Ot3i4iOtR87JqGCRpY7FVXrDrkOIWuye+
spx2GqrzVK4kzYf/NEycHzELZBt6Hfcphn55ci8Y5AM9pBgJxgvyVX48EJgU
kZf0JKbgz3TcJ2D+Ye4N+CllFoBtPaM5ql47CDte/n3UAyA4qrXfDgBhMBff
sWmVKGfFABtuZ+jrLO3/ZGJyaRe4L8CK2iP0AtAJ8rR2nzhW43KmiQ9jNC3/
Q3zWEhyew2LRIJUdZnxdpRMQ/VaW163k6NT2OlTiIKTBGniQFtT4ABYZLFvV
E7kbLg8pRNGzXSv7P3ljLoNjQOnRy5KUvN3Y9Szi25RyMczo9DrCgsX7qz9s
3qQf/TETH/QM6q/4QwbOnJDAopLHrTvzA/DTjYI7Oy16WyQuLK5d77IioodM
aEY8Tz6hM/ADmCdMzFJjQJd7PJA3bwM55DITNgsESL5z7oplrqPvdICfH+KE
tsfjOtV7qK0czgQR2Hv+toq3iXAJEOJy+u4z3FznDVhpDEfmXBdD5fdvo3jE
ez5o2Wo3j+r7+PeDYH6JzFShjlJjQ+IZOg6GJiccv9M/8BLt5Fwf4HrHfS2U
ikEb6//7OVRycSYTqhR2SGEwoq4HvvCPZXJwxxe8H481BFmhACyH4n4KScwg
KLrIYA8+L6bXDxBTOKUzMFXDfRZM9I6dXP/5MLiJEdiET9h+7brGxdo7Dtnh
0lkuS4M0p4+QMKukrRxWlKuqq371E7cseCk3TgdF5Zw9gylOwTs2fx0PCm4l
3D+naZjbkN43RKARSAaaeUaAskcZr7CH1zklYb49Q7epw5jmZjO+C4lFf9tM
ZLr/kxp+m3TYCuiJ/I8wZn92dc/01mUF0SlXRJlk1P5lOnU5YCDTBnyLtL3Z
8ZQJG8cXz+Ldia1B/ifuLQWVbZOPbZ65muTEHsvfGx8tv+iYB8JgVdk4DKAP
hcJ/QWIu0boP0T4c9P/EqqmugasChDmxoDdmjMHDXamZqSgB1166EiuU2xVT
MfvNJC9V3mZgAJaP4Zb6U48Ty/y9olnRhWtjCRhDXH/A/I+w7VyC6myaeRxn
RVF8exYIIE4GkTKipl7YuD9+ILm0IWXDd2YaDbCfRWuQgiwcD5ygkAmTveM1
W9k8zs7AlagVHIO0YILedw1vM5z1C1I009a2PABre/gaBaVSoyyGxMsfNre3
ECjWnLUu17TYvxkS+Un8nsZRKm08G5UQZwLqG4aowif7ZRwLMTue5qUY1nyo
oCOpvJ+A80gTY7SuRHiKmFvzImsxY7W95CYwy7cv14pq0ptZXUASf266sqYh
4+qSQDEaytcUvFCxwnDhLdVdVQN7nHR6xbi3JO9DWjsyXwCuM4t7POGSs4DA
NTl+79IkrTodsTIFB8k/t6jQ4VRudRmFcDgbI+ipr9mdH6ewwiznG8vXs5ea
BYZP3vURcZIhzRwlEncwbjBUJBf/00NQQ9mnr/13p0tU7IoOJq6zW6/0I5Km
zsJBozUatPD8n9Js1CS36f+iwnbdue3Z43pS2FPjnWQwx8QANq6MNns6AaYR
X5MoWrchcN2Hl7D1nO/+gvhtr94T1aBm1ZoBBqk8npdTavIMxiE9S04f3EZO
onlTqcAX/xmFa9gsD5CSFKwYjz5wSMgspGmhvsq1XiLcC0fk3PDfLBC4tTSd
QlTXYrfIjBR7OWhCeoNLkNV6kVUxcAoQEm8gkVSyQo6dl302MwUukEY1NEfR
uvKS8erAv0OqM0+Y/UBmx+Wczu7QP21RfO6urC9HFlnFVTJebTpcBOMNno+U
gutmL/SZNzIvIQZunXti/5WQjs1CqHW9IbVthvc/z4EL//MUgvWnPVYN53MO
VoSJE0i1EUXONeKpcY8S+pTGBOYG+HSHhIKgwYtVDWdUBQR2nJW03xRE5JbK
Dtsg+np8/Fa4Dy8KFC4wXOvvSG8FJKIYX3hdC9gCuMxOtpPec92/gmzjRqqH
5wX/7RcwhQDd5jEPyrCqczfsCPGZx1ZmzYRobtBKRLk/Z2U3BkWuN0lPQuzk
4nkVrgKaI3aB9Iw6kgO2zn0fwVFNL8RokZcxQ5uXlGN2iDlL1CKUfqeUtaFY
44vcFejPqlROGasV9hJoXEOYCztDosa07hzrf3R+P1qxvBvVQoxMAElrn1dZ
eWZvfw7oEM7t7Zk+AaEC0sNFoSPykWw4EjUL7mVvOlMMyl+nSgH2dJBjTmp1
Fq3mgJZmQX06gRIX8tthTPGuzw/GqNVDyFaop3wsJoBKw391gW4R69Cv62re
upQf8xtPhv/OajlOSecRYkJ9EOyPkmYyeYfCvULnn1qgbW6Kc1ZmcGOuLrEn
TYSAu7hSI0CufQR4vqmK2dcmiDdpFrZJXl84My4dGebYJDe/itPeIbAvCEwh
dqsLUFRKQHSItEg6LpVUbsoceP0C/EuCseGbuwFFetvs1O1sYFKS8c4p37hK
j0qcUJhdRsuWuuNMJxN8SdC4oaeElsW1oFfXF6bmLBgcPI9mRbPMEbX9qpqw
sNzuQz2q04KaBPm11vWp2D43slSir2QgIuI8z80HfbtXx48C+LjYszpoOEOA
/7ITbFJIARoI9X6peP5RHBwMbiuV02b1i/y3Awp1fp5I3/aE0NtWT62FsSk3
Zz3BXoq+RmbNLwEaIkvf1F4CYQEtORfuKwXmLuiuNMgKthbc3eE2BboEacVh
jNuewvoeA1GB4La8/eKaoA+h90KGUwOWkloF0n3yISOCvsO0qzQsIJxqo3Uu
NTgcg7/wcqxl+DlFIQ+dyTxIFGAINkRIP/MJHu7+9/CY+AYGE5lGPDVxVaON
fXndB88k+v3nIePqD+E9u7WLhdrdyt1cobcJ0wfMJwyctrRmr+JJ50e6TGfG
TA5UWWUerLpIwAEu8amELCF/8ZdVDJ3rteF38Dh7AGb/fqym4PZcvpdQJyvx
MQlJSRkQ6bWfrJCFH8l+nHp7756qHIB9sUe9uPOo75IS71okgZllhwobGkca
jeoGCvyLrmBJSndruzO7Vd6bLf3A4DKtRgQy2u13X0MD7EB9SSeu7k6NY+YB
XpfuRlGpsS3mRkXRqLtVcIo9/oqSY00SXeEz56OnoYyKt7IVMVXBZvLNsZHQ
o8m/W0cIoL3ck/rzeMP2Hf4Dn73QLvLid5hNfnFn5eWyCpRz3Qbj8T3OOtNf
lt3CwjF1fURc6J8rMwKdgK7ye8I053R/TAvGnovzDxocl+ojcjVgh/OXnBTg
W2jh0UctdkWnj50N8Ld6EnvODMWQKscWitVznSziSGir/nkNCkvzOMtW7pYN
YVgn7QRh4qS2aCyajCrMifMS6JL8zDoCNTaAg12+/Lzjp/vXx6/bPKtPq1xh
kT4W4s+URp+wxEO/Y3XJLNEOqoD2pIvYCArQwrZnfs1R5meC/Lui7vyygXh8
rAyHr7JXI6Exjm9+1idvgAbiv70laVl3mGcoc0qDuAMY21/K2WQDVfi9qjax
Zgrqd6vQqky44LTEpdMV4pZgH2h5eHV6Ov6hhz1twwId/pBjQtKFhAPZgsOy
7jv1EEMz+DEr6M0BpZdcS97kOMg2onskuBugdCBqVdleLY7aP9lPew2DyJS0
ch71tHo82LhWNldhRYZQg6k+BKWe33ETvKDPhn0+CDJQbbBAcRRz6UR1G5LA
+lYBx/tYoHnv/DSnZpswclge3LsUNmsnsMoeAk7JB2+6x+5w/XaRjCYec0xi
yDhLp14zFomE0ZmR85ZC2IkkuFGormaRgMdAsNFpZ0938juOKPXgN6xos2KQ
ibn5Uo2A5PPy7VxOsFI0JWI7j5eSzWvZyQ0EmZW2Yl3fgc3UrrAuJCMKmofj
4aey7MHVPlQLL8XbIne4yJg1H2RAQb9eFfVGqSdoOItCMuzYyFglkrJ7Vg1o
naWTb2cJE6RlqWPAbpQYmq8e5cSAwE9LZ6LfPfPnuhRlviNWO3QR5Qs7d1kJ
CCPdH0vb5628cp34IewS14W9kNZFaYHffczl44E12SKmcQ+IwlqneS61Xl4e
LS1R0JKKD9yLYSaGpxE0qcYpV541D7OJj1Sl5GIhCbGdJqBpmGyO5K1gK6c7
k7SyNtdJvBXDZl5XynCcpzlYwXJOwxQ8GLORyyBNbknSUb5gSiZnJN4l2hhc
r8q24DgIN092UCG2K63AJsDlEw6fTZNYaBP1Ua5LrgnubXKFSkSoGvtQ41HK
cUDhU6hwDZrEyV8AnhuG9piS5K19llRAffdNpVTThJ3KOC+SUKYQVCho/usD
JoURrQ29HTgxP6A+ddNOFx1KnPZ25a1lWuCbEiHX8DyVw9pGzBnTGhrROg3o
QBIV+CkXdULCFaJrGKIz1D/6ONc/BfuqEaYArlBZtoD3l98wOIHr88DPLcT4
0gIMS6hRdTW1Uz1eGIFSSA0owGzwv6+zn8FlRnTWpUoKmgsfLo9ozz5IkFDx
Q4ivDUi47xA8Ip6vuA/cTl7FREpRaieSQIizgFiSOD4XMEnmh/4tSfan3lDF
YR6xzfnqbBhc3iQ9piqbMDyb9GwmH5H6WF17tjpVSn5LYcqYou9sxJgqG92B
4QeMVoIdtxd0zTC2M39NOnjqBnK7nNEr20tWw4CeRLqKLQsEpzZI9FZMEtG9
egTbVQZrzVesqZRhuBcZRpbQ2gf2cRbdpSeZmgxqY8FtgbBNUEKnBYw3I1AM
WRoRvLIJ8yfXPjna3rVQe20S9HmPzaGLh4hxZRB2xqmlYHVqycZjptFMKopt
zVGhDGKIibepnLSjcJrOp3CxRrTdlwgBWS6hrm04fHDPl5vp0CQHm0RwK5Wo
LdEx7W52PmhYsxoXPkgWZCZQz3btQoh2yhWMKcoa+bNecxbuCHm6Ut1U5yWx
07i898dDvQyDsHTvtQ7PZNR8uc+xr7CsRwzdQT51VKrW3E+J8OooTur8Sy5D
sWbUZP2Xf/Ca6FDg9+8FhzlvafaNOrVoKiKmwNLXBhX5R1CqOzyJ3zJU3a+F
OTC7SsdbcoyjGIY1ynvdURhfkkk70+vzK49AzgGJjxW9UwrmfiUlZdxqErja
MH5BpumLzgDuALrkzbtWfjyV0hKXgc9Vsa2XopMpdRuL77G5mWzxWHis7UJQ
pmbfTfJvVxu73dxtiZiEy9ZWB0/RoYbrK+coBFeUIVBrTndHwBu7wZIzRALj
s5OlBi1kJgS3pStKTz30PONNEZ8XccU98I0cPiUSjf0ISos2+DpL5hhS0Url
I6eJ4xnOWA10uvSi+LJwi9FS5Z7YljnIEJkLLz1oFO6AYobEaeJ4+hETAtyM
Rq/q1fYKpeOwG4iiTHWPBl7VXr2jlMPBdmnDmf6T90aZX0qyxXnUrTDJ4Py5
Io93GWueG4C0H4fs2uERrG89Nx++8h15Qse+5FGC123ECOcsdWlwGB2/KHrm
sXj11NKSlaiQOVB5Lhm0gebyuAJDEVkvmNCjleFliolsbADW8EFQ67UzPNIX
5pyOqm3y9jrfyVj+Na6y0LD4Lxj/dwRnUVmQcZhGcG/P8FSjLbBWOrCnNEZ7
x/J+KgTb09w6sGKMbjdbxTtmta7/K1VhSA6R7YLdSi/Vyik4h/MS770R4ayD
jhkNju084K4mLU1t/tTbLucUrJ1Jtb8K9wGgls+tWpwsvO7n9oMllb0EJEbi
fGqrZhMjTw4Z9fpaec7UT/rSGMeVS1P2taECdJIA5JXHBLYYE/33ig0HuBcc
Q8FvIp8iSzKbw7rkdKQR7Shf5PoB28K/WkNPt+6Xk4X3JpEk2/wGQMU39f0L
iBoiQ75iX6QTk3GZNsFT+BaGSEa7L/p/0mp3YWJD9gvAKxoZhhO7N0C1mUTN
xbxnsul6zZfSvk/QzWLBtPItR1nfR4oSTyHeongxhVOgLAIEJ5TTYRd67hIa
2YqI7dtcuHVh5BuLKoHPk68ebSWvJsmj5wg/u1x824tCMCQdAjE00qeDHtjW
deH2R0PaolJ14GQaXszTsn78EnW0yOquEnOShxh9GuydI5yBOr9arZS0nk0w
SzBX0wJVBRHhSu8a39f60zODyFsfEO6zrFDsStw9bcVi8pno0YYYNmhT49NF
i2t6SyJwSxFGhB+/TKlC2oOfr7w91mS0vWnk0oJkSOHLCxigRnCTdh8+aA8w
HEmO5vr48D/fdqcjTUKz9ihA00j7ulTmoeXFvRDPwQb5dHU5xB/J7ZGHz30Y
GnFuHa0lcjrH6V5L9WMrWlI6XrP3yvApfQn8Ib+K5Owz8F+igeZFwWjm5zo7
inlrZ1p5wRfcTbrCJXixdLOKSdIMPlVEaC6MJXlPr7hp352ZIM4iNIx17IEv
9OXMdC/cWkOCV4IRjftVIbVJSLsARukNynkmXVri6nZpdXAhzhqd1rhFdYZs
qAjoqKee7zO/lARCJumk4mTKTqdJ8MLyYxvDN77qgWRgnvn2RCnHvfXQQZEH
oaAmdcKIQHLh6xq3arlMM6YzHACOk/jXhYDoa5tk3smn6KZT/TtC9vKLw+74
xcphwZGX/M/D84Suc5nhKGdm5O+V8EziVwx/IAAPG/5yOthBtGeTo0I8/fMs
PFHv/PWnzMG2Elfqmjl1nwd1QXJESqey3fpsTpwhW7fccqtiQ+uNF7M+TtJA
YSM9bHkVv+Ph5bLyIREXcpVv0U/nH/J3CodWPleJo6qtGYjUAQev6bFHp2xM
h+hncgEq30dSBOGSMlRitL9bKEEBR5nLvjidEeGZz6JwLqRV9W5gHA8n3T57
2Awl1L0NeXWIOG7GpLUBEuii4YZLYcvNQKLzfzOp+TTuhaOuD0m1zwHo5Mgh
PxRHcU9/3zJjiJQhalpy/QaTmnhn3JpCVbhKUCthojGcbbgMpLmu2iNDo9OO
hK4o/JZS+fGe6n01XzwvL+IXTQOk1RaI0kypq1HM5fccu7LugLIU2dWYwh8Z
jDtaZdCU+DWXqcKiasiaK5W2KoEYxUA4BPteZ2gu4LgWhXMJyTKJhyzxvleN
cC8XAgHK09+qws8ZC/ON4dEqBJ+A3jhHpJUoCjBytD4hV/Swzmjja7cIEKps
MmHxIze20GZkXBBQnod0BzAN1PhfaDlWZQeeC1de1VKleTfR8EVAYPiBtPJc
PtEJ4Bu0lul0g7SCnhDTtU7IICzkfJPIhg23BwEE+TngFJRFfp357LgxR8nC
5IuPCjQvbJk7U8rjk2c+J4WijX763haa36enEftyqOGqBcxsQ0CmqsmXUaGG
R4C7T3+rzXUbaicoONaOIOaf5btXVpSrYHkCgEUuxb7BSoCl83TTsrCFsNca
5zhDPO/8/2RsggwlBFnbje9O/CrOxucvLA80nW8JPZqkp/R5zYkh8zChbciX
eXgB5MYUC4LkUyA1Ffv7zHL/y5ODKrnJsa87Qsf3gJl/YsI1c/YN2725U1Ex
oXMQxqSL3iULcsMK8IZEUwm9S8xhmWbJSFfkbHJaOMmjAIlnpQbSiCEjWu8i
Gm4N9psIp9Jc7PYqobuh23JYWmcbtuCi6GTU5hxOxVMOD7q3XOZOdXAGWRjK
tHK1JDPWrhPpvJHXf3Jkd06dG4/0u4zIJvRqhltnXv04/VnVih816qp7QJcu
mfvlP08B7UBSc0wstHRDQ7X9c/S0bjc/TTgOE84qkNti31IxxdFFJQkDXQdN
1cAznTi0sEkJ1b3PBF5psKtJpgo5M60ujJM7FCM8RoktMZQit9UtIhU2Ah4Z
RoU6EplGgaZ2NNt6BUhCpiN0dK1qLIM7ZfK9paRUFWlJYdwqS5QKpGeU3bXQ
znQeHy7Z0EkSEj5CWXKZ4+ch8dgQQ2B4Ha/6dS9BvqLcCjOIjIcMFIXpdOwX
ZOcfPHOts+oFIJGqosQtVsZhVFVhyIKcZ4i4K8zy2ZYJB75sN26hGLkAnScO
cXzvflgN/z95O/2jMIEf58TZ1aZXYSqze36QTtTzuDjMc0m+G9/scV8+Z3f2
ly+cnehGU2PgV5DmlxB1k0KbpkkzepyWa9UPJy8j816/k15YmQtWVxysxTOy
EaZZsg2i3J9FL7CdaNQP56nIYlm1vITtHBd0G6w9E55teZMlWvVJDziXue/F
enLGAWT5Vb5zYur0r6+YFnt52dhY8qfhxNqFkl5IWMtyab/h0wib92NICUT/
f65+qEi+LDEP6riqt0feYzo067oJmhORe1auATn5sq4cf2l71m+Izg5Mvg5d
pCJCdZ87u6DG6Lasfps8topP7UjfDAwQ3UEhqzhMSPGH4fV7moUe+7/150QW
+qtLPM0MLGqaHUB/vEU0JWvGC33SoD/3QZxOzRi53HcA4LvE67833i2n1ggD
PPJhaX6WP+f2CoxzXBlo2JASIF9vYApNzeUNtnwbKzXZ7Wxb25di1YQJ8mu4
G1oZBoKVPsdVLXtZ6WOBfIu3DR0LZSF/Mp8tI6IPQ0mxSB/cxdo+S3NVfuPq
A2ospavlQ5Dogy//K3/ObHaFzN+cpk1gLDlu70b1q/vISlr3b5qjpPjbR271
pXFbsThPZvbF+4Gtid6FN13pl7Uec5xisZhdCBoLUnQIsZlhQPWZOE6MjBvG
30xZbE0QQcRI3Ro6jU4yS/rScJYjwgcEc5Zr6RPo88N0VFO81J2r5SS3KEgv
4qa1QWlPtGKVE3KTn4dNmaSU6EAp1Hwb2ocxMMXGat23bqoOJZcoeXoD4VTg
MqZXQPJhB3Usc+5lP6iNhhBJBZ2tV3ryQGImi9GbWAx8ex7voJGqjG5fl/VY
0edMzK5UUaOt6nxOUYn+mXezL0Evpn4BXAK1dZEhTLwL0JxkPnLXvWCH+lB6
TPA9NXqtRYwPPaqFLTaSaCfsuFvZfbjGmG54XHrJ9GFSBmuCg9jJJw/9wdiS
gxHTJ4CndZ6QUdVN/dpxUouG6SQp3d4XWvfihIGINFtY7Kzi4Rjp6NNpcOjG
+Zbv4NDxsD5n+PpjsolgKo2QgI306ld0nW1McgiHJuc9sVaEGuh09+jVXxfp
yVVlHGBw7sRmjoaun5S4d+ASWCVX7FzwDHFN0gBYDmIV3X4VoONSljb+xDgB
sjJ2vw+w6I0QHJqa8yrpSbRyObWzytWuK/pfCaIdq8NAqnmhbHXmBV772isV
Pv+BQ6Q8Y1q3YMU7kaWBWlOUfRxvXGvQfDE/YLttrNwE2OxWoxyzsmOb7kxv
u3rqj37XTCptwUQHkhS9RFH0w+8TDu1NfaGNaO/gG19Js9/NAXHTDFTam5VG
uaZKzyeejXmNKSlnPw2x+rsBnrkYfsmR36tDhNn2TYL+gbkeVMfv+uwgQfjH
NxkxQjs/nDBHRROq7egdA8Eweog/WcWBNePQy63vahbv3N9ACu0uyRiXlrSG
6kTKSRlYzrYhXQOQkISqHWO6lJNafG1qh5dmfIirLTEYalEZ7Fc/LxBgJxMW
KkT4QB52c9tfICoCw6qFx2YoKhOjWQy+QwtCThSiFibB1XfgCj30JMb9FJ2H
MLKaxpT0YzUgrRgjn/a1ZRpaM2XBcQybNXVitNa6+rROc2Jdv83dWIYNXEFr
ANu5Vf3I/h9xWU6Dge4MUIC8TPesdROlMtt8O921LH73G7HTI4/9x6ZA2i1O
7/odO2H/Vis1oXqDkM/QtLrdL4dmGmq0a91/t9mcyaUnzH0JNRZBiDup778x
Mspl3Djy2fEgclKZn94ioTALVcZuZWbrJkQz5UvIy+V24CuxA+vRCoA7jtCw
QodmCx1B/M4VkCd6s56GOu+nbZxVWVlwMjYoZzB4mum6AL3zlliFbjlYiB0L
RPmEq8PB3RzTI2klOR45H5LePYN+d8JOFf7dTZ1iYSMnkvzFF1bj0wZxGpGr
DGd6v/O5fyDgknOE9QoIPaUu9davK/2+OkBhthPTaJQ6rHxkYyVpd5UMgryb
jZuKa5LQC3UdHIyMTEu4Hwek+OdBkPIENyjWlLOCTY3dQAzE0r+bQITo75Rk
7SvQ36dkku52lmNTekktKwQTqmdP4SbjU8i7GUtgrpcUIljb+WSSlcNrMSra
I3bxvuZyNSaNAIfF2oGSNl853vebobJ5BYj6z3l61AE39TtIFsNHXKGWwb3o
WFTlK/Lv/Wtp3mlmHSpG4B3rebbY+GL8T1nzITm2g8+u/FGJj714GYkmpfse
X65EmTOixlVfymxRqk7UkZF8+ZvhWx9lRm1gCu/nWo+AsCiP6OOAeynj9U9p
GwSApO0PNFz43DK3YP1rG58QCpvVeVkxZ26JXeexSRk2arn0LrusGKVR0cwr
jbfVpZNyHjAytLfAYPqED23p3lDhMsTYrNtC/1qd189E0lBFcvHNgKfPBqgk
Pzj4b0vuZy/L4cE1Sr7Z5RBOXlEy2DWzfSaq/NcL+pDV3yDtGX2juwq5WvZS
KhKWh6qsv2cKmE/FVjTmzrTRuOmngavRt8Cz6rbvNOVuJACQWbLGSMWqKQxo
MIr66d8uHeMLvGKVucQoK8xnSvgkN1/jBdLU/yihX9kavwPY+zkU4yCtOwq6
4NvJOjaBqCcbHutYmatbTGVqbvClzas47c5BXAib3D3btgxW85bK/hHgy/x4
kEVNtp13GFGHVF9BzjXKLnmEqnkrs2FxrB9lN7bCyqFv6y5iD85SgcJLqHCp
kO+owfJ1oSescjhHtR3TEPeO68J7qBNUaQfV82wb00FvmZx0IgtpIMGxJ8Zo
diaTo6KR6+IufDhtr4zU8onyPOl92ElXH+XhczpG84aBP1jJCwrwCtPvxFKQ
qVXTI8d9NP6bX4FXB6m8SUhCFWxdBdd2uHlZqfRyob+8SWtrvW1EdmTtj62H
1hCsdsX7OIE3nb5m+B47izIJs4/8M2QiI245Dmd04kEPy8fCZsmwT06PWt5e
9cMuLIHgwrrFnTXcndvR5fHsWCFXFcYHR9/AahQyOlEq9IoLdSG3KiBa2IUa
HJW9EReWD2qgHpqQadJK0rce56Kr+WqZclB8eezKZK761811yH9UaT5AyQIg
4t9bT41SDNK0seXEvYGAIJYsdjgeUIu194xTrf24aCaKmZr8UzhM4o7gTL/7
Uo4AfzW+zPXqvnYVpEHGvyvjtJOjUafbxN7qRi4bL4PyXgXHWpi0TzRbWGCi
9s3HyLp9a5BMsUr98wRz8WqafjXxwtvWnHQeZEQ4uC7yJHUIyr5xG0mkkodP
Vk+5HEvwmeewBtZkj+0FBiDndZ+G/fucF/yTg5+YG/k9bE6r0kUQMmlCq2Vb
JVbu8Z8uW3VyZxLKpgyJAetAyyu/jycLazhs6+cNLwEHPvi/LA7TrDMkBvrV
p6DHNNFOkB6jZ2j9qmnLiKdQywssLLtF0FlbiqfvootOYshHGuPEN9oFPA4a
HtjTQCr+MW6aP6fwhgAsNdyveG4EPr3YxHjD+xQMR5hizzK329LVY0diUECq
YM4z9RSQgvT/17TbX5vFM6pHpQ9Wc1l/z2WQQuKS+LQObGD50BbPIcIetlzU
X3a3UAjt7EBMf1hL2sDqzMBv06GUlzR53fXPtd67db4tsAKgyGSzxI91MIlE
Qt8eS2XI5zcdfFTsX2QBleGD1AH4lEpC5/ABrIpbG64Y/ZZf2GCJd8ihLKZO
vWLdjRQKnEMV5B/L0mo//8K1mgl8VV5HC29U2eJ/v6HDyLVINKS5KpGE/7PL
ETvSk19PkxUHE+RpmbY6B7HUNlXie0ckWOKAClWzat5nkmt4lEgSqdzIfigg
wRjkw+z4p5Iaqh0MzsHaBSlmv8cCoj6GW0Ye0hfRSKoAYli8NBPZK35ZpWHT
91nPgf90KrejtAQ5sVSKtZwiHWsa+iRjghpnW6oPpPjFm1rlmWZ02UQiok5D
ZT2EllCoyoEZ6New0bKqFWdSn4OnRlEoZeRAvd8XRXkuyW9ElPLLneMGFBPR
YWvumdsocuqPNnWj4qsMyOeMDX+HdYZ/NbzRHIN/QIj919+qQDAmXycG4EvI
c1hRIQoBcQxI1+1Xe+aqobrbh/Z/g7/1/FfKTiKpw0wozCkyIFaMw1E3zrlt
TNP8CxEwsWSXg8Fw66x0LgFF+/XHuVoJEEAF6+vIkT3Ne3Zkns4Ner9UjQQv
CRHA7UhwNvf2MDsuELDUiLFaXopcYSKQ6nSN2dAf0SoLWAZ/Xrn9bPAjndNK
Sx+HsJ7MP/vEm0FuHT76HunU7xLPRFshsTZYBzFMSlrjuldayKAkZz/0vb7F
lxhyVctSHJpxKeLHh1w7EefCBCd+8hJWx9zeFAVdixh0Kw3ggZ0XGhHoryt0
hHWxhQjU/dlWwkuFBNIhBAgEFmaxWJSgPLCTq69kSrCA0+mvusEMTk3vglyA
FApsbOoOQBp0LR2xZVLH3e+hRzgSEwBdC9i6n9o1D+rm1fgPZdN52eqnzU45
pxP6C+i/vkBGrgf3GN2VrN6tvTKFlzeB2AMrppZ4+qyv3m5UxgjCR/AP3BNp
RNms8j5YDDXV7BHjMNgXpl7isLddYXaWijTYlK+51LrIK0KmRxbJ+HKBy8lw
By7k7k/MKt+q4o3vRCZnk8Jjti5MizT+/59zhd55cpjDNM8AoTKFvhZrUB6D
z/zWoFRvvBT6FirpNgCx8hP86RUomSPNXyLnme7WQnD6rtBWAwjhDX8jX0m8
OcMQP3rrR21UCDUBUJ7JJny9TwLdue2i0hOqW9ckP1lj55vig9r540h8DinW
RD6wLZIOuVbrTM4AgXXgX+K0vxQHwDMOd0t1goOEKZHEuRGTBgneqygy47mq
gJcMdGRLA9zhDP+CtQ7qa9ZkgMRpNDqFtCFkYf3PpNB4/8qoMGEETcSBM57Q
eyYc3/r06jOsYmxvm2nIkI66PKfXK2SHHqObk4wWZwyMpTa0ZAhmRahDABHB
kg37scj/V3Wg685Nc7njxGPtuK+3iL4tJUyV4gJnHWPwzJ4BPAb5eHsHC6To
JwbYNxkJDBnjt+r9FtvmVXR7mOxrGWm48icnETYFX4q2yWDJXiIFanQx1ubH
3z1tEGazlPQGdkw0YFiyIKlVIRDsHeM/mqeM5C3v8OUoO731ZHQxvgh1vdgt
59lhoOYOvHKT66QbqY6MYQje1+xOkNPF8pt1pylWSr7cO5qndJyrsceaCacW
9B2k1g1h9pwb3jjjAfFCFgWNnpzLfEXLi/W7MpgTvxLHUmr25ofcLJG2qJaz
Tbr+8XotIzPzrXd+bB9FXrGmuI196GutJic4bim+Int7GZMxQpkanfv/o506
8bGtXmquuGngmFXAu2rogmA6udR2ZykmOXaZRsd9xZdifSL3x0FnduQPFLvF
X5lEzBDZ6kOPbvguoO4rMYHpWch9Z5DfaHbbHaZgHNYodHwYz7Lj5MYVfaJ9
6KdYb+HtpNp30nXIIetrCWx6fzj4nW9jOxZ9R/cNhysQJMGFEaCrxRhZaFi9
QvXwz1C/GuS2qQjXpYdhciga6RWZ+pWdKxKo76WrkxOTUAvM0VYbPvIaTVxa
F+P2+KWmU+uzV20SXeXXoMK6/N0AkTHmiNLaKowSTF6UZ59nN0b2VFbYBRUT
PSgdFJo6cBrtqKJfNHMc2eCgjZ/b6H0YwBQ1tehOwS7dbpA+vU+riP/g7+It
Ex5lscmpKY+eRajoT67DxBdyg7Kgbuvzc2qTHbvMOwFMWVqwnQIUX1qrYeC5
CIR8Jd6bwni0bJVgCWDjBLhfv1GcGnjUybFY8kstegMRfkjWoNpCZwd99OWC
zWXAkRJdScXH6GXD4dPdx7R/YZsyrwju9vS1Anp3hBCeLuAesX9ibEAQQAu8
afbXFKhXYjTjE7oyWnRMD0lrc1pl6OCyUCkjhwGkLaJ1D80mve87pJgyROsA
vhR5chf3+EIftMGxbDxxbsvgYO4j19YJS+f0rueWChysjcqmn4kt1gm1knil
m3VmBA+UgMlwiW25EdWaf8tf5KPHuUXO0T9zMnQZuch92AU4xFWqC4k7u7cE
JvcVzu7Uga88OUF3RQxvrQlnaZpTZr2LEBQ7dhjov7NH21ghp+XD1042i+1m
8Yl+lHPVL0glls5lNem33G3IRP8yEnqQZ86B6vs5FueoGn8fZfnzmXrCfbv5
fuaGPrxmAv+vtcpsVFFcMJE4CEscfd9m9Mgs0t0BI5lz62upaZDNHHO0JCxK
8Kn5qzyM77Q5XaBwOBOPlb3jpgUK0iMTm2NPeG5Au10nEyyNIbD4/0y6+kvm
+eBsIib3lvwlpxDKEaqeT4R5sUWOwMI09q5yp0Xjhx5r2YaDt3w0G+1GnKGl
+q+alV1PiBcpHofr1XGoAeXcVrxvwMLDOBjAZ4GZEvb1wiXT82fafc6cyCLu
zSvnnEUoSGbotXBkqYTaaNsdkjMhuA9rILtXZ4eEaLEmTZSGMSLA2QLWQyzi
NummuScJarly+N6hOlxMowkWo/T7f8Anr2EkftJ9kaX3/1hFd/rggK364HHA
uRnjGIJsd4P6Q71o2HVikEugOkvmIQszhcxKAjhSp4pkouPaSXcUfo4vmhUU
OXt/n/MEzMCGh0fc4OxinhLSL394Wi7100YKJWolofl31N3gN4yc0f4BUY/v
7FHj6ZNt/5BFhV0wJX+Z/8g0FpWfWBPs9lW2LC+QbfhaVbEBfrbGX3oWOMcZ
eevGUKT4OyR+eMyTjuHZ4+2tHHBFrjfaIWTFEeOYrcQqZryqjOGFFI6RzUb7
iaNAOVgPdhiuor3hW/3XRJeusAzsBMYgfaHDd2mmZ5Fkysm8WYQR1zuxfTHN
9XgWC738d9BeCIiRjgegW4pUp+O9kkbijsFirjfAnYVlv8p+ixJ3U2+VfHqz
diSImDiMNiYQkOomUjF62ZxUbbPKJWlshgjMd24mwkc4hC2ZQWs8hbbYdmQK
cgQN70HWoEc/7+wD/zSpecp+T78LLFoI9Uyi0GUC7PZM1JwS0i+n0Mff2C7u
yV3LJjsq+rvdWN8cWsu9fMVw8HIJdu1DfYjFB2THkxv6tWyiWgYjgff7umrJ
p/3ULVUK2n2Kondoy9UKdvivmnX6ZvvS69a3b7CRTByDlKFuqVd/kCAh/6+u
LHRGGewr6HnJyG/CJcIJWtaZysP8Gta9FyBeocbH5C/YqOB6TCTb5p39Fljz
hnIPg1M1J77EEVx91bXJ8M/IXJATZM/eLK8oojO/ay30eTd8u9wfUAgyemcU
O1BpmwxYNJMuNhFt8v1vvZsarOJMKHfP9kCz2o8ncZLy1NhFpXfCMShhMOLR
CeHh9y/qbcur0gJksgtojdPpRrZcdkKtGhV0nH7/ZdNW16zPBzyGEzKBZ9Nv
arvVcwq5HRsI+146nZNUBAIB88xFxaZPrK+A22UQQLwpyzg73gSuzuZ99Gi9
YqGhxlKEPJLqK2V4prHDVa/gJGSfNmrr8QEYp7iU+yPFejWYd6VQrcUhpIHK
ooT8DWWYqy18BSKYw+9InZmduzjZxp57kXuUOC4/Y9uvarxuIt6avsiphBxi
ovptsqeDHDryb7TzLM04lzVMgFzyK45rIOlZ8qyHnHgPZRuRRuQiK6WjoOVm
MT3tSPQRXUb0JkKQAP2x4XA/JRv+E/q5s+FzezjcERTafzoYJZCgQVD4PE62
9VaI7H7CcmElMZ16wJvrF7cGgoSuzcLRxQ9FPgEu5hydXhBUMFxQ3alcXqaj
RFSt2lbB8sD4zWyKb+UpUB+QF6twR97t79R+wAp5RdfVatWGLuuow8bdze/h
hTj7ucFfloACCIuurVplE4OFyOMgoqKYA8e0M3gyV+hGIo0uPxolN7DZg7IH
UJg45wB/quxvLh57FlcJ5cRGjJP/RpBukhX/ErxmEgUT05dA+GC0cFE63LoN
u8O9kh40BlPR2cVolIVlMCoxG4WYT3NvEYA9SMOwkeQGxhFDLWnOPBRbB46k
JsyJ0sGc2Cv2u4lE+rPWdIh0K9rNDA1Gdkc1W/hQ/UOQKAbDc7Izkr/dkRXD
qjIpbJdj3ue/IpTPYyAREaQ2WGbFmzBd89gy0i2m4FtRa63wC/E5kiU56F8j
HVELmkDTJpv9eKonxwo3VdfrXLlsxcD7OOF7wVrSb8uk2+kKVWC+9vnavcWT
NTiH038MsA/GsKPtCmCKbR+JQOedlmRyJ1lc9fn3w+Rs4cyp3osh0BOsoH65
rAQQqMh0RmJR23O2NqNZDoyZJYXz4Rr3sJJWjb4WKbiFfMFWM4c0pii5o8uV
fVWQjf+DhaJm2+E7y2eM+LnfX3R+oQiu8yxXDFs+hf+YTzFJuvsJEcrd86g8
+a0QuCm0TLVnumLZz2V50/D5T4PcbHFgxb183C+FyngAI+Fy/Jp/jTcN71xE
TI18k19cBN16GUGEynJeecQ94YrIqYGbn/8g7wxuD0ITXdUtvzWyyVPK9HHF
qSq/vXkTAbidrsBSmGIF2dnqX/yK9lUH5now2SqlZ8tI7RZ3MwtiyEF201OD
Z3dOrMNkwAOOdbDmEHRt5OIGx277P2P75t47sMhAhwbWm6mBo51appSLEurp
uvCUf5U/YhHk5daLZQYhvNB2KdpFK6PRJZXVr09dCRcFgduxeMD+E0Kd94u0
WEQNS2K3+28yzWXbBxXZB0GvhRz69HiOy9u9WOJZTb+bpb0TTxurVObnSR35
sLOSzBaBYRQMBQEkAbQhIe1kZ98qlc8PkCkbxAuikLsyKV3Ly8QS/+4hrKCd
jOLE7rOZ4N4CJpNalFX+uQWUF610G7nrUPyVxVAs8J0mT92EW0OX8YpgR/uA
LogY/RBTLKnrcqZ7j71f/2dTJPNt9EURVaowBPm7W+PUp8Qy5Qdb8ijpbP0f
v0Bw1PDJ3/Uql8NoGDbj9HoCn31Xbj5g4QPRxsoF9OMorcogSs2Pxl9NLXI6
FLialy6Gx8MWRN+Aun4NsMY9hMSGkcz/6yAsYW3Y2E2ngdW0neek8uN/7MYK
yVSI0/f/uVT9cZieQkCsFqzC9Jsc+DiKDd3E27AbYe2TpMCesxGOYMZMkUTm
UPY+lBFAgqyJeThhOltvyu8lT0WpYwmLRNRwme4nz7g2ROnyM8DxCDcjSj6m
9aFlgCWrMvyHQWkyEiifr6XD8O4R0fVnbO99YED4eH4UXCfZlqtvOMWLIaTz
4EiK6aoeTUsweZnvRqQJAP3hrHi5JRWfiAwATLSfPv2cby/+tReain8Dn+NU
FxlDuvWrs7xvMTAILJKL3FuM8R6vvvbF47cc3PgQvX+2e6fI6kQ9zP9emxbA
lq56WzsKdVk4jWHZeY59E9ArD9XI6Rak24HOj+Tbin2aQRI8Ng5mug1MgXGS
G6n7yODT92uLYftNEI3ydsVo/ol26oPoP0/psyVHXSmzks3zDpuEiPYerPHq
PpUuUZEx4Lz4GMaom9WICsBtIXlAvG2XRrhmMA2dfdrVfkBLXxnq7ihKIKHP
Dq0K+d7mqvDmS+og5kQQURz4DS7fh3qx686BDra2iuXJ7mffjWxrgnmIv57q
Q3ilrjnL00E9B5yx5HgYsfZXs2G0XuUdsSt11wK2k0oj76TPpAJ7D2wMX3dP
WQyRRU//sXq8NJs8f5hTmPlnfJcgrT0e6Xy3BITKmjxuZ392Tlx4m0WqjrbK
LYOwW6wdPbkO/EN8oMk75W4prIhBOggkfp0mp7TLtToUaJjLahvFsZQfEvrk
NUm5fNYgrB4DbdZsMh3LoIBVtx0ljuWQaZpAWSVGDqiF0xKZdYIwwjd2L6t2
xg6DizaS9+nobOmU4L+mhaTSfibQBqpPGk6xEVUpn7PCueKHvjBZgbxJwjgG
cKHo5ZMy4WgxIFW31VlKpFjUHVajI4NOV1VVgBu2KAKPBw2NID3mCx0vehLX
dabmgoqxkLPJRou8kghZkGPq7PQik+o7JNYblWkZEy6j/93IrlIhQHGZ9mH/
LpPl2rYF82koDLvurvxSUAhYYBIY36PldOwEsY4JdMunDn048q8Vp+JqEis9
HDXk5W5vhIje7Nf6KrHt9DxKgicmTV1JZxvsbu2xKo5SmoHeYirlyfhlCq9o
l/53DtptX0dqeNX+k7lNoUdWuNU4lqXGVSSN8n3G2FUoDTp+Ak+eW7s7U1au
sZjrXuD1z6kFh3r92fmkHGb7LQDlOEPOB3iXkrhug/kye77aq5+BR0RjCy25
rJeGLMhOqRdxgDumXkNMxRZ56kJaeMoKQ0Tc33nVby+62t8bXtsWPBOr+Gkj
5mqe29bH7abkhp2/CWGq+JcdGGzUKmv4DpXg8bLR9HlZyQov7CR3NNRBRzUP
LXMBmjRhxLAtRCz79Z9apouWOB2Yotcz60qFKJAuIVkYvbcYdgNWdbgalulC
CNkLbv8Ha9z9EgkPCw3N9BnnMwTtuymJZM0ndUjY+OExVdq4AR/hdHlanGrY
tKmGGWRPfi0a3U/BkbWHQhuT3oVv3u1WzenlJpVzsHmyvcPLyiuOHSjCe4t9
BBxWNM3ruAZKAv2EOO/oRknjiLCnObIXc59vFqpR0lVnm/mkoKbHN6oIiF+L
mobQv2L6JBF/JQ3eV3KPTgD70GtfTZi/3S12byz5gmuUI5IkWLotTUEUk40Z
bLI7eSSHmmVoRbC8zPfH/vZp1Ay1GuI3ZC27ENr2hf8lz0lpmXojaAYu57h9
ldKCbJXUUH4/LeeYZg/Isenmg/wsaozQah1d/0SftrhjgQh5C6xOUViTHN5z
UdyQ5XqJq2mg4RPGxi0sBWkozwQz8jc5drvd8tEoYarIvOOwyop/BqOsvcF6
Gbig6Mk8hJ6XhBhPqNTe5aBxWxH8lkU/ySmjHiAMn9GS4cufhYozQc87mxBn
ZyQrx+JWdM3CpAKaGCYqfr9yKUSz68TQAiWl40N+6clTRTmJY0bp4pY5NkRV
h6mZd4/vyKfM6BW6LcvHJc3mIZiDnEc5Qiq79NiHuFuzo2lCGyFyQTTgEITJ
7xTHnodNCvmKzoNH4nyLx6cStG/vAoZY4VjTS+i/O8v7lrfDNKeyEy/gc+hX
ExNyBma7ABuIoGev0j4CK1huhPa2hItNHt2GRghlHVQ1nA77W9tTXkyj7EYC
tmYSLHLHOWKancve0vkdF6A2Ui/GV9ArIfUKpSj3GsVqa9hJVFV1rkhG25Ld
1pfb9adT7Wbk6kEQnyVXFgrawoJfWZArm+5Ywtvyo767XeGlDYcQYhtyw5gO
jiY5pqZcVjK4kLoxz/KbEID6M9ocYTIm62m7U1LQkCsrYguKkq48GkbmP4sX
c06tcXTVvJvpcKJbTHkh8//NGPvliZzLl83VLbcbKY305qJkwDfUjYqmm6bS
deukFDbIgoPu7XLV2L3AQW/dev3qFa1KQcX2c1zOPND/bMtGJCMeEKsfv5B9
wR/tXTyIiR4psDzZSCtpC0g+iR7BlfdNt6r5/MWyaa/9g1B8Xp58NeOpGO1y
aJPhtCYIgm24FNBkMIAY/Bq7llgR23XsCa6z/EzxGvDScr9+O/FmTlU1T9Op
2asqwU1tJDQ8NkADBESvP1tBjrne4PTJ5SU/oLh+tU54UxXnpC1U1GYRsQXU
Y0ryx7DH2PuW5qvyFDXqC9plw4Ry/NyUV5iLSmdeeFb1lXaXoEp+ZZTOhRi6
lGUAamIDYV/6qwc+vkLRpPzJoWH+rC/T0A5X21hEGWkxQ18+if2KOaKniDzI
hOE1F7dnCJBLuvfUKFKzzUeekooDeUHb6e26PhrTTjGE4QUzLvFNnGSxaT3i
U0Gb0zkmWJ/XWOloSBxAky/G37cGc0MxH3hp/gBtrAii8N3O8El2teObRVEW
zNikyjV5TvQKjYvc3Esid5LD1IZ2OwLB4fGpHJLPFTsaflA5ibjxgG8cECKy
sFaMQipj7KluOidGvkkqnw5sjrUkLIxuh0rwsH1zzB0cLHP/zTyPaJF7UT76
ejtnp7Ah297Ci66gAgkScbM+f3d3OYefL+tUFQ7xYbe/bMCyBKHveUfFo9NX
ro4dsf+qZH+Ux6mDYoRBcyKDVwNFvJsBV/TQZ2yBtPC0J1jzsc5aglPaNaA3
qslLbs4BgDHVAt4OPejiJX71aA+wqde6OHMWTDX+FeAyq31GWMjxRTiGfgOQ
gYxkdrQAfIuXdZDTFwOsU6alWdBu6SZ1qLEFIvC5zTvsPoT4itlk3IikmI3Z
SHfq+Ylq8tJCpYP2gqCguOaNk+9lEnYhUDrjDeZMAuwo1/6S4+ujepK+W4uJ
oiqXhkplcqcGdIw+otfbEgiiegGsPjShGNgbFcClFjLklu49Mf7xKoRwktCB
RdLC5qOZjrm3+zkDS4p5Vtw9GB0Bh9JOHRHHSN1stIBO11Un8mI0ehbtgf9i
ZswxOo+uMOkCD3ovXCGIDcASW4d+iW0A+7UIsVB5epnCX1NWnn4Sr9bHXVZm
aD1lahBmCAzsc8aBp1Tgr865vZuRoSa9feW/pCKoURUNHFoWp3/8Ou7LqkwF
Ta4X+yGkTSJGVYOt4iMvxfRv/i7bS9H4VcnUOkYpBY8GYFBJH2Fj9ZtjsKJu
p3+Ip08dO5FxnzLTrEPBNX4wDZfpOtjAqoafyIQdf7BhHiGXBveqr1yLhZtL
1sBY3azN6bCZ0x4OGTItSsithrfVgGK/+Pb+bD5PhTbRh4gs+Hy6qB9boMab
jUfDmp4DnEcTasJfuvzLweHE7wKqBe7CFzpxityjtxKgtXdLXINCTUfp5QEE
WrWh90/v8p9FMvbPzE21M4CH2oEx9LTk7ta6It8U2RR0/KXe6/f0jXer3dby
TuIwMTBivOFQKkAN0mtg0mjXfx7J0Eh6jPK8YgYy24MfTCiaPseSy28ipJM7
XvyexROrUwh1NHXZ5reMD77l6n+I8ipgos+UTSr9OkxZhZuHCR/8znotKgE9
61gQl8kXXjdwKH2+kDOzumzM9iS52NDlEPy4qhG99b+I7+t2GRgNoWNUOZbU
M91vFRzPtm8K7MvyptFnjWRM77cmzwX2gnMTbTaVa9O1EHaazq1yQo6Ncnp1
FXj3Qr+ol1wMasQpn9WQoRXoHtbNm/OlJBOHsvduB0g36EOz2NqN+2JiOt1p
pvRs+QAgIFETjIbgeLdL7MbzTTZBBIbToqKSD5FF2vdYU8RkLViDWXif0TnK
muywZWVsIDNZQsUt4OOyYdPzQupAJbvuFXiQYAycwPFnHsZbk0pt4/rz4xJ0
jgFk0Ci6fIfZuSSBJSj1Be7tjFyrlQ/mssqlu+pLl+CAQlv+3AKvktvCZC8d
xDB6Q9/TgYHWYwWiRal/y2tjaHUyQ7Qz+sGxv6xFSg2/ZDVuLYc+Mpy1j06S
BecLvNiY7IEExciljBaFtEm7heeOQs5AEJKS0cwKtXuR+8igjR9D1DTb16oB
s/Mf0XqmDrZ69T944WhwOtMDe5Zjcq1LjP04TDtSXXjBwjh18PHyoRS1y8nW
Pylgdfs1soM94rx4EMVMahvdEcW11QW+CHNxQC1eCoXJmZOT0AGsE/ji+tCR
KNjBwvolNKFzLG7Aut6x6hunHSkRsjzu83qQDCnN2KzespDtmmUn7vs0FUq+
CyBOMKbyjQezcZaCTqLMrWjsI1MhMNAUSF/FEzhkjc958Knsz4gGn0q4kr0a
+wiStL0WMCDippoDsqEB0EkpjVZZfdjq2ZdJnToSnQ9HhP5dHlh0Tuh22iUJ
amfSUKMd82qVHtRstmA0I3jQduT4O99rdXJXsd2SYItrMdNjqL1g++squBBw
GXGpLvxcELD3XL46chYOJ6CBOtt7/MlSLkEwh56RHVtcoLG1HMBznM/6ysdz
K4CgIgbuLcCTi0dVYC2hqH+HDONzQ0c8LDm/g2Wq/P6Xp4iEpByNauRN/KIf
xlodiS8JVdMRpbk2WlzKlIfz8/8V2kJH2IMt5pq26ZUpKzbcxI0CMGer9WZ/
Y1+U0jJXZxJ4GT35tYnwyaIccS9wz9+F72LTaPseidgfgZFZwV+0tbp0ddRI
MAW5Ii2sMie8ZXiuhyyeqpAd08MHCdkbe1TrvgyIlWG0TNt/WmXCuUXtz/AH
lF+KmBOWgM43xBOiD5M4yWxfdEG5vtdUOX4RBbDnJlb81R6Lfw1V/0Y2o4w3
jqOJ+QaBrEqFnGAjg3nVLbMLhr82LKaiSkVwq2MfUNgo3trSpbk/FyHVCgdo
8EFL5chzqt11Rki8SdVmgrYiIKsRMLUWuSm23eff3Od9j1SkUMiGZV88xZ7S
lKTmi5qCK7d3CpcvbofRyHPWZ+vEPp1+2riwlHFi4xK9opim1FMISrshAcdy
nVe6cBqYOkhIPv1CM+BawwivHiDyaT5pnY+ZRKD5j43p+DlXIxNRvs1YBa/G
B3UfVy/08yNWrKRKqLudnloYfJL9q4h7GFwYDbeMW0v1xBSAYFTB1z2xADUs
jGXkJOWdzrx1ks60dJNxaucFmkNadq7Ub2ZA4w8S9jH2x1AMYmExdRGAMnje
SWI0QL0nipW+VijrFC7+XlVd1SCb5nibyYv7BXGyI/WWYymu9gyaYLerRFkt
1+dxwSH0ay0kQ3fQYzzw+h30AYeICxmhNVnIcjcmTtqz9g8m374v4MEo5hOx
2Ieg9aKYwL9M/9cELNjxiU0/yY7L5r5Ug7+6tfkKVAbRWo1TyRYZEShrVCCg
ApwyxZgVlbdvBnAqqVKBu7bzv8nZJUKlVuR/gWvq5fu583oh7wjnXrEXsk0L
0cf/qL966LqX/dzDnT7zqKtVKx2hU18Ndz1bO3SilxqYdlXAH7ge3wRZw8dT
JEgLyZJ6c7SQtTY+8YzEzZKhuKhEI0y8jSAIm6K/gSZJ35oJ0P0EVR5dIzgZ
GLYPXJ9cxvQ/bEEc/AHcpLkOzXIT2fc2+AamuiWcY74ynt6fIgv7tLiWKuDo
d4lm+3ce6fJLCowM7Ga9JcyTi6dHV/Fz8NG+hIZEd8dgzxDDRIv1DjtrFmzf
CXSfJc0HjSJ8fMOns0B1LrGeYRSUivpnUa/768uxr8hNyDnd+5Bo6jiqyvW6
0GNSnKskvJAT0sOATPr3Kf1qx02a3LgE2YCrzrNrzrXwtPW4UwRIbfFMptzp
OvvYg+9zhqh8Ii+wnVjefvFKdKHfr6g8WHGknT/C1iH81Vbk+/F1EWFRtdnw
4Wvo2QABabOjvWSMK1w1U0LuD/u04J8xejHRMWvaJctBJonJjW0X1L70PEM7
IYQTPYe+fDxBOoDwH/gOhjkghKH1A7VbQclyNjlDCt+NZf415z7U5urQW8f0
l+Ciwzck+bTnRJK0An2GCk5L+r2cPV/v0z2F27Zz00orAPnyu9rPqseAko2h
CwPRn5s6B2I+BE4qthVOuNta+DMeLMs988JzwijCJuWDToxktGZyYWPXeMib
QDuVzDJsQ7IK1prOCJvOo6Pf31roLXNG8uSG6KVUXOHYkUEJBlhoK8YIQtuK
Rnx6K4uJ0dwdWroqxpJordP8Q8KzNB8iGHDzdGUHsbS+VLDtc53xU5z4XZOj
aA1b8kER8OlSA+Dbt9kjHmUGmc8W9J6FJG/QNhw0Pvxb4y1ELTIm+K9sCL+O
xDxuYhaj4/vWPDz36gYKO4rar8Hy9djxj3roijO2f0YdXtY8B9+zuEmGvWve
puZ/evqVh9SFss8g/H6j/VXdYMZTXD7ptp0aNLMG44Nxeo6RyDUCuV7HISTP
8bIVjROt5doKTYihdmwYE0MrvUyMsMGmj999gs1pyFd8HnmhB/pIPU3QOfYI
oqKoNvU0LZVNFVcW2uuC4D/VonqQvGribFrex+SwUzk6tz3OrE+PAIvoAxZa
7KKipl/fDpUO+GT7mnOkryTkwPQA3qN9pxHvBXmzPnv/Ds4lFmNAj7ThffTj
0CrFC0B74PAbOCACBZhyMdv13dca2DDiAglZoBObRyLsvEBAmxSh5MaTaQvl
d0LPJi42azmMlL1QC0hhIGjc/TZVp/5Re747cGXgD8z3oizK2uEYVHH/EuyL
bmb4iYvkC1tJqyhje/WjcB22Nc+ZF/1ETtDkw0XC16ipqkjAwZtkaVQsJ6r2
UbRMA4NEfKoaLORt83IbEK4ANulYUVnoW8SnFB+xg8bClF/8G5mMIIWlLKrL
TvXeSWdIb5IMArBQ52kJpvv8/Pp8TMLavqQmRANij21Y5xaBO19aNqhDoLi6
ERhaBuvggjgL+RUyMncDfXN6J/JlgnvSnhjygpdFnJa4NF8NpwacXM0FIGiA
HzpRsWA6cEB4l3G4/FpkkctKVeg922cuxryCTYFlVNStHMJFMFfPR+3wnny0
Fkj5NJjS1EMHN2SYTsoUBLUw5k05XxTknKDdsAifVrCfpkET3iw/7mFm2is4
MZpyFnmR8jHA6U5MH76ee4bH4VkS2S5ZvI3Lc0ISKy9atL6fH9mVWvqJVQlz
zqQqsWPt0HYmLvEBlAgrjpuTf2SH+YQAahdHNBajJD6dseChFOgGADrqAO37
XA0boXtk03sZE8moAbytdGA6uMgARcS4t1yHbngMcv5L6+YPs/n7NJjiMEPA
6OKK2runmACHXbuazae+nXizwzJw9aM0QSmjUsb71gI7TfTxkTrN7nYFIHRf
gNY5wP04dmBZOF/Mwved3P5+AaEGi4YQA85I5clUbSA8eCnAO2ywW5X4RvqS
r1+F+euXhK078x3R7gHi4DTdgYncPifWIDpV/I9DOWpWY+UYZZGzNAqn2CUj
NQOEyFYdSwPFVbSokpRGZoyFzox+QHABBAWPKTbuR21fEAn16E07zGocviuk
TNNW01aKtDS2VGuxS2MTlq2fDJ+1C/zoelPjkkEQfJI4bHu37VIOygMy3myK
93moHaDl15R4mLmXKNXIxxhyFpnlp03fXGOhrzpxIo4Fh11aQsWajQCowAa+
d2nAazmct86vhPNisrjDVi0DEjJ2s/WHenw9QF5NkcmjXWWfRCWTRpQ4RQAv
b4GWQt0t3sZhPh76OCnhvzM/QEnhu9uHTq9mRH7bIxQOy548NYyAaI1zgWM4
ROUr4cHFr62tMYbkCsWK6PSSdhADZCP9zqNJrMGY0sv+W/zReFtufGhcQurk
EFzzW05mMtp6aznwksB/QliGMSAuWRbe0SAkQ5Wh4ASJkGDFDK7z8aMKst8s
Wx0mQ946kU9AWUAbfAVPZOL4p8tVUnOWdRB+p0voIlmPuy04gJS8AojnlCAW
5L0eXLyBQh20AW2Q71hEjwh1DEYnwkvNwajX1CdO1gnHOPjF/nsGoBPDBIcp
JouoGwBv5r5HPOM7wl99mzwrmOOr9niW1ScUL4kzWwEmjWK4MsR4Tmi2qAo9
9SmHFlhor8UM99YgD5ymGnURW9oCzPw9F251H1b2zC4lDULaU1MjUFHRb4ZS
52jqNKoORG9rduan17dwmb5N9nG1zH3ZPECrblRYwQx0Cav96HAPwujQ+FCb
zDBZR4NuVn+9MlUmO/vTdz9qta95cr0O4MjXwKWi+9PnjbxhpbEuZoagDb0a
h/THpcCZP1UgrdbKu3lkht/iUb5albo4ETP1aklIEX0kOrfzCSPoZn0n9cbh
88D366hSj+ZTr8DNHm4a0hRKqgRvrV13wxNznJ7w6ctGanuRWuzbYW6x5slm
PhQtl5j0WWLIJJPrJsfahOwKvu08f187f8qh7wEHQrVbzEWghQ1G06ir+wga
lI4dHLKWOabFvqj11MviVFMfCuocw75xnaxW55k12gnd1axiD1S24zKN7bXJ
dxEIz46YKnfxy19R4nNHhncJPMNQWKgSbniY7E0id2juW6h0cgtmbh3m2aQz
c2F5mo6ytNymyJmVzB+jPMEqTcqphgbTcVY1r1pVNDa3vx+2sGwbqUymF3AC
2Z4ii2yoOeGwmzqxV5DnfjyRmpUJxGTwDPWJMkFXnz8KeF6wYXG59W3a84B+
DtzjET7vwyeSf6m6Z8Cd+3/M0JeDZ420EomQtEU+icUGJwoLT5ZJrAqQnkFS
ZteTm1cnXyzXxLb3Gp37cYQa29+lJT/skHUUtlzxhE9DtH738PNc0W/vZ2lE
l/u9Ee9hTqOVSQbOjiW0zPbt4Vyl3dfJBsv/ksGBuo/Ru8KrYxl2EA+zzHGU
2iSAud9/EXEGstL+sVQFpWes1nDffPd2un+BOA8977Xv23rEFN/iElc6je8h
21XxOF451xb5FZsxEb5k0iiWs2eT6uznFuwebcy9Plqerh24E+JinzmkZPvT
1eAr1ZIaDp5jowYmNG6xNGH+bV1LP3OglnfRzn0uTUE5/rujaE8gIoi0qEUv
IX32FX4GX13RTLdcQuSQwIVOgVC+VW0sC/oz1qvo6KNliQJX/T9+mQpSQVmC
ByUTD+8512XHa7LqB16R0tIDDbvku2/mr9cQ7LIfvncVxm6BPiThfNMKk32u
RIDbtglp7LUIAgmbQLrU4m7Ije5alG6jSLotM7NsF6W+vpEaxs8I/SNnds/c
Brn+2FcR4cH8/S7EpZC5UIhTC8lOhLu6ZU9pj9h7zo4YmZi4uSXbESlW5iAJ
rGPHPu46ChmU2vyZGZKsi3uMzLjaE4k1ncPJ03riyn8ZPLsmIaKMLeM5+4c8
9zsYcgNqg0oCyz428qSX78fngf9w10EhVGbT587xCoWPu0lSHSySrHDGxYKZ
Cs7zBTXGZsnYBHeGut1IhA5BG33/c4NcGvhr76QTQSkMbakigP7WZCg6fLQ2
BdiTi4ScAcbbibqEkzRrmCrmV1oSCkZLFBTSVasysI2MNFO+mrynPbmwfZcP
vrh6wHl/Z5KxXHxGRqwL5Vi/8La5T8ut6mxi3qQ/1hP/FaVAm3vZmc6o311q
1OheB4EnllDkV4EYAa4SYhLFR+J1DDF/ytRirLB6Pp/8SSgfnOr4U8KRpmIT
AyVGndl/Ksx88i32GcZDFiSwJttlwMp8SA42cogf1MA7apjCB3/k0F56ORNu
UdJL6W5KOZjYaVL8eXn45Ek99EQ3mRYtmCxj88jNzDv70m3dtHhnimsxWtUm
OKd79SuRuQP+/zrd3xH47R4xjT9MRQHubrYsZUo/gTcSlJlin3SkYT5LQB2q
+/QleoumeVvg4BVL+ARRcXXKMBV9XBBwkT9FYB6IJoTZ+NzFehevTQctoie0
wrm4NJLC7cL5IgoihdGS8LwDEJX3Cz7Pp+E3fVKhg4nONx5P5DZFCkBsbnbz
/KmaeMdr5yDRJj6SwfvUyPao9V8HCZeJLKcc4ejk9O6Vk0UIrWhQxO8OZd2Z
R+JiHmu4xrFfXtIxkCdC/fp4uN77uVx4rNXnfU/785n2ONwWD0qlPh0pkOiy
9AROzOIDoDHKgry3JogNnVytZMt+9uK9qynuQKR016VPRgwv4dH0Kk8jlv9v
2f8NRRrovUACf4R0JclpjNrFKCBk58D5oIqZwXghA+gAQchzMnB3UAlbOXDa
ALDtbo2AI39a1oVExOVt5eEsb7sX3di57sMZni196o4eWOxpzRknUNYpEC4T
/3TedaoqlPMe/FPvSkY8Z3s+vFI4WnyNLYqFSZJhvoaaFa6VEDS90zJ/T6wy
00/3g0yRMclt/NaHMbrvbxzBwpSlovS8zpsqO6bfml96pwdzq/Mfirwjyztd
zW4V9gRYnVR7l2Nm05yzN+5TxxZ5JhXR4QknyTo4vMP3u6Niz9nhekwQx7/h
k4Vd8288HlPutsHPssBb3duJLWG/ESqkcBiF7MZA4GauTckcHbNVYbxiaX09
syW0xDWPLoussueD/Ol5w+Q5t5XibuLDNdh36SVsyhuGWS/PK6j6YAZKmPcK
pEVJOvO7FC3k08Gb8rK+M2v9e6n7jvUXbW436p9/1XKZpYneYeyZ91AHMycz
uYxYIo/Yr1Il+J0Z7ytf0bcJ3YRd/X0N4YHB3J8VPTPgSf83J2y7jsIbls2b
QhOAizwyf4jrVlFCBKUc8CJW++Qm6GwkO9B4fnQCcXHbz9kdvo3j42DHVatn
ORBtIH4BUKzSYt5kL9etnMESvjHw1gWgk5UkY7/YImIo2gy774HuGAZYWsy9
9BAjOMxPPyIqK0SNe302HzZOCE1A9J2dgjoPIa9f+PNC690h6+elOvEOq1Ne
zOlVNhjQkh/sADUn/KU23qH2cn+Glmk56cmZ9UMK9qXs8BPOihkUCngk397X
BUItbzLEY9erFs549i8+HWfKxFsKqJMXb9VoaGl+BoRp5e/lwQFWFgHsbjuE
nnuVYZaC8bO6t31O/YD2HoloTAAO9GfafjOokWhBkirwSMHYAp9CuoW2fOR8
g+VAfRptVvK9BVhde54AHDBdpy8/calI5BAr74v34x54E2i4atQl0Fzc/45S
JSKne3zZxJ5vynM3GXks9bKvkCrGvcjhMWD6Ejh+pkx6PrhVoU11HTPylOcp
Jhe8JGAfPQc4OxXLRCA6i3ieGVdLRDtF5Rr1XRus1Q9jJBhGkYcevwsYS1wu
0MrlOBTzGgpSP7Rc1KnGkYy3rrjBnPWOol5fkTaLhaHTE8m6+C5bY7ZY/koK
MbRj6YCvshaeWENuJnsDbMr8xR6Fdm9O99rJT4+tBLllEFdCixL0dTHZdvWI
PfCz82QLzkJGz3V/lzk3A+3agC1TdF5nP7BMFGerOP8LvP9Y0S/hkiS679pI
iSey/lK7ZwP8wg5eVW5P0ptGtODKvK/P04SkQ+0fgAjIzTiaDazjs9SpOu97
ql4kJ7xn5PheMH2iduhbeTUj9vo6PZAvTbQlUQhg1Fqiypmr7NectltK5oE4
sBE1m1x/UVnEldvKb63NRqGcuW85+Xz0PPXpQugdRruKwqo32Ty1YJa2y07B
YM540O6VRiCVqY2QaBZPZZHwr5GOCkh86lh/SlGY5srMwVkCKGHZcWx9Nj85
8gdenGsYLaBNyVpn7jRr7swr7ah79JFSBtZIMWXgUg/j11mUgLp5eMzjRkFi
UxRFkqOsQTO2I57Hd1dgm3kOjH2lOT6jZlJMJ8jX1MDi6Vz+03fB85uzH8me
oo9rBJchUVETqv/bswhkh6yyxvk40MKPEcrOuRSYw8WByRKnDGKL9vdxPmkr
HVoJ5BxJvaeCwaawdiokNVTu+6iG2iaV3ELYhWycb4LRYASCcvbjRsHvssDg
QvNT7YuAbwiyUfEvz1WgsCXnbUuUtTvWvpN5U0IQOtnB7kxv+Hly75ug6iL5
ZdBv/7V7nLLNks6VruPIYbdkfKWkGXhKN1mKuBycLrW6EcnNsxRk8B0ZjKhy
Cn4k8jOs6DytIa32/MKXGwNVDlY6hZhrc1zwLuSEHh8m+0LgoHl5qqu2BRIH
uXwZEtbl6EyRpKGg/5Djl10gyzlk/rZblQvIrdDEP+amISjydhhkarBY068b
qL5SvODj0Vfo06h4oXcNmZqDFacZkFksf3+z4gYGhY4w0RRrkak2URO2FTbx
fmB6/U5YGomRCoN0GpmawCuwuhbL5aUgX6nzicBDTek5+Ie+zuutm1Yai2zf
sUXybiKg/844v2JXNqp43Ki4SDa5WgHQRMFP4iHKrpMq9TK5kGS30Xwf+MhJ
8Pd7b9t8MN1BIlHqzS56+ph2JNZx442RC4zfgRk5AaMt365NhIygITtoIsXs
4qktqDhzDn90AWPFD06n6dp/b9ttTPgEF9UHirn0JokiHo9BGkORBux6P7Gt
2xMxooTpIO8j+Uu4G7yVDAYKCIWMTbiMAvzlG9aV1Quiv0JfscXUXZz71uoE
6r4n77zYyOsDY0se4b5sEqLrDpX9o5eWOvTbk5qqc2fBXEcNKtEpJ5Accfb5
j6ZcqoRkC+/1uac4u9kIkI31dvznGQYr5hiqE1NODhsrC9JAOAFNtXuwKy+F
e+xlefNzpbGYXPx+HGjt7Xhazq68N3O2Nl+F7UxHPO2PETFU2S4omn8dWeap
/syd0C0yvf7cot1MerjqGrENwreNzYQNRVc8kDb9cv4CGQlxfEMy4wU2qnEe
ug6CHHYkRQGKLOmjMUcexshQvA7/mrM3djcH66ja4rMJg0ChyTxqpXv/j956
CcndWGCsnPzq6jh6XeXyoT5TupLrZtfpezKFAX+sXwtcczuARQeTBZ/wJgaI
3Tcc3qLcicmMovFa4Ptk3gubELpkPKz0dEaPUnz/NnF1Db+Tyggq2fZxxDcU
biJCqOqtkXwgxygnC2Q/LF2ajyRlLAaxEUV945aXCE0H1qUfmS/dwOW2IYbQ
vutIPVsUZh4Dsov6K9dGK2dhAz2wNMEWpEcwUt96lCvqg/fReafcvZTOTUtr
ihRihN+OfVomtz7LtFSxNxxHdTL0hjdkNojJr7lI4d7RW6HUZHpBj6pZLY1b
xHF24RIWUUX2DA26bKhyrRLvKkH6dG7ZTBYY6lGRPET/u3G+XlFtIOIk/U0B
Vd0XcTbDUnlgdc8UCoJg99DN7j6QOP/NrlQsaEKH34raLJqXDtUItt5aJSmt
zLox9L+yLcXTyAN42PF9Tb4G7D/9fSWhJ0oogiIj47+Ow11JMdvfUaBXiKzF
4SNDAzzuO3Bv3MxTkeJliEV2kPnwLDgwI1AW/S64mN8O1m2FgqX/wGEcM+Ux
ujjeGlWpnKpd/lWpg8GjQ5O9Tf8KU09B84V583j1uH4RjCdlCvhS/giaEqRJ
ftSqfQo5JHXpbXw94/zQxTg4RnnBF1fhG3ovu+MPj4zbhMSvytbt29nlafGL
0byC4NAxDkf5gFzdKxjybDB/EpwvfNpNVd/oZGrFBRhxKbPngPZrtM2vCR9C
VTQLhOH4hHQM20EefEJgvL9abfR7+ox+XZHlzlH1mHHhgqsKx4sXHZxjuwN7
rcgXBYulAFatCohVHDSQNYmS4VVJi0l9HxHz/X4DQV25kadCFDwZKFM69zCa
XssVhKZ6ZgSPfG60saP0GCUGYv4gfd50HYPFVKlcHBzOrncM3uxzUeQP2gQu
9pvLMR2FTor5TBPhjydJmyh5TKq3PcGodfSmDZqEQ/FzwAu89zSsczo72qXR
4Ie2jPP5zZT9YmyvudyOhftfDgrMJGyCKCFLiYLPQ/Hh2q9qXsDgDMxJ3lj8
NsktE0O28msU4clTAKXzfePDjCvYkoSNB6gsWPtqJXVmTU8CNDHAdjYLAfaZ
1uEb9g+uQljPOKCTzLChicWG9s/mlLeoSC/frF/e+lNx/e8Lheh9dMKDNF1w
fIannmUvyCTEWxw1TDPXi8zVXGf32iPhgoAkqWkkrRIlmlov1BERIuMYOYwv
AuMZQ8M0sD3AkWO7RNTl2GeJbSqBRzezUWUqyukizxjb0o6FDJ3X7PLCW8vF
Hk6X/EsZczUvui2DnOvHNm6c34bPpXqIj6npOrYm7TQilmAIkher393Fl/NW
fndgqIYHrvEx+IbYAltFj4xS9+muMwhrHu5Xxz9wpLRdaYBN40M21qJ+V1Yn
pg60BjFM+HuI4NX7xqduCZfzPrYlGXeQZOf6F2zZ+bXoevz6TfHP44InxJ6J
0NAuTZnD1cuUtTgp3hN3QRbmtpBm59khV+CtSLGmHjRpf7x9DwQj3aSUi1bg
QK+NRHTLFmlLzqSDAJarvs5MiGReW8qe1ucax2EcA2uNl3rdcs1fjRa9F6gA
tRGNx/piyi2kk9XMvjVpvrdmu9AlBG0CRm2UAgmWgV62n2wcz/P0SaTkO0jK
wbRiF1CbvQ/xbahO5Wm6VYQ82m0CepSh6jniX2omtW7ftVNVHUI/RpUt9LFV
bTi6gtE/hEXHK+dr+3PddJkBhqUx7g93izZsVBwZL3hDxXlmGqzQiUPlzrZ0
/vx0spoggoSbwhi3WY446k+mgYpDFhRZaidpIv5KaW5LVkBsffb8lVCoEn1G
UBGhxSlY6wvvUUCa6So6P59RNjGj4tsodozCKmaDuPLGmOHUiMUFAjUWhWBf
hLKoLcHAATVpq1O4ds8rwhjn2MxhMqT9Gy4gPTTQb/inEzPAOP9QjFPb0nRe
rXLbdp1reU08hHqvgsmE/XFUzPd7A3O9JWAnba4nK82vBL6IebbRlWXzmyl3
m8n5bm/6tORDE34+f5tZ8Jjbn0W/CF6O/TCk6lWt5v4hRFE3iZBQIfpq5tEf
f+gDs+XoEVkP9cv5ZXQtcD9m5xn0zdzA00IZT4hIhhOGxfFqY3Gva1Y9aksW
zjwh+KAWVGHjl3hH3NMKwkG1DMqshjAE2dHohLTyPdAJQCL1JHCqDjV8Rj/L
Qey8hxKX66e2zqT0Cqaozl17cuLcLcK9Clz9jng1LRfvr60GdG9ptNG4h9OY
oxXxkMla5ZGs74p97wIr+3iHpp0dOM7QJMMhzqvzXairOfP9OLos5PUZ7C9D
s453I3TPE4BZ3QOOS1pRS5ZSK3CkRavk4dTEEdveohwow2lIK+2yn86FVcJa
oq/Juslwnn0gjL14+X5YbHiBNtHnxD2WWrjeSblQh8keUA1TnzwjPPYT6h0l
63ZAWK0/LwkdMpYhFfIaIowLzul+BvcijRXu9gxooSBGncWO2VSbjdfpeYot
a7gMq+yvWGAnuyfyNiguKG1yAUx6fyTgDS40CGuJ1KG2T8oFSShphgKYJ6jZ
mnXyKbPb55o5GW06txaYv5FxWq1sO2eryduVvPWCfZTDD2O6VvH7xe0piMRm
U5ewEtgr0qo+WaMMqfgbunHagPb8xPXhy/L76jl9vw4FRukAh3O3UCBfe4PM
YRr4n0w7Zaie59zDMUsFAWTcrgHBSQIaNDX9gOAFwxpCtmbkAgZmvsX4Fx9y
2tH83PT+DgzGFGzxOTA1cbjzu4sdM5ScEI+j9ueFFYzTaEXfi5q/VnGintUn
VWxKVDNs5uJkvP5Gg92WamQouP3IcaI6FwmDreV6iZa76p4QsA1TMJP0dtHV
fkhwwTSBNRx1cUWjsJw0nHdMi4LgREeb1gt9twRoMq8xe69bwUUXxkDSpDY2
sOgzPn9MHNemkf5rGYhxijQB+DRnbTFFeOq1nzy4cny/lcsW5qN1VBGC7XIO
iwQW0roblvBq1qNWVXtdjKhompK0X8tP+0WU7GK/kDQyKu9zbpkYmKu5uI1z
Si87UJ9jJ9q2jVE8UnCJryBS9L7e+t3wzdCfX9fRTPoYlD7th3RDZQXOi0Fi
4sthVhJ+xxWj6fO1RChUcVbA+Nm2YwkhWUaM8+Avfs97y0GLGVEOypN8n0fq
jW/rDl33PJhKHuMHlPDud6AVUc+PILNRxQfPmz9SIZIvcuGiBsPcGjmLOm72
nxhxRNgMLwtjUyHu8XK8rx6E7a8QoVgKj6boWIy5muNpBEzFEfZSvqmMBS1C
l/k93RLFfX3zCcL6FBcbdhinUcuk98cSLWzuCXyc0gYQ94LVp5CzbLFFFpJB
UVPnTQFVwRpaJCUi8uS99ha1vYIPVl5lAIMtOb5MHYx50dqRsIXA+4FZcMQH
ysggYr57V/F9nXG9eaNaht1XnX8cwUngg7dslCCMhjK861Jl1Qo8hJagEicF
8mZF3We8/UmqxJewqONqLCgFUlqTwmcXD8zKW6pAj6D+r42E7G9/lKJx8aZ3
VZTebrmriMVXXlQYNzavhG6raSuhlTpFzqo/b3+118VM38rj+n1cdJ39Rbqo
4MZkQuLMIlL90hRKtZxMwiOZBHB1/K2x975Q8wqSaKXzXNCggyv/CU3TVKWt
VphdxsunP774c4E2PDLgHo/KFhs1dmIEdtlNQGfOpYfllzD7ZeWMUSjpzA6s
ynU5M7VziIbJABwo/LEs/04phYw9gq+ZvpVg93t1t3CfCNHo02MaDc7w/jDR
uT6rYGCxCbM/5K0mORT4DieAbfP3eATlN+xiixCtEfFb7nZFMC9IOlXPppQo
R33aoHpwgjFGQXphGc6pei2nRaJAcL90AW2Ay0BnGBzeDlvj2OjwUyi2S62e
0H3rbAjCTpIlsm7lhigpKdYCDmcPvUKt7nTcaBCt5FoCIBcTBGITq9C8mial
KIwp4nG0fqkTxsSfsoMVdZxInZRVocK7y/mEb/PsI3UZKjOu0Klawun5+rj/
U5GClZxbzl2+ReTE20oWSk1WzzFhb1409NBNVjluvfbAUf9FvCT4tszb1CEw
enzJbQiBG1rxENoxEXEkPW3vm/NVYhc01wIwRpgwR+m5FfQFeDDkBWEbWzNO
zO6seD29B+ZD/4GSoHCOARAY+15FFuweJTxvfCJ6YLn4fqW79UTdq9nNf3lg
sBUwnGrN52wYI59Y7VlEGm28vcHq0tENYSTBUNJMIjB1qq7yqSQbH89iE0uG
s+hVvjXcRZvcvhdnWQRaQp5F46UbZPpCurFqWRdmWyRhQJWpFGMys6uDtuwy
cr0sEY+9dNT8HcjuVgUgphqeECYtu46s5S4Jff+lKwK+BwawlnPPGn069Dk+
UyOvyNsoF2Rq6+3TycvYta2rEk8xEtdEyQsbQQzk5MWVs8RXxNoWYmpTzhK3
7AAGlapfPtIp80V2vrvf/xYrOxwxBfNWqtPZ1UZIYhmLSb4xIIhEo+8NizHj
7JYnZZWh93pp6lw2l652n5AixDm8aBEZBkgaidj07D0v0wH8f7/SMAveq5gV
6FnHGTXIHx6XzQbaf9sQA/l1xR3l20pVpK7nJIgmtgra63+KzH+EIuTi2bpi
kAvNs4FGldhIEYagl8wSw8eWLkJ0TAkqtGUrBSmO/QnO29y2N/TTQ6S/DCWA
WHTZSc7bHkmweLsnST4vAy8SP7FhCJlIcyB2vU6bYyqVfFECawy2MFzgFsYZ
Hqjm/04Gxu+aajtfjX+fgYw1JDRGop8HwElmO5+grUFP17mFhhpMZx60zM8Y
eHcuSyZWrfGSajIrffknHmEGRTVIn5JXtKB8yM6psLH79K1X5Tz+7Yp6OHPh
vOR4MkY5vck+YIur0vqZTmq58YAELvjdAtGQ7wGnmTCGW0q8A2OAmPBkWakW
JwzK82lepWz1akb/SUqEaowBkxXUfaSzPw5AWSlwA2YiADHXVOKvu9wuxAm6
SiTymssPIVyIcE9vTMr5jZ52Vqrb5AE8mpT5f+4YbGYmF7ZPzOo+oR38vLcq
jWfzBj9y990KHK85DI1BINT1khSqUZSdmlIudUQHb4uW7ci1qpiG/XxJjzqG
l7KbdAWNoew1elCKrpY9uL6G5pJpRkpGyW4NkTKwXQcIcNq2Bh8Pv2qbvaFv
ljWc9nKDbm8h8j9fPkTrdPqeS8vdDwfHkET81icWBKpj7Zw4NDDJLDObqsZ4
5gdYiRDXXkq2sVYrQvBfHYAOIDgtulWG78vwDM7eQHokXbR6NE+uCsFEbTEX
GxzQ3FGSWY67fO20LukJgDaUiJ/TTWAZRXU5an2LwScSKXP2CB7oT/70vrsS
BY3TD3M/CY90wVpNtRuJQaXY8G41G1Ob+tJVGDiSMl4CNqjDvHwEG6uCzx1K
SmOPJF+9xB8une/BuM6t7WfOd+Gip66nExuTcbrsg1SaG/CkIn3kq2Rb6l9z
ss43fIae1AY3WBdpEK1uU0c0lj/oyxIauyZafoNj/9AoLhVwspHCCqKfmihs
y5mPx9UMH6/8LuHnmxyM16N5c09w8Ve2icFxMI5ah+KTuOaJZnejwhHrmBwG
2CDmXZ7t4SdJhbhcfYmIOt/ayisuXGZJ2zyF6zKQrcNGltnU3isIoxaj+g4C
+KV2Q+Js+gHVl9sgrJB+3oTxOR28mCBIjKXGcO5IoLKbvHhVCHZIA/37WKDA
A7uFX4AMoVVE6HSd6fqfA2bHE/wrGlmOvKBTKbKWNB4D9ZTwAOsNP4GSpvas
RPlgcR+r8HPiznhz3JAxAt1ihdmGznXKZrqNwze4J6WdDJFBOGJBhpx6QnNJ
ItU30HwkOBVY6socsTHDx7K+97ll1r2C2VVcNsvhiRysL5h1WPK2YRWhMREu
IoqlHrZwaZ8dp7jIHZVyFKkbvAI2pyW44LR5weyE+ZXX9mPRuLZhiiUbnq3O
EaCU91X8NRUHgdwWTn2ycC7PTFP5Hw9xj/2OXEQZh+R8YSTBROjHzoi/tBhE
5ssyPSEnyZOK9yvnPxIGmkvtYFOSQrOoPn16OLc859sXT7TcCJ1P41gjqOxu
ItDhcSqdeixX9z0jxe3GBJQApS5BASIu8WcvKtfvLphW8OT5w3kFyQbnlUp3
7Tb2BkA2gnC1q0X36qJqNA7LTCHrB74V3AFckDkFP4k4f1VIXqvoNAavfTBW
iBSkuFKcCJRQGIihwalfeR+0xx2u8U2lMmrs70ZJF588PMRrpH1Us6U6QRIx
WsRilYvcW33IhncXkw5h6KpmmdnUQkCsRmPyLM+vbxI4++4aP9lY6+MFzcia
I7/p5+mju4Zimu22pbwZpHFVto+Ud6Bt+I5/3HrcmRw/vvO+2WqYx4vmTD2m
cTihImYZ05je+N6YkLNUe6Q2s5+toxeZ0G38p/LRIFLwUz6qqi33A+SoCje5
sbY929Xi+reTfvOSJbN5tx9dE0YvPXKY+ioXcXg87KFwGhac21TROr5d0Ru6
MA+oJMjPLaBA9Lywdbwj6x0c4ScRZzlsWQVOaCL6F0FfvW1FhI9e7t+JcNsW
kzIACg+8s3sf45AoTi0VAtWLEXZ3WJl0/auR1zJVhZFDWlb7twx0KA3na89g
suREtPfF7Zt9N2XDdQ++ZOeSeKUcIZfxbgBVbpfc2KvkBoHg9gj3Y9VkGZy/
pIz2nEA/KxuetNZ43QTJougzIgZgcdTVPoXBFVCTu5wE+0N+iUWmyeMaaW1+
B4vd4GVZaQVWJS2UGVWQCANhpeI8bHdKSqbzqlVRhO2+CMMrca1MOWWfPs0H
aevHZpiFLcGMAGL5QOu9geqcx60mzT913EVyHTbXFOB60cU0z/+KTpQYFFvO
MFvEf4cio18VWPm7B2rgTDYey3OPeqgtVSZZ8zA5V1c/SKHvAu/iFS3JNaPp
UAIb/HQxT03/kw7F18oKw5XbJSdMyKzha7sJsr9RZ6kX2FeUXboVYm87ezTf
JdW4fzGF/Vzoz5EZyrlXmpxhZNwLX/NM4sKPqPkC6MBKBjXtvTuqax1RRxTt
Rsgv1B5MAIh7rmzW7N9s9EvxFw8xorz00BASDvPYEnnEsAihGS0faNyFG7qQ
thk16leLN8oBSMLD/GkfvU2emZmQkduyv+ZYYX6DEmj44ZIs6nHgwFPX8kHq
JxOEbfA1xskEN0IJKA9l2BpkZ7Dmys9hzMi2/ZJ2WECrlEbQcDsTdPmvwCKv
ivDLrGK3VmWSnB15bSlSprwmNJCrD2eq0bp7KAKxrF89F48wraMllrhjxkV3
fcoFioPmjTcNhFdwZidrqSVD8nGAGlQBP+5bGcexhHhdNzOh3fuF77qlTvyL
dKyDjKnssrC/ERsqafkPiX+kz+KMiAvZ9j+lulyjJsXOkMzHjcg+37rBsWt0
XYHezph/RK07L8zrlmJlFKjolr79eHojveNZNic91vyDhCsqXSZMTmsiOZnd
McCdOoiz7EhQLCjOTrQ80sX3KCrPYKaEn5Xqz5+Z5IP0dSVPwdfLvKOn2yTD
BP5MXR5D/irsiIohVkLzSRCXL1KtoSyL4g561T7VxyEt3hiyXuvvMcbeQiFm
MxtCvKtu2D+KkBqrJ3NUlOxeFUgcsJaIc1j/5UbNKK3e7t19eYzbeKdUXX28
BF8cEOzOtHQkgiNAKjGID9FG5kLK7weiqvRR9ZlxJO3yWu4XCNKd//8yCGVO
x+AJB8K+sa3/fLwqDGWvk4Y7JxXoBlP45Niu5VGGfSPQZaPMEXurTlJk+evv
19AERzQFaIjtKvgZS9dVfHcOnI4PIeYnxkKHfWR5C0NWnESjviNkchvHDHzR
sHO22KD/xmp9PXeezgmE900eNAYFD1uwAFMEVutpiZAzkg7PvN8/hRW1MAXm
wXvvhHQQ+yrj7RMdfxvtMlB6wXVxImmXugSrUKl0enIzv3OznQj6OlJcBui1
SwUpbXPrcVPKC9fVRQQTjQBMvWS3NX2ALNOWNU0+ul8Kq+jcJc8R8IBHE/Dl
Hfbni3DioY8LMdcvbC1p6WWyN5NFZEePn+kEZ0tsL8HPargGn8z6c6L+MmSo
6d+ABfgx2uNYUnE85xjSC9tJJmzbktvLYcH37UzVikqhwGH0uEt0Z1hLkkTv
7ZwBBWP9fIj77bBUN1JFnpxSI08kmfZqoh7tQOMnS/PfnAZ8G62GfpWEn53p
SSzssp5vD9Y5fSPhYBtnYLto+jWR8dO+0q+DPe2QL7rwigzG97X3Ranycdud
ayHvF+TvIjVdLlnXmk+7PtBT+vuSFLZVNPe6whyDXtjb2E7+0Lrg4P9eJ/cL
jaCEznA37fZH82BoX1ari0WX1+TzMMbS9el/9A/qSrra8jMc3u3xeBiIv1GS
AIIxokxhaVkKEtycAYX88MTEP4eu9urclpOLv6n1mVi8fl5WkvtvZDtz7P0f
uIYQKgKelE3QkDHghXAokZ4fb2dkxqeKmiPDHOuZMcAfCdOwU2AZCKRFBO8p
fkL7UlMg4Evop6uFt7X5BYNNl+IhvwiKtuXq4SzVIB6V2R4YlDE4Jkh/Cuap
I1FKmUO22kBuQ2XoY+Sth/CT0qSBy0WpIZDTVbO7BTAnF5LQw1abZR76110R
RV21iJmqAa2SzjtLRivxmdeT8p3hDdAVR4fWKnE1vUqivYu38+KizzteOwRi
Fetu175u53wZMpsvFhbd711zL3aS8dnCI+FqbpE9EKDNu/X+pHm7BoFosrup
M/sxi1Ow5cZM/20/Rn2vo1fGAklwEHTl3FlwvrwW234RUK022HsoaYSDo355
ZHiCwLzhxLb2GvBIyabLIsAJ4Ko3IhksAGsMWdACRhum9If6yzUaxb0IY0tK
YexXM8D8hWbQi9pvmocX7PpaTEDB65beKcTI3LkCls0eiIjyWw1II6PPDqzR
PB2t+l4Xh0Uu4967Y/X1pl01uz5EnvZru/zy1aTqdGf96Rh1srLN81f04752
lkVvUnVTICUEiPoj7E1rXXpd5eP6tZuy3g2wjNsdehNneuPK1aMYxNhP1kmR
jTQvjE85IkjodCL7qzx+nFf9suHJBoMUhPBe/D0h0rpLS6E74u0BPEiDsdgH
G6OQ8EOsAMfYBMbbroBhpsyh7sx//s/WNFada52eRgZugpaLkkQr/BIpVNdF
BVdgJIgYebAydFGU7RDl5ylPYKh0EZnKcwXPUTDGHt22ctSs5Ig3qachMj5/
jlyalKM7h353KGDhWsHXDBGGgq4qpmQxuwkRWvneKdfKxc3NsuRyL4mPt4H+
yJyIe+VXFRqb3yYVKCH+XyHJd0Y1YeYxf3l8ErvXadZpWhelo3hg5nxifHo9
smwl8vl6n6DKeLK1RUyKpAx23rbvf9NqTObN04wZ9UQHEoiibFqY7X6/atAl
A5vh3VP1LYjJpZ2bzF9Oyd4Chbw00Tny2VOFPyGUNWMK/6ttlcyF51whsQ1G
LVxHVwpyc6SdqnbuZ9rUVRsMdWZgF5buTvB8tyaO1god2FNCq119RInP1tic
T5+QQAlQHf64FFnt5y41nJEz6ggPSnSoILJucT9PIIGMMa+/VBUNwwhiJRvR
RXW0dwkFGgBnQ05DKl1b7z4DP1GWQ/5MAAR0alQIQuBGHs5nJcEou/WH5Yti
NNS0eJHtHLrGysdvAipQJQ0ShyHcBAeX12OhvF8IszqZ8TX2vws6FPaMhM3K
4xZy8sCnnIy5zKnvfIFFQCCGnZBRsZuli9hQym5tLhYQXPCR3s6oDnc0/zda
M1vJqa1y9PLosYshhWq5bBbPRBJjmIRWJue+pwiPErlwFJXoIu+p6fUBvsKX
25+xfAGiL1Qvq5KvTahXQz5mMQWxRfaX/IFuQPLYrWIIS8yopeCPBSXiDMXC
s1+377d40KOfUzI/hKeTmTqQAUHPEa2HLjqu6cbyWzf3kf1C2+wxg03jcCKF
SRP08HKQo+NyQkYqrUiM9sPzPJ193hCfSV1+L+RC5X6ivqulALQD+Fu2rJCa
MrQMynmG7PjCCHoo6detkpx0i0Oxt/HD2gu0BRMSsUDPSKAQxUu9N3dQ8cpA
v/XP0oEePCSbWdCgeqxDaP9F9Y8ikOOaN1YtrxCF3gnNNuWhhQ9Cda6An0il
bXiKxiBrDNIEBFCtj+J/kKA6zwenPxti3CdeU1UlfpK0pBHQ3Y/B9VyeH300
d2bh0Mi//lL6/1IDQL3x0cN1V8Kf3GAqAVqkiGB+Oufmc1l4yFg3uBK2WUdL
zkZZXEWBJpVNeCGCOP8IdgDcNYHD290VeGZDRAyG7W74Urrsel0UJSxGLKh7
Zk2nWWSvhotrkKdAGFdU/j8WbYGJKeNVF0bqAM+fc1p9hwjmiWg4NNABo58J
JSLOhBdDgaKc0OHUqXvXg+AV0C3Tu/bmJxznMKudWCxOGZ047V++677HBLl2
59UqYH4z6xEo/WUXyXJnrfakfkhkKrTQLbiMOEJ3TDn6n9+DTq6yCsPYRoqY
YRMsYu/I7QtV3SDPUJKcBNv44ItzPXujwqD9LqBOdjLtxsgt4ool/BnZkZ6S
LKn8YkwB1wzqBuXSegDDqrn56+/oyJFAXmwUK7+brxCrqqW2RO1E0GS41bhY
jsEdx41qh070lHxkx0astfk3BumlE8A3OUiFlk5SpBBHCFH2pR+2CQveFqBI
Fb1UtawvU69sAJwK7TcNuomrQWMvYN7LWnI+mCg/nXfEs9+A9fhI8MO/lozw
SmbNdcN9NyFlhN45q+L8yOLkCQX93HFkRKL0qCOIFGi+gsJ/Jig7EL0CEAcQ
Xr7HQZgO7bIpBOA3CRnAcaqBblXxp8k9l9S1xEqBWxPWypBIFLTdIU9msIGv
JVOFUvQGOrqnRCJTEKfnIJiQY02BfohIV7l9v7UzYb9iPsHI2z7JA7ZJypUQ
7yBLvInvzkl4LquoF/C0jgnbVUo1ULRPCy4yMSg+RZt/HbRASvg0XidfIU9R
5g6Rv9FrsBjkmrosz9bQ2veuN8bpL5p5J9Rbi2uncMGf1xtYojaaUj7L+S9a
a7SJ8XipC1ktV/KwCmTtXHr7lzM2kYGXzv0VdBosFa+Dc9hc8WHbswrh1Jaf
p3Q7baUbVFkkXuJ60VyncsiA/Mv+izw1jAub3RzpCNsFvCW2Q/PFisUxUosi
V7oIPUe63IXSHt+2QAvadv0Tv5Zt61j0LtYFCgM1MWTNT5eIo9s7DJumLxaK
YIBo37zdWKTIsnbvoNJdShx5Aex/ybx3YQS+Xt+bGc2yZX3MmCgrm7isDXwu
Wg5fsBPbZb+Vkic0oeEI/k/Qz3bdHSFxyLuZfgAR5SL98M3BW0p8OBXrmi0Y
yHrNI3cb5TH3YDM+0K4VjithuTLPUAgE41bzkmXN6lc7sjAZJDbpKq9KneTc
7SuwlKNCMGFjd28n42wNg8KUFJInefJjbm2LRhP5AwIB0QGP4ufuvhD/9OPM
J4ymxCCcpu4mIUGWxi+cuJ/qvjBE2PAugocl00Fw/KT40yCsZF7cexb1fH1M
an9PAqIXL4fTSz0LX3gq94toTrUZlpwo4KxSdrKOBtIhK75gc9FEoO5HO4Mw
BhkxyghH9Zv3nRxZiXVnZHvL4d1euukvjRICbkrxuHSLjVpY9phYOIGmAAxi
Ef6nPvBcEIoYb0972xHojapVn8P8UWEPu8CU8sxyDWXNkOFQ5fi11rJaDB6/
zswBbprHja+q54ZIkWvkjzFOl4ZbhQ73U2fXuOGe145fyQzsKpM3VthuV5Qh
mx9Ez89ijY5BO5PWBprltk4z6+s70FPYEUPXKtYJAzbIJ0ZvXtQsc9ZMZrZw
aTTc7zPDj2OScddVxmT08vSLDSHSk1qrFjvOKM2BgFoklCWZhnWNAH8LRQ3D
5BXt9tWnzZVzVqOf0Qk00IOSk4fd1trSw7+Dez39mzTtIrrC+vY4uV0gvS9G
5CkKNq7Gvs6BKj8GZRJGzSqhw29MGTjsP8QbLcr12myRzrBXnUcjjQOkDQDb
099oqA5BILkYTFRDgWlCCr3nvT2TB6ReA7+2gMWP18AARfcRTHWgPUNp4dEi
ZlBEWZk33BqLnandpNtaFkOZKbWExCX9RD81C+kxQJmsDJmVniVsbvm+9xAJ
zgVXCkYlMtnzFMAJYNUhE2IpNfIRbBDPLlUc7wWQaNb3nfuf1zXDSvdlWrFu
WpmBmXjlURehTyNJu3vQeGvmFHfJA8NyYLVUJdYe/NW7IMS6E/1ogJFIV+5N
kq3YU3gTpAXWE2il06XxiADwGzgDEYjSvsmH2vOhXWMUAl8n4evyeEddK1kj
fcWT8Pkk9XBnd1fOW0/MzZNIu/d6Cn1PDajHO+xmJGeNIxIuAPNsU61MiXfJ
n0dih/sj4C05iGTnVDqJ4xKd+DrXhHLDz5jOGDgqZoTA6iZoS7mRMlFS7sUx
eYUl4/5RC9IhPGZLC3dpzrIKnQhRsRd/lw0z4FkbaNk18Tcu7ntFUOzynixA
1J5zGrJ1WW0/7iYhbbSdV6axCCgwerA0dmcMZW77TL3763hdr8avBa9tabC9
X6BubkJshmAVbO+Vzy4toNyUdg6d5c02/pTqnFdMVjjLjZQ8JG71Ptk22h38
DnMAilDo+RFzmKbMWHJP2I4J5aCcXGInZU6cWMVBEXQljfl6NBWl0JXwLTpA
cYmabYTpo8wiozFp5j5q80HsCSV3lsQdy6696yOZ8RFzk9+O0GppiBf+/kNQ
IhBbqJO5WLXAF8FjXcPrlmMM/iyLvmPKU0vuuzSvZvkEZra1KFgsZO6jtX8W
QXqK6fg390yxNPKZazmlFWoSXOM/nHIwFOVOrKYtMOakdgtELvooWF36h5mu
/Q++7q+RRm9d7CSLXkJ9O4rlBkDq0Ykq6DqKA5yGpQze2zGahv1wHl5c7mnx
O+jSedJSvyNXdiNeJHPBCSgx2xH3ee8shjNwfHQSJjuM/UH5Dn3ksm/vVcnU
LLeVJ5rObRnpsjtouStc1nlUGnlsYKo6aL4vPTCztUDea+WMIynhqmXU3PDz
hOOr6glXlHLksoL3aF0GOroEbBWAC74KIyuwb03Pr81xNscuygRaDTLj6ZCC
CbJFlp4iWgFIVCvRHgklOimsqpmF9wgf7O4HJwBPHzHZ0eYKf6G8+lfuDwnb
ObVYy4DXG4yeV8+sCc8jIp1XOYU3ai3A9KhWfhJLdx91yrxTPloZ7fzqyoJP
F6X6+1xwIf9gyMW4GAFqL3Dy2FKPiOaIc0xH/T0TkDbCJeXC3P3+wODSzmMQ
L7SUjdd1Pah1okRoiPXX4Ap/wv7xwPjVAKclY+X1FOI/kAuvpYiAWo9O3jW0
EjAaHxFiTJrYi9d4D7mE+/9WHTXxy0I8jTZPqD9wAYj9H7FK7NhVEQ0OfVxL
X4yq0wGLqICpZcKOh2BEVW/cdGIw+b1mCt9DnPMreDhxRlcwYjMdz4FKTEBC
ewg0860P2gDm3iZ+RQ042Eu+Hy6b2fsxmnnkG9T5z2F2zXEbBWYDiK//FnLD
rwke1weJ7uUrYa5Quyn4WyOaJtMA3hJdioWUb7p3WDj6BR8fMK3gYeP63gCo
HGUi9PVyg6kF7GgQIhFJO2K8Z7teJDBFsVvA321HV99Ke4ffoE5tnhXZ0MvD
OkkTSMki+TAeO6pDe1qXJ2Qm4yfhRCRUZZ42BagR6Ji0naH6rU23B/hRhgPg
UT4yW97cQc3ZnUAfp6eVA3k8da1WwZLbvYzB2F3duuqnr5D/SdFG6OxnvpqU
dj2szAbeIHBwjnHlsika0eSj8MTdod7Zmj2othJPoWBgfQwxyZeYcBYdLMW0
FTr32+YC5MHIuVxmKle/GwZqNpIyiY+yaTmvOJRcetfZouOYs9qpDX+j/INq
awB7gBtBeT7O0fctcn7jqNXMdQLriS1VaYs6W82jaE2brPpCABImI6vJpdFo
8+DtITQ7KWJ5MZ8ykzGflWcg1WOJfv0E0yo0qwJlEV5f/d1rxv7brUzdAt31
BepudyAd2T7TTV19UM1FLfxKpE4CbLAhF6JE1gtpWS4VvVg1jxUX3SsybyJN
/n3TBVa9GkdgcTj0XY+mIDZFF0xUH/Ol6Mlf8sbx5q/bkLazH9SngakgiqYm
y1fkrHyXT6jaazaFiN8HC8lbcR0ab8Gp3rwTYb3Q5qKzbL0PGkSUm3YoHub6
gxbm4G1dvaV6hNz1vTbKwnxu4+7bfJbnnyvV/TRpp41zlpdCV+o6MyOcE4ND
DI3qznyYon30IDElpeizBaG20AhKCTOcBrvUhV1YwanOezYZ5qModqZBekfA
5eAb4RNcXIEk3yXjoEFiMjBmEl2HaZGO0m1NGAQnm5nYoVeT4sETeWK1Iuo0
EQtlpatW5J5bVDsA81i4GdP/1ZAdMbdefweZe8hqxKuIiNiHtQiEQf5WBH8g
d+ceoGP7DFhJvljPq3rn/unoj5r1PtmjgVlZr0PwamotRwoH9IbNI8D2Ncd2
S3zH+y5XVTXBIhVhFY80sy5fEd3wHm8xYN2S5Gks8hrYBj9kAF3sXxXmmWOV
tEdSeQM+IAGePUGFXYMNcm162U49vdPsdCDmnDVU7EEY1x50dUQp2hhFZKc1
NZ6DMKaa88egIP/ieq9cemIzCrlP57nXsr4lkUMOUR22WmNIajuzUBczGrf2
w/NVbTGCVAI9+53FZaB9fYSlGAeDcenyccLl61xh4ehhtWSUGIUgods4BBip
Bw1ZtYW27AbcNWXyhfE04i4pGgXUUktPjlAk6PiOhy676Lb0MW4BwctGkVpe
DJ+lI3rtlfxXZUI26fJ1t//rcYjMQzWJjJvj3tva29ixfmVe1KZrRBGoR6BU
0meyAIQVRHWnoXgdXL/lknKlcw1GxStunF0bfBfHvv+aBMZ4vzqfXcYcZyTL
BJCSvrAph8tHb3l3V4yQKLIopJhXDH07kAblOyKZHm3feyznqyiaxigmgHSx
8ENuHCX5JUTioQnEAK9vu1acFLuJqLgXhDGCLegdqKYVJdj32wTxPpqHyrUq
/YTjHDYpQVdhZlHSHyhut+ITMZSCKAYSCOFckcdu+2X5wVhDaqt9A+dYHrIA
3xJCdgXmNqikZX5Rn4UH8m/bnG7zDOJxap6uHXb/2x9EL/osPv2ojQhep19v
OS5Wh2bTYQjBOxWuycYHU10BIqPxL06FWIFgK3yHcz/7Opq61IIm7UUg6+ig
kEs8QJCVJGS8vUM536k+cr0aoXg9AQXdsmEw+z8pjZJpMIjqpD88TZVth4qT
m+09dDak75AqY+H1DlmD2OIQpsskDqMngtFlk1shpBFd18b4KXAS8oeojGc9
Yh1woA83xZuK/huEduLDXF+6MPEf3w348zt/lbHw6Nps3EZZAFfaoaQwluHm
MZGP5S47AERyQ/7gjBWOLzkDlHonIxQfMvqAEC3hFEvhyDvuEliEQCTWhQmi
HfAJbOqpV9UEkwJxXyfpdZVxxVCArw3UMYKJNJHrdpB0xalDYMQKf7fK1kx7
54czPKpbW1gs+A8Zjs0g6iYZZ2rCQo2JQ8CPqXm8C4zl5omOknZK+oMlK3Ld
rwIhbTU+LmGLF9s0j5ZoHTH+8MCFiY5CDlqs+5NkblWg0WEt6aV06RMYqMri
nN1PTabAmnehPApMJ9u1XwdUVYXmch/WxsTNCK5Cmf4W0o7n5VgCekXJTSnL
kYddkl2GOz3VcBL4ag2FVME4x7HjvF2m1lWHV5TGwODlno55YcRuKKcbCR0u
V6ZlHsoG7Gf5nqvd2QOdzb6FI3yfAUmnq4YXjY9oPWfhKHAK5KXH+Xbr3Gmj
53uOyTpTRrdKmlM9dnkQyP5JA8VUikCymSkkkMV4o30ac+/ebDroV18/EX15
FBVhRv3lbPzyNEptTuo2mcB9PVQqiHinBmXWkiHruqO2BbWwNcKptSsqQ6PR
tD0eDJftcgLg/BF4IpAGJcXSdcfYloxPsbGXbht3Ji0JYDrq9g7Z6E940M5z
7u8D6wqJrFkR6Gx28OSOGNlQWCZQmXIvYDTOCqiYeNoDnrgTO6HYY8y7Y5kJ
dm5ntgCInAmK1HqeTZyK4ckNpudk3pRTkoTnB44T1XA3J/4WQDFqB+IBuOm4
RDQJ9clBnNeDNfqN0bt+EeJoNVvbYO3wgwDLyFhBIGsDSAs28zfEinKp1Dxu
RVdkHlGZw3U5Lialkq2QE/pT1X6S4lkK8kcZusEIAzbA1vnZhl68YooxaPNr
/7cQbrh6YWITdPeP6Zw9nepSXH7BvnxGmUxxDlpUZf7uNOzeD7fL6H0Wtlow
jp+dneTsfpvw/q60CXGpyH356KotN7h1zCvbgAuPiq57ankMYvB6Ua3LiI9x
SVa9kfRrXh1gVxj/PByEhZtG+TcKUYs8rsPYWIJlPYmtPSY3Uuu3hrpLLS30
viOaYZuCBCRGb76fBYo28r9Ejd1n0asZRG+U0N9w84XicBov07Z+tSaWibyr
Z1lBEuOXqdKHQ7Aqg+sLxGlU+zJ8PQavKHiMG0aFCk6VvQlnLnivFsb/Ufv0
GryySm9D9LdX8ng9kl++lOIBjZdwsy/t2xeDiFS4oxXMQ7y1lhHUJhwegJfF
uRTEXo3VbSCYt/NrMQ5vM2oQ4FAEbyp8p26pehkei7JsmyMUu5R3r2TBHR9u
CzueECYIqXYRfFmaqqNiN4S4JMvGGi2+kgVeC7JfzJk/sgVCLXeBOBO0+fhz
4BKWvM6/FboV3QLX/ejrjw000MPCgAb81cce5Qx6rQx/TGYc0cFX2WCV7Zkv
Iog3jz34KVM2GY2jdrCHeCoQOUNU58AALlQF/4OwijE9pg6eL7ShvYwjhm6T
wZ8r755GHjxpOesyCqf3vTo/Xz6ixGIt0GnJhmbKSSzWEJIAGPQLsDTv/6kd
/Nz5EGX29wIOh5aTl1Qtxgz469OCUeY7Zb+k8tfWU3TY7B0o6I+Ec1k6zFOl
tYP5gg9QdWwgoGniJUVXpJIFjOUfbUsf8zCKxKNg/uvhWegCvq5ebqQYzD4x
aP9wtbyD1KI9KZ0EWpJdr1/QM//Qir6S3Pgv85WrCEASUSt+bXm31ly9n+Qw
ZrT63N60iuEZRV/czSx8ln715DnrgZPBjs5P+VEwC2hog4vRcl7vDq6pTYyG
apDaP4bXhlCKBvNtQw0XMUzSFaJ7+vkdMPekCYMgHhtoOBJnXQhaaVHgZwbU
SLEg90g50EB3OVjTwrK6d5w+n0png0D03hAKQpv3mLDtN8TrJ7whIbXuiAVd
PfkOwMC96ERakdgD2z9qBZgAbjlIuxnQ550IRL17PlEzJsMHFbmaTdVV9Xzs
ly/SkAZiI+ACl+i6qBSq5yOFwO/XZO4QkZXvDxM5LT4jyAS/l61MOPe6dOhD
OqvShS2CURZwBRAFSKKHsEOEnFdtsro2U1/IRRf3DlLGwAc+BKffbku6Ebby
DimeVNg8LJl04c2VGv6x9ftWbENrq5L4iDyrjmAw4++OXWznGUj1xQDHZeHE
+NlnZVL3JB77uauAOA+nfv7meU639E0FeWUSQ/JCFg+IngY2b4JaCj9rPWj0
eFwRmJdEmFVgjF/0/5j2KfeLi5Te55H1EJUMIC1z2K3US/3v8G/RtC2c6M9b
0ptobB/QSVXNlaXzzb24cw8+2AbTjIxMP5mxAmAv0C0P5VqvfXgOKxbK7CJs
50cqwO37khjzaEyQeHtdQLDVXAmUi8xLHAvRewkupPPGzilFjij4rovfXGL9
vssekHe69G9Moyp5uP00fMFQfUAsGa+jqKAs32pxZDQBZ1MEwnF0R0TlAZHn
UIVue16Fi90LpsjEssELfhgDvv2pv/UVwJu+2gur5ABpWDH2pTJFXgA25z3/
wStvOPkVXao3FiCBg6vxoLfT3sZfIZ5uWBkaiU3tkhtbiRHdEEP+Zd0AtKVk
eIwc0EI73F8eGWJuZ/1NiNCcA/OmFPWFGqOu6+bo7yuPaXZr3AGNmnRmkPr2
8VTggSRSp8ve7m7sf9+HvfjxwokfgWAyCwplT6Fxl2Y6zOS2hyJvk0MXATHB
C1PUlfsNpGY9jR+0nGR8JE8y4YwtAj2VyZ227pgUriDGOTaQrDq8dTbFq0nR
gw5wNUa8EzWFTNsg7StBfCr+EzgVUqsltJfQG5MsfoxXBsA0L4ugh5fMQAAb
sAWq1/KK7FT+IRxaW6AGa21+O9fIk7Nfzke464XbXgdlJMVZyYeUq0Mt004y
XEgm65e6BkorLGaFIl31RIKfxe4YEGHgFa4v0iYE75xhiCn4k0Ly9wwgq7Fa
+PzoeBFLMkI5OMCW9ZTd1y6LAE6OAYnw9kKQUE8CPN+jSQXmQpQUu5iynO1n
+D8bWMknwI07L6sXgH9V/+48N7UsYHCyVuIE9Aj5PAzM0DcfFUdXx5fcBmVK
llhIZ+lEUVQkqW+OLLSmrs0MCC6BdDeLQwdFmmL1EzbxbroWG9XxqFampvIa
u4WKxtWIFPgjUkkvkq4eiYrhXBpRWmh08EmRzK/VZi7OLa60tG44yy9SNJBP
xfwCoCPzTNZSKuK6qQ++NS4BJSDj1z+YW7ojtUhLtaFltmnZ06gATjqraHSL
jmztAvsGrrCCowxHvpOjdkOXCQYoPsHPKAfH3eDGRb0cFZGDGvXvNN4KXu6z
RIwQqFxI0Q4eQ6uGWg5lAyTlr+sGkNydrJrrB/XBUPXacs3f76BvHniI/CwY
VMKZGYDL+PLANCs6fj2aNq+FFVpny6/2Ut51tgj47RThB2Ug4/O8ScUrCtQm
eLhZyl5EuBOpra97LQJkyFYdihFCwiJEy2iMeE73M88eE0sddB4IQb5vdxuF
62QQEVvqTqMu5HB4FTuS86/SVwAzf1g4UzYtfsqdIlq5Hyez5uk9bnqZ+Nwu
FyF341+FGvzSOCp7qeZmP0WcOcRWvjiqmKfHgo1BN0g0d6+907hwYPH0YtHl
JgcRXXNN0WtSmboVNJWn9JlKEpv7KSDN+I6C4LPIvs2DcQClyGTvKfKcDdMd
YgeTCCy5KcS9hJavPbrb571qgXMCsVp6lSj09xCvgdo4xd67PtmUYXC07ucV
9M3Q/0uDnVjMyVQv0NgJjGCssfVBaLiWyVXi8yf1e6sTfhfPrDpgizoA7Vvl
rI87qSog587WQEJma+ojfrJkcTNWVHoc5gbSRRyK6KHzz9L++lspPqoYmkzZ
0d29srbzu+7a/ynKhQWspxCvVBKiMjrPRHLoZO/BRxi0vbXItsFtGX9wMDEQ
STguPQI4K+uRcD2YzimSMSMkzXm81iQET8XBWduQEwRS4z1NcAc6rbJuvRXw
Z7CcAj675prNRnEQleEBsSng1pZvpy4y9hFT1AbDn9YQnfND3SRSWH43snil
p196ocKaSi2lx+qTTTpUUcVTv8jJ8a0A6X1rO3pXTl9ZxPWu5V+TBiM1BZfD
3+9gqtHT+Le6l4LqSwTKUFlcn/Z0fs9LkH0B92fFuDs+m8+WbHdS9c1g6Ypu
EiHPa32I1y+g8rU5lpF4XWFMCfKKv7u8026OqfP4oGbVpZ4UZBFp9/CdNZH+
Jg3xA1r5MjG5IGnpK/zrfiwfkJ5ld473jE9Lu3tQ1JtyHeNu4rNqw2G1vVyZ
iioZr6f8PHHFh/2IFvy71vLJzLmGPj6Wq0AtCcKRgY7HVqZFOMZHyWjiEfbE
q6VNfUVG17F9vM3Ag++jdiLZk8FE4oVD0oywBl20hrZvtyMj3OLQ4dB/wPf3
UMAC12T7XTjwtYPiPc/tr2hU93VYRBu2Hy2RJ6pJXpNnRDwKEbhDGDzevF1i
iVghTONYBiaP3HqzKtJIEmBn2X/xZjoKnNTV4/GNN+UzGHa/cdmA4Cng4Rh2
BslPQjMjdOXP78H+/p+2V9VGpFYclmErJt9PtId5ryFT/gY5C8vJ8ydJFBX3
GkpgVzzaT+4SgmK5KfN4qv5sGmY6VysZeT9d54euyrHcnRoAtHMFodkNCUnQ
uohtvndUkqG3p5Wxi1m92+2v+3fVdZ7WX9ZyEavxtQDCfoNc/G3NeFcadWk8
6A1iMcFF13KewT062dpeavv+wychomg53xRcKDEMtQryZJ10rjKSy84DVF3X
9Lmws/jBPzJHHNa3T4j5VB54Q3o/Ic6i0O1yKFLw7uu11shTvTFmoJCUBAIs
hAr6qeKCZ8uVvL99+i8sDLJEZj85P5TJoKfaaCyBNJ4WBKnXGR9bPCy1xYrm
Fj567elh9n8w+jXSSAPaa7Lv8jah30GCVEHo5wn1Yw3RlmGlOQ1qGlVK9hFL
mwcumSv3EekhlxojIdDhkho+cVMPYdkEJ9fvAeyjRmdxAdrTJ8EyMqDYnrik
iZbgQ5hAkg8FQ+Bd+JWXdgp66hb4pJXJGQv47QgPUe0Sqs1z7ZbSyG5t3UV5
C3qPdN4w9QIzpeiPkTOjv2yWm9b/5DI2J8wbIwgZVfbudMiYe/negx9w9PwV
3uR/4Bv3pPmFBqcOSDPibkRSqJXB8guZI3NzyjbvIFkBmlWx1uw8O8fNw/K3
+bo9SKeBKgUsojDLn/z9UwabQnAAQ7Rz5gDdVbIDO3VPQikUnGdyneFoZ74U
WKFjL4PYRwBlZIgN4Ckrd2etBLjtX4uO/G+zA/SvEd3uxLNYU3mhM+ReOWmk
P6lGC/myQBplpN8tXiRHtw6Bh6npPTj94/WGVJzyQY3i1r3tFW48zDtsGb/J
R8pdTHpLSEPKe1e8e+HFg3TUNo41plk+O5sOHT4v0UmetNFE9iv2pIyvu/xo
KeXKPlc6jF4AjGBGxNK3AJaWXWtH3BdsT+/gnxHM4Ty6jI7Plyl2uS+pjT24
Cux0zDl8dUuQGaAM873YWeRXiZx2BoMEFqKZ41X3bup6YLO3YGpGgRsSP1He
mHCiP9X/7llAsjZ0ix/JUDHBofaKgY/Dqj0CQPMNxpsaIcxj5QlWzcnYRhE7
kbOlCJNPLes9TVCxGGlfDbqbAYjBy0U6KWMc5aHA+EsssBZph4Zjj9czDuEL
Y7SE0LMFfxv2CEU+WbQIdbhb6y2ef8DBOjnd6qt7jVfVyTvL91p8zUhgSBJ4
PxjJ2/KEhS5YrD9KMC3Mc305IkAwAN0huzat0tuAanNjiVnCVu2cYEiKoGxC
ATrX9T78FBYifpHM8WDA8RIzWPqj7DEGBwHr1LGFt/6EYVXxReB3VlETy0VE
vd3hJIFUYQR6/kjgpXTM+KesEXlU7yZhsLa2+HqtyCJKo41FbAE81CJZ//M6
j9dzxpnBZQiXn+rHMygndSEWyIxBiMcCplrE5KbTrfffnKmL2XCrU41v8Z4M
G6UrnF+wOPY7LEBMuJggQwfGIIWnDBrkKq3vBgLbB3XQWktrsWJGP0gdO+f1
dlQ1Wq5u1xWQG/DNpViG6hrE1LdPjidjzcVU6tpwtQds9idl4fwrQXYsBEsK
eS70g5Ie2ym36j4QgRk4SCxSoho6bglVaJBllzkhM17w948fm6ophJS0MSL5
X5dM35fqT9oCcsCpKyMniVsC/tfwDeccNFyhRizYBqGXx51PwS4ZTa5IU2ft
oE3KVzs0C4VS2VP4OIQzHdEVeFOjVOHeDx4hzuB3yyPg88aIETdOWuTaXk04
8VSfPQ7+P0rJSVmlgDIcMYONa+ukFSnbKdF8SH/VycTr4bpjF8TSc7lINURD
HvEA58CL71ShLQZ6OLsNg7DGW3y3o+2PtjuWpH0f5jii9lFHOegnXwhQ4LK7
0mgaCDS7XyFppxuEgQ1NjbumkK2mz229zrmeFMcmiiP70jnBOixQjXcYpVdK
ZVNUjjcosFu9DQUDPcJ5YyNDgdepB63a3CFLQw+6JrOHPkCfMnCWXxY1R/rF
lTl+9afA/CxQS1SgyzAYN9A8ZEKRnpznAbVJ+o6MsDPrHmf0COhBjr+HmTSl
O10hgaDkjAHlOLmKlL+0AxIG9697qeMXtQIUI83SPaiEs6rbk7oYOk1CHUtH
UN0HCwU7PzOtEjvRheylcErlGuEtqm6qvv3FFfq7Gzy7VbugdQlC3SWvS/Dp
QvYJVyB+WhV2/eWqTsQCUEy0q2EUIJREfQWTP04pdEaSi+S6nLrQ6Ge1ijkL
bpLbPQz8WfaZcf8QxNdeTS7wPmSazudOIODlaI11PyN/TtJxVBHftEriJ1iH
hR3iuPJm4mCLq4izwF4Nd3SB1j1EW8Tbtbmzdk4QsDiVn05Rv5arl8G5HKwz
jjhCtnLAe3oMc+sQfTWFy4jW9e1mUjiHstayVm7wcruFvpg2o/p23eTZ1O59
gsjkJ2neHV2HW/4Z1GgpZxoZqSlISP1++cw37o0LZQQXes8igu3gD/uddZ+X
HCQ8K1SFsOrrmrdOo15Kmwod/RUVxnrH2t4gMNfWtbWeLoodLntsvUd3frHn
yeLxSBTR0513+86vHiBUM6JL5rWXGmDI51Cg8eOo17Z83QPlW2oecoPAU8j+
Agq2Q7fWOR91ZJwhaxZqrgsdottIhMPQDAqWnRAFry0ZaWd53pbBV7pNF7qk
zeloawPht3tDaLD3LbW8wRCopsKGvfuIsbzFg3iEbC//15xUYiQpg6U4bs+5
BonFjBPkjLxXkggHC5ooXKk/6wWSVqm+Eb+d4YAoQjHV2Gw8JSMP3vaBhbvy
HezqEocaIA8MKji2LNOst+il82GK9U3hzFVYcQKGYc7C88wyXEAvDVvhgLvn
cym4l+Ib31xlhjxoEowlKCrV58Aywtv5iVQyEnC4jNiNw/AAP6/HZKcMFOq4
yEG7JUJJLnv/KhUkc+uro37cuTNMvRwCIQHv9fIC+l2B7O3pzQt3u9tizKbc
OHAxYidgmYTe+zuo9V67agVTJbV3rDXirfm7QwiEFURmL6OeN+jcFX3tB748
JZlDVMM8/ZxDi74Im4xxCH3v2yP9C7DU2FHbtLf1miGWzR+7jCU1wtWlC9dH
FXIoqlcu8wceExOzS/nV/8DV05JgZPN4bgNJr5vq+B/fQztvnJsoR0sNdYn3
kNbrTXbuy/vsJbqeYPNmRvHRWBijS1ZIyPb+8UWRVbbjpVtpUrFRQFI9h3hv
yDtm3u2u69GwPuTAoronMtZwkHvv5TDZ91hm84QIANX+oweEHi7ilsPBNV2H
PIzuxlvdVVMEtLSWWoPOLMrejkcYTt2gz2572WlSEu4c4w0SRe+u83XuF1EA
RimNNtQ32+R1NEDSBDoYT6tbZRUA3Enscq+OSvnhRfgL8mXV+nQ3LeZIIYuy
QBTbr0zw/5gBUowhjwYE08plMrrjuVWNPxlFjthO3+X3nOOIb7hVX950Spea
5Z9d7DrqsRxrY/FdvNoZchDjVducacXRBxiZeZUPVnli0e0dsSCEuiRX6zqd
Qa+YaktdZbBs+U3gp1FLcCrEq1RzyeMqSDZLLmYzSRYUEjKGGMlHnw8oM/wt
CamM74JutHw9OQWQMVypZRhrOUilGSbb4PPdqN/QZwaEg9xkW9OBneat93k5
wb4PHDHoUITD6y2icEQUMAG1r7AOyMM6R1YTLQBUBSZ6+EZCV7g8oVOnQzkQ
hWK3L0znBTfQeOLyWD06F0TUd/9xxgylOvoHvs73x6OQNc49ACUPATYuwSrn
XAX2z/ofMlCS0DL0XRm5XmLBpn3ManXbL6dDor1VJlqbK7PijiOp3w0aJU3T
wez9ltGGwHqpkSP+7ikix7ByJo1WWAiAVhkgEO5bf4dRhjrqq82g0hrmwk/V
Pzs7m+4DODSE1lMhAUT+/ZunejXnmAJMsFEQedI8jR11EbQZrQcvVnf6tQT4
RJ6mQkFDIgGWPlOGSt5IC2YgUeXAuCNze5pVbzLqk1hBz7LB0PiWT+JT8cml
wTYIvNfsWko5tAoE5JEhSdnrLTRO1zSF/SortB3Zd8VAtDcHlp+76tMKgtrl
pNamWpjQN8FyVpaD00tYvLRHE1ZdIXgIe4g4i7+qbOWtmmrTdMgBjz3uevIu
KP6ZxMqxiMu3wfZGMia1ualx1Bsb2VheRyI3ZZj5Nv/jMXyKb5Yg7MKj6dMg
z4z6sczWoXnGDqLxUUmF38Fv3IlcE8knIQtXijbOz+ALZW5hBbvQmFVINbTD
ZhfS7/Tq5ufTuISvQmpSuqgTXC6chshn4YTzcWrgDu3t45sdliuScBynsWly
483qXtdiPPdhmkZ/VKa4mWXYdN45HByHITAs0p5uT7PjYKFTuoU+Fn0hiIBt
ryu8RSxSpYlzezNCqGr0WGX6YywS0plT0DO88c115ZGyczykdy+4lvD6x+Cd
J8dYSkDIJ8K5O3cYxO7xLP9akZlgThz5SWfV3Msfo32RrP/IwzHD+PZNSgyj
KuAuuJEbBgoXAVmE0NX66VOnYqqNoxB+N66tZXpFDj+hao7Y4JP4cmUCX2nD
LModHlbpY1D0hm0Wk7ysIezcH7nA0eJ1Md8PXXRvySBK0mYbsL1Ht0HzSQfI
mNzvTX7yOZl8LtMC2auEQYwFPDEc9safqk5HYv4yOZ/q2PMMXLrX+v5rTP2l
LopgKZB8L3knlRpERBTNFgJClqsrx7SjbGSLxZzOyZSjd7i/kR+1yaKpM8Rp
KZYuDPsvu5V3fNfHB2EnF31DaR9ThaK7MjgaO6u0SqZ8aPYi1ByPczSq1Uw6
2XmjSXVX4tSF7fnjmcm6oStWTK0CzwBJniTy+g7q7Vh0CGEVL5twoFXEyW6J
qTZitOV3hsxyYrhGdnemVFDM+SamVdUeMXXOWIUyM+nKqA2886kE62fYUwPr
FLukWGK/qBr3jY+ofnmgTjcKlfpQScbyHoY0mm1Vosw7sq6NoA67pHotPBuk
rDrNXcOMuHxK9F1ZENldm8T3iY0DZUaEflV7STJkDfglg+62bap6Q/kjNWAl
jFAlmPrPPQPG8LUK+ZBiPp78M3XhHSXv/CcwrnVnNgGkDAtf3aUNXUTdW5KB
4DIKetjO+dgJo2VhwL+/uRlSZT85EC1N2F4nHpPGzvTgct+dU9DsPCLX5eyI
NficsU9LqCKM0Ozg0AzAFA4OANMcdxFXxJ34aEsZB5izCTjXgLIx1ARZnr9u
q58eEAitVfzraH8dZIQWl9vH9O0Me5IU4PZ+xZEqF/A5DzEnC8ctDOwW6huN
UEDCiCxRRktiUupRt7ot02shuKwhf1Zaddorwdx8CjCn4jaRB0Z0KRjmOjmR
rPPIJRHvA4INIzyTJmx/Mai+Fhd9ht7Z2tgn4vP8nrEy81F5RyPUlvfaMRQV
7NFPZTPEitzTW+foRauejnut8jtATfgMjE7ecybc1jEgcoB7eHNil1Xza60Z
4f2a2xeNX0xRUXHIwm4yW3Ze3Zme7dOjgB9uGafsoP0/f/p1tggGwkYLoF+0
C1TdNRZ6NHH4DiVU/owo7vAC2TkzY0b0plDW+6mAlOrA7iKo7Su+X0r4wYT/
ajwV/zwRHFwL4jk6NKy4VlN522X/CpsKNmraU8IobL28PrSVeheM2Ly0mISo
k7s+nxxXO0vvJ8UPCKO+lh3SKTUEfJ0OsetPjUEIs9jJkxHuxQ+9YNk5Yqmb
717nazF5RYu0mSUAqgfq8UwPJ4NTfbhHXt1gk4tgbu2RSY8bOihahkRwa36H
xUcVCDmNZP9BvA8Lo1I9JnOsM9ks17GCsZOpxWu8Wms+ZDyEcHuB/5ZkGE7p
QW0x14Gl7hzmx/A+bkQUQ9/Ct+DwPphXEnRUvcGZ3sY4RqVe9nSnZ3vr4fDj
c6shDOfRO6zrZpd42nyMsqIeHpMdAry6eSaK5pYvFRFg9S2wZC/esvDknx/N
hpDW8GGubCl4R1CCxw0qUDTu7ab4HjrxXZ207jgFDRah7orpCf+S3lVy1t1t
Z5jtzQicSASaxUicVlxc3mvDUAoLayVPvTiAXBuJyze3VdvqP0w+BotqqqVr
qby5xWCKq+fVky8cA6HRlLPm5l7YbFl6T/zUaNzM6E73k+2t80YOtiGkYwOd
PO8cy7sP/MNpkTJCGsvuQtgs1d8IMWXOvDTZ/AmLTq3oB02DXsSQ8//qDt4F
7D5WsIiYIbJZrCTHuQhc6eMDQl8TzPEruBjjveJ8J9aNCzy0i0ciKATNCfvf
rQojPP8VHqL5iac250UPE2PlxwLYvD6h8h5JzI9YEg/nPwGHRjwioZMQVUX+
GyQBNC55l57JaTcGhCYXaEoZLj5FsxNXWVw4d9oJa/CA62w3ZGlvMpE2VtJs
exDftHezk4dgac4+EOkP0zy6liWVnNY12SpM3dAI5PwNaNmwRgE+H1alPxYU
R7Ymrjia6sGAXP+wO1Poxn6vqjdnFvUUOVJx5KBW7Ck4/OuyVX4nNVja2LMR
cidjSAqdNMSXRpSFN8VljOk59KOYDD8civbd7zEBzjgAjrrrcIgm4+8dOC5d
+GE7URlBrsXONYkH5sjNW9UqCqTHeWoB716pRd5rWWwZU0niUsUek5ixWNG7
ovcGN+u1k7tvyHFDSRQrX9dBiJfeYU3XEkVlAOHap8ld6fMWR0217rXFOlOt
RWFglOmEq22V0AMygOwKp6s3fFIAxJz8uGN+Yto/yQjC8IMDnbYwA1pEfh3a
pfYVU9KF9QJb4u8V6bdXEJyRQj/Cl/QCRzmRX5jamMG/8U52IcYjEYU/WOXr
WI8vWhSifymhtd5gn8HMucI5G20Df3Fpe/WuWBB7njpLT7ZpydXqz6qTm0ZO
E/Fbozf/mT1g7DkyMnTNAwfuKizsmBJUWepnvyxCGGKSocnuuxwe5TgI0oHh
f84L7viOIYvK35qZAv5kjq9okFXeEThr5+L6X2f3z6+sRiyx57/Jt3KzHrUi
lG2MoEx3dUhlhnOCHJpc1K7TP5RwrS5sUskl5GvSdhZnOP7IhP231z28cNmc
cj3mGM61oIHKAi2dsZSWjgQERA3H2XPSjBv3Ed2qqGNHd9+lmReCH+Czsttx
z+1kJK6lcZCcvvdtZY2+wEBi7Ifiek08QO1A2V8aLk9xdZ4HMXUvLSk1jfN3
WlZZ3lTlv5JkxF7T27keTvUOXhb4DyiXeJdaclZ5D+4TtgfXmgJouxRTZPaG
QHsiNZ3iWqY3RU+1fYwNYpKlLi/MJAWGgr4cCgg+o9obhwwUZWnxtPFbMKMR
/Ls1c8EuE1PXL8JbyuSqTdsv9wEN+4k58IxLf21A06fEfCsSAaBADFEZCbxS
Fb97aHNILIGkbo9Hbvh5ngx3Qz94sAna21zZyYYGthog66Ga+GBdl6+fFMQF
uyT13Awjf5mtAfId+OsQaLLsPMuoK2h8ekzwTbIyB4uT8KInwCguL3Pr1Lo3
lMFbSbRBT9iDsk38VyevKVXgd0t9FtyAom5nRcUcAn+Y6DzwFK9UZxsHSj9z
MFLOurOxnEWlWXBhcAlw5jui5tCbAGOKwNbPEo8gvaMk+QUxlCi6akRWmCt3
frwBQEFc+PxEHthFi5K6ZHDAcaiU/ILfBipw9Y0Y64UrcdJpZ9DNk3Cwo95h
NcqBPU/BYSxox2X8meDWiSFsBOSN2qm3P7At5kxWnuMl4iHvLJix2nid5gSc
1viGXzL13W01KN3WP+OnInXib0cpcgET54R3/oeQuBRVl4cLjO8X2CSOjlcN
nKuOJjpgcbbYVeyuvmQr35Bk8erURBlMeE0EKUUarQdL5nHN2ocE4S8MdWVz
ev86WdW+1rOW7lH/a+cSXngb3/wcyE77YA9HD4Tdh1p+tnKzjo/FvvMRy+nl
9tmmAF2bfum0FROwW12eJOZSjucus+s2feNAKTAGFGfRIUsiFLzAOZ1puiML
qzlLCRpxhfLhySSssmAYmw/6KIFgkC+E6FzUyLFwJ0WGqdAKbo3T+rSH6B5Y
dWT6fXcHuFjdew9Gzv52omcsH9m6ia9VCY/BRz9HSj18JgiLS3V1GYEqc8FY
P42QpKC/7ND9sZo5FhriTK4ZJihDxf5FNKpDireQ0ELtwXQalIiy1hbNzRgt
wCCDW58B4lkkeqVJcPYpXUm2L0D4Fk74ZYzFtVMYwFinAwQyIYi4TPTSGUH1
wsSp0rZeGv+jxHCjgDPA3CZDnQKW05JuhoyfhuWWbZ8Yd/9rRRGSaB6iHqeo
fcC6VVz3gZQxejKt6eBt1QOSvf+cQX4bilDgrNrVX2V10z+DT6x6TgUcz1n5
S8EmPFy0jvxWl+4U2OIsu/C2FKMDdtLulv+9fGzuOQBnXRBPZoV97AX7cZeL
h8udsnMBX+hecAUQlg5i5/i1zsoNH2LSNAv8pKC6xxCDQheCdAW3hkGEj1BU
zQ5koZem5e9HtXUw67K9YERiuLSI6E8dHAX3+DGajbnGVF+jbiVoBW/J9/1i
eAHtPGUAAL2vk3Xbi6PeaddlJz6y60VgleDnOuihHKqRJHFZrddgeaeyjraa
vLNA4odIGOHgljVmOtiSQHEghugu535S/jN355M5QGNnIp6orC5HoQ6zwFi9
iECzIyb6eZ5z3GpCUZn6c5SDHRYbFYLeSz3qx5F2JOfuN1qigtL2akhaWCY5
cU+J6AB+dKXxjKEdTv+1Qdj8kGIlSLrEutTT4F37XBkkyWLQIuWhQnsfjiRJ
ZVMTNNdN0qvBOPo0vetV7W6a/tvgTrbXwqFiffmpiydXmCjzyNF0G3Rw6mgU
5czsVQ+OhgxoIlepCINXzyxUDRFeaW1wbRUYXfQmiYFuJMYNEOLoF2zXBSJP
dx1rey810SOKp4a227dcGmezgg6HQMziL8VT99ErjNSpfDEmeAKd6ajmrVYF
Wetg467kPxiqTXw4J9DlQBkv1tV+NHEbDyjjkfveXO9UHJ3cVgj232dtcJcK
tCFZjKJrt3SZ6Lb3uNRvodw8ToXNLyNFLAg/i5FW01gNX7s/L96farT2wJVQ
YhTa/FDj39ZdKXapGi9E+7W/lFEEC18O21rpNVdwcuDjxyAD+akrAKChaCgT
aZnUTCZ7ZUY4jxbuOMznO6db2dy+7k7ZkDbd5KAsNaFGDMwGyK/c86EaZ/cc
VHJN8mqNdI5PG+YcmeD7bF20hb2vTqKFBMwJO3W03yQEBxP6c/575Pcyuh7B
nDbp1WmmamcB+CvrBeJfLw8N0Egcgo3M3wr+RrmPJLE9sRg6uJBADLxKdwnc
s5JKgwFKM5ZXNP/28q+C+8KZYBWaAZO5wuGq1ZGx7PEY8GanGKqFTCxooEN3
Ih4vp34NkX3NR5fFV3FticqIeDx7s5Co493ABGm1AqP03JJY7E9Y/YUGei2f
8iDtAzw8WG8Byk8CK9vOk8XfXLaZ6umXs2K3R4ouAQB8qrVt0J7rM3khpD8G
a6tobfmiDZyCxzIgOXBEY1x0egCAaf00mtay+UEn/hlbzb2OebNx/JALx2nJ
Aut/G6MuEfTUObT9d/2yPElRvwMyI3cNqGAppr1Ta8gwMAx0R9Dk79ELZISq
B6uz6A39wyT53RliekLfkoAhmk6gRvVDiz8vZjUT/Rz4a+s1ZbPUfSzykDKG
FS8J4/x4lZF+GSLKT1gEWwCvbxe4FamW4AZw+G2ZrHda956PK5HsGA0ASvuH
5FkAvo5vkCs0/ZR5K4KqGdMT2GEqrvUwq22DGSOfVnc5nJ528yGAIf0vVPn1
3lTnAZIpIeIoJCaxEx7krVCiyb4e9NLLOm/t4Q2A0UYcOECaLTTTkZEmMXTa
VAfQfU5rK6yr0xyChiAJOCDNEdWWqeuJAxzUDZ6Etsq57L3cKktNGFhF7GH1
3vRUrS/eXKnvD7vVBv2DeDQPk9wKYwUv2xd9F/edwXS0CbogxcGuZNaRRWu7
1+v+dSJ3noXKLe+gnGH65JrvSLJ1zKFHosUWV25qapmngHpXb6F7sMh0pBgw
YRzEA99G5tl0l7L2rJ2aHd2CuwqEyqOkll16gtmBbV+/SVgEFhxaY/IfHatQ
WNwFK9uz2JYfs9G5T6TNwigEa52Wgn5TXCFUd8BAwEK6hoVe7TkgoXniHG3O
BGU7RTeqHqj9p/XqLGzX+mST4N2EDhjxo7WyD8G7kq6BqTtjWJGzR3FKYwyH
O6Sphytr+KuA94H5uLrfkObcQw919Tp/nkdy3W2YtYZ3eC4osMoyh+Gd1iHE
cZaw3S7/tCI/TcHD/GSOTVnml+xlLiMzRRd9WAXU3LswUio0yQ82CIpKP/vw
aBqPCF/vgo5IcGbVqNkQIMUvBReO2J9mVAztwCq/Lrj9FWzA94nMt58XiaOL
Skxrp86hdx7NiIwU+NAtg1G664L/SnuBsNrtsRhdaRJuESuWLxciQjCvPtCE
+DS8zmSTxGSSRfgEXHT8V6d8ksrLYDnIYa6LpaJKMiJEKw29OhClU0Xba8aP
dEZ4frQkR+7r0vAS47uma9I0xOr/JL2+dvkvCm1IeoLOc6oJ6oKnr2rk/FVT
2eEVRY7GI5lTlLUWo/x+g9wCg3fMvZl2BozwjRZErC2GX0QDaA4j2JiuhjfH
SaZzk8HCAk6JIpmSJd4abZgV8W/UGCYQ0+cC62Zkih1ZjXAUm21aJwsc+Nak
X/q9qMrmSD8bUSjLWKlejrZtl0PIBLdMSHiNSS6AWRxj94lGWFfratu55pzl
Y6hBZrC1Sx7kCHjcisaFHm/1D5BGtKvOXusm9AQ67uZRtVQ6RtHjxqNsiifI
DG2A26iwU0mAzzD0ucxb4yKkyvkOpfALTz1LROvgDjNGhVJFWKhVPNVBcA/b
MW+fPhwrKWkkP3qMcvYKzhf+WEFIL+70Zntwb/Man3Uj6lO/i1kRmZS3fvxV
nYxkoOg1g4KVlaw1rwgGmpKCAjPCScIJHn9BT1HRLXhqoDONgXOmHIRh8k6s
K63HZRBs+XMdWrGG84FuUCBpkJzUcepFFETLmZr+PGiRaXIT3bxk6HBTAvWL
rvwXA1rPFT9C9A2qI5/McUS87q6oZ84ijFog60MZdh/+ef73/lm7xYmQc+pI
pHPcG/2ElekcSFQ2CTaNki78hghr5ykjcTX2VWi7YCXpEok7bbtC1lXXlr+8
bFS1ET5syz608BP6Kcy+68KlKaJaQ80//GstBBBCiLe+8q1o2M81P3PKqthY
tyxxHKgX47Hj6RdUGJ22pbLSUqNA32mIh3li9xpoNMp0y1/rVIbiKrEZpudq
01zo7xk7v/OUQMrcT8xGbphRJSGIqsVpD3P2O6uFiUDPrNjlxhe1durIQ7gh
V8MzwML9G6P2j6iDsLW1TFEsQINGZUqiEzBybq9T7E89AYMMp9SA2IzSuLwA
qdtxT5M/XBhO9jx9QWp+KfEeTSB965v0flK8t33QOrBHsXjBXSY4MlUcGgKV
ZVw4Ztwevxgq4fLQaImzx1xXLM+Xh49F5XZgGrsBzw0iQ4YqooReQqIdtMKB
9kkcaABPf9cOMb3FkOH6Add4O8TICWm1styBepmQTY1W7rksciBy4i31oB7E
4Ca6p9GvpZR8oFUQTnZxww+PyRfJOilr4U7+NUFwZVxg3Z0nNvpO6Wnz+dSC
JbcQe2Yjt6nVIBe1/OZTbv+XnN7C6YfGtdxpjclusC/z+Xh2kbZJbVmzKfQk
cTtilAvZss1rWFvJSD8Obkdh2lx2G/dBfQXZ3JZutIJP/rZ55jocoAf6t7zX
XFpCKkPQ7BZM7uxYI0ghXINMOCDmIbGvWIbtUEEGmLcQfA2ro9Qg8keG4xaE
pKa5Zfx9atfTcX1+1+ehCWS8AfgnIfBiwrMPfxhPYOJkYI7GyhbyfFN4UJ1F
6fOMSiR3Ae0kyUHdq1x32c2qae1EC4oOWvV/DYDUu9yz7l/tF5RAI/u4TNO9
WMWCmSZAYszoImODS4rpgncmcS6F3AJ9pOt8bVvTfQkRdvOuJGYGWVGzPWgZ
2ef35b88vAvI4ipTY3omREo8zWDZfsWEq1JtIk6HPbVqk13V8agZh9ycdVqT
j/z/zDfUeOfL1skQyQZ4HBWSNsGeHXO/8zrXSH1mnZH4FiT+OG4bdik8aI3M
1WOO28Xs0YjRENQFLQjvyD2fcnR7gvL1jSC44306BEYzdbJ8Mw8wwkhmEfBA
yiRrZn9bG+WreMOION+aiSw1bipY0LCP6i1iinteykDpZSwAvTiVySxfe918
7Y6GxPxWSJCftazqBsn+ZD6TkLybZDBS9hwzhs1KDRySgobuHohsXWezjrJF
Hd+U7xIfm0ge6geA0Ip1G0CB4Oo/qPoCGDZ9VUvxrUuGx1nsdSc7JcVdf9F0
PvyYmYxG4x8ZzccKrxlKAWonHf5+Z/luyImVBtApGNhSOAtFnA5sZTbFV8EW
HmRvJteT+r9FGzp2ccHxyqfpa/yykfRfnJEDVefq+27GGKGJJnqCpe9Pu8YU
shGbe5DDbhIaExbB52FlrpO0kWDmeZ79rp+rhWwAHMHi1px24d3foUGcZvFz
QqP/IJGIQXJSFhaweTiMeLiBT9x7jemIQrx4fLGE7RvtvQujSzn/cDHm1IHZ
vjwzTuNlOQBwTcZlwFV8vJYC/JS+4GHDm7aBewOrO3OqDKY9eC6IFkvl9UXK
MzMY3meqCJeMBrGbpcVd+DC+ExY1vGFWsC6giyMz7Y05gfv67i+63BO4XCMP
PM/7/AAXWjO9+N7ND1sHr5TRyXFJlvBQmu1tfI1EfvZd5UfiRHkLAmivbeF4
6Bj7mZIN0kBJeVF2iloxr7MeS8fKzny0CexiNRRsWO+ky+GDkSYb72jds79w
M+G00q4yyDKqF6uSSdj0HXORxVtmcE+QxbOYtWgMuoZy7lH42spv4J5m9hVP
89ljiIVB7C8ir5RcSqLTKXPBzcOokL5syUPASfzA0B4Mdu+th61aNj58LvKH
lCKb6qUNEfxNYYlCf7wQWx5vSmHJPXXb/MNIed0vHTI/dlDHzzFJBjNyyM/Y
Ee1SV3W+b9LFoVRS2IcsxpTIZDcG/9kAynFHNAfZ92n8c1XcD+4ZofurHFNZ
EIP8t9vZ1OBjk/hbJl8m+VU/Vq7lQ5sSzBQyHZRlRZ6B17CHRjT08vFX/0M2
lqpB2qZfXoJhFEsOMlkS3DCjqEdizxQ9KDpCTqqLQ2Imsi3EEj1/LsDXlfFB
12alOXgTwa9xOrVsJgOjbX9qPPjx/XtwM08mkIEXZGiGFEULNthBR/IHzXGv
0yuedKDh90MU/QPAahAm5xbE1xFjJONt/zIgWo7erJ97gZIGDzYcCxbHS3Yy
I/Ghsiyr6OvIBWVz2e50Zi0+JaDztsz0IdDmspeB7+3JNxn4ZGVpN2IqJP3x
dCYBKi3RrdoUtX9ynbmuZz9XkJh9lUhEOK9/OWsGyd3EA6SWmwLk2ySND1Xr
pp6WSbu26ffQi9WR3QTnPQuGpPIv425kyRHWqqnQWSFDDOhqZ97aOI1PRMQu
aMdP4YJsvOrFysEx64QneC1Ozg2ILRqFQ38VdfUXMjWZmo5f/MrBOTnHMOf1
GWY8/vcnJrmCBW8P5YYmmhv+ryUmIXpspD1l+y5daLQgXdpeZnEw1/5ZAp8V
wsw0HFRdarkB/6gSGFI6ULRX7z0bH29O/sljV0ZeK4Vauv27IL2eesZaCwe7
MG3dxpOoEQLkq/ieBI4iUogYOURkJ1qFK/r+PkPKfVUf52txKALBvWE+bA3j
XJv2AnzdGJfdeYZSTW1kLKqfgPn8tOybdm5/5XTmqtLGEz0nrszEZkSb/Yqn
HZPMZoXHLUyYr3akBNDnAyXMruL/J3r1+JP/ltbvxCpe1kEQWgwqRm2OABJD
mvGNqishqDya66BkQZE4qZ2Ub1cvGJQx0dDIj+jE1oHac+zQm5VSjbe9AOYD
Llpe0YQRmnM20YBwASECrrO7lbp7WGlm0Cl+PEu2l1i3XFYQbSXGldXT8tyB
KDOdk5WcuTRkGQ0DIJ1swI62ywx7V+I3w+Wi1GzAo5GgQaZWPToq8DsnJLJw
rR2BpwOGLToLcpTgB12YbxoTVpqCbqEZMSicZMeDH7172ojCDk0VY3+FfDO4
pLA+mLeI9b8P2Ld9wpWA7fjelZfi2Vvwl/tMENzitrT7c4dT/HF9XQ57VuEm
3iEutCopax4ofvgXOE22PzAIXlVlx+EQkC9FB0FqTIqKoXbYg4v5QrLY+171
DPW0IF2Gv3nFeGXhwTvxwqvMh7UmfE4H98dVke+tvkSuULVtiWqxr8ROCumS
UpvLhYc42E04GgzUwkFj2ih+qHKVwuP1cSqlWNTLkZB0Ih/tGq1dy8PuegkT
9VnRpc4BhM8rf/K6Q6eeRee9NvhZnO4/dpe4XFy3N/exBToh6w6h/D0xtBv2
ix8EYEeVo4VwmYUWIpVK+e4+1osxvPAfymGc/T97vwKI0ofI49WQqz2g7dFp
7t19hWWcTYQiP0pBl4IH9EaYI3b456SkIHEfNTRFcpLflkbwZsI+FI7anVq0
Y24AMXu+Il9ZVlWQev3gfEHEg+PdHzl/D09MDLJLLIN+yNcv2I/BG4v2D3tU
6qTB34YxnlhlHDkEYrv67R0RLyFdv2pdYioPU+vNV/pvr8fJrTYlo3vF9sJX
6ScexOJUl918vmhta35t/xeovFNAqDS0Hpz3I0D7dOsDkMurbGCTALu8jwHe
80e7NbjMMJB32oespLrd8keViGvu0aUy9cakkD549M+tpoz73kVGYC4+TXTs
oYACYmZ/a8SvuOy916d9SGFJB/ocVyYyjg3IGLDcYxEPw6b+hSzc+1kHmg3x
8jhSixWyaiXWkROg/c/KfLfgYxc9S+WtqiFfugwVDnLTkJtDHJfWAZYGqujQ
K9ioueWNSdEbiDyTCB/nq4B4IJDFf0nPZCFUrVFaFvoDvY4s0xb5NbGDctqH
ocSOEHaNgWUCYvDPd3akQlW5iL63q0aGkuOS4AYplFoSxwjsV/3mP4FjqcUG
5IPHR3KgN2TmuGo5+zxbGvbL1idmK2/EkG8/eqV2sczM22ok+KxDmgRyRiYG
OdCNH097ULh600AnjSbImOCTC04zXFkShRaV/Qo1tSKq0EDQftlsF2Y1wTLG
JY2Dgj6j+aicQRQsRe4uig2e/xt3ZnnFl29O03j+p687QodZbMWbvoCEiN0j
Y+N7NPAtGi2/ZsI3tdQm0F2eJ1ydxLZzNv2IK4wv3cZWYNN3q+xGwqH6oXT9
YhA+XQ2EjpLKPbTjSXDjFZuKZVzudX16lOc8MUZMPNnjinpxfDCsYTNpNL/s
DQycImVF7FKpomFmKkZoEccqIYmgKSuh3rlOc4w+dbiDOPCi/W+ONuq5D6x2
zu+f/VJNPsasg7+k+U65RRpwTyyi3GGlkkIHVIl4CeOY+QPbI2oFkTsAGv74
FDunKa3WKxx++KgcQeM2wMmGTz1e229ZCM6Zo7VuaMQMFyBurQnLkGmsX/mb
S/ITgFPyJ9SpRu/SmOrRIRVwxCZbV1/iBAygmArleyjjXn1Ck4pxDoFUe6G6
9lsPzyogPN8wC3AY2yMekEUi7UBCG2LGAM/x4LCxHXsPtS+NrHD707a9Dbs7
uekqjJ0r2pE51O65CUkHysU2DwxGRezhoJW4FPtEQjKncH0iY9gj/Z8iEt5z
G1R96RUc1FSBBcQk7WBT/n83e5CK2F5YHShb4N/+S1cD+BEkM/bAVRbThdVi
iV4zcDGqiBlN4ISp8pfhvCHemdIs3Oq8iQN39wCO35bPGZ/jDhsv99dJo9kn
KX3d3GW4WI1SRWwQUpCjF6PGVvWmFi4kNxZc73Y1K71pb3QX2FJMHryaMoaS
EwtS5AHZ5anZ37LFclA1ylipBtDSKID5YaaDaewJpIRFo1xUI1CyK0DVgMTl
mpmZ3vcH2/H7hA/EF5wl1Uwp6nG83spCGdKBBEFhiDQaSqzhn7ObJMuKAsRg
a/wZ3d36O3zq2JvX8eDOoS4Z+x5VraGZXfdyXATErBu7rxzNnjSzT1v7KVZm
sJTUityi7i2kOXjutjuyRgGzj62l9TzsXXu1n6q/wEDU7F1NMBEWFVllXBBS
EBX0PBxOrV0GWcsR00OKRtBtMGesCUoNU6jhoIGZevPHvkSb5S0uUGPzYqa1
pCnF1NBENof6qw5zwuPIjJl0PVzG0AAnYh4vnrkY3he0BOXKr4nLBlqo7IAu
+sDAnA00MvcuVH6zgmRHISzxtvn6MZq09TGamdIx78lUmhf7op+B4Yg89X9T
qphDYuM1MEc8poE8sLfyOcz1ufsAVS8HeANR/AsHfZ0YJo+zX9IEQy2Y2dLH
kcPUGVyIi4M7QKrZ4eeMVimIn+gL3DzD81ed+iHr2fK07qA173IKzmfcIrOQ
r6xS/fTUviZynqg0vyKzLMwmJy5wZ0IqdHZEw0Ap0bIV+wDBCeVCIBgTZBPv
qlOZf4tHzgzJxeuDIeIiMaaFDZwNbCmmI3vMmBOiFuiLIdxQoovqBweJvJVp
dTrasdnhvPcPFCM54plylyuIZlzjMY9W0zLKT/1jf0Sd5rlJOI2XL9jVZTi3
LxN86yeXX87uz7uz11EyNP5FHZHKKwy9azxCnTU3O1BGw/ae1omYv1XsD6lv
YJ95fkdp/e2VsM+JzRAEIuGBRHlkmQukSfi1bmxXgouzaGyYRFwPkVQO4sjP
dakj7hNaADyKT9qWcg8zpSmPnbhBXmrMBxYJwLGbAAandInGfbvhCXx7mLyk
wRi1kAyNBctfNtL+SZznPK/5BqvVw2NoCtHvyb0TfFQUmWqs9RyUmW+zv8a1
Bb9Ajh5PVVsCT43Yx1fbTbOA2dS5L1AEEjAFLh5nx/8zy5aoQLVYVh6UM+W3
XHTCwN9GcKk2g3ud7Ui+r9et8AF2atx49ptqedBvk30VDNkRukkf4jn8mNFQ
onyDse9DoRPZHZ73Z4wHxtQaQFIbKSorJjDejOHRDYvnA+nYXA0k0fKwpYj2
qt+iHCLyKx5IZRAnKoR2DntdA0KPNQXp0Z0BuCJwbPeItLNakFwOtc4XFDHS
PjsP4eLmWvAI0Np0Rz+qxIhbI8GUZIDA6bYP4AArYECSU6g0oWpCrD3RzhBA
FmK6Pt677U9Q6b3DqjDCeAqxLMzA5OYofnO1w8kClP8yxnYhqhp0A72TEoz3
kSkSPVDH66qiCDPY4oSwsDLGu3Hd9/EEqi3g9Er8kousMuOZnZsLBjQj9pUQ
tZMLfRBHhjusKWCy2dY0Wb4yHa5KcCeVE6hEs2QQxIzeDbTdlNty5vH+r5wa
JjK3zcMjmx6b2JacXIPWf8m8pLyhbgH1Q4t9TaHRRX7bbPYOdXZQuCRcwLF5
khQ4cR8zo2RLEORN2sb4rQoCkHSHnsD5fXfpolfg9ZBQQJy/WYS0YDKf9iFd
INx2xvjd77SlamdDTxAw7CmpAfVlq56UdWt/vEEpv4cpqneZVkTBY45sZPZA
4ry+Y5RB7LCzX9/LXxMOKp/Uj7ia2hyaGHCcTb2v4TI+vDfRCSPGRnNAvnRq
Z+o4rcFWzi1KtIRHUdUnO2aA5n6llD57aJqIst6x3N+06jkjCLymTe+gb+p4
ZaBHIy0h4paXjnitIiKQET9MSiuDwXx+vj6rHmrN54XO7EkZDUlep7RUeYY1
5Pe5IavZoSyUdt0khjwO/O+Z105OEpB2UR2DayGhEhJ0IfJgjDz/rjcsZZL0
MLvJwPX/96Amt2m19I1VHDHmQVHVwNaz8RasxaSlpixo4bAFhT5MxAYSjiu1
47vjmnp9vD+gmZkQS+stV6uTnHPKs4m6Avx9tJJR6kMYIBsLtN/wAdK21UUr
2U65QGAzrgEhtoDHAaGj7/h/fXkdisFx+qw/X9x8gg9i7GOdQS03O+0aEfIP
oGHCBfZWRgqngdc5+fAgzi70lnebAb1PJ4UJqKSHKtq6S5F/FdzOt2RC7dOY
UjxHGmFojY9O0xyXk0JfDYhaFT2PHN53WW9piRfX6nLGz1cRtEhUKZZtl5Wc
R76x0unya5I9BBUSijoqa6M4Et0YIL4xwiMdJu8FqyKshekH+0g/1tF60ce0
euXgVojtscFt6to2becvRVRY2FrfPv4DeMHC0THRguDtfkNGckWxWTs75xxV
q2s9GnOYxHXtKM5nxdKu34etn4T7yhHzSJTAPc7huqMDrbmWW+oLgd9/He+/
xdm5pL6qe6QFfqT+3gNsl4R3r2nMN7sESshD/RxgOF4zhCAXvLNfNyVpQEzY
Odd/hHh4nRySDPEz+oqTIYsml+5Y3UtPyYUPgj1BfIb9kpabpl45HcO/n8tL
3AbDiuv9owlMaQYwEaXocqn5T09Ehw5Ddo1H1JMeutwimFN2xhfKRn/Ey1H1
RkDTm9llYBI0qY6w5Gq72CKngvxTfBJrgk8Z8/ctQdswGUjlbfw73FAghmAH
7aAz+/McxJLQKYomA2XIyHBFRBZ/sbzbow1UEWKE6mkrXH3vMuY0V3w2k4lJ
PV2F0eaiD3zJCkGqXJnuP97CnEFFwGyqrWW6MTL+IuUay3x7CnDK2gXhIWda
t4iB5WODNmznqalCD0nOv1+9CKv7shNAqC90N6E3llF7zp/FdZSO/J65uLXz
Kq95WM63k6NGrJW2A5a44cnjSLWkSYWhYJU8KSBvmxDE/VEiWRhiPCJdxcs4
A+giA/fR2k3sTA6LuZcYY7SJB791UEn87NIfZgVxyulvrvn2O++//tdnq3gE
v3ImxXugfh2zrzJIpSM15FQERrvy8zlf4sxRLFxi9tcGadQLCsx0u3w+ndES
QlWMLUaFwxY5Pm/YhsigKQSNlWj0gMG+5VFIappohw+YHaRtZBjrXYcEloiV
+R5XOGUMQEumZZk7DXvqksLETlBf7Tzjaq9ZThCh5WeS8uqux6WCwKkzM9L5
CN9W1Squ89rgy30ukdZIAO0uUNJ3KK3Frae4kRs9AkrWFrfTI2BReUo9drHP
SP2cbaHCyPddULJLRGyov6ENw/glnsWhA1CJGXJEG/EB9dUCw6INm/Pm/DqU
eZBXfdcFiY2yv6/ycN3YWpZORnl/6zpVN6yt+8q4wlj0M3+B0rRQVDf39L93
7ucuTVCV6JSSw6NTjxlxW49gcesDvIG8J1R8EGGntvHo/RZePPEkqx6jbTAi
vnQLS+JTObn2/xGskgiUdrqwK3i3sJzgZqEXQaq0tyzZLaj9Dj14/RkF3bMQ
gfOLlIHBiHFv/m+98NrRSMCsFiMqsY2SMzyteLH8zF5B2Hk0walTIp4+JvWa
NVc++JLDjWKsGN6zkqxmbhmTCNiFRiWpMDT18mH01o7Gxz9u7NJt7koUrgxs
Wn3N20phwmQZrdh5JutlA8vFFcI3ihiBn7r05zwRBoN35XrY3YmShqbLZ6kT
+AaZ0O0mAWKtZbZ0mIZu9Iu1VnNJbtzqU1yhPnJX8ACs/61QvTRrWPB/ocJ0
qoJSFami/0LgqTWHQimHRt4Uf1u2Vdd8bmOsqAzaJi4i1AU4dQGtVWMSyU3E
XoUcCKJWfwyKLB+53yZe8wFwnJl+5hALusQboDnxdI/QaDiWqGBHNKD1kx7j
f5mESXK9dHKG5fQTvi6NSvoGIL4qPeVDy/N7L3NhrhotXEfvzpT+vlqigVOC
+g25Y/e0660UtkvUP9T12almAXPHI6A5+E4S8UZtvgpPx1ZoPPCA9PNTeaM8
jY2KM4rGvd9lQDqK/iDU16DYK5WCc9IHMkNQQU5V1jZQL4qfvIHslSGaA6CQ
xI0wnTMzE6qvNxjoIYYWn1XVQ1T2cWe/Cxmq3HaKf0aADVQtAWef54zEorXU
HZFg4nVP39t9t6kjFJ/rEHzM0GHVe2tmxySFcWyW0Dp4O8MhEj2mpTef1yhL
9zc1/WbPGl+dVaO1dA6TCqOMUwonV1pweVzcNSzZDqFYwb5vJ2kiKx1x/Eyx
M70G9fRg9YC5nGnffZTvnyKbuDoFRWqswSF1yG/p71J1RKwdy2PLsF8rGFZ9
bh7XasuxQtufDFK+t6bjhUCrwBeqt/mpObuIZJtTiDkU3U0dEAx/nHeHrmVE
QeAljR1MG5Hv6rwXDkpaTcLmtkVdD8LBhtxt06eGsVWhQPs1fUrqJds6lpzO
pW0YvF0zT4VxSa4455DTays5DLP5C/frK3mCrJ/mv/zuFTFNxModxG6V12PQ
0c1Dd36clR44I0ID3fT6KKamS4zTMhkHdiLFSVyLLFnlBsvp52wSoLhjXWUh
jPlAUTSHUOq3iZgkq/bmvtcygc1GXI9XaaSgTAvBX0RYyE/4oU6RjTjebB4P
cqK8sY4yfTz0p8TwoXLfkZ1z79yJXUZVMFHAtAQxX4Tz+xNz1jVc3yDJmHJl
m04qy5sm0pzN/lwkhKSBCQ3jnR1k6/MwEX+ycZBKFnzolG8j+U6trX6pl/5Q
DaAPrwKqqLHEHHgQtZmZXHOmqhhVuG8hb+GK8MDEz/lfvUXxyaxNlfqNOgaG
HYzrd2zQEjUIbhp9UQFWb6pTLAz1vFOjulKj8srTQBLQgByPJjaY1XyzvnGQ
EBH5fKDRv237OoNZ572KNFxrVD2RfM5BHIjiSpVwWkEuQXTnTnUZPKVV3pIx
rMMuatdxqnwNZBTml9f2FXj6hfRHYdK6u9JS9KeFBEWJQNl7iKZ12WUQTp6T
ezxp5TxLwDkxjdTJIoC9DR9EZBT/0M7jh4vYQPauVrOys1GKwwDCJQetYPxc
uvlagSvzuaDw2B0Edv2ZK821UrlA+MB3zkiUjMr4iyKfTbJC4CucSWAwtCz/
MzinaYf8KJxHhPHw8nHn0p/cS032JT8obRwkS96KFK8ESqsHmNtOWORrHNFc
/QIoczmwiDukUxldLJJmh87JFjAscPo+1swUYSepWKZ6uBvf7EypDRNd47dP
/p6qzrp3INijXeeRQEA/BRKN4BbTJMkpvTTGi3hpG2gHeDIiC2fUYdfEvJX8
3iIdEX+wBBhsJcCEFbmT7uzjMHKJjMd3aazfDgYZTI3aVhJ+N6louk0M1mBb
F1jQNk+6RMwvATpSxtaHTIBOn7F5KtfojRY/+dTX/7wgv1WgBWAj0Mzjedks
aKLufQOPr5wMmTXprzN2y3WK2HU5Y4RI7TW7Stx68vWpJQtTkxJQ6UgHyeeK
XQ77mNf6wrN8PNJRWYAtOJsfeZYZPGm0KbKXL3P2aRx7q5scl4XRuRBjqt8w
D0lsDcenTo51NTb5jRHx1Yny5VXnPAWUTZa3yabDKt5LVXKYYUpPOwC7iNk3
KDDtMsI4SQveE7AJtGrEHlKhaX9T08ltOOKEfqSXbubvm7AU81apBUo1MmBV
P25MVtyR2qB3QVwjyv3+5jrw1S0AK0Jij95Ld7SwgVpz/wI0gi3bFn0+ULv1
3+ePvRuAtBsySIBoiq/yt1Hx0j7Ezxst/SE8y9w20SD3UOKpCF/upANqIAbg
tZd+Z+B3JvZxMrDvvgQkgCEYReNx7+EUUwexBI86ta3g+rDV7ye9Tnu4P0ER
VB2RbpFFvyOWEK264lDIFP3twq8o2BVaKqZfKBWOkG7bpjoqH1ftSVWuBdWb
dHsSFLsN7iEqFpW/iLRpVOdDgOh5+DWLDCN9FY9TGQX1XuoJXkJH6GXDn4dm
aFau4oCcnwyrArk+eb8TfjJEfr0vl0xz+Jh1xTGeu8kvl+zBjFj8sAokeZtK
tMoqoRBlm2cNEmRuZoNMSX/aU16x1ietkdpz0MHXCOl+8Dhm3Vf3WwU3JN3z
sTcuoDBOeT6MYHuvnTVK4WARTpGxaa8pTw6bPhuwtokMep3ZzrlC3xIEY37A
DlXoprG5cFDCK3JuRhS04734Z9AjrBODFvthVZZXZPZ5l3l7rJqfP5tFMLnz
NqSGreWI8LocdbNcN5eD3Bm3l6kFpYvusakEIidyrOoPE2TmJdIz4A8STIBt
Q7NuUf7BlvbPdKGPh5R5mPZBIRtrEIrlW8Yj6oKbZzXUDrCHaiRrDVvS2uG6
3kYl+R4lAkKqqF8LSTIg00+YDXZRg2P6UetJgdkbtWcE9DM7lmcHRh6LNwmL
1Fk73e0tiK4hgaZ5IjOnRIvkEYaSpANHNMCGEX0dXndwPrk9dWhxe1HEoNFR
MiyRiQDvrAqWW3mofIYfTC+FUJvXKSBHXBMLsZDU8KYIOjpGRSWsB34IF50v
XxSRKPdjKXvBLvd+RFFASrSzAneY1yFXhXFDWVxrAjs+Al+EOsHz9LGkDw2W
/WQq8RV4nqfaxbtviAzUzULVhoprlzfD0M/Hw4pdo9IkpsbsbzNu56SzakMr
T0xT7ts3fDOYFCA5dKTIeiPU5UhQubnftK6I9bHQfEpZNqTqePVAFaHI+Y16
cwYx0KQWEmDvEqah2Upyx/1TZIkRUGSkfPr1iqESrU4GBxdTy9ki/zPK1VAn
QI3zpc1Fq0u0VnRz1lJxCxU5dDbSgk/Yyb3cCoSSA19nEQ9r236K4ae9Ynl6
SnDDyJE66SyG7neP0reSbc2v6ukaXGFbxXZWR9rc07NPH1+0sJTWOd5Xzc46
j081Jgffv5ynPeol6rJ8az48AOTFNvZgSi6VMxxLmK6UuXLax48qlJAqMIBr
h60jeiBeScznDi9tpXszyIJy5PHNAOs2J6MDxod8ZqlsnsDGDeUpbuPdYuPe
Mwk7oPcvmRtAjgY5+Jeu04rAiOTfGKAIgTT2NQVz7JvBzTvc51O6VDwem6vD
hSh6MHmOHK5yGJj+aJVW7jKxep0HDMvpZFx/r0bY9ZjUcb2ZsgtqSqQfWZCH
+8pNeY3lzHEttp8GmnC7ZbhDb1whn2CIDnd5zmA/7sm3Cl/Q4z5BCpH2/zNp
SaZTnlXEVcJJ/7yESeUkhT+suLQVGRl1XhqAnGWe0BONl713/ySPYKNZIHS8
lLbWkIUYogF6lX4AybIb1XG/jX7eHb4lW83vnQ6R/EEohHPhwcNYU9cwFHT8
FLgdDqoqKKBuV5pHRUFPz+QwGufkvXpMmq0y6qPhVdy94WIvGCDktqgxPHtH
lRdRcQbDU5ShUsmtFwm4jKyfpOlI5Lyy4AM2OFpsgCcSpurrHz3ruJFi6CM6
jgjQ5JTZvpCChtfI0SEjAb492oxI/dAtRlEXsxHCJ4wIYuvqbgrxnzSy2rRk
UjtM/4vvADYbZSGYmSa2Bqu+dOCxnIR+7mzG/a7y5Za2DGUMduzzL1VFb0AK
R7uqgwNzjIyhsCRQP/JASjtFdy/bosUs3dFJIRVTCm2ZLOXsIAuAkcn84CBq
1mSdvvIIQzDv81j9oVyedd0QeUFI0nKpYbdlquODKmtFNj14F7XjKtuYvL/k
uEYjaD1YAyNDvSG1fYdiCOuLo2S8MPVnhQi3gpPz309xQd7Db5HBauteWcGl
Q8m+9+JWGzz808t/Hw+tAEv3kS7ctZ8TY1pUsDc0btcHMXeZ+nNkQMCLTUaa
AIgiFJqmUGhhA5N6Vw3k0rRM3W1KspXjMcVJjjl+7lMt5NsZCin/ivonrKX4
uM9KUzaTb3OlxgigK7hL/+bm8iOamDXeDX/nQ7rVkqCEaFDabbn2QnI45yG2
ELVESg/U23rr1KRESUotAJBMxpWiHpwphbzPKnsuUojTvJedRr9GP01v5E+1
u92T1qXPhGySQeULIICc0WDg+lZeS0bz1zwc+4/5O93Op0we3LlnIV9ENp6P
pBRCsXls+RxOv06oQXrBb/lOsus7KyN3Ji/fTz4gFke2bcscKfDOkB9Crz+J
nC85UZ2CAaASIDrF4Y8IDpa6TdvcLcQnUEV32WTJ2JrcpVUnAZtN44+GuFea
MMAa+iUvkPUw9k7SvTowC2DSDWcCfdXM7D1O6dmzHtWrCgv49jXgYv3+bbId
RtI8ya1FmwEEzSeM606cKL1/303lrCmAkyLGcIzxlgrOJMWHHEt2pC7O7vks
01IjWNpGyaE8/0bnFZK1VsjAhRVYY/4rTiUVSONrk3a9nA3FNwpVovURHVvV
lZfLpHqNuMvQ81RROMjBEkswq2NZmfz244H67txfFQCZLbnpjwN6qUHiCmTr
lHNubPX+rNkUxR4lFP5Lax/Hi3KrjOGwiKmD280/UULxanzI1WebjMF9Ufv0
nuFC1cfz4c53ZAwvbhD96g0qy26VsPQ9YwxhI0V9uZmYBy/ZUcQyvMmmkojn
B6FOPfbatvd3GUep+1TRSS6tbxkXQWrvrKgYsYhAIwpspoRL7LGhf1DlYLa/
pHAiJmLNqUa+ClzEE9aah4gvNBzaW70x9d7Lni6rBa2l9iNnBa2rs5yy6Psb
5keIM/94h8IuMnECFSd0HqUJWxhKgFMoO/vNWC8kLtHzaUfzXg/MF/FLpWGs
ycy1obhfWFr+b6HkJEKpIeOhASVFOkPVqW6nwi2naWOUapY6K4nfV5BKsr2u
K794s5rKY9tl/fMLg/HXnUKwlE69oHvkMzdW4Qt2ox0J6GDfvp4g4u65F2gy
svSZXZLHqbsYND5MO42rsBvViC3pvYqeJtQQAk3zUvG48hleeyC09e8PNB5U
q4rsxz6IKFnp5Zs97cnKTVzdaEX8VXEoErj+PEsfPG2dd4c2Ys0Rdgtllxrb
pXEiRSx/7zM15MLq0I9U8lnVkdrzDxaJd0oCeu0kykAKcWKoYakpDZ4Wqv7n
gHSfLwRJSrKhnkCjbNcf0gEdynbiPjiKz1eExSWDlb+IiChSrX1F7sgb0e6j
Mt6z7RX5CRP2f+tEaEkA3H3410FN7jmI/uz9JMsgpNdLqyMnmClbRQNnaRrC
KwpufFOT/5tWD7LJIQKR7PKK+I0xyVquDp9wpzyrPaxEXks0o7p+LwDbLYmy
Rdp9/wUa8EKFEKfx4oMqk/+eLbHU9e33KCyr+0tT89Bjy3Y0YaO6Wr9svwKC
e7g+BKeWaM8AIZ23djfZ4BndSu6fqLijpmVdmKKefsei7+kJv1gw+CQu7ruk
/WyZ4uq15j/xgjI4LkYQWujXKmeR42E7NFSoLB6HrYcUOxCtbLLPtIUIaEe7
s61469ZWTWZBaL7SUNRnCD3U0EQ0EDgzWPst7yTJa2yBWJJfAOHrfSLNxi3d
Kveq2reyDBPiivMohoEOgzirSs0aXfDClx08Y56KkpnmEIcNhPFIW4FJ+31f
PaAnyeQkWIskXJFb7QRAhAdtakkACJYaQaleXZgOzngNohJUpH5C7A9ZLNNE
6S495bRtPkpFvd3EEewsKsjd20NmWsoW+wXlP8anjPgkOebQIKpYlSwFiI01
1c3WuzamzUXxLQrZfZLxglDW4ae0weCou6gykmgTk3empaGGjhYHAGZC+v6n
Q1BYyCxrSJOQ6kXVHYlyKRxpc3/L26eOMF2cqw/EQMiHPali3kEJFpOn37is
ZPipRPtHamnqMB34F/fnAVps/sGQTxA/tLSPpCEkU18iKWd+X6mG0IFEVeBC
qeWM7fKqNcOznZnpLhGxEWTsAVGvcoS48gzYiZ34VTrwWJ62xGADtfnCrwn5
PeroDcdvfTHY72iCBX5ntB96Sb3fuKLmG7qNsDHyEtFmlbop6g6Rd40lFS+R
th6e8tqD01bZGUfHYtUiidKmgNzJAOcVyg1lvuc2z4kg4kAfiq17y1efRpyS
8nlAcS2QSCLaytjFObO/YqrhYUfahAatfVj6XVFzDQiEePzz6ClyNit5D2V1
mhQZhJi9teLXSHE0GFr5IDdJNyo71iwsIOzTlCiY8Fb6zkg4/pKBSheefwv8
5zQnZMEH/Rm+E0D57G+odLw5lcDVlPDPP6uZStMUoAuxF2UcNNlNDCNRbjsK
vE8nn5E0Lg/5ucg3XM0bDVvHPg+E/KhXRgy2Xn6pEa21qw3sVrYt7t0nTFL6
llRmQRi8UobQ3h3TPTABahoYKcq4gg65NkoCkVQtbvnDqwpmOQaffHvTmJcK
fvMGtno/FC/tUNXx6mD00Og4Aj9vyQ2Wttmn/i64ngv11ScrM7IZjwlpZ2Um
i7B3wFFZtBASwTydzuWSgj5YbXI6cnAbomd+xX++uin0u54J2W7aeNYiilgP
TsoDBOJfCa+2hEK0vrJUtFkXhmayhKV7QKg41MLE0Og+b8DYK+Ke9XaeMVhJ
oDtZ8XXTXfjzfAO313XTYi0epUxEmxENRLFCYyJuZQVVt5i/SXk5pjGUQXnu
Qrfl05iEwRiej4joikJA1Wx7EWypx/DZTm4wLQgGZaVst1Am6s1HoA9sCM3s
9HVaTBmtKzj/ARlOnU17IN86l0B8X6gVXi5n2U1jTsnUYRy+rKEJUjT4XVGz
ivOyDYdWVk1sv6+yyufK2VHZ+c67F7Mq+yQFHJgfqqEg+wGS50aDvJvY3xwc
ocA+DIZAYmOG4fU8zO30OEn/dx+mrO9Zq+UYhtlYSWhUn3S3+PulceSlbvR0
SkihgmPVDXJbypHtT6BCbpigBGOOqD8intUl8Fk1A7t06t+4ffDQ1Jfg84ZF
LGDoBAMcndqaTuBONVqHJyobkWDKmzlwrdVWxewH/K6t+blVqYF0fDQCZc/J
vwlMXIM9eVIPp3sxenlLF7e1tIMratPwB1qPn66GfPbjsm4oTaaGFOGBvBne
GtKzznxsllLMqx5Op5eZIGLcSQYfARR6kD7ZjQjfzISslepGKex4Haj+sdLV
k8c+3y+cfla1lSmKjRWyuJMPYS5nmaGwG8d1pjL8fOwZgi0Mu04FgSFrM22B
uB3P5t8OFthQG0/ltMmPi88YgH/nIhbuzXc64OiS40fjaWHmgEakI/6+FLcJ
vtjqWYV1RcUucFEkuP3hWIUGwtQVPHytNmdaw+tA2j6r5ORimZpX5bvDrZRx
huXmqrcYco1u3kCt+P3LzEikYOvuaHc9OYFDqgC5WbMN5e1pz0zJqcud8j9v
LC31bVhJfFWZtAig9jYzX/2sv2UHrjHQHEWU2mTphma0+F60LGK2dcZY3mG/
vU2/ZrO1wOvNw16D4kFLQBhaL06201WnoKTiSb1O1T92OSgQJQI0Tc1jM25f
31o4UY+599ny5OpWVbRZBNCyh1raBb/EM/0utJW3rBg7lwxOO2OlNuTVwv9Y
wMwj6idyexeecplYMtf01woKzoGyQtFEJeDjo21pYZYHPVKuj5Yth4UrWJxI
dHTRU5C2BKoIrp3aq59+4bDmP+8oPlw5O5bqKkSzoHBS/5c+v+KfE8IRnQ7r
2eBVTTociBPuh+uonJO8B63x1dAkL4J0dwATgPB3rgMIESwEyHlQWtsIYeAS
HIpfg8KbcAKTO6Glc40Cv7SOAZ2PvBfF3aC3AvzM2jSVh61zgSY4RaKcdX7j
F/ty+tCphbKkZsfd2Jl1xZpzBzH+LEAkMJ937DROe489MvQT9PWMmHkg3SLo
+d/gVQOck38uXiDbsaUSNypTQl7Sz/QnNP2jYRUr0FcCpVBO35VZul3qdN7e
/EYpRSgfOB20ihw/Z7qLQ2SNksla7h0J3AqUd1DJGfbaDbjr4DGOBaZgih/G
SoSGkI5wq18ZFa9PCkorwdr1iskMiin0rxheBnp8prTqM3BBcYWDLze7jTZA
hhQdpQij0y4pMxBKucPIm1NdeTHMH4DaPqkA1n59n6Ydha+HGtIwiV3vbYH0
aVOzOQSK+df2kRNs/FIUiEdHHaQbIoCf+ujkW/LUYkgsyA1mLv150GF97gfM
ShrckUI+GjyCWLbGatnwAyDLHpxEPiNyTCWkxV5YCOgT12GdwZGJo91KuwF9
uHMxxR39aaMiz3V77Yn4aRKcCFEeGGyPEkmtN41oq9RxERwhKlsTAqXDmEWP
qj0F4o0xU5R4H+iI2nsVLSqaMJGr3g/6H/Prw0V+O2DJih32buUGVQXc7WI4
47S2oI6xAvejjgx82fEHvvuJystsS+VgT1mztM4bkMZRNkQS0yWYBXs3Fq/H
O/FjHQQ761iJy+9EqrbJfwx28PjmuM+ww2j/bCKv6dax1JHKFJ+FgXoVVeZ/
qKUeK3NbJ6C5FXdRjd/8OmVuwom/iWDuPQILgu2bU8cr9dYSlZUyJrzbxJ+M
B1wPNqPQlWhqikLsO1fH4GDk26A4xQpBH2Eb6w6O2bTbHaxKAAXTnLCDVu3m
zn9N3Bvv0i+0BgfXjT+XvOSQ6dAfAXpJT8P643HHL+Xj+bWoXmUNtgfSgtI4
2aaDKVIIbOeEPOHhqEYILf1y4fsPqHK5WHcYr1/pFUIFvAQrtHv5L6Qo0I76
2uwMHj1hIalt31MKzeczJiucd57hg41zfxW9+CfU9ayj0Pq0+/lvokYc7WB9
GXaxmsZHQ47o2ZZLER7WIISaS4bF8KURj90H/MlUsJzYgDhSkNiovJL50WMA
oDAhWpFhn79h2zCQH5xoEmhgZ7UyHugCzwm9fGlkx6836S64WAoY6+kLl//7
d75fWvXLdJumc+EGaxby6TXvMhc/TblMOD/ypWmZbcfxfGDEnwy12t/sdupd
RUSDPktAN8HDXT6T8cF2CBEfBsNHsbZEZuNBGBf1W8NIkYl9XOVk7WAs/ryO
dpwaU+eM3fhQKrJjuHe7yOpL9H4wWzDrmiISkYfQcOn1SF7N/C30gDoBrKnL
esd23riu/ICoL3XX2gjjNPM/6ZleMr5yj8i3t+TUGTaVEinCNRmtAp75nuoJ
xiD0TBj1Nt7+UoWSPPkLGfQVf7vaKvhJxQaZSOlcIlbEK1D5ICQSGVEB3/c+
eCs7E7ggo1v7PINAAzyFj49yei0OCn0aNyww1en3/3WkeC2BGaMdrDh7qoco
uTNelKIcbUO6fWKAAXmDcTMxQ6uibdQ3TBfT4WBLpXMpGt9qBPkMDege0e1T
hllmhGgcpZaHGiYlUeJ6n30c81JoTTyy0xWcLlpwBRI3oLyxbx5I/BJ8670q
IWiucIs7SP+MDV/xyd0fa1UzslshY9h/hOZ1IFe3/0XWChLt3yso8ZUfIgQi
Ka9rBgxYllJHedihTrKl5ocu7+0nGq/2cCIw9I1WZCPBr7MieoMFyMu3fGaV
du7/2WLbMA4A7dVWBROFcQgAlEbCk1tSJS7UPEvSy5iCXkvE4/UWuyUQ6vmo
xXEtXV2eMsksiVVZJDzTQgVUw0vW4UrUxWlnunqmTlLQI5vY24Jhcr/VWF8T
YBU0vo46nPk34/TNCHtjKQoIcZK2T4pHE74yVCXmxtwq9dcoHm0CqeC6yXqk
q70/3pzRbleVOvRAUAtmu3X1Lwq/omg56thrbPLZxOQiocVonetgO7i/2b3v
45FrCw2/Vl3Q+2ECgGfmWZie/G2mG5ZRbBrkGWJQyQLdw+VXuBqiCG4DwbWd
au/ucLKOyqC4z8KtiAz76kuaTtOKdzMLAX7ZdYbTtffjli5qahegZ8RSAUjy
2ltOjf3HaceiPfkXnSiWQNIuyceJcr26sRnLRUwErEmUzwJcSa2wOoveYY0w
snJiF+wIBYcLv/38bti7KVXtfSlOnzQ5nvm7lYOR2Atpepq105gf5/vB6QTm
4h0IEZEOSfg6xUiynES1EQpBMc5qk/NDNHkV0+NJXqxl7zXnaTpQEoy7sIRa
GNW6OFIOcmGDp+KpN5ThkMDGMYtbyEqt4y7zdXrT7hLiQ+nNcgXajkBsICRM
ajQqW6eZJOL9cdxRaovPu7rorQmmaf8/nxlvWJ/RmHod6R1Xl5Sb5q7Q6L0v
4y4wsdrZu6+FWxOKzl5RKxOTH8BEOkpyafHOSu5J8fiNDr0KKB45LgOvF4LJ
2Lb3asd+HJ/jDAzSplUbcANU1/OfnEGvugjaeif2fq0cszeGp+KdxBYkGS+l
Hc2t+XNtcS359Rs8zdP3Vksafh50BSom5t5deubAmR1xm+/x7lABjytOJ/VL
UV3w0eoVV+WXL2NlD741qDE5CmSMHkoL5dLNyJXsKl7IHDKmtUr3JtqCXcaJ
2L6C1ohRbm8ajGtsIxRd3vDKy1tfl1If5EgUNn/gXEd2dzGzXL735F4yg5rp
VberdQ4z8vw2K/nmMXOkULwUcne9ewBu7Eu1T5AureUo600zJ2IOz7i6bFUq
kexSze/WFvfp2jtM1d568PUo40q4w0G1z4oM3MuuXdzbSkmw7b6kpWfMK6fQ
7qT+RP3SY+c/4De4wGYyVYs6YpS9J1eVICzdBIWXDwSIhM40gzouJ4GfZXlN
RPqKvyuUAjr15w0IzdlxsjYGVc7aVEFycCb21Sq2PsHEvLe2hWJSS4gW9JQp
E+HOZ+TGUzz16qGtVE68S8dz0YORbd/XDDG7ETaOlK0h/kejGNmjeBxToLUf
fm1fS2brTZNNLJlusYBnsphWodCuUqNGzKa+e9JFMhCBZ/LY+CgmLAB7wsLX
9vLzuKF3WGhB9FbUBM7uOXxEhRmPSX8Kkf1lOW1KaT94r5inNUiSX50F8rBl
8aduX0WWQyu4InJ3tuAmbWXhXknYKM/JgjAls54UdhSns3C3PUI/AnlELN9k
2Hgvxwt5D3tcghiYSqT0nfbc+HJ3VMckRmNvOBYHnEUalkx9r8A2FANdU1N8
MNbgZ0tCVtZInJsytV1+sjoY5DwGMDjyTLs2xg8+Os8gae/QLR8FIzy6yIU9
E9YlRqaAQtH7d/qP6GFCevhwuDjmc48+usi6THyoyrZkifKAP8WqzVBEGEz7
+bWfNSDciEKmGnFMRcR3h3ycz6VHdrM8hwJEA5bVGnkT6xTLyRdHzR5L7hcj
XCXHBR05o1VORZg+v3qJK7byeQr08Hi1B78rMiSd85RGV4N2uaZvSEDEG/7r
SQTdHkbu+LKsI08bbbVAknt7T51odD7BDOIadESr4xu/6qTzHfikA7rB5OV/
k/wSJNcl5NXz+NIViZbMuQJekpTmNn/hLlTnQxu5JHRarQvn9cYcNrCv1d1V
fP4649JwtI/HdXthQv3kF9fiCjH1Ex3EYPFcWefw6hrHKjCfn9nO7PXmRXIf
/Re22T4iDPcaamS8JWS9M/oFYeLNj9ksl+K0SfXt8ho+Tnj7fNS3i+FQmWK9
w3MQxeIDhEkqGZzceOqKrl5as4E/f4+BayxsbLgG6e1ueCMKfaSOdONI6Zsd
YoRRC9tr+3g+JLihmKDBjWpxHX/QhrqLlGIQGkxDofegFLs9NLoIUEUnwK7e
FKcB1ec0Sb7zrhycp6kfPkvYK9hIFGIbNpTJJO8uoEX72R8SdRBqo2QLsG7z
YJhINaiuyZWsjh3jWczm2Z0RWp92FCag+QYeqs2f0ANVRQIKLuKGMiCSYR1m
qAleQiBlocRsPij8Bq4YzxAEiHmT/UODRiW9TH3/Glbur14aV45we5c1bzJ7
eRb/+iQ8X4oquqO1+xIJYcB7TmHcIIuszBI0kN/fjPlYTWKJTwOnWGoVIl1j
vjgaIlg5l0W3paDM77+hHvLQCXxcnX7+41iPX445zqiiFJM698wNehgNy4g4
iaEO4GezKW/JoNpjmB3WpMl1xAB6g/pTH5CN31g/jg3+roF9ocI+vJVta6tW
y0cUQwjhenJNZvxqsF8UGrFZPVpY8IflNdA0rqNKl9tiWgR61e8kMZI5UQXv
Fn/zdJxYCokSyisjkBesEEHy4Pwo5RlpV7/f2jRrCocfHvCMoQtPdaEVdRFD
ZTJKfbxvB9G6ei9aSyVqUQGypZUJDXLx30bQfLuxgOtqC03xFbDhf9DefFdo
/ixaXubnlyCDqzqm4oLNsJ9wZSYTAtlfAByi/OsZ219lRKJNnK2PXszAGqbP
NUz1EuVmGWA7oS41VsMIZiWbtEOxtB6ZQDZPIy6WOqBRqmGtL8mDqsVzuxi6
lf5UfI4dVrtAzfkm1mwKjwmVLe5AiVwjR0F7hwWxV1C/cCOsvD4urN37wXur
yj181WSm9CRT5fMYy8o4DD/znDG30DzcBhW6veXSvuO8JBinmIPgULX8HtFc
oAAshWgvbA1lbnDew6UhJEUx6PJvQG6VrZ/ai9JLLiCdn3Bv0ReRtJkb/Xa/
mfDNGoKS7MXJSYW4LQ5QHkJ2BvwYt6B/pR3vCTuvYYeRJVTic7AteYXivblw
TlBBS5PYWLCD75LWFUQ2Z0HOVT+enxmw3c9zWd+mRdeWzs10jF6vO9LzSgr4
v16AdVFr7SXYirTmAIPdTTA6/v19oMVFshGXn1mUAlSNRP7PwPjtSVwnFOfH
kwdSHsITpRBCV6AkixA6iNA5EXbUMF4WI60UF9L1Y0YFSPqvGT3Za4ZU6/xS
I/UdSDlLAdGO9+KKIqz36pgbOAhpO0vKmwNue6itlPOTi+jTazdHQpUzKPx/
YXz5XpfC6CS8GXGiAp23d4PXoIKKzab69/JdYtRIR/TJ8mb3ElE++EriXyjp
bJ8jR68hQIkf+C3I15M5Xq0zDzJ0sZ3KqGKXL60gfkpWaMtZq3PqDUebJhvo
T8Jn1aabDMf7t1wdoN6eHqwahjWMzV6HBL/8GGmYQ+08jk3iXOdMKwOYfkyj
yu0/WNJFMbA2Lymb/HmTyfB5fFfOD8fj9WZf/xiXaE6ug41KOg1KbnwXBXty
T5TBmXniV2W553E6YCBXCSwwJMhHjfCTbiM40Pw8fzmweMU83iAztEre19Gh
zmN8n2HQqQUeJSCyXGA697np3tlNWmO6gSWlJeMlh2XeZCvmXutJf5t0uEZZ
g6kFm+QrHybUd5OUv3btK5Dr+S3v1eT2FAajDIu7UVR6Nu4f7OtqLIlavTv8
4QpsAQbw3dnYvrXF4hIij0Cm2eWy3KLkEooXt6Q+7eEGK8bvbLmY4+qZ48X7
8eq6LBDaKTzO5Jlkkwj6TLFwjqnU+3uoI20IpRJ26OqJsWarDn1O31Bl15+0
1jLSs/OzqKz/78ccdwSlDHhyx3cQkpXyCvnDyTEzgZzkrxQNghGITDRqY1KU
/M+WdKffITnbjMCGX+xa+SrRgc7yWhImBioUQAM8X2Oxasu++AHEJJdzRoow
2opaluSHQ0gjGr9nL8zxzbNCW/y0UV/RvjHIlptduphob931y/dRTK7GP35H
6zqEhlhidkYw2gclkSAlJwnW/5AOZhrMppxMwRkkAzO96T0894KBrVaxI55o
K3U7w1m5Jr/3JZc5qq5AY+Et5ESwn0z9Dd960juEmE042GkKIp0sT3hh7y47
7HJPi+6KZDZm+GcE6dBznPtfVfsAHci+g/yXpK/KcznAJL4xFNvFFqv6ybi0
1swCCshe1vTOXynLf7VN2qOjuzWBjiwAMmnzeJSQqjReCDSogK65byd/hnCj
bMmBPOKrdaWP8/EjnqVVybAy9fUnc3THssImkfMgjiBKq/UiouuR1WpRzYxX
eaxDSLaBohSzKOLkLDFxvV+N49cPHfpNK5kodzI3Iwbpt6gOwP4zckd0pK/r
tcDdoZc/EHa5uHp4tIoqKH4YmQlToqEO+XjENlgZHI1B/fVYW15JKJXY1PY1
Rtg/6cxOHhRlgysWojq0DtaGjhOdkJjp4WqFxhlu/nBXJtz07nR7ZL1mPldp
36eLuC337a+HdPktmy1nr/P1mpY/YTW2ejvdkN9qofbxaoxnYLhPaptHL44d
JVWXKTsa/PXwUi1CKllF4tiC0hHlpM7UaZTF0hHof504rdr10qtXcyrz3m8I
V2RHfELGN43i0Aqs8bMtzLIAgGyyC2FbQ+gX7JLe3GsEYbkvRIu0gi75I0GR
CjEwV5SyT5vQQ/oI1P2CYPBxNypujwyeX1BiHBjqtR7F6bdWmWHcLv4gE9zH
Jm+XqdscHGzI5/+43me+UKie1ThWTap4G1pp2s9JmSHI60doqdn1bT748WTv
NS1OvvNyg9GpdY5SUwiBRvdoIRCMhudaWWQMDv0Ne/BAzmtSoL9slx6hjPsX
lTBkejtrCGbAtt5AbBGZHpk7CISRAzDjhc8BSvbcwncnpnl4VyLel91yEOFO
pVZ9wZMRWjj95QdA02HBZL1dGTjtchLt5i99CnqD/+EoQXaa2qvqeeOKA9/Y
qt16BR46A9Td/k9NmJ8vWhvotNBtZ44o7RVJ9mwcASpNxn9bIV7m22S7ALPG
2IBOvM4/U2boy2Q9/xLj+gR5pKay3Q6C3bhXMEwEag7vW7dLYLBDSPs3VI7H
mtZ+kkF9mGWJzFego/1Ila4mzaijMzCPytxjXwU9749Ppvt+8iQ6+TOJSGgI
PdP4g0sljfilXZ4SDJrOk5PclJ3vq2aHLI40ce+7aVUCSX3GOcPtcEmbPv1y
pxHgZ8GdiUW1coKfa8Go7mP0pHi8Zi7T5uT1LyM0qMb5kWQLu5Ei98JV5BPG
MbBnluDCurGjmamr+Fpnxoe3KfQVBsLIj/A+qQ4UiTgS9Z6rfEYdFyuQlbJb
ig+c24MRpyVgvviwUGlAI4f8J9wnn107dIVKG9xGWvQ5j7CllJ4idQbVEdYS
25EDCMYcmbCD9m7Mny3LKifpIUUQ5YJ/Y9eIfTWwO0LOUFF63qcWXYTHTaPp
7/F1ZHCJI6hltknjniiOlsJcXlxEUmX9B5luX7JAD2LpTWltFQUfX/kyr5ZR
qNx2zsDcq9vv3zLSpIoZCeR50PgaWoEYxZcy+V9b8tNcZiZZPGjB0aFgVLoA
xz/ByrP0SWf/e4St6k8rfFM1ETrZML1C9DnLNL/Wr/7wcdhy5kNDtjW46TD7
dG0Q0H9Yg517QrbLIvqQ3SfPAUzx8EJpp+xxs2lWGuXLkOO13kZ1LCCowa4o
zjz0XYxSwEwCNQbsCLrlc7uqORYqJ88Y4MzLbpwNc1FJp2yBUvLteiJ2yiqO
iKaECX9CMQMm4ERadHt+skDzKuIkgypCgMQrkznTIdEF2JqKaW/Bpnh+NNiA
pctqAVFZgCJ46RpyQCqcl3TOSC1ngLUp2RtPCvRhUjNGyih+Jzo4itRuC38B
Adhue53sS/VU6rt8NE6qAW+3YrIgFH/PmiFYyUdYoPN05wfjO1TDotkj+T5A
bTORG4vmRdmlvoFKfodqmbONVMe36fVYDKg0K/BnGvoIAGRIJeQ5gJwNAuYX
rEQmdnEnkCbTTBqvYBhsKpaoMHn3AzXVPqe/RFEE9PfPciL2t66rIVJ/LlAI
VvXde82+tG9KcZMwb085r3vIaExVG8WP7WYojDxBezO+HDPy3oEGUEihgac+
gMnh0tBi8yD0gt0bDOVIRxzcJXvrQ8VnJYdwrK0vZha8dWPEwlX+rJmTEGl+
4dpl49n3Z77xJhzTfWxOQ9CdNox5dSAHs1X3XAtcBax4YNi4A5piBNBEqwo+
RihwgC74S9szc01ztdj1vGB0k4gRYBM2FNskL3SPuKotPgMVNOPskHuB9oeV
CPZaTlnnjhCpOdNyijtMocj5AACm1z+gn01/JUom848NRAx8V0OhnNLghVr7
W2sQJ5ju9HtYT0FJKiE322WoPniacVYG7awi4cTCdWjbz6iEKccr/PiFxFkD
nybu6UxlmuDuachWlbLQI4XF9qw0oumcSuJCNZ8C8uOYCMndlTe72dKA9FbZ
BvOVT2PoxsZjDQ7cJRRlByVj27zzKtGsAAOG1lgZ5y7YXyNQSRZkoR2+mIf+
P7QM69/b+TkdxuET0Ficfvev/AKwnpkWy+keOlRLw7KFeiHE+vjBph/lW8wn
83y514xI1SnB0Pl3AB62/RQhbQYbsXOYwaiM+/dmO48oPkv6tvXP8PVNsvhP
wx9RynIK8ZMW8sUIjGzt7zJJFmLpDfHcXjUkkLk7E268/QXp4qY6mfL+BK6g
eLGK+I0lABdzYENF27PssHXU6ZV6geTx90KXh82euiVkjL33HxjYm5RAWdNw
i74I1EQcJK62tmWmtDtmZf+/2aoh++DuaY72DBDVgv1lByTw5rP38J+0PSSx
Ner6WgLFKrv0ObXgoytw2hlNJc9LRTpfWXoTTf7nX57EdiYk5FRP3c/jAcVR
+HjGIqZZPoZTvTT8isDKzRjRN74o3Zt02yUfrrJnHkHo8cIl5QayL5KZpO5/
UxiVyCSOf7tHZnjlgmJBqZOE0yiAr0yOF2ZlzeFeWebRs591EA9xYNBwBWT+
No5/99ybEeOyOpzGui4k4INJwPWHA1eWzGeP3i6bQ3vhhmRF2xI23iKOE1DX
RGm62WhUAkNkhT+ZG+HsahKYE/QCkbBowYUc6kVSPIAIGbQ8GIV8QrWx+tPF
DEknj10STeAMkpxvK5nDj0w12f4yV3SgaUDOzjp1/c0H6sNnfIm31XsHI3N4
ct6ofmpZZjJvfuFhAtBG/20cS1Qq8V2CNti89eiGh7ObzF+LpMIy1drS7xFC
WTguYeNbD0K1iOXxEua2t7qsS6AXPh3SkT60Tfj9+FfW3FtvEvQslAuRcsZv
Fo30ereqrIJi/oy0DQ/U+dp6qmxfzKOlBQyGQRR+0DZsfDFjwKbfVHEq3mHb
4PTU/X88P7hlkoAupC2pwL75X5qvJ3W0LsOLPiExcjsCPsuBAuoRVfYcaVTF
iGCQtrkizDvUwrCSh84/5KkHwDDIyZF4GT52NHFDm4o+qcyjhtujJuPb5Uaz
OQJN7F9HPiks7bZFBawgpHWeunFkk7GOqestdVn0URxkCKdOiU6P9kbsB+QF
X8330Fyj4eN/RIkEjV0kva48MrMHw+fsN1ohnGnm3wMnWEM9dJKHhE0qZmZA
iao91yRY1IMF3mrQZZGu/BhHsX2SuFxLpIsW6x1AKUelIpmiJNO/pMPZLAu4
yZdLAJeERcLJ0PQIxRzN5rVPgWRIRWjgXHrJIxTAnJM5I4HWcSdzR0yVubAv
DE+HbHN9ybxsWgsaVvynhXEX7fJharnVdUe+1h32S1jjzt+fqFGhZY25R9Nr
gY50h9dSSnYy/XKF1g5UlPpl1pgRkKW2RePyI7/9u4Y/2pJRMKozsm32xkN1
U8obidqsXEZazXmbO65eqyJNzjXJj7+By4LorXNTm/Y9K4BsfwuszC3anIO5
jd4gmryJRhlPG3pXh+eAurHrUaYGFU73NO6CBmCr4pQj32OvfAQfSg8PXf+l
XKMAly8yMDs41QkxBTFtc9sr/lgDPLM7VEqeNd1DK7CUk2I2wc5sGGDVICkp
pjvQX105QcYMxD+XbFGhrVw5dTTNRSR7ik8oYvaq3qh+Rj/JfmZZ5wQuh23a
+5hZJ+sYr47DmO80W2LF3WOVve1pmOSLm6qtbo2wDLotskzDJRdE/RZ9xBGR
byY3J4oSl4054YSgxJNGqbahAYiqSMwk4tQCdxS8R48dZz8fI6TCi3/GrL4z
29m1xxXwM2AXZqiW5kbw206WOZKSFK8+UUW7LVGKPmXDcgrMjZRr9EJ208YE
LNNUefcYFOXIl5TFe8A+OVgWjXYF92gQxVRg1ApEuPAcAW9yC1lqen5wsRL1
rDwyH9ifgeFzJGlidUhJ5L86EPBoD0z37FgO0RAtKbAQImPHm95pCkJQ3eYk
U+p+vLl5kPKIkTozx6tObOYTkJZkXUiJyHXyQJym/s1mImbzY6oPYaMNHtgO
gmsqm2Okln/aBrfZzYM3vqkp6QJjCrS9GJLQdTqI3GllwqDWoWfyI0uMgPZg
eI9dmQfSnIp7UG0S+6TneBY9TI+18Vq1F5vgCfmgfJKJPvpYVDgpcq+sa5XZ
Zyj6RYY24Hy2oRFezI81HqoFx5VprDG9pViOcq1mciaDF5YM0Vl3FGevXi58
qeuTU8PlqKnMrcPtgyrYQ0NB6PVq70hDxz4fh4iA0I0IEF14ZvlIF/rex3vB
+oGJF5gBGTKFLTzJzyeYsQqNPFqI7Q9eQbzZlW775hApTMi74KYmNjlpNAdH
TiRA3PQu4fLIsl0YDPOGkv4tSs7ZeTLGX1qKffoYsWCcM3RbBeudOGK3qasj
Slv2UTp/S60iDOTM4EfhZiDI1ebqoxtrnEcJfzHsSxsr13SXEc5zJA6bbEDx
9L9aIqjuRyvDgv5rtV2TTkJ4ZDChDWqriVgJtAMez4HSZqbGIl6oEsCNAF2W
CHQuHWs+WG2aNPCmYWAs6j7JgAzGYmT18raACPWPqSeVvN2duzDasEabSr+P
4Saz/LONeA4Q8WNl7oplK/HIAIeMO9K/fmQotNn3YWq++XvODks6WRj64rZ8
sDmnMxPI3tz4aH++Lv9HoOWXAgFWUQhYxa5Ow8Va/ka06zcce5ot/Eb11yDd
6zqA5gu5zW1pAv2AaBvP9783blQeHydgiAKzAH4XCdaCuXzdZ0o/1vwHHQX7
GhlpHNL2hmcqhOWXqTW4HjTLJPEG8Z72L+mL7V9mbvzfXN7FSjwAwirOaOWu
YGClmiZDoYbt2CmrVU8BaTw5Me51Ixk32SBeeVpLDwFVYwh7Wuu9Ae1nmebf
kYLEejX9+51B/MK35pwHxFCobDsxZybK6RKsAIwTa7EE1+iY9erco4t6UBSb
dBoZU59IXHedO9jzxo70KvJsQSsZYcdYzIhMCMhX4oJaZ1dsZrnGaXxUxBeV
FLWJ3PG+z7lTxwnusKsTG1tNscQmiTD7vD3Nlrsn7FOjeE8v3sZaYWbuHrx/
Q1XRzkYJPK0HHl1SFiCIsbwKRWnqNNULZl+henKEFD6kaglPTvDXCgNoxa5g
t0COrRTJzU+gDjRrWjyvGMLN50OG3B6o6qQTw2vzbjqV/yxjj/vZBRpLNHgj
oGsAZP364HBbQkA1XOfKaPf/egITuh2dBhJVA2t0UBqFg3r8pL8dQExOOqjY
r4jOw+IXtdKLQcZ3ze4IbMzaLnGVaKGyhOFIiCvXyDtio19sQc2W7wRN76Od
ozniKVtD0e8v+LpPah6p4MXt646cMvpIR+7d6lNXxNclDdThrZZgJyj1fxHe
yvkdhdw+s5L6txcM2oU5xb5DQlqzDt5wAPoiDfdyNiOYM1Ltt75ajjBEqMH+
ew6Oe0lauR1+aCHYHfvOK010MfiBpE1UOV8qlPNJ6hmqwZqJ2hpL/zxXQYdH
YfPe+NwNo9ywbNUR/A901iv/18Ntp5DdHkF6ZHlQvSD1+dflrMj5fPmGJURJ
fRmSXqAuVWW8UGvWmmLmkdgLovVFD4ScH16tudXM/kGBdgOWG5TL4hckJYsF
gRMcCNHXmVBIO7B9lBk1G1VuiIMSheA6SRmPBVUscErH7C0MY2NwbSVDfH3g
jgS+NDVcxnUs68oq1bsSCeDsLe3ZaMnhiNdx850baTTvc3JC2T0yNGjuuY8j
1nXF0cVOTuXZHrBa0l+4zYS5fID+TbyvEHmlRYZvQF4kP39/3JjFfcOTobJA
gAtkGCyoan7tWFAjV9c4l7QqLGvfrcZEG0KkhMDVBKF4EW+RTYSk9GjjIsfm
8I5myrf78mLzHL/KPt5QXPto4TUOQ14CsrAAx7vWal5kulccI1AHzTXo3Luy
wrPbEzhd+nLpbyWKDus5c44W4LungkuijJcbFElokAebTuzBWpC+1ELBNbGd
I2KPmvgJV6dp+x9iI9JouBUFqdKbrv9afZK+eO2yl0uydEddgc3OG//yaqKn
8uEJq2dDy+SarBA7QYqPHRe52GlgTTR5f8Pdl8Ym4cSTXBudmDs3kfChWit7
PRXNZ5xj6rfJ6yF35D13fovY7rRzv5RF35az0gXMYFCqbJ9XdSUNGEDB8fiT
sjlvejJVw2Z/Bj8C2rRRGgEhrd2u5UvmAKvVvHo7ZrK1L1okz/0Wwpr1hUPW
koNonXlF070yk4AHKIMSnSvAd0QInN9g0T4gOcEUdgKTbHqVdE+uHnVxw43/
fA11CxN8rwjv3fcG4l7wMC0Tvn7aNMq5uqkb7aPao2cal/DI5cY3dmd/la6s
34WBHGMsL86XKbrmfwzDsvUgSIZ0mTt9k2pkRyUV5APRb7AyMYgKzJP/C/oe
sDpW8npxbkOvNL9kvGqT240UP1mhz/C/yXAksrgW3ejieV6yAVZuuMO+sbx2
/z3m0/ES9tsbxL3n9YejE5vWmxQA5j+ZzwGFhzp0NHAecb5rgMB5cJtzegOX
sW9ekegEoVXs0fwBadZA3WCvnvozwWQxnjLd4YFb3cTPS9VY81Ye7NXBa9gY
HkNxmXRsXsWbR3zXkPn5y4hOh8P0xBTOhO2oogJahTznrbDsAXLXBFj7ZvrE
HSs7ZBEVRDc+aSk/iaVZl6rTMSli+wx4fOA6H5/CvaSMjEAXjWnmULSKvr2r
Hvyp98FhbS9+KMIjt9dVmnsqSX1kCWxDcIZ7D1vBpJDGu/Ks88fVB83OBmmw
Ds5x0CCzolusxBV2oX0T/aNbNXdvFncL/LZR7BsKVjlOoXjxCdJ0nkS806Yx
ZyU5Vijj8LRohC/rWrNZdI7ZzLjMtvXX4E//z6XwyFYR/jBRZQEsltkNBvql
woAsPGq51GoKNq3l9c5UEMiI2CqCF9Fr4Ce3giF93MTpXnPVUoOgtkrN4XBk
qlqJhDGi3s04msJWtQwQwJ2V3RWgLZcnzz7NWvosVdQYmSt6LUEXVKJHtXao
yHdwz0D5AiSamhNAdQ7U4JQnApR1mMbgceTfns7ZAIcKfhRbuQVYYQV6e90b
ejbRxKbKfxboZjciT7vtbc6Fyo3fSXQfGMwFqpvDNWrZq3vKTSyeB/FzuFJo
K74F8W1Lvi8DHDwtruQLrNugRTbPKOffzzL4tlSg30xDSueEsfp480hjzlDm
+sT1X7mKx38Hkctd0kMJ3Zgbce724nCnxSZ3OJqZEFI2jqk7bwgM8qlkd53D
C9ETPNW1ZFb/HW8tS1e6ngSvUILAbsJhixGE8ChNfriE12eoD17x4kud128S
oLTmmw18gCssI85dpxZiaiRCEboELNjqCPRBQzezx2zMVuMdPe/B93FcknES
bNRYKZ3/eAtfBUVVxWkVWA/02tL7LTycvjka75qfDo/OgM8MIqk6WMUi6q9z
c3wfl3ZvbzIfoc/Adm6rMiZLM3pnLAt/951q51/sL5uCf/XCxyq9Pq7j6AON
naU1/jr+tCHO83yGYFU/7LSIEA3vFF9bNcz31pkmcnFCJU+Ccs3ikI1oBZsi
iX/u+l4CKf4Idacfrs9+cnJYw6CUonTd65Ulz1+VOrPhi0Qg7rZv8CdDcHu1
5PlrNqFvcrP0oMGm34/nAaUXKTlfuXXqTIB5zR+5lsQUoXA+x3x3N3cy/MQL
8ybUsY9N2HtMnM7KNkpuxV+i5X6sndqTNNuFUB6AjzXES1cP6MkA6xnW3y4f
WARUnuXWGR+2di9xG9h4y/GwZle1s4P6rUzpH6wuUzRfzh71DRQ7+CrBMKpa
oXszrQs8CJGEhAeBtxkwvpsQWHGMWMctgeaAzpArzReGsnvz6/un/znMxY/Y
855uGkaOsT/T3KabewRQX5b2o++pgr5zgrIcLJkzwruPvOaObv7n088MCeUm
pwX2h2z8W3vw00bXErKXsn2qWJtM4WJDJm7hHwrpJqisxFTAvu3Ns7xIFmir
X6qSlgtTPzuH86TGrqF44dEaleIDxI4L6FVmcVEEQXnM1syH8g0eSZ9f1J59
NIiV6IFDfiFdVBw2py2OZY1kH4fNwT1GKPYUcq92K6Ak7Ho3STPvc4zKFhUY
CLsl8kFDpjf5Dygm/083CuCp6y1w9AP58KbsnABcilYQQyR5YSZtgI5tm18M
VezEBFiOfJ1ap6YxfNDPNPK41Apu8esBoln1QSX7Asredw/S7ktKW48j65WY
z5bEMuyLYvr297LfY/tPcWAlxmltye1hc+0iizZ47ksdldRngv4xm/gM99/b
xrbPzmHwGDJHKvcJ0KttMqA4VGox0e+GHiwpkHzhZOPp1K288GpYT3c11Wyo
7xNtueJ7sUj9UKyBvjsUeE1YB91oMFezf/yjzh/lfL0h4J6JFEoZQFdP5UYi
rk6iDoyEdCSo+8Ao99ndn1Y69og+d5zNeosF+wwXPN9ODZtH2m331As5/3qc
HURmeXIFlVNkM28Gy10+z5f6Nd/Z4vvy2cWDnmOYEmUBnYUZ0WY52bLoIT6y
r3C61vv2aZVNpWHyFlEScY/UVxS354ES9Hp+nSu48lczfqLJJ3gI9SnVohgj
1SMiAtLHXKflSOPMJ6OYg9EBjveCtchcVruWukT139ECpVhj+BeLWuhdExGq
c6O0HlChcQvozbxprxfpjqzwosp6uYQEKIOYbmLPyYWMey0kXnq165vicaWr
AA2vIJ4CHAyNj98alvi8HmExtR0LejdVFFcBSLQE05aUUnJKQszR2f/hm81n
ovaRuebDWAG9V3lavQ12QF0k+sm0lK5Qa8cjrAtI6h64D8O4/Vih/lISJlNZ
hE/YKFmTobaKIzHx7AdI0LjKd+wompxP2C+tcvf2gp1STnfEpEQOfUVItKBM
QkpI35kCpJeqqI0+oCYj51VJGw4wdhpaFnD3+jKY19NUwfjoaS6KP29B5r8M
rXulsblaF6AyXnyqXs5GdqqZfX4lMEhWkxVazDOuGMktbRoPnHaxrxTPINux
nOZCX0+MDrfrDlYpp8irYXzbH/81eu0sVIUPRCPe5rWmZF+RLE05K2a+tfoX
Gin62p/Yne3E7PudDrMg1f0oDy2Q4VhH9s3DF6ph1ldiKJv4qa3bsc8bzmAr
ijNr3PADx5G4cFRpgMZNW6Yjcuh3SFE+8rlPTkBNmrh8zSMg9mjd+Z9DzckJ
Oz1YDZDuMCq0zz6OwZyBmIbIiJPoSfjyJGNW8WyHM2VivhON0otBjOReC0Uj
4Qbnyd/iLxU8rHJl71x35AB/F2lnphFC7xm+fjBnK8HY8tmkDP3mqQxHHTpb
VPjUqrE/u4h+RwAhuk2QbVYXmVb6Mr64T84TFQT6EQ5L5aQQ4ZQw/mtMVgMZ
qkcyoooZ9kWZb8QkKz2ZaK6sX8lhVbJ9pMOI1iNv/+Nu4HrCwogrJ7op21f4
EpS63w+nN65ezCjAgFLuqNXIxSgfg39dLbmESlj5De4Bjv3OM3OgS7Un0YpV
SWtuMcVv0aYXNbl6PoRffCunA6mhhWAicJt6415jyKqxlxQpoV69lmzmBeMQ
lMx4ufZSgnOnIRdrdFrcD7natVZaG84TCZujB+YB1NPn8WLFM8iaglHUvUjn
9UCgsrPJL3IrYswvb0eMcffR8Sv59QE5lSlfC4cOD0ZiYSSpvbzp3Edj9P5u
lYrpFWpaqB8b4U5f+JdCBSx+qAv3sdHq3aIfhNX1IzfnFOdUEIVwGEb089om
Vn3DlGUCAEqTO+BHvhbEpxBL6Y4UhNEQIJWW/DLxTyB9RfyedniqAhmOvFL5
Cr37hVGiZwe+OZoKsg/TupTaBN33uJj7UohNZsTLB53xYWrMIbeaSWI2xotd
SA39May56oFiExwFd8BfLxBonMQGvLd6kfQQ1LgwDIV69ZL0SiPdtiZljw1v
gJJ/6OYFzC31qnJiB7crgG/7fU/flf9R4KlgnhTlJEWXmxZeIFisuzKBC9Jb
1wAQJujJJQVazWowp6+n/tETXDEsQ8QCiGnKSVKnzsHNXTU0mEb9clbRVqKk
h2zt7iyMJjJKXBcK08njVWuawiSyYpiTMqAzyQdxDbmEzKrhwASq1ysp7BBv
Fnw4H290ye1lbQLBfqa1DPEC75BfZ/XABjmH+fEacHrgUiZ7iy/chnoyhJQD
y4ldHjxla9e0ZK7wE7m6XXsRht0fQn+IcBKk/qrdpyH0XTYqaNqxnyIwMOAR
6QZ5a7N+PGkEG33MMfe/WF6V9KrTavZEqALQpC+4IVGSKxSfh31ak4ix8auZ
cfyBV4NnNYlUjBB5eGVFvs0GjC0ClzvL5I/oyBFdL7xBdr3jA2kUdU8SYHxq
cME+1hYf94R21ZN4bGf0zt9k+0CJoZ8pfTWZAmIjKPEbO6vS+E3QwHyyyYgF
fGh3YHjAwUiNwn2jpUkow5IAamt5mQl3QbqkcYEN7DAaftdSWbBqZNA5dijm
lK1DHG8rP0ht8H6S4Jt3aKx0c8RO3EivNbjUJVCzkZSsib+nt/TMrPsb3E5B
0zdx1kEOK0vZ5nDxAk3JIGBbO4PikZekWn+gtVrr9WZT0BId71x5Zclq7kFz
PKvmsppcaD+hUck9LiIR2gpehPf1VFsKc9zMn/Bta9lBlqVJDlHyARAO1C6L
a7DC2Z/n/1v0YztBomkJF3bfTaobM2Q0EFLti0W6oUyCszi2C1Y8a2zhA2Og
z6qiyTkwSsIFxgLLXspQFyjTTTlrz2jnCpLwmfcGRlqaDBjVOdS/VUMSSv3R
YPfLn8hV0nltGH0Sbgj3Z50YM0M7MyKwbqxW0fR+p08gbs7KhsFn5Hr5gn6z
k2I49Nbv4AAYmX9HItDLBe+Qku1+5aZmsxv7d34MS7oL5k5PJ9mDNT+fcwN8
3+TnMbIUiSOguQOs2sI0XioNaKRzEVHdXWr8o0b9vUgUhczj0kpKwQck5eqf
TWcJLPuQNPaA/uAQaGPM+cuxEbJXS4IIB/xQ+w6T/sBosZTNUIb4XpIRRueX
M7/oA2UnOVn1E49f1M4yq491uaLijM/57NqpFSdbznaLXURKNvlNa/1rhMCM
5vFJP+rSHxfw78IH8J8pIxOjGToAQb4F2YjeEp1lmLFRSiuwcz34dYHDgLrS
ETgHClvplDPUGx2aG2meM+CrLCxt+wq2cqTXBmy2u57kxGi/we2iy4q+Rzqx
67c/YN6cI/C8uldOsJVbHpoIMZn9v8I8Aw6jLLWsSpOO/Z35ySMCM9NdNfq7
uPCc0yT6W0m+92fmr39lMKnJBx/FEH0RmzdHoHZkL0dBYy77ErWbwpCFDx1P
zTg3zTg661kYSaFB16gXlNj0BRi93bMvwZy1NGXrkKIBU3MvMxzMLrSddUiq
TNuJoxrpV5CEMO9dWfs3IpEe3klHHZB+3x0qOXLC++655cplDZd2lOrWuY24
a0/Lnsi640ka9TIcSniQJJNffgRR4PpZ95dnDEF+FwLZKf9fy6V4cB1TSuXy
TNypZSBvBXM+rR4Fdc4vzGOvggkihlMeltUxkmg5xATCeIuQHj6XyTkvxXOv
v7qeBqBZXdgsQTte21xQx8yZczz13v/kWmOvGzG0V5l8s6O3E7S2mO6l7icU
u3hAXICK2lby0SWw0vrS78FuFEzL/wKd3UG8j9nr0BuTR0uc5TbWfDd1cr6k
91ux0eHrupGCT7hi0S6aNCymG4WbZCWRdhp6EOM6wXdm2FKb81lm+eX98wRm
EcnrkgoG7h8HzKMahsoLcCVEP1BOQIvDkKgAsN5KRI8OnWs4J26dRigg/wYp
0LlV8vc/lxT74XHgkzpCvNDWZcWoTuynbGwTXjvdudaSs3sjugoZlunpz76b
2O3UK1VDIfppqg1xaANFRvKEMUKg326XT/5PMrOSCXV7S4sHN/TFP20ic3yA
ICvdAz/CRJIdU6huxIHzaz6I/5ME/H7l6B4cb5HKObyYmrBArQQtjvmCtERL
aTDm8sDxk+2F7xmhS374cJFWd4J4VWRGXvCSFDQD1LswPzc5MxCGs70GGmRQ
GY8SjslhdlMFm5C+HQdXw/NpDOOYLYenqRVIGLSj85QXvzNwFxdRPwj6NAft
1YVV9R/bKYVexrSqkMxSR8e96l5HB9wb/aIKyxvOfHyxwJ1hFD8hzhv7/hAp
1CUoIhdarxsX8goaii3lcsTk7eJTTGZccmhEoRkhr8ez7GJfqDuwy9zgxXyV
/U1jgru2t7IUM+qSYtByV/0Lwy3GtFcjh2gqzc//cTHQJ5NPFhjNuDrubwXw
Kbz+UDYp8o1HzwmRrbgJnDL65lhIRBPdqj17/HPZAKRjNdEcHP2+QYFVrLOf
iZxLrJ0CKKHOdpZEVB056nj92sznRiZCJCZOCjQptf2fJlrdqSAWhcIXx0pT
wfjNZMsr2cMwK8NDamnxAF6vEvXwDMnQvpxjrLe+h/HaNcm4T5hW9AO2f2KB
sU1JGeBv642G5vWnvaU6pkvYsvnjPEvUDAaxHxwm1uJocv/kuI/9fagwx/m7
ApGLH4Vf+agdNYDEY+JbyK5z5I1szVNBl8Cl3Ipnf5hUAq2G8oWsJCrdOteg
yX1iAbvrB23LcyOS5QjYuyAMFVE99F1UbpeQ0UbO1D7hCWhAl0+P71A4jjJQ
tR2MmWOeMPkVMmn9oygI/ZOopDikHmzEjjmz+uImF5x6gyyYdr5aqIrRWcqv
SoL+BXRSnYI3ILBg+cXkADBCxgE2l+JfenwzgaKG9XImMOACK8ivChmENkq1
a63C/Ud5gtDQvof4HkNLrv+N6XoaOD4EX/tDx7qWDQ866vdomepbk2fh36Ri
9mkePn8CdtYlTHvkJD5OFchXs5Gitxf/s/1n34UOjbfZGtglOeYUAepYACjg
9huEZB2eRto0XZ5L9V/SjkTPrmnEPlAidce3+1KOdsVHegK6HwfzKj9InUQE
MWP1Rfh1e2nZRY87z6G53JqcVFBMOIQMWsqLGcYF7sxQtbRl3rGegh86mrGH
0IsyuV2Z7pxAESFqya4OkAoyMxEilKVw+NK+Ugadk9vYlIj9QnHzWJzeqXtQ
K/0PwkHwL558/hYDbDZY9l3k+RwZvrr4Up6lH/EqC0Kp2nqJoUtWsK393XiX
r+h2v7sjGtOt/cifXAo58umP3lQ9TwU4tHfaBOcX+36iu6vH3MOBWubvk+Mr
GUKBsm4xBp1Ht19M5m+ebPcTKVAQbdt0ugVkFbL3K2Eb7l9BNKjuaWhkDWK7
rVmkelanvOKdics7UKs6DdY2xP78mb+SmHMbO0XdjrOtNHKpMc1k0x6RYaw8
LthgRK4E0UiTCLsMYWAeo1cG49eMtJKrNUZBnITaCdyj1f4Yd+ee+jHU+zAi
iHJKwjZaKBbZE7rZophDE6qY0ZWDu1NE+oDcpj4Y2E4Yhoms8NH8FrtSOXsl
cxPF1y+cgbVERlLTFCscczkdArmV5gqE1u1SOowQOkO801yGH1drkebfJQvj
Ihe51rJO6xVhni5M7RcCjGEJaB7AbZtdYntwgJgtV7dZhNE8W94tHCcvtbRg
BLxelkJEuoYoJ9hTt5dClfLBXCdOt4WT0cpOsIolicyYnYYiBmEnK5PBDGjS
4fAedgHLFKcjsQ+kO4d2kDnHi5jX3lxdYmjNGwn5gX6JS4ROuqFaDYlyupSN
0e/cvTGlMdJ8MjOZpXSrl/b3N7OhmdmYd+bLSrDTJNd0cyA8c5mDhV+Nw1Hd
GwSXiKUxUz0sw0WWTBelb1UUsJxD3E6q1oq6Ac3XA5z5ABlPxGkU/PWAHExn
0FLOo2IIy54r3w6RywEzSDBRd/FHvhRVKvUfTVnDL6LlVgegMDZBEj7jtsh0
0UxDD1bliPW5ww5XMuVOktOSkRNR5v2jjv/90Jg8Go7FvRG1MvmqyF9S5aLG
ReE8Nv/Z19DEe0+8pwSEkfSnOPXNN8ZwDi6eu+g3cy/Ab26mFBmvZMsouQLP
haBAOZk5oyib2NgW9qYu6bC23QkaXwCVmBrhd0SdtaI+EJgSJXa4IgZ9mJNz
AY1y9xi5tVuA/2HiPAcdeyeTYLPsD3xVUodvul3MjQWTP1VEpgeq3g4SiFqf
xsvXWcpntL8SeNJ8NDKarwxFkQNRBLZGxQ9+9Ety859XqGGKMh7BVDULGsej
TJTYb5FrKUcTFUkALJ7M2PAnzV3a7AciMaK2SkOBAH4lh3kViTJDZilRW+ed
mF1cYJ7Ryr0e9KaOZRWLxtyHhQbdb2c+zaZ2GOWCvsF5hELuDBVywWBiFGgg
zc+9/k0nihvfx5H4hsJjnywQxpnkqyfqMRjBK4WRykGyVOkmpcBv5v8xkvfV
P+OYBxIeFxX4bbqwiFp1dXZtL9X3wgNb8LUuk0njFYnpftt5Gpz5vr1WPz5B
tuMfcp1pEOjVuGdr2cnnnm8eS91UT35xkBbOBj6a35l3S4TAEgZ6abOkQ21n
gCcUIbSqbF5it3oa+Dl+QOEfdNmFZFo28RLbZbqQZFjom2c1GBsEbWu9BMDM
jWp6ijmFU71yyAS6dBTFYmyi5n992wiIL0xTP8BUV17wrx/5o/fQbJ3akG4p
YeS4GPSrd8qovxU2AlgrB8/OES1gmv5JbSzitLLiEKxRQHPZn/CR13m10GkR
mtoYR/WL8KyRAJkDxvPKvi0LxTQh8j9JqYlW8yHaTu+lwjCdkUpLvqMtOECS
/L/0VvSpM8IGNLs9yUDK9eCCeG7rp9E/Sd5WciHs09YiMpOn7/wuLOLbWqkr
Ihg+p2nmww7W2pPyaM3x41qla+LrKpnTWEl+pIbqWpwLYJ0F67GewjuyJmlV
wfnbMGTlI2a4XpGDPNb9ZZXfOGBcLkEfWaTVgZQqWlQ+l3tIwnhFeiydlsId
++9c7qbsJgtbBjV44PDVi+OljLElN0erif39emHdwwYUwiFPdiyiUKcCiHYU
Tl4M66w3fNuhYykQW0BwSF8ximO9RAI+gXSLtJ2k9U159LaJUeNQAPIfYTwY
gPzTBTs2ZHKsA0BY8OBPuvs6cc5YaNuQEaeJip0YguHu1PL7bmnawtOhlRj/
uBpDNlR8cz1xBRv3c5jByCD7Evn3pCVyOjtaivjtcyUxLx+lnDGwd0YGo4lq
QxJqfpCG/KxUvc+MNa1yayrWkX2zFKW/U1Ubeh7qtu/zGeMqXrP3VZVO1XRz
rpX+KJnORkiPZ4ihCQyfSHFvBlcHlX8h3FKnG/76tduWyq27R7vSjrJflJWw
poK7msys7axLabBkHHurro+P4c2Y4uT7AaZn9PbhxOzvtbeZVTzmRQd8ykiq
sEHUx7qrDMyFly1w/YwRLUhP0tj0FzSsP5qgT5ZLbr16pVlQTDqqiRLSWatk
IXVNV0GyMeu6AcBdZf2J3Q4LYzs/90tUeGkmXooRk9rnwwY4j2rfEPMNVwNU
t8YGjt8JToYoprLTtJuMMEX6p10NdhGtwBIS+1wIrxQ/zas8OnlJSB8EM6tR
96asTHCUR9u6B9b7ImYR+dNOJNTK6PXaNtRB/CfHtds8aQ4GfMiJ3G2QHc6+
TqsR4fNQB2QllLqJ0qzqDSMxlwTnuYcRxHc/UZjLGKZ8Uaur6e8tJVJF/X/P
qjZFK4vCbPMRdt5qKZIH+Ba7xw++E/02CF+q4XWNRo+JIZ3kv0zytMD+XgiF
7vFhcEuuHHnLg3fDV40k+vxhAbyv6gqt7EX5MV5bKw5lIoHFYhzUewGttu9/
t5Ds0s4A867AX7kTZsdSeCzoGfP9k1JMnm8Z9xq2KlGZntxQMl0xp8FRBVqJ
ANgQYf2YzFH0rqB2qezs9nYTUI5tzN8K7EgiotW+ojqqDb/3imYTopbNqel2
T+0xWWiZvoXrtO8kpzKVASYQP5l1rseq3lEdV4ECI7vEFAgGgNyqFR8S48jn
NWR4+CSuT3a4wxPVJ97ZiP8G+I8VvOyWwuBzihuM56rMmf9kLuMBRd/nb0RR
btHt/80X+gJmGIQnkWHxuu+dMgJoD+dt9NDcyBkisdq0SUV8vyJo7xvb+WQD
vs/wgYA3uXLnuW3c9+FGuxquRBU70t2XWpmtLoMPy0xE3dK6y6luUWGeH8aw
8adgtm4zU6nXF4YzPXJaCYRuzU5/Jg9MUT7M+tOdPsg7DtQI8UB1yqZpKC6K
oaV1Ce8ZCk2favy11BnDGLACCU85Nt3m1OTKELYJKn77tyH4wrRUYl+xOzuX
tkW8d+YrFMoBbqES/a+oHLqklR9vPg0B0h9WAAMo1G0s3I4hhdZ+iJCkv/d9
Ni/DCCgb/Hp84428wfZArvEeqakyNkVYs3K18Wjg6cv1ATUHIyDHiY3tVmxo
kW9dfPpB3pK5Brp2K1jAtnnlJE9RYIyF8NBZvfzIiSs/DQ/hXl/k0sKxixEP
Enj4mQDYgM/kDYG7244HxT8XZ8qiKCNpJ254+PQnwya/E/62xh08ZdNz1b0Q
MsL4wl6JKko/lNq/+xYiNOT9ZrtbgG19qwd6rPn6sU1P9mnECAL30Osbaeqo
rgTUJh0n1rjQk9/JXnU0O+yx1RShCE+F6EyVk0OsjPZAOeLxw7UsO7oJUrev
B2Gj72GG2GuCtRtG5c5f9s4iRjUoCPQJmW/OfI+MziMfI775E2I5o0ydK1AP
vAuMnU7ISDzpQss7ndpqUtijpBU563TNu8nOAk6H1QR0uggWng5yF8bDGrY+
bwSJZzq/DbIF5o0v4EnNKJnfi78JVIGF5XrmhEcm78WDSYfafnfvAdC7etvL
AXmifc7vHpfBNXXphaaHBKfmg526wKInidxQJrQ7Ys2kFCaaBtcb1V0+NHZL
7Ivv99SIDtzP1tn2izWJfeyxC2Nvefx5NScg08xUQ+cPfp6fzhQyDgJF1NP4
2zAMgnEP5VGsl4EZLbp+Q+/rQHlJIB4xxgjIljuL1JuURGaStLrglIjmcVBM
5mRB+Jdny2l21JXQaTPdahIOtQeoAMYqhdl2/yv3ByedCLN3uz/cvfw+VmQF
8i/ap6b1xe74prpLyaWlBO69w8n5Wp0E4IJP0loyaZpeRjWJ6/yuiC5wYP8m
aFnCkfBC36eK4Y0LNnIplBIwCQj9U+lA7EIxUbH9zMkZM7WSDhZNhk4+ADi2
EeWf86MOUFp5WYIqUDxJDVbPAyBX7/rQvkjhb/SGIdlF02YhQqJ63LfpGHmM
Lr6dNGjVjULDTvphT+rSW/Q6ODn8w0r2yXY7AS7aa+eLBx+ZGFpYXORVKDAu
+J/uyiGDDugSJWc6EQJpSeAw6c8YmI7hZVaqF4QngvlbV+1Mibg41e7kH9Jq
rQi9Fqy9hvQBHZKipd6HVpLToK9adlsbexFux5y3TcTj2Udq0EOr53+kHdqh
nvGe21S7nxBtR6gd+FRg0L6mMF6CfEe7XoheNO4hWO9n7bhz8edNI0pin94o
CppmeokyYP3zAl1EsY0BQidy4KnFDz8/vZJzQQdEMxrSCezggLgVddLlxcnr
Oid+gWBo3+RJe47Qr4oBwvuuT2Uj5TLBe5udrSZzAECV1oORRhcUuI0dGUjp
rFBZvbgaRE8DsOw7el0ESfsxu3y8kdeFNx9uNHX3UArtgJCM/XQWh749VQDa
W0qVNwBicljM8DA0OtkUpUm+MuehKEC2PHP4ygRYBvno8i1Q2SoaMvarwwZy
LyuOIcDuiR5DvZmvNHA+w2Vy+NF9WHK2pPZ/wrcpBo5V4yzJo1w7lNYORixz
uWw/2AhWJQmk1YW7LaZYYCkgT05/phhu465JoO37clztUngMlX/X2zablqyw
wsvbQBuZT37isSafpVq0rKVZ/Zij7dJimx564RvBgp6D5Co/Tar5f1QQCbVg
/J2ztGvbL4Z5VNhTwA9RWCQpgAJR+FH6/Lz4+tdqWWF+NlsteFG0l4QLPrjr
XAGzDesXGEdw7+muxBzaRgAvaXFpkaKgCjpEaEIUjjOwuLUxUoWEPMg6UE9C
c3qqVgHkp577r7DYAUELXpxYrrBdPSBNL0BohrRHLEpMuA1IgkA0tug4KcEr
5Iq5gcLbj8nJBJ7DNJh8q1C6Ka3+vts1vIrxcB4N2qRUp4+V+azG/b4jZGLO
nfl+VEMJ81KA5fgbdNufn0fxaQIvU7Qi5zc7fkWYPkPi4mor1n3qHkwdcIJ0
cpyQM8FZM06Kvh5wCBbbLzRespg6WOJN9muG4vJPTzKCO+V7NwhWTfIzM0ZL
8FNhgm00npqTKClEdvPTpQVA2/72GnHzIFrCHMQOcvfQ6qQMYsiyyRzXjzJr
fBS2u3qpYiVFS5+6y31fYygsRaoKjXkcQvn4yel1Mn/YhdH+9Fy32agvD8JF
C0v3YG61IMsk8hKRlo7NGkTIcdYajDJWZ5K3v4xdvkaluovDqT3ss9CROv/x
gUG8BiunkJmBlMT01FcjIJDW8leaWHNliWsxAo0/vaJ8CMWGAfcHFmipEhHj
hX2u28Js1Obr/gsEYqVKUtdBMQi5IH9CxUAPVJW/iaqHZnJ6jYWTzRfgLREZ
0x91HcJ491dqvdR6yJqZR7lQFLiPXtmFQ8OJGdLc30oRwNziV8aDfk5zzMTq
3OWmsw/IWS/HD4QKKM/SKiNvua6ZHlxel0fF7gnqnmb2qFPGZkwySmv8CHSp
wzDnnxwgvI1yEj5NSB+enTEFsHE5C1QcurkonY64Yuzsmp05KtMrj4h9CZ69
tqfuSul0u8smVyFyMUGbw/wrbFhyBvyYFT+sL8gtKrdht6TBB4wUo1lXVO9/
dWHzaZ0FL9o0fArlBZi9/EHNSG8cftrxGW43JYgpFB+bTrP89zsjPfxUrrAe
/py3iWBgXlEWqDX5rQoMKyyI+xIaAIR+qdCUojjTbm8I1pqYuoh1cstS8hqj
o2B4TZJ5ViXm49AcweBZy9sok0Xr+8fM3PYMWF5/ZXIqmeEnpnB4PKfwN7EX
lggM2z4Bu9BpxQFUjIemRlP7YpPANm3ikg2JbRR5xPrze3az/gXOauPSIAjE
D4WKs6nZTI14zK+Hl6JoreKPzM7KBUQrx8w+JUJfWHaA2zvP+EGig3oTM8Z4
zUZUpQdPGGm96z8mL1Io6HclVCI0nDt/w2sAQn9kNOK2YlHjNf7IVw7hxc0Z
NvSf8IvIJpzC/lFI8Nrlr2Nsv67eucQxI1MebJ/3RTM3HRKlo7E0UFMsFdv4
FrnXnQJ5qY/kmKa7EDCraue/TzSiN4lkyVnLSctSvQqHZdV/e/sHX85oNjEn
3kwekAbyq1+pFiqs4P1KfIZX9hBxJ0LvcJibnyZ+SwZNOG9e0kpRzcOGB1IK
wtHdGnBbi8axIdBqjwSN4gcR8rLHOYuCiOz1HkZbmqK1MfM3CZmcqjGahkLx
n5kC+mR5d7/ywS76zeBVZKXahcdRvyn6pYsm3w7SpoQbe2xIkGKON/U4tqMg
UTz2zmlk2YvV5b6R3UfSisayibuXGIYNM+gSG3ReiyYxeMDXK9G3XEhrHut6
DKUlA+5Mj7/LVyqRtfKOSFn2YYVdz+pqY6UH6BsWI/bxTDV/J4kz6Jk90Vee
TQhBJPZPd5MieexKEUbNRh4r5BW89FXlHaIdwpJXU9v41A4Wx3Xk43yLyDUZ
ux9CVTRtwIdos+GPy1Q68deGp91nDkaKNSVvZhFHY2X7qtxarsRhnNwiHx2x
Get4eJ4/RFqFeXpcsyOM43UChKOFP1E+r7BFKWR2RwU3YlPCrHqInOxWXnW1
SAAaqN9zFx6JP4lFI6ZcugfD/IX9tnMug+ZeNkWBGUMDDta5McSmZwomC/ZF
pYqoVssSPGFaYHIWAc/518yzM/AdJY+kmV39K8iCpykoVnALwJ+COK+ogvsp
eJZ1Dmn9qqnVHKA+VAPe5FrwVPyfqtdipB+RBp4kViO3Xu5NGDE1t3UiNbAI
Qs66bn8HKwW2dCclbOjFATc166g5BAJc8hfSCAu9W7m+2n3hitGzoGvv/Vla
2FTQPay/nDPbRMQz06EQF0HLuwSvG4Csmofrg7ZSPvETDy9jhoTxrjzj9063
lBy7Qi9w4Dgw8H+WFVLdP6Y/j2USj80llRJX81AWBA6F1dowsihaOU27mWaS
ktZ0X2fQAQj20hoUwcuJPKTbOr7XxfPkxcdFqGFNJr/Kld0+iODp240JXjvW
AV5dwaLAgl50lx2+ffgc9wk7IjfUxcpIt/bk+Wwg8sDKqBTqYHgpaJMk68k4
CR/CHQoGoXt5xTSx4CGOA+w+yD0aAHPXHte9JOErWYP9VShNlFbE/LmKBDzT
/Sl1p7DdR//6IHTIgoZQKN4Zi4NIFzrOqRBIgs/OuTGWA7iiCtxjITPPkIuZ
IKctxVdryh5FIxIHrMuoxSSoKyFOEbbRcL2Mxa5ickFyZosHykO9OOMV+TPq
2hsX8lIz8BkE9EqsWMkh1MQEmptwVbDbI1hKYtxWqYdMELpJysCF/MYyZVWR
UBTkEcqwgq0kyhg+OQj/Ny4otnAPTeC8ZDj4ECdVJ7V2cOj4AuTugkGiOseI
fKBh568MEIhxrPmuGSTS/WS+9xZXtTeI4aNGam6S+WzgM6hUB9pFJ/b5MAwZ
j40nhCxBlvHnW6su0eZQZm3IA1lB7SimZVzZiTOjOQlGyeB1P5N63v54D92G
TzRjIRQl86hxnuhkeo7tBhjZBz37of0a4XXTaXNpwGemcUWE6sOSxFTcUkDe
xt8lU8hxq6phk4b7oqpDiNlSqOW86fcynXiCIvjnnI/wchm4M1qOY0fq+iwn
uDCQ5tWV0aZeB6eY6yOQ3oTfdFMvrp31GUlUiOwl8V97YTjswLJKQDW2WGEl
8IlZ+W9+UGQqlYUoUdjjx9IdfdxTIsER8qUC254HEmWAg2yQoNzgQD9g8K1u
mEhFEM9J1MF8ubBmP0ufjK86QhQNMTsXfieYo1WeKTbNgK531H7ii4F2W04w
8c6LTMaJchwv2bM35wqKLN3O/bX8caY4sjJV82dPzmWMC8QCHDvjCsEYePJB
Fw8Xzg9GFypel9iQrGkaqdEwGJqEq7kZ3QJViecSkQpBOOIgvhAgI6zLIqjx
NXjyI4NVI+SfO7TZ5Ve+WQ1Ejy6NlYHXaXnhRMBsMOWyWyhR2W4hY40uohZU
OaUcyAJ+DjqvWLBMVPKS64LSvI/v+6634vAzpYYIqSQjGfcNFF4pLff2NC60
JptPqqA3wKK1jILUwRLH8KGyQCkZTNAakVMJOd7BISsc9k36AxORkauKomMz
T3Zs30Eos7PX0AZKdofi62MSTW5hBHlPa8KUpkfWJdLxVrhAS54tg6KLnbCD
4SCCcz6+ELbhmoPzArSSzAkTfRDNtRM9nXObjWDkZsCuFohCu/Mb6Xqt9Zqy
4ab7Y6ucJ9hUGWYjYzUuiTe9kefx++SX7B+myy65Ta5QruwkCpeSdSr/Usqv
8RX2Uv453YrN1y9ApFeTHLZY5colJ3lqgCGKsEQHuvYGyl6CUVki2j2G2zrS
vOyyU//mCJ97o3ElqMh1JXzjAtv1dy1yKAlobLxDVgNLGgu8Bc5lPDZCWpok
VCyH9qdsKdypKH9jxiCUQRvR88j6lAT2QPRO3OJqJgvDXM15ffzSqADdqrvH
24P3WQUlD0/Gh4FD1tJzDCDbKn9QbD5DXoJ0jzmmMljPKzSOXFm8foOzXxgl
2qHaqLxBv3aEpztIV1AS/yAWC/ueC8eywIyNxZdBvTWfmlkGmEqbv7ZsW1Sm
dR1NJw4vFl0Q+lO9ynVd40tsLIiH/QFucu1tmesfGT4dShS6frtY4QqW3Qqm
3CALo6dJtVWCcoez6mvEymZfshoQ3HKRjY0+aDmuAZ52zmvfhZTvfy3tTpRq
SvAmcU5tBrNJXEUqydQ0uJqKDqeCGzrtOesCqETLxiyRI3HIjv9IpwmMuQLA
39YlHbrFXP6IHuqfTSU+5b3ac5NdmRqbRVWoFSWh/dEFhfb6UrYt06wws0b2
2tV6uEoLtbBaBxWWK/d1qRg9YPoaXPKYPDt/suYIm5AzLEzectZ4qly3eV6F
sdpxxj2h2lONFBse0D1ho8FzYhws8woPeMwwrIZ3WcugVjgKq7E7W0WCkCoc
FTc2d73QMmckn8sxCnk604klhwsg6sg+oSPDZRpuzGnvGrff8cPU3MbuYkEd
bgIpgRmwHhwqSC22uEyKytuHaTMClyZ/irawEwR5nVIncoReTTPcaaXMvBsn
e3Yp6FJ0QMiPulws7iUPVSMlTlPHxxWAO9bwqbHotVsoQjdU1zmzuFyhoG/r
ZIvtYbE7j1jbHn2vVdeaiiqsNSnEMJiYw9UijlCUE/v+9EJreoURlvJxM9wV
tnYn3qvKAx3J9ahKZC8IPZfLkR2BSFBcdmL5hX7O3smMBfjY7Ia+tJePjL/H
GWONCLd5QFvKp/7ZQOkI5qM6PVVFv7jOTFDSCRrttepSFlOVc8ehBXI0MxhL
+b/zsqbifMdRdE4IjGvWM9DgjBaveB47r0vbJqsbMbiX0Z4G6NudfgYGyuoa
7jGIe4bD4tI8uG1AhjtVdXhN0P3LBz6nwiV193Kt4LtsRucproPphkQ3eyTC
Hn8dzDCn3sEpTiE9CLyGj6kOxDastnrk20JKI7W18cqlLCB2Tl68xxfZ4aKo
hyaz4gVk1rEnop69F+PiJZFmHfY6WO8r3cNJCCSh7gYInEE/JvnmtbVDgwuP
ZsNmJB+dRz7U1MgogJiGqbUJtJtsgtEbmar2FWvAjXZojbjpDZnFjtrtXnz1
EeHS+x/Of41Vo+hsV4UEnQm8U/alocmRUx2uywIILaIy5k9OiwErhEyGv0vM
Zt6MlFsWRR0OhNceCmRv9ckIfwa0Pqv9Gw8Nk8uGkQELovDStUkX5zWgON0S
C6x10DX9mPH+KvJGRYahCgtO36IjodoIbyqYwgxKl7Hnrb77QNRtK78aVWyf
zGi2jrpZk7rKViv9e/EM57LMlCsJBMW7GxoZQPPv5uLDy0ITBex4G5/ea9kt
2iQmfxh2oCQUlB7C5LhgcrADPKa5le/fZJjmmyXj1IKLAZOnT9UfodC5bjYA
SCStodA6++APnkXzCC015gQjQpypGeH8xDQxEVN8vN9lE+aD9gHjQfoOvJnX
KNf76s+IdpvTawTe+jksFb4coe8wc//KhPmpIiWYr5NEmcnbqFUUBvGKb4W6
RKK61GXwfYfly+HYJFehYkhIlPGGtz5jbS3VtJFkc+Q1eEmiKiOiotS07hN8
ySOHFGUkcn5dF3drCvlMRcW4aZYXbqc5D7oXFcU3rvkk5XUzd2X7n9CLjaeV
ZazFkf3Bgekmhc8IUr93jWdg8Qh9rXGapUKA8dWYi2GnZbSVVjEYWAoOSZ/6
cJsHLnmtnr5aVKVAVpNhkVvNCymXHcQnzQm3ZAjCeWkGX3Lmqgkaews4HeNt
ZY8bF599vy1dXCnbqd+aueb1D3Sc755LdGQhJkSGIOg15iVmuMSaNGrmjS2p
/2ReYVfmnh4GzujhQZ5qrRd/KWk+bUgJ5kYm4f+85imA/y/PwN2TgoNs48qe
Bji4uKkcuVyGocboYHHbXbw/mv6tP8Y/F1Qcz/rKehnX4xWt23dXNIuZHGFC
A7qzooDg6UPyS7ENFVq737QFe9qY+iVSklpYlZBMifQgbg97LhTE0xGu3We2
372q3NUeFcHiiPiInf1W4LnK2/jo/Lt8l7e1wGi4q1lK9WNhnUzrurvuLvsn
MeXCELy2ccjw0Actng6AqMVVeTfwRAN/wEwYVBHupfwczuY8Fqc+zdAXGacl
+hzeDL5rgehdNVFUybs+bwpTItZXWaVh0d1TtsTNEESI2hJMzAKOF71VDt/3
TwEWZB95hXAZk567JXeAvu/T2EkFBKnn3d4mjap/HG42DU66YR4bUKwq2P/D
ebIMZNB9nac7RuPFjsr+43Ca9flVVqHqHjsJZ8aBO7z7pAhPtggQMJWtZd9Q
X92rX0+QJwAwWgWNzpxdfiQa5fy32iUHXKXYQrrtiZu1JrhqPEqM9ZwqkpII
WQElCg2veRm3JrFoXP/a7zrPYsyQ1g4qQgnqg+0nEBq8p81DVdltrSqIxG7L
lU1rXN5x8b0XXc2xG9ELn98e9qsPas9370jaE7W8amGlCfKjhlSCrMREfDM6
kg1V2msLwnp+d1J3mRtun8xJRgoTrQwQEZBjab7zRUK8nK8L/FqhHDShDoDw
ah6gmgDwuUemsqlinU5NMePded1nyiXI9SaDKY0V39TtshNMJ/caeTiBo0jW
LZRfahhnrJY5wQSbq4YsKSaw3+VpJ5mE0RTrC3g1TBXwJ/jBDnYrAupxM3jx
w19rxcDHd2cOIxOLPhP+tum7QdRsEpT2Ze2rMgxbPm9TwqF/ji+IVrQkDFSS
DxqgdRnRciXtoxWA57mRqjcBXGEdNdRivQqvQsy+PkJTOIZp18ie3SkFz3ux
S1+Qa5aYjgRQlS5K9kxQeXLcqqjCLfdFQSvoYUQqLktvmYRHeaoyJRW/tdXc
LlJKgYHTWIKGUW0GptU/fSFJFzRhXTQRhBKisjoTLiJ3IYJ3RVRxt+GbenpW
0UZrg4sSghvgbKh0LOFpmgwCxrQ2W4dr1kCsWC4X+9SjXAO1qVceR92kxDXG
h6SgOpx0ori2Xq8I2k7D/CAALLeV28VWLK5GRfB0dywnHj8hRxj7WS6Y0tRp
xS5ORL9Qyz3vKJQz3tZdcdxUyfOCHysL/0+xuGKa1BBPslG3+FCgDyr+qOCv
Z4i5nMwaq0sFLLlePjzr1S43gfiyrTbHe6sgAXPT3rj00mf4TpuAZTRf/R6T
1FDDe7WCXSh6NKuf2FOW/lSA/WgfFbOp/XO5J75kxbVkkmzeQa5cHh12+Kzz
w8xBIKzTpsH3YSYq3KJc5hpRi3qaciu098HstEF20tuj+/4bfbV10fPcIwJn
WL4Nx7lXSlAFxPZjd/9KmwK9rqSRl62nR9EVXTynCFbj2QByrrhltFYez++O
y87SgOwHj1HKypwhgpNE0uMGuVwjY5iZhXt1lysnE2dLZXs6Y/fJmxUkHgPJ
PkJ6wJ7xkwIewF/x9XYAvyzKdZcWIT0t8dagdv5Qq2vECNsw7OAqnmE1Ip+T
s1J5n+GVb+wNGwxy7a3Fs7uJOrg0pp8F3TdBHiD/q/LCBYUegS/+Voay307/
Iw9LdBtHM1OHG6Y1YuyDMv9PZ4PkrssCafNWdx1t5R+LvTMAIPpslGr4oToR
xsbN5rAKgL+YB2v27OaFNn54ZK0KQyA+DwMPOGYXmOh/WFRV42ICBJ0u8sAi
40TilKzP5OyQpm9OpySv1XVPdVzbVeQUXt3hu7wNZhV713LukHX9X3LikY1M
a3hTG0gU07K0auH5Uv2rz4uN9HdTLW2wwQEQW0W+ELBj7vFQ6I25GlDlQPpc
yHJQfcgn/3RePjCgFTfk7fSM4KDVAsAMGn3kfLWbk8GOZ0k8+wKzrFleO0Oi
TEqi+/LhxBLuj9Jq78jH48swQ4k36OgJAoNDmIQ0OcDEtyufjBRo+fKNIFNp
s06xwshzJgyuF8mooLYR1XorqTfBpJkeY9JqASrtV/LKfONvhcksbOxlxCnd
garcmt0f6f3yaKjS6KZpHzBpdZK2Qc9oKIkufsxwiIWiKIgqQKXgFEFm3jVP
1Xb9LrNxVfYcDQdJKL5D3/j5WRojPJbmOLnLxo5ksodKgiQcvhX3R7HbOKw6
OLAMlFQrmdi4Zo00yb8IsRkQBAYf24tAJsadZEZzHB3DNrgHat0ke01dtGLx
bf8hTvTW0T7IUdJtm2Rh9zx/KXlog3lK8ENrFiHYQ40l9timcsRgGWjHofeo
d9wPhYeP2N2MwPFGBo3dVFjisKWG4pXYXko48VxGCCvcrZdRxFVbtGdSiWTm
5hSWYUFvXc8jg7m2C+WUVg2PVnbaE9+qu0OUeAiVtFRi4mIhT5DVAbVhTX7G
zR22aHHrLCti+IwYppfeMVS+hZJ56PzNIP0nusL4Oy0aSAHQeT2o2Q5g0stl
6log7bvDSEV4bTVCU/7tBV7ebIiqOuRz7yTvg6m5dzi5aWv5cjEok2wlI6wb
U6+zAns7RyaghsBalUAae34X+Bdx9WIx+5d9M+MZ8nPG7UzX9RFP6XFScsw5
cEjZWcsUXY035Nf4Me8YdxLAcdPyN/QmE8534nCoVFwdYeWjeIvMsQlyQYZl
gHsF4di5y/bFfhUttvoR9Knwu/TfnG7S5f4ggq/b+z6g5sOdGiYlaKyZX1Wj
F3FMxdv4mXKXePM3TDSSW7xq9PwI+JWgX+CesixbQ/mGEbn0hzoPa5LdyJPK
K+FRaQtd2HmHfASB54Y3pH5T03lmJD6oSO9q2X0QDvQSF7/S/xa4fb7Xf9e/
u37HDOkgssnB2nQvlgLrK44uvhqZpLSZdgvpJyujgRHRIhfk+T41Ixazz087
yrAzLfSfzjPVznw9ChmsVCzLCz4IgRJKcFk2JjWvq6EJnTmEG7uPb3lZlO87
0gFOe1VOH03hLCWuuOUyjnEnJATKe1GfM5JaQe9VcmvJceXjgm22LEg19CO0
0e/BdXqFoVflXB8xyuxPe7duOXppsfZ0mpcymp2tayeW3QouyWYPsiJruarv
RrXhhzUuBiyd4dNnMZmB73VFkX+P5q43EK5EXHjtNDWa9fyGfmMXVJfBJWrB
lP6KJecMVknaKeHuz51EtTI0EsiijhS1d2FBtsSGK48inKhYETHveSDLwhht
lmR/l7xuIyGDpwvlrZvoexY59AbGFAGCji6S8yWUCUO4ayonZWYhccwypp+d
6ec5wgqvYnApMt2aAtrZR6nGxHrGswun7DgmapbjZemQOWav48LjVjKUNaDR
WJQPfs2Np7O39/YqdnNvbSU4nff21uFgTdbfhrBb3gczi1/tir/ypdLBBtn4
WgmMeWf5x2o0meq00dpCcIwuEEmghFFaVEEXf+0WABpKYn6Bal5/4UNOldkO
haQh+X4LptQdgjcUTpUyqzwPe/KPfbokn2CJxa9yQl8mo84JkPjKPbwKtqmE
9tZqHZAhGAp5kpCni9Wz/Qn2VL0DzG1nPAjWyuha1iua42l2p1nGUMYOhrXN
t6h3RwqKlp7ETnR5bdEzAjgIK+WpQIwaPmeiZCW3TSLqgj2Ozel4b9qHIdpl
JLsd/if2q2bn0LTMfV5/z3nwVdzDwuyRBIE5hEiYRrwACAJXKHpdlT7s0hMK
1yQPV6Ima8KkHBwLdID/YZTs8u6Mii8AQe4elpC7W81vgRXdzZlxJDyYJ5Z8
ew5kcsFvXP5gUskmxdFHhM4h74WGdEdlNCetLe96eBrjDXwrT7gXWZJt57Yk
UECB3V/CwM/QtfCv7ypNK3ScFg4OwvQc62Lv3ikxjIerX17hJHa7cVZQSSkv
byp0R/qpebMAjFVGh5/MvqdIBjLyNy1uJgdJrl+ykr73iou6OphXfbq+A2Ga
7PLD4/bTVncrbcDNrS0G28JwX3ixDFecoL0y45H/GRWAmU5WdstNUC2Ec/na
YMxJmalAhBwQ5i1QLYksblx5/kiKcUj7IUIhukTFNVmao5TLC/8QIqAPRfdz
ZSKrDtA+4YZLmCcpZTCui8Q07/a0ysYybrl52gsCRUs5DEfN12Hhi4MY1/rX
Fq9pnimmBKOpKEBfxQpk1PYlHKYrs2QOUGLHgJVGHLvzJgqESzga54urYr06
5zuocUAzr3EUY1XGE3FmrMj2otZWjBgQ0Ek1YIFp7NiKL/nwjJ/+BBxlqyk4
auTkUEMG1s+6x7KJJGyDynDBxPOinxSaJ8tbwH8CBW8kLVntg6/MmgQ16mtt
BJVeEifh8rtGWWJh4/kCmMLecxmC5GMtg4vFZA7duCjQqc/aWcvpldG+6E10
R/0YLKvZmkpaomuwFVrMzkRRf0MC7abX4MDO4T5Fi88TmThwFXKxesBIfCCK
xROMMOdohSyX942tiD+3Q5MujrUt8MCqQ2/xOkgb64qNO1TqNOF1XhoXjH+g
TzmrJZ7+aeZNjVesfazJmINEgXQB3Cf5cadgRPEyLvxVU3enu/D20GAZfZ5S
sohdjvLgGe3NE7PfSXnOlHYqVEJxmu5RoZhYNALXFIjSEaNFuy+EFf9HkmM2
wrSmdD4z549H6nu7ia1ZxEY+8axMIo390vPoJ8b8evEYpz9v6KcP9VTims1r
KMxtKr9TJk7G9nyepJldIqwKCo6FiK8opn3Jkl/5MwxLjMssjHzGvwh5pKRz
KUF/gRIseaIlrVSWhft9/DqS/3mFcc+t98fIq7BEs0sKsk8pEoBiQd0ILl9W
S1lgnERgs1nn9/Egpq0xy1K3JTGNLC3+JoDaAdZIJlkWlWS3s5YnRqPPoo6e
S0n++YtFDpPmcOeB70+AT4Kf4zH8ISMp+HWFA8p16JXFrg/DYVDspwW9mLuQ
1AEEG1GtnmrMV0gHQr0xvxCQdq8+vuSGZoAWncAEg2gQJAuFTvWzEW3hiPSu
6nUkJvDHVWxc8QjCON1mQupTlOOq07SCF3nUWT77KCAiB8q2+XKIRyTiW4u9
z/uzyYhejQb79/GC4WzJs9zZNOqdbzMD94QpLYtkm8B27WIBjzgdDgClQY9u
yiZ3AwkFxBMZqrnDKXpIRWB8TpoiFAm7z9BuNUzxlwrX4o/s3l+2cXVv2sUq
Q+coLLhzclWiv7s+Kg63rugu0keZ/2XSeRtMDHH0sHgJwjUBely0WoezLMou
EPBj1/DLsI8OL7fCREAkWRYHkdL1YUkrvbW14baByDx7glf0X6QEgzqSDm9c
vu9EnK9Kc0VRbXQVM8oV38/F6zLEAB4QYbkdp7BAguoMGa5AaQRK1LEHdqKB
FbD23yVYVaZJ/PnDS4o8yD+67esFNM7s/VLnWsbeC14FjJI5ZMf3Ag0dQeDb
F8uFMYLtr3vf96on9OBd8oqLwVs7wBofLkU0dv5XHNQohX+afX0RrLGlvac+
P3I6rcr2j7TBS0pjvCf7X/8YXSZAdWR8Y3Em7fCVt6I7YG8QPSGGpoiKvfyf
mhWSmcuZpgpNGdSn/O/OhWGwRKkvkG6PO+WtpcEpUY6mmRK7WdSY2Z4VrnVa
IK6KOMPwDbL25MxKSz/bbOul3pgrqJ2EsiF6RWLB1gYSZ+tu31vKzW5djMgv
CNSEPKr2u880mEAUx4r5KwgOlwUeAdudQJ/WQCcgrrudeqL/YzijNkKA4u6g
jX2iW2wxBiOWPPjIjZhd0qJbGsgXcO6gxJsYi6s7ZdQxAwYYlmg7Hk05E0nR
wHg22tfnlzy3Z0LtZ8vkkrSbKr9kVkpa1omMmi21MXttAHCvugl0Joi2UXDg
2s2q00ljJu5hTy8JChYlmt+kVpaS9yLluoNztA7WODf+of3ktR2nOaXiFIGP
wC+TtZgrZW6Ngr8avnlkjKi3suV2DQt/0qU/KHud0eEH3KPCCJK2qdxo3cDZ
SWtss1Iti/GXBEsOQqtaNM7KeQ3971R01EZs7m93YX91At1AhRIprLatTmk8
EpkPqz0r1A6p9D5hp+SrUjBYfP3aq7RQza+E8a2ZvQYV3+it8wMBXEAWUiwN
VpOT10M4zdEFoN9O8iE/CL/mpKxhvjDYIwAknxe+GxsluTovkhbtIYbLlsil
tlpLQs7uV55CorG5HWqKG42KYSIlgZ0A7Ul5WCfC1WcRrpuK2bZ/eNahZwGg
Z8U6yxBWq4wgN4msQXkzDWofpMt9AX5eRCQEu9ojVOzYO4ezJe9gBU7ZOBze
wj3Um0pb7npnxab518Iiyl1X4Y6b4yvIH/bD6RSaqgte3uTP9gnGnAy4VNME
/f6rbSBLZjMjMHPg3LTrBTv/V1+EtFJYoDoCdiIKcEBFpB/mID+0yBMH3rQM
hPu1Rve+fa06bwupJbwB1WP1BnYZbzRzW+fYZuKdQDw2tFRUICiHI4PHD3/J
/BQhPKoKenr9398h7MMCpYgq8B9qX1YnMXHgfbHnCIaMw8Yyixq9cKDTTRhE
/xRPQwtBJWCUIfncx6N860K12MnibhOQ/QBwfYjv9JRUR6l3ELjdjTDP+QBQ
PVEBnvc5agJpO+b20BBIlYJqVj1hPsaX1xNTz0h0OLBy2f6lH25g1BnrCCW3
nkrUHWmV58vDXPyYI6JMIk+Kwfu2k063dNhFG2knQi5HJSv35uoBUt+Q8Cqr
EJpbl3kRR3mdAQOp3Zqllw3oiIfWsO5Iso44FZLYPo4KJ8IsBj8aibCAeTVY
U1lBfaVQEi9r9R0hhmjISnYyCE/EAzQpjTtf1oUJ9/LroefkVe58I2/RfVkk
CiVyQZNsW64GQugWKTBhyxG/JTYV6RFueqN4LlUi0qweoDBvX1KVHSHSVYhK
FYr5De2XsdsT5EFUrdk+X9gywAl8bnpJCG5FAum2VagQxt2CgS2w5OZMpnwo
+mKanirAclHQyqkIFyx5FlTfz8V0SlmERMD+dEZz7GW+avMPbJ6imahLfvJ6
gzyqsces694agpxqic2Fx2l/bH2p3X23M302b/eyZA1NjV6mE+1vZD+/5tWe
BAVuSzZiZFv6C1/ub6PouL7g7BivEIBP0qHjYM8qEtXIiiVac51kv0iPIP8g
XhMK4pxGrdLOt/D+h9nOp4o3Tv87o1mC0ujx/OrKm5IX1+XqOeuBhyUX6Rcx
30kcQm4A0AmVGf4c/b/FKGH+3HUPfDfmpzKvau6HHhqd771KcOpzPbsYNfwl
xodQYSBSEgrBgA1Sn7kTPHankVHKsdWgigGrdweMpkkwCKa8ST+rIe/CWXR4
GR19YhYRfgwQONACXTDx5uS01+Bnf/EMAX9Ai3BqdfcaPuO+mEAaPPdFOysu
+d06WVioCLGl3pYlWg8jfLRyUfHkZJmt5yPZ//6LWbzqloK7M9IZGv/AKcKZ
Hl6t8SLUQJYTtQxIIzAtz70Pok/dQockT8MpOyEp+VQFsEfXHtWpyGmEzmWi
Xb1hX/d/pUQu7B5xWzzYSCPAgDEr9gthYrBOgiBxtatUMB6IvAT1gydbH9UM
c0d5LUgtJpi992rQcji8I+WboMaLkjHLrdt2RhjvwSpquH3X6E6NCmSP7kil
xtqSJ6mftlRb7M68Yw8lqwx2mFlpkemApTw44b+B6XHs6E5fXPvDwkHPQV0p
sBjUeV8IGoO+xcyxjSBdnyeiK7QNYEtBSiYAXmARX1iyxyaVfN2ft7ofBmt8
DCDBh0AiJtTTIlbCvB+rYlP1xq30ulAXl0w32IERZKU124ydOgDhm9MLDayF
aNPb3eNjBmfqd1hJqP7HEZPfH1DwdVhUC1u2uNtBxRLm618waLfYHPlUPjHP
VRlHOgTDaJupxV4Q+jRYysQqfpNkIbhnHLs4d23xZM+365AuqsIFKENYbbsI
ZPs9SbS/HRvLZhUatgZCQx4Ugc/DwYqebe+Q/YFjrF464nD23Y5lHXbPisoe
omp3PMAT7FohfuK2yffCsdrtuPQ1/4qwdJiT5PAjMhE87bFvk0slVzWWaFHs
Iwnk4BrtF/xAERai4vLeSxbkkoIaqqdpsfkTU8xxUAvcfWoynYVtXK0lqvOw
BRxuoLr2PNNaTVGx+gKHOzpbwDhNt822FPNAJy2T5CbrxY4wXp+yQtf0/kkY
ax1thX637ikiJIwnc2i8MrL9/ozGt4d7zZ8RA2HGk8XuoOKG31WBM7Rsiryx
rMNFPIvfqZJcqzDGPXbnXhOejXnFI1s+E1R2mOlR5E/YUEBTrxNh5PVUyQ/3
o/cEetC6CCQe1NGxOXn07xJb6yJaTZneQKqgis4KfA33NiC7SssLkPl1Rp8j
vsffgv1/eP3SmScRqDchxywChYjdJdFWxiQESW9JGYaVEfJNpeJhfMkPRCqz
lQy79q43GmKM+XapsnipHEv+lxHaUG+Pt2u/P/zmc976pDcFF06Eoc5UuSou
vczuPRgnhp/BE4ztewYGepEmQuM+GYdI1YBHaWhGdGt1P7rV+trxBvKT/ozt
RF9MzHBhUJJdhTkiPDkA9L7e0reK3WthcOi7ZRUEQLMIPCSJXS4Mpv0GJqM2
yL3fhTJxxE8T19M73o8GWD6A9CqUT8nGEU5WAIGC5jamOr4a3AMnMG1BAAkh
j45ZwFRMgprrjZDvOscgXMUgN7il94Ccxd/Q/2KdKwOCt3d5eZR/Lw2CM6dn
VCbN74Y+lw0Q5ZN5AjFrpodqjnbpp4En4Ngqjg45ctXJyNG8fbG0eZyvVSF1
yfakNSFkWfVYRxxP2e/lbFvtu/uwbeFPhvOxSqMcXPE0HmOHLV2VNYeLhtz0
OXTQlJvgzTHkmYf9GG2U884hCchnCXjE6bYhpZH659BQISBZJS3kMXUKbg/4
4Fs9GqVeEgNKviovtEY4P2K7PJLzXKDNoLXPDgoT3TcymH4woq4z+37dgXuP
Fy67hKAnL/f5Vo+2+dUEl5rAKUXaHfwAMMeiKEMsHLNm0Ztbi7kuRceBedZL
FXNO/LGLunoEIXUl7wptYsh6X/Rrf3McKIqarq+CQptDex0JxLwQEQrE+Wm6
Sj8vwkQb+kcXJjs3cBCvXfLth3lE6ClPZXrdAu1ylY8PR9PmdpXc4j9D5+VV
5GqHA6zLS/T87zmPcDrGvxywZWG+D/GuU66bdERz7lMBMhg2rNz0jyrDfVbm
GiY9J8L0Eu6Ag86O5Y1eIf+9gu+SE8pd7b5d99vkfcwEFK77W7rNn4NbwRw0
Yxzf+7+ORUlrp5yyMGGd2HxZTh1A0U+3oauCVJRhPhpwzLNgx3ij6labAU1V
zkKJgjUmPu9qFeqoWFwSFir+khRY4IaKjOQxl/E6R/LCzPFAid3zhVOcrEhf
zR1sx4b4PyXl2CKmAMmnGcEZid96zb+B9UKQ83qoUZ2W0x+fkpK19sZUYvAr
SDJaa9RlIpO6yEiJWejeHp5dwT+FFk9DLKBKtc/89p8lKxLU0r94KkAJrM6U
TEIjkoJY/Js8+3Rbumeyp0N6brjSSTLF8HoLsxn6iQhBvmjG2EXfpxDV2vRa
nBShFJBOef/AIy0kHFUQOpQje4hj2m02MU3qA+sPw9c+33AlNKoAptaDJbaH
t0RIXEQW7G05AC13iievoPWKZpk+Jjg9vnmetoi1QzJ3sjL+jcVhx/LFZmOs
bTU91fBc9gIsWoK/7ghBuuuKnlZ6Pk1PManZdcOYC/HLz+UfeCNicVVLlZE3
KvDFR0OtNtwCQ/V2IHwRMHQ2MicDvdfBfputtWOmvevDvnkzoU2CA8aP+FEN
spYXV2I1kJaB9AqFAmAy53ndo8Bxv7/uYFyXRgYH67aiXZQyu/KZxo2IlGJb
ROsVyawZNsZXPMgMtg7hqyp/ilc4SQ20LO4aEPtXh/aiHmtgUIF7MQicAOQd
jWBkK0hOfC8gumNQvbVJQOxPgN5/A/95aguB5zcuRj5Vj6EOX/pzbaV1+86+
7D8ILVYJj0C+5WgZm9EbX4V4q8R6IgoDjBHCBYKBRRStGOR7eUO+6Uobnj9Q
8ETCj3JSPpz0fX/o+4wVa3MSYjDNhYs+uTyTR/YMzjqkAcJ8cva1BEb+rYAP
3SyPlBE1WweqZtgzfxIdAc3tQGb/9emd9in1dsxzICaknqI84JjljHmBeUS2
gutj5QguetrSYn5dGH92DEIBXP85p9iGof0nT74r86XonRTfP3QPfMBg8/EC
ZJ0fnslbMb0eqxh0HTP94pW8K7GUihjBO2Q8a08A2G9VaV9O2XGY3Ap3mN3c
cCVLfvhKRy9XI2lUpI71ZPDF7IzX4JsTi9jAMVcfRrqSC1Hf3b83zeweP2YJ
xTt4FIaHsxdu5kGVIpEDeXAL2RhG0QLRJpSJ7CO3RrPiskjdGyVrugdC/75g
nNKVfBunL6Ofn9EentiQpmN6JFvhn7N/ER02aSvuXvvw9wMrhppRT2eJuSZk
v08hiCEyRTUisc0gpK3F+uA2rllIEOYMTwznrqojQM2RmmdMfTmJUnNTp5Ig
ggLWRdqKi9XmdM4HPJV/r5utPz6i8CHGVfWczzOlXFeH7w8KBrBZOtlyx7+Q
meEDwm7jUVCwjTDiQgK8CMJviTlDlSEdBvBTFXmD0zlo0Uhr+y9nCgLzlUhv
ESy4jIojFDwKZ9LuvHbSiSrw1Z4LyclgZ1YvHljuuiNR/quG87cqeSiQrpfL
EsxCUHTNDwuYwdu1TofciGJbUBoAmD2ZiLJA0zxihkYsXP4gu7cCS/ZLfP+8
M7audmlHlGyjICIHYEjW9XviETsFKMs/w9XruGGf5JFX+LitLnf8C3vEncYJ
vveaL92BArhfd+sJ4X8OajdK2cOdzJzzrjKl16ILlE7epvMyW/o1EHXiDAyQ
On0HwTg3RYHlPcRw+RyYevwG1NJD/9exalsAeIy02bwILVBvFIq++P//Nxcc
75z1Hf1kZlDffdC8oZwBWb+5k1A2JLR6WvHJnu6gWf4b5KXUchHpaGeszRAD
EISmYYJ7w48KBvQuH3tolLK2JAQjLNrd2f/HiCwS7I4P7Jia8ndbVfPR7m/v
QDgITwgP6+RaGrIiJbg0EYuQyteK0Jyvawd6q+kf01InIFGertstN6zxyZYM
bw1edUeQ9LyIO9IDKz+nUFwHBFm0lYuhjKI6Gs61VtvxHTXaIkJ4bQr6zw/R
0n7Ybj2aeadHRPVbCQLEG5Fov31dxx0rlHN1QKHOI5+Rt0RaokKFSmChVPFi
burQ3zJeblWGC/4vCEyTABKM7nBThcEpulli/b8KMcNdmK99brXHIFIC2CgX
hNa5+SdqPOiaMtYIkefJX7Ujoo95dreH61/tDleTrFPJvfvrSWnlIHO765vy
8c2wtaZEYbc+oRyxAwn8iCOT781TpCagFOsdJNtg7Nc26IPo44O5szX9IvhT
lfO0TWk46ugMbrToiXusDWsyHmk1vKiVjQOCwx63FDfzN/vy9mmM5+VUXQ/o
u2cM1JjQJPxvm6xlU2FMq35wfCXaPoXn8WG1xDzOmHanlEZuxMPCTjZi4Q5O
UpbG4eGfPrRgMEB6p9Ch24E0gk6tSRi2L3xZBCwmoNJ+tGZg6CbxVzAC0zH1
uPYK5M9nrjk9D9IhoOMi5dWY6xoKJsmxC9RVAZtBrRhSIV5m3ZiFuoOI4pSx
s/G3XGPCxeP6LmuCiRYhRF42G6J3Z8P7wBg8AniTtNyValVocDcEcJAskbTE
gVzbogHkJIiHtrGFNPm/7gUqG07VO/VIVNve/hvw7hAcHctel5PZ42m59tH+
rM/F3V/fAF0vU3p/4htzbTLR9Y+VaYXge3lmCVHz9bOZvXnMUiRj3gXlfhQw
oy6F1Thx1gwL/6SGVp/imeVYMyhb4cOA6A/u6zBglbcIsgHBVCmB5c+d7r8p
1cntMY/LffxAcdwZ0pUHxfNzXo21YVJpHhN6Z8Sdl3Iu6TkNrkWpLL0E3DXF
R9YN+jX/PUbwCieZLQ0Jy3Ki1ZOtyKpZC6igN/HZdk6i8Nuhq+1+jSFenZRy
0G7UZ0JYZAhE/Y2z1pAfJgWRi39ILPnXiviwJhyMTSZflFbqdECgjL/tBcaz
NslbwiZ8uLHiigUbzRWxxrBwtBgRXOzUUZvsX2HzbD5UZ57TbUiFEb69diSw
7pW4N5I+XbUf79lzM/vqUofGiesEyy3f45PzdkoolCIGddCgs17rEpNwOe3R
cle78wMKCzbD03D4VMO+Q9UG1KiCN5RSuHUJAt7kb2uJ31LsMMkxI1oNV8up
/af08ldC5RVPcMk5SzJ9SGnuPKC0vf47r2x9YcdHvkZk6Ughl10Opr5uRWAk
5OzmrBIb07JfuynhjNf6yc6OVdzX3jC3NED8KFFVyfu5lvVD9aA6wJ8YL/ux
p8qZi9GuWi3296EdAD2v65Gjv0oMsm+05JGHEFwBJzZKraxKFqruBfR8kyYd
fBon4Hc04OlLw6r5hCeW0oS9bSa1RMGDgCucyxORio4IMS40YKWXILjRPNSu
GYlps6FRslnkiF8aRfB5+cWG/KGLvjJEzYrkfSbdA8vjlpDoNXSTssIEtATk
mtoSIFDClYUpwmDaF0iIC6zDHYegkwwMfVtTn5knNAuOIM5xhaCvyfcViSeM
y/tMFLe1WxeTmSdFrww0cwvD3oykmYYNBqqmHRJrOe2umklbCJfYJJ2B+uYt
5PlyJ7y24TTkFVnHLB1IrvBJ+vnvkQvRQ50TAhyMA1DvaJVLpHyNA0FIU/py
AdPj4L4JukJCIcTigL4OvSdc9S/pYMn80tfC8spXVf5ie4lc0hEOFe5CEFPl
hwUw+sL3M3p9e4p64Es+hnqSqhMPdzldyJJ9cQVumob7W+QC7sAmP2O9hzyV
+ZnF68chpZwNbRglIE5TM+qX2ZWhMcrYcgYRq5twdW0fdZiy4Ry67iFsFVsB
/zcYnWCqf17BtXASbpJtAG6p1huUPEIbB/Dnge6UKfiMhPF05E0gkdx3TRs6
itC3hARjfaZKu0tMr/2rnE90iU3R2WuCePcvm68Q5ltyaZpiS11vpIX3pMyX
vfr6+XQbpnHILlgN446eUDyYvv5IK733RqZz9xspqSC1vN4batdZy5KgGf5+
9h5fpe9fePEyMD+FGQfFyLRciv9fBzgp5qiTSJC6u7EWSxlXSSbq9NYh6p0Z
g0f8X9GEr7HKL6DeIRn+Eg6BFkf65po2bHb6+RrBR/c1F8/vGoMOQGs54Kt0
f5J5UgB/zevD1GqMfPcVo0jHcNrqhgivEh2lbbND/5RJUZs/idG9gT7kOWvF
Sd2Zli5Kk0YNDjaN2+uZBuufjL+rJU6hNgsIaTtwcJX60wFq+3FEET7xBDX7
xK34rsb0Phn1YKjIGmjBJ2pJ+DQVKPCe6GdMoFWGU5k3NkKWYmUuPJVAt68F
AdHqpaS8d8JYHq9rD4rMgXVmyF0kKwG8Xz9211vAMovoPDkbfScqHDsfXtvv
v3/ROctmA1OuXvGAy0TDDIFNt/l+kpB8dkrHTJv9ecM+EvtezWFLPEOfK2Vt
t9rA/cdj7hAyUXp/Km/HVJW7ibDQK6ytnXW99g2C0rn2Gw3mChLFMbPHHyKj
6hI3v514x6MPM01Ay+k4OMTTn5JvlTiRkncLoOgmMvBciQ81XMtAqjReN5+T
uaG5ZWv8UNQAsxYHlEB73VfcHeb7cx/eNC2JnP7/silFwbMI01WLUgH5/oYB
yGPYD9UESEYVjvK/f1FqIwvuaAnsHQLmxZsDabuCllZSNe/Nh8WqZhw+bQmh
oZEmbtaAme9hA9PVBSB6O7Vmsi2NKwgl2QjG7h/2lV3vFvj9rxjX1bbgkKbP
FtZzVVDm19BP1Gt1FnTVea9qwILaeqeR+rvwwIdKm92GNcsN33a9ZL/STYvo
1oqz6M2K5GzVcF3wGqJ+KETNA30eWcWAW+sbqspe8fZIcxx7D2fI2mh+O11P
m+CqFuztP9Cpf3Ld0egc6C0ihOzYZml2xlOcL/DXdtlBuuyIv5X/uEs8aJaa
kjQFmIkn8+3Gp829GVTOfH93HvQccEYtd5SkrkfeC3gUyh7QR2S/uj9qFygw
z14olv1x7V8gwAawtMEgQY+ORzdO/HkS9JA3NAO0xx4mMXbAz5FiOhJlnLy+
ksLLpMkkW0g9oKqWIX1T+D2tsZmg1yKlWnNkhZ3yTbBFuEY7u1ZvaJ4uBNQK
ze+ExwzzSeN1PWVo1Iw6b1atZswdepxyfYXbLx2c7gCHaNqFjE+1Q8fP32Io
+QL7Qtq766OzBTMVrOjS+YdUt7ZC+oNFDR6xNv0SS0vl0YI0hFhiva5ZVHNB
SULDQE7N7xgSgEg7g0M85n28nVLSbxBLQmfrTFEZYh9epB9+sr3lKEnnTO4l
1wHEWJ4b16hOn+Labs6fCsDTKWt2THKFIpnW8TmK65FtxKSGWu58rDbyRGGx
xEp5XhCvGOLyJ+NLUWjZyjaOiJc1QBqmgQVyay6Di7pgSk0xZg2GnK8m9/XE
ZgWzc1KspO12uR13Bwx3zcfEHmN393DExTHGNT8GyNE6dErWAgFqnV4GuQI+
kEeXWG9i591f/nVQNO5giVqrqCiUHCygJJnpfezlwk52RbBv5noX/kZPMRto
0LGjRSC6EoZrFmxhvgvKJ1CYwCwq2Q5YCjd6bXiDNOtcEbqhpJGZqTJgXMla
wQ/k2ClqZiKcoRwM8i/1FTwXnFe6/Hx6MVvi1MD0QQolXrrQ4l1cqBPM/BNX
FTGnruRvEH4DqGE59g46doMF5vB5FxalyEkF8ywcLiUuMcwV6YUabl+rXb9e
s9dZ5ktOPlZBW7Ori+2MuU+KinmWk2YMxkcYnodrpV89dK9Ue7Odh6yTE1Xj
ZPRRfOYDKmqlikx8CSe00+M8aoSPAdOPH3oceKjcIro6MgHDnBLJu2Ils6MZ
XVE+I5XA1g5JzZMUCVvAmu4l4eDGkmlobB/jjo6gw1MSNkBgPNnoFtgnOzXQ
foLEUdlmTCXY96w5uhc0wReY5ihLZpjTQJKn27XR/lDpbT+TB7f5B1qhyxs/
NPciFjd4+Yo30N1TEvzlC2GVBopDlhDVIGqo1cTWwkxDA1pbz2Q2QOzAov38
WJnsoDlbFr9TW0UO7hYxhKlTnUdfbwlVsgRiIZejF4wDReSpdctS/oKF4sJS
BMviZ3JI9qF1rviKFaWw6okcsA6rk+DUqxKhGXW/DwOF1JEOvogf3lcBjuXI
6eG6DB4YNDKiymI1hunnyJKcYv1z1OQ3mxnEpJHvR4nywcviWsySbgkPmwdz
14d7eRBv9IFn9hz8ccG0wTf5ACaGXZwSjxByGGzMDv2DP9iQxQPdLWaNTxX9
IJ4tGhf9R8DbLxYZ9y1oPa10Ls06uOPFOLtYSOykCeTpllJzY7c9Vl6qmJza
99Dthb8amvI/l9yIEbripvxKsO4pEpDkX+Mops8mYvEvsYTkkGJEK6ztM3iS
6zAu4PaYTCVACydBz8OzeRDfaDrEIaRUWwk2FbgKYALHl+95l1KWzu002XlN
7vGnfDMmAO+2/zIvjUu+gDgyEiiGVDaJHWPgYOaLgetYP+Z5WEozmBQaJmPM
BP4NFYfbDF32mg/q7M8sRzNQs3PVJ8jjrauh+f9SanUtIAcfA4SI+LXZvBMl
koh0mQwZ56gOE/QhKkLTT7302RDOWoxJtbfeoNGecT533+HQDWTNC7Xe0cmQ
Fp5GM3hTR58xu8TrpmxYVcDa+MM/xVjOUmcRdwB7hq/QlalGfMD7tvE21Q3E
cVHtUip9kEmX5z/ART7ZaZBr49E94VBcE9xtaYSHc5SMLKcFE5SXCFc6i8RU
NzmAnairy1RdRcLUOclp+cKGvc0W8jUeyyhtIg9utrciKGJLMUxlxvmlBFOI
+9pQX2mdOEUU976gBSNBy/8zAlDYOEZ2A5gcA/doW60O6KC6K8lBnnY8cMYQ
Q6NHFskyNee4iGQxRCYflpBtlyGtPUscCcziwCDnwcdD2LoAp9neyrbNfPa0
S9h47ZOHA1JWrn/YYRupRVgEycBu0AN5omzozkUyPsUXRkiJhrGoPb9xxeuE
y+QdWf7iPKLW7sCN5WsAm7oy+KJXRmywJWLglSm77n09hErUnmdCX32U/00N
BrS2Tba9nZ4uakXmfZPo2oyosiAjye2X8GC72aeZAv0rjVkEOROBk6WsVkWh
0kZi6bJ4pRvFHXM7NMiRYrItMvlpcSSAW4EvKGVh+w2Z4diIJwtN+EKGaTPE
Qw/8uPTs4ktzUjHUCEbLzy0tU5wvE326cuKv8LYIECGkGYevMEGrTYCcqrD4
MRynu5IGeYNZ2C4lU52G2077uHHvIHoXHb6jBack1D8j9l9rTgLLt3zyK0f9
OBUdnhzPQ948XHLrm8I5gNaj+5d/O+B6tyutDrAQm9aObFFKLdNH58KbZ0Gc
Bv5EY2Kydc89T7oS3gnoe2XZ6EAV19UoklIfjb4/fzmtxrrLeVvmRyl1a9lb
mw/iD3hSQacxIC7Yp1TvDqp91MKEFUHg2imGWO/eX0mtkLxiOIhxLjJmYeRQ
Yr0hNd130hH3dCDoTpQHIf1nuxQ0tAiui+Z12txdzPVLtrviQs3K+WLv6s3E
X5cWdS09AqglsxxQnirYqeHu+yViswE/bG3nQ+HIRhi2PNB9vTFioK/YId1V
8Hq1lCjYIHJ/ot3vjZcQ+jF6CoXqWRIbXLSn10FhXMqNA8g8GZ8p+auQDzZh
7pKaRH9kFPwK5LRABtK754bDhPJj5JhbqXpjDTwqfxyzs3IA405tDJHz5C+V
xuZlJgayval7BjlweGpwbdVHESkhglmglY/M+nJVenfdNU8S6LrPGhPMreew
T9/UCuKjqE6WBhEvYrIn53cU1S1VwLkjAjAMkcJco5Vg+gUOwDyO+O+RPYnp
paCB9aNOLEy+uvgp3id5xdX+GlI69/YnwOqXf3cSg9jSJxS0sd3LX11p/et7
LReMZIJj44B/P/JoeY0aH0qFtCtnRaYQBHvcThCy7p9i1lOuzMhNuZp3f2iV
m2tZJSG2MNNX9PpzCpUhz7waoC83Mio+RzGa/yKWY/9Eqs1HG6mNhDxEg0jn
6nISMVwMIppqf4i+INMCBExlS04PtFTBqGFSMoM8TTj67C53/fXiuV2u/I2G
6dAe2uW5rXH+3GWvc1hKvphbcQQBuRNNr//jlUmV6pb+o0Cqwixf5IcMP5zl
AJVmDfJvWEf3rKnKh+6FhR5FQj4woymoFxR220Cp7H9/GIjrCju1nk3/gy+b
beUWoafzJ2Gffm01jpVRLl/D6Dyxcm+GRajdCo4l8gl5KP++6UdHIMWnStQv
3vnSJZVSH2AKcTYItXmR1ogUQ7WtxSeJZSFLaiRwlkmK8TXSMEmySBaqskLf
6I1+zs+SQkbIZjj5KBndlUe2dZK4/1dn9JPmkBiqCDtb75vk1pKM0dihy1Lc
LADroXHOfAD8G2TkHwwdhfu06Jn026Vo1rJR6442Xoj8+m6+GWJfx7JTWYgM
aaN85lZpFnQFuRONuRQjytJY8blo9qOHeAxN+Dd33V90W9lDXbbhaY1W9IJd
pg5GUjQjGJnWP5FB6EKhDZ1kz76X3H3fowJFix2jvUu6/DRxwuQq+PIj20ik
rXiXPRqMZU4wRsYYQqiDXwy+BL3J61ClE1Fj/MxMaeEqtMwMVgxM6kRzEKBO
6oCydpTZQOqDblmscd/WAVjwxbD4X4HJh1ImCSdBzPpCIwmK6TKegKb9svgw
c7usDKeCTcTyVwSjX+NO8L+ckBF4uZoW8Wg0gyrveEG0xyLL8cbhXFwheRe6
dD40ruAJsh0IBodgKoXL+Z5QWVa3wUvlREAZiBBhfzDJncAjyyHfYaU9LADn
sO+Jq7BYdiXLMuGwqv5kNj8e9vZq3USbPVssYFIoRUsCAZ40A/wXsidLybqy
seP/UpShl905lCZ/aOe5hlhVSQkkTUHaj6Rszu/MoWZ0+PsfDl0LwmU0ujVj
HpohTWyZ30P8HODpugyjDAEKTOdtLT7Is3q+vttT8LrEFGPudAocp7i4nQBY
JABi6qv7+k9ezUjSmzPgb1QYMUbjtCi7uhAvfX05KSHPruX/hiH6WSiYMmv7
XCuukg+gZB5hdHqJ1PcXBKA6fux4yM0Q9u67LLkmIMb3SB6ysDpUS615RWKQ
r5yBhOzon/F2+XpWlN2LH5e72pVcfbPUXy8F9f6b9KVDqYe3Oqg9HOIxiGbQ
9UH41sGQ2ESpoT7hZclev4B7MbmD+SX6UZQTVQZM4gd/Q8l5GN/w6RqDBF41
k7BW3J34HeR9YbuKzCpgxRjodUS+cGd995kSbR6tRs1zcmGAvbLSig7Vso07
fNdU56QLxdKhama0p6E9kkOGY02FfcN9BLeAapXsKLidatFbsyaFWPFfQvA9
8xUOAAIwk3jyK2daAIP0LYHUQTyqV2tZNNrJNxb27z2WjLQmlHC5OCTuSLz2
L44Hn/ENQqAHqz/GI8QeED6FgjHsPMsVkpkaP1f6nyNCwwjy48NHmocc+XnL
hnmZm8VAI/XihE0Wc6tZOfsIAphzGeQLzZRbJYb2iNEioKPxoTqa5RZ/fq+I
kDZgu/7lGNGHeoo4Rm4dkhxrGv+xNqJbseBD7XgsNH87fKeIfmCp5tcVEcHY
5sUqnaGcM/77VYvto36AoywYqkEIaOcNzAuF2muWKfkQ6RWMpzfRxTkrgjwz
BWrUOfkxq5d+zYUdd76tjpZlJpCUfmMb8tRZJmfBvCK/Nzruxu9orxLubkXG
TpdnZ8+8TzvWMlRjHT70Vo9B5blUpMiN9i6s2j0MzimDGDrhZyS8KHHwwiWg
I01uk4A8tnmuqveXYHFKsaECAf4bXS0N5jqAU68kW1ZGa0pvUMM3hpU54qm8
4vSwnRpGYHwFoh0Cc1CNQ/URWZOPfJfi2bvYM8asSu4lze3SD6/aVCrYRQM7
ZADMPQ7kDhHwFyiPD1M8JxtL3XoVA2fIK/AKTQ/bXXAG9ArScD0vK3swU2lo
MA5/cStKXwQ8MFV429cN/trx8kzrXI/CwdraLRi3/2oaR39K2t648FeoY/Fv
+ax78HNmsNqVNrW9iakc1sc5w+LagZJNvFD1seP5QXmMpugfw4m8hSs/OXxK
oRQEqWr9h9VLgqF4TJNZQy46AziY+cC9ywge/bRAnCc7CuU1VpjCY+b6m3+X
63L1xTmq0lr8y9MyJwGuIWNPFne1zGKkqupAN3H1DRdHCMamj0wja2NfIait
r3vXxcvrnG1fZpfLX6W0WNAlTyMRQ6qmM6PtB1Pim+onYZ+VLwc/OpgAIG/7
KFsnHLO5cBMPTFWFhbyNzqEOcpTQfOYg1/mYwqa5HsAHRt8j9U0B8pNamAxB
8qkqaHA4y/9Fo0yeehNgvFpnw7DOEgsHw6zBQR8ZeotLVNYCvIP/WYpUPNfk
8mA8kvIMiLgJfZG/6HPZv8QrCWzPpxVkUMSo7SfQuipqBzC3tN3c9rGODhG5
cbSJcllAP3Upx0JBkOqCVe2LnniaJTK5TyATa9pELd4/Vptn3Gw9huZNV/MZ
Hp/HYm3f/aSQ1w2LZkdn5Pg7CYasIHhGSSQUHFxaFqgkRLAhrRVNzgksdZMj
pa/IUZhTYm3ROcX+6ZiocAwjmbtWLb9fOauaqTHxKjL6shr0HE43qCMKPl1g
JYMat/CMqPFYfE1tipce3d3p7z7xL1/Bk+zo2ws2PELeHSh9A6rXKhtcbU8g
+8KnLIGpB7Rg8vBA+Jiv14rH9PQCM6OIygRdKrEjy9ZiiVMD7IbqnVKwuW++
V/rNHgSN2fPFMMlS/kHDhvYtYctUcv+A+laHWDtDVBKQMZnckadzqIEg/plZ
ofrlGsxsujAq/mHF9DMIoUDuzZ2OQHym8shKae+OZ2Vfs5KvGw7F4AUp2rIT
9EsMF7XWtnRgdDig0ZS+IS6r88dzqz9RKuupHSBnOLDsAUebN1hKNbAwU5hg
gCt/ooi03kHE9qGU43T6XhBy6WA+c/Rmmk5daS8IvZqF+I8pfu2mGsghNaub
iQZoOhbCDoj2eGQbGqPz0f/nJ9e4UwbAgerzfZppnmPTF4QRLZg6QH6QoGfh
deNZuJ2KSBEUHVpVy/wucZVHl+grxXmh68PXaU/GrmZiVPKDW5ex2O2+VfM1
aVsdXf7OjwLJalBXH5Zcp41Y4BBCw/nsZYtOZGE9SZxyGAzv8I5HAvF7pCkG
GFvcAwB7olhz6MujTgBcPxO7mbzhzn0JHl/W0teTClLNHtJHhwr431NdPhl/
Zye4zv8tNNVsNqxV3yZYc+vEYeVUrEkdJFmt2xYez+yOruNPNXYz8XP5/NgJ
G4hdEpfm9kGPaAigSOKLO4if4yJSgVtzyYqZTeOr+hIMJZSJjgPMrSggxuca
PNeDTH8U9vSrTiJNCuLIk5METyAy6F+dxHe8D7fK+ymxOcnrQOCyId6AM5tc
q6yo+3Q0hzQOrDTF7YFYOAR6vWQ71FTZMBzXgUhl7SA4oIhZBfm1fwJEoWvc
oOHu0h07LjOgImblsMmYYT+uCwpAWM1Ymyr4ZcFIHj95ZyvX10Y5/ZcAWTsk
9VP8FRT2SVEruIkYWj1XffMiccnrrDkTQsKr6Yrq1+PIY5Y42DZHWE8T0QSk
xA1fA+LKayE3gh0QhH6KUcFgXgeih2lYBwpAiu7yeoxSTxfuT1McB6vPRd4s
2TI6GeJO+uUNZKPD1CkAClxbT+jrnBEeT68sHNLJevWG44dY9ujuU6c/C7YL
BRb0VjGY2rpw+ShAUVD+JBog/gnBc0C001ZJB3b2V5wUTdn41sW92EgVMT61
BuwvVBxQQCqezOMci5yrlbxAGB6tuoEx0IIvS2ojcSWTkrV2GlNgHHRr/+uJ
okqnqMf+HNJIig8CC77p7B5Q93VR3JI8IlMGyEMAXaSSH+leJWh4dx9nl7io
2z2wariNbnCXzJGpztXFTD4ZT4VR12yxzSzPAWzSO4WxGb4/0jUCfkRzmrJN
7mrk3VLaMv2mLixvOK9nRb9jC0bat45FST43cAHx3KmmN2gcQVfpVczWnEH8
C3LrrLQJ37zj8nrLFkbr5D7R3tf5pIDNaiZdsj+9hLjz2xekr1bm/s4cF3li
+0KhTCv2/Dknpz+vsE4wpA0AwBzgw2YQocrpAuxhwrYJxTzPeBfamWMuxei7
czLSrkk2Qd+3nWaZ/xR9BE2IkEt8pvfLIebMPgJDjBrBPvveoeAfVt9tBpo3
9kHaL2HVU2f9XAv/GBh6Xrcc73n6dO7oxADHmhS1EsyDK8h0Z2+67NSIqTtc
jzvgwUQyE5m3a9vF56G2mp44DZ/bv8pL+PI/QBgDI2Q+VqnctZjWXo51oOSV
qRdFO1Zt6m5vSaSeQlEjaw4vmHf56lwr2qv4EB2EMcd3a1Qk5DnbgQce9iIu
8OvyEllrd4R6dpjcD5ktQirq5l6bD4W5Rgr4/jflb0BRXrh4fDLm1W69ta+y
eWHiqezUwH+UM1aiipfkt5yl5TAUS8hwlcNEOr2oPx2vE7594XPXket+hzYT
SGwED2jzc245sMvVZr1sSgrvZy53i5WlxM6t8OjmDGlnmJBZkr0yAMtV/xmD
nKxdiF/qnzGQ7gjOuPs4uD8askXLURGvHO6zsWJSPDrwkTr66/8tog+KvAbG
esqJ1eyyZvIpz7eQlynkAqe2fHt4xMOOgVkjb/SIVx5gAUQHkxNxCzECbna1
FW2c+vWdBOrw6ncQCirUIJTqskSjhG5UGQDRggX5VxyX0BcOwKSTiosjKoxx
70gEA4QL+CL68qIhDXcOZS+sfIfTOuoG0s/SbBNFqoikJv3zR2cH7X+RcCAV
5x2stnomyvxbOKyaWJxV53FjajIWkjZaHVis0mOljksjORXwiLP81ohKHPBe
D2Ja/16ifpHTcv6sgtCBWXiEfrojDtLZy5EwAFAtof18LpVBAWt+NcvbJWM0
PbKU6unqOvsbqT+FllEjlm50naofKrx647YT5AfeptYCWFhXu/rKJg5b/NAv
cSArp+Jy0DNXHh/Rw4YaKlyYWCKqfKnWhb0MpRgzIwrrRfWC5UoFqtCk0SDx
RtWV3vz7+yHhcvEAMBBT3JwdJChYEEic5nCvicVqh1+wLcalzI5lbhxch7IO
zzOYG5PIIuTKNe9lZW9yQBV1IU7NorTddsIBE4JxEQ83MsbYaGUI2zPSO7jh
zbp/e0Jz5LfHpacu76WqqSUa5UdjbsbOMgw7+eI8Oxx4aLHlDmvwEVmV9iLf
tjLlsWrHckZ+WAnnOkh6N2hf/CaO5eeunhpiOGNE5Sc/jmSIxXaPRmA13Jpk
Zrm0Ehkk+bWYONa0pdLSqJJY5DKrYNQwG9qHdN3kaZMcJpZ3GqiWDnSXis5X
3YiPwaU+WEoH9KkLe8/0M7sHf1bL3mRxugWU8RBzA3N60BxfnNqMvtU1RzUe
h8D0IEJAAsrGeQVlpVXYo5IHnBEdjdV3ib5KZ69mVqlGrnDCllqxMB1Ed9kw
6gsVyXO8VKzb+8CrG5Ptode3/UBo4YUxUVJv4r6go6BdtUy2vu6VxMKE6dHC
wQcsoUaVWMmQd3KFRC+/8h4sX/t8vZCX0zV2SMd93fMK6SuopubV05yE7zov
ZN4vMsuasNY46U5DH4ifS5l6w53T1tbL5BuklX7VT9741p8eLZ0I1fXD0f1M
g56RMlKv1VQHMtEKP86t5dk2TB0Xiq0PIHPspI4e8pq/anyZOV4Rod6opFyE
5Rc3QN/lIfg7AuxHxxoXcNkEqpcwRc2y2aJms69XQu1/A45d+z5gZpdtHCVH
IODU5uPWYlUncEjiacv9nl8+u7r87yY/BjsOb7ePBDOyS4kNDN/B0+MJEAS2
8WZEufnYuGya8wX+Venu0LAb/qfolWAPo2ZwkDaPbOEKoc8NQ8HCFEwj4UC7
rgGkT9viiUjGzlRHjgH4515OaM24cv3xrWGtaePASasQ4axTT9wnCSZqPFod
yEi66Bht/ibq2SeHHElskUy4dOVf+VadT4oZAl8C7nPwMIq51oQSDJNQw2h+
SNVL99LhIJzZr0Fv7/SbtZO0x0qsRyE+yPQQ3shurp+h5uRwJ+TJRxosJqgd
01ZvPFU6q4ljbdXD1miW51601RBnLARMt+VU8yGWjQUHMEW4Q6d0VHpOU0Cm
39xXi+qdpC0Es3L05cKDBIkdILKFljo091nYTLVh9U/LIyDhumDm3hvpEee1
w6ZQ6wDwLk/OvAsaIQefaK2K6YigGrLVUGqQwrjxXanWBQIKuXwP2n7OaiZM
/wuTZrZWxkKFrSDa+uZhmb4sUHddnGvQZg3c8oXw/AGtlP53bImCygpf7RYz
vK2KvIl0eOr1PJ1CHO8lyoXG6CYfYlHpkEHXaNEfbFAJxdr6BMyswqpQy0h3
qzfYiCUm8S9W7z5zCVzn4u+lgSHcGKC0PAfdKC1OQ5feLMP/NG3qIpa+k0Uu
UIQLyj0Eotej7SqbdW5j7HxTvNRtIbWHw9Q0VDmWAoNZfT3pSQr8R3XzpQ3k
0uRl6RmiQu+SrTAq/EdNxzdprmZlF32pBu1IYVJxc3/qbyhwDcc4+6hkRewN
QGKj37cJrkjjuWlvEBOfGUhQ6rtAelZJBWVGSf5Idpl2LVe6RJEusxL18iUx
S+K+GaQTzNpxdOsrU0N2uGMQY5jmQwk8aXDIhDuu9Y4YMKApDvj1tirzY5uc
Xj9f46GUz2L9rWHC9H2PNyLZEW5NCpoxqctwZppCCnrQTe2jsbgfiCdK1VSv
hnBuBPmEYOPxmFjopeWtjpNiBEZd5QxSdJreNWzC1g/EocexXuPU9XHU4yFt
sjXjVU8Wz/KOSYRRpMylN41M4j414Cm9wHXIe4a8xvbPNeSosAabTUrRgv7J
f9v5mqFFBF0GfNKKNM0cXFgoxTej2lX0OH0ngHOXWTr45YN23I3qeB2QuwrC
Z59tcrb4oSabf8mdf3SL9UxfFwblMuuPqm5evDuCoQEjQEUHc3eD5dyAs7JR
dCvFoKlowoCeVqeYUBz+1a1wWSSth9kXu5qMlqZM36M/w3TUZZXSszjmtQsl
1KJneyLNK2T6uBSvrbpndgwZ+2suCDmXlP4n0kjUTqoorfStNceRDa5Iiu6m
F0wXJEEYwHliRVJ3opaSqWGvMypsgwO1Y0spmkX8jEfgJa/cL06FuBXAWe9n
DEVCfGo6Z2WeaKORXKiw8QWT7Qfw2f3SbqUFJo+PVQ4JVD19mUtKIarnloCF
fAnN9Ib7QIwlNfCjXJSBaz67Q50FmNluRlbHgtdMnodGaC5sczNwMjXnRcA3
BuE9k0Y2OsZF7jQ2iIdlLChKK+TUIC/XxtWn9/tBR5w9b62iMBOvy4pb/IB1
m7h8lPEI3UEH+YNTTttVxkImqRRUxzUIAEX0GK9BbHa8Ze1U3GgjKSKLNgcP
owyseE/xyk2t40rOZzCiVFFf3Mgy6KzRHwc3KiFNDhmkTZg/Aa3+WKMzq0dS
9sELjqGh1h2f56nXDwqABSXwu+LoI2tMDc2S7AguI4/ODUN6+PoCu5FY8qbY
twl95FLK4RAVGZdWWiUDS9drfIjvGLWQF9uqGSjC4xN4uk9/WCX8/LGl5evg
7qQBrkusJsGfcvgzymkgeDw1kQWMtMWs/VZnNjlFWXxOIQ/jaNXqpsgWVSVs
4ni0I2x4pYD/e7lxUGvVlfO7N+EUm6SEtys3yyJLVilrpGIFTAaQcwvovllJ
WfxLaAGl6gLT7loTx2CXSedcwAmPk4Lo7LGYphts3w0Sn5TJKYXpp5oG/Qmw
bO8+4mQyeqgWd5t/2wCRxz6rASvPTTcbHxSC9jdoE3G97zYevknLuVzrcSH+
Jv7H0WIrgHE2NsBreFZSELsN6Afdj51c1o8svM7uVRbk8CwZTB8LottXT0Y5
RdKHY1h6ZnVXfo/FoPXy67vkc3b5bB7C8jmsuN2KX4a1+HeWWC+KQwDVQ0PF
ERA9+XZdhLwmUPFZjowkn8gLrY8bvUGhAZdoNlkrIsemM8BkIXAO+WLr3vz0
6RFnE2qHZaR2q/3sLGZKA2A5rg0kmi5RMargik3fIq5NNfY3M8yRMKhANlni
kuDS6+RCCyqdFUVFldADDI1EiN3yKbB+Kh4gBXL1VuDNncztCJitp93Tkes9
ULeSOhfuDlGVP0iY8W5aFtSp/L9YH3UCfPH2V/oeiBDkfYKBSTgXCJnWhSZ7
BEDSj8qR4aFpMnXYFfHrMEvM6tgICakozZ+LoWVYzvLYbb2Myiqc2JWXpp1a
fQwx8qcgPUfxo3C4otLIkTslvfX7oArDFL98/3E9u6fi/f2bWCVrrALb8gvF
deJvt4SUSS4QD9NhSsPFX1jDmWD5UbJXNs4ZzqVgeih8AR0069rCDfjvoWeT
/hOZg2HucA/Kn8/G34EBPgbnj2+/BOXa2wlT0+4ONMEPHftjyVwp/gBQKhU+
zZYFwRlW1irbjtdsdvf8OFJj6+TK7MVUvABIoAnzKq9ZGfn5AmcuEMzYtNIm
Z2+8zEw2gTFohsrjLSGq96AfDJ4C0xhFCI/oEl6Ag3SgIH6v4TPZGfWXq31R
gBLES+6wFHTxb7dU5zZHl2uoBU81C/Qn233boCRw9qWEDkyxHwuKGNd8K2+V
utrYwt6BID0OqlKd1gWDRUyQeAbGDaf3JwsTQsZXMQJj24kmQ3syGFUJM1jB
HZY9d3lMdy7PfPY9/ccxwfnKcy7KjI6pveOvIegH7kifv9eSXk4/aR/4WXHd
zL3B5c2gJQGqQk3Qy+MgSg6eLBVr6T5QMHIEojxs+KlzIYHC3mBqkLVCMYUN
RvTQvLOziQrIznk6OyY1S17bVSq8TI1+WomfkfrFC+SeuR5Z6ApKMxocr6hg
7YvB3XJZzMRQLJPD1qIx2BvY6ASvsOAyF/MMLQvpQ6BSFWMeI2rJF+2exfKB
MYDD1agba7ru4n5zIcB1joC6PoID9ZOYWvaVHnnfqyWW6SuaWz9Lg1qIWdPo
TAP+CpbY+W2SRgw3vwGNbnv+aGVmzWOzABKtT31NHgkMBYS57fHwEFG9PLI/
mmIswsk8DWQ95uLVOClxgzRPpN+b+x88TQDdrhqv+RsT7hOJj9Bt7eKtnr5g
zXSurI4I5uzno3I8aMvAyCNWPiUPnArUXvGkgca8EKVs0Yo5aWGN14fubwGp
12ZZTsVa5Yiatn+p/jel6rBB9gB3Sas1PwsxwSQnNI3j57Yz6YKxf5rXYng4
eXePQsnGQhGOD45Ags4KjFzbdEvwqM0KWbbqAhldRhNHr0KPDBTE5ipqOUBj
3b5pbz/sMSvrJi5u3+JrA9HSDvrWtvkgc9gsByAswMov+z29CFp722IMciRN
q3PAM7yx6HjWixMPlpG1t3uwJdJC2pURuCqybMcB5SNv4EBfkvuhiaa/QTCG
Zk38nOx28hB/3is2XOlCGVVhgvVNLyGWftiQV8j40z8zVUtu2yIep5hIfPoD
uanFlW9LnUDKuJZbRBudqHCvbM+eT8PIgwMDcovAFYNOapgztH86jV0tNSrG
T7ihlQsZzVsDMt+rs1r8CBeyTroVx2cTPvf6RJc5HsXo6cjNSAglwBV/2ujS
ssLmVZiswzp6BvXKTlzF3PLKyJtM9JpeHQFMJe7Ul5KP2bN1QcLS+SQqV1NQ
XsyPBcYNpgQf7oI/N4Xq8Mw4m/JZ2XeekiGWtWalHp51adJ0xQXm6rlwyAo4
+fHSEqaon3473aJKrq921kJJgHTf/oAzVKuWuJskhE0ietih159VQ4+G3QMR
2Zsv/tMVgEosCe2Du4r98PACk5v2jAoEGdxxGYe2gR9FTPU+eccL3ZSFa0e0
3w3+DDBfvSNrpU7MjWCDcx+XNEZCEbl+IS6dEVvt9Fp4FexO3eafCfrzBRZF
L5yFrmA1dABP9vDgP+xg9aZvhg59TMr7msnPwhK/hjQa4JDuNnWEAyjXHmA9
Xg3A3Z6ndLOnbSA2LU1/LLUdNTDFzNGTiUB28PAGDm/PFrs/Lx6J1HswXSuR
vjhKrB763DF4OTCzcvdxgwzJrWtNEi4iru7eSCXqsH76r3KtIOcwFDpjXRhF
Is18cGJdEd6CYFCYLJ2eKReB/E7dmkpnqOF/Nc22xCgvf1h/G9d9j3q0vpHR
UH7Fdpa7mSC31lHaNSM8qtTgiUJagtu9XGYLYAymSp6Qk6Lsv44HDKI4r6B9
tL2IajUiwdZNt9YtHDBsv61BWPUM+JFumn77CRcTogVmP++JEsP8VjXbAwx5
UjSs5tfuERNI/K3LPMxQLaVihWaUm0ckC6HtLhtJaAbodFOTgM4DoHiZCRKw
wsossbXvuuWCtfnzXLbZD9IbPs1S5Txt+ZrItvulGsv1N/NaKC7EfdGDwWvw
vymh8r32dSdo6sUsqvERhtzJw9+LBSOA41QtAjBVGFNlKsVmUlFGvFhtoS5F
w+CiXypSQq6jT7icuTKZZd5M263tHwA/zw2CmaZi0MOGOtInCUnz8ox/8ber
+zSR4wptugBwOqFAXFgMNMIjceB/RWywh+sSLkxQNn5qkp/13A5iWANCljli
Exi45DuFixKGkuZcFxjt9CrHWzdfuOqYXXshwBzUiXR4Rqwmp1qUKBOaL0sX
HBTVLYrrnru39vCthBhPFCeGFQr1LufcD0d4vjzQFmM/Om6RmdsGxi/0L6TA
zelZKHwdvmp7UlYbhSVd6V80KT+x3yY3OKbufOXeuwrkXTU843PdSEIg6Vq1
ZNMsb6gKVJYdRNNSaTeo7665z+n+nA1RUb3ZKmzBGn6Pn9CBXnzfA/WABiap
zLGH3Ae8B03l1F4oKp+/BgCJbv5nrzlPk2QTtQVGOfh1sxkein3OoCZ93IhR
/A78lWTCnLZy1GlEhh9Sp3HyeHrFFcSlnhCmtiKhW+qivrm0Ak6xzjM8EQgC
EemTDTM2VUE5LK3PLa8RzL0uK6HJuIaUvsJ4mAufB7yHV6/Y1X9mklIUoYNZ
8Mn/eAoSvHlJl54PlUSydSywhBay2aWjIjLC+7UaG/uUIfOI5fexiiJ+lUiF
ekaeaaxfq5ZbSAbP8y9qsq9HY2iCZ1DSQxUdMSUSUGeKNGqpD83y8O6CylaE
tdyN2RxzdzHslN/8/frne7fJcg3I1iKCQHx/tmpiGPWiCvmtMRpu+2gydt4T
3NGALNIkA7haASwIXgMNyL35o5UV2G37xOCmZFoeGuGOThQAWvmrzuNIj51h
iC5Fe48pyTiRgSz5vwJe6WoBFgI8fbylSlQlW4nT+DUR92fdvK4lxjmX2tcw
z6Cbw3bUoofO9PHe39LzLRJJPtmLw7X5dm89HlAqce6TvoD028uztno1j1jJ
gm7VeMjZ3B5D7RQAeecwOeKu9O1+vJDzXOe5qp97sBFa+UxeAIaYvArwkyy0
T5nX7q5A03Jz8pLhQ/Ft9HbsJVhFcd+p3K/ZHyNuDSWIeyfAFT7DQyb1Ty4Y
xz0q41Me/fJPIhkS9p/pGe1GA0iHlYuYv9HOxy66cPbfvri+JvVI6Chl5MMd
C51IECW53drLxU/Yf+A/UM5N8dtNcDXKmbbfceW0UJFQ+tGezNxo+MjTLQTv
ITjl1i4PJUK9DyZN9dr41w4/bAIZxSsG5IY6e0PUeV3IrfKUQwJl9bXTk1aV
YJxGuXsv64Y6mfGbSNLycfwVe2RqGCfkUfGfbR1c19PggSlMitEDtSKzN4nn
l3GlP9N1xu/zEipAZRd/90nRjdupSO9Jv7x1aSyAwPYCMXMJmzsjq6a7yFNd
EO40C4JGGRUKr/w/NZC6VBAGNzv/YZ+AA2aJIl6v8pE+4WxlC7F4CfSb3ibV
NrHYUIRmBCIxquNqAU4bfJf4gGq1pjaPFUKauZjicot13psUyi2XGZqtfHrk
YD0nEcNfdgMyZrPLW4liWruRSyFNXeEF6ONdC+5ZDjyp7Ag357V+icHy8+VI
FI5WfVHsEHYlbGgbrsB+tHkLWdvWmuADRJK9aluHJdRZ+/8OcOK7vbU0I7RO
sHUlDygwm9Vh88eFygCV5Xa5Gvdu7q5MbtS/NIotcceGskfr7QhN4X8uuWS/
I5E5eNOJXzDQCJ0DDEHnewuJG80qSJDsGP6oTpuy2kuSIRpDFGN+xOeG0t/K
X8gLRYJGMTvdpiGD2remxHaZjYu91K0VuikKn4GfIGqmwIPc64Nsj3IpTaMC
So8VQoGLmFavroFaMH20uYu6YbyR6Ol8qWxW/P7QX9vLnOc0p7x7sEzSjr0i
ixEq0KWQFmjG4jIjVQ5Sv2x4+lGj4+MPSZGlOoYwbqVqT1GU6/QYo06DYJMB
HHlEeJJWzc9TjKTXEQza5sX//s4MWDfiJszDKyPqQDWRZki65VyLNdOh9FzB
VlRGvXykXYmgVqqkAT3NpgcY1GoGt7y0j8N15RQVjdc2jSKEQmbD0gUGdXSa
FGEv3ZYi6hWNfkdyhJy339kSeg9QE5GmYcULScNGWkKxFTL7ZW62/5KNOcwQ
WAkTO8i6aBtw1oFIQa00lptAFrpz4+X0dPN922Hs1auBQYqPl7SIbAYBb7cs
YUPm9hgb+Ai00W4NtZCmg0ZtRVg0KrkigmJDs7ahYNgwVrKhI0KZg9hb9y0m
b6CjTxShBpGpspEXmVayRaczMK/IzM6/sOxAZzRSQiStsUroFP38zxOaAklM
H12qEJ7UNnZeYB33ObrQX39xFOBSgCFahE1ppKJquU9/UWyEABpPnlMyAgWU
6sNO75AS5mOVFK6StsJbq1HUCk4Op58rh7UJOuo24kxTw1ai75SwoBBgkuRT
mk6A2WVQRWpw+KhBAjNPyducmnz8RiNLhPzQ71m+RKK/uobfodajobM1Uzi1
Us6OIcrkZu1FYgxERDXFPXHotqkxS/58WC5fcNHjqNhfXdO5KfI2Y/v95xjK
JlcXMQH6gD4LCe8Y/4Q/ius7/aC9lFlqJ2DWXQ2I1e76+yEy8h4TriFExdYW
ZypuSx+dxnZUEOlq6+BzM0gdUIMN5KvaNqhNGYWbYbk8oKrZjJW3CD1P0w06
0kROX1dvZgvs7tueSmb7QI5Z57RFIkP8Dx+V16hpBQAjmlnv5o1Dfr6VatjQ
HWDmmDMdru8xPbMRIrJ92tpVwqJgJp7bnZdBKPM6gaWxPh/WAK7s2pVZlHLT
clXFClKQhow24A8ifG+YvArJpcglZGgEVlFoBdlEGzjpiV4++TJlPw0dDCoa
c69e6V9howRvsepwxlrAYaKmg4HmN1PKYRt70o8X2Y0YYkVi8EaJ+BuNF/mG
01NIoc+MnquocGmURpttAXVbBrrcW3Aa4crcVyOm5or46YHhhz7DV5yN+S8F
L9o0CB5fYPgvA2kf7VfvfrCaFuwPT9an4tgPCD9ripmxrRHsfE0hZL8HNh1G
eo2WuGl3Ex713aDV98iLNd2qk4+6rTy7NQLDgbHbGA41DBzsK2hiudsNdb9N
gjvixmD7kKzCZMtFscYedn6JIpg9LRVMp0TmlrypUR/v3NdqAHVP5vI6b38X
qdcOEDQ+dPA8eg7iW1K1hBJ9rx9YTK9/cgXtjOBh9Cxq6hEKR7HF/cA/YfO5
39Ha4/S8PhbrhrC3h8932+ammGsrD/75NpuG3J2nMbSGMGsko3WvrwEQEp30
rDObM0OxsfTLnbI6ZFn1oc9m0XUUGQkJ2BJHifrtbo6RL58HbsnsoUbvTMlT
wyyFBvgk9yWbPRV+fW3F1iw6Yo72HzyZ8I9J0qVDO25FN5nS5s4i1002LyyS
TabhiLM6D0ctCrm5BWJEJzLT/dbEmnRoRa5n6iQn96shwbW1yjvqF/02bO8e
U47GHIo84ydJTC5vzjv0VLfzixpjql9Y3Fb1BTc4ES6/j2VLGUpDeiaErtSB
NFkx9Fx2lOtzLwNcIt5UljCkuDdrp2Mdh1veaTQph3j/SIKyOBj6rt1idcHf
TM/XPFInfwsT+uItUt6bNSWInYhhgOmL1lY7zMaN8rGhtV7bM0HcSuBnN5A8
w5tg53p4frWDsuSuAblcMfauk/4lwlVBWcxY4dZymgpKg6wanpBrfaKLGqRI
2M7NWzD8cGtMBh6pU7cGviLnZPVz0iqvu6Zt9rIcbHkWGgU4yAK4uKmwSX+a
5uaudXQFi+7CrfxkACtzMElr+Pf0vo0ypRhuaQinRpd6PFhe5hs79Hl1ypaw
LRH6pUJD8a+sIhX7l28NfxUQ+U0WzbIzTL1WzT04KOCogl6/D+N6jKlW8hQC
7EsbHwTGp3eu0phkkRYQr3VW+gdtKt1bqo9waRGHFpMF5ZWPcyHh0cJAjjmN
tqEeCdCmMkU+MgkTph5gGSwRUfAnB3jcpNlMY/gRkJUP7nFL4bCiE/3DwfRL
o25bqQltl2bwe/XSbXg9rAEDjwPhtbps9W3HuHkeNWjX6FbeazU6D0a2rBWy
k/kyMqor1SJqdP/9aAzCe/RwX8l4P8/gxgaqSGNemn1Nxq7fuE4PMQWrNYp6
q6UYfOuwL89lfzaAp+02lqwJ0qE7UXsJfxOuYNcXFDJrYk882mZqPap82V/w
mbZ3FB2ou10TkhyMCrjdZH9zYZEbUQgOSmit7j0NAssRmohkmAYx9NJlEcj3
4CVmVEWi9E44YdZGlr9LUdlWA6xJe1Xy2nJNK1TbUyCx/+J3JumPh44ktGHD
dN6SJUrSNfbF6A3NEd0O6mM5KLcrQvAYdDA031sjwrnu/qm79Gv5yj6a4Cmp
ZOEzVtAT/P9Rbw9T9/H3LK1UaBYB4e5GzVsDYdKiV5iHnOjOlQ7189x/EPMU
9wxgfFX1XVXpzWk8gcdbZmg13TSyIzav0lLYflQesZi8N6PG7UZVfVDNIz2G
eN+JMnxNMDnh3VXlnK6CintTG1eEjQea811JK5/pC8RwblSapSCuT0wwJrEF
NBt60h/g1XDj1xlI0nQ3uCAiCLhAMQpDqY7lw0PAS4Lf8EYqthsHE8E//FKb
+J/DB6FGEuuIQCZJ/1K+GQetCbC45CdLxFs8q6Cngmb0L9u6rA8KsJf1r+J9
7ntDdKLQRnRokqjog4SvK7+wzsX/j8Ji7daEHUqt5a0gsDlnn/FnIXvThNYv
9i2SBbzlwQGtf2WNdzyQ8kyEsJ2o6L1mkVlXQjhv90vlJGyUFLyemXNlWTSp
1qHM/gYzxhEprmO58CCd1SeMhthPoSFekshNxqbC9LIuOXh5JxVkwuxYtRyk
u1jyn9hZLmJ4sMQ1SftadST2MgGChAUuIBiWdm/aDD5N8pEPXv1D6SzgF50V
BnbjtuLBnXxql8d9b5yvsQ889Wj2jY0PxqU3skVvHpkE7pDTbQg++f+QTXEA
d0BKvOQ38VT5TBvN8ti0rSGHuKZht/2NjfQveD2ppnEIzvPQ0YcRxcyZySzP
RDOiLmfjE12NOZSHbmX4VCiuOrRLe9bWiOkyeO3QOc6hL0iTpmBQMopJENA/
iPHVpLrvwD1ATbu7D+qqZaexTYUeaip9Hl0XnY7yvQLsW2T5AIzjktGnDSRt
EID5q+e4du6hQFCV+QnYaI13h5YzGxkzp/7TFcPC0WuxSC+QUZWifsWAZ6HV
akY7Nhwe2Sho/hIaFM5xGLpY+rNEd/xpRYaSLZpLOIBqreWj1GOGNjcY7la0
uf0TLjypTxrFWlwQUD61M1VmLsh4rdcujvmFqib3jM1rmLLEzyoXwDV9WrUC
7nV2uRMSWxrK8rRr1uoKeuNklWXwa6/Nt5HHukAnZYF+BmnHHpH0iURp86cB
7Z5G556G9NT9hK9u6PazqEgnFEnhlpyGqfKhX2pHzbPOdppu/2lssNJa263F
lH1RLhl5PVcx4P1bMPaC8GgaVF8bvuvrfKqwU40Tau7N9Nd2bw6eOXxHk4Cr
HbpPqUTa+OFDA6Ik8VmOqr4HfD33SlZtTK+yCIcfamM9uIiHOh82wFZ1MA2O
xG1RpJS2iFKvVJFldZYTbTFARDRA8S5Ouaypa3WXTapsP2G9+sUwNN8dAaOp
wU3Z8hku38YcmR6mIYU8CbG7MPEVm0xZooWb0x0v2+oeKdWwgjGxj1JkUIxM
Ku+sleOf9imWlxbWGYx+1VIcMNT4EaHjJl4HIe/XmQxqQwo8IhBsV8Dp36h+
XkH465ZItICerkb/P7F2YsgaEjDKtW1BZQ2gjgPETphHa3vsWyqU0tqUQIfb
sc7fgZLfWfDUdRFJjYnHQttksnd74Y9El8LvuhSLicCPosd+kZcEIZpMpyNr
WLFuiUGnctub1cz4tpwIHz4wfWWy4J6ii+7l9wSaEavzlz+9xXB61sWCw/Cg
5mNNyqDHo6b2DVAsVA1cxaR2NBeQASdCNCZ7rQLJuZrweeUhAp4FUyJbwB94
vZHQx6kTRiOrecv1n8+KzY/KnVho/uioDylVsQfW4pu22azLNYDZNxsaaJz/
jkK0BsQgxrkyH3Ahccvwd424snFymeZCGtOF3Oa/kCbganhX5AtoBIAgfP01
L3wO/e6B/rLdue+GfHr3BEcm69SpZajHGfejZkoAdQtgQa9XJlTrV11/a1rJ
WTrTve2lRiUYl1BJTut81dudCEMP4jJrOely7JkOpBb43fj/C3jaGCRWi+zq
wMM+ZHEUJUmkYgd4yY8VGAFgMTABWZRtCCcPvbyyDipquff2XjfL+EGfOKNh
wKW91RH1FvJbGu9GOmx8D7ZWiQ7Wod1mLSf33TCVLA7DockR/FPb82mPOSC0
piPx87SpFsaxgWZy+zN64+VmDdeQCw8ytvnYW5yop4a4W0YpylxKhEYGaChW
BBBRQbHClvuAYf/zAeO6c4GIko5cuYxUoiDwes1YTTrWt4gaF0KqZOY16Nm0
SDm1xVYlDiS5jsStmL4/ndfudUk8nHhc+9oZ4Kk81Z9Hh9S0eOjmCsddeogU
8lZcp0ipfK69/6AS9r0hMUII4gGRBqDI3HZTN7Oc9yBDbWtovxUY6FDDOb4L
VbokG3UdfCR83qE7Y5WIwhpwsvkqwi0GnA4jjYBbDanvmOlt/6xFGczXIPwG
EYtRPew2G5UXGfdFB6sQSvWx1XLjdPTBnKhqSh6QClGkASzS02d4eTHwRRBZ
l3lWQCarR967hiiRjSytvuW5NJVso0Whx5h1CnWVOEAwd31fvtWQ0SN7QHjQ
dz42VWTei5uTDcuZvn/q5OeS6uActOFCx39CsuP7HntoAZ5k30O+u5qzMiSU
5fgut+oR2imtL4UtqH4spFPi1jEEUm+5u581CLDgDNdK8C/TnFEpMl3kZohk
/r03yYHlnMvuEv5EwYxxHAmrDcFRIeImSsmpIL5GK89DL7ZhWZj0yP13YN2u
5XFhUZDXHqLSbYXLF2d45CyFlzHE29f+5Zy7JErhA6EJMveixpqOU9elShr1
bdmvW4Q/LrdeuSanCuYef6MpEELilxNaMrNrPDXPV2iZRjzm6FiuDafAJ59C
Ars+4WoWKl6vsq4ntCvSLrJ3rlG/aGtJ9QAs4NhcFgLkF9uOLml9JGKKiBe+
hsOR7EYxklCPVk2MS/7IiW5QjhJCPcGMZhbBBoJOjGqSk7C1QUSb9K5+TzBC
kMQIHbFKVs95b3/2ACcWp6Cfk8+yReY2NArfpK5OESlJsavFFh9LNCGARguX
ZwC0owOd9GHUd9Oc+9JmJqFzKjNEuV2vHRk7G+Sxb7Rv78PCvUx1VFxSBfkV
5dWmrm2CksDvUq3+RZSl7fYVrHwCNF6FKcT3jD0wFD8YeKmjqDyrYxEWVe/6
ImmITkZN51Jh0WBkixKYeXgDLDut+6gZTxr0hRy8hn1u/JLHSqyO+nv1uAFq
wT6FwcwpwJZK/wwFSsRXVLn253v47Jq2+pvaV5mHUmcvy9rCT5d+iyuoyy/N
qQQgSTf1Wjja+Scbm9Y7fF04XJsNGQ08A4yjOFw6mesTfEfzTwRIzgdXsvEZ
Y9foDkH5R4tFL9XAJagK6hL0vQ3Exedn5YFu5pwNgaRk990lYHi3ophRgx6k
WrvDPgTQ2wzgkiwoDI0ppv1MP3iCjehKJ+0Ld396tqQbxR23nKFWQuR9AwkH
qBqB4gt5pn3odedfDe2IvG/ArJZGudb3kPoJOjV2byZbHNbbEMohl6GBL+c4
c5Nw8NwEpVgF7eL8XPHNuW+NkHLhpFbu+P4dy2Oiqzwt5mSQGqVxevPYTc7K
wKjI3U9dEimh0jJ2uYaVvTSbhZ8o+4qZzsDWeHzDLxvZ21R+BvAfd5IbC3dw
p/DvzxSnwyeqrCQCipzWcbcsxeyJO2JcPWftn19lgXGryh6ltEyeJmtnwLav
iPCNxuqfwJV4Fc18zCZRBFD6z9e09rSUqE8u2KQaKCPXskJrL2v/Uniiz3b+
sBWQeJowOWO0faUaH6GLbIrMKNVbzuM4E9dQbjQojl2RqtcHM9+w2vxiFDmz
aYPgQOpWSnVuSpUQrWBifd2YAU3cv8e9V3zkj8aK6/xTDR0bSdPN9gzY8tEY
4FbU6WmYBMfu3RaQv2J9Q+le1kwHQIgueVz1V8FgAfPDAsqqYW5yQ6G4wofM
RmgJtK1iL5ycEUmzFyUzregSs3gCcQy8gyTAqus4/iawUqhtDZQo8JZQ8oKv
FEGDaYmM7ipcxB/+jly1hqz5UnzQlDlTORCgXXfuydqopWMJRVW21VaK55zM
mZ7EhMof/KJteY7mj6By1UdArst3Zn35fQh+8xaK6nvU/QjKQj8T8N9PDyOk
hRil/zhKdKTY+Gdv9Zg2zu6oxDm0mA4ixKv+2RMOXnIjReLRmTmJA3Uun7PY
U/KjT69Y6fFp0exjDB0GyvUhtkl7SN/E+2GTJElZuJw49TIjVG22hLsLjIp6
3XNwokg2aSz8e9AmFO1Dur7fK8xTcxsCUIrn6twIzuMljg83ayZ3M6iJVVk+
iLc1OjrO3hXViok/GnVyKAniB83U/U1+Vt0FsZdYzDsrVG0CGshtkHlJJHK/
rNZFStsGYRGlsX4H15iOc8izwb0AmEAVIQxHb6uo14aD1kWOdOSdj4KvwDeM
HR7cMFJ7e1K6rIj57YiPh6C2pzawocPI/xCnYaYh56nOKv/Leusz3WEj36sz
4gozNxH2AKrgmnXMI4Jiwb7i7cuzX+LaPvPXj752z9tPrp6Mubeu4X7Rxuax
VoR1ugpbmn6xdasnOFlr0nWVfUzVVipdWTXNvgX1dsI0O9cub2qaFfWSrHxm
GNfcfJMX88KK7q7IPy7cNTOb90S2bJisCYit7GkfyOirUz9f9lijMuyIiVBN
bGhrlCyhC6o8b5ibXM3w98VOv940xkfcnawEmJRhsq3U9QFz19ucnAukN+sx
yde/tRpxCpGqeMrpAd6C4NQcWVLComhEifTfsFUz090WzUjnh3ISbabhGwHU
HmKmNJdkrw8uvjbbMS8w5ghvTXF3JdeCbJKU3JNBqkYvflFEYhd8hweZ/4XE
Qm/McCHMaI5FMcMDRR4YEil4bplV7gcSZIINZHO5ChfHRbb2PNPIFmFF/pI9
Hf3BRgUGkLvFB5L9bhJ48qUYWgBkp7LbRHLi5t7yrJLm2cg+Rn/IyjjrLzBg
ZMhRebUzdBTDRHafsL+ZRunjVirNoKZ2LpBUChycUNykOkNpwCoEzNKATQ/1
mpKnFcFZos/DfgKwx2yH3ABvHQsBUWITbS7BzhR52E+VmtRgJKiuAWWAYO41
XkW1y3OmnZYCpQgdz0fo+HQ3UmfyKYeTJMtw0p+2WAq2Uv7SRtqjhBdP6bZY
7mZPW0CBDaMi5D4GQkI6mVDAg+NHhj/RgJJjkBSCQncLHJHqIKb62XI2AHCD
9+rdUthk6SiLK+pDDD4a48nKwooGYjIXwhb53RAPlJGsWF4S4xBK4jvCcm75
B/pTwI/C1+otA4DANlmY909h1Z3nm42dur6nOY4sbwGR9WA9Z7/poApR48KZ
fCqlNXDaLnv8MBFY+u7A60PLhG2eh2J1AyJCgOxqhMMBCpsjW1hQ3UO1v0Ch
pR7FDvHlPL+jsEvcZnEyFVTkNC/LYpdJzacyuEpzYCL/8VaNa4ImnL98BQ/3
M4Ht3QOXfnd9/l6i477fImb8Gm3xWigz9EDVZc+vm3xv3j5MdXcPRQj75UrU
DIy3zrHkKASKCPhiW1jaWtRoFRltIC9Q/6m9UeYHHTm8fcUtnv+z9Nt+xcjj
MBiCNcZ48QkG3hSbvIKZH6ZmU/J7F7x8ZIFoLZvuJARlqRGV2T0xoth+W1b0
hk/ziyPDG2e8h3c+E8o+WU/0TiGvCvZtRe7iv5co9WCwikCunuYNaNBHHsYr
/Bvn+Q8ws0bqVcv/3V9WtNAegl4ZCYe03hYVeRZlIO3V99CLmx6w+qYhxnd0
YufktRk0Kp5E7f0aw9DcAuOamJev7sHX4Ax6bvT5dDOD6wPYhfaFzzKJ3cwC
1qJQUrEs+rvmfYBGU2zbZo3sdDsejPjzgcdfhRlBUak7kBuMqFOIN0AGcyK/
fAn0cxuEEOHxhOfmIhI+QXgJl5NAd7qq+M5aHX3eP4HVEtsNOLNxZ5XR0xRG
1iFhumy/C0S7zIv1Sq8Ig/S0sRb5ELjfIyrRghuErK98ewJOynh7Bu/rxeIN
8xR0Otq2OPrrwTKLz4xyukLbx7qlBqt3eqtyYmIDOKZGtRjoep7fazx1FxFP
xkZvtwEeRaH6t6qqHxJ/OsbwaqrWC6psK88RMI4Nz0ly3/0jQcGV0W7N295k
bhw6bAVJK279QTZ7ChZqWHXjdi45MO8Jbig5mKmeQnFQfCYzGgd0uCClmfaz
sp2aerDdgBe0nOFlyIhTwoHEkPDT7/2blZjXX1LvBH5GN7zP4TO/if1v4DyQ
OoAxn8kCQTj5UnbJEef/0lDzxjj5RLEWGNsPfdApckmVqoMsWOkEXQbg9Tng
PCmM6Ak1CstrL5z63b7MRJJuEFlQ1NP+D4/kAGlTYjpTBpFz9/bfUB4tCslB
/WFEGILl7EXAXIivWkDLLnY+Ba6kL4HBOnV4zBZrZgAi/glGnOHTTkkWEaQq
U4OTpZKYoFkJCLTAZgyYMPE4Vw8ikSPo7lvbaNGjL8LcMJP1avfoFfOR1Yu+
dVwrGuhJJbg5c+Z1eO13BW0j3ad54c4AqmbmaPpq22Vz49nQGImXIlCyVgjQ
svDMN9L2lriuphbJcl21LCr2ft4GKr1lla4bD1DMQL0R8qvCc2hMmRSvliDP
Lh2LXG/zBEuJustxRnfshMT9fi8QJjqVdcXNj4KrlfwCtiweqOeTtFi0Ep1c
PGojbOQgkIPwrKFdlSFbl+BechGlrCfAY6NRJ+GBr9enhm7etPki9DGDDMvl
PFHvaaAZs2mocjz3tXYjNTZ4k6maHsltV8mC/b97bEFNknGdLxRHXSeoTnKO
TShusXGIFYEBJYWt4EXWXyi+m4f0LHSL5ZACMlfjRQ+EvGQ1Dn+FWqdvFvY/
wnFA6WcUzZQIOg+EeCmHNarX8iZKFAXeymGCc0LE8ngMhRFJxPy0ZXhB+bPk
OBDyN+xm8+BqYqn/rrEgiOJCit2HubZnnbnPRslvZGv35U1TG6QIRoRdD1b+
7K8cMu0mZ03dbI1pIvAqAPn4FwOHqjjoY16Vkmu/bxt7gdJm7aXHJnxAfrLi
F0T1nPAZ4zn+1dw57tKmzs1BVi1eff9F/jMQ4/t/AaBbrxhmxpeIfqZ/VNsr
NjxzVIR+1CVN7QWjkN6OaSgSSeiD21OJ3y97BTGlf2EtgM4joKeLanEkKI6P
MPgUZbueH0bqvOEpgkPyadWQrwNmPo0nR68/fhIHxzTBc4n5ygz0HakjOZwJ
LWoiIcK3bRqa3bMfhjFsL+riYU6rtk5puFF3J3wFis1U/JwCHn1ZkwYr346l
tRI6OoxzonEAYPZGoeG6Egl/ZJ/NCcOGutQy8SmmYZ5pOIZZEe/HfZL11iR/
7BPCB8ZFNWmpqoFQDbgG1U5tUpXEBkGfA5Eb9biuRVpaylO67XeA9blW/Jgr
6vz2AsTsEcKh3hia995Ge4l4mnre7gTa84Ic5S+UQaoF2PfDfRXYt5aurTq/
Fdm9MSZ9PkhueUGXa+VllyxaV82D18RrYuPQ9KHSoLUd/8Ubgnlioh7BjsBa
pkXr8yX08RO/pLl4HK9Lu9OqiXhJGbQoZ3xqqkTUI92C8TzrapzS8ebaxog8
/gmGlG5f++YehNcU5cRCfbWYsg232gwDkPa5DcyPmW3oUb4o04uEsWs9EPPV
ujpSQ4P8jaO2Ow61RImxDaRccz05B7SR9EMBJLc5m1uxSCRd3kja+1zealsd
PKOmTjYsdhOlCaewAmlhEPheLMJteEI/DnqKYXUNiUBzPIgQsdw3d2cNtSEC
zgk9EFlpy33sUUzQVLzuhMwnLYhq6Sqb7CoIysHH0JQdgHsngLiMWaURKUoc
BBNwy+yPekgZTqaJi6wW4AAtlPKW0j+6vx17FouAcCrSaYAaBeHCKZCfgyLQ
q+UB9kWPdmlr73QlaQcTyThcmHpTt13So8EHmYPFbRD9ItLTLphBMSRjDsWw
i6OIZT2Uu9w/Bi12gspLS2uuzs1x0DDoAE0AoedQPgRTIEPlfV/mNF0zYUAF
b+mGPKrh6HR1wu+Le1Oet51iybYUXg2SvVNVCbAxmvGiqrKQDvYdLyblZc2d
Y5MNUfrBfkyWmi1mn7xlEbztv5A1oVu3VS0LTAgGs0xzD+cnEA7RA96szTeI
UktMHG9tXWzH2fiO0ViuoOk0Skv+nMM0EC3P4qp5BfNOT2GqZdY8CqwmTSYB
wMlkgCQXQUE9b6AIttLNQDc1TlLCsLv1h9q4SqCLeq8XCgaOOryBYPNb2QTq
S4wTgvha0rzlgUsUoyadRfO2ThramC9PhO2qLgysJjiVpxMuv4gAzn33/dTS
a6qj4V64deO0VDZbRfOFEEki/uh0/+BQ3vFybsQ9tO2HIlgtX4/Cmz9ZDYVM
afUI5WReluGnuSnGvphfD9eGmdMxb7FyniMdKBOwGV7ATYpQnzdnta8mLM6b
sr7JjueeAcMwHRYg9lc+gAwTjk+HjEHzT3xuQUoByHExWezqhq5ephlHV7Vs
DDci63iWLh58brA5Ase67T66NactsNa1fjv4SMObx3DUynhjcZm4TuVjhDp6
ENN+HivPKKDhOmEW8IYMTHY2TG/k9w3i7Cw+ifNK15AVPsdgMgO6Bda6pgxF
UfAxnqob4xRqm8IqG4mcz+p/twPunFEF+J2L5ezzIrtswhrhDxpqp3XOH5vV
cVaqYPqga4V+Ul1mklP4AAmKALmqEk3+rZYNcVnr5jdBD4age8A8RddypCMO
QVl2H/nmlr0iGttkCxVIm5wtoJi+jckflAL1AC16Tx5dScl0Ujw4DYJHgeW9
D8tWNAEOhViHH2cIWOhm7LO/cBdSqcA1esffCsLdhW4W29j4sAInF/NKpspA
9zKqOXuQ9/UZX1EXQ5zqInWAnoAHzRNSX4oLiYyTzvdik6pTCslqo7GxkQ6T
oZXNaVtAlfG9ftlNOEFbm+FqCEf37cTTueDoOOWj1CbygtonRnbmEfqzklnR
lmdQNvV5moaG9tzmlumHTp/ViCMWKMHA/Pn/3TzWIi7b5pd2oQaId+QUeNQm
0NVooF/rYC7AUeswQQZyopZnlrJHG/wz1VfKbCbvn5yBd5V+Rv+upwASVMhj
PsYPHdsAtusYrwvk6ROD3LKPAiK8NQRj8+YhJfanBWDCjcFBjm1CbYqVvob6
ThqI2N9VpTNVjFKWTKnBVZbrNhb06pO13pFBSmQsln/w6f1FQngB6KGL/vE1
lca1MCQTZsEzwoizvC06WH376+sOu4dGBpy6VsEKWLPEPThM1tgUKYZPwKse
ObU+kQepEp3m3pu0nlFPNgTGwvFZHsLKs1tFR9Rx2EGlBopDNgususJDpFE3
VGZ1kHoxy4TyxYtc4+vkLPy3ukVxlI55Eqmdm1XWiGB0xNj1kgOTAFZsM2x4
IFK4DDrla8ZNTWSVdmEdTZFMf7O7NEouv2sPdXbtPSFgAD1S22gAuBVuYZV4
TKV4uF/hIoELqmRBCqAvS+cbfbN3eMxgSP2eXXOlfpX+Pt0rUMPyWsZ0qGg9
ptDngVtjCh6noFKKminKqwBb8Jyrs5LJiie2FUxy+UOGDEx3IoXjCOt7LCbb
mLJkBS41UUsxZvZcFFUnCkeU0hpomBmA8VrVcl5VGQU6MEK5x5c/6jUKWyD1
+TYbDqtlcnB5XxA2TS7WIcxbnNLPY+CQ78rIGAnQcKo/DrhhaXlbFpVnrRnA
rJHgT4hLPMbmXhijAkIQCtBqH6AXu6Ad49yVTYy8pnrFNoAzfn6YQ2JtVJag
BRtgz+2rdUzQz/lfGG1Cs0G962CqvU+SILHm2fFN1DlCitWmYxtCEsCMtlS7
JAyvjMFXYuN/ADH7u8WFc4dXbTfXi1HgpxZSnHOyKr+8TCYj6hnwUmKDFS9V
TcmciTveIcGNY4Mh0fftya4UvV/Nf/N+hcXqCU43kUpsKB9Wtn+KCEPlseCl
tEijqAzFeIw813N6TQsaOp9YqDCmho/bJxes5omxz4waTtez8e/k3xAnPErI
KK7XzICIaBY1czgsCrOCwi8Q4WuUDsrKROIWR456f7oYvtQIXEodjSRHZTph
2FyXgmIawvNAGCJJeoVI2B0mQEIvfv/TVolKC+uqA0BoDQdC+wLLK7DRHcB9
369bV6K5ae78iEMzl4THVjFsJBcaTYa8UOcZnYjQURii1HtJVi/9Od/8IYuH
cNaeb+AX3HK7k4noAzAlM9KMzd19i0rfZwftU89YMX7WqtK+LRo6tMYfbOiW
qatLWBB6mPtPgjCYdr03GD0tO6kTrO3ZUEzMi7d/5pyhmR1EKL9LTHI+gXkm
6mR1wgJlOOehSvq2rAdCMD1wbiKAxUgbdCMCx7puKw0Ctmu0WjwHzMg/gj0W
txPXmuWoPzLlXJwiXtxIafGMRqcyGtknIxBmmCW3mU50BstBS2TjYySbTFhz
5W2om0aekd+22xutZe6hyVAb6Ozs/RA8i5jxGiBalJcfOSShmv+Whi9aE4By
lTS57vldW0BLTGSQ7wmxStoBZyXWZEAyrqCsxPoK0nTMPsWogFHBI8RLLWFA
j/NGpxrRzQ0YI3K6lidfQzC0Hqlgrv8kUP58FzX4SCqZaBZGRSinPdJiWqa/
pG+17uqK2VfFJAVTVmEUBuwCEtP3/T5W44uHMUn2Yi2SG1Vik+a49i047Mb9
aiEnhgWT5k8L9fY1pWIZTGXLLg7XrMaRmmE/TpQT16Ko4z3OtWi/KNN4Dc7t
qXVtyCBmEliDbn/ga62ocyLi7+c7xadULB3VtQPG/tfOdJFVc2vUm3D7Aj5o
jrZGJ4D2wBzpYUpyzTNjrq4BM7rPogOg6GlZ5cYxhSTb/iLZWZMPUXfMAjFB
Ayr7E/gKDi41qxFu4LwclaiXJgC8mEb8+nGE2frSRblgDp3bEf8jvDbj11Ze
k6Wi1FSCJgx2pQUTSMGeZtpCL3/+Ab9GoMBU8xfZk2uWRIcnf+gsiutgkMVc
GbYh4mUXYj5kSZVlvpY/hrk6tUjCYWSSup60Afx0rcHMUqh+Lpza3DgfpeMu
iLAboqHYlBIiYxfuDo1s4yR62NEVuHzqkKuRmPLqfb4BqtXuww+wonZ5kaQB
XkM5YpI/CVCnI2hWaFqKzFEw+/WYLH2UcII8BCN9PuMYBrPoZwFc3CsAiQBJ
lgprat6vda1aKHxTo4sbf3IiBexQV6gpjdieYLP6wDJOHsQtxhbRUNTTPw8I
3Ry+U+XtYYbIZfQCQI9BMoG/MfsmcEAgZXf5BbDXmgdoVJ8Q3kmxqihlvBX4
dC7nzfcdUSp3mc/iBcm1mb1iwHELZa7ZoluE8eccXrIggTiy12vv9viwDg49
DPg4Bu1zuE2RjUZeuOewkMT2cgHFlvcdAU+7e4dcoLxzuZ9LyOi7xeMCWtLD
jMs/ia3/shSL7SReBFkTSM3LfuGDg/WQkA3f3SsDRoRUo4OcEfMonv+34jsP
dF3ifelDbc2H/bXWsF05vjztLNGSuqNJynjgBsJpAZx/+oEZ/bcAq0cJVAAr
+geqc83Bgtmq4BhUqt/JS1cmCJrIOwf/CaXzNpiF7CW4TXVtjfIbi5eJBw5K
dpzwqzTfPhaw6FKcirhDHxJmfUDB00bPMLa6TVlSpsmw5+hioUQ2MGRKUycU
TZFwFbKU97paTE9u8uP9nKUlZxkIEWCkBj6GY6y4IyN8eYtPK4CXAVqICMsH
MOAiscmbC2XQR+Ofrtfm5+ZoyyL8EsC4EFwYLeTCy2RBmaFkyOPm9Ednx8Nv
U5N0Ah38WiW7hBw0z7ehWYLVNo88GHg6rpBcej9A4PQEjYfaTbOqmOdbbaQ0
zEsl0fKeCR5R8p63V8L6c9KSX5Iuvi7vjkXjQ4soszoMuhb7+DVa1JJLYlrY
qiMABTJETplslYHxBBsGJKDHCqhzKyFjlA6MOXNGYQN2Y82fL2yb/76HEy9d
TIC0hkuXonpAKZAuXLqnYIxVjfhUOVPf6JSzR9Xdwj0Xd8ErQKL+znQzHp11
0URANignWHdADqR9ww5s1wPcO87+kiKy558F2fi/dyeOx/Ef9WEAhzn1t5gd
Nl2SRqk1XqLqmJbdV8S6W4zaUR1yjewG8K2kFfIYMAqavg7deBhJ6yJsYO/P
hUZijNqkMNVRpv04WsLjNs23vKuAQQVj3gwW5EiHNWlApftVAiZoxTG4g+Je
rZW5N550CfdtnMCcyBIzqqEPRGycK3nbTwrcSLJr7nFz61m1hB1uyXlMHXaa
iD5VMXa6Tm+wt/uckS2vXipoJ6u0Dx5m5WqF+eGngbyOkxB/cIjbXgYJxww8
qwtxSx4g6pGgjUqNlGTlcE43lByUu0J/ska73RCXUJg/+rrX/M9MjOHlU2GD
t/cyazTI4UMRUb1LgGsK2nd6Hz1rNwTCaPYwdiKzCh34cVg1rmGiaEeH7trc
ozXVG9955Kybsvat3eQJS7YbY/n3WWZsC9qZ1hkME0pjBBTEAVOdvlRUGUsp
nfTFjjkF/+jtkfhLSVhXbCG7LZG+T6PnEZTMausESGPvdEeFUUP2Vf4eujdt
dJrkGkMNB9AAoDhmQJZDphzP0jkvrTeEkxnMDIs0igllF6nQhW0n7RS3K+be
AUctnUwGU0gg28q3ZrFpp6QvxsCCqFM/q9KrbtSzy830fA2CXHdqoruL5q/M
KKINZMukvbSNlnfkZu5XOr9+2KvVGvlvDeytjj9oGJJ7q+NV/UbP3L/MbLMc
agsfs+xeR71P6/NpIvD+nhzA8cYs+hd7x0Mdg8tbExo5+d5iEGMbUA+N717z
h6CemI2Rh/HegSAjuJVVzopkCnNC22ogA7Ji8Q1lWJD3RDg5+EM5yfo8si/u
hbFaKlSakKkrnke5FNTuFXpHM7MGhzV5yi0zVa2xcHThQoMetjGD9n1sHLJG
vDHrFlGziAk0TE4wCHnEf7ZwOXOtuGJCj3R4akYjVmPJVo1xna1B1q3hxvaN
T2MD++PpcL9w/K8SjfbiwmgJRz0iQ48YscO8h3rWN6H5l7HcqD2QSjPzy6UK
J+d2UhTjge3C9dG9HhL8kynGO9twgF10siMBUxI4xGKBqT5zbgbtJhEd7ldL
orHTmVhyqUCMYmq/5AIhUP5wFn8+Z8kXYj774T09Szogs4DEV3M+GOpEk717
Hw7lqWt7TrwfvXzP0/kVlvmIdTkcGTLgBCD6bGjg5+LqtuRS9jQ/TYZYaOQT
C+XJ9X2Jg1zVnHp+/NXhbF78staCztTXte36ULXx5pHEjRhnH68XWXy5NHgr
6Hj85WH9Y0N4JLi4CLLGAwMix53sb7/VMEz8Y+YaTOTbvOvSHFYADCt0r82j
PDV38t3anF2GPa6HuETCT/v5Pr+hMEIth+hbnd6LJGeRd6/3bBSvBJ6csnEG
ckW042hVpt3GyN9ot0bnRl6LeOLk/0xOg3pHTbntDxoGeoke5POrACeYqAr9
L87VJdX43AO0dokKiFNFC+r0NRV9m6wKu1YjN8m4mEtFYsoY/xudHx/rDxbI
56sSWo6KRR81dNlB/WH5WGL1eMhcWp00EkzrPWHEGz+dxgijymU7Qpn2D0rS
dIJYUoZ40gYESBPqNNcusPEqj/YXeWgrfxcwoySwJTVQGUUXfhcniXTWq4QQ
0gXH4hXBrF9N2k9mEl7hmMAVnULGfIrmt496/3v5o3ctTUEg4/CgM2URURpU
2SOgCiUlRkkw4hlkvLczp+n90rxQ52tJQhZPY25V4EPtoonWvLYM+PHyz453
MZsEoea7Ih+vIdtTAD046yQ+zPJBuhtboroNIamraMa9+O7L2hAQmqJLRQU+
ToTKRMqn+fxi8pwu6rKbhX8SGyB8HEgMVL+ZFfkc1XvrB2gf/PZI6vk3LJDA
rj8S0qO1vlH3UAzqhM1DnjppipOJTltnjvBdetdM+CQMWMeqBBWssjTMrWVT
DUHR/egrF1jFqT0AgM9vBuyuH+klfjTW5mkddkAlbRihYFJP1ZmePd9bO/Dt
A35sW0wFRUd/XajaOJE6FpzXyHL7MwwPvAPYnU1DD34ZIQKTyiWli8I0TDiD
JSCQNyD+4jo/Cj0/CAeY3jXyuQwknSBNZm4kI5DXzedK/+XeS7iX6Eudu7bt
6il4SkXGsTxF1h62u9V5H78n2rTXVSC8g56nu9hpNlBt213f7q4gGiUNjlxE
lHXogMTKiQbrk5oMhEnyJy7BVq7/RgcRh6WU5NkBEQI/3rK1ug1NNJZ6K7IM
SBlcI3q0FyCCyrkkWso5GZ1c90C6AzbmwBJE5fXoagbrGVsG4HsUbrw2KMLe
MrDHHHPBk5hmZssHW6DPqrKL+PtIf5ruFHulzEAcnyfQdPxqV8jZzDDHwcEo
9wjGNboTqX7nBwlXHADFl3KofJKrPORNkdZ2n3UdPiuEiDv5Lk7Pt918FY+l
ZT7QoSEFwRMmBMusxxUndI7yoEtsOMRufooyb6ZZpeB1mn1WPqOi54a0vxOJ
Wo95+7pQ66FfRCOlf/TGhzSRY9CB252BbyrsrUOadTADhex4DILr9byeGH9D
7FubMJ3P6FvmidpBSa9imB+EIuEmE1lsUg5opQqdlnXj/CaMGbaYf9FcBYoH
4/s3j+uXdeXDKMcCaOgPiUObCf7eCVpbPARjC6sS3/LypTCHUUfxo84pl0xP
SFYE1UI1wZyGz1mUKiAGXEYkRnA0gwroZOFLKKdrEqc0YOzrVEmBoF8n7CbY
k7bMfpuvUb5DQ+F/udYJb+uRf62coRcQfjedAMn15Y4SMsj7CeDHcQRcsiZu
TjU4VFtJBA08s2+t8Dyzko0gICTwcT1AN73/cTdxVSAGOHhQo8ME8KcRgeqt
Uts9CqdN47M9YftFezOBBZXnM1T9EdepLdRkyMANaRHi6iAhu7Q90HG/X58T
qXnN3LgXnGDKxzyPug4rNxXpU4CUEImZ24jcwCPbuHCnOWjR1i39xlS3gEGJ
nRsFX6Vw0s8yh5ucImNXiduVO+5uXFcqCoTeR0A4qOYfAvGOZMZnb9W9vCKr
950XsS8+MDOwCMGmnLHdjQlCv/bQCDXPuPVSusxuBQUramwewPmzXyWaguGU
zWz4WW404FaKfHklEAWz00D/JxZhaj8WSTToco3Km16TVEDnjX5gRIKZSABl
a4SGxkNEzxY60eeLzvyA5N4Sez4aRhEaKElJ7NM0vcN45GIJc4bbttNrEkTg
9YZC3Gtp7Jvpo0myRxYwiD2pKbghTkqen0uCjPbOzMUVXj0xNASzfgfcVBn6
yW4IcLLpG6LXVe7/qn59SL+fZdmXYDfnpLQlulxq78bOmjBqrra/sCfrejGN
+vNuE2yeA3b468EHFhAQi9R/tJ542d0M2a4X1TioiG8YMTEFIJnQjVyVvt37
ZHGfiCP+ncbRuqznZCIZXCFHvg6v1mfHrwEV27fbkvLknP3Q9I50AmVgr68T
ynOiUjAFR4sN3odGXmVq7MZjrLkomyw54LWoie/PoCr7iegs2P1HpPIU4Yxn
/pS4bvAyqvsIPST7wBdU2fWXN47UHhornLA16MobXZ0jnN04gyISieS0hSnQ
NMr5BUBaJRKbjqyeqgAZwylswyofqsPKeZtTD/alc3UEzGcG1POaFJ2yy02A
ul/B1ZbiO8r/11G0Zvsl2oTxBclk9zki5uX4E1m+etk7zQFsy1jC8LjCxi2T
+W0ViViIcAAW1OAdoqGVqGyOsepIx0aa63X16HsSsPNRyFx/EwzWaaV8k4RN
9nZxZp4YzhzX4on86u+pyWHqOTWzpmOAELKqkM517D6yHLxYcGFjPq3d6RHA
vMYmIoKG+UJIXB4Y5impieuoK/kOq8B92yRM2nmOVAo3Q9tBR5edFzI8tIap
UXRnNoZTlP2GJFEcOQRE3ujDeoTyagLj/OEPwvsrNJBJJjF2PZ7m1d4cHBSv
KFwl2SsHarnZwA6w87TBvPAJDf/oMU6c6nFTnRDtYAc0Zy8USHmyuURrFLL0
QG6hGSUmtRu0FLixDwThENc/QLCxZigdnRjGkkIjxT9KzR3igSFIW/PLII4+
kb1fAdYFy7vGXtvgaws6SgR7PiCatJJs7IklohZHOIofRIo5Qdp7fStuBoeu
qyQEXsgeNq4fKfMeUWwTi08KsZR+A1eDn4JDyknVx73LytyI8aKJulLBn79x
MFU7+n3Bfen59ABBeZ1AhC1ozlPidyU+AzxfmjYybh3XGnHk7sfRTx/AKKcH
tQEECfhHSpI/lt4e/J8ZZUUpwPiiWZyuXvRlS32ZvCfI3IY2vN+kbXlkpHf/
wxUbAO5OV9gQOSnK7z/2bIVWUkhy7ToloVX227VO+GanZ555do+tqOTAcPJ1
uwBcM0gQNfRRLIk06H2667Vrc3Kwyefadt9th5eAi9Xh/pS0F/Ous6AFdF6r
4Vz0MDpc1S3WvBMJCXMVSBq6TswWL4NSq+SzP4prAUYEIXuctT8rKodivdIN
pdTyN4PO47UplmRVLK10XWmY7dOHmK4grDwR8hl2vaQ7IMEubSaeEBAZFM2B
2eWq9r388NSejz++MCZab4ETgFrGrRFpFuVr3hiji172lNcJP0/YJUrxAbJR
9Cr5BoJZiCLgC3Jyu/OnPa+rulgBendbRgcV+tpS9MMCEFi9Co7fu3Zv+uEe
q1ii4zfdqQduNWdbeBdRkwfbZ9iyK2nPII3zVjNExHySiOERIWxJSBAswuIl
E9H0iLMfaU0j0afb1yUz2df1EOPi1ovq9EptsueKNxwTXS+6WpC3VtX0yLr4
bGIy7bu5mcRWBAhjWc1vbAAYDkuofhhbXyU0gcVvBl1PetxXQCrG5daKnGWF
+4lmsqxaeZlC90GNl5mHqb1LSHQnYeMuMEHO6aaCzV4zEt4U5oiCVAW5ZyFh
51BLnjQnmqOc5Sjj69P5DdunSOMBo6ded5i9hfDniplCmf76LgS9bj6UC6sG
7lSKYU7NHUwIDKBvyucNRclzt8Vy/Up1aYDIl9qiSRvij0EjMxHRO1YV5E+0
ZYb5bFxTvQgzNrjdqhXp+h93CW2cU5pgOcYyxjIu3wnPY9EijZU+DWvxKXeN
TXKwDeD1LSyB+gkFXS2NLLOLb9YvnPfKZj7htqW652gvKZUT2rwNo9oWZ4ES
rLMSHDlinCXsxO4gMLa6rDarJ/2l4Owf+MxWbpEFTvgnKeC17exlZz7Go3mW
ZCYKRLw345P2jO6FJaQGYQKyjUjPedjaUHkg40v41cCAXMRqRQew76pPWX1e
3A00F5ifs4wsXKz/ul8Ae6mi3iIQSV4spfiKj0VweyF0A0YbQywTqDnEIyUf
MbhdsXE4mi5iVBqEJmc3pv7gyeFnjiSlNkyz73StA+WfY6b8UU3SZ3rlfs+p
PTJPZ/06sX7BddCqBEjsKO+ChznlwqXNlUacBXlteg1HtSs9/uspPp9iRFd7
mqR0w1K9eEiiDtJTKSwKMeUPrpK1yK/Hsj0pRg5tvEKD6HJlY0Dn2owvfMsf
oEDpkcV6gtahhCUIrlreYnRUznnrC+iLS7y9jQ4EPOAy8HncHFp5klmPq8no
fN+aMcR32LKNW0HeUmZxwPFY9UrNs6RXEMYhv+FyMX74zgmPurAshKcxOKQi
j21LSHk4RFjrLxHdIsJFQnPPkAAQ6xhieP4YLpy72ishhDyFMKXu29ydRZr9
/gO76kgmp35sYapZSRAW/n2cc9bIafp+KwL0N6cLzr6pr4B84refCokS5/qh
cGH+rNldO6BZSdjoFnc4dTHdsopzrcu50bbYSrIMXrqumeWqprYkdM8NJ9tZ
9decqIKTIpMC/r191yxNbBVkqoMPG4RtudTRvNOiiYgD/qDXeqoJyLLiO3tL
087u5B31+4EnhPs8ocrblLJWtqB6EwCXPMAyzvH3y/hXWdt/8txdHDqy02LA
AcrVFY6xwVrbwVLPdtHI8/jEWagRfXFCTndUxMJiLuBq3JGBrBzDEtH4t75Y
dHRZMOv3S7u9V6MjgLNTJcjSSE9FBTjODLr7sqZCO7HrFnUupxkhbiGSG5zI
cG1TG30yglYXKwnj8pHsTegOBxTf4FHgy1AyGFCBY0Gsq4CZj2cnWgcbPsM/
iwo4aB7eq1NgcaqRlrIG9xotRwJjbLZJsRLtKOJoYpahjhJWAoOIKaRCkXsO
hqlYZDVVkqb9LdEIw1V0KivE+bflOj1MSKFIrtEZuQM06H+QLbUiY6YbgTWy
ReItrqwxN+ch89AiL8VGQzKwrvfwTv//8Kg620z4GhUM2TwmADWU4+/wNMiD
jSls2sFwr4fC0fRVjs30xjnXp1jZQQHjwNGDLz7L7Fpiy2xJh1/ErovDNe0J
nlNmVSsZCaTL3fLSjjRKFscTcbM0Zjca0GFgUCbRFnz+C6IYvHn7cvgk6CUP
eeoHNd4b8VMeAYddMPGRb9khk3Rt8K0nFaNTVxZ/yFXON9ODNgvvxgz/eD4x
EVLXA1nGb2WRSIpLU0tjpB4YDXqAwasItKF1xDnF0ahWAACVD5yZxJiBfQas
Oi8noI83E24ksnZ/d8OLabwMdKKrV3x3QJMeqEdMK/YmMX8tUE/7DXjMgQoW
s7wB3OlJYofPg8dH8ZKfRybwAbLA4Q2OEu9T3Kn/IKDVTZFZO+sz3U6HmtTn
kjEgFBeINbCCMGQ8rNmYb84To5ciKUXi7SeGIzGSMabBmtHxB21OV8Waj9K6
XgAyVnqP6yel+vQ+Zi/jYha3+5XZxYGQ+02YgH8BXf2/um4Q8JIIs0P2naQ8
Im4C3GbQnusRe0eVQV6A05LaN2ANmDhM/T5QuyKR49zySnn13bQG8rOGsCTx
xuOAo1h2UZzMXwjjenR3BcUV4fIq9o95ZMpmJj5iqsH9Ci3x//tWHWGlBbun
LdH1vARqtrKI+CIEhw0AXfr8cQlOJjLazDOoMfMy0wcbQhKqsKtsPw/dzbUt
pOJYQQf9pWUZBSUJCj3DrlMqNiGLCaCANdhKfRSLNzJ6oP9a+lrPakb2HiVO
BIxzEwmjuvb7NYdO64ikbrEP8TtX4QrnPJAI6zWXnvFvNCi844ZHxoVrFGyX
tzBd42f53W5d7GaOwnsd4bw80HfvojlESDfcU4cwFjTnMt2xscyhMk7PG9q1
zockjkV2YRwlxRqgB3vOWn9CjylpKCfSrT4geMGSo37+DKib7SBVuw4s63Th
LVDwgZcQsQq/L0NOm873mUQkB56aZAiQifE0HCPUI4GD3zByLH2BlsV65UFj
0Pi2qoIEMNxj81qmLdZTYLDQlHpobu98gptp4yoXF98TT3hkOmFOS21auOok
hx9dxFMe99rwej6j91fbyyMc3kJ0EYKqyPVaLwjjwXMVeUVHC2IoZtaCYO/i
+QQEOq31vQ7hg8R9fBABijpGY5PwlAXvNxJqi8O4YJb4vHOWZSMTq5ICzL6R
SPNHOScO+YdUiPaIH8+fQKnVL5kLIgwAcge0C3Zgh6HET7TGI37+UGX0cK0B
DXHaohZVVrlVl2jo0yX7+MEZqFjnB/M137SqOXl+xvDgzcBTEXzTcxBh8TXC
htONBjlwoIz/btDxSiyrsX98NDGZSo15MXYessm5YS+WKSdJGOmm/B/VgxAy
tmDE7s11ihC0A+/MwxmIKSwwPeu9WShK+ltxq3RSVI+Cp9iaNqfp93qRhkDP
OB/RBnjvS8+LkVBZ+oPZWamtYIgiAnpXH5kXe1z7Un5AWw6uon9YDMyg9vdj
LuZ6ce/nHEp3lPvBWhGdIeskPWENd5+hmyXroIrQn4im9RZ1d9+xzA3ondwh
8RuLp+LF5cEpY0o45whiqQT1T0OsWo4OGeF0g/RX0WA0ZTlMm3HwpdCnHJIA
T6tMnlI6NpxBcJ1yq8bqNlGPeYqNLrIDqxYhMlDFbizY4dDSyGcrp4wSu4lO
c6MNTZg6oQDguhT1y0+q6rs2gguZkbjWj6g55pAp5sY2E83CX9YFwoyvixQ+
v6pZRwNwmy2zlnpLBTK1FlyHBoZeZw8WuhBuvQZy8Luy4+rXI6h3y+CXtTik
3Looa9zEYWdhXUyx5+Qd3fogC0CUhkSeDlqCoaqqOwh+1MohfE9u5V/6mdm5
ADGR9o+k5nq3zqB3gqXCGTsIDByHXQFnHZpwdcFmfd6xPrQ9gxJ5exJRnNjS
jd+8sBeAl8IiqI5lKQ7SmXrJhzoMPFFKI2VW7VHrLXj62hqPuhNuwOY8SbhI
IK4sL/iZisyCFNpXlzco/0x95efgZ6wUYO+Ee9fwYzrSYxWMI4ycfTCkSxf6
ZP1o5c7uzUCAatVEybBJSpFMyqMrQpOZp2XL+GuT19zDikGxJB3rNGA8aprb
li4znpY7wrDFBKernUBcGVk+j2zE/YWxoWg0U22SLuVH8eA6SiR6b2Uwcf8y
X1ZKw0Dw3dJFLX4yOwMukSzamJog1R7nUKwPovii9TY7wa0TUWwFIYPjHy7U
FfigHoX7xKR+BJ3R7TN9DHnVcAZphxhr6WLkh2MdvjblhTd2fUEzhq0W2xVc
HPE97rig8Nr19VsEN+b9CSSdrja9YKAle1UPbIRqtvfEh9pgom4A0Uh26ewN
7szgJ9CY5g3Sp23djBxdRnm+GFVjw7fOUmI4RC1c0Imn7ifMWu0umA1VcOKM
xUfzy9JoyqdmAwz+oF3UZTWjUSBDPr2GwzIhrb635dl7Jtk1tMwKhVbAb1Sa
KLXM+bDqk/mp1O9rNCYdpMlt+XC6gTAiBZ/zCHx9998WfQICUUzbgvFN2ucO
KMl+3y/MleLYqomdmbCanCtapaw8MUaWTMQrzHa8EKiDHWRJxQdp16RGHC40
gG6eacF6PlwubQVEZpAvL0SphMVFXDgiSoPT1UN/IQJoePPrCPm3IWh5CKVL
Knbc8M5SOkzk4bMCeFf9nPGbPFgUm57G0j2Sf9qTyVpH3I52QGB0VCVLzHdB
Q/aUAE9AlZWJv/BMGMJBFV+melGUZ9KfpfL6jez00JTgFNlqkLf15fATj2rJ
IH/bTI6OZyreaROs0gEUk0/9dQ+IsC/zIiPpCS+uj2865AAeiBEw9tVXzcUx
C/rlc7d1UsLiW7nWkJv17365qooF5z4hfODBzyX5IVMRopgA65ei/nqqXLsv
DYP+yXwCGLL5kEGF5mB7NvFdqYwSZM2YPDPEvfbmlmnLA+P5kZdEwW0jCJ0d
jhyH8/+qTy5LhzoPIFvabsNvgXtaOXbdxkb59/OKwolUA5RtYjKKmM0oykLF
rL9OkWDhR4WYY/X6BRKGXrhQwoD/Wbb3fzwP0zxwG+k6gyvQ36xE86BQLPu+
ULWfn1UPOrv1GczJHBzc+w40fn+u6MgANxRl3LuxXXr7N/gsDGPT/O/Z7ol+
jLJftWtZH7VQM7xIaa8DM3ht3SHeBTBkZcoz9yREUKy+o0Oq6ydeZSNzU/yQ
15+rRXxE++W/oMDYLT9nVZsp76aQkq/pJ62Y+Zqq3z3uIYjFJuf+fmQXATct
cDaj1NrsyShO1tiu8h00GZJF6aBCxNSiqLdU+vxHA499cY6cV5/VbvHmwHoD
+4hPZCf4R/K+s4tlH4MqkNtgoMT9UDYN2P5a/gwEY0nNKB1mS1G4HlgTKPko
aOiADH57v6uD7Txk1pvzETV2DijJ4a8uPM0bAzPc3PkOCCl7mpP33kskRz8V
KmWNLKgsqu8yVnNpCQPmPVqnxd8NiQsZf3WVF4CIwA68/8iROnoJrvpwrHmY
zvkpUVVRGWB1v3Mt/jldF30GXDrwJlzR9OHDmRvf0mGvMZZO6QVoYBIIKo8t
KINvlLBobn+GmZWHl/rHUrpg0zpUzF35+xzrh0YzfEikVgExV9TA7sWnklqD
ILGi2ixCGBKPa2HUxvRq8wA0+VDzaP6s9m99QhSLyNtOIRx95jlJsHd+E1Oz
gspTStGHYtRJrTsrxHgiEHd8WQFIIgEwciIVwn8lnmb3+rRTkDRMxKT3uyDf
wstnr99q6t5J9GPfpCleV5Md3+zWDiOaZFZjr2MxsdSh9jxpErLQFfgrwqXU
p0PNkxI+Mo6zlKAiMYEtG053KNsNlsQ476Ssq6isESIOKUKRRhaCH5GchqDr
m4cSUTPV2buCMQXQtqsRv44hzL8v27naBOOJ2jedHnKBL1c8UbHJRYQqy1P8
s+cKa0ZIW3nE1kB/kCdCGNTeznLJ0ZuDRLATUbLbUaZQYiZfCOeCH0uk9voI
K3UDkcLGE20OdLzuek/s9T0nW8P2lfDEIBQ8YCque5rBgXf+RqR1IVfmr50k
Ra1hsyMgIhMkEL2SBmYgFl4ZfDtT8H2e/IMwgw/m1G3tRCPmUOG7XBjp9mG/
4NmQRd/ASrFsstdV4JZxfy0o11quEg0x4jIs89iB6QuQVxIWGcnyURUWHe4D
YaXysmq9ujOCL/AjEsOiCYhYiGwz/4l6HA9n6gP1tCVvr7yGhkjYlrFAIbNQ
oiUc3df6zin23DRjBsFp1D8RiazDbFqBs84QIu4xi9+vXrWcrleYXF8scEVV
wfySeSXc57ruSI5sqtyUF7K9i9HMMzWBsY139M2Ag/4hrhlpoqM+7WOgLwf+
JOfhI5TiEkAX29wQCLW/0UJnszQEQ7mHuymir51YgVTCVGegLxLnB3gMdp0R
/xUpmtF/cMrxhcS6jYahI/sOF4ul9kFpvjwl8s1VKCFVuJhz7GD95Fdxw+3J
auZmHDkgZv93YjJ3tSXc2b9KBY6q1Pood0Yof5Fh1i7x+n2kCyzjqLfH+lnd
Q/jg4RBAMmc1MCKrbwQL/vaO0R++ha6SDBoYXZ3Jnsr2f73LuOROK6GZAm19
AYBaSv4UO7njJ97eXbwSSIIWR1H3L1QYKza3REZvpCHoTWzq9G3E9g/kecLD
Cdkeb1O0bEVOOcCPUK+N2VQC+lnfPfZN7kz5WLTIFfHYy4JEnk0SBWhWuVOV
iUa+b31KMndcyX8WVQ5sxnlkpm8e+1oRUHbc1EUY865V2ed3nLtybDCJH37c
sjMV9/Zcykr0XbC/3sN4gUXEn/DrdOAXMw0CqHfBnlKOurfIWpgEoRU0KTaU
g8U9cOtOJg1rlyhCE3Kx83Ajw0dzK5aoIYmLg/ZC1WTmOjpwn7aSg6RZFSKs
roAEoeKBIiX64HNR44aGGTFhrKC5zhLYo4V9tiBeMHJ/4O7Y7qGGy6zniRf7
5OWltEN5C67dHdMskMK6MqLdWJIa8j73Oylqp+7awKZtzzq9bQHvW6xV+nu1
TJTLt3r8X8TBovrXPREbfGPlJVcygykePpxN6N8udvmzhJdjiFw/i3ggwEXC
5Iyy6ScAxryP4whIJA2jSzcSkqqNxN8+IlLGqizo+ibDpYzNuXmIsvzWkXXu
I0zcexMn89rfiECN72mBQIhCEFFJLLN+xrZs8yP3ENdYBfGeTzY2AZbYbyjg
kOlKvjYjzxTUCdogQf+CZqkKzYLbHCOHpr7xnr6tFG8IgPYtVbu94uMjYTlF
Jqddk/uAAI+FzcOR244VDnQTTVIwnbwV2X+Q+nu2pYnnqkC2khs94qzF0G9K
ANaapPmtMvv6zr2SYI+h02y6so5rxGpkbsujiZn2PBaXYUc42HCHfiBPi+D/
JkwWQ4O2QCE4FDXEUHPg8LKi1/pT8mR5J/LQn85ervSRnykZdsBPqArNmEhc
bKEM7lKvTmj2A6BopeownXwFaRMT9JLiwgxpKjmEVsbs4Mbt77uhhWdzzJMd
KPQp7ZHR14s/k7LiFmjNinRkTh17MytF4fsxXr7SlBpGMW6WPNiz0Wp6EcBa
X9eg2hWyYt7MZp9APNnTfrZQi4+j7qfozH3UZrxDoSzrOGiYLTW9zfOCPE4u
fNXu/kEwFqnyBxcae5wu0Jv9emQLfzlgwVs+VO/ERD8n0NhuciMd9PFHy9GP
eOn8IQiwVoxTrywfFmGaoPDlZx/H9zRZKjQQCGEOr129LYBkdn42DXZORGYf
qT6mLrtUnnjizIZVFRhpExuRyYNYZlqYIMbrMDe5avqBB8I6xHbweBCM9Gu1
zEL4hTlIM/HD9qhDivHAboxsiTGY9K/KVsoXro1LaW3pkrfMS2T4Vc4ZZDC0
TcYj9SFoC6PMi0UtnQJDYD21uLG9lH8rX+dFjtVGPoB2J/Po/cjW1aj2Xywk
1bFCZt/Eh9sm71k+CToqY4vtnLxpR5oBW6UrapEpU+chIiYD1QQFWtZS2Zoz
ov5s3GJFeMJkKoqn02TUH3Di1cJfr4sQocFTCyerehiHeBKapLw1LNiu0Eb5
0oQqmYxv3j3xqDkp4trCivi4hV22tool2mpPRqV4TI72DA3ZRhjRLPPwyFBH
KsA28o9+Q+Xb9cHycvLlgYdWFG2XJkJxWvlF7KQBDI9lIt4V6n/eD3ARr/oI
XUmCIEPGQBJq35sk7CrBpvsIvvBwMhvLZMpBf3D3TLtWHicKcN5Gv42tB+If
TDGte5cG36u0LWHSEe4z5XxpleASdSnN+lVV7EacDloUdohuce4tysGoDPBf
p6zYcAzYKkIZgxCbmFFJT6d+ZypbXeJbAGy5nqoTfIfNZss8f4qc7iA2Kovv
TKa1zfrdUHox3KZ4f2h2VW2eh89mFupvwB5r7iVbfk5i84s14ASEYQ01v2iN
zq+CoIsUeJSja8Y6pc7btOZwXlX9KTtKS11whqKREBuE/7RxNugQ1WKoPBaX
RCnYIOCy5CEOfXB4AYIPXNfd+ybtLp/VO4h7Spisc3Ih0cYrGKhyrz1V0EuY
22v5pA63p4uVa8uThbEAuN6l4I0shIE86pAVDAK0Fu2E1TECn4VPzz9m4qCl
rAjBhkJjYh9swfZBlxzAEsTdkWVzuVaeSbYyuYKz1kANJnC48FBa4YLb6BfO
7vyAw0YEUCFoQlDn3hpAjYzWQOG+qJIVNOeIIRJlXJfk7nGNDx2scpbs6k5h
jKGNNlBjmJzNPpdDJ4Aa1HQd3o4n2ec9yZMbjd+mVieu6Hfspg8ypKzMnB2J
lSzJp/9asHcc4wfg0AOcu5yHmMVPlzGA4mUe0wzJFrQ/hfmv30kwpq0Kjm4p
LpH8bHv0t9D8X+LLEVAWWGIEYK5F5U9DWRTRno8qKQjW1Z8DeM1z4jI1vufr
upxULwRRqw51NjGI81g4ZKlgX/TVS7lJIOwUcZ+dNmm28v7VGXYQerMxKswo
+dYkqCbiYZIAtw4n9R6V5RBlVSBVfl1yLMUqZ1Fe92XaPl8LjO+KaJ9Ag966
molr0dcx9qFXuXeEcot12JdDg/QqWcu9CiqoK/LAbtg1SfLa8ZSDw3q4V3oT
8IiflqsiJM0w1RsKb19JyxzgbVf+xlNnJTgNkl2k5S+aKd9lQxMT8h/VE7H/
vZYtP5PAWhblwKwGN7Wtc8pFzgRzquWSOtCAubOKU4BFKHIAkFOrXSSycltu
AflQ6SRfHGwV1dzTtuJZkUJNurTOB3a5g8WKZgam0ZY+wnca/c+K9nYrSDi/
7o5GD89oinwoc7lTrUNPNx6wlZfDSKrSCzXAS0lXpblw7OO5g+a3Z4tnFpNy
RlcYyHbRr2vzD87QTtLBWZBM8zFspoYhT8Eh6c3UPwbHE3BtvwXF/j+ab1mM
lN9Wpokh3SlGKLJoCaO0T0hy/ykcvNXl1UyUfPlmXE0PgOvVSPclGahgjWp9
gPBglCEIOHslKmiqifWO4zLXePyCula7t1NkybI1Q2+RX23tkGzeowLIAM80
oH+CgVD3KfdkcVe/9HRhXhXiMm0ZxM3EalroVaD7JEydlU/qKxWPdpuuYtc8
049b9/NCYmlFTV377DCKiSF35tGu1Edc57Erq6CfZthziy5J8zTGXuUY0PtM
Jv4c+olQan0ZXgJdp5o0mlUkE9/8M5eeB9lyFdoupkGZZyrwLXP5082JSp6b
SQYESlpRmohNDls51USA3giU0S6IaRhA1ynZcb26237p1zRBwjLXGcF89hpO
7R9ayaeYI2xzMtWlNJNplUESDDSrKaCvRsrUnat4zhIyTW6ZuUf7CPNAydCC
iCYwuIcbhVXE4fJQqK0UXntc8FbAfGGIJKlLIkRjuP3cBB0Eey4qsWY3pT3L
PZRMr1GnOckXPqOVC3p8Q71Shfggt6xWBBmZsLgGwrQNKf75f7d2zeM30K1k
CR/Ar2GX02w/+IVRKwcDnS8P78147aXloMoYmhhLJEHCLP52S87BKuOJokB8
Ti6tcNtQTnfxlsoPvNUFHc+hrwTIEsZETWSYkAJic95+hQFRbhgskeT3vlWj
YkW/thnFs+e9YqiNubRIf7ERpkzjLM3Ec6YCF/lwtfOLT+tu5ouswvwrlPos
aLMmK7LJNRWiUAsmuJVrF4X2csrW/hkimA2ppJ9W9D4ojN6/3G3VUicabHXe
toa75sWSiqjWPvZ4LSk5QATux0WPdBgxYJc6nsSfzW9yspuEhFvzeVUCVG0H
OfVljnhMigqOjpYxL9TVft/PCDzAvZC2V45CU26YN0aH5Wxc56y6hxkBxUZO
hoGjrFEcrh8h53GE/lmUxUNWOLK/itbv+yOx/EgEey6ZvqpNoEmYemoTdHh6
E/eS484Xu2YefMp6EfNhnZyj1Mnit0QOlN4O5LALOAV0wYN8+LxUyYwN+tPW
se/+IxEvEkyEYQRC+Q7SS5N1yAiIhEjkyg1pBHs5xiXJvxVNVbgJQmCkimzD
VrY/OLd0KSzHmye9BkqIhJg98jrgQMu1Ibq5e2ao9la+oNOOcoxPbkFkRRIM
vIyPnLNFP37AHJhse6F++msc+x9/6iLeaS5QgVQM+czvkItEp0SjYsf9UfJd
gVVcdVPQXAmlHnEogxPJUt+0RW78lp9DeM6w9r4Q+zzJQdKfl114/7eoToFH
V38LLsVHOBcxuNtLfVBBg9P2qy+DaIpbx2NYRY6I3Rwt9DOSyxkRyXupkHFD
jMe6dWG48aYYOuzoKJrsBjENnPDWnIjIlwMj8N8f/UZBtlGjTY6HBmusgnzH
K6+h7UAV04RUUYlaiMEwnLnCKGwHguM0R8Abddg0qZmSi27jAJPqcfkjWKS3
3tWWP4/EFtGhvJGOVr//HzMMrorvYALNuVblK+ja8wym2WJCCfnfQZSG1FUn
QaTSB7CY1BvbfqxV6w/sLeGapDmP7RxQM335o2gJ5rOxgRBaKhsR8Tj2O8AV
AkZO5Tay3+0PrjGODAA5cw9B2GUEv/wLGFRyFXIa75ji8OsXVCiNpBH0RR5L
Ll/4u+sHQc+AW98YiLghAcaPGFVAIw0xk4u+TDytwftPhji/GGCs9MlLgg+n
5ymH78r8xDG+YlCYErlVCaQXrwJiNFFgLy/2D3l92q0qfd3gO+asNvNiWNej
7jqTPs5E1aJ4pPBK8sPPHnECR8n92nvan0P7X/Pd46eleW6gMWMrRlFe6uRv
mBkHSZENdEzxUqgU6W+tLRv9RaksgS7KIgdugk68gHgGKFhHvejfx5IZnHMq
/O4tXcZrdjNfpWjpWkaVl9Dlz2av9XcEtdwCu1PV95VqD9QBQpiriiJ8QB6/
AedqVXKL8BJNf4Rc+S5saLmwAMKFJdtx5hzXkbux5tuL+9m+gNipcJvlZYBu
+bUaPozyv2WRCv8nlodoDI1NbJTIym5lZ52Ur+Cyib4vJxblxATQRHzkvoSt
ksjAkad8hwUfwF++BUVwz2aO+j7MnWKE3Do8Fo43lVSLPap0qOrIfUbNvFgG
BAHw3sxzp1Nd100sII5q3vylNVZtjzaN11pqyZx7FR76usB5DSGLOKCtk95b
f84NP/P3v3mynpJoaavHYTf84CNoLanPIuCqLOFPDS8tJILhcPnWofpMO22y
zS2Z99aLbHmKrB/qMoxDk62IbRWhq5wlWNDaMWqcJybEooR5IzIJZ/Zweaux
n+fXL4XS+BNL+8GWjgDDr34Ojrxjh+sAIoMfOqA6rpykP4LNT/OpAz/fRO73
+NodseDqw2UWL/vkFRoYVk6wzC1vpyeTERLhxOaoHxln5Nxl+oxqNcazLR9K
6VykfDawBPqheSbY5G2NnQQ8D+DofCQbLAeLX/q8XyMqmbdJLIuCu87ndH3a
G2xqt+wsAXwBxUs+9Bjh3C62FbZeDT35/bgXHNsfls4GFqe8zE8JVJwX4EmS
V2qn6A4Weq/MRTpcwvTCH/WjpLI3FZkRq24Zm6dao8imnsjVH++IC69gwlR4
gf42QN9vnYuzJ9jjgvZ67SgTD2zm7X1RdqL1Ib+q02Q8k9xe9ldX52ZrvBcM
u4i37oMgLxgCOc8WURWGPeYZAhxPqglxak25CsD5+bsofT56vB0kZPtpd+Wa
y6o/bHiT2necg5XFlnHWn5P4SOlBFcr6kd/RC1vfVeiKTE9ikm2Gy/SVbnv9
qitESJUEcFGvwWp3XGyvvY4t/KmSRJW3J76wmXhbx/SQX55nY/MCbhGj9egB
1eNHSwqSfMofE926ViA/Dm0rNgk73VB/1YjVyotkMi71yfLGIkYkQFqJPNH/
D8bdtc8B7OfwwCWdfl4KP4hKiGKnXBEAgsmsWSio3cS+G53dveO8EIjtDbAz
WKUDxew3yF2qWH7Mt1y4NRW4D+2Cg65wHGPXegXVv3nkvMXL7rw9PZIaRmRw
ss8OJzFNCK4EMoeVL/AJJbZRNQuf3/GNgmyjt+0EccfM0CODKNjx34kjh/H7
Djd+HOVaNUrs2/WtD3iNMgcPSS36dT8whSJJjFAleiLTIdRgqlYcyhLe6aHA
ad/3LpMe3rT2ALCRG/F2EFDGhREjj8q2GokmYusVenudeULB8rOUnnDudneb
0WvWYGR4Y5Acv44NPzsdDMo7UglV2OA4Yuka9xFLV8es50I6grkWJp18g1/i
FwZfCCEjvf8AUps1kgK31Iy6GRkqSXTC4q/blSdrNzwb+TK2u8kgpnJ+R0ur
799/TkfjBEchnFkWpw6WX2DNXtEfEEBKouiBmiIvvdJR7dO2FAEYGbOKWgWQ
CS1pLDlvN4G/8Z45w6/iECOQ6ybwiDIJO1uOD3O8oX94l+0YUHiZTC7GzDjd
d7CbaYe6OyvYNVJtgmB0fZSKWvHvfT1eUOJ8hQahuPZXjRvM2m0PiQtFlWh5
lz7OY7C6/zA0Lbj2VkckQR3vCh/lExpJMV3KXC6QjOH6mDf4bhjefNB5r/wU
/wQ+iNr+VeqF0DeUFtSxrzCu4yrWfuh2O2kDXLUsuUdkiNyFpjhxWQUN9KmT
drUP0IutiAUFF3rWI3xP+7GIqEDZghVM/bCdBVPbAA9xMlbNvFTiOBQltDRB
+2D0qgU0wGwzYaA1eRONqQxq7nziRyfSn1xZ8p1vF2gfNuMwhNPjwtPaYMj7
pPhOor6XMJ4nlrBFVvYNTIS5B1AcqAas3nYnBcYZCWqcGwFBGEk8qi6yyJP2
gIoE0Su5oex7ibmTwZxXTyeRuK7LiSYQgsWHkJktoyX/rM7EGMhgfHSq4Y4P
bVhJOBIcDUSG2HpKs3pWZ/PO2z88j+jgDLOfjZOXlvWPDMCifoxtNVYFQ5Zp
vpdqWaZV4L10ckAFNvu0/f8k+bGr69PX0QTdc8Lu1E1lae32NUU815wf9Iil
yB/YnxMIYr1maBPyz9F41aUlqsLR1Niht2eZLapyMY2H2+JDla36whIZc+cw
hSPftoFQmBDim506ypquIQPo9bc2oAw+qAC7yl92dtEhpu0wfekWRETKnBzI
hUNSc6gTzCoYurdNU99XBsKxk2YFX1w1gY0H7A0pZlGOzNeKHrOv2rwZ7T/W
ko08P3148usJN6k7G0v9Hg+MsHXdIYTdVv+eJVwlP/jJr2u4B1meYLEbViFR
cBIDcycVLPwV/TDoso2Zv+MsEf5phaUmY6/W1AhXzcNJa7nMQBBn2pz8513G
j5ENnjLNBLbnGK6I5nOigJpuyq7vJ6S8pdY91DTdhANG3yHr/H5C1NMU2jBJ
rAdwPCg0g1eFivYe5bROu2Nqh31qzIYWK3rfZsXpXdQPx+IsRzMHbzFP7dDe
fR/gncOzEcxj1G15hUNiI2vOXm8wbNULNYQaQ877EZMz8/mpvt2LS3nyiSmG
OzYRGoZCwVOCKuu3dAQ55ZU1+beV4VtOyzSCbOXUOIZdX/9P9x3H1tkjaZnW
NZYSILBZafxEdU2yBlfNryNqt9SGqZOM7tMq+nQdOH/3eSxeSYF508GtEi95
zppUn18iy9ghhV5S7IeI9VL5I456tJCgnkcKkLmcc2H0+bNWMaSMpL1rAkkd
mpLfDjXbxX9a47UYzhe7rYjSbYfs44c8rjhLqK094SuAEDFdrUOdO9YyXbBm
HTHkhfTsyRSPdIVB/gyUugEVMfsYPIFJZhd9QRDEAznJpOcwMtM35UJPkq1h
d5uKsfrXYTG5fdEUSlVugoudkWP90hsGE58KfTgXVOEnCnog52LWysZ6KH+r
Z/bDSrboJqlarrrtonDyb0LZKuf9T9fUUf88LgXlsY0FyrUfNhp4PLo/0ede
8IH7ynKkcS+6atEjsd2XYDTRAahWm5q4t249EFLAggtoqFhSJTK7G0rUtd8J
dXZqFDMdGI4TQz1eS5z9Nn2QhffYSovfzT3u+UdXo5XdFxBkJz6T+KWBEOls
BAdK6swK09E5/ORxDFJtlxBISfuo/6jJ3zG8u8t9NtAo1XgAUtsmH+/ybxF7
JYbXA/r977oHV7gokZoLdykzKc29pijudgEPVc4auXhs+uivOhYDiwXE1lfD
gBNMW++vFZNcw/t5xho8R/Yv3qYDLqoyvINiSzqqtaEfBLu3LHpMzonRAlip
jj7x3fft85Vv6b1izWw8RY5BCSAfJHmapHe2BkE4Oivs+euJc+qrmcIciNHF
STaYNSZrRZFF4Gv5ZjhHJCvnz8cXl9P5PuIiwdFxbk2zc+oOdmuhUhWalNgQ
/bigiMPQ47sevUUC1kaV0WYCMufzExDDrH+iXGve3a2LR+1PiwYijSNibt32
0d2jJ6GY5YAVksVqrgdaNHgcd5pIMftMJEYwrW0PkdmnIm6CoSMiL54Zm0ZL
k3EyF3Kpzj6Y8ycbJbk2d/MZysRqbLqLnDzCfgPMQ06oTDFg/D2Mt+++DfPg
L3vxHJZLJVa56y5qMV7w9pfKgodwGLzIRsb+oWkosnDmc+r2qEXSmzsGdCRR
vBNsXUXMR32/3FMLFtVgbpyT2ucXNrTVmRkGrQOVF7e2rBUCTSC90TsAJL2Z
Q3OkHj3MOGok9Th+fGPmSmN8trCP8vBHWlMu4cvO5YcgQQ+LNFBw1CRw8nji
YQ7cbP7WKsYhHaRt3fgpXyZ1t6ZgHTjZ79ubc0uclGbiVDdd5stOU2DfnTdU
TtR/nivabHMxFK8Wz3fOq4oq7cN3Ue6KvTcIA9y1lmFGyFP4zrthghdMbrhG
rznXhaRlNYD1Zq3/mLu2Cl4TrW8xUZVanRKpXycOAuo2/o9f+lDmpWptYvM1
2MMHTq6goidSFANyd81tqFjbxpjmN3etb+D5YH6jjv7a9TKkSwXZ+vAGDoBR
gaDlKeGb/S0Hop7vwES0zgIvglEscQMrMnmdqqxjS8xeS2XWQBaAY4d2Uo0a
AJse6hEK0FApzzvwZnMqeLqJL9bsn7w4y3neddkUAsIFGePGGVW/4ARKQKDA
/pZ95B152O+u7hA3BofCJbzJPoActo54kIxBN9nShr/1SreBBSYJzPjPSN4M
tFiaKRTRSgLwu1XdWwx/usp26xsmPK/5BMeRGoE4vqPS/MzGdt32kibAAykf
PatB2MmVtkAA7ZLMYU4qrGNdGulz8Ffqd/SilJa/GOasXizgW/iJUxIshhnt
q57hNzax5zHtr+dHrNhD08UqhlYuk/r8RoUQ2wzcf2UzWly1jKdEY5rpGWcY
f6hg3NKioIrQPgcHOTNGQZstnNvK492y1Bxx+CyPME+Ue2bsmHw2CM8XySPt
C5bw4FPK2tkcE/ajEFn6FiiZcU2hTTCRhfnwTPO9+VlQiikzgRNi0wvHUVNm
s9LRY2mA0sz4lqEe5oWGIO95DL02+k9TOeZ9Gdzdf7GqMWXtnRRo3m/rW97b
qbZqTOzP8yw1uyHaURWkFKgCkr/RzP1UT/W/omEdpzikcb0ZYUdoULeiTpmB
TkSfBrpyt8NxqBJp1cENgbEaJvgN+gModGPsfiKobIsAkU1N5qVatF4wO1wS
S5mSVbqXp8vENaiS9hLyo6u2yXmCZm5zSATT6ftV2r6W0suhjT0Zz/bCfmfi
VXPkB5hTyAFRt2HO/eZ0qd21NMFrlBncLVUqHwjIhxdVGiiNMOZeYsWoceMs
WIcJ9L7tjuOVqopNkDJTFAylVQcnWYc3uzNpoyjp/7BnbjtoHmmKxqiOH2K8
yztr74uGMYFkEP6IP/Mw5lYyyLEQAJqPhSZ2z/BP4XevKjiebYA0sUUaAcVh
yZkBc+XEOp+IMMKIV1iqmzCcdaxjXhFzZzPmwgBRYmAOixqj/+0WEWRUfsLT
kAkHfIdKey/+u2ndfYmBAG7P8HDcnYLBLvZ55JCrXFEhMFfpsHB8J2n7QJCW
LSCrxlpsn5tCLIyadMv5pDIQXr/1wyBKPllKjLvtgheRCHYqTTtpsMeE3KXK
YqHqcwePfnzYoSfn2imowKITVreeIRO795SVxY0BCrDtPwsj0zWPUEeD4mDH
a4IXmaHz9K/FnQ7AQ7M0Qb0D+rpQckUgyQFPBmx7P1AWDKJ2SWvDkIe/bzkg
XLwZ7oVsS+bHXPSjcnEJFhsdCPxZ36ozz4d77GkcyN/hjDzc7pnnGMrs1pd2
lXnCAKQ4If/kUktUkU9mmdoD+WSZmGzBFlyj8k0j9v9P40AXsmFVlcD5UtZ0
0NidD0psAU0jyr+OP6BFe59t7N26qNe6nA8XuebIUwfYn0/YL0dk4Zpv29tH
scd2Y1Lyg7M6AA3wPQm/WzYAWmGbiSF+Dl7veLZ+j1MWcdNCVuRocVyvD9Ll
YpW77+d0SBICYCM1ME9BQgsYqqDIfCsvIv8yyqK8hXc1dMFSQhwUIrqWYcGp
yELKZqnUblCbmAYaJXQCgxyLprY22tmsScwnh+B1kMNygHnfNbLPpMLTWw4z
tU+8gy6MMZfr0t2aOfx41NvN24ljxl7suSVzoBybenHgSVOKafsZkm9KtRBO
5qAFZQDesXz2+oAhGKnG6e55ABn7E+TKhmbnsUBt+c78yG5PINVsGRv+Cj6E
1KK7cV5yk+PT/1rpJE/ryPryIJW5NcqPXpaJtRzh9BuYVNNWU6ZJdfZ49x1A
qUssO+YxDPh5JYDJhGsnafhOhhHQd68Cgv+aFg8fog6bJoQSkDT6+CgBfwy7
HjNKXTFcb0gNasrLZD0jxETWxwPeOzuBuEfkIGaaoCt2HRzzJVML542AUvWH
KOgLRhZ9XLfmFST/wHRCw/xNCU/sp/wbvFURqMttLqemM9+qDqk9fpIMJ9Iv
aBzl3G9KEcBmfzRCPIKs2xnxL3T7m+sR1QVT7sNKifWyH4nJ8JbtIYexVjNx
rh4wUAK2JINLfP7L1Zr1B8rppVQ8W4HKAXcrGD7qmefvzi8Z5C2YzeJBIfvG
CFfOQe2OLQ0MsWqZxSJ0QhIUI0gMuYR9f7/oVVi3nrMvfiloWWqjftpXDKhM
g4e2c7yvX6ABMArZC6TMshM/NVHzA/TCazLoTFQik2ht7hCwyviGsFX6p0gY
WCaopn2tVbdKG3TBM88qn0Zmi8LaOA2dAALVoX86bNxIvBTPyJUS6btXgwfO
A1jzl2kVfvsfbfir4D8YXNOLBS7QAMPpVd+RprsuS6RVxPlyZaitw3YR3d93
JcmCJlODGyuNo8AByfbiK6Ao6USdwqGTKUYxd/uZUDZ0BKMkUizy1YpOQkri
WbcC4rVYFTemWBkcQAo/bKC1DY2aYII+DzKP9uDSjE3YFagbn1VWHRMYtKbd
0jFbkKZo46dszd7rTSfvf4VXL1WI70iXgX/ytsIEXERNw2UpHi0Mgj/vQjkc
TgBrkHpgzVQlUoCpTkAJh9bizVOmgjVHL/evMyoeMXngDaKICud0pFbSt+TF
g4Gt+4yCs3cQ7RiM3IQ17hpE7+h3quSNYoP+lecDivss48Odajy1jsyOlHLc
RTn5Do+D2YdVXImijTuOtQzlSlHeTwaZAKx8doYurefhMmiq4UuX2VENgY9E
noZ94kU1X8UkrlNtuJpqLDV8Kg0IhgAUWblghuY0iZMgcAx5QHpsCEe/2HDW
iBDMVbWt1eJpiaNIZVPf3rh44lTvGMewtTVm6o92cFiBpY51et0fymqzTcAb
Rg5JI8A0umhUubL6qFdauVSGR7G6uiUwRnHN7VaNXq25iYaHginqyhJxK63s
GICAoQ+60KFdyu5Vd9L7i6bSz8X3SLs22/MI9xQGInyKybSwA8qUIUfNGk8o
/xYxIRAjs7fOK2IVM896hAADvLsGLZtAe2oAaaNSTHQQyPkmnnObUYInGsVS
f1Guu0i46JLX43Bzhc0cCf8wsOv/HT9Y7oWYr/uIU+plI2QkTUrQ0cX8Wo48
AMHJ53a+7m6uQ1EkjDOwSCqLU8VM8MGYZqAOlzdydTLZz1ot6sv6n3iV/Q35
uJwefy8Uu9640JnJb5tyy9bD8Jj3aw5tWff+3YrYRrOUF8rN1Las45dORetg
9wa9+Ye/ihTPH3nF5tbP+hKbVCTmOSuTXIPznEZ/ULeoiTw8gCDe/5+ZjDyQ
aPdUfPvw4g7CmmiDJyc5CyFEc3wqAgRIe00auRJ9OJxT4AL0dMa/EJd21jdh
HC5vZCExSvaLEcq1ecyVHgmWICSS9A/H+D/itdlbvlFbnfm7NknQYmPNuv7v
jQ6es4lOIKjy+S9eAWjxEsRgdvnuZDSAv4if3yuu6m+Cusgey93o57gbfUno
5ChPVjvA4al8tE6AYkpZVN57dAu/bhh/GU1m+XUGtaK6R2w/wqaIE9rz6KHC
na+ZsFr2qm45vaOTJ9cnOyBbQijtkQU5ahguVr7WBQ7Cwqb1B/Jq19M27pLU
01RQwpi4SCx18XYMTwUINnjnNwlggBib/y9E3/HXQ8tduY9UuZfbW4S7fYlQ
8+bUVjhNxe+86G/RQ/fVUtPOwyGSBzy+tAEW6E6WbtfGQgRWV34JXSiPClVU
uyNdvvjcx2+8eXAcU1q6uq5mKv9RhjTCEx0R41s7ot9iwZc+NSfYpOgwSxvG
nOXsAmeUe7oBRZAy1TBVbwDQhZ88fZDR4eoX5CO0/S6KcZF3j5GRk27umPNc
PLud+XnJeIH/VGOZq5Rx5YVfdZWRL2xcCSIOn8aFfZvP4PAsI0+WhYXN2YoV
K5zDXXUxnu2o+zff1dbzJD9g/8WTS4B8vN3US0qyOudGkC/O7xNQzAsEvZ29
9ZHAgFIYcjLGGqRaYdA9Hma0IR5v61NXaliEX8YGT5BsRv4e1suprxK7ZW2K
xGI6dlGTZIOqtXzByrxGmzDt/DEDJ9CEmCL9KEuZGYDpQcpVI2FQxsXHgMf4
OV/1K2kNL3S9o7qpAa1ScGQVeQVTC8sLP2RfZFrp5xjihDa+ZX6Ibr4kzk19
9/XCniVHCXT1MXoc4lPpa/ho/a41GttfosR7cpYm25OHVpMxRXfg5VMWAPRc
665oeYSkkS14Zc0AotXnjXVb8w2FX0TFKRADsWxz01fdXH+OHf1JHPVAzE8t
Y+RF/SAzv0p5YOuK/LT9TS5gua3Wbj/zmd4WgE4dELBXQWbkSt3d3rTHPvp0
sl6bBoSSwSDReU1BTbAqeE13kZZsxVCgMYt/B0AC8uDBO/fGyqr8zhRbRSlG
VMsOe3QelTlEEm1DjaAmlfAsqKFq6it/2yKT4hN3eWgwbKF7F5onrA4IZ8cK
kU4ZStunl6vzAHS5UdNA6zB1Xi5nqr6lYbieGCK8AQnFxl96+OGRxkXKPrKi
ipLUbJrLgyllyPQ2z3rNMttfNYgb38mTdxwsk6jOlx4GkN31QR/P2AU82gqf
j2KnEQXqUDDTZ5xyjkB/7ix8Fp+/pFo16Qgq59A5o3jGapKhNVxMPETZQdng
PSKyuF57ODSokhVK4Ekckj9/jgEprtHGadTJxBitXGyJOYIIyhT/eO/iWxue
0o1CZbQTeRkEtDf/qYhpAKqsyklM1p/+a4Y0WBczdlEY/3xOivr55sGsVyTV
M4onT5BqnkK+MJMyrdWSsfL9jaYM7+QbXQ7jkIicFIvPVldgjeH6RjHNPLJo
kFQqe7uOBZRUj25sMxY7TC2NURKKqzFGnxoJGEJBfrHN/xCLS43o5V70IGMD
xYBAeo/hkCgiBJu+m6sZxEoEaYxIO4ypT22pheyYJyg71QRBaAdO/j2DWy8u
he8WREOgR9q2tKXFc6ERH0O/0ObCjTDBEZL8IXhxBAw4G7waHDHP8NmCz0IF
o39SBYsoYUUbfA+rymBAWRnXpnwVDZInEljLct4ZaTSaNurpETE7Mn56GL5T
iF6hzCF4BaiSuBeOrzn1X4gWqj5TJPDCv0E9bMVslz17usKiwP6RJRN9OfZW
Doym6zcvVQ0Dmqgx4Zo2tlZPQOarDUyxLJLF0XAa0dnccxaFHJJ85Q7T0TRX
AFEWe7NlxtqpQ3TAkZbHiHDGk7i756g6bHBUQQ4aine6koe0oan8F/7eRSP7
+5rFWsjWbIA6tpkjVT76zLq/VjLjUxsWPtDJ++Dt3z7yA7QbmsWA88SC7n+K
lRhjYZOenaLlQ7bUyC3yoS2dEKj0GUPI0xV7SAzSzE7jl5D7JRFUTkeXxqXP
8CmzrGxqPwxu3+Bor3waHC2fCWwbRYUjXBcEl8fJ1Yyzipf/ijP+IapXhFHP
tnVg+frEfzTX8rPF8BM4r3vbuEEQ0EbpQ/YaiuvlrZjYzIKHna31mKMOT/cQ
00D1t07wMddjYxZzWewnFrEjoMnQEYH6nN0qOZLYKl8JH4SfwXYHy0Cx2eZF
sMZ9gxzePI8dcjXMS77h5gO2HaMZL1g8kMiFlwOhppYS6nOakjklJz8iTuxt
EUDTmJn12WMpgfS2ZLBxFl0cpHXS8d1FHbfbtjCdy8jXX94XbRolrXpbE7KF
DCnV+A2fpxMtsVm4X1RT8+vBAS9PazDnqwFxtTKRpHdwUp/X7ItBvPB9PElE
jiwM7Qhz6/CwsTl+WMZaAjKxEuF3KG3V67qYAqFEoIIq4wu4xM4Ovar3iVIB
IHI2eXU11O8HvheZfvqcK116C2hJ3LHJ7GLclxKI2wWDI9BINBaupT7EEyDD
ZhbMqot6RSq1Z7y4T8yqVMO+69PyRqeRKt3k+mUEVzcOa3rzmPQXcegPvwBX
+WpQAVx5fkfyEUpSssZxS7ult9t2ZGymE5nkJP+Rnj4J3a6tpOTy+Vkmm/KQ
T9ynm/+YGcmNAsrwbLXxOahbQc1riuG6524p8qPfpbiT3M1Je9mp8Yyks+bh
cXL452oyasZE9ksqp9ZujdyT+w8XtXH4MK7WRDt2dUHVD7MaD5g75X9Qzuqt
JBCXGJpzGQTOxXfql4+EjqG9bAg/r5k+2kLn+pGC9t7kfLHBoHpA9iLiNI/j
eAaZbrWNik+kiniMgGIIDB1nY/zI/KBihXmOFp2J3WLAzYL2AiZevEYYdmf8
BisApCGA5+jM1lZqYQzsw1gPx8f6O6Z9411a6Anoa6mg7cmBagFtyu9Lldj4
TkBxj52nq+Ef8u0QbDW5Wpk9whaGkU017OvgPPiGbCvDotbjwaNjm/MMxsb7
A1iXMIJhdS1kcIZGSUZzH4MOw29U58CQDhbkhMenVgLznP7Aa4dLA9THwyvJ
z3I9kbdcANvNIsOP4UswUt36qNLvrnfzVriYXD87s1ARmTbsXHczxdSvntJQ
mH2h8Ef7LR8hUGZ1wqzvNxWeGDB4XDzB/eNV3ulNnp5FmiLJ7DKWHAWtiSUC
yKCQmcH+szzBVAkcWiL0QL5ZnUY5pSgvYUCQwkp/adjf2Jvhf7xeTGtA47Km
JqCc6R4pUoX9JrYh0ZbIQg0jLg3B32i80vp1NdoNdF6W9SzkBcpKFJKyhrMo
ygL7z4O0Rs/kGnt3rbHpuYCsp8MVUGkHRTUI7nXLf7scu+Brtse6mM6B/fqL
kngAnHFTvWOhluYOFlC6A01bDngQcD2AKu8mxDHE1He6aMdS3polF6JgaUVk
xMfMLA2DMxa1zMtocqnUnDnS7iLfLuTZOy263FdXCK5Qz+dsqq4oewDzQQpo
L+86emH793atmWp+ArVoKFGDztZuKvplKzJMXlXS1ZQCwxHru5YHQklbksfq
wqKqjB68BPydp2+eVNaQH3PxIBI05Y2Z0Ked8GdcuALV+EWyKZQWBv7AzXC2
8Rnt9wpAReEnwwHIQd4OEiOlOAkKQm9mp+jS3uL1VC8OY4+73sx3qn1qnqDE
Hj8N1WLJMqWA9U9kwvl34Ga/AD9DtvyVMP4+dGWPt4QBJkc6dsdPXckTYJ4+
iR9UnMnGlnl7BrseyLNPcPiVYPXZDbHuR0kmuMST/q4x5RNSlBfoA5KF3hCA
Y0wn5LJq43yoZrfsqeEAhvvvM5Dbz8A6SBo9DslTBKOc07gcczJk4iWQy2dM
OmbwzeIdAylQbZJdX5XOMj2nis6fBwzwOWTbWT7tJxjRQFfbPK4+8AhEmbjk
o3QEqbXysUCFdJPL93pfBpWqPX3Cflqf59tfPjG4p0HO21ucgeXgBSSOnsdZ
Oz74I4wh3B9XBCxm2Viz+DTVUiu0itRyRgGlDOhcfVUyvF5EGziWEfF+iDWd
QBp5goNFGW5ibCtSqmrOGov86jw+9x21+0nKWU3hnIILvPgCOb9pTpE1zLGf
5coNCT7Yn8hTZjSHVQ4cHuhILx2hY3qVUe72giJ+1P0OgZBeL1xBC0NRMntL
io87vwmIUGcO3EcbjDf+o1QU+Uh1R9WmJZI4Q8f1UJ1D+gzcGq7lD7vxmGtj
bU6qgi4TEwXj2ypXtUT+0COFjO3//H+qcHiKhHkZsJoezjkPj2+btV0d3fsB
qQbvuQ7Jo7qVhyNpYwdNXdXVuXJ0Auaqio4H15eznWq/CC2o1gDdJf5wHXFK
jZl0eenzkWl+533uyR1AUnAXSxJXO6Z5xYk+yaGt0+syJgbdJu9i2PUz2ORD
2ZD5YpLofd5xC+rmjiTSxdgub57ol5LhkccYynH9vyWBClXtlrOzxqIMiIms
jgzq/M13VRlycYyyxWgoMnYAkWOL0Dm2+ZETec5vJjEUqBB6/rNm0ZYCdxga
TctUNJhS7/V5zKXdkuCZ6fSfz6LmK+k2Os7bvFZzd5+wNGWlCcJZFHDa92vn
jxA9RxuV5v9jGyzBhOpDYEpKXrZKl4SmAzLlwnX1TSaZjmok0/AqgXRjfw4V
DJR0OaGFUuKeQIpVkaJcSY2aMEf3vxblR/iyzUvs4ddKBCNUhKuFqsFS1oVk
fO/z+02TMwiEBlZbJfivstJvafijOy/p6Znzqt9L/h4ipPQnXTI5vyuJAhjQ
AvMpRABfoi7Majz0DTVr4Eaci3tof3M4kUkavuAnCo8Gdg4+g1FmCpBvljht
g8ZrS26FCj6xz/mC+/5mBZupAIIo8fMpjlhd7q9I/QQ+6MfC8A/Q54TF1PgK
UGOZle60P1fr1b5lU6mMKpm9+A6TNGfTVssN+llUKNOoMX3P9zMVPkfLZYiJ
+HwQeNr/yeMExkcxjzduBFEhJtvzba3CzNoaQ+LoMXNotWBrIC2ERahDgdRT
x/oPe7c44pwQzNiregEASldSccQeLSCQbm/7ynSPspL4L+N6nntFvSmF+3Of
FFVqLiykeCsG78YkNJ2PJO4gGJZPSo0hybu3DSuhwAbL8hTeOlMj/yCKGT06
knfQYkcimR3g/4enzDozP5CBbWEmgSgw6DC5HxKawG5vNs5jylZ0H3anuF9d
p0FitRrf5vGchU9RLs+rgcFe+xpWNPTPNp2vUCxHiTAKSnmYJrEz4DuhbHgl
/rQ95l73ZxgdlrF+7CpcYjoCSO5JF96RAcsmE+3cMvAq9JYfqc0Uw3n6uiA6
RyiQiavLeAxZRVkoge+1SX9i98f4NCSH23KlZeO/b5rpAbAiHFwBRf9OkUqd
zCR91p2HzGeeGEYzkXz/+iJamUrS1WNZ4GePbVsiSOEeRzDOS2lsipEPLvgb
cYe+lw4LjzefGXqfB7PnXZgzr3zlbMPM1vi28YQL8clHuTXG/rYcr4lfYZpy
1iWgzBmZkX3+bopwo8k8AOb6vF1Z4WwVc0VvbB3J/uXO+LlKfM1GzmMSpA6y
YYHRm+ErI8P46Ai+bEaPlx4NrZpSLf1/BxFeJ2cEJnPTty4oQ+cbIue6Gs/B
6nIn2FENSHfFpmMKF/otWpQ8iWJgTwZLM5L20eN7LzgbEGNTWXbf6fqQtZFr
/QQ518LZlxwYziMZe7ng0CysAd1tS/7FQ6QmFAKYZ+RXs/2WVjVkWnoNHO4D
bpHWUo2wW3aCBb0w1AUt8fU8ycKAquJ0xZRBgXToWyQZYposu87MEsvhB6JE
2KYjlaNXm/QCbRxxmDPUK2Yniu1U9jwMf9VreoyyqgzWruosC58D8VOQedqs
Ze6TipkhhhlA5FctjKCVMXXJVOnaz0PmRScsaSpHI7rimtMfkZz+kc4X/Myu
ErxVNXgNC8JFo8Db/MoskXPM6pCbRhdKSY/YyVXC6f6bvN3/JpTEtmFoS9jF
3wEq/MjgKB0imB6aIAVt1xehoiLVoJWqy3yznss2FW/iSstcs21ibuzR5Vex
V2Sc+yJp1KGqNpLdGuHdHwgydsZNa2g6j0yYJUXQ5IYq1lt862qclz30qWN+
/1wGij2vSUFD8xE7Xq5mNAigL7hykpJY9f6hO5sA83Pxa9hEOWTDFPVIX5rk
cB7Q5LzdMCxi2soww+K5izOpkX5ctu7o+/Me5/o76b5ZSZsQORbfuYHxCqFl
KwJAMpF4Qx2Mi2WXZ19x5g1TH/xBV+E0+j15Vg9UV99+lgR1xqnli64YCj2s
Hdxq6aConm/7Nh8U2FrwrEBJMHDrXPN75qEUl06vkk6MJpnoyp1g9tFKQO5h
ec99JpijIYEW+/ELto2x1EvvzHOralOvaKa2hvZrqQEOBlWzcUYP6ZT+AzK/
JVsQzywsZ0UdbO9OYJIPskKixSV5bOOhCxUWCFYKUBWYFHgExcxE283E1wq2
0XNM9H3fb4dDBs3DsqWd3YqwSUjTeBtF8SAHkzzD81khrOiiAdqKKsEnRF17
pydJ/gsTS3fjUK2Ow0N1oZI3psqrWgBpuOG0gMjTdMTdrKyA1IlirpY2ZBde
tvhv+XCP3kc2YSP8/XyBoYpUZCs3ejkBfVQDwQt/vL25B5KWGNoR0GqA350c
XgSr5g3/l6xtVYvPLPpXlDHJF8SEmTa65NkGU6tgcPJUS0OwVhhKflGALl/h
42EfZ7gXp9ChlSxTPSUbftDvMXBn5Uj1cfteIKRFhbJ37mto+TX3glrGPvUM
TLmgQJtk+4nlFNNpPPfd9HCsUsCLbcZvxDZRstKd1h9hHf40UveOmCWo+P8J
fHTjmDiWWyHJ01pvHXCCvv+YdMbCNwxhqLfuBQq3OAtnWQ/m/c3XHhWdzwmj
ZryefqEH5dPs+uDTLP5pOtNxd31nhBRY4zvgRyXdIooaNxiHRptB4Lzrhi6w
oBDaOGwWCunJYWCRDKIYi17lZv2A172e/6P8OEjL9GnT64HSRCTnT6K9iWc/
E7X26xO47USbwKrBaCj/UKXXeE2V1GxwX2DHi43gjQcnN3qa/o4vmDPXdKTK
EqoLpKwcpASm0pvj6bB6p+c8UxpgTZIgB/CBRHOWVkB9iLgU+yH+brEPMGjN
3A/bsYeANUZKtnB+gi2qqKJPexfMBTMBq9Ju7QkkbJy0SUsZLA8QmafxYSSu
bvpD90ckSU6iyungmilSRRDpmTkCXggA4u/OT+gSLfG45CD9g1Bn3ICTd/HP
wGAAdSBTz27j3A/DwNkzM+njL7ktCnAK9t9K/9LwilVQkr0w5WkMlnBxDSwl
QSfy+yrJkWAK2A0ohqqJNZ8+0MjZZmduqy5kUVVZqJwCP2pnKF/qI3PNnKY3
iCJpNA1bNGxtjgBdXe8nzMz+q4C4qnQv1Pq4FeGrJCJm0LihyHiXSJo0uniC
+8bmdb7pkDgnVWRQM3YJNs26tjh3drQyOrFLNIDcYWsnTDqH78IkFp0Ug07Y
m6/uFZZYx9HdaAEkifElBjy326fK41wFlckwLPEb1SKkdkmYhW3iMTo/OUiV
uYnPnb7Ov28x8Q8gH1W/VfI3T2Z4BjBN1hH4jBrXQbX4y6/4iy+eh64U+wd8
qIWJ5Cbq2xJDDLSuT2//vaJ9ALj943h5kOsny8UezUSC1cyYx86V24ZDiuX8
ka0JZgN53RVz8SD5JAN9ash9QpzUwpN35+57y8KlGDvzF54QUKXGDYhJzUAS
yKvz37lDxKh9mhcs7alnqYBXcvDtjZJAAfgwG+2UCbr6WGKFMjHJKmwMbJ/6
7lIVzzGkNYmFA9488Ko6JWUysDZ3s3r0fTl17XqY7gwzcnWOlzv0AHUOJ+5U
wmJ/ap3ob6HAslPj2M04I717XLWHSsg6sAOYqy002Adu1ktrVGHXA2gUFWUI
uAocj/z/M+07qSis3U3KkN8TPlpRZpZJrsjXoo2rWX6HrkmLaYFPjExtEbEG
T0y8fFZWhBhy8ahJlJp45ZqqRsCRmljIu79Vkc/ogsWe3mUslsEMXz8hPLla
LHHjoGk1fk23oElSnts1AtCqi1XGherwX08zPPCOLuVFlG0oP7ZlRBVvv6YI
S28MUlmnzhRe4RHmr3YPUAINIyF1+4gH0hZAo2fSLDnzn9pL/obc0A8a4bnX
lzOfePnZ+ydB6zR7nuBTu7bUmx1acEolCXo+zpmpO9z4caDzexGygyWtqrEs
bfoj/F8Xkxvps/1Mbi0haa5Uu4t584fhIk6YL8KrC89HHHxSYZEaIc8jdb1Y
LEwdQGMbTPSzyHxqJwmuN2J6zUaMQ47HmlMZGzl0g3Elx7rinfIwKqhVfuk1
cxZVj9tNeVvzFTGS1Ymraajq5tc8arNrBCRwQPNg58ouNOOVgcTgpQY5IWaX
IGEnf1JYohKhx9nntijiH/gmedDXul8BjIyGX29UFm/0DKsBrht7i4KaJ+i2
RT4YONzNKZuPKpQjiJwAo/Zh3Z3eJDqsBLTODrfLleeGphoxu1G9rxLMDhf9
iJ3lC9mn6breMMz55pzDjEy8pvolgv7zhr6ywa7EeNsZEJNFh8EwQiKnYUJP
s9exqnjojMDmb746rNFHJdRPyXTfzPCK1PIbzSfb7FoSQmoZP9n8zbHgMXg+
+simHYctIt09lwER2iOHDywJley5jhLKZsBAFCXUC7niFc5LKoABF7v+BqZ+
E8aSRhQsU2TMFomA9ZXuffEisENBe2oUJkucwGljuAXwmAgxFpaisGL0kDnI
zvBJ3IlZtPRtb8ibE8rxYQlYqxs5/q668WsGRJ/NZPiwz8ZfYDpGCAExNrgP
WHCy7se9ihnJf0tsAcX2yxBwAyKDGpARwGFP0pM/A+DEFT4I0rdc0QrUs5Jz
oDAm3iG3XpMzawyhFyDwKU5Cuk/U2qBGJa3ET6OqcVaH6u7C2TIy7I07IyOI
lWmszG3vknQNtGbXKzTC9K04+ZjXCng/SwITCeZ6fR83EDYiARBnuiRJk1K7
2738S+d6M0jUEKdVEMqGppRoXeOTl+dfUApLqOCTsX2FEVvqjgPWDZbyRegR
Lol12119WysTg3fLMuyDQ6Dp+89NIkWfyVOmLTLVS021iI9PHHc9laR1sBhx
QteHVmE7VYpmcF4wrU06n8A6PbkRGWsAaiZpRQxtzlbDBWONBTY9t4fZe245
WBfVLZBEl3rW+VrnXNBWCzlEw+zUvfq5kyguP8yFWRoSNg9yBacoBTmK1EaO
DrfrMbcGy7HsygrehNB1U1NiPkDrGshfv0eXqO9KUgu36ipt6WuYuj60uocQ
WbXbuXf50iQKu3H2ANP0u6Y72vvioLqs8JqffmEoppU3u5fC60YVCLthpA34
eXwi5xuik9yBHwXdbzS4rlewVEwKhDnFprt5cLJ6+t03KE2P09xSW6MkvRk/
87wT7XukWcT6Qwe9zACsD8c3Vh7/9wiLA58OzQ6gDJErF89SW75DC8pPuzmb
4kVzdsdsKCEQkprGFo2qA8elIcoKiHGssu3oTX4Wq+hF4/FycoT+S/UKmNBx
ypYPp5g/oS/CWXaTPFBbBQwNivtrlUCwiw4mJwqn/DJsq+ZD4g94KU4Lk0U2
RMoYdEUkeEB+Ch9zv1PyxjTXeRevK51/8bOIAAv8uApdiY/zkzo0fYmKhnHI
nrOTnEOii76A3B7Q6c4PTiDZZ8Hv3Pt+4hCE7nQvtjfiTObVbUq6t37zl8eR
v8BuXt811mMImJlHC5R8fjxkYOVIAef+W55Jl/nfQAU/IrwpUJkdQCizrXIo
yF6fSVeb3A37f2+j6Tf2KwzcuzZVKODQhnf5rjDew9yaroJOqK26OPEvNnSf
oTVkPKNzaghRXu2h5vZ2kOwZ0KFlGwSuycqHiIug7p9d/q7TkSsIdS0o0LEI
iubl/DBE9q5HaW/0W4az8atmYUmOdQPAS8jvn1k0lFfs+qg7/SH0BNNF/QjR
vlOmK+BINuQ8Nc4vRyTUnbaL3I4Q0aSlMoaAoqofG9wxfPD/Utw1jKGidVVQ
1mAwc2p8BP9+z/duJBJzH9eZ37S5jYQ3JzF2qGKyTF5xqGDrDEDPHnChKCKF
n6D//uLAkRbJOZdJK2sX6HJTUJIjh9xc9Ru9sgNwAMZKaouJpzmZKYxsj6Kh
BmXxwtsrzY0A18qWUmrubIhaIlikYn2IG//m3NpCmc2ouk9P29lWEZcSLbRy
5LEx/nLIkGOCPHeX6T699gntGCh3r3fHJnP2TAETAAjgAEH699mHpiy7zz4n
3a3cw8mIVjGujHsi1zQH6KL1xiFestAu4tjykoFFyLR3K769JQfrb1Mya44j
cBgwQOYObPRA+rYOZjzCe85V/IiJsiyzkVZe9fZfOxLYTiv0iLBaBf3YaRsD
soQNOnNxg6oHSRyZoSYrjYVHxtHDf3k6kVCWVjVsEwngYDITaFiY9toq1ynM
xrRpys54rWZsPK+bm6W3lmGJF/ylmmwxpOhaSZp2N9dpmpvE23pwp05EhX+k
mbSu5W6SouK5O8xWgSL1tkphq8b+hHsyhkYpV2OYvf9Rp+10Vd3RwCze08sP
ntWk/AIawjkwivnLhsRapQIFRb803WX6IOShBrUoVL+oYvvSw3WXaENbFQw1
fkk34zKpP3LSAELbb94W4m6xXhbAWB7Ldvasl/5aR5rwpMr0PuOH67ktr/fo
nGRWbfPOXea4DZovOZ929NpkfCr2UkxTvV+CfTTNoTK/TCAFTkWWNpeNRG8R
4QjXcfU5o86D/frVU/d990/c3fjCxjvVn8EGNc6w+/EnWfydt+uPHL4g0uin
ulXN73Zji1SRfe+JPhBUzjs9he/4D063piiWRrgb/weXngRpGi1mO8GNFUHd
i/188PLULfPhw/ZDUHd69cKi82YcEVLnk7NAentZVLK4em4/BczgC25FXXFu
qjAkANWx5gtdTF/0P/wiA9DKfs8zkBc7ya8umCEhqGCYoS/WVGT1FPraLgUO
R0IKWfub4jcmy8kLDjCLxZxXNxlWqjUFJCOAAoeWaaBdFm4hMMGg/90+ENyd
DPG441Ka6rnIkrTWQDkQa19wLLtpMHIn/UYn8wIN0Ty4Vzv34c5T8IjA4FEX
UDOqQRharbpdAopqNkGvIcLIdh9vXvzFhYf9Et2d7EPzZ69YeX2JVA4gJ1zF
6B6aunFWdSlFEmUWPH3WZAn/scxFGJDNeDH069WGw78uXHemLusTl9NHF00V
dxrVvZCImI7zugZO5jXZuB0NKo74RArR04zTTZOWpCVaFhdpUQp1uZ8Szx2U
Ei0mGSqbVr+qEzUX6mGssUiuXkmOCEQky8Oql3PEcC8MsniL1Cb4LlUlrUue
oJTuvcGDThhku02Xs95wEsk+QUJPHPMmXblRMTNXSNd0AEuQB4p0Q1VLIG5I
/xC+CtCIpziXmZzZpyJBtmmlrQpVkSmlKuc566Sb3honboWdSpMCYte/EgSH
oRqg0llGGq1uY68Ye0bJo38VtVQxkdTnh6ir7e8wjaSZBn8LADsN4bYrzSmR
DwtNjmOTvqIQBiWxyKUUEcizaDZn7BZ2SFQbie8rCT+0pxyH36YLT9a4p4Lf
eHDQAwZwHxoTErp5DI6KjfU4ycomfpL6Gt84oLHVg7wlQ1jg9wJs8zfkpVo0
FLVFhweMa+jr4EPGX3qxvoldbKbvLIHLQ7mJulEqjERvXYNhZSgMql+QpYLu
K4PPruxWsWpJ6Gusc+hQ/Q/G0Se8KZAGcWGHjhncH4KQ004u9iBbecb7j32Y
GqyTK/61141jFV9u9SyJqTCi0nBSeon+91O/LlsGzNt0S7tfSlhbiWHIwwJq
VA/49WBHsvY0n6jlpO7BIbbiC/fdg8rwC/Dkbx3lkEkoSWhXVfp7mD0jlOGQ
KNBxKnY1Rs96hR6BC/SPz2cjstIIecs+PivRO4UpxT06T5OaZ2Jw2+h9fADc
fY8XyTNst08z7ZkaY68e4ISba5oEOmOqnPiMDTDaD6nqrPXfdxfk9L4BPSeH
0LluAP8p+5ZfU5wjPhuzW0gNOB5u/vXHzxfgJphl1VaBhTWtKcFEb5F/jbky
56BfVZLymAz05SbfUV8y3g8DvoiWz4Tg7W7HwkzzzrAm/fxDu6pP9jKmLw85
I8n11f6SbUzQpDwKFseAYA3Mr3EfDmNP5MW9i4hssPn6ECyrojt5myyhSQMK
yIFKw9MfssasxMEkmeyc/p2iwz3CItPznZ/9k3hdXGkoqiGvZxnuxSUaCN0B
wNpLQsqCovbbyNshWaYUAu1c2EvP2uf3Z9JWGJo7r3HZch6PC+DijcfsgLgr
KR9QR1VGtwZBY3UhLf44/IacxnIFSt0+aLSNVa7X3BEpwyxlbs58Yc774Z4+
ccFVfLFVWvmCHc7j1wlE/hw6gupElA8jQQFLg3HvVy88LmEZ4g2xc/FkTngR
g0Kf11RtYRdTipKIbho/mDS/QERQGZXut45/UJsJiF2Odc/Nl7C7HwDgcAKo
9mWZ8BixAoPkYtK1LpNAe2Xlx2f4DpHdMZ6dVcBYzFTYs5F5Iqv2g00VloQf
gfsaGS/sxgG37YUlnE7ZdyIe3p8mrfXomKmN0mOtFGCzCiffpear1paF1Ln+
gRhh9Z0arx7J6fX1MwJJSRldbNQY/WyQbhSb5btJxTCXLGgA2le1/Gstesr6
pmV1/RrBHd29MiEV8503vE8Gx+dKLh8v5Jw9fwTK++Q9MtHnwS/DSH2nqIHZ
bE9zV7JfBE5WplVWRel0meZUwN8l46lGRvK8nnAMZsob7k1Ke86oNeHieV8N
5Wdux074N47fv2CBSIErej4+Yvc6t3zAJbXs/7jIyHHXsFKpellt0lSwLY5M
cgUwz1wCNY2KxHBARaeKX9Jev1VTNkXQMI8oaG3gTJ/hlhd+8N9mzCKrYAiG
HQ6CTweYx54BIkWPRS5iYEQm9jcaXu9iGPIgfyOgLRhiVuvb3hyd3NJQQymu
IIzCcDG8OeRDbUPWiAAdPNhFfUZVmC85OgrTIGbq4FQQSZXfO7t4AfSSkbwO
BpjDCNJEptnVYUofJvATnnAth84vRpJybmoNX08ydwqjJ23hJhH/dIYTWJ/9
kU4vOdaXWcTNs67UUjhonKdxB+iog9wWCe3ltmsPjXsUrhGKYwmBzkzReRCC
b7ejb4h6AHDjlrXDxE3dAbhfoupQBL9FzCtF+u41G/CNnhzGO7nuR1JEBUtx
76h/Y27WzyJgpnokAAYNB6BRP04MMQksWhkwo+8lTpIzZ0vvsqKdtVU5BAPr
akO1URp/mWo0ICzVxELF5Nt93Ux0JzGw8/VXUM6/M1ehFkjdWB32aBW2P7MB
YQCRl96AGe1ymzeebm3ImLvdwsC/7zU1UUgWVUalLVfNk3gh3mFtGaYOhwtG
13fuW3/5YDqZ3O38lkSGdUOQkcYZmFbH7cEz7tRXpZFkNaJRS6VWMqB7x1Ty
k/2g7ntfyDroVh38APXK/dw/FE5fMCPKvUWDFOU/UtfdIMOfzhyVip/0HE/0
v0fQkY1EqDxm2IvGl1yWo38WEzfdgNu1DU96AFIHgWDOlOiK/08Jq3NSLW5U
706Wgzgu/q+QHqFXG70v2NA8tfIpr/mdFnZwNgCm0+DPDyBlbfak7PcVG7dv
Be7RzKGkT+5SFKElUuHvMwNGOE7wQPuji2US4jw7PVrLUEuo7QQNANRCtah3
qE4lQ2WiSp6zXvzdy91uy9t0IO5gfh5S9KzCsx3rr1Kr8NCussNjiwCzyebE
jhqSgvQP52BijwAhoN4PaXY04+xoT5G96etTZVKMwoMAB8dY+Pvc6gW0uZMf
m4xahu5j4XUVeCZdXnJhz409OTJ2k4KHSm81vdcCcjl5UMfx1T4jsFspHvyp
vmj7+qYXqjq6g59U9gsAVSZ9jYjCCrs7h9wOEZPDxuE5aIYf9PnpTUbTAlhk
BKaTJ5x13tfi7TZwz68IkM5yZYNVq2zNVCQFdJhId5O6S0EZjAUIPGSc/NoM
Egp8iIjtJSufh94Za8uatc5cEaRPTnXWj82IGvXLqVQa83Gi42HZcEZ2S/Al
ih/9krCFj2vZ8Y0OSk+8Wa1SNOeokjx0zE819rvhbyOw6G9iS6vARUURXKjK
LMyeGsTX5dCoGveaZcAaOWr9OEj+GbLTGoqzL9Z48KgKw61mdhG/6/i5Fhke
4iwaVHTxdaT640rsJgELbG3WJ94EpZiydCdH1DtwShFbyN0P35jG6HKUijkV
xSL3AURYas1bK1OEuH8mgJBInOCpwRY6Xe/wK8Uyvtq24CnDf04nJNL3kzjc
aJYiGEB1FQOQs4UUfpET1Y1dJH8/X7MlV2p1X0bOLot66kDbFNgR6qkEKMvM
Ose62C6XXN71IDKymgP5HCAGqHLgPl15O4zeph5YM7wTsOoIQsr+bM8WU0vn
a+MUUvZuBseFI/79EK0G9sgUFEDOBzWO/uUORaNctHMzKcTJgGjc0NDkqGyW
y0nWEKQb6pH4AZ/yJQ2ei4LXAvEAlxKYP7znOYSSUWAhYlzU1UDkHIbvoqrb
EB2DlKPsai5qGljGm+W+E4kKvohmQojJGpH/7SQq7Ca/iZyz1mDqeoLonloT
7kDTtYJRkr0TUx6w2UXIXyD5JCqFKxC/DjIM/+NNgjsX7ZoByeK6XF/3t8BH
hhW9iK+BKXHql5flQtfsR3uNH2nWaI9L5s7HNFL/X8lpyThp9QScDvHGq3bq
pUba3gLkVH33Kb5m6hXa3UwS1/0umCiBGM35J5ot5r1Kx52nf5mUekmKwUz1
CtOTzFSJUbKLnD1NiN3lA4t/7+yqaf2tQV9YYAuqe7k6rUVXlZnsWa23c68e
/oPzB+xrshLJLRtZlkVkD19FMb4hUDeRpz7XItFAzGMKB4IUFY5cFoqpqLwa
FzkMwRcf3CsJSSALhZNwB4ARIYJPbuKmvA7xtAelKufK3GRUXyY/8/1MT0TJ
XU76C04KAaEzcVesPKVGFX9rpOpmLET2GlzSXtmgY/BNgwrwyEzELtHWmtCt
lDs0zRziBOejMS/0EwcCY70/Wttk5+Z1yYyexCoK6pA9oAyacbN5Q4U7SeZI
Nb37dQDi0bQQHzoaXrOJqHAfP1r0qsDc9h8Vb3iUd2PQWbKQxH1eBUmoMfPv
9l0pHK4yuPimhf0XGpTFP9ZBVXN8B73qlYbJRr6uU7ExgBHn1hmGiwjLk79A
5JzPlUWILX4im6OsddKQprxf175DKtivGqB5GQEQrihD3c1AvnWNX8SeUxZ5
S/r7rtQhP6fx3MRgYqheQnwEh3g81WpF4nT8nMlhkw2JivRulFsIOfqmjRXE
ZTGEXPcJwAfCoeWu+ZqoAsarFlzVVae5+ecKPtT4SuNquGYNzEINVra29wd8
c8mOKybzxQyiSkAGh4KXUJnkZ5j4mROExFbZMWyktSewtSFXjifjTg24BsdK
ZLeZQjXgJSDz9C9B894Z202JLkmN2v/FNY8w6d+/qZbnKTLvm7nT7ylGwvoB
3txZS6cRSWbz+wlGboT9FF2Hpa12ELszV3eK0asC3EJhRju6DeDa5UzzOTl7
EeNhOfLRYvo/akQWvEzOg1vn/u4ALUdpnXQPs3eYa8gA0eB57BDKhwBERdqz
M2/Ru/naeF50UYiYS7I7zqQypVdaMwOl9oNOZ7dn80pNBH5Sm88mlZJ2jISw
XXvfzXoktvuHm958kgqA+y4FoawdziTCtT+JPUFGBHq1sFuBIOKScznl2fpQ
15F0pJ8b8kwIQmc3B67tZ8SoFV2f3+lz5ykphuGCJi0YLLq674SdJMHc1pGI
GIaUHzYYc4+iaDjingw5E/TObpobZPhkGs4qsW6E+4Ha7lX5a7PySr4a58k5
1Z1BPXthOsuO2pu+hZqWddX6PNWBwqm/BDKB0SZSCYBmB8qt6o6yGt0Cv7Zg
uYkR36BLVGJj8KtMfqlsWPHpOGoQECLzHyUNAm2EsN8msiUpRKdBfqfJjaw9
pkBKh9rTFV6qa9sWmRafiL3RRVMDJk8NJ5fvJ5PYXLzpaG86M972OuIhTITf
CiDIWMYcxyDT2LgzVcELlrJY3k3lPhLMFkqEueYxyfO28qVSEo1mKIJU55UF
MO03gHbct6kSUw7AMKItyqn9v5aAdYGR44tYrQmRlIEKFgt3GIQkf7DziQvD
aljooOBHcYulDBNDyL6UY28hQYj853E3jwAOnKtssnjtRKfb/cqokzPkgqXf
UDIbu8SIXmhkQT/x7T8QTrp1C6aq/vtxK2eqJHn8HdGhaMYx8fWso3VXzTUM
9dG08/P5O6ZY3uTQEXMBFdcHa0UkE+YJyq3sEhUCNW0NwY/9a6sgwwJLnoCc
KXMCgUBV8vJbif8ks3MNZ3IN9mRPWSFEahzRDZWumqSiNqrAssB+3nt/Od+C
Wapyh+++nqTPwHOB8KazXpa/FoZm2h9uhSIBxUyPGtYiWX8PvWxrrGHAOs18
MQnC5Qnz7gJzTKpBplUVxMswaRHX94cmw6jfEJ92S6l+y9GllYCfXcNU0lbd
hsLYIbJQQ6jeDdHL+H1bPIpk01jtllEkR/YyM9eniMKi7O3f+Xaz1Q3aJQLt
kzTLuCOlIhLtGDnFk79bwB8oFvGCmYmDjZoc27/v8HanjsMk8BfOQJpcR9cW
D4SAEK2ElCc3tuvUzMnjOlWxsW5BOya/LTISCXQtu1o1aS6gVhQv+g/PpdJR
yZY5o7kHHnF56CNQvqKVARWHn5WK8YCf5LrrEWZmaNtQTZ8fPAoW5rtSomvQ
1u/qW3CQE1rH82CxUieQojD98S2qEjTKtWfXK77hEeAQLhqj1fO+KkHg9GHe
UyJBqkB7FdcpJfxHj0mRLOsKkd3i9xnV7zhFMwa8EcWp9TRJIAdwayMYnHNN
osBf7gLeIY7v0xh7oGLo0/LeNqXaEgrwDifJfL7/eZm+N10psaUGKSyFJGik
TB9NM1SujSeB+vXGZ5bvqM6MjEkfmZ227a5WdF9uVe795SaaG9MR66NlyS13
c8qmi6koEDpkO5uJwQ/Ohkntoy3bh+sW7Bzs/pKzoFAjg8LI8ray3oItQv99
8yciiOeHBAdu+JzxxmYlI592cswr/PezQnprz0PrZBWVSKsXKTZgGy3IdT6c
AtuLtRv0BA02KwMZ3F1JXQsVFg1zeYiFkJVEzx2aZjd/SyeNXSRPTr/CxdHp
RHp9mYQpUgt+eSjVtEFdtrtR69W/QlQy1qg3n/zzEhWRioxVa1tSDn0lqLlw
ii0BFbPyrmMwuigjzJKhoCeIzOg/7mSnBoD6aMJfLoa4mop/EzmeCP6DLu96
oGX7yrfLakqlLwfBvk73XXpMvzNk8Zps6WwJFqtPeWZop405mXD+VcLcXQWV
BIa4PDMvoHhPR00PpUH9t/0m1LOCMJ7XBkgkpo9r+G40Kw/KBHtD8hMD4yf4
6gJ5U4F2nPwa7tiwqyQ2cIzzA8guhrQcuvIRB9HacuoYFMA4SRHEoax03XLp
Uf7GFDbkOwZuRzsgjd/1BUTgGuk2PHpgS5EMYKBO/o9NH09lkMgJL7U4Ovpc
PSazuN84OCwvwj8pVIH8f5qaDsw+a2VD4ua8KaSU5STmP+acn8aL0fDrbEEi
xGveCfnmTZomiRNLefJGrlOGf6urj38HzYrDXSgPzZg3NZUmzyC6IL1YVgO+
w9WpsqyheSyvUz51sZEgxcKuZjVTreLQxxCC77sh6JooNsvmP/B37HK9/Kmw
EeonK/O5Nyiz3J7jADK7CQersOnXAXQvajKYzPNTZHA6JvMlUhlwiaV9sJKK
0svrPFBPSv70dprWi0E0sfXO75N7wCUZ1zxwdrsFiiGPrnIAmr8ed3tL3jPO
xd2P+DHPamxPihlkC5a2ZkmfKx/0ecJ8L8KszEgRXbV0vrZo4mNdyyWVP7wk
MhE4JO4DBTO9wjEsukMHBpfhB7a3s3joYt7waM0UKD4mOtqjhiI6q4mmb91I
wJA5/Q5AJ6158lqmA6VThj7o7+jgmQcE4/FKWWiG59tr7Vbdah07G+RBhuUf
CFAiJu93LsnBzTn85SY0pAlR5tB/1CwCo8GuFSD32VC6JAOLQzKTgEnHXO5c
tZdyj2wkh/8NxAm12IS1kCxrKcGmAcD3BM4wUHfwCVeyTO+Vf+x3+gKfy2W0
J4x6qZGr51823XBydjLj3ipgvtvg9beO4hokCwHD2F0UiSbUCu076+joQoAM
YAr68Hjzk895Wj0grVEmA7TR1bdrrH/nChsZRqGRcEi7hQ3NUIpBcqIEYd2p
KBXxVil0bQZ93acdYmsTkPAXogF1bEOgFquUaSKuuPpcwr8s8wTTBoTOn35E
LjvKEmSwasHpkC+s0LiKiM2L/Qh3Duet2jaMOplhJBDmeEL9JDSzmHB7AuZW
O62bUAmrDqcvjzj198UeT/6HJwMKnujo0HaQHBrjPJMFR+AEJqI0lDwQfr9/
KKK2iHFfwTCm3fNPRsasCm91xdF6UyjAsnHeQs2e2z0qLGx72+mujBK3ynZz
jWJgEjOEiFfnGPmGEZ5wZEdb9XS3SNorEhTc2dDtn0hUt57zAPJnVqnoe56D
E761H7ydPEsr0VZwTn5HI/CLXE4NxVfxW7ki+13WQRBLtgHrltplRJZypbzv
eUDPIM5TbQQln2URoUAvBQTwel5goq4hllY8wZVUfZpGxgRKGtPrUyLlj1ay
A0ejnzHZORw4mslgQDtIU+/ytUYRGw2811JRe/+AW+ciJTWAHvFT/xM0xjvK
I8EweOU8GrzYu/VdwFwnxLGDxBpvKvYQKmj+yXbdSZknav/PZ+vRvbtM6501
tonRN3L8X6BgjRylB62Fz5HcL3Vre0s9josnWtm5dl2MNcpz/bw12D5pGB+O
uj9EZeq0XcuN3RKkSCvoOGUhrOavi3HfEEHQULjN0/3pmOVUXvkoM7c92F7C
3xdSM4eYX45KyhoEiMJAs0Z1tsj1om7QjLTUMLiUwNfx+Q/LljMobMcufLNH
sRzDdu1+U1zxVLmrZpI1SX/DWJxwjJdADBg1Me9w+F6BRYCN1APUkuthtzqZ
4e39bVV/xUmkbYT3jiBnO8aSbcOMk2J7vVamTnnkOzPUz5VNGvw9+VEDgizw
HCUX4TQ6EkZjG3hN4MmKZb5lAmqZkxdUsSCtzrVb0LV7w/k1b4Q7TL2Wz9Dp
eQ4P5CLxE2RY3t1eImqtZ/AYuyRd1ufer/feur+PW6kQYgN7hBRYVWHHglJo
5u4N3UtE24l/C0w160dpaY1ok7k66909u5mjxdeVAbmR2BjizT7SeiXpKTEK
kRT75ftLKHxgx083ysuEteiGQgDenUKFPLpFmUepIlvlXc+97QM+Oti3rvi9
50OYUg4FtZpXoyQFbXq/tYn4rUHhOF+TuDLnR27c1ZwFXuyZgeICuW8GpQRq
pgxOJIkYj/cdF4r58Uxpazol8qCFja+nDLUCx93ebmkDsQ55Vc8rVMfdHZFu
WQ3lytHM3mcKkeAkWcEy2q33bWTeQfJvq3u0c2MC7dDU5ipIkHml+HqPmypm
LS1pTcayMBdon5MVhI9wHKIkdH9zvvvzmnIU8F5cjZ94VSNqkS6I+VzYUMx2
OIEfuJWxypu8N3yBYKeIgDRTBIHT7eNlyOxlWzqIv9pXCyfiAam+sPX0Vo9d
dNqdjCHbLhpLVo0KeO1q909lB+J2m1Yo069/znjLzqbkzEOwgpEAyJ7Dacjh
haMFKrqwGRyJGIH/iUusd8g2dUszFwUoHL02n99aWZwHrw6AwHnpejg3+cVd
xvWACGfMNw4+UzNO0ttX1b54YhORq5fbhgATGVt42elABwH/1qaZ5MKPs1oK
ReUqG/F+mZOYNOZODQ89QDklXQBtTXoWNvPbi6Mf+sgg2v4jEu0ojUAfCtZk
H1h42hWcUO90YFaLHRuFZTYNat7WGbazR8f9XzVBmwXD5hxs+nqb27nLLxNS
zDyAuEuAmNK8d/iehXZA2iM8CfO6YRw+tgPuzPNvdMBRW5p5VKKS/LOzvNwM
1oJTGBusjRZvwBhIFSZ17INM0mWZfd7CS9saUcaPCgKd0V7hro6Q6h5k3G0Y
1rJl2uKADsRs2tDHL3nBzKk7W3agRSKbF4NE4iN+2rNwhL1xsKJu5AbOmjof
hZv4UbFI2vc8SPXVP3yzISJjZpPXe3avzx12uJ4FxthcuN8VyrYZJM6uKq5i
lhhXsizFrWFZAjJflsJh6c1Xya6AuMBbOCdN1yR6oWI+1Q8BeRGXPR/yNxOh
tozJDAxbtoqxizH3uKZPbIH/MQuaLGTW2KBYNrcxkAHrYSVlKaS6Ly7FepXk
wgv/DUbchJvdiNS9rn96XTvhjGDSok1xXXs6C7mZW+SYtOFeM8GvpiWNgC5g
8gTfmRiLi3EWyM/zO9IdPUD1uFWMDgJpXG8MYEVcjdTsiCqHdsv78nBUdeZ6
qv57Ypi+CLkgQ+dmBbaqMckhvJ1DJKEKcZ8V1u0FhFjQLeEo0BrHmhULkePN
QQjz1D9r9YKlFC4QtQWpqaao2kBCXBxJC4giMdvWx4hqag7zp4QUgU1G3OBv
vTkkoNZ2+iUvmxAz/UN6KIM3hUuIU/BbbRUs1iJgZMaQdBTDqXrVOjxZXqyt
t1cAqVkNYzHsOq/mjpsiuUJ7fk6lCFiGbiE5joBRhj2qXX+cu6Lmdew1TaDN
erWfruVhMPNTssO+ve3ThPefPoI22ecPVo+7LJfMcXl9i+lgm9BF4nfLJbrd
ogF+vAIc4E5rmDje6qX716w9Om3GTYztn9pNzVTzHtLmOURUJhj1EGR7E6u3
0QeWF8I4+BMaXcb/PmKDk8uyAgw18LQxIL7USOdZj8xCx9RbR677BvSI8jhQ
gUwDCE5rddyi+ZdCycG4wwsNYUykv8adDwZLOz1TSwYDk9pFE8JT6EtPug97
j/sr1b3HZ8sZmUimhQu62MPsaGc5dPreT3wR+KJee0AmJnDUAc1rwHrYju5C
ffF5OAGO/YU2a0EBsfzu9QXSAmlRD/oLC7JLeMVG2v+ZlKo7j6pA+4NG3/p2
bTOmODskNFIpEmbrqS9xjBYb2UIIe3ELONIF9CJThczZwjbSsjGiRlMUUsSh
MgYEbVsp8qsyL65dZtC3vGAlpFhRTPpf19QsT5f9kYdJKCSUTjRbpBEvnz+b
YMkS4gSC5Ry/ehVR2MBamX1hAxw94MfSYvuMddddu/wGBekw7e9nwD72Wpcx
dCFahthxhJOtraZTjRmkOXNPAhP/o6yMfGhLV0/aeBY3eeDzhUK2jjqaV0NX
Y4mjvJXDpWLAtnfp3+kmlfkYwvCHAPQ8LwCDu+4YYh8bKuX3KZbqReiwr+4h
2QLQf7HxSH9fHq5AkZsk8u+xw0Q5dPrKAD0xABa/xYdUzdJgJo4f97WXC4h/
wdk/mN655uSWa2cTFzdM43eB+dRI6REhlSpE1IfN1VgtQVf9lyjptvK5a5fl
V+eRSowb1O/pvSQKcHWZ6w+hKCLZQePOUHZ2Tl1RsKbGExIRqJ1w7/Nf1ohh
R1jiUmnt9L6DQ2iXgrHGmkn9bcTl9ZnlpPLOjhcNrsVsqiK2vISFn6K1eRTW
sSRFE5dLeuK+cuvvHQ5vscj66Jq4jp25ut+UKCNXetZaEBDhlnHG50FyKpqX
GLl2azntR2YWwxF3x9dy1kf6jpxU7ESocyB45zhGtZy5YpuULYYh8Cv/FZ1v
Bn/WunokCqypzqfjbRIyff77CDftBYxQIykGTWtorCkhgdZEoryD6BBJbcPs
sSZUDk8USKL6PEbKM4Vl8P9KEzMIUEsquxE/1142GK5xbsiw87eP/g+w7Del
wLAVmSu75xj4T7Vyd5ybPSUuIxuFJgz5UcSsgHm6H4bMawMvO5Qah8HQjx7y
Ey8VJ1mP6wGSUuibObubXZdQ9EkacLUVfiw02CcNeEdR+RguuPwfpCaYaSKC
MKr/npEy8Tzt8sd/JuiHivoZQ/ylN5VAzy0H1aftrFwBoYsah4UFEXdKJ0qH
FvMXfgrOc3tc02t6k0XJwF09uuSzBRxz41mg9BM6+FbsYbza4foqYLfX+MZA
bE/aQVq/p4bFaDRAxCGDzASj8+2ivdSQ8maIUg5uqN70EPyOYCYHOb3cnDCC
Ka1NBpwkvjedRB/+HYD6U6moLI0ZCfSzIhGn94qRYJVzw/NCnLUZUr41NFdB
QiHwRBY6fdfhNIIQEKZZd4HUqNwoJ0VHqWlUsR7I9ysOOOoz4fJPZLBI9K2g
jNuaBum7GbhxAN6eNNj7zA3oZx0Tzy0IaTcbJ+PzuGfkm6RL4w8q9O/Wv+FK
nuCGHTJTPO1YvMxu1SL3uGxYFs+xbWkit7cEShVL0DROrw+5b6IBF+8IiAPA
YikC8gFXXK7edjWIriE2tdKgpmsWGqr/j1msIvYoPoKEdNLubIdWjTL6tYUy
/IfCwGqVNkGviFWRxlaIdeGc2A05DH26AC0L0kvePTTxF9Gb95LBQ6F0am71
hyWH0WLeQwRJzblnfq6GFb7SHnsr9cZTmLWOwW5aIwcltJWqTOv2zvADfj+E
Y3jIZOtvBQhzQ5IYSFCVS3HRgTgUrCw2AX3fMCLH3yxzov6MsmnlAxuXHh3g
2vRqJZCpLai6yGOSQU+4Mu8xFvQJwB0C9zRIVeANTdcRYCNXgFym/j5OkRl5
d4/5PUY+XgmGgz2e1gPohSoZttn3g2y+8k7MbU7bh0w0rVNyNQKKSu0xeFRl
Put7Njk2qFnmmAgdlofDpI8V+2Z7R/A9Q7lIo0zRyiX7bk4k5IC8g1J9LyoI
ZbZHI2lzK0z39EQiaDQIri1ObVRJKsQL11dORezONJMyOhZ5utrMXxX6wgVD
RePMbU+M5SwC5wL2l6y+88zA4oFilW7LQoPOtsJMtbPmpBj6WKj1PrnFkkGL
1uDVJs45GQEiEpzM7/x+Bfd5vG1WrqMlz59x2x76xPjPOi0Bywp00z8TuLSL
/HcnOWJumwYy8fnfIrkodhLQSYoPTuwfY2SN8rFXbG2wTFPvTDOVxxMcUOHR
/g8o5wm+iJlIZafQNdF+NY8XY2B9Wu3tU+l/CG5TSkrw/1UMeu5yEtd22q9b
fmv3inxSkkWDhQWANVEJJYJPfhvJbcc+U9C6emB6wDp49BE0vcZrnu1CFpWK
dtdWm+mEWQgYmzkK11ZBRdBvzbo289TzMXx+9kTPM/IAr8RfZyGZLGsl5sSO
VRH8sCj6En9Qt6HBv1qIxEp+IQsjRTNdD2Rpf7cCOH9OASRBS+qwPyH/0jxU
BYmPJ306MDHxW1MdmoHL2GIysl0iv9CVdb1u1IRCL8HsUvYQNygmDqVvklkm
/Voh2KL9qCpfFtpLUAOSoHfLXwZhpIqD0FC2IScQ2jfLSEvsKDcmiKZuyBqe
z5ozHaVd2og35Za96/7KB4nkMXy4jJAfxMoWfPBcDQL70HXZwv5916upZ4NN
/MeIFvgwv78t5Kr9qqEIFMHkeZCo+Iujf5emQRKXjdfcaSVT5/k1K4KYcm+W
yNd8HjFA3c2OESF7VjSqo0Ge8sp4ivS94ysHv7Kcbbc0Ww14Ob+QDxwNUgl9
2B/ix3zp/Yy2MNvqD5vBx/QcQzDbm9kJrYreLVqY8xJRXDn+JNqXXrAbfagv
2qBDpT7ZDmPxnN7SCHzeG+j34+rCl+Y6aHMvHgbzuds3gQOzllzW1pUtxAml
+Vm9TLBx0v/hTK8Idzg2CUq25udXVSO4z8t87uTiQLymXOKgu/djLMMUfQ2H
7yRhh4Z0AzrV5xBkPn1w5K0VipPn6PTqEtn/mHkdaPiAfzyOGDnpx8UizpE+
sOpi50uHt48okXDIrI37PuhHP3SAlx7oJA73+azSannGRQI4X6QkBD9/vXfj
RHPWJlf9wtMn2ZWXW2MUbEuCta9ZKzFAZhAHT7Ap8jsJUNC1JNFbe/GLVT35
+uf5eAza4ODCx0QyGKJIlz4e1W9JnHQjMLArSjnWEo8E3pOEtppyuMKBRxIs
QLgEjfnd7WezoO6O0b7U06TAKlGvymaoEpV9F1kz1zB5woYVkJORbpk0fS7r
giglBOnJs2RAzO7IaN1Pg+B8IXfbli6vEAPSZ+k2THj9yqH0zpTZFqN1i5bX
dY6oqdavzMdwYiupFzTMnyde4uyd17xfdTpfVSgUOGldEQ3BeBvsnMyKZeJr
stlf+akhK8v5DJNJy3mLhM/SHrA4LoxV4LsjBaUnsh7GOMAKL+tz6VfnqIWh
G4Zxjr6haOC0lO0qMmlve0tze9I//FuGV5+OU6Hq9mizDeq/PZug1upGzDXX
tok+QYBDk6Q+iVe/VKaB/DGW5tSUqlQ76Kvo4+U67M6cwMqgVBhQ/GRRP+DI
ZpgvjDHgYOJzaFa4fubmcjVdAeg39ewDDXGsPDIegI3JwNG1kDdhtpnySOVC
meDjFUTdznZyB5/e9nuRhUsHSdxiMjyBVNp7gjj2mx7FGU6y2AuIjypCzVCo
hTNcuJkeu1yHmAc5nncaE9W4OBlmfpcASt+1Jq8I4WnVvTOlJEN7OLe/hikC
EKIoJPUb3PsmX7u7AEOTrikkC59FStShcXNtBU6RxtZCQV86v3Ywcl8DJvui
BtkDW1EitlWR+KIovlEXFI4Qkb1E6RlFvkQNVoBE+Dej8kKAB7MxbHyzMlnY
HpbFniMLBPL9uQRCwi7prtO+lgT+W3jHv1J70LttEdntGJbMWMqI55d/4VIw
Sb1Tzea99ifRWXizMKBJ5fdhZJxv2+5oqXp9MpHZDC3s7mkXI7irjyWr3ro8
QSJJ6Wi2sk2p6KX5ZhToAbentEdupJkOumKf6CbL80Fp8OVI7EZxqZS3imed
w4mWUVTCDW+mcFthedvKXa0E0Hq1LIg+ca7eMRhheg6MfMlZCuyHdkyjSBUl
uJjeOgOnA+woLkkyAzRnAxO7TyWaG3384Ju6uQaLm6zVBmuCzdwQCKjmKO3T
i3WBt0R7gRe2hNo8sQg8cVg4BXyjFZ71cFjsR0hsXtO+5SopsvYUCm2v5qQZ
Y6ybjPLp0ep+3y1g3vKW5r28R0EoHWha7LKPWraGpb2cLu+3ujZx0T7uWJ4i
LmbkC+cn2a+Gfhg2kWXf9PFiCUAGBoHwY2gA/Ty1S1cyN5oNfJ/YVSigmtLh
bBnqNjZ+N/ZgbCBxkxX0umfZjBeu9PCAJ4zu/rctIDZic+askUjH0iqIZ6GO
3WGGQDjw2MtWn0AbbdURZ/2Sf6CgdQ0barrGefdFzZcrzTSyV2zxUaq+7mXS
CFlIdgeQOega0rwTnAzczX/igRbmwCG2rF5AXAwVqJXtroeYvDbfkonrAjMg
Q9MY2Nnu0SXxDxbJvzarWw9gBkRIDAfK86Vyxb0tCQW9rQtzDzawyjRRDfNK
A7rUrrIMO28HLXS9jgzHAT/hIyU9yXeXAPlgDaahG0Tt2fKvsXdmwkXpmtGG
7r1gm1ZdyYpi7k4vLiGLJZw0R6NoLp5aI08UTbMuPk+z9x8m5ip7K0t1E74b
5+agK3kYY2uHtPuRcK7Hj9JIqWdIN/oA1JycIkaa5anW3wj81PvexGvnx773
4h/wDeUjd8O1s3/qb15lvXws5wNiszGKjAetUqmaeg9DZ+KAWNHcD08i4cX1
pNaswKDpXrEcNbwKgjdw1/YB9CtX1xdGowbAqtZ+UnvLIXrW/srZSHsoH+4B
LOYHycfPnIuIbcjjd5bDhTbqqYVu0gHoBZa2M9zGU7B2fdYIVjlDW9pBaZdI
G+WTgIiY/PcUnwxuG/jyjOYSe4gqFxqvMW06n1favDiYO/HRpks1oYAnPtN2
10MHjhmCcGkocdsYSXVnUwNB4tFU/w5FN1reE/s2dUS0PmH4WzJPSh4PLp7S
3Irtht/h08fgyr+WfgF8QCvLWVozlERAPh54qwEtLaAuHF0lToY8E92iNQuE
YLe74J9raSP0ZVikpRLrQ8+IGgKgxrNk9L5/yvQ2FUM3jAy3WTYE6EIvN2kS
U2bIalhRWLDDkm6jyI39UIw6qbh3WDYkxuDYz7lXHBWXaSed291brT3zmNzZ
ZmuJVjSbBrDN/eTu3af1Dek1F7d0DdfLbz5Jd0ETjNGbU5+X6O3O+LSBw0sM
lLsLdMaoT1FctVMjqD5k7oAdx9SsTEXfAfmnG3GCLyvccSqehnMgwgh8z4tA
zGqzY7m+TVvj8tonooIhs1f4sx4UbLiRSHNw1y7dYXl0Mw3PObTgo3as6eP7
xmdKdQ64BbBEenTOzYeLnCgOhkXRLLoB9ieQ2XIwD6V5zgpBdwTmDMhyPxS9
jBEG+KqlCJZzKMEWAyTsUFIgE7EeOcaIcD1EgBEQSBhUniefRr04qkcIQw2H
kaqVAy523vPCqJbgj199juxsfnfyU+p+uw0tMj7DmKJ5Bfm9o5dy7kVBD74m
KqkNI7xgN/DeQIylJsZx4OTCh1ZO0ojq/ZYNgomlEMEKTLrFAlaayxkVWDgO
Ob5/S2yBiRUlK/aPPDBV/5Z+ZoaJ2us9jDTiUyB/naD7RXof92Bn5ammAa9T
h2hWFQ6ZrB3lcvMRXXpUkkcRGWBoAII3/0yQJDU1JRWOP9ICgdn1d/rYWZ+K
z7J68DiQA+5gaX7JkKRL/yL7gRPM2DDO1ST7xqVRoJlln7S0rAUh0a806efK
iJtF/qySz/R8iNjmQq2+XI1sMcjtLnErJNSbJYLJ3/45ZaHr+AfdtPh67AXt
laJE74OUC2dRGtzViFkrPA1TmVk8i22diss8ZjnnTXRYE092dbX29fcBImAM
zW2LhcDlv1UkfW1Wn7IHTHgryuo/QwcuMu5T0O6fjYds5SFPEF2MLoypdUE4
baoWA4Ak9rW4vPU6dalcE1uhDSmwcLSXfJAalI5LpIKpfXh7Uq/sBkaODjmQ
puRcPE4T8W725vo935ZmG3dCqoXWf2xt9Hvisiu4LBZKOC/tEGf6gEaDdqD4
dsNfA1JfznAjdjWXxv3yeZ7iI93hKhftLDY2urLHnvabruW+8EgA2Yxz9StF
PE7J6eEPu0MuHGAFKswUl+3ylPvPnikj5K2ehnF27tD54s0xVnWiZfokC5IN
+rA0RasMsTHDm1nOoZCGftaPppYj+OS8+EAQYs/+2N7iuvKv7fOcicnZGdnr
QSjAS/4D/mDBs3EHDfoSAXjCJ1gfj6BlWR63mlySWBgsvvs16SQp8wE5uN4A
XmeJabN+hdDhZW0+iSPV9gWMk1g3lq9Y2t+UvaOondAsv+fwxoAfE854FD6f
nWoSn8RfZAbtX/m3eYAqvrzxOWAvf4dtwcLZp1YmoCuEC7Fll8NRX22JVaz5
I7ofGLVEL94wR8i92nqgRPGocTUXvfEpn09/NvQ18DDWMwRVz5r8ciu+U7pP
sxKh4etzgYSd+xXaSoSU4EPCl5LfEMBHl1109aW3lm4hPkiqGmKTvtxdyz7m
C8LFyKJWBO0RLatXf5y4IZrPYJYjzT6BcLLCfrHBnJHNfee/lqwoyvAYqDwT
Cvb92tUP1rNunHwYeBwdKkO/mQqtTwLW5yNUmoiEiSL4o/Hlj2oxt8AXk9Df
tBVqHQYAx82PmkFVS6GE9AZOX9vAXE2dlfXohK53u9AS+rxuCxV5Mr2NMWWM
STn0vtoxA53DFwItuSEL/jSfcgKJKH/HjAf/qUFQMyRVvOlwlYu7no/uP7Is
4/N9jRzW7e13AK0zfiNzssjktL4XMrcIRK6aNOo+usNh42mqP0sGqJURvSsu
nZ+VxeWZ2awyZr2qqIBnXQsSLPE2SyPxuyZWXtnIHkyr8DfhLGogMbrKSde4
njKyzJ/rS8Gh63cEeVTKfqbYgraTJCnssNOWDzUdtmYrqCbOCfpLuPWpL+H4
5us6idhuYieJ5i65nhltPX70cwFIRNEP2kYIrhAoBADptOW4j5q30spcn04w
pVXXyRJ7B/gnXTuUGLakTWIaOPl/nnFv/dMw1vB8gNxtF10f7h5K2Fp2cNzO
HKERWoPeQ9YO2vqfl56DRDSCVp8eUeyUiOiBjeykFIBZOkbdqbjb9R9jhxwZ
CLg/hAJAy5efCQCPbpFowzaGgiQNArEz3cahhULbyWbjxYJuAVoruTG+8zUT
sWpAMT8UMpZCCoGbGRfNItyjEwkT0HfwRtfiJMzlVbL0fkHtk3OY5xssInHj
UfGz/zO/2xAYMDoKSuvPfM03hB03ZtNeFon0aq9RbGLPIYE7EsX1gMK895D6
ilChha6uF993WjVu/tVjxB8JaqvC+YSoAYBZf9bR8zuKDTE/9FmU+lQIT2A3
Vredf7T1gJPz5K0O+/nI1MO2df7gfQ0cInlyZd1f0r+XO+DUO3yFWAlDKHBQ
kq2grAzUJWSCnoJPYf3w8NXJ4cy4+8PZC0alvCl+l0wp8VZt9Yqzdzy4nsCP
0v5bb514ITSpHlUAN/2vd/MJiD/Vx9PxGgklF8JNZuCJST8iW9CR0paTlfew
23rqqxCEW7uLdyJMxvVkyjOAoNGI/CFJzXiYpLm/GCmCKNK0RAlWLtAKFBkQ
PpDtpauVn4sHNAdiFwbl2AWwOhh61FCYSFpICmUgpE2Llx9HJSQcqxE9/uMV
GqKwfUqnJwC/uVYvVhWLF9pxWiEGSKfjZcVYzdINHV5ZicjEmKDMBKVv8L9R
nysDrtbNLG/w5Gla40XJOnXj8nku2dLT8eI2e9Sf0ZK3fB+IQwGQqxkgMPC3
s/tLmPAy2I522gArLxZo1idX9Au3Sy98nseIpYmpm0feFN9arZod++B4B0qm
DNQKI9a6SATLNsLJcHibmc0xq8CjAGQumwo5tQUBYSSW3f2peoJ28fhsuif3
maPxSctTlU6qpmDathPtIkBwnvg7gwx6CuNQgYvMhRZ2KJNra0P5PFuC1U+V
Fi+HxNqHz3+FiHwjvixplz8xN3uv0LF/mwmgUX8V2HKrcT+yTFBUgE6T4irj
RGYFMxyNrTU6E+kJL5j8Xmji/cfFjPx9LJJX0MWwvEwKOSjrwzJR0qTVqDOk
ASdhm0jdyk54/Zv09mJwG0UPq/0e617xlDt09nz/NppDrsf5DVravcrgw07a
Wk06GcFRpeotF3Wf+haZYPOFtxP2bAwLmJtmQE4LyH6Wd/H07DsIh4iYHQtY
7U1nd7FyiEkuKLzXKtd0Y11Tw5qmhXfHrMXzTyOh4jT4p/cQuAYtht9sotvd
n1iTc+1nW5K1wqZDYxDJQx18zXCNak986X0w6vjRIaIMcmZALTjnet3vc3vE
9c+OZ3t7SLKXCIaybHQztF6U62Rmh4EbwtonvCQE80iLB/sXPwGDjkIR68r1
NT5AOOz2pmOf6iVb8wFSeLHewPhOaWd1lUokKCYAXTRsYt4VoHUNmlp5Skng
mNsR3lcJcsnB5HRhE8CpH6E1MTg0GwKKTtppOdyoJ7CAmvH83CPZ2umgPc/o
IGJOdobhJVQQGb+yfsCLsc+t5xWtSr0G17nEMlrVXNnm88zrE29fyiRIwKHP
IA14wTkw59sFvy5NEBW+07lHs6l+xDm97lY+VA0dHvbN/WfPMtRvGMjz105B
/fb4OrKX4VzXbOnTK1qnxMidAh7ldaTAXz8uM1k2hyNrd8smK55e5DZu6Emd
s38eRhPEhe65GPgJgBjFckQ8PblRp6kzbsHcMdTKffx01Yv9gV324e0zAE8I
gMJT7dAPTB7+GzG1/+7UdWz5mCUoluKE3ZokqVdr+jgceyPTqYylMpQFECUz
DJw3SDguSyHlcpNK+Uf1VycJg7nZC/VQVAAfu9t2tfAhgQPRpdcXGHlzF7QP
K60zHlh7FF53AO2V6eEZ8vaYiT6q5RjLeSxXopvG9GseG1vNG0vTuJwCAtXk
M8jZKwapkjUoSiQgXLBnFQRJA6U9y8JtAdvcdJPGs0IjG9cPwyTzIbXkizJr
NZ7nINGLxNclPyyPxiQoi3lSxVMtBKXR3Q5aGVSS0Pydb4EEoEywhglDr9Zn
+4UhHCNwKi3roPeO+jqUIgrgyU97OnsDC4Wd+u/kfKgqPxLRklCbo0dqgL8G
M/v1qekNCimWL3VCcfqKW3ZwaiWfPQ6ETqiCULjFNeel7SAAUKuURzVlZclh
Qq5Dj8mV9esTVgCPj5OvyPzic8LcGQtliw5kQLyTMrzV61j42jVPkFqJzmPU
qLsU6gCCICkHtdCdGqYUT+vi8o+HClBpl7FvxZfKfLsxzP6HMaXTQb7xZKE+
MiaYDQAxiegKyoGzFqZXCmJN1XumJMpY3a8xD8Z71STnvRHta6ylFsp2NGhk
XgAuh5fIrIqMw3OmX4hFNoD0eDB6NIiwJx79DSdRAnzRmf5G+lj2cdSxT7Is
Vi1hGHgdG0HY77aHzqXqqCD6VS7PSpgx0grYxDiRTKj8SaXu59GbEaWAofnj
dTnpguyToVEqkk0FzHsfRRGWYNn81lbh52eyC/7ULbKqDjlL57YxfvEuuXZn
LxL3WYgeXbPxKre+AaEPZ9NEgGqF+qzqOkJ8Zw2ir0wKz8q0Nr1OTeIHEhKw
yT3Enai2Y98V2g3Va3VuwbZoWZl0/P1PD9mAXc5OhFKHj9uOFmarvvBRpnk5
RsnOdVa0YGConkgF97lY/twL8sepnWk7eKPlCmextU78HIw+Cb3dhGo+kDLG
wQ8Hdq/OuSXWTs8o9HAL5ouWT9/I+/6zX5Use0voSNz0ogkk85nQQjamxh0g
6UfTB6qc7sya0DawJpuFvxwYw1x79HngkiaUBeo1i38XZKWcOhGoB0irQGzF
BSrc4BajhItPHxFfEbA8A5Uc9RYXXIrPe5yskSEjguPAWdoQK1tc5z1x5uEs
hMKIubWLqX1tRROq61Irmn9VIEi3OC+7AOf4w5RMV33QrbbXKyItzBqudi+M
f32eesvOl9dq0NMBM47Wk26VUd/HRAlC1FC3h40UWQrZds9TNyxo68f7FF/l
SHLpycomThcwSisnyOg2FFdzmxqJG1wCqphj9YHPV8MsnkpRnIzPa8h+mAu0
lR0WgUfYeNqXDBXzfBlfNqGBqDroJLZkDemfVaJiLaEO063w9FhLDuVd82p9
e+yWrkNVUUzAUIqsslZSPS7kVARweegvVyKacWbsBauydHafm3hy3Rc2kjQC
BXzxYnD0bGJI1y3Q6PS1EHpEMQ/dV2Kd7Ne81Y7pV6Z7rukbGi3qBZp2w0xB
KSQ10hQP4/fHddnFUodNj0mv7tyRElybXem0LIi5a5paZ3bWzNh4L+JRyWyY
KOtwEJ2ojSnG32JNKR2yrAuoZ6w2GG5fCEzvVkITEbmYszM5NP++nF3IFnu9
umeYvqIJeGVvCHZbyA0fPZ+MMIHoygAhdCPShQ4aj4oej2UYY+0GClhJuDJa
QS3lq2bMp4O94WOUOraP3TtUMw9gllHTMHT1dYSITEepD7hV3VC1YepnxryY
SuJPABn8dyac3aNByMmOpU500+zJzzAxoUsCpCX+JIK/eL8fsDwhTzGWKSQg
LwSQ5x+NsQ41Rw7ln1gdbE/i3hVeEgty3WPUXie/ey1wkmhEPCqMuEtTkJ3s
hNUFNKQ7uY1hIjkEzgwZCaTudOw9XW7MvrejRSlI1mivUh4JTBThF2qgqIEG
G4fnZee/fyatneX413ROzsIaKwf+NtAS2/msgKdH7YAUtVqUsULECBpmmauv
xP8lJRTqvZoB0LWC7+JxAK7rZ/7PLbOE9ru5UoGpl7ZS7RLC6lHLunwNBDyx
TVWkAn72dei91uHm2fdwln85GfoceTgwywbwwa/1UjSS9aMaK+zHqV38OCYZ
E0ZLmYd4S0Yl3j0JowvTcyM0ksHNtxMbMfmkuQgQQ96ucTwYvI7PFMZsB6TF
8UgA5xKB8PkxlaOgUyrD6drF5gXSsHJtTA1sZKuPB54PCL1gUIv5F/Feas0g
2Gd11UBGK2h2PJ+MQJ0RN2B5gMTYCePBiO+ihBwIr69tbtXIHXMR6EF9dNCv
Fvytar11UwzYoOHBXP8jo3rePkRaKqNhNypIsoa6yvX6HA+dW2b0LPuKUlmj
XPfAM+5/yCGwUjBMUrgHMwHqK633rqY3M01xSoXyduSAKMGCVh5OaNWBMEFX
Uu5tpWOw3J7ZT66Z+3qkbq06dPq7AI7difil8z0U45gRGckPQjUwRQidndhv
82VTZSC8BCrNU/kzrnhzMP0I0JRbj50jcgX47zgM/XLJP7L8trRAojyAji6L
cQadMyKgJqNiDQTuXv8yQ6OVsG1Cn+2xUFUDg42cIvL+eldK0vLiDJTERQew
ZBTzPe3AXqiqRqRw7d1w1awI8RPxJJuDeS3clJf5I3UEF2porx26j+y0un3c
OQqB0kpxa0aGSWo6FQE1Me3L1ulkjViyYFvM5hnUlkU3c+AlvPyRe3vB2NGg
EOP46Xf2TM9NcIFO56IrOq/mRu7fLh2tBfLnDJ6tDNCmCGhNml0xWuT8IZKs
OnCxwwsIR5l9rPBecBMkLWMffOQbBCaN4dllAj43j7JjfjNtAu0uibuok/LH
D51xEZJmlzQ8H5NJwRNOXaNyc4G/Kb+s6AeQJKegkXNB/lG3hCit6r8i9SUf
VKfV1fDhRv4sQsCQPumDodcuFcuOBCwc7Wl3lNSp2I+0gm0zvPgH/f42prWb
Ut8s/qiaao5asSJYRliSTIsM9ZWDTMYcLEAOKJfQR1cBp/9zfdKI4KfiVnMh
aZeDz6q7NEhGXWv6IjFfGKEgybBY//BqS6AUiE5ndxY9ScLJ9wH5lngVfHtk
szf1ImT8D+ySixnB9z6Q6/zEA956/CS9MKUGu/hrKNAMW7c3wD9yM5m66yjl
bPXKPgh/+gEl9ozRFC/KDkpx3MyIVksQ0K/InTiukv4s4l9P3mC016Lyq+m5
2kfTBNtj3S8PaeFRaxj8NOICNIpyUxlrmDle5CfDFH1Qv9x5nULOnJQSFTHH
1q1fzJQYb/8KmFmhatd7vV5vsp5FeCCusJ0JIgQTieIQ2Z18tqMekCA4/8yM
WBdgi9gd1P+SeKd26eIODXlG8h+Nm6da9N0+Dagp/cJAq8IdNAVnZu31UGZu
6ZYAb6nU4zhjbC7cmAniQzgdOsLO6Lgi0A72HNsfEBHxmTGUr0r5sYjJjIQ8
voRDaF6OUJLJ90G1RmrTf04ZnOiu2tuF7yU6g6/eboYiSnZVkk2iK4GSGVDP
zggd6Oext9b4nvpAo31zE8lIdC6N330MuU8hjoX5QMc1+T9h7SYuWJJn6anJ
Oe8dew+SN+AZn1rdjSj58H2RG8SqY73qTDS5vdClK4Z635fEcyrH99WNxaqD
x8tg3DzB7S6j4ykwmNZqJhRA3tyQgcfqWfqVI/8ey3NTIo0OlDSNa3x0E5uq
XBX+4bf/HUPaTnlMvD9JYJsjZmRSbwcIwj0eS0W/CCEXgvKkXFyygVjgYhhZ
Vok24NVqrL6Ad0yqKqRiRbXilvDGjnHee0fo9/eO0C6HAxULtMDRRKqLewIr
4q826sc9Rp8mjB8Anr064uBeMX8A5n1vhe9JnaowyWOHCBwCKmQZo17a6YMY
yOw56Id5T0e1F4aaJ1uVxIRglJ9IiUmRrSZywNsfGQJrRJJOAghCuDaE9n8k
i9SESxEUhdz2pkbx8mCONbRpUbghC0SLUYfiJtFqmny0OmwQ0pgKznIbLwS6
D4sz9y4JJJsP/S2W8Jt9I7+35vVTZhYOd2sSnx9BaiD6ZKqaLmIKdbKmtJKr
qfDLg/cBXfgn5tPfc9NHPLNBxn0pXfNC04IG0fUvOCCP9708Y+z9JR8IZzym
VKOcc8AOj5ijFyBuhRutDQLqbz6+zzU54RhjW0cUl8HS7HhJcwRZFgcDMrOt
nPT/oq61Cbj80mwve7EFRp7oTGKXpRcr53MVpPCFgDsAEDkwZGDynUG+Jdik
pa4CjjMZkpb/S0Lim/97Rll5edPziaVIIewxwepMtTqzTNIgjk1aXKkSPmoX
ekpUCr7OlLGdaR5ys8JKdstQTjJOMsOggPBqLi7gQ5BNL/XbkyGnaSikt1ty
t6CXb4sHdk6SPtz1Rlh7qH7tl9kH730bBqAL+VNVaMUzzu2I7RRBkGCSgI9H
rhHFyEzPLux1mPO7ChxA2mQli/M4r77yyne6Tvc7T3F1v2sWKvfss6u1sCu1
geg9apOWl3RhgQ8TdNqrvhgjZAx8WjAggl6bJr77I+9rIdNYr5T8zLYXME9n
L49Ian4Xr9IDojyOfPhuP507OxK8akOJl1cjSHzLhfIE102LG51x2tKFq/U/
bzyZABHC77LZhtDC7rOpGLIEMVtlmkZ+Y2ff8+Eb65PPBNCIvromefOiKSKo
72+m22qZoJfKu8zrE10p9ObRU8qZT4m+WtJ/72gPam+CEP56apfeU2velzmE
V5A/qYd1pPeeuKXmGZV/LE3mIGOyBbtzO7/btcHC4dYBnu3zBkKCmq4C7v6f
nWiavqhFPIxqgk1+pC066WjfSthVL29TRXXvsX7EYK3++pQ34Tg2Jm8o3XON
EcTHkKcyeKGmIofO16lczC+zxaEZp0/vg65XFL6YeWQVGw860wpinbEufadu
IGEYWmchp8HsjlvDLpyjARs15f9MEh1tFP8DEvlEgiDMZRZ4qwYyHV05+w+I
B/jM6sZXGuq+AqveX7yHZ8s76R5hP1LrpXIVEAGswMyUMzeXwlJmUWZf4x1c
mn+pycX/eeqDLNE00PiloXt2wx7lG4ERSKBtOXJlMscJT51AdCqGqJGMYDCg
kaDC99Es+60izJo1lU5mg317c0nmUnqNkmiH1ZgxdRbW3c6oor8L/ofvWYX1
Vw85VNTmKTLithxEwXgk06c2VznY3xfxIcCM2OZp1mR466uMv6RvCVbq2cXm
qmmkHyhLtKAQWYk3o/IY72Y+08sZ/n/xbKK8Einzk59v/mR2xuBtPVWYn5iN
UX8ruZCE2H7A9rbmLgUxIV5OIBIvUoj9DzB0poh1xjkoO/X+W3BiHS/nlrf7
7PXMs5dwSJ4x5NoeK3lMxgVRWvOeq1Er/k7ccTHWenu1bjShhrz3/c0fiOFW
zOjOLFIS0Uz9BI2WiW8rgraVzbbz+W12uNWR7io2BYj1IxuJ+l3QmhnQzmTN
NXAaBXPzdhjHu6H/Gszmr+/25PkEA0JBNdzPXOEdlX6g1gW2TBt4RTuHREjz
I19LQ9KCJhvOORuXYD8jBtkdqpqji2U0ZYF6nb1EckwADD5evUFh8+yLHKmC
aXaQjpqDU5RogzKI+op1wdABXDouc1OeIZbYAm+cSQPdbYlgwUfhDJzUZc9J
Xvl014BOwMczFLHu3wkQprdyFdGbg5nU9XapOHfCoeN4+gFDgBjIUEF3ZIkf
Q37d4DxQjhT0P04BFMzNqp7Pb+1UTcByqG4f1aTC7irQPbWspsAxrzoY3gXR
gerROQCizOaSx7QKYsMCsyFYeJgGZ0BGKuFcrEGBNdY8V0hL5a2R5KRA66Qp
mnrL3Onv9iiXJuimJ4Yc/q4xcDUrmiWMorVWf8i3LnBqAZhuuUYTtU6U2GKm
8U8RlrIbPgz5BVoC/JGeYcsSToqgdFj8DSHwks2RvkaMff8tC9G74zy/bsyp
gA46Fk9qOMkgoSoLtvH2vPsFQoTJjCSLnHf35C2DdiTMWHo1wqRlVp2/1bq4
f6+JToCNY+72pS7/EWPi7rhkJ4i6faPTY5Xfc7nQ20em3WIPsALiIN6enm0v
xvxdvegK/rjPkx4aD6Tw5ksE2H049Mm9dJrBLvrrlShJfiI8XcKhs0BeiaIz
1bWS9dzhA2GZ8KUKpeK98BGTEWw4UrXeReuC/CnL/nLNCLG1HpKn173DvCux
sfuBJGnktp91h7T0igDYhIsx4BcMnAwuNd5dz91ocj3V+JyEPZauNeR8I0K5
+q68AZABBDeQqmRA6YdgxjlsCXZ84giXMo6NwSfRRwOur6V/O1TXXv8yxHDZ
UDgzuYjZLeur4HWuznszOTltE1Jy8UTLcV3abrz6LHgR5ibKFDhV0SQOFFTf
OUHdpsmod3nwZiMWkcI5rJKwCEB1CByIrWLIqztLqGbtac/17/ovuKW/Qm4s
1550ewoYhSGFocRK5hMYjDzd6HQAnsU/T8f5VGOv+lW7KQRm/R7KbU0Fq/pA
9AkgF+fcyX3K6IC0IdnE9B46H/JahnXHbsSBSX+0G+/OwpcE6ZUgCmEbIvWJ
huEueZaSegFiys00vqJ7edajmbVAaww2b9q0OhaYxzswsyc7Pk4N/RUaU+xv
mEniks+7geJTDuz5XNku7kyTWKYZ/zmGGHI55TC/2dOP+u54vgARH7dvO+wJ
69CbQW0nNjYO6OW9/qnuHP+I6G6hG1DQeT6SP1PNxwAKAEHlzRON8/B/K2Zq
r218JFQ6CuARvpZZqss9MzZtKCtJWrlXp7N2+gK34wG3+mrgD5GcewXpIElT
1aF56LAx4QR8iWXBhoKF/UVXTB0IOAtcJRosLOXv2PbhseQTDU6NuZ03nEIK
0FAN4Cc1jE2wpjsz4HCnAp6fdZK77RwMVsrKynWin+Sa1fUD5PZhii5vKph0
DazmsF3UubxICobIwVe/ImWbs9YBMk6tYM4fDAbl5fiMSSCJ2XXgAq8veMu5
loemrcaKlZDguuQvah66KYUUr+KeHQ14MK8nXK1gGfAMb3ng5LyLstFsORsY
WgWCaqZRDMYlqRoCdV0qKE69KR4ixOQj5wJNcStCQA84zVCigE0Klmu7YOi0
tDKEtSthrWqat46UuTHgI3vjDu2kmiPV6igDXMt4XYKRZWpMWBI5zMizLPUf
WJnrzFCjcMw2GBuYj40Uqnef3/GDEyMbQAIvhwlI8niy2VV3UviFOROjVi0S
r8+sLHt8kxc2T3E2rVJ7PDBXAkNYrB3aVJ60Lq37uvfceL0VJd5EXVKmGtr8
/mlyt+YR6BsRAZkHHsBrsBON6xBdc3IkLPqZa0mUE8RpO0bDTTrIjKRMWN56
Y4JoPy45DbSRO9kHecEpvpV2bfa03ueli2ooJo6e8IL7GQIo+JrqWcUXawtq
6gQSwe64tFaS0ndr+4QYV00dolBZPo5w0LW7k96m9uzDACJaJZKnUp44JtiZ
KC5rivUcOdW3u9lByd+E973TPzxXiYFJqJZNC4iErWc1xjTL4AQd0FFDIRxv
EnZzhDAMZEFJ1imls8VXgsFci/SE0c32+QLVOYrUEVSRAFBpIZe1cJBx1VNw
lPNQJ3cE2bVbq6wXNn+vgU9M3NrldudzXuBUFeP7LKUE7jrtK0glEA/6QiPv
YpNdKtWanS64iA+2L2J5yTqepHExjEISZMQFfgW0lUXWLgGdl+oJBU1C5c6Q
M9zvtsV3vt7XhYtPjXm2uHTyUZ+YiaIVroeXChbot4an2u8WchzvzFpx7kXd
vE6spgazk3v8FwIuso5TySfbUmdP4TUk5Bz/yS9ylEjclB/WuOKHq9rY9hyZ
dbuGr9ZX+zzySP7WOUaN7S5GCCsrbtcwRERZK/+vDTWjmBjbKphRqy3hwlOB
U0pwknwp62USF5vdPW7nxY0H8VSffEQlQRrBy9Ssjq/4fSHA0UAca6d4ZXDF
uLiUgP/1ijfn1VI+0SY5MfKbbCfDQRCW9bir5007kaHNtiqRN1aa2Q65subs
ql1IxQS/6fupzNOXS+ixSmQDW1N7ty+a6t1aQAu0TqKd9L2EwG++aApXyRja
FmHfzITLdygq1MTXdVcs5zkXf4Ji3X2Rc1dAA2KcGTj583KbPXCaUlHIGYk0
EtslyLq/5bd9DzpNeP/ckn/30SFiAvjbI28DAJf9+IuzHtX685I8eYhxgk6G
A/zoVOIqOR40a5iVr+x+Vy7KsdRAnsapxWlDtgvR7hWhxF2ZJrFkqvhAzYhL
OCep74RTNHuxMBpQNZx8p42fM8R/e2uQm9b3sL/ToePdYJBhyZUgTW3ygX0w
avlnNWn+tyrMf5DThqW0mou0NgaQlCd3z2DeJWICoIZZWCYz+fMIZG8/cu16
wzJtbdtepHClF+XbzvgiBfHqBJPHbgSVwGjzY8ioPySxpSBgVx6As68ByTwS
HHKtGOOZuO3e5moWaEApuASfBokW+gJcEO/O5b5GseGElWr1GPnSmJ4KcVh+
/mH9SyFiGruBwMORPI1FPMesNs0MlsLdsSCdR7YUArMKrb+IzKd4coY9dsfK
r5BP4+CVZXopaPCz06QsZjsWBfYl7gQOJglFw5pSRwrQoZX0h8uk0wmv0iaS
tm1OONa9oEigHdTAVTbXlmCqX7pKJkk/taVZVghp31eBVgby6ZHgZW3pux8c
ruc2qNoCCRerx/N24TTHxxMEsPjhJTUnGntvCRtfnqvGw1mKnmUJmYvXIsRM
6fcMAvBe1R3ejaN2jw/iz2PV5nLb7B3aPDrYn0E5+8dkjqGFb80RJKjXwRJ9
1flfNZHI6TJ5zom914TTP5Pvc7pAoCF4oiSnrlvb+Jn5nCeVdIMDaHfnk+0V
zDgIyI4JoNEnYhvGo7ZLLLAAHIHaOqscZNMIf7tmjmx8Ly3Xcua5aWkRsJFw
EBYMPsrCQWM+fV/l/pADPy3lPj3Z0FAy0H2+2V8w75y64QlnJdoNvpHABzCU
kzZ+yFERQOJqZPcdpx4LoNDlA6sBFHeRY17v/Un0zIzRxIVzE5wf5bAkC7DT
Bo68x/XyPYjoxyHLejR+6bkhLMP1NJya7myoX4OqODpQJwf/dr8iO/jBBYye
ny78Oa4dhSGb2Ey1UrKHZ1B9gKtKwlgI9BXPLQtwLcCXapKmuwpglvQrbiy4
1ekwOE2/+4mTu7aWoWevQHTYmq+4C5zTcp2Z27Ykqt27pmf5QWbTeal1rsWB
VNRXLoPEO8mmoCXaJ1v1zHIAi73FjxieBy3Lf8SLYREa87BsFPzQmezS+/z7
rN90Z7BKjrYdZbJq1V1MXGUXqxNG42XGreLXXnT7ymFzTci9IUcBdq+uhxif
6a91PqwkPLThDUV37hDKMDIib375HzFbG2gBfxpeiZK5jBnPRsVkZ0Ubmrbz
ZSiNNQ9VfMPjqq89mUY4Dk2dqhU2x0Ua0x/d75D+19vpFlE6zJ4mBNiTuLlG
Sipz0eXnh2vs1V5i7Zg2vetnxrYDIDBjjxMdifZFs85T7dz/K4SFENnvHDp/
PAHKc268cp3ig/wMd/3JwIzylpLLievjCWe4kmK6kl1r/cQ8xDpci030mEAe
LlZp/coArKB+9aT8H1+8P2sxVKoGi5BAVfHls682HID1QhdDsdZowDb3yW9z
s3q7XFm1cxuDtqLPxJk+Xid+nYuLfuYrpBda1ttIFQvsf9Bl2Qbtq3hPFowG
IundZdX6z0QcMrsiBy73zByW/b8l+14sKouNumNANFQehRHB2+Tn6gfyrY9h
DUi4I/W67KO/FpR9mLh02mPRhGpwDby3uO2jrbg/9Q7z/IGujZRZNPccZyr9
4wv6MaF+7jC3VZWINgkMp5wpwpGyX1K2mD/Mv2keJ2CHneR+iPstqsdIrVLS
IXjDHX1rjbQ1YLSkTh56cYVcPVmHfO472v9Pil1yvwOv8jGXLHa5JIOZjyKO
gUWxhv784NjDf7z3+YH2yPIXfkE4vpufdlms8kQBH7zhLGYETguSXsAmtqI1
Jb/Jlb3fIz6korcVlHpaMipk8V1uBcRb0aKYsOu6JFJNRlEMiuMFcB0VwsZN
MWdvzPDXBK7zf8TxzqjDbUNd2Tu29CTJ1f7mpI8sCwb44KrHE3Oj8gcZsZX6
fFtIEEnWWrYmY8/Gn5DN3RSkwN6JcrYGsnPRYq5DAflWoqDrTYPuAkZwgfUD
8Anz6ZLSOYaNnUQck+h5uvF+n4l1KyIz502HwZMnS+cS9MDwbvqgXakYpjLp
gOJvh0z/8B50LJJkATqDm5AgslCbsZAGY75aVl/x1sldxRYVZI/6tjlJqVNc
N6HhVYyFrW7FrRO0YMdtGZJeySuS2YbLrzwowI5ylgtiFRTdENrMC0+Zllwo
Oh/ZqQ1tquVG4Fx05QdtbHLdfahiV5+gkJdhWwwm20BMm/nCUJvrplEiCAuN
kzsr+0A2z3Gq8LOH6Dt12gvJJCYlIEiYo6jmMMZ17IyLXkY32fXZftJxUVue
ol1QqjZQtrwBFz0TnzQ3ElT+TezWNx1Q+2vAhyz55GfVoG3NKXuCKsetWzjs
//xrH+wcHOfza+oclmQ/RDoYzyFJnve7/UtXLNqlPbgkCC1RXz9ZPdP08W1X
NvSN3EKIgNqcumEV/WQ3G+6oDHIz2bhf2laETTPT+iubY3q8gzzm8exy9u7H
2xRp3pApaXAYrINjOtNtL2P8P1Et0VJC7XBanLxTnSIb68B78zNQxtoEoHAK
qdosxt58WBVnpnAUJlBL2hKR+vDK7HJA6fUlTADSMunRcWv0cOQWyc3pK6uE
ONncLMcl5pVY3Y/K6i84tiP8H11yj1/UswTCI0BjfNScaxyhX/06wdToq5Ly
bdnS61Yq4kidi1Bzhefv+PoWC/7YN8EgJI5HbJ1w8/fHRISYaYlISE7D5A29
CnHMipvcW6tA14gssJWQYlsLETfT3cK24U6gWGf5KfDhEnRPb2NGoA9daALX
23LBiDGEi7uRoXOrzULriDP9zHWcqAJ1zMJ0F2FP4/3Ffu9GWzI/awFgxiyI
zc3iGhIXBElMef4LitPLVOx+2/PGaZFhzWOkcUfq0/ATReR1NXyM/VKph/Cz
146gArZDuSMPkcnXzrbTlTJXjWq17EBjm9n467Tv3RipdrN5GwumFDNIqH0L
ow4ulqpbpRTpzlVf2ANyC0jLelemfKaAqw2Wg+cPsQ1zUd8inRf2T3y7J/j1
TvOHTLAtUjYgAVbfXc5l8rln3HPfUiBGGdEMvlc+aLBp5CrL4Wz68CCP3Yvr
qnoWGCBYwuu3OasmFJDHjaEcHuhLElXculXBMcJZz2ukJE1uMt0RUNu6fX4/
b9NT6LuPVxR0lO3zIoLY+NmvsOpNlWQG/6CE0B/u+H4CDiSNRGVZeQyDTpl4
ircRc6hWecNSq67iYJz2U2rhr2zfR42kWODY6+FLkaxL1wipMj62y5BSyOSl
6LJJpA8DAZMYhAOId86fmxAG8vWyMUNXL12zwtIyAQu64W6Nq3Xki0y/VogD
nXiACRlwhFyd3L3WV3RRQtHcC9inyPMFgB8pZBzN40EfOIVJK+LjxIwuPG6N
zrgKf9eY4/ahSlRDx2Szm32Roa4bAbMrFtPRlIeDq/FdZ8fn0Xu/SUUoTZkH
kqUY3IOwSJ2y9Gw/BkpN4ql+Cbyl1fY16fPYhJgCrPy1gtTI3mGjgWSUONsE
68HT9tNtaLM00S+p2ZJDTZh/LSrD2S3f1iWQ335nljV9YKClAZviVK6I/t5p
A8Rr234U6kk1qz7HABTvbMtFVfCKwEOOCctodjp4zG/pHCkWIp4MQ8DprzzV
1rwXno7KKFanGLC9nQA1/v6xYxesXyDr2o4dloDQzv41HW9ITCn9olYgEphb
S+Ro+7X3CgeOQ6XFfMqGJc9lbJCD8wSUly63GRizgYSXIu7YGhN3eoETreXa
xAQ0KMfky41DTBxRAwVl/tn/mIUJNK9083Xft8zCpWt9tSjo0zPGxKqLxtlm
YJCxotyRxe5ls4pl5vHBN/ra0g+Z1FnmJB25rLfYYVDsLXO+MU8gf2GBlvH2
DGUGzAqsCoPmbRfR74WizP+DVinGMJMp9eT5cJr3HuDiV4X2ENLYROpUTbbo
CvLkunPS+I5vnUq/Tea4vLJZkvrSEF+Ct4QtYtEftC4D8QHx+yrftNmrBWxg
iJ7uDYXymLDjQKfYN7Axkjhu6smkhG8pfBMpGvfQhjRrjg0bbv5gfzAIvM8L
ZY85Sz1OZlfYX1jJ37YOOVbMnt9kgaxR5sPzymgYbzqYl//tRFw5cGlhajua
3XHuupIE51yGC8QA4ZdUnUBb27bZcXoBapR6HOavMuRb7X2AbwlNNPBiH+Uf
BO8wXBga27Ap1iJ/xsj7BKmpNZWT6PjWboErRlWlSN7gUBzTEC3lsWAsTpNX
w2JlMHcQzr+hVCKN4BNQscgE9dUj2I4QcbhDliWIjvCtLe0Z60kFuxckl8T2
nXkbEe4yBunOOx2ijibDBJG9KUYq3/09/Jxl/wr3LUhXqLVPTKzM74Qz19jB
SR1n9qnqB7IsTqsw3kRkJMAXenqukCCznmBw4zWNsjXB3ndw2aKBdGuTxK+z
XT7PgcEc43RrWduqGJuPba3geuopCyPYdVXeDMXpF2PJJVaspxsTzzLL+ANF
fa2IuNnDhH+nhLzGLB62cYj9foj3hMUTcNJSAHesuJw789sl4QiKxMu2dYYU
vSj4fL2CM8awVs2i3uHFPeDQOqqJ1Ef4u8SQeWBlWhYdqSW75c2RTN/VkGjE
68lc+J6ou/s0pseJcaEovZmlowPvT9WXv1E4PLQ9egEYaUO1qYdRR3O7FzvY
uZmpin/8W0pi6J6ahcxvB3Se7MoylWRT8/AmgMTJcypvj4UiYOQ8ITIP5wJw
i197Rmj2+ix1qz0cExcpu/7Y5TbzsP7dTDF8lMdtJj5LfZTvVOZh1WYUQkZ4
GA6MOS8D+qDP3EF4p7k1+RNuJU7tiiw/K0CDalcTlXtAX/T6PLup+f7wFUR6
s1bCWZ0pdOU860jYqx5uk0IoygSqdDAUsE6fLj1ov/xL3Nd6lk79v2KonsNR
cZmneijY04uxHb+4QkbMUQ7ch2+En8ToF1SA6efCbvBEv24uPCjJNQV4vLQD
urwSK/gIkpaG4EhHuFy0PI7BGgWoToI/J+Khp5DVfx/oc1PW3T8xdlghakW9
gJGq8Yp+Nzm8zYc54kNY6/RQTgqjQlB8u0zXZ9uXe62x5FoYOj5vqW+YVUuo
Keon4uPcsRkgfVlBYL8S0B4jO3lNpDXC5g81PEpBPRPcaNDvowCh56kstwUV
UyCEYrZ0QApNsPl1mCfJKJ48wivotwS0gvvH3RsniqYvTB6SbH026G9o6Oxa
DhJKC/UVk3ASL73DTFy9DRTqGnCvcIMpkeazFhhN2XktI+sxSnmuv4i8DQLC
AQYGbaqNMzHzJ2T/QgHXzEwSWmMkfF1ES8kFcGgR+5+Gz2LkXlIo+xJ+doDO
aGKhDsLF4Fv/bgImQOa2SuBvtxspb8PlgZO0qq+AxCq8U20mXQTQqkgk0aPS
Tempz1j9KAGoiDN6UiBfHTIeilEt57nbn8+g60eToDbTLxnC9uVx/Wq4J+7P
51pP350TdSUAbfbjy9jd8ney0/mspB4TzGTsIV5LHO9oHpXHA3QynfN8Dp/Z
hiFS+ePpjhFq6DrkGu8pARtgAEpi4pstM8Fi83NWUXa1FXC8eQPjw/p4lHlg
L6IZTkspD9UB6/qkVyRxqYzNm+Qjj+LfUzKzWcwQrM2FZmTSyHPSazwOkiSD
utu03YQw+6dW557BlKrjggE/JHt1uhEBuRiwTvab14mnA0VNAq/fCgsKYcvI
sRjeQeU7u195KJ3py4jfwqlZ3027SFzqOxPDeGwMsryz0lNSSqszepzxSonF
6tUhLukpqrpUIJQrdVfQaJKoy1ahFXzh6Anc8nASaXIY0FAngiKjtKIY053I
iN5Zz7w6lezWzNSw5rGwA7Hq9/fvrLwV/UlF+yMb9bvqv2DN/IgApmsDfEZy
hqLaPHfofmqK/tyLIEcJco9phLkMB9a3f2pQHKGWkaiAFSULIQLdnhkL57NH
5KBsmNxo65vsXQp5OnOsupmAZN/u1HFjFaoL2kEnj08RZLWxyksNqnRfTMWO
gJCZ6LaYgSzh4Yy3nTSp0xX42fI8AdRWpxpDe16cttDBQsVadfhqvLVLhlbQ
oMm4kJtPfQaI1Bejha7zUMa9Nj+dgykca2DDJFTSOVhzFyZCuOcJxLPKg7MA
PVrGg+nO1Eo0z+CaHxbND4mCqDlQ/PkumkNMWL3gOoyilnLbeZ9vTmcLI3Au
q5DUKICF75f0BHOBifybqrxVmfWYZP5oVpQqrDOz2ciwWpW1Ae+GHqfs9tUY
s60HyCl0vWkJXJWUxlMYH+GKZ23yKNpHDIHGu1h8P1vyNdTF6q7VkYqllGHM
ApkYXxUd0K0qkZIAT68/HkB0o2bMnbGbFj8e7MI0GxUgTmC/7b/s3ffJvf3G
nyRSGqTWlTs2CicToaq5SgsrzXCoGqo7cBBdRUFjrsC9xYdCts6U0mdxDh5p
V0eaNO+voVtP5fBeRZ8UJegEM9c2gOmEnhIpojf3rT/i2M5eq7JxJ1wIS8Fc
+36Q1Y0GrlQtho22t3FD+pe59QgXqkveM12fPTtjhj3xV+qEEHR587nIH/Dg
Pt6TGsrJPnQPnOHKL20hiAVPhNxNfz7HRCXQ/pVfhl0UM8nH6htv4sR3wRFx
aKKeRYBU/Ej69fBKi3O9hsJAWNhGst40gVspHiSAS0Qh4R6TwwyOtVbwYpMp
GnbIlnWtcel6dy6phJw48twjttPIe5eHZF2HVtbdtYIrrgQf0ILAoQ/xLZv5
UKzQaWkCg81pYF+37zpuH/Zz6uhOXIsCh0CAojAF5f9VOpY1CaKwYYXnx/UI
S8GXaJu+i6YVIzuCPL7Bi2k1ZyL50sWO5ks5ovZa7P/reDdYSMo3BmhJUQiW
o2Lodvp8yDWuDa/e/vY1RCZGfRBBf4Xue4PFzSP/OUBJMS7eBo03/L9L3wRq
Xq5wqPwBJyX1x66a8G2ESRXBkQ2XaA335EZCEzjy7ludtSZgAyIpv7qlA+BM
BSGxsMFalM7SXBhs8AAnpmA529ScdkjZXuDvSpBZzYiygQRBdcTDKjaVMzCF
xljWu90zvqirLhIEhNWGiGP9zJtGr9m9sk+FyEvKTLbatvbSps+ajIhlDqgN
CyHCRMV08I2wgf/ps/LY7upNpopBGVSPzyME0bCdUZW/M+tRauG55T+LPsxu
G0vJ6hRiXtu7+mh29hvVibhHa8ktW1Y4tyA2oZNlnjGjEEp3UvC1ZEr93dKv
QL11rsgYcPR0QmZ3axYFzzLCECU5KmmQr98cQU/HBenlE7eiuHshRHsZezZh
8AC3ebbeEstOJRbTYRc5VQ7rZe9qHpmgwESXHG/B+ntBHxl3pRZq36OK3Ow9
cIXF8V1wuQp5mTD9WDadgvW+zYuPE59uhLwpoLKZzHtt7CN/6OE71wj7M8fU
0X5PY3k+jlkjHAK29AvxnibUCbMNEEu1EhzrCiGUHngA27208tVIR5v62MWW
stNUwXxCloIeg3XTxQLeHyr+4JyADPBc1qFCZyOnXC1cqfphu+yYuJLtUj9z
efsyJ0pyTJ/PCBAVQbhQv5nFc9f8NgHjoa0R447Mtp/GLNWH6KfLaSEiWxrB
zZfzjR9qo/FFgXXN4t2D487LA4OhbaVGVQiDi3UVGa++gzFOad8nhSUGGEaL
V5kVK4GuoiqvDHGfrQv+pA/JJQyjruIfUAUmYz4mqkR6QJp7GeIEgWE9b0FA
3j0atAOex8qtm0o1yWuO0yFmu/G0r/AF+hnVQsjAHuqGwEWJcU5V+2o2X2Og
m6hfGDOWIwzq5bFkzlmcgraN8ZNaL6USLzrIrvEXWdURmqJDzBiAOcUnOvVf
uUqtE74OOZOr7ICqVI2lo43mVBcNKDgzyq/HQg/4mddqQFkK46Tm51XYNvjv
Ov7zspxFJ46TWpvt3+3Tee32/QrJKWB/zm4/H7V0DoVXS/B6zXmzck7+3K1m
LdJFCoZA8fjwhvHGbtjOvzu/1waqxtd0Ggo7LHfCNTM65tZJRCFNCCqFo6P6
khZ8eYbPkq05+0oGcqnzP5hUJEwC+bx1Ebr8kvLsio5CbNM6FT+DYUOow7pb
o90Bgi+ACWHXTNVLgYdOx8XtrQkNxomZxgt0bJ5Q5Inh69RHoWtyWOSlNGsY
YrzwPKMfDlGCAe4t1iubdFQ7sVr+V4SRpJvR0BNp09OGHBpjDGzpkFLH5teQ
boDJLTsqkR9rdmmnmoJ5K6N+qINrFDXt/KJejA43cy4j6h0OFnBwGGpp5e2U
h6wmQOvNLH53nJL56kUyf03te+7rQW1RRdTo3y438LtLzJxDTwI9FyZNGV62
2REpD9j6KuySwXuXpQVx2f0U04ts4DZz/c59VeqwESl47lCU8SkKmaq28uaL
G9+cFXfBCSh0OX9jqWS4JWo71azH+MxHFqcReJkqTxerGLho+NRGbqL/iny4
6tGvw1lGSyYgEhykHuPaaWggiUBQk8dF/0+miHbDm4Pek0y2m+gFVOiileli
XOWX7aA1xwo8jeiYttb2MS2OftY2BZEQ6eqNBJv97jGrDX/193sK5GC0BUKx
UYVecdu8x4eYVCyjuMAjTtvpWwSSczA+Vdxhl0YdnXjZYQo+aXNp6Ti2l1vs
PYGvvwMx+9/C7xthQOLYYHN+vqwnYScx8sqYJGcUuo2fjoY9W41Xd7eQ8L/Q
mVTqrf7pmbz7+SshP2uFHBxTMpMFR1Cx87PSteDg0L6pjlmohhEtrDWpvETN
oxnuKQQAPgSX6p3Z2YTik0HwgboLx+QhD/A1TauwW8IwEAR/7jJetCRxZ/VS
8DifVpiX5Uktn68HFhWNnuwbMEl1UWktrhFJHxkCYvB11Zh9uGwA4JrSRbQG
AISlHfhQQ4xe3XUxHcUPuKYbotPF17LwK7O2Bjm5hr0qLOXhqczIFAw3FxWG
sMxcXl+BtfH4orNUgfqqJ7r/Hc0cM9PElDBq8fhZ4ka8450RTWx+xOjEaFt6
ZhUXNIvK27qJNwHKQqMF+qAP0ZXKv14t34zwvt6TPBmoQrBzUL070vzLn5M9
TQfWennyF8xdGV+jdjShiPaxEvtq+/b+6erfVElv7tpPqF+LzCv/ulFdTkaL
A2C7fcPcKP28sV1NKwNIg5yTxE8PtSLw8Ueqip0A/p0B8b/QbdhGUP0zVAC9
MqBhgB9So1VDbd+567fS51CRxRUR2QSl67vP4lLP55UUQuAvAPf4OKmBm984
twrfl2TXqTzV3nrRUubCjj9b362EBkxa1misblKFg58W3UQ31+6lGdpOWFRg
QSCiwfrRnG7sAHktz+/sFr+QoJnPXlbNnPKs07OIUeHIJY+ST9opmcFBmcEg
zlobGaSXs47gs6EelqL/dxdYj7Qf0C3GBJlozcQ38ybHAVOoVdyHjx2TeJal
PRNSo/EBadV3rbzJpasS5iwL/KlNpgyZDqPSiocADV1YZ+UItFzJ7P3V6CBc
G6UPQoHT9aj5T7/sqFqS4nEKoWUiUK5HxbD4S9AyeWu2MScHlzXlQ+0FFmPj
3NnXRuKwT7g0jVshirwqpM1aQg5R0FHh7yteTPcgUma4DXSOGFNPyKkhvejh
hYfTADjijfHF3wSticn6SMLypQrYyDXVXOFZzHLw4Vny3JLLH83XCQ06L0yX
2N5ETERyLmrKPmQAgkQLfe9Q9FhKIjYtYYXpu1CUDfmQU98AvlC+TFlg4mbm
ulLS1OdeXPZHRsE61KMpQWQtkgbypdO+P2h+AwS6/dLSdHynjH3hJmn/jccq
T+P5+vtPM01biJlbCUYAr1ugJdQulvAIn6+TaVwPtCLzj/F6QOVSHhvXayfJ
75XNS9NRA20rw5sVhi2Hd8TnweAA4F1YD+/HhVm/bLiMCk4Wr7rsvd3Jhn7q
pGxk4FLjYjsZM7agmoMHYzf1tdfMrHvp3OpBvjd4s6GgJmUBHiX+msVHYAm9
CwZem/YbnXjr7Y37XrHVsBBNqvtLX9RxA4Dj63QbfXyehTr3Ry5Hf6+2/TCq
N1SJX00pfE5LnGNYJGGI7fJNXjlOCIYBBx2pYmgaqi6f3BIcTXdrQjJ4G+4f
GbhW7hTONWzCapSkSCOMfMPeORdBjh6ybQ6yQGN7kYiDS/4+NwZMxzgsp7BJ
3jHGrqAsROjxXYadnLxB+ScdYKPHAfiSTchK2fPzr5wuTvqjdyUQFzBN3wR0
HrN3Sz0aQdqj3ADXwMkDxSc2qIvaB+EaeIwl5a94DPI0tBQnAk+XUlCUuhBa
Bf0tokWfp9YjsBcgsCNnormJPm9Hu08yqipYc2wtfBEpxNXkDLbHbAQ9l3OQ
UhlZYnrr/3KsYBZNj+LQInn4Cne6GvC5n46vZ0ifWSuWi6VV6z7y3ECIupP5
w9HEMQqHuDXEYLZRlQ8g/AtOU+R3SRh0BDIDHWKYw4RLAMJ6oIY/Ie2BU8hI
Xd31lZip0BwwReGgHbkCpYi3PrOwLybdDM6+aRs/ZNjC/mQEqdeL1ILc4/oe
vubpSEZFbc91VQAH5OwtTeANxt5s267vmB0aPjs0jmdmsNDjjQQLlWJ0U9lw
22wtWp9V71pGuJf8PjuXC3lCNpuT83avXtR7AWMiOCjwFjruMPNerZ1Yo8F4
fqeFCQZSa2CygLFpRKdei0zLRrF6S4IK1tif9ONiM59hIUyhvParevGSOb18
LvAG3sR4bT8z0X/S9ynh3U9NPNf4ZzT7Y1WtefDWsFWDPswtK20pPaUaSZr2
LdUInhZVWs1B1RRGml8vp5UH02fKmBy9zpxmGvAOhqeWrnOB4FVDC8/TsnJq
4lQUmrczNqEOCBzKmC93Ae/nubjn36VUASRALTGjj0O+Y8YEeq3Vj72RJ4jQ
5DE8c+TqdkNVZsHjWQMaEUelt18qBtUZFghpXVCBh8Rr+hJjuy079tDMrpCr
s661NCRsFB9Q08WMftm5qb00r2UV3UJSKjv8FJGrCxQvTE95ZReVlJfyA0ME
vhqxyuVNB5RAkb34IaIAY3ri1sn2rJQvsV9xxziNztPRGALjVuUSMR+W75Ik
UZxDklYJyFJl+smWCe6RSfAt1SKHSwMXCOTlhXX37La+1yVQiMZT39sAUiiq
nbD32G5AJMJ1uqvOvZ4bcgrc/LePYj4MOxxekes0XCNBnwXpKOU+p20F00v4
5GL5NIlcossPxoXGDBmgNR1TXlSfhJVi6wiLvUxmU2Ikf4Pao24yryiFFN0j
D42+CIy1aNMqmBxsJZAip5IX4NgwYUccT9dSCCEAkr21/DHpef6WuqmZetbA
/uwIzfZKfsSeXfACkIOwl1cN3Xa01uii4V+pzG3UxINw7fb3WmV6lWpCirEp
3gA3Hyg/44bS6KKwnO5IUFBJyeKGResdHr9IeOZ74Uyp/qWoA7O/K0X6fvTz
hRDcfHUt671phmHJ9GeqMpTSEklA3WBkp62PIsf9OeghhMEIACUcw+QALWL4
0spT0I/CFJ3h/XVG7VKURpUoDBapPafYquRruqgejTsAaaftkLQQdXYfdyed
Nruw6dCZ/0TLX0WR5BBYu0mZR0wMAnBPnDuVmOXIc0VQT7zzpr49DqWgH+Ty
1gAYaKmL50VuJ6dkU57rWUxSm+10LwdoXJvNfsRV6ZpmKecnRgTjBxoiAGhC
41nO9HIKzJkHm/oEsBtTR186Qq7Z5YmxFYEVK4aOk4m/3Iww2CdsdPGw6cbm
V6Y0QDYucCzIufg3/5QkfvhP46hIeRZO0jC2F1p4if/zSABgR/wlQeCn3Zvx
MkY3Sj/4FVYB+yN5rneC5w3lE4DbQ8vc89l0H2m4l8iBEGy6W0ofCgN+L+o1
VJC1/1R6zII0YXXAlh8ifEP0lI/VNBfYMV5Wo5MLUB8bcFr7s8zyoOI4Cx1J
HuqEG12DNa3xGkWy2OzCo6Q9yvbh3g4HHGMnQFdPRH6fqVGVUf86Hm2euipv
A2Xy1rwXOLN6fFRUYYQlD9uCJcQ/LMVyKMRrhjb+93lpGg1GqF02hYyqWyEb
cKQHAd2Codj81/6oMVf1ylOCKr/m/Nl/e3TKR7v24UCDVW6M6x8ZNNjixkCo
Jq3TuHvtaFL+bZLAmsbpsflVy4pfLh38T0u3AAxFjjM5oHviSV57/IB2p2tn
1PxN17j3d2ZrCjHSfm/zqjlPM6Df8v9lFDkwRzxVldQM1w1xydRyX/5I9mqU
/UZowSXPhzc8e4AuD+rgy4AHryb1jxrzp4vmr6dJdgk7WVLZRvf2Dk8068PX
vClBbMVl80S4MI8Bczw77fvcBbDVrMAKN1XemU4wUrjejsdEHMDC7YnfCBAx
cLbpd4/yBID8GyDFVkDYkzh0awctGkkjs0wPC6u7Pm5qzsIGc2jUaKPsKQso
iTErZYYZ4/bCDu473AMWm5Sl6aNsA/Ab+fCouxuDZF4REzcqwtqzWxqKP2iI
NtSe1330JZFkioBF6JuP7h7MmlGI74+qTqTpPH6z5/cjuScrVpAi087A86Xc
oSCnzaTa879MSfGmy0h9vVtA4mVwy4KtbCyu/uGC3r6UYYc4aMamWKZfW2w4
1tjeJF23G5RqSbiBoBMxlYgyVMZqoiKILm13JMI+99ii8g5fGBacMeKFPr+o
6J0WrGULnklwNrkZANwkfhxGrVhzJkCrSCkw0yXb/c4IwpMd3RXO9aWhbd1p
1rksL3vKdmDW4PYGK18VSxk2nGZxkK/ddH20W1bEKDgoeMgp83iN0ZMrBawD
R2RXy0XCNnlt8lSPjM2DP6soYEBhNwwyl/0qIn9GYhPDfzNeCoy2ug2q35pZ
val6FJPTKyqhCd5uiTlR3AhcJZ8xjX1AKlwGBWpayExsPo8Y/7LB57aO1aTt
IIxcGrAi3YdTQNLxNEOhuBYRZRWs7JM088eeU8egVOEu9YaTx8hVjKgI3CP5
lF2KvK8ki5sbhScxigPtMVMdw8tZ5mjDZB8Gx5qMLDQGzgZPGU0gOZUfkn5m
akX2525VVJwfocEeh9vE/mytYNKmWvMwDzJD/o2LcKSFFdDwPYvXjSTHd8r0
7I4SmcBLLI//GIPrmOw8JE1+s3hp9rEycF7ef6V3Wg/7T2Usf3r0i23CgQug
q1PYEF4+QA6PR8ThI/PlWlW1AbuH4dQmoHV5laF7nw7kLwyMV/fU58Em6kf7
dD5vDODeiATGC+oorzjtLCf3L3KDoPdTj+sLpj6zFR3MOD0Pb99vGtIolNcy
Ul9gkAq77tOc2Gd+H8bCuLeFgAOffcU1+KyTQsDBQ9AXpbnN+vyAMWrxSEsG
+XskolYiWTB3zQjVbF35NUSls4r2ctD36rri5I6wPO+rPNy1QC2NQuRrTnIV
vxstOggTHiYrSSLuDWBQ7250icTQoVB4dTvlmk6fsiygTDX5dWqzEXSpvGPu
YvZNx9hzOGy0uBVYgo5njlcOus83MJkx22befjhpvoU2hOb4hrn0zdVX5htA
dEb/4nruQJDkNTsSKABmdKhoNY8afD7ON4djCeOYBrYVF6CLsbfN53Wuh6cO
0ila+o2g7aIed6GGTW0DwdDl7StTCkVU5rN6j9xJ4vtQ1zk7PsgUcTU4+5bA
hkLiIMm/bdb/2X7WargkgrNw+EaqpYLeVS+3f/C9i+coSFJb1HBFVZPLlKg4
kIFXscosLebFbEv55ImxO7aFRDmMyjXpWAQ6OdXlLeYDRtP1qniB3yPNDZSa
5r8WBA/oqbeqOLaH0tEeiBJbctNx9hi6Z8z5ahPP7QgotqpqmRHpQ2geKEgI
KeMv9iox44G1SLEYrt/FC8MJjDqeNOIinIIZJfnIyck5yQGw1bsVJW0I6jFU
a5qA3k0R0mTyjiPhQ8HIPOhT+ze01bYzJCTd/QSkhfM8TrEUBLBJKURuzis6
MOXs2G3QmZzlAHo76J9Yxq/9tRMDes0Ylr5zxXsgMxpvTos/ROclMKbMgFPe
zvkc0iaa4NNrSBuTfEt0L6Va5lMUuaCNAe2tqPzW4QSmzR0R27Q7B5qZ860x
FJJ3x2a3fn8LUQTSjks+sTBnrziCPIl75upAbkwPCDAhQvz+F+SY224Bkk4a
v6CoSJHtuznJTt8zkAY3ufN7jwDvtRsFn6UM39qs7XGszlps+Q6MxqXMVTLA
QRVUm5prdf91ViDo49Oi2SxywYJObsyyT8G6BLmn4M4apE/bbKUjmVI187vK
1YD+B47D/3ck+a6fV1WZvJFDNc9gqJM2HGB8/WfxrCJL5KvDBL8vfxLoCwwc
O2UzxWjUqcFtOlLvhjEtigReD89cGxERshdJ2RWPwI7adU9LcJOByfYabsgk
G9ZPvbJmEyZE0Spu2G3crN7DgxeyVA+5yAmn6v862Y0SNu8wLsjy+hwswNsI
z/76dhqvC4WmNHWcpyazxxRnOLAEzO1SCaF1Y+FzBbMWcPXmvmGKeQ4fMnqg
9CDlG+9+hx+++1AZ9hKu1ofIUSMulYzYYdYFukDIkeObCyQw+YZuY/RWb9Uu
Cbm+ZOjdIDP1yO2WI34HhWKdAk86ydbmVAI894saO60YRhEgNdMQlynreqSa
n7GvM6uNYw3d5lXNdZNS2hz0n7TnWrspJlgfQwd/OwWg0e/gs8aa2vWZGUtW
LuWsuO07bBZ5BB6WjZOtiVtZ2c0zI/ORF0ag2T8FsJBuTZSf0Dk+mnxKE+MY
d79SKrfrIc5OJ3O+pF75tC40031Geqgc3QyTBX3p5RWeU35Fvr0CV4kSgBHf
3xYEiFrBWVB2J7Ylbm16Xm65CEpbbdx7GAmBOsmXfgJs77vo8NHEbx59hG+B
f8+f7wmcjSrc182K53gJQ9Y68AzusvUmHR7ZMdnDytv8IVoVyHSMo/zy1gyY
2cKu2GOem/tKJl3Pp7VbQoDuDe4ZW8ioCLZTA2HXHIKsFYM0mETCBYlVb2nw
xz/llW+6VNjodKq68Sv3L2XvDVhGURWPfNDZzfCZ/6ZyWZ5f4mC4czu0dpeT
bNDDKKEEryIpvyXYBieQatH1rhy4hAEiaPMGW2YaT+o73mx3HqjIpiBZOkZE
dXb39F7GwbNKjIs/28QyhilJd/GDfHIx0/Ija8AwDRDSlZUHlXixwpRJIcJm
o8fXNcY7ugWbPM8VjqVdwmeKuH2kmEMReYLheS2xKU6JeaEp+Mymy9f8y9I3
FmVbTdTu+BqZ9fsi2dvDV/hcBbq4FbJZzUfoefF7Eq3W8RKOw2/9L8n8I8wt
gZq2d0Xi88e5Rv8AOIeLMpqYzE9YiHT+EbkqIyg3TihnMVEsn4J8YqOyZ4uA
iM0lT/g4waAEHzf6kaAFor7x0NEzMtxHAJUc4yIRNsykzCh9/kq+gq3Q8RJt
pfbJtf6WQ7mJ4rqRFLOl2CFD5Ty/QdrmUgyz088WeKTFMH0BGmOczJVbyWIM
NgB1khYnEmUetNPb7Fyi05d3IaKXxBPz7Af/3mG4JCqU8P23EewLeGQWlZR7
/eJTd5uZYtg2tvxoWuXCdPMoPZRuHcExvCURl+RWj4OtNYF7+F8erlpB/lXK
wvXSN6RH675ogDHgjtomVgMXMALbC3i62JtuTvjzEEi2reDPCk+X3gWjv590
O8M4tkJdp9anRVCKwqjo1fgyZs4PkErN/1WSNVtVFPcOgGhu1dwKIUegtq1K
9wa8fI9VjTP3dpewpaphXldSUrs7HFgpq7HpCBeosh+7AAep8b9W6bdB8OpD
4yfI8NBRGcSrFUdBt448s2FIDMNGMtedfBW2SPBHLycr0IuQMk4ci+K0FHzf
aWVw07qURFRJAXcQP3uocmMcyQ4OyLfdCDuEcrMqCWMt9Y3BmJIVQBaiYQYo
OhX+GVPf8k8sUiEsqqmqgB9HmqlV5bwN4UsO4oXfAnuvOS3W8n9YI09rKkS8
TIWpeWhuglaYAkAjnPXvUzBZTRYohRKUtAtlgQk82tLqQoapjdljgf5v7Ui7
hrz/DyJ/gCG6Zfw/HY2BQgIp7/3XsOhGbLcJ1a2a0dxg81ySf7NwjKZh5/Kb
6dRfINRDrHCvUJTacmhJym5evEr9DVQyQ4p9nbucD2juMnDkZNaRmkQ7750v
QcNW0NwLCEL2JoqJH5J1V5PnOdD0v/OfUkOIAu1bSmrbpOlaS88Ong2Xq74/
U8dmANHLc+3NqtFqHk+A/5smzOA6qCgFuMKqWXm2/h5vAnBGg8qX8Ex8MIKF
pEfV8osSZyv+14kJQoiWSVGjXHraggUvf6N4XjKF6ZRxFoFd43+6D9XYo54n
3JFgDgbxaHqiO4UURDUPx7nhPFFdt0gG0NsobdxpIHnIV064oyO6+ehHAez+
Ur5vpFjsc53xwlHOtm13lqLUU84uzFtF+2XlLACgx00ZeIuQNLZhliHVHa4H
V0BhL1Uqn7KFkYDS1EDpLIa17wE2Lurt0R53pVysXys5+UNSkT2hrdWPun9D
+Nny45SOU2kr4A8FBNZ9iJGwMbMzSWch0r5I79mrt7Ou3uyJIY0+RB0/hVSj
2TcKtWGB+QM4/tLBXufrNelhulLeFPDcfkqs7WqsXj6UcSvDDV3aYSpctT/G
el9NNW7OzbmLnsaO4h8PPyd35U0TS4Km0JF3ja8DOUnL9P1Q1+Vsp9TVEE6/
XMRay60AVhp5CNwrZ/r/xPCCMVdP85seTdf3m6TolyqS8LGmPs9I/1fc25y7
eYxgR03fpVSdiyL5ZY+Uha8XHwPX9Gg0uMlltsgD3trwVeVP+P4z1MoSsTUX
B/VZTDW221d9qg/uEP68STomU7HOaPDVpDWGsnqrqB/sVDwp7lveHmFAct0P
kxYiw+LmZgibX2aEnt8KwT2VL6I06pJAeDFN1blDUa3rj4Vtm7Y/ZYtC0mGr
qMA4Z9P/xgJYhITwqNWgPHjIq3lAewmWYqT4b7Ji+4tOmXykGnRNecfrQZn+
NBMyOQOsIiD/RmydS5RU0fYQIMrS5ZuWwnKXQ6JyU4yk8Xd76g/chi+IFlW1
fQJWJrQwjkhhzeHhgRppLtdVxS5Yjj9STx2UwXWNPKIzerhCNuKFSOfYVGrw
tiD+wfpxVfNLx7AY2Wj8hb9ZNBHe+Xctku7Y0ZOB/mBYfmgAHHVtawPVFD8a
Ia8HbeqPBuPt6z5Ulbz7eX82pwMxbXIOSQEPmwQtQgPNocEToCVEUgVqo6SL
rrPdxko8+NWQvvTYad1s896idYzyavSUcUZaO4jrnuJcQxPe+MhtMZvLP3pa
H7HdX5yYEDiYtQLq9HkqUtS6DDRf4YjG4WJ/M6DPhC1FLLwAcUbCD9/SC4HS
WF4bIGGZjDGtcbYi3xEPdcFLzaInFj0IRuAVre0rA2J2Zh92DGY5/mXWD78L
Ocsvv38RDolhAelH57gd1VYD8qu+qKYuO5+aDGZxGZQVKsz3va5cTyK/HZP4
dbLOddT7Kuj8yc4j4MF8rHgMUpIxU/Ts4qI4spSjtG1JEMQ1+qT0O7cxA9i3
hs824FYOtWRHpRlaUlJZngVh7XpMwASe5aZubYrHIh0qX0SAjCzFlufiNmO4
6bMuvFmEACfBK0TU7oWq+OBQXqQd0CUMijoyD7KbW+UL9s5rZe1ebZ/Ut2vC
+QTm4DYPUuhhfKfyiKjGkiYVrDvxQB1WCfQSXPxVkXqI+9QQqMvr6tXw6lwI
oiYdZFyGfjlC/RgSpUtbxl+SbNptzuUw3pP1FWXK5dRhA20oSVm3zjrn2xmR
hUpmU4OMLH9A883lHR6dYSA2G5fRZ0VGu/H+iT7MYCd7DQTGS1Z1vSObAOtn
D6/TVx4Q4oCAbDdL+AXqNzkaC4mXh295nLzvOo+FDCbd0GMEMWRfHmpNeU1I
PqGb6ZD9FxZnp1puj/eSUP0Lv5Xn6bYDoO2ORrPyoft3DU/bpf2LZEhsjCRY
b7u0N1EhrWQNTuQxpFohl+OQAkam424U2mN8bMi5WG3ZPOGAFnb5Za+EmM3Z
R7nSzOEoyXkgYkWpPk6jvlu163CHeQp8WXjzKh1/Wv6iL6bkyLaz+ATKsduf
A2L7xYjmDvYvFW2lWK+Yk4XAvgh/sgTS1AlRUJyDMdhCMNZ36r9oPweLB0WD
FVHkeklvWa251OKUdYPN1MyAPejbnpy+MBOBuGqbC5qcRnkX4LRMPo96W3AL
Ju/OrHZPendXXP+QrNi1Xc+qqg0mWZZQfmPJgI7bNN6CruU7OiCT3vuur/J9
RKMMwqRrLx691gvK9JIrISoWeEmnUBbOxestqAPRP6HLKfapgjZfSu4ehklD
uN2ONBPZnjRAnP+upn8RWHdCtBC/3Ai1HbeBkiz25dtsmmZQHDYJqorYr37z
4622aBzrEPi5efmpOrEY+rRhzzI2WejiJOSP6JbXmwlIpL9nVNxpObI3+X6k
2GKLU226PNwrXY80MwPvZLvLDY/p/suzFCB0Qb1g5ibyiFPDZV9Nvd4zvq/H
UwRq4R/MwbW980YDABl6UrEbK5vF9imFaOBcYzsCGDi+WeX/xhJu3uJGU5yt
m1bSPz/PMf6xfMtRLLsPRy84ls+dzaRqug1zVY9gaZBhQCNwvwxr6Tt9/cDS
lCCDNHSkW+PiqF1UV7QBROzQ0WXD89TeLFqraOnsHtolOswMNErSgZpiYMBx
3cclMORnYZndxqlQR3nRJ7fBtPbkxib7Rp5imEIKgYCCgwAJBywRHLwrigZ2
Q0+XoCOwSuOASo7/kzGipMhSjFZUkfH3LOzG3dWhUPJ4zuY2OXASH2ftsDjk
HJHSU5M5s3zfcukJw/gj2Bx4ST46oaUeIf4BjNhm0o9xsPOPITN6lNFUl0yX
2Zdm4E7zlQQpw9WWw8ezEnQictdzVnP96n6jB1AkOE+6bEhwBaoJz4vwGzaE
8nGztWsHN5ercC8PCr1EBuvcxFBFTjzabvDoTu5iW4X0QlYr6M5B+x11kfNS
1v/531LSllW2o3/TvSDdSd7+g1tUeeTHMp3vZxlzd5snryCvvUQUoRRDMjqF
LI7MQ9cF9Dn3qhh2HqhQxx85aLUifOk/IZsNd/+Afe0RH8QsXpaCAFfzJ01V
jYHDyqm+EshjHnvUT8+cJb4T5Mesw8Qcnw1ufBaFlPpp7xCV2u7O8eDxGk7v
ZyccnFlaCd03M8/wQ8FG7TzfGmsoWuQJMugjWQVH1/JBARTVosRuXgD9nzh1
Mvp35rpbZdsGXFbGPN2vKcuOGcuhYeGVF2pvJ7zgDN0Pv368AFultgS1q/Ml
tn1gQeOnl0PMPnW+sumpVnFrvENRy3FuoYqO/GIyC+M4pzxB+JLAskj/Fcw0
f7dV3KP4oh7BeyiaqFmT8Xe7kc8wPfdmiHySScm2ylmYY/0nZNCH5zmM1/We
5U2+zApndpmhckaMz1q7DPFlXojaTkcJOYfsEfnM7KcYudztaJu2QX2NZnhi
DHtXOrPEqyXqvBqp7IuCDugLnrZnWUSYhTsPzDR9tfadn5zfKtglvUdqWu5M
boOqSUHof5NGM1VthBtB6lwTIO1O7y8ZN85S+RJyi0YkdfCFD2fa/FFxYzCY
GTDln4GtnzAHfEw2Q00DHdFbAgtaDMMgYv9PhptYey4gpE+0g2NnhQ5IEZmE
CwJq0N+vEDiBd/9Vg/8BK/rhFqB+5iqDsc0G+Y/o5R5eJlKzMmwwIZp0DWke
XzEtvCv/uEF783zApZanvE5iM00uRJHmZMrSaV/kE7R3nHtP/JZO+OB0k9Xl
hx8GiGIczwkAcL5qiF4Cir2WqHXzKd1575a9PO02m7ONk1UO8FVComJA3xUU
xxRMwmppffowAV/JMSy96q0Gw8oAzy8i4mEx3S/dXLzGK1rKBdM1mcobxmz/
8VuqHGQl800y56bHlT5GcLsNZFP++Rtxpa10LJ6qJWxuamYmTH5XO5kHF4RU
48ixKWZbV9SoqwqZdj4C2YWWUC0Dfp/ZvJg7xuNiRsI3S84/9Mm5c/ZyTlxD
gDClDChD4zTND4Sk0xuisvDu5p3i9k6Kde1DSFirsAw3B3EG6EN79kYMT9fh
v5pv98tTDSgNqvBMsM7v1cnaWdAMJd1h9s9lw+VpliRZ40uE4uno1q2CbP8v
yh3xolYuyKR1rjHsdND189lJus4b9Dd+JP97zd6x93D5Mu31ChDAP+w6+tzy
Qkpe6L4BJ/WQgXr0rbnsfICjOE84WohaFA9JhYPOqbE78vzRqYDpMu0q/wYX
89DjTn/ijsFBIaMfM6nCMVohtJJB8CGPoIxDXQqt3FadmYZQa5AJJmAgJjBx
yvQVQZWKP6IY+gz/GLW2rdeoDIvSFMoIHGd2xhh6iX82dkNg0oVDmks0QDWR
yYSqG+ZWNiYVd7T80ljZbx5bXFGE4RcUQ8u9VXkk0AcDQ2Zm9eVo1G9XbGJr
+pHcBYAKgl41eLcfAtKRM6G6hZk0LDkIl3tQvGxyod81IpoPaeooymZdqPpI
tpBc9CdA5/sTssWU342JlvuOX6LTpcHM+EysqT0iSU8oD2BhAYsh9JOKz0wQ
4ZG2uEE2p1tzePLEMSyzxaeOG/7b6IJGiBcGgQxVCuVCpCe8v7yMOUUV5Dd7
jpeLq9sFau4josxRjNjyEQGccMh8YyBLH4PjgXIQXgHvBmkipLPSSPtibrML
hcuHP8uzhfPKtL3WQNhTNLNi+sy0wqqMOUBwu59b2ZArn3gafN8key4Tdto4
KrotMjnrLB4NlhPeaiNcBnR6AN0Uwo6wM1ZXjidEV+SAZomDcokYD76XpuvO
Z0goohlwk9jP2w1bI2YLEr85inQrdcBeTazjoNCaRJFcpxT1LZhFP29zcCMz
Guj+oOzqvb7iIW96wRsP4qIKLPkcHqlah2XkINrpPk0g9lQp1euSIgiTcA3M
A6LuakJMbj6A4XbL7VxvCOz/Exs4cmVyKystToJ1jOA8IpWrSlqAPUvEFgYD
Tr0P1erVvVOtjRzWTTDqu/6s8+F6hd29gySA7nh9vhGHyANuiN7G0QnDWBZ9
B0U28ttlFDkvuXlTK0EMUJxTOdL7iOapv8IbSjP7iS5DuzMD6jYFJ3umt+IX
uC4i7i9GMdfiGqwQQfBh7luLOFQLZi6TVI3QP0AVeOEUlABnHlpWxzw7q5GL
hpkQO61Ii9tMI2bOR6az42nAOaNKv8NJiQTfehYmx8ILs3pxhBKpVZ9+i5WA
cU0teHyydJ+m3enrlxvwfebjTEPCPJao+CRNIOTKXE6MPEj4ir9SMloLXpO7
dc+aVPEnE/I7ePUvk/UPrSCnAJpoGvrbQbOQE3lWwEIgsu/XyHN7t5zV0VZn
34DccJ54j5Jo8NKom4CROumyepIbErFWfx2i0VWGwMjG2tjh75dXWN2fhzmi
ShXqO6SMjrejKtwSg8sLwOtJZFXQzC25TN96SkkBvggOIIM2Qwoc9I797rM8
Ns0dkP8CIsMGCEUY7pMZdq6hIZc8ZUZIbmgbUH1iKBCUrmpT72KEtDzIIX+Z
BALJcjZw0PDbN8ky++SXp8yPKNNi27nXWBdKLMToi38zePz0BKaEFaf3iqjr
MdxhAqWx9br8Nmnpqy24xErHKxXAVXPtne9FRFB34vQTZxNCsHT6dK7QolCE
94nDBMtqcwEqTx29yUewkRndCuqAGZXc8eXHV7wsVAoVIqJoOSRzyK7tKbKE
bT25XeuuK0UB/geoONd/+NtVS5dLFS2cqsFcpzIPbKEe00DDF/gBSB6hDSNJ
T1sGlAwfVhtEbd3hK7juRc7YopeEtnG/CO37kzMi40rYf8VQ6xt7k2EcHmq4
GJSg5Fh/PU3DOctl0zeLi7vq0+tuUKs6ZaN40z6hmb5IlM1ayALolZn/ayE4
bDwf2kUZtKIYldgD2LpP6kZ4DHyFfVTh1XXEvkOs9RTX98uTk50+Ru0iRet2
dajmR5fC3VW4ARINeTfY010irXuH026u3N5RBYSC9rAvobHETlk4NxzQST59
snUy3y/ESP3f3PTMgI7JcoqTTchRS1EwGmf/lAr8+XGKc//uJS5B7HJn5Bjd
/HodQh6pzlAI2aoClMH4yVOP6mbLloaQqQ+5vtdJzQcLCUJAEOjx1AAUQM0R
fVM8pzXg/P6qEaC5hUnxVtgCwVq9fvPl9HaMK/pgfIlfjww1ixSScOcSo7XB
BPbMQ/oBhvG9iHVEaxjUHotC5PLqOs2k7iZj1ag1NbNcFkbZzuveZq+3Jggl
BYDqd16o3sE016dohl03rUBiA7mkYgJo2IoOryPHlxexDhxyiEgpO443yjoP
OQp3GSp2HGqiUN2ic4aNyCelpwsQRapVM30/ELIkdtzuAXhTsdmY2PR1JZlJ
TB3sOkBG+wnNAFPbIw1J+v+4jVq0vh/JUh0v9jVMudDVHgP/WwF8iwuXCLT8
KeBlKAq60hZDmCZyHL+qeyO7HVtOKaQLliI4+gW1d66Wp0Bk/aYLmxXDK32h
CYpJZLyxslMnQwTEhiGqJnU07bBksfV/PQN+S1iEWAQEbSmAuKeMihY7Zqh2
TCCELUqtieJNtk2buLUGMvpKmzOjTQ2omeUa7G3BU3onS/6wPHrRGvwPTvpp
gmMU0OJsD7OJGosJGq+bHXcwvE1vYc8f2fDIHFEO3Lt4iL6U4rQLvQqOw2Nb
YWmZJPnysA9INh7dtg8ysCByXAcZoOQOkYim9pku+m9jtbWCs2RNPwT88Lu4
MN6fBY4db0fJQdalIAFAtICbapQUYwWyxU9CHJAmywG8bEKDujSXFUtlJh/D
pt0AsH7mdj9V80sVOe6em2CBaxWfVJ4k10U/4xwMDCMIVYtqu40+tdbjSa0p
zno6UfRM4lK2nbUFd1WI0FEcaZCg2/mMlH00R0lkZH3nzKLarjj/e/zdXGoc
028XV25upMdy/KVj9xEPQlntCmuFIy6uGME5b73ygL4m1AY4NRp3vY4Gz6tC
wv83u46aNzoZcFHlZZ6KnL8hpOi13sJO9ZU6PsQbG8dN1g5qDR9Qh+wPM6lI
JjKT7MwPd2Z3mDRkpoPjl/Q63PfdJ++2xuEPlmcMMT6XZHZc4KX4gk4vP5dG
ryp7RguLVFtu119aSBUQzS99tIPIIG8FggfwhQLGMO6StXtUWzHwaRfkwAY4
DsqzFWNEFb05Qv3dk0mHtbsJVxVdg5VGzGcyIeDj5PLkY2M2XduOybD4a0sq
s42zOxwsFvoyg8nK1+RocuwPtfW/X55PmBMjxHLhJxyeXAe6RNaWSdTUXhLl
XD56cEf5l4QJd5GBItMo7boXUqrsWjf4W7i31wHu/rtnetcoAi4k3autGDtE
T1qUiGo/dH0Nk8RvXK7D3oFAmA2hp7qIhvhBDm2suAOmS/aC1gqDJV37miRi
SqEcIPxGWJRuHDgp+n9w/nFmFkXkh6+23Z9Mik0HsYjreAkVM/oetmbPE/Mo
v4jtR4CH8PsiVSB6swNj3cxH1KCH5uxOtM3lvtBKV1wZthXw9yaGKiv3TH43
L/angHTzvdtU/vGqq7YJbyGZWajx9G9AFY/7dAFqEgJSmNUAw9tOX6iI6RjE
AqgTWFSv4/ajyita1G2Wnu4+z6JwYJtT3KmoHUe1GZxNbkjCx1X33+zrNBn9
vIZ2GCiItqOUwXj+LE2ngVYw7kkxrvS7QgT/Wsmph1bSeAvjUJukENGXYLt0
PzyRETsFJcVZUhXwN2CZXkIqDcuvN0BGcAgxU8kyTmhxu2kt2a0x7QBVFqo3
uGaVIf0kD6EofTgHpIFvGnu+xxI0Ahg/30MIis/kbrjhBvt1ulEjslHIdPyV
9zCTfo13Xb8PqbNbBb4X19FFSoTEskcvMFQhe577X3SBLhyPLPDp24grkxYY
3KDzrfOgMxApEgPmjnY3Kvxn2G535ipbpTVVl2MLJvPkxFUrMXHiD+hFEasn
zIpNTDc+YAG74FDwNAQkCgxKr+grLCfe6JDBezM+0i9RNFaUx+FSu19WC4xL
BHFXbM6jRHbKRa4dC1xI6ZC31g8B7kIRn2BE7oHmW7Vz2o7+psijrVeYWCf9
guWD9SryBtEuWkcisGXYcXIKEjVrauwwL4+wQSkK5Vi8SVXqbeZEWilySqIF
HvK3TJ3LAfZdI4aUpx5nhIYnnWGT2D5WXcMhI6bPhf1ttv/FX8FYk0RD9BdJ
0bgY7wAbMLjxgPLH1RS2MwYfkEJLQr9eUyEDZBqXoG8jAvRiI/xKF4tFbpwl
NljIkw9zofxS+nDwh2uYgkdMwp42X/6WAU42pnv8ElUrd7N7blLxqiYx4Gil
VF14Pwmo+8D0ImKCtqTgG0/ESdguZzuTNn7NwO866iI14StAJ7FpSKPCx8Lb
txFyiCVoWfI0mI/5JECRaRR+g0UgnGYqfVVx7gL8dHtlTq+UCN3rf7ptAI/i
CBwGkT6Z7iPkkHg8g0W6lEaNyk7LYoqFNMz7A9AooenmXdhBeXepg/J4hafv
A90D4Tk+j88e+p/hGoKYrAA59xVbKRDKOCVGc6N+rM1iXmSuFRvR5qyiCPOf
22+ZgBlqzzMxTECsoyIplfY8vigVby/AQ4boC8v/H0h1+7ig0nAopnzPuptH
PqnEAfskbLNZrBCZyo43LXQDtmJU94P6QsyjXX8QPhUgDQtAaJSApvAUp3tx
wZNDbdRCSzusndyFk9XgZFRNYAhMnTJyv/hwCUZHlhUUIft6vbAnQrpmT6Xz
vR/4WtGE/I62EAknhnDRLstrr09rCO0nUSgiT8BS+CRiA8Pe5hZ7gijRyFC9
wG2phCq9/d7RrUU161fCM4ddXD5llGby/2bwb45ktm/7/z1MnA6tOXc6cmqN
DDktPjoAWn+4vm+Ocp0rTINYcOFvoY/WW/+FdqxKY4IkSvA+98kCdSebhJzj
EL1J32QUp1oU4aZSPR58qFkzWHeCCbRsvhXp61RzsjjiDxonromClqruoabk
bkyMQxnO4Il34gTjgKySkMzi+7/LMtXKtiQ+Lc5ZK9dL6untgXqZV7ITUP3G
X04EbkbcFEIwFmWP/f6EeTqyS6Ofin16lDieM8vW1wzlaPqyiiPHrKT3PbJo
bSPHV9v9ETb/4LfxU9fu0jAlE7r3rd0PmgxAZH9bzq0eMfnZPyHCQkx29I90
bXmDK2ylc4sr70fiohgPQ9yV4ZDfAWa8Q1UwNpDlI7S0jMSry0BshyUYUkKW
BihK/a9AjvEuASsq4XpPldnuqePDqok6XD7on7MuDDIeFR7IBvkYxxKh7ZwW
5zW0/L+5lQSDKsYYG6fEI2gnScZYivf4vC+tyaj8mFjwahs7+wo7UW6p/JKI
ALo0HOBV2TtbpFb7PSXe5Ktj1KquXKbFtxLN2ezH2k9xcGRtLT8yOiDO3ilm
mz57WySdLRPYi6ZWB761ZVKBqf1h8ALEpwx1GryVLXuvISbwvHab3w+0ERmO
u04f1+FR0QmW3n25DjdL73/P/4fGuwULEki5Ql0frXr1hzWgdErBn1ZI+SDO
+GN0WHEdO2j8P2PuDO27mr6C0MQXpZfc1fLBIFCgKCQMZ1sj0gRnMVEagp/t
UIAyoQrOWhlQjN9Zo8vkZc92xu34zOBwi6nhIlSnm1aj8aVLIyornVL6j/nw
HwUbpzPVLM0UJJzRFNP1ZCdqkJXdLEr+t2QniBxV+f99h45fnzEiryKP6Qqj
ivw30oGJinocO5cvyKEh6pvRiaty3dW9zLWuUfrmP/OGwd4yVRo3W9W2MfJO
P0kG0b7pLgF2fn9rym5gA7KL8smqnq085ypvXP6T5dzFHa+qQGMgm4g/SMLU
Odv0nM3Mwh5AhejT4SOeJ9/H8oVsRPejbcOp+IUKCCe/amG8Cii3jj4zTwKy
ZxbkrDiBLi6hPICP3Am1zx4LDSUGNSxUzE2/+7UBuQsbbp1cKkFlnNB2EMoL
bREejdLCeLkOmE92Xr8KhvU7EqCND0fn/5e8G/Tp4ZOxoBq6NxMv5NCZLoFM
MrJWlwtoDlowNj9hy38uxDwXCDBUtMlMX05myFSBrRm6H18AFWjI3OS5TXXD
KW6aMBABc58tzpg8zH3vQ+IZdxiS0Xwm/G6PxSSdvh6xJV/nDpnzNOUJIdod
VcwYqs4Rl8ePKO3riaLf7ixgsLxq5G9cW8HPzvN7MH9TgUxmX2jbsVM/K3Ue
VgqUBEPlp1Xshpcxe3hpqVo2TScn5JEiZenUKAV+cGtY/w9Toh488jKU/A+P
hHJhXBju2GTwxxbZP5pPIp9xc8TFT4fBMFiADhh87UnaAsDzt8n1XXYA1w0q
YKctHf+Dwz6gN5ADCYwB6yXUR7BJx1QLU1ac1Tk1gmIBKNj0sqBzA/sEiKlq
iR/KI+zktDFPUVy9Vb7NCMfyTl2B8MxYdFTmGE1+ikQfMsKo2Ce8zkuMLwSC
Nzz/EJ9DbXQ4gxYLL2CNDyRhZd0I/oBEjvewcwyCM0LPCb2wV4Pxz/zpU+9t
cNPevRSi6AaWfH75Lf4LMbXNI0Wrh46kPfsErRQontmk+Jz9BKCfW4xe5qu3
buyRckCTXHFNyqEqerUK5V3nntyonCTHPDyQVe0HJtcwzFXN3/KvStqFtD/4
wmdWUW7K7q/b03ffSjCzSC4pk5o29CYHxf3ufP7uoybPGeMForD8ow9oBWK4
8ZzyC0epHAlcau898kVwmkGB1uY5Xpt+7gIug4xgYdRjz+gSe8ku8KsBbnVk
Jw+MYIZ6jFhO91dqzxdObb9p5lgUInlF/Vh9Ay5JdNNjC1ysBGI+YCFoUL3E
1UvCkIdAyw7tGOUVZ1EKic9GK9CVSIJPGYXVV0HITmS98VY4fn1tk5Gd2VS2
VZ1qg1ymcMVCoK2ZvV0hRXhYlglLw/FT5vrwsOZg4RkHDrs+h0M06hz0WuGO
nnoeuv+bJpBLR2YQlekCkymynFnwWBqBMSZB6+uF82Du4NoMLtPi6gkkCiBv
+xvfSCKxRXQ/eSWrhGVXwFnC7N7xIzLrKMjc4kybdyNn+8fgY6p9EBQT/Fsd
4lXAT3zryy+h3Uyn7pbQOsiw7wSS+4G5kvb99UxMr+LCYYyjw/2UbDMFIfju
p2qgaCV1pOR+0nPjbWzNvWfkTLKvghap+Ier981gPw2smhUafaiw47Jj+fMI
FJeGd5ojV8lcALnibC7TFBHmugAYCICHNaFsd1U4J5hPDZ3x20Gy+vHWK407
zZlwl143e0VVKGjqgZKp5ZPvSkYZCAFkmT1+Wo9QwPwboBC8qKMGz554BsSc
sYewNqfI0C1ed/OL6uFyWQ59rppb0edwZP3FImkDwRceSq5AkVh33ssx1waf
n7L4yqYv4ZUFUTXvNMbNHIYPek5drKToAiDWzmcwaC4Fa2tux3nUfjDxmHys
9J5hOe3wgiUJmdq274306S5iNJbHcntR0F2iIPSDVLZf1rznw7o/KZHqft4w
Qz0xlz+Ohso/LhddKMflyS8kXRv82O1WzZnDyh3Z3EVcNP1hYLUQuKzsPsmt
PBr19Gdnh/S7LF4rrFBQy5mTHjw8tB81PTQSFOMQQFDq3L7eRRh8clRmkjN8
WOq7LxmTPeSgQXU75hnCOBjpv9uFmCbvY9TBnbU7TzFQ/iujpf8XhZ2DBzM0
YJtxmNDCQsUu609IJ3x9nQdE2x/V7AxeUGd0vTfB+5HRfljI8oZD6mxbbYS0
BcBa3j4elEq2/sA28w7pCOJtIbO43rZDsA5SOggPCDBn2xhu4IG4ZWhQNU2E
vz5zD3ND87/synfJLaslLxOgcVRTGyzUHY2u18ZyGYR3OSZKC1FUSl668Pur
LYd9XGooRlq+BJ31Lup5aVn6L0t3WLahlyQZiiSXCtjUn3yjyJaDIfcV45fW
tYN01wynNHhphug32AsCifuI36KP92TV/T0rBTf98R3VEhm5TRlrdgPktNIg
9KmVrREf3vYup5PuZ3pgivhjH1957tqcbfRE1/K9/HEpyS0J3sNDlfBg//OH
r8oJyPX9KkhgnGsa4/vbTJmQvOueXbKJjrRLFOrQVvqcFT7uab/8UZA5Y4pF
NwCWPFYkMQhUpWY7Xf6yFuyrXMreRmdzsFeAt+WiGIAxIOsCyAbBx6KiG5cK
7tmRUrerPC6gGfRb9ydYHIhXLjX27F1uZp5XzzaKY8fgdfN9xhJh2pXUHWnV
VLIBOe+/XONqkk32pPCa9YzyR6l8h7XdlGRbLFtdjGNKYEeNYFKLGXUDy4aD
sQxsEPozJgY1GWBeHKHWvsnkYvEHbgOS84izAOlQ05+MqvGEbWtT7LoVv9ia
djBkRDce9d16gmfSsbyusqcU3OvzvwSs01R07znnv1efrc04dd/j7XDE8US0
3ix+o/CrpML/0PE8UpfywOPqkkOCN/aLDwHzHC+C8VJl53sP4Z5/jiMSBRNE
tYd1n9T/86t36bM22hWeMFEsOi5rEAT+JS533cCfCp87PQiZl/VXgZXMNvFJ
axaHHq5pw4ObP9KcnMLHxLVsaD+KxAd/p/Jgf3N76HzMJnXuBakfrjPRR2Ds
5r6M8erzxkP3lwm6Ut3D4NGjxKrnQjYeFB9T6Q9TRpf5kS2bDMJPMDlFKG2s
hUazhtHsDhB4a6Gmdp3T27nFP8Tv2621ftrD+n8Ocj2LiFv2zySOvdPWVL5u
fy8viZPaMkikkcjwR1aEMSjGJG7gVfa9W84NGexpLvFVd6kxBqZqMg7TkGon
JG5Tgh+P0B6vAqWO+yId5OY4VEZ6uiOioLItcVy94U8Lj63Wb1er/9yWhVmJ
VFZjSLrINm5CA6EtYNKAjqLYOTJvuNwcCQeh3feEdX8P+4+PTgQ2FuzyFU3z
zrcwW6AohiFrcKPgqV56f9q1CQcDLBAMbNXB3wUlCKYop5WcTgEyw47CVq2B
QakUN2UUWYeVODGigDgoo9bAxaJ1pz93IRGiepA2lYObC1cRvDo5pA4Yffut
8KQ09MmPv+gjTLClWOa8Yv93DhTp+VtEXokPeUlQow3vyFPsXVT5g3Refs8s
5FqR9JCfCO6+WDlI2bJ81mV1X+CbrSq+qB7TJeFbBp8ETvGoP9l5ru9iryoY
CJ0CmDnlqOaSKDvR+G427HMZ0T2i2Wn0ZbztZpOKLRHkElcafg+z85AyIBZv
Sqc+K7wJZXP25zQsmF5jOyQk9Y6fJMHAnj0T+uYQ70qIlN6Y2ZeNWkDvnjMR
4dPdVNsvl6HY7Mj558oTK8gVCMpnwjL28hOBxvr5fIORJ4xMrnGnQtaflXf+
BfdGJMsYrG6XYJXGC8CgKMUt+1nV0OPbUhb7DbeljB1uTbXdkbaDE0oryTqM
73vZBWRTpjgMabHrUxHkHADHXXYyXLCyfylc2m8ZTig8pg6X1meu7j1Y9sv5
UaLDdxZOkQqjHiMyK5TbgNuQy8FLbDlNsMpdvRhhnLi1Sl4Jyrxu7YEkaPpZ
SjNhgHS/GbwmB1bTiEtI73DCTk0WnRyfs7AbmOiuJIqi7PCArzVSfgPpl1Rc
t7vpBzZ5MRcEP7cG3/ZLEqYe3no9nYsXjDoAdoXKtIMXcAVtLkeywm/wmpPG
vLjF8ccYFYn/PxhvGPbWxX20lVyonICxcb+BW1rgj/nhceHuAokDxMOfRZF3
jvdTlbzZnxDnGsuKSD4mIqog8tZ32yniTDOZAwwrsWDcj+oT+QFuCErSxkAI
ow+YteARV5OTlKpBQqEUlipRaMSkCeDv1XoX7xZcLE/FQAiDYOqdHZALlCae
9YnH3frPEn5ZUfhDYIugnrM00EAMg1LaE37w/pXAtHtElBDa/hSyzsPnwZHE
kI3MnAPI7mzrA9dBkHrb52T/3pWjuR+A7PWYymHZfpqkX5+TtsHTmxIxFYSy
XIdVk06r3cdTvFpzssNsjwH0qnIIOwtf/sLrADn25F9hgyuAe6DMumbacfv0
Fd61b//dVrD/xnNh1cZVFsvH7skZEQigkpAY26X/j+Y+8INLyQ56xhJyUMS5
MwhLbW2p+BGfpkuYvF2Tty44I9ojxBZhNxWuWwM60tmgfgK3CQvjVF56zok+
r5lZeXl3idi8egUF4LA6bMAH2PrldO0VjLfQo1VzkknCmq81zf7GtAopWT8I
xQ0O3MUpKveN8WpJm7sOqv6E0ewDUyhnqff3HdWq2PIWErfwjaRQZL/UnFUP
ZggTZiZcrCInCyrSiMPqEIJShlEI8gKhIbimLGy7Ixg7YStSBabD3mCjqkIr
hCx+gnAZ6yRn+/KNSHMQPbfn3nluHiCycICIyk8M/HWOgMqq+Ki5P6SpOUS+
d1Fwj2EnxVas35P4/IxiFHwCPOYaYVglQ+uctmohQ5Hq4F4UGPP9THedL4R8
z701KUDtA32pFhyHl6ETchNzi0MPbGQEDVf8Gx+bUpr9gDtah/zDrFELw0Wi
PzbIxSpuHYYA4gWxJKkUb6PSVzuzbjXeuL+zA53lNRv7RQrEWoNWuhoaTg5x
zP1zQ5hX7oiHMZdvUisActcWuArgoovHpZ/dOzk2ybs9A2+axYGklnh/oqTk
PmaS9TyTM46/H265CVFBb6hXC8qk+ijvtlRtxZn7pVgN2zS6vaSxTCyTIDYg
ZbesgQfieWLS12nSpb8yeg/cIRvQIUC2EpAdPOn08q2eGhPcDigS4nlkpU4P
c7n3AzV2Zv8J9iqAUSrX314Tgh7YVKbiplduYaDWNgs/Ft4s0BpjDuuK2O8s
ZtP8u3ktMwNgiZX78JxPEEER1jHMy6j2zDPZ8OTZ9lwDW9/cDNE0lSTTyLuJ
ONvKgj0LfNE5xjoZAILz2yrU140ZVvQzvTJxNdJYtf0SnROgRBsOay8qu/35
+P9jdq/GhdVjq6Q24cCgK8R/SUtXuKo2sEQD8J6XwxQ3yHpu6bBdliUqgdJ2
iL9qGKGZ7DPkeWe9hi83hilIQvg5rQTwl6qZOZ46BfW2/fAkO8sc4+s2mJB7
x1EJrtKbX57pNGRn6oYPl9vuPzRS8rEGNYKoNv8lU1w9eITBFeC0TT6OwXE2
jn8kG25OKJq9z2CKfd97QOaK0SatpFs//klupdN8SFP5/EMcADexjrDPVkXn
PllKMVxjaZ3DA6GGvnWFtmnE/HABnjiG9rxdc+OoguDQWKPABb/JDIHOFuoQ
DCSGNkJ2gPi5uYQUqiP2anTeX3zDo97DpwBN55cUggdA2hThUGQW7V9LhN3X
efqjvYlOISiLrfyg6sijsxQ2oxSDa6X6xqUlooFHz5AqiixL92mumgJoaIHu
t83lxWEGWcOpXkawtKOa0b7Zw0qwYVcHaYId0IlzgLDBYVxZCWC+9r9bRIRE
WIzYyeRECLXhCM+ve1i3hRZMOip6/AL6DFSdXwhgk23imSgnymQC3yqbYJzE
KwYjDuQbyj49rWw/1O6c6MTYryx6oUogKrYMTUaw4ZVYE0e8AhWllKW3y8y0
kohuSoZ5LAsd0T+rWJIlqkBbKOt6m5a22ZOdWkbYHiPHC+6OmELhtvsqfn0D
wv/jux98jOWE5MtfP66MvIV3EaZmHrKfJ3RBhx5ML9qGsSUuL9Rbk9q3A+jP
pZeXgsqR7hmMLCCXr+f7Y5SwgE04F1MYRtbU02HMRLeh5GUN0K7ZNZMfLPPr
pKPZ+pN4zRS9yj3BiBUFPzqn8aXqTSWF0czQp77GvJbytyHckmGaVY2Ze4ib
zv6C1XiPGWRMAcltoGx+di4u3Scv6foxns1JKfIqiGDp1zn5crshQYSDCtwc
n1BsXttUO7dX56lRkLHDtm6gFBHZbuSLYuWBGWBLa+gw0LLpmW5UarLmPPO4
LTsLym3W0dUEWfvVOVhBW+09KRBZz6DZdQL25q6sh5D9AdDROHtaHlgtF6Gg
8Me5h8COsNYa4WKus3odPwOk/17q6lKFTJ1XVwoPDxjb46ubanVXGFM5By2d
ILrvnGNyf1J3rkqNYVPzpO3Tp96DxL+Mk5Udrlb07Qyo1LR9/u3fVBiCL5M3
VxG3KAHdaEKQIFZoIp6GRxx0X0G6XX6b6QOMqmo9n137oaa5WaHomSW62rE1
6Y2Wt5AlVgySkDVr/eA0lUb4+sWsYZ924uXtX/T62hXgAYbY3HQstTiR3/cq
vIBxjFmgWgON1JZ/gHBn0H9P4Nfwrf23X+kJT0wuXhCFUWfyCoPeTN8Gi1dI
jH+oOJ+rS28wN81QsGDaOJTW0+HsqgPplvwty1etkOkc35tNVZISc/2t7kyk
mDadKEAnp8Fc7wqdRJ5wRuLcu2aQzZGi9DzQOr35rI5LUuE0osmGcdrAORSD
Wfabf72Hmuwm/4/EMGNn1AP0ObY3lX4bDj+1YT8UqvlL7JfOL4E84RJkieqq
ui5Hk7L/u9QhZDjT81yO8CrSQI12fmPEi1rqg753SbBBktnFG9zElst43MRm
aDBNoME+4Q0VF6yHrzqgjcT5Ivzfu/Paa4mtHwcKk7Bms6hi3kamZLB5vbUR
UkbeoyXK14SuMLAQrBJd+vN3P0ao+zAwggx361FjSWTqQlU58bzgC6nmL13v
p+VJWWvt+Xmq7nHNZz3CqxcrfTuQ4zwhxoJK2acLHS6k2k7zQfexv9LjX+GN
g1vyhsYUTUaA8ZOXkOIKJxVFCEh6HqmRa5HAa0LBmC+Cbdq9/M0XpvJ0o038
PUlP7ZDO13oYlnem7n/gof+zllNGQ7AcuhOiV93i1o4Zqpr40HFZH9878kzz
PpRZ8BWgVWJut9/Kn/qjXqvXmvnvn+/Fbzd7Vte5jhtm6h+AXVHCMsbON3HK
zua9hoWaQbb/6ojFsamOerrwjaGc7+OeEc6PWIwEke2to9UK6/8cu1+rH5Lw
qWs0kzrxH06BWMeG+uc1iKps0ngnJ/vw8EVgL2jTIoGbux7VkNx7EW0wbURr
GpGxtpbYSkBOBZjgAXWf2RwMAxhv2RjDNMOz1iMlbiOvGEjQosCuooS3VL+t
CFsN1aKPUFWqgCngCH8kNB3DnftTxskJL0r6MtmfJm71JJfBAPqA2o1uLFcy
eB1hmlTYRAFwtGHCCFM49jQpPBECB+qLR1GI/llzF/ExUl1nr4qUxKtRwVqu
ZmHtp71NtPlV9HcAzEEl15qK6ftwhs5mZQVwth4LcGguwDFHdyjFlVeDUT/H
tPfXpLzK1I6bQ7XMbmvl5ata99TmtXqLTrHAmaZDGqxpE2KRRxjWY/MCnoky
vNIT7IG5s5CJuzUjLWXJqFXANBXA26KIlsODTB+/2XEdtGQ5ICRvanNflXwi
Iqp/uEe9tVqFnYmWXmWvh68zn71qJaFqy3in9X0q26O9KaiDLHnDK+xlocqF
Y3r+FnYc6dGNRPXg9HRLahvAZV6+H9+QdbAXdVedXKk/Y5MyI71wLT3XuBJD
BdVZIVLGFbndOvcjDCO8anEzgy9ueGQ4cHTJL+Ub7Lo42tsrKSAbsNIEwzTx
aEIvnEnNyC7BLl77Q6exGpon4ORJWB6Xoi2WDB1oaL6JJp96xGCXM82WQEU6
RSnK6nmlYQfQ0TriymK0m+ezsFcHaTebTzZsmJIsminZcFkFqZM6OdeJJbHa
HbvXTcTmMNOXDWdAeWBRnQKCPYjAzTBmP0xxN+tilb4SWbQ1SL53CiG4yQ/K
ubkTHjiTVytk6UP4Z6o5CJyay1QDqNOoFk8jyzIWhbAN4J36eGxfWmQLlIcd
gwZpbb7bDuaJoGGrJNGVXCh4yUL5YeFWlmycB9l+fhI/l8wrV0UPV/LQkBFa
bK0y8ZwFXfdGg/tiHnkR8NJMwHBiAUxfCeT0XIBiVoZPOLBH0miXkVoBglQM
Iz1F/XXdBieOHaOQJwnu4rRdibutynDJvcGNCj+HdqNOKyoG6HAVxQ2f/Igv
99Ohwxq3BLGoR4cO2WGhNJ/4l4BtlItXIE9JRwODMx/plNu/xFclXfH3lu0L
AFWV2xAV9ltJUWSEdYNuUN1n3twAIHkwCsbswGBNBseWipWH9jdAidPUXadi
vOpPKpcheoEzmh3sjloYLk0VpsGRch6NrDduHhGA29RxJnP2K5aPDm1lTyZF
Dm0tPmVpM3AzWfPkEe+aJKDTB0OHy+5tlqh2mcBfplNMLzxFTLLwJUNunAwH
tp2MTQSCxE6afqksr4nPdY8pONA4zMEvN8ZYi/42Fp4MVgEfzJprZjhlQSRT
ymaXkQ+eTcngQvov9tyxbmrwKgZDi4KEbTZOCh13Wech1CDL9Hr1EAjuCpSp
WmFjiNN0rsyxEYchtMyuAi3tKnP/wZRms5Sgbm3ePEcbBip5wvsgvJrPMfnN
aZ18tELpyQjMcpayNlvham8Iazgat4JI2OfFthbmPmxEfT6jZoILJfrpkJGc
bzpSKkQqNxrB9/E0Els3aOUqETtxZXF6Pznej62lyVuDMl39s7UHE8bws1cV
FsNM2IkOihNe960p7AXw7CuAoG9FppNRgnJKBWwmAALA9A13H09M580SZZwP
Pnk4IzLqYPHU+kEmkAj2UHixi4AsPAexk7PqbsgtnFJEnNAgtoFpEiOFVA+Y
ftmJKcxYKwApu12IUWg3ITwtKgEUGXJIPUtW/C8ZJfqP9HSDgoDJJGSJ/YEf
qDbY18xufjm85Xeth1m7r9MDc2KS0/0GNQkXNHD6ImPNw9BypF/eRJiD5JXy
WiVU6YqRWIuKtDJNLMJT5FfA1nV3GiOATMc03TSDbmjNk1eT2SeuKVQX1Drm
5Eqs2/k3D5Fc8C8e8wTj6AJSqV3b2UPshw4yHvp4NmdeDmYfvl57+z/YYYho
yn3zYM0CaV6N6waRX7bwWLn1eI/f3/LUH1LlrVG5PbIoaLQsTF8kWwJEiyOw
YsoDLQbIg00C5xhXF4fQgWTr+dXotyiAYiD6tGFFO89c73aVb5YKo5espMMe
NHT6kqrxsmyVLn2DE5o6ZSJ3ywDP3dp8C4rAqHfiqKVTA0lrp90X318I3qb/
1VbWU7/+Z6pMIVoKY+HPjmsyCZ9pmIFT2g/8wpmPEabuH2VELh+eT/JLPoBj
HVoDL5dsRHaR34gNicPwHZAUjMgdkR9KLcX9PWYVEYeoy0v6dn2MbtRhoWgm
xwu3b0++cKcD0fi01LXJ3S3pTlRoNwJDLNLCtHJhr/yQ2Vgsy5Q0oj9ursaU
LsDntwVV3utej7EqPTQNI8BQjse7sp0Od94/Pp+HZaxWB6yLyjB14+77NUjr
EAMGEtlsys5UDlWhzFBTOCStjJvTKHdRvCxCABXjzmDKb+IY2ZHgW75Zn4lM
JWJ9SlLILTHiZdhHYWZ1axx5qUMNU5mmOj+Vc8nG+lVPnYGvKLrJwo98cl1w
EwitFyij5bGxl2tmC1QX0B+nfZaFWE4vPqpaH/7m+hDJPr+Yf78Vb3ScABfO
OGekI6xSh+KV4X0WVwxTE2BDdkOMzM2DgafDGUMNTDLMtWG7a63GYMutRRrl
ZKYPTJsCdagYHLzAHpNiWq+ln44UWiZEOuKYgRouhHyjUkYJW6eLM2frSFoX
L7g4CXtAKGAxBs9WEQsmgXd2D9IMeLwEvaRrvzeW+ABJRTZTPQtBe1SZ/LQ0
9ZWO+QNG+J2fufDzDZtQ2vnATKgNOAe51ugTpfz+yXb28uOnLQj+zBTfS4Qa
BuGdQFg1fQppope+qsxr/B1oHES1w0HEHb8zQjs6lZT+7ZvKRtTOAzsOqBSU
Bm+aHPprsZRX6uIIZi8ftI70yRczRKhpU0XOa/FTR+J71uSYiKsnUNeJKwVu
Ty5psv/fEsiDlnriK28MztYA3uckj7ST7QrgUuCe60tXm0Ih7sZRag7AeCaF
cEsBHwjIHcGjTBisCe6WGJnrF/rryJmkOVmsRTJzan6G9e/SvjelpGco/5Xb
mJqv8j0XjCPc5oqSuQ4f0fWSgm/ICBSQodX1n2Qo1JR5V9knAktvAU3KeARa
GEtgUi9fQgfhMG3ba8aPhlW/L8uxQPJz7ykIazUtcRpItlgEMZ5+pxbXSvTj
5usf8XnBc+WLiy622WygnPgK2YDcAa8kOWDxUZYbixvCjPLXzjXUKfJke04Y
VbWeadhCRVT7E9diRB10gHoYvA3smfb7ln5xEnhf/Pk5aRBBLhYYA4ElYFMU
CzT3zIlSeC88DaMv9hyRPRh0Kv4ft/V0Qzh+Ig+1T3VJ4tvW1K4sxAujl0MU
ceo3tFB2bbFvIJkRh+pM0aOjI6KBVgwYPxM9PE0ukXFdxMCBxfj6GpWrhM0I
lmhV2OqLlKG1ftZwd1w65JNUso7kq7konUG67N0Su4h8bsW6zN7hRWO4Nj8b
sfg7bpuC+gj5EY5snfETvA4z3YRd2SXBAwmXdF/L0YDBV1k9xPOX7jg9YUWt
MiReW8YIOLe7bLSxDEi8W1gf5yAfJdw9QSFT6o2v+phoei0eOmkkj3fp8VKP
GYbphiiAih3Ik8TkODeQl7/85yTvzp/23Y9UGdjKNJPsUJvuFVImFSEEAtIU
NLSuQt9NHXRgujqV0w+Rv/Wyf3Ti3cVWb/0Qpy1mO+1ETPLb0DYbKnufbret
U4O/2+U2PVhjzpeyZTvePetvHEz9TsjdKJ6+lhYd6JIsxkOGaAVpHZK7n27G
GNZMBYdI/lRYUGRxS1Lydjptun4PAajCuTkK479palSuDKRVmEh3tkNGT6GY
AeGZ5caD043Cn5FK1SiN5wat/Oihp89n7xIFH5rWbXyRqBdwMdSMV9A3jsit
/UnEb0b5PfRI3D/TTbre6zJmMnIohdMdoV1Z1UJ0TEJ8LQcKH4CWCBTkhEgp
fY6dCsWa/YGM8Sx+t3NJbihX2KGBWJi2qdMq4aUt/v20WYyHHmZIzFgYGnde
VAcLAA6hx4BVRlghoWYeVXbum3YfJFggyqnM0oBuhb2zPeneZ1px5PZcy28m
b8jXU2Te055uYrsCH881xLxOeAPvE8o+pdl+kPxe96dXWB1E6DPWaj4G5+zu
e0lVx+qdcdUzVbg6hgSAWjDzfNeXRp2lZPvBbd0+SSe649plEEgiSvQIOtfS
vZ8F5DPkkzTlNpUwk4qyAEEZw5RQZ51ADsy4rSfCo1yfxSQT/uTCBd7T3fzS
pqfFqJnO1+xOqygR/18fhCu69dZ2xT1xeKEo4fWEiPXrabJYO6h9D01NRg6s
nFicPvj7QS9+pVG8Fi/YlG/+uut38j82cUUkroESE08suD/SHyvnySu09QQI
qJtCkVtuGmyZaZi74f76MpJgIBcgs5nZ1Yu2B55vtEcgJYKtSR5s7/NiRGZX
M8QwfEuZYzl8maIG3IGWsRfD9H8978ZNioC4DpLbu9fadMQAzNyc08CQ9Bdr
ySqRn6yvGw1icqGxfIOGFmotD7ePaQ5O6r3fVuAFQm9EY+t1WrXaJIEytmQK
38NBzIx+iUod3Jwr3umFbRrwQ/I4RyCgKxfK/0UxT8coquXisyWpswMPeZnO
T6y6x8ih5zrrnfAet4za3Pi5BMQWGIvl9S594+H+BdP5JakrPRmeQUGWumfl
fgAwN+PNuMORr3vZxHJO9/fnznoYOfEuuYsRlm8nLhenX9uwBt/TSbUBgBh6
lLoo8nYNHW3E0SdFrumnixICAV4VwZpYgafY33CG3dIxl6hyImNJ4YC/toVS
5W2cdU139mBE+jKwLgr/7FBJiQx9em8/kkDR5E+vWBbPYWQAo+LRwf2r/CRE
T+k8xiSe/og7pQWyDDAIT9qrQyzm4wlghJSVTA/n/jn1dIQPapTdgMBPDS6A
eOf5I4m0TZa7FhjySzzN0o4EnT/2T3FjLWFhO4s17aJsnLd+qNQ2DU5vMzXH
+x8qBdXhUWVTjJ7iP6ljTgWTdowe9dERBQ5AJ5hP8EbPe0f703TnI538GkMv
4EuK3hANCAxIf1WRUyNPfd1uvmGjuk4NVTbrGcpbNNlQCIGNWknlzfixWqqp
EGKxCa2QyQONB6hunwg9aCalhQy60BUkwTbSQ2dv6+CthydumysTEX2mwh7l
DDvl77JoSdCx5cyGvZOKQVOYVW+M/LVK2n0RhNr2WNWzfCI615tfOVjwB8dp
DXkKhQQdRwaFaDX6exSHCL8CD7wyf25hoezgZy1yjyKK0wiGV0u6sPrh/HIO
uny8ilVhFETcYKWAEX6ib+PeZwPnD2/Xsin+k1iQ3Dl3fxj0upZ1R8yx/PAa
YgIAIwiGORF77eUsB7kGL2WvlSBWAA7FabZkavVRMvgzE/oEumFhqRityY1L
JkiQbjc02+iaaAkvUB79WexY3tROxy78lq6APekDXjCwIHStNQnbd1OEeJYE
UwBv9ngr/kkgFIVFPdFKdXy+CjqgdEIkyc8VNH8FlA/AZDFJmRv81DpRIOL5
5bVM/fkLAciI6EyjhXPXS+qulnPbSQ/7UzA6qXlNMj2Khe/BvDoNAy6TcYmd
eOZisfYEibmCobHtX4GRWWN0qtgotI3y2M7egQyAaIxJAu1Y34mOeyXKCNSt
uzbhNm9LOuV/+SB1EkQZReB6F+WWE80r/Lm2/AghMGDwDzh0Qp8sImNTb3XG
hfc5ULdLryBAnqVBrwJaPAt9YTxGJ1hFqAMPv4M/9cASb560khtEzQPUCBBB
xfhkBI+5xrBTOma8IfM2YN15I1wC2lgKW4MrRnBA0/9EHLHWbLQx34hzHB7e
rnrnl2+5a0ko0SDA13afknmsl8VZcUiJmEuEH6cPz8c0l4DhEYLh3xnhFR9+
pTRor/6ghW4gKcciPu6B+Pm+xLD2xUgpSsFHj46rexA1O8AmJmjNNoE3ra63
ybI4GYgWGcQ6N0hIK6BQMEqiEBykgjNsaH1A4acdQNXh+zUVHrLx6D8LkOQ6
kfn3fm6XxO4JW6slNLR6Alpn5NK8HuZUfCJPNGb9V17pkILQGLvAahhFPfgP
YdDP7DD0cCM2wFFHtZRlDQpvmBfgOCkavCjan8kWTXg3ya2w1O0r+aLH0VJb
XnJV7ZfRsO7YWrZurEye22LdG/bL173jsL3R55RJ965T83VvXpx9qnRP7FcW
+nf8/1r2MsJOXwg9vlwta89z3QmKcm2JrfezGjStP6cehNLBdUEeeynVMV0d
KyGVIDG0OK4eJHarULlJooJhT/Vj5ZLEhlZNqaLcIos8Qk289KaCZ4hkHtQw
ubeB7wGwUqnbz88GlXz3/WjaUBzpQKNJ/Rxz0s947nYq4h9iacFkL2cF6T2E
GwuqI5ZtHwzJi/hVQOCWCp2brcpsQxFlica+I4swzEhJqtY0xrBa+7fgYbY2
PdG17jhqqr7WQGK2wJz/4pf0wIfiGcFFibHVM768hjXXPvVTjqAxZ7Fh88Hz
Kztjcii53PMyJdl8Ya59KKMy8xVD4I6Qxkbx/CH34lBeH7BSJbUrUKX5hapf
Z1tBSqRgiJxEHAdyelw4zcmGCDD56/CpmwTC1YqBakXklj1NOZdbnHnh0Xaz
QWdAjPeaPQpZk+oQat7y3DbWg0mRIAEgNUBYlX7oBcJndWz5JKX7vk8WvLlw
HXFGa1Gery7q4nFiN/X3okwVIrrFj2CDznS6coZ6g88lb7E0fhoD96gRguHK
/OK7cq6lc+WCSj3ngrkHL8vAj6vYfjFQdWPNNbbkHlh6tpli4G0x72rut2Ko
/aPeeXwtUkpcsy+6UaF1qU4N4CQIn34ncGIC5LelfqdxK2Jj0Q8hE3YbJf2g
OH+0jWsR7kxe8Nbj+OhQ+xt/9W7mEPVI9eucxr3lZdE1kkhLFBe6EqLAEAYs
POJcQtmZjdTgTh8JB/953zuQHJM3CnaKFDVwnJY/nW2I6YvwUzQ9Tlp+mYQs
/CUIcT/oynaGHP0ariBNELnUT5OtWEOrOcPXBwtaNkWq2BwvxR82avR3CxII
8Rn8XZ3dh61Xq2r5eFX5m5wrMB7EFto4zb7yVVZ72R2iiaUWq7WZuY803Rwz
txiNwshWZIaAdA6yadt/qZgvKZ6pPTyPYFCpajsUF82k/Ivaef7v/qniDtp9
/oNFyDgrHeZ9gQ0LWmAWES+NO/nllL2oEj882K2z0UehS+wuOzn9yyBFi1kK
WUrl1+1ZhvuOQnUpT6NFHKIb4w/31h26gGdCN6G4Gyp4XLfDg1nDfmPmOsQE
i0hCiFsyMVtQWEQcCto2yztLAjsu5sZasKkbr7tSXLFUZEqNERnhdO+DPKkJ
RUjI7i9EzCJclzGj13BegXHkN8sN4vdKeNjcPcN2Nr946gz2tXgbc0dLPd8n
kHvLuPlLKGXcjzo+h6upHxBf94ejfEouXcy4nYxDIt1waofsLeWVxe0CBlgQ
vZFdaVxSs7TC5v0oQyJ5+r26rz22SCIa6xbw8r4BAf+cJ9VpAc8sPVqiylhL
ojfWXBVs/a5RGxmJZiBqgd5MHCyDqw4tW8xVwGsBpuUksTceWSSEO7GOo1aG
n9nbxG7uH+2kx1cEL1MEV4SHlm2oGQu7G9QHhxBwOIA0iDSpfaR3YygxiH2+
JPsWgvoGjeSgJfQnm/IRxfSrrxboxABwUikRMcwmYNJU+rxQmw82sZqYa7G2
/o57ZPQcPM5n3C7XMZig+9zqK0tFCQoe2oO6dU4FWMIVEZ4XRBezjSAFl5nJ
lY8JuUc8IfzCn1tqG9wCQ95TIgcFxPhZwg/CLEmEkDNO1nRJZs7HRo8ccGQc
jFdMZgA9Yoc1Gr1xT4+1yds0mxPwiumt/rT/Y58GtveVPuV1hcPg/8VFi0hK
HjoereSTtPskHDCCmdRdiKwUVTlblDQZddM1VuECtkFHYivV8Oo6lRpySWpm
CYvcl8VIi3qV87A9dwi0EzKSwTFMnt3ZXcXGCivKJYf0FXRFT8LJU/qpYEs4
j+bjuTn0OZEXzQDLY1Hf42M6TLiyaao9My7MOX8r9wSZWq/dTg3rlKDFprKU
QerfMam7MyhB8HMDzAZXzv2HO5VMmdTfF3YUQIgl5POefjwTU7OGqPMsdfJt
1aWxIaepL7CK23f6uZpnre0VizNvw6GSxH70OPHTK5uxqnkg1NHTARI69TzK
mT4hVNzxirG7f9shmrr3qaWaJdQyCprhklVvdgqkN6Dr+nbLEiGA0eWQk/+j
Jx4xDsFGOY8179hRgWtFk4gZsdEK3SNQg5KpzB+u6HhL9JBwyE5dO30U+5MX
3+CH/zl7q+/9+rL52lxi7aSmhVGo6fTa73fD7NU2uhXVTXczepCZX3z/tFsa
hkfaVgrCHVal4EuM2FZsRW9yrst/skoNjFbA54V8MOxrs+KIsuh20i2TWXSz
pqgL/W1ZeYktOE6iaY4Av5ij8LlhGoQRnR7Zrk8lL+BBBmxHoKI+rAuSGsoK
E6sqYx69QHtxP1t5+ptWyVrImZsrzvWXYzhlnWWXKeCHIxbhNHBXGlhUq3HP
0z+NTfnPfFxbWdoq4CO51CeaYtpVgD2jMHcleAniB2Y/QTD1XsI48IPSGgCw
6IR2wpucpqIfRknEBfE3Q6mqxkQ8+yXkOfb4hCQ0KDtrrOKrTMLe0maP9UHC
nkCLgPAchumYyqHwijuH0vs+qF8TkVAh7EReAEBBFhoh8oBsPAXJR/ddEETF
DxybfT1C9msE6r2vSiT32XANW5HaoS99J9zQumFMLH4MApyDw4c6YpmaQHda
WuglpWPg6KQAy/ATA8oGvArImXSP+Kdqw+2V+J9egt34qdRYAoWT91bOYnTE
QtMHiO9i2ud58atCbDTlfxsO0xRwHj8sW2tMX6OdjPV3MrnbvO5ad6qwIW3W
eGDwp24bT4T1yOrNUEjx9cj6DX5CMOyPTJKWhHuKsFYy2lSyWnMsjeUaB6jY
AgNCz2Q4iaBkpese1xfyEQ1O0YKv0kwmrIjHziQNbHnNb53SkIPLI55hlbQm
Nh0rDG+XD5/SzkXLBaJaKWOrQNlrl6e7p445+w/nbki2fw4hGxy5teYNBrgs
LWnhiZGn5AcUXRNPhCl2GXT7qUXkXpn4sG/q5uvBuDeGreG8/X7UTs51xYz4
cOo9uUTSKSUX14g/FeUS/h73wlNCR1rxpiwLEVIKgrJYMbjNnpraOU5e3nRF
Jj6PxXWAfDS8UfAX/qXEvcnW8OF3KYWm9xWf3nTwmRwBzq6Xgacs0zVp9263
1UFfMdA2l4D9XfPr8v1nluSPSRAysFXApQb+ooRVWIY49DkDElB++w84B/cK
8yqno/bZZKf+ujOMhNMVDS9WdvWb+ldr3DbO2rEtFpExN70s5vHIxZFemsZU
bmIyfhI+SRE9V9Kjxr5/A3LZC1ko/8nJ8+Tpo1c+c0KqDtoBne8cXLJINJko
7BuP2wqz/k3JtdNtJy3P7wnt/b4AIcXESYGTgHmcnW0HPmBUTx/bSAQgJ2Ru
J77+U550aVg+Ep3QSpITOAQxE4OWHjIlkYW4pHy1k9oeEKLkc/74F3oLF4Pi
2YeOnTBPF76Ioc4CaGzZP/k5pTK205pstN1Ct79DYM22KLKkqtLY9eS9RWfQ
33FZMtnARNnEVwNjvcZwQ5/ZrQiR/jLbHaJ5suG/GH5pI0p5JoAOwZ4SUGHG
g1QFIM66aFdx3OqpLNrZDAc366LCUZ0SjrAVqpQOMd73lEZLKOGnJT3oX0Zg
QffMudt8klF9h2lQJxUn4ZqHL1B4i7+8inKLG2CQ0RFhA6wLCU7dngUoPviN
VPV/negndqn0Dbqvf4SSI+vZcdQWcXE+PXPTSCF/Bwja5vZ/f6r0EziafiQp
jnFzuSG71lQdKoOAbATzKODByjvQCYJudyeoBD4oPPwaMMIqyvrvcxESZ1bG
BfhX37ANP03HGeqkobg0E+b0tp9sI3h3OEdTlhZfGK9xuMFnc82O2MAjMVc1
FIlazgFPQowGOjwLFcpIrmZ/TgFapzu2cLAl2X+jbwoG72sNoaFYq/azYCOr
VAgjiH9w4e8W7RB6u5DC/+AhDju2RO/ZyCC39CoOHWLG8nguBajpOJLMJKFh
o1qRg4i1NrBN3yeU5ckbyNi193dZX1/Rf2aaEvmc+zdSyUnpTCw/+oRPWFd4
Rkbp2eqfmf5kQpIVjFp4x07XqD0DGkB+yZo43ycFymzcPN7vqiRH+gdRKnDo
yFHtL5en+nysIeJbZktN+Neij6X5hjUmTYPK6xbZmQVu3GPc3033v+VM2rj2
hwLr3cSH8d2Ih/rQZDW+VFXSPm4vHvocRB3T+HZ/hQUeSa56XkhXC1MnIz++
MgY7oDHxPtDv9m05NZtttCXbvsgeq2snKNHOymWbrOOxdo4s1O3nAC1vB5o3
n6PxwsJ2HAV2o7DDKKaQC3HUap+8ejsQmJmv8nV4Fz6u0KTnQB5orc20bI8n
4ZK4fG8vCHQThXvFuSUxh2Z7g4YoL9izAIuFx346qpXf4Y51zDZJ8c828FyQ
AXAuAX91xRazSNTb8esbQdhk2gLE0QsrZ+gEu0jlToxfxhXE2HIqrYVJfIu9
kFoxyIIdhWG0PskqTzQcsgSf07q6VSY1W8VHfdBw1KrADjXR4Rt6O+ombLj7
qHY4Vk0TnxH31bUaAq3hnPXscNdLJouSKINzeliUOxfwzLvh1SdqpCgqLeAu
uDkgKpZf4Wz9MaN983+sdLy2twGL0WpviPB6a9sz0ld0hQiRTMKT2Qp+axR0
qQlM+KOyvq5VPmyTzl1X4alQRTPupad0HSFJFJ3E50tq18LnZ4K9X69eSDI0
ts0qC8bWkxBQ4JsVyLsQ2Ucj5X9JhMhrCJGnKbSOGqnSLG9xq06rtv7iPV6R
sfF4LsrUplPypMZuU9T/Ync2qgSWScXMA8VUxufTCxjVL/nDcxr1Jj0C7vjX
kmxhXpRtx9A71eKGINuFOV4HuKgBnnTW/exFpa8O7cfkuN3l6IIuXifjaDv7
tt9DPFNZDhw1T2pvyuiBHxJQHSvVCc5nFBcLEA/X1SPGftFzHDSC4NNKMXq6
JyJHXunC7BqM3hVqMrzYi3jALa4MwqtGGxzvUKFWrWzHjU3aHccHuE8OuXn+
fRldBct3Tb59OidAY6G5YOoYOCoK1YJGeOlGGO/Osz0vaGMkA0UQBgtV70aY
2fm6Guimyb/eEy0hhIdWFO73PlsYRuHlDaa9dJsTcXoxecqHoKaXN6o5DZCw
+XBTBkUqmSLMHcjqC3IBkbhUAQxcmOQF6EeNMU9vJjUgtMrqfhlaxG/SnO7f
ikVyWUcJ6NVKA7NnaUHG4R/Yhot2egskX5T8y8IXceyKH31rhAXyx489qTa6
8JzOq0UvHUY9uMisZF7A3Bk88J/o99AQDpDDQfHLaMSl1xQqnHyP7bXWrGGs
JZDRNbSbZXQJ1QeKWK0oZZEV4w+tWwWQKl+i3WWKRaHoQL8zRwtnAsjD8wxt
9q0ndtiUQvPcs9IjZyMzxicKLhosh/25Qh6fjirnbeixyko0fxR51Xt8wafM
go/mSg83mnW+Aqa0sosfpq6Qj7UizBTJDkUKVS5C1T8jaJu7wxowEaGXXFp1
dMTOG/X1/nJ01K2dF7GfTwKwlAQ7TBrO5vvc8qRzYGvbLeviGTVTJNxtmfSx
PQDqIJ2S2O/2cN4l9drnVDQPuwSbF3FXMVFu4mSn7hk/b81PqjbOOsDLJ0wx
zmrj1pnWbhb2+K0Hdmjxl+Z5iT3j1T/2C5HupiFYJxEPST4XwBYrgpfiTGqJ
K4tpuQsq4tdOizeOSJwllNTq15/jUjtT4HqhnmR7CD5Bv9YdsCuBcUMBAYk/
WDka29uvEjx6SdY1oGR48KzCO1Q6hZDi7SM+CuvdlDGhZxkNMwiFhY3oFa0F
F/ETKcxFjyRqjgdv69+m0QA86hDcNBowEYOLJckMVqFVBQRvHHEdkItmVk3d
mfcn+/tId21WUhJjqNneAKl+p1D/mUvN+68Hq6Bt0+l/gXVWzE6Hy553RWA6
+yeEUFuSKUofCY7LH+td1c+X+9JN5UVEDQwHZEiV+GBeZpFXKfMp0lMedY2M
iOFijnvgX9Fm6x3ZY5fEs75I+RTSPfJBz4UIYvQAOWf8CmNJL4jCaSSslFG1
A1vNefAWwlD4DPL5YFNi61bSZF9DVB7ikzM4Rq/UHg9MLugKQrD7SnD8+YOD
efiT/GMkJbsmemVn0hVPGQVFAZip7U1W97IH0+74+Hyu/tTbBZQjnYivkLs9
/G383bt7qTf/PAnhxoAQSJjwcMUqwc8JlDQtE5bjT3XlWM4lT+TFwwnP2uEk
vsBZxE+ipZemUEnWynje6nvizOtL6SvGsoRG8HjQjVEchdfov7OpUx9zIK/3
t5RK6LkUKzodYeMnkXiudRxrYG/oT2zXbAKgDSi0fgaatk8JuzE1/RZdp8Rt
b9VhA7/3oWOKSi8axNlPA7QzCJEPRc+3vIq11GNv8DNIhpXGDiXLr9fX1wZC
tT3yjgU58cs1pL3Hm2z4sEdQMuHHVIorF4qHlphiVwnvPFd8yUkya4Xj89Gt
p2Eg/vQ4lRdZ6cOWMnjr5BQXAlXQ/RRV2ZnboOz3xm1Wlxebi5drouxRM9ya
aboeXxfqTxGNFpy63c+lcXmS6wgzqkg4kyyWgIa56kasu/NOmIYR2BgAer8W
wHVz8B+kNAk5HE5p+JDyx8QN+4O+Uv5oI60kkIY11WCPMf+HNOAEjZO90CC2
FI+NFnb8XaxU/d4E1FlZ31wsftHiUJeTN25qR2luTwkWnVXpRQ+R8eX9cOGD
XNymE979TDFKbTD6Ix7tV/pUzwG9wQTs/UaIKNSFhg8P2rcYuWGnmyiLuAM6
mEKbXUutZQHrlO+Lhv0UHiR2ss3ilsQwoulUfF9Mlq4hPif+6usCOXzXesD9
3TO6VWInsD6GJYvaYKP+3VKcRMOa5DpHrqJE1k8GmH+bqvK9A2pSkihE1q7I
LcKVK3IzY3r7wzSR20hnUa3kdj5z/cuAoIwfNNunHwztkxanB0eX2Xym7K/G
KTcb1tDMGC/C8MZZ1JwLRiRVlKfA+XX/QSwvD5d9Z+UdX63mCJYdlENF7YXr
+jHwQdeGTMkdUtyUIPA2F36aZye8BzA/vb63hwH+EXxsxFlGfB9UQ8N2Hb6M
jvQHmO2aRjGUkYkWTqVCCgvAOaeXKlHJy8/UGlSTaxzTqciJDakgTiew188G
0xnHh7REuLL/ScVAyLVq23sjhP83lH+tptxRH2DrDZjVNEl24cu2FzPtFj44
hXOxLnWT2oLI1pOxOfO3Dx3HOwiIuXQ6yxt3cEmlkNWEy/vepAODlhIxkZdo
TanHTPVxs2STYjjG3/zRi/oZWWAx9lIRL2iG/JwJpCM0OhSwruInwlvJIpNJ
kmw5M1LiYw4wEPGxpKZ7wMMIhPy2Jr8MHWFIuf5oUyEXrPCgQrmJGR35ALkh
HGzOylYhDvCoz8PnojZ6psqim0dVfaCBTRDoX3ghQzoAYIwRWJeBVpzzNFER
w3EpPzDKJ2oyoGjmuGpkATitUCKY7fNlOsyz8T07L6cbwtL5T2YpOtrR2Q1J
m9M9m/TJg93m6juSGg+asVTeL+/ymV+AOAmUm0rKvwX0NQvORulfDBY7yC0U
TnbFe0QBgxpGUQYIW2UeVbFOSaZFxyfAe41AgbTaVcja+vfKw9rI3I1E/P6x
m9inMD5rqFpBKMxJDb5qITZ+eTvjiYwH1qmv64vsdxt+EM40qexYMixm1pPw
ZaXzMLzb4JZJbSrMBUfF3VaeFySRsXecxJaFwpsypJ0iVrJl1pVdp7mbJdaQ
u/3+k2tSKQI707w3tDzyNuVn2O9dCMqj2wJsxbnQKGmYrbU8UMH4KRB0I/9U
qKQhuXcbRBbmBQp8jGNnhkmjlHp9bXqFfsRaW3LKCdX6/7sUOMrO7WvmJ090
2S8NEuknhJ4vPtrv678BHdvYNSGy9vvRJyDmkSMdNa1Gb8z7+ejHDPUpHbVs
WzROiFIR5MTT9BNya02BbVnMf6Zr3BpzdubvI2ecImsPaHhrAuTpkn1oqLNS
mpGv8BGQzOwaFAIj9juGLBlEUVKancQ5q492Pr9+DxQw7fsyP2P5d7ZONrnK
HRmq2rVLeZzPVpPxpXIDz/PAErJOd2M0CVMwW+Huv2e2RX94rqdCs8KsojOF
SpzS6CZ2Wr0Kr6gTB68AAnhYYkqB4iZGo9aEmjJn8xdaQdi1v+aE7WwncOVd
Iwx+sZcxzYBOW66ahA3BWYPXrNSl063uKmQkcE+hn+EBcUVI04J63y6AI+8A
aFO6vzrrgH5PLjnXWiXXan051U9HsRfyW0hSiww8WWtAdeDr9iTG2eyvZjuw
Q4nVVin/0gFSzwadC/eq0zTYcohuByeyF+HWkxgqrcfsJIfTyf31z3SWRTii
46tTG/x3qUNofj4QEOhtEtOtaFzNZutYrOMEmzT95VVnfMC/ICUfzo/o+XZ/
yrZaSAUZyCNGgmhiMIbdYRPg+jla/FzXeaCBS54tdxW8E9P2Y3SSlaMsX6xQ
g1nWqcgo3nNvKSywPwRZZfg5zOhSPgPH4axDWuwa63/2Xk2fNvZyi1l3giom
im/9tVsLY8BQKe1VGd24qdNJvaZflvAfIip0O9O0M4ZKSzdkDFayQHWm5LMK
7cRdDsVSO5KYwqqzFtv5r24gMXZ+gITGGxiSV4DakgZki5oSdHTqr5XQtYgl
QoUIht1hwltJIZmQbzWqWXJpwxa48UX33VssrZnEe2usa4jEIX84GpvxV1Mk
/lJejwN/v6JgCZS5TStoAt7h+MWbT2HJNIQack/oNhtQlGaM3kYMrXpyclti
iQF9MD67/kxFE9NR2bVMOIc0+SjhA8RhRSHnOBSpjYJwRVluX8AXV0ot1ClK
U3UmPxpKMuKEVX/1yBA8+CmzbC5d14peFre2Dm87/kXsnkulxwI+a7lBRuJ+
2pxND/t6N4Cv6b2rLPvXci2ZTf8/4ZVpIxZPxHkArsUBeKhYxsOf57CIH2Hx
FbsZTsa3gdTzImtjaCn12qDo0xDhBQS8XXpi9JbyQnx7y7DeoGTzXV22U7vV
iRFXHUaqGtLBfecNxGsV4i8XAAA7q7l71rBkHtSHsiC0ll9dfSJCrbNtiA50
Wnr1id/4BU18oJVmJtbc1tvR9pdRJRNlYwCfE0q8tNJrU37hdaXz+eqFYRYN
KAP7UW34/zBdbodtWf9tyz9Gj+1A+chXLB97WkrqSWQhWGz5xow5HrLjbRjN
EkxCMT5H/mnTRPWdhYFjPwXzOX4sNT1gFj1V9GEeszcU09ECdeErH5QyNioE
LSvV1P3lB4PVzpJ9Kr2hCk5fNY3KUGNGjY6deO/huLhEmqpNlnam5hSOziWx
LIiN9kavMVA3l+nUfSlYUqmhprtfHHZWMxX9ZK15+irGDRI6b0Kaj7VWxTt4
+px1i7K/uiRPcoXOhYR7G/tDNeTSDDHwzbVpGeid+6PE9XtNfcQET23FC/pC
ZiHYvAyWnnDhcAiuPdRd3020cBKlt6NliGcPxMBFYOxFMuDamT5GiElZ9L4B
UHRWV+JlzpMaxxAwqTvD1CAvnGHtdCqCDolMcolNtRcmQFiIXHE3DEY/0chS
TqTj9Ji+77g0d4TTBMqXC1lhF9lw7LpGbOKc6LExxeBCeHfhsTzCmTTGpE+8
Mjec2CuoGwqpw4d9A1r0ESFgBXy3N5lQcZEUMZyRtUt/JDnfyte35mn3C2f0
txsM1dFxfAXHT1fd8Eql0sMFGNDYQfkS4FIV/tQ4vm3PSWdQuKMF9dXwGhfB
eL6n8pqwo50vCEIKAmdwdvuU1NtpqHFAcyiBtioFv99Y6NR2tXLWUFIPOeFB
B1DQdQPSzyhReONNXtnmX2AcXCa4omP9HCZjy+QE1PrWrmDgL+n4GGO8OlUD
YqQipN899oDAJY6MFrQmdYzTjZtIDlGWorHyWsrykxn1LODyOBkr9JBq0jPc
bGykAxWxRZPy2eIgmgJIJa+SxpgewrkSj7OGxkqBn5InboBxeUDy481yx9fp
Dng3fYy5bFsWMWYEkVembZ+ONAXHt7w3H27008QlD04P15Y6PWa37Y9EnaWR
N8na8ohQrZmUGM38VObkbiiESV/igkGV1aKMeQL88saL7CPT2J7MRZ713Yil
w5BVLoareIrwSA9iZRsHYjxQ3AWPPKKAUiIeRH+dPVHLe4XYoM4VNsg5450j
SNmnFqnesHiOh2HGxoaUBXFOlFCPfQlmgBoUcaWFOP9c7YrP3IKhvgcXYxrP
06DYCFLOrNncTDV96eCrYa4eKGljcHlGEYqvzWqIHyMOPGnrweT1QFrBreIk
vfPv3lltm3IIDpsq+4EaANgYRQX+ASaRUcM++oP0BzaViZY8tMDWyByEq+mx
opVDxDz4QSVes88f0V2G5824BOR+e7bscmwvu0isMRY2QCCyhYH02gC8G672
ZRuj84yBqYz9Fx92QbSFqfQU10aeMO9jXiO1tDMPGjsL2iS+oDFTei9Ms9Pt
HdzaTqNs1pZX6Jo8bxYu8XQyGvQfJjGufJzKbbTrPNJYyJAwl2x2RgAQaRqL
CEmkk7QPQTNuLyg2PmBdE2WqqAPK/Srq0SE2I1lQshrJUIJCX78K5o1mV5Ou
lVP0sERzhjzXfb7rj37rQSuXrpalASnly5xf0O4FsdBlww+ACRkJ+idK8awW
n/JZtZyTJnTzdXay3TBdmtkp3ol/OnMNE70zwiIUwrMYxRNfnQ8cizua5jl8
yWfTRf91VyDLn9k1HpeF7S3jgtGwrMVUJdLQb6ODyR7R2r4Z3xNblIkNW14E
wV2CjK0wTsd4H9DV7d1cRYJiFUllBTbYZlZWReWfh1hmN1VBTqUTLN4l0GOW
vGxwUU2zzN0JvNqO4XDsfFqcdHy7TQqjCuNeoW0oZBREfhYbT+Uf9ydlrYbd
I9DVW+9Bvpbg+1Ju9vRLgUitGMCnFYyZLq7NtWNuiOhGIgLJrBEMnHGYMOIQ
7bYsFcNaQSEQukDNvZz0zbp2/skgeT1SrD9sAfikuQ4NzAsP/7GUZEsVpmwL
Rwb0k1dTRTc7/OJi9E4AuZDS48lacVIMPw42zNQ0UcHxoXOSSAd30quUd4lm
4cr1HsIflt9ohu6gVqIK20wbG9PF/gV0vAQOe8IM8y2fCUHuPwxmFJYU8paq
n0yk0eE7PJpU+6BQxZNQhQYQB+7GS37iNyphEeYzZj8uFzV/5WA3axgS3hJK
F9vImpwykivln688bJUB/UWPOtO60/rpSPg3kU6DIlG76yeNaXgfwB8CvljX
mbHqK8pRabJyg/rQ2NnjPuESlgQr671Tly8yfTHwMHuy4mT9CJq6Q+9Cvnux
14nfW8oSIzHSGT7O5dixYtotckJs3nAho//vh+QbhvKiAwQfYORJo9qYZWI0
BTudxKnL6OfFxrmO0/8f1DlOgpsffrHWbXAo3xuV3pJXGw4LXy1o0/K7CKLr
DmB8ZHS4Lj4soHGCmZO/9as3gs/4E/RoaUbziKeeM8+WoHqxYOjV/Z23j1p+
hc1/1u6O5dEIRFpuycq2epcslFU5FOmwSLwTpJHY97vBNZekdgklsBYGCt/c
/7aefKoXvskkQLY0u7mso389D0PBa612aug34qUwFmLyQSzv8MzudF2Vv6k2
jz2cAeTTrw4wXOUpKx5hYsKVy86i2luj1O51dWyK/A7W+Jfi3GogLP4mVtkq
r0BgvE2jVTkVjvpnghnLUrsQ9UsubjOIHnuzgPDSytYBt06UdVDxdAcV16zq
GpZGvcTp43wiuwZZtdi9GRZ4/VpJMeUjIYLjhuW+D/d8wm7YJj0WoP8Yikiz
OoOYD/QIyTONojzQbN7I9oK5Mn49hfQyK2kmiJK/QRbPR6MWVc41eyREv7UD
36YNdHmh8a27suCjROhEfjxlUuY1wFF29C5Suy6RKE3ZQWATtOuWUqmXeE8x
NxjEaE7bc3h91AzexqI/lfwPMVCp7ibR2W7OUIpc7scj0cqQUo9/6kIAl/VQ
7Dt/67yspoxDx3BzFJz66sjwQjX+XwU1CWQVRPGsbxOmtiWx0fuzYNJdoU8L
Kfqp/IItJWS4HeWykj67k61iQlDz6QBmsdetzHb+iDXYSKhx/lVsEOG1DjCv
xjvYlCIPGy2Muc0wMa1uXxMVDBaUbOEXj6fkzwUmH+EOZLYGFwWnRWURRW5n
QGAFgo09ZiiQaqvu15nsFbiUkk1N4ACIqBe07zoogr/thArE657A4fZDnd0F
ZH0JyCWOzjpVfuZ2csN9lXS9R4Jtkt7yVoHwyf1kaGxVXepxM7h2wae9mf59
+OI8atqS3UwKajdzrAgQJEVe81fbgc20T36bEXbiGqCqhQk7xMOYwfMp+EwW
KzNi3kA5/yqkRJkgPSx23ACE5Wi0rK5SdAh9umxvtlHswXhf8mjR/Vn7434Q
kiW7muiWYx7SUfMxtWCY0DmEogiTCYNYkPQUXYN3bdat0T004AO1E3yeH4E5
HRBjQiFWNb5BSXMyGbTMTqVclvBeduEI7u0Woq9OcfyD7nHc36z2oy7ts+Lz
6mMvKjUAPVc4M6WfrWE/UvubDT0WYx5GQDpdLLCvZ0AlpJv49K5nSsnMJSup
glWKr6ySNlLQe0frwRqAvu1DHdTnKCvN1ZdYZPEKbhs5UK0U1I8P6T17a4en
md5fa5a8wI4RNoFGEUL1vdnhzIEdEs5MFHLmu/e3LCz3PbCYtzm0EaciZ6jY
Ep0Ca1IxMVN4jQkF6dMlFy5glqJXB3vSZDUEEW6xFw/aOS7yMIs41CJB46V6
RkBmcFSd1Ot7M5giYR6Luou3Gnd4V9qoqpJOJBrACTH6PtPDd4uH/apgdbQe
l1ND2up4k3qQfhtO+Ze5+b2fJfMdx1B4DJ+7FjrIRWz9db3dBk57lzGO+I96
5RwhlLveNNRzPUg+vd3V/yeiKHWFB0ZhPahQHqA2Xnd5znO6RL9j7BR/RdG6
hkQ2uW1yxI9zgFXyprlGyygFspSwPQgSJg6JtlOpozta9y/kBAev5mG2JuN/
mg7AX7UabeMnZ2JXC5LVM0LvyRrMF6b9LkzHAfJHESQRYbu4RUEr6vQ0otYY
QkL1o7iwY/NcmUXJre5no5bugZBxbDUU4gokIx6IIp/ZHZ0kYB/nwF8kxs86
R2ERBNXLP5yOJTtenAd1Qtq5n9a5iPrethoGeeAJJwwEjrPBYSYWBQzR+tIh
BpFLw9/PiUtdK5e5mkrzU3zIOtJ5IXox6qGyz+Wm22knwO7h8iJpsqxF7Ock
0lgap59lCsizqDaX+YuowpxjBew9PgGgoIe9n6EBvnFguwfwDzhe3T20HdMP
kfh+JDcb/244nSk4VY6oB/x3La59sl6j2QXTPhz1c/0+6I7Nm+rzRioq0uxi
UG37F6Chd+d5w7ioSBoJ7EGiKmu0MZBCV8Q8ymbMzb5kAMrEp5yEFUGRJbWf
zxdGKEIJ0tY+B2chETb0kJ8xLPh6Ra86xWet4EWMmV4Iq1xwBxcOVTkyHguA
AeO9BpBMjiW7hSJisjeRfjGQIddOFKU2qbSt7VIUnnNvoe6zRfNAPJnqR4rV
tPgeiIOuedrxzdvXDqnCnrebEreqfNeho+xLIrj4Gs5eSAMKVtZvo9YoGuEO
9xj/H9Pppe4tNAQTlVgkb4DlgtBNrlxwYNktw1YaOuDLT9DoXP+b2JljWgdP
Qdi2RGdMaufsSyk6HMnqxW9lkQHCrdq2Q9BK8Tr+YDEd+C2mqsf25ItYhEqG
YxyxdWNeVELMgW0AJsc1qsSomim5LA3SZ4L/UBeS+aSm4isXG67gxyXlSVmj
/AMiBEBFTpPj+uRepTSyP49EH2O/wzKGc/UTkypx2+cjUhT/CUxT1hjxKTnS
zJBJtQ6Q6Sw93J/dR/wQf6SD2ZsGtZb1k+GYl0Y0YeLi+RiuHEVZUhLYsWdn
vYUD6ZT/0EtJs57hkAGLu5qV3V+GIZtAYRh9XnNfuY5DURiWMqPv7dalINkS
2D3AlNjoSkJ27ZQ/XYQzr8ZPZeChMMxMMOgKVTDs/QWlnwohUA+F4jFRF1W5
Dtmu/d19J1yXIZAYRrhccK3+t/wx8J4lv52kaTP1yHAPZsgfhg/BmE+uIT4j
2c0cX0qQ19jUSMLXlOQfdtRr0lw1KzgD/qfLve4zBB8iN8cNKn44Ev9ZOffZ
Kr6vaLZmLPbaHRoC+hlClZYWvRigPja8x31Z/aT8ngV5cM/IJeOIbsG7HvVu
noilH/Co+JRacp2pmLtxS0WhSoV2a5WHTYsnrN/BZUbEtZFWYAMnrO+fqv4I
Hrs4MBKX7L/cEbzT0iDVn0+oVcYb29u1g4FJNolcrgN1Nx8UALAgeniibwOD
24fybUbGM9xDYNjc9rzMjs4WPTNEorW9EeCJ9dUBemz1kwdjuT6+FlLnALb0
QULrqQ9/xo8InRBri9uEXJnyDTRXAfH7m2VkPeCH0R+X/F6tJXsx5rz9fC2w
y1Dil9aN7IzH9vJ5WJSCK86BqE3hVRCsfptHRnD/Q5y7U0woBOU+Xb+soUCw
GWpQNWRZHasXF0Wg4TQjBUIXoZ/XynFa/DHsA/AnjZghVlmnpdSpNT5Ieejq
ega3Be81yJG7/0MFJ1tUA9IH84qfRCHKczMKuM18A+oOB6/wT1ZiJV7gRA0O
XPw4ECqDEpsNHnKRfePGIDQoCp1y6JYciiGsKy5CXXlEdPMkvJsDA+0gMip0
aECyZ+X255GkQvJHYsVRNLYWbarvGUB//UwH7xIB2dMrA1aMwUW4Q38R+jov
LKPsCKjzngpcTNk2Gtpj7G6jiqddqYAOrHQCjFp2VNhKFshzIe86Aln8jJi9
6LPkafo6lL5reFBbSUmRK4FWP6d2eIjitoexRybwp+HhaP4ehr7WqYiV0R2t
HZE4uE70O81hk0sYD0zcA3ornZVZltzaVUDMGplI/PqjLl05HCZwxx041Pvt
rpeeR2ybUL8bFC+AW7U2JAv/hinQEQkwR+ffY4vHL9LaT2stJlUTLZ5UI7B1
cibVYzhXLYvCmu1G2awkWnJZ3jY69S2WHCG8c5g4RPMB7LfW3DP5AjrRvIW/
FFeaE5kcnYvxtIzET4vz9vNVqkSLltD2Eg9sh894V/9ced0in4GHBJwXfEiK
rOMO0oopWrSRA7XDrVfspugP5ZqDT3d5Hhm+9vdxwJc0yfmMmUZ/tycTE43L
UJZltOu5ZijlugkbDYzJvCQh7+kAD90RseeNnj86QxcXpLQCSnR93QhIrY53
e14H96QFCppDdLf4J58WVf2FyrbIhaCVkBCzM8bE/Ms0aMHb+0ltTuQLjK0s
nyO0+tTufqCGWolJkSY8CreuvfpUZB/X12S8dQ7QyN1cSd1Fs22JZ2OlKWNk
5Oqk3WQf4iijhg3IlcYWEGq5/+yabEQh7sFB+PyJ8gZW22OcWhI3RYUYS7sY
xKCoFywdfYTx5minJFqYA+gvIwRPIAHsJD4TRxLgYXxZCGagkDi4z6RQuU/z
6Qb1m9MGe8vsmSqvfBSgeVRIkKWcc4015sf5GjJ3M61a4at4yx4eo+8j3mUy
StIkGqgEk900Ii+Qbz+J2vb8mK3zniB0MEDibf+K4Z+859wdcseTpr8qv7V9
+v1PE4b+TBlApjMjf1ngpzpjMk/BNkxLF2MCvYEIU1X+kaTm3a3EQTkj7pc3
zafB923PyV/+CSy1iHOSeFJ6wwpTNDle8whNsK9HnKZIrlNcS18SG4926+kj
f/ZTY2wd+eUv2AkbAxWVkT2Ynz05qRTXeuye1+/uaoIH4xwol4e2+pDboDsQ
errVHZSu/3Km6HA6NaWDdhlUs9+oU+nhAls2Jo01VWfAsuvDycsFf6B9wTZD
ozbdM0d+DBQwzeYYwUkvz9/1mBNciQRdU9BPhIub3OnqxcXBQ+Oj5kJ3Fjds
gPkJfUa5ModXMzpQ1mWbo/8Vo7oyK0Ydigtk0I72hgmIsvIfzXbM6C2TsX/X
5jnZx60vsDIoecTukEokkc5nkWzl+RoQoysKtKQjzQBeB7StyiFBlrC6/g2R
U1otnu4QtMxnbHxHBLmiKZqbOLCdTsIQUMgLSNsKzsA1a5hpd2TpbWUWrMvp
EZx9XlQS5MaJM9y+5/WbE9ucLkzRhGO5bRQOxKPHzopQ2kVipFQrhi4W4bvP
B+M9TYP/eiN1gVPzPabHXtinAUpv6QAWOIluSAwrwyJJMRHHl8D6xV/NFg80
x+cjkGTZEs3j7k+qL07iHavUaNGOYU11zzU7Cr9SKlGTzJLsxeJtvkHLR64o
YgVRo0ywhdq8GfEHpQBJdHUjAM4qrjH1ah606QbYBx45JKQq9e2oGACIEKgw
F2BGyuv2Tl8e/xPNSCqlnQ12wnp8+BCZRRdZz1yHbhrBW5CKfLbe+JqKAp4R
uEVl9n8H/dy9uSlaLtwhdx8LKKlZs35NXt+ZJaXLVQqDlt/xbNoSe0G0+8CD
sIB03YiwOqxIxyq75hghqw0u5N0wBljE+7G0dlLbUVdkn4iGrdiQJKy062/f
Bkgn8Bg6Fn4bYgKkgf7s1d1o6oC1PY63UZgLNuqUpSvlHGffUrhqSdAvjgA1
XlRw40khb+iM7z3FMIUeIA6vn5sHpS35TeVSIoLmFKGEULK6Ag1jnJ58utYT
rym5k+2d3gcNIU6YbO1mNoPZtT9GSliWFGaOT4em4q43ESNjpr9ycuaWi/Ov
zqHYT2dal1mJKvmBeo50L2h56W2BOErFZ89Gm0g1p52qu8RGpvi2se9zrzmh
bBdWMa6KesuOjt1pKp8pdx9FlabbifkWQh1JgD1+vW9zIwP/qX+IvkAuxbKJ
2wOxTD71FnvLwnrzYMLtkiMF1Gd/YQHsnwZSv73Wuq3KVKgMK9lFbLQzh5vj
VudcezW+Bk5k5eJ38lP+aDOEZA3XrIxjezb/g/l1by9f+8vmsN8EmsrxPglF
ORG2rKbHKiV2nkB/vI4d6Oq1xtY54kimq+KhibJkmtq2W5HXgYsgEgBtw85U
n0IYwIqwSCN+/q5Iht2gRPn3b7yJc4ZvrBkMawPn9hIKl1w50Cm7koobTR/X
ZToHmn8vjfH2gEl0YIsVoJbcvwuEKO3lqysKB1gBG0ULADYhXH9NWv9gEnUZ
lIaCTQ4zoqCQM8AvadlvFiDSCkpvMvNzS1+E30pG40GLcBS2tGvffq4mQ2I1
EplczX+41bWO6IZc/CfJnSY7itmHYsuVIdKbyZnUq/FKTbpUXNUh/ykZIJul
rojaIYEWzViuQ8UOsABJlnQ+E9qqRHmjv91jwKkkTRjVbMVPzNdF95+9xZj0
7eq6mMTwWn5rEcYKhltyuFcRlDW9/eOPl5IEz6dix38+Id62ONMXaxfruqiX
HtnqauM2+Eb7olRHYzj15teVMDy2V9VRG/To/6rKNff08Jwk7CpIP1zVzs98
xKmoQk/IPSMKvkcAQ6wvL04OzV7VoF8VunMYb6gsJNAVRgvzeYfXFGrIfzHo
cCon3MOFa3jxPPfo0BSqzXLE7dzx28FXm3/1LS3XPStUPJ9hJtncfT106sLs
SaJlKe0lADmGkL65TvT2B6NwVeeeILLmohyB5ia5tOM3+oEXbodcNxYSALWs
HasB/UQQbYGT4Yxq9hQuYTwVNAVUG5iPOKN2E2YXu88aliVLhQdSVqBGdvdL
2NVwlfiy5Ezs6Y2X+64DAfyltzJBq3uzFUmHv7VnQ/EHz9i81ncZ7rtgvEHO
TW8Dsaptm1Qce4oh3XB+lBo8L59EZAqw6Wi63HFfH4CSIsCTY94fHKzSgDFQ
FyXjW0lE0C3IVTst8GGwxcMmpHR7sdSlESBSMKMU59umugtxf7cKl8Oh9cbx
E+tqanTOFmnUFwRUvTGTUPM+37W8YZlPwjMIKfAuAh/w/oIkJWUWFtl0B2FZ
xFjf6bshPVDSwlCvOSbtU7+UcYtQDRcqF+/yMQ6wSE/iTy1d+wOcdg5MHmri
CyckiFHwzf7YZW+Kcx5wsFH8BEMH8Ib+ws4fKS+LX2QEnFZXEQgZ19k/Wsk8
5KPm1YY8yIUQC2hHlizWK1tgwGzW+7CKhWewIfTTIcCaRZHzipm+CDvVurIC
h+RYjAxVF2rUKvL871GbxzACwkBqmlS1GXfyxGLIUvcj7SfMdyYL5CaAzR7q
A22nXfd3hu9FbDS5CdQQ2m+PnFFQuZNtATOSnlMAMLxEU3LsErXJxX7/3NaN
dHi2JE45zl0Nlz0rnBRmB0J/NPQ9fMA7SBRwqan9H9BVFtec2RTYWOGRcdh7
ZZ3kt3N9QpW9mW96ZEwfe8dKV/2r8diljWD3rmoRt/w2D16gZtRBnlhv8D25
GNfGmYpfglRA7S75XOsscVXP53ZNjidkByXgXmolP9oSliqqoexHIMpGMqzh
V2+4Mlry2WvzJe5g0wfOJ8eNSPROuNvGS2jlSPAat8aQVOxWjBBfk8h/tZM4
2shLr/1wEJdtjdSBZ+TyFSU8ARY32nYLyCzmCRTBku4kBEPI/WP1wM2E3iNv
ALGeSgmSJtTQeIMMOCGa8hKhxCbqs2sfBddeiNlSRskIvFHAuEHSQS7+nngE
bD+bw0vco2PBc0egCh6zQ7KBDqJODZNumC5If+ixvt8Y3dCTArH1bRtzEQ7f
jfnavMg5y652Z0YhvhnxNbQfjZwq3OYg61BaxXarR68duKce8Tx8Y9B6+NlA
lkRS2fl5AQPEDoNmE1nLz0lxZNX+uUTVNgNzeBCSaI4VlYr5/Yccda0z8Jyr
DjnyZDrQGDS6bOvS/wYAlzRWt30GC/egc1sy9ceJAo4Aeus2nZ/hALacfGhe
zMFOvaUUGlciZoDTMP4PpZoHmC0nnof8d4uEM6mk1WQqoHcwLC4G2EzpecZ/
N8OpAZmSl48c+U9cQC9MOGmGUAgew/uI1Jh3vbiYgcArN2Cz+SoUthhuZ7nY
rND0X1RzXNXpzY+gD9x8z+Cqv604w7Hin510/ZlhYEbBWZ0BvCv1dBmAxomB
Lwe3QE8g0M5i6clW5j1Sq/fu4WLaMUteDQ9X/RIHuNGvSPQgLa9b5iWfL5WG
U0CD6kj2k35uMan7u015XaWrLgLkOxhxdTnCO/akyYPAj8QFgOuudDSaM7lD
4ptog8HrqnIvkPxBlrt9fzF9MjajZefP9GYfrNqgeDM7LfA31T+fpU4F80+h
wUBwtzj0Q7ND0ed4qQ/5hTGD407cTD5hLl4MmGJOtoHp9ntOxgCXQ0JdxoBQ
pmtzdKhfgqviWZPEla0u27fny5CWoC2jX5XS7sHW9WTHoaAnrb5x63Pbw+un
upUWqJc5oIH8KwghbqQ3RI4SXzm5kZGhXYuKgS7q8a0Zv7NndLhKWUFWjAZm
6qx5HxYJbUvT7bkxhmIq1ciH+8JtsmQ/2yMNQvd0/cPVrlY4iyfdKkS2d2Y5
4Ac8Zzzx3ZT2Jb04IMdpT3WFHCVfsbaAI9YDZMMKhSWctSke630GPM/U0N/e
soPfJAqLsftqy/tCJdxeMdEMtGhVeSYgSZnLPPNdftrU6H+xCy7Yo6JlxqRb
HHLetQme/pid3BJuS8ADdl86QDZrQ96RvhjgkbJzlmgZbRoJVCTgMatUbhM0
bX3zwDNKQn3AXC0nr40od1ml9VylPffWUapzIBevOXG+a5ERdwG3/zk56ZTU
qojCx6v0ucffZ6qzMoqE7pySnPGpb/Z6RusbVPDIUimzn/2UYZAjbKZvZzhP
uphR7UM9nk2qAzbJi40vGowPnOlZFEOlYFPdumqXXKjoA6t+fb723N6o8WDS
L/D2AN+8LNP/rNgdaIYOZz3U7aNOKXI25bXDjW3Pr73NH9lr6LCq8OI9mBl5
RmXyyw15zjNv50R+b826nk6J5lDNyNjW3d6byRht7PEP66VKAbCprcE/ayBa
ZHUGSNZuAFzKe+hjFc73XD8bMIgVC+b0Vl2mGlKdwP/NUSks34VzazGhRntR
qMmn6SpsNW3r1tokMIfYL95RT0R0woJHk8ioIjgD/0ha3DXbyhoC1IKw62Bv
7C4Lyvpqj+LruZ4gJm8abbhjYYvifGAB7AaZBpWHmaQyZTYvLklBV62gGIDq
Y+Usp7KZZIfSvC9NkdMppJXs8AAP8pAhrU0xTBNokMevxvzf5PvGQ54K4GNy
nby89CTvpGcNiH79EMRoeHdMh2X1Wqr6PgS4jAoV+qvCAh/5iZu7452X/3r+
or+uouAkhIBpVBr5XRXHGc3HGLbFoV+K9wzNtliVB8a0XfT8foxi1zVhHhRa
OOPcuPFtSPbQkbuIMUrl88q+59Ay7E5Z2KGZUwffsVd9skwx5h/cKNPWtGh/
IvaN7z9UxtbSJME3e0bYlafJyYntz3eUIsE4E5CmbXgdRDSa4L4o8LZRkxKe
R38gqYBfalmDGvGEwiUrc9aYy8MnBg08EE2S18KmIygv1ckf3i8dtdE6+om9
Ts19orHU8IpPXf3o40/+S7i6heuGDEX/0aQGceVnvavqYhwzDbtwOPnp7X6f
MX1NzmZ/csIETYmCKoog7/nyQo+uQm8CE4aMvH0PoeDdIpZ/LTJ5eBY1AcHY
XIY77s3aVKmGvvATPvixFYJ2QN7vNGsxizxPQ2bwt6/HKiU3zIywVHbjOtuS
3wqszthD72pjdRJObfMx8Y4Y0l0jzVu8ZPhR0FJoF8+AXqqEhO7Hqz0Gw4kh
JFsugnHIK04qAuz2p7Pvun8xyLtOIza5k+RNa2qegsxuw/Mbgt4Z8a5VrzyB
BaZXS6MAtUey09tfUuauwOj8tlfiUkEdmsitH5xEwVyJaMfNO51V7TLWd3Un
/iPn5OhCjBa5DIFP2u4lkgzRAzPIuazXyh/ujBpPrSRlsRi0Hm/ZdP50L6Kq
LvkH37tA4js10Kvy/Y1iu6ztqL3AeFiYk0NUN4IxRNz9IaPaE2oWVh3a/3VS
6HKd4htvsfhw7d1McK5BeoQdYHdESw4t9+0DscUJrU/uQfI2UxUwTDgpl5UE
zp+qRc5/xU8JSPywPYDwZD1yeJUBQoDIFw9ga+s78fHlqUkTxjkiSBKWzYsW
9UeJ7FJpIajDGvxmnZSCRuu7V3lp+4S+jVAJ1TOT+JSNAYdjuFQJpnwG8dtq
yKH6EFal5pXtHN9BoIDJrlD6RmRiuVN2DJOXhB9+4z+VawwTlM60xg7pXdbp
RRETrRfEiLsgmmGbdDNYtUnRi4mYHCA2wikTxBW//wmF4Gm6R0JzV+gbazaM
X2yeA6jVIYFUL7rl5XHTAr1Ik6Ia+K0F58pbR9w+lTkyIbd6mmOK/15V2vkp
Bzfl/Ew2cti42lBXV3Na9NXCUvDo9XrO/eP6YuIIIv5LyTxyGJaxN0hG8j/Q
zZk5tW3u8uSaKqjjTAkaOLFKvI+JlTkpFet2GUnMeBVaxKLQqx3KnW5ZSdBA
kdOrWy2NmipgkCirbfjYBhS31w7kN0SBY2irHTREm/rALtirSz/TGUUjpZtM
2KhUr9sXXFMhV2VHW7YhdQeh6RT396J+wfSmqi0wc0HmHgHAayLxRvdC3ghF
WjpbRfrWYvsjhtXy8uQnq+jvlEL//wUc1XMKq4U8ijjg6H8eOakWoUm+EaaO
eKuyxtfaK+JAoFDdLslXsE6s5ZEEFPReYIkbSc53D8gwQ/mwcTUvm67DNQfI
wrLYBjx9QydK5VclzJ9AYIwW/IniTel9AKKD/q2FwMur2nVjtglmc3VCCuwh
QIO7UU4kZGaFE3VaykULLnMg2nfkHv460ZXHYQncgE1yzHNcn9lsh8jt3djO
9XewoE1I5TaIQ0YGtmntmhskC8AhJOsag8koMNgBQZH4EZq6ht0alyVfX9OR
JbT0qoS+dTSYZ4gu4CUZF+aFvGCcwkfrjUUlmsBGeqHQmVohN3UktAVMo3q0
mvWTcPDVnDxREoYknFUzhF0QszzFr50H5wFFQfVuLM0DG/om4vbPtz+hvrs6
Zy9iLup4UNUuz/WWRpjrYj6hmY/uzPuFcDXUFp3fSwR5ep3XMzBgcaiJFZ6K
tsH1r9jhp0gqZAYydEG3QJ7a1iOq1Y6uxjvATwyu4pem/xTlLT3UsG7vodoK
drZf40anqM77gO6v9UZYzuoQbjEhigLu5tqX6ro4fsZ1EM3E9BCd0m6zDeK7
L1WLOT5kp1MjIFIN90CuOaoWwOqA6upQGNJf2gDMLSO2N+jJ6e1F2WMX/Hml
X/a9Nbd1cZ/pxZucpfu5Ms82da7QDyfy7HLk+WB7ySSadfTiDhm41dIWHpYX
1FYTXIZDj1DRGy22L/GnG5Q9BD+QhF8QZZUH7S2686v1tUne5SNVoMexP2HY
ech98abTYJVc+PFFQOdFug9QVOhFaioyrr66tLT4pKLG9xS6Z0wHe0xYbRdc
60rK8LOVYZeazz2PpcJJscR6yeq4J2j3GmKe7v/JJrQStlBzVSML6wProouN
JqaCTPvtVSAJdNkDyWKggWp47bUq0JOJ5zaLNv4l4faNyTymrCPzyPDJ26U/
ZyOrP63ZLjO6KqxsMj+ItYyjGVfm+t0i4giOtBGmTdc5SUAlbODqYLHOWJBb
uCQ5Gfj1Ij/67mA5rnuq2eCmuKCvzoSWw2ynHkM2OT1mEpMJ75KiZBuWrmpw
hJ6BeTuADnGU+t6CBJJodaPXn60H+VwIP4jLzY/ByssklR7Xj39bOXwOEIMW
jszUTAGpMEYpIRnwMXYleVJzVuvl3fmm2MBCmXran7ifrMaVrUo0lvt4MTZE
YVQebn3k9vdezq5STM92A0h5S75ckxhB1dobtGmvRtZhTtQ4mNTIJcAJ+RvM
yK4bXpVehErx00SKNEGi9x1xY3Q/w2Xjs5fZfICwmHD2bCAGZwnH9VgiwYDN
vpoot2KHBnv7fCNaq2FLXWURxrZlKFdcJrBNOuIUOPk405Mutossq0xWPbG8
cMsgya0wcPpEXjxQql80JHhNv3bee1yfMgr5hY168YaBMyqrHRBbLckmaIHJ
b7QyOQPyd6tkAgl/69XZojXcqCht4hpFnlsuJRxr4UmNMweeJlCxnYbrnsSO
l2/SfMhcZBkDRvj1kKfyABb8FuAjxU7geBIyV6mG9P19J45gMO3nCfvcyar+
A/XPA1mW/YDo875w+hAFt6RBCEpFhydw0BzP0TGSpxyB0lI/IDlh4Q6S9DhP
TJrjAcHTsKfffmO8LmT4wmEXsjyOXbqKXVd5kZArHGgqXHjW3lubiaiWicp3
alawhRVUG3AczgcN4ryI8AezooJUDx6A9CiAkvUmEbRvhJrZzTrEgnZvW1Qp
ufbXKa+LpDTU1R5PF1JzzQ23Ovmwk69bD8DSToBNZPu24NTF2Wq58sORQFAI
eOSgAXOpjco8dVU+/2HbBOzmLfqh1WWfjNNkB0jfdMai/vRvUBuM8SH6fNp5
l5GLPx2pVBlw+5HCywrSqGvyTuR/xR2OeWW2e0TWdBx1LwnU1939DjHjl+Qg
AJVlcbomIRad3ivNCaL3olwl6p9OMyXqJgDt2oU6PXp098v+WonjRz/559qi
Vl7ERascehuzShw+jYVnKg5KhA6Ew6OHxoGl60/reUaCjOz+t7ecBKOmhBy9
jUQLR+EbYBscdE/fft62cFPRmBy9YrFN3FLgNm9RFir28ReTamMa5h934KSQ
15jLWCQgg2aJ5oAaqWBdIaLWKvfnt7mziqwbEaxD6S6y+oIzq/cfWlS3euU2
8w6LoGOuORAyuoRXB1RcgPbMPzZQJqtBNHgseBrXl9QWqus05Mfn8HeObUBD
Rwlh59d81SNuEBCy0GqPNSEzNdlL/98OK/W7+mhhpYS/aJyeddliwTRCsdES
0PWyHoeuhIlfGyfgDRWoLdlKu3Akq7zRhtk3Pyy3GU2U423fDN+tYMx+N03+
hVN/8ygyHzRMRLqwtWoDmXo14XJ2FhIMYzEJZb9wNbJYmaIs75dW0DICpqkk
PF9ewVrrlHmjcKOV/zmErcwA8YIMbdwmjYQCKFksabXaogwzXAxqh3AfWkuX
8/DWJeXsdz1HINDHAfjYOdZYgAQXWljdySmyk2+X/5KJJ4tHZgQA5XeSpEte
yYcSSZ28Cxu30iZml0kLWZOEOhltvv/4FS6pa02FyTsW0ohsPHRIUEyLOs82
YYNSifT6OOJVBGNSlf8eTTnjgl/LOnI4fyRrA5KTV2PoUHQnSgtlB3BOJgOK
QI2fk9kd1n1/K8W9a/0mUwP4/KoJEhLEIESPkw6VukNmHswwj8YBfyqx/3oH
SrtfXwGPW2QnLmNnwQpLRU51wxbltO8dKLQFvJgb0qfk1YwMnfMWaigmQmvL
8SeO4hhlVUbZOQz5iSOlXHIbT9RvcnEdcUrdSGzJsLr6AKY0ZYPoFQ5h7dtv
aUMpBdkFu/nQwICDjM7bsAwbciZqfau/Fy6C2hpdlCJg2xTlYn5M5O7/VkvO
YzKPIdktrYFIOu0fsBcbblJ+u9JBnNSnmFigrEZ3F9UrmdChTi+pDf0aIO0U
noHT2qHNdDS2Vu6knTNfLzYhdTumrbCmuZIIxy3CT1XBFhnO+dJQ3Zr9T1Fo
jxfpKBFng9t/SOZwmNP4IQVi9oMXaQOdj1rjxv5A6dxuGLlbWjZWm/M6/Zih
/MK00V7LwCd+eUZVnjatxhLnwB0NDOGjxYX+RCGsF75DoLuUDj68qOvCphVJ
2esWhhy2C9WwO9T1RLlktbwGbShcWDoHd5o0aVaJ9SE3lK853fpgZDpR4Hao
ZoW1pyZHqPneHm7VDVcBHAPY5kcBj3b39rDuyAJYzmowpKmgPkz+SoNz8NcY
I8Kzjx/VdmStkA0nvmDe+Nq9iGBkrjfxq4zr/mLojIZwFppuKvztVc4aBgBw
ERHRn5HBZovnQ0HDFlEXYxLDx7u0EytFTlJSA3yV7Pz3cM3ljGjhta4PlKZt
GmX+oCXUSgSkA0EeimnDQWlwBIvJJNs0fkERMz7iwIDIZGWAvEW50Bq0Gmnl
9F5lkbhmq8vdQMftAmtDLr6INaE5AVN6z4/EE0yic5xeOADcopD283JJIql+
AqK7mWLGDjC5Xs3RzP7aGDaDNKCx/EHvIRoMYLJe6Cqk+dh7p5cl+1jzGdYW
1GAxmr9hVKdebIbIzYGTHYZk2VQUIRn/uySPcOEwRxGIRYegtXifCtXFzp0t
CPJEzfpjB1gh+997hQhHpELKPbzV3/UfiuPas4RxFNuzxJHlmmSWj8KSubTq
5EBbDnFnoSFOKm9Nr9vk3CgK5Q0T3oWmIquFAfAitsNEMCtgstgAp+D4g3aA
g3pILOJ9jxkDsxlCjFGJuQ9jErFvv6bAyW0FWNTSimebA+zSlVXwZe3NiCnB
LZ0zZ+r6Kkb+Frq4wsvdPu16ELq1BgjBHD90eQX+WKaZ8lB8ZLvAOAhcefoh
M/HmkQMHFfV0HvmC3Xnj/N7SXbUHyNtj8Rp2hdWy2yt9VPRtN7ROqnhJW+Nm
cHo5/zbnirq82ZQuda5ppo1i3bzWN/dUEKvH6NjQrl1L3828j2OKLl+1F3fZ
j7HbxSN+XOXcOXH5A83PX+Ox5ZkQpOUCB6bvWSKxrZoH/WTz8Rwpk/X8Rbtu
NhGbZupko+3qVk6muZEV+VJ1M5iWFiBc15mVMrHwWHxHoBNtoo+ntzzVTtnH
LER95mnKRKS20TOKs77lWOAO6ac4ZHJ8yw2T9rZ3D1g5an319FwCn1RKpPfW
Uo5AA+eZfE1fMcUF6ZQtvHqFx1YS8JCZjFzzyk395hui75lubtxDK/qvP8uY
3dtL9mIJi5E+ub4boLkmzpZfC19oXMA27Y8Ci1EwqxcNJDBZSRl9b893uzfT
5fPR+XLCZ+QWId/gqSj5rN0QLRlivRA2kKe8x81i4eSuk4pmAjcDdzYT9ObI
jmGZySb6uBSRD31iWnWNz5p5gQLP9rdAyf9OVPj6H6FFTs7pDf61zBwreGzB
F5TMiRydsXwS2x0N2YyoolNxs/+bCXm8Ze8/rHLH8UZB4qAji66cstoKpxqj
zod8UlPHooibtLo9yXgba8FOuWHUmcJ1EL9CrNWR378MCqPgsX2i4HrLw/O/
HZPGX9ahWvMXc5KwSc7AdiKSCluK9jcAXpBZd/FeAXy7TBM0VzEG1THaPgCH
xKP6ndqqo3ZevoXwkWYhuGUKvUoUuVHk/UaF0ybw3RvBKuhUJujIrXnYCNNd
DE5a37E7fbHrNCygECgfcKyUe1deCZ7lSgxkmiZTnZ+PKsSR1Rhz94dafxjc
AAfV0WLx0jNhwASOm890YOm9hdirnPnVr1egeNhJEFH6CJhN3ZuXSDsXRbwZ
hOaaK+7ytR2DcudFW9SCCPpt+Zh7ORqvYOtKn1rX/a5o+IKbLyQgOP5WQyhG
ZtUkcjceqpxeGyvnHHk+EOrNocBi28PvyZSAu/MYz6LldiJIPSFuPvd7MR8a
kpDUbrfTo4Uaui2V37gyyKoOGruetPUmNBcTeRo8RNwdwSRenCU9VzYB8V4f
/P8FugriVfVIMT+R83G7Dcs2tcyEMKvJ9iMNFA8w2gAMLNgpKEBsXZmdGxo+
9nIo2XBVhPB5L5s0xLW1Vr8l9FXML3Us6dyq1EsEv5mALvV0/XxlsPK2XGwK
vn1DWSn9rvRM5F6MA43n4Cce0Be1IjwBE8hRAGUv5ZFvIcrmM3ZZ7XVy5KVF
8Y79vJH5funfG+d1qQDTJcYPBAJ5EeqTZU4S9OU4r4KkYOBMBGKhEKQNruyl
K3kre6TfBqdDkAGljKnc4xlHDZHMx/r6dUwuTFaCST84mQvWLFZZabP8VM5l
Y1kZNy/ppOVqSU3Ft4/pnnTXHjLbcP/pw81C2ZJ6Bp8GT3360TknuhdRJOR+
upta05fjUTgr7c+p8KOwDsr5o9d8jbZTJv5aaSeuqWSsF7lFol4yYYV/LSOR
n8Gk7TPBKU9uH8edzIH6pabWXLnVXM57QyQkCkI/F3cOJL+rPr6IhvfnI6wE
BtGcsxSqyDZXH9UZ3WfRiIxwgFVzaGcPAuMCYo7LwVOZaVtKIefRLq5BvQNs
i+hZ8GDYToiRxphGuajCSclOaOLOsZxwCU2JMtZd6YPRItuektRgTWr0qwDR
vpKEtgmcNXWJU3oYYKVuLABBZ4QZnviYToD4EUwqYAlqW5ufYYHzvlCY5qTb
uLSk0Gp6tgXnWMyTOF4zRYnHkCm18j2BSYCExiVowiTbUXT0MVXmiojMF5Sw
a6JPBYJBkze8IrQNaJ3uxPmp54/Uu/Bz2R1PT/sQyEvtPa4GcXhM37PaOSPj
0mZTwTxXNTmux6MOyoupfiDTdEnLTklxGq8eKNKJjZS2TUe2pj5N0YXgh+6V
b9zpE0cQGOM7F+PqEOQfi+UGKS/h/VxYqDihv3l2CBFpKa+f+Rn+ms1YtwrM
NLEp56sbk31oZHd4j/WomqCCnWBd88sPaEn69zBCoCx8afBDBxaDcB06+efC
2BEfNy/bOVi2PgAtX4XKmP+UONEe/x/tukYJdjCVXjQj2rV9RjpeUDeU9OVu
JrfvQNV00HTh7yRHHXcZZcHrG+UlmCaxorqpeo4bWdTT3wLKlzjKzFoIYWPX
zJVoRaF8s3mZSvl1UPObvYR8h9+teXrUrt/6g2tIm2YRfxWJMHI5MMCNCFzD
yLrKeZrQgk1rjvCQiimaJZ/QDSFRA/YbwrMFSd46Z7haKVmRuYlUtUms1MlZ
6xsVztadq3a+ToK62iykvVRZznwGKPXKwf3B7XjFxH+Nvhb5EJtgQNLa1Tfh
iebgOCpAQzN6mYWP1wVCKz/eaR81qw2in0t6oJIhKgyBb7fSn1eoUM0k04k7
+lIGATyP6i4qk54AVqq7uvs1ZindbETNZDwsYdIjxJTcqhL7FNhGoLrdah2K
fTmPOBPUYrJFkDoVZCTymnVLvsUi3uJf8LWNYUEDE1T64zPRKnBKG2E+rHRH
KRrCD6jsVvQJIn+P7mAwOomyvYbmnHE/nIwpsQpjmtMbBOSsIvVBzdHS8fVC
AAMgN3BheIVVmzuhTBIrWBf/6RvI8Di+cqygcNQ96VDTtt47YToXWIlcvBKg
DxkrI+zk42siRLbBi23n3mtRYxuTlVzpO1VYiIJa60vwgfuO8wxM7pLl9hPp
Kz5+GRHoeZ6jH+Rmo3brXnKFpM9hEU80sPGfcHVZhZLjWq3OwgwP0vTJ/VpE
+I/K+UxVyvk0cRFCBLcz1NDQd1x6PJPnXttk4IjMjELKzuScvNYYWNGrOz8g
eT3eLeW1jntRQoYNKPXOaJ9UTK20+S2O7jM3cTi/Jfs3AXnSOz7LVRw7+aKr
qRwUAALzC4nU6tOkaJuzV6hWvZizFcNmEQH76Sdehq5NpkzLl+BeUgd19+Gm
m1/0iAnuwTyUtdk+xkN3LDqwamvPKRkpdhOv+zX/SeDiNBVQDU+xMYDGaMmf
bMjTbR86KJcr1Z2JdVvqTqiUiKExL7GZm5zqVyTBju2ALljra8yKLQzSRFLs
5Ba4NfdZaa26f2l+3nlG2863D+DcC2lZddQbhlls1sKu35vWGzqh3PLmlIN9
aRsKUWKZkXwuyXb1/TjW5PexAz0moOE4ro5kenZ6hivw/vftv1vSS3KNmh5R
FWboqPWIVZtapm2LoSOkcK5W1Kj/F0CfGr3QlHH5GgeXgGPRF/K7Jv3kK+mA
TLR9Ig4Y6s24W5cPLamrHucKiFhGN8FCXJirWAqRLcKuMeZ08N6cj2RczkVV
ooklyhevdzs7Ua3ww/+7XbQFE30faLJIeYz4XigNDgKi//M2SYdPtfhRD/3T
VNvgtTZ4d1XZ+854xjM7a3VcURZCMcqmz1USpx2S3tPrHt+rhhKEks5VkRx4
+LdmQxBripRcz3XOdC6/A7o6BkyMZmEo5vbt3LZJvSWfQ+DjxObNtPaID+GL
kwMq1Y6pCWu5a2ATsN94ohCIs5sSisQH3V69YvSGEgZV53WzQq/aAf0TEj8G
0ZTKOD1wj5aGx5jAXBemw5E6WU7AYdXLc106kkWES+qzegr9uW8XsOPw/1As
/zsVzaEtTnSlhxsG6TJMk7wF/ijbf0eTmiEfIfIHpmmLdFE+g7QELmV0cBz1
adMOD75UGKgumGUmWbVwg3KZ+YUnkwnIPIZRPWDTqrXMZuAsV7XBOAdGz0aB
ESlLe0LisTQHEx6yXRThZzqHDADLmk3a1jSjAkwcCN6SwMUtYrw3d5UyiTOC
hc7QxBgQ9kxkA3d8oXzkEbPQbGgzRQ0rg3dw+m4oTmKd/DeXOQ3sPO1YOtFL
KqzZl7HfGYywfvMPnk8AZO2iv5Ik9YETJi98IyR/8iA6UghNjWrfNhXPQcHt
Qp4LX/rRNixJ88gP8uEEkMVWIy01TLhdqTnVZCeRIDCSLas9LGY3FfR9As9W
RlEA16pMCNTjQeQ1rM3L+PvUDDm23v1Y2oon+s82P3yEWRzxMZ9t7gnFcEfz
6mC5qYp8aRoP9MPOWGi/wC0JPZlY0cFa2yGrgQa2+N1rVX4rxlc6L1p+IvVz
5yuGqjC/+AKGeclHV3esHsUU7UNyOvpHz19+ZU0ATgtAJY+nGeC3CTXFB8kR
qv/X8U8IRsO2qxhiJXaae6xLp5UGlUwmhrdInF4wCv1vFCioMKUlETpltU9B
2Dv3dis2A2Pd4zmRUg3ebDiemvdUS2YBA7i5oNuSUkV9NMd5tMKJ8MfpjftO
YdwIlNsOJHF3mOX7JvqQQ5tIQ8MuSfzk2/dR7jDkO7pzrpSVDeVPut6+3UJ4
TSw7RDgBMoY/dZkPOfjAMuQpjGA8WtckMyGsTu+OAZSQ3NmR7Dzy6jiME7UQ
s3EefP/MECYRMvSUOMDV/7LF7Vpb4Eu/pvVNRtSr5uaAdKyHyL7IBzORlLQ+
d/vjynZ7K2F8bhvREW5YR1LlJGuBVG+T6Dsd/HotSyaKDrVcQXmjjUqKGu34
MAMVepXuU8NmlFFFGBoxi2/7VYCZidT9o4G7kxitiHuiepKv+SyPT6TAAWHj
x8u57EiPiJzCopT2Kcvmd6VW/6k0HcWNqKlyhtxLyRZElgk7tdCQwOLoy5x5
pSarhHmYrVnZNCl2d7+1dHG7filV8iSBmixsRNms7m7fv5WSabX5/r+k713s
+vWbxX83uDhbFV9uKkizaiE4zqIigrD6owJIXoI1l7w38rmXenIcogZXn3uS
Uxsz2nzwr19K4g3IX4pNAwaDKNFqrFfOsur/xgP38OYyaHlT1MLoxE1g6bvD
xhxi0ffyN8KJ208QzVDuEeJ28PfSD0RUj3Q8VkwILpezQgvmYC53xTpUgq8m
5YKFK2QBcfgp5lgTPb2/aUrN9yP6lQtb7Hthqy/RPEAsq9pc4R/b6GzlkSEJ
oUmQHOneUjs+8gXTRi06mahIsnpAykQJVuxXqIIElTgflWatO+HUHOPwXOyJ
7D7xpfvugEqGDvZfpGKnjPQDXrjVhs/MYaQU4CHyHhxqbo6PEWkbc49/h3zH
SV8S7y4LXYBBLOpIlg8tRmb6vPaq2gNEGoKGUbVyakfQpcj/DTfGQvL5xs+p
XnsV6lzzPI1MGQM8QnQ7arMmEjVzaofRmhLY8/9mc0Z16D+LiL1z9OvU6aQ2
b0uwqCIWjVxGTb8liBivWme/tftIjEwlLvZw5aemuJCDbIc1a+yDluGK8Jws
6tFPoKbINVZL+cUTWKy+HRX6EzP83Xsa6ZZX81TD1u03im0a8UEuLpIiI8p5
i1X9aHYr5riPL9STIGfYs6fFenyJ+dPZL3S2+Pic6QuN8grow7bH6LysfcmJ
y7OX0b7w/hhSn8FfRHdIg/ty/bAX/GZTiTcBkn0DK7LVSr+aOBXaRg9gSeDK
KX6hxSXOJqhexoMULd4uCsu/NqIGGFPsMlx++TJRgkQX0MsHLb9FUIFwNAN6
8kA6cNdaWlj3qel1jfm23FRsVZkLRn3INLaWTP7bsYAEUL7CRiFN1GXJf/bm
L99HuPpfZ2vmQgMNTJJCgAbtFMS3zpVwiZeN1oRcneeCDNT//dkg//a8c588
xciOCyk66B8Jk3EZ1tUD8o2CsWG4RQaa0+OKAnMAQPwCJQtOHtdSQKErSXRX
N/aAHPc2ZlmSQtbG6EyZo2A5b5N3GN37rqAVst/+dRvc0b09Sp0ZZ412M1pz
jPjCRTJDZ88zBIMgtWYShN7n4M/iky1l4TDgh91e/+7vmjtdo4+iBpZpyjst
DCPCrscZn4HbFxwl8revo4/uNJreI3FPepdG3tWecfysRIPpDybBTFInpgWv
DW0YQRD/mfCwkkoCfqoVq/sflkHJlujjeIgLqc/AY/L57L0TmTab4/U5oj5Z
v8oX+IqJGK05YQat0Slv/m3Mb0FNldsminLfBKEJ22MOqDiB4oUXIo7lYmxd
Chx5Vk9WHbfh/UjQn/tgti0qOzr1c+mdZA16zsQuZQF7ZRVM+dtI5Ksq1cwU
i0n7N+9EUYaE8S709wY63X6nr1JGGbSXeaeIMmVQfdnAZ0W8oA8OAH0qWN/O
QxRS92tIi/EdP1fKbp+cnVEWWaDEEDA4fIyFKg9KqV/mlkcgrcGXnqyb76KO
gIE91XlRwhpvjYft04fd8a4U4oeSkZ0X9yywAl9q4XDpasWmOPwPppuVohAw
JKeMO4biiEcoXMy552XFZ3e/HZhqBpJ01yxqY/umh7cFl0Bh6FPubZ07iK+Y
beCWRi4wsUxxfbzK+a5JZ8tmLBYEpW4fQEHuj04D+/rNO5EaNrAmKfWTe9yH
OPkbcgCR7b1J7yTsfMVFq4r5L5leKP6wQ+/3T6GZkNHDEudVO+8UulLWTpdq
bMgTSfkumvI5fbm9QeGrx9DFfvY0fbj6Xj+EDp+K//eVv1HLG7Y1tkPumREF
nmkW4koPNs+4NAYWbO6fYDwwGAfqnO8MTYC9eDv88X9Lh6LFtX+5YEY9DM3l
E9wavpRbRMdTQSctVn+hEZZY6hWVKIL4GHAYUtg7yUi7LTVfYlgWzAriN/Gb
WhGT1ZvBTXkhmVcIqJcX62oG7di13FRZ1kjtFWaT/F5Oh+O2g2T4re5YXXdS
Q7tnMATFDdbQRJzk3TSMrK1SzG/7SuJpLe6/o2bPhh2Mw7hIWc6NUF60/IYj
PBz9AYQROaxsrSXMxLXf8qlQ0VEe0ILn2oUfcQWfK6zdC7TXPaHXu233R9V6
hee6M20hrC+bpJB3bg3GfhHSlIou5mOp8MjKvMXeYy9cnCJPQXoPTvTsAqih
ah6oA5bRFhZnIleBTR5dYV3ghyyez2dm18UMzquMzDjm2/PYa2vaGvHVWjdS
/Zz13Y9bYAgfpuzwxdnhRyIJTkAz56eh4cbM+tNsZFqYZ3J9uaOyxbJb+8YS
5WLJ5Cwd/c5qZIiafo4EHwM9kaj9scUalPf/DxQsiA1CJrwv0AoZegqVW/3l
9RL9rYRK9pdtKWxfWo0nlvYqFweT/H+7RbRR4pJ0a+SvjsnI9yNDdFK2QMqN
tAnNCW5/OYD2IIVcGm/1n3KwfXl9gBNbNcO6IDsc5l80bWU9ta1rclB2vSxe
d6qGvOfltSbGBXPkZHFZEE/RmOQ9mD9zqv6hYO+nKKkjcwrZ5qlLgCVCeNcR
ZBghrwPtcypLaJoaE37peDdRBLVudby9XBYKansRve8EJptjkxVgbBJJtO5D
H4fv4q6ISjL440TafC8PVx0YhtxEoV3oN+WAo7zxLXwLMGixU1sliB70NAPE
bzg9A73Xe+3mId5F0kxxgiAcslK9oIL/eOt2Kngm5pMNjzdA9tFb+JEovrhD
YGy4fmGImnwNwWKkakq7IC9ghj1ZXbwMiQmmcI2x2s3+EMOKU5mStoH874hB
hSV/8is72S05bIPi3HQ8lGivsyxYiyz43ZvfNpOxwlzBtRWesspFXr7Lxh7T
zrgATE9gS+X6eUhhLJLSfwlhzT2+tPtULmPfZ9kmRd6YAD1h8wdh1l/De6M5
Z/OqoRQmNp/pLgE7dOrEnflI/WGPSlf4DgnzUTDLAnBysMKpZF+SB0kuBBDS
JtGHw7YRNVLUWNsJAQdEs0IWbJeihWsm0D6UobGW86zFn8ZpcZhK+z7tmqen
EarDnWwq4/nHoSBMd+QVMScKR4BTbFH4esqf2CPvvYi0JVlqKzbLsH2FsjDu
1HRVMK4ZxEbofFyfE/WU7sd3mHTJk5ptvqPH+gEZD56uMRCuXsph3tWAKgh8
QkfxbQ93wtkWpWPw+Ydlys8t9W1akndllsziZ8AZBeV7Lv4dX/pe/lWfK21e
iIXLaE96Vqr3lg0VIVDaXZrzjg+23uG3KgiBgvTtXzd1ZhUD6AVrGc/hDX1h
dgF4O5hDiUCgurTw2iVDLmnJcNCYe654+SIEhjIR/9IOye2hYV9cLmr421hT
jeMPi9DgI/sRufQP/+94s8wMkuJDXNt2PA9xyWyTEyC7QP1GSPXrsrO3aYzY
3jaHsYOPSsAeLaQxYkntKCviXz/wDWCH9tpXuNnO1G5d44PD9m37LlO6yZbH
7eDhULIOR9XWFb7QnyEBZLXustpDRlNCg4DStBntcVBw7dING4AjQLcRixbB
UXzhBlVtBz0yvpPlut4V2PeGwoEv5ilcQ7OiwdytRYTe4WL2bnVezWelQ2M4
+i16n3XSkLKA82a1ItdXSo6mi4dQFg92kA5rccp27YH3aFsepZ8uGbKjwiVg
qmuPkPsKTSfdyL6n5UeKpN2Wh3Xs4+pGAJSP6Cgv14vtaAcy78b3WG4z1F/k
HocAm7PfosQisfjLcdVYzk6TWcodpa+2CLFobhD+XK0epyY3jf4cmfvfr6E/
Fk5fPzkZKK2ATK0mxmYbFa4OQISAQJryoz+aQQWk68fGxV/golsohWlGTjrr
mu2i9dJ2VNNN8XJSXhtmEYrnx8SUHZkQcYl5oTwgU28nFVAPXC1qOzVfsWbB
H1p+IwCrcj8kTMGKmqZoYAmCnurH2p4iJ31jmWroj8UbL47AHjdYyUMzo0YM
hWdpgLVwcZrXupieyQPsyEVtCkfdSXZqFvJ7ezxXdgiANFyUDi/iKH9IGWqe
WbGgoMRrFmrIxRzZrbNuu/Ukf5MQV8vXITcc4jvqo5ihDGJouJVLOg1kNBKq
n9GRkXe96UsYKq8X8L3i3F104NuiC5PBqZseqydKXFJ9hIejvmZGoLjnle6E
c1CgoUxyBgQF75AUJK+X5YHtysFf87y11jeRWg2ViDVzODN30UzZBna/bpig
g9zGUWRqUjXkqM5wZY5IyY/YVK61TI2I0J7ebN5CxY5QQX/5hEFNm5Yi6p8E
juceEd2Zi+Qdlv8IsJrYN3pLEiTPPoc0hLFIHnoc/y36FSqyL0GSbB29p0DV
K08zEPphhSY03BgMb1lbx12ed/YQbwRgYn76EUpYVGOjREcl0U3AL8CDGpQa
ltnzcnSdHXA+cn2NcqqqAOaQuzDj3dzrc+BF7xBcIU5Q1ARtSDltLIEXj/QX
pTgwOz4zbVIObeXnQ6msftVkeXK+kJL8PCGJyGvzxWbjiGZtlvwCWetPZ0MC
+qvIzDknWllUWM6QnISLR2p2MGYHi2yYxTsM+UCEvmFOdM+KjbRJN6MPVHbX
fDC51jSH3dbVYkgQeX+fG+/Wh1C2M6wJktLC2ULYJ5K8WJqvEXhP6iCw8rqS
1RSwayiFf5ZR64fJW2/uPXp9pFWY5wMOzeya4ob0jZ2Ijxf5UFVrx1/EYGEe
yIGncB0REcLhBRWLtTXErjCKNoqyUoo8zafqAHZ0aytIog/l3r8yUD8SgLJY
2CySmhAAjJp6M8nEbfwwY6gWR2kssLpXAmBPg9vMOdyydykB87AoezeOs2hL
rJEDBMhJ37OOMov1QQoQpZcpWgeq3wZ8p6+8kZlqz5+i3KJ4oU8zn1nvvdhu
ZUagJf01BCgeTkuCEbUBVrf7Z/3l0Ul3IKyoTclOeVcKVKoDwSicuSezTjiY
jn7749UCvhukwHdrSYnUyXyJj6HhEEP78YJAZZwSd7ndtDsLkZV2nhf4BCsm
fttvfERvGIKh4ZZWsCZH46g23PL1RMrS5hIHRmHz8N4GnJPHugxCjVB2yqeu
B2gyhIjZ7CRw/TWv36imutoo60Lm863O8LZBr30ZKCkXmedTETMjhqx24q9k
yfYdPicAOE0pgCvrbVMjHpJpsR+UoPM4uiOhIBMLJ4Qn2Fapz2cGi3iqyfaD
nkkW2pMZ2xSPvwTIj2ArRpL7vyshItvaMUpIX5eawdSnAXdKoyd8v5Ng3x+O
+aNYDjK2d4RJNr8KVjD2OIyClLDA2eQPsRzm2Kq5Juq9LJ9ANIKzCDANfEFj
G89u4J24ZlrQQy19e/IdhRQyu3OUCGdrDQ8uMWNoc6wwkpiOWJ6Zdu8jPiTM
L/Vkjc+k0HCSAB3Hb5DYZnCmMLtqwH9KK82bEJCOyGcM0PuaYXG9xaLIUYe2
0roT1GVjKEWTkmTR0JUa9bl5pffmSzLnoBw2I/78Nc4/HMNpQS+S21tiX6lv
9TkkdjXXUaictmCC+sOt8NykvLkvgL3BOjkRP22dRr+S62tj0xKNVxGRieCD
PiaxdNlMOwZqZEMN/rRTxbRUYjsAsWQLS845his0OTQbuvyRMxeXyUwq027y
hCV8EOxm654ghmwWPBv868zR35mMRHhGMHmBD7yz79ewgZNHErM+KAxNSJjz
2PkLp+SuiTFSeg1RPOzVoyGNBe/u8Rkb4HcmrYBU6h8mOwvPEyD/lVzP9Tik
Y4n0/+Ptrq0oT4CdLC0u+7k2lLbGlU+c5IbIq8c7kEbwRwGS3fEZzTjm9pBp
ffq3gBUXGHZV28SsKYQI94qpVriU7xLgzQ6vz8ouTs37ik7+8Rz5dVmugeaw
pGztkeKgILDwApCwZCADFAvdvPnpSdVRTU1OjtWed7ismW+q3b+6kpkdkV71
aH9yzDCeKfDYDYypEUQMChnh4aSxWiUj+FbSVKsepiFyUsD0DJwUXP5E53jQ
THzpRoIuAe1vZeVBqxbG1MGLZ+FcX+jdtr+i/M86vDCf5/4vrdXeHqrgxNmK
hV7H0UH1V50SIRhjOctWorag7Z9hhLodFIPniiN92vknb6nQUneVdllvqk2d
eUUQLwBtxsFNdHdLP1KnqXUpf/dawQN21FKeN/l7aapW3AG41hyU+p/OMiRy
MJQAgW+bnqZXNLS+qTBGu5TbgW52iWEaWc7F44kl3kOTeSEOnuv0zAPPgz76
BmIBIrqyq7VEbPXJIFyOs0WL0VyUVpBKrEn+4/ngtUumIGlkgapCQ3MDweZ/
LeitXmU5QiGD5O5/dBGhjpLIR6smtqdr/chr1sbO8h1RUs/K53WcgKRdN5s2
W+TRHPQuXFKoLq/azNcCVuTRXeNFoXS/PmX+w3W/PcUp1r8ptvBBQLkviDeA
STQTHswDqqR2OvIfPUNy0kyKIY0dOmSr9a5E9frHSIoXIc7NgoV7BUvWr1Kp
6RN+Ns8+f17COMRDX1E3TjW08DyJysBGVX8S4TG91KxL9LjJVSfrGoWRJbwJ
EM0J1l8x360Mv3QndljlltH2NW4Y23ouPYjSj+mKXhkz8LrBnEnvOY+cLC4m
DSIBr2njaxamWB6fJPYnuEZ5ghMQROc4A0YqW9kqr7S1Xs7x/1PQwz2m+0Lu
9ABFXfpnhZuwB3woN2q6ZNUn7pumjkxlV4oYZlm0BKEgXksn/Vzn3ELFTZjr
4bBM9kaYnLlozknx+zNp1R3MWr7JM7K9zL7Dt1vHLWT4+fbd2ACGR6dTMy2J
T0S0krcNUMfcIq9zgRi9gJsAUUpfh7HxAzeZpzA2NqVgLBpwtthti126On4z
gyAYqOpJhLQ5BRzTbwHdMH/y18iQdY4t0MM99e73T7ZwQEIZBvcRLKQ8NZtQ
uAa9/yiCHMvvCo8J0R/+iGI6pgv635J+Ikiv91Jh7kP+qby2d58QSIRQJ2gj
6LcdIjth48jMeMqHGXfFVoH+UM9OKr7NqqrWdFLY6jt83fW140xamj/GDGig
WIookiQUTQTjLjZB7TYtkZcAneqSLttnXclIr2MGB9Cn2sBBxEsesHTOT9Fr
F/Nhi1GT9JnoDEeEc5Di36vOoVHRBlvh0xpu2G7yTxox5GoBA3q04VbiM7Ie
HlwH5KbOTu4+PUiskkRBpNNUVxCjl+zNs3mlkXdyHTnnjQnotsuftBqUu9Dk
/5mlLmZztDordpdpiVEw23iBqVEoeMaDVJL5UMxIoEDMVqBEE1K0PNt3DLV0
4FQPOhl090iIQuzRfua7nwIVNJ5dIaTaDaotK1Q0jW0shEgsZVQBvH/FG4Z6
RSmxm6+Xae7NjzRdI5T8ppzBuRjocPGLxPI6wp1a9XyFHoR2bTcbSfpB8Mg1
VoSfvqVzIw3q9dqn4a3/AiA0TLBtNIvlYVbvvcLOEkhvdbJZeYF/FOqnspQu
8FmM5oxy8ikrpGwZ8fwdV9wGJeroYpIhNvaGjef+lL9q4ZOrBlJXZLzyO3Es
TGpN4tLycarIBre5qD1b0DORqSVGFF9ecJlf9XafRcpngsMSYP3ji294XSWN
M9dqNpCmTlIsNspod9JrgLnIGeJpRLA2fQCD/Pn5fYEPBOorFiWZqQGtEkR3
Vlw1FUa7ZOV6tjNmywogRj4GVfHjTWjGzar1hLAWw+4T99+Xvr56EJ/TknZa
DlHGWCxiYMHrock0CXVkoI3iTl1GXotGTjm7TaH846LSg2/Y8sB641EpLlUU
cvHrltVYUxJhB3nQSBMO6iTNsu7rgWOtPEsPJTnYlPM3MSOcOVoDQbG7KDBS
hyh7kzjTjR9OopXocwCxolSixvJzW7hxniKr/xnbmfc9kfuD0Lz8ia3Vs3bC
zhdgf6D+f3QXHolme/aj63WJEzG3l6guL/t86AfzOnUmqWRKBNuxolUnhXiT
78iOzzNUro93MOmYoh1z7DPg7cax9g5hJXGbO24V2FogIiMhue/REZvlowEJ
gz8a5HZXG+SzG7r2B51dkKslIHJJ3R57DskaMTDQU8RsDBWL32pVISU85FU6
TDey9U52IekkPsxC/93jn0SZSANJkxhwhOF0S9AducauOiFJqGGzGR8d17+B
7KdEHfL6cdKIwFYlympVrFdZ50FwgXjg/Hn4WbhjBilEx8YGZwH9+SCQCdkj
KvymVqq+lqspdR/7koxwtwHJmJPvAE8m+0kZ8TwEhkVPt007+k6ib/eKp5ej
MKkp9Qi2dKwXXDh7vEhQsfX1p0Ro722YwcGAVDpomq+ETY/0/LV0YauciIgd
wndlmZh7wgNgEd00oNEIFOXSx5EGW6ivZHnCRrYe9KPJmfl1g05JGu03S8Hd
9/zWZw/+n2aRjtfrnW4THk9xPoI04bxB8g9czP1ou92Bzk+LipAYN8L4zZlA
4C1/ltWSuf/SHpQKQdJGqN3QKqajB6/1KuUr1cN5e9eJzzCfA9MUFbnc5IPf
f3SLztPX1d0xlURyved8M9UI6m7xS8viJhFmeenYGhZLITwKZD2MbV2ZWu97
B6o3bE3IvFkenJLuFYZK4lxgCwaPpu4+nPGRZBRbDvW845w5nNLXHd5IlkQk
a4CKm+3Gm+prdzZ86a6cJsvRFqXW9tFfvWvEtXRmlYUTtvtkbsEJVFWTEf4b
lQtNScsHYAUssvFKeO9XVARiTR/9P9kWsw6W9vHR0is3Nideql7whVa5dnHc
/nHLCBovtQlvUYql5ueDPD62L7047Fh/QXkp9+EvZcQ0pmW/XwunLP2p5lmy
QKyOxa/lfgjjrBUHju3c5maXzm/mot7ie0PHZSbNv8bu8+aYRGfHGhM3Ctkt
p8Fzn4A93Xj6VFnjSU9SJNvEyw3YctWJfqV1mV+CZa+uqIVUDM0tFwB7MeTw
9zksu7VOthTGDW01PpWZj9ghHH6ob5goKUipwi3Uf5RMl4fqbLMDg/FCTBNQ
ObIFrikdwgbXKbU/1wzegOOKqo7PycxS1He0RD20/Ua4fd+7ahZ77wpBDAtK
F9hvYcNnQDv1FkmJi5zHqbW9FQ2LoFLMs27/j7vmxzXHOCjnQQAuRnndrs3U
0tbgYKBXdQUtgSj+CFPkNJUMNnITIjD3ACwVGh7JZJ0HWy1MVT6DU1yZ4OHW
9KEmFwe0ZJNAaSPH1GqIir3cWRkGLQfxHamOfrmlvPvS+Vt2PGbdbzC7jiAI
T4kanxwYU5SNv4RqLPVA3ybHRZHMsfdtvlSmsAE+kOrm2vVX+osfsZkDQwJe
GbcQpEFuX801pDh9/+KTyhw4KrV6cO59hrFCmpbttcJ7TEEmkZ/+JRroZjy3
sfm36jt7wIRw+Y/3I/LmM1CLiSNnxrFdyP1JCInLz5JMVsDERU24HPKSLmHN
GPQvvfZstvuKI0m82QbxjKn6Z4JkB+e5t8rmbeL0rLzgl0PwQAAnm5I4SMxy
tOXFYz4Sxsyxm7MObE7oqk5ek0I9uQrDzKY/hJ03SD5MZq0wyMvaUzufOfjl
/paRvzrXJf8y8r+szeKMRgwzcqCU/GOwAUAzBpQUzSAzRGHL20da34B6u4k3
xqGeapDbrO//rmePeHm1mkGAaIYBaDY+WAm7oVUi4dci2ofAW/kWQTSYIfan
Tix+X7La4XlJK/R5CabB2NXuAUvcf//guoJxFVUXLHABNCFsP/gpAxF4paih
aeqBIgbW5N6dsc2xgeYo6A5I3ogGwvynCffIWVpf00P6YxA/mNPh2kKklzZ8
9i4qPMGLZm6UMX9ZYPWx+DRVnqh6Jh+6bEd2WUGjPNYjD4kFu5H5hi+vgBGR
DYWGPND2piNYFaD7LpTD3/W/X1a2nXMb4XVxP+sgfg1PBlfWgmknBfL3unfE
xAsN0fELvOfxbCa5jjsRDjJ+RusyKjJRDxFSIVs7sDThuyYGidakH6JPb9Dz
q81T4U/IZeRJJNe7ipYaYIts0996A9CcDm87VwXfyF982yG033i7ujtseHSb
zUOPFYXeRyZAARcyo55lfqCCJFymQxmV9mkX3Z6lO2I2zM6hqM+dqG27MvHH
yMPJUGX1e3vMNDTrjvhh+ChTazBYvHj2DT3SPJlbWQ//K7zT3/XaXMnG93ow
TgOe3JE1m6Ph8OaWpAU56Ks9cSS5iwSqr1B785VQyP6DhYG9pilew6CFZtJG
KINYJHcPvCQEjzDrCZ5RX/VLxpEhv4rjdbNjr4dCP8rN+rutnombq3AwgWOM
WUQ9eiGQ5QTk3uUjlRAEznPYQvKTMN6oSZEn4DFnji9dfeyEroHtXlwbUZVQ
5kIfTke7c831984Te8xnvUjIICqYv2SLlB8ADiRNFV9NvW5C7/h8Hyml4VoE
2xQQFRznq+RkgI1fkaJkAqs8HHjwfPCVQFpdc9jHKu9Gsao8fzt86k0ZgAGR
UoqKGL3F8bhH8XP945xoOmXpKJ/qprfTHidiZZDR8erM6ErC+/0USIB/cwns
HYKcdF/htSOGBelNcMw1PIk1SCOtiADJZTpaGPXwXPRYFB62np/hjuROsQwW
a8rS9G2SPrUs5143Hny7l1Ys6i0Ocp0trhhJTmKFBOdeNz/Civ7CEywLTomM
NW7b9YmtfYMaR6eoH4WlN6b8y0G3Hd2OjH0LCMj7lbFPZnzt0LFl8vowyXHs
bcG3XV/B7GMLS4azTI1VmzEJsuIl+DQYTuo9qVTM3YGZXQf5BtUQUxjDZiuF
f/15/kah7U78fXxi5bzUfx0t9aO6Z5Ai0nncGAFDCpaQiMluKZLBQ12j1GBw
8WVxC11Jwpu0rIgTYjXJhgQf2Cb3bNU4Q7NS9qMDhqUHva6T5IfQnETnSbWh
CoR3QZvy0fRuf+DFSxweTgDqx8/d5oVO0ONxijLNateU/57mtAW7XfIZwd7V
Y6rycUbb7d4EvFcnqdq0D4X2zlLOc3hxMJflhDqWWOp34w8WoOuQgqyQ5vnM
qs5mzmbyN6I9LIuKTpVgTZ340jjBBq+AyIXPLfQf2sUL6xbxNJ8v+BYtOSNK
MxZQPi0uso/vyY+aR0DP1UwCQwd0iA8CsgPsg0pKlz0zrYbtpUzw6WELDxBY
k709k8zh3ii+oEB/ntkutcqNmjXkt33xRwKVOXE1BtLnwu45GDgJHAJ0LuWd
/oIapAwun4vWD94q/2r9tWoiURaLJwLolI6AJvRScZ2yRK8WgHOfhNnV3kt5
LS5zzsQPQu/Q5+KFaV/NJf7bWnySl4y3moMw7w5xrv9zD0Et/hPv+LkR3Ygc
ST7AX++q1AKmS8npc0AYIbbyhIVUJDAA6XsXxr5c+pGqy7gTSx4RlhiLfErY
eVtFH8tJ9IaXwZWAvrMfRgTLREeJWw1M+rAUyKPhA/1+Xuukjnkgm46udAyg
caWO0BgZ36zKjPs+W3jRvMlgdiBw1kGel0tYOQcdG6Hpb0OdopNqGTZgF1vz
1TqNV7iN7lgRS8yhNcUPtDxRNyD4Ho5+Xn2crXdACiKNDMfY/3Nqxvam2dRB
KzajdAyBST1HELNTpFnVuXI5Tuj3Ex/1vivePzjah0daBtrpX2iBPLhlMEN3
RDHyCpVlYN+uPjbpagkSgdJSZcGtWKR7cIkwXiABOoyN+tiC463alH0xqmAX
JWUNzVzDEVCkBMIdoaJF/bTfLybhwEhjGSxEpXv+rhbXSmWDxdKi+e+u5byw
bzzUqEjHl4tbJtP9Y+1rtKM+j3Q+5uokXg1qsBG55q3lGRJQQGlnKjk7Yn2A
MOOAXdBY9v5Kp/+Uy/D/GzdcNv6y5qLQcnC2e78njg+88pJErnpKXErEyC+F
MYBENwKIO7gQTk8UUD6obKJZEooWZcdvdjBQcBZOnXeGvKzl0WuLMxtcrqxA
9Z3/COx2tAHLHjRl4bO0uh4WeV8H90/2mAkf83iurzIfAvG3PG1X861pPdlb
beBJK+8rUptFlsQhhVnXGFu8nPqoKoW1ctU9jfGzuGOapaXCZ1LVl6DCV/RI
xmJE1hrhfobvBpuVuBsXIhGL5sFaGZoJas7hvr1bCYxH7mk36dXXbOx9PkXj
mZfGFgLpBJFRQx8wAibP39H6yQGyETUTUh0dMUsqo0yH29HzgrDbY4gaxsmE
ZE9BQC8xkUc9NbeYOa/vQcBUKs1cGkpZqxxaAfH0jhfIe6aJwlT/5YMgDZkr
2tsBYWPRWQ4B9ZofGzn7fU2f4VHk2qSEJe8TyamhlR7Wu13PQLlRFG3zWCIS
J8KNRBnSC06HV9ggHREdTbE7rbuG7B/daUFlTi7lJNbL3pRbpec2lAgyUUVM
a4SEJuZpTBGI5wwYG7JkXZSoi3XKQvRcczHRIC8tBeuzQtNOg4hVsgybC/50
xh8BisId5fiVQr7BLuXa91JT+RjSs5GFoxUwk44EVKykWyan2hIaD30dhsuI
eVMYTnBQNbjoAYG59v9yFzRKm3ILNKpe+nKvu/O4HoOc6tw793/alOWLvwFD
sgM4AoaS1mJ26FHe7rgXFBIDZ1AhiUQ7NDIKV16wonGnyPx6ocn2Z5Z4AAiW
tCM6UgfErYidI16mbNFS1mq0FhTM2pxBvSVKDVS3Sca+aeStGsnBsN3OUVAW
qV6tkiMYj4LlVqpSxbd/Ta9dMyyZI4DKmClmrJtqQbFpaGWa5WK/11Ql696x
w1G40td8oG5jwIfFXIYlHJLOoTEgmstIwIAOy/o+rUd1NbeFNASSQZkS8kLg
rxy+/trG6QPkrcVo/TL3WX3sIEVUBNZ9QiZOGAbqOzSuBCxJgM/z4OE1zTgs
V9513usbBwuiALXIZJebzTTDL3vsmc/eO4mw3UuJyCh4vBXOnz1Wf5A+H5sB
Z+HQO0brHes6yINakLKkeBeMRiTERx/JrY9AiswzQDunM32pSoFd2ZCgX+6v
qIqqbzYfd154Ov/Tn7m8doEPOuI+MHO4m4zo8z/5S1WlO4Dg4/9zognetfio
staoNNSSFM1t0ZJY7ghkOo0GvWETtnaceXBPtZBly91+KadPbpOQn8VvRo2J
f5XvvhQR+2wUc7yxZtP4pnD5gAcRNAABL5gjt+BsSnTgtJZ3dzi9RSdKIiXw
yG8hiC8+BP7tk7pDm3KPbc1ayDGNEWw3LB9dCMMYkeg+8I6q6LT+sGWcEJrj
NMUpfBUrpv5LB+SCC5rIgddpkJA6JDhVlnta1NJebthILU3T41dsgg/TGBEg
xiVajj4XBIE5qhiljVoTdFeldmtn2irZP7O+1VQC97nCjgM2kzedffTpOGSO
2bqTaxhKXb1Fj0k2P/l+pyclbXSoOW7Eg3wpMZ7E9YbxkqtiFhCZWA1r1luF
Tu6rpbDLngjW7dmeCiqGeEYljDJUqUkw4NdO7xeXlgcMazR03sM26dz7Lnap
3vId7oAx16WRhd60hqvPox3aQLKqol8ikYDC9zA3dPJ54saKDpe5xO4t0kQY
K+cwiuhaVwnxHorto9PFM/x1vggoNwbsZnnwEVt/4NyTx5ICdCzw08tkAs2c
sDGDWDUSPM35fGwlC2W53Y/xHxuYlHj5YQJpr9lTI2fJJetXU5sTDxPF8UwL
4tbF1iLhe1sDX58lM7Tc+vKvqPi46+cmfu07P9WInCs1VcwyFmE12zRAvcTI
POkKEc41MwtACBk+d/2JmiPT7yE3cA4sqk2y9qB8b6elnpKNWPyqWcKmZO3r
/MHgMcAVEpMDP4ZaQ+b4sOBFzaaQ0M2oSf57txy4UEKYDEn+XCKY26GH2Bc6
cn8S4Al938zgOdMK1eVWIi4jrNPQ44wuPhysljEz4OK0ij93xX/1ejYRCXZ6
FKrX1XEFCO0M/93DdIzkBVQFIGkQbP6yqLFf8GitKkt9w72WGie4po7vuUtG
B/X2rTxtQsq304egF/EzDmS3Sv40owSg5WYAdYkLsqsKk0jRQwAfpcaKTj3H
kdqpo6NfvmbWCF0M/kQDu0OeodshCsRkfm4tE41Q+d75pBe8fvr+AOj/8EK4
pEsyopgpXQ7yaEf6REE45+lrdsS3yAnxfRALXPMQZioZAEqW+4Jnt0h/qBaG
8Nd5GS8JuJtUcAeiRjEa4wYktWmF5dKx74X1DsIcW6sA0WJRD5nKunu6fcNN
wBROmDD/T2amoxpgW9zhppnnZlrlC7J3TRwmj5FzE1ey/DXvh/bylvRV5ZkY
lIEMcIOq9AgxAmpyVxBE89j5LDZYpxhaImcMWZzTU0ZUB8TzpsyWq8LoDTCq
uNU2XoHXqc8+eeE5sBv+6cCs5LpBxLHbv8ICx6ouvVByKGuKpWcVpiDc8CKh
sc4/+ND6HmIZzweXZew1xUhZo5d31n7ZQBSKpzK+3SrUDKl4ax92N4+30m/n
Ww6EinsTar4SaJncWqksOHEU2HCKzo8v2uGqbTwmrUeGv6LvCY4LTVc6iY28
MNE1+y9bE2A25KE20uXD1tYvTgJWItMx/xHHdMsiC0SBkwLalVs1bRDTElQH
8kCHn5XutGQEmcLCXzWIMSuPOIGYiw2pbHbdGmkyfYeMyqsousPR/+szWP2c
EzM9Z47zfZZm7x77RMuIKSMKIoa+n+m8xT1dT5a7Zudc92Tii9P8P/XIgqer
X1ksCE5dbkeW3lIBDnNdWFsamzogkLPYlO1I+Kn7kXzx2s2XfZEeXOC2krvk
jZsIdluJ0fLGUzhCQjPPkH9ST56YOtwRddFdfXQ3i0KUTVa0ReexvsHHuRFS
PUMyQRrudLHSRMGHD++lF7CLASTvDUmUsCkD92H9+GdhsK++JbjYIOeBA0iX
cwIxe2DQXBAhWoBA+OEE6DHA5RS9VM2vD218fvuNrrNT5NFwW5q3QSJ7Yqsc
SurfthtDKDxXiuUuiFe3/eYj0kiXHmMnDuAcExntTNXVs2JMCzl7FegdrYA7
4bmfqkKWuEyDmKL6J1GokuRyw3lXJSy6ghU81VSoWNyrobyqkvpY33MXVNka
/I1HpxsvpUvg2wgb9LG0sK7JbBZ8m6PjFwQbZNiuCQyeHj457ovpLgcHSv1G
PreKl893FQPg6odfE2qiSc+SoG8jW5qdPNPHkeHJFtwNI470jzDCyCtgmzS6
zPgoFbqu6WdmpfWUC8xcvI9fFG8Q56vdU/kOMm69dWIp+MPtcWErmsrELYgP
Ku/yC5AyoxaGRCL1aAa/QjPXEUoxf59n+HeBQOM3Dcnb4HkrzMGzwRThb2h7
kulf8ILNGiUWTA4Tg7mE0lYSaHJQbyLi3oyU30Txzy5JV2uw7trvvvX2y+mk
Z61n8N2Qgpy2fwyApYH8HZKdbXtsR1ie3PomayIOwjIgBlOjb0V0PS2Nn8Hc
oI5OqF15tmL8k3Kj9yovLv2EbvKaUP17BmNfeE+f8l40hjnPsGCEzycH74SN
QSl1nhUex3/nAlhtjg7At/qgVERcU1CwEDhfN1ulyoMh5JDluQdiMMgvogn7
msa6a2uC7iQOVR5Vl6H7W86i6+660dn4Zc+N62JVCbLYQJXL/dhQybS2eZSS
u6S7HBG9uk07uKUerdvgPWyPBDU8yfoawz2HyOnyTq/t3k0ve0WrM5Ch/bbr
GkyTp8SImZt8utY3U8srtTBL4h9se0jxUZHVRRgWf7+GCLeZZS2VAQe7E/FG
U2JxlimI/OlxFwlIMJwpCEREttysLLo9spAW83RsvF4gl+HYgitibCmBLByN
QbnFrZnjNmbHz4zGlm4rlqjxPw7wTTTP3qDqDb8KCga1I5aMxMJGAAmHZi4y
9sQYOREYbD440WlzRagjHo4QdXG/FswA/l8yNmflCST5E4VNciRS7IexB/lT
yUBf7O8WOKe3udK57DVsthk5mzFMT/EESGOI7IjQfDQj3Y5lhf1RX8rj9rEg
k6Ffl2PMRmt8BQs6lvr9NZF20m0QvscYr/IpKePT07oT3lv8Im7Oc4NbQO8x
Z/bgX79Tok/CtBnBDZTGN08Qs4R2FUO4guV4oPXJowlAT2ZIDs1AcENebvhr
ZFp39egPBQA82sMj0MP9rNqi4/bCaS8j/jYM4qX5V3Q16KcHFjqC6FGeIv5T
WpO8QSmzfitLMHz3ipkB6ahHJmLQhkjNeSfPgMLoiYgBw0pksz36De8DjrKr
46862hajrhhdFpodg6p3+2itOgeiJ336Y76HXFe91Yp+ae6P5XnVEwBogYY+
Xt1zs8ACojoVrwdEBmlN71ZMfZ4YdfHob3AAF+gyUMCYCPufuX4sRbHZaGE+
KxP+Dkc0NDNX2M6ZRV4BT6EuW3qJLnxdnwL9U9wcdw4ADvd8CGCMbEPiQZdJ
FtSxtlLELdhT+fFenlmo+oEBuAx6S4DSyvQIrWSarQ/jpOwDKPWKTJR7fmqc
cM1PvQhe7cccDeSCGxvdPaNOv1o42TYFBzU7J8S4o2XUukIvn0xSMs4P1KSd
n4IYKxIwUZgsJbqB3oyhkgleLBwDkhpW/x18LO1AtJN8NqSnG9WBGT79YvcI
I/SiCNOwL6zuyNZDcRza7r4gKfZjewrMc/xOxrxPNUNVMKhW0W/eM9UgG/zV
epV70libas3dDUlHNbpVpVB7o7mF6l8fJMKKp6Jtw9i8NXC4sx6txOADnaN2
1YDMhvG4GaM3nlR43dDr4WVRYi081KmDbpKYU3a5X3boNQdEOG27tNmZB26k
D3LBYvv4gcmJSePDyAV2Kn05Ng+5YfjLQcphO4Gpf5qszY+ZMz7ouSxHRuoj
1WctrzeKx1LnOBxYOnPPiMuL6bbqaDlxpTLIkOyP49qsVrrYwWLd/Fs9B60/
q7pSO/AKaI0ziVdj1cuXLV9lW2zXKErlepbuL1/B1MIId1lEUMSyEpHZYE/n
U9UUMXl+shrqut7h9fuiOzh8yMHLCccOXyiIhsf2YnKalBGNRU72D1E5kF1p
JG7fvqXV8Vm1g5l20yl1jJuUpp+dM7Mpb/wVQWOBcKbQB3EN/PlbI8oAgtcS
UR7mUGrhFdqTggoDQr0qx6CSGfLgnb7EkAJJQ+t7tSE9pNLeT7ZoeVM5ObEb
X2PMOCHIC+XeuW0NqAD5mJsoyZHpX0TXo1MsO1yKwkp+2UMbFgBTIJsMVk4i
t7k39/PEiR2hUiaZ5Veq0FZrIfC4anTYpB6CoPv4yQOYSa7Hfm4VFH56xbqG
genlc+lwCSRSX+H1JZmv7JclOLukOI+MYSYMeUfmJ7xml8vJ44QDzyiZ9WHx
mW1lV4PjdvNSJngSjFt7F13hCnqV+gUGXuQYGJPLYWnkZUQALz++XontH8hm
EmsoAY9UNyL2NhA6fqQCSkp8YMl0DAe1jlwy1HGBETFBE1RJbM14VUBDJbQG
9lKVcF418NOiq7QlFTQVgedRXk1VYjFGrkrvu901nAlnuKA7P2w3Dpeu9qzs
vuBQ9jIhXlPHlqD1APIx1bOpACe+3tnZr6cC4jYKXJmzsvPYMuiZjMSEQbMD
0OTqU3XONxP9eP9DDiA95qvNRiNbdgzc/rH2KvPmDZismUwlUsqz69MM2Vcu
UzXtJRHcWBqTxeT8pQIaPx/npAMkD/Tu8/m/05jMC8PiMcYbLfdoFTZGI+Jy
2zLG/wj6W8VW7TrgxgZuOMi45/yCLXg9fpNhEsALbUrDaj+hPFfdyVfWXLgP
/xJ7S1DinUlQRITb8DcYHk5/CoX5fWqK5e9gv8jGJsgUjw18XDHfJk7Dl9AZ
Jzi5KnRvvkiMEhHZKlR3t4xOiFySakLi4d+dQe6XvJOI9Y83KVTgq8QARnEV
6oO9qjZ2W5HX9Yu4IYUeKdw/hAhUp0E8pk4ae/5JMjhmaPjz2Y1sPZ01Y+qI
vsC5aWi1VSeDuury20vPuyS4fiaPQso5CSSucv5fsSnXLJZRFDOLgFn4A9zP
1bt7DEHKrq9I7S+YghX0DQBqCd8nGLl/mFEqWcy/fX5BN71kGTbHxNSqGDag
ZtQDMHZ4rgiFBjfCoPtmBVEOrbsRyen0OfduCDi9IGTw7FKpXQ2QH4RORgev
L5jpEHSzrTtGw9IPnAs9jqFBJJonVLzPScOhSM6tkZC7wviz87ePKxAhV9w3
gEgJN1RreCWRxrgXbdu8o9rt5ZYSEpNHq5E23q3a2c2kpkpXNMLTONrHAiNv
aDI8mwvwHSMKYU6u+dXpAZI+NYPyebV8vhY2j9JZGhBMFSKMrtZOuoCleAoQ
v6VU27zBSfdoinpiKxmLYFvD3/Z5fctHlAAn5y1ltQsqYNCRhR7TP6/Zx7rB
7UYY3qf2Jq2EDeVz2eRnFeI7Pz2E+JlfVOVHAWlikwsEVqKS6mMh1eDU5ZTA
gjG9uDKU86T6PMU0Mu8uxZ3LKwm1MYrlHN00ikrF8NWdI+/jMVFEFVD8gP0X
yMErQl6N1hfZJ+zksfZLF4eA41LTTGKDGhcXc7FZ0My2ynE6J1r1SnP3hjza
5F/na+qMlBDS5Z7P93h5d8sMvK0a0O87HUwbvrA32a2FlzIVS8TjYxaTP3Pn
StG5+enTy75ICGQ4GEqFnxMqkspRdN6VdTtE+TPV8qmeEKQ2cw5VwEG9IV5X
vCLXrQjUSSVxF+cZUO6HEoTfHFJb0slUeCoanJJFvpkck4y4nn5oCRMDcJA3
tSZHtc051lcNXRzFD9phAtJOG0nY/DQHf4vbspgFSi6VPqNNAqu0q/4/CJAi
eYZCh2W3qF6xx6QexPUxCqnWDvs6boq82y0K2MePaLI7i4y0w9jvc7lhIstJ
VFNIutnB/MnrvNtUKbCwFUZyP41DFkLRzFxRKDY4zQQUGp9AydumwSReo2CF
/AbTUt4akSLtL3IU6tY21c0KfE/8REFqEz48fsKt1LWAaaVAuZbeKyAs7G6K
hzPCJszaHKXjDJ0rFN/WrnEkaJxQlu09hVWVSl7iv8fYXx2yHSuE8ep+SwwY
LKRlNe1228lGKRW5cyaQKYMOaHtFPAPMwwCh2/mLRC4RpxRbq1eoazmSvpdV
vEB52n2ymlVoBEuU75ji/UoG/jjzdX+NZjDr7ruebbyU5eJKmo/wpxfT21AA
5EibJeoEFHyVEde73HwuUhf8NUSwkcsTuDzbUdUDgMEFKiYhlc+901/mQEIO
5O3nKsiD7ZcdThVDnWn/d/ciC37O3MF75gec99tlIMr4AsjHACAuMCoJpiHf
/bHwUkqHU+1GyIpyVLF/XxDOrhUf12PzfuWYcXI6W0evWuLjY5LR8fgVBDG2
OTOZ7XFLFJnYKvNb/ZsOFcQnK/0CCk/mDMbs07gytklQ6wl9wsxB8IDOlrYm
k/YPWBZY95zf0q58QjZqNFlnpF65legY+ogepL32kmAnjy3022eQYxasLzZM
L4zuyG9XPsNdw2wo4EBkt06iSlxVW+qQ82f9rNtUa2J8uFqa3fyau9CIfSp4
SItrhw1eT8J43t4nfao7sofp0AnHl9QpFmx8mFtX7oGkZ3iWk0wglC/mEqzB
Hi+Lv/SGr7xIs34iqpAqzcI3fkZ5j+Ka5ZMHEfBVvpkf5WM43Mds1ZfQtbWF
/QE+xoZvuqlxkDr4/EipPTh8Vwmf4B4yaRmNNla21Bb0b98PSxLD7SiXQ3A7
cGcZaqrp8P+8ZLieBhMvpKmzwxRIB+xgERFOlrwABhNr/G09WpAryaHgla5+
jhfloeGPly4iouwpYDv67B4LBa8mJvyss74LrC/XB8wRpZGrsh6v+nvoI9eW
6H0kkGAVhpBwNT9+n/FAF+gVzYIBdjohQo3OQZQsBvWdBkN5qOafcNcKLqZD
scaBjZqNwxSy2XwPyp5+t/8cEzaGqqVMy2eGS4jcDgKTkvg3A0MPm+gORCeW
TDQ+/Dn1GlYTV3Yv14Ga2In4dAZwafmyZxn4QmGUxJzlu89RlJkqFDb6hn3F
v5GmxT22YYcum4fKqU/Exjf3/GDT/hFly4AlMSC0UYeM/LEXjG1iwIjQRamd
tD1OyUckk8hcjOnDU28XJmOkAD+smB92cWx/C/H238w2+fBaAKg0UJ7zVaaK
3YN54UJtsAnwEsAG4jp90gIVIN+1ipknmUZzip1tGBvaYjk0P3ZPIs2bHqgk
kh79yWa/JJ7yE3ozMkOGWBTOxej0f/NEfXS/+x/1ZNg7tDB/iPdjbN7Ob8ZI
vhr3ZS5iX9wEmE779Olsq81lT9rlbTXvCcfyr1NQRy5Q+T3xuNau1sdfq6Qf
giH4sfrvS6Qc66Yg5kQ/6xROMGKcguAkq9ROHp5rHwdgUD2MDDiluf97zWJI
LNbaojVGF+L1kkzgvuK9d1Wb3Li32gnvE4L331Zh2xt/DIKxKBD54aQL20C1
1rpXCxBzxxDAbupLgEbkLwqnev5iXwz3xCj+9xYs462BeElLFL9MXdK6FSAc
AxlHU3kWvMttHRAF9Sxvf3wgNkYzjw6NFCnFYX7UMv38YMcQjtmvmrvpqUY3
yzz+QH7AF0JIEgjS3jU4ukOru8Fz7p/ifLz2Ayciy+Pq0A/+FAU7RhxHwg02
RYcr4TuTEZvxZiCGMQ+Ayt9/NAObT5JiI+0mqbO3yS1OOLKUKNwF7NPOIX0l
Z7D9J/hfYixodv+6mIU7S8WTOweyIXspZ+EPMz8YVHb5L76dvpvCbf5MI4LS
I5/4qrcRYvVhtf+salsFS4fbtJfwHJRtOaiKUXadl0aMud6N6ioWpXCJderw
ecAXUUDAkIHlGE8YAHyfRCAKLVc+dvw1L4pBJK4FtcyoXmQ+BeCUBVaeNLdb
FcYu2KuhS+N4fKunsIfciNQlRUTz+xqB8N8kYyknMQ62x5JtGf1B3BErYrob
5N1HPU2oilI9w8dYsa9wJGjcpcol0emYmeNLXyouqEz4DkSQ3zTtaH2yFyEa
YIuUXxnTtrLyuXupYHwb9ZSGkQyQpW4xaAkD0tZXbdtpY2FQrl1M9fFbNIgM
NtGAy1Jx86/80fu/m8J+4VjzMnVE8St1DYUx3mrLY5F8KP9+kEheMCwO3ryh
xc7M+4aK0N8qXR9yn1z1jL019EKKsA10kARofhZHCdCiQXCq9Kw6Wr9QGIoH
8KubzmtnKN+/eSH5k6MsgrU3r/eLox1xlekIOKGqnTCPZS1ver8BhJu2syHY
c9jHOxpU2g1hI6aH6Pq8Uqpn/y+HMHXVUh4IRMdSeHn7tGMTfwyd5laL8JDX
C/F0DVe5tmO0fVtev94ct0M7Bmixey1rybmQn1K6dXPhPRNL0opPYteBUMrt
Vg+4nHTuXGJT2lb8Al582OCrHfM79vcBhDooPcsh0Hk8PgEC5zURqORtROHs
Ay10UMAc5ECfZjs6IX1gT/+xQXvDDxYLrNuDL6eGSxFVbWUFAuotsvDi3Smq
rcVxiquqXw+D3dWq8EqFBPtIj2qPBx39AS3mXJgDEClX1x1XMg4Yw3h5lfs5
6/KHo+uXJ0OmnBq0lmM0iYT2RRTTvuORMw/lOdRHFydL220XLFYOBJoOGL+9
5oqGJMchGIAatHcm2Yn707Yb8vkjCuA9ONo5N+DwtaRJ6yHcH5wvaw5tYHyO
09XmxzaZPRJXkX3vm603mIcdACeXbAfT2alc9qrr6jKSnWVXUvqBESUoC4X5
Ts8qsjfktNQ0Ww/yFvPXFHlarKqhJvYUUFDOIl3/47LUPVE5yhP/zagd5zFB
WZLR4ZBgOMaCIEEDXRLMXsQUALh/S+H44XcztmSEb96wPovVVxNpVvwBlOOC
K+dSAzsEHlKdc1i7aTemv0+ypXMnJkSKdfyRSXgRdhpTUx8QEHc7g1ppuTsz
u8CMdnZy00uoM1FxzUSS6R0y7qNyd3VSbw6ryMAaMkSE3fN087qbdAO7nzS7
zH2NnSbTxgn0Lqdo/rq7MjpqK1Vsme70WpAH5IcW6UFyZYjtewe0V9JOr7YN
LRLFHMa7g1WmTg3f5dqwsjOGsS0xFLz3eluOeE5fAaUuJaUBMUwpClXTlagi
o90o0bcOQTBuey/ixXwDEpeiirFztkUtxYGJM9cGwb21ADbEaml09EIHSKoo
ag7sRMLAbywJI1QyyLgPb+JhN/CRXBpj9OSRBwjgUw9mzCIWmEg0FE4u6Uqq
L00YDkv/AZWcLqQaKRYsSzJisTtlXEA3Ck2UDor1WWBSuXrwoeaHSiAnLwKi
vKBY2v9c42yZPlNvai5jzHhzogXrTL+Ys5kk4BW/w5w6yfJbcJHEaiUDlCWY
yRkl9c3zxLTogUO6AapsLgle8jRb7YGOhkLafD9v9vRA6HyP3RRQBOom5Vw2
jKtS6v0Xpm4cJZPkDEuZXG+PKKiaHI1uhJhV5hH1Yd/k3Lk/1xkUbtyezPNz
i8Rko4NEX7thuv1f/Wd9mj95NBNk4PcyeYFZvTcGpEyxj04/KRrw8ndpDC3r
WpN+75U/BoRFYJtbzki+mo26sTcUzrchF42kQMmE4RDEETUsvOuY7N+FApJo
eFzBLC9ycXRr2/Xh9GOMLBJ0EMDCoUQ00wOT433V3aJSCPFwFQMYnrMdZQuD
S2bJhcanDIBf7eMYXdKaHl9Uvuyn0u6gFUnBklaYKrCfKHtHdHxXNhyd+Xjr
44jS6P+whDq6X9cr50McwIdVb5Xtv9CeETfrTKWKWBbj40pa2dossSCzxv07
04TH4u6l4NCuZ9IEuQVVPlBcLpBdfa2nEC2jRefHn6rz2dsIFX4y3g+MssHy
ky0YMm8WSdD/iPfFh9Ix0LD2kCyiefbKhyR+tSeI9hmJG+IfCC+o02psc/7i
O6x6MLeibsd8+/+WHHAVAKQWrIadHX8yIqOHtquO8wEb2yhbuu7uiDNXsfba
BvQJnW09L2YzM1Pe/D7TuJXFPqhDryoe6v3rqqbIVfgamlgqQVI2dXi2wlIz
KfW6yJep7i77X2+pUUY19p+LXOTab4UtHEAGXqHv004HEBeYb90wN401rk/x
L2/ybNrRxEHK8r4fEp/GlYYLXYrZ4F3B1boxzSsugEpNy8f+t2HCHtX59EYb
R+cF0D0fLco7oyCLRQJ/7nUYnw83ARIMfrxn+3/gnlIoVQX/166YpnhW5El6
xNdtKEbttrxI1kIx4SzxVWuiiS45BISjajXrbmnrIyDPDE9aBxnwAiUAAiG/
1/bec/BFp/DVM9DkXQiVrzv3NQVKfl/Eyyq/qB8KTcfHmp7cxmzraSafrDt7
04xXXxAntg2wPKaEW5y2GZqBayr0884yAc+qGxhuahytQgIudB4wowm//x7J
pcSwx3UtrXxxJToJzkAw1jZJnQE2Wqhh+s0qIlI/db/jhO0t06qEg374cw0T
VWzZUQjSNv7JHrwVnU0KQ7SM2AFHvMsGj6G4wXWhJ08TfQcK0sBt6eLipqFX
LXnxIMMaPWfjqAvPpSBfhQTBdjzSU8+8QZI/j3W5xVo7UUNS6k3cMx/EvNKf
J+/bEdEkY4l5UQOFcOXVOwYX0ZBNU6lztF3mEe/jWoz1q0xQp5cQWuibN7PA
SMg6xs3G8dmRpFpc4mTuEzW8j6Tt9U5XE96wRrnzp3zVc+tXuAnSpnpPJ6Iy
O2xEPYuY5byOa4VvUBv0JpZMz/GWD1XX7GgQGam9l+6nVBYqYqEj+IbJBHHT
gyVQACHUwaz22GL21zJj/8eqd2V6I859BW/n5I5I2Cp7CEmQJpBYIXJERaUG
b+5PpdAZsdATNgOfzwxvhpOf1v+dmbwi5PoM7osdpgi1INUTT8VwGMMjsEnJ
4e0VByDvgANyDTm4Y5mgMDZ4QDnSjlnpeHtQlJugThcYbry8x8dCIbzUCU8e
fUtGGl+b0kJeWjnTkOwBkEvg6ovOjQrxw5y4DwQpfFuGIR4AGwCIw9tJDLVU
gs4AFOF2F5CnsMsFkBHyqPI0famEkZsG90CYOen1emoIF2Fl2AcQuuanWRQu
tUj1A6divAR9HVWhKbn4X91yat1kwskBGmkMVFRHWV2nha/rpNdGxoK7mmwu
O3XWT5tGq07tRdTJtU7DAoBMN4cVpsVjIRmsoLG8wvlz2BlZ8dX6jAmFdyJv
tjxKLBhmX5D4tojbJTPC4XAN4xaCVTkM5tQ3st2ASY3vW7wHAsU4pt0x1jWZ
z9tR8rvTScRbxTidJXlvhgdgPXVVMLMqpqM33nOtlstNk50fk9ZkVbtJ2sRE
wPm2DVlgi+6VADtPbZ0D+XdDYzp3nJeBb2GLoajZxx/8mTF6O2iZCNo+1iTP
FeNiduDn7mWsKFk7xAFDG4jn3+89iPHMIzOkwDSDJ3QjXte6XxGH8eI9W5Vl
TVsJhczAjp3JZuwjbfR3mujnLccMfLHiuFqxs0nDom7esUQ5bAh86iwBCflQ
e9VVrSeAv2FvQadeQFbOPJuapbljsAZZBxex+Pi3asnGOE6XRTEy0Zh/1g2f
2s87jXI5Hn+bcg/OtUO50uZH5+iUlJsru7RANuCfiLvrashbYBtq22xvEHop
6/pQIelpCR8ta5KdGqQHr8jkZwEmSPs7KPn5ljbPUx45rIUOrFti2eW/Buv+
3Tu37whDyjzMysrhyGi7WF6+TRt7/qeeBfA7pB7PmCr35uc2OPjNhjbf3ueI
VclVDoVDgPva12UmZIFXGQdQQgMwHB2h/fP+r6/sYpq9uBhaLCXVLn91hvvZ
la/7XA3QPrP8mpNPd1iaNBRE90+39PWP6ne4acKty0VKJcxQuUrJEiPlRUR4
TI+bD5UqmcYuKpKNUdKcMoT0XTcopXPXo/rO6KNxyS4ejTw7c6I1SJ4ftfl+
+Lv/p83pyN0CL6+1vBvFhDdZXNAfnfRdvo432aWi2B81HRavaXUWaUfagFLU
pZiRfrj2uJhbS7Aib9sdIAhollg5sQM4LRzMmGdqxJoGAUxnKhKVhKkcZ9er
Ecl5ABtGjK4YD1KNYJ3Yf3X5dWOqZFRBgYkGCj+e0wBTrEs87h21ruwn8cdq
JZDS4Q+LZdl1fHMfrC87QDiylkkTQmJggO3u2y63TvTii6/GMPMhYbncdjRO
/1qX/663O+NkhcuUIwvh38ZJhzDLp+xuQS2gF3CvRirVGgoGu4GRKWxSQwIA
jXU6n4SKCCjEHRLu7m3kfrPmqL4ohTFa8KT6dOpJ76ZIe8bgDeyL8ko9EWAS
e1uV236fI4erUmImxoqKUBzFnakr5IO8mUnd0yglA1HSFbjV+hvjf4zPm8ds
jHs4RbiO3XuLDpc6yiyiLZoU95dLfY/DwmMwctZagNVWN6mRv8eJEZYLrJO4
NwCgoxkgtWLppIt6gyMvyLU5qFhsJ4nlxZQdKYKhrGFs6G3Dj0MZ/JVJVMJl
87bjj9YhGs0wRqSBbmayzpDBrYAO3LZbZl2T5b/uRXip0LnB0h/kquCimZTS
qumxKP5ySGGDjA/kV+ko6rplfOVWaZZiXvNflw0DTgB1qyPF4mdaXFzFjnsG
PIpXUm29Dtfmr5/sVgmOMTU4Q2xJ504NKajkxQZxbzDarYKPox1vl9SGiF6A
KiVhdzldVw7OWJSz4orDLWpGN4plhG8WgpGq94E3SBdlTWLyrjc/PQdKRE9b
/dGfXlKd7NV268du9bQ/ZWibfsYHRnRYuCRw/VmhKTr0fTg+B9PRAMMDwCTi
SAY6rniaLPCWC4RGdHj9yJ0r3ICKx8XF/FZMrsXbR1MZ3EHrrtLosx7Hw3jt
QXiXeq6Plwgj8co2RNgieujYaROwlI6pJ0BDzI/ECASezdMvNuc9B6Rg3kEn
DgDOREZIOaf1eSAbyv74IRBEpwC7dWpjr6mgT3RcAk8ssFDVaoThWTDF89Hw
C5++I2Mun+d83t7UKN9vQk6o+vbArFuRxbd+jFFjL2tTm/D/TnOHiKZbSrx1
ge+fgp3XVNS6sPFyMcmr8SouApBANyeyWT7BtBjwEIYR8/CBofRrFQoWZ/1d
ZdYLNnawP4u01mOipOqgCPvBOe3CqRSHxtuMvU6ZFimBtocn00vMvl9VDPr3
Jcg1enHq2DuRjpCBV7b3xjTeyQW5MuX4Tl/waKlW+sAALMfzS4T1XpCVVEZl
/0H3Krv5RjYUaiBj4vyUsG6nG3DC5mdy2VhAQmbItWD4+n+JLviV3hXz4IvI
uhDVKwIciD1CG2X8vk8AMVY4FrhspOxrNsbNIvcXfzDYPItUKJy/dWLq0Sg7
wggUjeFaAqQj9p9L7/Lnttqlurd1+AU67uIX95rDmG3zr+N+dEtRS3KSYr0u
pa/Lkh8nMtygB52SyAQix4uZe/xfrcHurpODMNkwdBPfBLXbtw4SBB2i2xRa
yRIP38FjDZNYoZ2cqiuVB7AjAMHhuv9b8kjtxmpMHjXjIn+Qprd7bxufvPp1
OEOQQCDKVSRw99yI5W6lqFtdQ7U9xVP1U1T4ovAeU5iRFk8AtuvP7iCuAqR/
3kTxInzo0rfP58znw39Sk9QuQIBri7XOgJ4C2AZ9wro3OKUoR2qU03ksqGHm
xV3OiThrr2KdSwgsmFOQhD+AS0CYs0NdPa3e040JpID1F/swutqTRmkbPUGZ
gAGpFHV/hAMURVZDECRFxFGRKDf5exnwCZCLv3s1bPm7HpoFQeKFmKDS1Rn6
DqQ9GCBS2WdHu8rdfcyEYYGxigUCUCfYapaJp3V7vZzE02mXsabyPaAoCinl
1BH7FBu2NP8eOO5p7D+yiB8+ihoEnyMpsstRmrz7h1jGtyJzxb4+3PaPQNsU
e4JI47aJd1n2kEaI1tBrfpU3yhMXi6Y6pG57Z53FgkXd/fetUpq+wHEKzkJv
dSqX8lVia7jnTaiOmp/tkAcHHSLG8tLhtrAu7TvwTXa8I8z235BBWhiSkVEv
lno62QKKzA+5xpdKGnM7v0x2fw47yK/BErW0K0skh5ejw9f8ZR3YPht0lZwO
n32HR53phX5Gjjq+R0iWMgX6ILX5GAeaP+WHa8qx3cnLJUN6Bus3oJ8JLN2j
pYdb6w0xY+bbK4xJQL56t1bR/D+yEPmaawgwfcdv144b91B1YlUaVNoNe+Vf
hTKxE53fxvngAsKddAb2RRtEYaw+/KleNOOG3pxcW4Dqlk8csK+c4gCoKH22
dkChSNwu8KpVBMaX/HUKaPg1vxppapabJRBS2c9fKHefs9lt/i/94vI6bR0h
bYPMn6p+X69yamnV3V4qoZpItW78G+cjawAOyCkkaahDl8cwIRVEZSw3WDYX
ABl0FHzvuLTHQ3p2Bh99hOQe8WofVUv8+7zSkk9nSgCZO5WXEueaFR/yH7J+
acgmCKwf5MT02QA+DWwA0mo3NhyLfDjNoj7tv/nSHlSZQgTc7H/IjMfKRnMX
/LiowstoYjCTdTESc2iDBHe5fpVa/M+czbykKh9jzwKd6mepq7meauq6OUSG
y/vy/o6F4qHhOxYTAYO5Q/H7iruRo0otOMCFJ89A7RRgyA/WEOcV9zLCow9h
54MaGMmjKuZjmJ5C5wVWA4ctqE4o2FXAaLIAk0Cpqf9dIXG5wdp2pxmxB6gk
F5xviVFZWTpWaevaT4nKcvlqH8CBwAz5dS+FF61y6U441fGO5zhoJih+wYD2
h0QSI/ncFSueN3yYC4qXjWyuAAJIrMiYnBmFLdWDaG3Wj0t2iGJ2ZfrrmcGP
nOJeQfFZINjkYY8wzZwFs2ueBdQsiOUrDKxmd5RpgL9tXWZyB5QH4h83jPwo
X8IdCwbyXRDpPDxbbxTtY1H5IHcbcBsMxxNTYAEv2yYZH5rb1O3xm1rzqFxI
upOWLlvZNS0HCup6p50kHWWv0byxtiF+Leuer3hNTKnLz3ZRTba0eTOVmQny
nmQLQx5VaApEMKVGlvV8ruFwq3vXCQslOAUrDHdIowZIwxXupFCi2jl8Qnxy
kbdZu2bDfynRWnAecWwtA/ftdnSBmxn5Y2TfOFNy0M0E/Cn755u8zzrpowHb
H4uoTX8iaijh5O2UWTIDlYUlufvAugxyEAatNWL0Cgi2hemsNC8nTyMW0VbZ
mjwC7ScNOdykCxSzaRwqDayAnvarbjMaTnNKMHAShlGjpDaqTnVnUevAB0qQ
KwVqmJ0i37xpPEPkkyoZpaAP8v9Dkx6XFUkeii1BjXYmSy0/QYNXG1rYsdKP
PaNEBO8pBvvhNmQbwEk4Jt68wWDjaf/LS8iRNA79NArTJaSmw6MLgGytjz/R
MK3cr5qUT2bDOP99euH1TeuRwPanb2u8AYEoWEtmjcN1A8Ixzz/YQUNJdlfI
m8A1wk3x1gfzREV7fdgEdlyfu9wjKZDhqmbPiM16BPfiQRfALU5EkdlgAp6p
Oo6gD4AZJkYxdq8hWtJPTTvtZngJZ34nWjfpw8MKN9PSdP5ERrr9oeFUL1Fk
aR57ST443l3ycbmiPSIStZPsjIjuFwVY+/Zl9cc/t9WCv5+P0dKZZy0ZE92t
IEfgkwyBEl6B0EYXs4W+DR5Gm1jogJHOD1Osie1hZOZ5CKmnPbXwbHQte0ju
6mh3Rw3aMpi2w/eg1saW9mdDNBiU0QKK62spnt+FvW5aX0E1hDZJ4ASCQB26
2ZkhsSPen/NLhW1hu4WZy/GqHJ6xFJX52HCZgayth6d/MTFUAA035iinYl/6
hhMEaKnNWOL6EtdEqeCk2/gfNLJV1PnycJWBzT/ZcJQiO+5pA6NB5Us+vhip
WWYtnmnXoRQZnMPfJJVeUTvC16tb9t19il3zPx/7ARPl8s0JudJsop/iW12a
fkrA+WMvqzp8fjSeR1b2aTi4Y25KQtpzYUfvOU1oppUtZ3ZsWaS/Yg4XrfDz
34g0Rug1e6sta69UrPbC6aXocOjp1v6TGXHsTkMCNz2uv3eU9qIq6Bs53wq+
fowjG3EMzYGtsLhQDIBTsdtcHj+15SkBU6NLcQ2SGn4G6Y0vYIoZL2tFssc5
kc5hsLN3fDq66/QlRsu3nEQ3OcpBgJO47wCYJf9ll67Ms7XBxbrtQeRzNpGA
1a49Rhh9EqF41ou9neMaQemwtVMOf/Xk42FCHvnmvuuvkT9vxQ41swOuoG3z
kJMAoBcNPcTXP/f+b8jnZAp/iz+joxpGXhXytgmDKxiKJyZQgAJjBBOASWw1
/Xo37Ri5dUDAIeYnXWF2aGq+JCshvK/G3T6s70OitHtpeWfrJfBtcr4BSceM
NIHtNazBWGTkzgzfWWsZ1eqXqgnuXYfXpFZOGytMtLtvFvPM3LNzfbyj7Qfq
5txxXPCoiBgwYyjAUfuOD1fTXxJvEyvy99nP3zEOOSgR9Z5SKgDY1ioC7d3p
xXC6d523BniI8iPhQxYQWQxbWL4wgDerKes4ghU+zut/Ohh7ABQR06BjToqd
y83lr6mL/mvF/1ymmRNNTWC/edZDlIkcq/P7KV/6CKZgheJVh+tdH4sfZ1DB
9wGqyy3YeX6aKXD+sJfmZDMCNHqMjBNynFia1EBXZvvkY3HwkgJDWBB/1Xon
gKOKojenMLaVGkx6iBU+DOqvppEXc6UoiBlpV0zIXPERT7wxOcyNZvd3bjLR
4sRen4taUKKRR+LtVNB3+oQICnnmYN6ot8oOmNYTXxkQIdlu7tohg8dlpL4A
3Xi4WdBQtWLYMtX8f5Mn+uoH2oQOif8uFPuuzXqMwE4yn8iyBbgCQSZBKTA9
IB6fhlPjRjAeUZhXiCd9rp7Ld338Qe+NesJG1Slc04H15Ul9ZOZnUlSQch2W
ivMEEdQch1bxeoChauDMzL4rJxq0Gl5DojHmA8OoAvo1uRZuLr82RX1V/PnJ
GR+xLTRH/LcR4jtKi7B3zQyeEphTqdbJwM9XXXGvriaFe5ViE9yky4Y9xx0i
CesshnrblZ9hD49mgeKxrwWGIHBh9/RjwShEvBfrmP2iwtaqR8TPhW7lSdWb
8Unrk1xJfW4E09GsoWq7RS73tnsdGCaoX8ZlCguEs22GHtHuSpBI9U0EZpTN
9H4WtZAC2NIF5ZA2SHaNor+QkAkHK0bp17o8S+n8Vdz2J0MiKwFcfezOPXRA
HI7RbxFUqqBGThNrBCJ8MXkOzNMFU6rqJe23jr4yOd8ky7qli/M6HZ0rsu7s
Yl8QgtXOguO+O/+bYYOI+Qlie6XhxSdpmkoSYS77p2lqxTerYAelYHkOJI0z
F5dbGOQigN4XmcYkiL+M9bqMmIdI0V52tSCoLfX4oabPq86kaxSE6Iy71TVW
mVktSV/FPXcBmHTkLjnm6cXongja4f6WLrRtJaA/QKjMHDQATLogbQRKPln7
Yl9di2rDv2tLPY4LmGRcAu6c/tyaKqK7oyoxbbZLnHV6G9hguoJHi1zsPh3O
PtUxOFh2kuq/0SOujfQ3brXjhIyZmQ11C1oZ7x00ar+9ZKvNBYm7v5utQFRP
/Q+NinyGGUG7LkH1CHCvtmbvFoIyigJHDjxG7tZ8FtTlD8khEPgqFS2+4ZpW
72ToC6K6bVJSnNyvhRiqvHg0MAiVF5VjumyPPXT8oygslNa1BaOsORWGdbbV
Gq4HxPsqHXwlvgAQfssDnGYQgVHiSJ6oez++IbP/6K8bGAjwYP2ObWD5+8sx
w/R6meuI2fr0MlgqB98p/R4Fk90uX8CjL3iOEZdrxO47ZjD/f9R+growbb0z
keSCa6LRttMG8inpchATWRmvqOa/0VaJ11Wx+98dqB2sM4dO5/mmw74e4m6N
tUoyoTXtiT/VhfHs5VIwCx6F2pHHpuSvbQClLWAwZ3IizqYPMSf8XCzyWHW8
K4ij1dhYUeVxUqQLXqeyA83kdM6ERmsArj5QchDD/b4lEdY+uKtKk6t73JSz
MxhMY1V08iVnmfardFW3+w59oiGaoXQp+fY88Y0e60ZKR5SNYE9/WDHYOyUx
2oeHDkTZ+1og67iN4y72sWBZo1p3N3Mww+YeIHVgN0Rn0IgXbsTHB5TjRkRw
KnJ3GQavWs53K/wIY7HzRbo+5ncT+UZgmhVNlFRqCWBDMiFmDE4k5lYjvrqw
VQ5oFA+98GIH3LnA2zJAoag+gC6f7mY9J+nOoEjlPpr5PWSvrMh2yUrKGbaz
jlr5eAulcoPJgvDAkzRsze4HsnEUr2YyFo1PVTzEzYLJwmofH2uTkDFPB08y
LuIcbKSBJCXtcmYhDt7Kizh1XlEnAOUUiFrkiNCAjmUrccZTXehhvfik+jED
Kfr95v88UQSZAC40ZWPc+0cJkrPTbkQ604o83hxZXy7OUB4n9rfVR4I52H2f
CyKJybYRQyvz6LsAhXGbPTtz1Wwex/43YkshbwgFdvLdlYS5JLSfMvjR/CEY
XyetliKhLLf8gSKIosq4fb6zPbT/ho8y/4FDZKrelwZ3UaWwS3CvZJVAlZ5r
83jYIMvhp/jdzmpKPZPNl5rAAZtsDW5lhVZrTb3eHoQDOE5xORYOBGyP1YJc
MN9K8t3CS2eA9++SENlMVJ+Bg7Q23eBME9XCQW6UVToDlU96V+sVmvwKk7Ms
/4SPGJq//EyVNSsCkYkUHA8lvFUhbPrh0IsqcYMXypIkFlZHwl3OtUQHsnSV
aDuDNq/NA8ynblrFv+jCFGVd/gjLc/ExyegEiersdYpBgOhWv1TpVaXdjLtw
R/Nci+HQiAvkTGVj1ZdbFND50WOY4WkCcqP6JeNjBV/pGtYIOkWUskho9UVA
q669AD5vfhWSPAd5l5WV3cC9H1K7+Lh6Rewkfutno433wh11Pmbic7nO4pZa
cNaZ8K0sMOJaps6goeOrTVZ18VoC3sPEyj+tqq5PXc39IAv28K6Ui9o6u+MG
xk0Jzb46C2fJOoL92f6wakcf9jrS4VV8KNQJG5DmOc2rWF0fCTSLsY/7oWpI
MMUFiYy4dcDQo9NFznYTcVZToz0s9U6uWYWSPU7kJHlmMRhnLgtWTUmikdoT
l2RDy8GdCCskJdoRNEqiD1fha8+G+Bh51N8NDlWgdCT7yYNGscRl329dCHW4
zdI3fsCgGO5Wv9W8jIQ/9I49x0My3oxslGKeE/YffBAAbIJ2ZRr7YAIm/Q/5
3lVaoBdEnqhjs4qDYiP5NkZbpKEpBg6ySk9kdX8EWQ/cwoNf8779oL0O/Zdq
UGgmXxqivTVLttn4Bs8bWYGaVbibRuQ02SSiXQem7kr9vN1nwp1TnuSMIstu
DX53xMugR7MNUTtLT+hofwCYOI/9tMr8i0REZz7tJ6vz4gT+hreX3J2co8O6
5Uzody40d0DfSszdTWQTu4L0nrKMPbTcLkiCrSF+lF/CRhjBmiuQfQO+uHeG
x7Hcsa6JUYiEfTQ80oreVKULjTi3T4ty/vUKmbhtl8lwDKftM2bsSG2mF6SW
Uu3rfTRx+SNji33Qx5z5EKJP6i6LFsJWsBeJW1dw5k4w8g28XUbZQAA+584+
pqpmkpcxwJdtT9he8ajntlpLupCg5+vwPi7F35rlLLUXdpKkpmIO8mxxxeAg
oyn1Ww5f3U/b6B2R/rT7XiENofzNLax7tIluJDDxi88stc++XCpcBtyxUsol
IflOLbNwmPGW8m05nfo65r2ZD/DRi8Boz15XQS5Q6zkGU2c0ql6uwS/H/arH
0UMpIAKRt6EBVR/Oa+h/Xta6Pxqkdwa/iuKXVGr8Jh1Dj0+X+FcljwtS7STO
ciTOKzHyMRtcYEpPjzJIhXgjR6DN8lfu1gff8LRm6hy0M9Av33ZlY7W9eP4O
UxDadvHA9XZWgoIUdUme9es9GA7dCpa6hbZU4xuVnQdyMOyn672tz3JUBkoQ
0N1eLWj9pCib+va53v604xZoJj5d+C2Kshfzm/pOUvpdlRVcIzP7UzWD3PmX
+N3fy9yEqr9ulmaUe6HSuPRot6kowm+vc9TKItdgrlNogXWnRO9f2mxy4+CX
IbID/t3eFZzEpgUrfH8XY4dGg0gsGEPaaVsEgY5vQVGtV5ZyR6FVBFiHaFZy
9xgfOFuHWYVcNjPHNf0csJzH8M53D5HkGL1NqISc+RTPgnFbbUQdSLFHjiV+
Ga7Ms+vGdfy+sYhYZUq/hR0eICiF8Wv7K5Bg9tZAxVCkXBJj4g+yQicvfXD6
ggE7qzICYHo4VXjzbAebV+wqz9Nr9O1Gt0Nw7DcdVvtiTzWd0ZafMeEKKjQl
dM2llNWQB5z9PxwleTmXiPAfFVHPBEGPb/F/uz2OUit1mkFXwyoT0NL/5xVD
GTfZBpMsBoMd1/OAMq6pD/t1WSSbrVyuLoCApO2LSMbbUPX8L/tbwK5q5DSz
5xp5JP+YDHE5nN8L/YRp9UT4DAt9QmHHjteZZsHgvlBCfeeZv0dK6+hrcWCf
9UmZk5sWuUylQY5I4pondBEDwJydMiW3nS7XRORZSdUa7UlLMNVowsd4REkm
gZiqz2soRMobgsihd+zVaf5/9LNbN5S7bUc599t48c01ew2/YX1S+JSA6QBq
IyS6fTAw9eavHZZNRahyFVsEFPoIYtG1QSviu9RKzdi5tyfD+KgH+tyO+iPB
4leaXHJNt31U0ePRwnVaZoqIovl7pqI9scCtp2c2oFI1GkOCuG7FZvYHM4jO
CMt7r+oY6ckCok0eQCt9f93emflB3P+vnDj4yr20lv0IVlpS7lAKpq1j+AU+
qbROiMJkYvrWLOYJif6b53wT8F3HXR5/S/RZ/hN27+5i+dYj1Xz8AZj1jgO/
BLIbuzsti4+92kBWGxZQzV9hdVd0+n4ibPyjU8KvMqu1vU1Rb6oJpUbsZnYj
tCodAJrIFS7fCdOHpNRMCwW2MjFBReDln6I96FEzUo8bJJWvknZ4oeyDJuIe
ELyMqgWUsec8vVeMFqKCYY5DV5p20cS3VEIuzWAfCN1IxAiNpAd9tpcwpSQK
j+Ck1MZTXN+P+jlnlRPFkdbhSApQrgbcuHF5zHPAaQTOvEPcOW9y5Nx80BHI
GCKjXE/56f+lPiJcQdGtBZIv9QKvZFaPmd8puQwggRO/wJ7zlJ02nwD2s2Dd
6a9h8xDC1n1m0y8cgM1flU+0duEF4fXODvyGbdKb/Y4SLeBz3WeKHUGTjF1K
SiojRGDtB2rwGWiYtP/M6OPzdwo2xY2isIj3pNgqRk7xMna1MhiWai2vktQB
UJyMd8qGAz3yr1FNnqaT5AqdZeysTwDva2Hx9AB9QSrl53pRphbbqwAG7yN1
ky5COvDQZ3gZ6Uif8h5jxJmX3sW3RkOj2BB1IjvStK1jOI6CfDMkGwuEajJI
fWm7LRZT5RSazlCoRjUpFOoKLQT7t9qvY6C5yaLSd6Ulq98cC2BGZAsGIHS3
reITeGsHYrpW50FgQORb1rlbEY0LUixMaddVDyjp4/XEkjQt+vJ9SsRlURFx
GTvzujpFOiFY7HrzNyurAJRapynRM3U6nGLyyJiNW8O2lcjXemPNk+u0506I
DNCDTcxDjTVjfIDZH9yvL0FGJbcgZTsp6KjwLBmBdz7hcQMuDjk6iCfe19kB
z9UD03q5zqmnXNhzLOyh4RX2iZfIBgbWdKZ8wyQqR3jScnEddsZjpdWudEZ6
eiw/PP5tmQCf0xMPJOJdIrX4tvvNEHfBFsT3wNsenih2ejsuLq16qfZSR+2I
feClngXMgnRGs/U+CQqpJZWyfV0b7qblpcfpD+2bpGdwlI/A8f1Zf+N1MK5P
MwHxwdiWcE9mrLCcnYI6gjmBMqdAbLaCVb4n+DlBJ/s2w92FAX9a/AchZS5l
aK30akBzvKpWkzBLudFtKD7meuXNC9vte44ii/pKxbZ0gaQotm39bNvuxl0A
7muns130hAT1KCm4zxgLoCT6rFCPAHTHB3qE0tPAozuNC4yohu+08AuTDfmk
xxLJKY0jciSeT8c8f7yNwr1Qvur8rCZQ7Dw0sxRo8r/6X8fqh+4rn41UNZB/
KaGjFWkHcsxuCkOVgA8OMF17JuVV4LboCNOiLgkJ8FFsgMf3vlOSTVSz3fqr
qvG+Niac6eWvXCzVmJrfD8sZDpFUkFNFLQSzntF5iSNlhBggbR8qpgltlIlw
0+aiYP3y3Ec5vKP62LBtEUg1ddRySlieEC1PG6JdckvAfUZdE5UJ7RKPxEFK
DEVwl/t2weZupzXBXx9XMuJ1c4Sc3RpkRju87FqNdjw/2vqEjWLALuddJLKR
GYZAEC5gRp3BGMgNFRZAHkSn0Cfm7Ykz6E7KWBLhyTN4//7nqiDdYbwK4u/f
Z44qRdcvCTlPGp8u0nEhzOrxkJ0hJVl/WO/kVmERO3xn3RNwD2XWgE/R3JqV
+yUbRXBjO53vcGdvMwAfedGig5k3u9vsCvYNplJ+0GL/KLlz4rd9PhkiJrp+
9br+92jwzUCHAs8MOIC+wB20OK2u6CkdfWt1bg5Mh9vwRqVheX9VYpOJm7a+
XTaLy0rlhNASe7o3i9eecjUk/YduJV8hNIf0/xt8KWNHTnjM1F7AP1wpgEDD
uuLUIW7p8x0xI3mnFnfJ+wxM18G8tJJnrxa8VzFGlk9juQUpx3XgKTi9uh3F
3Tx3tKsYlpYkX5yLpMT8THSnzuw09jPStqXfZ9U8L29/UxgZ0qS0gx62KZxe
rhPozOCPNzRnW0iuIukV7afGqI9bXoPdreQdiZmPRCPY1y+00wJmV8mCiuTH
71kOeAXqdlV8saXxBuhaymdR8AdOrV3GDFgbsJFcem99wlrfaMTHk5IbOopZ
R5cWP7uXRi/8MU8oKALKMuMCPTTmZBh7k1pliJL+eHaKV/j3pHT+QR6DhMSY
pRMKa2KKN+oHiRQ9tn4Nsem57Td9pVCzt4gArMEgt+SXnLntbx4gcs3bLYPD
Yo/WpNECTdvyqtQDM+HSaVM3BK0EYo0rqJRj+guH7KWi3jlnnuSK5AFihRBL
wlm6cuQHY0CTpdoG5+oTyKxCXXR1MEH4PesOaLLiELC3rHe1pVtPJe2315fd
SycdSLD/Mt3lok+sB6RnZXhWTv5AnHXySeJW7Sca4lsnemHgfRs2HfqHSd9q
kL+F0yvfrVoM1nZqk2tXArcVXu7WpDNeGo6S1uZXxiG7BQ6yzAPwHYfWn+uw
xKvgjUIedfUd9+IMTZsuR8t2lp7EJrvRyY35ROHqo6T9GcaPfMp7WTP50g53
N68AmGZyZynWDkO9IjuPO1BK8I8OqDygZv4EXyImywQTIGX4Ur8mcjPXoRZF
PxOQc30D5beG/fE6cG2GpocugXThbYP1w/70HQr3Sd3hn0pGyoRpYEfxHApS
b3mOizSrqOSTh6LNsfFFelZQjxopJ0DIlgnilZv14BAan6H4Y18neqlsut64
NCLuscP1cvlAv88IvVuXag0R4QzHYdGaZDA/PT790bAId2odt7KM4LIFk+fO
GEo5fm6LiRoMxtZjVGkBTtL+iq28xIPA7uzOzIVyPTuHQ1PuZDRH638Hal+z
zj9puAbgIvpN9pkkbm9Qlfpp3ySSBhe0380RYi5lnu85Wy4bgw8AB4hRM6yx
WaVPRKPkHVRtLv3kYOJiW9QE5TA3MZl2DwfapO6nLskeRpEE/QDCb+LB4vv3
6wCx2sKpJE9yVqQzC6XzF/W6nsxi26hnObl7JS04ZqeMu0U8p9zBrDeGKGMk
3GMGCL/micWi3YUjqp6Iay9t87cRtjq0okv3Yt400b4NzdSDWpPzO409JX/N
Ff7Gd0Z+KUOxYkgKLH+kvXYiMMytew8HxcXXaG+G8leRhJCCLK8wvrJFDknH
1U2BnfqFlyDFsy+GwALt1J4dgB3c2bZaBA/BnpruNZ0wA4vgAPxpRWSEa4hH
dtHt+bn5BB6wTv9RN90jWA1sTcL3h+rvTn9E5eJQ1Jd21V/NqON15CL6NUEy
j9GmdLwZm0Q1vhqljtbXrCqA4TfHIXD+52XGDkIOAy6LZoeY8U0I/ku3V8tl
oJEr9tLl8hQkv/5J1VVkwNEYcbAUAQJoC4qPV1fThtacL2kerSNTQOu9Yt6W
0y20A1w9D/EGk6w5t3sovVQcRfrZBn8vdkzZUtjZoDNfDdUIIcK0PeBXyt5M
98Psr4tXhiftnyfVm7dAdtLbrZGi7VCxO4B0WbqIV5i8E6bJeTA8C7QywRL5
B2kFlI+yNfk6MUZpewBVMsB2/ecsZcRE+ssayhyAh8UX2Owtkb66ytzWZFu8
z1lStsXdvILo7wwvIexCmLw/JUIHoN5DSyjPWbRj2N14CJ7Tp2/LYiKOD2RO
WkAza5DiSvYOasCV0KZGXiFZhNO3wV1VIodj9I56jiyOu5axNwvOeQbwFleC
lxeYZy3mQizI6kZhrggG9q+g/pNI8c2vr+Lj5pjuG3QdyOOEqkKgreMPRZJy
CpqecJfQtPR3WvCZj4PN8XCbdEKOvj36l038jsvh0zf2MLeKXQcpvVm/agGm
dCxGEaiBjsImoGNZ/EEYmb+//4DWWiZY0fH44K8zuADQcfOyVT0z9X14DvFW
HEqS5XCV7628OrMDuLIK61Bg0vmn8mfUV4bsZ/u44KBSO/IwfRp+O+/AboEN
22XkaGO6kNCcnNDW63PI/rBB3Rh81l1N4quaJ4rUzpmeT99exn63jrSWq56b
x8DLKmXpVAhMAQi/RZATY4ecR2DSgnVVEJyex1g9QIoWhUucm9JCCHTUx2ph
n53F8Ys7qYAQViK3KoqdAIB0Dby8VKIJScWRj+oPaRACPArEBfvCd/iJniBc
mtWx+0mBAUJ05FE4GSYlCv3hLZCpPGrBsUaBsvQ773QN3P2N+6mz0lQ6MV0Z
WNGx/AkZlGvl8JnYGsxYNUDW7wWHDeWwSnRy7wH9EBeXsyin0282O6WiXW7a
GIO6oQEqc6gOJMoeR5NSd1aA0muaCxBZp+PH5kpmWA6pIAOfX32mXRfQajKz
QifGjRar1msN7T7+4aSLCf2o+C68cRSW/hqCDiQ/fbo/1Zhk6kxPSYPDbugt
hlwnGHyNcM3i71iQ/Pd3fqr9nNXFGCQIlHpbyd6P+FPlXTp2z5KPLqxUtWS0
QR2ZQ3c2HTGw62lOlDRu7hazdIL2JSLOHgUobilVtx4nj7LEzqLnEwY9TSEH
uWAmhbmaHwul877O0mhpjZ3Bs0l3zO/8YDAlnvYEvIxbl4NXhgESS9Uxtvoh
yhA7VkLXJlescYOlrJ3NpyBddFT5HY2xamiLKmmIxL8Hq8UCYK+cJgqQIl7L
NSYjbyMxn5RSPPmDuMSEKAUTaPH6D25LAv7NQjyCdi0lkzymzhj1drnbpZia
glYOCH1QXUXDz+jniNqZho2xqhJrS1pwGFGwiUXziY6pZ833uirBXQNYew7u
L51TBw7nrELZ9nFzz5GZh0mN1XpcdFb+Zf46SAvLKrYUyZLr8UO0+nf1ligW
vgNm2baiVl9r0GFFRWYmuGoSD2J3GnKKDmIl7XNNoTAmjBEOrftZiCJhtVKG
iS661liMQTwjRMpAsl52WW7X158TTuJim/6pQmpapKI0okGkhSguaO86aMks
zW2hPWbPoswt0rWUsESekE8RjiZcYSEawC5o82i+xFBMOv7bHRa07DvXa7Cr
eOwnMDL3SyjVP+cEFMccTHrSRxYPbcgJmY0wxXsZqDGNwELPJ6zvgn2aWxgM
hecHaGnIsl+x8K0Tt2Bfrgg5syteWLdPgkXZ9T2txq2QGujpDJE/sRsvGiCJ
PsUpUI11qfN7YB6LSn3+fmG4umUjpeBb8FLRLxF1p8JuaQDclB1xbkv2vYI9
VSS7BUIqlUjr1FWSaYQ2arW8avtasvtbW3Fs8wpsNs0QfKH1isINNIA+r2qQ
x9h89oozPBShQJzRSJzx7j9CwBUcEO9wknMLWGlfRpe7PG9RVmjt4praHVMV
hhJq3HaDMBUYFMkrcv7BoraxDmY8M2XNQvtzAJrZAYzm9o9dfI7nhiA8Dq/Y
+CNKIEutpiYjqY28k13vwa8ZUBXjlNeC94F6G+yt4ktcvENpWl087g0uK02f
RV+2yrkfXescmYSBl/E7Zwp9rlg65orNZrf1Y7eKuH6edV0gVTyTqLX8dnTY
oB9XwG+fmWdQfkjWtHvuVM67nNlU/xOAr8aroNSc7FWrfMk7dUk8d3GQ1sbW
8Rh82ZmPRR1k06gfr18jfMLDSpLHKi/tJupIKHIWBZNd/NRBOpzZgAjnFmbn
Xj3Uk9D1B4Xht0w9+p+ZzuH0eKpOEWyVi7i0taUqLTCp/q15tBJ9uuaMbAdM
8G4v3UcZvfs60h8ny5z69Ih1Cnr2ytSvQHSDQh9eM5tvuBnyfn+aHM/VEvyZ
HvpGP5ZrpP5IwRPofU98OoM8Yth8CJsWD5CtBjPBIYgDA7fdvDW7dEOailiy
jPKK+uU/S0nlfXx2nHAeyruTxjDIJvpu9QCBvZWf7rqiQ++Tn+mw2kqQ+6gz
xCyDi1k49kJ+l3DuHh8Ci07lga7MCyMSiVjEtHOxZnJp9tbLZZqIkXHSQ2ME
qhE287aWQmlrn41u5vmcC2a3+Fo6gFG1ypVn1tvzrPdq1fSkYpnI+lJVDhsj
7rAXzXCvK4+m1SkSFbhcALAWaxqVRTvpt5tFjHt3+OK/0uxoU25LualNAstb
OqMjzEN8JQTnHqqfqmYiDCUsY6iphKjzp/GeCxAvdJA3tTYLTOFbbGt/l1fN
JY2AKXZIeFawtMmbCWpLUP52YQqlyflqKOjBxIdYVV5dOoN2ko7Q1yCjlYx7
8k7RSW244csFtq6+4IGBTWqKSJv3yV8PgpOPUIQgsvWtpS+9F+6ddjWkFf3U
/50J4Lan97CoWgCHsA1oyIkr96eWy/qhlj1gtoaHIoCCyK20sicznlk+L74I
Q51+52ZN5X9jqsqCxGg+eh319cMppWbENTC3dOU9JRkKMK+g48Nu0iF82sAn
ZXnTwZmYkywqwuH7YbPHyLyUWpUCtb8BMBJwa3+EBgs9UJIch/wHdOgiGTJ1
1PFs1tMSmKZhiKvf+LS03DdOIPDWQ01aGECimTuOBeJv7ObWlnWmWRI1RMYL
1S1skYJFYyWYWRk4dhgGgxAgYA7+AkxXVoyIPWI+9xJeP7ZIOeYO4hHZBVsF
wz+mPAY3N2OeqlXQT4PGEy6cmP6/rYJRNYrEA2Qpdci+ku44PCm4FE5Ep1/r
FGPn6Gjt1FqnRJKRu20AcELcTcK3Yas0b7+LJyy036vXLTWz41yqaet4pCs7
l63aLzGBvw+fXvxo1yyVQnIHeTnYwAlUTIZxysIb0MYKIjQNZsCPCbItEMPH
FOCKpfAPcOrBRRpREKWIT1BozQ/xMqbEsMX+McmdxODSHbisD07MwF09aPmW
h5ctZxdU/VBoAM4Soobk2wKVGWl+O2YcbG8DT/PTavJNe/yPfz3jCzrd/jIL
9Je2K3hKUoEmgDy8FweUtNh1HRS6NAZLxREs3fH/pkebnBEiD8k0PL49u0zD
JIpD2BPKky87ZKTKAgch57L4s2fjeWYp6HAmYYFSa8jvQS9HXtrbHPGhJOFU
nMKIROwZCCqxZab5YRTbmlX7ZYjYykMM/poBFDIuwh8f1VwXtd0EBfBlYCkK
JYpjd/rm7aiEjp3gDmOOvA9b8MMQoNhgwi/IScFn4dQ5YrU6X0PPOx1l4zQ7
fF+SbZtLEM7tC6TQQhf/96rD+Kyj8PEnxJXsdnudM/RaoT1gav7Z1ofesW3K
wye3qQXXiKoiYsWGt8Inb+fiHg4xkWeAzpbOIDQF91D1rMJhnxDU4C9pkZQV
+QaOlZXRsoqjKkRR+XSw3nOqtWfC84cQWID8m/2w4nXET5G253yney0QBkhP
SbzI0HvuNt8kTPw/A+0DuIUY2yw0Reja5gilnPH9yuQvS39yunMbOwFoXUiW
wpQ/5JNg9ruvZSfrH21LfnQ/qSoLTn261O+CIGMctZo2RJXB1fhICKYjP8Zc
OVbWY9fm2z7D/5+jemVOWuKRctV6vKcvfh6gWKYG9pJmUGUYx8Vqh3JzvIBt
HQAoPtoKhOuFrXfYRljAdQIrNExFDYwJf8BjFP6SD9ibifhs3gxRyoclQsYk
5YBgJoqTG5ZK5DvH8yQvtwomuyR0cHPeRaogUkFb3olvDoi6LO24ONWo8nAO
EZYvvDvztWbw1rdGWwaltOxnf9Om0N7rA8+m8fp5Y1hDgnPcfHsRsyycodrm
4MdYAwMzugNPpV4WDwawEuPw5VL/bhXJIzEfGafYaheMTsS7MU+Eps3/7Kq/
qL3BYQyhP/NmYB2+BJBRW8/XRATk3T1TGmWwgTy2SrlMI+lSwczn30bz4y/U
QdxUuwsI44himXjph4YMNJgv1n706MRY/TAKzegPTa/n1UjoUlXoM7pCuR4F
YoyFBtXv/sEqv3XaaUqVFLDxjT7G62V4TrcWNU1CRWTCRyodKU+cnYi5slbr
20Gw6pI7lInsusQHSA8UhzjoSaKxGXP2qScVDaVJH8sUIbXOsSQyXQIxBHH0
kEiiAC6SVKAZaZw9BghJ07A8y8xEgJNfkAzIFYvSzJdUJ2+srVB7BTl4o6L6
o/sizAtPaMa87YinJuadocLJt+aA/aA5wE3P7WZv2HgMx0eSFXfo4MhxspRe
5Okmz/8Tk+C00P69rzaiTdoaFye7vmTcS42pWj35joHasO9u6T1yO66lcHQD
n4BLWkWjBlvm9OQu6hpzKM2bcbhgs9SiaJCnILzyr/d0m82baaXvK4bk2LEe
956hKuw7Uaf+2xvGc4ulkfZeZ8bjm5eEsZX6PBell43dOjwuitH2JilYSQJT
7+0dUk4h949ehEe3zoukbvfDUhTWZAYvyc5wS0QRyo08WJw3AUNNXieTCgCd
1cc9Kuo7dbTWSnghDquaDwsl/PMN3ooiPRZOPkWnBwRUXTFBXRHmm+p+jC8h
zpZ4Uyzp4RWHH1ZpZfL1alzIiEBAG0ETonNFk48F1612vHFUvYwHF5J8cxiv
9nNybMyve7w8iiu8TBfNtA0BziqsfgAciNshVQxqbG7oJtOBu98NmkcdpJ/4
9ErM56FKyIY1OzDoUvDojJo/Q2xhvjFoPOhBzEWhBlaiTQh6uc3/bMuDXhOK
T35VAs+FyMua6E0cZsh4XdqVKrBQVK7EgT1x23q2dQPMXnyCZdgfILknFAY8
oCKQ7SL61sEgsDCSVPqNKimWkooiH8SV/9LopefOMqEmTb5JsWjn/XnZTzxj
4NGkNJ2vGU5rsKDNGhZNaTDBGCtqYB02anfVFOJaq8PeGUhZo2UmOq3OFxJR
W6GF0h8waaBF8Cz5rG55PQyEhWO9mnLih87QnncqYvRd88MtmMbB74PLsvyz
2KPXB1QNPC42naoh/PvnHaJk0zk+1/iG0JvWqyeprj9FnanBHAzVXlALeIyC
xN+YtD5jfVuSoeAfUbnPV3g0q/hxXWsJDIGAdN4oQWQAgpBK/PgLeL8YdVP1
Za8fdcfWAzPoDdEf5neGE4mGkFiRDZk95EHZJQI99DAFbVOOVaC3GOpr4wEb
V1EY7/T/UGEFQfkioUqorKoMRpRCKPLFpOFQYSulWmMiqYlJHNIDX1kZVtG5
AeKy5sM+Frsl71yR1cUO7B15v0GcrMgGQgjuCczwIdzJ//je2gU8WYb5C1Hc
+iT4xyW6g/UPmKGrwPyPhCeDbyuc4K+/Gn9vW+6ukyLVxvchfFDuGFbWjnFi
n28Q6H05A9HdzYkMTQzyaWWlEYJL3VaHgLvxkbewujyyJ4bDf8n8Doe1Lo77
ixfHXCM03EfstHqxHCH6bt1qXYmle4bE1M7pONa5qN+YrhXUvfupUgR9/9v9
YhfdqQrf0s/pEL3vjZiElXaY97y6FVuZZ+NMDLfmct+mD/oYygSpIJrSSR1W
xco+A0KqDdi5tpVqydb8DsdwkWr+7zQ34KYgACIVm4bf2lqFL5BULBV+P7hU
flK/I32jp4LkAGVg7T1MyFcWHN4LYac+HaoGGek+uxR0fgaNAeStd3Nsn1AS
1pw1E32Tac5U4fUSNQ+/rzTEW/L18gvfzro3NtIvWjyWguyWoilVE91CWDMq
bxH9uZZBi03hXVuBdOYIY8kN1jICCFIkWU091x6t6dZoW3Yyp+6MV5bQj7nV
wzMTpLuR9c7xRYB1N3oKCLmQx9ldHETSmpYo+ByIdVJwDppMLEwbjsay+1zu
aTlxW4UIet3LcWEeh/jo/zEldloNzS77mHb+S8u8ywrq5nEw9QJaY3oL1CrA
wwWzASJbNOmVSC9WTODRlYErX64mB2+ykpi2i6fXnu8ZPwQTdAN8TVn1CdtE
LsXSREN7kKngGGrruiM0vxetpsn2NyUxTn7wl4Ln7/HoBsS3ktN5AidT5lrx
fBTjJ6YpyjOzvRLQ45YF7E0d/XQlYrZvgHTkH3hFx7ymwc0QMLuPmS5L0OEu
EJZW8H4leF9GVrJ5UgljEfwnO3hB2lcsdFvhw3GJ66/TwdDOKRcwTbagCNd+
w8TOGx3DH8n1QWLmcfyYVfBMF0foldS6GisffE9tWKNdyeke1QPnKpfdNXDy
LBAFL7pSSzV7zEtxQvKakZtmmuXuBr4iRIIysV1OVHR66JJ8+GGkIFll9pIq
dH/aw0vmxhnpjiGbXAOVOJgnpo3jRJ3WUxRwkTVmrEhLqRsH+wM5UC+kpvXI
bEUM6deeGlmq/cqs6acZFmZnZvGUQXhKgCK9UWEqIel4AaSNq42YOrev7OkM
hdRF0XZkgcPbzTZBsh1uCQSsvYe+xYT+UTiAtEbAfnxsjO0mkVBf8aoaNOC+
jlHs51v2g7f/7BqDddyZQwEjATIHlBeGVlvZZNMAKx3gs/ZWFNwiKp/YPaCI
8AeIGoQX67W9C0PanHfS3m9K/Ixi6ZwrbsNkgeErC9RnWEmVA6W3VClNBLxd
LegH90QityExeJdyuYqMzJO9j5M2/84svVdablEI2iAywZWRJhxQKYSZwsz9
fev5NmPabhS2NawHYPtnIXttwL8ZqYbd3zBKLK2Fvt8xI91vZKgFAuy9X8/z
tVzAi307FVMRqI60h0135l0qu8SFyUTvpiv1elNCwe0fH/1rcPXtsefgsgZ1
PBYmMynDmoZA1eK8qJ1GXEdZJjh0FbiYG+LdBCyRW8jDIYEScBZ1eaXOY6Hr
4cYnqj5/zyI86SoXl+xcrY6+aPERejy5tDm+gYS5XhM144RnL+Gv7CZW5/8d
lcC7VXD9pZo95zx40UEuxGtjfO4PWAW0FHlpqJOE7B7g3bvHG8fmj2iCCBkv
DYNeo8Ab35g0aiO/VuzX9K1FLk/Gg17ngLLDk7nD+bviibBNmwIuOlwGaA12
wCmsxyUfTkwHw6fhGcPFqc5A2YR+w+f6xnpqf8Xf5Bd2oRIQKzXKPTf1bMHO
Vbbej/KLiAStI5QqKuU9vSAq77RdTSvlqke+xyFu5aOKcHLF5M9pzxVW5sig
IKamw+vrpCkgfSeFjBFFKJdWgXd/yHgNEKsKrPlXlXcW1CDb9iy5rFw1CZpx
saUIJcV6YiwAjlCypApY6Sr/RK+84Kznn882UjBxi2W7PFbH3rTss6LL2iSF
kPNi+3IqdyQavfbpqEidyEalKPvdsL76pMJb0SqGW8ocKPGuEu0+bOUt5+TV
+IE3eT28RdxRLhoJZaiahRo00MULFyarHCZW4S4Q5lfcGow2wYaAD43hiT3I
M3dCN15fZW6I85d6bbD+TmyemiTYbqpR9R+wI2vS7dswvY3hCrNCYYv2WxiX
dKltU4Atm33Wrx/N5DpssM284/cdjS7v1zZ+58RGX9e3RQ5Zdmz72vAqQhrb
mJM2EssqTrk8ZpWRVE3U5KcpkgvlUThqvArmPTli0RfDAFzqLgEJ6hyCDiXV
/rESdh2TH/94Ryohkb4uqFVA95Y4zE/ciDErvClvVu5lStrkESxsjTknKSbk
AtckmGCZsrKMrMyozoivYSHAAMSZ8BHFVdXnwFiPNyIvgzKFB/2/1KUSPVuk
MGxH1DhPXeaaLuZEhNrJCDVq2SnWHdnQPlpTUW3fM00f6XL1TDEclmSC+HbA
ImCcGdFs4tc/dpxlBO8zRXj3mRC5A9MlWJbIXFod7aav1HOGgNLhHcBE5Ofm
QpYjnx3A0w4Bs8Z52D/fFsjnUz9iAjQTXptOjnsMfT86X6OgmCbPUvWk41SN
knMu2DBZrf9a7fnZDsG6p0Jd7TdbY5+zQxIFuPixSwYCqcu4NW2VERkagbHn
QUQSBJlo8QAy896zV6gLFSDsPirJRY6bwjC4Kirlt7yueTn0Yp7DQ2dBhNGD
YI6jH28Y8xVGCG9YR3gu6Esx41hFpZAP2uFHDptlytOPUZzNRSe/a0mtD3SU
e+K+9I1zRItwpscvrMs5oHZ+Pluy2Ar6EI1lQ441HYuFt3lzxFiUexaZ26Pm
GZ4jXbmUHO+eOC+YXhvHiGXN3ejQ5yxMEIHbPRHhNenHqL9JMuM4iYFUSx9z
44ud2BIrqQr5OP/8ak/6NLNfqanx4GEaVojOu0QB461/LKhTkte/CueOyn8Y
P9R1CBN1x7RH25+8pcSJsxTsEGtmg2P1zujLjHiPE5rvtPlE8Vc75AIk5W4s
s5rh5kg6MtVnYdeqqdAk2bJ+j21N18C8q4CQ6Wm8sDAp023bCjymJqzs5cKr
l6qp70YImsL4jZ17Z77mtjkDvDFlCw6ErXxyDxUhOx+nw5lkqHK6OGaJC4en
ExurmWEH7gTZk4jtv9hEr1FTg6Y2TAAABQJumwba4xn5hOrPtGvLQq1aMgYg
GoYIWdBZoIdeStROMN5c73cqUYAVUrmrvG2pR3YmO6VcpsucrfFuh5MB9Z7M
ZdqnWDaydJT3bQhbHm0ba6t+RWLCTlCFWxiuYxRF/Og2cKhc9qHaqDo4rU1v
xHTpAU1NkNEV0XG5ndvs1/6Rkan/GQwLJib2Ft6/WWrF2zI6MJKVrRqiB2oi
vzSLeNN+jzQZDaydnp9lgxWTtWZJt0gDWwOjSkvcdBO5r1VRZKYcDdF+gJ3V
0h+/DTJpfoS0BQvnLuB7vYi63rdBOKDAmxGztA2XaWm22tISp7dL9fFkbpgl
eyE2Upqz8LxG1OLUMByrF2V8Ozfnj2QioVgRrMwLzehI9wYrEmYN8gibgUd1
CpRRjYN6Tz3tlCizs4edFHXX+btYVqFO7Bpx74EO8cLJPFFeZ/PlRhbDd+Gk
qaG/gbmB552ufMxCkWrKo0yv2mV7imtHe4GXV/yuJdpYZmXM6PevoL50Fd+k
LDjB8qbWUGf6mhEfhUtpWPPnSxM1OVkQGuMrA1ij6dc29uhHSViYQhF+gxbL
gCq7JKxlX1ynrueOYluPPf3Ha3wceEj6cu56GFH+ePYIaGr9JuyqzhslHHuL
z2odKnRmqviDdigBEWJhz06QczMwFB61qe2d+E6L11Uz4eSf8RermWECZZFA
25CjseXtpP/LEdjzZza8ZETaZmB4tQL56eaI3DOuIOWmdtiKOKiJSNEIWcUp
c1TIJ7byBi5eJYjHGWbTAX4LRjajww5OPZvnBQf5X3RcnsAUjY0fXRpSbPqo
3yMZAzdfHSyT2++Hhc5qg8a6SBcD4wh11JFkInCVcNY22FlTwY1a1meYpR3O
D1/2QXlotFEKXUPS9gzX7wAZwwIhFjQ4vRE014+cHGYGa/WWT0izrTQnflbb
qfLvEJJYHA6vOqlEpNHEtKVy+b5YcBKmJu1LstOshPbdWehhuW6s7TnrhzfU
0F7xzqmQQpImZEiL+jLSPfyKCo4kuM/W+46+KX2hXsLuW1cCMKUfv9yF0ppO
E0NuvxwQ3i7da6RBUi8wa54mW98V0b0eWKqwbWn3ECTFLrnBtmB1uqdXG2Au
onwabc0yr6x4H1qJHPsfcvzQZ9hHVIW8qvaizdlM58otafJEcM8Ptsa9Vy2X
Kvlk9xIXxesSlVmEPWE1Fuplz7AMfEHYRLKfBpue2D7p8mMQ5d9lcxL4BduT
i0yk4RSJa6Wd8VVDg9PsjExXFT7okaCE7SBE3QCn53CWhkCzN56Q8vtNPX9i
8kJhTyBAE9PR5fQFyOclAWJ0b5OSJoOomnAxslV0mFidtSf2d2usjyOqmznO
F1m+4l4BJqlI2uIyD79CoCMelROnjB41oNdzhZpfGG6zgKQtfNST2HwC87Rm
ZQUZqXtathNOzRHn04QUM4+QhHjRDGvYVwsdJOUBjO8YMjFsWnJ5WWIejS++
ubH8WAMPApZZXOVZ1jrwEHVvcmHsPT3PEPXhQnCxALweivDCXnuhtN9qEqOs
JaI2fnF15mEQ9rfvJimsmvP4v/xCy5LgtdPF0DTLE09MKymiWBGbPktSScUo
+QwKK1ewBDTv+U52KdExNbqJI06snzaAKRvh03r6aoGXlQb07cQ5x8jexJPA
VqTYuxxlZD0mJDBvkTmD4qvrgZdwggt0kQ6EBWWk0e2cyPmw8FyBMk6zaXiJ
rBM3iK1x/kNix02lGS82T5cnP449jkGL36rGctAuZ/ydWyzzXw9/qswd8gVu
HtNvLU5mp5cLKyKzlUx7Pl7rI/Ta70n58LPVzRZZWxIcv01AGP/EaYRfSaQ0
zLfRRKjFMwDjd7sREYTULvtaCHkoAe1Jcg+uRMIDnFhyC0du/Dr7hMcpNEZn
uH2ZayNrg7DT6sntOnoQAkbCyW8fzVPVSTi3XH2/KGVnSqQji6DpkLKIBal7
ouMpSl7UosXFY5i82cgmRKaef4oCqd3MFx2lDruURo36qset3djvIOu0pIL2
GtT6QqJGFgTRSGfsWeGVRCcsn0T+DiRlTT5EUvqgIAqG13N5E827TwSCLvGr
nEJlu0gj9G/L7egYVihZGEIYCpV5RpcW1E8mBXkIWIkPkxwHCjq4Ia89EZJZ
+BNO6rXHX4hTp04OTqFa53zVwj159dDzdZ+MzH7tjFUXDqJsXR4Zlx/+OecY
p05D/R6hdaLWHoIy93a1CbRnomx54WznO7EQDCQ4pMsW0dfCjGlWnJ7HgAQr
ng9tZakGXB3ReodeFuq1RjVyuF8Q7FhEynYgdR/l3zQsxxItGtFpTjFU1C3L
87W4LeOLa9r5IBXntOE37s/RdjZj5TKvsjCYExhsjY+5wPyldsTnJJmC04u8
1xlcJSsS6orzSID5u9pbUpB3946OW7lUARM9SKogTleJVRrGqVkxb8IOcY9r
OCrkYkgg5dPbbbnAHfvobpnYnQozQasfQ7M/u8Y6Cc97SDK8Yp/AFUMK1ZGy
0UgvaR94QbheHAENsAVco/UCFUs5nwKY0sgOrOPPocLDX/OSGT8fEV+7sdca
Sk2hnNzLiOY66dKvATMGlU36uQlcpkc7sE0VBUrgZw7ja9K5Qmt6YHTbHtXm
3DLAwTR5/HBSU6CJaiY6c1dKeOK51lrGRpYpVGs/eWsTRcH6VPysKdpftjxN
HpQmIpeLC+cXWCsFwOCImMbRAwbwD+e827O869OXjAmhzVkAbo/ch2ajm5cA
A5roUpQ7MHYVedQp7y4CFdBstNhWNgcxgrgh7O00VMLjBFf00+sXXl2lg7b5
FRQ5XLE3xSGUEc0sQPKV/JazuPP5tLkXngVR28CuFW1Unh/COJqzmxK0FfiH
hAVvPuLrN4Oxljpsts/Q9D4JohV/xXPuloc4PtlLV5QmKKbAk7lVqDdRtByf
MytlX45xH/DsBD/nb3Vxqzrw/aDQw55+fD5Pqlu0geQfsk8e72ftrF1YUEyC
sHd3VKf0sZnZrhl2pxxHznUnCTXyU3u3aRc1X9SIiKSRbCC2vNcinOsVXLNp
rW6nfjgHcbnz14SJ9CXRHOqGUYkyHVSVXsei2m+2QVqadX3N4Q+bIIYmHMxP
WDkQnsIOe4J6nRFJdpZsLYzPXX0cRjDNCuJWPuU73XhhmzJP9QIJXgye7ckF
pQsNPcNaqg+LQceyhfmbg3DWEvzBIBJ1yRc5cNCHUD/eq48BgmjGnA0CXTTp
/Rx1aaHz2W7E5yKrPLTm0VotY0sq7LN9rI0H/TqoHrwacxS9uGP+USFz/wUP
Uo+b6FtfZvYzr32sY+MyX9s25+3vLxZIhed18CjCa8z3Beu7qrrHG12i+wmv
7/+V5lkfRrZwv6JHD36TN1kGHvNK72Xot7MTn8VtwRutPAFDpk9+3qv1awOt
AfFwVHSRNIrs9y/0yGciizNNltgmcRO5WlztdZjvKxIRk4x0BmGc8P5xtwB7
Os5NUR34uQWSteaDKWJhDizpYMnE5dhLrE1TMk12fW/VSC4tIHB3NjF/rKfD
0gvbOmozaeb8usr8q57MU4svDqKoV0nLv8qaeLKhTZ1u5Xmj8UeYUY9y9A1U
+RkVUc++lXkKhr4uZh5Pgb7SMhwTx+YPYiSx3eefnhSheBs0hO2HuJeXwCch
zXcSqSTq6TRowNHtQhh3Y2mV+vAyVeg0yCo15nfYjwu9aikyZL39UTKxEnbs
LOJZH1pTJzkk931sdF/+R9yBtSJILgFxKYIpEa/mmYDuVFfYCtzwCAXqWA0g
V16qJppkEMV3sHIMOkx26nPE6mPLfB0QG857yLy4pU8HLr7yyOt1ALOBc+At
lDcdSNzBODS/YYzsnrJwFdBfLKwguT5vfZywigKWRSDRNB15y9OVZC33PXcM
Jdg95biXShTDaJ6dbCqZKWvhHbHNk2Qom2X4oXXIQY22lYqvabhjPWbomEyC
C79h3oXuxBxJ5SZxEQqm0YrNt+ijTeTrjy2UO9Aziee4oemDFLTx78l8p3Oh
oYBNmXpHfVtZ1F6caToF1fS5aieUk9CrWI9nNmkZblcaz1K+gP+JGWtQabxd
caEByfG1Je+h62DQr7dUosIdX4603i/sQ0jhjASpRLweQSRGf6ouDJuKjWDW
eA+70NVD5ATfiAh8GLHHEQBV/Ezg/TRkqbVSSJpRy2SiMl/A0GFaSnEH+nAE
8vaScQF0e+gs9kPkg17qdv3z2zfF6ZotszPoVOMISWgo1QxabiW++jhSmdSd
eZAmOU7DkfCHfuWkkEnwptEHLG1oF2XHW4w3MIspOmU/Z71xOazeftOsWwV4
bnS4sZGuUXm6I4dxeRaG1wRjQV1UKhA+Iafck3ArWO4qSh8YVm/4sYzd4GzL
Ykxb4H/iKKfmTCKX9Yo08RAphvDZTaqNwgVFTP91Cyb2fzznY2aFVCpsJ1Tr
j7Pzpr/16SWfp/8qyggE6EwxMYh4L7oL2wlRKCg5LKk/AQ1HsudWb1i2MT8U
ZZNICBFFdN2dMWLvxDG6rWpk3jUz+g9fnXZ3qgaCAswjy5p7/OH3Km863Wm0
airevfvdc/QwscPHbTOExB5VvhvgNOAY9KrErmeVn1M/RmUh2ZvDlk3wD40D
R0ZS6dZ5FfbCjTfHYWy8o0GWtUP/lHQ9Hkff7CIAUnOtbuqSSjmAYvhepNXW
5DKEIQEQlK3W8Nw7TuvGrTyxBe48nVIrXMfLTo/lh/BVzk4ULHNoIzfbHPas
cKDsVPCfSMBPhmhwy5dsx8eHCXewVpgC/O6CoA+d2J2A8ZLKnrGtISGQKmno
MA0TxqkPu+5N1KnwsIBfta7el5RI5X23hbsN0oD6UZuJTxhg63QhTUjml7b+
TK0BC5VsvJmJ1o7eIKnfeC9i6gZR1Ge26Z3YrxYDUe6AgB8a07mMP0kzgJiT
ouVb0XkBtzsljK6MMR3omG9cw+4GDA0ABf7nIIGCikSHsNx9o93tY8vJTt9m
EQU5bAUlWrtJeLN+pRJTHJgjydLI2I2hHrNuyaYwkeb6uuKD307XtC/5ZNRg
saHOnWbCQTEVaNuLkhNAbyLUZqOW5+Fj5ZO5eCrFuamkVINvZlUVPA7b4BSK
SrwEwgWgB17Yae5TylyKadm/pnyuHj62QD5GEvsFlBFmqNQC0PCMn5efnfui
8sKBz4PSfXFoObzj48BdjJ+UsH8ApJfj72ygV6Gud7FAd5kai3+jtKIP7y+U
6BWXE4/DDh5CofZWxu6pIIXp2ToZh4IpQBCYsYSNQ/WNy4ad7HHwPO9SIYW2
I6YmGELY5EWq2WBiSkEvj0WyjD3eemhXiE+zdCaL5g56MgRcYBMbce4L43GW
i1lAHAzDBF+oJtsVMc7D6WIa+6tTM5Tvyb/r7n2Ykwa8tgBlhiSHS4SFHcUt
Us3s9dJH9pTdwMBEugRkQBWEpGkQkojGLyC3ZKIPxVXp4V1D8eLzUQ7Wv0ra
YsiD/F+G6uVA60RaINzG/MijnEnWNUVC0hZ6ov8twB0kiUedWSNrrLrdo1b3
n86ge1VjUuXvVjsmAJoPsPVcfijimU4G1hz0hrnjgORj94RDFXAhgst/i5qu
3tr9ble9XvMbqGDpxjVhtrUYJr9EdlAb0i8/K+IcVGcfBWobHKnJKT7bI0jF
/i3dibVHTVct1HPyC9i+i9SjWJTXzH/eFViHR9JaP44+qhyrTHWyTxdPkFCr
+J/DzO6IHukFRJfLQE+0NGMW/jmS7Hz3D8uuw9KsTDPbzZj4XO5H2wU4ucM5
qwDZv+fnx0sjOsiR4+HS415/1WOl9gvNpgUxOToyU7eN2dY8bGgb5HKJfviU
/7uWpBIpngxMKoIK/CTMqw7clKhVB9iGp733Qq5NkZcciLCrGU2Bla048by8
0NkLi7keI5KqvdNknt3wLCy7ZS7SF77mktCqBNYWlnGfZPH4mRHii9r49tML
GHI1VjzJwNg7AkADRYwRrRYdKq2nN+IH/ZRmYXIqiuzh+VjzE+++S3nO2SpR
5Od1leMDpfoR+PV5NJtdPLYZC4MgbdrT+IxkfADWjOCYesoVJl8N7SAVX71c
N/1BgflcuzlwQNoyMJh9ZvcsmXGkGmX/BoTCRQQxVKS16BakuXDNqxmRsM5F
F+pj3yikY6TXMcfmrh2wUq25xScHSqgDpYX9/1QnzR0PyoAc3xyxwAZokuhQ
2mNI0TX+iql4xrqa1ZEDZIIJPUyJ5h6lDEp23zzZRiLQ2mGmQMSXmVOqxz/m
RDFrX1NwLg4pPeRK1xqqdQUq0q2JoLYOv/FTumoMlgqvwq1sY72PUaexJAVk
srOFdvcjfUzSDvUayN9pvDSiGrZGgQNyGYlBFOiIwGzQkth8RC6TjbANBzhg
aUd4m74P9FCiF9nt9YYzMClChAXDbQcyLgMU+RzA7F46A/ZjnaoDDz1fsjZy
Mt/8fGICCxjA1pO2MkTZZQsAGAOIjoWmpQ23GG7nKC8agpkbyVqBgn988ZP+
FPUYhCT47O/+mFxeHL+rqM0Rk6l8bvFcqp/VZDQqYJ9xOIDQ4CiAoE38Zd+t
fd4zOOQy3fJPsG8g3FkQ0a+SrcAFFpLYi/M1RPCPDRbiCP7XXee0iTws3W69
G5mk0cry8jSpwwq5CZW4rOJ4wPmFvRUXCYYTosqI2zmUdTVZ/jNioO0mUvG2
Os9ofRVsySfXjEuI9DWUUls8Jt7ACMppssd2iOVvDfzM/phg6vCLnIVgk1Qk
+5EwghZRxo/ArhGqh12NvGfWuAttn+eWLqFJRIU6WDYTYzYgrfUMs744QKO8
Xs2oZazi7JRt8hTxnY4HisiglouDBcWRlpMt1+A9qUj2QczQyQGbXfLBStXD
zXt0hLtXuD4imghEC24US2pbTD8XCLvncYeeejdQrq5b3fTA//89XPuqQ71m
14k8m8ULuAoROSaXVTWaREKVKR5g7F+zqBy3h3tSxnKKFhDSdeeSaNcFLxVn
SDjGZsnUFTYmgypN0nW8FBLjDSY9Wvs4pfZZ256Bd904xW+ZlElHqyZVrw+M
dMuR2MOxoxGbC09hYzg2hhSXeKE8WO6/cp4Tw3F7qYcYKaFUvhk1ngAvMPB/
gUOGEjwWeQZ6lDhPTkR1Gs4/wxjP3CIJSjHQB1tcx+YkHTAQGrg4bbxgppfA
iXfEVer6xysvQZaJO5yMD73pSKy30rDoMX4vY5xHynIiCY+Og2DUxqtYeSB1
UKSqGPh29OwSwZOr7iDZUQWd0DVkk8alEM+MiBKD+m4RMauCaNmbMUImflK4
8CinFm4E7QtEHBvXCUcMtQJt0U635i87LEJwkXsNU/QeL2jR36okUXP4Wcgd
yk2g/wIMoVotsBQnYvMaF2neenaqFenj4QKYzFU1tZzoO79LnC/t7bNioqfo
n/etEdKyAtPf3a67EUy1PFsbWTCmSw0vlly7WiJLZe14AsRfa/Ombs7YXLkB
o4t25OnduqjegMuMjXIc1NzPC+jGINu1MjCD9u4Da0dXprVoYbeZxGzRzyzO
lzzu2guOslMeWpn3G2yYJu5ccmHAhi+V4bQjuJpZByxD9TfoWO0tN8yH64SL
+1cHbkv9e11PuC4je6la23dsEtkR5HSgx0rZNDPH8+KIrRYOxeHUlLoYT37t
IUOvyDXy3/U8Wmq7X9ufGdiNOxop/3kP5N7+XhXQb12upLFRQjhWC+ags90Y
dZhPpSjnzd3zYQrmtHZNyyY7jwRERc5uJRFgGytdyIhdL34nWaGrQLKVsL4M
IW6j6oBheNx6SxdKRPa3ewN7OGIROS6Zu9oDOj1QLlZtdzbx0ZYT0JCjCOz8
kCEIbZxp23qXc4288BNKkhD/g0weeqgsiwtll7+rZ4Ih/rjXINWIegdRD9Zx
CKbEAcrdNjSYHu/DnY2lMEbYJzJKlvZ9/alqSolnkryfr/GLWWW3NlTKD20u
vVb+UEpdlWDDp4lJwgbZLdvRswGeRvxJNuv156cWeOlBcXCOlU0dne88S6Dz
rfUvk8/ynq42F3L1W0suZhsfMDdVP2oG+kDfUDMzaQ55NMImnOoIcDhiUSGn
k0YAE4CChKgoJng1xSBeJyWimcvAGRQMNV1pUti3FlVdl7Ltsnc1jSJ6b5gQ
qH6NLHV4ycsn30TLAjKucCT4FR3T4kDNU2m8QaXmLKeA/4BCUsnVEED7tb9P
X2s7Db53riqdPrBewuRCYpAK8qxP162+TIiJpmMIIL4VSV1p4FZlb3FesQa9
/weZZIG+QrYLm+fJ+CmCk+7UcN2TK0UqA4YcJ4E1Xvl2aKeH0kpO26u9SZ9G
cOMIjT6rBo+JL2F2qFJEBpx/kle/QTzacNHlEfAsTmpBLlQyMqZ9KdDK79lS
b6AFyjqw/AmVBqU84t2CoH3XB1vc9fPpCwGAK6JL3RVDs3YUeKumjLBHSv59
LIOxn/l6pNVAPzDeLQZyZmZEwgqPZniSr01DAm7HdYc8lXdTnNBYtBdndFQ9
4raF/NC28xJSLgepG1xcM6zsOpsv76xnHRFLZdz3gInOGV/aS4cCktZgCTix
wYeq7N3yV38eCGBcLvwSCRhkQADTN+X8fSZuxbXoZB56YoUvTUaelFMiQdqB
kIhVP5cUyJcC99FrJLuWTS99iD6mzbC1ODVJ1plMbSBuz3uKM4/kdKwn4ILR
BEHLVwB9e2IzvY8I8cPAUjBkgJHOo/SGvaefW9T6DXX7yHrFjfRnqwIkq7wv
O9T45jr7PydbmIZhxZ7lzLuyTLf7/mxqKqBX9o76+W0FW0r0WNCeJBr9sbFg
mdshevq6JaMZORR2gq1ZFWhMkW3oeRGU6TNpjeCBn9S3VHpp681VpMnm8jDI
mFwpi61bs9Ko4NiCvX0SZWblg4iaOEvoC9fBO691eiASaE1I30eZ/AjlS9KB
/fbmsVWHF7/tMp+Z3ZKnngVt7HRwDh2AI8Z6phX4iArKQeAoqGDM8F+1AXab
P3J40dRLjNQhoCpZhuT2tMrQGp14k4dY2AZRiB34Ch7LI+6Mcp2ZmkYYcsWs
aDppQNiP+arY0wdqD34EOG8BkAkjbKUgIWQk3TtXSh0fw/T82tsJ5RYCEVg/
eRjyv8XU+/OxvgYUKqSGVuMADqo+QNkEPxfzFih3bDyfJk1AG/vMr9jogYmj
YzcAfSZg2GXiuj/bbGRDb0cCytETwdeOPtDs/YMwoL7Pxx0nDSFsvq9eKAN7
ACn8F0/7xRGV0OVpbjoY8Ji1KvzmYjssgjxwrBxATRdtY+Gw60j++yu5jxxx
Xr9Z1uJGVJqkVcyYZz1f6/4jgYsm8LmSHTcWe65McZG9QtPqEO2spvNV03W/
BhRpmXyb4nMW/aJDpNc/42s4W9UhHWmTU0vwLfCe+d3PsFrATF/iYWVhE7a0
je5fq6jVtrJRpKNUF77531Xfo5yJ2XNO24ScTq4KCm7W/d0U+qfC7pldbqbl
TutJPN09D6OtRJ4YbVON16RzIaqOXQiXtGyrRGDypxwUIBazYCz+j3YFbmiq
dUiA5UjEnSkLqLIlkHfoimVEqD9ksJJXcsdKdpm1Pn12WDZ5lPku43jOc7IN
yuSyL8UL/JLmYXMyHDeZP33VLTfCNeeTiqS5NqC/AgpoqB2tW6SM2P3vqNeQ
6b6rF/JaT1dySd2cLGvliB2FEkD0piorkJYhptUApNfG+qjEZ3ZgkMTKMNXa
uomTQRz+yylHTz4LQbUcOkKHjHEP4ep8Tb8us1EBtoT13J+O2bxSJbRoRmKi
4rd/0IDTXUzIrd0NTl4CTj1RGYTb2mPUjTU8rSxVulZfhiCepq19TKsMZO5g
uu3mP8ButdWd4S7BVkXBD8YmvsIoa6ONfXFFvhUiGpSRaKmb5F/Fu5n0eHEX
RH4HkjxEBfvMKKadZwIyOXkIL61tPpmfmCCKzTuuHvHftC2w2t742X9XTz54
l8oWpHuMZYF1MfRreoGoXlgWuj8hHPG+UbfOfTHCAOwon+B8BeBAIP9t2h//
kxwDLrhuCs0ievF0G8kWZ0VXBMtLj+ZFZMoGGN3kiLIxnKSrtWtzhwFaTfpC
pjH+zsDU2kOKYxdJ3/43mhf4z5UP1K4JaE+DCPDkOGrnCZLlh0k91jhV+M8P
DzvpyvzO1tBoWwDkOzfWzBTj5eumYZIZfGY/B2S/mf6AWUQ+HebfBaP/x8JW
ttnOvWwm8YB+G+HEcPDqqxu1WCEZ5CFOw0bLC0N13weZWHeRGlOXjERyIdII
OMQLt9yx2QY1KpljEgjHKTr3RLNt5jAB/p05WnypbVCNPwnn5z4ttbu67ldw
3RTOfpRbYopQfzf9/wdTm9vyehdfX4EnCTzXpsh1s5f9nl8dM8zUU9g8VmJd
KSmjIJhq09H+AB25oNNjEbiWgJmG62K2dZbVOi3l43s8UQTvC7NrYcG3JItV
5UxIS15qGoGhrzLpRYQesHgGYh94xuvmkMoxVRQFkdHZs/kgv1J99wH7N1UB
RQGM/Mv6ZBP1FDHUtwI7qT5gqF7TFGngW7ISzCdI+mgPeaR4/mN0xyTGA/Km
KGJbYTSQqD4AYCCJCDqYHmwBn0YtemsrRZHu8tgZmMJjwaSM/tMWRbRrBWDZ
IHBsimm+ig6jXdbRp5TplS5vRcc5iWWzWbS8iTwn3bOZNEEUaat0x7kBP+At
5zhRhiDLBzPwuHlG33p/qUrdARK7of35/lsgh+jLUDG9BapOTXV9q9NSPJbo
DvWubC9dQNjLO8TFG6qAFTHH1njKe+Qmez/j/IO991QqLINxtr3FLaCryFEm
2XEZPTMU06VuqR42mjvZ3kJFUKdiSEvRMvOGmc3sjFAOU26H+3AQOOQVP1rB
2tpCgFda8O/yrOVg4rnncw0nPfKxOKWcPZwfA4xy7u5w8Nymta3tucZ21+On
FeS2b8Yrenu9N47c9t7dJEr+A8RaRgnkjg/DJKLpDGUP5bINAVAn9lwx0DVR
ek4zl9bGZ+bBHZS38U3vbCEhzb3OZbUlqhMaOam5/PSPqYsAQw8OJX+w3Ayw
iiHGE/lNPjNUWEpAQJtReivriXqZNcYAnf0wDXrg+1e3N9lz6UbTU3K35hzb
qvfME1BOqdFwR3vtbl3/1yQyAnybJzD/WSENM4LAdA+7UckLcxgZyd7WuczK
zOW6mj/2BHDnu6Ba0YPfAH/K42ay/o+ipq6FbLCjOhyrTSF0XwDoTqMGVu6d
Kq0Bm+pdneQZ4Zn7s7Bf+cuXs53u3ea7DD5Ad+I3Qtmx78dBAxTge/svlC1e
D5itR3tFF7TKAq8ideDDcJ4DlXNDctMsyiqPVjKXDgWPasEj/ZTF/ptRyJrQ
hRkL1ny6NQMzGefp+pxLhmINc78JjBFuPR5db/bbLhGNWQE5nXDA5D4mioi1
S6oolhtcHV7RObvZraTSF2pTZJXTWwTdGLiYbbC6lp5eLbGgZ6i9vVO1kiv0
BTXMoleZ0UdYIvJKcv3gyMuHY7Yc6ypywyulIk4zzG2+pUHumiUQ9fj6Tamz
ZS/NINPxcGjVp6nuDMwqyYJx31wB5GwCaS46E1CFg7eojylMw2o8377kF7qf
V2+OsKLqwjwksVMIBAPu/m6bZP/3/QOVgcLsrZpXf6Zrmr5ndwA0zWal2/cF
ypxmVN/ZMLzcjD6ZsxsQvUNO2n4bcWvx72QVAbJZsMnt4ZsK6a0hXGfh7dO5
xhjv+veLVphqutJokFMe8ajtS0WgXg7zhSEOpvWNyDA8lUqKRFi6i1jzUqeF
gU1+aDHcNEVuIEKgoXDCnYTJs1/6wz6iXb5J7intgYnYYoTvWCz30J/y9fWy
ocQuhYKv90XvxoroDLCgqwSGKUPbTUlULOAkAaYIQjk/gCR2rMhslOEVDyOb
qDAFNUr+5OY4YHE76+YzdnyurI9XrGze8bO5VhCbzBtpYHaD1HR1RfaeXeVD
6eN+HI0sJMnWObRDKk5/09nwUZ5lcU8MWLbNBciFGvzAVcKUl07UFQDZOJXk
xxO8lrCzpu2/WsCWC/3q+fCIQrbaV6m74G3mO9D4C5gLbQoc0GgJuV8+kw6p
d2fcer4G88+dK9+M/FkjxwuJ6tkrufJDGCqCZNaHhfCh3KaeXFHGGxEccvgy
1rIlXnKP8cy4c4aQiK5m3R5HEyTLSSEqXS6Z7UmdmHrZYTznffECHu4QHBVI
b6euPARe6OnU76BrF7J+62F/ZkqJC9hkZRDbjMj8OPixNTDjBvxTZtfy65iX
juW4zAkqBNpD+0Nb21TiUfLEdh8Y1FHfdvAD39r6rogZ51nDSimpHnteMfTM
ISVFBhD4k5LUrmUL35arD1MGDpYnEJPXBrxhe6Hu49T+kiPYQJMbF3UusXuE
a6g3I5O04v3p85rduFu8gIV4VAer0jvrZLbhQDu8UcIuTVF6v89t8MbpnQhX
8Z599Wu+tvff1YMIOtKA8UsCe4QP1G55bwUrKCj6+hFcUjPyS1Pei0MFiee8
M4iYn5B7rIgMh8RvtwpxNhQaojzYDeu8dtLbkJpN4eQ4TmI0lNzvhfn9BClU
MEUYzzqtaV1TtDJzu19Cwqu+kJeDSB1pLnGSQNv79Jzul8HsbzhD2MP/nofk
d94rX1mYl4vTAAnR9HrsqF+Kb/PV8FxL+9reWwIiIfmnkllx13Ild8BrCx4W
7x8Q+aDYrTy3chRDKgMRfULOdeCBV1F7Jp5xj0Iv+0dxcdWwoceUw9s2yi2I
H7oQegKyqaIdDfRmEMSVvlhhu/X3E9VP/oEe8ZsJx9JhwYxglG/jDRWChDw/
LaTTxshKJZVrTMpRUlOy0zBoMGJjpXf8dN2KZqkitYtcqEyXHIj/aD2wp5C1
+pZ+WOIEa9G6tIsERQAEQK/4cVfrUNyN3WWqGq/T8DgtQzPkBka8yqnAb5IK
MB1j6h9Od4mktCobRiDReuQm52NhVENrTegfNdd2ZX2SA9jE9Tv0tCwoEj5a
LAQqVQi7HNg0kgzHCQ1Sjg0qJY4Kqw4bWfxv2hChYngJtLyq9ULPRyQ0jzPN
xbD7VDQNwB8NAfFNatSZ6Z+BdRX7NsIGHZ16/oliJzQMhICuzyF7n9/nl/EX
bXi1uoe2HFAXEeI7OltQ5Mg5K4NFMaxNxcPX9dK4x2T+Cat2bG5VReoDkX71
WvtxhU8TUbKlwuIYRhHs+yv6W0FE1kHH79Nzf1z7TBN3XxH1pM3+0XwbhtjZ
xCSho780KeBTULuKgdujhFj+/CLizAdmGlYaw8ex4y7MyQsSrixAM2w1xJu8
qDqOBU9QGN3YeJmIF4I8q9DAPHmtk4SEE0FFO5FvIfguphHoNA6n4p9DfxEU
FCxv+IShr7o1AcIbGJ3igXYun47rjfV8YEmJc0ajumjb290FXhYsFJvTGhdD
tELSjQJ4qIU5SizPp/JbKCvEtUl8+lDvr28gL5XR3BIbcvqJBE6S2mT6gBPr
uNjTB4BMfXrJKPqBKH0/RoLoeqPtxZsQNymzGvin20xWL7Cm3B0aXDx9yZud
OcSYBwtEXgmqsN3waj5gryYvrZfFDyGrWORViYnMC57zjayPALbDrm/ZwH9b
+Y18kK4jJ8BcMmjxRbUWrAygDwzaCeBgqgikxd7ihu2gWZtLRkwPw8BwKTWS
ImD0For603FxTSuOmzPD1sXFPO1V42WR4vHzT5f1ORSy2dd/4fAy4vWffwSv
M8FIbEiYz6uMDe+wKOVtcnPWYpUJWC2TL26ubV11TSDX9q7YmchpZuQj/17n
6cTctffBkgN5bM6dguCWlpWnhD0GkWuTwaTnvy5tYisHlb/Fs22Nfq9IrN6O
Lip9dxBPxjGOPUt9IqhWTByjVzBcSxg4YcjqxDORggINEnc3UxtC9b9NFTMQ
1kCbgn01yxatC/dV7ZPIk0GAqVIwBObGedBbCxF93nSl7mcszfLHmp1NhISm
XsZS8KAw15Zckf4y9JDasWCrq6b9dOZMgoC896fEnqJeHGoVcy7Q6BKUsJZ9
4nLqltvekz2EKSV5U3x9/j6xhlyuz03wqtBvU+IjZrReJYdHKUIKTVv8QoDh
uO4t/VgJbTRhHEnvsVR8PgUsFekrf7k1xNYJBNho/Z1y6r3OkLDLOg594eyi
uf9tQtRyLxRok4LZOwYvD9996OKjAbF2s0CNjBu+jqrYr4Flw+mrWjHOadxg
My06RSphkUy5hXwnmJ5MCbCZ/UQtGNroHVEOW6W4Exb8owNX/rH5nMuhRdyB
ERxsL8Qt0lzH/TAudSKeiGfhwJMFZSxs/wDX4H+vQ4Yo3ZrteVg/yAcH+MdI
8g2CPktvGyjJzli8Wx7lkdWBEMRQjuh9tlCBwAXObtuk3nmjevEL1Vd98HqW
Utf6F9N1CkMqqUA9LAzGWFSW2THCy69DbR0KmWkWoL3xNnU0o4mOjaXrHxTg
yPv8QSKilUKg5LjsAyY5qlH7p6InAeA6J1+3+WNF2fpDUMkiP3N73aoVOah1
CCPHy++rj0qbPvY25X8afEUxXpcrHCADBvCsmO53mRXuvUS4EtD/tMfe8WFP
l+Ez4iBgNchWWvkzBryNukIXAIveR/KuGrCQyi8L5q+bMl/mxAZWBYwxUjMh
hoKNj0TjZwzbTpMhvP9hy0eWwC46/jwMpiA8TnOxbiwO2mfVqI3ZD8TpkHLj
ppn1yxFbr5FHzh+CTicTw+uqM4aDRth7sYYBTuABBFZnezOjcxdLMKdeQxr6
9/s4y//0phMl9yRinWGF7vBjE3087YMD+IbEDYfBYq2CITokecKP7xAijFh3
jifTfRdWiFMZnnaxGZV2ZiKAwK4pE8/0hXZ+0peqgTgtWItIsVv0CkIt4jaN
HuOCgmy89K6ua+GLEX32MkpiuVxOmyhSdtyB1KhZQ+yikku0LQ0stVH4j3+7
ul5IUJQRSgWPqPRl5lc5FuBboTe7OY5loNwqd8lmFyb9aJYIkCdR7WS9Mwhw
e0YGQzTbll6RXSdCD3PVSEDum+canmODq8KTAGqFCjEYKMA4+REdiQFpbEUL
j7SF3cm+aZh2sRBgICWcBgkVDIcJH1UPj19JO6171azZwfQV+G1J1oKLqHuH
zAsKvu5MMH7ZPY9iKaoorg+XKXr7Ihx/XX/LT6nBkHTawEVxqNkI7SRuL7Dk
SK9+tIPSpcLP/NkQguX4SYq4yDhiWhTJaDurM2suwWhFIb0gszJlaspUppC+
wNhg41Mo3hkK3BA9NTNteJmWobQB76l1WcThg/lx+wjviC0TxXkwlOEPFSfP
qnVUJhWz8D3TKAskOD6fWXdCUkjjhJlaogfY9TAL4hzPQzXubL1BnduHZ1tu
3NUCPhSHsX9yXDvGA+Rkun2JEV5QCBoDm5WUwzC/14nUGKo1S2M7gxef1FOv
tcOLXWtwtIzdbS8QC9oKAQ2AcBcHoinvElHO9lHoKH8v7JnxgiCWUANYxOWD
t77iosGNrXEA4TcD+ICUDz7EusOG998zDq0MTKCK2XyUKETm3Yua9WTgZocH
8GClyVBYtQnwzzQei5C29BEMVIQHmkSEU0T2AfHTVrd0ZiQXcciMb0+GZGXV
OYKKA1FJofAwpKjHrk4LjjzaYGZ16Ys44nOinlHFeAEXXx//EKcTDrLmrr70
9YG7/mDUbiPhKFku+6z7xpkucZoODsT5v47PpPWtAyXmNK+DFYGlVVYnqyfo
Ca8eC2nvGyF7WOGrVSDaN7g9xGw8pCBMajAb1r6Kzi1II8qcTGTVtWkIoKM7
GxeAffTpt8Twtg6kAse/b4iX2/xmq8s0YkjRVCTdSYmuHtFM+p/kr2gRN0jw
QhiskOXxjGxUhWgoNs3caWtbkjW/ZUckGFlbpvrluKR/cwV2o89jvPUOWpPC
ad7PlWYFH35qHJJrlKc5dO67G60YuYCYFcjixWWYMq3KxyGt4Sjkpq9Wemp4
/78tvFknGVigVlpvassyZWIp+r0dXgz8g3xDsHbCw5Y8SRCDQ8oQffPTo59G
9V/8DwJvgiTPYIr2IpB2DuQwPkh8vS/GTGUzJSA5QyXM7+e8apx6MjT7HM7j
R1Cbv0FQPMOZSt+6c75puK96BRh1n0c4n26YCh+5OIrXW+C6LcqmWaqKgSZ1
/ll3snXwj4dGX9mKiBMwXjyrawQXJT0EwNpfCksQGsxUD0Ru0lqBpRP5mBV5
P/YwJKA5aSCEAhLM/5qHzpCkBNiTQg/uLKzLc3mrbvaOYZMtQnjifMadQOw5
BPAfVtPNmfxjJ6XKl7SCu55lOwXlTi5Busmh0vXphimoBOcR/oozb6aGy2E0
u6x5HmR9TkiRs35wEkbU2cgOfLRvTa/5j+rQwaknRYbIB6BcdmjbyHds/VGj
9Zazv2+RVxj4FtZk8P4IH0u0BgZSmOIlQhm/f+xqE4zirwm2yBbn9L5AiQzv
QajryRFLYH3I0rh2lPqfN8wHiApfmJ+Kcid87JKeraGkkfuch/plonz59oZA
euxyTUbVQ5JqJnFcf6L4QtBWArGZ8M9cxZCy/c5XyvzYs7bpwRSBcNymRsUI
tZrnDUrT80eMFd4g+bIbBBtGXNuhdK6HkciElzXO8KXiVoS2pF2l6vG4zrsK
mcObmJfk8BrYn+s9rSAS1RjhFt5vIJ9hU/aiBxUWRJwpTFA1HOcnr3OFPu2y
GM9HFOuer6DeLFCAjcA02AWoJkaAcx7AXbRHcwZ+GNZcOidfefP0J08zy4Qr
jmgpSXRSRE0zyxD6RnRIfOI7Jmg6AiUZtrCFduNGPoiWqF6tpr3uXNdcbz90
CZ3OetW1kE32nS+6C+qqsRnS+VtZuU9eS2ttwP4ssHRHZ0T3e6ISy7qKh97m
ljbRPV/hJHqt8SzTyemaYVLaZ0NZff/1fd01Y+synY6gAXoqTiBkXPYXbb34
ZXEybqdoAAAQ3xCoxZpg1EIyMppbNWrb6FQsNjwObzQw5YN5ybXs8kgUxeY6
voxn6+EpGCYWUqhrL+Lc7jMrrIBLLb7mPWr/NNU4BjASAmj/3m8vBlewUob9
jmPUqQikIqtd8xfOLqT6dXgJBGtY/sB4BQpWytda9MnyTzMYu9cHlamz4y5o
dsMF974TY6AsLUIUE/9rxD/5HzNOqQyYwFgjnwM5RcsjzrdQ5C3PQx/lxYLy
B0Zp6/pY0FycYiZoWaU4C3PmzTMIRypBY0dujoTNwKyS0uBzIlYykb4tU+AJ
yWLuy4ZiJg5Z4xgCxDiL6G+kPRp2uwQxudRAOu9Z3hufQitdrVPSjMorBh/8
t4PBVQ7h4af+ra2S+6G0LpLkJWOHqMFIJkRYGqPAWAjH/kOUcyh9ytkXb9hj
jDvyKLWYTpewjMkzSocZkyntuOYqluZVTa82knVc8jj5lGiMxsohkjWSDffj
tikROVoZpCf258LZ70h0nB24ykXqWGO6Kz+2WBISp04So94th2PTv1/efUj2
t/Dt5xPJUZYr52O+5oz1dgdSZbFQfj3XWDb8We6ngmfASapdoqPWVuksmM4/
Y1q0Jb2RNbXVpX8AXA0mY4o8pknaSBxV/rOoKuzogeB1gTeW/6/mY3kooc9v
j0Dq9t3cf0Od8HTD33i/9EUPCOQIIfSncyGTHmO3nmGT6ddDqrlpNFLN0u77
vmq/cZVpIjSpEhWZSnYp/7+EPbl2wj2lBcpaQNJlJzjNr86tB/5ZhgUDkAnp
JGZixHcuYandsoN4Yu31WpiPEj7t0hgovR1ih3BbIOmHKkPnEB3/yBVv0D04
aH1zf8B4ngFa/wTeAqaMLIoEfkj7PnS0CZr/cQPQSc9rfMmUFiqj0WpnUtAi
0DuDm/1detBzqiQbn7bNmBZw/MRFfePAV+HRfrU35TJMwKQkjRjuDTl66IBJ
hqgiZ/55LyWq9Sn6cwKVghm0k2acUYQNEOIICjJa2lSAXQFH6daNFFUFS8Qw
5Skqi/zSqRhH2eUxSYNnmU7HKQvLq6okzZTVUoYnbpbO4GZv/E1T6f0fY3h2
8bzuqYERaljjT2IMUyXD3w+cW04pDu9FPvFXIZ1QaARuozQTuJjOR/V9+lxD
QmvKl3SlpVKB0mj0WRyhQZWbrzSj07u8dhoTblZC9EXYl3fMNCP3mlBhD2PQ
hKaeb5CFMk6jIkVrqXbnQpAkM9a5xy4gby3VaOROoZKg6Brxsnw1suxGL2iL
Ec/69geaqowfoZoIUhoQ6I7K/rHJBwSo/19pWihAHLONVwbWJGtx8Eplmvsw
gWiEf43zfNK5mk0QtdzU6WTdWbO2hBIHFzKlKtPg6FZWyVNfE6QCVEhASJwG
Ax2q/ocYED6JHWEzFuiBe49dXyvMK5p+SCGUqyG41Q2rQjQBcHsXYIsZxFjl
yZU77leH4PKjrBDdxH98KMMm9dSXa0lhbuCsPN0j3pdQlXgeYT17RT4Oh+mk
HBeqBoF75zns/1eSLkkq0xy9AlJoS1uTBPS1EfHEHiPOHMxNSkvSj0/qHMgF
BFmEuOshGGihytDIGVKXIDKm3liY1hrnvm0zk6CzxEeDlz6gmmJw3U6QlJTt
CBny9jpleP2n+tAxIgnTNOEtUjessk7CXdLYel9IqEh8SR2dwWtPN+QExGwR
Gsz/dqhagIDFr2NO793qo8KpD2c1IR2MXbtugtaIv5Jhi5eCVVFtwIb+JG3q
blI4yb3MAymyvGD/na/87qaYUYGCY0i8zrbwFsk4Os2hv+oY0Q8jgPFUByWc
edNJgdYhieHVyOX1aJiopoHoXMyb8yMD5ZW4EZpflToyAv+8f1ZnMxxX1NoE
Bp5Pr/4ei8nHigkopbOJMlHar4MZw2ugjP6huCbFaI4Vy1JHuq6t5GIfoFdi
GwRfK6tu9J13FG6fAMV/v0mGD2NESTGVNg1DE02OtRU269TX6N6bNq4E8o3Z
LBuwNVW0u2isJHxmag6LKTEDgKuYC647Zn3rAcZyPeSajh7IQkpP/RipA4Fs
uOV0COMf+Qz0kpyhapMsIIho+EGF3smA0rChJ8p0iu1AncH1B8qreQEnuJGy
tyTN2bTZXFDv6MdZ+DRTtR1Zm4EUGj2kWswJ/hNo5FWVLnax8mEvEDAcz5Wv
/LUrDkmSNSTRMnqRno2ZgoKEnALmjPtJyoAeHv35Gj9bqHh2h3iOV0Gym+5k
xP7x+y2bl2I72znK+KEqBKBpLYzByuSkkIa85A518bDT/4IsHCIiboDQGTtC
egdZKZUWGuC/hAXpGd/cqRLuGqGfPGNsHfUrYw033Wd9HAOgybZwSffEPxS3
+4QVmMuc7qK4/RsWtPonpdEIcWEn/v+v23a3381ZUCK1PUatAYY64aW5LeE2
yxjv1xfGXUI3GN538ZT6SXux44oRdjoBnaQeiBzS6i0DchfxGfH/hfmY5b5n
+T3Mw3BBv2FD82aPOK2oQZFYJSNmEInMkam9nsFGCUflPiHKEQYD32Kxap8v
3joqQCL6IKvYBTzHTjte90CNJznOgLJ+q4l3vEYJECzJVCkVOK5dmyd65a+M
qTgkMHreWK6rKA8e8bl85L4hSeY4Gcg/kNveyXFQ6b5JhFFpNKCd1frTy1ir
VyXilZ0l7AFpbakA7ZFpmWmmOQATCK1o8QQ6lFy7jyCuOSuvxLCLqslWPJcM
PJtqb1Rq997/yimNazCK+PIHjGH5feSLsTzpdCiDPkt/2hHRZpt4SrJY+crd
ItI28GVWeojG1OJs7joTPRrVhN0pLtxd09LnUH7SnucgOoTiH4hoj2W5Lvnb
vrwKodn/iGu+NQXuM7UbweWSBOc399xmqKQl4VmGoaLVaeQX38JbwHn9hYF0
k9KbndUFKNZNt0BlEJqEO/vcYrL8dCfW/+96JxJUnduWdD/XQcoMNic1zsJ7
VDrB/AV4izMMU8k3onarZ4Z0sjpdB8qlZcJEtvx19mYvQtYFn2IV96qfdb1a
RUUZwcLWOamReO9QqCZhjs4GF8Fz3Vq1FaqTWX1IqlBzOCJ1TgV39VJGm+Uu
0W2brP8lhE7ffh9DrtC4N3+lBO77BECs6Dhne7ouzUKYcumCaIghfBJkGqEf
ApXfZOTKUk7fPTccb1TS00fUDxlrOnExJOtpmzCTnx31jPY746PAt0sSxAF3
sh+fXiuQLa5i5pOFv+Ld8tz+P+PoKS6sM1aOAodlU7ODWWqg0IRYBatvpC/h
Zv+TDTDwQZcqP+2poiqK9hKjiTyViKCA+powbQAMYtOhbv+GYaugP549QGMG
fHJmHWnjv/8BV4Oz5dNBL+SD5/0ID6SCLJdiDfNFFpHvmPqQ1s/DXZ92C78x
iITwmOgfoleSXJF4Kh5Gfk71nLRQ7en8V/UU53FDtJpAlpUbRURmkaZZl6re
w+D8OJH20bxU9P2awnP9MYQmpdBKsE25T7pwhIjO31PuN4U4pydRYgOrq/I4
S+pUCgykmcTaKUHuFU2vNQSM5zJKpB7I+j73rqIOXR9gFnZXlF9aWF8EeBf5
g5pxUkER+ygh5nhJq1tmUdkGJaQpVaroMqn0CHYySmVfrCM+bqJGQfq/hek+
CbLVeShJZQQwXu+mHOJF6ZgX4JqYK/2pOTCDRz5aes48JzMf4W4zVhBSqUNj
E/LKxmxOJENMQ/qtvGcxiBP1STeT8ESGvpojXB3bOrzP1RVaECv+iJOb1OW7
f7rOi5c9fnW76yDviNSoiqernRwNtPirDPbCArdj2dUuioF39zjwtqIRyxet
6Gsdz8LNEIl/upRHrsScGkBulseW6QKmbwOFflS89FSZnw0P+7yl7iPhruL8
xcrkvkudEKWxiM3KlJtE2hlNGRs4UiSBENVn4AdirZ6LlRPRC3QfHl2LREjY
1QykERjETQtT+Mn8d7zNszYh8eh3GwC0YFqWmsyvLj8+tb/zFSq1dVEnY9Vw
CkPdmzayPNcxibDaC/Ght8u6nRcmMYA5w/wh4pjecQHZqjp9uv/66sDQ7VOJ
W82hfqHFtQKec779Rj65a5tCPHd79PAm5VyjbHCpsRRxRvRLpxrgFsP0Jd7N
wQ6l0I8un0ItYSJribTiN2Kw9JWfk6WRIelnUtwFtLfHzB1ELcVsA1BVvHnD
i1ksD9Y6wC4at8I3ybzkeMPknbOU+WnJeaO5dqaewJTZaEQc8a/dF4K8ci9H
0w+DFcb1e9CDGyfpsfBFh43p/8VGNxH4cbpOflUwLajalXTwyLiuTy2U24KJ
kCT3u4nO7RND18pd6BKBZzV4XpQt15xtbhsfV10AlTdrv/fQjflJ23R5ykVs
7pEYbcoh5GCXWm9wFpb9kgfQDav70OhQyS43i9TvmoxQPzyDmH7oF4e2UXIX
CGKKuUTextjv32mYSe3B9ao2DgzlzmLsRnuXGzYAWDVBE8bPBH2jcl29t82A
oEWQDda2EGsoPLIvKxiGB35Z0YiKR9/k9uY1fAqY0WZVaRfN3HHA/Nn4s3U7
1wAvy79PNtCADYFPa2U/nRb/D2Y2hup1FEOIigQQclCiMwz/QlTrKy8P+CQk
hzSSjJQru2+IYSJNCa9e80WlC7B3+tR23Wnih2HhWeTbqN13+94TRqCoMHah
eo0b7rgVtsFyYZ88Gteg5Ae+3ao82uk3iTK7adpEC+8U78ypi3YwV8fiK0jO
aiCI54uF86Q/+oio3Uis7lP4GK8af1FjXBbWkXSn5PtFfWjBU7h986CxsWwh
u6lGnAGURcMxGZtYggt/z83iZUBVIpvrCcqMXAZckd/BhfnIHP1qZWJMayK1
fSTITbvBFMklfiIrKKaBsugcAloCCvIK0xIv9hgdLwztecg3lKOqYmwSCc+j
atITj5wB/vIBTk6kPr7eQ6/pzopLf/VhsWB5xXArZQpH8HpKxoriT+oTHXBP
Q5VpS2kgHl9gdaDqvgwcTBhpUu5Q5Pb0CEaVzXS0tAK0JXHsxMBvIlADD1Hp
B1zYf60zX4xAfafxBSMnpEP5fAPkZT6jT0cvzCqdTMNoAh/fnb2Nf/8TtXpy
4aeb4C07BcfyxP0w2DxzItrHl8T8e8m4B00OQa0SO6z287MucUhYoLnHkR0c
ndfshqiHF7PTmSXgUnw/5S+QNNBlvq0x6dptOcfDVAV64Kyy7PtI2rhmr8G+
h8cL37kxQ5T7T7nrQY/1RIjq09Z02rzuP54uxOgq0FgmzDNy0U0tki7mmUMv
0u37kutuhZxSq0qFFt6/lF9/iuQPC+V0JpvpNvtz2pdf4UJNYxyt4U5+ux6/
5tssccPZW3A6jFhss1VLzXm7xKoW2oPi1HHAKp8VWyBGODo6HdeYvhJMmZT1
3jA1jCdiYzsCwmhGNdshqMR8lwuZfN7IIV/6o8s9TmO15lkZuYm5+ipwbgnl
F70sSDm5SbPdLLHsp2qNJgKMPRb8eNfw9CjiRa95Tj/O6AKRRgicfFF76SYn
LfzAcH2yqLJw/sjfhhstrBvFAww6zWweK66BaeIS0drbGz40Vi9dH6bmT3lb
ngIicVxF0Vz7DyhSLccuQf2SEbyCOW+ICn3Rs4m6qpFi3t5Rxk8l0XxvbKTX
6Yne8R80mwCUj4G1yIK41wSHrnF9Zv7hkWciQMHQCBaCuXcvoZs2LEjGMc72
WoHAGlHUdF/dJjnjoHShmghmhlB6H14WYH2g2bpWHwMQ3b0CQaP/E2UaUf6+
XzCieDTiarQUjncd/aLofLRljD8+x1WuLl9LuO0ajWZKhAf//ka0Iqifg1Fr
Zi7LdRRT5uj/4uNR7qqu//sDWKC4OpOxShVjJRfMp2B3AUAsYMXNjCm4qOiL
Pe2cSCbzMJp71B7dMebZJJoOT4EGzTq+v6Dielsa7EG22XpFR2b5vixz9rx0
bRyjz6L6ElKFmxMP/fR1eaLUaPItzcW8VjapUibb78KJk8pe5gyz8WjL8Aq5
V/oV953cOgllgQ1Jd4v2UejaiekQubT4fsnvW8aLjO7fHaw6ktJVO2Johce6
yE8eAd1nnKll3BNVYoJzN+j1C2EBatYpTOi9lWeK45s4wSIurkZwGXhSCWZ4
LerPwhkvNbLt+28lqW00EiAlZ7zYVS1SMI1v16eG/Zm8QSxvKaWV8mEPLzQ6
qZUu5MimvXL8KlJ0tlenvRyUg+fYYeRJcSSYIF++Eb/Yo+jUS9DngyfO2+og
WPT0fPHwFSqrY7SfBX5Tf/gXVrWa6K2kug7wJ4pe6+s9eepZtV44j71dHvGe
Y8irr0UVQsQvUZpwYWn+ZmYpAaxGoDklajJbfYMeVg2ZA7jVz863/welWR2n
j9wgcW5LDbnRg9fxurO7iTlXKHWqb3hsEE/liVw6gPgfVGWGE6dvy4Wrclux
CvWMH5WNxBF2hDgnzV1U/sa3ZI8t0J7oPH3P6utfoVk4CIQmBvzxR1Ku3dUi
LCahxNPwB6OLQg2MS6qBrip5x1GJ41vMAbVDfkJgo7xN2/JRipG2zkIfhpG1
JZG/5np+zuKx+fVWBdUTh5cFSPOcCk20L2DGh/G9Um0UoGKYb8NCaVu8j0fX
Emfiv6g2BA3qogglue8IY7YZzrIy22CcGJu8TLxkPVJ+5hB7FovrQ80xS2/k
QTeS1cuc6yNxiwLbRiyKvXZyVPl5GxE7P8mX+WUKiMwNaZFQiSQ/i3ELg/qP
+ExLZLaw1gpUiZulGOsmo4aol3lknL+sGoLLprjVUtodayopk4GCp4EyGEBE
pWIQj1S5cEo2O0ML4Us9zGPFlkaIfdGIEKOyDYrY3FoJklDmlg1GU3rXtkVI
di9R0Wsoy9su3kDHmu5NK5Wpzuw1mDzlmwaWJg5fcbxDc0/uhfqzoh07kdpb
Ka2eqMyTWvQS00N4Drwee37u1LGgBP7NN8vyhimbM2tvhTIDRxckMnZcmPw1
TDrKGf5e/XjTMp3mSxmSCV3rpJ9pSBg0Vxw7AC6JvnrdSjVjKk5TnO6G5QZa
IjFzcDLtDMsYa0W0LtpEidgfg+PziB37IBjD8aiMGFvK+Xxz/OF2R1mH9Cw7
eNaUExdHJKCT7l9cfdNUiMCTrxPtxBZ5vwbAC7NWylIUZNNG00WKJD3iBQJF
8bHxhGlm0NpVp1DqgpexiONpRz+nu3NqM36oKaR/doMgiF/Z3FXWAVJ5hEQH
vZLt4HL7G2xx+Fq50AhEZWy2qU4AQKO/a1sTHdGXB8Ojd60HGcbXDA1SPxpw
Yl2KkU3ypursB1xQPqDa6+/Cg7rZfUevHFBTMUH6UDN6dJz/jsjyj9kOFKEI
mpFQqVsQwE1j6fAz0fUguiRUwhrvrZWgDXQF/D681kcs8YDomnaZ6sJ+bYJU
NOHwfwYS5H4QtXnAELn1OIa5WGgAhPR4WkYxnZvKrZf5XdEOrU652jh4klEm
jMgBKX6PNKwMNc0KWFAF3tV6XZFN5b43MBWfDzxcKFzfZSePyO5M5SxaTwWF
LoueVJ/EK/jCLlO1bKNGZMMf7kAG4zxESBSwEynvrB19umbo+p4GX6ebBct7
noFBOfkgncJ2nYAaHRBa9kQRkRVNk7Vn2zIbG5GbezjNqS+JSPpqwMVogLrY
IaC9CmrJZtX288+EXoM3CyUFPR8k1OsABSqBb9o8atSUwdhV8EwOUdTim+MY
Rkbs/Pp5x0KMyN5u2u6AQ7QopxrsPrZ0kvXOgtTowKSFwO9UUxN/i8hcgIxN
ULwuIIGYvyunlkIFjGyFxx6ioVjboVLrhDMTFpM10csuq8LuvDUhFEqYi17V
tEZIyC9SUoe4YbbFv+Lv16gchUG9dTzdGM02U52wAdmy1exjpJTcugWQWx6x
T5DX7PzcQQtbJYhKMSJyEORASPZBhDdgVSlZUEhY5becs0Ux932T98NrGkcM
CdMNRORqToU6sAwZ961Xw7VgjIQqqh11j9JVubc1SmyuiuB6ckfPDC3NfRk8
4nR2VgYyNITZOY7peBvqKBUl0Cc9nu86rBn3i3eBwl2lTSLgSjPc/ROfDJTm
LbefCFP9ha/eP+tFwzaVypevfd0NowOU/LMzgbtG0sH0OAFrLS+Nq7NBqcEd
Z7KOg/ItAadW4w6Pg9o0LZsKCvFT+7PbACURk62JQcZuyH8U+kf/AaSmokc4
Jjdk0CSaORFJ119gth9flqDSmVtvjq+uuQ4J3KRTkL5UGr7wWZnDNGqUCQhS
PKrWI71NCW9qgRdeq4dCBxKc8LqQSrpGZ+7rp8mZC426/YJoIQObGkm4BuYw
Y42q+qmxHy+jy63peD80sxMaXssJHdb+PvsPditS7ScxvmqeCTKlXwhpfz/I
hTX0Mp2NcJJx13GcRlxny3OarCXbkP3qGm6wSsnPzsWAn/BrnwToqamC6G0B
C7aYy3z+I3PaUITpsWmx7fW2yP8k+Tu9cPs6YgK/s9kSwbEV/yovx6peYzPm
/dgbouCde2qG8VoDHUc3B/Pv6ds+rogudlwgfjsfY9ZOZEW4keR5sib3rDQN
5p6ISzYyjS4wntPgyHNZSpa0yKEvPAU/pnJT8r5xMaEgRx5d6E/tnXt4JVrD
VGe2IFvwU4CvsbzvqPF7CrwRyc/Kr+uNpEhIO9XpFZMmlsnE5IfEH0gYgMX0
gFz8T8q3ClS8dqfmwuqOmB6s5x2DTC7DQVjmv848e2FhxTrGWwqAUHP+YDtJ
37AUc4ouGqC5Q62kGFuqeamwQWk/VvHsiE8G2rnHBJEzZqly7LRoVS06g8x6
rP0YhWnu701m0HHMPH0TvQni2yApbk2R7zhPwIh46NHxcuWT0s2DwSqaIXbY
WR0ztq5SRZG0hXjaVZ2BqKIIvHMEj++ouFxr9CHFe+R+53g3jbW3uQqSzag+
XO4bwvfSEp1udCg+UsmRp3kiHupct37VpmIhgpe+mJ43FY2AssQ9loG0o9dy
WNhvYvtxC+jkiuttin9u/+fL5Xj0aoWtEojzOafcarum6FtWqhZJjbykwIqA
9iaVbSMUbRcdlCahi4v1FcD3tP+4lpKmDkZUIN+NyF1kyrWbMPCI40K/994j
O6Ni2Vy/+5neODEhQNcyLt9w9NXY3tDWz0X6Z4Oszzpjtkc+Pdm0GWMIFgxn
FR1AQWcNECzwWETYmDPKhvC5Jm5gMnocmUipYEMZzQ+C5UrLE8j/QUDLwQwr
6nPHVQVqMgKqUWj4UHltM4N2i3N1H/0nZlgAbmVB86gqBNljLOlzC3PCMdM+
OLN3IQL6WeW+65aDkB6tKtZAyHTpRpWcduDEaFtnJEqgilftUF5Ltdo5cd1U
3/XwJZsdawrouWG9Yz6odF4NbeGO9HXJxK8X6R1yltRfka1tYp5PbqBfEUgM
JaChAJBZ20vf19lL/gEjaeCaj5n9DwsjRBgQLWbUvz6qi2S0vItas0ULmV1o
EwBCIOnpwPat7ri/eIhJGXkXRA7v13UjbLUM2pFow46UFCNrOSv70mRprETL
j2XkHv8ZA9fU9hfiOxm/qyDgvH+ALsadoR52UzR/AwguCjCwoO6jI6AfdLVj
Dk4DYgXBMx7PPM4lI1WZU33seWMalLkNAX24t4zXR5LUgdgOyuFpwqRrd1OF
FO775Ka8q8m5mnWoMyCQoiqooc3k1V/PPfS16PVG90b7m+k4hvAUyaIfga2l
u/xDuXitG9gDEpTZtoBgeicqgKm9bYH/qNmOAbPcK5IaEHM9FFhRpIKLZ+YL
WKXlPATiAmwj8OFm6OEtAd/B4wBFCPNAl4Fm7ler36cMMVEwHfOe2UFHKHU1
X4kW6DPjiOSmqtyCcTsaiws6p0sNMB+pnRsW+WEVoN3pVSxQO15LdXrS+ABt
7RfF30rDHS1YlTvbpcFE3LqB1N9RoyWWqpYvzCi8hEwIHm/MbaYyfOW6tq6F
vTAITbgM0OlwTAveWJEKI6YeH6qmmqZ07R18FpqR+1ayQ1ewbDvnri6xZOYo
a4fQP4AZuzN7GmxlV2cvauhFGdIVcqT8+GE4LvoLmvAESsrgoX9p1NHFoC19
RZaZGEbQtL/bfoTZs4Em68AzY8tSFfvd9h4FoKAeXdKmklUybs51t+EBjnlG
6la8nDqOElXLXOBagqKa/SuNboyPPvKKBeTzK1jgdk+HAbEPyrZKHq2zK1oj
XbCEySDUjHsw7T6wiaBm4OqDZWk9mVO8zAWVm0pxK+FUjnXz6/PJt/VzFuME
1fBVmE2d8HFxdPHoyWGaiCc2rpS79PMBUNbEQPP+JZ8wBPi6H+NZtg4GJo/4
9pwZxk141PmAzPB+vTv6/RwmkGHYlFN6eGMBSziz+XxYsktqO0INU4u1TUvH
HTfnNZZMHu7haXCPf6U4EYjXw/ESANJTGkydTRcE7m+igmqlKwIlmoatMO9Q
3njA7KVnQKS7FcZc/KLgSZd6bQR81nfkO04s1bMbx3luZ51s06ZYJ21jlBHZ
SPRlk5qW7FJgksHeas6LitrGzPtMbOIObYBuFP6PEcJTz9S5aaFPNhHaWYFz
4R0Ehj4VfRq9aC7WcwFj5EGfnJlUf4icdBw+3Nv3gN2t0psEsB/iVPEr6xtg
QN/0gl7PpJWyc7b+Hpr6e1lWPcA/9+KhosQAYgfnA0MFFOakEUsxdtXtByPd
sT5pKjlEEa+qvNd7G68VNZOQ+flxhdSgxig/SDRr1MbgE7m8+6IwUgLzQl2H
imywuXQkLtu91jZZ0rrS0vU1NZfPrGCaGUAm5GAWSbQ0VjkMEx1cBU0J1Wfz
DbIbypjGDdi/xgsw37b/sFooBgofsRncauuC9hB87WiEsDjh/soJ707/bphr
01qZ2N1vh0771zWIcW/Wnqw6U8UBWc33Uiu+FlUYsfX48Xlx+8KcAaKwCffa
U5zR1qC5Cr0Flbev/LfdCbBkwpF2/OX4zPSv2E/Z4F4OKkHQws3zLXMUeAH6
YonnA7hWFY1KnsxVkDvG9hEmmhG/s2JtVA7hJovZuyQOVKYrSnXTsCXEorLH
WeMdgVvR4YWbWgbNb1TQzo7ot5VgZYSUQTosUa/FfN8NHa2Id8nPL/EuGOG5
NzRNedbhnlbboNIDW0yC9Nch4H0jxgQ4p4MLMkcKUJG/xq7hEpDBEEtC30ur
XhXnezo/ZL82i4YLqsr1KxOLiJt8faiK8DRXkG6hh+OPu93GnGK3otghgYNS
GzDIzxxBEgaPOMYItGWCGgOaVQ0bIMmqsCYbidGb3RhYvqY9q2BwoDFJZ0Qu
laqzUDNPLJGOpQs0tfWeuGItoFE7Pq9JMeTLaJBxBq+M/pWwJX3dpwjMFD36
VisU19fUuz+sWuDqt1oVphJGp/BkFRxjsz2MyiaQeTDuOqJLjHQiKg6YPmND
l5EWS8NiEdZI7A4iAKLDPpsUgcGpPeRGZkXPyONR7RWRHdZnFIC31tSZONmG
gA7mVoVxAqxFL9V7rQUI8PHNFx50NiCh12nGjE+SB3iHyV5yLkaOApmZt8ja
4jfZwFMb0p6K5sENjLSc2LaYgfLg3xyzvJcgiq/F4rX18XM5WSoK8tDCvVCr
Lj8JcBbjHi/R+Wx7SeQbaJ16AC6bjgRF1e04cd8TfjQqPEMYMV/EjFTSSvFf
/Zcma0u35ObMBwgNK7z4r7fzZUNh+69f5MxgVXCS0OgZwCF991l0t3vjbAn9
JvDCvxxPdzuRNq+cHr8qLyYAS6Uf3dHvm/08G/P2Nhp+7O494PwKL8cYLK+o
ILnB0drZf19yLELtA4SjaDip76uCAPdbb3tzHfk81gPHPQJblViJ2D2OLUUh
B1ya42hdlgpcC/IdAk5wvbMPI6wUu37OLlYpdRZNnyt7PbfTyC2xcgi7gR27
uU0VEadnE2P+9FOGtz+iwdWxfD4VdoxarDEhpHckTX1IZ0arCy72Ier1jQGD
P2NBTPeZkHkWt1ds+/Z0qdhJDgrFKotzCSe7ZEUpNQmW3lSkfwNSuiglW8fa
iiqm03MhscA2l9Bk/KL+PjztxiVXeOyihvfCGr+1xVnChJ8LUgUOG0bQ0atK
dR7X1WD3OipgSpJljIk9Q3SVuxeOqFnyMRLq2e99wMvwaAtcJj5StX3uwbRn
qkroomn2FU5LIpzn3mTiv8+GJhdrPzpk/YDuXmuxW0DFJf1m6pbRhK4eBgdA
vPT27j6YoZcJR1uXGBhl5wcLdnSVQv840BA8jev8eWSol1WGDZgHFcD6lpc9
BtgsGVtfwv5AKwpFlYN+bK+fHHpWS12w6TID4AYwFwwotryuNawx+FZuQKbZ
Fg31RfZu6GT2NEMEsMTYe30vgAwqqcRNLlCONekpmlujrVTNxuDfnILnv6Td
v8c85i1ND6Sf4Uhd4vHJ6mlkgVw5DkEehBx0iJZCYiOQ1E584Jq7rtpOdcf2
z5FWJbHZ+5lbk2SDx1RamrJpGlMiZLZW2Oo7t7SHs2OFpxCoZuPttxDsHZ4m
Tti1dwmQjySXVVEa4BH0KByF+B1icHo/qYckVtlmJgDDhrGP3Et/BgcqGmm1
H1YO3uU027T2em/w4gy1+38UYT59rKMvpBIPEqQ9n+UpSPLedP6aTOmt4Elr
WlcJX2x00jWC1Od0KS3ubSIEeNt6DlBvVsQIy5AaEf/Jzhr8ndKfLJh8xNfs
+Z0MuYbKri1RfNIXhr2JQlurxzzZD3r3VxL556r8T+dm6J2xsMGyO2PAsymb
A3FOKnJ3vqbJW9Cb6mmZOaM4jNiNTFr2ERVdeyVWFFG4SeQmv5YLkk1VGBJ1
+slCx1erl+m45xGwJn1sdVsbrS8XKzYOYmxE3Hz3yDsvBnKHBR1+ue7yj2Rh
1RqfkneOf6yr+ivrms2a21q0MMz0yykTtrUjek5SN2AO6WfvBLzMkwXUjMLL
XP7wdaWAGQs85rsJnwk6Gq+Rr0ABXUVGiExrAfkWea6TbKPsam+UGAnmMAmp
VsCSU1beaOmZKjvzP21U2x2a9l3Cg62mhhhLympAHIAWsMQMQUkjOiAqz7Dw
9BZvduOv7IntmYSQkNIW6OotgvSIZ4I0ho3u2dif7Vr/14Aey3ZxcCPfyeKf
KtclsHRt0SUKIWYa/UjeIUjH0+Np98CPoK/cvvmmB8eqdCyJ+QXFK489KvfU
zhjMIzplf/jfep5hf7qziXWxvYY+imDFhZuczt6k3yZwjov2/wwlMwMUd/Cd
HAZCLV1UfTqn9hfPl5P/WZ0QHhdRDtdHAuUV6mBpgClZHMenBmQQ0VoPWDiV
cjrkPO1NoSQCOrU2iwvfmt9r+uW/LkkWbxiX75MQUfAxujQgnsdaQq8hCuxP
mCr15g0YLryU0KeWrxXOOFq1wf8ZtWwXuC9kqIMp6X19dVBUZGI1NFAPrOBA
RAKadkMFZjz1OM+qyyFSOw9/eiuMT9eJ7TXea1g2BVhctdND5Si0IttS19X/
x/ogODqYxDwMxLbjta6WpnLY+A+Mv5W/f9VeKFhwx+F3IIIcvhFKmFKC7NFy
FE40TAk+qsOPoofqXKkBcYVdQJOj+Tdtq2fVbJv1+xsZ8G3oTxX/jom2dLde
jORDM48W5oY0LxzKH2OqNEu4ROXnf6p8ZsK5Re2McK03Dv/9DEDPja1DlkGd
G8jWSUvRv/s36xEKrG6y/CBvnGsiDXyXxAmX1JzuQQZjoSdKG+Jkdo8HyRJ5
+hNLz9f0IpsENTlrnsP/xaIagXfq85Z3d9QoEooeoNwL8E85kdPzjS62Pthr
fR2z7OQbtt+LzJ/BvKN4JKlc49XepGtRZkpyEt5wvMUT334Fn3xVBhDpgyDZ
Kxwju2tFepBjTHnNCI5mkV9pHwXjBmxH33gUNYbaG1xbo8iyTA2b22DbYywR
SVmVQpBidQW0QNMcqryIuXDuJPmBZc8ly8QtWW3Dkx4QLj01+UQyPhx7AUhI
7Lc9F90ywB4cFmFtJAzJ4yX4Nk6s2/CMAf8eQ/ckXKoVjQg12IUm48wmf1dy
Llrb7cNs+LUppgc0wx6csW67ajTNCgVAXfeawQldzIGGwpScY50gFv8J1qj6
rZm8MvKZQL4hqp3rb25r+NMcN8bhtuOOr/+34l8nvIBzuLH7ulOXtFJ9qcuE
wjeeUVa338GCX8/4pC6g8eQW6PfqUmjNwqiBa4fHIiPEVIrvUB+MMN2tFw16
1aDSNAKoPoZF4ULfvkyBMdpU2IlyV47Be9vL+R9HXbDDfuQafCyuK9Sp6H+Q
2n4nOGT//GawtVvKHrdKPiBBmLMKRkTz5kWQ35UaacDMwV31RgYyP0pd2Puk
fpOuoob40Xtc4QiNXfHYOKXyLE9QCH0x4cpJ3IPrjkTY19Ot6JJNIHdCX7YT
7Uuz8q+OS+PTXCEPbA2Wo70IPIUN2tgVB+RTB0LZXF58cQOeeoi6slNrb9lJ
Oa+KDzhgdVONdS+p4uHhIlcGHe59FAVZ01mvsbpCKZxYnWOBl+LwNB4vYzAt
gBYzJegfcK/NdkbXyS9e+mRTz4ykUObwTN1NRTQeKJdXdp8AmewIJjrOmEvb
GKK3g77zVdUtusBt3zx76KBDSKFmpLhPusw5MfVyI0prFZcATJKvuJFToC+B
jqpQ3m8MtL173tvBTBQVE3nkoc7L9LCD5P+++Svf0FRAf/RudGkTUYxKeNRB
V/BjCGfZLsiNdNcZ9QvEn3aAz/AT0RMkMSZTIyYMoxTEr3QpbJQ5Nf3LIV6x
ez1ZNa1HPqSwQTrjE67eTLu8ivp91k5Tk0ly2xO7g70CHEcPl6hNrb8DKoyF
nUQl0oPaxcVQAXCQV75jTa5TEpIHhTqHhgN2dbdsWvTk3ZdyoZMiRq0V8AJ6
xR9vOe0JyI9WDj72jT7hsi1pdrJVt+NXRRHOeiVQWPCTXfgAit5/YX5pfTHF
bO5MDfJTP3XnMQRGCrtvI1jm1Djt6z5Fof5IoWhbjdYK+YkGrvG0zfqg8LJh
TeJ/3iJ6n32VUzZ8IhFHX5FDLy0DYeFZN2PnXw/qEVj1X+U8uAxJ7XrJ+PNw
H5WvEC3MQLasAX6ygTLJC76f5y5rFSaCSkP/M1taiIEMV+FEkVLmf+SBRg0f
HlhnpH8wVNtocaWSdegMRU1kGw9lttBIiHjgiKwkV5YiPY/XmDR2Wm8f7ZlZ
xLYoMAzXCNhE3JaitXw0vtr3zS+RUA/TfNcELKEVOPtcTAYPsmUCNZGklwJ1
LLxJ0qP4+A0QZCo1UQI57xooy86EM/TeDX5LIp+o2j209wcO0nsWTf+9vDPU
BLpyiTMsYnDQtPRnbL4KV7twFxSTdTkEP7qsFjrHPHyEHM1aSwvMVXpz+1wd
qv789VOeKWs4o1odzFPrEzU+DA6SyH9jhtuvTgt7CiohZcrip63nM9uxOmrP
1uV4GgyHcHOCSE2vxQvnjtwowLo7cWiKedouUv7xXr67+CYKWl+MUR2o937B
4hnc6RdlpJYFmuKVWjz/26uhIsk7l3cfENslobrmDOjGAOMX4oiZxW+n8kW3
UGzfSXsEJfcbGcOXOz2gRRsDsTw1gkrH4xjinRcrhnAGrB86QOJEB/ik4zrq
v5tpe/HyeQMykdg1lqzZWQagBb+GD+IslU/CSt81Ba5d2kLQ2Q6ESEyEAuM5
WW6LuKojbgIxzrTXUQx0405RrZ4Ghy0RY59VGttAqgXk5XmOCK13YVv7rxhA
o17ZopvSDIKwMHse6cmG2jU2vxSus7XtbQeVyF8dIue3n8t7vOPNvdI+y0l4
he5LSr9WP7EiTuQ1p/c8EyLSu7jOczNTabhcLqgaOwL1RbylhFrPL0ls5Wxf
SWhRTc116vwmavVkdLsEpyzA3l2Lz7T8I0246t5SPdWTGBxoETv0rQ2dQONt
lcc++1s3wxGV007rN1kG5v6eWjqQQCFcWmaPq6GDgpG9ZweDoLLoj0FsnpeF
+cQ8tS1yzt2Mz42I8C1Co9ptGP3D/3aiYTyUESEH5ut2Furf+4lMC7GZzgv6
dFOWuFVNLD6MOZ4azMvxHOZ4MW5gZPkLqBOypHeY61zEAbSSCD/3v+1d0F4D
BR1MqNj2j+qawiMmmcYS8gCB8TICxiFuxfUIfSe/FyQkblg9e5McP268FfLw
fPodSDH1IQofdxQNM7lYf+zfCSn/Wh/n7GuS4klkBFe1l7a6ZBZRZwFY4qWm
76M+F6vPmR7hDXvmMF05gEaIkXHcgcvRhd1+undv8gw1Cy0Yc5M9ICyJrtrg
wnFTAHp2IKbdJ589QsnYtI5SfXqfb40IwlbtN1FfZISJCiTNPmNbaCvdYURs
QJmDXwrKeZ8suFRIJtjhVAj3vG4R2J05oi6yOEhrvZk5EnI6sUKbMk50QBo6
BrRO6FWWC6v8odEVLvgTywHfej30St6Xn8QJGQqEz1o1243Z9QKaNQEx0sLD
4LHoqobDwvTM+OYmwMXMv1BQJMUkLFSwTsO51VvHmikKLcQf8JUB5u/36s+x
iOB/V7p2NVslJU8lMayhiTnXW3QkEnKdrqgRNKx6t2TgUACLO7dFLUz0b+zh
BTrl2MR5OhFZYCAy2Bcn0EVUITk/oH7FkULa/eiBUyvim3cAM/4jRaE00UAb
VgiXCdbn5g7F+AtSNnL4KzYlbFIxHmPkwO5THy0WTbicIp5JuTBYtzR80/tp
axm4euKSZ0867FlJPA969jQFnhZthbx46xZe6KyNFTzftVo+vO+nwM9PO9Xe
ZeKt0DBmM1OXS94V5WFtD4mN/Woaypj7VIFroDUuGQV8DyKCq7woqTO3HkRr
/sM2K5ESo0ywiwEKBsSoH/y0BaZXzK7QJ+LK00bTBHhsX0hM9tBjRcQdPtHs
Wb1yOtinhB+O6pGqzqDXiQbngZkLPsW56VmGoxd9j63hx2SXKV9w+B8ZXHMw
YRI1t0Ya6MyqgWq/mQJW2XQESzc7rAaowMoNz+xOqn1FaLprajiCbh5HeQAe
jjQGfNA9zwXwXJeLEYIXd4oLYOeg+GhlLOz3ohz17mqwmZFHpq5Mt5O5pw+M
WlsD4lyIj3oqpwx2pn4M2qh6q4kMmTvpPKaijdgDyg7x2stSYCh0DBMOgr9t
kbse5aocunjfexGuKAz4JiOJrBFX4htvgpMIshWGVFhUFFF7Ryv43MMK4ebm
4FMojH5GZl8SWcOGagp8xqJuFu96JsQYSRRDThUFV/Nwh+8Ejr0zASvnGSkU
kn+0D214e091ewUO0A+9MH4nVPPrho+4fyRxeuqy8haQNmuWq1njNBd+gQ/t
JBDA0RmnnR9didmVIrn/B6gWiOlWRLdFVIdFjH8ZjBGU5ZgURobDXHy/WHQl
NYg/X9LQmrm+4tA26f5i9OzBkR6s+6ZMYoz4Qe04SJESMRaFAQoixYGDix8f
e9bHVhPmt0pflGa7XAp9h3Hpoce+QJlwO2ggib3SIYjIDhnCF/8/lxe5J/Xr
1Q4nD4F22Qlrzb5TiVVMpnyNRb9acPL4LtPZoK1odVVzoAM4g7DKGHLIRBIO
jH924yx3WhTxLavXq168xLstnGGPt27ZoyOvilM3xQ83vMXDOLBJqGOssTdN
aDDToMSchw/Yd5jGgysMZcr8q4THxMsWwL9/QuWWzVwxwgTeTaRHgIAP5n6O
ow8Jbdb48nThN3jO9V6yAEvsnCWpR4embVR8wmykY+M7bkk1v+R11t8XyEvs
QuKAA998PpM1gVxNn/JIoIlA+WivZUr9Im8DwyEFgNpWyvQrHiivlIV1fdRL
VYp1u8TgWv315RqRo7Y8SKSXFNQWnh2Ykytp25JDvInxI/yodT/BCagrxoJY
IwMxDaVo394sC+haboPaToGrznb9iOgwbVuFZPMvuyRt9W9ehrhaHRlycacW
W91ogn6bCHTWojXFD4MKXqZA80Mkbm2O0LWMwQv7GaWbVr3nEylaXSz22l+0
LIe0HUfMLStPpPm4vxB57iqKWAvLsrYMgDFxe/AH1R1MXt4Sov9BMNCDUtx2
0GL1lfws4C6huVENDaKOk93nFUvJNpF0mxfZo9yvRn+oBn2TMb8xLtU4t/Rn
xaT02gZbVsvXdH4V5CxsqFVpM7+Uu66Wqmq2B1GeghvPQG243+qd8fHia3ej
2yNNjGA6f8sY5vuk5Ofr0IM9MgggMjH/3+Wm85VWms7rzeBEDsZVaIy3RViI
eGVO4EO1ZMo4zvjdIUMh84S2vl4SgeMoxbtApoJra/Ka545swBsZeGQKr+0/
UA9rmDypXqo7/nv6zHy8QQ3cYidH/J4fKdPP4xtBviWTUW+O9YxqGhRnActf
VoSwK/4IUNlZQNr/NZVdFVxwL/7xFKsT05GYr322lMUet+5bj56SopGNyK/E
WIo1HE8kyUCHmEb7oysayQ51BaQv7/YYVHsMKe70bzwZ419zwhd1TXjr3epe
lj6IljxIYAXWGfZGcz2Xf+yH5hbGQJbgp9GxlEZ5IaK21vUgh83M4JLvIAHu
SiGG3/JAoBiBhR5UfPCTZEbFBL6rFsRs1T0DQ9y0iyAYrj2hs4z96skJXWuI
DInzhlKXPG+XvjUF9oj2SLAYfB2POCZzpP5B5BOIWFG7/Ma9RJVSnIXMv5PO
uQnkf5HWO54NZrooimtwI8aqEwdiMwREU0xeXVUHozZMa8xT6Dy7Uy0YHeAv
5aHnLTVlkYPpaBy1RV0c2uz+8d75IaMuSrwvsnBnJMWTQthZrOEkn0XY05b/
FeD9YhSOXl2BMLa0ehEnsuXz7B15Wx3V24tEN6YkSMRnYtDD4yWgRzCta+md
S0KqmA4Rn6rBF35jD2NAIJQymUf2K/Jg6qm4+DDcxtesWsP1BAyyCsvkSS2D
/xcujTTLireor8K0HvpklGQVsOO+2VWV106QauEctcLIJQxxNEKn2nxvA1qd
WFCuw6GrayVWUeFJ0sCQcqLlAHxkqjMl5irEQvT56fCq6BcxTbuJmCBIXf4G
457zKI6K1B8i3rG4dLbzfl0nDWHu1MlGi9PJiaMcpVEpR9NI3lu0qYoRw9jd
mH7ODDHQlgmt1jb0m6NPBKTbnsgTDB131gAZsIFXoWygaG06LXDx+uBotSht
l74Ikd/rx6aXUFaoESX1QXwLnwm/c59d5MKtP/gLWmGLNEbdFi4nBpPUgh8y
GKCpdC/uCdI7vYWMX3/0wMtFO4CKsSEY1ZxzuzSjlDWrg5xJ8ufGEIhtGQ3q
hh1dLCBODR2FzQ7PFERE5WFUogKJ1T/QsYez2LW0c/jvE0+P0P7SbR8LW5RM
dBRbRTy5RdgdsCiTtKONIt8V26ylBCz8r8403J+grVjvjWpN1eiuIHpRQMQ/
nZP91XHUPzlAfp8sIC2wq1dFGJu+pqKw1ppbc0G801wFFKqwBd+bpvjb9tzW
jqgARXvyaNP5RBNC0lr/A2kedZBuBNP/JDOMjlesI/GKQthXEA6nM7GfWPT8
wfG86u+UJctvKgDLOqqoB1KfiM1RcOi2YM0uFZWPMuUJQE81BzK+h2n19mj2
guqzdjk9UcnzR76YHd9UlbwxjDRBqYk7LLMeX9O+/D4Ej9LZDGpMwq2f25qQ
y/QlXHem8NhsX76IBRtYwKI0aq4YCQRqbaYr1UisBzTQIWMUjdN/G5S7piCM
d3wlsSKKMb2DwLWxogQiKLp4AxS/K0vMojUeqYorusK7Qb9PQgS0P1V2wrcQ
eukB+rldlrebIgcchWPLt2CvOL+nN9rLzcPeQOCaw1+9PwuoebcYf/z6vs1P
IfhtqUt/P+HwUtQwOh5/HNJ8jMNA1syu5Le+LX/R/AF6bEDiAheFJAm9+QF/
GHJJElwFVyl7KgV95/7j0W1Xq331FA0NtamvuARp59lhthWTyoAYaVWBMROl
92sDoNFTITGxWAXdD999hKTT1yt5BGaHl3xJPixgY6B7ZeR/NdqyGYNdmNqD
vE1YD2XRSCvzF8XMfUDctqmqXohlTkovziuiQTd1ciTSkTU01aBiVL3NDjnX
UglM6pFIzodUmMwzaSdjfnvdIhJfqoszO45UDOtZo2a3xVfetzxjffGJnfYP
tn2dOheaUfW7jEF8eGLhuxO9z48GB1rLr+HeM6x4445RYDZgVWLO3P806h8K
wNfZNc7ycIPMGhw5hQwgyPxbukwFd/BQk/AarQGzbaTScCkp4K1Egw5jn7Bp
BAAIz6k3NAKhGp7CEIs0TsLCXM7qsBTLncJw1HRmVebCjWd+6V2l5WuEQDx6
s4FUdR72uAnX1ODR9lDpw95zpiSnFivB3acz4wyn1/H9bIkPTIOLwNzwYBtx
nTMgBq6osqbFiciOKvfj5jtnvJemFDTnukpQF09cCB59zDWzvCU2Fmn5X471
9cchGEIbu2fIb1q+rKT613IQY9AnFprlshWn9I0WvYZLfXc/oPx7wENPJlOM
QidzRh1S/nSVygOysWaslzmX1xfzwO6POWLvp4cjI9mYTO/m+747McPqzT9S
aH6ZwWSzl/TCv0y/g39/TNgoNQjd0cx0c3M9ux6cBpVVhEBsgbKHegP9cgWj
MhZbiwFZMTzQbrNyejv5a4bg3Bc0GgrMlWKCodjBHvXz2rsCDOgBta9Dvi30
bKLeX5A8lVKcZ+UG7Oni6CiADVeER4Bu2QGmqbg1FiNCDPMj/bLcKBss+JsS
g0Nlz/Uul+T1EKinjDgZXS0HAoFCQgWu67lR95Zma07ERoVtH+t5z63OfgO9
/bdsCVEoy3V/zjedK3VaXrAhKAwbUCv5HbQ7N+JULUbLXjIVUpdq2tXPcIEr
FQLY3RQ5QAxZcaGZIVQOEjpnHNP1R0axqxEcBsEAECCU83V43BV+W5e3OYLd
JPklJx43Hksvz9gG6Vejm22ivMSAuqJXCSHIqgG9c6/78v/rY312p7D2kdZb
Cg4A5cH6OGZUPyCYo4wZwdLXGyTSmpNe8ZITP1pPGwC6fwqkCxRDAYGjsCdG
+yQ26NumCacUozP6VY7fn89RsNivz04g5XrSaNv7+z2D4uraY2cQpG+skPE6
/y4YVODS473LHCQAVmbSQ9Z619jchDg4gwJX48NShYVdaZTfisiAXPSWaUnU
UWbfj7gjQ5JTYIiAmlRm4nfC4vQrpKu3Rx8/9EzO7BvwBnV1mOR/X8uppRMo
Olka8y0HDrBYBNqIPEN/IlmcVoE7Pikp8wZPvfsnC/R6y5x+hCcFpUROx9Sb
ZWDJWKiGBoEYxnrf0YPUEYukQfD2l3Alrv8JgJNPwJr384lYyoK/vSoefQO0
/kGBfw1ToDXD92KnckJx7PX4YVqeJCFULU3+YNeljH6uI+FFO2OIHwZDzOD2
y7DBbKu6BYQV5+ToKN9fxdB8FNLNSzJxUskoWYSaxOVwzszLvLcN+QtISoGC
jJPNrzdSgNmiF8yADpBTgFEm9oXnSjmWS8WRDHAvej7UlOF8MlDm/OK/AWkK
oJlfjafSNER9VzfETzdtsnlH3OcEcUqBXRB8+vuJGs5eOUXtq5qdNTx3fQoo
VfKBHupRV46PfNd+7i7Mi90KYUVO2rr7kbgSvzF6j8kPekyQzsMnpqOpCe7E
YxyUMFAJiAeHe585j2nG3j1sIw+VW5346aGWx5NfaNZ4PpElYYtZMh4Mz8Oe
5v91MvV+MOpRiztB6qw1UQ6h3CwYecxRvoGd7lBhS4rAHw8lU7Ze6E6AVIaF
/P75CZU7ueZzrmXlhoAL8k1cIJB9P13Xd8NDoVXAPQ1uSysGY8LJoF6xYwPb
ebN66s3WmprZeZQzy0XXjpzZEPE136MsAGfkAWVZj+vDPaCteMqxq5RxZRwo
nxngPOpcEx6DmkEmzdYvI07zbtKPhb2yPqNiKcWi+kpbPT4ZL8o95b9ic1K3
Y1OZ77gIr9ZZYK08c1r7STftFNSlMcC0kpVyUWQ03TP+gK4n59PR3TRTLQ1N
xcybIuQUihED90SHcPgudRBCy66CWJBYZtM80YSKPa0gxOIJpsGzApLgqSD9
MRPiovvlR9g5RxlpOUworDVEcQhSYGqAzWFev8sPSvJwIE33fDb0yC7KH7aj
0ALDfL6dKKIKbAJ3CXat72wwNhnYPJmNtUZH/LsMu9FPX7yZ3teUko97QRfT
mh0AAKWYslz/LZ+OSvkbUGToCoAoHXUiYdtSYg+JdLT3mRh5cFGP41c1JUw3
bCWpRMtd876jJuUh84KQDdcix04Y8JqxFxC7k17TdGoLrIle0e+yjYOMeYBD
YZgOd77qAZ6fMubgRxSWZf8NJ6F2QozkumT7Rfjwz7BvD4odHCoy5/JzBODW
CS3dlC0aDBiaqJ0fXbNknB9hcAFvhCwe8GQheddMqqR/UwtlevE3OiMcoJVB
Zbw//5lWNnQZVc9igrvt/ZdBjDBsl/FKv8IhMm0LnwjflbsrtiHsNazvmkjh
MA3r57aQhlOt3NGzmOSUjcxA6LGnduRbZF6QbOH5xn+ccZxW0tYKz0syiRov
8drFhlCBekRHGLFAEQ5m+lrAItKpocwDAXOGcCTFoBJUEuLHWOzqUtowY2cQ
0z+AzITRJziVnH4zZdoSBS1i2tjsuMunVxmNy9RXluE0qefuJpOlo6MFjVK4
F9Tco8YNiqhYDaiceakuP/6bvkoKYCx6mjIu6Cv/KFouTSTXjA2/OcMJFQyP
fDng/DU3iKjhlpmf6iRw+Gt89Ha5VQrKzgGKXGtFvEjcZcQqJwIVg8UNRshp
bhpW49SxGNLZzg8toBpqWxyImLTBGqOfablQm81wZU0uinEJZ2/OctbQIqlJ
QgtHQLbweNZ9R4TNXtf4PGunaysoSPdC4xkcDCv5eiQw7/JhL0oKqFS8ZLXx
nOcnqgoe/khxKNDv/jLdcIFay+ivYQmly4BqEY/Y0q1vtNwVCY3kAlgeeTr4
CVLwRm3pzK8am4Ee86AokUO1bEvjCKggEx+g6PokMHmh72xGgpx12bfY72dz
cYoCHle4j/lKksNzXJkTSQ7Ac+swRDHa6k4+KtR79M8z8qwSPDpiV3embQlY
mnLGsnBUTCKGEcstGNcmGJCB1KEZ32Tr8zwTooLZz1HjsNHoMJdNMrBFRSlt
H/LkJQwmsWbABG2JXf1TT3mv2CLnToJe9w2gduHBl6VaSzHJRMBz0A4bV2Lb
Ki1rzDutfXrTogsfIeufr4xVZlPQ5mDMAo219kPXje+sWrcAkQDaAF8iVAZ+
iFXWUGFisnYz2CW6DAviJG1mA1F7+ytEKTgrEgZ7C5F3l6dEDBNiKHKXWF0J
V7SHmXmkeeDtdqQs1+eL/inwtGlFM47M8ciCy6WQTnN5tXki1WSkSSNMy+q/
JP6Zsk1XAivbnrpM3FZ7lQZTsBfcEXq0847Fbgv/ct+gk0Y4CK8AuuVBRFUQ
KOfQtiofagUTxAxbTVBIc48PuOTVy/tskE31G1JcB9FraxHTUMIj8Nx5BgXC
iyAVx5vFf/p+YpFoYZvCKouxr6+j8U6PHklFYsW6dzfH7Cqw3ahfA0CuDU9b
tUnvu5UaPLyzg6zXuwsaBLDX0x14fUBBsuta1KiOmoHlNXucchQhpUVUr4N2
tL6MsQXuBdlPse27SEvBd8FohDwsGtR0WCcjEvpAy9CTcXHNcAhBIjxHQ8c+
TunMlS1cJcT5dTlzT+AjvAOzoYs5ADwqvRffdIMsSiNJi0vIsUAkDIhOloLw
/gWiN3vNGnEPZwbW4xU2ScaqaiDf0O6N0KbEFOOQEuejT2l5PAVPHZPe8Zf8
XUMfCyhxbewk4a6XFpMgpztKnFhmRZJe9fFvErDz699qgIi5xGB07Yf0R+L+
0Oy3hnpeowxjIrhqosdPjgd3b5dOg4EO5pix9FZ5INVaVjr4PdFAn6NxmaP1
2WJeuzbT38B0q001DXLL/poN0awopxpROhLKJnWg2yXIcdqU9/bJ+0QqZ+BQ
Fbnu6HDnYd/LoPKDhZusLNcoy1FyYA0YaRYSDNrOBhBEI6kzc/MKcM6A/wGi
9JR40e4pWENgSWBFfNPez7yeg9tJdp7bx5HDDzNhgN9nQXGPz9W6HBs94MhK
2xwmB59yL2t9z+aU55Er8Zjh6sjdqmDbT+Vb/rmJkUc97h0L/fsj2aus2F3d
35dUl40snQgfaTY8v/y9AAchhIX+rpTdUoKfeB7Exb2mT3OUoRUaYy0XZkPo
ljdqLKoocpBwKKJ84WEG1QwLQO4eF5nFJQRmbEhzsQsr1gMTguNrtgdtPCpx
t/C+lYXM/Kbyqm47ovZJkXGPoYxnnzSe7reKAgJMxljN+XPh8iUgvnzI8KlO
LcxUl7VTQG8jyCOjo2Z+N4+pjbKVPrXhWbpHtYViP9oO5dqte9VM+QI1wYcY
bDCWTWN4jknVFbHF5jyK00jJaK/b5UfgBnp5Xd5PQ2MplJGe90a6Qa8d9G/p
aXHDYsrT/G3p3KMRmV3qggZMSojLy6W2E8OiSZwAQyAlEjYjt2JWEW99bKhx
OCySSC9cYuP8AUFgy8ju3hlJaCevWNMzhEwDGL+DZ5Cto4xpwE8e7U9k46hn
+bYU1+WfZ6ZOmHifzqdVye0qhZIKfcRgHFA2otB6CtdfVhcCEzaGecLKEYMO
Vu/HYdH73fuEqbFZEkKBNIwMZd7aRm6kdY2rjPhgWf72DpcTyraD1bYEyyIu
SCDuvfb2QOF0mAlzaDtw+OwLIQwJJ5Y+xK3wJdFGvEIFspeH8GImYDfU4q1o
0PaLLJe1oYPTRnVabtX+BbcKp1XWZ/nYvqWZPTNGuGtjBHTgeATqmsmycgiY
c0hmHxyMdiirdAUOOqYi60LO30+rpvRSnU9rx+TdMVbh8VAJLQtZgLZDGJgI
6HcNzyjZT6mFkj6rNMkGO2aMun5oQ1HVv+/yjhPaAt+BSSUUNT0RO1eSknYg
DFj/FzW8f8bIs///y+BPb2VMN2KvpyyNvMjIlx4BPK49UROmbzEtEMEfYJwx
Sgzd7m3OG1wtXPNYbzTrjfTtnRFkBdhIeVrGUEis5OSiTXlvUnj/4deRIPLv
cye0wwJ6XlaVPRqzHE6i/fmcXKgEfHvv9vCg03DTIkpwWgJNf/q1hOQbtiHI
Qp20HPre9kCJBlN1+VDw74821IEv3p63NDIMeF/k9P9yNw3QChUjIoJiWz24
UCc+DODLpO5ResEWeHuwBeYRUgPBqetng+TW7BAzxv8r7pUDH6FNjrd4AZez
BgHetYBgdmlN36vESUr2xXJePcl5+FROaFLOOHA/fSmMBC9HnC0LKC9ZnaLQ
rRlvRDLQA18Xj8Yx5aePOyrJOjJc39vKxvPlCdM9h36LjjG+IPTFvFRrgQX4
cBTBUkkiWzjCXQzXO23bCUCb7VDLUJj+VSTLYnFOnJnLz4sGJQdqCz20Pgv3
BSQmc1hTfmHj5ne9kArIBunDu5OdsLAUO61rEGqpoaitS7tpjEKAmWNtLION
ZAylbJC+wJ7l47ddUxi24AzMjR/JErgFJScupnr8hMFjHgo+YRIx1WZ+5jF2
kVpGClVx7oNdtJl0HOxPx5bvhhaK/K3O21f9DmKlymoX0XErDVLsWlVRA40j
ETY3SuiyCkb/l1ejoQCW9+4mYO+WLiUz2zv7ADQl2g/89Stp0tFWoITow2ul
PAvrIiqEBMRSz16cCJUNYWycoUSL3OBL5KF9EtKN8UccGlkbUz4aMw1irwvv
oR7j8Jy3TLZqt8Xdd1BlxorfbbIYM46A+SoBOjIzpAfzKgNNY9OqqfP4tAvH
2/aSIw3mQpw5knWlLQUTgg2l9NdD/H2kASkrXkXStTSjKBhjcvtbNk4xKGRH
D/yIwUjQHJAWd3kvzNHhYr953OQaV+4B+3Ycck9sywNpVmLgTkLCY6HwSZA5
VlZx/b7D/tuHbhg4zDeXI+MZrqEQYPRRcO/kVRy1g4DzTpi7d5qERqHJKHLP
LsDnttR6YE5LTq+neWen+OXeh4qGeSF6uptEZFxgxe7eMiS24BVamfBAKY1O
Tw17eggRD+PJ5PHqSreRdGDm9UgWrXV7ERTkhHmjMuZwMNZ54wXrhpZnfdrZ
b3fWlTQUbD8azNvrxbdVAmSk1fW2HSl41ZlFbnfsynAfwDCz8XV9v82iWucK
2JrUpLHWK6gN3tUHACY/l/davOyCzWlC1Oe7xeKzgBbADxAMiYsY7Imq2J9Y
wbtaTXfPJjBcbynSBBIEJTZV0nCPFQxujLsCeTqqVkYlZu79ejiuRUZHzbQp
nkTPfOGzF3YOC52TiNyMKdTF7VpLJWH+4hZ0qRdOySRm9U5ia1GAyka8lkDM
5c9GGJABZW9F9Rsk4FGFuYc64Cd++kf6K2LvRuhAPHhNa/0Z9McX6rvlzIcq
QZ3BMmOhBti6mInX0f48fGnZSmjE5QxmqWwF0Ye35f2j1xybvFifje9H17gs
UBxu5LwXVf4EL2xrzMCxYRcjx4/sf9LVNLUlh4ITl5ncEpNzoLIOmgJttaS0
KIjvz46xP40OPA7j/o9q+XOcssHuYzn3DmD1yZJ55ZVXL56olh5UesXJiLiG
KEGDDNMHt6rijyj3ffd0FItl0iyzin1Z5R6ICaP3o9VZnn8wPJ3ZYX25nWvJ
ar9S9lziphacDcEjTUbjSdtKNmyxb9GFVlSDodYGSucZHkGN5VL0FP5hjRD6
SejTeHniGMCkSQi1sxJbPRO7jX713nfhE9Yu0zC9YSrcnwqd6g9c7tg7gAfk
qLIQlGo0/WbcujdATb3VdDUqMPA5I2BiW5JK+q6DljTlQG3SttYNvvbj48Nf
90Av8C27MZxQR7ZQLLNx9ptMGB8eHLa9AhEhy0VtdTuX4RTQ1vUIWvKfpPv2
t44rdpI+vZrdC+ODGHnX04t53W3v8mouZj/IjmgZCNdFCEOS5Q2DM6G61cfg
wb3BrgZs6VMR4TRnjD/KG/YzgLxSa31f96WVAtJcZEJDix9IiJHyE2neKZbQ
OFE/dC3UfQth3IRgj1rW+7zB0YsIhwE9Xy+xwiJ8A41exG22Rsr4W/e/t8Ck
vK7GXo71tYC7dn9Hh60vLwScmeTIDqiHoR50KfhwTF+K+F57YDudowzPM+kq
bc6yc1B8XmM1gOjGkm8jNH0mevEBRLT1yIHc7gUws4b20BMx7xLYsku/oC2a
0vWFSi9RhtzSn3aiPbojxDGd2dJXflqqOt+3Znhu0rqVh318ptu3kduqEgaF
T+k8EO18gwDIMWlc01VmX8vra0/25Xb+NCNKbb+N91fROMPMVoBx9zVfCPLd
Z6q4MRlZgVU3Gp6hkH4kPDmJ3U14CZ896N12aGmvD7dnjWckRKYTZyJKr0Ei
Sl5QXZazoogXPxnJ6FGPm+BOd1uHJ6Fexi7pEnyc3e3xs7XUKI7JmYiBWyun
YWxj2uNEj0SlU5UWcq4bxpcpCuQ1ONzBQxmQ/bgbGPlXNatm3/9rJJa6BAGP
tw57DBnDeNptVESR8AeOkR5xHU2NVy/9/+PCwArmp8kJZtFdX39zpBNWub2L
jiAVI2ALrlg3YtvlPLGNem9QEs+KAkG1UQAs3L6AopAZc18CK4Gr6XHge3DY
yonTVZs5XAUq7PlDlyLIoZehAL7IzaCO+Ib5OHRx3fzEEbyQpgsHMy5MseTJ
porfX2ImE5YNpWF6Z97ucceif/NYO/TZYKuDNNKz29u8vU+23871dG8Zox3l
wEzbsJ+woqDjz3nit0DiTpn/DWfg9D2XM9iqCCrs1KZlUPxCMAjYBQqkuDDO
CEMmwcs300qC/7ZpwKaxTx0EaChsYjSUJcxplpR8XEBxOUX78RVrHjr8E5IT
jhyOfp8dvl9HXzauhsEkEzk+4IzpPz0gmLXtVswngv6EjQSC1rfXa8KTuPxc
TA20T7hSlDqtUd47sDPpjdppLZVUk18xpHoI2yXFLyjCgyJf4EPgkwDLmvyL
5XqxMD2uFgnsMtP9mP0LZM+t5yakhQ63EGTtvwPGOKJwc9IMhMe+O1JoxJa4
+gjj8os7S0kyNGYzdLWfZIsLc0AknsrsXNrb3tstbv5+yGFZ0z/LOOuGcIW1
Ywdoa9baE/vVJb9XUqv6WpfRyz94tQzS968zUJvvieS5MgSp+lyjCJcUFz2X
JKM/z0OL9lYsNng92+xUGe4apnTAQRm4oW6n50O1pcGDzGM488QVmsue5jBU
IUhCnoBPSACme4fgKWJ6dpGHJKYTtNRR27kzRZt7VjtUO62kzPO/GtkcFoPv
xdgxB3vT9/V03vRh5L5YyoZPVWluU68Vlcm26m2bfcPdOeHsdQQkjgrQaedm
Pih/q0RkmvTt660ZqwTjORWS6FVGjJVfgQmojK6XP0Y0jlo0Y5YYrA8VTeGX
/vtTqAwgGj7knWgnkty8ZvNs851ocnQxxJ9YG2jhSMhLkGOvxB39W/mS/N0t
pDfV+TfyPtyWEvgyV/2Dc+ESokA2kV+D9ojop8xXAxq53/aqfqO+TlbMV5SV
Tn7ippY1oRm5laaux2XJyAwY2D/radI17TpbFzTogpH6ykyIVRejby9MEf8s
emsKS3l4rjUTb9c16VyFgUzt5/AOTipTHT111cUOXrK4wWtO0h9rI/WRQ0lW
McxOpy1lWiegKUxqieFpABtuxoq+mS3gk5Fpb6Ts7aMXiDActZtWP04pbxo8
x9xCN6fCwLDit9xxiC8O25nGzuhCjLhsoKDtHAYH28pP3aBnh8qC1utPM9Vo
UYArZh9/NdIl8UV2bigstnitXEUc/8fckEKlyUs4vTxtl7yuAqNpi72VxdEe
EaUfqktDymo2fupHF+HBg1zO0kCOieOQS6lgjoy9UwHzhz3t2zw40QkLjhMg
pzmomUMRwHFtqrIg5j5z1fP3iXcojHDRyNzOJcAcvT/up9brzq+mdM6KoTG7
NjiGEkvwnJ7Phud96qubd5KzCxs2t+RTWYp82tkJMakAF1U5KbRcKMSZtXbj
+jx27/2i+K/GHv8p3u4llJJGjuAQpOEUeQOMPdSP7gHHWyCWwzvQmlbTEvo1
zNdzIycipUJjyFKCd811dFGEuO+XmX1GN867kZA8tdi1BO/SV4yajyA0204X
CdJpn0Af7W+3nUWghRf4ZwjcDjyjDLadKEnBcugXv8n4x9jSA0FzPGlB2flz
6uIeRExrrp0doYDg+shknHcWeVqAmzYT3lrqDl0kK83lbsWwJqVYBg2u+oOP
xYKkrBVx3jq43lpWpEwIRIxIIhFHgXxK2+TM58LEg8ku4lDxz/EQ2WLoIkoA
6qGGsqQzpMxBmXbHXZ2d2SaVWXb+Qx2WzuMnhOX+9LLqcWSA+BsyGAXQeBWr
qOnfPBSuE6DkqNFT5Qi9Nb86jf4Y+I600EgIIRg58IueC7JrIZX7180hmqCU
VbxWX58Sd7d4DjS1ezUOTXjFMnLI74DnMJQzT4GC+jlI6jz1X0t0Nz6S4ttK
pQblOAXB3KGscPWfFDcQL26lSSrDZMm3HRCv3OJVc6mpNRZfyMhY7WKaVroQ
TmvEk2bfS0SgpYxgbg/unEwe7apQmMlzIiiUcasqEIJIM7aqtlLSmpCjThkF
r7QPVIjVHrVGbFYPF358Fs+28BeDxi4Sxp/r48EMI+G8KJp1hbjl/abPWO0q
1n58SYOD5r7BxukojSvKF0mfXoDUC27LHPvLT92gu4IezG812bCbNx4lEpos
9piLCTOAr6G37PHzcB4sTckgzHOQFov1QsTTZj7KWd1XZAF6XOvzIpT3hq+l
Z4ZMEJvCmtXwtLAcUDzQX4b6n1mNKavO3C6MZHEYelxnWtVLyWZv5QyQXqut
Xpb3macG9uqlBhc63IWnMUu0kotHTxUnw0Ez8U69R24RbCDUcXBcatxkueld
pGvnztiwFn93y+HZVJyC3h3mJEEv1mr2yPXtcT05keMx4l9bYn6ieBxBt6EI
HaQ9LfIDFWLWbBOE5lZZFapBpT/ir0RnHvZhwp8JkGlkWg5lXaPRMhxOgya1
C86zk/UlvU4HrKo7DTHhwAKQtmAOQDcUVCreagSXg566bnyrGlnZg5tXn15g
ojkf+whxWX01U5fTb5M8ez6uhmkTS51mlMi0PW5ts4MvgNyrcsNrOmBbiqrw
sHTQD9JvxuVwPZ2eoIj+cbr2oU4ZyH1KNXdMafH1kcTjF8jqzKTbjOizeTjB
8fZFTesWnY6hIqxbYYFj8/YWW+wCh9ZJ6D5pu0DqKdI/nhuWzUJlVEH1vaL1
AXDwOSmZMZp3xpQ5yZQVr7wIJuW45Yxz1nSzWZ/RvirxsjGjVroNOVH2GwZV
FlR+lIYUGeGVQDU9lk3baFmqC4tMXeqyHviQwfmOjqlTQXfk7Dfl/u0V/F89
WDMo1piTQOZ5ZdgJzHw6uHctM9SFK4KNo6b8iIPF1GncX/sWscnRx9cI6sVL
/MauI8LoyP2qv3KTXKfD0Pl+U1B/2gapCY6n7kpd29FFAgr64TeA6XGEXMu3
kls0CnQ7fzC1tKOXby/fdmvYbZXMSTQH73hb+ODl4nS5aDsyPk4ySzFApBrl
Fke3kVha5dxy8ut5rapDiE8ArRH36hqHRM9ZhiuN3Mxj6LPh6zmnQhls4yKB
bYjLUupYWlHCj62CucXSMnqoGBy26khbFoGMApbQCMaDXfZU9kKubFGzrvJa
FgEJ5dVH5Nmtkl65JvpWBLUEFC3aK+kJ/p6G43avy3Ka1QZPfjuiG8cbuSKW
B0a6ftDxMOo9dbKLPPYmBiq+y7GGKB/MbeN1KBudA7JpOEEHMv3urp9eEd7S
0upT0TVNEqTc5ODGJo8PZqOCQgdedOcniU7SrLUfHpu3/Mmm0Z4HjsX6oxcg
8p6K9u1FivZ0iiBGuaCO9OhNot2hYzFbG6uYGwx0Ru/LXP+HVw5sBi5xlvCY
HlywcVErH1j2n2tUKodx0nKP7BxBmGaPEKmtmJbx3UmN6mhK/CGu/QcuRpL8
xtwfui9vFJ8lL6hfekh+EdGC/UHdwiABzH986esCl5+c1DMR6C8nJjAlIpYq
syvDClE2AmdqXf+WCZVcKYJSW25mKkjjX9gHFv+I5VnunWPbfxuEs1bMFk3a
/uYv7CKpiXJv/h/cf07i1djZirT7LoXOYz+xdLKSJpnZW58R3DgqrCMA2/xX
e/Uks8Pj43ZlkEKfO6Fm8nWVi2DSB97SzKMPdSyHKo1u0GZe43GU3mfcsjdd
B/PGdsw2lfPIKslJQRblZ1m4PqXhiM5nrxTYiVizWqYVBWFRmolvlDhyjSdG
Tqn9iT05HpHe6y9XpkR4OhTvsflNQDRvKq7/7B/jT752iO09aJeQqq2quFdv
K8IpD7b8HG0PzPebA/Em8/10uVNo36u8AHu7s27DU2GYHvYHrR08tjOCRTLq
OBhFIe3/hCdT9w9Nxu4DQ5UmyZfA9/5r46MU4371+yJC85H8ANogpoYMEspj
JUfq7tZ1E9Wcyvcmbage2KOgcN+w3MsiTFCGrklj4wYQdi8Uu7xV5ZicNAOr
wj5/um81lEmvNDYudLD5n4fzrIRch2VnZlkXx1MYBHZ6whciA7ABpd1J0QsN
CG9JIfilyWf6WQD0dHH8UxG1KK5DFpPxEpanhfnldEmXrv67ZicwFPmgTPiz
UyYiTmJPiZ8tfktieG0z0BAsvxEh3VRcjCu9BriHKo1k0YWFS0laCZINWScK
BGZh3b0XZSLxDOToeU85OrwfQqCx9bU3ZE3tUPpPDCmN0VfCr3oQV5zqeBiv
m+amkkeJuGg9LSKkYdMZN8Eab+Amkw3k4Tr8ZweJqxDWNfHarT6yiFa6ZPPs
1DrOXIm7Bw7xDmUAnSXE8zn4HCwKxiN/Rd6w/8RxtnWpIiG2aYHmSeMDbN4c
zW2BDDnLH/mLEhaPTwTw9h8SMUHgPlpf0D4g8bj7ael0kIDNAaaMl1F3Zzwr
xLtBfhBzR+j1OLx7yXhVTUUf1UQM0jxi4BguBsWuBfOD9UBTyhfAiUjllTSd
8nAPTUZHYSNK2fvomywsbDGpG3HttEgoOCkFXcxgPf03LsUmly9sc0mSxfud
mJxTDYehkwMYHBSUPNeZO24sUK0h2nl+SVeD9iSuU/ijsLJd6HMENIkdBpBx
pEZK5yxiIHdoWBYawDcLlkS8Kmv64DKk+UMYHo/odvo4hOAQB+/i3gnwEQSm
NX5U3YIycmDfg1vuAk5uu7L5DQG0U0ZebJrTDwiSJ+ydX+yJnLWzePwkPDXC
eib67dmhO/cpAhEPjhGMhT6D+Cm8WkmTxGTNpAdi7Uor/be8bz53DV41D5oH
RHZraEjI++Vtd7zvhmWYK9kkEnwjyhE0dyV1RG31gqBQOsY6/szCFPxzORGf
tsJVhEMgBZQkw0i0shOAEBWhRGDlqECgwRVbnOzkacYQdf5mXkCknaCiey6R
xUbrF4yDbx9J5tX8RcrZowet3cVoSOKuOQB1qRzbokqWrkHOzQnqTdfWOJD9
35ud/mlRGBHxqhePkRyjpy7Eb62SxyU6pb5NZkpSaKpLup5Z8KjhnkHWHc0F
pgfIxV3l72GELvTboGgpCL7jQBOXf6FAv7QPI1de34Sp2u/dsTqyUvnarQAY
qFshsJ9Q+mepTDrMFrafRTBbgEAFY3OSQqxuNS1g1Hkrn+csakvLvgzZa+8p
d34hUbFUkd9bBK5pt+iAgzibFWPW9hfKAv6Ps6Drq+u/MxgZg1PJbX6Qnp0v
hZfY/k87ivq9MwnzvdvvSmFpCBVg8/J83+8K1sJz6SbPIS4lpQeg2gXBeXJJ
bLogY/wxUrhprE7bfKrpNuKL/4bNr3/iWrL4u3tjb6xrZJPBdnltjxWpLLYs
k70f7/MLps0KUNX3J27+JGaIHavDSCJur/LKcsXbBwuOSpgT+yzegAv5pgrR
/upgLjIaVoj0Xv4SFixbcHAG4RiqHDdpsNkoxWM77J3aZhWumdW7wy/ruZfT
+VNJb5SmV8LeqD9oLAeC0kwMLPt2Sd5Ep4yniYB2LxJRSr6Z2PGazooLNn8n
1LBElVHwg2ws+aFbi90uH+LDOcZbKPANBUSF7lw8AZ5rbUOVnhX/D/vQMJbz
G7f6sk9OGAeYZ+WNO5qkiYiZy3eEXVXM+c0DjH+43I7212uTmJjWF1EohuTY
PbBELzyI7DC8B7jUbjPYQv9E+g09RtRN42amlBwIMwjQhYWNZ+zhza0LEHKS
wdioGPRYqF5iwfeJe6JiJycE7OxkEELZKY9QLyOnMR3yzvugdt5hEqsA3PRa
kd3/W1u4Fd0WUWH7R3ZdpAe+86qT+L8zAV5aJ/chVh4oLZaGct49c+VIiRzU
Izr/xZF/6Ndv+dtaKLKqh3ZgjHB+B8iNwVCTS1HG/MgPsSZhl7dtLB8wuwsX
1Kte+MbpKry80p808YLSXqvI+k4MPknqbhGS+8ug4bdhLMI5/ZBlaw7vY7rk
jBO+Y5VsTTIwUM5ZQoG/vLSpm47DdeNDyVDJp3/fezDT+B6DTo/i08POLq7f
iSexzcVIIEmhv9oKxtYcwQ6ShWsFmN1qUivc/qgTDyQ/WZjU/Ob65TAufPsW
3TBvotNIE/6b2wlwEZTO7tDC9I1XljhUEmFsh5go4+OtuZ3aemcIOPO4JZxI
7Hh/S1WQPfTOf7TG3azGXd10wME6hOVW/J3yqkuTv4EwPQPVktkiJRfKMrOu
OBiU+LmVGj9zz/R2oNVIlGrBzLpB+ngYcHJDsS/CymH3Vq2/D86vc5rlTW58
wwUEJtWt71ahAlsZkK3UkjMIldYjWtLa2CaUuwpE5mUPQeAwEwpUKfPQN9jf
49FXkWBhhMmbNe4YxJxR74Q7Oa863TvMzrY4FzoHmsFDGROIUReaC0FGOWix
qdxVdEH/+wXvpc6qUkV2Uc1zTwNuf5QeFm4YpzlT/s+F8IYRHCLipkj9gxFV
4ao65UezhLia/ocvCgnBDz6Id5HwLm2scr7XXu1ooR/v+3ogOXpEQu/iG9uA
lyX1wolv9btYWS5m3AjljMHwFTq3RxW5V8WFw6BrVwUaPnEA0+v3ofIhJYjy
thR+ZuSwCQNSgbHSdP/ri1HI34tBsJGwPYS1baIFfmO0dJ/B+0dOjoPIdW/3
uFBpIlG6PvwjzlOU9t0D5XU4g0GJeGLCVHxp5w54B6Um5WNIDPF97yTlyZrd
5v37nh/G63IEd+o41d1mU5QGu955uL/uvjUVtyeOw9cWioHR4IDR/Svn/tpp
VwbWxEKWUhj1A2eYtpwp4mzR9sEKpyF48eMs/SRv3Un0TOlEWi6yWcdE6mHK
v79jkpK3QJy8hFj1JTMZDOHvrB/tgc1il4+oy6UTxGvUtiynaQYA2+i0ZrGC
xEYy6Z49PXolPZ99F8sibjsNdc2q7EQuqbb8fcp7Fs6JZUOB2gdlpnwECkY6
6ae09Cg0AChmQ4lbIm3Gc6JYv6gk+OVVRHVZdiPodsjsu04AbPs+OCzA69lN
iaQyFu4h3Gtlze8FtUYb0QLaxHkwolhikTk4dQmfseA5772arOPwLoNDAWxe
zw0tC306u9jZnlsViljN1gea1h+4WZX+s5HahYAk1ll14cOrLaRBZWYN1t+W
+CLv9zMtpaIp8fQ0fQ3zW8JQoI+Yw1uJ/VhLpEKG671k9xYhdm6E0pGqzeyI
FHUze+zO9rIDep0MTkw8CSFe/dpPRXw+mSdDwWU5XCG5+SSxrw3XwxIZ8DKz
+liT/34ThW1dci9nkNB8mA8YxVk3FYxeSzEuyZgoOLc2Z891cHSosOog9rux
1Rts3ljp8ftRDeKY6EGyNOCkyfAiL93WyPiqiDnhFaE2IMm9JQEUrHqLgcNU
vU7K9d69ypxcd7NCuwJerzMJ5HroFqITAJikqiaey+c9VVRhV6pnrTMA1v6D
pkNoG8kSgcj1ZO3/5/n1ovfchw5b1PGJFCFUkOkZIK9SRqAzbFT0cyXwSn4w
NDT/tnGfo+wY6G4In4qrbaC5KhRIEvWBPGfxI5X/0+NgqP2aLATrwb6P/ZHv
vzHcqLvnDLT8kY+48hywTJc1f5HMufo+5Jg0NwhAWqwj7/qY+ehd+YKoPk3Z
IP6FlQWFS55UEwAc5nMZfWizjlSp7u3aQvsw6XKjhcp8fpSziK50fRFgx5Kz
4Ot/pf6aWCzoTQuEK4gOaUDH54TvpDwUAd7Wogit7wBFvLRRX/SmtcDRWJYj
qZm/fLR3W/DuXvKF5focOnVlt+H+38HV2juLtsXTqwkrE7MQXSAUT64w42Bs
4Tpu+1GPt3Ay27w0BpXQvy9QWd41GzKwgVkuDYg8fT30igP2fFtaosi0t+8B
y09VLKUhGN5y5agru4JEqI8Z7hso5TMpe0ELC1bA2UjbiqxZ1KHZuz9s0zUG
Q8r7+Y1zLtUkZQXUJc+naTCzHcJ2sM01uoNo4Lljj6zU2ggE+yxs/t6ARP1V
65fZLBFYquzV9jxT6sKtIqyshHgXPHhshJcUr5l38sYj0ntOlkygQSdOK7VT
6NGgyVDW0dTIkgKYFnkN8O6hSJsJrq23oAEbtl2jQwGLEOptoJ1PfaH0eB8w
Xz5OjPWkSfoyT/LM7Xqn2A8F1xC2Uc5H1Xw7tWHL8Ujzt9t03OVtwoPn2vkX
x9r+L/Ls0XJC32NNPIOVmT7Kp4u1w+uH9vs6ynMP5EPS9KtOzkUmXCeiKmt8
MOcChNsSnCSxKUNcDCpEJMIbNXP03x/nRpYDfujRuzIC+vvjOt1PNM0c290X
qv7+ONlhGu7eiB/IyFJdnFslLIgU5suHgTJr6tn3WD58Buv9ewwLEtMrhq/T
G7ixCUMnBlhcpnSYgToOEBUEW8T3X/EVaOtrs7VaNFxnrzUxvgo0os4Ja48o
5VvllyYyewupum8OMVrpB7Cwk189RNI6yy3yhCBOifYvCv3eJm1Zf7I0ps+Y
cyqlH/6QNagG3JUpkutGdhbYeEPqbxIUT9FdsIhC4kuj5xSdD7kHuMaTHOB4
GuP4EAFcvMZvElJOp5btzVA5GP5OwzWKiHDgoT6vyCmM08S2ZrNzqigL3Bvo
DGYglCq2pb7ZTMZW6801e+XQ18XUDgLZZGPuSCzhwzEtsidDsYvRdLw1i9bD
PagPxcBh+tA18T0ipvj9ZmXQPBoLFgWbVLOtnYHGtRYcI0VGFUtPulCEQWYV
v+XD0GEsOD8U6hO1NeArRwEdUHOBn6DHsxnvarF8lKDZZzI01+kTBrOqqsyD
CNjcLSuJBSeqiJfvFPG41rmbRBmcLfR5vdFGUunaf7tckx9iisDZU1xtsy0f
rpNbHo1LGsnuV2xpy8j9bZuY/1+er7otl8t8XCSupDzN7lq3ixAqHDldy7UV
h0/VcmH4PN/TeLtutU/QR1yPG5T9Nu44Y6UhIKk8y/r/Dus3Xf86M/Adgmt4
ZaSE9JYpMGCUIxO96UCOqvKqlkvj8KJpTNadWDyhs20RXOp+u5ifSfq0vovR
9odHRqXa5LrX5+wsWKIdis0Frlqk1+WiJSdxxzI99NQlOGZE5exVKDr9az0r
qihhFiHgTQIJFnPOS2FeDmw4k2uwX9yg+rNFHr5MWC0IRU1a4JI/mR549gH8
Ehu8geJ9jnlKl0xgpMygkrcGagH22VnxaLsutJOHL45BArYQjbvcKA97zELm
jEVwV6VjJp0qkZ+tiV7Ke+ShJ5OG0LarHXkKXfQVmuBWU8TOdSMgRpfdSEYw
nL+Sq97SFfBOoYahKXuNc4W75FgbLfkLxbZCc5/AYnAMV6HQKn+mRnMfR9qo
2Ni9miAJF58e44yJcXWo+HEW8+qinWRRqrxuFXJvQaVGCyJNVhSL3aiAPjDh
zOJO5T5w9Zmx3dHfkjZB8lZC+kKX6SoLNc2Z1zxN5WMskmcM/IY9tPL3j8xX
BwJ7Rffx8qS8oFTD99XSAlPhlTzAzN84OccoFFgenBXOFMMNZ2r8GyuDDN6d
19jYGu1OgRAUO51wgh1FCALGNEBvyN0Afy4YG1zAqhVaRiKb0Aq8mUCUJ1uo
WbwChzbk8pOwZFB/v3PM+Esxzx0Sk0OgdQ3EL18vj8GDvUXC8kI952Hc760t
xBwCd48x/kEI4rHZ05ka/feVRFOba4vORdVdEYbewvY5A7Z/uPGtjXiAn7l9
M7FUAeORER1LBCExeAUyTHH/zOGoy1ue2Q6LJRG3N8wr5m/giD8+zTwyAepR
u9S3E33riV9D90g01JizEvVLYJ9z9DckADDPOa2poGyO4tNHATUdPErVSJrq
O9c580XrP7BQ3FL9THz70ltXYeQeNFsOlT4229b0ajwb7SlCm+8NmlmBZY+w
jRjiwIjjfIDqSc+sp6AbtPrZGENLCj2zdvYf03UDXFaahAn9k4M/TWDfWeEW
8UyLLvV6WJ6rvyqL8znGqcwfqZBBe3tUOwVvAvsFc5OMkNWD5OpdUlJRQi7b
6YvkuI1AHUZv2rKVKChimgvsKPaCnRULwqU7xeTkCM4R+5Q+CBxS8LHzdqYu
XDwk5Y0gH2fdB3nbr3nDOpKXBC8X3uIHnLUBc1fWq8T0KgMawRC+m49Sgzs7
/pbPhzo2ZOkLz+UBc5paq8jHwqXrdubp+9IrbE3+VzizPsfmMMK/eFZ0j6u3
kkhSxPTylkVPmkhuXPb8L8wtqHpBznHwo9yb3mHYtHWEZe7ra1djLOQDC54A
+n9QeKT1UN6NswUCv1GZzYgcTU9a96xKNEnzQZ6ALdIEjIQC3ls+TyyyfN0i
cEORV2U0q0DM+cDtevhwC2ZR1O8ReaTWvkQoMb5tASLu/sI89TjoPQPUFmTo
g2LZ086eA9CVHcKnAmmTLuREKcmJXb4jFIt3BVsXvZ/W6pcS27iX7NRCmtBG
ivKTXz4IPdvy1PAi4HpoIbafeEjvzaFZzC2PwH7xDRkhtEtMaqF3GiZSuSQ3
W/IQfCJ+u7neftyO4/RhhodRSR/PrtmVi/IQ58aWLN+0bSyJxEEf1xw0gS85
syflZly5iBmkLWPDnvrKEymgiitz6OZoiPg13mGio1aqgrMYaGpPc7UURenz
Z+dac9GbvF2rDt2h+p0Ocn3AI4B6FPsTA8OKP1GnAE3pqx2aCI66T2Q4sXrb
NyKQaQenqmUaGAowWFpxkkQ+dyPB1SMOBFy4elcNVT+to+HhBIoMa0t68YWA
CqrkH4tvLixHEiWH5ycIFfGsefPhiITvTp4PAUiF36B59X47VYSylPrZl7r0
CFgvv3AgWLrqoykv7fJvF8gL4tSiZZDAR3G3N+ix6S7Zge8Za878kCKA7rh7
cH73XqSN//NjV040eJGNEVtkeu3RFu5EaSAvI8m6uBNaa3rmcB/9CpjzOxbM
XfgwVZbOiCjz/Ccj+hrGt2RMFmvoCcCgCrcnjKx2OhuXlfkmnix5S6hzALUO
1kulHgZ3YN9K4iG+7aCuHmIQv2NX+LbYW5jogACFO8N7kk9EDh7b0fQMPqwZ
ZqfNUM3w1pt/8RPUeqKhNY/303/yO6u7TVZyVbfez6CCY9H4I7GTX607b/p0
n+dbUmE9ifS3FCteg0tjXyFBSJl6m4wCSWjkcr3V4mViWG91MkUxSRoLuNXa
hqbXwfE/RSDIcdMr5GgBCnKCsCe+R1m5Jvl8oYHzyFfWgZGHWS5Ld96+q8NN
j0k3UBm87RhGWo01aW2ujRR6MQwbgxv6zB9vWvCEYYoMnQf/huCf5ATxYskG
PAgviRekfuQL6TZ8HesZKkKXzk9dTaxxoxG7Mv7nsI1Gi6oEeBrH9x8J0I8M
P9DYMZy3L4V7MqzMNivt3cjATLZwmndCtyuwyk2Jr1WnQ0RETlKXWDKn72re
jSXh8fAUvbqb1VOO4PAI94d2mVxCP6Kxk9igjZSGJH8m9HMhfxy8ZD6NdLTF
XhwsOEsE2o/XuJsBuYcoWhdZ+FQl/DfCFOa4myNv0Av6F1/qabp3PAZk+cH+
jcTXC8LahevlZTil1IssMeakWWrJqmaStKV4NQqMXoENjSMJEygBflN816tY
UFS4sTyDqK5RuAizdX4ja7Y+hEYa4N3w+bWh9oo8W182khFZC3+/Z8eYEHqF
VWKK3jcl4iWdhAuUF0PCOmoF5mIRTTfsmuAjqD88pVdiozip4Fvm3bBikNnp
cOrYq5+sWp8yIyYbVclU4aUPdIa40QyjUm5nh8iqjifhUJ0tO1WJyX+ROVmZ
TjKkMruqWP+779EwFOupSmxzwUnlYRT/ivQod6ylJOaam5nDJFH1QJXNCcs3
XtYHkwjFyF4f5LfphL2HPgjhp3UaHUIey8CS/UsuZ4BOCiWFQyAvK+Otgudn
82wmji72XX78YsxaooVT2aHb5ERZn7Ok2nsINDuQsaqA55opOidlEuCtSpfH
wPRrWXVhrKN3UMTBZhJQ3F407hPGC/LJWI5ap9/SIiWEcaHIavm/1RwlqCk/
iXKrLfKVgdV7ONYrq9SnWFFJZ5QDIRdFZ4R3naKXEPA45aAxVhzaUJdBg/IL
n7INeLrRO4/c4mUUkjbiDtnd44M5kdcexxsWt0W6nI01QaShLSqI9p3T4N3o
q12JD3ZNQ3UYYgvNU96pB9I1JD9yGJz2Xs4EBnl7v1T3oFkdcJ9V72PRgbGH
vL+cir6/YeaTUIcvhnou7RUdzShsYgXCrDiYVTHnBpO30hHGBhTru3dtQcuU
H4XP16E1pea2xDehtV5BviZTofFA0oXMGzW/FL7EweWGOeQ/OvXl4IQUENmC
stGunTtxK+wnp/IwKBXOizlJK3SUzW6axlA9Zg4voEswfptWhRQHRtcqq/h5
sthz3vWLQavgWZmSA6KDFLRSN314LrCdqlnvT4OqpRtSmsTZXUTzkx64RsSE
tCb80ZEjylwed99HjLSsQoolO5eep/ra477EnQ69U7Q65AQodh2voO2qS3CJ
hfyjBgUXd65W9jLomQoh5apeDj1u1t0vEPpNQwyOL1ske07qUChgfuRo/zKR
d+gQ/FqK9PZRw857XoGufb4wm//eOENqvvqW7XOG6z6dENL4bYdpz8d8FJrC
2pKzrBBVC1+keLrXsJwGldG1AaZXLmhAr7MqazneMdiginnUxSpkAn6hsAGQ
jMpF29++EgcKObANOTdiETVuhcFFP7QiNllPIrFQSGod48yaC90IPTTTZnD6
gZod3eHg8j8PlMroQkL2ZzJsFCywzsa5q2XgqkOwayaSsn/zUb8JNAzYW8um
1yen/I7yR4Z6mRg9GQ9c4+SPG5nrPoIECXwMjtRSzXka4/7vHCjkEmfK6zTY
yMFd2MKgbtbIq1tuuNI4wdSu9+Ci4zqMtFjMj9Kx0OEeW6fHV9xKFQt28mtk
ApOVzyw+kqgXaDtWFAG1w95/E5tAmWSxIlI/cZuo/uYIGDBmdANAYp8XJruS
vMd+a69jWQrBvvuzww30dlGSGvH7mRSMm/k8deYM0H7VG+C2TH6ThshWdXXH
oYzSYZSKASdLxowwI5gzwUSWAViXHxcRLGi1a331MdYcXTcqFXDry+e3oShX
4c+cSWKZb2N4CN8LooCgTOn8+R9JTydw07s4hcI+hcwaazmB+yZqUsOR2/W5
x/ak5gG/WwNqgt3JU+o4iYKUX5kaLzXZWCBOlN5t/XZ8b+Iej5IreQJxpmYq
yki0j/SwxtQMwXWnxBwifZHXqNqw4sSjR3SklypBBwee1a1obV0JCK/QURHM
Am2FwB+7mxprxcvaLG5zlzoWOgfKU1W/KX91G8H0KjHFc/LeERqv/RHDJ/CJ
st/Qu2tQ/dwwem/m80lDr+UuzlCRFw/wzIdaNBO915387VBnquSA0oPAa8Rl
KwEE+utOkWVIHEfoY7pMCOQighl/wi02ZD2gGfHHD6N9bN9Fn30gmOxOsC50
duGUjcDVmE3+etBTsSkxx0015XMLJfJNPD/ZUJTWY3TAr32CujiDmTYCjH9V
oUnZR5fwKaSDBY0b9OWVdbcP1Hwjg6sMGIlm10DyxGlYV9ojlUQXM9Kbmk16
7Lluq04IgXvVmQ+javeSf/MwSTe+gL5ytPGEB8Mb67h9cda1hq0GLpfCJD7b
uFfcj74TVqZnu1082WtR2gJscbihTe/vzu7iWHhNw1/LxthdH0yH4GFy83HR
PdkCcYbamwbUnN3oxMrIg642OKqi+XuyXReN1mVVcSqAIHpVoFhl0gSMEpsK
ck60FQ5sqjLED9Gd1RG027YaHocnloBgnG4VynSRlxo1ppzYsls6eWpR7T28
05yW1qTCqGSsuN+a1Coe/g9N33+WCG1ZQb/wBDgvZxUHiX3vF3aLfYZtHB6C
EiBxpblhGZoLKCpenbO6NvItqCwLTeHfKomsSbPCRvm4+IOmzuZQVsw6Zcof
pyTxsRtRcKJaUkBsmtOAUsJU2E1q5sRZlFlLW8CcA8Qa1iYTAk5cRIQbjxZR
GLgB7S6f5NfH8fthrv3idC5hIV/ODLxj6Gtm++LyPMdRnUdKU4weweIWc6Z2
V60QHn60jWdWghwc9Ji7lD9APZrTAy14nO6VcX6oUdwu40d6V1+CkPnmABRG
ruCxsyhmVEGxgAvC0uXtfOCwOCefqY+yK/BtXm73RJVsn+FPJUlqnyMFSh63
nMSJf2XDT9xuNmTIKJq71clNdGXwHwA3ogpEISrkA1DnzFLxQARYwjOYVrym
YdLNZDpYtF173SguM+eYy57Jd7XP+q3/gChRV2cQajEIgKrzEF0uLwnDBW8f
OtAR5/F0SMTBdlbP4+xZ2U/+gCo234xl8g41VCm+U9YohbmOg4/4KsvaRKC6
REAHR/nUpcSHlwvULyYRhRmFPyovZXu+aP5tAW+noMp+2ORe3wEmnd53mD++
xdgQXyxz0W6TiOl2IJ9c/ZqJjriQQAP+z0PWpdfRL2uA3MRjCn/6TgimAYtK
oU5dHT1b3sclC+MQRTRFtywROMidhUuN3rXt7+0k0m55WKoqGLXKCT9g/gvJ
0rd/FhtPEP1wLB6093oa8rJoGmrRd0Hqt6Al3E2IYTNeXOQgR/nxOFyDZm2f
tNUo491zNN1sYz1tLZBAMuxxUiK+IMkGIFfDg8IMZPFqnwg6kK56HC/+QByS
HveNVbAKp+ZR3XxgZA9InUMNYxrD5RVqViR3EaBXteVXgW4WTarADCNjis3J
iU+QIsXEijFGSjggo/cGhcIMEzV7qjDQSYnwC0QFOt7VCI2/gi06SV5iSHgJ
pAHBD7EWielSjzl+vx8pA5RNiKEkt5yFh6DL3H/ME2V1Aqy99mzluFKq9Ggu
ioQmj/EWayOd7wC9HR06od2efrTQrzuazJOv6IO7PrKWiY4mYLzOUGbRxLTJ
b3XMdnzllvBbVgWPg68gXCz+BWFgvx98ueiiA18MmBa+Hjtord9GsIMT2/E+
8Q104l0f63hl5g4fxeJ2E/NkCHg1wnnPO1h77ixrPEH39Ayt1DX0C9BHEoff
aATCh/p+ekLQI2UcV9bKxohjjl7A1RAsc5zYHH6FPXvzMFP4lwD0HaPRe47t
J/QTuRTdg7jbs3zh2MJNutZs2VBPuYB8F9lfa3ISU/lcswH81gIKOib8lxz6
DECQzag5OIqdbf0wNmSmW67DyBEVysWqLmfVdAJl/ZXfF1pZ2b0GX2XhEByN
xuOAwA+8AdXOf02ru/zjaWm5s/CozG4jIenFj9yeKdswNbH9n3OeyBb8MldY
fPLeoal58TCufVkqoHlgi9qrrg5O4OzO2ixjB2TpN5PKbF+ltgwBw6yH4Ngk
LhN1e852bRXtET5fLhT/XbFjapi39eP5mlsaqXv95RO/Sz3Z6UP1aYRoNfIw
jghfo2lcKhlS6erIaG7yhqLh6ADwJR6ostuRiMO3gift8qgenH3RCBOhdR+/
vk3oMov1NNizh4Vzj6m0TL7wP4JX2iO+YRns4LU0jY6BOQefSNeYXScWeUVE
7Iae9ZIUeMvqp8xNBiWlUR++NmJfRREVBUx8/tTAbePWMFtCx3zkxrMomvkf
MyJU2T4MghQePLNbYLZ4gKEYzf66dBrP2WkBMwppIaY2OwnNkpVBsSHp0cNr
PivNMDaqxlnbyiYHtj1yMIgNHEHPVQPtG/Q0Mbc64eErmceQNs7tvUIFGUL3
E0yrOtz3fqeAF4w4Hbx+yMqCk7cVq/8tp2FJGDZSVbDUi5o7JvehY91cP9gP
KA2nSlRdeIABSNXoVwUjAzMcjTenmGvA7twVWpUcZJSelHOTzEpbPT/p0B4+
K2vPkn5kJr08snHzkeMZQf8V+jq+GkkzkSsKAQVDmJ1HL0Z6+NYYQ64SB/4g
LPz/7gZYkYl2o9vBKkTmx2vcnVqTOSyIyoXeDULwvoJqLgYeI66MNHvrogpK
/of4yg/buTrYPxR9e+PxweaGcHAiAGQQNTI4m6r/J2kaaT+XRHdWRnXeiFXX
YLiNMvUZQ4r6A4SRfa0YR8iHkX7MYM4vaa6+Ec8Vx/ioRzu2OJvge3Z5R4Yi
qbDHpCQVm5kDIdGflGUwT8lxmXr54NIG2wbRsEOF2pxB896wJ59nSH8s3KQD
pXqVK0Mrb0nt4Gji9slPnZWxGF6CBkael5/0zhUjGlTfzNjq0zblDen7jLNO
ELze2GiRlcqHlloOSTXgvzIVa8os95VuM1UY3zw8aq8yGfMFu94Da7/vGT1n
wwVeiCOd4fT9rbw7ewpUKqrPgHoXI8pMrMrXIvasc8sTop55mIa+/Y24UWq5
Q4iCYu2suSXBJbo2q6OO4OuuE4pMymFlH4unCFmWpDUWkOXfvDZ8e/Z47Z4k
78ODgzvKTqhxYPieF2MkJm23yvnLfLvRtpWcWTV1ZtlN5OuPRo7l0Y/uekyb
Hpj5K7OFjfSOtaadUlnaQ1MLd5MGilv1FGPz3TR3iaoNv/I3H6TaZ46fUhaa
9aai1PTCfyDs5USmspgo+jr1zQrLMuRELWkIKi/NLFI7yjtaipYqA8j+cjho
Vb8w33pBhrdPELyhj2Kf7rC46mp+5r37qVzT8liHKIVstSGzscWOHaniusbc
qR/tc8T1EWpnW0sSBThVWpCXD30ohhoX7NnV2FKFaEuH+w6FTjJqvIqihefg
lgjTekE8Wwj4oiz9ZKPgyQzh/pdIOk7lkxaC1QWiQ1ud4ubOa1X4TCMpztT8
Y13zFWk1mwqQkcPYb4lMsnwACE+JkwhDLRBjhyYoWOItOvmGs1NsCwKiVBNp
u/v7UfsWFwo3Wf4bLOyVvjasZ2jpNgKUd1noY8qCj9lbP68U1TX0H+sOLFE9
8RnlsoK7vvAXeS5TCHAxETyyUs/3GaH5J4aFRoc/2vzWi0IIg5gQnLL+ztlq
uXiXZw9WDTWt48gbvLRLZbU40JFzQmzNuKIuMwudGBYvmqdls5lcayyilhch
Xes7OubHUxglQQcRravFZuFCL5ZKNcH+9DkSIMQ9e+kv1XFoX6quet0MaHu6
BUFZjijoFAyunoyXkc1rgog14LveiCTU5lRckpr55o+MImyUVUruf5D/kiOB
wBn5HU/WpPUF9l7H8A0po9zSkgFER5VYpOGYi1Iehssat3d0kJOnhyPSnbt2
E4TX6sBm/R2uR9Nj7GYB63q/1QQBDh8oLd0latSMmuoPHj+BlImDJo2ZOgJ9
wK14ksWqmlMUmko6l8j5KnquEKosIcH5w7cKyC8DIPLwKwGeAiqbj0bX7pyr
2inLxor/DZGpncfZGUveli6yyuT2TNistcEsbMIGLpGA3s9/WQqLgOstoZqZ
h11ieS3NYIQL4nWSxtmP3mzAJPvNfehWwQfMbxLJRiDDmUiEHEyLuSUiht0r
Kf016++579i9oRYyFI1idn8pi44e15atOdr940UvAxkX6JxvIxvCkFT9EzH7
RIDC1sFT3TuMFL8L3FCK7N9QcFpGQ2sWq6f5EfyrlxnsZatLxu6cZAnTM29P
cjlEfjPK6lc2AZasaWspG6xFu0kOgqCbnhjrffEzM868GujEfQquCiRVSB36
K8xv9Iy99A7PDykXVM7I+B6ou8ebDRO0adXr5/klYLOjwCqy3g5/Sfpe83zX
Istr7zbkqAt2VufgrmpuiMjudg58ZzkSwLFJkRm7p2O4FztfoZ1t8Z+Tz2kp
pSF+o0uewK1JbIvD2HL6Qg+Y410AMmi7KAFyiLHTlmKP0NaoJ81NzM6L5yj1
Ii/BMkkvMUUycgyzf3DgJEScBx5/zrGyl7SwX5BhyMfQ1nRj8/TIRc2InD00
qyqSJfYrGq6d4xqK+3q3qWAwBOGKymlq9tXNS8f0OfBz5QS8dWiMLtSrT96t
ZpAKDFSxbmu846fEWNJHDTbj6lY4pe/6Tb+dRWA8vDWHVjxYoAyu7WuCjHMU
QhOurYWu0s5sGoLlG4Kkh43jPBn7NHnREfk9S5tjOTVgahehHkfhj/cRcROP
V9aLz5pMNYK665WykipnU0qjWSQtDRZtMXNQjh/FWHvppa0KBcujufmgsbkp
E+6PCqqW7S4OXMNzPcDP3umyLRH5m5z72JZXwH5nwCytsXkpRuHZdKFE7PWK
OZVFoXxpztq6uRyJp9tEdbNFEdrZdiJQfFL/LEEI27zyqZRkPZAfb1V7Cjp1
zeCDRtziegqg4c4wY55Goj7JB1ctMyYDhjdSYV0+lKKXBmeBmhP1Gz5SPvLz
Sc9OSwZT6ksCAtD34rNiF8ORDc89+HVSa74hxztlij0TkpyLhTFgStPzsCId
CKUqjK1MCzwYdI1jVI7NYns8S9WpasTOzEPnE6kZXEoLksOJpK1URNibE/ni
BEJv7KhGs7fKLqoO4haBt2WwY2UvzDWqvD47zpjaChmo7ytoJhia+9brXWz1
tTZfQ7Vl3DJuXc2Qq0spgw9O6qVAo6nz6hnQ69jdE1mTsj1CP7TcA+C9/4lc
Xasto/9sBPOxiILjtKQISl0xKFPEUVlZIwVmbb2kYLXdr3SU8pan5W7Unf7+
1jDW7Y5O7J4kCn4frdPXEGkBF+Pa2tVIswOyUtVvm6iFGTGhdvJIb688dlzu
xiVECX6ChaVxPoc1Y29ENsM5GJFVZq8nMlIOZKwRgvbzy8xCvuIVD9mJN6DX
8r6ktfB33aWdo/RabOBSo9hdT+p03DRCYU4Qj4r2FycjAHA3QTIfSrTaoXcN
5HU/8m6d9BaZp+VvpFHc3eVtLSLJnz7lQmagTCUIzLLABF8xeePFFPZHRyCB
RtNvOvUJbXMRDbC5aAavMw5NTu83FSCsvWrXQFNiDwEjQaE+QRmnZr2YsZQs
pR3SUUHgGRxFQS6p5bxFon5xGFyoO+n5+w+ofJsBs/JlklrJJ5rX45Vrhhys
nqcdlBc9W2k/MX3leoP/CvWOE9sizYSTTEgcUrIVCMaoIECfdcAEn9HOqhhy
DYPLGgU+hQHCWMEtzPdGxVcAZmLabLKYOr2hkb3roYzRKPkpfXnuRX/xSVR2
FTW6PFI6drmhfGAbtppbZ1TUqTbHrFGoOsqyiAWHvE+uG3xi6ezpGgnhpTrl
vJTabaXr7lSYLy08zfiSsnxP3bQHYlgJ/VUjQHFOLugQhey70MWBEHZ5MfIe
OCpgy21YGC9I/9bxxJXdBbUNfs8v4PokjG7o2i520atmWNlpRVig2VZCun9H
hwdTsIFfXkwHWXXm7TBKJXS7hgk9xzR91hFyWm1LWtGTWKdq1BPf1R7zdAXK
ht3zbCjnQE0jVl3dmKJnjIezx4vjNA1hRLXW4H6fEYwwkcM6Eq0poUMMnSfS
qfgWz56LgLn8YO3VZDCjY7+bULgEZ0bKnaMWeYdtKsYn19duF6XnzffJNq3Q
PapsPKQgelKn7F4eGM/EbHoNV1q2Sv3LXPrPyq0xQcYxjE/HZGuRxtW9edST
BM0+Sn2S3H9j0T21ismParh6HHRRxrm6HHmPu5PsqzYtJJQAAArgjuj9z4am
PP4KHQqW+OWBPzUL4sNcWs+RwbuUL5/ztGswlTGPEdu6fiPlE63YAKnPWtyI
bjOqz3dzE0RSZvxZU13S7IAogfr1boxJgDLqXD2tPRgBXREClrCPsrB1nSLc
EPNo6qTF35DUVNfIfbDXBC1F7eINhwoKZQcCdO2YUxo6rvoNykOWcJONx4fh
kPRChyqaCKVxZKkX4f/UAO01FNeRoR5ovL0oA++oQUzTi2T3eG0aDK7A10LW
JhX1LBIIlnMGYXawpjmT0B+KvQAk7mLQNKC85zSdx2s/NhtHRs71tQ5yy3Ak
ny/kx3/dKFOg8SRjSmR8SleqTNdf9QNxovap+lSdwxQYCD88RRpU9TEY6pnc
14z4wvJj2L5b7Df/5foryGzro1d41T5kU8SZBzj9sFlMQGHnu2tkegVRtJag
+k37nGLJP2UBvKE0F8+kdGGxzD4/pFcnXy79Xq56TAIhcb2wozKtwBslJ+X7
UY1nNEeRmECQJKRDuqOimTSjZFsNlPMn4puHNEqjN8v2o76rEd7aJ2hqincV
A2olxygM6/QqRD0yamwjHAGHHE19tUeRHRFG+WF7KoMlmHCaRZyoC1dourwY
H+bXiQZkWWmPzsHYS4w3UqDvlAFHUKOpL8FpVRrSs6Ap+WvmKe61P68x3BwQ
ncrmKwUqcyYSFtV9xT+HUawaYwbLtEXWWHjtPkBkT3n2U/Dn/5RL/cJNcu7n
VxRA17oHipSQYhNmSsb1JztUyzKoTtACvmNEiZZesitcpp26DWVoJGdbdSPZ
MTdy8H8YsONNv1YzQF83LpM6pt50Bad41cxQPKJTujs+fbpoayHXfsYWEux8
NjloaVNSsXDMyMxCep+5ShjbpfNYvVSpNPWjpg1JXl4AUJ5EFxHiecJ28/1j
8vE3TU/DUZVNekcBbY4ytjO0DAZK9Mrzuq51V6rMRyWyzA0M3CYHUMwi2dwf
VQPUP/ew9doZsiY8rfGehLT6v/f345gEOtqHiLSag4Edi93ghpYsfdI+s74y
YeCw/mCvTd66xpDHeK2Qkvvy5xFCGpknxUIGSLXyp+IOkMfyQhOw5zzzdw29
NYXEgG/zRY6x31PXlZn+NR1JobPyis0SDt0mpIVF2TjUBcnxy4thlT5l0gHt
P1v1cLJ0xNr3tzfNiORDB0dRJ4Z8cY5miigG/3hCJYK7UwwdTkygzxRptIhj
7FGziS8smiNAjC4s5bP4ZX1TODWd/3x6n/z5wc7FCnINjDK5zcF9VdBmgfYK
iFwke9Z2ooOmQ34TPearXl2do9P6e9XNTA9h5pGdCSKy+tXbLQnhHZRkGKKx
otCTY3zFDP5xYfELBgudpV1KirjkEpf8P8YvF67MMAaavXzEqxYr0MDGO0GI
4E5Stccl7Ggksm/WINpgGtggzhQI3kyWmckaj6BrbJFVAMSIqDzECv0tu1T+
BfkVtFKPbcJy32HIQGV1AicDhYGZT5v4+6aeIdsBgMjAD1OnJ7xKEMHo3jPb
MMfLydVmVauJvP7xV3h6xNY4rTtdJxyg2VN3BO+9vQ/8DCjpUjYzlk0pXbHf
uOZSefTsbO77Q5yVqVLwZasC6JQ9v8b+HBb/4iWBbto4Bi6HZT+ED+tnOuB5
c5uv/Z5ZYsWGFnvMG3oZJoTcWYQQPFA13IR1oTrqcf0/2+RPMXr6bxLOoul7
LAFuCASgADWbRrC82bdea9QHXqt3JKpEfxpssViHsFYltFWrEYWtfWf69YKk
wQ9XBKgWeJY/+L7IvU5jnkkm8IVoTmhprVMqNOqGLyxuXcB6yJibP82ws0Ib
5K1ykd+85FJgBRMG72ZOg3Dk5Vp+H3k2z3GrdiVK8Eo5zjvMNgGMYYntjiPk
Lplq24dEzh5l2/+ND3Y2qfokhs8V0JKqRe6ep9XhspxUr377pNzafFSAMl0a
7xhyah6ROaomoB7++8JTWrLZn3huePZwJfq81iEiwzlawxHrgZ4EtNGYM9hH
rJPHdquiH6RwATSTFv5j0MmujHW2N57D2uQhmd15VKIVFB2yfNwulREWPmzG
yG6kznhVjD06UnHQ4vPBWZ12EMHlt3XbHFS/WETqBMxOhMhrAWhAyFH7hUb5
VG1yN9ufHayrt1TQxfOTiFJIH1jkTxaXR8/xbkyQ0infgfBIxpKmGHlPkrK1
rLWgBFPCte2TMH9hkOp6eWfbDjV6h4JRlHhXi7+bIpuYroUabUMUY39WHzBN
z/f8SPJLAXgmnA+dH4lesGTehy+LsbH3vKR2woBHclyVr+3ZZisWz4DPxX12
hpuJNh5gE0Bq9EpOoR1241YuN78+eOkQMyQT5iNNKHjQK8aBTdkUDTeWlv2J
PzkVbUNQav7a4v3nWEJ4865rHc2OK5/URcctWp70gfY6gJkC9qPzO3rMbsS8
4Z6JNWxU8MfEHH1Zwh6KJ1FGHo7kgA1+glXtE8xHCH90b0/PpSq80ewmxyNr
M1c0mltPwPizHHil5tE5XOQAUmb5edJVQeJKH+P/SalZl6hqAw0gDpOSAA1U
qMg0EexRX1SPbT6UPRUBYNa+hK/xkzlIPwKj8dfkiKS4AqqxnxiOLG8eDsrk
0lZuLS/8/rXC03LIIrGcg9rB3S86yXp/SoJHctp6qjDOE3uPNlg0atnci6ry
a1SLtcWLSHqZzCmyu3tpDSkUyDpQ+KhhtIfvo1k2jKO+e2l+Q7GqKlfOgGgc
eqkbobdSxjmDJvTEkdCjDQOfH6oKjWfX0rHpsGA8K6BumcCOQa7j34Xk+NM1
/j2NdYdLy+l6BdLyC1VdKVuEn0mDWdN6dxFSpQYuM7QiI+QYiikvrIdSMFZJ
xPip3E64ua7XC1ovLLKUd3mAjTTrKGOxEu4WQcQ1lCRSKpvktMa+soUBupmD
gRXn/rZlvXu5k0H1KP2oiXWpbX7GXk/m4ePf3D/9AoSp9PPO0jfkyNtVACK8
3kUuP+23E4v8JE0vxfbXV2tzxg+R+Od3FuyJPDwZP5ZsOZEbBBkH5gbviTxv
Y9t3khPxSIH8OsdeAUC/+ziBffgQn7GdycCQRwGYGWDL2gG3QgtJky394CGr
eOPILJ0cVxwsZj6kLYKWM8GB2Rs7ARin0qo6nBPRvOKN4Zxy9FVMuZt9wuNt
G5zUqHgnUE3JipYmqRba8Gx89YD+AdLBk+gxbvVU9NXlVfx7JnsHoLt2XRaE
C/NrUYb/sIcmxUvc8IKAb22WpsAGWAhNwBVhbR5eyaJzoJ3C/8laWqy6CTKl
cNXJRGsGVWp3TvRb7dhJrKgLBqZwDfewpU9XA+UfRgue1ntuPVQlx8+5bGfK
NiIdlLgyFAhG1vTA4G5231pjsbX+BU/PfEn/KwyIpU3x0zzO8vH+eDt3bkVD
gKO/gWiNEyG31+cImPWNKHMdmAFhyXJmQ+cZmGZ6hNdxaKXTRRUNAk7vA3vl
omecrZ8sNurMtPAOsQW3V9SApyzaTGuY0El6EKK2bfGzrP1I8zxXS9PJHaY1
RAoAeMnu4ElZ7PZkyGmAls/ntX59wFvcejJ4k/Dp8kJ58JdYXkgIQQoCQyjw
Zxm80YX55LD9kzmMyREVQD11nZFTituv3Pq+4nYNk2TkIaYmWl4xLGdPSrid
bybfLEUqoyccyoPS3hFhC5aFMhYbrDyMYigO6og1cCkOSbqzc5N1nMMqotF+
U/oenp0OKKVw3Zie5SZnYigpxdLGoiqcGAUB14RPQ58ZTYYOEIqIl90/gSee
kuzCC+C3hxQhcf5cYbBzTGV6T8vtCiAKeFMGr5y0M26mxIlqIU6t/4Pb/Wy5
1pI6Yfks32mn8cdm65yDtGIb21MSFcIDyXkUom/kAMp6qt4AobzCm8q0pOEd
0yTIE2eQEACIX8FpfWasg/PClQ3I1kG/HW0TAAbfThlQ4mMXiYZwOtwqROzN
HPiLYQkM7WtZQABReXjsxq35ugd5RcEqJS3GpBFZMsMSSkVaVefX+gztlGDA
v5uiYBBxXkyFD1VZbR5T1GdfEl34uis7/qd7VT6wNyJM2surNUpxbVYq79l1
0thH52dR5Ot3rQcRnt4TEYKEyXNxTSShjbGS5wN/Z8yLkKJj4GMNFKlxAFW7
P9p35fafiJzLgEjuGjKGhu41/aS5OLBqbjdqMZtZO4XI+03QeuO3/SsHA/S+
79Q4SDsI4zGDOfTSKfjabTI7ADJOr4xk6I76pYqRhlEiJOYGerVUqmHhn8tH
FT4gp0mlPnyyLVfdUsJBMS9G5MrNZdmKkGur8SpHrImUsLAUquelauZMZQ/m
UEkQrEmNIE/SFZD41jFJtw15DuL5537o+t21+atV1r3N3iGYsznIzKs7Keb1
YeyipY7DDSCPiGEQRc2O556rUto+fy8GDabetIUpu/epFSSoKGHL07KScwg5
sR4ALhpfGSaZGOCi+faCgZ5uGJbe4w2CvcqAdh2dOjtQFg8o6T9vfQxvldL6
pdTR3vSZJjzA00H6w/HwRS516fcSpcBoiCv8CREdgl/qzLv04fAeW6QsQUE8
pvoaaE/iILAvXsh4aeMGUPJR5o2H/Xxe9geKrM3I4tJiZC66VjPnb9niJynv
ISjtMcY8g7O9PELi/vsru2+/dIgmGeQsB+m67JyLoAmktfQA7LfCa1IuEWnA
23/9tPR9PK56OSNmlswPBzmNdSPdulkOaR+QNappFvwrz2ZZMV0BVL80ZZGp
SpvfCRuO1HBaxvVCmPxcnQOEsy+iWlJhgw2AHdqKKfE60GbKdyPGg+mWWwhw
twQkD+LtaXNcUpaqzKHLoAZzmBssuB/KTfGBZFdvDXpHm9Ad2PfSHye2QoQB
4Gqvb68VWPa3t0jPunzVA2EwsO+mazEvJBBM6cPTEKWpWi3MuRhUnZed7M1s
VNXgG++bpcUEdbaubLSh8ekjJGlpCR5If2xYCbeGIkAyVUEkPxVTRZtMJ/TV
Zz6OVJCACns8gOkH3wPf0nK3TJX0oH98IYiJn++bM5HfP615a0+jhFMqe/X7
S4tZrF5V96l32xweI+4XavuHaHuZp1YzVOkikBVV7K1N3tjCaW0wIAc91v0Y
Pw1NxEjfRMfE32vwYkV5BOkrM7WiUABAhKxfXPQJOQdC1BWH1xhZC59+mUw6
IyophailtvoKqZLV1sEAFObnE682lMRPCvTIxRwZ1yqKoM7huUmHdXrE4f/7
ctMfcwafGL0yUwUpUUAguvw3UpojxO/ilaPKX0raRHmJUFKvIb0SqPtYYjcJ
he1zwt9WVzUtQKSUJe0yUZ2PfDmOHpoipNfXeupcCnXO3XmrhSrWJrE3nn9Q
cHa8bX7yTUaUGMjV8E55RyeJjZ751FlDwtKgeHIGpIzQaeBLX1NXDRZ3+rje
+TgiSl1CggdRSorQV4Y+YuanshdPLcYYFfQhbzVjF3408+Cd4PmBSlY4UDkY
v9s/7hZDYwJ92taWk9SpUMUaP+f4V1FZoh4TvcJB3CQM9QBMkGwj11kraA2l
qjJ9QBJgJ707K6uQLWbIrDSyivZ86g4riOXjbbNK5b/WYQAbO4w27cZr2/6W
G9fRTzXFk9EuDnkJTZxLH+fpZ92NuLw9712d9flbJcKc9nl0VsUvsHMaHrjQ
W/d5NowOCjlI0099SQfLYiw5LsRt9I+joSv2HgVdC+4idm8ITgHkEMHPJD+F
o+FFlg1DUlOYfPrK2PGaik1aif1smY6rAwVCU6j3ZzWzwD+sazHqB3KlNleT
78Y8zdEq4NNHqPA4fYnxa1+4/T2yQ1Hotlv/11sAcumbzLrzgd9P82vqluZg
b1zlyIfbpJ2eBG6lpwdIo05CmToZElM40ZiJuawoQr6uy6Z03NtJEM6dEk8J
/2uEj3KjhjVG77Eddz/RpFZb74gBX1TNAgP6mhdwU5FHK+HTYUfnM6D4wfRX
b4YejAf5s2XepkhPMb33htG9GrfSyy1J5ZjUFa/R6eWHEZZVZnXNYpQNTUqP
d+AobAz2JpC5QjMuEm+cdphn/gfTEnhYLDZ130T8GPPj1Td68KIAl48tUHJj
Y9z0ddsrzj5p8TmLOiYN0H22Mdm4FtBtN6J/0zS/+eWWZM51MQrq39gdUvx3
Aqvx0DZgeQJENkAl47VAiHB1RawvRjNjjqxwauq3qTARn1xGF5h78reDuBOu
Ds+0Mg7kI7Etbl07UMzmYlKePvCzraPhBspchQyiaSd1YaVcosv4BxU1a2pI
EZL4BVa7NyvAkdS2+258CmjE4Ae9bjbfXvSft8I1rHlTOtwjW43yuSSazAAH
NtjMBjkc3l0HFJELtPBlxD+PMH+xDuen7l6/sgKGaKOVygprTRmJsthkyEAz
tLqRWmWZNqS4xtIaXYIvHV5H4sQaW1ny6aBjDGAc0DBm3w/d/BKxYCLktpyA
hd8ZROCES4KGNflpZXR1D1hQSL2z2bbN2ty4f/oDxj93Cuaj09SEmwm+46n6
niU7owtXNQykteuOeWwhWoF9+eE8mqk1/yc2u9VSwr/1e5qKyFTV7RQ1cJcK
nC6M9K9MA1lNYtSBkjeaO+sjb3M/Cldnpr+UZ+TAgWDSdT+/mHkOeeYBvqRs
r/24b+9QqbsFxK4nsSebm+Unqw/b/WBOkkPdZ9528bMfPgW735zPpNkRI79H
xXYNColN5EfZpqabI2zU4iZk5I6nzlvXCn8I8Z7r+87576GtdeIbOg2Vh8/8
jeNNV4vSrs/teEUR0Spmyh11oA0US6bDyqS9OxPlimoIfyoSISvT5mvycakj
3mInGtBfyo1heHvJHKingGCG3P9m+YItFf8bu31drlMFSw8/JNMLxg/NLoC6
qV5Dm77/ghmOskUXUl3fXni79MTCR9ohiK1c5u5mGOSd8vd9V5rAtH+NmjSq
ajzNQWr8Iw0P3lYc1gzjtSnk+pxu68Vh12PXzA1a5n9S6Qq/rK4H1DNeTg6J
5rFZ+s7LS2oeRlqvZZyp2q1Jm322rjW5kNija65sM7ikIDZE349ozbwItYmy
jsuNLEkdRV9hNMD1rYvYky64XRMX05v9TlimMcpS8F0z9svHnXunxnk/Nrk/
rbQisFOFLo/RNKEm10XrjLgcXo2exiieGjrxMO38gaLS/mF/1sjhaabG/LNI
FXSFfOgkW5spgDQEcKxoS5wjY4CtLQEO7qt1O9ETFqxVfP8TSM4JmZX1GSVu
7On7eyFn72Q1i+AsLczBzsVJe6j8vBPjP5BRsPkbmeUVMEmfMpunUCG+Fb3m
sIWNbUz4Qn1lFjPxCIP4BuBnSkV32VyxWWDmHd8roSCdOYFsPXREAd2Ip0MQ
CdnY6BoxIXAEjqCYbjY3tpTCxl3xgZ28Bprz1MVjvhlQrBiSn+3p+VfaRV0H
CNvT+JOjW/exB9EDMoLVKepJQK61zvEGHV3VtYNRXisLv/SczIbhPUQsPI9L
rL+k8DBVEOmFBcVOKxQ8pVTBjyI5pHqvycZMdhda2DWOOPTFwJdy2CPBqiFo
Sc3sG6lWc4jQXYRNrZdFCnXQUSRjNBwzTWMjuyS4nZJKROUVeFLB96MwGiqX
aG784vV8KffJ9n4mepZHveDxDV4z+5xIOi/j28QC8KpNiNPFRR21+TjoE4Dw
xbbwPNx1cp1CaJbhk/FVgtrMbHoPBvj4QT8bcRZ3D+ngHbsI4MhB5X7W9dGT
BXaEivk+uoMqySFfk+YaZfIQ3iXp4thPPT03PQuNkvJsRN4fgmrdcrshHW8f
22Lk9bCBXJCfSj0s7vT8ioPu/HWpqk6rECcIsX1+PwdeR2kgJDn4klCcYkb3
WZQOhrXuFiKR91y3Wdyq4DpuVjXLOiiAsA1jw9hrGM2LgZ4h7vV+9ZT7kQ+o
FapsafV8Lqn2zg/0bgo9yYAyoM1dq5S6fQs75xkcjox08g/5nGt+FacI/YVi
keRa+nd6zcNzbmm5KSub0w1MLyBbvLF80u156oMnzlBEl4o2X99479eFTDYd
G5/TKTP183VuwNSkOqbkC41HUFI7bM4n/hC0yg47a7oNnrmY+J48A76HXzFt
+FPioAxT9wDX7jro9Egarv1S457DLOPBSOzvfZ6YtrXwa2sYUreUKsutNS0E
Oo9MZwfo3hXCi6nqQG1ljPIdEiulA+dkH+bV1/ISOR4dzvulo/chGdB7CuiI
k9GzhPA4gfEFLmmugjdyRlK2LXmSPJFLGzHiCNZ5SBIG5Q7JlWOcnOZpBKQe
LS1QdF9EsnNFUNGx8DAWPETMX6IBQ9bhcdW5YNrYutOnodccqAWcPPBcjE07
2ofG58V0ACTwEfujh/CoKuNFFwUcS/loK8zglme1fr6SGOlC8aPmjtunomKy
KFEU3cFXqb16D2c8dITcfPTLjZVOoLTqr7OBUDJ8ZabAttUfUqmFlYUasykn
Ei1r6tyNEkg9g16mmKiv1rGTE1QTeOgO6B/FzIqfWxBwjjnPoStPWD2+pBjd
bvKw7CtnSzX2lmL7SJDq0SyyH1QZUjbafxDSx5tu1QC+Y/L2vA+BYGxKm5LB
674GcC5LgDMX1bMEjp2cY9cPiVUfA9X4CT/bOVwE+0HP7bx5/MlpQ8bkQBbp
wJpFcVXMARLQLBTnoKTGV8zZ9VBiKPCUR5LiejVJj06Tqr6PkU8jrMrhm1l8
+JEenUKTg3f2ENwuQGGhpq48v1VYTuLIHatv2Cwn31ASIzJHRsgMsJr9D2FU
xnYVoO/53xTWL9dHQhA9WjiYdTsNSP6vHlrs+pwOscyLpYmakA6ZqA8qW3//
/8EJeyKumMu+ikKkzztVB/+Lby45cKgKUIVnfeZUdErr1Cg+Opt9SaB9ZkL/
r5ZxUGJ+4M44TW6XRxNfx+zWsO1xiZnY/kQOhdn6aN5pVpQmvQd20ZNnO5aP
Z1pwwuZK9OGhqKDwp451qwYSPW5vtLiOnP+OwwETYaYAf/jrEK5+7d7FvhpH
D9cS3K02oro0U7fe0J42HaEZrzPz3p06a8lccjIiVifAl/YcOvrR35xS/uXF
caLSEnPZWeZuzcYG2exRhzj8cw7VD4RvEhoBQI096vlGcDDz39uOlRxTvykd
xpNftL85Id+CMax3QrasDYOTNJBrWLGQCrWtZ8qI9S0gAsA3Fn/F6V1b5HZH
u+BvfHYDLVXw9wu813Y/RvubZfWuqJMG0Frr3/cliPJI11VKP9r4RlEk7tyF
/Agl3qpK4VXhvs/Lq4O0ossp5B+XVHxn2Mk+0VeyKzSJL7PK3Qj9VplDv0wR
w1trky5FSPtATABB99lWO6AE3gm09Tn3gql3bpsYvPRfHR45IV6DZuFzc3Mn
JqvXgULfOdyIWQ03UYy4CPA8LYXrWYxHvC5wpoEpAnBidTp/kDDZ+DhBw3EM
vuEinallXhRAsn4U6WRA48D7hWbxGx0NfhoKRmt/1tDaFSFMAS9nXVvaQCTb
6mT5cufBMZikyqGPR40ZVE8DPhbJaxUCfSP8S97IhHdyXpmQeVS6IA3s0h8R
ZCPDGRljQqy2sN1R9KO/Hyqgq7HurfGMXbO9opoRtb3iU8F0cHFNHid2VoFJ
8jdM93Y4S3fWWJQcY8mnOGy7wE7Vsog3yPuZ4hOnQKQi/qS64Z8R8Xj7bogx
4uoB4K9PY8ZV4KtG0j+U0+VTBaSz2Cwem3ZKL79ibYzokoBJSECa2kHGxwae
b5spFaL56xYnEhQsnGNngMRrN9iYVAoxrsJ329Oso3y6xXwQd6aWbTzp5RZB
Ia7sbyEzovRk2mz0FqzMRKZ4JrfY7AkoyLj8y4uFPe9ue3rxV6BaJdR2NoAO
5GmegSyaZ4U87YXfmhV14wq9MXK6NBr3emqffKNTsZSRi1NAhlqFqRIklEfs
uTINH8MBVrAJijlzqq1MBWHxlgPAbijzX5O3t6OpkNdpYq/uVLUn3oKs/8Nq
ij9VAFbo2B1jskOjOHqih4Gf/Bim2k4F61p6TBF6iq5wLP2CVjTjg0FDHrSZ
iPSaDAdFZlj+Cwpp8RkTfnLMiEGhc5wccHZ6Nm6R0ISwuhaCzqAQHRtadbKm
7LLdMjwxyGKBLmWqDsApMLdyFMMYMnWNaPaRs3fZTYCI42t4IUYzHGMNRK0I
u1JrD6G6fZ4ZrhpBHU8w6G+VKJzVS30ycx6MKPGzM/JAjasBGWgmCmDSPP8v
fQqymgrLTsA/lVcKJW1Amw5jXHam/G26MzfH4uPAx3zJUwYMgTGs8vB+jJ4Y
7gpK8PyC87hPVVzEd4g41cC6icsxVnYBiHz66bsJv5EHzr2JrapBaSNlg1Eb
LEOGUHLCcMbPzN36X5+rooPr+nbYlPRVQCNikaiPaYiKjZwNDubrn5OJDxzQ
80U3G1D7HKt1afsMTYgHZ6uzQ5pRvdlyqa0Bu6bv+j8Sth6da8SXJPnmRP2k
e0wuhLVcx20xY+SFY+dDXgGCBHz/q3igf90h59kF0UDc/BOvvp5qfIE2L+Sw
waHQU+4cGz8zDeuINQ+iAIGbIDDmQu1jANJC4CSoJPSswWclzsCoJq+QaBDY
2SacVXpiix0yIYHS8wNQOMWAwJCQ/T8lKjmvyr5bQoj1n4dWICJGbIWM++ay
fu28C39y6jP+FzZLdztbtzhvp7Yx3bbVIJmEAeoUYm6uO5Mw+/nicKUD9Slh
aaMARDtams7BPV/Tyty+9xAvjfhKyhbqa3vBNtwE1auzTaROswMUuNltw/JE
xgvQ4RVzwqDH/0JGjGKF5rm0TRisX4pMC6038laTxEYCSWvMGwIW/egBEp1W
imL0Rfy/K5K/wWOPfUEPlkdjohd9Xd/bENvZIf3dhGqUNcMayoAXpWNbAUJu
ClyYOPNJ6y2rtIpwdQTo9McOTrx/gJvRHkjtVXbUetjRZwu8JOu+8TyfOKv7
MdBLbtmny1JbA4IKtcHKPuvrn5VHXE5ixjq0+Z076OU7dZAYWY1pn9hG8jP1
jSTywTylUGJp2SWxtRfDddS2XjOa9XVXLk/aNv4WJkALmR4ovYRFcq3xGbW2
yQbdt2A5LWuIvAdiJFolwRUXQfQ4E7bVJPXrKaGqeHUoD1mbj0cMD5SSbnJV
wmhsokKR6JsY8Ddmxuy6Zj3AqeE3Fqjp3KwtZAxO9zItoawdfSBcukS0GV1b
DU1Sq+Cur9fLt4y9ygYAgZP13504B2xkgnJ5jKEtFcTAFGG/vyun9KmnlWN8
f2J3o9f6pftDyiUiZy0OwDWFt5Y8stahS9N3Ma/rcxnZJN4EfO9Uoi4vJzM/
R7ONzcANqGqKOgyauW0dURrRtiOdGTHHsAbfMzlTo09QbYvCE78bOX7DpgQl
LCfYf83jz1vnkCjLlDTzoXybFikG72u4abgtxW2S7UrT6395fFXYSBEuEBeO
FjT3tEX7qasXLGYT+Nz9xeqmwmw3oI/Ydm1QzfD5ju3PepqH41pmnT1kwm3S
l77105vIIG0PBzuhsqUlsdwqtvTva1g/1n8l5CCXceVmiKcovecwe5XkoUjz
5oVccX0kgtEZ5h8gODUjruus7WiUPhW8GfD4BMUyo/k62Aznc80uwLyO7ofY
nbYlWSQJaJxx38GFp4HZCKua1Td5KEYjleqRPgT2+RwqoQ9hQcVwROJrYDXg
LBZcUunEriFNBCFbWLZlhYhPvQBF5Kbx8UnKJ1Qv+t9KsDJAeOfP/Sf+mqMp
kiJqA6f0L2q+rVIjs8zer3afDO5MadNf2zTxOAQJ74jPUrMfPv1qHiHE2eJj
h/KF1gAgUnPMlAFUXe+LyQUaRXtm6MtC9//S+Vg0LZdrldrtrpqn+R1zpA3n
rjzWuYg2MeySHzctHT0m9mMUBSUqrQwJUnLrUJSJ1YlLxzqwtW0V6uiPrPXG
2fQmzB8DEG5S3CQkpF82wYQ7xCAZ0WVwKVqJm1qR5sxoxkj8cVZm56MuuRMl
iQXLamKRBVsBUTPf4To848y9HbL+ZbEjgzikxCHgInTKGR+uVYXz+9bEBEq8
u7d1k9y8IhrT0Y+lf2ko4ASHaXpds5vXFjZB1q9GKPvTEgUpaVA115LgueWy
0nxTTR2Uf+/ebkLJzL8ldRIDNAUKZheArzNClrSdXQnSsOLLVy1b1PuLAR7r
eGqx0UgSn3PBJO5eZ5MOLyhBiVjCiTtEdxhKwwBTZywxqxhD7Om/p2u5W61J
bQQfq/0sq65mjSAulvpqlha2u4TmzEn5V18d//Y7oquaZDT+wqge2D2t1BC5
D91ELvvsJwWoxjMnBX9MhRBBvPFJCoGA148U9zC9LsUmx8aMvEetlGvS7NQj
3Qeab3algyuIWp4Un+ayAGQYgk0aTmVPeEgqvxxr2KS9d8299aAMtl8TMTJW
ToZIf8or8EX0xi1RqEKkSg+sBN7nxLrBjPf9IbYyxIDQjqNx2N//2Gy/oJk2
Wcd1Sf6oG0g88czpL6K3PpP8z9T+1gpOdb/xM7sEa63r/3OHDPyTKB2FFDng
8RxemmU12bfj8Ur0jz5Ph1kSCsHyI/gw4ac/jdpjtXg4P+AbwacVJdHr7n3v
PIxstR1Drg9fDF02vEfH98RUZViYxLZcwol4xfQNHDPSaLvmU/USS+BHtI+V
obGGTo50wTV526Bv7sjZ08uxQTdC6G96/pnzVxFgyPh4jmzsToYfKoX8/f1z
iMF8hXxaIuHO+aywE3CnesHuOrZfh7LKQUO72gk2ZABCCmEbN/DNBgJpzjqT
uEJt769f2j1ecEx+dqzmytB39R4ZyP1HsG+ca/8oJB83zo3h8TJGevVH5B74
OFexLSEBS+Yk8DSwpwUM2+3DdOIhqeldYlovx7Loqw5hSr9FMrY7mVyM4IBU
cNxxYVjaJsFhpJzw8HR1DMYIw2R36ygbSPRRN0/Q/N3uG5Sbz3eEqQW8R2q8
k0kszWDiFkrFhJzRSXLRgGX4CDN35LO7an6tR5KmYa8rYucUMtKYABGsAT0v
b5qbNGMPeGhfhvqcInI9+Ws6RXmSNopo5Ash2cRXnwmxw012ExIq3Yrlztbd
3Od4HJIgbzbLVWydkSE8p8lEVGqKF4p9LXGZ4au0ZavUJS1YuwuWql2F4tFa
AAoYKQVVzlGy2mgn8gEeL93vWHSgvGiUahqb6urp2ZjJhI+iw0rJPxghMUaS
7kC3cHhppSWv6eDOYEUv2B5e7Ope9ZJv40rs+ymy7niLT9/7P1tlUpTHneed
N5EJPsbO63ESQaXVc7QzrqxS+P6LOEMQU2eQDKmsyc5twKd0D9iUjQjU9e6E
+4+fTNm7a1sSmQAYLtRolvwwVilUpxEnJiM2+xo5qwNZyOuMTzEewZK3vWVV
VmtH9qU3OeuOFYkEwHk7+8lCzKyZJqCRx8yz1WvBThy6VqgbJ/F8fiy0Rly8
mzmGxb8TbdfcgYoshHqenLJHmOw2q2lIQH3kgi9s82OD6/Zvmp6XrhVoCZ2R
XKoB23WPZn+jFPjC8X/cj5s0qYZ2ijvZsZqM5NSJAISMdPAEL5F/c4p62TRG
fGeru78rgEKJfQShJUceSHuQoDq35dA0L52B0DyALDP3hxbVOppmYit4rdOc
vpyEw9Ji7ooP8gDlTFn9xzR5qj/DPA91YfVmv/zGEpRAIPVtiKV5oBvmfDSk
h42el1ntxMWy6xDIKiieADC5IPzKCnXLgRj9XHySBRqkVAk+IkWCgit0431Y
YO5IgwG82wZeoMCzhLSTZ3zxxohu4NId2CAxG2z3toRZJ29l7BM/0Be+yJjB
zc1rNe/1Pq/3gy1yzmodJwexKje5KKoxXecFQGWg8oq7ejTql1PM9CUpPHsE
bOM6p1TzSpeJSmrsuVThpffOt4pfFpVNfSG0KC+d0eKBjNqcIC1o226SQNg+
lxNIRy4nd3mxnrcKW/rdK9AeBySf5zSglrMLpB+W4iiO8hk/TWm0zgjGFbQP
J09YqKEm2uWY4s2rfmRFu104ChHiEBAV6P3h73Wdr9I/mGrC71l2THicc3oc
kmAq+488vhjpGKQYczzq+b1Zt+VGiF8nJ9vuMK39NI50Dgsy3t4BPUL6IDWJ
8eL3Noax32ZI6H0atnssHNH1SWj7+1lW+F7arqj1U7EXA2lvNKQ8VPzi1tPA
gXxv2w1i3NEicA5XVWi2IpPP4GQoS+IeGP2oJy70dLSQ+xVWGALOoPR4Dg8o
t+xZIJvjxh5R2xTJeE54OXvoQsisAxT/KceCDRIboeK1r0vSauJwf3zlZqbh
3g8RSo3TyNyV2RFbZLGvpm1dZUh5YVcZNoVrdeYfzyPzFEdDajPK/PIexuZ5
nngTFjODQaxtCN/Z2MCi5eCmo6zfWfXzMKI5EGH0ieXXFAuzIPjWQL1TIT76
16CtQjZYZXhkEVuHnFNLceB50BzrBSqR/iYXhdjAUlSm2+uMBSfKAOBoh4M+
u/FUBk0NbzQBCnwtIRgJMiRD+jFiAssvQcY3eCD/bVps+I3+SvGTCCwARApe
VtDjA6jVhGc1uUOQtT6+UZ+kGzrlni1ityQeYSPP7uQiHVCl92TCjiabg4AP
6+INzG0rS5LT21ARDClsbJWvIvY/kye58SvEm1WjCj4upSygPQCw+C2uiQk7
9aeC93rzFeaZbwX8lwQY/9Uh6le5a0vnkISlKI/ljjB1MpwKYOaoFQytCH2w
ey1bWhprA4kpm1B9WIeHn144/9//ccKYU5FHN5iYZ6BjcKL+9Pu3Yjmt1BcK
Xks2Nq1i8vdvz/h3NFdoqPSb/FEodZsk/uwseR6RWN8QRLj8hcTlEp4z/9q+
Jt5BwG531BOU9Fz1UnVOMS0xB4KxmQw65Hqr5PjupZut8j3RzJCLu4E+fpgv
jpOzVYU/IU568gDOkuV4Q6+ifxTgPDC4YmreKVColIJZDKQOM/KrPfnMbQgX
R1b3P2hwnIHSCQIICvbWnx5fE4A8N5lD+FKR1s8xHbYIF49T64F7Rnrpg0Jn
vnblw1LUx0qDIWTJC/ArEebaPe8z3rLUQV8+1ue70ZhombScPBoOI9ywQa0x
YLdjJO3vJN0fgO9NmNvvnywpk3kNLxB1JmoofHLD6/K9lED+IoVFXr1LuI97
uSdjJCQY05ozE8qt0210Xn+otE5iVVXUPi0IZWIk7iQLMBn1+HQ7X08dg52E
jVZRYPZtQKoL947YXzWedNjzeVXs0IjRP54tn624AhIPnFdrB7k5zbRr5Ji0
dLA2NmA2NVYSyRcQo0eMMnjH8HH7gJ7E0DtdFiEtzwwFSQYOgKu4jUUVxdBx
oqk/yI/b2MTsif2aSGVwUm+xDERkECnA6uAx/z+gpx8BQ0UeW89quKk+dkH3
rgSRQrFXGCuylhNbp23lNSWpiPfBnlsCbvj3UI06CWQ6r0ZrbDz5CjtSq97a
4i5QmsHnyV4Ia7tH8iZ8QHnckcxwPo1MIiLOtXhUXEP3rHTMrWuWOT+MPo0k
64KFe5Ztx0vrvcCZOqawU5XsFE2/4WaUBCao7fGeOGx0dpfct/y4yLy84n6m
/ZkpC587P2JdZfBlYnX69N+RMg33oP6PMdYLWU4Q2HkdXJhrlxF88WF05pj+
xTShaWrjb0+eC166RVvY7S6ifzLM3N8AzdGIYx1Q3FdW6kfbsOi71JoQOCBR
MapQ8zd8LarjVu2wKKLFlHhp6q4HReiP+GeyDmU7TAbU8/g3MrNXQfrI9hj9
WMCYk4lG2tnGuuT5fuzOMBURZS1v9lW0xhKtG8sACc3CgQ5rSz/GnpbmKICA
xyaFJwpDF02jJ4uBpBeQIses826KFLOEhnuyglIl7lT3S95iAZswOwtBDwaC
XyIoHCmfjTPnYiGrY1DXOoIfi9k1vrextYG2ftiQe/dRBArNPztbMKhuEFLQ
kTEGz1U21KNi3kC2e2Liv94KhOUiAjKP17YjwE9qcJ+WUTu5ukNpdHnzalj0
UO27TiGE+tK1Yib119dYYr+ye6mBg1/5vKYzqJo94C4AMAlLfFCkDkwCNycx
o6Uc6rmrKCZKhRdzspZKVPsdtZ+6F5HDvXjH1C+c2Vci/5JgyGWK0G1Q9CJg
iXhHaw0Pauvj/RA7eEgXaQDsnzh/4O/AKSf6tyg6djCt0eEBhoZP6xp/zt14
adWUsrRFJaNzMI3pmL+cRhHzQyBNlV6vZ1eSntBAgF+e52ZWYwlPmnbqFfoz
DcyIvfySfm7zuN72yywlC7lPy65FjyiMtEf2vWJt2Ls++wOkRniClMywg05z
YY1NvrX7EeUTijVywdDv6xT3Djh5xr/cnGwE2q6FJJ04+3/MDmAPEGurwMdR
8ZTesFdZaxwlEYCNgZNivELDfiQGz8VSpaHR7a3EF7e//zN1z15KJV7CUiq2
s9JijAC14XerKuhKiRFRFMomvaF+b46IdC8vcyOU3WgarCbzF7JWXGeu9rg3
QmfFoY63YQqOP84xNaVFMrCle1zNrNUBmxpSi3/lUKS4zOlU2uDlJhVTRQvo
cWgiv2WwE+JprwlLVc05WBC4SdKr1T5+3J/Zi/KNBpldmXPgDPgOQ/5/tUXP
VRKtT+vvHXGo2ob8at5VG1mUgjExPbK+30XnoDc6PKS8UavmrJ4kgsFt7WQl
c6iHFjTRjiUUNu2Tg4HCxmLY2nbT7Q1O2/auiEREUTuZSB7fjt2hTGS3u975
Fk5S1nmN3bYqFs8RiuFX4hf/Dh74xhwrK0ooIueUCdj/08x29H8BltzZlqS8
YltLY/zSQiFS84ir4lCaUua+dNmX6TpVIhQIiOEYSsL1D27Rt+Yiomonln2u
6d+gZkCb1qK1WT/FYfGTy/2cYMuyN9bOK2S4rT9Ps4CC4Hm0/VPTpiGccGIO
0IqcfKT4NuHJkYj2BFPnvulrrEEItcMb24KA1end7Nrqj3Ez8rLizPRlUDce
+Aa6AbVkVc1DU2So3IxducG/p7FyuXl5xOF8hdbA3g9WsK/1Wa7rikCUtR0K
KWeYZ27GpNKX8VIz2AiT7TGnhN3xH93zk7zC6/8dTKgIbTItJQFo/430qHCw
+QvdYNwE0dICbOzwGlBgfKMijiSGO9w5ufr0GGpIU30Ox/4bHgMW/fbYzPnb
7T/Zux4v+lD1lfGz2uXlUGnTe3crRZg8OzDlZHpfsZSdoviP/PqFH9YBCJdD
fttCEV4qLtOdCB+AcPZfZQ8HZfCZw7c0/WARyG2mTPkfD3nqhiYOYRXundIu
eIJrUpZd5jo1qrhmoGYn51AwdR/oUUJuc13g3EpMDTsDeBisI3L2eFTK53c4
SKKRBQec/EY6Hs7RaVq3pRaaASB0/zfNqQ2kych3OKpLyAgYzpDK2JQrwMoO
sn8sLmhsxee00gcG/152VkhFpaDLfRxaMfokImq0Sxs2SPYuhmZSZYSIJO7J
28KyzhgTsSqGpnDz/kCWHupp2cOQ9DxXTnOvv+IRKg/ehCuVlmdHxnh0zqPu
K6qCAYnrGx2FcYHWf864PYp5Yy6Z6zQox14kSY96BYI5pKr+Nb/wn/6nilP0
0khObRaGghvgQtNNmfrgIiV0/rIjauTnefBTmOLBNb4qb6p+ooHmzfh84xXH
aEgL/PCfIzC52L8EFBzzPZQmbStCMMjnqq+9dGK9AFstt12uuFuw1F5d/HA/
k4W2O4/DxwpbpZ4G3KGSfpYRy283EA/DJ1gyKmyrinIcFhxj7UwqVGosXnya
dSb13HzH6u8Bfw1CNtmx+ljUVhu2vNL+cWE66tI4RfDQbuGWCZOn1lkgm2B0
OL2Lt+EcXj3XPt4IBSdhlplNUL6wDujTS2tE79RObbO3E2DN1INVOtvRtsxl
u0xqdOUWTr/7FdvqyJzWKZPsjmpbsxvj9SADo0F494WHiNNG6AkHa5xOQQ9w
cmoSy1UiukJ7Up6LOXCme0PAi+5IPiGGG//+7698ZsO2HDSuMKMn1bzN7PBL
wfMBcGHVPUFa1F5ZhvWM7OurALDxfSmbKqg6r2Y6C9kZr8w49bmmG/jmjdT6
OFIAw4QdH1RuTlrr12yfAGuRG/M9K3Wh5TiB83shhp5ATZN7XKL+fhBQ7ySO
6uAnXEfNYsgBONsDY7JtrF6ffmQJkwKaqVgmJC25Vx6ArpSG8oUfA/nTD5u0
hU/0Pb6C0XZM6kmNvj90inHI2s1WzoraEWkwcwIuxmOIPLUYebJKEhhj0Utp
c8aQx3x4anPhjGACyldAcz5iCKcjqp9fBEi7RR8b8FBgnC4GOaLC+KeGtR/c
sWcDme9dwcBYN1n+r0U0P/vcGZSrOI8QMPKV7LsXm9Wk9TKaTfkj389kSFdV
i9NJJJiamoRU3BF8baxHOWxwjsLh/Xt6SWMTzXnyCRgt2t9yFRLwWHRIRvwW
L0qKzZw9khaRkkyeAyD7V/TwiGZUDGTdEy01/vrfATuTVn0uFlSK5nE1fgMe
yEpdMRTizz8xlxhPI6WBjSco0Qi7QE8R6WMNbX7dnVbEfN8rCqSoK7F5Qyl3
QVN0LwbyUilZx14ysZFNjgcFusni4w/cG7WLchpiDV+7qUevglz3M8BeAwIb
B3vh9YEAbaX0HAOmpJlAnG3VslUN/PaP2BZfYhoPofdFc+TW2H3IHYU/YE8j
A3kD8YTDjQoGCr8IGc5GPkpUQjEISMvA5z3QylNKveHwT2pRtA1td+RytYkB
fZzzuUeyggMMDmWNpmfSW1RcbCs29hTUMwxdgkv7jAj7ybvPfVLG6cNqhi/p
JxIbdhS6YRfxWn7zk0RRs2vMTaoiiup+45uWNTy+7JfE/U5JTbWH7+Wj8c+D
MPLSerKmpK/ogpdenah3IYMoVvsXyu26mh498Og3yCREHDTlHqvvsNM1QP+C
OlXCqiCCCfZs0UG+QKX1st096j+sr/OlGxVGIdg2e62mPrUFBa5Dn5Dlm4F/
khmQrzSF2TDzcPhdN3FxCciM4B1jGyS3itcvwZX4ulV4CkezGNSi5fcdJn58
GAcPzsggt2JpbcbXHi2DuS40VVXBRPs1iAJ7c4h9soUFv6QumrxYUjlIfphx
R3p9SyQ1F1BRa2Vb589YrqdaG6uoOuEkCFURWlEKkwgUiUvwcoKn3KXLluyK
NUqKU/To5brLZfbNSapbPwQiCXRc8CGvK8twTOjb5/K3OKgUhk3d07eJBlzE
VgtR5oFuQYLDNuCCsDjzY6CU1EDV3amYBuKjTuLzz8FRmIBjpzBktmzT4P8g
TJQcAs+mU7SblvTEFCbJrphCnn+d11cKdSOjKMGZrPuO/G0/ZASiwlPpZUpa
aWhrxeYTPkuyt9BDaTf9J6DIsXorC1mJJa8l8HfvKc8RXD2b6gujE0SidDpm
u+O+o9WwWiYSbPiWxeOzfFZZH/U3zW5+hfhdb7aUbHmkI+TGE/17mdDeTtAH
Fx4nOLUFhVzhu1jvRI1aGA94Mu0omHwPH6Yap6FVhu3jWrOevb4L5oxpsKjy
SjSrmckOKSvO+S2UFllbxl7O8zBp0Awj0p7ksKzQ3rA1X4pRC0rr+92STD2l
iKPPLvcxOA5bIi3A/LHOAgKvSGMqKsiyAH4rhZWAgonr9PbnPCnr+A8EDB9D
ldt3hrDvIsHZtQ7eW1DKL2lW5tYjELFvUL07HTUJXle7cxECLdA35jCqqndJ
gWEdMrQtLn9onCIFC8rX6DwXJg4sL/3dNiQe4JVBVTN6jIXGnIODrgoHW0Vk
6JT6cz9d5l2PcVScDrXdWyfQ1Gl06JS7Byw/sJQLcaHf1cXx+1PyEMcTNZuU
N47WXkK4ehvxXg0P8FJAROGYe5XZNVqQnFEX5gwz4xAl12sxR2AsmzLZ4KWL
+WmMhW2zasyLj/PjPNctTYgADpgdEr3mwOtAvq+YkGPDxskZDIrRx5JlcbSx
YYQCtJqbfEi4DyUxLrVGxdvWyvfP+AsNS7fM/8A2NSqiJMqinr7uZN5aZ8TY
XfNgWhvrNiygaLGkn+AboyTCaTFMoExiwDcgVgOx3lDADYm0fyGTyuWmJrD9
unah7GAuK0ptq+jc+N5Cpx4KoqqeFj489qNaocqfdIn67nCLvNK9jTl9qB3L
ExtjHTd+wrzCazoDrf9lHdwqrH4Z48Lp4zs9Wzz+3VUBPod47BjohMIPzd3i
cHW93gX0Cokdb9krhKY/hKsYWzm9onT/JTjZEGuPd4EOa5gggyL/ZWydblfT
Y9tg8m5Bk46aBbKyDZ3b38MsKsNnBO1YaTVh1grFIE/N1eOzdKzR9POn2EZt
Mr9eCHE8sEvwBCZNL7Ey64M7mGxla/V1Uh6HYRFB7fAAFGh3Ol+iBz0r/cWW
3TWkFxLKaCNY7XMo6BjvDZ6a5vVOeJhGShLODcVziCAOM/R5M/NLTCCPIUbN
81BbsTNe5SQSsVr9Y4e0ThHs/VZfgAfA10Hv8ymoD/NaP5w44rQNIYYaCYHr
KQk1dwQC1U+bqdKF0EVZtsFfMn80ffuby1Gd50vedcWhJ0/723HDOWVES6M1
KKBOAyiu+NYKFmBI4nDgoXOQ1qzraZv72EgoXGeuYWYnKj2ChAtYFvdO5omW
M1rmiRz/xahc7yFvZ483k9/k5DWbO+pjr+B8Sv+Z/4+sE0rkv0RAv7NFmNZB
WTurc03VLVNf+jI3qW/xxHPekH2QR/8ztRPWOwQaOLPm1unN8ptmXUl5ca8m
Kue6POAK0U8OKhiHQ/fYnlijaq34I3sV9ONYYNvbaIGfCAhxUYTY8G0ZcKBz
V3DXVjLn+c8Gz7J2NzlH7QiwBpgSHFc7/H4aGZk5RVT9ryvsASv1bNf1v3Ju
usTx/yvWgBruWg9CppzL0cpm+OulyDBfgQR45mx5br0GOsErHcGJdGSG+lOd
Sv6akZB5hpF/5NlzT13Z0kTpEc843hr8dVBYkvOKWsj3mE4zCd4HbC+42pPo
WlDaZumDvCUpf+RahRv4A+3Oqh4TWJBOvCpbLZPe5431j+NKDnIjR2WNmvJ0
gWJMQ3qjWPxBpIYhULqVNcjrZkCwYIylSBuM4dYhmt+BypsWffkMX80W9PtH
FIEV2FLo9FZyQL5sGU1MNz7AIBFxLn8AslL0hKbl/WAOXXlRJ9D1vqB65ger
akY85H3bumNlOOd4hWh1+XTXII+XVzlRaQK1gJyy3oyQVZNw/r1An6ugAipQ
Q+vo6JYOAWQqXvzqxw60HJPn4jr6YcYLd3AmkZSZ4cKPmrxmfGRUKTy2C5oH
oj7KUZ2QSg4+kOL9xkn40t0RWQpWLO+77wAGWQmflp4QqkbYtIj9lCj4of2O
wRyTOWJ3+PcE+KbYBnz53LYFsF7/BFvGfGjw6PqsgK6NVNjwGMvVsAFiOVt9
Nqno32RqlsOrL1o5k6Vvh13JhqQmzPNdlA/zMFfD0EhRt/oYLZn8KwVOQFOx
e4wLjvQ0k2Cc04TlgAAlp+uk1/xWZvnR8PWSmAUB+7FbW2Xucsfo6ZhSVh6p
aaBJuOABmTaADBtl+qRflUt6c9xLlSuX3nGGLEKUwhym5SrPk1dPFXYXCsNj
j1/5N02aY1m2pViTYrafp057iRuNNK8JVJM2PJKcey2AhT4tpdf/SSMNz3xy
Il9f0ldtQaujDr8btk/B8t/mblpnF8sPpcfKdGDLVPKzbVhIaEqrLLcPYAIo
+NeBHmZ0B8373vrzLobOfCxooLJa8LZfCwu4+ptJJS+e/4TTrgoZXfk8PKFe
v+qIYQfjyeYRleZ5elmpBGzSDprc91YwkJ2uiqKPYXvg/U+i1pBNvZLQYnMa
w0mYgl7PtHutwc0cZBR1GIxFMnG2XjoZhRKoQfzxugp+L4kwR2MedSY9N1Tu
wf46i2Rs2qW1XI5eFBAt44kcz0a3gnpblkq99PzX9D6qf0MxiNrgfbyrQTkI
iYGPmk9dulIrtUZt54Wuhi+8Xnnuj5kAGSWATkUvlckJCzE06zhGrZHrrM3V
uDJ2c5OOnc914JwW5wQftXa2znus63LWrbm7u300PL7j1qQymlZMGoCZ+L+N
5/KCkfdPe/rqHIXzqrftPZ26qlWNM48CXyNKzsrijU3br95XyjDucLzDvYoI
SzbVjcGXsvvd4fgkedItFjRNL0xju2UFFZcgYeaiDR8bwHNGuJdgEgcjFTh+
QpEGN9aPqvnWOTF4lzO5T4+S+i9nNPZT8wqGVgT3NKVU30NE5W4wQoXOzjXm
+2M635yzO8zO98TdtJP4clSQwhOStFIzWjCKE5jOUfMsVLE32aWI4ouH2fLd
+8pGRdgaGiFZ0oGj8155K/thnDoukvE6T8hShd9g12PCiVcf1UC7f+6yUJGE
SqNaV2wSZBmgv/uK1qjCIdF7+ng2v5fWiBu1Vkv90kZggLqd8ZAyoPb9RNMX
CwSNzTq9LfblUjKRIF1TaHbXL4zrcpMqPICAg2Udq+eU0j2QuHF9EvgS8ibb
7qe3SBiTQiyVWSQ+K+DkPPIjRmd2+Ot0d8zMaZcnnb9IfdJRF1GRv3xvEi19
nKcjgr9uESyrcY2JQcxiBLdE74ul1C9Hu3PiZUOBRlHsv739YDS12oqIG7f+
RBp8ui8vgOgRRUOxAKQOrNdNm0h+xoZ9ansj0/xSp9hKPzoTcsv5ABfmU0L+
sn24yxw4prX17MxEFsqEZajCVB47AKOvrVBFKjlAYfepkTgHDcN2Tle1DvMg
5t9W9DQd1EMi9BPCi+k+rMmZtk2PNmhYsb1US1RaA9HZPBoOyZRosunXzxoI
a2pdekH7nvfUftBUgp6q5g15yGprKPyjCRjEInnPqet4KYGx91bMpQPRajg+
u84gVfzWtQeBc1JfG78o07CZh6JvgAoBBuwHkIKGkifCaU7mM5QXDEo2PRfQ
hSbl7TEi7zRYgretaMHWRIGvwZ5AujRSXdKzwAq42mMbLDQDIv1cMeTeNoOY
7UNJaGcMihvFgbwnfZ81Q97IjBUHDHPztZ5D5HIr/pRaQsgzl89i/3+mxwDH
vHKD3fvjM9X/+2TFjjd6WgI8J9m1CFNdEMb07iTyqAozIxZo9e/J0q3gAeyJ
RY1PWarf/hu1LKsEf8fLLYzfjmGSOLBnA8c/BdEql9hnjMUjgscffHqoDy+8
kSLnjOoFQOjAc4JYVlM7jnEEwFLXiBdY6NJSvjGuKG0N0LzCIAC+l7D8QFeh
y0ED1PQkzkgxBFG4XwqxC74R3QD9bBWlLCPZsrsXm81xY3OiEQCIigQp8rHh
e89kOnCGtm4ojBgtUIZb55LnmBT8GhJxzWD77HA0MIYiGton62/lgv7HEpAN
PTNR2Hw67bbWvS6oxQVyLrMowvUSL/5HSBGd2WF/eZcBqKH/Uh68GhsGlDU8
pwS0iwEnxzg+E2jKFQ7F+ZW816HsAp47III5AWa15IlHkfiaK8Bs6nYOeMTu
3FbG19+SuYfAusWrbUhKa1QLNu6wTEIiJiiZlrgm81g+O5BwtAgr2y3PcjVE
XX8PB8kYz0pbSN2aAYOq4w8YmSBMootswR77Ee1O3ZwyHbVAF6RC7aoFCivs
Qje2tHGhQW0Wv8dgd+0vhsS0xGn/6KBNWSrPT0NZ6iusX+kXTQN27gPf1Lf2
SSBN5nvVj+OrkrkpD9QIeSMgvgcg/GMoPcaVfrKOgWiHKZj6x2oqorAjI1X7
qrfFOZkXb5dJt1Y/23Jt/AzeDF57crgUSxgL1GKNV5meK4qZn+ImEdqqnJc3
4Iy4PYuwt9ighzeI7LwjHufeTgq6XU5xo9Qckx7D/QIdovMUXsyrwVuYLi9m
WylATQcBKXuew1eXm8gjmJaqMS/sA96GnwWNlm+sw8PUOOt7F3QlZzsxhhLe
KKB2QemHrBmO8JCDVZvmHFqU4maCc9cj9YnODr6YsWPIY5vMSrq5b+MDY94h
N3+RfdzGFa/CuuFAxWxQqBT9K9cyUxpaPji0vdw8bkCDQrteM+Z5c07Txgbt
IHiYJWxULy4rL4lhs5vZz1Rv8XJRpu/gy0Dl6hnXYE0rfDqteSw5eiPFRPIm
1xNAeTcSHbg11TqEQsbv+XUyxG9daW5CHMV7NDTTa+bAWtJxye2K6NsIFIQX
pigTBk1gBS6DjmVTuYQIOuCdRkG15n8ZTfn0eK7jD+/n21EUGi7D5GuYZdEP
qYRs0r3L7KOShTDugnuL13lg1+ZaU4SzsWs3jIGeP9jGuMJoZfOCIZOVLDvm
c/abAF9brENuo5D0/8vQ1m0yFwj8mu929/rALQGxnxs2fgUH2cHw/GSbG4wB
Cvyos7bOGsXZpHPmKKPD5KQZlJguIV7x5yB15+ipp1L5jRiVd1nNG97an9dD
O5kvoIR23sSGLeYCJAu0EzSTDdhmTqkqYGAiaWdi5UUpHUgLa+KwvukwnR33
ANxnK+bXesa4EtxeziDANQS/aGzhjkGPqjKqVLuin83rTrlRlcxNuIMDG5Ir
iUIqVPUReHpnhvsH3RBAsxSRN/DM4KoSs49wxuT2WAu7kDDNNzaIFSpXe5HG
Mt9jV4nj7Lkp8kGfgNfmeg5ZKIUstcu2PunI8Q4WttnhhpAjklJAgizdxOyy
1lrBiH/96aOCjc+xaRP2VQYRv/hGfIEOn0OYeS96afBSmaMm6CymVmvBnaQz
EOt9si5YRs+PS/xwGrM93jfSh5Rm43DElu+B2KXKSigRPNWqFR7C5SUYq6ip
ZNoIvv80UqKBIa+m4T3lLU4y08PqW7a3lrh/LrDKVSyEZ2MYyjXo2o88J4iO
It/eKHz+qWtODpuEL3ORw+Y2dJTzqSbzEnqCBgc4Qo1SpM3CeyS9pckTNzgJ
KIjx51/CY56Q5ntTxrT/gFJEdg+vsVFVGoiGAKjScpXvRtOyvIDvTJ8awgcO
S9SqaSPro67jUWWqVB5jLlvOD9bpYNIYR6qUq5L00k8+lK7MRMB1NNfC1oOa
fFKnmvsp0snXlx1DETIYv5dHrq/wOxmcwz41bRTaCFkjQClgTFtFM0ZK9Oa6
eT1KJBR0tWThJgqSLi9r67VLxpwUfb6B4zGgH+X8gkDmZ9J7WyrH0v/rH8zM
THxfDLlnMuTIkHAPfz0GEsFKS5sw29VmE/6wFrNLWX9Xz0cTMn1RHMj791PY
ZtMzFbwwsyGztnP5irOI+75xUqNnwSpFIdcfGk7fTp7GY5rJrrai1qfOyzky
7N6tuT75ENPAO0U1UK5IeE5QdU3GWNXJ7vD8oSqogP/f7ug5YXbku/rYAuKb
9Kch/ODi7nZrWGYHOsbCyCuqm9cn8ziC5HsvvmRaq8hVSkkoIg1c5/TvMpBB
fOmNjbf1jpJQSp24CCtN3O1iOgSbF4EScRyJE26jWIu9wDJ8ALHBNC0s/a4r
qbPh7ZsUfVtCb+2DbCP71iZycd20V0ijrqyzxJFsoypLBlX7+Oc/nv5+SJ7u
p6nX4UKFIYoNoWtZdGK2Zo22A2cbuDt0Gg+Uw1LjxthWefsVltl07rFnpUid
kCMKvwPbe1i8kZPyeaC2OGrrEMr2+bnycQYUZAM2TgehmW5TiZu+mZ3ohykT
SzTOguOC4CKFhuxm+KBU66517DzqQh4OZC4Mt0Wf1QVAfmaPHTyy0WpErsdP
6FsdDZcSXVDUzhk7ajtZPWOtrOm0ATtBqC0TmkF8b5cJ0WGCwtlE4l47ZB7d
okouIZ6j22bj/loI04wGzXCAxHwlDLfuhuhx70CaRIwlF6G9pSMJXGHuYZYl
bj6IE7sJgZTQODGoo2ingOsvCwF1utWVFOCKo+dVb0FipcUjCOMKVs9zAWNj
g2vs2NYbGlHJKzHWSE0B0Wd61Ud0gXSNdj877q4MAx5IfmHPdEk4XQK8/zuV
NEohi+1IXyCtarvcyBI8KkiqRx2Z2yse/C3IziNvZMKxiqjGRA25ad8InXjX
7VWV2Z68iiXJyOu/woyXINWPtUbimREH6ZuolIRslxSogf10fXpTPUIt33XE
4YZp0QAR++V6utXnN/7zlepvRwX33kyPtteI+eSgfH7HA3+ztBOP8UUyaBWu
gyfwsY2UGiLvAcP95g91MpHlqI2SI5tYbaMKs+jwCEms3PCWlaCbO8ok+jKt
WJx6D2/flEcfbYNMy6Xgb7bJq8f2xbOXP2Vw19qddZgFQqxqoHc1Pn11nMd4
AuBI1FwKV9JnnqAi2NPQID/mkxFCdG2tqpioLE/nKTIKNX9lyxLILdGmuTBV
iSKnETwqAKOJM5MB6Wta3RKS9qpFvcVihffOxaImpg0l8BP6UG92SEbWHYxD
e5y+JVeYNEhs5WVjbaki17zqSPhhWRp0jP+SFPfpSnHBpzFlcGPaln5vQJC8
qVm84tL1Rjujasml3mvJC4hANf0cX8kP0T/GPB569HmPQKyQQXuFi+LrPhFE
5TH05Dwm2a8R4g7YurJXHwHLe2xgTpIPyYfNZyq2TveFBqq0XhHEo8c8M9VD
MG3jd6HZAzpbK8IYzEgbXYOOPcHP64zYB/BNIgwxZ+yfbWU956n3wU4lzIs6
t6pBMoVO44zpJ2jrSz18itX0xpfNf0MIE3Z91UXOoFT3XeRFRYNTn2i/bs2E
TM2a15BDy72BSj6ii30RVqed8QAqwqd5utzNU8wFo2cMODD8vgC8CQApKJq2
sZwzvW0tNhlcwXKB9wPeJOAsQWTeCwGfFCQPmwlCkB9q9r7+FPx74GeWo1eE
qZ/XDmndIF6csNhFni95XKQDV0+s00AGNz4zXzuTgR483ywkFADGePAL/hXa
e3j42qavEtrVS0AWAJODRgJnFlSEojhAQVmL8lnms0o8PX2CxJaU1qQRSz4s
gPg+gcq/ndWZAhodp31iJh0TV25xOP9DtiO42OmMsrcUq0egEqxZHKLXFtU4
St5ZT3QFefrKMKhXja4CxLPKA5eguT5XctXWwk5bigyTM5rPO/x5XVfQTWEY
AAVOPKt80K8Q0bwvpMAu9fYzbT+W+D6B7yYIvazdbrLLecAFMRetnTQm5tXv
BfomafkKNSQyXF3gRh3tHht1r0Y52sgcIzGG55n9XaRQpOtt1SlzhYRuJU4r
MiMb7WVhowVX3GUX6NptMysvRdoa3nkkkf+pBT/A/ssq46AdZmnk2U4HXIU9
TEOjABZb0D2ubjqQGwIcIh3WRKzejxhq7jGRaSPMAYWZ/Tr+8oiehx8KV1Zc
XthjWDIBGRkNpNBhNXiNUAteVYJ/KfeNKjE27aX0WZhV3KcAfOBkAM1ssmDI
f213gZZOl34Lr1Drv2kevkMrFL5Q286K1UJAuuZ2xz7m/TkRZotEo6LzzNtz
82G9G6eAL5Q1kELjk2jipYnJwnIw5nmTrptRtfDxr41vvgd32EtWntp94V4G
Mm5ZUvEl/1SCtLeOgNpOLJARZtGTN/i3rjOz9+lfbZrS12c4eeR5dOTeX/uB
vnMH3+4Kvh22jMXvyiWp8yMIQDTK1iU4gkjpUI7cc6Ubx06O7ywmKo7Git0/
Wnr9ASulaNYBPNocYE6YQuvdwhM8avPjmtik4L/gUq7zjd0Wzo3RNViBvuPa
h708UTWW/SrD724A6ZZ4uVwihjdXj2c2eaBmbmnqpMUOEUQAh89zvAn70VQn
MwRy6Tl0cHxtlzIZUrhPBE4eRjtExGSS9qYxXCjCsguh//wWMTo1Xqt1qCPC
ezhf28Ag77hP2qTQGyi/y5dZTvYVYp+/s6Y8zxjQAzNdU1/N3em/NL44TDnD
3HXsvqxZYiuxRWTgveMm3yXciUMI0jePhG/mHqBz8rIcKsnQqV1bLo1eHUAB
qIltmRL5EOQ+dCaqDfvSRGSGTRhrAQ5zVNWWdfLQ28JZntQyquiexofbNxq4
raWELYXxvhz8rtRk+y/BW6f07nR5BDeCDu77F7lkvDOnGZuIJVxnkPT1CKNE
lpH7Pqf3UBgHE11e76E1foTXN9dD67JO73/f6Qb79ZMVUqLirVhE8uyunu+Q
Pw0DMWqKk0Ttr7stWXREBuOTUDdvoMunivsjxIs3qktlNYyx0/wBzw9LJ9co
dPmx+UilziFpMdQf7EsuDGzgBbGFSbLW3JqAvgPw5Px3zeJzfQSf4Wx9bDCH
hw1keqfeegpPBEjHJ+O9xheJNZrMWoY4ucqAeA1MglP8F8Y8EHosBC3Oq9e0
1YesVU+uDoW0pbIe8v5jANDGngrvjhM9tenWRrpaY8OQqLdZY+bP67QgpkcY
adL4RP4kWCAcMHakZb0nUEQvhC5FeMS2FiH5UIf8e8l4VW/vfNWCRmM9VfOA
MLkT8X5LuDQ91cJxv/eaNPtEKLl3Gc2BGKNUzfuJDTwITEFH+Z8fBm+6CqRM
0akQNmksxjD8AA8CHOp5f6ffsTyBZKbgnMl8JK2MnttWVbbBuNAB5W3Elrzw
/rCSe4McWEORdhWEwyQ5/g0BacKlDFAbqY78CyEqlJruuxTW1ksn0oEdYiiv
0oatg7IdGQNlZOXS0y6twbRujlqt9usij19E8ILd9ZFa9Xxaas0wTeqJFQ+h
ABumPaggWWOTQzYD8/Yh7TBdSF/sm0KoopCz5ot2A6d7VhSylCk5FYClps9s
ohc3rq0JAF6jXvf0jAMXOa4ei2lRwggZjT3+clxpTSe8BnvrTuWDWjowqLMp
sHb6L24vvoV6S4ag2TmezzLL02wG0Y3ZMeoUHfjmJ5NihWLfnXkWoObgopwr
FUle0ud768P14yppGm7f36jnfXn2pfKGGmp2Y2CGSjHJGlcdFAEgkf8YrFhj
Pk8rrZaZNw/zxyowZmTeK4EmomJCyWdh729/Vc+C9CcHd0lUh6uCLk7mPDmJ
Bm4FDP8VNwcvbCmJyWN1A8QRRr3t1o0bEO4ouH+OLqvP484rQyGd15MsQiXv
7O306/EVNHxi8aAwrRKDk4UGO2H06VKzI0RspNnzKDwV6wxBipZkeJbXhm2z
KWgkRoL/QOXRqOLEx2ZAhWQGiCM998VTzltEow9ZsL/mKHKKHoQvFWkBLrGu
t/71lBkvtefRYPkNhZpWPM2lPpYC8XbZwjqg/Zo4RpCG2dxipNLooA8BS6qi
BluB1P34a1qChe1ffUfL+9jyJiDLRKsYWoweoTR6Vmme4yNQcEY8pWR5c2u5
PAKQMRcujJOxEXt5kLRpBg0DNwmYqIw/i5bSCsHovYKAPXuW1uVFev61gvOu
nIhQ9e++ZOuoi3n1jEqFYBviBvxsxBTj6v/mlImdyXp8m0WCCqa1svuFMPqc
THTVeY4nkZIOBKmV7AxFPTSzTzbU/Z9/ILWbA2bPWRP+MSM1EzX8Qb9uapsd
trxrpetFDJr6eLjcqA8mkIuPe/vto6na4RV0f/C2plcto0HMlrIzeGKM+Q72
lyXR3VlU8vmyMpFFC+yq90jsmu64MKsVCR2vI+HBNtPxkBy7JNBZ7x+9HJIK
RYTeip7YFU2giuwFbFyd3/z7gHHmxcuIKPLBApyqVoRpHiVA3cR+NUKovXGJ
ndMXzgo4gqOxctiSRkGw/DWvdTB8b8ElVlq0EJ0cLK3x3VxjjhoRNSlgsiA+
UuZbNk+yvEiGECPO/3P3+96cfRVzMi98GOT0cjYYTmFim0h1OInHyiZ2M/yD
RGbGDILU/aK9lCLJlSpoBgmVuc9EzYLK7M2CiyCL7R+Kc4qIGwl/FnUfUjLW
+nvpbCBfyBnB7sDg4LYPQQ2zZ39xi/l3dtZH8O5NszYvzE9MqWIUxk8E5Nmv
n2IxwzrKXioFvfGrOeR1RzfbefTJw1EMDX8auWlkmkg23HrEdJT5pZQALzuA
yLRx9seS66XYTdHf03hsrFNn9a5kjbfR+bJtGr9tCtHYg7fcYB7coPWPlJkf
smium1zlFzw790bVzYZJ8TzkImimXZIqbVIAS78XeF3ti9cwRAJ9pumJ1SEC
k+9VuCKpamQlrUl2e6JKJc/Bqo/DvIuloUGc3flK0ptQI14sF6uHY3iOgaQr
CSjd/vpM3VMBKGJ6dv36kj7+37lCBq/7+3dGag94lk2piNAZSUN+S+o91sSu
ew4Y+ON5rUneqsxFnTNzMawIJPAQolsy+BmNCoV/Kl/eaN47gRIknzxGGzX0
akM8yXCrPMEyhLd6icdGUwwvdFhWjDXQ+iRfG3FbuS4uBQdAtum2rDyYn+8V
7XuPynBQu2PEDd5WcoRdtgIA80o7s3wYISQxuUp9JWrJAxbtmgtXwmD0Hu6j
M7rAHUgHgY8sCrvxzUmvJjto23+Ytcx5nFkC+GkVOAYzXmtUXzDn/WnmCwzo
6uSDNfRUoYp6Gg3IVF59BS36FE6A8KX7o6BX4yGYshXV9/GN1JGvqLEGOr2F
lX+Oavq7jl4gw782BqBVRQJGWPuPePPylCzHzj93RUh2CT+cY/2mGPo2xuGC
dnD1dHbAeGVLSTufSsw03K5hHwAGhmOhasjKMhH6r9wYNDpxA+d0wpAYBncY
EQFST6cYNBl+fBhk0J14ikxYF2k4YIYeMlmhvcS6fYFlmxqDSwcMIQMeK9HB
rgP2GVTMHDyIRfYn7mkOmRJ/30RsavDv4cbh54fBJEcE/ZIlCIysdmfaMxSD
XL7qfedphoWua9Vves+WRWPiBRrSGVWt2Gyxl/dojFJyTElS+kwINe5KABEY
hpB2K4Iawrsu+EjyiE85xMlkSinUBNBRFL6cZfRHQbhr5y5QZlqr4bP7b8yN
fb60Jd6YicamilYj+WJj4GNKKnVs/aHwxU65RlKkBAXfAWm0NdQForUXlAhh
Xv1RInOgbtlx/vmpuZcECwXhLoNnTzNEB3R6Mehn5si2RoZEA2Mrn3zy5W6M
+clF3SJ4AJk3vwWL+hOibLjQhDHZJ6w860G8YEMShCeOsC356EAJKyb3qoTE
jE4DF2EH3hDC4QYb4TMyhY2RBUquJKU7HpWjCrxUc9SJtIaO76Z22+UlLbMe
1nLopkAOD93A8nbMGe6BYxwpKdIrsRSIm1v53iKkXiYiViaR/KMnCU8wl8i3
+gwFltUpxJvdXlELnHs28kor0CPt5QxoDquQgrfHfGo5DD62atAiuSXLoiRk
Yff3Vk5tGQxNnXhHRq40+fE8MmmCegf75WBW/VlWvXiOyduP5cpCfQW3GZg9
gnUcvSG4tsIvYwV5SbixhG5jMFMEWucfLsTdb8ceP4J4zw7R5JmoWg771Ry9
EJBcmFKG7pr4vfBqYLLSOBDbBaTkd+dSRaa0AZX50E7SfCjAnmsFvyYmpZM7
+08sozpqGvqzszb4JuCGEVIVhXylkEhNFUyaDJRJskl4zCT5UcKc1b5RKRoR
9ErlmkvT7NzPlh0TakUzLgTFXRItWPXkTjmFV2f6qJnZ58WTOjWKT6snQF/m
6ncdfUAXvp3zJULp7gpNtE9MprzyeNLGnDlV/mS/hTfRL1i6VGXhE5gDjsoD
tZfiU2qtwmZR/HIYiM62a9rEFzpybDHmJ0BNKahBMpuTfNMIQ5u28KXseZfR
AMXXCiTxs3VNN54vFFdUGQ7aPmW2dpTHTUvSqE+L7R13OHFvgP8oX7xl0HHk
CxlL3NssDBwPrTcwz2cSlGfJdTx4Y8fUPGzZZc0DSK5fJpirMRdl9tAiprdp
n99+QhqG4fjsERQA5y3h5lIQ/GYsHi8lZqNGl2nPu9tJ+Hd5A0Jql7yAQAcd
G7rpu+tsDTd+nisMVRlYbipqUepyZj2FhvZ1Sw3g0+lNKJpudlIJissFGi+J
UVs+7Jir52QQid9k9Zrr4xycs4UWfVxPunDIfTFkOKCtNojL64xZapAJ2eKt
3L2g4C9tE032WRPC/6/IljNM2oebVWjf873MrbFLr7sDN+xYC/CxgeaLoOc9
I7vDkFxL66DnleWYgyhRhRJrEyY8IY3jrjU2r5Ea/Ls+QUJd1mrb5di6K+A5
ThdkuPjF3uFGpcIj1d/e+9hfFCam8Rb+qPg52PWfjyj0nLXbKQH9PVU8XTJg
InLkvwyE2xwqjVcKhmR9LRH+eQ2pfU7u9sPkuoTFM97rIt4agc2xWUJCQiuY
i7NWv0gqcQTQpj1vQ+7l197LGdRw7eaqVUveT2dwYn1vMiNvjN2CodZcGTJZ
+QmwDK0fU1QzwUVAkibnP5JIbjip27UUIkAvstInsTFbHen6Qq/9EBeJ0uxh
OnkzniRVa0XqILT/xMIMls/i88UsuAvR4ybRoSkNaq5mwZ1E/+Zn1e7kOA+Q
z1JquL0o3S2p0rVqgTTqg8WOAdaCauarcKR09E+meY/uClFfGPEscMYFF1Ss
avwqx++V+ymYF1KPbVjLbHzuoA6L51SpA15Hyzh+GtnTYHM9ucRB4sQpVVAb
w+Tk/pX7Pi6YLu19ZPeiJ97ITBPm1YydMQCZpYtanSf5e/l+RS1aWhIM55GV
tx4Bc/+XKCqZTJg16kV2xR2NAdGe68rHh1BTAZDE58OIIMqkt5of3bCmtbkS
Uh4Z/pbs9v8xx4vcS3TXCNjIdYC6wjaegqFobwITt6NEh5ztqdYa/6b2cZVw
2tGVuRU+dZdIKxWHDsykfkLCLRywQEBq0Ms5+Oh26IpMIApIW/ZSMeX6+rGo
pYQb3JWlYgeJlUTaOQeX2wJEIZcqQcWA+CKhLZaDGZUWzjdvqactJOXOZh39
jrbfxptFGnznFUzjEanX+KV/5yEiKFcNrYYMt/hrxpFJoX5ys7TTDZpGlneS
AMydnhRzy2pDB9BbUSLuLKt4xcnvKhhaAD3VAJmPhU4foXBI/AOtuYv2KEb4
buotiviwD1R3wylg7WHHGr60tWxA6opZJFGAVpEk5JZoiYEPJhECtpBjzdh8
pv4ieeR/ufGC3+IQm9AeyIwcnFNNi6aJ1Q3CUS6Xs1V5w5W1zSXEqGOd2HHl
i4mJZtBXiu/vUL7zZo4BvfTQnvzxR6vdoSJxlZgFbGzc5klFs0P2tdEEcVMb
nxhl5HX0W2X6dMkCUXX93IWdVmTWwzjHBoHeLcBC4Q820ttDbGnBJ1JfIjCy
JLG9kDGniTzFmVgzpDMizFffVD/7y6RE7GW13jmx8q3JTIGR0io2ynax/4G9
lJQxIRMnL+WhMuOXo9/dFxJSTD/k3XMeBVk8w3A6K74VfOpjOQRh8bEXPEW4
szlXFCA0oWNcUeQyGU29oVKbJ4p1dTbGKO/qu27M8ZpZcgUnk0fyvWUDxO8B
Dlasvreiulof6meTKZjerAfBLtTgBLGDtubXM5Q0iHPoScK1CjgPX05Pcpeg
xUke88E0mklStXlGzCafdNT3SnycnqvvKT2UYPfcAPC9I3byO1QFTua6Iysg
N3/xqVXKOUn+5uy2vqviPqzawCHDkkucbcwvTXef3zSauedY324L5I+0jLf0
wSXz3aMjUP9hbB4xcS9RPbZSAsJW9/KaCecMIcOUuUYYdWRhUeiokCp8e3F9
Q897hoEmb/y5qtepmJ8sk9gUW+6r0tdpi7q2EliX+1QLDPVlzMMTLcKHNGVD
J7ktuOLxzlwUP0YMFUnsiTUChY9LZdZLZZv5BwPnr/9uE8+q/2m/7be1gGKR
mM8wiez6khQgPQ7S4w+AHl9GBVMQ3eQHW5fpw0hnRISvu7tDhvWU9xQne4Sp
wfjD4WJvI++BT3c83HsmtvYdwtxSnJIjQXFYfd9YQcabAxaWyqAAfRge9Sif
F9kRsHsToL6MI1EFbthWbUXt69gnSICS8oNPh6tqPZYwRrxySKxLgU7GOhGE
AlleaXTAGT4rVdqQdwt4gy/ttIK2UTPhrhmDG6n4vEStF2+cyXiTLDZT2p9N
zZ3wP+T2DPgdy2Bjtqv5kyLny3wLTK21uByk+y58KPkqf1Wsp3ChYsSJr1O6
b/VyKHmfzVmrR1l/itX2H68tdQ64kFYXBDYomr0upKyjmuG7hKtiiy6xh48d
5kWSEZhvWMZqAwxs9lq5Q6HhJAgGReqOWW6nGRdHzp6XW1aT5Fv7NvB3cdFj
lHyqaQiTgTsUSB2azGIFZZzxfVG8XohZ1/YVt4Jp4a1QkEi/OIjVdnItb8YN
XtOITNZXF0M6PDlGRqmvgtCanIWmr3M3/BPQO5bB9Ct/kJwONp0hLSzltvfi
WBGUmncuk+8DCesQyNaRuHTtu8GEKTVKEwF/Kbm88rb9nYirVKXB/hfVwTMt
V/JG/78jYeQ5xfL7IPHjma5Sg8C5InkzGK+sEPeCGiI9XlVOjk1JpwsjafnA
GRg+1UWjpRCrc2kFpltiHV+LXgMRn2QJ5TnMYUf4O5/swnsxNwNGNHCl0AA2
B9wdx9DLSppUPlKVVWxMR8QUyaj8+ETkkxKQ0ZRb6Xu/4HYSCyPTKOkJ+7Rx
nsUOJZqM8Z8OQfH48TybrruIhNoXy0sq235cus+S8LRmZT+zHRWjmd3KpM2E
ieo+M7W+05XGOhrWXyyrD//P8QuUK0JzMwhpyDeyiny6mEkQFO6F43mWpkUs
aiLLtbn/4j0erWq3cRcpcA5eHnwrk7OmAzgXXPlwO1haaBN93LKG+TaLKRa4
qENeX7PIx2SLeCM8XQfDWPyZFLavM8mMfo8ROK/KYOpMVtoWraRNIHGvqRKy
BGda341T1j/jx/RJEP6QI/Xb+GadpMZO9ndb1afh9kA2rOUdKSE5HRH2AhRz
bGKvFRJsfpxnCrXw9LCX25L3gbpyxU2IwVSmImSTE+1TDF5nko7+fflBdmqz
kqNhQJc7DMu3KfgsBXKGZIbY+XE9BM052E9UtdTobQtI8V3gegnVnmuCFBaj
jOVEmv7daEWsqMxaQXcBh97Snii+f97vOIluXf+FegWJqnDhQ+XM9DO0ut/p
LlkCKRlxA3e57Bj1tZiXlT+9X+OkOwQQtPahV1WNTIkzcrHjbCzELzXKVTRD
4BT6SbtG7hww2oOgm4ZQRxBKL3fK1hUcuzpOJqlhijb5xa4ftqh2L6aVTmi8
mPhy1b3qGDT77Pfqu5XfN/KZCqj8QDtliG246YChGf/s6/vnFH2uevDG/2dq
1uQOTIq8KY7w+WvVDvLom3r5kybYinqdeCZnsiUjJ2bEjAQWkrI66emN0Z8H
FJXtTyQbzkYUxGWizo9tCFFfyRm4+C7oPDaiEUjM+AnKuXbVsyAbmyxLLtnx
q4KTWc7lWT8tSMuy8ro5zv1qQ1yLjbDD8RoTM1yu51Sh2JKLv0G44F9kLUa/
pIHqWNRjD20sxIsszCC28Jam81g4LcCFacD0BoZiSa8DbWnxScTef6PYghKb
j2A95lwClIlSI0A3kUOEcK5nID1EKUTlbhPztsYA5IAApNW+yrkB4p9itGsQ
xqd8iYjosn0u8hftD1S7mV4KQ2jpo3RoFSQMiyS/ONvXI4ftfVb1RU1so4sO
FpT3Mu9ViCg12wV9TjtaxlHp8mPUH1GumNJcHKX91lxd2rxkr3zjhaMMl8Uo
3TNFsqzvsEYg0GRzGV6/bpNVg7dXIzXzKoEgzRKTGBw42kmMeNl53bOj6gUm
9nJBUu/tDsVSdLED/2MS+F8xR2rVPU+wKQY/Tw8/1pX6Atj6lzOquTWfs4WJ
niki6fFNqx4+TjI+HGzuPGYfAOS0u5Y3YB/nJQb/vqxl4HVeFhY4X+9KSrds
OKYhFchjq3+GBu5CDDdPdkZG01/SQqk+wvBt/kq/k1MIS1WURa981SHqTG5Q
UU/NklqYgaTNCZFu6Ksty5HPitV60j7Se2WG4n0YTUnwePiqQoQO3snuuC22
Wq5iAn2iyr0dC7GkLki6GjnTDZH4cOB+6oUissoA/LfzqymRRieT0g6S2gbL
ZfR0VB9PdUvk1ZBB7Zke+NxTNHt5ghK1zX8FN1E2kx3GiABVOV4ujK9RcZVu
55gT6+5gIWu9mIY/0hxH/Vdow+wxn5n/WuvA3STOtuWakJmsbZU8+DxHQ86D
hjC5hmSeiIIQ0/nrXiGg3FUYPmitVuHizUzbGrpRNrCcnSlw7yoGgePR4oi/
NTWj8v6SzjJmE3Gpr9GHslMNFTAx2nju4FoY1MdQfNBCvQKjoylndfQK6bZe
rUBlLSWaDXpNa1OXRr9Tc/bsafM/vTWPEwuKXnVQJGnmT0iDfcRGSD+RB72S
twogrfRhGtZPeWp4G/IR8gpvrvZvAEp7FmkRfXlhtTd8Wp6Mb6ULr3BkcpwB
XoOl8+jb/504Y7s/ddSG+KvtSyuGvLTFDVjWZafNQP73TJTFEKz+Yzrc6Mfn
yNXRk5eMV/cEOhdo/keyTBryzUTHafiNvBkZs8POY3xkK5dSclaeIm7APoE8
DsaNk0nUrHWOW6AEABfL9fEnFTZsY0nf0CqZf9rLFR7ccOMFgPKDPslk2mHF
Mel/oJPRamjqRVacJnnkkjgF47+nu6c615co7OM65qzuQYoaoPkJPGpAqbsr
2VDLngRh5cf5JUkqwL5asiVdQXVMKmP9h/hdcRnabeKa/39GesdiyLdTMU35
ROc+9Ky3o0Pi8nfu/M5DZnSgZv8Goc9wG6xcEMHS3eHdHpDmNAdoh9HoIsTC
IoC0pkuIdytF+Jflcy3odnyhOQdFYDWHEpPYcHOo0TuYSFygk2Fl7mPYGfQc
Va0PW68DPNACgwTmx/R2z62RkaAGKhhwjYaerdC8OOTHximJLfwwKKiHwjri
sefO4ud4CNUCdM2SIPKUHLSLsVvyt0hQHTJSu/xmmk5Ev39NuDq5/rMAjTBY
M3RD8jG1Bqib047q0wlPIYUNcdSDDf7FA6RjKDAAh/0Y06WtB0p3xzIFskmn
CmL1rTD7HLVHfDRNeMEfmNO19OKnVOyYPPs0wSAkGvGoMfhKHaPiLqSMundu
f7AmGD7fdQsjsdkGZDEM6Uup5XfX23YQ3+ZU9ylEJUU2sBKUX+J8lLUQZCwO
c3RUWPoNijiq/ediXmJm75QoK8SNEj153DzMbBPJKKIxSNuZKyqbhZXMmWmB
Dt8OnVi3d7SQkPGyc61mbkpM+5OKYggXudDhwBnL7/U0eNfWgk720fKWowTE
CjJWbxg2Jw2ZsdFux2r7Sxvf47PZ71mO20mcafiF+5y0OE27UhCuFEs/z7AT
ru199Tdu8e49lhrP9uc8Qq3tE99YXbC83FO6mavV+Zp2mq/BFJ+wIFQdvLJc
Y+OYccJw+PSd77oXy68Igp6e1apUyix/SbIiUIUw8yj1LgPbNLikIMCTWL+2
k7b1hiX34VMZYfPSHIFUciweoQYaFvqah+o2vWG9nW3NhStY2h04R9xfe4l8
oULBugHVzfOdYPlydH5J9zYjNgWl109nqmYCLSx+tTnCKdLfaHTDMoH2SFDD
6TKsQwusgnAPSzlzgJORxZiRhZCqUEy8UvuMTRtVJ9ifG8YTvRMjBmB9wdxC
+TyvegSv3sCw+F7X6K/oknXPPMeF61okZvkAKLMgZf7Ovq7+75lTRqoHN+Ml
mcd4Vfp9jGtIiGg3egS/PGq6wdvc5bqE5UWfvFjMVRYxWd8rycvrXBi31mr7
hMMW+I8W7dftwHE63887AMWVFP0gkrbo/vZVhYhlq2qtuT+nvCSw1BGitiPz
4spnHUNAz7f7VaBHHg10U0MXKVcA4BP1GK8KkG6xt8EYJx1nE2gI1jiahcwY
y/LS1uDiylI5oGPzWenl4UkPVTcFIU3b5Iz9iW+hSS43ETN1ZGThyyw0UJ7O
MDlZ1JJ87d9vyfIkyM9O0mdS2xvbcFurS3U9jILWbMkxy1tfz21InJihuakw
iKYF4w7PxntrcCxEOCTXuO7YS7KUXYNQUCN60fftNrAg5hEukI02dHYEBlGv
3UAorjwHKiRllzoLPoLXV6PXU/ImgV8ZBGMSTymuJa6Qyq2ZfojdudVm4XEY
QaNsrBWG+zFzTrOvVlEgLuftN3r0y0jy8n4END8aIzFXYedvJMqMdbQCHp7f
xooHLfGb9L5xF85GuZJ9YtZE39/BMlJ5q49/lGEt2q5FqXqADG1HrtOlAO42
K0J5v3lrXCmaKV1tfF+mdsiPwjCYJ5OTnYZhUOV7k2SAqLYFz0RRK+5o/Rm5
+JmVkeXrDJ6b3GzNsTRIc9U8E+E4K1OWmwYqqrjqUojcmHjmCQPa7j1KWF42
emeFMJMvOU0mAt/YYvubVJz+0wmxoWbhaSwSDe8+ngCHVNaA9htueplIJmi1
aUOgfu3dKykr3OeQn5WFF9PhMkCGJwOH+j6it9AlYtRt6jSAbGh3BZM+sP8w
MiUOfCYcyQ+d7ThG1p6Bkxf8PMDXRwsbuG5b9bLMhr0e8OOvS54oKR1ZyUn9
2FtD6GNohdwdltUZB3ek7sR0nhnE6sq/gybzPt9nHU2/K2PJ02vyayvkuEp8
54fZChwoTuM/aFM5aj/27Zoq/USKDQJl2BwR9SvqzsMIBLFbiTv++AmNHLpu
oqJiUS7KQN2953gfjpV0604oJI0HotYHVJ9qw3VF0z//l+QQy2TMmTaMpaUB
faC6wWPx7/ysr2u72BhfouJAu8r3wZi4mVWUFWiPCCBRApeRHdd57C8c66Yh
CS4FZTSe1UYHPUC6CGs2kudWaJRErPiMphHqHuPI3vxNdMq4G/1E8dzAyty5
H9tjj4C9M85OafANKv/Jo9aq3drI7guOkUdJMaiWQon7K/bPVZv376uKQtx7
h8wBPvNLhbLH8KZEhp/Ig0UhR5pTKapkwjr3yOaoGHApAlPVICM6L5jt+rZW
rxfsXppI8xAaw1LEH+3P1YDgB3/cpIbv9khq/P4fPYFWxoXawV5ownyKpP/F
dN+xal/yaFv8qq8TZDR2bMurA1lcRw17JYxts2G9/If3jhoCFzsTft+bRHc1
D2CeY4Sx4A0TSDcZuIbYhKEbhj5wp6xrvBF+t/UizD5T3zwkswt/GDZE4iuL
K5qacW7VxkJF3eH37ZvBRZx8n9hzkDSpYKycbtU+FbdJoAM77C3YsRdgAS9s
3vgXXhdAMhdCEn5qRVI1qQA/tqoz4ZX4FzvFdKX1/bEloLHUqLBkjIml2QQu
IiCX7QhhSNoNlg4uT5xP0DCnNnfGYDoZsYtpVA0au7wYxJvRAGSV7QCV8f9v
GWRLlJNLnHd/d0AbBKEItFK4aCr+XLR35XsEnGbCh2A3eBMDPnQ3/1YBi2kc
uB7O7dzOzBdKNZOxlIpzOYy8jycL8BemwnSDI6ik0vxoJ21x58bOtV21Qyvf
6BCxXEvLVwj0secJhyXznJc3upTU/Ce6Q0HKpkD+pJKBPtm7vOyBmP9daIMs
hejDzkY28qYHiJtLVDKdPIrU2atO9U/FDbE2ZIDoGjhxMw0d7Mcs/eCe+Wvb
n91AxhvBjBMa6KkULoaw0fAeNqcNFPYP/W3o4REvg9X3UfnaWbtrT7TQ2Q/W
pZuNefA/bY4OvWxZVVmAtB8MPxuGM6zMfmPpHPRe0g3kDtobPJF8EbftfTbg
HN7TppkXxV3vL/6sMNp5pJz/L6cgh1HS75lBwP6oAeu6ZtDUe5MsGxexm2eZ
6oZIvY1Yq2ngPSkU6Nwu7dWxmj4BgNlBiGbQwQNq0swoGJCadWVo4c60tPl2
euIx67tTT3Cbrdeo5VZHbQ+l3/1G/WmsmVpNNKBbLxUSsb3SESjOrDyIZyN/
Gcptk6nTAzR6BE0jFA0Hg4FMIXcim5sA2LIpdDO0xZyc6T3eAeYDU8wWZATE
tJeviZnxazIdi2oQnEQOrbN7dL2p2h1Ng4tugiX3J6/EjDdKIF97akDaVAYm
CupaRATw44A1KiFDvZDuKQQMNIrYdjcakdg2QrbR9qoW/bi2xF5HbpWh0r8J
a60i9xu/E6Relap8nbSJxO8HAU0SkIjXodmyG0kT5FL9KxVfMWmglHwQEnuK
zMaXXy5wetmGVy9qDv9ue3lb62+xL7sfIkhNwC6O2Uw3bGjXpW3+xL+5wRrS
fLQ5AXpS04V3n8XQ8ab28jWPQtDPlX1+1Df8295EfKyn249AN3TfKRJM8i7u
Ek2cBWdtwY0Bk+M7wLBuoh4V6Z1548T2A/js820WW/HWpK5OkQSFeXNS9Mxg
bnn616KsenYYvwbZglOhp8medEpuEs0Nkye71+qdNxqcuerwMxAGOUkPwOrl
XKwy6HbJifI3Pj5gkYjTgznpaTao/7OATHss3Twbj/nP49GxhP0ByrFIQ4vJ
60dA6JRtAyFroGUmP6XDsT4m88HE6nkWuuaHVgo2kDOOscSL+9EzdE8Lur4a
MMSzg0xHD5MYWfzPneIP4HCf22xP5nvlohrkLdvHtWdj6QmP/I352cQJXzCG
c3Clk7UHzdFTfh83hiuJl2uvE/qTbJYvN7hjurUuSDRxEyow0uRykO4PhB0n
6OlhQ4sxVMkyQhH8FIKhk1Wv/0NBjcj9D+crKbd4eLWXTYILAwOBa/mmOGfb
kG0fgLe0oFvWsPbB/fa3Psa2aEyS8i1vyZ+9VnkR7rf1HKsBUdrvmE3fZueE
MwHHdPbym04hwJfZSCrNBQ0o7HtBNvxDf3gnyn3h25BYaPbgbGg3mC8/SXV5
Nbzkb6jZS10jpVYVP+ouydS/xeJp1sumS7ldAn03NWYlDI0Y3//nS1nUv1uc
mlQRWedvUtuJJanFVEFP1aekZmUnjNA7xBhSfFGhwmCNsCl+yRlR6sagnuF9
kb/ylfo36Tj1/ON41+ZByFoxwTKDT7J2Y+q7fKa2iBSQDQAHpxtPpUij7dgH
YDFLrH3ualD45WipikBfBjtcb7QgcSTr7XeY+j4yX7XvyhNp/nToitysOpFF
2ZVerSJA+ULJNn/iZssGnytuz8VuiE9/6C5ejS/uZX4TThxyRGfwS9huapUs
cIA2mNMssGLn/eOMMcKjbYGRHGRTIAEmUGO3o+ODUvYaObI0VXcLhPwbsxob
TXpMnPYRbKfikclq6cTUdQtn453L3sZeMHckzM42x9ltx0po+6+pISK7XawF
0d4Fsq+iXs3UbXZUYpdMJz4gte1ttVC0FBXfnMwjU2I0DWOAT0PJVC+cmWwq
DCu3OUNObRI7+aKMpJ5JlTlk6ILgzb+RYD2YZHKQGaNn3IIyFFaHtVU+pbOI
337svo7NjmUH85ggIUckm/6Ont1A6Yr8r5d0KqepQuut5GsnZxqYvJ7D1D4M
nSz4nF0/mDADkPs61M7teJs4KoO/uGS0qx7fCFWtfjUeCY+S4jKRA9uFmvqP
Ln6C4/75RRXd2fzeYzfw2FUYtptGesuxZZupn48GhUKYGZn5KWEfw2ktIUAF
CXwUXhMCJP/X/LdTIwSz8RUoJZfK6WOYkWGUQNf/0GaAIzj1C5JT8QOlXw5N
miSUtpYnzMNRUC95hkt/QgzmVWQQ0UM7nGPq8ESAvk1eNoDItl6naIDVtzfh
rTI+ANAx6DhCsi2Y7WamJ++hExd4X1AYDvK5U7/YM9BUbvXk1p0npi9ZcI6I
4xNQahonsnSqbx4JQlup+osc4hPANm+VHJR+GhGqGcdhxjz19k2dt5WWcon7
D7WnIe+IGu4jJn3QK79536MGp7r6M3OKDy/OQwaf1ayNQbJua4bWpVOaWpRR
LNSxOzlx7IYTYFfhlyHp1XTGfhywSEb98ru/jZrW3a59pdP2Mj3HN1HCnYAH
D+yoiKhOuWMqCvi9inq4VLtW7W4abcQEiOejG2zD5RiQ0ylUARAhDyOOAjpK
X8i0iyycXXyBJx4J7v7W8Rd54lLJdHn/Zdt/AkPcHtRzu4AT4U0XQPmPjZBy
5sUwz21/vGr4M/2g4AZYX5SXxsmBZR95iXHjEJe1q1wCIFmgtH75E5fDJEi1
XpGOYPLmcNI2oQfQ7HoATYKacXSoDV5MNUwo9KO2aYPhBCnHjR9mMhKkT/IR
WcIeD1Un4dNqj5QKmN9LGC2KaaqqmjZKNfD05Z5gOH0i4fw+/SV3SgoAthLF
LmhP19fLK5uEkCxF1ylZa4MJ7O6UQ0itXUqZVg52fiqKjc83eCyWupTurAIJ
X8SWY/4H1Wv7BAdqVL8tZ9I6Dy39nys2kEyJ8RyWw8IeSpgtp+YYH0HcQegs
61+k+BdBs2pIVwlSCS+7zUXd59WvtOmW5gR/Qn5AxEAEncb5tFS3vO6DHqYV
BMLVziLpDawt0mbvAvvlXkjbtppGJgaGqTS1c5f5bEJKq7NgZQ+7ZcXl33g0
X0Nz14jqETRtgA9xFYhj3Bv+BAWei5PdIX+HIG+te0RHyYlhwpwtFu7CaRSy
l7MuxTyzlfdVFFHvWHnFkucn/DdRU0WOpd/2HPU1F4DM88SzmR46Pip55DJJ
sgwaCtG3E3u4gzzqeNaGHdn1fnVG/0mBsZsaNztkSoaVB+wLgJUVfYZJNHGT
W+8jOMeLA2G9a9pgiWerk+ZmUkarlPCeoDdE3cbKsQMtUh7FZHCjosJKkKcC
FTf1IUfqfJw277P6Pw1zAvknt9Gsfal0/+EpWk+HDRcKpOHdUvHUzqF4oRL7
3w7CFLZQjHtrzxvl4S/t5bmAfF05cdaXeQNOLaW2oRb/IGwONR+7WcDP0Tjy
JeGMxvlYatmEwvNPov4SFHRp73XEI10i0Gu9MFCQZNqvJn4ZVvAWvQIL5Fxi
1t/Pd/DMsbe5FbGGofsP3/eJ6nbm76iLeyk7PPkVSdxB+9cTJR2TZ9eDU9bF
CMUWnkxechJHF5ts8a3l3WFzCuv8NtTxJmwF7HVie4E066Q2dPo5ctJhnYYp
mKZRNpT5GvzSh4UXWOh0qs7AhbjcNaRkXqRzOpk9hYKAIJf5J8ImzIVLPZtA
Mp7K80hrrM8IpffBmQAD9cHlprUphgt8TAs+oahoLpUgNqxEoX98ehAyv6pN
wX5qVIiFd7PKIeBl7Sb/GF9eUYfces0TnzIPVdVVc7Uebe30LHoxVAxTC8Jh
Whcfw14jQnzeoFtpCZ+R1ZIqmF7dkxvNSP+CgDGIoAD7zgnBWizPklKXfP/z
edcVt9Hl65+QhSCWcIfSfjiocO/bL74VW0WTMnvnAhN6scbflw7DrIZsepoi
d3/ao7oNTKEOgviKuUMXECCMwwn7zweYSF6UcN/u8aZM+N2w+sYIU/V71T3E
iCqaJkcQAZMTssik1R2hqOEHuMtQpMmCqwsoSd1Mij4SB557YMXiCXvLktCd
98SUr4giwcfn9drvFbLUWbV1FWXM9kie6OfBMbA/zjFuweXA671vtNkGtCmW
MGoeoP41rPLsNSnspPceXAtrQlPWefsT6FoMDWz/s4BQ59naSLPL4RyZH+hq
fd7CBESQxrJuSH0+SB0AH+wMzb3lbhlBAf4iXh2NCFlOwak40ByIL4TUnDZU
o7MmQuqsB0HM8Pu/3A+fb3vxHEwjepcmZY3NgT3gc0rN2DXUNhZeABqcIGj0
JNsfRnpOrk8SZ/Y0coRGZ4RL5hsLU++0c3IQCgxL0h4EnkIkclUSbHJQ0pUL
2GAUZLdXk6h4Lkgl33Sbz4RsE3sl080fRpJWRqx/1eQomFj3jBWDEblUJYIk
mLxhyiwGfVUJj0BStagFHMgDtJPLJYlfopAqB1cFBpFJFdgqtvU9GMpNIP7b
smk99ULPxKw74gXJ6ss5YnvMRnQCGRCW6i5XrnT8kyAYa+e9HdSt9jzBypvu
qMVNODq0zzQrG+Y2DHgmuSSIGTdzZ7CLy8iT4pft4QehSgFO4UsyXuwCrwYB
ugIDLqtefz4IGGOEVWnaF5aT2wDsh4ep5QHWlQSRGTpJZoUTK3Go878IC05G
NX9g0mo85vFhFBj4KBi72m63WXYqYhsKJ8ag12Bu8SkzfSVeLl8udOepz9dl
mR9XRG2+P0hkiZju6B4SJbUV5wGiqPQixm0jVeuE4G8U7jqy0RA5y0pnrVE+
huiwQBIl4d3XFh6rVnLNixqM9D2/1UjgTQYQ96rE9Br0ZsfLRcbYxHr35Y7A
28winhXmaksS3UouB3vUJlRwu0mvBB05BvVGO2QDkwkvVzIBfGjx55MCvkgs
UeVkpg0+yXiRYaJZQ4qacl2W4wtggFuxK0A7aldc1dgfvieoveLo1njWQGtD
q/WbB8PxMEJ+gvHyOz2tVRai/AM36Uwb2ZTVIUg1KwmTs0You6+bkAmTwsyJ
Dc/PQmvEgbWLcQW0WVxVq3et8IkvvS9PPJ1pveGg6+uJn/TgUqmYw20cI937
rNQW0FZn/o7+fvN8vXnBknHouw45ekckX8zNQd/j/Qu1eNWGhbj5j2bOv54d
sioHsf67vga5bPfMiJgqTeSCHAf36/tWzqZEiai0lxZRRoTzHRf/IJ3xACb6
XX35SbepjkHVGxsz6hCXIQienCoNUuyy7o4bvRKjWDKq+9mH0zcS1fclKldL
ckWMueAqEABDddxf8o2dmJlSvimX9DtDdHMGP6nPeedzFIyc3d51zS2eQYu9
lbIHYZPAiILtNZgjS+Mwobr1GMm9i4NK8OVMcjJLNvBTiQHg6HTuCIrw8jTA
COYGl+dHvdMX1VzVfUVGIEiY+5r1yggI5iUrD0GdGF+R5QTeGPl7ZXeh9GxQ
ncFic4di4P+HoqVlYOcxOrhpYC91wvNeKJnDUe3KMINFbAlhjTGoWn5jaZAQ
ypt63NJq5vvHEomDLwwYSWKupw4xlbxkiH77UScxfGoFcKP8QG/WX5Enqxd9
dL+cv6h4e2/7VDc4AtfOmqIU+dd5qCL7ZHBhJI9XZ5c9kwOTdT+Ai2QFGZi6
ZoenJr56zjod2jAnF/sVK2wHCaG6NRFkS6woTIRru9/Ga4cOJK5Bc8ie8yJB
Pk5qyofnruzp3B/wsD3LJt/wLnoW7TBHclYWbJhTwq1xyU6Rvz9nf9Da8rYP
fLjpZIpEz79uWaGbl1JwwiXbKSeWGTFY3cRufkNzfZRIlw6XQaC9+vCj7o37
3FKGdR+FNDsI4+EMsixZr/LVfgRW5exYNwFqmOgTRB3QYIRnsqB9nZOj//yr
JqsG9x54o/wLqtr0XogxuzaR4XT9QeUhDh10gnH1QVIVM+K1P9bB8SuDTEOl
fgiKuSmHGtLvES9uz3FgPlZ0Gf8trvbL5jbmnJ5820hLexWvJoXnf/1Zulil
kD1eJQBUUwyChqMTS4GAJZmnbNqlD+/vrMl/Dn1UUrCBTS0lzV7yGLHb2Fhw
aXuei/ZUlqefFTKhVRj+7VEoYnE2nCJc4DPHEwtIfOsI71CvPf9EQfduda4c
CUgpIOeQWQbbwaneyCe7c8quLKrS+NqKUhA9Cnn/y4CDtjO5iw5SqtYMPIFp
wq1JlKXVV8kYwO1tWyrp3PfapcBBvXhraz6AT19UL12RGTyJ0ylMFEP6GQS8
I9B0/4DbzSRX80yZ6qzV+uAQOySdwY90ICHfpbOXPXC3ZkY+NTeqiuoATSLb
nKoQXPq/rRU1huR22SJggzZUu35TrBOePT9gzyLauo/ZhV/S+cGk+lPN09t+
GVEpjjztnEk0vKPAfweGN3tanCbB7Yt2s3WI38McCwfEICq66MjTV27s/43s
Dn0ODJJSEOmsAUhVHqD+9g/KH03CCaaI1/2guHfXgrNvsqsEBSQ5p+4lkr4c
1XxnjZZRqoIwXtahdWnXvPTSHBMiwpv0lZdM8uFPGj8n4PUrK80f3CSwwINW
Fo79XruJn9sClSQzH9ZzAz7TNwKihn5j3eM/hBjJXdP+PyA0hqJYFq3aKp+Q
t6MQbNWi3XI/+tSKZas6degTCHuZGhohLrVVP/BB3uBavY3c2v0Un3kSQs3K
6pU2NFF2bcbVDHzgRQqkjhPvRi38yzruGLUz696esgz/F8UEEEWKgZbEegAm
neR7nKkkssTU1phXs2FHNdWPDl0KN2FcgmvU8N3ooyMvokGhTb2s5sNu4fqQ
j0zBDiuhMKmWdr5a6aNDg+y5l73s+xXn5NWOBujHpRUhenw2HeS7DlWjntpT
HZyyrd7p9oEXxHijQZBzrGA8AToHHFY8aCKzwHaR0eOLfK0qmMIELkhqRD5U
FMGHXIBDyd/lYle96dFeYteNCESd5uHTWvDvAsLTh5xsSICA1hC6IS7M9IRA
v7INHACmpRcIOgggrXjusH2Hn8r+g58lmOSIs9x2CTZv5nIDLniVAv7sAfxl
9+FfzKirfRLryvy2sVw112vmHjjjXkM6tvzQBNlPB+42LxpeKCxQ9VQsTZzY
v6DA4Sq3nrT+vcL1gkcEER28bO/VrSkYwQAZiyB7pCIZLpBDQ1ER7DSgEkdR
IAc5SmCbByFKwVjUAIoPtv1m+Mspl4HH2tdfO2NDEYnihPU/UJYWrehnLS3/
Sf08PKo+msR7QfnNNHKpZE5Shooqlpt0tKHgoybxocWbOdlQvukn3EHz831y
HDPDVtUQURhQZg864HXyMergJtMUGhsNlFUC9LxJ3e0i/UydxO0LRuYMJFFD
dDAzWZax11KR3PfCs9z8KqtwT+wk74O6GAa2yKmiZs2PXlQWqAIJ1iricVWu
sgAbLY/ZKegpFc2L6OyjDXEQaIwXkVSVsBK4WJMxTPRlG+/1OyWRHpVxn0xO
Zk+wMGLCTu8isZdfP1MGZmmRMt11H38tLld7MLYX/ecxq3Y4TtkLEyFoKZD4
IAps79KSryjEsrGHIted6ssiVBycHUQ1agEG5IUjxrFx7xmi1lnUja2tTlTT
U8NWYJUcclftu+mSMIKgWXEa41QXWwGvG0pAxKPUnSZbS3wtPp8FfPqarpau
D1qKFmq2RaY3oXzRmOVEaYWoC5g/oRap0TTfOGswReMtR6hqrc4aKDLagdLF
Nq4V9OZJxSN3Q3Ttp45w93B4AQzRVMC/L8EFyNtJlwvQ/1eFgsMDL1cPVH1I
Os0/wfHc08hg8HNWLO7XSzVMCIXgtRUjhCJGPtknHK/h531FHgmedSfWIw0P
rxhAghOS3bpBasppfa6kWggHWmsS4fq2wwqfBgLZQk0DqWxpDeJ9GNlklV1r
HORGjEATLC+xUm6pxOuH2R215xGPhP5d7bxfmuehe+AFISE0awoYq/PE1aaU
tjCwXHayIFMbQllqrGOhIMfURpM++91XeHziIa0fgFByX3YnNRO+mu8oH1Np
XTSt0EpPxKGzJQWfbtOSg7g/miyQsrOk+oc4fGNRij92eOzY7yp53M4o3Hz9
dgsMa1vEkgTIyZ6xAH+LqrtJIqK7m7eje/cMIUhEsVvrS4U4vH1Qc8T7lrPW
0dqGEuatYfInOQZNW8vOUN0chBWIcjCbGarnhRd2emf0qDyGZaewOAYIoblx
+/9LksaF024rBDqQ2kok+daYIPndT2vULfanonc5D/U7FsV++uTZK83bVPRr
qTnJivWAPkuYuuPSPonxJrgPzDEJp/pSpALSi7GnXFdMk5v3SXYwLfCDjCX0
YT7qCJQGZwofubliI6MrgKUO1FdkEaYbo/LZO3FatlRZXpW1bPUJcwdZQx5b
mQgEgpQPYGC6rgCjGXL3JhmYNHuWm02oouIrEojsUwiLdz1j6vAoRjkGJNk6
6BnCcgKET4gNn/io63lCV7rhphsNNRIyj25EVQvV3hnG/tQgS+uJOdopMEoX
RI9jkoCKbBcKNqluWZCpI4tSWk5zG15eVRWkM/nLXaaWfvNtzaoUeGN4YD0F
otGSegQM2FVHoz+WP188A7w5TbASugFQH9I5kg8WS6VyAuX+waRaplZsqZ9h
KbQ+Rilg/NswGB6McWkubSL3wjDownzPcMrfUEDdi96ykovbchlQk1hWR/PC
MOgRHPe7hX9SOvx07XvUGEnpBCORxH5FxuFWkWag6Zni8M2m+15PE5FvyRcY
Wd1AGWFGiI+jfkgUX5nKYucZHRtvj50VVjfrubZHSypEGReLyMuSFadvwwVx
9hZs9LLpvYgISEo1+/AFcOjxKn/FNe1u6ZJS/bW8nJeE8wPOVaDGfsmfDYcu
fdwCAj4W00rCYEA40bf3A21eZIUjiESW77VDOYQjwjexzrl3xcHzEwcstrHX
5Dmz/PqwyLMjEZbTPXf6M3u9OvSjbE8iDhYgYJbzblcjcDPg/WN9Daj8rTRY
CvcemP18fP4IbKGM3+Bdtrmzb6lGL1Hlq10Yteak9sMcoX3ZY302aoNYw1/7
Hz74qqSwEOAXkJ125S84D08sehdiRbiQEZ5soO/44ViTVBbbrbxCp56MjcIa
g7yOXaUJOesII1SvbFO0NPm9pfW4+lyfVX+qeekMLbQCFHqXmIM50U1Sg7bu
+NZKA7K1f6iHgQayq9ySIHLXEUm5W4gufKj3d2fXt7R4VWuxORO4iYL1eltS
KAw5KiikJSxVyFi4uH9SK+kax9RGSgePofo/lI+1AnbJ/ruHTQ/l1UBVaEmC
MxVw0q1TtsFug0/RFvF3m9Z4fvaw/beMq8lOT0LtweDtNO3FLavorlrEO2AN
+0yKBEJowIjWcYKwTBqF/KeYhwoa2FdQZzUKVzIbLjXkAjz0IqR19gCvcxSy
tSLI4se8rraE0GBTbVXjLRQ1zMvDM8zsvmIDkGUq/7cwLkmcN0ZywO8PrWzy
zaDVuG2KZlJZfIdBwEByrm8ku7c+nRv/RA0yZQtsqIKApz/CGZa9vEgI97Kk
eiKo24xDovc7CZuJdarZAczrJc7wsxHc5PW180agiDlzyd+OCrluSQmPcGYv
WljA79eKKsDsnvwmPC84bdQDRODIKcgUq/1HbNNPed/2wVT1s48tfStTIppw
IP9nBhkyBfbCl+vgUX4FbYcJ2uI0fsHLtWuva1xJY5K7lUOfUXBlV1lutLsn
q3mOm294vWGoFmOHcvxVZsHxmySHsHHQHRzJXiDvCmxDXmDRhtypoeCjLKTb
oOHw0kAwVycMsjWq4+dePvkBtxMfrmjTrOvsjkN9NFRdVMSTpDwCQhpBGJX3
yvqW0MBfLNvRf4aVAXWtlL71MartwWmdU6VA7IQvh2H69Lj6HPeAfpqK/0gd
iu13jqPZpsoZYM2IYVqEgshD/rYEJIqPh82p5/eJXUlY4d/IazrGqDAGV+Y/
zogKZEZkFjETrQcrtS+LicIFTXhCGrAcMonka/Bv2d+kjvkkM98lPt5Gzi2J
IM2ewGhELJkde5L/+Nn8oxJocKs3wn/pomlXPPGSzcbslAft5x0HxPACeLRR
FweFIfeM2IE3TxBnmGiS06m+pAU999q/57udZbdZDl7ZN3IvWtDq15u9CuHk
WWlGXvV8OV3oi0eV+mj7uBWiv23dBMIW4bzBB7ZaMi4RNCmrWybJMEaMp0No
JVB0uwZ7LoJzMK0dnWYJIqDpboRQvFbJ0IvdfFzVPTsRCopTECJeB4xJ+y39
DEfpkW59LyuPsgy4OOsz/NHGcKxa82r56ahrkYS3dAdsQf2OO2F+V6vF2Udg
kywPMYaFC2WopQsoRfzRVUc/PHCFTSe5Ea/g40lhtd1I9MpQkBmfS+5lVzQs
9TRwB2d1fLPn3K+nW40w04q3x9u+xC3ZUjMi53BzO12gqi80mNM3D4K4N03I
gmZZN8udLaB2w5J1+M9rFnbIOPZ8uaXdMORslcs73Dlej16mqz3ZWQvgnqwd
iMB7yNXBmJMhckfsv7opZkGZj9VMAXCZMwlNNlJYgQW9RsUuiImyB6VLKeJ0
Ej67K9OlGXNyCj4bw9SNidvlgnSg6Ld94leZKlPC4CyDAglwou08DgJYELN6
OCQvBd4iXH+r6R/EZdEzCxQVKrpkrpEtVmYT4tx1LBtwcLvKoPWIKQiLNd+l
t4TBaeviibI2TjaPtpTMyF1VeQ9rMModejyaqaGxoZRJiF66BWdSFjOdR1Iu
LTP+AcjBWUfPc9yrrdEwVtRtXaHrWbRkrsZyO58wzU9Fr7tFa6iJ93z/myxt
7EcAEd+qMs1oIK3DHxfKCPYoZI4rJj8sgxp7bayrLx0omozNNwx7wXZ9wxL/
drv874kSYDGb+eaphtFJS0JhHVUQ/onk+xv68Y59Pf3W6vwQYPphNRscL+Y9
CKu6rA0KWHfHGwtlB5ND7C90HIvsQheJhZCCNjaZoMUs0reQ2PyepIYwDiws
Z5849Efzrz3csrzT4YVwIfBH+sAB/OfsteotH9orast/upRhr85eJiF9cwXB
HE6QVmLoOq5a7ucXIcPa33SECTZB7QEFR5svdCfXB6S0llEbuVUhZGoFf2Ol
tgSCdxDZyf7jVTzkAzVzjaVxxRsFdw6ss2A63IN976mnxiSrnNP6FofA0aFZ
qWYhw/I4ADS2xV7EctErigyzIrOQrKd/mUD0Uezz5HDDCsY27zPuhuQVejB9
q02xX+xnnaMH9q4soriBlmgpHoNrTSlvnPo/oHDFSBKNqsnFCCkl1p0FS0jN
kreHvl9LddlPCEWZreXMAED+/In0VJA6wZsDuqfID6c/q/AmfrFdNmu2fWRN
x0eSD/zyjuwJUg4+NqbYEyNATBKV3Z3OJFbXXM3pR9jESIV7NjoYbl6Vm1A2
hB59k8sLtjl1vB+E5PsGwRYkF1XhtaIt6ntgn8IfUE1tz2Nd3aLNvbkze6wj
yXA8qDMcE+yzqrDRdz2LwnZyOQItrFEikaegFEjz/sPHzPdEqoiNUr7bAmqQ
GdEEJEJJwmR1No3KCaZ3cw4Gfe6bZIhWCC31wj0Wxla6vC/nt2o+Qmp6KB+U
u/UIQcDExzls/uIaiEuf1wK8RabV9sWoOYfM2JtASvotPvHAQBY7rwOegaRj
4rz43NUthzbFResFU0PivfBHo8M5fhNdL4oPjFEbwyevOm6y6ItwX3x/VmcJ
ddaGP06uwXgMicq1p3tUSEQ4wtGyH43gNIYUftukkcGcMUuLc0ZJIV4tJSGN
0NKkfEdMjnysctzin/3bhi1JXdlPdQ7uwDKD+sgKMCdzSc4umWdM/k7Fx8t+
BU2gcxls9Flk3bAGm4PDv1et8Nm78ALkQRvNj9hX8bp/FBS8F0BAZWOjG+5v
wjFrNyM1zkT0lt8cyJXFrO3D1QamPT3l9Zr7vBm4WVMbwui45Ky8YwKJ8Zm3
bBf+r4uo4kbC5liTH9d7iddTlsJ/XByxBPW874KqutnolCDhlb9XhdG2GOEU
ffl6nhmXdqOfENdeDJaFbeuRYGfOknpnVS1UnhkDdwfpt2XL3pFf87q+52P2
aLMCgqpeghN696RZHImUJTPBCB3gzwnn0e7IpNMtSXG8CZ/Evm61ycKtPtYw
9LKKBVd4qkRhU4dyz+4o02L76wCy2F+BXjwoWqTNhqya+r+Ja6F0jGl18S1U
Rg661+AthAlVvir2u80x8w09cwwbdZYq6Kgf5AipQ956R2SXOQlmUc7Xt5xu
Y1srNzsORR7AC/M47Ipvgo2FUHTjoxYdVRozL+gs3poM9AJ4PwHvgRzhorCa
ihThXK3TRlSMYqn/cElnLMoqDdWBUTQO4F72r3P+3ihcpW90YgwnaH0ED/8l
LwR5OjFFVEyGLubIp1B2NAYhHFm3qjwlY7btgYxewsSGxqN7izK7gUV+9BHO
4E7+SoMyOfCN7j4yE4j0D+6Et4BZ662MKsBo9PskXEbd+OGpTxIRGZ5+FAbk
HadkdDdLgF2o4MlgbaSSoUbkRLFZvxRnrUpq3M+0GRAspHGPmKgL6/D0FFBj
p2taoO4OzaanPh+sG0KFQ7gLE0QaGsGtSOKbeazEgIldgUhb1Oe2CwJ8nJq3
+DVwcXcbqsxp/a8EMzDwKUW1AYhBqPnfLxs2hjqUnN66CAXkhZqsZ7aw8KOU
drQOl+hFEED0egmiPEbwTAtGIO5NIE1xCFaEqdDDzO+2DXb8Td3TQg/trTx2
CfBWC3IDJq8oSScnMc1k3Lk9D1WzwZMHePKdnN6KYXDt94OyIoGNjn84ZVWs
5yhG3BA7D6Wp/f0ge01r5Oj8X8Te4cVrTMOwJoyhKGgcXTdHo1X8EGItWTcr
BK1bYfi+8dCfskmuHtaWjIUAIaIMW2NzbgKFhnwZ7gSxHvRInRyi4tmusa7u
jF1Lyzn5WjGqpDu4L4ghOKqf4iPO5vBs5rpLu8wKXCK+GqkwFCTF5VEHBYit
Z/epTQFWl8cwrMn1B07etyas5ioZwRh/vnyMsglE5wtUZH1KB0p6M6sxQw+y
14Yn19AlNh1IZAYnMWd9BAquzZHMmZ1BLZi5NPpmj9Ws1dHVPO7+0rbE5iBi
JvPX+ALeRujgS3KQWHkPlqzHBC4bFFFHHvSkT72FyTYLqNP7JvZOzdYwlCwS
MBFBoqZercbdd9asxZwgoe87G8wqYiPErhCUnMJpSkJHTJJwX3JChhBZE+4k
9SYXXF3JUTZAboOBXFwidJcQX4GEOV09HSn0BGMjyYMEvIG8uLfa+5B+egZY
NYUs3Lbsn/Fy07cSwLAUo+A78j+x6qcH5VpYzOibilcUlP3GrR/gI/iAFpXt
gjrWb5NCJq2MFT/v8hQTSjIG9Ty7PELcQTTjSOav/vVxkOj8Qu7C9W9Xjmu7
3FsgJOlsqHx2tJaq0ZaYghjPaBNu0nKrPdMMpGIMR5R+FCuRPS6fzmK5C2mH
vxqhpE8brlPMzlZxupcqhMJRiGTwknC+4weFRe6HEVfmU+wJJYB8wkvjIrh/
QBjSq8Vtt6RYtSRF4UZ1+aGOOGKxAdlYxI2brn5pln/3mVsuYjMSLENVKjhI
d1DoNz5CbEv++++j4rF9ghdHqiC7IKcQqF+xElvDCrXGcfRyQrLYI7LS/CIY
jn3E2odv4g9zGEU0mJczAB+ECdSj1HpifmznAQwG42axT5JSLmjKkETGZ6Ak
j4okYwEmF9FCyyixTz+ajvqDnfAomeuAJxm3EpNW2XS+0rYA6e25+PRfqrDA
Ei1nL4OYQGTaTE3fYYtj4pR1s0pcPH/FOKPcJ1CsqaLIdqhn0BqtJBdguekm
JX1hyfGIY/0bxv58nAaEUFReYCypTQ44vF3DVmEkWK79TcKKN2eUJPyZ2Q6+
fZ9dJb5BKWbn8ZY1w7L6m4ZBpa8egEykBC6ziiXmPm6O03ue6px51YXFeb/+
bbpTgg0eNqJRkBzltHsXL7CYmxYTBMB83flmV6z8CmgoYQ4JMyM2PxbvFsoU
CfuiKrnD5ozrULKzgLY5ya7dxJ9yzCD0pzr0KxBMautn5dFLM9fNG91v+9X8
vA7vQ1Vj2Q8CAa6tsC0ZItlM17UsnEgM6FkypnyuOClXZ78erJRVz/K8CsP8
erPf2ztUNrVTg8Tk1iyggxm8r9bOyMQV98qpGvV3b5X6BqcGJqMTA/HX3ZsF
8VFXNlpC3flF8c/OEpx9yA+YFQqnUh5CQjjekw2jgfnc/lwxr0+ztqZczvlY
8W3K0sLavaz0uRi2MnWjO2Q9ystADGbWI/YNRrXLSJ7fshJ8LFF5UUaFr/PY
jMVdlCMrsinkhobJMAadI+SuZwvYG2/Y+AMxiV7swawPTh89oIH4rCQ201wY
3WT/uOi9khv4wZEpahu/WyL083fOUjnVfb0gaCx3Ds2TJ2D4f4vRASCZ42S5
RdVwETuihdqUcqQgLrJZWy2e7roJGjMwOiL7OTb+4QTFP2sRXAvp99BZdI2o
MgStXpWBgT2151QEJvwjig9J5j7zK83/8MHOeWHuO2SmZQro4HywEoA9UxNP
wLmQy89/hfUUHXEEyNKJFNKhbuK9+Q/NVcA49x+p7E+JxhF6thnpJ8Amw8o2
J9K/+RD3d0CuCUVpgKIR73QCxLEDZR2b7ANvmP7rGcpuVgpEfZygC5t5WAIy
GMZELiwjX3nW5Aul4K60lC2jUlXjSnO5kn7tG8Xw8Hr759EalEVT3lBH74hT
ATw9lffObHtgvzs3PFa+A2dS+X2S37b8TADzmq9nEzuv1XROLTkpB0/ol2Q1
fbhJnOrBequW49v2TU6mV3SRSL0cZvpbis6YO5ueqKL9XwRMmZ8zyRndWZsf
beZZbRVMCImevO0rcjq/1KATnEYK1Rni3zNAdzvOvC/Y8377csx/xrHq1aWP
d+2lPCa2lG3AnGr2dtuRfaJaNWWGquYeE4Ei2WBmruV8Y2L+wj8p9El2XXW4
dUNdPH/K80QMCMbRjJfvp/PT9Jgtu5weR/OWpsR4Se5dBojZbxwehb4JDAyM
UEljJN0W1oR/CGj2x0yxDBvNAP28I8fr4xSbvL8xGrumULNBlt4CiTPLao7x
8K60JsxcQFkdggNllS8oNY8akbfPvr5AwVlvKonNaJ9XAA+OBUqfTf/nV5Qz
C7iv4uStPMLsUfyEXnIpOtCzNEycaPLLPxecAhJR936Dw6PTdS/5H4sYs88C
N6saziWE4Tp02a3/6ECDlUPvSpSfMbbEZt3HewZVeUZMQWLwn4HZSrNWbBKi
Kz6VwDoK+J8R7DC2zMfOH8C/bPOazIZXkHVzM+ElPNRvvokuD8J+oDnRh9OF
Q5fljrb1gHbdebahDpafC6YfZIBkn9tATmU8Qnp90olkex/DD3lhfIzDs56B
RWtS10UC2qdIK8eMt8eMq97CFYein9sS7k/S+TS/fQkqDKl0TD9M7uja2y99
/llHU2s1F7uYVBI0I27wFF4OjnRwxko6aQW2HcAQ8IDKLlPwmJAc78EsWGzZ
nruT/yDhvA3GOVNJUohGNqVNnHDtwoJHxTocgtoUMVoT7zbyS718lY/a89+2
sS/anj9rnRBNIB87fMS9VIN1iceSV8KkJ5Rx7yKMPnBPREyduQNX1iEq/VxB
S3myoxW63iLM779gqEAROVuLn4TSiYI93XXU9YnrgDgpluki6NEOp2QPBoFC
2zZF8/ka13iAIrDA9eNpdGhs43Iiome/Vlq515tyG5EzkilO1nGMDVgMKaqX
E1yc+Yf+wL1vNIefhmlONP5K5FrnT17fjcSYdvovrYtIdHjOI3N5BWYtqqZe
XIXtU5CArzMqW7ydFwH7+bWyXmnQqBGXJ8XQoeLyxR+gkpzQT3CcuLMwiqQj
dFZzTWC5KW1uL1GPqFt8BM+xQ+wLZdv91qed5myjkY5FV8TNNSigtHzQtN7q
od1MqmwWQIIHkHRXKajoHyWe4xvNK83d4NwApN1I/ZDLP2zOk4wvFe9Vf5Oz
HD1G115Gm6bRY2WOdo17ixK9/J3Ou1znvl3E0xaCRVD53I67eAnHHNfcjURG
E32jwCfe6xtdU0Gw6wLmbeyuXsN5lom9pdDnnHaRDmH0RKthILsqYuFeI3ob
FxCbjXBgLIORQBZU0To9u5TIXO/RCBS1B+GUJQ2qFou6X5W9CIOUZr0yMiEO
cWKFQhAONtfyRKbsqnhT/JNq0SK68c8vIEv5J4ceX6Pedn14hmPwQQNpa51o
cN1hKmihKQGGVzM64RdY8dyI91jlm2Mv0Cb/knTYX724Cdlw9y5BAGZ35rrd
xo/qkfLydPAC1sejFHu7KWfHM+nj+myNUH2uhDKMkUvAfz6z1LjBTQq95sMx
q0lX3RaCdXW1UebOnjI51+yGh9YhFX5ObvmbPIpJ/ZTRIrp5ktYoXNRQXDh3
HX1z6Ybi+MBg2KPMLic3bX7AY8V0n7EnOMXxKdGzskGnevnUARqRS7tBq8Ly
xm6SnnBYp6BPueJ8dsGuB/4FhcXa6p/ATN7VUv3366MnHTjfOynOF0txbonD
PDpSAJptWeu0dffaYdsqhMYZTGu7Yz+ngtEIHREi2KR9VAY2FG6fsmS3/jLJ
HEKrGNH6echNFT9iFLchY3ttUyJueOpYYwBz9e3Rq0RX/91tDd4q1rd3NBRK
rRIGA8fjg1EX8bEj3TAFzBbvAhSoQAjMnY10M+YuTcOIdfm+IIiVOtmMJaLw
ClcjV6Fh2sx+eHcGU12AFLUSZ2BTcqMlArqg70G+d0ro38EOYMvxitMW03G2
nYVLSQyl/gLwJxM9FTRLnsalbFb2xHQuxfqupX+NmwKxnu4ypcsUhR55yxps
6w9Vf9CFP9XangiJfYufFYtRo3C0oLIBb9Ydc5oChQKKH9l65TwvzxeywCZC
S5O/1sZSFaXUu8NqqzwE941elJpcToXTTQp8ZHrhxfW0R8Lx+KsJW+12R2Ny
cvhZVAPAqV/OZCllo5G8k3d9VJff7U+SgIWBEQA2garevl5EruFgFL99pgTK
Jb/TVrCUvM+le78xsEKuwdJDriuQQJzVYcASPu/N5l0L48jjxFnuVJLw9UXT
n7T3r5S8Ru4O7uyoF9h/1hKAD+AZJE836fbsDeS0DOPdubCaoaSdF8hPRDOt
QQ9+Ff0BTBFF+/MJKNK/dLfUqGc+745ECx5edd48VVs8G0Nb3aQ8VC4+54UZ
gBX6ctOjVn29yHA4u/Ah5TyoAL7FSQX+4520gn4oqjOqH1uQTJH4rAfTNOgD
dbcpzZWXG6Nwl0BByyqxoNZridwGPG5j+1raad1Lxpi/EsLdVCjKBi9ZU8LL
o50cr+07LugRWT/IzExajc09+L6HCN2z81r3MyumWDc//pxNcGV1R32eZDma
dtvaYAt9tfCshEiB/EA0E9GB10VQffo00HUpQ03kOUlCStCLjTogZRX836nN
KtUO4BThTyNpPS1hGaEc927toN0SGTeAfrPrBKYihOMNICvOFt1dzJgVbYza
m5w2TGSilzw2ERewKYuKUkWXmTz9hMvae5Y87n4owOHSMBlAc7wjYYp7mY9l
EhbnRXhwv60aMwROC+jcN5b+DmHU1GtIXOddksk9YXBNu1/p0U2Iip2qnC+4
oqnW6/TwgNOSA0UpSOrdwvulh6fPiXh4x7dsoETOWfcaV8ZbDu+AtSm2zrPi
GMLvTrJdZifx2PcE0OR2zkoamEqSz5nCpSDrXO1TMJxeGsO/Mi5cC/JSLR1q
AQUZXYSlqhlph3K0RHfDsBxTQal1mFrwqW3bDxYQr73ySvSn8xkuIfFd3UYB
F6IF2DATXRYPdfZOkU/JF3zECfLYumaCb6WA5EWsVSTTuaaiaCPHRb5F2R4X
LmnHptZ/EbaOtSB+z2pGN6bIWtzAZEkNeGtOp6ZIxrrARQmNItGw2i73rZnN
PumlCBoMRWbmcv4aBjFFGRJ2YGGWt549SGp4gbvgM23zQyKQqidurw7OaWNe
rlSsN4BQVJFW+SsG6RKigbseIL1rymTfCgOUm2uvI9CmKmCozsgW7HmKWsV+
H5IQD9lgn74ebaPoApoPbJ2QD/AkVJJRTlW2GtWCBDyaU1CFYYE8f4PY6i29
8mXpQqVI/CY3xkhraDKthbFOToff852zPVcx6Wf7ZgZ33UWpC7VjPjgmFVSd
dKb79VTeTv2VTk1mk2WZLz1lwWuEf6ldJYMcET+EPIp+dfHl0At7MMdBesHs
t0B2b+QZvdmkFRqWLZuCOXbiKy2Gn6DpZKwW6NVKZ6Sm3ZqWKqpKmdnUs1uF
4S7rT0XKSuh5238aDuc80wGh1rdMVYMbHQe2ciAYEkTJ3HKZ8SjL5Fw+lC5k
+d+ORfop3U+dV12V9NW29P/TQaZnNsaLqCtVlvU7IbhBHxrWdhQGgz6y2CuF
iwCH50hCap0imjgpdisuBT1nlCCdvAeB4tbRQ4Qy4Vv2gnQZusdOBbVemKxE
5Zusy1EHYW94HOQq2r15g5vQUZp4FmXztCsH15+aAnJ+op96PJ3Yv/Z7NT8S
dUd3M7xMLPTBpT1cHAG2VPVOf72ghpYRu4z6E7/VUY425o6C62O9qMrGCg8y
fXOC/7T2KTYz1m+wlv+0Gsxg1uLJ0FIhZI+wEQgw9ZVgvKmMOK2lvSCoySzS
tVowTFGipVPgr8RuZQf4KpGY5vgiC+ZDAo3E62DS3XTXFFUpKeTyIlpxvJuH
9RJxc0JZXGVuV0q7Kp5j8rSgh9mczoOKPMgcwdHpgPtr/WPWtRKqNU3a0qJU
HE4ZakADQIhw1UlX81SBHZcqlVoqLHpyiwXRSNmiVCEzR5K7AgsgH7PQNe1b
lovPUdiU1XyBcG+RbiL+ZnjIBO05ZcRflDItO+4nltE51xncvNSVV1FGEwXk
xYyyoohFsJU048yzRtkdWaTcEthquapWstP6kJBiS0mBkjOMiunPBHXaR/p3
hcW6jGGUYAB9jnqAfYMeUU5aBndgudAdU5RUM8clJC8zUJYjiGyzEv/+dFe6
GF4cczxU1pEAWu2AzOnrMa9bovuBrMqhi7a96Y6tONpLnFkSJmhcQ1hMFFXS
XadnrHI9Ygjybv2U0DI+LKsyvBZCEJMSKpsZ/fwi3xzHoC20yHfXdvyi2NXp
U56HYmritz14fG6uSerALGnUyaz/ngTMvv/2cJe1AY8V72NDmmy0g9bAbVBd
XEBZSE97z4PSj9DCXk1Qb5QIaaU4WNV6M6G2z3LeJ99t5kim6E4i6tIEgv/U
YR856SMUn5e4lMDa1mI65oa9Uoy3uL2tFR0Gk6nmaKJ0uPdlBDGAQzvm+fiV
wcCTkW4efBM0rKde8wsNwS980Jv7OwrDmNzlN1bm6yUIe7BHBpX2HxG9wl1u
6WvjHBMd+lr2XLPcUf2Iig7ePREJsdS0kNwqOufU5IZRtiCxkBepwdE2w48W
hwgndu8HWoFpQvaa9CmASnhs30dU5xyXxBUA6eG73N6iTVGfk4d3NtT0i7bj
uMJW1SaxVK8TFCAg2sQCUgrel7MgHFyzAmghJ4nbaO2sRes8VDPWytjA4m/n
JV417Z10lvZIy4yRcwnELPkZXwXdSgdfslW/m+cfUzOt4bWuksRZp/Qp97Pz
Guy/q6Gp+0yEjOB3i6KPatR+bcr40EihUKDShGSOamsFvfK9EaVKkv2eWYak
DxsAJCtBjJZcwwcb5bKTzdxomp4IKg8DQ2tg8eDQUD4Jg40gJapexrOJvLhX
9NPGVrmlzvFZMQODRuVNu2bnvwyl1ybXmX+zbM1drkxNhtLatXNYWUJzJhQZ
SX9YR9AxITub4M8v+LeKuYxHLZ4MyRg4PjszeEt9noV10QKVr1pnEientcEN
evRE0woctq86xUzINKnr8MTkuBUSWAgCKb4OcK++WutIebgJJtzC8KW3oluk
p3eNAzGSbWG03Hc3zo1pNtDkH3eSMCDT4mQYBu02+mRwepRwkx+uA0COmHAD
eWsxbEZPgOet10u/xHLAHm1Tn6c3ii6BjdZ/lTPZSDFEaba5VYw4Z+pHc+Y9
i4lYEJ0g5oClPptqLMzgafjX17z/2rAQzOpJYkCkxM4YRCv+hH6miCpwvzGR
rMJFsglmjuZHP65zpgcfw9+hwQ1UB3zvNB9HsGXxMFX2FwkO4/zgIcaZOxJ0
Ogt07eNvAxk8R6fuNnYppGTyOevC/L8AuIZ3hbnoNizQYxKhcqe5cNgUJDIp
n9P8qszCM2Id2d66AM7qcFs5Bc3eawpvZRQwF/pUvRbAYFYHRtr7yAwlvMhm
tGOe0MKGUOTOId7+u89i1hrNQAAsU30ZV4wMY5iepaGbl0ntAmzD3iSHMhae
Y+Sd4YuBjSQzL0/ZTGyvv63hV+INf6s+H7wg61qMea40rWz/9PB6/2u4oqxo
1LlBx8nQHEdAAFsePJRG3LiqgPT6dyN08PIAMy9mCA62NK5qaTT2LEpqnGBH
X2CmpUed4Rt6Kg/6pivcgx9v9za5FNPh5hlYLEIIM9KqwpGwYps9m7ToPKji
BEmDSa2hV6Z2jIXLZtjseVOEAyz6rtDjGBS62q1gcQbKqzmtgBhzXiO+85iU
WDEM6xMxjhdkVeL19GbdA4qt8vowDHdOayg98BAlgeuZ45wts2KNvd6Iv8bB
rmPh4UBq2YMaguid000NnCRdHFTVhxkCYb13C8uhC9J0a3EF2rgKq0Nw+DXD
qjrvnguNLuPCiqaRccBfsAEfIF2zNHE2WnZLwkDafKqAo/uYgMu4xU1KSDiF
FNxQobk5xzAeskxI4TLx0MtkUialVUaWvYlrPNZOLKn+Kg06Q8eGS24s4k0g
qnzS8dn5+8kMc6uo40EuxCVQihAc6p9wetNMfNGxIHMpKCIoVvQdX7UTUnFi
k6IawUAffYepTM+U6vpG5+cVbIf64qWG5nbVCdiWLeGchzxhqt5nlQjVUIQc
S4ZL4FOSqPMBPJrbN/HzLpxCVup4dZv6ciGXGtA6kCtWtBz+hhzVEaqgnxRc
4f2RZVLFlByLagPtHHHwOgrTS1TGl/M7C7cSkoY9VbKENj3eAHhBv1dJThBd
TaF8WWVOL9hTB0Xz06mXfxDxV91dEhLAFw6/Mqj6rDtS77jgXU/Lk59o/LZh
UOXIajQX0tt/rCR3ar3+8ikF9rcBIMIMNa8L1Db1wt7V3UeDZVD00D5jnLah
kgryS4kSypEilRLjYFCol1Wfq1JpBX/wExHrWxI5nUxRNxmuc1dkOPhwT7Yu
eYjB34GaWIISDO6Bd3oYzJH7JFY/TYh0LlfR08heBUN0X2im2IxaexbvTqI5
u/4a+xnSKUgDYcUk2QaNgJRorWYbJ+OhZV5yRt3RyIhh2wQYKDbmt9JHypih
DOYqpImUugneRXR1aHgT8AlqjaxnnmnhaluLqFxkNSWJd2o3Yr4u1H1Vb/pS
NitF8jUKozKkShpUAv2JAiZRkRoc3It0Aj5YetK+gCrwOrOHp61A1mkkVQpA
QpQAHy1UKWQNUM0qLBiJ1E5qyYTAtWGo5HwuUV4jIxMAazl2gUXg1pfplAdZ
nMYPtrds038LjAYaQDFKvUknHbF3jN0mYogzZ6hL4m8qmsgv4lWaTrxD8lwv
UWWXfPjQCrLxl/jE2c7iangc355Hu+q/X8AKmT9ZslJ/ZCIxWwdQ+DJytbWU
4Jf+r6cBRMjbdHV7qpBjN9IiMyVgib/oLPpCdwHYU/4t+hbusekjhiTwr19v
lVCsnWnF1m5hVUHD/amlUJ2R8Q5VlmjfwyuUUCpf0O3BEQ+i5JWnGuezEevE
bpMnY0GjOfbuRzeH6UotLCPzWSR9kAA+1d+NYvjpvat7BK9nKV10O85h6iQN
ksr2WLQ8nwgv6ljMldLzfjOdKnDbOZYGR/IM1PcQAq9Go4MxOVEq9y9ihmAr
4G5wipvOETsCxXt//vJFb49246KqbTowLTmJYz7MeLrQVS/lfH672+N8ymE0
kRzgWqYMpGi7FHnMP6UZjeCE+ANM7M1FLpw5oPdmWoj2AlIVLGw+zgWiSJ3c
X8bwfQIntZTwXV8GBpm0mUyrword/R9lljevzu2pTQfSBs/Wo2Wc5P+ax+Sh
DKVOih1C2HM2MNivwGtAtQE0VU7VleyUvasmAcKrqkjMI+r2BJZM4utPfHO7
fqA1YI5wUVtjYIwb6wvL62jrakzl9af3zcaWfiDWnQmd5+ZI1liNZyBWEEIQ
GGppyUaEBOesV5T3t/ZeKVqNHBCfzlNbEUKWTdJgIRPBN/k3tEtmncmFQB7t
0tH3DFbD36cS513aLN8lQk3vQVIFINucOmTkccs96kf4tKUSMWTc396UHTWz
2bQiUQRpB2p6SkgEs9oz0XtwajlXmcjqpUzaFVHi+nPFJBmRf8tTJtrKOnxD
xcRqi2oT3O3InUCdIh69fz16Y4AnsU+Nn6xz2e4ss2Re0KBqvP0JMnRbGV9U
gnJ8128ObNcjhSgFWc1JEfZ++FROSj0KWekWu9YX0r++fbPeNqol5ZilFhBw
rHzEmq/mEWvV+Gsnpvd4vhnnqVd5pmdXA1jcD00O5ITAQOrRCg9GOdE+5NBY
AQ/v6gbwJ6AC2hxL6V3Ii5+TwBOxYRiE/eKrAirP8xQd86OGAZ3fCJLueZGz
9Nh6gBUSwVjaJI1VjthR6GKS2o+HV4TWxcialmOnoaW0+dQw2Ph+0eoiJuH6
kyDft9oi4cIKrcxBwO5pbgvQOpjbYCzn/LTjsxSwNhgU28UfQKhnGr3r0bF1
Sqp9Mka5oZf+UZvsAO9ucaxkgveLFWZP5ePz17XkY8/kftu61svWmsBxbJ7i
xkV4zYyN0zXwCGLpGKyxyLPx8FJ/veWKntRlcoof/va3H1jVuEXLVTmCCtgw
QZgERM/ckw2LG/Mm6nt1YPgjBGzFoyqmUuuv+l0tuDK2yGO2XGhVyja5y7Jt
qM9AAl+cUo01ikzvYwV+nEwAZyvmOoiciQZDCQpWwem7UlR1oANwxvTeXaXY
cs5dx8wTJlaaMNldSyQENKESd9hCuGBpBed82GA+x6VNdzJPTPevD927JyGz
iPUSbOtKOGxEk2qDd4pmK51gCpb9lpeIVh8K5SeaQYaEQNItaQK8lJ4xfIdF
dcJ0mTD2zwok8YeZwb0K+RcEqqkV2hEEqVO495fDi2SwRb/19HWZwEwjj2DA
j2Dc0+z/GOrDBmdxMbuqKY+pR1X62BQNEF36ajMlZ+mpxNYjoSeqgtHUSqFO
G09dwkfRsZbzj2IzQrTfYh5i4+zDsGBbEx+itXJ9XntSSJdCcm0L7mBRts7u
Kua8HlYy5vkxoW4xLsCIqlbpIF3b8kT0UAKcVAL0baxvxFPUOVxueKdcnOQO
pbc1xayWzmbMNXoPi39+5JKZFrLPzp9T5imkpTuNPh4LpaI9+bmKvnJ/nM7Y
E3NxjRfed/1lPqLnSEBpdggWp9hCiHrAEjEawn1nfJfuIsaAJr8Ez8pp3RiQ
xsBOmI5IWs1KR1ZX5VcOkFY3HPiTd+yhoTS/r7q7vXvB4C1Jx9wKxikuE6bg
Ne97IPwUWTPc6aU6fl4zRwa8ym/7b5+4KiWbU6Lm+P3AIMktGFFtPmPjvIJI
JfB+YY3dzKrcoa30qEMUoaTeGhOFYvxxljTWIUgfuUl8UpeQj6/bofVBK8Ga
M34E8cKhW1/OzwJ5fOKOgk8JvxsOcU/JggKmN5Amzmt+6SbND8kIdY6LaAs1
x1fZ+BYsjoSn87k81pRRdm3sSKfrkYdorjq/PH24z3pWD6qrsTj1tmusRo7c
61F26NiZD5LULzrHnaVfTzPTxk7YoJlYCgNzaqPvP17Ylqm1BNGWDcbMQIes
YDyWFOLvj1HfOq3cr6Ur2USdaTwpJrDcVIWmzncg0e957L+QPhp7ShRDT2+1
BPq/n6RHWx1EHtqfbOryDd8Bhm9IcslNmg3TfL2Eq88+7i3pox+O6sjXV3hW
zIFH52+D5KG70LnGiaGBOK6NPSPyA1dFmvMHp9+vXy/AahdQ4i0c9dmCWl6z
nmvic8Wh+0HeKwwWkL0jEFh1AuBkZ7Xfc1p/DxTO57W/L7rXAe2oCDwSO0Yw
u23ALsx0g0BlnH04dC7xUQlZteU1xcRfPu+dgOba0DljswGwhG2JvovKQq4j
c1+hXz8hmg3HTTshGMYsIbLKmf7Sj5gsSbWaXWPKR4AVTjzAvmCl4K/IfmUk
NPL+HOquoqhsR5uYvDhuIR6FJTT2PTRdoefBcFZWhEIxRf2G9j6uL6+ZDj+s
szBebWyerq2WQwPEpggDtCpJZpOpBJhuWYRTlJ6VpcJzF7l/hL9b6wVCrKL1
hA0egtz2VBp8zuqe7Rx2Wwq4dHTb2x9JQhjk03xBpJX1NJSsVbykyyGtFRQM
7LVFi6VsWVtIDNHsh69rNhVNbUnoqfVtxTKgVtDzOS5rnxTVMa2e5lSQU8Mc
ZSU1Ku4Jz+t6dxQo998O3bntOabAuLFRkae8XSzNH+XAdF67QCKzQmILPw4+
wXvoldgozf9jUujUL6p2beT004u87BEYnSu0etB24XMWISG/cJrs2XOfcSNm
frRAP7uzZJvVzFSvjMksREGIEc/o4i1VOACaFcZvM3UiMMF3jmZJnawVE7z5
w4Gp1lp5KXn7noyokAyQGUOhQ/R5q47x/RzYKpGhi5hrJ1alwDRInJNxjHG9
E+sc3TqS3zWxgwJrPlfbTdWg78sfMqx1RPacsZYAJn+SX8W1bEqqQKVCVY4F
dl1bwI8ZhmHzvTK+/N+a8L5OxGpBO1xAe7I0Hmhink+at2QH9exQpyiqm9On
hOjx7nPUfNkz/csCj5bctxh5tTq+XGgBhAcDB5YRqklOOeJFh3P17VikI1wO
tMfTwVQLP5uwr5jDPIwdMGUhmlAHSQ+y8bJtgQHn+4nBBGqWPdlkCL8ey0bS
Cn+wjFK5Xp6powudtHZAq05aovub0UapKpPRfq7oyeHLVy+R3UBQuOH+EOSZ
ZjVlu2hV5XEbjPHtMBlwY9jzTH5/RIiSuSpriNqyqQb74kTodXK28yKOTUxK
5x7Kk5npjs7IZraXfCkE81ArRTfHaYrl9L9wMLoSxPZG/O3OeEL5guv8+WjG
sebNKUsZthmcsg7jbVff7aMCmTK3EGZYU97D/X4FrfdGMtxkpi/AHpq3zIG0
o5UeJCyogUDYNpSKnAAbVBkfXAixoE4FJ5BCPBocPf1MEevHSq/qLH9D86mY
aooz/RHFprSwMxI60iN2m4IT8q4FIt5H1Eq9IvSWiAfd/jjwWsUb1D09sv5z
8MI/2xBwvsgVlVvhvUMIZz9GaqqOW7Z7qlbGeDVf5qzl2t5IFb35W3LguN6d
3Pf+npYXyJjmULJr0hyuLhmUoxMq9aiAI9DBxwJu+Vh3bxTk5gn7wg96Z3NH
gonn0MmgW5ueOfraku7zuFO1OxRJRFXwzbfyYVfMCy0qN32w/RMJh8R2rqrL
fTDWMBDI0FVN639sBtOe+0uNd+KmrUPvFzzVx6/D/foGVxQsYjqavvrhxBiG
bJTjOnfwFyeD/WNpkFuD/GxNMoQjaQYiJrdKmRw/rtVx5xeMUpRNaCXka706
V/22jZaNTxbAxccZaXx0kPW7yyOYraIPW2xNhQqNWaB1WuTtXUBk4dMLbSdf
rQXhIPUZkYXI5jZ1xCmRHGn9hzXu+8YMcqaUPsbxSstbYwjLfYjEROAJZ2ne
rj0ELn88DskIqkBGJ8sGjfN5THQJj37e6UlRuEK7mGh9Nv4/CYjR/AMv79Ss
kfPL6L4k5ZVVKZR25xLIEX8jQdvTxkUxk69CLHYYNX1gK58j33ZxEaqeUH/G
eOD8NvikXZB4xo2pV/+b6pj3Pa7+x6+Igv8BOs4vo8j+/BBpNmGVbTkH83Rv
ALe+yfv/sFcxIIZ+g/WZQJtQQd3RdhfoCIcwtbnK0JdLtXJE6i0B3ktsUY+c
qJMbXqVcfgpxvvdPim4zcpYXPS0g4WQ8EHfTNcIIcGiMQ+OYn8td0zKc1Hsd
YzfasMiTWzFcFGL5z4spaI7extUFZlV82RdQ+BNhi5NVnQ/xBBfHl2uuCl0e
K1E6BzTX9N0we82MZBT12yGI/m5gbHchTJZxmmI5GZZSvqHhynpHdz56tXUA
mztjGSiVbJzoOy3+coZ7nRTd5D4gv4KYwYNAG+OrSsxj8LWtVFdS4OBVlX4U
9e9NHaYdR3imnNQND4fa91myZZSyPzj4CW3nspiXumJ0hFjEyQiTZnUYC7g7
n+dr6si2kLr7ihM12CCX+dqSJavlu0HXqT73lydsRdg6maNoE8PqmnKqiBCT
7HoDbzfjEa18WXHWYQYiRumq1y/4fi5hMwebvVK+JVtZdVt+4IRlf/FMBPYs
v4h4f0PIDociLKz8Cw5UPeEExMcJMKnp6yuMfI7OhLpGYkuHNHHUZWTGIx/T
55UAM4YRvSB1zX0Hph7CU0cTeot2BJH75/rydah876KXCZZG2KFzmQATGkUP
lQ/2ugpI/+hthWVjh4CAV9gdEr0Rjkw0v4hZXVVQS26mu17iz4HahW6FzDGD
3MgeKOf9UamTiLwneqSIKhBLnPJTVSv7EF4Ga/KAs4uji3uQ/Mu1ST4Y7vyb
1szCtFY8JOZLTjkTC+ylM62jfAZO01V+mbDh06/i4FO3N2xqGidWObKxwcez
CKGfAg/5U7rwS17eycjbGZnqjK0LcofM4GdvXYTZxOiZGMfS2h47ItOVzUnB
K+2q8GhG8zubbQF3Blxbq+5HlESeZvZlZ19wS7qs16FAZQxr4uVJeFVKiEba
fSaKgWu8GFpQRdvRreu1IYFnxGqOvVDyGqCS6mUZDPUdLgQGKSfVfa0MQz3l
yWXrtLYDDtNvAbqDlT5FzBf0lRoXhQvAIDdtGPrA6PcHCzNWNWkJb8CK/X+N
/1c+advPk86gyz4rj8PekDJ0EtsB1mJZxWQlIpPHeQYZktO6wh1JU2ahkuV1
V7e74MCKNWbPMqR/fJIVd9hlb81LLpUUPvwjkseexiOP8iIjSUoR691OOttS
mLboRzQdKlj7qxc7VTWFK8a25rLpXX9c5VSUWnp8PFrksXwJNXhlvS5ULk/d
DOwbzJisNkpAe6GQs/IvAVH8yT9SKN2TQNq6cMKKYylxMnYWosOBAdxsafVl
35rxRVcKPt0M2BisVEQMDRBZoOvR4+bw/bc/iIf3ixI0MM3mcFXOP/SsPFi/
zRdUohg3dr5bMGvJqOGjaiRNsoLfIo/zzCEtxvfMpMUHJB0Al8BiiR9JpFeZ
x+l083TEbptv+DQtjNFyxjxjLZWJw87gyb7yirOgE+yMXmdz1EL5f5FDeopF
ho5+jNQs/milU4q8jmd8L1cTLQMgbqPYBw+fXUQlKIqtlAzEM5hZlaTvmjqc
dlpBjI2JvRxPmqFJW0RjzdGUlJDweq0BXRrF7Vm3PBCwfR03eJ3I5jLnix6D
gbbT4lkOGBvFKk5mEJ4W9gxYkRWTwKz6rJh5Ujzkj7ETwplQ669uSxAXnRjZ
L9JajIf30Crj0IWe+wcwvXZWO/pX0W/umQJ71cJ81jI+WubTL8NLwHBGY/sA
h1kUSY1KHmGIVvXbpw1j543oXivwF5LAnvUdgmzzJ4Buj/2TrUZaaKgKXxqd
O53YHnaCgbbGlzn/SyK63oS52nR1LPzLAyIs3WefiaP9x9TCrGTKgbGBxv9E
+PzgEkJGC5ZsAT08G8WiDXoS3ijravbPsQZo9xFcYGqXfgKFF5t/tZgqbWGo
bDDNIo4/RG+Cjvu4Xn6+H8EOK5MygGhYuEco6iK3IDunpZOMjMMpB0mle08L
A+G1/mkZSx3niWaUVS60n3Gn6S5ztU62P0aCK7MnXRPhHm2lRpFAegEcegiD
B9xoBogC6r/MH8DnI/PbpczXYFWVd1Okn1/3PXrcJfKPePxRKhXMcx/BJ1Rm
Nuss1QMsb7zel/9+1b5+ZzLgGjJTOdf4mppT1xB23C/k8ujrdeCJk5NgXEDk
V04NlBDp1mn4LHT6IiLF4M9Ic7hxledXWA5nFFhJ5uLV8UabSSN28Qy35+Y1
0o9F0dJvK9TzQKGpQiTZhXnz5b7bTBdRqnY++jSeSZ/fD4c/zxzu/4JC1Gq7
ydGOC4Fsgqr+X4iweTsiaJG7mhuKw53UT7wMx7MjVH3tbmAhRWsyiLJX36rO
EsLwVuV1mq1cmuYBaS+BwSH0UPPjTh25GoWg+SnpYV0hcIwV/bWJCuZSJ4QO
HGuNVQl5xPx2D8YEtwGdUPRRR31lhDCzcC/2Pr7lg8uFvuOx/pJz+AsaVb+d
0WTqMc5wWIIhSQWQ6RsJsMgnZJL5hMF0hGKoZ+mPgMnAgiHR7J+X9I6UbydG
lN8k6axctyDvYFRbvuE7eKOSYqgCHT+DZ5bkumE3Ycy6I1rScxznH6oKUz0V
c4F+nw3f+6Xj9z2n1WRNkIf5DwRKCJwUeg4haGODnHYW2n32qid3DTm7pzq3
aqIhjYiVmV63aSDswtgLTHjE4nRHm15cJRLTYZQ32jakxxbBmXDn2oMyMYAi
NDkCwIOMLn9JQMEFPWvDE9J47TQmBT/Hbby5Xy4eVCK3awdwuE90tS4A0vjy
XaSyYofmWwCvpv5V8+iBNV69umX0tNXoEyBx5AP/7ndmSaEx26ybP32hLuYo
5ht0SREOEcZL8oK7qhvs2sGS3eO9F34M5HZY722noc7sLLF4lZFozwT0rQM3
HSoHjsGzkeAscS9dZTRTrDWvvLkgJYa3VwcIJPKZMRhmHFK/YGDUwMukhgaP
FKdM87uQSuyM/uzUYMajSbIu6G4fFH7AGB9NkmCxgcRD/oqn1b8gIx7YrBzz
LrfwFI3Q5Yw6SHHlxT87gU6nyVgjgNdEcPzToC5KgsvDHjMEPcY+KKm1+wcG
BDsvse/tbyJkLDqqlejImx7sXsci9N980nBv/RFcLoKCevdIyfbzMLIRdWv1
46UD57emHc898deytWMP3Y8tT8Iww3hGi1YF5Ixf/bA8hbnyxGg4tz/VB24A
NxCJbzTZrkIFPx+l1E2WOtP1BZG4jxFfYsWOnBfHPDHNv95pXUY8DUmqj30a
rgi0oUPTD4foceUpnPCSD9kBAoB9jHpcvJIGTyYVeVzq7WYuS3BfRSZbHpgh
c7YRnRRetcQhcmPQDCA6KfLmRKh/1REzQbg2ef/FMYMcf4YuZPWHh2Q8IV2L
dWYukb9+TAOpQu3eg68aR2GLaVHgtuLTKjvGbmLolvhe/JkxTtbxwOZ+AsTc
l9ijJwDCuMwKTCjfMY9lF5pb97ULAZliKZE6wftneOn6Q+gNDEGv3+R0Mjqf
i8ZauJVzadY2h9WqeqR94igj3PA7gTdePLIB2/MN91f96Zbd07FuVPamNvYM
SfxcievjSzziu9CM9wO3qxmhYyp8bZdThdeQ4OMKa3npqKKe0zSi11DvzPcA
QrCkou2X4yQha7ukEk32JKMQ/HroNfYunUy7c1lPTo2Yy3Ya1TiGuAiVcmpF
g7ga2unBaKhwT5kn00iyCi/YkzKMThlWQohYQpsyoeSftjl078yrd033imbO
LwAssFpb6HNsiHHjXZtwIIRmDwwc43EsAcvzpakWDYOZzxgyhxDNUSvh2YF/
GhxSkdZ0A/4vJehFJsJwu3l8/KRzq7O6SnslAIjOHL77f09gDfyZgmwTiJeU
jVeLcVpdhwBR4H5osk0z2C+KQwHfOaq4nG3KHgGfYJhpykPJepuaOtia9Etz
iGU9OJDHwX5AD1nDIifrGJopWKEuy6RY49ZDdkkmfnxnaB9OMzJgp4+scXck
0TbqOfT89jErz8S+dbfhEhiQQ6RABVZKwQQ528Z1Ln0spFJtlyX4ha17iNl/
SOwfr+GK5zBmglCc85CR0AcYhtTX2EUNyKE13KQlNLuBN8+lwrKikP1alDMa
qeFAiyRVvkgPqXrBHCI8S6PylgzrkllPYwI+9TTcc39kxRKKwN6qJZul4zEU
VxFyWRjWkLX8DfIxHhBtpeo4RJhZvBvsjJ9BaJ5FS6WE7TiIS7H2h0d9tbES
9eSycgR9DkQTlz0MRNsXbJZP22rtx6kCfHrj/rcvRbPPSEjT59ytopWnQTmB
oOgDH1X/XtImnrLYeuoOv8KVNcCkl4cXNGErIkbgcGpMzW/jV6QPIfIqJPYC
0uhjl7SdhdQ9fa4qjKXaJnHIrGJVt7a4iHwWq2Wg2dh52JWsKVMuHi+mnnmd
eSZkOZuP2+9SQsCFqWQWEIoE3juYSS4JjdCS414RzvNu/UiYsNiAG+dCb1Jq
RrAN3OAYIc0p10b0hnUeW6PhkLGtXdJxPdokrti5VAIHy8MmH73HOJOeRF0y
pRBgLv/m3tyowY3dI0YIqIO3yvKUB64hDItgBZzd+0uYFrqDT04L4wITk1f1
/njmtjcsKbvYioSgHB1xKqQOwfvnJXc8zmk0brvA5bR1sYRM1rsujJ+hRSAn
daBg1IL7A619UiKk0yI80L3bserlUiVUEtwnYvfD0eBDm7ikhTTEp94xLkXM
PJxoNVyZ44+aIH4VbzbbF9X9mMJPnoukqtMz+xb2iL4OTM0eqc2N+VfcB5lY
VUFybNNWkKG84gda0Uor28rFkvQ/xH+ylRlGBjSycoxKrag/gRkSoFwpDUNS
4w4eTqLRx7JvOpOFD1XUnP2jejh0VxXzKmt0xaSoP/SGWrr8jj0TzdgMjQKo
UXxi6RFqHuc0mb1wdP1BXGV5kLAG6SZ7SIpLhLLOcBWrOqyCVmbQFun5N8Xg
7upqNmlQVRoEEVqk+rSka7no1DjBNuKx9YYr/hcKvu18gDPFXFffPooXk8/X
wKEScTUgu+q0WIhS+3SFwxqbHjRqBPb8oQe5d/WERLy4M0hIQXnNfkXCkWtz
FgBZZ1vyOeOeZWGT/ZMqLqwDQJQR3dTXZ3wxTq+lR0dtQKcJyZBtghwKciED
E6WnN2gQGeiGn3mY6PphSp2dEs0GDl7sKWFYlJYSl0OiGidXzeJZbRz0PPeo
6mzKAwtXDc2G6wK9Akbi+PKMSaA603qnHkOyWDDge2wJxEhe6W2HSyyvJ4w2
fmPWalmK25mTzqeR8NCW6+Jqkq8JV2X1uYHdk7CsWRky0SVEfVp/waoj8qud
QKcbhRiF+99fp19sex7iO5Qp/rkVRgX9tSHbc/jyuGdKfYi+k8b0EQFjmrpp
kEi27tAC7nAP8odVmd/jGJFU55uG02q/33bU/xuc6T3KoALTp0ZQRkzjvGTw
LEe0SYIq4foxbjKt7PmMHBlskMD7LqNOHQAvRb6YmgpUXd98WBOYVznr+XLj
9gj2tVQtYQva5JBQmieDw3MW5N4OVhtGApi1ejR+/pJhSjvAh/QLej9wzuAj
xDzzSnFSJdRRBqSsXShH4bCHwBKVYj3nfATepKdlhSLmEpvmqd5Vvi3I2DnY
37lAQnFDhtslZveutXwcbY4EbOi5gXKXl7E8JREvWyiqnJBXlbWxXPUHq+n3
w7sOsKd4RPTNz0paRd75p/Kyqvv6bSIULgoMqASNNzWMJ7KKTM8hMJZ21iG+
t6eY+3eEqJYzLMNsoY3hKUDbzycNTE4kFfzag0gIthvxmeUTDogNT2gDBK23
zet2Zr2s6S65I3tZjWPoDzfbdP1fcPul92XOGY7r2Vqe5UWG1g2g0LjwrX6W
CWWUjiW8ZtmBt8AcDJmCjbJgnt+sKevtOWC7Y3YfqXsJ3Kw8t81GzecltpzW
+TP/qGlsls0NRpc1ewjia0zW81z2e+SZzlBfT1X+SkQTB3AchfUCyy93TI/e
AC3zPSSDK+Mt6DuWMG6A3Gf0r5VVzMMXbJ9UIOWnVYUIwHozSobn4c7AyErX
WbXNT9wdU6WeCLLwVYB9/ZWMBfuM5v+hJB2+3QC18Pj9+m/V5z47VeMwQwqu
prsfQsdgHm1t6X98mUW4C5NDgedzZ5/J/eiozWEOhOoi6QRP8cHon99rsruW
DFzh/NBnAQL1v9+4QPNSQ0vhsK0yW9KKvI5XBoSQeg7uitHKtd9BiFXL6hH8
MhtqOKD6bUMUVu4T74t4kTSFcDHM53C9y1zm4mysg6JGessKN8gK0pS2z9Id
dzeoUnOH7oIw/Bx2u7HwOXoxByBCkjBRI9nxUn9FackFmo1H9dovFIbLgaZ5
a7VTmsI0bRNnCbCcb6IZTSfiVPkH0/ahdJCDKuum7jPTxnSe9/OSfWU/xTBS
nnEFX1+vLd4P37CAQPrRr+xBZrTHJR6kmlEoFHNDHr5GB+KayGizDFf3cA1M
mkFzzjmOsvVG9RY6Ja/86pQ3LKR4cUgMNpUpq6PJ9WztryCa5PByRPqDDcpu
CdTQlvY6P2A8GIeg+glOmOhO7/HmECfAFDbb4iFHPSnYdDk9Re69+FOby2hQ
e5wlUUqq5P3+TUZV+l0QkbC4Kwo5LSOlKVh9vI9f/gY/DgAXFflzRKdCtlG2
/Y/XzGTEKkmY/qIn4v+hQrAykH/aeWEnkivG5NnBVGIxwqlntg5AyKkY/yxv
RmTn9NRjQdUvMU0BJXKdKF10PEF+k0V7vuLo0ZpqETJIbZmJa2uQnsMaSMky
YAKA+JDtg+wow4ev64DBKAY5Szx99iliISuA6tdwYQGe5+NRNHUEcJzbT0wv
eZH11PvH2aumeGRbrcMumStnHRxJsyb1Cod8qnALU92zXoJMEsK/TUTr6DxR
KNOeWbxfRWx9fTScfWgbKZ7yEvLyvWa9Q2GZm8GzNiUrwf5wMVgEiRsMDbf4
parkDjVs9vxoHy/tZYI7nRtM7/itJRi9EZNsO0tFtWq2QNjfanJKMyHTyL+N
rlUdhqxDvF7O0u+4G8HIk80NRbdS9HhX9/0Y9BBaFpnPop2BDUu2GZkx+EeR
OeIKOHfK92m6kbXq2xkpF3UtUV1LIb5BFqsTnq+gF5BPEiFG2Yw7NN50pCMY
eAop14t84Gh2qZZdeETlFAPC7uHFsulzbm0fm1/micP8KcqUSF1WRv/B55Sv
hhRfIG5q4cui31DmdqJ3WSLxRV5ICYVjti47aY7Acq82XEnP90dzOFHk7gBg
X0eq9+viWMbUjbh7Vc9FwV5vuXVQPKOFlgbN9Lmojhlu+Tmpx+vhysbv8sH1
BVhlesMjerz4OvHPV5HjlFv6R1nMj54wrhb1NSr7sOMxqXskN5V8pQmWgeZH
BaE34OoaPffl9/URZOlmJWnEO7uMAi+th3XK5YGm7wSmXqxPzIXTP/cHFoMl
R9Xfb2/0Q2JY1kFUGPe8LHVcS4EdW9tD6XXkeeZap+J2AkgA11vAyUTcNEBI
4xsYIj3aC3EvQrBPgT6G29WsmFOV1PN2zN2YvxjVS8K2vHH6/WigiHWB2Uik
XWddUKfpQJFv+UxdCcdw6w7nI06T7NqzyH2+//JiCVUzvM0Yqtg+dck0kLn8
MFdJmJLYtevgqhGAHpmOJS98LKfwZXNVV2tzKp6qyHrvS1nIWzq1Z/JcC9Ok
JtRWC+f5XtjTdgm+ZI/tLcnjBmLsHp22djibWj50qTr+aWxwQkgqP2k/ud7y
uof0igwO2TMjB2yKqW4Sb5rvj0lSMqrz0PymXGVXMYmnaYM9SrqKvhnaCPdN
DhrEY7uJ9wNgTmPs//mVJ7G5RCnctFruAaXSYsq3YMxyBhWWGbayJtS/ojOi
dx+7pDENFbFf+XuQ8Jh0V5TNhTDK7FTKMpWY8xIdOF+dIrerYSg6IXtFr3sF
oIsahoc31nlQukvq7gCrJkcNQ0dpSYY3TLGwnLaTxZdqgVBtgjQp6AWD02Ul
EqFoYwxVN2aWbhf25lncrmndChaXgPi3VEsKlId5s2UHjOYzqvvqo+RKIVra
mTRl83ujxHvMVEuZQnsYmGjJa2eECzmf4kjthWnnVB0wVk2/pWt7hEIWsUiW
nMmv9n/Ezh9cDgmUju0E3KdpWzA5EnH00xriVVT30/LVypJbCtpDZ4TbBwa+
5ZE5yaMw+F67VsdEoigagVq9jAWCLAfpODfQ+tb2oJwvvDxoHFkHg53TYKh9
mK+GW860W0ZyH5v+ZhTl+gLirhULwO5Z+V2LbPM5D3DMCf4/TLfzh8WfUJLH
6f4sxMZyHhRSzzZlb1P/0GwZ2y+TeWN1jvrnInRMVfmvbOz7kXpbcss1E0l9
Z8oFPM/SsQaRM/8um34btdWt9dCb/DG2lurW8noRNuCrCiBIHvsSyB3o+rA0
nbTCvRuI1m2iM7O+Dp9GerpIKv2VktXoJ75sfqv2XP0iA9DxNMaaXpHI/Q2W
8rVuNuKRZ5EuLXvssZJeFbQB3HKvjw28Q4evScKh875anxZJB/ZJ80Sw60En
5SVB2LDTeKmtB/E25fyc22C3yaarewjPvX5x8f+HFcEA9nTxtTJxYhLl7pur
/H1gwOz1OwAVDGEBdHQpoSP5Nm6/kzZB/ODDOGr2NJVPsIrUSkGxryr2UQWx
cgU8qK9OUFnajjUJKwz1Rt8JS7lpmG8EDbecyJIuRUwI4HNUCiATcE+cwzY4
v/m4mRks8MKNXLHbENu68+Ph34zyNAChOiQGp7gFWIcf1m2T3kaXuT64hPBx
xOlBNd7obLyyT+jXLA9ZLjVzp8tf1UHQ0so6G1oVBavMkt8YhY8IUVCfgp9z
8/wfCv9qU6T8ykDyfTquEKO05quduFAugNWfQL3ubpLY5qmp7YwV/Vw8DGyx
nnH6uasbHNW5rDym12dOMDJTNY47MAgM+eVjlqqVe//NpvQESbujvWU7JUFP
1NLwrD4AFFOYI825Xt8/axL/wk1iOKdYvEg/MlKsGi9WlwT36BppYWULxOdH
XokJlulWXlRgkITSRcUyysUcwp44J98LG3Eiuc1YkPj3e6QfzZNkNsbR4PZt
OM2mVZOyheQcF9ruHwqIGS8URAGNyaIjnCOx/lyv5ZzbIdf2Wh+RrATdnz2Z
cDJseLl57py0PbXdYy4wQryDkqHirZoIq79y+3pbVAqMn+7IRzQSP3aTsIQ4
x/87TeQRHkmP9y1tLSB4AV8001vVcyge0AvsN5ZQ2bymuVIVI845VZWHPCDq
s1zAWgPU4piAA9Q0o1ZghQFk9yI+QExxBT3rt3arGeeS+ohZJMiW3kZZrmhE
jd+fHJv8guH6xp3kpRjTn1Lp3nkyrUhR+6zBNO8T/vvwYU47eU4PiD17xlby
au5q0LU5PRCr3Gb00Y22xAIiP69Yk+I3WxGUrAD+8KUKiDVLlpQejQCLEem5
h/9Hq/h+rAp2VJnuVQeMoxeBPLP4Xx3FJs/i5PWcS4Ac1z6szYrJjEbxg2W/
XvYtyuMdCJSFeyL/7r/9HRl62VhdekjWXROfUy0zEnfk7/Of/Pa0Va5WzBnt
RzX9OT/go+zjPH8025ivXuyyVtIZY7bPCUCA3h4d3eN4pdcHsyojNc3foht+
mTs/ZFBLfR90vGlCfXYuw8Y5ne/BndS/MmKUX9T5Kr/kC9VvuA7T0FbFBCgR
oGOzaxzOb0Y8cCM8hQ8Z56hBQV7J6gi/vHIDiYjfcC4L6OjWU9AhBb3s3aQl
49vp4vUcwzDAlJTbkE2d5v5sBEmgw9R7M7kQKNPyacugRF4gEAJxuGejJzhk
wBu9w9cf9l34yyPfZF9+VlFeJUUbMbVEUkV/ZPTQFUaBr+7ckToNGFXSXtZO
L/Y4H32qQhuSF9fzxgQodF6ViWunr6f2GSltjTTzvWrodoXRFh6bH4G4Wo4U
npK8aW/MEQLrdSHxXycbZeUDebAYSrd07HMWRdPCqpUXB1GE78LLrRq+RHvA
3qB4LTEe+93mmsrS1KspP0AiLZeMP+lNTGFEBy5NNaDbGdJ9y6kXmOANsrCZ
Kl6A6MnDTVkzexIi381ONM1jvyOQaCjf4A/zXAlC+YRJIpzU69uBtRj5GCqy
yHWQgOVef2l6ZHSLRkOCqUMKDQgpl9RYALd3YuxeWhJb7IA6744kD9GUXjBC
XyIzgoWEBFv1tDpbEtt9Y4VqDsn9+A+fguHxpi9K/1fqql7c6xDK3jwSk6XI
n/9iOjSvr2IP9jEgg2BQN/sosryb/ZL63a19e3yjaG47EMQparLmZD6CPMGm
5ns1ccViUz/pUKu+oj7MkUvrVwU+z9DJckRP53BmaJgAt8JAe3p/qeQQwJZj
UQtAvFVoYTxrZCpT58D1slxOx4Xeybl1NCdgpSXlusJZ2r3xPobGPOf4241/
nm1XdOPeR+srUywGMO1wGbFYYEhNwJrEapZ6RAhwB7pWzIRbpB2UFnYa312n
X9cnfY+Nl0Bk4kMdyNgLVhvpesjw00j9cgPOaC1kSrB4zAH9KA6fsEfdc9Gw
l8o28UyGk0ZIjwS+bxkj6Kc4zZrQU7GmoATAJSv53E2G/n3RsdPzUvD3D10W
wXZy+2qIe8RGYIXoJ259bDz5yU4jTZ3pmnJmv2V5l2BeF/CZTCSDCvdEgDfz
DAcHGzZRwP/qHmo3UevH7kLYIkDX8btDpjJ3td4P2F137eENFfPtbBDSxxNi
VBsvQnexRzh1fdw/m/apqreKCvL1gsnu6JUlyDr0lpREZ7ZpBTn5/2GSt7g4
4dj7RfpwjdwRc6MoW6wrRuwScH5DW2cdJPCX9E8Jm1U9e4clIIxUPy+NUHcJ
uXdfxj5WG2/837kzKbeNvi3kQ30gEhW85QbQEmjV+MrzwAlhHrdRIMb+PDZg
RoQ99QoZJO/WoHluc8u+/BJISSu7RCYx7c+iwc+LBmDJuSgba5CFe6a/s8lC
6dqyWMhx2IVX8FlKrXvtXM0PeajGsANcvMStThWR6vfeb6FQak/A3C3QmmIN
DQrOcc+0TB66ocxoPfjqen13zRY0WqTnmYJ0GVlsdBAjdisQ6dNmDjk7nxR+
d5HfSJnnTEt4pc9FLrmyu0sicGixx49CJwb/WJMSgqzZx0Im+NvolRz+i9Ox
2GhWnynI/u5kH0y3zlc5Xc3ZUuLPdTPI61Z/ZN5sE3WJjhftCYoHtoM2AgjH
CujtZa1yVEyN6gAH2bsbAKP/zh9lyIk3afilrAy31/melSOVxALri5p7gZ7Y
z9QHc6TuA/wIeesvbIrh+B6rK6ZkW7khCX2JhTvbDWm1iml3NiaDG24yVk0Y
SpD9pLrb23RYx3CBzPfdRa5M5cCKmKyHXCfHJBXNOxEtLvx5hkgcfdRCEJqL
7Uubvw1bWyJMNmEjZpVRGCyN/lAojwV55jan8qVYwxqJ3lPFrdZFvPcWEIMw
VfbH9yrslefvH8uvmnrFRhF2SK3TxsTiFF63W+jf8j9uiArNFogYgeRG9qie
/YbcA02V20EXnJyKpkGPD2T4JgwWqNQjXyC8/Ehph1GdwVNfSMKWTQB4HYbG
MWX7o06QzGfhOZgpBjSyR8fUOhq8AXkRPt8EPtfCNG86xUD7cLfVzyaBA2JB
PJ7zodNkjhMpTGVvnVYgL0RjT+ndJJnkdLYOVIH7TZBboPxAPAC5QxRpBVir
IlRcX2O0bEbBaxLXnuHM8COVbfx2jGe6EMnIkMAwYKl9kyOH4AEE3hLBVWkS
9HfuQmtkOdzDzBh4xN8jK1KxsqRG/TeIAVhc4ZyaCj+SWPo60NQQXisQNPe8
PmgPixBSr/4pfwW3Yfi30/GXaWQBxZgJpbBo/1PV9O08aJoYGssjiEzvSfqZ
uVzHlerPEa0TOT/oD3wPVF+EZnS2ggEUsx26hqyczNMWL4IC4vTt7H8ucK4p
uBi6jAKu7sLfViYqWDuHd/tsW4zKKyfWGF7MveIaQ6Cn5AzOl/BL2cAdkVmH
v/wYxP4PJe9qtEPcvIP/OyDEwi1L8vNxCkMpvnxfaKYlkwRf7IizKGYsvKjL
XgLd2NVl8QzVqfbXQAaua6eia0cvN2u0eXicrmGSlJodMZfGvIysLPoxibF3
+M/OtumpZ5tbq2enIICdSLQAXyAVRNMGYSv9YUHulI+pXKhckg5XPhOnLloO
Q+qAGPym6N8b7Immvwhk5NSYDXhID6EGx05Z160MbyX+5Gr75D5RCnxhXDDV
7YhQQSG4KP/87gt0Evcg3n007uOUZBkd2cHB14lQ0stJBThwrArzhoY4YL/e
HnhSlErOnLWYMR5/2ln5ikCeYe+HHirqFb+q5uuQVpCUlWblIMS4tJK/afvA
LB0W1HaLmwQB+Nn5qZbk+nz2lX3W+93lLoAmZmfdiSSqiRR0cOWjmGakAySt
4Yv2tL7dEHTLrSypOBFOaJ5ZBjjWF7+czwccVcSGRPH57/p+DLYBV9DyTzYT
vcIL4mv/g4okFw633NK0eq22dEAI5dwfkE1AjD10neDGh6VRfIcwVJN1xgJz
P1ohDn3gxRBHCF1axYSFr00SQSk4njqFrK3J36QzGEjQ5GRzdvIsoydJkXXE
GPex8ZTNhQw/MWzDMtDMu+Lfi5ICHeP5K9IjnR5B6d/rMWpjOuDzmoGoIiP+
MeQ2tnea5qVS5tcrUbB9litD/O9rMm0GSRnVNELhGhbMUxM/JEuXqqEZgjcb
mwXusIpi4EZwkcd9hSHPaJBTpisywJkIK/QtOy/eo/O5sivSBi5tbU9g9nMd
2VQfvvz/vBmgePYBjGMtNSaLUT3H1pnE+7dRPBAcqoo01JWWk1OpXQSNr87X
ti4202XKoLIMJ6eYL+IXV6QQ+HlB5x/7SpMoRg/2iRezYda6AOzuK6Nb0375
IqHduzNMT3GIVzOsIQ5cF/lU0B6nDxxjt4icsQeNeRH3Qd2gZB3UY79on9C3
BuFS9WHXsnR3InQ/kxEokRaXxMaqPC7AcbK14dyneNhfY8cWRvZX3e/Y2PMw
XGn50MXcqKZR1nvg2aHGZWkPCOdrJHktAZIOkVdo/4+EZCeXlP50Q89LBKGS
GSt4BDdrOsO/bi4FMc9p+mbMWB21Fj75A526+7ncSOksVz2jb5tPpKJzz563
O8cKuZtMj2I1tjoTnw+1L335Q1vgXSuXIWZPuUIuw49/WJWXl91bozGV5Ws+
J0PTxL/JVs99y717RRk2zQ9hVaf2wYLcwdab4b5umkYT/YDSTWs/assSNanX
tGVlMi4NEWhacD3XfWQHvv+cmuOlpvW176V5V3vsDSMVv3Hf+36bpAcf8rw4
2V1Dzx4DrlGLG+v4vD61YFBVSEteJ5x/L+FaRgCxEgj7cmKTISfGla+LUJoM
Af8OB3GfVcNtzjtmEpIa8KXWmANRbLXQcKzr6tFbty+MxuYTdBD71rGFZiNA
xkCN9csU8RNennEHcN3psWwFlgsirNlY7NcdoaNFm8g5IBK0UuAwGOvX8+p8
Eqleuvr0EowDPXW4sNhiM2X2NmyB4cv9gh5ju2mVEbngUGw+QetLOVmsMIqv
c8XzuS++7tsnYiRTydhNXX/TU/8bBoIWDIGYfKc6NeYekYyfKo6q7eMhsiwd
kmkE3wFolv7U9gjnQoAIksXlHYVg5pY0jV6PtcMGgWBg68ms329QcBtXUGUy
Gnx5qNDvm9m/AYElrae3iPxgTcNTAVrw9s07ps+08ETPr0/VdyOEu/pt3rfi
s1WpMSt0uhPWD55WWw0Pz33RroUPWsv/w07+uw1nKE/Aoejdx1ylqkK2C8h2
LrVr3wXud+IKeUHUryZDBhzj7Hz/4ilrgBwj/RaZF544kqp3ltTkE0kdr1hr
DDj2AmAkOCtX/598KlYTUOpC9s6NTEkK403KEzQAiESTOaskraMgwh0CzzdE
T5KnImfaS85AKsEO7KtSusn9gl83wUgLax8ba+xLJGEQUFHDw3wh1EKgiZJC
UErci1ZbRB2EQPQ7JV7lKSUpYq3ux3eVNGmGFRwRSjN+laIq2faDmSgurVEW
UI2lp9tF1RleVQz5WuUTIA6/ujNhAHap1Qqjj054cxppbtoYrAMartXnOnSv
VyTcdjkW9KWfO9q2UpsvXfUaOhBZly837bEaAQRl6iz1pD30nbGQtY8VmIjD
Tg2YGMo6Ik3KRYGtTeBmmifhkBIf+AQiffZM3VnokulGEb6RZLreQQR+A2e7
kBZITP6a/ScAIVmn0H9+IuMJVgpyTHtzr39N8KVXxFmJeOOpXeHCXGKzChTC
B4XEvqQ2JrfVsAT5VClvf1ZjAV2Rsl8P6y6F08muRtJfDYKznKrrl7WM8RMk
/9e9+tu4pj6NaYS2sh2q45EnGR888DEKyS7hdLrSB5ZeV2m5qdDF5ZX9BgMw
CoKGRn4lv7SG53QfZfCJaGvpI6nXypTnOR0WiPGuSonl/u7OlIqHLyEPhH1f
/r3OOawdwAXlsvMWqX94dVY6lTVtRM9mM1BfwkKRyfs0oQSibXP6CtgjFLB2
dY49nL8ejXd4cEgBz+cmdv6FPs4ozhBrytXVqZMZm46dFPCyhG0CVV5jd83E
cqwG+QpdUBOKG6aFIArRoELjPN3KJqW0RGTOO2jmszMel4dCmcin/m+arr/a
hZWQdhl4kJBE1ouzOXBVoE2VE5IbvzNH7dKnLYkZhcBO2I7fg4TquwdPD8j1
phopqye6k3JAzmrRxgCdwc0QEDh14gQeq4XhSfhDtr6T5OEWqrBj9ebmXnGz
YWm6uNGUY7C9iITUuwKXyQtiNb2BbnRzX0EXXhUfyDJfm07rtgfkRvFt52MD
Eiobk0SQzIXwMc7HqgUqDm7uWhXzAkEwCjkZAEQr7QqgnAGa2WqCJ3ZGJKVm
2EV1WdCZyP5qpXQSttmV3+QUiEY85EduxvAzeYyJyufPb9oE5/A1FdJAsV0z
w6O027Yn9nGKcic/T+XgflAjmkw0/q8KW6Wt1k1syp67Hkl2f1ra95trjKY5
HbEHn1Vu9R57yOi0kGYpxHePnOq5KXR4yWWzdmsBYwOjTOqvaxEkor6an8DG
M8SYoaIky7BhX4Z3eGUB+Pirt/wWll8YwBGh3DMnk/TBb5b1iFVOST0TWr1q
rYHN5kZom6UjsP/UmT/xBQygufMbwkxLD2UkW4cS6ViL/wUaq3nmHPfGD1Ff
RYlp0SgLFMWSAcDqA7Sfjz0EO/dVG6YpGtxVWyD6ui9bWNe35CWWyhKYeVDS
fiEoU5PYrlZNrxyKOtbR6s+tM2gh9PO1X0lZF98V1Ycy+hvQjGNKHPOFM690
lTqKX4TPViJnN59yr1ZAKaJX19vhtzHiQLMdv3xaBNN/Hf7Vkzxr6rtUEQni
3Ag9gohAUaMG1zofcOe0wZypp/79FuFcDEyqAl0eNaI32oDWJnsxWaJKZ1mn
HIYaFlVYCvc46E5DMzsEI3/8q2WlMZjAsp/EyiYLH3ckYownuS3mX9QhhIBN
BwlnqajFO1LxzwhBZRB9X/WJrpkzZiOh1vXEO1xAhUMfBOxH4Bw8ZwXFSHRu
ssRpeK3Ky/bolFyGCEOL+fAFxexs5T3NS+FEUQ2gJ7EROCEOGWw/P1O7bNFi
tv77KKIMhaBxo426wpRMC4T5VMClJNZSDetEJz1TilSjVCNdV7TWka5lRWGj
BHUmtKU/jl7JLpumI//EDbT3hoXONUYDlA0rFPnSWxcz4eDQEohLw/zS52cg
VaHb85RxUe9iLZB8BR8HBBfXfAt7Tjf16fShsq3Sm1CHGx5nX2C48ynAiCJ2
vH/It/EgNCOTYq9E58Q43h3ZY3X4+3vGJ52YrV6PtlMPq15Pa+UWyyRaUtL0
OnUaetBO6W9ATdP0vryjUccjs9Ro+uCA34Y42F6WqasATa8R2GkH+IWqfOPj
RrlibZfxf+rXlPCm2XqxFpJnC1rWuUMO5nWhj2ZAgjP5fSBqHCADORvPPlwK
/uVVB07xdIjVUwgV83caMFktUqSoEriZu68rxn8/i1vOGrqq0IOWutpKocny
hGcWOVdhRwyBBWnKZzxkDgFqG497LO6SogmmHPP0XXbLUe3MlnXTLpC5MlzU
UjzM5PWar3tW8kYz3zR3DCZjNY9WloOKDfZf96RFpGQWeysci8pDaTGBGssP
pA7IhSrVXOM5ozoBtt6OQgoLPWFSvuhilMjcmsA7Dx2qxPI/JGM66wz5BZRE
ucBjGhu+ZJZF0wMWfvvC8xA56r95B8yxT/duHYbpCj0l/9e9/udzvx5aF4ql
TbiEqRI+YaJf7tiUDuLwmEI6dvz6YuMIwQp2y808qtHOaIt4hEDyuxTfGcli
/dpL/n4ytOzq+483o36lnyXKBig3gDusrBiPM+/G4FSBlgxVy9t74W5wzSsx
pjXPozAXzEFU5m2KxGtNTcxZba+aVQ5LBloVVGj1qz2cA6MujoR1azcVbAMN
hhQYPXxf/JVQ6TIxb51wOcH2jW6HUIHpfmU8So6s8t5Syyfjoizu0JgqzO8+
qx7Yx22TukzRIpscSV/H+9sVgL5x8GWbJERrcNvna9yohMB/DdHewYQFp9o+
0Qc+TXRMjLPtM+nED4AZ6T+u1SAfMPeKspfb3Pu5G0PtmE88yT95G8DWzlpo
9eCrwNTTNiVYiiriWLICqj4mTqNmuVJp7i1nHDO8gPW0ZTW4CL7hQP5MpPf+
d7stG/QtpaOWMEJFqGY15TfSwgu4RtZb+e689xVBF3TnalhwfCmpJnj7Riiu
La7sS+SqSxp3yTtY8+MIgxHrm62T+r8d3TRx/P0aPYpsH1wBjQ7gTKQC5cRR
DpNrqViPGh8cVyPrW8+vtKHAji8opTxcS2sAvM8Ua7zcBtn9/KJJ8o5hYSCW
u5Kk8gMy8AkrPs4Gmx9Wc7PiYH3Sc59WHC9HWj0GgiupW0L1lrNtbgXbnzSc
QKLm3EM3eDc3LRjRavJNpdyUIS2nISsngQanZ/DFN/SYb4UukwFauFrGZM31
iOJMc1bEFbWtEzIIrqGNGOCsnpcKAQEpdHm1hcyC+er7lGw4njvHAk3nXsCK
pSMlNYs38f9yHf1Wuy/qur84HEjSIOi6x6bFr9PNLO5SL3QfR0VPZRlo2zPI
A+D4Yhu9Ds6s/jGXJGvY5A1w5ANYUgGuqH9SiO0C4+Zsi5/ZqTZVaDFn00J0
IDDIHWbOK51Wv7cU1D78nJKVGalGdhT9pN8n+uib+M08QNO+ojccVAoQY5nu
TAqKKqXncvlrj/iFZR30xcMa0Ld7dRDtU5RH/aYuDNp20mZ8CX3b1e3UtnKG
IVHMjGrHrmFlhoH01TfnvA7Y2cUrfXONBmijo1igO/sXjvvayg3q/A5qUcE2
kxlEl+eFbo0rl8usjc+ZrwuE+BffAaI89KnzLiY3rzgWNsBWvTzrMjc3B4IB
QREYoDACGE7fp4JFspgA7urrGAbjZjGIj9akOUZINEHSnM6bBO9Bzimvbfnz
Eu6sRiFB15TntjHs32rb9zrf9OB8G1RmJte8yUeV+BRNAi6ZzSXnDKAKCQSF
R51UGtQYqBEvkmjCnqvMVZg4YFgSC01yFULjqcRtgMAIcIQdSZ9bPxPSM9q9
xKhCALbZjckBNop4iJIhF6Uo1CEU4EKzoHp0X+1YyQr28q5doeUA5yLYn0ZB
RqoaubJekughTSoycnjnFEs9R2c/+uqZuywq55JgMlhe5kekCmILQP41cTDX
4p9kCcOhqnhOgg54syZRtmZIxHsAMpHVg8mdzQSwrO73cRRd9zOK7X9wqMTX
hajsykf1m3J3hkcGChp+Bf9qTh/z+02U1wIt+27oRqAYPCHCusKKGZ0fiSyA
jQrZdnDsyQMp5xthOJlj6faXTDKuom36LHuvRtJJLnY2S9LmW/Dv76Xr9PF8
LTmLxm8BDET7Hipdlz7IIUFOyv6ePIiGSpm9Gq53jMyLKzku6jbw7cPx+iVv
YR3SBGraFFeIBUNKOXTs590XMbKtYRUhCf0w/n4V8cw/UVuSOKiF6JUEx732
bOiAd1mSAGYVVtq+K3/pGM8wfGZd9QrRMlMr2WsTXyPussP8iXFYYoULg8aI
jsjAk+cN6hdWtZ+X799mSaL9NPjJsTElJwK0Z6lUnY9VsnEfVUUlkO7F4n9U
pjQ5C8oLe+OxYjSHUPn7HmSrTuP2YbpgomautvIyDkOTGxBaxKCxUXUuWr2U
gDxNZ3AGatNbGq2GkLD06HPPQOh+bv2FpEKoLQTjcrQeX2BsisKFPcmMD7w8
S5VbkI1upTyVngXjPUTqqBmaxvlV2lRuDAaCdztKwQnvFKF1RC8PAWYxpmU7
PinxvRTJFuy9AvndY6PJBRHUYJvnMvPCd/YfqIZiTRo4BixCoCNOGvDcQtdq
Z+TgyyF/ATuw5MBXdZ4RQisJbdouXOoz01aKKGLUCisJupR4fYROw0VNnKPz
hRAc+3cCrO7l7lYt/STcsyykTJnK/TVjDH9C9c529L26BR2LiXMMu/Nmd/fb
f5Tk4j5qTIGO0zAjVXI2TtQkkBi+/BERN/F0MbziA+dQ9Um2f69ngvL2oBzu
vWZdCIuJoTvZc1J+JiB20CatTznl/y7lhbuffUOH03h40sp+tZVRDazyQpa8
cqZS41Mz+TSF7QmAG+e+9aFNa2FMr2dRBR1yBQN/BYTpl340+pYyWIeVW2ru
na5eb4b0NCkLbO6af1IHl+lbLcqSw3rn1Do4S98bHg1pfeDuYASC/3lsbZos
h0yt8fjlIU8w/NdVShHBDePc/xdKg+MgNP+73sb8pJbsAXy6wh1F8Ei74mR4
hJiai6PzQiiU+kVLaZdC8hzpEYX3qkJHZ83FGsYOQ1Wq+A6knQUx3shxF6rV
B09iC6V0HzAZfJH6psXwOFh5pio+58wLRXKCGN2XzQm7n53LbAcArCX9v2HX
GPGGSmlc1cJPm0nb2AdSAapA5iYVqIL4uOd+eshHP32+3hPqSnblTdTBthsF
gfJlYaowQTxbBy55tMmuwcbC6zyj+SGxyWM+/DxbY0+vciDdQeVOAuSTnHvc
lJMGraLHbLAN9EubblPL14tWONd4zVS5W/pOEqzR/cYwONuOXhPDA9dOUwGZ
yocaWDhcaGU8ZJOr1ip6jRdd6kSUdJXNzypPex7CCaAXyFvv31FAwE6kyR0p
CE+fkFP/SzoO5wVfoIHGlQbR+0AUsGbxHAWUlLBTd5NlMoctsVgMvVh13CLq
rgy8XfS1maJ1gM126/myrYch0zOM3/p/ZvaLEQZ+hHEWCl7MCiDt7tWaEPuq
sNQ30ZVSX9NLkSKV7hiYoKSpVZ8EYMi8tOiGisS43dn/Xq/oUsWwhjH1WHGt
vhexZGLBKmJmeFeSmV/dZ8QTYE4ZnguiAhib1COsgjakZ8fzTSFvPFM40h81
yFsunm/NbuGlkW/qWpQHncuokJZ7BHQPXTpCbzHh9Xlyoy6mHAS91sl0tgSY
hKip7CDUgZ6+E3lYREzuap2TG557Sfy4rNCGy0fMNvxfR1N4mets1gk0J9gS
hmYMhg9THCCdknmA80ThVHTdposqseQfynzHjWiX9jlvS3UgX0sWac/0BInt
e99KXG6g9RrEsBFN5CbqnE3Ds2N6O99Lrl57UyBAjhq3+Cs7wnnSQg9fASfk
jG97verVKr1wJPurMFD3OCEzX0useRg8S3jENfAPY+1ClunRDhIURuDAxfX0
TNFldd/jiiydopgf0AGZKmL/kP6GHc221YjgDOEXkgl0VcYAs7xdffrLEmRg
g5E8/AN/bO+hOfoURNN9gGyAUn1/g5mW99V2l/ZmerCmTIkIl5Add2Oadora
sDwlg7w9BBmVfi1OVy03vzytoJybXHoOhr1yoLTpQB1ZFOoaIsDG1K9AkQ7k
eke+fF2VcGLjt2q4Nb6pVVvV3ZGA2W2n9/2sMM6UpwMuvQFcfLx7u/UOui5G
t0Zv24CzFjKjCTkqwN8kc2Emi7pYALnZDefrWRrqZjL+M5ia7pI57K9QjUuP
dXZewQrjQTApGqy6DnizhsnclZRPhtm0ysp1CyM4TkATqa2ZAbayR4tWC+Ie
NG3kC5XyC1UsXElQN8rAtLUJl2rbqvE2nZs4OV29UV8tFNYoCw0sfm3TqnGD
ip5JyBcRDhc0vN3yUp3zWm8XBL9Zr1ZAgbBNVW1LvJ4YZD/Sme2er5drOzk1
oqyK15wvPRcJ2QQKrPcbCRwSKR0OlvCDVUV4dEqX/uxS0ReFE5176Sch1tGJ
wjWrhLCMoQR04N65aKxMYL1wX15V+rodjoqlexWvUUmbXrFx/RAEFyk52BLY
/3r0FeGC+UMdTLbJ3V5TASW8RS8wabrEQT8pO0riLhzzrtU3Og6Xe4Pi1+cm
KneRIURyKlAgXfAlXswzri4UwfrY5IAfusEU7RrapCb3Z7Bd9UGEuYpTat4O
OR9QKyAdTq+5FusVdIuksOfFmn15uE1rrZBxs+jG3nDHYzHfQBkqwBM8OXZd
Lu15sSq16+izR2P33v6qiX8d2Z/gzW1koEe/k+w9FOMp+dwqutMyogKd5ZDg
pTDEbtQt+6hJEgJY10sgHKcga/TDikb/geC9dtN+X6Jw2B534OiU+4uN18t2
nWBQXkfpVXT7gJtAdR/S4nUpkh8YUBMJ+KGiw6DCqvCCqKjioajrv0YhhBNm
kDDLUMpa1lCDJJLvXl/YFqbnbQ9z5kZwDjeGTzThV2lRzl3clO2drBSEmKBy
PQtbfk3+46rDnEioAZ3PPen27uXMFmMz1OMrEDTLbGaIYuhs+7YBZUgCEfVi
Kw/UHb2//BSK6L41MHj1ZVHks+xZbdMb82zpYl3UpZcE+ZVG9dPFKJLaeZw6
BxF68428U2F/KiIG11OmAc44Eh/YiBl6b5l2LRozbSQ//FwbQmWT/4d6VTpB
tGcIizJ5o1nCUr9GCuBjeYPY9e52btmPVd0lQQCEhvho9N4FlI5xB4Ebw+j3
Oj+pYQvf0r6i9++hrs1Ni/ARRUXOiDZOdz4mE4AtlcR4vfINijIpSxtlP2QW
k5Qk8XY5SeDL1YP7Va2PyE/PBmPD1YeO/403uDaBP28OWr9V+aATipQpE3Pa
8llxkHxGO/XTwuvi0dG0g4YH/hzumplKtKfXM81XN7eL1PO/wudRbUn6hNBc
DxJyveJXm8sxOEFdo9KL6p/wVBIhS+b8SMboeEJUWBv05/R/RXxTB4USRezS
51OpIiSHK4T8YfAf+Xlr7vCjOwc1feunpJTRkcw8CkG5QtThp6bx2klW6qZ2
RF6nlbdi3N5ktqLPlfe9SWCWyhYpzDGg3z9Oggoe8myG46pKUy8r2VUnX09a
pDAJMwMNe3wLJMBnaM+v1OhlKQZDrmI75CZEkl1zPi5hMMc78E3CETdhV6Qp
lnwoV4r0JeTjFiq1ps52zHouX+L52e7vyOCBtRcLCAGUIowdVtc03PrX56Yr
b9N+bAqevv6RJgcTLKFdxBZNsNyLeOjnutgvVoqyxpml7KGMlHjdYlEFoqBE
p0yr91y1s48km7DR3r4mBjFs08e6lV+W366I5eJHfs7cRkQ7Aivp7h2UmTzn
zDPH3et3bqw+TquN1DLwOmcsCrKAfjBRs49434Xc8bjCu5vknl43edb60kRX
u8ZrQTTEkFZo8i68agz6IpqAvdKyrR4TbStJp1BfKLsN1dKUvGYcmaXtmSiq
QbiYnj2xgsfYVSm3sVp6t5wOozihOCR5IeYdh0O4PSexT6YGgA6F0nff6TD/
SjvcDPHOqgUPdLIEZ7wRJCVWGDSGTSHty/QpR3UUOqCx33YnLkgYRY5WLZ0Y
Ldrv+OSQkqKbvx3SoTxW6E5suZcdTxapdiuTmc/FhrtVZIVX9Ryt9X1A1vOx
/M0LZX4quGvtmefRhDjEfcO+AraceGkV9P1qkA1rkEjqymRoKo6TFZgnrtUr
HjtAR7mxhNRN+euU7oW8oDDD3K/f4SStIhN+aSpzSw85zyC41RHxrUNB1pc3
Dpd31U7GAkIbb1EUWUSKLvqAyKM6YAgdndU5h74Kek4BYGPs/vFa62/pRtQv
kqntf5C5+m99LN16cMbzHGaiQWaY8RuXSaJdsqOzDCvq+0smxa8oRcb95Spj
sMXceCSGRCYSv8J6fDKU47E99ObuCmkspWN1XeyGVqEVItG+iBevnJ8t6dNP
Dka6Sy8bauj/zdLOB6122p7J9dkY9YuNXUNMkeX5VTMWZg/3KZzqOVgbBhKm
oNplUpJH43YkxheKHtLnG30K/EbBzll5CTG12oz+nfqu7zx/fNyBuKNl3FyZ
uRkkhuBXENJokPdUt/LM40AAAJ/u/gD/HJjvzvA8GklDesmRDpg9aTLZEvv/
GDMm1LmMXCe5NPv0nd7oeIvCxOzkwN0wk1m+1liACL64cWbTcBtM1VuzFVEl
bLjJsNDY9X+iJVqDgIcWCjNpkzpr2JeQ/4kXk+d88ebW63KzlMa07YLbT+xL
AM8M7mcD/ZhAQkPflmVr2KBAVZbw4sOn2e99iQPEBrkwWOATso/HUD0psg62
0JdvWLFrGetGJ3xm8B+6YnTLvRzfx081JCmMl8BowN3+/WZyj9k9hz38+hH5
l02gFJukvG2JVej7jX0duHZGTDKVT2dfjoUqFzEB/TzmUAMwUYJYOWMcWAVX
z0EEJe2T+bECMhBTwT5VS03G3NgsZ9xub2msc28b48AFCbqEZ9b3DxmvN9lU
tCowN74KypllyhY3nufyWIYCHvcPWf6DXTJ+blQluOdBYJm5QoboXuDDysST
Q8Wge5So6mVYFNqvjnP+GyDCO/UNCNgXNUCQu7VK7Y6UWkEBazEJGzvEum1G
D88orkOuJTe0vflSUDkBj8s/04LTyl92SP7zvXtkenba1mwWU5y+UdD7ghCt
JdUvsX6+IiAXCf7eYU10mubj9ZMEuchIzQHBbfekCHneeubmOPZhyP3IYh1k
Jl5pgteLQaZsdU8Oqm4X4NsDoVpty4gTQ49bgmJyY2Vwsm54isv1cN7BkUbQ
e1Ur8rC7VDzaySWcMRPsfdkb0d2hXIeiox1lwc8ZWUdZt6fVo8IuI+JwrlAv
Qe8OGMYlWcU2N7soIA/V/EuBeyqsfjZ7Tc6QdK8s+qGYnAx+o5DfZ405TnYE
5FV8c3/23+kqn9Ls+eP66yWMrvHpFEc3XoJ7Bph18hbmwCNLWGw/zAZGFcDW
yLOgrdUcEqjJfhjBcdVDJGja7En69PohjJor+BkCXph0EWprEw3eC8pf9/+B
+ng4upbgz16hh4/jgCsBZd6/xiJnIIy6m2axpCvwQOmuY1cbXWg+Q1mzVHPD
avLKVmr56HT3melVouOFzVPrugsaAnIWkkOk0KczVkmWiwqeZ4th+uI+DWI8
CuAxuMh9v21Q87JMnRLSwffbA1cMcG8DlmRhNx3Z+Luhlcuvd/e+2ftAiV13
r4sFJbB9M235nnA+dP1dt3vxF9MzGNlDXwb8/KEb3afrYBB7T7wfZOKsIz2o
acU3gRmlBB96M9zLfQAp6Q2f2JljSP1U4HbsJMM1c/PjNzSpW/hQNaWOACMY
5SzdC+Q8B9MOW1pghu4uY9CCxOef/0ARbiohKMmZ51POw63r5DhVe0S9zQu9
fdv/IHGw2g/Q9QnwUSCY05SGIZAmsktbidP0SNS5sjRGf94RGLuP09KvbtBz
FDVACK8GtUbzm7UsBI89xkLacOpFWs5/h7Nhjhv3e/M+ZbtV357grH7Itij1
o3c8akdFuCHr/C3F75dRnZ6tuCWddiUzO2E+c95pN8n1qYeh0yUrmVp/PMyi
6Mx9tE8bEJHf6oH9QQ5SvuD/nPyEPRYQDbpu6gE/09QqJ8eyluPxoWgFlrgE
SL4wSXjBsag3yW7xIlyHSSmHF4kA6n2oOPso6UaGF7lGWYo+YUeiN530Ecyw
0CHAJ9wzeiGaPjGpJCbkVlj/wlF83JRO/smojGN9Hp8XjDdlT7UOE1rPNldc
L6+c1THRzp3I4CkkEuXV+7FDwdbxxMuevUorqcR5i9KmTQzfr0WEdY5SDnxN
JGMYUxn/V/8OmiSWx/FNehOYz0xmCCkIS4Ti2IhUBLfSxMa5jV3NBXeWMi4A
HooHgLV2wi1sm3EYsYa/q+U0uUts2tL/yjgKL0XevC41NdlRcVHgXXvIO1T4
w+3ZyPdTv7im8r/o233CjnU00wypvcX9KU2Ni+Ts/a2RoFCyww0uFKBGUbz4
fyGW4jZ5ooeAIDA1WKbDAc6ji4XAq+CGR92IpL0uj1e1cI8za04n2qoSllaG
MV+j18tJ0kttdgyMX0AKdf8uvsrP0TM22cBcMlII35pdyjwHiQBda620z9EF
OSIJatnHa1qca6omTan0LAicmmwuoYwyEq9MDeJ3zFqgpMNusQ0J9S715Ctw
rOXqUbgoySO3m9rMbne/xk15dQaL0j7zTzbJSfyhizHqGhohBt2YYItbmINK
F1QMrOf/0N/gWlPalgxJSVnn8s7eqPb3H+DOEMkYKXB4UPYu6MNXqszrJ+8d
eD2FMIhkyPvlDX7pcHukJ0kmkOa9Ut9HtYqXShSTubCDKzPfSHw1N1DnaPLb
6H936CamgwxE9xC+qk4VIITR2sAHO0pNxj68r5/9/q8dYMKIOv5zqNmw/hpk
tbHKBrDHV52yJBUqkAoKLyoJMih3zToB3GFo/CuYcseBOXeHQW+QxnRABH8z
smZ4bg0gQRekuAzxM69qzBcJD/X6YW5nVOg/sOJm0UzHBgOeik1qgDBPdFXu
Ol9/YvHCgJYaoPfkPFRZirOItVbwKOSdCCJAqXBAIbGhI4xE/H3zID43xh3L
jYWCPmB/rnLzMY6Jkv7sGszfRYhvqpfm+UGZ4yx0sKpIh33UtsGmVedyVnnu
6pzBNPQwpUkXidLIcMmSac4IM2bkZqEyzsGRyFo58eKg92Y1fWSU5UB/kHcG
JAsTbPKEzXKojCFQRQQrw90OJHB26a0QhKfX/BWKu4Ynz0naW3Hh0SflvSy3
GtlPt8R2A9d7zP57j4SpFl+BvtzXC9tIn2EQDv9D608oR/cA9dQsTYNNRP8+
5m6Ogss9k6dUXMF0tBa/WFkYQ+GQOSiyz7Y7khWWg0obCeL4G7fSwm4Uadda
iQLcGtQboSYcHMlBfAgjpdp8u436uHb0Yha20SWOI1n2Z31wWU3nqvuzvMb5
eG0TKrCZjR7j41fkwuPlrXYM33aPO1DBCqABZZsFoxxbWfHET0tK/dkWLFay
11Ughm8anIhBsaEWl8gPGCS//X+VSCL/2pKR35CvZWDHqWv3ncFKZGbo2XnW
07HehkAkVn+YCk9ONDaZ1LDL4TmfvuBhzR58nKaDKI4QW2zfvTqHdYBobQ9+
et4bzXjOltvlx9svVT6RdMTrg7b7yjqql4BzwG4A6mLtEtEl+Mt4fBPrc87z
LQTpFjSXHVPZ/nKTGOTgvFCIBcCjDH/gAfb5FyZC215qICSPOKio91LH1wN8
X0FcEyQAlQ3pACCB+lxROAAe7GVPswzziUFT0MfpYFMFzzDTr67xXPo+nzh6
3SePkRTmtQGsUp/9AHb7m0UDtjjpdKlRa1DhSfOrxy+PvO6gXaFZRpmr3WdS
MsfG6ptoPJPzwXWaLTs/AarOWy4ICe2Lm1aqguFmxBVUBiTA8HRhuOfMZc8F
iU1VRMljL7NNGwSTzs8GZbJMJW7OKkyrRD2fTU1w0OYiUeOU7vIlhi4x0dnA
qsGkJKcDsZeqwCcD6t2+7xOXCO49hazBZhq3BhfhTcu1x7nJhCGkYMsVrN64
czP30S89FtquWomQfgdqaT5zEZ+hjQhqyRh7mQ9Q2KJVQBFdjPVS5nzF2znu
pB1wH0mquWJk0/12jX+iEx4VwyuamXlf6a1LfPtblqQZTht6MU8ThM87lx5a
KdRXdn/w74EgAdlcaZ9HdpmChyZOqYS4Xd3U9CwAYM/295bJRrh/QcMdu8+0
Hgh7fDr8/mP1l+8rk9v9ku0GzIOoCHSH8f/XymEcz15MzCXOEnJX/D7qDgGI
TP5IPHe0cOeAj6qBiTvjZRwIBT7M9klCUyGIFA+YYKroi+IHSCZCizoySzdx
dF381hFRt/qQLnknPRL/gXAeHZiq7BLqhOED0eaRW1gCVITFmnwUaxzCSTdu
j9FMm4965DXIKvYYE1jZfzG70BV2MGpFEsbHe8iJzpcyEPdJPu2tvAkTh8Dq
qqHqPCx3mBU4dKzp2gHkoo2VQ2K+UJUYkwOIe4Ptmnv4gOzmGjdUvqGAnOOe
93r3eOwQSV2fry4zmUyYvTX8oeFRjInAW2V39/CwF/5lZJut8nwG/mVdSsuE
A0aO/v7gHRo00blXzahlubMcNJl9KJEFcaVx81yuWdWvCwK7cJyyyr+qWp9X
HcXr4izWT+e19QnhrKaHdAmdiFQP/dZIJMSLUxyJ0xlmuJFaq4nTxPcTGLpC
Ws2mZ6YJdXIAtdZJyqphi+vGyRHd4Exjlzl8YN5cAYSeFeCxnKwtOkRf8Knu
SDtYCP6mhejv2dc7cg/65AVUk6n/dIgywAaZQx7xcN8RWP9Tbbx8iFf8wdo8
i0HdjukdAU5JppCp//qnlv2DqMRZoKW7gI0qWEjoWYciKmvv7jJeeh7FbzBq
RJN6VrrRRQhDpiHuxWf7zRhmuUp/EoJRs3DV4ixpwdsR+5wu5xYp+88MbZdV
J3KUzE0EA99QNosKYsz3F+oM9mmE31qV7aIOy/fhTlzAQoJAN8ivBKOjX1at
Y3ZCp/4C1FrJfnsQTZzUcecdnH8aHBqeWjJ+keTxBtt9jpHUNLceko+CPuMP
ySV6kUWuKjMtOCPJunZXzMCN7FyiNRd9xlu/vr+LwDK4dEK5IcXFThrxuav/
pQNZufwNI2s+CFXdQuHm8ECtVBVKsFDflPCZKKkjPEHgJ8XZmQrN56QKTUhG
gGyj5c3B5k0ndeB9O7M01dW/MQvN9lvcdDgyLbHDVf6DAVUE5dcUI1iqV3Fh
idL2cIHaDy0x7WDk5XDHHEPkLCTxx+JlD1FtQwiyiM7Da0C5lSSZ7ZgGx4T+
8z/oOogWQlaVf/bU07Ev4tDTjr1NFP1e/JXJC93d+nGyhUb4gaH47Ax23ZC/
/o56SK47hGpsvx4JhV1XluB93CVlxdLLNwkdWtO4ydi3e1bvuwrZoHIavAcP
p7XuwyhhJdXNG30bh68VvnI1Lg9SSueUWueZYqMsj+hFcGuQJlkVFZnivex/
bphBboSR59R0nQ08MzLlnf+/iF0aYwYlbKE2nvn5HXn4lnrd/xDFQn1kXh5U
dKCkSchZB/mvzmCNfK+95m2JztDsJWRP17NYs+Zf66TU3IDcNaBFBEDei8Zu
NcsVw7z+6Y8NmQuxFIWU1yTBUjNLyMNe77yHrO+8iYC6nkLLn/EHYtYQIeAt
uHVulNSPNxF/os6JAqSbKUvlQa7nlPp0BjJrz5nMN0WYrQ3MA9Hl9up7psHZ
Txu834nYZ9CA+PeXEOl0yeCpc5X9epjCz1LKJyDSh4nA5v3u4fZ9Ie0GlDw8
yOCAIVpUy/FsXaOgULViqSFNUFd0go3E5rfily1cdoZXApPD1RbSE5TMiwVX
23Bjj5fLlJnbxb4Qhdvruq/dhgV0SLczaU9Xx3uDAdtbDB9ulpY39lOc/mta
ckRBOu0hz7h2ZfQaHc0pL4XVx4O+LnktSb+KLrnY+7n2dXr8mwtG/wbgsEzW
TTo7R9BhGAlYQ7Iugis6pDe3bTZK3WkS/uYdKUsZuL2WEUx7mqsHPwY9bnF8
ZtXjnbB5KFxB9JSGJVR9xRLCdjSpCDoY86KG04gwbtlZt3eWf/f+pKENXE0B
g1MQrd8REfXgHeRq22opJaEANyCYXWgAPzk7fB3V6C0MXkkMfj0tlFEpTiAy
xr5lUZraYiSMRA7Evd3aNwRL7ADFpe1o2mseHNYO/Il4filygOevdA6FqY6t
ggmL/BeJD3DxrbnXPqyGU4CpERaywtvZj+filxFxCMFbr9HlYTlZ/LqtC27s
+t1vpdjPYNcwo7d4jJ/MxA0nweaubXMcdHXqfVaRMAjoMLGjxHgjdEky2FZv
WCOtjhN7Z7bv/KTw9J46n7nHdFsXYVCR4DF3eMr+DTNGKiKHw//fEBqXAIE5
WKSXYu+QYfZHPAblUS/NmyXjAjzx8r6xtlLnRgixhKY65bfTHmfiAYi/t/U5
pGBPTKB50BISNfTUbEaKLyGQwosDrQ2qAvJ0uDJqTHmKQo8D7cjpzGO/lXL/
PRtBhQOLgYCLIkF73gabX2GE7fE8Au/6Utqu6Cq5uQVmKLW0WPSyjnmrifyj
lZTz7oqQvRLPo/jO3Gi7J+WU+k5Bc3VEsztcVyW7/pt7F1f+WPTKINqVUvv4
krDNk4jKgX6gCaGYxbUBQ6+1NjpldH3ijJPBAm1QtrfWiYYAw/dmDE4SbJur
TDthaX3eHyZABzkg3DAmEGkQqbxnu26HYAdSPOTPkJqvy1Jjq4EY7IUgYN3s
rBNCIJSlYvyhfRD+KTFpVqMAbfjW9OoUikyMxughkZ42JsIMo2Atl0doxKAT
hIy08G26CT9Rv7OGzjygpN/yRXNiRcT5xi1p/662oXiRu7STlGhHib5AlLQv
AoKZtcOlSKrXsRkkxTUJvrEkm6ms/u5mmBtCsZv5QGqyhJWO0UrApanQdnk4
fFWdxSz9HBd6mPDOElrdDI7wAiOilT2HtJvS97uVA9+BxTNJi89P6ARYI+MV
uWEGOhgVx6iidlDgMJ5eAEjzK5ULlBqWekt/ovbQXLwdpYPdpYx78eaiuLf3
JJ+8fmavnLaBKeL3vZwdpoflqeMmVKgIzcRgOev2mYWp4XSlj6ArWZnPtZrM
HP2a03OWahfxv96nMtQ7B+My7fBc1lXviwzACw9XZH6rp+LZ6MhaY/e86eut
YSJNVqPc8APLjmkQgKKtpAo1vBXNkoA7TqTAdzZtEjZNzwgCHCLN9zVH+ZR6
eqhRO5ogtsPORaekBBZqxECF2fjhL3mqcuC/Lx9nWnaolaHVcGy2iFaQwljH
iVhdomOsbK+AZ+s87YXoDm5cMtHar9EmkfSf15aTYkQ3z8j9EkhP0M7xMy+6
Y9lHBW5V0j6E1knWUHMKaonoV7sHod9JdxI36Vh59Le8O6/ugZof42Icj6JG
am/8hUT3lwkkOgsVKgfRIEy6npQkOSEM+2wIaDfM+gqfAe7CHyArO49G5zYf
RIsgV1eCd6Fhmv46RChdGZrMmUJE+AJd0CV8cQU94OYxizlEYRw843R7zT1K
rRdLsd29Beg9Mak/Wm8Arh3lgv5RsE7fdnMM4Pt0KpoHYxqRd2lL2+AL4ofc
5LwCvPH8j5eqV4EXSe/hanhePr6c0mIl2Wnm+6sd/DlUsP9aixG0ghkFuth3
4ABgYN16nfRDWJD0u1iDplQyj4czpbrzCFB81RFy4GkXDtYA2Rr5B41tfvo0
Vmypl5671Ig6vNPLi15EX8g3gNJzH3EXWS5Wj8T/NlZSVYEua4P+ENX9tBS1
NcwmBEM6kggY7on1PQNtCAR+twy9VsyyqW0iR7BXatwo7wXIgRcaC+tDqxia
JIOWxaRQSbB5IgPM7+99zk45smuk0Qp0zygb3l9hjrx3ADjWbor/rGlWpXp3
ldxbPyvPZCACORQXfwa6x2D21rfLDkV5sccpYzn+4z9ido44kw9iBw43VZd8
DuzBMAfgW3NTJ2Y9NQPvOKuvi8KM44mkN81U3LBkY+dqq0I04qt/861p1rRt
MAVIeiOX4XVrixwer9Kow9Ju74khb1ITU6C/tyM4xoZQNGchyFqBii5ZPGPb
InnDmNwey0oyxVAI5lccJoLYlwoY+nJHwYzRThtFb9Jr6/ESI1cEJFOo5mxO
Bwr87KxujlNWwxVzgQDtCcdHdZXUjYBC5BBYHBChgznSG/L/ya2a28+AY9BT
i0aBXsgfAa6AgIgMajZ9L/5m6xFRgrcvtjwBQlTBabPILOjO2rVAFypGA5US
KCcMxcXCGOkFmKNJwydjqUl4F8nKofUhtSVW7fpbCMX8bqtgpwirCz4R7lut
2PEXDs4PZrvzniiiB2Mv6QuPP+SX+RwJ1I6fAMhS+xl87OrgAfY66Hj8ctMn
G2TzH7patqXJGID7Ev3laeT+ouPAUJXZ2HMW/SsMiPRJYh036wnKneZppz80
CSxOri2lccT52F7LBGgGrTuESbl1Fuprz51EILUlHppdGSNyOHzN1pCMc9l7
JreLCzRLige+PovmNJn96ZH6VXODUnjPY0/07XuG9jxfBgPaIuWqPqyBh7dy
AL6TjS3/wWxLK7wqbWrpI/wqYnMEhguc/WmG2SJLIOiTB8gkV/FVGQLUyz4Y
EiqJzs0jNqJKURnCRUxALa3CJTVNwt977OUlKjvpC71eya1KSD+GONbuQpix
voPeG5y1TGud3YIIXxW7sBE9QweX5fM/3i/9yWK3BklRwoJXXzsLilyErmqM
4x1xCJ39e+F78DudpWqgZPZp9cnUVBvJywBNV2ofdnJH1rqAtrrAqUcKMa7D
FqZI9Hua03O518IQ05eH0wfdjKURB8vSY7u7mS03u5xJCrgWMqcXJooZ49aO
M1vczp6kA2fu5Tw5bCf84Jmbh/aJsnWg7XmWGQ0JMJWmfcd9nKGhw9YgGHPQ
glZqRhP5SDhnFAa4LheUGhcXf6vpmMbmfLrX5+r5LFwCXgJt9HvNzWS4BJCG
PrJo8ZHdHGwbhs8TeBDdGCsdE7OKpQM9BAUVGK3Z7jNK8S7bcIwB8uKsINFH
b3XZbGvvsClFugeNUgVlfajemAQJKT/+UFCCBDAYSBGVb3SZMj7PA+rGIKpG
idqCyL2Bhzx6DSBV5Hg39yPwE6WfAH+vMtjMtlu4xQe/eVmfekluTHBRY8/E
pb1VXIgJHmRfFc0YzYk1R2F6gKUhKiO8U4s1Qi2MlHviA9QUfW0++NY21bLN
qSBkxa6qg6xpL9CU0XbWrXMNuLxhzj7JS9FL59jFc1vGlA3Prz7JVlDqc3vh
5iOZkOmM0Ec7hw0bI4VbZn9YGl/jOEQG2xAmJID6GHtw3HvCfwf8bPGbl7Dc
oWkODUMLtLIVpyLy749Ryez7VQlJ7WZNcC9R87b4UVUwsvGxNtzFbjyij+9C
89X+sllWxZxNP7Nkz/DtOXZHYZmLHGOudKKzrUt+W0RB5v2KQKHLYD0rIDwN
yY5ej/BnaYguRNr6/4C3ap3Bq9wx6WHymaYCp0xh9xdoNxSd3gGKzaj+FxAj
kjBkcW7ji5S/oRFhNl8sw2xyFt7X5UL6cG++ZzJ/4vOlWcGKjoHNLDgWC5qU
OeyBd+GfFMJ8NbabL/R8qGgMfIQgg0hRjZBHWU6Nk3vO0mdfrUESITdZ0apb
iMt32FBDC1XnzLeJlqpo1HJB13MJA4pmuWSYhtWTXqU10dO9k77JUvF1/87W
jRzJRr7hhTi18mmhIik4VrSb4ek85+lX1qftFC3LvxH/4uFjAm236xSiDHox
7CfPig5MOj0Kg8eoqrLg+9RSlgm3oX4ILOSdaxDaf8yP7egXURBmAUwfIlks
NBsYGHpxy2Q543XjYRxDyJfvO5251gnnz+oPSyQhBXnXxY3p33zbyylRufln
k9GntvrXg880r576xUiQm013r+l5yX3BBK5NkRkfA4lYKa1nBOm3cQEUXcID
X+3N1pUWxgGIgcj0wgt4c6tU5zfi7wHK974N94TznUBu5UKQs7DoXPGk3M56
KtKMAqToNwfe+34lHG26fvpziuTTTofY4LulbjVknzAPIug00IbosNaHSk4S
BRrAQOPBwMJRD18v5W75XeSpfR8cVwn3yGa+WG2gddQTF5DLt99TRUTusxDU
sMI2nBY0+jJfBgB0ZbUJtUan7rn49aVWwqjcv8QetVRaRSFZfK/jEWyDtt9Y
gb7IBEyb6cftGlqpgX809a0I8wPKoZlTYpkVJZHDaTi6RqKfaPpbscdZncNg
9hMLz4VFkboVhoR5tOXpFBvXrKx2nmzXFUYCIe5yUW2ogl99uZyZE2/CoLu9
Y18BVLJ50TFX+Pkr+68KGT9iOc2P4My42ZRyZOV7Q12qAow2M1SX/ROg3QoF
GvYzkW8HqK/xTaHHoW0xH+GT6ZEa5PB7nEHMDZ3jGd/2CvASpUAd5SsJgweu
opaqrhqlfi2gvCXwgzkNjoIoKnj8jLB0PFRi7DKa3rEGAPykd2QwcCuL5vTe
6ZX+yUA5xVzT4HLRjaEEK3H3H7rz7wZ+xW4UuZJmKB73689YMWH9BVUIpdgU
SaRwtwGcST6X6ilYG7HmhJunkdiH1wpWKKbjLbDEt28oRCohJB0LjPyrqWEu
FjJqzPJvnGRbGVfI785h5xjTRacsNGndrvDXdondgbTrV5tE/EMKrQ1HIBxF
0vMVTWC33Udn/93Jg2bMIpvfJRiFkgKaueG2cvuyP5dzyME14e4Asdvu6n/E
Xgxd3l4BGzSlYOi2v9VMgwaC2pgfhnPZFc6hh5vd1d65ntKNQdkysZlPySnQ
q3QYEf5xTR1Bu4K4/vdeSvpq4ppk9jYznDCQE7nWrm/GNEPelliInhjDtITQ
ISeNOUa+bQgJ/u0s2x1u4CutcykzxYJFPBWMwUeZeCNDCyYMAaGu7/sT3cBW
b8qnk0Z/ItsIVmE7RuhZJs2xhSbohGHWdfooYm9JC2UeBoE309pYcRLLy7FP
DdCVBe6k/94jaKMb3epqRnoGkZwQ36exBGOXBqdcona9Y+UZuTrTwlkD/tSl
XUchzl+hxnHBuOMmTqt13mcBNgElMuSkr474v/b+OMXhfd8AvD7JRvNsgNGL
oUeV/HehBrklKWZLg/1TnBvrrOrVjDLYBCD5IxQ+qHycMz1ClcXe+G3kCTzt
O2gcGFvkrl2g8fRSFdqERvbsCZwlYxnkkmcPcOq0DS9ex18wmQ9ZHdaAJrAw
nJ3IFakPTnRV8yZHwduu/8LmdopbtyCW7A03LsJCqJKmb7G0zC2dkjx8evkY
2dLnCDiPNOEdv6E8ZqwPSsNR5DAJ31FMGipf/BK/zCncLag/QHmoYYLOkgWu
4h1M/NUYksrP4SkuifGAwr7UqizHVSKcqZ/EWj/r3d9IYoCjcWyqcB7RyjbN
rDLG/qDKfVKxQIR9x5J+pqN42z8Gg33oBAwkaHp4M7EDoFttVfVp3nFMmT2w
e46TpAj1LW/4ZVTAtCKzWNe1jPjZBiXvR1iY8oSU/+a9XVRi8H2fLmZWuqR5
rgT/JogqegZWAu735CSfNoQhau2jVOpw5SbbboawGooiwEy79/NMfZkOKxSQ
zvDHyrlFxa/NUk73MLuggRrpr8hffD5FgRJQ6RAXnlALYdtLLwPLX4jblKvU
XVRVyatuWjJqKsP/nsCf8l2Ed+6itwmfbEECrP8B+pLi38aKNuFXWFvwR2G3
ujLjfD15vqASCOrJ4sYbPmNntpaFd0pmk/XnSjpWBHKgW8kMauxXEfMb4D7r
0xfwChqrcPxhCVXGzYXx611xQ51I4ZcfzLpCtPy0m8Elo+XILJBbKzQseMUA
gjHYsXL3h0hJKEkbsJIQM+Yp2MCWbmN0BzDKRQwFL05sH+/yGKOPENkL4uBA
tCuXiEB7Dh8fKGAZMrWywwwZLCZXR1QL0I9ihgb4K275gFXXKhxD3qI5tZlD
uXzfcuAFYcxcC9Uu8v27j8DN8YbuRrrK0GobpmYN9iUy1YOUC5vxojqf/RKb
qnKOfsR3+J3m7WjkzCwcnBxQOdZYpPCtZohyvvFhNBV3Tw6BMuXBH961f42+
KtIE6z7fKKgDeDXxesY2EJo7kMAws4EVLGXjcCJM+paNp0Rg+gVQlW997UEk
phAVAx+Cqg3alb61EML/So/lArvkfaRoCSyAJNLIt8ExNZ3Vp876ZmC/5mnJ
bzUVnLnY0kdZO9EimNhNmtsp5yLGXYQCBjg2K6NaEZwmLLyiVcq73V57QKKp
Or8VhCfMQNYUBgx7H97ElEct+0RSO4qPTA6A2B1Iz+kST1uRZVuqa4bC8DKA
+ujoa9Wct7/25eqrcA/D+Doj5KbZuoWVv7zK91tMNbkzb1E6GxLnePlVzoNh
WxGOnSiZYP5g285T0jwfZa9uliFm79alKEX9AluOQfk9PLfNoG6Yr1QGBKWZ
DiZCH8p0QWWJRINPtSWbyLWAm/mLP+TC9Ilckv2plwFI9YuyesUajXdb5rnF
ZUQb/dWq2xw2KNyKFGCPIyZEhaAygawXSxjMLAdYc15gjPqxrNDDtq+WyU39
AELm6dnfr2XILuny28kUXcj/w72Es8XrcZ4X1JOxs8Pxm4duACsMgPgmlSuA
xqAY/Wa9lF2FyXIl6hIKwqkXGvXAhCFoMp/RW40ig4ixwzamu1j3EFNQWY8t
SZEM68h5yCf/5JQap3XZZVmwYw7Eic+qHIJJyaPMAE2al6YWbGgsOu0/bxfF
RhyG25jg/+59h0npH7fy7A0OO4yPPhlsRzaHyBtE5YbMPvjMtRC9l7kRP/5a
vhG/7mjLKkQzWe2JDagb/VAnI479J9r8FO+aLhqwPJDGFlEZKErWcnEHXkQC
GSol7nmtsdfcS17efo5m2DYTvPQecl5XQtoXfXfUkzI51V2NMrxD6SC5uQIT
Vr4fvzH6TcyIm7Kf05JvYJebO7ufIJ/e9RJRC/revuHy1s9DDfIluZ+slY+g
F074Kn7uLxWKPXLKbXJC7Ly11dlKKHuj5CiZKnnqvIbNHChCMdyc5fMfyuVs
X1j9qEx24NcP+U8RrMfhoko21HksluR31wpUThI2n7ghdxXrMJJYMN4YG041
L0pKaoKS9pdSOXS5zpIAjXaD5zjyKB3QnrmrfkNocPpaVnGhy6aqgbMtK1Cz
qMx9+pvpLPpDhOmOJ4E1LhtsPUl31Ov3h3vBLija8vgb4OVGWOYO8RTHyfo/
0q4eSaz7U0blPrN7VDCGsjv1Iq1jhgwj7E9IVI20T0sj1xZ/n/52FC1Tn/cM
GT4WeywVqG6vSP2AYITo4BwyF0TGkRUeB5p4brObE8CkVCT8+oy8anTyTaDR
bpl4Q4igBfumVoeQCEpsI3JrFp4fKb2eyRqwIHnkenMtoitGm2tBfAB182MG
5g3hHOPP5BVlMLXOiHyyD3HdolgzqYD2w750psa5w9d5N6XSB4r20EJvswkQ
rJx1xPSVhwumok4ahoOoNFrz464340BKl034lME+kyFUSWKSHiJHu+I2shyB
4u7u9g2bQvEn3qXEMcd4btRKj3YLn/PEJnnCOGN+fGvD4Af7TGSd/5ZUZKjd
1lmCY3vjl2pR5EI1nxsHj5O2pwF0F2zCvoU8ixkbd2p+LeromGGWBopxllin
ZcwNTmtKBD0Q5tgIc0dfnK/2Yi8LE8sb9GWkzaLOgQ8Ij5HjaZ2ObwggOvb+
iygT2Ni9YEhwUUVsXF3yl3J7pSg7/ZFHUFGwh8I+4ezfoUZlzsF+Yyv17rRr
M55k36+OvSdcDrqL/pNqYIT9ni+UMh18ffOKc6eNDSwU1pL797mrGrLjs90P
Jby4Qy363X25iRgXW7V4pG5t89bDTylJzUbD8HNNPAHzeFtBe+DDQvott8XR
hcPyalt2TnDHKD+9yCP4x11PLKvgibeO1QaJoSml51zJA5QmfZsXiXhYqrLr
hZk+5p+81yGIJd0BwsitIKAJI6gzQNppyYVETxgoCGN1zsyl+XEdOz6zeWpz
WeVQByo2jELBZS0zAJENRCqQ2HELQN2iAlTmoOZVRWBxdpUQ7jJCqFmhC4Ag
/DALMqnsbr5pkolGacRJLQIQP2+YC5w2/fOCdCxsgenEe6qBeeZl6eVCr/Ku
TOcuEh7eDvPgi2NKDgQrodFQi992+MctP9dSafQw0J8gZGnJZCRQw1FYv+Ga
mvf/8yLhyzig5NeV/dWWTR6JrobSbXP9TdMxnOqLVDOST9Sns8Lxw7iZyJnW
L/Z0vTgEMPxU5wPt7EGZFvUJUAQdxxkRlLDB+SB2VjjN+Om0a2r6uXK7CeKR
ZuV35VQXdtjgIxfjAuTp56Z9pEuyfbtAGYTe+PwsrGkBrXw0MeROOpJfdaeM
PxlGG1OdpVFZy6v6RUdo1fMcyiNKzRmpVK/DqcvztNVUuGLzfFjlMA39NrYh
4HNfKXoQwv7ChGjbEWhfiu5PYu3+VVuXIQne1z4WlY6khJl7qNjcyrBC/NN+
4yOWowy2D5OU7ynpLqkNijAc04orYl+5scKz7N7gyACq/Q6iBnXbYpGXoZGW
XfjwuXoPwYkxM+dVhXECb/+kYEUVqNkBNTv9EfA1wVMzA6Ugo+2YbDO1tx5y
YX74KGfxxtKicqCOdcGbPtLjkU6iQCSrBfXbXbCMRPCm1EYSQHsHM2SukiRY
/+2VSv2NSdnnEZtC5xjLsIOium+Hd+X3bbJKt1gMDfxWbTt9nH6U2ubYZxlP
1n0gYNKz09dOV18UiNP8IZUK9OXpLLczcandW3F6jZlLIGTp4ddEXyDLkI4V
yCQZUuoU7vLZyGoO4LjqpwzjFr6KsCfo73GNUtPlcA0qy0AUB5jzmAMKddP6
FaIyNylp4kq9QcglhaQfoE3gnOsolhCSvEb+TyC60faqTnxEtfSJqTOGWODq
9hi0xT0sNPb2rtvwvvcr3QMKik4h17oJj9Xx/24ldFR04JExpOcrpdzD/RCa
PSPzBNVyv/MLWzHnVf5Zr9hqKUwyAhImGfeazhhlt/JWn00vd0O4qnjEoGrS
sRntncow1U2Og+ejglXAgGYGCxZrPU/fcSO2Zf+AVcfSxxXJA95oNuTf9RDK
2YKcRKlo5+PX5XHR2ry3EJ2I4etIEwO44F/HhiqxfNmLNAnGNrVoiyhV0PDn
yrPG4GZ3TN1mSAi6ziJaJNCCLeyGplwuYSCfrbZSlbSxLzDZfZ8R0Pb2Bz94
JoT2gCcAXOWedxMY3Pwq6DsGqa74WsALAdn85FGdqvRGlPz/+vS7X8U/FwRi
OCqkM4fGb0uSqwi8d7jXbdbmBLCZ2OW18WX2R9P7kINF00j3UV+oAe17L6I4
aWua4NQ8fTwuRXoSP+CcBHvjH2ErJEYYzHH2vldlTkZDIm4WSwFnROxAv/Ag
t8FfkCc8Ruufa94SKGHGXdlLMOmH98+nfM3tb5FZHinkYLXq7G21s58YHqq7
W9nnqr7AgG33FqIronkgkt6KmgLj1Mv0Fh250hhSo+Cu3T7bZfBnMDYpIAgc
VjZ1E+syJZ90PX0E2AHUFgCtl8VtVX1d+qSksV93ky1UyskcwAWkUkpT/Ptu
Mm6+Fywdba3dTqmww1rtZk1rUIbbwBdDcJ81qSqZSuFjrJFDXXHldOvCMr1R
iB4LxffJCYtMmnpTcCv6/FiwCfXXaUCNd5ZxaAUGHk4hxSPCh7PCE0JanaxD
pBcheHbyXKWWXxdQ4d0FqMSwYO5JGMm9RYzQ1j+Xc9HwvoTPdAJTd6fyjeUW
3837rDkAcLt/XBQ7iqttdN+lMRMVB7ydS8mcQpl7pqMIXLVrfRc94Nb1wryK
RlCvgoUKi/8izBi8RUdEwKbnWvXSNMxwP3KFAhxSIcrrzNt/lwsCMfIC9KpM
QoaC9NY4hPOmucdH4vsv/a6aFpp0PhB890MvYtlSybpl2oQi4k/XGxBQYg8n
Wb+nT1jZvF4AZEywlx9wG8VajG2bzNSDc5H45laTwcHQgf6n6ly5RpaTC9uz
R7g2XsWKfnoRHQc/Keh7JNwdDtNq/BTFbuEUqN43tcaW8oRE1NT+8Xb4lTAF
S3Fryk7OtB01E6hbeqDC4FLZIwGNmVV4scjayVw5HuQhTdnmsaJ1I6mMOSe0
b0/7mH9C8ONoJ0yYQEl/BqQh6Rmvh2oJN27p8U6Ksc2RfDCrEEUJxQDa2oXy
T1nZ4a1PcSiriWHBOPfrlqGokrnIqjoczFWTR13LmUD5blZeTQJ+JtIlHZj/
n8eaDuyZnX6tipXnwUvlD1ZLPhxfpdgAnhEBzcPakx/nWSntslhMEF1vWWHD
VoQhj5Gb871TqBCwb+pjMM+jA6lu9+pTo1ylZyIBVfzwAi4+iB0h5N45v46T
SqWjcODV3WAxm7mTpb3Q+O5rnOCV0QiejwTqfPKUdccQl1dTKUKc7RKtYfv9
b4yACQgP+x39MENkK1mWBjFu/cZDnHl54SHZUjHAMJq2EEmbRioplh4KAT2k
XTMVtwsSSwjZkENeexuvqBTFVDsVwCfNhwYJ50M14Vl4EAxSfN/ZLIT9XA+g
RkG72aFjFVPVRsRM1gVo1s0aFaxTTkf3+G5WRxgljFx25jPcKfz8w4M2g4SG
JuPqAkAe2ZbbGSOlx4vMTil3eWDc44U7qiIEN65/6p4zSLJmm5kwtE38qQjy
1DHo7BX3KXiS69lNqsLDMulr5V16rqrpHBwvHbHzs09zshv60uO4uik7aQe7
dM2QN7vRDMc0GNS35w9RCXh74uZm5Zesx6FsPcMlzC7TTHd0++XXd4lvxoLp
Lus3QcxEEZLXwXpeRHrs0AFYOLtuetqLUoF/J0WJ5L4Kb5gGEX+rHkCtNep1
CI8LjARzw8i+toJBwehUHmlhZtaXrRPOzmE8eH6hpIqU07WLp/m2A9Pjkb5F
xeU20+XHG/oigGYNtlhPqsv/1U/AMgpq798cR00JsbmKF++Sgt7GWNAySI63
YOV9dMNkiFcfwPjPJW/YSPxe4+0hZ7hQzoJ7OVSKXjr7vkA06Xpw7RGEGSbe
jTWeC060xrkIdb8h7UksoGTB2qqT08WjO8AlFBguDxBv5J+kU8xDUJpZme1A
aqZ7VH1tRcmOPjyD8TnMj8Z6vFhmupzEBAUDmiKQTYFXE0Y2mX6Y2nQRdGTR
YTP9Nu3sbCoWMVCSHzAxe4vqdQ56kLbCZuQ3UEDEb+FvGa80xC1Y+Zl1iPlU
p7gBOrUACqt+Zo6zdPVAk9c5AyjkuRW7xoeRbBK8b6vVzv1qeHb0zpE5gohx
E9wVkF9fdVszcMjYmKWly4rSjQKA/RGiuJFfzNteD+pg3ZgxArSDZPr2QOFL
k3/2lOu8jeyl1vE1BlA31HvisY91zFsn0Du4Dg8KJZmk8ByORDkVyx8UVYGy
QDLl/3B/F5ax8MhTVN/XQbkpKKWaVloj9btL0j/C5epNakI/mcEYNRvktjzA
KO+P+qMBa9wSiDX+HNS9ELu+WuvC97wDY0a8jepIay97HKPhmF0bgyJtQ2A6
t08ZrWauE9LYFOCAObnhM1o8j6UuycswzRwJz4ZWcelFrE2LoDbNUluloYfT
vxkpz9PjW3ICow0n4cPCScqlwXlCghgctCF5QRIuTGX/vKUCb4qggq5MWcRW
MEAL6yPtRWK8ULanzyE1Lkqkk0rACxBw12FiajlbdFWAIYB2mOkY/ap05S2d
w3KFHIxPsrZrczNXOaBLWmBMO6+RRmRAHqs5udl0xuvbvrQEsWAGJ22zAgEr
7lJxtSiYBW9gtaJjMu2WXMwINW0nAFXRqAs5rsZDB92jbP0cBwqF8vU9KDf+
96xYAftkkOWsZaIiBMxi/kLk7c0ONCevzsLQkw0pGDWKGV2YCCnqGRhR41wR
4mbw92fj783hbp78CilQyW1RWwHqrCMDCWmiGDKlxM7Z6vHErGQetrTNPSin
YMgVdh6mBo22KvJj3Afat8V5B8l9bRXZG+fxygcHGBwymvJcL9x1RP8RDM5+
QBIKB7iY1F+f0o1urYesd/nzJJt+CZo0hXFuokfHjv6Aq8q1ROiVHOlBUF8C
nrR8uF+OjhlWLJPktho+0Ca31OzjV6nUnI53qiZE7FJRlos/COelrM0xGYqn
eapoU7jeDXyYyj4KA6FaGUWja+S4ZSk/kEtmv9TE2C1BGICHUD0qLdf8Wji8
OwgvLUbPf0Ku8OuXc6FjUN0wOH15oQ8Jow9BFEVVe5du7d/tjR4Y4xPrjgSb
Jk3VRuCrzJZbYqaBt3xPzTrlxrZj3rB5nMrP85xGhdOXF4NPLZ4Bi03QyjVS
WlYKGP3WQ5XD2alcZzau5NqNMP/Yoi0QIajAPecI+2F95zZ4ZNs6I2k15SLi
QpzgEt2jARWfWmRPOk63tiu5GDmRpExwAJGGSiqUD7XUZoRnUoBCgwR1oFUa
iDs2SR90eG8C5OFxLFRDeI6tBrH8a23x6J1JSqzr4MpTRDAW23y29syeBSBw
AyiAThDfQTuJaeexTB0jzChdEytnyW7T1ZmcSvKl+y1CBAAt6393laXBkxnC
RersM2pAymfo9A+KWamcYDshdVishdDW1zyVLApI9GqrE7oJmeRvBCEKPSEK
MWAe5jOMM3cG+0TRSbI3gljQX8DMTyVUsVG+xyn2J3HtV2yng60rMt2tXIOw
oP0vIInxWE5gX5/vTLmESzEibimO0/6E27Y0rsZFZyr8iVCzFkkvCWF9Ot8u
9AtNximTCD4ZCDvbe28GQ35CJC+1dP1IQuhfJQzjCbXnOH1ITy1wVrUvbgBL
m2SfD5oyI3rIWae3BUyA2TJey0VtrtB9tZ2H+wYHUW3GgsP/IwHJz/mp1Owx
FqR8LqY3Gsqj0rQy/Lxa61+TyO0b6eZPbsuLdTiAS/2P12nVr7nCsfPnc+dI
hKjRJn2W7vRfglV8v64ZhJeuhTuwxd3IBRuFCOiUR0qwY7eD4c8w3dJfaAUn
C/UUvur09ygh0gC8qy0OSkHVWbA+p0MbbkOxDubDuOBTFPciVT8X48pg2g7F
LU9xK8ne5EzJ1FTSvPhn6ONZuwve62YvC0qIDeMLBzcpdDVUU9cyz+ZHHaI0
LsLJrlccKrf+hx43DY2ezZCcYK01LSUSdRrg3NjMCuO3pAiv/u5N5tcMlLla
bwJI/FQN346j6kyByVoQIyUcBPS0ExevWZ4Kbpm9DSlNRCUsWLH3kri03G3G
cWrchUbE0PxJTTtMEcf0JK8qPWaHhjo8cbxxB3ZMzhgfMkixXrm7dZxqACJz
0LTjAf0gMDkbNkPcsZ5+R8frlaTldyWCvnetMmfeSTj7CazPKAkLoqjdJhzd
MfbkfXtSUSXBmElSoXUNNpEhWAe2wC7v1gmNmAj0ClfX2i4Lyax0UqU73vZT
x99brZodgJ54rfhatX58x0/D7dpqJWbFBXvoNgVdavQOxA4mBSZyn76l+7ia
pP46F4WNeIF6Fgy9bM11r4/doZZLfz7ozs+8UfpRzSG+/viS947OGUCrZtQ3
EBPDvr1PUT7bQWbTjAhCOMKimXIf0Hc3CV1pH7ThLJWA1kxX2VKIXH30h9/E
oK5wX3GpH9zMaZ8o+8lvF7L4q202FqoPug9BOsQKqG668oShkV3FOGSakZTU
eTki9ehv4RGEE5KRbi7gnV4ELhhf2QXjHA+Y/BgEA6eIQcsydOUtEe0kY3/+
72XFuDZ1bwh6BwN5VpGYPwvn2e3lEao48VTESl6mH/ily3fqngUG8QGCx2ZL
tULkHqssMwn48eCT2yPXcAP2+bnSGTT0j1OIr3XXXMbazMRnGV4+bw2OmXfG
xboa6urLb4k/Sgm727vFhtgaXsFR+pqYaH2fdZ4fHN+Fgol1ToLhIPnoP399
oqyfKj00HhiWcK703Sn+KHOvRuta8p0WsSlCtXrekKSQeS9Zl6Q4tZmlI3WH
CtedtT9B0oCoNd6LzDBdD/byg7UTjTOKy5ZIR+Z85OAbwRp+MgqeHk4MVelV
80xRCSd4Dgq8+NxkmnVFqSwusfVrRnfa6ILVv1Y9PhCqyBhAHr52972N4lFm
2hVaJx7JpX1/pBT6+YZq7dr3nDD5poBij+2aBqIF8ck6ImqdPVVFC7TrYcxX
CWph5JdrU5JPujJSDFTGMud5NMhbPgSiBzKmYcwxgvn3eTT+QlNVVAczS1eB
GecHchOiyky9+Eltx6e40egXDtgueTkgq/czebQ6KxMyN4G7ZM3GNHtY8yoD
ntuRXtindRM3Vkm+KoOYldOlUm/y/OHZYP/AZadfAlxVhjsqMIcvQrfmuXRM
P7tP2hGmS0daMpLhOQQSTrwxF++4BxpDI4Mj/Bv9XI/O4k6s3IM+FdObhdXT
GMij4zfIwrJCGncqBfVhKMHSNvP0Ofvbvwj8xj9HLZnipKVUf2b1nwWkZSKI
h2EFfzv+roSV8XWYtUi3h//7h72udBNJNPYfiu67iTjK0feQcNPvmLYyhkLX
lsQ7V4OVLnTw75qDNwTPKvUbaOKoLuerAO4wt1xJUZE0Eo+RuPUfSsqFPlNV
BVtrK8BWXSN4Sob3CRnDWSiZN6AoY43A1Xg3b6rluk88fcbbo1Gy9l3qX65r
zSN3qXQGwG0wwKiqUNgDEsgDOj4fE0/VtUJla7yBx8GIVo5NM+0Z3q6/nRY/
b1nqaMCmFMT2bpyDFoxvRFjWkujrxzQbPj1loHrmECv38CEsrSmtYVu7dP+O
LiniUIBoT5pDn+JTFA/p90KNpVlAfsCYo4VVoOdUwQ2nKiyaRQyn7gal6egf
zeiraZVNwZds4tRfwG09+K9mX+jH2n3ohKzn222tbYsJt8MAkTU7B9vpfgd6
qX5TFLGDzlZI3xw0f91CeBaV+kwA2e0vbmqy7XUdEJinJONVqtQK1LnSTMmJ
OBBxT890xRQmFfOkLNXA+LnyWb/AndQz8QNFT4Pcoayo4VibuQyoH+qNq7iK
zdsqc1Uq0FINRm41nhSDhFexeiOXP36NZXFANIluCqdI46lFm1OvU4sNH0Qr
zjXBjg5hvHt/kBS0iQxTYyErw/LT6/zi1Px2o9KI1Pd7P40VfzMeP5zyoOUZ
/P1aRdH/p3gYbUzkwhLIB6KmGdh++oTTvlX5TVcJKYUK15hKsxfaeZINhEYZ
O+WiKsDTIzET2cuzmnlaJN4lPEKMjC+kzDQWOCI+262lFMPFfu2itsvr7AS6
+izCgSL6AwL0F1MCUH9/3MIa9kTGhFV6bvTigQfvoxtg5jatMvQf2FvDLlly
FUbOqchSCLmzuVvh4EUyXsNnzJKu1I173DNQN7Mjg2/20zEF4sxMdL3dPeMF
JyHMCw52NZfOpbQWn0sohsNkrjAEuKCYZFfHMCtaiCxscFEqlULXjkopqACt
nANrfw9GksgDVIkcwagskgcyyxFz/a6ksW74KERRJD9ZsJVB4l5cyJLffTge
ZQdPLSZSyNKzVMWX5P8oaYlV+bW77JVMVGsal1/4lH1wfsJJ7TgtBHywsV8H
51NlNZHffF6PWHIFFHrQ82TzadLlR11W6Wgtk8eJ0CZf6OEz3vQgb7CJO9Ju
dhVwHR/+sMWMWFA1H2yc00zSG92vZkSRO8Qx/SaIveWPND41G7My/sTQJuzY
w3s9CUwY/YX6bhsSGYDWMNQNKZc9y+5e/l0OOkUXMcRjbme2ovTehqiUr4X0
Oj4OYMVeHUL2e4D1Iq1W50WpLvJLoWLeG/hVy9nLeHMPJX3PlZu5dXgOefSM
rSVHkNpsvTWQDXdsHPC0TEa+lU+Ft1gQmdWlsSGwXW2/rc+/EYe15xy5dq7k
JS6LB2DSB4qjshmj22XHTV6qHV9R/sg1cOyqVr0jqv4zSiwpmOWLHPcKeftb
p6Aay5IdoMQk1/XU8zaFqeg/oU1QKUxLJpmfd5hMhY/6bHvl2nA80XFk5Mma
XAwvFV8BItDxCqdQqknYIU/37UyfVDidOEpXG2XcUwcCSezG3gKQmdH9FQ8/
XFG7AkmhNlM7TMozwaHeO8pm5WlZ4EHeZRYbpKJeIvBMsM71OHNTvcLTGqiX
ucUXzimsEB39sTmifo5TcTcWcNEF5W0KtUER9+EGGrOvmwEK20w1sITza/5c
LB5jlCHce2E4Rho8Vy/42bgiCrlSwZQ76n/73QGHqDe++2StfLR4lqqhVVOJ
V3oxty3wk5Tl5hlFJkyCM6xAD9Pgo4cYI9S3BjuhhAdN6yyszGIbNQvOdtH9
VLttuwP3/UUwrx3hF+kufCWXKLPf1VlQhNT+UqwCr3lYSxMnT9Ffuv0ikP08
RgP5XsLA/JMEhKn0KRUqPpaISyuoacFNScrXK6yQbmASMGJIn8g0pdz0J8td
J229BYXyVupENmfc/ZPzIwjFy+NEfa9X43+8Apgro75u7oC1JzPZpwdwoptq
33afH2+TgELo4Y5zHc4g8GgbJi94V9TsmO0mrF4hFvWG5OqTwLFUkU9IebvJ
yiK9kxDEKqPwjWD0X/ZT0ncSCjksGGylwMjjqaFz9IcRKw/pGSy5h2cDhdu7
BJFqgq9BQP5S4OU8vWYDdhhu9Us1s5aI1ALze7p6JbR/Y3o6PaZJVNE3V4Im
R43Ii40ykCrnA3XrmGRnHdfQg58LvQEREFpfZ1zEBy5kqp8zVtUVHCrZl5Yi
90gQojmPnlzWnbgMw9YrRj8MtKtmUF+/p2eOp6/VnmF6vFzZyA1Lj8YQKFH/
+mZLVdzZ8pApELa6jkEIazsgXkNY2b2FuhKfKX4eLqO4nb7gB6HFUoYpC2f3
LkiiH+MHr0pvLw6e6PoJV5RVighGMrd+/NKJSq9F9TmTIkrbPdabQBkiwjW7
6AX3CzWiR9z7AdtGyCyLJ34Hdo/f08GNh1PvC6/QbzCbiK1UY9KAqTTKS3eQ
hwcifM1KZ0axxP99A5C/eMQujvLVoTTZKb2LgNsbv4G2TpAcbcPDl1qA/cq3
nNL1BiRj03ChDvHqHKEUAnUas1zwshF1hqCAupHCoA6KtNQQd3YfFKhkDAtV
8JwY5CPljReTctZl4z5TCMWt5fCmNj+EQaAUWwA5PeAnGHhGIdBmUnDFC5aU
YQ1F+C3L+lXtUgv9y/2/RRbEUg4kN2BevIfkUpOOCEg79urBuj6PcnvDttqm
bCX3urV+Wmxbv/vOdYW1R/aSm3h/FUsZn9rxiOXR8KhNNAeoTIMdqo6m35M/
7r1rHSn5uwMk9ZqRSJOmCB5D6RHiTFhZMaNevL7vCaw7heJM2yrCQqtzRk13
ePgRwllrJLe88dJMC1SRIRaR0Md7JEif5BwmrPR6GW8J6ehaeMK94IReu2WZ
yG3NNhqY+F6ROWL+jf0PDhPH1VT6d0WLuBCULHS7mMcGaGLEGgnYUOVFuEDV
qrJv2s12y6vSao46KBfEx+zsVrlQikANYG/1JuO+oNu51QfYkchR7DhdTKsW
vADX6scFMqibQrrLn2XrLZSh0sm2Zm0ORvlhSr58MsIfHynDw8vOynkweHtH
CIGdiwmJXo+V7FjF0VhLCJDRuO5gnNN4I/x0kn4XH1M4tK0xIqeLwZlejC4r
aEKCesth8RqXmrQM84qdVvnb3Xq3eC8VnXEeioo6e8kHGK9JI2rIW0g67wy/
y2GxuRxhgU4cGIyD6ISXQlGpTO4CrubNZ420UrD7TtK2/TbDgeytbisr+QUw
R+S0lBM1+GRCzoHXjJNhnwcwu0/bn6/nLXfo9OLp8GOgZh1QNkRWd7bmKOu2
cPy8/D16nhpZSWIOowAFmiK0JeIHxiyiUiyoJx+QEpbmW5bxym2abZQaj/Qx
5ilnFJqnajXOkw8Hoji5vbEKTM5EOd77xn/SU+xRy8EPyMoUjQFha4egfcqM
6233Fu3g8tJIobgYLMHXNhhR/r55bPuuopsqzt6aY6DfivxQb6eaREBqUOEa
RlHr6IZDFdHgm2MN+OyG4/JbFVNNHLRzoI9XIUpYzRkLOa/635ivGfcomyRJ
sIGIjHHEAE/Xr4sphVwy5gzUg93DzGisEJYPWx745j0Anz8yZ+tp/zLJzuXp
XaJ3GQR2y3KqXgIoDAFty3nM2x9uvi06/N01sZxaWZ3b0kxZIfWmzqEjMj14
hfuvn93LNe43NMaLLeSBOmhN45lA19Fo8EqcPMD/L/lW12dKcJLPAB6zZn+w
EkcaD3bLL/AS9kbmmWgngitThGfYN8N4K/5f7TnLqz83aTEVnbB10cokBmq5
JAn2ZAFMcdaPQFfxbt99kjcNibQryYNJ1P4qMSxOP979ha7OrosGHpUc17y2
+E3yNLnTuMSufshCPR2Lz85FdSnPjQex6+zvj1zGUYfoCnG7rZI/9YeR9kfw
/ubqEEJQtTBCxB8+rgA1mtvFK4j0Pxc23DYyW8jtRGnJ/uQNV7ELS8QXXBsd
uc6iAqldeN9yYGi5fpFdONh1LWeTs/Nt4i2VkNJYCit2dI7sLcr5kAFPCWxB
miuI2/pvEKbRlQDoVWPwUf7xq/XwH7ZOKisp/QBIU8Cu3SWoDh5f5XKe75X0
z2y9r0J8xxUnSQ+UcFBKqrPJgWRn1B0vkZrddR0lcCKDKnVmuGQNEeteDqtt
9TWQYfhWRuZH88RzDOd2mlsOnQS/SM5KikSPKj+C23hMEIQvYd2Wxj+Hcvgs
EElnvGt9NUM9tmsHxUQ8e62dRTQnHasaW7wyCwZuEbuwind1UmnNGiNj6NGn
HEKlGqnPYSSnEaJOaw9y0p6Wen27/LXipDfjHCek7u/UTHtStu+27h2xVIi9
+ZegKYagd+Jqc5YOWVrQ4zrbE3JsmS0/YCx1HTUbuCh0z4o4yN84C4PfukWm
6tPiSeMfgGWEEUctNHDpi2BL5Xl0+2SZjUO5cKgrhOv/OwVgPB4/Hi87+v9p
utipRPODrAW2HbEqgM8VtZbiXQN+dpPTIretsS5wUHO7k09PXfQgnk0vZC7c
BYMaYamycRObTowL2S1dPC+q50S2L/Wc4RYeF3YxdceE4JsMe+Lu3cX7BTG/
UZj9t9E2QnuPrxD+LWrDxZemkWSukS0x0UaO8tjqvkIN9tY9G0Uf5/tM9D4i
cNTx7GeXorFUUL1krDXSvRR1nZAu/yRp0Og4uWDlYCgUj1ykda8phBupoQlO
z4SkCHtyzCTkdgW2lwW/fkFPjiRBSwhfNP2qtPSyP89zCsNzGeI8XfU9/E1y
L8R6d2IOJnjfAqyJV8QJd364Tv4x265wXzehBM/5LCEzenYMjbNu9mB4QrZt
Mzaq3dc6hVlSXe8PgOIGLxwRGs1DdcefF/cqnQeEf9CwrKkgYgBO4FZxNHF0
Nv9Hf4JCEUH6Kn+w1Fpjw4mHgiFYNIKspNW/0OCa2a1iu2SOaEAnJ2UH8viQ
F/3QYcf7VN65KW6RLqOC5ef0/5xPYTviAqxx32inqNj5yoQvMfefqPkIlOQW
LQKBcM7jatGGH2yDZY9iANL+Vsnq1UmySOW59DR/7uKjGnL05BMPFWBp4+5Y
b43k/04LvIOq6JAiZZFKF3dIVg+waOCTwlLftEOU1yvAxIy/2r4a2zIVkjiw
BDM3Ritop8D8WqYZ4KBDWl/4Tu8XBdKxUgBgjFU2RaIlbtAnGj4e33d3bo9U
Fkj4vl5PUz1rrMTgXOBzo19gjH16Zu7p+e32D0ki1aQ4Bt9kWPC+F5ZoNDpx
vJu1KKGUrXn3B5515z00HBLCFHVCy1t7aJftG74C04nbV1XzT80Jum0vdUDp
5ir5+UmCoJj8XM15HlwtWpOMz9sRtcjME1pEyHd8c082398I3Ge90eM4D/Be
I4IxWlM/1i7EIZHLsSw1YIOP+j5Prpq/kFim+SHG+bMit4AuxcVRmOWZjhFq
O3554UF9jkrgzNor99A6EvvMZKneGSVL75qgsb8mEiZnoD9RrJr7sbGG/YL3
oPnhP23pfegKYwb7QBbwPyJnuzSzJcX7oyKbwAaTVSoib/uDMpfyKutyK2BZ
0zAbWg0IIk8kWNhZKZe3U5K8wOhzxlZrU5mdrwCTmhsxftHTTyTMmUWjLHVE
4pxE/KTKqStLeAhg7PERnUFw2r9+p5C+FwZ7oaCBYih1l46ExW2BBIIRLcnl
9D28l7zAWUWkevE+9XmTuhqcc8+UYtSBBu+h5zZZyazpjWLovHxKL/2hCEJP
GrkI9/Rg6VNWdaxzO0fJZdRrh7WXc8MlHonvLVIalsL5+3L2LmbQr6wJom+g
bZI6BTIj7XpcAb5liyT2bayUcXhFsvy1ulsiXypvku39xzhme+aQ1D9cZJQD
WyFLzREBq3tgMG8jDCXlR9kT8mk+495p8am2dWDSWCtBc3d/nq/13fTemZ8x
RTSId2AwtZaQUKiOlLGNP5505Ln65MJKNSss+g0bhKcwksoJH95Q5q+hFG6q
0LYQQSWa22z+v4IazoX+cqgVW6UKjciqzA58mkuD+ACviH3FtQcxhN8lY6jc
0dAX9/XFLRkAl1xbcW3++qIlLxXw9OFOcl+k1mq/gW2Hfl90B/nU8vIF8t1Z
R/9X7RS367ROGce2eD14ULpmt1247CxwF+RuUV8SUJJOsrrR+TeAPCDanNCV
xe68arAwCLk1HPMNcA188wXWR1GsU2NQ3aLlgql8JzV434PX9OzPrH9kQ5FY
SzfkeH5ZsvspUbLVCYAakaV252m/loUiqEgE27G7Bm/bRIxxPzFQRjWn0mfK
8WncLmDwZEnk4K06VmfTXY/IXoQXg1eVrQdIKmBnJEpQZKtoE1cpe3Cj5tqd
cstZ1HCpwEQTGEKikeur1yhvpVY+Nn4RuPuqEvgr8hOLk1YEEim/veQl21QL
HdwxceDR7G9ZeWzvRB79a9QwYkuaI5kKivvkukscL7KCgIDBjIXDqwcPozeZ
rzKSJ9UwvEE4Hd0fi/bkIHaXoA4VQPAywWW1qfrEu1lxqRDnzYS/MhS7LGGZ
nv+JFGjii8/Qzerv0OUUct0dqxPOSP9zuIh9G7JZRQHqbtyW7VmT4xMabQqo
UvCDGLAythOy5ajtynCH3khjnWzUEq/LbrSHPUoVhutvL9IeuLrIx2XtNJAG
YgmGNP1ty+DHOuyMU9ohocUm9kurdaJzNumEoy6fIrXC0Nb2Re7/BxLC2KC9
sf7R6oDlPEUzS+n5iVPqXJekjyJ0gHd4RYMkrPRYoqd4W7sTfNEFE6S+uqmI
hNH6Xy6k+w2Qi9LUu38oYPeoIzYDR47hjiEYnTLdbhukQezM7vLw3zBUR8sA
9uhHl+uSwXI0w5yP099MhuJpMa/2QYEv8/vsO7TswaaTqApEsSwodWzOlpGK
ACiZlapOdHXD8ujbW2pnb7Pik7/0QZNds6yChi9JlD7fM5qcZjv/wl14kziY
Zlsshp6WzS7I3XCCbVTVh8ijyRhfOVot5qk4xcICTyAEzN+EnrBXEzpOtKbU
y2jtfcNzMrVslS/goW7VBXp8/FYzEMTvV5HnD2xmPr1trSTORWtY3+zrRg5F
28vbMU0i8ZoRKlXm7RrtaC1cY+k0sGdeBV8UqXAJedSu6/yep1437JuCR//6
6NHsiTK5MuI0pDNBAAP6tf4HcSi1LfBUdAETERcYY/v5kWDUBRFh87WRoI/W
YVger///EFI1mJ2nr+lgNgS6DC/Z3OCrKVjD2CA5Y1OG1idiOZZakG4Bjy2X
VR6WsadbSDb3Mq5WAFBi3sJKtrJBG6b8DNXMkSju587R1B9odNZNIyQ91LM6
97I+EjUUrNIrLUzwzKufbGGjYW6FVO1dfJFxJ1R69nNHomWtdat0NtnyW4Nd
E6D+VYX/PEFxlENU/zzLY1jFa17iXSifjiCNgXR7x04opmlEwP2hV9pF6rii
PoLDLnPn/YrBarcd2RGxP3zhTbYNtczUm/lhw8DYInoR12OjnIzPwB2seoYA
sUmdSEHnEc9WODDxuIjVpQ5w+aAezWP47onrqb5YSUmA5IJPto0Qw/fZma6a
Rq3LaTsli/GhjQyHxfuoaot0t3Rp6KYW84uwVHn6+9U8dOgehJofAH/3IMfO
ivZ5S8u/1CKFpc8zTkzqdKeOX2Z55bFQ77mCFsgF0kVOo9MAXmBUhlrUSzYU
o6XaTz6bkrJih+oCywABBfuN4UepW827iL/vpWv3uuzt4BFU+w0JT0DpncC/
UYvcXURJ9wtPhoxTt9Ms7jWSppZZDfgNZNY8Xa0CEZeAz3UYrl6QvqRZYcrK
I0J4YjN3jBHwskQDpZudMeL3ALz1s9j2vn/ZlQSmIe1/bGkFBjFBqTQoVaay
ZDKDTXUIIJ7GxKWwA4umBYyPhgDnG+vKXpXvd6eZmm90VDTktYvCg4CxNEWx
CT5B4LoLRABt3Shn5zb7hqewVUnxOZ1vMw9bgtRxmlqa8scOIAc9txd8pmEJ
p6AbJl2dc5W+2HqlGgO7xhb2bl/lOl7geeeu2nHULaODaegLlMopw8LIepdD
pqfMONDP60CWNdcmiSJXnJpwkkIwNUtwy6wCyqFnMLyLqRS6pa/zej06xBky
4KqPX99PyNj6xh1ZeAzOPj4b3OuJNT9tgBeJfSoPFQvjL0jyP9540E0IR3VP
QcHqoXdWj7fuwrXZ0tcB2DQVLg1eYO6JAN724gnEQ4NZ6plAaigtHzVeB+7I
Nmz2QBM2s2a82UvlBY13ylZA0IGAnLswNW14vzwjoch4N5VIz8Sda48ILthR
Sh4gZYAjBh7Qgbz3MtMmS4pA9sROwQlTVeeahNsbt7DJgqr26l97XD0rCZ/w
kyqNYHStkjhAJo2ezPgBB4R8yZycNKsU1dDjvX70GT1UMAc4bPgQeYrlDrD+
OFxLj/wj2S7QDaEFhdlF1aL+EgwqYrnUM3VcPa5H/xd56jyccPktXxGwX+Gl
ACCwTuBQTvrjDVJNLJyYpcVp5wV0o2ixgWIhVyCoUBjQ7ZmPVYk4gHA1JGtz
FllmLBfJaFSDkc5HweP2ayPrR3AwLroIzxvQUZEWAihj81JN0r1eqzFbzeES
nsfWyNGnojD6ZiFvB6LuZSYONjU3OB/NH7ZYMidaVk6yneF77Oy85Gdb93EG
WLXXH99nhKbxg2VuE75Y6gZQvW6u6m/g8/RGV5RUfRjijOv//gBiK+i9KKZ/
NOohYQO603KB/T9tdlKx1wXgZADN7ewdss3g4+ledveh10I385Ni9kNsWqeT
uJqcGvJARA2sWtwxYKcNGaLOp8itE+/SX8ucIeJoSseplf1ZvlHRh8ignuoo
Pgm3a7Dk+7rAp9pmPprqaBpCwnj9kxNxZCuZUObfVEeUDtiRRZP1rlkHd+aD
5WaG/wtKA0slluCfIYDTu/KrFnWn8eSDASb9yvTm31b+DeRZMNx7zDx+frBg
ZNTa3PQex55rE8tAKxd9dasGA+9MGxHXAje3XFQWaSdj6Y3NokFxfePaWcos
Mh8SYMqfwgMw/2IqrpDO7ReNx3PjdDhqAoQxqpH8N+CiYd3MvPbxTeRdYGPM
XZYq4r83fkq4m09a8A1W4WAaveqiuX3MqWM7KfVG4F7oetfUAQtwNPN7/xH9
zxI3xc8UBj23LsspzMs5g6kqIdrJynqsV6KjrlICDRzmXgdHvqZUMOENuvfb
2xTS70FKr11y1eOIMRWS6PPWguXctEvFysVfGgG01LB1eSbKYmOK8LI8sDoO
ky9kCDQnC3qiq3P0HBttg4NqQ1ZHeLCmUZCL++6P5fbZC4Xdyu14TWX08VWF
k2uXPacehIQl485tIW3dRtQrUbXaHudOgLoMqfc+uF4xS+PAzeHk+Mg/GuUv
SwrpvCFrxbcAMEas8ZG6lJ2+0d6Ww4zxhSBrOO7npV3oLs04Ied7dDlczWGG
ZxW9Us69IVZ2piKvIoCk98zm+bqcPB/EVTh16aysiCo6mjy9Wiz130FmKDB9
WgF4xqUcVQu8OhJugFnMHhx1Li5fzzhRm/t4NzagGTEydpIwZBFtjihucysc
WUmMFzk9a/Z0soE/rljrLJ7VmBONdaqT8p8+ysUZ6WGEHAsf5nih4UbUuwod
pJluB/BY9jQaM6G1ShWfdeEKGcwAtyL+qIBSlfWgl6PmG6KnptI9non7DxM9
Z7vORfZe+P+SjLsbTWqRu6ohi+joSLKDhDHgdnWpUKo7kYAlftwXMw9jC4MV
exz72vNyRmPZMZFllAPiinnZGBeyXgLwPqKocFDt7EgGNSuMWSDLeSzZZbla
80GD/rDRY2Bu2/RK2eKf35MmMZr4Ida0k9hhctcNWZcZEqJ1m8dmUWdGbklt
sdOokvALNjp5/UmqaWL9MbEWkQWedaTxlEkpk5lnkf92fo4mpdi8j6g4vuCH
8CW94xnEQHdp8LaMDx+FV8SN6SrVVmMAplxtt1ZPWSnUTm3UM8Y77+3NYyhy
e46fwbTtRBHtKLy3Rsz2xm7wzEUPAFiEwEuoiX00HvTXkZonqU+mNikYNEeM
vxp2qBGiAzYJJwsdNqMBeG7Z8kKEPWpHpKXR7Ft0jmq6xTV26D+A83iwv45V
kRHEOF7GbM5SNTOtHFwzef8uOpAPoMDS7KwNrbVE2bFHQ31Wm4AIPPeXUeMw
ScHN+ezzwVVyS/XT5rb/LBRji6ChWGpeuRAXPic1tS8/dwJWbfH4WMFIQpcS
1EBNEmVd9d2n9J7A8UO3AoXNyGbPge3PNaXa79Ue1BnxH3J4m+vNI9yKv5iu
j5j1jMZZpNBMhXLrA7RKDHMU4yI3M/O7YfQMG/SmDNUOlH19fITZymWW3GoI
xUGZr1d1gn/7Mr4ijzhvQCWGqKNjKajApMfnQ2e9u75Tc93hKkjVb+lQFH/c
kmylFfFt2CR4oqz1bSaSYbmXUuFfyyJjoI9m6blokgXhTls1y5lbqpFHa57R
kRsaereYV+YO4r0HwW5LozTMDixr+d+pzpI8UTh2Hb031JYAMBEo02apBV6Y
2FEV/GRtnyAFsAeI/9/YJGlZRMfnqkz9lt7dyRvqHgOPgpsPpU/8StfC8iu4
1EU9DdaamEVDZVR2nRn2BALXvKVrfTTDFH1+DA18nsP/kD3w3EuqiLYekkgs
WIC/bGYq0ulIcxt2q3vVVgPEou73aS5tziMQFOVQuUfGh5tTQULpNceEwY6+
wUdEJ/BnNGDR87VrFYA6LqJm4brLh8FYQxasKs6ovfA59FEN+TlZbwuztdFA
e77BhPX20jIWJpI4BoWjE7EmGbooRnugQokMY/IrSNlmkIYJf751jbQMteuy
op/NmwzdJB6j9yi8hP30HpnPG4LZ0PMUmz30Xc/3dM8VUwILDA14ruw9Uzy4
0mCt1Kouyq0H3qP5oxVm74Kn8bHzgl4G2qp4D4CKZ30M+CIY7KOHONmMvrZj
s+hdoI1TWoZSvQbFgWPf/kp2UlAoi273A6GMXHqPHSAJwKsjpskFDtqdNSfG
r7iaHMw2ysT8B97D7IgxL1gVqTy39LZfvqZ7GhgoZobUY+Gz/hXU5/sS6VFe
4L8BQ8SJcNZc6XVgQ6RM8e1TlMCw1Esf6XftAmV/0mjH4AIQlcCc8SYO9NIA
gBharrQpQLhYtC5/+ixL7pe5qm3gPZao955lzZz5FVKz5d/LBQ16BXAMfj+D
8MNYZ/ueSilvTeob5XcrJkdOzH1WDF8h6yuAWxEQF1Yu/EKHbMF+anMpenjF
9po83VHY+ZOAInP9HkycEhJEpx8aA9D1NSCtzmE0izAbZ7BaxvFdFGs5Rrom
HVNfpRjpB9EkwgS6gsL5WxYXszIDlsjvzedUSVjQaZF9D5MUAHHMSpqwqKUR
2W440Ai94bfcCSSlUAQIPhwunYaOocPZM6+KmRGSIimlujViLpHbrODSTL2v
IXCRfK+57aR+kQs4U939rkngNrK6coWdUJwLRPfEMQPfyR4K4HsII4mpPR1f
xbp35RoHHL55j9qlEUgStzCkcK1paE/H/4TN8VbaN5F0zLHq6u4o+SoaQl3y
l5oeGUPymNUTpF0BpZIIOpJrFp4N/e/TvbDH1S0s2aUkCbnJOD5NnqwO64fR
zDstCTVJsN+fnUXQocV4B5A+z3NahUYpmODkr9fjTwNn/o2cNRDIaEabzada
39PYVS310FZJjK/iknx1qoS3eNoWKQWUL1jnNT7GEubo4QQkvhTcQsY6AWBb
OJzawGtglkKoMzcXtsVs4QQpZDEjUBl9lEULlFdI0t7FjV1jk3dAwlROTmsL
9vnI6Q4qj4Bt1wNy28XHOqCe2zyfH+WJYKkHXFQvpJ6YxC4W8uHbcVtAP03O
3YLlKYrBrDuGWjUMW/QIVUzYncKuxeo0zwnyfc8TrOrwwEhwvgpLvZu6Etqq
sz5PHq/qVtqDGjijBncHhhxBejIDIDYWQ1brysWgckftKZIkn9SeuJNAMel7
dXkma8rkp/ESrK4Kfva4TsMfw09h86OnqJ+sFTgcezwXWWNdYiOSmqMME096
m8O0YvF45O5H5nCgAaIJoRHvuRmnam78mKrHtWeeUmD3cKjVD96TJ7FSk0rw
HaUOCWbJzhK9oDN07YZy43DcNIAdWTmGi/4sWyF3+l+NZ55442yePOjJAP11
oSHrM7fc3K+Uc4QXF+5aaahCBAY93+0GhnwsvM+r9MvjWk8i/BGX1casArDb
Se49IjUal0IvxiYfOJBdunoiLQ8STp3NKDC63L9QUr6JOBh/DLmMhCu/Ns2K
rfe7XDb84mYSj4yWBb5qrDtwpgWcAOnbFVfdF80JVm+olfuxtzU88vmn7w/0
3mQvb61soGBF9wggbmh/jrXhtF+yE5vCh6DyfAklgWXn4iatdfiVXlgTbvsU
siyTeZcLq3RzQtkMVeHfPEK4K0umvy0SQQZbfZ8HNgQc861cjusaaE6/NrmF
vqVdNzXrpo1U72DmTrgRWDVJfT5Ukvvsko2keGWrFiYqY3ta+5E7yQQW1jqu
Kczf8vl1NFUJS63M2KajGHQx+fUAUhs6eVz0WIU7G8azPMUxCfypSzAjWg9J
wBvh+iWFsEanpfOawvEv3D/iq+pQ2wDNdzRd7H7/aPUVXm+oy98qMwwoeHKT
2nNGjBLnnjGBsN7qYIPtdmv6EL4p5EG+t9MJ1fQhWDZTVATkoRLouKA0oGN5
xna/iUpdHghHk81X8ehJf19I2nnecrx4EQzw/b5+ZwF8zRUxHk3896Wd+Ymv
dHCWlj79wAQSpAiaPvuZpaJnm1IjP0Wt3RK5S9j0WWhO+NMuVM7hZY62/Bcs
pdT9ysuPMOnqOndiNEEwXHg4lmBczNOGo7grkTagd5sK9zQ8sj/HiJkYWWBh
LbyrEpsU9ComFidorEtxoC9oxDt/a4vy4AD3xc03wXwwErjV6OJAFlNx3A4p
AVDUjmF7wGNBIqdVVCj47uLCq+WBBKwOaSWDy4UCpYe5gkugWxoGmYm9NDPA
4ah7h3iaGIqhNR23Jx6DCLqCcgmkAJtLpNcJJVIkyDV3nvcHT9Y12bM2cER3
0SMULSbhTitQDIUJROjjdkdRhwM0cndH8UCxwaPLVro07N2mBEdm7Fb74j5J
TjqDyZruN4Oj1VDltHtmqZMb/gHnY+qxH+hYlsF62Dy7be+MwuvCFNXrf480
NXyURML9mrz/vmQieqnxUY1NA0qcRXjwfqvHMloWDvoKmv8idfw/WYVvv4M9
PUORtXLVVMHsZSohSfmxLJTwn0SgZmHElvE2iR+hBHEmNoXfuaNSj8VJRfR1
OFlD2QSjq6rLVrQh1/QoTVuGmdsbiBkOQ/tbJb6q9ep04ve1RFpDPVzGr1+t
Nan7OuaG2Z+J3VXYddBRmv8QbJ6g0MJ+9tG1hmZ8JJgJTOl8XFoKKTA7JTCR
7Zim5hk2t2K9tPnwZ+ofPPyFYd1Wmerp4JPHI8cfgzdhvbthan3r7ww2nxK2
BZnejLiKFiTODuvXar1tBDsrZ2JrRnyyR+jJVdwPCv8LwiLAvHx0l5557jfx
Xn4kkUxAxlkQALc+WAXt2lsx9tNS0o3pdRVhm+Xk2gVRVIsyHHj5fDq1+tew
uFpsoVlL4g3GOIFqLz+k+7Y6AoQ8bPuA93oS6VxP4wumcyq8QJr2nZGjoOQf
9tELT3SQ2qTm0xA0UyR/w1OkmP/45q4kQfHyAKdfMAMzXRosxa8BMQUvnmlT
XiIZnQAgmqQb2xWyQ0x5N5mNViotesW9WUMeBXkoCAppTgfnEd+GXzvZczG9
DkMGwewAEyYWaljXEZaM+580kmZ4iuyPQxCZ1NXiVjWf1A4kxig2aMBjxFY5
gv5WwBvgR552/F5LMiQWwCuWOQcllqsTQ9J0tjTS+Nu83kl6QrgljLRC7Ey5
w1WRuopTf8gg5Sa9zcdlh1vgujnZJzB22oSBZ1Xad9rQboKpBrolhZP80/pL
K/H1BymOpQ4Qk0Bkw9bfd7EBhgfooU9230fkVfOiUFriCXS2w2+ytzEl7Iyq
og8Z6saO7xl1sw+YWJOlPVWBz9PjcAFv9tb0B6LfmrPiVd+t54EmfJ176850
jL7L0Cx0OJptryOu6rcaF7CCONx4daLUh3C6E2VGn7U2RtRk66GBJ9l5VB9m
UXeQ9xxmSuET8wkGD5wVZFdwqLt6hDL7jc2/DJWplzJwnq01kucf9xtscPXy
yzSHa640PXZLE1RhOSLju/HUFkOnFektGyK+/jBDFHdPCFsyebNrpdctKYLR
332ibQMc6NOCA20fY1lRHOCmSxBiXQ+R42Iv+TCkrL2P9Xblb6b+7MLcuXN8
Rvp55MZ2Ia4ZvYlNT+ScFx+8iAVbeMbjU0V4uDMDP5pRp4bjhO57hUYTVKly
ySkifYACeydG1q8cuMyKNZ35tjuWppuZB3DVQyAWvrhNHjakZia1d0rU5iev
8Wrf5k5xgTL1aUL4rpxoV6jsazZmYhZlJRlzcOZkLpfDxkv4r8vzVfQs393c
VOHdp9G60/XV8OpdtN8yytNDrXzhuQbeZ2dOEfW/JwzBxtJwc+Qk/bnQeaBT
J4u8U02RPtr58DdLMpBfINY0sje9aRUphU4pNrU0rlJh/FHClcstSKazeT0J
VzfRrztmyYl7gMvMWxGUB/H4p9sYGcfJrOVZc8nTXsP0SVGde4t52MoZATDo
F+WJGONdhI19oPmsaVm5XSGnggUT+Zm3xM0zd67JwXjEkHCfnRHPB8ebimYx
cmAGUMncPYR+l5EfuZ2pQOhx4Nj/WhCzc4GS5AcSSVsySOpy8L6caPJ8UieB
IIvp5It1tpNzyZwP78gVkibOMJmMdMP2Vmb4mmHnS+MF7+8SyOuRXuMPCmNM
FcMTLvwvEkjMVWFG3zASEOF+YBSJ8jitUcywf1woLNWZ55/Y2d8G2yDA00Px
huNYztXGW3Zgl8JGCSd8d8ctu3HRT/eQmGg92TCezrRYBTjm87hJNG+8Yj9U
Jz41HSfT5JW/RC+nUp6ZmNAFhRdRn07mwBWWOhYD91bbfWtAtDzZ4P1KKxfJ
Otj+m69+0sJazNbFxkVq6LEN9FHfXfO8aGwdc/k9B5ORxysMqKGkjbxtnAPk
F6Hai8rjX7vuJl1Bd+vuO7WdaClL02XvyZxt6qmO8RtRiqZgIVapVQgXuKRY
YEnMxrb9qa9eIcbzVN9M0r1kqYQ/nqV4pFZ27o0TyFVkydaKPQbxi1V/DWpY
E8CqeW/K5mhJ1BlByTrFGaXzAgQKt0WC+EXDp2WYb39TIjDXzIvkHgLrogbA
1OzlhN/1d004ZL9Lwjj43OC6BM4M5ZVjnOxcRgO9ENS6AV1mTe4CRj/R8Sgo
MOa8eMHkOJ1WrUhf96BT9tfurQeRq8LD14gi+Qscs5eOHct7aRn5WbH3aY9U
5QuCajGv9ZZt8MmcZggCglPl9TocGGuE1f4digPRDHs7vHGUmfkjDiJnPtt2
FgPwpFQJvRsQaPz93tzlQQ8EU9oR0/0EnXWTx1ketQ/z/rUB1lCGd0CYJ28x
dNEWvHqXDGGvwO7R7m9XyH4VYnw0dlv3Q3cGvpg3sto+mxJ6/2XrZewYUytO
9GjjDzYZ8uJCsGbM4BnXwxTY3KYWVh9koLKWpjF/nKfwZPH1KEwYHKDEKg4o
yzQxi5cyYJkmRicbK9ZyzDEwtN0XY/usL6aiv6HU4gyyLORt0ZFydCQrcRpm
SarEBvC7XiZd2FCSB6pSa6buYpApwV6pXIlWjJQvIGY4Tzl4FYqpBu/7K2SX
FzEIvyXYIA0+VGaCOWota2UuuDlIO+nYX45UkTghpqk18jOZipC+WE/7fVG/
AYyerdj0/jJS5qx69pS5OO+Aez4BWTJdr4mplkf8+IEiM1hwcLY0Gd6aeNU7
TuEcynVXMENsELE4i8gFeD0FK8LQ6iw9A0Yr19UHMQT8HZZvG27eZyJ2GbQK
zeHv1WxdK4TcnF6HEz+u1aBh8UOvfJmbe3Bw0zucCIqyqxn7D/9okPwHese5
CsaWESU+TFxWAIrJlcx8gpVeoU7LKfVjlhPGXNvIrkTYcXQGHDcNEfeQgIYJ
jXFQGeNDztOQ9uPqxGp6IRAbEfjwBaaRfJ2FGgfa/ASQHvbDlFbu4NYIOUxB
EN3ZJubKecNOM0jGBushf3gX8ne5677palLF0RoKGvN2+1AkM0c7feNKS8lG
uswyHEepI0ISV1PvocTCO7JIV32xykuI91nbXN7njNhKPsOzB/oiDXQJkxcG
aaYeWbxSdShVxlQvcYzLDEnPWBh0/8bcbOIZw3Z9KUw/0SoSC/AobVRcyHMd
dSIaInKyE7OAg2iqpXlNajBKqprieicC7dym3UiE+VI0H9+GzpsebhBwDxLh
VnYumGwvHtMhdHIdhXWZv4JhfUwn8ZGud447kTtf7wG6i6SyEcC7F/SNN+O8
yGfGUDZXr/HLzGolcELECi2EMwbKm7Y5HqoLOG9gxRblDiXFaseuah3KMj0D
1ZADOq3fSM2jaO36qTdgDB8puPlJCrT1F5+8e4/sB3tAOr+x51IrJ1zPiRBR
xL8xdDmMIiSKFYtUMSFZiwEK/N6N8EcrOyblh4Q587BpYn2Y2e61JpcZe9qT
Wdktjem6N1/7vhXIpograSNm9C5w4EO7iIduRyHY7O4Ls0SFprYc0fwBnn5b
0cguNp7XPMuxA900GiK4w+48oPUFA8T5LYabPhh2qP4gqBbTRcmDCBuZ1PgC
WJ5kCEnqAoJ9MkRwbfq2vcraXIO6haOE7jRbHEdUkl7msGB0RsInGpuv0347
XSJ2FKiZBm9pn4Efg1CYqrvXHrCmK7h6OWOfDI3IMH2iORcAoYJDBjhH14+p
wr/urfn8IZV7R63xAWWgt91BVoM11/Kan2nSK2qmlmpF+pDQp4xDTMuHITNN
LYPUx3cmoH/myM4QAmOZuh1PT48yr67t+OI+zTUafunIjrBJZPxSpdHCx1jJ
LK6Int2tQ+wye616HiK1r67P9ZOeHGL5vsMPSd1m+cpsviAlWRSLc8nFlXbi
cTukBzxZvykEdUdtTeFzTdHd642klg3bbOWgCF/LJLXWHgx4V1ocUKhIL2No
x4kVQrKDVEFmxkRd+DRWlFHE1Gv70bDAFdPUTldNcMnmR517jbtYimg26CT9
sOd20B4rSjLa64eh7OyjaQTvb/we6aiZSZ4ziX/svhDZ1jjS428Eq2MTEOUf
7DP7NRgbAfwyRATiN/geAf5fGAMFlfTIvJRpcES5wtKvuqmCe2kCYfMCqyIz
Qy1QVGkQGvszjmSgAhS8fZTPwbGvc/gWOcB45j8/RVxoYtVwH7dm6rY8Lx9+
8lJtDk5VxnnpFcjcjVVj3yR3trC8pPcLbbi7RZtKHUCojKaNV2+7CIRQgNqp
8vpGOb8VxOVO4bFKu/+DCX1VFH6TJ+igK2Gjf0nb9Y1PEZ5MUC93ZVN7CPh4
HW8R6IpYAipFCWnkC+C+UnRaYWh5CnDxZw7V5L2i0D58vMP7wnTgTQ4wkDFK
mh98bSh+FXHq+ca6pjLgrca9UzHy1sQW7S+kK6Wg5dJxnWNYsoMUDoS0ikQ6
iprGEUXEvokWea9MP5Em3lzTurlJLC0e3HBHaikY/o/nQ0pzl+xiYo534kgH
1u/pt/F/RNGvjXBMrslyvJmokKpcs7D8fx3o6FpoDw9lhtMv/mh0kFapNbNg
NRRi0muOVuGNX/AD/H78t9iagAkGDVi0Bg/xWkfR406x7HrXWKmWdHq+bhX1
cG6VT/GwZfUKBbnRz9E6KH8AXzks0HJJ23GNC17gQCoOPQ2GX55KL6uiJz1m
f9vS4wYLUG9TZjZQSx9+ORl6poPUSSv5iHHvIaboO8V6MJjIMGMhYNRFYv+t
QQ/daNYCd4HK4H1U6E5+mppZjgnRSkBRcd8lbCYBeg2lb469oNtRCUpi+7O2
u5O0k/ca+D6P0R95W7QLrmq8CH4tg5zh4Coax25zG+nHE2VaZZBQVY7CcdOZ
FD647Bh5djonMAvUBarbqvzfh0prMrzXsshQcncWs7aXmwZTtpTVWMDOuB6s
A0DuQ5RYa6Zxum+Fp3oyLcv7JFKG7E+q1uFrwLeJYPZ+P9M0Nk9D+sdzAse2
rjAOboroNvEvvWZ7QJY60QZoQGW70axFKSxuGAjhhl8/MyW/qG+SPA9YqFtO
xlcvdeVYUvdDXAT0ijeBV8UGMOvSWQZSi3ylq1kcdn8Kgu0jxVLFkRACQlHX
xVaobtPwbr5tGWmsVOhZxfKq1eH5t+AIPWRd/XKE51mveLiCzp+8nbUTMcXC
adyiZmay3Y97VS8V2rp82uWuuKWGPXDhH/QpiFnHtYzUaZYJSvbIUUO9Vm+2
KuXWpGL8u9FvdglvEDb1ccAo7XY2ub6PQAV0TvdlRRK49MU4dvcwRy2hsK51
menuI9m0AY5j5ASAYw+L5/ERSoeG+zyWjY2QgOss+cakg82k1PMZM85mkVqq
92uO5Jg02YywReGHZPO+xAoe9oPAG+j6qjPiVpSWWvAnltt1xxIS/FdZhlxG
ztrd51/x8pGy5dDEdXUsw+E/9YUClG7G+A6o6DW/g5tW9y0FGzHMJYU928zD
RIdJj/1t+SIIiJ0W8DQSL0K8InbwXLnFpO7QWL96s0UXP27zUaNdy2lxnOZd
VZnlqGtQwyFWZPo6qABlwWWnYQtKxl7t04TmusIopbRgh1W2dOetAoeKc8JM
tnR7OuWilUwJI3NGVhc80uBrKKfyv2+CvXE+YUopMQyLALHTughqi1ukFCw/
Vjj3sOnKgj4q0AGT/fJoO08mRNsMl2xKjinl0dSs4PQLzYHnc9BqW+Q16mnz
Tfi9Z8CAhRGaaD0E9KUuWcPinbPpt/lUitNcxeAUO0dg/8ZCa4VWCV32GMF0
EsXBt3LCQVWCH8TSbbuGjUHxEQKKWHtpFcEIwtH+sz7SnKeuUClrfNxJozqF
wZmWHalum95z4CWlaQ68oJKiwpcP9I1xRW7SCPoCSombbwR5vx033xxUqlLv
vYn/u2PgGabykOEcG6UIg/zy8NfB6W+WNav+qJVtQg93rlWYjWoBD5nr16TI
BfQmXKfJUgd7kWGSHc0iy9BJSsV8UooE8MM9sAdAsp+f8C3oSXIjsuwb0fD7
uB5gMHDZUs7zPFeM1ldB4Ih9uBtq1V3hzordIW9RAhGxEz8l8ly8GY9qVkNW
jiYf3bcJfSo+5y7qhNdr6yM7UPA4/Qm8OqiGgHEXCOA/LBQfMc8OXKWuWvzU
ftgteuto4RBi4Qo2nZy+QOE9F8QgJqgc7dKoJCT9VOamo8Dr/jnx/rGhhi6h
URLU2xjPLW7zGnx4lF4oVfk7sZOYHngb/STdGNLDqNAFxs3INpGrMCSU22KG
svMB8HCZZCIW+3dma7crqBOHFrYcC12mmX8aVYnlgD4JXbJ5lsflnXo0cAOY
x0/tRbMiCPdRbswmxhfM5HVl0krlc/ky3wyCjtiihS0K+BsbMOJcGTehk10y
hasDwxTbrOX+NL4cVHH8jUC1tkhxi2NHRDklJApsQpDe8/Q0jQuQ4afNa70+
uTt6xmDiXZxISpMk9t3eHUApAKD/ubxfrgv+n+8K92IAcIgTrvW7VQWcWiQh
swX9txKN9EPQcTxixJwA+d2+4R4rVtdPPqoFUAvAI9mSvUWXB1RUYB0gBWMA
95Tu/4p1kSX9cMiKoJdou862jZqgniiVDfSYMW9GRx0zPF5dPpm8o1zzGy+V
uAOSAelpc2053mQdFGSqWP90/1UO8lTlZomIvpC3Y5qY15cKGgXycBBwuDOb
AoyUBKzJt11cSKG9KBL48QvIRKyUW87R78tRJJL9lM24mCGg1+mqtR+c5Y2O
ETobA3NOQav01pVQ5lbgvS7SAVWdwN/yGWHpC/uMGL+9W+fApR8kOV1lKuu3
0SS04sVKTmOxk56MFMv8+uvL6T0I90Kc/cnQ8FXwzOwO+5ZvcJKM9JwnaIv5
6CW4oAR2ONThJYKXdYSuAJPTpnj8nJeV2ql4b7B8wpJ1O4MV3inYk3LzQeS6
8gB+jsISp1eigp3BhWzrdLPrvYaXSNDd6ds9F2eM5nGmT/UFXZHku4u5+TYg
m7CKyJ4Ou+NwTn14MsFeh6H3z/XYN5dyrfC63/5BXG5R1H5+REx+mCFipXHs
3dYyKk5+X9YfdNT3q3fqtHRMKOXB9/0iaJ/362JtjnDTNrOnliiaWW+3QXTh
M0LmQLykNcuZhb8ez3h2YadGDkghv9kYgfWUE4fhn2JAN1a0EVdU7s4v8nvy
FuU+JPsu8bTgERhIcl3kqIUBAxko9tAFw3xRXsM1wuUjPaWbWHDn1IQFqVAi
ZPT45gk6Uq4nxUK9fvQtaTeUf+TxHvRIcz0hqXT+2CY/K2n5/SdjvxOBvANf
Nh4+XhuzNBu4IKsSF8thN6Yxcx/IBBxch+uGYkjogy8io98Ih2bKWCCQ101w
YXDVAIChnPXLEna+5W+wNj1RDReuzjuBJx0vCLjgeXab+VZozFOEx+FwKLi4
MZC41WBz/YXw2tmWenl5d+OGje9ZGuyWRsWCZAoQ9X+kTi0+z5gJ0JTG/oK5
422uTysFCD7RsPcyjTlZiDs5/WT32GQEbOteaHLMy1OJto8kND5Lr7VzoN+b
1YGDhthrVatu+u7Pww8qpoEgKnw63+RGLul/ctA5nmhsuaCm5nAWKQpe29Ex
9TXhJUj3KzsJpwYX9dF432+C+LIFJIyicBndMQqvuLl8PgCdDf1rfLywjH1e
P5wqTwTrngFgjoWMZqoBIuq0777KCAj1CjYXRbOVtGxSMi03GVc8kQLHTLBe
FIv311UobN/O83W+Z/whskvK0A7o0PaGEzCuORXcf3h61hcagk/ydl2zHj58
urwGDqLWFVUgmZh0q0Af+Y0Nv4jKk+inVVRS/ALHz4vZeP0Jq3PgeZjvvmQ6
3vGZ2x/uZjNSYVMuf5IfON9VB1EeU/aWEl73T/z7WiPcmpDwJdZMbZR75yuC
943sA/1l8lWWeZdiJvsaKLuqDa4zt0/25x4nGbyl0J3r79WKBvSziEHOHuLG
9IiOB0ku18dDhpwq8Ijiln+RN6IMAEx4z8KqbACbFxbCQz05raTahoMi74HS
fu85eB1gmJx+rXoB73qbGH9YiY6ip4Xps8HQsOZ/attVUx+oyjZyXeEs+VUB
2oLMIyxW0avCpswcUC8Q7VhfppVRRnckWdTX9uuh/eK/QFxLyk1ItA+X8Onm
OceLc/qWleKxFxJNj+yTnBpGHY7J0B/JKFdv1nZDjekjsUIeVTy/EyosmoBo
Qn8RR521ytu8ZkhFI6XEwaY80Z9oqwrmNypeE/Yb/FPLbZW0oJTxo4Hdn56S
csfwTmoYVJ1633OA9rhiKNYCjdOLEhYYFnnDUqvZvzlYpMczZzsLJWe6GG1L
Rzz1Sq7aYOA+oImwMFyexVes1//WPilXVbaTVkuKDvi8o4lR16F/4hduyPzj
/vkEUmXcXi4Z+77zV9tWgrTi9h7vTK36z2F/A28xKlZhglaGwVY8HLq5k1BL
o2o5GGsndJkEg4Xt7M31DUjjc9PiVtHOJ557Q5I8+QNhcI6ra5w85NqbIpec
iwLRPWDZFxNC8EVsIFtHx/91IGuOrm0L0LyQk3yGiGYsj4QiECoqfLzpr3vv
Eq4vo6ptYM5rvM3G/bRdbhNcPwirY9ra2cEibBSNQ0g4RrPF79ovKLCjzisl
HW53qO5jjwJiaOzSTrJTmAc098ASO8lVLbJynvJhr5wD1YV9a+e8qtBFUgLf
bFWcyYtjzs/PCfYAtFfa5D8WLhPRISsGHoX7xOQCCupx1pVbExIciRL5ucnd
1jZA+dFvj4NbRx0hZesWlb+pRTeUZYhOKFNRDn5gprBaiA0k0Q2kX/c1YBc+
qwkgKTnRiL9fD5V6Y998VJ4jM69dcaqisGJN1uk/HuAG3N9RclZbK+WMicSr
r0f/6wWDH1Vh5KVSza5Dsmz909MhqAQTE0h+0ZOcPceELFwtlulsyOdLhofD
W21SBRljDTJ+QaVY26H8ZgGV9TZxPhytLNQ1vXjtvPKXl0B2fpvB0/yQtB4t
PimoMyLV0QtUlHqtJa8OCma4USsqpfsCtLIHwC6GADAzPblcxE+2Ydr4kKE2
gfTpyMBlz3GEIpqyZOH+bwS2LSC3Mei4MnXUkTyYOSovCOw51Q8Z/ps43ZPr
PIoR+wdyuqoTthKQR0/QmmVunPR9DIjkODvJPTBUWmhdHkBRwll8/KD5g4iJ
ic1whBCtqEaPI8xYAtbt1/r2LDvLoP/LVfsHcrT2AIERmioyKMz/96mLyEwc
g948xeW5e0cubkf3E36LmN3MnYWbPTlMt6ktW10Odib25bSUU3RFDPjdfZpN
/hLC3dmm9WTlxKu+OO3yM13ebdu2D2JFEDoVgnkPkBVrde1bwIKNVgM9TGuW
hk0KIy3YfGTjFrD/JGtTkQsIsgW+dAvOOgdL6ZmEJ22oUAhtmo7LJXrYugY+
GGkgPgHMAOY5GmW/Do8hmVshQJfLKwK9LXFMVzup3GmC+eWpuNVFZC+Kj4rr
BqjO47JVXPwqMXqWGzmBqlm5PQC1qJxtlUlcRIQpjzgx5jOEd6jE6Uuj/Rzf
DIljPv3lU9Z+cauf9RLDL3UZtIJ6dHahFmGm/jGcirvcTkSezKgxJc9sMa+I
YimzbXGn0S5Ui3tDrjtG+ndbveNk4TD4iBrIiRNln3Yf61nOa0Af9ye6lmiX
D7sruEKcMS5YXWWP3DYV9B8p6JNCRvzakIjQ3qMxRzatK0oFSDvhv5ezhhdT
HNXkNMoP7mUWei4vIchdYXPyWnfdgLCDq4LZT2sBOO+w6eOTowBhxMKJnChT
3awWP6nbgz7J/US8GmZkWcvo+osYm26BQ4aBoax1bOcPqQ7J7FAXptqFVx7m
cmkSfc4BuypV//qCEqmOqYxOVVGX2Zja1W12sQYNdokx2D2XRjW/dfqnNNz0
nmiZG+wtRy07Ebaqf2B49wRhzYdOvO93ElRqr46AUCSGwgfqZpcX6FhwGR7T
rpyae7AwIZzn7Q2788QpTItMi/6PzfhA3JfWiUx+6rX6Sxrwn/d46QKYW3RV
AT0rdJAHF9tVW/eqLwz1InPjGuihy0I+uh1qD0z5R68poqK3u+5KI2rWXXqg
A59DPGFxThe/2ADichkX3FHvCf81kpwxG0yH78amTYS6Bxvxsz88kOJlJYTI
TsrSJq24mvJdFpOGNzKC3ng7tq3OlDapi4mwpniopd0AXNG3a31FRSARpRy6
fTyOjD7SBPKDdz8P+40opHfuFTkst6jv+rRy+qYOc9r70y+YfVm3bpmyQhIi
uBt9C4AP1t65ZARMcLxKXdmmA1xKJAQ/wnfZySQjzy6KmhcWZFo3qOe2XrD1
9gD8AeivAyQpbUWpQ7Odxiel5CQeV2gIGbk7j8HkaIyBNeF4SQA6U55a1TdP
/4BWfeiEbdE7VXb4Nw5yufxQjGTzR2V91lJ4LJV2tV73JMZxdKBBJSxcz2fe
v+sn88t+HxVJyAyjr0CqeFD0PBTDAzXCJM2GITV/PhrXtRCgC5N0M3/YFUCW
hdaXX620mVO76udfZLYfkjJ8BdBhf3PM3FuoJ/3AblWLnAsFsL9vX0XEjd/W
LV1smxarMNp0F54ESiQmln8auFRuPAdqdsC25TKeoXMYroRsZ5oGMlZgP5in
NnC/88B0tRjPhbZ6QRhf1Eehapsc7oYZfGhZCV7jRVFsZyiGq6ikEv2JOexs
D4OMFpwgt61LJJxqONFQ6C0UotY8elvoiCKLwH+vCZuT9+pxAkaprSSVW93+
7D5f0LuFZc7OW/ml6CE5eOZMEjpdKYsslNbad2Jb7CmY/ms6eE7+dAchhQ2w
9P3VwfiknP6776YIgkiJ2vfhwLKeeW1UksPjWlFumKud4cniOq95KbT6gNJ6
jYrVJJ2FUnKbB/KrCYStWnsqvOs4jY4eT4lYo4PbzSxU0Uj4gA/55nm/i4SR
M6GZo7bQyag0K9Pjx6e+3bPTrCUOb4BWXfHbytODYjbbhP8Es8x4q3rzappn
I2Ev+pkI4pX6XuVdh/y42Q94b00ByiNN33sT+66Yeeh9Qy8+KzQXucf63NNk
WsqMyc6V6RLh9/AtxMRQ23DYxNSh0TyCQkhfRD03/M+XmM9zD19r09rZ2zsZ
NlZeYiS95Y6V5JDAt6m3W5sOxmpMfc3rg6uSEYXS+O4ph8XWNRbXvtzEV7qX
sOpCMlDE+f1cNut8COLQtZbWqxSYmAp4St/QiuwY/DmtQz9YCWKfdmJmNDzF
oVTSE86DgSR/ApgywSqx1clhIoQxkUoCPvlnSVdCvmc/LC7599BsKRbSDsx6
QBt/zEDM5CfiZssu3QaRbwx5tZhvwp+M0Op8M8fPo1KMTtfbUI0gU4bIMm1F
BJrFhQLmqkkWlRwdwYN6CS6Rkw2mLileMAsHPXpz6dcee/qg4K/j4X6nN0YM
eSURKZ35tT11XQrjZWwRs/sLIzTbjEKdeKELtLuSx/5hD1CuFc5XVxF8tGzD
T2kdiu/YdzzmGpiqPlSM0VIGEQCoTFmQnp2ZbAMIi81CgckaZbcLwYk4DY0V
C6wtkP2nkOmeuP3yd+X5cTQ7l3Y924+ryx9Ms7AoliNai3vxax8fQ99MrTwq
qX4Q4xw4Cdl6CIx4SsPsQ+ujA8Rc52saK6tM2SeqwML8Sot4UAGlXfeNzz0i
97W5SaD51+13DoUKQ94AnbcT6+0eO8rWPjAse0IIPVHPF5pG5H2A7K07Di5p
FqWI5K6VdqsgSt+faHgA3NN0F01F6bQab/1+j2mpKKDrZI9xW5ntyNuHXFiF
6FW5gMJSCmHxymscGFEeOz78s7lxbDDW3AEsC1QlLHA+/E6L7z+0CvyrNYXs
Bvw9nwGrF2X+dS+ZXo/vYCmv0v/rrkEzn95JmmpO/YZfo8+ydWYV4WIi0JCD
PhU0kZXRqTHXFCIwk2XSvYXIMLaEjjlSycgePN90JaxDGQJWnSy6u3+2MrCC
nw7S9MkeTRSCdQveJYZyIbS7URsDZzobb8yjlK+DHJLzkquN9j5QmSxNxi0/
+xJazpe4tCmRwhJUfdShDsqar8jy2AUxEx9HZC8STBIzCzuZDox0jS174gGs
1JPb1BxP/yuoJFcvomO/G0/PnXRDM7jIFLjGVKcqROeZSQwpbpYLNYQauinA
42YM4kEr5CsbWy4/rdWy/lWblbPO4COiZdZCbVe02wD7ODuAN9P65KjWQey0
98FHUX9Kotx0jsrPeH1t9yvAD3qNcmo8f2kkcQHJToRSMDHp2YOKBfN7vAeO
KH0YpYmB3JydPw2f+l6uMdxeSp5ULoDcwDm6ZvVtaKhak+ek3YGAF3H4v3nP
dQq/r7O5WeOYgrxfAk8zlBGVgogYCviySFq5e/meKHoCrLF/gvRxLO0kNg4E
QbdUjg9izVc8VWMGb67+4YNS1a05ztVtZ1maGtHDBngb/Xy8M9+cpJf1dI8E
YnNIZ2EstoQJRgRkvxSuzBlUbXsZ1TBh97HyptD3E7C0Vi4O674BCZaYLH4y
REXsVKrMskopvF1kRNivGPixqTp63zxU9YiNXamXo7FZZIEfwrBA+ib/2/7h
dwQuevha0DkmMjlhqe4BbNSzLBvaxOJEDYgq/yY+t6fxNGhnrY/GIvZJ7Xpz
CJJOuS1PCC4MHacwfLRISdALAwken31fIPfGp5sZ6OwKIBbZbp81/VvzjROP
3Vn3S70Ay7SzPvNGOIrjvDdyBTjlqgoc/J2S/trTBElkTbyWog1BE5HmI3PZ
d8DBENKq14gH8aeILlHqGt8JjVccaEACPeXhtbbCSSKbuL0pfbW8QSxj+BK2
w4j9GE9CAmau1p7N4qV8wJ7oQ0jZAjcZhfuR4nBe7/OfzAsXlxaVCLu0dgwE
3Qk7gcnYK8dxmh8XQD6TaF2Z4dqpuvSFntS2wfLwB2BAzwNVJr2u/LP8QVSK
uMR+We1w6f114tifFvfRKyqgmBd8+YD1uMf14PgSM4rf7TqS7XOp3Dx1Wxbt
JzFDFXc0Pdhpti8NWpx5tYRofb3A8X4gA6c7zkwf4SSe8k1RrLnngMkJZ/P3
irS/x9GZ0aiipg3qlGhwfvViO0AQk2kU7DIsSRsiHKFKgPLI3V6lK5jIeUq1
Z7K2deEi+up5nH0vTJdNbN43yI1pe/R4YpXJlRvhxiWQsV2WqnhkcnpylWQM
l0+bZhf+tOfkWnm6Txgr/J0vkLW2xa54SNYcoT4tdiJChh5eNUIELbJ86ybc
zwkdNWYrH6ia9fQhlmVCg/ir95hwWWWW3UeXipr7eXjUoVZqFhOezihkLMOn
v/Os+CDxoogT8gGclIx8ERUd5QivLt+p7ALF9nLnNTY0cn+kzz+jFwC8hA3v
vmU+vcZe6IgQznkCrS4GZBHkUbX/zmbFQBXugsywRwg2jjae+Ee5GO7xLS6/
E/JngdzJc3796pak3DZ6UwagY3nMbO+A4Plpf8WgvFZH6F8uCv66eC/evoIF
vRTCatUwBM6V8XDAggc2m43jRAA4RluY5qtyBnBxFADEAagg6V4avVuD3rJW
XNLWY+hCzorPPYzJbeQJZqqG93F8brl+0w33r+UKFsCzMI8dD1wBDhc2ztq5
lf0rXkLiEJdF2Y9v5zvByma6ulmV6M6W6oEPyXQSD54U0Jmv3hN3XV+qP8fA
PRU7c3TP+tI/d0aM4QY/Hr+CGDAHwXZdKjbqxy7jtn/qzsYmw46YYaTsMi3D
1EPz7Mr2ixMwsjap6TjQO4TqWYLxntakdLtTvkj2VFrFKKVZSXVR3kJUhGhk
0t12iut5sL0EVjbSMKAPpntGJueJ04urx0JmpdUFubVuLvN7NrknQtukRcq/
4JbPJY6W8bmS70MOe2D91Kb8CQyF0t6ClDnGvrcTl14T6FqE63ud55rixOtL
kQCUtpVkvjUCDAh6SwUBkq4rlDWbamJnFCg1Y8K+xXDeCh1p8xu3bHh6A+ZU
nIOjMV18S4rHyO3lRoJkWDiwQtmZYrfFPTejuo+h+g8OJu72n2mYe8quQH1q
+h2eCBTyLBvLYQbm3dXFH19ZIyTmxKztD4yLseGLxEbuJ7XQNKtuk6/IFua6
oxLL9PIraVMV04q54g0wugxxTfdVlon3Pq7R9fK3Ka1sieo002AbYaqi0N5z
45sYQET1AHbYFBOMVFUM2JB9qZSM23bJNg7x7Jjnn6HzObk1i/iBhOSKmb7V
gI8FeNovfD8cYKNJ725VCp9HojRMYttG4D9CunXA8GsLosaYJjBOE+xJbAw/
6OBzWYYsf/KsBumg2PKmzdrSuQXJs2MYBTpW6gZJOCbRybeizwVDwxJ+wu6Z
wAJE4dy/6demewhq0Q6b0BgImH3vtgLwjXzX8SDkPL+bs1KT1SGGISes5MbW
N3o5Chdjwl/6YtR6ceKWn0w+YVfLrIPT4tYqYiEvgd5wj4Aynhs3a++NHcUY
uB6gy3dnR89ipvkaYn79RfSIpocKUD09QQrx1mAWVEal3v0M0kBCDdI82hzL
HbY1RsmqsFMrFfmo5/jb7JDXNm5mKqDI6UrxCC6/7eL6Qow40u4efaq3DUgL
L9GBfo1loxwOE+FmSfZXn/DVufwOAUbI9fFulloXZD75ZYbCJex5KnEj+t+I
OKS5gsCcQ8giuv2BnJfp8823hzpKFOTPwagNHJirQQKz8mYHX+mI5SZINLrA
kcH5P2mh72FZKNp7DKGsEL2LWfo61jySlpfG7Womdn89Nt6zN90ZtdS6RMGA
+qLMw054JdD25t574yFxk5Sws7fyVJ0gX7o0imCLbE0QLDTWd55bwP+f7rql
HRGhG2a6tZ5VmzbLfcq8UdS5fRngYEULTZfUJLMhmlvRsNlKEGkiKSSWuwUz
Czu7wmYOiuZC9N/KZMLzgaEvL7J77eVi+D08fuZFyZQNH+X2ATPck70w6wOc
zwKo7gnu8XFJBhKOdZbz1WNib4LY53hi45glEIA7h1WnuUaX2rSNsLC/YjNa
nCI5Mz+zYzoMw3d/RvoRnoXAttP87rCemkBs6lWR6hLSLYU5SnzLkyL8+uQe
NjR+cgeMu3xNuy9G13UWawR5Sffx8QouaUhV+LOkyPmrHNZVOaZVKpy8CUJT
SqGIS8JnouWe7UqFjT64aX8p2ONcIVpGdOoZkOKXtEgWXQ9t4T40MmLIQTar
N5Dh9cL2JZuDOXo3DD7JGmL0KsgzyylMPu3jRX/mw0R3irHL0vtlGUJ1DAwD
LFMtdjpjV44T7bLzEZGX08RRXjTKaNjJvw4w3oqvb9ihYCpL6bmskAAJ9K9T
uMaGj7h9owTwgAT9lmFaacBJhIgkGr4QKC09LEnOJCmMX073iYErR4Z01ipz
4MjcxpOAzFW7Z1Ia/0Pc/uJemQ5ZE63jG4whY8Xrte3RlU+9lWyJlQa5llQj
549b2O2YWphDOo88gDl7WTda3Xa4DpBNJ7fDkMlRhH8Rt1+wXN3b8B6x1cBl
PNFPaMf+0NVUmMvrgKf8xTWNNWWt49IEIPYiIKq09a/MEW4p8XpnC/dpkeob
E7dyLYFXn9yOljmARtUOVNzTshPR6DISYn45TiI09TjYJy6xA7VNOjt1+sSx
f9rcFJ3arV+CUO4vOomyzLhfmAhc8nw/0ex0QMjPbaHNUrLF+0kpAcgPluwO
ibKsrAg1QFyksoERPH6ZzNz+LGggS31JziyTM8M8R9ml/Is+qQb4aOK3KDLS
EZy4A3lQ6Z+JqKbT4b/fhXeTwKw/p51mcN0JrYnj1VhY8pZYaT1fZyYmuIIl
DHZ83utCxsLAoml7hbpL/07n/32VywIxfDJOS0SiiX/KbwomYnUABMvOtc7E
70yrHX9rcutiJUlJ+xYpeYtzLa9SzImTCWOp9ksu0aJP0jlMC9Cto+GsW6Mb
utpDoeGU5P7PrYeJcmas+dZls9DatxAOjJZNowo3cPNcse2wr9NFYCZClkzm
VBeZ7f+1s4TvvQRh6KBTx28ofyvWIwpKN+ZhFIuNH9OhP/TSycRBs2V1ZNf6
lfJ2USDiPCzj7+pvIMhvdFmwfCcr3uiIecUREtV78nhWo7oq05+4nggduNkH
Js6dc7mqAl6tAA+iW8vnshNI7Nn42M+RauyhYq1I9x3OwuAEUSN/bru8Qo2Z
pHgSYPlEEZbfKa7rcsbp9v/2qGilbV7UzqDIVlR9NFsxU64RTrEOSdnXz88e
YwwouVrTHa5QLoI7P+oNZ6Cmi1YOH9jdD57BLs+eCGHx8Ue80TJE7wVKff8o
k3ete27MuIwKNldAu7rmGg9HfP6DnehsVZky3zDOfQzG4+iCjDjET3Z1f44n
c+ZXaDm4isjWZksY/vDo9eAg6KMmcHmRyMVCiiujzgVpfUiM4TkCijo6kMjj
Pyl2ITLx7yPASlP/rwIPWWwfHQFjy3uJgeW1TEYQCYE5ANiGKQsn02oEsqaK
0FY3ipGhJMMIR2lFim+s05bvI2XvGgbLC0lHSTYk99PqOh9noC0rfhZAld9x
H7vq6Ycu8UjDvfqZERv4WA7Gb8GxZIin/k8AqQCQNjzSOtCVesnPct5MTo3y
PP8oP/z6XCuI2TiSkvzjoUukNh1ERiQUw11V6j07BrIXWEJNK7F05NIIPo1k
atvdfnpwHFoxCZH9xiI1qSzHPhAC5DfeUYJhSg/zLxYL8ZsmdkSoAv0/o1n7
u+WMlezpfpQdIIjKE+9VI2yn2+8wGKCBRiMIBEnria1p2GE/YsScXTGt+228
xjwazOwVSVkAiHfCZs++Ac2DT25scmv/c9Ft8WlGBznwJv+hhUsj8tqDNgyy
XF9tNiMqnpInCpRqwGj4Rr7e4KgXouSZxlouJMdDuwdn0abB4pWGtnf/bEWa
AeYaWfv1t6MS01xPzdt1KMGXx6Qpo3/ySkiwYU7q91HJGyvfnVoqj2u5uVTJ
tBUNkFC7pE/jY4QD+CEWpD25DQpuVdQ/p3pej2/OUwQhStrCF+obWWTKHxjO
Al/+7iWFIEv1Hnj/eAxEozSBMwReVUrSH0AaBU43QrPg8ONLOmCV7ts2WcL6
vcguRSrPhbLrtGqPJeQETIbJnSEsCyzr/Ll6SuxneYZLEfIpZHktR3a9WmxI
xiYSaJsYOLqcEwpKwd+wK+br84hzOWEHLOGFtF8k6M1QSgb6ktdDStWIm72T
wVn0kvqdl6LCrpzzYCpl1Z9+v4xdowe0VhmCAZUy6v+crjIi0v2ZSSbTEpY9
8vZWXVdy9dmbROUtxetYCAo52+0g0Bhzv9TxzvL987Xn/dUo2r6gqMaFswrX
i5EN+z0fakbBA/5CokdBlGcyTxHWPO/BLWHplAxXVeRcpivzlt059C6xMW65
q8e9qCOKfXSMsEhMZiuSmq9FOOCX/UaKOeigzGdTggNBKbfva64ojy7GoUP4
VU7k63KKWJFotPqhQ3fqH91EVxc4kEgf2WqHM0rFw9ZtXIGSZLW+1QlpuzmY
Z1ZhxfBcstx0OOzI5sUHrrr7iAjsdAu6z1Ris/X7qHUH1lAjtGa3gGT3386u
fn7coAuK+xRAQTvSH0p0v99khrIDejxuNpr5+dLVdhd9AZLzjkMIp/XvQIVA
4Pjp+H4zeOH5+OYjGp2plIZ2/O6qkIiPkmuUQq+Syw2zp0bKCkNN1GYtlzaW
rnWyseyaPmIeAxBxvrYKZ810EA1rAFRKMkS9R6BgSjot1AHlZPQcGBm+tSPG
rBkP1tGWkR8GkXaSPbAr6l8dEjKbq7WOpjgwO9XywqAsQS2vYgy1XDtab2HU
wiMoBzslFYYXICS0SdBMfGa7UDTL5OCTMdQjIPACktXFFjIqpLHmKQ4DrYN7
5U7N3sO6LP95bB+ghEVcL/2T6suwRuXKlDgc3eiceOTD926x0whXEhZdSJIS
/BorTzXfAprTqpkyKnDKE1UKb+ixk9T9Wu35QPgExD+VpuV08bEHpwHox57X
zgo9BOfLoMhWzXRRgb6KqxDnGtZtFRsNHW4MxcTLFRy4ClA0RI85waOIe7gP
hdVKqk5ExkNxqgQtmxY3EMC17Du23wryKPHokHxCJnHok7PkWpjOubYrqOsI
TAH8+NvTUdWN9pMVDjSZHRlB6E0tmb0zFh0uMcSQQTLm3JlX6IFoeLt+AH9/
ZxL1vtHoIxLUZ/2ZJKCczn5OuQqCu3Y9wBUYT3aDgbvvkjgHQRI8EaGzwyaG
PHvPbSHU/y/3CAsjzBJ1AMQILyFRkfjQxF9yktQ/xIN0GOFouMS27VKF7Iou
L6LthvDg1AtIyBIx7e0QHwYId1+/0hZznMJCcppLYfH/jwOgHhvUMZyEk5CY
YceSxcLSDK+dkpBCeKtxiIHc9RWtVHKDI6ThRl7jMhJBLvdH0gLhylwjI3uj
kWnBO+yKNxXO77IfAuoHCmLoWlDmtmwUIyOB8s1qgw+PnomOUXAd35UXsk2s
oLyqc839/QXWYcZCBCnOXB+7XCah/u88AvMAz0sFGzLegwPR4/6YC2FQKFsk
yu5H706mTmlQN6p3vq8AcKBGjr26Fhc/DJ/+fJ/n54m2xcwbs+sd5AZCqhxN
Azg2xIC4nW5p7u9S1EbSnUCvcerKrVwDU4c1k1tnNrY3R9rRvvEqOnQlQRzo
+OMSWkF6ioCJ5mGHPLj3osX4vh/52Qs/jZwJt5WJDXm9DoR8IiH+GOOZzOnC
OB/6jDBHMzi/SbsyBWrASDFlZ1nQTqEsVUGIlbssZZIg1U9w4tLXVw4ksNNf
au5PVhdc+eMcwnNz6rMd2i0Vihv8AGxniySxGJiUsa5QvVqLoFZNSN6FVQJq
HEIFwOp/XxcWKiE38g2I7oZw29phQR57IoZWwQFPijFDYyu5Uh5bcalA/jTu
kyKFW1u7hLfoIR8xAoHHI8jebe8hVu6BV22JKavCcj4qfQZ5U91znt1xNJxx
3aXgzwcnt/za8ExT/3HMWiGYtHQ6ioBZfTnZmBm86QcSJawgTk6VqbbTqnr2
P0n79GX50oKXUomIpu4xyzH81kPAqT6tLlG7+5Bs+l3FVWwKhLgMs9t5FKx8
EatdE/yzvtz/DbK6oK5rxUEuL/s1ItV5TJie1qfFS8S+mU8qO4XIUMxbOx1s
OtyW+tNakl45ka/wVD5OUlc6z6vC+9VcJlUUAmd82mTH9YTqPXvjUQth59CA
Bugklwzo4qCoqHIp1/ahF8idnJ+1QxjI/NVvpQA+YyECcqiLE2v/H33wN+ip
eB2QGkchAJ/INxtyIGz00n4vmgH/+QG16lBQWsjIjwCeMoLhIdwmoAiQtXNv
XRn3gDPPcxThn5eXR919zYihOOhedApWzfD9LceHAEr6J8742IJ7KpxhtVtF
PgkfyOjMgKe6CNjAVlc9nQTXqhuj9Uu2VqPTwP6qhYuZrLBDq1KR1bnRhaAi
RayNc6lRkcA41+5H9Edn2w6v7VdaVWzUNlva0mtAYjFQQKKTcrgXBo+eemHI
sBGM2e+oBkDvcLeSsx4s6YEY5JY1PLPlpMzg/+DlEr/ZNEhg2ga4wIueX62Z
ei3SiGrADMe9IvwrRzyFJhB6Rt1cdtzNVS1FIf14g1VdsnjmDR+aCwgC4iuN
8KNeecPjQVmhZ8/o1W/Dd8B/n4rcZXZpD2B6eKm5QDXvK4RqGtw9+MEvGAJt
TFBnA2nbkW8CwGFpqK/w2qkXDGYa4ZqLcSpOWsOhmL0tTWqaO6DbCVrYXPjv
NTGNFSx2Y/EZew/KZdoz4pgDlKlNFboZopuHU9aFpxHYqMsQ+yCXSZQEJ2zD
xCbpZAZJ6C4YVD5asWVUsBuIIup7IWVLGGW+IU29kc6HSV9CliT5NBIRvBCL
nVjF3tJeTlX9KwJJdJdf+vaVge5h8f7wYb+QfyKdJnYlHg7Qk9PiFQqShJFj
4bJgZ27S6mK3vFBTPWTyfDQWyyR+VB1vuf82kSvawOGJf/ICVd25r7QowtoM
ZShv6jx8PZ95BDJCxZxg7MjySbYLIdCOgPvK+xolvKg6IsMsFMS0HRUt25kw
6ob0SzuZBtHdwMNr9SQHoKza1fkmSnySxn5BUFPTZp+VPRQncxnRA4zlyNAM
1XmlDPklVXPOH04TTgq7J8xokxJYDVtLoK62qiyQEmr/O45AYUSaVz5/yhBB
9FoDl7Ip0ChGb467A9RuO5gqxSWWVh4jWxLDH4Nn9Te/UIonwBvCK1Pj5hQb
4pxN6D9HA7TA4hkuyHPJLVaP+rvI/+eY+o3odREFs6jkYUHF7srjnyfFx/nV
rCrPzruUYOc2mgFrMDy2KJxRPQ6ytPy0QtVjWxjC6AvRgIkEYZEg3UfJxCwp
o6oy4nJbFp/CeDQnXWEhVIk2ZDMJLgpv2/YryLX00yUfpKIAr7dzpahK5S+C
dhiao/V5YFjHk21X+k8IoJeoTh/M8SmETtg4qmjOZQMToP2tUscNRDTXvY6Q
Z9RaODYXd0j5eqrAOx5zAFhfU0FnA/4wos00gMP2PjfCOC6I8xubcHzwUNfv
69v9Hr/Xynohj3jpHPvPYew1nY+s9oQfzc2G7mi9Jo8gFjcF7Q0tfNpDUgx6
ltIq6WSAlxwFsJBx+1HnXVJRKntFJf6K/ltbjLD1Em0xh4uV9mEPGQZ8MNfb
l9GVuXFjULGaOGUfwpl7B63DNRk0AbTCPOz71GIPDX0689elDq+2PRv34DIj
PGAaTjaFNWVcQQQqlcKFPEDpv36uDMxXusjL6c9l9L0thJVx4uIp/s/8a7uv
yev8L1iJEz2PrtFN9Jcq3Mh12GNnm+lOlVxvlLd7Uu1uQlBrjwQmBpbvmw6/
0L1R7DW9xzSmRW80z/t9KRSH+rPFDPgGKfrJNsKvefiCvK5dDxHNBNU20K73
55XxdB9teu51ThsmOYSqdxQ9EfgGrWEIOxlGSn0ePsuX3xK7xr9fmmkQJlAm
lFxMjuZrufJ1NqM49UNeKSR7e5T98jB5gng78ATt62rw4Kp8eJXI894re0Xo
QaAaTiJpTJjm6x5advWgNrf89hTVpHvfA+ITo2+wFkxKU+AGEdylEcoVZiCg
F+mpOP1jCXZouqE/Rm6XsQXnZiA2G0t4gtUCj0OeJX/NVBzvMzWFyx8l6NlS
fd8sllFOrKKHy2odxj44QY+MjcXWW0c6WM5EHr4I20XUSOwQJSoXzjzrIp+u
Wt+jmczuGCwo+Dg7DJUr62cgMRhG9Lf0pV1wLLOTKDS7lDSgOY+5ESE0aijU
z61U1jT9lyH+Tqtfc97y5WsGZHkOYDpBng/5fS8xypY7cFFp90orGqgBDNI7
0Q3T3mQBAoyKSWTOO+4SstAZv8s7Q+3snkts2pciL0l2EnZPfSqF35uFW0CB
LGoEJv76ex58QnLL5M3a5ZJnNOEXT3r9ysCJQrPUZRlRz+ZOnuddmBKEllYv
HsmLVYPq+VljofyIT8jjmZkx+MPnEde0pUJsPIqLSkwmgX/F7grpcGSZ/FDU
ZLW1vcCh0BXfZwAnbFlFWt7I0TKKseu+3OiH4xNf8EvD/GVgr27OlYhTH/jl
MYzwofsP9XbpWkYudwGMX/kJR18v4AwyMPoiUW1BLoudk4pPIXGDCXFBNcS0
I/uKe2u8ZM0L51AsOfGoKFWP1sR/2xeOXKDUI58LBXkqnZ02xPHlZH2QY3k1
I/5ntBmMd/uvd7xnQG+HoTcyitQkqr+JnoI0ebC4UGOol7xAI9uKkGEUbyNG
3KbHwaIclAJ4Apkahu23QewAbmU2cDg54d6q+tOupXkyFkIwGKkHHzegEtWt
2gds2AP7PR0i/AgNen4QF4Kjxc2h0IpTkN8VE4XFdECuakA1NlxP8OOLuBrr
cAQ7MRkekLI8OefGOsyGa5fDkKMIwGab6Pm+iLJf3/Pr4TJuwx+zwQ/oqYfK
khY7WnylU8swlE51mVhzh9CXL3+/ovGM7Ol+vQ50moS+ojpkoZqLsypkCyJG
GxpwnLd+ZwFIwc7T16yIbqGLejpZxkNTH7uVjNRozfbuDLyc0VtTY/eUnkZf
XygqLVSrzLmIkSQkk2fL+ffcxZT2M0MtIsJv6jl9oR77p2EEeCqFMtwU8Q+Y
L3zZyrdydTAF4k6G/pS19LSQnHC8Ohl0FK19fxMPQE6bAoQE2Ea56EkJtYAP
Rz5CComTfzQ6zVNWlOJP3G4LpofIcFzcgMN90iLJbPcVvIazheHqwtWKq4Qi
DB4L1a1Rq2DfT4Ca78CvfY4XGIVCX9cnHCC0ap+DXlcnlIbzQzXpQSeJ/rxZ
9QprfIs6c4Y6u8znbVBlHVQz5fAQgaQvKzdCyacTytgb7OAGs9adrOepJ9b0
0OSHqLptJCx8OQ2VYi8bLH/DB3YzFaCBbqTzgaJd3ILwI/SZqKkkBKbZcCag
Rj4ZhD0NrVj9Ay2c6zCT8xL3BhszJvzB63Xvs72BcsL+2vwE6V3p8JrwZKwl
un345wxdTO9wj0vywVDS85gFpn32MzmHwYsGJkk7rB7tidMT5Ll9P4IepdoM
LpxkJlUVJdanwYGVIdsIPiVxtXjA+pV9LTI4Z9Urpm5a4oVYrXCjdKrnZk2A
WZFLZCV7aGB0B2d64J+jz0uFIuRBcYhJA9Lh75lnMOc6h2MINaG1uhZwQncS
TU6uw3AvGf/zzcGFa28CCm59vOe2/ZwJgf+Yif7KeKryey1f0jksRvjhSQNy
FOCQpxlCeqpArfcKSwlYtZ70msZlaSTLD1vFnRiuCXr2g7fUB0THaM6qRLa2
tLsjwHpjHTbj7qExltccUzR404Twosq2Qs1UCyF71lKNVuEAum7WyiMdY97D
kZBoxWrro79UNb1AvfBnW7cVfZJH3NUuivHzA1tqHCDQMhiWb8SUqRY+EaJw
6NzLiIqa1uCfAoWm8b4Pn9r7VIYiMYCJ0HHjtyL52YPx2dYf4c00oFNuP6Jz
r8XqFliMHPyAd9y9lwE3+a3Ks951uUU3SEHCjJxdL02fJO005AzCqiDsYwfi
6jsT3YRbxgayEfKHN9MImWTwZ9AMuXYSbAJRnxRJVmfaY6Bwl/JTtdnXLe9b
A5IljzViI1EVOPvGTRcwm5OPp6TjhvlnRp14PpSYHI8cwcBOoFJglrYQpo6+
etrOYCzne2rA/vCMw0yPfNeC3pi8D/YnezgT9afT8o7y/rL6opb6n76TKZtU
fmuM1EQLWZ0N1hMUwFYDCJRGmo3qbtFMJQ+8PQz9vkiBpnNmezey2fXnljHh
n8rPfY2mAtnQU7TDvX2YyCuHnooSbuyX316RBpW1NRrQ65aUPqq6bMI4i5ZU
FAmAcenUZ4DKNbRLhNCxdUxqvy3rKLn1i3DNJC90yfmBoyHnpcT9D7zAllOe
cYtnmRj47E4le2kSmmac/mCx2lugFbLCQWyZ3DE6H+IRq+GzA7wJZBvgJlvx
oBtqWwUGZu6lfqew/zuF9v07eWg19cAMexBVnRUwWtlWOeWEH7R8YX/DbgDi
1du6QwySAoGRtAjVnWS8W0njZQvukxdzRIzlo9f7YzbuO5smarz28FBF6kzq
9qjUAj9j2HUafwRwXcOcUJwnCgzS63nUJp9Vpz84MnhrjIyFvTGKSYIZ7txt
EVUHGxgMkgIIW8LYL7oreBHe2Oow6Aw9Tj2DeAzxUli56RteFu1jaisklPSL
SQHfz/kmRjGeaQSPgFYb9QZcTNFqkviBUiJE52C2Yr5WE5PCiFoINGUyzGkJ
0m/luTIqB1RoVkkq7OSDAHEXGefmF9eyzuvK0g+EIsocRrrKkMII8AQJyNu4
EZvcHF9Zxy0zEFVWnk94BPEiUyyAgM1mThuMXbyU9N/8DAdR75XxKNalkHzs
V11xbMoFmudcCC2IaFAzznVHoWGTDYO3pVqGvGDiNsmhhuRsqIWnlSD4Ydjf
3vY5YXD/oSLfANjcBbbAX6tvV63N2h0rGzSoHMaMyaX29BRw3u0dkcL6qcCy
WOGGy2QtVeglq2QuP2d6HylJwdoCrbEgchaJYqEemXwappisAnSIRNgxd/Ec
jJ8NMKxlXCw6UVwfb+lpmXtkWf5kR63722oyKa3Aqjd+fq7FBG1BXRyVJU4/
RpSlHl7h6pc3i7R1FpERbZR+fcmBEaL9lbZB80pmr6zqiQ7JpzOiF4XHePYI
//swxdUWkLTtfCib1vRB3GqgVF33Yw/8FRfOWIAOsj/LUtelrqgZWsSE/Ydv
zL0hITH1zIXyuUDBHqJxlVlsolQV9CYQlMPLkgoaYnsZOn/03n9ya3zU10Iv
jmrq1xvmntSxO2R8blhFqNDsVQGhJxn0UrWPpC1FCBR3h1B8qDfwHACnoCuA
yjHgBm0s73TduVrglBLiQDfPjpds5014mgtwG1VYu/wkrhvajsTR76C4FG/X
mnJoZza2A8MMO71xJCG/vtNeg1KNRulhuC0vf1s5dmByPVp2NXNut1zTwQ9k
033kT3YQTTzHaeMxs3hIWtsGJ2T2otqOfbANKEL32ev/G6gaq6a5lmxUBzse
kvLZuTPMhdw0rI3ewcG0oydxt4zDRMvuGPAShZW0L8WO2pHygtSF1pkC3yVv
Ew8wCRbHkeLJMXpA+3SLiY4RJiaT8DAmZ+5F65+mpEvI2F9UIW1d4OKboe2n
t0d6FJhul52SsmF9uQ6doEaGW5M7XqpP8HuSGTcZAL7djKEnW0eGDlVuojH9
u22C4MzTsUDWfEsA5Y5JVV9AgejXvHpkw0M9uX7bfrJiCNYgzgP0jPJpbbdN
VH/JGn8eLSpz0tl8TvCCUd+FjQoEq0bDbMC3keDgUVq+sqLQZwKg0gVLNyKT
sB0kvkICp3JcjhM1NsFcpbpssM7p5fdV4WvTFCsMVCVgpVqetHElsY2eYZ2S
Csw1T/rL0KDiwVekPg4KBgtVoMQ3JZw501jRV2l6wYeVvFni3LLw/SlRmM73
zeK7MCWQDnrzOdpLiNTq3HsvyCexZYNLv8m5Wk7KIo/ZEj8Gn6Y1wk/VtL5U
cCQdUw1r1Hok2UtKKtHHRXvv1fkHPRAHqgz6Sw438c6ZzNVS0eNghcqmRKxz
sd2iUeUdYKoQknEkNufrT1EahGo4pS8agbdAKeEWA0egmX6S9zhmUuDXjLR0
m0Nv82wyc5UfWlztqq1FjpToO4mloP3Kw2bpQzKcFBsYrzcSnzbl5MSQkuSq
IrK4p879YWFXDadfn9+EnsZYU4t8ORK3Uv9W+aS5b+KNelnPGG6nThAF9pf6
7empbL8EJ8W0SCKJPDSRp6+i0cHVpVtk8IYP3ARzH/qrKzcj7+zJahKjH6Pj
xKK6tf2QkkBhw47Dd5gUIihdF2GMljONBQMxhjqwwrm8Ka2jTaW6Wt7t7sY7
sK0wEdmJCQRuFGLdNg44uVsJV9rKymXZKLqfWbJvpzs6uGyHQyiABnJbYDP4
RaqkZbaWg5+aqz8w32U+VDZwffe7FRUetD80j8DQ9E5WpJbOyEoJP9lMpLGg
iGqJIzJLbgqIE7CEDz97/jmu8muWt6yNhGfu9PAArkpENqmdWHl5QKJVmlC+
Cf2mTLJi0HgfbNIlQDSaDMpJk+GTv3c2XKi/4VvK4BBay3Y+ttFdJLWYU820
OSPj5S/WbMtczYALADR4MbCrMKkeT8UgIpwUbGxl8OpS9PJAJwLysl+r9aKM
2nMYGBJV5PJKV2/WArd8khlbyu5Fg5IYtBLMBVKWm0122nWrejkJNk+TA80V
QfsB19pA1t6LNdcebg+0vEOb6BoXYCt5vduKQVvD54AFLAcED5ONYvZLoGEs
hFlhyQ0jba+7OZUqbhib0qLw8YUb0Dza59nc5M8DGUgmUjIYz9nw3LETE6Xp
3PuZz6Nv1kvUsbmRbjVckleGnGspeX3PHXj/2DaTOvfGG/rqKnk2wf8xGRgr
iQ965zcPhf7+q50jYyCSJBh9S2rh6Jsh784b5a9jrCl2/lNRHMD9lpnXKHl0
KYYuqRs1CeI4HVSZrS498VGdQyRbDBowMYX7TuLbjqS+Sm3xxou/QnYzRcFI
NvjQc2C6hT+qZfhx3ffi2B+l3DlGei1TQUYW/fk+Bagry3zQei93/7G6mDMv
+gdj/9g6Vz3u7fdcAWAoX/Ro4VdI4wUqiXZKVXpCKfir+oIUdl3R8Om/uRID
TVwlwve2KI7nmfvKAYEgjOSt9P5EQbt+Q3MwC2KkZ74g7n8wnUiyFzNL/8LI
hB6fUhS0I1PvbVAHRmlXRngtRRfzBHC52jQ1VrSh1iK7Nyrxz3saJdzl7FOs
c+WxBcm19M6v3aA5zhY2FVtrZVN7VC9gqj9yqHHy73vo+zH3S+EBNsxRz3fN
6CUK5/IYGrAn0LbH870T3JzgmKJX+MdGTbxXC/rlZLzlKYVKTdaZZ8SmIV+o
WCAufTpdlVjHZ5nh3AGWtirWSju1oHJOo6JJAhPRm1iUPhcqz5l3QnZyT7yB
HwClk3MLNLJl0zOJ+kC/sy1vb3sqOemDgVBKHToJuRRZZa6LohdwukWE3mrY
w9WR2Yw4SwKdxiTcZLK5eArv6fshDKW9rU/L3sGAt1j2WngzugoCV8V4v1zB
vgGvveuMBFk6vxwXi/sGaL5Unq59SbKX4O44KkUvdAQmPpeUWcruCzwWyf75
tZBDxvuup+ar3JQOhGKnWy+d6e9Qalnv8xX58j6TDk2lXbnQmm2+8YBYK7ZG
WrK4zhFqdZ9aN+eW/Anj9ZDtSHx6l4p6++csfoki8DsNYVMw6ti+eCpHCtjd
Uygc7jB8IajbrRn9xr0ZRLR5NkpnZrOub4b7e2GrrhM7OMZty9pHnHlpFD0P
NZJIs/Pdz7FHfdG15F7BI4YZAezh8NpVaJqaZDR0RqmhFXGDGARWnU+OkYUy
5IYSDM6p4Bzv39mV1c9l/505bMJ2eNBbiimPoO7a1CGN/yOMiibK6+36qbk/
aMvMTwmruiIKBExqvSsM61L/FCDR5qpwJV62nhcgpuJoaUsHh0OQKo5S4juv
C0JOuc62AFPcSzdEatJNRtty5PcknGWjOGCWIghR7jAvibVGZzs2LbudD4ls
XOr7SYmWiS3JelhCfbnVB0b0y0aO6a8Wrnh9xSYvEF0bqvlAdisc5UYKXDKX
/wQl7jbd02IyWlQjQo+PZ5oXWsn5xO+pDzTd+dl5Md45l9p+TxPzM0GFFtKg
FRj5QtUT343JIvG+j8COsMwGXtCSCsQ5ebcB3SL1Yjjl/XwCkbuaQKkACH2S
hrVuKyUhS4QeUFC7jjwNWVE/KTX7fYEbTPTNurU5zBiLEStP9P+lrkGUCzNN
484xDyU/rvyiTS+dFreDAfwSzAHFJPcDmmU2/PtTNKgsUxpeJQpfKEjj21TG
ZNq4GUUQnWSLy358/Ho0D4Aga6qTgrcK6CHvjIv4zexTqmjtX3v6nMy4RxD9
D1ZX01XiK6Kf7s9JoLy7FA3FuD97IUtF0Di+VzcUaSz6qp7oz/H6b7b3ZdKb
khcnhikAzjDWNBSqkWRStm4eMOuVJnN1PWhjnmbSdPRnMkH1huXhMA228js2
JTShqLoIPYiiyZ07a3cBjU8yKWo4tFpFM/WcV26VcjE6BFYMUfLdwYPXQ4Dz
34UwCtQu4+OmDg1JHaEVFSpFEik4EFUSuoO4yCkc9O5Agx3s6ReP5EEBY39n
QPNnpHwvxV1sLGJkmKI0gZHRvpRz/ZjwZo0EKNlcCRKiRgaEh/acybCvrKdt
zPtY55a5BEIlgxkjfi9JW7MNsoaqfEAb+O6WHhmNph0w1BBfl/oHxfIFGPd1
WUPco7qe/52+WDqjRB16k5qDbkZqcHhEiyRhgFvFNw8G57mbeY6IsgcN+ucu
MTODDg4iZUfTtm5PGBk282dUKw4R4l6GKDQpawyOuEiwMfitUi0a8TD3o5Ff
WHtY4tTTU30FI0XhsrvvlT3jTE/g9S+7aps3l1GxGiFKcW3qQFaueyn1mUzo
EB9GCuaRR0gaHKpXutGo1nXB2LGxkLx5BjH3JGPCG8a6ixk/EgLfBDMsFw5x
rLS9AhyCa1v6xBRA3tf1BBIHmf6auYlcP2Q9nNeM52FqejaOjg5CMq6Iksbt
tAJD6JUBEby3/M9KqS6VFdzdlEWnNDgDr5oBf6t+ezj87VQdwCV2miJW9stc
lk9KJFvVZAOejh8xOvkrpChaTgAjWh2Xf8172gtunOZj2bgBwPIOfAyPTubD
0NXx2Srt0wTSPbZRF+dsifS/d8vGO8ijYeyetmALblSlfnS87A4Vn3urzq2t
c9l3R5hIRtnJ7Q9ZGboCKmxz5XNr8N6j6/riFYJmfeUwtIviBVIplHjlfAZv
P7JG8CWxOvPiH/+J0Pf/tsWurtH76LTSRpXJoqdc0l2R5+gQE8bf2aRlUVFo
Q0mSZNXr9mFCEB87n+t6W5tMNlPYsQgAK5ZHR3gtXMujVjDdhzh9EvbP/NUG
bZ9PVGUFfLilsF0VH/mbAIhdCuOunS6maCNxRZwD7Wwnwm6VnHTVQ3CTGQX0
6rlQyZ2AaaJc1Cit1hYuwkClBAlgN4OddEARvG3GSXvpJrq/F6ZyxEnX2+Gk
P2y8Mw2xgg9ogRY0tKv/X5KrF0ZVMOHdbGWwzEGOVeLI+cpmXhB7wb4xnIdG
1E7fXpAF6HmSsoXICLb4e8loHXmdJ9tFd0Fhd9s18sbEhsS07IAYJSedxEJM
a00ihF1CZyZImrXB4cl7vsZoUTZTRY3JccKnFS7neepLoqnNeOX9NYYLtqog
qZhyUplr8tC8P0W0ZxjfP3c7Doof/GAa7XvHBaAtsDjSufsk8moZQefdUma4
VLdDc3yZ1TGtxYgHBqbhPuxSSw+NWMsSI71NmrXcWoBRoinXB+qT21Z2/iah
qu82OiobIPQkxT8p//V/2NjxQUU8WJ+D0fpkfVUpaXiCYzCTDt5bj72LKukm
D+Yun5iBFg4vw4cLyq6wtKle6ZTfmbEh0q/9N+MYEx42dg0CpDPnCdZrP5Iu
As4oQw8xtxQTGD1pyNWotVjjxwOpg/UdUpfrlUqBTZB0wz/XXUjjjXyf3+1q
Ica/m5ZNKBfcTuu4RPa8fXR/1L945fTA6FcP/8l7XqEj4GMWiljWT1iQdXdW
lQ2XCvP6dGILdayS6ZoDA4WdgEpn1sMRumQ+KWJP9jzNFryVWmYEnmSz19aR
hAXN6vLxgXNU7enVv77TR3MgMP3VgorJuxMSJ8qbB5bzbpxG7dRRIDGRP0Dx
pLxrPuLgHyQqlYCTbuaQfZeVpOC3YHMovNJkSfErvx1oLJhpsG3EBGlfIv2C
H4TWn5b5Sj1D6FvQsjrqP1alabSf+nILf8EBPtUvVPcE4V7sPXG1HM6i76D2
DYBNI5G3t413/xd3C3MHUCA5rtNa74K6cENS5IOA5MkLhlnO54ZtEHxYeIEs
SZzDde4OJbpw4M8Yn700zZjTTpy1xCCnBaDcssoKU96OOQpYW1nvGTq2hevW
HiU0sdW7JVgQVjKKaMpWMMpZN2bt8fVbZ9/5BVrzSjAJMvKSfRlDJo0cxsit
qECeUG7Nn8ZZxduXVP25ccYCSwHgp8vBwF2waGX/gT4wGrwi8fieS/xDFDh9
ikKaL4KRfCXXvjjxb0F1kxDHBVhpAukXuTkM6o+PRPWWZ3ekJgd0MMkCzjeQ
sdpVyTkhWGGanukOrShK3xOgZagcMbBcg9Z32R661ojxAlKksGF7KZFNVZQt
qC03TuM9na6lB1gS1SJzbxhllh9OibNrvWZjqOh8sfhlZpYd3dxsNIh5Km3N
inbSH9/o8xaZCiu3ET+FKET/q5Lc1U6RxqY5rDCOPGRICOKTPmB4ikRnnELe
ylv8R6Y8GwRsd0TqU8MkZ1sedMTEwTfaQGZ9DzQT6E6bZL6xV9BHcVJYBC6D
qu1+mCG2Iamok5xx/UXKUkswwsc4gS42tw+B+6PFJZtlFP0qjiXTx5UvM2K5
Y7Z6H0tnqkgrc6dMdkBbky+zzl2S3NCRvibK7etrDaxG4KfRyb8B8UbOb2GK
DQlowSZ+VUzlfAqDXLIPxrV61wQzHZR0ZBu4DtMfSWjpxBtquQucz4j19l2l
536UJn5ICHp4Q3mnWwOjvph+t9B1fQMyfOVsVDcxiWkfQTreOnwNk7ynJbJo
ggvDhRhFf4HFsLIutJloclpayUpaVkH///NrWi05SiDiVGoK1ZiN0kYK1IfA
0hzfktIqvakbObTqglbNK0aOfrtd0JOiD+EyKjcfoHEjFJ634IlhXo/ksdcT
yPkNBCbpXqIhvURNm0oB3L9RTFDp4ffsE120OYwhjqSsvHHBQ2o/2FgbcZr8
c2dp4l5Vkm9ld5UMMwv+/oCOxHh5f3Sq8FnKtnGZ4TIYR3wliu6GI+KYtE6x
Ibp75FGhcs3JVaYbNP9SPB47QmdHOP+w/h4ajJ556WHMOeZhvTjO/EGijJLc
LdX1ybYe9NeJeMrbVAfQbLOeY6JlZdmQz5nEtgwA7F9K9kLq/1xoKtvNVs+k
vbeCkNdr+PsJ9VVMH1oPM1jle9IQspaaM/nBL6H8DwaMiLq49l8rbUJQcq1G
PHeinYE2+T2MECBfUbn3fvoPgAXCErTYKUb4+ZnPL7YOrAzZDb1OgU3mF5VY
6AavNvsBULRLwoJC039Pja8yP/cPgdnQ8fJ2FXWv1zOmtfHEIlM++x0LxdK4
5mQuw2JDyLAmOtpaHsGEc9jFw8wSXjcBs/kW5WdafPUw7heSeuX8Fqz+nZL2
pD1WMBG1XTIEBuy0hWWjQ1kSFYYjDupXkWJIrZYG0cpx1qAw/hjREheiwhS9
Gny7P3/nC0IJPXXzbBwM45R/gXxwBSSdW1nhgOIM7z/cjvEEaxM8MUBtP7pV
okzqLxPQ82yb3kQT2lOl8lOLSVxwgJsI1q0eYuMCC5bkmZMzpjog595z8gG/
mQJJC0gIeyY722X34ZrVOuaDcyALrtIpdGL5nlUASa8XIZNfh+kxTLYezTE3
HIdZ5wfW0tI9yd5nr8MLQkjLBoF/ou99QCfp8q11VU9W6rzHlUtMQ/5cGWx0
EEGTNxgMtjvbBsG+pPqcoIitWQlB0ncNpEAAyS/PAwPm/NUXvATgyYHh9AfQ
BNRqajwEmOsIWLzMpO1y2hjRrdPB2G9tN2Xavpku9CU7P91re7rzJohNuz5H
pH1lz78jmGQnFyzHATISlQ0WSsxJ4m+JFTAMSCy+afnr4WFIsYKLrpz1QUzp
V/8rKYcnO/0xth6EubGKWqeNnLcLCOBkU5MGtMbURqnpQuNnbIZMDBxGMLmc
bGJ3gXsFu5EKcjUhSKL9/3L5JTZclsNEGrtmkKfohhiljfiE2cwLrZX/+L1X
Ftc7V4FRPS9BbbihSB6LQzHnUon3L1fDH6ywFmY3MhE1h73MNaF907J57pL/
v/fjy69qg2OWgH0ttCf00JeRnN5pQB44JqRVtzSwU8xxkPLGFBgeiwVnCpnj
ujLS5fVEfTMPo79Cb5WOcPhlPgEHoyJmdFVMDyazZtVYB07cZO1PZQYmGJ5n
QdxkYcRNl/w9HEDNh9dWNBrPxoObRaZbRYvRDh35oTSTk3X2JPZ4nLrpnrmr
xX0AB657IcLVgFB7OD88CXczXHpamTqg+Zifwbh+jw+ZeGxAzDuYCYclUe9i
bUHCEtXPctfPP+JKZi8O26XkmODG0O7X5P8r7PFUwbwMvPrSU89N20tuWcYm
MwRRKOc5NCyV/b93L2UuV6sqGEShjKEDwO+p57F3919x5WzKHjnZkd41jTif
49Exq6+KRp4f838toCUrDOqySK6dX0PYVx+dtDU6VAiVQO30XPpL1ZRR9Z9G
QjzwCzHFi3i0Z6tiNp7jkuaB34Yy+pjl0JynKRitJRBVFPxro2UyTg99dW5u
3EI9wWV+psjGcPYvSfNDswaVIvnZYg8QFuwBa6mepVaNixD/Z1cl3mvjShdR
+fvOhnHSmIimUj9VzxvQOKOcvno9jnyCwLFc37O9JG35/VWSJDOdQlbV5m5H
qn5pjEcitQeDRF0YMSLSerYLHMJYqG3lREtMdAQEzRtezwJhl0FGMIPtUvKm
5AYJL3wrYzoVSi9phRqmQUTQfE6Pz3n70EYyBtYUcDmekdkTkUgaO+RnPfY9
/KR/Yk2KnTXbIiSqhNLBCfFUnPThPjdPOF2rc7Ggxr1sBQ21swu7Zx/ta6sk
7HL0GJmWFMpRbLPe/6CcFNxkonW25LZaYup2+fPNIORwq5Udo9yoaOskskFa
D4TSQWyMABupvRddQAOIAVcuja5bm/cGSDYkfvw2ILWtg3hW0HDFmwKkcdNu
ghYvF+JrIhPT85URRf5wGEogRZLTUnP/WkDCTm4VS0ALwXGj2ul8dieUvR1V
gvTQuOArnl/CrZzFYgUUbIA4FHX1+uugexPMgHBaBXQLxUyIgRb62eJCi8B5
gAbegyNoNXcoOSTkRGYdWXc+ABMk9qs5ootBtTQravoIQ4sP8VNdzh9TUl1g
yMsyZufCV03nKhZQGExRlU76TzaKvJeRYqWTe9kp1YdFtQN8oCea2lj5Etso
Q++6q6ZsDiFwuwK1ywHE2Jue1Hn9zNPgI8ZrbkUuk9gYK0CSvcwGeRlB+nQ3
8p2aEqU2taxdDtGogdlqspyUrWyAYif9zHlE49U57FE7//22Kztn1Qn/HS+o
pS/goL0ANbm5/9DDyVZqaPZqeP2Pee8SnRUr/zceH4brrCkWw2nsPXXhBYBw
TzNhS9YYfA9CaeduVg/hfzrorG2Ur8WWeUd4ePwWOOKPtcd/20jgZULaFngz
4SlkEqx6TchLCBGWVe+vog8mQmRmvPvbNdFklg+AAYDJ4LxxPE1tWKrcqOwB
ld05pM968sxht3HYfIHmV/oHycczLnpnAsi7MRLyCwbi8hokQ5+CC0pc7Jeu
QcReHMCvSQ0FWdHsonLXfEkzrxGQLSlLDOKsBPoKTuIJQTbS+2eZGCuZaVFC
dIkZWkEOYOeZOHs9KhZ58uXMtKLouwgLn4Ae/B4qi4xWV4o9pXL+MmMb+gTi
EhUqDkrpZNhyy7wWYNUb3O8s5nRchdWZMKGtqdUTEoquP5YXH9qS9O5PaIxE
QrNHcGD4r5J41nufodfRrn77TMUFpMrACfJqqQRnkNRYXN0IohGkwSBxjoa2
3UlN4P9w4mD1XZNTwbymZjdj0EeldXAZB6aBPim7dZ/703QgZkqm8tiUyjZE
ifCNDd4hXn0KoSuBZ/WCfBazio5AVfnnlS7DbrxjvS2NOilrOoT+/AE2k0V0
zKM3tZDwcKMhR0s9eRWZvfls31r8EUnQHe4iLevewYJmHa3HlyII+Q5zZ2V1
7vm6YIw6qCH/fhMpvhGkECOKxysC9Fe5ZvPFBxCZoL71DYx0BuwWdCXkcMUL
1mqAMs4tcIxnl3ERO4Mu75qYUnYv56U6sPxwEhS1AXFTmR9E49fF6Kgki1qC
Egw4ml/lzBUmHRUh4dqtENvbufEoxYSVB6oIsuW95JhQ5bZDpMQA90sWBAZU
6J2qw1xHDZZTc541nztRydO36w58rubbni87QEFMqGodMo5rA3crP0U7+O/r
3rYYQm0lffyvzbIfkvuZ/cBSuiYLr7iiQ3MMjXvd3MNoPBAXxwzFyHGewYZj
7vHQvSRnjHrV79z1eeE6EAjkOtrRqVsOIn+6PCc0R5D2BJUIIxMufb0+DnLs
mxz4LaDYxq7RI/olovorh/FfxWIwkTTSeqwoHYowitHto1xVqDUzRnoEAzFE
XfQnJQ0FawCPa4OQtqqueHj4V2p+IHx3KFYcJBcALQ7jbcriUk9Hs/QOiwau
zzO+kmV0n75qZTCw9sN+SHnr5VGBrvU5wXH0QWNx84KYY+vLcBAnPhgBRM9i
bhX/p8JiUmVYkkVjvC0Ow6A8vs9YGZeHi3lsUgbGHh0F96jhqZpr7IvHos0t
FnFBEHLACWW88oyI3IatGoeggUxLxNvQt1+caZtJSDJfQYwtr4Vj+8LJ/rL3
EwM8VajurJX4vUpmTuDT6KolPV+y7a2nsk4tUD10shBolNVTALtBVlpG9u0e
aNjShbU/YzqM1x2K4YQR5GLqC69ceulXd0iRfX9Amj3Pz2ggaSJR9KHtt2NY
QmNF2gGVv3hbHqQBPqquMiPuLEQdOTRu+3mUzW0oSt86U9HLDV5qn/Kpi8AU
mWM0XIbjsLdr6ytJt1Geqa3I9RGCBbSBct6Va343So4HQEI6kRXvy9KKltgZ
rlfyaOqu6+92t7hb8vzZbbbN3zyjsd2BRQgrbPsBo1bvMt5Pt1mZR4HmL0cp
g9xbrPn/2H3Uj8oVtGDqqXbsCf4sjPVm0kPJ7ywFF5RJYwoXyo+k2VTQRBhI
Q0vlq339F4YsZJbwABt5NCyxZEWujLfeNmuJn2CE/+/yzZ+EJAwyTWf+0v8i
iy4KHfu4RXSNc9ClaM8GH5V1zgMW5GUZpZV35+iax0zal3e4Dtk6QeIZS+sK
z/8f1ZhW8xddqsDKYul+YH1whS4fhQ6VvLsq6MUOg7S0W2oStNV7BqDeQ2a2
ngboqHXfT5fm/5lAj0KKI354ulO1LOHmz7qyAohbr8MZri2rKcqz3quamTjT
BsFZ9xnBkSRhC2UZR02HjME805QdpFuiupaKbNWk0VXbSdjhu4C/BmtI3DS6
XDHwv7td5iw3jN70OeSX37KMO1RZLlcOpJ2LiSMzsSFx16qf0uX5IeTJpO3j
HRqTz5Wkml9+DrwKhxGwOFdt/T8Zb90IPc8nO1ts9hKjJi+Ua7ZGt2rpyKh/
Ex9b6XHFB22cu6U/XbEOShckr9MNVb3gE8jmeex0lgJllsjo/PF8bcoRHhY4
qv4wbo3txbOAmNievgF8kBmNb+muyEh2Pg6HhgiRifRc9PT5mVk2IXveHL+u
BqE5OKmuYUV6IaZGc3TAG0EzU5xKPcE1QSSv/s8/1NSunY+z2yFpNXI2Cfe4
Vf82T7DXiD3QNNORNe1Xn2cBGfNOJ5fAD0usVpdpesW6sgp0qBE0xqajYa2Q
6aSGopL1084qziCDqzbo4geMF5f6StA+DbVocJpxiDa22vO/wi7aJp+fkrAU
cFUswJ0/nQm7y1Mzrr7W0eGD5VtK8Bhmd3BMZ666XzQXbvxjn9flUnboqYNf
YQ8dL4lYHxtTcpgk7JfHMe0egYtlvkfvaKgBWjhFl0qktNoako0+GEc++yQ9
8OrSJZ4breeSCCjzO4h/9hV2M/uzFuQADIePZJ7N9S+zR5ZnYTeJy2hrVqR/
SsrXCuU5MWPN50NZLOS+X54gVA+5am1BFy5MPJn+3mSK4RsFlAVc6L3RFpuP
10GFMHSKr430+eULDAt6zQVSvSzn7cYTcZQ2DcwlNEBxj3IFrUNy/vmh22aL
IsbsdvATxEqbboD5OGzc08pk/jHRDCv/Q26A5XkwF0Jcv/3Al+YHdLhsg57v
EsEQwpjq4TOElwTT7VFxx5HYM+bwwWbfUBtxt1W276Rc33ED+cYzUzsBh4qH
Hqe5QOhnysUpdHkzS8cpgDhr9zMSyGnAz/LkpvuMm0i9cXRCjloB0Uj+huIY
KZozl5c/3IqJ837kNmSgRA2PXkcEkL0VkEAtETmNlmcXNn28dwJyVBEqAarg
xOAMTTcBOK5CNmHhMHUTAhjGlUb3CbLmALsyoNQnph79sYv7wIY7Ql/amMSV
OQYGtCqfPeH+I8TCEaYCGEyWxhexUo/MR4k58OZgBqrf5KwdTbhCiMq/oQ5d
9UVoR0Uv29toP6U3zE5q+MufJRWO5dCBuqFt4YK8gWkcozsG0w3nBp2tOEgI
Xl+05UJxSpmclXNT1/k6OFv7m4yww/chjUW8cEBMlI8mn5PKrQe6eJSkDAGE
hP9HhsRhS2JzwmOkOcHBCpg/bRKoQSC9ebXjofdisTgjVqjcqZ/7OsLnIsCN
4lCUmwIrBfraFgwlVOUhoy65qW5D+7WdjlZchCnwUpyNtfVfwjlEGGkXgNrp
67Z7hhOM3YpgnjKWzgoOpatXKsZB/nZAuFh05eha6EhuM5h8cyG+6+bEVi8u
ALnMv+ORM8jd82016gQbGq32ckaaQryO6vCrP0T+g9EO6ATntrGmp0HAZmur
A+cbFKBy6E0f2CbdbbLEZLEjN9tQoozkP9ngMs1bzarKGHdBXo08CCvKu3kb
KcDRoOUlxO853Cyc1x+DMpPKURsypHId7TnVbShS1d3xZuv1PkW2NH4+X8FH
WceRNBt6/oQUv7XTjVDTniDlJufy6Rhsp6EO6NQDitTGaEqqfpu69lZdO6cH
xBi9rm/D2KgCsJiXXITvJmrHcNJOWkcKkDG2lbvm19BhXEgNDq8xW+uqDNkj
NNuxwMYLmJDRZrndSM1c5HJjfmsNfpo1guo30pMpNUBbH1NzFWMk2WsqZ2Zu
hE4TeDvWFQkDwgF5ccYEl/S2U+0IXTb20/vmcbqL1ugaNi3aocBkear1eEMN
X7r4UYEWqUnjT8A8jp64luxUqnAdZfbM1qR8x7SH0zu+VcPGFdeN+bfA4idp
MUz1imdzIqWe+l6y6mnSq+IJ7zw3BtZleB33HZLr3Ntfzm+WbKAsBe8bEr5u
dyhUSEkzmR8NtQM2UUMIr7hcrr5IBulcRsRRPKZWQJJW41NgOj3lZzi7LURu
jwSUTb4v6GIE9WwxLSFGnGKtTpDpp6iw+MmmLRI3VnIq1aCYHpjazrKV7xwO
j5nDM0hGN3C16yzo0rfC9Tp6/H5T8hu0j6veeq6ohSVhecI81GpWjrQ/NPiw
lc7sE2/uKWF4TD7CET6ELSdqQIRShCBKyeqTq/sM1iEl2McmaeIoUSu/FsO3
tItYECmblhebMiZB9cwg4EeXJKVm1TZ7CniM0LNygaX1qAFVV4jxs76Cb2R9
HV/JXh4cIc5ChtKNhEgHAB9+K/3UEPDAeSNM2zyLCChjSdQNxgP35KBO2Bo6
OS8OzUmk3ncruSR6TOUItD9Mpn5r2pbpJjh+d6JehYS+IhVctbFTxGoQK2Ri
Dgg3N2AjzC9LXFMIqLtpgbkrS67ilpwbKFWOrb5Uvs8gTnoIEPsHyCHVyBDP
L7h5qSOHkiXqIz/CjgOfSy9XUcvSLxpbh236c0UFZ24F7OtHUdfdDtjCYx1x
NCJiPYW7RKgvimFgoTnUPAQK2O79Tru3T9kocBbHA6mln7kwAVplo3TJ4jnO
btCDrNfwUdloljQHQkynwhqyNh5EXbhDPD2b8O5YdPKQboxMXntQrD0R6ljv
UV/NQV9Kw8LByOQ5rgnrHbjhjh33zcmgtImjujaybNV3eXQYzRkmbeIh2qm8
sg5xw5y2JIuKg9zP7V4g+28vgasN1xcNZcodYdFKtWkfXiUxc0Uflvku4Bzf
DlDYksipRnUicI6DrFJ2tUsDkoJRWrnvSdZ1ml34Su2Ci9vsmR7ss62UcqDz
3iL7W/OCIvUN59LahnPuGOAXeX6WL5rXmZIuaqBWbpA66miGxXiszSdedHPQ
oMJVUNOxh/GfS5GkVlD8mIUP9CljH2zpYgvu7X/5WnxO39fqEfRKcffStk0O
l0I1aTi2SGQEAdyLk/C0HH+ikbnCrQN1lBlqJXMwRKxOfsXP/gfnEUM5r7fd
ARDZSpbPdTcop7XR12FMZ8/c7DDx0rOHredNqZny4LeWiqfFc+9W0p0cOqwy
uKfEQTtiYWDuxdb+y3z2d4Zci3IyWb0RD8z70wutkYiu9K8VsQCfmq0x7gZa
dqvWdKTolli4Xm9gIY33fLTP0N1myPHsPW7gSdrJtz3hwJiw/FGjrVUMU1Yg
p5nrZoAZMXXf7/laFvkh+616SqQnIdr79lac5/LWU3ZRIgVMVXedB1ENbaaH
CFr1yeM3q9USEbfQdHDCQybB/XitNtCMENtZGG19FEzE1H2DUydlS6ujXxPT
jsofeDLNlLEkR6LcDtgYjcV8WfLbbh9DXs6PllpLwwjorUh0A7t4cjQ2zVPn
Nfdsnlw0H1QgSg7LWFZ0LU8lZz5qsBP5cI6EMtLB5CyfHuUfV9pbXHNVZ+75
gbyZLnxlUBKNYtAiaDPy1Cy4cUvpV1BQ6pEZHjFIv4CN+fxG/ZrD2hF5nKlo
NCdomc7ZoAcN6AIimpAv4Yhyr7ZRo+I8+QouycfFMbyAbG9HTVDmCSm5Jw7q
i/pc2nszTZmcnRuOBIMVf2e6WgHvBH24sUquPBNpm0wGOk/zyydXFZxkvCva
2Yk/Q9kyiB/4CQnhnyu3ioLYc5NjJ6MieR8wt7ppBARukvE73InrzXxjDxK5
/LZJfaF6WOeEHcIrBjPW0z0pxDsQCGfBDP9KTqr683NNi99WerDSOkDi0YUQ
Vp5lj/ZQf62uoNaLk5xET85QzxQroKInCbAfidhuE4/gRzMBCbGPLzQTefpF
S/2jt/9qn7Xbofspj6k3bNU2QPn7jnYFanEdne15dmRN6lEN2hfaSMLYu7q+
IMxA/nOtk3lTmByCkLK7eqb1PRzZHTZgPIR4O1/sOwnAR2f+axMkO81XjK5k
c1OJm/aELQkuUCqKP5KrzkgH/0csAkbKNzVh89vnmnyB6EJZ5PmD/fSTJFU2
nt8CaW/h00Tg3PP1ms4ZXNbOjp/GclFjxob01tjIXhAC0KBGEkAzfkievaEb
vsGRK64CpaMGoadX2grbJsR/AnYCcPhFIJMEudKiyyITzU5bAX8JHmoR1euB
yAS3KX/kUcPJ2L5cJZDa4kBrWNSDLgFhaV5R32RT1nUKGAbKagsVFaxJD3na
8eUEpZbl49LDOJluXPKSMH94GPUhJxd0WLrG6KLLDVbVbfmrgDnkfy/UGW+q
sM7gA/qv120Oo2zD19CWcvmopWs3RTljwMy0Hb21Z0CjlcCSUz4ypfX1uRv7
msLFh5pSw80FtEfHrnzmtleFbhuK4yeVLJYeUTSYfWwQvqOw7X1icYfxe3kI
1i5qFJMsA580+5elNr9XXElS68iQIlQakCSce2Dc0G2k1cc/3IZtlOX3o9Qm
YNgrOa4+4HhW0kIj1OC/knTltUbJaZFAiAf2kweSVCIw0zfIbddAkApuAS/n
ZeYX9z2peWqsp7YIvK5iz68MYIKB2ExkauGyzDM7SSkWQENy989Sp5C4BGF7
zWbAcFPfkiuNBtrdZd2SFWUNHuq1VXaHhP2rh6EfFF6orXeP3btBSJbn8uqf
5CL58pwbZep93vFcS5QDty6NL5WKc33thR5v7nwdn+P8CMABk64jCTtJSJCs
NbI+DRAOq48b6VzeXA5M67OmLTzwRV3nqj5lr8aiBdke04fFLShekwboDHvb
S+uP+rBNZZR3kdx4KLW3EcVube4SCAkVQ1lCvuqWqbsGV2XdGEdZMd33JL5K
NWQ/eFcM5ZMJTlB8V7H352XA1k5O4hW0FpAjybbk6rLoR/GS/NB8RQk2wBAa
6GHl53jIp/6l7JC2vOqoYChXAD4odOEq2cG4Zz45QYUdYr+HJmpkQZrScH0G
EfWPNseTQZiQesb5KLf7wSi2g26j0BFeQZfCMExy1Ji2lnUtW0CUJ57guWL3
dxmblM6uwl4RpgeAE/cCIDzamaCwCk7XQJvqxqExvGdflAlj5Dru+Hcv1g+i
n+7QNk6FSQMGouBMrBfenn57Urd1esIR8nRd4eSmvOLzAM7dS7dzpgjd9rYL
LN26t/6DpNPIoievAoSx5wGSP4SG9wAsSIOYFfWSPI+P2i3Pg96CCu6Vb8Q7
sC2SjMsEEAdzpVohktXN3QXJiHUgwuIOom1uUbHP0YKVbSd4cmuds+PcWu5h
SKXo2ajB6O7zz/YCir+vqIG64ZD6EnA5i1gl1Uwu1HV0LiTFy2M/rhiVDhws
3mpDlGBhyz0/w6mzexkOASNEapluY0y+E7yxc8GuF8FRaPV+XxrIQG2HwcZi
bFXFJI+6sGV93UvjmQx24kqjx1tJtJg3b2N4M4JvwCYvqQepAoYTG7iDvgJt
uqdcRaMnhQHVNWeu05ircdXim5MG6abxgCgHe6dStj+DoSA2hoWVuy23mNj9
rI/KjmowSCZQvMN0ZFGIW4Xrl/I6AcaWrcc/VfK+ABEfMJ+/qlq+m0nedLik
xn18/ZWsI8LLKROlljnKHRwOARDqkF6Q/RQOK6VP8m+vEqzAg/Ug4IOzrIce
Y+FZsl+k5gWpS+2THSA0ELOsLokscz0FZjCNjA3o8r/wpXY2BvhGrG++XTBc
lj3ld2LORjwdqhwTrKU4MIlzD3VgtivIoiJ7Ds08E3kR95wqLYReecnEtRDn
GgxGfZTi1MXZvp9TiRnr0mPF1NAhEb/aLGBdGdwT+5IqhM48DKv1jLri57Y8
AtvaciTXOdJqSeknjWwptiz+t2N5cJZrs7QN9ZfvQPZVubOCulY76ugoHEZK
nh/yTdDM0uq414PebNMVhbg3IVFCX9FDGL+Y99Qnsww/+79bvgTYhMUwDS1q
a2yMjJnFgtzxwgz8FwSOCNhkXqJRCwv0BMjcZDgHvWDVIxgF9y95lckhsnT6
PhODfoqlGFESPAYwLVBosxpBcYXL09X4nT2qBxyUqYngd6aL+DvJ1eA0J9WJ
cJP6L4Rish6znT8In6TX6/EJ7nmueyGJ5+lLWFhUYtIbpmf53sBgwsRMs1Qx
fWPWLGdJUlDYV6FELyHKZPDeGOuzADBhoobW1qJaOIp64uUsMLODCowP7cvh
i12wksxtopkYJlJjltvBeQOQOv4V63lAUq8rjRP9AfLWFwqAQvMh3NfSL8SV
360DtsPecdLeu6oA2d8mZFRsA74aptLqQi0BZR0cTz1AEOuWAFTIvEGt3LFc
DsPcW9XBz9SJcFG1zZNY7aZ09rhoOSVYQv7zx9hhvWNPOKAZzjAwKuFN+3Qx
Dfzt0aAkjFumkrL13fnIS9mroO14ka0wgFPzIqSqmHybedLeBZK36VSWpgg0
N6CY5JP3sPoSnnWq40h1Po2PsgvwYjoeG1p9XeWSkf/x0bXy3dz1G4eWHXpC
alZLQWjYj4TB/tdUvkR4WLywCP0/r4U/zoWw4qsPJ5OF0rJNto5mrCv96AGS
8B97AkplI5CnldWRs28CyRyYOIe8qBsnQEJH9rvgCMWmiSi7YYseR9t3pKIH
BkjmOYn9BnRcsLQHK31YISFqtCwXOm3LAw52dIpbxOR7WdGGTuZoLzSWuOdn
WG5OzYNvRDdYQp7WpudaUGMB0HzNXHK1WfdLw6arzFZ84QmcPBILyKljdAmw
w+S2SpHDKxtRZF54U4D7f3NrL3I2N2M/yD/7V+4+QHm0ksQubaClkwVuPImL
kQGCA48bAumKfM0mVriZqxxDbmTfKyxtN1rsTBZEK7Vp+5u5UUCF2BOZmaZR
HNDWM3yLXMjPRrAhMPeA5d8g+4cihOhjBZ8srWU0s8gNgorO8t8I00m/gbcl
WCLydyO1HsxL4iY9Gp1j7uN5M0kyX66/y8wjf2GRhcv5waRlQY4CNNBXsu49
M81IsuRA2/ylJ1uGv1qViSPsHUAQP/0STnHl50G4D0piJ7dIv1DrtlfkRZ+B
X3g+sbmyKs1vWFVESR1FhrTEjyyjFqXM3V71GxWSYVs4Qak3rROXGwl8Q4Wf
G9mOdnb8kveZR4Ustqky4p6XTwj1qUxJOLGWjpU8PQU7JMMg08Ht8prF80FI
Ki9S2TgT9XQyZiwsiiZGlvVVVaiH/Mcygtf7iT3zg2/jWlDwMu905Ls6FpCE
XV/dRb7igHRsSSobR3xoWp+wN4biqaiAgF6YM4JLDUGxXhplh6Jdl1e6orjO
gQ9fC63LaEBgl+N0fw8/XhB5Qs4VRS6GjlJaf7mCBa+llm0fqRrNJ74PmPDr
ZbAsafaoIrKtFx3bedD0Ug7boawKlRhkwapPe0OGpaLI6LdU5jh5nDnIcKgQ
yI5K5YehDIemAikskZjwFPwDFb826qOI66gp9PTzagNFUuaJ1YYMHWCfTJuk
Apt1pCvHa/swuVJqBKW3jO4F4iWtd7NqHMG6re+vBqqmMAxDgfYB+DeVXxI1
+x/5DhagoV+zA0VH/ie2FRVdWqqVbJyYMOtBBQaif1iJiU49An+hXL0c/t4l
ROCKcNIaUyegIu6G1quGlUnbNmDcv97QFwZoQVIVr1nQXlbR15Ox5gTxWNYk
bb4M+hFoRH+KAaftPBSeIunJWNx2nB+Gmmt7htqNDThuXVPudf6zZKV39Pox
phyvq3rG/FVdjBQ0I0yxMArhDMm4w+SSdufKF50Ug+nThip+rpFp1yFxsOn8
Vrew+B4CxIlVXpMfRckHxIMp6AcjohiIPLKwahQYzy4VEoLGNgrOH1vEx6+D
Ia2XZeXs5J7X2W5FqaheLheWo9WhkWq9vlW2KbW/13VaVX0CKlHi9nSY8+d3
Ni8mzvN80Hd/I44R70Zf9SgAuifdwxhK8v4IVp4tIQtjynF8UpqP3KfxQ9Bl
vm2bCAqII9lvKU5EDibQH91Lqia3Vd563sDrASTz/x6iumLnG1byJKHvn9RM
RaF4mZQ6a7gKdZ+RWH2FC4yiNPvThJOWQ3qiYb5yd0wfqk0vUr8f2sm0QY4K
t8yunSfbStSuENAIoDLpB6HQyDnKC8kdONRN0+ahAeFAahYLMGloOlbUkIRD
a/Pe0iTcEFckvTkXvPkC/3Y3/vaysCwJpy3w5MiKSzXWFcWtjGzfyoWT5Jiv
t2UoOVr2PSxs/bXsAOhgVB8S3BTPmJ4qvi79KI6oKJQJM5IwWIA2xL5eVDy1
7xs/5dCbK7eRd54Vxikj0RvABeXhciggEMN8QTQAcZK4PL4MX3djAvDJ69F4
Mj5bpqwuPpg9nlgmoRkZzB7cspGOS/gvxpsYDFZj7Fj5JeQWasBnLjCwn620
zF31+xRMo0YMQFrZuKF1dMDA/4LnagpzfKI2blu3uqqINKLi9+UEv4EG0Yeg
v+ns0rxppuEKyQ7ZgwOscFoQ5n2mgn+jftpT5NraDkBRAyGF4xGktv75f+6r
I+Zmu5ZJJJr0puPiPQ5n3AH3vZLkDEq4vLWY2lrqUMrpQ17kyAVOQVDi3O6a
ijmOxkfa4TNCQ33eR62WGsQcnsK6I5zTy5otu6HGyAYWrggnQBqkgy95HK+H
u+E+6woIPdJSsmG+5XNTngKlAx2muQI2Oi5U3QYn1ZYB4oR1jJL63NdrDehE
AfaeNpxsCxIzbbMFTr5hCd4NcEdcnApJs98HEOHXgEWf+WKyyA4ihYucZaUM
yVkqPuQdYBdBzXwSsT8TH9iXH0yLEB4KkG6kauuVY49YJSbyb3+GfD5f7C7q
cPvw98eKbXVlyVaDe7qVNgVSurTg1Ev8p+3dJpvAHqsKpYqm5EoaUS5aXRd3
7CHAV22gi59+sLoy0Ht+rjA3btN8UbrIJVjcJ4Bs6xfrSOj4zsRfA3RvXSbp
MNtfVA3sFoMyx8bq3D08ubLpmdt/WqgcioAQvE8Y0rPg8VUMHI2Q8BukN5DC
kE3zDzYrrh5/LcUuMorewXLfgFNTbO6lkH5FHpZrUWLC8YZPZB9+VTzTvaxu
gIRvsGcch1kGmaI125y/xt8DHLgISGBxBZnjAVCe9xwPyPWjDzFlIslmSMgZ
8wELt/mio62LwFflXAp/X8qHGAjPyR205r+5uxRHexvE6wOyh07IMs9Ewewk
rSrVqjyGszT1YCWGwO55CQRwJnstRz9LZyGAdNdiyhNcYzfzmVEW2onS8Q1z
JTjE13AlyQeqojlKgUDsAp9OM2ub5RCgV09ykC+aFGUs10D5VodgzR2LN6lS
nRlrYQOW7GIGv8mBXofqf29myNutqO/wLRBb4qyJp1Tnja8zTvGGHui/YPA3
M+LqVc5VhfzGYPn9oDUEf0J1xN4FIeJlkE01tqMVmJsDtAE6NcKk+3ZG8aDu
IYNjxf92Vn0p49zlruUGB5/mACnj4TVlFSTyTPqhIrQwMGojYU7PDQveUgUJ
odDZ0qoqc+ZD0F3kcWVxgJHJY0058jNHzhEyzx0BrOJs/puGeMXWlNvwpQTg
XPbQv3fwlkWJovRzrH+O2inO6kx2whioq1lnvRvpnfYHVCfgTGf0E4nGssSH
ILg9LrKGhfohI2aUBhT5O8fVSldyhlhq0tmZ6tyXzRE0L2jqURoROi7GIxF/
lMOd8m+NKmvT4hR8jD/vKykTTff5mmD6iIX4CESjuIsxBDsM+RBbapcEbBAX
NvIYyLHWNGnqT/XgqAl+1VNYHhORvgosCypaYhquyKENw1g3dZiOWGQ6JKG8
9m9a+OPq2eSY556mYjBDeWfRfL/BMgKKX36nggsmo/lLH0NlWVFlqob8xQuy
2dyQMvDW3BF0Nk3JGIi2lC+OYOfLHvWSwTx4FeF1hAWTgLGIoW/7XMXbWDJ9
V9HA7U7issJYgLrZvbc+FCXuD/eEXcHq3lRydBj/e8jNTWT6KEDCTa0678PU
HHiVVeoyM+2sJqUpAGCOaaY+aYotbJNiETfuRQFD9MRVFIvL6iZo+jTBtevu
Q11bRZlta8w6BDUhwyy/ppAAUt92tNGKrqXtC9IqRXKQkiIG2Yv5k/ZdUK37
g7h9Hncv74rkzejOZqhyZZonxe4+mEJG8lD3eRgUr34Xm/wB1mzkxloxVrSt
/T9LumJMvhplbRNTXlpZerrt0+Au2qehRSBfHFNhSkaBdu0VZ0EAUp+zkjjd
r7TSDmSOlxEUxtGEHb7Q4WDEEN3f1utFNEIB/NP0NmGxTj26C+NPPY+03DHT
ILcBNlvyOnMdmLQxRu9ohnjLRrOMtkltn5NHQKLWGmyZ9ubQmDXfz+AFg87D
2qGNpcZ8IICbtqkiBqzwgAXXNoxo1KjXUsmgD1bJH+vEJPNmMSqP6p1i91Pf
SKej5iYe1LStwSCrfPVHIS1gd8dpy19FuwivUm7jXmZtWQJ9SFVWW56Dn9sN
XUQGjMwiM1ptfpkh0H8rRwjqzxNO5Rnw6RY8ILAqronU/tUWZa0HSfP2EF5o
0LeFB+JDjo44A+qXdtcadg+ve6F30/rqViK5JpctKG7mRRfauQVs8v1itngK
oGO1G+FM3TL4DagEh1Gd6xXDygGl5UlrRJVHhq5DYh281R0yPMThmatBeSdI
snloWmjK0c7E+3iNF+xqCearLzq/acdc/7Jt7hXCQ1hXeq4wHQCrSHp5MELt
dCKaXQ6VBfOF44rQaeob7daBZNaWU/rxhm93mzgRTjWsmla+ylORx8LjMff8
97RhBjVswdGByP4gcsla7YhOXX4Tu4HY1jAW7SRYWApPjhStsNzOpPgTxR54
E+AzjneFPafD0q+q5WyF0RyznWw0BiADFTMd3mPYuBDBdb3+VEHilZaMradA
rPpXYNrXKttqooT5cLAfdfKBGBDWi1LRXMq6xfMgzJrkhyEUyrccCiDop63K
v66MTHEH64doMp/m9wSHUWMEg2SGgDUUNhlrbRDGcgH2Dw0cGUpf/ouefl96
aCLQpxclT8dxUwApneSC7/1CNV0J7MzvfCoACi7H5dp41RiBw6AO1Pa3O2Wt
Xr+iIrCNC+9j++1C6vsclxYG0dngXhJeILcASYi0AegLDaRm1PnV5AlIweEc
RbV2V5Jez3a6R99T+fzRWj5j8GLx+rAbLtBsGKTMJb6SMTxLTGKK1ztP+Gsf
hvdq3+G1g7Hgvamy/KFuibrFWa16M4q/mmWm/pG9p2fpASUeSBhX6pU1uGTN
hd5lD5SKlDqMAtyd+g9EvU9v+L98PURc0inwTPJThUKNyY8VxfnRXWT8IGNa
fClGvIBLeyNEQTktwJB+RoeL71eh79Q+rUDJNJSoR2195PH9n4gp4sOOLfvv
N/su70BSJETvNBv0hFFTZcZHqrDdMhRlVterk0aUXc5k9nzdjKotPoV32xI/
63qLUBUaJNL6qY9ZiyVdZ9Z85HmwhMAtuUDm5kjEL8UYYorJOCI7sj5Ch+D4
ImcIixf3EqWhO6m6VigYwK5qE1loAOluZ+pQNi+XXHjldkR6BpyDW0xdHVLm
SmtzC3CVOEJap9l9R/8iJgIhAY0ZzcGt/+X8U+uo/3Uej/CU2HAvrUo1EGz3
5bj7JjPE+sN4+47lAyMcK4wZe1WMoXMYzdj67M7WxgOZ4Y8DVJjpmVgbwHDo
X6/CDQzsLtJ3yIoSy9QqzN0pakFghW5nkoBNPwXwWuEYGyoYo9fcfwsLZqQZ
w5ggxbXAi69w2/zz7fIn9nltY5mnB3uxV0kn0N0AfPqANMMjBxEbFHG4O4LO
/NzZgMEMFazodMxqm+Du+yzdHBQy4dUzfR7hMVNlvYlys2wHo2ULQDuuHGQI
Z/LcvFGWkgO2gIHlZE/OugHbDqhoGyonbGOyJHtSkLDT/lOu7ym8gmyJDVAv
Pe9xLrqcUuaAYVc4/Bcq9GNf70/PB4yznUhjaa5yUGepqSQ3M/ufPuvPDwo3
ik5s5LhB1zdCh5rNpScBrQPEtE+VtgEs8mDKTf3QrVNc+n9r1YQ/POOUKIDj
P7yrr6SZKlAo2ggOvDNoNdzviEb1CO++FKkjd+dAGWCIwBTEiDmUTewiF4Tn
m/VyQSk5pU8P2NCgwR1CA8lf4RFTZ3vuj0fHXy/jkldpJzUTSJvtMCqKS8rb
v/BgKtEdnCZ9tmMcT6nxLZERh1erVzKWNsNx8kvP733F65IcoPFx34+vzPzM
pKebbG6K03ivo2yjeMIUl7t+qTgyII6/sISHlZUnFmP82/VF4bVunSlx3/zu
K8SHJsHES52/bNBHpLM7R9CZ/VWQG71dOkI0MZWLbeTL3sBswcctY2APdP3P
mHufT1aEgSm6KNAa4XValtkyatEpYGvB9pJ3z8Ri+Pq8nye9k9sSuZzTUgEN
0OP8qEpjZOprby60TE4HVmh6eBXMfKWaQWD3fbh7FdGjSqDP/Qf9SDADl7z4
SQdu5x5X9c83RxODRVtAVf+3z2BqqhStGLZsqqtQvbRThfsRv5CfDhoad8Q7
HepMLoK/R4MyyXgRGssHT+zqveMhs/FEelcT8AwfrZMxIM4r+trcvot/MWSI
hScaChSwRWD0smmphiYd3tjRNeV7sVayMUI5OoswGP6hRK88oRf18IBTGxd9
TvYFGLnA32NKcg0iqxHXPD58U/Kqhowcbyd/Om9gPfVCWVmuQiCLIJr9vGRZ
87LyjhtYw7Rnqs/13xTtuRDnMJVXh+VFlqdkrPk1h1VRExwa88UNDoDmkXj5
/nf0zX0I1NVVniXAr9OKDDN5gZ5gZAdWiThSB1RO6vgostHiG+zk8AVv5ub8
5lJ6Qek1WLjIvnPhZ+UfCcxl1tMtyXAyoCnhBvQnjrL7FXwA+skTT5L+R8TJ
jZheL9gc8kGilE+OrrFl4c0vY9VFzqEXF4/rfA5X56rKrBOu3AvNY3o50Iyb
sjF9noK7MEfhxaMZNZ5LWslicUfQw6ORHTCd1Lqiz19kpTBsYl5dxMJoYDgs
fpEVNfEtvi7pEpPqzzR1ukNBZGJId81gZUrU+DSrmblbdlKa04aOCNBsPx8f
9Zl18bl+F3zMGsYqzURLivGQegz/NS8CGCKTqnVODw4Xxk42Y6wKZF+q+Alb
S8MLX5ZPZN+0ZVPJqoo/kUa2xSKqSPV3KPnFLLa1MmyvS9Mz//SzLmxsQ2SI
M+JkIsweGU5ZkvJdLw06Fj5YcLwPSKriY89rbvWHm0H+gIpoXoN0qAqS5f9y
RmurW+ax10pGVyvkmnBWb5+0Alrcrlyt0MUB5FxJlb6XPyADyYlTN8CQRrr/
kQOPBLZi1NuJrsZxGkYcbhatb+rF+G4ffcxSzCHR3A6yp5NAtX2w2d0gTB9z
pfnq6sgRRSotf17DLLQqBZyv35toSffgZCovs+5WobWstnTeKxIEpjavrAFB
D30O4brpjUihb6na/E5W1CiaB3InyiSGX9OjYulAf/BKnmyKfuTko4nxgZkD
edMMF3Q/VjS9rkIU2JApuFQNwSMUR5mfTWGAWz+s9k5YdErgVOIcjCdjOsEh
XGPUzEGqiKTa+ZDJJzCH005AjAeu7iFtpZ01icagRV8XGy9+jGBW6YMfDQwJ
2XGQ9rd3Ehf+hcrMvJRHmsmw/1oG2FbkERYDzyA4Fws3zirOuokDADgH4fba
X3jomo6+5b111NhnymlFfeWpxs2LSlQggx3zPP4m+PqVzgiB5P6qJDwVvBqQ
6TW1zEzaLsNF3J5yRFe+oOL0LKvPKEauNCUPAUoRld4CADbUAslboixYGGDP
M8JfMWZMqJX9Y7lXRkMDlD6LFOvqgnR+8giJOSUia+ldtpj4irMoZilmhj2K
h1k9IU27GafI3kZvWvZX8kaioQATsXZCOOh/UPvEJRWI4gr595NnMBIn8yB8
P/mBLEo4HtQfsi5xgkNHH+RG71PeGw/OiWTvKKBZgkE/gGuDBuy/C+l6iIKz
58e5jFLrqiBmdgZTteVJyL5OrkryOhhK1yqyHqSnI0VL14zm+GDST0QhmKRy
39kO2gmSy5VMbdjJhpshmiTBGIew7KAnmCRgx+qSI+kW73sd8j0WWvCYQT5r
AhlhcLSks0agKMsnd8tkQJGtdYXnz4YVIgHIidyBzhw3TYdtTOFNKCuM7iLA
E1WWeafPr4Vdk/OvRZ+f/GBWBre72jXCll7vPHEf79oOPuA9TC8iHwckLOVm
Hbhng950gUf0MBYKpxiVtuMXcbZckAYhbbc4iZ0n+KrmsBsCTVX2J7gybvSS
N3/1mcPvexFowUS4yd7JNfFQcpgwDpSVcRO38LCDgPxsOp/bAIYwtcMiu7Ui
42Izo1OyW99ABkt4TnYAgRJ5gLryDuyQpLnhM0hcb8dpsltzX/NTrVPIusyG
sCZ8pGBMEgXvZcwVIKM0FW2MhLS+Q5tRWsBYCsaOMXb2U9YeiZ2c6zOGturC
XiKvFZfFpi9zloi7Y70jdMx8HfN3C+Jlmm24GZfE7wDjA9VeIYson+v8F589
EkeeRtkoGmQR8ndox2sSb/pZD83rKa1aVv/SqRA1o0KzU7ei10FUxJSzdfTU
fXssu5TnZ5AyPRI/mW81/gqb7iZTwl/0GKiPmUlboyrI5ONRxpuYPBQ2q1F9
q+Al0zVir87qfqnWLKx9wPMvzD/g61uG319sqZ1aDuHX7mYWaiCfYT50KF8I
RRJ5bXcVsa6yl69EEXYRG9QSULkBJqsIPfGTk292EMSl8dLD7/rEII0pSNRh
Q3QPoV574cS7c3GFsCF49+xxHH2LsXpumph3GdX5I2Y4YO9Q3tsx6L23JMiB
llamEJ212NQb7Mvsg/CFwrWGwOvV10s8vuXoEYtaZZbbAgjV3OjP/kn/XRLy
cUd0d1h5kEKSkc0wium5wjC0kStUcSio58aFcX97OKIE/OA0+rU8dsUr+BWb
2hKpyh4baskxVzoTrLj16xTDHdaAqjH5qcuRE0VthK1U0jXGZiXz/TLAfYao
PhOF7IcB7leANDJUZgfMf81eZRcjEUzXwgdk3uJLa7uKiqI8wz9J/gLZeG4v
dkjc9hsMT3FE7n3DmLRuLB4LBw0ytqX5Uw5q4sihVBy7JlppRL/8BSXcC28H
1njY2YZP46vXJeFhnCnlEncEAP6xPbxPQ//jEaLNSgbxSX4UTbo/xaB1H64Y
sLQd1aRb1K8f03qXtOWcmSPwXIMz3OL/b52FAfiI7VRe2mfrIDKXMaHoGVGR
eyl/K8xPfMsBK9PUETqsCFbl2To/pqcOaBHt2tjgoJ1VJxQRtNS1mbMGZTLC
L3NPHhNjbDDKx/+AWj7FTd1G5SWVpCYOAb677TSNjX9+fCziS+phG1y2gHPR
4wPiecaPg/JWHssXgdZwubOzZR5/OFno8QlgFv9Ah1F5CpYo9O6I8H6CCLUV
0E32S03yOOm1R7TW/W/WDKkbHZKSWsMDkPCR8C7AIyMPuThtXOWCkxLLLWcL
5ac6rPnMFFv38ExMCwcBus/iEYnbEPhZLjw2kvlTqWM5vjHq0O2zkybzaX1x
Ll/40WQYmVW49nG7N1An19mdSY7cJKKHBuN3Z2sG6j6VKZAhvmwArComHnt8
HGPoH8aicmulo9GrdjoHs5cClk9NP5sq6kb81OgvUZLYm1fQOWYlUDEl9XIP
5NMTXrb4yuKfWFMcpeZnjbjyPHlbI1ncEAFWp2JsjvqRZ7nfauwn9x0cXJzl
Eh2ixHZNM5tr4MRCJ9/e7QqwMX6tRPufSGIYgD3GQmvooFQwihtaKERxW+LZ
MQKrwele10QT8L+kRd4uHKwOTw0xms265XUM3ylNB/g/KlxRLO3KUH7iq7Vj
hgje1rx880QIoPUynNZjYRmmE8JOAh9j0GL63IixICL3XUK1pIQ4M4AkNd3F
2zOLw2y+CntYDFZE1V+9xGOgpO+KM/MalE+vJ4XjXDPr3pnxoCekGQ7ZSC51
jbNawgU1p+Ivmy0ML9GshVZoYYh896aoblX8borKPjk0RIjMArX2glRwqHec
BV07AoF3Mn+ro1+5MzXCraTQBawpDER2fjNcnziTL/xO9ma0kDmW7obAyko5
k8NF6V2ZtkqVo89rOlkjRa1TiuE4nd1QL0/nwv5YthnB9hvgdUmydw8y8alm
0NGZfaCRXPPsBWBWkLKLjYH3R9BaawTDCnKoinxcIa8IPhEzf9BFB2GEM5R8
GB1cuAq4mqK9dy3qn+1K9jKyQAx3XQKRsK7rMPHS2mzqtVjOt3SkAFGeP+wi
swuMMmv0OQ1rkob1WQy15pRkPNE2aDx32qV8Mo9zV9OiPzWSTY+LKgEGLpxS
pbzLQU58IX24wR71CdwzTtOtR4N9BGLaTNRmiXEO8X8ak+/VbzIwFws1HTuh
sieAEmw/OHEgX2I7wacEEt8hbw/v3Uo0HqzqbhDpepKx0evPuSmc4MeoarPe
jhZQTLMuL+PvC99iSb2gymdUeY9cdFSa9pZzOX5ds0AGROZLPW47uD0Rt0Rm
ZydilqbgAjG7rgv2v1LgdiXlnNR8tHzD1DIwPLmTrv+gpgadicC8IYfgOzVR
jatrm/ONjTRNQ6E+mYK5gGVu0Rn5MKPxmbxNr3DztxmAOOVZmE1OHW8N3IyE
FSIqO+Jc8kKVMyrOkdkJbT3Q0OJED4JZgCXuQSROQO9vPRYvlMZql7THJBEc
EXotzlQHYiNyPcOzBh6AnZVXGnMyRHqmj3zEZ20qIRA6k8M9zqnros46CbwS
hbe+eTyS7BrA9Yde+bmaty9x3T6M8mbDDkv0bCwZp9eOs1wZwtS0dfAZ2b+3
ZyGUClVBzIwKQw99SeMBcJPR2jwtZUVoDoX7TV5Yk82j4s/pNOq15zBV2yzk
i5fxlPTj6Ab+n7efEuaBgujQX8+Q+7Lu4uLFmIvQUxscT1KL1LCFVkMM8hgL
yi111fA3X1+9Xr7NpGM1U22WsSFmBNwJqw0szsS/G9C+tc1Rd+9yxqkXBLAK
ihBc6NMjfOHZZM5Li5ZztxXVP9hFYuOTFVoYCOSRTkdMXgLZImuMjvBG60HZ
idc4SovQAsfICODcFIHkuAuJ6HC3vjgEbFG1DtAzP7FGrgRXS06Htcj0dRki
O/+MXXd82Er5gPLKcx/vHwBIZWhdQXPNYoqxVWsux+JNJ8PELpb8DgIGnzqK
iqW3JbvazeWRKjs5n012OPOsGB1lg0FiU0z5aqIxSPEzhsNnEW5pvM5LMz50
kSJXJAuszMz/z9l42J1REjKo3k/bctAyXCDUFebEIJK8Y8FMGul++EgZfrSD
1JyW0rfX4Esln6eCnnLDWFAzKg6i220pMbxKv1KHETOkD6AkI4V3w2k9a2MB
znSCBQuPUxN0sGX20eZ4jlJOPBKisigyO2xMLU2SYkM5w+A5CYMaQ3r27e/L
j6aQQzt6Imt8B1VAc8jnwD6NZvvv0h/5JpxLd9ml6z0Dc6PsHIXlDEYbCGPe
s2mlQy3Cxk3ELnl7GorBJzS9r4HgBiG5/z4QOdh3X/vFUbf7tYyvLhF3Gian
3JSoF9BSJGvbFphAyGL5vOYenQHZJqTYRD3QHXL/aLj293RrzuPMO/EvrR0p
Z4cIwlUk5GJj+ceInwzQOs6UrX5Upp1bfnwYg9+QbPhdzYK84V3TTACGdQ+3
ET8nYNTerLQ69iW2s6XT/BQF/0creDf8xTFyIQOdA2FOXs1Lfm9SvJGCI8Gi
LTpz9oMC4bnfCLQ7b12nJmLm86zW6ugQOXMnP7o2WrpSPqyDTKT2bPvJeTXY
kMj+MMm7uz+v/IPPTmOEGxd6xB8gMDgPox9vVWEUCt6lmfaKqlCxqY1oy1e3
QPyFfa6Kk+0MicAYhjJmRn54Ewkr6xucq4Jn9epb7vTXT3AaBw863KFkgrQF
QsqXRnQCGAbNGLjBZh8xXEzk/gcNdGVfNiro1ej9F5y5/Te9VrY6FJp6D4JK
R7wf0HnKI9lVCiT8XaOgjiBEMcSfVZk9GxzUA0BOXDhJwtv9xWGxZuH2ij77
qFmcCwCSM6sRJTgjzCg5zU7iUsYIMoXLIjw/K1h83rxR1/38ytebUHzONz77
Z2ATdV1Szcs614Z3ZeSBFYSt02/Mrf//+Ts/OhTsde7bTREO2wthSFKvh/WF
wb0BFsODk91zR2gdrfDGMT4eJ1tWFrAnK0Y0SiiW1eFPo/lVSoEHxWU16IvT
wE6Jq8lfrZ2AVGzYJCLSTwNdk35GVoTW+GpDgPp4uzYZQJ8iBSVazkXWkGnk
P/0ABgCarfJ+67JwRF1dvOzQwIaL7dmmU5tQ08kG6qCFkxorErEEW+0KdIkw
zjR66I0fCLA2wWb9dgPzxVdWQw6N6CZz9gBl1eCd3T5YqUZaWyQaDwJBIKG9
0W3qdtnCn9Ji1/vvuvR8pfHLwN6zBYu8RShYWkTqy+q6wRcHE0j09M2qupk1
Lpaoc2ZR5NEJTZsz5SK1lAfH2fWslE0jS4uuUm4lKFw97pDPTZTpKZqlKRZ8
XwZ7BtL9zOjcYPYO0lLqBW2OBhpe97RFinGOn/cmnLKaVivIs9xDffXpEJC7
av0htqlkNnbmtkb8AbqZGeMZyyKRzVMaKze492cAFEWfXG48LZOz1RWpVigE
4VctU2UT8FX3KzcK7BA/nJ3DV3ZWz26VYtA1MUMXybUZh1OBJwpOyYCZ54ZG
swXvKfMlkYhXoyDiNN4wAj0we61NqekqqPu0yTykeBtmpM8TbqOlemXTlobl
XXZn5rdb3upqK52UjVN9R8S6KeDT0l0/LNQOz+w9eBcsMalRC0eAA+RdGc7D
fnBPenO8HOUawZcKbk5ealBhKXau0vLHOWOslmNaECXZcpBiYtrQpSLCZVJC
dmVeD3wB6fVE+BqE62IXXHKVun6Hj9AaD0cbJbiHDLoTOL4Rw1tDrPcdyA7z
n8jtmKMkxe9b8icRb2IoVhxHe4kDllySpLAxTFBHIHDwE8yPDGYfu17+VIk8
zR4KQqgUGG5mb25OYh/kUYGXRv2n/r6ciHHAYT9vBudcEy5xbBD5lnMeUC8q
2ISAelvmmKmjvxSK+QI2EwpQiIa7a6yO5adgZ3QK+JPW2qq650XSMvEn1f+r
tgjFOYwKEQNUxjNgICp7sq0jN85vOEKqSvqOPOnll75JFExBctaYwMAk6CAF
UaCmQSiWlXo7Dmt20Be9ceyv3r6RQ3PY+Qw8xV++dZw+4mpr5RZNmx0Sh7yX
IHBUCPCWths8SzQm0kLH5wiH8UCzS/D27TNpZCNrs2AXraNx4RICkJ7V2dqf
Qfy0H/ElIhInx/k7wwwsLEdDh7uQs+QmeVewJC47bjGn7TVJGeYbOBOnNB1L
WdW4Lg13Tp/smscKmQ4EOdLSi2GjiAjVZNmnMlDB6nD41hVQI457+FLGDtY0
TKevjD/hCqMs38T2bexrpPOkeEEmrTwYZHRc3bF8P7bi1dosmCPAkZbckmkS
0jzlTvhi0pwEfxjbg1I9kO+lK2N3AU8iTcSG/3zNCVTUWsOnJpRmuFjx1v5m
V++s03o5At28ZdkOhHB8ISrWDsFyCA5bSCuLLvjcU00PvFvwB08xgXo3eL+X
gHJL8M+UnWe6JiCwqbAF2LLVsLN8EXXElHJxV247DveFRN+q+EVzzF5Ln7pm
HU56I4sMX/JiNc3IR0I8Q4tm3prbSEuk8PMf+CQUA3yo657ChjwyyAOrUfw2
pnGfRXiHLbfDZYRPSnO1YD5fitp4MF+fhGGIx1fiZbUU31UPt8f2Mn6bw4XA
IHoiUAOo6ZEPOm/g2UAObfayD72aJGgIVYkeP9jGX6eokPn8UhJQTeN3SYOC
44ZUOi58xTasNaGNznds3tyXRfT6jYQ3pbitv7Oj/gTVbQG+FqVgYReTZVUb
B5s5eMZS/KawmHvIKx6I4yBrXHOiRuQk/K74B5P1ltg7Q+kUgdilDR/x0n1I
FBLeJ1UkaOo8bZLhw0z055xlWxF3xWoYC/O9EIvdiHUI3P9Mct8haPanUU4t
3ELtWDV5ZhqPBomB4DTJ/+wdh/dLhxqIeds6HexxeWowA/Xy1ZlEQrqbHSv3
BNVneNkAS34xi11hFyQ2dB+AW1kByK/UTxOyc4rmVdZlMZQ/8uXRXiNVMAR7
mM/6D4isbGw3dvPSM2hAfJ2W1h3Lpnct5EdGrP+JoY9C3alK9PBfQra5VOiy
+e/W7e5GmE25pLH57j7x7la5Zvfu9hgWtLr7pHxmFAL9xHJR94fVoLH77Rik
10JfAlHrPZvxjFsprmhbes+lB/q45+1kZCqpnxZW3BHHbPrJO00iTeD5lVMD
22eQRgGDGyK8qWOFXdwRu+81qkevgCmfnUp7WQUdXuGFrdKqrfQ+4iPm+tYP
OWLWeohc5zeyWlS9mRTQ2xa0X/Thv9s25ty3s2POu0P44VQeo1AY+uD2z45k
LuX2VgPPhG+xrluvW+lBW3XICI6gZtRhJHaq4bjXSvJ1BWsUxkbIGh9oR64n
VnBbyNcWUloSOAwu5IjRgEf6qRKHeAgH3m5sea0UXUvvEcLKLagUv2dO9/B8
tobqEweN/7EGpgnSPr51nudaAFyXyKOof7wXlu/3bP0TPfGavNIJKk5dQH7c
xTm2vh/x/qjQFvU3zjS1YdjqdnMKhpcOAUsgaTzcWIk4ulRh620vu/8sglvN
cnA46RD3ZZYOQpy34quUux4oGrxx8I9yrdvqzX6S6EYLZNNg6mAE/2k9mEPL
Ar8J3zno0QfOEr/e3Zk8vQbfAQeXz+d+3xARForzec6tnApdFo2c1jA1+wGw
0h/z51KBn3h2e1vdKqiTQ603Zt83MR0gzBvJN06vfLE33DlKpZH7iU0WNct7
X+qDxt0DNo2TYJdTbM0JV58D147omXtVMPbPFF/qosK7fpmQWflFMiFXUBbg
Vppcj3Sdy9m6fMVYySRdMzueZaWaElOe2cQfjI8pRwHxAXZF6d3LdFjtuJxq
A+7Yx8qJb8CVyLEA/d+FfJJHkrJN5ALPJszK+WJ/qat2jruJC66IVEf+VEnf
Gl6s12An9Y7WJegc3sfX003f6BmYoDNBQtnToI1NLcB6X6CjWkgYGUnEjiKY
mREKeiqe+37OpGxBor3JCWWz/nqKsqvrewJwrEukGZgzKycocgf+nllU/Hka
SCt6uuPL3t3vChB2WSdkqy06FVb37xTBmp5MWbIozG42UgP2ZtkzSuwqCgae
yAQxcdHSF6/upgYC1MejXY+hJmmndfrXjPfzPIrCllZJpF8gba5LnRSasXan
VCgslvvv04x6dmcwR+SBqquNwgcvGxqGkJNZgDtVMrZfZMATWBt/MFgEgE2h
5+DbWxCk9HEcNbbyeTBYQ+Og3B9MRCEDNiOdeiQyh2HjNztW8uk4tZVaQW5p
VAbx1BCX+YVtfaZt3mjGmuPGw9wF2mf6SivfgnhLVKOsJnVTBCMQMJXWqbvL
wDAjWJCmX5jM2ZsW7mvO2bVOn7AiFe3yEzBbsTg1NKeR+z7KwbZuJqmOM+q2
9o4N5LFE+FCOjlVhlOEF2iyJlXUcofGMgHZGtDLVVWKTvBys7bOaM/NzgXw9
sq8jJGSuyDgSy1zg9mM7uS+tQFWyH1lc9Y7pMktmBAYumgc5VZxwXNWHHs37
h8CDbq9XntSiNFPwbFln3tzqJvRdoYgcU0S8cVfK0xP0J7Q2kkacglYYzSef
m0sfgF+tu8iw2MUroxOXcL8snTu+pcB5UHscw7q+oRP98glsItNeNVL1GIW4
GaJD0/L9PLNBqHgcuXG/WF59BqMIibtz9KEvdaz7LtGuxa3HPM/HqU0XntUI
2exGVa9vL8XCCEneJ3jgi8FBkVp5y8AnYDpfNQZZ6oBXEGQzDgcOWjaCo+7W
py7kYv1ZmQ+p92euhv1IiaxtFMDXZYjtjB9Jo3Ps8ZuimRITFB8Q+K3HEpD4
NekpzEYpcmauzllk7rgrbMMZl+G+6cpz08ykgjSeRy0K7XlstXf3RT8kTwxw
5u5qDyek43NLy7AEAo06jaf5BP22cnAvdPxY11glNbNziwXprj9ZmDqYaSab
VeoUDz4O+XkwgryfiuXnX3sysjXlnYXtGp8cS9wCrtIWrn5ztln2Uo4IkrFm
+qCmfJDP6vdFiTUO2E3Y80ZuhL/ylzeh6rmoEvVNdIL4w/fpecyeR/90rz+W
aeQqyMK5Cq5NwIUABjSg1QHf5weSv5lvw+vgXpDhDSbywtz5fDKpXgmdl7eJ
FGzkNDVN5LF82yItxxR/8Dq6w5GOEkL/C4Nh5Plq01ZtBixo6a60DnSl1D3e
mRUfxmUeXgvTS1TgWs/74LAmG5IOxJ7P76egZCeYfgtOyVvkTwYf8tlP7kie
/1DnbLmsEwzUOsR86I25h4ILRzZY3011XkE4RGHJwGw57B4sbdcl0/lirgST
EF1GZtfmxjTVT5+O+wjg2J+qpwbEJzmJXV90u3KeWCoK/FL54RnDBRGk9G6q
tS7Up3qBYptCkU1GwKY793jOK6Wx1qNP6WCtHOBjzlKJTuP+DCND5XzRhDg3
MgBgKoWm4BQffBYdTt0PnXPPDNk8SrwOsZA738D6ki8e2a9xeGtY7QWUui52
gjk/lUupvrduQUmtGl7SbnkdQZBWqhfsYDdUIFQsQS3l5WMouuHArtivI2oX
A47JSuRNaOpZlvC3ZWb0RHZVUg+wsAwqbMklrmKDqG1asSjO4aX7/x47UJdG
yV75kA9eiyyDZkLahvxEfQ2ALVykRZyk2BYnS1FocPU8c1Ja2u1H3fR2yY6E
4rclYJQPYx51jtnDv5hX5KZ/faTWOoG57fZQ0DsdiZWI1xQQY7N1VPOzIQRR
AampkSYkiZwGgim4GwyPH9+VrAINcc22FpJXnl5RhUUDeSFgxn8vmxwFBOMJ
8fhkxvBuMElCcmVALv7R9tPF+urQsfKc//vab+aFStMXniglcyPSUuDvERrp
U3/VzVKLz1ju0DRCa4jeI6iXewe5uoShDWiQSANqqvJHZrASlRcA//g/xIJn
3dLz+SWRURyS5BOrZ/Xwi+pxJOfZPDWRn1NcZSqg6f23Ud0pujMa2XAC1jz/
YHdSFXNUGJVD3Nbd/Y/u5Zdd4YYF4V+PMlX3z34u0xqMiz1BUo2z6eSgj93l
3+Kf8ApPg4Z08DrkFBYeS947b0tU5Kdk/rrzgVbgFpjWjiWY14+ggx7BBBRr
kKo6vIiuUe6OH4JCtNj4xbpZ3EAknwj3YbYnpDrh5MPW3bQumtXI4CwuuIjL
qpS7A3JEo5DVmfdK0qqQ55EBl7IeJmkJ+ahcf5xIbPP3BLFtgKH8PRDwW7Q3
cwt/Uqe07Mo9iLGRjJaI3qZCIc4ezkcFYLVXqWKdEridoGsrO0gjJ0Zubyd3
ccciTAk5w0Xdp2NzAreGiwxiHHRmhqWz+xjYhdv55xXn62Tdb6MsL11lDNhK
EdaDuwjlvuPwmwKYQYVhJ9QYtLhyiutQnV7m/HLP/7F2rTV3QyesM6tPbk2w
yBcCbqTUIzxmLMwmLTL2WtSbKE3q6LO4JNeBYIgqC/RcukhODov/9lxjjyiM
sDvVp7yvF4buq/0qgZ9wI5to4TMRkJzEplrgtqydOtLBWHtuanyRDF8Av14S
trvtAcRkFlR1MsiP9HJhkek//g8EFFLv6BXeW/Foilo4Zp+8pPvagiQIKguJ
GEs+PM/weF2OxnTq4WTz5IIjdj/A1V+/n9kGVCncHyYZ7S/Ydm5DAkHcVjrh
CQS8YH5m7yAfY0HJvZWIWMNQhe7mNpot/88tNLXgp/AbrTAhJ5RCc7hCn8E9
OHkLdxRQvPqNy4TVJmMXWTbW1T6DH61FaRaoS421LcM7gFhgB6VehbYB7PF1
5f/STldezND0j+cRmJZP16XdxN9LMcbXjUsMWQGPidOSW+gkbxWWKNWbjnx8
Sn6etgDndfZ7rtW3KCLKl/8pXoNUGcRnsCPKldOxvQ5nbj27toE+kDCPdOZF
hGwZUN80KsVoegL4i9t15E9P3mems9tTw5BX2gYpRVzVp8AJ0tQgIM42h2/r
wylDvTfEnzY+ROUWtp1ximG2tF44/bfjELCA5zhDL1Ma7/w70qDKSXR+nAfx
Tmnq1U4VpMr1jYPaHG9AM+C6NdSJZ/AVp2oiSIpn2ln+nxFFLPcBTdiVUc2z
62rlpAYPg//h1YmNVkT7nDA9iMCG3qT4cXzlhtxQnSqMcwup/c8CPpHLXdBb
nnebgoI9FGD21JW6Mqp9WvcPi+Zy1avOfW6nFWbZwXiNDRrHx6GfHU6opVEy
vpAdrtDQZMT8xa/QGs/blBl3sdzn3lGBR7xPjCbq2IgHY0TKugPDO2nN4xaj
hz9C5nx2R6znsvQOyiI800zvNdFE+nyVxK7uqulWpQjSxWgP8KyJeAhbdbdw
FMrXooNRRgGMY1CsjaXYZVyM/oSpQK8ATfAKt72px0338yvzVPSWmcLOo7qK
GgXMkUAI8vhFFtxlTT44NS+7PQed5iEFcEugwoSw3TKHjU4s4ofgonWcTmyf
dX6NDXh5q/DW1FQF77buK9U5EEHBHn/f+Y3JWm92UHD3ET6MXPPHyPaF8EaG
1NQM4Jnn6ktGvPHKtH3lp28kIcdNt3YuMlQEFEBszM+n7KFAfPhQpZnuO55f
/yTremv/etvTbEtwkLQ8KBEMyDf6fMmIIYaUGr3aePmdy8bQ6L6BYm833Qel
QtC91yhEkSxqWQxBP/0WtpRwp+QiHoYuYM/6+9IilMosg1mWm8Tw3d+0Lr10
4/Wg3DMNtWc3RCuEeyvGxOdmhm8GB4IXy28bG8Rvf7RStrVMULz4RsxSDokb
Arw+j82Pgj31jbvWDopCfA/Kxw+oNreCWKF2Xgors8jDp+g4j5mP6nfIUyWP
2uRVDW+S7EulRlTetvdgmr/jX07l4a7L3cPv1e2IctRtlXtx59D5w4yiAU4H
YxsWFVWdMio4r5ZKhhrqWUsehMyvf5jLszE8fvFFRzRaXJG+epBa5tie25n/
CPcacPV67y2Pbz9t/jMZD0JpVLSR83dzKxrEji9E+XwUvKj7o1HkWn753AmC
FrVo6g/P4qBGOhp/pqVbnEXbFjjeRQMCgAxP1CnI+ue0iipW8TnWShRemJCu
IvIbne8NwjPeD/YoeHSqL6AaQRch83b/82NokZTJZseMaj5LkSPI6RD+2kj/
0dO/irn5l2oWD1tXRdd9jjF8o5bEmX1u5Qu812GcCYvI509yQK2EAQ93XCBY
NFFNfQ8yUxoVTnrbrnnsO76SzbF7sk3T5vHa4HG+DAKUXteVqgXAX4IWuP4d
nBB9oZ2+kEN1WJHmrFWgApZEWiKo1Mgg015U3wVtied6Vm7UpPHMMgb1qi10
RwtQKMneJGrB5Yp9tA3mkwzBwp096YzCJcShps503H3faFvUCf7cUHuZXX1v
pd84dt7OcMHAqicFpamwjufDmnSVxR973b+jB89u0f8pog8lGOERBPz0coOd
3VOyugCjaN+2evGDBFGGIvD/plFrpp9LWuy/85Mj773itftOXZEtG82IMGHH
mDmgi5/B849pUyAL3rNorYUTiR9lMQrRmgplxIGlfQIwsirBi8odpesuBJwJ
LKrdtai46pJcLYV3NsshkHpwl3hk275JgyoMJeTpAseYnCQsIVExm3CKIWMu
nEFGLiNp8LpM2o9ypF5dBb0q/Dln9iBEi31OW5gXvm5T6Qvp2YBzZUFoLHfA
Jl3570r4jE/JmXWY/lwmsSHHrdpXALv/KJjlpZBxCwIGtirlAPlCjT0igTXT
nDylUuxI+XqYRELBFgUgPvVHoxK7ivdvWeWinI8hBH18IvVKaY9cEfzpw2Ew
jvBUYZIod89VPyGCfu5+MFU/ICdrxGA2NpgpzF2JWzDTOIaFxfYJIs2NH9Ow
NJpcNb1YQbYBK1hUD8QEgyhdLMZlbT+CosqH+uAckrUh6W364ttXxWl+efPc
ZiP+kmRS/mYk4m8bZtHetF7qNkmjgHOhXW2exQIl3kRPW2isATA/eFIkeXU6
VQOGtWassxb1PZaPjw/UZq3tp7vS831e0K0NhSs1BDhilTKDRzxkcxdiWgXW
yLL7LTDaYBydZo6Wr8vyUJG4YPKZp/n/2a0wZPJgfgb19b7LV1iNR3f6RKDz
JcDL7ebvJTRQseyinsj9xMiecQa8wMR6zC4gdeHKpl9g4EhCBFoMuEfD5+2G
699a0+fQx74cmdNPUBgaF9gx1bggWzIXvm98naq8v4qUN7Im9s50x+yI4cet
jhFItq9xtyivsFkk1vhfLcjmdUYkoyP9uYt6JEqBd4PfgCv4BHIkpi/DHPKO
f+NiDAtUBZDOvSzwQ2LaQ1MfY8ABYxNqML34aoJieli64Rr+GQwuFCIJGpAx
aRXLLgdoTc3IEvPChyPr5CIt/F1kOR5HGU5BHvdIxUDySpPjSmJrgRB4UOzx
sdH4/C8wZcdkXVeaj6wff6279oGoA5lvGz4xwvz1dRwmFvDGeUmuK99IGg37
H2mzvCr/eCPMEZl0b+UaO8m25G7MHktvHnimJD6bPXHF/LKg19LzEXvhkbrI
XA8py3ItqlhpuwxeWWr2wwL8clBcmX8R1K/F9xlwFGo5zNGOJ03rTFt0jUN8
RTfBPX9rI518QvK5afWQ2wVxUE/w5Ny9RuExZxRHcCvrQ551WWCg2tOuTKkv
4U9kTbL/2fAANv+IAm+byumbfMGpKkZ4obkbpcWhKbBf6/Q1O5yQxqenDQYz
LYiEDq5l/JDG5vsMBPcAJKFHGjLFt6xp61ZGWEOpgGuIgI6li/43vG3jjuub
WalONGSuM0wMaLfTGlb3jcNmBFjQSt98+qOYA+Sme55WDjHy/fd6DKdq0kUL
9twlK205PtGOR/QEp0h9zB2KBYuudYMNiQR9nJ7Y0BtsHCPba+dENKD6hb+4
5jLTB9h1pF91K/bqFJROGire3P9AKT36GkmCTlm5OHOuNA4Wiwlbm+fBumZL
dt4oW44WyPwOIMLjklpxRU+R2A5bFI5t3q+czumB6gRXMb5yOCK1A3VUli8C
HiJiyYjrhyp8uE+3iV1vgq08pXR/te51VVRdajmR2Fq0whg02s26hwhxJcq4
SQ8IyASfS9KULDCBcoRFGbo4w9Vh/lUAZOOFzOr3rE9Lae/lE7HIvBlxB4U2
Sv90uE221nFnxCFsMcNoYzNivDpWHewOeN+VwSuAyjY4RraPaxvsMtk4iH9o
WgsJ956Sz67j0gNK/reAb/6ZmiYhJNTpnOYU/Q3pvze/TKkmrN9t1RYfZc1S
61Q7CtXouwk2QuUWqI6MJhPl0EItWFa7RRFS50ODl3zKgWIYDzn8/kgv5zvK
D8q80ga4cFLNx7RXNVyoeJbNzF/IOK0EKMAjixownCJCtlzcNmpjfnHDdRzu
H/C/wzS19y+t6m6QGTaqgQqguJzN7cTHrC1ud4sWeRQIC7bnen/l5dNXiGQ4
fxNwtVOssZBNLqZmxSBjcwUcSSs7L43+zEa4ZkqmoU1C9Uw63hFQB/RUYxxP
6E5QhBfGjU4e7YdJrZmn3qo70S74BDfE0E0auarD2GKfBoch//mYGH1kBNkT
KYBVfht/tQFEJs7bKEUOUZT7d2XlIkyWfffwXVbkhtnQJ3JXexJvFJf11nRn
Pu+CX58vUCIYUqHHlPEEn1ds+TvMwT43gxep3RDflIAXfczmnzV2PL2jkmg8
urnW0IBR6qKFBj1GVWOz/v1JV/3snhfNLGr40a6f9g5kjZaC6Ohk90Pr3pQc
oONGQjebfjV9976vKEuFT7PxgmiwD3r4/i5aXuYz1ISRAdHsLfBULHm0iCKX
CX/cBxkBQjYpN/g1rRloYt1ymiIB57hwo+ezGfIJpkm2NoF0Rsc2kAFwy371
W8AKF87TEXIK70Po0G0VMS4V+8S6vSNBGQ/fqq9lhjjaeZo/RSuyRY3jph5Q
VgvWZqKuj3FjGW/taUNJXkM5dBN8tQDbJjR6U8mhwW/TLGifJy7Xhhru6rwg
MRC80LH99IymVQF1D0u0asBudOBhUECqfVYPLHr7QqXrrDTCeS0B090fM1ri
oZIpIdijvj7DSaKTkRZtvCEwWSPXbojsPOEmf5C4Et91LHZRMx1CIxn7wQe1
g6Z2z+NeI+Hkk/+L5z6IvUyy9bS3+YOw40jwnSOI/pPP3R1rYbyDfYtJ2OxM
XcMm5MxK8iC+T5ja+8ydg5Fq/O8oyD55cw+ONn249uHI65McJ0i7aTqCfSC4
zoxTRDcVKZTpqZm9Hh6UAQ8xflvP9T71WKAr3n8i1rbA6N6diEbE8O8ZXQZw
cdj/yDm4OK2TGfW8NWORKbzsRk1bp/NJuBg64TWKqWJQB93+Q6qBHFV7vJ3+
rkV1GeUt80mREBXIgtlWgLwTC1vItSPSltwSpW1BfXtVeRMULF5Ex6V4iKxY
38EZYocP93teM747BmOGNEh20KASFcsA1Kd9N78g72H9x/T+dP3zB6O8LaDH
EpnnFYqr5cMgP9ea8TburS5LcFiYPv93jxgYCr81uNGavRa5iNmre9ynwGul
bkCvz0tLZKWI+W/ayQA+elNVwKdjbcKZxXYqD9x8QisUSJGuDkyg8EAb6psT
IBTRdDm2Tz/uKLqcY3PL6+jRbnvmgdGoBV2Lj5ObfXHT1nWokrrgfzNL/thN
97p3cBLXstlODAsbp8xA6Pkf1pyTpTGiSgY4tmVQtb1njPk84e9QiDI7dx4h
TjkQS4I2VJ5rUJ4mx1miu9cmU4/Giay4GeDWE9oOOPXSo53AaRUq+L8umLUv
mtauj/NnqNQ8reGwqEWBpR7eDliSZ06WTz137gC27HtI2+T3AK36y5yGg5dD
IZBISRF35D/QjJSh4bEXtXSxEIfsAKziUb3BxiJ3LOaJYbKGTrdhDqxG7I+M
y73r3TXBq6lqrIIhbF0Ot3zT8v0mVpooTu6z1giY3TeU9yfPSIyqTUNmYg9w
KwTkjpZJKT/Tq+Ilh1bCii+jdjgfmoszC4l0tNn+tj4M5RDE4amD1jYjUgMi
yQiT3NsXiG83Z9yf2YrbtIlZteStItu3d/x3q0mqo4mgJZjBe5jsN8c3x3JW
DiHepLQiZE9egkOzUwxpxgf83PoR/bnI2DjBfcLu7fYrSTLqfRhn6/Wojqr/
GFPtOSpc131ry2gyXLrELimMrR+WFPm9Dru+Vvxqbp1YJ1mnPVD6SaEatiQh
/9+50h1ZkfHwDoEte5IrXm2tVGgvOGMvo1FTXK6UL1+hc8RBpQkYOSH/MLr2
KX5iLxNN6xJmWSQ1brIkK4CJk1pWu2ZhUfP38tmomWx8BlAv+CPqXiIUVA2h
ElLH753CH4qJx9IUOz8xO/Y0z0qhVgjM3PGXjp8/7ZsKDQNSB2+UVTBnfLRQ
6OdRncrVmMuVHLjwOjenqQdLuckk1nguP8NAGPxWmprc+EPmc1N6HBgErQFb
gC3UB1bK9302FtQG0GgYo6vi0EAZXLv6srXUKgQH3paLZ5vHjjOlVSg4xM5e
B2pCJlv3J3rFECGHblRUToEnp22zXeTHOVGIWpWDfLIejcaNhabDaG4hyI8A
SJWTVgOk1caggrIPg9RIbxJtNaFo+kzw3e+VIvmNOy4MYQXj62RQrHl/KyAG
wcZtzOs+DwofPyyZ6cii5ugXhbA1psvRJbDM2aUcbCmQQYu79JiyiCbaHYdz
xhVvKj2MFuZHJL5LtmO0ojYnLZh9nVb1rv1TuFrWT4m3EJRHBjEQuakHkng9
LFiRWRoDQijgfhKxvtABoYPi97Pn5jhqMXq4TfeKpytbgLkQXyR5EcGCEoO3
jO5sJ2Qlu23YsZd/KymJgHRIalQ6nLo8BsdwhZjzIer4A/tEuqYjQN+e0Maw
2SZAlnD5toBQBel7Mrx10HLgowJo4DGPNEwU8OqPKDqyKwVD/8F9kZiziXE6
BbCnAWq9XatYVoe/o6J2HP7qucXx05AXc9uXmSQ8x9FkHCmPpDkMLJuZhU8+
ZksyF+1gZNtFb0cKHKJmF/o+BY9aU+9KC9tMrv7G+BvN9ckndFp5U8Uvi7JN
1Py7h+evfEkBAtnvVM29MMuUXUlkYhVzN+y/WtbDer1SK7jwMBxl4E2AXo65
bYzj6Y+CpMbvwH+eaqmGHG6Cd4ZNP52We0lz1TYs6RpfF6GQPH3yowETJlfR
Cv/2LUAkAP2327N2jTZlamsVB9b7e0YCTG2jTlC6dJLKTshcRUQcCi5ABCG4
V7zMtW/VzcK/dDxHIO8pdWPCXzjSwBBqHcKUPltxo5p9a9JCCpFiOy+SHNsX
Z63Kl1M5m5Wr0l9W1TddaG84HuGqr5/dwqNapALmGaQ99dJHV8TaixnJTCgZ
otTPGbau5rZatwc27Khojk4ZZCmf3ncnIM/EhoTw/K5PJRdarIJZA1GQY9xT
JMCreijA1xkEnQmQ9yzMUx1Xmuc7Id0TrS5qU06RyNiA3O6feWZqijs2GiUw
PplxOqtpWl6/Q8E2wgAME68W1FZWyUbcUM571sCEZGvW7RC/w6zL4Z82v605
n/9Ma8Kb896kt97qH+TBbYq2IUUkQG9NATVVv+bIjfUL4JtHCQs2VfY459WH
gDo5xM/PKr79xS2gufWKvShLwl1NUdx0jXf2prHo9t11q/F6ugVCNmj2Cih7
J5s2mu1xOb1oK/lkEHurXSY0fk+t7Bsr85rwjEOxU6EEWUv+c/OC1X61vPf3
HWjyAKQt8mhAvHS1SX8q9OIBrGP0CpmibMswGwFkxEBSGBzLeJHrIk5oZaI0
ZfeLANGtzHuVg0LW0YWXVq0Z57E4JSwy/2ZsTI45YvyNqxXeClR4KcSfO0h5
Zb4J4Lcw38A6rBoYwrfKyV+Ru2ydRBUovek63Lx53X9TqM5g8P/kCppnB3Ky
XRJZFqzRSZgnue5rmIEnbyhGMgOjpuvvSsCQnFXOfUwLs7jIG3eH9NcwjLUM
jFq6xDKY4cq/C9K7ueDizhrYQNmpDxHn6kFYIl6sLYWTFw66Aa1zicvzSHOx
jWOxzLLDI03uKFMfRRoSgO8kf3hUViHROmRfpNUySQlkzB9t/y2x/7lpZ9cw
q5H5PVv99Zrin5Eba1Yu7bylqUzxQljjBkyZsELXxDYFWhWyz384eRu8dyHg
+NIV4lxzlP1rFmjXiBXu0egGb1XYgaoryyUJFGwct5DMA8g745DME+CqU93a
Ds9XbTTVwBHCDBzeouFuIiIS1U2KgF8MdwmGR2BM/a2TP0Ybz8gYM1k4vQSz
cMEau6aPZ5agJR6jr4NNjjoXQfjngcZPm1LCWsc2FEWy6pNtYWSVVzvT3ovc
hcZmbFMOGzRgnBYqwBEnYjZqhbDyPIu1Uz1kKRj+gT8jmvFp9wsNxSWMQylV
o1JS9xMVWNcNNuAFcvdvLqOCqQdxqRQ4Sr0v2VDaT6yY2CAttb669BbM56Ns
lBBnqDZZ0tLH/ai0N8ym6AOziAaTGLvqwuto5Css3gkvRW/NZDYVZHnanrMi
qqpYD9evVivdFmEJBWhwn5Mz8Gp6+p5Snfws/3x8+WFr52R7JkPvWHgyHpfg
rKSLHeH/woqG8ZEU5b/GH71kE/NYXzJjMC1lZPG19dtNJcOyOstQ1YFrCO3Y
WtnGoDXsaiH5oUyyRqJgxoqbQ/JkVvJBxAREz3cckN2C7so1q0MpxFSn/iQV
7AXIlYQqZcPLsRSr0+8uN//B3WhitH6BZfC8PU4hDCzcaysxpHmeRWDQ9u5A
waOTtecCHfoE6ItdsU+J5CJs5ci3+f6bnYYjl/Ac1CiASR+h46kF02iaDQHi
o4ya+kokq0/s19fbfLhCKFK2Vdnlu2ORVXZ0iC8Mz34v4Bvms9Usi22b/H4j
p5vYpBo6zoVEzproOc7w/uNOngY8JkxmewSaJOISq1y7M+vo2NE/A+oNeASU
s2i9EB4r+CngEmBWcbBdc9/U1sb4mjMMeBTMOopF9wFgMVsMa1yS0yIklmKI
PanlFK3kQb5Iup8omYR+iJ8qXWcluZxDrL1fH/UcGDiBxG+qRiOwliCPQ/HX
ug32gYvVY5dRkEdz1PawcWQiW+I6MMatOd7mm47jBQJpHEUHqSKKSBd7+Rd6
FvRDeFJfqyTYbTUYu9xFQQIOKpSXR5DV/RsMN6/kjCZs8tKCTh1p1qxJ5loa
5J5D4WnPlpz2Y5ZXjMCtEQ4mkL1Uwre0Ihd0NrRhTJWOLcGEanNeCzSKNhDX
6nRjZi5YRcQpZelN/vWMuFKUD+Cl6ujXapV+HNZAjzEZBKbr8kOMXNo/Ikct
VBaUEH+QJAmBlHZR2UcvHvblPT8L2xBfTpB9HJO8Sw8fKt3AVm5xEjvVgG5P
Ax/rsp3eK9IQDJlaTtZPRgFBfu1b7bCDZ0dgzotjUDv2x/e+8o6BO+fuPnkl
XGJL0BgCiSGvwYzcnkh7vmviynZDdRgBNANFCSeif/YieIgOOTkMzjSIz2ro
lLdWjaurONKLFrSiy182RRxrc3unGG4QAKFJ8UgLLiHqr6tAuJsE2KJPG1Sj
NCkI05oe3xzGunbgNzf9qWMFU8pEZQMgzELPijXXBlbsRGSjcZj5wR3wDFnm
7osOzlphganCgSFmFk4q5qBz88HskpHmjjFotpbPo77koPlM/GAOKxk1zydU
NwmKKAOlfG+MJX9oK/gdghYP0l4WH5uUi8Ns28afDprpJgo11beOMN/MdFqG
klRb9ScexA2a6uGJXypTYkVKY0KsA+gNoQgv66HccOl7bCoWP2clSdcJcKYE
JlzO/GytigGz66h/z98w6CZmD1iZUQpW/KvGGqnJTVCwbA95VhVJWfS4MrnD
XmMsoPziLOu/7YSzh9sd8Y2NhMiqA1sSjcaWaM939Ks/Pzhl9bk7Q7upxa9y
9Fu+BxWCmKZsfrNwjOUMg76u/QRDiYESyuW+tXhm9zEUuO0qys0M8kPC6HaG
fnmq6j9XiGsNvzHSIGa/KypQgxdfh8vohPuER6h4tfP5llo9nd1L73+uqxTl
v3t3ALwhDbu0XfKi2VrMHfqWxbLI+pjvxTYE+NcTZ8yaObr/H2rTHWplKDpp
As9eEJzhONC/8tz4Rak7GY5dLVFs5wkzbQpP+4XYeKeOmNsY/QlM931q0aHU
xcHrkqDx0/2VFWymbMNgRoC4Lmp8oPEN4cC2BcHxe9Vq7H2CFVnwS45gy5ki
sS5ZD7QSViBvpObACXfWM7zfWOjbYqDUC9a0ATVW1anY7o7pec4nsrZw9Zz6
vEqWgRL6/1pRhHGLg0+gUBA5ZwtvkkfzwaG0ERhNrxdwc1LZRLasDgEwW4ot
6gi3+28+uUZICTU9mkyULiPWJCMwV3dfg+UGZhWL9SIrsBQRHpZWdiiVILtw
6g3OceXoa1wawBTR+l1ftL5jU8NCnr7WA7MgNM3ZHEPCNL0dJ22Fo8G9NvMW
LuDQqMb9lBozsRQQHpaW3+6fdaZEhTL13J5Les0ylXu6AbDL9PMtC4Yz+Ms9
eyMgtNhYjUw744eOs+zTh757jMurIyGZJUO50XsfAS9FHMFQRguA3l+s6Ykb
MNEoEicDuNVf7NmjLAzRlJyE/RvIDxEZew0NJOzyGJlVK1fNb6fi24en3pXZ
lRSc/nk9lgnxqWC/uByWPkQUasdEsAo2Ls2DYevv9DDsXFMPXUjFgpaWpHHi
ZEHkP1bSzmKLX9ZlgTLbbdLJ/sRpVZ9BA6CQZoUrVCcflrJAPLgyRqrjOWst
PSsQinKAbZVJi7Z8zrgY9IKeleA4VHcdW7c0WGBx0iWDPAOptLTPx6b9Dsrq
gF4x2bCH6LhZvz7SaN2Ih/wn7Ryn95vjNpvrb+eyLi5j7ezhRYGv64SAVjhA
IM3YMQrL2JJ1ppjpdXLvqos4vTWlYKwrb4QVCNpEg4Btibl85+7iHlt0b/dB
c4rVsKJEdUdodQoBtDyO9W0PfTofiiAPnLOScDLIMVvWD40hcsQGAjiCP0F0
53jPdJoXvBhaj3od81vDa4D8uwiUywTIMmYI6nw4JtvohfgR1yVrqqCtkz5k
Bv+QGID/Jt3xZlewSk0o30Mf5wUdAdDjKs6I7kooPFMJMpWB1Wc86a2xuYub
4UMcSDjLvRsQDLUwLVE9qny+CXibL5Lqt9fnh9SofVsXtNl0OUDYrwOjaLtP
3MUyCB4vPkyKzAuh2KODgThD4fO7t5nTwJUxZRpdZEhQlRVVjg2WIa12eQc5
T3i0VgRVIXXWYuPHso7d8tUg5eHYf8cQz4xu/RWEmn0m0UWbs1vAq7d2Vyx0
gKjGNmq2FtJb1rI/DMbSiyS6zi14xMexSMUswuvJeKBAP4qMIo3Iq+VHztsJ
t6uAZSBCk2Uiv2jx6CxJcgWbeBVZ4XfsawNNatVEayfGUWo/Th9CXcHCJN9d
MFeqebgZAmpXnRP7hNuCo3xFejio1w3U3hidn8Wi87C1VgZWO5TEqW6EkdYA
Cha1caNEfdvnyfpn5d01Pt/nJjFcVdrjoSl5USO4wa8sHaDVoBaSwTSYSUPh
nfivbGXNhWLOTt4W6A9zFtxJ0womSQDv9dWJ4gYZDp8/BhHOFEOW6PECfUsd
aEIeIaNQo0YQAi6GQVAUUXE99UPsj+HOIBkwSO6q4GmF9O9CTBUFKtEpdAkh
vz9v7KrHQRUXhlFRfk3M1EsdyMHQAZ9P2b1/EN1d702qf5ZG4zrdZsksxJlH
+b/qW2C2kZ6Vck9d4q66qxZR5FIKPcn5mJNsV9phBbValcUssHEvadT/8NLM
aB3Q+6sq7X0AJ1H8BsYu+OjddKivJ19nhLwriqXXHPcX+rlvXP2r5oBpru0p
aY3TO6zD+8b7+wCHa3o0sESwPKNc8iNyzY2zFyBZsT1/Kq2xav9u3WjSVSCG
OOaRUgh6LF2QL0PcN2iyXVEXXcstap9efbVBXy0qQIAhr7yzeV8cG6XnsStE
0fOLXALyvs7rlFC2bzj7LS4gi/uJpGlPmW/L+o45bJaHdfj4YaMGnovfIZCB
LSewrT32CApqaFwZq33QUC9YpgsYITTnR2e0aRdNVnnqSIGWRu2yDNrY1hKJ
zFWc2P7Ju3xssfN/Yb+EzzgvYwSqShWA1gOV+v1gvTsAQLaOaP06AT9bxYNV
ftQS01TFRXctFN1nrn/7+sqHSYO1c9iTw1EuAuVbF8ZXXuISKGfRSJsKxnsq
5vc+rIktly0RAfvfoebk6UrPmFdcIeCPvbNzzRvyOcC/Mw6WFoV/vud/Yc2y
VEnVmtI7IUiwnt/LgdwveJq8VYgFQfpBIN5Vvn/iKKgBHvAuzcXC23dsfSu9
KA1JADikGsZhn7rIaDpKklv3ihhwpYNqvSe5/19XI7tv1A+kh0KpT5/RyTAd
wXPRrSN8N1GSlgalAZ7JF4H9/dmY2IohokbnP+vIagK2WwvniwVU06fCbE1T
GWmnrLc2ruNSXcGLXQd0HevsLgguq5cfF6CD/HyFcbrH2EgkbhzCg1kZRsSe
Ieb4l74/F9DYtQB93lFmx/+GICHedJOu4H/k8rHq5+AZjqysUh9aXIdoV2vY
qcQQ3P66CNtZrmsHAzv3rmz1pZZfZWAmznqUtZOyK8SlREABpkyNtIo+LCWz
vEyYctzYiGcdWfLmKpCVk3rxrq/pZ9j41yUbGNL8n80+cJmN1kZXNkVdCp83
68Q7BiBWSDy5DZUuY5HM3WOQCUHvmtEIQGOMJN1rhJ6AlMotKtO29P4zipH8
WGEfX5+DepsWkfa/2K56GPsKP5ohVKuwZ9w8nzaty/d1IGY6gZ4oVHtpj1q+
eGWRVXQZwL6QZ4JGo9mPoiD+RSTC5m1ysGsmrqGSUPmVQjp6cgTMIUcui0G2
TSYvKovJyEAOIIV8b5D9LTl6Cvs2DArpR7ByjHKtdEafBztaq+dQySugCnDN
5AcMIyY5C5wflI3eJc3zST3nX/wkerYU5Q7mkXxZGdEv7vQ1Ec9/KP/bJU4B
Yp6Xa79J0a+uS5cEMXK+cy+NWaLW1ptpb6Q3IqSXMW27XfTshJZOlWeNMR03
12kdJt1Mxfb59oAN4UgRW0tk2hl2iyp3WomzfgLKOrL2dDkXYFQm2apWaQ2M
RaDw/+XD9XW4s0ffgpsMWTwRFGgPyfrSjvHjohHc+f/WWfIQlu2ablPn8BW+
9fJ4rqdTn+UG/zCErqSrfZPmsbFv0Wdq536qVlPCgGY85o8eTm6sH4edrJTY
O3j+8aFw9w2AjVsmClNnM0QWkhLbssRmLF/T66QRln/I9ICuOe9hZuK5vmWl
luwF99M8llMhsvZac3LDz2zLbTtUbvouz9Uq771yRZvQVZpjeYD6RnEb8Bu5
ncXcJU6EUgoH1zrBJv/ZQSE1CJVvzccrYKkdlTGyshILjzm0x2O/g6YUsEzO
3zT0X3fE0ukIsiapC47btTO/Zi3MnvArMfuAnU4c6S/zIWCOHIpO5mDFi276
DL3rHK0UEf82lc74eykhRXs2cV9J6pq++HmDpWPdjvyHB1RLsbBI3pgOmuRc
ZKTk5LFOw2KB97kvRZfbWUq7i46GqvIOV3SobJ5yPAauzPrxDck4otweOewF
q4C8NxPEDDFtqr7VkZiRg2zs6VWZQIm5O/2mSbd0R5Vc48sucevEV5XcBCzy
KpbTy+Am8U6B5A/fcpAvGamj9bPOpcaOXy6/M3S9wzwgb6JCTBSkmkWuyqmX
yN0leMNvNmm6j1MWVX82IUAzk/iX61Cau9OSm2zqn9qB2WbVHk5QSDIKZJ6p
9pbknz6p2MySgQqzifBcausFYsk8Ag8dsHrTZNLtG5u9+1k9KrfK0g4Z6HxL
NgeFqjZ5y2+vUP4wbr21R3t82YcH0ovBwDXQW8DdVu9C8bjjn9RYNJopHwKw
44TcePocI3uRoxQQSjd5/A2YRs20PFheuYLxFuDLstfZTlj8cV//x8X+DjZf
ck3Fm3zr7HS2LlblykcjYo3td16Q/fW3S2QUj1sIiHEkcKHfMD+n8mfGxBOi
sU6d4DOKMn1UAfwRIT2SMTWrNF41sitdZNWbtzEf7njC/KJd8gKmmJnOVXNn
tQCn9Y8uBV/xv9KgMVQq5Q1ys3WXIFwr0QBIlMeGDYnG+ka+RBJa/3nH7H2L
20rIt6hvzt0F7fAsTbjd44SU4YEN19cyrQW12XfspT2EyAYv7FRtu/GxsQ44
s0TEPcRV3HvA6lOOiByNf+WCvfU3DW4mq+eEPNalxgShUFEyKIMcWEJVDfoU
noy0jIRwSQTsD6X56IAjC7ctCCAIhkA7/zck4+YAa3k2D3Pme7klbqKPS5BY
+hfsIvU0fZ9TD8RLsIt6KYUxZrASZXESB3Od7kg8d6mr/1cvL0mFJOLwVM6A
KPuvtqRdYCz026539ePt/iEmC6kwCpUce1DTvJNZ7dRtMeyhKO7NSVRuv2eP
U24lLzI5eq/PBFgvOXJzhkG4wKmh+0M8PbB4sLNYNw7fRsFr03EoiGYgtj17
sROCeE8S2azCurM+SjzNNl49EEK/3d65h2soQbhQa8xndDchH4yLf2BWi19U
LAjtblluvtlO3OgsBmJ2XIaivOOKo6YOqiP6/FVGPhQ7rBwPQ73Bu35+r9la
jhLI1gi+PT+YcxSKUwpHK9ZNIA07pGK1uWaVRWeptwPaS092vZE/J1BUioJf
7xAwHQ6E3xwLE3VPee4uaSSb8kkx1ff5D69Q/ffAptzl1uL91QHanmxRheva
7E1mzURQoTHSkDTipvJcNx5PxfEE7FdFz1TWI8/Bov278FXO066+v2yMS2ma
0/1+DnAMRdqi/kprl+3DeSLz2b56241eO9pDJaHQ+fY4PqTP1BXIPb8sE6XB
+LqTw3orvma7N896gH3wJHyILmMrJq3JPxbICo3/YNuqHTaWIWGDPRFyFo3C
23W8evPLOgBJgoj2GjxCmed8N7vZ32e+WvnEEw011GsbLThDygMiKJKP9Mo/
DS1yKNfT5bh5CtPOLBenGKWxwO+wC941/mcNqdJ5EfTs01DsHy7eNcHiVR4K
MnQG7ZQgAkofxbenvt5TXbd6tGAo3Op82TzLCfXuyQ3IaGaAvyzi1HKJ1BRk
PEQmaXnLljFFBHvzJ2PMR9maWzxuNieae/qAJ5VY3z4plNpzqk3Sy8qv2W9h
O3U4Hs/0+3+O3/x6jZVCUfwiYWx/VpQXGBWxzsszmRXAyEnn9xR0X1Rdyhhh
Stk8HVy4VFD3+JzUNV4sBV+gtgfrMWEDC8HY2wobwkKegAyqmweLrOCTkUPn
H5CeBz52CV3K/fKs1HQwP+FVtKYPBW+dBFeSeK0IPdWmsucSzdpgGF8dbvXC
4JldpaR7w83CiHFhdVwwgdBYmU3xJei8vrL2SnYspayL+Bq7pG3kz7I/ye8h
MW3Qk4AIGaYmdgdz7p7g04mbcbKq9zx5jaTOmyI3sZUHfn7AhloKOpEWMe9z
XOmEb/f88tYivpAWItWsoxsynLCbDHxQpP7LjDdwEwPHxPM+cBxJx/Xf26fn
iq2izd9qjIRHxwGgcPTS+yAzAgzh3RkUuO3xqGF/NKpBfDnurTcql7s4+0OW
ehg/TAdEXeWrFgG/pYvpp40KLaMvFLjL9JxzQztB1/TPcUdoQwsOJq8K6RlQ
rtTLFjVCSFmIgXZXBk3B964NoZQWaGkN/uKESDui6EYPduXE85QPXXzhXY9u
UAnGVPbalu0tTW0uaYwdc4Ra1SBV7KH8W44hpbnCtqDpkeQIm/aLEtdj+9JM
L5IXENT7+XwdDMSwci7/+38Dkb1Dp3we0i8gkr/cv8a+gUmfv2/t4TQOBxha
Xzu0tN287zNbv1aamxwNuMFYmGdxy58BYxc5OWQnDJHYa5KEv/taRJ7Dx8Z0
wq/b+kw50q+C70Snow6cNZqMcnXiQqW9bFSsRmH7OupEkWd1gy6SEw5E4SEs
Ayn9eL9vILydGfjkRviVbFGTUtUyUG5jtfIgcLrXVy//IRK5UeDrwspSaKGh
DQEtumHYoZFXM1j6pimivgC5UcucOjAz4zgyqnVT41gU+IKgDRZ1eP6TjOrK
YYS4UzAnux5mZ0tHatFdN9kgornPqDpznQBkY20OLqFKxzfW33B/16rpjz+B
pu+NSATwp+KQvKS+QtOz7qDZ2IU11HRJSMJ3ZJf2Zhe3OZTRAOaSmLi8S5Rc
lklJJFTrs2Q9dd1aDfvjbKWxvAhneFe2uLUm+gR45spyd9vo39JOlnpSCQYj
Jo2KAjlGXD6T2BKglIfTHI7i+U3s0rKZK72dYiVliOUdQ750kZoVK/li9Vrz
uEPu21mT9+QS+PcSFUCUlPP02KSncXcPH92GQcToK1KSJJhKpzStC9czs9cy
qNQQP6UmnDU2nZ/G90d7babGLIZ98fiu7zvcQklkHyR3FI+pv09l5alCRwWO
ZhZ3d3wUb45AhDN9+S1gdlItaUt5FvX/tVC5BEot5Vc+p6A5xgvkNUGLy2uE
JMc9ZK57ok2e7TjMpWePTjbWBgagzPLgghG9yso6O5lnypmJz6s4A5kyPpkS
ICJbVuqCe277F6wbezwUxXyvB2uRo7LTrBFiBeYkFAflnSv7xm9jE3w2rswK
2WO4lRnqWmFN78zUcyatzjsAi0Y6aoiHPNKaTMx4G4NTRZfZ2L/5dB5ZUot+
k3n22E2KNUcfuDi4ymMumlSTL7paP5cfHdGoDBsMZF/qvKZeGKrNMMKcccbF
7Rzun5FXudbzd3xmKy1Iv9tV3JB8ygbye/HUGXG3eJn1DNXYRBPaw1K3ZrRE
mXhFUEPwNOcA2ODVFLY4X2tQ7pFVgsVzF+z2MDFrU6O2zqKbi1tdZ1q0VHP/
zaNdmYs+w/uekFzr7uPEDTN27e0x2RLiWMAELJEZd5piq+kozDhD+eQXso9N
CnsYnbHjG1Yu8F1pMlt3q/aiHGxRECyMdtdl7OL96c3ScAJny+Z59qy1Wpn2
/DIM68pHsvBrzHOTs2vDG4ksjUi8BXhkYDV8RkEFEEwBvMvu7SDaGgDq0aGl
e8hsVNi9ey9SBqvrQYYvJXA5S2U1kJ1xaUdTKWtECraNlX5W+B/wSS+pSF9r
2lMgfUpjRIRmCJbqGRZ94xFe6pojm70C2xQRXUppLNfg6Tl2m6pddzNO7fuD
G0tUAJig6HvvMVT9xEa9csM0tPTVpr7t2bNN79V7Zqe7SZW1C7lbyGigfN5m
5GEueuEw5VDil/Rkw+4xEXR2JAwHEPlaAG4mkn/vKp0wQF+q8uGfpC53T3xx
rG6PBdXh1E1HJOkPDEemP9v6vjQWXusDfX7Pd7Ie75L0xqLQrVqBjV6SbIfa
jbBpmyaf5ON33jEZD2I1XB2ARLz8UAaixvA1rKV2SmHguahv8HcpK30S0jRD
m0JVV959jjN/qTnfqDqv7vJLO5Z8RwsF+Di/2xfnAogHNAqvTAv7psxozeKN
wt/1jGzkROBYv0DX5iTD1ruOKMpCSBnGG0hOfBvS69uY6u/D16em8qJesnXH
/ndc7ym48Hi7IrleSclmZWV7GkUNSLpUPdGgzHZ2Su7BYl92ZLcxK5KoNlrN
AEac75LmOBCe7G17juPFB01ufZBbfTu68mwhx+EVTjWGYzgf04ofKC/tCgKJ
DEHI3gfSShbScrVdWERGHuuVtrVH3ymdEou94wVR0t8chGVvBDANry5hBaTC
zT6tHQlYh2l8pg1melr51pt3+mBoOCuM6p3iROyLYyNUfnucToWClF1QWsFa
N+2fWScB/U6u7B/ZoKyr4CRXpascihS3gZ4Tznw+WbEXQVI6K9115epdltsM
qFEWUWhktiWix8EbtwaL8irdsOJLdPLtxDc+iWiz/ZjvJFUUlKIgw0wXtJfN
9b2NYCAFFuEdUYFk9umYXFUWtQff/+NfJiFvqGX0RW0lTLlx9CZjWc/jIZVP
+RgpAwjq07d/csGf37diodcr2lUodN1nN8YZn8GXcC3nwWwxkhw8o+6tR52R
591WlNQZMP2xs0PiH/APtEHLwWSgeW6bN7LdqwnyvqDBdJeF4UcTS1DXdUUa
W4YI7fdxGUvUN4Sqde96uZlvxXHqnXRmrl6UGZJ13pH0XiWTYrIxJXXKQLOQ
aZtgRL6LZXS0A5U35UJllo38iUu8FndD//CoIcunmPpDh8/SXZJXYJ1P1bx3
2p+L5bRpwCK9XnhKnrXbjhsHb7jIoZWaxSLtBmmKjknXnWYcV3cLu/1fuEK9
OsDFlPUDR14joYt855ET9okDRWvT3Zj05EngllAsvKuuOdHroFHpngl+UOxt
cBGjdswW0gArd64rrukommTosDgLCim3wjnD8FD8TJwCP5unZ2IapoXcVbX1
/z9FpxRlI+uCVozNo/ySvawhSfE2mcuVUQ4XZePJngAOvFevJDGcLgiK0owZ
sIJwmt4GLoofUnc1l23uk8xv5Kb8KGD46kTsQsAuFv1vCX9H+qJZhPntljzp
AoiXinRtELgHSnGIM7I+psZ53wsRF6v3hI/t09ZPQF3aRh6Wp5H39F5jm5eq
IFeIVPcQV64ONWc3/XSs+4Np6HqbQgABAdHbK+YJDH1S7T2Z9F8EqqL7hpq3
hm48ZnqPZDCeuqJ7DpAzDp8S+eU98d/KipardCzVlcqVla5XNlsSjJG2FqmU
mGIhFlkoQzaqzHKnsK88jh1jWqlwhUWaQXO4PcMtPaCp07XI/avQDXWhA4RU
J/FKwR2TsajpBz7KHyjSprVgPTJTx306hnaNl/tTdpNBIrLMu+wjLWYxEJxd
ppxjIN7Ol3f25tC/GxVotSdACe+qCPFzNWI7dqs2Lne9s7jVCb69MRST5Hzn
wcZhnQdUjb4oH1/n4UNX3cvHEPXVMoIjY2DUOoquIPr6G515Bu/jsuLGoo7+
hdoNm6b5f0QTfSfP0+OzombHKXmaZcOM3eKSpeNw0Yj1Rw4Tri5fogGieZDF
9GC+wHx78iVwlct5NQN+X5x7TWBN+CfK7yEQGXFbe/+OB/S4XazdIpaTPXlw
62bWLgeacMFMIhkVTDdY3TxBHRU4FLO11qqpwHw1mJMeQLGq0mi6obi5oy3G
c7WTeEmHCLd8FG2M7hsMs1b3tZuTq9MEgKSaszBPf9M1wNFdAqv9lSolBbDG
TgokgaSB6BMKX9xGejAWiATmsrbFQWbwaANksleTFflnGeatIqG5khEoVgGX
fVQenc1I6Eq/4IvDSorj7QNgFleDyCy6gin6Z7z9Sk3J0I7W1K6t8/ZZIcxJ
/i9nORPZhm/Roeyhpk0PZ/SolIXocChgchLpNowUsE4gAoElBTv04ptHEMZz
40bLMKBH+68TbBl8FEoW0Kr3UWannS15UXbopG5vRCS3lz6fKftp2V7gWnyp
hYWcfFPbze1f+dkFh4aC8074FRIuyUyGj/RUXRp515GSHQjh3ILPCO9nVlZw
471KnCzmLSKcmkKc53sQPj9Damg1BzQDuJum2wQ//rifrrSzL27+qtkOUm7G
nOEleuOvF++4xCMVBUbydf0qVfxtqd1HYH2GTnvTaayqP7bUxzUT/5BFXr5p
tTnmJlAOvtZk8E6KnISk3GCZA17G6i+uAqlSjPFQc88zQddFI3rBKlzOgkVA
LwBkKixU1RFLuIKe29t9kHqbUzVGt3cwUOFGdig58Dw5yzHmva+edcwkqXfv
Oc61X7SX/ybzVl8Il5tvAuYo4T3cxFH8UtpneyMBVIE7VTvUSSsQ6DVjuDrh
yoI9ryBCRXfX8Cno0wzglxt5D5oQDa4MO0gloCkZJRqKLoXPjSEPS1qu5hc4
p4PN349NrTUDpFHqWXrkOM7wXFJ8LGMUtvr8fCBJIDLnCI4vwK+OtqUS1XYm
OPzLF2uRyCghUlKxCC7zjtr0H/EtHS1Co8DJCqh2JmTa4KtdWabFURS1Eicv
W4XL7X2FYJZULYOyrYzvB77sijOIgy8UeW/MujOU+RiWeG1JIdE3KR9fke/Z
gJm3AkmnUBeMF+QGsE1ugwOOo5fn0cg2E4aZyICZ6JDIOjT86kK3VRT62Mgg
6ZDIOH2NAOcSmZ1BpFmgOpUgOyp29Nf6zg+/8SPtwAYKHd0+iY9oO+uAfDwT
WsM4yiWXz695VA6Gu01eiFB5Z6uesIZDWTqtOHkXSEvsoxEeIH4Ozm577scf
+8VtSmxWNmMIpKAivjeqz6zdEaxDg6tEGaJGaqfO7bwn4Y3aqAWfFW4a78Pl
9MfzpE7uZq8mh+a17Dfna5LQr8dc+sVWTiL98tDAWvSKeW6Qwd8oJlYpe4if
d2QMepq9eDF4IDSTSKACG48W8dtmxHuJEgItq/WroZX91wkxKJyM6zV14phG
ZKnK7pjYhLuZOMDOLeBk55TcJ4WdJ/mBRH+WXiS8pS6IRY7EsbpCinrJyDaC
tLmcok+1F4f5NYjvpuZ1Qk1egI0vh1lk0H7p15H8B1bYsh2M7JUN3/yge7gJ
GPYUAS8xycfGR66Jt+S7SGpeFaycwNLCk30nZtYr3eDh41OmtsRr8S5UdaYZ
UwyNA3rRHgplb+ic2/rRmW4dgq9Ox4jYPK37MtUYHax7KJP8Tc0LIeA0yPm2
J6wNdDMAQx5MswUIDHV3OXOmRX8nP+Ad7MKfAgB+9XQXy97gLgLwozPV9Sm7
M7WflMadHmr8zepozB9JXWvpODISYpbJq5ZZ7At3yoIv6SL5B+NNW8XlxLAE
L80uH2vpbnkp60JW9hBl4l08OBY4wRaizo3aIwOvkcHZQLh+GS9CL2sChHEH
6JQwn7WM5SmsGZ/uinMlsM9hzUT3sgOV1rShZEEDufifDTqtd3SyE6ydPz8a
VBPg8ps+7E8aqiMq0lJz2p8VvAvBHnAu69VUc7uW+bPt8aRr4j3uSamgOCWm
yPT6Wuf9kR+Ryzzd0ghXgPfHIZXKmyyo7NKqNIf6eT1dUUawcz07z0Afx+vx
xR04vO4IeBHbz/hYFrPxxhuTIl3vi4C8rSkp6Al83wj2dYT2o2PKodwpOOF0
5tKUB/dR4CqMBTs/MdQ2pCe7KIMAKtcs5/YjWALJaw2gt4oW1QX4pt8dhLWI
CncDVVAVpRw4aBGH+0MUUwhzvJJYy1s9cfoe6TM0Qy15UG+gbCFdqyZKMl03
dEva72wE0pvTb8lhfhftGS0AyM0VDA3tiHG9V1Ipu1bh6GNmpho/wwPedluT
Jb9LaSmMhEVNJdndic2Y6Zv45/p8t+gKIHxWNpoN/R7nRHOtWgFKtpCFoklh
vm8B0UQ4J+fw4sf+xR8HeaBSs6h9ZfOB0mUgRQ3x/ldvswG6QxSyvGacxuu8
VFf4QWaL8byPFbDwR73Tr733Etoyr4r8svXvNs1nLT/d/7v5oR2Om05DJKwG
Rxs393PELg1naQyNT6SYFq/XXlGwLQu+KBn2UjmXrAgYmjq+fMuz6NVzHW5N
WFAd/+jrvU+y2PGvtKtDb0YoZ3l4kS+ScSKLpweY1jP+VTF9EsykL6q0Vygi
WgdfXtZdHDh1msPbq/vbutwXL4CQUkDApq425oIKMjMJvdIzsrpiwhWbLoi/
d77VHCMalUoWv5Im25wHfTlTHYel+eKq0rrUKxecndgalQPLjEAj1r34kNrr
RmzYzD8DOt+UYt/2XM6WSQQip7p7nHKcx4D5kq8V1MpRhDDtRUsPePDLMNcM
LbraxlcICn/mosmC1M6JnoDptH/wSQDwwJLbeZVpb5L3QXRrnD0mlPN62vS4
MG6X5yN9XFS33A8Jrwqv5KkKmwVUre67rmIwMnd4IvL2f6cDBXYQkPoVf5Em
4YslnzJu/VT80zUTpcLliL2AnvlFUlHGV0P7UFyYaM3luZ0jOjvb15GjyFos
Vvm0Zq0Q4lEW6XSxsFNkmVfHx6gZSGASGjK5u1AITPQ3brwC3ftH8Rl6RiS/
ZCL9N9gVMk34XXFp37c1kdpW+tnzxPq8oBxFR6ALXNFZC3Q/PkVpwVkFJoC+
eqQduwuimCeA1xRZJyLTRtGqzh4/8adXAGRPfxaM3caPbYNao7ReqhOVpN45
fvaOlFOI0uPd/m+NrsX3YTP/gZgGFTQwosklhVRw/6tTxpoDujkJbaojREgI
fx3fjwmj4pjjwErWAlzVT3BDpggyPxi/h7yKuiqEbfl42Z7NVkV64OyfK7aR
i/NSSAObtITEnjkHOBt7MG5qyWyhyS3pEBtzPHEcKKtdEk6ZXoFiKf+kqOi4
3XMGM5JphzMwAWOBy8RfZhCXx83xr5dyCn/exXmo2K73HwS7Io7OABMu9662
FjYrN6VOc/fybXI7UoawNaA7d4dR/yGk2QgZo//2TLGSRclfXb++jVQsR1Ip
q83aQ4KVpGdClSwL5866YkeooyWGftMf/tm9xCyu7gw4LPg07DwphRj9GVz1
przedD6BkpZ4jpu29nCwn38CJFSEE4oaI60s91NDFd6GELXH9hy2OGjiyXTZ
f8RoJX0RLBA5uan/TlE1u+0Ap3FpMK8OJyDsiyoBYv/P9M/WKj4nI/dmqckI
qQmJ4gQkht08RTuAAC83BuQtnL6aOt2sEIEZD4NhBldAN4C5J9EDhYHw6QmI
TasLGgmDb5yqjobLLUZmbitNixeBD80Tie4g+7YvBdcaT6hZSAIxPV4P7qw8
hI3PFft6oj3Qsz5QuaRn94G+T34YfMC1duXBthc1AJewuU3yJUugmiB5Wf76
KJ5BLP4CeygnfQG3zE/2WNuJZyYqMWTChNimFusNMD3ofVWprNWfxS4ZZXAG
7jDYgDJsYi7H3nTGJU7se56w7EJQ2ckh/qnP4sC+/QlCz75fW2tpI1fXUhfz
uNxDCUUmx/f+5J3xmFMbVyDcxjwnai/ymCf5W6HZlBmoG+PugxN/5u9cIwgM
ZIbeRL480QN7atPIAHJxNAWWGsp1YGziYdtd1D5xBaybQuziRy+8wcTRszc7
Zn2ipqLO4bNWHw8f2IHSXwF0XTxlAK26zIkC7jMM6lnnY58xt+lrRRavldq1
1cjVWNgJRsq5fHudrkRCLyIt0YwJ5xUnsL4f5HhYUz0OZavudntegy823vNX
hpvQLaGM3tC7WbKKDTfohtGoTys9Mfn9PicLjgZXAbn3SieaqPFzhhqgrlhy
E4z2h5XbcCfCVoEwsdPH4ZWypIaKKy55yuxb/0DOoplaCU3LtKNiXeWwx8SR
elN9YRqpiNrnkuxJk2qKIvVoB4zogylzSRAaTrbpXgTz/AQ5uMJsmMfsAe7H
4+OorSrNJwcP++7W6evAJ8yZhDBuE2wOXTLPV6UV8heI8pypjZKTxtJT1nqU
rB2S4qUfdTmHmxCFOcG60xNgRnUYps5nc5y5GHwNcVWbrlmJ95JlTcsZdAEM
vr5aH5t5PmzuVfHzxTsntp6e7wB2KwaKr5idVz4AZH6y1S9VXhiA6cxyFUGH
U8oqtAfR0SSBFVdcgxdAHzJFq9WRO8LcuY1XUNMHaIdKnDAmicgGQEAArFEi
l1Zh0EHZqeEfxkteZPJ0TneeOCK1TQBYmejhtbENH4TO9szhLIvHQ6ncNt32
2OrkbcbLUb0rp4P8OC96MeoYvHFcCpKvk+qqLBkMBUAUtqu98mpvmf593zQk
UIdx7OROVGLBSkI4ewx52BdKwjSye6tDa9eHrOV0XDU2hrDCRGTA+ZoAtnCX
jgRNP0Uiwc/lV+xa2EYZO1eUv8yC8K9E3Cmv8Has58opecDj4ZdRx71FXQAG
oAXRSrZLAo8J5hu9jGLjgLavAgrjDh277uwsbBf5wa4lYemHRH6DCENuUhZ+
hQCLGT+NCbzZtIPezkk+b+BfSppKVjsNYFBc7AZckM9i1ojJNeXtpZyvO09S
X02OzvN5zRwqLywcbnbOsjPRyl9nm+ogTsUNmqX1JNROq3ysv1fHTwmRUNNH
kay2jCeGtgtmvGz5m8iQAiM0IOLKNni1z9wEGSRMLkirpw8WmEytKKaogFWf
RKnwc06gpdiB04+A9mg2zwy5OuGdMpkbwdTYQW0rtsuUfERnFjArPFXuZnS8
/h9Kj7l3DLS4fVm0V75G0HR3B52RkhaHqJEEBS0TAdBjDpbin0gXFWAFDqS2
GP4MemJtKMwYPwDlx2rZvtxn0UuWxZJ8HilsBf7QThDHPnJH7ovUuM6hsWs/
RDbgKSvfQ67OEXcFjWkr9Q6gWxyXnKxm22phR78IHvo7Hu0HJJyjsK1YPJIS
1F3oocnK8+MXcMfi1krUixUkk1be44cNHD5r+GCNwEOr/sAENmdayvPJNLTM
8IJmQP5t8CDYvye3t7RFZcIe2yiwzQamYMenhVq3jLSlAmlHgCXA/ZqvkF62
5VnJQEEQzcvdpxqpnxLufb4EM5T9NfmwFbKaJ+FJ9oDe1THEi51RvrnhSawr
T+FJD9oFpe0d76EHouO5Ol9sfFKw5aOY35wKGT+YrQScZA4RqUwTmLhzfnpk
DFhGWeNT/B1HjDMZM2LGZJEj5uMFa1C3jlCrm0/3Pq+b3WJkPhBsbfzlT+mO
OWNdEVE16LsLiG8mTatTMWAZzEEYyNv0imYssE/v3WBCVkfOt9baiYM1tJsq
cwuw2AycSOXdbm/6iuwWrv7G8yjtX8RuNl4qk/JgH0BbqphCcz9v2s94kNvO
WWIXj4AfSVREKR8KkTpzXfd8Xi6JhgFqzSMggzyMTsVgI14fq8GZTAhQydhR
Rm8BVbf6C4FZazyBPajIR7K/5VGjCD2/qMyVcjVdX5qWogMDSyWuLRkeNLsO
IB0tJKY5q5uxgrV7LDXJl2stGLZ7aixmoHYvyfehwk/Mkr21BLfzIVHXG/t8
3vXFPsk7Hk4Es9qWcMPS6GWpl1NbPoMoxiFjEsWGTtXi0CYtiymviEq0P3px
o0cyyncfYbwF96PEpOMYoi83kRmRt/5fGFkqNwRts3J6HmPkaElvt9PakJL7
3Vn6ufS2oo+itrJF2bHXteBWHAbXueF/0MfmvpSHYopafnxlAeBKXaD2tJXa
36YV6LhJWtrdhu8Gc3BX1115SnA5bKVd0dpZsjTxALpqfliysqoFNjM8VSji
XlgZBhUozNQhooLe81ae8Xtz5ayvQN8NDAbYl/1oaOhZ7JkefuX4NPU1+66A
K5k8fKmr/pwaDf0dLXYkfroyg2nI4sLVJeOWLG2Yfw44fsog6IlbrybAG/+B
uKb8w+fa4hlRMBrEmttYRCyiu5xDW8txVRE4yBIYwzRZYqHEkiw8OKPdoTl8
AxYarGa8TFKFbRKI2gMiMrKoueeiNQ8WCTKtkGAaXdlafF6MYhusQ3hacSNU
7C/Vz963l3nXyCHKpEdH6ahaJxz5M9dKtZGvhXsLYqHsLFAHbQp+ahLgaBow
K831KDIECervNla3vNYp2Bqjb3jIBascqAZEAtB1RtmrEdExEbW5Cu0xcTru
+yyzX9e2HMSN3kxCDbfaMwQu4zOEZeHRvlbudA4uQvSYv6y3GmjHZQgaLvFb
8rzYtT5qAIjI2eI49+BeF/ngWMh5n6FneBeV+yM/QOjNNH4ly37705ybcx7e
cYJgum3+BLlsj7FStDgCKGXHmnPFIsvVgYacDA8+dUSEMW3qjptS1jcN1mlA
c73/3CI3MLf/uPCzVRJTdPTS1Nbi57KA6XADUu0DNMr6txxKId4YlamB7PlI
nMF84e0DJ6tq/WAlSHtn/5C1Yb4kd29EBcBwTeKybwpGB0azqHiCPBI8txVM
Cl4tMUNyWCwJ13D5AQGfhMlDqURQr2wrZ3eYVfpZu1bQzYhXUCrB5IQjt4Xy
OOFF3jCWC4w9mEx+yib1il8fePwmaHFxFiIUFqDWUMPHyRMRS7wIJH7/JmMy
ne2p23o3JPbOtof0/tvFvjdHM8dVZ56mB3dbsHtubNhfzk/qG+UiCNd5j4f4
60n62ByE1wMXNXQk33yPEfIlZGF5HzljnEfsILTSrfsWDFEpbTfTXuLOoU3k
jQJ7c7AIWxd3sXmjDC9OGcZeZs0sDRkkqYwksLL1KXEl3DkZibHkbFAMqiae
XWyURFo8U9neSm4oliqAUb5jlcIb8D0gU85ua/wRA9/jinGek/zoVKxjbPN/
b9CNhPQL5ZqDWqbIB3IispvphNpBsG7MAeWuIF/IAHwBqAmF0Pklt0JNHvhe
lvgclC2/U4R7I7c6tuPDNaiXDfFKchXVj5802DnU2uNIRmfX7DqxkcWucXGv
DAMPL3h2xZdCshELli3ceT638g3yITTrXewZvXMD/fxBhLoEYZ1nWnoMEZ9X
RXn+FRjZTK/MlSz9EP2w6r+yIhivLFdE0mjMZ1sjWIZmEngu3UohRbxel4M6
hfzs2tco2PNabwyVm4KlZuxeRMaoSfMOPJ9rPKdpXBVLLYAqzDynCDjSTNsr
YWZQ0LigyrYE4bJzOd5V4HOldI66skHUIlEkP+m7I0gcnLDUe5SBGtT9lO2j
8JDQ6v27ZJBUybpRfKMDiMKt3NANBzOfSbsqCCrzPEFsoGyVvjzknYep5u7z
+/tXP/8saz+0OIJ/OfBwxq9yGagDS6slN/SPlwxzB510al5wNYIhrDI04Jl+
ArgBVbXittx2/JSzA9+r3ZP6NMj7ttjrw6PxQAXusflS6Moq+zZynphkgfIS
ocFrlF3L859Y/+dOfjwmBbWL4w3vX6aUXbFPxu8NvGuckGzFcXRPjWsoR7z/
+3jTjid1PgX23aZhhUnNrxw15o6/yMRZO3WdAixOHSc6yjh5PU6AeWjQx963
VS63cWLIWvp1AT8mR+tUs7ge3xIRqBtrR2Si35ALnRAQFLp0fIl98dCdFROZ
8/axP18JfrOo9VxUjb7sAFL36Ytjjg/Ga8uLFDoMUtpxLFxrJVhmx9M2hz4t
ipFqWRNshSjpRSXm0+9bLLVU9+yTaRQOKy1rXM+lIzdrlaZQjvLfQmnozcUB
fIO8+C638z2o0idzSKCk0oC4CJaKqdiipdPG4ezC6Ri52gGhNRJYVKpLQneL
aoVBdDJoq3hltJEp7lNEbZWpDAanA0hwY7VxUVge6KQ7DfALNntw1NyWjRjp
P7jvLBnRl+iVDxTYkfqjBU1OUwS+ruGncBs55CYyRCWH0k1hCbqbSjFl2/xs
35KC8OwD4pnMG5LTyiUl7rsKAtXG3Fk69TG/JyvCBQnih2VLNvdA7XwqfSa5
ctMgvk5XfZSTIHOHQSxCAvlWcdMbnYPW8LgQ3Q4uH3VXZe6sMaUfUEI1nUby
P5NuRZAgPbAMKnT6yGgVmmLBjruPZ2EKAvoiO64O/FHpPslzNs3kvy30NLjh
dRn/EfGhp2oFBx3bWi8wsaA2/CrySvwPeAFaiaKTqMgbWHalUunScssjjgJM
CyC4NJBXaJlv6JZ1hj4ruWQwzEilom4NtWwYrTXRpQEVg4m5CqATuzy586no
5G5m2tUdrw/7nWjgEDa1GFZWuqjantKM7rU9T3ElicJ1q/T+eh6T2rYGL+IK
PMBu4W65W4IuUe4LYGPe2Shaa6A4sgKF3eKaEsadtc2isLCETvnDOEAaQ6kd
n7ev9AUdyS8I2GCys/tj5OJxpz91sWAqzhIpPryRL4mZ4VKz/E49PRFB0nOQ
gWgAoUisAreFDvx9xQJoYR0E8rmufyut8OeS8mq0dQCtTa96UPdBzXt9p42Q
yaR/DzK/Q4Svf684CR+zur/eMaM/Zyt8UkeSbn0HXbgrv4swKwoyNBV2yQqK
iZFcHKpanpvussD7As+5MYM39TpDYKZ884b/mlsMiEyk5fyqzOitCvLtPzEB
TuMlq6CTBA4Jiu4hYw+3OTSgdP4f09E/K3MNNAWrzybiMMlp5tkP/lT6O17B
v4AL32qD+QCeA1JTbsjFXDmsWVq0UcIVnc03zQoQk1Gz/iHKd42C0a+RggJq
DNhs0y2umm6AALN4fFffActwy4dKkJnwV3LEuPpwGYfZQXabFT6/nu4tUYY2
095tQeEdhRsWOe76G1+/Zg4IUY164Oj4n4WuLnffV2N9PrfTMupAb9XsmsZq
iVBCM1u5uxOiT8B22O8Fu2ca1KbMb1xvMTu4Fej7+VOnTR97CN/Obl8r5OqV
7b/ZIzMiB7af9S7M+Ta+8HLpa5HNRuSmgXsd0QVkXTHY/toKyJMPjMfwvfu5
A0jL07GyyD71yEZE2EVQTiBr4O0BCD7qvU/uEUHTrMDR+RCFlpgKZ974Iqqw
l6/ceRWeRAKmek+TFZe41FyJCgbbogXx0v7FPZ24Jalra0JqgAQl6I1hQSHo
ZilTO78xervfRs9pVN317m7TaQ5KOci8CMwLaXybDfUZ0b1II8DDoRREEskw
qTiXu03PuDHOz0TnVzJhVrbacRhTHdZTlnh0jSKjeYq1OGEdGznkeCp2cRw3
Xq/jlkhbPe0IgR2+sdj8422PC6lwigS7jwc/TSDOse4ZGbofSYW0otTuwtdG
jaqkRnq6pQUiriO7YLe35M+p3KnwMCspCFp+e7ZKx3CVv2+2i2q77TlHGaF2
pDQitu6Ht6qsedKxcjsfGBaOXSuosOAWwymcjkyFpxIKKErQ1DCakS/j3j2c
rV8fWp4htC6gS/hk+Ssm4Hq2enm/8CCwNiYOQHMKmjQl/QbIX57DNW4qAGRb
Sq41os1Qv33EoN7Bmu5rLCIHJ6T8PcTdENY6UwaDGULu26oHvA0O6sTJCJ4+
go5brEUdJUPbLzR7fBFDLPvO822whmW/XWCLFiUZfJ4erUalKNYXtRcJp6Zf
uuTSI0SifhZSbzDVplHBGs6Ghfr23WD40RtDUBNpij2nV4LN4nhlMObob0Aj
SQgcN+oUOs8Qrcjg9rSfAJne6YpvV2Jfd37aYYgSAARSEudNgqJ3MyNjZkee
yu1Oo6K8sqXtfoXjcJSgDXfR5/pLmQ4VxufPxwCLUr9Deb48oa99Ves+ZFYK
PLyjbS16Pseok9i6yyL9JrxbTkKv9Lr5FJFRwuw28xTD7pa0mFPjW/yQbFZN
wwKhLfcCnlit9ZwhEK7H2fGtTiy/wRBpLidqXhvw3b+vQSAYEtwK2Vz2gNEV
ydaACQwUEVurFsB6VUwbjKXDzvVTfB/g0jHOKnURpi5lGhPmZCqm0WQufiPk
7m+onklHwf9Msl3ar0PsFbXXjxYNdrzhsGnBG/ioGskqsrQgA/kpkj2vLe70
G8k5UPXCugt+Xa5QneDTV69qQlVHrl4xxAz2RJC3h7+yPbkGuOw8BrAL6BCI
1REWb9hY4fR2N4EfGpp8P3xOJ/p7GukaHEdq/jNM+c6VUEwBpKCKVbXkHFZ8
eeKNWeEXpR2ts42pqXRf0eoN73NRjY2H4NupbYf0Qa2NTToKeAWti4mKLTVS
y5zH3tR9lGZgKfmJfTfMhAxZQm0HHv9/OzbuiIEy2RebvLSyaNoGBsB9Gx2t
CZrAvH4zinsC8OYEfFTvJ9WGu6BkuYTlmIHuBrctgcBVVpnfCJpPmsXuSE8C
DtLZSjFvWFsFpvrAHsGUYG6tGp1QI1zMTLMtfbD0jqQ2VcWDqIhkYiVxjH7J
uyEO+iK0qp1AxCQJlJNNsAbPMIwgvzrCsqJR5dlXM+lkIOmARJzpm8Omm9YA
eUzxyLSl5XRiHxKTboad66FOilu10GgjGZ2V1IEe+PFJoyfXEhp0qNcB1CGq
p+Z3XaKMylEj9eAl0zuHSUyDiyUJZCvOCmQhizeoldAxn3Blfk/B+F5q8sVv
k9xi2MJ360jVONm52mHeCEuLPFkpx2KzPe9/QpmPNPmMdyX+3NiSphI/pAZ9
GkzAoZ6utD/yV4Co03sZTjtRnuCMhAd1ZATk0GQpbzJ4w+y42jf47FajXlff
rFqajJhjTR3l32R1XUuHOyn5BcQKTdCi1KP5B7i1pw/e413JI9UMLu/84Ogz
Pj50whtsA3jpz7Xrq7K3hFw+P0uxf4zSKQ2CMaHocPLqztn8aY6+jNfZB3NM
k4G8N7ByOMKx9EsHQ8kb51wgTLbXNW//tj8W89aY5I+BNE0qOZg+oTXX+5/D
DsfwGDYCAVIeFaY6ylmWQd9lkwQZNCZi/iGr/NQVIgTSMRR58MYr+Z6tfVZi
MDvkJT2mBMTfDGDZUFH+qtSo/6KO2Vpd3EAb7LG9vzTRHHn3L3FeNa/uzbDH
7rdm0z1DufyVje4RcBQo3Kq//vVrXBv6EKTreIC8xS9lwgrDMpVkqWO7vJZx
q5QAc4FGCHlh7rWAbE+KaEzwlt7p0xFWN7qWRZvwUKZtn8Fo99ZzaK6lwf0L
zDji/rfGJdVZvj7VwM1W0b8zDCtPiAydQgBkpdXepAPuU+pf8SkYd4jh7yDx
JIYiq5Ie0uhPMewSLfKp9aQTQ1Z3MmrQis3jvedS9leaUMla2JhnzbWN/Z/Y
eCtvu72B7e4FZ0NeU6b0elSBCiqOZ4WsvHivuKLUanmMj97R+QETAQmdby5n
j9aboe3RRGf8hPYPb9Xp3F7JgLjK2MeEBCflf4Dd/1wFYzYL19OGMS9+/hvT
qwImpljQiTIrxcTVP0KgoZ7zO3Ib6ghZqJAmk7IfnDwrId84/4xti5VAHURf
y8pw+UE279zjvtTgKe3K3Qj2BTRNTuChZYAeHxLq1Jvnljrc0kZznNpfskhB
1BD4cIXkIGYIu++gl7Yz7RZUulCyf52L4rAVuJKJuULRo17f+3f4Cn0odTix
Ori269rkCc+IjJtP4zPCKQgZqicZnaC9Da7eNEae1Igt8qtF5NrZoSRYtXHR
7p/cx8qSGwfZHAWUKY9egz7cDzMUvBb2NopgEMo33KtrKvP61tSE4EFK9/XS
pgKB8Y/2J7B2PhP8iBBZka91j13MsD4n+qRnmQ1D+VUqAGODZc0YeWplL9Kt
umr6izZpngh4b92aQHq/qJiTFNuDNy9iqOK20m45bQp8guNOSkXY46GPAz+x
xHdmHqj/hFCTU6R+/HzkNJ2VQ+e8u9DvQh+g6rGLXd55+PRovu22vYQ8OhMN
KYyc66TnlaT2dtej0N/mvSC02qTjG1GruvaUKCD1OnH6Ost2kDvKp968D+x+
mRyyrIFdJLhc+etB6XVLAu3B0ls46OXKvy0nRnWv+N6UPLDsUqjESbKtcvRp
f0t6w/oEK53X1NyhtMCOURAiNeCuAxTqaqcnCEXOwyxUoaBykmbzYGRCNM9O
6qkzXBrXKNBelz8I0FfkOo1oyQtKea5+1uob7tP9j5c5i67U2sNNTtNe1MJr
5fNeihKRhhLtf3Jvz/nOm6B9tPCaTDjMof63mz3lXsn8h5EgSEMj/yvznvlD
vbNkUQN0mtqcf1mB6tBsyTO5AKYHsY/wkMPJdlPKalCCGQ1qhR2Wwnw5IdC0
moXHNL4BmK5Z5EsVSkruklaXEwNZqKQdPwZpSy4Nfitf1RH77/xixu6+bSap
TAgt6ejr8RKnK30H1BhEvBZ0HPWgDfuqMrQ0+CnswAc0A5oFD/7sSrGN+46G
RNQVSAuLmQLDXe/TPeL0dZIGiOt+7J7gQcC1NQIKpsZ3J+YuZw3i9TAjijX9
Dju3nEX5FIllzUzDlhPCLrat+D9VsfmwZr2D0y6y/CWdQME9KQ62Q74Pc7uA
m+DutE5ombdlKckNHw7YkQT7zsV/1J3anaBextsr1yY2G7ovJSTEXYuPB0M+
DzjNv9DwL8FjedppMl8xVCwZi3A4H4nA7rydA0ZXAgybbDSdS4zruCgS9nr5
yUpY0+AgJMBVJOqa2PoGesyD0938rKI9RWT2ZaC/SzvSBPA2Qd8Q6yYlcrNq
Q7uh7Hh4AMf9SLnfN9rd5NDY+FKp7ZQsEqVG84xNT7IwazwSMO8ESfuYEM2A
8yGJFXMqhzHnHCAszAmeA1CxMtSSeB1AdwO6Av3tDR03pTwmxeKIzwxeR/Qw
xLb5ExNHc4aJbk7mJHTCWXpR0kJCf7Oz953XhjmSLoEv7l+6IecI/r3YqddR
U/UviikCEf28PksixQ77awSWEDR/d0TcVCmdZ+cbn8EEy4LWGCmyz+GQ/7k8
M+f/TAIzyiokqkSfgYFYAxkFLOEUqti7M/EIEbUI6paroepaLUlFoaeyogjP
Oq6bgM8rT7er9FtC603LMQeLHAU6nMAHrX2BYKqyFWXXsIkRVplDe1ispXk9
tvPdBJ6xENZRvR1cikUQjjccBIhAjKyCTwKn++RXZYJexLq6GRm3CvJ+M8Dl
QTu68lVgZAURseSve+HYUJK6TjhK17k555fFakMcZ2/RVtB/HtMxSJh6u84v
LdOXVV28iWddATU4AvzIK8jyoGENBakzvc3flaT3CFIdKj+oDaAseNlxRga0
J7/hjXG/W+y4aKUHv+vVIAyGldC5+13208EtC7IOXzmEtx3E015mqQRgH/IF
CYqucihNjLJ+1o8UMRQNRO9kL8MH8e4okPbIe3Ypqi95z0+EBrFtaeboE5SL
V1L0/qhTS65MLf9IQN99jmzoy2c4HL6WYvfh1HpcQ3SO4ifz1DNMsXiZ66Rk
BQzyFdfyZjZJsi0SMTTyln06xF18u99GWd0vTgd/4l6/t6KZun/z5TCgFLD4
E/GkZfEFHKnGBGMFx7HL6LvnS6Byg+mRFGQt3JKtIN63I8vxH8VgTOW6xrPb
HqSTkDjLS3DPBM/OOxDLkzHUtv4ei9wLXyhi39jE4t1hIRsIdtvX5EH0k2JV
2kuuW1qcoqs9TobVnfJ98nBCJEIowcp0OoXziugDtxBGXNuEuyBjdOZVfla/
etRt3WRGBh96GFRMIkvOFlC7f65V2YYW7WkkcdzpoFlmqMMrZf6ncw9r+q/a
5vF5hDEaoDGpluXMj8XhF0Cnm+zH0eqACQ8OVkLkQUwC9H0Z1ez/Bk8RFx5H
ZBgyfY7keAtLQS/mLOEmMzUjqev5neBlR88S0e1/siYXnkR++qvr6tvZb+fU
ESXo8KQeomdQ+aCc+EbB74gqF+WD9dyw91Q3jq4lGdusgZAnXIec9q3eoC5f
7SD0Zf5uM+SawBMZ9dWICfAnGXBXETitek2OToO+00jXK1YRj6YCZGIFsQyu
J5YcQsMhhu8vAwJmqK+AASk1Emwmaz1vpR0rUgahBPvtMDlT24sDR/R8cBMX
dodWkrslswqrcaRBXQVcqRLxzfnkU8XLB36ozJZ74y75fCuPdddn7qh8/PgU
AGgNlZAsDWaJb8KRUeONMyRdcIveoCakXeiKjDe7avx5QlPEN2X5OPGfI5HL
bmxGNyGTlYAgzAeRuEr0RV6qGGRurP9Ama8aHHOumk0Rkrxdpb7nwmG8ydb0
7wzD/aIqqXIsg2HJxkjqSBNQWPSxc/u4qH6L7gm5VgLwho1cs8gYGjLMEO0q
rCzTPY90wIiZgglR+en55Njcii8Wg03eDa0u1IdXCd0E+0SryOOC3/ToMRxI
XLr90Hi8M/cE6nRKceYhPhNqwvASBcE3AT0vqbdAhgtcOjEnpIu637Gh0wvZ
Rmz4G2/7H9Bu4Ku0XFq/OnRkn2q5iq+gLGbLJNGzaIVkcvzsoebUK02s+B7h
6QuSBKn+L60HIPl7ROc2+Sd9r2/BrrNYNp7ikEV142XwqG4keDIdszXneGuI
9H1MFuo9TW/mDrLtBEGVf8htghIMJhCHfbJVernUB7vBV3zkmzYTy2FUZVFc
zeced96mqlcIQkI+SIhJMQTBPz9p9k1eSk9J4bSBU+h1rox6JLQ56HfpMopT
5XTLNg2tCgBxjyfdOL790UPqTZVhTZW2a3GDg1HkqLeQYGtu7EcfhIdXQcZz
EO8u+lrzNCy2khcJbXgARBoWDa5CFK64yTXBDM6lXOu7IKqm9a8XNRopLzYR
WYEtKJdhuhAr/ukOLBknZ5XGFb8cSi1M+i2MTq2qSatKEd5M3TXintKb/EzL
qCXpQFPN0TCugQFzWGF2JU75WSRTooFVZge8UPZJkDoDLsFMZsiNifYyga2E
vRiJxk98XfBnqwPHcocrxjh2WnZef5NFUGZT9dcmu0QDZ71F4s4RGPhvnXVM
BQeVkKLLAMJPKXeoBMRDFUjP0XRZOCovaswfytlQOnuWr2rJ3Ps9DJF7t1IQ
RhPw8FKn3jKWrjpjWMkWm7AhokJAbUl45WhKlCJwH5Ogykdi4Y8/yR8hoIqX
nJf8cLLbav6aHWHMNGvie8kC2SoMQVprxL3/+rY1WjU3vzw+tTpztKaYqnE1
b2Z4Z0+vuyyvjNtkIRgxZPR8RiDL0tQcgl7PPg2QhiN+VljJAdVJZq1VXU1X
9LSqTcOvHMm/B/AQyiF84xpv6H52PNSXwHtgmh019gdEzVJ2aJzupUl6oHea
4c+2E1IlSTBpYBD242CXenbGLWTHo48S+YGpq8fMRcHCSHsZ5fYQNnEUSMub
nwqQdy6DZBd5y2CrcVYIwTs2iXpxhMPSqwIRH0eGteo4k+OCVcYoVHgpPc3j
f6CMDsH3z8LA01URgxoEAcclM4tO0iL6UZHUW+FNouGDYvdCVXakC8ua+gFI
AgiO5W5WrhctHg0Ic9c3kgagAE4hMlv69TB9P3j3BHhLMbobbMFQZGQdu9l8
h/pXXgtDDuXS1Dqe0y4cGLvsaz6wX6PC+7aOYxUH1wYiImNVCY5+WIgBKPGq
C3BLvoqIYUOOafcHQqaXuS4BCaBPCAJeukP0xB7Wqr7q2lJvOXZJXdb++ZlM
+hczoZqnB+wik8LMVN/oweIWFFhkDCPtq0CIVJrnxGHO03PYX4hIHIeLg9Jk
lBsDBznr7R4DIBfnweQNyeab6CdtXvphuzT2s9GlbL1tUc4H0nO0za7bEMXX
1s3hl1YbeCb5jPCc4mR2ci+tGdMYCEbncZziF9KPkbhGpga/uB/NdL2fIAH0
yrG20oMK0evxnXEFCe9Ovy6bU+FwbOEwyrBpBOtpTQhQ/tzwMaVpJdYfICLV
sF6W+EHKDbH6f2DjMG8i8DXEwcM4EnYnrcJnZap8Ou1PniRlT555C0gqBRHG
Q+kTiKBdf23ZBadj24R2lEhnyrwqpeIP5qEW9K7V3JawMJiykIF8mxUK1kFv
4anbFmtM46OUGmjouLd0JbHOvBOKUJsgxfodskPmsIFWNIkSRi2fk6TH1m1Z
1NLb8tKIjXBrPB6wQrV/6JSB/G3lzvFmho7sw8YVQe03itSnxzBseskbmHcE
bSAEDNNPd2lT6ArZqz7J/4vcfgoWMEPXe2e0x9V5BIIWKprHVatW4HLj79Oq
fcz/R5/SjN2fxxwbRJCKpeeyzgxsTmqOCOSqexhVxlfx2y7B5DVHJNCNzDrx
PE9cd68sB9tphrDa8jyXeOEkkI8p2zeW6Evp/c8Vv7WBv3emN2ztW+bcGPGJ
w3zofBdckByCcMyY3/UE4zOH3gxukqsLh6cbvVCD5aZAKn8zeD9YK+9Ri+cL
4/OJBPbW8BFR3LYfbtdr/b0hDII4QvRvY43roy0131HKR6oREfDqT0o9aBm5
qGOgPhoD/hw3kOzEHk2cICDNcKZrfxVPObcln56Ms0cje3tE0QjZES/HeyJz
P7YoocMiP/lA1IPvatL7Btwk/nL+CsfuHtA0W2qaeNSTJTWlXFGUurAy1wNy
kvQ6+fBHPtdlGyqrhTNLgxGVv72tpddVhKPpyn4INzKdi1Meesivrz66NvSk
UerXtQOgiUlZqdb/kOAuZcGIGSB67JYcTdoaPSJLOqOpX2/kKGTwZEef6tT1
nCs+vCOJfUB2lw0ZxKp2oAAKQPXON81u0z37iTh6LIsLDqA7wh1gW38bB14h
CK9WGDXeW8WXFugb8dOHGrAdDZ8JFIxBo3tVbK/DmJB8osFN94druGl5UXiV
171qTWUSaIHLUjc75pAM08D3eklSt6GhmnxYe0bKXJPh2VDH2G2BaB8Kqldx
3fhposbRgfj5M9+GrLfXQ8mqp1ShB0olWpYLvrBd333DUy1L/VRzJzFhUcGA
FcsEr82Qs4t6OlbBk78+KxDNrwn61fPGw8/C0LBd3Urvd4nwXJTtd6G+oEKq
dyaOPFNIYzrZGdl00fmvdDdFx2waYEG3UOrTujKR0hXC3KlV0wQbR0HOdlPg
YnsD6LcvwCy/JraVDQhCT7Lh1hr70B1Uic47RFg/ysDwD5nijIRBSmtmSvcn
ws0UMOnzPCz+pQs58L0WXqDPx4z+vEYkLHcO+D4lMxrwJpFlgr/WxIaDPaSn
fzOjBVlMjtpjIUBUPkqkhZRsSkGBBBUM5SJ6Trbst66EIZCP1iyONyyJycR8
0h3deXEsjcHSJ88ZjJm36uF0+dbNwFCuiFTBp7SxjGBmfCHF0oAxQ5Vs69B8
JmApPWS2sn9QeMoAV5wpqndVmsPTYEHjp80LmQgNkcIN0/dPlaKsRdNPtN/a
BxG8PFJuk4jNPngzXHQ0+n+ePSsZ1NRER1Nd/ZccI2XXjOOk+ZzXdq2Xmh3n
EAXlzGFYncgFz9IIiPXAQUoP5iTAAJINJOFAMTKqejtiWTK1811IatRXZfN5
N3IbPrXO0c1l8AgnPwPe2PUGUhIfNHlwQrpBAL+5wJVCUALH9SHJ3V4Eoyv7
j7eCCCY8/A/UCuxWWeAgiK9c3oRM4qG87Wqla0/uprblKczAXEdxLoVtV2ZR
x4wPQmaOTbdtKA6Ctvtxgw/rWX9Ei5DrOJV9HJZqgB3nPZz6/135J+vuHohu
CwBISgKBi7rn2g0IVK0c2VspxU3t1lku1RLAktyYFscsS2uCn9EHsyzGpSdL
WWxmZCwNgq4SmoCTsPqAtW785wvoE4nsMq4th3HVsEeVhXUBYIT3qOK8Y7bB
fgiR8Ws63y0f9T3T9qUJIxIhu0X7kenZ4DNVpz33bjvzKBzSq4vprh7miNeM
bEAzfIzVc4j8u/6w9ekYpkNpPp7b2uGghuytwwhS5Q7xNN8kFiwUziCRzl5N
T78PMUn5RaP2vrD3caR5jI8gv5vNNyKUj5XTSPq10jsn6daq7it83jxd5ibc
1ybv6R7XHVRPodKFfuNleeIcjxpe1oOtLdbO7yNdiVddXFDNwkY1mExZPdzi
gZLo8CoRmsM/nhArojUbPKphqciWF6x/aCI74DOCvhfGC7SsXsym1+Pq6dZf
k0dDGTMNp2Gv4oHwfNAaR3JHZY4wOM6g07bGwrb3UOkZSFcVAoRBLEYKMQ6M
dOZFBiFGCElZjGqEgYUiu+DfzezjFffe9eOUiEiSl1DpJxqJzugWcho0rMnC
ngt1JXP/R36pT2HAcHfSjo7EeSvcC3cW7wPo+iwBVhHYiVarZ6jQpC6fo4FH
40ihPBAR0b+Y6PxMrOYX/yx+ChCVGbtKkY6Bcbwyd7b/Vq1pdK71HMvhIVbY
qQ/LprsWnp+gjQLUUX/NB88Wz+h2jb1YHFrnBwABj1HdeBs1++PXmD3ptwcL
20Uk+RvVvrsbpwR5m+XTqxiVJ6ipIdaaDqr1uqke3MRmMD8Pzhp6u663/FOH
T7WFa8yVpl957UuiesLGHr/1ERemampskUplM8aB5IOXc8JOTtxF7RuLocOd
20LF7tTATf6n5EUvRRP1fnL+vQVfxACHHcCzsKqdz+brDbhhUL0ingTD2m87
PdW0a3BLsZGUQFb8po/mkFa9+dy2y4pfSAi8Acko6glqp+fctGwt50jkJOuf
fOxJnRSPKwRY3xCtZ7lItRrsWWPjGMlOr9yGsD6nxPKfOYNA1Rei/KJIqjyg
+rUCnWz7BmO6kTUFmAP3WpAd2WIhR9/l7/meqz3e7JhE0saIAhQoxMt/3ZWU
6GqwD8F6sBUqh+FI/ZIpZ0foFlx+1XOgT682uRogWw85imjhZ9d4Ui77Ndil
jBKiIhmOYgMI1pJgmEhZkVGd5euQT7e1tkUYL3M3e2JviXQLLvO9RCDd3Hce
b5TOqUCS01au87oqoIlHXhIXxI2893x/js6Iumg0VFM+u4mlt3UCZDrdUvVD
5lCbxZDkfqfJysBZJrbELQFNlCtTgHQ23y9C3AZPiYEDIWF2DPRC/Dkk3W7S
GbqjBX0qkWqiwiIyVZ7n0dD9Sn4XgAwQbHP2b+03H6zr7ty+0RhbB5iDVUuC
DWpvmRYfGs0cIWFGyfPfm/yPBtw6bFSQNFt2gcukGUkK2RNXx0Tlc3cWA9G2
HZD+Vbsae8IUERZ3Saa/XhOBV6y1IQOmirFCqEOoyTTbqLaaUnzq/GVzhjYv
w0eOg6cd6GmO4dfTDKaB3PcWuPAZfQNIclcGjQKgttff3zQsoobe3Qa3vXvY
ZXqyjkTOOap2sQdtgylRvEwxbIX+6jfK7D5t2leJKAwVc2g02Y2KrUx60ahW
jDJGAAIJOGbASzAtLwkimglj8jFLjTlXYBOILLELYDE/34GDCFKyH79/YczR
lNmgCaXkzmQMZKWdddfPYKrfesYsyZ2jGy+p7iOJUt28+NjVJitQfPB7zGb4
948CaW+7lHL8eteDA9jqPLQAOJQGZW3KdFf+XRHhbs8gBynSFcnuCDOZVTv2
XCCeDIRZ+6vTe+ZorFJCVUBsfAsr7jeRlIrcIed8fBqY7eVF9g5DSKHjXX8P
H4WxHLRrxQNnKFNcBh1uxhFw7ww0O0F2SQjLCzV5OF9bE8Il39cUdWoU3MVF
ISw2PKzxwqya7hefMnhwcmFda0zIlN19EmZ+nKZB5VgtOWARYDOeiXQ8if9+
065zS9pcBukMVHM9hAAvB6DYL969xiIhbS7aSqO4SL5yW/9WEjZ38EEGV7oF
a63TABWheIMvJbnzcT1gl32GmBX25AhLERNtR/CfPWMe/k8dCjyrr36iqLf8
3SGOF091DMIC+5BZ5Wq01znspdbavyx8mpKi6l63Z6NuUUIW/noKrc6mIOvv
oCZItv2a2C70vQwNtk5qAecHBR86eaVDa2M288qwdbp+uc2TUT33+gXbCiIz
r7sgFJaF5xWerY30oiqkO/G+HhQGtGb17Xyb7Tmwfuni24Ga0r9k5j/BqdFP
SzPVCcgOForbkPYGAt8RJaPgHZ5njEX8gyd2X2hINdOpmuDSn2l16vAuobuG
xYZ5ZF6I8AAlSw8+wxsmqvJlO2H+lzFDL5JitpLKdwnVIwr33wVW+juHBTSr
qc9fDfI6RzeREseHTblk6vuMOLxlNUGhNXCIHWZj1gZcBbvLi1fT5sbVl3Tf
x6XQJpBFCcv6kmKwqHcpfxc/jo5Ttdvy3zKrRnNcVia0HIi2bZpFvTI+7j9/
ZVTHHLF2B8Ph/xbukg9xwfvyKltT0y2udEcmAxNWZaPvPYaJSGQi3qoXSoFc
jrBwTG9AxrNM3Lt1+g+YZQ/F2a7h/zEc47rboJnjK6Adul54vLseFXybfJz2
CBX8sA32cPRMaZ4TVnRp5Dx0RtnFPXlohkuT+GfoCzhiWaL7wIuTxFQgheQl
y7EllFCGbXbYvPsOb11RTrLjRqygQIYnhvSJosHaOiUlJRC2cA88NBp6SQVO
a/PRMah5tC+8V/0jgA8JvpT0WLmcJ14fLO5RGjyT+Ad5eQSF256NbrryOT9o
8VfRXCtaueSvXliXsuX4uRoTdOpAip55F0FAJT9bvWl8+OEhoZ2IW2a4glCT
28QQ0U/hi/kfuSoEKF+BCVpEgNt3nau67WLuQ5M2LR5OxCuhZj0c+Si2YIqr
eC9hwqZkhdtsZ0Se/GfQu5KC/C6khEUQD/VUgqOczRp9ZwgtL1mP7mvfDfI1
+gTfylR2fHvv2Qb4NwEqMMB0YBjZIbDfkMgXt7H+IvBsLP6GkyTw0YCan8JS
ZF/Qzn47YT2Tjqu68LaKcPcqyXNQ3bb3WkDyVuQN7sWWNXVeCO5EBl5WYBbs
tV5RSDEzpncMXbV0f5XyGYWbBvM692AU5NpCthU4EuUYy0dGaM5VrKb6pY+h
WwZ9xfOgKCYJm5DK3MUnNfWPlyNeoxuWBUVYO6qqKNgVyi8t2L3nej1uwnBz
JQfzeW6cKlKuXx++pDtc7ydZ1tzpqJ9C8i9Vtpk8bLjFjPhj+LeaG9oS22KL
1bxPS7d3kgyu9hOEPlRuH7uJrO5zx/j+S93gVyZ1n4Fv06zZrMvEMj6MnH5e
W8kwVIBIT2E8seJisXIkTgddPydHerIGmfDRs6aUOxms4CFuyhvnIkMpBegV
h1cU95vycF1xvOwNFqqSXCZHcMfwMAIPFI37YHv+eBV46h1Bgv26TvWaUXLA
CNhSHw00hBw5myp+xa9W8OTb+SKw2Gxk9Mhxgz8Dt2DaRn95uDVI0ScGCtjr
6ExIBN3PbE2on5fHoGimq5eaXbS6iY7VNQ/2gswfbIcv8llQ/R0DXTUhJdXp
AH02OROBAXhpXYFwT0rQ7zdAFn3VvukqIMquWfn5c0r5bKMWosHjT8nbWjZ2
66cGpRCSTy1pB7/pN2w9c8rGVVQEO1Y256ZVZD+R3xJw2lTPl0SCRPYWFrZH
baunSdzuZD6DCztDIlkw2Wu2hWfn+YRNpLkuzllXwcEW9YpgG1YY7iApL6ul
IKadhfiMsE4KseB8bMC5H5q+iXG2R+7Xh5s/2C9PMr0DU8TaKUDW+yRcq+dL
rQhp+7JVAMiiKGg7ebH6U3kJJ1o3FTsFedWFykiZ12TkgPYiQHhVWRQb9D8z
e9GO5Wwg3R1GQ+LSoxU8DLxkoc25FltFaEttU6ULI2r5FmscVV/B4HOAkpGb
6/c1eAhK/dhNyIRCLmXuVf0mU/D5K9TMncsrv236cOsbmV+4LdHaJLnTN+MB
GtLUqphm+fT2xXAQCMkXjGjKWCTQdjLToBW7CrnQf948ug8FkV9VCiJ2ZeQx
6eWtFq2fH2kLvAVpzKGtcmo8dnk+bBiyYeS6R2HkXYiBJoDyl+IDOBS0trgd
goUFlr4PI/eXM9O27SB0nmSl/DefyiZlRku1LIXm9kFAP/J+7B/4Md6lj+ku
qL6xchr72syMtR6G+k1toYF8qU11mLmuhKSiNsSnXbqH3B80E0Oe6FcVVuEm
kyax/zINkj/bQILb/rM88KLuhS7HvtTfq9IKbAvI2AITH7nMxkByxyh1bcSs
o2Re7O/T9gK0xiY8qGGfdpy3hJjAKbJm+ymT7m/pI+BOd7xJVilxsQ8QFSHH
3Jc2/6qtsRcnVJvsg1yx7OCy40YUaRz8LMreYQpg/n7qwT42qpemyxWwLaIF
9dQRNzyAR4OqUCDx9YRUx1d85VWlT0wQNPv5z1AXKOwMjgFZVsGBkn0oYiDv
it2gnsMbDvF1vTTySpMzXRZzBfJ4nqv8yb4vVJD5t9MNpprxUMf5TwA6x8/k
rS6/DN0iIxpRhhvKNok0XNqmXwZR6Wk5hP9runMfSxSLcqxWSQUS023bMf0U
T8HM6m8252h0fxliN/c+E328Q9LphmRIY2RTK19pdbOXjdXemSlTatuVYH4f
cW5kGy5ByzHauf6EeDlbvYOO8y9yXVTSwY7wor1T9Bo8zLY/oAMgqoGHf+R+
Fw4OyV3VgIWjgv2Y70JEW4pdsmdeWUAWneY6XL1x42+N+Momy/AG54rZ5wYP
ND7VvK8B9hBQ7GnrMTG5JrNjaYKinlWLegcBebL13iX2AppjZfhdTPmvgEkR
4ZHZTcU2XzF1GiFLbMRv0IEGqnTqMwjOULLWFwHY8d78YnfsZe9m+prGOIJP
lPecj4io5kB3j4O0gqYhGVuFBeyOHd2cTGd7/pFDd9SDj7VMcZnUaLsbP3Nd
PvinZVBJC1tYvZUHPwQxF2Yx/I1uyN4PRml6Jck9IxfoFe2mNlUgtI7aW/Ky
C3ba/V34YOfBXpq+t94ozYajEie5fO72EZPuy5gOp9pYrY9XU1Kc6Z2qcHY9
2Xjc3u0krH0KXJPwV/le56u3gPPScBDQ/QlzhXIkMqcwV/JGe7OObGDjb8ea
7fBfJedDCj+q56HL1c9V00Jc+EO+V7hEMWWVl+6NzPALZ/uFRKhaTko0RJLN
zMBwvtpuycjpDjT1vkgli3RVtDV1Rl0nXVN/CUUiHhBUw/JPyh/CsOctY0LS
39fp7xd2KiCs9zpfEDV/jPjBylUwYGm3t37PPnLXxd8kPewg78A0la7u0v6M
jKJY28XSot2npN7jtydlmG0GyNvPILQbRybde32oVD9wp5VTEJlNt+NFmcIr
MXnb/833n/PmKnr3OeI2AzECKp83YwIrT8LGWq3OF1HBX7YC7f4O5Y5A8sSv
WmtWtoeNBRxHCw8eglWol2II8RDli6Nqprr+zSPqXFyuct6YXuUbSTw/l2gt
o6Tvx6hZCTvEIGlmdxktE/R/JcFmtphH2zzVqU5CssXkzy0Wq6kmjVuMDY8W
JrXDH6tSFMGAeqnZx+04OPRrgSHzpQbrj/3u5L0PSMqT8mNZAaC2Gs1Fe5fe
/ciRBgf8x5VyS+q9NbX311uEpl631I0b4dSP3fI5APz39K3I0FEvviZzYvlr
EmHxK+eBZq25dOhfoA8sUNhSMFfIuKXF9AtlJ+DgboDsm5tQTtEOGLks88VQ
3eAfXYSMd83LOM2zK/A0mIP9p1HQxdrLbrhEYke6WCQroAfnUj17oHqIlTKa
6Poww18KkOCjCSWpv7y9fH7vxuqZ1U4+mI0l0zTEYHWF175gtMCiILM2Qegq
Rsah/lKGNIIYIc1sNeMsr+JOpfFEBgTvV0syFq7HADFHwGLFra7pp9u8dB2k
S64gqN3Nz8B6rb3HkdrmdKGtwAG0k+zAPtZTImw+s1HSW3/uMO4HoPm6Nymp
Npd40gDqde5qhJHUPlv0mh081cCq7QbfWY1inGVcyMXiKjxqMthw72eF3HMv
QXyPjeuTR8jWEITh35swLIqEXqQwHf3GSlIPVSW8fnn8MQnwSxlLHmJ9TFMD
IVAP9UMWr2qZnuY6kjNzvZu0XjDINDfCMbRWpAPzjwPymS3DVpNxC5SBqRrc
frNiR6N1TbhjDdJoviug+8J/YJB9MiMmejRQBtxbuKbmI97uI62GT6RnfIef
mm5+5aQsBXl11Ecg0Gcj+VZbTT7MYtCn0PsM6/KR6QSDf6OrnVv5SADiYrcJ
tSV8gW8WupPlidDxYnYCmZdhL+6yDXf6pVOsG8LQvcvQP14t6aKXlHPLbBDI
6kDclFhRKjCxfWjTN7s23mrFVVlXng2jQ3OU+akMqEwyESv1RE/F4RDK2d4e
DyZp++eSflLE+Hr8QynfTS6V0JC4zmAyNqKG+TYdFYzJ7zVTN6pj/RH5vXj2
qi5qwW27PPtJdSEzO7e8vOsEZv4ssmHruyBOSeVJEQ9qEZVYcHVoAxruEJjb
R4fPnhhTnI+evRIjcRCMjEcUqkq9kmbfrtuVNQqCvHt9qWQY2VwwFpRf5/4j
OpJZEKCw3sVKmHtk7hg4E1J5qa2iKWqbvZeuTYjTj6yUAWtfa0xHJWHhp4NK
eA5+SB9cDdZPZ0kPSadmD129yqkru71t3JK191S+TEqyFzoDcCI78Sb5Sv10
SiSpQV//YlxhNvm1tXQFdm6mNNcm7JX9hhqgwa/qLiyanuiCI16yXZGM9/eE
leC1iUJqy67wAlF/RzQ/w52hu9w2wixscSipgBLMREFWbhjRQX88kaRObU4u
BQXcvQNEKG+NkcggRhpVasLPl0xosSrK3pZczrDD93AJozHZpTMqXgLOkIzK
cZpcE8NeIiUcg72z60ddn22LcpdaDfgFGfGsXJubzcdqPDU7T/eK2NYJN3gn
bPm/OjT1Fr8xezdhNUEKmk5ucJz/nCHmQrw3ygyiAvoZlag6LUueu64dxMH/
dnHGGCfc9hfAXsFIRZlKs5XQ+hCevVBWAfzY8h1K3r4wWsnolRVjyDhfXZAu
I11BwhcngB6MFUidA7uV+2nrOtWWlt8KBmgcaYEgRBVI5hwh5IAMtX+Ych6f
gcAOujnwJLG2cScJLTihw159JdbeGyiQlk1k7vFR4ld8SkEnopSVvopTMnMf
Cf6rKCm1j9GF57ZlGXIFVVq+OQeCHpvjmgUwWVLw+CXZsn3VImpJPGTlLwAM
jdZ+pUT+ft2dTvJ1aakZFBppZF6pGtoLNtsgxqTzJr+/fBOoLJR4nB+F0JV2
KpKsPPzKt55cBHaQ8ovCt+wUlw5m6kX1CcGadCCZAySAlCU5c2ET8O2y+8l2
yxSNhYSMt9mMNubjumeTD4jJlboGyLvZAAoQDPovSvWDHPGaXmn0hLGbmeBz
3bEeBATKZER84h2ZUZmydhVQiUXHxs4SYUoCsHqd42SXf4/VDkR/adOo5dMS
Vq5DFiU+8tKgTisfGBbqRLMpBcBVIjK8DIMwVWYzaj4ZuXpfd5UlNExl4r/F
xIe1qHTWu74ytbn93VyroZim268PnGexoRchvuoOCzXwpO1Jkce6ujt+yISR
8RVPPwZC87nM40pGxqzFO3F3nTG7/RqPbgXhwL3oYYmVeuaKBOGFFynfsl04
uAZDkm4Hdlc0Qb/C09ngPCrQIg6M6gCI8YAnWf36B3gmBFYLp2omipIVe1XB
aedHb3xa6Bbv1IfzgmtN2RhIIdQsMNzcE+vI023V4densFrCW0yBD4zWBkLC
Lu+1xycuYYquH6Q9Rj+aoEMfCA/cqBWobIInm/Du/lhDEgoOD/xbVa/vuhVW
gV6nlVjgB5HSpTtaHVsJp2Jp2nBGh4kZ5+Tksj7qHmNALf8AIuhN82iUfh6q
wt84sjpaJrd7rv63vfz7gTU8dYJE4Nd09StDjfFEPqlC3hJokDCfZVttpWAW
qJ22b9YMheZlLqoM0vurPDQnj6zBKH5NzQFKd7HjpN/Ocqqc7zDl+9rymotw
NoceDeWegufdJ//Yui+e4nuxdslAKA5bwQrf2CehKxw2E7pJEiFy9M9L+cWL
2UpmdXZr9IWQOYNbfIyvIYpcHkGK1ua/CPPFsrhRl4C2x52il4J43YSZw0Sj
YlGWxAWLX/i4SiQRRCgDkjYsFCR4m26ke41GTNKZxyBlse6dDlpZonoVRRNc
RQL7zucQ8yg+D4TiFiqD0OM9xKcUDObug2/NQjjQyS+jON8k/RyCfu+iGACI
7bk4t3Gf5p1tqmBir5zrtJ9QBw8Dl6Wx3fWOJTCu9+GHMNEYrGNOlfPL97z/
H7amkBHrgxf9gceBdA0XSm5fCz6ANkzEcrwFWgSE52YSR7bcdqns75dj24eO
PPIqRoD5C9j8nRQuLzIErWIiej8/NAQL8d+TovaLFmvXRtMoOSXTDq8ZthRO
nbNe0j2/dxuQy+qoBURsRfK0o7IbQyYO7F+dNDPSuncwdDoQMjAR/GpyD/BK
lzPBTRLtBThqxe6H1mJNWjxVkYo7x+j/Gzc/mR9fzGiQL+P9Cyh74qX72tXT
qwnk15+uo5gIcrO+/gNOw9F/kX2mQzBv7vhKC+1ve9vVhU+hwE6Y8tOnRbkQ
cAFviQeHjLBnF8QcydFfjI1WYqlfO3Q1qIQETaoNQmllIfRQLL/vZzSFs2ay
oS+zzishmT1q8nCbdhzE8Wle1Mro11RFdEbBPHUS2dQAWxyvu4Ku/W7BFzKn
XYRo3THRkEDfluLkAOwjwjWRx9ARll8WQNIyQDdtHnhZL4x2tuOZBgm9Fq5N
wB7PIBa8KR3zgAPS/cKhBaeVnLEcbWlM6ZmMd/ZwcUUqQ0zx+REKkeQ3Iva3
bm9j8C4z7TbW0QVQx62uSZEDuRtf4LJUsp3/5YNTHH8s6ys5C+/1/ytyn5Co
Mo03Zrz8g5aDeWSZvZi65zb7wI7cThIlu11LZUg672mjBk04DAx1cWalpSn2
56UmrMNJKo01HpDzSis9VR7xWq6n8jzsAKKILbFWB7lieGLx64RxYObv98KS
mQy8MfwGzTyQ9JlaRjOtkl+nwF1VH7i16uI7VT7RK7A24HkcpYkx5LWtsVoP
w51HGwWoYczxNSAVGWDBTDAj5fM7MEYfpyHy8hQd3rX/v56jkvs+WSjckl2X
Ne8SomookaGCL/ikM8g5Eq+Fo8e8Qba4zCRrpqHMMRVzg1ZFFfV7lhozZGEa
3v2pSrkMgFSEUTaw7TNf8PgWdqkYWbQ6wFZiC4CuIWPw1BA8AFblSgUPO6Ij
249JvpEjc1F3BDDvpY+EVbqAKBiFDOXxpU2Y5lxCZs1gIKJWy/0j6JXUtcMM
RjxijxLBGqkEGwiF9llIK45aP87+ieqeSbF8DNtlZwYgjaBjLIKDHgkIqX+X
6rBvdD4KrTbskai/THRf+YYDdNuWLIcgUJAg8APsEuFxwFDwdN9LLxt61OOH
x+X7tlOnGb/e4y0TBI7X/NVEtj8QShjP0f+lKuFNtC5s5aYdJk0vKSIw810L
4LAQH1Flq1wC5BIjlSGJJL+Mhrg5hPdjxtLUxXE9KO0da7UrpL8x3fJr/XUc
EI4/wkc5V2uCdZvtwmMOoWzO6LpT2HyIlDBNEishGYWj0lASxN8n9mJT6ZdY
LbM9Hx8SQ4OLIPdSOdXNJQ679G8Ip5QHII56t1jg3ROZ7A0Fxcn1E4ioZs9k
0G+rN9ZG5q6fXHsLq2MlROttTSYgWydkZPul0ayk5Ex1cXp9QrEhLmRPwTX1
LIG/XukKqdo9zxEVS7RGdCxhNTNQ/2njxA2umKoU9w/wm1Qe7RLHYaPqL8e9
64Z4P2V8RCLDzcVyKGy35pw1pckaNtTkVv51HNyoNVs6j2rYH25Rr56f6EcM
L7qQD3YgFm6I+INTXkfxshv08Jxe9ag89EXuIkMqm71kQ3Q4IDz7l62JIbla
GrVr6J0MqXipXvjLgJoNvQD06EwcMZmhBMd1ceNf0nKZmKZqUrJ0Bctenmkv
QepjbMSd6fWRPwWXJYgjaF0kZ1Oxs1WiGf60IS8tyQVMod3blM/M6qIoDeeQ
dHWPppI2FMnvOIBst3RUWOS6wNJkMax6wPMaW74wgadccrmiswirEJOD7IAu
raTgllSxVIm/pKevHernkWzscqSrVozwguBDNLDDniBvcepzt7P0HwTofODl
rCegvxJE03vvHSSEE6zdoiQ9FXih0R8CL/Cx8JGd+ua3xiCrvar3IyMQ85XC
pH/poPbpfef3A5fQIzosCxTXYhWmGJOvJ7E+JKODDm2GIJYOx7cyHEoCe4LS
7mQoUgVs/UyMAAggVC9cqw6iW4IyK5vXtdSzfciwHNqnxPOgcmkDxUMsNQ+T
e1S+gdzNiAz1dKjFCtKBW9wjRJLNQFtanQDohVYkdIn/w5rwT4Dy6Cgi8WjV
X3HEWsV2nW/7+91WxMqiNmadoRGeacjXQiSF1rE+IRnfuMyXeysTZeDLDNEn
SlMBrHF7NKuafSEozYrNEuuUuQuW7QUDEqaqJjaidDK+ujU1WK158Rimgetd
LwXWqEBFo/7YVdLpIG5AIQZPsjhDMbvUzwACLfgUCnArozXTkmYXFLut9v4I
fY6a0lFL8++uqhNDrcXfeoKH5h5AGZDE+qp/Y4GbsntOhGrNwhhL2LUy4ypz
yKuHcy828k786AFzaZabr2GizoqdfBQjE2bh2P/AY5MSAkyTgQf8+/5JI5nf
Sy0uxShD8kSvzL5Wq4bgzL4Q7HG0s0qHrLPAWEbOYs641iqfjfHbBlsAx+BZ
qpjW12zCfO9XHU+VaDgqX1OsBXrPMjmiKIvh9fQgxiHLzVnxX0CYy7tVAni6
0KDaxCDxwTSrFoLpgGDauAp2ex6X5cy/PVYh3rXXw///v4q3+NRWibZYTMba
rKVTRkxExxKjJNNkaDyalkkaZpbeaWxVfVo+1iTzrKZtM1X5rGn+5/6cgf4W
pdzITEDK5DHIk4WX07khwHy9uT/N24ppF3rewKC1XmRF+ILfNfiVuL78Gr2Z
q1RKys9fAc83iy7bUiiaf8Annm/W78OHp+XB+afh00XXMPXkyO+4IUEcMZqf
OJzla/mA/TsUNanAyPV1SrE496ds7CqlXOTVao39aXkZ/DozP9sdSiKBHlWW
jo3gUBbeNxU6CHX0qw9WTiO7le+TmJ3hFznvHL2kZWUyYZNc8tsiwGGoEFrG
wI/vba35P0jjfOztdzyyZISggxRFJXItUrCifIbxPfSopSjbaUEt9P/gCzG0
DHyzEgdrMsqPhZkV7XLa39vsdlO20ZzFttvUnD15XxYPI3R8Ol1NQKuPCwhv
HRCCHvea73JLsxt3rfMR1lJz5vQOaTVifV+46IzC33Hwyez0UHnE0Mbvfqn8
uiSAWYg9ONThKPfRD9+tBwNWxwAoDcN02xDl3DQLLzA66p7vTd+YXh5gJjXx
2+8hE99h6XqZw/tnRReH/2+rYJsLY/6/wMIzfqn4wfbTfCHz/hYeZPm0ItrC
BC12HvqrqV5/iG7WzXOTKP0mGPxksQB6AOKP0G2/OJ3EmsNkQKnXqaP5WlIW
ev2vQw2+JNaKSaQjAEK/KEVD2gsi/C31m7iFG9G1BerTNzluE+nSdMKhjxHr
fHq0Cs0h6jctbwRCYz//Rp6y4tqjb6ybO76vghHcTPpSqJl0vzuLnS6Bx5OE
OzwO8C+WaNJbx851T/GljBPGdzCT8IvCoxC2our9N5xmzRXY7wc9L69NtV3I
qm3/IQlAu0BS9KDFEkKQlL5msxY9KCzLZu6BL0X1dpcqngwe7+WypySETygs
04w3qy5RdtSBXmGW4qTtFSx0krPgPrvOx7kU6Wzi9FEoAGwwyoUvvtzlzF/O
YHrXjendiAuNKX1Y2RjC3dInW3Vk8p7xxAjc/NZ+vKn18TCT8uQjsLqcZZ6r
rVYs6KzkH5VWlRLKe6cJzoGlxI/BjoXzQwVpVITQkfHQK+2gjo7xJdiIn/BO
Z9x2uIQA8gW7pN4Jfscplv6v4AX7ABEBPGUI0TZIug3Aalp8wuomYCRlGEA1
6ZnfPKF5N8QOxqM+hOEjrwmSfrl/C+A9K89b3VMoKXsw+2J1gwyEnCqMARDr
poi9zgjhGlw+gBdSIEcuJZTllMGw2tDLY88OZFwkBNoEIQ4u9riGrKKmOzdg
FssbpTzBWxVKs8nzah2zwypHOBgK/DxykP9emAfTr01UkHtngWFUq3KetztR
0QQrcN+b6H6xA6jF0x+jUhm6lllJm4aaxw7xwJAp+JlXEPo/uPX/M6/d1XOD
3DHgtOk/AmpJTLCHu6lRHXms7XQV2YSOjPr8O7oL4fB8L2hHJqpI1avvzXve
IAozgoz4lBLI7bczVOcyqYW4pWP1HBH6mtdffosvu43/S7+GPodW7wPJFOrU
pAhJCQ8oK9AhnGrYDCS7bZUaW/pYxGZXrpidtnlPND8+WXM9cf/PIXd1ISUp
8QUQFy3Lo9eKcmnvLy6VQTki+2uTNKy0xScltkFY0mog4YSEefqvuw/6fr0Q
813lLzaP1koCixnSePFtTVUAI1ZXJeFtlInYsET9QE7H9opIUFQmhQBA42Jo
bewLHDgTmMwnS/k0aHXMjFRQcoLXT1R0RFyXMj7hiJV4g8USbG5eVq9YkMaD
nASKsZTtzrHwuJcXwSGmdTMJ8I7daanNaAUvDDOKfILRNFmICEgAG2OklDit
MVCQEhQqOn5+HAuHArf3BpSjha+Mqb1rMPTqMu2yNq/q+KQ2M5rfdp85a4VH
UOQeuVhbTKuaDZKQa57kyt8Ou/ME44SmQOAUG7950fnNQ5DGjlwsOnHZoBig
wQQ5r9ADPelwQIRLyDxtjLvuLH3yZWgT3Sj49yo5V6yPB6DlWxwySgXBt3VG
adLtKW9yZxcW2SUKi86C4gEZ/sLZtofLv/qgBKriU1ePxrSUDDPtyemP2oob
cP1W2dLt56Ov7KdeHdKH+kb598xBFOiqnWqdc33tdrD5KFdHrSDlwxPMoR+f
O20T1gSPC4yz8GjKCVbR7qvOYuZRYvxk/6eLwcBw9sBCe5OEEYTXzK3/tDj9
2NPHUfQIpTF5WugBMJeq4oNg8jJJeTtp4FhTC7NCa8xbtUwBg1cqxFHit6UB
GtFHz7A8oNTPOW7FHUVPmXnzMmNdHlorqGNcxWAXHB/mnzeIqZM1S4o5vBtj
uYvVSsAfiTTWfLIVQSGkYUWYg4QKci8RfaF1Aq8wt0gulIPW6lSEug50Eu8f
Vc4Swe/naJc6ESMsu8REjrIBhgkY3obcvld1qxZ7gPBL1X+LA8inuhm07wUI
KwWSInA9iqptsOixRSELE58A1iu+9QLZFxHt0jYUXnc6l7qke6jb9+RKQj/n
nns+hMA9hhjK9D1HTGo2R9UcGtTzHEYRoEtq9Uvveu8fwquLpYQmZTgtnLc5
1jtT6DmPCNcLxrioAx44KrlyJqdRb1O8v3UwnR2ncAGo1gIM5FchVNboNhze
xLLqlnuiTkGqrNzYpkqH7K13Sjs7w4M9QJ8BK26931axR13IMTdIYmnnUXyN
79ySG343a66kdubTqGBXm+nkdxI6raPH191dR6H7ZXZZCJ/C+vWL7LbREqPy
LT878bWbtBygc/u7Cp+UDhYQqi+3tn8qlGafIjz48m8AXZYA360ocU8zevWP
EbNrAoTRjPd3V+FiG4DmwRaRBFYhR8eUOCJGE7ueH6S+UwZMlUUgDp5sGCR8
syMC42jaM++CbAQfTVtNEAWWyquuGjJfyf7eOJmeRkBJgVypWMnWLhMi4gg7
pCGJ/VyP0hv98QoZpTEfwAaGjMVN9nZSzsYZ5z9RPbEx7ImmWG496XBkeTOc
f0x4sujLJyhCpnJ+pXeE0G7/FvI04UJmA/v4lFDcG/LHpviN+9arvKaM1fxj
r3N1zK6WvLzXshdTK4LKiG9EOEQP/3PT04QdtFx56ypNasJ8Fxa1RVqBjTVv
aSue+WftNdN2mfh3flfpT3lhj1QnqKu96r0zwr4gw2WDwgvyqqdAnA3kbXhz
pgbC34SiGNsAy3LNKRENHHigTjddZSqYW+O3MMN9Dtv/lyTpRdQ3AOebdyDJ
SeZAMloK7LPW6LkyHNR4rjHFbERPu5ikE0Q6xm+uIon6td7mLyty+49VI1YI
nPjfBWjXnE3MHSs+Pyb3/pFj9djRkqJUG0dWCFPfrat4FxJ68U43wUr183yD
CCzmFV4Onesu22B406jPw94cMpSO1yiYkU4g6FNSzuxllCuzUlbzQyJHVJon
c2kNR0EAOd7q8eku7nt/bPjtUMsijdv02bj292HhJpP1N63tFy9/JNOd7LdF
adiX10zvNh8w2V5BkJpSpOzNFCm1fuQkNwB48+C5mxRjOpTKF5bBAYJzshBU
W+0hR2DcZwmN6DPLWpzX8w+IAhdOx7VKxwjdf2ym/ZnuFHfi73iqReHXEV3c
HyjWIGMx6C32FTHg43qkLjx83Y/TewllfY6JjlxXcyAovWfiPPOW7qghODJO
GXR/tWeHBhuqVQpBoQm2sXsuIEtwlf3T5RzEDUQdQ34VVDhAqdazbdL5WGre
15FekvrzhNnLb3BGKX672jGXEacRD/WiVLl1f91P9s/nEr2SPQ4jptz0w2vk
UvVmvRHls+aJmGFsOxJId2EEioafr5NHqYVuiz4GWxYRYe5bcxVsW6NQqaKX
ZfyRFH+L5iZgoRI9oiZC2oidXCmgm/D6/aHNkMsWW5D66RbIx6RQ4EyOWB5h
WV5f5ukVYpsjpGRCUyCao1zLNVC8i3BKMV8u+fthy6ifFR8t+p90oZcC3WuX
zYMpEOOmUPArdzUqLi68wBsFFdZx4QksITCS/YvmRWx7Dh+vHeQk6O/WRtDj
gwrlHFY9HVfbQ2kbM3+t1zPv+gQQHIMNc1Gc82OQnC4ToBNJPQjEA+jjW4wp
E1H4a0t8jykEmM6fP79GKBeruY4HyheO5S3z8vSpg50MEqMTcQ325fvAkYaj
QlwK0bQAen+yW1Z1K8SujQbEAeWcM8SEl6ID0ter9gjFWa7U5+7k8sQr26iq
Wo4qTDM7VOFPJBFkmW0uPmqFoGo8hFg9WmfB2AZXkKraWAYiP4DZq/kJO6up
xL9QJu2XWFn0GQIutYRa8Y1Z1cqA5+fXtjlXx/Bq+gfCwY2vXQYCBxR60PEZ
IXQYc/PZdg/mqc1WWuv3UdapdgUd6WbErH2qF9wsqwT/s8URML3E+PUGCGrr
XeIwcQYVY6RzTNOIFn0aV/HLH8OEUGgYAdNPcHV8IE/LWKOO6x7ixOy9B/T0
S/5+S0X/OXLEbzTkb0mKVbGjas0NCH0ViHxFlBTw3QvN9d8sEsb0XwYbnttE
ILWndrfdDFP86XXBUpBY8iqBpcNfSQL0B+n09E9Vw50evJwuL95n/DLOs9jm
RlPSCeLJ/Ye/84ZRoF5lxjjZVNUoKpQ4uzvriC8YroS2P2x5RpuPnUZyK9xO
G2GG4dQlDCRVyDKIuz2jcV/VKLazXn5ZvrKMPUveAqQHhhEywMEGVWrCZ9Y0
5I+qevkz8p0uP+if4RM4Rl5gtnwkHLbunoGAaEIZauhB0WTchhl0VDamjuxb
jqoe6s3jTZuRXFzsJhjsqtXAUAEvERONCQ3eCC9o6ClbjuogbqofSom5UAr4
PjLqoUIwf/MmQlhJoRozjnDvMVZ9P5IWhp7UwdDFhDUj89bYJXjae+vi41IO
2nWrgr20SGXotEmLnoXfBY1RaiQVK/JB1h0C3FT7k7CLOI3U32Rjopb+G1dI
f5Evs+3lZsNVVlvtDnEhvc5QhUhHDItz9+B98q5hPy3LR0ZoF/8Kfg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "221cqLfSQtZLwpVKjUxAj0azxWo9qWyTHel1yyBq9riDaTa7pjyEaEdGOLLz3wcrK5rHulca0g1g9Zlx/VJp3su79bVOdFJFOSZrof0/9wf6C4nAWrw+2PgJSzMMKpaFLO6gpDFruW5083aTh1M+Q5KnW16yLzHWGhpxtWHi5x5kzslfPRMwe4HyZUYh8/FwJanr1Um2jvkSaUjUKvojtHUTdbUpkWg93bqHvMIamsncpBfseSGa8zqZ59qzsXxKoiTVgdeUr5Th4jrjrrxLu3ubE7mkwL7Aee4YiDISphZZ8EZxzDCR7z427GFo+6sMdbXSR/A+yR3y4NxyNrm7T5x+l/4AwT/VA/4HntwT8O5e6r478BOSRyIbr3EV45bgHjGKjx2cDDt+m8PCiXiRkbSAYcRapHB994+P+7g6k2tu1Zpdeus2XpvJNWuwqC0Dg69MC/JOJ1ZshBL6OkdKuu2pn7elccKzQpRFZ1H25N0DqYPsu4ZADewiRNZbB+kdMcQTolU707VQZ+gk8aBu0t2pMTpKzAHnuouB0MZACORVYydtN3OwTyaqAp+DjDw9foUDf9+XKZc0n5hrkpgfxD695Tqg0Fk+wz//MKN9e4IvXWe4X0XbGayCBzkL/i/Ez1E9pJc/ErsSrNkKQ/+4lm4x+1HIA5d9IRkTJBiZflyYCzMIhB36MnmIdPzsaLNIiR/BkkBSgTC9XVKmyT2XRnYf99NT8pFnjgMJ0KrD10EDW28ACJ62BfYxn1sm0mRAAwWafAO0wq547xIvgahOMMS++HGXpS6dYwj10S88lSa8krAZ8haiuhIcyZ2DjKuBWkJaFKSNHZQ9MAj9kyYenfyMR/M4QDtwDhDWtJXdESP1llv9VBLsYj1Kv2Uzzom2tlWjiIFW71G20a1py6KLrv8vl9NhZ+o2dlicFdV//24La5K1SSc+xdX7GRPqpJrE5iv+FovxMzPkh8onck+TIrvSqZQ6sbXQHHXA3IhJaN2mFHrv0Asx9BjmrevRNIie"
`endif