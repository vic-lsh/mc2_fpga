// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Oyq0KhNjFZMoachcb+oafZjqEioJpGhS0k6v9i1NO1wZfQdjEynapWiM1jTR
KmPyk6isqDdvva4U6ZnkrQmXncKhrb3nCD4T15jHM5XxRz0exT/rY94YYMTC
r+jO6ZE6La6mSEGWotRIF3dS67Cq5sljftQCuXGB2ODYhhOoUpIlwWWpNqay
JuBIvOarcPWFsDOjPfJj2WsWjvMoEUPL5huAPIXeKZ+8Tj/FphElxdf0Ef7x
SHWh7pHYa3jhuA42HxKIOe9pEhZc5ZaVX5Cz8zgG5837I6psD3nItdcc1Guh
XkTTJj8vrVqnxJu7U060Syxw4DSM/QrRKY1uugqmyg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HEchtZv9DWx4K2UiIRQRPBQaZPMqoY1sAEzR8GEFL1dYXzxCE/VBTxTvo8bV
PrfRQxVz1ljo9Fz8TQomBEQ22Lzb7gNxJ0ucWQplMxiOojzcOJZYjPX/5OnB
av1IICgvjFSHkdSwA06ab91rDfxZQzbXQJ4j8Bv26UzN0t+mks4j/K+eVswj
wH2kImWeDrDnsURK02TYlUo01BN3eERTeslq3juy+PDHN6ESpTByFhXLJo5w
YNluodelTwURt46yQ+bqGT9cpdqMUGiLa0S5WmF3zzopGgzVfYxJaEoFqqY3
E6V1lODhXS4UiAZ7geVx9LQ6onV3kElGfTTnlkGA9w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ihyQwGmzrCKtPgLwaB3PjZYiRZM1kJo37vH/p4IpVZ/sJVzfgBdnt/iwUKSI
h4OZLyUl7GHYb3qtsMPnbubF9/12G94NktVg3/ussbb7mr7UbE/mh2AMIiZU
iFxeul6tNL2Q9RfDYu7X2nUBzpNIN+la9+zk/+7uA1LPdcrF4uGqXWe0CBvr
qONklqlp8yu2kTytedxdLni8PjJ/30caZC/oHjZ9t5qLdXInviw9OxhN3JX7
RcsaBVH3mqQvuI7E8GbV3NuJ3s84Z1FOgnAqlh5CytoFkkANeQQMl8cjV6el
cUJixMVDs/wXoGW3Va5y/ohksDbwDOT71uzSycX5eQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l/rYae25yCXklPHAs/dBdNkz0FRfLvp6l6GbBBZ2q5jDiT28fF8h19kISl+t
l5douF5qHM85T25U+q+AL41YulXOT/0Xakl5tADvGFj2BMHRpI8qJbgC3/U/
80eicCkuquIiHerYSc3oJg4UXA8CATGslRj4UXIabTJuSfP3AygVQufxsirC
ZR1MHQjNlpQZYuWxAOH8zBBqF3ESNbiXtuM3Ggln5JBI5CNPjgpfCo/Ylufz
aV5L2eBEzygq6cgyGUd7guDoy51JpoSlcc8I1RDB5xHfDSbpWkbsedGI+C2X
W+zIGBPOt5R6b1tM9HlwlXtYABD/GxORwEFfLP0t3A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a5RPc7TKk45Q5fOIahe8B+3GwkPSdUfaP5p9XQ4guqHn3KGjsa6CLIexgQ0C
CwV4d/TNqaOnw4bOvGm2e89aEs7PSe7d6dX9WKJcMbmRJTAOqM2L4sc+FUjd
JIVxKk8XEGaI4zOhFzYk2csavmGiB/F232ZPmocC/CCvjDRLeF4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GCUM9ct/BOcroPJv4F+LliYnjwrTGMxH4MfSNOe2BeWpGlQWErTbxQ+fjg+j
s0h8DB4kcIwlv43/Fnm64CzlDel/5uBDYExvespS6ao2LpxAfH1I50Mxau2l
1TOpFMzu9b0CZ2eh1wahg9Cr5qCtjzLflPWNnOmo1QECsKTuBYoWGIPdb0vl
jx1xaccio8OI3fPlL80YU7649flEzsYamh6YblmdW/weoJ43LdZUx55U5Jsm
F4ivk5cN7H+OQ5Y/yzF639zlE651UzQ7zHQhZqVRu+fVAORky8gfXb1UWFz6
fSEuGCY9MrBMz4DcCiDNuPl68c4dQuPEayPSvmruJ/LpkT/FD2mFd+2liKDl
l3dhHxXtAng62plJ830035QA7k4DnCeq8cq8y5ZLBGK0U6kJqrd7FF9svVIb
pDVD/jgRzrjquEJuZfzHdR/wRyk5q12HZkelQcmkCUIwrX2S+bR0nSXR/UAt
B3UJtDmitqrC8AR6e5Sw/7lzYUr351kS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PuF5CYNUdAw91HLTXBbPWfsDdePg2YLcn150IlCnc5sBbQiHgFphi/4kKJ94
eeK46YkZDU5ojXEQkWTCyALr+oVjZx94lbu5LlXuteopWkcnLQgXbxz5pM+I
At3Q4DbP2AAl5joFRlcrKOxIvmAxhEvnRZJ3ONlKDsFuGQpG7P4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hYe2NtmV7HPMkrx/+N87nwmAHLwWKcAYHHrF/9glkyl8JuF6k98g1Z+TZggc
Ndz86Ai7kF+cdWE6d9GJMikKTQlfEsjjNtrPIklCEDxgBPaCpZtwWTM36qSy
6F44fGAR9v1OS1i+3nvFp+IzvrL2oXK40ef9bbgq/KU9VYj6DRg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28432)
`pragma protect data_block
dqg9H/r4VjDgzKO1XcHa64IV7btf6TMHagHEqDoWemuvE+ZvUpEmtXzTP6wR
gORCl1ZwfTGiF1iCg15CQ36W6u9RfH0LMrzTxZaIe5mTB5rUJdhwhdDLjQaz
Go3ZC2d7Z2pTMOnyuvOhIV6cRe6OzPgPXnGW0j0C7HltGpALkUAaW0CfrFRm
nepXooRUWrKiJTMocTJeSWnp0W1RTT0Fi94ERQYekWA6Qe7aBNgjriA+uo8T
zmPUnkxsqykz2tv1vLlKdhgCvht8yPYfrOk3aAC4SO+7mU3F2dn/yEvZv2l9
QIp/lLIz/wGgdJMD8woTqidwLtHwtWV5GLOUZN3vI5hbBgOrm7Cc/ROAN4QB
ys4g1LcR0e6HmtQPvG1hCEfL3E8t7RGPYjnPJciHbqVbQJmUsG1MANEdpeD0
EO5yBW7E+whq0eJipFKtudhZlhhQC6wu6q+v7PK2+gtEyVD0q+OLF1eMJPar
F5d9rqV2PbTbxaG2zfRhWHZsVqo77tglj2MBYJI7Od5x9rVUapoSyedtpF2I
12Mlhz03nISeiKswU2GgPDf5kKJkL2ApLOHF8LsIZ+7CnrYs+7CnZxgpQD2g
h2xDG1xv7S0QPzcWAS5V5JFGk96LOq80MaC81meWy/wyxi01JQBHroe3zapH
JLlaB0qMkUS6DRqb97LrTh0UW3qSN1FohuqfbOkGxgaTRscdaWpCok7Fu9Gn
E7V5G4szWAwCZOf7pcklxcR1z4KUeYhqJeOjqqRwHBfdWErmifXYrPaE0E/L
KKVec/jFWCzOZCDszDhip0BrtABaqiSq2i/ThLxxBEfXyADPiL3oJqg/RXtN
Q0S0ThrV9O7oEihDJD5dClqvg2Xx+FkK2fpBmNpQ9T4c5uSURiwQpAcuEIef
NvhuzydEcLS7xEQakyLOhxJ6JApSw0z5nBt1U4CVGU9/viIF8KqOREznm7N2
DNh4Jy18rAK4tkEXGsT4ho++euxoS6BzL0AYFBpldhoVNJM8FjOWu1Kdze0Z
29qd/nqkU7QRUXk/R/qSsXrwcKG0sHi9gDfkAtCx67NtIZGOL1DFch2T2fht
ZUYUaSrBcA9RV5FeaMq70fVgmVegdobCZVxvuLu8R0el9x2tqrjX1BLdXbwX
lOnLuVnrFmxzFkqxqKMI5W/dS7tnBlzBfNgBU3B1Y7xWKe4ijGv9QtGYMWb6
UJ4DXG7B8yEoXJD8fmIbNbaUNxjS3ecz68OIw6QTZXX4JUrspNfF/Ifeq2sZ
KXC+Lm3qipjmKbOGwK8SwcOsjsHhlFPRK/du7UYWP8xy1djkGb9dwHoTJbx2
c9LpHVL7R2lYMSGEqZBr9N90GEklKIfqYNTSMNKnJLlgqa0gaIBBFdz9rO9m
Ylkk//PbixNFEgsTIX/sNZOVi7JSGUSisNw/eGGe9jRn5RJJ0GxnLcmDgi9R
VccrOUMTUIOXMyjRquGdpKDvOzl/LTIbBCIO8TILFVRf+a4UFSJsE3iO5Gzf
0NGo9RxtVTT9MFyf4CUA/ZeHOZwzN1uA8bzhWf0wmtAlO8DBbUF2NTNi/Qag
1qedVltl/j4iOBcIwYuYkblnVhc+yIoTi+gdnn7xDUWZfTpk88+1s4OX3ajC
7aLsh8T6C84+GFE4ec2AgDIvbiM9x0lD3yY4/23cVrloca22w/q4EQnyZaFB
BEhvfo5PRPciJnhbS++Ix1lwXBk5TBffe3MQyiU6xQW6ibi3r3cIPLXPZ89q
mcxlY3K6NljxDnI3J5A6UmxU283UPwvShpE+6L1vAq6Ez5FB/vb10OZef2M5
++zjsHuE+v6I+JWzXN5AyjEV0eCGLYWZiWPcEZQE2ByVCHtXGnppJ7Jh/hxo
VFDyUkJ2jYUNcmfPnWKzfI9u6qR3N8i9dS6C1MS9cJlJ/toPVfjxNaSbgsr6
yai1MyAMnJkwdi6mjyXiRe24VfN5caSQ5hUDpDJXSPeAWB6oEm4K+eav82RE
xJ0I7dBqYG/9gskuEXJEDpae8JAfGdeSSu8c6TjEw2NxqbDLBGtaG68QIdZP
GZnzTd/P7hdHmumwKhqADotkelpHwBl4AGvFaeJXQFA99rN6s7OEiayEh5sI
n4zN/KWzYSnvs4BMDmEi4YErl9n1QkBl3YP/kYreEtMrE7KzTk1azc+3QVYH
UKUIHI0ahUTIE+QBx//4rF8MmoxT9RQ14ea8rW2tgA40Sn9BQkzCmjO9IoeN
i3v8ch+voPSEmxDuV2XeGooFEpbJjGt3N24ChexYPZivwIW7Q4i2vhUuOSfv
fTQExorgXkn9YN6HoQFuA1oaDE5vWNtOUnsDh/EEzTOy7VIamo+OcdmBHV3S
vXov2Fv5aJjM7nURvIDUd1puJRbf2Sb9xcF8/NPaaCUG37OTP7zIdHHlpFke
MCSStUmxEUcMH0JnwA7XoOUJA/BJqx2rhllLXAjpJqc5fBTAVKQDtv3ZuQhF
0gIAB/tw1KZb2DvrWLBscINMgECYpdAkprb5OIYmkF0iFZOmbmjpnwtFgBt0
kb+fuq9mAj7F6wn+5B554sY5lIq45SzmXHnk43U0T5buYWO2ZlIzGz/OJf6h
b99RqlJytqW8HalApxRZVo/3JBdH7ughLnhs8T7Kywd6Uc7O1fYfwF+BMW3H
tRSgs5/u3XctATm5UBWZkvm78rRx83uyy4hcvNwJQHubJfa/RqCPqpeEPf5/
7v7B39Ez3/WUHQeFEP1N7Qw2xRCe97JSpuBufA3IiovpvqZXohR8kSVszdRC
8dTvuXj57Yl/5/Pz9UpoCx9ce9SUZGXMkNQLEkfn3jqsJi1a2UzWYfw27YuP
yHC/jJkksGgYlQB0zpaJQMfHaMUw8WzV24pL3ieSNytbISggocsUmadAYB/s
LIhpsdZVkqxqFkOJdJa1ZsHb4U9oDaVhaz7a0bTOUzZorNZCXIPi/BjP8LGc
KwM+UpyF8F1BP4UVoh2n03E5kG6/0cs/CUNALWQGuck91DyntID6FIRcao1/
/k3icsAQfD8WNry4Q1Ynrd0XnnfWp5ut4fX+h86RLJIFR87LVXlfLRIe1FLL
61mVEtfvmnGt9VymC+C/DIs74kvHYpKHUl58pTaMqu9g8cFcC8awZlKAi+dV
Orzg6Gw2Ccn4dGi/TbMT07Nr6eBOjzEala4sZC1nbPBgck1YvVLkAhokrRRz
2plr8VRBXc5ko3qV1AbVuja/G2jidUaz9EgNL8IuGQJb9qATe7a4awteXviW
Z4gXdvGammJvfSsX6pRe9q7aLNttSEf6rVyM2poU0okY5QWzNiP+XwjegJmH
rpRqH800v6TUm4SGGxy7RKqPJouUmOfYuMl+Dy051JAXYFQE1fu25nws8W6J
JDYKDqMZKun4Bv0mzaxxAxfiudHBghuOdu6asPmyptP09H9QsSspDH2+AGHX
l67rgOWfIXPETZx6tDWVV89COEC3gYA7KEbR7no4seKEFi2TvTo++aluwaYo
Bp1y5BbG2j9WsRx/s+OR4ddw13yKjeHOZyA2iSemptXOABVWgj+ZubrqXbTj
AOmLdOzhRlLLKzXxmJwvsRRA033yMtJjaBixGcMMUeXjUXRXnjRJd73+EdeF
IU1x+32ixhLOInTEoe3aWwpk3axB5KLFpPAQGj29oL9vPxzpNyVX23mYDJpI
LLhGP82Qdb3Md/hSnGHqxXMC8g3qb2kWgdCmOye1c9+dwdXiyO+oJr1ui3W6
B5jnQ5xPEBXtF/uCaR5IJ+rviVpkuC9w4BuPSYaJtK6dIxYXKtNAtJo57z5Z
gLAm2UCwGx+bbz9rW0Q0nOMqICm3W6wsYLbFJILGMgJFO+l+Wgu7oHy4QWoR
FIrJHUPtA2WWjU541qK0UH9mLDMnbJ0LyNU3yLaMOflm4hkaJN72MpfJOW3O
EI46uQO4+bDmlEcF7JK2sDsXE7ujGm9GhgB9mC3hLaFVq7MWz/R+Fvi0Jk2x
sPAb5OFGnpV2RJ2sD+vPu7BptGD3THrTeKUXOBOVmO2Bq79tD3Pei1/Ljg4F
qTUc+3sqHZUAnBKAahNmULMx1EbcBOu6bEavsNasu+4dUjas5L4wgOoGN8lU
zOgGgBKuV3YUBWZ2nTHkCbhME0swRNbJARgUrcQktjzEqV0eJZGTxoEwXfFN
cgv+PAhB8jrptTBJ5HbF0FSZJsc/HNw0WhWslsWhuZ5X6eZ6TLkUHIIDUg/C
Vov4JuhzVGXdRETxoVR3MDUF+YM50u90jnXp8mlFgMrxlOF50LmXP6zCC8Nw
8Kv8vq03vSiHcpFLgJQOlmsCONPvVTqjT8L9vH8Lqh3zVJeUieqom6u/G1Ir
6MwOcAeQIWyc61aDUO5cgM4G48lt9CazyeI9yZVQtPLSGtXw11enZUcS8xsm
GKA7a2TfjG9brfpzvV6SYoOiqGMvCnK30S0E0qzukSMaoY7kJVIkYCcIGe6Y
9n0+5PhOxiq5nO25jKj/tiPtzLgXkW1QvV4o6jYMVNhIZR8IVQif6zvspqlt
TzaL8wnaToF/2vALrrP4WcFKeTpL7+k2dyD4wNWFLQdfUOoEyeaXHCymuHkE
y/qy2dHaoAua5nl1JenQzEUGII0lnBtF8aFYWJSXHr8fh6m86Bpy0nvdK5U6
56Uj6ccGmwgvn6in3dXGIBtGm9gwjKmdaYAO5NkZq5Rs8kURdfPWfjxwgEN0
4CHo1Ctr0psGI10Ykrc0G/vbCHmkNwAGcPeTZaogKqGMg2TWBRJ7XYy+3VSS
zGeSmvIODtmSc7LS7EJCFICS4BWd09wRAVcYPWYQE7JDzoSlVRG8LtODrphC
11l5wjADDCurEY61GGEXr7Uca5YkTWvVfoNoPGVtEEH2i06hyle8IT2S/pf/
ej86j89akh6e3Pi1RlqGA8qD/d+pofkKY4LteWEaPQjo7FGkCl7xLV6hqn+b
n8JOyhw2JobHeIAyEXx/1LWIOjZrBeyVvbf8TiSicrVzDiC4tDmpUmVdkmDu
2lMpmVmSP9s73LaR4PZOi/W6X3Bd02uCqbn4I409VgJjI+C4AK6wTSQkwNzj
MT4CKrvMMXKsaTjkmNJZiih8SPuzdllexdR1PYSG4xD8f6ow9+i0m52+JUUG
0B/A8CewUJbGkcPtbQZvRnGQ+kSdE4d+ep3QYxt7P9jNWtj3T2XS4ao1IIao
DEQ4Bc2Islgch3WWS9Bcm9Y3m67JQcZn0jmPZrLBOdNsGozhYxox+R25Il4u
sS+rIx1suI/ttjVeKXQsoU6SdnZAWS4wPTPyraFHTCenuLUxN/L953tVHxHG
IYRX2V4w7VWdGFARj6ae/MDLSwxzMq6cIno/yZ5P53Uh0rQObkzBplDyXZ94
GMBQOUCl94UUL0GIhwsT+wKrpQwBKwU2w72PBS9XeFkLr/hNsI4y0/0lLCmM
lz7JR/A5KzL7OF48r/73RaAj714JtQQLjcO9QrpLYv/MT52AuT8YuW3YH7Yx
QTC3gD5oFmYdLl7i88JB8r4QFk4VvAm8xvSizt7kmBO4Ohvhzd6WYFMCyQve
mVjs+kckCj7qr5OwBHIJ9AyH6wjPXYmGS7fDI/qfUrJGZcs8ZZMrSChSoSxA
UxIEa8cZ0LVQY+CtDk47s7C2Tz3sTEas5+/ytqXPopjQvG72/vTJE4hCafZr
hpaGz8viSk/rqqet88vIWBUhQAXW1JEuDWvIsOLq7Dg8abngfkL8tvm/ybV9
LYg/5v4w7WD4XVjtFclaINGpTHpwKsZjFe9jBlPL4L7Ggjc82C7ZGvvSRQaL
+XQhNv1lICDOGRE5QTQK8Ruav9olalXWOFEdCHBNb+atBmyRobWw/NkSbzfX
SI1pooYRJLo8mtSzeR5vYAXCfWgFTVlrRK7pEVeN/LjVGpFSmxoqH/DiGg6M
GFjh6PtwFrejqAZf/1XoXx1U0++eUWrrQKuTkLcOkrivotTwduGFiZInOY1j
a7rieCCGkAWrbTLjEnIiQzZFP37Hm3ZnG1uwuOy4Mb4nB4+YK8sqnw+0x3Hi
V0CmrLS/8Ef3WSv/vPGcvKNrn5Jm40nbXUmVL5MYXfSQKaUECS0VNjb/FqMb
BVMaZbyoYE3AYS65ca5+0xjBjoT8pUDFG7l8Lg+S6hj08gBBRXTz7yMZ20pU
IejeTFERY2Gof9Togil2QF3zKbyS1Sg+9WUmP9vGF0qET62BVoxr/ku8qCEY
o0y5yK8Uk0WCLUFkFU772F4kEzMcyTZNxgQeYKMLYsyDNO3t/qA4Y1Zys7Up
lHAqrtYYedHybMZmZvuDywdzsOLyeydOlId25133C+WBiFvcdPXxX+UfSIyd
WK9D5rjw/KzBR9pJaOnrXYtIdL8hnFzUJyfI1D8bGWQXVqXfhNY51/MC1vwX
wPqppOvvWNMkkuqTgeAXegIlI6IyvvT0NF6qH4IBMzCxLMEvp4tChbyOV+gg
9YoS6YwF8kG4V4KVsZftcygNoioQSFoBtGJpnTv6mTFkU8YFb7w+8l+583ze
nd1wJQFKRF0PsLKxJgFXTEhrL1jHGTb7KTHYjEGm267JTpHtyz0mDShIMv82
eHk7ElzhtrL3Ahr2bt4/dghNh2/fIPrlL987sW1budj+QuBjDFdOxi4rCux+
BHYk6EtDEBpPf0moTC+MLxvdynXhQI0XXrRSkLwBSpmbTXc2GHAuMyKo6yML
boyJ7G5KkCA6GUP8sq+OxnPyScYPI4rHEowF6WtSUm7YbKXRJXgEz12UcF1q
rWbC4Z88S59yps4VbGxp8GoH58UIB5D/o21bSiMncOquwadmpAIYykq1wBTO
WlCWcPRfGHUCXSCOfpt1dhx6mh/BLnr5fbZyMc3DZiMNUE8NA9wUjaQCXbsq
KhP4/wu+Ms8v1SJvn9cGb53ZsmEhJt2LE+3MSl2VKWUmjQnjfwhwz4gqgLhY
HRHrf9bh8cewQKPo9btMUDNuopYSkXygda9B1ocXxAIzY8DLQByQTdgiPQoL
99nyjS5hgZpE4RsUyhW1ccvOxVa0V7u9sGaQMuEqfrR88IoZXuBj9dQvXu5p
sbu+6/5HInGoaTWiG8QtcC5T/94ZdPaXi2Sl/y8HjRoJLc46sc/UCtGaHuzz
jMTpuyFqjGfPd5jU4W5NUQEyw7THbmMwv6P1lWwO8i5kaq4SF9FBZyI3hnVs
Pl3sdVzxOccrC9lRQGPs4qifKqB4OKZCTUA2soMbpwor/VfFJZeB7NzClJQ+
o/w11/Mqhs39cFb5Wd1QWWglwB+Y8e3Hn8XhhcrOZKe8dEWAnehhZ0iD3doC
5fGQJW1YnvO5nH2gSaOm7+WFFDpz7N/PgNGruQp/xML/vPG3jFRa/DcBr5ij
Lq8nYNrdpjgmFJpkvF0KgHI0jxYQfMHcTupBvKnlHBgXyuJiUWLMWr2maDWd
YbxUg6S8J+flkjGWie3xU4VYjycSqjOiOqo83LM3PWBoFXaaWptdSqkznsoR
QNTQGal8wxL6PT43Tq3QUYdqXLFjk2nk3y9LpKceGFdxUIMx2IAPd5iuD6id
k7Zungkin0wXXH0XZckJyMnE7w1OGAAeuWiQYWLWI0tN8sjCRqB/FaYmJ4od
DqEV8eRtoHmaahP+bDzuA/AkTp8M0pVHGEmgjPlzbTBfZinmxSzm4gbrFvP8
F8bDnpVfZ/g+Pnv+bgbo0MpIZSZjwPmnrrmgQvoHY6tMUOBEgW32qjlN/JU3
lLdMLirxp/X7lxqGUZK33OXePX8LapUdIzpjLZ2dIyQQobnIw8VI+WN7Kynw
PMGo62PaFDqg/gBUAofFWV+TKVyR7q0W0Wb7xe2jNAu9nQeqtbrISkqkm8CK
diTDlpb18Gm4q1DGO0HujvwvHtR01NTLYXBjXTxASUV5gSjhnJxOq6D6yUot
jvA+iD5mQ9rPwEIf1TO9WeE391KUi8HKlGfyHRUQYKurBme5QnCxNSeQ7peJ
m8WnR9PeHfpH+a0KIADU5EQpG+Mbp987qCTfDrfyRmUUpYO+XMmy0by/Oknv
Sjy3crXXhqE0p5J+EH6GSwcFhV8cz+xztSd1gdSY4ElH9kfyU2jth0x1Qrp1
IG4kst/+g0MT1HfSCNUaH9pQQFqlrcFQ5NFFQku1kTVYGR2o3Vm3/6k4RQWf
luZPnjcIuGBcM0Ph4idx2xtgJBzHr6Cl5JZLoBYeIt+Hsk1ZCyJPi0S9yrqE
P3fuBqcMZfvaZbL7Am/T+2G0EtTjLN7EFeDiJ1okVjDtZlNpYE+ySNPuF+np
kY4vWEvASs8IEErEazU0keVyg83TPV2VtoKZL3KOssQBckAw2jIwRWi8o6Aa
kBPmkPPK7hWCCQOFchROPE/Ae8r+5dyFs4C3tODtc7oG3QjjkDftEuCCqANb
BBFywv7V16T/e2eDHSUjKJ2TyaG+mxTe3Xml+Am6rTXmns8uIccHf6w7gYE+
aUd+qa86eNuG1FZtOjldOF4K+8m6jfZCd1Mr+JOOtX0gWZC8GBSjjllpkc9Y
vecEuxR1tprbWqbQifahRlBbc2/iMdyCNUaKFrFhUF7jxL9VtKrV6uvbb6sI
88W0vZH+/PuQBeX0fZ4uoCJYknqDP4DpAS+aaNisDfFDNeIV9ywhsHI7jDig
CK1TzOFYHQabuJwepIrigEoPGlKtPqfRy86Lkj7tcSLsSezjEYO/+kiNCbNl
LkWEM/sRgQi16RyPpMkVeFEZMY63LQA6OCXRhoDwX+OGggkoE0FvcNPUITK7
xzM6ntGOF8cmJfOy3YyZYf4hyheAhJvRy+pcFmdrVDJIlcA0idZleV90cD7R
J53utHuOVFc2rgbTRe/GHCr6ydsRAAONbHsrdHxKuSPBjj8XzVeXR172zDcY
rGXhoohIIgqwLM1b8/+/orDjQFs/TDhiLyDkfnhR8flbcspvCcF2624PmW7N
+MWT2zIeR/bBaMiOZ5pB6w1+yfeTWg/wEyFe+sGQT2IXXbd4cfwDpetGtoMO
lzUd3yv6LN4UaDbmnONNxZOWMuj0X56bYkmfRvkgw6AdB/kcEbiiAmCLsPO1
sycAvzVVLSPxafEEWJZYd1Y7qzpo4xmYovKZD3Kb+9KLAJDBPaREmVg9AxSw
rX9IOp5So1iv8vFZLiT+Zgb+QxUYZkMmak6Uqnd+Oiow7TiTwNuRMs1aRAdk
2DizQES0MTRDGUuf0L02+/rlKdN3AiZ9SHOJdnEmrjGhfPekm+kXzEvdHp5z
sBshnxkr7DkUQS6Xg38SoCU96O87nYasN2RV0mbOPLM+XnXQ71MtYBb8eB6e
9NsLEQIYihCDCJc1PSqfTpwyISH4P7/lZeYkb5te1YujC2ZW09pb1kd0pwv8
/jWrfEt7da7VqgW1vBumjpKl4lRIT88tlanPUYvlTL4InZQDmab0mv6D8pCR
9txoggUQge/A7wXUOEf2TyHdsxpNrtTg01f6OEV3NCu1MZi+YxUxeTTpcKWf
vTdqjXW3Sv2Kq439JPG80B9Ejb29AMHsIgZqqE9Yrcl+MlDkh4AYckMVu6iC
ZTsoc03ATzuJi3zavmsHD459pBiglgFJicFWOY/KvS2fq2Jkw62JFG4nWBOD
g0ca7vaQ88sWkhc+i94/eqjOETwzmZ5wA0fLV1d3DT949tPPL5aNO2g26IaL
zrvJVTNm02E1DeXpqWBw44sG7i2f4mVKwhnGZVWQKqco42XfrhlW9wWdk71I
A+aOQIVuKmbS8ltnJ9gqqooEn1NhxeIsmzmbfb6fsbcpFfMW0llLH+HcLP3I
GzfWv4Rw0WfeSV+JRlmT8813od/1HN39uXZy9uKj4Ydl/L4R1kqUrzVts2Gs
18Qd/rsZ9MvjJ8FhrZjfzFSMBqbQ2NWxKtIhWiojmNvCWyX8PeaxORNZL7O8
te9GraJ6y51KUzpp4+0SHtzpKmgUC7TnoBpJRUtERkh1j7ay0fu7Ax72hSJ/
+bM579isd0BElT4c/iKPD00Et2AshmSoMrOqwHiVy+w8J5sW2EYADEDf7Nfx
oa5kXGYGNTKKCdeoKW9BZ/OBrFPgab6IsNXTDy+p5DnjHJbD2Gs5Ad+LsR4K
9KXwXK6fhHDV9vgCDlXd+DyAk0cnwaUqiT2gBT2JFnLzlnAlq7PnuU3RKUkY
RaO7Nf4kCq4DnT0Mf3kdPLwHnfbt9RFb7vVwUZ9z8EKmMK0lrpV4QNy8d3gK
2fLLvTfwOD2X0bUiC7CIxArks8+vb3+ypafsAoz1fvRKduiAczz6+ENBeIGh
vZMmujwq5fiy4yPnBkliWAkFwKx7Bdts86S4xKJvnpfYTW3XGhIuESxuUI1+
rvIlJ/i09I5qjN6FHMBiz6VSDT4tvZGulmpIdS9KOPv4uyQPsv/xvfCyz9hI
jBBRtvOU1Ai1Si9vAz3xLnUv+SmTLLTOR4vXDbbQFIKNTUd00LErCcJWOS/h
Xmmv5rGjowo+rAe0qUkc2nhoXnt5sa2aBZCMmjHzoikiOC34ntEqgSpkHjVf
jgUDbsxbJzNXJxTk/Ty2M3Hf761yqC15OsR6GfHvJ4H78CDyZDO5ATDdC5sT
iauGF/sEKXWpGd09UDQCuArGPxuAX91yJxc/1HZFHDe173L2bFNoGPBXtDtY
861GsRogPG2QrdeDavlXNwMFx3Ae9FHISXb8AwUdNmAhuB0J7cUsQlePkUfo
9UCYJSl9S3muNjm1AB0BLP3b7/DmlphsrADrUJ/zRVtkWRME0fz0NzEbLchp
c7w/Vxj5WSgKGnwl1pDQhQCa0Rcyafbcix6wQZ/PmeRytvy0VJ+6yDfFieW4
LlzsI1u34uN04I1aQN5wl16fSeESUexDYkWUhXsSPFTt+boS2vQjjHRKIMJi
+mJWRO0fbGDOEhBXfAzEPl1kfyd2ZkN12/iQfZtkpYX076xEHbdfKlogdAMT
qPdbHjqfrcrd/T/0z8rmfq9lxmR0WzZvdBRDS40CmILzrcAn8+nl2AYcNbCW
JwVeIwSvFxasum/C2/Q98bS+ZBeFgXLTyOhKBn4FFKid7zy/0nzFUiV06jO7
OtUO75yH4o0bqQ1/tpPxv3AuAAEquoctrmptfxGHKYh5vaOhwPUlSQxo/7gf
Y471cRNWr2Iseum+YBMUun3fuK3toMcRF7wgp4RO/mLLHMXITfFoI0yPll25
qFDmZ/Qi9D3C2OIgTs3qzFDb+lthfEL+hvUNXca2oNcqY3xyZfvitmhHCiHb
Xmk5HcfBbvkTLdotjIxtpRBclG28+E2sJziIQu92g0UwqldFBpnG09lphTv4
51vyn0VLQOxMeK9yGzjaHn0SPt2lYH76gETTdvVJ0tEDrQS9Ld/0e041XRhC
f53XVeJSuWZ3TFk2uat2whrrp/XGzxUr+qw+ylKoTGiYB6qmtYZRfTbyigam
DKt5vLYTmb4n3XQsTzzlhpOKQQiym0Rb9Ge8bnV+N4eG0yO+K9ZuxmHxt7Ft
UhbOVj867pxsIzoGrYqAjhBOMYr77fVxIqt1QNyyzpVXKqBLseI+UfbM0Ba1
nxUrWnQLTSFPGtSt2l7ozZv4yTp1QXeBJTDv5gp5dzbjZAantAtEbCUzG8cq
guDH14h5iNUvZqVJ2r1BkCw/dXg2kV05jupETAQa5WtRnqop0EyQuw/ChJsU
xEIwZmrUrDk25K/bbfjzX+moRIlD2/6fVO8IQ1f7ATjsjaR8cmB+ALLxuJk5
I21UCW3ZJnInwjJ/GemztMfXUez+2314vTs6gZw8fIY1GhvLVMhB+9yL5wX2
ys69jhk21CzwMllfP95nyWXF9TbSj3ur5OikANtRP9j7hSnoO4mctaa2FWMm
hJnxjPHJ2sfeklCsKR8RyZ6kdSpjNd3oop04d5EzxlnOGDBEZzK1kDtjyOC9
nPiHW3KY0l8mS7FijtbOBZHi/BhYpWR2sJ89qpeag6Qfvm/1EEuYTVVGLLDB
1AYd/BDgwWzELvlSnAHDiyg4655EeueST8q0a3crFMKhFYn0WITQm8ofyNYG
xA3GFe3pRsSauGDDXqtQoGhd7Rloj5zxbNRqyUTC9e0JzER5ctie6FosGZjM
mwLIpeFKC3fuuH9p6bzVEgbjMdOLvIDCl0JbQnd0O9u/1DePvtJYwvSRFkPB
ZyBGIBaBUuWYYWINO4wUfSNZcNWoOU9LKNkQObPUMSeNwkkg6U421JxgRA77
jsAi880vf6S0O2RDl6Kxnx8drZOhQyjEAeqVsHwiA/1dw96xvAVt8rxro/rX
mWTIkIUBTf5el0klWrPw5pQj4a1iR7pVjRWg9/MryfQDDo2R8DfA0od5F4Vn
WbVh9vAA7IBYjKrhXcFIwAsJm1USVKfywDSQ5O1F9u+ZyVzWduy/4S2uLUa+
JXILvT6U5bSmi/J16fv0T4Qc55SD4agjtL08WGZMkgR+TyhPVnkPtpFwSQ1n
wrd/aj5aoNK5IDA6PNZANPdPKQk8ui+IcFYfJi9tWjEnHYASK/Ae+NQ/4gSz
mohflg7jfYVmRYQrS+E9xHwc9/tnz4L3+PxmAzjv49q4ox7PKyMKBVG56eEq
xNWrYDvpi4pUuJV2z9RWIn0iRzv+fTKzK8lGoVZovGY3NjYUxq8zwlKjtjCi
RBw2JZP6Czl3n0EkP9qwIqQsomBAKqn45VQQQsFpF2tA83umQuB+vxcTeqdW
XQ0h5ZftGtrcj/Us1Mzw2pd26TDAUDr6euW1w8NvjkOqwTh6EIYIZ9R+GIu/
+NFGHnHO8vuYCIINYqWv7yzG5Em4L6Z3lKe3gEAR0+0yNte+15w3yxHiiIwI
7FwGiRvt3cAJ88CEpT16WVMSPfd56mOy97B/rFCdlwTi2vXjTP3e/TSdk4Fs
xyuFDGsSPySkkYQHqOeGfALuAGlBdEl1ufT6I0cUW4dQvUOk55hhzUQAAzss
AnpZnfmt2rQTKYC7OZWUB7qhV653eK8neB2B9Jm3eSo5bA4HB2k4fwlab4QC
jWtJ4ASokNx/jITy5eUNqb9UsARHoLNIKS/mGJwoMqk0kUzSlUSzapdik3ED
zNWS0LLeUZueYYiDMg7cJYk9agRn6QJ5HWFtnMI8QvyRuQOGykWLJzcFO13o
tsr7a3GEEWxMunzF7uUQzCgCOk7v1lwqRu84NnCCrmvMwUPeUn50YsqzWUee
ak0yyhb8M0NGzmrgQeRwxHWg8k1Af3W0HrdW1O+tXJSfB1vFQFscnUMWISaV
mndOUl4hM44TDcoGIJA4he/qXh2dYA+oUTwDfaMuJI6RK8mRRkPOiEjDx44i
C560/yPl41bVRv+eGf5nirJ8zBmn67kze5fOl3bO7Go9CdM+JcR8uYCdZKlu
rTyP/H/lvfMqKA2LPxR1oZCzH0tIdjSP0McHFbMAPTLWVdEmqaxFFxcVRufv
a3BOy42YT9O3t5AxER/OqZX43TuUMcZJNuvvGkn/obDavRQwnlGllkDAAUSA
nGYx2+sduRDxhlU1ZJvzRVrRpu+Xsla4/ONzszCyRmNvWphdJjDrlPRHxIB5
pmkVFgKQIfN6qUQmV80j+T53c6MfrBNOFSqHaTuh4DAQ3k4US4lB7deX4+3H
s1mnNxNL0xiSs0Tn+P71ETmyPr6eEFnlLb7NvrEkuZBRM5iOKfk+2+fWZNHE
14biUyos5rXQoQAUf3z32xIrma9cQ+J11Vw/7SCE3vKUgAPzH/9qwPpZVe7Z
BY5ttuBPbkEsH7cCLfuBPfmfRz/8zqzDjkyPdPx6c3HW4quFZTROMXrjTA4R
jM3a+BwOFQfBZq8a3Wpg24pdHWCmECQfVUaJ/tG0nRzCil7Bl3LGxtQ7yqA/
oGoXPfz/L+fFWQtFVfM4hmkD7OfXLHVmSeDlBQlqRNf6c/McZk+0WyGrsRoi
slyOpo6wpewY1Wuen8HbGNN9KKQNOFfVMChvlLt1hLJZ5aYVJCPAh/MbgKFy
m2k/97I1KNG3pt4q7BJUC3lpkdiyrHjtvLkD4UOFLQ9Y5i2bDKZTIjTE68hQ
Ay48GcFUNkAsle7QHxJMwHpF2H0KoeABiPvJcCejcY194NNNK3youdYjAp2w
kIsbqgDciK+v+gzBcWg4pRVn6KNiz79kc0yK82LZ5UYXlJmEJm3xG5kdgHGk
prLSovN8L3tmF8ToWJl4Qlj1vVmIeHcbSMgkTJjw9h2tlmirP07lsra90HJS
jkD85wfI23hjU+C9IF7LvzLgXTxPRkCxI3d2t5dl8n9pYMnH7AFNAPM+Tbfn
dQELehbrIslvfGyed67/Ft79CNPqsomITvIb/RfXZtYg/DV3yaEXGVpGwccc
QmvHstrADHkQIuZfah471e32K5C1oW96dC4wXcwJvIUhvauYBUerx4w8oHYq
ojUCPMd2ghIm0gNjj6ukWlV1qC873rAn/90vxKRj8lOPUdAe0YiKdbKlwEYo
TZiEE+ICT/x4GjQrMHs58/o405/n3lRdsOcMLWnj3QbbgvSZo93A5Vyv+VD3
7agg38o9f4U7BREAtqd5++e+q22i6xXtNaajeYMUyk6gsAswJoZMLjr1e8/o
P75oXqA3X9VuMfRmU1olP94JewSAZ91dmpBLEv/uIsM98nsF+0yMqUTOnMMh
Q1B8x40CjOfzV5c4fhdFS9mbRNCVoKGm4Q9I5i8B+o8QJZzDM0yxuNx4yk2z
+2k5KYOu4MXyWggdLfmC0GdK3Z7d0FImzLYJDa+kqgtEIU3O4hnCefMlUGDd
KODisKswvPmpLXS4x3rc2QdHXNPYKI0upvkyQhyhPb3g9eLSaA0KNHwtp85p
YmBEjQEVEWAZ2YKlD+1pq8XDqt3F4H6NI/fcXsGIipSeMNebygPnPH6PeQJ0
6BQuzhi0but8jyHSMJE82dMXg6saZ0EO1Hs/n8HANZJlt+xz7Uwjn8CqRDua
jZS/o1XgKe5lvoxcITOfCP0fwK90xgtNxLJ/oIYaB2iK46VID/ysckc3QalR
VKeqhrWBw8Ga5o6rxu2HUSU/n4iEVOCpO4ErMMJWTfoIm9FxUBWL6nAXjrQl
vGtfd2INHcn8NFnbRZVrSsJUEntjsWBLFROzUnW5l0B9hKNHBauSCa1GHyKS
VB9pSml8KA2J0KbZ+Zd8XvI9mIs3ljk/FFNtdQWaJfs0nr7BshHOmTfKSnlX
6RdbLpRuJzJE8D/VIYlczzIloAdzGEqhG2HKIPOqUobLOJ80o5oHYBuXjLcS
R3BDXumvYb3acSpWxsKdRpd2iJq9345clrfh8Y1eV/WcUiHZJkIyNefcFg26
pEHCLfbS/HUg4LRXi6txMBzAzaH1kHZ0eBERBnyekOVhwQ5IPw+uHV9hxjYs
Oa7no48aYIOHuP7IfcKweFeVBlT/3/nww4cHMustTllRg8SkfPO1YFnrQwdK
sjIK2nmPcl/rlWnA24K5925AP7AmvuP6pvtv3WXtr1fz1KNX5yFMmLffaWpH
AGW6TZzaSes37h2+kvkGPOiOcxVO6dEmfHzqB3jAGkIlR1UZ5j5GSQ3FpHJq
i6t2DSOcEYim/6eSjAZ7Sxs4mUhGq/WmfjjM2V/rI0BICREgLAPs8vI+ZPh9
UxNyNlnDqyJ66lPQGm5OepmHd2O7IK5An5bH+7a0EmOV4urVZIt/cdwVfTWM
BTenx58td5R7O2OEA8Xw+jdDxUzXaBbICqPpNxxlJgKwPwZXzfm0OMK4ojAt
i6B/7ulua/8bDJ3XdlkO/t9p5fkW5Q1RAGcTPXP1hbhaxoFxYMWpUQ5ToKuf
bQ/7Rv/bYBhEtKVGq+d5RK3FQJHd/sJW+8I0U8+ZvWrokuBYwRUxVMLi9stW
qie/g/q9cViIHE0K9HZ5Ha+RppVNSDDUjmBFtFV/qCyw7U89FteBdQRHsrPE
R+9tofN8ZsFaxB8pG20iXCX/YCqhXnEeX6hJrx8EgJtVA2x5ctAl/KhxTp35
B1yOzKiDK53zbnUpIwiuW0wLK8/M7u6ynqTZLqxPQHHdb1JUPNUZ37u2ELaT
a2M4bg5VOG+Z3OcoAliVv+Y26VDWV2bWfc1x5UYtqqwL/YOxlo6wA03mTtlo
G74lvJtmxeH09UAk9VqEmR8BR5A1SsXyLgOt0KcmZ5ychjOK9rsvZm8bNj28
uJBgMeXxeRE41Zvof4nMFb9vy9uvIZ49nntdym6HzDMmHpkbsmru37IYQKRj
gNcU0FaSbsR9ECNQzqt7TZDcJXDlyqTJ47U2EllYmBKpeEu8aEWJ0q9GM6cX
1Ew4FE9mlAusN8x83PmCU9zAkguQ3DPHRhDjBuTYa8CXo4olkOgXq8m7mp0y
VgCOvMBwllpaWTbChy7OHmv1Hysw7horyhTdqcyN6RjO2HnQRb7B/YUgzVv6
zVE91tAUS/VdPJz/PSal57uNjwAoXlwPdDj255oX02yK2qR36rY1/O3Gm4YI
J8kr0F32ArviWXhjur6yCvQ9iBtvy8qmGTqrr+f5tsOIG1GuZpj3s++Fmfq+
Q/3Xico5L5rm1eQuRbxVrK2lQcC7gvppoM5EQC6iFA/pw1/3mAtK/ZyfB0lw
Yyykjpaf2HOaG6Z5AsjyWTFrG5eHM4cPjAUcHbMbo2VlLU9ezdfuKvR/kkYW
1NOD6vrHqmolEI1+YSG1rL7/y8eVq9sW617JuchMr2cpc9vNaPm3lz2lxds7
w83P9xTQr3+VdgcPXjLJlxP1lWH1NNTMu3E4bvzLGWdhqdPvv6DHYpHbhjz2
HFwBS+Z52bhD2s0rVFElPs4MCM7Z/rOAGdu9NJJO2kDgGnl7zLGYtcM8faw+
I9E8r60w3YEfIFug41BfmCdO8GygMsVAAu3veoyc8VkTzfCZSlA+qHa9IvkQ
EQAjvmRIhay5R1OWcf0bqeytkIfqWTOIqAo/pHuPAVXDDSkwHVubwSFJarQK
eiIoWzayVHqZG3c8VfJsk7BZVwFLmLb+wmW+V2QDt2eqzSjJlpAngwcdQusB
pN7lYwy7G2WYa49680c/52lZuNbmbS2dzJ/hxRJ9+blACnZcnHDfetwL+ZqN
UKv8K9JQFZCZUtsPNaZxRtR5yth2c0pPF4dzeOXrAFfA3to3wx7Mqf+Zo7Ot
HIyn17k762rU0rgH/eximWjT37Y3ypd6gfGmpDg4wIuMfXC2+UzZC0zoB1Al
9wR4+aOqpRBEILeVqQcugCj3M1/1PwxZcKqAamVv4k00RZ2qMjJE8pM8qq4v
FYXC93kyB8b7g+GeIF9seGhUoWziJKJWuipY4X3f/rMjB1B+y//719W+/Wv+
prREpCjrYpJPVOYmNTf04XO6/EUTvaHpLTacUDbwk21yc7jKZtp3r7nVR8fh
UORiq/aFaS5qLPFYxqTL2VACvmZPXXgjR4imBDuwCkZqMSRoPABUjKBzO9zt
EFj4SA5bZa4aGLJuWN61VDzbwx2KtDD3pl0xgzFeV1oRJ9rP7BS5jGCnInE3
B1aLHvIXup8g7FuIpWptjVGAc53iTpBlIrZTkEdlvoySRcM0fDZGfMuwvDAZ
1pwVCam1EafocwVBmcSnNOET7YmK8Zg9WI2pMw/+xLrmirQUOyHroP8+Ziyx
Dj+FwYC4q4D5M8O6oXvx9YIJOrJwSiyxCmPUCVMVUExTpFFakOYqqhbuDT3i
NVqNXamdNYMAW5DlB75Aj8vFtqxTSlqnvGsCjPDqhODdelbV9vilSGLt5AT9
2wWp0A9p2T4i5tSxbJ0roCV1DjldTd0xU1NHhAS3mgyjponoHcl7zA96LvO0
CsFnL7fKngN3B81MAuwvkeISWpD88LsmK34E1i+NXomKIHuorOk3Y0Vr6Nf8
bWHOBNOPRzP+7CyWFQBe3xJ4FHznWtfWiHUnaKhUNAFo9kOzEUl5Y52aboDv
pLqIN3jYI+yd1emswfhub4/I2qrDFNJ5X1293yn9L7kRHdjbcy2UAtoYyOki
788Dge9XsNiwbAOLawq3dcwpz2OQxOK+ZRfMw1emBP/mqP7P9NBQbgtBs308
6IrUzNsNm9rlSJ5mYO/IGhJiIAWJ4HRT+bluW4tPEZqy5tX25MWy0ys5mmEn
S5lgamY2+/ro7WbS/wPA21OOTbSzCbN0bE/VyAeMky3bDLPc7t6d0dIwEfGb
A/rFSAeRD8j54WdFVY6K1WH359YSUtywtNtsOk+Uhlv5N3bwGvI80jLMUpyC
ZoGUkmXgGweaNFfvogwMjlaufGTYUydcLPG7T8YeoHputS4WkWPtKClGq++4
4W6SLpRhg4AqXV8Cgxd59aL0Bi/oq6kwe9Nda4wz+p3m3GdChtpAyTzIm8KC
4vCWPNOS4VDHEIx7t/s8d92GC1JaJyU4x2QsppXz44dKCrpLZJxsOkYamDS4
2xWReKElmQJzXx/WiV8aXRjJtCgAS37Hd4AASqYUv6DIOL6UlEx7MPYDxcbu
KcV6a1TTXNDhrVf3GXkyPUHk7ofYxyPL42l+7hisNX4Su/qAVYSN5htaxmH3
qpK63sF/Oc/Uk75Pm9bMbEINNCOoq8qmzWHe+6iucCiYTJASbmfLEhHxSb1c
jMxYAd+1nWjRd5O3sBO4iic2sCfHsWkIhYCzHBPkQ/4kKdyVKaa2WR0oAshI
LHahpYmQ/7NftnWmjufhdXNliF9qewAGfX03+C5a9opSYs+oq/NSrjBF8fyJ
N2awAksk8ckCZJofD/d0nHs3ipTrHJT9gqUiHKPdOIxcxS7Tt2aed8qmlfK4
MgKxCLkIQK/F8W3hxyNn4AVQBWIDTL7CQSa3yAesutJucfJPZpCv8hTRVUJd
cluqR0l3qCR+OsfKU8zxA3QS/Bl4fCbUAYR1SfhHbBi7vXdqvLKt8iD8m71U
Pg/sOHXhjnEnroFFQwMlMRjUes4u46tufM1Qyx0MgX3SPBi0UHhZ8CXFUXYc
221CjoBFacw7n4hw4ZPSpvqzKtALqJN2+XGR+0beSM4niloTjimrg+sWnXA3
rcgCp8D7SR4bWkOCeCFwXlGyEigbtF6kCMMq4MImUsHXNmhXBAXQL+aaVpTe
Te7p9DJ5xGbZ1TfYC0sEWmX0VkDKdJmvZtgXu4kwIaBwG5rcv73HZ5AyI9ZR
N0bKf3jG5E0bAlHoh5pwb+dBmYZO67tmWoZndI4L9NIz9CYIxH3sOXaavN0m
xVu01d/F+j6zWWBtbWx+HWmfuzQkyG6APaHJ8+xdXbtuSj0r60kYigu8HnAn
Mr1xesjiRCLxA8EquJnrryj5fZ8mYo04hPjj/I0ppqHH+RFXCSMfqXAL/yGT
qzn6S01kSsi+rqbvrz0uxfsDDP3N3Ylfwrp0s84XYW/Z18WzNBKdar7TnpXW
yOfOZhmf/oizXxfxdznqnNyITHVB7jcdrM08PDpYAZgI+Qk8kKirQ4A4Tpcq
HhmMGYRd4qyTtCXKw/aNQ2CI2Rwd2j5/Ia1BalVrMUOIereCESmtsDSRrmYW
g3zQ10FZRG3kv3WhwMtrarJTmXtlodX6NcohKiDbd7nVPghQNLKDQjZf0WWM
BRQkyDwwlonb53CcopKxdOv74rzmHN9nuP2kZb6ShQVS6Oy1qenPUq7tTd+K
Akfih/fVJMtkTDsdcWVUKFK+Uub3Pv8l0fxLlfJjLf1cSA9SA8lAZUbdxlc3
XX+AMlAh8IzNNavbnWzxxgLxH3IgtI4kw1Wv6j53JtzW7LYBygyJd76o3wBi
8NCSs7f1/Si7WeMKgKtDXX3DrC6nO4YRfQFVFVRxXrEaguwWSXJhAld0f6SF
LHdnr/kW61fNLWX4IUgDxEgpzznuqznpK7AO5BRMXtLaq0s9OVtqAOyUAsjH
E/N1YjzeACEC/VMbOBr5ej7D0dE9QBHwIOqze2NFrJ/Xkr9QbX8shplpvurZ
wN+i6dAH9jAzJcc/XL2gn/oP0QvnIYtOpoEQh6bzT4+f4E+0FmPcly5OSKbx
C28AeIzr1kppQ9wb2VCWqOPnQmYH63PCFc6m/3Ek4o57j/UgDJiQ7Nd4eNeM
+vUrkmy92Bar4XFj9RnmbtL99lFatAN0HS9XbZDFyftCXaKmcm29xSCPKARo
yEGW7FGhU4mW4zF5xANurEegac5a3ttL6Xz0SV/hVqmtBihElr8eZKDUAXOt
oU03U7ZuAs4rO8YS4z+cm4picyovkYTUXDOEL+NqjFyrmuGgtiehJpfLXI52
CmwfdORaJHKKYxdbYaWIaOKN9V/8NpGzR+G7dsY/xHlrMJjsVyCPzMFdAFDj
hwKlQ2DaWJTGrAW2xiZC4Cmvo/YiQEKqzgtWFu3718piiO+ttE8WugIWzzz0
14P4dSpoZrpGhBE+0kJcLky4504LYCKsmESk04ulMszJNfrnalhCb5MvvJmK
P2kfe6QGViguMUtEsuRdbI0f7YiRXZ6/4gOicLuMQcmolJKoWXznoTrEMGGz
6pI2uJI/X9LGBKVAt0l138+1SvYPGC7Ag1/Z1uDe/eawNzz8tu1NL/3H3t+/
tgZRo72cUffbzzqjSFSa8GWz0zupkMv77gZLvHzB4Z5i24xtJ5CDUpYGiSbZ
/706wWtnoOJE9qTBDgC739xwrgcikwQ+tjc59rzjTrYKu7ngnPdeQWtsgnXJ
bKQ1DhPr48w72nIut8sWgNWiTFrNtc3hk9SIGRjJzvLpx+eufcVkas4n7VKk
xKKKOQTzrzjB6wiJj3MPud6OrZ2maWkuUkk3jeEoGdkO5298AbANp5KIxFPb
Lu6CLF/3QHygDCd5VWzX/7Ec0NI0UOvSV+SeyCa8rv4q+CB3JpYm1iFU9wAb
vao5PmiyTkGb425hzVi96pPgdnHA+7wDfuiD7myVdST/j+1+cDnS3MqX7q71
yvEJClXfuhZNKL04NmCODd7UCM4zhDz/ZnZbDc+hEehpco15v/tTwnHYAcaM
PxfCkS0i8IsEM0g4bSpGc8Xznkiu+2XEdviziaFW3mOf1BDJS+EzCc5fkoCn
+f/FUh2QJFpoowPrW1V0RCveB6vD84L2tLc2PIQcSxvyFGtEY0v0UENGDP0P
2yEVK5fLNqdMPOSPW/sfh1zjJBEcWvmjgYBxqL6oO/dkw33Ix/TOrBlnJ6xD
KLQBgOWotZyAz33+L7Zi1gAePIlOmexdUvRsKZG30MyWbn96FlhKc4P73cG4
cy2+9q/zCOZb+UhWkubUSCNaQlY2PP78Ofi1YISDAT0igPh/dyqwV3puVE0e
CprGED1xHPSfFeXjYe/VlpLUTPM16y5jVJQkG8YDTUxY2X1mo194aFNiBY7V
24hLVmWGTCaRILyNAon6jLiq+qBZp8hYlJDz2OFlKx07ysZc2OZsWsCiXJQF
GWzCVPBavliggslGTtswXaZK/WUZDnvN00sBUZt9eWqz2n58G7E8023uLakb
YlFiY8XR702exWetwJjYEAybuWNPlO6q/NfROWO7yq3YYrpoclJ5t9hYhZcJ
pSkqCU9klZ1wYR8ptDLidUMR8Cpj7av+gMnCkrf3mOxfRiBSRizm2/+eCJP0
5Zee3TcoF+iwEMqdM47A4DlR3UGRgy4hfXaZsUM3p93AWAkmyxnYQkkClUMv
7R7/pDWSma5iO96HmLGb/IoNyp+a3gdsitYxC3g5w5GS+LiNojxr6KHaRxDS
5trPB2vGYQ23gwjsKqKps8latQlZVD3bOL00IDIkIcaQMSP38S0rWhYaCkDF
pk5+aoso5V+n2punYU8bnh7DR3GSGozVLMyEFkQgffUVyMUcJkIrIBYWz4yJ
QEm8Q6NDTE3xJeGMA1GEZOTFcWUAygP9MMtoen74oZr8u9VdxUsLXtqqvxfV
sj4qY4ymWDyQkotsaOurMFHfvIQwPdJvS/fCa2gxOnA9nczXToDNxqzKAYCe
VRWF50nri5LWv6v79bn3JqyAnx+DkuET9ia7kGcl25WoylMerPZuzvdqO3fe
ilbOBmvlbjqT4P5TVL8EVvuuf7/3N7oFNVJV00Z0sa2XRpS55dQ0TITXALrn
M5wBxB9BlWrH1zQinTBeZ3TGO4VSuUzpJdEsLJ4wtQu6tsBuhw2nXqxsCegy
By5GlohkVk6JtOoOD48hRM5yUhPbxEY8U6z89zMDO44L9E5RhOTVZzL2AWdi
/Wn5+h+B/qzMm3qH1DEewnewSSAQMkGbhN9wNZ1VhaogT4IM48e7Djop9vgA
LUS5nDzXcdi2qYSuIqJE0lcqMH31zwjnmr8DBpcHr+IBKcaRa+BV8fhpqkNu
LP/1/TayQQj+a9z2e2s7hGIhqBm/JdHmpplbHFj0CSEwR+TKb5zl7k8Q283I
62ZSVR6+eUKbv6NDH6S1yLFwhYnzp0XRHAoa2CgbjF06HzXyKXDg84CV+lOD
/0dg/lWuKzfui386p+X9PZ5hPovxNAzwXaoeW5joOnLwktyU3DODkS9XPeBu
klFVovorHfiNnF678AdEnI0tUdeIqIjk7jYj41a0JVoUFaQ1W3L6kWEF0HOB
BIlBNFTBtDmbFfbewA0n1wCtnn+4NQfU2tUH1EfKPlD4vxQ2knUr/ECjf6sK
jQFSjPkliFUR5liP6Br8duV0Rifa2n1degw/sp9Zs0oWSSLUXyv1eCYu4El1
yH9LV2JTSe/YKxLVLQzMux3E3YHyixN71a8ds8TqhEWMQNeM5xbqq+9hTT7e
T0nDg1YOmQYwaRFk7rL0SE1pd0WJCO2Tl6smdb8LOkCuebT6f8wI+lU1VohU
BY1V1YykS4fdlTsKl6mrh1YpblJA3N+6WwDdSm3hM9WoLvMdlsNnJxrcgUDe
JEJFYZ4lchdLeUPncBv0qlPgdYK9mMy8wZldmkqcZtStpgcaxlVEh2A/lDbV
LpoewtSDlFq0/qSpCnIsz/l1gLNH5y0e9FzmllD8kff3BpCXDh+X4I9NOzj2
l2spfVaL1sNoG7NcwpAuLapgf1DZU1wQYIfAjZ0cf5cmmJS/vU7xnRhhvtqR
tGmayN63iN1RD078FumbvIyZn1hqypOWXlLg7e7PXoBU+WHdRSmaiH6KK7Y4
/f00iWiDImcHqmvJbDSfWGHCoh12P9MraGjDsiYTFO6zpDYO5GA+yTEJpkbv
jCbrUNIvT6kft+FYz83gsVkpsdergNIijzwkJm5IBBROYRB0jrLdEcM1Mxtm
sLrWx5a7RdczRtDdhEbDdBrLaFmrVLZKRzk8jFsD8waqm5g+47U93/9e0xgR
hUXIibPY//CKimJ2DrwBcdSW946C7DKPtDTaxfJt53RfxQHxfZ6ju5hxeDmX
g5GCKDFgzO0QK0DPluWuqAkluaMxrkTfg+lop8m8uBwWd+GsDQffJPNnvblC
gSWyvV+PtC6Ddx1q+/7Rm1acblP+8sOmue5XysEEY1TMSPMKBX4jMqzPO+Sv
cQRBdNcuy6txR1Sbl5A8ATF6Kdc2aLbE1yR43XTiQ7rI7zJkvHnWBCJXJE7j
x/jScsk6YGunWkIEHbNJK0pROOj/T6So71EubsAcizF/smiIXdMk+JccSspM
Dbnfj+FIoZyED/s093lsOvUt9ofKxCuCB7RF+jzbNQBiR3p+O/hHv9v4zI7P
TZVJb/4iCSigVwwqqRyEDKgs3EEkSxYUieqzlH5y0KXMaVLYJVgRvxXwoNY2
59cBUMTrl9UUIjNs6GnB3QB31yJSUIjCyLPBkrkMwiEMvnM6L4HNpyud5szB
GmcKS1saRydQ8je4//DUQqptyg5LN8hk2rv/dJcAtslI6olUbY4Srvgc7Dpu
GATAiv6Gbeio4D9TdgqA4H2+fWNXX7RChG5xbIDQzbkNfWGby6pFZF/NJtiV
NenDJ4GgW5nt24Z7BMcimYXTAxOz5LJ25cO8F9J9ztY/DrclplaJC9SKEKEF
XK0oEq0jvt2BqpYuDju7rewcw4LJzO0Jz0NTR2NuuwybxHa2Kbm0n6RBgQYE
qSEqo50xP3FvB8pN52C/AdNAeuONMBdD+18xEiLJsNT7Wn97/rWuYhwImB46
NeqLyl07z8Jf6A8SWOHn341OZeaqOifZgsaT1uVo6HlsOr44xQDT48yMfmBY
hiVcrIx4mFh1LX+j9gHXnB9l9PtkWwa4L2A7q4RTuB4I0UsC44p33opG5qrz
jnfhDs4w3Rz4qV7qTq8wwbEQk5FhjaUWMorScxP36J/NJqAYuOADZs9dehcU
oQhtpiYYU0PsD4vY8hW9Mio6RbUB/ybCRNENiqqySxOZjlx3PCmSyilIUS9q
BrXdbRkv204V1tX9RDQcYEliUDnz7sdvzUE/1X2wYF9Hm9mL1FZyHUWUQxWO
qeEg5poLUgvyrpSotW4JMONPA7ydkAqmuXKSMwmQR2vkFwTgcWJ1sDvWlViB
TRZzmaRvftFidINc61qgol5BFpRlKP3kW9HevG8TnGOzat4tSAHJt8F0i+W1
mLEqKVGfb/Xhhs8GZNGgxZi4I8hrSWrRr2lhxuVnsT62HsYS2S2+d2YxHARs
krNFGOg3X1Ol+QB8GVXbsfrNvDGW49r4Atgq1kYcx4nUNtazMj2eAtLylw0Q
FLFhDUOGx71XB0B0O4/bMBOUeIJLY7iAN2jqeCmRmzKbU4AXLu3HRvESmWw2
XewgXwtGSgvMsXlc6PR5SUDrPH/kQg8EuyzfRSfNQ85h4iKYeOMAUdK5l5i2
CO4BXY9jmeuofJ4ez40xZTxoCLEyWM6Ca87ZvDgltK6+cvP7g38Y7I+GzVJj
WQoG10wkQPxdf3rb9uwHlMftwtDXPyqQW9eS/hgqlkSojBxta+9FfnrN/jO3
0csdHBG/qsoPAgT8sUx63knsiDoRY0NWrbP2bsCPUGTegV1gF3FRoDCOrqsP
deU01yMcqjZFm4LMMNB/k4iAtp/A7IhmKnLMipijuAvzr1IyiFG179i3ttAR
UC7juLKQom6Xc3pfBkJ3qRTa+5fyFCoSFX41TiCvGep5UNf0xIk9f3uKEomt
EJ0uYjCVPUJuMRZwMFoxMfu3WI7tu2t88Ee7WKOVZcAZ0WoKGmiiWr3MY/XH
5FZx8af+kzhEhHq35gg4Py+OICJr6UKIf8QqHx3NyfKsRjr9jMsHo16QY6+B
loMsP+vrkgGGAFbDgSSBOvbEo8+xd3kjDj4cBuqNzqmfdJpQory/DkYFv9s3
6YtWwvuann9PT5bgM8XxLcWVwCWMU8zcng2QMsITLyM1dBz9Hp7ZLPl4PBUI
CGq6n0aBBL36uAdJgGIZQfP8RkxAQbhoZ2qksnj8HUnWG/2IWP7RZ93BkNfA
IUcvg+m8AXjjXv0eg8ZeTNn+98hcdU31WuJsU+oJCBkDwO6wvNK18Gepr89w
PHmYw05hI37VpyC4rgDIPkl2j4aHZ8vjAPBIGE8dW64anvOk6icrc4hgLN/8
LzQeHM0yKyOQmjBGFE0EwfhZmdAUhvsxjuRjAa/YQHYdhWlvkvV83wpeLLNC
p/KhpFRE/AXANyydlikSsyzizJRoGycOkq4DYWSDm4q7mZFM0yF3PJkJRAWR
YSfqpPm2tGSzGzVTBt4C/67z46F6SLv7MnmBERiDeqneqqFvVBaZVw+DxlP6
D6LFULNiNJtNuv3+8855yKNJAJdtLtX+/COy8qIBUHOJyVPkplUSSs7LKskO
LHK4JarLRiIU/wUEiJrXgBuZF5Zd691QHbKtLdcp6MQIZNfGN3GqaZar+eBT
Ma+mgGHS6EimgyuC3ZKKGP8t61hgoT414YDDj+KPawzljRz+oX4fcfjY+SxN
QxbFZL5/rK4qf9XPN4HWdX91L08Uhiy7PRoWLj9X4UHQW9jzl/JNaevq7BMq
e2OfgJb3cJfox8YjokHekpcKQ5DX8wgHqpvrGBNO4dEhKl61ag4ushd0jwou
FEiP7A/aipA4k3gNKJC7SNruTuGLLcoIo/2z8iPO/eBMbRsR+16pG0j/pQdE
u3kg5vKgipxtGfCNnZjTMfrBOuPBK/rzT0u8mYAEYtnT7P3qwmhHTW8kmHkG
Vu5bD3I3pnM4dO4K8xvXWjlp0tP2YtvHA/xH/8c43q0U2060uYH2OV7FxADe
4T4TAi3eijtbi2Tesjn3K418cCxMzOAHkT7sbXOfRUoh+dNxAp7wjVyJ7J10
b5uc5XG4qUxui4LnvsnKnZ45i6FctLt4D2+W2yIkcu40dnvBX1nGPLiECodP
KI0+boOMaDE2AslJ10rBxiqivhoZOaPL+Dk/DBPDkDx80yqN/JkviaPlZMDv
pr3abhb1DiBJKNYuQU52DYtIZhyQRioFTEpCt4WR4bdMfq3MrYTJxsgoy72i
cqaH9M3iBKlGiLGhDgstqpCao3wHVriSWAS/AE92Ya1PHwEf+zmE0joNzyNy
hqU7gTfGpicCzx6SJ2aoujzaKkG/kOcWEFRuBozUus0z2U141R9GHXGnKSYU
2eTb1m1R5du1F+B/6fhHkymh0v6Kzm7J4WJLWxnvgN2Vl/EsTdm84jFCho1/
UbHgdkxZ0zKfkoFFeoIj5TFp4sSuUwDBvMyG/hCxDQltd/jpdYMmHWzXR4Sw
u8DY3bsX2FT5E8EwKLtBXLTPQCfwydd6LShhvHS5wcqqkOYv8wZrTIhwiMh0
POdwh8tBuFqddrLyitBfqwgoEgz4fVjTCbnNdkMNTI6ADZltAHt6W19HLZ1k
TmzUnMqWRE2voQhN8i5hId/anRjBVCVRf09q31Tx4e8WcvWiH4CZUVGsZOCL
aMCsTnFd6R8sN67uXB4qvLdy5CN7ouEJT8OCdzgoJRxpEdhboqtwB3mhqt/S
y+Redmepjou28nWqSbzjP1uEc0uDckJuBgTvrFkayOiiO1Bh2tMZD5OkQgz1
y8+IFXMtz5b8xNsm5vk1a13xe2Lo3Zf5rT7yI0QnAKHmfY+Yt07gqHDjaxCm
0LMqwTglc9yBSVogxys3WPBAsThgDWLJvDKb80DxaiTZnU71ZKPxaZdWJggh
YmruMqV4OpJodyL0T0oVLROuWjqJXCr7X6T7emnnMplq3sps+kURhBkA2cre
NG5vNz4Rh6No69jnT5IDk81oC1MgBktzTO/sdBlYSqx8ueoMCSgv2KJq5/Te
9I0hmz0kwUd9fRHM444XXwwaZqyk7+oE0J8RHNeXBxR0r5NMquSYoMUE8eP+
993Us8FgV4Sb2K1RA9p7mvjl9NWTUfi2hWHSzK1dB+53metPLkJZfgS9ZKKH
vtCORq5jncgELO6XFC+aeTLHalQBR8mF74pYnmd04eYTwsxT8KDVCOTti8Sy
siGENZkOPKutd7+Lsd5FLGnnR+0NV3Dh2Xz1V6mbHtXLaHOYpeJrn2waNGV1
ANpV2XT6qG3eysFWEKhzDuPNku2vJsKl3ksWhKChADmetNCQugGeihcwCSRR
yQ3mJyRtbDuSd4pF5X51K9+26gXP0u5MiHC0NnWeMh4wBoVBLRGYBomGK4MN
FCiPEixjgEXHtv6cjaFdK4N1rLZXKBbF9vZo0UzOJ+MWOocaOzSw9nYpJA5L
ueUQaMAIgxLI6y3//YXUxKtyniDF4YWXJxdRZKVwNxBxUDoYsWqbR7uAdqo9
I7xsSaFbFjf3nx/gHq6wtHgYjpNp8WgMPbPQWCbTeXgqyLk4oFqm2L74TWHp
cAeQ80eFnIQGJK2UERJCB5HZyLX0Yodpcxz0xBPfgp5ZLZ3lRjRVWc7cqZ9/
BEbsLtObpbEsmwFvbVctJzbR4Qh1g1AZk39aP7jqHPdXVKP2+/JeQqMtZYeK
+eszO1BT83Qi4bAodqZC2ygKTrjCVb1uAotxcEC8w7Ze023ZPqN8JZSsQ6bk
aO1zfvr/vsIZjQwrgYUY7JuxKfQjFDmlbQa66EjTLUfiJAaH7n9uidhgHDHt
ihYmb16QL0imTdX7OrHG14WW2jts47+wbMmN45BB3zaflY6Ei0cATkQntbhZ
MfI5IVkzEZ3T5pmTafs0GNZv2BPwPxlg9e6/ZCK1wl3Jes2OuKHtBedyezuu
q3hFvs8JRqB2olfc+l7fNyql+u5za5irCUsFngwqaKaySUG6n2//aW8HPMRP
C77IUmicwOPIBh80DBeMdfTIYhGwzhY9c/KwUAR3qHH1YRl7/4IC6zD/Pe4b
o3YOzv9KpDN1nK5ykBgdOsF3w7NhqTxxOh+2Ddrv4HiMAx4gxoEZYJ/1hcWz
EWwZg92pC0AjXu5S6/D8hj934J89TPRpQ/eaEpHqnzNUizPfigAmtLXSIff2
Za/E+6T7QrGyAA5tAPYMdujOP78yG3i+cZxTEuVs0D4s3cCsCfwZ1s+AAeCz
grKcJABAMTjKKAcmpKnmXyVPeDEmbfFUjdDX761bIyx3Rnw5kOtWjJ8T7Sf4
jHmoGiqDkHywDpKr161f56gFomk50x4mkiDubETqgsJMR72bKBKkYKi2swVX
9PRkVsC7xuqVkP8CpovUpZtqn8teKkKLhKnjhzhmtwp7C6R27D4vs9TeTCuV
TX6bYMpQRjZ1CjIV0Kx4uZ3EAm4AAgtOCoIbMys8kt69otvpRbtdPZGfQRzW
X/+Cyo+9+8Kw04SxrwR98Tugnv79gWXhP2ypl8zgIDHO+KyZoctV4wI1ybkU
ixFCUhCrHpVuoqQWkwpf/lIdk6KBW6tPMrDBrgYcOp74hUfbGxJMZKmpnWfM
SRjVC/f38szBLEDN7S+/jVI7OYfXsfdycQFTv3l/rKBkukc7JHbsqAvAfKLL
+J4i8EzTfG++1NWGzUH9/9DHcfB1jDluMZLefwGwd1JeCxuimJ98rOgQ+XuT
81oauKeseKOgt4zzNCtlFEwMGdpEAgQ5Tus3xCf+8A/yRCim57+Ll/N6ZjcY
1ShWb9y0pt7rjIVUI8LF+V1VTZv/I+Vd2mgJKFoSxty3FLAcDayj1ja5IpLa
0Lke0yEgF21KOzT5HA2+Yz/ugp4j9wcnhGRe/wAAmFKNQs67xmB+OkrVyStY
BH9pP2FLeclEtPua+FUmg6o/7bobG+1eiQtfyRWXYwQWk+VlbSGaquybOee5
QdGktqMIpciHAhhrkRUtAdjlJMvbCcbv+8Dp01wL/BD6lUJenHyDeIkr3wC9
Zmm/TIauXA41gX0aMxKOirFYZkm/w38vqXTqi4mWy6eezSzDRml0ESLbYN9p
+QSTUP61WRmNSmsZGydvVJ47qydVukb2QGTWyUwrcmzwmXbLxI+ahyu3i4Gw
O0pHbOowY4q8RonRLOFtDRxK94Ao8fwiGWc9+iirBhe0/FywtdL6C09Lf/Bf
s9jn6xwrIQXgeQPaoZIJ/xp0sJigisT34x2l+gpa8+yApcKDja6t5IFdzQVu
MGcpByEPDNuFUQ6/YBpYfAI543tGs0+SdSkwuiUhehcA6MnqueGicotnVYOT
iK9A/RPPbpWfb7RcNZFXpaKJhXvHncYtoeNlWHejBOwJiPCMoG/+PTpkmxU0
cl3on/7BrMZJ02Vd4+ZhQ1p6ze4FZDK1i0NU5BtC1y4AR18vS0AuVJjYO6Bn
CLPM8+rATqOMbDEJoPSUBud33Jr/dCDk7/kIVptSABa7ZXEQR/BlB2ea5yKW
a5z7eMxo0AYJhtzHS618p/mvakqxIcq9KGb2GFBufuhhCgVIUQAuuyjjYOql
juZIES3BxScS+7zX48Vfp5EzFq3sAyk9vD8jiSv0blkiayNGYSfBdZV1OgeN
w9mnZq/Z1jjwpkJwqVLNC7zFfyaUr82hXMZj1t8eCGbMlv9n5v3+RIRQfMdx
llm1KmM2Mx1zyH5s9gIxwMMjrzZ57tRV2IqIicxo94U8P+jbGYDTLMunujhg
4U3FvUMX7v6y3wFBR1obJGhM+0u1mIoq9ijs69DF95O8kRex4F4iwMNYdPn8
MZWK+ikhxvJBXBYNRTNHJdUpBwDEgSGgF0sWs45fOn1AnPClUcDONFaJ69pd
196PWO8zbPNw3v3iJ85oHbudKAnMvUMmOm3VL29Kb/lhhYIqm9/dUJ3k/6DX
SY/6MOL7bui3SSnMx37SkoR3KLkiGgxzTAZQmVRhXLoEQJ0Ibo4JlgWJ2+zJ
rGmq/nWw267eaA1RVMms1sIvfYlJBBpvU42SX1ZbbUY+7ZhnxiY0PxTFx28V
YYy9K2HbtR6EWHC6iSvnUwo7fN1JWK3NnQRSAlR/Ke9F2VoO7Gk8HukddtA+
O4PbrxsbHsdnFV2WBd6Vxe8Z8zaPV2g2rh+V55ggfPRozmX/6SnB/ps790xC
sqZMfAhwySEGKApj7S07KsQkQffuFNvS5WgXeQSeo87/b6iAK8KYBAVi+DvJ
dk5kqMkTMOlJdESidIfz49cwvlesbvGN+xN1pXalb2Jbc/nhpQ+lWnli7/OT
oZRmWRTprBtB+fxO74pN6VZGczwMcoXbfLwM9xdZk2qvmTM/oTeGDQrMEoXr
2kn/fBh9uMqFlZTvpjGwB1u5kjNYQ/9jZ6yVnvDOUdA8Z675oxsIaNQmqPvj
DzDiDsUu6DqkI/bS3Gu9mb1PlIAy3exTWUFz0NqZmDpgysck5TqfEOh3nDYf
Am4BAsYYRvRFnPKcTVVsrnGiZsV2YKpbdyJM1DR6dbm0ngQcxGmQPEQIh7+X
5Wj7nZYAcJNUrbssMifzxqsc0Mgk+cTJdqJFf0vBGRuUBYIFDShD4h1zWeif
FmbZneRHwXXdpuFy1j2QzRR2MXeYG7pwzjhkPObdrTgcEkLEHdIUU4dSp/Xc
VAPZToClTYsInAOx7O8HIegVowM7g/TXiAleQvCBMyVTBH0qLrt9L6wj32cB
QGoT9HReK8tkFkzpAHUStJu/E0kzFKNnjYME8O7kSh5mho36JuCEdRj55nA7
Ai/LFdbg1ip3KM+fTOhdHUnn+4BUoJon0PlpSnH8jo0j6kchrNB1/WeO6BD3
ezBmEbQTwUwul26bkVsr2JGM1UQ4J2oVzbra4w/1Rab52XI7aB2vttU09oSu
5VVCc9vbxhaVNNLlgYOxQ49b88RBd01wJzynEa/IYNtT3SKiTq+ABk7DlKSO
Vq1991TpZv1tl3otfS+/QNDtAM68xwzAYeOFhT+x/1Ei75unURoJHz3ACylZ
iG6hnuvxlYmYhnHt03r4GAJ69VG4GnnJffI4cBLGtUbXonSetBarMfdH9TL0
kf0FkypI5rGfdmGzQOja1wTMCxm/M80oL19p1ifLKYjp1MZMcN5RO1DyYKOD
3yrt47vpQG9h5tAaS67yf2tvLReaDOWgukohiDKwyIYjvkZBLRNxLoU5mst9
iK13gpFFc7ZjilRP9B0vpRJUlKjNkCTShnKjgIp2u1yrHE81GOnYecKMILbz
8M8y0Ksbjq2euvL0CaEkGNMCNbEfxNaoDGIBMGlYxU2jLNLpr2nQ8Wsp64ld
coc1bcoo+OE4K5zPsJBVycxyuzzcweD5mADfk1nqOkoezakgkDKjVAJQRReb
PdIhCgJoOTdT2m8bXvpNyUw+1i2J0ourO+mZgHIQzH5Rq5ixtVB0bi+Ackt0
gGnajDq7LSiFlNhpYgEfqn5+KP9XbD/Qv7jteRQr9z+VV09Z0cPt4iPXsiod
hcyigSXF7nXANMlLJBFjlqSjxP8eV/DxPw7ig76gXVbh+8eiYPFWqFkwFTAv
3DtuJu8hCriUi4l/VAk9SIpb+iH4++EKi9NqknQVBSHuESAA/YTrZDkjavbn
0XXkHbpBY9uH+KyopdUsYjzwOc4F44uMyjm8ntD18wfgKaZ6Kc64vNdib5vG
i4rX2Uz11EDf8dzkNBjqmNGD6gVZImEu0IdT0JSdvPWt5p01I4v8jqfIYbGz
fmfwrk28qlJtLORTRioMzMaWXdwlW2/MINc7A0kFnC3a0L9EQ3BkTEH85Y+P
GAWsusEBQ4pjS7gK2/q009uya4gB4vvIqBCrK8GrzWw9jaGUja0G+LEo1yqp
pwRF+AZGPUKyw9IVUA6Jtx+PseYw8hwpfn2CmPzWC38NBdJ4HzrxFdhLYJGz
E/5/gF1Fp+AvPERB3G0zeN2AG3tsXHVRG4QE1KVQN5U0OQucvpcKTYbuhGoX
No5wlDaUii6nI09MoYW5Jq0ahMcEZlTYFLmbrvXinwsTqGXt1vNHIDS9gwr5
AOnZcoQdmCKXIBv44riu99ZBbZP5+p192ZJhsqvnvr1gfZokq5gBR+mdJJRn
+yemkgpwnyqur/8vBAyhCmHWYeAEZb9ofefaYF0gLwyfd+F5KbYITDV25OV0
lMnF8PAWyrN89tNFP7nNzEG1IHfMde9v6KMmj2IX6cg/EEDzuZhX+TCPm7z7
OypTEp232DnD1k0zhJQChz3mqXQICqVCzFt3amwDIuQaFSfwRlJa96k5D9ll
egZz+jAZYXz/n/IDpF/RhfYUulvZKbS9PTvNfNlHqibKuOCl4+qFdxzA3P91
H0Ex7/55tKBX6fTP8rh5nf/t5KCRZECsgYYa1dffQ1SC3SoQVxIpdB3nsJJK
3UQehr2NiQvyF5DN7BBe1z/hu5G95XqwfgD4GtHAm/Xj3CnanDIwXff7ZayG
nF9S1/cBLMupZWb5dxswGGO+Hteb+VyoydSqhFqw7m2XyOXR18AZsab993wm
+ziqpxr80r+llp1an1x5xn3+GsiykhaMHOTFYri40UE9bmrjGIABB+O95gEi
RjkDenLRCcNlKNlLxaVkn9P/4uqpE81aQ6w5vWE2cbEqJIwdULMXnoMDZ+86
U64233Nsk3N/OV+TwodkdTF6pL8AKMFnt/YntMD287wBQfXjmS0hyXK8xVSX
AL0v7Avg1w89BB9tQ939zYKl4L7Dsad4j86mUwqhkk+Zu6TUZNXaKnH6cEnz
Yke3LMgkdfYzDWo8Vq9Grr6nORSiTvtQZb426Bff4Nnaij3JFMHjHVgMSw/d
YZmyonVUt6R7RbJ8Uy0doViQ6lcDQHsdAUNnCl1f280faYoYI3DonzDpzvyg
26bW+tvFEWb2G14UojWK14gKjAERCpmmYdXPLYyM6cJ7qjiNi/Tx/FNOsqcz
cOo90o+Gnsy5Ci4ko8vhwL6RbVyQZjEmJeJD+F0q2UZE3t9mTwkztIux0KgC
+w6Y3SYoQG6wcc7OQnQ/BwD/LEg8hCOtrgQ79X62Ry8a50m16do7PQx3AuMj
cidlfuXBuj6YftM09HCVap7Ald+Nf7cyVGxUIophz70G6tCm6xqZRGGI/4iO
1RqTKToNYI/AjryxVEHxLhQZKuiwlqLxv5qMVEOHtEjUYUCHI5HZ4Lbn50SU
WnDZiNw/Ahm220JLHbhUJnCKedlppPgUd8HDFzqdi8k1kVxoSlC94i7oAmoe
qtWf4WBJmXb5ISRxx7T6oznmspg0so0ATyGVMXXMepM6xyHj9+hItfH4JD7j
49erXB2pAukgY2K/nuVm9SH39N8mVamXoPewdC2DZHs7fDBPum+26Oh5bEq8
v90RzKxWRGcGqNUG5oYMY9NrnMEdALHvADPsjcdBMrsK8fBsw+MUXBuYDxhA
0Un9CAblNDdwmwjCvOShxMZaw7trnlmmh5yxpmu/plw+3eq6XGD1xFnTeMZm
+VJ/XRqISeiy9v+OdgKnP6RnsKWHjlEl9FgcnPf/6AAc0+HuxtotIkl3+QeN
nIExV0eB1TpmhhI1iUvxCyu90/oEi/EPyZP8DgzDlLA5ZxvonHkOVfJhlmBF
6UWZDNlQPwhItynOXCBvI3qNWAHhj13p6Izgj1GhGAwC+1KnVH/423BJaH0g
tFdhJUHM3Dzq+05yBKTOWvCQaL/qIcFxG+Rsm0K6UlWP9QTIlwOMsqP4qxy2
Z9uqQjxy6BCozZmW0Tf3GsKFt9RcE6VvNEC3i/dNq58XiI/rPdmrbg8/8DJQ
u3DjanHb5uqyAw06xvfC77+F8qCAFjQiTJ/7ineJLa9jooEyHLN0bHPmFR0a
cj2lobkO7FYVWexy0MVcCSNDQ/qTgm13J/ewSnNcEFGzK7diJlbQhY9W69uy
1MR5jl0TotshW8WIv87fYuuPmb/EP9zI4Oc5WVeNtwLE+nhsbKu8XRl3WwXc
0QFtZgPzz7jLbxnkGxNN5y8CNYqQVZoV59hNsuqkM88gd61PmRBRM+xLKYev
hXOnwvoQGO6xCTYhgrY00dkBlRKjh59ovGZDG/pMjHvqj5tpDIoAIL+ngXo6
R+jH8fz4Kv+6M0lUMiWQ7uMybxxcoPaMiTTQixBFjlK2wahavI0G6IYJ+5hD
Pcwyb/+XHcmikQfzV3RfupGxooaEhS/Qs3YnG8DuY7jHsdNImC5CWx8wBdkz
apwUrT74T0cWssG1J3qwljFDpHkf3KSnIuDVEWstnrCY+lfzEUP0ZxGAZggm
nn1UjYkO3ThZ8heEaUPb6beaN61mq+DW0hoAYyVji+gpthhk5U/QFLei5nCv
CoH/MhLLqefEXHqaq81A6o7e92iVMn4atm16S7e6D2JD4iJzL9q6ByBhC03p
rcVLkYe7Eg5q5DMmw98XkxkCa0erUmDalRKvYY1AlS9E7ZtFH5OMFpUUDcQI
xYqdx+heg278vk6xbDbMHS/3K/WjTh905K0oYDb64+bgKRRalmkixtp6bdSn
sIQWa1P1SQPEFCZwuKDlomKktNr4Viw7qRYXm2Qoq7lFkBTpkBSz0ojx8485
X4ZjvYSu9T8gQTdRNVgHAxst3Tsnvb9DeTru+XFSPpFcTt4xodrNCI4m1vdW
fNrmEAGPV0EwRNpmNg02UmVKvFEGMvT7hE8YBK9gECj7TLG5bXyzjodUMjIg
BNYmnnVU7FF2eK+4zZM+LsRZDaIVkoFPyD4yHPXdKjEg8xbJTqT557v8PSSb
3BaKeDgdyov5dUs3rHFF/P3tGMoqi5K1ipzJ+5aN37jj9ck6HI05HfMtNYB4
EuYfCMhXrL5A0Dcw8gtXyg+Mhg2/OV6hVB9QQp2OaoXfyjti+Ozk5EdgWIoM
4KzH5RMj+CQhASG9fSxDbQpwU4PNc5IcSYINmvGHVQ4AE5k6lhZG0XmkA6mW
WAhDI4YRAnVezC5KxgN45xTjgTurVOV1RxAtiXhSkvqohvcqo8SC7Is6963J
80ynKpc8WwISfbsxIjnRx7zZIJ1Sda5DJNmStuj4GDeSknZSWrnh3cy00m5y
Tnt79NQtn5l1C2boe5OA9zS9lkpNuMHv6DNzWj8LvPAZwrf0BJGLEF6KCpxq
WuweGz58qBTJCEDGPOngXuFWBLzqKwm7Y2+WfSVuse8jEPtf0izptIe9OD2u
ptaw3Xkt0B/DAamk5uGvE+11Sk1/Dn1q5flCeMXCPj/47Fu8ydsudA2bWbad
/bRkzcASoaHV/l4lu20OehJQKD3nlq40cOUSLB0Jwxob6x4lF8OVALd5CY4j
Uaqu7F/a1vFi3Xhw77WN5KRHlYJqCgFZuHqSBoRNn1hNL6zZbET7Wgkn/SZL
N4OM1nz0s5h6UDENTGyMhsOxV6SF/YM+xNs4gpLsGeanstV6eNpgFsst+RUd
tGNGanDLXI0JKJ3tzE+Phdbl231bPgz/94kc2GPx3HvKvSzI3V3ytmynuhS8
WCiuCm702/L5RBek3wEQ0vjKHhqqVHLPdHG5D2OyVgnWic3kLgTGlNoNY6hz
9151yGnD4/ixNeJVS1s9q61gl75r4fkiRo93u5QpPsPWqO5kWbGeuRB9NRWe
hn17NoAYremXLPIkgEHgxgh50nqnQTJCe0jMYVdKX7rzAQx7NZggnBCVWT8D
NquAa8r4apbJnQkkazBq/sy7jql/GL0wbroLZF6lUHPA3XMXCI0jVJBSd0J0
EzSEvRcSO/GQUCLJPoJk7K4fj+EV+nsjhTROGozoVAOiCzrs+T4c9pyxM3e8
D4jXJuwQ+mBpRexsazG+/Auojqi6nPMV5Yqx8TIlWn3CW9vFiMxdNqJX7IEn
OwJcX8CwToPf6HTG4Zvep0CF5tCsuINr2FnMsrRfQkuibZAe5HgRrBhOOjwK
ipl7wVLU229zNBZGBLmcqgAzfR/d0I6kw0BYWGOL9IV1PnJ979mbVqnAegd0
dJ0UC7jxY60q1MTAcJIq8brT9B6aFLdCXswXz7rus3P8kyPD8UYs2aob22fi
muciiu4qxRDvHY6uD6sSUzP9MxJZuqLk2nuPGlJYTs+JdZehd5fmQFWMJJm0
Ht8c8fCp1qkcX78AQL4bw+rh/1/ZEAXFQKlhMjRF+WkOfUcJJj9RDHd8eWr3
gLJ/I/H6xLt79SYR4zEf3A4VGKqk1UcIEAoCpx5WOtUDdFfTmEgdmh7CZMu9
fZRrWX+eXH9pcr4zg/h1bYKommUkB0v6qCUiSFiYD1l/gA7aJVIwP+QEwVEz
UDllVNcvnC0eHD9C6Lk+GY82IOUUu7a484VuWS5/Ul6cH9/jIEIpJiCOYZxk
k594j9+zHGP1iRSW7dulkEnqzsOL/WWq492lyjeCsxPp5vh7zvGF1Vq4puN6
l6rdPKhdqXmAtqSrtEpHKy9wPGMg4vHxyJW2DyX6ILTLbRXaN8QFFgTyUbED
Ax3jUY699ElsvvyjnCVQf/5w+sbYk60IP1VThh9S3dj9lgSbhAe3ZGhWxq7t
UgeCtD3fsMF9ABU22tRR/i7SKay3TTR2xgSCbLanOLfBbGy10HK4/gQTdTYc
ziEoKG5u6Q9kK4+Q7jX2EVoMpSLb1X1DPUkbRRh3ZpIJ/y4kFP237RPK6qO4
wECId0dc+xFAYydumUblm1HiDcvEIpSdZspMashLyu85ZE5VOUBWiQG62xi0
iSENLiA3TK6OnRSyluj4JHO6xuSVM2xQWiDpURwegeEstAwiHnJmd6TX2I3e
hFkfZrhEU2ajOigRLGTAZ/zmpisp9GELizLE53UCH2WlVN9nAxBLYin0kjFs
lawjWGPbsN7xENm8pIBhMY0hIvy0tWH1vxikHyGJzIFOSGMomYePPyo4uhdN
6aeF74tZketLobStYV9xRR10/F4HbmFYAfWeV3BvVahw9D7LlBt5jIO67JT0
TH29AuEUrIItESz8nMEDmuRDpesTqJnkJbVYqDaIrNyFWHRzIgHF81Kw0xYW
Zoka18LWoTGuvfXqIqzyBgt5z9BxXy+UD4ksjt1q6YnWJNVXN4uIENv/NWny
lc/mPXAFprWStohQ4fmnHc8zWqlYT+Phiv+3+7j2ZAUykPJlRkm6gSyESOpu
xY9LwpecgCV6wfwbMfHM5CVwkggBylQJSY2PvWCF6AeRIc8Y87pmahZGwCEU
8O0SSOLriX6xLhABM2hs/9D0vsg8z49pdRp3uoNrpqNVt+rbjsu58BWXQhiq
hryXSUaZxc8C77Bd1ztdl9/7PioKA/TosA2iyZKRHV+Uc7EepxZwVBnfVxOl
uhcGIJoBDWegbOtYjMYuZZgxqjiN6LDubLid265tR0vmS8+8kg5CJfwQKcDo
qHOSD3S6++Sv39yN8M/gLjQU/VNVfkitRZ+I3+CCpoov2juxTZTML/fGOuNO
m+DjL+opekMpIZCyJdZQ93o9ulnwpdqcu1WA18NwsxviKNb3goaBSCy++rtS
gMmpKUU4v4Ai6/oCwgrpSHp0jFK+EZ/PNTvVEbFxtcvkPXa+A4q86GQS7pxd
3bcOY/31FFv6YXvTgXb1j3bPEv4OTm2oBz2MFpPIP3IDXkhrcPQH31JslZo0
uQfKrzDf7Anp7465f9w1fHIKATDYSd7WOLSbG5CbNzvn1ZuYQcixPidysm32
7eG9Hjaq7by4xreJZ7rWm3oTCbJSgHSPqpiwGqFrIZHWHudcG/JIB7s8LsKJ
jH9bLQzkR+Bn5xLgfqhgQ9ZcYMyTkoHHSZO74tSh/99d5KKRxXRIebZU8bfM
WMbMtXGWw/a3jGGqeXPpSuzQPVPK9xcN0ahrxvPgrVfjjSVfzP5CM2Gojmvo
IB0nbXFHBNpF9yYU7RC5oQ3FNOIAhxkK/oM/U8MGcdlxaA0LSEupf2NTi8Pf
dbb2q7Le+jeflztjVQklvayhfJFsVkxXzbk6y6bgIvhIH4SU9TxayRp4abJJ
c6GTbBOzTM8ctgrHqPXfl4fDj3PtJNgIFJMnR32MJ4jEC7U10WfI8Ua7ZF1K
aTpJSEH8HOUGavxkQICDLBw/Ki9wXK62urZgF3ExusGC48A2q+poVYN/6dKu
SzEXhpzPoO07nWEnpi+BzQmvXumNptqc/jkaIJtjWvA9TmgkXQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1ITFcsoRrMpijH0gJS4gWrIAtKbsGwEUK1u25S00/3xY9TRsWT4xms/tB29BWzQyMnlt1AQScYfOpFocl6oEA1gO1Wk10z1W39q+T0vyJmm3InTBMHozQrgdnb3iNp/P5otEXMxsbulICZCKEJ3JCAEdrDIHfL83iZdy2sYVVNk/khqSfAtQyRTFl3v7lhnxqvvcxgGo7stszKZPoxOu6y51ef06KKDmMtPKMLvNmskJyUdP/iZr5QPFbjqTSAtA0VVOVNPGS0/NVQ/occ2O3YxmhYmw3mT9U68vG1c5TWIwXfWKYmOKcb0KIcLx0kAPpZuBwR/Tq4bo+jNEuE7/2Fk+FlEqwWiTOvAPp/zTRnfm0CvhBX3Bixvon88hLazyklj6jbj50M/ThuZEiWz4wu83g8yQm1FqVPhTB/eW5o/0mTHbrup5IgFyJ3LSapYO/aB1QsgFzgMnIUaYQmf8TYKumxa5zTCl89/tbVDOD5df6LAZfD6Lkmx/UPNY5+mD/532yySh+20rjPELVMKj9bY8j2O6ZeuWpB77LHZPEJPsyElQmJ14+0yz7J5VGQPudMoAN2Wk7VafeEGRk0hAix3/A+qsXgB89XQ07kUB/rGihNvWBL+YL7BEGFfeazMdeC+kBMVPVbPLq1b0t3Lq0+hknSii+Bd4ESpK5lPhi4Cbm0zryLe72LSFfcKz5sf31WwJmPz2wxqJyzNRVKJEUmkwBFDB629uF1dFh8Hf15SygqO68OGsYt3BvriSZHolJLEeVNQV30tgBCkUNdMh51e"
`endif