// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SMs6XTiJSCSA7KgT8Wjms4z0IB7LZeRPaKoLKY2apmHgttrSUPLKupaUEOcO
eEoG/93u2vqioyaqkuiNfIW9makR1F/i9vQFQTB88CiNV+7o7hB+inkXDpH/
CwU+5ZUzaj7A4FHAgAU2RS01MavnQbIUL3ubz/ve4w9Y+bj7WwZmp/8fALip
i1j494/vCoQrEEMlAdfc1/YJB+mE9Wdd+D7IZmp97yImNgzom54Em3LzmoCZ
tdAOsOHsfp3BZgt5bnZm3VzyHzYauoZOyko/NnVTdpxbuA7Pk4PajHdUu0dT
ou7hwHZVQcbgoBsc5rxBgTgniBMqBz1k8nPXXA+NuQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HDRiWScCL8MZNscKJankVYerxUl6FFUQyimOE5XlTjzetPEhgsF8z+Mq1Lwb
spEvz8ybEx5xYJowzRVzB4H3sEp6Tl7Bzck8xirGjDwVZYvIs0ktv6HioA4l
S79p5x1jwGqmZam33kXstR5xN6vatBa5ASVABKkANPzWFkRlO+YLRx55cea+
uGCE5E835boSTdF0UBvpDCwapggbOUQ8I10zYjZoOwCwBEz47gfua74YeFlb
qwKlxLlGYRo9+cCloPzRHU1HZ623VkLKt4w84MN9v4ySkJJmfGhOiQRgGIyk
P1lHWIehPXUwZDRBEHXQvkE90tcPfF76DeM+WsI7Rg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GTFgJInQOqQTJxxKr3ZT+iN3ep14pZpORDSi2Iar17dcEYzL2ae0EZw27gcX
RU7LXPCzXS4QGSLrpONZB7RDRsNL3TkNrYWND3dgaawJ6CeqRbbrDKw7VTpj
jm4hTQup4Wpkd24WyOdOzw8GxvVDDYmnz7T6s6W2sYP3JJWPBoXYtrhKnAjL
icnMQJKQGKooGClTGvw55ST4fdNkl/hzQTEa15Zlobs3GaPCAjl3IHWtrxVV
5JhESOBMD5HG5TbCGDUdXCGcPRFFjOznhOvZ5U6fdzhpysc1EsmkowJAfd2A
zj5Kl0hcFgcVQj/Fgjh/5JAiMscFwIH6ILeIZozoJg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SqtcZTqke+uoXfJyDBQubKmAXsv6zXLH2XK3lbhIwiHh2wFu9iEtENrJwMDZ
0Koqxd7bIJixuR13UA632lQBN7THbpUGuvvTe9wnaAR7ZGBFcywnxmvcNfW+
/YQip8AHJnZ6RpsQ7z7KOVy+1gvc7rYP9a3ufMFg+GueyJEiPVRmYi/FPL1Z
lhFqTCffdJXiNLgrUOU5WGOG6gHhKC09z9wS/kOnW9jX+ipTjyPPt2AaOyK8
2O4UUF5Obl0kDmdAzzglfu5KejWMORVAi17T+gke4n/iOe/dicMlUmd3Ug0S
O7ntX5pxIZfuL9J0nKqpDS8ymnAQtww/ruMW0YynjA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T3LJlP9uPzFvo7BNB+bgA/LJ0P3OKWRJwxHZ/Vm2ydFveLwgegz5/Vl535fU
bEe32jVNEvdAPR31Ms7qnhV5jEfJoKYYVBEUqxKzXn2g94NILlW1z9MaWeyH
z+ckpUiaBxEObl4CTkPAURPEcIS/+JEJo/A7I+0nxfnUuntLQq4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Uvz0SzacWfV6SQrqXRQBARYe9pLw5IKWJuARQdFv2MKqtXXBZ83pVp//0gEM
lWzXFw+7PjIKNl3WEPea29KFNaEdXWneG1KTi8w+vca+TNaC82bL/gNm6nnh
AmXbURacjmaK7n676TRt8LLB5Tui0pdcm3JrEGqupl6hEPiL/LSGdO/xHsM/
B6FqVKqV0XH3okai7JDOqvJ6b4kIR4JX9oWmkwg1ttLwYAyToqHSLvhfdCdu
G6XuwTSCGWS3/PtDLeeVXfBbATk45p+1LXL/GCAcrUACjq1mgKW05G7lzXMS
huSe3rTC8cvvEJuQ6hq/xkf9mXcvrd+xUDfz/OEycsoWjxGsapj6QP3UEBK3
r3UT2Og2cVLq1xYNXPT/5KZo5zkla2IUpUVhEyA6y264p7rVoZKjQoDfi1DJ
4rUMf2mLQcI140YLzEa5O/gS25fh7CF5FP3q8LqyoDwMi9IcvTRH/KHVOQl1
4mTqYGLfu2I8nuoqJMWzIikq0m5dXW21


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kgt2TolE2EnhVIP3ugX1oKSSsbQSCiS0X0N8K0HaP7YWkiSaGHuk0teCVByA
B47zCRmjcsr0XOgqSCIGeaDtvP8n7RSmpZc7yS3uKHtm1K5DqvBelKfHJ7Cu
VY6oTFEfjHOTBHpAVn18vDC1fQtTkPZZ4XVO+bchbRpg/SH+KbA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eWgOf4hElg1/TMO8SH4iGQpolo958Boh0Jc4TbDxH17ZFSYobdfD2C5hcQkb
qpbgMpHqRU5FBwo9/TupvZaFNgHNKzvQ8CEXypTzvGv4T34y2HbSqBtzTKRd
yvFie706Tx4EOcfTMYpPtYgLJOQupJP6WXN+kER5CNBm7Ic6V0I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1056)
`pragma protect data_block
Y9O/1h3ae7ZNlAljU8DMqKpoRE24klLwkuShSNQagRl7zMepIvmweuY+iBto
E6TpxnBilLPpTwM+D7ol+KJOb4oVNrJV+oAzH2RSUjeXRbTB7jCa32t7XRzP
4f6PbJxIB5cgV75aVVDk7YB/Xy0t79zyiadCZbXJqJgUXb1GOeL83Dj+zCOV
tEt+v4//ZxX13KpAZk43lcclsplphcEyr821i0DS7tDLvdTory7Yf9YbZecm
LXrUxJ1yu4hb7mOJ8nM1SlCKa6R3RPV7pSAwNxgjUwri/7lUJWVCB7lfhx+C
uR4mEmAyomzxz0pVUrgRoqBZThkU9btbrK0aCIegACUURayG9mrvTKmpppCO
gknFbGaLqLEu9mo+RyTbI897lZamhGev8800wnHMFQzmZ8kf8qXsh7g4lmHs
k8cysi+PIfNOjSgbVoamaBgFGso2gt0o919nbXNe6bKMwvgdcczd5tRKYCOJ
gsz8fF+l+aVQvSP5XBb0vGQqsmptCjw7OK11gXQWjNmaBIo7ojMgfcs8jqgv
7mRqpo0iAOX6EUsphp8zj+g5REpqn4AZYKsA4dLeg9/IA1BbLSootjfZKBDC
Vy91Cq22qG1afxlPNbI9ac6R70LmtPa6SzEnTT0v8wLfx3I/74USk02AeqwL
LdJHKYNIei4ytaIdCT+koi+NFL4bTbwBfMEHVP/A20rWwICY2ISwFNVv3lrp
eQRbEuwjEd+cwBq1zSNskKdTBm44pLaVn3zGRIY1DIh7KmO3DbsvECupXcAh
w8eFp2BZgJiRRK78ZtD2A/uklnuXnPtddahmMXiDPURXoOj4ROJUphqKbcxh
+nijT4z3beTyHGkItk6eRnlIpdqP3Kk+lnpfCfr7BhjHriiyj3r8rCR9eXoA
RcATmSK+LLJEcy03VeBldMLg8jHjso8oTQnjOqWjHObquw4UhiyMAaRwRMCE
IP9vpkPbxPehHD2KxA1ZEiU6GIz+TFqTtlvJhJbLF/BFRS/KSSgeCeGUC3eB
s3VHMlDfFitZRXUVraxreMzAMt3EMokkbacdXsSbM6qmBLZEK2BxNO+7jr4p
BqQDuQ7cmwnO73l6JFO2x9G0xLg1O0jrZ2IJjcVGaDpVdo7QVHO6hxFs6szK
+KdndvwBiVUhppTVOYWEMZBtCJjQ5re/A3E1UD8aEsTSQJSb6zXJBP3dTnUs
QR0+sFiUIr3b6AmkYnbPPBJvNFmB6NNN+N3iCzp9sva5tW+cDEHLBFH0pQ5M
8MDBz0MUy6kIEfrrlGiibCwyqxQzyNtlf6dIPIc6mat5V+jU1hZ0U5Dxnc+R
j4iSVg6jOmVu/kmKOSYBNTKmgiM66GOu4Q6KndH1Jl8X4vJtsFRbEkqIRWih
reLW5T+0uTrOIZCwDlAOU7hFY8tK

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdiSocHTcTfMWpsYDEBFvdyZyCuNCD4lLuMKIjk/sQ2hxaWEkX8LUTrgfalQKYaZ5B6KGNafOy30CvSC4PUfkahfJrBjOKHhPpSBJ1i/mBZzZCHipH3jJfkCApPdQhRQWdVzgEg8iufFwFXKUzyIzkHCjgkoSmWPkzMuKSAgZjNcLwQAPzZ/2lnA8JmEX8Csrc0lbYlj/soVd0fztPHslFKUSUyI6zbmGriNO1KzALq0aleRYtPuF3ribkrzgHigxcZOdF3TRLtfyMh5dB3YKh2mbiZ1CcddTD0skqpJrXJ6tJoSKmdFHg+NmJFZm/71QPFCfW6/H4EIPDBqVS4xH+ymZUmiytHMimhBQ5NvLrQy996Yy5sf2YYckHd411f7OXzvbuSBkCSSmS2GYdfur9PAPNFjXUU0wxyhAhRv+wH+CzebA/pr4J+048oMhmbvsOJAwRyF9aJ7Kb/Wkqp0SCm6hIq6KfgIDQV6fESZ+3L+pEhMnkRBkw9uU0ZntRLEWdmyeBE6MTWBQw9WBbno7IbP4Pi/24EyS+QwGENWQQwI0pOESHpuBBTZBuy2a/zLMFc2Jrs5pvg2wXJ8Df/rQrLfhjlfBP9tOt1CYR2Ma17zyFoafh8AEcf4iJJIGTdH4HrjlOrL8Q64XJAlP77DqPbyWpz9gPd3fl5xMmsBtMhr7TTJmMMCY/OLI6Sa6x8rmGYFmk9eVeIQeSOAgX8xXeeKxckmd3bDkZxXfcAkRYAnCfMQdkKrkraoLoc1mIKEj//XG4cA1DD7wPeFDK/jRUT"
`endif