// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DIikyy71nTEi20MrzUZRmhwcTv78Am9rSGntH4I6spAQ3z04gyFpk+Xyo9VK
gn4MdxmP90HITizLoX65kkJVKXjqW12Bxns8ot8LbyptKji0Bwak3nbosNYj
N1o4Xuh6CVIshAG29uZzo9hM6TzC+xuGjAmcnTvGdWYZfoXnlINd+25Xt/gE
zrMek40+o8pCHAHhSHywYMmd6/SFnA2Cxxz6JO9RZ8upBG+DqbxnqUZ/qAil
KxYANeEci8F103o3oEMCQktfWIjDluZwjaGeRn0/fAfwxQVIVr6bKC7Oywqk
dMO7sYg7PNVtP0zf2zWUzs+WlNUgT0ueAuVf3pFBeQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oTTAx/ak8FT+fR0q+YLZI6GTjecwuhWgJMP5BsBddCWfLESRovpFRW4kgo9E
bKiItXuC19f/S5uK5cZs6g/Kc7URbqBFcIMpW/qFr+JjbK1wfEYvuuCe+Nm0
xJCq7ymaFaRzhIo1TphhDMkIU5xSQdx9k+GiH/CkBY/ba0UNJc08CHShCjl2
O69KCqUTdfG/Y14OnasCo8PaNq0XLDi5TsP0OVGQO2vnuonf0cnojAHGRTPz
fRFXgcl2nm1Uw+UbuknH4H828RGIWhKZpMxQlKA2b3XGRiDJvd3Uin9nJdMe
jB86bw4W5epMg+9wEzHbii0+8E74L1h8dFeXlapeQw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nofQgxQ6lIdwHF8gOqcqvsRg/ub8xg5urz1w7kLZSLAAqJonyFoV5CnGMtiL
u04C6fRmL1giSHmv2ZkMjhWZBrs0zehKZk3Lm6Zw+fvbHB4hYRg5W+FGLvvF
wCjg0Xv5A/kYJ2NcBxVd/DRdxDGB0LJ5Vtet+Mmre/t9DMmJ9WKMtrG5ZuzK
KflNpCJ41dJ9v8g6Fe+296vNqI6i9iMGr04ag9jn8GA3NAf49WeUl/6fdS06
jQIiyGZYC6/byVCWQ5LUaw6rM7vDaEli0WWDlBZpJ/0UAB0g8bEECWAZZY09
x206dbyl8gKU5OevsFlKl+pnVCtJqEyEslrj/Vo+qQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XtxzXAdoW9KIs1R/4/Ws8eBXrgO2HkCYKTCafGYFF6ltKn5BSMSfor2l3Ap1
gUNaeBdTk8dcQ1GMRdZh2osBZ7LXVmx15Qw2yvPtl7o8EQc3SkBzlXWNnmlW
5z0Lpy/2cHqSOOnoDo/3BiDWBryOMd94JaJwTYpydDu0LjQt7z4TsG1kM+wj
UENLc6RhjBOrWAdPhxjlWmWDHrCmpPli1v3PNN/TyqjYkZDoPxIGmL7cidJu
g4jMms8LOpFrj+op5p9rqAkyHFViQgN6wicluVPwCdGOx6QWogCsfrIm95uE
L+O9eVEO/BR2XlO/y2cXxk5UdGE0eOwwcMLv8d1UBg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RJhQw/H0C0Gs6BhRN69okNQgfQgn+qjLqR6rYt4RCONfhZiSfGR0z9vm3FT6
+l2zzk1Aubelxbz4ItFDcnnMXHmnumcxaS67lcVACVNDaJV5hDej6rrXEuER
bVqAykLpDqo/g8x1qxLkQGU5++9eImQTMABloFxAssjAein9q2s=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YLT3Ud28HRHYoVMA3+TBADAcVKi/J5TE+uw105pI3zg2AysWZ62ioHfexmZF
4A0iy6V5pMuTW0gtQ+ZZ8/pjNTEGEaj+n5U+eZ2QkM4TRvBJDnoBkek5Kimu
5vmrtz9yFUac/ZtLUggH7R2jt0j6q8A5KT9UDxbXH3ILKDu6EcEwFOpBDoug
/Owg0o90ieNkvahEvhv7KPrTiNw7G1PrlUo+1q/GybRB0ll+GndFpUTzh8jb
7pKMuwb+HFwLf9tlo0UEwo+bvel34TZ8QwhNHXCFhqWj/u4EFdxmOT+WJEiu
kdkY9FchoytWl6DQcvBudtrFanwaRdPZFWTX5mxhdwuHiVWV78E0V0LQULAe
/bdLDin/OUT25T9AjZRoNqSt/tUV7/RX25R4c0kctYGtWwo6peIADJGmZneO
A0G/61Y9GjZ0ZyyWzQjymatH6nqK7tiEQsvdCr0QCQeD1M5bz/yZ68ZvJaBD
GXrE42bue79D7Bm5osW0u1ECG4DftjU+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OSSTS9/qQ/jBZIDoqNt2Nw9nxQbOkUlFLxFs5/jQwkCBlRBpkiXKXgRxOsAn
ciVvTyIngRI7iIL4sxFJ8YmoVQ+DX920LkYXVjHzBUODUTrNCMyLdXsC2Cej
2SdOuyIVVLP1PI8mv9TA9MSJfrZ/kUDOiXVm906/OIyrUeP4tH8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uXDBk1v0Ldwu91M03OxzFvnoGsFoh0Cl0FigrK+gV5uwqbE7EmQIA77J7aLM
2P6OjeHWuaR7A87EGxO4F4q7y0RUTFwBBioR2dTnPpjZpaTm5Cn++BaV3swl
XWZ52KR0OfPIVp+aQA7Rj1feG4sWJj9Z5/IrbgzKAA2N/utOUOE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8480)
`pragma protect data_block
JZWfagl8wPh60rlsFNRljKQPJXeO9dcYDgbfdrs7o3B+S+3ML2jhAnW3NrdM
UNx6SsFK5lFp+2vjGftxY9VvvDWCVgl/jniu3MLTIsXEt4iMnDK9sxtWwqvL
L6MvLs5lohvjdi4/8KGW7u1BGN81LV74/AZVKPBnShSo887sEkUEmlaceEFB
bCsR7pb0xer1rvHpAhTP2abk+0IqUg6gd//MiPGM8Yd17RX3+RGFvuNxcFWw
pKaDOSaOBV8LlF1JYV6ThTkcH2g0X43hpjlFQemm7Xg3rZZejmDHolcAuQ9Q
RYxK+WkmgMEidl2BTFX1aROp5Yrzw4a51PPMs5AxajIvDWltaTot3Q/Q6/IH
PcOnObYsHm3ZWHcCf8dmVb57Fhb8lB1cyznS2bpBWwir8OZgVMHHHemfem/T
FynEnDvNKi2jmVFokiSzpVJL3qDmFui+fiOlkLdoNfhWtDIfsLdpeAXHDxtO
B/BJ8B0J+7UbK+SocmrEWKuUPrplDpiLKPwfbj7UJPOTIG2K1Vgaok8ayYYG
9VBYiS75ho1WNDoK9QUHxIS1Z98xrCjxjpLS2a06/drqNfR8kiKWj/8FzFsQ
DW7re9zssdJmRWoQCgoGXGAD9lmoI07j8KmThPCqlHDVWEQg3/rl2j93y3O5
w2xFu905RnZ0iIE/FY/WaeAEomcr/W6kRC8TbEqff5J2s4j9WlXlxLsOvrSr
HkyFcJf2abXKpaW9PwLqaZKTE114syjgjCbSS1nUJK9Z/eOgX9pL3y3AnY4F
b7jtsYjMnOU5jiOonIYQTWgnTagMOZRdbIthsCN4QOlm+W/VPC42wfp7zE1y
9NsOHFVMa2uRiSfJmdRm/ZdexQ0iE07q4wdBPtYSH0wTt9ZIJvJwXqvMu/ds
b9xN9Wv2Nk6Bpm462XFQiBbNrNade/BZJy3ns54Rme7qT9FBGILZ9AP6Uvtc
VIfDMzNh3VQxzdu/tq1ITgWYy7b6E+B0/codokd2iEmMXZ0d0a4s5NR2n3Mx
GKQVi5KpokAymrg0W/2gAs2W+ssi6xk8NLMnWTHu1P/I92dN/IOsk/R6Vt/O
GhF3np8J+qlFrCHfnaiUTY9ssOUtdEc0fIh4NdPSwnHsMNTyIKuKk/Xnw6Oo
O0A3bPHi13ECCmvQOnimYyF+ZRAA+h0W7Ahrzos9l/cH/opVPBpDdyOTTBiv
1eEsb+LfgVDukJLP74HcEpNxX8FLDn1upIPOBEqkMZaWSdzow19KElT5s/eL
GclHi21KM1kWYvQqxyKPkWLRFE43g1gmoKcV/JZW/RF2YdVd7bf4EYGqxrbl
aDl3/HCymkvDpaaU6ip8epxUwdMJN0f9pD6MLa916RO37ifThKpRA9ub09i+
VYoiW+AIZGBMhT289kvoYFkFE4Jx+uDzWChDQGgvfimE0cvJep9Hnb8xamxU
sX1Fv3Gl/Ry5xh6ZeN93A98Js1WYd3BfDcPLXKo5FjZy0EqiNxa/3C4D2t3a
uVb8YOS90bnBopznVtho0wLKPV0UsGM8by5SDRnTccrW2z/Zj8NktbeX7ppQ
PD4vNRRkJ1DWYlg+OWBk2/dhqvu3jtbfkGKwPaCdZemdVhZ+HgvZlI+wJ4Dx
0YJ28pWaigufvVqirkExLQOVJLFTVjCxrg7LEep/5kNOGJ1TDCGUkTtF++bF
i/SwMs67fPok3bJObsH7aDTLdWZf0PRJIoyl9NebmTCpZAxWrOxu/P19RVYK
KLl7N/H1t+wJ3I4TJWdPZq8vGzYJFDxgAa/u6HbYWFvop2dL+uPJ+97Jldir
PPf/S8g2op+5LwIW3u6d5gAeljel6Z0asFlalhEyFYoS26DvVa79ns+bs0n4
QF3uC8cTRt1ZIUU0z3owaCQsFstD1WOUP6JKE8kvx1i1gnAKMNp0ViHJqn7K
0okyu7diIyrfwLV6lhBdQEEduQYD/xTNfkFU4BRX1pLvfU42Io015hR6uPbO
Na1YEjgXrDZ9AVAOwBNfMYqLZ+RrnSo3PdIWqQEKRzpijYbhSzUU2LkbLl1Q
Lw+dcLKnmaOIOHijIM4h0nM+l+Fuk6REr+eor3inXV6nC5RucAstDXL8phVz
MmSq2h01c1w1Ao7Atkrck/u30a5ItPhww5sLywpg3aMNQkb84yZk7GPfH1/v
RUEhJ3ozeKP3kc4DPdhVzJcJrFo3rMiCOQzp0/GrvvwO+U+aSv6aM0wQ5+83
P610iYWzaHjHYGcwFuBOa2ttnktzh68Qqk4EzycbOVI+gqciWJWplVnwhdgZ
A26KIymHnyN2lnz0zPZygOW3P9CxMaQDby3jo56Tbk591425bJrGrO8wzu0J
uRX6xGA/G+BQnAdo38hS1lAc9XO9DNxiiRi/3x1GFp3uPeTlCN5VRwwngSoi
ELtuUcm9yFTmVjfPCczkvEhdmSZ4Xfde9Lm5LUXcvRTNt6RGO0maiGs1h06X
KPTo8oF7t92gddPXT8cg5Toz7IOSCOQTDROIHIm30cJ0fuE4MnXtB9lf5Is1
Kg7ZrIDCAF9Serlcjgvhz2uvJ/7jxkKxBQFaXyW3eiQL/4Aon0m5qHFrCgsU
uMfmdP3kiMiiPROlQoQ5oRjnC/dB4zr4Zq7FV+D3QCsKZ7kRpjiXW42s2zcN
85VxexuahYgeWLW2VGBjr5cBVfNrBrv4Ii5x0bHN2CkzQBvJS86rYhw+Hi4p
XmEksKm9eNGpquxe/yglFHB5RvZMBIlyaIgRypv2l5Zp2DKbdjBJMrdybq5L
2ey4loW4qEZ5rPS9q9EBdqqnxmrweGqMwV63zZ00rr56ovBFl3EGC4XRsuyX
qjkIr7nOoYmSA4Q6v/UfgVPbn4btggdGgugb/Z1kprXraH7CgHAxl7UjVHQw
dMYBNgLKrzpjKc9JxDP2NYSrHuYHUDKIVhTNAnFAEMqD1Qvr4pj668OwfWYQ
erJcTSIc+cKzDvCmdB1PeLw4v2wjt9Ry0Yj/VBbClCn7eV+Cpmf/sOIe7Cvo
+mjFVLAJNju246GhR1qc8TBSl/so1/FXfrqiCyitfdl8g975JrARnP2tn4fu
tthqiUzITtZTNgUnFEzyDHZXDGkl3kPN6/1kBZZ6xSKOYCnQdqLANJaIzVhE
uhj4Uz/ujPFrcc+aIiuwNgNTBZsAJjBK4hpj4LBrlAkHsKEkROLTOzYaYyT5
m0eLenlkOGpzHjKHcXD5NFlqY6uYKRBHKbWz4By5hzwl3exuPzfRF5TBOWFm
V5kHG5b9azy366dR9+F2BiyMb1RgCJe/Wy6ER1U34lUm1UEcJ2a8L6NAVp16
9Zp018GOJ23L5t1SxsHHH+KvWstKUfRI2aNKK0ODN3nk/ECdqkCUOzdQKRcV
QysW5kLtEr/ALycWYgNBeiOn70Fu9mukyr4xJrW7LgYCsA6Hp+FqAPcjRVzU
AIFasbV3L3Q66uV1R+tM+xizjj0xLkDj5C2U+BXx96O33KJwcSZVZoefIjAB
7PFUElHQQMk5EJuthcH9t9t18DHI/qLtfzwf9BvVcRpd1/089CfabaaG0/a4
yKaZIe53EWOmaahK/XnBmIeW9K4TRTDFaZRmSHS4luoWIdwcyvxCyFfYSjOX
/htqD+EAoYeXmhtpxbFjp7sruqUUeB5wY4WHpMJOyLzh2FxKdrA7tGQO5hxD
bbd8Gly12I+tPXV/fZhMDvIvlxPxJE5g3R97t36bExUFIK81HQTY2JvIMNHO
29+GWLpOjc3ACy6mUv0r8s5gYmVrDSCRaKX2BIrXFG5HsvGlIxi13RqTvEe7
pCw89Zho7+2L4I3ZomSGeLFlBIhaML7DGuTMih8Ij1Lzx1P41SOispcQLxKC
IoShFLbwJ2isBoc1qVduDZObq24Ghl36CpAJfA6rEXhnn+yQpUse6v7zTRut
OryK6An+9dKDepq63QF9QHatXGcVCR3cqP0Fm4cGVhQ9gEzPXjRbl5KvFx+m
WDMdf8q3ss9vtex1nHFVht7am+EvPFPZ/lusdUWJ+KYUpeHBDvj+rnJb103O
phSccI/QFyD7Vc6ngDfo4bZYiAkJaXf7ZGOELg+ZvhB1dkegxu17D4F9qJ+Z
akURTD6bHXk4dn8rr18NBU6bwqVVCJF09JJDmB16QNQ3+QsxaCeoZg7i/blV
C1pRYefLBNbWmalCURVEmIxI64HSSPVyrPsE+YIDxJsPo8Koa5vHspI1lFvj
6zcZoE0UnyvkVLxP9eHFgMsv96TNVgZHgaXNf+JRK+DSNk/iqyB4Km+Chy1I
zEtgaDCADp4BXx2Nktd7bO30wykUAwJw1dZyAZ83fATn7AxtB6khg6VUcmEy
gyQrSUceOWQhyDL32xTozUaHWKaied8b2BFtdVVfluVajQwg+mOW7wjUjYdS
hBOwPh8X9r50IV9mF3VED3JFJ3z2H1/a+krUW9khgLQ0Fpa0m1QehRCceM3e
NButiKWtq/okZLecylM2e8j9MYiKOAqYN85XCozxaiCEq31b+YCi2teTg2bS
K288w9LcNxZvi+afxRrniiEJM6bvjaqynedf7PL4Jl4akzGYww1Oj//33qW1
TAzhLCT3x4SMjspOS31/xkka4/wDmiBvuUcwOaDgofLv49eOfTY4q7yGNBqj
3fsrcUi0o3v7/sspefj1KKJKLm/EwhHitn84aME39trFejfWDwy6Mi8Jf3Y9
RD1Iu9lb+wlVQd1pZY7ucftLcJlW1DXkEvmQg+to6LuLybkc3zGF4jIgy6TU
m9LUheSGiELuEbiCHNkAxtwLcUXIeomvLWM/Z7gQVJFQ6st6XfrylZI6dNqS
cRhdXgNmqyLuMATEOreyx03ZrGH9boREFE89M4Uw98lKvqkZXQtVltToXUao
t6ROQjnb26fpPQNmtowZA8xq6zHQ++LQm5ZnPNULU7oCrYjSlPYsEbK6RVzA
Ut8UnyxFwqRocaQI3hwXfN3In1BSWEiI53smgwP23uO8I/PDM7V1r1UuS2B0
kQplNLfWIU/AqFwZhliH2f98RcgAqWuub1EtLjtrh4i9Uw9kOBDOt+oVGugk
wOYS7ThvYtC5ZcA2JPSnuhGzboPgCjxMqKi7haN38D70w4xV9oIetVj4xWc2
ZxwHpvxVj58YYu8PQrEWp+QSRXi5AQlVedjPokHgqWKNwRhjYuD9usWN1Wd6
T64nnq1T2O6ZhWNOv9H//PWjvqfE24N+6J3c22AsEiyzsZ/2o9++K2pRbZ6M
NX8VDYClL/T1nsgBR0twjT5drzG2zXf7RKgSHT9/2B+xYd4vmempOE7z7q2q
JMfM1ij5VN4lHlKSAOQA6DshCjpv+JlfmwlB/8lHuPmAOEyw0Kwt6EtcyA2U
OANq79cDk9xw3vArWTeF5fksIWeUR0CrnzYIo7w/rUie4SojaV1tfB/cxtE2
14GDlyAuA3teJVMeciK/EsxjO+yV8qf4LLWiSFyzsp8OkcpdTTRqmqu39zJ7
QOeXvqFUBFQmrNHOByunpHU307X+ZSg2xP1/kySu3mq2+2tn0Co4oIhEiCpc
HM5pL/f7iCWEtd/MlTfLC9mv1J3abyd8j3gOihmT3gtl07lWqlt2oo2cY1Oe
x9KqdUQ7lyoYb5UGUNto2fd0sR7pW4+lsTR7Mv7DeLR5z2Vqe3KXmNP1x32r
ZbH7czFMx+XISY9bisNFONzD5tBWemwiMmCBom6q9diFnL98e3baYj5A7Zen
xdlIikcb/bgux8jAI/SrLSH28zXSpU1t35ockfq4fiWDNrB3Rp2QJZ1NBICK
LMwgqOzDEvhwIuX3nXScXOiRiyN1Dl9/HpOA64lwV8VZU6Ke+hbVo4iql8i8
l4wVp665hw/XtoekNaBb2uUmO7hE9Bx3h0t0QpIv7P1ZGE+b8cQxjya1aT3G
5Bot5yAlFFnXwW8KZTAJ3xY07wSbezz7rFseqpzEC8gSs69reuJ5QpPW6XRc
MHfK7iRhkRXNcIMnvMaqz+LTFyWMqTFLIvFE+2Ohq0kQYBrfTBl+R/a8DlF4
WNs3RodXiuebXVEBmbNGXTerciL/vbUdYb2zJBQC1OWWrJJ9rngkr8sum6Gn
B7xSRAaf6Sl2yxQ+kX6XNWugI/OF3VE5R5Q8JLrMn1o4tAv1J2FAOWfbVvDi
2oMtsydar+ZDOZdEsJ2liKbk1TJmafbtqZCxKQUvAV8GNsSbD7aPnH/Yokpy
QV2lDlIR39+QaaWZS3VaZvaqzcGUEo4ovSupR0lF6ZmjD96oKmIC+8M80nsk
Rt5uCqU/g3h6GDcmBpumVpuwriZ63PpXHXLzdMefS/7OxIVHUz/u8mqiTNbp
xucrriv8A9HtHKugy7XifkLWJhlCZtEovTMBp8+UJ68QVY3sda5TcX05xRPN
ZsHsU/VapEpl522uyqC8C3QLEEfUZRjHuh8JWzQcGeEMYmi50XFtIi1tu5DC
MIu45mWIWDzG5w/ARSPGS6uwuWsr0qqe5Fh8tJXIZ42R0CA2h6Hjte5R8CS/
ci69W0UvNwtAEQkOupC+T8TTc8VHi5XvyCciTx7I69Pt43Wb2hp28Nn/SdRn
8P1/NV44IeTMrQuRIf45kgbfB7MuiclQYJ8xNwKeraxouDtft/e9Fja2kKqF
DKBZNspVhOYS+IeK2B7CVVfcj3J4WKjoGSQN176yStdhdDbGj1tr6YFuxwqM
6Sw+m16UKh2jA1mdS3EJgtMWPm8kn7EKPQULpzuc1mreJMphK6TKsINtIaEJ
cIfS89ZVFHl9MEUCeJOc+qdkPOd6ptrH5Re4CKPqElvJtlVHwAxwU5MT4vYk
AO1Z4lLc6BHpzbicrTF7kYZM7aJ9Wc6V1fdT1NGpSu+GV7sSEKKCXqKxz4NT
XmOIap4dzOJwxhymxNMR7IoFldYyjmdk/knW8A79t6enx5zjokZG+fTmbIy+
zUfZZkltmxuEUkkuj0kjdSIfnObt770e7YS8GPO/buPb3XYZHbsKMkwSV6GR
ICgCJERrDAypebHQAd09UW1nWrcXJlZAiaJ71OADd825loB/NYQnZjn/6iHZ
t5sMfexqzNkSAQhVGgo2LWCrH8IshhJAWNCMBPXrWVkALshx2GUvUlkPEZAw
R2MwgPS6WEIzQl/jy+mXPjmXt8fOGKd2ZvAY8cc5G5MaZFuTmaRhPZfk9oeK
i0Ile5D4MTSHwunQpO0HQP+f/OE5NnsBWhfrT8ViRti2AZb+RC1jWyeA+nLw
TloZ2jM+fd9WOFfXKMW0ynYICaxYSAwRFarx3CxOhmg6hJj7/lRWUGiLPl2K
8toEYHaTrgAzYJjK12LAkYp7BkqZ/ye1ZT2Ojex3rH69fyhT0pydsQyi7UBc
NlwMewVNdVZYakp/mxFvP7rJAUrpZe0w5SUFeHfw7jBgZKTDrrE/A1ftfXWa
cuUZxyl258agIQhDMycX5a3ENO9VKw9Sw3lmEKdVyGOF1yR0pC1/rUhic0B8
Bvcb87l4uN+3QL64F7Cu9rAvvYFfyMxzTqGeNm4o/9YPIu+38+Dzci3GgpwI
sFaX/ZDDbwvKqDaraHSh3NEepq+v2v+gFoEUB3Wa+YjWwDw8ushuZdIFiOd2
/gvPZ5u7pvvXuxYoErLMAf+k1YfL61cKSXnxzR1SgaFv/OKDjtbhcasqzuTv
DVfrZVytFkp3w1+8gMorJFweAx92tzShBcvtLftds/FU1I4yYiAweubaAaP5
O8NM2YvktsuFX1mVZFXEkMVRNknvjK4VJlCdwJlgBuda02XWoDNQgzwGdZw/
TRA3yeURnXr8XQjsG3f43A2VRmNQoPuFPjiSxKC4mMoP069Mdu6AJEIa9Ya8
nCzjBTqoYzqLfntCmYOm/ml+OCehn+GzYZAHO+Kk11yN8hIgFjeYyL6vLUcQ
bRZBGrwoV838LEJ9H41bQN7UYN7Sy0oTeDquYkqrXOWdAQcR3pKBb1dd/Tgv
QWwoasEDfGeoxua6Jv7AWImYAMkTEeaP2tINtOokiyUUERmaAxmYcZRrkOgi
voLkCf/+v575dN6zkObSFDo94zHkiMfbuzLoDGGagK01ZzeILT6CcB6mz4M/
j/iJb65ah5VBtbrcmM21so0hwGVLjU1dos5wigaaXVJYeE93DBzWy8/6dPs3
8mUqRkNrhM3Uthaq202svuTIIwfx0eGHMfpNdQNF2h8x6mzVitP6t1GE0mqR
gHJY25eCadGNQW+6kry+Asis4ki1dq122OO76ouMV5i+UFMDi4PtSFuiXKUR
CVEwEkamsiXEzsyxbWsG/Ij58VGHfEQ+n1yNhMVKZQ1nOtzw1krvgxrSwRU5
dP5f/hu45HOjUghZXqaeRLVpOZx/3tddrIVpFblJkkOuMhKhFIR77Fs3HdmZ
0DnrGSRXgsEDXi974ASibQfA6ahvi8X7rNSVaFusgPuZ+c2MhBpIYAjp/WZc
SR5aSsH+zk3erg8hpbm1iTlt0DIHXJMy3qssWUBO09kDseQ94WF6kxk8a+eA
Nre3OyDeKU4OP4+qKPIMSV9Zfh4IL57mf5hfeL28d8akpZNIlO0AKcRMBBYK
3D0vB5KOR2xof4n5Gj1eocVV9/isowWCLZEP+QTWbojFj6i2Ay4Qp/7xPdH+
lfLRwOmOn7JMpLhtrimork1LJ9++w+r700/DtiBEswDWbMtINgwTQ4DiaHLf
W26yVrk4vHxjKtxkEfduJAD0B7BUUXKFyxd5UpvxBzsmWpNg/Z0F8Nk3yGnl
xMOy/SCOhyMlLONcVxjrki/lhwsJj8u5ffwdCdEoRL7qdahPa/rouZAsXeg2
wxq9qOO5jZiNX6C7oSme16Crci+U1ra7KA42IEOizjKOdjLAvW+RtiHchOl+
TTT7hmAoPFz3JUHwQ3stI2i5CxdGX1EBiTnamYGS476DnGIPln2Px4BuVvRx
GzJ+8bl724vyVGIDt7sGbCF3wYMAjEVNsQECQMEhnPzyFTRTzdLd7s3P3MhA
W2cQLaVkLzT48QspzF0PrGAPjcVgHXfTpIdpjHUr6BpXWAqTH7az8YF8Vbq8
9JJy3C6VLdMjleaE8orE7b/LwbDrXA/kOA9IeIF5UssVIuwFez8rq2TCntEi
0bMZID23SygMld1Mqm9bmIG/BaYbF1tYrzD0uJgnKVMXK0x1sp+wwwE0ioYH
CB7/NbV7tP1K18KQybe5F7jEfjjO7LdGVysrhBaxA4kedti6xWYdepj4sLTa
0siyu4puu3TxwgkJRYxK/DV+oLp5bjEBXSGv7TsNiMh3diNWgWFX0QnjJTMw
UJUVNJk0d1oOkvajuCLwXMfSMihip2vd6TKreQPMLyp6i+sBbfnU8Ik3ttS2
0/J0tfkff9GWpWQMymuDU0hr3wUw1/9VAshB0mQ50B7mt1qt10bWrv3Tk3MD
eRx1+6cYJO323VR9oPGtgfra1wAVfqSwZ7MhOoX9pjqbVTtOMzezmOrV7hIV
OqV8DBu0EAzgAlU9gl7em/dyAZqg4hV/3MM769CIqY244kMC/E6SoZz6ar8t
2Y19QC62Qe505blAP8T6YbXl0GAhqEVI74ZYPSMc4WQWWqxorAXxA6pQp4Ma
g1wL2Yq95BxcqN0otGfXoaGUDtPvAaEAVjY4zfvi/ODtNXmj0ZSBvrW5wCZO
zuavSCpm8MvN4P432BsU+Ogyz/mI0HAPkxJjvDNVs7OfF4ODe9mvlVZxSESp
7BC6JZU0Iy+GqQLcOv5TXc1BUFYT/3LuaHt6SsI1w4wvrAA/zi8zMWJhHzGh
+le/0rtChJz4aH4cz4nl1s5l1TxnDvnHMQi+X1v/n2430vTbZLjkUKaDbYxI
g4xc256Ie3275g+Sy5CSVuIbmVugpivLDTPdt7QB27Dh+yVpWOfrv4Ytytze
Bi3xAUI6nwuJQsotViODb9b2tP6njbij5jewudxJjcFYdjBYlhkkAWYUKfJG
0UkdyiaJe5CamkTfdotHiq4ZFYuLqTzTBYdE/Kp9N7o2DnVBp8ExJykeEtSH
hLU/hWloHF1itX9ifdN7mDh+F9OMVPHZfW2v5YVCMhos+Zx1l5zZLO6ID6Xk
EynZoayIrP2n56QNHFK6kaq7H9c7erytX7byIyrCMrCeIFCAsEhUkYIdeB1U
drCGeBK0e6v5t+RD68JRjQmB9hCjFXWlY2fqWiFwUS3hBmbGYSifnDqtrA7s
wOPOROn6aPEEjFOImd+dUOnQ4u72kIF7XxYfFckkEHtYRvcWU4AVltZ6QwVf
M8cYhyexQcKN41lWHInCQBK295/nYmiks+S9uCwYTi5gdgX/Q8v43h+SK66P
gO+RTY8FXK9cxuZl1N2AGL1sonQuN059oxPKyAP0SvRkwh136pn0lx+htfXF
hqle95k7YXLPMX/nWXC+03yKaMQ3EjF4q0aosyIdN5G5+Z8tTq5iekhq0BPu
egfywVfFZI3phhOzD4rfjLnFFUPWDyrb4dSnpmG5gafDGe8GvffAzJm+97Z2
B7mGutZ5u7xFtwBm2tQFSLk3XF/KTSkl//yumceeSNJRbJavzDob21aA/M5r
4HzcjLJAy259Jn4Uqh+E14ifKwYZxWYGlEe8KMbmQqSrF//+pcrFjrWBl9Wp
t+mrAncRt1UHAHMF89w/MfjmDacTIG8W7E76X39FTvSPXKP0cYAwFI7hyt5U
0ZNLeGNzTFIOcJzxU1J98hdHnksg4ZPSe2rTEb8LhUaS8eYpZFwJZZbid2l7
Iua/jcbJind4MEhbAXlT2LlLH77fNVmBfB0d2vbfyMhTrF9KBj2lRErYhTAk
L60pnZyclEjaokVncywbrZwvk0GeXJ12ojo9ZOIJWeGBAf/GqB+DI9D4C19c
BojdqZEHv3kpliK/W9XQlBVMyEhP6v3366HEoUKiwlgh2lHhKypByS0/M90E
run+vJ9cqWmCVRNEOLmUHrjvv9V2Oj0W1v4PHLtSd5uyiyeg2jHoqzE3TCsm
yvSnv5wj9qFkSZKE1VzWrR1brTjclHph70mW93HvuJnnpMKnxOAgaFW+zyAQ
8zK1dQdSAT9lHidkGHSGQsvgTNlIU3B01+1lA9FwlePueT+y/uHSLT1Con69
fQss4YgNFaN4ewQHZb6rvBmU32EbxWdokciKXQEW6O1BEQzXdR5AAYpN4iOn
pjDi6nxqXmKLN0IiQnaKAs9NTM8Xg+L08he6JqLKLMwIHQmg36L/S/a69Ecx
fhlG7gwUqq1E/PNAEw3On0qgsJ/hX+yLZgQ8q+df/ofezi+aMLVjyxZbrq8J
96OOb3mHHoZAS5IacIWGTOwr/vcoI0TTHTXtd2RCgKUFnkmK4bVZQpABnEyE
Ms6ujBIKGoqwfowEO0qihYkZd8c=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Kc9w7Y47B6jV1QbgnMUl/sq+eBW7uCmd65LZtWmnGyB87iDj1tQVmvgZqJeOWP9vhzWhKuQV199rKFyG/TDRWQZzu53KFh14ffvaraS0MlnW4GpOC6d5JCkfZn9XO5UuMoWUJvv6tTEs8vkEhRmKyWjDbmO4S3RE5oxMPYN2LGW5Sh+pbCSs91ZoRpfPyDn4JKRjm3/T+K5hfTHrA4G+lv4zMkWfWroeXjoyMbaHFzN9AqpRSlKkEoKflDoNPqlbBZZ5+2YWSxM83uao12CmImCQe4Lblz1YZW+5KpwrWiGKmY0a2j3017sLpuj+QRjIx6v6MV5fUF22iI1RIgEd+leBTiDfH9lPi06878Uyd6PMiuUxVGCW16Iz/sV/NmwLcTWr7ksOJggvapDtKkBstVVjgUhCym4V9LE+K8bgHMrJYTgOmd01mHI3cJzUuqS2R8avFJshbxpoTU6x2F7wvy3eim6doDvzdjmW8iYy2wR+g+d6fsAVU2ZZ67vMRDLETe8wh/BV2o4V12H9Z5/VOuuQnkN8mvGPke1NDa3TFFYGOCvyFH5FRqXAC63cNSKdTcUTj8DJ5YRPZ82AaSpsCG5+O0LP2MsJh94P6wB/Wj5bWGkCL1N/YyqunzsjvfEfjcE4Sf45n5+8chWFPSalOpfsNFdgsxFubvRzqpAuNwuIWLhSOvP0l57/+hav+RgM24swRSGoAaSBjuWz4wqnZP/6mu84hGVUNExFwS81TILJmzWlL7521jPQLJtz/uN0G+jrOlMhJ+54ZJMLG0D+dr"
`endif