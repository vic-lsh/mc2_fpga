// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tv2DnPz808LCWwjpoCKsGv42GRhzSXT0IoWyaEZL8P0kALhoTg/yPLXluT6Q
8rW9Jq2p9fG3c7gbgfCwmxHUXDVmmgFI19mM7oh/G0uOtwTvLrY/2dvF3I27
Sj1f6ieD4bAJhuTvpiBbXSEfMtI9kJ9NAnziSHttzuReb1kB4p4a8v2rlB6E
bxJlt90uH/CeR3sdgxNkO+B/sxevnfiK+fX+KL0u6QRQE19rCqrDJVJsas+8
CRk7uAiyK5xlDDmN0IAgFPzVmsBIhSONBn4FucrS9+NfNiC+VLECE9+ZRcKN
OQMRTdZaK/aGucEW1ls21Utj9a5sj6EOKBRXz+WamA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k1KhNkgoLbYSXdYyshPcYkW29+MkXsZ/uG4zlcY+jnghbOLwP3Gx96j+O6Jx
LPQEi7tXAweozKGClHcJI50P97jzVNESXWcWqaMSHkhuyaGr1ombVHG9Tcsd
y5/62F0VqajErvrYsCPMDkvV/pMww+eqSJVnsFl/r0GJzUMbEyj9q4kq5ckd
87E/D/M8cN138DphjQ8q/yUiqGZXnLW+vym+soRF46uSq2OAY33g49Bm5P/C
9O1sBbuHK4hiWar52S8f7aQFAktIvOx941RkmFsODYNSTD6ueqxRiJA9/isI
vteeOOOVmr1HFhytV1aIBVacDl8UHeMM9ShpuJE36g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t8EOkjxTvGeSk77JlRNsSYdgNACLnTRMKV02QDOYruwhkY9qVQW59jpYAGgF
qsOX1Oi+danyyUfXBanrWLBv2VtCZnnLxBfvsvNAu2Ini0DIq+1TKihofKqa
sl+mZ/Q1irc7LjZpAZM8iypVM8L3XrTXY6wBIEfkwbbqHmjaaCah/lVonxZ7
FUgXZPiT+yCK6DLuxU5MaDVtcZ5fL4yJ+cYe3duAVlmErbWo4Rwm8fgTomfK
w9vJBo0ph5n7fU3bw/9hr5ekYuQ06oyzxJxr2J49iKAuzWod8hOTz6qO2enT
vqW7OsdqZ3MzL7RugP414KWUCUGT54Y1FSYbdJhc2A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jh6BkJlhOtBAw4XI61KIgXC8L/blXBqFwmgO1oGnu84ZZpBE5ZgQUbjRLXuB
Xk4deOvQoAZ78pBmfbBCHW3YxBTwRpHccKs5huCS2reuA6tnC29qMPk1AhUx
/xiNx9swQNjg8pj/L3Kd5REpjfKcofA6s/jxlbwk+MjBG6WhL8dN4+8iOAWX
OR4acfYzmT8Rgruwo2CsCDcWb7TFZBq8FeN6BgOS927SIlIzrnL6c/S2dHsh
9U3tvOAFuOA01WDX0tQUyImwuC6ryd4qGBYea3sMKZ4l+3E9pTGdIjFgJpKd
l+Shs6Wc8V1gaxPTlKzo1aPdb2EZQfZtzxQM5zuRdw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sefxSA+al1aeak7hQMWHbT97ra7fC90G1bW+C7/hNtDSNjWB9OMrBrZsz8V+
05iQr5rPJTKo3cGkpFBqwL86pWZCXLQa8ELcLKgGpr2M36X3emD9DwDgXXw8
Izj2LRc8M2IoqQdOJVtOTOVgHFycQxlCi/UB1JwR5e7H3lADRHY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PUDO8nnBddfyq9nUMk5fHA8ExTO6rLcXZrGHNclhQ0L7QIhpku+yRikJCKkD
DUocE2W5knZjIs1G03cyVsGEJVwwLl0DB52dSv8415cVGZ7M85ZE9LZsK0dj
dKMy2C3QeM8dvWjMCHGE89gdI5FaoXAJxeoaM2JVDamZ5M1ptTZzafxAHjzV
+otkDVOab0TywXfgHsn/bjOsKtY2ZuJY7e5UWArMsECmksALvUCEzRocKlNZ
sgONO6FsdQYk6uaZ4nD7umHxUMyaJQHvPYD86sAo7PhtH6pjb+8T38OcjCcn
i7Er2ZWvG4K+d6pT4zCOeODVdIj2GAk7HhhdXDttuCAAKccF6OKBnf1LC940
RHcwtI7JJckpF8/CqP8b3JOHzCWCsntYXHYA6qy+G8cXRgbDF6quKqbWQ+jn
1xW2PfyPB/rvdePTKsfJAWVfbwkS5/5PkcKyW+2eNCafE3QLoMZE6RsZfLRa
WjReGwxAiciQ6BncKOq6DG17mL6bV91V


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tSKEEJTGuLzC0aUZqnDQ2VQBWnTDfo0ISRE05SBXNrC9BGd2aRHKjAmtuqGD
LBhJpoCMDw6kdK2QSB3N8SREgl/St1ZXHCvpanxbEydnG6k5C9MGCE0+pC3X
M+MFhRNBf7cV6NT3bRHzy3h4UcB9Dtftr8pGLvn8vu4L2gnfcGA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qO6xCiUgeuhmNVJwsaIEX20BjjigEGtrchp89TRjORJDBXBUAB8YRQyvo+07
/z5CtwFdiFJshgwPHTFj8Kk2J++1hdKxkyt/JnjTrnX3mHQ4TgIp1YpJDx3K
mFhfTk9w0QLPqmgbqQ5OORjaUotF3llFrhfkBG+MLj5HsrCNTk8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27536)
`pragma protect data_block
P02/U78dVVMgZtZ4G9fmsGz4chFyhQ8QN+67Jzv++iuUZ2IeHJS6If3jDY+M
hCT56zOIGXU4UJqtZaDg1JlEpikwRP4IF6qwyDLZmeBs1qyVB6k6InVoChuh
x2SohU2y1qO383hg2jMlN4ZAC4lHsdHiCU/Dvc4a7QBSgNBGtnT/KmRyZV+C
zvo1xik5/imQNCNWPpG71lzsO6/94vI92iEfSSYCUijvU4umkHPt3P0VeQkQ
LQ2JR3SjMXvP94p3z9hKnXIjH9MkSs44UdnBR389IjM1X19IhTEf6jItwiQi
JQXFN+Mr9pl91iunOQBI/Cgdbq15xcyP/HjwOIaAqTORZoGibOVEqWe+VWrC
IVd/L/0naKhwGsxGq+pQlNjCTCwJ9vgNOa+ZZamIN40SxYWVSbukWMqYX+DD
8atwYQovOd36Q7OW12FQe8bMjwvbSKtgPEA1aD05NBPD/Onvj6hTNw+uF5UF
LaL1cIG1ohvhpAc30tirAjgIvLvDEslz2JvN2T4+UIikRB5sYv/w0fJi2wZq
BewCNCvSHZ1m6JSKMwxW4DaRVJj/pD8p8xkVlN7Vz3DW0Xl0uzcyNHVGLO1P
CipuufA05qZ/VkSbooC5YxxSDudWJ3/pzEXEOrHJdaYI1LAF2nVIph+1uYOG
nFsB73nlTuwnzKe0rnCwkOmPqOWapmoRHhpUiDLSnRatAWS0JFQDae4zUKD/
1M/J2Z0NWB6fdVtjl/Ve4mvfQYNyH24hfvroERWAICaAXv5cJOG99PZY9cFX
jGW1KUONCFUuJHd4wGf/tFjf1Lptlk1zzNDWyHezb9XolWseBVA8EvOpD6PG
gcdTJxOQzJQwu0BR6xMijtqIaT5uahAP2cxZg45hbZRm86vttsZEmXnyGV13
mvUgLygZprCHYDE7WyEFP74y++3B7UG4uHkNwzNPWIO6uL1xnv27/37vSaBS
6HDXttxOn8szBszFFoLHIVHByOkXpc8BJSdT36HsVmfNjjOHtVufMqbyGc7D
8u7t/K1QTxmwdiMsLvbZ4E8z9f6UkzWmvFd1uoxzwxRtqOiuAWwgO+KBTzSm
9ptket/Wm0Rd2C4WKrkHdMLyq09BAPfIXiqHPEsQZv1mrCv5W/fADqIdHVkC
URshZcZwYNZvDNXRezfAHYrp7uBun501S0OCxUz3x4tLc0fgpb6krdFdvPhP
3vDDe3dXu7fjCaJowN0aQMhOdQo8yrUrh1muIMXB7MddZOJ8V7va9/0CSe8K
AqNwxaBBVVMpoT+apAb6R/4gr3m9ntEmLdAqofmhPCGqeboO6DaohMtDzeh/
Q+Tlkfa9BTOuPzkn6oEIHlJuzflQVsH9j8kejp0NHSl8aHwk0gyAfUqRwIcw
J1VaXlD6EAbt4Qba8scPg2DwwSGJPWRbNzBeXHzk+ynhL87qk2/gkks7dNW6
SRm2v+OqFJUG8YxbokjKadmefeyMPBBykgvqJ/KyC6GzLOp8xr5IQ1nM+GeX
0f8u1NTm6CVzSjtc6Tf2vECJUOWic6ScSQi/IPnvCn1VcJYkYtooNwh77QsG
0h5xfZsA+MJlhne/kurdV1gjCrluJ3VhrSUX/dew2kGfVlHYcX4WuNHvApBZ
elwjdomjaJXkbpdO8Zawe0MleR2Wzj0EQG8Z+iYRYZ0yXLjSKNf7SG42eUV7
Q3uGhrCwGSLLxtthhx6luBE+0nPa1b3ktm1/avMTl3DaLxCvd5GxpE0qR6Qw
AGQKcsDtEiI7zjY35b15UHaoNTWW1VwJOclsB02S7yfTy0qdacbbnBbh/Izw
M604n/Eteu1v13ZC9+8I8MPIMdM1XdSQf6pCZCL2pXm944JjGE0lWJVJMC8I
4XUPD4q0C411Zc1OBhR3C8HrSW9Flb9CQ5Baky2qfKntZtZbOboKNduANyRf
BjKRVj21i8KJgMwHBH47O4+wkiaYyxKr+45dfWc6+MlWL2+0/0Pwp1Tr3a8E
8NQn0w7PazbVfHOIWdSvC6DmG8hCaIRTH7wpaeWWBj4cBaHr4/+rYsY2bQS5
RW1gf/GGqQdTYZoixgdkFklZrHofg38k3t2zaGiOWeXnziRpaogbtBQhCoYj
YgTk8mLaCC+xybNQpp8nFdf8vhv80npEnxDYrnvqYRSFsnFV4+lk1O8rQ6dY
CF60hkffg3NWPRnbXlA93xjTrle6zEgVVVl8Y0z2hJoCyTEOR1gEeEHjwHE3
MapdcBJip27kFQ+RSjU1lnOGD12O25/boblfIlLZZN4FTevn5Ecd0KJmJrhv
N8y4Zxnao0ip4E54WrMKHoneimCuzgt+oPDlNbiThrSLZMbsFUK3VV8KNmez
MqTbKC1IUBRjXgYPawtRVT+ydJ7i+k0n+SV8AI0s23MUawTz1w/mX5vAMljm
dETeXZKEMJsbcxQ/ZYBmthzriF15NqgctoO2elc8ZdrJP38TUSi2q7wQ0nOP
xYveI0w8CkXxg1Zjalp12TjUUoS2JCMegOh+Jo7swrEz76fCOPM623ybHZAG
0bAL9/tMKyOqUofWUawYCwENoTJLL4d3O5k7+by99IZqLVZ5pC181Ew3ZrB+
c9cbDW4MeYpWrthewH65NPymxBeabSv56KxxmjDU7pAfKlmSZ6weqUB4O4bD
MWSBc7kpId+gabvNZT3XXRABe1grJFLgZ6AdLojLK9sNnsB1DDQh8m64srjU
DxM7a27PgtWciIWLuQR2nMS8L/jC/gcMde7jOwaPlTR6lA51YmM/8fem0jPs
rDKHMVX0lDflBVGzDLTyJI2Y3PgdfKBX8KpW3GAWHVrnidLDb0A/d1Bv4jZ1
wqEnNfuxlJvIEv61q07nJHfjbJSgZhF7QQvSLarUc942FRg06WCAARWBleAv
6FzkvYUuCx/tAF3p2dG8meLxQRfdjNax6bBhKH/bx8ycZQbCoQOx0hVThx0S
FUdXWGOXnWApeStF3EAeN5n/aMoEq/IVbZbqiJfIPTutM2jCfvLnQBqpmy7o
8JebENDyUbSmdEOYBohg9tSYuIdclTG6YiHUJjGwN0iHP7fu4SLy1Cy9dJGJ
zJNjDVSQ2jfeJsml0Kc+6zhpus2/ZT9mTYfdwveJh1iBDj2MVO7p7asG+0dH
JPoXvC8Xb71FtmpfktJFUxNJXXZr7i6RCZ8QT4D0VBQvdkwRw1KOZkkxFsHz
pk0Hy3rOygUdrrvtxPcEN7RP5drdFYinlCfVCIhDcJ9z9HYjmH0VB5bVn5qr
4VdCMedL6+33a2D+a9bJWiFi+/Izx3D01YLImubzjrF775rYiPr0X/Buk7pG
eGA/pLPUiivSxlh8WP1i953xG7aTFsutWkR/RiqB9YNgLPLjw44x7PL8zyQT
2Epvmf4PO98fezMKEV9eScK2rg+xQOYG9bDI7+x4TmULFixrGP8BGARW1j8j
CBeeRcA5LNGefoXWDZz+bFwXZIgt5uG5Fzu7uqGZIz5T+PxeAY8HfVSu7u1h
1HCLXE4/cF5cLiPgHJ9aP42nyifsYarqz4+9mcZokpYf6BVq4flfiu7wgued
eo56Mfdl1ZV6s6eHgDQlswTPM2vOowXLxxfHGkbNc9QUeqrVEtC1Mt7f9M7K
IHaXM2YTzoYmajoFD2OWASaQbaj4OLD1u6zrjExAUyFDLlqyN1aw6kFQBRE2
Oe4vGQLmERCWh+idRS9S6P2sSo1ZJXCdFsVqnOgK7+4JVLQ8bPJbMenn0FfI
BJAZKZIaXrceLA9FPawF4SFBTH/eUvDE/ttFIv/LQTjlTB/kEkfLQDVyRhl2
GIXT8+GPZhSwWiYBbTfexlQRZlMumKnaNypT4bJzxaCns1MGh7E5fcu/lVff
Db92FUGiClTwTACU1FHRO0MpRUDWtTpRyCvew86aZfniaGAkuU3oGtQ3/hEu
fxxESToFfLlAMiYG41FPupfOejvujMjrqTK3WC9uCMGvfd5hirQhzuABZWRZ
6lO86ybhw9io2uTVEPlTBsrnbMCUZ9Y6w0z9aVOEijiDaKEUbKAanf4TEIau
ap/3F5pZkTDnVAs7Jb9Ax7zMezBIgkC0Dgd021Dbmq8r+v81a2yzTFCdn2ta
Pud3hZF5XgdutH1+5WGhuwrd4zQUQ/SIcQ4e6sswJiEpI0NVE5wAYt6Jxd98
zS+GkFeXgpEjVRuizfaoUTvHf3jCLyMik+wvzeoegCRL7qjYNEoTwotTmXgK
zlpiOAEMdCny9K2hIGSyPGIDSvff3xODf4pSIeHiHJVZlfN1Q0KQpleUsurr
VF6bWafNnVX/4VflseBkcKlRteFOULi9Y6xGkhl1WEzPqaPl91/SMny49rah
wAOHvVJVa10ZvfBbofmrWipsf7mTWnvCei6QJk92WnA1WKAglqroPxi6jBm+
Lj59ice0B4qnM4nA/Aw5AJpQ5jAXXyrmaYXprn0x2dIYPqOBr8t7D62wT/mW
OoQzvLOJ6Xoq62OsyOlSd5un1CnMI1hwzJPLfnjbb1EOozvCBXadCWt96yTt
hZGHPkax8zrplE4T9+Y+7RP/J2P8sVjM4fhsWlkHlPMX1k7W+sgkLfYbuAbf
vyVpIkbQecDZ1pl0Wu1Z5UyJjW+uejW3HeimFdRkl5gN7babpOaoKMzSnoLI
bZ3Otmmm17vc3EMF9t2Hd7vZampKvNfJV4TFn9GVVhOMCpLbm+t/cRpoY7IY
gpFnLQqx2lRDUjCZg6n4KCAdnbnJ8KuoY8XTbMmufRAirYlDg1Z9EiO4C2n3
zcO937ajDdWlqpXHCAFMubBYR2SnPE4Q8BrxZnn54kC27u/O4u2khJ/b2xEN
1H6kK+qNizlFPNd5TDASNbd9h6Zf6bfraSShwt6/GfxnisMqC3yJ9EDa2DvV
Bt7AvKTdVNaqI9nUYS0Ps9V1ugy0GVpY9zB1lqKGgSUdUjhpMfYtBxm8Zn2H
Gs85En3+Quofp8A0C1MXDIoq8K5EPwVYaPpJzEoR6KH5+Wdd1xTQBcSOql3p
aDycbn4tjnZhGdfsY0+739hGPSmOFfPfet0lMGxUuKUie8D1bxcpbaOqzphj
us9qpyAkqpmV2NxxRgODMe1eT4VKiq2kZ6YES1hozkng/ugiMf6B6mEVzQA2
AH8ErOMNUPSME7N0oUPEqW7xAwXqjifeupbEnX+kz3X4+B1YLAgkYLmHdnge
l0+2oPJpLiQCmAGeW3IpkBf++7XNuc7yM8KtigWwukxQ5hyztA7IrACqxPGe
c6QYIwsAi9JhD6rxGiTtpC4Xd9yB8uU3PmoA6y8Jl3Ie/FvYcl4ZUrmcztvL
4OLt66gt0Ijak/J5ojSJdtGGzIXSXAkxR9RWYRsh/rZNKHLdtAyODYP/BWX7
6Y3kQn791VkZ7RLVqAbnfb0o+vs8nNlTAc0XwQkquKd+hTPfVowGdDhf/j/A
ubh19/27kcN+tv1a0p1KrFUvPqg1kAm/GD2SeCI/q7rPh91aQK4eZvzXq/FF
3Of0YYyoMlSxd2197eEbWRrSQ9+Iuzd7bgLkdMvfERpcNuDL280j93j7Vvjm
VkuBw003vh7qCeoLzYbjJDKJ3IOMdGbyL/sQFKIegbBJmQd3pvtLfDT20uzN
FfQj1dWTQMbtKnTnW7Ec883dSSlI8+acigaSi5qgahxYB+QsC1UReIoN+Kd6
6IN+5yi9B8OoFSGQ4wy0Mcv6bh0vUlY7E1PxMXvf+IEcFDDfoK/uFMTMFzvU
pvXspYEWu0bEDXUAYEKumU4YCi4AFk875Oxc4MAVFAMi4jy96Ca4vhSzUZen
8d9y1wK8pnAz+IrPOCUNnYojOya4tdfU6M58GZKcbfXUu/ok/dmNTEaWyfi4
0kmjxe6o86riSv7JnFCUJy77ujH2kx6YLm4n1MJECehSb6tCRpqCJdrwReGC
p50Yr2fDsS1CmThlkTIP5idODSqEzddEujv9UlK6qVPAMbSnKzDON6g8xFBI
/zchVP02n0Ti7Gtz3SA+afhnR+v9w2PdKtlEofRzt/7h9++/uVj91V2B8EbQ
ZhNxe1M0eC43YmMxAGP9n4hoRNVT1ApNhjDns2Rh5YmbkCyGtAcCkNzwdxap
XsplxM+tKjmmXSIY5F43vFi8t717swueuvvYJosUTw53bkFBiJoMPjoAT0PD
Fkumqzt/J17MNPi6eo0Vt7/NXbiIBIXX0LvvH0xw1nVUM8pcptkBsrfMkwhS
VIewiFAkEKDwzFUt7IdCRU5oWjfOuwu3ZbC5R2GZmZFmu1xb+OrXSTvhMMQj
hDs9dlybOyAm7VtOQtp1UZPKfv7MsdBaIT5Wj6TJg0fi/yaFLATVueA/EyJ1
/4ODEYBc+nWRHvyAN04asunEmHk5ZeSGkwELRWltNWeutIyyzpKn7h5p2OWQ
rJq7nrfbD5OZaspSRgp9JW23/6nVcpt3g7zrb+UuJFg8AL2Tsw73CgvuLRiH
zQ7MBTe05Lq0VcnZ5pt9I35rRhHcOQCi5a8IsuLDp5X2Z6rGXUc9CkLwv8g6
Ez/f1GlqukxAMvSYDdzI0iFKrVbD55EzDLoWL733XHGF7j+nYq/4DQw/sXP1
RSR654XudLNufQPGmmvOw0ArxbVyBFw5/ux5I/3xE9SEd/ccnZjtAU7k7rA3
kYahYWsMyuaIlI6WxDSEpDCkw1ZZL0gJzBzwqCWe8Nt4W817WX9PrjZCou3t
03Z/Bi24cgqduPGW+/l2+YU4sOPwgTUjBIqkUZHeeacsoGLCYlZGpjF1Rxei
V13SHJuG4WOfu9Pt/06s9U7EvNftmzsg84kLrJv0x2RL77XGnbR34W/lzNBq
SawSJK/eQ9fs5ULfjvizDkicvpsKJcO3xj5wf/p1sYcpVVofq+uLe6bG8Ke5
5lWnlwWGgKKSbj2ITogu9d+EuiIBwAH8hW8x2C0hh/otEiMaOQAYicr8YBR3
kKlqRsYyG0yhfPT9Mjv9onho9Qv7iBy4zpYWjBYAKqX7aCBeTcMVagrLGisY
AthPvVflvPRD0/LDXt12jWgj38Ift8J4CJdDoHIRzvrRJ65Mb8vQVfJc4zuc
kFM8k5fEyhvLy/OE9k1TSzGNgjZ/+Iziroa6djce+kEprAqGqAk6cwOQIkT7
WkVyXc31nwjI8NKmWC6v14bjxus5H7BOw4tWat9eVfVBnRIPnpZ/mw+rdPmu
rAY3Ta/+WsEqOcrzXbXMTqV3QMAmQjvpPV2wVKMxtRqNEpeCCJ4qDjnL8JhS
aaF7t0lxBhDCVqNxHiPHEaGYhOeufDQ+q0sVUJ3rBJrPjNdR8pJnLx/DrL9V
iKk1hQqcXOCqhu6js4EEMBeYmXUuCcu1LN0d+NSqs+5AxL16WZbdqBa5KTr8
7Ngf9PoyJC74wGwUaX80uwlJUrT1u71qy348QVk2TTAoQObEjFWOH1HYncSJ
hseE+cV7NrRyqoxsvh1HjMYwPGsdrl9jh/9IBgKQ+H2qTeYroiw7MsT2EyCZ
JNrahpFBvCl8DkYBcdJftChVSVDA0eX0KwnTuODfQl7gB0a+KZ1YBkZzfZZF
HXs1JuOOK4NDq5NcpYYGzBnrOWL2A/tWkRXivZlLd+h63AtTqjqpU2QgmUzm
03oKmZ9Uv3EW7AF+uIQr3gOJ0lmxyfthDfLOQtg5EPC6/bCJ/ocFhah6Uvqf
VvV4qHhOl/mRWFcfc8eAhUBcuNOB6uPNSBYXVWMEIuPfnqPyGPY7ChFYkeoA
h5zEMM9zG/ZDgGq5l1N920Xos2un1P8Qm/NXk2a0EyvhjAmbyb9bkcaSJVwg
3OgJK0or35TsGYC8ZWdacD7O9H+ybMsHIcRk6JHsy2PZ44q6c6s0cdXlEBNt
1SuikOyRNjC+2vP2LBNQDEiGEN2kjzgZwbHb82Zxt1gGJzrWgDiSlRXBgJNy
GmIfJryyviUQkZR3kbCic++ao0SqX9WLB+NSYulS3fLgn219ioAmp87sqccz
wlSrFLUIkq/bw5HgUAIHoCWnvn/xL2F+Jpiav/vVy/1cg9A0DBE9Aijl2yQk
r4D3yR0IhZFsqtPhIonTZ+91UZV73zcv/3hZMIlAKU5n0Yhj5s0yno2PtZkf
80CzaVd0jJKmBsqpo8IRTBCYAGcJOUda5syyI1oqFw2rBYeX9DKjNP2rV1gH
2AKzE4JE5KK1AjfaOgl43UiqctPgM9olATX73qMqqoeUyLNEPhM6+pzsV2BT
96XWrQYwvgF4hsOfz6e0VWZ4os9ZRcR83VRD0fcATMZ8/QlR9+Kg0H7FAqD0
aJ9CoOw45Sr9gyYJj2ZHQpuhEutTgMPY/6XSZs5+GVCGH9qhBsNg/Ew08ZCe
KEFOLVD7zh9Ud/jTJO3N0eWya+FZC91YUEiKdQyDbakDdYj8ctS+FDJSQlJe
hbKUKaIwGzthYk+kW+wuWKw8ece/WILFLoMD4zfOR79mpZTJ2S9zNe9V8kq4
IKqrKxIJT/8nbT9hPYpgDspN+eULxsCbfrwW5D+kqaPJchvyMqSrOtQq2gG7
UQKAnQZnOnnz0l9im3PQaAICvuQ2aIIjmik1YQEzeVgb7ssxpINrzS5uZw29
cm+MyEX7sFtBKM5G3jB98opkajRB+kIV7DZycoxQ+FIK19lQ9dI9XA+mk/9s
lf264GQM8X3N9O/GQjlI9PYkVsIWqFLX+DKN8Vs3OV4Ab0iRrtb4iaGY0rQE
EfXaC+1TP6IGHNL/anyfvurwmLMNTchZYfID0R/0kL0LRK8K5Cyu4+021Tx7
VKG5G/exZlWBV1Ef0Q1GHpDPnb2NnCumia8vDFoWdni7FSUW3Y8/z2IX6Lc7
4pfgHwrtBAG+2VhsebU3UlOF0ffYYW3tmwGjf/QXfyvSQn4ZV4KeBR2pzFas
JuhmuoktEdUI+4ShNw89ny84Qb9iMQ7bVV0X68glB4AbnJnQZVeFA3IK6HMm
opEPP3zr2zU7OU2g6rwMz1U4orUgtaM7URrjMFYzs0dyr0XKP0j8wcHUt4g5
J37qkMOdol8bZrs7E3Zaf3oNIA8vYvTFHxa5YN2H7Bbylql9rP4W+92Bwld/
EdVrc7K23i0NIQProwEpddXvRFdzxtN0u/eHJI+Id0HIfQQzAtKsHCzmeVkz
OzHN3iPtyY+CE1Yp9yyAQPwLbPxu02ckt7KK1XjPOPLgZmzFqvKXzlbNPIks
ryjgWHycGzaFajtT3DrP1qhP7dSy5NKn5QqLDXSNgaKz8uR009SVVCdOXAgx
nFjVAFbMQFUA94yT1FaoA8KfBUHe6BBJw8sYMNhsMw7jNiGzFeiGQONZSbP/
seeNEFfXOTb/s78ipGVPlM/z1s7tkc63Sv7TTq3UEwFPar/fdZ6pLZcHkzRL
zrl2KLybQTkK/Z7u9HhScPPsaPpJE600BsBJkiinOx2i8zz7FztqSuOa9Pd5
8e5n/9JnRf1ZU+rF6Iy2gDVMDHbZBzLkV3AM6nucEjCyTa1tVNivQ6WNXkBN
zCt8HVYrMc5LfPKgrlc920WkJ+qgA8lUqTysMhRZB7A7FS6nnlhAf81mW0cS
+Dqah0m3MvRvxEqwXT9TLyR1VB2Djq9fM1uyZNXjBiFTP5AFtb6KWdemH2ZM
g9Qk8sHQC3FY4i+jjMGUztCcSxxNiv4VVw+AKO8+6RDvNVuev9bvpuVq21Hc
ZZBvkBwH1+ECZOesRtXDvp1joRnb+5atEZMQS3tYl2SMTfWw3dTzG244IxYa
X0L3Yjg/nxXuhecieEVwhtV38xf1tefggCSo70+uupXjic5EUA/PL3zqVeuR
15l0fqKthXdYcoAJbBeY+cH3WgR7jNt2OUI862N94tp5cR4THA3ND3CaaCqc
61FYCOXecCwQ0eck34t0RfFzaQVPHobi9iHz/yOy713nzXGuelp6kkG5+DiR
319fYkiWzzfOjHWJh/0bA8rppbkciz3FkvQnA8u8cuCojcxfyhQ541M62eIu
65EAPbzUkhGF4y7mhzqlY4uVVocjxKPCldAzcAlQIY+njeWquuohrh/cqRgY
UzapG8pyoXbMiwygbp2LVUUcbq6xZMfIJQnssRQJoflPqB67alfWAQguQ4C8
9N0HMyWBNEkLFmIjcaNCcv3CEZ+OVstL5jcF1oLhLUPkloqP94jPs86GG2Pa
9cRNF3OiJXF9hNN72MEDzvNzqiQswbhObFjW58mJKDwiE6Kk8gJXoYW8ymnh
vbNVDk9ZEe3HlAmWOhos+oNuOozu/pzOIx4MQEM/lGZKslN4hnLegnl6uU9r
OuqMN34xI7N63XFBQH0uQZtrRo96tX4lZF0eMWQtQFNWO4erZlcOgNpAcCr+
1jUXbu2VF+vZDQEwwEfQyZbSPK6CdgPB7qkA4774g8bPj8ZxFH42PuFyQmFk
R+RcG5WYUnRU8DsCPNdl3b5Qzalh5fVBnd9SOXAODIKuseTdlEUS4hen9fJ7
3UnbDY6y5INlumJSraaeEnamumaKfflIl8keXx9jPIItXyXAEm721giis4oF
ebl5XTuXhZqK4WGAxbWqjnsZ/trWAoUDpgr89QSz7iygVWKly4SPucFDF4kx
QlJTz/OndUwjjGoQZSTQ80PtWez2/9AEJr1R+iH+IrnqMYNgJnIWKiQAxoCY
EqQHCeMh3Y+mPStIWD526YwCk7WmGuh9FyJCAecHj3BoRMjIIEUqNjYgVXx2
QXWUw1+H17qJiVh20kUHrF/jceONEASi0k0ZNkgE1eI2OPHHNnBBgHRDFKhW
z43wIIf8i9MoIm4LrhYzBdrnpLPOu1wFOVXHpgqY/l4IQQQ9S7zh3EUfPVpZ
qfhYrDE3FOqUAiMDOr3bC4jkyUYVRONeGbfQzlgaAfjm95853j9/Q3N4kRR4
8GW+xs30YMp0t60EfqsK0gZvhLtv/ZuJU7v1hZ+/ObKLxMpTJ2+3IOTx/QcR
wIO8yuQU47xIf4XaU30B4HEcUlSgTalELL7ZrD8JrPGETI/F3CKiOF14d5d/
vp8o68a0KxlykpuH+HP9DvPYFwLTIGa3w/qQq7CdaJlshv9nx5KQjY3F21Cz
cTmND8OUi8cw5RLgQaOko15QiJTAfKRKBRd+JJc0ilZe2Oqh3DBmJWU2gZfF
fkPYCR9mC3RxFRUD1WaYvS6fsEzPEHCfjOvLK09sHqZNDSsIcDYsO9EtYaYY
KfVfEqpWZCCtkG3CevtCiuaCNZTQoo8ac1U+N3otFHRmxj3/BIMExjOVkmfM
0qNVuJoUwzj2RMYoxNbyiheuTf27XSwVnFBSe72keZRaee/TR5QmvLoczY/0
FU9m75XmbXXZTc4lv+PbX+uRqMvUxbIdkV8hd85cHIrEak/CQYduEQjn4IUZ
t3dobKH5YDUIbCjYdK7NACTsKOTv1/CgjAQxkSIViI82MPQZMSR4azB4cOXk
aHV0NdPbFSLaiRHsMY5KK/rN5dSt5+ToEyMlX9/mdw0crMpDn2OeYZ6DLP79
oj8pVKyYC2st3uyd2kYVabzK1RGhSx9kEfogyDGNAhO2QgBBFChp++5hvJc+
3wxgBeKf6ZvE5sm+I3in8LbGH1HBZPer3Kwt/Jy6L0kHU053XdJnWzXplJBX
jAwa71xdOso0U58ZehIvhqovNAooqla07uKqvpIOvyaqEhCagW2cAYz8DnZQ
wCa2PaRD9nHzQlJH9v15NLwl+c/jlKPQIhi4bCylZ9K+nwePvMxXycn+HH8J
kF+JJ7t0i3nHCYi/8Sp+JZC/XigK1gLS5j5v1E0GOXSkxTidAM+MhBuAEplN
WHCPSLZ6a8DqOk//PfSSoieTIxh6JJVadvjP816YeBPSJYbtX0iOuOmNli5z
+qZEdVNHCM6hAd/OlLwBhwJWDUzJ0RtT6Wur9HnWfTSUzPGX6gEbchFbAIC5
bnrVipbDzLGyT6GMeWJj36twkvipCxHd1S3sGgA5YVWRS7qDqzF1EFzrzFHC
4mn366suzcITl2GkDadPgWl74h6TJ7SNcLfDO9E6JgG0Gh+76qNDhLa2Xmiu
19zqgdGvR45CHHDpHIGeyELeqajl/eyJh6VBuQzJWRPrJsZkcrfHmExDVijy
Sw1rNpm++hSWKasjsiibCDKfSKwsUMh/yrjO4OwJcOQGk3ho1nnP72m9JYSn
2ECUknibE0gKM/HieQ+2T/PwDitOK5/QGfkii3JN5k4XiaH7b4ISMeIuS6kf
09PUTV2pybC0aYftC5UUFJE9pDxli27MD1/+KrplBAC9wE90mp2VRyeX+Onf
kqU3OUZl6Aq20ofAPSt0T1ms6JhHvfKFuDnNhfD1aSxzPJUPvwqF4hEH0mBu
KRAQ7JhLzvLXIsaxO5pc7tRPZ05/fUBM2T87YVzcnaCbSnL5aXfKOjPb8nqE
2b35+THOeY1cuK4o239f5D2jtPMl9DIzpgCTVzCAjtzc8Rna2Zc9NxZFHeUX
afZWKjk8VnHxAKOlIVFaVYfMD4k/rP+FWnxBKBQb1r71YUeZ0L4KBhdYZ28k
M0xtW71AotI0YpEISp2caF8KNoYuHcERqU9oI7Jqa52yKL5Z2eqUwcp+49GL
cWk5QIPvdmKvS92lbNRU6SmaEKfZ/MgO3NYLtpCgPNoRJVGefigpiHXuARza
7AAztWNJyHE8E7nio1L89CYmGAShCq221VDjZ1VWmWXu9K1eLBmB+9LJyuUh
zQJGRcTox9/STE2Ebkg5Jgem/FNrorgQU+4fUigiadCmikIlePv43Oouhpm6
Iapdfb77OwloRiPASPYo2NUUCzBOGCsG0JeQX8AgqvCs4DZZ6mrjROFqS3jT
gNAqcHKgn6IUu4mTyvsV9Qg7vm4Q2XcD2KSoxkZzsgnSRIkHUI5D9dU11CJD
uBXNye0OPDVrfx6R+wz7CTVZGVRCZm8QS1rd8ndcA/7IB1Ym4uiMGKGaPnyS
kUn1vIAJesG5tpbjUs8y8PpgVln5YowOSB7/jbZ9L0iuaYuPI7JpX6Wtmz4x
LRGSDeCXHyus1ZdU2kCQrUWt8bY45CwFF7AU+2cUV+tLdvEJ8cgLmb3aMIn3
/AnkB2A8NR/JnExeUgNhIEc16EAaJD8iIF8tQbjWxg/uq9V2LhXkN6aA8kGL
pUhiIs6jMhRbnu4a5pzo9LEBGZbQ4d04PmSxTp39j07QRTHVvpWzjbSsvFiU
QwkHozG90Q5uwon7ruAJ+vACkHzeE6nHluXrp9Iv0tfrC4hPR3aYRL8v7t71
wy188xMbPWAQDYFneevMhj3RPRAP0Qe9IVjc8vylmmR2fR1IhKkhVtfrHoUX
bS/UItETBOeGO4GAI0M1dZmsIk3uNH5sYsJBrWNHBaywV1Xh/acQOeLEFYJ2
Io29LXZPrXS36zu/ljHxGw6Pl5cqI9evMuwhYvDzhcE6zyUL9gU8uEjnt8SF
6nuipS+FKgXXY7bu8wR7POop6W+1RA6CJE1nBvi43NKCac9UP8pWOYCq0vVO
Buowhy8RX3q4KLkCbYnPbUoefmVfNLl+2KcfvsmDgbWmzpw8po7hHFw0zBB0
wjbp1DpzyY17+ERZVDeJJFPwtv2nIuvmJyvRqpMYz9TLhsnTug7moYXBns1U
kE/tn6ZXkYgihAAq1ZqpEhxZ/L2BVGNfzNF67n7NgKbOh1og6MT+sb7itgiE
gJlNxA26Q87d83vrBhA7/zdtWatYsM60xFigpBCn2r69PBXhFHmv34y4H83a
D9PUNAybx4YF6y3EONFvj5O+ADmvMWBfogWMk/vHdbrkyJTvmf2U3HMv4VVm
19Tsg6jeQfrwl4yJEElC7bwoVuvfFYu14S3uBpm+TNGXTHfpABbKV8pxjZzi
z65mA/UDKcCK3x1Yw2JrD/uviAazbOMS9rZPeZR/622RTqh6Wn9knhy713aq
goP9u9UIPcRtmfsCUA4ImvbuiXCX8mx25ys4B0XMWq5ois4WQJa1QCsWJMcm
puG20aCfaCXFqu0NYUcPTvjRZkwggBL/MBv3Kf1U6nU7Bt35VSj0TnQyShwF
LR1HRwCkly64L4UBNCqhIIVNqdPsuJX9X3wl2md0K50mqIGqRAqNYQz0ZO8H
8azVYEPLmY7umalDBt9DfZ9KzpipHhaEhZCxCibSmlxk3c4RFEmQSSiDvHLj
tC2jPtyOPed/Zr2XgP/fppNHhTItlzpy4OllqWM7vukgM0pGD1ahKkj1VWGw
xugblET48zkyje/8HO7OBHkITMglM/uadhSmFhZS5uxgTZ/z2y7gVHXSnraZ
E25ApRBecwjQMnwXsnsM5keNjFmCh022hMNIJdh6MXwGHjeNR3qWunBbrjUP
J49viKjYZBPc1lKu2GqG8VqyXQAoJX9tMVBpmlZfIqQsuVpwXOGrS6IpjwgG
2+FEotMbRSoiGb8tObYhjwEHAGtaTD3xvuKdvk8PKdpgvk17Tc49a7pMdNrv
mNN94vmQs23/JICnuKM58ljLqPrLEMjTxqK5+AlxOd474EAOlj8AX/pEVMgp
OPx49yKnwoS6FPB6b22PYGSGS/RAGWH0EXGtZZ08Ia4cpYEoJiguasEx0LQk
DgXBW7ViD/xwd4gVkAM0IqWFXyM/ZKlOk6lUumkPo1I1/+7zTW4ESo3injLU
MivLe6SPL/e3a6OuDYnYSwH840IweM+rPNHScuPuh3bxvPMLGy5tSEcnTb2+
V36XtclbpNzRJw5phP4u95RigS5htO6wFekAEzjzjPV6A6+BIEozUpSTRVzd
aYi6s7KrEWxBfLbmd9Cpm2Y2EQMFeLjkftn52CaZyGXUkqrLFDgehhrNFGZe
YTRdzKJqikbH601TkHBQ5G3skfAtfOhxVOdPhBGDN9Lw6Hl8ocKQrWVGxeid
8qJkm2g0EAIbC+6af5MSK01Z9p3cMbyTO5VjV5otDx5WmxrwJld7NbelaQFf
/dXmsMYyquRs0PlGYCFHamF/Xn4zAo00vHMzynjzS8W4irAtwXhn4poTMkDm
NN/7EbB4VvOqLM6OV6AH1jvU9Wa+NZGgIiNMjBatJqPl8ITVz1vlgZPMpGmf
YaCYqkHXv2bNPAeVE5J/77ddF5WIOU8Ngq58L0wFWs5FyXsUblOheTKht0RD
NIQrNBZRpWznfKE3QtFIgSEpeVnmCg25fsCW9qDlTlWr1JTUllJn5Iy8G62m
q+U+t8EPBJ7/eJmDuGDz9/0xU1Gg+xq0iLPS4wPoFpHRT3ycazIftNGZpM1T
RfooJZbK+5hbEcWHwouuB5xVUyroDGgcP9XO6rqU+WWKbDgdr/l98f6enjig
BwxQL7RlrefAIQXGdiaYNO0T71uAo6a9xhq6B3/m0ZE/16NvoS0PjNp/5yDU
rBOD6K1IaVJGTLxn6TtswKQnVujAsx1bFv4nK4kraBtBVHUT4MMQUnbQ4OFi
GOBqOlkwNWm8Q4mCssUFM6q16J7RMdXwleEyZGNh0zM5SonSxcKWI+9y12nL
L9ZNeQViuvUrARzY0DQLd5lsVt59zcAnxlgvasUfQvsPpMjSZI+N+rly+F5M
dQrkhWSbEeWFvg6djT5AFIi6bHVaG2BpiXjriaBSs4dtbRvbxQ2LXy1HgEbq
Eq6U23OzTUVcAHVJwXHqv8rr2igzcKArgD06aU40wTkjDPUAOAbJT2eYMMx0
Eb4MYzzGWQTi6/+ecxG3Xl7zNbScBgAW+RDWxV07tvuP1gu52lgPxbvqntAI
5ZcqEWmKxa5GiatzLJnxNfKSeLgQWLJE0bu3n/f4YCgd7gPD8XWrOIBhmTao
aqTRIEJ2/03Asp6c42dUxI9WPWTGU6Zhbne4ZDit1ogLyslytq8FWH4srsAl
XsvtHL64J0sp4jaikR8HaOBN5i0onJMcc0CbwD3KJEzT3iQBVwPrFKYiNsSv
04UmCf6gOp20QhkaYBeyi4Tlql7Lzsk7+eb/rGb2kAsnU9UAFurAdqj0fobX
jb5pnzzMkbcukaBe9568cspN4I9CNVjhujxvu9OytSObMaWrUQD+idpbgpgH
WXQw6ZOTVcaBsAIXjMRBct/Fm5CDD5TBrzC/Nhrv+HqcjP6eI6jHpTMrpV18
WRr3m4NG5xbLH3PgqwPjn4IWbDWoIJV4Bqmxf0l2otLor0us6dXzAFcO7IVr
a3vBdoOOXTmo2qISwKRQ1gotUXWT9fzfY2f3jEJHr0taUDUZUFZ0cI3jTKbp
oy4a1Qm3r1/oCjeYH+ceq4e1I2YKJlJb//u4HlE6+wZWmsRwPIGXbtiq6zQn
dXYTP1bbneCS4yZl84RIU/6yadoMUL3FCNUp+QREmpOxxaO6811X9CbT3et5
LzSQJJCTnHWFW6YT95RhzHk9QWPjbHWXA2tLz3C1oOf8gK++p2dLBF2+9rO9
o6Hyw+FhzFYGJvHi8DfuwJzr/RZYbc+QyACPmSi/pWsaH/cbw/JAeg2jffte
8T1/uINRtQi5CI/W+5oaLxtzLfE3VnX7BPa3hu0cwhXvn6AH4lSUQLX1a8+Y
0Grwii6lgsoM8+OBq5n3EesTYadOhw7w2a/dElkPE+Nrfmeo2CN/0wh9k5r8
58Fe40S74tZx/k2c9gS7DFlkfqOSpauJbz6vTOCOakIshLRENd3v3TPKyHwr
vdvI6BN/pE/0jHNNTVPph9exvuNNPtUbd6OgxbRcIQstX+G0GjvulWVMneLG
Tm9SfnkdzsmMplsPQ1B+Q5f86EBMXz0sc2mkqkEDfLNjkn9VieENZvAvMt7v
z/i7oeRw0zWR22XBbQz/LqMyLHjjG+gLpdT6mtsDsefBFvdOLRZ1U+t+567P
clY9ZSKlE0ePsqLfCXg5Nzso970x6zjucOmuVKsxhQCBbcYgb0AGZ4w2Ssfm
yCkwQyHhGGoJigOos4Jiu65852kqsaYlUuprpfaoke/ht1p6w+yETatqyQzW
ZAnTleORYXQPX3r+2VIbXu/1J1tVzVV4zBdaAMGjrzxpySsZZ83Ld/qXN+Je
FHPsVkdBZOb5nAcq7PdG+19Pum/D8/IZlm6btOfiTXGpRYtFblobiftIfAOp
8mmgHhbH/3VvA9ara420Cm0Q/gKrquuaDI+YeB9PB7H8KxkVa0E/pf2S5lX3
daKXSdBZmTf9eykpGYV8g1W/dHEEdClDUC78af/bZz6WEmYtISXRLhhTsFqR
3PFhwbzzvIu2JdZ1SQmiRul2WDlV7UglJfVTF3xkfPJeMiEzggguJDC7y0kD
MXu3o0NdJCUZdGO6nIu24R0jCRVtm9tBIG6Tmr2qQtmnPD/wl2jjfCAOiPMl
pIL2QERrN4syz0ybFY2NSH8gF8fXpCNjr+2O1Jp/9dIUQdDG/xSATGmghof7
Exq8t9OL0ZUZ3RtFPH1MQgZN+DZfujSzPGEnC2bUp3v8d4Oi0wtLJrIX/ZIh
+olm5XiOKxfaLRfpfvQKi7qLkPEh7tuFoNoZD9oh37yoDnmGpyR6eLLsLfeD
xKJn9MKz+4eiZbBmM/Wl4YhRODXdyKEIjBIGGS3Ohi8apuwoLtcIok9mVOXA
lAuPshfGS4I2ZB+DCvn7qWvc6mgog8eC07POvjuKI+Fc2+2Griw5wJvqZLl6
Cgq6qOqfu1qqUxdgVJh5JGv9wkONaxuF1ae60ZxF5c8sDqsdi+zPU31k0Y5X
LvASf/2WlBkTa43/0M+AMvZ7gJTEstvH14Fdjyc0BRQn9ycmrp3PdfFJ+5LX
sliWulm5SUdzXBx47bC7hCzYXh0LKXwpD0FcvRybynOsLMLOMO7VXJsNjJ9B
cBYn0c4ZiCF3HXuBfQmTFKglJ5dAJIg2ydNmYJorclM2zIZIvTLL1ZJFpDge
qK2sQvtfjTmcpqlcwExsRL++ASUDRMkbMUkmqp3bmXO96I0Qu8xi48pVjX8c
hl1LmP8sESMgq4SHLhCPAeb72COBuLsEzRuUvsR69TSnEltjyNRrQ3Zm6I+n
T47xsXfCHRkQUEjtxRTYJnjgc3zsRP/v+RIALEDCnM4bcl1DbXPfQ7fbYAKU
YRreDxvJz2b0dMB7rHiGcOJUMNOymYdnaVcjUPvrvY2chXPQKTbpJT9I6xAC
SjEaxVyfO22ohYmOep9gcqGyfo0lBQ6t6WwajerrlwARYc/LIQtSin1EDDZO
HHseXc5Z8r0ZlUHvk7Wiv5TCTf8A5cd0Z4YjVp3YSu5Zgy3vBroF76/cPJKU
FK6eZy/dXj3F91mbata8bp8u8ZHF0+HIdhv7oYSRR4nB4tnuXHCo+MMWP6T6
6eOgXswhos7Vdp1eSTn8hUBTaU/LFxIqleKRKaeEVPyHRsFmr6Fnd1u+32GO
NCqP0U1mSnJIB0I/EEKcdIk9mSu5Skc8FMzO5fdBKPVBgzsn6rQ35Puekeew
4tr9bifYBH+8EnZReLQbntG4y5l/kMGAAqVTiZ6dFl4WtfKXsDqyd9AhYQE4
u2QWkwZI9WpRHs6uvSsDOLstAVdaJA+RO2LYhBEozVtzTpavwrTRFCqCyZ2e
tZXDhrcHp/nX8WSFcV2o6ZlbbnnY5ZBWVvQvYkPvam+k8N6MJ7SJAVk9E3Yi
Yf+e2lvOWiIi2WmeiNJrWDpWFnTrKIfySFzdvJsRqPcJp9PReuIlo5In/fpo
R1ORu9aP1uPBXMG/QbasrfCWzCiz8i1R8QJe9BKLW9/CW+49TcjD9KF/ybbU
bhd2LbXl/PJ/oMGKPRNUy9hR/AJov7dHrcN5FBktZJslU+4d0djy2fvBHUsh
qxsFS3/GHbyXcysoq5RN45wXY1l4D8SzmXMmZFqZnmqQx/0sHSr/GHbyR2bt
3v8icw6mx8r4DuOKGofMCOrXeTHOxgdKb+BTrAUR1sCRRXvLEtUqRSWrHZPE
z00Yhz2qBHTcu0ocsG1lwUKrIUb6mDLb00qxNWiL5xMJFVAJJbHt3ncRWDbL
zeoEeP1AUnOZbyxDkApozD/GErYDJ2Qo72sSPAb8q/9S9KWAn22RNe/UUuPC
Q7Z92bvFRiNelMRfKLXKXeZkPCSdjW+mshqiQm3LQxZoDTKy31b6iaHnrjb7
/jFge+i5sr77uEvTqRPyOtOlb2Si1qINrAs7fxq/GGlEuwgOONpL6aZmZgC2
eB3U37RFCM8XKWolgfqY/zw1RVRSoC5vAbUNhlYbPLFjc2EDWx5MvFzTABYO
35yxnMKezRpNrNl8LabZVERYc/Zy22ybVcYUNotrlXC/tApbTNnlmfYMTFmy
4/viD7IBx7E7dt0dyTj5g3z8Luap3P/1DQ3RIa8tXK030Av/tTcPr4Zp+P1/
yUQKLQLg6vGNMmQHWuCnhaYEMwVUYbrdv9kXp5G/EnK61fkZCcUbAtYEbITO
u4PY/6oT70/D3bvucY0ABv5sBg3F/GANd1FSPnv7N7aMyy+WRxmBq6SMEjyR
mRYCKyOIQDxRzIAsGbe4pVeacGnDWpZlwbuZ+kjC+99FTntLhTu/iP+/Y+zt
RPfOaoEiSsvXVbn8MypErCpUS5NkBFJTmIfC9X/6mf1ADgbDxfAcurNn2sSl
acHDZtZzVcHtaO08YjsMCFDOgTZiwHn3OQrsSac+E3I8ocuPNqFh0vSYD7UL
WSyo9E9EodVXH78BSgsvzxAL5B99XNS0/MlSW5YNvKyyL+U9DYJHLYIWGnEx
pIUJ6eQYvzPOvmxsDe2H70ZP3tHSb0yY0GUpzkxMtsxB4wqUqlEcRnbHGteo
9u4zSV+n9aXYqVZr+eFq48WsnomEDekayrpiYRI1JvUC/q4NArC19aorgPFB
wQriSLfJAFsuN03YYyx5mE11qMsu/w4VpwVgUz4UomwdQAyACr4Zhxy/rvzZ
f0+LIaDmpxQK6shHCXcgMgiFYd7B2TL2HjthpeXaLUomPZZCvqNIKx9bU6jo
uGAnNMil+wZ55am9RCWnlGBQrCp1hThK28RWROxYM5oT6jLbB/xpGMz7lNyy
yyzl4xUGa2PoH8xw13FZtAfzLaT//hLH6UxaSZ/BBZzRYMs2ThkxES/fjgGE
BYzgpEy8wJWwUmetslP8NLbO/s2FpumzNjYtQ2BH82ZYTsRUuEJbQ4ps44hv
D4d0iPkzbnmOHii3i0/dAaK39OVi8QukBOSifMk6tb5qKWN3uK0zVXBS4Gdh
D9QhRu+GbhWGI9rJzPeJwxf5kePKrsFThcAdIRo0O2doq9qq8/KWHpMy46hx
vM1VRoHijUODUnMznU/DjRPWjapHnQ7gTnCZZdSEYyPQJ5R7IeeDjxv7FvRo
NHmMLrH66E+0xQl+T3Ixf161maXq6WpmWWeTfmV4Ze1DDSuYSrIRn+kwNtin
9SdITXkVmpw77IL5W+LkJuYD1ZZfT7mbW9qhl0yWzrcTNGZGhJ3VJkDCnN+k
mrUuGGAzKddB2Z11TPZIW08s7/1Bbs0fzOAgt28P/3cgXbdz6OBlGmP/28JM
TjXxi6rLR699TUlyywItMmy8u/qJ0nRoUh7y4XwwxrsQ4eGARYS6hZTD+MCc
aZ2c5Ykl6EW4R8kvNkpa6GQqYMGktkQEaFMjsviJ1bJ++LW1QLRwi/uy9SI5
e5GZ8CAcf+/roitElvCmalM7kIrOP2F/JHWah+w2PVaRLihkHpijVsiRRDLz
wB53Jlq1mlZFh8XPnga50YKZywKJmt/uknN55/P1cUldYQ6NLQoP8CvkegBc
89tClO/lluKIG1B35ew3z2/U2r+8WhYekdIyMVk/I8LIyHFlfgqmXhifsVo8
xkw0OG2DheZM+XwTwy9ulINiMidR4T8panyuhjvVRuzdgARRE3nfrnJM2YPY
Zs2wltIK737Di1ZrQ9g7FUMsqmW7n2tCrv9KzyoFMWAYlZjYy9ahoFy6BKAu
zIRkbegXLO4a6d/wy32psfw8rp9vXreAoue/5yJuORcaUU8fyu+r7xFeLdtZ
X3DjVdt6MqGYl2eniwVjw6w3PsxrD7eQDCEL7mMjMQ68UBYA7+/uhRO0UH77
abIzYp4COzi2r0pIDcOKkrn5WgWn5oqDvjKd7NsSCaL9deH6Yo/vR2N7eEqB
qQNQdTXVGhRveyGQk9wncuwKdoBMXZBae9m5ewMGj9aP+S9h5wVCTRDKpF8Z
OXWgLQdKhXu2BI91FWme40/IcRzMoGLyKmsIY3VyxzZ9S1C1MthskFR0TDaV
vKdCQcxTiJ8TNI9UVOtJfmvLGGJk5ypLerba2obxmUb1zjDgdNHkyt3uFHRg
fRZzc0tJNLcnm8bQ+/f+FN10WYbD3Z2hULM7/EHA23fRvswZULJxXoF/VBJU
DRTMnuRQxCEVXzdyrnRl6OAtIWGacJviVhq3VLYFSVVHPwxyDL/mvXRRADHj
jlvx5ThvygC1uQ5PwzBQfkBKg9t4oINPytuJxx8eizJUaSwx0Cm4xeu5aGZF
jwGsQOfUxqywdvpp37L5HSLyieiIln6nkJZsXehkGbfsrgFZbkSDdpNpifuj
aRmVm3tlZc0gEa1S5Q+ui7ikyy/F8TOxIv746TShmvYtNitgCTHNy8ibOGW4
CIByfmffWDlQkoQf9+PEzh8zJkuKX3eT9cSwNUozz1qUqsAQFPRpiaFYqOwD
rQhwyygG+KT0+UHA+9jcEwvCuxP0rWqywdDOrIPXDr9lMSfilpmQobNK+L+n
vgb9qUEVuRZk65OUW//Es2x59dAi55ZaO2ZsimahZEVWkDtcJaD3w843qO7u
kmhJB3cKV8KAydl8qteIMGyG544Zf5/7YadwOqW0yJ0cb9yrS7barx0XGMD4
t86d5gGOMLm2csPuPMpyh2tjKrBjDysKIXpTgGGtplMX96jOQ9HQ0Sunumpv
qFPhKHNEgiK98TzSQcmwCD5VcIKoNBeTrKqCQq+QC1QMk3XE3001iUkJ0mpc
SD18tjhWxpuHVbzH8hb5RbZdGTiSHyEKZWppuJ/qb7jcYwse+hV//DAcJXnm
zNWLo1BPBTa+rYLtyoK20sxROAFQlGwXLbh31atRInytPL0qyr5QIqqfvq7E
rayGs5wGBRW7hbAd/L2kq/mE7K8mP23/YOnyAw1LKaJPL70zcpqDMwEpOZXL
lQMiVjQhhkSEu5d+Bt8cnx39uumJ6diRQZTSFXjJQTYJcp5diRE7q9M8lFCr
QB3aOPU5XDLs3IDbGcb5Sp4gqbTEvw42xKzK1vFWvQwa7LZ+qLDG6bl5h+eS
mkYBbYSuTAEMXFvZipdPMotbIswOZd7Xkmbj/VEyny+47i4bRWQbAZGS9ox2
3Ev+d2O9d7ltAP78lKXUk3GBCzcMYY3v+3Q3nOGW2VvvaC/pvqgkK6tHTxUh
cEy+Wj6C49hjGEKMhMkMeO7zWjN/6UqprJ/ZeTOzlpdiwFpW+KKW6WBzUWUM
IZJYpCIc2k8cCzRFN/GZOyo4RFVgJMiMw9ybwcfbaCi57tUyVWcoUnYEZBjX
6qi0Adm+EX6pU/RDnoYtZ0V7c6RwoNt/oPg9bACmRFVcastmykT8SzGS5scZ
kYRl/10J5bB8LYWFSPVnQk9NXWH/bqFTXYIdBY8Bx0e0QlptKvc/OotsWCY1
0XHWPAF06Zwf5z+CZ9+FXCZu7oDxnPTabdy1iWqRzgK1NpHTEvCjdJQ4dZlN
X7n6wwCPJ/CwgdyOYFQ2Utkm+NQ9sp+RGv4SXh0doAMmmqs0VkKI3kIY1TTL
cFtcJKwJPoPrFHs3uLgdLdqJf4rZDg6iNmlrfjHP+fOTJnFKqQEhY3d/9fgg
qm4IdOa+PSaTtT4yOlRG26FzTT8OUwmL2OMm36qU6u3M/gjYAHs4J4M1PWBm
P5a/XsRiNp+QVRX1UPAjWVZxeTR2z5oNvMXf9sImtrrZQ7X0xdjYk+fNtG76
qJzTqTgr61fHW6xViboXSSDJmrc9Z3+kWTw2tAXMonuBBKsgg5A/aByttTTt
lQxnLQ1ivV+D/UD3ca79T29fQDSU4sZaouJcrN/HUGntkGkmCSNF0z/G70Fe
CYjuqTxjC9tR5wNm1LapXVwk4vXuhBR8I3PFL3T3d3WRfFFX6A4RTMBFSUOL
g/alMV2+x7lxZC7uZRhXT/+75nl3ucalidA0uIo3DjPBoGSQixiqTT1SnVU0
3HKc0W1pcixlwkXV+tIwgrkTcrTuxodKLy4PBWDt28H91tAaitvyOrZx3Ucq
GWnhupfVuOLOYZCl3qCDHNTm+oidqk5IsD9ImLqMDUfx5+vZL9xTfXNaHXSz
BG+u/jMcy8+Qdjf+UFctHBIBoW/fUiT0sNBgXwVwo1c5HJiax8wQd+WebxsH
xKNcm954q3x98qkexwZgtsBDbhWlA0KWbHYkkM2iyhs6h2aG+un/8e2ESud3
vOhwzVfgLuECifiX5laGOOr8P3MyfYhIs/HY2egckAD9roAQ8esGSlaUtAz0
iBcXjSNKBWpNrELMpbaKOUqrToYcbKggB05M17MpNzzmUIkjUZlcCV5S3lTz
WezQnypS+lqREu8bK4Q33Un8TYdofcaYEJBeuruIkOpt37d9CRDnnjMV3Zr9
tifzkKxynH1Dlk2rZEfRZ59cVDM1lx+bMXMPnOdGnmXFIi1aU51WFjxc61JQ
YuWfaUCZ7FY2W0r6FtxPCI1JbgQXuC/6craCoYC/9sUPrdO3BcKcAh1fD26n
toCR2Lr/EBMVRnEy7REwiaPFsp18kclpdPTBVyiAn9Z9cBKNgWJGG/W9PBCt
fF7tL5QYoMSan7UGtNGLghsDQdja9nn3SVTQ2xc5lwgEiOaYiCCeh7wCMHIX
TbMJgyaCRwqe/MqlRrcul6zBGgcMqSu/IUxXwAjEOlBI087lwAFAHoNhIoog
lBtypM6hGgjUNImz70ixHDi11ZrOdJEp7xP5008TLEJVF0XIvmhaIkiOoTOf
qZ7MVNPnYpBzVXpPKvfB34rI/U0TCKF8DsQXHZZtEnCiFQoGeCWnKX4co0SV
XYpYupnA8PsadOr3L8+WhkvRLbmYDWh4gffl31KoUavNN+B7+yRCMX/Q+bmg
KC4w/e7/7OiuTVqvLVqxSODsndqeGz9muzSh7VxawEXP4cghjtav9y17iI7y
DhfT8/H36aYYbEDMa0xJw9dO1iRY6ta/HDO1lEqi7dOIbRs/p5lLS3qQjJ0i
AS/voMNJ9T79QO/wkVylrquJY8yo2kAWYqV+IL8jy9o/L1LKiU0icw4uKnms
WSVqA9ajV0JZ0FZa5q7CbWIUV63clh5CA9fNxLcatf9yGq/1CuPbXBZSuslx
BEBcR0b4yZS9cJqsvrp2UZV8iA7Ix3bncNs9oLs889mvVvgwRnRYVED2stQX
0n4Ia0uP4ffhQA7txnjQeX3t06LMT9DbS15ledO2c57F+Cv/4SrIJ6HYlA9G
opmHRSbd/5O/DlPbLBtg5aqPG1QZdE1Chn2VtmGRm2brhT/lSmioD/3xiins
0R3nF4wH0yS+g8FVbEHQ7SniKklh99i87C27dg+D3SJoJ3lDqsuOe+t3TOwK
8As8tn+LO4KcpwlACSrfuNjwesLzPP6wZBBXD7NTwmHvOKnYAmHfHvTSD6tj
/hgiphercAkcJcr4oFv1WLgeMq2d7Fw1uEMOt0CuFga6AZb2lgCEJJKRDUhn
oYplPsGISBte+aYlhQjEpOSZ3DL8HlXoiISigttb4KVARCcjfZcesyry1bKe
tuQ94V+VE1EQZDSepr/J7tCVXmO0fEZeSqolWxmCdPJw9kMcmqqwpRKt98PK
Vzm4ghaK1HZFUL4CCUUIizC7tTdLP/p6L+f94vpiln/SxzvtfOOz5rDa2vvI
v77u+UxY6FD7bZlpp0LQSGNTrzYZnv5I3LVRq3D1UWl14aZJ6tORdnAl26wX
i4IDWVCjnYv+1KztW7iLbf39FMeAcT7K4wldl8a31wr+LZvpZmBavd/lCKUL
ip8UPpZPOl50I2dncYfvMqPBjGgNmyez7NeJwUIrPrzyEhC3/LaKGbS/40Tc
lihBpe41aLu6oCMxGTZJPzJTVAxwX+q5ehaOsxY+0IkPsRfpd7KiTJZDIaiF
PWhWvI4XVqg4mVyTfkaV0WZGHqdJv0LKE62z1WTY6vKYAchEYf4lsJZix0zk
YLdc4lCpvtLMorR9xE9rZYqkkNlkIVwSBLQKUn2uFvMmpJMtilfMVawFUvsQ
0tUGWyj+D8QaohORcRiA47ormfRpyNr2fUb+9sHDkNQZJ6dSjZYWT4f9O9mJ
5kFZ6rJ80C9Yx5zbsga+XpEplINVEYA+ZMaaKIUabbdSulX+Dvequ/SHGPAQ
wHfXpgNYwaFfORacZfWYGb/S9LeYf1nQlA7CO40jfqiV9JX5WoJGpDvSvQB5
6SM8Y29hTAQqtt/o9a6QP/D2kKad1HzoqcpaFUlqZukWbMdGTDIRkxQS91G4
SAP9vIooRvBJrVRPHmUy/Btj9umoFsmhpc7KC1z5IJPToyo+hRwIR6ckxX7Z
uQXhD789TxEZGr7M4kdz4Yql/QJGA2zCBfuQPjOBseuVKLA3ARYpYsXyy7lR
xv04Rdw/5Zxoj5h4PIDmaY6Mx8S1WL99TTdiXvtqFuykHgRbR9qbAPufs60N
u+csPLXNfKeHnJ55HdBy+8bcGRcJYpGdl6t9WL0Z/Cu9maI5V4I8Cx2b5t9j
me8UWK8K/wIKUO85SUBogd6eoKEp1jp5DhaAQj+QKByRiUZofVIb7vL+lrmA
mt4iMmfkk4uJ3hpO4+TkJpx4/qqFyeqD015dM3bN7PNg+oMmUFyJs1oUqYdK
yn5NqvwcAKJ2WW7Phr2WEQXm9VUmMH5Z/UDnJXT9YBPHvj6LEcZpkOn6UOrj
VkwzzUPlApVC9ru+SIJEnENAMN/2jRfuGIlXdYOjEWIVwzWjlGBIz9Y4rnVE
EfaLbt15mebxDyUyGoaA3tf3QzEi7aQ1RZH/fD8g6AFH2jBA+zRoMneVvubm
7VFNRIxBKmvijTZOfiPyJtDphAyZmIhUCI/XjXPeWRX3FpO/SPYF1ajibY+b
QXCGAPGRlDPphEQnpHHPtEFCbgOrfT24hjyG+TpfjD/Du5e0W3xD+kSHEEgZ
KXFJHWig7oidK70korDn3oVZ5qO+ERNkznNndb7s3vLyxeSdcLBhQRPNodQ4
rKIMJclaiIIsdA3Sx8l9Q+10HnAFeIDdafr4b6SyOa6sP98PPHy8ViyKYdZa
yDzi/xexWVvc/TInokTKCCt0HrbZ+BQMpNWJbqvhEHJObnY3ls11tj0ENZKx
CLuL49lOrowm1Ry4m0MlSrr6mI54v5Z4JLWytQ8iD9s0Ak49n+g490AkO/+l
dYmV6fRWIMOeLNxGMJHCE29R24vv3Gap3xSOrDJECX9XyXxiBxpCz2Kqy7+7
NCCv1EV24ab/klQ8/LCOCIw/9twCzgTTFveEYlGUBJNuo03/VIFIaUljpR06
PZxqqci150EuJ9QOqPIFAj0h1GdeeCoKJNlM8tilxdlBzQHYoPUtUcXLJKW4
RT+63HL/nJ4JMoZoQbvA8w8Ic9chJBSl/JqmyAora6EWUPWPwhyvx9wQxwbw
n4PcF6gTrtzfjRr7OC1zp7DsdWeW2acDKO4hZAk0S1/mZS6lZ/iV1N73Ie5O
MsM4+K/F+yuMjFzAz9g+PhGCmBZ/gJ6Oc84+pQB5LzjuaaJAphNrTfHTWDBr
YR7udy47hxJ3qhziVd4JGf246RkDD5Lr1evl1dXYpMB8ETHA4ry8+XVq6WFN
PkolPhrjr5CsDTpfwS+lLe2RARY5EfYEsi9IqBOkz3Wm62ZI6c4VEGyVF+aZ
vONF4HW9jxNsudUMYkFQxzQYw6jpK6S4spGjSJ6L+rdztaICwwztY69Gefa0
n/fqjr0s3t3xVOra+5KtgsnXlHiYrrAsOt/uCUI5vnnae0r7iMAxzNWRXrPh
u1NkCyXC3vryLKUYX/WZRjclUOE1rrZ2kBQCikAxgHCd5r8m0fLLTiaq0zqJ
1xlV3NXAxPgHYr4Qk0OIJbjSzdDXJv7+Mj+cY/rLGiOwXd/ztiUOyjScp7hG
VOU6jnGuqBFOSyUP3NlJ0lk9QcRfIFHzc195hx2XVI0Hq35M49SIfJ33dIcz
Q8LkSo7wzCw7NW20qsN3pilwEmZ60tT+FFgeSefniGr6mpuQaEFeRhN1SnQO
Yuv5x1X3EoLxTUjEa54fW0FTIfZchr14Ml0V6PSO76HhQio7/3AWO2zmvOos
0p7Ijr5tnJpXnQ1CKUou0egKeHvxPMmbdt2QWCbJsaSjEkTVDKv98vOGY+Cy
14tWxyryi+lKv2FPJ5oKFgMiBI3nfA5fhSyzIChjTRXsz0ZAkshwJ6eNdn0b
pwlveDBg2GENOdBoGw1gnLMJRX/Qct8y2Y1VAn6fFnvdc2z9gM7mZg1EjyzK
nTQt4eGcN+SqXUpCyjmWJ1Kf3LK8JLIf5oQRS8FK/akH8VI7KHmPB2yuScx5
hVSLm4Obf2Ulr3B78RZQjKa/rDaMFAuZ4NzeyaeinOLMCXNptbWBQuBf/A0s
LSGcbJp5lIUZWwQYIm5xI0AWxIC1SW4j+FY4buiCNcOs5o4QqgNvE4hDAS44
a2lrozErNeKqePwO4p2rAA4U59qAoWgHcWBspncLW/ABUNxiJwKniyQ8SUJw
ZCinrZsNxQdHISTESPQ6YnjeXsyLac8DEhWNgRRn/XH5Eo3JGC9hGDt5jA1N
pcetom2wjRK1TwD+riH8de+tWKyR81g+EP5aOqNzTK1TDF8f7QJxIYB0/cki
zqfrvusDjCPiIhHXgIrSWQgDO49934/ptVaCZMzBPWOkSkiHry8du6sP3ybe
5mQaP/oyC/oSgGTO6UF4cSWvshXWVn0A6OJFLxKVyYCtgcVX8FLbYtUIUb5m
Ahd1Jafwoc85CE5L6nr9DvPXGAjy7sD9H6aNIrLcC+6hfnREhejll/lE99WO
GSjb2I0wj92otdbSV02mtTUy0TxT0PgyBBubfQZEP9/kH+FG/mfm3f/JhQUB
sfhEs/W7B5qnk+oFIGDdtpHwamXBbOWeyc4s6fOAfUTT1AKb4E1KZydN75BD
mK0Y+0hh6r1DcxuawFN94trx8I8km3P7yQRO1Ctrx6Cz1NGzJInnzg/9kuwi
jWY1/+xS7A5+L5JybH5OT7gY7sQDzw+pHh7axNfOeE8bw0asY2jbhfQ1+8OW
Xnuf0dl3AQ2/aRKMnEBfi5WTxdZEx5+HEXsZGGB1RgwcfmlaPsgxeDz8S7y0
e+phFWufND33JAmubgOILCNrkn0LDW4vf3nZxQI/pCauN1PAj0X3Bo41WtIZ
pMf88PPQG+NUpvFg6bm8J5VK/M7nSrd2xTyLlHEAV4olJejxpCdOLUGLaK9J
7Yn2/cCmX3toFPcy6jJSy1xw2k2KCF4Kcb6fH7qdGFgF/Hb1L0urzqChC74v
ol7HxvaOvB4cJkZyFc36njj7+jhlWGdAUT6YY3rsVpKrPph91+z/WtO1Fvdb
I5RAcaDJeEypx2J1X8xTIezZZgqHqCCwwnG6ByCkikGPDIXGVGEc8ulSpss0
RtHUdFtnZFSK9KByC0glwtow40Nt9bQfKIX74B/UJECYQ7pSXp8IClHDCOdG
rcD7grErkQCbtl1Auv8lkgzh7dDrA38fHnas9qj7MT1lx/J05suk9z919Bfp
XaZnS17vVcvhN3QqTMbQA3wq1ife+QERFqeqIS9+u/SmBcLMn5DWULfmFNAd
we+HPuWT/drxSGp+bUGYMdgLyPI3EqCSgrDP7xPOMqV4eVVLne7hA1L3upSf
HTD7104FM9aXAG/sSZtW4RJ6aZcdqoKuaTtLky5h6iBmcByvwCRUPMd3FG8h
3r5wVOkIUzI5+qmfBD/Pi5CalqlEh7w7fYKNnnigIvu5s01s+UjocgX/g2Fd
vY1o1kjcMWwsNtWmt3LkDWXohuJIDuCcx6Ju6e1pbQOzMUw9trkIROgE3cOI
72I4SR8SrRs562v6Zi1UEIvZdeSzbznznEN8Ai8uHC2YbQN3cnMrQVV60ouI
+M+rGbJYGZLRPOb9/zEw4yraL/zX3SGs6oF8QewXMSC9NlkupON2oMpkJkf+
xaQpvhnzF56zwB4I4LGETA9HZyJsj3ruZUZ8MF6Ddv3ROt/V4W/BdL1ZTMya
+yEbu/4hWw/5Do17DYj/oRlrLkKx0hh9Uden3AntsrpZciVH6algFqMGxDpR
1B1pvbFsHwXls5yK1dLXAdNmKpYtNskxExA7M0JgJ/CD5bHVCrCNAxrnz1hZ
pjAxHlY03ovLwy+IO0opTMFJvtVLUPtPdHp02GXQ/CrVZxLbWxZmCamQI773
eOt9FYjNEBaLOlJnr8uDRPlBWTqLo+xBzd1V1rO1+EDQ2+tkxvDHdPQGU5x9
WW5+QJvBMJjbEslQcV0gRBrSPNwfygM2EGklvBM56sbmo57wq1uCZdka/r82
KTn0H0w3f9iS5ZJ3iA5TQgN7uiSg33AVolUlSpUFkGPpvMUoZY/55YXnzETE
SdqzctQSJhiksj4eOVRrVBy+UsIe4BMzshmgG4bs61uSbz5DfYDGcQATFWeo
gWW0hCueC9irjEkI9Le0Sfe3HWIAuwxmDXgKFvc/bxbDs/l9Njjry+z8dN+w
BCzvej+gCMShCGi/zBu2QX1xQa9FJaiMfZdi/vMmh0u2nSycfHiIq3N9+Egz
bMtaq1CYSfu9KDBB588j5Gsb3CgivjM8qp5SHN0T1Nqd8WEaKfNwzGHtIsE8
x1p8kQrziWQ1GlUKBsxL3N1mNcXf9UThiqkQugs6eQ2S9wYDH2wMHwEYFJdY
z6ysp4Li1XesJSpar2s1rQhrVO2bgHQ6U0mcIrMW8soGPUKeB+rmAoVYk4aM
6uzaIBxLOeKa5hjuwHkm1m0Odvb07sW42bNDqbNGjbqJVVzUVXcHDHKLtDV0
iB3zXdfEgRK40W4fkWAjBhuyLewa6edag8a1OE78gX9Sdc8Uv8oszEBcw9Ch
gMT0ZZS7ez4c5eYjxwhuUnWsVRztdiSnsaRl9zwramF0Lj2ViFX1uwHBdEga
EzqwdhBVf8KS6i6zjNFMVCGsC47toO3+Ck8T3AEH3D9ydJpyZNrn10abCqc4
sDWRuXu+X5TUDchjQvxZNQu7bnFLqnYMPBlM0Rfae7xJ0jmH4lVF+u9kEE8I
D7BO6ys7iQN+H7alnrUO3YEnAzbWayjGGQvQijhy/Lds16tgr8AVurH3xfJ+
mPcw00PE+/XNazx7UY6LiXiiOtPbZ5maQV/rU1aP1n324k7tM8faaoDwA05u
EY1qZD5wNefTyXlA3/WS6oeGgY6KrpQGgqIBd7ccQGqlaznJjNXHd5AyhaFF
rkBUE3Ofel2JfzUqC4KIjDwVW0I/y2bmpvEzXQJYuTijT+pUimF75M5wB3Bo
Tblqw/R5VPPDIeZDDR0eK0/UilEPwTYKNKqXEUQzD71VTbwkXSz4nzOjdcrf
ktAxXkFf0CHSI5QuOmdpu6jB+9JXigYn2WewuGywNkuEcnzi5MPB64/ichv4
/qnkhom37KiDBIrjubCh5yYGgljvCLj9Ca0t4QNWChW5Q3WCiUNpaV46M8Tu
iJwWR4mqhsGEi6zCL7QOGuz5iWHtPFWNr+7qNbV1GiradVxzkDr/4eOa7U7M
EIwK0vFUqpV081Gd5R1azApp8nOJVohHRveBt2dM5JsCpmEhaOesyIc98lfq
OwcaobDoMlLo62D1BXyKk6kIrwbKsHQ3dqsOQmlkF4B9aH1QYqtA2XpgmL0X
x+pJqSlNWPSFPfdKJatQACFJlZMpL/bsMGYGTVIVG1n9EQi2HpZXvZ+Z0i1Q
kmP+64YTOpxHasidV79Nv0Vw806w+U3JNclPVoK6xJmdm2n6IhfDU5FGOdeP
ztsdOlnVRFCv6BaFzMeOjv5ttR5/61lNWjXTy1VY6s21pC/i6f3IyFZ1dhwf
Zm+rzRfu5Y+INSj5pR5nrT9UziJesHT+Jk1YKAECtk64+KOy3q7FWU920jrG
3JBCCU0gs51Iqg4ISOvFBrS6MQBbYq+g2YjLikuylp0RbnOidKzjfXaVcgrA
EpEByp2MdMI6qF4No2kgLfV7VZLNxeU3WgBHp4SkUM1res/6xg1mNyxGQEqN
F9V9zuEo6g9BxQ9C067ciML7zKkBBK1jURMv61m64eVyRSVeQPiMfmdiskWo
dVZXb+/6ynZX5d+EVON7pVrGpa7a7iQwXbQ9Zm3dKTlI/lCPthjt2n2JN1B0
Dqj29Zo7ULg1Y3QIx3WcHwHj/b54GWLd6KW1GUesV1wVNtqVTDP1JZc8JtJj
nA3EBi+uh7XXsFN29Hh1S3YqHbpo3kS92BZ6vwV3Q3hINEO27f8MCjVUMdl2
ShRfVqanwCTacrUYfeyL07/lj6jan3MNHrPuvK+0JXGJGnQzkvV1Hfr4RL7w
vapIj8bA92s5VP1goE3YRe+afJrnkD90Qy/yScG2NcEp7rU/Wz88jEEtyNsr
Nb7aDRB/EQGfooTYbxnG4TOebIWryI5k39ybSxQEIHLDCBRRZRagaOBrBtGb
EFxs+1mctnoOBRbdtE43GI4Jw/LgaNoRVOArmCyDWj3WjLzxe+WyAL45cScD
Y8H8LWindfRfLYIxAPyeytcoGaZh5VmrUk3o/sU052LfJrpS7kpyK+z5LHvX
jncs9YLkYVxROqikWPLdWedEx/FQsEXsOog0/CcG9ZcSsGCDapcM213e3+8w
3HBC1JG5W7EQFynjZITvXrSGjlV3ZOklpCPSqAUQ6L1nGg4FP07XH4RNKneY
V6eQbmxij6D1MYpSs3nueTKq/88AG7bCMib0W9rtxJHS7Dzmia3WcFg7iaxo
yRb8BEV/I0RkgLg6RM5hQVXd/iKIm9DTIQsGSxrVHLg7ybY/59X8d/AtMNLU
gJBbHmNYQ3KyVQNo/bbI0wZb1rqqbCIUi76wUXShqUQw2nShGAH8Pmy2E5lP
mEo8SvHSg93+T2RAY1JPe3mwbCj+w4qxvzb9ltMXXvOkajC4sFdQTDr0wvHn
bDckBtNHkpECZpJW4mGTOjdJUxrXp96zRhZljiHiSeLdp2JSGm48ZSqJ8ULt
0NfUtP3Y7SijEs1TMK/lARiKPbPeVKXwsJ2denrbRzj+N8yayIuYYOfU4Irh
Ades5igHXQPn4XRJjHhoyJzpGoPhcz/Ef65qfxNvL2RSxBDOK+LpM6iFhahL
MGPBqP+dyY7pCVMh3PMglLMQmYwHUwXW7vetQDP7rA+QkM/7JGoSP07YBi3W
3QtiYGheFTr6pSMRMIrY6FZVBRIPkCWXznWJ7hTVhyd8Bk8oW/xkxi7Xvi5q
md8WIJmhNtyyHTXXwDQ+k+xplsUpGzYHweBcTeyG44OZasvFKR9hWDXfP3Ax
xwm0EmF6TTO3dpLtiG8AD+oW13P5vG/ImwrBjNkDxPn56Ow+LYtkH4/dePus
kSUaWLPCRKpryzMs+e9vNRN3lmJfsYNlguHo9jY0KhCavEhegLEowbXNA9mE
qiH8Tzip9caK972aoE61WQ+OWz24Hw4D+idQf1+nZRpR3lud+0r8231keDDr
wdykJt1+O94rmZlXcfC+OhbQypWCPTjz2+krv9lJrmajtrMEDT38HHRZMgLB
jwKnIvcLkX66U6MwAl0u7h89WpaGX/wktQVnQ/A5FJCNxUu+dxlVf/asHgP5
Rb2FKZhtxMD9i7cC31QCehTrUyv0fuRC42rjdrcULHRUEWXr11rtWVZ2nITv
uZLGtnCuOgSjbLEMxcmWwoF+GWDFTLU0eP9i/8D5q3MxJQ3TfaEHap37n4EP
b3jSyJSq/CLvTpgYTk8FOdhI4qEIb4QBoMUt6F7jxcQp+H6uFC86gG3yJM9c
emZA8FtuTwwxxN7ioW9pAmd9FVXnbQyBuXBWVlg1DqOUgysE5qjfnp/R3owh
sSxQM30dXPFYBkG6DHWCM7YjIB4UmRqcJJ07MrDvOWnqOR0g0yeCaB6J7lRz
ciKIg9mD3Gnci59HpDY2FqEE/f36vAQ4lTe95r7p7QFF9UiU0cdkxWZMOLQi
ylWKjcGtAmIMl/yt1N6ZBTzVZH1lqaNLJLx2+5HN3v33J56+hBEXFqxZCL4L
UaKMemR4yEHn514BhUYwB7gFtoOGRFQYyCC7Z7oCeCeTqbu1C957EIT+A3jZ
VpOFLgyrbhIrUr6ZxuKtlR6sQF3S2gjJu6QUh8cCwVDUUiysr47ywQERV1+V
tWUAz+iy/KpXKBY/pLXtiaZ/3rnEVsCgMigjEFzds+Ot6KkbB/KfnE0CmTqn
pWulk0mvpHoFx4dlHz5WFlcmHbkoN9/zElprIcLk8qed1/xdQg5UUwD/R1SW
ubdzwRMKY1qknzwNi5a7r0BkGjedwfRW/HdvFlPeABBE/M3mTsTaLqNshCwK
QEA9caiBQgcvdT4Nk54s5P8rkniDcojNOMao51HKo9U59bkSpkc3aOVo2yF9
KQE7s7o3AEhlzAXlewXuCFEbGT8jS9zha+T11izfMF32/k29kYJvAaWmE+Pd
J/en1zpRoNBm7JrgX8Zcz7x9WJ9iYv7wIc4M6QBlXX3BUF8erqsCfDV14NgZ
Kdm1pfwdAgrE1TC1PZ9cU337rCeUV5Vb73/kNJ7DFTmrXKT3Cm+6AG978mle
6vqpMrzwSzVdaviHBNXLb7CSTo1zY6c3P/pi8JJhPnNo2l0PGZb/JtQE5HlT
ofPaCQ7+ghTKXuh9X33XERz7btlAfQMS7FXSyQdJinL6J2zTNvmA6OiPMbeR
RIlxEdaFzYiSTgiySjVFLlEiCRc1F2qCZMUOlqIgULEqh966oPDvsgNzeP5U
qA66+tvDQx8FTYW/csraj9bVBkzo7OBj9XZEBcTa9teYUxcc6YyMRR6RUato
gsZZTHag7QS4tXr+IuZdeWPS5SF+67RYBkGv8e4cW3qEIg0CJVrTObbsZM7F
XSooOR1XAjGMlrnV/AUIrh5d5EN91NhgPMnt0gT+HQ8b+iVWgGiyeGY6HAne
iUtvWc9XcocpbTOj6elVbkhbb3/uDapuu78RPmlL8yAuLV5Vv4wdhUJox/Oz
y4BiZiVl5IgZkV43/811QPI0MOc6vhfgby26EuyPQYkayqe7K82Z5UvIdO0/
blW87o/HO+xbOYed15sbtoQAmnBwC4tApj73z5U44HTltIVWpdSXNMTRhzI+
6F9U/qWZnYEYeGT++D6xFvvPqrzstVaX96ifOA8K25ELIta3GSIEPtBaNPc3
3sWDnoqVhlKLYBC//J3j5FJUcD8MJ6dKD2xhaRwwdJbt0G8w+lp6YZ++2ci0
ikJMt2acY0RuqCoxxtgkqciY9hr3E0zjQVKixP5IRcn2inTWgi+a2rqqfHd9
K09OtDU9dEw5KRomkqxUMbrTzgztnN4j7FtXFXTbK8ALTOJS6QO8UarIwbji
3xhG+dchTSqroLZzuON4Pn6jMok7tKLZpm252tgj7rXC9NgOgAp1Ne5lqEtL
h01g2zJ+tOroBGalVA2sJ/kRLVNzKSnGUdN9G7dqY8OQe4plbUdUPV3MwhCl
pfHvjpYUlWtGJYwbXbaL8TYh66oVBFOIUBXKAXdMFns5ne4gdLXPX5uxI8rw
ugL2WUyl03WUOPMHcYgBkpIMLwxut69ChTYvxo0L5iSycaGSRPSajqjSbhAF
Vx36E+EkIyK+/8u2F7Nv+rJgyfSS3mIxwSoaKN8DEhBDUv5HZkw7pBQVqdFe
nYnuG+tWCOFqBfPLjgKuVBcyWKNvw+1MuTQtuIqKbLGNIwrKJ5bO8Z/rmiJy
kb8rOSvjhdUi+wf0gYY/b+Ic3GR+NbqPiKB5IGNpNpVWsQwZBEmGKQmf1EeF
1P7uvu1hUFAuW8IP1yduV0WQoR4XJXLzJ7GZm/8efhGClLKOKRtQezXmC3US
JDYyf1GbYtAVleHaWHzV2dttDrrOVnxX1vFGs4+AQ6275VbqDTcsCSpT53B4
okT/DXk/zMFHq3f5e+XnzjMq9e/q52icuQst2jJZ8/zoDKcPirssMdyRlaoz
4V7bloOycZrPPFcZOV6eO/SBgbqJzMyp+1+PcDX/7RKcbqc7qxV98tJldD0d
l2xLkhFn989XQGSegjCr5nBoqdH1Uo6gj0RADAscWwLxiS3IYrLbByuWJRnL
Tqg9k0TT7aSQnYjDP6jl9tClHjB5vZKfZH/+QVtw3i0/XCnBQyP3cc8dxHYL
UYxLbC5curJGRLm5CZHAMycnVCAJn51ruPa+UfwFwstkwbVlBR8BOOOJWo3e
oj9mgL2OkYB+UWZ4CrY16aHn4EtJwZvm8QKPjlumF8NStl7LYaAZOKDmEj/Q
J0IZYWubDywO9jD4Pbf5QjsZqnSypCkhRQgy9gFVbmduOMWvhkAMrO6Iz0oa
3VNK8WzpPB3wEGMUkUbzxZkjruBxCwxTzTHAVVqGGfB75r4SxuGqH+EmOybP
DGa8qUN/BWfePoa3ChKvpSgyhMnvRS0y1u6o6gow5QmHjS5xsbcn7HBqwCXT
Skch+7ANwTihTk0Xfubh7C+yvkMJAePZnlkqcE2kcBYAyMRD+1dXOVZLhaBV
gJ1LuZBj6wtx9jPOk0+ExBZfV5uryS4kWWxRnyStbqT/orGL2KwPtz4uxDn2
61wocWlp/DbPEIy03J07ksJ04d3IHV4ZRcxoQbbrkTnjRE2D2Ukjr4lKtPjo
eSzt66b9+H9PCaL25sn/RIoROuNF7rvDY7OVAR8S4eTjZ9mN76ldiI/E7LYU
/9O3yxDT5YYRTeu0DXifwq1ktAXLeNImpRFnwz264uvXm1gZz7c2uV53n1uj
HXJi7ZphtPamz8Fq4R9pkFwYFo3UOdYuZqqRmWbnrU+CAlIfdATd/zHhCcPQ
aF83BL7QyK4ncArvdFRsUePPX+uNSOUSg/RlxH2a6njE/blMkG4dVNfwK0oA
IqV4OQ7WemJqyKwcJ9HdsEiEi9HFJoaGAT9/N5HDacpO2ZjNDGs/0wiVeluL
UP88kzHsvuIwgvJjPgV4pbqGMMvTKBzEEjiKhThlWiwhgSFlTfj7rU2fd8Bi
E9alNmO024rzC/eLMlfLjIItsWnJaX3MKbuxNlL9CPZDKugUvfwe6nTZ8I9k
asg/Zi6vD997LMGts31ToGgc+/+Z24TiTdPJ4Rvz8+Gs/3eXM13D/OiXijPz
JbWMSPGzu79XeFxe+u5cuNOBfe/p2/3wC8nj/5cjHycS29PNfoXvPansOVM6
hVQ4hmgIhMzYDacWDTaugtOA8fJqcBNkWwcjuxe7g1TaYwz0hygYTtqKUMsR
KabSQtN7n/WRzRiDJyAStr7xuYnw3MPkzz4sxWQoAyiFqr3AUgm9XV6xq5YF
rGglRUViGOvStlqO9ysW+HxvNgV8KZuWCyL6DWRJS0BaKT9MoZx9fv8yBF0z
7lifNZ0ovST6LpFLVeoaPPl+SFu2JAyIUVYilNeVbCoWzS2kEUuxhw2lB5xA
LVacSLhYd2xX/SiZ29elSMajmhBmvGy2CQb/kHDTRXN3N4S1Mzv2XvL9PsCE
67MS+7Kp3djLUWefnRj9bLTnu0Wc0nbpeR++2kyGWwKDXwS6yG6GX++RApys
jLzHNekV0fmkxeitz/2EqXnsumV6fuMqVdAv0RzOyRSD2G7ueQ8GSAAaHNuS
c4ks3ppNIKbE0b23pfEZ3GZTTVryakP6viyyR2Hign7LPE5CrITUHlU55NUh
POAKRwyMTKImIUCS6SG6YNSLXB5NhikKduy4NFvXfDtDv2U9O3U7ZdYOksb+
fyNQUMVoeNu+4lbdy1KDgUcL7u9krG9z1zn3Y0H0/UMjqa+r5IQClcKYp1CZ
kBib9v4qP1t7hfVv8AYtpE/KcvoKTz6LGmZp/3ZRnaFyvRpe7k9uaso+g2XH
mmjkdJgZthXKMmmOwPmoTvKI0NIIep6sM3Yb0xeVqn9ehbZZIndUiD0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJfRn1ssieXjQdYzAE4fI1yiku9x7EJjs5MtJBJZqIJvK8BBsQLvYk7DmHGLdro6V/lV0gehkOoTCT1ixh/QR13tGRr0bHfKakYtq2Af2A1+DR9rUaDyJqGSfXq9eL6UEEPaehtFWhDfAAks1fAcm+Lvf5zDR6X4vUaVAMOUxCTAdoPkwUxc4BTj/fpDSYijQEC9afKJ8LTs86ETc/6CtVXAddqDnL9TKqXu6WetlZd1DAKvmpK72ULd4PtMqF9Y+C6hxW4EEui8za5LizKP/v6zJ8kluEKPd9KPXzC4cFmJmhRsICcCNEL8a/Josmoj3xojttZKjj/9FPLwTppENu1sgO8RkHTycQaEnt2LZk2aADHTXR0ua2VKwWGOfkmzDkhj8ZxKnB4LYVqLr+1qjcFCqFVh276HvOLVsnRJu147A/xHLV89PlqOc4KGMW8FPXIWYcKEWHmAJNPjm1H0tGSiJCCmRq7kSnGanvyL1t8r4m4EX6bpwMzqImsdRdUZe7qaU/vYNmG1OcLx6Wv2oWfWzSlAie0uzHm3oqV8E9mTOOQwp/6YSHcgWi+cMXG1yxX+fYsR4u4LZf5a665ChHbYIL021rB1pQpXAMbT2jfagEXkOoNXs1yXNxNaS2lyp66p0MYTl5dlpOfdefMgbLt1fLVeqKg0We3bSPijj2nKH96jYfg8sHfXvFzT3J8NrKNvw1msWyFzjHC9hEgRfaDzuVQPB2mErb6vzx6sXYALa7mPygaEvgk7+G8+14/a5V6OFHCwON5nAAiPycsu77/"
`endif