// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FTvnPpZawdQWDyG37pSYebImpbV04TCs4v0IFNLGSEuou2Ya8GFvgmrMtSFL
c+JhbgAzVVnC3WtL87KtBtEx98cdhgWfUSyVZYyhVXDq3jE6h74T8YCGg91Q
5OwIb5MkfiMn/B4BMAlP7x4lHK/5j7g8QWl6nC67Rurs2CppIDUQ/LhOrwTA
qwlRomjjbqXcElwpgoBMkHNvraMPz0ot2dK9Cd3S3xBlJaJGuojz/WzWxr8c
plVOA7FD5fy7YJcqeCZvZbGUB5x0i5C42ndK/pL7HS9gFSjJdD2ThSedZZBJ
jdCOoKxBwzvXtYvP5Yxi5dhke/WzMwvn2CgAvlXBmg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WaouItsSmXWo1pwgsTB73jvDDv9BCzCgdS6FEirQQsRPpvdbmmY0qFAtG+mN
Y3HZrvUfnqjhOCBz3GRqtyOXtEvgvEgMDTg7QG+jYpNqHIlSUE2//l7bp9m1
gvXu5tW1h5GajvjQjcZSlNA3A4tAkYRKhsMiMTr/iSctUJxAPjP2nUhaZf3T
iAUw3HP7+R9fthFd+k/T+lO771RKh5wmoWKnO4irNVGbhNjm+CpyIAwYIVUJ
cN15nqo9AoDt4woNvHqn1MqOeYQX1BBGq97YInx0y+QNL5ZKYFPWPCc/T4ei
TEwTwh+ATRmdCRq3psDqyN1kXtZ0dOBR8kXRVZFLgg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GdzC4HgP+awGM8NqSBTwh7XazgdkECQOhWE7PUvwvk2R+wfyM5/53BtTIvHh
rQNpc/+mMKLth+pmLdtdfoCPiZPXXy4PqPYiODiBAX0Isfw0wTkEhyWkuEw2
kMOfj4uzp1Q9BIOjiu2SZ6cmViZrkqyqhL80ulERZj+uekHke07wx6phG6+H
KBBxMr3jJa1pegcm31FiW8+3dZFzRKa/MAbsv/fi4hPiNdJpNDaTTOfi9Km0
y55oMlFYC0WG8n4gMDhxeB72X9RNqSf5XgT/pGkcJyJWSKSbmw8AcInYpufh
c+2uFwjwdOIeSWKB6H2C4B/TjJNN8pKK4UsYg4Llhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A+K2JGnqL0cO2cBpe1yWbvV0ZTh9IkGEbil2np+p0Kuq6yga/KA4b9vuoQXN
zY0LaI2uecOWZ6iwl/W4i57rHV+lqm54s+sAAzxaB6Ts+FvtAXD2doPdD4WD
kGWM2M+2dc82nC4KqS84r8Fcwvs6WGstnqdh2f2ZMyhOiBnYH481aNG1Jzkp
D3vIUQjdBkRgMj0IBmgmc4TXmCcIJCfqNT2QdJK3vZGN3SUCwV5SghukU106
+2pC/xbJUhtKFafbMsoOJ+98F2VJGSZlFI4YM+Wa2FGbg17NVIpgKIz4D5ix
sWKEdIQ6XJwLkeE7Pq0YIaOVuPkPVK/oOmEnIEZt4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MpQ6V3unpg5NkKTS9aatREAwhKeoCmmw7RNUd3vbT3KPL8xBDOF55A8SPFy0
OCMLdHZEkFmKK28kPZqzo0eVtW/yzYe0YwQKM2XgcptqC8TUleRqqF1SjXYv
RSt7tgtGGuyd4Uf1hLKfaZqMYTuoHkiyagNdyfzvOtv++1iIO9A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gF5sE3+McVfNU0RshgvJ9XXrgnIK5AniX9ImSuGmt7hyle0Ag5up7ByDrLCE
neyljkERdRvqrUETJ/sh8IpcWLmXhJqGfMmQ/Iz7kvce6KHhXO9PvVJ3jNP3
dgRmbOdTCor//+blPaRcC0v5UyBD7XNP2XcfmxR8VJ2boywiphh2QVvMX3Yy
98TbtzixVcABPy/cD0GbbiYK9buAluaoq40nhPPupeLnxwd4J82KMX74hHgy
xSupyhe1bkpBoewOpQHlWljoKOrQJqLN+3f093cLSt/nxb2kpKD+WO+BMksU
sYitj+ltRNK/TgR9Ks/Sr5slZIiruhTgBFXCziC2C7dH3LImscKVEl1ewZC2
iRTw3r03TtUTt06FwcA4PcTYjPwI2lRYVevN1hwx/ugzugSk4kodDBGhNT21
Z5v6lcd2vvqNMt8piTmVY9ATGcD1XmRgLvmaLm3oaW1zsD9z8FQx32bFuyUL
+1Z36dWIGQOgkFrhpHYVhFc0n50IgzMh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QRYY8pSxwZ7dyDctvOdHpiKxGZPDPc9fYJyGtTLWSJSu0CPtFPoCmZy/6UE2
nLSMVFlFPYNdIMNfL4EefMZ9PfaradckoYbf6wiHyLWL/1w6e5sNcgCIJWUR
HsIXBk9ukr8Qv745HPIVs2mkU4RfJdaTHqYR43FvRd/rJaBz2H8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dzCXN+qHRW9T7pzGS6ZZLZlvTg8RkHWpylqda9Woh9TCynU25l1A6qRFc7cT
gIaGYgnYYe3Oq+kMhkho/Dkxk+eWOmiDOL3kBANLCMheNh8jJWDfVGH+U0nf
86JinQi2napWXcOE2m+blckzfveoQ+ZfAArd9LL/jOueux+sINw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16704)
`pragma protect data_block
y/4A+Up8ZLI1p3OyvQY/qMZYRX+d5UtvQSagwIbamIeRgJ0PfseFdp276IWf
sVJImntBitlus3Gs3Kos3NvtK4rYTUeU3Rr8zSWbr0oeMWWIfWsoxSuEyEm3
M0DktK11fBKiKO9eA4bZLjx5zlChv48oDBM5Uh3A8/X59Ua7EhV5LeL/1xwu
VYt3xiYTjYnMWbz5xqAJMPB2F/4qJSM8wN5opwkF2rjKb3HpyEWYvK/BVzg3
2AzeXe7XctW+BChCPXM7eRZPs00+N+3SVfR4PRnUh6sjYygkU7+uYz7esDat
6xYE2eKV7XjYpw/HK9xYG8sEs3B84LtMGQvpeQfs0+fKSOluSedJaXqcZ6FT
sdctIrGupTd4BrFzkn1dzfC20nhj+qyGt+bsmS6dXfW6lQPEcu3Mlr33/3Qt
2a4yNyhKmZc0sX65+02OQZJHenpI5V5rBEfhyZzZiO9yoSPB2wlqcq+G0wLT
a1dhlQ5d/sh+4K2CzfOlI4OKVwvgQ7Cj5hcg0WV2MYouWGzb6rfpoN5R7DNV
YKkJFk0sgI6NpFQbMoBakexUe8Celn2REzlG6Aa+eC/1MQfDdv6BsGlJooE1
RIpy64R8VFujolqX2yABP4GERMxQBkar090qOQSMOUGYWG7eTElqkXWzpr2Y
GW09V179EVO2MbpQNhc9krQ336rr3/1emLGgGEN37JcmmdavQ0YvjCNd5SIz
ciA/54G5W0JoBKxdad4satsheEX6gBgIk/5uZObgUxT29vKEe9YULglcvJUK
+kV/HYaypcrcyjeQ7ur1r2rZBKkKQVpP8lAV6osDQLXjb0/3WL8hO9xDN9D0
O4ku4OcfcuH9jRry48YTVuAg4O4h2v7wBpEozvovMKDdXdz0eiMc8VEMc0V9
u/3fenBGgH/l+DODaXoH3azmkRYwIj6l4Vuy/JdYHLIUyZnzTgeY/BIpLI5y
GBrn2HGzn5V5awsQlC6OO9NT07OAi8p6Ylra/yrjYguaT6Nl3ZAkOXCKqvR9
dw0ze+ulpWTU31+vV6tvo+t6snkCsVKr2j1TyuH96QiTsdlSKsFuwA5x3w/D
H/J1GszvzHp0TDwvBTtbutnkZHPiL4dgFUh2g+UlwZVE8bY8FHSOBxdqdTPx
X62WnC5MGS/8xnwA71CPdCzkoHSjfn6y6DEe37Im4ObvYrk7SbOrlt/I7yoy
HTZS5cLnjYi1wxm8cq7J+J3NpvUenObKAvEWHcMHtY/Ij71Lct2ALXqKdS4o
0QZUvRtXFZ3a3dxrc10vFpPxxZQZSHHyW930ebq9z5kq17CCuAVFwLeSoJFt
qYHLYPp9ibWXeTNwfzgmVYmRaorRb8GXM6KqwRq/HEzkwx7swmbv3x+O0SUh
WJFdsStdg3Zrx784R2hrQGJlfESVhGz/HUOHLmNm2HEPyk/zwNntnqqU7n88
o4K/HWRlBETUzTv1eg98yLudyvSMqX788a4QoZ1PtPMFIuMjELdNILg5wqVu
WjZFTm5r/ZWaBt5Wcw1PZkCwHn7jyMqLqIqrI9S6WB4EyLwUCbGwuPtEwl+k
L9NiYXKivnKK9N4L6sZS/DcZzdjpne7LPzBFYYz/VgC+tTXuLVhMSIzLNaBQ
QvrHP6HoNAti9mylgqHSmo8ElkkDdlEZYWDxwqG1Tt45vkUPOEB/LICFecuz
KImxaK5CBoTp8Yd5cW8j4oVYF3upQ3lGHIDYXFiDl9eYMPnDW1cnPNt+3yvm
/mUplB+PW3ZMa3LxAAPx4NPAS1nOzPQMwhS5usRsYmqRcDFwxPadGF3BFpKt
G84GH74PCnF2U/ynRL50f6ZolKorNu6VYbbVssmyV9SRM2QvwOxRziotafdx
awu2xZndMEgzEEAhPG9TUTKisH2jSG+RoRwYuy3mtSXGPk6Wuv2cwoJvoFnq
BdGaks7lEo7uYJebXgnPsVKbZkdkg/9dlmOR0ZWx3ScklqM/Fg6/ZSzHG/3e
Zb1nOhY5imfoZQFRkLu5HUlfl1FEjzK0NoqPwLClj/miJ/wDl4jB7vYoaHPY
9iSxzcfmotONuBtpqGnT6dV/XkCscfHVHX3Pui1qvUAsZyCOGG7YWHTKtduM
5dlnAQbY0Aq3Uw58bPgbWe3GKA8akVRkVYVB/EwjNsGUd22RjAhJMvImA1Gc
mzpUa+i3MVAi36qAJ06hmHeedsrXAjuJ8Hzvb27n8AcnrlqNgUXJ7WSd3iWq
QuPXC7QVe39cl2CIgboLnIS6ZPzoK30WW5QPUxdGGA1dc/4SVoUltiLpiDWY
TD46sySJLLT7IZFgR/xrJBoAmZ6tUjgmfyB8bB+/gDHzsOSvom55AYFzs2Je
Xsf3ziG4W/2VPZcnx9QRPgA5UTtsFAkwoweGH0BzGdG4ETwckqCmmj3/2PUf
DR8WUbEVcE6gntSQTrkd+HNWAaGOTKRTgZVzTPaLpVvKeVliTSd6clPw278N
5XbTXF2jzqFCfQIblPCVipQ3ofKQAHjlONKIol8d/RBgsKxDLYuBmlo2hv2g
9LwzkRErRk7GLp78dOTDb4AxsI/hnrr4TCIr9froiCgroLUAZ/S4LAkVoiVc
VOuCvjlAg/91pQp/5qghA0rZRjWbMTJuK8dV7SvBrBa81A3mRqcQdydhcvlV
zaYz/9nuNU+iAC9DFXs93D9VcOQvATL6U9s2dwUg49T4DBDGLopsRKa98rMp
sqnIiML/BcxWLMyoSuQioFk0lRJDQinVfx2zp49939BHcpP1jO6q/a4cp1L5
icl2DRv7I2tj/+6syoQc8F8TuhUhf1PiKw1BKwC4pa78ssBHcYXgKnsooJ8Q
Oh6V5PPZ9VfQYFbc+kSn2JYjkejUQD16kY570MB9opTnK8XmCz+LxGP1gAV9
GF5dfRApmAg+Bdq9nDVFFovRYMG/qzM4z2zZfJ74BdGr7sDvRB602ClVy6zt
TWWADGEVBhPg/1VmsdndeZBH0S60fdfZ2ozaF4mZ76354PIMJ1BbuMExe0dq
cb+ym6DVkMRZHha9Qo/0lKLTg6Z+C2y1savGI0ESQChcJKBOhBw9EgtoWENB
+NkeWov02Yn8VLuadGkB8HSgppZb4dT5uZHyVxjtZfFiL5q00vQJp7j9SAVM
g7LO+iuUHwLBfnpcueo3gNlcAhDTF4xrhwXuOw8BiTPYLwdrz1vKCK+yiqEH
jmB2ErMg0IeRr2wM7brXXUfqWx4sqkSSWB5KzlKiF3Hh6/rIuDDuYGBn91w2
diOeRIEnDOjHH8MhY+PKINy7TcAeeYeLBMF9/3Y+6WoY6XSj9ZQEqWnAsmZ3
l7/GOBDSOfOXOjH+FK333yoICm4rVz+Q3dcUNHFSHdU3Epj7EmZGmEnADRJy
tSb2M45/PuMveB5Ac0ACTxMd5Wk8nQm3RLPr6KIgspWs4LZdBAbWqxQKtRh8
HOEFVyOcx9kdFqrOJBNKSW8V8eMBXuLI671uNVh8unzgLnqhloiqFLQxf9Vf
8mBSQ/QBkyTg/efDxBrfAqVomiXQqAye8lgh5VJXFl7MNxB39e5V+e6wjvPD
RozV23IshLKU6dEbLqBR2DuPrSeWNhdLbcZA10zwTvVbEnHPeE0wENUREoBr
gxUveJ9d1x+T35mp524HuBlruIkpcaRoPsIs8EOTh+/vvMMHawjf5dTWYjFi
v/NgssqmuNr7O805gSrWoifRNOzEzYtrsSkSEvQ9h/PHP1B1TMGwR+MFkcBD
p7P4rHISkuDCequjOzTsHylQ2t4fwqjEb+vOL0PeqzOWE4gU7YMQEUmDFjrB
HK/yl5KjHblMKK0okZjSkKMSoKNgW2M4ka9QbLpW1rC0s9l3TqhTJAxXOOYX
uCaJA3d38UQOQIJtIRnrgFUp9J4LqFUJEJN7skze1oXn9NPCrQ8MKH3phiEQ
aWub9qhiiX8Hr5b0cKQzXSQrRiIFHg5thWk1zB5rbAFIFPADecjtkLMpGH/e
7LyhxYAtVXuMOtacCY0vsK5XmlrOSui1W8L4ZL4L4nJHvTRW8k1WGVqyMUHp
IiSJbgKIYvs19MGFZj07lPm6k0jyrRk8hAUr6LuzbNY5N9VVm1dYpDMmNRBS
8y991trhw3JhXGwt2mjb8XsVp3A868g9ITAgoduIsY58WTRbi9G7c2sVnUsb
MUyiTEqGW/heQnjUmFXjNHSpa5kg/LeR8RXbUhsklwnhoJwPr+XXGDTFdzlR
wvlOVjZWw9iuCOmTmCvQdZY/fbfFqPm+/4ztp3k1oH8bNa6WguDS0iG4N4gt
LRjSjiHnFJRQTdi30Y14TllK88fPUmietyIJ+ULXkQL2Q7+qa0wn+5TDRUQu
VmthABGFh06hmLu9CVBBoqP9QEIxPs6M/pTA7hLSO3VyRVYgoukBWWSXYT01
JTm2IpeANLtPBVxiL3I2Kr2IqRx9jWt2zx9iXpTBGeAc2FswVLh5FKsMydZ7
NI5J8l953pSRSbkReSwHI6WxtzhjjTbUiqYn1aLi82KXdnialOOMp9m3p7u9
mprxvZp6ZGnV54ECEekdV5AJYYruP4G/401+AYYxz4Wjk8NZ+oKbxp625+k0
lfiVIY27zLWAf24+UwMS/4oe9oEcisWAZDOSU0dVQhwukFa21HsNQA6+ZRt3
MO32vgh+Hgak+2AVa3s9AU1E3nSSnW/HGeKiC+HidjV6FnIfxEMxDc/o7BWL
txsrZu/EhbUOCYymWarD+JFNSNRSBDL2KZpVWC2Fy/10pg0MMECf3tPk0Svp
KAvgPMHLxNQipgjo1y3v4PPWTihSBrn5OShZroTLAEB3XUvJ1sTgQE/16Ytn
/N96S9MQ7mzDXy1oSkhtuG+maa12oPAFXcuUm6X5P1phyktGuaMg/41/5VzO
9QYplRslToDM8tdsMIwErMkb1gaQ3oIoTeIW7VygU5NHBuSxeOeShakkjn4S
1QxAKPl1N6wONND1APOEaze0v0mtVNw6tTgdkSRBn9D5pWTzSArhl0dJpK6o
HDhRnnumCZklroLTKq4rk2Rv7UA7s4pvAICB6k8gw+EO14BGzFmeWxI3vdWY
X0Tpb3YxTR/I+SdZK8IZTfD5g4huG2E6T402c1NMR85wjz3yE5gaDcqdXekX
9EiYwYXGeH+E08FSn4FsEURe/Y0OVF4C882b8lz+17+wBT4iOVBWiss8BSiZ
e9fkKNYQyWkleZIqcYssRq4PYgO3yQoAIy9hQ7uzHoWFE1sm+Gz6S/ei+Zrr
N1qWi8NYVWxdMtZ/lqT8D+les0pRct618q2r1VvrQPQRTXmRDU2ZQXDhJOfB
RYkxqnN2WTqndHakjyDJUtsM67TU2kv5cQ1PVAvA0CF5wVFbx7FU5pqvyNpQ
sEfwXv5xRrkoUl0n+K8vZv6Sti5XlQ/0xx5Chwky9M8D51kxKLeWYV40F/p8
Jsn0Ss7ITpkU7aShqolO6xR+QpSda/kpqorj6Yx9DUYhN9qKbFL69fAYEFoM
eC72SD11BOw0q5gqIg2Bf/FbXt5PHhdtPe58RaleVS/rGh1opEZk5zTQJLcf
FsRDelz9HhtCbZoKtVX4cIVpGrTi9iBYRmTY9hHjVZSXF69FIEzji1H12/5h
hlw6vVnO3+DuH8bhQ6cYs9ogyOke49MzpNdwKF0prDNmHyHI6RsxHFzBwp/L
KRGHI173XB99HHpMXRWiV2ArK0sMs+/70SvRgU5dsb8oVFmgDwPmCULo8vV2
MVbGqL2yjp3ELIQYNXdGxRn2I3kW7khSmA4TmXKj7gbbzd1rqCetU4UuB40f
IazFmGZtf1zvpX9dQlJcx28kOsE38YyR0ni2ajLJQDLUeIgpXcJ4UJKSWQSX
tXLAmPsR9F6EJ9dItx40iuT5YLSj+6GGEgDfDpbuLPeCqTsCJFuRyLkIJMiy
7BXLrTRe/9j4heVncdpzf01yCa/z75CsCG33k1A4KHHfl0P1/OTfpZcn0RFp
laKQpFAiVVFNCBre1ntTTZuIGMTNNVvV6eRl60nijXojvT7st4SZw09St5U6
ECoq1ATIpxu+6RyK7Nvs40decTfsMjLZSuGw+SZJUEJ9zRhL+t2ZLvVEDTbQ
DXBfYpHdEcQI7XIpBBsrkmRVcBEBmQX+h0hVGXgQukYjyyBXaDjPVF3ImsM6
noc03J8zoZOtLuXMPeCI+5znQi3AGLP8FkByWqU5B9NNfyLOPwAdkQih+zU9
VuH+LiNzfGY+9QZn0BNrY+1GMMfnnn2EzH3yDhjPmW5ESYqD2WnC5cR0nkkW
2ZjSNVEHVMn+LOtBL8DARq6eYy9Fp8pYxztWw4fhR9cE5Qvu4ZjXIBVospVq
mLGilOznb0SMAZ4tQ8rufm4iyViN8Res9BwTUrsPCfj0tbyZhWHyllo/Hy2w
BqBVrRVj6hCtYITjnxMWpstdXoXm7c7YscMQYPxkaEezmoY1Kgp8jkeGLI5D
eWeLTocIRGJsEEDrD2WsssebR9+wnEVJDcsapsMStRcgktl6I8CDkraeg3oj
PI08FMJOJR99KWrkJ22P2YRNIRnXNEeU0bnITqbV66OU0BZmiUmO2hpnRp35
heGBl4BjAflpnW/AmzGfXpQ8uHOWVlpz5aiMhwnvP04e+tG1L7FDVjS7pWA1
3OacAEUmMf4dKhgcKay5aE6BUipP7zWrGoJf0tjD4Eo4T1dstJFoFxj+nR43
c4WyyE78l+SVcjSgtoXDtxffR1rDH0AhXs8Qwjv0FSE0PHx94FbHEFRmLfrr
s5WX4vpZASK5qigSrLI7asfbf+hOnLTTm5GSBGPsa7edt3AaFRg8RZcvbVB6
He9VxEJVh207YkkkmTWVkYo9Hk1h0Id1SHKZWfpDv3v3TpOagRNMqH7xl2KR
VRLFChXZ4nMFwGay6kK31ndoRdSH2ZOLOKPNSkBzBgbOHylatEhRTkDhAeMV
7HsbkGaochRkSUtDMCskaG0v8+NiYcVMqvu4Lmro5z9YwlOZzjZQBG+KEOP2
V0wHt8xhYYCmL14W3y/nXKYlK3GEXGzmHRbLEoWlqWOBkvcDSPOXjBG/P8Q7
tjJlG1JjEubgYviwZo6AU2euhxtJDVRbFy4ZiatgLHzlsaFwuW54g1mMCyw7
08nMAE82Rfqq0whKGMXEWTyVJ9GRVETByVEV6kF7AUhZTC9/Tsx5vhiCE01Y
vIW0nBCC4bvitx/SgM8isNFJMsZn9jANkjnQG0yHMiBUac6z2WSjvSAkRDIM
RmGJvvRKiD93MoquYhNCwCyrxA98DgFQMjVDfguS9VlcM6bS+3B2CAxjAATm
4lbChWSBWeRy2rMhwCgtNbZoNMP8GrKB5dCaI9qdMsvHt80tzL+yIDX6ea2o
QwSqLTp52df7RI/SJTyddlW1znErPIDPbyATun/GXkhmmLpiIfRZ6THFPlW7
8RP0JGz0Wi/qwsHUUv3pMIBsnbszuvhPn8Cnkv03zEQ/AClop5qK4oGrlJOa
hgxReLyNUlX60SbnwQl7pyvoHKr93MsKpTjqljo+iwbTLUE7HfF8yWVG5NTX
PvQ3aqTbJaJIEFuPm+VOWdpgy3nxs6OQtnTCvl1GZRmBEDnJoFboPqefIz7W
dmKurryhed5uQYhRnXYVBrfZbnP7OisEuV1gwrqkHi4TF0KB+BlnkeNmb3s7
W7g1GK6RPQ6r9ZSiqBExHhxqbuRcUBD5eCq5tUyvGTrMbweConEEUCOTRubM
EAFeZBVQCAqGnvgWT9HqcEXCt3nYIYsR7ic8Z7FdGYlCRG3Lrwozpox8lLHC
cJIaFYImNmPqvbrksrFtQbUMGvLrPS1RmBm8Tfr5aVw+rA8bGYUZOAUpkA8L
m8okj4/BlfxU9TqkDALDihsMsILrdjIrqcNsavSfatiO6dFHS/DcFF6qPS7j
Ltffbh2QmkoFz/bvUk+m7IoDtGInzml12qsDEcEcJIEsrmzT1Bi22Wh5akBs
MOOEcKMJ2FnHyvCl+YxuU3Az15T8fhLgbUxvCD6P/fLPHqqKBdNlGyJUc2WL
NVuhzTs7rayZzpVzO3gpu8fo4O/9FU3bbLvbcVyVXEXbaaWaCAIzD6AEEmWH
2KeWXl1/JQ1rnJLDnXsagkRTzrdaancitePCYqg8yuPFklSSATxr8U2Ugi8G
Is6SGTvSEV2RZhqtj/2wrQ+VWfeGQn0o9Y/wVIv4+B797b8HuS4YLKGYzBM0
I+mOwMwKft41YJtVPzNCKhB7XTU3nECvRw7GHAGn+MooipznEcuOcwZmbvO5
zyzhqbv3tnr8obCQwaooyAnTdxWjTppJt+8u9GktMuIGkfvOiGxFpZJmFIU1
BHT/Xx/o0sAwKXU7vWeHHV17DkEjxsC/NloyREQLBNcSJaRYAO9K4t2S5V2S
Ko6Q15N6l0UlhGYONZGs5EkAIUkt7YIg5jIQtbHcLCAn6r6hqZers+JaxJH+
Kc/fluUaU59Z6S/1vWTpUPU2n11BSGi0KuTS4ta62n9UDgOBo/w/FuOwxme9
TqYvIF32Cw8dbISm6SPHLg4oAifrZwggo1LB9UH2kyBX8wZogsv8r2vgoPU8
u+F2397R8nZdgP2FBvy1qZyTzWeF7O1WvFoV19yMt9JZEqoDpNa/92bLFmkn
baf3UelxFU/UgYoMDhn/5GBlIlcRENI8oSWJ0AlnJUoMtsr9wK41qs1CvjDh
OLpQ74bEf9OB1ut8xLMnpyZlW1NVqvM9WwLQfyajEIT+HfysS7dEejwSdBmQ
ct2ivYQgkctAYX4BF4purRf1HLnes/CXAhM6SFSuRfRKE1m394szUSX6aXqo
FpWUFaqpqxBDVel1clxJDy784AuRWPBrFlbutcpapXd93Pf8Nq69boSSth+k
5FAgJh022XwescnaziPXpquB4W4mPFHH9OUJbNh+F3wJ6QfTasNT3h8xuxFM
efuuYrhIAguIATgKBHCjIEqR2oDCEMledFAtKRO0dhl3yn+m8slfQzsmayfC
LqHWy+5PC618LiLDnCOkAAFyGfgYtFe2vJwRHNvssTCzBvbvN99kyUyiVkK0
q6iXi6AegXAyYQWscJg0dE1NB2PmR/JaLKQ2YaiU/nWiBHxErblB+HbD9RQz
BSdrHzkxA4HwWOJ1OUG1zddfYZNXSynLxFXNSPG0Qwgs/XdvOwRRDW/ridfw
ae5jl1Q36xmHIZnTaN4ZCOTdc+6C3s4NyhCNPOE7PhU5MI19gTiALOrBdv1f
amthA73NjojLlnkDO72QzPWvq/IEA8Q0HZf4fNUGpEFqahest9Cb64eWJMrm
FNXFQRFHl65KsrbT+v6BVSmENZgB2DyzPmOKiG9xZhBCbjkJ+v7LOK93dkmD
xTwbdSps7QKEFUiGDBwVyMSXbTg4tlrBe57Sc8mXeMLv6q4QVipb0saPzmNj
NhmycaKQjrGKw7+lI2l18EPnnEhFcGBMAShaf6T2H8QFf8fsnMG9ojjU3tuh
aoG+0dmxzsJJDF0Zcok+ClWmAGJa3JgUsCAuiCleAmm+UTbv4+ndnXMzQaxm
fPtO8Qkch2HZp2fYv/a4ykqvbzVDwMVu0tEYzGG4j/5qCqDwOav/qtJMjOE8
gis9vgo0VQQwgnuh+/A8srSC0UM86Yihbo1LSzZZDrjbSgrYhDZGJBBKi37x
wND+ADCLOJ1K0Yez0EiVfBWEse/nbkj2VIWdQpnWIP8H+f8WMtFEuG3u9Yvk
YzqmoBQegwouAMc51IHa/Qrl/GMUG4ZRIIWfGaaycZ5qiy7h3cax5HYFGmlz
CVNrf18Lp+dEoEVWZBrDP0MEd8eFAuux7HkeqZin9sX5dpDQu5zfqVGVTrpw
RjFBLOvip+XfKZC9b51qw5GdfNvf68+xsP5IFyNzOaJAs1jshdsU4OcSB3O7
2FrJkx8KGrdrnqmki8zUcKv7jsIS18Cs6CAG7XpvmFk/K0ZVUqZ2Km2AxwWs
NbH9jW/iURR5UZNvy8JtKRHGq7/qSR0iJ8o6DpOLIasxu8TOP12vF2/zebfR
YI9nuGwoPGa4RMqqfBSltuqETT8Ezwq9ZN5SIrfUfygcbteUCOka5qf3Qmfo
EfyeJEC0LJaFM9VlaNtyYp8MZCFHwl+J9rJZOeR/mPiCi1WAcYBRgwsaFu5h
TfWB2iwkR2JvFwMNh9SMuFWRtMZzcFktS1onrAxHTumDOBWRCn/zeBGv/jt+
q4jBPrzfN3ujSuAGn0NUJsV53NawBKusiwoAOLRg5q00aqSc2HpliARPElOt
Z6062/qR5aEbG7vtnse7TMLVs0A8wrbzwADiiyrwbePz8U4gYsrIJmwG7etT
uclOwXdCH8tRsSFzPOozQRDevOBmeiFin1ocOuu6ZafiVOqR8qYCkj5OjtXo
TFEXjPlBlyVLinxzEAbz+ogtqshVgCHKfAvpGZ0dbd5ZhGnSSK6H+zGG1BoS
lW/ihMyJwWoBDZlNWQYUksIooL+OCawKi+yZqEFokL6UlE0Q0FIR7W9h5Y6S
IPBaGOoZKqmAXdJXUcQb13vDe2zsbF2Es1EWdLmqM/csc87V3+SytEEdjVzO
pCRwlIxkk8MR40fEM55b/RjCuD4/3faJ8PwgE9e1gfpIMg1in/5TIkZL7H60
1t/N/N6icfoXUiAkYPacXGq6ef/2Q9T8kB342ZAM8VfUcZGrg4+4hdpAQMTb
r9SdxHzqQsSN0U8pY2ITpPRJIvk2mOA6LFWinkJLWchwi4H9GJqdNJqndPuP
M2PLEV/ZgqoHP1BovweiDtYBsCHb7Qs7FuvqThY8jiI2qQhkd02gjLOMdkYU
8lSdKIhUEYxht1KtIpl5Bw/RF6SlKMqBPqTYzY/DmAd+uWuR/QSUBzeE+/HN
wC/SyxGmHz4bVSD5IYDjobv7jHy17Mi6Yt5eU+bC0hif8bSs7C4Rr5yw+Xe0
whzFg2/FbRQfcuA7KfKqCmNl6Ueu8A7ag8txrNBn8bJ8o7Ha+4jPispPxjbS
PAtb+N54xlAf9MC8wDMJENbkUDaiD2f9KXPukwGKDThVmA0RXBJ2eitF+9oX
xyXfqcxJEGVIF3Ysa2BA8S5W0IcbuID+gWATTpp3FJBB6V3twgptkAhzd8+5
IgpYQTFecHVyMLu+QXlmMO/3neK4hh1BkM3wczSJrTGzTGVBYD3un4yMp9Q8
Otc/QAb/MmLIFjaQz80bmJErnYN5IApvPstmhd7TOlkxg8pu1uPMf8RHcMzP
caMXB+K55/qvWn1iMPQVSSXGH5o20BtHnPsp9VjgdTEe45XkoAwkJHqAbC1y
sL/1kH9+6zRZhspLkK60XnDBrBAK9j/dq/X8FT678rXRH7oY8hM87Jnb20Hv
QRNP32Ot1sFHwSwfxBLrY5qJobT7bW8bcr3B96WKYJQpVzQtyAOVFf77BX3Q
Kbb+a8fm8LZYKbnxEyzLeTjyMXo4pyOm/8+erk/+c/CBMmKOnPo4pw4pnkMh
hkjlvGMIe8/dV97b20ccqKIUeTCxoAOq95sVLuAEqfwDbtam3SOds2WPAXYD
f3u6XmDM5MytHFZ2BLWHVJe9IwfxboUt2G01bwhrqt2YtAZrmyd+S4vESsLR
JaWoho4IkbHyW8UouFSxoFzTBxsxVZWPjP73DxiwAMGmp84+8iSt+IwNqkmA
q93sPwDr8i5z1qGJGU+qpfTwfWpwdpKJ0GmcQQchhbVx3PDJ6oAq5UIrhOMc
kslJaTY6eOUVIO6hVXqZUYmLVIrF5X4Ij/xC/zWZEe9bdtAMiosPWXBeqs/+
x8z1paPVLYi1E/UcyG8DiBKkmZiBcVC6y7NClUuzYg1/J5fbLvZYiHHIImP9
EGOxqggRc2mOVqSXAJ0uSmpDgcuzGylLgkty57wWX7iUrKiaY6ZNA5xJINkq
geNIF4zPDT7rdwf0JJzRbVNLqG0kTAR9cbXYgRQdo/3ApBdXOsly4mVD3Tc7
Ok/dQO3krqKRnzJrlCtZoYI4ZS2+j+AmYwXdv18rd0y0IBpfeTJsHdS8+G3g
/ZyknUBzUvmpbf3TzSue3REqITUlGKoVEkp8sJTVGYi7ozFsh+vGqclbZXmH
mGvVOOrwdegyvte4eKqQhE3Jaz2maxdWpEbDUEoDR+55ureJxKv4Iuh1rByY
JMMj/R2wHnB6c6Dc1Rc6JEOcz528ysvooDuDpkhzb2aVm9JFAJIM4FkapVVG
NrZsUCPxbFeWwKozilskLCkhMnrh2iD2V5MvG3+xPP250mMNIlClVuuU2qJ1
qvOUBgVp0/biPKzm+htmhm+WcLPvn2zYgBIa2e/b+0KlOLrh9pyhWYh4vqig
gfep6ME8KxGQQT1tuwG6St7U1G4R7XGY60p8Weslh9XNpmW1qIbBnakV2tAe
rh/TjPHtKWzCpWHV/Aprzwnr1EQ6NkclUP35a4x1OawV1rQXfBJlNZx3m00p
tJFurOoNV8EaCOLt8sjqpIk/rnALRbxaiNF6/AUOzkylnGbW160L4I0LjgK4
znX+Ak6iTRteTXC2GvHdr4putc4E8K3Ir/e4OqO7luNlmoGz5lxzmDOXmmIM
k/fO+K/vuW6EhLYFZM5C1Oco4UqXWcy5toyGnK38qCXMM3hiDjmEHehwnp8F
424piYmtyaQqEbnoCE1nDPdxVyfv4lzdCsJnzBkuJ9gC14/vLrgyH2PB1XJU
x1PjjB1syB6Bp4gR1D8EmRvYL6RiqmGgekJ+6UclxzoIYK8aR45YOH/S6OJU
ytd2s5hbL0li3VJnimuO4/26AzatEbbTSDVP7fZl7/7I9evgUWIJJG9gaunk
S2GFH+VJRNllWwH8185qT9U/eWjS0V34TrhfpKpI5AvHtJWbRLecPumUE9lX
F8NA5CWLCXdsv8rmHl/bWuXsuDPba3uds518LR/gMei73tDJ18ftSCiPM4hb
M96R8N5qRFgRNdmh+H68kCT+25YHw1VWPE6a4taZh850tugH9Ywlq2PW4K6b
0o50/0Obj3mUMVsY/BjtJa+u4jtItLfY1SnSnMOjIVbPcTLekP3v/fu9QVmz
+gjVOkoyHfUcY16EeZPUuzKpcYb+3TkZlmpIptHm4/8EEVXF3ftuu2heu0NA
tnP6aGlbEcjfxfGCjul91I5xFDFjns3ePFQabvDOcNVLS7ZSo16oAmCBXoeq
5AP+OWppj0Yof6sM6LwKLMlddrkH7fzl4ggMIVsUrr7iCmSYa/OAXlKJy9xy
5nEEW3bse0fIu1vTY6jK8/ykG8YzNxR3Z9OMOtcdiO5cCBGQzovTq4h7wubc
/0trOhd6CSyQjG1Hh7MS4vekwq81Pdk3OPbqtxwyXRvnmdzMyyPbrG4KuKBr
1kYZtip+a7DAOBMT5MPotTPiY8o5gb6QapuRjgaXBe4FMxXEZ4k/+m5QxTz6
Iom3ZI1DWMQtu3X0reUwDrSOm1DnDMKOVrY04tarSyQohipCi1ST7c8I4fF0
L7SYUxHWhS+bQhKHbLZYQCC9d1Jt4YzvZ8dmlTz55oRzYZfQ2RdSFwQ1vpe0
z5Nuz1ljIslt/5Gmleyz1v8bJcJCC1iSx9zRVdeadrdYWIZI9Y6+5txWZ5E0
JtzE3zW68BFQIz1DLxcCtctEitOemLcKgkrTDzoVzgDFe4c0Xa4rxeKF7fjb
b7P7HgsyV5Gd2w/OpPA8oIGiVWdHLJKp5Usbr4rG5ZDu/+5j30PtH8VKY+Xd
mhwrIaSI1nCpvdLuR6oB7vCaWiu5gjwWwXMe52mwlXmSoe0glhMrNjxMo6e3
keOD0xQRJ0P3XeUx/6olma5oTlJtACBa3iHSx2o6PU3S+pGxZwKDZRATI6UJ
nlZ5+M8fIVDXMRsWMHR7QyeiguPVqPwnuXBN/CM8ZCWdtC41/M+VRyV/IPcH
4amYTHdC5m7UXywNlkrmp4LOcLDe/Svvt2eTK3g4o51DSu3p6ol225TXZUhD
2wMu3Gsk1qlaE1G9AvMDvNDhz6Ajf0st6gL7yGkv7EPSZ+NpicY9x73UBLRU
TzCVsvo3FEgA3YI0R41T4jkvSrOdHPL0pGzkOQGomaiSE9MqAMKfVMF4waDO
iyrUzdTkwSHHVvZsFP7XGKew3VfOkXtEff/w6VA0K1SZyVCpd8hBq1dZY+iH
taogSPmMeIQ/XI8PMYtEgt880r6oTspp1usx3UWdFdScJ809IciZj3wMs98I
657I+h3i105npnEztSDUk1CYBZiuuPVNDQJM1oH8k3N9U8TDyMM3BDkdhHMg
Ll5V9PzHgzB1kulK+YVlxe0N7dDtnxx3pxBLw+l1wKo7/BkvaKFQaqATB8aD
fLxS0gqurUiwK1+0AF13HI/WDMh2zKbtougTD7e/F6X3nIoZEIzD1fPT4juY
I5WJtqdjJ5t6zPmReoilDwUK9LpdQqUvw2jYqu+j1TN3OPXfRZ9jNn+DFLjQ
Tu48TucAeyDwVybvgS865bkhKyuT/kUTeCv3nFBm039ARVThoKBrzeKUsknO
8SRI5gbtp1Omt/ejoYtn+XG3hieF7GbEhqds95B6/TgkbjyPoatCk/REAceM
brElI8y6vH38Ktb8FE5AF9xRWDw08lErt/ULmCTKWB7hMYE588CX6wG4wIXT
VlLacDYEunIk7Riq9lIXsaK4pKhefPG8TeTIIDjym7K7hT/sFjodrm20RYOf
d816wXrxEXAw0j7hFRAwzghXGCvruA0NAojxIcIBrgLdfhE9+rCs6mq7y7oL
Y7LEtBRFHsoftEalNloS056g8fQu+lpTIU+oKWUcbCHuMVGtnfsWkonLf22s
ngfyJhUE3TUWD3TZCZPUIuvxqZlmAdX2bTXmN7NfC7Pc3cJbuKP/fXjOB9Lv
DGXNsSHhHWmINFI+snDBah+wtRY2buwgHwR/eZO2WviralZTE/VYHcOmQRh+
Dxsvkt2DgKFmKqsJ0cxVYU9pZj1RPC9mU1ZS/ZkuJDWhs0a9oXy59wqEkjPa
rX7MAlzAmmv5OPZU+EAKgkCZgtXKk4wLljf7/ntKJMvac19J3O8nTlkT7rRf
mrbrZoqUD4PIpqie1uWxsgiQ0pDiLmeF7qW3S98uoAWDj8kScT0hNZOzFdOh
9bnYSTIxMmuXkEmVD6PA6Inb9LkR9k0uGa+E6rcusA4Zwf4j0CTWRTOw+KQi
YjTIX4xK38pZ5hP2ZQK9yTxYCcC4VBRHvmDq7Gf7pZ8Al4ETTxJaMp4mOtoC
I428+oHZ0nCvT4GwRAM2j2DHs1XHARTJZjhn+rJy6XUzdTC6CvRruRFugKRz
71JXJSgFTxCaBVxTWoVWW7YbP58FMzB2jmCScNL5SfV6eQpcQl/r5gO7VO1n
8wkZwNzyybai9md+7nmP8gR1k96wxvDu7WlXeWUPzl0GOrPowFw1Ne2loQ9e
f3CslNf6oHTOJyFQ3e/O1pyCo8GyIewu656wKMNU1BHEDwYhvTmXnX2z5PxK
mmhpE568gyX2n4bVo5Rq14h8Lq0HaA5flwT9IeGEuInyndG3i6FpPmLj6oda
UV1g3U7kaBqz8ec9CvBBbjkMr8eRAe8p4kA13d0LPHKzeQYEXPM1lyMG4UoD
qvk5cGoffWw+GMt2KxIrIPkMaKH9OYA3CF1XKD67P66oJgx0+SHmpkBkMIlE
aIlxzRX5dVnJXylyMV4V2vttoryqK6LiX0JTkTugQSwUIkWfK6x33eKrWMQv
0s9BUFak+Dk4NEHTdgw6ZEBxQh4x2KT2G65tAQ6rR+Q8KWwWfr+WZBvY5DWN
m9e0minDQ1A2FwXE96HZu70OB3vggsCjjTiXdcvqwJ5yY3C7PdvGlJApudBR
T2R1dW9YGJsRWjtOgiZ5L5vHnV42EFKfCiZaBiTB8KuFhJE/r3i+HMxRqDZK
WdLKzZW1w1V3a08nJopb7UXgg15aPDkto5FkI/Pre8WJFGXayFpupCRgfFao
75l8WaOpKO+SMFgQZ0y1G6UivsAHSU50Wai9PNTVMn7SVdtS0nQO9pKx7DW0
84bhaCBMvIxBDZ+gKrjUAzVlmAzIbNZYJNb2EozS9G8OSD+ydKJQKlco7npn
nLkBt2vQEzPLfe1vGl/2GWmmIlSiTx6NAbyeGw7oXT0XsJfoMD8E2jwPBuf4
xLr1QvTwacI2aUUahTWsi7HZf+Jw1wyHq8kkzs+vxdkZmROAEsZCnO4ednHO
fhju4c0AMcBv6C0R6/+4J2Iczhb2B6j/UjxZCvEnFuZojRJQbX3QewauStxS
TgWpcgIXZPjNclYGbih1OocanDFSel6qc+ckDbBD/HjHuVEiALhudpeeGCZE
WOUajW41Sfj4n1D+YtannrO/Mipq401174HPRi6AfnVJWdCSih2moZ6pw/MX
06cFHJ1g1TATAA9VIwwIrGrR8aWwNeR44nJP2OWh3o3bPmsSg/T3Yr1F71Ke
1uEOGvCBnACLPWYJR0T92I0t3J4sJ6oaz2TOBSD0eOalyaAiWiKqefgY1p4H
1Moeqtnt7Kx/J4jTqFQEM8cSzP9lUNJLnfpyqSox2uYC2JMTWwvcthTp8nBh
JXjPjsVwuDInuBV6zynk2AcK0U5LJdByZU8T4D3aqeEpkiPNi+w0biw6cibW
E7PsTKanq7vBhdAGk/nKThOxnQoegr7IVbSg+CG1uTGtINMY1TEyt0KSQYK1
zClAIKrsARZ2ykt1TBQUffSSycW9d/xciQAVdJbPY+NXveE/dOHbMvSlOKWX
S07eu3EfbnqdqXIu6xZSoFbFBpxDPZ3RRE189JysMfShZPp9Za8HC0CzHXEA
0gN9GOW95Jkb3H1GtL0KeBTDlKubg0SgAmf7edpfdLiuoWYSHI0AajJvFwJP
xuCpPLOrgGU30scCgbIL+HXDlcyqz8OHrDQCkXBCJgICyyaqKr+mtXzHoJb6
Q0aMV7pqIrfHT/c1K+e3bthgyjr8eTdunKfcTaAPo7xv51iMqh4GiTI6mcW2
SOGLbyuxjaZYaiHTQRT0SgONizSGfzDk1fJJl669+zGV78/v+7hPrRdHbScH
nV4Bx09ZR7y7gxA8CIPjK1714t/GCXDc9nAlRve2VDGQUoHjV5dlEJuMIEPT
hQmP0KuzLokAlYzZVTJXcn6SqVC8mhCXvkBfhBq0/mHLtU9TGFJDl+JvowAJ
3sof3AxdePjRpF2TSloQfKKJ8JGyNAQgI3kFJIPxameDhKWl0TuEMNNwODwy
woBjG6g+NKjuPZSuOgzvzgN9UCauj+shMyWv/pJuZVSuTSusEbf9TpZHBble
GuaSic0hB99otzHxBTpRUa4OScwkQ50mszoqB3ZQTSvP9Se7YtHvzVjMOMjf
aOZoA2lbSmHY2nNX7WBcNvPO73u+ZgicYBVptjhVJjAcCVBzNy/wNEkKLwSa
HM/DqcCjT/yICi4Ff8iZHc0fau+zyZ6ANluqdikT4xnwPSahaydLKhNiBvB2
SGsbDO6fxgCsTiLmeLqqA1mLCGX0Gw2xX3I5K9mQmiekRHS8q/U9oCySotEs
bVylMgcLwgmzrtStWqDPYjMidUlA83d/g3YjbOxoFSgAeph2WKgJoDMJn6VK
vxcWy3mJ2h0BZnMxrX97Dk6efMPstomnI8CXpPAYL2dnxALR8udbMlXEg8nv
az3xAjsyf8qI+vAZnfieZbpMMbj2CnUGOpnPQ3z7Fi376BafLk7futrGgZ9l
D72GyY9wRV51NqDaS/FzpiaSKFbjdW/CjlfGuhkW3DVV4IEnHkaffNaDjpcW
yioKNhP4GHXHcmzOhp2J4TYk7TAHmZYvv9PJZUeDNQkdtLsAvMFK11BHtCFG
RBlbk8/FpGsmwouyb+ilIYj2SoW1BDek+YRXA/z+/aWPZzlT6zgaYcc1XcZw
r/IpjEmpUv4DOJa9Ad5drWu8ixmjIjgF0FBhsIDW27S7nxmfIrwws0fFkgft
eDFYDt3d/x1ly+ZWHdtrXZ93NrTcXCgddj5aIfT+FHZSC8lycjzOdTwh+m2Q
MzlhCjCod/qQ8JNQfkXKSAson7JftrYn3u76k4TzdZW4i2UOgi5aL6LFv5vf
YlHK86ztuRxQcG0XLEFZgX34+mS1eY04dSr+MJNffKmDuMSGTXoVW7MjSwjX
T3Ckc9RJ9PoYZywZcsOXBg8k6p+mYJ/fcz3KRJPfkjVWsVZroDRJx0HkTVKx
bUdAPPtAIMieIn4aQysp6PIS893QFTOHS+pJPg1VB8kUlEsCFGSG9KzB91Ij
FzQrdCx9x9WrBYMzR+trzojqT1oJHHNQkwCzWXq4GsDc2dcd2+3obmINTkbL
q7ijiigl10OkhxdrlEy6gsh/eZwAUCOyOxfhPT50VVmi/yPF2ipxhEnFL1rI
7dDT2iQaCps56YYtWe4coil0GxiSV5neE97TcPlqtrRAIvCOpXW8rrRHgxMy
QB2dsqPuA/Jxcz94nffxRSHgpQo7nngznvkJaQmnwX74KhR2PmlVP5fls2Ba
WbQuYlBPyPJ45zuYk8XRGPIfpmjTxigAqL0TExOIEKCNoUefseQycEtvuk7+
iOcEjPqQZedlcrJ4cKPQCAwYu4OR2Z2/lrqgCZa+PNhG7ir9uokVC0BOv2Jz
w35qrHc3Iah+87AAhzm1CrN/KSHvsOtPKMlXbW+m8V+zGMBBh4d1EEIPIr1n
zrgpNFAQak+k7OCryhXVCeE1dDZN1cWHC24Gld0WnS4mMSW4tEZv077q+YjW
B/lCL30VOZjH73TOj0IGCHH4qg89M3MNhtR/0tL7g0wbmfxoLl2FgtR/HnU8
dGrJ3F6gJmdSyue05BDxYz3dmDxmxTfx/hr05IiMSw5LRbRfeYVud35tj3RW
/BdBlRZE4dzAA/cowYgkKFNrKcUi+Y41gl3NZtQlBj0ettHSPdaNKjKOm2tl
J1a8DX1LPvxFUuUmLzbhbKPhRtgFw7RNe9NyuUvzUEvDbGs9c9RVPzr/8jS1
Du80nb5JDr8Ix0E33KG+NzYpaFRTBsCwaoyUp7BjtRfO8YPXCOhle+oXS551
jAAud92kgMs2E5PWwGPjc1Rs+KDH/oXV/28Ga1TPH7nyVAjyDt7FQ7Wod9MC
F6nHdXEAitLMyphKK5EF0xBFQNEDIQUucZ48ktiLH+iBqZt6//r3Mvgn4UvO
yWGzt4Ef7X3VcqHu/1gRb7A3iCLvg10C4+7aX0pDJ5WVDv87Z7kHmoB8XSkm
CDJnnoEG7Gw3wWqBqr4Odffk4Akgq2T3mRrUJ9i4tYluqlbBlX83fPtptAJE
rquWj+ZWk3hF8KeVW2KxWd8cj4TbNYZ39WjUs28Ce3Fvco2LgfGwJaYFX+Mn
EmfsCoisbuVS38hcgRjbMEDnWvLzDnde2aNSVUgjYCYXqjoP9q9vMEFxnQLZ
0RilgsIWt2kadWBUoq4KF3ByBlQGmD/YtkTmfXZGqDeolh2/MSa7ghVTtX08
TPKhMm2nvCqood4tx02JfHaeqnLz3EwbJp/1rBkAwM97GqYNjgkqHiqlvRFe
U4E3eB9Hz5+Yg6PplJdkn8dvG7Z07A0YT8EUy0s/JNhAaX+leCzfSP416+j3
z9ZVxkCoARu7NtGKU9pQcrJDe9bk4X0QIoUykwTTpZoEWXC+8Jt6ZGXz9dSl
waRPVItU8s3yzEQo4hZjwYsVJWErmGUj2ozGPM5YGmC23VaPb1Fyvz2qFGVY
MVFe3C9s1PpsqhdOzVO2rbRBxPRbXlf4RwVWPIQ/ERgta6rtSAko9Vkakbrf
ZS57xvljqSNk0FAU+Wb35m3aNHzWhDKE5ssaRCkbrVEnFukx6l9GiuhT7CUD
rksu3AC/2I23sQn8I5PGsfxksbqcj/GcAI+m1fOKMTM2nHbnXBrtgJhWMIqG
+bAU3teUvlQn9C28T10saJTWzEW9dO7D/OPi9hXwZQRTYikuc0TM3t8SqbDU
nkI9yzCfD2kT4UU15eQYM0BzfgxvuyAFKvLsF200Vf1dda5j7BbGwyzZ3+kH
4NiDtxv7KyJlMoZ18hNiQI+rLipKL/82dvU1pS7YvabEvtfHdhpDSPO5ONb/
cfJZX1dfza62xd+9VAPGFoRG59AzsJWGhaVTRjXzjcD+Ey4cvrm70el/M+U5
SttcqrO/sr270rF4/fX7UflhzjOPi/4WGDWSrcZ7O/j/QRmI/zsFdcp6QOh8
ewyMi9ObW51LaEBxsLsXAyMwqGxpperHHCnGFn70+udOA4OqjEWwom2ACUCs
Dv/355WtKJ0fF+BszHdsO3VUvImwWAiEayTP6982hJdDOMMIhFAO8wYURHTU
h9oFEHfABYmfCbS7XrcxOgXNsAUY/o/0wExjGQ57R73PnWIq3SBCjinmxMsz
a8e/KSkr58eqjqmRXen73K5cCbAz0oxlxlqN5YnGU9IaJ/W703ozYZJd0h8u
g9i5Kra280k4+xnbXMWYZCDLhEsFGaMX5YZtnl+wBSacbRcyCGZ/tOn4QdGc
84j2J8J5rXEGNgVdEHikTr0qbtiQPpjASA9Y85R5PRs799T9EXNDxCaUqmRf
j/WPGRys4Nr8LGySlNVRFoc2ydoXBjeet2Cy4GueyWGnDEwzKuOCDQJ6HEii
ZuqNduaJGz19vBc3SLMVeMp4iDdUb69MpKGqZsRCdTb8SxGHTfIzmL7pH1YC
vrQt7yQRse2+jKnvvZtLqf+woa2pN7OXCWItaBkB5ZMCaXUSfDElY6NximxH
YLxuTJHex5cVUmvUs86+P2Invc6Mh8Xn8WGdJzaTrZhFpnF3+NArAge0DAlM
NaisLHPrFIKMlRgJ39+mEme7x6QkIhQHhMNxd2PjHppKHJfECBjgpDCEuhvd
+RzCbOcq8610otRySfO5OX8XNXcuFKOBwl26P3cbf5pEGTW8OPkqe4yPTHtb
4+0SPFgb3h0rKqbnKQjhsGzCbLiAevTTtRsvAt1IknN2ikS7XBW1iDEa35+v
NnjZi7gFXhAE2SL8XUimOX+hqx8AeNMX1wnrvUBMFvMs93lBbqpW8JIrJ/7h
8OM+CGAUQeNug57F0CMZBx3XGlDoM7kTRTIPxUDEhm0lq/kuYIOdTezfB91R
bO0hn2Eg8KIdJ1xxJ3ukt2Oq6vYumfPAhAVjR3ZTs2dHY2FSEythz1rYu7TJ
wVNoC859uuzHG5xRokc2/0mp+Sblvu0/QhEgLmHsKMAQOt1z0KHJMi6DGElU
EjZOqkMUk7JQnAMyRnTfQGERqYth1K/t03zLgnVgPi0ZIkGUmot8b8MSYV5B
zfeWPl5i+TG7bS/Xa0Q90uyodM8/LJLpr6abO+raNJXSIDhWmLpEUk2zJ7EJ
nPxw/JXf1TcodrS3UCMpkSQK16quwUvdAaUSwZmdkR0cr3PwF6eyVDamJge9
zDy/X2IQwi2brfy0TMCaMLMl7z/HpWNnfDFuj6PBXcaAt2Lx8QuxsxVNucL9
VAvHnD7kd7cUEn8OBCC32v+hI6zyaiBVNXzi9UPonTVZB7HdUxAQ0c6UJUuK
uO+Z2FRoyTe+5tHNQ+UyeVDbt4/gyDhL+0688udyOeStq1JF3PVSzf5Y0B03
RgIxqWK+2heyUHTzSgO0R/we+8OjUodLF/G0su+ykTNEXP2yC+i0eds3LTEx
Np5drAOMUW1K1CcntONfki17AUvMck6C2QpugC+umZUdCYfYgzHjYugaX27k
e6HzBNe3Mq9M+xTpsIb3TsuVKquXDIUix7AQR/dHv5yerWgTWWrFiKHCZE1L
0V5uMILBn8pk5Pvdfec55R99m1vXwRb5lIwmyNnsdILJBYRdb5fv3Cmer1zI
0ziJunpunilKtQD9gBHARgFOmgPd8k9m4sNeATHXELHQdF7KLgYlIVjnLtCa
sxyjsM26doVIbNmW2d0PqGmVFlq7hD9Gsf3315i8dXNdrixzkriSYbMeyvX1
If2LmVQmvpT4/5Q3vmcJPYkb4Q4E7d57BL6+vpbsqT0NY+Lw0tdc/gytdZyT
f8o16nbZbVhk/9VHno/DD0fvJwKAADgY85ZTL5AAX9Cra93qFRMiviJ8kbzP
Fe8jUGQx12U1VaVHIkmZiufFdUjg5GaqSJkviykm5w94+daE7mGF8ieCDSRg
OMotDalio15QLDNfOPh3tn92hfQAAM47hsLManEQ8CTMJa+UEF8Bl9/ZOHHH
7tEgyxh0+HVDkatappyDOO4AKYPW1vSpc2HieVOjhwdLQD2acsvdcLXrw51B
KP2FIYq1xTyoEpjHgv4UqWxlmGBy/W50dgwMsYAHrODSxCeegbTyr419+Iiu
GIuz5aGfEPwIV3VeY9/VyconGAurnJwn85EgnPjXWDex7QCRalTVT2JOzOOw
/OyabCgf3iV6ZPGUZAEdnlXUPW9EA5aZeEtM2SzuI2vi3WyX+gZRtMU6vHdS
SYoGujWlBnwA

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1LJkMh5kz/fkanidglmNkoUZUotKtYsVloV06zUezDA2rqFfUWIsY/ZOVF9SMAIIVdQ5Vtydrqhv3vuOM76gYPT0jWDTnt8j2lymuBtQnpBnHTJ6bFi81k0GpUgzL32O4HkL7U4aZ32hmSRD7XqeRSelou76CXLAZ2HOzSi36Ga0SmXXHt/QefRTHKsLvD7AMnNx+PD1NP00RGWJXzQrGKRSs05AUhsIE0vW/cNRAjmJgh8jfGYbdoun0mh468wL3BP7Q16Qj+hpF3dx5UKw4Mh5HSZ8B/ywFNU+zKkRbaaoMn0elnWNbvjA7IprNRP2VSZ35hI2nNTqGV97gA2WcWPucZsaAKZt8KzHxy1QciReG3hmZ65ZCBA1scBOoFeRJTQ1fC0F1mSO+VlgO0Moe1imzVfV6FVQuuXQfWTVMAes+2C7gJEzZCw6nWa28qBzIJWzWUe4ibIXq6p9DYBzqdDIXGulBh/RXT+u5qunqjq29lYh3XKvGRz8lrDlawlLlgCMvFoG2GmGC120w+s+FHAD8AtWo/K0J/h3FjJyRan6HYduI7Z8P6scTTVPBWpEqXoLm5AOo5M8aSbuJwEafF3sZ6OyRZ6MjDU0KZKCNCknwsN051UMKv1jyNwT+bLhtcEf4Gv8u/NJh5V6wluBvmgXivE2Y//timt+HZ66hlqrW5AObMW8RgoIkcVxaI0SyNXLnoF2lIlBTHg23RawXUKkQnSPwRhujCxbe3CWcAYtOwgQUTWOUjKZwQs+J5BPZPIrow54H3EV55lvJavHRVL"
`endif