module emif_cal_two_ch_altera_emif_cal_iossm_274_psjm22a #(
   parameter NUM_CALBUS_USED                                    = 0,
   parameter IOSSM_USE_MODEL                                    = 0,
   parameter USE_SYNTH_FOR_SIM                                  = 0,
   parameter USE_SOFT_NIOS                                      = 0,
   parameter IOSSM_SIM_NIOS_PERIOD_PS                           = 0,
   parameter SEQ_GPT_GLOBAL_PAR_VER                             = 0,
   parameter SEQ_GPT_NIOS_C_VER                                 = 0,
   parameter SEQ_GPT_COLUMN_ID                                  = 0,
   parameter SEQ_GPT_NUM_IOPACKS                                = 0,
   parameter SEQ_GPT_NIOS_CLK_FREQ_KHZ                          = 0,
   parameter SIM_SEQ_GPT_NIOS_CLK_FREQ_KHZ                      = 0,
   parameter SEQ_GPT_PARAM_TABLE_SIZE                           = 0,
   parameter SEQ_GPT_GLOBAL_SKIP_STEPS                          = 0,
   parameter SIM_SEQ_GPT_GLOBAL_SKIP_STEPS                      = 0,
   parameter SEQ_GPT_GLOBAL_CAL_CONFIG                          = 0,
   parameter SEQ_GPT_SLAVE_CLK_DIVIDER                          = 0,
   parameter PORT_CAL_DEBUG_ADDRESS_WIDTH                       = 0,
   parameter PORT_CAL_DEBUG_RDATA_WIDTH                         = 0,
   parameter PORT_CAL_DEBUG_WDATA_WIDTH                         = 0,
   parameter PORT_CAL_DEBUG_BYTEEN_WIDTH                        = 0,
   parameter PORT_CALBUS_ADDRESS_WIDTH                          = 0,
   parameter PORT_CALBUS_WDATA_WIDTH                            = 0,
   parameter PORT_CALBUS_RDATA_WIDTH                            = 0,
   parameter PORT_CALBUS_SEQ_PARAM_TBL_WIDTH                    = 0,
   parameter PORT_VJI_IR_IN_WIDTH                               = 0,
   parameter PORT_VJI_IR_OUT_WIDTH                              = 0
) (
   output logic            cal_debug_waitrequest,
   input  logic            cal_debug_read,
   input  logic            cal_debug_write,
   input  logic [26:0]     cal_debug_addr,
   output logic [31:0]     cal_debug_read_data,
   input  logic [31:0]     cal_debug_write_data,
   input  logic [3:0]      cal_debug_byteenable,
   output logic            cal_debug_read_data_valid,
   input  logic            cal_debug_clk,
   input  logic            cal_debug_reset_n,
   output logic            calbus_read_0,
   output logic            calbus_write_0,
   output logic [19:0]     calbus_address_0,
   output logic [31:0]     calbus_wdata_0,
   input  logic [31:0]     calbus_rdata_0,
   input  logic [4095:0]   calbus_seq_param_tbl_0,
   output logic            calbus_read_1,
   output logic            calbus_write_1,
   output logic [19:0]     calbus_address_1,
   output logic [31:0]     calbus_wdata_1,
   input  logic [31:0]     calbus_rdata_1,
   input  logic [4095:0]   calbus_seq_param_tbl_1,
   output logic            calbus_read_2,
   output logic            calbus_write_2,
   output logic [19:0]     calbus_address_2,
   output logic [31:0]     calbus_wdata_2,
   input  logic [31:0]     calbus_rdata_2,
   input  logic [4095:0]   calbus_seq_param_tbl_2,
   output logic            calbus_read_3,
   output logic            calbus_write_3,
   output logic [19:0]     calbus_address_3,
   output logic [31:0]     calbus_wdata_3,
   input  logic [31:0]     calbus_rdata_3,
   input  logic [4095:0]   calbus_seq_param_tbl_3,
   output logic            calbus_read_4,
   output logic            calbus_write_4,
   output logic [19:0]     calbus_address_4,
   output logic [31:0]     calbus_wdata_4,
   input  logic [31:0]     calbus_rdata_4,
   input  logic [4095:0]   calbus_seq_param_tbl_4,
   output logic            calbus_read_5,
   output logic            calbus_write_5,
   output logic [19:0]     calbus_address_5,
   output logic [31:0]     calbus_wdata_5,
   input  logic [31:0]     calbus_rdata_5,
   input  logic [4095:0]   calbus_seq_param_tbl_5,
   output logic            calbus_read_6,
   output logic            calbus_write_6,
   output logic [19:0]     calbus_address_6,
   output logic [31:0]     calbus_wdata_6,
   input  logic [31:0]     calbus_rdata_6,
   input  logic [4095:0]   calbus_seq_param_tbl_6,
   output logic            calbus_read_7,
   output logic            calbus_write_7,
   output logic [19:0]     calbus_address_7,
   output logic [31:0]     calbus_wdata_7,
   input  logic [31:0]     calbus_rdata_7,
   input  logic [4095:0]   calbus_seq_param_tbl_7,
   output logic            calbus_read_8,
   output logic            calbus_write_8,
   output logic [19:0]     calbus_address_8,
   output logic [31:0]     calbus_wdata_8,
   input  logic [31:0]     calbus_rdata_8,
   input  logic [4095:0]   calbus_seq_param_tbl_8,
   output logic            calbus_read_9,
   output logic            calbus_write_9,
   output logic [19:0]     calbus_address_9,
   output logic [31:0]     calbus_wdata_9,
   input  logic [31:0]     calbus_rdata_9,
   input  logic [4095:0]   calbus_seq_param_tbl_9,
   output logic            calbus_read_10,
   output logic            calbus_write_10,
   output logic [19:0]     calbus_address_10,
   output logic [31:0]     calbus_wdata_10,
   input  logic [31:0]     calbus_rdata_10,
   input  logic [4095:0]   calbus_seq_param_tbl_10,
   output logic            calbus_read_11,
   output logic            calbus_write_11,
   output logic [19:0]     calbus_address_11,
   output logic [31:0]     calbus_wdata_11,
   input  logic [31:0]     calbus_rdata_11,
   input  logic [4095:0]   calbus_seq_param_tbl_11,
   output logic            calbus_read_12,
   output logic            calbus_write_12,
   output logic [19:0]     calbus_address_12,
   output logic [31:0]     calbus_wdata_12,
   input  logic [31:0]     calbus_rdata_12,
   input  logic [4095:0]   calbus_seq_param_tbl_12,
   output logic            calbus_read_13,
   output logic            calbus_write_13,
   output logic [19:0]     calbus_address_13,
   output logic [31:0]     calbus_wdata_13,
   input  logic [31:0]     calbus_rdata_13,
   input  logic [4095:0]   calbus_seq_param_tbl_13,
   output logic            calbus_read_14,
   output logic            calbus_write_14,
   output logic [19:0]     calbus_address_14,
   output logic [31:0]     calbus_wdata_14,
   input  logic [31:0]     calbus_rdata_14,
   input  logic [4095:0]   calbus_seq_param_tbl_14,
   output logic            calbus_read_15,
   output logic            calbus_write_15,
   output logic [19:0]     calbus_address_15,
   output logic [31:0]     calbus_wdata_15,
   input  logic [31:0]     calbus_rdata_15,
   input  logic [4095:0]   calbus_seq_param_tbl_15,
   output logic            calbus_clk,
   input  logic [1:0]      vji_ir_in,
   output logic [1:0]      vji_ir_out,
   input  logic            vji_jtag_state_rti,
   input  logic            vji_tck,
   input  logic            vji_tdi,
   output logic            vji_tdo,
   input  logic            vji_virtual_state_cdr,
   input  logic            vji_virtual_state_sdr,
   input  logic            vji_virtual_state_udr,
   input  logic            vji_virtual_state_uir
);
   timeunit 1ns;
   timeprecision 1ps;

   emif_cal_two_ch_altera_emif_cal_iossm_274_psjm22a_arch # (
      .NUM_CALBUS_USED (NUM_CALBUS_USED),
      .IOSSM_USE_MODEL (IOSSM_USE_MODEL),
      .USE_SYNTH_FOR_SIM (USE_SYNTH_FOR_SIM),
      .USE_SOFT_NIOS (USE_SOFT_NIOS),
      .IOSSM_SIM_NIOS_PERIOD_PS (IOSSM_SIM_NIOS_PERIOD_PS),
      .SEQ_GPT_GLOBAL_PAR_VER (SEQ_GPT_GLOBAL_PAR_VER),
      .SEQ_GPT_NIOS_C_VER (SEQ_GPT_NIOS_C_VER),
      .SEQ_GPT_COLUMN_ID (SEQ_GPT_COLUMN_ID),
      .SEQ_GPT_NUM_IOPACKS (SEQ_GPT_NUM_IOPACKS),
      .SEQ_GPT_NIOS_CLK_FREQ_KHZ (SEQ_GPT_NIOS_CLK_FREQ_KHZ),
      .SIM_SEQ_GPT_NIOS_CLK_FREQ_KHZ (SIM_SEQ_GPT_NIOS_CLK_FREQ_KHZ),
      .SEQ_GPT_PARAM_TABLE_SIZE (SEQ_GPT_PARAM_TABLE_SIZE),
      .SEQ_GPT_GLOBAL_SKIP_STEPS (SEQ_GPT_GLOBAL_SKIP_STEPS),
      .SIM_SEQ_GPT_GLOBAL_SKIP_STEPS (SIM_SEQ_GPT_GLOBAL_SKIP_STEPS),
      .SEQ_GPT_GLOBAL_CAL_CONFIG (SEQ_GPT_GLOBAL_CAL_CONFIG),
      .SEQ_GPT_SLAVE_CLK_DIVIDER (SEQ_GPT_SLAVE_CLK_DIVIDER),
      .PORT_CAL_DEBUG_ADDRESS_WIDTH (PORT_CAL_DEBUG_ADDRESS_WIDTH),
      .PORT_CAL_DEBUG_RDATA_WIDTH (PORT_CAL_DEBUG_RDATA_WIDTH),
      .PORT_CAL_DEBUG_WDATA_WIDTH (PORT_CAL_DEBUG_WDATA_WIDTH),
      .PORT_CAL_DEBUG_BYTEEN_WIDTH (PORT_CAL_DEBUG_BYTEEN_WIDTH),
      .PORT_CALBUS_ADDRESS_WIDTH (PORT_CALBUS_ADDRESS_WIDTH),
      .PORT_CALBUS_WDATA_WIDTH (PORT_CALBUS_WDATA_WIDTH),
      .PORT_CALBUS_RDATA_WIDTH (PORT_CALBUS_RDATA_WIDTH),
      .PORT_CALBUS_SEQ_PARAM_TBL_WIDTH (PORT_CALBUS_SEQ_PARAM_TBL_WIDTH),
      .PORT_VJI_IR_IN_WIDTH (PORT_VJI_IR_IN_WIDTH),
      .PORT_VJI_IR_OUT_WIDTH (PORT_VJI_IR_OUT_WIDTH),
      .SEQ_USE_SIM_PARAMS ("on"),
      .IOSSM_CODE_HEX_FILENAME ("emif_cal_two_ch_altera_emif_cal_iossm_274_psjm22a_code.hex"),
      .IOSSM_SIM_GPT_HEX_FILENAME ("emif_cal_two_ch_altera_emif_cal_iossm_274_psjm22a_sim_global_param_tbl.hex"),
      .IOSSM_SYNTH_GPT_HEX_FILENAME ("emif_cal_two_ch_altera_emif_cal_iossm_274_psjm22a_synth_global_param_tbl.hex")
   ) arch_inst (
      .cal_debug_waitrequest (cal_debug_waitrequest),
      .cal_debug_read (cal_debug_read),
      .cal_debug_write (cal_debug_write),
      .cal_debug_addr (cal_debug_addr),
      .cal_debug_read_data (cal_debug_read_data),
      .cal_debug_write_data (cal_debug_write_data),
      .cal_debug_byteenable (cal_debug_byteenable),
      .cal_debug_read_data_valid (cal_debug_read_data_valid),
      .cal_debug_clk (cal_debug_clk),
      .cal_debug_reset_n (cal_debug_reset_n),
      .calbus_read_0 (calbus_read_0),
      .calbus_write_0 (calbus_write_0),
      .calbus_address_0 (calbus_address_0),
      .calbus_wdata_0 (calbus_wdata_0),
      .calbus_rdata_0 (calbus_rdata_0),
      .calbus_seq_param_tbl_0 (calbus_seq_param_tbl_0),
      .calbus_read_1 (calbus_read_1),
      .calbus_write_1 (calbus_write_1),
      .calbus_address_1 (calbus_address_1),
      .calbus_wdata_1 (calbus_wdata_1),
      .calbus_rdata_1 (calbus_rdata_1),
      .calbus_seq_param_tbl_1 (calbus_seq_param_tbl_1),
      .calbus_read_2 (calbus_read_2),
      .calbus_write_2 (calbus_write_2),
      .calbus_address_2 (calbus_address_2),
      .calbus_wdata_2 (calbus_wdata_2),
      .calbus_rdata_2 (calbus_rdata_2),
      .calbus_seq_param_tbl_2 (calbus_seq_param_tbl_2),
      .calbus_read_3 (calbus_read_3),
      .calbus_write_3 (calbus_write_3),
      .calbus_address_3 (calbus_address_3),
      .calbus_wdata_3 (calbus_wdata_3),
      .calbus_rdata_3 (calbus_rdata_3),
      .calbus_seq_param_tbl_3 (calbus_seq_param_tbl_3),
      .calbus_read_4 (calbus_read_4),
      .calbus_write_4 (calbus_write_4),
      .calbus_address_4 (calbus_address_4),
      .calbus_wdata_4 (calbus_wdata_4),
      .calbus_rdata_4 (calbus_rdata_4),
      .calbus_seq_param_tbl_4 (calbus_seq_param_tbl_4),
      .calbus_read_5 (calbus_read_5),
      .calbus_write_5 (calbus_write_5),
      .calbus_address_5 (calbus_address_5),
      .calbus_wdata_5 (calbus_wdata_5),
      .calbus_rdata_5 (calbus_rdata_5),
      .calbus_seq_param_tbl_5 (calbus_seq_param_tbl_5),
      .calbus_read_6 (calbus_read_6),
      .calbus_write_6 (calbus_write_6),
      .calbus_address_6 (calbus_address_6),
      .calbus_wdata_6 (calbus_wdata_6),
      .calbus_rdata_6 (calbus_rdata_6),
      .calbus_seq_param_tbl_6 (calbus_seq_param_tbl_6),
      .calbus_read_7 (calbus_read_7),
      .calbus_write_7 (calbus_write_7),
      .calbus_address_7 (calbus_address_7),
      .calbus_wdata_7 (calbus_wdata_7),
      .calbus_rdata_7 (calbus_rdata_7),
      .calbus_seq_param_tbl_7 (calbus_seq_param_tbl_7),
      .calbus_read_8 (calbus_read_8),
      .calbus_write_8 (calbus_write_8),
      .calbus_address_8 (calbus_address_8),
      .calbus_wdata_8 (calbus_wdata_8),
      .calbus_rdata_8 (calbus_rdata_8),
      .calbus_seq_param_tbl_8 (calbus_seq_param_tbl_8),
      .calbus_read_9 (calbus_read_9),
      .calbus_write_9 (calbus_write_9),
      .calbus_address_9 (calbus_address_9),
      .calbus_wdata_9 (calbus_wdata_9),
      .calbus_rdata_9 (calbus_rdata_9),
      .calbus_seq_param_tbl_9 (calbus_seq_param_tbl_9),
      .calbus_read_10 (calbus_read_10),
      .calbus_write_10 (calbus_write_10),
      .calbus_address_10 (calbus_address_10),
      .calbus_wdata_10 (calbus_wdata_10),
      .calbus_rdata_10 (calbus_rdata_10),
      .calbus_seq_param_tbl_10 (calbus_seq_param_tbl_10),
      .calbus_read_11 (calbus_read_11),
      .calbus_write_11 (calbus_write_11),
      .calbus_address_11 (calbus_address_11),
      .calbus_wdata_11 (calbus_wdata_11),
      .calbus_rdata_11 (calbus_rdata_11),
      .calbus_seq_param_tbl_11 (calbus_seq_param_tbl_11),
      .calbus_read_12 (calbus_read_12),
      .calbus_write_12 (calbus_write_12),
      .calbus_address_12 (calbus_address_12),
      .calbus_wdata_12 (calbus_wdata_12),
      .calbus_rdata_12 (calbus_rdata_12),
      .calbus_seq_param_tbl_12 (calbus_seq_param_tbl_12),
      .calbus_read_13 (calbus_read_13),
      .calbus_write_13 (calbus_write_13),
      .calbus_address_13 (calbus_address_13),
      .calbus_wdata_13 (calbus_wdata_13),
      .calbus_rdata_13 (calbus_rdata_13),
      .calbus_seq_param_tbl_13 (calbus_seq_param_tbl_13),
      .calbus_read_14 (calbus_read_14),
      .calbus_write_14 (calbus_write_14),
      .calbus_address_14 (calbus_address_14),
      .calbus_wdata_14 (calbus_wdata_14),
      .calbus_rdata_14 (calbus_rdata_14),
      .calbus_seq_param_tbl_14 (calbus_seq_param_tbl_14),
      .calbus_read_15 (calbus_read_15),
      .calbus_write_15 (calbus_write_15),
      .calbus_address_15 (calbus_address_15),
      .calbus_wdata_15 (calbus_wdata_15),
      .calbus_rdata_15 (calbus_rdata_15),
      .calbus_seq_param_tbl_15 (calbus_seq_param_tbl_15),
      .calbus_clk (calbus_clk),
      .vji_ir_in (vji_ir_in),
      .vji_ir_out (vji_ir_out),
      .vji_jtag_state_rti (vji_jtag_state_rti),
      .vji_tck (vji_tck),
      .vji_tdi (vji_tdi),
      .vji_tdo (vji_tdo),
      .vji_virtual_state_cdr (vji_virtual_state_cdr),
      .vji_virtual_state_sdr (vji_virtual_state_sdr),
      .vji_virtual_state_udr (vji_virtual_state_udr),
      .vji_virtual_state_uir (vji_virtual_state_uir)
   );
endmodule
