// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vzM01p2cUtEOQV+gqxx4132HACxLrmF72mZwSfGDM8B369gTzl4isy2Q/o8H
3isy9MUyG89DlJ+agKuDKESdzBVU0T+VWt0J2inmhknfnDffQrrZi8stcwcr
Otg8giJELAIpUTou80SwHiHBbsNgoKC7sQizNQ9ajVvJNASYjmAHNlmU/B51
L7mK4LlcD1rlgLfFtNfTDijCOsDdd//6TkVcf3K95i1AELInzjUgSBfldCg0
JD1nxCA0c3dwjZ77nxfrGbU0rKokkybDxm0B5R4WGAjL63bOomqrqpzp/AZA
0s4I6SaihsCflCYCFTYt12kZQ3KSpAORebpwkWC6Bg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e32qGR5w7jEN50FTi8LdWc5xRH1QAcp7d9HoKMjD9VJZqj6AeelRLejRLmM2
qxuo4r3hvolHXuIDnx/gB2KRX/2zpmK7RcQjbLnWajUnry0/7hLCy1cjIg8/
c2vxj9ouGYa6AmW5yW4PQgutu1dfIVtiIgRLz0KoV4dCryhj7DviUJbaa2rT
KoipprvaZvzSR8KMrwFJMbyE8Wly2jQxRgFpnYBH86tQRPe9JKWR1YL0VHqV
ZHQALrQKDM2TgcPqSvHBBIQGvgelFTi62w+GA8ubpvVm4PiuciPK1eeftNjk
3fmyP/et34rVVtgJ/VIN0V/peTcx7Ccp+vbwIAiWeQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ga7sE4W4FrWFOxHw2+6pCQepGNeGpuS6odT8aXpib/lKWDXQrGuWenD47PFM
Nqhk1bNYFKq6QbOUjYlNWa7IdPOoZIxj9OZkgYzdgxOV55ScNyIaSiMRNXVH
pM0sinAf701Xo+aYqAaTgT4+upji85OIyK1K2QyUt8d6MsRnux0WbZ4PhWol
pQJLE3VzStMEgC55nUlNFxpv1MQQCeY18vaaum4fQu0/gsalQxf/WU/A3v9o
HKi65qAIqYGReE0ctTgGNGczidF1ym10ITDn16e157Yl6lcbeFrOcMpJ6bKp
PyVcEHCNI2bwH2pag/dBXdtP3qQn3lPiKLnYjBafPg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HJhl6/YRoinRTvR92RBC9i6jlzud3QLMrumlNZ5Tct2OnhPp9SZlenO2YYJs
VmLzOGZIALypNlBzpAwKg57uFGio3QFwH8/Q02IdBztailW84X7vibWZ8d9P
jNVa9lRI3v4CiQvLLuYraxU5tz+wfLtCvrS5nwuXB8iAycksp//3x1jmjl8x
rZIkdj237f7F59xneWAMtDDqtEzfAkWV/XICIl9rm574nqkds5pdSg/v/1Hh
GK+XpCr9pJPw96tOzv5hj3arPlVc666cQX6JvOQ3C1mVhW2gE4aSkbXoukB3
4au4BlQ7jLHNXdpC976JLuk9mx+tCgpAQ62OGA7pgA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tSsKaIV7dpyJGwiE8oDXV7qy5QLMQPjkib2kVTZM3/oVuJVCiVo19feRjeqV
/6r81L70F+Pg2jM1I0KvHco2KHkybLV2mEtf96Kl/IvdPSG8YfkSZOkappIX
xhHsZq2LHvVHYA4Bhwy56kd3wjvdNAln+uk2D29U8b/Y1sYS6dA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
otuTcIFV+ggrClJ8hyOhUOk98GJ/nC6H/taGqhntI6LOPFcFwUudm1oxAogL
JfYlUSi0oFamRo32X34H1yvgCZVn4zzDWCCvGdwTyTLM8LrtkNwwOhGRZlRc
5ltr0EoVnZRVPgoPnmCQFUkCW6pP3J0ZMGRYv/1b9dvfzNFpkVjVdYhOYkwy
NUPq2ujkgnQcK+j0lwMLKa5QnxHP9Cfvo3lqfpskpCwzWoguKWx3+WeSqDBm
qmEttuJoyEPKmoYRbI3dI1zf8hsnJX8RjLwupVWQpCMjbV6tD/RJywhXgtY9
VaoE3/6hPH/FOUGpUcwD5GIXyHjXlxi0g0G1LbUeT/N96ulrjTO25t9xuXdK
wZnlTVTYopH7QIahiaC4dcOiDoTynqBKtiSacNOdT9jv2QpcrHtWZteEAGJ8
uUOWCzaHhZJz8qlAo+F4iAPXDhigsbpkeAdy2H0J4VcaBE9iaolUVXhFNysC
x3QxxwT39cEMuuUefVUcU5ssQV1T1lcH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JUMfchm9b+7Vkg9gx4kCGBndSsV9vO0Upl8NmnhVMmS3dFHy/SgrYLjeA5sA
I+fAkN1oEvcGQZnODYJ4w6k+PlEgtornMgQc29dNoeMsH2v3vCUsOiWY2+Wj
IBeqFSwVzEDpJjWT+CNlUZefjC55I0nY9YWdH3Ip+on9KHUwd04=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e3O1larhrpOgl0F9WmsfmtjSJKO5bKWlOFz2HOkstdNZSxYBd2/16bpTeuym
0PJoPH0pBgabVXw2w1KFebte/sbHNTmzCdrVf9/+r1g5UKqZhUoVh/tzrrgh
rkOLghEUa6C56d+blOGXoN1+z2Of080out098CsqsLtvuAiJzvQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
rxqgdAwe8xq2d0I85vaq3VxqmgArVKLNo2sXWLKAxFHLeFOI8INJIgbkAb84
on2jAJ4iK7wtBtVn+7W54fZGU/D2Jo31w+LqaGLgf6DrjE0g/80bsQPJs0Mz
3BK+stZPb2wbSdSIZkuxZiOlUZFgQidmES8+B4/xbIBnK0WHBGGVD4GGbhxe
Po936o87b12iNyA98ghbywQMpvheoaFCNdM69/UORSPYyxY7QdXgt8n29Se0
2Zmc78ksYQXY8IXFi5Yu/EGaXHWmpFojnWByeUp1CrVNcSIG+gnGbUYumQTF
93TKgmCDqjX4LAl64oNhAHRi0RfSKWApdsOCTy4+6oE0z39JFNnGWW1rpzY0
LpN3RFvDlF2ytfUhTT0Ky2ExPI2HEDHwwk/YSFp9LS81fHOoinmbv3ofRu0k
KoVztxCY+/YAxumUe08DQMr5b8usJKb+bVSJfbNXaeZNvxGm7EaCj08BNFe0
ME8cYh3stg8Vki+a56U/nF/yPQQhR9MPha/dUysSUaFs8+XxMktwkzqpxI/J
z3ld0KppaYU9Kt5LXZilg7gmmu6TxZgKc3sjZuWC5KmsMpOBeGH9JtOeBvQi
m0s2XFMWzvSUbQHtIDp4XM4MeXZb5KHDPo8zBTtgQxmLAxl2L0LLrit0aFOh
RfcJyhi2oVNwNKrzB1CsEfRywai+uCReOwbw+l1uBFG8JAv0DmYtHBVXuHoE
EA33ysq5L4QbYLw6YS0ue8B/ozKLwn8s9R/UD1zUR3meu1qkxYDS7d2kaLRx
mjONALVGWjBUYpc+eGwPpswtlD55FI/ruDXiy/vUDbHjzl+pTbZoPbrbiJ/d
TuPfYFsU8COazbcvgLKnc7Rq+fUVtbyrp1EHdUg2jn9XzppkXPDhWcPYECrc
ZnQegq8kwVOg6sX5YPCPufTWXfzVgWW3Uu2jbHF8IkbueQlzxU9S3N+Sa/sV
PNkUXVnSFtdLzAKJbAcSvxGSoCKbOMhfj9sZRujNIxfYlOdK5vTgqflYSEPn
aAv9IuBXz+J0DBHhrNLj9rIvNcLy3IJnIaA5SbF+PJkDHoyID+WT4b1TNFU5
PWi3psuAMnjxpqN2iZF6vsTFc9U5jWdgp1CHDmxhJOExRKDeWWsHIt/04JTS
0MwTevduejgT44nmndIGLPOQVtgpzAr55gQlS74ApAaIxi0iIJdKTRwpgsie
ZtE9XmCarZf8dzJNYzOJ/K/2HxlG1Knk/bxww7plGdPUqsL8KV/ql9UZCjYC
P641duhq8QzE4u8rUlepcPRiVviWxz9Q7jJ1XO7VpNJZk6L3Uy4mYOGWik3h
mquBQZh89QDNdP2eY8ikAoxE36OSDTni4T/HYFmpUEMqQQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqd8J5hY2UZWznk42gZn/LWeSpQ4xRBgssnYqpz/rw8PnoKyGzAdUrv6MpRosQ+hmHtzHz201M3Cc0FUosn5bYICKYPtUwPgon8YUXlY1QHrJ8PFE/rWa2uttJ/G2traGnlTGvHT1cKK4ubC3R65E+oux+GjVb/btE8U0D8FGCuT8Y5nt3Gb0+j7KJWw4AGcVCXf2PhreJUXnPi4YAxo715aq21g2tHjLjYCRW0vDpYh9hf3JrZJ+VL5c6eLfviDGtvi9c675NOTIKpuR1d1hI+32YIbZiZrtJB38hkNLq3gP9WN1v/pDDVbqPIth6uf2Aj5CPDE1ZYJw25s/Y7q8W4jx6FYPAI5rdxnIdfhKtRzjlFkBeer7lXNgyoLh0hS1M455ckZM7Z/ROhjmh2YCQgAUGvooV09jpXV45h1lSGtmIin6Xhwcj+8ewFH3bCsTwxBpz1St9HNseuRc6WsSmD/yhgM++K1rOGxyUOY699s1jwhK7hFySy4dwzrZTVests1404R7YISZ//HJln6tPMe0KVNDAE1aHN2tLNqXtsgx5Idyou+/vmi5thb80EFLXPkPCmI1aFmwLUFYmT9Hl+NWdVKh5n3VOWjCozu1VUE82gtAFLaJYUNT8Ke7+HjdX3sQDeDdjKEOVXK48wlG7zT6Q8K2Gt4qjZxT2AL23t+VpqAw4+uu0NUPE4BvLCTPmyEPWp7GjYK13VyjtSuk3K9+XsQqQmaQkken1HSs2NvKd4LuqC0pqlwx9sW+qUk/pZD9U/EL28fyKfIk1pHMYRs"
`endif