// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UmivB+FFteGWvenNwwd94hvsm2OOZixnd3je0VJY9gy4pBan9TuKUtGIf65H
kMiT7SYuEdtgwoXQzihWEiWK6jyY+DNi4C1Tl20kaDTMRDiXYuESwiba/8JC
w13gdqI+2cyD4FRYv6t+os+tsNSNH6Oe6b8jLXk6Vg+9rWUN+sBoftDryXc2
v1MA1fnD7RpUdQje+aDIc0wPGszfssXMNl44KU5o/DBghu3GnGES0EwVaN35
ZYwRLyRrpXta3KtPxSjNEIEtVEihV4x7Z+Zqw3/OcvpKcCscxO9zvDnyuP6F
ngDebU2JI2BeCIBu2Nx/aV1J+5vBvcqHNsOim43ySg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UQk9JUsAF0dhyIo4emXYbtjFah07p3ohWC7jxk77ViQqLElrtgiaYOZGFdGK
+/9cGPBbIXJlr+qaxBMbPTsy7n/w7Lo7yJKr8ynHiHWXu1MfvPop0UEKBiol
zDaqwgU+hvpzTrjNNnkWmcH9tdXaSvImwCJdWHplWr0uzQEhJLWXbJ799k0w
4BqULD/UdlW0Bc+I1IjeJkg4eBWw9nKFmjcIWTjzwHw5rFIknHDC5s+7iq1/
2Fr2YcCRnvB7X5FecJOU3YFIMJxK/EOIfTRY/drTrP4Kc0vZ4rdjwbtOOjxN
OA9D/E6P+qtebkPK56KzdYbtEK3ZTutG+aybDqX47g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mmA5s7bUDWGDdSd1aIXh2C0x3jhPFZVs94/loU020rNlWebhG1kZz3ByKbnf
yuBYPIxE5iqaXFYAooc2OjbI2viKtNZCnhPFhAaV9Deyx8hvK3MVBcqrVRlC
sekS4+d2jYGynQmod2irY1Mlp42aBRsoULWZ4qAkAU23HZMKLjgsREYl+5D0
A+Fc0t0d9ySnLkV53xSsLczXlYi1OtHHeePwAfh3mDM3Ab7S5rp6/q0XTT9U
2KDaK4x7L2OrdDiDDs74Y5jz3fz0lLArq2v3WlVZMUaCNXX7Ek4f7YLed64Q
0pEu2668u8fCLCNj7S823+gPFd5ILOzK0csFAtWVpw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bSoSYbnFLqGxuVWZnTRLqWN1hkR5c4ZgfA0vIIC545a29r1GH85lBe0agl2j
jVp5Emj1KtRbASrOtX3BNN07K3CjMQ5B/3dpeYu5yzNrj8ao2mX6A82ya+PV
+rOjwpNokd4F9CEs2qrS3BhPI94AZmMVI4ekHLR6RROgOE0gAq8xE59zJIK/
Uu+uQ4wsqSIPRsdHuw3quGY3g9d/ZQ68oDRuZ6mZB7H21as/qoG5iqIhZHjJ
wRHcyhn6nJk8we8Pvwa6e0S8JJ6CvGw3Cn8E5k+urxn6fAGrjrkyk3BYeecB
Yly+YEhc+eqhLQyGtq2LkQIjzav31BNebNxHfxSYSw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CzU89tHHc+16Me8SYDKbmSc7HqFKpKbhUjQTRndr3RZRbfFN/zzjkbJZcV6z
Zm6wXky45Cnn2uulNnw5/ttUpnESLIUbWXqtKDO/9taPfAiD5dY+KEC3uGAG
hXBXQVLKHN49qZnmi2QI1kY3xSHuOViyyQd34PIhSjVdTz5g55o=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xn+LB+y0D5nY35WE0GxHXBmg2Ysp894XtaAKfLk+/8EqWzwCzeXxKX/V5GQH
2t8vqg+X37nZySfDQeOQnuAfL3rUqmqIRY+smyWyNgSO8cAmOMoSeHECLSCv
nzQf/KNb0ftg/ECw371y130jXgaUbLbBs1DLgECpQhyv/u7tf52c/59+Pfve
1vzeJWFXXAWUa9iXshnun0lQB+XTcRAilWqEAA2g2ItgPd78AcTvnfBwB3+o
tEqh/UuXN0/um/GMECAdF/11ednYGq6TQoPTAnnBhZVT7ftv8xQEel4L0YQX
elbLoIX47bfTcAOeXVjwlVl7PS/LFBKFFrhZDHDca/FaBnLiU8ax8Q/IgeFp
j2cjl0k6W7XcnqCbwCMSBfhrD+qXp67rtKCjK81Y3nfnmFsB7KrXTZxtn4p/
4IUWE4U1W5h/nKTHzaFLu1QaKHsbtFWR9i849GaE1viOyBA3k7NahqFQm53Q
BV3BkUkfRxKXu29saXk6MTnDPokKQnzW


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kHFVZafU/3FWbYg+PMImgpEFvv+E9Rn8BQHV8sk4sSL4I7frH958NxW5YuT9
gei/M+P7eZPl/E1Bks7TT6gVIL8G1Ue/nlzqWlwWV7dbgtIOMvztLik7Vcaa
qJneEQQerOcnRLsRbqrKVUOMEOLe3zajMCZ7nmiM+U07P28izV4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R7VcGJNBVl5cdUuDEzUsNmoUMFrZs6kDp5hXA1whHafyFGwjjFyuC0qqVAMR
+u5nhjpJmf0zz1XVf5xnKiZOm5brEEY2TKlNlhphuqRn/fqBrdvtawZGmH5Q
1slQ6aWMAMmboPTJ5+RyydJlsAxt+XF/bx7U8+l62ZjISZcZ32E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 20016)
`pragma protect data_block
gKmHV/2A/Wstb4kuISLNC26CVaYeyrl6QSu5SFZvPYhaAGGgX4fPXRGyYZWP
0ca4cGLOh0kLP2Cuzvc3GCQcg8h08eQ5PrK2obqRb92vN5sBbS/6AbTNgZW3
d42/fsynQyoGBGDF8wVyTnRIgQmVJea+aWWDvgN/gqPvgeaLFtMYShuu+cjS
IfC22wIgkyCxYnKWCOIylrmjhCmoDFJo7BFH0ECnK3EzsfCbOTLG8LOvM+Y2
0hfDBZPEW5Q/xJ+uC3yshVpST4dLMSV5bjPZDXVkNFVnek7lliFLhD6U6sTc
sPvMKeK3R+URdxh2HYTQd96VlF1pEDY+xnndjstkTjMwdkgl2ch9rEYgd47G
Z0OpxWflYJ2EMtVn5idbp9SU0+GntTtVB6E9qRN1PQKI//4YDksHZf9Z4FT+
p+h4I/skBJzWLs16Q8KIuKJkbizw7NXrzOq6tILUUKcBUujWDD5EwN4JGlDG
rBcFIg0nkJOhCiK8Me/4C6x/1CprGpc9qh47BfrDjxkX9EiTC/6y85al2NwG
yRHdWD7aS+uBWlpRVMJPe7XzmXzzyqa1l25OsJp9Rxrgl3p9jLOsbr2m2v0d
h+YjbzanvCRmX3OhucWynthBDYj4WejEkloIBQllS9UWxIiEtThSBlt9n3wQ
U0sUwA4xZdo2iZ1wNWkd26fHQ09QxPvVkjuY+ZS+rQESU1HT1CKGlIEYP1ys
G4LTXCUzxatpxBUcx6HChQgC7JIG6G6Jl9n3i+BVItE6OjbV2gOgr82JVmfh
E+YxibVmlTI/BHNllKRQdxXzOCZoktUGE+BNlcnL2ZS5rsaXyOjd7ShcRbBd
LnmrQAS1SB8vra9oh49hFOos9YPxXIfBfpedKiHEJKpHl+jhlH8hJa4x7Wa6
DaWJXBT9dQ4iHjxyP29Ud7WOoLevbGoBeF2332M7doYwCX9yDllqPfK3KAGK
m1uOmi0XoN4jNgOpkn8ASvwHIFFX7qIhXWF12goNh8X4c7pS5WrKvg7HF6YO
OrfTtFhZQc7iO446kMpbEzcMInZbDjqNIhUFpjhtGiY/nud0UXf//1oXrLJZ
qTKhrV0RKjv1WVkyRyYRM5dzILqvHhlft4iDmmI/AF6xC3XMDDBZc1oPAL7J
epNCgJt9rO1j4nYsqTNm4Xx1t9ORwsLgIb757IBqBCTQ04AAg6ETjbqWPngf
8+Le37NpiXUrukglpdVMNeb3Ak203Cwad4GEqdRAGOqUYpZh1eKzkEcTO80X
4Rarg9F4spbHgtL5X7RdfcfUiTXtMY/l3hPkVMcShzJxGwxbkW45sJOIGqqB
mEYwlnIJNmNFh/+yVJBK/k+uxbH4Jm+EeDJF/yf548+ekLOzDIF4FSuyMaS8
cznDTWwSbNaxcEB028tVt2ysWvG5i2/t0R+b02jgPaEhkt3k/EYRDP5JqmdR
tjdGyVxPVUePWoutaRNSWG3oVQ2qNlBvls4xOgR9gaoyx7Nns0xptxxpdWiT
rN7jSfeWHZRAE1wKkWv0Dgo0obCvvHVX60tu8c8PnhWtglgdZsoXkhyw7U2u
bLNHjTJenwnDfhyqEGG55/Enk0e1ulrKqMt5FtgERYVRBp6zO8J0c2WFrdEM
4k1MAE4vNsTttAbvQLBwtvnipmfPIuy9ZXHYUMG5LMfswrSiT6snt+OigQT+
60TLQ+EH6HmVxghp2DSjFGtXx7O7b5UsrOurenuDMhHbDVZuUcp9slVWSsy7
tMl0VMUJe0Omi3r7prrUfs4pTaOG4EgCyi9g9W3zOKMuce9htzDZgPONAXOs
yzJwLHyQ4L5JqFHXGMaTXO92pM6E9o+jkk2QNo1qtiHnnUIHzJlMGSpX3sDi
W8BFOaX/8VEp4i904+D1mw0WFhnFeLeYm0p9uPI6RJ0oJ5oxf4BJoFI+CLhr
6hkmBjXLbR+4HNqluex1vAx4Ofxc5QhsCFX5QAPJ0I7SJ4Rn0K+KRd6Dqr+8
3NTOSDNRMi5pWBSi91G1ppaIbvk03gs8C55MXvYJ7yz1bsKEKbR6+iJfQ8fU
zKAzc/D0fGwZ+nCjfV9yFBiQWzcLMgOcHwSYf6Q54yNRxkW+yYU8NOWE33Lw
Yfo04qDBNuAmiqO06fZVo1G9L2aW8zSiNghNINz/uMQx4uD764Xyx6v4+5XL
nT+o5Sy5J8ti4SmRzQDbA4cd9XkzhqJCrR0IJBzXPwxn9omi449Il2rEmybA
RsVrCQgoNXO83YTUv3+C19nVndUDGYjclCvx6XNip9+gfc5NDHxpafza0ZBN
urhEN2kY82yzUgJxwR3xVXjxUAGEzVZh243U8TqVsR25waFu4M1VtOru9hgd
JE9sH1zJFQCuxAIcWT/a83VimkEOBkxo4C0ZthzstWasUjHrpVUc3MMAVF79
sj1EmvoSknMvkNEqq+sUiqa+QUf7e+GWgktYexaK8ivYtWjyVAsklwwn3L67
S117M+8BEbc7D3CD9/WpcXqaZv2GUxTjRNTf9EAh6HJk43YaMDIp7Y7WJpAP
3/Q0z9QVT7AUQZWiQ4XUcufLf8zbbE2B6hU93WarV0IJA5Y+dBnb2rkN6Hax
vGadMEYKpvT3AObmR8v2A2ilP/yjZFda6cfOuNMWRzlBB8LLL3C5dJYORBsH
E5J39QU8SzQsK6nwPJBRZ5is47LbgsREFZSdZqyesNjlYMfSoyTB6oItqtLb
okWVgTAxWgReWqLTCgs8Zx242heqNfyMzbab8QWXw8wTXLL+HppYnRUZsOM+
MQNDR/W6epG6VdSAlfHeb6J++3q0QG/7JCkxhzGT/AEdaBoTB26r6KkpZCVt
rxui7sVYH5rK4a/wwHpO6en2Kh0JnW0+GkUL3cSA/VRE2jtv3VloJViynxfL
cKzkO00R91vXw9oUoyjYLH08OGCBdaex6lQadSQwEUKKB7EtmXBlPBRw0VI1
cXg8wZPlLs/8Dx1KHuj8MgS7w9hDwdbxSXHtgiuZPZsgvYvr6/m3PpmrfP4s
d10myJDrHAAwumDmw+od70GboWolKXpnaRJBeNNOHWua1tJUqXD1RKOOUiGf
k8Nz3b7h2Tu3qwys7Lvmwk1X2m8zzqifd+1Kq9UubblH8h3tIPLAqay9Nr6s
9R9xQ/SxbYJLcNMYl7fGGGV+yxFnkrqVNrFn24J7wBC2JdDEM5/L4m8Ucsnn
aISkWym7JTfcmLip7hF2I3nyViUT3UPUxWv3TT5om8PSrW9lQM2FZdhMqfHQ
5ql/4LejPa9jLMvc1A+lua/VwqFJvUg4x4PjVJQjrzhajygXj/mQx3T5OWW0
SovHSfK89lS61Jm5IK6N65AZhKXd8RlEEIm5Blg7Y9NtAt5D3wHt6HiW4RKj
Dq7uS09gxAqrnzbCDhWBND9gAmCqeCoGIrASGJZcFe3i+FAftOLyUNDYU2P5
GVi1pEL0m0xUpvSOa9KHDb1P6YB0ntOSLW2lCJY8qHtmLNxtxWUAPL1ohDlz
0kPFWCeBJ3M0I0nelVz62W1S+GGXTWJzJezRvyD8fwqQf+51S74MZJlYleKp
M5U26EG+8ji+lZwRU6w4LcugXGKoyMATNJGv4ag676glC5R3C1bAvs+snlfG
OrITbsDlQZfF2Z0lnYJqrsob8IZ2+O1vrxW2L/lLbMtkqaVN8gzSELsc8iju
47/50bk4FUbvu/4K6NfGDQC0IbyeC28rXh4M34Iy52qPkXiZQadrTjsQfxTY
a8PcdV9rMWWfFSz09dBrJpMC+Phjjyu7r/Lp6K7yFDiR9MZu6RQ3F1BwPI/z
k56Qd2HHrc0EKjrlT6P1vYl/Ea/dMfBrHWXFMCEV+yZRu+8hhhSm6C7lGMO1
NUPm6jD8FehsNtSFUfCsBPvWxgo6Ph5d4vK/CxP+Zg3HiHbOSlnkXezZArw4
wjM2CAV2ksGoAHWschk16FfhMwc3WOLxzc2lPXcbVtSZUTFgEKe+OYjtE8Q5
oqIiWl+25Gb48ZQx6CkBZG4AYQzjeWRwmWYv/bR8TCNWDi6Tl7lVh2kr8wOB
5kzadu5iEjKDGBw10GMYbgzDNdfmQF9EjI+HPSjcH9ndDVPvrpJzBCXlpqPS
/05g3fk9z6k98AZ8yk1fGFdopQExyU6FF86F0RsUDaVxyExs7EIELHhQDoLJ
WvxwG3hP8b58D+8BT43DxYSYu/2aXHJ0H40qhh2m3j9dnPY4uA3h+9mpONBd
ApUOkvrnXqhBnlA2r0/HKy1sb5FR2qbaVgSpZfp3xaPxEkwlxbueR9GRdH8b
ez9kft6CTCVUjXwNr0eSewZeO4hPPj28Vfkua6AAP/0pJZjNI1j0zEWTzL0G
G1x1ZGS0nibzaA9vf378QkJupRHR6xiREJ2xv1NxVFZQsZIQ2CBmkKLTfP1X
lE15uH3iMU7dhl5nrM4l9Z/QyY61fOburashsvCn+oAO/JTT0Us8WfU2ww/x
Q9S43jlC592Pz6d3iDZjEs3qvbflC2FkH2y0pnYHm1zGj+fjmMJWN20Dilwi
zQl66Gq9BHIybUFzMp640nd437nrWorFQUsTcsdLblCEVrSdwuzRdI2oY1Wq
9mGYMY1UC/n3AAPAK6yUoRsqHLodNwHmfS8D/ZN798xJ9tsvWa2aRFnEx8xl
alEnlONZSXw/b6GuNdHaPq5IlxCWd2gs9nJZv4ygFZ+GVMT75TGDWH8VjTF8
hCUr7IsoTWMVrtnWxSKQReMCqPIz5fNyQaeu+ehO4GUOxrMXD60qXdOMGnGA
jkWGH38QV6z+f27cGTjX3nDjlxXFqrGt1ZyXA3lnldBW+N/QOcVtBpOSbMKe
TYsOBQNSRIcwdraXaEtyPyQwqr4YPkk+l/LQ+7370OwyrA6PCq86pns44Vs3
tOpPGR3DgfHv7ClPgoFFvqe/wCuGoWQFtSuiUypHUj6+6oQC1GMqSk6ah13B
KnY7yK8Np/7XXj+wdxpa461TfvP0Ap1Gb6axnjEV4lKJTpBrt2gjIqx327ga
7J1dLQhdgktc3/qu9qC+RQahP98JiUeFK+/Gh8cUlUaAV4j4PUFdHiSVgRPd
1UepQBFdFUlyBBWPhrj2cV8z6K9JcPCDgYIj+ulLW/rZduyhK+x05u6nox4F
wIIJLCTu8nQ02Fo7YvDlCO10Vqj1jMx+1zddt7GaRZB0uEBwtV7Za4r4rgEK
Q5g4jn0io9A9DTR/ot5R+oRMjsk2oMHUiNfctuugYpJ6PBHbMhRy3dHT/OhO
K07XFFUjQOz2nEXjdW79M5zt1kFAZAPCRSL49UZhEdR8R1duiMJBC9OiUpCX
OJAYYRCg/egXRp969Bn4cEuVjzI+JOKh25Nsp4DR9i0BgJ96fUgoXpCsoRqH
0CJPoQdUaLhPpKkb+dq1tUwOBq8wALT6d9FJ920TTXpNz0/hUoY7x2MuUwq5
8syT1dZKp3aqLSgPxq7bUIdCuoQFn+9VYgdyzt4BYcITGEwFkBsFwYPHm8D5
RoUuy0oLirJBMOoQFtKgrJHzuSm+zgNUwekWsiltynRsZpEDeqFZ/xiJnVFA
6lNttig/SlxsLTYboBJzJIiZNsrMB2gj04rgCMh6WkKOqYMaieCUu/e1cwOs
x15bbfPbEk7YuQ+mbOTiQLjFkn6IUnswiKZGOsU/GeVvJje/fi3mNPi8nsKc
NHHRCE9wb6WH8fqsYVM3ZU5bh6hGYxIIVaZ+mqjp8zvepabRMCgoQnpo6SCO
+umzxn+/4jbXJw3rQpVb0qrNju6eu1BQu760EHdvlOMZZBRIM3+tHDVRvGuV
tUYAMCS7WvnMHZpUw4NcW5RBvwK6790qplC2LI4O24+3iBnCtj/PBPcP9Fi3
m1Tw8sd44HxJyOM8QDd6kk9TCwJtgHxfYR5ew0c3xmoTxsRX781vEPiGsMQe
neGTwS06Gg1vld1qVjCfvT2rWwpM2431BHOFpQoPxmn+WY35ZMSGydOeKCRv
YgOhJP4J0W0W97RQOqtTMiawnIC7/UQ3a0jSyO/ZNl8UEqF7tu8CKrLwr2Ur
2aUBuNtjz9XgANcESuPF8FZBUhdssujK/1mqufUWAglPhWM825gSSmSzzXJs
/uxdPkjVOB2zyaJOmTQRb4tfhpBt4r4FtLKP7w9VspwxDRwerGMomxySRBe5
W1FZ9WwJER3lk+hyjZEe7QGAqdYsbq27h2CLTHWDHdlyrwxdKUPlRifCNDT3
OT2rnV+uksD01xusXMGngMFWUBrH35AG7qQ/4nVbezZvB2XDDYWvIxYnSKYZ
IFjO7T3VJDRekd0ZfcBWXgAaUdhb4F4ENxlREiY+bS2hgXzeUpQVGrrlf4UF
n7qIQLI/8ryyiRzpFT7tVVzglawLM1ZBv4zVvi8iWL2NUKAQRYXxKzRYvEZi
MV9J5jPme2+IBw12kFaGVpzp7HMojhQsXTCpHEgGJ3XcilC/Phie+ZyghvuU
6nxVWJUu2PQfDC62vG+EOBWEWSwtDtwoGXzPQGGpJaqiGe18gzcnCchUXO46
blZlXEV/XVxokVv6uW3h7twwpFiX8IwOi15i2qQ5r+xDMAu2aX7eV6Z5oV/i
dyx0OnD896pccHaUK/ZWXB3mQSUQlRQRAaECTXjieglvxVS+nBYa99as9oZw
8EWTb9tVa8BfAhtA0i5u76eY1dxQrX1lBmx87w8dmgdx561j6mH4Td3XqRj6
DnZJbVmqcmy6BSyNyFjMbJMgn9YNakm52ogT/0l705WpjVtek6ZK/vuAUgkY
GzwOYiZeyyuLF1BKdLCkMGqaxiNOMdFnBHJEFnoeWGw1KKNAm0Zoo1a8GRU4
CTDMqJvbMEWxDasknOPCLoGkNDPwkgtiaWk7l3YWTfSTj1KLNdeTKuUCFGVf
ai4pBkwTwEkRhLdV0cmKN/CCkX7hQGjhaLdNjkYdUvGrX4B2N3NSzTLxJ2qq
uHZebKj5o47UW1RKpJF2LDCszK4+B9Z8GvAKuBA+9vW2cUHXqvSjgqUD3NMN
EWhWeXja309OESXaC0yki4eIMDMCUxsSBQFpBhDnK2KsVlJAB03TrGbwhCzt
pDUhx075+b5zQrxqSUk9MoheJM9fHzXYPciIpt1qIcmIcMU8hQ2jdZLjrhRW
c3oAMOb0WPTdGTzf3AB+PKerqBj6gVRU9WHX0DC2rJ+If+BZBoU3X7o8bzb9
AdBhLaUsh1FHjrxTbh1d+ETcLkrtNUROdltuTfmGV/U5aGQZto5KcZMV93RO
EkgaUF3Zlyr98jQc+kYzQELtH//OX7/X/B4lRGB+hk+d6Znurkj/Yd1qw9e1
RXnkGn2yfRfOsERkXT/l6teSDMMdkvP18+7s9Q9Cty6pr6QnZ8Xg7KAaMhjP
XtoDaAOfSTI1+Y+Rp77sa00GSSfh8ZV1HWJ2o0FT7GrEPNdSLJFaAJ9Rv1j8
O7uCYlYnB+nY2QZmqz9se6CkL8h6h8a0wwjl04y6HuqrDYcRRz/wxp1dignK
qfNG8iwk0Be1PMw/v3OoD5PJx5ePTAeDCATL/fCrQWkNFbDs+gsPPQjIJZ9S
UYfkn/87bRxr3S7pwBc9St2XDfU7jmsKzAccv6SEUF3aECb9vlf9mioKGa3G
ypLCA3niS8wieRSlzJHbwTFEfF6X4RNg2YpKNcDMDMPZ2AQUgKfUvtmK7Dm0
o2TW/NNnB6hw8vRvHz7Atr7xNYZfc7Iq4KOLuC4zEiEU4eTwDg7Phc7l5jgi
mqC8CX0hA4ujbV2SVtoAu9se15JRL5DKCR05L6N4NWwsPWo0LfGcYIdfN4bE
1/gT65/gJVS7JkbD2cvgmHcl+1vszldN3f3HCBgoVpt5fI25iFZzG7TDzPH7
RdVvQDfRylRahdlfZdg01ULozpWauioFQ7vRojsQODB1inlopPFIEaj4KY7S
Iu8BQFbiLG3qshu2j4IRJMSkRUTW2EA9tRSC8drtXsgNFLHDkNtb7WeJY2ht
NXfcufiQ4arpT6EFAe/Efc5oKha5IRyK3nJ4ImMT38R5WOdX8Ar21aotamuO
Dr6y9GfZmjVLE5NeabQYjMFqVgPYLXTQKx1pBt7VTqVIrQF6zk6qeICb5SaC
b9BcBH8EmWEyRu7dBRehycYvyvSudS6glulAwEOg7pyco9QcpHKRB0q+Y/Wy
aLWFGktr3HK8LF1fC0smjvfQ9IaSR7pJyslUCjzSoXBVumVV2hhjENpf5UtR
V2ZXTCzbjAgRdAzOHmGt6KvyJB3Yzr7adDxjsJG6wN1xg5RsLLyPv2YUdRl1
bEu7eoqIALzEtV92EOSx1WhBU495hUjeAtt+bUPcZHHzvF7/eluHsWsiplbZ
nlG6Z13LvjrU+bBZvjGk3Q0W30LDZwarfPANU195D/2Jc13El+sRbUAbLjVO
+MRGyOFJTXpOHXh9rktFJLT/xNY/bWGrmukGT+ZtWFCJt8tVhCbpzmKtYXah
R3cqqKWywCb8oOq1JQdguDPoZysp6Jq2BfsVkJjcCRxKnvGckJ5nLG6vqx54
X4eXDzX/GWTdG44stpx43pjXq7JX1SND/dpq7GbUqNd4CRYXyQnRoIKdbz4D
Rx0C/XVmAN0vD7KK6DutEyBbbcX3RH2I17ONT5zwvPjsd3ZFrufKOq1wFIIH
katTOmhp4vJ2YjRqK2gJ6cxHsyp5n+LBSDLyIIQq/HNU6cZ6JF96Xayr1Kmm
wQzGBfQTfy7/abLNpru3XuYfOHKy0IP7E1Dnl8fiSkQkuOMhHnHMqCWyqE2d
vXJF0fdXsuiBvsw3YlAaPki4IbUzM4aaxgbSZmHN6UGYmuvkGDvm1XrXVaLf
Cr/57c1M3uzYwv6PCjomBD11SuD/qtEGYPWpHmMfuGQFgDoBJaO/xjUE57tX
s5nNGhlG6ln7D6bWShXsYDMJbhjC4iyfswUkU4aOUJAItrXLq4GQbK/RG9wQ
bdpxomizzs+ho3o6cJYKqcE9v4ODX1WB6eLrpdDdRtIqyhcXJd0X/+CUBZoI
Aq8PRWCvLAn2cNKeQAr2sH6U0OCk3CuWcDSh/6zY6BtH7W4XHNUpgso+mGNd
iotGPZIyaWRCZoRxQlKzIMRmcu3lWP3kN7o4Ot8F+G125HqvChhU9LZRD5/S
QpEr2FySnPN3uOQ3UlYygzh8u9tZ09ddz9RRgqoLEGJGVDzbsfqGVei8pK54
4B/GGED6+gawo6oIP1zjkv+mOCmvN3ZS32J6WAurLOYi9xATRV5kj3b4oGN8
GMVnzZqp5G877uPZBZ44t4hTXKyS8XmE/+UI3cOXkVLEAeu37P3n+/LA5sJ+
hmVBUFM6tQyblTq2Y8/+e9Y+RWS/bwtV0mbaODNHpoNv9TTgAkdwLLnYjiRr
LLA6DligGkC6g9U+CRMarboe56H2pc1varrEpTg/xRN7Mrpht/NkZ8MqWtTb
/qkubGJCDmIbpycd0yqTup4rSb+hCXPB8Ckw9k9vG191528Oq2voXsag6U4T
oScYzw2x0UnRcW0AJ9hN+hjfn0CDR1DRBf3zr7l4QPbdJZsm82c4UOX83QCr
ogIqmvf+pMg7i8Q4TP90MJjtZZqzSZPZBSnO1swjjEdiN4z4mA922agZQUgY
1HtVsahII1XhK972AfkEIra/g91ien1IEzKrhfvVaGUDd3tZqIgo9QArBpFx
d710b8Na/QbtiD0ByyFDqu/aMUa1v7d7dsd1plnxSkmHRu32GVCdNu0GzsvP
cJeEuWZ88jnQbOj1/jZ7cxUWpU1qzdDF3W7HscfKoF09AY2RLBJQFhBHzJo9
FqdBVVnTNnAWIE52mvPnMwC2QKfa8DDHE46wL+vxC4Td6ntjyyBxZICRNBga
w8Vzjp1WjeZ/Eh4dhr7d71BaFnaojausgxtyism2iwlKvGnRahEQIIhulSwr
JXzZSHGNR5M0aobRjoqO83fiaTsiRRyKD8M1Osy6MDz1zqgCMQA2biH9+VBA
2fPT0+DN90LdEBROwGjwzHgiu6CPuw5ZxPq/EU+RIgBGQL7L6oxzRX1PVJdz
ib6HJc7gRGPB44s0g4JFs5qc4JUsamiXQlw9ugFbnUEZj0QR4i4rGzLlAxa1
KeXHUIi+YCX8ooOFvDJosEjoV6ymwk/6tMQCGLBZActpjD8lk+iwls+/8sSI
vpi8lldgLbTDQ5vvkU8WWQSQsC8DJQn0b81vZdIwS9AX40UZcp5yyDbPMZE0
04PxjWyxJbiaKdY1KFXitWvL2uLd7leb/l9kL8Be8L9uZI3NTD9/x5FcZrVk
0ZN0zenucN/tcldsq2pBlKr92Rme5J4NUG9dps++yprWzzTp+QGoRoSnUOUV
oAQeH/C8As+T4XZkdjLjZx6c/DJow5wD/RlHWoks00CXf49kydnMUWhMv2jx
uSALkdgdiAvqZ4tJ2LqyvgQ+14Zu7t/CUbHSYUOLZXOfq0yC5gLc1okZyV6v
b6Ua0+LawGFrcpA2vnxyhwmiwMROJYUW8UqW60bw5cPda+j5+XyklarfUliK
zbrxXf425uTG9TKtT7Jzd71ePprj4xnYnTB1X3ukm7XrgrEHjhboeAmrkckk
6RkEyPtKRzkCLvxZ73+37825oJAfJ4dVOzLHkEeHzkk2DgWwONLNJ8mzwLLM
s9c+h68L4OWro7mJbNflD5h72xXUb01ZqxvabueM+4N3GEqj6NEpBlQng9PH
aG1tl8QSrvQ8Fm0Qs95yDvvyyehmR7ICK4S/HjfcjaEt8vUXjgdM45CM1kH6
MiTSGNAcEcbCZXkcw9TXwOa2spHEg76OxAYIWiU0IgGL1Bvj0kkrh4/wVKqh
OGePZBOKkuMuI5vcp7rU19K9gifbnJ3nP3wY9c+7ISsubIdrJhvDMTo/fpKX
eduKY8HBAnsUeQBbFkFnD9P24JgTW58chT0A4IzE/bdbAi2HCGiNZyEDCBy0
lm0rTA1CSflMoNy8aWCLn0XfwpdQSF7vCofQQFYB53/s899URWXSYbDH434e
xZRXMJlkUjLXVeEhqw8rwc0zQB+byj5obAikZs3Co/EhQ9NwFcPiy9m98Jco
03/KbSqUFVdGecHCub1dLp4yQDncp0gfCpevHi2f8JXsjq6DJ7f2Y+5jT99M
ljDob3LhcnA18xNiULjfUqV7tPre6TkaWTjC9NuTXaRZXLtjoCTND/alpyQQ
vXjHP7yCMQlqOYl8EcRG0u/GMqQWkRl2OJjDQNkydYB7/HIYXjJ8Et1XNoF5
zEl99gsAVE87xkt5AMuwdjPFjrPXuFG1KU4fBn61ghmq7iHBOO/fEnWYBgX3
rfT+MShDELVlDM8JGwWs/bYj4XY7tTuKxYnreLWkXFYZ5X8Eiappr58lG7rd
2h1bHJHwvoqT4ZQBs3HPy2SJSSXwAKgjWs3lK540/hlPcVhnxqCExrDGWCce
ixElyOZ3WgBHRitQMbmtPwNvQhla+sipvsshlpv0K+a6zOXufmdEESQnbR/8
5G5y8HSitbAWf8jvXvG6HlCGgqFdlLf1z/u2sE40Evz4sBkWFM64ps0aZTeo
ain1nXlkYOla4pLmiGeoIqdHd2UOmBLmqcQCwbvRWnuA9B6/iNpphlh1+U+W
CifVJ5wLaWafNYn1Dp4iUTomwTHcIEervecA+9IBfCOS362dw+yPyLNuwHJZ
PuAZ22N4xrFnXTXkIU0sGKOGJRWbjECRfBdZ5vpo9xEpgtNhbPKpTerykpwJ
N+CXSfmWf6Cq+Iuw+VNdUjFx2sQd5Dy9gGCt5jHF6T7PXKPQAhdKqVBO27vG
eCMb0liyEFrKTCY5uWVAlLqVL+gidnzgb8zFubsC27y/Ouoxyw1Xl5SZaezz
Ngyh3F5ZJkHyCwq0f8FVispSh3w2u603Y4CTmdw1KnEF7sbG778zrHyX/Ctr
uLV/NXwxA0oLrRVUZ91L7fWOQAS019uua8aFlCggjz4g2MgzLBMif+HFL5Tg
LxpjGXaIQDV+GeQW1n/51OScUJmBpnJCnl9SHxEzcQWuI2HXnG5Rk8KUvzKq
oaNDsS8zq2Uif8m5OHpY7zpgQzh8DSRrLWv7T7xUd+Y7b+qJQFlscLV88s4l
3HzR2837lsm6QdDYpCABt1YTI4HiTyUnvudAQE4V//S6Zl6Knmn/8XE9Co4c
N9a4nIV/ZZwY5QnIElvfrVHoUB6ofoN6TegY7i+EVSUgdGwMO65It5Sp4kGG
YF3OIrRGmzBLD/RT5A8+3raywzdmytgb8bJ/HhPtZ/m5hgQcGH8qxuE/KcHt
rBALljrHRDJeRLMMpSWOSzDyXDcOugoepEAfJ5Yhyc8IGH2PaaXWBJ41q5DX
KnAMSIfYM95HgdHshmaIzm+m+SRlVdiWLDUE1JJqVAJPHj4i98xoKmTl0faK
uJGbrTZ3UmO8ZcbGopQKsy+QuEndJocS/ApMwc3L8pFTLVAWBwtoHWepfLdY
Vl19VplsJBKNa8Nc0vd9BoJIuFAKfrS7CCLA7Z89GkKIRfHOzLfeqFsipeGb
iHrhs97V0/sxCwEV3KMuwgwStH5Msw8AYavItepSYH+AqobfkmpIeCuVeRwC
GGOCG5eAXrWZ2Bb3VkMqrGgcmH8SuSnj8zb2zUCjEwHkU5IJl/NdzjUkd9Ls
Z3HDtF5OjsIEFxtH4b71PgEwpAfQcp84b6Gk7XAB0lidR178LAyDU7eD83a/
sTJgn/ezgQIUvgMBcKexWezowk4CGYolGeNQ/yfmC08FNKQ46TNhg9yuLOL5
EgGQICgBrqnt0StL/3tDyHHn23JqCO4KoGL5hJ+cy3Pt4ZmS7sPkKdrH/XBp
kU1bZMFeaAFYbEmt3Rb3u/1iM+ypjAWbpISt17NsUlsfO4juc3U7i444VEKR
IN2zBOUvyV7zs2FxyGh5raQNnIv0PWTafN8DiRj/OlBXoj4IESaCZn9GGaaQ
am3kVgpTcN9Y+3S782Gde0kcRtg78kJD4ozRpfcwb+NPRrjzH5KJr6IGHaSU
2wmf2y3MozhNFMfM+c4lOcEPG/rjMHByaPQTdsIRSFoNarCP1L0/U7/KUtFY
D013Zds7EdJqhb8SsRuIXSaSUgCNNltgGP+4SSBwLA7et9qd+bsaKsc7AKwm
/wZpC2fax4mhzjPnRxqPiXubFEpEdQAN3I8fYKifvEoV0RmvFrkFfrnf1put
agP/5INT6M1e6pC2JEYqy9YpG4OeB2HQKQE4p5RYBoQEnawuKMRO2emZFuEQ
nxdE0yqUk/5dV++FAKlcuB86CYTjQGu7VPRlN9lSYQY2rFBULVhKFB7kpJ6o
yHX1sRGezhRB6rbNvETV0fruHOlqH0AX3Qtsi+B9INqzAdw3K/7X7E0pDVEG
BXk+sWOuEzF+w5P2sZIbDQ82y4y13QJiuNDhd7wPPi2HzzHIntU/Kq+YkFWG
FdZVo42RkYUAiMcXrQ22Hddk/3P+lnu8rBLnM2v3CsNLcHi1OUNMlNgftJMV
dco/ipPrNao9RZVCGHUe78wCY9sCIKeYfMmN9+bTlp3rzcaMLljCaI2gBsnt
Nmzc1tsus5KlYmU/yDy9bQfTHJyYlOc+itar+S4MnPJJ7KhiE7aY+jMX8JqB
xyIUyjc8fBXy2hl10q2xj9IpEYv+u1ohNRzWRKDTcInLhRhwRkpDbupU84Cw
gTHv2rQQp1iIbTz7WJMYawU6YeMtZQmI9OSkZK/QjPIFnL1PXZCFghEYhaD6
vPey6gW2MciBWL5PRE2/7jDK+MViHjwXMTUGLT/EH7/ZiPOZrQYd5a6599ff
IYD44mwFq+qUVhpPJsdB0MiInKcPZxg9YFzo96QmoZWLkX1MYCRjtjY1xiW3
6mgNQ8pyg03YT6QNQ/0/KCli5thkWeNfqp6um553nC8XL5wBFpxCFIOsrI7l
sltiZ7IFuxgewZRe1GVXEIuSAAfGK32MKfGlB6YCmAGnUl4eiq3YLunNIG+s
Ya+ON1m+tm/xPgiiORRay2na5nQ2eqp7dwDcPbMHPGy72QHLmmTkqm1PZj5N
Pp4ynvnJ9M5sjHHq4ZJhNro8hRHtVRqIo1TM9vx1g4W1nQ9xhlOP5XxKHsdk
Fnx9WC5irSv428CYjeyXQCTgjrSdY+0kw3SHTqTdILT8VBcOeGbBVniY2E7e
3xZwR/kNUWOVVrKzaq6RhNKD35DK+gWa+4rL5vYtRiXZR/D2PKMz3w/6dhsu
xlF80h9Z1wrftlwQIwDBBDQyzGARq6U04kIyVFa1kPaEbI8+HgBsIb+m0R5q
v5EvNAI8gv5fKts3wTkjgnaP8J6FDD2bjPz1in3ehUgONWPmCPsSMA2c20/b
o5KwoVocdTP00dzI6VWXx1B/Yj5F/4XiN86R9ERsCoL+pKeHQHCZqoGXhrv4
chLtSGn8vZCqCoCpt2os1RLxbkpC1nh/gEtuS5MmTEQTXVP7tGIuoq/oM/8w
pV4QNgdtwUSy3BadNDuBKC9kyeWtZd7H05N8APKFl37Sbj2UGyz3AKHmswRt
DdI83qsgVb7xsCfVcW5SGUGmDWwDNG4hoGS0Bb7Plk0OSRwardHb8oL4+7gi
D3zTeluyqENSlzTfzJ3pxShxyLcyVNZjjZssndU7M59h/m9ANpsfF0/l6bDN
zsnyTc6TT9TVrzHE6WuITm0HUWpKNEE6/xxPIsLXa/zZSnpSWGwn5WZoGpct
vIg8Tu+AevwCazLSXsqs5yC+5FbPbjgGgxNSEoGsFy9hSox0W1nAotyq+EIp
BrMpM7MKxMlmObKI+jW4l1CjV+8rQm+5MzKH8fbBCWvpFa4Cls4iMfMgg6Qy
jLQ70/doAHZke/ivuDvHghehFY9xu4DAon/K7ClhDRrgXh2Y8b8xcDlcru+Y
NBDsbVbx1Ya85uzh7yG8Yh4EEksd4JwhwJ6u+3E1lpC1QSTAwribPIJaF2ak
X6YXzVRxUqneBki6jpy5DWd7YwO0AvlS9EnRceIK8cuwC38utCK0qLGUdHMf
oAe4IcN0W3u07CkxZOyQkCXEHE5uIXv63jWQRX8KD7B++eh82WQ1DqoMpEGq
9bjBFLdKWhtqjYukjvbRCf7FoSXfbixylBDdKMLku7/k9WvLVt1Nd24M3Afp
zNI+LnJdeKnvjZ2G1RQ7LmQ4x8je0WyKiH1ZWmrmMbovabFBYBtRvlVMiH9e
5UEqFS9CLRCcYu/uFmpg4nQH+XPjqtqdQNgrOrmj56yhpjvqUb+ImK+einMz
UUSwH2JciVjelBI5Lc6nPd8nfBhSIKkpsZVB4Ir5hxHfwE16xfvgrF6+IyD6
JJvvMgJzrEz7Ig5b2qQ1s0TfORSfWCeKHPJfYkG9DFk9aSvTA5YtAc2ELN8D
uX+nbfJJ7WDtrofmL1o3RAHLdqPppHHbUS8japFKEVikBY6FB/9MvI/Ol6GS
Dlmfc6HgYNCNf77k3pa9ISIFQf8pYP/sqCH0yoNZTQWq0RtjAe22+jB4PD96
Hv0gnRW+wOAuEjymb89h1dFWKwPGErZ92WWfPUXi07Qvs8mj7gyL6SXtuYga
O05DpRKEnKBECmGMwWliFBnu2fZvPOqhjrAvajsHRiv6GcdMxVbe9l8eDouj
fnTX1WiUJwkvkdJei/P2k3WEOQVAnaP0EbqW4Gx/yubPMVawsdf11uWC2aMN
dhb/CfIZZWrfESxTZHK+I5uad3HP8ktI4Q74cnm2c3EUodIiuowoKTSsPrQx
DWnodYEsz5mv21YvCFT2pwaQEqLZPXfRdMwoStO36KYr6nzIpSUKnso5D/6r
8F1xq2eU5F2u7gkepCQIUuo0HRrbBhqfR1vq2VCZg7YTihxMDtkdlCtJVnow
FxD3XkBc7UbwA16yuCkLFZ9+Ji1Jj3Bqyq0EuakCiakBxstR8XFTcE2+1Qa3
XZXkKV1/bEsNKPpFlHAqGktflxzzBpGcgrn9+S0sqfrb/N+hV51pPFuUkird
nbsJU/TVVkZwQL2PA3zUZVYY2DmKrsnSOHnhytj6kONp/eQQ/o0PorkrZiOC
LocgczQLWRiLvWAxWGBN0CykDzddy4UQa1IMa19FfT7+AQcciUxeJBPhaiB+
n5ITH5CByu5Dt+N8hf1r3nJqPmo8iX8Nq76w8PtS7Re5O6Exi2UZGvvinFN5
rrWz0wcws1fcgieStEUhPtfPt2jigTqocRAPau3y64aYFLEbe88ukC+t18Ln
pqhXPs5EJ9F/xVkO8vMBTvBd3eGueCirpbsJCEi3UNhOB0er6XPmuEQgaHlD
kWeJ5I9KbyojK/+OAWJ9SrQTbggmEscRufOT7QD4kgKmJBQ0evpiFZmksYcd
1YgHL+vhhAS51TQdrPrDyMcVgSfmHKH/TEeuCOdknIFaqezsW0+xpF91XoJK
XfZN05CIydyntt0d0xzSwD0TjM6/pB0dV1PeA8K9580gQYqvX1fn1RS4u140
JFe1BhrmISRu3JfsDtmutT2Tl2fD+JNb2az2csNhyb/eRV9Ju6Ew6iyJoUlP
sgrbkl8cr4N2o79CNYmAE0MUAViLGhUyvDEvVQa70ndMqAB3+/eEybZFQQNt
F64rEPJ90+Gdqznq9oGav/Rggw6aAVUUCb6V/jDIq+GzrzXu/XGREUk00pVK
0spw1DgnNZqkq1+M8z34Ok0P8l/c3z0SuL4b+ebQD1xsLZkpRE2IBedp1bJb
LxfdBN0iQTa7rd8I4Wr7CBOm2Ijms0f0m/62BwpnVM3lzQLYfU3JNiXC1Szx
xmq3JbXhBwxNQACYIfdnKSud9+KOlWJ2O5nkRSJenKlPs4z3QPwxaFuMr7o8
f19pwjXCJaBMA4Yt6QVf4Khnx3c5dfmS/dvoNvcPXQXjk7g+PDK60Xy+8vB8
LvXCT4xQLnmw8MpX/hl1fVMaERlUepnLaLIh5mHYdzR6KzzELudX3lsfNkk3
CrYTnfkuzvRkVWCAJIV8qeT6UW1d4YlAGpdHp0YAbCBKNBD9f2kWpsdaSmez
ryIfmlNa+asnAU6j57OH5a1GBuLJ5j7KcVVL2OSOPAayrKdhidsvKoSnPexo
K5CeAkhbsnlsu4tOsjgJ5mo0uLRG53YRFcGOzykP/+Swy+Pjf8k4y2wUUXx9
XmqPLOp2leUSpcoUOCk84Sop+UsYppV8+4UVT2QSYPwLIGQ+azDrG0zuYxqg
ab4u68AaBQRV744F4SkusTZDkFMPvLAcnPEvTZG1Lvz3xzKC3TdnCzdf7jb9
PtRmhpKVBnGh8vWbqMptQCSFdNK/SIlvaW/ZDAFeJq8zbje0JlBS70wVXgQm
cbEqg1t0x62koar642RAGbyuPzgcEq9lu9pjGqfsDAgRZyzoV4CZXe0+AVL8
GtUCD1982f8G/EmQiIwThx9bH2gtsyEHEZxpwd+85Tuu+N+M+Tn+UNYP+Ho2
yMmUQ/L/F+MhMGiwcFDqYtZO3Lhv7fmzCNBh7OjONr2Xzpq8FIlbY35UqD9x
eCyLX8y8jkNWlqsF8vMqj4FbylYeygmzX4MbacG8n+DvgGmkwtvxWX2fkLUb
Jsi05IdN2vIe7u9IvjLQ2KQNcRjbi6apF3VE0Ezk5I0/SPIl/s8yHE/o4TDp
Yrlb0Q9KiEVizperQunAv7rrxUhamqWb8ytgzgcRvMiNMkVpUYW0XPzNw9vm
AXsSGRYP0ko5KQoCUtfoYs32nj5JsAW9KUCFctiMMrTjUJ5F/BGFRk2TdO/X
Ga0opIo3A6NW0I7RpLNYZkmTi0k3I1BMVMP0BgM7F+zr80PaN3vQqYN4+y/R
jg/0AqIO1kN9K/0L/XnWruFZM7oQ3A335/CDeb/HcuDVKMa1t88Yf51UQkPe
R8EChM7Zbu1MqSZ3FmlFkWAMyJmaYiyxhp22PVMlUnV7A5doSbtbTILae6pM
CIzm2mkACMd5rGbCKDowtuC2RM/KDoU5pVNz3aKGoYblytkqpSBP+s8DKrVQ
w5gDL2QTwkizoDwGBOws9KBTMoXE5hAfc9sNy5W5qd7eMkYg5xQQLityjOmV
6Rd4xm3n79JctwAUV4ESpN7LrweBLTkE6feBN5879mJa5cMyOrF/8a+0RhPD
jlw/9HxjVHjAs3y/rC5wS/i6Bw96B3ZeiZWvhJBICM8xVNGcNniH6v6EZ2ik
cceYN7cqJHJli4cMZ1sUnBCksbshWB8g52wH794RQjPMaJ8ors9Gl4aDGaO/
DEgAn5AFeheiwHlJikuMr8KgOekUxFES0MZ/kVJ3qrpq3ok9zdcHmRRyZ44A
2B1GAgLMPEz2RDrysWU+6TSr6xVkwXwu2GTXZk+/D0XOLGV4TUArp9PuV51O
x1Sr8r8KVzv1xqmdXg9ZsjSRJKdzvkgCgdKIy9F+/cKHa472tvDaYVe/ajbS
tfewQSbLqiE6VnlruSTsWHhXdT7MU96DmvdWm5jH0+dbw/wTsbBIMkfRha25
mIsgcpGGsmaXD7B+8iEXcR6HOyDdKrLFxLXTAjD0fySCs3qzo8pRZIzMhr1m
gGbnhLqZN4+FzTk4fRMDXoFMYUoI18GYJp2fzoNTLPUdq5zRhEryacXfJ5PZ
1wtN1EohAdiL8Z/SfzaIhvmgouytfW+i73ak26vrKqKhCrE7XNKNvhyVeMDK
ePrl9WOAD+3gvzJvAXYCFPcQcs9Xr7y1FlMzk9f39wQIxdLIIjrxa2xKayil
SyCsUZ2UeWdWM56D2AtrE7OyfXi0zV8nZeFDQ7Am4OB7mCuFSWEWbatjYqUJ
phFiic1voCcjthoGppgfVBE+dS/Fd6yCORhwjGCy0KAlf66t+iTBf/kQGnHq
MKJmMTSVVNgjzqbJ3LGlgV5X97T6CW8YSCmxyFIDHI7EhwnX/2vRyzj5ohkH
FpH/0rcjVvvd6JSZAt/I9I/XMcCvBZUYiOCMePhYvrGCbBWmfKgcI/hS/SGM
hgIrjK9dWWMDPZAY2Hul7a0mIwahlUguN8eAJAIGI7twy/3QUB+xCor+pK2B
phNe9a9//0AG6ecxtg31uzZDlKOdbDCZcsARe2/y2ZgsTroqZbKH3iwO1XND
wJG/HW58hs+555/vreMmrM0pL6RDPAihcZtEPpjRoASnJNoqqrZKxg6B0dug
/uPWVx3heFtKd5g2i+xSe4dNZMY6bIVBHb/st9KCzxUYf+EqRdVONfawICiG
mGk0SMaFZJ4R+ijardqhHjn+KyIIMnqMjiCjRYjheazAqYekXmixkf6PGkPU
WPqhR4HDC7Zv5CZZeUePWpuNOT5EFj2jOBVueaNrt1FAkaOSAkvA4zmf0cC+
f7XP7O0qimuxvztCK54T+USSscnKAEDqgbf4aTehHm1wVmTZFPa1xVSeKCo4
YV+C6yKyapdt/dyRP/D01B2zxX5WuHg9yZgu5UJDjuiPzu5Ph52DqVgc3jrA
lDl5jJgs1gO43VfTVSbLpshCORwFsR2To3rsO54cYo/G3xOTXdU/xxej+Wwu
6afpVl+/26tn173r5e6oYf4XllYBdrrUNo1LxSg1zrCuhxiau2/5aP2fqRDX
KXIkrxbpVWvslcJqPAM7EcH8EGCmZaCUoGe1OJZYT6DB95cadAUvLcL3TeRD
v0HBnWcG5w2udFHsAX+eUsdZJhQQLPWRrIRM2Kvy6twpjW850ttWibTCwcGL
6cz8tB/mJy68UxoR0e+K19awjLKrwgv9sNyEPIoiXsoBIJg+cMy3ui9w3f8X
Rso1HtpErvkTfD8Z0REv65KUAumkIrgbSDRLkLhLrgG1+JBaWbAQ95SpJAta
6cjHJ8BZriMlDHaBb7H+WHZOSAjJfIj/bLimucNrZQ0DJFvh9cEZZOs2SiAS
1t0+2MyR14crStMPAfNy6KZ7Y1GctX9a/dq2mwczMgZfTh5uWAXMvCW3vdEk
RgkKFjcV1h9ML67Pj63+WKtU9mUATLCrdqOjlGlCbPp90H+tbgtb+wMQW5IN
3ZwlPbhjkxu2TTOg1UyGFK2v/EBCZDZ+u29ItTLovcvGFFRtP6DvP2lGCYwN
bbv9uU5Tyn17iCRGJJZYDtTTThol7gv0Rcg8OlMGqk10mRP+zXPt7gxh+5IT
b9DWktSTmIa3oBzbGNhW505YMjiB56rYiK0SBfgvTDIOfExYfURSX2TZSCAg
/B8Xlj7qw4dwTPi3nXEqumiDYI8TmhIHM5Gozm3/2J3dfFBTrNIY8v3GUUOH
pSyKZiufwXG09UEHHCZOleUR6oG6QaBIVQIU6k63ezouWtJPB5m/XwI39wdU
9HPIOERS9mqgaPmpU5WA26eshxAbBGxFia9LB35heaaYCVAV8uTb8ZQq76rT
vB/U7s3vaqieM/NRrjv4C2YdY8b6umoK/q3zyGPPBmQBMi/WA0Z+8N7c9+Gg
Aosykz94j4+YdJLQSGQvcTfmfNwC/oB2P1ek33n23A8gBup3LzkYbvEZP1Ws
aZVS5c9BHcwqrpgmlReVfg508q7sNm6MmOeczXOLxCtz/P6d7wwpotyw2fBR
l5gI7CRDjwsQApt2b8N8j5cJzM4UVV5BtSZTA26XEB0jW+QuFhUpQgQ9oVfA
Lk/mjtHMrbtQis5eC1m/R/wCCyl+twYABdqmMfeOzB41lfbbIv667e/VZIh7
JyDdNlzygYsUaWbFV25kOAW1fuiYztXF/TrDc82w4vFzVboa4iUJgeK3fusY
MHuE1Hb+3RIj4QAIvCWmBQAXQKVHA8tG23Big29bIJdUXL2GwlH9z3Z3NNq4
0cFM7ChpB107FHf4Owk5Lv+U3WWMCxciBM7cyMRDw4g72Lz0I2C+GjhL1pSq
cS984tzay2YtQv7jpb2Zy1IYxAkSuq6wh+Ia6vkEv6BO49zkw0taqYgWCsgJ
e84fS9r6RxgzpHM4GsQtUI6b2MlIGjMDlJQsQfx4sgAKXzctFbl70ZRexsPZ
e4S9bPwdNM0zDB4Qeo93qk0gdaR4WQ/1AHDAuPjkyg3j6uDRHwB1zHztaRfX
Ady2ZslBTWxYrGLnY5SxAmca02FZTqiZpHMnrwbrCczTuiA1EMlGpPwXq7BO
SR5a0iPpjtzNLKtl+Y2AfsP3inoQqNq6C2sfCogqHimP666PYBLHx3SU7Av5
pEOa4I0xXeDkwmKnEp2ZCOS3IHhba1BpbENpxXxZ1cf/Zubun1vLmy4ejzdk
B5eu2LVHZtEsu8PbPqA2fXsUx5AYNVnCHhmC2Ld+SEDi5Nr4lIYpZUcWikpT
B3UH6KWHBpZKzVtc69kGVxu8baQv+yQ3WuDbUbSTMLZPCLt14ea7UaYSIs5C
0LkPg/YFqFPsNRowm2G3l5BEaEmC6icloAOPXd47Jqu2RKWarEezjG+0prVT
Sxs3ZjACGyZbWOwSGJYApycv6AcfWp68J6Qmf8AGyhTPwM4zjsXPg42ERMq7
jWFTfuBfTvDsrUvnljGc+grXHl1HFNfQX8Ok8Jfvo6dUVv31do3jJKCaAp+L
YcFmxSp+oSLqvq0v4yZi1K2HlY022TVVm4y/ppZeXmwa+Y9pAq5+pm4Do1fZ
/ZbmMtGCznXMVdgcA97bH+CJPAymOeLDmxBvRG/1U/erKL7BXIyfL4o22FBB
X6iJqy+YOmFbSckSVPZCUUw+/Y58fn7SeBq+ZdYQ4XeM6on7yMd15+5pcjeC
tUlnTftioDJtdK2kkSk78BONi6ndKMdYXa9dFrCrx8n9+MlxcLMyHHpU0eYy
B8Q/D3UqBCV2Lw5531/oG4p1aQj9kleqfuNedJRj6AisdSs8/Gly4YpNUv+/
aPezFdzVq3YZTlPgNNhB43qBRc4zCOkEgYsKxo3qoGaLTieZyUGCkTlvWwGe
FVoS8NXsX8LIMz7qQkl0pidn1OXVjru+7PATPna22S9MHO/a3bh1VcVekggl
AVkV3vVLHBGffDMrwGQpZf3SN4VwbV4Q5fF734f/c5gVn5ScKB0eFCn36Jdh
ZTkEvDDhBge8NnyoFSLQwQr+Tu8sHn+HFQqhkW6XdYCUFmx5GGRtA2rqYtBv
DGooc/TovzLDusXlRmDLT5iSvLFtuK8TGJ8cCVaVfX0vxjd7lofKeCKHm1Ve
yDtf1oWWwxQarMHRy8qi++qoUS+jWkTKS/fnXMCl+8n4tEfBoltCDp6hvBn8
4BmefnY71eh705mnGKNMCM/a/m9t9AdytjvM32AwZRPUpT+h+8dafDrxQ1Pl
ztJSN34zoiqF2hSavCmUdvCCS9qqb+rN7TL3bQR6EWlvCPNk0Yfv005eZMEl
3NX/tNhNgOliibfsUCZhHNbgcKMpPlWcZ/I0hqhqL2bvtD2X3/MQrQMlc8Wq
T1EYNWYHLW3hf97QKXqQ7ZkxYmrvj0KhnUpN8rFUYD143yRtt81KDFSI6nJ2
vAlyCQNrjIgotIUWnxcAU6Dx+vKxIys6I+u5Cm1IJOSedj1OoBNbUGAerb4f
5tWotm4YVK/ZBMR4w7e1xYYQRKBrl4QH8wm4p6HSobcEqER9Bi925PC5FFXm
StljMe5EFK/mnKQ/zy1+ldLOgiz9kJgY/NF7/HpklbPFVOpobxP+zHX6jHyj
PI9Qp10LnKCEzSpAzN7Io378piKjyhai1kHL7NQ4wvRLW7Gx2yAsIK0QR9i7
S2hERbbfGf0aYm+DuOKAUCo2m3nO1WqVQtsoTy7Ga7ZstVLV9ppy/Z3fzvOx
XTO4UKnN1hWwEwYl7SE55+OLZfAmA57J80jEfUc40IL4X2CcoDIs7NJJUCRF
y11aHlUtpqpRp//9Aaid6UQxORzo/JZCVoTh5+19yzAFMtNJh9+a6hh13K5K
Mvmfgk83ZrLSwuOXfBNCfAsrB1IBifU/OWp00d5nRwo98FvzeU84QIi4ZeBI
yBnuvIpGDwmcc8vrE1HzOYYfgugyjtLDJq50XKqDWM9WhuIexNPxow1kJlOq
3HAQefdW0RBUpI/P93MV2bN3NZxnO4IFUs8VtsxXl9+vS3AV0u458umNMQJE
SPfGm46Ro/2/kO1vSFSHODw9c15fvGaw6m6IB88jzQ9ItxOSSETC7uRjqBWA
gtDFbjN2rmt9w4gP3NJe98+AsGodqJpEOva12L7bxxodbXF5LB1JJ1N3guXP
vpMYCFmzBNMq3rgmdmyJ3pQUAh330HS7yidHA0S/Vp4+VZ3FNg8jGBugEVJp
JXdGUl5dGuUp6Qu9sYGSu6jZY3UnovzY3aLAQ+WB5D11uip2P9xNboAH2aho
5VE+8JybH0d26uWHVOYLRYwkFujR6JI1cYCTzehbLBxonpe2fDxXhajbb3Hg
k/GP9bCKMTz566YK0if44CY9opT8Hx9di/FwRSGgrZBZSRbNCr5bHVxaU1wC
RufOMJ83Cm9CYcj44AV34ESTkqJM3tG+/+aUAWqJCyzNrWzHYg1mmkcaaJz5
W3fMzsxBma7a7/aDhr5sXKVjy9g42QVpEu9av/pT4rCSvtrWFC6A9ibROLi4
w/sJZI5mZzBRPz3lIb10TfeVaIYvBF5CWtJFUWK1wShpTS52OtwBDTvS+1Fs
TwIfyOoN0p6weR6lgfogmIJiQyxq43Y5oeVY7y2O6v14bu8WzywodZ8Hv2/e
4Lzm0Wap/CgdXtvLTXvKfirsPTxLfWsiG4liCzG67PK0SrqiRbVr0aJMSiik
tXwIh41Rm1Q+dz6glNmQdgeF7yLkUOLQ/Gfn0FBnMYDaguJN0yTm+4J7qBAO
mlHhHkGvBqM0fBf1Zib4gfB6oEvtSycCLFopND+0GKa9Ws0rbYdNvqJXtof8
9N6l/TFHZh8ua/uT+h3nMInHaRucrUW/LymQKxqIhS/iMfYApqxDTK3dztVh
gjJ31xjAaPdr1SQ8xxotccO6XJHFT0JLbQD3gGjX+SCdXOvP+CYRvbYmn5t1
dlaCJGc89uz+xj2/R7duNz3RH9fKKu5fcPp1RETmdif9j/BW8VQDO0BuOZ4y
E1d5JkNLZZ5hdoPD6Syeq0khi4UchtTW93asuP4yJNc0+lvKIhOBwIxMGI6U
rHFlsGNtzityM4jZG25CSWiyDwVdEaTGyS9DMMdndrbANM0OjhuJvVR9O8lr
of0Cu4d52gSIdFQS12FxF87rjrgJM8P5qLm6PwOrsjVIii9bs8sDiE6TPhkW
ZIZ6KVc/6l/FzaE0qA/GWEp3kVc2Un94/8QCk6M5Nan9kfOy+b0ZwwCfM0pa
Scs7lp/v/vdrDy43wuo2GjPNWEZRfQxAbnfgabY7zFwM3lOF8Dk0vV7R3lxW
/ziFIEY4bQ788UNoaeEuv27LtNNWBm0KywMyVZ4I1Orw+t8byTcvDDBoGVa+
6N4DjELM/FCcQzTMEtZeK7NRG9EsbHoj0myXDCZ8gzvxlIxICozLvUSkJWPQ
GmVZCbyGCw/DJEdnyAlxSLjdtPkSgbw8o9QLrQQiTwVMqyVehBQ4n+o/AgtH
AvTY6ukODORpThD7/o9oYDxV1uIWwIDu0FTrXoOKf2+JOta9gavE0G4tNWlk
W9KbkH1Ie0NSalnwwT52dQaZldg3sJA6RsEpgUidg3kDilU0h38EG/RmJwrS
2wEeFPPHHmEjua1Wx0OWdHxlUWFLFIPHguZetumJTAwXz2JwYdG3O4gJEI4e
3fcgHE7So89OYxJG2HEv7rBiPiZ4oaEUck4b/+fdvo5MZYK4znAYL/alhi61
aY9z/t3fxwrhqWFm2WDWGXBIBemxS5hL9R+9Juogf0s8ndRi85/coHn6OcMy
5rmu2MozZblnKBuc8uTDUsdGiAA2r8uZE22WGpj/eRro3fa5PohpmNiIgrY6
6eWxg4hNHqf6zcpzKUT6OgFhmtrrOCpbQVrvbvmFwTLiad8lcUgknVn+fJDQ
3W+7CB6WoKN224w5Bsgsxpi/HPFqvqiYxomf7yDXbfcLCAjwbXrXCOsxp5v9
VtZtigvFJy9PvPMOuWAmNuT4h5EZ/F+VLDNIXOWFXgc6tjHhnK6zHjWWMR0x
3HQJo1PqHtG4OopwXCFjsOCsv8uVuf0SboORU/ct3KAYDSRj58Tk3B6gRfXo
3PFSDkG7HIh8KTDH4L2781jTbfgMIzNHZb1KVudpZU0+evN5hc5b7YBUbYK7
3ABN/b08yiBJvzaruwxCnEsnLRZLdrueQYm2D/O1H/rkl16byzSBZqwBB8ea
PkZgWapqPRJnXR5HV3LaAhaJz/lSEDRlQRZiy4GLGyHPHE6FEjvheet+mLT7
ZeI2O9wiTEGUrf1fhBNs8yFM2Ax6LjIiFevLFmVE120kxSxG3J8oFRUfspmW
kUJdVc0HeOgDfFBBcOlPUbOWsP6gXoTwW0dBSSIvzQvfQm5BtiA2eMC4heIc
CRmpXmvxLhBNfeITf9K1awhWkO7iyWIcXcASd4kliDItlA9niujUgdRnuzoI
fiMgJB9toefwNptJcDH02TrQvf3pQJogH0JeDXuEi5jiXqr+D0z/ZrcsDcU/
AqBZvkZNErJ8daVtW0D1PoKoPw+/bscEME/ZCm+JTtPa1pqCWZRz8br6f8+e
EJ4pDf4pkl3C6s6UDkHfVigkrAVGNVOfMZ+Hdw8KMYLLYx5GtJD1V6UW1mXo
vdFQ/tslVtrWZ+2NDPVvJjyQdGXaX27gxWAChjKjpxXA1cqAt4n2y4yJfq9b
vhcaGyjrM42XdF0laBrifGBr+i2MEfRlp5aFl4wzzDaOzBNFNEV5xMosXl4W
jPKZ+RoQSWw7vUyRBW3x0aUdRR4qXLqJowNxNSZcbwuRl71Q3NJ8WpzHnmQX
Lr5hh9SoQPTfPpps+dHcQaf2tuc2VuBcgBBF9GKGSZzpRavi1Ck1+7wtCy0w
xDAtlSGtmMqxwD9mazjIb6nRgiL0fmkFa+slRTw8diS3Hvp28qbrP7kZxEZb
CRAhUkmf8tYBw6V8Q9timxqofPL3WRYUc/oGqa32hHWpirNRfctyJaCXrDPp
0H7cO8v7+e0mYRtjva7fqmPdVuhnoVM7yQjL8K3KdK+PrWWNO4TeD0QFUkg/
cuWi5Sg9t2iQwrwUSWRmazE7GOeF89C+fVYgZ/pyRHYBSTgJeVUE51fL7Gq0
VtuMVy7BbDX9+F6HQupucf5lGe6uTGG1q9v+1kj1AOg8W32Aa/RFiVpOvvlp
Q9X1t2fifAMtUfrEq/9TuNRZc0Y6p1woEVSdNYtZJHLqbmUzoMWBDfOE7zSh
KZ3AvdKCLPx0o0mK5KS2X2DIF9LGNwRNSdetlHjKZg1U+WX1uah0mGvPtVTp
YCDQxQggn1LMTK3FZocNQGsQnhEUYg1dODsGZnpCqljfosGlvh0XFnKfoExR
u6Xh4reWWKWhLfMIMlPdJ60QdLNny7G/vZbLexhF6y8UXH02qFqay6zPgkJZ
oYKtL6yoby9GofW1h7V/NHthIpO9XTWu1vJMp7W95sjJq8h9mPn/LsVswuL5
hFV3bdVFwvPkIFYgnE45U+nU0x7lThsg0r6qZNIOBU8GKk+juuZkp/IMVC27
r+7YLy+w7LHqvPpore8WV96SYagCbQFqScqyXc+nMDMt3uA+bL/3ZWqrRln7
mW6Oz/NjkWfcI5qPPCm/K+GfGpPpIpopT5YKyg/2sklHYEJmiJ6ZwcSJ97uj
N1+9GuXUB5H7V6dKuG2mggrnj+A50UuIocDQ+HvEOuHj7YyTt/l+4lvrpqVR
QcESblhsr8Bfzbapdhfft+9W/Xr5dD4WUGruRG+CNPJX+DUDppbb4ou96NsM
tU7urfA9zW1GVtL8hNMcMpLqS5DPJzsSoOuLkk42ozPZUk5ysaCXShz6Ju6Z
sLv9UUsTHOvEJPRKoNdKBQ7ibU3N5Gkbbi2SL5K3nHd/nPEickDBnnYmhjIF
ANctkGEM6QDKTsxrfpEYjRAQBNHerIWAqy7uS0R4ADbcBABR

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzeqTjf3RctLbJHvV47Ssn9hX//GEc2QgiFtBR6RnFGdYUKzsRUuQpkCz+B2qmkNyw3kPCkkqT1fwiRcLeascQSWI0a1yMhJLNDc7ZWosRh2oxpNNrUcAXjeXgC/hrtpM2AODv1SFghXWiekxGenmoYZXq06gR///gnokg2+D3ZSf9oSe0KEdjcuAhnv/zY3YRVQsSIax9B0294qCfU4+ragTjW5YDlKrpDKyazw1zvJt/vJTKt+oZQRhH0SLD7jgIQ8oR4Rq14BWwJ0gfoGPm6SsDFVmlbBw+f1tLCMSErgLbMsv3vH4mC/Q5E0YThWco4SvPrkfrmuOyWe0BGwfqErhlNnhjCUqaUsiHMgJdMr2mYdlFGDMcox8AoHao9rl/R8KXvF7lXDQeja8Ow/2Zr6uHFC/oIxnnA1AeGB2plCtOxiu7M1mS2pVgOkrZ8S5LSRvX7F7wPrlPPSbZPihS2QH1iZOoSwyVHbXo9OJJlcyiidfqCNmAol8MgeTs79SuAucJQp6NPK5LwcTcXM5Pn3vYZWAplpzzXSvqvcX4qhhp8OJosHNOqT7HEtwxXiHC8+nX+tLzO8zKUP4mHPJvfN7qs8jED3tfq7XBPo487GxR0Jz681p/gwU8AmzE/KMbnO1aGkwIZ+eSlxSfmek7k0jjShOEY3YHm+kXQ0EB9JF5xeZI9Qs/IKw5wFo3H9mh42hkpjBP8D2pZHkJ6guUURseRJYacXDBrEm+lsxnBhXhn3O/WXHgES3M6cl6oGCO13mBqoDfK6bM1iZCOLpzST"
`endif