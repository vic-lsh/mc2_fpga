// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VauNi+juvtxgQrL5jkbXrFWXXBXFw8dHnBpVcO2yTzDZspI6fId01DU3DWk4
+9y9dYVt7cFU6sBI71ZY2kp3ifjKeI950Ppd0/tjUzCF3vCsYo1ao0alYJKo
+FeY/nvvHIPlFsed7xyM+/d+0R9DTE5ht26541HHhJz1Y9TLmBTz7CuaA0OF
mEfxTeJ5xQOAVLoCTrSqv3RUshIy2btoCbLmaiDe5+iR+qXT2oKw/hpdSUlF
vUTa0bd1FM76151rL20wx6IBmE8XKhlsz9HetaAlCxYIaNIT19QgTuhSVcVZ
2aAU7Oet4BDTLURY9mNSC45XYUlVsluI+b8VbGtPwQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y4Q9gtRpBxn9q5jXJw3jAeidxM1p6KNEGNMj3SVr/klETJNl9HKzDiaedr4l
qnwvZyZJ+zBEGt79re02ZQlTUgCw/7Pc+XzX6nlURr8CASapAQ7MeugFc2UK
QDRb5jbeVfmnbrQrEv9Tlu97pt0NqFlWUexC0HOB7MKwKSrJjm8nCr6lAHtJ
nL3DoGSSE3BB4uIWnCEqle56PqX5ulkCqRsQeKRmBxjSLdTsYzJFcZbtt+k6
gV2dMSh9ON7f/suhXUKV6ZbghzI+8xeYRrUpH0duPN6fkKveN8XS0NzUPCnZ
HSLiEFukFLj73LCKvios5gNDoCOpq6KpKJesN62KnQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RvMngiLmHer2/zjun5VDV+mHn3eLZuUCuB/0pburZ1RAE0u9+fwa/bKE8drN
YGhEfAy+dKBTcOEuL56bEzd1o5UrQNfDAzeyz+aRc2iNG3C90Xkm9B9edVmY
QuHMzr4nJGwjguAzdr6oYFveFpflOJAk51D6awxnmBBoc67pYO3bK8uAieHG
OVVRyPryoxGMYfIku0YRf7jE3kx4o9Sbu9FWuiQzMF80axT1IHfp25muJ5nG
1gJDARew2tEySyphOBO2xL5xdrHmngZpqDLIO85mNrAeK1rZW7y9wo3DUuAI
53uQia9B6kEEm8oELVxgs8eIPBqjm/xD1kjLVjPJjQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qLXw8qutWT70nUCXXKPuGd2mPrSeCD/xb4j0IPMxv7eLcbMi9hIC3FfQQ4DP
ZQbGi9i5vjKglAsWMfHJSb/IaSU+76L6ALJ7sLN9yHEUNnOQetWnwvMuzCUK
4jjmN5JPuEE8twDW1ZcMNI77/DLSAcyTIPJ/1iN5KdKdhSw/Vc1adyIunk5B
ZFjtJYKMpP4B3j7LOhqFXlpCHRIQuqdXY+7jSUVColozxJXw5r9cxtmzt52U
8asKhTUKpU4CA7P0Rjif6pQXleQPFd2hs3U5lPLTG4JYDbEYxfecGvxIpA9N
itn0gGFdBIj6ygQ/EJ99f7+bIBTRkBTIMONzk5a/cw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B8wfDUYH5ju9B5bSSBipQTtwBHoOmTQPlc8SnlSqCUEU5RhWNEZgcf81LXD0
A2V615tXRNK/Nh7JtG6yyNUmBCvW2DL9ePDeOT31YoFwnKNbjuTCw9hHUDO6
7iSnLZls7S1SJSgw1jM6Xj7HQyoF7xoBePR5F5HgjMqQu3JtRl4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MWJbg+0G3Aipivx6CWM/Ppot7SuhkiMjx643CjGlTt5Uc3Of+RngA0D2Vak9
mFm2VDHaAlY3rY5ut1yVplIYnCTeqwli+tP6X1yrAYiXVW1LJf6fPcOwjtP5
p83FFQNXiYXBSPMw3wj1IBtU1QVqFFgNpyGOa5vrz91CqG+zOiU26KWIkyXu
u8cqNcUXc71BhvFB/soSvajUJ6JCIMrfH4JsbmBw1o6+HTe5T83iTF1lsgxI
1JO6h2ZAV4Qt3L5Vd58gdru4PKujyPCgAdXIfCNo5u1eX3kbEd9VHtDfQMGG
q/1W48UjlGJMkV693UnqQpcJDclz/k9IYzNZgCQU393+CzTVreqQzddeF1+x
Y4iiE6pp6rDZL13UH0KUwgEPzjVzgrTAk2yXzQvOsLuiSiPIqyQOz7tWhJJz
PVQaJC8sWxvYVvXiOukTUX+wmYh8oguwmgmjj/w6MKdmV0oXkBbdGMeJop5e
7qk1ysjzYnzzY2KBwer9PgctnpdHk/ye


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kQj9SLNw3+6cVutmgIK/XQecjJfoB8zppjCNu5tjFJvXcf9gKRZ8r66jpOgX
SeDKUbc3ONy9KtGksNmFk54ktIVSRyF49u54LxA6w9vTEuDJqFMlk1sYD0SO
TIqo9gRpAM4Y0iuuJbluovDJ7gQOBtbHrLzuoPTx5YSc4rTLvWQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Bct+N7vsI6iB5E0DoXunxlFd+9u2PeOD9GWMrDF9ConcZbKl1WhvsjbxL9Ed
r3HBPnb0sPeD4+NPVgv3uqpYg5/KjE+dSjJHZTL0Jl2YT1QeWXeaG6m007lu
gvwb4FpdWYQy/4sh1SQrmph29+5dzFkPhH3VT8T7ksa97c5flA0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 689456)
`pragma protect data_block
I4/KEH33KAWk0CreXKoDlpb158kCCoHuYJ22sfZp+pSPjPc1vX4NiEhZa4v7
ep7yAnShzX89aUsq9Fqr6lm97mglSx21vY8iyKF6LOThTwKKjU+Oq8J0yQao
SCEo0SPLfNq+wuznjh8xltpVYDLPnz6QyWk1j/axZkNHXsAN+H9Q9lJldxKC
7w0mwiPNeRsggT32vMLSoc+yccM39dNyScjqRe/O5eIiw7LChEFrJ8hJ1L1Z
xsupLGAxv/Ri/W08/OS1L0Tnmozc82KXfBhHSY+kcoi7LLsFolAs3kdgCWnS
SnP+rsmaWfCn7IC9brZLE/aa3PG+fX7XzgBhMBGRQUJyuPKj0YYJnujNS+0J
TBeyJXSsyuGTtW3zvE+gljhvg/oj+cY6mN7FIKnvUd6HDQ5SF1wiSBKL1C1l
sjzfcuCLN6xcDujxUbo7mhzTW16J5+wp6CgibMC1nabXnjQeQE3cF5fVS3Ve
f3d/gcmakKH5c/gkoVONxM8Ht03+iQpvqlODhBa4J+0XjQWKW8BcymKb2k6q
nwbPPzEmLHxF+xwrYU3sgFCVledQoaucv17LFGCUQPDDZWuVKGL3IxHcr8+Z
lt5hfK/c3bRY9yaOH1mK7buBZAHmiLeGCzUOPGSWddwlpStewK6JF1tl/u3z
rKbynXz1I+aqb7CZTSSmLZF2loUYtulV53P56iUWjj5xX/gmO8x/SQ90M6MN
U+N1siplJetsS7yj9OaklsVkpyj3848cF4AwGsIfcxGR1Khqsca2ngs2xcDV
okFPH8DX9kVbjbf7/3AR3/gUjdFIeYdJMcVOec1YggWMi7SXfiE8UkpBUDd2
kmuRXJhrkrIs4mDV+Qs9Xuy124FYf3GBqRkhOKKo7B0VDxRa1Ri3iupp26O3
J3AYn05GcLdxM8HoyCRMtytbXsLivcbB2lhS3aWB07+fg2nS+7A2tVaR0YbF
m5oLxPc7pGxxQukgKVhFyLdEgiC6gMyPwolp5tV6WMeq8/a64xVr6mjD6PwS
XvVTyUQNeUki+JJOm3wtA3F4WILU+vkryFGpZXO8IMvSmmaPwFBs1P8TtXkn
wmTkik5nDoe4WN/aCAI6DX6gjqhMf/9qaMRDRNx46s/RnKN84fHleX7ho8Dv
OfM99EO6UEHjzYaSObyVIxnlU/8qXut1vUi/QmEhh0zKyKpWn3H2jIVTjFvv
R2pO46aqMeHIdfoK2zLu45zVkFnht4u+dt4e/1DfnvbEp6JOvX5tmFSm6p99
SIKeOsW9udzFp1A3+uok10isl/71tjAagloA8NB2EtkA/EWAtLbPWQ6t7fRd
fwqqLhXp4O/R8Q4J3eL67Rs+AWNyuR5OgUAThoK7BelSHygOeNPbdoh96SfN
4duNJEzd3ynqmCRZ9e3+wMDcojyJ50PpCsoR1xyCsodAEN2oSKiFhiVrDyCR
XnlAZAO/x8cbJnT95ouW33HDK0V+RyMN0GmQAH4jD22JnoPW/oekSqHjq7H1
tO0Fq94iqrVsJF3VL0bBGTZcD4+/yUEKSnpm9AwP5TGc4m0ShywxfGPhqfXN
WLSHQ8xi60Ermvr+XW+fN2tSdKH9cYz0RKpjjugaxdbBg+FPR9iGHYzJ0Qjm
khK8ltnubeA1UT2Hp+lKGLIxOkVXz8XuGY04pSrKrj562+HBW/cN5BkqrFOl
JlC/UzPTn79qQjdTPge0KRonj3S5RZgNtOyLHgz3yVwGfZlpwRhmXKB4EgqO
ZacBiVIabrDb3PRO8QRM7Ow9YvtoivGGkKd2Mp209dnVmCyt3nAsVANjbW+H
hyKMHpymhx0l7hAFlKuypCp08J8V78UsoZbDfImHW4rKB3uuNt5xj4/KMZa1
eTCixT2tuGmCPVuClUSAuqZdyPkrGoQbLh8aj16Dtg9r6XDW3qOsZaawjc1X
dF55ixE6CayOTStUP5Vo5+kkVeEOXu4s3FSDKepe7Hw1O/8WnMifEC/vL5NX
kJQeDVy1110hvhujs2cBfD83k2KGGtGsQOdcrJsqTqvA4yqK9EEWjvlVbICs
dXdpFma1H7YJVPHV3VMtVAvWoR+O/d7TI8Uw9ytpyrk25OmMpjBAMphFwJ5B
oaRm6FuCi0l9NyK0uiWj28qWamFfbCb/4CRTaxjKU3q/2GQS9tJbSg+YP+M1
rlyhTWl+yNz5XszTl8+qF73DBeANm/k+QSb/FwBLOgy8gLFSTbcmLQhfNXfc
xli4XbzXC8lIwhtfZj4IDDOgPqTwYpjkgsSqAkWK8A8V7za0EgWtPQBgfo9I
+fFuBYWHEVatP7DdBABTkTcQX4641SP+DEenLdak6xJSha09jbEBJLGoo/Xq
/8Bd5dY3KjWup2UfC87JRB+Drql9l70Ah+qCJb/QSFGtkx3HezfJ9kqFnsyW
efC1UMOyvCyrRyEb7trctQ/Nc4Lli4CcRfg5rgxkQ9Tgfymvaaramm0PjvOy
/mFI8KDyh0DcUc+PNvUj/SeDwM41d0vsbLjiJB3232qSoZqkkG9OEmvASnlJ
/DROdc10UgeTr/LM14wrc6nqAWjxof0ZEVE4U+TrmyHbjcFiSadQj4Au20Nc
TqmZChGRyfA8BTGvRACPF0/FsobVZZnEL//DasY32hFXWFT/o0gAevq/OW7n
bisoR8yLcmytMBXPhZmaErYs5csC5gfOHRpKicFcYxQVmJwnLcGiJnYtlxMj
hoi67/4J67MEPCYOy6/EgKWfL5KuSkwl1nijKt4IZtru/eqtB32WTMMg/GbD
uzOzcYdvdw+IP/X7dh/t6hRo+Gso3+vKOksfGuptiRsa35S83LvRt5wxJjkx
vwiqx2CPLfdtny9KiuV72d7dSDJHsBpcHHRoL08z/49IBui65Ksu179JxuAN
bmvMcU5+D6ccSaxvJ4Ep246fUNsIsWBSt54hkeWDX6dsw/xG3fA7QXRdjvcV
Ek4Mc8b59sx5D5/+RzT9A1WxazdqGh8g1hwWvLEezB9MyjueXSRVrt9IrGqs
zAgPjeahfwpd9sAR6jrlebRZl3899BNy1MJk3F6VDySBpXTJ955XpuS0ML+v
zPYDy9CTDjqpH/loeFG9eBD2QaA/bzlRQaMFT43HLDblIvDJJ4eovJQvdE4F
v3/lzrTbIrs/pCeRa9a4RF0XgogiIq6ajZ5oJUYYycaKE8f6gwBvOIOPHu6F
DxmF3udXr3Yxm0d0sxEJfR8vZ80py7T/uamtjfH/G+Ax+IKpYQ1mdTG0zhzF
PfNRvEZV+4qV643ownTvj9MB3ZQDbJ9kGxASA+AIYR+GUMu/C//r+desGVSq
QyMU13LIBeySHtenZV9fpV0I/tJdI8NQAhitJT20SvVv4l15ZGimUjDZ55JM
JSJ6KfbIOSKqEJeEt7lRz29fWj5y37d8XWbtJmzlvV+Y04AqAOcbayo6cvvf
wq/l/LUbto6PIoHFCipP7+EixCbUcfzl8xG/JKoiezs4X60aRA6jWjjwALPb
5rSJcEcNkNYL0CtdfiQugG5h1CsokIhM3EOh7+QhIp7ZabNAsLNCfh+MpnVd
qO4VjwdwwEPor3hZ3y1bVoR1E/Ec3j25lgDjk10VXgZw3/PBrDU/jMExi1pg
EPbSHE+RTb78SkGOX9RPKtYYKIJ2VR76N0HqFxfUtUDpPoq5mWBt1QbaBJfR
zkycSo7W50wDuLHpmT+a1EVKgbuBd3NLq7gD4OHRPTuo+jbjb83yFAbHBNlA
Xt5G0sceaNR4hx1Irkgf2nBqEnLRS4Z7ZGbQ3JvjwtCaKMOj9G7pailcb1R5
26rNnC/HwazY121UO421nAM4HjdEP43t0PH7NOhBJkAAF4x/tj2M0xulsTBd
BYmXRQN1ZfbQBCQ2yREE9XNaq3O3g0VTHMCYvNHAYMO+Hv/dAlfU1tOadbzh
2/HYFYv4iBlB7H9hPezU3C//5pktLtNKYPrA563WsPSxOKKAK0xPFXA+w0Ih
yGZjrUTeS5+/QQTSRyXNReXftFCrx1O0f3cVs3CwN0cgast9eIGDZAtUQsEH
dT95UyvHVJlS0Z6HceUVXH057kM61RH5X1t71nlrJAiBqzYkZFeX5Aw5AqKI
TTpVSV52OT6I/q5HebIijeZvvbofYFbybEqyZ03c7V8MHcZehcjnoqxMHXJb
5PtISP/edFrhFieIivW8u8zeNgkHQ8LGu6IeLwx/mTz1X/QVcJutyrgES+XC
18RkyEetUitjVhU4B2NUKW4h58eFR0Ag82nLTQGgrjU1tAa0FwmT3GWik7hi
03nBP6XotE/44Ep77W04Qu+BkaMSen6Pr7lrkwbUNr9hK44TbXusILQCPuaA
Aq6iWVpGWP00IVMry1ZuXeSyfSNgL8dcnm23RxBRMzB1mz2D1rXjQlDMOsV1
nioQgEB4xQmuZ7DIZciMXbrB7y09DKkpyEyH6hxKRrbjQj6zCMpVuFis5gaU
d3cOaRef4IAGVKdt80M3bw/9w7HEtVEcoMEtZ+8uLFtgrL2NXHmEmNtQ7f1z
kbxVl+Sn/anVDXFh22679YenJGwrCJH0kPL1siQaWkQbrJ6vpRxqAT8dREzM
RUlYDJ08usR0H+VFevhsAu5kuLRmlMGlWHV0cm5sCDfWC/ifaLC6CDKgNXog
25NZBvHWsPgF1vaSv200QxJN2kqVo6ekCeSxmgbJNjcc1c2zh1HA3cawaLhU
AxZUqu4DqkMor3cyVD4TYIGwzZdP/GKYhOzvrtNtLiFd8gf9pEO+qNB0bYUJ
LGRzQ9lfOZWhkry4X5/+tZQwgk84BVJY9dhlPltgWepkCcuBWxGe6OH92VDi
lnKue6piEWrc8XPblnJa0I10MXT/GR6s1IyUvnotZe9TM8IHVSvjX/MyPO6k
/u4K+PUZ5nCnXhSVd0qmMgGs0PZS+LR0eUmjIMUC4Bw+TxpNU4zuCyPKV+5E
nGczFMKossV1wKThW1zhSfB/3rfvkUjPilyWToIqwQroSjrfM78Ek8QF1I94
8A0C0gC8O49XJEF5Vbkcb0icWLAbAYOFEpNcJmfQLkkcr03+E3U8EfvqupFr
llXLZLShdPwRli8/PmasSEDOBGb1WcF+/BIIp4c10m4oU4PpyOjp2QRn0tmf
cIKlQXy/Uk/PjVxVmr/uMD3wjuCjlUt53/aEGR5DgTtj1EthRbQf1rBFxrhx
/XvCxoTpJ8ebkXZGeRGRbQNX5OjxzV3OdS6G/dRk5ZqqkuWETqJTcNVClXjH
kEx+tzyZyob5CjyL05kO/uJXIm+EsKhPrx8UtCgkt9QLnAXTVqv0wINTU1MR
WEd8L2FmReFQua/7Ny+jdJTmCpgLhqNHEZ9dWQ0D1w0QJ3MyGiP4ygpCQBQJ
1uwUIMXqIhQwGop3KRJH5aOSVuSpM5b2fB0WftVmAT5h7xY9Z8tHAm/EfoaL
cOj+yfCnON3LhdsZHIAIkiEghFAiUlXOFLvK9Iqa59gauRoKdPTQ6aQ914Pv
sR56Ks0799w/8os2sxkzCGiGJ7tjSuyMaWkCqXKGEpZL1jf0SEvTn7FpEws+
2wO36zcCMy3plAq7TNZo9h6rmO9xS2XFLM0Hz/e4wFLUB/wcMiWjkdT9T4GG
TNp2EpDzdziWJI82Rn0ouwpMqmuVLfphi4UH2SHtM3mvBG1+DPQVJ3N4w+Ck
nEGfk6ux76SXpBNkgnCERiyshF9HbIm/b3gy5HkG0QyoZ3S4Oh7EbFSMGkg2
3DANvPmJJZA8LPQm5scx10V96h2XkruhFAn4sAfVi7g7C43PHZGq8HlUOKUr
/IHqxaASuYPMJvs8Yj6NaR0IzBfOskdi2ygwVYSS9fVok2jPNYls7lTAeJpQ
8hpj9399r7Bj44I+dR4LS1M/OgLYJAuUI6iZ6nWfabRM4WogT8ak1SwVGMYd
FuCiImCdnS6/+nivTcdyekyVaUrXT7YQAc3d66lj5zq6ere0w4PEvYyhj5s6
h+IkRVxjUAYDqff+zymY2GUz9EjNM6R7fSb5GTwMOglhjgYQsN9u6tIR7ne8
+Ze88uCl/9BVwm62nQhECnFJYKc2hbNzjggO3oke15kkIPRszZhTKuPxbunT
GrlPYc02rsOi75EjOe8ORcegapijDFxWi1yZDoxCsJPuqjR/LysM02EvBoWs
wK+OPjlzLyFEYJ9xcw2bujm4bvXYm+0HX0QxjVr0gS1hGK0hCYxUQrj8yU39
qiw3BDkoi4Z/VRzlUGwiJNV56AU/oVdFpyH7oMRurvMMGFnKV1ODAmW46tAR
08uz9KMkE+rAKWKbBBGqTpyWLNz5nfw2ikTEiuatUsxZKNgJUPff2QpzTmLH
x0n+sviAO2cqOQrSx4ESWBQBdmbsYctRbiESv0WYIJzXe1+ZnShJwrBTxzwZ
KfpuqFPa9E0QUDItA8+B+P7wPukMm7KbZsXz93p6C0Hepp/ShlM23gvikjlT
AbNBoYTRZqbFrZgHGECaKoQRr7UJ6ba7gI1PVnLL0EsriQeyccub9uEHWJCk
qiDUqiIl+BxGtsfvSDuCAZA+ljHjAUO1oW+3YwTNqwYCZl4yKzT5BdPerOHF
bka1FjPp91HJ8rJwHHXeSu+wu8jKcfXvQj2inD5e/HcOBYG+gjUaYIcALGTe
HIf4fltpA4J7ehUK9qpUZd+YNSnoS72uClqoutKXmQ0JXTvOsV3BtWyjfZkz
xR2WP7A2g3sJVcOleII5yxoglB9Uz/HauAjc4fOX2OAI7Z6D0xRo1ti2lAq9
tNeRGlQ1CY4434iaEA20PAvEfUDntdCdehZYuHNw86DE9wNkOHY/KdEep+Le
bBhUvQBmNE7PboAIDipDqGrwVcrCEtXyxBQpyiP5LefFypu5b9W9sTHlaoU+
Hh2gP8NI5QIysooHpbhUFbV4O5OpQV9+zoOahL2HgFDgnouyg6uSYg40ziLM
bZtSchKaEMpDuGkHc1CR08EhhEB3rxUL5kpFEfnr2KUPi8CZMb9i/ok76hUC
tz/1pNj8IDrFpN06xM+tTohg4V8D4Oe2RpeI6oNJhck5iFk/CgToR/SeayQu
WUACdTqomfCwizTFnqWy6gUyrZ615kH6cimiJs599qkaLDVRMai23naRcLS5
LOI/mEeha30j4UO0CuNdcUNHxaol/OvBLZbI7wavz39KaaFXJmoEbaw1rLbS
AG2Y+hEreJVWgPMAbwUVbUlWc3MWDPlwgNtwQUyyBihhz9dmdI1spzEV7qPj
7BX9nkZaLlspEF5BepGU5ZcA5InXmzm2n57Tn9aTP9fOBxqz8piUmhHa84ns
pR9J50pFgbsHYIEDTlJunmI3IMpnT7iP80J3R9lyd+uY4GkTI2XsqcAPT9lZ
nc+14oVcwa9YnBheJuuV6cifefCPC/iu7v0dCS3+bI5ikTzmbuAuIGv2uRcL
I57RvLO9VCOwIdOPTMlyTpw3/p+A+ryVA/PbT2Wns4KXxqVMumhqRaboG4+a
YRcbXtjikTGY9f5IQwrLshu9FLwbvzBaHymttiJECtqpvt+BRnchXbjs/QDM
8ZRiMCHUMpWeUkVqRTUrwncF+gDRl72680rs1rrBn1FL+cse7uSug29UwhSk
QrDL9muU1IqYgc4MlbLTGM1Q+H1gSfwQwCKrSKafnASo3jBj0zwYfVfzmD4c
DtqL8Pb2mjOL5VaR68vUAVzGq66351r7OZFpjB0mP4beTY54fcj4DjddS1us
kJnxsejuLcF22dWEsKPMdyIfbNH7sDaBzrUwn2iR3n5MwJUMgQuHQBm3Sx9j
ltviMEk+BA7TosMHnzaTg9hI/zkuWymEe7PsT6SUW7kr4In0MnzHZpE1tbZY
JS/ZykttpftlErVpdGkSzr1JXBtQsQ5u5JtpkNZMSc4bkUh5kMTDdklgIewO
Cn6UHMauqq5z8+6WF8FnC5clI3uhAHEgF8GIOMNk1flyOuFeli01siJM2GNv
mhwCf0s8BvQFcuDtZuD/WfmfkQE8LPk3H9UaPAAe0I6/r54oxqqaQL0t4549
kTiF12V7lMggFQf3UcHR3F3cvB7TpsMtvlyXQCCdwGsznHsvcyGh5f+BlTdM
L8LGfG4frgCJllsq08snupuQin+3IPN3+ZCZn8rPj+MYhSgadJvWbp4X1za0
Cs+iNZlfvxowePc3yDbJJR6Bip1vMWXjw7GF8qM6qJd0qhrtd9S4/iMmnPsK
GmNc38XBxT8kK7IVDoEtT0YSGBXdT4uK/nOBu9fLKxgpjmb0cth5JjNbSZGS
yHX73tct1cEla6Oe9Sbn+uWtYunfHOiSTVQPEvvJpiwGXtctglccpcfXnrYc
UHThPkqh+4dsJn1wKeaEuMDDaktgQWVnQ5hOF2/KXYxlJ0ea6OT2EGFXZTN0
daxSoCgxS20eu83wa8ifleePmDA0NuJUTTcUODSXEZEBXEbKQ/3aVcUo9lSu
i9MWR9j/45LH+e5t78/dHxzcMmCZLFBM1Esdt94V+CdUO+BsiTqLjIkHfeGM
in0R08oOZyiEXxgk69EZgxy162J3eVqZl7MBze9gmfUxhHyn+MoyMephM8Gd
gzjIRkjgHSF55qk4iNrfyZeN2Kt5m11kTKx7RjzAkbnVd82IoWru4V3XZMii
+uvAK/MmFNzDOSjwHqAf5WBSxlqThosouqvdD1k5RqeRSS6NhtUEAZ6uB4Zj
a8dsMHCyPTBKWMyLok0sqIy4dGfpwOtKn7OvecHYjJ7JFIDasc6s26nfbGc3
M69Lh8DJUgy0CyXKTIQwQtRI+L6fIXxCldmOXDVyUpUOVkU6hKyTdgavOEvd
gUXIILFaz4I0S8AeQYERuXXw3q406XyfGHIQdYXKgABUQQ1XmucUrzK3tNz6
SbHPaOTHk+d8guJ8ujsaOiJ6nYPsRZdXMuqKLaSXbxrg4nhGTh2XDa70SefZ
xum6pc7lGlU0WHMA95m15VQIrul5Xe7O7Vtrdiu0YDel0bYhDOqof19ytK/n
fsHhD1gI6qSh0jton/t2SulMzX63aMtE8fAY16vSTO50QiqwAPC+u0bzWTEv
8+zIGqqD7lCx1VLlAowb16wU5yEr5llSHm5oTtPBR7WagcTQVV5EYjdyKdgt
EI5PWqf9Oo9zn0KAesqtN3b9YYX2ZSeWy34pBViwGTBuoHMn3mTK4IdnPHXr
m0ie3LhDo3ezzyK3DCqo3wQ39yD5ZDBCaQhKgNm3CS7p6lWYnXx2kA48x0EK
e2cAyF6SIdQq+zio1YwlYJMdRJnDktleIuok43FtfcmyYD0GYMeIg7tIAYeR
+ARAVbmVV0Tndc2ij1YCbIWjr+y7X89gpzVX7TlegMOEPGFCHn8+vYbiM6m8
KKXAhJP6H5+H11OsPACkb+/PlJU0mroG6RXjVA6IM2t1d6XFzRR/uRieEj0Y
oq5KTuRxLqBTMSqMnQIB9Dx0h+DhridLtK4wElhj+Uc6u7GgpDKoi7cHtrdN
T4H1g35pv5n4UfUNl+TQfd6YOwIGjeJZm9Ghz+3VAVQvvfCPI5TJwwdL0jSo
pCMXb0e7sOP0w9D3e4Z1hbgjCz7uuOo8JTOhqaibVDgOAvyW6QNlZAwRGDUY
le5Uti1vAFt+xdP8PETsyRWTTGKhOc+43UDlTJKYZvPUmxxOs8pIBRAyKwIz
7kkz7YplY62oF3KZup1rajVMHPU3XPIwmZBiq7xj2yuoal82WaqMstVR6Yv7
cDPN+fdya+zo5dMYxE6HykMOeSwhTx/JAoniUCzN0NEtnYY0zERCmJj2nFH8
PY+t4psni8Tjg7+PZywsO6Eo4qjRicQ3MoL1hyHHStzIVWno0uy/QYrdE41p
ECOqINruNOqNlJskQm9b7WY/apqszhWZ84vzrMWHPneJgoYaKv0RC5SHUExi
m2Joy+vd0MoqJCZePUJuV3F6k9Y1RUZjkl18jsGrFNeuiw34GhzlAxX15kCb
AM3DNTonXBiBcCmG1qk9bWvZrjOm2tTMVjM+yij3nASESbh57pt/9GIUpobD
C7AaYRLunaXbAB+5m/fRykvO8DFy4iMs23IdBXnubl3VEaBN1tZ5vG1vkXnx
HdGSkN1PJMkr48qP7P8PL3nKP1c5VZ0VvvUTJlQz8Ip5KKzXgiW3qRz521QS
FKGuprQNuWHZts7T3vOEfvRI12KhSiTMO9bpWZ81syrZUolUXjPVHY4eJwmt
LaojsCpOrMyrCHHYVjtyfayq7vuNq0SRCK1YPeJZryD6jfVekZr82HyiurGm
0M34XBTT998+GMhGCaj1mqNLT5w23dcSM80JPEcS0TZX1qvKeSaB7pJ67mmv
oWikQQpUpI8lKPusHTF5A5Zb7o/pb+1vREamC0nFekjBO1dxwN4Ew7Uok64p
ptwWJYPAXRh9UW/0wtOSiJnPwzb4iDVP3yq9vwk5rlT1W4TFCXYt13yTiXAN
aCz+UoKANFCKUbKJEV6AM3b/8OlEs0qhqdpg2TnOqmOxNsl0VOdFgJYYGagm
qRc38lJteftr8FYc5bILv9QxA5v5WvjPo5p5rseAgbeyvU0KMtx9ueurQ5c1
uNxhqPP9eHtdCQjsMI1EBX/58Ixx/L7B44AvJoawaXi53cfxhdRlpZZlvjbp
rPmUIP2fRlzO3if5wlAxxqHGwV000mCFcNszvMj5OmzluERJxTj3w7VYboKR
HER1X+fpjwubybAmhe1TJB5fIN8i3Y4F1b8wFIc/ol52usCWUERc5sbNjFGO
vBIlqlwRMWospfkGLvn9v7jrmgR+N/fu2ChZQHmcVOc2rznj+MbZRG5i2Xye
9sBsbAu+YzuTX0iNQq7wAv6+OKWuWEI841DbuUz3ysBou4PArjOX7LbzNr7G
9AVmLizGhSC+Ns1T2v+JTMnKRs4A8IMC9tWJP1jyxqtAhdurUAoZq4oFbZTR
wYQ2KymbUu2cKTKcoTaPlAzdHsUrzV04vWiitTjNh1RdT0x2K2q39K0TIxPJ
0sLdQLxEguLx9D33iBTLWE11ijhCZMaoUU/zmlp63Ct5OuofhJ0cUhpIEEq9
sCT1fC4PZyfs8LRUbBE20I7+1C9v3VExMHBKFjgEzfH9sFj8lDEJwqhrSuBa
7DjS+pbfof6mgXS4WaoH4Y4RNkJYj31ZsmkLqcpqdMN5grBb2dxci1f2pfIt
d4PweNMUCORpAWyo9jBGbxnS3AGdFsKg1vAOzy78CZexOm52FKqUAKHdf0fG
uLlYY2DP+qepf56O8uLhJD3/OQRdx6p+He2hO1MxiC98hv8UYVZ20/HWCoq5
zMoIseW9Y3qpGrWQb5PH7QVWCcd28kjHyNbnCAGfAc08qibzYi3zV3YaAKLz
sSCDWg2zVuwiJ1BjlTN3bHY/k+J8pF/WYnWaa4/1GPkxpVvIe7ptQR3+TCOh
weP/KdWPivEqv8tlY3gy9nbbwe2ljrQkblnzfpegjhaLCANCT1wwz7XVxCJS
UYCtAeC6z4c3Qo76v1acr9n3GTcVLME6zI3PYx5bp5CgF/+sdm79QsQBk1OX
GLMEh1L5kJ3JR+DOQ5BwhwBfzqVdRGj3VhG5teYjEGDrnfqCUpnt4KeEVMfl
59099/qcmabUU1Kgf61GdMjlX9U0Mcpf1kC9w3m01rihZZskLWrF7uLTMjSC
dz791KQAA95FfyfLrmR8bb/qXnBg1zZZh+KsPOKe45DqJNuVEjhpWpyCk9R8
7y1TsaqoQHYGmImcsf9GLmxwx3gLEsmYO2rtevvUN1laaOPL4nYCE+nIUEjh
+yF/jpxG4NiK3693uuCoGXzAUFa8hmS+l70WnVJF23TDgEtYvfhzasmmg0DR
XvQ1tncIbN0o/+bL+vUVghVAX67f3Diw1Hsj8TmHPrl2AsE68kaCjbHkkNV6
bAsCs9I78KeeKZ4Ts2IYnXfI9QAnmHCjWYUw+v4+2pVuNxXVXDjCYBcg0OoL
hOgmvsvmiBKm/iaW+TkQa6yKlBBGrJrHJXoihPttr2nSLZDMyuKM4WWJn45q
NU1zqXvHVnTPDSR1lciPv92RMWy1bv9Aa8n8Y0MOIcCM2Q2jIYXnTSf+QGnI
8u6oQsGD/hsGmuqDleh2OechUjA56p+FKz/Kv6mzeKUlvJYqJomKZYFnSA36
y941EH24Mrg5lqTYaeBrI3/0mUGgH/Amvvqs331SWTfv0Nj9+NcpqCQlSuSw
HvAKU/Mv6QczWhDwlEhSVAfLk8hK4D9vfwKnMjtoyPcnHHDP5EAm0mjaHQhV
9s8oSs5TJYDpVewiT9bSIgjU6iniqPWaMEre1vCls6fJ3Za3Ff2ABtz8M/To
uwfbFja5+hbbx3X42v8Eedy+q8G1IHnjpxAttoAGb1lvQM+ucGzdY4FpTU5o
l3PNhI70D8veaZ1u9tuk/KOms2KSQp+4DA2h7IhBzH1LAwymOfz1mU54+evC
LGsElgaCp+LRwDomjiLM+//TV3JACkn9bs6+aZwJJ8BuubXxi4DpOpJ+ygyc
f8Xq1nA6X4NMHOx8YXkNDuK+EIlzz7Bp8nrzWtOkKkSTArq2UGCVDlsSFB6q
PedKy2PQKcylxFfXbpSDMw69EsHP28Dsi3RnZeo66POjr+MbG1LbnVTRS1uo
I/Ob2KdtlVRa5ABJVz6UJD7nf3ZoYJUlg7KRYoNpTLZltTCgaWEy15+cx+px
jZBkE53FI/7P6kMOXDSfokhklLPJUeh8BbtZ5m4d7QYe86/0JOhVMfQLs54s
+TnzFQDEe3hBNPUqw49xBaHrGyykqlS8gWypEA7EPxj2DOdQGp0LM+DN2yu0
huPeIiyoZf5SzOi9GmrsiQ3X4w6KipRjahcztvNbpimo6lTaM4DpkUswNeNr
uhmCUdE3Qk1BUhKAXCVWS7Vg1k3cUOE85+mWji9UYp6z7Ubf41fJCEOtIQ/K
MtwL7CxqVkhDvKavOYVe711v5q0uIbLAYZeQ/Anz21r5Sz8kQB3QngAOO31Y
dXoyFudgKTL1wpPRytGGHpEvFx+T89i9+qLlDxUZNRf2KoU+ECxdARpgfAvX
+JCwVReBEyWc3EkXhS/IFg32pTmyU0BzG8RiQdV9moyLbvvbBk3GR1uT/0VT
VOgTx4on0GlgEZPmbgoQKdld+r0DpL7J2FkZEFvQ/U4sWHJJE+HZP4Sj1tF7
I3+gdIvhBUIRR0aJa2TZaP8+loYgbb13qFyEmR/YBzy/SDsIxLyz6rSVAeDc
eRjBdqJ/aCrBVm7IZsyefPkCgzvSZRBzE87MAmVpAzSekgv0AmtfFts9ab1v
4eYebbs/XluFD2Xn8vDukeiM6dFFNsuTu6pu4bcmd9FvjLlHTvo9zfNCno/P
3jX9c1tf4kesa278IRWqVTC/j4Hc2ZU3JrFeXDcQkgrZg4krlFH6E2NJmlwj
DbG4o8WQGFvUATy4h8LA8FVR3ZC1T1NGCo2DVcC2y1w4I7gAa+RYi72pmaFK
uxQIO6PNNaEMWTtgGbylTwJww7uGx8Iu4jty10Nhvw5U2L1DY1KOjLHr4x2A
ppDEkdH7GHH8UnrX6Jvth/pF+5ekCweKtIBLtBUKRqL53vaTIzZEuefr515i
wOGqT8rLzvbu9CrDBXy69bNNg7nrjloT35l81Q/hjttNDdr+tw0D756lAkx4
cmT2260VUdCsvrLMgaN4DExIoTz2eAZdke7f1VkwJ4U4fZ/23iyUwGQYHEMN
/iDPKrv9ornV1SmTDUrMT7HO+ON8vIBKy4W5yIEnq2t6AxABK6+mKNnouXzv
Jan7v9Txeq5H20VYjnTj84SO+xFcG+dwQ0o64mjq7y8zWzVSGcUIEB1+S2jl
25JzriTfZ6/iojhr79S0gCAoxBVizb8H4Q+zm1wL/rl3SAa9UVJur9jCZgTj
OrkRWsEJfQ841AfrWEP/Z7MsMEAaedQYBApVYUo4595e5uhUimIMBIXTRcUW
3dmntMUnTjH4UfvaL/9EZBf0oWs8W9OFmKjh7HasWubyNV6WiL3a2BFTeXL8
rx+QwXTcWURu/5zmLMRUfSb5aE5CJazP0XiU8YJ5tHZdXOC0QgoXaOWzpxJn
jn8moUsoU4FWeKOfdrmp93Sz+ax61TbSQV5hShju8AB4ViyZR9RLlaRQI8uD
OuA+ODAiSWZP2gbcjsMRwMSfKrYQsHvCP8FT24rmwLI0cJ032NLfe+/xp0H8
ONgC/oNMAHki5Ov7UI51YtIdvf1E+EUg9l1TJgUIB+eoyl5FoMF70YmQPWgm
lhUgfQ99BchfIwuSFYwcC2v0ZmnAXxEcG1bJb4kwsd78j182By4jWu861olo
aBIymgCkt8fzA/jGv0twMCmzCjqxMw2NM1fa9FJ3N0fW3M5hRaV1BlwIHXsJ
4fBKnAVa8ocDlAPFSMlm6nirNkt0nwheFb4rFEkbQCXaHBQ6d+gAu4G2E41J
O90TXV/LwXAJxJpy4TpQg3PcC8/a3N3PJw/GuM3lQmDjUQY+wuvH3MZN0tV1
xI/835SZWiGRlnjwi/820KDBrlEZR+qC+NJWVY5FB7w18CYwv3Kz9JzZ+mWo
ADK+BRLn3Gw3XSUdwvmRdPolX7fBJ0sZ55zhU7w9krpgKt6ELpw1RtFWcD1o
DXQDpphpxetyE6k6/YAPb4GRMb/RUeZYL3NdMaxGFwBLBN+2w0H/Q1lCCVI9
HUevEafxNyNKJJNAt5eDKNs8IjedAzHGaY4Ul5JKYZKwkEY12+54gW/pTHM/
mT9yIgOWfvXCmj8JnX88aivYQgcUwgzudlTFkoCPJxPyi4cyw43KamrhRmyp
gpPzNoerGII+zFhFvZgEP6fH3qMxKVOLHRrFS9NMzrxM8iBNkKPcWavmJXHc
cp1sX8SbWsIHKJcfNKpiOvmSVNWm+5NzwzYo4mqiAOOt22Z/waW5ftXnTLKf
lBmUf4UZy+fIAMlRXwe8gew5y47BQxtG6F7pWh9BOQEV8TnlLA1GLq1azu75
lag9SIK/YIFZLSoou9/5qR9sGkIXcf+r2ElAB8WTqWUGXKs97BwPpLv9sGLz
9LA6C2RgJyyM1VDf4Nrff+jh0q5to/ar4z4GgcLUekM2QUPFT23um3/HgLaI
ZtUuLvZP3tawHR87pc77DavQ4vuGsXh5hJnWSZg7hbf2lAI5XYd79RAoKiRo
HMNlgPJ+0Hw7HrsP4S4WEDywJlqqPnBlGnXOXestz1TkV2O7AAOA6W7xXrhj
bnGB6MGLD2x9j+eY+tXhpe+k1LrQ/L1au9XBT9b02LYCr/51cy5vgaDWe1qz
+GClGnH/xT2YJZ4GMAo8NDVFL7stfEng41UEklFb2e4pTy7stvmUrUPo/E48
4GK6CysKGygKSS+Tj1UxQhAUwhgdaen/+GqcnrcB0nYAMwgM18P+fO+ixAkZ
Bz+6E6y1l+1/0/TfgReNChvDE2Fue+cyB2Fz3uQbcSbdBykDWwuz1wIuAi/t
8+JpLHomCmWFICNicWpLfCOn8NzU9dlAuEh0OvtOp3YbS/d2/KW2ed3dQMaB
3KkV2yzTJBeYJnYKUO+pKO98nAXThIT4c/olwvRC6GpxE2Rf9S16lONd//wZ
abJ5VDUPLAIDEt4Xrtqc2+oSCDKIfjRd4rF0iEui4mdhQrX2b3XOrOyu1EoR
DynY59tUT3smUpSfGM1RDIYtXv7VEwUQlEY0og13lix43XPHjQpscBZh4gjS
zQ1A464VRoY5BHq9fZwky/wdi6H0AvLmQlpvRzQNVz0HiquIOwsrqxBXp+D1
Ux+uNM7oBcJzo+OdpQZanQpXkpqmF7Q4pt6eAAz7QZ6deWjkScf/x1pM87Ja
h0VURXfcOevp9uyY/V+BTP3Dfrza00Zr2tU9Lr4sUHLh7WWbKBSfQWhaOPq5
YEX3SmWxzal7beeLLmDrtxJjQ4RtLlCkKhu2lK8OPfWtI35FfC96b8kJ5Emy
xr8SPmuQdkjm6ug4I3dUmHtlC+RxURG9v4/YEr6rtSJiR9JTk3erjF40CeVp
dD89pQZrKv2HBok2BdKvU6Fjh0c2ka/rNN/iUwPZhwS4TQvlZBlj7L9zY/X8
pnwsV2qzsUKxpaHC0+l7L9Xl3DoBsf8PVcDvKprVd+yl3z2SHXNUJUeWKAZk
pjBCdHfrUJ3Uqc+lFQI85EKQX2R1lK5aNmNedBKckjAI9VmW0Sf6BivOefHR
N9q8cAA0YwpqodKB2z+DC1676uDM3a1aH9ImIMk+VS/e07G4XQ6ixl2Qev6l
vuYwnu4LEVBArMcQpnuwMBOiOsEhoTIcr1eBGFCYAuBH2atkQIoxj/owFyVC
Taf/lI545s3JoFB+uOOmakveOVn779o+4mwAJtIHAGqU8uGJ6QY6AqbrGe/s
2G1Apg7nR/d8v27OMaDIrRl5r/jccpdbLncROii/M1Sw3ImMIb100+Sn23J6
g8x0ukFv5QmpINhpBw9lQKfUAy9kmTkQkR3pMD9Iy2JAl0u19yDaqMUZ3OFH
7YMsON7Tnx+6hxHh41P2YlLZJ6DCCR5EZx7qJcbYqvGjZ1PUZI3U7JemqRlB
qo+7Y7XH3njYU1PUUnJUo947+zk657NUOPM1C56JCtJB8uLW5zwEwJLQMw4W
wVXG+aMJufMGxxh5jN1u4yVbMazVdfrgpSZzTq0QiBzwF7Q+gFmDt6WiDxUp
O72J2fcySX+zlBeooKHJoRUaXEMNtXIMtLfDXGZ6QK8XivYm+W2QOLYDUy8+
2JdqV9yk0vCmggW/RjAk2lveSQZ3VVztvzvoUlJ6rBZENWlVNDFXlQX6GpBr
xo8c9Tj6KFNV4jIK2BgIuCvcuC8hM+13viD8/SRqzmHOYlYr0UFtood/HNC0
As10Pi44X/7smlEqz9kMw7DCN39aEgV/TFipDYA35bt9fyL0NnRPd2Gr7n/x
MQfTdrH828FaqlXT1BW+lq5GAIT9vlOwh8DXslMfYiIBtzkRtRQfGq7ChUIw
HDWDc6s/KquHMemQRkN62c4lx6CPd1epj0huwJavM0VMC4eME4n1KiGGo7w6
OTWLleYbDDw0ctsIr2sLLJhdP5nvXcb1z/XEJFfubUB0P/4W0PiekWnrz4J9
UKLEur532DcIaw8Ig3uDFWBI4+dp8aZy7092Wntyv5ZT3KgYLRKAK/xH2Y2L
H0MFTzqlRnMwCiL4cuSANW9bUCQxCx0bRT/Uz6BKybFZRMeRVpX9R593bYOp
iWli1x+RzQVqCslFGbq5HlIIhOtuCh3yrF1X9euZcocceooyre3aFlSRfnIh
rXfBHMGib6VhfdzBECf88YhUCxDOsMsVTNea62IuNapv+YxekjjROQkOXDxh
dyqrK7QBYkOziBFsVqfatfmT3/m7PGtjliV5qBeTRt9owguWNiJTpBXkFALL
1EhtiymIlZiPEBxKXWFA3tguvipvNagwrMvhJzi6qENQM93jcKCbkEwXNXcP
DrnFFhSd2aEMFLK0TSoe9sA8zVXzxd3skvvVdP0swP1G/q1F/N2QV6KA/0ny
ZE1x8QtKLGxlLVa0Y8uKayRGq/fZm5MGMlhVihJM592l7NRn9GcDMBj10zFg
wwkqKr0R+cm91zcEqF6GsyX1UQ/c+YnKzhaRkK1jVKIND2rV/5Zd5jwe0YVz
wfUCwQnBws8pLipDwoDqfzQvakPdNiwN6ds1DNzDp42PhSYPkt2AaGv1Vbwn
RnDYa7yT3l/xaLOV2Sh9Egt1Sj8s+/DbtP1lJQwyziE+BXCGc/aIyNKxx4cp
Wy5/ejl38mwzgg5LRAVvNfEFbyGWb+HgL2oIL8N97WPKSLM16XaBWdjXcmAf
GXG2k2hwi0tX7PVjM4M4ZkwutVe9tYWaQ9NZbCn4WFA1nFH2zu0esfquKa9p
0pk9UDiZSq1iN8MaguKkR/Bhc2wYUNUmHGls34jCZ+mM+Y/F/XQCQU9/knQb
vz/beJoxx4gpH5bGcrjf73e+cHNt6g+Z0fmZjZcTFi7AdhMc9hGB+E6xZpSC
FynveLFXke5jiyYN0h8vzlKv+fdb6cHtai8tkt5kUK/RCYrKY+zDbXsKD5Io
x7Wir4ge4eBlFE5RcbRy1pSfuuhx3cAINjD8jZXODCv2DWjyBlho3Sp0GORo
xNAghwGqK5xp253bfo3guBoUmSYJgqzoMaGC/aeaw8uh0WcYj+2VSeZmaScz
mZ3oXoLQQeHl1P1KjXJ/fhsMdeeGqrPAODuUi7h1dX6Knio7rqNKQPk8G1Wm
UR2VEGzTLSnJe+4ZoiToCeuK7z2dSdPZJJBPCJO5LGCZYfxbm51FSEQvki3e
iKrxSP5R9ZwlDzOHxQT+v/CZlVKkpbokzOfO39jjuvmxiaab63L8NLbHiIs2
PlWbv4PpsQsIVwUNGohfYWvAaV0xGmr69Vxdgkx3lO/SGBXhZqYkTkOwm4hG
1JlDz5t4/D/sBRzeXgiV4njrR7vO5FHPUCPvghiL4dSLoSc592ny1QfeJC3R
ew3omiNyAUwsKm9fSakmVQRG7pbihMQpeCoqxMvH6dDxzJovPJAbkpLHhf0g
6X7tKErXmFutgc16CjhR43kjoxkes60yWA/zo/EPNvWyd70wkvixElMVSmAT
TRdYTLuxlYSYrdFilYCrvLS86gvtr2mZuk7m+1pSXAfcOJ5PkQrsJ3eP61H6
Gg3ma7KfKwouPoXCjjIez+u9jUY60EBPWQboZZigmgJ7yRrYk7Yl7jUq/Iry
zFeJvWc0dxeZA/SKOIPt740xP9ntGVt/aWO0vPxqiowLAW1Te1qa7JBbCawo
CbntsgANevfnstW1IckUuGcFYVx9bpbTUSk98sUfRVZYO1a2e6to+fIuRKNJ
4P4C4fvypoFToKMdC/FYEDE47OCf4h8T+DQJ5JmLxMLFIvN4+RgNLJx7t8FB
ggXTAnHl2U8LECtw0Pzfw8PHs0/ooRL7l83co5a2OUXq5uqciJ8l78SmgN+q
X5jdlKxoJIl8Knz5DWPQxOv2BXmGpCL/SDL+6DMv/PlMly0asPzUjXM2GkXT
nC6izc9CjAdvaYWgeplDbA5XkUd+sicTOim2vJzuJIirq7Vxli1j51JPsJO8
2VoHrsb23C+OeRG3dgKHKTIbnNOOpcsvMsq1taffGyUk0xVFweesRzpxWuGh
UWcpwZJxgx+ol6d5E8Tj/xiVXueII9/yDofESbEZoTXcblhYj2cCx7kZNpGt
xx7xz2RN80xNzR7PTd5EnN23zbYaULL2Mpkcsrjq1lQ/wacKiM10yFO80DnA
Qe6wm09wgThtwkU4oTYTgIYWng5AWPJUqODo7GOsYby2gN0707vHBr+BKc0B
FM1os8kvPc6/qz8JEzSlHhCwT67RTY8+x/NvQ9ARTrhwPtvcKJZRxAE0T81l
JC6w/kYRzMiN8FYNwwxbumb1e/a62bhXc9NinoRPQd0loqi2y8dzr5anSDce
WUPiTHeZv5xgdWRLonBLOTEPEmUy/EhdCHF0Ya6n6E8e6UMric/mCjS41R4/
DlLoc7XXx1f3tfyAIkwjTIt1wiwfbkjPd1MoGdFFH61vWyRbdmdb2X8WfkcG
T1z0dop/cGl2G9SjrF74hLYVtT4yhnb/6N2X1IR+PfLDUGztRn/KS/kNwSoQ
1dOrDGUEIfAONVMHrKZU2mqEbg2hUJ50R1RaGArCz10Hb0v3m48JXFCyeMGk
VCm+CTRrZYLK3bi6iblAX4agXu5qdaWTe1zjMfRuU93dvr+vyjl6TSNPbHrS
kvW6QoTJWv2rz1u2vVmuE2Ip8i2e5WvPfdYbJpWgk/Ak1EQCZQQV7P3YhkU3
Hl1rCLYbCfcChHD0FTvFHa9tnDob3usJ/ugwyFYLASVpJm3+iMfXvL0s2KCW
asubYaUgxmykkdDPhOLJDRIq2vsKYQfQHgs1ijw54zUyx/KeNqFzG5jfJ/p0
VmNUAmOkqzUSjKgjCG/DI34gFXLvPWgPHpx8lxv/ZGiTIqpi2uVkW+hS1M9T
+LXBFVb6OpaFqqyXT9M77mpSZaYbwjXdTReHkziUCk2R2RtAntGDYZj8/407
b//94dhHXHzn6vOfAOxGrSAMI8HiyGI6xkL3VXKZZcn1Nu4SduR8NtsuyZS9
jL6GNqszdX6I2WwNNCKzHIwpVY8YEuHPDg+YrNYy6UzfooovokTH03XXGhx9
03CeaYpb+rqSiTUrC2KPAoMp+WsQiffQF1oDP8MsjehQ4M1GVSg/FNIOWFnP
l+6L2LWasHzptsB4bYMp0Rb9rivNUZrHJXaJlo/ctGpFDvyRvm1UHZGsvPbV
lNbGXtiba/mcx32AC7V9uEmeG9OvwD4UFv8jZEsmphS800JHgUPxB9B5fSKJ
FSQOUeA1jHb7VPA1ddw7c//DIpdG2t7B34yIGUNmjWtBatDcl4WjjPH2LEAP
Qn0sM7HmhQtsHbRj7A9kjpBMHGuHjCVIOTJ5PD6o1yKphErLFGGx/OOGFWcx
tnaYjeUrYGMVIkD7oGCnq6sr8L+I0ax0bHVge6Exz8DBhprFr9PWnercPVCx
e5ypuB8YgOL430OksEh5b3cH7eXSXKIFQfOVdlF5iNFXzTEjZQe2HVU1NexS
G5ziI67V4OzpEQ3KKr7pJqi7mQ61AYXr8U9jXccs0Gyu13V53tpaQFExcR+N
xeMm3TaJEGej5B07R20OsxR65rGMEbfG3MGy4YVmwdz4adM+MPChPIM7BYvf
wgCLwTBGY33CmlMkf3dxYKWSVxt2Dl23b6dQYZnnfwCAFkgeuoYZNWf/VpC2
zIW4MTeyTpQCRmrfQBw5pwAkIF+Vma44Xbl0TJYhLPO+oHMVfL47fq/V0/p/
QWTxJFUXkhEzyVGyfo9ts+uEPNuQK58kwake0EatMwby+0hEDNHWa95GUN+8
lRv7MjX7d6yA0Aio7Tco+zybjjqco2rqWiZV/pcjXbI1Evwa+brwCxiX3MTH
9LQ3VhXWz2JlhQy+6yHbFsx/sSbuFxFpIaJZAlghikNRnW2PKseVZbQ90jxU
T58wDhmHcBlfPFjEo+Wt8k9qYn9VU0hg4ZtbNisPxVH50OL3sKKa/KUN5o5m
qiHUwb7MvB/c4nmK6rU9oarEQDFS4Lv2kPZcYX50tf77l6npLnwagWDfECGq
fWXQ2/kYPVRGlVQdV5WRQfjG5W8E6vIoNSiKvlhaSnU9b23k0xpKmrhh8WFr
nk5wBv99Jz/WfpAeudO+8QT6qNIrecTfWU0+LFMV79e15ViGIT3PFwXkHfaH
9N0vV4BTftKTOwFwd1/ATjajj+ZmVGuB2QQPvCXCxKjOv8C/D0WPrZBntYH0
J9jTVd4yAktYqO96Ad2zYZiDXijo1//NRM668ILPTFcRBQ9Rm0U0+VFjVDCN
cotdl0v6eA5rS/H7NYTLQqwfFod9snQq+PMIeftddG6ywEsCyHLpjtw7fNIY
mi8NmH3TBrmlJMkK5utsc6xDVVjAfL/gOg8m47DqA3/NCcDpupYI8LgzxM+E
5zogi40dlSeCxWcImWLKShzyP3Fa/RlVgwehJX2w1+OcT0rNISazNJVqI9/2
LDQcRcoYe77OgvD8MdkkPFB1WXFYqpMQm0S2FesHk61msTlErpQ96FUKjgPa
NImoYPJCGEsHt2Mgz4/LCg2PEU11W3IcL4sDrWtzphYl4jl5hlzaGm/rDvxJ
IHAqgdO2WEfYXsFxAFRV8iPjimHLogNnB3/xADTREdqhZXO56cxI72lt1g3+
ZL+kliQv8N/n0F5BRttUut74tR0lMo42ucSs8ZeXajoXiWSwR6UC2MGoOTTN
pAovNWTnqT48HPBPRlem5URZTxoe3U4Gz2vhf51X8HH9H/vb05gkyyU4hP9f
T1/PFa2WUDCQguX944KvvzIrOGuhGyxYfy+qCKLsSAb85FYDVa/FJDWC/x8f
CHwC8Abxe+de4KZSed/d+rxcWLlrALEwicp5PDMvgtpzKAdwX/BOMlt5wNUn
NjqW9svVAH491QPkiyOAjnXzYY2h9HBhS++yt6zGLKMn7gwcXU3R8tq0iOpj
T1QsabuOhzwQp2O0TUy15EJawg6yQ0y558q/q/V24Cm4MJ2tEqfwrfUAl14v
b2qaYuVLLFlM7bVKfX+oALqAUvrwDRSoKF+2vUb0ubapCX/lvFLuXnyq9Qze
cQlmzQKpH33Fk918/R9FBf2siF+64vHBZLVtj466Fnmms2HKtpGHeitUJZMO
qSvEN4ejbOPCweyj4nxa+RGHXV6MPDgeMo30wSx4/3iFN3oj9i1Hu3ccmeK2
9xVxXVd6UJoiVnIQct/FF8fU4hQIxjNfEOM9ifRMH8+Qy1aBxMLe6wmvEYWG
Wgu/0dy5cDUP1o8kf1LeHzy0S/7h9ZrYU0WiR0El9xEyviaEjpCDh5O2pHlA
eXeL8GZ32jXQRbc+c5N/dT80F8nxSIb9iuI62QzxSeKbUKuKGyCg1H05pGpa
VJi9l7Ho3crG5hf5T6qNdhlEnPZFaunu1RoAvV153arzHdhDswIkX9XQWRKv
uV+mZZ2k+nuuZEzvHI0avTmYydffo6QDl1qa8DA30q/4SU6zsEthqPiPOd2K
bBGhyZ9oJ3oJYppp80MBjDW6KF3LI4qeJalMmHN6QTjLbm5lPBXg21WFUaDs
aPMuDBL5G+qBb1lSIzAMPK19IYc6qOqtiWiSive71bsi0OJ3TQKuW5HsT+Od
AgyoR24P3j7fo0U9XDfDiNKru/c9N/D5LSBQ2qTmIRt2Ujv4hw+JZ8QFn6ZZ
qLeuI9D1W4w/mCCDE3ZpB4hIrAzdywPg6Z4UqJrSVHaferZ+DgedXaoTVYyq
964NXC+rMps58jbhlyn++wUrMk7tDHJ3KozFO42rMhb5DQuRrp2AD3vF85/x
VIU2oIk34rzTzd2nhxKwi7HSvMaoGTnmNX26INgRbAXHHKFqspxHLbRvvfaZ
V8zkKdu2G7DdduXIoz0Q0pAHGZOZfL3k1HroOo6M4jomTqvXFXfAOGsXQYeM
7nawUFdTLbpBtUiDOAKh0dw+N8dHu6JUoMAf8yroCQnY+wVK+H4S1pg5o5d/
gzpBAq2+oM4EeM7Duy9hq+eyK7xcPR224aXbmFs2Q1IEeMRVKa6rK5mG6cAK
bfiaeu2vAXpv0DFqKwGBlGCw9SfQD9bV3zogXNNBIIaw17I4gRuDWinkP354
F7wdGh7S/cA6s2MqbiEF83yKSrzoHtQ6hDqrMNk4m7Z1gOYnWEBLDFTcwyKK
YjzeD6kBqGxgvfw7YsPgp87jUsJGJQoTZQtCK1bWXaMb4WavOqwPxtnyT0+c
sfUHU5FAAVb3Gooh9rL9/Kxlk9ZteSqZ8qFHvG6ZnYYUxwwVOy62eOu5pEmS
l8nvPb9aAMFuGfH59HImUxxB2Im816R83VpOniXY/zBf472eKAskCCXa8f1j
Bxz+S3mI482D8OqDTIH6aBDkGZBaGnJk3vSBpqVe1xSC8spVOaO86a8hLTAm
UD2LFvx2WpWX0Eovf4dgaQOYM0UHGQvFWMVfPDuYY9SjBQ51gSWtc4kmQU7M
/MfBzKlt6QKleBPJPdJ2b4AkVrgn2+2hhRkIIH+FQRRklNCLBhs+Qhs4aHO7
MdiqLJUYPDyWnh4N+s1G4lEtoGBm8h8iprsShkJbc0hUlZ9cKLe2yAlUGRdW
uq2tZpQsyHZzEYg8vxA7iVUSk1A4tt5KS0sTruJC9/9szaj63X74XyVh6q5f
2+l+8fa71e2bG12LgGagAkc8H030z+RlVYvpOcEzaZIZE6iO5yOJAje8QmmW
wPFmXoagHNKpH0LQyaQfh1rlEBHkl8d20+RoCsbQOxSNsIyfJX1Mns2fSAUx
dqCPG6wLT6uH0VxcpiZs3OLDLx7/h4T3x+9hYXGzvxwXsL3bDSvZbWj6dx2T
ToUKrTQWF/Q7OoBF5uLMTabWsF/a2hLJcP6jeSmkPDY5atMD39cdPEb7Az22
/DK6XuAx4ntyzGuihXebVopo+mKTKL9re+yMcJegdD6sUd9opZ6LXa38saJU
NIj8wjTkw+wOeLcxIEc8ZJhShpnbQ0wIT596nn986SYrjXQYB5QOoXxeM+Dd
qcwaRdmpFgjwv6dCwfAhH8/Chqquq8ADkiYjlWA5KYZ2MWTIrhmfNvS6pkGm
yMkk7uKujwQq5geuZqZgxk2RTBuiN6mpDyEEN9YhmqpYh4RrT5rGHDsN3Ro0
8BRHqkBDu9CL3TYsncqasHF/ntQSY0kKjlOPYz8pntZ9pOj182ZuljPJutFb
r3FfunaeAtdLHUeTkWBMGby4IEVQPMpbeZ/4g2yTNN0uZIH/BaGlXrh3lP1M
V4kEB7TkIukim7GMwYeWAN3m8WosBm4NQ53WbQZBm9DHjpUn+1pXw+ZEN5za
xRp/q7b1V+CnR2xVabAf2OlySrpCwoUZEACjRP+3OzdSyf6yJKUleJKbJehs
5L0zf+MtqHfzj8NaZoXEgaic7O/uoCTkS4YSScKoNSM3dqgr2tzOPZsMnvWj
CqfNpqwYSMvZ8Df92g6X40w+x/zPsZdCjze2VhC6Gclm8ngAJP+rSkAC/O9z
oRsj207LpRNA4pEU1ekdN+Fbl05NSoJr6Vyj8gDm8DPo2rInbnyTi35DRMyj
DraKK7UiJ7TmHPnqodtawNnhzfFfl/P68Z/iMpiAgJh+xKbN5IWHiyew45T8
0Hgg+LQViG3h8JXM/WxvrZM2WmAwe+NtSd4EEPIxh70gfUrkkDqDXJ7BQTn1
AnkhYFRjgOtT7VGeugRNpt3Ygn91pWuawhyHJqUMdK2F8ThzylSb77jGatvX
mEGBPIAIjXtmtCLFB9XvWQexds5IfiwSftA6UXnUjL/aFoFhfM4hkGtB/AFw
cBCrq9750Z0MbPQDB1S5rklGjHgqCFJkWZI4Q+62CnzhE3MO+SJVpsnCHKg5
fLxcip93In0VRzNLeyZybqCyXZnu4066Dbk4CaPSDzdr0svbp5z78NfEJ5QN
UALTmF1YEvmkOt+8xcrfkYWqdtG1XIqgJ0gBzPPlBPIj4YqbrquBJKB4k2s5
EeDK3tsqtg/jfuDSDRFl12H45mxRLuBQoXapQWIdT+QnSoDXvXANwXNHHfnN
CgXjLigiLbvAMo5x+umj8LazjUKDvsMQYPSaC3ndHhEu25p8MPNGlxp7CAML
CGcc2CFyiL0E1iUGMeNPFSBwmZJBtLDn2Bi/wrYkQ+006jR4Ab0FAXKUi8YY
T0aMsClOwhDTQdu3B37TLsA+336YbJI7bUsO+yn8Bn2YliG70scwYdneH3tJ
e/nMoGDYFqj8eTffLQNSwkYccuzXlgccIMr4tLi6abmYFiqaBYxS4/g+PP1q
DTmEB9DZvEGJbZR5nkUqTvzVqCM759c3jMt4jOExmnzba7jnDSAYTTpTvXt2
SLbsJagMx4q2QXuuoK0Y7XWd97MEU5l7JPzt42UYhHna2Gk3wWcSmiHc006z
umYqpw1zhKFtTF0afdUWuyP5Frsdpql+UC6USSASwtRgPQqXiIewbdVBvmBy
24hPtoR7598Ib3NJkZa4Fb8aoSiWnFv9q/IiDtkVwXx/lyvmLpyP0k9v7UJE
x+wyenuttPizN7U6JgepW7e88KhFlmG1kxlhb6py7JcUPdJtz4ZokwMicFL+
yiu3qmbjSGXadGE+LYpm0dggITbD7J6OHhXDvwVAYCQG3W3rqRtoOxakEVIY
kD0Pw8H8NDlcSRovbddaSsxEUZQBJtcneLwqi0ylQDJkRfoBWBjX/wRE+plf
Rpg7lCE1tr3IGZ3Zs7puRPnqfo/qT9C0WW7g5Ex5oFw1u/Cn/UFqjXwyDRmF
xqa7mw8rBHQGsD5dHXEn3jqbEjV0B7Q8Tj8faP+WTTJdF74IwewkmN9Aavan
WSm+rgCvfdUinCrVkMwtCwCCieVYawEqcKVohXsHJOezlYFDLFbg0L/Fyi1e
uJI1sqpU1KGRVBLt59KqiddnFG9zyOGQwSKBpcMk1didFBtmouOyHYMGlnE2
bJ80TZJDel6GtjWpVc2CViZJOKZm3L/ANcC3dN7DMRpezVqym9oARXuLgH0A
6TfUk5v7rCaC1KY7ClqQPzevDKfEikLw70bsFV1JldLxMck4sso9voLh4dWf
mH8bml0BmMxkZwXVGakYFl/0N2maHnzpjhk/307S35M9eWOOK17yrKu8huux
3xDrBW5C7n2t1we3k89yyqbJrKQlUPbrMuCZgqTqvelbJDwwqiLjSoboqO5V
6nBe5d64tQ0QzwTuuMmbdQyz4tVQaQ4+lT5zQiwdfaTDKDuXO56fuc5WMwpX
mnnjcUnx2nFyYp8U92zmprqXJS8tGVxgaHjLanSLQBQqg6n37F5EAhekx5ww
KNqt0LzPGqJE2RHbTPFrj2xRvugLM6BtkC+TLs0bU48oLfq3RYoouLb2uOCf
6npqux6WJX+TqzHCXsTW9Mfh7/8UgPRXMrw5VM6+ob7uO4xbZiNluALOvKEZ
IY8rx3r68V4GQe1/kI8MrlGtRyEc956TL5fnIIbbkNN+Wp813k6iCuchfZHD
XjHqSUnTJ8dkvebc9dcU4s5wQvMYwDws4J3Hr9MzHjk6P5f0m/HJd2/j5DZW
56YDZNv0J1hYcNrwd3jiUxWpcneJd2DYsncBWWnDjwQ9c+fTXj7JQphAGNao
6i7VuwDco1D02WPbsNnRfadHAAUSovylq0T2N+BEkhyDoEq60MEoMU2nGcyz
i1cdCZuWRE8eSbCR7DaiWXXKq5F7NQZMcrX5PzwAbuo61o6q984ntyQsuYAS
iHQADeM4l9vH6qgt0WXjfs2MqHQBWHZ7nSutMPARrSPaD4zBe4NCxR0IiFzu
sQTReLMOsNJxPGF1YfGp7E4j+0Cv2QOt+cjBFJFNchuGcGjdJ5zDkqmjOwrE
smQwkH54u+RmgcgAX/U793wkuYpGrzUZp5+PNpODXHoU8iiUZjE8wNHjqTg9
T6+wNNhqEUw6d1L9O2u52nsfj1zG1mRrr7gL3eXsHNbMLNq8qLTfbPCQwMcD
OtFTtIjpagZZtvO6M2ICGk0juBfAxMAuwN7DNxR1M6eDnyC4qExWGnop646F
mXixyilSiWn8XiBjwVQJyMPFXt+ym3Sl1kdkd6lEq+LUOW5FkUGAZD8KadP9
WeAiOX+D1qYJ6Qaa+Mx9WaP5oT9WFNdfxZXzTqDEEmeuOMynb2+3DWJRfrlr
99QjE7C1QstyFN6Zdw6bQmgKXHUEo5RJ3jCnEc84G4D6AG5PrKw3WMTkhqBh
R4lyMwRSugSzNxLQzJP5s5zW4fd/2YHAdvhG0sO75XD8kSapK6tleBVgyHRi
KzKmOOV4dVMT1q3BLa62uhz5cS/OkTQnbKD2AQ7QODReXTrhPzSuN2pBzz9I
w3L1kNuKyAYhaMeUeNO4QbyCb18V7RKa0lpTvbNehZMD1NTwHlJ1YiTQg09l
LFMR/b10dsVbQTpIjL3O+r4m8Oiyj7vi3RZ6DNdR7HikeMnh6FSl3hgX5U+3
zQHQn7CyLcwNDcN0o5A41H0s7dgnPPNhDeMfZA/G2wXu2ElggtLTKRDjIo4r
+u7ZrsGLe5+btfBey9zfRV5Vev28j2/6littU9VFvicW/VK+I0D1S+xsPJfw
fq9AnZHDgcoXaDJPxVVWSMg4f+nsFIfrQ5BrOZC/iAVaCPkVqON+0JFzg83l
Rp4sFDVzmIlOU84roR2GGorX1aorr4pcpY4YYhMEw8SBn77gc8nd7iChGK2q
HfzuTe1Pvs9QmCkZzibQGd8VdHFbKxlEYpM4h30G1s3aCA0FJW/+ml4Cnawd
UZMb96RYxd9v0ecuTdlV/n4aX8/0yriYgJrW7Q5hkllYDQY/RjplfB2XQQ8a
2h6qNa7Wl7aUN/I+T3S7dBoryoPzwloGYDXqAokRjrongVdDAzpip59B0J8P
rj+HviAzuadJfaBUXO/tMDB6kPrLRrBiVfXXroH0CcZwOF/tJ4ZaxMBnyPDQ
jiVipQtrqPU0f4JVAx8nP5qo/V5UOOEdQGSkH452KHwFe6vAfEaRzBfMFdkL
bFwd/lPPnmuPCvWlkFxPLy+U+d7o0a1cOUgmlhbaW36nlfX/Od/I7ulQEnI5
xh2Ve56xrVnUfYE9HCRV0IssHMVL+e8wptJwY0/v347p3q3XArcVawDnelJ4
phtaIJrbqUrNuqo+gdSHIw0GkUDsf+kz1IVlxvOyBGc3qWNu4lqcZ88CdwSB
JU2rRQO/nwSHKDOsklOFt3e76HdKEhw3VH4bK3vl4TA4vcJkSrLePgxTcIR5
uSoohWYmtbjmPE1K5KpxZjDrq6fQvWvYzzdh1BfrodrQdOfQXcjyumSkrW/6
rV2N5/g9jS4a6gF4UnVgjZElCre/RmeE4fIUj4+tCvcua1vMQkVoL3xo1Mz2
g5YaiGleMoa4UxBE2PoPUlha7BM6rfdKi46azGhr0D1pwK0YBZtE3ra64TLg
oqX+r6OZBH+6J1DBWQDluCU/tneYLmDU+SalBmXRwIryHQ3096gZ9V6Mp6hd
qnqY3geSbmkWBX4s2CAkA4NBmlRo+XlEOogOZzP4RM8GcWjWtERcHTDjpOV5
vBCYH98luLx4KJD9GhaZZbQw1QXZJpyzxTLcLdglq9aOa+moZg7bvgBbnD7R
j5K/q/z4rBIXelsph+X3H9b+2ZNqaWnQKZjSp/cIp/QUkCM0NMe6z279KE42
EnDyq90ooJSYU1NZWgZiGAtQjsMug/Y067ssTXbXtcU6YJxwIWbCc0/WfUUi
BkTjL4U0oIaV6/5Zdr99T34zwhWSpS5+zJtyr6w2x8m5AhZQGIua9Fa42Zi/
luovhC6+jWYNvUlHNxk/7zh3iPYXnytx7RyLQdtwc2UtLKK3Z+f0Y6guhjnh
JbQkvU+pMpll6d/8FJYzt1ZU0q3wqVlfBgOIXunknMnSn/7zarBIugfWYZ3x
r/RN1OsGFxNfo0rbXukL909dsnnbi9hvoQAxbFg9hX7qqjhylU5/s2S9//1t
dnauXfUHGJJh2hQ5JIzbdTEYPcikVTX1RX+gvdVDYSknEyEwKQIvDLSVWGUu
cEFmfcAJ+0S98wRzUKTBOrKpCh8b0D6EOfKrAw4VZgN1896ntcnSUtSZF565
pePT9q1CSdRonF1qYbKhSZALC2GF7a6Bi5umxM8gOnhKNSEFYJm0oftflKFN
pe/s7dUbY1yavOszRXFedzw90x8FKCOJG8JuZxFxhyoiSRpDsAkbZPfy3uov
JguFNSkhTlANs0WMux6wi0ULS0xMEopjRvjh+jxjRCFKLntjc2+ZUSi1dpnZ
D1qgoHyRZi3PrmM/e8FFOM3gdd1y4mX1v4/WBobOWJMbVDemjSxkPIuirJNT
F/7dAaDBV5tGDp3E13Yy7vJzLBcljO6+/MLpFLp0nC4kT1H5FFuvs9c6NbzQ
WHWhL8K1Tx4wBzjHrfmt/Et6mpUoPOtjcAij+k8yyGmE/yOmnQPN3SFYJmzE
LJn9Qb4h9GicSGzYdRgShr97j0rmxSoeIsghKrbtjd8Wsmq8m6ifXGLT2Vw4
z6SiFdFCjNO2j40XhaZ2U2yD4HlOnHPM24j8mUEZc0Ev4xTRxs43SDO9qkxO
zMaUdchL/yUZ3h8QWOo2NnK5Ie0uM4bz0iNaoRfcUpT5Kd60rS+WJ3TQEr80
ZHbaWtOcWo9tKBzOB+rHXven++FT3RF4vCsK8IT5Y4FwjNoLmEhCTc7tU8oX
MwAyZARQpRGDpLHNoYvCYxyh1XrNG5aI/lNVMFcW/rvQ7SeCTgpRniCT/51h
/n+Tpjz2/mt+wrlykZbOsUUhYmHPZ+o1KpF8b42GDSV85CWPC7nLRW3HuutT
41GBc5OEKse5/ANKtLoxpeDGE3T35A4gUj4lqkl7edeYLuYABBosn4wxEWkC
mk2LXGiuafvsf85CkDf8Faifr+zL6njbKk+w95sKuHg0XdZSbowQyq6xTdk8
5mTMO7JUT3LgBfNJjxH/TmM6CMsJ3a4B29F+e8IeEbFdTVVT77qIbncfVhN+
AAS2N7YAXAGT0KH5gcEivuV0lTnOTOg77LvRU2+WzjLX5rnV7aEABhOVwOlo
AZ+LcB712Y8ia88RpebS1sIQCBLXIPGOTC1ZfxnjENHS1j8xPVAkicipoOIr
+b4htEA51NwiLuEA/qc50wxNiG6o6deI7QJE1taEOtul7mZ4jgczrE3WqNjt
wjCaX46JKYFZ0Tws3egzGInUNtJ9DDiESOz8C8u/Gv66Qb0q0T7c7Q4yfCNw
mnK2hM0gpseQ+VQvX+UkryE9h0OJqMr5gIksulQQeDrAeQt9TV8x082AeG7g
qXmXLm0mOg+MKuesWyzocuHrCTLackem9Ih9pMl5BiuAzjTykl9Gd0EHtjrc
EdNWv/o7zGQq4ofj6Jdji4oJpVqLyuEw4yLb+EiaiN2/UlphxqpCNV6MobZm
cEYMXtiOm7FjnLgHuTsa/8mj1bkGA3PoHbGjyOo2rPODNUor6eI+mvjCicyS
7+R5vULX41sEADV8F0sjVfZYQ1HipDmoTQ+WzZfyrPTmNvxs/q389j6VDZaj
N+p4yq8fEbK7JYFYDzV6DpQm5/AKoaUIeT8au6G4M8A79326cTwrLKOQsGA7
kke1FJrq+6tQ6etBPgvNQzIrXQNtATgrB2zzHXyVQbTwH5SODQagCLMy5hdh
eHsyBbEFRnmQWBBm3JEr2RyiW7fXGJ+jU7PzTVKXUhINpHJUquiUaE12T4lX
WjGojbTkgxffjfTTkufHmD8CGpKHFgTb53ebmypdA6b/aIWHsJ/XjFzYtRsK
q14InxdHL46wowZyCZQkviKdFih8j1pWZZEprqIgOSRxI7ME1FoEZm2vCu8g
uqLfqk5qpExpxGgrsTB58IRuxnmnbcp5zjY5IUqzYwPevt3i5dTup//fIf5n
feG/uvfgp8svM0IerQFkzThna6j6fCc33vIE7JqVRkkGYM3tlcXQXujh85gF
mXkfLJcDs486js+75pYJ+AVoyU9vXymTl9QWrlu/h3XY+J0Ky73YIxWiE3LJ
r7KT8z+x9pwwLMu9wx7QFYSKZWm6K+gDuGgdSA4qcGRXyDv/SEn5jDkqHget
9+P8Ngzlrf1VLzIsX2HNer/ePhusKEk6+MJ74PfwtP62dHH3/rtZF7FL2z/L
roD2Jj6TUZX2ADQccrHxLS511EMep8sqWPAEqpOgxjID8UG905UJxngRQfa0
Yc37WKs0/XYoGe+HES59Jau51v2DbTa46w2DUl/j3HTUBcVSn9v+HgTRB4l7
WLEoK4VnYRjqyryue7Cflm35K94Z98x0uevg4dkGdO62feITHvWsgyGu/yds
j+jyNvyF9NKVrzcZ3/Viv506Hkw2E56LIvw10jPrPY1pRwIpB1S5U3op3Mmz
m8EC1/RspRMBGDxumoNW6GmYrkMp6XN1vgb4On2gpj8WHSny+GYA4W88emXz
8kfK65uVoJs7LdJedjkd9IbJPnKsPKIjKs/oj0PAF5J8ITozZnTMw/HJuyeh
B2RnvtIZhNN74ZWv+hNvx+pPnnH3yunqstxMgFBA/R825prUuOPSqiDkhAxN
l/xq0+dJBL4AQlnk3L1IUoIRWK7018FELxnMxGYAi8Cmb7W+s9u+lW0g5ONP
ogtywGSGte4x6LNZMuwrq2ge9vK824KektcrLn0ph8pE+K3rMrNp+N9t6KIG
lFmx7n+FYeVn3ra36X8+DgFCog53aLGKys+lYmFPHf/+KQnEHvH4aipp20Sd
ORfzgO+j+3kpm9RPeaK4O3rstRxZH9UZCELALz/37bCAFdfYw7ta5PWA4HDn
EgujY1zOZhupTLKsbbkpGxSxuJFafhCn6ho/fs+DJDfulSarTgBohDJMYTsw
34ShfWqXzEUFvzs3fOcwu3frh46XmduAGmrBZnlX/KTCQfOUXaywXWqwWGmg
UpWU95kwLj0mRoHNKz1lMOm/It5EGdKjIG4S15xBNNuxsQEab/zZ86ACFEOV
iqde2r8hOTrqbv5RIloQC//UFKC8tpUoFVtkPz2U8OtAPpIE/ybKqfmwSwd9
M7rBV9gbCHAop50P+/O9rtty3Oj3HzU/dpvN/aK/XGGzRbSjN/j85mTd6Um1
hxJPSLXVL3n4T3D0VRhv1kCm6tmricMUzipWTgtzsb2tro6V1rr0YEwI9jtz
1ayUBOmjhSEOPL2wwHWuxzoGCSBnOUjvo1dQth1+nNHFZzsDeTRiKesBQVAY
pSM3bQ8QBDT3hklP9B3Mu2EspjqfBd10GwUvgGOZCrQN8JGx0lY6EW8PInOB
7Cgu38QaniUqsecsHmKeLkY/ci7i1gCudgLsbCaa+wSyf46mIrnMlbu3DWJb
fBLW5IQwqIVeVPy5VbReLOIo8wsd0KxjFZ6ic4nYMhKs88GXzg015/sTfWCJ
k+top2bOLDE5rJrh1z9NkU9KldP0gRp5ei0kppvWCPagDFijK5pxfGdNYTvK
oVC+AQ+uFET2i0+EDCSUjNWMAdH6hVd1zH6p45i+S2PJzu5OSsNal448QOAB
RDqR4Ie+y9Wjpmr4dkUp+VVJHoSeJfplEgJeuf+/AL9ziFKunlFTKT4QpfeN
Syv3cRU2bEZJhHU9FtymZUdSpb/wHGB44NJOrnlshWees/wk5jhms369+Lcw
7FP3BkurkNPTQbbmLYwhA0InFvE4p4AcrXREDPZ8LQZCzaY8TeKhnphfvycY
T5/hABfR4qBcr+EL169pRqWTXo2ClH3x8MwP0L9RXS9xPKvfeUy89QPR0pDH
yz9noyDSDIX/lorBekY/N0/PBzDIikTD8fMjjS0Z1XD8g+t/uwcwrLgiQDPa
RzrQJQEfn5x8wnBN7SfbyIDLkuBkn+2NcmJzBg9ypU3/tT4JO3d6RYlpQiba
xE0Shbk6lUv1eDt5Xes56JLltjxE/L+dxMYL9gTD2qMb9hP/7j0D5dJWZdq/
c8rz1kVK/hbTWiQxGsQAZj9IhUpu2pAt9wc53L9qIRxcSqqThpcZhm7LNzWW
DsmiJpzicd0nWFlNmIoiqv7WqAUTcCIOWgm82q28Um4Pz5Fmx8XGkivm6GM2
cvWSi1BwAX82lH3uXoFvgLIJd4y4+k5fwcCCwlgk+ZAqds9rcsukkqHtqtSZ
ue4UTpeNUjj0NrHelIAlZQ60uPQ9S8m8F/F3QCYvTQimLfjHsl/7r3cNLf7x
nsmCMVS9akXIqf5dPOwP/O7Vut3J6Qd1SHirfjvB4vuo2GXbSA44dqvgl7aq
irbiZDtddhMTfkhG/JcZw5E5bnr7aZ+mw+Dohus3vh8Sts0vN1G3WVJVLOKL
Ca0eq36ZRAqLW22Vevq+bqhCxpGnIhYIJ+6RNFtiVMugHAeQ730es7fjNl/S
EbQiHroKk4iwwPH3lopiplCbMD7YOUelzCGzo/AJMuuPD/Z1JOOT4vzCdtAn
OTGp5dhyZcOphsXhhCNanRbHgtNNMH+1GgXfM/1jk7X4d/CuxMoRr1/mC9uu
Rs6qYBUfbG+alSIycVrKkBO9OamqiHj08cw5oIBRRAHg9uqT4qc3dkEfX/N8
76uQkuzlr8TICl2sWIaER362s0/HF3Az7DY3ZzT+cn3dIn82KGpxLoiIIeMt
3Wy/oBVVXPgVJhW4lLP45GKRd2LmGGdVlY3wmE8bvwaR/TMKrBJRaGObcjKq
sadEBy4cm8cWRLXifDRHIxBhcFeR5si+EogU1TTd/0iJmYAKLlDf4+iQtQQm
MxypQzSqPr4miyual4ktBWEfODe1OLXIkkImEYO0Wxql6RaI5tnrre94ZzGh
/1gRl3A4P1CjnT4yg9F5BlRjcx+tEpd5ESQMuj8DLYzTgP36uRg48/XOY3Sd
nZEJI2BTriqZv3AClc2zIrmDiASR/+Px4JXw9DAbCH4GZFbij9ur9itE4BH+
TunKDvCVrj92HdQ+MaPimo8IQwF1Yhj+KIEVa2OtymVc6yfLFgWKdBzoh+vq
snuAt3SVjpeZ3y89lpqqlhgkWuAQvT8rRIab9j/RxFq88xkQHCUmNf4gMmF3
t5HczntDtyncgffaxSR1lp1jf7pURjHovVATMGknOHnmWdg1fTB4EEoMcoCV
DgU5GAp0EVdY4AEUckA1wf7CG6zRyKeJB4GUs+rbBUwLPB0fF3MwXVK8UdR0
B0DcLysW4UVWz4XPN/TbhSgfvVAT3M+Sl74oYUsDP6AF+Q8CDkGDGGgLt0Vu
ntRaqawVOFxZQWb5P0uK3ryEHoDNzFJmilcT5f7oqUS4L3Di7TTPUTh3clME
GirBMwuPmTIZWa5rydFQBch8gGfb/5YbIX9uIHDf+0VAthrnllo9gSmWb5Zb
WhhcDf8EyLE6L4ru4BBVnDJA8zg/eY7XUy2qnpSiu74xQR7xuc0FGBIQyhRd
RgcPp7QAVapscgxm+79hLRplOy6uTh+DeB3umpK7hyJH7v9J3yc4DXCCcOdW
5VLo5TRKgOlOS7bOuKnQiKO5CedihrT+XD2o0jCz+ezBnLxCTf48eu9JbVwb
rxcfMEKjidgyIclGXIflCpvD4q3mL3piKZw2LGLpSnTB0UUGipYSE0azELd5
0ducjrBdoZ/ZhvLEMMqfbMa5smyFBKoVwwVD0uxITJHrtDVor7GdQ5MR/Q4Z
xKXhmr1EZNGsY3/AczEtjDfAJnQw6EXuqFm8Gzk2KEkgiPMDEaU/DqQYrsRw
kysaK3u72wzZnv9dI+IB3Aki1cDOwIqMqNNolbAtjXqZNX2AH4UlBgBoLd12
HKwfSGmNxK4QEt8FISwUwH+ppftGBiuqusE50zhcVTUWBgD4mTns7v81jnqH
v79C/lTPPvXBEqJvCSchxN/eucMzpi/F38a2nQUY7O3LDCKmkdB2HQKu4H/P
khnQU+0GRP7x0G1/lfKXItk1LrhHBvLGOXew7Ly9TJwI6+pmuueBiQQrq5D9
x6VKywXmZIcB8U1buUgY943pSFcw8/GTRNr6Jhzl2R6NmsSYd/Zkphry2P5/
VwcOb15a79KUa7MA/svl+0xxrXeRrNIL50QmTWpPsL+qcQ1Uq5U/dVy7lfx1
H+ejjbUai2t0e4nPpVVQ1+ycrQM+bU+YHEO86tc3LfqEnDomsFKO9m1ZIlKl
yO2k5Yfc1d41E1HRS+cW00oFvKcKW0luxi/dU08B5yMcZSy1h1Y/d+xp32+l
M+t40wd7uaDYfQjXK/ahRItDiDVpegqLCjMDC8+1zy7bRlitL2i8BuLm2n2v
iJbvOjL/HVx6qbCsOfest8hGcpZe6BqvDobPKNv03XSV3arIrMCh2mEf1R6Q
WKAfiBYF31y9aWsVwCJeE1Wz6dEehc8mvDUxFnGNn20FoL8Qk+QH0T5ydBHT
4d9/PkqsrZok4yCy8GtW4grpZuWYZiuUqqJGHgl4xnd5pzwUfBnhqslZhTxk
lzd8VuFSTTNq29u9ljFe888GTPOp6TEsdMuNHgrhAKG0ZuKO5+RC3N4BvOZx
JLY1K6KmULh+02ph5wLCQPvUPM8x4aDiNI+/Ek2ywdlw7E0d5BibW7XozsIR
KNpRXzUdMFMWPgKGNJUR4vjU1JsOKp4vB2Xvt+fuYNTkuXZnSZQRpvOMgbC4
PxIrIO1kVT0gUZuTLHqFvSVzNn1VPs5Pv5cjtQ8APWXA2kHIn0Tj7m2k1pUw
FFKqEKPCyW/3VMIWTIwhWnQMyMYcbPw30E+Z/pUDr2cP4//Wxy4N+o6gquXa
keXpfbNnOaOx+QwiiHhIspqHENOwjK01mnG7qw/1ichOzHq4Ws+HJupOY82L
QEN5YBhDABKrRV4CpVK/lreusGuYcC2QRai/rmryc19wNwmJHB5/ZzrFcvJK
4MFzc4jTG2ebD09pjcX6EjG7u19/wCTFTYl29JCWFuu9uXODdwzvU9jlxSqU
Opwzo6+kVdUJkCkO2mPTb+iEqUeocSaN0zDcNG+pCd9i4zYcZtSBUQyYHMBE
v/MIEHy833KZ7M0TTu1SEeHFebnO4sp6lbGvSp3X2uYRXmfpqAp0k/OtQV5z
gMppAa75J/8Ouqi4mmOByB2GRdKZkPopIarS4QBwv1UCfzyJgCNl9mtZXGcs
LRn8R5Izh4d5In/M1A8dWNDFTsgyh0YyTQ3nJD2ooQ7M3rkT8LzdelJe0pVU
2xGpAUdBIXEMaEBsmxKDgFDw0laPkPKiaBDzm6wVat1x+62SdQKdoDrP8UTV
ybaNg7vp1nKu4CQizKrZjiheeRHku5+/qa8RjQ0qeRT3y5GoNcswJfvdtpuD
grtJpQh6n5szGsBuGTdUaAZxnxiW86x4CdfbKZyvbJjcF1zNWmMVydyQg+/k
z7JemWDrWmE/t9yoLmqnp50dDAICZJgQaPXLYX9bMbPSAROwMCLZa/E2HBxe
/wddGiZ4YuIh5EoC9sbJ5bOr0qtY36NB8o3/NAH1PxH1hAlrdd9f6Xnh0j7Y
h2d5UQVVyS+U58D815u+RWaePLGDzdWyGNzHeVNbcdA20luc6qzMrWZ45op/
Zk/bb92BorfehJr/sgWlfrlgbZ+qJc8lA5bPMpPu9NHpHxKJZ+cBz3/KHZJv
bUXcC4KwJ8qL2LPjnnLOY6ikGV17YiJv/3vmEsfMqUkomxlDbWYXBQj+k9Ys
Ev462BP3zy0GTDdvLB93fXRlM9oG39a6Phg2X2+KuWIKHVbMWfe2Y+uOoNqR
t4JIvA3Ujs8p+Si+8NKCSwayHuYrnYb0aVJADsrFZd+ooVD1+vB71jxXz/X4
lKNJ8Egio8bUDPHdWPbqy7mcJGV+PMcqGgkCq2lyT98hvE/UZYgrAwl0ikiW
oFuJdv3T1pQRlem8LkkQZQTURw6zrgNW3ZLxvvOnfK15gx/+TPzX2aii2Xt9
N488N+JfZUp9Gn1BaxnExd5f+76Tj2yrXqbSgi1h7hhIRFZtOzozXI7P8srn
yT4pGwo2jE3B3w9CK649NGhhYTKD9hZuLyuHtn3GGAUrMXVpDNJIIfhxp2j6
DRvs8cw1JiOx5DHxoAaoHJUpAvS8mG+v+dZbgRTXM9qHnt6f/paR1jYHRRhT
h1ilqJWX9zr704rIC4sHdL4DUFMB/yqPJs01ZnVoj9dc0rG9s32ogtiKA8kS
uRQV5GANyx//hghmX5aXZJGhBCElvrs4S9qUKRZdZs7KjMUWhfPhP9hlCEIE
Hp2H5+4ev2nsFtbdJGEw2VECqfR83DxSfG+ttokhTVwB+pM1FXW6lOvD18I4
1dY9+v6LAmkw/Sw7k8dVsTZhT5qLeoS3u5r7aaoKDuVWM+peC4W1fsRxOo2c
OQKvNtWYLteXbnR68Dkaj0N4YYPGZIHwKehkmeoSHQZ3aK+uUtGiTff9OZNW
ikiGwJKu0rw6KdmR6taY/I0IK6hLEPIJ4Yj6u0qiGhOIzi7mKfkvhEPdZ0sN
+wpl/XROqmjgP9+QISD/byd8s34/5ezUUpuDZBJRby7TLIK/dvuws20vrrjj
ixQsEUK5O9Hw/CT7LyjtfAwnQsnNwmfFzOTQ9mLU/aTYZSA1ggQ86vt/GDrj
SIzXCHi0mZkgHw5cNl/aM8K5kApVO2YmyVf40ERDO+SXJbv9lv3k6NzzaEYU
tX0XurWol94YOerLBQ2cnu+E5bE2S/HJf8B+PD5MArrXYIs7AMLWkUHgGFFu
I1GsszmWfCfLDfdxqgywzgNI6uzCfc6/sdjp+oB4ea1yufn3xZ8awxh0EgFH
+83kzisa0okQCzLZohJBztNa56/7jhiD0raTedJqSqBWrUju7Johpn0kzHHV
lX2FRURUSgWPWoh2S2RujhpplPh4gnijpB8xW3S3SGfGOZxK7q8ffRHTKQDw
alYtPxP/F6DoJNvPRkbpFNhZpN2dlCUlFcBVBKHH2pxzP4HAvqhBnuKefOGn
oOO3n3onjWT0vyfsM2TBG0bb0uda6gihd7G8z9P2WCeoUYf96C6/DVtVLAew
3W3dt+hvNsU5TQXwKVy5w5aaNJkj0/KKY+CutmP+PnzgA2xO+hY+LFRufY7a
7dwXwafQaFYkMBf1QqgLJ3+FYmgimyUm0US4LKZ/RNnswGK50UXofi8p+AMs
NT07frnGc0Gz1F+unlS+W7tq1SS78XiZxkAXRvSk52MS11WQA/9LxjNkh7KK
WF4hsQGFEpYRLUXGVD+eOPaYvdFV9vj++KtJ0x7s4CddJX1amzTrGOBTVB6L
F2gyOCEIQSCL2kNybvwItI3KC/lXu5kBoRxUnF4IdfBdrSFfnISKNWKCQRSU
cs5CpbEdfnoUCZl0S0gGqs7ygBAQhYrfhN5VKvGrBiNq2JqJuqGsWH3mJV43
1qMD0sMZQwPPkIcNy8J0LZ2F4Isfi1bFKyLxv6JTsinlxkeeosqG63+KvZS1
hxw8Km5uTI8jm54+JwodeH5t6i2e701rw4HFXvhNJKupyUlZ68LI0YFUea5l
+1PjbDsXgsa6kjolhtsUWmn0cQ6aPfmEfATYDgRF6c5Y/+Tn7fsHqS3Eg8jJ
nJXRYyBjJ2V9NLIe1huLoyICFPZY/ng+xHh/JYGVRhQX/cnvCVe2QaKUqBOo
ld+RtQCyqLG2ds4j25JTfXfi9D8Ol8yp9z/oqDAhOBSI20610npqOfKNR5FR
HvArNxPD14X7TqZFer/XVYJ0ylruiYuUcVwCoZ7+qfv8letMgFX3s3nSgB2U
g6szksZk1zhnRkkbpnIhDU/dE3p4ngqDLfpkXrE0JXtTrqC4goAH3NnAIe1n
8jX895KkP5Zp4Tv9raiIfL7F1ioIOFduQ5ZzSHgodF0z1npFmr+gdSK5G6Va
6ZEUKFv2G5t9uZ4cx6Gd4H5D6VYurl5cm3d3wBKvTDWEhryNWGKofiAjGUjr
yx9P+EUUSiTIrPxJgNoJ8bX1eGxM/+leqJyp+726u+WihepAXVvHQLUpO/Iv
XbiicJ4Vmr9m49qIS8VFqCtNpys2GCjkdny3FvK8Le9107Y7v7ckXyNj5lzb
Iup19FTHzaVwPfhaC2x0Tz4PM6yA98WX+bD+YhAc2McgQ+/dVyTCVHXtLz9h
n6HOMLpSti00HWsGOPcNrd6oyf6HnFmYMAuINo3AxQv5NrUdqJh+Gh74QP7B
Xg14QMS2Km2HTd/beQ9S5e89QQs75mJDenuSfh/S+gY9BqU8j5MWMo2hkykz
sU2Z3qYY1QpKw4Q5ImdChV9QvtjJ7fCWETBCYj0GRAyVzZdeD2O1jhig/CpO
5IZHOyDbVcOLb9ciYp7s4oNXpf4Efff0Vlw5yIMHLkg3CoWmdcADQwKI2Fja
Zvd1ljun8W9frk+VIhkdFfO3z+O/AelGIfoHcK9dbMpnWMW67v18oIuqWsfc
7G/txQg0cm1TwCn1Nfs4LXvrl15D+d4UeJ6rUtmzVY+udE9H3j5TZDSHocWZ
EXj+DtwpIxApFvtvkiwH/MjqAS1/tf+jU8QWOGd8uqYM3z9GgpfxZzsC39gA
7JLsOfjLWKI8ab05/WG1pfGmZzBzsNFALMfkKfpzUcaL6wOFJ8v5dWZNVN0+
adaj4cYVZJ5Y2dpxE6jCvryZ/D7muBTROAwErziY7uIuD738WN3mfc4eg58j
H8tONbext8cnvbzbZp6FA2WTayZk923RsT+PSzVUnyJLuL8CFsA/qwnni2+k
OjcLjN0PhErDIyYfSSlEmUp1QuHoRwrtmjFpoOZzUb4iya16qdmxgnwG5DYD
lD2aE9BYet5QhqIio4AlnPrObRTEhpdoc+WXGXbMkfslqtgSr5v8hQ/51n3R
C4MAUwax+USeefDAS/nthrlSnV76JjJRq25100+ebMjeG/HPfXY2qr6aOwRx
RB0xJ44qApjK5KiTOQG4jHvYwPYYCY46ulAjdb29v9OGVZbSfxWBsrz3DktQ
fzFdZCnPYHK8la5cEPpIVan8rnqXGtnuw/VSzBmllVQQkfgo3+Olid3dTneu
Up8cLCgaOPZI+Ko9lZTxk070D0sVvOSH6G4+bT9xSsKMq6NSuA+hrqFXtxGJ
1IvxfDlTTSTYN4a86QLSS5cmOsgbHP84QzXobz3uKrfuFIoCAJH2zG2ArdUI
dFO6IIjee5xjBCGBKz7okV8xT6AvBlPh6F9z9Nl1aOSwCqWfIfZLYIGrstN/
7sBhjR4j686hGUoL7k1hLi3H9Jnp+p9L2bNGg3YHfi/KR0ZKIUnzZ4nVca+G
Fb/nMfbqa/WopNw/mmUGShnYmUyD6dFlRa3gssW+1J7lg3q+2rTpmZAvO/A+
V71fFejRdGi21PSgfl9LzVX8GhzS8B/8/Jmwq5FzImk17hLh/W7xrYLtHWlL
xNMooTqCk0VHwGorJmlwa7TQqX1/JBmkLbAF0yIJTP5fjmrfbuXW+HxuQcPL
NmKsmhirpM7ZAy73bR5XgPlmT3id/r6IRDRtgU7R9guoRJpPL8rgXB+GWVrv
796FY1Ja8kmkcIvPdBojYCXkOZuAybbkV5+24Sr4hMlhQcuKcYnON3Sz57/P
kkw5l1P/KqSKHRgg+xXcFgoBgTzn5g2eQBAtslNL0tUaNlXh3/MjUz0XVW0A
vCxzEQIOy4363a9c39BAjeDN2eed/qUi4vDuAmzTDOZHHxhQE9ZNIpE/MU+/
2jlZpIFdgfOSmhluGQpxEZwTKqEquACAI16aCMFAj4UWHyrLghdVKzQ26gXE
tV4O96TYBeccM3DA7bd4uTQFI/JL8zY8Zkwr72pab3DUpjkoBhlAHRykwyGS
c+qWBrxcD/6m4mWTVE9uds+uwZp5KEVe01QpjMlqoQ0CaCPYcMXxyeT0+X4H
Uqz7JvvoytiJbqAwfGt9SQOw+DlintRmLrG6M9zaVq6zYQhHBDGeQh7yz8CO
DGUsXqbqCYBpkDwjwiG8s0FPAN61W6jiw4EY8qbOdi2N/1QHESNWqRkC7nrG
W7G1rV3tnd1yNIILjrbRzzwdytRoLCa3PtCe1TwH4qgI6OXXT4fbUh6POqrm
EqXGC6lYRy1OYYIe40YiK3/98nUgwiJ6QhdLRshJ7W3E2LTCofNJ2vlsqCJC
ESV3fudmRpu9zk3hcrdlkJkaAdxenoHIJZ3jIwHP8zz4FX33iro9LqQ/5ZtX
924zaHTZSe7ey0CvlFvWzoYs6I2s/wrrNAqEjLs/W6JbjuofG+gPe5DhAahR
HEEYv9l1de0vx9hpq3kfI8B6zEMFJvARtaQPf0qzX4/b8g2T9SfcVIZ0Vk+c
uaaRMDJhKiwXSZhGa6/RlTa/u/LLDcv2QhFewUVmx2ynUhZhUskMOeIu+aVw
D4VNTWvVTAv8cgmCaRFpbkZv0ckzvzqTRSm/qkOFwGyQtegv8o83z7q5rHek
TI+GbBNlYhwNS3686bJl3MouzE5w9JmU/SXgqCS0fsSOTDn3GtQh5FCSRaNS
+bOXnGw3TLtNChjgI2ZfMtqmVSa/C4y8y+weQQHlQQbw+ar4GjiashK30Rpc
8pZBSuu6e8jUkZwlGu6ZcKu7Qr/zQUE8SOWldfXxzy1pEsSQ51yxJgz/kyPp
AGOKlTxix0li3ZTz8n+xY2+had9P2bhdBT0UxaH6Yc+XN38bBhK7g/xllVX8
0D38eu/LdVD/peG8w40vRXDVeIPhe+neaigcP06axnKeD7kUJPB+EmhfAq7m
P33wdjQIM3+it2ikq+knmtO04tyynco76OWkhtJWDx5vH8JzU685WpFJ9Wc2
DpEV0ORtwC8czGhZtaiA0WXhGn8osjBkbokIxyJR1GvFwaMZ8VhTv+Sbcv1n
7VUgRDSFlzd2apbffmOme28XPWU2VrFoUzYIxl+88fzrr/CeJ0IF0QZWnOPW
yEasRvl+vvl13A5PcDr5U+vd/CgUAqgrRuuX2SN7030hKge3uoOvwGMcCQbH
PQmvyzFRfiCyIuZz6QV3nE87ZGV7DdF4C1llL9WWiA/Q8dkARAtZLC1S7em7
4oKRiQP8zr2Hey9DeYJqKMMrVZlFmXrbkRUTuhN8VhMd+eYAq/TAw61G8S0y
bgYvlst9HMpx7sHWnTrplhs+D2U2Z2bTt30uHtunrLDVVVdceZnjyCMOgADk
FOhon7TCHTRT2+ugsHzCkGBgDInIYaaDBEQTCpyfwzrEGjSNu+m78m8G7JH8
ZwKiJLTVQqOPL3NAJSScbrLsKbFWAqISDySRNw2VPb9js4pWbdE/ir/c2kaF
Ntp/ag/EAOaCe6Rg3neDVAObKHCO6m2Tx2BX0xKu9Vo9BN83Ju5F0orPHS8n
vIGFsjRtGvLLz3VtK5SFKLTlekGEmiBRn09zBfkUW+ykYalyTRxgSKsDLpvV
21vsLff84SVXMRFwVfcTla2F727Q47Mc39kJNs1iXi1ktXsijPVpXhDkgBZv
FMXx8VS5KPNOdgTir9xEbZifItIWLOmcQmbPo0tLqmiAYIWlOiYAtE/pY3H/
MRDf4zDgdQ59yV4LazjBbW2DiyMt2t5uLM9folK5XxgqUV5lhU3EeUs2cSce
QOpV3yDIxI+ZFMMnNXqC44KnyZ38ez47l/avgfv6UauFzVsKgEhyNfUIE1Ij
hbBzJQ4zeSntoB7I219m4kGsNDFMdSwedM57OEZYuTUfedL9lOhmIvrakeae
Cr+vUMUkSbf54QV5ZTiYYKazv/3IK/bwA1MqkP2KeARhvyNJrgVHoWCRtvJa
uR1qAGO2Zn5QBdKirTUH+aX9HeDzCQzmZhJj9T5Lx61EmY0Q0oE13stQc1lb
css5w64y4c3A7hNbZhn5mY40JnnjjssKwYrZYCkcQjzw2YQiDGZ8ZDHNzJjA
FKXLpNF6Ibsw5it83wgPzUk79UGxFwKJeZeyt4yjpYBEow3tMyTAQVYGJykl
9scIP+rMKFQIe/Gk3vCcyQs3+TtpnSfpEV+obrWQDCMsS2DsjZoYggPASeXj
HhqOCNaFLzO83qB4e7WymawNGcJVtBceCEjw8gpgAHg1J7nixc6FCqFhijfd
uQ4xdo96p8BnBh1VPqnnl5hg7YgA4A8BP8GO2QFtVI2qZOXCIfuuTr04W1ES
LVAOxZbkcGbntpUkYi3o0Da1qga205ANPWnnAvJ+zHZaRCgnSMWrY7ZOBrSx
mP77qtTdcAvir8pP1AiWVQtObYIPFzq/sxHC3K4mmIKPDVGQd8qRo/yQzrzq
1kw+7sX/5svOrw5LNMQoH3S1cUdMs9mVckokOitWqQ37/ynHGbdfn/7yk8k4
zDgeOOm17sLGo/KiBDcJ+SNDdqz84UXiKRzQb9CVHyb1LKdj+MMj8+jeWYaw
NpccZ/mppLbaV4RG+ETbxEHnafYRqqklKrjZwurm+QC6YA8miptpTprLljAd
e4vEKRYetQ7vCcspRAuby2BXdI+D8WZP7k5gnrka3GKeyd8sFEryyjbYut1s
tTC9rLbJHOdhkymJqvHHSs71Z+Dd/ONfpvIUjBekjx8spnLX/ybtGCAfvjUV
lmc2oXTUQa5fwwDUosGPYxnFlD2fcZQd2eEe3pzqZ4L0NarMM7jwxW6qciFw
RVi9UtL72OpDcjqXIvbDH0FK5wES/iIZlhqz3xrj9XHzA96ZH/fNziYtCTO8
Dp/JFCwJ2Bi1Kg/0+pd+RHrunucbEZJ+y8mblz8yL2hwPCrTZ3NFCSIVXNoB
xvaA6wLqivWf08SdF163fFfrhbTU3kIx6g23ANiChqtCZ3nzOH2LTb+Gqkep
XIvJ3BpEPJnGJ1p4I2JeR3ndhVcQicKxvOnlkUdM273x/tfvQNLS2itnebIq
7jMLW1R3tpCqGLwixjDL4EKEwYVyMvPVNULbHk0dCoGSIqoW0ml1VrfgyyMM
v/zbXIRr3K7XEEZ6HXHNVg18w3Am++ucTvy+SzDieFwdvCoyeRLUe23yzfPT
bzaDGe26wSzQKBl5RL0kOoxFY0aczTvjkIBY+kWQbRus+D0KAq49EJCNtI2Q
PQffexuPWU5ke76IYZM1DIj0JapNY3X8acqFGM+Xu9XCK1P+BnWuFGg74viF
Sno5KOLCscEHv8R0Km2qewlv0EKsgF+escYqhgF6Kov6Zhq1YzvcADG2zkcD
T8+Km8wOxQEbdyEfx/y0azyFl+3BC7bVTU3sEUoxks5pk6MmVrPGSxuEkx05
SlrujP3EZ5Xxshh25zmvJii/ClVWRbemxU1vjY1P8NBXbo/joRWQowUBuyYf
+0wwKCdvKQ7BQwvPWN+GXzV+ltTmjwLWW5Uv1nn6TH41pWxyw6gaesJ0pyD1
Gh6xRTikrGdSJ/MPrF3tn4cmvNZRJNvy60QzdY9afzpALZQHnH3nWv6WWQun
4S+wrSibYPVGaNM0XNe9ICohkMv/zGtla+/IdUOUo8kKBOmPkOcMuRK8y5NG
of/oJFEPgqYl+pn3sZ5mWdGHmGB60Fm0yybBJ2XLGYjxP6bsMCp5bZNgdaeD
iEUgcSRukB5u9qMSzENdvFqJx5l5x0ChJCmatq/t/dwHIFV/YqXkXvhrVJrE
O4C4l97xW/OyOSmzsLSa0I2BXQ+iiiM5MFK01Xpy9dTIV1NEmY5fail+SDDS
+1ACYXb159AI8GT6sRbel62m007+iNJ+FIzMlMPU2mTlHqfrGwYEQ9XlsFig
6XjGsMv6o5jJSMwOrqY/XmrVwoamoH0QQ3du9mOi/331ce+tZkoQCtnNnu6p
qG3lcq6JQDMrbElLbm6yxp0yQ5LWtauMKLSyA4qLSnYaLBdkI+Djb6F2EXzM
WRVepqKB/15E2krPtu33nkZyDk78kK/q1ea04CKjLJZ4D50eCZ7n6OHGN221
AjDZfH8/g8GpEWj0J4UGNWZClFeSXFBAesgbIvtd8B1dl6XvtlVJ3ybnmmh4
8kyJrazzQdmKnvZbwzp4KOhIaMxQ+HNA+i3gTN9a/ObFcBA9YEi6ZVQVF6gT
kf+ElAWF5RK2jNH64ulByjOS/Pyf0pVeDNEjWVqPAQ8UeOcv5K/Hudi0UX7w
RLusZJdgBfXrTHXaGTq8vfZrKMlYD4HgawVGSx6yMijTbzX2vxZxE6wl2J/M
TEAy6g5VzIo+HVLQ5X4gCOod6sIl/RpBPNpppDcDe6E+haMjG9uq8mfg14uw
WE48bfk5t42+KHm1ZOwk3qQUr8+qrHYUVfVniK4LC038lYcBCsLeU3vxIuJl
I6o2m313B3/ZQ3BidZirSxep4Kdi2L6yAwWg9F1gkCAlILa4p9V6wCdpa68g
GlS6l+KoP61b5jdl6j2AO7FvLQSbvX94uhURjozU+gfb+4WYHB9Mi2ZUupKB
W5hFT8wVlWlpc6omx2Zgl5yJbCwSOL9iFuRRCwdD/ZGWWYew52I440CNtYO9
6tweVyvIji2QD4f6dlQaW2sDlI1bfFUt1mVufq249Z+AjditMixgbZaIKNH9
8u2BcTEh2gQ4qDj7S3G4PI1y6kLbjjVeIMZ4eZ5BU1smKFFHCZ/pYhqKyIVT
9TCVQDGAmKUdX5cU9cMCPHN4fsua2OP4lHO7m4Ss+Vdn594N+IfaAwBSc6Ep
8apSIMom+ib/8SYJ0Aj7Nqow8ehjLYgG3g/iKkvB+IOBcqzi2VQ+Tx67GWqh
yg5QtIlzu6qHcclTJpHaXZZsMz1BZl0COHxZDOjsjP9VNoW+JxbsyBa6cEI8
LiP/Jb9vz1zfU1+9ZemP5ykxFXhA2an9cRLpJpwv35lRcIYfjhHByyw6E0ub
E1WXGrhM2wuPh+T72e9RwoFgESLRr1gadMX7leMxWUboFCkg/CKdcF0+mdZ2
G1jS2TpbT774obURH7XozhE8X2s/tYtakmKh9YKrf5DTnYE4U2eqJZLhZIu0
exEkWtl3QmMYRMqpOtMMTLBvC4QrTnpEkVDfyyjRzU0fpOa3G8qXXIfeQTVO
ynCZWcQ8KYal9QC0hcEhNpTDKChcz4ydB1EZ36iKZB7/NLAvC2cMeEKMsQhZ
9svmsxvi5EUB6tfDnC8xh7FthYmzhS+ERMSIrcRleLtkkhQPQS6wl7HYe+j4
au/SRuBT9pBpHUYPGLIEmS7Gq/D2y3cZyl2BZn2b2NI2Kg7uqY5TDoYL7xi7
UfS0oPAoUH3nfOSSQRFGztWN7GhWbjXqURgDkIw+rxNqgW2mI6+e6em8Sqt5
dhxbAVZieOOKzqrjBXG40+zSmfs9Ir7gJ4PxFmWlGj1fmBkxrWyhjb3dw3FJ
QsiNNawEFXh92fFM807NNbJYj4+lBiqz5vBzeFZxbFVXnhMyGHzdXPbUvK6X
m/7Jb3M/LGsmmC604Syaw3Q5kI8IHI/d2fZ5ZQjXHVyd3/Uv8T3aoE5rcNfD
Cb+cg7riDjg9/PlelytZLq7HTdp6lv4TkeN9U0CCszwe2aEf5nUe8O+Y7WXB
J9HsEAxk31UsoezRt8ROHL7tv71PKHunc11dM8cztkIEbPd8ZlhzCVENzWkX
hRYy3hw7+0BD4+l2SoX5rFuXhM4InpCqcXg8liXwfvHVV/PRkgwVsLPWGwO8
0ncLTMDAMSzLMgtl41+ztpH3ZCqtAl0RFHEAnn6eHCGEvlEW1Atb1RY+gOBF
tIRx1j3mm4R1CIvr5jrbCXS1sJxei2oHhwGEH8IybBmsoj/8JAul01rBQ5kl
/7hrQoGuyGuc7RwnLn6svdouPS2Qq+r/ZkjQCaZ81Wpgh5HdbvfzZXkUTjXe
9td9bk/vocyR8GiLc2KSBLBjHNgfShX8Hu9na2BqSSkccY5XQUsDFSt6pqdH
jQqGSDBUanyMm2pfpTh8C5ejZ20B2/ymUfH/stZWD7y72CgUcH2/D72YWgxh
ehsDHWgWZi0E64cYtxJyCazZvHc6NpqsDrRlHLoTzvQGiNMEQRPFQ8Cw2U62
KWDqR2AejfGMiMDt0yimDRVsoSGexKhk8MfvDzlnvMT+5ldlObMHla9IE+lM
okc7molsZ6cRESp7ss23cqIxGYWg1PJ7AdSnrwjIdYJQbg1Zhx4jkMmyO0vz
V1EOC6HetpZRN8VQM/ParklEAEL9wtxgcluAPtHnCanMFQrpfNIloaS46lb+
cdmJMaIqAxSlI0VQroNdz0AQcrI1SdfDt1YRLo1X5ZF8SOKZqbT+RF1wvFz+
E/QDS7hLPMvD+NzktG5HG1cIeL5OWHOrv54dAHpBnS9QWBEHXsYBJ6js6kEy
6wT4ZTgnWLO183D8cjpp8RnSr5+CrsX57e1Zb73SP/V08ogyb9U5a5ccELbe
O4a81xbPEidn3devY9CzyYSMXe1k+6JHw+fvxu7urOJQ/WV4XR8GGng11trh
zZok7f/1fwBisVXMRT2X7xI6t2qniTIF2Fd17pnJjQgPtAD7EGYMDm0d1KG+
+0yFh0eIEhLbe36X9baRzjvUsEcAFH4etKKM6x3zUySdZCXXEdU3fdb3Trhv
RD6JexMv7KLXg8JkEzk97SJtcr+73k//TYjk63U7nf366lr1cj5jMHH0t6hV
u7ZQ16HSZFOw3wQzKnPLhX81yy8nh9OltmqZhWpnwAJS+p+DXQ+4XLPNY+rj
vrHqn7GZoV/0LicFvQv3PO91FjFe868Fp/a9uLwVQQq2O7TZUm1cuocWkmbL
jaeKBbuHrZW+FFN0qTFJ4BgKDXVaepu5AoVfadhAZMNYAWOUcOaBJ3GzoUQU
NOuOTx5Z8mfU7WQ+o0KsKX9vTg6Nqiwq61GKGFd9I+O5hU+1JvsZ3mv6eeB2
OpkMRGkQGYoCX16wCQO+taDXN2tjz9irEERi3UV+XGl2lmMENJu5RtZGidOr
pvM6/kv8TwPxBiJyLuShsk4FJdlBpt+RT6QatsgjcE/NQ1qQ+u5Fl7swPdVM
5tWCEDkCbiHYtwSr/ajzP+eieB40nXLbRvnzF+2baTClX1ArHXLhKnP0ZP10
Y/9z7SDb4LtZpnBeo0oL5FC5vW7MOuEopJdwidzfrwxM1/GGX9Vh6vtUfCwS
cNTeqPeId4ju1q1CvhcLodNmflSpp6YoBsinh0gObJS2zVBBZaxcj1MpjwSl
31rtMMOfmzO+2CwiKybBkeCkhL6lI3B4UA/V4sz/Nyo3gvJc9tc0A8sqqYAT
g+aW3/ZJokPNnmJbkh+nWHRA5xwFR+RktUuLfsi4yCU/mZSL/LBRYiLDByfV
ipmKxE0Ev3A8KUw75rbfQnwmFTOrg7qF83Pwt2vAcbmedhz+Mfek0RPkdZg3
DFsnlRN8iosr3idQBoWdYGIcnMAF1SAsC/KKjzQ1Ziwa7PxtUc8fDWmXKZwr
K1g1ZrbxCfSz5BqsZCiktPGzvow/Ef0VVymroMGb3+y6rCJmSSAo81QN6XEv
s0+lv/tySTtz2VZ1+g0Yn+WDAa4Q+8CyRBE/X9FmBVYZrd4LYtvoXoNO/KL7
n0VghY1wwjuo11xtuFXlcQX4K+2UJCBGgRINN6ar6/dz0Lxxx1gqAB//E8xx
HkiBo+4K/3lAL6YeBuQVpwzL3wDqQImgTBR0BbZBG4hp/1rKP3wYs9UrYyVk
O0ABL6zzaH/4FwGe2Xou0DxGvVfmxzf/6s2qNSYLawMxrAPcsIssk/7WjHJE
ISDmn9uwoSpbZ8o/2RWVmgudduRktJg6niyrpQtYWOV20h1VhCIMM458DL62
WmI2gv0Tp0CZMXR6iLL9bXh3b2C3D0KNZnVKhjEdapi7gCyhNcaM7wc59Jf2
15MBb9Udm9hatI5uenFy8zXKsnJoLxxDhbe3zH6Rc2Mi6BiWPYxGc8VNBVLR
XRnjHtfyNncd9fLuvqAvLrWJDZtZEdB4LMbsd3Sleyu7a5RRRjeniN14ME0A
A9sjXLPmoBqYa1BPV0/a63umJnlEdz85sncrId3HO+1KaC3D6XoG1p97+h2r
Pt8vUhF9KakFq1KqVdLo079W27x4wvsS/fILlvq/Mvu32CFsbS7jPAc4WUoR
Fkw7C3kuOTIqMg1GF147p/1tFNOxjqFzIT4JYDAemnK8GEVKsWx7b0MC8ni7
9GPe2aNlEBRrPrG2tTinOzPDsfFYcQTQjMN+6Bhx+mJ2UlMoLBynJ070UdBq
m6deNrNuNAyn69TLj5UTKIa0pnxQDkMRzX1GUkSGfeym6Rt2rMe4fqEV6h0g
k0YXNwTDWzq0qavrwK8AFlcgQ8YnjZl/yWgsgc6moc6vKcOcVeGodcQK27+P
8CtX/g0qn0WBUiFO5zzsu6jeSBW/LhyO5UebDBSAILr6ooOLh12yvJHypVqz
UU7EaOoty7wc1WQIl1eVZBqNEdj4uEGMaVfpoNPSCZKkL0d8WAHfj96Umu3K
ewyM/6xwRCOXko8EWa4zqfyowgDTjOFZlk6vRFYWQKBdvJIf5UeGU4x+pSP5
VAtZTInS/FAIbg+kx50DbN0K5Q4RJsvU43pNPQVxrfi4PgiGdKG/pc4s/k+I
HRxZkmoT+iH7k4Y/d6x+xIASXe/dCnsE4fbbeS3+65+uoAXgZr0jsqPsiDnd
QoOZ4hoJRy7glexnbpxdsAoO5lPFr+LmM4Ewu+xrmcToR8KK4puIkiFp/iDE
mAADFxBkRl95ldDCEhDssq9Hyia95ChljVdz5ZjvaLrvQ2S4O5PFGCqlayO0
/mzzULJVhA2WaTAv35EXEeVSXYgU7r8WLacy+z4EppOrGU95N+e6KIiQ9Ly2
cu9fjx20jrPSjeX4n9UsRFj1MwNQF71pmuLLJIbj6IE8felE86jTxyCqNbog
GY1KRk96tenUoWTmZdqyNisnru2+65/rj6ejKMJFDV4sgwuQjPnZGzkaXyoX
Nk9TbmrkR1ZXawio3X8zilwo6Rp133NTY6HztBAJaOLmgStZA1K/gfED6aiZ
5SbYgTMkaNdCRITnnfLQ7R04wZDVJG2gbnhtcxkbig/j86VW/4OdJJwT3gDu
EYUGaEz/WjkFsZIxJRKO0AyPwDSe9SLihckevIwEFrDleCwKQHhqNIjVZF6f
DQZUlGV1edlwLNifYmDS9+Hok/8aHNs7k35spRLgGuzzIBSChYAoImLl7uGK
aD8h83INDEyrM+rrGfCu8WpKbsBDVqfw+f4ExfFay99fZhI4D1bBvoyJTya+
E+aJcdB2eNaSXTymnfojd60V9OMRhqT6OGCJVp5yGb8DhMqHKHKsyzxcA/P1
kuZ7MkAW8weYAo0SyPi72A5fz+A6RKvEyaoJQT3i5yKHgamIFkLiZR1wfW1B
shRbkNuH4ouKsmHJEEq1QQdwDCDeOCX26DLbrXD1nTe65jgZLIJddQsPnti3
IaC5vGpSh/2q6iSr4hiEZ4W6H9NZxoFdbKBB7rITEvD27OcAq0QB3MrdDy6+
0npWc74tGuz+tUiGpJ1U5IpsxZ48gx2k0BqFh3IQRUtjVnme8IAP7h9kBraO
oXNa3KljaCwyHYgl2lyEBwH0h4zIU8DPgO2UqdGQljUbHKFjqslu83l7XjhU
+5y8qubjRBfivEgqNJ7H6OElQqAqa4SSJbjU+FB3ZIq96Kv024O1vF/k2K7S
hKmtitJsaV/KPdlce7b9SD7ptGuAwtJPMAhSfJ0VFYm6f0fJyGtkqcGGDSsN
D2s79MaU0UHe1473Qjw09gMpJjaLDUsKxF0gj63qgWLQdxuQomxnhZE/KrSk
xWgCPf8k8v+V1FE3fnxPjh7cfQM+LbyzY84wRXJrPxpU4OINCZmgvPinlhET
ANRNVjoP1xYU3zumiLHHGUbnV3lYUbVYTvi52AQoqewlshD8NaLppQTx1C5m
ymPScYsQM5vkSmHGI0rYA85G0ytLI+TrNSobH+BE8dcurtsJitVZzDVST8lR
LuWJR6tFVJ95T7PK6aYSI7Jor9+Ene7zO81/UiznrgczTjkUwWF6hkG5CTYc
pCIrjkA6/y9ux9PA8VMCQ0afkmE5yNjYhdNAGo4uWC3+FPzzIWufMqk+VyFi
UGNQ4ezf1luY2yFTGHqK7MpaJMNissfvO5TbYhttYNEAppIpFOlQWsmBcJ8i
BA3dTQNd7sF5OH47+/9Nzg9FhJz1MgzxSR2Sxrm6UQOaPKnO7AfKa6vJnHzW
8wLh7yhDMx4FDQrApo1/bZ5QJFzf4n3G/aOq5MXh/JV3ftJN7xG0vvXjC/L5
8PTeOQjXY2daLlN0uAFrqZcOkbvV16Xau1X369nby8DNvmZcaNm4KJhOcvP7
i5i1dgmTx1Yq5MWUc1dMZtKOXq13Ih0ZUkmkWG3vO15oCj3aH44gu+ld5V0w
D46pweV2W1llH9BBccYq2gHK9XvuUuQNM4UY/l5rdlQPO0i21MLl2FiUwcCT
X6AxRbJE52b+XxxI8LM6pNeFz9LjBCyENBfaBk9zDibBr3PhP7+Oyistp+Bz
GRizJN6Jf1iqiDtw8sp2Sch3l3noePel06uU+96RUhPScpPBHS37nKRBuJOF
aFjNv7EzcTYsR3/AoUDJmWYd6uRfUkSNdK6xyJn9fK9hKqNlgX76dZvDbOmG
sebRjkhACo6o31bnxxu8CRzdLriZauQT5mFhnHNaWtrLIe0JcotGk2tD7upX
XRIvbGNWs3xtMFTLcTJfwSeAE1L3/ANgOPsa0qpWxSyNFCe9Lh7DPi1jkRRU
mrfz14H+4TQgFLX3IVIsBiHphaXRoTMXY9Wivx4T2JW5GcPblAk+HNpbYHjj
f5vpmbBLRUBmn0CjXbxB3fwG93a8WRS3jAO16UZfzN7BhaQTGufFm/dzy7zS
jV8DIPwdzKvJe0DumZYOXwsTxM6Y0pnELYkzQEin/QqERiaP+DdtP/kmt8Oc
UeQW/M/Y3ggDE8nSBO3WTta8y6rtGYnGHBTDSCYM7wYdBhOTjiU4BxvPYu4B
PPDt3/wt9gYT4F/A+EIamAyZngOm/27qoblCUOW9ZQY8gK3hgzl/DbTcpfvA
AqOt/hu1vNZK7hrI1oz1hvew2gbrbCtEtbJWyoCB0hcLsGfWsl6BeQoWmku5
YsmLgfnNLKoTHlVofq9C5F7gOdASxjU3OS5ue7ibrYPohgZm3ZRTXzxPgLs4
FAGf9aeafqMLp+1FVr3RZdHraz30Bcto7CXBhdkKdfnA92dWaCXwMv8d+LQW
SK+aNDWzeYw/Y9WN4K84xYY8L6lD+nVHUMenE5O/k6jdrck14R4LP6v4//V4
DVYzUk+MMrc0jNdavtbmZdQt8Vm0D3WVuTkhi1o80V9+a2DRaISN+zZ20Us2
O2fWWlgGmhGmLoLSxQwDh8hzwVse8tJbCmhoCgyQZfgyMRxm7VFLZvtbBOlC
3iPeXFH9PdI0dmPonc/8YhVCWBtjVVGp1yLBbDv4FjVP2Gej8nGS1h2RHF1+
+Ug2RgfN39dMKbzTvLMndQieSXMDxI4IjlPHyvoRVCpNANau3xiMtlApGsNW
MXafatj+0jGchOqcJtJb65xSqZRfXfB0JtdzHlagC/4L9y3k/dpEthQOmqha
XwmltOtuxx8FdaxpPYY/TvuO18v52RajFiAtwFkRB/0ryUXpNqqQsuc5vzm6
h7nxU4u4tNb/HOi5otQBKkf+lYOAypqnP5z3UH8xw4b5d8J/tjsyHBto7nEg
vd2dvR/1rDNPMs6Ibsfj269443KZMXlMh3VfPUtAbWJbQ5LutaW2dX91OL5A
tnowMMUlsYRpqCjH0qOac9Mde8ST9eLwFcYvRbQ9c2k35L8p1FInvWLXIoJQ
G6PJ87HE1PFU1CSUo5k+cqTAy3coAzk33x5xzcwfY2CxWT6fA633P+j4JcvZ
UZg+qkqMBX/t5PipUZHQlK8jJTiTuSN6nHlfZhIyU62Rfv6kXwff+DYxiFdp
twaRvomjMmd//4JTTie0wJ7ffhMOXRLitaHJNxKX1NRMgEwwe2GfRyz7Domk
bnXAXMPGlbigDaykO4m6Xva8/dStJtc1LVoI2c4Q2lCkuA2lnQ38sOoFtsGD
RocAd3xEXCmZ25zbY7YUM7vYtGgtRQS7zY9wKDdchUJBKpkVcxxiF1SvA9la
nZjXV/IanX0NOMtc0YwV5ardCl8zDwz2hUY4PimSohCHGfEAQaXgIL0HYv66
Kjs/zj0T1TKkMQ76Kn/L07QS5hyoBbaQq7K2vPfrtbsyw1xMEo7WPbxniwTl
cGq4Ep2PrCdY5jmT3veufWsq/CmKkGGsfsQLPPZ03yUlChJkWmJVFbw3VPVw
uZq6cSi/w2Vb7mjWUXQpnCPKMZczs1qgJ9wT3PkyGINDR6WOHA8Jp9HCDQmr
5eZitYMNtkYQE3VSVFm0rFap0XuwlNmcv8mKL4KvPDmW26c72aj2bl/bV7Bx
gfn9bst4vEi8WAfRnfOWSQUCeV973xZW+xLBESb9nenEwEgRBRWTXZd5CeD1
x+L5G4+gVVn9l8JqljRVhoGq92EFBBbxqVNWtsm4U+iJtdntaEkhTfLOV/mh
b5JvtC0uepFlC5do2D2ijp0vqEMPtx1vwox+Gn7PBUv8DAAxUFjiRksX1r+X
Ig1w8dSwSdnp2/lUC2xmvxe9KVJf0iXlFXu1OZJ/C/MjEIJITZuQoXb7WnFA
xizSSKLkhCmnXAaZ1/TvPhLb/7a7jaX1zLDe8mv3k24Ld1NbV1jwyjmpDbf5
3IB3pbFqsNpLvxn8blaNohxCSQANqCrXLVwQ3aXNSRS7RKSsEBMZaBF7Ouqd
Fd/cR++disifv5fIJ/iPcCE45SJWcNsE3C4Q0/ot/tN61f0pnWjegQmlsxXG
BWSpfscgxEf+cAlNHPnG8CUxYRLZul9QvGsODUtRU4UPaFqR67+RyBzqRfDM
l/uRfbjYSuh0kdr5ICEiQirKQyJP891klj+AUpIT6INjB9kTu2uh87WZRV+6
gSsqI08MVx28m5jB87qKKsWf0NuDsoGcJXufQY1oprZT6CIKU4Fui4CgqE0O
meEOTg+3VcLkvxuTZOn4dYyjUfWUA/f1MxUxHP7ovuGoMRnZN91t1W4E3jF7
O1D/LutSflWCJihmbVwqqLRB6Fl3cnuGc2r9hE3pqxX3Gx+coPz6+85Vkj8T
X2gCLiTd3lE4/zS6d8QZOsFv4D4+smmdPMdT5J9I/fuSY/k1hPG/LzC4GBb8
WUAlnNZ421NIWao9Qjn9we7xXPOAHqc8yR4sODjmxx2eZAk9nyEac1EuY0Oa
Qfg8AyTXxrNwmbwuH6BE14Pfs5L1b7wjOTvUYfJIprp0/x3OnSQxQEam5A2l
9gqmxkS1B0z0UscPCkIUR8yJRL6CWnsDe4zXp9F147xBTHkCDmNWLPFHf/gc
qwCTGdMdSxZhiNscGTO/UJ2jSn+NMIEPDOR7YNOiaVR5EYpNmqSYxIOd0Sr4
z1/X2cxJ/W6szEstswDxiqpzXUH3FpR5Ab6WrRcPirGEXzgGSpdqZD9fglHl
XOoUV/EwREutdtRgXWT0y0VjnSMsnCgIMrwAID8TXWFJ9n1M7I2bfK8emHhH
ngpqDFlz2MnNQtzM2rMWY73lCRHlD0NnHhTZVyoCvaYotaApHNk8xsfEoPOr
4ShE4uK55z3qqaxDRCM+PV0r7mj+AOBTd1OnPKIYZluUE63aSBo7U+1VK345
VvKYfV+q7nJ9T++55/02jFRdHkoI1XgRun/pR3SL+o4s6HEXxiMCXKaD49Tn
r3VFeotKi5TLPtr+zb5Y4nHoUCg9B1paavKipE1c1RA9o/gdv76I1i6vbzUp
E9ZI4B4keERFJeuh07UZuN2SF8dgUXw4Olk0gy89pyLZBets7Oa53CwMJajh
igaudUf2QPpI8fW4csNGRsXrhw4QhvOM0/YxUeRE/SfWVxHAlPDs2q3KTm48
WDQ6TcONRrjCFbRKnVhWW0E1EM7/mjww5wDV/G9Hvofwda24WhaPtqtOHiRN
SYRfP/B+xWLSOIPWMWRY1IiCHD55h8PLMzwubGBFg5zCiJl3KNlNpfySbcix
jo+SOXdc/OUqBQCnFyr58xKa5EkMFfu+eCeBQuLKdeWjvlIIrZvCrZs5gBTX
hu2BaXOCe4J0TKgZP+wvuESOM+a5uS2V+PxVOQFlZWy0bAsqSggwRahaAMKW
bmQTHsnIHHwUvYAyodr3pw1uMSL+a1pjuNlcOJW9Y7ZOvfPVeXyBm1NWUy4I
lbiAi99tjljZN2Ep2zpaqsCUI0E7nRRQ4U/Iofesw91vnI2lm7nO3mZvTaj3
Rrdh3Rpikjo2g09utImt1K1kICvJvEI5GpDNu3gt6AZo1yZyHgEywqUOfIY5
4oVKDXxs63MojlXsNxr8Ktdx+QwuE7X5KtvmISHRjMVc8QtUDq4YpDGVGO2s
x6KPq82k3NoEfAtbxfgrMYlFZJzScVZpyvAB9OlM+5SsZ5cyPE0mrmuHahW/
tnN1pUn4kJdOhHTTrR/rvd5AtBfzxuGuW4+k64uqfFMkdA5EmHPQnXfswKjY
Lw4X2Cg76rSLaV/y5jU6bk2T0CNuARK/fsMYG7KBYXehLo3/kKwdoMyjSBQS
D3NVbcY4knj+PtSqrK12qzBeFiAnoJhEdUfDFkvVOMUJBWktFXi3bFDgVMiF
R124fGV1zij6R3zCSGbZ0qYuhfsTRFT04uaGk1NA7YxFG+mtBZSNRfpxiomT
SxNe/TKpE6GIn3ZLoNi/nnldKnH179/owMBH5RfYMMJ9s+zJpwImP2dmrTpf
HQ94oK3cANi8orFIznBXfALlnYWdOjrBXfO1t6DsVHYYKkq4fydmiVXMwpcN
eTC9P03611TrJGmDKRYRQnNnEvHH2peCW/MQc0jslQNtAk0mAerY7NF7wtiV
WY4gNR/3IHctitYZf2iSek8CKX5y2siaLMV03mELjyPvSilxGGj7BGE/x8Av
RK9LKChf0EVQ5sSiPMczBNBL5xOK9LhIG3kPil5JalYf1t2ex4ZWu24QO3BA
I/Np6dKyw/xSXueVpu7KvPmv2MotPa4qjh5ZJADUlsxoEq6vlG4VS3Fc16ri
Ri+MqxQeG/CePaCte4FSV5IFAC9uFbd17ArYYSqiO/05b1n0wk8Sie+OOmt+
4r8mR47eVKljDQyX/USCfrmR6KCGlRTn7O+1Rl8vc81SW7TsyNUbBCpowzvx
OOmrk/RfCRk6XgPX/KPtZBFWCZ7wsCMdAgYHdjhnffBGQmpis5GuiOV7fG5G
Z+mxBh8OzJ7i7XZIumlJiP5jN+7Eo4ZK8ORIwUA2qYxEqFTbRbuUC+zhZaHK
ig9AQkCTpMmaYR1wj3ZRQn9Dzc+e82wqBzpKPmjPkoTNTTw83IbDwVD5DkXO
xZATC2LcUC4Jm3yTBjXk6inbYXvK8SZVHknJkp+WbhSgzWr5Tpt3BFYF+sfi
tdbIwqf75Vf/YQ0uEISK6Y01LQBemZLPhnJk19ZmeXhpG3ClAXSH9Qd6dZvw
pi8Hj43fPU5RboVxGoGZ1AVDcSv4nADc9394Laj5oCghzzwN7rwoZr71d1oB
STEZYBXR79ptq2mlmliR5Im/g9Mw8/H7QB9mrN1lGLB1ytBHU+JgouSUBl+i
HbYnAr7ZhpKyUoNBEcDBi5XJCqBBMjQSubbPRbDnYSQmRGjKYMH8WUwqQqQc
AuT+OB6GDF9Pj/8tkZ0B25vizIQmkyM65il8EFlscWapxNsnF0t85opBr/1D
IZ4/rlg9ObLyA4mqGkkXUN/TmJRtdbleMzeDnr54kteHg/YgQuFcF124j60j
h5riNulS5paC22doUOSD6IEBbtE0s+0E47yAHYkcAN0O0iDX6szGh2rR4ArG
BPCDnBE4WWcQ9DzfU1qcXCCVWgVA0iQbeaVBFpR3P5B407irEeeXCmNx1snq
olPyE94oox1jRvsOxoMdXNanLW7N6aYQdVqSBODdBRksQdWr5qMAagu700O0
d6vbcXLsER8zgy15PnbFCe+vdGbYFNTIOjs70wskw0rLACNl3hiaOWLtfsSr
fsxl0VYt8ddsgubibbekMQgYR8X98+hCCS047mcM7Nj9eahSUm39Fl4C3HJ+
OwHCUPs0miq5pV4Hd3R1vv2JP4wAQeglNCGbPNcNcstan+Y6Non29eJfZ43Z
QKOgw8q7Q8Z6I81+ndMh5uFq/6HkgudFlpAyCbcl6pEC9PG5CcVKo/xjbmPc
lB1gqDcafUDj1GEiAWEAZhlIG7XdlxsnDrpUKtau2+9wOblMu/TLPLIyCgyd
jd3wlvahHchXLsA5IP/RAW3wxZ2yAsardM/EcPwBEDxn4kUnoEvEnUo/5tF+
BKg+hjvFV6bx4UBRfSRN5v3KfZv4W0w5TBybZ6PSz2HcciCe4rjPYW9U0+OS
07ZK70SyGA55hGBwHYWu07AuK3FHFnt9QDdAgJzdn7/eZjzdcB/c5SY5wE7G
QbLDZ7d+4LqzlPAChUN+p0MkY+fl6upqXf/He3U9xSyS6j7FVeXMIT5GbYG3
j6qNMkNeiHW1EckxyrPOp2La7SM3SPw9SiEGxKvB1tvAAZeICEVTGY2/Sg/4
eqcvYbQZc4RX6RSoyuS6blKoLLkbt81c/vjoJxdbTVaTbOh1Z8/tOlbJt/r8
x9VOWYZkhtYqCct0L0lJHhSzR/ITCBA8PYOBFRnpkmJ/qZDqgZCuqHJYPFyV
XYQmhz2tWx41F32OZK43020V6OO34aluP54624Y5QvWjMlvq01SdG18MP/bu
AnTcuGoyfaXVozUz7W/Ysfdrqk+5zfcsD2FBvhYdl2MeKnbN1QPzCTDjP717
T0ZwhJGUB/uqWJC5LnZiTygbTM7dP3+1d46p68bASEJurem0SUGoMP479+XS
TtjPAMlVMSzw5ZGlyTKxYUqKhAdRWUW7zIjMpvIWwd9fCCXqR7c5xII3Yx7P
bGUmUEsqpqcuBCDhZ6BOHBWt0akPNxz9sP1larAMEhWLNsHZyNZntP9VoYFU
D7FEjCdd1CRkDNiVy8VwXHs06nlTZd5gX56QhaYX3lhG5vqZ4Ske0ynoFARa
1e1H9O3J65PkGh+HGDB9ZJkZWhKMWB+ZlTbGHLlXO5X0hLgLDYLsKalnDUrU
kXFYulJfqxcL0GIWrvQ+8TFnLlELiY1/Rqnlq7tBhbAJIZ7ilmPfPzRB29LV
qf5iBADRNDJ8btcwZIhwPVdiXjMcs9GFtmZjO2oLPYXb+8fGJdUPKK11zH+u
c3t5Ugp9lQp4HAALsrkAtwx2Wu7oTGia3OgkUFfCObTXi6wdUWS29foqnGJE
c9WlgNFwECWJouV7AwgAE+lldXdvNAJXeXkXqbRKcQLxMlCobdtYkc6G0YrF
lMEeH6ZeAHDyLUD2QXD1ZKgoqNwxqEaMWjleRLf9O8/7o9uGeAf8VvaomP8O
pNsrUqHlx4UP+nCRpMrKi9WmMZnTMGTBBo3kkWsNc6vPRVy1U6VhWTPAs9Vm
ZgGtWw0Yf4Gj+2791yOL0sv3AkRfew2uwn2tAKCCBPupsxvPYERKMyiHDVGD
tgNrpwdPgYF63ygJHT/m+xRdpE5OxUhHViP0bqUcp2CfkQFvZO4fKU+5+fIV
AfH3+sFbcfgMXbKocRlRTTX3HjJ1cwX/5KdZ8HEsCct7n6MbiF+m+0A0hmKM
yeVWWP+aNMN7jNOo1dCvHMFEjWZva4xsEgkyDC3sMao8I1PKzUIx7ASpTq+7
VYE+v8eBZsc41zlQA9NAdiVlanLXZazq1lY2QJHramYuMdsAH2ZwkMkO2O8s
50eXl1dI3pMSfEQGjIgUprI/Gfhy4omMb4JES3Abdr8y9l1I2ywFYvQQ0iI1
HPEH+t5dvm8S5bSs/nmguN9/Bx2AnT6uY6iSMvgz5cT/oCbHziuQ7ktLy1oQ
Dn5fc0CNezgb0DYWnfZD440UwzPmvDJuLrNIfqNmETTjmNiBSMMDsDJ3+Z72
tvLG50YxedPdjvx1cxFY9VvdNNMKN7u7/rXQclnwbRoXA5h7hqrjTBYcFqpL
vqVxIF6YsaoMGwQZjad2TcQcU5qUQn0mgX+Pjw0jzh3hFrZeZF8lgPk1wFjj
lNO7+TaiHj2qWUlGdvWEGIETMxiMPAPvHGyq3ocTAD0xIoA0OY1ulIXffRB+
agy7sbBoh1F+NVnjRJy2ErlET6cwLd1hrz8oiBQE16QumCSZzSjYxcSPp9Rf
ShhqPSqQQfFeknvSoK8CGB1uKKDBmBIGoPMLCbVO4sdUQofwcPKE3iG+ohDB
V1J0fQcR8UlMqy0fviK2DtyUMnzjqH1M+9cUCfDOSaIiuLCUo8SjknZprkuB
2PJK37DVBO/7lKHfO7Xz1N7FrNbmMG1gTjweg9J71aSBraMFK++6het6+fNG
1chyfgP7QJ73d3fe4st6/GbsVmIHaLmZ3gg1CFWvjd2zmHoVB764fSvuCn/J
xsKcts96dQyrdCoa+tUsFFNgqrswWdATaIBq3/bmz0ZzWjl/W/BDx9tX/lz3
krpjPyGbhh2jVNPqQN3Mz7VQjTQQhgxjPFz/PRCGm2vrvYl8fzwjX0rYPwvz
qttWQSbHHRHBNz2VRzsywtNTWz9dpiererfVHHnqqsoQ8JcWvahP570G0aZ5
7ape5BGRci2dPKNTtYfoXH8+f5dkAz4lnY+49DMG4CAAe7wT9Rbs5FLwm6mO
Yf7I5NQBZ9oWFQUZlae/fPzDVHtqio5TqX0GbpobD0+kVBRWosB2Mv1nmjaM
NjWKN+qwGlaKXKrm/12G+1vTtpf127oUVoCLb/HtH1f4WT5musl7BbvYlFHe
fCcPsDS7pGLKRXTB73fc7Xeigz7xnH49olCa0mA/LCZLaPpMsZ0nf4nVfXFm
mNGQFxTNnDOFSK+RQqKNN5GxMAvb90s88RT7LGVkXMuS+1tw7U23eqTA0LiX
3pLeRjh7YW4aC5iORSAm3fzwFSLzLYjtTu0aCmc/XZOZd3f8cfc5KSdDYLkA
HcVd65+nD9IPaNsm2XVZHdcUYj0psAyJRojRCSWE5UqxgXi602rTLwuTpiIy
wBwa3ZfFL/k72SwLXUTcD2yBylkNTkfkNzOpV6eU1K6v2SPPEUzN65MKfIZO
Px0qrgXWp9cLgZpUJNdgxdynNrs+MoPsLL5EiRmd/dOjng4K6Cmc63jqKdmy
8CZGxQjl745O5blvJR9eSKZbOnVawDk3zsz9kq65mkRx0mX45vJGGvpnxqlt
ltfMQKuPkXUXFlpqujOHI7JiFlTAFPL5tK0dMN0NJk9DHOJ6dlYAnl1vAUwx
97IZZpZ53hY7N2dx1EC2Mpg67V6bejcmWDSeEtUtnQgT/S0AgfFMPt9nJWzK
mXsqpUBdyeinjmtHUFpy95v8kDSF6f3zemU3DRowOxK8RZSxvPQbL/AJ3dfX
mwaJ4jTmV2NeDAoyFbWKgfac/6kGDJUZDyQEGzSx9/DMmzSKsIi2hVBSoVLY
J/WvN8R8qfjASlLZd2uesCQUv2Q25y8ObOGzCjvXlVayynq0SWd/ryc6MXRw
NGeZ5js8kOhMEudeV4A8ceFR35HMZDMvipKrAL74BZe+V8wYQkFKmZ9biO3C
XSvTw3LFlO6ppEFnNRI4j1MV3gokFcRzo5EGfOamcrGxMe0b0PcN/5hmy1oF
IhSJV3pTfDwVR/szinamERWy3HvXGSkLHC4LwGthp9QHaQqWcbilyTObkvy2
2viQUpbzAY1R0oywX5ED0NgSj4YerwVGjizzfefPDff5KwdZlUqq3DjRz6WU
JAKMCcVbaqdyBkWJ1gNh2LImWXrhBu2yVWj5Q3ZwKSPv4o+eT1q+l4bONxST
aoxZAPMeP82HkDBWtmlObxr5xhdfKgCj2BgDmn7zg42t1ZWrQ6Yr4dmxYCAn
kfBAlbvQy1TP+jQNMiPMdR1fjKikiN/RireZI2fzJAR8nqUkHb+IBvuCceBb
uR+OyDUdz5X6UnjTdG38TnTj6empX9uoqH3y3aeDcAWxl17ZI6x/Zt9QQ8Q5
Xmp3o8Vy4BFYEmvXROMFaxb+FmVZaTzFc+afO3RLVbsixBzVgPolR49fQM/9
IM9ej4B4ZL2QhPYaeY7RsAdikNW9f0U9CECroztuAlFOA1xTtlZ/AeowWhwC
aI9UCBgA04cjn7M/UUxvafeWiM+RQA8PBUAObr6oJGY/DnhvUfabN8CYH0h5
Z8JGYxx47yg4vHgc5jGLgp+TLUZaFVav8PZYOEXyTfh5ZL2cafvjZZHLjX55
2gtrOdyDUvypQ+acJFbiM3hpDzP7aKeEH3OByMyCyc7Yk0DU83F00HN3jXqO
ilwN/borvgfBQtxichHWX1MnDenvNb2jMZ92S2OzSJvUUuYbwdfsyOHW5qKT
WqzlZZ4pex3MSngYrpmAjLlVkKNlib62Tqo9aHVOR2UL9CYmrgmpBiKw5qhc
ZEHinMDeV3BoFfhavkjKNvfvq4OoJG1iplFaMvu+n0+wpwxWgXHW+Rfqs/w5
et4wHOrrlKzRmEAi8PcCx8HkQ2uEmmudSPwTjTDDrdPItyQxHPOlCYqy0CCf
d/f15M9X/0d/6OG9AlQOwNYzEVoPDvyhqN3Oee+a/Gthdoni1CGnp7iI+gE6
Zt4xeL0z196unnA8aDP3dyfVgKUeVrwBei5xxmQ9Hdve07R6IUBz5sYGiuT+
JAWe2kCRBP5KlGYWTqSRACEENOJltaMF5W0OZ/pehK4Ez/szv61XVKplL+7c
+bHLViRimi+ZuGFWtlQlOiuG8ScntGmJ9ZZcrDgtAqdVA+KaWesHSHzF81Pp
3Mw8tsZW64ePX5IdyT+6BW8JDY7kRQ71e9T9DFn+PikoCp4ZrFSZUuiGo/c0
ag87P0wYcVyKEreFFz05A28JTXwX4CoxK/FPYSAEeeG2jv1hU445qDI+znrc
no4icx3PhLO8xGZjMWIJQsy/bTFIhJiGShBKdCpBWGmmh4PAF+v9K5gpjI1M
pSXX+chHC7b2Bi5U6eCJxQkMYfYjyen6CQxeUSJ209ZzNA0Dae1SgMjMfeXK
0b1y5uwppXVXuA7GpD43J0dozhRLH8GwFDG7zNnXp+MMZCeGJc+/munnIL1/
K24C3eSYi8EJCvHe3EHZcurM30sPi0ZUq46+xYjER6WXENdPbAnbdrErl8fb
UHyy3MekwXhKKKSZwaY7aMFd+DukmkWri483YYOwu/2nK23k49mxGf3g/tn5
vScKNzY7Ou3OCv69I/CFH9E6nhJ2wQJ6WPKpf/24bSDyRnXo9HiSfPYE+ph9
m6//GvaBAAYgEOn3nIgT5Nh50OU58aoPeNMimQgZ+GNdbacgDS69GF06zR5J
GI8+1HF4eFhVoE5yBQt2lDdPvACkJmlV7h31dfQYfWnOOPigTz5rqMj/kSmK
GDS1sX1WaK9OmIdoVf4ThEXQVslUvPpCDY6zrUBw0a2VuM8xMFT8DvhNL/1j
sdobnwAh5a1Kpj31ro6IEyLqLPgiFp73j0TuV0Ckt3Iu9us1157s3JsyX+D0
tXQ5ANEp+dN/a4Fh7SKNPs9JOlIieKb9HLXre7+TewBE1M2yrY9l6gqvZjwf
5Db38hQ9etD1L35LeP3JMM+3OAT3KpvPU0jgPGfPM5b1VWjnIBrQA3AG3Sue
5VIZ+QZf1KKDZtANAFNB+VtAauIz4kTe5mTiUgzl4qEwbM0T8kEUF37mGjHD
CSjj1pcMLd96YI4+VA2kQBCi9dlidKxZ9x6S8GolTifTrUEPTYG63OksiBR3
6VmjO1wQwD33JRI3vkEGEHLIGYaXFaUX/VWdslh8NX1wNUSRU/BftY3Y25Mk
MtI7R5TUgBIU53/8mxziGPQNzmcGiLcg2UjrrJ09Y4dBebSzJsqoU8o4y7qy
sA86UsnksiQj5G/ZIWKyIOdt7CowFRFaaueTWdJ0hLzdg5Eyy1hgxS+kIJi/
4Y2N//XvDPYvs6vmmfcTb8s+7GQrj35Mt8+4ADDqmUgQOvq0N+dFl/UEOClk
T7KRbYBw0OOL5AtmPuuJ1mbsWBX8OJepPYrokFgINY/hJpbV1INNSzAbaysu
FC94wpKwMb8Bvj/jVmeeSaiQnxpc9YiuqWw/gdkdSuF8kshrAvDNvEOyhvj7
1mzPV3NiB0U3x12iS18CFBTVmXq9YjMkrzlPpPvqj7amAa/JMK2U0XgsLkdg
oUyv19T+kJyOhw1e2arPMooEllz1xD+xv3aSBsZRppNsiffv1sxolyOJXcuL
LdyfO5Y1lCtp0d2U4K9u57UhS/8YGvUX9/6Id5akLaCxT4k1p5nieh596luw
9NcYoag8B3gjaGd4YhHg40+8kAMDlCEwfDmwiC7s6mJhAiIXvRZel50EX2yj
WO1Rwk+IKAPc2lLpV3MPAV5mcZGZVSMuB2R/MxdHv5i8WnIdGxY0X91AZoGk
884naAPaWWeL6BAikkcrFoKMcF6Jiy7fVP02moyuJIELYJfMU8UtzyEjm/mn
lBdBOoCH0+4nJQ3WMFkPWvhIBInsxYb31g5RTTEC1ApBlBtu/VPPhv3wuDUb
ggkauMFUTbcTRm54L0EQ9JoDtIhnbbFMyE6hcxrOndkT3bzlJM2XknP4/Qup
0MKpUQGHtRASifPl5xJpE1AcOZrySBg5e0m6NRppqax33/t/QLRlRWHCkpIp
ndVZ2vxX8bdY9KtrsPOJRC69xSsx5IDq6+bHytxfxmOmmWh64BauTY16/ty2
LwCLj+0l5qCGYIXgaQjPlU8e0aEbt6+F7Gdg5YkhadEnG5oGP0nCaVBOb8F4
jyyz6HbOWDf6ANazDdiRxSiLU4+Zx5VkBoyhqLhI59Uf2Luik+/RyYcVAo4N
sguYSQ7iU51zxs2Qclf/9gL0YMQkRclWurLaRcUQLH8ghxIaNACHxdBQ6/QS
lmJAElJsnf0lMSpuOlcXzzsDEQoTynOa1eT8rifz1FUKW9UH3gGFoXvYgped
woyYyclmwQDLJVeqdi2I4PtEzTmO8xckiAlC8XUqFcmxWaTvJP03UmYb2ttb
A2v8tYM57GmzV6dINFwfQa0sFZSI8knG+KssL2SPsivVriPI3iZThPfHIkF0
C8usr3U+MeB5rirpEdjIas7BcSh/gItk9aya5l/aizjpiyPNxPWS/IuU7oYB
zYWAZA8Ta6dcEcNgYsIgVoaFHEt+NliH+Sls/OABTSRaluFgyOrjsu+FiAdp
SNOLT3wjnOAdVcbLfV6ZLF/i7Pqs92uVq1E9kjCYjm31fzfBDp74xYhBBhNm
TcwwzWwkgitdakNPrUWbJtpWYw4DoQWs45qP+szz4G5oIdgXfApT5SJT+xaW
MmG2982guVGXEIydc0+gwarBvjqElxFhGEcexdysh3yHXabiWdSxtluPZk6C
Az4S6jDQfNcNzWHVS/QOg0PGyFoaZGkMFbslXrsdUTYlAsSzUz9AktmCgVe/
dFGOht9sKeMvDFN9D7GBCTJoHZV+NpoBvdyzzdEYaH6SSYh3nNrA0XQK4Pn2
xOJwz4K9DMQL88a0eWnlzBgn7FleBS6sWEHR7M4zjRVKw5X9dRB4WRWXWapN
+tUsvTB6F3JjzZDqM+RJVrEXLyMysKTJU/AtnLKQvqBuaFU1L+HomRZQwUOq
HESoJaE4bCdVGVRywTGbbLml/wlpqJ9FNRsX4tzsfEj3y1TVPsiUaI1lvshQ
SJYW6bO80AOOI4LtXqAQj8vMx/FIpn9BR9mw3O1FVoPw4rnDzwxQ3OnfkZSK
D2JEtNPH5Lo7FQTWbNy6vfoCpvvxvMJBmEF4pSkJSLmfx3QF9HvkWJNvrH/C
NI0CPapnue/mg7yzsBU4uAgVBsC/98bHW+Rs1NXA94nrX4wiNrNPWi0QMBSY
QkTCbE+7UhmGwqcAEE+SJBpYROALDZ3Ah5pf+mrm+f9xq4EYpzbZzDG8oBx6
YR57a9Wvfy7vf/iOwGL9krJvZLGVD9sV7xV63tobH8qNUdaVnjPVOpsuA47S
mPO8HRvjZmhnPdFfF+/jD/qyrhrH9YgzUerg3aSOOijMwbiFOqSIdynCCFHr
DRSuTU02va4CaDTQIYWiZmZC6xJ110xil3n3qGBwA7MBrZJU2GXYoml6KiyE
0ByPnSRs1iQW27x8KjGpzNx4DFL0XIykEnmCt2UczqeLWEQHvKg/KCEz8Xy8
0w3tbTznHMBY2FGpjOiN65tsCUOK7z2Zr/2sN7DSIYw0tMynIaBGPvfaGJR+
YTOL05Z+RavchKpFUIqyf/sxSHkrNHHfYDsvs1u/b2CBcKFZ4nk42Qnpcw3S
q4gWn9GxQdpsJ57l5jR5uAiO1T8xyqCoj9daSGtGjUWEL0nZx10o7DoNBlBO
OpejdzYYhIlg5ja3AehBI1aat+lJoQ7/o07wnOo6jXDWVLRacY0akmj7HEsH
LAKVn08EDQLKaZOwxFz/CO4hsaUzBTw5DEBuj2Jl99chtgiHV8mSHDCTSH1i
fvajv/SOqF62XUEJDoGUl+R/p8xHPExeQDpSRP5dZ7WT0lLFv0ZvcS71zInm
/TyBsRR9EhMY/JFoGfCNWNPffGav/Es/uPrr9vCXqF/3WC4wHUbTQmIxZ/s2
FXmwhcdtA91a0R7v1UIi25yldDGT8HuaQyXEMHz0w8MliApEYfoDno6P3lzM
GgXG6i1GnmFG+/mV02Ced1V8OQv/kM6Ejmcom3bi/oWoonyRXsv7Fw2sBalv
PO4N4hzi2hPcATpd74DSgOV5b5dr2a3bfsVnWHcQwIYAf2/PsS5qV1mM/30h
CzrR/yk+Mm+USwGSviWdVB3v4/0atgkast07NUSI8et+48WlKPptT6yUyjQ2
9ygKjXUnw2xzQvfJWg4GOJhZ0hIm+v26JNOMhOy9nI04Z60jgZtU7QWU/wvC
W9HODgstZ0dBKl2SkV+iXvRRwXh5dwfDi5oov24WqWJVhY3yZLU4FcKh3Dcn
wA/Rq+OGr5xwRgQ8nPkC4UF/SuiVxZuaZ9VvfRxEciy78HlRFIkn+JZyCB9m
JJmoj6m6nHUqurS36kNiDVSVLAiipaDYkG9SsvZ4V0jX/L/nEnxhWvLP+Y7G
a896J8uATkH0tCvZ6G02kMcIzhHccZbt+sPHcytsjPtWq3vNNc3A+KCAhe5q
hSo+Icr/nbsYXDmvoQZ1f3TOFVdfhQVtfT3c7lUG7iCSD2StaD2fQ38bSAJA
WteTnuiuJCa3dqshD3hMTqD0Kwv5Fw2CBN4hk5vQMlvJvPSPAGBWXzRi7v07
Gzec4HUciw7jbtuHW/iRzFET52/iRfZRpqqzJ7WDDbmZTUGfG7gx3L/oZPz5
aYucxKBkuqKvFTwr2iFZfrSWCxW2jyXh4EpHoz0IQa8VH3e08l3Xfb7OHWTO
TUyrjE8/1Nx3GK3+5iNen7npJnyCYsQmVgFnkwp4iNYpEB4IN6vTQSZofOfF
Y9cKrLG6y1E6FIzQw7pb1ocQcciwJv4U4mepY/U+ALxUZ+wJJ+JiV/q91w++
m5d6haZS0RyMaijFxTqNXQEm1kg5RRIByiWO5UxnGWG/1EQ7w9rCaHUp25jl
o2Lo0EealdE8GjuKxtqxAXcAD8evpFmpAlqHSlezZaC1uRJL/05tNMBaN0A6
LvVe9n+DL3H63a55ot/W0rBfdGF1VLHbLpZRvdBCKQSAyMuDp7mby3eEVAra
tYoRTK6tCrv1cVCayGz6/YjasOWgl/gEmkcCQnDyx3EVwImjFWunc+rtuqui
I4qhXLmKcgX/nYlips09+ZR2fnE1dkJTO4b9kdc3s1g4ztDp8/Whcvh9cAhl
8qoOfJ2h79DcQr2WGgCCxcSJzBxqOuKaFeN3dYQz+dJtNm5C7ieUtfTvo5MD
xbKrgnp1eVm/zFhXSnBa+Sr1mfGQRtXKTtYajCYukOhsqh1kzagLpFtsi0RM
JpODAuNwOrZOD9T0d/hOdSvMdqs3iO6bVBsB1bk2XBfHLdA517nYlj2p1VaI
nY9kqYd91BwaWwUWFfh+N9bnbgbRRAicFmLXjUUJNEIrgsxWpMFz76Xsw6Ic
rUzouppfYb1GvPANf6Q339uBiYjucJxqmxEEtajZIymfG0k5UpDnPh461XIA
VS9B3xe+GoHOlqsYkEh8caVdg/uHTmzBCDZrIiN7gsLWZUAr2A1lvCrVGz15
Da+L8t9zsWnoQBvq2Rffeb96uMTovMRHxp690LteQ+TDxlgx+FfdN927lbig
TBN8mx6BP6ciseaBAj47tQFi+UOyWnlIbp9ZMCzYnUb/qJDYvMbpVpiwNZ9Z
U/s5MeisWtR3lJl3nVt0vPXWppIXq2MNK29icV6JqqQqnzc9aPiqhRSAJlZq
zbSgftKp9V6+cj0Zuh8E8i8VIMTJoIBtektjKMhlSPU2jRc3hzbQzEgdjISf
0mNc7A5eTqDGS0wscy6DPRTGKrgKqmsHsYS2iWStSHfDCOEqWy+7F1PY7Ja4
PL1Lk45v5pe1LM9s4KBmkwHOQQbO1a1RDTvcqt3S1xOzPXvemPdm8ocResc/
GQ6n9HDkQsAJuMNX9wMBb/iBme3qOwNWTSnVbHv97nWfsE7Fki1JnLD3+Rg+
lL8V+Jkndg3ow1OX9IN14PDjoXNysAZCDJcoDLWPLKLYahJNeZTwKHMIOtrf
S/F2LUcSfNcUqTd9/SEuC3QtgIhH/nTfux+rTH4vuntscyPX9FLuPjxCZUGm
KycmROzV/9ODGbeaQ4ItgqVyXQi2gyvc4pwb02WOG/1WygmIxYtjmNuXn6C2
miQySo7R53z+FaNBS83EsIHfcQK6uhrzcc5tHlu7iDWdPAqV8KSijVbj0LQj
uYvzBTi6CY1Mo1xSWkTJw5qt4y+nsUgp3486QG4r9C9//LZk9Ps6+MsCKyR3
MnEnOoqFiuRwrclFsHO/iWut0aaxMpP5I7AlDaiaSx5mH0MeteF/56JSObTt
HqSvqBHw/2QGmOo09NSz9uAYSQ1lTcdbfPgEU7YcJ9Yas4Ac5v+GcmMkIPA5
D4k78Tr0/1vTYHcm1Sa2wFL0EBwyXnAA6lgyZlgDousi0AFbwnOPFGcDnBGO
3fwL3vsXj3g3HFIlbl0F2SrL3zV5mjB+A1I3pW+kFJVWuq3SKhQ+w8BRGtZx
Rgap39d749S/inFNhzAOKp90LNv+zKsmLDk/THkTO9jgic73CHl/bxEFkNZV
vuhnZBK7eYQGFTVxfkwOGw4aZGgUH8TOT+ivC5pKW7oikrXZcLqTmOYm3Lhg
p6Zzn6UVPVx+Y11MXYQ1Mw7Y+mIj6qD9Mt13lX+Dm+kzilaDp3sRK5oI/Hbt
eLPwaBW123VB81zoDV9Ceniib2mIsiNBAJrkSvYUOn2c6bS5ZXo9QhTDX1sz
90DmZ828RzYeIa3jHEzdCKljpXQ5bX1784rG4eMR+HqjsLLFEXp7LzEbZAo9
EtevH8Uhs1zoowJhiXzg8uPQ0Dztzti2LD40maJYdRVO8GOU3Rjfs6aegVtJ
sJ5wz3ZKoCVaJeLgY3aLgfeZSixVtNqUd01ilFGeJURHOoiRdydjG3UsB2uA
2MPxjkWR289guN28UtRyWbqvuUO3rY5/JwIYL107kdINSYpt4jY/LjqC+Jcq
HQYfHyYdKq5YRq3u5CJ2NmepHQMHWdHMpQR7hbPIC/r5Bq0AvxyAbb3Ie701
KkhpUR0hcfujAOBoxIkiXWjA6nYJBEq/PoWR8q5yCdZ6vqt964jLMveV9nDm
8rl/QsBK/l5PSdcLwXqv5hPQwtmp6kNDE0Hm2D3B8olkP+qxjol1slprBCp6
MUxg3bYZ8yKgP3qYkEr07Jx0NFmR+Is2zQvotwC3QQzaNs+Zq+8C3W+WvkL0
kkqhMNzuQn0ThMV292nyBUf3qsaEersAy7Ac+ddLt5h815LuGTsfqtjog8zu
Ae7vdfSeWs4BxVRnjy5cbRx829knEtox75k+hyqMiZIGc28pAd9mSJQ+vA5z
k2eXxEHx5mROckAy1s9dgEp13BEbpfPtPRLvD8TW9rEXkNpMQgkP6JX0eiqa
zhcomXy5QIN/PkQ17PwdLkh4+VU0CimDPPAS0SOLC/xtYDuaMnDA6c2bkvZH
9QhaLSxEqxk5FnieTAG2Lg9fRquZ1j/Xe1ZIGaVic8nEOUdWA+vBflwnj42S
C1Q0/PWbd6MY20e+q/MjIIaVS30fCeLXo6tVPr/jQw3zQGu2wK4mGVmjk63P
ibHmtwkPSXqthpWLrEozUSjNYQfpe9RQGQmOueB33Itg+qeJADvKZH8/cup2
vZg605vYphuMLk96yuOYDy5oG5iYakU2/UUVJk0HTym7Kp4XgDfE1GIcyAyz
rT29qq1d3ioi2n+/PFreEhLzuYJIhIsot7gptFul+nlkHuTwBUkSMHmmFeIE
VQMaGu3DVwkf+bz1VgQoBQTiinrlyKDoTiqYzgEHJHkdl7xVS3h+p3p6Ndus
WwnT+m7JBKBVduWOK38WF/isKZJlrZTWA05QzDBNK0xs+T/HdhEBfQavHlQs
mazABQIcI5zBjjS2u94aT+w4dFoR43ttoZpQpw4ZS9wOU+Z7P5Fq6GEQ+HCY
yt5jHYWjPc98628tDhkwaC9s2Yz2Wrr8Xusx9VRvaphO2p4KUJfW964zLtpz
mh4MImPgN2Q0BBk7eyXhE1xEucIdDYCw+wCl6NyKZoIbJY0kj480+Iskn5R2
+MUv+8qKJ+5KDwvd9ateu2FGNRxLpys1snpUBdbu4NYFnqOj1brFML+Yvb70
QQkT+sNJxH3nXWFpSVi2718isv37glCG0XzmoOiLNm4iXCyPNySdnGfNEc1C
8gXWPxpmyUK8Hollcm8k2uoDlj4G+E+O3OqXlv7tw7ljwc7dpY3uHzEcoV89
K9Nq/lkbe4fNfkhBF662ZDNUsQ3Tei43MQ18VlXqrgdGgZE9CJ7kclJda1cb
zjoT/SC7aBXRl/qGvNUDVYGgrXgiAiaCXTXR9Ph7v+KrIeFo9vtD0kfOzcgL
q9ddszwhnwcc+7+bvE2uZtLOVD5nwUGmDSq5eTV1jKjzeCpk48l4Jw1PyEFR
P/KrtHxTw6I9YTJoj5+bVUhwkYCA3nokuwRt081c8aVmFe8Y7BqUODGLoC2X
Aw+A3ECFmRDEtI3YLTKT+0FU+IdXtiKpF6Qo1nEQCel4aZbr69eh0jbM8ahv
/L5rRxBZ8cGpflv0HJzmvMs54l9wGpfRbRrMXh/hkpCcZBZxfyjFa92i8/jq
aR8/zu0WYZSzQ+kFhkrWYxzOdQPyHI/s/t07i8OgYYgqmsgMZl357X1U6thE
h6SBg2Lq+RlCY3oXBq8TKLG0pv8gDMyCA5flKLCnOysyy2v3HovUmjEM4hOY
KF8uGvFc/+usVy8indbIYo9+a+bKQeaf9m7HlESGaZoMzPonFoHMkQF+ojP0
CyzSKXyzNSxBlvgOaqMO9ibTIylwH7VVIpaPG5rYzQ6VnsQPs/ZU18EPL1mm
L+y0N1mTKE3w7DSeiGVPZR7pFunaUyNsis2moXKG1UkxB5fS96/gBWfwmG+g
JNKeEs/cJKXp5Fuq+M6A/a1dywVQtL9I+yTc4mEVk7+XKonYinIdtdrqLJ4Z
5osINbpPLaCvGo80h1BLehlA9j+kWUTIk3yuum44Mc0xkg5QczXaeQb5VHEr
yVOZSh02rAJwRIRkRKv1fjn2fyhxkMuETzhbmXNZyBuO/Mpkl0FSYC56v4Aa
P1Y0ckkKKv4jGbw5WUVjgsQJqZLkmLtNbc9RBhRP7aZOEG+ItmJnDLSz4f/H
e+2FvbaDzO+GLYP72YUPrj2DNt9piPXHWr6hEAYk8nKYWP9AZQq6KZmDqgQI
gGl2RwM7XPXVniyF0PowvwYf2W/TgvISZXWRUrckW3e6RD1BkQB9XbfK6bkt
P7xNHAmyD60jKa/9jcslhli/7V5cKGpMdav9hRMtIh10ZIZy1aPfICTBJgob
8S0A+1X+19/JZfmJmUVhKr/jx1hgSdgW+kb20lum6USKTv+FZhgbiWQEgvGd
nMyRlLnM8y68AD6b4MPl1tvlYvW/+iIS4DRaq6qbvuAt4C5VhiOYxGBIP0gB
HOu6ywXaa5kC3/5COqJXaLxMY96C2+G4e7TkKbR1EG5+gdI11rGYD7nb3E4D
DdhFW8QSoMvOusTxyEPvy2MpNrgKs66REI+lwnI+OnX3mCFOwm3looMISK7V
C/PjKHa1PK4srk1vjo6q7lZenroyO0ETkSHxpmYDRPirA6njww+d0CJZGyRo
PhjLIydyH/bIZa8PUyIocKomv85qCVewV4F5OUwboEg8rBEKfKNYJIq60SKP
yAIOK/94QG+9gZhoOAwgJ5ZXZzsy5cPd7xJaMPUDf8kBqNsU+fF7Os1lImWs
MBrHUebq1MRHO+anSPXv2QAg7sSB7zhmebzW/4hxR8Lxi+fwzbmYSSpP2xse
5M6P38vPhc3FYVdfWiDsyY3kH4jfHaxDCxfHe8aoi5ggGTa7TX2aZQITk+Cl
Um5dAKVQxbHT0Eb72atfhhUrievR/p/3UPFhY670gKtxjpRG3yQtt9fIP8VF
P7UPTQ7t3tG6UPVx8EgGvl/KWoSILf+h/xedMk54SM0u296DbcjnPYWjmRlx
zaeYofD0j7LYC8EFaeGlQp4y0OilKVy/RZO2ZuKK5v6syF0OodE6uqXccEbS
0JHbOc+dkP3q9e2gJMX16Mi1Mbbabcc3knHmtm1yLIt2dxKCXlfEKsIn5f5f
jBUj43CmOYIuCu15L92+VnkpA8kq/HD9oVSL4ajXtFL/8HLRDV5wIlH84Elv
xm2/DxO735lZoh3Ff5lqM8p9OSzewOBnHgK4Jf+61hO7g/eVxHnWtXacVWhh
bxjgs6IZ86V3UHU4KwUM8Bw+pZA/QzfOqe2OILTrU1Pg6g1smXpFYprE2HqT
QsDowBFqzbrTFkjYIvko8xUa8HZbX/D1DVfPRjRnSCmVZUfvAwo+8tf1rEaK
McHszb+MEDXu0OstvMGQhv7bPubRjJOybrKn/Trm1dt6xi40v+q92LmgA23R
f1RLnzc86+YFaRYlUwNyiXy2nA+zcyTG0gHLyxrdPlmqwMzRYCltlLkk0gMv
A9k5ADgV6IWEVQqRsflhkvKBpjB8SotSvHm5YttH4CybI8QU7L3VQrOl/5Ms
6QEMZLdXFKjEs5Eiitca1gmPWdqnV0gazfplE6JXvbFjnt7yaLdhMJ+WnX5G
YmYoeLoU/UfjxSAsMliPxqMBxOBOzPy+UI14va7eIWExYD6sqi3xBVvEHtvV
TbJrBbtQWHZWhCoyZm3h812WTxxF0Rnbw3Hfc39OJICC6s9jBO3RceQ5jo+2
WaICwj0GFPcM8RRQlNEj3kwC+4aAe2qi3RfcT5fX6kzYRg7X7KQVj7k3Uj70
z4zFQ4Kki+8SUXuaNashyFOMCJM9Clb/HbiidHPjLPlDPhiGGLjrqt1uS1Vt
HX/oDAQJUGp3iiKXgNWoDBD1as1Hn2jhVvTc+9bEW6W0tgR7KyuqB76aK1tX
EF8+RK4kw/PEjyLKc4zSV8pft2WbIP3V6tq4z0V9/hWJRNVm+OFpC74ml/Sf
YrYecezSPxkUKA4J1l0l14tqOND349zOPHXvXnvYbAzBcdXJiN2gUCHq1eIx
sI7H13b26Q85L/26WlL/SUSBMapg5uzwizMukIgqlQiC3juxTzmvIjRfYzjS
vJJQdqtYRNkf2A4lyI+0B7yQOORDaE6tpN+j8bFsB4c+eFb5pUa9ZsnhzZoM
/NqYQtf8r3W1fs4vOVgUipOBYUD/eBatbLqjZKKDo2brraua8RC0/hIs5NNe
jBmIYB8K0JiKdmm1r5NX9qiFqTglcH/uVUskTVXCIO7/QlqYMAHLQSOYP74I
PGGIVzO/06RFP2y7L94dvw96klVUbtAuAMhVCBJxhDDP73eJSJLQWL1fD7+M
cPYeXEdgNcQe3d0DgcCmSIcQfdLUeLdTKx5/CwNFYTAq9GgUWuKqCKpNbR3w
Jg9+xPTNynoHNvdC2s+iT1tJgah5Sfn7gyghBDUcNt/hCUZagEJ+w+OfKuKZ
OkLaTeHU5EsYr8T1rW87/6Xg9ADktKr/aVg8NOM0u5Bby8C9PYIY6tJqMIyB
l3NoE4qBTEzapxoqLg315FXu2vnyRWKEhqxgLsk15GQDtxXe37ujhpznJfyU
PiLusSJ875PwrzZ6C+0j0TaNJVrsNancT2dyx9gBdnwO3IOtI4BC006QRbFs
K6POf2spZ/RJ4HUon4xxkCkEjbVUpvP+3kF35LyWAI9cO2ewhdpTpgfoPf1g
IWibiCAHEKctrDCB/G8Hp75LIDqlwt6/zLeRVg+cKzkx/XoAk3KHBT/ZloWP
8KEzFXFfImyurpGnO8xr9YCLFv1kK7Q2vIvAuAzM92llRqucqXIlFhz7/8g+
yLaw/KIuYnZ3HizKgCAeCS5arrVFbXbGQWkuEo0HK0iHO/lIB8MsLnYkgyZw
Jy6wX6HJ0x6HZUrxDNZFl2o/DJI1WAjxFn6Sb2zidd1YnK2KSEH4BN74VBB9
Z0yr1Amj0ernXaW5zrcSKfp9HL8Om6B/Jx2aaoAoGJdNjx134NWFPh/+m8Hk
tDeCJo/1k8AIO56G7tSt858DsYxYVbqjYwvXR5ddRxdoJSdNttblc5HMSAMA
sL6SBGXlhmwEYv7W9zti5RWIhe50DhqSgxoDzlVEyugIsc4afn4O0+Jf6HcA
AqAEvew90qPyR3wB3UahF9NDcbxl4Z/c0zUtPzsuP7nFa4sETYWpv4wBP2zX
wqkPGkPxpVt+2ZE4IWCGqW99S0VFjXTgUWa/7zbxPIQoFEHeTOtNEMBfzNGe
YA7lXSibBGgpZHRRcv/KZI6hyHcjVdbp6IukT0geu7GtpCvl5r6mHBicOdlH
O1Xjzx9ysyyv92xUj7CEawLxqZnCMqcbykCZJqfYZdw4EsZXSalQqmlXgEf4
0dD54ZMzuYowfxHppkZqchtTfh3uFFCZXFBwOhl2yNlLdgWidaMn5WSd4Nb0
RAVjG/NP8kcvgt8mMFSlJz0AGXb1b6da8Jjy9/L0geeAvCG5NpzNbfZxZnfN
kpBnuvXvVHHUOPgfwfFJrH1x+3Sqs9W6FruL06kpvYtdUWtn8XVVy1dWkRXh
yylaSWsiKnaCxayYjOYmR1BYrZGBN30R5lYenrXEgxwkWloWImwUtkzEU9iq
yuJnlASGYjXS7mSFGb0MfpcyWMEFVt2jXvHQi4OJVFRobUf0yhXG2VVxNBqj
20ybNp/PWE93doMQ76Y0FwZtU8lWDXqhpHurmygfVwp/EjVo5VF5fq3IFV1N
CwFEDoPZnH9PlPeSCCM9qGJ3IZ+JRflKAvLPP/TtOPyHjYqy5WgAIgRxcxA8
+tSzHyk/WS5K8eyhcXPHKcHqwW+lbugQT8jA30g5IbnOyaM0f7xgBmGmDv9A
1nmUwzi4LaLOeZB4mXtlRWE+75zJnu+2OVClquj6TEd1XR2wxARXhLgqtJu2
6RzRyACVnOM1L2ZAtUWmgTd5kJwFl2VPhIeG5q0ZdaQ1zZEc+daAKLb4+qJa
spHuqbtI0bNAp5w4AfAet8suNBGjSSiFydIpoZZRp59cv4Xv1PGhzes5k8VI
pLBNWvj4l+C25+xE3JTLw2LaPK5OMOgSvVsJKIsuDp7sQXyNpCZUob3pWS0Y
xSvOd3bTdyA0BATSN9KqRfWcVDFnJA4ieRmckF0Wc6mCyb5s3pjdoYWtBrdg
Xi2GNdPHEuEUzy4f8avUM3P9NPEFLXU4WDiJbjhgdGWXMUviPiht31chyCtn
8485pzVSWZm/6uDFCJKUZ3pz1XFoXYpTv8PfUn/+VxbQ8X8N7/PsUyuYd0zC
2FIy+JBJo5i80CMfUUas+wfPdgxEKXrGi/UdU4yZrVahCHdaONl2+lfnZdP4
7z1WzWYa96+7XkiOJWvg22fG4ysenX4nJh1AMOXNAF5K24BnxtI66WIfj40S
16s2m8S73Ss+hyXvLpBfVwIXgo0KW/v54fAZcszzVnoLQttHD90w7Ct5QqHa
06ItTZfsYcki08t475Lu5YP7iOKMsCxqVZVSBIfpC3KCj0l8Z7VldgUQH78B
thfUkWgtspjXGMifeynvQydzKsb3K9/zW4fxfBiDxeTSWYa2xifHucS4GgH8
f9EosdhuObhJzOYEiipNQMAQTDwBOFx9QlAj/kyq2Le8cq3fZNNPuf+HZ97d
t8LZop21oOWsvVfnKfbgOmwCiblJn7CV/ENXqM5WroSx4OIcqzCC0uLMeUb0
kEMcq/EOtPYycB7wDO0FkiRJi5DAMxV6F2k/hzmXgId5Yj6S0I9pEmqne4KK
lnt3HyvIpjQauDMJzaPzs+87a8URj79pYmDygGbX5RRR8cmmrxG29mPHH4tV
DitPrAmFtXm/nrcjELh7GHUxf8BusLSpAwgSFO1LWVbNpDzID8z7xTzmzbu5
REF0/6wCRRXd0aXy9DMQ9laMXkNdt5KXMymezINeGaTKl3iP94uznPkcui9Y
/RlE2uUWwr7oydi3NNSO5xdRPQOvoxr4MyIULx9dq7PxvxGo3w6SJlGI9Wzc
eRBITTXytjMX3A2ntjD5cRgMdUv0Qt/7tGbTaZdYxtQv5H73Knbnsh02ek8h
RnqKT6VkPTmrs29pVFZTaoadQNLVVs8NJKlN6eTyzZQOh5q6GF4ak/fRHe6S
gWdebYSSlU+h27Cl7P24TlZpnfW7lascVpFJ0sCD+Bkdtrz12Sj+VvQ37ik9
wRulvrwIQAChUQIHnVfdr7iHbbZs+KvcYzt6uCgpZqS4Qdv7jO8u5W7FfoBt
f3yuQ6VFzMjaxUMuenpvjVuqckDhksxTXnU9CSdRHW3ig3BRsloNqsXuXa4O
4DYBr58wPAEjc/N4zWrO7exBRuTCiQAlcdVZvMrba8Cs+3vmYdCluLUWvZVL
GJdp7bGmaV1YD+HWxYomkCiMBAMoHXMvh4hCLpzPq8BQoHtv66DBRY/vrAot
JtNa1Y7hDO1lM9upaTmz8dJPK83BNe93yA/CXycA73CmAjAFfcBDCYxnKapQ
dZUmjNKYJGotV9uczeTAB3B7YsGKNRre9MYqvZDUC0QecFoFzLK16UwakTgF
54QuG+zORQ/n+nNwUzd1yKgWJ3lnPcyZmEDRqrFi+DMXBZQe79nVh+zksgu1
7rDyljWZjwspJJ7CUxGXakN5QaolWIVmSfFlcSsuB+lqlIMx1qeRUxk2HE88
JCKvTHpRPBZMVX0AbnH4QoFYdDPs/Fnty0W//epnVP8m8zeVmzliow/BLQhe
PgRFhvYY5NrPFzD7ojqkXoBthbGTXT1x3M3P7iEXjrvBPJCgRvhtIEyPsnTc
DJofig4RuDmSwDBthdve/dOS2DJXJS+/qUnj1M20cFwitQ59u8BAhSxXMx7Y
aeFIBnkgm7yuqwq9zmwnAGkaU3i698tg6Z4Do2h9rz2HlAB9pV2oKH6Xi9xL
dF8nkREq6jECo++E0aA2kgzaFMyO5mL8K/e8MBT+XiYu1/NSKjjNsla3YE+A
rxL1c4bNb0VG+dhQpVOt7nXTRa1MHUAFNDPCSbSE2XSkVr0BfYvBlf9dljya
yPUTrdf93UJqaMZTHNE4sAlVtLNLFUyJxBUUKnn6em8jkfXDp5uMjj94uITa
2h3kIoNb9D7LTVRy3kZezzfzVoU3D3QXT7s4grZJAEbxQtuzQHNnuv32iHuQ
zkfSVPA9cGZCK/u6ddkHK7jwA++IuS/s/mmgOmVLvP/2YWSjCak2hGIME9km
MO/kenrMqbteau8yCHwagVIZueU5XK35iu9YTee5MFIVz9rlYvtbv7YWOgTF
JrLO4wWdQmrWFMcHQNZB4s1iRroIU0WzePcb396HgSm+cxE9HluICmToiBbi
SU5NozTIpIhUpqqP4YOhXcDgMuzL12OhH7FZUVL1m7NzWfIjn/Nd58zuwC7o
iR0EW4syyO1841Vm9Z1YyHgG1vcr7boOHOeteobY1mTnMM1q5wL0EZXzOpPF
O5dpdXrxuLoUG2kuRQngwrXlE7eSiNZYBQBo5thKzHt8Mmt1AUVZARnCFLeB
ct23BIFQrPpVjJOvIud2oCnDA1CipNoh0RWYhU+ti1qGOyIQAdIM6o8G3vHi
XZ6U+G1kS8vRwpWM/97jnd/VtK1iaUaaOA3nbgx6d5OUPgX3JQokN7gj2lML
KbOg7eFbiE+Wn/E7ao70mCo7SC66n0UJM6sWGLXb9B026cmWPV7a1XxnKPxk
xXgsGfQBLUE9j1qmOqrgEKempAD5bKC17o7S6lCHviTvYXn6lABN8wiORAGd
pz+rb+eAT8NzEdwK5WFszcdRdTOKffvTn9HL7v2ViljDDStXGkle2mIGoLbX
xP08nkqryugTDXPjYTNkbWhf0xY5DASmu7juVUmbMNyNZY3xnf8sS6cO7BXg
NiBbh1cxNH+/YcGvClE0onWj4f68913QLm3fkTVAwbJ4602XPB7ie2IfmA8b
MpxrvKGLyrKcnvOvGAhlo3Ss1sGFYksqjr0W6PxfC1QM3M5Fixyd5x/UV9JJ
oCTnw94JCIIiESxlX+dfGAkQzdYiEtv/Bmf0NyEkSOgG9+KGic4MbUgjQm9p
1yqQTvqd14gjqhCHBMK5OoMnEI6jBNpMIppd/dmr0zAqJXTJZUGBTryOPpb6
lH4UODPe8dDYkqjNQj0vnqHmSds5tSZc28O7Cnf938kiKe6FChgisN8n5uKL
2F3LRbX0ohpGzfpYSx12P7pAL+nZVs/hmMxCS/2vugsy69OItI0KMpbCkKiz
nFKNszmcMI1Iuc+USnfrRY7FIhNVCwQ53dxM6jCPkQ+sPMUa95FQVHVM5wtj
FenCP/Jfra3e54tnOUCg/iVEkaHv8k66+r1mJ6h5Sj3h7BLdS+G7YBHgQnZJ
c/7dCj1a0de9APCOXNARamH5p4tewu0CURXrnjMmS63/cOsOAv7tTK4Z0VvC
L/0tN6GLb5YdGoQJXpP4I4rkSEAaUgzrZweO6C0qO1eb2+AF5ppnuWE62vNX
mdIXv87mgBLY/mUhQ4ntaJNF0BPD0YUeiQRoQvdBRpFPL14/WWAzsMvKrqKO
JvO4FxMUu8ku0pqjeMDwIAIiI0cMoPc3415USxt9b1wr6NETmOMJxmSvr7oF
656/6OQ7yuRL0J0UQb3Ts97J9LLjEctyDxGBzGLQLIB4TVDz7K29zKivJQSu
zO64Fr9yuzTr+Mb/d0uuEDY3XpQ+MzX06VCEGGPHRHLFlGrkrvfi1Izx+124
nl4saru73oY6dXTyPMogPs2Lo8rYyzfYYdvmf3ImUpRGrMktl48LEsFnrQBQ
XTe0mHK4H1+gME4KNbcF+gmaDHNV+LLDVMr8dIQjbFbZG7Apq3zMx9A3ttko
QN9IMtIfXEj+R2NjiBkpomxnQoptzjPQ/nv2xZW1FNQWDuSD7siGQ2L1aJHI
TH+8+V70+ETPezEb4aXuODATggeCad013SOuW6R9AJ6+fi6PQAlstV56uS9C
JNWva3qQKtltGvC4ifNKtxd8rZxDevGe/MUoftVCPNW9m/greN3+HZWY+TAU
mmxG7WPSij03UhtwV5XtEqnHnEbRgkRRo+/jRVbulZU01opLJsS2NYLpeQQm
bJGB3PK0WhYAdJdztxqbQg6lS+OPq+0SP5K/NJnqVO9lIXrMIPq1YyVKpCJJ
Q+BYeuLrCrZu5D0oOrneKOLmPQIVxbz4Q0PwE8YTFDhZDQNGC3NyADDXNKWu
Ah2bQ55SbqUMA4A37h8TBKaxnEn6V8s8hRRFdawEF0isyql9Ce0Z1Z1/9Ren
mVrDEajjmeCDgeBPrCRUugRnrNrcs4BWLfPdhQdw57Vde3XLWxfgP7bov/0n
M5wEoIQGYBBqUMXVBYeJaw9MKs6KPrcJfXT1N76WXjzuxNFuiWPmFKamemur
DmSNJB/sCBmHI+QZWzRyxf0y1LfkRFR2+oJMCWL+K31AfitlikWWn5DKUs9E
9YMM6xmMYhRkBZ2A8cvd68TxUHEu3FUed+reRaN4agsOvVfNL8HC4jecnjh3
yFkHW7arx1nEL3s2LMMCDTdojPyRXsS4FkIfaQuNDY08BIWyQJxYgjDen7YD
1Uq538gpFfIf2q0ttvnm1rji5E4SyEIUxA9DNenCB2A4o9JaRirR5Dd39QoT
n4FiTqAURaR6WT2OLpo4YG61auV10V4dHFWPHGv5dmMqdWC2wFYJNR1f1F6o
AiTiWP+ZiLiP3IUKGjH63z7kIl4i3oF2xhHNpebdm46BqGRBHDYDVDrTMIUT
1y3gFgnQm6lYKjfzGAL6HHRZClnZemd2IsF345dzRM97y0mwrXjrOz+t0a8j
ZdddH4BTM1vwuClKnpMqEOk4tHlpemrBiDwbijhGqma4a0PVWGHNBM+b2Gb/
JBRvl8kSluidOkCwdo3HK0bml3gj2Nn1AbAu5UOZ6dA5GOdxCrLKqanpH+DK
DBYz4PMvShN2EK2Dbu0XbwHOe/JXV+gtRTiLQMaabG7K4RZIoLYEFTy5PtIL
bOCSSWp+jJ86jOjFISWwlfzQhWOGqSn3sk4MSbikpuCgR86o5IMJIlLJ8g0E
LhkhuqqQ34O+R7iOvgK4PWNVidqur6oBwgPMxZybE3Kxz9uOdZa0YPdhGCDz
/0VdrXxB7I4dvP6t8pYxphGYsrt/grK6grR4JdnVW+IFF4zhpkHuN+NqIrF0
M/7Td2LBLgfE7nBpLLqtRNVR3/E2/IrilV3k7X0DnmFiICyVkYlFZmfBq+K3
42+6M5339AGRSFP0bIlkIVQCPDdO4yvx5+Hj0Km/SjVcMre2P9xQsiW8V7WN
bvL4+5kaQf+XIfGKLKuF+GXkkCWTo5LwbZGG0AXeu0rnVVBMDUSU5rRiwmzz
9sM/L3IKHpQE5S3YudPTpSkh8nbQD4eJKq2yV2TdGuG/lPhczGTMeA9WxKtJ
ydi7BJ1T7toausmOcZtWXfv/v/7dp7QG9lMO82HjplGr/pcPp3D33Zas3xD+
0/QTnz5MQOwTn4GMYtCZl1d+YTh5XW7wCX8g9n9AL89SzarZdd4uNI8FGrPO
rpZcrsi2D8bb2Umj9uLuIS5guf4KVYLlkEVZCp03LwFBCmDuIFy2hE6VLprm
lyCdBTNPGi52I4R4OmBgj2VAZxq+PqmpIFVsBS1SMKz3WvHs2Jex1PcTiKJv
8lw71GLv70qw+nBmDQdaYs+SgDCZMj4oWqfgtodAovDe9yEHlKWqWK7cI3r/
vX90pG8P77nRg3xxtGimfSZfuUDrzv1vaayFCCnO+rKT65NjXR4QjcNhvQXz
XQnm/TqNnuy6769U4P0/l2KFLgULHkYf49XYYdsVq6ary2azaHkrlPf7ClTv
zScad4xObgAZRcG6BsBC0m0sKD0F+C7J8EfrI5ft6tLQ4sdcsR5PrVfjdtWJ
ZiKw2TY8cHtF7NBJf2uZmEe8H/5fuaeclWSIW462xl0rzLDgCEd0nptXVYtJ
3zbc9bpbpjNUX09s/MwndSogq7/fxMhm/jOve4R0JZm2c8PKkhlWvJpRUvWu
7pLTuzJyyB+f4Hjvc2ukFHWMVeUJ4i+htqBzs9IDAvagXOw3aJ7EnIjb6+Ll
oiUZilqCDQo9hSKBRt0bqh6ZQ7ZEosVfalGozgClEioLcNptnaVXeKpIk3Z0
QyHjWKSLT2FadL21yQcHI0fhX+3gXnIKPvlGaYLjaAR0tXxdIkQMeIk0povY
DYLi08GUwgSHmEMUL+fHrb0L7Au7kexEdL8EAa4s0EJnQPQjZ2PmiRWiZ8bA
UuWEgV5sa0OukBtyGPdsW+Idy9VqyW5LymKNj8BtEO5qje0Aiytde2VhCn8D
76oOe8agioe5G3zJyTkRp/3soCa1s9YcXi0D4mmVzmyZk3HAk7J93mcO2Tcg
wFVw3DKRIF+9XLHcp+bh7ZvcOFYzcztnrZchDu/MdXd8Y6Y402mQXKkxYWIa
3YsgCVJ9peP+ECsHYMoGJtC4x0P23s02r0R3OMnIrPrjJDIrDoJDnYGS5CdV
LOXAF6ECpzRmMIJ03RCqxJmKeTpP7iwQPuMwIIOmJCvOESY9vt8wL389FDd/
QeQziGZsenT77lS0h0/5R74KVHhXXgIPEYJWNjlmYtaBGxBhnkofsIWNqWCC
U9nSdVYycvXQae/+QHoMWGSxjBdLaEeG3b9+hiKumcdVc5OKFTQz+Gipb4kc
fXJ/3d51pfjwkCF1/IRXauamf5xdOFA7BEveIw0CD4ROKPdoUIsh2iPDImaG
1TKnvyG5gNQ2S6dlXJdb/MeEiDz5R7WWmb59d0vJqN3GsNYG1vQqPDg1jhMP
YlsFnuaDecNEroHE52t5a0sbVBVGhaPSLsTNFxhHSxqUYbQs2ZHYGcSz2+MS
NR67WSnHFUBW/BcYUP8Y59rr3Ayttiwi8SzUgLI//ZePQrrKqg+akMiNNhyx
nZ/3hckYviK/Nz/otepqPD742Zjms28CRQhM21vf7iq1eXCdqwKbj5fEQsWY
XmXDFhWl18wigmJYriRFXzVBfg1Z6Vk1QeUDs1M2MiH5VH3cBPzStvYFMUQV
Ee9kMh+ewzhkHjwzOQ5pPva31si6DnICHQaBmAUwdm8/cuoTdtz552+IUc+2
CZ30AM93B0ytqILO0AlJuVqAp6vgQRbtQ7xj3Oe2em1X4gFn3PLsZW+I6anx
qimEITvVD/4YW/Alqze5AcMLIhFRiMKMuTiNLyTexieNdjUYeZ1LCv0hZtjz
ixEoZO+jdEjhmhwJGRG+DZq1yWuHliGLoc8JGYTsRn6Wyz1Zw7Zx8u0pjOB/
KSjrKpXIjNmP6jF4FmmiSMFi5vFDQLEWNtSb8kQIYTaggZjN2uoyHstlRm0n
eI8YaP21dJgxDtbnjJ+jqPDORTx+5aJcChbRrDpvVEOXYQyf6gK29TUhQr8P
x8S+WxVtffMppQgawt5VEwPq6rf/QYsL689I1FnLjYxOcV+iL8L6RtD1XkDd
zE8Zqk8rKlEagLKmMfvDX614/o4tqTxqUJKU84YjTGOvaHhumwFi/2+dezsS
oYVlHFZpM0ajaGrW6xOzkGHaccV2uQX2bsSqnBq5TxuSwnnM0SL4WTT3o0b9
unIa9DPfrafFP59KBURrM8UXwsTfFcuL8bKDWE3V9qEU08eXMxYQamYVvktG
aha9Y0kolUbksUToNQwJ6jMBg9QBwDVktTKEIXzVk6csm6qw+3GHAD1T71cu
jtnYjnC9nSsXo2DhrSxOwpOdGuESwX/m8x0Eazrmzif7V6BXDryTNd3FaJ+r
Sd5080+4cm2dkfUXYXrF88bWLeIELQr7yrcj1GpqJx8zxNOqUjR+4qOsnKUl
de/Byp0M4u/I7k1cqea0LjEu8JAHs5s1chLtn0iGnjaWfJRNQFRSGES9TMHb
NcNq//w1qPkI+AXMFbSt7yeMxTg6f8QgFnjbr8aF+VP6FfrucFbjFgtBrmpX
NWeay0abElLxSCCRmSFrUtuwc/mJUKjWuIR3xRyCIfguMAVvq7syBrbyTOTd
d7oWKQDPcvc9ZyYCR7Yh11AHQDOfAo2zoUccxBShlvzgIWP2TglLNGXpHp81
pGApEgYQ9PGmV+5YPmVDmJKQBK9W21iiEkZwomAAzsvhtOQ219tKFugepB7g
4k9AOP8GKojpxgWce4DVYDlATawuQ3BCJnJDoJ9xqb1lsSMvjN/6HJqn44uP
Lm6C0PH5Azt45bn4jn9WFirlxOF0LkNuojMeVBQ4CgPruJN7oVoe5ofTQnXP
25NYExdnk+8N85N35FJs+Pq+RsLqAaRbOTFf7Zl7NL2uLzrmXFjcPkHWso0T
N7l5031XIJnNu6py0ZU1mcGx9f2lgi0ec+hVvD6AUgH1E/sfXnt17H+FB6Iv
eVjxEbzHoXul/+cRHHoN1eMAkO02QBWGtI1SblyIZ7/WD+zJE0j9KO5WSGR0
7NyhoTgDMQHdb1BsZJKDQUPml/JQC4U+rSnLN28ViqSFGvLa8F86ewMYm8Nr
Yzs5nfQNMhDL1ZMXPnBEyjRZa78/KqywNoyo9DG0iRX4UBAmZDAJY0khTNKR
xOst43mNS5eit+0sipKmzh8szxpYoEXG7JS6SfDdnExX9NI3pEuUB9c14PvO
L9p/HZAdnoLk8BNUKMLu0T2B9pXaBajaiFxgoXXx9hD8WoxgPfUhB8V1CL/7
k2EMNq0n6XHa8/JrN+rOTP0wb8CTELIhAM8qNdJZTxnkwLe0C8FMav4oy77n
DYGfGbiaMXHNTWQKj7un8hQoSpDw4PpFrflRlxfjXcQAMSd4CvFAoQ2joTC1
hYktV3hUnTf82Y3gmNWUXEYq7u3gV6g2/09rSabNDq5wPjIiv50zQk3W/2/R
zI1Pik9Ox7H75ACUi0ysAHQw5vaWp6bYg3pz7LymdfQFTkSWGzdoCZxY1Du6
CnjsvOXTc4XDyvJyrdI+NForqGa6b+HZWBEhRocujcYCPOF90TyXFTqBHYnl
pFQuW5AV2UHmjNL7rf0bLQYWHaotDA1Vijft/iJsBofcEKZc7tWP/3cVXBwF
DcE8JkMqe+e8JBTW/o6/9Z0UB5E8avuprT7iToN7lC+E2QcK1Trc3lNckVgP
VUlCazFuCG7dqjVyR75iUbryxAVTPnD3Z3CugnDSaT4hDd6qs21nQTbcbYe1
OVV20Gn716jDJi0i8tST/6jKr56/32H1lIrU/RxLoOnYa916gUeVUas+wcLb
3yuQ16syUNsuARpahsTNljcK8FtE2UATUMY6sCm8i8w8UB3IeAHe5DhYcojm
4LtcOWlc8sVUAQsjlL8EcpdO4bdQAAYIY9WB2+cWwUsF8GxIpZCMxZCk+Wd6
2sopxI5wpgoQ/pBfiGNE38qhlTFDoauAnIY2oenNtbWARdtWH+TbJaObDFLj
E3FlxuiCxskXxSZZkNo1qdOqT7hg/WCrgw8vnyhIt911bgx3N9WBhFeH8boa
iCK/rL394wXiJSkenhL2Ewh2GrCYZKcGbKwHFfW1lhCGrXoN7lItW1TMykYW
4dDpHtK4dgqWe9dt+Zd70+GGe7RP3eHB8Qi76kfEOQdLtauu1EKgmY4DAmxw
3nCYVacduR0fRKOYxpZPaeRCz9ut0eTfUnwe6v5ih2vXO+IGZbLHO2j7N3dQ
PCcnNWsXW33mudDxdwiIf1FQFoJDMo/4gdu7+KJkDbicfVbYKIqiV8lctZxA
ITolQOkZWlxYUYjFZT0FVkGWTg+cMZWF2GARGL1QhFYZoRV1fgcz9OW5koZO
YcwAJRAvvR16q139UeN+we32VE4uFsq125LplS6ScUEtaumi/bXNG2Uq/VU2
FMs2Vl0ZxUQMLf1bdf6OtjkF3vbJBjPrbsMmptzExum+uyz2ENgFhpsBJvAI
9uO8PqbX8Zpi5f6YtA/3bfA30UOdPklJzcGXvp+j7IiN5A/B+3DIWM5JtoeU
nOk4+5Drts7Z9qOXNTv/MGU9aEJ12j2iyvj4a0CS47IyHRt+yLiXsR7AJ41J
uiNNHlk/H559NCoCr6KGzcui2Xa1D7DBAyNyvbCJeWOJ6lrU5zgbXaCWy5df
uVdoxvIpiYzHrY9Z/6Il6OCQgsjVV9vOUyOT8W19NLy8aFu8DCYGz9J2B91p
FKcHLULstiZRV2+xn7OCQJlQ4kwjL9DIIsIpHv/5d4YeHCOxukr0Sws7KT5w
kqvkiF+D5FVwt5nZOFCxseBoSdoiJUFndtADbS/OYSZD/xtjIFzpehywxtLc
og0OukvVUhtg3sqa1/r2oXM7PNC/TbUu71mII/aXKP20/L9FXSgDrWZkSLlV
jYveRG2N9hncXhG6QGzAgE1u6wPCjuq+pTLlBnYLyxaRmVO73z7V/5MbXHMC
doU+Prr/V+cR521csLOb8kdO9zwnvL/RmpWRfjcPH1UnkKkzaqOo24nFkygm
YqcjF/QnEOR0hNDJRHK5zcK8BbbQG8pM1BF7i8IzgK8hzA/wKpNrRykmb0tF
6fUYmEVcGoHai4QJIT8+twgeyGPI2XvQbagfMjlAWtm7nRj5AQuLyVPdSENy
47uf2wk94ZmFLoOvLb/Ch784h9unNQOOOjPVuFoId1MoA2OELPDkYfSgBP2+
lHiBoXkzsrq5bLpnr/FwPjhNN0Vk272VjFOAMcn15hDQYZm1kn7iHFqKN8bA
ZU6H3R+9ALbKT95Q9TIg2kAUSTvAziMADfEZ4LiuebZX+8m0//KYDz2goBDv
75miMLce4Q9qt9pDZpsVMeLdrQFck5E95DewkagYltdiH0ovIgmoEgL95WFO
qd7ia9E2p0By3B20dopaUmFjY37Kl02DkfolUZaixK6gUnZs7XhDG25wvNvC
H/SQhndIBaJEODjQP75bJr1SZs4ttA+54Ygy2UWEbG4d/AcSpoiIiqdur4pW
kDcqyR6yiIKdIdaFSL5JnCYQF5O/Lh3B4ovzScNvD91/dtKvcOPF79NDixFC
liPgajRmHr/dieRwQJ9+qIplzGX7Sg/cwbnoZXXnmvq8lXP2IkBOWLk30PeX
VzUeRYgUci2+CM8NR6KxblBQgo1xHUJhD5ntPcustIyYsQKyDLFYduYdPjWF
hP8k1GRjftDE3t8UqBUHBtVLLHy2e2ATZJ0qtoD4Kuj1R2DBivT1LB2yiTIS
mVDWwlHxqw+2EGyYE+L6UHXbhncbhHQ4pOArnmlvvVWvwDz3IZXT02/q4Xd7
kwc8g4eKM4Y8rL/ioDQsT+LkdDi3O3AiZGe4u6uVquQFnJ186ymVU2BQH+Pd
Jvhj4Fi9Bj04gZMevSDh+AdzEdl3lhoGKNB5iu+Q6x7fXESpKquhcSD7kyn8
hk9QPIIM4WTJMaMjO4NxQ8ubmwvDDemar4PJAgxsKRGesApQJ4AO9UPQsVPz
D3pROnDiIKbC2P8vionYnGEPOO68WPII1f6g5Q+PY5hz+S+Xh3/GT4zJ1yHJ
RDCQ8+ud9WKvYCi7oLAM/Vsw9MbbeZRGfhX9iJPJJveDz4sVpkufw6oh8FqM
qV+O2T5h0J+Ve2n0rU31ukWXVGs8dEPnK3IiR3Ri7n/kj7JPDeUNXQ7mMIER
idMHG7Ze4BXNFT/9bqhs9QzGRk4FabSiFYihYv395lxgiFPN9Cd7TSM+1pNQ
YJWEPeJYsz3N+VCtijAq1wOsTQwHvdHQJjJGlFFII7XM+gJ/m+Bu7/ooIX1U
YAyQTmahyxKZYbka14SgAp8KDVL9OddZlbWftUOdmMxFBvnP+e78lX0pYyOD
aRV/eb7X6POHoK9L9DlI7lUhC3b792AKMcXISWkVa+DTP1gagexFH2YiypHt
NwBoK9iea1N+OOPCC2uHIL03hZhVXARFG6M1eh1IWtP+8sHhnZ4mHhU67Ijc
f5f0smQXBYNazwigXlJfB+/OROayW85cAWMYxwubS5LXMGo7GFWDQz24heF1
DM183qkOhv9FOOMWSfLIbXo7JQJt+CWH8W3iYqxf8z7uypq4w90FVYDb2fIx
vIZ66/o4jZ6qA2EvSRTM0JrftJCK7kWC3N0C2p5toP/DaB2za+lqWbS85Cfx
AOrQCL62ig+T/YxK5MYUJ+3KRbpRS4Emjq8s2EdgV/D5Xko6/vncbiiOwP2I
QInsmj8zwsEpafwL9GuD+z7kEdnjjrrYJa9xb9y1x5yBPet4qbEmbMHGwZmS
BqhKMWeX7qbOGZiEJ3wOADaxtV04go4mgZiDD8+8ALS/UnIbJgs8LPhiZ8RT
veLEK7mf/lztvvFIfMPDnqC3cMiM82XjJ02ipwTtnzDcxNJJP89Tv3C9y0lB
JtJ+2JhU2nOPQKBeFACqh3YtCgBQUIoSe84N1VDpUN59Vn/ZAL38yqQRjyN8
F6b4eg4jfab/WxsVjEb1pElr3Mtx0cUn5WOeorG6zQR1zPFBHRvqgNGkhZr1
lsMDg6q76E0yp1kgf9manlgiPmBaQe5woAkkKfJG7fCSyed046kRuN8OfAnt
i3r+6aAHo17OHXpPL4T3YhRYWuwzKK/N1g+sCxrbNcUkLGf8eLFXKgBpWCzg
hy6kmjcfBWDHC6IDWMWl8DxOm7RQrlCl+Wx6PsMQQlo+/6FeEa1GMApPNgf3
UiaErTXXq5MIdV2Khn1AKI35uWv7Mu5CQblEKhQyyveH4fR2iwUY55qQ1Rc4
RdEWqjcFDI3q0n+/9IbdfaYg1cu3y1rg2IvGhDuvh54ICCEnXru0rIaZaxwo
CDq/7fJQCIh3kuR8xm7xCOUK6ZK9VnK5c2h7KaXf390AQUiMYom4+v+ZE9sC
8u/lXwuUoJhYC3SnJuMJNi07ZrmnLWHMqjZmbc2x9WghUJiJZF9t2GohROAM
/5DVByf79uYo0MvZTjVNTEyua1AflBrm0kcQAxVx6rH1WK6NQzlWi8NQ32LP
KBjBX5hozX2r3zYPq7p9OITbwcGCvtwfbpdQaYyN8nn0GfE4FqsLWerh0HAB
QZT6E8vj+1lRQXi0WhL4gpoLDiJhm6dErgyHwnk+sIj90QDYtSjJrWimPOs4
b/pcZz1klcWs+/1+nSq8R3svrO1lf3kKB6n5/69d60x0vY9luVTdoB3CUwaQ
TVhOzRA7BPA9lz0xQBRBPUkqB+7lURGUGUH7IbFP/pcBs9YCpWAS0Ey1WDic
ttKJKvMW5GQ8eqxctza9bhd2wb0WW4lIxS5U5kL2Ta0qnPY9HpT0vVZugkps
bOeMBaINtat0FcLKsEvSQ/nDZDqujDNI47MJb4zZt5XVv5usUev5S4Ur7oJj
deYJylpSnyRivWj4Z7u0GeCkeokuFMUdVa7EmnHX1HAVlhvGLGOqPJsK+cc/
osecIImnp3G1Jv7wZZqA0BeYvKNj5hPut2fbGMO+qVL4o/yFPv/cvFc+6sY5
uTqJqL0eMUbu/mpHGr5xpu/iMnKlNLpkmDBkRABnnA8XNfg38mzK5C8MjId4
xl5uIVe0Uj//VoYQAkMhx1pHdE2/VaQh5eG//ah9DQGYO41olWqsRhY4y83f
d7t4ijijjXxvlNM7NCxT8nfIKqXwwTAruNJLlZ2rECiQcF0DyEdKGd1daQUp
xlio1ImjhPj958j9Asql7eC40mO7HkJwRmiX3/Nu0O4EZ8D368pfH1jsRkWY
ut1rvM1iflEYWuZbCDxTHGXOOrE6bNUTjWUxO2XfPpQbBt2+U9NqQJy26+iG
mbE4wl9VtN0/6D2z+HAOrNP42GNC+7iddKdJd929jEboYLCumQdjmbOSfIun
8eJ7rHNNsL1299i845UUkUHMgkhEoOlZixiDpg0xxEHwkGgJ4ATwnJAttxAv
W9j26diGnypDKW6fKs0e3Pp2lYvpiIv2wrDVdkr0JPUXs4gNHq23+UVvg4qM
X9v9CmxNylrxRt8gi2LqQfhBDx2A6rv61/eV0+SbHd2j5wwZ6agaUX3L9RyC
OGsecXRPjvUF1Jt7ITP9Ghw0kauAX0bCrqVWsCs1mrHd2eVe4hX4gFB2kVuh
4f328MfQ+7GZnWiZHWyjdivMUS9XHSQs6ulVCMEPP8fs8ROwh0Jiw1JGAd9R
h44ulPQkIx70UnzxeSvC6Ska684qn9MnCu8yOp+cN5fRIS/GDoMgNlj96Sov
zta+VTER5okudQ1SqfxCs2hAHO1tUnDwU6Qnfm822QYwGqccLTNaMaAI2aDX
D0Hpb0tY+uW/ihU3unQgGlBl5a8aK90eP6PiyVnzOa2ra+b1CKcCQ7NYdOAt
WXIrWxOJJUZPUFBP6kBbrs6pixUI+uMP+llR6hcIUy8Uw8cOS8ELwGC0q9ed
b8TVGuuS8Dd6ndYQfE+hmZ5TtSCLijrg/LedL0VcXcpbUFuQegJjAQTIANin
ewSNkRXYD/M/aEn0AlxuwoaIrwEaZmxnWwTDB1sIXEHzitClO821kOR7mew6
xGiIw6AFJ56qicpAJdOqUp9FgTE7HrvEeybR6LA1hBmrjgtXg4xgZ55g9biY
EtdBzFPeUJvgIsbWhEzcjwC5Zhcyu6rbFkl3NfjIU4FDR81Rh7V+0RviFQ68
/8fGtoHM4GXzmhmd010IvfFU4Xg4ZqYNu9YIQoO89s6Kh+Dg40ljJ6RJEUiV
PEcefwLeJOO0Sif9zoqidBXeczAboeBWjkCDlEU3pGCIOVuol4KQaQe0xLhP
64E9Jnp4l+KLjJm6Hwl+1n99CzES4ksJBGkCKmuEctS7H20BGFeUSAmUbzZ5
OG49ajBdyN/UYvnPj95cYeTQ0k5TyrpFc3NSWoeDMP1nep25eUZuON1UVQPR
lk/ZQ2AyIfRg6eWN+eiXvtVtNCIL33Czkx07woSAb2LiPYhLbV1oE/G/UV5Q
OgZNBhSaokDBGxEtNq7usDvfUK43VvTw5AQYb9/S6cMG1Q7ckKB/9ltdVLTJ
ZSlsVlSFoyW+1KJCJAOIk2+mjbPot93MSA1+tmcf1ebRRgRGpfa8cCPYRsqc
jJ1FTPWDlOFPYvHbtkchSF5Bl/y5dkn15CiP/lki/EO4IbpDeVKlh+oy9HFn
0Y7vADgj+2QDlOo+ZZ55y+M9mVjBbXgufNgRbJoZZXunB6TtPJXg1Hs64ILS
QnFozPjsIYeSETvRZ0UUmm1xIDIAd4JEGI7JBeKMCC1+ZgKiegS/ipybq62S
qfn17oef31aW+6De55KTTuBeSOMqE1DvVamTkHtGuffO9swQCdAtYkPgT9pI
v90ArzOLy4A+gaURg+zZKV72aDTuUr3LVqBtRaQ2p/ddyNMYpHY3ruYfZJQw
RA9oGkgauje6JmclfwmjcqHHuplV5fqadpIvgI0nLVHYvbuCENIygD4iApR+
4nk3uLnTk3sCkS7MWg8EorkftPZGPQbmcrKJljiFHeIttuFcUJri0fINP1fJ
xf+K4v6Du49v7KuY2WvKwCJAtUcR57jS5vXYSF6mFfpVqbepHXPyOsKlRaUb
G2t4afGCtIXhB9aHV7GvFN0byXfiH3Pz9z3X3ZcJOi6fE1ZCTr6ppfwXGrgW
yIBGpBSQYMwvWHaZedfUMBlXbZFx/ox6JPvVlOAsCvCWJwjvFu0UFogxzPa8
sbQA+EOOu5petfkPzl90nAi63b0OwyiDYZZ0NaFRcNZsyOr47Q3pgaDt75tB
KGCO7uDiKDJcrQmMphUbEf8dxNgg+ey5S/3kjnEP8szlimaUrYb/txjR019t
q5XRG6ZqrKkiyWq5kzihFQA46gubJwE6XMnSS/M0ZuRvzKn7ssf7GkS55BIE
rD7XgZzpyXXeXjkfmgwxuqZ9woCB6p+wUAvKZuTjUNeYYxcUUKgfOQ2kA15V
vOa6xy/KXLDmeAfm/BNEKS1zGFOZJk9eOKHytrHVHIhKVQHEKmVkjwxpS+PK
k60tXD/0ebnWV7YnvuU62DAdhq3UR0ASpb0BuN9OW5d6Ub8UGemwx7aeEi63
OU4VXawJlReW8Wr/QMmxjnbfI4y40n4pDA/NbOnmUO5eAQeHZSNaZ2bbnGUg
SEIQfdoVsvXVEYKpP37w6i2G45nmojuXNw5ST8+bAvLWT+oIatJPrMHtt9ND
hFAu6qmjgJMlh6FcLK6XxSgoR5/lKLL5I4z2xMzw8Kl7xXEOJefDaMJfJhCc
R0ZuigOUDl+lu4wmEotp/La/zsYZUJnz6xZnczqzW3rEbxotnMpfGNNqgETe
jBTNpBnTPv5k4LeG5blHh07Cizb+yx6tUwOcDw8heDwAuaCOIHD7Ib9HCc1a
3bFunX/4OVAoUhya7GybngjFY3vH2TK9urXKfW4+4zQg1pI6b949/kraQ0k3
ZLV9yPTG/zPbsBM7SOBQXdQ0k1OEq7Dumv/lQIg152iITWu7uXCbyLqf+8Ej
CLhJTUJWD5wQF7gFNooqCiJ2g8mUXtYMU+c3EcgQD48s0axMN5hCFMHzlozz
zC+T66p30NkYEIFaVjEG/72tJ48XMWQ2r7+3JSjkvFlhR/1ZqGStzblDoPHV
gdQVmcj4YsfBB6RAYEBqGXSYD31F6E0qSC0I633OPzjJePKQAnsHZevCUGFV
DkS7kgq5rPTmR575YoigvcXjvTjhGeJSLtHzbhyU5s/hUfyBmNu6mXjWkzJU
iPBtBfXx1Ux45Z1Cz0K6XN+cYXSFyiC0aEPb0K1DWHS/K/quPJXB/ZJOHWFv
XlljicRCbyr7mNR4cZ6F+Jyc15Hu+ff0RiWAe2cARzvBbRVhEZwer/yRFleq
e9KprmV/VODZyP4VzdRLcag8Wi+LhBG6vwHNsVPndOmgqqcCl5QJWv2w5jXa
yUj2VFc+lDb6wX2jeuDQzEaGuDdLwgkhUVO96Jc/XddpAO/7a0Q5RBw6rB+f
nnjMecUdpReHoZjvvl5wpEeJAr33YM/SPKYa3WpLJK2GSE316tJrlITLdcI5
LDsEpeF45Ck7C+AmSxCUJpktnxMYGGJjEu4QZ4xI0Vyxf1A5/56WV644V8EK
ZnASLDkMDWG0m+Lz7tOcOy+RUdNWuFOjWd9jfrJpz8+F2yksLl2Td/Y25es+
nslhCoLeSp0Fk+P4YlopomPdEWaAyyLTA5AhqzB1Xkm53NW3zk2TOhdmnRQ9
/4YqgSTp4Jwy+cphHm6kUT5+66AmvcwOEOYFkaFfBojIkPqDO7/5XR4e3018
oQR6KqaYfz8BuvBrx3khldrbmkhXkQQftIqsBORC3r7sK+n1OU9OBhn63EWG
uc+RDP6PIIqU+2Cm3ZelYt5E9RXWfpyQ5Tom58Mta06mIRYY1QAIM1kVikX5
N0AVYyJEjnQMnlRR4CfT8XVGrUp8OcqoXP6nJ0xSDbaSAzcKADruzGws4BKf
RB5yHvFB5J49/rNmvF9CIaYKT3XurAgt1YwL45XPZUe1jPcAVw6WOa9v/LvL
tFX0o/ecROat3GvY6AVbCYyut/BJiDAMBWo5gkz8o7klDzIo8Z55zQITGpHt
J+09V/mTvZSnbo9LoGYb6GTUYWjQBvn3vKV1sycf2sEb6pdrqwbFqjhp50NS
CDjlvcTZJRQe2ci7BTIDKRNtYkYTZeQYwLjprW3YLe7CmWUh3Ia+JvPRGPdH
mt2W94YSTr7ghL0Q0m1P+uys+EdSUOIxE3eTEDyCo6ZC/DzIRCM4M468J1SO
EXXfJU3jNr7aK+U98+B28xc5LNmC0rIWzMqcUvOlTLkbWkAEOpwL2/bqP2Sl
C8+oLh5MawdjbiGEp+rKkuCSiDGwOtLKq7fmsrzZ943KzSkZZjaDm+9zFoBi
rtSsAYwDu8w1UnZvyC1X/OIwGwyckRcBegoCPjM08lQ207UbzlyhK/ysdTLg
pwIo8qlcgtIZx69QmcfMNXjDVtUp+FAkeTw5Sy0a1Wn2rapIK0sw7gQP7cRU
JsBODtEO/NU5Ludj9ZxZxCo5Zy6TfkzR1GtmNvDFx/osLm9/uod7C2FZ3d+k
6f8gGeF+4DmWtuBtl4WaoEJrIZ6wZ9wS6hoaevJVbyVCuWP33wstLjmqyil3
RBhknKAhwurRBUPr9d9BXPCIc4guKw9WhmcY0kOgbZ9/6hDA5CPaM0OOinFh
gF++RdeWUp98V0/MQ8e5VzMHikSFQPwrFxkH3CFNAjaH5k/vPalR9ehtrJUK
vIKMUVorxzIpq2yMwSZ0BWHQp577tdl8oqzmy7I9ADqOY0ayq8mgBBTk84OG
mXLhCKOw9y1KBvjaXTu/SR5pc1nkbe9qzrOG/sg9p9W93X3lsPhP0e7D/EeI
tMb9QBMUKMYNz4dlj+5wjoqIZCxketbwJg5xLzw4+LENKbLHj1tQVeBSYrmr
NtJvzlfyZyPnKhStaFqEQJ5e9ykkgNvtdxoaKqk6boJ4iSu/32fhg61wvxdB
ASG8YxjD8rWlo96vVQg+SWzjAyFUk+J1NS2Uk4VIb3GjcI2aCPqIbgby4lRt
J0FWy87wkEcGsWDiAtUxYqqZl+P0tkAWYWDUNYkbp4Sv3y7gbd2csi/AmMoS
7aeTr/TdgK2ltc1bpdz/P8VgIC82ymGfFfLVjZ/daA3fTDKKC2+WeKiQOAyW
+fGmfR5om90tg06FXxQGdl6paj5IroEjPkSoMUGVZeUEx2n+uQF2eM+arw2D
pIg8LI/te55tiS+IK9LSoRA4ezHzO1aMc/eNG+LkTiGtgBdw0kgse08I4PPe
0wWUvbpmPGUYVNtUtCi+dDgn4hsjNNTZkfJO47xuZNNk63sMLD3pmaf88y8o
+1Y4JA3FRoZeaEYJEOb4mIDudgNuNnllHVbHggLZ0lDUTvHIYcDRu8UF+jF2
w3BwVnguWHyCYyS0CMV30RZSfKPMbSNycRIU3A0GbU+K4RVH8WybFv1aFjHu
vixEVBeuGWaf6pZYjbKrbCxw3SIpdy3HsxQ9HmixXBXW/X1eep9KtzGkRhH2
WLmio2fMiaTg58MQNhE2Kyc5JdOF9XEUGiLLkrqBlnKqya64LysyckTUk+TZ
zQWKu3BvAtsqpUo2FOFzneqec+elh5WYBgrv9oRgK4xa+piqMmzs6N8aqsQO
GwQrr3OZC+LlACdwQTyoc+12cZrdrScDgblvXdUeuSaps8YgYDKkZasgoukm
5gFklVpOrFjQBpiXrEm7vXXNFOCV5WfGzMmxpOoU4OIWhrROwd4Tojfcvf7N
FUWqvL/t9ywOQH8pXlyM73isdtgCL+dnsTlBxNZ8iCKfYTBzPh+v/VweLycL
MJAVe17nC/SMrOi5hUp2NrVeil52r8+8rkmk6Q9jqAfQ09iQmnHtHWXS6FpP
Mm4R5SpJBB75X3IyN+prSgAbdAXEUg5ee0jd5/ZOQhVMwusQXZOCZs9hi6dk
24CxcG2sLRhGxvOcX78QvDNmgUsNS7U4mjJUZoJk8ZQf4fOT056C9FPEN24c
CdHb1emWInEr2oF9BaYF/6KeWjSVclvM8VvUXtOUzWTTLYvZS+W/WkwQwhFX
rr1WErt5j9GkxGP69KHCaYlNdgol2sbfNWLrjaLxNWK5HKEa1brYvF96eWwc
islWM7WwgOs+xjeKJhyKbYIHRxzg9pnXwKZnKk8bHSjKKgjzDHqQvKq93bKw
YLoL8zcxZLjFccz9+EQh3YCYuaP7qCCNp6D9TJQt3mFDyAipKDqBD+WdyRGu
sxEAHvzZik6A/zNMxa9mSoFxvw+g+O3Irl93QSqSX/rb9U0ArB4lg99FEwmI
iYA2ootROu/zAPUeRj+Yg1Ows9NhX17FJrkKmCDrCXh/TsghFZQEmZFqQ95N
JkC0jkuslk0jqqo8rpjPlVCvHu/HZuRMkJRI3Czw14+mKfXBOzFpahZV8orK
UrkQNnp4qHPtOrM47WBgLuWSntH+euTUQ/vA5xe8FT2Se8V3CoXtkl6NEWQD
chvzx6amMbcaQTM66HeK6QLnWYYMQppEqYW0cYHeDg309ttw1UO2PCiTf9dg
Y0i6OXbNUAsgqnGxP+rkNvohJdkEXpSqav1eyFt10KVVSER39q9qlyL4XOQc
Fy7jNKQH3gIcWpwKfKhXwOgfNYBO1koAhhrLwafIuywNvCI9xEgchnhx+e15
WYZk+Uoab6Cx1HiWHmSp8iXwcSKA6NIGfuIeziNSJGvmh/Msf09+HjStHoTx
ev+drz7541hMBhL45QrtI1B1nE9vYX7PAQF17pcdGkpU205xRYGdFN1efdYP
Nb36v5zDLpNhC//fLzKL3cLG2xQYRgHJLvWvfJjj7q4VNPXOEaEcEVR7OpKT
xfiEtbO18xtqeCiwyOiTNa+Ljj3WikuMVc+X6vY9ZODXGFr6imCAa2e+TjLc
jDMeFitnqmQpmZuQ2nyyDyNZ2+gKGcioiHzv76GoRi7AOyJnyXUBOb1JPbOx
MBUhdNKEiypkcS28gdmhamsBagCkFCtIEQWEYfvaxHYrmgkwoIZtdfmGVywU
5TaGLxnDYBwKMEC2EKGXDlIqNF4OVI4ntYhf5bSPpy00cYje9PW2hIjCeJj/
mcZ/fGxwWgRjfcNmECUihpeeklFxYxxAXCcATNTFEgGAMNVQtRaZe2+V8Rwo
MZQiZMf3uVyI5N3glUaZDKzXEFHWs/t7pwRIjJssVOz50GTBKQCI+AYFyKMo
dUCzAslo4Oq/421UM/Z4Nve6G5RndOCd5pTQSoTznSGdr86vi8LuZM9QT6Vu
CYsIqVhSKlVZUAWpFSbrRatX+zEcMhjkj3qHU3EH7b/Zd91YwlnutuYERh4O
zUxSMs87r87zaICmx//8TJxg5M/V/aOzx21UHjqbMW6UfHPeH+djUlrpDg/C
kXjAJnsjzlNtYX9Or812gr5IRRVUJFplEyrrztLgWAXmtfMOE0uXmhclpUs9
u5N5H0BZ3Rk3zKmyOYf+Gdk6KAfmw/Igb8FozcAvITctlfAVZ7oF5rcwcUuS
kSpFlCNsMvdUIFUVI3SY2fqFi/ohkKBoJjZ4iSvR4ZMS0whatz2fr5ctE4/u
/Tx/J/dRUzD24ggaZr2bbm4dV3B4tzGCBdmhLHFXB46PqE0cuiFgW6sXv7fY
uZ4HezKAh6H5d9LotXuY9LQKbgZFc+uV92+jw2/hsGpNenTw3QPTGFAKEnm/
kLkJ/lG0TCNLTQxVrymm5mctb/2TgwuTetpNBO0jcnyUeKRq7rMEPgaNYda5
snYIhDsiV0I0a1vVblkGX2AUTQYuFwBl+elOaHnnXOVU9BvzKIimmU9ciLP6
kzniBWObk4/fv/ULciqZv4stf6gzBerMA9bNPmmQ28Ol5UnK6uYSQDELYVor
28+3yyDDcDFr4UnY3uJT0MjRSLAj7Hzh+1MAZqVhABQAweQUuSgoj7TMz1Lb
idTQrjDyfMM8aRV2lDw3uR1OKgKAMipDSsFVUk4b2teeTkfRmDNkNWne+50+
PO2b3w8E9NOgsd1wMxSTH1aI2+vtwaFNWk7RavHenjqPasa2i4a/xJhXRUnh
RqOs6QU9rywMl2Bx/oYEXXMIKYbwOuHSHu/IHnPlSsAbvNXYOASPlD85K4Nl
G09XX8nuIbBLz34jKOZiSLVZZb24EpCrI/4ySmJJxAf7DRYDdH68SagbiouO
2qO7EBpqzm6HrvF362aMLvkLxGAbKw48uNmrUkUZChLqpqHFCgjfWv1Nvsth
fGQiec6J55XVLhs+OLGlq8TZbKp4NBIo+IcfBpEbAoH3iFAavBC2Bni3JmT1
dnvYcf8QB/zp9ZclUxqiyP8O5O5CrBjDjQg87QyIbmGwiDxDl1RNxCcuwFIe
bHlUbZWgVaPLDgee+gAhG9oVPT2RTdoo3Fz+kiDgTtQXLrj9e4hj8//exdgM
Zx4we4a6MTGL+oAXtQzZ9V/qyNw6JqQ7bGDsdiF077RrsMsflM0ybq3XUnIq
2xCaMV17RYzk/vtW0nQaUGWjdyQBLZ7nNKcW5LCwx/kJUGuSWW5lDZh0G11j
Yz04fYU6+2YRzdZ+rp/7AKwqxqhDhqG2JMIxQm4aXsb7pVpOHDfwWqnC9XJt
js5b264P5oRN57shX4pbLWVD6oSkRuKBlfrn85sDuwrSUS/UGohgMAY2VIEf
tq220xIYQdwpVHY7j+52DfezNJ1pBLQkcaouals8/W0DUCwpTl6m6m2+86fG
pWPU+oZyQMvUqA5u7dV89MJz6RZid9AMJt+jRSArYg2MJ+eI7nBxWq3lHfmo
1U9haoasoDS/RSOohpHC3ovmybSoGNV0BlfrBhybb94Sei/srw5SpPe+N7VE
i6v0zFpx3TvnJ0d8xgn5mlXoLewnoRPGa/yR7bvYiRfSlcCoBJnQLjcn4ZR8
inW5sVJVD5Q06vELTu8WQ+HYhDqhBXTJCJ+LKazCZtG8R4tdxcC4qXNBvhdz
ONuVgatkmzYzA87iBG2Rs61v3fcdFJIA/SjJCJpsYjNm0Gob2nunnyiOQAg8
WV/pXorpyHpJUwldt4kuGuHUuHE7x0TvwNQArhwKssfselNOXaP0CDfiYEis
EZTq3UwUbKNJVBCh/7hTVIUIVtxSHxMUhSgC+jzZ2548GCxgqocCYFAM0b8g
XB5DKE87ricy4a+ehPQgjkf51PqtgFoBGRK6UZRLPje/q+7aHbmnfxwIyLSS
2STTaV0tYm5kTnBrcLRfuPv4WrnQ0MFeG0InQA2ZJKe4ylijRxA6PhJgoZiW
SjJld7wUgY6KUtRnpHpGBK5/9Rqd1VRkmw9D6pMn/+IjV8khv35+YPjHDGC/
54LwiQhkJn/f83xtmnxuWts/AA16qw83xm4103HjZ7iVlmzkBfIDCeJAI6jm
jNEZJAJJeDfm72z531liMzyGyGNOHdd4mmUQMtyHRKbUGv/2sHNXPSCq8phY
jnVgG8w2fpRavWe5E8hZg5emGt8SMw3s2AVjfIlGDtIfFQQq3tceDrKzpE6A
wdQa/AORnJQRKBV5Uws14T7TqmVe0DBJfenUm5uTa4ZSpNvlx6miyRSmIJwI
PVfeb5pjLAA+eOjMeA9WqM/vR8VAs1O5gFMBqbvLY75Lg9O8lCQXHgsnhvNy
aVMFwlCyNPSWeD3Y7esCZz6QufJD6lvUMAhxu5PqCAa18tIejC47cWed961c
NgJg7C8phR2TiK0yr8Cxt2p3lCYkryb/HA7r3hmBxMgJFxumw89ZTsbUV7UR
QGehJFXH6M6R1CS7vVtPX6WQ9Sxr2WdJXYqVcUFWh+in46PvheMCPeIXrH1x
1udMZrsm/ONseTtDfOXKCD9ostcLrznZt+4qSU/I6kABpuW88A5XBZnTwcga
v+qAzL+Vy/iS3sa4loiDn6j8DTAJ6k7AwSnkHEAjwwYdigUld2u9FoNcnp4C
UUANqXv9F3Dp6v4rkA8tTBfpXvMKKLTG03FHyfzBBbH02L3VvawJIEFKa889
uMj9TuxLgPwFgToKCSrp3TlXw7OGyPB9auQ9R4pEM+P17AMI+D+qnpDIIiDi
egRxgPTy8qNPqMTQE1Bbfre8t1MI9/71OPTXBRYvicvzeXCgb/aKY8SmCidj
YUZivGBRo7+wfpq07rcByPASYx1LDY+E/BUFPSE+Zw28z3aIx0oaLuaq84sZ
9LXviNkSriajCAlGpr9q93OGpEh/FgvIky29TKunpXB5/NhbvwLiULGQx8Ka
4adt+vBclaLfcxYE/Q2ktZE0HwGNebrXfpBI8fFcZE2dqUgH0RcSW8XVdX7h
dERQfe+DxQrdfx3iQ9nKFahBKoBeCxc/0/J+swwdhN3CYFV2dOKIXxcrDwDI
K2CnL98umZ770fe6ru7pfRHeKQnWI0SFdMAgQDwPBY63SiDF1ggfbcCtBBpJ
q5QOeMVYeihsUU8NLEw6p8dLiX49MyVCYik10IjHtHDweJYGbZkVfljTehdm
NDvvef8I6nLKAIYOElvN8BQObB7wrKvOG2B8/bBK2U/eHywMSysyReR6LTWC
lo/RwjMu0uifiiqZFN4F0o4ZGJQi211GwrRxinGfwzt//6cd9I2PhQ3845Xi
tMoXRcK4ZRDwQCMgn+JGoJ2rFdm2BU7KlzMtqgdGUnkz2HAtkaTqOk8FMDca
WbEFQh+3oN1qlWRQciFaPLmuwmXGfYaZEk70Aklng7kFsRdLVcknlhTKYuNn
4w/9unLJjvUfoMLi6vQa1RzIlXOlVHCTOzIIb23j7C+qc6JgjKHjWQ3GNa17
JZEqzaCuMrRy2hSAwZcRxnBe89CCpR8+GDN/bM6CdAgGd7u+mpw+0iyIRAac
yG5MkzzA5qMz8RgYSbVMnsAT45dbwEo8xkCJ3Ftioovq5QHRXKTgeu8xJx4o
sXUXw2VAJXRjjBU0kQsVL5OEO3aA+CgRFoT//8UnBLO3LV7ZOEPydOPAPHgx
tMbmdee5AbUqqGKZxUU1uVmXyH25R4LmpFY8AFBUJiIAnaC5cx2rg4zsKaHb
2+ZI9DKU/n+pN71r/GHX60QwEyNJ0o21VU2y0dlmnEKrXDBb7ex2t4WKHb4Y
eXCrAxfMBa9R2rRtRrMWETwlDhhciWb5nTK04e9XyH8+cLpdi8j1vRJwMNxW
aIEOqnUqUzHpCPZQEBu/pxDlLDsRGyNC/QfK/gXSWUxGxnFd4cd8YLbwuGST
VxRHFRUg6akhPX9aXnCvTAcD9OXRLNAlLnbvV7vMr+IOQ5tFk8K7J4WyzbiF
gTjmvuN7vTNSl5l6VgEHaodTan5/xlPkNe1IA0ooZuUZOQY4gpvXegbDltAM
U2c1LFUVTgT5NqW7n7ISFCyEhPlxydkqR1NY7UpjEhkNVLg+X68woBj/wFum
8lPIurIeVVSeKDCxFkYZRUsbNoxh/KV8DesOCftIvhKhfxRBfo5ik9aUuQw0
kmUGo628oDdZ6nDMuNSEWt6Le/d93Xeck4LZbmAkONmo0dijZb3XTwSLmMkS
UoAa9PIRiBNh0CoX4rvffEJVWqnzbfWbcAT6YGiNXqF9kwPrc1+0LB7rxTsU
zQ6sNEeSsTgxp69uS2TpzuYa1UzxRtW0dYDrPfZObEV8PMWFAJzsHiDJVX1w
vLM+LO/GhyiC03Tp+t/1dIenPPjlihKkcVBr1RBie08u/IxtYtZc5P2YZ9B4
AtR6AS8xGQBJuxmOCV3DtO5szbR9mz9yEDSsSGEjB4COXYD+oXAUs0HtrDli
fRTKiGEyqj65vHTqF74IpZYr7MerjYPp40rcCGwXKubvGyDRhQIKxQ5keRuW
WqGYNCq0funl7i2eYv4zf+EXQt5oiwV/eBGKnUVIHiwtflTn1l5oTA2mxb82
9IqKW4mIsy/3VQoY61LbhZ8MY4RDHJh4/ZIU+nnigA7pf5Y8P+Pz7/tOuoys
MtJT5xUDXCNagM5xD8QwsNbyuYAKXw+wE/q26WYDToWtVynXRhyEGVZZJI4K
yFlONuubnDG5KifScr99rxWm2Ri8j/2ZkO1VHI1WNM4D9bczZkPl58BJ2llx
NrVMOYyEruukCRF954YOaoJs10aBGCKuvOm6+iCT64y9IfziUWW7vRG6u7JF
/ap9xHV1dLlnhOVlHei3NPyu9rWOYaVxX1nfPfsu8XeYqQX/3cHFa0Q8Ogxw
zMDS+UC9dYxztaqnGDa5LNXIVpvY1w2mMSsOWogCtha2hyugpt4MIzbb5pe6
XLZSEE2TzfSDQum/E714vT2NPiwhiP+iuGCJVHVl/4C4HC9EfCTMlCZGIXMM
z7hJfColTu3wj6vvBWxjoZZaikwRwhthADtfV/2yCUfpKeSG3IpDBwLCi8uo
PnXyjWIUtutLNf2sm+AEnhjRctki8ODCQ6XXSFqSdl3xR/pwo3Ei0T3eyK9P
AwlNgeiR9YV3eyIJc5sl6AZoGfOrpfyyN1SbSdsAT8J9Y+8hV/GM2y+uxT7y
NhOb/zNp8OwMM9/VEqEQvHYaURRyqnZKHju8kfS20ywSpjZLKTy83pLZlGt2
oLI+Fp0HLk5oqcO8d7gzBFqqMPTjkbLgjr4I8uj01ZRCOYfY8lWl+xqDTIDv
TbGFieEXjI13XphLzZ/rM+vXMxMz6auwqZugIxwsTzNmd6JaI9jgmraoMwOt
EUghJFwDf7sC/Z8CEMmjyGOWFX9gr2PCI5oxhq1Mh5UDBDmypqJKLmiaSVZt
qtrNj+iv8w1vtIAqF1knwfxOacMhyiSE/BS1sV1fohDWx5kjQ1Md3Lc9E5Do
/aWesaLtFh1/HxmgARf9dtq/7xRuqNUp78dlTTvtikBYc9qZGtnXLR5hCQwu
vBPUm4hPQU+e2Nzf3pAX1YMBr8eLnZ2PQQGxBU1smxnZtcNC4OBv4tSfShrk
lIxeMDtxDYBYnPiIKihhHyFY+Rjo72wnq7Q3govpfWRzt0Y3tEymNU+SZnCU
GeMJMZEeHZ3puUnQcYz1IXfYaP+SnIjop7WqEWT74Hh5f67aXnmMmVV+ZIdl
253CxEElvkdyKqSY6jYvqYTRfHN+cQLTLwmxYDojFz0Z1w5mhaKoLVHVpWsM
YPoyZCGCykbYRmIbRynYWmB9QYFnY5HeBQMciAP8lJhcCUKIZCpF2RY8NMD5
gKfg8O8UIxtSdj6Qz9jnpTJbDkKaD0/jPtHGjMAoxvOoNnQhBsmuc9IrBzrB
y2aq+zH7OlGrdLxU4roRTsnBZ2rte3tG7ozCzpJ/e+BwZAvx9iw+Sb41SKi5
2khDKYNdbjZ4LyVIF4ZiPS46WTtkFN8UJ83EO2bmviGIshvLQCos3U+GZfT8
OiD+xisI1Rl7Xtsok77xKJKGoqETpRfBXDHDUcGBLISxHZlcWU7EpcIRlSUl
+JnsPkhiDBC4UwzY8jzShzQ40kSHMfj27TiOOIn6DEr58FY0zfCJk0EQ2sEA
aOLjzpCuu5Ifagng5LVEyvRycTi2kcS7RulMoKaO8NsNRkk+/Ml+Pop6kDKp
QQYpBZ1oR5lDidKlLyJ9y604QmcndEcE3n04THr5rhRiQ3u6Y+yIxU9hY1nj
zZkM1jWT5bx48Ovun0c0i0JrmzVAHeQrANVfh8MuUVXBDm8aEf+b0RLeRS1j
1ifl4br7vAYs/3Ut9vqW263hUGX/T6m4v0GPDMXYwjc+R1eikg5cvAAWl5Xw
j2isDgtnygUhKMvxojbOYfWjs+PQ9YGllrAIxpInrgxpQPAVCtLqh8L9NCBi
IupqNe1Pjs/Bp9UMOAiWzWVVv6YpGqjLHcmKCJiPNPZBAfdG1NvqdrWTpA+Z
b2iNCaHHzgHVP4txBv1g9QA67cR+hA3WI44cnAul6YitXt1uDdpyc0sxFVzo
ju4QDEwOISaqMKQVN0Z+N7ZO1ju9CTlWV3iLc5Ta07gLHinmwzOiRLuVcnMn
JdbtMM+vi9lZGnskIQfqwxWMEBAMDotP6QS8OB3LAKWMxZI0s3moMwwXbQ6K
5v9aqqv9OX5q6gN3Y2VlBoc2R3/EXJuLKzJfv63uki6MkNMYs4uqKR3ItOFk
knJTEXbKfAEAc1QTVfoG9Hd+rCViN92N2krVVYwlMp8Gmizu9qIHDwc3uqUZ
sYngOj7sixnHbHMN9Mfk5ekDLHw/Akq8CV/GAjq3ToWDZsIdF0B20/0BMoZ8
NKlomlQBEJdITdJyWQb32B75HOTRBYhIqAdxvF2XtXa7X0E+Ha0JhX8c7Nni
Viy779woqGtykOjTOqtN5dH1w9jQLT7cDuQhHz7QsTRyoL3QENQC9LuNnzpD
SZ+UOYXF5hz1ccym4JbIkFHXHE0xWF83c0qltF2MjxMqjYe5KmN6HPB9CT6Y
VkBT2O41GD/9WW+C+4tBeP8VsjUrME6qRxoWMZ+cMwwQpCrnIPyU4+CZpkmF
sNgtSA4lSvHkNwqCZfQ2CvYqIgif+/iTJ3o2qyr3TZqYFGF9shWF4DlCSSbo
6B2XHVnANpCCOweDFA5mkkH+6ecTbxQqR5NWyX3C8UxEMZJvtJJQBlhGbvPG
v8PDq1qo98D/xlmu3c4vdZ5kWdmPT/4gAPLNoSUmm4FuSndW2wlKXuhyOxsp
3Aq2HS2ptDDH/kYcOd1T/DyTdCDCHqxJ+Nm+zPCl9bHPzPU2hGNnO+O9QyFR
RKSkRFC+jmLeF2vMi4TBrhfKaR1aCpfm398Fpx8evTqgNeGFp/uUJZPhNQKX
yyKCMMWlmQu0Yr5ugQBS95qHJ/zRRpOaVrEFZXQK73+uF6yYU1aznkNshTRD
uYxOYzHBglYcKfC4/067MCIiJQfyNWIm70cRzCtP1e7BINROzdlJZJpOOjQL
wMrlIWsHty5jjJ44k4h9U1JKxNvW4kNPYYJ5ff/PrFmHyrLSxUquwD4c2zBd
tmb+tV6xnhD8Qb4IofJDh6n/uZV/XqrbLWd1u273P5TKq7u02zHWEeJEiKLz
vIEPQVCtMa3yrO8t0JUciTUv5Nqy+nC9asmjuyYJoKs080ACTmNrNdwhA0Vz
KLBv6oUABIpLb7tl09N40v7BJmM1JZSQLiQMF2fppW34+10ttTrmOI4F0ScQ
mvBkoaA5B5LnPBGOj2nnM8jhRvDH3tt0XK5fPn9r1CQy4gY/cV1onwUy1Uat
iRpzONSbaVcT3WPc84CYy6CtMA/GakY9yGZWS7HEQpUZNXV1guG8seMdDCZz
+uh+RLG5SHhT/7u2AXMd4kthBYeHF6H+yn9Ke6X/Qz0wRi3FexBtRudVc+QO
z0D5zTy2JltTZRpAW181uHsEMPHvyivcU3DvWw/MElaOeTtg/8aaXf/uuXgX
8VjST1zBY6TwS5vtP8DsmtzhTKzhIDoznTvGQX0d9bQKQnE5LdTDDUvao3pY
4/dTakyjUAVBRVPUfVITJKr9i22ZWSerCfeeJz8+xF54+7Xy5SVWeUbNv5m0
Wjyq2Ldwb+RlWJloE0xW1BBdb1d2Y00hT3TuTRhA37Fr9FKZCZdwcq4zw9DU
n5MscwD6/opUHi90Zs+DDOyh/fjEwu0px5CEFGQTEIIbWlXYEyGHWFnY84GM
FzT82jM9WUNC3KuEBoy2Tv3Bb/hmlSUZP9B3ERBick2egNIm60RL6oPuyJMB
40sY2D4pXHZrOihin0RS49JBsVC6nI4qsSPVRwjF9PitWPVWS2M3w3iU2Ybb
iIysPj7i/P/gEeU3hCF3REL1vBLB5OqhubL6EFcqHRvW20yHlSrKKHSsPTI9
eQg3NtBOEDhdjiyIbnpsOgVgZu5YOnMAgKwNuyuYKei86liD1g1ultBmRJZe
w6h8sVYXEmKMZ4MBvrHsStJPwb+g3ipVGmY7ZFTxWYGlEBbznawtdOB8BVyI
wKHNf3H71G0hHQLmWiC1s3/cgIFvWg5+rSDoXr7somK6ieXJJgHbEiIRqXJJ
j30caEJ9UpvNko6mCJIparoPdilyj7PSvKv46Ya0qq5CgLYvbirYDFSyy4kh
BCoiHSbai2qFPdeo7khl0CU7CMS0oawhKleduS+zClc2N6sfck8Ioyofzl2c
lYafLV7tYYq2aACDXrRxEKWoSMU4VXT7PmuuG4j4xCPtGTa9HI8kKBOWh9Zt
l9/saMDrb8fa6jsc0k7YWpJFOke9Wocl11/AFnOOBFibzukBgXjFsLelQK2t
zFyVAd70lF5zPcbjq3Ph8JV6o9x/E46lZmLgIVQMwPOLXZZMXu9Dw0R2PNiB
0Y0w5qFxtAVmHWsVDCCkVDRCr/VKtse5ivzZdatLQbXQHMUXqbZeiZEQYji4
tn4t+w6SXcXOxfJ4r6ROAS9f+KP4m9Lf/wlNLvt27rwgq/vvHBTwy6c+ZtFh
5SJkSTKjxI5sEZ2n/y5uUx5khpJ1o5dfnBM0EaxV9lsyqIGXLhp8EgBatklm
hGmdTw2L+NLwg4RXyfEzVul8jhgFNdmciBpIPTQRLiddR9Kz9VC7LGPBhxJf
sXJ+6Rk9BGv720Ra06PP37iC66g7mdvH+LWT8utkeD2/Zt7G5NFddidGUPVQ
PBUP8NMiEEYW9t3h9PkJ6sb3rUQE7o+EQLrzmmFfalun5ZGQyMt4PW2DgpeE
1B5AVPaa5R8B7SAcWo63OWTiQeZ6cP72R1KIuh3jr+KMHc9yAEbKKcB8xRE5
VC8tmMOOYYsc7cOilRY/HjzreH6CCa6jZ7+2szYd+K4w2Vfh7Mbx0SESx6DW
IAtb0fgVB4BLylZOl0gPHrr6aTdofQOfJ6TUGbLH44uvI0bZk1/xv7e9jBZl
Cb8binNdK2ZFS0iOSaknErWPnlXXm8M9nRXyW4vQUFp1u62Lup7eEcB4PNee
ZnoOf/c+MLBA5sUf5ZDKS+2xXEoQcpCQ8i4VT5AanSsrVFf0PGZeGnPNY9Uv
NAGMUGUlkLag6JwHaulRbPUrj87BYnWyAxRShKqqcv/J3gJO21p+H2g1SxCt
3mMTlDNuoUDRCU/zH5RJwEhg/+cjrz5k+iOVHY/V46vwI851Z6bSEFxo3lR9
0NvCVx83ZkNOjISgS6K8JI7vkouBMg+FopVoz88WJjkErBOacEAGfPWZsZ+a
lQMY14xZEe3Chj1cVmzWo3THG9bR9LO0u9jBBtgPjcbMDFneAoVXBGvx0yJy
q4HSI++nZdrjAw/vkyETS4+3N+bFMtMTXLuFkTyfSTLFnXu5EUYw936sUhcF
LZJgv1gJ3D0vEub8O0A3MPUlbHgPAmT3BPs88+ynfMkApCawOjfrh9dRIGHw
2Gk5/WDf+SFUuXSt/S+3weLCrnXc5eSAd+2jfdbFE6EUJzqtQ9sQ/6g41o2B
8u8/oKharDf9q1SKSHPa7ly/Y5irg9kzVOPutoMYoXgWZXuN6iS7xaCuv/wp
Wd0cDT/RioN7hC3kRZkFEhx7DJNJw9ZRri9E+DXQxHKmL8kFKedVgZXqAP/t
7/LV++yorBQKUQ93vFV7k8fj5DAaErVvQ2pQUlLIPOwvuvokjEJzbpbwVLwu
E2W8m5sA/E+cIYQfXpeaqW9RAAdl4PDM4YE1SJex6VabOqM5WhIWKd/z8YyO
AFp8qblZy1QFfFI+34R78b2cu0/5DEwlH24l7aQLXdioy2MhNm9uIawP0smk
+WGO83ilSo9RiPdxB1AUU2aXlfnfUxHGs9Bcgu1q6cv190pHYfocaToMDrjc
ifWZgn54LnVhFru/6y57sNkpXemaCWw3nIx2TfmaSCy3FUfKj/ZB0gu/e9Ms
KPCLSGN0pwWrPlGaMOI6Fvxb1vDWNlkVhutCDoLc7u990QvWfnUu8vclkZnq
8t0fOIhJjCGzkdfBmjVOh+eFkRwRRZWIJ/E/V5cvkxeZGodXqar7ZniupQcE
t/USL2v6XidO8ABHHBNtfh1cPbQ9UWgDu0kwCOjKHhpAcLp7NRjs5CagRg3t
m80l/orhJMyhesDi5r+JMwMMNFjq+W9xmWH7JD/b+fzObYWzl2MtIigor5nG
vETivcvA602ZxS3exxmOZ+sOUkLjmLbfHbiPHiJzmLzrOYIFifyOO4SVL7gV
UawU6YvPcd5qWj0pSAPgi3gBORqKjTp7KJBCm0zKmAZRfpmjdT9oQB5BXfA1
9A3mmhwUo48Qam/55llStfxoaDSNGEAzXZn28TdbVS+XFqNZx8kJDDtE69/5
pa8pg0qM1fcsRf3Lgpgsg62tCItxjMZoCK6iF0G/4fcBHJFqQK/cUKAOAvZo
oASyNRnG/HXXUxLKBj7dQ0ofzotnd6r/LA2WdI2WF5sdFgl88chl3cezXDnz
mtj05+nISUksKIQJhVX3a3+oKH6BgT3blKi6aVF+q8q1ekP7VMgvF0I+Fr8u
CWH8JPVOBTVYzrqgqU7ko/bhDTN7MVzKyF8fE2wQ+u/Q41EtWAQjLRonvDYq
v99TuCzXIEYzgiqg00Y9S9fdaTMfLro9anWLh6tbaeHfPvIElWvodJSx9Ecv
qE6GYLtWJHW514p0cx6eyJBpfB1Up0bowqcEN+u2KV7AGM3oVImBUMFeyW+l
xcA9cBNObWw7aTSUxnpacv94Fw+Q78KHeItitrZ6S1Vt7jewrVHangMetCJf
wFqtjY+80XWqn4ydGkR97JCG29Kr8uUr1X4O1mcAgdbZvMCFqH+7V17TPk4q
+xI5icEU3sP7gGYSB14CmXjupE3RXYXxDOZ6SPL5s77/83+qPdAC8IL9miby
NwqUZ0OnfIXGlmCcspL4F0KzZBx3/OCl3IkSkUPLmDpe2hbEHAeKscCkgpmx
LTg5Ytm1VJm5NHYdFqcg3gZwjC4Xx7vJ7QB0KEWfimxAyCfi1j2H+5J592Vx
Ic8npK1BzT1r16QQv9DLBeceDcOllx8kUzoTP/RCilp4AX7km5rC1Z1DoiWw
RKnlHon+SVtMY7mR1SKc7dvxU9uF38KeIQm/hu8n4p9Y6Eh/GSmJhKizfF5e
3yCqlJOAjvYIhqYUvoynFekrd2TeDPcN7CzhiBihjsu/CXd9E3U4BijtAZFf
XjByuRBdxkAjnU+aIGtuo3463Gl5BP2A3/TGFZ8B3XOCI9NztX4yvj5Ezv46
toqDitkKJBhjOGj+i/BR5/nEd20fIVx92+g/Q7MloXY4tOfvdijT6uy2jVus
hqY04/nx6xWC8ifYyRqSh4ZAohudSad2SJWh2G+BcE23zzj3taM+29Bwbd/3
5P0xtBq3MNze0bUDP5lCueZw8uPherz7sOKdVoiAlGVajw8oV8RedVL1i6Ke
piG8R36yMBo+tDBL5yfsGTN0hL+nYoOySXVRARcNd9cmJfh169k7+7RC8/H+
4TnJ8G/0acvXg17V6JwGQXkbO3Oip9nJTFRJRAGJPwcEohxm5qRTmNYyvzkR
+eofvfVXTnT0IUgNTjUMf3JWgarICcBle1ygRwI9xa8nng5fLWY9HzuqtDNc
GCUvnAASgE6Rss//xXk4c16CrYmUE2nLo8YddhX+a0e2ppoI8Nq4xyQqlKtI
VrLHl+WrQQlVtezLTkbZXdpspJ0NMO/z2CWortx2jsUeCVxb4Js5yC6SP/Zd
6Q13Jd1rD8FcN9yIyDy/r1BclaTsE35U0J75+Gj8pzDi9fTnaAavGi62Pw8x
pFMo+JlmcrmlTZMIFI8Aym8M3ruVYyVSYjLAMmgvGK0XJFbpSQYmzVxdz7sZ
S8fobLA0CaSPS4KytuWjOYVWicZPUB1PKJbR2GXHcLTkwkISPzoJt1Mez0Zq
zm3RFxFwDFC9t36VFVNRcEy9ZbiAY/dAIuO5vGA24kzRSWI0XKPlkfMdzZqI
hQ4gIj35HCrDO9CxGszhWQxFI/bTBVnYMZrc81qGsQyBwSuLcNhf4JIjbxHr
N1sX/n33tS80MqNuQxUYgK6J9LdZJLmo/41pKneEzpmKo82fnB5K701x3IJ5
kcTkANMj5B6F4ekeOKnK+OhsUjQoDsjQISxJiXUe0cfqnMr76+f1nbbnyR6J
q8j4hvR/5/vbWhttBm/oroeTxWvRhS/0vL3i4e55qGOzKBsPgaNFcF3zj3jn
r55l58cLviqcDxWNwqgWRdgFFxcxcwAe6mAnr26CIh+3KdMjW0hqdQ/c4Gni
upyN15Hr17aQWEhu+N/KT7c6kOSzCo3xGCDCHhtRbCXT6WYl0A8MWZWde3n+
SXszZ9ElkWnqIf2rBGpnrTxKGkOHZiPXd/BbI+naqpjosK5/e4Z2ZQJEDGxz
+TAcqhWVRFsqgOcXxU8D6igUQCh1o2X/SCwu5QSfHygX5R/MuB/n8mLB7wRX
ExdaXtd3lp2jBhXKKsarMQH9//p/S+2uCqDLpzaIe0mxCiNeXwFDIHRGM/1j
1wAkZaTtjTMMmXmVwvRlorSOXv0i/zk9LYdM+6u1ujiXFsoNlZ/nzN2Ed8VX
NlBQEztQepUwcHbw4UPWb/uCEgfdBuaEPscMJGwrZmZhtL/VODU3A0TE706j
xLpzm3OuxSHvRw87jyitviNpeCgBDi3xwYUdLlCu7t4ldUnfBxQwhVYwJe94
2BpmSmN2Kp+oZAkR6eBmjNbZieG3lw0MZZ3J6ONwKL3HZ6b59eL9zJhcvdxW
C0E8VWuC8uVC7SIcEF4tpXXOq0ZLqqzJodBu2r27xYf8mpolIfnPkgvwl6Wr
xSsTvzXVvi+9Cbt01HtkrRlUR1NfdQco1cORC+Thze0diIPEjUjMmW0k1IQu
eQ1sugJWEHTmziCTyNkeb0n3RgY3q75Sqv0bHiN0ClpfGVyy48SHLtLEpzWQ
0vr7rl1EctNbydK3jMsdplw+rgKgt8SvuiSmy4Ri5ifHSGljt2VTU4lJVmmC
ftVo8YIrlechOJd8MaAcQ/PbrswZlM50fWQVrORFxj3dJ/fQ+5gxJd0k/UR+
MFDZhY0SthJiHZIGDtLpf1iSjTP59i4A6k2bn3A5ATr4vVhelKelzmnW0452
QjUSLz53l0YpBlIRhasKc5XxH23GheD6vu+hrou3gXzkF6UjyHNdk7XBau40
NTtUUHbK7bEyTHIly4Syy5E+uW0khXytB98N6bAIdZc4USSd0egejly4/oQe
GA6Zc/lTIwhsjDEsCz062yeUGVIXKpCcjee7IDhtyhvaQlBs+auzSA+dJsTb
JFHAdbjWPdqql67VUnQt81G7rMB7RVgjP/7eV4ack/fjz3KPEjnf57ryw6wl
zcm/a8Jo1zUe4v2oFpf4SouBUAq2SYwlLHepL3O46rMQC1OXX+qT0yu9mWlJ
kzfcoMCbBooxkJFXdmm3FurnSooyiIEP++ewzP3k3+CV/zt9BftnQi4LO8ZN
QDZBHLt2VplyYQVQ/BK4McbgyTuhxd22XSQtd4FV5dfxP3EMEbFmq7NK4yNn
7ZpNFreeiMDucbCStlvMmHXBWKq57/WtjCYk8C+w1HRfN0mJN7xnc6i4lAWZ
fEkOsKVqclUo45IJx2D05GZP/ywOgDgA8lWweATIo0LKfGwpXHPZE2g/SGdO
Jp0RyLxdhdyf+nJQ8XVxtDYYDA2hYwNqYZ8v+Y+CbvOYQJ25kk1QGszS4jdt
3z3R552Vd30tqRFptywmhvNftFF7cpSyEawyq23++cCBedZ+bl++89W2h8cs
sv7V/Kmz7jarkw5pJRVZpfXncrcqJzji5EoK1/Qv7KxEl5pljpvM+1rR1pye
BrOZOzch/UdVPeTFtj+5rfe1Ka474KPa2MKvTgER/OoRK3mo2aCL58csxTSQ
nvfhuaGVLltiotED6oxCmFqI7mjl1MptvtsP1MjuLVzC/DLIqQKLCDI6J0of
0mDtGraaYUaYcnd3ALLPlzrvXkGICM6wqaGzlfrjoO1oUktdkPnfWHhhdvX+
J2VS+tyU8nUfJIgKtKfH+UMQZmBSvWU+z32DGIdBcQVCGLWzkT2kYekolTdm
+o34xHI3fGssDunsQR1yydxYg+ju8ZYecj/8ZJOF2A8Arvcx7RqLx4XBJoS1
0dI7YDthaB0anashoe3TcHjPQ0MFZqDhvjKZH7Nufb2iowUZbhzl+yUVWn5B
VyM5IraEn6PYsR/p57SKClOG2N7YHBfyruc1cfxtfD+gLEIWHMq0D1DVtDU2
DILu7XrciNU7RJvNrpb7cI+NOgFKNCQyQrHujBy03WB1u+GcPwGA1TVL0tg2
6KzLod/VLWDGc6iAYVaojglARs6ihNLxyB5m4svK2p4b8cU89SKVSsAPh9aP
Wzi3/5l0m0gQkZqvkOf6E5N6rZ+tKOTmB2o3bOzuDLBzQ1sHeGqZFwlh/B3C
T3ot7rF7ySoUtps9XkONdZXNlQrrpcTGBRbibHlqlUTodH4uSyZlqBRfXTCZ
ra/KW+uza5ZMmWnlW3U2b5bvSPc+csHE0CZ9x4qKhl6dJyJvF7E4gGgKDZlW
rnQ0Cq19ufDbyguMsgphJa6NsPMl0UtQ+8GX4joS1IFluVnSLXb3+kJiuVSX
t2qBs0/Cdiy+NP5gZq+sy9+9t1CqaXF/VhArWjj9Ztt4BX/2K6+ea5AhRyDk
0X9FpBe4tyNNH+xJWzPKbqoGHMAFCedQr/4Ev9KNGnPk7W5tFNX0qn+HygHH
UcYVuczT1Md3PJ4ui8vGOuFlZifHpubIW95I0SDxmi6mM123pk53iat0Udzm
GnH44KAV7aXGd29iY67W3JUq+iM6eeLc1UapaVhkXqpBmxmo3qRL45cJ/FUg
cfw05IRb56Nb/u+UchSjkdEAYPKWbODwK0Us0WYHkqyqIb60sdWMyOSJozA3
Ld6oyyyZX0eqNpRziw2/kRVeur2/EmuJ0KrUumx7rQ7nDx6/1WNrYRFAdu3w
w88/1xlwQLUgrSWjMeE/w/cSebGIs7NfnoEDJzYaCUM+76a6ThbepmH45YAV
QNBGIsYZTOpY0VB/O0DS5SVkAnyrfRnoffzn999sKP0dFtH4Y3bV8481OiRa
dsEiyTEGpQoKW8QU/O+QqZO2DoEpy6XfEPpqfhPh2Gfm0YgcZ5a1V6/1QyH2
Bu0bSlPSdvBTBYyDRUxjwQx2lMoAmHZR2gZjcrpEECVjRXvxNQYDWF1fuATy
j4U5Xz86NrbLpznCLbbUf85iPebBM1lVUgtoVRurQkh+uqYdOEfjngBsjIUb
8fOvfc1JO0XRnUywy15EkOeJwZKmFQoPEj+SKbI1nxGpsQXiLVq4ywtINzJf
rULop6MNZi72fvoJmEvn5jj8l+dSiMQ0oQ8u0ZHda9JyN9Q4HNGQnxYRL3sp
zebYh02o/IIxbyN/HkLXufh2oYbY60GkY+RWQgHcJlaYchAlnnFWWt4GKrmY
7k29p+gd9uLWI3TQF6ckrkexCO+LbXKSX0X6JtJYS78Igrflw/WDaLeTudsg
BiNYimkvvBMdBwsM9gnw6FLSIw/fMnCrBXBmltrsEkqR8fIqk6oak4BRuvhW
7lQJtlUl5PVcHGktjWR/lMb3v0brT4c6jsqcZFotoaxJ04TanPuOBUenVr9c
1px5yinTwl/b6bu6jMPa5EM8U480CmO9DSD1XqqRO95TDUpqItIMlzO16HGx
CEem7BW1KkGTc9ftiOXUYwNAvQj6uWT5yVDB/7NZ0mLYd2Yb8MyA1EuwemSF
LmC0bdBrE/cU6qI3XI0g9kBqC2AeCy2C78Gr7EdeMIVGo1BL8u7eEWgZNg9T
QWbntivIkH0+tV5fQn22MJMAVDUxKTLoy9QcMQSkjpQ7JBNfNRG0iZsrStT6
hoA8rGtSe+pQmwceqf7CRspbsuL/VMPvbGiyY6s7O1fGxe/yPe0tK11RHefl
3YV+PR61xpG9jjO1fo8P7WikIhWwIHL/WqjMdweegEMs040kHPthyT8ACQvn
ohz07GcuCut7W59t4WeDmd4KtHx2/6V1ERi+sbNxeKTWTYq0fdkvIfqbtJqu
SYP9pKQbXDk5+GGeVh2oURZqD5OunTP4grmAKT34KHsLNDOJ06Oykfs/cmRG
IxyrUKAsf55bfLSWqTBi5F39y9pOO5O5i6ys2WYPR1G+igF1f0J+Y9CerCfF
4cj83U63zoTtOIVrRT6c6YAr/xRg9/8Eh9bKJ34FADRpPnlLfsG/cQChR3ZD
1lb6NehjbOZeRG/n5sVatfQqTnmGxiZZUuaYeaoJW2ggOiOY7dF9Kx/giPLa
YVN1X7JLlajzA9wK/3nzhATfeWoBgCVDecnMaGxJEyl49ZkG8OEqgb+gPWCt
udic4Dph40DtoxGfev38RKhL04Wjx28n6WB8KkpxVM2snlTv/9zOELE7OIIM
9ZPgh1jpawB9osKkH/ttcXlvxumYM34oLBAMiDyje4B0ktDs+HxNPEChFL5Y
hJR6GdOta++o5aWMP+mRgLOEc8rSLBNnQuzBtmmkHsx1igOBGq7rnq2qk68X
S9pQBaHkEhUhAxlJCtuFdiCqtJngIRu8X5AhwIyf2kXzcFenGoe+/QquMQx3
VSswz28mnrRTlFWVZz2t/mLytYarJj0HgFVCgXaLSvKV/80SinpbBhrep60W
Lp3uFGXKXf56qxBtXKZtvr0WhKp/fNZhTx/Tf2FoTo7zctq65Snw/jFSZJym
Ly4V3lJbRCfoySjZzXUH/7kDuN5/s1icbYL0FxV71pAkwbJGMGL1ESXiUIMc
Si8Tav97tPBBAx1BN2fcoJMFf45GLQWx4DCpOsbAmN3mtsMrH6or6URsVzbn
8nq+4nByJX4XAM70hykFlMY139aY/ANNrR3bAVF2r0OsHar4IvwwF5cURDo1
0lgajDDiJes92mmpc6yxP6HoauNqVWtf7E94ai5FyonFmJUWGlau+Ph7gQ7C
VBLUm7bXCDP0Ul8bQlczcB03fw1yWmAA+VZT/f7WErGK3na7KlovQlMIi3zP
NWpSyr8ZDkfmenlhkBINC1lV9jH/bSt7cWIl1DUY9lpSZFvy44JxGmlJVgw5
fXD46oelz2X/PJV1XsHK8DKJmRupi2QXGDeWeMMYR2kRKJmxuNvD5EQaPLYD
uuC1VSu6KW2wvQGGgIs2DiWn54v/3jIhb/CvQ4XqK/ips843bGGsq3Gxq5PB
TIgDUz5KyvBNQ4Z8RnwddXqX2/6+xS6RxiBIe4kjqL9A2B2BjV9EkRjh6Quw
0HVr6YpwZmZD+b7OyGzM9wbOevSkkUmDN0flVPJKkxIw+NW6ZZu9UFlObDTo
RgxRp9zb+0QkETrhM7LE7eEEaTUhazWsss2UjJoMT6R4DAqJ76C3EVZ9jXFn
81iS1DjcbKK/yGfeDO9TCWK2zg+987gLn0MZYlxiHnIeJ3ff9OrGfNWR5Al+
ISBn28kxKfOjphQkzd8VdRlfqzo1uyBANT3HGnv7NMkQ9uEfWyzPKNUpxzuK
6jLF6iGL98wuv4PTNIcCjE3GNwsarLoJJMnWyjGkttutzKn5sE7tnI6Yi7EU
iFiXcZdbDZTnr51q1vWJljY3PvPYLyix2nXAPr4gOrSRYZRtDizEj0XH2kZU
azwgdtnpG9RuVNwaLEwrFQCz2OVKSUhfHrag7l32l+u9FpcQKxpPbEJ+8ySl
si4aCKBG96YbWrl6oWWM3b6eTzEAEvpMPFOlWHayOWrpmrnZyKIE8Ak4GQrh
QDBkYlxMI+5Wm0oa4qTCcCo4hBI1OK8ruh4TltVhA/bfoxqubvjv93R3LZRw
puJanf7P4D053lE5GkSiZYXsSTHU8o69m8pud8leOrldJxhRTKbwf8KG8AgN
oc1Ih5QIsoW6dNMs6lwgWbz8hcFQrMWsGQc9lVjpEVkUE0PNmocFEpJoaMXO
PtEW1PVR1B6EK1s7Q5kxA0muBsYeCOuFr+EhrqRJ/ET1ZD+Y6QizsliMe+uD
r63f6jJdwqYGKiQtk3AmLOiPnyx6+KoGw6tva/+IVbSam1s2ZwQsRes4CjhE
b7fidTsa1WVNI3xvzPYIrjII+AbLm58OMsoA6WZCyZbfX3AT3ntYhWvOp4rd
b8ctWlnQXwngAi1bdIjy+zZML23q08R8BSFOjsiEgTp2KvlPszQuNp3/Ntd2
Cfp1iFOv1MQ+WBiu5wXUlWBfxj3kOD73GK8wup8z3TSI7pTkHxZTNbbGJx89
Sbd61/b+3L20RoiUQ0foxLPsmIZa4TWWmTNBsLhoBwv/VuODinR473iyhFUA
JuT2H+RFySr4w0r1kqKGO5XFd5npdOCuJ8NhX/w8dX2hNWxknYmvUyk2ckTR
kEaUKrvUs8cd5QTXno/v0lshZhToObriiqAV0acqSpAQ4FTkOKZy6MGusW/a
aYBeQY/JianH1Hd1Iy1Gt2E+F5bl4sHECc1Q7DD2WQxCCv4JcFsFiQl/2HV+
4Rt9/dweDz+J4CfrBN/tjwznyAvypyR9Y4aa3hjfHgpxDcgwJ0zLQhUvPItp
X1bPWokITN8bgsEzdgjxO2pNwv2Xe09fxvClifPwatvetlveAlAnLT6fL3Kv
jIrb/4FYXqgZdZX1vcEwsyZMNdgJ3aKU3bfeZINjk5R6THzJUFnPoxxsxPPe
FHOBuTxzpRjWaOtXdT73PhLnapR5iceGGkNZ4iW93e7EgTwdm4F0wm85fehj
sQ5Dfk4RAIMeqUU7eZeYZ+K5gqvRKqU5DuMDfT5EUtBWUv1GJK7B+wixg2Wn
QmvVgtVi8VciyGoACgcFfN8tnc1ax1C0kImHRnAFB6xgeDLG3JxC6cKzavzu
SRO9VVUrIVN9avMKMLrmD2WGcuWEEJpfiYvUtZycTvvWvtTPnQl5FKQMVfoK
21f3rMCz5tX3YIH57KETabg+YnhXRKJmd2Iu5hpblFORjA5/HeOdq1m6GhQc
cJERr5/xtJ8rDC5jFMg/ayO07USgLVyS//+e43Dkmci+RyORnl9Oy0LEnoTk
QhLCmKtcG2Mk+rTnUusNdhfcAi2iM8l3d4zLuGaFbGrm+19m0dsONo9u7NMX
EPL42LQze+ZHqxY7IlCOl3v+LsRgvsGnLqBTs3KNQRlgk3O0T+XphFUuVQ1W
2e2saVRmp+a7Ld9K3PPLpsziuJ54fNLvUX5vO6v3pddG1rrJ0q5oDLz4c7vO
6GY4EQ6SVSyvhrKOlEkJLGh8GNm7rOlSo8hUllmZJniGRyGzHNUIjpwWJvJR
/J4dvyol53Xo/3dT8w9mfFLOzRAoXlubS3ox1dZVO13w2CTCkISPACmAbcUv
+cIXUVkD5ofeIao6wn3QkT7vYLEgumxl48UO7WhXbzVX39s9ORSPE5CZ3Oi5
QGuGw9wLEB4v7JKYOdOHX+Hd0C6pEBNSRmk9YvcdGLK7T1Ux0c/FQowRx+RG
01/1/xtbaKGeOXwDgzN7NvSHd+KnuYNMAMO3w3xbHr6PPAg9HVimoN5EBDJC
oy4cBpFOqCSk3iuwAgdjv+OWUCMdElqGKbugD/r8S9ZdUKqGd4DAX1U8iRiA
xRAWU0fkfMhEkhATw9ufuL2Hb5J0Pyn3Vl3h302RZc3+OKavcmthiu41vXxz
JN+sHlhOggi1yd3h5GegzIQ9lh4oen4iGHBKGOk4ut9NyGS38/aLLbDp1Azm
6DS9NFhDncbpwhre1vnosYAxFL4vo75tkyGU1PVOIvKrBOVSEGE/QeDZnsh7
XUT+DXHYJalSdn68jUcytlEkeH2/zK1tM0bzaKqOPQZ+qjcaYhbqQ6VvTOM0
Ty+jajDHNu50Ce8cTlqMrJXVGyQnKW/4EUP73eLWC2pydS6ZKLv+GDI9ymU0
ky8k/GJYeEi+cf1+HokhjfNCbuTYnr4cUMV7MmteEQBsYk1XWINrg/TR+qAy
Qibh3xJl2e824ib7O2KK9Odr2JsttSr/L9H80zNn4Hzval+gBjwsO0sgRCXS
o3u+UJ7FQff9Qfw3Jfaz+IfomgVpv5cMLLJZmK/00TJmTDAiR+IZK+DhMDJb
m6vWpX6GduVlxYacgC7EfSIHjKeTT/GxkCpGe/iZSWLCVakrIy9BPNHF6meX
J6a+sDfNmw8IqgDsjDaCHTqDyp0Ha61eL4GdN+wR3xX3dPFROUAlWpJpqvDd
AHs4TQKImom1Jm8gl0OrcRbtMojwYaJYprdbEXpQ4T5iY/4iqGm9XSqAWGz2
plAuTo4Dd2FCxIVAAGZeRwjV1yY8LL9mY9gwBcC6jDiHHsJlJdnEzvIB3szT
J7qk1kI6hD1A7GHvSvSj6iDwQGV3ocmGD//gec48WJVIVALt8N/g04oTUuTg
VIu9HavDvbZgJHdpwcbvjqXgKinTq1z5yCG9/uJqSxmSkqJWA0uvP6Rg3OYd
Y5jVa1ajhw0xbcYJC/6xXqAP3NzIHwLgaAabhQd0hsoo7BGI1zvaGP/K6fBk
8n5sgfBUxsY0WZlKUnt7cyLMb7/UCojraCNAg3JO6dD4OioRq6JRvAFfCS9s
fvW0uPTf8b45o5Sxi3c6p+14ZomxWfpeTIT/laFlnis0Ne2onpCpInrkpZDS
2+LOG6qC9Dj6576Byzx4+4ZIf4vQyEXa8jl42ZWHrdQ4RsdpWaDxBg+RbtN7
A1H7HXP5CJhj2CujdjPF49IRMKe7PWwsT57NqjUa3UYmvneaBPQM04YZDNIO
IlYYwp0pYc09ZStyptAKVAGQEcrkiSOdkNX6xPGyBqmiwL56oKZnevTJD11W
ZprdT/lMdxxQaQDdOEyMbjGGAthKxkSUHF3HP31dTvqIuUOi3QGLQez4COfv
9gWaDA+zmHGZ72H8qThPMYodQjQF7kHnhuUXVko7wATXq3Nq5ypYNIht1vQn
7EO6XxZhMpMrQebvsGRfhMDG57M1qaV29WBPUjxggU93CJJ2vZzTJAlFC2/z
Zsk6r0EnnaKb0+ys2A5WbPLBjcNtTcB56E3pRhf97QMG1UGu9aaEeYHd426O
c2eVzzHo4NZhF4CXsnsN1x3kzIM7scwvfbPsfwBbf/e0Rpx0aiK76HW7vCn3
XrKfB5ZsFni+WuHQedyiUTZptz0VophZdeE1fg9GG9QMEb1LLOaCWH7iURz+
DVpS/nHGt6LFLdKK4hbLxi4axAQYs1a32BULMWLW2IKVGxCO+mwcsMU59GR8
brHvj0yaBgonTWbD3hN6rLO7O2TIRsoW87FDdsrpzuQAMvq8HS7SAZhf6H99
F8sPZmF9+Ji42sdD72t6iMWBaHoep3EqdWUgTAhQhGOG0yEORiq5jBvLj/a8
f31+j7eWOuo2+o7uJy3VlzdipDSCzj1aGlQbqL1ixNTDFS5sfuVW9oSqRRad
vdS8M41DBPq9OJktudOE/XhtD5daE8uxOd8iNKiOHZMldv+Yki8IGYv0BkpI
KD1DIoluTt+wSpgckycDzsfCfpzmGdnnox9E37/2zGiTuPn1fgF2dgfIxSeb
WGq0926u7UOEXm9K5e6aHHCrzTwYTExPe1sbga0NLSIy0lsfdZr4nwP/IQyi
5pSfsfitDKIXJQcQEKMCg1bbamQ6wuZkmaGYF067Km+JKBbiePtUCJBrQM+d
6+PvXe8PNmPyv37bbWpmYQtVG3pP+3kjLQPhCKPNub+o7Jgry/Oov7T+Mhnt
twxsIx0RXqYhTB+hpcqipLTXeseuIqKhNus/DaU0i+nOR/2lAzpU7MVuUE4K
ai9gpS9FaDezh4Vf6wR04YpItgZoWhkLSHmxDEfJGK/TOHTXeiPQ6fHvLMjS
1ZFsL1xL5Zhx/2UoLz+V/+dx+b3UnQrPXdUSlOX7KdTE5j+Sr/Bn8wYplZ3W
3x//cKnoOqKIngR5Jy4BuDrlQp8MyXwFsEFqffweWXZciQd9t2ckzGv4pNCC
+kmfvR9b8uEofEklhQFCgibc/aOJvqnBFkxtFlB6/J4XKYjKuons347bT0Mh
rs5Lmwx7l9HUFOiETZY1TkgHhHjHqyBktJlQGv0fligrcFMZwuSwv9KJ7TnS
JtszEFvraeNAJEURae/E/w2OPzkPVPV0k8RD8h+jgYLc03Bqz/mhBGec4B7J
HrP3vklj9HVQhohqt00Cd+x5ZNup3DBhD5CuE6EF8RXxPvQC9dWohdOgC7Mg
zrI69YSXPOB3ydGwWliEHf0rfSfczSlMZiG4bUCRUMwEQIV/iBtgplbp4vnn
cP40f7CiCELfCtNsBVO2kSNLwMYwH2fa8AbQxn3u7FTU+Rnh875wV13/DS8w
MuzcAcI3Mp1fAMvZkIJYyzsiFczIkeSvY9NurgNviva5UciiTLsb4AjK4c5E
Ap9TtHXhJnKv3jqykZ/Spxc9qXAjY28sb5t3Xfk18dISiDqYUIKefmdzRhii
VthmoWUk78/DlmmZA9QvhDyq4VqS6QVFJm/iEOcjSCeOH57Y7MbuDRTy+yh1
Y1vlit2HxHcGTUwI2c8JJ9qA0aIY6WXAaaVn4OvpFwURm/cFptLZWhwSmPjU
k+UgbhZCCbWB0K014rLPSwUAf9MCTc8BDyHl03aqqDWtk4saScndQant8w60
HYLYaMaudhRkmBNpsDGeKr+vEdeRDo5472jo9JOCI+lI+sGXj+Vq7b1jsxxv
GbTvrqY4k/UaJIeq0PZeFgODT2AblH3wn+3h2V3qfTlvtFODNF7ak/NVb3PW
pqCFfR2D8yr6wE2rYhUfqI+AfLY5UJ3LVUBJdSso4GXJOaGn/4Cx76G3Fjw6
hb0J4B30OkoYzgAQe1iBWfsTadUrBYQGEL8+JrY5z7I+Ag5ulgcvZ09gYP/n
f/DNX31mIaOBTOxlauw0ipm1U/yHzPFrC/pIHibTRlcTjQEqeT+PilTztBW1
cDGqX2g4C+mQpNV9Az0pbNvJFpAG9YQl1CaMD2TYykE78PqqKNnUuWk9DTzt
2/Ls6SeaROyKMdnheoBueq0SsfUSlM5kbHE88jn122UdJ8u3LtxC2TxtIhxd
mUJeDARljdkqrGwgUZbDHJ00ll94hU6aqgh04gFvDHsE1jArfl98V+3fzDIb
0L962ePxgPO0k2e5HR07HsvFSOvM5++7nhzQ9ag7UfxcIoDXfaJwyq4ILJW4
Ywk8/EYRzX5ONtUiZOAlwfeEfuNJhQDCBVMy5NJPI9UESgwHqGkEsHrg/f5E
fyeuSzINSfyjtqba6u9Zy8yDf+2OnmyvFqJ5jo12pfeDvi8QHfgv701Qis1V
4hy2tqwjlx2FThsWm5qTnoA74VjT6zrAda0DY+yVj+wSBJmzBtZBWUZHU2hy
CYBT0IVTeroYlDWABJq1tQvKqo+d1cwYw2MBLhmpRibpL6zoifg3zazPe9JT
OHgwARotLlB5KJ8Labo2+jPKBKEu8Iqhd0dqwFHdC0lIeoiDesymKG1Ng9jN
EFGce94kD9m4SLXiYNzfm8YsdtllN4M297QbUAaAiuHTwF979vaJLwYt21CO
j9ZjmQBHgnSXzsjBtdATIwahnDjKGGrwUkvnHj/P5dYhrh1LVZYC+X5zkH6r
HEa9UT8keX3S38+MocK1Ll+9trl4yYTqd/fAmMPuCSS9/Oq59EMKNEYDryse
OMeakAh24AIMrTTJXs3mkqZQ9asRiOV5HKEJsCi/V/r42LIRW/G9QOn+HVuk
0ybNOPyZoJS5dG4+29HZyTfZNJDMeIoyb0Amtl55W8nJye6FzwGLzOj8ZbVf
0Va2bSl41h+IS8qyC+ft4BcYCU4sa/8IY37DanCTAS15rSZwskBE0sqxBZ0o
uK7Wb1OneB2T+hCbavJbxcJooOepl9vRkRgcyPnmc+oLjI6Cuh9b/wAbsPfZ
vE3afP1vY0MqyW8gu5SQ+KLoLp/Sf+0Su0g1t57L1S3MdXZDn29qaZ6w8vDB
dChQVKlot9wKnjf5522dvZW3mzd2lZG8ajJlP6iWWllRFu/wsBFmGrPzh/MK
UkB/NI9d6PJVZBCaecJJyLFwp9Qo2B1WqPxKK2+BftkR8+k2O/l7B/TYUSDd
Be9VKPr4bh9hdP083x3LQeR9sde/GY/p/7nsG3ji0dHZOK3uzYcwfjoEgOBO
l4a+3nKO7FGUhMwXxg8rzPknJ03mYlve5oyY/u43woyqFfa1E6ffYU1vlMr8
pn3zz9gqP7Lcmd9ei7nIycMj6vF9vIlt9whKltgTxO1xkz/DbEjoUTGklNOJ
wM6VFV6m6P5kZUK5t/TcYMh77G5ENr/w+q2So/SAes3LTEt0V3ZEqYcwoZK0
0pPFtrWsOhU44FRF/gNsYeNb58U1at0seJHwipskbGfwDXpP4DECtSNEPghK
/FOsFFz5am7jn56ImFlwSQIOI7+isUOmht7p8GVbbZDufi/r2WNbjMHU6NlY
wX7Tk4O71XZ1d2SyfnfFq9Z8oSAq8uMvTEacob+EpiLG9YGVR8UqfUXjv5x8
SlEBb8eEc7N49btCgzZBXZDS/4h5G2egwt8mN7KVlbPdjJBvO10yisriLRP6
mKTmU6BHZdXboVTzdQIaYlFsexChiagB7leEnWtDFkBm18LXKkF/opTZzBu1
aZG4jK6No7E5Y0e7BtZ8dei4V0zOowbEeBPWSc2Nd4Q9avs/q9FbjdDfA0Rx
xMozAvQJMXUlEMRx76+kOopnSuPZrtsXSdt4Z48/csUZSyynPu4Szs+TLjcT
+skJn7SVsZPOMDkxbLbuybNM3aCDFT0NLGS2nfirFVfT7FtAjgIkgj43GuEz
fWSUxVhkcNNKA8k1+2AmgukzIwlgWUnWXuhkop6zkmSrv37/1ekHhcwNOj+6
UWplRTT7InOISa6Q3HxIKd9qR/wMa/+6SGqiCIT7m4ayqLjA7lOtWqKK3/fz
oYLQbCJ1d2gl0K432X1fVWP2o9T39XYIL/VtbFLPrPlBCzWDmkl6EhAtCQ1W
zjcM/ixWe2ncsp8ig6xOn50/wcviN/JldF9LaN9nnDo8xBjR1ycm2yTyBboz
UWBog+ayctzYfL16nw4wdYmUJx+yjgC9SJpSSCNPnzCxxKarb7LVamy1142h
9j5hiY8PNasSouyD1Gi1jl4MdjEduMk3cCri0Gtn+0Y3Lr/e3njq2ulgNoB2
mXYlQLgZiIFwokvnMwx1Uj+oTjOjaausxytDGR6avAmBe39ghz+NkIC0o2z+
+jnla5LatfbWjmV0syZ9bUJxEb6MqHaAmkGLX+EXhLrLgMcn2uOd2tkwqTgZ
/RkULu4LXgCdBQyhNbjtuVBR0Za97bqTPjTQsdGvPXik4b4mw40RsOZgqWqP
BxkPRGpD9FLIbN/3WsmmZ/tOnHhvf8+WOKd2rTLSa/vpCtF+QY28AdjjBoLE
Kw6vY9fJwP+xVuUxWVMFM1X3It7rfOtGzMlmwd4eNGOXLy+kJCSV+N8c9u+4
dOgVDyCIhxoJnAbZ8LiAM2hY4fVMfjEuuGWkDREjGFKwscCR+8qD5J4yu0C5
7QkfyY4hy0sQFTrI/eotFzYIRBrbpme54TCUAfvgYcVPgfOFyrkNl10bCVsO
5uiGZ32t3ag/kYZqCQ7lG+g9openA84wkKfuXc139VP08OQuRjoQFFaBppGn
Hvt0Jpxdf52x/oRzLfA0cY5d4f5JuR2Ay2wUpSKDFEbIcIKh1DFSCEGAbBCi
1ojyWIhpkgH03N6gIXpdnsLMCSXRYyf5UC3CQg1NWTcfqoauGNw/Uc+t3YsG
NTi9LNcUEBgLpKY+mvyynMaAyALeT0Bn8/78xualV2MbPIDt4NXYXU5yaN1F
MoEn8TgJDYPVMtwO9h07x3+sb7eUVpDUgtvI2kSFsxhLZb5WT6YqX6Xk+6ja
OOg4okRUw9qCVsSXtL9OKd6YSY7gTf1vdBuhKnlnNbzCHCee6fzerMCgM0Rr
qjRJjgrlkOghIWAtjO0io/xVk5U00OtLKF9oxe/LHg6z3UxsuoA09TRgoZci
J9SQt9P8qh/Jrf9k5G2HVJpW7RQQPmwHC/Wy4upxtfhAaECLzPNpUvxt2CRh
UFnRfWh2bDATLPVBR2fKs7y7uI4Go+ypYND/0ZjSKrjHndowBEedYP0OOmDH
7q0zLgS6b7V1IhF95txIxGPpwYKmxNKgodaO6wX59Ve8VcPq5VnyUdjj/Qoh
x2SQQ8dr/+YpBEBsEpzA1NZpMK+YWGH9Wz9I4iHRKIY12xpEvptA7pcYpXlh
M6VYINvuAI2M7lPPSwlvONc3WqJFwagO1k1V8VvzKyUsjv9NYfOuk4fxVyPc
OU6wjauG3xUha/2IBJOE4+Y3DTxZQBshY87T7c1u/YEZVe8yVOw0xJx1l3k+
XiMwF/3GP+oOMk2nMSB0upJPxbbHkJMqJz0R1gPBj/KCVVdDAhGfItSavPst
WF6cbuxfTCIjmxj4yjgGLNFqbVe6WYZcqJsuEXlW8rg4+6/fEviYh4z9Qj78
nJ6D7RgfD1gUWpN+A7Xksz+GOoOqvLtJobXoWi4ubSU7s/cURb69XVquz9A9
nitYfses0wF0GZ/uXtZ99EO789l6s1MuOnFaUhmug5zGunBM9jTNU6+qo8q7
m5pf0upjKP6w4k9AUUYKCwo/hRWRyTE7caX5yw6WmM9UopPVjVy2j88qGn6+
/3FPTNPSVWmn/EOT0Kga9RAkuDpEhMmmHJ6Yob4OQyCP9LME1woqNq1s07fP
vEg+2UmCC8RLYgrIIKkYhCKH5ofnDEBXpnHvP1unpKSjrKuFj2MsxGuxeMtK
iQMMT17zdoO/ZAL3QP63KzPIXHQyUR7u4rHksHXrSvepTtT9YWUM9KP+m28P
XndmquYYiOjDkzDpPjJN8Usd+E0k07Swce+YQ5DnRxss7MNlz+WTffyCqg0K
y1jod8DWOSt1ErwC1gQX087ivIsToOAY6pdfQzZo3BBkga/JjpZK4n+Tx5yw
i5PdGCZ3sKde1Etq10v+FG5fnYY/pwJdSVJ1FRc0NnejYASHTAaYtyMzfbEo
oomoxzGvD3eN6ys/5TSZFfx5lqL/nBSGmN/PEMiBhaT76DvSF85cYtWitYjI
8kgHrhxiqmBQIX3ZiocF09w+EbY3osOSuqSCdFrwh6P9TgeZb6waThVdlmm8
RqYqvnNy0Ya939S4DwAJnLOHOU5EzMJyQ5nCJcYy1c6CWL4GZnEnisUmFItJ
/gmPGGkipcvKUPjIZPxn02x61/wqtVusq3w0xfZf4r6vXSLQrwEfgwtuKLJd
kfD3NzE3b8Tba4TR/ZR6mF9/qmbAbStsVTbwDpEyL0vydHLKwscgdu9TxTkP
UOf1ptZJOOUeORjA8Y/3iLloSFsX5O4/S3qP2LpdzI5rQiJtYSTdX/tc7w1A
quQGDogTpuTyVvgNAXhf/tETUTo4+2LD0es1K98wOVJeQbYhysosxGM4CI0x
KreRbjV1hSKoHsie/NAgp2Cg8oIvtMtP2rgx8SmtxSktSbDv2/L+EXyv/rdK
ACm0ei118A8PHHDLki+Qnsbnko3FHug6OxEUeloxse0jeaPNKbMoXdm8tEF8
khpCQX6B60I38NL1VEia2/NI4YdR2vQgLl0L/VzzXC0Ov/e/ck4FYFhhi/Dp
tH60SwKO0ZzQTz+jhGE5xPqaalh7wB4YdVReMo6a+AnkOZ3Cs2VeHo0MO8KM
Q3/kXfGK/ixZoFZWmxfSSrT6HVsbHeeLnURBZxfE+mDhrDzcxaLuPCWLNfae
Q7yve952AZkgL7OZQcNLALbtc3ngRzD7plkzAGnWcGbFOAmH+Py6MbcfEc71
BQ0hLp81UTfhec/Sy7oxU2WWhwcAP65bgC2tS9+zZUrG+OKUpLnU/XY9EWol
ILwPNBz+805nU2+yoagQPzmEq9amE4rjjWAO8YI6Y6PpDMRy9KimrYnExQt9
tOqUKgCkRVTz0n/7dKqS+4spknK/JoFs07YkhriiNeTQ0mrkczrT8O1ALR7r
PyV8oVSTrMEajewZSjFjDADOtnkI8m3RVWKHehmW8H6oK/wlKpdJ4Rji7kxn
n+3kuqeFuubPep3e7ucZx+PXx16IofGgfZ/ZSY7FmMNSOwuK1Je+Lix74KFV
1z2qttTFTg+pLynDQ00obDjo3BJ0irTvWlpF0X013mGOXXxAv0fMZzMiA065
LKwvlsJUdZEr6d12eqVhFk7EqB6Y/sBgGAfFfUdKuVnDIbwGGu9BVgUPEAuo
zcyvMPjG7BX5aBaj5M69hdcogXD9ONFwSzd/lR5VLPJ7D+TxM9Yvi9V6GTNG
3cpv/ykmNSlzZDLKjOYEcNkzs+6hNVsVDpJmFB/txJ7pD7xDF7l54XNMRdeE
j+V5G87xFgshTP7+a+ESddeRvFgFjEqkD0R7BGjs4dSCUGi2iPxRcfcDIp7h
tseFmOKMcKWUgmVXdVF5s5aWNx/NIsEnqpkWpyXXe6ZQ9EMiOujvf2KXyG5P
eotCnpZMd9jJ6YblVwhr+jgqJTYCslEW9sHpYzvyvumJGZxKJItWVIU1w6DY
UJ6cT9lh1aWYdKTFQTzWYAY1EaK1Ic5Tm9EbTgRiXQMLhzDL5GhyLwlGqqSg
yCZZq9hChKxw0WsXSCN1eaYMhfNCeandQvHDRAHneNXbmx0/D2qO4/7hAdkT
fL0Jlo4PG6uQvk1yZk4G2z2DMakJSAI6HlgoOss7diDjMaes1ZFtjZ1RUvKW
KXpy0y2JBrMUHmSwNG90bHGzDY+rkO5guzYMCLL3EsaK6NGC3rT96p5TE+Bu
/PI/f/z9K+LGNBTwWxiXEbESkk+Pf2mWTbgVp9UVoGdoAvTxiXPyXcGwMPY2
EJVMvPAcpwFZzXsESFj7HS8fCbUoGvllgdEA6EaDx0yOYL2r9QnMSl2XZxCA
2j9jWAv943ioAbqrWJ421E1QDCqfDI2tMK59Sr7UjqX6WRVx1VsKWVN2gbl+
JN0Exje8G/1pW1gBGFBJhF3DOWlcpBbM8evJLu8p/kmYCk+QNGl5oK5iWyxV
6xjJX3cWaGbdPLxvgyS2zX8ni1dNzzdtyG+XTwD2fOVMakvwZG7Jd2lwd1OV
1TH+bEeBLK3atR5VaB3Ft9aGW3qCXgs6rEH/G5MCMh8HecJ5ItcZ6BmFP9lJ
Y455X0utoCkCDzKlhTpzpemlv0Mo/mLyOK2a2HEwXVX6RUs9YTJpgr1iiazw
zYSituTDAP1yA1acVG9Kw99wEbZu3nrNd40LYYEPuLEvlxyUu4z9dc4T0AJM
rdmardPpjfJdmlD075yNWQZ+nQ2BaPN+e5Ie5jYIjFmDzZNVwjzVkNoVsl3h
WIkQ1uowrMZjznhpUQwph3b7CyYaJ3exfUZUaHrFijZ+rSIWeIrAIi7o3jHS
SaPLZOnfV2sTJeKOGyAKobshKezdBXxCMGYijabEUqbnSOsg/P8tXkirfqfV
304CV0Y+OcmfB09MHwGGv0xxbnpjvK+5V+z7oxbiuFQr+1zmAnVEkz4R9c7i
Zd6mx0gwn2GltZW66HApy2cexemblrEa6SctjwkwWqlnpVg/4BUTiHl0vajX
CV6C7PiE8WVCcPBuDU0FpN0D4bJYc2dFK/lvqJC4Va2Ww3gPCtX7Szpu/sin
fPWmjCTN37AjpRphyFSXF9xf2ew8dUqAps7QMG7TAXxeYmT+dMSi2FwMLMea
Cfy9WgbqyHkxwKZopDqsBNUGTIWmCtJf0bHcLa1yjYvznA7WCXTJBPFe4zDx
omg9FtmRGUQ3BCsTmSgyczdAsVCg/7gSI0NKMYPKnamDee/92XOR5Oe/sMS3
Xj6hJHuIivviJxMnkByTPSA6p5YTsAOvm4nDFLy4CYqc3GVgPr3BZN28FbPK
sPE/QCl5XbAVGIjH3XulIUjUNNxP931OVhsnKgZihEkfJ5rO2Xj1ADbgjzoC
8LFGqmXh+2WhhUS9QTMh1BJfkVQ+aNNtPJZy79Hi5mNgs4xrmUZ34/r/DNgQ
8ducrzOlsR/Ao/QJ39NP8WlUAXGaHyBROJKFmdcGxhnr4ZVC2i8UMIrMFUES
y397aUTH7hq3PXt31riXcyp/GpLYE9DAZPDzWENYraXCMvYYcr3d5YZOaP/H
1JfkDpt75OOyjOGDMPMLP2EkWneftr1VB3UjiD8pp/UM0bz7GRRA7IQlFwZb
breX5sL8RZkr3/Y5I1mnUnhzLWRhEn5mP7M4tTuA0dWUic4mSBlNZ8qnmwPf
9lbb7v3e8VBTOZYPazwpD7eqTefWMAUhehQlsppgtNjwaGVrMuRDx10SJ3dp
nh11V1ozLHazGRbZBaKFOmUQYkbA20k+B4dOmWQFYH8BH6s13YDzyOFV/s3v
pRZYf6Yfm1RZQaFdIEJrToHWFUfp+vxw025sEL7ZGsiNZ7gGFbEyEzlBUKMi
+mTehrRiKJvzPUf/bh5PcBk/1OnL142B0mkcsfU8W5g9ZPP8caZmlwi8wS9X
xfzt4bR1edQ3VRNW9rjSLHqeMN1D66sEV5mGQbgFd8EXGZxKRM1P5jdpiq/8
kV8jnnVl9n3TLfcd8wcK4BiWNdd2Z+XW2BNlmXR5gxf2JyKpIBD8aIf59d5J
4sdN/6FEiF5rw+ryU8IgGGue6Ai6mWyx8ZJ/iT9sN9abZVc43Ox1wg6GxasZ
MtB8VCrwvq+92URLmlD7zHjOmsvaNdzHfiZ1CVefJjFMD01biTrsjrfqp3al
T4sz129p3mOShL5hyU1qZZ0ot4Q8jwnX3SVYRLWN4TlD+N+VKgh9Uw9dTJqs
kwDbAe0h4uTgrNZUU0TzjTl31Rdy58OTs1Bl/XouHk2IyYVH7kHS6yQJsk7Y
wfSgkKaUNkHGS213nWrAY29HUUALEKnxZ+w45a3+G2reTy6CRaBhONCwPFlf
dpp2H1uKj8EacKOE62chmfsuiONGZiCIuCXkgr2un2TyMN1iGTcY7gekYRbC
lXOP8tz6sz+pnOgog49DadQBQWmnO2LQQBsacGg9lagMIzT1NfN7aXI7nWku
3tuxgvGzmS3tOaUUKypCO8Whu6arjxGow0VZlwzcob/sBgtGXyCQe720CCSF
CW6DewIdT/+lYRDlRoesYEhmCsGSQt8hArv+u7jvz898/L8Om9OmV3zNvneu
uKB56awK4zHlNXBpImCMlEl1+r6kI1sAUMxyeLv/EaG5czPmuKdw4KuHAzh+
MaRI2i6LdZbtYYkclLfi1SN86G7R/AQfoPixQskQ7c7HzaEqqBnfRUpU6moi
DualeExdMadFh3598vNfW/upmzW2KItY1GxOXsVZ1WB6bd97wFT8eWxjKPUu
s/Ytdb9bCeCP2Vuc8h9p5GcLE83L7LOxNOIdSUvj/dlffisDyvEPCm+SF9Zb
1Kkd0MG/KyIvx1s2k4QQhucl9ieM0cWBJLmCcvJ2neN/gOdmsEjChDh4RNHI
VUZdzj/GrnRSPllCwgq6fECLJqpdxtNqkb8oEDC2hpMwaq5jtmpOykbYsMgx
iNXYb5OPfcw29QcOVdYRo/68RBdKojPxr/ut1fVRvTCNGCM0ULR6dV9sIdN/
6U8Hu7tB4MLPId/k0EG60XlHNGshMPeGclsJyvc+h1quI47kWR4sm7sImgc0
DUs0PdFcTH+ppPbgVwMBpNPrM0YGMORDCHo8ih+sOyXn+2UAc97aR+iztOoO
WLRZDb8dqOipNBOZbN/VSfxV2hKtvxt5YYMrPnl51hxhWS6h9MaiWfTqCTVz
pcIP68FyC2SvC5RkkVcyTIpNDoc6KxsR9an6TCIiwNc3NRDUK9yVuz7HzaPb
s6DrcLP+Gfisw4HT+TshFUxvkm4uBz96HOLkG7kKjWwkg1P1l5ybuIvF6alQ
pXBB3PwaSKaUOIrcUj04ObUwiEqYoFvfqMYSV93UJJZ3z2yeS0UYYxYA/FWq
/TOGr2IgSzJtr7l6fRnRcZzTk1804WSDQwTFeDYIQwipgS3IYAwppLIbJtTe
aE/nhmjk4WBZfRqNTPXnUvPOcn02uzPfbl5Id19YFqCKQHWPfCv+At2BjG4l
6QAdf1tIFAoZTHH/QNLRREhAeznP6b6/kIcNsPOdaOoMvlrqm+h/PFJouAvF
5vlKJShjxlLTetPzvnkMPjBR7UAFtdxRAfnkEtsC7ff41clxucQhtwHcEPIB
09srSQ1wnfGu7h4ENRea9JW4aSJSrxqXNs1yS+juflcUhGYa5zVFgKYY9UGa
CnAAQz1vjTCwij78jHN6+LTY+WBLPFNOeDVLuYWzrFqrOMDlhlUrbZKLbFOz
pZvbV5YmVUntnfvw3j3ZF0Zd3cjah3y7ZMClVJ+TH0E0akMIz/gGD/KZe0rz
YyCKArGI57Stugb0dlBTG+6hT417dNpzrpdcwDP/IBwy/Pm3vT8sdtbQW7zc
m83C41Z8cPQeneAeiJI5OKE+q9WOaMnwiM8iTReiGYWko8qtZuS29QyRj5Ds
mtGkpSoEPoRs2RVHzxueixxCJMyWJOJv6elhvw0ymAxpg8irAZG610FTZxK5
GFMJCWqdNZcsOAF3zzSCO07iZbEEqzN7xKTmKpeUAiW6cLlbhVtY13ZF/iaF
DIWPiTddaPgy812DFHktwokblB966Fkmp/+9wg9UyfjaQrqK6tEsgeDkgZZ7
XBrUy5jwgp3iEaRbKj8QQQfPdVehNW5h8PQmF3WpEVl9wSvx7p9e4tcsLsJJ
sdVmTv8LsHw5cnyEV2RAKl8gvDN919OuEWV1F9aP9FeNhW4QBaDqhWUCfWr8
rUlbCbngCLhTlqaqlJ6w5zdnO1uoQ3S+obSujt+jmnTiNCdAxe1VGeQvGDJ/
H+UA7DDpzvonA7uwXtxBNAqoqYqaM5hsw5MZsaGCdUzujizUf9ZHWeTQfWRV
1Hp8llFWukxjHPASnW78TcIf4UU1dXlXcMf/tKRtJCPFSgcn9ME0AWFNlClp
3szCBPAXlx79lN4AkgZn3PTo5au7XJRW1sqRFsnKR4s5ccbUOpb9JIQ8XfzE
YKKe07OZbR03lKw7stv5tj+tHT6lGjWi1ICMSjynaghnP9NmdBJEOkbitGiZ
wrtARvMaffhOWyE+9zl2+HLNcDmggG4lbgktqlM2i55p/Ah25U1koFWl3thu
H7S7oo4nF4/vS3wcn72UdkOi54qumGJ0TprRWvGSh2Lb8dFeTEJvLQgcVNAI
/cs6Tv/pa9jmZmJXjVH67jFiuD6ZyzNqBj3/5DRkIo0IHdnTkz8in4PTFikI
/9WELC3IBNQr/bV2q4g2TFNXQZiIkSQv+Mup7iz6Xfbf4bTJ+MKkZ+wTvaOh
sDHRUsjD9Ppdo7E7r5nqTAGfFlJJt6kztS/I2gsSvRMPbYiEUwda0bKEoUqR
cCKwH/sn3Vzs1FhhZhikIQfxKpBRpACgL3mJeCEck8VEKzQmiTNra78E7PvV
qZJuBRhItHV6n45ZM/mLqhObldFll1HeKZy7T1SRK8yNfdrD7BR+DwPto8vx
QBp7QdX7+U6KYtsd8CN1Msg8apg0OTw7IXBfpnFRtcV5QgVWEdS+Cj2I/Hlv
ZqZ27goJPmuY0YnlAQCKq8KN7vTbiYDXhrWpJXZ9xrrCkTKw0gTk0nlwHVvq
uAKrtOa3sDlojxuZKLqpBkuxONHsxbugVp/44Z0E9T1r/nRQLQNAqNarR1gV
7UArwz9TlWQfYntQ6gum4UYwQIQIOPMsH3bnc1KFHWyUGpZazjiL8sQ6stnW
BbvGlmw8GuW7rV95rMlpLghOKlqRY9s95IpzKKvNH+RcMGOLC1ao0+cm0PnR
dYy5iZ269EcIfk+OzpCMTwMvL/9mQOUtYAWvb7/Uh6o+tORVh9qZYuHtkrqf
kxag5d1BuMkX7iJ4tnsW14Lx88EeEVSsHnfTjlUgyFXkHqhRV+9wpqe3ZDMK
44m4DP4GnYgslX3imda5OPHOJ+ZmrQlbU+85wtxcv8Q9FWpk7o0kGfobAvs9
JLpAQV9Qxy9rLlhTeyv683MIgunR2h6ZXo7yddodaXZheAmh4ofEqk/IEzZG
oHPYtn7QHZyoyji4SNoYI2AXFQTMdTZGOG7mK8JVCFiCc6LfRtLE9oVF/wW0
RV0qu3au3xvT2y5UV9S5PL4ZnDD6u1DazzuoRCaShUle+5Aqv0i73fbSQKcy
RosuOEyhqsMMDxp2FFymizES65F7t0W0+IaGWGcKwh85/b2ndCB0VjHXvqth
57OPBtqjW0chR2uJOS69O8l/hcJCguFGk26TF4nTdxYoNNG/XkhexrZYjwt0
8la4TDP8eGrILntqnqrxJnRaWz2Jnh6PkqIfT/hw/u/ceQZXKVb7wfqwph0S
QoQTM/gv3T+M3JqlLmmvlqeUlknfOVinXZneXi7fTxgep7vBa3VxbXbROlVI
5WsJEzaNNz2y/Zh+cvdkjF5iKuVRVOlnIZCy1VzWNpQ6BNlt4sSHgWNq7Kep
NKEEbQ5/0+i5//TIeqt1tgj1q7fgvuImcbxpQq2q2qO0dtVALluQK5SMmISF
QgMBhzP5ipNa8WvdDgQmhn+Cfy062Lfli8Lsh/Q3lZk8F/AAK8ABzhHnjKSN
WJYjw6xciKvKG6mcw+4UaCW8xih69CNmg/5Dyjth86osQFsuv6PznFc1HltW
3SNACe4+P2K21SE7aJ7DNzk/iiwU/vJVFsp9KJpPZimB2TAzyx3g166FEus0
KOeauiRb3SwkEBPCFPE2y9O/Ij19nNnXlz5l3Igixv1VeT7LRtLGIDVCgZPW
MLClB5lmVAbVFNcYEzIqc+AIqLPTjA1ni+oGu/xa9Om6FYgGRkjBqvTy6euC
edLWQXeQvXU5/A5sPcwUloc7Z3Vo8I/pRtLyUB7E20ItnkdWBJzZ7CDjuIFQ
bRxyDvwtnzT15O7s1luTmR856LqCocdqYRcPCs6E2JJ37dIVcI6bXJ2ISVl1
7Rta2diEa61RmoYAbIlm5HM/aIoxiPlDO7Ey8CqwY8H1y7jv0MWjWREVdEm9
tJF+E6UHMJOF6r/W1zEPasYa49k+Gk1lWXF8wUq8YxYTDG2hHazN+1wpcU6I
8Dd3Eicp/8ECfO3XV+1fuoAnqqwRSRNYG3MNBDqz6KOEzaJXTgyqnkuv6lIt
lmrKe1TLmSJiXrpcOkAZtVoO0Uym2bm2ShmLNaxBVyTyQ191f6dw+SihOtaK
wtaLrWF43CVJtgInWR/JeV17fjuIjcN8By6eO8Bh6a7hwWN6oG4zgUGzErau
BfXF8C1YBuIoADLotagpM1gmR0SkZzUC3vxZcHWjiBZD5wD86I6F8wBSK/Dm
GLQBFMXuGO3dFOniFZQrcwdkttOsL7mnU1nJARgRJov5YgbBiOlmcZ89FjdH
rf1D+KNLOU7uGRaN5m67x5E5MsLYDPIrmMAXfWtst6TRTD7x8kXYCZUza4UZ
4oxFk6IIFdJnUzHpwAsUWqtdpDtmSY/IbzA6iFwy+z/5mpWxr7DXGrlLpN1r
C2tXnlc5J0RQkRxnZmRrKfy9gJF5BNs1ckMb5scWdI9KEkQhcejrr1tM5zOE
jIHArE9SLxmCt/BsALq6AWN+wFAxH+qSkWq/5upmejqfroha7m7CDOkqSpGi
aqGha4pVMbL+IV2SUCOIzC2sJ8tjvqqQWcNGsmtn7zoSSIc7OVPMwCYisc7v
mSNRqcyLb+GnqGlwDFGb+0eecDbJPI3qbYNkaWoGJ064T1Kka6Cp7lec+MSw
GCqPgOP8lSFJ+1G04B9Prg2kDAEfS0IocBlmJtBXl/AquYbu0MouBITMykko
0SW8l5Jkij5R312dRaYqhK/YNdQQTh4g1LFWA+mgysOrysp/+tpST+Q/Us2p
EC8+7EJzM72tm5BjJ70/NpX1MEGICrEmzdwkl4k2ssfuNoeDhXXBQou0/Rmm
7xobbihqc/ANF2vHOpRoppaW+eHdHq771E9hanh2lufEHwWbb8VMMdpY705u
4OJyCxLU2dirww5LYqEa96RKDKR3/LN8KR4nkGPu7NhFKqme9B+zew3HgUqM
rVskCf+p89I4dR42PZd8Jai6VmslxG9d4I07QzmG9OjKWBZF/cL65giq7vhT
PYutv26XS/0AP972rpZVT9/YoJea89qoc5AXqEftF3m4JUH9oDCg/nvmZK4f
F3lTVI+46+m9JRTFGkVkMc5ioaouutQY4mPqh5GvvvasjIDELf7sA1XbyjMj
d1EgOS0IgBDoVboE7ZGWW8b/FNOfx6BpM2CIQTRvNZq+gm4OaWlTga5sSxZN
LuSl92P/6Qwu6GUbMK6uyS74gO9scqMZJ38EVt9Wz7H2w7LV9RiVi0M92FRb
rskSP3VXIxx6LoPBF1pZnz3XLMeoVAB3GLAvQPwtOytBsrUTlIvNpayOSqTV
/t51Bjjay+B6/mfEkkUZDRFS+FCQmn8ZayPGSxXusYod8T3MCVkuJaQFLc2D
FJWMECwa9/tT8LC2luacCJi135zW1s4jr71/9zo8lhinTFIzUO+6K8KGIpKr
dBo6ekZNgmfl58ibz/Jd4GuTF+MXtes4nFm+n/pSGe7zGG53HO3udkRG32q9
zoCcwihG2YR95T/woH02Z6EUzl/MYktsIM6O0Pn599bDRQe7QyyJ7Q0GyUAP
WtIN92qU7185R6nOMY+LJ5Df71j0jHg6bLHKdr16PMWZIUD7dPVXABiVRHAQ
5noKAYCUD9GvW+8liucgpxoNj+ozrLsz7JnZvTlbjBN9cpB8k+1dkVVMvk/5
WI8wGXww8tlZET6noQy6z6BLzAtglVLlAFCY9mxYN0lK2M0mcs9KvBTpDhSJ
jumsBKQ7fpP4imQDq9ctrdUilhAzFLpRYDR5zFj9nVLcJ/MpTI1BH5EAf/SH
rsWKoizuuyXucIaERF1lJi9l3sbxnU9MBIoCNWskEnJ7vpUtxWkCKigd40Do
73XzUFOi3gfV7383lK0G/08n+Gn5GlmuM6gmRpTbukstXUVoOCqrGUK1rTg5
NjeJojyqec7//pcrpigPv8GjVtsoa5rTMM0yz/2NczJexQFug8qu45pG8A1k
gtbrEMlQbF1clQCW6XpB6fmMren0WCs2QLPMEmmAyMycnFCMLCriCKSQ+3kR
D5TkeZkdAtorRU6jScimoOwH5blhN8H1fG2+CqpiYdDrmG89HGKwF+TpYyN4
VCgCgKQw0BukDx/DngK6q/gK7InKWH3iBsyes/0hKgPKpIegyQg7ZYHxDz9x
/l6wFt+Og9A6vvslHM5d0OmOUwbcYDpYtoAhY0pY3Xw/PmtuMriyF9KUSNgR
alxbaHueWYHpwNWgRFIPFhZlAjcVfTdbh+vJRmcneSZn+Wl5tvWSyYWSjxTc
DNK5t8RkqGTBGNLzOd9EqXRTScGFRnOxtDBxBMxh7x2OVHgzHTg9bgYdipyf
livzkE/+H8av+3uOLsQBMSkxYwF2bACQeFgF+QUEgVSXgSBGpYIU8r0y+GLE
gO760wsbhR8p1se2jQuD+PAVyipKWJXfqnDPzYzptKTH5oUZ0+l1R1w1QYJz
TXlODx5ovHQZ85dZYas8fxqSZqJ1T48k1Mmt6kDLKSx7oFHdQDHbwVGmd0iA
iojprXtqriMtlPqkYxqe40v10qT3zIMpgOA7NmI66W1trxrJ28ez3u5FmM67
knSRo8ZJoH/bDZgZrwigXVFVZuJ2Cw1teMcf7vmw8a9sZnoghPq+omgaFoIQ
d1KOTFnBCRvRXKOH1Lu6EDs4vHKBWlvYMZkWV1hwlVr4RwnDz4DxQq6HdOIX
MEPBIZ37ANBNtWjEZ5hThhTf+EFWtSPbja84bT2Z4maqv7wRH8VsLpp7DNHV
XGlvOS7ihlUvntzTKSfYeucnrGwRVVG91evVYXANtAbprpv9drtvBdvTPLLy
hOhB/+hg30KCA81+Rmar6G0kV4/WPU0AvquU5je/aASgX3ZZhOeDHaRcumVP
lZsK+ftjH38Dt1A2x9betHklppeGS2LGxggEtfFx0V63YVEs8BWYAbbvuG/J
9ft2C7KhGqrBMFcsZIeGpghUJYd+e5aQA7R9GwgN5C6g+j6gTCkBxLAbRXAj
R7CDqcLOjavSfKcxYg7yCopS2OpS487fK+aXUOmHNt0uoAZK0+rnfJ7iFu7a
A92Ng306/i5bThXWQS9vE/VeO4IIKMOTmNTQFN28P8NfpXEaztjH7PfXugwy
DbWrUwM3on+eaIqJXRpluLjUTSkjx8nugReSrSeWVdGlJdm/hcRWvU7BNN6N
AcJshppVCwNd+GyqPaQdyPaxZGotSMgek0lrBClYC04Bd5PiLWcd6ef4yGhV
eX5kuNE+zJIBR1sMgc6/PBmrkldtGKGIEklLLqcykkcnF+hywryVPIuqEoBo
wPaEyAH/KEX5WkgkOP0jLd/U2WJEki5uoFskfJ6RbzQadRjcIhA8Plkn+Flf
V6X3wZyMDlZJVbjxFIwuGRrmSOmEfjR0zuR/ziOIVq5BxcXF4sY+GqsF+5KE
boY/aEslfZnKpc/8oMsSvCva9nYQejECAIlDRA4s5boJWEo+bBihXB0fuzBa
irBT8tEgrUMs+0/vGhCj4cHd/FAKMAd6ZzSnE0E44fRCOzcTeu2vlNWX0GPh
ktmqfDWzmZcvFEYjdGoj4Fofcaiy9/pELt97kFiiFSxZCb2GFyeVYr5X356y
R3hGhMLfYAgVHk7pC2RkbTfRUCJoaEY0FoWn1FQZBJwsKQNOS6NK4PXUQXEa
PPzqKJIGpgTMRR4a+Uj/JuMl7gwhdQ92FogPcvbN/cf6taWmjL15srsyCwQO
3n5SgKlggdN6w/Fqwfb6UcbbcAcwKb0iBc7vNLrqPUBfkbBqhLgn4KElTBl2
Nvyo1Oktygd5UMrzlSr+xtWHoWzv79/lXnhln2lFXNKjbtTqAP0fJuf/Ltwp
8chns8yGSQ2xbm3qC6+RiLFxvlSIolwz85kNF/XBX7a/OgG+9ljz1QA1aB2R
yO477PUnrwt8QSEe8ai7NIa1BPiIVU9/RG8BeM2D/fJ1jOQRkpF4Dq/6yaIN
c9GH9+pbKz68s7exB9mIihL4+lduXPp/5N3K4ftBmx9uckY9egvn3mts9NCl
xzHWb9qoorKo4TAVQ2ux9HBbwk7r9TTmsd8x9zmscxkeZGy4t2pHovPhCSkn
vIBZnnsRJCAOlwKUWBeT2JySRRtE0fdHaxyPteuU4joxeZM6xZPzVX0XzIaN
ibLyhAKE5GwhHy8HHbxma4vTqSIqs1fBFqug3zNY8qfhYA3fu06uspxAuXET
HKeQjEM167LlK1f6IYThaUyinQuRaU8SwrdZDL0vR01GbBSWhRJkWSFhJTyL
wpCFiVlu4uzn+pP54gGSDroiqyCa+sR5glTLU5NJAHc8PtauKWaqyBjlR3aC
wk5TCPrLOw0GWl+oWmSVz3zXLdTU25eBeXIo/iGKIiBkIMhUeE+Nnx8N01Qd
cmzxoNkKDyo9BB2ImYfG4kFXC2fyMAYpJPkUs0Y5G7wffnvhCJG/EMbGi6p8
gHBATLv2WFoguuDV/g4p7yDAd73BgC1KfBhrxoEb3x64z8L3yPoFnomHkvj9
DCc5+KsMgYy1IB3M2exnKFlrbP//z4qWGjGu4r+1UQRP9kJX3rqQwaLLaDQB
NsCSxUv37E2KtWNOmfH9sjF671++wI2RcE44265Y96er/XJCm60BLjt7Hgqn
+tLC/nWOazVTxCHtIvtYUQKJ+shtwcwGU4pkgGcuwPPxcfvl+IaWbso9FQol
u9YBnTKiY7PdVl45B9bcfIVuwPEbIZvxInkckaTkY5XZk3Op/ijRe4xRLk8m
ZvM/TVzEkBAQAJ5gnTQZKU/hVrReswnl136DgSWsjP1wa7pXTnCLLJBNe9WP
j0jDotQ7p2bT4WJIU7GUfGNq3c2GtW5C7zaHsjSkY2K/tj9GoLegCoV+DpCz
IAVcZli93NJZ8nc83+PVZj5LLL7ofulIMPzV8vgN250c4eY9R+cLv/1S6Qz2
dg4qIoBX9AdxoQ1CbTjYwhEYvSTV8itlErz4LPdmWXmHZ8QRVzTRIuzuYYU1
PwcAkt5Q49ojlzgGFlZSNu18sCVnJiGC1TyF7lF4VyMr7bXbR6kb3VGiZLT4
/WhadwWlzvQhPp+JrvE9KYB9nC7HrRH0FYQrV/lIBacrCL4niNR5hgEisSbk
5TTQZLqdHoTAiBfzoIy1ImAklh8ABMDRfa1fUk1lQ3f/wJHEaL8yznO/Q1Ph
iDLyRgGtSkaA1fyiWprWnC5u10tkhOnqjBfR5z+v57Uwf9Q8SevaGB2dE1+A
elx0ZgEF+kfKA5Y5afRd77LZU+mSoHF8+cEe3AL/+xeKzGVmf+qa0KVAdQAC
774aPutLgZAIOz0m5Q+FlepYbtgS/JWYicI8fb8ruYRrT7hvczjYKnrrCWBT
3ogDeKyPYV7H8aiu/+16V5/XOL9/uLt9mGl+zxWQrSt2BpZrlS/Bd4++WXhW
aeBmy5pPEr6Ivymrng2hxcx0cqMpiLUOIi2dHO9YiM/1ZcLhhY5a1o/LiFLm
qetrZOWthfqiYAOKt3rCM5G1MEd0tKbeUgd3pnRM8LUSuZ8cprWatD9PP1F6
oRAzHBwZdwaFTP/fUGNEnniDNmgxlLpNdY1L6X6aPnyVOTagWNNgo6FBkGpM
kRp7GZKuLEYL5wMX7lWf5AdVmJiTSFvusGYR7Cd6ib4DSNloFYYwoBrsjGFD
tNaItZJBWBJQ03cQMF99D0A3au44DkvDMmqa6UUoo51FZZ+Zu6/lW4hIdMFK
bmiYQMREhgQ8dLm/2oIDqNiLr87PFfThgOdmHiK8n8TQFrAuIJB+LFbC57Qk
My17jNXzFJIvw5wnXqZLD/cNw/tCeVn3Sit2kxvJiMhqOuBUYFm4k4DukYQ/
x3QYCYW23DA7FAe2cNTf+2Pr15/S27Z5pqMDhtPWFfokKAWaIVQYLH85JdKZ
CJZ4+gc/pTTQvOPWA2ZDB8KNcaPq3kKA6lpjTpZ+lr8mWYY07G0w+A+h5nyi
at6LAFWoFaiN+txMKyRbsn4iWJn3I4BI8NufBF0zYWTyVpaLDJB4I4j3URbo
vPZa+as747zVghBX6Z0+TSS4iibKviayDHdwAq0MIqLK6bLuhLHosuHM7JB7
1PQmjH4bJ0Ypn50rYpYwAeTdqiOyVls/H2r0pyFB3ExvvyG+bNjNUjEV742c
HvXCUX4a+wcLXFp442DuuhY0vBliQlH5M+Ht+dtUcMxLesV6wNc6q+lEnXLi
i0ouWUzLNO9zBLLmMmRJPBd0/8ULsAg738wr7QVWhk48cbDHauSCMSmNleN0
I7oa1oR0U4D47OUxTs2JR6I/Jy515Rovc1HbkWbkIQ/eDFMeHfRobjqcpb9a
tyI7XL7cw0aUhOGSRDwp/5TecQmI3wh3qf7ucT+Mpc7QmtFj2RnsPh4YVSeD
T/BleEPsUDoSbAIHlEHLV0MG+VpFjZH7Z0fiTsYyqkuduqAW1YGXu/fJpjN+
wXME2RZqVXQ+RUECrNULmGKc8ba5vajQ2NOD3vX4VzJhMaf+pd35Pfl6L/Bo
VPo8UbTkL0eFC2TpjaIfsu7VEri23gYh/7gDNQlbe394r9qDY5q/q3siE7zo
mTm5zX4b4n5ATXGIxYsocdpXoocFLXbFZrsW3cbuskn4apWi9UUGbXORZuQl
g75+zTh43xFq1wx8SFjNHrfgWeiyVxGON5m1d1/f+9LfvnPQ+RHchBJgx6s8
S6TgNGvN4j7/pmvOpMbGvGR5FQnFv7ojuDUw8xSr6F+oL0Z5RRahKSNEZeIN
BFmY7YBljavXI7MGkJ1KF6/WtAyz85uhnDCWwdX5Z8lWGW93ODNc4cW9kb3A
MCVyy61Jg/kHJtIGDv7CJiYjOWAt9ipHfwmrHlt+JrSrfUDoiIax6+MMpigo
qkduQfgpTSdkKWpfvIRgBBvL3kUAA29U8w7et7bg/rGff5O8OQBOqP1aPonY
1ONWxUrhJMIDJohLImurVKyUU8xTRI9+dkaYsOAe4aqYdj1Kt3Tcf7PX+kR7
CuEccTwH44H81DvCWE1jb8I1svdOFJvJi16kflzCaSN9bEud5F5mNrPbH1uN
ExhBMy0RpI8Q63hX9sDX+y7ZsObGfi8N2JvL6zMk8LDt8d/YhsQvwQEDLDxu
uWBknppz3gGg/WS8rQy/6wlSfFsrD8Qqd4iNETpnv7pJHMoheUBtKws7wZyY
/w7QAvGHjTSf4lVFFjS/sf49dnRcRyXSQGSBH948e4Tgx62sDwhHwfYk5672
jW00kWer08tfK5jqRd/DCwjKBrxj2evEnepW4oWa9oshqOflXUmYgwiAQPld
A3m71xVhWsBJoMT1v4EH1vqzkMeG/pH3axcjLEkH4op7XAimVy+1mEM6JRqD
yXol9tMDqaK5eiOZjShOTwTSQdxdjtBlKdkOFWlzsEFYuIlFzTh2gSafa3gy
tFTKLmsqgZErPcFbWwOcN9PenUgHw+oFLQAQny9dYnp+E6uH8bvxvpUjk02A
SDuIW1J6mzi+9fBdDIhm5SX9+Igdk9cxSwNXUOV9G+R8kSlC2KukodZBvNI/
BrirOU7wgoO762h8nM0BBt+vTvSq/4W21KhG3gP7uivOPCHGNbpxWKZv7X1k
J8dY0zJtzdhtIy9JBYR4zF5CPhv1KP8BYuss4MRS6IGxJ6qPbiiWCduXUHYc
gnuNB92nKsvRZ1wffPt/vlAz57Al3pnCUu2+PTrMr378mSvY/3VMtww0/vKX
hrc48Yg55io+sQ15yJscHX3NtBCYa8A/6YgxYPyY9IiQcb7sVchS+YMK6bxK
tfhjV79xmZIpuAKhPZHclQqMCR7J6L1aYvowwXBjVKRO9VIHhhPqvflooMpM
BcxJ7WqX/yhylMnXSKhCCxHsHL7oV6GQEhqoBL5oMlgX976Or8alTdiSl+M8
3THnjvDksR7AUdJxLYaRNj4dCJhG5JLIwO1BPYSEizPWMAbhKnne/SZSaus+
DWBfG/26mMqcOUoQ3d9yatKql3Rn+BxA/SAiyUVASaWHcARXwXDZzDqFM0nq
4/TfOGbTQkAd6qB1HfYvsUKqJh/Xb2/nNB1ij7Jlqje6uXx7q9tfW7gyY456
MJh9L2Ka5FESzGGd0y8X91OC8CSeICdXz0KA8/EP0Y1DMcL3ez9PQoly33vQ
HO554f8JbyhnQ1bGbUvpf1qFMNgW2O65rZLFfPD3uVkhZkVHWTxSyRpzPFNU
jmiaqON4YuBxqwWBdFXm90qmetB/HBJj2hmG9ohkbQDbvFvjrZ0kydARDgft
KFpuFg5cUA0K3tmze9rKsDc6dNdQXie1suT8RvAMqjIiq0ZiND+jyJ7rqZt7
pTAuJKk0Th0dDT3NlnM1sd9haYCS/mxJCuJtdvnVVqnX/uZjbpWGedUiDG2x
s1rYBbS6ZnB/81c4NznRUBAgJdJ5fOSYev5cIjWcBHiQDqBCu4sC3C98Gxax
OFcqqBF7dH9/NJ+uUiwDouv7yjs1bu/ZqOuHjVkQB4FPEr+LiJ9pByVGUAgF
ox23j9gaoJZtoNM0ZWkVdkTYoL4FvRGJ2x2TOS+bYbJ6MVbVN8jLP7yukouv
cj89HvFDY7wdyYREchxQ1PsB15t+qpSwAR5XNhAqi0ghYW52CG4iB9vrzmFw
m+Dn9rTOEVbl9d5C/MBrw5ClTo3x6G6/yEFjlwQ9AyBgsQuo9cIhRCcrkjkJ
A3nKrzc7EIQ9xIBKW9J6u119Oi+Ya5yUWiGi4XVoCZOu2R0IAFbh/eEh910L
GLqKqgrCHo2DRtjj7Z7a/DVT1tZhYJjsnb60rzH5bgPDFKnJxN4VEhklOH+I
QG6aoZoXh+sb9cvAVGFdGL+mkYEr5TTvg6s8kdQrLGcVfQxg7SYac1AuwkJn
nwrIktgycfhbjYUWJ/poXTp8OsHy8YbxUuii/wvalwboik/p64W4Oq8V7QBL
4r3ikXLlhbqedE09uVHtbcJxSLmiRsA1nWDDrDgZxsuV9AlOeeedf7nYYI0U
ZfTdjISVN4Vu4r1oz7SwOwj9eMTV4ZGtARTN5eonfcXwHvUVyee7Vf1avSf5
eUPpSpoMkt+TMCGEWdSTltY8WTCkv76vYlstH33eT8jQ2ulEpwJT9H3fj9ev
AWMTfk3U637npkJ0KL/Bmiv7dd6+ZNIcVDCsDctNrFovGBLnjv1g1rydZ+9p
qPRHk2JJ2swH2Nwsad4MS0X+lJ0ZwouNFwriFR3yKPr4J2j31iky9Y8HzqiQ
TLVJiRaxce5MCWSfgWkP2Y51/6j7oW82Qgys4gv4GiEpqgKyNmcB5qONACjh
YHRGN6VtobDjPvky4fQv6kC4nXdAcIjlA2WOf3EkE0l81r1NqZW3Bml5A4DA
rVI3mE0syGn9bKxGKRk68//8Y6IIpc3NCCc3am+j/DfHcbkAIebU5XYc7pnj
YRu9j5N0bAos4HQwakA4FtJz2y11GRWALpVU1TBFDga9wSrku7NhFgq4U6xG
zT72Zmkuh9mA71yL0PHlIQt3Y8uSL16nakzZjO7uT0MC32wa2TWf0b5rcA+f
75ZpjTFxO/E4yPCfw2MiK1W2pecZIz3ZbjSfvRaxhGzsr19WujojFHVa59D+
+a5EXGLadBtgAAWODp6pgv8tHpIbkOPgCru5Q+uj1aFnT57VAQD5pV89RLcp
EJyAKIiO+X/2mWCwql0UPZhacZWJMxD6xlj2KaT16YdlKRboAbrWIDhaq1cT
KQVOUN9VurSGqL6HpReYKRwsP33RUFNIadw13F9tmneGr/maY8gcfI8mipyx
j9kttzMKmzK+ZOg8fmibGYgvtPE6iaGP6fzNrZmx06UtGLoHqVcDsd2GmFB0
aUqSs93i0JZnKF7msLDndDXRWwoufFpUgFrY1uB+EMGBv6q5bQQpknOEgk+o
chieRXJN9NZRpVFPbuP0c4wiiNx5G4NpN2WLmN0gRpSDddt8ZcGa9/rljQYf
aDqsymz5ywuDscXqSb23DQonfJRoKPMkxZpGFBABfRavQOGhatO4vsQPEkqJ
nYgqk1C2CCkqyYsHB3qSy3NAcByM80G3CGn4ZIIdAIKWEAWuSwFOR7HD6lV9
tKwbQi5bXdlMUaDigVcmyu0nF1xSuAOqzUJeIrYJzfYRBmV+/yBPtMC9hvW8
/mzhN2zWpr1pHCCQMEVG706qpOEEPudhOycHGCsq4MKrJHxv06UlSYYg1zDc
CK/inu+4j1QhEhzW6s92d9hYV/1/egMsNcXPEAkWK0j06a7rSyXg82MYtkKP
IcKKL0Yw8Ma1aCK3YmMRce3pl/oQuZaYSqMYSagMQzoIY7iJQUyNqscdsYdN
mNQVBhVAgzHao9y7RqiIH7L97B81S8ns982T/Eq1Y7At36nEUd6yMa1BvIR6
NYar/8KKGwppJowWx35tNvZh6P89f90WWeV89UuofszNZ8khhbdeb0VTfJ3U
lcvZtgSS/4hhWiap/+JxQuSQT3jz0MaKKzacTpG5x2KUN+76ylBHSiZWzfok
lQhK7v8t4orr1WANHbA1jhw24fBSfgTBc/5Mch83r6DqJ0z+/h8qK3Xp3l7C
EQTSXBQ3uiM4MOUYMa98Pv/+7PkRrq1i1BFQ+02MRk0ablma5fypBxjPwU52
+UDNB/fGLAc47yGM+k0YmM3SMGvFxUUmS5d99AthzWplB4IJffmqUiAGvCL2
Mzz5khsqlbCpD+l4Ox2O8Ip9P5qUFvoUDBSGHi110UOOB/nXsosd431SckEV
5hBklaRGW+5LXIlwEL64QBZyVvTOqwW7TQfT5hkqM1v3n958YlQ/9n7ceuQB
/aiBdTq+RVr5NxpWHyzdb7ymwhPfDo5McpNvHsBOqgNqofBdM2WzEi2X0Qp9
PE2EkTAg6Wf9w8wU8LWj16MS+Wgs6HT/KeZKp0O+XbL2Fal++bxWTbv5DWFz
IfOiHey4QXPN9XH6PfpDTH7ziqddvJwx/o99qDEJ7NkJwCEWpvQGVRd8cnP8
fyY7YTh11fA2vYyQU5GUh0EYlQyiql8jCOnxmOuNdONNzTQ8xzE2d1cR72Q1
YDjteeRtNB77D2rsyETMkjdqoHRws/cNCmVNAnx5uszuBbcGtTgavJ0KDVgo
0iTUFn6Tnc74E1T2y43n0mKKYfNwHaidHVUhkeTNy2m4QBya+FXoucmpNHz9
x3Hl6uUiYaE3GaKUuDaHCHsrXLEKpaQskF461gWo77DC6vcJDg0zJZi1WthK
UIpfNr/rA4w59F7BH0TWcrjUYeT1/D2h7+DeDHY+0B5FdNM08/AUU9tYaDtn
8aohLU9mgivOwa+76H8xFlJAUBEuqb+12s1BtnhcBL3CxGPeKv07VKAZsaFl
6cXN0enp53Bb4vHHj3x5BL2Kd02Ey9AhYJmGgQUGHuPvUPYAbkTWXONLKrWW
tookwmichs4IAQUm8c5Q6407sSmGCS7wmL2wX5TB1fmNXAM/muBGXfgCbmQW
4Zs+yaPqTAcJfOy+Gmy0WBRscA/h0hqCKxo1c1xxKAmBvwPPy4usnlYXWUyI
huIOELiUS8wuaQnDLZ6tYy5unOc48rdmS2E0ZUeJO2sOWtdmqzXT42eX+A26
LPrNm44xbmdH3BMIkHeiTi0aHHQT+mPqdT2qX71jNnTFOGPgtL/WKB3LeX1O
i4lDCeC7lNmp1N3lr0t7I18RH5CG0JvohN/PDMyr4I4L8Hf8c2/cfy0GmjKy
0QEoeyrMSlkOoNvTvhij4zqr0WEfB7E3ZgltZwauBTDWkrAiO7Wl0T6FNKKF
TX2yufl0FbBLN8uu548q0+IHXklQzjBIqPMV9nZsyj9KmDlrQCko/RJC8bDV
Y5CRVpsB8asruDMytI/4+iYRiHbsKMKpxE7NNJgf/NL9av+XBejNkEhdvnGc
OuVQgzzLQk9PWgczouP7NvGxYi0XNG8oKTHeoQYXHDxj40E+1wWN7Qq5gXgD
JdAgtGekbQwYwa5pVS8CcmYX4ZsllrKr9hyT2wtd5O+sjmcoiVAq3YOHcO6j
hn53h+WWoZ5beW6UaNhIyDg59tJHwFl9BfZfsLxgVahxPaMuq8EKBiZYfe00
7AGzEvKjoMdwka8Fa4fUDATrkLU6GiD1Q7awkiN7B85fhF/ZhlYNZkFC6KEC
CXJzyaRXF2jmdKXn97RIYOT6znM4x3+ymReqSHsKHhI/bcjiXH48zFd5JH5x
17sxhg2R5puXeqO3mzUk8gd6xFuPh2PB/NEhhoLGwdY5izwPCrbeIbxVD8C8
boo2qN7K27BJVg6UBDdoJ5x/Qb5LpdNseUWTHejsZJF1WDJWTaDMMiso2m1e
s4AWVY+ktqtUPSr6ofTkvyX1iFORlCqK1vx7Gs3oMPEIutH4rM1u0vaNrdyx
A7V997E4E8gz/3jTBi3TcurVRcaJpIYGHBdks+u4vjodL4tSur9zY2BRFRr9
Jt5489XzNzHzurRK0W49zHSH7Ud6wHLmpBIJ/CnrXs2JSocjdxYYpItuntBE
QGtkqWiqopYR9by3Wbokkp5dbeB8SBcF5kEoOJg8iJwxedPxEfFuYX3qyI+t
OxaI5dNV0AT0MyGjJ+4KdP8v+o5JyZ36x5vgmDbsl0H5pGIICOLTauYOU+rZ
mLDsQ7GDwyupfXzV1L2rLA3zZztK7DE5zY6bZydezJf/i8HlvFHujob6BWaX
y8pYDrE1E23IGwecBa9rQLmpE0pzU/nTiFEAdXwLNelKR6W9Mpzfseq0VcMS
gWw6h+iYh9nDL1mK23jYFVS93DzCW2POc94UfBEMR6xY9uIaiTqWhmHBZ8xr
nNkND036Yld0fsVW7IKRAHDKayW/di7vpWiyJjM16y9+pN8omqIcReudp69o
OzkoA9//ty5P0f781zjEs1VkVM8Lkrz7vbtsIdwSlNNDiR4MCZHssQfaqd9C
cEAT4Dey29DRRK+mqWm8aLkg1D/7R4QYkzclVC4ryxmPAXXuu37A36750XNC
XIUWHo1e82ADBgIZOXKn7JhxkEcjlDmCUs0a0V2vtNxFYVXmsNjN5HKdMybs
e1rbxmQzhU3flGm77+FsnIFFFFG4l4I1x+Xh2kJwc0FO/JMFm3PHBK1nRuff
ii6C2IuMnM9lIrlSxLAP/46xZ//EqPrWl02G3NwiEKqPuu/C3XspadUtZmcv
zf92+PHM5t5u/8pX4C1xaIQBQ76uGKa/RygMbVhRlASKBy4w4NwDhsghJ5IE
fBTC/Z8TU7tz6hNq0EzvccZxDMZtcpbCGmM+AdtTo6LJmqSqEjuVxBS0PQQU
562yQf4zbfA78AZOHnGMZ0h7SpVH35/RffHUOWms33svz9DJnSTyc1+QoZ6i
Tmqy2ddBhRjG/QgtSxQsxlkUkQy439GW+QCGY4itJ73XQntlGr10Cm7MdR8N
HzeeaviTHzakVapw0IlMKgTORFMoVAVIkS4a7CjgQODb7L3FlAsALp0BkPoj
eXWd8DPvKVc8a7nEMUV+P7ZtPTMkkdYxodjBk5iDA6bfxex/RCV/XlWiZFDg
xOoYYtKntHaEmX3VJpX/DTmIwXD3V0xEWw9jQxduY5jgc7eR9HUG2DHbLVm8
zsj9f46XRLhTg18YwSw2mj78++yYk0IKq8moYcFZodOSGMn4cK/PPP0Tni78
hsWTZXm2kPLv4VhL/TL3o7tJBhYHymE83rVFIdoJEdbm+GxSIMiFu5QjHRYw
CmXU6q1UA+FvZF6V80203sZMKBNz3oUlE+OdQVYW2OOnlAPSOvpGML0ov5lb
jbpkDTosK6mID5G528Zon2qS1M9ABQYa7mCRp0Jy/pB2pU6zdyBruN/6NatT
F2IhBwgsffR79d8fuyY0NtadqRRl9lclhKQ2IbMAzokCVuEbjCmhgqpAmhMN
b9nLcqVVvZYGVcF9tq5O4vDGAT4zP19wCPOhcCixS3m2JTn2XuJlXrg7r/wW
v2ncKLWUCnXK5kNC4JoPhV+XwXF3WcnrN93rQeTNuviRTBUbtLNONHwf2BMO
geDen7a1iX/a6Rp31XOo8NG7zDrAJdkFbO8vM1r0rfT0xdEzWYFSDTZy5JIM
VvJf0JZEjc43G1372lGCwFrQrYJfQG2kKTxQ4vmtwsDBEqmHnEKriG/tyBgN
/Et/9T+8mK6sjmtLOm1AN97o0x5lN0AWFTB1T5qu93WaIsr0YqtpGgUgARod
6MofboqepMrIySatncn7cnnJEVj7rWIBxYjaF4+V0guBnLwgRWRV8RwoNRDo
emUe/lPyFUP6ZNvkvFMGL8Jb93/kXj8avHforQkKEzecqD9vU+AfUM8wTlYh
tJMkg5HF34HA6Q3oF+HddQ+8jAbc8kFLA0FYiZOQ9YK6ShjWZZCUNhvJ4JQg
DI1krgtQbpebnhDbiyAIgYVqbu5Akj5tTORw4D7/ULc9Kp5jZ9DFlnlZb45Y
MIbiEbM4wKfXlgtGOZ2tjL8mPJJrKozPNiDTedWoYDhX7p7V2VolYSh1Vgzy
I1Pni0JHvq6QzSTp6GBME04IUosrJ7sP+YEgmiXrcwkLCxUNd8AxQfWO9z9h
15HsZxNM7lH3rv1X+OLWp4GdoaqqVRyNADEsdC3zvECh0yb55agxolpEveXV
NNFQGYWRzZdynIz9MIBJAQ9MMg50nwJ/IkzEKkfKKE5M3bhwGPBzxIrPvQh+
UeUGUmxkc7hlSTINKgEvllNsbx3K7GtkqgqROux49XRKBY661pDihLMRb9Ix
tQgHRFoFpeJtJ73h/k0wK0sBQ6bXHVlC2jTin8e6casVFJzjhQ0TklbluBEX
7He5upNGKBRrPQ8ShtDKkWIAIe8hf2MNrygA9SxeBsPPkYJnfwMIPLqlKAzy
P1vT8XouxvJkOy5Gg5UFZFjrBLmK6rq89W73xeTFH4iGGsKi/L0wZGzYbQRP
PbiVAbDviF8Y732nZJoyoBT8Zl7Pmabhu3UB49/RV/wROa7ZYIP0qfx/nHei
i9icENHMT1KQN67owVzSVdAHvsRFHNV81t5G5nYEJF0OUBctHZRmmmTbs4tE
geSY22YzugYAi1kvjyjet6LX+AH9BODYO4FnQDaFDWVuThFKrkbG9Q7nQFjE
cgN5yLSZYZ5EJf6r9qODmysqT7Ft6cqwotoxuUzEE7jDxrO0qbqU/le6BTpG
JoNV/BGnuSwJHXAtttbCT4ssGscIEaKbLVpkaFRpXNZhGNR7WtUT3lZU9B3Q
rVG7fF0Ls1FqeD4b9C4KYWQyDxDntcJB4YrLTbFdQ8AFJ47p7EnlclHTfh02
0RENfUaqA+hyobx/qhbdeqwYjLElscnUeBJZjbibcnfd5KTf/1p0lPKSW3GT
I3OODhDKyTj589HVfbZ/w7RImpw8PgHxScdFbGfXR9b+6vd/yAluixWgIIG2
Tq0VF+agq5Y9w97yiXlJOnAzX9YT0r1iLSFEnApt3wvtgDK6pzL90lkxNKI7
yt3mzbWNWKMIi0OYsMfr9oiXl0Ss+ca3itQbHX0IFtCXLtOiMHG6TobhN0F3
SBDxI6LE0XpMXLJ2PYeXLVzwnR4wx9HAUwkRltLpw3iRceTF5+pnPgE2ogA1
cTgM+fGi/QmA33zj9ZlgkExvjUIG8e+Nm3HI0M0vZqG+glzESUYBM92RAB/m
AaI9PKbMpyw1KwdpoYZjiB5nHU5wJEUVv1MEgI0FTN/sYmVd6X5KWSGvfCCN
RjgBd0L9TiPdZsNXAR8LpY2zwpGawofMWrYFV+cYeJx6C4ClABUP0+OEUBWC
ypI3NZiM4YplvGHSLxn/62/4ScgEMUDDcsNWHYJSiLCGVIdzTEnwMCD5njb+
OoDhj868QykiiSUxqmlv6bM6zrWFLgORff8VeAwstBP+5LYdGeYB68wopk5R
LwJbnZ6dV6LlSYjFaAuyXMZcXhmMB4aDVXbW/akJw2GrUsAiK6X3GmhtEBA6
Ueeap9yzwnazm5sf1KcBdRXbb4pNAnClRr1KJwnu76jbt83Po8fj+YY40yB+
25D0q1k7byc7Du/j+DAowoDicj1TpuSoHau38OyczndVf+mscMNypVidOKmB
kSFL/0IDNrGbdaJBBc5+u6iqSDY6kfKsU5vzf0A+GCAgIaJrFtBoqzdqvajM
Yt1zi+DQmh0IFNiG4E/+Cx899dEMERE6wTwzZDggY3oi+cum39CqDQruQGzw
VNidgciz334oJS2VPlSkRKyrGLtf/4uaFRIRyeSvBtA/ugDQk0mD0RTSU3My
fGXE3xzBVjk//5dfRk49eT+0lZl/Ea8IwuHwhUUC4CDDWpOheDNqwJ+Kmh0C
cTdJRGZbTsLZVWJ3xHzKyjXiXgWxxoxM07+SaLBl4ZJ79a/zPPuaQc76f4KU
21LJqD1tyarzS+VjOHs8KYACsYCh0qymgAAlqg97vbMjCNJygUAtQhtfbfCN
rqy/nYJR5S6LvjyKIuxKl8ytJL7QVbOa2KYjQb2fnmwyo1dgEBRhRfC17gUI
+aXFA6yMZMwckc10hQ+jnUX2x3c/iUgX8zDuUQ07EFYx1DSmnijay2uUzneY
+mjEzGVdvV0RCnAuF3MQfUZ3AbdcQcCnSuwJdAyHr5H3VNqOAtnGZVuwEbWP
AyrIWgYju3DrRWl43cjo/aNGbYDdRBnBEv1/6OvEcF234qYfpZ+YGNW13/Wg
MqEO7UFPT0Ss9LjW07PDXC/ZP9Yh7rkPrZDEbU6/fcLZOU1C5nPdJ6V1KJ28
qPkKJ1Dv1AxV+18hcrh+dRq5fSEvDqxkES9kd4ppMWj6e8L3zpYRbaydEQJh
/VwOeFsq+UO4WvSdXJ39cWcSelGcLFER+/5CzUeP+p7Ie1myIDIXoZFyNJoR
bH0BrUHXLs6stOVxIMTKZU9QcGBMagT0GY42PxE1ORg+m0WkrLkoMdRUD9rh
ovxWTKMZlFbSvLtZWVeYBbl025ZjQUFk8FNkTpthzNsGMoTdC1TlMf2mZi4U
C3W9irWEzb+67ZcG8iU0HFbSJ/ONOat5hKVI/+ZVoSEp/cVj8hl1L79m/o1O
EH0tGbNdaQP/Xo+2vfrSdnMUFGRUMXaQ6kmg4wTk3dJLq2BOE8pmfJ7W0n/5
L4gDR3yv7n3uRuMqhazoTLe1ogwG71e6m6JyZ8ZBcDgKdC5xyTIX/MLlXpPv
lJMbFcigsH+oYUZ7pWBG5CZY8fPM7hyfoJ+gczUymVEaG+/EunxP2/j7/LMD
Sdc4lzaiFYz+0UiD0eWYrtXTJda5KPV3ne+I7sx4sICy83HE/0T6ScbRRzX4
WxXQBmtqr4vQABooaBMFmBx91xa3HBI2Lo2h/KEcnfyWvMxfom+YYdyCkbDE
938XYgSiKfVtUUKXgGa59+XSdUZd8expt5NvavAjr/VkoLwOc1QGkTR3KWVk
ocAwxb7Kqfmkmvz4S2YtPTfU3tM5K4jZe7iFQTm6K1B8erwH09O6/DIQRQXo
xFExsYKajZQJwxBO8pEo1u+iZcni9Sfkc1RcmihKXIyar587jm3iXBV7HZn9
enBwEfSs5Fpd9zssUqkL9YGe0xtvDgki191lDcx8pNAFE5m0Jf46AYgqZ6Dt
OqZQgO51Fts6ZpEx/DNklMk1L28qv++Nm9doPbIqDmdatitWsYCUTgQpAeSd
JPbe5IkDGHjVX4crqlVUI5s45OYhAO06arDbhTpUb5/ownHoQzViw2kAO3o6
5gnpbtP1YGIvXf1bG3luRxAhRrKUuwgD2Aq77omTaCxdzpRmaXOwx0o9uO+4
ZHzh5VoGfH/Ij4Z2rD9F+cAZsKaoAJ5jMKWd3WAYPkJR8na3H20fc7k6S4SE
F2RPteG1B1536TzMtcjMVgeTOZPKBP3NlOkCFjQoKIvYqSJAfJI47SIcHv+M
Nz2oVjSavcbUygmOiJdFpPBTFNj+D42MuQM8HHwpfJBbq1HfYF+kkjJo6rd7
jX/HvYOeaq1LqgqMFMDeXYo/3JiNvT8Ewfqe+VckVtGX8Im/OtXNh30vkmTP
G+oTXTS2GAF6DTNo2CyXBHNk8jh0ksth9CWlZftb7ebqBqsPoXdW8gibx2BD
V4Wl0BaG7gmc4zKQTLqBXz5SYbFpCIpliVZ3oiIK49hJqrJm+yc14PwZqOLg
YsJ689qbM+w2Ky0UcU/c83R+ha+a4LdrLYqlCsacKliZjQTTGkiZBaf+tMUN
gciChIk2YUJMay66aVB4hXu3mcn50BsXUEwZYD4vNPk4JQAdGwLJx8GPkFRB
cTx9mDbFnVlW5jm8xPQpypZjwpxR4MjGzh9ep7hLpKlVQ1f/9Mf/XD97I5rD
DCkanZokDOO69xyPcMKlEj9Dxok/IdfYi8tIEUSkRQvBZFFUvuvNv1V+MuYc
DShACrAztNslTT0hcnFWCUM435z3I8dz800sapsvucjEX1BGnFzZAwJErtx0
Ls8V9uNL5t6f7Uv631UPTVtEY6bt8f4O4cxIkfw8KquiSnZi/72UNDOA0ahs
5SL4fIbi1iTvXOQ6NwrxIOAj4c/j5um20bze8r9nDK6ctN4vH/M9a/7r5Unj
US7nN1HZpUosDxWnbLMF2DKVbY6c3U/8ZzCzyuOXOcQDzSdfUBoYmhmXaq3v
q1rMCL1PZWW/72eUVvBbunx4X/cgDl4S+hZvYEMoUgNr09Es9ri+v5EquDdF
EZd08gEbbbFkP+sJX8AaolnTxLMmkFFrcCmk/2aUEwg9gTtEeSaNd38Lcrye
4h3YKC0IJcv/TZzoxAJzNGFPEU2tOimrtJKEiWbYeimFt2hvN/vnMMUqKwNT
GwV3zkG/4LBxnBVtcxiCS9fF3pmjRLl6RvNyQsAAJpO8XKaZ7pBdEHQI+wtm
6GYp1LKhTdYGvzvSyJ2mEGPfg6EmsK3YSknpy/luWXXWRRw1p07U0mjBVs3n
LnF6VPJh3Ar2wLDdW86oiaL9OxscJduyyyQpFiUB/x7x36o6Of96rgJMmw0D
X2rbUvhKstEqlDnDzaJka2jdMgq3kd5lVCjlqEiaRfkWdRGov1lTcE2kYTYW
PEkNP2W+VXm8bwH4EiC9w3fM4Y9vqGQl6h+gLMjbWFMgyg5cl+iiWa4WsXfj
hFQKI13uW+oBBryXoaEVuPfbVHh4j63cVnAq0B9IwlD/2paodD/cXAW0JHNa
o/ogTnQ/nk/R3B51vfIAhGm+HARrhtVY3SgPwz2tlcdk9F5H9es+dIoU/yWO
AiZr2BTzWwzzLBLwpMXNH8cNsi9JiVDSEojwRxS2rGqViNx/hvsaLeCZnUzD
Kg4+1rB7b+vgZRs6CEC/O8m9fUu5+qwnySRqRuWgXHCfaYqLuoHkkRfUAJdF
W+c4baogMdPvdcTErmP/JN9rPu7kQ9ReHw8GWeSnOPnyh1ng7zXtyM2DRlnw
M3xychuED6ViZ73Zabg7HdH27wWKlRWaHwHRfb9n+SuGWtAkB1mx3ltem2o5
pDohzvTfOgptzSoW52NPQlrze3syHP05fg7KxYtIpEVN0eMtxXWQwk+rYT/T
t/iA49xAtFhJj5hEgh+14XEdensuiVEM661wTYa2L0rB1excPzPJBJFD1BQR
7ACpqSXTx0x6BnDRWVqogGo2rWN/780us4tioiy7zgs7YyWieZ+Pq5NNJCsu
INuNeZsLYkkQsm1c2QmyiG9M0hFJB+hHxETkjtCfOA3xBPKhpIWrD3v5TWvX
RMlAC8dkC+jAod4MDC3qYlYI17xIRQjRlFPJh6o3PDjVnO8iVwV6EVM47yqJ
It6446LvBysXNyPZJqvZB/pSWgQwEHJyKLKcdc9BqLHX63BQhYBMjSU2aP2z
bySNUMrmhXDZQIrrChKpkf6+rHt5Fc+n3D85Huiw7P07qi95KPdPZ5/gZ2no
qpL7H2o8NLkMuPNHGgIXsXD90Xgqz/ej53b5tV9Gk26RPt5f4VaauBggFtFX
5WFVNv2SWn6nWzMHNwZZVDJqNP603xPGQwEMI5BOZy8OaHcZpDnC7Xwqwiv2
X+M/TSMLn2+6LJsEsTfr/R2+aWrWAfKmJ39cL8Blg8GnW+oq+DQsF8ffUsRQ
ZJS37c8HJsq+9QLiB6JKh7d/Tci43ugPIFVQDjXUoeba4GzRjldssVHY9T6q
eJ7P0if9mIPTqJ14HlY3Ua3pnkTsB1ps/+kRBcnax3DkG98qunbbF0pDqTaM
EM7ryabriHCiydxOLaAfWFB/py/kyyvBTtoPGiFQlfJuD/ismjaKRT8WhLbW
7Ukj9v6QvmeHGGUoL+UHYlIiAS/JsOgKA1+LV7zG8UyInkfvyH1y84ED5wmK
DfNsSHZLa81eVnRC1zhdefCU478TABPgYO7HTSIOqtWzLczd1Sdwt7zxCtYZ
AqCzUiF6zyRgyDKAcMQ1I9iGctS4wa72DTSxNqbeDe0EoUj2VWCcITRlkS07
rIZrdbLkNK8E3qXbjIMLOgcQ1hUJDlgz6Ta2XubVXalG1M5OtKItFdCZu8Mi
j/Y2v2oG+hVw54MPc6rOD1F1rTnLRUIRNg0kFD4FW4NuaAwuoWZehOjCYiW9
ezBizd6yIF+XV7zoTmoD8VGiFpBVFanDWyY+oAVrlscoJLcIigGTTjesRTD4
xWvpGfXCexzDeJ+rtS3wckrH6YGr1HoHyvc3lSaZqnxAZBl1Tl+EL5wt32wO
wypsSwlTB1uO/URBCQF1WAeWTCoILMvmz6QizOcwKyC/Dx4+MegVCUAT7FCC
Y+n9J0EXoDxzMP/yTlavQ9JVDwHpKnHodUGEC5PCv+XMBghHikqjeNmkhHlq
fMaL4FC7swmjOZBsEXWeGMqckGCvBIGlrqHdn/2o0rS82CLUnzdMQiyMWKPC
TliMYHLWbbkiU+2wD4rMy8/PVSl9yaY9SW7Up4hrvpEscXHF8JSVd/miRND6
+wlgkCc/S24Rz0SQ/LsdOUDQJqjkptn6ZBKNOG+z2pNBprDsD0AUvLHZPOEY
f5+gTDa8L1DYwa811/41/d4mZ6Ikh4SkcLS+SoUTeTmq2IZlvGXOfpe2oUjI
7bXCWej5NkhxDG8Ur8b80kmQv5KWb2b9HXS3TASo8R4FxnqM8lGaR22kh0Fw
l2lyK+TSXttuNh5gFzzuBwIpBFPc0bRCOcn6Ooxa83wTsDiUJL9fMIhlk1WV
b51Xg+SGVsYDcGWBKVvgcuV6hEE0olg3CR7QRJaBIytZOGljAEECUC3CK2BF
R1IlB6RFCbeJRBtFVvRZeOY1r6hpITWta3WQekwl3qTj7XH/9oSyk+oSrJId
CzGvPyPJwZRuQf1kyb0X8M98CY8GypDnc6lmeb1ZyrO60Yie8tLZO9H30WZ8
6zszsJ/0QvNzW5WurQrNRsQF2wxvWC1yDO2lsgYIhSlegWHYI6VSKzfWrfdu
6rOdL4XW9BK0pvTlBWKvGVsZkXYkFYAlOCTp3F4CNb+WPS7R5/bHCj/AIVPt
E3rXajqL4JJMCLB9anwfKvT7pjXmg1gWPDKfn/ROrkGZz56sIoj5rRYFBgZf
xtMY/YfDgbUyVw3q7sJhFBY8Oud3LpZDfv7nU9HpwPB38tJd8WQ3Ei5MApgr
kwJUBTY6qx1pQfeayVZxyKoSnG9z13Dmogg9v2kODlDuJnj4bD5fYU8k1tV9
zu4F5fGpE/Ke5komTVJ6pXCqjA6oP6DTR/HdIVLC0Ub5dpVJZajsrCYSh5pZ
xxLVLJ08HJeTk+br5NVNTIFTMbjD8apF5BiCU4+Xqegctlqc/R8+UPqOQBlH
GwOd53HpeE/iF3UggLLwvryJgLcIdZVHQa580VswFpMXiCF6YNqQ7X789Fz2
O/Sy/oDp4Je48UUltS3UurYY7iKnKcAbhfjdW6Xr250gJNrmKCuFEUn5hCKI
GuNIxnaTC700CPsG8b1TKVhuCy+7gVKjg/+Jjr17JP0Rc1uRIyRg5BqlFgJI
nZK8rkAKhNI/dcaqe/4MEoKsYIDM/iGp8hhU0YvnHv5FcO4h3nTW+VCXJKUZ
ZForFlj5t9G29FlwcTFEpKChMjxlMpZGzTh5hboK7efgAd7+Olp7vq0eAssR
FhmJFMSpIXXCycmVczZLwTzpwxhPMJ+lFBiQXwkMt9ZcwoqQKFgbYnlV/s8o
1PkHhW83obIOH/7QsSbhOsv09zJ8mO3htesNU8ASz6EbPbzbIggXHv/JCTIB
ycWPeJmgaVcZ1UHFG35ymH2XEYwFushUjf8/+7QrNe5FvBwwHmQYcLvrmwr8
UwN758q2/uNuThC3IBX1QjRJGjssfmzeRAX7SHgaxGaieQQlph8Z8fV6trdf
vfXQbHaltBR+EXw7L6bspa2zzwxGgHu6pf6bT4cTcZipoC4G0zx2y9bT4NVJ
Vvnrz7lHY/zpjNUCebsw3PeRS9i2CnG/GGXZ7Rm5kfWYLV4DKrDSh4SPOcHg
kOfyMQ/G9baNQjERLRyajU3CShlYW6PwkNAS4MudzP3EAT7PUCNGwhpW2ehb
gHIzKSWGriler3FFVPsfdw2nKlbxgAubkGrvc51K09qhHIca7TSJI6h0NtGb
kmjXiBzd52blcxrbStjkAY5hWu1OxzfYNvS5E7xNR7RQAUh0NawiqEXHvEUl
GGuMFJNmOWT1G7nrpoACD9xVYCVdq0ypCR0o6jdlLNO1JcENKWADL3bM4rsJ
EbPBlaaK+3f/lv4oJ/Pav6sGVmFInLfr0HaejFsifQStcfJ1h53wofGm6QXg
33YgTLnwXuQNa1/b65W1fN4Sy9aeFHDd7MDDTHh+MVPTmYhaNGwFuYZDXd8A
41sL8bCdwYE2BzkgwCbIDkbH4c+/nJ9trXBCrOnJg0M5GxCpECm21gpFJ9Ez
qcAtekpRcUfgYcEYQba+9+bHwcdsD/kiSHcVClhkIIe+aM0SCXxzBwaZTHoH
y1GxG69V0KaF00+rRJvVdeVUwMfRnQZGgw0LMofHO07sHiv0NXvE0aNrMqXh
wKDYDTSEPoXmuUMzrljjSjkgFlF97e0SVMAWTMILvMe29BmHyaZMHlnbguRr
ibO+tRsqe0dIdfdrT2MwvpAOAFM2xJTJix0A/s/3IOW7A7zRAU3tJR4q4eu7
/ZPzJaYPzKP1G5xCMd11Cm5VQw9NSr7arlrD0doIhgl43NuimrjScBG5JQMj
wg0542AgFRfDobWFRC/GqSaa2QKzGCE0yHdXNpkA/HRXgLtyg1sE8cEZnH4Y
1DbbKslkXx9cTdgqW5deduv4W2hl5Kb37HgB2VtY66ecFivVAtxRiixMSLym
ZvYJDKc22RGvL5cHKlyYi8pJO7dhuXk3k18U2Xl26//8FmA/6trCByy7lJsm
7r9sheO0Dkk3kveYJMsK1PR8byhcWr0Zurb8QvzbeIn+q0hmqx3IbtXutn9W
gyJgL8qllN1VJ4Z9QLn6kC1dWgW2/yAofc7Q63GyW2dqSJaeDIlzYyeF+Oms
F4v3c23BU3qDvfM28gVnmvWLiJZELFxaiF6eAfvGXgh1ppoMO2h9y2uM1NQM
5Qgbs3FSFKcpY/SiuEs7ucNo4EqHciyvgGPjsQ+L4v+aVKqHOi+G5QJ7sxTF
JXrzQ108AnMSZ8Apn+AOAB8SqQtN4lhbMrgcFIX9mR553iTobaN/Ddzz4zjQ
xw1hXKSskm7gUPBTayCO2MHowoYBvXSW6HJBP2NJdM8Nofdr1Ifx8dCjPkMI
zimkpEp+5DW1aoV+G/hB0v0Alvuy+GZS5KmYa8SrMP/h8gfeb8svWC79RvQh
5hmBafoCNDOX91pi8YqqvyPy8CjeFGKQAsF7HWcjmWq9qJugyGJ3N1RtA+lb
Okv4wnfR85mhYbm+IiZcZQK7vN8+FSE9GV2Aa2qpRDLkVLwvcNtPrrtVbL/7
QtVAxp9yeJgit91jpcztM8jo3fM8/v2pAB38fSOs0aJNPiUCSMR9AZOuVfVL
z8YE8Or+IN86OA4qURm+hmjkOa7Ya84ML71XvFP0hEaR4M4z8762OOmlQ20S
t2z9VPOvtm2fLBIMoBWNn5wuOmyknQI0QJXm+2bPLxxe+OQCy0DkvZ3i6r9V
cCtMolYISu5SEeKLz2U8S0GhcBEhcT2No3W5rUktZUir+d8hAjt2YNhLF+BE
vbnX72Uk7tfWsroCz5prd1HWhihCBxUe/m1uM1FoUZa24d0INM4J0rmKQP0d
Yx5482qbdObwycqI7IZ8FgqwQ+K3dXNzAtem7JbgOy9KIaeWsa5IwrdJco02
wNlObZH2x57SIxiCcMttmcDHxnSVvPNQBvcsC7fwSbq/6StGe/QGUJqHfGaq
4cGO8uMHxr72bWFZWqOSLVG0Z+wxeLgfdBdxJ3JvpS0b+Niz3q5TOdQAZjXq
roBjtN5aj9+5mtAoqLCLIrMRVq1S7Jjv7wAUEUsMvaTKycdbMis+K92xKPn2
Lsi4anvuhHJME4w6PWBZ9mzTFn3PTOwfzKK3aIw6e5kwhQrAEGxmb0y2QZzL
nPLeGblwOrvOrUigyux5JMbblNmjGJx/v9gSSVkogWJLyw3HFMFz413q8kpk
nnmcBibLyaSgNcXnU2XdEibYLzhaW223oZLof6y+qOSQWEJKUH7JBjQDsgcX
KgsQI/VaByaL+FmOhk8ddnbUQjATN3Gh+VQn3Y4Tv3hvAGeyKtled150z2+c
44XhsVxIaQKaj/WJi15oR9DE3Uq3MqK3nUYTgfBMC3sC6xLN9yD/ovtC/w1w
RLY3vHWWs4fS1BW9irOGYHkYru7fCvDUFaLaVySULT51za6ZST3KWK9N1iLa
f0o79D8jq6oThEPdIX7RWuESj2+qG1F9N06jeqExiXzBFXxvArDT355VeafQ
b0vNQaVdcTB+rtCMj8wmgnvkwh4tYwkndgpndsBiqG030K7lcuQtyBtmzjpj
mtGNRYO+uk33eQrwG+8RMalfJMm71OeNsoZI2+Wp63XzN7ltLCdI0NxxZuN+
lHOxsBFN8+uTA8xDzp0t8DfCt4sV3mMTp5Ogd/rvGr7mOYHgvd3Zhh7SfDXC
p9Vjuxe3rHOkZaf2aFFpDYPPEBjCK0T6LhkdKssfBByOj1ORJXgAn/G3td1s
sHOYzRMWmxXqUyJUgRFyYKIbsHCNyq9dhBFfY7APuy3Cdq2ESBm22ROapxy4
AT0M7gjvZqNuNW2l7hwad4lmaBzkny/DlMDP5qVFVFcErB7kijWlRdHv5Bh7
O++BljeuiYxm20gniWF9CPFhiUXdJV9dpsR48M1zFuEAJFUK8BteJH0vdux3
YPVCrt/ZltITIsfm0XkYoQIUQg86lp47qCGlVbs+4Jy+4jrwRvV6H2E470Qj
wQBnU63cXYpcf7+UI1vwazltWQ3Kp697+WJnBrv/D4ARqIAN27/hLNF5hYRi
Wm8B80pqq7ZCgz3wjtJIdTZiC9el4wnxkxt7rzxEx2Yx7GhNNQarJe6J0/Ew
8eQvORMwtVXDQmwHh+fpb5XJFxewBwezOa37TPx7+JQ4rcexx+PsxA5Ql3Jh
GMrZgBfMH2mmpHQslrgKR+vV3pLnYS84N0CpUOES5MsSteq3vqiwkRi3iSP3
pi9PvOAzP8gYAHtNPeN0uF41Z4oQr5irgeOdJtI0BhypPeix2zzI/bXSqN53
SvJmZQSgmqQt2IVN2YfsfFw1GcOooMvu8MQRIEpEGZ7c/3ddd70T1Wdvn98f
434XYo8k3eW7ooCes83gC7mUumK88gARrMPIrLPcbbUsPRHH/I1/sMcSmvvA
Og5p9Tu3n1gsqyN7sPS+6j/HVZ7nMxglp2vbEgMikZfeRqIJBepbuSWW/yIi
nCzATMBFL7CqCoQ+FR6USE92AacSIIswS2aIzJbMQ4G6TbXbSB1N7xczcIlX
JHrR/C/unr+KnCggMAADk2si616mKWZn6qSLYkjNvHihvKdTL9vAAUhwbmbx
l47Pgn0lzObbqeXs6hvqdxOz8WZ64JLP8T5d8hh0Zbf0gZY6zm9wzB8Ee5qf
k3FLV79R8pFUXZm8zn489Ta+HCUltTGheSWxy04YGtXLKVW1S1TbJ5icdUx2
VlVc/QZHnFSe820x6yAozzJhQZOkoFdgvJd7TdzpVf+A+niC8irM4NFTlpiQ
U33o04fym5mU4eoodHDEVSDUu9rnWUoRtrxkO9v/UVvTsLx+YRmCjliz4Eyc
jRm/Dzqh7jjdTgcJVURai1t+5lVbBtZ934en6AXHDm8E9E0ziIuNkv3yQWJg
MkVK1vPg0dTs0cBvSA4I2quhqcWPeHhLYGorlOO2x+lotti0d7Pyr8jSrxtN
6b1nnlEjbcUTrdUr+TaBpYEK4fZ5KAFT4L85w1UEBRfO0h+TxJgvjZEHoN54
dhccisoMSJ6Zb2Ii4xThUFR1spWsmnoU31r0/Al5AQSJjRBr9t2sHKAKQR+i
yXZEFcY/mgX19AIOstwsym5cLE9n9oNUJOnljKEgHbdaOMP0AwmwgF2jvpAR
0u5vVAXaskO4ar2LfVTRMlOjYlzcjP9ynDAmiUczYAOoje/ROI/1ZqhFPrdr
9dIFoI4fF8EWqSA/nCH6DEc8SF0HRlAEkbXraO85Ic8PHWBhnr6B0KHpccEE
airbWXs0Bmm2kYjo4QUqWNXKDb7IHoI19KoGjvJSn7O9lGTCDcvyuUAaRM0n
+I4RqahShueFEidOJxmdbNPN00xT1aQfMX3JBlxmNd0f/sT0EQuP4Px7/KDF
USCor9nFlwd/AjC2rsGolvf06RgeEPSBQgPe+igFY5AsFQ+S1qYtkspmFu6b
FeFQ11VdLx46h4ryle2lwYcW6VLgrXWG6tiUWIuASORzKP5ssAMzRtG9qxrx
oBEIJ3me25qpt0uyemc9yuVVuVbjRlTwViyINhDU+vIo1gbnneeK2EFtd2Io
rnQn2sgvjsKlhgJzf+M1NvdP3ocyKNfXg5esR4tdc3aK5nD6wQho/1hH8NiJ
N8xRqLlg3rXXIrXxvJfr6qb3Myc+ZLQvJxQtIqJKZysNjH23W6rJyGJVpsD6
6tBOYaHkdShx7aklVWBwevI5Vz6iwQAzQ8dr+GblLthZEkq8FIxNpj1cY8U5
J1hFUEcZwE0mMcowkbMXoKvm5WVm7JFrYyHXLM2nOaKqBpog785wJ2vjY/Fe
o31aRiDwvuPG1y3Qt7EakDa69KSGiDavRObYUQZtVUaWSxJPNQRH/TkTEzbd
r2BvhFd+YsM1Dfz/tmQd5U6iFL+n5hDcQMDYNEaIPG53IjhIUg1LKMzoAqpC
iIYKf3XRDsweoI8wiQJc0PxRG2RBZl+jKwjc8SBsc/wm0ceymLlYeTdTYTGv
RWhIEI67ChsT6QRVkNzKJHz9pQMiaxCZ5g4QAzw81KVl3Fspn+aHpV2AV+zH
woVwmDNnlROsCvNyTLcr2Z8NGAwX6hV8Y23M9Nmgg/RaU71Kq6IXbp5FROdb
6g+UQUxwC7ujYtiW9YMM06BYeeeq3WgOQ5tp5tYOc1rJzY9UaJztc7dteKEb
qGQB7FuOBR/nhzYclijdB2qIFkVXXvGnd7AwayiNzFS8UIRROU57fQHeSQdi
X4ZrkF6svD339Til8xfv/w6pP/M7SQxEIz+OCAqFdRpWj4AHcfMtzwbMvv4U
N9tDCMt8fiaG90PgQnUW+6wKlyJEmc3hHNXmHAjLtEvgphrjh9NOV5epcpZi
q9GgYOgFpJRAuvamJqUYDGpVkpCVHPzjsF7LSOMlJPzWYUER4et/JPykFhhI
czpwtUZgOom2PpFr80t2vuLpR4orUFOSooGNphy0VanzPC4FTTO9rZ43IUlK
/xeN5gRF2/itJ3xEpXjPTzq83ELPUp2J2HLhwOCS6APKMFs/ak5d9N8eN1j9
dJ8EIKa0go07LxAg+isF+UTrrGNVAxPW4XilJvhLrrdUDCIkkSUd9DW8YL/q
xN8RvPslceYb6M8YDs0W5XgFP2zDDLjZuZmxVl+mieHAb625UbN514/qX/3u
1p0C0e1XyeC+KNSg6FwANgWm4rpljQ99kwj2grLayyELklc153yzl5CP7DrU
lqBXdCuFfMMoO13BOKbhsj96+IAK8wm6SQCIeLp+MsPw/ASfPbcCvaZte7kB
PIYdUygUo0Ghia/JS3S9KMuS6GM2hf2Tqd1boJt4WwyK6Vi1yis2+EOdnCqp
e7pzcL7R/dyb5k5ptK44T7XgEFz9MWwLwRctw4vsR7yeSwHaM13ZdzWP/V0G
+kBRAQfknoIdj8M9W2E+Jk9FWrbK2zIvud1XHerzPyXvrOpOgcxHzri5I8Po
tJh/2VnW9pqOh4vdoXZbvthcl86NZpyXHPYnSq4x76cDFqwcjkp0uUHIChDP
PJ2KPDivg/SNRc5lwB9DPsKp1psJPE1GYaoAk5NgsS3CjJIWIhpIZwyLkcxx
0bO4wUlRpDUyUknCZmqv0Sx5n+oATUCjRx0OIlbX0woI6rCNlNrUu1reqAs6
NO1PIm85CRVEwaK7YZFrJzU2YwqMahDv9/8fv7230VzkSIDs9wZ6L3j/KcvY
0oFxUPhEy7SaCgD3rfAjS6Q1ENexEyj4n83fmiKpCYboZZWa07yBc4FRZ89n
E4ZheqaLGVphi27i0HqEy+lKXUQ+vA2/WxFQXiun6WqMfsnc7QToQBEASm9u
HG+N1GkZnKkgxqf9FoExvs0BgRhMXvFAmG61z9O5tMbP6YmRudQJ2x6ue3Bd
DlC1SiCks2r56Rw+Wm3EobeU/LuNlOy95mkUx7OS21yDsiEdBU0FcdTgR+mb
vhMWvBP+bNFS+vFlbyBplR8YF0GeQ0j9wbt3QC95KI+OWcXF7qNCeH2DrWMy
bnsp6WcZ5HoEitEIe+S5K5XzDT096eyyzWjwvjB7kccT5K35My1z+Y4g3GNn
B3iq3iaJNmyHs/tOHTfqqPinZ4VkWyQirtdnGqYSbXKbjHs2LzHtO/ap4Z8j
VQ6vKbg4PSrv464ILUbxvgLcSg45t0c53Z13fh6xTMTkQewJiC6qcDSoERpP
L68NwNWJlNnk8xmyCOPCC/Og4mM4sXnSvDCuTKkqk5Zm/2DWnFfMEXbynJxR
u0tu1DrJwQm+iPiTshodw2uLUctSyHPqC5fLgNF8yZKEgiB/gE/VFtCIsgqu
uP7yKJlvyldp6ocVNh2j8KeFB6SwIh6935h5aV/yj9Iai5M9Th8gi9bnsBlC
J2nSY8wDAJV/Vrzt+ab0PTAVYXZDzSiN45fWTwSPiPDodYOrzP6FAOPS+t56
eIKynPoPMl3of+IcWt0uhOwAD31WLr1/XfrPGc7IQAsfu3AwpIvwBgNqhhX0
s/YPanRyiyZqPRVAmGK/DNhcZ1PSi1GmV2frVAsy1sYQA9cA6AHGQ2Yyax7E
LilEeRiI6qwmIiRTIaaksPyvEfxBNO94jA7ZcsxMK3rB+27TZSl5Sg1ay1XA
S3u0e8slN0ggy/HN9iiIZjAqNm6hexMb0Jt9XvozqAtpFcCO61b57VOzHe+8
mKa8j6332jVt2Ww2SLsPu/6i5oD1Xn+G4+18joWRPLhInJ5PQE9Sx1oRUV5S
eN+77hLBUwkwIbOrjhg0VTZJ9v1Kjlv98YpDw9LYb/gqEo1zRtAtumGrBeZT
i/2yUu6frkzwlgbkNBKs4hJHNw7h9ftmxeOCK7cD3Pu4pAu/mpnsFfKWiTSq
M4P6zwDAJuFR8LVTJNmHZI7zHYeE0pbsLNTw0utFn9zS+zx6/RgQ9mEuDZ9O
ikMGhy0g7P2OfaNrjVDOWCbRcUv7Up6FqVzAsDe0MFCjqeH2HnKAn1x8ECxk
wGNAfi7gP+C3PH6xifwGH6ye8xvm6OVWsqQ+tmxq9scTXKWUjxoBnR30Irhn
e0jnV2wspr+oFJmPEqljH8o7nHrfYVqlPUSvz5KhA30wW/wAqL64ZY1AnShP
uWEJZnW6COBTHULn93DU73+3lFBAS+b/ziUI3Cv67egflYdcsUOVm4dhopsI
t9ItIfIvH9D6YJ7/5y/yBxJ4/8YBl7N4kZdpRm74KXLyCFKb5EKNIp+wVWfd
QzTQnbwgv5IV8XzixtSCH9tHZXJarF0oMhnfyidYzy8z0QxTlihKF4JDErKZ
xdCxfhp4Ty/XisSfGkNQEkDghj3slfxRwXArgPOrfZdkUwtsq37aIi9a3P7m
PdEVHi/DSBWFDN0PYKRBA+QTmZREq1vFnbQBtB6RjMmXoVHstVgFEOGf0IR4
YySiIPXtZP/T4bB1cqiUbFs8eVG7ESpc3xHiZ6IoDqvfxNoWb8Hktgv45yv+
IVS8/huzjMfAlJz8/yQRAYxjdweM67IALAwAtQC2lU+4qOQ9ivS7DZh6Yqk4
DjGREH/G+uZogb51rT73izahVQsNG6Ievn3voMTC8UQo7TnjcSdN//xztQiR
HyLCqgMxTaYU4LMpL3KGbuCSaYITs9YXVRFEzB2KRZpsQqa+KtoQ/ubdIPdP
Sixlgil7MMEiaHmz4uxM0mryOS4qs+hXEB6nmDit9gJed8fEIbJ8DfxOE6i6
JKPZxlUt97IBSgge76jhccc9s8ygHNpTZaXSv3SQ7shNnPuNRvtpphX9Ynt8
woSraUCKteHfp8iuyaFDTjE4HNGyaRHMNLTp07DIGN6DXNrzzNQhc4bkA4ET
V3RtktdfPvBLdRBhQHxxQedgetZyCqOWt9CEWvzGWteHBq5KTLbjIwDvMpGt
+XmIRPbS0K3/pg55LpAJhLBMpFQdPPRRMb9sQbZOl4p354hzWseGfItnw3fo
savPRPXELxUSCy23VOBdhpVSei5J0qDULN/zKe33rxddEawdBRQrEhovy9Y3
OGN0h6Gd9CGQrr/FMOcodN14kmJuU76qn1ATdWx8rDKk6WIHjtJ99MPnNzGQ
XvIIps315/NgnvAIB7MK3+grGnJiwTQ73kjFYwV6bIR8pgW4OuLTA/3Dr0Dk
BR4dKQNUhujsAa35MPvUFepxb0tPvEZQmL6EUKoGJfYpSKJ4td3nctWswm23
Fu66nTaCEoTGFTX7w6ZcKL+Ldy7k7OdZKXmsAwRYj+lGXlsNSaT3rbXygD0e
ZQVAI8uSgC/Qu1fhpldarMbGylOEpQLEbS6h2rSLzfMb6rskPJ4sZR4RNO8Q
q1bEz0OW1SgwjXsQSDAs297TTeTsoWusMTCaB9g287wStkFnTpJo5+U0dder
eXogbiISxlFmG0h9vCjyBy1Iofx3vP9y6pv7N8q9pZ4rHOe0NUGXbuhO20ZO
kwcuJlMISrCTfxYrxXoomIpDo+p95WhEpjuu4XwFbPCmu1yH6O2cXPNAN2bg
/hUT6f71/qOLWW0gT66Q5N0xvhkd2iqBcFf+5sf6qCQi96stu3qR11h06vqP
pUiJFPS63FJAoHz5C7jlCrEjvF7WhNesE9AKR/xvckuOEFeaKGJOFxN+Z7/o
7/KQnxnaVbdlpurYtiGB7wcUB+ENDzRElbnRNjvLCEOOq37isfBF4zVGj47x
Uh0VhNG43Jg4sl/mentDzpQ+8xGbLO63Kk2dH3nSp3z6TKPSlPClTSAyoL4V
8+lhSZ3MSq9euBxb0pw7ZlMCzR6euztGVqxRH4UFah48whAh5R4j5zPbLUDg
BOdj7Xz5aVGVv0Y66lWQwu7WAOeTeL177xQtVyUZvzYei6quuD2eo+sG/tIL
pPWPFLGijvTxeBnfQ6adBNV4UQ4pwez1WEtBHfmLL4S5Q57YC/PQTk4fsFtq
HxZ+DAEYGUEimjdjvUhFf2xrOPeU9nnqhPkNkYRELvZ6k5wm0EckYUlS1Wve
ACnt9udHmowN151deNNnsVDj7J/Gg8oBVlkQm3Sp540gdrnlTuEMlkwfkZvO
oAASxrDmL9l1lZ4kS/xC2QOOLEdoGahIYM7FAKr/j06fKxJsIt50FX59+JnA
F2w5Dkn6Uib2kvnB0ZbRfIaPHlA53TOWnV2SSvNY2fVEWvmJQQ+UBgeXdMit
7JsUiam3hcuwlEkwTAaAfYYap/5HTuwDvuL1/PRVvEyj6b/Vknmh638VTYWd
10pjm7IwqGOg7Jr6flCDku+YC3SlP7zGh2Y0ypNJjCyg3xMXJWEcR5pvnXpZ
CM3vy6kLafrPjkRUzoc+cxqrfqICJJNNXBCPNiRq1DpFldrVxmMODJtrerct
O5UAHjiR59wtEIBK+Gh6ppPJ2rFqdOLyUD3Jx7188j0bpN0M54WCkPszGwxt
sL9mXaBIAfFxcUyiI514URp5mOP5xiV/dJGkjD6ECkr9HAOKfxMpNI4edzlz
PqNTekHjGQA8zxtAlztOekQp/dGFY70G1a5IxhLTpv7ZMvmmnKtSz8/c/IU3
G83RTDByHxM52R5zduuj6AejarGxGgn8WsolV1th/02eRXlnugd/XmbkLBld
6jL3/GRjYou6hCkgkTOiM914U6OplMplCIaXtgWYyNwLwnuSebvhzeV5ZnGG
uK7bUux34fCYa8sl3W1m83hoEJbEECRXTkjKm8RLnAmqAu1oA+j/BmEsX6qu
xLg2gReZ7IxpZcybIy9N7vAL13TIOBoLhJIDpYGqwgGIR8cFfez9UAVn4hwR
Nwg0C9WCdixsEPNlrF2vHaP5MnN/lSbsFqaRMdIcAsyua23r6ZHUsR+dL2gk
GKzIkQv9cn2un46gPz4MkphjkVoD2RfGs9jubThAxf823XWUuYz9znL7sjeA
mpno0u5QRoIcNcXlL5GhSeskyogM5rvQL1Mm3OlR/tXdDO5jXuc/3zITKMTa
cHc7p5R9H9KGu0OWHfGsIGb6ZTgmN5L3vaueAeJ1T5gzMqzpZ9riD+rP8rPc
CXXYijURFsuqwg9GITJ/k683I5JLK1W8gte77WQwn2vuLUoM6lcfQ0EOb0/P
D5zVsQaKjb9cYw0ib83frxvaaRmk5abbEQtbguV4Nr/Nfgkz2a8TRIpZXOxl
jvfHyRZrTRrqb1yANt90SfTqmLgaC8h25dz0BQOVmaD21iPCTevTTyN2Jd4I
M2rgZumLksAvwhuKB22PnOmx32i+sFxnhTAY/xAGkoZmzAXFgqIQxFBR+Ywj
vhXmBVcP+Pck0tOHmwKQ0ktcO6flXC6cH9HmBMhabWyr+J5h1GzHRErwsj6R
1fW4CzkbVjyh6A2sezsXdxZqtciGDt+p1EOQ3eNoSfPwxn/JcG4aI1dZDT5+
DOwjhDQChyVC2hULXS/tbBX5lB/yNIULInd5Zz2nuD/xQSHERbDI4jLjUKHp
T81zz5mxNUlKegh42514+QskvYYMid+tvM0rk5iZa3YqqmAfIyb24VOon+S7
WONWjNy1VrnZMyEtKiLLEMfu+ALp81g0BqIhfGLRGQsyX7U/qVeHykw2WrD1
AIFWSC34jba4dKFvw8aEfnL3wZPnQLz5LoUdadHqNpyxcZ8j5vGFlmfXe9jN
NhEyNbNgjxSBTJmyXGAmuc6z6VAPvbPqmC9V5IVdNyqZuOQXDgCgPka1ir/7
PEugWfaDIPVS0fM9mcNJ9fQvmcg7POlQyBfCamEx9OglbS1nEEakpAvVAIWz
2iAzZZe6G/bCwzli8RqIoiNeiPbTiisFds5IHugwgaOiUo0UXfLIp1HT+Nx1
7/NxnGsp0AsIJWZDrH2Y4Zhb6rAKRpgVfdeFsi3KiqYdEm2z20a5DajeqQYb
1KJ/82VsMhsBLFnz75niW+lrKg5DSKMzx8d5ijXGEbO1XiVfydPrRgdP4y8o
umcbZecmOb9T21TL69s4MJrzT3uLCzlt2Zlhjm9yMc2edSPILVzGyvSUhvaH
RdtHYknlsd9hcFcPtehpeLwXPrSulmytSKN5DWZno8PWkSQiGdxeHoAZI3YD
M2L/MRqysm5vbmSNx+WfP+Qdrbe7NkHzPFD7JIyZxeEXQEKG88iuGv8GA0Vl
azV5JyC8drJQT1pNRRpuvotd8evre9LX4N3l3CIuZBLIiIcpBz9ki/02oNS5
LJ7vQmG7BZCcMfaIsD1KaWO8k39MbVB+IY2l0nfONGqHfQlaNGC2v8LRWmUX
yQPeq/V6cpbsuFbOtxDvouqkI1IewxeGcTHxP1M0MtliI6GO3RtIrm92UoWz
i18JlyHPp4YuinoCpabglqtRAFlmkD0E2tySdwSeJe8p2wgA7Uw4cJq6oreO
E6f4vGsxBF5swpHBEzToairAF2xy8hvgt9jj4XDnEhUhGZ1/C4JFFDKE1Lj8
y83klPpFdMZC5dVRsbSGVm14nVFy7b3DNGHR5gtRW08KVmeT0B60ZPgTsp8g
xizK2uWFTpcLtam8NJUFCchZSf+6C3re+QZK8MZooWjMLcBpaqw3j5+6J3OS
kuoIwYltfKCp844Qgiszh8+5P97A4sZVywuDGUb/cr9yqVE7xxgMaoft4UXE
7nU3D4tolwHTL+ZN8Lf3Yt4Mdgg7CwbjQ04Y7Jl5X7td4xGIk0digNOiWxNW
LrYaFJNPa7qli0vQHv+N/eP2Qqi2drkBvml/LxLYMEIiZtgxqYRB5nx5Ysot
ptIm4o4uOZt1AVqZ169YvbRv/2coiIVtCzleG5/9k883zZKM+1eVW5m0yaSp
jfyisIu98ljKXu2BLS84F88fjIzCPtVA34C8iRooDSIgzZlCUMMSEPPq4ibD
FRLmUanVOn6DpNEuVz8wA/mtPMOzYwYpuXaG42DpRCLE4vjxLHvFIgemBUpA
+HVr7wjHdpjZEkbiaXpZJWYvQ7Nl8E1f45gsuLxIBwGQc9Y9QByXVU+6YChI
x9ECj8pkzjBBTD/l8HsLItHeIvZMu29nd3S1ZL/Kd1DhrDfVoIJ0HE2Il4DQ
LndjqWauxw4KAyz7csLmwW+Rjy+2V6Ec7+8WGKVUOUQQdDn0rBBAf+mnKbwa
GCyAMDktDJ91pyReBOGBW6hecpmqcM4Vavj4AZozhvLLtQ2Iry1QB7CAGH9V
Tk23nElgvzwbyTeHY9AutJs1uaGtVVQt9B5IwzfTXB1Xjf3TbV0bWBFZ1j/I
xPLFuaICoIYxF2K6EHP81uvO1ko5kjkfYINBh5yB2orgnd6lP9eJ+z4VZjPz
co7LVgXW0CjGn2OnMUkohmJKeAk3XOyyIVFtQfOWf5lWRqOGZZPcVPQeNB8g
pyP/qoofrgHhSCZutTN+pMKUrxh/7KwdjDeRCdTR7mcx6HFTlfdKOoaisSPZ
v7xPWqF5IR/L5viG8/mYiYCwsHm/ctfzi82M35j1WrYC0Wj6c6k5KilGFGN7
PScraEvxiM2KtuVi5U2rIBqW05k5R+sorOwi1TQot4BiQSAuqMSMzMMDeFtu
plXwa1Bl4o/1DdCkRR18Gi/Iq/Uuy3x5MAh3CUlc/KGJXb9getc5CGwBK9yd
03pnzWduL/kcEQY4pwzuWznksQfKHaLIfAxxLjF40p2SNktF7+0PkoPpQOxI
M5tEadwO46S+e2UuvaJIKUSOMvWEshhiFjbq+uI+IQqwslBp6ETET08dlNEz
khVEmoA+9/Pds27rAUAqymCy/h0y9sD4icJUeongyyyCvu3g8Djtht2neyDe
3TnhqLWUWoVdQHlze9y/XUN9Uj7Fs3l5NyMoj7j40pCOWiCVuLIix87s2gda
m8xNLJdTuGOpl2MuRQDeQFiGgad1LOjJqYpja7pw+mg5EVz9oHifllSpCaav
p636rK4HqJyWI9PTLU3RnV0tK/foZq6R9DrL+FowKTmjYs+/PmnhL5V38OAx
0kyI8JjQzAa1fuw75NFqCB9w2Gr2mOgtirR/qaCrSwBYfmlXxK2+aC9X4JOG
KKwyNO3xUG819xuJRdyQ3oneA1ufcXeaLtyhzWI0eE+frTyqG5QbzVohad48
J9r/v3MAc8725ddLakxJHF1i3k/zhOlUqMxRIxORvRD7M+XKV0Dp76uaFeFq
zhlWBZNCEcAaYFd09pV+70SdRAhL7Q+1FYyRT2+4cHznmz+MVPLvWXZ8Hqg8
0JovTDUGkTcFTMPf29CuNJtOaSE/KFXglEtqUl5hGB9/TnaOVIzCEcMJfxrC
KWRV2DX7b3WMsqTRQZt2/PD5cKKr6enjiexZ/dx8xvJ7me8UovystB8D0Ye9
+aet0LjD4nNQiBmcEkvNeLCFpP0q5hqED+zalRz0GoVJhznIZy33Fa5EaXPZ
7zdm1y0f/M7aPxWZJBCjIH9zcrh7CbuVs/HzVpX0WvYVoM4MISjXIPkVgvv9
9yMCb+ifQoYpO9H5RJJUkSlV1PR9qvNEEhULoraMiAoXlZsmufGLa0EUfK9H
t26k4Gd6soh/eSOLsDmLDyBsduUTFWVo9LJaIJfhdLOYWe/ZrKqdvRoYThEQ
9uqG+23xnLu8IGztj5DvQnQec744R+20juN8Ywz3X06/8t4K8xAVg4CqFlw/
DMib+5wU/SNn9XyQvLzpyrBjdLBgpvS5k5Cbxi3LNDT3X8Y3egwXVfe4hzy8
DTPFMawQ8d2YN6v4gXUVWkZPwMhEQxPC/rju3Q48MIrhOT72V4xyCZnBmwIM
2NiDXk3DAlQEnC73tVaBZyrOQz2xB64owXg0vztgi8J67RgZyZYmXMuiHsDf
vGwFRYfG5MM/Nm79tdHkK56WtR5CbN9Ui6iRl2gatZkMP9A3hZ4oNZ5mzAmr
NfrNr6NhfOtZBC8zvhT6+ErrkGoMWuTolwC2QzxEfTlDQnteZqWi9Dps8ux2
Qy5cLeCmIoZ7eo2fHYcuOq+IiPNW6GNFSx5IOSO5Ql3pmlc6qwPveaejOMe6
SK4agwbQIr53qFxRD+2dezESUB8G72zFKGbe5+87uonPpnNaiCJlLhXiJjPr
XZcr5+OAO2RnBfxueYXM8uHjur9lEx5MiPw19ofNmpbMzE0/9XdM2hiFkwOj
bmZtVQ3CQAnFxAh+/ld2NThfgFsxJy4Tb+c4jEYyon7Iy7w3vOR/HOppI7SX
hP1wT4vASLg68RWvUKLc+j/hjTnC0JURMSl/EA8zSX01p0BWYB+a73GRDuZN
xigVpgPCAtIwqU1Ktk41jE9t98t633x9jIaS5jJsb8eui8Wj5R+AglJJ4xY0
dpQW+RAv8GXM561caeDBUVpEM4VXe4z72BbwuhxEmER9osK6eRFpRtFE/qA7
lCQQSYV/GNgTvw97XSPlUV+PJAPLq/jI4T6eb24mhIETG+uglBVIGLE67weP
Bgyy9gX1KlQe7GWJcPJJzMFknSJgy7WQhXf7ymOKIFoFzGZ3Vu2vhEDoKy/d
Wm84ua8jg4SeqH9L5Qn7E+j5FlRwa5gXwc0JQxfxdNIYGFwiy5rJid1+8XNX
ss0GTFnD+xmhNR4GgBw3Ejs2KDgLIl53wniEQf5+dyi7j3zgvfkkON61Y4b3
vxB/SxfVR1Z5sOE1KUOgBwdS1BccJxvNDYH7G/RAN/uXVvJ82wBNZYnKg96L
/W7DcEFvHwOF+BCzxroEZjL3WuUqpof///08dbvYmp8IEXbpGZnsispHQInW
1vHVA5vKqCnh4UwwvhMwV4Cq25XEJU7W6XNVZob1YeX+7GLoyyJx/2AquCis
BIaVfKafWYVNy5LfuPX3TDQwkkpoP+1ntb8l4koRr2XANWq4sQwFKjt9kG6B
efkuU0v9oeJNw4R5OcuaRZ+fPw0pcnt8LHuuBr8CyqbwU/k4dLSZwVLltTM3
XLVt380gTq+0SjX1N7Py5UUSG9d0/3LtPmFvViKRug+jkspqkF3RkrGAkcmN
AspJYfk1c9Dx06zGmiYwVouqXzszwCk3bqOWAao12XKMTkIaam8l8okEhNyD
Z5A7fjWNiyRFm0RyojHGgrEbT//IHVOASXVAlsHnZC1rryerLwoDNfMtDgp5
fdWrm3V+He2wPoSibHCSXpRIIDtZ6uWG/b/SuvVm6MSst1fSE4BFUe7KOTid
XkOUEJeLk13zk+NKfg+9d7CWgn1sCuXk6lVnvqLxjr4LOpfBrE6n3wYb4kgb
T7XfspDYyxypQ4IFX7+0LczzqHPiSCi5ivFWUm05fbwRg5FbALaHjNiList+
nBEOYt7aLXS5T7fTzZGIgfXlfS5AzXDQrbTub/8B2WbiX7E7G5qnFUi+/ysp
E3oasAEPjgcrn24AxRjOhVJhtmmqv3D8oJdnQjvBB8KoP7cmgjP3iIGmulkb
M1kP9SPbZbq8FZrlK6Wfjph6J51/Hue4sXlcQm96PmiZNXG9+thFP8evgRHf
hCG9ntJvdgFbHyOZGSGevzfrWk/dird0Y3h4tEGG93MfGfNSItnPAssS1BMq
+8D75dKJ8KGmuu7jQ907C2a9wKP6it+7LHw5pWpOB1kJwREmhu9cPpdU70hG
euboOUFlzbSmyyj0747duEWcRhkcvnsqWyPQqSkBTVVE6qnAtWBzuvpJw9fI
SZayUID/8Cez01/P7+FQk+lw1LIWa3GW8wdF4+Z8OTrK+25VI+a8JyAQfrKL
oDeTQObCRogT6yEBeu5SO5vdDRVzPdWsdfIZOl2f3cAwhQkNqfQXa1brd/kJ
6V/xAKRe0raM7v9LwfbZunPPzrxpAxmv63t8FOZz37f5D4aQRq4VpEiqhSWQ
sKpukIsDMeEQtx9yjp+859d4MUfonlNH8XhoM6bqbUce/y4kTZjE6LFANawE
xrG9H9gudmXr2OKvaGfOYq5tHJwMWGq1g7nWxRNpHpAQBIuNo+yCr89ES7CK
J+o6zgO76IwI8igIl6O9gOxdzxTTz8Ld4R6LJJL5ImY1z8FnjSI1/pzYQEKC
4OeKpmQAY+DV4D7Zu9wXB0zfIlZaTcqpgCDiLLiDqw6zPg5bZSGWpHd3mbPb
PThL3kl8StbIYA7DnUMp4DyuSjuw/yQskuWmcpdl8LHymi9AaVzoypIVZsx8
05MZQiUly8kRRlsrY9n3UFyfLRUlf4Z42KDB92JVPeUnmVqJwUKT/dO9H1k6
72Teh/ygPIKriUegk09dRAv5AqYtLQo3pcHlL45yhmPicrTXPYe4+h4F28pk
dWkyq2eDEMj5wg7iW/QR/pQ/bmBo5zcaDN0i8rWQtdUeFCdsrDYhtxPIb9+M
7rCi3/HNryUwXIe3R8pdkB6NI74pQ4DE/k5SbXKhc425wQuqcFoKZjl8d9ur
uXPaMXjIKW9Zp4EFvrT2ubR5eWSotaYn+GgBiKYLQq9/a/MhdVJIbaAfS/qH
0ZHtkh44IPhJ1J7n9ChedeXQM+9I9cRpYyCdHPnyyzKlOU75fvM0Y6uy8WCI
3PPbI7u2/VMhbYqft2eBYCreamN/m/cbg5LJpsa0WqXyyy6Pzi/DYJVb5F2F
FbYBHxG9puBuz8idxMaKIkKM06pHqp9AaG24kP3XIAoL1YIROyJeECBnrpZG
MTv4k1Rgd9l5JeRKIl/m9ho2vB5osKBSJX6BnjWAIq3Ue9RwFzMrZJlFG9cE
Ml/eUlTyq4MvMx0TSLtroFtbH2Jf7A7gQAvhSw8xafwSPoARlsMe/nVCfb8a
iUHTwjGAQTU9UeoSd8BHHAKJY9y49kNgq7vQHIdyPl8PugCa/1CfRibFMKyB
xtjbopuFESyYJ9cFva4nenT4YAyB+vf5yvE0Pww9HtFYESSbjH3XF9hmGKd7
mbepsExI0/wdA5OuZD4wf9D+Gl9IYl+zgnCDpGljxZ6CoC+V/7bQcSy4KYdO
0DpfkfUtqMWUYEQePXlH1kOAqsSQu+Vx+r+ZgnM3PB2R5LvhhdXcjn6nbnfF
s3tVud+3HXezxatYd+FZkwWylltalBWdZPRDjQs60bOKhA+6nBNt/0YoFBCB
mNmTZvbK5S9wsqnvJPZjgWvKFXZPOK89BB9So0RjYUzL9rHtXW8qKv1LT/3u
TMUOrJ8OxbbVZnMjfzuCKAzQKwvSOPw4F24+qkZ2jFfQbhh0km1sOP3/KaKt
4z2f+8JvDj5CEgvxTdcuzD0Yhcde+rOoeBqZZNHh4t6X3WJJPFsO/iuiY21E
M/XEi1UrlWArQwuJhyR0mRpo7KlDXf6tSnzfq8iLzT+xi1/YZBcerVE+j1xT
YCm8Qd0STO+iVyy467tAu6q7guEndA55NOTjGyrnv1DDoRr6bUpMGW+Fwt78
oEj1nvjjWbvNakyn7oG+4Vp7epsEfyrnOlrNcX9zwfAoazc4S8W17xFBM5ab
lEzAVvZjMFih4elrfUNzN+1IaoHXKaYFT4MHgi48ojkvrr89SQBFYIVtvrNa
0prX1k+mF2BK17ZsDQHv8fIKy5AKfSrtRScW5a4UvEQHljGW6x6EO/TXI9W/
rum+YBuzmQ7BCHS94GVeqrBqd2Z4bedeJ4bIDeoJRAOkl1OCdj1/k0AyEMfe
g2VAedcbeR9zqGMMytLiiTdcLPlJ+eiGItbMx4p3XNDgfb2ysZzY4ppdQAN6
hZMIoyLRCelGAEjQTVHYfOi6VUzfmlb9Ibj3m+s1r2dams/2ijNkOO9+rSCx
3ab/dmQuPmycg8wEYfAf6DwxeZjKv0fgHVK4aypmhdy2uibmVIo4CsLGoQlk
g1NcXNsNcYW2h9Fx7XIWVJ0vyZaMoV7zsa29fdfaHsnrXwO9gndnXN+J+9gp
L0L/FrFvUPXaw/d+YzOu7Zmb6c8h8U+0j81ygK4/KvOf9qjs/H3ul2H8sfYF
X7XJ13Ya+bb6pl6Bza6qXaqJsof5JPCUqUqVWd9HtZbNa1riFQ90w7W9WwZ7
M7+wpTrQr7zYe+2XIVUa0gN2IXB52lq+0ar4TavPQOp5veYEpIQ81M1Cm8Y6
3FPOqW7svSptci4ETphQdmUs9xCTArcHpQfLr9ipy9eQg9Jcxg0bCSzDAb5S
5tN6tuhzvwrIY/jG5VR78AQwoOIGtzt8YcMKEPwBuaC8QLPddsRUF58+SoYn
ilVaHCWFM4M62xT0z8Ag4lXylgba5TzMDHgHUdZ6uyCy5s7cFVPG4f/rScvb
LuYXMYaO3suv8TRGq4/hmY7NiIVOy2mU1lGZH3X2jcD7s5jrxFzNGYch1D78
BvpvowJpxajEiGY+pzN7NC1Azp1GDhsiVlgNPgdIdfGEeXY55TcqaeVX6nis
QiWxNRZFgAQIt0IjFldjtwgxAF/UK6f42JNmN4aGo6yeHxcoqze5gZUKbUrh
YJmDgDxy5glZ3S1bOyvWvC1MffBj7uE5K5GgcdKGPOSJA6sN9He0Ubld+xHh
Op6F/f5T2eZHvLH2G0sJx4eN20M1AJxKv9SJ0O0oQb4wG59cxwDnS1rCv5Ab
YS4vOZKCH+YSD0z9a7UeWOCLtgrmddTvfORAG6DE40k96NOJrpMgZ8cPi91S
pC8+hf3A0+RVKiVXLZFr6G7BvTZb8tRzZ3NJszp5bLCmkGwFSxWWliwCA5g7
BeKsgtYcHC8G5gddGkIrvp5wSAwpRFDtOykQsDlAjPfKe1KZqwDyoONnT1yS
2TQj3SzNph7dGBUthTF9f+JrZ/0ILyEYyEz2S11wtzuA0ApZR5Ihy/doIIxf
U9HjqVp2aKRTkXNDfx+EC6qal6giO50pFcI3GgXvg2dECb9gdyI1M1XVf9Z0
6aUAooQgbqgXPAX0bH+G8HArZ/zk0pfo+rZENrDUdN77LmiWfXMt5AEAMxlh
mdWZq6vFPYlvMw1GflnFXeN7I2lnroFKBepzBySlJvWLfmlzQceQKiaJkgSf
MTbEa68AE3m7R0EWxrNNjTAiOV7PHd3sMklodl+4EmtO220gUrw1qietNs0w
gjC0ISqAejXrKEWN0fwB6MWFe8HTHUBoD/4fJrBC7DFMyc9BASgy1aBgl3pQ
6kzRFsvd0+XBFcgH5TcmRIfBUOthSzC0yQU8ohYaFnkM0AwpAQypdotPXrrk
q3Ui13za/xR/xrOTkmUIRQb3uogHR+wDvNaav81t/Z17pszs7Wdn1R3HfGLA
ZTZHobMMMYd7D3KCzmGPIR2OaF48myEtqGoZTAPVTte4gV0VpxJmkmX8aTjg
8k1G8HeBP+58br3nVnD7u8PLk4okXgChrWnY/tNb2dyDgoqWastxi1MJ0jeu
zgCNonqflTiBjzsEoMVStFlABBlB4uObujkrLRttAuQX6Rpsqn2S/ZODCJnA
X9xTvQ1KEAufzCWhMxvkLsFoKE150HI8Y+hGifMu4Xb2V52u5I1JomVM5hNL
uPWsenY0wvTtn/rebJvuGHTkB2mj5MbwrDY4r7PeN7vGWEocBlaiTY5qjVZy
18jLoLo2tP/vBDef/+cCGmkl5bDRLoZCjPqu8ip9Uwg4Cm3fK9hPEB7XSK31
DdUbjHyT3TW5+4JtLXPBbU2gYZMfNbfFddXouvxDHdLUWg0ti8qzHcwXkPOu
o3yMNRXLQpJu8RfbWP7bWdt+ebS2wjE2nR5sPe36S1y7qdD1cQZA8lA/08Qa
8fkst/AS2GhFy4eNjEGYTDn8A43vIzHA2Vksd7rPUNMYk76kxEdARMasIl3r
0kMCDTCO+CC4gMO/+q/e9F2/j2CpF5O52dyYfIL+38j5rDICotm0RP9DiIRU
t3UZPoQOdVn05Pi1np9Uv7OX0lpT0lhwnC+aDAcIatdqR2rzhyixwpwlIIfg
l5jR9fma4iOK4nsVv8FZ46nSPrtTh087SNMdZQEd1HsF3yYR3qrPF+qCEzb+
hQA8YFy8KOviUbiBxjxwrti+ApdTjkoSrZovpu7hgrWHsVDXEZNCqDyi6mIq
DewC/URf14oSIb5cRC6I9iDMuR0K3XawllJSom/KPPfkJZJtIzLvSYYCvatm
SVnNPPU+mzes1+CXFP0qIgXXX4vDBFL8NhGx+9Ca3OW20cidIjiCUF/ys8Jr
j7MQ782AcM32q1Sn50I6WSNKSUFgz/mY2V5ijAhjbjedk6meJBzcMjU22XPM
8K0Za156Q099K8HX/D6tzafXselLgBo7eXK3sow8PXIRqH5fAY56dKwBwObo
iiZSb1VimlhsWwLknQwp+ulI/kCy4UN9S8+TWrK2BrSvQ4ctxpVuWTB/+MsW
njHpIO/3Jx7JpJZ+bb9QQEuscSmkAiYHs1hSOCf1pfLRTclUoxCyioCWHLrE
ltw9nk90WQFWsES7V8MlWfKgJGbqmmb0v2dzGJfBE2itwwyh6imXAJN3iS41
Iz6sZ7gYgDmv+lLp+sZFxXTtX+LkYcA/fgXrACHQLuemk4VVLzuAUFWDDmf/
K5bb9NNLrvMMIayvVNR2z0UOvDBgZia0QotvWGhEAh8m8onQgxnZU/0h8Knt
sXR7Ime0zfO4UWy7CXo/HlY/3HExYr5Q6W2HX3pRbNhvHV6wYed4hoganvWW
c+R8yPVljdJOBOCPETrLCgkWegyw/FbVkkBf92C+X0LkeOGYlOClHYzKM6sP
XaLenqW38w7gGXIg/eMQm3W9CZ3IKrrrR7O0cqbNQ5cYT4X8jBU9eDbGq7kd
CUQhtyq78Xz8rrnTt4BcNPmpUafTkNDUGc+nFTnXhUvkIZzRTFAJnAYUyEKl
yeEbS4E4yGw2GS15TqVzuZJ2wtKEmNR+lgOFvTLxH3/31T8XHzZZQHCElZ1j
C7XeJVGoO431A0KDZQVSLpQfBP2gg/sWKLRvEoBV1Y/jdQXMP8pRQtYYOMD2
SHrgMbVzeEul8XYMX7KrFC0WvYgoKdm10ALVNWSzp10YhlxxM/pc7Yg1ZB4H
yPrLG5PeuPIBKMF0ir9Iu+/Z8Nw5j3rVgvXBF1wHw+R0jt5umvIEv2uNkplN
HKy/pEDELFnBsxMwFBavdX5m9UsGV0mEMqJMZIrZlhdaZlQ6Omj1vPE38Fmu
eoe66B9ZYSXhFGDw0svOrF59n/ETmildCN6CxpbPK/FW3mJ8DulTuq55XWyE
54dbBsMePaa+/9XKSZEO/ritjHI1m8x4pqD3Xk7tJZfOqBpBeXK1n4vUzsEl
ZHVk83xlOrFcTQyc8u/OPdyr2D8aB6gOtNdjfMT0aTuwzNqkXcYnIshN4ly9
Ml5ZtlYUnJyDIvrQvvbxRkq1TFg7+z5jvaMLAgcWF3a17WiJKAIUtu/j1AGZ
XUS9wuGILpoKoO4CYagsoIORH6Ozpt/1HFHiosTrRsBo2zRlf6CDriOnVqz4
NhQsHY7WBR9s89g0Vflefyzt4rfkMmFfeqSp0uDf64ZKL4LePozv0WehEzkL
fCYmiik7r+1JWvpS6WtZLKdfAwtIjZFqLhY1TyN1rX6d8JF9vJbGQ9Qf2C7I
VcJNtOYhgPr+L4Bd/ai2OdCH/4xtiZGaqFeaykCUTbnouYtcPEnThJv+PR+F
cGsuyIHGC0WDs/dVLh5CAo3ZkwlGvGppiH248/hNcOJw1HHBIFZwGr6Ii5SA
6X5bdfFJu96ocPfDH4NBVowxx/JS8AxiNYQ0eLtNeRRVxXcLPD8N6dyxhIF3
ACZzKnn7JV1Z37ES7C0e2UYH30b3P4rjf1YvdULkTyaIkPnUVpXzdHbDqsda
reuSxFQp/r6hKu6fWiBzPBLhzzH7fkW40LqRlsp0sZkft6Gm21vW762cfrvT
Y9NHgLMHT9WJj0uIGUm7HRTWw3hVuLAhjRmL0sN6o73EMMqukhHwamiww8a9
xQT6iPfZEXUrk4ZkdPqTfo4fTsFpo1ainBsJu6CLqBafBq4i5cngy0qfCHvT
E76kxxpr5rSmqPV5b634/LnUPzCvUXOKvT+Zi4tYoDb4ODOrxobzYVgYA2W7
UEqWVz47m/2AkiqwfvxPINt7z1ayKXVJJujd1lOISvg6SbHyCBJrHAx2E05t
IMeMkeEs+f3DjCjFX4RqhKOJParvBHP87Bc5U64VjBETY1VQFX0YNijyhD19
1RIFa68V+7nuqBTCavx6O68AU4hFQLiqJCIRud0Wy6o8kl1c2On6ZIRkPa8B
yE4oVrYMSKRdKdjJfqx+LRfOb2R4ZuixMxiiuAhSfDuIQ6grTu1EuTMS0KM/
cNvY4SxvRn1w6McfcSawcq7bAz1US1ycDBBZaWYmDPzaDG9w5bU/EiQrrLaH
ZbF5+1sZkmaswEwg6RLzvIWSkRs1ZM1yzOKA35qbU/Ch3GOrFZV2qnXpB8EE
u6liK4u1jTXOZ+HAiW/Z2p6tIDVDhx6fDOHJlnOkkfno+k+/KVQwP+6YsYB6
aNgxXK9PZ3SHbNgV58xqMjOsCstbvmpRgI8pSbWVWmQscph8WYhavu7G+OMi
M3vgjtp1nIurUc4rIMst76kSZe7DHcxkgyT4o/U6FzrocRvWDbWf1ueEP1WU
4Y8iEYU6oOWPaCyrm7FJpnzCa5Jz9uIkVLAFZ0CvVLubiHK0Im0D1eY/KLnS
BKc2pSwcyLrhuQnhWYZGsmwYM/3qsgxugYR872CnMUK1sUmeiT4MnQVy0jRD
YVP/QGmrYZnb+MHFDIAkYxUjJ8nnSpNBFLM4+jLSleiMlj/+USVds14CfSqT
4QelKsoJ7GKprUi0w1UAPiTc9vsePN7NduoweOm3OIDQAn1bM22KDi3Qw/ki
NkDkvtShAH8ZguXv25Ac9bHBgHzQ1D1MaxA5aeyaguL0Wc5zU4JAh8OSzPof
uPT0O2G9WxAWUnTYJmSWN459qkvhmdxYHMOfaZgwkaZHxR5zcJ55fsqpYpD9
bWP+MEBwBi604EQKuu7Wf6JZwKC18XjJ03gnR5aOZmmSzL+LGXmzINY9Qeru
sbp+GXV2AyFuO9EsulntG+FgmAOVojzTPZFr30mj7NpfwjBdqN6bxbO2RDHW
sXduBseFIx/+I8juXQyyaTTgIZI5IBykh0/+TyODjGCRNWVBBrMxuf8s0UKP
YGwElpna9ChjAohKORpthaToVig2NNbLLFTLAgpWbul8kHqM3xy9liOcrwD0
7QI3Jd15Hg161Jvk8oP4+EwOJgdN/c7QryHmrbHLhF+5Cvbnq52IQjpTAimT
Dde4wH+arBKZcVICKfwRKZTdIBHe1mOPzX72IO82Q8AyLKTfl9vq8DoFx/gh
rPN6CHayMpyykdBGeSkkxzd+/3bQjOWD3FTeWKIM0hudxeo8hPR3OIHpJgCN
GI1W7jmnVingw59mntup8LWTn53/g4vlTzRf7lEvtVkgLTqnJkxE8pqXBiLR
rxe690aNDhdU6nKVVNLjHLUVRlsFMN+sddXdlBLpb86eDhifQzBN/emeDqsy
jHQNbaGYN1+YxXM3HfZX/aoXxwkrES+ISfi3qWQWleknw1GdKsfagaPSf0+B
QmGHtCwtG5bOnH0qfgwR0DFkzlKBWDXHk5jUeAIdrkXWlGOi7QLqoB2u5eNB
YgqPEklGj0TAYMVSHqzx1ZxRr4pX94otE5QhA23gnoavrBFsEI6yHF3LaEp1
CYHc+f1xyZrtSmEFd6v4xmKHChSfkmRaNPGuySwmPA0V5gKn6OPqjEJTEP5e
slN1wKz3fEQC9fmO4NmPKkXgxWNByjA1WX/xYSqJjVppkrR473tk424VVcfV
NJAP4OA4wjXH5I2zGH84CXNSe7jpSi++BxxtNMmD2IOIMXOeIgSB/A+ueEQu
2wVLT87OqmufULJ6KOU3RzMMBtXTpB+ZSOBlgUFoYE/rGu0C4BHthZomtJ80
FyhT6LamMOSxBNT3sY1z5ffRooJqlmJ9vVosZNUJmReA08JaoBEhkJ4Pdw6A
DT95U9W48bQ8MyjTS4x5DJgi6e715CW+WhIoO2gBE0UDMmi5RmYuIx0NDe1I
tk2xiJgzTUp8/mc8+yca/ifW/5p0/B5KFY1UOcXTbHtjQJkBtU/quOj1+h83
q/yyg+GqBKdSO5JcfjxsFiQUB7GsltU9m9n/BnByKXj89MyrKguUUQwdIqe0
0Sh1JhF5CchyCpASpEu+HrKmioUP8U9AXO3DqfjTockFbEQkCSBQB/AIk2se
Ylxtp7L69S0VZ1Sz89DcFfkDeTLGI/EFAI/63PxwbKid8bhCeRigy4Sd2gtR
Qa9xH6FokxjO6GJ1x5bO28vWXSYJps/0+d2EL+bIXnREZF83KjNp/PD59Drk
kw+Wd3J0bwORZnknaEuU6d1lyVvQdKwg7x0HfBoNgqJan3pA1iUwowe4wJML
wGPUUYdgdHYxYuDdUT/1WTpr5iVuBp5wy8ahad5rPdozXUN2fkHxHrKQ9+i2
7dpJjK50BtoR9OpduVtDt+07u7wqZ7RegaFZKZHcTCj5b3bBz8IJDdOvMeQy
mxDr7ZcZfBLQOx1RpcJPAieOez3LRmqjgDooyVIXCKEATOs7oc6tdOgsNDnL
Z87T90M1yYQZZVJN0vyrOi9XucfA7rcyuk7VfqU5QJ6ZNZJtxedO8OErp3Qv
yw5meyrnU7Tr9BYx4Eh/m3PH31RTpveR2p8DNvfrtqcnFI2AWIWFocfzd8kc
raF2vOvmQrRc2BCC9JgaogbsA6mXm4kF5FEaX0SuR6NxsanMBO/odbZWr0Tx
GDJVQ3/tysx8Tau5MTQ2FdqMaQD0Ag4JnEL+fhIchKHG8VqMLuoVmDJEjWpO
O43Rl32skThG/ttEWug3db/JEnrte2S5Tt1PfZrdGM/alg/wX5hVoO83O5WH
puLJv8/aP53cEmrlMsFBOUY2REBfd1zcSAp7MAdbabOzsFWqOyTt3j68GGy0
A0Ei1st9aM3dJTJp1xsS+ybnSlHTiVVMLOlhyf1LmsH8fJ4LDMnpafEO98fM
IHqlMtSwZG/6tYvpkVs+S2nHe5WM5bbh+jusfJYLouZkSOzDLyqFFaFPW/KL
Rk9EDgOt6E5rZMn/pVH+acMJrHlTGXsl15RfxR2jnabDe1YbSwNh/PIVU5Gt
g+YubShPfCQZsiPXW65UxyO90EMoB0rkDby3yVRJrvT58N9O4ef9jvl2iF7i
blr6CqladTZ7m43a8NI1WOVkQf+niXWblV8S/qsLEbArYgREk7zfxQTYxm/3
D2mdQIKsa+hqJU6ECWuGsSN2JP60eYXV5isToUSbVPNXb4ekIsHxMlH11YbG
0C7MbBZSN9caiL2GZIzVu570i6Jgw8iA5KmE8+1fpxqKB3d0VyoqBwYch7pu
7gX+jkS/1Miw5o5vB15mucyBjt/BHd45p1wuUOjdbO7cburlqzTyjvtd2srr
FtZSrYrvU6luCtMv87yErdx3E6CZX2lLcQdq1pzBmD0zvtj4i0JgxskXTQDF
WVNzEg0ZapJedGOaH/VisFZnTnMAyZFzl8WljOLdwiAIcjGZkVFryYKKaW4b
LJF/empJeWplau8FAXLU4j4AjSuvGFOYKP55BL0ix0EGljKB/G3iqnWLL8Ji
LUWPjnDvre8uHrfyoQKWPdEsrUVqCEx55ZMux0ml7826O5y4xJ9HIUP8x8oe
A2dhbLYEnOKG5htFnXU5gcXxP1nUx3eLDvrwBZcTDnhdB42/jwmz3oaSsicZ
HKeipiuj+W0PiAoHgJOFwGj/ata/7VLV3jjZmZnLkPtPG2tj+Tkw8jbxBXUg
cPRc++HLarren9tuZfV4JXBmkTH3Uyc531ARbB7bMI+9C0qQF/Elw6GL/diH
eoSQSDpZN5GQu0srFZKDvfemeaA1BoiqiJ4YIpyMqMHvjAzY0lVJxRPaSA8Z
mgP/vfi6yyJ/NJwSw4GR4860kqS7dQxVYVmAuYx6W+ymuAuEVsxP96hmrVjU
Fb7NxwRTVceXs2NOa8fQ+hlv9Oxho2KwYjQQNcAQmgHuBxoeGKOkaF8NTLbF
+BjvFFezxfJ9BCsDwVlt1qpdcXReKFuE1d+Ca5sPldNW8X/ILImMtbloXx/G
329PBNx/wRWOq2UfbpevxttQynVj/RtXLODM3yyhsU//8l8nt5Fm+V6OaWxz
lAZZ0lmDoyPqzQCw8cCebAxw5lDwFO17CjudSz82cPW4s4W4ve4el2WRwvLL
UmCyl3ceND/kF+3kJJzeOuiMk18Focg/cVmpo6x/+TLrkpw3Rtbu07TDBkHi
uI04Y6XXk2JeECmtKNjs24L9JYQ8xFtSFSnWBlOsXpLyWe8YlIcngQ84/xQD
OUezd8hMaeEZVcNym64kUaDlJ5AZmB7QWM7O2t5s8fi+7fc5SlOU8l+k2Z/W
ldz5Juru88akQNXPvKCR3haN2Krsl9QHRLnhS0YNIqpPOhxRdxSBi6n1kbki
2F3M9HECEQf2hBQhyXvJH+9oq9LNMAxsJZopiOZTA23twpP2uqPsUYJAH3Yv
HtEwBa98PZBtEaTR+YLVWMm7wjKVqWM9+POBC7xc5qUXjv2MjmpP3fVdDtvl
ymyYGKqGCzM9yxk0BJh4lUQLXdDOwgb4EDjVeh0zK0weL2jvxMqHxtT2lN4C
S4yyKPo1Hsx+RjgZ3lbD6nAlRQjv9MxiwbTMhM3aHXw/sx8kkc/nET41VjdO
7dVx9VuY1eWjzoY7sOT1G+rlPAlRnfVLFxsE9eXFS9rnFZNagvlEt4/EtUim
wD4qL8US+uJUM7pQ1Tg6tUI+Jqw+TlmSEsZ0dOMEEenL2WDHQ3JzcEGE5AG8
ljub/59RLmq1f1GppQJbB1aL9XRu88ACA05KZQ4GNZ2BXXxHuF0BW5NBnAbU
wuTVd2POzMGeCjVFYM2obxdM5azTjramkKGu9Na7u2XuONLpCHv8S99dxhgn
nmT974m31+wAd6Xg1xPWiJGIsZBA8IsrjKEAo4VacEIjodtEASD1Zvs+CbZi
alqdjQK8f8qtJHrHLp08fFEOHNBSBm22lzk99ignNuAJCHU6d5gE2ZKC5UtC
1I1IcjgZHMq72nOfzDztZbcXXCfBjTknspAezmd8IfONjnfyYePR7hutZi4I
jORrxBYI+7OQDvalB1y02ecDALybuBdwm0NNB0eZpbwyDxFL+ysj5UqjA1QF
z/4DQjAL0OHaWeg3L2Sp2wsoZWZATPNsLsYVd3Ypf5842tkCWCe+quuT1EXC
QZQJim7xq8/bRm8oSBLKkSrHAYnNf4u1aZb2yEgIuwqe7xwROuOuR5Tog5K9
vVcVnDG96BeTNP9DjRPQznqgRq6YnjVPvzIhnmoBzmbTtItfhLRc25IxvNas
pjEDvW/UEixcM3W7gA4NVlZF8rinCxYP3UNdu3A0qcH/nUwCMzu0cwHPYE3W
3IsyLK5KGPp6cWEpw1sxh8lAtYky2KOHaQAlLLy9yiY6G0z0iDvK9BaBvFao
HFnxXgTy4pfMMBl2f0oGhJs7+brxHOh1vXV09gJ/cPeP6o+tYrgjPS4DFAmh
LbWqZadckFZVsmKDK0o9Pza46AJUjjO9QoU63YFgiNA+bDZu+47XJgrYCuu+
+cFjgpD5/jKMZ7/8AdCt/FN/c9rY0g0PXFuVh146JzCjnJT4IHWElu/LITly
0IePRchdXBCYyhSDwsynPlZOsSi/PIK7HG5+JNPMWWlY1PXmwJoeOelE3ktQ
C2Q6rK+ePukRyMrwQTLZQlGuOKibsa9RvSBvKTKwy1UJxicJfKTXcttoTwaY
MSeXEb7O7Q7iKtzKLgeHufP6DBbn36DpW1GsX80VF1ispbaMHC22z8pn9xIf
BLwyGoONkIrx7yLWhcOyJ48MAsgInuM4aLI1jxYDWV/+X4WLkLdzI0/m3O/i
bilAAokEkuaIjqfBJF0ITE2El8q7pYw2RPzJ1qzJhGBxItEym4yEPZziyyFy
CdxOq9Dqmi9Pg4vjII01JJ2D235U0HvgAiapKZG1Dj04dVn7qlaysq5oxnb5
b9rG50sawaBXAFZggSxmpoXFFfTEhFXBrnSIa3zgNwUNBWl0faPPIKOq6qG9
sCF44Lm1nNTtp1Kmj3v97gQ/s1l07EBmzhDDpAH61DH3PMgcmEAGSUwZ1W3t
CM4Vh0xPnsCiqovr8UH4JRducEVevFhssiZWD0+mZNtt0H+CcqTTpZMqaEjZ
5535IEAyUfiBtR41TjSFuzz4ofQAXT5/fXHfWh0err2ZIsUbuFHWRVr8BbNy
WzvyPgIGcLS/QHf+DsT8pwzyvxDi2TM8Yss9ssKqyIa+A0bvavsP5RjSqX/J
Vcrb3/a8lFlTAtRRarJpL6lbfvvjNR8l0mXuJwifEhOnvWf4H0B2CtjnnNIC
8g+Iq4bKyk+8VB4HMb2YLAjKRfi55bWPeC/JWiFk1PJI3fkzVDJ+HAlGNTFx
/qP3h3iTDE3mjd3hda+nb+kJFSHH7XKKrw4Rq9z6hjZccI7VsmzF8P6LzTbV
S7aqmYXiZlk0sLjEdMds3rBQ5w4Hk8PQCsRu4JhKR2nLq5kBQvLHPuz8FTT1
WrG95bVVcTnjkO5OrWzq5lUv4a1y3w0neloHrfBmYB/lURgpkm3CddBL/c4q
C0zzZ5+vvxqCdzECI7WQtXyzT8ZaBty/QzmnrwD5N9Kjro2fmUJWbrSupk8V
9l60llllSzwj1ookCuJWcvrup/RQz8L12D+j/m7Yrusqog5t8myghBAZfOJr
QwyZpWuiilstPn5G1R9KHENsocnzYFPiSbJGDruR5t1/cZb5qhWPfCELqErL
GupRXRkOdNsTayWlWrUkZpcqGC4lGEq3TMbzsNSDlljw3bovxpJVaa8h/1we
I2c/C8L1NILpP9CymSqrenu24s4dLGBhhtkAh+qzY5Oj+15YGirBSOYwOrIc
Uk5GoVg20eycVGyEe3eMZqUBlDyiVhIu8Q6o+0hcy7O7Rp93QterHstCNjg7
EsPinOJduuNs9qno6fw03SDxOlCXgjpygXBnXgmKsKRoVcR+sPEictvGCr9e
vyboJpDRPI8EB9UrKo36TAgzOOOsCnGA0dsLI9H7uAwwWIsRZ3b1Ee49Kjt+
CDzQbFKWLd3P+GsHv2UAPGSMeNLZGXKzwW5j+G4+GL20afAD/FH4+9MhueqP
WDfTY2K6k4pOuv6bTVkJioBFUyQlOHpJKyZSTqDBHS7KnotVFO+TRVgu7en6
YNAJ/ngbRZZU2jSXnCOxu8WJslDUY3r+bWt+TqU+u4yZguZBLXmYg+n1pkoo
OgzSs2+QOTrUusAlzAsMdwvAViZ2lD9VVTNorWE5GPfdFC5SM8OLm9Py+9vz
eh0EnQcCEaP1oXqzTaWumr4CSGxYMMhz2pR9z/jR+3Gww/yt6Z3Roy8sG6b3
iv3vMPLezdS+5I+JbV3NNIUx9OhIXbW2ZFdAQa7XWqgqmamb+WITmQKkhFP3
dmXB1TXyLxmXP4GsEQK2JKRto79KybaDkRCQXCkv95SNkw/Ql5bRZOHXdn2g
mN2N+974MS1jlMt7mE2Gu8KpC2lwyueMuU8cfp/UDXcA0f14m9KmM8TjrFCh
zNHAm90quK5iEjks+Zf9YkQwvqQB+qWZgdisKbgsuXgzJDWQGmC69Ns5yzZi
3b7wZDMkzVm08oaouEfdCw47K8UJLt16UCXcVhQp+b9CA+f8+8KcBE1s3zAV
++svlNofJ/F9kgAe5zvCE5vAyANsRqZElNVhFBNx95fiwBQcgp1NYkFM94bM
CMyc18kU0Z8Xs5gYXbXfOJcYV+qmdKJIhO6xQo9eUZH5m+/n1W2McXAGrRnc
jK34TeG7f7PQUBdcXuu3iUxe+/JIIygJH6XUgBUbNmqD4Hq+eZWV9EQIJsO/
Ns0T4sCXUN9iOXp+PF+Ad3j5shGudm2J9V4tCH1aN+z+PziSJ6wthRMkzGpj
hvoxBTUSP6m1kM6Tu8QnAy+YGV7wDKmy6joKOHQrxJ4seETfyDS6PklW90E5
RAex3o+btkzV8JZlSyOTq6ckboCbrs3Y0CEojwTijBxc0ipOSnqct0mgzk1I
u3Uf4Xghwi3QhJbMXiLmOEongQpgD0IqBYGypuetukqpy72kbSKOUxOpkfvV
Zt6kD+ZVIQa1xCIwRni2mhauYqjUX0X4MQZD1QYYFIMXY9RdJi1NCmx5n+Kq
giTYe4plWUYL1GPJVoUQFHL6pUXu0O2G4cVFQ7ZYIu9oTXIZuLPDMjkTUjTe
1taK9zBwZZIV06L5PJdSHEUDcZIIDZ4PnCq73GxCLAg6TBQD67M7Aq5wXPik
F0lrjGpb1ij2kR7bWADfRX/I3fObnyXhaAU93vnIwP1NBjDccx4G38Yfxpu4
YgEskUp4CRyDGvOEIesZ3nbfjkiiiB0Lb0RTc9iMNyRIB4xrlknFFREFN0CY
W9mPaxycrmk8QdBSzCkehDN8mGG63C552xb6GPXrXlhVfWUgRJMqy59MqeQC
yJ45RluKqF5WJzOcwmnKy8w+lyftMOUwcZuNeLb/VpH02PeuNMJMBU2+WMxa
OHQJtVQFbInER1icWZrreWeH3ycGZ19FudS/ff9mCwPZ438JhFNoqgCP3pya
65C2v6A1YhWGerfGzSYWllpHSe9ocTtjaY02Y+Ac7rDcXhh3IXGtx7jivRvX
8mvZgEF3m9/DXA4zD0Ucj9fT87Ue40kLMDPLDjMON0jaJnfZaWtiuDz4610S
lis/ZEvC5zeGgQw6zGLLusAIaYr5NO4iQmI7AWmN+0/rzT36sYy47BzImENP
0pvxJTl3cF1oa/wkPzRWxguDfmpLfLKm/hCHs0wzz9gqj8izpldQ85khkGA9
MTtwK1PsqDvfv2jx70dnvqql3NpL2gEulkHOr8GxOyN/tQEY3DDlJGhCzGOT
qoeoiIsqYSSHMml1JQubCfAVMn+uBjA5ohxP9ZRpsNk2EldQE6WiYAKGUDqx
FAB/9rHj+B/3z6V45keerz1z0fjZVKp3IIFa/8D0FU01boGDUdpU5S0pMz0o
J3sxlEs1d0PWyG+ei9PNEz1RSvfXT2ZYvMC85BzQK/NzrgSVA19ztBabLj0p
TqRCg6O5CnAzLfyy1eegTAxPLXZVloJSFdl7ebPzXTp/OE9NjpTaTB63hQF1
SJklGpinQxRV32oUtIFrRZWYfKWVmhTst1hgufCt5lyyougjkX5gy/xnHdAY
Du64XcmJd7FxbQAPUceD8nF2+1DXQXxgTUC+8oV9fRLa1j1SDkBq//UgjYjw
DejHxHwSb2tfzZDgDQZ2aoRg8M+tXPn88kLQPjiIOPNH64I228BzeYg0kCBj
D5aNZlpBdo+3LIs0lFm7IcFc1C3Nx1OO7uepMbMGSxv+QlAUHcZC1PcNXOsO
GvAcxCyb6xTPjq4fKCHcOTmd9SpdrHDK5Ql7iSZTB4x9Zdxb37FokA+UeAnH
QwWjmow199wCBh37gr7juLIT7Fbo38atek4mCXb3uyaADxbnaXpw4BMS11Y3
oq8KuxxchXOnF9qDC4ijKgk94PICXvIOQhXBQlMc9KErclD52EljnUPT0ryQ
rADkmxm1KbkzEuM/1ddgb66STYzqKp2W354W7mfuXfHXUIPX6KhAVN2SEr44
8cHH4HQX8XV7Q4+dPMe7pxOg0D4fw2vxCNdf1aQknt/P1kqP8QxaHNXZAMPD
P0Y6jP4MbRuL5BOiFbejD51U4+3xZicWpp9L4XtXDXKmh/yVSWQ47ceXkkcv
wKPmd2E7KocsMFs+T0C+LSlYz/Jhn1gVjX1a5/32y4p/1oRNv9NCTLObVq1i
s4+0IH3QnSxzogLN7SbCxpNnqIqecy+FytdmTRaGx/ZkdOOzh4O+mnnns32M
89USzXWG9cvhTIk2ySL5kEkpn12Hi3vTZjONM5Jx2eFhC3vnxajbyoRHPf8w
44Ct59+t2O4OkQhYP5iilR1o9xX5qELRrU7dNnq4A3Y2TNdmPuyKtYY1+Ev4
zijl+TGDx7CTyc5306EaTJwkZ5uvCrEqPt3FRlaA4Sw7qLdtaQWEsrT0Mj7b
oAsYkc/a24jfHONXVP//27Qe4CJYRCDhHjXu1bpGPKXK5BkPGL6jE2X/9Sqx
m4R5h1oYIUdTt8Ir+02cr1DkFfZR4SAku0HVbIBxFCg3QBolzVOIhTXfUfog
RdDtKjUOyTTMAuClLKH2f3jNpCgcwFJww8r+ed6DBkaaTWYhiZunzQrJrRxD
r67/TTuedr+ilMTvpIkiCi2wbucqHyqEDnpoQ+YFFNud5Jt/eLdWLC8e4Gya
m0I8wrDJfMIQv7JA99EvjDQB4BWrpT3urncwwYKgXCDYsL4389w8HVgp3/qS
33ZEh5v+irp3x8i0NPjV7SiazCoHJDWZmL7r3a5e0dbcsSIaJ/olKFttjw36
Qu0SubFppDEPTnl2B29c/QhBm6o07HV3NwVnPXwyEMBmzNF04+4BuH3NuwaD
q6n9ZdqnhjCAlBBniUgu2gz+5ZGh1tlKfXL5z5llzoQCe/1eMJzUoIQIiFjS
hI//Ysa5+L2g1rJNFpsZXGa7ge/VQpXLejHnl7tjGqHTKDsxAwm5YO8sU6U9
LOVeWzkX7tU30UkN78Re9XwxOGhopbyPJ2xjI/1QltQ/B3+FcptwEEcVeWC0
nciaKfIsWxOj29fpz3pa5/ubI+Wsb9+1fELMprww+Ggbf7+3XXrHgHTDrJvV
T3C3EiiD5zJv4fTOvJQODG38NKL5MqnopZsnYDh9U4pfEZUt7U0ifEzhWNK1
0ciUxmMRoNQ0iy3wV3VQM3ubV/IefYKhSTTbmup3spxjHb/Xxt4llnxIMITA
OZVrqT1H5gxXVZVySfxnGdDFDFWnryLvxgI6ePwjFIG7o5mJD3DTC6IOVL+v
tYl8FvunKbRZenHe/PNusjSPBD0YlU6gbfozABNnjYYBigItBU5jkXBFhynf
OvoGi1/rbGh0hxiOFhhbd4uQqGvobM6UrXcD71X5qCLRe1MkBVnnx3a7um+6
3W7PeEuHDNhFV6prHmM+IftwQKYyjjr44EdF0sYVq+e1M+wMKINkBXEtO9/Y
/bMqnZXg+aZ+Hx9vwmxo9AXxp91QNYamAxBUBVa3peE/XBlKhrWyO9fugckU
jZoqQ/Q2T9D/vgkaa2nCswXwMt00eQUhPKXhCv28z3fXLIwVKkkoD9mPCTUj
A6rjbP9JqpG4QgnjWfAQHl8J3U57vW9HT5PO2zWTQhHQWNZBLXf6uzA9+c9w
wNnBu8K1FrKiTC8LV6sk171aUcLCffpwdIJ7YyFxe8pHKWoUWFs1Q8NqlZsD
kusfN8nm896JQzgcyZvpUirtBuL1KasDl1TzlIfx5QMiunENeQLPFnUkF6vk
1OmcaPyW228zw5UXt1ZQHADage7cxFuAg1O8nr1z3PB7xp+f2gY344e+zZ1I
XS8Dgj1oj4uyJ4kdW03y1BfJBvAjQ1ovajNP5fXhBozC3/fDG0dF45KCH9o+
c8TtcEUXkxADVPoPcz5JINiRwOdOva5gXS12I86g6n9vkXp80l6J6NAD3AJM
s1Pd5faoSZidRA6w3FvlSsN0USUu7666ptzSuXbKqiDh4wcFwI7xyDJa7dq+
04PVL9Wv/bZIIECmYdX/wkZaECYSWssKvGmvcMfGTE8YfnF5tOGZNWfdKsJh
xum1P2NIk8DCAIl42sTleI68mSyVWfw0GjJPxJ+ATTP4lUh+B2780Qu+0Pw4
G8ldqprJInpJw+4pWXCjfZ4kRKvKOWtHhsV9+lQ5nYH8vYgXeyz5bT9e6sHo
rBfv2iGdIc7IJ0Bfujb1Qan6Y46jRdkl3aaLmMWaqmugd1kcrvA8eV0DM+Xf
50fjSL540on8vImb2aFIV7n2doffqegmmIevLO3Vg2EhUfHKYWq7oDQcXjwU
pAN9KfKIorUKPoxFx1jZzUOzFuVEjr5+9COu4F8dpKiuZF5MO0SbdHGEd20I
Mml8fRfR/frHTc/C/P2M73LEFrEjDv5DhjJZk0/YeYPRsVlBdMrPzzxGg2m7
roVYdo0nADO3uT7LGuprXM0MwoyJOe/zlRJkvlu+nWPCACsqD6+G5hd558jk
C1QUPP1vRdXM5QljkOFkKLWulRh6SVyTbrh0gdcUi3JlMpGVrdnfLhczwt1/
BboDMzWPr5eWhKdX95IPeauptJijbg7R6XT7b1hcs1VzBG1XLaBr5OSAqYfb
a0zu76/mafbQhiSVpbCAnVrwOlid24pV2j/U1QHjs50NC1RCwQITCV4A+mCV
XZGO3nZUQbfFdbHjDGp//AhtLnNDRbL86iAh7FAmFAGXookJy1YFiBNK+vsO
VtlE5PfInaSZU/SqMuFQ7j8aQw+jJw/2NrCT2T6aDvEOcRyW1lZLqSHCJAF6
1JBsFsuQITd2LNhfTfIPEHBoh3vDt0zRRw89FHezcAPXaM8YjvhUdqGmIH17
oWX9ha86lNGk/tP2k4W6nBvmvV9PGFYYxi2oYrlrOX3NBkOsKkUwPq+c41AW
xCn+VJyZJeBIfDOduSP2NuFWQ2kH2H+mfNJ4hu4OvS/Fyq1z5r/qik/Rd5d3
mA/UY8I98RZ72uR4Umue8VD77d2sp1TlbE5vvO6LHtV5SnEpPnGEMku6Vgms
wlcONmSPhwT0Swx1MTNbdX42a31YyB8X0Ivvm6s11Kaj6j41ct4br+6DpUza
E9Da3MZm+uWAs9wnZmmS0soNshjmYxBgAeMjbU+ZNAWPaICzkBXp7PB+Z0QO
ZKnI5o3D+dQgOBpor0gO9OOHbTCEcuHp4OvHCd5yKV5tNgbHaBdu22p66dmQ
ru6OsELOsHFVVtxQcAyIRzGk0PVCKWfuNqs1ECfulmM5tU5a9yp5Es50rKov
ycXubA0Dm0YwoZrkg05IqLMGy4A+UHxaawQot6yDeGAHpTdUf8wWHE4jA3mZ
B8cWgEUSNAgrU9bYLdNZfLt+lUNTH/xWTbmdEJuOULP+Sqffcmap12Sg3XHo
1E4B25WyNL9Kf1p4tP6mMCAIwyhKDTOg5xRy+PG6a9h6Z+6BuQ+eMfbshld5
bcDXSgi7bliFunJBtNIuGo/JflqfOaCapRpXTlBJrQdZ5ean3peZyHYJpL2I
KGBdtK9LR5vu0UbWwnZMg3YdlLiw3HbTSwDYiGrSi2OuSHIUjQoOp8F98T/q
CbflRIlflz3IUX/7LMu04zJZxzLBNL+Q5aV78aEC/nYREt3KPbMdh4nMfCfT
hq18uWGo5SzRiBHW88KhcP45c8SCl9q4i1cPcud0dQCqGXlle6BgL1ZZCzIL
rlyQNkWBDf/PMANCmQEpP0n1uund7vyMgp9lQxtCSPj+rOgAfsEhIY0TPh8g
4MFfU/b3QYMIseItYU0iGw20zCZn2L2zJtE+dOKtj6vem+ajs0ntNo7G9eDa
ywmIKsMV6FSVaMuSjqGg29OIIRvXLukQFRHLoqVJCTeKV3xEv71xiyc7qxyL
1sVdqqQb4mJ2p+14HCpxsUuzg+zlTpVOZhBWaKZjuUVhYXn6bi0DLJ5D8LMx
KqQ1SrfoVQCFeP0iQ9ShIJsHlLtWpQUxiWy1XeeJrRUmdF1Ns+mZsSlK7fkw
x7Jm7FxAxtJiOJ3cofr4O6yMiAU99iBgkD3GkW+dshcoWkNg3jD3NnSkP4TO
lFc2lugAkJQrUof08XawRmi543yCMnWEfCou+IsVe9ANg0J7PSJoiKk+ezuz
G7I0eRf59fkFQmJnrzZ4vA2k2cdek0mQdkpl1KKkvGeaN82EeHDQZPz1/Rio
KqlXpcbYdSanjJdaZSGml1Z9i4hwfjxzOFMkidSroaCnJo7sitf9zCf0Y7om
cYd73vhnQhlGwPkbY0rGJHhQSmnhuchUou7vyoTXV7sakobQ806fbJNbQ/vl
y9KLrOrKdoZavZEEuagExXd2KunkVOiIJ+nL9QyUkJsY7hdoK83tGNj+Zx15
wCgZIMPUeEFL0KKe+FPShvuZW3QfmNBuhals+F0fNDBUxGFkJl+HqKsgyNXz
alGM2/PfaKny8LNZQwzQvCKlR1dSxaTv767Npsgnlu6S+DKhG1uPoq8mknFq
KwqAduUuHmRzj2oxujQInkqOhnR4ZCLGa2ozjYCBG4FRcZYaFuz5Gnc3wcCX
ezYgqojoVKF8HwjENrKnXTJe3yLO9bMEhb365XntwFF+wQQFYb9bXn8oMcJv
9M1+/Tpkl1b1vNItcSHDhqBP663Os/ODMiBEwA5WjP5oHDGsTSWcDKcOobsu
tGkCg9amM1q5UnpZ8cu1miiicj8PqfRlpN2lJu/QiQQExGt4XmGp3cZx3uYD
/Q6zKmPgG546XXsFrhSRYb9b7YG1ibg0carSavIdn3xCIF8B4yre//Vydli3
RzALa2o+ly5G2chlULJddJG/xDuLzUJfbtgb1mQm6W+zd1pz8yEkTcg1+VMK
jilH93QMCtMFDAZWThCFp4t1WCQKSSP55Hb4ReJ94HNo4t2oLfrufDlsYlV/
LmACrDeT4oPW0iQC3cw81KWRdYKX51gK2uaqr1vdWbIGOY2rlGOjnDMHfxCZ
iVKhEdKuQW8/fRkKJJu79QBrc27unJesKhwMlR8oxi0fsUcnrTHQYwiiR1TM
85NiROodrT42E/fF/w9uUMZ4GwAfG0z2kD3suv7uvOIHuz7jAWNKgzRJWLq7
n4pcKwaVeVvl8rqTC6wT6mqJ/NLcLy61I6r8uDUEH6lRM1EbiJjtU+TlkBi1
q5vzVNyRwVhFuDFOU2NsLX2YEajEY8HXp4hb2QL88bxSSf5dir7qxmdjY8Ro
beHfjLJKsh3jpZXjiotBzlzc2D9vQ44ahLfwsLRZDsNjOG8KgswO/0N3wOda
5Q0QM8ERkLjoNnkSSqP1rh87yJ87L2B7PZeeie1DRXgJbDjH7ukQmnCeyMCW
YcHM8DUlG46zDH+XibUzVOFkSBF8qOHZOVkYI1GGmArzGry1dAi7Qbd3Iaid
OjmhyrDHe81MLF/ZXoxULiW2JftJn144h6KYRplmrGTidQNhVQAUxep/iznR
WXtVfH9UZm6z1/TnjcCKqEkW3nylcMPjJhsIKZVpaVFyY6XQriXvI8K9qIcV
N48hj53EtFUBwMT7M7fOhy0KjUpLTVFEsnT9giOsq45tnygQy7woepW3u0Pl
PcTbMgG4Gr5C6Z0riXF6ipFHnzNxqfFyHUWMO9Tg0GDoELjcSW9eERzA9YOV
fHcEqcNYUD1FwWIrULWVIxoONYq6H1TcHtchL3j59NpbcIrSK47L1N58WUhE
VZEtFxFto565aOn+kwqDLRAV6LqArt5owqyRC5gRgSPG1a/TCo4E22u9+aP3
vRrFUeu9imPUELg5FCyJi30DEG1YOyFLMAVgbZsJ8DSmNRGkXwgztJmTFCQY
CD6c26OkF1l9tqOL2ruzL7liRYY4PFpJg+PvPGXRVUKx7gOnGdttgqNOFvGq
xL08QTvMdGanuwz10vNfexVZjurVMdc8jFyqaZ9LBVSbyMMKwcxcQOjLcJ2T
jFgNWBCdZczSh+EMPPBx5HDhWby7k7La0p2gUJHjXHYurirZpxPxTImIbDWM
hBOyU5xemzsc/Uoq4KGEt2OmsuWMqgqAu8ow1FMM5jR4DUIaZ4tZdivehGMZ
/oI6K6qq/3a0TVGodN2XfI6IU4aepzjG4SiGl5pf18gIVYb/stUVk0fd1XL9
RA3QuNltwd5Jf2YqAjMQlM/DO0xRVtmM8i3Y7mgEYPXfxsDI8JXns+TRMVGQ
H/jjgUD+2rNvsQXKXvhGeQuemOd9NzeAfZm8Ru6iGp/ppK2ZB5jvvKDrj/kH
wXNoxbpESRTN59tyBnuQNUUI8uSNAr1X+JqH1Zq6U5AaSc0YPF5s+c7wHAmc
TpnLRThrz7EY030nsWF6bZtDOQ/gW7doItd2lETpgPLSBP03s+WadPPf6YPG
m3/LKNjp0yWt77nnuwQUdE0aI4wFunuUU9rA3Ao9HLRXFcjVJ26T223rARyj
ObCw9Cyy5h0RPzEWOxbJRYXeJBRAsevo7c3PLK8V1qUpRslxDEe5A/1Mr2Ex
1aYPgIsaLTazNFDYo+XEOZNkbfaByj2OnMPVpl7OFSNJuoClaAKyg9V+7yyI
bIKXG2gbFyGg1p+0ngvzwYXyJndnVme5h71RX77m9vMri1geNoZsjtaR2glw
P3FqF3lKZEvHpKfc3A8WU/bI5K1lJPcj0zS5QQkwWGxpDz5+UCH/XiJeIMQ7
HhiPKnpoKRaV69G3Y7xn3ShJiOTMu6UlsjqWIc/lJO77X7o4gLB95YVTFIS+
F4mDHjQTp+aiqgrkrffdSMiOaEiJKKjztT51N7g+OxMLZVgwRJvU1YzMY1OE
P2EQkG09WX41We2rK53LOZT7ZxMxlHTLFYeZoj7+EoPyjED/ohm/eOSd60bl
gilCPFmgPXlIxOfc8WsXcjra57H/RryoQF+B890tsV8q09W5rXRNuR5j0vIY
rV4/wKGlRANj/sOofi+R6AWxHoR8T4phJ7zXGaKTehBYr/0jH/vSCcvMF1Gs
aCi5DlmnHyxZmzXPp/LxXKmTtI4dCmk7eEgjRpxX/nZ2bxpJCuq/TOPXDmeJ
gdWQL5n0A+zydp300rdY9Urn/7peHUrwxi7Nm52++EGhi200I0R5DXvAQphs
KE4uqdI+uLEL6t8UNE681pVPvD8GR/HoEirogrvMqmu0zIr+nsGE+MTencWf
cbefW8YYvpGSEE7L8tTrjpqsMZPT0X4EExSWq4GCroGHyroH6k6lAVtEmOdl
CM4T5YSKOY3QdCS1ZKQQRi6V4OCav6A7IJ8nyWOBjtdaWxhplsLAsFhEiGyq
1M8Jipp8soF6+ZuigQENieyxHkcCxrYiKTtbUupEDN+QK2ditSDSIdP09puJ
/KrhARO5N4rqNuUZH3CuE2EaDEBNzY3b3Yd7fnk9SnYQsnwVvVY9unnT2O6s
iS7BKY0anhg2nliunJIqzrqhuG6kyCqsG2Ailx2K7+CR5hl+95ZpD0Q6/IAu
JhpLXggJvKGv8awzA+/IrXYDAONMYn+sEWWy97Q8fWMplRbEZRj7fa6yhV+C
HjJWPBKW1V02wQyfuqY7CKiJBZeLtBtQGnpbkC1ARLuvXycyoqR2oTCNlvxf
qLjZu88zUCTlBF1n+CVwfErzyDdvvnTCDL6yDj9pgmGMy/wSfoofwWxIuIlt
25bqI6bIvdAZZKPIN6mo70UeZ5n4T0Woa3SoZ4QSVEKenB3Fxfk241JYDDTy
6+UUQNcqJ0hNhFGZKauNLDRS/9TXmic68pULbwl9hdenJJrseUXIoADPiU4Q
ybJFj/tFRYWoTg8aIeUQWalqVlQiVvq2uf12R56DDBND/LFZZ22q6oGImd+g
XE1DKPnURn429jj1WMqNwjP1lGGGuxv1WgjDBcXM3dXWFK5q1KKdWVOo9D46
DeL2BFklfwbF/YUKE3+qUyRDePDLdy0PbrGVP+QLAsZOuEM9vyKvzowBtOkx
FZDaoCOCnT4nUYOPpS18UFN/WZWx2jdyIJO3kIiIoQ+C11O/j74ts309e9q2
ZhNTAC1L+bnZh5qlYB6IIVYF/IOkwnla/U+D8xfKwNAZKAFsxvDl0h9mHmRe
PXQrDQVhhifGy3/ui8/pcXBLtf86SIMXzMphc853pPPbb3rGHGLxMfmbNSSx
pqmypUiczkCJrz7tA5Z2CZfEwMtA6gUJrXMx3CNL0veVSb/ydErL94Ayp9En
ctE8fKbfozIkuSY5ZivdCp1S3ry1zelL37tAymV4nbnRjtNResn6THzKRY78
9mNX1fyNMnzHEalPkLUYHWX1Ma5Gb6M5lHbkoPJ+sLmklNr1vNK0EsIrABOu
3+MgNFC7BAQcOxYmN+4/pouLVj64w9xR4d3t1QtDEel/Ttk3JyndUJWlKmoC
2gXbTqCk2ZE4vp+hnPNj6i288tFb+fSqAN73Th1DwaKWgqE8k7lGkRKXs9pa
eqhQI4k1CepMBoLWYY6x2dwzGaaKCSYWMtOdtX7klG4zr/TViLG5Fv94XjL4
/0NOVFFKj4wFbJTaJTTo/d4pEhY3n7b4bOrwnw9JRba937HiJYDCQC/oyzIH
GPcjjQA9DDVs6InGs9t6SX6GJ+OmIBaVl3qd1BBsvan/ey32DpcQBBaWm8Mf
Ep7OKUUfSq2/hAg3jaGDAkgPryHCJkU7DIirCQPSbnaI5W76PQaQpng8hfhq
dgCKEwvxeweCO7iHtM3M2i9R1qG8x8906saFByC8VQrs3cm7ui6TKY7MvSGU
6S8q+8ON8QWYJRaFOEgHfUOPuMbtfqWkkF1IzbfqGfhldL7xMkbMPLkH1sb7
2+NkUt5Kumu4d6oG/EKNrSnw7QCMpO3O5735GBA2vpBo8m7ZnnIm2RQys/sc
b1XNmIpqJQEU87Q/hNR3ima/Wzpkaqidpp1QAAJOghXcD2WKYSNY5sRDDBU8
kU9Z8uIgZ8m8kCZjea/gWtnqBchczVVR96AB9SzAGiE0bT90NxylbKaa1QY/
jBUb7Bi6aepQnuMV51e1tZwvvxdzZWYGZypg1mzvhNUdKihFNO2ZrWMEUgf/
mw/XAWD8eELlTt4HM2jr3kYX/TS2aStE/DCkEznJh4cmfB0+Et3Qgu1BkkRk
0h3eVaVtG6dL9P8OlwcSFy4b5Z8YEAdoflrf0SYwDQnfenrpfDsYHBHwmdwO
ley0hWvO2/FbA9b3sLXxHJK1WR0n4YRLno2Cfu7ZPlYLvDvaUONyLgjZVaCb
ptjjvScDR6fWhMQcKyx9r9qBWD3orJCBOiXBkBh3VPGgSl3jgAGuqtnEZxDd
UnYvG4sZlmzo2DQpgkjONPeZKDMySsXD3VJ2WbZ5b+6FfejlUGMOTT2KLJLa
J+3+/pBBba1ZItknYAXiJeIOF3J+XO925OoKxtWblT/SVunN0IpggXfJPTPi
L+yVuK1/Pij2VQ7hxvdGCsZ31IxSZ4Q59oNDDP41sXrckM8UY79/nU6HYMJa
fYWie+CeM64bfswqwQtBdqGUMXqZeJQJHojzsmJcTTZCm8j9u1ZkSB37lQM9
EeMfxl5baNS8kSyrkYgnLJoftqZjwqP2OBi2qZBDGrtEEHsPubnFhCm1QZ3w
KqHVIWLnJyOcZE3aybxMrMk0rdj5u6myMQnSbwFC7WAsJP1pOECiRjmgvXQj
vzxFAjkMhhhoQB0WhfyMoHWTfr9Go3VPCQDwvYFEZC+xkvG6SBmNqLajLARm
OVexPNBwUPRB4KS1263gWW+VAYBL/Y73qHK021EO3SkgNbJHB+YoggLWnllO
EVp9P/U14wuuEXjTudk7hdn9hWO+AqYzp5MAyPQU0RzP/87+0EacM79+fzs1
2FSemO93G3zTj6lmHT9eqINhwUauTkB00YQ1ekoms9GK/SyCEGkmgvqRLFfL
MUqRWlfsxK8RmOyGiiIRq/6eINnFeqP6mzkmsDKe6CrrYe194Lqr8hT63+Ig
2kJHzkJeY2maZx6gpkCxx1PtYidRC6/HZITSoQlR+lRPvRTynKr884Uo1/XQ
adbuOBJCZx850o0REb4hye9uEQoBpWE3AU8tY35nyBReoXysp9gMMgExPdWX
iIRhbL9p26+ewcX36ogL8m6hxrCv7eLnazi4UYKO2i2WOZ0l/me9O1JAOVlT
WSBSfT4OgQlJXWwozL3hhHhh4hf8JAwSC0jd8JRBbak9uypK4bMMmLT3CFEC
NWN7JVog1h0tMzHciplg+pQCzZoInjrhu9+lZ88GqvXUA9H39RgVTYXKsyBd
QVpzAyTIaZEpmqxuY5c3NNnHSct05Pi31MrZHGk4Qd9fAR2rpZPnhTJb9uTX
an+7Mytmia8xIPXEp3oh5X6G/E9WHCUHtuCvJ/OPkcpHBFSOydMmZs5KiZPW
fL3wFNOHYFNB/jd3i5srQDPZBpwiAoskVmzSPLhJaBzKicmQu2v5ZCG3WtPj
rCBfSUs+mJef5+2D/PZWMhmmQPTMh/xZE9D/MSxFJzsYrCsrAnNs3/CV9YFu
V4Pde40YPrpKvkELPa0AiFD434RXAN2oCRGCrn1fxl5krtbqoNgF38c4byjR
W9PE19xxuoFKczNDPP/WghBmNWundumC6BFJeq/hCsCRIweQaakzn7rklaDI
BhLlDW2spI7MZX0rn9kgo/FKOG0/OFGJCOK/jnQpDqRxiAySHiL4FVWtv5Ri
l63Sw2GsxVlfGVtdX/u8cxnD5eXM/pCmVTAdSv1bGpS+n6siH09nd9nXBh4a
+0gniPzY0X38yKIXEaDQjISq0IaOUCZ49mDr3XU+Hljf3bPKBOeyBydOyZ5s
k0qFsd+pCnCq8Z7x3rvxKqP3YUt+8IvTomR1YAiHrVzNQGGffb1KnqSqEvvj
94ryds8b1vmBVTZ+E0usLSNYSC+BewfvT1oUfkGoZcbiR59twATVErM/HhNG
CIYjolO5elgym4XqwX84P0sS6mIPXmfeA4E96SKlbHlxVgwmMonAG99LP75Y
lnVDHq6beCPs8Zyc4x+AyskiOyyA7wAgnuBFcPDMGxZ0JrxPid2C31iss9P1
jWv4Hg3j1Syr7CaZPk7d8ppVybWSc3/d5I2TIa5gJk5KefaEoScOZSKNb9C3
fn1bfu/hMDMax5CIgMazqQCq4I/wFW08UBhkV7cWE1BIehLhBXyf1bS0HRnd
0E1cyMhap3ifofqtRMLrFpB0OEoyV9NLsiqEijQzLBHvtRT5IPoQlcTvZTF4
iTYszLBsJZZPYGU1o2sarhh4FG6GzBxYcJyDlT8Cg7UvMVnITr+R8yr1tUsk
qIi276Pv+2w/7y9DM4ZK6nYWb8ZY83aBtPiPy6sUTwWmJ9m0OCsmV3ct5XNe
6yVb/G58RA3yPMZ1u1oBKwmAp5hFR/nue0PY47t3LVkt8+5LqNZ3Z90yyXfT
cSbWz21FiwvRjcr8EBVRKK9eBZUb+tEH2PQE54Lh8SXLY+K6RnOHX5DFjjMP
1leBi0cUElyDfKFWOzVvZOy5BwBygRD73KQ1VrG0Tuy97SiDAPnFqUEb0Srt
N7fUhH/ah9BwzKKvSrCppq5m0Fw84bMe4pQhCo+BBOZ94OBJi4Q81C+dCNup
PLZcTYTOHVrsL8RE2Wucvap+WMeYRLG7bB38zzt3/rSyMVuBC06i93ww/WFg
FzzrponlCI53qwPTFXvc6P6FQ8dz6KBL8cCrcxwAlNtB2DwXjFNQPaLqLmH9
u76cgE6wNIcWQzojmNcyPlQCUSWrTQevmv/zlOSPG2jXbx/gsqQ5ihBdaVJv
tXFv6KZPVew13iUOax8dqR/jWaCPIoopwDA+ff4iE6VrXUsqn/dqzoZif/Pv
xwvcjw8e+08eItIZmJ1qPOH5SbbIkoQ/9qWBcicajCCghQ1Nl6cLjX4jXuE4
/XBynf8KUqElRvLSW51+UlEg6J0kx4B6NKtBh52D8YtMzNkH5uuEKVgGy2mN
voCE5nn1e/F+RuGQWjDBw6fkZ8gbDQmcZsHNAyG9+4i2i2Ky5nGsPX18daLH
RGFp+oQbrWjaUb2+7U81wOcyaxRfDYyK6UoJiRpeprYDPuHWAdWL3yz22lyS
ynjLvX0gNZYZi5nhmRTuGg48PydJOHbw1WTiveNpl7NPDJk/xuuYV45nal9V
CNPKwD4KPz0Sh5WINdSdwMcydN6iFqBLp0RQaN+j8CJxnS5AO3WpIRVDCtT1
17FUhAJ2vTRLv41W4qwnR2FxNHeDnn0DWfhA5fZZLxV72pTtkDLjDPP47BYQ
zOygsfX2lipq+5a4CwaRPkKFWF+BwWy6SOfry5dbWptcZeXSMKQAFRe/yZAR
pjZeoyATE1P4iuTI32i5EI6tLEdUS9mktNZkSMD7nMu+7g/E55q1ngrBjbae
N0HJPFECxTcJC2IiTe4acm3VHG5L0QlCt+dk2TjbZBbtS2RSlzJh3viURjaQ
+S3y4PqHyNszL8oBHZ6aojvBDBcWXm8wZJggnXqoEKIzKs8579IYs3nfhnZg
KZ9lgoy7gRVx+BYWhbEKKi+4qG/KEdnM+FGxA93CMPYVJPAoyP5RGsjK5lmc
l8llX5AfG3E8EBKaK8DYACxc+uQ9GncX7fJ1y1gsxnUy9pKYDmwJQw3jPt/V
aDJTKLzavW3Ufo5ObTRB3aPyFPcaypqW6+TJHthwiNhahr+nz0yDLmQ7K6zq
q8KN6xhszKMVy3dx0dSYvVqBie02/bY+hs89FLj2mZTBb1A62XBoiUHITzBw
zYsIfQtqG84jcV1wuQqy5VUqOwqSHUy5MWrxfc/pXbHEmAxsU0uc+8vSZooI
3jT4zNlcQ51KG4sf5DQxpA6VGD2OLJHdtCN3ZQQHRTrWdYwiXSNNMb2yevnw
MAzPzZaE2KcpWcukAmvl1aY1tVP7Vpk40qKB7z/Y2I7M1Carpic4c+xHotEF
Z/F//IvA3flKxsqqEi4BRaO6Z12jRCGYRSmQAMqQhIvgM9tj8kSVu9SZcuwd
tuxC17zdopuXNm9lM2H+pkQiZYEruXwC/B/JktLZRsgMmrHxS178EVgdxkPr
HZPF8vTaUXeEw82TjI9SUVaqFoMHZbe2QLCWK8m9spaAs/Iierg1htlk1wo5
xKma/Y7ZNrYMg/eL36uj85jw3UwD2gbE2NUOKvN8texi6k0ow6mdWu4vfrbT
6yb3yaTrOAq8aXvscUW/81sD8gTcRc23jrnBAgazyhzYEr/cOgM1d4wr+1rL
cW4Pj00ohdigz4wZapal7XsaEQoDtPrVeCzLttKOiF1gZnhHo0hhKFIxhxHq
vmcB06kuG4dOdIFGGnFZe+zQYMhkP8/7MZX+65+uGOah4WKPWhgCWxmFQxgc
ML1uSrs436EeS2denA1Uh1v17S9St+X/gxoiKcJBNt2Bad+1CQAqdIHYDYPb
mWw10WCBIyLnnDIbvyEd/4VW0sD8DISowAlkiQHO9TLSfjkKU5u5ugVvg/Gc
qH/9qo6PXlGH5ohnQY3nrsuQwLhsIgF77LkLxlvKg7QJ9dZUuh2Ib4DfiMsH
8vYG0eLv3Cf63oMmjavGV+ToZMFAtyItMtjKOISS9aEmsuvFTftNBl05YUdv
Sa/EiFDT16RB+hXlhkkdnizeBrwOx+o4+IMGrHj5rmh85c0IZJQ0IOfwUvyn
ztDzUiqiy7HihXohaxNcKG6DtZK5p548ZEkKr8HXf8rjjMAzDWfhPYhJQuRP
LHKoTujKRatHG3rbSEp5iuNUi4Yk8S91r52K6KyjrFGuCRujDp4YeRl1xZDN
BXadKFrS0POrE4wKbGHnvC7p6Viekxes8qu7iaoJvIHdpQR8CrJBP6RmWT/j
xWRqTKZK2HRwTIp+3DqyWlVNaPRutLKzHl8Bo30qI2c1ZuEzXM9Zc+/TP8zl
hPwkS+QO9Cqvx883hzjIdehurDwmTegKMmmsDbxh1ppOYQ8Pyy0wspbQ2ASZ
6cxLVQzqNK/L4nDs+iJMl0NmwYG63B7/RoF8jH4XBXO49ovJNEWiXX4MRBms
JCb9dE3QcaOVMeXd7H4JA5JSjhQlakhBalE8afn6u5aIbe1e+tbSM3+WuQjY
oKxjpSPAB/RpxJKr1xLLokCKEKWc4hdDBFDi+aojJwKy+N+Gzn3juxvPa3Cz
kwQiVfMA9xOS066ACRuunx1BQ6fxBeUMS79in5IKuDY3TYvT/Ftv85eBciKH
G8Y2OTQjTA+HJQtegaYJykbBLiCDjGJkYlxSMWgjs4Jqoaa4AnFek8qLbDOK
yZPDFXXB4IO7AG1tB6Epqw2dX7KuPLtnlv6B8+u2Vfi4Xa60l3o0n5stB2z2
HcA8AvaoSZ/AgKuYNskvsN0Wf/jGEes5DsF/mTPCrywljxjjdrULTHID73ZZ
3ox3cWjK3wZ8DtVI44nOzntxG1Wz8cS01H7zhaTyhCKPLPNoknRa+1q657un
lCHwK14FJC7dJqdirqqAHWQXG3SQOw+Y4bnmsfx/wSsxj9KprjfvRApidoHH
tnA/z9Z2Ox4KFYke0KsyWFzbLG0Bjmxmznh3CJox5LdnqJL6RMaAxVVjdpNq
fk4aNzVWIWkyGefZFqfCpdJSwCLnxiW5rwzx4E7IktpDPSTAcvsmvOodDaV7
p4UBqwMlnxBvw9BfD6JlP9qgEFE8x/9R0obGU1MBIeeZ8T4WMf6NYpx1R6SZ
t5TpqJfCFo+jY1aE0SfKt1+b2R8pC5vckT2vyDQnL/JKy6chLfw9PMI7CZlN
NXmUTbI7XqzMKIIXi8BrglWUWtJ1CqNCFE9sQEHvx6u5t0iyUIGrukPrOSKk
Y2slXqu8R9MkVFMg/Cj3RnjodUL7zPWmO7zuo4AnnIO6d1e0v6dtYzIa41sd
bc36/fnf+sd+P5xFlSCKS1LQC9wjHfjANwtVDQBmqpIUTzuSm6PNi6NHWifE
JNfo1/e4fj5WNXzvDJuCt+yTsOkS/77ldzkCXNkY78lZ77OXN7K8ocJo7grj
3HymI8T5Q5vVDgj0AdbDd19filQiXR4jnwlpA8r9DFFx8uqC4zb6nfgFRCFa
l3tCJs5ELkS5slc93fPSJuCsNYLqwCpCvQh/uBuVn7unIzAcSdnX3xTplMEs
2BbCnihawFxWFthGf+4HnzKP1LNe6AjYorMALwGaJZJC6NNCEmml6S+hE7i6
M+tyYUeNnj0H0Yy5DqNFOFfVXSGZH8KscrD2Qjs3bYOYLEqHXtCzOu+IXYwv
Kp8ibNR87AVC9WlI7+im1vjzYikL6/DN1DSITIoWKqTZKHoGW/pspRHy+f8w
MToMWSsTNce5F/vjVtYBv4A+EaO8hUqdMwQnMep9vTdXVRpWiFKhVjlH8Y2P
JCbUBW/XyYLS8p4oLhWxbPQXwIUj9lvZfM2AEvP6ksdZoc5bKO5sWl1cHCrA
P9iKf5Y67wQAPsS8YVDzlUpFgGlpfe0jz2Ebeyr5yuzCTLEkEEYANE3RWXvf
KJuho9zqSQjKTrPFkhpmbdrVZYj7RNcyMCl2IirXyGWOVrn7wMB01RXAPb52
SJhC6xtfqN3yFV9M/4Djy2HCFaOFnr204nKyxYqP5A1534dPRXvRGausD4qi
TMi/dI55DUZuWGgk1YCSvLRx+jCsbGxcSGGen+zFFtykw1t/iwKUtMpew1Gq
uRekhGiDq7RTCLkx+d9w1TSm2JJiJGqRvvb2YGyqKBxCCoT7VnAMUifYc2xY
G18l67eZvTDLptPsG8LAqjFszRsERp39WIcsa1ZqLiojdOZV95DQJLsxvyPL
tZ2rp+4tW7P9SO/eaKG2QEWb4LW4D3sQuTz7RiImUnS6K2EjAP/FjKiQluVz
hzfI0bGfCnblQmaqf0q+KL9gSEJ8DHRBW1voVDKc+IbkvtMk4EBVmEEiSpqM
9qb9jn3uhgmIjwsxexZ4kI26dS1LbtuRFuyIWFJwtuYU1SF+bPWmooB5arMa
iv0J0NAfg5J3QR2rK+m/iE3w3GlIcTwWV19DNsgVruf/PdPFBsSutDO2wjoN
lO6FSVrEHCgJCj8zZa3yu2Ic+DmygBKvqPcOPdBALdGbelG8/NT7FrzMa82I
PiN5xs8wcSd9CIWcbXOTQqI6QtvqM7GTyAumjQ1lH4CZ9ygVfMghGe2t2sv6
/ZgnWl9S9Mbt6hEq6ND1FFbS+PESML5EovC9F7f8z/U3GiF2O5qq0DEmJaOd
SEOVHxHpNj/wI1L3kBMgItWkQBayBbIpkvYmYvgsnJbE31TRR11rpl2+Oj3d
EvIPLdjPbPKD8s6VRsz4APtW+EG785PTntKQGQIvjJJBa3INzgRvoFoy3wVU
XWt1UyDMnGU0CrpD40arl+fVF7piUaoeVn31Qu6JyUn6P2H9PjyDm4DSK40L
rOdUMhJTSHdWtc81VlKNO1OFh5/QHaXDrMt1va3SEcSThne17r3jEx1v0Cft
DZCc6ZB9aEij+OdrTsW7WBaX3IzTNGxh1iFmWp06LdwfB8ntArou6kQtQZ6H
IBsAa8XWjOcE8y7TXo4xQpGO+Yk+TpBvPSvLfktbA+j4CSBTBkqCgbeWeBCn
aSAadKUPMi3PLD5ELy8/TfBhpLdRbgW/AftJ3xMNPk9V2FwbOidj3yQZi2gZ
U0I2rRKYegbDZ+KETFOmcIaJ1jroelOj0v8w9uvDifaWT7EC9r3eiVJpTJhc
wb2oEDPeFUIEgriSEsV6RpQTyZcqUr7R8loerTnT28F1tiosCArDP+Qoza7G
P/JoQg8O1TvSWSFD6UPeif1ckRD4q0oys0z8P+cUBdROgVm1ouMQQhHuanxy
1y+e1Enkl22xMyGN3BL0eKPwk+HqEXuOB1HP3mVYuO+hIIkEA9OqddC2NDWw
hND4EHmoSp/L2CqlrUPnpO4MuTjVLs//0JpN774l/8JTEQvm+2Oif6XotRq6
i19mhclT8SS3ONvdKEeF3siANiiFiRHOsI8MACaIUAaCKo1sPLHFBleqklDd
UcMoxqbuYAOXEo7g7Wb7NBEWFVn7eIhCoMOQfkkPtWcE4YuuX6iq85amYEVj
2eRGMSmEnEAjKM1O7qcTTvIYMGR+ShGN9DGub/8MiI9GnTrLzZBDvekxHCWo
NfVwpztDRQmAuocN4iEvw2BShxHW7tWa1BX+h5hCxaEjKPLqWYAKC5PPjTQ0
JbvwiE6oCss6CyI485FP7SNMobq0D5QjmvZNtlUYAdlCwlksD1k2ARytUEmJ
YnTgzzg6cbsODnziXSsdyZTaZPPJY4S7pUryxjZS/Luf8HDuYplIFxRTHR1q
onWXaaF3AEvZ4M0gFcphHm75n3uN4GM+5nevHoHppEnmEU/3EfMhaRdjM7SC
2GEKHyjcKV3WSISZnSRQPgnETrJl8m+LsY1wd89XQsSQqqDnRIKhq+1O6El8
2ezM2paAzLBT742lgqMTohtECwfAJd+E3Zz2al9lFtKqdOYOpZSqlyTfj+xx
OiiDuz/Tq6qO8LyYDdL5tgqwOrdmTZOzLyjcp0dhZOSWON24nUrJMj/8J6Y/
Jb3Kl085iLQejC19EPAkPf+vYpsKs5/w/3nbPXPEOPSIyczm4gk/5aE4P+Vk
vPMNk9jO3XhL3WJUVIW2W4/XuZcHPAubqEvQqDPozwiGtrblvR3cbSCJHlsj
ZC2Mm9lxbPh3kwS7gUohmmMMVMm+4g3ofAkRA19i62XwzB5r9QyNHiC3VBh1
AFrSnIEfZ6WEbDnXbOBSbFjNSTogU6HtKsvONUGThMrtHBBFopb6O6nAq07d
IjyzbWNrHbEbQw1HR3pCdSgnPdNs3ZnAVKPiElEUAgcPuIj1YjY0BsyYnf3X
3/oHQimBybOA5LzbG1uL9YbY4mcKbmalbqSKvgsy9yFVU4mzMil/CfyxDUqj
pdhSntW8nmferKSYmF4AY1xBRXMKZGH5hBZhOmRVNz/CsqNC4OSOgScjfRUt
2cBENcRFkHc/7IYv7WP/GRAMPyKXQhwW2diA9Z47C3noHZosTS7gD6rcV2+B
N3RvicDmJ8uONOzr5rh9hpHabVMe7H85wiv1s7OzgFfktAdngY5mSOliwvf5
SJ8Gqi0oQafuHz9cd4DbuZEWfADnbyAJdPYZrTmI4LQBnsaOOo1Rs3FSIfLT
OMonuaMSPiVXU3hNfc2YlcRfUiDuVh4gKgDNXiC7yxGrMXZRLUm74us7Kzu+
fpf1lxcvfPi87MGLNdQtKR2at0nlD6wE9h/G2wP0MNs24lo/Xg7bH0pqOzKQ
RL4oMu1vQKvbQrMZDAjQh0RR/iQvd9pk9Nx/xz+JlPunuBkowiTUkZ9lrKPb
j8A85T8yQJuQywGm0DsQ7PY9mLQ6DKKUD2xwBmFIsuZ6U/Cl5gvDRfuHth+o
TqpswjvrJyDg0bh4G9aWpMgZafc4V1HJeal0QO699/E41BBu+m9Ame1P1h8Y
ywZd+HP9dH5nCs6sFadu1tMYr7JbXY9lpDtlAb7wZ/hy3vajbdFzhK1qgNIM
/J06eT7V5WGqcLKq8ikjd72mU/uborzbN49T6RMF82M3wKhHgzNPEuf0bB3o
VS8NTtVraLby8H6Lq1tkgEcZUoGTMTTfsTbJPYoN7ti4eBxVMVaJXzBUqwqd
NpoQ/m3Fsbn1Z0Wp7ULuboPiyE5+u15nf+eUdZG86ij0EFwbie36GRe00S+w
8KtpxRPUVFkH1iBNcLMYPG6+5kUB/B3E7KyqZmlhY0AuckeKXLipXLG3c+jo
MWpy6jUwEeMX6NcJmjqnrDq2Dd0IrhTK2P4KpsM0/PWoYxjMFx9Z3aOGvXO4
TUgnoNEJnlFju5hfVtgUXEAmECCyVKb5iHHx9p8aqChzLGSoOPw1o6CTL6E7
kwhy39d3h8FAy8HNNNWqHa5KU8PXGnZ5w5uNnv4MTOO6vmhlntfwb5mI6tKe
2ieu5hsnCLPgS46r+4BtxfoiGLV8yzK+z6guMU/r1vOViTX/fpMB1QVcAgOL
pIP3u3xutHyIb4VXv+eXfi5yH3iwdW90E2vbha6aoneZLHBQ+YyTFP3hktzK
QvhBKfxYD+5n3eAgfE9rrvRuSDe/iCQ1ijMSYXxe+x/S6JGcAvYKjaewStfa
c97C1Yvj4pAXPLfqXcoEjQZJeAigUEAf+8n2e1Ul76LoeejnTTTpAoMz4jgT
epA7ED+mFGr7gaTxwld7rEwA+hwYczQqELXqTwF+cACqfwcgG1Wu3mNyAs+h
DZdLlBf7OCEQvhds98oiQsGZAqSKIxpwDyyHNYofaZCa6mz0Atf156N+dFpT
wcr88303akqGHD5F4+pzg5psMRi24A9jeGFxP/FWzRceNy68z/NQkIf6Z88O
5i9N/+qeg8vE4k1QHvk3honogfId2ypZb3uJ3hot+0LJMpwCkNABbonJi4vW
TSXuQ9RCahJIcsJ1iPBmUQfudoHiTVokTYaKJDBdYZ3Xl70bQmphgi99TsQG
5PSpjAB4tTKsWDNXS2Y0esrSTG+Y8ALH9+cH3MyazfV4SEJvA/9xDyZYo7UQ
1yuChkvYqnWj6kVt1r8C1jV2T6RPpdiWLXTouGZF84/FP5yHBA1LHA8fdIPA
LTVzBXiFm51IZaMf9xFRMKFCLrLP8IAq3IBZyy+E7I8IX0Mk88jiH/z9HLV0
hjRYw2ksWkltMg9eh/Efhah84bHuyGJcB7moRYUa77XDVu0T7WQBoZ1xmDYb
afyheEcrubaKQ1q4uIufeHfCT3jgjIAlKR473cFNXcWF9zE3UASLUc/E7TZa
fg7atx/IX6lUvnxEu3fTKpe81VnE4u+uYPy14wTaSAG2gGqhuLPrKo8Mph3v
IkZPFffmFOl5YRaM0c2ZKTJ604u6snThmIMpkblkMUkT0SAg71B2QPXFRYPV
0lqWKddvYkUQu9mRxvyNILSJx9ktEpxCA02EudVcYWRVUNM0YfAgq5ETAfHA
B3cMD4raaJAUaqSJH0BS35h5YiH26ezs3MTVWCuUWxDveRbdEtPDTtcwe9uo
6lEyzFFl3R5Ov5EE8UtrWcTN2rJ7JIfaRXclTaktW8Zdshs0pB28UhNxEu5F
/fMfMHI2K77OrNtrC2XbuUGh3eBHr5TyL1cwZJkQEcVSKfmjM6MhjBqgVPC2
WyxU/N5AuRqtaZjw1uWyJ8+K+Qq4p+Q2hKnJVvrEO30vWcIzzmqytVqzFsr/
Yn4WYVhpd1Wx+dMXTLvbYlo097XI3TRejyUCfg110164BcwTmbSCZm9Pdj+u
MxJjSn3z3AY16Kq1Je3dI+giZy7WZpCf0oYgRRod0VEv6CBWcPzwz3zZmZ8H
g3xdMfBb3O+fOHjTHrDE4esNI1f0/ma1twIIkdrCX6QmM5513OuKgo+ETitJ
iAxU4t9IFwzna+dxWwYqUVAkWB3WC6iVfmq9p8cX21V2zbFIUbcEvLnlraq3
ozUKEiPYhLjlXL+srRfSWIYOu+NZ5YcXX6c2WGhF+gK+y+IesxH12L1SvSk2
2uTBHQ5v3LrVGenVzp2mJD7cldHkTHqGK+ZCqgCxlo6528a4jl7grIegf/z6
KX8Q8IeFT2ZBVKDv/fCTX5I5diDL3gZqH6NydrRFNQrcgm987MTjRxlX3P4Z
/zt6T3UQj4suh8ouRXmOq3Z0FNUkdp0z+aplFb9XIgVpSrRIk508YU3sXPv9
tCzCKlQEIahWzTNU5IbSQg5hkjTZc/6wd2Z2YyrwxFc/Esm2P4bbHVsvxC71
yQ0xnubLGQcPSBMDZ5kQcW4MfKHnsBSApyf/s8xgzvnKmdpDd1lZsS7Oj234
rpZmt5SOfEUcEWbgN0QT3iiU/a40+DrNJvuK0IxzvEDcf3LPwlP1j55eaMdQ
8Uo0NfZDCL5Jir5fu44ZxBuCCV+0DZRzaOrZ5zI79Se0w2ZPlNuvhUxADxBb
C5Sh/jsaicJQmxf9G2MWPG/2XBs9A87nXfyi+oAqecan4v+wkq09oEUJHkxh
y5UpvBgz5dOxGgdlHXf0DY/z7BSEAOXOMfODQ0D/PeD/EWFw3qpK7emltujm
aJN1gQoIKmb3DU75Wep9IovWrgFT1pI5o41lwkEp5VPykVPRU7XwAbP+VFUm
7zOpsXLhnyd3WONg76McozdNEfUVAmWBB13R9KsPOnfw5biiT4rNqINVM4lW
0hbSzrhnsFWJmjJjr3iYXzVgV5TGcqWrxZVFUVh1CgFwTGiS/soMBmYlOKkz
/usGf7c8yT+EEzXurLivoQdVBssPeeyCt7NymAJYAvotiPedStbg8AytuKyU
LBcfB0q4QxCHDw4PEV6gvSbB6wRAXRh8fuSHCg0kS7Le5q+2ebpDz/csjiYh
U+3qkSzPDO0jcZ4BMFBOS15L1rFW4+Ad16j7eUT33Xr2fps6Lj3fNVQ7JtD4
AqwPbaSL/hm81eTsz60PLURLCvlNyC5Y36E7qwaNl86v35kPBLMGSx4P5NTJ
IoDuJf2ojzCrilkF8aVq3gooBQ0z4fysahjFuutQLDz6XoMEV/ObIpZpjg9h
0/XppPt+LG3TqyFRdzI/td2ezL+zGYUHR+LRAv0uZonydlB/28vr0xj4i7AE
plhOHOQl9AUZuApTWDE+tNcLjQH/RaFYbZAFAE9ig9oU3E85Kuj/QygC2otm
WFism9pAEnVQ0sS0D6GJqnt1RPqKN/M4Q+NqidbLCG2ghvNxJZXOGMmsqSka
ANIGhgeG9BrSNZAgb6brYLyvSwP0cIhZqzMWklSmeK7vsF1KmcPLCWl1cOls
4mHFi61d5RbUKn/Sk7sgFG9a6i5bM0g9dAGXsW0G8PwziZfBTZE3M7RDA8Ju
SNmbeBOgelXSzeqWT4UDEO01J/VivR0ZveBcOquR6lDITqFRfH0nbuV+a7ZV
cGBPR5ck9FZiEdOYA0LJfDr9n2JNjqCtWwLBWEfnFJ2YSu8XWvaiwRmRd2gN
mhGwkxv1v5FgjyoBFcrzP/t75MLzhlVTvPsCKxFs3mhZiz+F3RK7LDE51Hx5
avRLTBWZXfRAT9/UdqnYRccR+PyYTnkcef75y/HjWtVBDCqayGtHvTtkpoJs
FEPRgwlEmLa4JDMtFJm+CJgTJKLWvRA7rUsg8gyFhJwnor82fpfPMUOt7Bc7
vfsqYikDKTA5YqTDN7dSrLylDVg72TOZDFqfaAZCe7VL3S+dIMgEVUq1Z41D
Rof2Z1BJnV+NHlV9OJP3VSNDfVcTIzr6Urgk4TUKYbyQkAWKLyHI6VxNZ/+L
xLzUYgAcq4adeIt43ISIIG/re3xWsNLCL1M/wMUHv4ajPhPHWrKUhwmGsy4R
EJyegnAc8frOakdwvGaQ7jVO/Kc/zrd5ajAb0rjfuw+tRCLrlUPUCRuI2Gb/
rlu6GRQ43eEp+yuWLkEaBequJsKTB/XPhzeSfiaReCUmFwFypJW8kFkWvM0G
sP/KJP459Jh8W0phGtMKnPOPhmgDXKF4okM98GLW2bMVRRyb4xsNBBLm1cTd
q58ZK70GQpX2UDAtpsRHsNTjxDgSs+MOis/bXISr9cAWI3vSOcUcdXRJm/lV
S+OQLEmuAsylXkEpdo6UnOTQyPzEuC3wWwzDRgIpyOoekaN+gD7e6mMznE0D
ccDJ52+fh2qmRxUnqPBGsdrngZEuoLbBnJ9eJYAl3QLfF61QXOMEK4cAvXDi
zsqXXfE8GkhT0kXsFC/3kKlwcE0YVNbmnk/SMYL3uV4e0w09g2/9H6lT/eTn
082E1w7U/O1tjKpXqRWtbvGNbMR8yDQ3XOgPjcJnWgyO8qOQzQUQLWSYcDK7
+gsty4qo/QELIG5GCggwNnqFy+DmtWNoT5YOdimk8TsHqPetA6ewO68QJwZR
TXwvmJHzEoCcvkJSCbXBAEsB9cLSoJsnRj7Li24rM5OMvct6c5hEOWZKPHcp
LyqoTE8LciPHZzEcz+LZnKkYrdTqvoI5ZtWIUsjszndhd1wjOuNGQqTPw13u
kUQ9ikj1X39CQ5sWXQkZIwxsw3tRjv9ZM6C5wb1ERiAYgXCuSmyB2BjMs/xF
k5u9fhXsc34e7EIxJ/4ENVIOGPFdu1WH6KYdijTIxYkh9VKaJTGEZWWW7Uuu
kh0DSwJNNah8sewVb7F6S/Y2oA72ELHlif06xdpIAG8u9Rmqi72pInNOEcEO
EIZwp3pBdkbN8FC1v/Icc47ZWOGj75a+PGc5Y8S9YqLgI6jizDn1+uvyosb4
MoWmfWobgCyR2C8yR3ILIcz4ikrHi0lo4a1DF1kQNPiS8qT1KBODgAzjS9Wi
Qi1fNKg/1dv0u7M7/lm7N6HoMDyB1pGCltqNiimVHpKf92jokOV74uln5qyJ
oeg3lqPNz0co0J2GANdGWe6FCKnd3f497CW9iQqzOxLHH8yNQCOET8x3+C+j
Nx51LA8oQYchQ07noqU05MRieNLr4kzpglXgwQQ/I85Yt1MQB//WyCbfVO8I
fQme3mITxxlLAJGDMN7XBy2cZnfyO4aZP8a29qihtce7B16P5en4VEbZENxZ
kxJBRDwS63zSWnMs99zhhEqyiDWes/iiagiAl3ztf2hu8fqllhhYqVD5/1uE
M/X64cSW34rzcxSEw0z1RX6jSOwkcmhEshH62rcXsRT92HGlQAJ4btCvlKpn
IPz9dgZFiN+2WfZunwol2W8jRAOtvm2Xx3E+uRS4p6j/GxgWITEfGHcvwQ1A
x+/ij8gm2wXMlpqk+pYnvNhSjfs9H47CIZk7FaKL1Ssbu+twpWMA1ZPiXAL3
gdK0kDm7K0H+SjIhCd7YSyLbtciR5Rsc3umvJmcMadp6PFDDW7opaLNHemN6
vwLMObxU81RT9uvhehMSnk6msnoKxTimAuBtDFKzXaFlu6OzRNeaBbcGo1Ul
+uixw5h00ZBV8VTqGcInkF3KqVuLXLG/ftalEFEDOo4FhaoKhdl4GxsJBTvI
PsmDZ1YPBtXNwS0gVSeUh/xlwushIbfcAZ7TfxD+SMoV1QgGc5BsFsnPU26d
OyTXJqhkCMZN7trMdeeMrA6VVv0vQL7uIr06dEDCAAEZXsYFoFKDwBymhbLp
BYkSbdHS32LlDlbKXzGjhNbMYgjrSwqvy+eAS6o87F1gWHHJcTuphQorp213
LYP2fJ0DcSYcrsuacDIRdEP+7DDtvcZCH/aifdno0JsGFdkoEM06ol8sdO4z
s8adikutVKf4P7/iGn28pPJpmuGnKbRgHDSRoY29owWmAabp7qjEeYpvg8v7
Fke2RlGLwAOaSVZkrZyKpoYaaedq/TOc82YUHgIc4zYycX6i4BcXYgiQCcje
d8L6HMGUBn5L1x1WRqux2s6ohWTQCCRWRIMiPh/nSg+YcLxMssUAF/GKQKTY
K/3zX5GKvfDigILp/s8YNUwyDELXFA9D4kT6saGtLlBkbqZsJno0t8B1d5bB
XArRVEVT9Y2j6liZ8nC/L2UExoaiAHsCXJ6aGl5Eg6PxoiFGWcHhmZoxbllA
7Y6gSP2SVhmdQ+k7xyiLPcUV/7AkYvHmWPxJzKXNEhy9J36kqvBNUTiJE/ye
nkXlObjgngC1mHACpAjeEsLDny5luBAckrfbUcg2ep0O9JvZDUovdHHfUCU4
Dt8SgM1em/HqCGKs9qrskgDe1fLMeDV5uIVfjT0hSRT/bbULAEQxB9I/LpkB
q37ghwhBT/40bRa4kiTQLulFYpb23FoAdo7DrG9qjTbBgNUEuSmCeaB1Ea5N
2S8kkjyA6Gg1GBoFclrdh+SvjQih3qEVykSA/jTL2eonCIwWNXPAHibgPkPz
S9hooJlNEo6dbzZdv677EjKwinZd/ugX6TsOGcP+84Mlrmw020vGwQmVmYfS
YZM9uUt755LmFfL/i1z2jTh2/L6G1k/SE4qZetE6zIU1iFO+KLqYlf1WCBGB
14ro+E3TmTUksgELBCGPa0sO9/xE9bTgdCsqEYEp62pC4CZ5miJ8AwaH4rIt
DyC+44yLmpkiZ1lcskP36HcfZQvAG7PC0I2ZGbKzZnNodRvXTDjKvNx1g7Ag
dJir2R33Gp/Y1ndQHJCKKLJKc1oP+cPe6/672xjlMSthcZk4ipKLRiEUy+KD
f9/XWbl/SPsFSTnKpakpABI8WkTLOKwitkugbHXTzvv7I6BzEPnxgaob/V1E
i5VxXBG1sXOZdnj629+M/bGIBM9g8xFiNiJ6rbCJ8ptcwFcnZHIGnh6Odxw4
LWxTCxYnSagRJr8UWmMpAqQJsGXUnBDBMPme0eb9onMp66vKuoAxUtQ4ZJ4Q
5h+4AedQ3vi0LQXUA3mq98iJp9Ut5hrMLaesyGSXZoEtWjk0H/w4GwFrPJqc
UXUaJ5MWuMdy0zNWOvknsNKNZGvmsapap079tiUfmCTJfWpVwPiHUcuZpCZx
z3S0uAYH3dcDnYBf16j+5+hUoZj/LnQOSngWcbLKjSusGafDCL6pxRmYKpc3
FgWlGI1hkKBck2Y6oFFa6TFLeJS+/W5ksRqzPhLnTsOnzF7UQTn2PHxnIfGO
9BcGHZVW3V/xtQBkrVA32M+nEtLpA/bEbetqr4IrGz5WT8jO32u3Lu/BZCy5
+IcYNXdCHSGWh1Yz7IlpXlHRsL2Ceh1ZCtuDe6hdtwXgGMM1dZl7OkPi64DS
VWM7Lvc5LYl1ya008g2n/xrv1G/Jh5RQn3gbW0BjGsyZL1DMs4viUpvCXRJA
wL7tv0YzBrLH3rDDCZzTt8fPsLHUWNWvNPl6CsRg+nH1mZxDTSUI/OAuTrrn
ndzZTM1yYYWmhmMZ8+bxWfCOBfhrZJRqttR2MeDBhtabh7s4YHnFO6TTAdXO
M1eeBXs8EA0ZCtyCmEwVy+Go/gLQFQveCQzg58Yi5rpW1pmOH4NyG2ZJRPOe
0Dbe5hxm8DqwULq9AZ2O5GMwZPMqomS/BwpWM4Sl2ua6aNx0vxNY/n15R8yJ
a+w+SpaE3E38MZUEDnvCkMxK8OaqYYWs7ZJrto+ttezABcGcOlIP09GlFIpw
fpn+XjQhAKNXEpSs7hOaoxw538dXqlpoDaF7f9JGTKsbT8O4uYD4xwNQaYjV
rsWpFt88E6Vy/ERjlZUuVYH6Iquq3yjR2R4ilLhdnPYxp/spFJRqpzC+XyLd
HQ0F7HwzlO7ETZqJpZVyIbxCd75+zfm7HK8oKSO84ddfYqbZXS/3+a/SJ4xB
+XNySwrq6L7OnfVOH+bjDf+KBV41EnR54XaRlD0/9yt0K/jWgNYxdO9Z9aY4
eLQy5CDKj7qYI66NXQGIZOky/UOYzMNQ+wrRZHdTkrtD7/qkfY49EAjOPqKb
86BGE+N91/XsDp5eAu35oA7BiwnEHC5/PnvQ0korbpH4TDi5RA5e8GAczQet
R6/5C8iX2635UgV887lhSpx5WeoAvYgy3N4scGRT3jWnwMrZQ2oMIh8Qgzk5
1/83brY9tp9qKH962mPtrlQUlmSIhn19XbiRw59ssAvKo6HYqo+1dlkAixAs
HJMfzKiKEu8vwBD4f85Lp7mDfi+PGX/dTiGV2vuwvNEUx+pUkMxBsH7yUIDq
oV8LQ8KXCp1vl8Knb2IaqZvQ3qyI5eNkvol7QOnzl5dXD4A0VGbgbIeEctHc
hSZHVFXLijXxwXv5sMB40RTIgp3PNHPP8JvPz1t0xq2OiGGCznK1rjK1nni6
AJ84XQtMvD6khQSqq+2qHBZ1ZyUxlzDzrRfjMb9Whg5o1SgKqthhnLBkjyqL
B9+aFdiqqakJjx9SQpuTaFyIysiyUgxNoKfTyPoeQcbr1uXaw1Z57zhQ452e
Qesy2lrl+5aebo5poA/WKMrKqakfNClgvlCmTUsj1YFTaadQCUJIusrWpvz7
BhyxS4OqIB/1Xp5uEgfwk+wlMFio36Q8U4hruu7A4M74uBtasNP4Rvv8Rypq
Hw9QINvJlolJY5xjvFQ+YiZhoVY6W6YRnVGDT4ohgCJ9SVQPKq4fgphX1aVu
ydp/xSiCn8pJgFarLaVGtYtDOCauGrhHyKlD5qj3U+R5x0zmP9dzMsdhDPpd
67gMtfPWM2AbN5W5BGxkC+MqiNN8j4YGCcP8pl67h2JrhG9+Ux1kzh2K5HDG
VL37n1mNmF4bBT3U1+gFkEjPgTROwNDs5VQHXZJRXSHEPyK4ekqGK5rnOL1t
ln7+3NWlPdLBwbm7lAqo8Xti2gmv4HFYkcf3rdQiMiImcQV1fPEKzoPoZLax
0W8M1miO9UFZ31SMTSpaOu4ofMyOJEErF1VUmwbpegBnJ9ZQg8LJvFhfjzAE
9vF1NhBbv3rEMtM+HG0kgTvYuzMqZsS5q++0/ASUwX+0GaHscQd83ulua5ds
cmTiBktBAva8Bc1vNYnZkEsMHkMyYs9tQKZTzwJjxNxRWUZnIOmKRDZjSK0+
5oZWWndqVQo5Nvbf9RziXGw1jovcu7kNyakUnVEeurvGm/DkNFac3qT+7XdW
eUjSCUmPfYblUe4HKzQnvSKJy//0rgcqyees0ebEhvKTmAd6r0mkTSe9qIcQ
0AMWXf3HwYOUdovCRWVVFNwHRX7lEWuNBqoDbFBaaRYsVN5GmVfXESFSN5WB
gUWbe0po2ie4jh9PNM2rWUIoRK3FHJp0Ju0vaa3lM2m/EeVZG4iUQWhaCd7T
qGpoDBAgu3lcfawtV0W9gcZtNAyBQQraizjA2TZeRMHNCs+DbBqw/uSOhzhf
vj2+taqVMNrPVzw2a2fcyv1VMilJBK6kJ0Hbq3gdgay+mDIcM7cSIsFzmdMV
ReHvGY9D9rBU/V4hM9/zxxiuQd/TADi6M0RHvVw57zD/VwUNeLLQHyFsmmBt
49ioQKfKOdqMBEhurtVw0VdIIpMNp93X4OJzzpbC9CwR9PCKQYiJkA/+kPUN
SHyF9n5DEGFFTBlHovu5oK4/uWcH776ueaxaPk/4P5dUaJ7VTEc6dfY6qaV4
A0z5HEkNXATzsYhIv896ZzAvkcmiUYVfQ7jUjvu/FdxOEafUCKNzmdA0muLg
TERrpjyA9lfRkcSjDGBrCsyiohMxTpO3Q8PqGAF7azsKKYVZ5YkaH1bcaaF2
WAiRdyrM6U2nXz5DaRKJU60UR+kbXpB9758/1R3iVROCXjHScUtNaV8esepf
1enIFXmwOStTIQxd+ReAeBl5WikRJyKMS1RPKa7pDus+PUVQPD0ly6uHnLn5
FpqClfjXAnzBZa3G9Ly0z++skykZPjjASzIZAOkNzcvXWSC1flXJxoShKPyo
p4Kr8+b9wGt4PH4PUpXfch9GRiccIqsXaomUEWJ/eKYu6FBDYCjuQF+qOeVH
6XTbD+32/D97AyT8tNVAEmwCORsDTCe0wJBxie6cms89zU5iYJNHpSbBuRoq
i1zOqCd/fm1IlMhbqRDcvFH0FbgA1ad31YeJgcjjymbUfte+gMelwEmSrU/W
IIE7+PyX/QSbMKEDBtp264ZE08QVzusUYWW/3o10h+qgT3OB3FkeKLngIOvg
A5s2tR0BqBB1vJdWlUfGxigNgwiRXD3tDrF0hShOCQL+QMzsOSigN24z+6wq
e1ANzmaWdWSuiZzY0BeirIcgRTxNoUz8d9hPqvc7AkiYMGOHl/w/ck3nmSd9
UtWqVRHr7pLFNdmGK4a/Uk9PMtfHXmb5QYMDF7KsnS0MrdMX6P7ySvOWL7EW
vE01QmBsPmmW/6Xn6c5auc/X2uXH0sfX4a4WWhvOkvrhKyrT0Pib5mRBwB9S
tisOB2o0qA0gqikSBX5iWmPiMgkciCjxbO3JYNC7BP3ZxcNDvWj0wGc8MX8L
fa7MTQA/pbAffNWjOKM+by/6OdcCrvWXWxn5NXUuW/L7jY1b8OT/tEj/fWcI
ngxo+IHgqielSYZaz5dRl1MIA5K6Qu5oXQeN1AMgsr03Aty+mPSWzamCop/l
Is6OCzPO7j47skCQrepHmA0unEXX4SvH+qfhUdcBuHaV4Tenz/kwDQ8N93Sv
9pNQ++B9mt/L8qrA0kLXJi8A5seqar96iirnOHb1+e6K14KblXO/dPbiYLIp
S4FqHEkaSFBfa33251rXDA2tJ6A5RBTZS+KhpIOVZ/vtOKvATYn95T8oTqK+
C6FE9qSsZoB7dQCyyh6V7Jf+Pzm+nFxC0Vc7fMwf295NUwt3biDzxuOBqZ7g
vo8dmL8IVJcSmjC6M5hMH7XpxXkExEomS+h+x+tuspi9y7tO0Sz5gYgAKKNY
N3SQ8SaVzObVH18Zn6JUd0EUub467TBWnVW5qzTwTOzRVSNtE8YMZnZ4jn2w
wh5wzXsrlV9PYivLdOtiLqI2pOGgMFqejN4Nsx84B+tPm1CB6uMYNZgo9LBa
0GK1iNOTgX8tddH3KrO+7BEWEXD6cwcpBddGifvxR3rJvtbTFY6L0BmWnCaf
qxN7uWUJVtUBJ/QZuRshsTfzUkDJbj8Aa77f7GNHSUhK+AiasOR1ZSE/b7Pe
p20rsYJPJTLSUH7OXnY/FROzftRkMuBEyaZRha257Xb9zMJ4E/N6I8IWL/1z
lXs5O/vHIu6/a4kni0TRIRF3d2ZjrAqTJxjtOeUqxrvmqX9O6O5M3BUsEB/A
wfKg+RHC47SEIDtprTA56d5GB5l9uS/WP8SokMP241GgCFF7rHV3qjkLEJcg
SOl8ywclvQVDGzx60X5AdZGeHddE4zp3MbM9yypE/Kpvzx3SdvvSub8wXYNY
icIVoUR13crHj+EBYk4NjBCoyNvWV9WViTNEV/SJVVI1mhG5RiHTxc32J/BV
4Fj7Z2q9iwW2Xfzzo0nYsoEIzhXTw0/b0Ij/9s+OCnkKKAxMRIsE+Mf4nJo+
2FvXxD5qaVUXSnB1CvZ0tlNk9uK4yhbLNXa6K2ZNEZ1g6B5Q1cEzeppvkbUD
EzCrhaOLn0x0BR1r8R86ueVlzL3vyt1MoqIuHt0ZMKPxkxE3TNlz3Pky1HP2
iOclPCDW0Q88yP/xsJfwwk4B9W3GeeSZ/6t1/vaMLO5Gs9u8ncoPX5cDbMQT
v3id0XdKfOE1ZZmVkQ71mdk4E+Bu6GiP97yktXDCoejgbE58MyMQ4eZru4B8
aXqJzEelhITB+EpIzxV1KnhmlgPCEQZ8arJhoP8NLrXr+1IkImxNmd6fG6WW
O3kqKk9Fai0emXPXNBpkEKeCsUTU9L/zvawLwXSwiEdmmEYwBpVQD9fdMnN8
rvP5D5/4fkBNMAdBq/vcPkMJhcrkjDeNENFGmYSa+bH85EUjdVGTaQ6SMp89
zmc+nZ540isqff73Xn82m3Jx9l/G32jyEyj7x8Nw6fbwpv8J4FUjC90SrdoA
TKWRMMi/nIKZxsfMUmes/PcyOUhQtPX+41R3jjAOPeWQTQAFqqD5Rhb9Bvo8
Y9CH2xKWYoy7/K3cPfFT4OS7q7qMVq0MGAK53WoXNMUVmPuSDoLm1Ycfu9v/
x9CpWi+RR+uwZ8DaJJUuDKRu+dEU2VrgYVQnFxZzkF0wB1rNFxE8J2AQN5M2
2FSKfQ8g3kV/u/fe99bXvBhg9ma96dSgv2sJ9CoDPBvxSy/rosIZhOprtwCT
dh7Zd/48IKrDSSN0tnT5aVeUqAX1nhZRo77zeLkzwHWX0d895gmnJvZf0xYM
SwMX0gq0FgqCJeMsDDOtkKTlUx0UraMQpcG6aRb/x7bGwIFDnA7fgSlgvnLm
JJLuTfcdDXFF93gOqpQEcMLRokxkSuFoVpBFukCsb3A2Al0RKVTfjpVJNxpF
s6fvtd9AOY8wsS1wjhCsrtrHVERed4NXk4Irb5o2ASYFr9vo0HTzuhZJS0rg
hCn3QKbgZlQ0ei9/N+gBH9wnrck874m5eI8I9G1qhURQnTzUedh5+5AkX2JK
N8axCO77mJ3+gDXRm75uVJkUWXl+JcC99ae63rYOSwgbIqkt8Nhe0Xt9CzDj
qIYZxfnPeL+T55xadZQLqINAu4mAkqOUAhbSuBo3FQVQEQi4+9f1aWn7Ox/l
QVxCaZ7vPAJupmfN7QJrpshpnhb7IW150jnBfm8V9pvw82MVPYHPLBtMmVBk
WnFp0CjLEJc6uKDSdKk89edFt1k8GO2qeXXNe8/kZKqyfmhe/dsXVuF7Nw/C
YEndC3aSGdTH4jHq+BDo27qGMV4ztEtmV185g6qAxolCQtcAAwoeOffyUCaU
Me3O94aG9F7c3tuZR8jzn8BjmvP4CEknHQj35dFG0ReMqP23TdKZXW/2JPak
LVY9iOF6/tuyBpRzT15PhCXnAuaBUtDeLuLx6TlAzQR1Rb2tne33XUsjSBkU
naLpc73Yp1lfmjxTxAovi7G7u+wNL0fUt0lIRsRlZJeSYh4kmDIwGjs6CBP8
FaI8wB89giXLEsJ+sZcyQshc3ujEtTpP1b6yzRaHJsmZqyESAEa3GIF/INJC
0k5Tz4vafrFGjKnEMqdd3RUkpJK0hZkKrFG26vFVfhbsnP0XCgHQKCP7bJhp
Ln2IzSZoaH7oDehRux3bXnmQqxCfOdOVRA3TMN1Bu+YgXvyhufgnO03NxSYE
2SMGX8V04MlQk1WJt9X7FziakM2LUZqenx2WLTHpAGg3bdYacQWZsJrOEEK3
fTuXei9WkxnubIZgEb3BqS1mn/dhCeo3xhXERb3Cuf+6RTmhmjXGLcnb1vxn
069dPK0tPQs2m6cHFEnI6/l2lhQoYiCPdmYjUrql20vR5gaVBUQpVWOyFf0f
7PpUbD8i9/HvrBoQ0osFvUxp7azcfrRiUiaej5wUfh6xXgkwc6wS7Y8m5ZK5
tME1M4KO6Fv2JU70Bies9q+vB977G9Jvf9NOTrnBzwWDHNUV1pem+G8PIhLA
LtR7AqSLhrt68WnXzrRi9AgllOF97LIBkE923/aPdnwwW2kpUFdZ+ffnci2I
+6cro2MxaB6dpEPFZ1uYL63ciCZj9zpBq2ZAlqkQo6BylUOwCm5icr/gsCoB
CQ8nPHNia1hnWMYDK0i8jXPXGMZR3cxXdSc8qcfgW/BBPPaf/lf3GrMlCGM1
Ut2FbyOwUnOs9vegbQ+Qcv211Z+aSqhkWhRksxQWbwFGCN6a54YPTf++Pb3o
kdi8NROi4EIMRie6KBtpLKlveEOpNzz9+yKwQsPAnI18rQOgb4F0wMqhIqmk
aNO0yxNYXJPzR61bhucVv9zbiW684HHHFynK1DDbpCRhYWBLXMXx3wHa/BFT
CoRUISW4GoFjsECNRtgKPFsL/9QdJnkW3wwZQipYl311idEZ5lm7XsP6rx/9
wplXnm3fqAGyNJfiHYZS6/diHO4GwYgnRN4CAP5gfSTKoEkfG/goxqMw4IyD
EgAhA9sBWS5wg3pC/pZh6thU5QUdqIz15eMsLfEnAri6QMVc7lLUmVk37/fb
cO7GZHJltmcSixRZWxuFdRaihS1ly288fUqfKsdNJbvdsYAwQ4fRSS9aI9nZ
xDyomOGYwF7PnQGWHZjF9Lvh6N+OiQY6Fq1eYdyJVg1G0MLWTG9mlcMD1JZ3
xLOtq5BxCD1899Cf+bWTkMNOJDSCLS1t7feMQitArY2cp7hIo1ZCCTuIhOr+
+Z1IMyPfkXkh6CoDpcAqWgEk7avJPEPopSu+/sYrIdSS3N6f2xTAEtDm1gnP
9UN8JXB/2YFoVCyG1B9b1rOQiiPMnVZX7Yy/IfQpQCJm0hgHbfhMg0uGEteR
fhWGSLviSnP4Pla2EKMh9Q4Gbz5pP8GFtSUPUB/sEokklUZGN/QNJ3kIGZJH
xX8npbj66O1utJ3sHRwCwkp03szrR6JjIhR60UoQ1Q05x+KxlVRpk+mHZHQg
9aq3VaJWYdpkYA+871n2dkEasDXDfWlJ42ieOwp76I9rOhnIetDaBCuUF2y8
DU9G3fjAvsGjhDqJ77Gz1Xr5WxiDHDi7PIh1iuJwim9a4CsXSA3WTelPPyfk
lw9DqN1iIPzk1x9SW+JdZCDXQWmzjDf/fCDg6qmpoG1gP9wtiYK3l4bVfHRk
ZssvXT+APVzo1xHsI/JBZ+eW6Y+xrOzuwNOvhSleza/ShEvuaK59TllS1o4a
tZKEi6DmcQe9lS+uP7ZlCST0X6blutDwZxCEUy58IFe3Wv4+i0b2fd7vQp88
+aAd6S7Y8HEstX4oU7yLKBMiaRJBj1c7ylpQBGpD5LiMqe6EcFwBhSmI94Y6
1EeGz+9WI3Z0vLiGQo1GJlFbdpy95zdtKV+3rWH5iEwlqStQJ8lioOTHmIcW
jQJTHibxSiOueLgjeQsRB48O7PXBGIUT/LRRKoc7txcAed+o2U3E2unbTtMd
0x9rQqVkcaYShYq7Vjl0F2kwLADxfW7VMnpvetcWaH/BKW3BOqo32QotfibB
8DZWmGtKdO6XaCxdTxJ0kCe9SxgC2Cdf3s4gg5+CNy9VaEm9UEq40+HEeZcX
cVRZPqW4zhtZfcUbf8ZvzI82VTJdoQgkoOD7wBt3ACMjF1lrP8xyBxy7hLHV
Hw+PqnfLzmkbWpA5MBwjCp/tRplAkQvt1mu73gy+KEwJv2+d+i5r5FK11Okg
QTQ5t6+4859Zlnx0B1UgngmBiXGMDp2kxNkm4rrnR1u7Cf2oP7JrlnSbc2OY
S9IV3dIi/GiqkyIO8b3dqhiFrnhMxCUDX+f1j0h9C1+902EdbtJshoJFzNhN
F/T3LeEB8Gi7iuA32p/ab5T2TbeyCbidFIr239gQaBKxNWcwMXmv5tkJyT50
9thaGQFd3G/Rsh8ooyzWxTTpfskHtrq6mIr3a+4Frm5TD7RRrJ6/r8XMWVte
eVvhyCN8PgF0BOeEZSk0g0z2uqIODYYSW99AHKix9C2EjiEl+fIKKwxxf7eb
Ip4g9qIu2Y2svYEHiHdxHmClGKmGL3BCKKNhHiGuC10eFeuWzxaHBbiq9ZcO
11AzLZk7TxdevYagf+/LqH2EqDbq30fvwarCls0rhVRQJ0KM2XP+Prt0zS49
IFKRz2T4J/zIc81n7nTCFkXgP0T/gu6PtMZLBvl1cPPVO5AsYt9XhcQ1qVdR
9M6Cb3QqHHTepoD2CpAGZT6IKxe1nqlsYNUCtTNLE5jTjBj9VhmYhpiCb8a0
rYXYtaURPOYyePlStvI6GcDwktm3KhiriHxpB13g9cDOYv0x2pJyj0aRQz3c
1AXo6imVPSmmYY5BGMTJthl6nMX5oacHMIzGq9J8hhwOh6mSE9aer3lDMCCW
DKxBu/ZZf+egot76IUOgheqr5tvKMwRBBUmXYGvy3Rx6n3tysnR/y80uxvOC
QgoqqXJRx0b6VCTaRjoz24Z4IRs8XjvvMKnCsEmnWzs96FCtHLWq3n/L4gJV
1zZ5ECdJcYJdG5H+x6cPHe1NH9rrnSmDtXGRql42K5nUMlwKIebmCsClt/rm
crzEP2dwurLsP7HYt4jRsYnNOLYZh2Zkw4a+UdBen/PdILDqWyZIsKddxD6Y
RGgpGV/jZiS1mtuEFLATHkqGynjaLsQ2LxYxGWPY9TNGEy18AkvN535//l70
J4tj1JnjK+PR8/3aIPHDEiGHyntLyoNoHSoXR0QwjnQBzSjzlRCSFQ2Xoe1E
QzqlV7ZhGI+tMSZlXYjBsj+Ti/NZYDg2i0osibzqQqDQUrVj83nqHC3tWz8b
YMVWyyusLjlE73zM7oGDe6iL/l5PSkErZBedwDkJc536VmUPbrCWZymQqasR
97YRIwSBqMGb7SqJsywFuV1biVaE4rRuX3twtxf6usI5yTjUXyNI4hz1SGHI
dGSG2xBhpbnnNQj870xh8LSV0DAoGX+GbNmK5OcGPRNZpdnXHq2BBWS4pNeA
vLXHl/mjqVrPzyeBMoZLHvwkf/0ppVSQ/uNBS5Ya5zwjFef3CCRUI277G9P1
D5CgfpMThSg6S8mBtfm81nkS6YCjQKYCBKR0l+X3oiGnzqFaOSIytUWbOhUQ
29Bj0/7F0qFIViY7WzU1Bnv1BKNad9/JVSKhLqyYG7/qzjxABFkKHVCk1isU
sPGtmzEWlbyPpIJi65mM3p0THbT+Zin9j2mC4syL6Y2rcLn8u+eaZq4LiZx9
l01V7nO3mSML1naQsxdJuw4AfY64RYGjr9CGKzMD2uKyFYgMXZdcIbiv3gzQ
cMRsp4C8rxmKHUxRi66n2QSRP3fjvIitQuRMz+j8Z3k5laMMiqAfoWAa6kKR
spshZmtFadyQ/szG7F7/nrcIBX6ZDkuL8QSjnojbFNmN7TWcmf5o1KWg8Z8Q
oVLgDk5nvmkKPzIS+51jO2LuoIVJLmEkSxDrgkprO7y2cCLpxhbaJZVaQQJa
RALbFU1/UhAqOhfjFcyZchFPozp42ILOchgXyWs91NF+RQVRovZxBPzpT2wg
3FKvNGcuY1z/iGAPF01iSNaH5O20uDFrz8cKJo7ItGPM4ikZL6OhyIVw8z9K
GZsB608QtJUZs1aWCUKccd86YUzyeulz7zSm102ss73gWjqaPvr3EYGK6rtF
PPNfORcXVhIuCY0emjVbAhnq+01Sq17zTa4V/aE3Zp3yAq56UEIyV1H41VUC
TwH+M6iSuY1sIZb9qIllEQDt8KijL+yjwmk9Ea3yEiY+08lnMCZ2+WZNv7uw
ZUQ4+5ppFXiLakRfaDB/GMb0MvT7iYeimZL/Fq2rZWYGoLrMGtKtd2llk3r9
1gj6DPbJlNhsfWwp7bKFZQY7FHmEWLNesD4BsilWcxcubTqX2DJMjmLBv3Fk
TcIMEqiMjwulZeBkTnaMExx63aVlHqC9PioYOl0P3vnMuxWsmnOfeOeAu0UU
MSG47nAjxGL70099RKikvoHHWyYPZNFoLNrBZ3OYQUIatMA34434RbM999CK
GEpyPomGAVbxdbOQGedC+x/DM81q9aC2cRhrYZRSmg91ylbJrH85WGNBgSx0
lPUg//lUAlcZUVAK1mmL/Wdc04M6vFVRaTCoYDzqF4QYv524nZ+FSMuyTDwN
AqO4tRHtmnI7nuk58bE1LqMl7KcXm72GzSb2NsxDZO9mkqw1y02VM3pTbR3e
wuVSV5G3BqhbmgSvEDWvorKhTafQ5VyyZ49nbdXDtAr2wlBXw7tJYgAhYARX
V46b6fRWf1ZraxJRKcAIsz8qF5n4C9UA62TK5z+YzuZCVPq1c0dPrvz7PNGn
i9iR93pqj4pIryUpXhCsEXkkyeqgdv/4fyU4HHA2/YJcHUs2CDxWyCrrox4F
835wUWUg/mWOB/ROe6JAgeTeVBUQM4/7YPsfdMFyiQxHsHPUCqvxlr7/yqWr
G2a2ZJcfqe7Hd6Hs4eqDNXY3PvGYUq7H5HafJgT1ypd86+SAxME7Ez0IdNXv
WjqIYhRkQwU5p1vjr0LbxkgigJu9BIDTntdo1MlJBL7Ck+tlcLcy5oMFZXNa
T/81KS5arg6JS9LUyPaYIsZaXf9Oq3cO+2k8cEqsVjSx/rkByXJLlkRZiG9X
o2j70c6D+HjKwXKn37xLSzMfhaFnobYXcMsnVFT6kndbWMtt3B8RpAsoADS6
M1X6o7xmt4c9KFTFfM0UrbnEQ3Gcy++CaizdxFDxinQdbJpVakxCSqbzzl8N
PtOcIITPaHWlNOk06XjypyzBPpwIvL/k0U65OSuwFSZpEQmrRlwjZ/f5d6xq
NwqX1tVCbMyoHHSl6r0oufeOt8y75ddezw1JYLeJFH0SD/F2AI8WuwkO1ru1
gUrqya+Nx63yB49Z03OEaHvby442R7Zl+uQnEiR1vOwwt711FR7UBkQDg6Dq
sjiUGclzkTOBbebeQn6IO+G3J+GE9reh/KQNNx6kradtjR10XigccWkLCNjh
UXk0hOvSHdBtKldrPPv/8MiuAICEdzhe5/J/ROArGi1llnU9AvltkdYUanzn
+XniBzkFziC0PbnDomE6Fh40THZe0joZT0llM+XanGJ/+3XuJiNtfmDMcydz
UFGEKyAGMJMg4AuoYeZS5DLTzBlX0Aa84bBKXodCAB6WsRHDyNLTflEEnoli
jT8pza++c5vigv0swM38hUeKq3qFZ4aU9ITkoxHReqdPdguFmZjpAoN/X89N
U77JuX9LHZ43o/MIMXAcOZSqgz+f+VSTFNCoKJmurOgGzBVPkjqnReuCgFq8
xo4CXA0EYTXy3tIDMv/bAPY63Gubep+1vGd9AlmccwTaZF4vlTZ7kz1dHZmW
1QeJ+nspt6VBDpw1VtH1L2GBDw+TaHdXwRRy8oK5C/ZikSj/j/zE/dlci0x6
hs9Qew6USG5dHwYmM5QEm/oQAN7cKtl2u0Y42qodZe/oOxVBVM0Fhlt0U0dU
jpEj10Oh5wUhrUwKO6D9cCbk6Yw4QmKrb6ZU+T3PeAhroH/ASBF2DMfuXf30
DR6CvnABbmNv9/naFS2GPY7mexHNbZVZYHOTh7+C6cuOdb9WX1C2PdApV6DZ
USkWU0c/ualkVEfD0Os7fatQeEIUQSwmbVtTp11mkqDESHscbr7GU4K91XMm
9J6Y/OkThZqBIitYB3GDOTS/dNJ4NjMm8Sk+3IgYPI6ZCWpv0j7mF9Jk///3
MyjiQoGq7+zTeVe3NtjuvOnlgw8+PTnC7Ws4SDh+NFDtcbIfkngbWJgpMBmW
0jQUO9FCS6ul6q/Ff2wQFaEZ87t6ruj17fd5yViAtSpb+2GfRRckSuUJrz+p
W69DsEPBjl26K9RvJEd22C5Ierc6CpJldWMz5gJR8xmm4D8Ed/jVdrgp0IJ6
HQxBfilnDd5U6cz40Cgt8o3sYaXu77a/aH2ZkBXkhkQhWYo2HuuozDUDIN1b
8SAMTtAQb+Dau9MA6GUvnDn1ZTR4s3llxnPEtn2Ur22ou1KlgT+hccQyymzD
0prfqI/b0qC1WoaZ6mne81nY38/4dWKC1ZkbFFwiVIJwglyl3gM95HbilTGq
56EH/5ALJfNqI2JcNlDIKPfr/mxmjNOG9kvMwuyJUaNrYPYkeT1Dh+H9iOfR
Vpgvn27GDjqnQJPj+0E9XRAuvNutm8RIYHFMuwA7yDvJsDN0fhTzJW6DJqiC
dSzf5GOW3ePj4l99RE831XD2crdc+zRE33+y7V8jKYW0xeagK9LcT/DH651h
+5e3MO2P6fqa4Fq69TEFPLuOY24Pc2dJBYu1k0r0uRpEgufSP6eYVwHnPXU7
g4equz+eke6Y87kgi8bQsA+v1PEUod1RELVV1kif01bvrhTIc2UuIYJHHi23
30z9W07W3T3SbD0g0P4iFqGB4tL5H3w4gmySVSSVtnkDSA5swO9XI1I1IY/Y
55vFUF8uuSw3na/voByW6/3vbMrx68WEfn/oDPcdsmpm2EFUdWwB2MR4IALN
XMAIh95kQwbwAvGkvZ9Fn2S3bbU0LeefZKoBsq6OzAdwV+Azf8ijlxCJs2VY
CgEL+PjYBeBnzcUi33LDuGFWc/3kZb14MvdJyciYC9qMqh1xr6ltzNfT2YcB
OMvvRycA7yAuGYs76xde5INw1Fk4VzLxSVyyfgvL1inJQDqlAh0DBIeEIJ2A
hpusrL73MOq/hM6q8CRaMpsHUTM7GaSvJyRhOXAIpx/fRafCvNWjxQ2DgCzW
otpYfolgGkYjHijqz+og1J+kf4TophpxqauXP2Eb909iimxoAnjL1LdmtTUz
3eViDdZp5BQDvKxSAaYeBbdBNjpEAmzVnMHKCbKpMmlr7bzA6z7MoefoRaEi
qGydH83TdMHva5m33ResJvVJQVCcXwGxZF5U9U5mAzEQxLmtnT4cVIOaJY4D
RqVGlheWtapVHEyamLfO3O1drkW6u5cQXFi2q1chYZ8IEJIji2/tJpUSjMER
3Fi1gYwvhYYvu3dDxemdLrrCHfE3dlBWkLH/e7Wyz075hZNPXL3PcQUDaC3g
V7me4/f0OdaWGdjycRUSH4bCjBP7ql/1Qp/+j9T9tBJiS9IyWDdbFNWVWj0H
wLO7Eo6cTV4qH+MH78VZTsgC7wRRaHyc4VK1d/YC0yiNoaurupwF4pTrWsYR
5SFHluC1KgeNuzLk9Vku8IuS85RBzAHYPka97mALL+ntK4wxkwADUiOVNDQU
evKcNDXqwphvdxptvRe0HjSHDZYsfaq14Br0J0NlpTjbTKgB3N3Zsye11/gH
+W+es4PemGsIhra64G9/ZbP6D/eqAUNV/J7LvItQE1J8c1792gJtMa5sEIvi
zyVCCH1XCHRK+nb5TFEWq60visR5q5KV3Q25sYoJH1wsARe6Wn6GzRjvSlil
fGqACaO6NAczLWfgFZDYE3zH74Vr1sXqNuXeyQhfpKWcUuuiDglM4yDbDL2q
4IEl75UAJxhPN5mUwqvEUD7vfDv/fQWt6vqAZqRTLEGJ8ZQ07TRrDY+QJRUW
xmuNAQ+RIUAX0VqX7/btMsG9NxAZTj6ssFDk0CKXtJ2OOKCyOlGfAzeLwDhO
Du0kEACDU8Qqo2KMUJWw0VYs3VwNzBRwy9vvXmpDm0Pbajv9vyBXA4M9tk9C
doMDEwrlCpo5uCTIzjzmDDd2tfj6vgzgvzoXgLGj6WJ5TtUwTecegbnmnljX
lskXj2I8dO9PD7ENpBcsvNX3AxPO4+ESHCQyk8VHjxeO82Exf1OxeYKBKc5A
KcJl/QjdkXmlVaFapRHoezicVzjsMWRMtYyyxpqZnYWXsspZSJkrkCRe04pY
eY4yXqq7ELe7WogSgBJ19ezkTaHPyvr8Y3GOqckNCQyKvEqha9+f+a6Ftf79
B9yIUCvHHuqM/T26hqh2tPB5o8wpRyyD2q9lENaMwngv+iwZo22FKO/UyRnq
OMkHsJwuiWUtgjpu3uiUd6eA3S8yGhbF6YF7XuxN3CuYsFowb0Yp3k/CQdn3
MEyBrCxdNb/vK4u1pNi25D0OgxJKNTNeh+bUwj+uxrTaJoEjKzXcnw60ZKMC
OU4+E0J/dvCuTfSDYKLjy1gUpHFaarW1K7p3OPvuwqEUave1x6J749Q7Xm35
SrJ8+P1K1ztNVaphjE3m6cg/S1y0WLaLe1o0N2YzBrg2Hm1kOOnEYeImI1Kg
PVqmFTsbBTweVQILy3Uvjqy3KDS3qz1nYS0JZhORrh+Zld6EZPDaVPrF9oXL
WIxsIPUzLzZpKmTZzgsuAFBn93QCbxLQXRK89dIj0onFK7dwhSiyS7c1Fxh5
MHIML0RP+tXLPfG7GP0s34CTX1LEL+0zXNPyzyn9dTw+o53QJdLOKBCEHjLs
KWG18PQV/DxwUiQ6BT43LOjfKfi7DN4O1tzYJLj1m3go+y9NigC9iPvMqChP
ff4viyzcQgZ5kA+J90rgCBquoAvIPNyiksHR33McdV1368G6cDoIMyIMj6yZ
VbXedgqQ2i8mKdX5fGyfGFf6wdDW4TzkGPyhBoBwzV67KJFGMDgWqatdpQ0C
+ircbUUeDYs/ZwvIBvuCK00o6k117juwPv0qtpEqhXCgTynWUxAek0+v6Wni
czAoqPv+hgvn2Yh1dB8sSvXD8ngI3Ez69I4z2KQvsbBIic+TkYIw8ph9nXt3
6AEuN1VuP4rZyOUAgQQHirAqjUU09EmRcYfm4JMigiCMdxi+ZtgvS8hs1nY+
/+fZJ+nqPb447p49vhXKBDxSN0UHqNdT73txPema0yY5MODHOb2kHqFbRZ3W
0yGsticPnia9wiYsLZBqH7/kFhMPS7qAzPkD2ZCrVIuwKr0QR/kCSBhIBAve
JOBuSqwqGI4OEOwFIbzxdeJvG5/lWurckc8ZNrDSBEHSVrJHTEnlIFNuLBoM
20BmdonIRzfhk8dXRjGvzmObu7BcO3SWLBpxdE1VtzxdU0ir3iIDN635d4Nx
tmdR2VOmfdKUVCP3QRVk8NxzOUjx8kccP8ZWejES09IvQT2QN9BcoFLFEmYJ
22z5AHxEjKzlZ/YbSQvzhudV+abjW0YizijTTXYRzYIUzUexdu+cgS/yBiqo
Z2iZuaSWrLq82DJj9x1DgtF1AG+qsyGdwGOiPesKE2NKmHyozTMBGA0LB2AA
GmR7EXGmIRvp3CKA9voQnjZiRJP4Lv87Grl36RSo2kDS/Q2QHlF2ZCj0L4fr
dsPCXlJszwq0bDoRF16oNR+xWFTF64KiXh8aEzCEx1wcS8QZVPUsbpPlmSgd
Z2I9vwTvU7E6cTaHjY+xMp92Vjde/3rkdIey95uUTVy8FVqWid8ObIY5SAQy
fPrRxt08RIwWeY6Igf8+1LgfGgO/+uj5exbzjSA4ZpIgD4X4/I2fs5NYaeRq
dODdYScupBgDlVllKBJLgpAxe3NUBBmAS+jtXlBF2r9YUiVEbVQFszaa3KZY
xEJ2xqJOAsUmzx1gPC7M94MukStI5IiIz5lEEEiafJ7F4ABeeKx3Z0pklynd
YmyH0ogrDchfLJ/xDy2er9dpHLFQWpvwC471IMk+K8BlLKojWsFuITZYeHYC
alh6cHLwW27tE/u1mzz95JUgFTwG9W0RIkM33rM0I9NR9PxOjcrwryv590HI
jSpFFYDUeoNpF7kTlhpe+HvvNBK4Vjkx32M7VSYYM/fc6bKglIkeZ0vLzQFP
XiyZlMO6ZxFbhW2kopFrNR9Yib8n1qWok5wHG+HU/MsegPRlJN4/uOI47z1I
eWkh46GLfLrcHniOmKVn+koOybcJ+3uLwUuMk7E/9cGK+NgSH9QsDKBln2KK
+4xm/YT9gK5/SnAD5CZPFzAGoMvViBV0ECBRi/UVLKICbvJB0Wy7a3OlCqQ0
f61/g/I21X1raDyM8pCmrgU9whAF5JxrvozsQl7q+vCsNt77bNhUUQ2J8L7S
rVRUWdx9bnsItBY2MDZgSbBZeHgPDX//KJEDRszmuN3elXgmwbscQVwnj5e/
DR4X2N58EvOO60HbU/nUzsockNcy2tgwq4w4ClsOF+sRcScdvpk8apuSghOT
ne/haSMhn9k6cMGjW+rSWNAeEYj9+2KqeTfCV3zmjpR4gIrUqid/oiRu+9GB
JIut0DyU77pghEA/ig0fucylsy/wWM4XIzKfnyvYXiWmsqw4VyCQt8KrqIDY
cIMQPap+Cv35uIMCaivPsAYNZzrAF0c71cwog3zZIrHnwnb18iIibRpw+3Xw
57fY+Vb4E2/4ENtfyoR8IUEx54t6lDRKkUbet+y+wvfjuuFGMZigLthjdu9o
4rrGavf5uNYhLYkfbRDhPY9lLvRXoQH2jEOMIz84i3WRVdgp4f8hqcCRTFmz
90LMN6ygBoDC49YLDYaLU5Ix1A64s56JkzTm+pxGOL+1G96Bv7Kl9HsIZ2R6
Yv5KZOULDw5ZaleDI50O8BPkuOL8WuyaulyLE+65KfG10UPNxffVuRuSwQTo
c9qdrL6Byb4wYvPUOfKxxTc0jmBhC4EhXd13/vzxLFLLxHaQaDG5GgGgCyHb
OAHwgvqzr1z+0jQmYn6XeQsYoi6sY8lVDS6OKDfHNYkvjZEjpnRdUZ1aSp9+
ag5HLmbDc0wrdLRXi24Hd+S/yLK6N1WFHn8nGEkuxk79NeodLCIMEStzzn/n
P3aLc+BSZqAFIqJ9msp56ze0fn+FztRWUqdW820tF3kN4gJu77ncM6N/N1Du
jbixzMvkyHLwJzpPBTynpF0VzPaSwvwpapqfw5r5ni3/uHw0npUJL4115YFo
/Z5j2ZCWfvERtvWS6Pmf5izZua7mk/V3WFaEYFgi70pyG5qhuGHS+AyellQk
wKiDmQSnHugPlrWWXjjhBjq9o9vTGd8q7054OHK+MI8GzC1QRuyJvqoy4OSz
x+a8qNMWlPm9FP+4xvG7phxeqfW9DLanYa5oXAaU2U286Ut7r1PBvMf4Kp0R
c3YE7Ah80xAueozIHXgTYxqIy2vP+Hbw6Zpi/mM3aeLHXxNELRfAgXcJGmuT
DFDrrHSTLCLsXSFgcZLZ8ay5gYZx14YCRCXrftTokE5Rd1vK36A/+z8UO+FZ
4akDP25ijJR/XcztwQtqR1OCWRptKxEini/Bamh+U7Q4qSQ1Lgu1t/WbftZn
PTX/pQw1uI0+wwL1TX9bePJfuxG0MeGNxrdgZhdYBkXRg4rUYX/Oajfuw8uX
Ivv98Si/trowYpnEH0I1Y7k0KUEhxHYwKfSXH+Q4eqhF9AtcObv4HkXSTcmb
hJ7nXe9EkTNLkFeYu5L3Z01qFxqu0+K/jnuI3kk/3MesEhsrAyHBeE5mUfy4
+53E3zQg9GZqhCkysjjqzonBErSl4L37LOqy6cc+7o53njdUQLg8aaWQU5PJ
h7L4Ej0DYJ/9XBpk+yCOawNb1uCikBjp0B37VZsDsmmIRLTKFGjXtFKaA0tO
3puSY/RXNNeYYOkPdJvk271CzhsM6p9QsB6YRzYojB8IuefbHBQuIfI87YwO
sE4+Rn01zMTi9/x1G6I7s+F+/ABaO9dyRfWWrwjpzzi3CVFyljGZWgRmfxzz
9tnvt/a0SB1mFAQmNej4Ye9bN8wf5ZcrybgAX7ygo4rhuSbxh0IBG28Vf6nm
nO7BlslcdtisDmB/RR1wGI+DMB0Al4IEX28z8kW9pzqfst2w5YnezWsgW+yS
XUhfefj5V2751uSmlNf8iDmz3bXGmpMYfQkPwjsIkge7MCeuxOHr9g8A822F
37pfEz4ndcFkyf8UrdO/5RNfZ01nYLvN4HAoH8A/3DBjklZDCNnlJBR8IPIs
g71Qf3URmA+AIfxQVRmm9gLRNrKduu2wbk7IoDJILH8/+ptpNgTRf+KYZnbj
Kf4XfBdWN12IvG/I81FZyn6oO1L4T1ekfspY45nbAbGDxbcKMABrrfj3Hl/6
zfPZn/lzdiwCD6Y7jdk3S5aP9SJzI8IMKf+ZpbzvOTCWu0dRkvIumNt9SMSS
lsZerAbw5XhsTIzhAcIsg9PDZFsnOvXtM4ZKqQgXQgZLxxPHc7A1FSSe72uh
0vr6sGJ+UYO5cjp4c1kVXyZFYUJ97Qk9cpkb6JW0X8JyZMZRi/lgM6TYd4Cb
mSBT3HBXveOJ8qEhahucbcv30dRLnvZVnxMKT78XmDpj+/Vf4GuTDJaEVGtV
dURaAirbv9arVIeBzUaNXSgEvfUA/16GB4Mput5ob31mKSoqkUif2Nm/DXqo
WT7HLoA4zW7Ia76mwvzMr8Tt5lxk2LKVb6Udxn6/rY7EwLqrVyR2P5C2ec+8
RvsOxi80NG2Ie/ubGJRT+49QQb5bQV6vtZWJITj7wkerOgCajMRByQWtKc6G
OjvjkgXiLomDmmTdvre81sz6otiHH5IKdn1HPJnocQrxJ0REcIZK3NhImUne
x1RvwnaI/ew2TAmHcjgd7UTb/jmCkZ97ZrA8L+eROcbhPaDouigFv4o5GjRU
5sJqgQgQyq4x5uk/EVmsE0aFA7yJQ83SiBDmju5onUQjtK+anaAR8Kt5Na22
q5hGzT5Ofyj86Qzn9t0AcvIbtt5DgTnTRt5+dUZf6ivxrlwOIu2svLme8ZKO
cehmNq8StGYbgUzEbQx539Au87C9MKSnv/M6UPNpzpJF1oFrAyEcztW9RMz3
dDg28tp19MPFYZeSJu0CA0fgceMzKrLz9xxVBeucIrutO2Q1HzmuKSf3Eu0h
0vOGF/uiAvANRLzamTwq94gXxzoKp/EZrTC1/63A4yJndM4C7guW4I5Pt+ph
4rotLG7nPCf6DkPrX9yBHfFZu5q3Rt+p3Cmasq4gMiTQAOoYrrK6sfoTtDJr
8ooga/hUATbSUfKTzYIdYsOtRoHR6QnVjOQ03vvTccMbNnKfHLWXd5awBDci
5GKSwCRXvUZkz6Wy8m59Qgm0KgQxCJ6IeMBHBLKE4qBSpaACD4SA0wWtrczR
8nKfdescVqmrzHH7R2v3c4TmBTzQqRRsK7W8OkiXgMKDw/1Nw9J9DwMe2Duz
C1ME1Su0jM4+VbAnSu1V/YRy1lU+r2D9RtlU3wd8yK3+PYZrZgBKpWDXdMn/
+IZEeXLLI7uO0/UOdwD7ddYI/lTup8Yks6jX6nBOQI+6Zp/xTYokoHzUPF3j
1VhJ3N3vSbIafzJLHjU99UaamBEfRgXI5NSzAyCIW32FcSKl7uNFIQOLpo+4
hspbUL2owPBALuBHsqXsFrXphSdW2lA5Q+0m0N7wX37alMuFEs+t8aLeD3Mg
LqIVckXr8D5Uj+pewn81E3oL5jdPh+Wfy04CYKT1Y/dL7qj3o++2R+mYzDVP
FuEcEdcW+si/3eunaL2J650WWchZa599ykrM82kjxYnINK8vka1DDo0fyzaR
KW5/arsNLEFcOB/bJRrgR5diRn/F4pUW/SBVhOCZw07KwamJlfaRqR8dnh9p
I+PsNFrD0ZNnzYJS2PrRFoqLxrBjwKQrrdA1kCK/yMS1OxdpoSpZUBUyxVOj
rtDk8qVjOc0/MMxx2hgSGS6uMCda7m94XqlVt7HMwTR7jig+NRgK7c5xtkMc
txk/a9idrCdsy36FIGE43JuXbgT3gpXS+mP5t0Mem8OEAFvxTvrHu3bcwX1B
dR+dzBF5m8aWzcW97ct+u12uO+XnqCNJOsk9ZLOCX5Lor6iWuX8JRgQxZgRX
hVxTLzLdGnzMSvgPog3AWskzxUmqK11CXhvQWGoP/m/ae47l8S9gO30gUwgA
gk8wj6VWX/IbVMVevRlLTrNmq0TI+AY6XeT9p5VynvAzlxLjjj17GQzNHnMe
Zxu8mNUfpLamLxzvKPEtihHfOvF5C+e783WDRGIQlZY/kcyGX9ugDM2Zznq2
OTrdJSpZyqVA2ssBySrEHYS3jwgxga+XqrHQpzNl8RkqiTKwhwSQxyWNLFfO
kGJT6YeaWSj1ivq7AkDVKBZCnpsqml6BWPXknDkn12HUn8/9I80Xhn5uHai+
vnnSlrBET77labw6PyMmC7Hrtix3tBszhdYLVUwmhJ7EikaUZEswfqNUAoJK
v5XGkKDrl6TosnftBPhzBd9fH7Doltu+oyW9r3dTWOdVq0lntY31RWNL20lC
z/hD7WwKSrSOktkO8/nKYNNkqcDMZxynYboBDTch7scqvQpODhw79FmX/SrR
/SupTmHGBC/qFyfa6aBWW+g/9Q/90FhWrA2TVhchE8Jai6F4dLHED345k4mp
WLsw+6Cwzo8Xuhopij5/gKtZhdfNuK8YKcPTFec5Dt1autOhoUgMkPdmFcgv
BVP+2nAfxWfr8SAA5EVYPCzKoYvYNf2LkTYumT8kS1YgDf0Dj4ie6vuftCWU
7ogiqJ4JZ5vQf51gRhQqbTH+sMUeazKQpv6Sbu3oWb0qeWS2+iq27eDjvGV7
TldIMVpnS8gGi3KtmlK9XbyoNjvITL1dxIP6OV/K6QJWKS9g9E3dCCMySeH2
FXtMm7C4ei3eI6jlFrhjiIPP5uKkRRb5RxcogjwH9s/8kaDHtXbLuD/pSLb5
zQxWoEUks7cchy9VVcu803fnSqioBVajMGXdTRNLG2TnsHegr8crcuuMayom
6Um/P6zQwhRXmom9tMw/WFisNRP7Hjx81DVQY4SGwatMd6HU1AobKlDrib0a
d3ZY3nOuBsmBz5lnDt+G7vtNvP6n7iluphxcQEMYf6pM4rMHJDP9Qm+QxmLD
SEgqGWtMvP7F4BUeqtx5pvqDGKIvSX+tiDtgQm6G5HWhHMK7x1jet/ietetl
QtQj+0N+/UK1o0c/MaZCvY5zbH+o5rp+87AEOR+/4WoAIHYKxkXI+Lz/uT6E
XzE+Habnr+ZWxNuaTahWR16jFFoDUgUx/7MjIBuL/g7l7rfrH9WqfzPREUSD
FiczRMRXybTYOxLSl+jNqFWoOu6JZSK9X0Y+HW83gOje9fOnrQXlTlbDKzRQ
0QYnCcs5+D71sFMRPBihBVQ8c/nSeBCQJDzvy8IRdi32hVOb5rGtiTvMKb59
jhUvCkYXUj3CA9hy9cs5x35mQ6SQCueZTdSEhA7U53+yvcQY4z5MYGm79Wx3
Ki6vae3gZmfphjmYxRZGZf9czpuu6bHU/240Waca1NBvTaYako+E/MkM8LbV
MwYZEDAVED5G1OSQqFBMvsv2ztgkJTZQrRgJaYN4lIXBBcjXam2yFK262Er/
P/bvmpMU4c3z+Q1jKfY8M7QyJYl4Ublt0JylHGl7nS/ycApVw74wbWScesJ+
X51sC1FYM6o/Gv1FCVNly6zVN/UCbRrlxnTr2lfefas78dWPwfr65gpcmC1s
GscYycCy384832aNnsmoP8UZ4xmtEWBqGzC3tGcM3MLJdfNQKgti40fxQb9t
tyeSDZraXd/R6o+MPCUr91Ro1g1iXmX9wrZZWK3LeH3NBflbS+Ua20AgTzU3
g+2zuqZeY2IpRnUaiSpXjVZf4ZXN7JLauR7jJPQ2amaWqkXbn5fq5p94VTPL
1fnHPyB+mX+7Rf+vjL71PjoK4/gwuT8Ld9cdAzHwERPfJfS6WvpNXNsj945l
myjXWCGsDxcXvi79fIR4RdxblVaQC62VGB98hx724/MJLgF4YaawTl9GYCoD
iOftSfEkDcO5MYfd1Cak7hg/OH5VU/WNdBo1ggV0UdZA2Es/U2z4i5ZlISig
Wf0dUZF087vRBey1vXKoa30dJmA4UNoqE4BeC0omH8f9pvvU+L2eWLNSfx7G
G3WhcjejyKRbGCKcNLh98VHOiOPgTYp3opv72w3hl0xP6SOdl7Y1rwHL+c5F
lcFjbsElK7NO0MH2iM4lpbNMQX8gbfYIMK5U5DUAZjM/Rj+Bpc5GVQhiPQSl
JB/A0Aw6hwZufFMiWtKoPC/Az4BuQqCAB8seNOlPfut46+CAsF1UWKCLVp2E
iPoiBwca9iY3L6hVc7fLxnx4r0ZQbyZ1qgTT9uFuDiDpgpyekTnBJcHVM9zk
05Q+b9Lv4N3czQ9yjBGfrjzkIcB+gu827q5hstI7J8GzFx/oaOEqY6lmNSSI
2kyCkDt/fpzMaig+DZPTiCM0AWqBCAQtOBiTTmZmmxJlxcZCrem464OfJ8H1
XJ+zDMzMfHqwu9HQy/YzjtLrRjIOeeRw9XzAKeQUCYq3NBcVGLNegNrtwgOe
euhbDZ90l7tg67CzaZ6o3DL0MxodPv847+DI+MV9CyRkYCNm+TZwI1GmiAs8
erso7Nr8thW+IpsI/uY9TvZwUqfNSdwchh6hAS83vZSuFP8cPHH89ExyTmRr
3QRbcArF2sJNYFxx3YlhuuoRiER0y0kbhAL95XUSYxJMHBuj0g67tYYwQciE
BX8UnjbHKij7vDXzQPF71D4S4M1L3th/e0ZC91L+B6G35hJkyNhe2qyICZ65
DDtkh93ltLJw6MuSRWfnKGNGp1Pi6+xI0eFAt9FtEA9ZjFv3UO45YTrNB4KK
KmOTxLGRybgm5ufl6hC+W+/KZmQ1iecvjXJG5ID3197A/2DtEhLewfAtXjP3
Y2nU2+V+Qm/DBzSYYI4dWqpruj3vxW/Ix7A83d2DWq12UGihCNNHwkDCwSRn
sh9lC7oIfTMVwfwByZGUEI42OFb7O47qHrJuJPhIDWosobrpWppP+PS6FMl1
Ag3wiySeihvCkr3BS6aFaI9qBa4wlJ1WXPS9mtTJHC9SwhAEVozxlS9+SQs8
Tx1AMMbvdMHsgyXcEYMmpojpT1FhiTgbgujONH3xK37fyGwt6TqIWFBLzx8w
VD5lJMePKo1cD+pt4/w+1qS9p/7wX3Xm1tWBNpUX7hHQ5Ip+TUvLY7LJs6+c
pocHp1Zs81xVXgmRpazC8kD+xFJ2kz5SUE5HoXKnm31McHUUXh9LCQG8NgQ6
c+yrasCT8xumFGXCAci9ioLrPTyvytxBXPwXE/Bnhyh6Svzqr1vgyeVCl8T0
rEwTTdgqVBJ1dFnfJZVTra2cV4xPTbqDAnAacAYUksNHI01HZNsBHAvw+DFS
Oz+ssPHlx/QRXM5S3GV6bBsYIUXW3dOEFbZyTpPE4DmJdkyKYYwEUgM8WoWA
9ErUT3qugMfB3i5daahuK0q7sQY9edN4PT39Iwn3+c4Rc4zqzrmmjX/4BOtP
9gUQsi9fcGUsQJNpe3uqFy3fGNZD3zxwPl+DwC1anJ3ROzmJNoXFkg4L2bpu
A8EC/4iosbFbYIp2CWRxe7j27aMpZ4vfuwVYrmdHGYsRm56qJMLViHMyNypv
DXQyBrt7/+fxstP4BTMaIraY5hmS6Blf9shxTGIy8T7sriiFeIAU2/T43Df+
ZemqKkX9BYd488pbEQt8jfIpv3Vkacf7cRaCyeWyAcc7bH0pMZAdpCVF0qB/
UJGkS/wQIo+jK1eSLo1XXv1OSrbJR4wVe3RyOuu/1dk8mWRT+uKZ/8/QicgX
XfUQ0rwCEwXfhi47KjgyRfc8ylyodMDTgKrf2MY0jy9v/NWlUZXySjJUj1DA
+HPgxaBu9RbPB9VGAoEK977GcYJh4CNkkKPJziy21Fvv05t8YUNf2Xlf+o31
B05rSvxYwqHcNKyEAN2DoHk+Y1CYa8eWjI+WO3+uUHLdcM/PTQnSDNx8/3Vb
f0MCd8kAwPeNdTcx2725zcsxigEv727VhQRXkp4vz7Sj2s3kUnbSGoBIUtQ9
DR65Tdx5StRlabcy08rjlvavwvg+IbMIVTMi4jQrgp8kgoYbXXaE4Mg6caeM
ykF24EqL6GjRpmV3HWJZ808wx5UVfXHfj9yAzc0K8szZIqHNh+XAEV1kfxvn
NZjn+QCjWuxoCaR6yKxUVosrJZXkye5FiJPHOHeN211vAmiiTI/2NYWmcpFM
/3CJKfB0It8NorU3E9R15TBxbv2QppziOs2hrGg9WT8pJ3HJ2JQxRojBPo2f
NNoVs2v5AdC8pJ4EgxiGotRao70I+gBlvq3HtF9QQrtzxJOWKaLQqhJhJ9VB
SS7zO6F55HtUsKivLpp+mHnEiplTImSlgi1jGVESbpVGFveG27p2yMZa6Gcm
y4CnZssbxfPksbwLTe/00GOtLFRmmp0h/RP1VdszwBQOvXGdZ35vq/xQ3QNz
kgE8SOdaLA8bJShcQMZBOyMuKjvYoerJuK+xZ7CMdqOKDBnLN4uO7pJsrzBx
nvmIgKlHOqvTZAo8m8JSOzvhVDJAWT9ULAtTU0qkN+ly5JFzFhJKm6oBsyzG
tKAXonZVKenczzuDDakBbp3uIz+xIf1nvJjCwLfK3YWC3xPE5YvuBT279wJe
QmFxam8FnTC7hClB5mwVUq7H8xZnKK7YIKwh7zQywFRviX0gAOg4wCrpVJhC
p3vbcEg/bzffVNMbdH65WFc9YBQQkDzwe52uwFVLO3AoVaLxqHCWhH56CJ3O
AjNPS93NKql5XEXWeksh/E55HusDZXvPaVMGotmlVfH5TpikFn+IqinWuk49
9no4tM4Nq98y4lQoeucdgV1YD0XLX61F34zr+/v3smMiQ+cOEUy7bEFRVkhE
gziM50VOTcUAdomJbpaLRCNYhc0by2/fWlA8AUI8KGevmVBYSpCyrO2hOZVf
L8lz38cEDo6TCGaWBUShvBahcgDFX1zurq1ToB1DGOAuy468A054zKrmyi2W
rMJBUJ7gI19KEUwBn4ZxTFE3/eOQUgkkcBeAfisgfDNICbTJh5aWbwYnPp9z
mCGs3nQzcTPQJ/rr7/idI5sI3flfN1xcqGsF7f24jIbsA78rgGjzY7hmV6z6
2y9I+ap8/MyjUlpmyx9JpCD6fiELiV15uvpqiMD8uDymVT4vwe5DMVzwadp7
1Ytj1WE3WHL+yvZZypY++qQAc22BbAql+OPQdNjur4WKe599Aj7gjtA4haQ4
6gPYf82lYZb2AAR+ECoqxwABs2qAOvOtLopr5FU96CMzhjqOe8vhE++2O+2n
746c4a8lhdlo95UoieDe/th3n10g/PMsCFXxYJTYVF0kP0fqZ5hLkHoGI7lO
w67ZgobDxyWggpFaX1sPt5So3tKjjD+cyL2QcbA43joDxA1ErPeDm8WxzWfS
QVCchY2Sl+zuiXct7CTu0qQW0jomaGiddn6C4xvHJhyeC0MrV+/XZhzrWMPR
VaTzl01odf+r8qNGIFDf7vesUlcHlwlyNR4MWOWiWcN2a8+cT+lkNulxoKI+
MkIKsz/GfiQuKF6xh148CJ9wLAmueu4ddoo4kxwqbx2yyFwsPvtrapvPb5v1
qfB7iSgJUwnWrauHL70MoWRN9bvQk59XNNNFdLPKyLnxt6crFSRTErTgLM1e
9DTIqDBWGQCX+ugA/V/wtgF6U98hDm5veotZ9KZ3kM42SE4NRLH1X7GjUoRn
I/Iyn6wjIUsyP8LNiG9abEmZdqrTal0qlOFB/avRsOiq02kJtc26X/dDbEOK
BypN5yE16+AnpTkV535ZgP5jvAjbh3LZZdHZrUctPYQN5pszzFVNHejbQ2jP
/jKIXmFgo3n5wUr2E84eEbtQmgSp63nYCgd6UsXaojdQXjW28MO3m9FGGP3o
775HPC7m/4T2VLjFV3lgpO4KYiYkwMPPK2ped9ZhgrRO/pDBMhPz76Za35rN
ySo0REy68ZtMwdNukKE+Pv9K7hJocsXjX5bmDJotbFj3Xi+Exljf705deXzC
tjNIsGY+OmVROnLDAiESC7Gj0RSQVqILQ6pC55ywdapuELvS5W7GRXNZUFPT
nKnO+e4pk3C9YekFFJZMZUH8o3Bd4Bp3Xc/KSgyzhrB8cvVTsSv3j5+HQmdJ
HrZzsJK1ucHcMtIvb5mTRtfzdAxNPxl0+CU3xeaeQwvHgv194n3Ql87H3MoY
ZR1L1Laig4NtFP8NMlSMOZoYpXV+mw1YnCPFC+O7Hqztta3c0etkNb/F9p58
Q7lYXCqR8BvmvaXxEMTHNQsWMai5h09Amkk2c6gIopER68liv9RuiLmXfTpe
vggmCHyMiq4tyKprxEdMBGYaeTqqvqmR/QAkW2Ao2jIBDB4e3RZIaqMc6d31
KQmSwbq5hqFwuzbSCWym44kw4j7Fv7s8Dnv0AgprFocxh6a/JgnrDCLK1GK5
YznjufbH15PLWvxge9hMSEjyMIB5bm9yLrVPmHs3LNin0chWcJkSrzNpxAPR
o4aM3JqdCAQXiS6IwkUv3PpdHLm2PmvqDdOT0W2lwJE41QfUHz9P7eKUz/H8
3seAtLeWeve8rgz8LCQf2PcegzsaaxGBpLwOA61EmzObLXi5I93D8bz5Xvfj
EaJ24kS2QjKR9AgsgBPMLzpMkcigyAbH5sYer6W5nG4fGRQfzyYIJXNV/O8t
L3I9NMXDL2MWUoGwg7Wvy7QXjFxYa0u3uOAFoxmspIVhg8htFyODP2LS9kAX
eauxsVfkiFPc67OC5dSbJLmOfQHNWe3prysNATgCtHf2phf842rXw9RT7aJ/
RHe/o072n1Oi1B1Zzbnz7lbtEbJnwxEFz8Csv1LEasNAqMKiu8m3UnQ9uIe0
ndB5joFC0emuGH/ihvtdz+rG7db3mfcMetnAhWw7XdmYcBYW8RYX4ublMiNc
RMLYzE3rmtIOiXX1Mhv9IK7DzMK3XUP8MTjk4Cc5+63tLetdw4qLGun5y9tv
U3Q88sAX7PJChp4wG4Gq7me8NHir8qp4ULrsWd6cb1vHP3VaLVi91RVbdZBq
LNfgHDZMIpNWeEORNuX3sj8aHKWU0TGDIXg/lWlwtfZh1PWASlrIqVL7VTDE
CpcfFErsfg7R89pifPKeZkGtc2hvCjBLe2Ct0dDWzpvibNLJum2oeZ31oXgY
BFOXI8oKJ5GbvgMVtyC62wxiLNdSlJ5PcSv1yXWHB6GlG3qyHgyD0iU42gWU
u7qw44DOFrnoqQvffvvEQE2WBYtHBCPA0OnQgSuiEOCM0JCyFjnBGkTSnIRq
Jpm6lekhAtDDuvge9mECPhKtqrHWh21haRdgq7LLPBBPyuTZMLO7sNk7Lvo5
fVknebUIRMgqaV5s2MsL0sYnkYYJ0pct/jn0Umzg8SKMQSrdluwwzqjx8rF4
jvmoCL0Fn+BhHYfGzU6shLldm/5bkTC5WvicB4HwH+2pl1WpNinrrJAzCDIc
84+5J5OyQcoB2iqRSkFTrkU+VqeDtBLGZ0Kf05N8dOsAs3lU6l/L/GuH251d
5rU2TXBGJ9DnMCGQ+qcr9qiV2X4I0HwR95ZF4HQ+OVKsA4zZ0rajttUwzoyK
ZoOyPpRHxJY+WyMjo5EN/cYWk8QH8e8xqJCfkNfiBLGacSTEge2X2tDDIdwX
zSo7rFJIpBsQwzJYGLkCPAzysCrYgF2eZVri36vDXCj+/aXVbd2IHKQwfhF7
AcZ7T0Qx/fq1pwN5lqe/3DkJ4QjPuVT+ZkhYN1tF87cJKeBxrD/o0hynTEcl
1K1+vpe7QF1LMDYnqSOMkIdZFQBcKHbI6LGcEkzXmZdVKvZdufvsSvrKotVi
DX4VaanQ0nC0E8iFmQALoPveA6R4eyj6trjaKuGjI1G+VFvhfg1WkkUFPP4u
L0dQeaz5nBBcRE0GWYqVWk/dS1u3WAkVyQBKcSlOVuENygAIbW7wSZKK2UV5
kGV8cEHIG9rEbFhJ5adKU1RUeP9JP+ncEwqjHcD/cezif0uflClvNFFqhp4r
gw/LqTX84uwKV1YQFGIUcPge3WhvD6j8vSBwxceTGsl43oesc2pfWSyV4KDU
MtuU2FZj9eC4Xby3g1PyrKComWd0VwXH5OTB0I+lQRsJil1i1Wv1yllYfC8q
JxuDx/aM+imjxcCAgBC9RU1ltKmvP/r0N7qIG/xVNdMSdTd4qutBrfAdo6pD
UroBBx0aSKsHvLz7qDX4znYNGZ5JqeaPBi6qq00vJn7JffoAqg/E1KMmk6mH
eFBl87/FD7sLEDITEFS5uhbLVyUW4Qpd12vAEJf4VosnIvOz7g//vyBtMOmt
i4ynksRzIwYoQJsENQ0MvcHKBPGgBtOctSDATITMnhQz4odwPBHNQg+RU3h4
TbUojTQsL5bheCZTqccNmYsyrtvuMAdfnpsQh+HnxNDnf9HW8YBtb596oAEK
kF5aQtzURvJ3I3Ikp/IqOQKE1xk6mQoeazhbnmOstsGh/8VUxVaXJYEv1Ad2
D3UOS5WmnyejrM4roNtXhdgsb2oSHnbJff+yzW9n58ApQiAnsDoihW/3HvUT
NovCxiBED56s5K5VLDi4Q+gC38uo4uRuD35d5X2cgasP2vxEIuNh3a1PpgWl
ZtPCPR0hT8jChfejUQUPU+4fgVniqTL16ua5t4ueEFFnSPol9jQIyVX+HoFs
LKzqPeAZcA8phvgJSCPH1ulf+jFWY2iivcIap6xfou6CKE2mRXiom6KGjCf1
kXCM0gkN8d1x8q7oOzzinN23TA24PToBTJjTqxQo2MIGftH/VrM6uISPltcY
wkwOf8yn5KgJvHi9jKq41bgHmaP2tSuWxkrjAeGPEPLsodjFz9X4f/t+sk6z
dn2fxfyBAjAHAw4wiF4/YV4KjmR0Yutzf8DlK0J6MqJxp8RoqFpWNUCWM5qz
T7j5YAPQIRgbpxbC9mbgNHrlutBgfyjTdDw81A0n3iDrC3t/tYADal55o+3Q
TY+UTj0A2++yaG5NuRg0X541fIIHfpat5wPWd3BDnFb2ws6v5m5NU2EBGZJ1
KHO+FPWLk6wNVpcYh3lQuSgFafBNm4eQLdJCArjp0DjtwcI+WNdap5Yeb9o3
uuxLc+D6QhFG1WxPJbfsDHilVyVzPNkcf0Uqj5QE5Y+tBWl8AL7TM9C19qR+
LGVnjgJkqG5FVv0WBup9NSCPFZstzPgwQdbWAENiKr+QbCnVG/PxNjLF/XBk
XNsB0peT4TeRhgp0Gt9P87madN+nZDUvpGrMKpOk81WbHOSw5M60H9ZKyeJC
CarI3WGNRL+NlGhY5HGYmIBfvHO7selyq/1IPxOxHYHEIWsTLdbhrOM6ES0H
rUx0BoKiepgRCBs04KKUXzktwY2MoBzkFLXJ2FtQJc65GJcYjopgw/Jv0NpK
+zu1bZEPHaslooKn09hCUKC1KtnAfkNakAWfXwmcM/Xh0wHLZdn0cgiG7qHz
b42G8jDUcnE/ydzlX3unueUHb77cJvbl62X9+NyJu9Pyn4uuQtAyXf1qnCgK
BAd1az6EqdWCw4s0nB+Lerxs+dwfxOUJLEsBt9cKCiu1XEkiiC1IyhSIbipA
0KayztoZJo8fD83u8VCPdvKd+5GtCviUuQRHzGnrfpULC/WEu/YRcK1QXpur
cJqRv5xE7bI7kGawutdizqcEt24oB+Jke5iij4DeTzWxUIRU2DV3pdZw/jAn
Kmn0BMCQ0VyTlLIT+3lhsDb4eIA+pFXkSJeCVfLFnxC75dG6IILrFT7fyqgm
IL30U6iAbFIbFU9Af0Jwtnfk8CTJUwz/wew4JPtl/jJtofElS9ugmGE1bz5U
m1jHFSw3Fc0NpMCRbXeQZrzfuGtJf8PX2Zhu0pOPBki1kwdT2W1GKAaV5VCb
GxFoLlSxPI8EQEPefv2np8zSPwuD01Va5QblvJDQV891jUcvFSfBlgv0apKd
NsADqiGeaQUTNN6+CiSy0iIl0quc/NlqAixcgcWjhmnpFpCYMKbkGhxPsF0A
5/KCBa8jcAVFvw72t7TT2lXW4r79b0fm0NRWjlBf1EIvO/oS/Wl1n/3uTlp/
Mu4weLXvDIA4lSsXYG9PRYzkUaLVLVECjQYQIKoruzX7dINX8kUpDdIsHmJ6
aAf+K9LrhrDHpxHY6U9b0kMdzSgbZXbajpOfYnJnkTWNlDYMR46QYB6eZ0Kb
N8ZMQEN/o7dRuvBNNvOGwks3eN7JwFYhpsvgad3nx/HmIrGLczKnFE/6kQy3
8j7JqOqar9UpdmXi7a9an6anesjlGEsvAWCTmN2u4bWAvvUcKYPKy/TY4xBk
OLdsocQTe9Fom+UIeHMGtkQ5r9Iehoqhv6kBqfR/5zZedoSugecOEeGc/nCY
xJ6TvW3sTNcIMf0Ri1f5DnqnVWBmyBKrbDMmE9kPbqfaEfPlQzJt8aotUHLz
KjdHh99AwVQyoYDcx83vGwcPbwj/jwrR9M/GYi2LwNG505Kudju5gIM7zuEE
74z6/xGMZtQb3hp9R2TbKxc82QeSzt5euryA8XPKoblGuoBoUzUioJrnebPB
wkw4aowQEQ9iTG8WNwfVCoqCgUesgyZ9rnLSgMDYhLobsytPhuf/fneZ0R+l
tKOqS/Sysr40zkqDidne6rCmeBzlGCX6wTal7Qg/DwQijrjy/eXtW0Rw8oli
P+mXlJIxU5I8km9HCqqNWf9GFTBMavKpUcYOok0PUdptmBgmzv7+lKzU33ON
7rYIRg8Vwd0CbEq+YK3GIudsZtva2lfKnSiYbAjKvoSGkbZHhQlZHjnWze6d
Pnmtu7PNraxYFEh80Tfhbu/hTnempeTV7kPx8tr54U5toAQQUT19ni++KM5t
DA4PxqK26Baqh8u6rwrCkHl3aIKyxp3HJjTl+glJnZzOe302Sy0LuT6NXtAD
KlVuZZ3CyCJGiqVNdJwX0uEStikIcmDw3OcuZKtOKXCPRvUd2HGcEf/8JAHs
uK9G7t699mIUCS5PgtAARBMLQVUCbF3FHuNxbmZh2u3wOMEVM4ws8o/sqOCr
LpfAWxDmyJNj2O52WPmDnq3kHotbsXQlTByLUPE6wWChIVRMXYt/MqC2RAC5
s8ZQ969qMi3Oq5PiaxXH+n24J/tjC3szp2Iag67WNgJZfmcCDKOd7SFIFg82
hL/G03jCwz+Ytrkxxa0s2mu1AwNgnBnNaB+J5nn4/Dp554hPJbnIkw1wTLqp
Y1HKoFYbw8Ybl6D75250GAqK1w3uBPT+dRDQLPitcmc7bqMgULDRldx61pBd
n89kuDeQkRIzwZzcwB3OjkiBcQKZZVTmcRvja7EttUwHZGYhzhjuXqIUBmo+
8yMMaiMZXLinztxtYDC4MH2hgrZcTMquw5w9GORXHBtgaCyxTXa++/g36+8B
yQ0+V8pX/EDnRTpENCCbZi68aJ3S99TQpRNxUiKgCNC5Wkiae9uxkexKP8KE
qGcjnF4jNidvK4CFY1SFkHJ7nzmc8xfjePXXtMLnVBBmCvbXTabgOChSodIv
H1k6OeMQZ8zqhl0AemtbgiUSEQfYXTNFR/nKWEE4zy1OxLeValRTvqFZkARw
Blc5hxbOaAJS/060jEDmyoAAacZUReJVHyArlbULtDImGcr6prPeWQdbtvs1
E4Z4a/fqsyzyD4qHBo6NGrUtreQzKFuD67HROMDB1eAdOOimvha/nyRuFpEt
b+ZXlCqk3OzCzEOQc0Ld2YT+g9Z7dg9Gt8EDKSL/iMGBzXXpFBJrEWMout9l
90huois32Wj6NHzgWB5Mdg3f9MIafCbaN7BEhpMyHXh6krucsMlp6VNEGGed
pC22isOmZpheG+9678Kova4PmoOvb6OpKVlzeYNisjzxfV/xFmoWSg/0R/dQ
wWdf2gNXRRxL1KluGBo/NtyYFtHVeOqZyviP3UYdkyGaHEhrremxGXPPlI5l
ighcaVjHfwQywSYELBN2dXPugc5oU9yxVQ7fFoCkY5mdgObo8REmYQQoWuje
L8fnkvlkMIjmNhgGuhEvPXCXSt6MXN15Gq8skV4FS3liCHST3TggjDPW5aH7
c9CLKMZop2+ono0Nf+xlD8znGm1r80lOItbr7xCeRPdsefK6clmcfKgZMbbc
c2P2ekkGLG8g1GjjlTDRc/ZbM/RK87zk255RzMBNNZDRQ70PIWGvXYNQUrFL
xXaAGBD/oVefovvUVRREPb08+lv2lrwyEAuyR6PwTwfCOPpg1L8ETrnBW1NM
SlMY/eClOzNypN/geXWqbqnRSslh3qfLzoUeATiDqU/k+ru+DJY06b3Iqht+
3mJjsrKCof0AFRtZ1vS/R+o5FkpQY1RWY6fDtypbW/33vAty5DWALEpCG85a
rSZbei4dB1tgdccKD+nL4/BUNm8EOE8cpD+Dgk/oanFjoCVF0FSwQUprDQOq
PPXoMDeutBTE1Pnm6UGGAWejuvUeHN9m/CIbtTeFBj9DnjcavsUreb7gT7fX
FA6fnggNHx9hSBVaXxjTcp2Nci6WFCFv9+vNANDvBaAgpiTzZ2Ov/uJh1Lwh
zHZOg57eKMiKCOmy0GDM7dFrDa6fENfl/JNoNt9dtlNYWvLkCJNwYPnibVVo
mueWjBfcASkZUGpnW/FD0xnmFquS21qFuTjildXAd7VDQHP92oG2JgYAhzvj
SDmOjEbwSlbeX5E11PO4vgSisBLT1bGP/mpLsrCGLD6/GMzsTQlKn3yBm4dd
f08Ww90fhchoAHB6EViGs8opSa/DCRfahZDcZxo1WB8CORvl1phKLdQ6df48
188IU7/nEetLpI+XKymHkiV67CS7F73noZgux/oUoSBC1pzPBGmTqw6cbGPn
pT5Kq5JtJYkVf0iTIkqCW+Zp94OlS4u5K+dhMvE/fBQxRtYxeERx7rItPKvL
//GYniHllmXYieBLjVZTawxgO1WP48LgP/9EKlYAGHBpt40Q1EEWWc0/DWOg
0TGgZ38pm7KmNcsgZwFK8GLgQWtWzuZlpFTf3YtXpFCbpcqEvPO9/vnAFqXi
KH4U8cdAu32AxYLctwcv+JoTp7btc3WnT/8gAuMj9XtsgVZ5jArCw4GrSSJe
xtYXigMEEH8xZgcWckYvKXFGznwnRt2v0mle9HNgq4vhb86/biSJt3ux4axM
VU8GVuJ8YcP9QIvMFWfxl+73x4RYaVEiaVT1VIBNtinFUTP7XIG500yjXZyN
EZcPexNBYfD0XYOUSkByoddyh2Y0pl4JnybdsCYzhBw/njRBXjIZGa79uASG
D3txtDtQVyJ4id+JVZ46o4jQ9NZiKuZiyfeijzoYIrJeD0ZOLaxNEC38Ge7G
K2/n8n8pTPuJKw55hzkZzUI5FlwTDvzs4q5P+w8hzaoKn6n/A31nuElvXgbQ
dBVJl9Gi15hshBeQB9l9HbDUqeMYZCIZtOwW3bIr3g86v3AiVWM2Ef4SCtnQ
4mOTmHjfiUJpWTiY22REB0Lrviq1qIXWsmYwkMJLlkGcM0QLCti7TMZ6QsLy
dDm3OzV6agOLhuGMdvsmILvadrpTzx9jr4y8py0Tf9ZDUOgWCSvvumXXia+n
bpEPpGmnWBAPGxEyvrlUI4lJ3IzBix7l/y9qbWfYqbXETgQ02kT54Ec6LbgP
aWgChvkF88Q85eNp9gNyI2FuWIye8E4J7qgbbTtpi+pzNtiuC9i5hWh8OF4H
PfGDzizqOGFdsNV0DdCjaViUzRavfVVROsPg38neZvVXY6opIJHaGCDWMsDK
lUROmxxyHMlpZGKKt86OChhvfvfO8CYGz3y/kvwn4JlpFjwLpJNBLsbSHt5H
MG24/cqzJzl5MSyHHoYcgA9g7SjKVY9fljYCcAS8GSvfF/iOpnySEE6WMJjg
yg4dhBmjpDDGw8FjSmDA1KUq8YL7xEHfR3+l2sAD3GnGqtNsIdGKsB0u6pdv
YXwgefvnN2dTGDuC72XcnPVA/WjXfUu0phyjLTV1cXuyiI54FQVVHtOJtuEi
EFtAA3vtAqc3IAtbWuNtrTOlT/2LyPTHCtqa43m01NUmQStfbGKaJndYYDmb
wBVlhDmO9UXgrRq70NccPTJHcmIvu4WrzWO2lq0I5czYux0ks7/pJUfCbVS1
RNtJk7Bl+4xQQhj0CoSJK4zimZ32wUVoAUZNR9PaST8BymEu8qikiUlRGR2A
bmI3FIZ99bMtAoJ7fS/bbYpdmlN1y8tKFOC013tDoqZwe9LDe3D4/0Mubglj
8JaPqeIZQxIu2hRnAWIbgiej158dezaZyqV4XB3bnj0KvUyxiWPx6Qw46yd4
AxEqSRIu/0PqqMyLxT28BO88zwaOx4xDB5B+H74MrVyroxmVQC8TRLmVntk8
7D7zP4yKj6b22cMWCCj2VvJEDAODqThOAk0yUJSTyzQLC3bHs6XpUDqvtRHV
bPV1AeTHXwrJ+Y6aLDWoDQ6R5GbgJv6xQThYhzMEFADqvQZgyyCTFggfpKo3
m6s15DPFRJLKsulpYamAojo53S0mOyiJEMujZJfhPlx9Kh17CMXieiTcEm+h
IW49WuXdH2rby60zxEHbrqJkbZb4xPeLIypUTRH/fIBr0sgAqd4KO98C9oZY
FhMVvWKdiVThlL95aMtq4fQnQK/o74t99ExNpyT0VKr3/K+uCpYWRXnpaNn3
wN0OifuJj+zlS3VoCT4imPMAnSTG772ttb/aaWS/B1jmYyK+erl58dLZj7DJ
C9ofOboJn1GI9tmR+5KML6JAo/V5A5IQptb3I30jtK4zew7JWBMSpMhsEb6z
zPkfPemyBcW9/8LB9yfUJnDoXmkDMvga2DJDQLdqS7Dp+f3o+XMNwBK2t5m2
v0avFBVB4Lw4kRWMAHMcbzmX6W/9Q7Q8dvsaoIm5iZ1YZ/7fu7pPcyN8CQ0e
yUyMu/asN18+L4nwDXY7cTjbAvlqXLHUWoArTcJoqo9mDTmk3dNvaNN5q6ix
C0cHESbtKJ3bQ0ZDk9tG12NIwNQeOluBkzvlYC8Mje7xVRIqEVyOhPN8cGDG
6wvEuU2yKl2CCnogwVxVn9X4YGbClQMMVW8A63qNqsM+7IFkQC27bFGvTCLX
WtU81gG+qW9OCTO8bKhFoikw+PTW8vhwaoAoHtmZ4QOvr9NZE58vyh4fdwcp
gGqrNubH5gk3oCZcZGBVrc0L+hrwu83cnlcRg+E3mGyM+VXB9Do7CyovHDNU
AzSII9PiT3ZGatjOLHcREOVkG9x0/5xjUhoiKRltP85axFiO/b8RBUoHbis+
w2Yz3osq1+rxaRKjEWWJiPqXPkVm5jg97LNp+XB7ejRfUoFucCgrWeUE76Fk
K2DdtO+Fz3DfaS1z1OKnh97uXJtreRqUKVN0U0HnZXrRBJpk8oDaD4fwGTSV
+OOkafpGWxW8pQ5+yMsB8xnLGKSESizPU8QIEhWjhmhxU5uKR7EWhSzPCaF5
xD5YZpKjnhlYf5rG/HUekLzE61BNBa2ivWouVrW7XVxJeuN6xT//k3fhbVXf
EG9IsFr3VECPZr28v4wKvpe892NVeU36guTITPnEMyoMnclvu42I/wfFjy8M
cTxr8r0cv8xM/XxRJ6wAEX43LTho+FNJXMjKhMRFro3PaMV9dRuBQwHhj5FE
pJY80sMQ1xpQm4hBQVqkS26eOSN/Ow0fFcHWNiBpQFAK2FU39yJaZNn1IrML
7AwfG0DqXjsON6fKbu/aR/q1QXYxgJ1DOlbM6pKFuUB8nWfaIL/1jEOY0pLm
pC+EGh2q0GGdjdAK95frsvtv5vls2Ludvtx87kHSWsI6lOzaOLH9Be4g+h7Q
kLcyqPCX3JVK9Vm8LHWcKP6kAHI0aFC/WAWJdvar4Mmto/LUpX7I78Xo0HoM
ktBQ5HO0tNyAeHY+UiRHtArCt1+rFHzQ6PZqKB2H6T4tMMGLGQ2QGiI6F4HK
jt5E2D64OhbvmpJM2R1bvOmGxuKziunZq+FZU4NorK4TfCoxI5z0iZozOlTy
jAT8PxxskkiwAhnxTYjTUftwOFaQRRgWy8H3n6wNoiyaAMSBP04Y0OTgXN79
dwaSqqC3ZigHVBWqkvq7DoCkHbiCTmQrDbSTKuHie0xRjnQK4ZIOZNV1cBzM
WUSlIpBEhN9GKrfq+XpK3JcgH/qfj1r6GRrJPSsGVNpoRBy2oclxI7sD+t4e
9YnBZiFme61jgipCSsiQCDjEdLo7wVtCiM4TCk2yd5EmeJoF8cs5LXrUCL+A
1v0MoL8jjLxpmZpxHkvtKiU+TS76nbj7vpSZT7gFAby5ZzxlWDu87GQH6Nnu
AttxD+WeVbbunGMusgGZUnQ+ZfSYRG6LjzPBlJXBmfVn5zHUglUB7SQ94y+q
RhNrKihH3bEHujUQGsrD32NkuBBnKhz2jXpkKxSnxLk6gK1ZXWqvUPAAQ54Z
A++sxu2lSaYiFlqvp/BTqx4bExrgVjb0oyj86K78PQ562rn5Me/1IPuf4PJL
9yZlFVPYj6vv45/rfTwb5WCzoTU4Iw6HWy5OjujVZM2vpO4PdeUtcisWlU8S
wOVHCELVuAu41csN8CAqk5tHU3ukP52Ne2DEWUPPmPYgw5E5pbhkqyhkEWZF
k3XJmQJLkl1RXw1Hz9u4VK36Uul4pKDdBI4jc68qHw/Io8hu5mQtsMVVW2yb
JAgLXlwp14AjPQ3EJPPrFHb9dX1DbpDn0nG5HXW8hCj3t+FH46wLkT4v/jLL
KQdVThmaE+51vimqZyIOo2Nexg/f/wpKhswOvqzxRh+8h0kwNe2/POw3/6de
Vt5utEV7XqiPs/4rSCACb32GvRm6e5DmRfQx367sZhrFHIrkDYmXdBTTBK/W
KW4QUYPG/YMbNjmZuIw9hWi7uAjKkiMc2usx5oFGmXhw418eILk9UdPx6keV
zO+4wS0nk3SKsrWCyezJTYhtaM7zdWygeTTpZ9VhrqYLe+SIK7VpyCtMai7J
HyDejSGtHMaJRNgtwx3Ruv81+M1bC2RZoCRHDzkPTQ7TE2vrg5Ux5aVmOy9h
VzKbGyeKdFuc6p0qsBmpj7ItV9PzvyQFhgQhaIMFQwdanAa8g5GAfDCNXsZJ
TrG3Vzl7ifD1sGDriyZH6iCfF1osB2s5fsOiFdWzjPQCnlx7EytWdv1tssRY
jtdwLHgmPkMy0g/gEwcNAz2ZasX2jZvmkUvNY5VQWY7yMsAV/EEn2pChJW2R
1p9G1rJ8iFrllnJVv77UvD8FJbtxI0M7FzYJr9xdcWcaFuJGU9rhONiWPiml
rXIxUPe8fvRt8vVBFLejw7j77oHZJ1ocQsvYNLGk7FN0ggpRsPipTIBXvNuX
hqWwCgbHfudNAoCtQePUytHmf94hsTXpfAgVPcFDn0V5Ls4+k6y0st14FuEX
AYZHJ7k4jpK0ebuZy7I1F5BoxH4FQJWxr84bZk3JicxfmCmFL7yXsdAh6rWu
MVRqHNxYhucXGiPiTWBHCVdOporV57X5R7hCpmen98Qie7jHSDhCqL/IRuv8
B7CDiP/ynmVQn1EuupPUnvlAOmSvc1ZZKhhgen5nUz9t0sDzTIVhPMDCtfMF
/2T4cRFcfygmW5Imj+HdQ1bOQyLtBIAQVQL89A2LGVjNQkyh3yw9OcCTtbnU
GHtnB8aS4pvO9hKfxlH4Blvcu1QZGs7AEY4VShHOtIN8mYHJlVHsj3nn/N2o
JLEsy6akbs6vNCCwSY+/sjKrh7QKjVQqqrk6P8Rs1dLQ/vMbOtKX/LrWA8HI
PmZJxt7fbqD6HJE5oqdpZ0njlx4IphP67vjI/nhrjCfcO0pdEUzyXzeOfJkV
lUPSU9dZ0TqrANttB9t7DFzj1oQ0SMnOHRi0W1Dh9EzzJMOrINXaEISSw1AL
0UbbyEbiAR/i4uMA53lJWuC3SJYiN0ThSInXPEHUH9+DV9Z7/qbHfrLmqA2c
Egv8NeGJeSAccwy5bw1mhiNuXyeNy5qvbUNl3yfznftjmlDxZZgLfsm2QVVB
p5sgI/TSV9uMZUAvX4i12DQkGmyC53tr+kMDTvrunU4YNuWJq3k1VqQk2PK0
9xGQZFupETPB9sohM9Vmd1jPotPbGnqFGDAk5DuFZHXxch/iuaVnrMfnWfRr
CVUL07mTmSutWWqgAxdKSSQKggDHDz24P27UqGnTRgnt3SynWo5GU/mT6j96
0kHRjOia/fv6A/Ool5DmeQzI8Ht+jnaT2IVmL03DC3Et17sO1IX+ZQqL0RaD
JXybLsQ9sTNNX/RDRQbTWJizGioQGvLz9bMsh4kq9Shtl4wMz6FZMCtIj9Up
+cF/PKyYVnyn/DPZukfpvuzsjzmXA1VwZZU+MdMkYApDLqYF4+ONtTWsxJaD
qYugrPKjr+XSSjvYo+L5Mdkn5djaE/YlU4maVzcPnN0SotVLU3ZQr5qM/Dg8
R9sJNegXaxu/qP1wQ2Yk7JHuIVQOjBm77bnZCXiV/J4N26eC+jO6SZkd2k0y
ue0yKMDNd5TtCDvrCMgtbIn+nXdmBoVzrtRIO9n2VbzdXGQBLIMRJZiK8U1B
iPBGjTP0WI/zPlgt8KKO9otiIsLDsXQ/ILJdAufXCfb/jAXd1jq6LLGQ+Nyy
Ynjil1npUaHOjaanhwmCcP8SlA6pADcx1GcoZ6f0JFvHfmJ6pxTzaRd9Mpkv
Z8PuY4SCYez8/JEeFnh4kzcdLtGeahy5z+CEvB5RwCixM9uwdcDHcbBYQZqb
F7/79S2qIIjUDKuRv/Lv6xxxbpaCzEp3N3IBcctdIudUa+SFCd5ibsqZpAwt
EGG+LshtBCxfJn1A5f3IB02HCeI67KtSVH2VRWqeRshhGDic6kR2gopUioUQ
U/VzVikh6UmjMmJlxIj6tIxLqoxrzvhdgTDZWBEBdTcr+3gF3Vr+T1INzv7z
h/UQXhNgepECAVVK4x6FxQoYM7UN+k0u2FeTU8lro0F7Afhvsz3UOpwf7y/F
qFYFj59p2njsLCJt2ofIW4dhZB59eaSTunD4t0R4OPmjRB5hLtQeeq66oCww
2Y4oVrXMg4TFpUcK3/1UAclcRLBorgotDVkNQguV+tAb91uefE2JaKZJidE+
NTcSVJq0SKiySgszfZqjDL7FJanQZhJ/3MfjR+CBRUL4JcdHeRjxV7nCPLKt
h6mnmlJ02ZNWg+OctHEBeqmhZXotluEyNxADGVdT6kxl3TylUgylbhhhbToB
vcTTGn0edZnwackL6xOGBizb6UmGdupWRchxEzWgvL06UWjpKCv8ALAoWSNO
3WAuwGaahnXZbSaYmCwZEIMf5yiKz44W0q7PKt2ozrJIA4qtKdlTD2KGg9Gf
iJnsHNRAQUAtSCEsZkLSzL2DSDhGgfR5su0si9VtE1aD0YpUznBCGf2Bgpbn
FLvMEbCFATumnfLGbH71kWI+I5SeJXfwXVbGUYDj5OUhffm6XZIl94vxnU9T
eBCkK4iWmbjUuX0o49aiZU7miSbbdf+yDMJ29jebc6IkiJCrwXvjJIuDDx/2
F9DS9ubxw7x9fTitXDzIjb1nJQoBe9Ykhy3N237aSLYgPcMezKQ1SVZEj7+X
EXSiSOesBRcMGszqh7HAr8Rec3HC5hkm6cxLX89xiBBu7qSkonYSFjYN5S5k
310n4D45v6N7gh9/NmZoluF/CkJtWM6ZqgrTgP0klO7IZ/Q4rrDPvCOkGAnd
60QFZHPDI9fzWxACtb2zLzbMhxW/kGIruT47fxgYVNyNEKS6MBf8W16gfgMN
3FPReqkuwFNNUOBfq/BnbaTBsoAK9k8DY7sQ/zucj3OHUOmPw1zKoPP+VWMF
pixFfQclPFQA6j7GKsMFJgzvLfJUdxwRO0tj8Xnk7mvpmYnkBJbwSJUMkVFL
TqitXGFDKWeIlCQcZkuBWLCtY82kxKb3DClzyeGmOoteOm075aeJeW5UNodI
Z4rBnUjNknVMoIsOwaNQFrILOsyM62VqWzqoHBf07IYG8jsvXbuSU7dzIqYF
jpWf/jKETr/iONN6NsBqTzl1qIP3DSi/sK7DEEZnTnPTivteH+dV7B4DhWk0
eoIcLjR8rlR0330RxQe4v0f9mqQhXc7egFDjOyR+1tkb7yGgxzngSlCCMXZt
uu4A8RVJurW0X1W+pO2oPYUyEB5bxm2VaIFCPP5rVzXF9CqptJqq4usX+vtR
XWHVKWEhpyoXzx3VhrhdiPMS3zegXqElTnvHwO2WG0pOoVsSobptxKLRU6tn
RTcczh6ItRd6EopxL/LxDRksD2XjXA3tkp4riVuyxJMAbyPci2qET0R+l7VM
SI8zwhrOQgmP7ifGWVL1bcotR05fWJl30Tl9STPon/AwhZ80+iPVzCeGvy0z
ocHGOC1A18FYMJ91RCPukoy4Ugm4hITcN8v2BL9mu2+w+wov6xQ2g0kXchH2
fjyvheJvXugri3dHdB2A4+oFupG/fMjZwis/4h5CeNzjIc3G95GC3772BjsY
adzFNA/eQXCw1TcZKFn0H6sa7C9pZh8t4uWMJRWdqoZXRmFRV0BCvoWBV249
Lmu3zHVkfz0tTdqX5ElyeEo0d+cVXgxL3389E56pDfGeLJK4dqRF0Iannh/m
mWClq290sh00dXCO5t/OLrO1bU9G/OAtatp6XtH1CdkcfhzSu4bOY9Va0484
N6jfv04iOwRyp77fIQB5Yy8oTOLzNtvyq0ustSGQCVNpfqK3UHb7P0uu6hIN
2KhUVAtqCiXTr9DOPKoZ7c6MgqVa3egAQaLrSinOZraXVDfgZbPh5m7K/bs9
WX9i5Imd1r0KWUcvaCDGRlkMaDhgZbXPTzUtq9sVcBu0P8shJnYnsVCEBSLu
ZD+JRLk5UrPrdAijR2Y1bWT7JEvHmKt2msV6Q9rtb3yyUndpHN8zzFsZT+bv
qstcXRam6Os0kre45ZmLRf3g5YCV7/9CRoQ+CTfadjG7cLKqSbd0V76Ffnaw
STjBwWKPai1kGjmLSdWs3kPwnh7h+Ynp6RbHbL5ZnlTQS3GgtPxDVSADAS1C
v3VHs46cv6n1Ddh5LF9j8wrlPL+Ot1GmPT8qyS5dLCHzcV8sPr4uOZAuWvOH
+J/RpYuQma7YKqYWmE/yKrnd5E70lrom7uBfhV6A47zgquFM1roqR2swZoll
GHxlQT9t0rzLLypueWQhHGAEI3+rZeu2w6jJc2KNkIUoJQUFF6A3djlRGEom
ZYc84QI1SiO3Y7beRUace86Xpq+0lTR4KKEpGEU+FvrnVo+wvVI664Q8onth
0zfPa3segzJ9jIZLiXMOPckT0UVhJNu+XqtBXV34oACIgTkvTAKUvKDVPwR1
NqyHH4HfeldYw0kHGwdfFHxePQskHZSNTOt6hdhzsqwFcT3dMe/IOkQZOimb
/Ef83PNkOGR8j1oSYwjiNE2xrJtRCD8ePFAppWRPEhuGTBO/qPW0KaeENos2
VaXoIQxB8KEzDciPY0zKpUzLqR96Iz0FUHhaeJAxvBKNgR1eheGpoJt8MehD
d/U2YG4sl2lsjpYCj0NH5OlfqVYkbJ4S/I2824N1F8F6ySio9ApwKFS/lAUP
BVubng/5m6Qil5XdSqfjycbr6g/q59KYBZUil+lWE0ZGafrjj0xX4lIrv8uf
4WA7T9RbUtiga7+jvUB0Hhm3PN1NTnIxlXy1aazyvdLvv4fDgACx7Siy/qaG
aI/LNLPkI1FxfEvbryoHH+00ACc566Ztdv8tES/Jk0ao49xEleOiVb5o1/TR
Uc1IIRIG1DIF4Sj/Tyo8IsJ7GNIYOyutazO36qNageIUvRN1WvbM0oEvc1eO
FZ9P1rRZNqS9MKWJ1pEQXNE4RaLhoHMRIbOdDWlvueBIeSGDxQAIGLlXiqaU
uFkYR1FpxPO3xuo0dLCBPzculTAR49n9EQqQMiOnfW/ijad0cbpa8HRCxNY4
5tlLLj5U+QWMlTWG1FGaaKl5MpDfCDYuDX6QMzIt5V5Dmsz1F6+S0u7tR5lB
5YHj9WXvokIVxPd+q9HhioOOz+foW5tQBbqLD2zjBr76Q7xkFCPmYzlh0Amv
SVRO09IegSF2OjAv9BjYaUB6ppTxxmU2Y77Azbw4YbRmkhMkUxkMNfM8kE1Y
fKh6rrS87OIOZiiVebFNcumRwkodGQ8YuCLIenErW5X2z/XGQr4xMdvpPG5c
SqrEoMfCv0J/e2yQkNDVGOITdfZWFuVj6fJkwAkotUgkQFujfrqS2d4nv6OL
cQb+YC+liosOeKGVX5l11lkSkbrmA6LUvahS4Rvq8wLB1XPOZ02ft5n+GtIc
IuGod3vWkUqGD00IVgFYq3fev3aNWUznuF+gXOzlz/ztOZuE81mIzrL2KhVi
tQwAmvKD1kOjDoGTfcG1Y0vPezNKg5Bd6IK45hsze0HTCFnr0c6lU/xAOxZq
kXPMILycwG4ObVvQzkla0/XqAm1/tg6glGevT7ZJtOAtXtOTYfcUkkrA+glJ
3XjtbkSfW8LeyIzPV65lFuvSCKmzh+T6+yGoKar8AdASI4jpcxU4o7LfLbBe
DojEkOwUxxHBvLKKbyAxXix/5++z+T3XEcaTz/dgp7A0RI4jCXiHXTzrPF1M
kf0w32FZWu6XRhbAZH6Cup9pepzBbrQrsERSMWMpNcLXEV0Bw0QMDWb1XfLi
bkgcYn/bOQpcO2UrQEl/K1IZa0GMkyZenyOY7u1WVvdttrub/0WtCLNLcDln
w3O+S1kQp13E839qD6UgQF3ZEjJBAJScpzuNSImTDBXFfPPsfpfQs8735R/s
VUSgUZLYd8LrD+XNonfsW8ZVPx9DZu6JcdlzLzKvUKhzSVnHNLlNon35I26L
9g6IcESU2pj+mQVNEIZR/3boqIVcZMJhjdg8woqOvWx3scv87v5Gplkje5Z6
80YslIGVijKFlKiFxbsYRWkf5isRBqmwtC/vEe+EurfAjALvN4hr53e3T4nZ
Ozn2cU5mgPlfch9UfanqLGnGrvBoslE7PNlnadXgQBsNr6dnlZ/q2J8MYOQz
fUxE01sBd8g5iyvOhwelWfysI2lluaOWX1lqvk7WLGvqJkVbOHPlAkTg6Kxh
SsP3PNlkHs5cG6HL0BOrp8onl6wR1JgrSpn0/jczBOOknp5sEvyWO1PFWWOm
T9g2B66AeZjuEcwkmYFwrjZERonKVvoClHodzWO6HyFWsKmjdfYpCPhBu13n
BQdIplNV7UdFoSzM/v/0YTuQu5AOWAx0A/81KJhl6Cmf5nNqdulDC2uHjsRd
3nehH/iIcMiaVzW2I+BJsy8XTWP9V5cu/lqJKZ3WbTd8fyDCcs+8JidP9wg3
7rCZLn/xDJy2rjMHq3YzlbRnHxtD+/hGyHSLF4SbJil10XeAQhjNPMlAMcze
ee0NNmVvdpoiH5uS66gPKZsW0iFwClALOZo02NkN6k9A28nUAECM0TtQGb7a
F6B4gsnSOk6sx5NunwzdD7pI8bNTUo0lCiQB4mkkHgAY3kqh+9OrJT7lBjeZ
9Ffc6WQ1bNEtJDY5xzHuGKKzHbPBpp548unnIcfu7a4pWNHmIIvs57m0netw
SuXUAxU5zG3IKrd2N/dugTB0mNRpYYK/JuJWm5DQVVgU9ZS0mqUrIJq0c27S
WkcRZOxK2CGBBTE9sPS/nsJMZctV2nTGDGTm/VYAlAyL/IcPG/+DiYj5Hpvj
6+z5tM2ZKVo5QFEEbpYuSeUr1BuzNU7G8LwmS4aboAsPcRWJKr+ITqeuGOzx
47u7iAoP1bhpb9GFw6uthA74IERbQIRiAb2ZtaewGcQ+1IBpd2jCc9WDMWHo
wXx0I1g+rphGcrCoZpt34v2wdYOfHK/YR3FMvSX0ljOTmL3ybnAPQeGmhTrq
tfYyAkUm7Q32RrUpF5jnp2gAyUKfEfK73gqDe7Vp9eClRdceTPXPGBvEsz1N
V2eGcBKybgbji1rBoUJEYjIOL5lqTgt8iibS7qC6IGdmJsHa42RrS5eq9viN
q7F6gV5U5zIi+CFgaGitbGyFU1iCu8ucHr7nqhdNv9WxxnktuNhxYYTj+UCo
9DkluBEbLUZDtdm13v7hbFWpyFzr5jikeKp2pwNdqaYciBoPElN6iUb7nVfB
FQyFBEfzWfCCOk3qM7kAjXeHcZzKD87IReHpMw756LX+Pqf8G+IXeH6d/cz6
wDfAxLt981hGrFDZUdKeer8LWo5yY1oxHghSyL2JWKnLD+3YWyOGfEQ2PfOr
FrhCa2ijR5HsGGUnAZuRu19FsBkB3up14vVGCXeao5UCq3MKGQu6HO4KclR8
5Ow8w/TzkAsBLP64QBYPQfZDR/5sBNESKtuPqEfKkbS62U0s3/vY6PnocuCr
sMmgjqH53QoY4bxW/ozXXTyT2W9jZh2b1KqDpdaacWI1/+VhT1Izn0OHb/xZ
+psXDqcwE2dYHv/lIwp4V+p66i83bk6dXmgtfA7p0calgRx4kfD8+n9EoEDT
nE6pT9PMuGH+IOtngEGQ0ojKDL/na2hwUXP2LSjTaU/9gvn8ajFOTSUFBRfG
4S/j//hMeKisnHOMahAqvSOC0H3Hb6xEOgy/XBiokZpMYUPRR1FpQVChuAeG
ZwqqeldldSNBaUQFb5a8AGkS/yCN3NHKY9hkl2v0v/a2KwiWapqat+GHqsaY
Qw6Sj+BuRNEnnxTSaA7Q5mHip099aasvKitfNOkRL3lq7AXeF8TGAbdN5WIR
6Wi78KKKnxSkx+8yKj3ap06gQu3bMnSNOOmYo33pvbfLegXo+UgKzJ2025tV
W0UQJLf6Ap6xw3vsthcYlhn2rt25oFmoOBHdE9AQAiUkeEGIbmGHv5zNaCft
P4yXjdXy/flawuqtViP4+QF7oclIu+GZ9zRBkbVeaTfgVcOF1S3lWYDWK5FI
FrPbhDi8zCOlEFNtnto/rajaudfL9Vbw2/SWioFaL6vOKZLO5erN3D4NB5xW
hRQA5RyJf8snPgvyz9nLMx2M4/Wajyo0uqz+M8NjIEFoCobNUISZ3N05XWrB
G+yJyivNZFKTXtZT2FUL/QalvcarAaTj6pKb32ixd8XYWqLdisyeDBt4B/Wc
/aZTI+m2/LWsphy0A/C6Er84oi6CcjsLzMyU91oE00EZnTr1AL7FOZNrG3bR
p+v/8krG7NM8fuYotGH7Jkn7kCJd8McqEfxHUxBP3vzgEoUYcHpVPx9FH0ly
HN/eggT0VBp5bcFKpWOPANiJLBciPouQhabNSzWFw1Op7nJo+eeHQBirXQxM
LiCUyO6LH0c3u9iQRKB7MU0AtDGb0oJpZkcezJTgGBWtwOBVnjUD+HggaK+y
A6a1kCnhuRw1slagWGhMjr5lLBTwm44zGIaVy0LPY5oe3gUpGvQcDc2fq+P0
GjERI+U7Bk335j2w67q/ibkMWAjFKGZYcKgtSL0tnblSiS7klN7rSbniUFOB
1ZHf3fsp8bujSyMpeuAfJpE03/Lz0M2fMch0wTRQTU6VqyrKjgLHPmpM2+0X
gTkHpziwzt+CFXrVEckVPLYd0UpsePNrKAK50MYzFefZ0P8MCnm3Fo69LVTw
xr3Y9FLquPI7nKvsDS76FjYjQhbUX2blq94E2caWjRu2lH08OjBdckudObOj
ZQgAo8aEoGkbrHoVpjnfd+n/dCIEVQjWZpPgT+yi9YVMPlTShFsRW0j+3F/k
Sp+fP572Jzp+F1bowcEYL5cITTGkJ7G5XktX8y7qClesu7GdQ4nSNLM/eosG
T0Y0SUw528bDKZAe38xpzfSLtzeu+CK2HAfeHKQyHGQ58a3fXgRVmjIVl/hH
lGAJLGcICtD00ptLJjVOSD1xI8RW7IzeS1bZcRjXoIxz/OrT84c07UQHYqwD
1Hg+aijzBNSSu/gMrF9wjR5ooApO7KI44J5l4VtCeWdK49zizFIELMwI38zV
hL51lo9vUePMAAM+18/TKIUfQ5rPTAIaG1C55ePBl+IimhKiHpdwhWMKICjn
j/YiG6j7idVTaqGGBJ8vmOL4Ct0GZZAvl1elAOjYifSqjo5hIMW5igMWiRMJ
cPMz3yXdRqdZk8hyGrMx0GxfGXFpLS8ynRiW0egMsaU0t5N9gT6c+BIgk2xa
LcmX09vsiEEi4mIqyUzKRjvIxZ2WTadDkihnc0xsCb1jwjfgijkwr2Gzaxyr
DtvGD0v+N1Fj8Nu4jaiuUB46FSbHIgWnOlj/Srv4zI3MDtBoTQEZVBJVlJ3H
UiOHBNNAbfYyJRxk2/QWYhovZhY2nnfhO0OjAf2RCGZlZ4l3AQ4GJN9SsFXN
Yvllf9/bcRXKJ6PXJXND6SwMBQ5sjjgL3tCPM+OEDECA2doKL3xpaJvOHQ2L
7wdNorOTON0zeqgETsTFcT6k2Qwv47S73x4n/2hkyvcWe+/qMsS1+XTmFeKd
w1BV01Ledskf+LNahxWrcUXirHWxSFKElwwkUWqOa8sHnNM+phQEOxMwWpkI
d4pDjSGDcGW7Hl2icJUt+oW/79mF14GoSlJ4GppfUzWQrD8kqiwTujVCczF1
spGTxwjTCWalCeAyCzIOujvte5LxOIUHddYRzEjPceXdBJCp7ga9cNrm4ZXs
2A46isNIt70Ywvin8k9cS/3Bo3gPnpDUth3kIWrhxJeyUbPmH1dTf4VKbrYR
YXuKbKKFY6jq5KHUuuOPRgIVFrzO2/8hbufVnrGxnP+zE9A3SIvmxNzw/UGJ
fiqAic16Z1sLDEGPuJGxZTdpuDaD21TheIemtLwEIC6QIJ6XNmhmHufARrdC
7sUS84oRzfCvSAThlzsXQ/Sh85avBSzLP7vQJIOzkEbZ+rnmrqJFOICMGWbM
DEXfFZnN5Y9TDSJLMvFmU5xOkJDzNad00ZqkDU5878APEfmh7lCZM5Q9Dxj5
+STR8pFIsL2p9mA2tEwDqJ5sn/KNukGs5PlpG8jkNgKtsnN+N0JPOhESUdW2
IRVS7DXeep/xOqSbSBSwJxXGMg0hGJxuKp6JrWcVUOGUww/OYig0jYaqS+v3
nsYAmpNtn6Wyg8cpmaciiMV5KYbCLGZkQLq0D4ud3zuvmQAb/3sLs0Os5myS
2CLE5DRB/pjmFsxkhP80ULQZbxKBi4stgHnDacNxPJhIBX1ge0CwrHal0Dkw
b2/aPyTznsheMKU++zous1MsJGBFIpU5xhOUjuqKBK8g8aBqXce8e0VFa1x2
mrnRG/Qy/YbXCQWNfrheIPsPgn7n/wXvf3M6f9x6f2qUXE9/KbL7RmjEVwj9
oEu/md1h1LwXjaEQ53iQumsrQeOCIVqsO/ZZ3jL2G3laHL6uyUA83fYZPGsR
3TdNMetr+PxsW0ZBNBbz6VY42zb1cdz3OH3EaM6Mi0xgyjz/YvLEOwVvZRpX
dF5T2P42cApQDOOJXM24NrHuSmCP5TlQCyDIqU+NK6RbCIY4F/onokxGsYa2
P2ToZ+Dvjjpwycf9ONtqlOt8dTYuaLYwieE0NVPXG/69q4ilo5yTtlJBRAx0
TFLoMI8/x0ycRmEHYVh8p2V8zPPanZnsrpQ1A5SPB9+p/xCa963qay4q3QAS
36WQeekqHrNFcgcfCG3tcSghOJhLhsDkcHv1+DnYLCfmf7kBhluodl3rxywj
qWzLMHskDYhMKozj5/aAp67CWCTjKQ8Cb7FmepRnT0YmdfTXvSK6cbQA8euD
8ZYgmfysaXrzxpBJrgwOiAWVl7LOM+qz0uhWRI2/6Nq9fDSCPV58tLaiDfBp
1880eGcRbObUAMqalT3uJ/g4OWxBaoX6QaMTBQZvXE8TmeeGTwIfsI40FsCV
V0z3sTG5bocX43orZzbxO9+3ZDPsfADVGZgKF148mqzuD+8DZD+rk7xV8384
PlWSAGGquWY8TPPQBwD5y18Otjb3rnd5t3qtYyJLmWkumfpTwvPD+cRTG3nn
pv4DewVj5hI/c55xymlKZaOyVCM3t8ww7tIXjQVswSYR+lX30OjIHhxHiXVp
SKabE7DDFkgMIurORTLbXIN5iy4kiDXBJwJIurc4n1Mu8tkcPMKejkL9+hgt
17wEmV+qE4vVvAoKZ13w+XSBTlJ3T6MwcHoWmR9v6mDZMOIPqwvNOFJh3wuB
nEkumA7AarPU6jwBSPLXwMvxg+Lge8pTqC32TA7D2uLyDy9r1JICQIuy+ghp
0s5OtxPGmh1wka/an3gTA7IVbHNgVsEzlpqvyoKM11+q8S/lSAELVnyAryP3
sDExurdTn574P8xzSXxbrgfPbRS3yC5ladjUmzFlSMa77W2CoKroKLqTvCIb
7QKgTNzaNAD6Z2fi0zO1SXZEZIuOzy6b5BiJmLV9mH1YDAjqodtlRDJo+Aek
nrdXbZstmUEtSylUX4XN4Lb5T0sP+rOuPfiV5oyIwNc3S1gsV/1sJ8Vu3lbZ
6PeDNkX/UccvKI1TVmdDrdUGFVyTxgeB9zDssTwrtXbp09+G3d3h8miI7LsJ
kFxJ1fNdN9SxN6MMpLwP/MHVQulb2Oo0mICKtmw8PM3lbGtAMr+29oLVdOvG
FWdwRNKx4eCZqk4s4vIq6ZUn9UYywGOqrYOousuyih8+LH1tEGtqQLzZuDcH
i6Pdd0YYeEgBZTu8vcv0mw50p4uMYBQBpYqITmo+33SuC3NlJxiOCdvR89yg
M5avRmSwKQEduyXbwb5iNd3Dl2mqtg3d0hpXP9Xyh//MPKXUm2EZ3D1EvSRJ
g759Jq+qCJDK44mp6/RYpBC2p9tJMvzq9rO+6NQ4yZcQUp1Oy7zSuXscrTP2
TBILXr3L8hIkH4Mpiko8eQ/f3gl8VusVCyQO7A4cOrKl5mTDcMDjCdGvfVBJ
e6lP8H7JEFpbqfABm0hUJSArC4+K489WNQyE8PTFEVVvJS1ndVOLm/pdLUjJ
7tNVOxBHvdmV1GJZ3uawjXjHx9yuKYK70sdTNUs2IR+BrBFqvxtL8h1HVuR7
pF9OZSpxD7Zo6Cdd/px7UK0ogdwdFBD1grWPkJiCIsXYGzPTAQRV8YvfNZSN
uBFpap4HeZroMcGP6cjxTxBUCsw+UK5bYdytrAVunYEE27FqugNA5jfkKQ4J
tBYSd/3oHGBezua2xaYK+qBMbWZu3VEJzYnOp8CtE7ToMrdi45ZgXHOuXixP
bBHTeHsegnhca8DrmwaEWu6aI11ObBcgMBHegY7v0Jh7F8BzZqocnmThYkmF
wPY3Ifdyy2QQaBUUI5WSau5kF6ziWcAVPEEWp1kWp3Zw4D2gr+/AB7nkT53S
JONx5IsbzBtnBRLl9A7dATgJcroZeWP8AKhkqQUILAv2QTYrb44IcLD/kCnd
Hh1x1esOqTTiRHWDDtqcyYOLJdzGz7ha7vUEsVhpPOH4lWWVtG/ZB6buyl93
Tlq/wPvDlU+lg3R6F3bzYxnVV6qM7ytSpSRb0K88pSIK+XETmuVvaLQvFqfr
tvIGVhCUrjCVPBrO6Bbjj4B2/icrcc4QQ+4WSg5OXHxjIyswkObsNOkZr7Ji
vHuiMgJCBAk3wKOUEPN+UKtAsvfx8ItF9zaNfO95hHLhxpAge2jPgpQnVn7t
w6mJ4LwSrn+gAjPpz71s9cfdbvHlSWR1ElL6MlU5BYcvzSKDgL/pzdL6u61x
4TLFu/nRyM0YVaR7UGaDK6N4ppGoldDbZyXjwvksS6Z5UjPCGXW4k+qBZJIi
6SY/H9DJkoHGTv1V/UI6KQ9AQuJ7cTmKtzHXrb1yZ2CsWtNtxE8GsdawtA6S
Xd8s00Xq4lezN9F/IblSDwa9aPqC80koOONqkjBwwbps0wEXewk2cTPAvJfT
If7YM35TAc4MtWShaQPg1pBUbflzJxYmyDroklcPQpg2aSxmusN1u/D1N67e
GWWILluaBZ9uyk5en8nGS6QZcHbGp8obD8BLsJ3Db9oWETTGHeyr1FTa1rOP
n4FD81oYcSgSA3LkDXyy5ZIKR8WhNqGAMciH+gdD3TNEVl0BS1iFEZ/4VPhg
5z5lEqOp/IQb0WEwooofT6yy0P0iwwGXILgsF57JO9URI9GDHs2RJnJ0Q4sx
iY92h0CqN2yWZFWESNn+kFKUBTaWQfrof4PBkUNOmPeAP/7y6yb9vWL7fcIU
xIoqv47LlGuY43GAXs5vjo1W0YhapnVKy0UORntUxJsIpFman3hYKOmsd6mE
+WJms17uh7W/SOXnlIjUluOZP2yx1ZDAXXvMrFJHFNaqo46CLfM+/uyImUuJ
f16tr4TfEuhxAcuZ8OivVvOe7Rv5BPPuFa0l4x7bI6tqs9mYoe4UJILC/bo0
51ii84DxFQxm0Rt5HwNlyDwE9m1E1uLyQhBniEhYNnVLDeQAyl23yPSP0G5U
i1fAcO6mLt21lKoWl//vLeamKxzrGYmzmJy3HZT7Gl1JblbSZM6W78/roSG7
Hpm22ZLyiQZNOOQ0MnLtR1KIY9mNMtL3ps8iDWMTOPBYCIa7EKvzArUwOi52
GlVNEF/AtlwFurb72d6m/IKyHc22bjZnD1nMFEkV1bbqyQ0B3nNm4/fxudFk
FHBhq6xT40yivbrchLqbQ4lx3x63GELBwGzip0c4pRl0+KcvIDcnWYWba1/G
EF+Srbl/uLgvoPCyyW+d6/wfmRZRzcyja+r4VMP+++dxp6UpUutzg82JcHaY
QhoFJTBTpWkMVjz5g9LDifAxK72PLqlwjcR9o9UJ97VzkVVKhonupgICol11
JfKGJA2sb+VHoh6NlHo/n1iCnZE2LML3wAI47gMb/fLwSw4vCkdSQcc53eHe
donWiM/mAuz3sxXS4X8Wk9bUA6CPnGIuwBPGblJkcYHMrmA/Fusuwl9TbtEu
Rx1nL5S5mpqh7wMy04XLzFy4aeqgObOwg5Cuzl+yqlzy3gg1Mmg+Nmu1c0jy
BbYF7lyKIlTQJ4UZLb8SG7iSlfyLD2ZBiPNnuf7uStRtmVKiW0f7qsnq6n/B
PYfbjkkm6anMp70IrBqs7/mVaM2lhp/3laLOZTNreVJ9Xg6Rov6pcEpH1Ml8
BfaRyxdaclYxuWKXX7R6UqkpxpWJpIA/WNF92E17bUzvmcmhl9B32zlvIEWk
osXYv9JDnloRLzrcc0Xrk7hzt/lzp+Hl0AIeKEhz2rRkHDsGUtz/Risb8inQ
t8mmUU5sUYBhAwiiLIT+AsYtz7XMCOw6sUb92nMnlLgmH7q1TNKhLgAndvrr
uEQOfTj/3f2l7ndwpmJcIGVkFgGQEPwN5CDnHhTa8LEWOlCwXVgDSyj/Im14
WN08TPBAgGt/Ih8I/Q8N/QiFMwL/eTDVDAEue7bs80bFiZL6/5pS2MqjK6b1
8y9sAR/kJHRgp1+Kx5sjm9/xCl6uPIwWu2Ko4We0tX4XxMM6IoU5D0ZvdxpR
lF7NhUa7GrK89uFEUs3AqLuyzoh68gnBVTwAgLG22Aw4AUjFr0gzXa+NDB8/
ySH/T4noYHAxvlMej7NVKIetUhGjqGEQtDY/OyOtkzwLmhYCl2O5R/B/e5YM
5jmdJp6uo4K6PpTAjLPXOjQRh2jeOSu9QMkuO+9rn6nDV/t3xh/fvKKrKPyL
Bl7l5nG3oFnI9VK9/JdykV4Kk6aqV00QstnNyf28BfLugtxgrdRpIE0Pbr5O
nPgOCJYfdg9YdGWf0ql1Sh3xa4ZXgI6ogivarkwUS5chi3luWiG+wforqZ/6
8qHZDcxK8GUbFAwoFiJOyv5eP7t8JKoTAsI99okjLT+1PRuMJdZX23TdStgW
NSfGA/SiFuXFeBY5dGG47x5yvCi5G6K1XsuOfbLTKpPmWsEYEsTEmBMlLXRa
dhfGUJhgOUjaUZiSNeUStxDpSvsh85EUMgUnJDV8/uEYkFHGntqa8EGPlWKo
369yN9nLCbsA5MUcWWT8nNIfL8NBZLJcx6LU9qGWF0nE+zLEinxt9XDKJXWb
aWtrK9v/qSjiJwjshQu3BQ2yDIQgtLwT+UpowFSO41KUy6aCkOQ2vmSwlZ/i
oFM2/ZXgcznsKvmJ/o+lq1uzbKm/swnsk0Xkh/CYNyvCOB53/XeS5I6+9+by
iG9ssgw2rJHXh5iz14MQ6pAjbUuPv5k8AtharnKw8MToWBCnPjEOXbi2qZZu
O018pcJzpHGcoB02SMltFuFJtGV6MdYQ4BBNojvrngaAkxtjaNRCa4TMSo/L
3gcPX+Yd2IymyvKySMMh1nVkg1oKu+r/tmrzDkvIEs0vQDIf5SzIsqlwG2zy
ChJ8B3+GPwZl1fEaD0iG3BUc9spUfIVByl/YXBGEvrPPkMybPrRT42nz/5xc
WMTMreqr9l8udgdhOxFpPtECiawyYvhhqOMbpZOXyagal5c23hxBoKeHoXjN
y1s2xCaggOsNkcsZL3SzywM8tL5BqrosSgr7/Inw9JEV/mW0I64EGY+SEfN+
FYzY0hbsbBCM9LEplLrG4KgE2i5FXgyvxfJ5noZN2eisN6TJZXl6/B1hRUTZ
u/HvgQ4AJuWn0V9XXEzGRU1d1MTWFLwYnDUrIVoKlmWNe0B6PQgQvU0bRsg3
+na505V74eyMPBEzrG19CbZ8Tq6x/WSXQyhco1459aEOKE+hKCOLGZJW9oNj
fHN16djb6+L19fNDCOHY553HfuBhssO3VmOjly0dsEiyKvYTDPb6Uxdkd6kP
bC1PzPezEkHDdP3GBPX112M7M8FrE82z8fDtzAeYljg9COoLa9fC1jyeZnQ/
+PoBI6kTJ9y0kCkSgwvW4HO5mGA+asWbC+kREfbVJgNvX8kb3ga/ISluRu3/
VZipztS43X+cdcnIP5nhdE45K1xrIq/8++2TlfGEUx6tFpKX/yrihAfzhRka
+dEFaJubVcQ3IYJZ1p/l+hm3N0ADdDIf4nOyBEaWF7rSNQ1ZbCKtYgTFDo87
YhKC8/5AFGEHfkmKN9zUU69c6N5G8iLDkTkoyOMJBd19r1YjiJZFcJm4f0Vr
bn0LNQYRICjvj5OM2aLUMAyJLf3PKwdBCu8cdmgN0RO45JNBJREZ0avwugiE
JlsGX6RJeb+lm5QUynjvqeF9dFXwToJcdcMb8cyJVqaZHiJ4PTpJx1e4Aq6G
tVubyvpcPaQyZdTYZX703D+XCeJK3X8fzTMTHGOngGlpe0u4MRfmGKj4oxqj
/OitXy7vdwrIzigyCkQL+YpYwOPwk1Ke5NMbxkGEIRYxi0sVM8jz/64riGzn
/jM1z0Iu1cgjRssNjMMF2rDR+jJP1YpiMSGGw5vyCjxqdXGN6+QvLq5xUNHO
MYU3/gVDW9rJJimysx4pCknEKw/aOj1uxs3I6wJVfFJ+5v+O1c+Vu3UL17if
FRxVCndea4+H21V2Ta39bQHGgsL3g+YKPKKkBZzDowpOgE3yi5D9CjKySFNK
Le7R8ww3uma7E6UCdYQZNgcf/irYOPGxP+AoibiyMor7G/2AuAEsy4td/+II
wRVxoLPqFWrYXGpF9ABuUEljHBwPPVBNs9pdJ5QCG9w6evUU8kcrg/EWmZ9z
eS2Fq0ijVaq4JfyFSdJtR9p8mVdOA8gOeOQUefZ3ToL0Va2UHITLgaY1XAzx
D/3/V9IwvDJ4H0ZJ4RX/+Bbg+6fZQlZIqwwenehw3W7b7cKC/0U+RAiFqLh8
KEtlNixqehZP2mRW43d97mvKTN0G0fWnH5pS3/eUbOO2rSBStFhP3+wf/lZV
8tqDz9Zct+X0GfhUhOI/l1APFzEBVfR7OGlV51XnI8vDllAPbGyt3+/QOKWd
LJyB4a1Dsl/kT2iFNLaHjqhDGx2nyK6r1QOubIegx9803zt0Ev121lBQQkGK
2MFj5RDpk32y+8Ot8Zdmtg/IEOmblAAdr1/Di+sdsEcfIbxPI+d0vJkUAn4F
hPKn5IA58Qvss/+VsmDMX0b3C+eX6ZP9VBpoQnisiF/uAhDkqw61+1Mz/uMU
lxzOFj0CN6BS3jazBILnH2UfY2jed+sQd/4kXVBC160GfWuIqLwJNgvx8pw1
8U7xA6XK/nWruO0IUMzITShuqktv0vNLiioz9nWb6uOuGQnXMZffMM0yThR8
6ifscf9SaZlz3/IMEy4dc18KLvgB56RIflIwadnEpiEQ6gIi0jDWTZCZeRFG
jHx0urXVR8gdaMZcftGdBaBMEgTwAzPjK/avVAEQK6Qlyup2XjrwlDT1OGMj
xCRe9n9XaDa0d0VUnBvZprkeMUbxsGUZosZ1+7rE3sSUVTcHD/Wnawu3yEMR
l7G+JR7UiwkTqTUaP5Cf47ozsAKJymbpWJyzCf3XwZcvOmIIF6u3Ucj+VYgq
fbfQZUsqu0D9cHkXfE9OlYRSRqHfymVIwEpwc/iEU6b7BY3DyZ/OZuAgP3yM
+lJ0j3pNLLgjJly0tXwZDX7rj6kqWFZ8AEtD+YA1yx6m5WHcllhE9GfkqGu8
C6pc0LkeKezV+jJxofFLNdE15gT/FxVtfjqFV38fPYUzZRKDFBOYFQZ7A0u+
LVKOb4ZVvsBwhu15wKAPADtzfyX3o9kHmJ8sq/qMVgmZ1VsQx9b7C70jNdqm
o/j5s8dRk4QWR0hxL2gp/kvkUwvlVbBT02hIneEaDbQ7NKjKB+fuCa3YnQTh
ZKj8lu9v501Ks2kEwL9WACMbG2g14Q2KfcjvKKi2G/CZg0zNnGbYR7H0wiiV
V4MegKlyZSEUMJRX9opj93426b9d3gcGs7ua9vUyu/oLaMQty2HC1CUdeqFx
xpRaFWsht84wO8EMooGz62RA4KrZCrvBC0S9FTrUvK/ZtaezlK/b9mefzlFn
I8Q3Pdo3oPA+z6iKV1Q3+80uKAW9hJfzdbawH4hyN8wb7H2zypYVFyDCO700
qP4TQeZvv7Wgyke/z6ps1B4rFLnqHYbamxU1K+Ma4wV+QgRDUgr0KXkSW9D6
ox2X76spnKJl5852wtPpA0ktDVsVg1VOdeAZURiopBw3T1r/ZA+IG6opSqmS
wS1DuNz5lw4DRtHT6szVo1FqVXi37AScufHuzrjnX68i8TGKQMYc/6iFWLE8
Mly+KHtsj6OIIebLzSIIuG+xHKjxidON3JNKULfAPnzsJW7H7ZaDDwhq0iEC
D8iTDqfm+2n1tCMRmHRbsMvzGL3hW3GQ53v9tazuSUNX3cuLfBneoHLJUBcH
QTediCYn33chDpDN+JfQvoQa2QzK5ZLBFFCU7zj26j96Ov7D2LAhpxoD52fS
xWiwmvVFATXIurPwpN7lCOXa6n5uFjmo+n5dMbn+5+nAO31J38gm8TaCBDZo
vOhZki1jfzUPvACQKBXILhzjwZoes+rjwE9zjSYMTGDLLRaIz9uZQAj5C1OX
yWnAKlJw5g0nmeix5Zb0ZdhKkL0DL45EUKMD73eYtNK9uOg6X0ChkWskg1pO
/+YXWooQueU3SirCeq4yZM9xdiwn/lh1EvJAIt68KBbkfIIz/OvVzmwQJ1rl
+o2UcEJ3pVsCWL3CBqTluJCwdhdFU6gfs4BKercN+mVDnoLNDf9qM7vTBdyo
P5RJh1LyD/hAwaLX9kOg29ps6M1TVkRzSlZvxc5JzcfT6dGiI4jNOKJK8KiV
KnU+5xoOLbdGW18fqXQISsQniIl/oYS2qKLjmb5sqzh5RbxPy6Rg8vPkxJVU
qv1K0sUKh8ZmRKuOG0pDGO4cHja/NIKD4DCb9ToG8y69ps2GykBQBgMS73XD
qOWQPHgEkWRTfC/3x5B2R3/v9vX2wBssG8T2EFohoLseT06PiIh2dIilBRpY
7lm0BdOGypjy+L2He9SF4piv3laDCc/lNlonVND5TV7nrn3Ho8M1ngbcF00F
RQ6lym706ucgK4tCG+VvaAhqQ/WbutS3PQnbrIAfEL3/mrYca+VMAcXWhzun
lFmDLQa3n80MpU/bxhAJUrbcr96oLfkh1OpkiLUbi4pmpVcF/7bWhVCT5VQg
cKnPfywchJrSp03nt5TVXBRa+9eShoScD8DuEO/K4lbvSdD1uxFQxHM2YAjz
KCvfMyGoJbuMzHW6rjlgY/KAsc4rIzxTcv3JotqitFsIWlQJ/+M99odRySuU
3gZskq9Kw0ln+SzmIbhIRMMTCs4DSJOAAVVeq1lBd/fdLoH4/wC1cFOqYjIx
agpvPQrGsJu/ooWVj42VCNOcaWfun4HvGVyrJk4qFxjxrhO7W0Wd3h5bO5G2
nGu5dKd85kGXBRZ05OGC9cQqDxl5SAYRbL84KXRY9PzgRL/Ri2fZ09gFQrUt
cUVQ+7kPKqZM6cYi0jH49uJgdsuCmTVeurb5Kr0cEWVh/e81El+V4nL3hGsa
K5kykeu9xfjelU5zKIDoaSguhxKh54UYTmHMcVhH7AuoBm4HMlFFVCzuYyIK
DaSwDKM+6B/yI0UeyLjQJfuA9+LI4b5i/QqvJ9e9g6t2j9KEUuogRgRmNW9E
ORyAxkU+BG/7jwuOavBqCFDTGdxDculrNBvdJwy5aHbB8oL6Nlw2PO7wYQpS
r4U/tKeBnmUUOJxu1D6JTRlBioAhuRe/LHWlGlqN4clVPa19tpuLOjglGpln
+QHiSPMsSH8u6pyRsj3Jw+gx4L4OTygZ0RTevz1xId/yvippwZQIdArlx1Kq
WOvqnoPl+cIn/vmeFzDxMeHsN1jfQ/WreqaOky6gRAk9XO8uZBpbe7yqPBES
faOmhZbqGs1ASkbuSqOegO1ZVlYRgMTdw7+Y+XdUoa3FH3QScTM8B94p4e/2
A1YrE+c8B3c/klueQGbfCB8D9Ic0BQ6lJxMhjVJq1WBqaVcgk0D9w1GdBeR5
NKPtG28/lAPz7A9J65Qnwb+LlDILJTirTEpv7l05IItOaJAkkeMHYuZlE8N2
JDN0V22o7z7W8klLA3m2cHEFU7vGShAVDL2ljVYIKysYBEuWhgCvXmNiXqOG
fLDbMTbfGEckyx7lWyAS8NwJ1FHA6bccjl67zffl+JDBY2TBQf8iewjiwqoN
PA0keRPojUb7cjAQ7tQzXxg6b4IVHxw9KQ3u+w/EPqetqjtJIk5CNFONBo1c
lvwqct/FDCratFm41p0yJqUFkV6J0bP9qWQUUgnZYrmXEtaIsJf/troxNVnd
Rq3OKP52tzSxs7/U1nsbWrjexSByXn14Vt58o9smdccKHbIZNMAWPViDk9JS
7CvvLk865T4uA4vOd9JXnVXHdNt7wLDpM+vXFeLWjuPfBonxBBdOZElB+8kT
mJgbUq3FQe/JkPUZdbvpxlrFOTOjxkpIpUi6RRJB4NYPDIsd47fV1YQTAdk1
9uNHBBMzhRKHOVEDTCcxuJK00BBgVUmWGOeAUuVQfQdPhtl3JBsY8PXN3azD
ZEfB4N9t+VRO9GpcQqp6rgLjRK8v+0mFfcbdjJDVc5gpn1lh0LciybPRL+rw
9Wm3jYjmFvefFJ/gus0Te/zuLB01dEnIROKYTi7qufxc/7DB9vUb18JdXPDq
VL2mTe6+lxyLalQEz6rzxJzc3iJiZJGnjf30gcTH9ZY0Vdvhuif6WB7kxxf9
So5D6ckW5T9deX99ct4/0shAlieNiqkT8Du8dmAtey38UZnGOESSR3Z1Cf2L
ZbVGRRp7hIhvkvicyJOSVyiB4ns9qOLwjfubSkU8NLTVrWmGCAb9KzMGlrS4
wNxbnagQ8TjDRmndpTltTAw4xHk4Uk8k5ZX8tHyy1ATKf015iGBCCs+gcjcP
G9Uycs1ebu7WC98nkJyKNxL+Wlh8KEAO88K7M/TF3QgiWR95aeVDBudGdpqk
pgHsFM+hXe4/l544IbMMc8p6WdhEz8utN2TC0+J6+skTkJYOcUZCBeeAp+2B
LepIlLPMj8poTk2GY9q5iANISLHvtJ4FtL53dgx40l15lFYX11uH5hXuXG/o
g4TcNgWhUvnI1aPZbhDgfb49M7JZkvHtHCdFZRCVP9egh6MAUFHtGueTrMAe
0SqPH4rExigkCqBIzJkBveIKTEgKhOqzH1MTcBvUPJOQ+43mP3QIKMTPdcWG
ZophxepjmJ0jtD7uPmpErAL7H4gTNaRZjqqwYdCvDKeBs96AX04hy+oLZclO
YRMJ65OyN8jzIXIQCCF5J8VzODpvCHoooy2trhsTyLJLh6c6Ii8X1asDYBI1
eASwC0r8MNZc8lH1wzbKq6AwjLVwxaupQwiITmlLRa2cyYxq+xhiM7rgVVRo
L1e5PpWs33GnjP2venrFLCk3UmF+sTbIFjlQkwbFl0VO5UcOpQobD89Pu2dP
mEbhVLwz8v48Nql6jxYh4eJdUVhsRUgHpPe78KDzGRRl0ydzlKTFXAXwLvRU
gOZKaPT/QTe9rd0GH+ltRhoaazXlxJCvPc7JJWXmwkR5itruOVHryfFtqllO
hW5sHE9S0xo/fV5MMJ2PjvUC9Uzj3BkP2J3VapesrRxPf3lM4MXCznMU91YW
hhAIi7HmkIaUeoXzKuPCB7QuQBIImswG+L37iqkgN5aJdXAMd1h1BHRq9pYA
we6fOhPj8MKA//Dp9j6j//5sKdcg6e28n7Ekaf9kS/Fl0NRyw6UDEY1vt/Kz
0B4trSUFPE7UonMJqDefSdERzRW7cfe0UDWbYIQPWcJota7RxhlT8Yll1Lvy
eYehJNDO5h+8UKxeErL3VxTGQvji1HW6s2FQks5J4L86Th3j65/U89L3VBlV
iKIujO9+O09uqfNsNCka0x18CVRizRz2yOpT3VqzDe6iXXXSIKT3/SRAX6ar
aNxKhIHVvpy7CglYThK1goQw6GUESmiNytEIO1o8O2OPgwedddXgLAs4B/1a
1+eSPmiuoyrcQGOr3LbHtpqBveT9vsIyKhgXGH1w4hwTrJyKLAnNESnd7NSc
U7Vt5ZQsmTV6QkWiHIRojGUA60RlZhxwtEESF2VojxGGGcyxoHBvgiDm/shn
l2ec277AozatknwqN79DNn6l4Ta3IJfGcDY2gDn6Q0LDEN1FOMT5smFvsX2L
2ac8/kFh12ZM5Ped0dcOatD8TamfcF6QG7caQrSi1GHajlSgl2yPKxYRRa8r
K53yeTtHi8vGi6QeFPg6OZYT7NBddPfOujOJtg+H6wvfzD6U/tgg6W/DfM9H
2KkN/UdM0uuF6qGppJl/0y/CnEGrKVJ4Sjo51VMz2kWhSNDv+0p8nRQrB+Zh
yDra+bkL/6nhTuysDpZVHTyrhu1Vz8JCldva+Oj82/ZrPOL+lo1a6YdIJsIi
1dFvO28ugHv5aIYQhmf8afTwkTQaABS0BmnaNi6aVkrkW2hPAgrR0ojdNIPS
IwolWdg725bBwgQsRT7g/KE/WWoLZFrtyhAlu4nvO+zGaEyoAXpzFFPixe8p
uiDPbcS/u8dC/lRvakDVAJww3+S/++L+1ZQIB+eRZPpqwcEuogkamgR4/eEv
T7eT+F02o9Oe+Yq/KRx95RgAvAzu4PMRxAA1gCYrfGmMx8iHu5WTagAsWrOt
ksXmii6d+F9v/WT8krwn8bWNNoji1TjSxuA8xmYssIW/ZwHb/cQ7bKMO4T8k
1VqsCRVfz7vDjXJUy63Ho8sQ315CDK5dJy/jP2acptzgtEr1f5cw7cd5LKS8
ycqBfze79X2GUPLf2uK8ODOBKBDAtgHtD3VflqryXZXDvFUQECnv157fYokf
gSwgQ0XG+AkkZtY4PEOCRcn9gCwV8gCuaaKjtrHo/IQtlqig2/prkuLtc1xl
x/aRyV2TkZ0kAdiPGBJNK1paPecZqgrMVbQ6V/zTuCBr6EpklrPaOcrJ/ZCk
6fO13s5PWlSO/oeQfscUPbRBtCgraNOPiDYWfZOlwByBICIIjMh3v3E0eTcl
wibmrHODgqhDEXCApjVb5amykWT+YViEy2u4GaHLiG+v5YVh92Pub7tqBI2/
hP8xkTwojhcFjn/+5x3tvl/ov+WoHpuhS+AaRXFfdTWk9hmECuY0lkIDy5tn
wS9bWNBecSIuY1j3zK24iP9Z9whf3Lny823Y14csX/SMIJpYKffIX2ayTywp
sRxs+rTziZMg6tr6d01bUcbyzFdoBc2ImQIgWfSV6VWxGBxyMdWka2W+T4nH
uw2fgivkHZ9fM+gGeRCh8bNIHLhN+7cKIeEDMMScAH6ZgB6FeVoTADaG7ZvL
BbK7FBjZKW3xirgTHrTdd9bCzfMvirEbjXTd9DxxhPD/NSO82kztKdxGv7nE
1kBmg6rsYtg3+0347XJr3KblJMgXEfySO6qce62r5oOaucdzV2wZTD4vRSt4
01+9jafIhZNLCXg453rGFP4oM4S+YYMnk/3P+ataEH/pZhG8vGPUmD4otbZ2
pICdvXrS3yQSABy5C44sIPGBbzKtL9WJbJ2feL3s4iT2Y4jk4JpGZ50IEv7Q
gJb7QIjxWEf3HNH/HuqDhI0+Vn4tKFegYFKp4wfD4MkMgniDOWLrt9rHORGS
f4lEfNRf9OUX4yncP49UUAzvgM5WMtzv/troBR/WQejY+IDUzvZeVLmDRKym
bgGOj0jP59HQVjiYcr5yzhVoV+0cEZsnHPxnioPL1o9wEQtceyEfwiUvT8th
3WfCf7RSQ8fGk22OJSnUkPtf+ezSmI6c2Lb40OfD4yrngaTLpsUY2dG5Fnwj
/kgWX/I46DC60vtC1W2y8SPMC0easGjD5RzpXmUxnrPWBUAg0JX7g2fa9sdE
ntPmJBuxxl2+6JBKOQfW7zxLtrIzsZJozNxn8kX5+Atq0e0S6phqDeeSdxpn
QzK42bLEI310gaNBasJ9pDdhrTdcZiDKQ84MfkR01+nkvj5xPj0NiO18u81J
TIYsJyFYUOheVKgbTx4GvGlvVfUJiTmeKbr38Y0S5G+0MTH8+HG+nl7MitX6
EukOhGxuDHUZmZv+qNYb+shCaC59p43vkrdBev4VKEuPlx3d19E6Hkv03N3g
znJw8o+lVIoEpZ81DdLs1Td5voa2NjV93932/qlVZ9c6R5stce6zHDHv8YMs
hapv1i3ioCz3tCkZ7vl75HfFf7izEFwTxvvQ5/703KpKmuHjwveFwgef6S8d
ZeN9laHXqv74V8FFvJjpAVWWGmLagmr/3q1MJmEp7B2q1enTZ2cpTa0AMhgp
JdwdJqMYug9+kjK+BU4AZ4s0oSsC1UJ5MfaWCZyuPxym91N1YVrBa4KdVh6M
v0iwCWp9b6YS3vcgOfOTlA9utfh6RdzayzLGntQTjitJzk+VYh+kFJEdYz5s
5TUt326Wbp3ph0U9bj6BjHQ3m42r5KK3HLBGLz/+HqaQpZ4aUUM9Oe1fWKHi
deWPhVTsIBJpieziLwxwx3R+VBax5dC2qhgPF+zL7bZ4bXiyhF/aG+gx2nHE
KK8IHq06GxjxBg7QTgbSACeme0vM+TpLkbVztZEpKoB+auhQ+qttdoGsikHD
V50hXP60DSsqUyG1K8A23J/rLzybKqGs8pXs8zDDqLc7KoyreybsjprKkS/Y
H5Z2l9iShKuCbammks9B4T76udpflQaoNbOV+PicbWHb+Cp5+rRKVrA/Xk09
YJ64hJOUIrSFUDMH0OPErQsNv735lYAsl7E8JPz8+W+LDoq+JwSzwV1grd0u
EZThp0syha8MtJ6X7qphkkYvGGmS5Xy+zy+mxhR2cdKhKqrX+9vsPsPk07wp
intP7PkGJMg4LTNkCcebatoMeOUrtMomRCOXLo+9ZUDX8jxoU4Ki8UQAFy8x
bDm3aR5zmXVR3osyyQOwNIq/J60e1P0bUs3wDblMNZ/96SmOIg+8uzg5+VWc
wOZbH8QrtLE+Mi3Tu+y2Dzg0A7oRtJKOel3QxphgKBQA6I8cOnKXh5QiUsZP
GCLByzHOn3U4kv9BpTSXNR+EajcGmP3yXhCHtG+Fh5yC+O4vLcrimd3mtKKP
kimeN8CTMNuTQb3N6T0IXdzE9VabDu1eMaIrqSA7heT2kESyAhGV5QArNxUn
7GSUndNSnGJ8+5ntx39wqxlxV8uncWpukE+5ro7rLhDeVQT+0/5f8Wf2sAtO
KVJgAOz0o2leELvS1DF27Ai/x20lR3rvFYyJIIkpUukwDUrH6Leny3aEzsDO
Ivk03Gp4Xaae+f5Yr/5katoOVJI8X0wG//6Q8HkLHFlm4DfwwwMQJNv2nn7G
vaZRor+aY8zt5Z9iLkG+PFoU8YMJ0TV2o/lnn+98wIYyVBVXbWQUL7/MUeCa
GTXEGbkczHlFpBFlz/bckWyv/1p640clX+PGncPihyZRLP6BZtZDC+V3kva/
8pcqd19g2ySjcx9kAF28THp/cJCorv5/Ad2AlfZ1FcY84JlWxA7LY9O8CvkH
N0Y+rI8rfC32oZjMv2YT6BgPwSjL9HtEgbPAomc2dQ0OF4odhTj9hE2HagIz
LQoqHU9izQf5tTn6u+cxdbYprpbKw+F2fYYR2YmfC65HeKj//3Iv5pG+foTh
K7ccBwXqj/f5l4pRumQS6FWqpg2YV5RBa2vReBn7N2yl8FI7uVXMsBrTcR9J
r54a5J//DIVZbvehBsCbQ32Belmq5RzmvgpBPeakIC2+jnR1ozbQmxESazHi
YKStxrBhlJo75R/Nf1Qw4wa8bmB1xTVQhDZdqBTIYbMltuyQfu4z1caWUDQk
LT/d6ma9t+CMUT7HhUgDSSit3PwjG5wJub8Q3U/dY2Y+5KOo1brzQsO2hcIX
DEP4l+84eE1TGU1fbloePuAd2tNMCk9QifCGL85vOTCwaU0n5GZ4AXQNXzcf
0GYQKQ1Qve6fbR1LXNYHpyIh729v41RjRqtb+vcu+0eaO322ej2i0kCwQpZU
W+QZM/cDDOgYgQfuCNtT9UKP9lWCu7WBk9Y0XJY9xiFXyUYzi8Vs1PL/jiUS
O3Vmw2tSqHR6tkyoE/Wlek85DOMGgAVnwhjrWqGw9eszIIulxRWOTOnfQLfL
iM0tUkOOQTxwVVmm6dOFrZ8q6khbl1tjTOLlJE3WjV0wgoc/YsbKZiBAsEPn
kFK8PWTO0JD0uaoV9dombJ0GatkLmlYWYbr8bm5td83FLpe4lPMXAF1vPsAi
2LVknIQkfJpff0KXS4CfOoS8WdQS1yFYzdebfSj98ULjwrRX/8djRF15hP0e
t1K8xpMwJ6RLghBYxYtnR1AjuSTcsz7oGeZtmPKoM+cQFmtRdiQDjGzjuWbj
NCOlmh7CFjBoQzvemcZ2cVQieLaTfuTqrdQDPqLGmjw0MP4p3u6Pp2ZJJS9Y
suxaco0TuP2kDh5XxT8Q3Bzourmk5zqlhrjh9HJ+rdabe6Ia4KyrbeQm/xI2
7aMdKRuN7XT2AMOx2+NtWF7kBczcxXIhRZgFHGGLxIHsbw9WAjg9fcHpJxeG
yZQqEmdVXY2tR0L3irQn/AynQ25tXQPpZWf8Uqz03pDvmgWQqz+3W/4Dkdl1
hErqqLbQkvritCI7NEC8gwPS0/xz8Ut+gwnEPxSTVhWtvZT5RjAhJepqFrBc
bstfVd3n+pPkXoLF8wFYIDqQlZyLBCo8iQKCO83OnZP8ejx8CrBdU3ui21/z
MJ9/fDMucQ08dDC3CGIiqYPxrCwMiRHGu/SXucypVgerUEDi+2WQl+5voOgc
N9VECUVbHeHTKBkHVxKfp6+sAT/0Dw0mxPfyKvcKnlV00loJ0CMRLTB00ePD
Tiaw+d3hesNcOZoZpUjPt5EVWO+KL7OjZsqq939W1sR/Mx+vi8ZO0WvSuJXm
nJfryeTiAxfF4aG88KPHlnt8E+8UkgcY2wAtSoz1yXkPJsYZ0FghW026O3mD
eU12gay/t/x9Ri/dlKmmAx5G9ndaJEzPYh/9Z4kfwcLWFe1MO3E6PmbWtp5E
25NrXKuT+fz9BBjc8+kZI705GTrMvWWsFs95P29lG5m+sP2qmDi7IVud8GHh
0UJI5a0uzm42rDvpSKDLbF4vMikQiFNSFed4VQjcNrQ6ulRIp2LAe1X0Nmde
U1Da4L6jw8JsmYzB5qUjtUiwn5LRvyhhmGeP7q78HuJhqaZVjPaSZfXuOUMj
8OTdQlmT6pVl7xbYjkFshi3KZW3SzhiBTDc2XE6/OBzW2uaghDgXfvuP9lef
uEca62DilOpr6FZaZjCuTwGCi1e9ce2ept5/00A2qEhtNqbAIexy97fKZs8w
eP1psFIHVv8bHK0iSJXUTXFDwozFv47zfUaEhkaCB8o9feax1y6Fsk1pNdh5
CRbLUiOKn5ixYeXLAlj8PbFWSME/4n3T8p6atXTGyp/F4GVS7sUQrkpQ2jlx
+P5wbUqPOng3GaAF+IvBsO+p4WPS8g64oxVkrNvP9DnmwiRQ7kpDcXUielBq
Y+Trlzk7yEVmoM/7zQPttFh4Vuy96gaiHUskcIRHarVaCjm9a4x+WilgtfSt
6YsfOz4U12Omgj6L/bpRJ63+owDj/FrnTy1lkQgXEqG2czkH/IoXArzOgkwP
Lg9U977Q/BgxsTUtj6LfpuLt5ALewg1CWgY1UVVmwS+oXAi0hFbqsK3uNJeG
woZp09ubxvKtsfjtEa/1p4WtRKHHLaHIvZ38Ys7LQLCxCk4LYdBODG03XJZM
Llcinrd/fRnp7olU6ylc84Vu8yv/MdSdxT+uPMmh5QvmpGUCto3+SuryShVS
mqPhshoWt7twpWbM5/9GyhvzeTdiDW2kpuXn+2G0n4VCQX833kRyjOU8/OnS
u5vZEqWlH69Cb/oKinTzTsCZXBHCtR0k+seUmI3Pdydo365uMlQf6UQIqhg+
SD7+yy80XafS4to3InpGcUobxS4BEv320PQEFIpRSpj1jzbanGojoP3CGTit
uGQ62gO4xnKmekgKJP358hymAmY3/NeTmoyPc1NiCQzw813KEFU2fcjMMLQJ
FE2AumBdKFfA+7RQu6BZxPZQOq/pfaljCXJ09VAgT5lF0WbV2nAsli3JEoUN
smQ8YCVowQwr5+EnXvnZS+qWGkGV+Wt/Gl7N3PDn87KJKXBBM8cNiAn9faZm
2Aky57UXxXvESC5qPj6217EoI6rXoDx1pq0SZCg2JnhMMHLZbiBpcEoVJaSw
fyeUIp2x2zdIctodatkWObmVtPoUvqDbU4N5SquWz5lCVr5OR2UpNUq6HFYR
t/JEEmihF5VthEbaIloB5VUIO16aDp+/SolUU7JQCwxBGPa4Csho57CHcY7V
fBErOwQ3zn0bc62bbp5vxFCepOeYZjDwfebsnm7Hr6TGOHTBCg+mWekVSBa+
l2/FQmGvjFvKQkWiKHlzm3/w9HE9X5CiVoOQuuioPckGzXLei9B1jT9t09ir
TOLg2rynDPOtNo1Dm3b+RZh//Q2M6rxbXGr82pDLfNmZMoOF7kiC9t99skvm
PkNFzS/iqimm1A4iNIzDHMiJdSaxYMlHHk2s/DZx0ftjin1yy7a7w7SzsalI
ke8cCGL5fzUaphpdl324R878m/3IUuoqPxth/cM7mee4l+tpGy5LOH72OL4g
Lus1PDWwNT3mxCWp5rxUeQN+g2yTGeqpw4JlNcwoMsLs2s1JQrRYSg6cSdO9
Iat+VZ6SggCGx0PujqUK9q+gCYRl/kEVQ7NCHPlUQWg3miqamDryUt4XeSr8
KtS8jf6yQxeUXNAYja0ViYuNvEOzQqe7DJpfO/u9UMydc39qSl/w/1KeLPHJ
HNPNsqGy+rPrskqe6p4FPKDLYnxlsaQjg+IjZ5MDpKANF5XQSMyc7qvZFnPu
t7rl6RweRi7sNii0kD5o+iHEqN3C/7Gd9nt22jVnGr/Y6kZTgIMdUsDX2j/p
7wb7eek4a1dh6X39r9YXHiWB12b/RA9lfg/2ZzEDq+oNRMklLFLPm8jdxAa1
d8d6DfrSLuRSb8246Z0YxVfwuF9Le4qfG772cpjNBKevuFIqzc01ijICjuDT
+YoXcOaKTMGg7wA6vUwifEhyyU/KEJSXFUXy0Fl9RnOjAU1tJl2tsYfovQHq
Lyxls+kcAMW6r3ZqP8EXCLxPOVp9lCjI7Nv5Kn/qVYyxlGSzIhllKdWzdjyp
Wfwgr0w02xuw+w0WP5WwYrESncA9x2Of6ry4xxMzz6SOtn1P0SYvporfk5Ss
vx+WwLP2uReBH5XGdZhL5ndX2hc0O/Gee3XXwW7dgoWkZgcMoDXQofQN3h+m
nTUFM/y69o+22551fhBmG7U4yJ7pEuP/7iDumGkqUVt9YInWO3L5R5LV4DWu
meolxbalapgZf/whVoukcqrD/+jm3+gR95nW3AOEK1DgxonVHhl3zkyyrKpw
xk36/WtUpEMOm8GRw7aY+ca7JDHx9WpwvY32rnMuv44ilPUn/bBgDALuOvxm
Ljl3znVs69Ipn+CG+RTOgr2Imfnk3Tf96Ni2fmO9fayB5sezivNghFXoL+lc
8xv43TRIXg+km7Oz2TUylDbUSbDClIrqKbwkdh8OeZReAIIADueqdDg8I/Er
98CljLvyU2tgLuK0xjdntC0H5flKsBCU0pQs2/HeD+eM30ylUbeY8MsVqWmd
UCIvM5ZpRPKdWKe4G/xYdgvQJsZXW/a2EuUbAaVnngWTylmQAfUlWRYFpfkK
Yr9qFJPti8MkLnbinv79UQrSHm8hybObDNBI89azEMGCZebIJTVeFYkNYGn2
YIGG+DanFqxiDSrU14uuP8rxCGr4NpPT5n5b/lCgu3lsd8Fx/1p1Av482bKu
8aKHSc/l3xzJfTb8JvxmBwDmrPoGWWP1HlfNZG+e8fZYWnP/2TR0skJiqlRU
fkg3Mz0kqZxRTgClRK+Dp6vJq3ypEUjHONGgNaELFdCbc7I+BWtY1iNvlgon
h2wbFzlmk9o4z7ooKnxwYfnWkEqE4Js0Aji1q9ForXQKIW+vzh9pbkp+ac1T
pEeJx/7Sc1XhYnglPJFugmb5Z7k0FnIiQobIrZ1FS1zU/nCWljFLa7A2EE7V
yToqazgfk0Ql5FfOnc525Ujj2JcMWyJhfcIEzRAPsyNuf9nonK230vJNjXsV
ZANfbYL6G/7l5MPgTsNPNK+Wqe4lZyGqhdcjZg7cJX5msCsricjtPJc0ftXt
ypqgRveP4P1rhcl7XN1x062JSxzdVZjjU69HQvuGfTB2HSGbimqeHG3d1tM+
JlHtnWwwHPyZPWkOnc1J/LjkOVigcWWgdVi6a3rRWkXi3IlyYUbjSyUdBUF9
qQz1wAfUeU06d4Y6PGMrPrijjFmcj/bsTCsNZmP864gkWOE0CvNLxY3bLnxp
3AtazTnwjnHVJRHMovgcfX1ckDKZ2cgoEHatLlaD4hRTFluqt/W58zA/sFbM
2CWviMmnwTHdQDWAR4APyM6sYIFYiW91TkqaTD0BEdEms7xQ2GBHR6srh8wl
qL91NvTtcU+kWTLjujj8fSxRcG+PvrlZ77RP2LSf4v0wcEZ4jpmuggrYhdsj
5EX70Qiuu1YvLrZ9VCgYWRbiyn2aQdm3WzUVaHkM4hRmJIwGPbW2dHt5QwKH
Gj16d1dAVQhtf0nS1qoDz21JG6ldbV9yBFSvQ8ccz4fHRANYl0hR0AZS8DAj
2DOMGzFppnhQXsyFT8B0OKMSb7aD/NZszfmhIIMzJSKJVSZxGzp9W48Wvwkm
d+o7ORio1lVXsZ5UABmwWKXZWQcrH9DiwsBverLt2jmuwi2PPp1IPEmo4DAO
L149culcSaDxFu+Rhr5XhctkDZLYIPd8Uzjks1KeFVf0PVUGc9GZeZTFVgRz
c4LKDibnpw/dJH38IzsnfaqbT5CMpwgvjMbjLKcw7epePN4wgkwzg2v7Z9L3
y5pbiRGkiHRxKeBpubXbfzMJuQYx6jqGBa7NEeKUnz4nCxM4WHcSvQAGAMbI
8FzrRWsZiT6dmLD4eT/26G6swDKrzlgX8cQa0jdQVrFPIV3nuK0X4e16b+FC
KsVrXBwmoq/1XpYjqvg6uUTOMh7K+O+cDZhL3IBhd1JcACq1ETKT+rFueVah
vBimlO9uLL80ul+BM6wQnD1IXBZa3FcZNNv3skEWSq++mhWLS1Y4vrESFZYy
fSB4Gk2weQZTzqdHlcIdPdXN2o//HURwmiAyYgpvuXYpXZZtxUMiY6kiVlBb
KWwjby+t50UFaVo5h/FjZzrn9wkWlwtkfWc7882K9RCnOLgxK7nSPLn5PLiP
CYOC4Mlyi8jRHUv+657yG8jfl6E7DzmwHac1zSjijAU76W1vpZkksb02Ug2O
RyLjS/WWPss7PUKjwvsV6UCqBMLbYvNeUgyb7CrZkaj5bDwQ4W4NuARL+5GI
jQw4L+8NC56oWR4be/7d+KwhQ9qQU58xJgyF7VOb+mNwRB2VejkpvZJe0dmw
fUJKdiSmskH7MF2rSNSmVa3Uz5HUrhigVuIBVoa82RsSZZmtk7ebVM4ADI4y
wAO/4CTdvEqKdE9/sBiji8uAyFSPk9azQlEtCt4vzjTmWckgKyXmobt60KwF
ceU1Crpul9oX8sqa8RluyKvT7yik82aX38X3j5Dzxn/JeIfgqFPZjqy7bm3Y
2eMuSJJFaGKf4YrgnZajlMEZ9SOhg/JK5WCm31tY809uuf3+Ng018PHhfiaq
6vM/mfl6dfHM5lpnVmPs7+NOg76zVkPyEV3COAy2wsRPaxFoMntBIBDhGTg7
JgZfRLaXcSGrrjysWSZuXXW5GySFpjTdVFQ0hWG2MsX2HUlzdZOXJfSCEGOt
OOiy+tXoRVTXOP154q9sDf2JYTs/wkMulj3qGikw7/aMhB7nbyW8R9GGXYet
VkKDrI0uL1dGOjJWq6DwTzNaQFKjAt+VbjR7U2bUPjurdwhRvl6uQ2HFVdfv
ZvowHZHL4tGnf/myoQaG0xQHTgZtS4rsPiO0fHqwsATIjUSGknKU77DixMCb
KnJ9B1eF7T7R6UJ8+YOk4cpW5+EHELli53wcZQJykrNk3ex0lKupIj5z5Xrl
IyKSFKYKtKHcOT/5CASOc+eGXMwAJhe2g82ts33HbujJ34qJUwqJyft3JoVM
CwHBGx9W84h2kjJHVlYQoVEZ5LMcHf+yRppcJUA8YlXIkWHVBvOVIz0B/+Xj
/J1Tj/j+gx6n88Tzjpi/Dpj2AsERLV8qE/Sp89Wl8LLK2UhYwqBevk4hisJ/
5iXXODk2phBVsbUu4zhTFxIjB07vlxY/AeE9reaYnDZ5nCxHYXJoT2FWB2FO
KnWOM81bBDfJvtXBxFNHMBPRv8zslk2Ypz8h9zMJ5ynylfbxnPf+RfH0WZxx
Ot7wP9/oZcSYColRda5PZsRONMErq/yMQ0VHoKb2HsA0FRVRiEFjRHTSmDw4
fqNeIIpW3fOXaGpFDEu9SjrsJzcp5Le3PGRzhDu0vbcERF/fiQ5dYJBmrfy9
gFF+Dwxs1N5j/51zSPNmp70mMy9ZYsaJ7s2BuOCjUaNXysUWpGtNwHWuzSTF
n/YmtVX67Z7yuYc11iI3kzuybXn+QyC7gyI2SzDbkPlg8kz20440BX0TkeU8
iUuuxAtSJeX4EbRi4Xo/eJEzASCyjkmBMtFlTrE5LdBtxfu1N8FTUXvI2g1s
ECjwIBc75vVtC96ERWCoJu+Za2CMGUUodOGtE8EmaVF1WO7OLMLsHmZdsm+h
ajqpXGcI4UnZUnLVIpWTjYvEbbhdHc7lO3vG6RWEfg8LtbRWisP5QKPl1LAy
pHfFGxSdt0XeAlASi+kWOPRD+OfC0XDctgfyF/5005q4Lx5Hf3SPS3dWL5dF
DHh9FYxKHsDHACzLKZzZejgcy+VFauoKwiAAhASGnNyQzttpIU70HmpN+wQS
aUGK5Ekx1ePDzdpGVdVvThvvkg54C4UggtXowgAsIkzxHZ4NQLiUXAzFASL0
W5NbQdti0Cwm8BbbIJs0vIaUoUVYAYGVHXkDJWbRVmjNRumEh/Ip5j1jk3+V
pIR5Ik+/eV67NWUk8mexiLMnE6/pyytaK2ImKfZz3XqLVzcdW1Vkw0l8AeYi
V0NqjMdU4BiLpkZcj82TMaW5QoRgW2EtIWdZoaLH9gNmcfMqSAeYfkn3WRNt
4u/owtjuYL8LIMpeQGIh0Q4qqVAbnpxl839TtBvA7IcM0YQCUwz7VvFB+P9A
N39MZUXwJEKVHd0Ntm0+7N3szFxsfjLw/erXKrxmDLCsimh643oD9ZVEseLb
a4cylkiAQzwPtd8sQ+O+FiLVhaZ3OFE0OE4oRWca2vrGPk/XBubf/6rpL9xc
bVbTmAJeC+If7/FHLR4U2ZeAAXge4cfg4UW+tX6ojmeiEACIsNhpVP/Omwub
6MnAMhkOtMo3n2Ed8PTXBqHjILrCEsA99xfOwQE5EaxuxAEf8QeEiUhKHWsl
+OczzubaxrdzSe2Q/vsFe9bvkMJNtXlT5ijgpr48UAOdspk1wELKouu4EK1t
1dg7MBKfwN4IbWSxvGGsvgg+8drY35xn8k6Rwuf4NaayWaPgCfJiJOWawrtL
kHsk7NE8oD1elP9Fh9u28PR8ednzmQa7htGLS+H8pXjAnM3ceTyl87kpgTvC
0pr78TjwqjB0OqSfD/8zF5MaY8pNX9Y05qK+TLjUE5DfiI9tKrFOuQPBu7IO
ZmMz2eWAnN/1m1E2oXmsqQUA0zN2GKtj3lkujolXNuMLLI0hvvJluYYvxGL0
BfkDWvCcPlPLruqZO/IZBxF2ZLeQCl9hLOEVCOTp7OBJTT1TtsXf+Pz9YIo4
3ZenuNSxU7mRXFMJELlmHm19iT3Dv4/UbBvRrg8+SWRg3p2G3rHnO9sFVPvX
KZN8SrKuKsjn9bz4lAxTU+XcWhT8bETBNrRwOqjzzqcgW0odvuJm/585bTKC
34WUvf6q+niwadXHEsCcSL9euoUQoeKXuSkaEgzvTSlrV7aj4+/zhpfZNshE
ZhzFgwKtSjrfoG5Hn10pzi5bQNCxNz+VSZeiTGHstm3CWqKbhtjaTbRpqPDR
SNAR2IsgTc1IVr1CR+3T9tU1s6XnbEUeN02ZYiogNkFVLLBTJCcIxXZMNglo
qsJQig6+TTm3doC2RgxmTiNjcvmVB5n5JpSX/NWvLkAeIWzo3Kl8hD1sWNj6
6z5jgrmy1UHMBiQQZfUfD4eWV2Ce3QSm/U6G81z/MNHsXEkBd1qZmumfQa3S
aKeCQAV7PlNykdXjFJ3pT2SHVIRRU9hG4kaQN5DRcDgmOp9s7wYojehEr0Ne
LYBFsQNH48wnPLgNzr6XpfBnlbIRMSTSY7P2m/FaLAF7ig5ZMma75z04NccW
fkiScU7Q+vuDqKXZ8y5Lf6CROSw44ao8cGmW/5ujRNE2BaXK5m0RcuHlbkV7
JUYlxjwZnwjoudm7gwKJHUVwJDFVnrBbX7l3buGv5EqWJwUx39+kduk7Dm2W
0ikXR9lSQ8f/hlxVFqHaLJ79tqq5FGDzOCC5OHLJg+Z89Uwvno9R3zbhbAzV
bnUk+b5+W6jOvs2YMRRxTLUjw2EoUH82ZWkA6I8uJXSRlvxt2Ss1tqpeqEjg
QB50RoLr8KrGoDdnW9mST3eCQ6MM1ybtbeGbB6JcpuN1a497nwGxPhvI8O3Y
Ieeea79WBXLjnZq411QzQaL/8h2dhs/XtyGxAz1ePKrKJpgXOukQUvb0sMnk
vbDsWdtab9UQTqOnhDCy1l7tFik0ED8EXGavbIiTteRPD3360d+7lSGhaw0G
xQImwyvaAHz1IKRiCVzlwx21nQAqzVsVK4FHHPtbRSo/DkAq1264yz5+XyyP
2CzaTlBH4TFO9XaymYMqiXGaRfuU3yM3F9yIipeIwsHkfCTpxRWQkEdH17cZ
Rqnt6YCZggbB2gGhM8HiTEc0gynRl2KIjy9Gjr+tMpJPi2+qyjUfAoR2GCid
SgSazb8C5SJuiNstfd4eiFcziZRAG0+mZCiaUC/JE4N+WGm2elZ/7u0BKVfJ
j4DR4hfHoXSFPHa+CdpQNR1Z5353McCk7Ub1F0nprpQZadjA8qEhaSh1BANi
LBV8yGgLr4jrNxom5UdNHSLUsXHyX2FRB7WAIwG1aW5F9cbycDj0lnX5rjWr
g471P5XR7Jp7GRWHaDODQxFTgjWherKd620x6iSbKGR5BBw15UZ0ZTq/l4Lz
e2ZqZUVLD+BfHpYmqbxH2erkM/HzdQhSWI2JPNQndiO9SybzzECYRmNBzqAi
gqb9plCuEdELortBMRcCzZTdLaIKL15ZaVIwL3XYVksVTs5o2TjZ0JIKNgp8
pe64yxDV+YS/TIxJFDj8s0lHlVYFSDG3LHL2ictY6grcFi1p5UjbewuKc/ER
p25P5iofu3Q1eHk4KLZdOlDO5AhADhwNgF5OSWvsQ3JJuMgxjQXHq3kQtOGW
xW/RMqGaykTdtarrykoE+qg7/MstgdzNaQNoM4svRDWbsybNz7dk0jmAL8Wx
vAhoiq4sQV9ZnNRicFlvAzaYwmd4ri6mBjRxFSt2Rs77ZOU1hdW7mAmZ7vOx
tIU7fxy79Xctx962/NQkmzdIDztK3S6YBMFb7/tyHfPNwNm+OstkquBDKYcU
QHupTVt5RLPNu5N+CCRP4oxzhqNkeH/IGDmAOfE+D+DFMD37kmD67BaFqgh3
u2MoEYP/4i0kOpKI/mtp4nXZbNHb6Ay1gQMe3O7NFEafzJs13wojlqaGmqVa
g7U3Bxp2hwoLbde+gw4LMkpsD6g0mUuU3d2Nq0AdRf5n+XFPAMGyULbDXn67
IxT922hcK9NTCHcbD9Iemb5RyQ1Tg0o/GczE9xaR5J0m1jD4RC8954WKxGhR
7crAyRHFcmQYkqJJOEaLbLA2BEN7aWPyk79YcwCk9cCq6R00MkM9KnBoWekQ
e7BGfAqPM+5Vyagfk49/7Llv4iI104l9qtbSPr8qGmOPq2lWJMbNuv5mtG6Y
5IZnuAsi8esp8uByNPUAS3Jioc67/7KPNbRzLvv7VYnTi+rRMHrw0q9fANKr
lg54McCAz67nAfS4cMq3sv0jXaWPPHEhLDk61AJ38gf7N8nb2mILw7TG1RMu
MCWwdbdxA9YLjAA+NaELp75wP4b6YnMnGlhb9sBC9pSy2x/7jlPmbZ1niD80
ui4kFdBFAUWVrRIYoIAwcHbPkAko5Bti4kH9I13znMUlQnNYM5PT65if2166
9Pjb7/EBiuFtPJBT+r246cNJaet5LPDUqr9Q7hpZ0iaSi5Ik/NnoILQ9K6iX
nJFnrwA0qUiX9q7P6k7bJ7sDj9lm4kSw04oxUE9MeGJeRnRbu8m3PdqsGk5H
xQliFFiYt21bL9gB07582hHn//Xy6ihnoojYwg/nfLHHDwRyB0t+E/SRsH1y
HphfpPleqZlcZPlhpzCKgN6KPWgQlqWgA0ZhsQowc9PQkOYU9a5vJ3HXOO53
sWLqiU4jHBAUAeaylweO/MMqdqKDjr8e5nZJAe08voEikQo9eqBF/HoeOSv7
e2n27BTG8YWcF5AWfR5de2iwag4SLeXOlmMcq+GIZ+XY22MYwqU+PmpVphMs
8LErn8PVbNlVqPqABoh/+Tm4+JvJA7NLdXaklt1IgN6Lan/9s1RSU1G7TDB+
MaH9bPn7rf+4macGIP8wHHAZ7ZeidXRnJOpZimy2bpzutWJAzdeYRWVb8vge
ufjVBYVPEkS6iX0U9G3uxnZ8CHKsTj+QF3uCAichGlGe8mPAOssijYlfUb3I
IZcDyWffnzIBLN4XmNaCkGWSn1GNJ5r4FD5/p7FcfSyLD3dISS4JVOd/eyz0
AQC8TVgkx5YT2hilCQzalzP66QifvEQvu9xSn7LcG+qlRz7PLq9VVxEvAvPD
DlCuBnO6pIZjW8LhBFtUv08DNZdMCQZiHq30xkmwpOo2tayNUp/fBeLbbgHV
QTYO6lFNiMpqIzP45Ni4iSnva+GR7hsPFupdG7NNKLVABeWX3Zr4YpGry1b+
UY9Pc0clzXhLnxQNGT6J7lCd7lBPKrQhAFGAcITs9a9fRiKuTYk9styIhnIb
BbEGSxM/CA0oPrsO+8TJ/U/WS9PyGQ2T77l0YFHCqRngQmo4rg1PpOOIZs3l
2ePeiic8gNzziI4+UwKVioTtPfWUy884BcDyPHxamSx/Ybu3EBlYWeAtsjiG
r9O7B9XK58MHM8zeq4h0xAGeGj3M7WKwhT8PFrGneL1wavhvXQkX2p3g3ZCg
qDAiOWyNxVeuWczjCZRiCT5ROeqDJlgI4HmpQcL4lEIAuYGlighhG5gAEJlt
eN9gi1Wy+QZ3rQw9eXJ3U9dg8BC7jFmi6R4oAMA+QlvubJf0u68OoH8b98Sr
tcYDrEpWMS/8vvAxV7/h7hUZVVs4RMU+qsuf/AoOqhq8TmxLs4vA74qmQTmE
hL3Gncy89ODIsI78MeHue6R+2w5+75mKJKetzXc7Ql4zs9v1I0MIALE+tuUW
3gLeKIUTbNtzYPt7yyZhk/IlXVqmrNPjnYHJPV3LSUxlmIApwggZiAlUZWZj
8dThndYieD3BSueVHE0AozFyD86uAJXDEoyINnQwlib+S+7KvRlD352C5PL9
wX0majEu0iXdVdU3puZWesaEmbiCkhE9rNPCK6opluw/XUUFV9GFSnZfTueD
5muvrJeAh2KBVvPdUD1wCqevCJh9mCkVIAwQOr3TRmn4jfuLO3OeM40VY8IR
ReimmJsoNZRpzxksEgiWhrZt1q4hmo1BB1DaC8KHw6Te0uaEvBOdIjIkw/+G
Fn62rXGoNIwNUsJPL6IZ3nbfhPxVUWGiJa2BAGdiBkWjx6rVymoxreTwQSps
xVMUNyD3s220150KPUT58Z3s7Di+i3fqrqpeV5A/XGVIoxycSP4lYa75JpSI
bNs+ju5zwrhj/Jr3iVi//gH2G4MQLKhpdKDWDwJdwWJGmyawxnxZm/dIeMbI
8O8JsSNOlrnYyEMcKCcl4w6w3XpvNZo5ZOpsqrt/G3L19xe+sk1q9a4gshmb
MXAi7sDTcrcp4eUj3xMb9SzZ844wy2doVAIrHHnfev76b9KziNv1seY5Xz9e
yBGoh1MVc34t7UK3wPMY6W8nITdVX5WBYBaDCobkxE5KXzRvN7hOqCFqWJJ8
/Ry58kfML9gST3deYmGD1jM4cqf8U8gtTHbQsApic1+S0uULmKidVR4ykRDB
LbKz0s5WAM30PM+lh/TE1PxMcnRC6x9h4OYmeauBtAGW8PGmTHVf7IhQB3ew
xaBDjPADzm/bKD5Q0kEK5j0+1vBAGfs4Y8uYpdP3hHLITXFuZCt5rZL2KDV9
FZFqAjXeqh7Lv/sumHCJMtqhs0gxJAKd3cpi7QX3rYDUHWCHVKXnwY6lXftj
942P2lQrw2iHMIHAQ50sCkjlleYxzAXxP0Hcckm2yWz60sOEmXVGrOdfWNNk
3wKqx4qMCDUmZvsjaGfxw/LHIodqZ2zB1o4nBYqb3K/l0aoKPyvLid3oIqQS
KI0YuEDoCg41Hu/OdwwnCUJrcf+WQLol0sFCxD/pWt1Wu2L2vg/XNPF1lnn+
C3wnS4xM7SEUNEoP5SQ0BVf8Q3mJTxLpy8p4UmCeN2OMmnvgI2mLUI0zsn8l
idF2nwZW2QTcegpFvML+h7ZbeN4dCOeP0xIWNQ2nrIvthygns1t0xQHO9ZfJ
URZ+sxe32E+UYsfdz+VImpuv2x0BDCz5Q7XstKfeM9kSCRRdd7DfeavUtWgi
9UzvsWf4k83SwmHdR21FUjH2l7PghdH5Ud2eS9jOJUuIwTLgU6xtixZZfcCQ
THdZYHBcnL9jiLpspdlDDcUeBXbV5Ggp4yabtYMldZIVSNtrxnJZCJ5B21a1
jLFsql3zGiPIIEW4y6+AUeZ0dINOf3VcOGupQCU8uD02iqyiEAdq7mUHV4Rw
ZwuAwFNGjYTG6T5FdFKPcO5UfD5rHCgHLmNn1FklZA0MxPcibDEbQW6efnZd
XMgBxVKyBWca4Q8a4pjdQTtgbbQsffyyfNy5uC74iOnx/WFOb2OSlPB87gZg
8Wkigtuxv7Ns4pcR2SL1VJhN/kfPGbt4PptLyGpijHAG8esMimt2QjxLp2tw
ouRESmqN91T9Ss4PfwqdLApkFrRqSOzszw7Zt0iWC2P3uoP8trb3fUWMpBko
/GUsaT8r6GJMTVvxPUcTUb1PWkDsMm1a/8wR6KbnoTjrCcdoA4LJ6huf6wKk
nMrO/i9NUU0CwIs4FekClnoEY5nuft5UHLVj4Oy+A3kloYjtFmfNeee9hK4U
esPCd4EXASUYaXExFsMl4LKdSabpmX6sajlIUaY0+QGjmeZNv1IhMeWhembK
mtWedMl/zNkRQUrWm3rTBCTaF9aRBEf4b6hBN529A8pI8XSH19FQOiC+xVnP
MQceBd+cqbm2WCtluUnnRwRG9XYuGhKV9E5gkWFR/4nTuwTqZNDe5AUilfIt
+4G2z2IsgPMxAtv2QgTLE48fOpBVyQF/fMQXB8YNn6KaJ1KaphMiZtqUTV1K
wi+DwQTmMc3iIyXRQu4rbQChXgdOqUpzMeXJk8BFogPx5/jWIoHQkWH8anoN
zQ0YXZRZcQM5foNtdZdDMF9rleE8oOuAwXdDHJQbb7jVr+DopNqPr/1rh+hA
mKAsRqAk5ihkOMlmGJBIdQ676lmC0CG0tV6DjfHz1B/4Gcw4edlfuHFRQav4
y49djlaUi65XZachjCNXCcBrcwliTU7lUbLBnMHjfHcUChOU+K/ib33nPBqK
rdrZZEb797jYZAedrCucglyADbZcZWeTwvhEWlOFRe09DgCfi207cC/bZUS+
VdbjjZ0wynu7NEGChgi+CP//iSv43S2Oz6aTf2wZ29a/RCg2q0+XZ/yafsM7
MQqipEvZIvD5Y92r8gfxktVNQCFMPoS1KLIW9qL9MjcijjNWwzwJ3pscAGdU
39liELo+vLTiB/qPGhWadbY07t6CD8F1Tue9NUTN9qG8w47stUpIEOJMuxl/
xDNwxuF7+uAqGrypxHQO/Q5l6rFpC8Qg/gCjOPNDwrHQyKH/JUDhOtZYDHR+
72ovqWuFgfspbN0c40xukqE0CDRoOnKYknZbFnYo4onVzlhT3wznWqwQWH6i
l6DMXq4he5zmUQnyR5f6JfCvYjvDc0gFU31Zi7cOgdyIReK0tAU8ym/XdRQl
dZiEEVhwu3l5B3ilQxBRp7F90wYrrRkx+N9JRpot6Kebvm3wjcygea2q2zZc
lu2mbPepBVa51wmLR3+niAHHmGjy+3q8Ytj9idPU+x5xKl2EZdwrB28z6735
B/PSXnKCwatpUKZz8kMMhLTiS7BeFS0sxOSIQOX0MtWi95B74/87jm5/M5P9
Jp5BEbWZZ71e+lSFBDOcwfnhzFOdn8CujuLzmQbyn8R5y1V7R8Q9F1niK5OH
80//2dNulsvqLKyp0Q+xM76HtBUSe7L6NyK9Z3PHiKO7vjxsAbVE9B+ZIx7Y
2rHZhex8K5wtxJH2ns7Ge/jNEXBX+Bm236RdlFg43QjwHhTWiSngLD+QUgj4
WbBpu/GigdwSpw7RRR96D7k6IdHrBUB7j+nRDcb/i5Z+aacWwYKKIlgIbdl+
VcSE26t53YtRmvkFp9QjHT0Lkr3A6C00UeNmzLFbXYm07ogFn9WRzEIXFn3D
EtTugVRuce3MU9aTX0BhZdsINgx8sfXboYpNNlFjtmzzbAianqumAQUQ8WP9
6oyvNcoLd3A3mCQvReitqVB0o4yYqGVpAZSKCAJ9p30791zc8GMEXg7I6Q1G
djk9q8KHgZS4l3PpT8jEC99c4aRZcD6+99cN34ChDgXFcAqz1Eu7Uh+tDm6Q
oqIay+X0F6PBoPcjCde/4Ua3/3pM1cPjhFfDSTIIw7R4Xf5kUehyjSNDhm2D
dTXJCCmVFXWlzonHAZ4F8FFFZBAHH6LEMxUqqy7J/9WZL5pLih6DqG/kXE3Z
/BcddKFL8V9cUmGk6KNbiz6AvxcCuLHfOaVReY+W6CWTIT3aNi3+8H1VyeSV
j76GMBdjC3zzAyprXsh/xDsiHi1t+U+77EBsFYYmQyGfmYjdSZ9rygo90Szw
BaM3kplmRjJDovI1zMW8Agfj+lwN21nTOJcYEku9I6+NpIvNV53kldkKZY+X
O4n+TAVOXrqALhxn4yxwu/sgUl6RCbjbteSxHoYP6Oz2yeT86BKhYP9hJiOb
8+v+YAy+xyWJcepflUv+h7d/8p/aR+3bFuwLKCWII7VHmT2CSIyuHYNmy489
FVvYdulFckpv6tALWSUdkN+iRPBWayUp3Sma9Bo0UgBilPODAZBpylsXG1qI
0/3WtFpsyXdEzQKwp1Lnirqf7+DAi6jYc3znviz5etLaRjH54EssAjYEC/JL
pYXqDM2E6Jx8c2yl1mYk01sfPQqnHEfnCbe7rliazVvOhAGncCKZFLEixmO7
dsFPMJaunAm1WnIs+a/Tq7xK/FtpP9hRxcZfiZN1EhmCLHw537x104wQAdRc
TazQJzuzScsqUBXFz+lB+iTILWrrxcy2GTLKtTTWRQKufrqq26ySfmKwfhvf
aaupknnAi8GtMk0hzN6cAb4T+5irfwv+N7YO2jC9ig7Wt+CsizcgfMNV8Oeb
2Zb95BCa+Gj+Own48dB4q867JPF68Y44/awNigYc7r5vdk7Op9Fj9xK9kDZm
/agD1l4BBez8wn4WKjpzN2fu4jkRSP12g35YYlFYk0ARJYgV50+hRj5v0aLz
SYRvh6d7775nqDFMbjnq+v2VEokke7fkwBZs1XYdKexceIZE0RyXsjGl27Zi
X1zAxi5GXXPM8CWRyK5OKB7eXgjbkzgh0auOVQqWVmYKZgWOpWroumD8On3W
11rd31Wr/2xPxV4NgmIu0U+WtcYBverVwMeNrG6GuQQDpNbaMX7JOOpjGH/Z
GOTMXWp1dS5p5a9fmkOKerzt/VBtAWJDT53RRHXy1ovvYNwdcZlDS24d/HEg
5MUtnF3B+n3oJhx4peuNCVtaoO6K9owM+GCCiitTS/lhjmaOPlOBCBJtj6mI
9y6JWSFqnN4FbzG9l2vWvjo0f3th5PKtIbtOInoSbuYKgAf0LoWoz4viiRZx
1D8lBx5Ip6zpszb3BITXbBejWkeihOWrFwGsxuyD+RFSvAUNsakbV4vEVLAL
jSsqqBueqFTCzYfC52zop49Y0mTSj4aky+Upd6aLLDJ1uAPA8Xk94Z9QQW49
IoHlxmklfD0ZUKY+BbbSeTAQOwvxsO0SfinmREeomhyrdNLco5fVai+YRxp2
L4Z+IHbUZ7Q2QGDI099SX4xLrH9ZkIwlN98w3l7z43XU3MjjoPb2ZBv3KF9p
MAiyfsNju/xlLS0vgHcxgmMxY5mSsukIfS5wAsHMvFZn0VLi0Z8RIoaJX9an
PmVWx323FXpFFMZDVRdqIESyCMFk9e3MZZQrAvKdoR0QzDpklDyW/3852bup
3LCPz8fbdhc5VOJjY5rVkPGHDJ3NIjg1wYg//vLX180XMrY3qBt4QEpHYfdu
b7lOruGYchh6Mmb6VmZFOB/6OzQoUy+p9qfhRs6RbY+PQVxgSSJBZYWm8C0d
agjqkJ+PgtgNEwGhq/xBpgknXkUJdH7+ZHX38hkJ1UtkFo8O590SwQD48vyw
6ZlGMOYmWqPJcUQxQUBmYdYhEVuaFLbndsSamE7D8w25/ruYgucMEO4ovC9p
nE7M9+u6Hme8/5XmEKm9p1BqH4D7tImSP52mpRhnAWCCiDNvVoBXtPtHbdcO
dWcfcaWBCS++OAfvVuwJFekoYo6v2S0vBTDK3XmCwYq9d/8kqXxlxqJOWVuG
+v1jtqINOF3aNIrWMW1TPTLWhFaB3zH4Cs3/I2jUYRoUwYj3wqcwOA5KTCQD
tDBSjCCDMdrsq298yCJ4IKIrRPYeEf0bIzTiu33j+km5GviGS1K5GrrshTs4
hdFduL6rgXNKEYTOGXoR8OR9QdC8N7L7mKM9DtXVMb6qsGakTFyOZAhnZCxU
C7xSWQAkP9W7h+DcFP5S2QhpD63yXXte9kj9v6kktm7SV5nies+OHG6TJxMO
ZpT+mgXS72GGbAQGE2C2PKTK9GtR4MZrIDv8u78Z9WACGAIMkm4KRbq4MAHF
sZyeBbSB2kDkywKVxlUK3g/D2bFDXnw7YnoiNUIeNUkTp9SGM4h6RtvGP7Kc
xNgm1l4DmjnauYhr3qGoZqjQXL1i7m2deEQr4qXMz96TpSXLKckMaBZ9tjae
tnCwDQgVlZt46Md4+h9iT/rnm13NTRrx8PeiAakVlqDuTZ9amADQ+R6oEoGG
SKZT7/Zv+vqeo5Y3QjZ9TZvv1Fd3McZHSG/J+nB0ce5282UApb8Zh3hcn5q8
JVh3Ps4LzWJfJeLxJCZ4B0KpjpkpYd0G+18NbsEsIz9n18FOCqkdnHm32ZoI
aFs2TP7IRQzEPLK6SLUX+8FB4881KwYahiE3h0+lB/fbwnu9JRY1hYGzd9+m
dUCVCT+Ll7Lr7jSguQWa5Mb+eu6Upkfv+ZX515+s5uJAGhC262o6louEq/wg
JvzGBNd0OzCom10xzQ+ioWSdhIdGqKuTxtQwOAyWwf8eskdNw8VREv/r0Yey
o1XZX4C/NENjpqQRC5PPzvPx/cch4aeUWCyMNE8Zk3L/JLIU4b5sq2YzDYey
pZ2VZgI5qIPDW7zUreLAHjtc0YMl4RDSZCib3/eZlja1Gh/MBrhHdXqWqs+Z
wilrgBsGKEMgvn8l/wjvJzAjn5+Q/wFBcZi4VJYoiM3DNu3qcjUIBA0oT4Kg
lw5kh2Zg6L+yqXCTd/2rQ342a5GVaAVhiSo+Ba09tRfmmHYh0EqsZ4GNj2eF
LPen9hWxDHvsJg4VY7hKXd+JV8QYR4dO2QkWD2H9j1mL9udKIQX6oyP1RzuT
gpgNojLWRtSYsLAs+gAa9DOqt5Q87qcMGpp01YW5882KKyY6RnAJ6kpUmZTX
wiFXrnqXHjYqVHT6RHaBwQC8fCIiJ5Kn69WfYZ6ZAPDW02Wt0HdsJtfgYab/
xNZETmZoQhdhZ5VFs/TLCdDUupLtxhutghjHwZ7MBsERSstYT253HZCu4ko4
Q9OkaEubOzYpg/YiNm3KNxk5hzibPhTheql4diz7gTUVQp+Mzg3R8F/hWkfX
Qcxo5xVzc7hu92m2aformKPkaSY4rbn3z+kY7WmIi2mjjjWHIswuZoq9/UsO
PbCwYElLM2VKN1VOtuxdGfnoALvs9DkwJ2qOitfswj4gwm4vtpl4yoPrmrpu
F9ih8FU9O3/mGjHe1iWN4ZleBgdnRLRcqkrStlI9XVV9746bJGhGm2OQMICQ
obB0lCLK1/tNX+1NGKjf7/J+AQuTaFdIrsZKIDpqp7Tb8GcCyi9+AbXpiE4J
bOWu0fOm6DGIrjS3Uiixvp7VufzrUjuWRZzt7lVK1yNRu2spZ2CaXUHQ5eSZ
WwY5L4o6VYNbANRcuRUq9w0m2HoQ5ucdGDWclrXE5PbV9vWbn+uedHEd9O3p
poAy/pW/7h24OBrW4FfDSXfu0fXobzoQz7A4GoGx8TaJTTmgBBKGTnKzmbrJ
XHY4AqZayum+gmXgjBFD2u5PJ1GHsCWv3wIGtrCTUvq48ac1AlvhGQiN/7NN
mrdI1kmOEPTR0I83h08oVVd39CTxMPLKxuXCGLy6WEh2j6ObdNwKcNG4WXmC
9igS+rP+PXVo3m/wYW8B5X/25LokDmXB8kecIG4ZHCXV+sym4A2L0Lh3gP9e
ddNAyna435vUIVpwCGMHmtzInNc2YyBZTxMsZGCWVTO0JfK82nyNxY0/b5X1
MlfA/Sw+Y25/iQW85cBz0tlo2cydvxw+9UTgAx97iP+4mj+c44FB/vM8Crug
PTiOIHcWvFOgCFhSIow0ccNqE9NAPIPgESjj8uIt65Gqr0cqWWXjr2MSTiVn
0rUfy4Sl5/MHiOxp75LNOO7iSA/YjyDhjAJ1sbaqkiHH1TEJ0ZvR7AkxhfuC
/0ztucrHwrt8WcN0Sm6EJx+fQxAGcoO8OCtEeDKQO/zxSfpaO6JrC3Als78h
BKFpT0v2pERMwSmodurnIw3fLNnw0Qudkho0kbHPQyluOLMFBPf5M/Y9iRrO
lyTJb5I6VXJ6JxOTmm8eN8IRIi15WziWN5F2y3m9TsuwouVQBRTXgdUyxqAU
HPmS3SXnuGd8rDB+D9CXlx4/yB0jtHwEJu0AvqQtvq3zyR3b0Fjqeb1704+c
GlwX5SKTTAucp4+Z1oER5hRKg3kK0FTOMlaXDiamrxjp3bTcsjytcSsMBQSI
GKB573hBmWBB8ZR3BPdJzawbHmTDpwdIL85OfFGZEkzQep3RW/SZ760tEiwM
9lWjLSxSYqJcqmKKmMVFd1lOcs4UE6JBmxWZFyGvWsQf18nrSfwFtR6nWn/v
g3XUMkaiDSAIOyjg6veAOhHJ8X4crU01DeJnR00SkF1+xpXIh1mca6lfT4vN
oZrOymln3ts93GynsujMh5m13tvY6VdagVZHbgr7jU78uCA48nXirP9HC8+y
TSubyqp4eu3QsjnWkDI5gZSR3OJUn6mkoMfPvuqQBWsNwao6GqeXUohCm5qN
bkgX+61/zhUPG3QfCyU98wsCa9cDCWVQqcI1yJi+dSkQYPTUPX3KqR/ZCMBe
FI0zjtjBSUtnwOrRuQPoN/Amtju/40uGY7hGTur2rOrkvvPNUdrvLV3Vadro
dNODcXW6dOtm361QhZlu0ucy0EyrfBcAqSK8T6iXQVQSVeHc/AeSk4NUxML1
dXgNQJfPKrVmUPExw269Co+TlYtOlYKnvd/DyNJpDmOLJCo4XHz+BEoWh+7b
y5LS372djEazQaWQ2EComE8nNnUCkfmAMufXdraWHZ6PCnn04pIUTKePgxA0
3hV5xpdxG36pmNw2V4g6/pAxvA9X/tmXozivey57eXjFp9X9TyssNaQQw1mG
WQLofcpO5CdhPHgipqyL7e9PIkvyDo6Tlxl0nL/JQUL+xTWIiRxTutWq/46F
wYfAj46EuVuFtFm9nkybb9qaY0kxwKUPSP12zDDj60hyGHlIdL+n1On/OqRf
ladheLim4WOOkDQqprzjeX26g0e4hAWSBxv01WW3PNCc1AKf+cT0VRjtleDs
tUeycbyXzn1x6ifYJ07HhrueokNe6HjHX8AujdLhjVeDmO9FkdxiNgieCwiv
cha0SsFFcUZAGNUZ/Yu2eRLv2CKzgho+jQp3mz5iAzxa3l2WUDVwXXDDXOxe
YrHU0KljVEvNEj5IyxiaZmoUEYdnycYvL8+qV7DMje2qMjU9E6UAFbOM2SfF
mpvDBwF/9bKWuLR88qgFwmFEZN/wcja9V1k1BvwhoTK12t08gy6ePy5J72eP
ShBi/YeQWzrU3SITu07vqf2x5m50Z4l9j09BVbigualR9ygmlu/Y+q4cT4gu
aCAtsuCHqs/OifH2Rn9Yl/RJjB/wgVJ7DCOg0MSfs5znW0t5R+La8tBjJeif
payooXJV/ZDPF50eQX+UtAhj4+/wEftgoHSMs5lPqFfqR7WZmOevtpurxKjC
Q64Unn3ZYU07vFGU0+FyViB18RxaXQy8TgM22hcuIhQBdL0MbOoAPbm4Q2QJ
SOVie5oh9L8gXDe+kBKPiy2dmHibfPjWZ+duzJUhrYU50RiID0QZ8BR5/4dm
8ILjHGpPj8JCl8yoZJtYIdoA76cblfbV4H43pM0kV8gUxyNE55AmmmQHPV8y
ePxVA+zmpm/Ru84yogL6uDfKqjh6lCEfQLto0gRf7WGrG8QDE20lw2I/3v3n
LZpeZU8EPWp7bJHpwzVX4eSJoisgDnq5ACgz+fxBPkav3443w4hhhHCyfacE
o94qQklomIeBBiS7QA68S0Vw7xFP5g4VqwfU1JvqxZ5gy7ZdVhaGjPDE8gYi
PRY3c1dkAdys/H3FRjvyoTcbwqe9kKw9SBte38GzUXPTp9oFonkJQKQGb41q
jQUkG64gj61zHclz5nVU2qEX/1Y9eu4EmTaQOBOFj8kQgYAAOYB96dIB83Pf
XvzeR1sKvJt8Dpv3jGQWjhGywpClVUi2RDWaBMC5/1PCedOZ6ZgoKi5eGlyD
PTxJFgSVDpEkWQE2XHcpIAePQfAxCux5nI5epU8Jt3Efapkmb4Sez17R57Ld
i47i5/DhFYAOh3IRi0J5vGWE7/y8s5MfuObW8EIsf/eowdO7ssGo/v/qjch2
JpbcIfcwc2Oadq5wR8IdYh5JrcNIuy2QsicG14tdbN3EKpcXeyt5OdW/ursO
luGaaQfh+XP49nNwzGVcsYdiSk5v4y7efJfsea1KowZi22mUYNLuIGYe20k4
jHxl2hgvaYumLHOY7pQ/3rFbf6OtF+gvAIFqiR9WteYJTfga2C4VlW8Yh6D9
RdLFfeEHwZPUZr7fMJJjNAFIoGyiv0KKOFAEn9Kd8GssQfeeHzGubhO8XbIi
h1ULo+nHjiZD0hs9rsaeoR8x9Ks7tWy22ntKxLzZRZ+mOsFGDFFrJg+E9bwC
IMWYYuhTdV+df42ngClWI/XdihIhu3Jv3oXKyU0VoY0MdtqvjEa6nx9RoFCZ
1bumUeBA9R6RqH/1yJV5F70YXX1KiVuAkRp9fc4wH1zdnmY257NRYHI9hfkc
97/GvxQGU/GGdTuQcpADAshm0RQ1RllWn7yGcyFlCxBpKnNsivFo8aNWiMJu
bRcEQb85NJoBaDUWdJOc3rPS1RvWOIGagNgr4W7NaZ3jgDQevEA3Ihc7l34t
7Y1+OSk/pgy2xDt3+ASUNKxT+bBFE9cJPU+nU7OHmjYzAhzcE3GuOT3SC4Jd
f2X4Ul8bUy78wKoKiPQCwRnUptWaPHXG9ktkGFskQeOZW1HwzO31b0vmOJpE
+PRPzfr23C1Q+6vy2jFySaUMN6rJrP8L1TYIasU0bUVds9cAcBg6sqImOTfB
e3coOjgMoARjRhivaGyNdToVVCG+hOLTOc+86zu/6d+ozQZHbfBPVWvk3O92
tE2+lEcXD1X7XFbyQrm8Xtyn0LtMj8LsyHkl1xhLJoipEPbK69YWPZHTZ630
rapavWFH88F0a0qbsOMd+nnHdHMh2f8g4BRfbRgeAoQxwq5FxIDUrF0zCNXk
PSnvRK8iQrEBrvNKkdJ13cTKJzWxjZsDZE/nZJjlcITppKnpsL531yzZin/N
agGtq/24MjJgE1FlcZldV6upAPZif2LjnSBPfalUX3pdFzxMQFjCWiSmb/J0
m6y3b2asKse1OSM5o5Ohdw1gqDcughJsg8vstbnbc/HYKRSko6Lc5dLLWDcl
rKU+/6sNqO1t2ZYZwII9Kt1zALPjbBRB3Itl+bLuoeS9m6knWErgjRrN3aMv
3tHT57SuLxkIJU3SjYPp0CwPT8TK5Ln4y4jUZTmUMQVxepoxv6EstMn/nLxQ
53f/BLF0f+4DX66STye3vTB0qvSDinyUHOy6G3uzAh7NCHbBFGa0rTiPigyY
9mOAmD97uyEg9Nhzy6QefbYIMqUf2s3ztjPTYjKSAozz1bIo9b4RxEzU/5Ug
g267sKfS2xQ1j5LHK5PRyi4FBCUwEATeu7ITT9cw2064cSbuh/QAa9VF3H7k
AWqSg0NLnqqLUWCqO+FGcdGBy6ARHVMIUsqFgOCOvSXM2VqbWmNSqs7hzn08
m0yKO5YJNeWz9dVB2SG5Xutu7qsAwSUfpjReKE1XbVwZkNuY03o03M4jGKow
f/USt8JZPwvbTNFLk9QmHrhJCtVGuKcnFrLxIYixXmv1p6TscJmlpMWgJy74
D5/RrRRFQw4776GgeRUyM3pOeQ0wuzzCtyZb4wh7q4yxaOLOHijnBjkfkfv2
dJSU7gbBUxp9at6YaN6RjN/TaUCd4/k6vCTEUpCOpZbO0slT7VlfJtQhY20+
uFgI5sRdlz6PM03noppOTfuHjNA3MwK3lNxtviPNgrkh9SNmLUD7rkUtg0VB
9AviJGWyVeQ1jMHjVXZHe92xgQHg3rkaAS6P4xlmyIx1/85JFHTHi6gLZ3m5
+dRxA+yEBmviEUCxTBqrh0eQDrmDt42H779hLyUz6orsq2Muki7uwz6ycu8n
mrgYz/o7xoK7x5IXoWK+skz+b8FzR9SvDJoBoYWCY1WSvWR/SWaCXOSq83jQ
CK/XbkhEWI1UnkxuZk4a5ZOA+784S0rCjww7ROnWWY7ZTl+fDh20DlZ/SMy1
Tlcki0UTdGwsEUWpH3Dxdv5Urzd/fBr1dZdaXEeEyOUS3lcb/rDYAIgYq3uX
BUSW2GsOKdWr2jQpR40G9sxWU4cqwqkUnXCOTNvrE7pr9yGAFpjbXjGnKG9W
oIjSXd36/NeCAs5gvexHij05ya1n5RocPTKtSb7IEafI3aGgqJFVmC3LFVPe
aiIhCR6jm/dw4GWBaflO9ebPEicEe1WDJFVc/0Q1kTuXJ4uuv2SSHkAGtERi
UjiqvX/yPkptIk072mi/wdOAb78Za/qenLqxoftKFnamV9NmhLJ+BdNNmf8v
Rj+6QzjXnlW97erhYfSfJAADZJiVbpAPL7wx9J5PT59mYJU+zS6Vh31pATWn
T3Lyi745AE+oDIdyPTygNEAU7ESvGmLWUFfh6zjIO4gyrGGw4oyVNlpLmOzc
gpfO3GgEw2yOWaMPQAqUYHBvmJg7ufgngA5WL+t2JVazLagwYIfeoiaPV0zd
R0CDZ7vsg2BTaUiVxPj8HCTUGxZVpwW0Tl4BWDqjKHmbUzznJ/+PqQ8pTpwa
0b0GXEKhLQyD9/Rxej45edLcGE1uVKjsbE42SO1UvhbKlK6hfKOBUnHqgXtG
AwbrmtMEDFYPvbYYouwaGrIp9dpkPEM9r5pBUxkrU9YxuZ1F+gEhNuoOuaiT
iZvS2fE6PtlvJgOLTsCkL0vihpdotKUy/hiapWMkRh8E4VD2tbmsSGyfhdBd
Q0DHbA8TiDWe5FQHWTwRWq3dP4YCVI3FxZTkP3hLHLk9+aWZzadNeueXzVdh
N28J840/s/WIQ2XtIru7Gi4x1m4kYWhJ8ggWM4PH452WoLOBxuwBzSeUymz+
YbDSxyPZQuwwDVhi97rbPyEyS6d1fiYT8/ym82yEYtr+S5WLyy7tbQ0iRThN
vExRUmYJSTptIwKlpjsLEIcDe9u6C3Q4YrhlZ+QJHX2RjHfLtGF6gBQMSPD1
6TaZYLCiZ9TErmGvlLcTQpFh6GEdG+hn+wkHTaAgtLKQTYYJV3PCPhRv203b
wOO8cdXFymSRMZsiQrXeLiypeScNFUDzE0WIFfuqI4QhQuI/g6LtCcxZf8W8
Xlf7uDewB3/8RHfE0bz5Dcg7Unya9CyLci2RRaJHhxL30ILH7Mk+RyEynrEz
PNYvhtTPXXKn5Y1xFqZZOAtrx4DNjRVmlBquhEfLfhHMAJc4DSSOad+4W+u9
xP/kjlsqEed0aErFHPArzjFw5MpgDLrsepmaVi/VR7QqKCWvONpriF/RX0Ly
ZiBpq8qm6iNHaO7bWDX13KYrAU8GnMDBeuzEQAgOycaroI2eCYUfzaCj91Vj
Ln5Owit8waSX28AEuqqj1OUvWVm2psZX4JwGv199feeugjgXSyCevJhGSwb8
VYA92dMvtaj0zYPRgYBGnBYB0lmyszToNdo4O2KTbqLBL12+UBsPadsJYYIM
hehGkc67nj/fJoILsZ0FeDBjzCQM07k9gF70Fk9UaQkxLb2a1R6IOgF3RBzz
nGNI8trLHo4ty592VlryPGjwKmEFfJpDCCNfvMI1rw4JPtPicKYvSwOiysio
18YcTlDy0WPJC61hGNSy1K0jf6nd7eJ8jMu665iw8KnvM/yKZGHtmFevXD0n
OjosJXliBI+wgsjG1nm43wPQyuEs8HO7JGUzjAqmjxhi53aAxmOrMtE2WGLY
xiEXrXMi5CUszqYVJh8cakvFZolzHByF/2f0JRXGTRMwgfT4ZX3Hlh5UDJeJ
u0BzaLhdHyl9KJAHNOHZlEBdij33ue+AqWb2EDb9A7btam9zvtk+unyVOEHo
YYAGLoayq6DR90FdgoPyrARNVbXacBXyuLjD08BdfMC4NqwR5ukoCXYjimGF
vOjLVRp54I8DMYuLEpNnElp9zgPqOKtkNYGjXjb9t3Ndhzlo1qurYMxRWagy
8CgJTgCSa9I10WNCvq7pKSOHjeHbRB0FF6aM8KlcqzTulQUz97Gtv9KaXoRe
I8fdQ7fRr1rw1Re021jNiYJfdM+OvjEs9s78ewrFak0aQKFaWDiLK5UB69ET
/HyEzUBVTnDAqlq0mB0naKniZ+LykSglbp7yRmkAcV7OcBo1tqMV5bxdwZ/W
M3NMIQ7X8OwAK0gKIsxnmnckxb3wY/tZq3kQ50rQcPbWvyBkCD+XGduVMGif
q84fhSmoGDq/Nc+g2n5QznldPXPfp9DDZ7YRZ3FpyIuwvQcHJBjTmEZMZgT9
F0hWfFajbk2lSw1guhauScrlOXOOEWQf5A1xdF+a1isGK5W0xSVXcAIheOy5
gr54FFpC5f69tR3hEsuaZQEaphFLCO0clWpsEg8HTTmWsZrtkiBPYqtEONJX
Rm4GythdPYPxhg5i+/9D1U3FW5Fet3zK49akKQaPYJjpGEK24oYlQ/w4B5P/
PPWGTwggX12gNB7Lh4yWsohPf4Bqk8BVb9DoV80qQcPFWnYcFEfn1j7Iudip
b0e71LQrhey0GfIA5YA/V5NSokGiL3xcWlxGqyVUEjqRPQ9thKHXQxpd5htg
jj8Eu6uvgSk/DViDYFI4y/tY+vL/3IkZl6AJNrKUYh3Cm+gMeNLSyby9n1am
J8Gt1sXLGQRoxmeP5psXZhraau2zErQg5KtcgYytuKaUqIX4g5NcYwew66TP
FLfgi5u+8bF3Wbugzt1sph0g7ZATss8maW5k8vH3ZJIqnEhgtC7plIBjRYAv
iUhvdTHMxruNfP6RYGeE6wmH6goVnw9UvDtgQjVDpjdR9bCCj6XTUEpWBJuF
7wFlzXuVyA8U3+ySTQo6eowLJ+KmXvruA59ueF8M3IU3A6auI0oo+lwROivd
r6d8hgOZUThA6ErzMPTvqkCLoROXBu/KbvAZ5s3vjfCFSqSpY2x4cvovNqV/
7Ekv2UL4gwR20aQtXH//fdLigZhWY4ZNUk0EA6gg8NV5WWWt80WVjSpUDqzP
/TJ5betBhoK08O2ahRDEv61uKNCINl/akHJhamfzgUKY4NXC7PcuBBj4xq/h
kVhIjStbS+26oTzqUMG0D3kh/iv8SjiDK1w+wfrk1KjF8EeekJhAX7rMcBR0
EIYZXbSX7mCcfu7DQ171NvqVo0/sYmje5q92n7DEhlNwWgXAhqjw2NOoKd5J
YjK1dFJphNvPK7tjphMsQNuUDBPOiaov/BKpW+LBuGEj4Y2mMz1BmvPcW01w
lI1Pnb+/dCY0XkRcagj7kKO+JirOTYlzs0tOaOCqJc6lzF/5Yv9fK5h5ypHA
uIrvbSQatlIPFPl6AhIB+FQXP1gd12Wx2Z8uCLW1oMf2/UZ3cbOFVuygxQfP
xQknkQpqEbHiKopO12EcmYRV9GaH93elYuYJoD9olSvQSnBDl8z0AkybmJsF
8z7DaANOfmsgr+MB6XgXlj+wtfO54TjUgaGfbuYS67IPW4FXucv/Esoq4MrZ
KptkcfrZVBPvvu6VsaL8XvUPNxE+aKgHxs76hR+2zAB5NSGwtGKtmLNazqyf
oYH4/bErCYRqtwXwph5ZqGFjhafyVCrC0OGMEzd5f5FeUzcDOS2NM/stP+Yc
JV9GPo5EKF+qnC/GJlqWQ1A6tAAlto4VJOJk51CKrxzxMcoJFFz9djJOVbUo
joJYnZ4pvfd0/2W7I+ol3d1epgpYa4wIQXhH2hNNislq0d8DlzxAE9uX7iAv
U7xMNFiZNcGOXAG1/Z2Vk3e4rZn0pBRBiUn9kcFxAEW6hnpzf4+Xn6DuqRMS
KyEYxmUmII68IVHTOLEw2fIfM5w6cLZfTrrjFDOpyvgyt0YawX9W7HuxWcIo
EhsxqOcLoioYFOsBM5JOZvARcdRAQGFS/7k6skIz0gZD79slN4hrhUiVtKFK
4XX57xHEwGzw2fBcdVAk+MfSIXOCkmXiIn26Z9iXyqsL9MnfCvnCHiXWYGfu
08Y0kBYWTgYEUs6k7UBc0Iyc4x0akOmLNsQVygTfRuSInRZdTQljpV3E+2AY
/FIGopr+TYH4T8nrkuJfwGNJ80B8G2nsDE5054ssEQexCKJuJJX4L0Ak32Jf
lcMZBQLIQJ06crfJtFnVlTZNS88NMvRM9LdVb+cjLt1LZhOGk/A1Fszh2UR8
yE/fZfI0+7g45rHzV3nbWVljCydi9mRDVVC65i5YStyEHCz1hjSMA3Y6FBMW
ZO0SpP1FXLIexj8A3FwLPivkAFVk6jR9AGM2jSePCaRjZGva6fZfSJsTT8Xs
Bo49A4GY3YFZU//0Cx+zECy/Uk3uSqvKaSbMJEHBI+aIcd/aht49WGnGlrqN
gGftFb0LQ3VOp6LppcB8M24YTuyHvR5sBTOuROGET3M5FEbjCmmJQsOJ5346
ebUoAA6YP+FAN++DGo2S1NfEjFIeOLkbEnQAQRDGtvY4ta/0Ui3oW+EmcDTQ
Zwm8jLXuo48AR8jYx9fJdmK98VWPHKQM/9WnrWasZxyS+o0evWAB4ItkcIvu
ZI1MDi+aAQYINHRJpdJEKnlvHl/2U6KitDi5Ze0fIxiYLJfoTZ+yXIXqtnCy
ESFiEZE5cxJVFplqNfngYyxU2TrOz2r3DVFHL/UN77OyJdfzwN/RkTUZi5ik
zpuCpocNA+vjqg+twnItFaH8hrRrAMDit7rNGIhTvuV0DCQscnFM/rcOB2R8
V+/TyPzXYfAJ+y5MpqLkBpTQPAqd/mBFk7MTlrM4mjGiDm7NPxYnMUqSt6aB
6WVai/2lNsOOQAuLcItSu96yzUHTUn5YpwG9qF7qmTvYs09rNHtLYG/dkO86
lcNUfqrZUsdttdl3+Ov+U/a7G09tuH9UD0EJNhVEdHlRJNwMvtqd0xFwI5/G
JTc1YXIyNVdghQzBzq7CzcTFUR9YA1pZ3RWgfexFaJYzFyLEO4nG7R1m6BUV
whZ/4U+y2cpRke7uoUfjJg+DJTcoJ5y763kNBCCGEBJr3BMRCV2DCJ6PuaGo
ykvhYmt/uA6tyP8xKNK+qZTEe4PLJwZ27DqxCJ58eClufAqz2l4xj04UrpvN
bgvN7m3UOq4ADKqWGufe1XHIQpO7c6YToQxWhKnnUyG6xl3iH7x+yRpDOKTA
kKQzutzy6Wd0ShJyl+0A0UWwLMbE0chy1/Z2vgR5TvBCG2mXTxCY7qjDsqOG
jqnvQ+/LIkO1U2FHPLwGuQqF8yeEpm+QUPMSeVDhEAaD+WSBnz3EKytWam7m
oYNv7idTSt/FRH3rwaEzvK/ZrKIPjUNq6jUYrQF4zsEfoNwyNe1wHsD9c4Ag
v8MTuSJhTk7cg0Vzyw5p+fTkCuzG6rSTp/AjfHQDl8bqhSyBxjHEMRqZZviZ
9uEyKi5Vs2Nb1Jn97l6vI8B2NT+yrNCtHK0yQzL/bRfaLOx9lug/1sobvfu0
S/EeRfE2uqldfQZY1SbKX/0ZwlMa2u7ZgSfRQjf7q4x6np1qzakaV1pyfEib
gEjBFXnG5Q/GGRxG3OLOKESjaGIKtA6TW3QfEnLgmBPpyxtt98oBynrdOVys
ctK2woUUYWQjy0R+vnkwiq5ZH1A7+EdAB0GyArmfKHD+k2RqHCAEURLVojsW
M3zjht0M/MzRsUEk4Ln+XNtw6Z8jM7cbDbWXLg9lpj+TyE229EpGF8iNswM0
EG/KpC4Uywdp1K8jOWxbOGLXN7mC4et7Kc95w4LkrUZtyKX+FgH6nv3DPKHk
f/xojzBQ7i+q8XeXiZz9ZY42vPx/fhqvqL5C/YoJ5ZOEsPOpw+d9SFwEoLZl
jcdQoP9WmgjOi3SvhDNhI0do4LVdrJzzb/DNhA+JdeQbugz/o9jO50cFdoXr
h+6QGnVqBotGcqSCitd59ZWPhcqjMoQ7zsd8+F1A4InoWDzbH90NUDTerPmO
dhPgf4Dt/T7HvF0qlR3TEKqjfgZX/81MmNXscjwYeKZWIGtPCBCPDDbAAQ8P
UZ6Vde0HurJ592fNUTE4WlIQx7f54SCq5uG0K2sRjtAFJQB+0xKXpIUOzkii
xF+H9oUrtwkONM/kbeXPyaxYRb12vxZvPB+gTV/fi8qT4x/y5k/JJupeeuv0
inyG6DmP53qIo22BD//0ahQLlhToRIHI3ujaekTNlpV6gmQZcRr7a61ZL814
INS8T4CactWvTw6odPqqLIeN+ObnIyWZCDjHHAt7NuGTF80CKGFPMYttN3IQ
pROCC1dIDjgR+9/a0Z6GKSUvMILvCQO4cPPO6rBkWKmkWXY+kVA5thm+UxJE
5Vsjv3/1LUvv8N6+pypC0j5gIgHM42WO0nTfjAgtIgUYXKqWmbNVYtY+BTCD
B8ENIH/SfAjG9Ri0q3hAu+OsDPK3YlaOcT9Q1BrsN+2u/Mqe5iuZ5/5NJX2t
7M8l/Nhe7+hggZeUyYDv57ty11sPTC2/GArKQe13zSDSH2j9sLyRAPWlzsz3
OXNezuHRrD+mh0bgsLa1xAA7SYs31L7nH4v5LuzgK1s8H9CcDA9cpNWji8qX
Gw3LgpZm4s+RPVTVFxhGaQxQmKjujbteKQTpTDdSA5/RoSMbQAx1m2u0roDc
Z4hylNTh4/m3y9N8sb+mpIQPlGMD+NSeNkNdk6jCvgUUnXetbbBLpjPPgV5d
mHNbWmuZEBFI6Wg/SQUyJNTfT66I77z+Ekc8SmCJm6EUOoQMZR0o/p/swiNF
RI0+1WAvkhqp/eoXU1+PMocTRHOt0kpkUkLibeGnNWB6kB8Nb8N70Saz+k3A
0pwHzcykf+W11uPP7hnDB0gu9Z4k9U+2k10+cKqZ9VwmBSZhbO4Em9N+m5Bu
iTXj/aZaORyas6iwky/wIsctyF51A6/JNevtKNURG9aJvbY2N0TyYaVCpHLL
HW4jE1W5ociqD8rRDFVVYB2CT4tqqMAdzmiYgrNyPOcQOnUGs0Fe7BIffKUf
WzGBihSFA1P2hVl3XCzFd7mfI9KfWuUsof28qXspEJXVzpoZizVWlqjYDhRW
iuZhUVuNSDVItti2cLUHUNmSpg2K+ZSCc3ajn/mm99AMLFXVyb1DNCFWJCQs
bEZgnL1+my0SfqqrhpTp/0KXLjjKS4nqzy68PzmD1PT/hawK+3ElhzlA6s/X
gY/WrJymsjyVZ+rKu+YGlX5zbuXyQRVvAym6vYGQ33sMvxD12NL1lfSBwSra
3sY3CUcmJbPSHyBtpvwJMYgD51gWrfgEIH6E/cxqWezxiqffoDa/pqINWZ8l
dT7putCkKSp+lwNiyOHt92LgrL+3Vg2moh7ycf5SIZSgyML66XH076Z6S0fQ
/jj/Nv4oXDGogmZ0IbO53wzCT+so8vVGeQ5Z4Q53uUAKxN1DRVmlgqc1brxQ
qFGjzb8JeyK+k8Ld5fkoy8Ga5H8yAPooKeYRArXP3r3Pt9iSJw7JU9FhG8LE
WEpiG0ieftHRsGVgx3W3fMI3AgOEdUDqJeRPk2foRK4m4Ngg0MpLybE+2xBv
+H8q1vVbYHN98nq7BrzHW9NnQCpORQdPT9EOrdqc/VQF+r2FKiL9I55QfSpH
EYjhALvTBcr6aXT0tkkHYVYxCmFpJRqUbv72mCgl27xudx/gZl14mbSYYmkq
W5P8wSHvZo0mcGvdBGVc89zIsjCd323m/jLKshlDUKnV32GdMI362K156QHD
+6iDsUAgGxK/PJl7++90483gEUhFcOStX+G9N1uiCqVzDW1iBTK+NK4kWYRc
Ub1aBaRM4p6JZoIekK8LIG08jOIzZZblSXSlJmuqJ0bObCm90Lom4PBcF7uz
5QQKcyRaOhfJGPvyIK5ppemNgOOBi/py7QSWW+7IxFGDVMsZK/dVmC1yNjsu
rVny9WHb3YIGsJkj8XRxkZh2FoL+EpKMrWWWZ/S0xj1h8s0fJlbc4aN2jZDh
iU8SN++xIsA56lcAOZNxO/qPd1GCno4/iZBJcATBju/nblAqyKgbUFxXqwZn
cVFAj3Us+XqEkpS5BIkUW0OI8y+q3cLfUhB0HLdcDjeFXIm4m9OiG7vj7paL
dGUvuJ0xsSQsOAt73/A0upobypWnRm2Xjt9Jt9wWcKByYgJXO6YUJemRqfuw
ABvPqHXDw0eL/SaYrZCNTCLU8oDqbiOhDsDg3MW5kArVpm/9NIXdelU7lY68
weVnuDLOuXkSWsgan+0xH9oAt8pfaJZnI+GHk7Xqyow4bM5cUDUmNbclbFOc
Y1sbLjYctcZxbsCXMDExCgIFUfHurb9ftFpwah3lGIA7wZvSx1JPIRmnsCq2
+LCyM+gsNt7+2ZIHPeb8MjokINREjLVxBUrHiCdbGC8Oz4nYruhtrqTHtEfy
PjCJpZwDCW4I7mBP7w+q7Y/YDE5rtKmkZFKy/IoMGK1ljXsJS0WWqAbcuvqg
e8ZABGt8gbB1jRGKZFMRRJHfFgq9otE2BICwaGj16NNleJHcVBBnkQNtY/qJ
qw5sFXexe2kabV4Ep1YxdYauySE8PnhQDKyrbu6q6BcsqJwOkwJ6x5u8auSn
1s2qZxmAYYnMlKBHKVM6ZTDHSv+M3jBfQBuUpVd0oFdwF7ENuafdfxAxtail
yTYDhxolBrSwTrjhDineno1WihFElJMyvA6lkLna3zO7ds9XCbmlWhIp9kL0
LlXbpAlLLWsvOnWWGx3p4I+JvWwH6xcoBQboHEUXgis4ue/UPvnnMsH6/Zt+
BoHQT4zR8Cqv3g5VpXPTh2CDiHlrPjuT0K+YgWYdsYBJwZVE0G7sLzzyiDmD
+7tHF1jxVn+B5ZbEMoH3AThNrgPeFSwtkTVBJu22CKP3F5v594IG+j46n0mF
c6sUwQ4l6cWuWItRIiFaAlxcixSUNmHx9ROnvcc+rmDa+umyZdmMLW6G6F9T
kA5oxVfL26amINzCoRAN0lV4QiQF/NyZcz9yR1h5qL3YRq2z7ew/vKldf8hG
I5xqR8w9mZn6uJjEbPSVcofDtsNNZvxcDdEMaweV7tiKBWAF5jZF9tCL4uF4
SvLbXYIMn6B+6F9J6vtGuWVIV0A2bKaf0pTE+Gy6/f4feet7Ma+sjFBKOMI5
BeO5hNJ5Sj7oJU9jZA7mC3ir2C+hJRjgGUgDUjqGhKwqOTmrASq7toGleDHz
p8Lu2Tzy9T3G4BZlquilooOjo+Ch4JKS6AnpyT/9UJT8E7bzPZGCT+etWFhS
fQ1xxbDv8S46t7GjIQrAfwlNtrG2hXaBLKneFuuruF6HDqhVHMqPiJsHBp2q
lQugsu/DU+QPIIWOs4K1buxdkx0B58Pp9+6xRtiYJeW+wqTvxSyr7anOLxfG
d736AXeTpLuwwd/dcF4V2TCXoqDAYf5DcbCgboMtzuOE/8Xf47EqXo2fomYN
qY8Y3kRigCxCXTTT09wUQyHQHd1Qv5eeUGMFXuFmmcgg4m9HlJIulEINciL5
KswYj9KAAfPNwH2//y8+ribLOIwE2NzONtdqxcvZkAB69mJIiIwhZFh8r2zD
KkRR8jUn0cw9CsV49Ebycz8M3BqxHnh3fxkBRbM61/yX5mxYV0lUm2ZMPF6t
Ng+H2vIzy73dC2klS35Lj7VLwBUZmPLJS1DriQhVqpfDXlh8qIjCD7XFJfes
T/Qd7m8r80geyWWlc1b754fd6AbZ+IM+pyuvPj0yE/Cv6vDCjof1DiSP8mpW
oTpCWY+v0eBE5G1aHc8KEP8B3MXdWflcmRbPFdEBJIRIQTz6hPME5dw5hf/7
Gehp/VJHYsQvdjIXL5EzUeNH+t8LHFhNZz16BrVVSJEtxw6cMBGqbjzVY4B4
Qfl/13JAfDZbBSZy4OgZ7P7ahrvFISDjDgzNImpd0zXEATzfjEoqCNqfZgxZ
wpnc44wRVX1yWUHgpu0d0Fj6rEk4mi+X0mE5S3yr/2nRtzqTb1xX0rKd6nbZ
CoOFZLzNS/QZRKw36wBoaas6rjQqixxUz6/sl3jbzm8M5RnCviC3rJxFhD0Y
LrhVjvUs2QlaIAmVICAfJJila6qW/JcGfb/I9/aLy3WiCGUeuIqqmvZkKJQe
U/jA7asEDdmTY2TSBx+FW87/ATdmGZNOk/LGOIl7tOzTbo6lRv6dBVOHtqkh
D12qG+rzGRLVVjRSY9/KnVk11zm/YzS/EhDVjkEPo88modNavAVWMq4VvtwT
G4E9lseIvSs3oafpcf9Coki57VktEe/HacSzxV/rDj4maJ47OTNLP8FQlEyn
Qv9A1spH+CI1z/QF9+OcKuf3bO1Smekvkh9r0Q15JdsXox/h46wqYVD0FiU9
Kww9BG0mKkSRziDnyXUOUu0GozEG0UogyCqR62HhCzwvCJAPLvqB+Tc9mwLO
GXB7wbN4L+Yu/rh+uFq5kmu0rFbCJi7oUhub3rVh7Wlc1dOB7jEbrEU81U3h
GwjqkaaBLtgtxrw8tJSpBVsY4dvN46xa0Nerg2gdbl376VIRK1CvRNj8bY1d
RGi6XJkIaxAzze8SK9Jtchi9sbZdjgpDdrBponf1BmGBQ4+LPdSa80n055X3
1HJ73/Ta8OUZRLD5LgMCvsi1L3q2ipAwjflIKcQY7ZgiHklY8tBSeblJqcTE
/v4yxRdQdgd+KWFvA6FEENvSBfaHQjYmaDRDPqPA8I+QunQnXFFQHmuXgj/Q
iEiso9rpx6hnwPX6ZjQmRZfPhQcjD3k/8b+ydUZq20m0VUHKqKlhwODrEeZ4
B/N3meflnDR4ymQlP24NHyNACjTO15qfOtlrYQ5QVIi8XqYRmd0HJV/toxFe
nD2bGkA6cwZCp2r+/R53Yv5VMwSXexY+HCH/wc9rmj2kH7P/ZdElwzkzp8oI
wqCDde1YdH7HhBmiq7f0ela3YXhWU3XMr7LO2rJbcbjmQKBSilRVD9Vh56YU
dnCRM1af01r83usDdLudLCxsi/VJp2IJ+kwwusgdeQzahyQukonLiF/ZGvhp
OtJmsAxGyz694rUg79NZe7imZpresnF6YC+EC9L2IN+NOFnon/FJxwCZv67x
pR8+y+JStPlNhggT3NL7DoTSAGIqD6V7BOcE2S3+qespYq8dKL1x5ddsKvJ2
s35AaZQPOstYVYLYf5vk33704mpiuECaywBJ97Oxk+uC+QkVrBKl3yD6QQzM
K596QaK6pMs5cIPuUKGJoOsOLB43pamE4D9v1z4czcewXITJ0XrhKTCqJQU8
MSE2O/gOKqZMaj4+k181KEwPDdOqY0bIvR127FmAwM2oxRz9nYHhIg/zFoGz
V0tMe0MacFPy/CZXgJPODp/NqtDr2mi2aQbOOUWOt/ffpJ7Y4QN0UJ2f+2Yo
xN6SAr3j1i9l+AqqrYk2rFFUIDL3kEjnlHaIrAMOBJ3Ww4EOaNIZcvMDZBNc
BRFyqGiR5eW87pgT6792E2+ZQkleEaC14hWVOWtpvYPbJ1E0Y0l8PhbKoFsM
UCXnwtZsFoGNGlDaPClX24a+69cNjhAjw8PU8cW9s8filG9xqTiWRxmbUp2k
frXn2leIB1kGS+q3rsFV26bLWHU7uc6df0d8o7DhKUTaWnb36X1kxBuMf1iE
megyQ1qGfOhAwI+b33aYlR31lLWG8wbFqWSwNHJhPOYDg+ypoHuyXKUrzO7Y
KibtDWwFPRHkEr3SPL7XRRyl0ebvfnbHAiw1eNkw6tt5GMEzGYpllANhtQj5
WFZ/KY+fbPRm+hfAFdRTjpYAn20VHH6d8J5hDFnItZpQOsG2dD93LDanE8h1
O3K0VG7Wg3/GaX+qGCaR5FrhZBkHoPdQ2TRkKV9FGWiPDmfThqX/pOD5AYCN
qZ+YdKzlKG+4NWFXrNts0xWnCnyF21gjgG/2CeCgwe+HAdidprpZB7YI+YKZ
qN0+XvVXi+9HomQ+OibOyxaki2wX9JXLsWsGHg+sgFeeJciJ8JI2WCEsGFTd
bfy0ZwmK9Kv6H0rOAfu2xgeOx+0E16F8VvAFV+V9pS6O1fw4+pDwntyAtJ3z
90yUP9qF5/tUCRn3pFNqszGuQt/E1zaUDyGJdGn0oxVmQJXmn2bAX8NqB2ll
ZI/N14078wNg2caV1MXx3esHivHu5Q0y4mIOhWc/zDSejkIbENcYGCWE9doN
A9ca4l1lZGhQXHJCVSMiwzPoq/qBgbS1olZKfoOkZN0YT1BoS8//O4PX0vYb
ZyVhIg0hDD9yjrXZYPZr955+AFTZ25uO8zADNplLJGmz/kQr6Pec1+vzzvaE
cg8QQyisIq/MRaxOJRO/0l71RomnIFbURrkdcQ+w1o6sWfTKXD2la8I0w2B6
FwuOAm/RhduaBcW7yXxNuMUj9epsiKtW0dfwdetTNlqpUoBd+vjfUjfZLqvx
4PkstxKyfDFC8uKO/2hB7nCndrBZfaS5ZzUjQXks5qjW5EoC3n4hOy9Pne+Q
eT6AwNNTHaVY+Px+ikPCsZgmsjwU+CI1IO9RWbGUwVPQcIQmSay9joSWBnEk
uk0xloj07w4aYs7/cChZaAFMnA/aI/jBdkZ3nVZt9aCZpbfti3JTp61o26G5
NhpKJ88H4XnEkGXWiPYY5+hUchJV4hduiMEXV3N15/L5PdGclE3jBXlHk7NM
RIPlMAB49f2QoIuFGJLkmkUFXEnkHkAHO5aQOg2sDi+QC93FeOfZMrMbFfDy
IRua7xrLFxo+NnLaVqNeRROp1Q3MvjeLelN7MI7SEHhzZyM22bpTI+x0cRY9
bNZ3RGsTxrhsGM+GmhOJjidth6suGGNVVDZHpJ/vApA9vhct+4p1aN41MiRu
0CJC0Qpp8dpc2Rz70UKmzU4AUXyJdCFrsHJ6yJyKwdYAbsXoNyl1G+AjOUD2
6dNKCR23rZXzvGpdB5lpe+XCTGSg1jwMjjmweeMk2VTMm3usmv4teQ9T1cf8
HCqQ5vmcs0/6t+3nllpotQC8X7Q3UtSYK6m2AUdEldgxZ22lfz2bOJhfcu7r
nqlBiDfw9TxS76XmybTPwu5DjK2wcyqa6EpxCUa4/EBwh6pLuo9PJ+KBTfOV
aMwPmekZhoOXUXABz7mPvb2WZGpUUWR775DSpUpRJXddquJIfw+WraQFJExu
GKL+DkX4FYYLNadWfdPUwGKUZrot5ptwJUamNc44ODgG4onMIcecWGbgF7Mf
c4mhU5+d0l9XcxUZRIaffUr+2oK3SpWnGn7dVtsArEtASoiRcBe0mssk9Xue
NKj9qJH5G4SoPM69Gb+FTE+/WQCrUWZa1d3vW9RdqYoDGGF6lV4CJPk/z0Hz
jHABA2wf95gbxLgXYAPsnXdN6nXiPyxMtigY1ScWEIK+3/aCinP2uu2YewVS
3WOehLkSvH3kPBrBW8BQkQX2rpT7VPKjRdKJMa4u04QFFuwwo8pfiix5aGgF
X/qQjPYOJPqokdFBqH9TUTmR9smWUHD7GtINEuYYvaRaNQduZxmrK2X1hMcU
H696sthJ/jvwzosd/9kwGb/u5WwEL6KbrD3zPDo6d66CbjC6Sk5IABx21U1o
++5MlPXKZQcE+offUPQfoQy1CtaLH42L8/mgyBcHgeFjML2J84WYkVuuHFO0
kRwXVne4Y8OprpKLeYG+rlK77Fcnzdmp5UHDSvck8S35Owux+0ijzI45m7hp
I34hBrXGVeaQUk0FyLKvv4ZZdTAO/b2XU8fzloVdqiY0KXOs+QWSrjECRcNH
72VIlXd/cjZ7+lguPxlPqZGhvDUWcAmy67OZ6Qqo+o/nDaXWXHdhyL3Z8dSe
h6ePFmUtT3xVrCOqC5DT0Yijt8m5r358eUb2SQRkJ0gi+RxllvIdbH3vaugA
ODlQ8yT5GWdGo1bWpUmxC+WlmC5nZIcoPVuBOfv2RdLVWkSZmhM6DvH9vcrq
HAle8hyOJ2UBBGFwOvRZ6X148NvrYtpWTn608cfLq/31b3MqZHmCW86GXpmA
dSXzLDCwJLmqfj8Dp1GiOCDS6ndkpdm0FwgleJmnshy9JtkUC5Y45nlJlomK
LI0P09nyklpf+tku4MPFbhW63BDDt5r5Y/hYUiXf8YqzZixL42pYEIqKgwtq
pG7N0+/IkUTACbOCOHLD8Bwl2/DRkJ1F6XwTCDF5xDPzifIpSg/QU9P3IhOs
Yu75Ya0vq4jVqc9zrKGiTVD3eyNqaU3jfcIZ3r5SEj5J/IZtXdFrVw3zZp3t
MSOdVRRFy484/TuQxDnMNk4dB5OO6lU0DSQVlcqUmvsytciZrm0vVmO7P5Rx
KlU7dlk20oEfYMtKWjAcNPkBVR1SBRrBvcXUnW2s4HUAP98MoZLp3Xa0iSkQ
RTC4u7ra/ehee/pU0RUUQ9gFKYi+rNXecL+1cpvXZVKER0+HeBIvL+YMADJq
JOyh2EeYRPOsQmY4bUE6STL3jfwIPMkOnVbDOtsIGiUTNuiT/XCOfoFiFwN7
P340fBYbjSDgrFdtOLX+lGd+o5dgMeKeQOaz9TsVZvClC0dwk7GXwQgF2sWA
sIQMrEmcVwvmtHAW7AQceO2bN91qSSW085pwqC6X2JwS0WFz1LjfRUcsDJyI
rwZfDdvPvueOXq94ai4J7tqOECFedclY/RxLk1wUTxmnP1bA7kDa1ZbHXs2C
0pCOz7JfeYPVxWG/WRYKjf1OLQB5+VNqlcMoQVsCWu82MjQ19EKsnSYB2RDe
deE7RNiz5UhccMq10CPwVOF0XRlvP4t/FFHlDP0kwgbN8yC4GqzOu3gtodDX
nq/odQwX8RvblgQGg6wqWP8mLw87uKzwkSEg2xdiucg8RQ7409qsHqEC6fEx
Zv2W6IE4d2FK6/fysyRoZazTGuNDwCrthRg0jp2H+nm8RV4QiwijZ1R9NeyG
wubIXmSOlrWIkS/HLhxSKm8givm1o+VWrmv0FSx1VlETvlBBgMkZHJcBotME
+vBWLfwnoiKHgLz5H9s9vxH382ZHea1Pc+YXtfmJw4jnpgRdjRa4Crl5fBVC
r0hO07md+IiffuE1gZ7ygD63UIZKooDMDwymBzpbd5vJCM8DdpMLnG2MlhsH
3PpysfUY+YKOOB3cpotubP3u+rm80j19laxfkgFEXV7/oPANcOgABSiWFwsM
2LQA3JPaYL1QN79bNghW/IOr9dYltO4RqH6BvRgYPqFKQspv2JCjP2t6Sd1x
ccHgTfAu2uaHDMfQMD8ZhGmtspFD1ntRh6YbYrR8pdOWSTh+oAU8LDH1FQ6T
4JcOgMdgALJLOfCNscy3c8u1ihefmL6cj12CDF7qIYEUpPXrFYi+sf4xrphs
Pk+1GI4SdRiYjsosHmWK6HJySwC9UhKKc+uNTk2PQI/nZz6RjsaDZvZFA9Y+
qDvlt8EUETZQ5bAJeXR5KhLNFDyQPHCKPG7t0m7K52xJTqZS7QkEhWXHxuqR
+equbIMISQnxcj/OgoSvD+uqBbanarcJEE/wHds91GoXdpbE+JWYRiCq0grs
0RCWI8lVBhUBV82X9TBmlzxTkybw47XZGeybFeGL9e70jwqm/vgOmZD9zgK8
U1FWYdBhf7IKnlEKGLswgQYhqcvvMssOFfcK96Osy+rd7vhwPwLQfIbPaOcw
nPtyJG81t2JPyBIh3qN1Ox/Mp57xw7p/RBT3x3x1aaR9RVuzzVrFO7ETdLmh
kCZIrEM722i6z+GNXsYVCPVlQ9oZzu3XfsQPqhCEi8Wbr25paP5bNHBaQCHB
+3StzUpSkpbb3eg10jac1sTMH2T3jau4+SW06XGxTbtXLhOP0cJjXVjbZ06B
IlLBQYm82nKP1svbs/cqPojZ0xE00eEwM8HG/HrR/ckIj1JtaGFNnVQ2BW5j
PouSGY00TJ1waLpkFInSnT3exRlRPa1qJSoDXmDE8Oib9qzIpeEHcMYGHOQV
R+Cet9XtbTqHg6hQwpnOFHWp0NnoucYeI1YBTFniS3hQTnx0Uv34VJWLU5pZ
j4WY7zb5TrRsWbT/Jc61kCsa1Lx4D/MRpoS5O6lexVI4Sdkn7Y8Y2TFG+nun
BIZ9xrn/Ii1Zc3WOBXlgJi/jug2ZCFnhAzIDg941uEiyqD24JKAs181m1EjD
QCeFJxTlyDI3cP6G9EpgoqUb0JZZVQx6/dP0rT7TTFr8r8k4Iu7WzAHMbCzJ
HS+Zi//45CjU7uWck+/l83MvSm6h12FyUd1F9+4YEF4tN1DxznZUYHlB7K4o
mPEdu6tgn2NdlwmYm84IB2AfQc4Wv1y45mB2daXA6roZDJNRrCHNiwJD0bdZ
G7V3UYLLkF//0BJT4/0gbYQm3/jSlAVP04ZY7MO+lmzW5/4T1ljX5jnaVeok
sCuz+KLe53c7sjOXP8IUJbKTdnMxV/czody573lvVuoGyuRrfY6jDCCHw9ZZ
TblDzpjFDhaeEaxl2j7V2TvGe3x6jakHBGmh4eZ/4m/lUDx95H9QOSlrBp+C
muwC4dnFMPbLGMGa4HFUN6vP++23TTA2TpMwoVF1vkmEugj31bAnZIOL21hK
nOYrgrvs63VMLviNDJEIgPONF7eZgS6Aq1UIEM1x7YROIbgJMK5nRyY0/451
jRygeJxnr0oSoeIwmre2WWHWQtpPNR24VDbPLapJ4xNLte6fBAPNzmaqbL3Z
t5i45d7gKjdoClhx/TFtD23gmbk8Ldah7Rk4mdcV+aiAU6zzP1+jrUlxbQZv
KlooEfEotY+a+ZWceM0WcFQNrkGofhf0BGd8rlZdezCnzRwbsLsMjWAhJUXE
o5y75QeKkjKpYUGAs0SFF3ef8j6We9JvMz6ddrzV3mQzQat9qI1im28IOCI1
vQcBOUcTa6hdh3Psxb03gTRkSNSFuL3l6oAVZsr4QWfAVsIPRUHATv/MrT2T
QCnyLa2r0z6XkVRUnf2Qh7mq00qOAa7WXZMf26JrTlH4thkdzDu2h+FL1RBl
a5Bzv4TEIOab02dCQtmy9gYoqxX7ltG1xnXcH/sdPurnpS3NFlEiYab/iNqb
uyyEkF+/GQHIgDiWI50hCMkosfl2AjEy8UVYyDMMbwarIDMNT5qqbjv3Y9sL
J6rIBpKomer71w6A9VlaR/nJOf5lelOVFGXkwmpE/gRxZ8QScMc7AlOjncA8
AX/IHmpE2R+gl6YLeQL4Iv1ieZmi4xdNdwEcEz5Q0NCqSnXOJNO/WRb2vL43
TV28BD5jr7sW8s0bhZuGDd8VbYkUFdjCm8uh6aSG0g+kzKDSTrLTLJRVAGyW
Ji47nsNQYGJP8kZqsPkfzajTHaQyZV5LYTIsvJ79diegnGzy+k3k92ItMKag
I9brG4V6FIxTPNjCh0ZPl3xehbeRf0Z8ueKcXP96LFEXm0URxvTlTNZu/RsP
5or+O6dOMbt0otD5FtN6Vl7OX/xEJ8o2CuSVL3afzHyCBlfWlKVxMtvzOPMh
+y7+jhkoP0k8vh3sPOlQQWqGtRCJFm1JK3QvqmGNMigtOB12yJ8cEMDn65zm
IuhK6dR1u6aY8SOBrOHY9IPqevLxRtv+AwXahjXMSttqhKSfSf4qaG2vBeqc
T20tbwgcqYg70Ssp8agb8VuHa1X+0+MP3R1jT2kPS/21ceJpKDyRyeSYzwE0
0xuZ5ziHsXfUXztHt3qGNVNZWHm0Hqpkm5mTKpx7zdpC7+JdkpFGBDo1UtSn
oubSlZ6hmRUNmkTjAUzGnldjqsTPJAnvc8vnUWQ8yJ5AWZ7/gBnoU9X/Z+bE
1x1jN/fJn55SDl9sobb19y99N4jvk/iKe0YjGbCXqzadLzL7gsWv+HpDn9Au
JtCMZH60I3t9aweMF1ErdJL5I1uk0J/oljxTa3EnIX7j7ksDYOHNoXCDQICE
eVK27PpIxH50MXo7mVdFaX2EK6W3+SDDl7UlxWiI3P93EeSeA9Z0Gbdeabvq
X5Ts4Fw7FDPx4PsvbHOAJitTH2Qf/lNjTnmwLXJN6Mxe6ZKdknybPWEFrYvy
L0ok04u3QHIRkvwMa5ymUtqtXweve/Uxxvsz5d+hp5kljWW/mpLnpStl7bly
932/rZmWJQ27FRpKATPtbpmi0qtpEkhMB+cMcfcBJlmqR3w6UEIEP5fsRk87
5Yb0GDgx6zaKCKVk1pn48yNlqAvUBrEB3pU2bjymQneIQ+c7DLZZu3lHhSXz
BGhxt1TvEEz9ldrdLJBpjXax62XcSiYzsGHcTFeykLDNKD/iu86sLM2Ggt/s
nv2AOERA7ECB6i92qhrS/7ArlXiRO3UUj9AmqcL6QyrxoJ5KV/Yb9eXMqj1b
XQQ2k0v6ymooTZT1t4Ruby8tT6F/4MpjcYz9yy6Pf9RBsG25nU4//fK7GGEs
/twNplbP8Ojtdd5kQcDx7ww8+mrh6ZS1JV74Y9goWuST5w23kRXOBfcL6UKG
AGJ4eCl3rVYQuG0l6+g+wrxNAANEtwcPnacmfYC5G+AxiTGAhw0z8f+4bHiT
RvxBJOFXQp762X27+SnZ93OJpBCnE0MOhwe9izdRlmYOgshMSRalKGOSeYvu
lsPIyGO9+SP3XmrCn5iIOZU8X5Sj0FxafhQhbjAE3h9676mCQr10NYdDzLkt
eKHfqXlrfbjapPClw7jcCoOEGDDfFSE3fwPfl2zyq9DnJP0eAyaWIdfKdIdQ
QPL6XNP1OcYEMzL5RQSxr4bnjeappP9td5BzJziFmNSUgigFJTAJ4G92MXdJ
P55TZb6kS/u3KLiUf4i2uxzzOxS46EO8T36o9luc/JD2ct/TRvuJdOkWwDnQ
hVND3wcHU/SG7ywz2evNvWqYfbbMFKG9Kru1dJ5IzDSIP9WRqpF5vpr+RO2h
3x5a/lX14ksvSrMfAtchIHE2FWkL9orqJQ+m9s6dwiC20w8Jngnm8/p/2evT
+mi85SYgNFyuBBbZnNqOb7y/52Vk9S1mlBpFF1QlA6zJ3vzt77dstoqkvhAS
5DhUzpvoInxNLiOpLlF3YDwsaP0BqB4pWGucoNDDDpmCtR3dXSc9TIBgv3Md
n1d8cDp0RdO3ezvkA2kwuYCySxA5ZzQN6SqOUv9TiuNYweCH1zpdRPXCx2Wr
QkbmcnDxo5Zb1TUygWtAA9rO0DvP+ebN0t3+NnwjgAC7apsg785S2H0YYUE6
onqlwD5wXhSrPE8/XDHjkKN1twyvLC6liKNXH6ACQTrUdEmBOyn0K9yoFXKs
PqEGZa48Fknm94D/X9s205nT0Z/iNOOCa3boPYMh0J0GPGLb4Sm0ZXm2w/2f
8a97afOHVbSGIP1GrfP8U4C+fevpQOnytI31SLd/KNm+XrpEmcq3amXbj0lw
2wpMygXuhOvu+l627XGHAFBbyXDfPNxKv8XAGzEOwBP/sEtzYLfQXQzVYwU3
l25wBuYg6BExlqP5YP4tES+A8WrA0pjQYU5qvsiYLasn4BNu29acc+R+D13E
tFB0hSoq77EioZpqjm5xP6hqrLhY25bLkdu/FHSVm+AwvS83PPPCVS4z9D8u
XECPMiwJ4BuVuVPNngHpnfx7U6RDD0OQRaXcFzYBlbY4cefzGxuVKPJiJwc7
XaCy7aYcdBNvoctG88rVegZMK4pbNJjpq+VO+M//R90wm/Gn7mm4SnZOJGvA
Pm/EvGXEIOLZW78siZ6t690SXOu/kFmwuKs5t2y+gYn0YvDFmPu8wtNxgGdK
1tuuyFyYaqkJafaXRYSRK51ofbGXKMiDIg8W6/ujDOWAr4gZ3QDHcyoWGHWx
8K8WGt9vAuISf8SLnzNLOxWcqXWf6/ljuUsJLB9jqmGBPGIunk9GZWPqk1FW
6BM16VIg6BQe7nsdfmeEPrP+r4qYSVRnUyvXcaIaeX5yJaFKZCDKJiHwMq50
Qc4Xm7HllLzXUf3MbKCk7TxVn1GbgLg5Vs2w+CRAcwjt4vYlYwXcKwQrlB+f
5VmyUPOWCCMBumHMkdr9pp8AR3y89fcfy0uQGoLmEitb9k/2tGEkAHkv/Iqt
/UAIa/5AMsye63GOZOBZWi1flpQWovw5ryo7pMHDwlhQb4wRMXs8U/rYvRi6
tUMqpCc+r+fGNDypbcGSz7zAt8nG7jP+odfoMVMmyimwipVAtGDRyc+Cm+re
+3/7Ny5TZww0twjrgVkgxJvhqOTefKdv4msC7HzJbxaiMTjmV8dXR6eX6jJM
XzV4gNTp5EdnC63QdAfLvA5YFiQ1pNPmPM1pPWQsz4cst6vnvWh6yuXQH9U7
y7PJRKoyAhwzRieEofdn2LT1PIGdx/OjbmKcLmhq0EHDOd8s8J8mcOvGHXBG
jfvSpCzMVxJbUsq9rD9TMVr/piAVnw2bUEMKgjjasUViu8U6vFhgNxRlnRw4
Pwt4D/g20b0fGXmwFtj9RPLA0IQYjwLDTzLLQ+uCtgfs29NlxnvxPQ1boYgP
wkCAIDUszdBILIV9xOKBjvu7hcT+0OBKSvoA2TYo4ECb3yHVYfGSqNwul9b5
55Z0eAoZwcram/rdixA5pC3khUiwMYuIKMxWNarcNqE0mgnHdy668KbwPtYN
S4KRlOkDWqpK74mdXTFWTfV0YS5YQRZXJqkceFZrSDzsoy59/3TzUex3O0fd
lbpW497s7GkDGnbqyi8gmAB7baaLmWrbc0PkLrLEO9pgvarhKDtW1K5XLCPv
cXpF1Li6j53UEZdsF254cTJ58rJltlb7qozk4DGg3G6vH2SnjfX+sfJMBJjn
7kZBSkqiny+ZnxlYXwibyTC1d1karwccUDdZG5PiuvUg/RxlS0919xnSn311
ho2GgBJFn7az++efvH0WJ/RPhBG8WiuMVqTawGfqhf5iCiVJoNX6cPFuNfkV
Glm7cdD6O0jpvBoDkIIG+igHw2Gh+pJOrmDYuWQA8upk5Ta/lNh6ZvTvZN4o
IX1zh85uDNv+O0GF2L61cYV0Gbu81Bn8WMuxaOKpf8/uWC+vEj4F+grEyliu
Hfvc35cISvqRHCyZx9ma0a2x9jk9L03DwQK8BKT1WraX4GAnHPStwmjp8aE/
lQq+jZvKPlxTLT/gildnDpdj/10RbxXUFazSjwktpVXKPOI7RonN+kaZZyqz
OJs+STXB7MjVBMpT6etDi+XR2vvIAEzkx8n0O9biFBLMjMs8i9kMpB/UIray
jOS7uk6dRmHojMjtyKjEf08YmtwvR2qp+ZnvHUr7LO776wxAp4jnfYjJnjaK
qS5NwvWePia2RDVxrvxwFO7qsPAMzVmA6nhxfMfiY1AHhdIaHrzKEOEgiwYx
Ow61O5bfgpUyEr0BpnbOU0zljv3uTwmIQRGOJIdKnQdNvjEFQ4+6gdVt+Aeb
YA3AhoUZWKUSDZY5LjavncCrhKNmarn1JXymOmIyz3EIbzOSPGkNwo8OMtb3
nq9VAD4/CbJgcdjUgYuVibgY2ebmFULP/18eezpsFZzWhJ/AS3oMNXpgh7oK
EQB87GlWpomiUSipt8SN8LMqMf3iECMAONpuHhuhbvGCTV7VOfnPFWf5ByV4
xbjJHbNYp5I4gkz/Tg1KtQ+YlU5mXjKwF8d1dRPJ4MRtm216L9+y+hnxAFlG
XeThJYsCkXRQ/DYgUnmCgUj485vBRxIfMro27eXL6e3xZJ1n0CNyBr6Ie5Sx
aF6ZSw3+0CRdlFCJFhYHcDmjplfvq0GbsLy8QAhOy/FRNCO73rS6RybaIQlF
bIhuNiUOBKvsEU1isqmGEMyndF5oHzxFUul3wjq2pnDCHqz36VqwRsEAQ4Fm
DDAVx3h18bECbKIDjp3mR8rBXzJxu915tTF7DgzzNy9/aqju1d4xiBACgVVK
WxrO0vYEAo4mKVc6SP7SFl8zYO/k9N4wn7UkAvQ+8TGdfluTobs97flbM5kr
59SrvcL3YmnvKixzmBIkVQq9Jz8cf4NTkgVOZ6gL8lBU7yeudZRe1qrrD8Ls
K91fao6MsEgr/4VJxVTmDjj6B3L2LGsiRlXFJa6WOfR0a0YzXqbkDpfnodqH
gwQzxOohpnRbY3+ZwjHTmiN2CoBDJ4Evqu/yO/6C6AjX3KwY7ya/O5ADEoFK
f+rFUCR73wpG7sbBRAstgxGwowr/hmzaMwAIDCSz3oVKBVH8KD0xznte+TPW
ln1VRVkb1EreuoaOleSK63AsXUuq1Oy13kGHWsjfEHgN2bZYH04jnSK2ZbBI
2DppfBmoajCcZsvX3gd69CQQj3TTbkvklmA/1JJKjKWV89/7iRfWogeB/g8i
iIZAzFxL18WTHWg1s9QyO8mpXUfwctdRAsyET78V6U6RQpeQElOrlh6iCqiD
aAwnIY8XENrmBoWWD9S+w6XKnCvKXb7AcKRf75jHV57wxLzWaLDnGcymrfYi
rswwiaantFoMK8jZMkycA4ofrztQokhsIFsbJujoRQshOkcplXAe0OT3i/29
41o48nvGiN/ACGBA8RodaD3YwWr9l4pvSijNLM4YF2k/w58Z0AL6dTOrRio6
gJJzCrcvtPS0CUZMlmyiBYiO1A+PY4pzM++rpTRUDbMyv2zgcVwsQUNk3Fhp
xzpG3Lqo4ZQJmOBShs04JSIZ/ybyc/BGRkztJ+OOyePPowpctZeD6f4uMbwo
A6IqDBMkRtlrmEtlfN6DdBQFHqo0s3l3Z9o5viZdn87KirQKIzRzUGMmzT5Y
gQX3nz1Ui/aYi3fcXATi2vV7n9qtVk9/WehW3+nFKxzhWZ7v0Ye1m+4OiuUf
y4AKfXzOPiUhqRXIIVu0PCiETivU+4K4bbkA7als6HTCMAWt0torI5AKJO64
ROxCXBDvSeswNBI1SycI8NMy869mn0IrIm5nkjLvJr8suCB840+UYPv9toOT
CKBMR3oEa2FNu6DSG50iaZxupLZEx62KWz0tPdEsAP1RIrQRs6cL7goFpKBS
JX+sr5LnqINXx8sQc/PdbgYBn1xCN0wIJ71z3Fc2wmqjRKt5AOT7jM9yVpUd
taz6YiPQJuqpsP6wyd9+FtKGZvygECI/FbNUohDNevgTqy2unW96AZG6UxA/
Bg6loU66U3JgBzoUGXbkcaq60ZT8yXPOVFAZaIEE97ZdIuxWEb9XlOG5FdHR
lcH4rCcjUjP3xwq/uVugzSHhNsCN6bn700avK2k6RRZsKFxM0ROTFHhNqXCn
JOxL/y0BSbeAuYTe2g9uOvcJzY7oh/KomPYT35F8eaxk+3ZFDW1Il1ghQvo5
Qm1YC4W+E4STLL9soruxYGe5W2Eh6NE0GbT3udnaIQG20fr8ZEmp66wlGr58
t6VRmNui9MM2HKI6hJW6qg4yR7/DayUxdWAIHA0cfSq435iXgwIKd5qyKPka
Zk6qUNOYcXSyyg6yuS/VNAKJRZgzhxT5yrYWlJHB1BWdJvzySyZNuRF7+5hU
rVFLI+iRDqGmmeh4tz2TIj7alD+sc0WWEF9z5kYv+6C86i8JnHgBsWyTuzGr
H/XsMHib01mRmnusZhOB5u34sbaGwhpWOuxb4btbDN7i+xPMTR80YT2O6Ey2
9O2KRzmnGSPQOhcaSgUUMSgeX/C6AaQi9Gz3rEcOk00ad55sGwNe90jnw3sS
BbS+6lRh2PpqllfGDIrUnweHc4wv2Ql0NZA5qIwGi+U1qaZcrSNwfpEzhU+J
jep/4YwnF21giU+RJ5HfxXPzGG+bezcHhoiGn//qytNua3UcGJy/HrCousiF
B6x7ruOmT8S7Cz1t75mACLjV3O4dVUS4zl51bEKynXbe/0stxTty0jwZOaW/
GlmWp2EfChkwXCZevyLnNrf5+lf1Yg+o6ZRDoE4NtIT9u1ab1OxSiof0hmTa
0+pSVlJXc2dLVCFw0Sk8lsLXL7CawiiIX+oOR8S03Z3wbmWdka3GmY8GICAH
oVL069LgKRdS0WJ2Au+LhHNoWvBXQ/jq2NEBB2RTapZsg+KARDE1S14ijm1/
jac8WsGiPWwZU3n08TxqWssAwZ9VBbNwQ9sUlB9HwAWb1C5Ml8y6m01Kn6ok
L5zx501SjziucTFPOh7gG2E4IUOfU2tcxVcoGhj3TeMqxAVD8Rf6YE+OM99L
8HGgUTqWCa+hbiz3qDdvAYe1NnK9cgijx/xGKZpEnfOV4/gkZjsIIRSCznC+
uAYBH0Lq0z7FgI0/yjhY+bCu1eoxojBiHGQB3xznuuuA+ABgleEKyv8rWwFY
IppuMxIblSdTjVQZ1hnDdvlrCxs42GNL/tnw/pxXAvNwakEUap/bpOnIC56o
UrKCYPWccyrhoFS2TqXFaTJFuAY2lTdP+lBQBVVeXxpeRxjgb9NvLCqi8sz9
mwqYWpN1hVf1Eu/WFR4r5lQuINcNyWFvlGN5DtoFJwLDkZwFhWSic++xebM4
Mi1Vb5E9TOqOCa+ZgPPpAF/UeyksGJoTfYISHXTDWihf5LG0UKFSPEL0AedX
pjzqzSs/vp6uklsBK2+IiIWcBeICX5vbfOQNc7dtN6BONcdxr+Zri6w3GI9I
CMlXFX78ZB+o2TSnnXBNzNp3w6SR+w6IYZXdP7TMo+ozt3DV28DJkCwB3r0L
/3BHToafFYaGimPosToVMyq8GARN4ajLDehA0UokbQF9kxHblsMFWAFosT9K
VvNkH3k241jhm/Rep88uRAlJ029Gy1UdU9OQbcgMlSLDNqsWzu8yyLvPRM9N
auM863jTaP/p8OMb4uyNUvSKcDVDTtDKERm2zmXDxkoaXbfIBcAYBDQVDuRF
ycSkFluq9B6Hhy/vk1vOsyiuvVkNL7h/VlBv7P9yYEir0p9VN9Wi2oYyl6MQ
Pw5VhhMfSUf1INVHS8YcHCFjFATwb+hWsbhNU0W9FbEc6bFgWEklvZai/lw8
LUYEv8E15ni89e+EBObvj9rEKNkp5JLnrO0W3sXCY+frGyf31z/c9tAr7e+Q
kS/qmm4225vfCMmKCDWWNhT7pLEPPWV222KFtx/bxO8bZPYjESTCLEgxeDwR
9RDC+O6rRZKV11PRH3e/AMbkyuBmRyvX/Q70EJvA4LbhXfKJxEtMtszRFv2O
DaI3pN/cIUb4xHZG+0RvA9MQ6RsRkiAx6tzQgDxjG0nAFxSX1pRKJc5Gn7vq
N6jaNi9HKLIclnOCzrZP8uWdCGElf4VibeMxdIJ6WiM4DROC9EKRQFAurG0x
3JWY5x3VS+aQfBF0gE6WSK4YYTW3cauFjVDF+1Gywg7jBBy4o2lyVdcxaddg
KSbec2bPMKgQyvv/A3/nEhPWYwhaEt8Pi5Y4CCxNFbeb04JKHvFn3C5hopCU
JWlRGAr243O8GxA41Ff9DdNk7LVg2fZaXRELhJow4ZMAQB9LaiFGnHfyJkBo
apJml5ELNj1oE1QdEkkbav1VT6CZ6wYIwOo4a6RjEwy6b6KMRPeyZ2sy4DCr
V4x04HF8Wv5+ftM6aIoM/jpto77v2OB7ncnugmnPtXZLOWIz0EfSWey7Aaeb
GhS16rKV77XVlBC7/vNZsMH97/p38y7iY7PIJjH+N6EiStYZi7I6MyiWHBSA
UrnpzKFjnvj1/zkIpvc0T9gXE0u1G9lhbDfMI+kTqq/s345klAEPCCUl8XDk
85KFUGvqB/OqF1WSOr0205yOKaLiCIWVtzqbFWCNGKBoBT5aDxYqu19RLdsg
d/ApAJq9tvNv+3UujDyotDpLqjrB5Y4US9KDH4HtIZ96IE1MRKj+fhU+nwGy
gBMGgJIm6t8YGgKYSmnzcwq6E8IQFyBariKjDqjryOM0/7DyofkywzmiNN0V
uCNH5E/PTTMmbna50yBEupoCgaOwalhN5KAkJxqEXmqBOzCNxw7AC0a+u1IR
WxDhdHiGMPC2BWnrOsbCEKXS+BdmAsXyvFK261L1MVskJ7wknwWABMaKpGbL
id7ZMcDtYVI9ov/Kuvxe3kkWA44TBxY2lrYUyYQgp4hyCkgUjoy0lqkVMUf1
yqi2SZMnnDb/CmFG5Iw0DwtrJJICmMUXvV2rkephXCynl8vwiEdmCAOUVOaC
rQX8Jcj1EU0CWJKxBY63Kk61Gr/otWYdtk7gCO41IMcAW1xrahAfLNS1jqr6
q+V7OWoO7PA1GBm7WuZ6TBgEgtl+e7f78oh7F46K9EbE4AWw47BqC4XyoZRc
H/z3+gtqiH/JlME3rZFeqbNo90iE3mhqjZzlKT3vEAuBzepXe5nwls7mcYHZ
ahnwFzleQWmt+Ex1mmfX/EgHm81i6vbioKzj9M9bofB/SaMcIRVd4VgmtDoE
pJb++E3LWpJ8XOxh30DmBZnOuiS1YFn2ll1J7Y9morK2Xx1L+I4Z0c5V9z2m
qyJsi0MDYfmJkzpQ5Ji+TdJJFKW/lnbQ+hNw6Dyc64Df+cOY+0IBU+mSOp0x
BxMAUA+oYGYVap1leoGpQrnuM1KpRvRJcY4DoDJN9vwXkxPO8RzwiXAchcRD
4nXzWYo42NYUiE7be7ylCBuN/J7yY22VVaq1AQ49VzD/5JaYNQdYT9fIjShC
TklMnFINVuCfzBY9DoT0xpibcSHMy37F7HZgP0MZkZKKrXk/XXiEpEe3lF5a
WfkkX8Uuy3hIecQRO2fJ9qSC8N+atJ0MTe7PDSM6Q2IQ+8ANHWfB0AugrMt9
HmPn1qhmyHqaTvPuhHrRD+eS42FHaIu/B+LNUNC3GR0+jUFIse4LV/nPxDvM
YlYkpJV/FhXZy1T39fHTXAkleve+Ka0FQo+4yTyIFJDBS8pBG23nxhU5gXDG
vBBFQuQDxH3SCaIf98Q298FLLdnz2ssoYOWhqmgyzTOIYIw2EmwSCpbAs+Tb
nfvmPSmG+P+2t/lWEnT+SwY3zMQQbHiHI0Gz0n6Jky3o4SjgXK57UXagaCqQ
U1MSwVquDUr1PMdozLtOKWe0bg1mlnBbKrIg9Q7JUS73PyqurG15wRxMrCgs
mjuzBxeEfbK9pe/kLHiWjHyFhHoxELw9APv+UUyTGNhLruOwOW+DKzzgzhix
MWFLebLKf4bKTwK97SCAkSnyAEigOPtjFSSXxjitt+/Nlf3D5/5FfIYc7OQR
WxlehEOyCbvx5/TYiJRZz0yfXRlTDCIt2/M/Y3BI7MiSW3kiPrYFthAGTeDh
vn5/mWSKe5k4FghwSHtUjwUeiNxZ1RBOiFGrRZ57wfDErGaxR2KVceXLqUig
m3eYka/gHgrFxzidbQuMGIIZJZnRxh4NHu5gh6EFaccvt1yt33uW+uTan/iN
bIpsIumZUZf1pB8R1DiQgGsghVPk2jY3UayiwRMLXpN0Md54EI5b02Gkf1NX
C+hI58agFSzUIzUepo/RUuasRZNdOAXhsKWDZNDjzQlOYfr0BIZ+XJxToLWB
E99g0FHmTWXuF63u76b7jb8uBzCjgj0DTD6IFunM2F/bsb8ANgFowxOry2OG
hcLe70RyJHzIHrW701TWxSVha/KgjjEqoRhSfLCq4UPDzoKq4A/nxSXf54fU
IP6kOmZr9trU34q7QWuIS1skYSRyiKrZ6wNYUHhhO8gcklDjjwXkj4G3ecTM
4fYG8pE3yR5yzEv1xFjEmoAf5oLNYEQhOLZVaB+r0KRUcgxrA3/mc3NfButr
HNfaWVtv5+cKFJkQCRXLolJqdZu2dUzIpvc45oHxt4D/qWD1PdY68tIAZAut
13nWraIHtzIuWZk9eqTvIrdJOql9lZ1O4neuCShi4+eBB26nFy7GAmbToZuQ
mIxTAoZd2YyRVBLatwEH/2IP15zEB86IH7Lb/SH4VpWQJjpVkN0bGRRrQbi7
adJ8WcOKJiL8peuS5pz5JDYLGpJUU8KrjThlBCr2SxNXmfDnQ8bgZjueRs/d
+xp2SmTpr3o3ucby1L3ufu92o8EUXU70X9Cr6eKhESpTbDgmSDQyjSCgKxgI
vtB5cxLVjfatRHIQTCNE6cseUix93qjb1JLXNERLPgZ6pyJTDYmRbsRFVDYU
Pcfui2cl5bmT1La13akOazvPwrvOax+fVB9jdSoUpmTTVqqYfPmOf6/sVmUo
V1VnzAzfp27Jv26kKVKlPYriJeeUFY3x5TiLLMKKb9063roo6X1lOJal0vXg
0VEHoz8V7Q00uHlcI+fjyMHKDBvewSuhHkfYoQHS6V6q3zx8UFdtq+0QpyGz
2AsvP4d74kkfKFxbCd8yXDeFdDzTKgkj78MmAUOq5URuGERxduXmktMvzIzj
bZsKtzpZrT3MZiqBaLSMIaeSdN6sLSr+G0vC0xwHNGF+g5XatI2aqr+WjQUU
gP1iDImz9IWJjPEcTMm+ycQw8T9IdResyo9p9xH+Gud1PrXAPthUSsisdsU2
Wjq9gFkOZOd3OKBSKMXH2fdkNwl97Pvxk97Uz+olNUEFb4ZPJVwyQw1E1ASN
rUudLgds/INZp4+N+86Lh42ra/UU/60JD/ZYO0K2c8/oitDX+Z3g/5F+P1Ue
cX4MLNSFoAmZpkHN1BKaeth6L9ndjZDHft3JdOUQqp5w4bdul94R/InEvkSZ
ii717CgKGuhIjRGor9mfDKhWTkv7RI0UW+EkHHDIg+nSj7f8L1kKIKQZHY2J
JHmwLIPLwTMqbLMjjAxi3NcAmkpUmOOLJDAHH0O9xG7vVs8sYnOMrx8rTFp1
usMOTgUOTx/9Wr6sEqlKhugR/aeTdmEBlb1yw1PMadcZty6mZ5t24D05es5H
dEUq96Ttpu5RKy9ejtImhKqQ+HBxpqIEPKuMG3dHj65UYBPJdNP2d21T+aWY
2EHV2ok535UDvN+X8l5iSIy9G2xVHvFjD7uTYwOeoykp3TY7ByDsGkpu3biv
X2c0vXtVJzwB9auWv7ZyNOQM/N2EeMSwqxRTmpiFUxiDrFpjPwlACG+O1B7w
fkn+qE5O/oXLSxWLUJwwV2vuJ/hyYxgMfeHWMsPbB6fyIZyPrASyHkEnWKpt
BuwrGdd/2NsRUDoI5Bmit5w8mW2W1U2ELZf72J9pj/2brK55YLK0U3bB1GBn
sYZqSqOIS/PSdTj6fMtGsm3Hczw70DKnEdU/W2uTI251lbXvW8FjORerxrF7
9d3wnJyh57ZdyusGuHxBimv7NY5T5RS6BpqdiDP/4e/P+MpMTumOH4uECCy9
CHDI11wTHub4fGDSSfy2gFEKakkQnuK/vh85mKGHGcJFRX325Fnk0I5+LduU
CSTrySpZF3ibq/RmJOuglHrkB2WYhcy0Su/qccNp7Ufz5dRVfScUYEX10aOj
AYapcEyN2YnletL2Hl8I9jTwnucW5GIg7g06dr9lOwpfa0KybhgB4ZkpWxOw
1Z5pXMKIZtospGYNd1tUTxn+oUPlStNbKpGOhpILo4J0xGtKtcn23vluTUtA
4pr6k2vgjPd/TOukURRBufShA5AcfqjDdwEnq/gOTVo5ZhsUzNDd3gYPPIcG
BLDfejldM3mygnAd2BmwJc9d+v661ppZ5ZnLO7nvvRkuvOY/5eYnqWO8EKyM
h0/fsdb2OpwoUXQy9Z+yLKOBc9xJ/WD5QsW1bjZHJfwAlXrvR8XzqX9JToR2
1mLisKKqeeT7+/EIJTEi0ELh6PMGqZNz0TWkdU4aoO77a2gFvn8pf+B4KI2d
y5vVSKvfQaRRXjw9LXWw7WUy0ZccMl1iwydQiA72XnogEptrIszkgOBJAJIK
LMDCxzzRskV8NjP2No8AaqKiewtbaVBRlc5/7RpI1mvzsnZOgjvDrBSS2I1D
K4rddkA430oqRKV7NrvibcrVBUq0um1cjvqPrF8Ig9+s385hOGoquiQg+qyo
rkvpnAnyFD5wPfDXvcSNx7sMnJVHPEozCMM5L36ylv+udlc6oriczTROjCyJ
SytSLiDHgU4AO4se/K75Me6grqySoUXm1a+QDTq6z58ukOyK5NlygZThYbKI
gm/KP6BfNfBzkBcSmzClum1J8l8c1KuxLW6Y5joNFvYB5g7K+d+EHgr5ojuc
rydShOY6ucDolk+HkDoXYaXwwePI3lc2iq7Ul2E0hvBYGbk4fzZAtRzrvkaG
HKdDfbRFYOOw1LIeIIPiYjlrx807Y9ke1AtwK6i0xqjU05VIpFh8hNmNqFAk
csvcR9XBtaQ3VjzBdjR7SOJ5njtUs4wUIiEAU1d0WCNvM7rMEeA5Phb4LyrU
9X+meqKS3jl3fC0kiZakbCfxIz1vBSvLUAITqtJa4+e+XQigELdIbaB19jjZ
q0VJwtjpkhY8wtvLDvrVOM11sfQa8OLwhYnCBPHYNfUJsdeMKUtGdPOHuPBP
ef0zlkJuPCcqw2XF4J+J6jBqG3Pplu1OH+1o4RjT9dhvxVSCYMF/4jP00hi6
NhTWGmaqcJX6YMYr2nYvmwTTkiRol/nstNYRqYyzs4KHr6Yy4YzJxpigV8lm
Gu9yKt1Ov0dy3sedb/I/fMGmU4bgNiJtDdpsit82HnG4TmeNV9tvJI82zYuR
phLRK3Jexk20lUYPPKqOcFChxpApjkKlHP7U171ylGfN0KgaPylsV3TVd844
WulFMeglRD9sbVNn8wmr64DSeX4+Vjc5T4tIyBwTaaRi1vLMFyeYloOs2RkS
g4c7H7siBgAgQAWQODcyKfAk8ggtRmMi9032FLtSaPFch68cjVEXmRSQQAt5
2Iz2PW7vyM/NE+rJv/b5ONAxIWAyK7UHtymuYgBJ3A27kyktJRIpXNlGsNn3
irIhChDKDZwdfiZ3tNazZRf1kk+3c59g2ivCfLFRHoSQ/yZAeFSoU9ZXjar8
uHdiJreii1FHBDDPQ2ceuLrbjH6Ivd/0gykYwHX14qs5rPVXr0diekzMC0mS
K6CnC0oONv/liMGBDQ5Qv6pd0s/5gBj2ZFG2inVaGDOUhiCDb6hbTI77KAEz
ElGPruYRZr7P9Znq4jE5wvGEmJPnubSLUxZbEgIz9qMg/hu2iVcm2aHw5Uro
iUqLxINmuIUFBt09gOvFpj2zN8/3VhOPtSCD34BI5kGTJWplatlHbH05HR2p
jGjGpzzYWRE9uMvF4ElRnvpAVFwAGjgzYC6++zuasTto9Wik/0h/bquwb7hI
oB6eBGhJi9ssAw9mF8xG9/R8UQ4t27jbEtcah3To7QkEX8vvwYQgxtu7/aF5
ONDsz4yAagK6B11cu75lvVF3WsAnsiUNsLhPl6d9m+r+sRnNnzx62tAdAjx7
Roov19YgelewYdeaS5GgFZgPTvTEP7p3KbAHxThUg/3lANUcmvM34DzNdPTK
eMuoCBbAcAVLjYIy2ut6z5qJn4hpQUtFldmwfoC0sqqEHaIjdBMWmY+U839K
5zJ4gS4UDGZmXuHauJYPfbbnzzTXY3jaoOzKFcGR2b16YCnuFHPcrA4I1VLN
mnT8nccPcBOTjZgqCpK4dc8QyF6eQVVC5mSLEUsqUqlTfQIaXkE9efBP8PW3
+e8L+YZZ9I2zPVXpfsGTqKhQqzOGQU/UGkoWu+g+++hSeDadLjO+QjASSMf7
JVsRpDBkZo7FBQnQTbrwZEQZZQ3LVrWpvINix7AHVNZVyCwse7t9LW26+zHQ
efdnQrrhvJMfRwuVoVSxMCBjOsa4xgHI0AUj8yP3bjiXnsMDHhJyCR++tKh+
29DwM8hG0pjgSfcXda4hHqLu8LjSD8ptzy/ZFcRstXNztUiMXG2xbYu7GiNh
lNOJg6Px6qq+KDsPSYQWl0ZeVABcgc0z4R187YEg63dx+Cswy6ZqmDz01MT+
6GDQKtuM9J5fbHIcyaKFiPMkHYbN8ZNxjqMRRqUpXrDviJT7JtqqDRYq7omQ
alIVoG+bDZSBRz4jmXl/EC3bsU3cCjvT2UWjEmRRXKVvKgQeCipWEBzoHIrR
WUej9Drl7snHQaHeSV6PZkkongGX6DTRj2A3jwTnCid4oq+21hZt5qoQNzw/
qNBVA46zHa+ZiqLANLIJS8yHOFV7QMvYUy9o+s2lJ6/kSPgyxeQ64rUscKCD
+qeW/MVN/aMzNkQFlyFS2PJ/+992qm+RlyfK84H8FPsMBZxJdJXKZDKIIKxh
eu4sQpYNG2/bNzy4aJRX5K9Y4UqY6ASbO8aH+fVVzDB4WmoK9O7t1JCu2tEG
/2tagRHDH72P1VXLEfEAgmx/oT7t6ZnTwdcETrupd02Joj2tqiUvqGacjVbi
cklPVx+iafIqLFg0z9LCsB166zo35F6VhdmmiPabdHzjeea/zbx9B91oUBns
vC2dmz8Cr7dOjEOk1TwIrY7xHY9SI+o98y7vYN3oyyor/m3OBuVuIjdccTPs
8DFhTRZHi7aIWdxgtw/VavYRx3MfajmXpPAfYPcY4HJFQa+MOOFR9S0k2bGk
qabYBz5dWjl99bav/NilInQwKfDvEDBaLZ5D+HzVyE8/KAa6iCHsSIaR/szj
pnYtvTwqn7ktICaMNPsk2rwQeDUL4ntr08j8/1MM7X3dYWYIufcZOri303pJ
0olQIyVsqjuVZiLUmNsXyF4/yGLu8BJ38DLxAojrEY/JuSgPrs4l9MC0HOoG
nE5DMUC0UbNUYVs0gofwF3eHmvsf52KDbkgZwTiUr8ttUiigb7evqKLyzhvc
+33gmuwdXW/ED8W3iJ4FgYWMg7RMajya0qt32QA3C7FNoH1BO1iLywEJAJHN
7c6lzEJ7YKcmycyPqdJn1wGZPkn0sqIfy60ofnHX4tVBpf5sKa6UtKwOzBPp
FqRFpmzzhv1eiYgQExnCf/crbw2G4lLCQm0hcV8fglPkjYcA9dxmA9b3rNuD
CXRh5BDEaRCh7Emm9SCMGeH0ehcV0xGX4JeaNLGsc79hfEkxpFrp9dj8TL3B
hnZgCZnFYXVuSKwtlmOmlqNfbiTuxhuy7QGT7zoNOvb891r4eeC3vvGBZPu8
ZVB0CQmi/tW1DgZUtsR6rcxJqWEHbWeBKYfESGhWOR1k5LMQHooBeBj1z0QW
t43BXHThryPMx6BF1AQySnY54tRUUOqiEXSybA+sMIbh3lhZOO8794vKEBxg
qGgT9sWcuIF08F9dtnth7R9syzidaKol4EnzWXOQvf4YNW4ZLTKdj0otWmhi
6sBtRBHbQ7TlO+g9dIYWCCml9MPjutsCqCYB6I9SoF0KWnDZY05oC7/AUqoO
Hi7ySDFrH04LiVud34ClAhsEZkJxiOgRpp8LeVadO4C+O1ni9fAie5NfY7SC
min8Nhr1oZRMsHkpZJCpyEbfLyKMec1UIHNORs5VZ+BI5ijWTYOjL7WqGxrO
VXqTk4E/qxyvs1sz+GG5sRWWjJ0tpqkzFN26Ra1mZkrZZqTobYONL+d8DXwG
AeyDJWB7yadGckD/vDicyeZnVX6RC3I/r0YXRMbND0+HbszMrLm5Sz8PDIvJ
f+YkPdOU9/ml6XiQeQorMgfM2gkOtVpJ96dYOk8kF3qnDW1JJdgpqe+G6c31
izM7ov9MYFFuSQMvlUiRVYxLYPskAkfvagYoFdjuASuaq0etaO4mz3KzbgNK
i5dDZ5mtaWwX8y6+ewp4/1GJE87eAP+EfHBeeSUxdg2npkWzuwvBJ1i9NEIp
nipWQzKcxi6kKlT9Rfy7VH/AInHExbE/zwHp4c1epTkO18ScJfsJjNBIURsd
NPP4K4/rAGSWAmr1iM9IPWjPEMToDBQx+3QUX1Cw8BblRNc3SyIFXHmw5oZ4
x2ZLNuJXbEucpHdBSnQ7cxEj3X7hgFhA183MAoQ9I04yqiu4Jz7yAlJsVwU7
KsLpejW+w48LxAW4YE2Hk/yVAG6DTUqntmwIZePvl58cKaNYKGwnB+2yAtec
EfYddL2DPia5Eg7X71FWVZuIQ3upNrj5YvG2cp8CDbKmujZqkyyHwRzbko9Z
gLJLG+qNAEcVD2NCDh5Ew8ruKvIubLyPoUC0m3mPHg1npcZ2cBsMrN+0MeCV
nCwSaErvC/EjZ5j9L7j4DegKFRA7yWxJ3fkmGjGq3is13c2uiJqO5z95MUjJ
HZ0yVT9tysRoqw8eG1ipfG7wG9hwXsXhKWV8QxmsGN1o4/Xv0SMLmrxZhQpG
U6MRVdQCICaEDIk4Ni3kdG3t0/fBKUE0IpCZBkxB5cILQ9GMmS8QZ7DMWK1H
OFQCW7qeK6YJpSQu4tZi2b8376DAO5ZXvBKLFgs8gNcE9wfwx9FnSLgdqCiU
RxFQa09/AEHiiqsoVGAD4uEtpWzx8vjo9xMPx0qLyuYfM3lfKHu7hHKZz3ms
KykQpgR+vXXWv5rRLZJxm6HdMXAFDMMNA1/zs2d4RvxnRCfiCYXlRtVbtBEv
gW4fbBAX6NmDoWz8AhElU1pGJuLRFM3hroi1SxMnZ8of1N1GncSFphu/S7Vr
rAzcyXsNGgk3pYCm3vaelbzudayhZ+NFs5E14661D3hZRtjN+lC7JMiB1DoK
NdoKeRrtcru9n6DRL6WEaMqwc7bLo88HJARLESkwmGzbUMH0ijJuNxBuBICq
5EJBZkoVPleq46O+e6xOGDBBKGtItnjMIUdbVfS3XSjqzRUCs0zWvpdV8w3O
T2oSE892hzq/OEKzgz5/sqY9L9Eta8RFBh+Y5+4xAojMhKhAyEdGs5W688mz
Lln135tRfnv+oYf+SR9RolIh/o41dkvUcdKO/NaG3xgHpWmizvD4ins5C9Te
0UozTpu9EtO5Axke6qWQskpNRUwbHRaak8hO1Yb87HpcE5chueB49dwWZc4C
v9+T1gDFIncs0NwoCHrsi+S97RB71cdUsvyFAH+4raNj6CCToSvTXP3DsFGr
NYnjbAIcw0LW9UdYp6XBFFzc+bcyK5gaNEquo2j6+9ymYT0trB7n60jWzZ92
SsiWK+E2BG40e7Xp8P6SlE7TMUFsoPRmoDwVPRZueOouvsnlCfDWPKWhQYWC
d08k7eGzB4Ew5nrzxCsA8YISMnGrPkrPQZ8peUVXyESeh+o4YH4BVFfJ7Dyl
3giHe0bCACpDtBlS2IQyEgl1aBUIZUJdePzky2JlhO0oAelcC1IzWMWZUZ4T
xN9PTlZThD7BJUScoLgPF0xOzTymsAl0dnPqBDs1Fje7fQ84zDRlDkxvqA0v
ZxKiiQaEtfS0SHQF1NLPRMU81MlZHEgbaARvHRYxJNoyGl2skhHxJaR8rJSd
dV8vZZM6Mgs2Ij7IlmZOoNBWWBJm2aUEElaoi28/XwyPENDDRW4ytrLMfHmt
FMysQL0CZLYNyme3yHM9jtjbT6moyA5Za3fzaD9LIG5qky3kRZyEwFBIQNvO
Ua884264qSAFV1jfzLWJHbQz5T895Vgz21izDs1KZsU2wKI0rnHcFe7N9LZ8
OB0RhPNaHdbRFlKN1NIEUi2NeGp9eqBKNTfHfYeVpdqDJ4NfvpqU3Qz2TM7S
mMTTwY4fSo5kSaio8vyiT48VNGR7Z4jdqy4Yb1jTMKHRY7KfnaRHFJsetU2P
rhO4Zyjsm8pfXwTnxAeaRs9JDEgs4ouKZNSQWbl67hi2GPKnQzy5xTU/A5XT
caN5XtJqcEzg0lqFNO7D1cFaJ6zx0y1zdI0TF6ZxvPYHmJcSGRZr37igBnap
46qCfsI1ffv81IDELwDf8gB9yMdcCpUxAWbwxaV5FEThUhKPY+YVyR4xheqc
quCKJe1cXLl5S94BH7ssssfKUGXHEJpmmyo8XDIHxclG7iM/G/gwsILBt4Qb
0Hf325TLz8qJEA7F+WuXWXrg8AwJkT8WxAQrjT9pfiLK7t0tZKqeJ+yR65zS
pBxj8gGgyqUTfZVC0KaRAinViLjZ7V7otvfoRym01IEhiqBPP7TxW0x12Tr9
H7SHy5sxsATymyLmAxiN+r+3p2J+JIq92qcqL5t1P+7bgGXqOb5a1iMxG1jN
pWw6q462IQlc6NfLaHmIZdfcnEA0tApSk0lfC+6uSsKV4Pak7jVPIOOLRR3u
IGo7ACmOEIK2JdRAS0olteCQorHQZkaUXC9P80FCuMv3ivLewF7TkQLyz36G
SWlEH9N3PsZNkfocJxexmJDlqRTHQuo76GsLQKI3tMLyOC0ndWh+0jkWtscZ
3tqSE1Hm5vancl4Qs4wRPegkTgRNPD5AwjpUX/JOimKif/PIJ3bqyMb6rhGf
OqdDU2OECAuyw4mKjKduaY/N9O8JyoWYQtd0RhQBOTv6BiYwAVhIZTu718c9
2MpHhOg+PbZeOrdJklZURwJkoUqJTEfSaNmTctX3uZK2z43vol7u/LwGXtro
vejThgxGoC0Xb3d3e9plPpoArqXSlmGEV6p78+9sxmmaMEmhH6ujH2Cl4YqV
CsHj+DlPzoHkAZCMh04dqpXF3PaSTLyuDp/QJXEC75LFnfrVJpWmfSjYe1iN
DrAxEn+2EQwS9co5nMhKk4KYnJ56UR1oKzd+jxLRrVSq4Frpw7WWrlgHLqQK
XNq2aiBeCQR2MqJLhQb4vi2LHJDki0RGISMLDLlqe107KjDAiuP1QcYvDEKe
E5u736H/P9zVvs39QlUDrfD+LNKe1fdavhEJtLta+ElLVUS44kReq2lHnFqI
YhRPjEPO68I1Efni6MUYqbPq3mY8FXIXMIuvABF+4gve4SLhBkHad1zkErh8
/+bjyLESQO5hIbhqsYDfAi+Maq+tlGrisvAjZjRxYJD2zU0zF1ixBGZIoamG
2ie4xhEYNehgVGHzg2aB+/OQS5ODyWMRyUp+fUZWPOmI0YftoEmobYLm7ovw
dM+ucLuVmZ9yLFnbeVWwojx8zL7VCU+jCKtCYiD/6LklTCiuvJVW92DwNnAM
eECHA50ii38UpZ1Se5c8LJZ3jSFyoEt2k+eJ1nZGGX0iS5stN87z4vRuy3cO
g5RaQ8XlItA8BGqycOSRfavDbNyPuvQ09/U6d+98DDvqCK6VQchNYqWCbQ6W
3BiJYIi/ImmCq2LA0SR3aWMxqcnYum71uW9FJYpO0T9V3X31enJw7jfya/4X
J1LkntJEGBE90mq4ZSL4nueFLhdqPrSgTin8TnYG5ShLbEpVuSOVGcde+HlB
+i6ylQNW2wAlKFdIXRSwCH9rPBPb4y6gAjqQHbbWQO7xiyr1EwYWWGltfHRf
t8GQZPD9Xo9sXCsi+HpO7KHFqhqRiw0C3QTyAjvLCTVIpeeDPBY3m7URs7nI
oyWiRPbKHGo7FaKc+sZvQrFrZhyec98PVVr+vWM3jj0zsiYz+eTfvY4OpECh
stAaaJgsexEm6MJuNc2vFp+K8Hb059IATG46N4+sqV29uYLLxuj8SZo06GBM
e4gmPD9vqeycMMxe4JzQpWwhyRku0OYh7cIGE5bBXAMa6VEntV9823wvjEhB
t/5HfAAslN3WPaUTTmWqYT2JFJeThPb9bNKMl7wdqJhMSO3lkmj5V0M1iNTv
f6hXM6+FAh7g0g+t+iGSK+cRi1xQOuLPAIu8raenWuwBfODV6wiga+JyR29p
s5HCgRTUeYSstZWG6RmweQu9sN34pEuPSyEdZe7d2aMQbZ7QkugJLcea5FxV
x4HwlkbJTucqhfI43H9179YHNST0yLpCpm36EUmhOHcr3GHqXHepnJ1GrK8I
RwRt2e8sHaFBUHOr5rOekVjTFTUj1vCZo8dEgFoIVTq0i6PXmfr+37VEZwYN
sxWDlh+BnCGBg8NLaUp249D5lEMw5oFYNJDEJqjEgyhJ0Teg+3Uq7Cr952f0
/WeLRe535WQG+lPOQlI2cg77ygr0c0dYWHixvlkarH11jZZTkl83JbDqpxZR
llsxvUq9j8cVXG2zsQlToRBTKu6t2Mgsjvl6c/Cpu0HAhrEEk41zjuiPxCxr
RDwOl4mlR37/Od97R+DkPWw+IQpLrjfE8v3f7GskeU8cBjWDsrnFUrH8N3CS
nk9+4lidqAIrZZ3RkVHgjY9QEbgeWu/SBDYrrx0LvtsBFlhBf1fdHsjCJc9x
s9mXFHSgTkH1GpmBCOZSI1adKU8ULYn7FmXUOBWVkSYte+fLc/DaLqbwVcsT
+ex9agj2A+nPgUGlj84hP+PhvHGte2/21Ssot3qEFznUUbYJKq6Aphd5cAGp
qlZHlxWrcTUrzTp17sgqzqMiDmIlP3kgzTfkyiFNanF9ewam2DiXpkhz5o6W
x1l6gQJgHbh0wRKVPdF1upJ6XdS2wRk1dxgaI1xjRGVzXLdobwdcB0md4e8W
1+3pf0B4E5DkEjjHEOeTrdGZP3z/GSngT4SjhUvkfRRbs2ECnVIfAGPvR9pX
I6XhSpolvhNDAIMvoTAjpJVFADQOl9lswkRalmBg2WGPn70mHFcCe2CbON4p
orwFS6rT3qIDSYaOjNbM2JY+DdZLrInhrcD32hBhe1bV9MBMz0OsvdGzyZwi
ZE0zZ5HWTTzELkNa094+byShTqDp5us3Nkg5XUS8AZ9YbWAIrEAzCIhMyBVZ
E0XlIJcwhbKpdEY0eripM8yGOGD37r5kQLBD+n4CIBvtB/qlV6TrNvCLEn2c
2JwJ9S6N5CVmG9spMKk8l76q6AtocGpyFThvTczobs0FlEvkL0drwWIe9fNv
tTD/yjCT4Ku9fFygBUapgIeSHpJkNkFZqYyHfejAW8U4GF/hLr3Zu2afFw3K
qlkMjaihVjdWv4av25zONuqOqvaq1sPZ6Il9jHI+6Vo43sHcoNkMQTPYDkN4
ljfj1kZO5c42GSf3TSgslWYp+f6veCcwfjnOu25e5PZ+UADJI/F8v0pLlHvb
PKCeSpYFQo8sw0+Zwzg3fsG/JYHvdr52MLF+ODpKsQqDWjWLXv2cl1evm5w7
85mQqdoJAFC1AX6wXjgrZHMBo5RLfPt6s414mNGcyRe7f6H4x+sAMDiqSqh2
v6mymSIyvnPCn4thFz9mrLSi367pIU3dSa5V1FGDMI5NfFvX/JBrU3JCyl0u
Pn4LAuNYmaKrK03fhLStw5CF+igg6Wp3WaeGN+cu+u3cSd4WUTFVT5eRtQ+P
qKZeOO69gbvDp0ai3HJtt6VwDd5CEf/SJea1N6vvDSmAzevM5KgSKQEV4oFl
bXXnbcDSNp6BMs/uFkLGFLpj5uq7VToMjYdtgoe9jrDuzwZftTUmztOnuFXX
QNVjVepNdBwJBgc600yFeUWUYt648t6pZnxRg4zGg2HFd7grdPUnG5pQKB7X
r1FTRFhWF6JT+GFYgDVKEQLw/NI+KhpJ1kY25LE5SMR8z7ujOe4QDYwVFPVy
f/f2eHOzxNM6trVSEb5gHy5KZ9XYJgdBbRxKN2zQI+tLAQt6FV3xo9p1/CEM
M5vhUd1MkAt9vxEBMJTxMELuvlgihCsyR0XL3jP7iX8ffrBJ/xY7lCFqqpq7
ABqpslfK26qSBtn3dw6TipMZPyDNC+wNbC6Ev9qZ8l2JxhM3xWBl/NHAvIZB
aHhKppYipMUa3KN9y7Jq1ZN7I0Ro7znrjjXLq1BIdJAY2FEmvXvnYEFmUwy4
Re0Mz/4X3O3G878eMmD73F9Btu01VODdOAt6YXohwSWcUL+XMe/UTWfyI7lW
qQ5uFy1U4EbRfDh3vIW/sjxkhH6xCrQSs5NAQhjCtORgbKNvUlD06+Nai19L
6GUxNvgW2jfE9fyIKkiKguceade9o73yLVdyb3r2XtgS/LnnWzR9OBScixTo
olZQ22WABs02lljQ4FcP/yKIuxNrOuWYgney7xssvbrGzyaFI1YO7h6/Chcr
a8WAgpM8g3g5Qd9PDD2nj+JAW4BreDj3WxyTq/Jig9VqUcs15rL0uaW/DyIu
CZ1DQRhFoHwoerQ4MBLVQwgdKRI8yvDpEy0zpA32/9MexQZTqsNVuFu8MjeT
v6Gx727tupRUUeCokpMZUuNeM3f6MYw924G1JX88HWtPTOM9Vbtsl1zxeuSY
qZLgFVFA8FwuF9tOVsOVWbyE6zIY0c1hmaNKfcwF1HsNk2FrOP++Bq+IBKlP
osliSjI7WQS5dBoJ1CK1MckgbIKOJ3EA4HQclGGkquXjoH51Mh0xaSF9IbCb
b5dznjdz0EfC73sy8ms3mFzkM2/JTo4xFjBCETGqBMWFlqnfIvUhJNGFUkkm
m6RWJxuRB8ksO6PMEwRLa02qtiXuv2TJMYwMdOVy3MxSQHfdAcjVIMH2ualK
tD4q1iw2y2y1mQOvBNNtCwXGFFjCt/l6/6wYSQoIEq7j2hn4xSlgK8vZpHIQ
uyYuOFNbGQqqSus6DQhsDiqEUbwNETP7PYCeJfIZohzzK7JZCGNwCXKS3PZ3
H+87yl3CXJyAl0C6zSxgcOEVLo5dvI0S9RzPXrQDk3QbPkxzJ2dAY0ZixKLP
5DuHl4XZORiAft33q5CpM7D28aElwXFFZJQLTwpP97iJcg6mpaB/hdJKpM9B
yPly4AjBxKk5RNpSsgHmMvntWfTNVNqrWutvOBAeNJVms4SYC/nAGRNz67l9
2I/YZPYrjR7oOXgNjrrpf7k8zr2uNsNew2oYklLdyxonlmwJtNmuLrrUTYlh
0TQhZuKartonSC1LkxQ2WTC4Msd5uvKj8vtHQBoNxQPTslZIqXV0H8nNlOHO
+XU5D5TuLLb6zuUuPEPHJqd2TDiWIXSaTLldO015UUiw8q8SDUnOnDfLOY6U
EnK8uDFFMIRnW6Ou5N0wQ/thlys8tQ1hsrNVn//os+/GhrCmvAN/7njfqozL
mBHbqTUPeZGbRmd1I/HL4B1lBudF09lh8vv0pn+ENMs/P4Sy4m1NoGvVRYoj
9woGrpM9BUNtXnYPyeJfM6LS8TrEJAsNWsIXiY0dbw8u+aY1juse881NH6PY
25KYzFlEgYndmEwbBBSPfs5dxVfCA8/CZRdo/nZW0fPQjgniBif8qKLYNvAk
1Ovc/J6xx89mwpQmatPNEvicHTsVIbOGDDt6DGRIa4lVtMQAR0toaGUL8Mtr
1D/g135E46eYWY4UyIHF3DQne/PjiK74lf+qndmHXvUlrRwL6nla4Km3eEya
EoVYh9KVGmdW1krY+do+Ucf7YIPzwDLKWmTgwdR5WJJqSku+h6MOm3503uPG
fOsE4TJHw4HasZnOBoFSTmihAmWDUB7pqEUlpxmdibO2y9YIEAWkY/wGJIfu
5PZNKb+9R9/22pQlNL1DeUVbZ+dfqpBr8REKTm8syK8HmAwA1i9YZ1X9ePIn
s54TjTQ6cqMUpRnpWGafMGzz4+UB3piPEg3kgJVdPXJPuSvTxX8CMiz1oC9L
xvVbAb7PIX+ynmaOgNaaiS1MbndRkaTwbAcgvX8L3301THP+Sckj4QD+LjtD
bUcAZNQVoFcWmMslA1gDMkXfjS/Bo4iljoJwLMWT88J5UOx4Fyt2Zjioq4zN
+GXAcaVKDgW9mRX01vzS7EUTTpDmmVy2Nj7TNxb50xNJlbAHUsu0ceWdMWpu
9O9HRIUE8N4eTi0cn8oPAr28est8zqbiReP7Ne7VYTMkdw3YS0M9E9s3GaB/
DNARSyhmGkFwRIk6CmfWOm6+LKaRsBgkeKZbFs2kM50JXi5Wmdx6wQmbMUo2
79uUKDIOSpIxrfinnN9V5slS+B5tPF9sbbClDbAFrYbPFXUU0MtYBXmc3OSK
6yczjB4pdfdXwGCBou4hAJDCvFFsvWNgaYBSMvo8ovFUcvq0rXGuYMR/1/EQ
EvhZO7unIuPYfGo8ga+Hz+4OBzOriyBYEQfnmORSA3vGcbmtQtD0IrNDsXiU
jYzQoN+goWqh1Q7CV50/00NTxOc9kShD/E6zxK7zKGmz2V2WU9Ovo15QnugE
5cewr+mEJtkiglywI5Wpm6JreNFDPynOUUnMrxgSmvbj1C7i06jQHetFt+Fq
zaijPp7k5J8d2vjv3tmm5xCAc5mBQlQHiPD8BEWyANUAFD8kRj+9GAJCZQTO
RqMPLvgtPbl+QwETWiJcYWDgTDaxv8qH3tiVFmL9XLRTT8uNhRu0doH6Jr1P
7fZpFZBTjy5l8a4v4UvEhHuW/S2SQBog6wuw2NApxY3WhPD5pp5dyYJkivw7
tQqmzTMzN44HQlfFF6taCt7EiTUQtZSrV5GiZHDi35P9Qdg479q+CKBIw3Yw
GgiHjxgIiw/rRf5ca9NoUn5q8emSxV/CLmrcIoAdbzW5L0YTBJ8mOI+fhBjd
msUR9lt13rYulLdbaY+64hwNfaaQJn+gQmM4QPpZUBleSWOfigIbYyz0kRwd
9wFuQdvaEvepPFGoDy3YL2RKg2uXY4Qp2I7fI9gB5GWLXsMMboMKHpgyKwFx
qrSKmaoZ7n19nUUW6YbvBPEPjTih0CFkXBZo8lS8DoAWczMyH7VD4sT1nTJn
BUlxnP1hKzE13mLclkPDyHs3jLrXDAZUDGd/BRotEKn6fAo/FFEtRKLm1Bj9
fHQgkLr8yzhpL9gzpttjTeR69AFqIJl6UgbJV5CdyRIH0GLRKEFXsHPi1Jm1
6WBP6+Fre04gX+PrQ8ejBE2968l7xl7gpVe9VU7Rh3Z8e4LHPKlYTbq8ikdo
Vg5nzIkY94h3HxLGWQaGrxbqCNr49tAPWPptTpLPTubHJLkQeFE1aVpeVQff
gxBjkegxVCdxXemz0Q27NnxfKph41Y44c/eGNGzibJl58i5dEUQih2cn64dx
RUuaAMhKV5TFvVZp9RcyYpQzyJpxraETb0SYO0UaQbGzlkTRGjmHSHUdlitC
5ttCV8za5n3ZKlW78ZR3OLVfXE4NOEid7FF7oJ4Sxf04pjaiWIMtMMyc0eUm
i5Nf5Dr+YSTcSgN2fLyMjqDgSVF6/8chmtJ19L5nDa0ByinlmOAFmSRr45SP
y1Au9dU/CznMqI8x4q5YLTTBryKWdzGbHTJ51TVUGh8pY2YZ2Beom6m0Ush8
TpVWD4YDBLyM+QZOgIb3aPcY/7TMeJy1RG7o3FmKwSJ6CX8ueiF9SjPcedPu
Ld5xBnEUE3bQGmMGFnl0cbPhYugLBB6i1ASgzoBG+unfNcrSFh5T4zdiC06E
KDdijBcySC4vC8d5sgd9aByftUvY0bS01EMqeSwVoEd36hrYm8ED7zsYy2HB
9SbmkLxgOr29cEZaWwgIQc62yD6f37GmOoLolkpGbNvhOPqZclnDC026yzOE
csqNNdcBOV5GzQBoDA6IpGXcl0PsCLlRwonyvMU75JHS5HDHprCeJpSu7Ull
y3S63vRG/SlfgeLXLgSLMI/DQ5Znorw64+Zg8v8Xc+MXv3JWkSakrnJjspbA
E3GMtZWwmFytZo7YrvC6A0tUyORrIfvbDcpjtFB9d47vAUreYE6wn3NOd+b3
ehMctGivLra2HHzja9ydhQlJjMMm7eyAMZbGbFNUzpareRNDMKPLmqrkO7ag
ojPreDo34uDUuAIHcgGSOuBiEvIN9XAfscjQbuECyVEgd4R5kG5tWwyd5n4+
vwN+6+gIyJGH1XTwGQslhWOLGfPYkuMHIkphTMm4ZPBASzfSdkNtzmQ8hTbp
CvyE8s+3cas4MIswFtX/nC+npoypQxnfDHuD74CLGa3e+loi6DOkwzIUDKMu
VGD4YBjcM0jSgM2GI/lPA/pLV2AKEihEuzwznCHejUd6liCOaWuS5ZKRwf+O
tjvxc1EmTQDGt64AYzwTOu8bR3B32woMZiOInsqlAwmgS3ps8w79/KlUFTac
FfzI3vKubLeXeXUunKdpmUekVXPM8cv54yW0YlUzSngYZXkzFnOXO+HP/7qE
SpdoigOGub5WbKznTsq1FAdRFuTZXw6UMUAgKV4SyoZ3kSRs18e34GWdyCIX
kguzPUOn5J8wGGAeZ/eTLT7j46TPQi9kyqWhC62h2Xei0bPfdGEAzHA8pmgw
iyc6Jf9Fgn4AvWVX08VspCnvb/Ax+h6HOLpV0DexCIwO7uoDF4QsPTLBRQaM
64hGH1jFDoHUX29y8QmDVX+Wx8bHrWnt9nHZVRVOi1dUwITm/xT8R7BcpJQR
4d756/OCPDZJMlVjnPNEBqvCXJmrUpyLJK/vocWg6dWoWrcCrjs4FLwf4mwz
rNYG/2nMzOxtkmYArpxo1kGsjUbqVK7KoZFvIhn6M55uvdzxo0BqXu8XqPdu
8QOazr3dq/IcYpxzHnboM/4343Zr7Axq5EGVkEBgPZETSxEzMAUHQLuLsFaC
66FtxIy3wc6+MR5BaINb0T9F/Nyq8wDS87LAASuD7+QXpXJw0ehIKLfTm3E2
jepYO+GnDYe4TTcV6s2BR+QmFuVxnXFJi/+k4UzERUs/nhSoLRUbcnHJGkDk
ywannvwuE1d9qy2OVtlPMcXHoBw94IVMecUBJifN3vd3RRxNfEBXgAq4EMai
jtxvNjZku/ykcQ3iWLANij/UEzkc3NoYEL/496ByDXmIOhTXfvYmwqSqA7Uz
XXSlSdbvQ1wlxnEr+X0Ajj6eWpsXNN5mSQFd3L52C8jADXNP46995t/05OnZ
sMH8lr8Wpz2qCDridqHiKEN9hjsSH74uMYAp2JUr8roE227+t79B2TjBtbhx
lSO1h7vUDi6eBYdN8En+4tTgo/PZeEptu0zx2XRpGjcoXlJUfhiOBtxA9jB/
qCSZ6Ftup5tbc4BCu52oThf1KzYmpgNRCtL4UNrowCl0M7ygVp1aK3ivCViU
ZsaYTOWxOARuIak8SokvlErJVSj9JQkcR1UwEIcTL69TrGNqpfXNHLfcUW/I
6FN7bBsmgUVpwubj25kRKT4NYp3beJ+jK0248X3xmgEW5HrVTj4BT5/eV0tk
Ajqoloe/p5fc6hz/8kvtuV1Ny/OPXbnsR8oUqVRTI40ak10PXTb7yoEtlvlq
yBFUwVvcEcZb8ZOoyxzr59GNxrtZ1cTzhc8fagHS9lhKRbZR/uIAtzLXB65S
FnK6kjPM4on9cfn1HVTG/8b9l1ZjkHaVEP7KlYqQu/H/AzesaF/WYXeS9VAF
vIndvohYsk9P2Ot1koh8ZdDO6721fDDSGF1HAZ/OyT+c1K3ZCglR8aUltJ5G
+k0gw2a0QBX/UPuqfibrFFox+AdqAIKC782Y3NeUKFFRDUl7A5uk1JXdL3nv
sP59rkvzHXFFbeVhCXrKbseaNb5mWOgeqBhiV7o/pC6oo+fFw+zNjR94eRlt
OtNsntq8D8HBGFhdt/uEncw+dEoEMAB4GJ3RyJlPe4KRIK2Gdgz0T/5qJhtP
5qa2USmL278OXAVFzyuF0GGFNn90LJqnr9M6GE124x9UP7o9N62UP1eT5tm8
StVLCg8DdB5Hy/efbGx/yMdxWnacVXF5dO2kWthLUHPftfTx4Kbj3QyPAujt
EgGFSTSTkMRxqvzFKXr7U7WzkOUjLSHZDCuamcYONV3v/NvXn3lRwKNGLV5/
ZMosoeAHkVHT061tCyxmQqve3lO6k6pAdB3fyfQSvOIwPlQZsNkx3O7NPTmp
a3cwDyOv1VEJWrBLi3ENh8pcmuyQIDv++DHmUOGDeweR7uaOtdNGJ7wOzRXL
uua4B/a5i77momtFRP2tVlWQv1NNVU+nkaO43DKjtS/WtvtiOty15SiYcQld
4rZkl/2fF3/a1mGdd7etF+zIDe1XAbw09BsWlZ610n+2t8UjJ8l8EAY715Sv
YNrKwCTlbrDXge1WC5zRjrBohc5cOhQBo7dGZEvjmQx6Vqtg6D8KEaFnnt6D
9SAGO6zIQcaO3pxXpmU9YuoBhCD04ENYHZX/+MvYTTxCCMhOodsEe1bxDfZB
ds017PX5kXpnwYQhO+yd7NJyWSPj3DSrwgc8OIwPqGMo4tJE3EZjkHRTll65
vOvD0mw7bjwGl+yfeBx06ciVXTQb8wWALBBzUx0A5CZOYS/YWf/JUyr3vCQv
R8abr11DK3lVxE5qRuWVYZcwfr1cBtckidEXP/3rg+9UPT0uXlicHSuuMYg7
uhlr/Re0C1EjnGSNFsGgHwAXsdcUZ6hqhN+OA0QBi2p5EDFWvsLniOD8mk31
CG/wr5rtLVNi94fRlC55KgTeOu8d8C2eOIRW6EfLuVR61Yf1P4A8tsC2btk5
NHcaRQRfcYG1eZleGCe9KU+C/LKl6ztHcilpbZGUrxwhn+Hk4lH4aBGvCHmy
tHctunkT7lWMpmgHEIpYdpCxMOevDxPK8gr84i68fDyj01Mic2+ueMSSPwmc
0r7M0Dh7sON3MBZUEFsHw/zJz0Z6X9IXDZFZn3hrJo4vn8dZTgImwEFt9fbP
QlmxEQsdi5hC8G3QCCEu4Gd4YXmBlJuiXZZgyF59RRyXRrv0NXOwNvv4RAx2
jx6OYzCn1Z8qVrmLtDKnaOFSt92d8+qPnPYVCFEUfGgfZMmk3KU2pYHlSKD6
7cxn4zPQPrDyBOwsPJnXu4R0OTJity3CXM3Pwjh9TpQHKvYzS5EXkMQooqrR
QQV6qGocQncd8hjR9RzxVXeBGdQbkjkUxQnMj98QRE277scx3awDW4nndkyb
MeRbhTTTFlk0mErrZCDXrUuMzohYo0H3xHujGgy0Ktz6Hl4hTEKKuZXjSbeX
HnMAp/DBlzT2+VZIPR6aPXs5V1dmTK5rcgGIbPZUqfjzSDMWMz3r/DqjDsSA
d6+uxKtyjZp5SKxkg/PyvQCjz2NtV6JLbcSNPuEVCJ712rNM00fvWVT1/Fvn
dMRMCCOd+ln0YjoCN2IqIONhYeixztre96WhZe7NNQk+BVj5B8XNYsAGmzDX
yNschg3ZaRAXGsd2uaoy6tH/2nLy5vEh4wLgZilrCLADjZccNxdnJZKMea5F
oxk5OtChEHc49V8OLkSyxkec85kFy7DNRh3uyNCTiRZvuKM+6EJCqUhVoc9Z
BI4999JyAGu6DoVTZP+qnFGKFmgdVp6WZta/tlwV2lhw+QD1jVYtyV3Oc5Qz
JDJMQYW72Juhq4yH9f63P8uarZX3GfITtukSJOMlj/7u+v1iH7mShtR7bxcV
WhMvcrXytNpvbmZwMZtl6A2mIQnE3d5u2T8CSojNg5cfhBdZnlWnWngeOxYI
nHqg9w5zvdDGumSkWXX5wB5R+5mmcsQ2rArqYSIkdlAsPgys094oWpE/QcnO
B/gmqYjYHigL6I3hByQRoVTSzc7BJ5LwTzcE16kSbPyopTRf2v0rdL8mGJpx
JKuqED8/SMu5J5b27YWFedeRiEkDFt0P3vamm8Zz4vO67HHzz3Jp8sanisxB
K0pTLRHIzeolj8HEjRHnNUZOAf5IkU+DgblCFDWLqOUquflogR0muNIVUFhj
H29a1QhFxu1/IRD7qLHmCphrxJea2Fag/L8SHCet9Z2w3hh8xpA0iMu3XqfU
U19ow85ev2/s+7UIH4IFYlEGJfuoZ1Ypg/jH0EpLXJcJoKW7nd0P/89VyS0V
Zy9XpfSben30+vnkRiDpy/yaHG6wualGE6Wd4Cu+jg6V6RgmH1P60pzD2xMt
1xQV9Hd52eZUAjojxIWQP6od/JVBD8laSJ+P8cuSXDwHcsOt1u9jBE1L+Ujv
KN1tUmeIEL+xtjsy/XWXJvEKVIii7Uf6KCYKpVT5wSdkjBVrjGhXyyhBD6ma
nJAhDAu+oxKyKwZLkP4VwOrSD6gUyP/CFIWwHPfh/vEHESo6F4GurgJgSxQe
30CHr4nrE4A9k4c8v52EU8D+9hd2Z5ihWomtnn6xWSxr/GXcwFPS6FbcyZn1
zD2mfLc1e463wqhxg0ir1nWTQ7zyc2ut0EcPnFtA/CsOJRdcG3fBp+gU71E0
9AjgPqmdLLMDAWm52y3jfTGDNhZ8cpULAGWf9se8tsfKTADw7YFxn7azzDQg
ZfhLk/n70twHvLq/HM6qN2VTfGZg9BOkT2iZs6EzDNcD4B4OZOLo9xIbU5i8
8pBdxPvkgOgLtjmPjbbLCT7iugMKfLR0UPUdpIms61wi5YMjeNInJTtGRjB5
bhxzRqPlLvbZ0abAxQCXNB16OVODaCSUqn472HqUJM3Qjpp4oVZb3MMfh0df
IMNSs9Cioy5T79iWe6+xodOe/tk2p61D8uCRJwjFzcYmheYlCsMx7+9tBHzu
j/incvj5Oo9wF4r+0RJpjkeHbbmiIYCql+fK2m4jvyiRgZ2WuGKLP9Mj5WVp
4u8RvpQmDUSMpKOcbIKCzCTWi9aiEzKTlXrtMp3a92Ql8Od0K9dSgA/bhTQk
tkehHU28EtymEPTBI9AqywdACb8hMz8Tu2vwrCcyAlFsyLmkABpgKC62/VU9
A8pARwzyP7qjftk53S2cLsHuajlU353osMsCXzA3QeVuOuYqkzhfF+CbuY0q
twC7ISU2Rt4ol0b2dCxo/MES6uZVLH1fe0TQaBjqx/zTjSKF71pH6mWFaEkn
evBZmspD5QOibCpwFcrGPPkyNmeufIh5zowB8Qj6FrHjEcE3JweQipeCDQ4p
SqnSJfAmp6xbo411+EzmS6+EupXFWnIhGnnXq0VF1+boNC/WFCz9j0IU/j4K
6YulwKZrXUjoTnfOR50GM6nSAm+KEd2wmxB8iJFlTfSerXmuVup0PIulxjTr
ggcG2lN7RnwDWX7UXzM4NFSb9SjqqbI9WRI7pJmcvLl/zzJkqDIq3oFGcZVm
uWMoKMjh6QmxkgFm6leR4qFFl3p1WhUT8oRFYit9SS9iTZ48qhO6QwT6Q0dz
RD3tjDZRSt5/1BLghHAUID9yI70apNaJftyuuKMGEsJ7fU+2DL0LJAFtnnzj
7JL8t1zOXW4kP4N/pwJLN2rgBCi/CDE/K4eYf4yavtiBHT4N7Fm/lgL6IrZ2
Bwt8kmcfEpP/gW9yxXQ3yHhPVpH/N2zvLUxKEiN/ZDnJhIURAqTYZkJbwB/D
xAWjehv53vw8NallFEBdAVrJ4b08Xg2suCzsIMGvIfeBL1P5VlOgV9ewXCyM
Np42mVXiE3Xr9BfMfftCAs9IulSf2bz+fet+5NYt2d/kPqC2Gu/gj65CJQBW
ToohuKULnAphb+N8k7RHIYS+RvgL6rbnOjexCeKmUZHfi7/bElKpW18JCwBm
VQpWMnaITdhj7l4Ya2fhvLzjDZptcSBPpfKg2ZzswXacvEZKJOhO+FtZ0UN9
6fqRBBfcEp/bvP175TkF+NLVVu6tJpYCEEOwey8Wp3Ap6fvJTf+SCyaYWmC7
J+9rIjEQu8OaUh4dHsPKlPHa0GGR9O8kvppimXcdxR8gde3xBFQYVkwYhLdZ
0GPg40QfzIjAmalFzILjpbqHvU+ve1zFJ+K1Y8G9nx0RkunNVK2/2xhzqscP
Sj4wDaCAKoMn5ia5IM2oo/JZ+ZPmHhMbv+X7NusOb6dbzaNdhkDe2iL5f0VH
KDZ9uPPx8nGm2gzeXX1Oih+HoDptSaXN/cSOXA6MPdwJkxGNwibSfbPRvJzP
uAWSRELijKyUlMRBTMADfPKQ+l43uzJjJV832PGCvOImblkEKXndUW+mjGys
QuhTOZkQpFApc+qzZn5SmfVDIM3+1Fq3PFYboNuuD99N+k0ON81+q+3yPCYO
9q/IzasTzIUr8QxcxBaoschQxE+N9vnrEQM1MjqO0RIyNbYs3uHJx7j3Qg9W
FeVJz1N4CJScnCsA/b6UXerKVUYIu2LU80BGRVj7NPVGUpcjaVa3OwaDHGMd
D2T9Ia9j5ITN9ARIfdcJgkqKOLxfLO3PxAu0WXmIv7CeclTt5dVhCPcQapFx
RGO7ri58iPivdRE4+ZEdQkeK4pgJOZYyKVWnwMsKX+3ZHJakt4CYf+l1GxEx
sQucbJ5BlKXpLD6u4lRwbto+pYRyfKIM9wmOitb50MRyjqYOnallscD5Kgge
m5paIjxFkBpYlz1fDzx656IGJOMB8nH85QUYO3yXSzcEHrhYhq8tEKUJecSF
EnV0kisH2dgV4zoKjZVFcPW9SwxAViHWzMKGInXyJeoBQErJhYw9ZqDHuqtB
nCA73aL0VoxtTW7xmqi08TYhmbG73bqSW4rq2WL7ANd+Zu9BR11e6mXoU6Uq
7mrhHh3G7uGh7ldF1cXczjeoAveN4n+/Qe/pZjKTgTRriN/WUD7Ot/SezgKs
kiaVHZxQCR0Y2TAa4JC1BeW5n59obbDb9ch+x/TEdfCKdSXVX8NyZCdcs7Kx
nKqXKXudFURm8FQ8ObMjRIuMpwqEuaUA0EObHFE3F3Zu/L1mnDkLB2ROaLr/
MsY3nqVccuqF0p8iliEFngSs9Qgg626ys7Y67Sn1By9rbp108tBjx5iadwZo
H6Oxw9VVOOSjRtNyzAzYZLLAhGLOOZo50c5nlJpb7Y8IJpy3Rf1L+w0NMHCx
7bdEHWHdGJ6wedMVpU3RQSQq43jUKycIfg60O0i5oaEhOGhF4bkUxgpUGneE
YkJ2qfzjc63lnjiqHFjEB2erhRuJEqvzYNAihy46fLKq5/Mm555cpK5t6sd6
+FS2i1be85kVifIr35kPJffwDQZMADKVB/lk+L5ms29gGS/bUI+Z5EjMwYJq
yf1tubJ4AC9Mv2lOmt4G+pMH59Ma2YA8hRojEmknE7OsV/sC0yLQyehkxZqv
+pJwGfDxwXgmt2YYFfn97or2pZroslcn2jYHFweoemJySqSZplKGbVe6dsbq
xFqjLLYj9x5ORdV9pv8u2ZhKxSkohyNo9fC10LPQh5T+Dt0C1JhGOfgCf7hG
Qhy563CdCs83zUoeFd9NaO7KGiPep/zXGS/eOPwtjI9s7c0kqAJ6G3x/4euj
SbB+PjUHuxRuwu1HuEk6vanWsD9A6cDS53RjD7PFT190YQBiU+VoQJm9SQO8
pedSJOsGWzzxOX/YzGjhw4lmBMuugX7TGS2DXNXmXn0YnrokVOIdRgQMZ4Fw
pLZP+RZUaXAJl5s6kpKbizL1kGLXwsVd9OWd/3+C3sbmfC/wJATm89Di8LSs
7qyyN1coyaCcFbKdi57B1at6d0z1QvTUMqmUZQMW4XDedVrbo1gPNLnn2yEU
SEXDDnctzk9AsdJD7oGZFG2hOtocOCkuVxBWQbxhgOrKYTQipEfhvaPA1cyB
AByTHwTnEp7GLBtv9DwNaat9l1iOSPKrAcjwayPc4VqK8K57roisjEsIuMXm
J1gIy6XNIOT5gz1V5/N+jBU9VHH+5SpvQq5DfKqjLz4v2c6Tb0GUX7kos5xV
HWL0BcqqNn2bUmiiWuaJ4YzB7NKklgxDNOTG+JHGD89pImzhW990WPrU/3iV
EjsDAXp7fatVyUYkzORksTmejnoIM2ciTL9i4GjMHQk6hZY8rfKqVgPnwrrv
VT9ndHX3WVj8vTEl51z5WIAKVZh6B2yzphQ79dAB+KtBl/1djOZILUHgwfLu
sGR4MJtDtoSkx2r9PDp0bJKhtUWR/M6pjmd/re1dPRaUlnpl40npqUF74l9P
gT2tjohRARPJpyZqrmd643QXGZ3CPQjv8rZce8wi9G/UXyGrnaVZZcy0Ui90
SSR0WyzF4F+4cl+MROuFB2VSW+sbi4CbFZ9K7L5lo+8PHCAU2niiLk0eDrlT
a1QN+QfCsAt525rL3DAv86/TVnUeYUSW1880Eee1230XpgObZmDrVSAscqiY
Gu4Wqc4bipnQBkM8JOmTThw0PzirQaIzA6gFWbB1arpvMjY62x1fwldE9Kex
3Aar7owLVOTuAFXl6PKtyIGmLGixOjyrkDqGnGVZi2B59rudHD244HX7o7yj
s5G6MNM3tGz9BaJi/qs2xIm5O7hbm4qobAetoifa5ca1We1o5iHAJBRD9r3B
hwplwAeX2zwxZYPNlmJlK34EyxBMyeucoBi6jF1NC5JvXnGR6ixp01Z7VRUo
S0bDCGnsCddSW6yKq41XGD3mJvbZdGu0q3evDYhF82s/OdxLs90aUc5ojZaT
93w0sB3uZsaNfQ/gKpnLFfJqfb9joHFDEeQrG84tP2QDsC3tmfpFrG5gH+hA
UpkMy89Qb1kA1WGurL8CW5e2GwVCViPSp+IvdIlwxRCmgtaWJGsq87lHf6CN
HryAsc5ZEbtKxPAC3kikCPYdBJVhnAShWG4YMBplCaU1Is6d4bEciieDC8U/
28lRpzU+1YY71DDV4kBKk8PhCeKbKWfw7CFUTtuuIaTfYVHT0KxToUfPuNAE
rv/ZQDWWQkxgH0Fl2j5OddtoW38oCG0TZekBolPtDuTY+iXkATviu6I3Sj+8
i/g3IOjp+VUsvdztAzWwXjrqe7u6ngAULes3rgmTCYoPgpNvHeEZueDfnOHA
aUx2EIdXQaw3rNLoxmujL4SjD9KGDWio2cio5HuPykfrBZ6A+ICofFGgLr+J
dQBvdrlzxyg1gAMkDABaeYa/6PMhfHMrTyK/z5E/79AiePteK6WdQngXZ7wU
eCOrHWjI9tBnNvToMvpwoQ7T35i/yDGhmP+spOhNPxtFF23/O+2/2twSei/p
/+rlTM6nCH1K+C6haYZJKHzn9eVtLXuRhwbOOR7aSQaNcO5HCG3y78siYAF1
bY0a39ggxgS/AzUPi5DQUWpZTNeNffJitHTLueXwGHqfRtGKcVeLZuin46FP
wrztdG/g66nQvqPrMG0+Rnpn6ZKbCFhGHX8aNJYMyigS7OEG4uS5lQfArrQt
Jh7Lg2cxkOcFuy90JI27slb8bQUFuf9DAcd5WdX8tZTcZbge3cdS6L2YZCTI
OssLxkOe1/Ahlj/g2f+wTQoVIwy+9mQ3bkylphaoV1IJGo+y1SVTb6K7bqy3
+lsd3Vli7WLpAUvEF0wTv15fvnbj/cguCiQF7ooI+e+SLmbct6gNl1LrenSO
u0fYGkgY5IQOrDGja9jwIQbCbF27tkG1y4yprW4kMVNSOv73eGp9QAsZ8v1q
ta/n4AwOXDbgEIBKr5vwO8rcolCIY1fbh2CXq58hGQtwrjwwV3Di38ZPklVi
YbZlzOSh5IBu97HykFrimXwh9PdagQ2MBQjbT5N+6cUAWGYXRbfOzw0KovVD
2rIPtwibK2e1AjuaRKKMXAa/FcwK80QybzDTloMpTKRuy2TQ+hY21r8oQi+d
0a/gk2Ib350uoY++Fv3zkjSSSSIlZf/L6V1ULSdFh83ZprcZlzUr33XzXZUX
v1cVANRnDTH+5rzJsrFsC/JNum4IKR1d0CbAavG16UJjUcQtmIDzNVmfvuFr
N5Z0G1iCPYeLjhwKBsb743ABw+0REjqY8aTF+Idg2b1xLY0e1tv2Ptuoj6Uv
fjTzvhCfc1RS6egqrxYcMovFyzKm0QQQvRn7h8rFueyr7NePK7XSWcU2PToq
XlfEhWtwIDOcqsk9kliVpahCJrZv3i1NB+My7lsRTdxhQN7IAiyIZ3PnH4SS
QLOHiSGb/FKbJjc3TIh2irShp4idcEqg3QZ/fq5F1ZobNchHB7F7H/6JDby0
x4M+nLBv1yIa9jL7NtIwDYBpVlTYnpfylZcuMPIK6Entn6Vq4HAIMg7K+hqB
57ptNQna3ym416FgrpvFsQlW7J1r71fXR5o5W9o8eqtcjNZ5SI+5UKt3N6XH
uq5djNPvUtVKm6x5y0TwFbNARKkO411QAkgYEmpDuZgBDYhtVSmBgQ7FrnJZ
5zp2OLjz+PembbPCGt/PZi0IVxddIUF1h6GFyGGfLZM6Yc2M0ZKxtYmnyNZy
uqMMzIVUEj86eElIPhnCggxdSrHrlkszmw8h0QP6osa+wx6+DkoGIKcq+5lx
oa7RJTA3ICwdrapbsy98k8ccC55HD91YYdRW+B6xs7GvBq9Tr82sdOy9ubcU
6jMgBfTs7X4gl9bFzRuuO1dUS4jIDo1Dp9eeiWBY2e3KQO+K559mqHFxdlcN
cZHLvH1XFWt46NPvbv9TmplgEi8dU7HGy2KCCboT+lG7A/zLqZ6yfi8dRh8T
/OYxp3u1w0E6laKYxLzSSBbqSYfNYG0N4Dr1B4e7ghc5X4v3Wnd12YbsxrAC
1MV/ilrvgndZz1WGgpc77/EWAdgAq8fsJP3zgbVdwE3Oqx13cgLtDid2rpfJ
evwolYyIhGL7aJIgNgSDdcdDtu5Ctz9BbUw3YVr91P4cTIXKxPFzsRcHRjUL
+9SSLfuzSnYsyplMhN60mmnDacVlkpX696WCM+WuR/JRu1KnMJ6yiMDLfqqf
qmZ9MK4iDLSwnjKotKEUpC2VIwRbAbXszw7I4dUlMlIHJZ+bjqpyH30fVY7o
n5DT9xABCaI+F9XjrrUFDsAO05FLWTZMMRvcdetYL2tQok1Rh/3THck1WM1B
wieSgoWdj/5sQFS34YgmOpFFaph0G0zGnaccfMAsJZ4qI6G+Iuo79c5YxRKi
tO/eCiYvQx/cdqHgiECCzssHiu8zvq0w3+rCbVnWw2n2xfWyKBj0wnGwuxle
JWq7op/8SY0qKzgUM0EqQw1/cOjwGSH6b4SwviqtD0IjOcCymzJHe/JLaoFG
kmUAqO9h452TZALCcUGvpvm/490IUCFR1RUDcmdTElX7iWNBSkntPzRNtstW
XU/xSZgsfIAKqs7OgpfyGJv1w2T0bN/0dMOBSGKgsAumVXSUxFPbwz/kb4xc
NsG7QZDVN1goPPq5pjTUmC1YETJzJ5qx32UA8mfVM7Fr35uI6i4lFzh/nVOE
peGSiYJxtrb48/DX1ANVQCT0c/WMDmox/I02kzA/+iBXXtoKYoxBwWjdwl+I
vSdu+8Qfa1aRUOY2hkypjlgDze2Py955UqlTDNoI6pr5vJg+mEibLzmWNeMH
MqH8EuPVxIT9j6Z60DRRwb4vYtnZu6J/ya8h3o2jlFKE5PX17IS8lGDUhi7S
cPa283advKCMgIQPniUeApKJllfhhNfxOrXTZlzWqY3CiKRmrdweVsdW48on
bMo3DN588MhiE5ZmShApfLR80VkOlGK8xrQ9ZTOMvzxAnS1Bpy+JozE4157P
A4Ud3h1tFFN3ayE8zCXH2jYOFby/ZRHnV3YQ0bwxA5H9YvzVhk9LLt2IMN/S
Ru51IvMQDdMTC6sa4uILrfx1CFYcv7BAsTOmyO/phPGQvUmfzQxgZEtADxJF
TNiD6yxMLip70u6+I4so51seNXttNEqCuK6kVjQdBsmc7O/9dY5HMpgOixUj
A1KqeX5VQaxD+UFcQbQhniNmPfkdaTLqCS6w579eIHkC0gAWHXlNd02bNsCI
+g/QSU1rp/DBF+ZimHZ+riZjFYorb3OIMdVqA2pkuRkv0o1XzR0xn8cZJIs7
ZThSnBwMx6mvlgCczN+l1qkBom7Q4ssC0c3zv02buqHB2zEHMwZb7JcXimlU
0qkOPb8g1tCcZiQKJX7cnvFEoM/+/OYq4bsbMNq/9ODKtl2m/qYkWxbiaikp
ynHJvX17dHOLEo8ptLvWN4E0LclgWXY61H/fvbn/bMTuw2QCywPA23N6qEz+
DdmNF+suDBizmzIHEhnzTjFAR1g+WX3fRIu7W4s2wZGSV6Uo38181GllSCwM
BDAAfrHqkSbQRWIKUbad5AmaZlPvu6XppPzBeuD1c+JygHK0+AvMpXx6K5yz
ZxDUfCYB2ya8eM6YC0/YdVQhscZOkXvnP6hII+SBfJMPI6MhQ6yqauuw3xUC
2dMpvb6dFZI3GUlaYvGaTMJn8fU6CVRSpdr2Hot3iQn0LzVYOVZT+NgVonSJ
rR4ngoiGCTDhyucdaXd5P1Crf2Flg1L6jgrWe4P3jrZb9fVIxO7nhHocb6o4
z5jV+LgTfTmYvd4/s6BgAKt0PHCpX3woDyL/dz/TVZnfhqupo4CK6D069SlT
0LYjHE1AaUOcsbqc/nZNHXJHIqbmN1NDkoTvChmgPh8zHCCZx1K2h4WB/sLz
fX/L8TcKhyx3oVe1jE3PhV3ino0mnzBgX5U2BA7jTUGaKLNhVzji9ghqiu/A
Qqm+fYeDT9LciVxHv1q3ayBLXFZsQwsvRG/2g0qz/TKYMUJzEuyLfjWNr3t6
q3i80Ggma94JaN+KR7tooYdVXK0RBGoTZ3822xuyJ6OzDh8pAz9c4rf74Zbz
UXxJFGxoFuzmb7lPyiU1vmxjJxYR4mZEkWE/fKls51nDz5JH+dFf5fK0D7ZW
MQ/uG9ANE7U+L7zsLMXKYrXGBqkiBm7FWVxwHSOnyUfrNa0KS0sjB3lyWxeB
lmGXZ2W59LFspuKYwyv8r4+oQkekgN8QPxnmtDGjGRPSHHmpvnyM5eik80IP
qEd+AfNpx4GxfZIm1w01HoF9cKNGYhmJVJSFoGZ7DC2oDd+BtNXk/Wd9YYwI
OX5duUrXVSgjw0vOJUdAcYKPjrEHe67rWld4KSrBhNfJ34ZxgQHSv+/mYa0N
KbbM4hfwq87qwGmAiAN96POllsG4uLXtivpK5HN2hDJTswZNBkzy0bLGkRrp
bPG7EPd18IcQUQA1WJubn2NsY0Cgqkiei70FKqAZOtttF4XO7m7lV3iwZx8y
ucasfRqnVqhNoF3faAyQhz9+iQWokncZ8NOIOwU9oXlFesavgQGJZFI0Bkpx
SBpR0iRmFJ1BpW8dhI9mfZGIhpvxUSh5Bkut0lS2ZLfbbU4zsCGnqSnJ238+
lvRHY93P/GSO7ZFSq77JY2ftcYR7X1SocECmhkMuhWMXSGdRnASSwVs1sk8U
VDNPNDnvZoXHCt+Ue48PTePWxDf6dst1E/fnQ0PGvdL4taTn9gaKlEn/30ZY
pHc0iNSQ4vPqhPLH4fW0Bb6i1+5Gwm7RuhPBcz4Z78KfGBkjCGqDMpDlx7Mx
RCB1UJys+i+s/RcthixyST6Vyd+Ije7oya7MTRswYb+aVO3LZ/P9yL8Rh4C0
ZwU+qrSa/z2BxU8OqvUqbB2sQLiktul5lIclIt11k+HiCiiIxsrcNnG9bSWw
iarJ/XkjH5DqCc4h9rmvWLThvwSxSrl2yrxd7+HD8iqmbOp4Ov3C+moQKRew
SywKaG6bpM6aAQ93IoFt5p66hPoVkfkgE2pmYtESNb/f6ea9ZbXQrydi9kkO
eI4HKZNKWZYIvB6xbswl5zTn2oABt5jFPpBdRVjoLI2yVkSaeo3AzB4MS32K
T4oXaj6naIcb/bFjfYEwm+YuQEo/kUT4L+IndsH6Dv6hwOq84MCiM3sjdgi0
Otz4HMS5N+Fb2z5zuzgn6ysvJOYd1EmK2PVjgmorBXyESS6xy7G84IEyfv1C
LcqqwTLHIG2iQXbLTKxmnyI2heL6AXv/hCS/ijg5ZkW6fQfirsUvFadYwRDX
XO5fK0j+TwuCYqBcAmfFYCxyXvT93LRCxA7Jb417dSI46usJdUmeMmj2KnbR
xQDIHQk7LL/4/qt0eoSNbAUXIT9OkPv87a7QhR8KveOx3xymPC2STIypWuuI
mPb5u27JmvueDdAMhoUDrVhHmthMK+pq/GUJbjgrXkEzvJP+7JIoW8AYusVg
ZZ4rUJDmRX55c+cNCmWx/6+kwmAoLtzKAXczEUJ4O3d6Y5NX7bwqLuRz/x2N
LV5Ock+wWD9z9j8LHEKdODgzyceVpQbN063gpPdY/L/aM4kFutbMIcQDsBLx
3JLu339tAI2b3Nn86eKtN2bwLcWvlWOXmUtK5G+47TxPm0cqid/fuueOUWTe
THKyY+RDW1+/ToOjZUm2hbH3Xcxpl4r42RFasLj5QIQvSz791Zn/O1hvOBYH
vIblfPYnjg4b+gr134eXvZCek0cf7OzY4ArgnWBfF6hhXzxh2olf4/mDeZ/D
w0pi+St0P387U4VgoJic48oJibiCE+Zt1VsbGcbl/CG3NKWcm94+rKaG1BhE
l0HKY4KlqdQF5+zKuOue9ebsD05Jvz87WbI8bIAZMJlSRZD3ly82DZW/QOMN
UriwgeoKAt2FmFgwByV9siR2eO5Cs45RHeS2ATpYJVLEGp/M7e6DOjKZjHB+
DKeS8hbgRYnTIOz8P/7mFBkAy2XTza+/8Kmv3BnVUj/4tFjZBK1h6xP6979S
TivIxs4ZdAwr827R8AGNqXiYbQ58aeC0PZms/C9EMHdYs4w7qOC8ahcaBGho
y4IPQDq5D6WvESbY3suFtXlewmXA0Q4MM4SYJd/oB0+kV0sMONXtzG7lQ6vl
jUqGZemYNYGbjaJamcD6nmlyRXfeJdEWVzzeuct2r+1BIpJulrImvVb+JMQP
T5A0S5/42GvrWKZkNZK9hgtIKlltYZRkeM7gsEUN7hSmGdr95q54CCnGtQdt
Ghv3L1xFFK0qQN5fYQWEU/mc3CDpsPV0HcEcfOXlp5VrFApmWEDkZiOSBGZh
s/EsloANZmUX++M3+T8czW7O8cfYbCyiW/65jeuUkXamh+4i+Z04Pn5h/63s
JDo4RfVikb6tgWFECTR/9IMnH70URliOAO1j9RWDksvtkgywmPtUopgMeAe1
FH39cRRVcSuM6hrX90g+kQpReUSA8cIojL1f8IuQaE0kLFb5RnSjCeUH5Zfq
i6zT0SAS+FsooZldsaWzHAszOthOtK26dc018xXMtzhNUWwAUQc79jtKRRWy
fF8PiqpD+Urs7rlwSHX34q9+ncnHGI6KFmSBxmDbXOjwT5rMaEydaiat80Cw
nK/gHS8ro3M+NN7P/HTrFAPHibZmwrKokq2Igq6QAt82+Qw9/DOek7hFDaJT
RBFmExpFCP/4p60VunuFHW5QAnBbLowKXd6eLv0O3jj/XVNj2iquVkAcW5nQ
7frYrxhGKTvS/Nv1LNOYPcV+R5t+KaulaIRBryGHieMw+NI0bMpDoCWBBDT1
jj93r4beADvNjEXetXkVTLnOqa+GjyYVt90Kx9xf9YWNxnLscM3DLihrsG2d
VrM1220jCd1arsoBP2Z57ha1adsUwKBeXsrAzxH7GYx0I4wqYDvwRB1QFn8P
GAQwicWjTfvJZIf7gyu6+PjlJ1vReVL2yUSZ1qrpvk1qMiZkosC6GNgjDchU
IGgjKqF0OkMoE5tI6uDu5E2U9QjvsllRNIfbAb10qaGvjTkroVCEPXMdWD46
Tx+JqNO2FR5Z1UNMa8F033KLXV38zi93gdLdou5jBkkpiWmyhF5xsaWeYlWv
vTORzqZmqfbM1yFgRZgxnjHXkW+8BQAjr15TtQ15Ym5lYFJrzrGMiV48BW+K
bxzvqgD3wdqTrVSJW8Z5sgfIao4dGybLk13ACZ06sTJstvcO4m9VprgW89+V
x2MsrITJAb4BjsMuzCH6Jpp/knfmo5TVxYD5VSec0lYSFTBeo1RjM3kpRmwz
03nQWLeyFJwgcw76thq53DmxO8gbdcU2+5OLIIhgm32wavgxQ5wY3pvouGKr
C8iGAckqfNQjriE6QKu34szUR/ESlh5x4gt66brXV6npOv42WuDE1ckW3q2o
CEpR7C3190BlbX/uNslt58CyssVyInogURQo/TGUSeELhlCAIOl3JwONMc/g
ieNiOAg74IPe9u1u3+F8L0oHWvjmLhXcXb5BZ/KM09wnCt0jGpDNl1Zvs7XH
L6dSdqw9vxoCvzJ1SJ5Lvzcz1LQiW505PuF0Viiqlm1+a8FVSzepinxhP3KT
6ROlaMKCcwjbEwohl+AeL2zhUu/wfpT8iyV0uoXWIY622Db26MXGLYIhJALM
a3y7szLNoI6yYjE8R8nLFyTG9SSbNcq7c93Aqy5Gc2uHviXhUkP7uOFsRzmF
7gY8ZI0Sbr1h/OywmOBVZR3v6q7E4Rv9cwp3sYFMldpq/ZJA7RGaTG6n3Pio
YKydHclosgZcvRJhcG8ew/2Sw78GydeAvqgOAaIV3ax3XxL09eV/bFL/LE2Y
HKBmpwwQiqcOp8P9swMivdzbLmNsiXQZwfhWdRhN6oRNtPlHz0Sn8matoNgs
OfyFE1H7/D0dyBYIs7Y05QBhZnl5kPxted/UCh/ZZnOFekbAlzVJEsND5PP/
Cqg/e+iloEQpEzWSNYeODcg7WXCf2krEJbFjUMm8DHRYzofTiEqNTtE4XF3a
iMF68WJ8J0X7Kh0hbgcxLnztRNsEdA1fRENIeMB5ONhC2x3DBZCe+sy5RwHC
ZlMyTTmG1uzgG/h6lzm67wZo27ZOn291VckGCljmMx6Uw1O3v+F8VjTnsfJY
GR+D2d1CtgN9/c2GHMXE83/59kMs+C5MyMisTWwQnz0d7Sep4RJM2nLw/z2O
VLuq5R14ki1hxAl1dgWB9y6gqOAWMTw5vcUtOsAN9n9shw8wNL+EQAIBkEia
L5M1Nk+jb7gX79RBQ6twjmkgHJ2vFcILQ+2AvN/e4uAUUdYHjHJOtmfJNPrr
69SHiOSZNMmVo3rWA7B+ZoD2qd+3biOksK+sowpLg6XWV1S/dm9R58lO6keb
MRtTqv7ocVguQwGGY5vzA4jE7kZ2C/tvNCcp6uUyfoWccQpYnt0WmLECgY1U
nUI/gbMQ0aXpJqpHxA0vkp/lVElkOaxjXBtObms5smMYiH2mbRxw4quu1dj/
SmZN/9rE4QyMzLJsCxpwFHYlMyVwZhc/NtZxtBW0nVKFMU5un42pU29ENJWK
ujRjJvEJWDYXAlHCsKnwS7C5psATw6/J16/9d5u9YQF/nkMPkO+wig7q1ogG
5KPHCznpWMHUw/vr17ZNTSpoS/Pbd0xtJLn8J52Q9PGQKjv0mt2RySparGyI
suo7+64V/G7KX2PaKfP9ihf04JGqoS0zYjS+nuhAwUQeA4HWGHkTB9J+Et5a
0S3NezjU465XpI25W4JWNLsVqbcvd2b3jMDBS3j7QPYkcWPS3apVPOHpKpvB
+VQbD3ISoChQXEGM91i20dLgsSAGsu9aIBF2JpSS3GPIHoxiVYxZRjBMUo3t
ZiNNy211Xjoz/o9Lio05noyGXxA0aUcgrp4Bv0URCUvvBYJZYYsxs7K/VaBC
cp9/7LxUgfDpBtRrr+AKa1i2MJaPg0vSa8ORlt8/izhfOmk8HpCy+Ud8b6y2
AkRlp/Yfb+4GZ3+ulVx8jSxhPk7oZadt5bJao4gTnnTkXRs77yvasMhyJEyD
zMc90E+945UvJO9zp3gthpDqaAia3KZdRgTOfntcz37UtRk7Gzmv9vcFl3Z6
Nbc+l0/yK54dzDtzd24cyhDkvPbosQcIZ9fQ9BGELZEYlAlJKyrAFRvleFHw
xV+9JSvkijcXPGDnRge2OZkHNJKazc2FBCqkmdKOgpTaNoVC1ttcDSfv8z/5
2jHDjPRGtErNDKd1SYNknHJgI2gX2yxZEgOXOiFr3ohoAE3psPG+eIRXEsQA
0MFIEO4Vdy2jRN59hsPMw/yIUMXpVzIHsEM8TaP17L14i4KM+5mVNrX21VQK
Ob6Nm/Dgi0jho8nBMbgZGpHVFxzFyGdR1BkidtMkvy//0MOvwPH1s69ewlg6
2sJDzqyU81clyTx8+InRoJUiHWUL17G7UaBulPFaRfYUqESUb9BNUM41DnbO
ZKoslkCbKy+cP/yS1VMMPVQb3OJ9vFu9rBvaTSgX29EEMh0M0CeJC7WteUJO
youYZfhbduWzrYjD11UvCA97vDoon9sx/vZWXkBFqzDCU4DQoUGQRkfj8nIz
2PDP8vyYY7JuhK38kBm6vTjWAuMjn11lW+ORLKUHrDAEr/PKsvhe+maLyYMP
UzlMPeVSXdIpufNeuhGZLePnBMTSsYDHnqrCk7QpYRKXJEOqM+pGoTJr+PNg
9Jb5sYoAdApf8IMzg8QRfgWPm8olwO8BzHok2chKDYZGmgxmEE7ZRwrpHRnR
isYp8C54hOHx84xNdzZQJD5fwaeMugpXEXkc14y+5TwbqJ/ybaTIT5Tgiu7g
KeYSFB+9dmofIhtMRuG22c6EM1Pd72Jtttfrh4ZLwFUpJIuKiBZ4dNznGf5N
t6aE8ZmIhs2/deHg8f1kWnNmCSxc8t7oIyvuVYRrfDTiJ2Hf6ZH3LmIc875N
9gW+2k59Wfvk6XGbOsAWEOgMZgcRxm153U+6FAc6zztwLUk0bRikifpxl4G3
l/QeDGmCiBmW5han/5Pnnh540mkaB7g/P9DiP2V/jm9VBebgEq1dHVEvor+c
zuzCs/+B19pFaleljuGfYEsZQjP7GPQGU1GpxCVNDPtnUVvQd50xEbH/iT/X
dyOo5jrZxpxAb2DEK+lr34RGUbekWKIPQNLhqJA1zObIkYP8N5lgD17rff42
FFmOnSZfk5aYTTGuieP27kWkahVW0WDfrQSklcSrqKOO0+JWYbidX+epdUJc
FSW8bBW02wEeDCJCcTD8XZTxRzeGLrFl0egCIxlf1O1Jnrqej8LvHa+IGH9L
KSq65Hn/PokLp2hWFhcMTHhw+BPOXOo6742xvHKVzg96alRQPELuu5SvC/w0
Ttf2+0kddkYfCmqKbFKfAQMn5i2bBzVVX7Dmt6m1I+ksrcfto6yfgaBT6t1m
P1eUSi3V3SUma+gGxT3DR5LZc/e0+iQuPnJi7FciPG9T3TP7MbkET4aZHp95
jRBbwrKhX1+aRshsLlqbpHAlhcIvnZ61+Jan3W5a5yZQeHT3CAkh6VzJZfG7
mhiOyExgFOcmKMBWaWbTFX74vx5VQe2+LFKAl2YqKMH5W0P2F/im6Wsk6K1e
cJihQG/7MnQntNfDiOT0RUOxloXqggOcbZUV6hvnQZzDrr0VS24a0279Zqx2
+my9bCB8r35+K61Q4FjzSaxh8LAmtuHUGSYIxSrH3t2abdBbge89upwSkXEN
o4DcfkR72sj8Q/DxldfyVZo/p/pYCUMRxRsyNWM+WblrQkhGY1uOflIK6624
VM8sea8Kc3NBHZaLDKt16bk7ENFODNBfB4/ZPREdwIG2tN3OaxPVLgfDU4HI
vmONe96FWAyV/MNpFy3YAkVan77WUMXKEF+Zqr0HQ+zYxlBoAoeaXY+dIObu
6knXVSLNmBsAJnaKvEWpmn34MqXMWDaSDfgly1IB/RbEntxfX+SBGUyL1we9
SYLewJem+YWKujOyrOoNeFfCeRfC7I9avIEdIcezM7+uGwGq4LP5pyN6ZFo2
OQCMHCLlvzap/yQ3vUX7cIUY1Qv2o9fFlSx9Qmc0+LZpi0z3ctdsp2gXCFEy
7MwX1NBVEYNzi55fLo+gyNGgjoBpXAAzNtSEC6AniAS+p4fYoYvyDLZNCBWF
f7HUtoUt91WpLu7BOiZ0LMZekvY23jB7XtT0nqftgvIRXeuhlZKnRIjdCTAj
4BSK1T5CYqxbXRy8la/6js/QvJnSI7Qr2zZg52bM4XnfvmVyI3Vhi3H8q3+y
l5fitA6wpnntbUrxjVN6EZ7fX89X6gYEnItvAsDVOrAWiNVURgAqk56Wv+9Z
6FDfiVHz78eOhwzOLAnrk5wMwF/bQcSxttq+9qY1nW7CDVgfFmBAAq4ivQ5k
OX8lDn0WXehhdOpEkmspEe9pYGur/P8GbCKNCN8LV8JdeEoZkgn3yDrCb3z6
YbchOpRLqmsMl8YunE7S6kCWjhlP02uwZ5bobyocxdLvYc3+YD6MIo1KMpbm
LPoLnhbr9e7/A+mfQjqOyS1fl//89I+dfQFI4+9/A7B/8dfzJQTjOKjrLyQc
dGs01cB8L7i7YdMvoyT4RiRhHXX7jEv2P8Idc7uISbiyD39+QFd37vVbmVjV
E1e5YfZK9vxbWlcI7fb/RpXibht0OjEQ+GqUHcev3JtvV4jx3gxV+Ri7+T1P
jjkS/hpYfEyaYbiYMtizr0srFpyvPZpBRL3SJCS8sKGsJtstND7qZcMhQe0J
Q3iK/hNeUS63pEBtzL2zbQMk+mpZZ58Qici5SWH22NxLQCuuZC0lveGhBhgr
sbIAm5dsbZNBEtDkIb1SjM7GqMqTosdim+A0Kd3stBApu++HtO8otxqBVJQY
r3jSiAi6SJiXbC3cugE8kOcxkrK01DwLCVa7VbpmiCOfR0xkhr7Oqj85HkKn
aaaB3kT48X2UNQ7x3XWkgh2ia86+3oJWGskko5/aITMypj9kw21Tkwm9O5pp
LF6RHhe4N2aLCnF5sWCGQccG6WzMYJ4jXCs0vv7ovVWfeWhRGZRGUrJ/mMuj
R612FNAlLTc/dOpV4W+nBLcZeGQ+yMoOUgOGPWIxBvwZmHMmBkkmyEU9bkSQ
GzbFevw7KqC1IqWRtp75CHKlXUK//64LJHc8mTHt8q83Zl7FvLT2emXmq1jE
5qYrYW1Z+BcquCyATKK6X+z2ScgiR4BIlI0B9kzKBtIQslBFRTl6relnqEDy
fle9C4piwzYeoVX6xR6SKoffaxr0nzhXd/yjgxxh3SL91EVFhaRcOGXEC3tb
arC14sLvqAcvVFtBSKUMFQ8/BYjekJ/d+lH8/ghDf8c/cADSeiQt7yXSajLb
5FsN+m+YAjYP/E40cZKI3/Jzrkeg59t77TFYNsFyMGRUzCDOU7eiCJUX/DDx
QXmIbsqjdmcYoi2ZIya+txifrZ3OBvjoNaAF7Mkkk353Qr4D6ie32vJF0MyD
BhrEQIYqHIDE1LniUkZ+zAzVXhQSbvnYiFsLX1/uPLPe7IBFPP4/0X+HIBoD
et3LJ2pDniknPtQMQkjJGj2e6dK5SO4zwPGYBsyBGMRMhjl0lf0NqNEC/E6c
+8nU4i6rEqpiuhiqx3CmQ4M85knSx52cypz70p2N2Bd2alhIbbNEZTPOgtPb
PQ27IaG+SIqINllvvf3Q8izIW/7R2VTofqXGHc2wr6qa5NyxSNyJTQ5t+g3y
lc+fLup7yXymBf31E89g/10ytYqV1aFsakHXvByTg7Q6cjumpZCqCaTjj44t
mSAsWQWV+qlo5cqnGbIpfUAXYx/UTJNSkwUlL9i6ShqxvX8Gx2Yf/2DvCKzG
dVY4HHFLKBJkoD55W7xgbpZ40rhdeHzuUhjlegHoHxNfGfitPROHol7axOJ3
+u2NMvd2DgYG22OCph+QxxmOXEjb+8xsOrA+GHS2Yg19bGh33MWSUraCmbCL
Qm2RJAQNXU+BSEoGy4A3aYEbTWRrQVOAUz2SOxycYUCOxGZ3t+Chw1odYwcS
FvRCmP9J4Rs5AW8UfAAwozWfmLwsHA0UCSS50ZbeP2vVuIAQjb0FOdakjGB2
kWSDMQPBBr6l5iR5d1h1igNJcDiO1FDZ1E60hSuO6cIQ7TAcw4mtO3BVVjt8
xL+8eVuUVMzCmdQ7/7NMcain27Iqj7jPdJc6vdwJ3CrX9w9oSx2iN11QbOjZ
yxBcbFAyrq9/UW8OzZsA5lCDn+na8hSqlVvKkrIPz/8XAr2cpuY6CRxVSXhv
wjiSfeW4PBfD0+vRgYasDyy1TiCxNj89G7lWFfSLRZww0kHyLtICyYTwG4Pl
XhMYeqjW5VLLBMvqWs8sEEgrqG6YetzgamJe3EAKuhtCQwK1M4T4bucDcBSX
ghOwNPhX19Hm+eWAt1qYZyuiSmaRdjNeum5ZMMh08tr9zx/rcJs3uVwRMiUl
aUzLovZX9RZE9UxzoI8/IvGWN/H3npRZ5Ljp4pGXh0P1BhFB7BpMN8Tb/P7n
nICAK94M5htlSZyNk2CwNLLwY6TolE92dq4G8Wkh0Qf6eDDo+K2NgxRB6gMB
lke+765A9nBvhO0lVHzsJEVdtHcctGzqYSBiQ+Jpi2wzTIqMmRqCo/3lb66g
N50EmvOlMkD3Off20OdVzbmA0ICIkQ9BUL3hyjfQDqg5V5/83bHljxR/L8D9
SLr+bNyAR6IyTGeQU1myL6qiu32rqHQhPp0dglipa4CTWmzbRrIAW+VoC29Y
nGlI3zTodBkfLqLPgHzB5DF5hInL8cYBgXR6DL6zM6tvzfm3U68kRfJ2Kwxd
LRiSZd1UEnUwfqvm84thzUqgJjzF9XOeVuM1j1QC0RHY78haml0IoPBJq+Jz
vPZr8bqyzmdOjYEJ1NJA+ArrnBw//p9T5kEdJbZFlU8LSpxsQad3inek2ftg
7Eauqd2JscoksYHmrJ8yt452JrDjxWGaWOd3sQJcvJ1JX3zFpEPAuiW9X+WK
Mafzy3UlvEwYOLzK2hILbiDqaXXZ9qQjFQBxgdClawx844VPWzmVtVB/6oTY
Wty+xlmIPRBWnPO/tZ/rL5+Huxn5+9p9uH/H86j8jKAIejqDqYJ9CB9BgtER
SavjJSTnGuK8NY4ts948Ir20+7f2ofNa6EbKJ10sl+ZhDRHSJAgtEIMQWj6/
ADyzQcJIz2ya6Ohpuh5nfa5Y2Neii+aMhsM8jgHlgA9qkboxzqsgli7l+pxv
vBL/Qwp1G6qGLd5521B5N1V0oq6HdxsEZhvfJIVMANrtjUoASZvqVJY2323V
0dujKHjNMUIJHR2cFTuDQ6QFUAwqMSmhzrK/lLH65tcB6TONl6nVieZYIGlk
2bXY9T6964AdSFuJ2f2w2WZ+GvsnZhTRY0E7/UP4e3sJfg4breAnSN1I/LMT
onpKyzjBjye9e6aMJ7KRWTiQYhp/jo4j434OTGEau4h+VaPS8BThBPzrKZWC
oEId2uxiS1k/pttK5DRWFeeN0B+Kt+0NvAlIHSVTchNO1iwTSArOX6OAFMWR
9cZTjgaXPV1ZHb3l76mR2zFSNg65nOi8sEQbEY/7r1orQV78MBwnc/TbFt9R
MTMTQKtC5LlqeeDmWBy68kky18r3CQovRix4GT/++skv2WFJHEvhL75HmT/u
5v/M3hD7paMxEV189oVsXVzCDAYeOY8NtCAL3QB+0qBXhSp8RNK17h3DYUwR
rCS5EXL2uw5Frj2gjXMzyvqU7upG+dBJ4Lmzqhn4v8zUDHKN+fLUqxoSQ5BH
d+4e4NOFxFmGHWnqvEH77LAm1+ohb5cXOSLfAI6FoPKCuS5CagBR96e8lh9D
AOp6ZCGQmSblgR+1s0sQLL0fafU8BXC0N6cMUB8V/mqsVMWAMurj/Pn1npSS
OPynmfeieu+X57qp8OyxoARh/8LLNZfkDN6PvvK/CgwS9ISURfUi4wrXTQY2
yF+oIXoVXGkfEuKHN4hSc+cAcRMi4FW+Nr+/97FuUCSeq41BOzGrM2T/6i5Y
agBG/W23DOouuQXnMJqI+BWN4NjWMwoyFzkCW7Y2ssQU+sltBETz/gmABHJY
srDJIWBHNp9cVZuq/6M30qPzeOvyHgkQaY0UN55Ul0XIVM8hc0kwFpMVBHyz
hRY4GrrjcysKJADhxPsA8yEasL2SA9C4gQ9UJ8TpW4V4VmklsxKgY6pGHs+U
Yfd9+NM9HSJuKjvfvOJt37fX4wqDpoWq36QwOJqCQXEuYtYqpNFwe12ruLNT
G1eboBEUWvbXm9zCVIX7fjMarGFCv5LqiIvh0/Krr5V/Xujm6TetZQ2TSlnG
LpTCipOXrRTZsYYGCscd4O6/XnyDWxNFjcHEmKKmeCVK7ZylHLRBZa8pZhFV
lL4TiSE+i6kbPnTHYebbcDk0xQJUwNic9HlQWjY+eEGE2toylChjDfi38Fv5
uVSBugtdJSpTQwoaDGYCJWH8/NVKs098n1OzCm6kgRm7abH4zYUOmGFG4w7P
AGHdqvdfQJ1PPSKIeM969f0/mGLuS2KhzLBxm5unCvJGYA8tprT3g/Uo/G72
4jTIddTitCh2jhgTrd3NYTgjyqh084ocfO67FgNFSMbhfatVrHQF7OcOTaGI
XdAj5/3GkId83oob7l1IX46N5vNSLeu8/jrMCgC6wLoXH2L8aZFKtY4Ivogk
13APu4/ac5iaqT5rX7I8bEyHbCABBeshuNrrO4d5fHKURw+D2c/W7KGI74xQ
EAFwdEbpkguYoruf8Z2kwA303IKK0wEhInDqyOrIIl4BcT7wdACOmtCX5o2S
p7D8iC2Dv3I8JXKopD2YieljZYaBONe2QNz2qc+kz+gDr2j8jXo3KcTCrdsj
QMNN4004h6INO3NjvOAVkkwAN8YJmT2IgN7KnZ7TMHdBDu+emY1LBIQWENZW
/46A9OUh+WPphIFSnX+O340GOTwrycSbfuO0XD63VGvLomIE8kJOSDWtJPib
xl/8HOY7PA8+avvVpnyRdAm2KDd0fLZ2omcFm4sj+NTmKZ+LvrTFpbT0zhai
5Fsa+CTWSubHoiifnMx4fzApwCRKm3lOnbuqyNkHiqR/9AVvxutuZNuCunUA
EaVYT4Jf7dw+q0jjYQc2U9dIhXHU556UnDFjr2S6b4gf6USVlveVKFouUkd5
9yoiW1kvudXKnejJpuR93hXFQ1kkCU53jMZKxSCSjasjodZeogdc1+88AaES
Ma0cNnGzYCY02uLjm8nzJAAIE04aStjT086coRH2NmHD/RMJb6ZfZzmMaHwj
eUp1EK6F2hUq5i/DWX3gPKnZwiY28xYeh5SxiWWu78UNi9Ff43EbagQmWcno
pKlZA4x1yRXlixQvztuTUUagwKd4z37VN31T3lqsTdhINZrv+3NchqBF2N7B
DjVndl9y8js3gAn6NKfi8liMj0z2mDFi5rJvvZGw7T/EbQDr4EoUS7CTK9wY
ob+2rxxgTgr3s4FBsrZBJwfSzgdHzQFwWMPHM6Idqls8UEHd7ThYn4n7+RgF
W51i/cqDLJ1tvyN3ufescKlK83JlfifzBFYf+2Aav1Khs4xBGaSrs+IacUrH
MvqCrX+5zqHXZLKGxpRt1656248aN3nqd3ThE7fclBlKeZXZ6qSLK0egqn2C
kYQNWmFsgi7QDGujZkSON7EaxYuXXbGYxJ9jb/gWRqWUk5Lmb4zadHNXSZJr
Ts5bufYaLwe00XqwEHTDvQCvhI/dTT2Zfu+eQqSGOjA3KfUBodA1X4P9FtoJ
S9NBdhQWG4uxAbCzeyQE3zSfQtmYmnPEKF38n8U8wfEsYyj9ZX07f+r7aEmm
4D/fC7RRM/kNiyUzdze49MOLraEr4H7ujaZx1O/JfBfJjXFijvPCCbKbHEfW
dww8f4mN314PY+j0xb9WxkiZITwIAoCWHQmpJrJJEH9h2gQPo6wgUjMjvgCQ
cUBb1VF8eLU6+FCcPQCw0c0a2VyX58B0Y8tDUYK1eyJd9B+ww9SPjWtSycsF
0LPMm4AAD4xSc3IM2jM3UM8iT0SE/qQRL57IXBXD/Sy9ku5J6IDwpX3Xjw4T
ewzK48ZZ7+3hV3Myd3soIog++qBo8i3wDGvooVB+UiV2f7tHEmX7hoL9IwzB
+LlyRkENfn2aQrFQgkqDfDDPY1uQq1tzSkKLuUfCnaUJNL9NFkRiddqQ12/X
2YesipDLtzFg/gipv6sWGknG1+ewPSkrMeKE1BlepGoBihupOBGbNAa90US+
h2dY92j/z1NKJTKx2zc0qxcWlDPV+EasjLa+18hqjxLwCCMbTenS/X60NjVm
cjwuI5V03YqN9kK6nJqABEXyDa+JcxSJBSPi6o4bQ3vj91B5edHd3kaTfZvd
R5nW8vttPvLzUwcWS7Hl7bvYG7vqW0sGXRbDUuqw1LfuCpIKPq/FLcV4EggY
NI3/Qs0WsQY4p0FaYETTidUC9ls2/qhurQcNxgKQsMtzTzo6v/1U130sfhQN
IineyCGmSSQML8za4NZriAB0LPWeabpU81GtEFs3GdSDt1k+SuYQmCcNwYVe
oWDl8aezsoS2lpEDK0+fY6xiZARGDLeTFlgSZcsL3PuvzayZvgCxWhM1E5+0
t55f8pNk/QI2POorLzQc8fduaEW9sMAF0j7S1C4mD23agYrqUiPNgGFZqJH3
hf4j3my2tSXdpQJjeJKxKl9gPjyQc5D53KLoMovIZ9BjStY5ImNxs5txvdly
cJhz8bqlLloszm+EJf0WoyLE1UpJM27vPH2BaGNXIfp1hHkcN/qjQ0d8dlKY
fDuQ5IJXNOIgO/dbiB/P36XU7n+0rSKRpvWCQz9XjWDczLzFzc6ABsWYnyew
ZhUXQs028/exCUAIhkZF5MU8YAOew4/58ZDkT221yzQfIQN+5PQY4ptHVrek
kdyoaldOJZQurQT918fbCldkqv+BN+WLkJE0JvSgSOv3bWRmTleWgHv0V4AE
j3K0ewXgVZZ8G3wLZT3EgKXztcgkYXwUFXgGRLMSMjM1HmEizKSuf0AcMCrE
uPvuZGlBas5ILB+UJ2q5/5XFViLQrOPhQ/a3/YM3A7vYO6GvEbZPLMo7rNJY
aKY4uRoviZRD/ezBCaEcYTc9uWZqtMMMPOe3DmuPZg6Zp/vKMjB/CzceD+4g
Yq+qPH/Z7VFGjLqlUcjhwZGx8MgoQjtXdI9mSuahHbJJi+tbSgf4c/NeEkeP
ySQyYlJLfoCbjt6SS5gYO2Pt8d3kqXJ4HrM2Hj0+/DEWksXFtDjZRxvQbiZy
wTox4cQoGRVSKCz3LAcfZ0vGOUg+9mAkV+SkZcNKq38+ATCXYsn+AE7RvD8M
qAtlp1G3GOD0kJSGw+rVOdWk1j17Nsy5jZ5VVPNSgCxrKeM7JgiFYKV+k6cd
OQ5ashVMdn+p9WvghEa7L4KYvsH749fVXCEJv2fGfqbLyO40xVw8l6ula0eV
33uYctpYwKcL4tm1dpkg6/mCdbLc0d1k5K3g9BjTrhJ0nqQZsZS4Twn8j+C8
gRxOQ/cNg16YcdeG155vKbJrU7x+763rhuESLK3a3WPtmCMOFZ604/C/BmLv
l0ROPlVfqYSI9xaUXmRvNsHAQZb11XTOU5jcWqfwIjuJ28/9V4WJ4aeaeCyF
VbDPxGY3ghKmIcmgVJG2fbhMpiKZ3qgifC14peJs0FgTsiZIh1Zu/sY25NLG
0OatyhmIW+mfC79XwibBYzHZJ+DGrSSd7NNQ45o1W9AeU9STseIU4KAa5Dnv
BCngMNu00kw7PJLrD0wnKWkcCJR6lwsyv/0QRur/Iw4CYopH4fO57/4F9917
ja4lgWgl1j1R6X5a9ykLLHXcyQDkuTQr98SWeUznIFA5UEgRaNrCx5MbYBB+
FEqLOVGnQIaylFKIRQ3KFUeFW76rcoXyZx628HL359tjMYFRXOU0d+IodNY4
kF0my1W4cuuh/XikgCEPY3ASKKOvR+bPB/yM17QpjcFsHqFr6doKah1O+p3m
L+X62HtW9tHVM0qjhr9bbreO9iHMgP8dn287bq1IEpVkV/IwJUYeMhg1p+hd
vuRYe5UOnarA+O3NxTa45QiX4j+GITceIGj8IkO2L7Yo8MS+wN7ubxOFOm57
pQvaExH33yDF67TbXfalFF0/A8Q2j7FRco9n/XgRD9NeXBJn5IsATniPRD/C
IO369Sa12j6e57y64tXMOIwFmP+6JMI/RCerJu2k+PBEmidkoBCSnyd8vdRa
t9JkiblAsYfN/MPBbITv9Gwn5nd/1rFpyrBbI7hdrDBHKzYMQ7j7tQFKjJ+6
qqUPkFkgJEqmEHjQDRpUqErdNBVqF5HsG02FiwHHmMNCaizfI29+UAoZbtMX
pLH0fju3qRp3JC7CibYQ1Ps5DcmsOQ3WKWZRNzUR1AQOG7MeSarx4wYu1wna
S6U5r/PozqiWObISaungtkKZv2/jWI1cknI4movClo/2Uz3FskGG9fsu8OZe
Ai8rNxkeM1SsiyCWXpAhtOb30xrb0sva4xY+vfbPycZvzRORXzZ2LnLzO+ym
7x4VElez4Eyg3QrdwmF8c7ZglCNIByJUah4ewwmqMQiUHv1N53yVtQYN8Et3
n6meTe6LFFo6AiHe5xeG4A9Qq76U+DQJe0E3lINaiUxxMdin10CexrmQ5Ckk
ebPBMW5mtm7TSJev9I1Le8LPrKXYSunkY1tLqpa6egMyanBIzcbEHNwA7fgn
5pEqKJr3yfrjEP2+98GfUpkp595Y622zcCXWvjfGkfQs/v5uakQPxPDonZ0H
+VqKq2LgJwZF0h950iz9SLrefyj0VRRflRzzS0e+N90UJfo9p2eFoMlno/md
uQIsq2wE5mM4HTXWCn9LyRu6qiVfhczdgB7f3F45k0qeBTEc1LvcthhZeXph
0Qqjuha6R9HhcfNoV2EkLKNUGqim8FBEgilEg6KuIb+svjxM9sLGiQLtlRix
+9gN8xXrIr+rQclxElciDTtdO92LUm0GUoqX1OUXQs9brkU675SD/gcIEGmz
P3dTwXZK2wLRIA/Jd5QBW2rFz3bHkMFtgqICLIv1rJbpZ3LLcYk9aoDtq5y/
yhs4QKhG0zgY6yvV9R95gJvi6j8LIA/KoLBUKpsfLYF9SvMajkd3jXOlVL6g
+2LaIYFNyWUVZctG51LilCnmKlI5VSz3XlBQq9SQ7xDGCTkN63Tjf42aOujE
Q+0c23fJbFHK/VK5Y7wkfl5SzOXkI2dUudfB7SHiwsaa7FhMLtZTcu1GrK1J
9ZRysPbmvAVqCmlbwF3iwvMnsHV7MnL4IU8NRA/6A/9rljqOg5Nmx+Jrns4j
b0cpgYOGtI2HqYpvP90IEXqzd0HKVJEe5HV5bi9rAsk0hoGqsYhvnQb5IwLu
SE1NIuj/2V3NVs5CSj08D3POjPS+OYHVgNRP/HjxRoKRXnN6EHDSTjcaIH46
7qNe1CRDFpbC7lxIYl6x8qq9kC3G9I7dBp3iIZIpZqBaL/ECmlexm6prgD2L
7zOJF3zmRRurYquHWt6bKGEng4LrvMvsk3dnVSkged1C7w5ZvaMbFUKxD7jv
3g0qpt7yR8a1b+RFFSazIJ+bq0su6f8xiXK+dwIkFlQ7ryjpWzF04wwJZWi1
DFPbLL8RNBFV8iuUFSZoeSQXxuoY/bm9t4yrk0yZThNQDwYSxwayVBiN6Zhi
PPfhFk3+Gv9ZmE7BkusdurPoQSlYPuOm4IX+pBPkhwKnpgKsj9FNo1pMJXIB
KjbGw3j7wgkhWqvGe04ftKJwUwaJs3YD6o6cdjSRmkJO75flpY5Zn4JiBq4n
vPmVm2q8oOHL/MdVTq2t6wAkRxqaV+60oDD6AnMYJeWLjQvUHwbf6RUBjqDC
qwigpbnZWQ/Tx7grLQzmGPEulozcwngGIU/P23a9/hvyeBKp/o4f7C/b7mR+
6WNE0hzXTKHKGXyrpDcT4M3VZWglP4kQWqnh0qm+XwQ7qdt0PyclKCbmC1V7
mG5zro2yLT/MwS0ye/sUh5Y4pU8Y/NZQg8hOiNRsA8gt92VZm/gYeTm2WfSd
5kHj+woYLcNZZIXIhvngQLtV0YvYNpw9rOTRHkOXRPFdBVoo5ykfviqjwaHG
L8ZQUsJmnP9qO1NYobxvkLnEf2FL0WxNUdGJ8Nip52YleAmxcCUUAewPUbNV
+wovgAz+GAbABYi0Zsv1uviadoMmOhxmH1gom2V1kJlUPDNGjwJkpRypf/Lo
a8LNoJCx26Jvdx1INwZjVjUsEEQrcMcYIrSUqw/wPaJa+hBTAPNCxwRzX/R6
1+P2/uB8zSnlcT0RFT+2gugtRbQ5DZ15wJyJgHR2Wd0yx0PAafn0FG7FUFfW
1qPJ65avfdKkRBaKFC4G1gso1kCF4F7iLKyq/9vNue3hPo4vZ5ZnUAcrhcs0
DoRh1LKRrKoxbQmDxrHgNOTgDcCSM2N8WV8Uep0iwaWXU1QPTVx//gmZz9Bq
EAEPtrcSzIN+76ar7BLMuRcOUFIqomodaBel6f6hbKLeDrP6tIQdEt92iNXk
YZ5Ricn9kI0+1vTvHpUnJP0/gyhw1bvLMQqFVJeFNF7/k0ruwQjSEzTOyjct
dHVnEhkjYRItUMbezH2MV8N2PojMPn9eunPZPvsc/lnijuFACWIElOgKozTs
kdhaQDANUSHA6VioFkoYziIfYgy3YmZUcgpoSMfob+hrjUaTlv6G+Ujd/2j9
nP/9i0y773gbSZwhUrOsbRitgvd6eWKxxFq/eCknq4IW4QYG3tZkH98rR4S4
0Ald+hbArpztCNYZm8U4oUhsx/0EaVXQLoYIrwwMdAU2JGStEKZUHKSRN8cU
ZKi+LyGdYc1ediIMH5BJ7H6SIvItwD/yRp5/Adq7fUK2vr0YpNWSRZ8WGe1G
salJd0BDJx0TMLfBxDhKYXYfLN/9JZA9qSPohIrzP//GnTS6fpWUqGn6SkV3
TFEPxwQawVY8TMwu+qUpPKhchyN/gI0ZHaoA8kB1PvmEAIvCKl2NGzH5x92+
NOyp77FcW1fyu7T1a6r0urL3My8XW8slM+l0KRHXmZCBR54BVTYBFT9Dmq6z
213va8cs7Ed2McVt2Mpij5GuL2mm0EMrIq1oHhIcNoBV1vM5Dq08lzOATqj6
BfbQfsnvhtWVfM/Bfi9vUEtdGW4E8RrXrdd7Ms+UZjwxSwAVxJUMnXzMRlPs
YXEmTrqAMmPHr7PnDyB8JXQRFWlJds05jm6l/idx1urxxX1eqUZeOUrED8KY
PaLtf8q95mnmCX8Yeutfg3t+u3P4VB2yXALyMQHvb2zyBiPUkCQ4wVvXrMlJ
RorP9qh5mYjhaPGhNdDykM17izasn8v0X7YJy71HiJaiFD+D1BCWjBBsa8U/
2n6cRLuH/W0uHHkTK28uPBJP1PtNfih2YxNbyANQQ34wysrGa1VKM7Xtf7F7
Zy1ZxVuhMQ5czIzHUGMEVd1GS4jq7ELiyfX4iMc4gktz6alwNkKUW1dQJQHY
Ym0lB/ksU9SjL+Se7Qfnz7MV8lbSmIQkNH2ev/JP5OvicB5iGovjWBtepEwp
cBx1Y+ooC5R+QJJRzA/4bK7OiiyScbvO29tnCJdQcTZuh5NMU+om+iszgQ4i
ePGK2Xy5KWhIQZnAzcjpULGbsVGcAUurhUKtMR3wPisOCL3pt+K3a3kerieX
R7PCMLjw6K49UkMG8xl5BrmVybeuYXxBa1gxBwP1aYBHtrjRvRsrOlT6chLx
doG1yTwMihghoQIkjGrjXgcHID8aR+/Cp2vZTXgGa4yLXa9DFjATSewPxq3+
dJ+A0LRQDGs5CWoSlrXmsSy0Tg1yPqJJ6n4Fxq0m5zIjyH1FdwURpArydyX9
/7oOIjq1elV+yUdcVMCrdzxECpjMfPTnt48OUkVefWjzynX1YM1Qnc5p8+bD
2tPmaUPyvf4W4vih+7GZaSZS/IR1mDQclf6EptsdqC3tK3QdmFyT99yVt0IM
dvpQ7jwxzS1TwMinvvPWRRtdKmIrQNpxJL+ivGHSlWo1TP5mVGzX0p48RpTP
6K1wORHoUU/m3QRn7QXjbffX4+CC01KVpOJ9oBr6FBtS5tCkkDwEiKKo3F+a
zXLSthj1pO+M6UaaoF6YizLZI/zJ5wV3b+iQJxyyrXc7dJRc2x8TbSXJBOIH
mISzZFcWyWGI2gxQvjD0WL9vyDJSHUFWxg6ho8DppkJnN76FbnqyBRfGxG0l
IdCrWST+r3O/mEKdCo+5ps0dsWJrAPZmU5p6nfz6NRJdZLVci++xLyRx9EL0
mvmNNc2r9Ft7J6zqm7DCXUjNiC0op+JIo4PKU2HqkXwGKcIY7EX+OLTfzON/
X+C73hKnPzCJCOgUO/9EKwMoyq+SCU+Cs1H9tOkG/o/zfitcwPc1nzaKm7kf
97xMMPg2MxWCfjpvvSnoeqBjKzWrW3D+bDKZhFKcrZQMZLwtDrvAUja6Dqmk
9/vHUqp+HmTA9AM+Dz/OoEX/b3/E1E3TFW+GpzXVVmFvorBOUP+E7TrZeTbE
HODegN+kHPL/iCgylTg4pAcr5i12CtDYRvvOQkenqVQFnLgXNGrlt/wVUq+g
Y22b6v84/uGFsmxHwgsE0ezDLskH3nLBfXta8OloSyUju9DtQRlySfYu8+WN
nl/nGXR+Jr1y2XybuU+hUOj0xexuYoE7Kff5nevjQvzw985KDMrIj73iXfLJ
F1LP/HfOqXU96WPyDFnlzc9cv0cvK+TH6SqI6cQkxzl559FAk36l7wtuq2jJ
XYbLFyRFr3K47Q2uAYNYU70BK2pjTyHVSPjQn/wZ/1nTFOgYfEJykbhBKH6+
V0fhKZ9pZIVJn4+NhEO6By8XNP6yvSftqtKHbE+SHUHcII2UeTMvKwkbyPXf
tKHZHI/gPWLtb3oIWjnfiJZN4ONZVXl4RIZZw8idUBs+hmQLEGxGAsX/wBPP
kIStTlkzs+J8ws8DvOxsluQZGyw3+/kRPNlLV2YhhDC7pnw0VnUa/QqVE1Qu
an5v8G9/wDuqSecBEjy01G1JAf06cgVy+vWOTvt+FlEpu3NyevBeg0IhF/TM
hTnZJ0GcN9WKOMP2joS1STLSVUqhkWQacmJz2vJEU3I8nSEBAfgP7/+TY3km
H6UjZyaCYaHmFSvAW7i7f6EJFQaMDJ8MAnVasLt7YSsMm3KhUA2PDJ2Ne9CJ
PqPYMfqlbKnWyUt9PdxMl83TQLONgiZziO5c8pQCTkN8pKGERS0hTSo3bjIJ
3lGf+8S1zdd4FT1MkefOu2MNnXTu1v5+OnV2QF9x+IW9+4KdN2FP34MQMG6M
4XjIIRXKpTJZnD5B/ecTYNqppFvxL2IxTiykBRXB2o4X3DCotSEqc1BAyAod
xMANBgQj31HNl3W3K1PB121zF/F3anT0uJ1GcXzA1GPQmaulFTSLmBn+UZVZ
dQCo6nomwBIg6T0glh2JrDxeLMuNd7HD7ggMgQ9IZulo4YM7venPUDC6P2Dr
IoSOzblS30b2ZXljrYPLtJVza5OyFuvyxffhfqwnQMBBcNxlnSe0z2cpLgJh
CMP1Wb2nLFaewnWDTi9aVTRNBrcYvSDIxrQw8gVQXBPcw+nYOgN7vHe4IvFv
LfhytKuFlLGs+WyluihPF0NCvU4ZaiI86CeRYl6+x0sr/CXRlb0pdDDdtEcM
O//8PF9VbnOLHI1MyXspFguG46bAdBIba1D5WLCAOLWSWMkQSZvGpO1Q7F13
e/jbV7qFNzZPnBXfkZAwQLHyy3o9B/8qZxBGNCz1/K2Tb4yvn1vpnPmLKHkw
G/OnVq7j3yUQr6ywwDC49q+O8xOJ8S3vJ4si93W4Gs6xXKiWyVTcvOwWk5fM
8j+BSn85qTKXZHX27fVpDOu2S6CGHE6ANxqeR6Dxr/mAbtx6yEXE5QDXh8cI
iSg9bFQBCYYXcErKQYpPhb+RYbL0V6vvwV5PiqW2ahjWcSBzWIATj960s4iP
/DmdNagap93ltSABwgQjieMo2VXCCXgBOjzhaiNDSvzfllc/2OGWhUmzWad1
U4gP6svAYmRy59tr17eBQkq8srdboATnN3D0cyb/MrBKKmtyV3cATRFTm8AB
hYO2HegA1AR2B4q0/Ok4ZT0iAu3H+OMsca7cR6rdbFTTDSPiFplg3U5+YPUl
oEjjsCHvfOS25zfl2CtXP6vaFPFu9YWHaT4JWeuoCoOd6zJe1Ib4mmpqZnk5
7nrQhu+EXkAq1UJlszVGBevfQRVryxIsATnWFCe3XwEDzYQVtZN9GVomcn/Q
pjTC41btLXl2JCj2yBX1txnlAi0PcEOZax3lxM3am7K34J/+rmsZCPm2UBbY
GzKqRbjeF1bdsg3hVU+IoqmbDE1hQDJmNK6TG6108qmgHke6aClZQZAL1K4C
T9NtqLX0IOrdXzMYkRzd75dqxigGch3gw6P8JCm+mrYS8ae4w8A3w7Iqh8Fw
jhq5dN0Dm8ebcS+wjPnaJAjOs4NqTXBBRzzf9S0yiBVFDKZO84X6v0ZLMgKQ
9OgKPVL92TA9QsGF/hnWFZsW4yolzBcf9pTv/Ydg5tHWgOzg1pQd3VBdaAv6
rWNqrfz+h1t3Jcn0IFWneT27c6T6E/ybdy8qdg0BldE+iEA9YLRrDVYcLMLU
J5LIXwa31bOoOYqtqO37nl92ofx8SfUTawVUuB4prefRflP6z9eFs0/jik9p
3M8xbN3RkOVwIp/8A9aYWD3HoSgiymrySm9Ceg27pqSQD0p204Axd5j6QrrY
C4HHR50LmY9iLwR3h0KOUirHODb0toP5NZiAyCQrI1VrNX4kRFFAiezhyxsf
PCI+rBZKnZDGlACdoofdw95b9MjUszVcomfCNolvehTyXsPF9yRyeA2dNdgj
Gxx9uz5lt024jWQgQvui/lnet0IckreqV2V3SSqRmvyjuthw1h/G2OLgBYGS
Mgx7J4muXIFVQPIUZ2O1WvG/qmCgz+kfivG2iguzybLJsKf4HOt43oAABW1v
Io1bKMTmsWBgD/kEy/WSrsN3rpl4CfCTgCtUksKmPk6M7fg/L0ryL84BQCuH
3MGgY+Cp5yEvAtLcM+H30FP68uYsZCG+Gil8FvWJ4MvZ9xUce9zj2Mi2chsQ
qJd2cJI71bRejpYHXTzCWUDNL/EQ0Ud7Vzb3BZBk+4JdMNbWEe4zKycJ4EgN
FwwALKMfdEjsShuksAnqQx6t/sPeTdaOoa6FldArcRozsYp3C3dkoau38q5L
UU3/Gw5+467CeBKovBdKPiKF2b4+pabzoQHwDXcJlPy8/yJOoT+kKGyX68f/
ooms4tqZqjBg1i/mbPipJJyq5EjauM9AJFdQwul9OvF5kW6MawpRHHlUOC4d
1kgPrRYPhd3/U7l0kFxoKkoamo3u3lxtphZpRi25TCa3ylizJxaKH7zBIdDx
30tFPyddB1eSQ+NplAgQp0UFKYQaHrttwSSI5FH2SNRywwyy5EUNIUVkslTo
vO9/GRKrT+z7kQEVkTbtcSNBDkJFBleRuF077p2XTd/wBIKFuXmeRWuiFcTv
0O3Yuho0t3ObdZ6szlVbW3Vt8ugbdCPI8pfYxarpeeROODvAn3H4Tgf53XpL
spEsg3dRG+COQ++birRskcFqkXWxzee+zNfbpuRe+R+RtUH+hT5WGEsYx0M8
8FIil5KWrscZfGf5DdHfxBKni4VWl6lp9QCFKz+XcB+lJiEJ6oWua7GM0qs1
0qAh0rV6ghsxkPqY7gP5tRyU2OZRLMrEG8GT8vm+0V/Ops+XPWeSfC/57O3I
6JnjisYitk0nTA+tTAT+VnqY9BoqCF5385FaEW8z/rfX60h2dYowwrlp3Ro2
3XXb/8h5lBLjMtShUzEzRyUX/JTAcMnLXZ2kJlpir+gGvkhGAZjxBUAejI+b
FGp6RnHAgwf7PaiHOUNMZQtVCHjc/PVDG37cvpaXUEIwhGwBYzsDA+vNsFA5
PdN2A0DcsapJHYuXKrgk2wg3ZpORrlESC/innBljUH0vQ3LFKD8hvBPzGimG
pTYJU45UxVzL0zsh5KxkYgZTcdmTAsIJ5PNpeflMzxFUl+1ppWw4q2TS2EZJ
fRA63FjBpxljuu7ifoOqF9440Cz/orasmFcf0rVmGp++b/b7VeK6MUfRM+aG
Naded8zF4zsnfLCXn0msAu8tjj54uGZn/RVNTsJtFGr4emFU1Jotj6cjpOrJ
Ms0F06uQd6oNauqeqWoPtPEy89mpyWtkz3t9nXq+NkA+y/buTF/UqY13ZEyf
MCkFfe7FoQ4H+oasIBsXIl5jGfUqCRVP0lE3Urjjtu9bw+oa/lcQr+tWg1xV
LN/jelndKiIXI3hMDeCG2oTDQ1IcKiGNg1q5m7cAQZclMARGwVX/ScZsLJlf
gQRUfjBveqilLIu99jeOChTE8mT9p0KLWsLueV/v9ND0w6Z+6qtleG0Nckvo
IFbGu/mF6XB+s5i7jEEPj+Da8ADZblOvYLoBlg4T+r0wobvyL4evAERXsUUv
gwD3+k7G5BUsow6AYfROLLIplyuYDtKW4w/aQuG4nVQ6hatSfac4bjnyUU2z
5foKaQx224tnLY1rkudTytbM5aHfOeB0ynJEHHGkonGT2ZwIqfOCUOaEJU/o
x/ha3nVQ9Mch4LpRorxyEZj6hpxAHhhs+BeYye/KB705VpZqtZzAxOXnYMsA
jp1c2kqhXtFdSl1NUjKUdISBi58I2XqDuFh6/yI9Eo49lyvSYH9b6GN3yog5
ewmDaPv1hyYoYFao+7letakbNGxvdvd4AKWtr8dkVMAzEZUc7yZ7oI7zxa7/
YYyObC26/FkUiCcKrHaswznLd7F4S8xPZofvzTsroQgQSws322+GpSAo3sIf
P0RFX17GdFQkE5Y9fsfi41Q3qWqWa8NnxhWjG4eQ+iCQHAY+Yae7Iexjcgkg
Fa0GByA66Qtlv/AUFFS3QZwwNorHotaaTt9g8wVRE9S+FyeXMWBLarwsaM91
g1idLjaUHaggfz6in8OppvpjS/GaOjoNYSGS6F/xaQU4+TM3hiVX0XyoIvca
+HPuEdYYvWvJXhY2OXaP4raIkELc4zmihbS+Ebak5WI1reNKovfK8Kq701P+
Ab2kKIhl+f98DSCbIvj0xWQN4w38I0noJgPrMzerwlDKr6LMWMaYaHwLzTQR
kaOWAINwj8qpjA12lLQl9S1wIlqTVpdw6Wvb5ZBIuCgAyC8AuuNBJmaiYouw
QC7iZDd9cmRnfBPEcwd2ekR8wdmoGTgXQ+w0SCeAcXUo5hbzixjUzPUBrgtO
p8BLmWCsOUve7eHc4EZqiAvbQULDcORmg1ixUZM/WUy+Illgei18hOrS+8Cw
ZoADeNoWr5UfGOqbSSExLQ85wJWoGadzJX9LpwLtRmx6nXGK5tT1nI6S1viJ
S4c73JW7Zz/2kwaMM+l6Jcz2Okc6vGQ7Fi6lqv+DagCf3gpjCvJhTe9SbfKA
Ed+R18sA1eRC6oVa4IoIUHDJ0nrxMyg2xW8xmDD1PIulwEbQ7BgWbBo4r2Ij
mWXZ0Y1C1pNKxwuwXQJhH5ZFpBZ8iCW5HyZS1sQRpVYxhw8Ws+LeMTBjtbQV
WcO9wuff7MnCQ63rdH2IMo/vtiP69aoU6wPRgRhcZArG4rQLfepvuA1WYK7O
zoSPUxOqmooaYIIfXdKoBGowzI6OVtie6rJyYiYGfZ5sKEmlTSs/E4ifoJUd
2PUFGrIGOQ/6U7rrz4g8DB9FICCnOyfDj1Ga6/5lS1UxH5RyX4I3qRXsvduz
iutIiROpvvkrNknwDG9jPYrq2SCLrUvaFCpQGXxWLHZXpv4NiD7l19AYZg2j
ck16wMT+VesWLl+UnRpyJ6Sw6mhLAI62p2HHh78DC5o0XBEUDWdZrvanI2Cs
De6EPCaM4nyzJwqpvCtLXKg3QVTD1QEBCy5JKzRqOhHViACNGQ2QXfLu+MGz
26oa/H1uqyHXMOxeqkuJWmaamZe7LoVnZshPtEdMUiB7trmkQp/R6hlu0Icd
tvEvWVEbyP3ho497ryxU/tFnxAvaWZyf1ePVdoi4Xuk76/sySNazCix3HbXd
ctHpWDqjLnzgp+xqKppNMtmuqzYB3hKWvCUdStpx/kXfhwm/dFxqp2mFq2S2
iJHotGoqkL6WhOM7Ad6vrGH6B/ksmwYeFPJlZeCvmDptOMFuFiCnKOKyq2GB
SnBTv+OUTAddBzmLHh+qqjXiZnmN43op/QEQwwUuVgI5/V2qt4JqRq2lj+0f
lLec5ksjdKeVRlK1Oz0PXYXnpUXYYGIs0ufdJLxXUtpwAZduFLCwChfHRQBZ
eIU2q0N3FKcvILpkJFixWIsO9fjDT0blEYagtIo4Y1fqHhisCsAKLBcfyB6p
Oqd7PQz1p553DpoTdiTNERLS7EelDIeLY0AmV9reUDqd7EPWW6QuDJpgus3Q
/Df5nwA8Vu9aB96KUFrhNlUszrVrgMlG9ZeNF5Jk/DeHBN/ADoVfxJyi4ds/
FedGpH+csge2ogGyh7Fe/n2bEgY9SCvZRiF3ul+414OIi02oYV54tJVUN/Zy
8xV9r1VsNZ+YZjszYPHGZMjJCW323zVdvrTuAv/RuXA5/jNPz/EbrPiJuUVh
v1l2aXKMAdnmNWMnIn/K2XTNB2u0lq2ynPHRWaLe0mM82ibHEVErVDZyJBvB
77QSvHQ6aODnBz6sTziR4kstiD9q5EtTWpQGO6oRnZE/fENBynTQweUrzgm2
WdlxHLa9LwFdRycroVwFxOi0UKJHTCBsnsLzItlD0zbjSiFwkWgD0LLV84B3
A6zKUu61uzmJrM/xOqxlodPFjXzvGUUoOiTOnAWLu+o8tFZeNTMWpQyUXOGw
+vTTZ9MAbnzIGZVxsdvGba4/jeLvLzw9NbQff3uKF9Rk8kV+OAnXSBAZVV30
ze+VKRmSLOjAHkvGFNmvfMcDaGOfnqdbtzGJ3xpE/8j6BbiBprzF53iY07Fz
VjkmeRbeOpiGmza8ls0gI224efSjPA57UVg7beVRkRCr6p5ZVPukYZ0gJgCb
zG35+W0/vie0S3GzJzbk3vBUvcSE2Lws9yrab1BGinfOwZ74A+3j4VtszswZ
2ThAO75v3TEdSGldyCFy8GjNizsCFCGaZkIj+9GfQssT1KU2aJWZwVNSTxh7
kbRbqnW3GemTXnA4b508+OH3rAESF/fZMTHHyMlO2jOA65RnoSzj+R7c/QTc
lzF3FuFx5sdPNTdBVKmMLKD5u57SwUuw9UiFN13PHVeggk3C3t/yXZdv1Us5
IwlOBolPlJM9CK0FpDncm1wUVMLYB0RE5nPpr2Ln26pyTWhSNvz6fM1bBL1K
zD9SatuYby42yRAdhOm2UWA1rHt1TnzJpYM0kMXznr/eD9y49p1NxcXl9I7q
cBczXLKQ0F3gj6wWm5YsA6QHG3YO40ooj0aSkLxKCmMltAw1IfNAba3E1l0/
C3dYlEHqybZ1+ZCU/VT+MqF3HqgpSVaeuBF013mQEBnM/xbN3Xwv6cWvra9A
Q40fCQkB6clUCeKlKPAItjVmJHrDOEznCrVK3uBPzDWFJwnYqUvl591OEani
LX8SlZ2fZNVvL/7OmLBs1pC8kiQhdMnKq6XX0I5aJ7tX+LLAVVqLZCBYujIZ
3ct/r0rtQPlOpxnijyTl966YCdscx6Sk4wu+Livk/l2Jkw6tcZWCtithTO6g
QE92TnRRUliu6w3Ik24QGRlo7c/pVdRyAWIX/DLJdP5/Tl8d+dHe6uE7lubG
TidAYBin5cQVQxdiFVU9zf66xpPeeR3HtDSOfbvi2onm22mAt0lgJh+ut2i1
ItO8Rf89z6V/Q+9QjZVV0niyO9sg8kLH40VzKamSPOdaoouyHBpQpKJ6ApRP
YHxx6pFnTgyQ+SwWcFan8YJIQSpcAiQMmMD4kcYlQ+24XXQbQtO44oSEmc0O
HOeokWarKSuBJmtoK4krxGEwTT16B1Iw+Lz9iAsPRZrDquj3dhwP3e/5T29w
/lLalsD94qf5Gr4iPtxA82jIBaoTT6DMHmBs42IR6gLOAagxbZ9lQTgGWVIH
FwX4FQu0+yUG0tDeulE/z8ntsFsIRI/X9WZheUyc4+B0rp52p5yIK/TGDqX0
TVAjFQCvoEIF52P9M8rFyRJ0N1EcmI/aoBEMG9r9sr8UIPINw6Qyn/Bx33kj
xIShsomrobN8f4zXG7+PmtkM+K5evyj1bbmMIsByK8t+37CHGHuEsFi9esXH
rsI3SW2cYeock3YbsrqKDau039CkGnboq3U6iqjGSLYlYHZT6q07w7CvTRnH
XxcJ/BNX7hAjxdvWo7OjIdIJ2bf0dXO+PUGHKHnS4nO1bEzaBZszQ1nfGbZj
oDVr0kMopgJVNf7RUDSw6HNpS+NSRBZcUluPYnxrIfJVgg6KOBUyGMIW925O
SRbfPvx1lM02ntwkx7tQCyhLlSvWQP0t6GqM5Vw3FG71PQqO8UA0z0xOJ6Tv
fgt0bXTbr42fTSSBuxd7Z05JeMLsbbbFWhZYConeAMDGh9RYRDM/tagR2/Yx
zXuy9zWUNImxuULG05rXBcqMw8S7eTpZMVjjYQa5NJNgOfy1OOS+CIqu1l4+
a6p6cCuSnZ2mSZc+M6qHvUo9byMmli5YK0RYHBBL3S/VuucH2NKAUMtGWxOW
r78yjG+MtXqdzFDBgy3oS5PbqjqgyATc+sxpQtNxDs2OYRHweTx/xTl0YTTC
rMvC0eOiVV07HwaEBTXuTYEFkslgyar+TM3nxx2cJwpSXf2STqWrEAOL9KLG
h2UqQb25CR0Z13bUIFSAgp3SNi34CVkEPsGG0OeDr8H+voh4CbQjaXdnbWMP
y06+U1Z32n1d/eH1tHMstvp9+wvZ1LPzMOZbXTsrXCjttUvag8In5z5VFeje
bul3NaYY3drCP/5/zeDU0DPiaK4zWAFdShLo0ftkWQbiRMh2WG+huN+5InwP
M82KESBgG16H7GT/gOPXm8yXYgq5qZbWvyVPM+L1cwBmmHW2GeSPAC5vr/Hf
ZHsBxnzrP6aztFdvIQ+orazxN/v71baOpu5OjCpAo8VLTOmP3zbd3KkTEAf8
BDh5s9uWZnqRVW4N66kecqtwSigmor2ac0LUhXYX9Q3mvdRrRHexUODQlvKW
Xec0ItaXsx8UiZSDC1TNYfs13OLZBj6gmMpvJOZJDrupKyIRqxKFwJjGLwpM
T6lU3LiWywSl6YrVJykhQQQGsUGcB17CERNHpRBQT3j0wDjmx3KsEpGEWv4j
V+90AWV+teeJzO4Vl/+spoMoO2iOxa7iXcmznP3jLKeFw/Bi0DM2nJ4MiYDg
+3F7A1ihikfPPKezxVe2VGl+Niug/xboRLiIJWAj1q+VgSQIvVqZx+gPGRbI
KcSb0OCxBCpfRzF/29CtWWvw29Lbm3LikMhMSsBZTux4OstVYSsaF2zjgiyJ
0XGaU+b5u26tYf/rXbc7fTtQ15qvmnZfOtsIttMcRv1kj04rjx34hZCLnHF0
eRm0DCJreA5gS9EvrA2Em6PwhwGiheM1yblfQDqn7JY+K90/lD5aE0KqMrlc
ArTLWApLRp2OXihXZ4ftpsrpGPUoREBAR19dGzyPu2fgoEbtY122wLnrMkyx
OcTftXifWUpLSKqythtiLuUDVzLQ06p+cxHuJ5Ym1EQnrPVKAVmqpPlrnG18
dPWzcx0/d49+vFE3jEktUOk5F+CJhutnVxzwpEuop6CAFcU8/wH/OtHA+w8w
ZJEKvMgdUpDJuDuk6Vc7vSvjxYKbSSqAzUvuwRbtHbloeMAAK6mXMwR2fc/U
Wq1bWdPqoS4nFe1jj7RokRRO5Cp7o3rV2atFzhlsuS2i640ZDur2oMG2X7fV
CtHfcI/Vl0DDPH/2qsVSqgzpT+bzpb6pa7kdF0kkm+OqA+W65uKCRRuLt63H
iKi1n/Do7h2vj+eBZmL0J0NNDzo5eyv46DgacuoPDHR4vP1mLekaMcVc0jj9
5n/H4J5l9rvB/9UcxDTcF9yBR9vdzVOSNG/L2s83z10gXZow/znrjr6DGhQH
AONMaqN+z09vDoF4f3G70aBci6uD4OJUBo8LVMqzL3Epu5mWH9L1IDExIHoB
nWT1+FY9oQHbdlzuFyXN/wTfmjIubNdvdESKsE5QoW1e6ijOhPTOSb6z5stn
aceIROTQdfkUZKlPA0pir9NyKcfyLsPRXFis7+ZLIfJsf6q3d9p3mHqVYE2f
rPIfifsEadZ+nJaB97OtVNG8A0AiLxybUp7XKvgESZ3FGOZXIfCWWiaC+bHI
qRFYc5ntsznwZXnPE/UrJ8nqQmRO0WSIxjYeCx/WC4Xl+YmRdOxn+JuuFNXh
duApbz5I94IcQMYxWTlIUr/M/R+FAjY2V/3BoCrTG/Kizxdubzsh6+h26Uev
82gMhWhxoVsaQXo1zZ8jSuJ+QJdB1IZYvM0ysRLjWyoo8RRKCvdjTpe8hW6X
q/3/fwHDNJeD9pfQb+G1M8Nb8ixtjoyy/HdxzWjI6vgygAT8kqAjVukKhCNI
y5YD91fn03wLVR2IMljAbUl5615IV1dSnpblB4v1MAlnuvBzj+D7U3c7eKcm
E6a06HSKNlZ7egnh1vFP6IaI3cy1Hyi3PggHpsymCNgjSwO+c5kYEPDet4ax
wT2DQT+GPuoHQPO2rjTThuPQWr7HkO8UufOPjgpIZwgBko+GkiThgo/y8eFr
3GaGrUwfv3OOMmChttRpcfKLYUoYrJpnPTFwXOrNXAt1KAPMFvXRlO7tXB8t
BoyUgG8FNFGMsg+Q7Ro+Yncs8Ur12OCV20ETcRuNOUxkpNI2MNsv7sukKVIG
f/AP2I1bZAMWRZ4QagE7ZvHLMIlCJ6HzaRcByCbxmeAVuAm4PyV9zOGU/ene
MIoWFqBpEFgMYnkrIDN3u8FfXYYxZ9Il6q1HdWa7bN9/6na9sc052NllG+jB
7YYmV9BsIpyIFLi0UiEAq3poM/N0NIVqxs5mKAdkaCzng75XEGYUDMUe6G99
XK583xM5z9hlgkWFTyTdiCwgbxbVWCYgitFWlWeua2BVs/y9H+6uhSD+Ku40
NLhBmOyEkOXjLQFY31y8jRkKOMsTd3WOjIh907ZPkI6itTEbRnNQKaX3yZzO
F3Q4Qj3+7hqLtPkfEmgk/eqTeyvvxja9oujRiyXDh9pJszyl0O8M+1zC3iov
pFInmVodoL+Zjq2uZwamTWufqM8MREFQ/Ae73p7UdajX5RTFEtqHfqW5j9ve
IxkHe7x/Sc/l0mSYPI1L3dRBD1QIsn/xpziPleIav2cM6uLtiFpxSmb56EC5
8MCzGtK7d51VkrLzPOm9g0Thn7HNJ6Rc6OffeCZLtWlpmoK2btNIJDjcrk0Z
3g+eSQ7KL1KUesDNgjhrs4dG4/lzQSoa3B8xkuLnWixRc1zL1fTxLtaqP4qc
noWYKyoEXxvdcELx3O3FEq3onSYwYrDsfugSqLR9NYe3Nsg7XRb7MiyU7iVa
GV0E8AHwILlonrdgsIjbvltGMHZQjCyKCncw19I4AyAUSKB0SPy6e9IDVgtk
7/pGC0tPtXVyDlZKCiFESXPYlUkL7I3dJLHdz+8PAw0nUrULt9Nx5zGObsdd
vKfd3rPJhMfAPsgLac/38qDm0wmASHIla+GKKVUpbIr5bLbTPMdojxuz9IGd
+h3V0k6nNDvbcfOoo3siRVejjPol06mTF++ScFhMfAsx5b6janQX9IP/s7SN
2OiYZMnIdTjjK0deC2Uth5foeyBOpDLZqid8OFlrf8EAym10IHexXOcd7Jln
j9ldmnPHrKm1bEIYuDzoLtB/6iZxfh+ef0qhu9jN5k/OOtwNjaMwYO7qZ9PQ
SZw0D0b3lTGCBkmO5nIxesStZCtzv9iNQ4wGGA0xZzwDiGRklYVXvLC9LAm7
unT56m/Kse+xXlVe6TPruSZAZIEwgrXPskA/Pkc4kVKNLMyhOSURrWxVE5g2
R+z8rvL26wcqEn+1nuqKbde276JgQ2n2YT9YYwj/f46gkwCs8STevfe6dO6r
0acaCWJRZTik2nI78E5ZtN7KI6O56C2WkW/EKDobJcR/ztqmqBgZoQrofBwE
uMz4kibGveuBwUo/8gDLnEe3EDGlx1qkFGCJ1jsBZZDWy5LVM67BEM1y0f/N
pVUzKvyNY6PffaOfv2qIo5J5bboR79un0K6k3oZ/O1ETTOV5+RexzDJRQ6mr
6DHIt3mfKbCBg1h8XI+6pr5vIJkxaPryMJ477wPogbJjTezSbdkYaivCG9m5
8QCuL9oxdl91EJtXO7sQMD0gzJGWNIdvPpmj+9GQUv+xJ/9BQdVQ31uLFsx1
ab8DcqydojLH4HxGw+XAf/dJR+E9sW46s/FTWqs051IgmFJBMaIHY4Q0hQZd
LxVV6E0P+1s3pc4thLHcIB2ma16gOM9kxZhdn+bhg+XakunN4Y3+wraGJ6b4
3xCy/O3iV5kUtHBfmN9rzr3e9s0Y3IyLVOyEBYw8ZnbFQvqZ3wrehyOw7mgN
b5PnBZm9RnoCn9dOyZpuLcTAflqMiHAghygyPfR0fLWWCghx3PRE472NDIzk
b1Z6xecHNiWIirNQzk4InTqqoXx+rATFzmkzEHKPj8lLC0VH4u5BHgOpC4sQ
ckz/9ujCxwPRPyzKeNnFPxq5enpMVhK/ONSKI9Nzp8itV9zDXMQ2ZhTRmFKV
l+iQvKYiXENY1yJz601svMcQl/4VoGx2YqsIBXCZpNdnxh2sQeu929GPypUV
z/E9QH4NkRgSklOQW2pszokWFQhCQpXu/FrUDxRjatj+aljg1CXv3VCUPM7R
CKXfBD6RcdfWymXQQnYMmXxgUgq9woYvQ0OQdgon98TLw0WrjPS2ynzlA0vL
EecTxvjiim8/vnFJ6wRrKeCnIP7cDuywXSNYA4Ln1XZ5ooMknNK6DzFwvS7L
gM5pQOxtYKx/ihYQA7H4HBsEbglssrSCZCiK/6YhP09K3KLsq3+Gh1KEAUUR
7zRZoWKrQykf33VIXcJ8USaSCKU71ZH0WKglJ9oHddpkiHOB1pDncdm3U76R
HCVsYTAFSFKsoqJWMuB60z1ICCvsF0zwyH6q1Sy3RIr32gWaDrpDJL0+Qq3n
7Fvu8nAP8byNAaxvfN4gPjnY6P1KmbmxxTnDeb+dEZda/lYs61McjzXe1ZrG
nXMBqcnpZr1sgiqbm+6arl0sm6f6EWbT5DvtY2aJriz8M/07UzF7xPemqBtm
uRvZY6ndPMZr3O0gYZcs3fG3ChkAUoq4DNN3/XGjPDtItnZTjfiTonxDHWra
vKwg3CtH8Xvc/2yGKYpI+7bTxH54WVgt1OMlh8wr4QiFNhPUiAOgBr2yV8Fa
6PjqHmgTgizrF1JYGbSR1DtywLO/tGohsQu7vp5Qgc3RmBi2k7Si6YH3Hrpa
JkBiRm2qGwlywxZCMdJD77IcY3ulCabhLu/+AtxznNI+V4Fa69HobwRGTxQF
PqT3doEKOL1Fq+Fadxsq7BF3BBzFDHNqNAK3SYbZTYwhWsQDADzrptNRKdR1
UsDr4oztclRpXys9n7+1ooD5viVMkFfwEK5ZPVRQ/LuvU8ABJsPuTgIfWznv
LgEoJOaAiPR6l/A2VtWMWAyYVi8W2FkHPyL4Lm8GgHmJXmf/1kV+6CLMSPtP
2sPuekawW6gbtDCz0sjKgYBxhxlrTIDpqFhE1KKoHDkP9nWgsecUP7QvEEnY
w7DGv7hC8i1ZOKKUH0apgcdoU8x4jBXzhTwbqybiYTAM5th1fUh+eIZt1JiX
yJ4ZaFpX9advmQC3aeP2ne4l5nuQYjNclmNB9OasEtcBLHl/Lg+9muK5GUg4
UCBIZLp91BzdxKGkm/z4eecE0+iTfikVY70zKo3hHKIh1U7r8t6lnfrXdSAO
kVGH1j6sCAv/Mfwi8g1lXVBOuRXf84eQW9/khNRDo8DTuTycYW0F5rqiMIf5
n4E0sJCFVVT2dF5oIVCX2iVPnVNyyduE6rk69QNuBtva483vaaGkzY4oO/nI
wtLtiHUkhiYnw4gJEXfH+mibTiAZMaqmPHe2LdW+x75UcUufUZDO7kplr9q9
U3vjIwXzOHltTQSX0DeZFVmfqOz7aedAHUgQlMrxsfR5toC2BxNijaMoLsYr
rcThyuLxJkiYM8UY8eEZg4eu5+3XI3QvvdBOz9qXBcZPd/KJdLzWJtGmBdmV
Rk2ruxy5kw2sPaezEldhX0KBLEG9jWzJZSNp3i/bRkJbtbwgwiEonYCa2fph
IiME6qsUeTgKs4ZrqVd6kEEg16PpHtdi4YEmer5ZV9dPS7a8F8D0n7DJPb9h
WE6HDF6eskgHfuwp37HjTM5a58Z7++8v1sJ48WVTXBj+0Ep+Y18LhF6jScZa
1Cc0YUZVwRuMX1G/YRIy+3zHIQuQt1otuftM4eTC0WlW8D4u1+hQFL+/df9L
t2+WAyHf0ybUNsTkNKgqHZnRaXWkdPqQMS7eZXXh/juAo0G5H+9S/egbJHek
lyDXJPtrr/HRDIXHHGhyVhK+/83/dSYWgRWxpFOJb/IlneJZOFawBU6RFsWU
G+5UTsJfB0SxijS0TDIK62ty38dFwk/hcNxvxdAZO8tpsHzfIhHzk612jxYf
4Ezy3AjW8734JEJu2xBcR3MJrgymQ6ssYk0IUOIqRTls7IiKEu61xw6avaL7
eaMMZjhTE51KL5g3UDGRhutSdlsApiFTGOMPbnR13S3C1vDeGgMPL8cashT/
NwYb1TiI7D+HUQ3XnKopHBRUvS3GDPxs2vyNf0bCWSI6xix9Pb7kxn1u8Lw0
v0WKHGoEoiBZq63kUVn0z4XsDPnXjn7lK+JfiPaJwz1psmjt0Jt8f8QJHq3a
hQjgRY+uL6NZz1lKKXPYr2HBYGTFCA6EFoUTij/3z3mThxGAJ0RO+KWewwJm
oqvw/s3Pahr/XyyRHVaUJttnxEtbefxpb5iV0vmsH5Hj/QB7nZYHpox7c0fB
E9983DiglH7kpGOngKT44MF7tTax1PrpwtybCq0Y0gH2vqbEYvVWphUwXfo+
V6vOi9q+ED5e+Fy6urjjJMRmNUJXCSQLu3SCCeXji9P0p6wvbmMY8PWzZXkI
m3Bv2U62fH1bw7vQCosFYGAON/uiitTdaxTdmpaUGLLRSqPHjwAHFXYWEQf6
HvlE95bak+8fvzqIefDHU89UGMO43kBDo/WsR/enTI4inxSkfAOa5EXtboxL
G645GtDwn9lPYYlFbKLBTj1s1vcLsLF0I69/zPflki8NgOo8x0aeNPX0hYYs
khxvUjoX9y6IC6JDKV/wTyZchQlqkfEF5jeNw14IuLK1Hw5i8iJAV/fjW+yw
FzTXZkqWcpa5Qq3fsuGQ9Vy5wVO07Ds8/gRAFbOAEMhNXAIsayKqJVJD6gHs
tXiLl6llkHSwFEbmSPIBjBQWjEuX2YqJ4g9JlHIrEVG2Aq7XUE7BiaVGSL1B
OvzJ7Ft26ksnBlEe1jOLnkqxvO5V+5rO59+vqvC33/fzPXeCWz6WgXHVIyja
E5BKXhJDWpqJMVle/dx5xWed1OtYMX6YMJSWnR74lAGVtIfrZ24JWgMf39ga
NRKhHoQoDdT2EQzN5+4jBMr2QdEMXp1NeYVXUlJDn/ktKbcpCntGbmE5i9t2
93f369z0xVjRUqTrYTlYkPHMhYa1NPJa3tv82bdnNxwMuqjLwKt+RxFAKFd8
Y30bjSfYj6WmgLAOIWDAwKBtxlePvkFHhKFgf6GWN5gmqMXNQ8UO9lNAgw5K
JU8QaDnPJzPLfqo/AEezMeccr4ywIdJuUssie1a4FCDVdGExYfY0er2X/NZG
3st+oj3nv4zX6knVDtQuOtT8QZIqEvPYkXSpdKFXd1wjHp3l1HzUKUDi9w+V
LvwfIU2L4qkLN8ISy4IsU9fLWgI0Bt8MiV33pJ1zInoTXT0ubgl9qEr+zsue
/TObyhdPToQvjIoHuheNWpyhLHCo8h5lddfg0e/rTFJbY4XrWzBEGqriSEM6
JeBfWjj3CU98eOOrjDpxOeETTq1xYFSWOYOMev9fb5APrC5uV66YqFA6m5t8
YknD2ql5eKfEzYZ5h8XL0NyI/dUmsrfnejnpYXb2mdAVNymbKeoJvx8qoOuJ
ow8s5+oUDfDDz1hlz4aZZAf6ft82qYzAyRV4eyDVLv9bQ4DGPSqBZZ+0MPnA
A2GppJGJRr5TPu1/rosWqtJpi5omIzYvk8RBDQXko+er1+n9VccwedqOhUME
FKcdIkx4wJbFnlx3F34OeOLFaX6NYbTl4na2GRaYUWvTEkgzKglYj79+lPPe
thOQW58YtH93PIR3IxShtIVFA7/lYbnhglw9atnapmBrgsiU+1eUdUiI/7bq
r+WkxMHv4SRIdwkH7r5xtLv1bPQthWiEJaJc1JC/OVRnHA8sSTdQE60TJSed
IJsETmghlYMJC0YmA1RY9rcalkN0XAgy3fdvgnJ/7JfiEqYLshJYXq0O4Pu9
OVkK20Jr7oU3iOHuHpbBfY7BtNKoOxNEvf7RkGj7dGbBdRfYXQAwudyQM3W1
1wl1/21O6+hodq6n397HDdMqQWsJMJ3C6Jr+FYFxfcPFIjHgHxMsSFyqgPKe
xCG6aUyXCslGFRCvL9r00Hqi2WZ7fxL9gEzcBrgw2TNgatpI4YFuVXnmzq2p
YBJI89OveWfWb0cR/xE2onESmVLF1zky2E22aD+9Su5AP9/UrymuYqVhxfXo
Q1zGCFsnIKGKgzUmihPEdymTKNAMzz5QGWjixE+xZllWWe9yYBssUZathJp/
aPiXG05p0iL/zlmelIbeo89XuV5KhfK19Rqh1EL8y0v7/BvZ896YbZISJAqS
chLg5hElKTmxMY4ldaF9VhrDRe/eoXJ38VpSgtZrBLy9kzZa/3zUNM1Bwt2r
tLa9vH2DFBysJ7l4tGPCFVFzsKBiRqFiOJkpjLaGAF7acJEmkLtm+U2YeHQV
HtMkOJdGD0bgCjdnua5nQOeTkQECsWt2V3PYGz31usH6+r6jZqISLFffsVD0
qEPuNBexxgko5l+6otxicD2jAskrJwWKc0DsYmrD1NdbUUahRtE/5tG6wh67
G9vA3TR//G/X/QOhY8KjgNaSokMU3ITt3k9e3SBAzTdCHjn5N9f+/1f0H6WG
+3Q4uheV3Pcfk8HJdA+6CHwL+93iz4WSpjojm3OuLKPFIE7hH7RiQBynG6Pt
4VbLmb+CODMHqRsUsbyxKo41SXddf4SFiJ6ivX4X7HEl2V4iEmfupdEG5KR8
EyuwZUpZxgSMcEhmmaBJpyQsA8++yfkUq3kiIGENlbmFiHd0XSDlWao8IcMB
eAC0YIJMx1Ln/7fzWJgJbMiJ42U/83qEEp26hGtWrDsyEHMblikGKNwZZqRa
TC6yUTIFuMC74bQfodIzeofOjtRj9vxeUW74Fsq1nWexL79B6jViu1MGtLsN
iP+Ceo3v8D7UmBlPSCi9cFi2VyNrrleNPSfEMKkftO5eZI5ucn/pphADS+ED
9b/Nusvirmg2WU1/sjjY2m6EzCv6WZZWfM2b5JMSYpxLCXcsFvM3eaovpdKD
IIkbMrbRCtOoxAagx8y5XnPLDC6EIgCEMuq31FZHlpIBaTusesXATaJPqwli
Eb7xXezNY8FTpzP/EuZaDNJxICy4DOxn38iRvTBijFWtKQ2VrQbgMnR63NQ2
aFK6vgg7yBQ9Vs4yY5lwsoSCq5aLeJFvMExve/GbBMWXv1j1mAXycZJr4zcO
jix4mnpHgg1EjjFT6n9VB+ISlJhmyvzh7Fzo+nxvyh+Rv5i4wUBHNK20zXab
twujmsq+EOMCc9apWd7lem/b2ammscezjMygoSiE92egbKYfBSiS7EGPACP4
mNURimuu0GoHz/V81OD5D0vX/LtRzifLSHyg/kuL5eaQVsAURBJOb6rAgtgV
vJp6d6yeErg1E43eF9iHo8T1/iFyhI04BP9j3/j0uqGbkCF+n9PkcUI5Qn96
24GNIn+MeM2tDpNkGjZbAwyDU/bfS+jYPkgwBCU0nVzZi9L/l0BQ+BlgAgN4
8mhR33jtH43TaU/EfTssp095mcrbrPQZXzBjFeOarrJFEnvtOyut4zG390b3
kYHfutq6pWWNjX27F06sBUeHvGYhGWv1BX5G0GrQ9yEG9F87xsxZtZTMsHn4
8vHSuIoNin/FxTKwrn1Bm02X329gC/A4kQI0dwbpa9FC0w+mx/vVuGPXlKDP
5rVQByLtsAmUbJWaHwgqs7SQIBrKeyWDP3B5Nv5l/Bhj6Mg7tXQXzg8iGcLE
d36XIqbk/XxFNDYpe7tOMFwRdf2qhIowmwMrxxcJhi5xDjlKs9qZBShcwPU4
80Y0cO6SmSfeAn7EvBKy+mCU6RHttlY3u9r3I8B/ER67GP3fa8nmuDt8fm1K
Ij+PDVz2iFXJZyRhvyMZ2YsC1mWP9r8tl6sHKo/46r91JSDfaw9OBh+KUy0W
DtLq7XYRr3SpYNqJ3gmMwlXi3NowLavTznyUYJaBl5rLkHr2tlzQLHmJhLu2
5q/KiXvSLszOJRBKqOFByXL+3i2n+od2YBJqHsg9T7cZcREUbKWTpZzTw1jl
QDZKbUieuNV+IPFgikNKSRdMx57F/vUxDJRqOv6lyfzDlILWrdfMWhl7EXLW
gaGL1R8Tjw6RcMD34oI5yi9B9MSvgBlhjkLJ19LNpu/h6j7IJHnP47gQa2Vq
udqJPxUnj7QB6CfGOfjJn4r1L7qevwOE7hjtq3NVHQQvO1AhG/AQfT8yWFKa
yvK1jU54/8jL11tGXsNga40X4MGnwLoiH8kajNJwWknmfeHvLXcl3ZkRxrCX
UgEj7zDXvJq3kmBQ+khVtzpkZd74iIy8W4+wZtORgNAL5doDOGvQ/Q7If9RL
jF0mDfOFBoIK8sV33aT1wv5zQLLa8MmJ6FIbGWQ/Vrl5ph4UZn2UTZl89z0U
MsLkYSMjsBVrw6m0FeKuNf3DkNHha0kxEfkZ0fiJv6mAH2t7mj5RxMXM0Aok
wSq8qb9ewhW+8DYxJAHBZuJkCYUbaw7FGG3RszvXqyT7PRpr9GMB7glBpqK1
mlTJ0vV/ahoHFY0NGluUGSW/v9mxYJ9w+vX5acZ1/WqGc7OL44TJPkHuYCRv
8LC373xf5mfGfhALPksdv/iybsZos0V0YTKOX9VKDIbLRtN7PUH+LwS7+U7a
nhhUzHN8a9cPaw8AqYW8Zjuz4EPAwa2qpjXFja2lAg69d9nwpIeAbBwu8fEj
YWDUQMOCSm8ePUGNPaUi4X2iAkAgbqIYsLOM/TE+lLEIS5jC7cOOOEs29peF
XeB2566/WNZQstHPfNWNzqbUMwZJrb0ml6/DGxYrJOLPlXbgi57+eHeL5k12
zYveRcDBcEPrr0C3niUEe3viRmZIKKdV9smNN2J+/hWwzJKKXyACEBYd548Q
+yFWpDX84V6suykogdIwVZ3dhYbalGdyyLFx2US2Ab3NlU314G8ROrpxQ49n
+TDfJvityCc4dG0gdvHR9y11WrIODs1fN+WHssbN9U1wGsX7aFuBseD/3ZAu
ko/WX6cd0TbXiydZJFHFhIQ+HpaDl0A5YwvgZxSn+U6txSTD7pmK6GROWIPq
hvOrdRIsH6QD0wPWCbJ96xphDN3Nj9ByAiYaruhfL5ouiig1QmIAo+1t40pi
v3uVaFNKDpo58/kFTEmGyMsMCnBqUIBYhz5fn1MxUCGD217F6SiuO1QQITiD
4ZR9FWmwItJmad/qGmEr8fdHlq31IVSsJFwbpJrYEYDKZncrbvZdY02Hs2hl
cqD2UGj4JiKidkbj38D9RMQMJCPvAe4qnsKYu4QtTyJsB0L4urkQa/EwqEBS
W3VLljSk5ka41seWdYUI31njVaRzRhZa7bNYXslchkWA2I9yDvfd0BNULIK+
y2qrikaBHsWtq5lxY4dulyeH4M23+3RfLHeQP5kpCT6hMInCFOTYrTKuOBnC
cG7t0kVPg9NxCfrK0QjuD54wYvCm7nIIuhn3M19b37oeRtY0pviTVdw2T+sQ
Gw9mBzsj5wu7zq9OuCvcP+kmlVrDe5F/DoJOWp2s5Ze0hhaDVU4CyVz/HOyt
70kVpSUSqaepxLxl62cicgdFKpPf6kqbWhbZDEOp8EEejegF7XJr0X8br96e
ek8LyiDStER4i9x4vbmnnH6cq+WRU3JM0z8U33RnQMhopdfyuIqZnF15IKzx
L3+ckAh2Bxr8iEmAENg1gv5ot8WhFXMUjCP8XdClIwg9dIHTkFRGAzLvdCMq
Owh8IFvw1JnQp8CQWN1rgwFaeM9L0YyYT/Xo+nopjjcC20uTuWrYX0Ya60IL
cOo9XNNWhGUsg9nw4O9Z5Qo29VWuZeUkXjxSJrEQJnEM7UzCpCf/tVpVDldh
mHrRPJc8qR+rzYwRryd11ERiXDkVCKgT7FbKxks5/l4I604oQvmoW+u0T7di
qJdlX6pFG6Qx4JcvD/Lz5beWxFjFy7/RLJoBjzMmYEQu71IsEEiqnS+FiJKW
Mor6fglwCWowTdpPMmWFkY2KClWNjbjohXunSMENc4fbHIsMvPP20620jUMt
YKeoRvBvHhbNA1pv+4jCWLkbRhxiCyCfQLiLtACGNs3BdjWNu6mA6H+ImX9Q
Wxoxm+h42inynwvfLhJnh8P13eVG1hjZCBq5uAdHDQYeiBXnFcmtDAJFo+/V
oXJiLK2HcH2T/Uf5NPnYUY5LUczxtsT3By+udI+/AhCCFDQ1GcEYhP6Z5U2w
mHdAcyOt18p3367k5vVighz/AWtLGvcrZDuR+u3kBaI+jPy0JjQPJlaqlfWF
pIqLGAH7+erMPTmDkUqAU+rP/kE8wYcKIPdVVfaNgHjBAHIeVpWChxUe21Zx
2uvxBPGblN1ED9uhLD0q/0ncZPxSq2y+SoGmcejBh0ltcgt7git00vX0K0+k
HBviZZ9fyQ6v/oQZFkrxmn+B+HUSDgEeIPhBVB50flWo7bp8d5AZ7HvnigZT
CnOwT+yEs5ey0+NELmTHTIqdU0FoFzr6Q+MalYQFahSTM1s+GrF6OsfWsVlw
mYRlS7JtTZpjv/2X+R2je7XiO9un09G7+jScYfiI6OI25bYAaov4j/I2WvJ3
pdCfOVn6ZsQOM/TTL0D81WoAZVwosT0ohiE0hYIveAtD+EXEa+ZRHvaQDj0U
HAqh+5QVuMnzgUx9DVVHQXsoUIz32FJZpF5ogXMx2TRNjcE76XzppJlOn/2x
1K+10VRq2ecPw9epG0PBSd90fO9jv/k/5cHku/r1lcsReHlC8URGnswvFt1K
iM170lG+C+qELs4diuJRhCJN8YLgMjnxNSlGHqZm3FEolmlA0ABsx2zVXHWW
nLaoRS55VZuGznFTKUfdd4bnmj5b6a86al/fG0hyJ3w2s8lTVKmY1bZyvb3R
mmLduQ8Z516n4fH4eMhNiGxr/W0QemcWbdP+YVpc/4DRE6ND4+UsPRxP+7mY
4bGE2zW5E7t+Mz0cXhhseTvTYlYydRvoHTfyCWw4ZozFhOI9w4nNA4asDIuG
jR1qVJohYsEBR7jebgPctX0ouLmjk2gXyzY+WXgeEMoeoTWjMgpo3wrA8QGM
JyiDUx3/SudZwAfEkU0Ex5bWp8AnOLhe0+DESIBbTquk/Wl1+F+fohnTI/4G
FXT7Z+JlPl+DeEtLMzQkqTizLvWTjEybdyMcHepf8fiXXP8XtKbeag2Rh8/C
NToHQL0sciv/4YXTadFXK121q7Vqo7SqVaZFAtdMmpXvWYl1PloD5xX4zsPi
8hmpaGULjpyotmnWPKpz7T8cI/77+7RtGYqvbfOHQEh9/UGRcShPP8WO4h0d
7zWFwUgm8hXkghWYjGfB3X95D6sVkr3OVgftdw9l/DEmGJdUPQF8Ll9362bm
Lqc1r93Y80GKe1m8UCYVQeRSdAMBKcArftVdMRf1+HshaRP58Iuz7+vIWFUY
c6wIs4H0ZHvVBOIz/iXUIoJA9SSBD5ZILnCp1cCPCBFuGWmRZ+r2Uol21Zs6
+O64rcJgvrYUgcBT4ZIeabWsyZAwzolHksbOYDoZjoO5KcR1usVm93wHOTKZ
D962B7ByZFdz9TkX9szEZyQbXVzVepaW7pCuG5wYHQ6PD6ojLLm/0TbxsPWI
SD0xg/ZIDk6XtjfeW/WYMtk5QeztPv8Hse7y3KOZdEdQk/41smST3OZ6k+YP
AC3gJ4Q/AbFbaQtbF5lD8hNOSddQ9pdaaCdAM5olAHLF2Bgf22+XFVeBa8PZ
+WRQHOoAsNaLOZOZ4HJRe9vaupgwp0tBm0ifUjm+5LEt2Q5/KgcHTmfykTC8
TnnNv9jsKUAg0GGdJKzU9PlJVGIbwYxxqFcbpDCH6PAqJYqdRMlaxzqqyXt8
n3/KPg0OFZSc1ZKy8P5efuw9gxEHK3nSFaTLNzzngEDEVcZuoHK8xhD01jAw
pguXiXYNEmjYVoM027qD8ws7RnfeZwnnW4CQY2xa7qpONrarJ2C/jER278TH
W99N6etm1XDna0S/FV54yJQWMkI8RnvJ/WDWCak69dnfUD0BRgro8QwUONao
OTiw8QBCGg3/M0QdU4b7rRET9c+icXCHuZlJUd8c9eBZ+Md93umti1tMcE9A
iTguW069ls22wlsymiubGG3CTctks/nPPX+rod2mOFk6nY11DWG4lhDEf0cx
cccwpi/Y+msGfr6fYgO2Vs7eJAxVSMiUgtq968OQX48XeZbfu5a7H/q9C/Ux
4K1j6yIaLp1k6ef+FRKyJ2KRqfXa13a/dmsgOaRN/xvjER05E/CcnfIplSMd
hpAK+x7+PsfGIDLIBzGUCwGUwo3LXOPueMgRhLzpMkdOgoqqg+QZcRy8D8UV
XsO7XkE6cGh7ouYra9AMsVOFSUx6bgEUg2/sufm/fJObsmyjC26vWdwIgCPv
+/ctXo4yNmABxqZqbL3uKROeXwoJAh92GZ82w2FOZmgd/BaWopxJxpHJnya3
guM7/hX99sxv730pqbA7giJMLXns6XshKW/OzpN0zi0Yq/ZQ6FrqMdw1fGXF
HbGLuAVf5Ddev1LKsQSMqLwkK+qtXLklh/4smHvVxYctD5U8lBArkqJnYm1s
3j2wLKbrrQNTgseQiqV3d6FXZPjOqddNO1e+Y96T7cLJCgtiXBwjL0zuV/9V
K4WWMtwTSWb4uYOXVnqXS8u2V/WuXjddnzfxzJ7G70TuDphghtlR91EcBJ/7
PC0VYi+2pza2ircOj5rcvx2aUYxmUXQNNlCYgchzXB/ZUD3PXkp3nsBWAkd2
5GW45vvH7ix/aLLpHW7pTXN8XFh/NDfQydhpheVEcBAH5halb636AWzeDTTj
4MqC61L3no5NEpvy9vrVKk9x7tc38u2ujOxsdVTQN69W0ORjeGN0+sQUBEKE
PusiSXaoRXhcioH/7b92nDLrV57WHGwVXTfaW62937SkdXboXlNeI1CgYiAO
/mdyaJHQE86YNSaiW3oPG5k9RCAfmLivqTcnWXMsnysvvxGLdbkrgxonyTJV
MPrN3Pz5GuAVSnNchiMc/pPn59UdxJwY25y23EcvKCvQyZr/FAVJ+2hG8cye
doYvDhSFkkHfvR8QqPe9cD3sjl3UPMXRp/auOU35J/B6NgkPRcK8Wt5kdOZd
GXVL6koJBqUAeLMsynagcLZufcEpXw1h2mEOBZmlsDJrLRixmIcCFKSgX8Gv
OfZH8r5gSI2pWs5EqAhlF9cyIUtu9S+l8YWjB6uddYOjgkcSuI+cJos22jcB
h6r+6QmxV1cTNdubxjBqPrQ2cGvieXWMQFu6QKr7BHaqNyFH/xOZymPs6zsj
LH5JusiK/is4E8iyh76HZjXdw8L5NB4K98fdH+mRdWH0QLUf+zsyS3x74Df4
gSZw/JLUk6tyGRG5HIK/QleSV7ISFgdMgow7cZRHNrAeUZGf0w1ArRx7dwTe
de1NPVuPHM8ReLylQwaV3QfoG2d6yzCaGkHhwnIq716x3WI7fijgN3xF9lh0
XL5Sw/2zHJlheZ2E9qv85yTJ0g8ToKkkhjINnJ0IHro5LNTdgV/Lz16H3s5I
a5PHpGCAvQbbyxKe3FFLtKyjVO0kd1S8vfaCh3oK0+ohxyT/xT05rpWF8nLX
8qkiw7+TqWYHww2lT8/ZcOi6lg4AsoDQgRX/kYvipx2vNTw9Djg7T/LKXP0b
jraGsfAXWg6dEtdjwwwwWzofb+BBpIdTb2oNFMhS1un07bR4EzFmbdIVx3XN
BzuHYLcC6WQANaFueyWndgYwEz2N4K+RGph0GC316oAUSVWGIXYHhKRmoLwz
bLxa7WSUmJCh3Enw57ba36nNJQpzqsThBrJX5iQ8kuzAxoa7ShojlD4/4LdA
/yqiIFh8+Ty9udYsGniCo7R9nph0STZD1rR6x5GRSijo++AcReKU2vzEYU2s
TaxcY9zxH/UKJ6AY6CLR4BpEHJ05nmAqvqhEXP0Nn6yENsfkHNJiKVmkaNEL
lZ8ufKjyWoNghp8dEnX7sMGugqDD9/5wsAZ3UgjS+mD/XWA6SPLbJSsOUMOa
ivlIJe5UUnenj7hiT7nbqMPl7EFE43uYiv2smLj1KZm2GBgMNZ2i7I6GlZJ+
QKKb+G3FKzNN2Q/VBTW1eyIVQXI5Zs+RVzDdg7UThZL9bFvZ3mNo1UJm9ESj
Sm8PvyCIznbZG/mlD6Mlg/n7s++wOgA+BJyZ97N6r+hwPCcHMBXiOP4SFw3h
B+ubS02XujdGtI5/mP2CMJVKLkU6rnYlyjJYBIC2+Hn4K3RzJyd7RekD3YoI
zo8dQwIFl9U4OjzA9Az3ZlCFyXCAJ0Pl+3pOlYkRK4RJiq7RwmHbKw/xsiSD
peiL7QAZxNJWMuNaFvPap/jv2BOQjJqwDZxbJsUmgWNRYa1yX48b05xyuLn8
K5+Vcdktb+RNarWjV/vcjnhRX+cKQRAHN6k1jbTjbxOaQBE1L8CIGP5YGz9w
5s+bY+LV26lTMSXUeJcfAda6BpSqAaTqzgLUiJL+7boGNzS42iwR3UYnrbkm
Y5aji0iQI4GdWGSGCrIVPN/dkHHqqeNBhEV23y5v7gbHr8lOsWtEGHP6EZl4
Dxbe3iA+rZjXOw0u0mXc1hP0ywUzN4MJWxk3uxI0+dcAE4ZtWJoC66cdrB+g
wc7q5js/qxftWqc0Gk27eYcojT+oswo6tRfFumBVmY9QxtQUsubyfIlJGZTR
ir4xwnOCZ+RcW9Abo2JB/tMgpgCZj7ffuELAxYKpSKilTZBdeElN+RTSTk2/
oCXHV43oiGORan4TeaypfF4lU3PM6JM7cDnrlAdOgv5RiEWqKyN/KsYSZz4j
QPi5AKxTET3gbGE+qJ0PAZ8XX2/ezmpTC6MkLn3GRd3sLpoNUL0DVp1HKlfK
wCxdicFTfFDYKucXeQpHJegE502CmNSORbHFNHZtQwR49NIFKg+eRnT4Q1Zu
6NVyjwY8TEE+nLrUEpdNyXn8qjlKObOYoFlhYBwyxZwNjnNmgyNQ8R7kltxC
ibzLgAU2waedqkJ6s3L+ys4mysRgkIpLpVJ7cl4LTucCQPdGIEx2FKDe+xEY
LJ+CjZaqdfCWaAkVSj47lpKZxVaN+xGu9Y5cWsDrfPtMpgY4HCh2xLewPhow
9vcZ0pzWg+99ejCuEzcZT3QHSggT6zo46u4eUFJvqBGoEs/gyd59Z3pp3zVe
kQe/PmAZmSHXt6t7x3qqUwE4d3ZnEA7SEzCDXdVl+Po+3rP6IX39c1f8HoMy
mXOq+Fh9LXQRu1lH8yVOuqhiOJoAp7hy8owYRyUVwHrVxZaskqbQRwQ+B3l7
Lsb0w6/Zx4Kl4WRlQHJuX/D5obGaMDJd3YbSrFh/ItkbjYycaevKAIype1o/
Qwv2fKZD5XdIdwlpuu8J6NiG64bTRe8Kq69r155Ok7qqq8XLmFEl36EEnsDv
173fZMreG9zxQQPzssFR0LQh7owwo1Hl8+GByJy3Aydcxl7lmdm5Y+xoxv9Y
3u7EDmJE6cwKSbR1b13orNEHFSfRkan7hcXIDWWQ+m+Hl7v3hRmZgwaYJPOK
4XNqq83/J5rumsN10ZszD3KUFB+jWgDvIrGo63yXOcf2hDRyWG1gBVMkTDE/
/SQNcGqKpZZneSFjkWdyBGYw5fHOpcoAD4czeK9m1X+8XTI4yB5oiy11VWk8
ix74Fdb0NSu43qAnuwhsmBf61lPle1JbJf38zlLldMZSjKnR2f6wy1pD2eSP
8JWYjUSDDr7KaWW8azyYqdy3VII9ZaPJ6ly+6pqSXTVMfj4+QhBYdFcMcQ0g
afSWysoYBPq81SKaiBffGJThxIxR3ZRWrHunNNm8tLOiHaXRuRAovoVT9CMK
3+snmfeRY837FmCGI+amC0TjyclGj7kSSFgDuchPkoHSAftYQdBs33TzckH/
vLUWQNkV9kO3GyWqIZ0WPb18l7cLKgByM8expCXO2PRyo/AGx8poZRDJ0XCm
ceCG5a02UuzpkiqTf18QTpMuQaDJdElPwyf2mCJWujhYQmhmHwf09MQ86G2v
dEguEhI26fTOWUTT0OE63EdEYy+2tCqfM2mNH8FTYEzZnN5lSzDC7nu0vKHx
vZmWLBOAZ1L+KKpYDuRzFxGpc8Q1u1L05ffmv4b0ohPS7pFn1WPdjo3pHy1D
KAHi0vuMqWJJvwvbQYSFDcx2LxKPOy+TsLnU7nD2C9XzV1sD0Ls4/KUwwdiy
0adXxQAoav1IBLu79nYnJfOHGwZXgLBxDlJOMnSvJKciE87FfaiWn3Sh8/f1
jMqsr0qm6Z11BDVLuzm0JP+1GGz1duDc9p4UrS0AsnUBOVOLttKdCn2lNn/z
BRnqY2mpC4I7i+HUlHAE3G5ueR9CeZdbTqIwseNeBcOc3KiBVXGX2hHi3CAA
xDfajDpYirkdPqeSChnTKTbLfG+hiZIYI6TJCK2dB6XIMqCE0GJ6QMI+AKXo
r1FTm3g5OeF7FU/fJAppJY7zGKrYS8zviG6MM8QBc/8a+tdmqUQzLkimEab6
zz9qJC0StyRb0Htm1VtYqgPUTcchIpxX1uX5eLS/1S4voUXr1WdEkFKTINwo
AgBZKnSGHyUTtMDjcTbC+YyHRlXYASu2OZ83Pv1Go7XVZmOK4F007XUXvzyp
9jXO8DeqVtcBxaf3l1kz9gV4jGwPNWbS+gjQtAXRT63zI78/4al5wlKhsmul
oJqMzX5UtfqO5S01NNpJH1MzNxT/0qzeRn8Bmn4mGPQlTuu54ciumITfsljd
MforXCGjAjU+69tcu9DCoghCoLiEfYI25SOqnXkv5UVEpEEKOL94XdGtF2il
0jkXZzHYDmJZ10L3XtEwbG3zjYAAJbdfZSPfF8a7PfhxMH+K9w6bcfjkyGq6
l04xzO8lC37otq+v3kea7+X7P3Vr6KenQh6JKHc6Zdo52PugDIfhgSQSiDwV
m8PiWxj6pgUqHerl8iEy/Tz4ZaimGIyXvKGDfyLv79ac8ImAfvjNv7NWMv+V
9WZFgr6GhYgsG1yYqTNQDO3B1oFczFe5NKgaO/CAtFRnchin420KNbPXEazn
mFaZczXNChwxf624c9sYiqISvTa/5uG8q40uQIKBfItNK4cfiN1O28V32N5p
MxPm8RQzxy8p4QvZizLBqd4X0MMemHUH4Ud8ezRCAa8l51FwaQKCpcnTCvXi
kQPc4/hdAPUlgg3+ZIQWKFoe/3xKJr6fPKGsvQ8I2vtG3LQxY2AmK7oO0Wep
a87jrNkQoPvCSOPVXM2FFitpv9JxY66Z000GoWxNzsZhrb9p0jYXiYWgdvvi
X3QI1fCcOa0lOiqMFpxi/0cYIMgCfHuNCnQikW5WpMQ1deQKiluXLN7OPQfd
ic6LLL52DtlkKUyPSU1YxGQEi8zqTNxZRF5dwoU9F4MJTEPd/1eUCIZd+EN6
fURFVM/IcNjnOaAsBk2tWV88+U+p2DXvjF6dLLMlp8g7I/SkgiuKe+egBEs/
GRBvZ7tQKme3W4mdV3tmhGgrhXZ0oV2p8RjDl93BAagS2U0/U0PmcYAsSNXx
B80XLIrT9sxXhmJ/eCDMO/+chbQ4XeucV+czyDUoT4Sg4JZO0qeg1mElI+dn
3uba+TVG+0zbHXjRKzDxZYgqrBgTsyAUiJZ5QXxHldPtY93vuhmpbkJ8oGx7
393ZNAJziLEHyQhDwIdI0Sb+z3x2BDHkSt9urit74GvnxiXMpDvLxBK+wGY4
Yi+JNegAQYmjiTmfIngBRStZC78WD+kBdl1scsRKIj8EMk7acZwB4hNlGBes
LBCxoSvAI2WDIqn6jv2c3/caEX8ircioV0iPZnCc5qXYa7pCEtTuwz05+HhN
qUeKKS89g7I80/uggC9LxTrpaIgEri8MvyhzydhcGhCypYXVoIY9dLM/FIL/
iCMfTLArdus2V7LmJZBPCIWHG7CKOLvw/1XaG06YEKFz4Kqd2pqli1kov9SJ
qqcvMb3bqOpvjecUUUHtWxIj3VAGuizPbV/laYhZ9XWDgGYZqEN2NWylXhwF
aZG7o6urQegBjtdIQCi3TVRimRHYMOGr6sfqIXuKJJ4pPoRRPOauLnHZAtXd
B0LfjxSDulKAhyJAatDHzSSTT+0yLlyR7yEmoPkyXs/UbA2dZhyWbBkcdxl3
s1BYrFHp0jANYrDASaWZTvmzMgqMu6wjmpETIoFa3YKhTqT2PZhCFEy8h/MR
+kUAbdv3GFf4R0myofHSPYcl/YVWRuXT5ZX6LUfB6DnmaUBNigL79sQ8Quu5
fV9O3nXifIUURUCt8OciCFgddsopLB6OozZ1jaFQSqeYkzPyw9XTZeY4SPRm
rPnYgnS2A6dY4/pAZTuT+SLmf4sEN6z6UeKy0kPz3JDr8WFLq+D7reketVpz
wWxyAkQhihRzxUBHxlicLxKTHI+6hRdjXUMisOUBdrDGpiR0cFpsD1vGl9UZ
eUI7kUI7d2r0qyfvbnET59P4p9Q1DjnIXkPsk41E0f6eBbhfHZ1AmPOAJKWV
Guq/1i8XTusPGdVHPJnHEhn80/3rb4/xI4VHH4OZ8leH4nWD/i4oNGzSu2Qo
BPxoHwT70kg8yRu10kDx7LGcTJwqQhiiu21lBbzYh5zUQkI6PlczAAs3IuF9
GOJVZQexV5pbUe+BrooOaNo7Fj3X6ESlDG1erL4KluStbUeAyweDjDQNqEZS
9xCSEkCuzJGRDB1KsbxJPx2FALop2gHFfWqCdsIB4vnIhG/Wsld58HK54X+E
ve2vLLOGyNuWlbVj6i1EbcsS+bN1HTbk4mjbmdr17G5iEEkLMl7FBZpw65Qf
YN3tC1h9jM72VNKh6fddGd3X0FzMCJYQUKqPr85z/R7tKWazyOePT00X1Hjg
j2zSqVZU9xohLmySMUNDa8IvJtTE5qXePBUg/N0i3iuIlejiA/80Es7a5WFr
Y0Ar3soIw8MH/IG9oixsLCa3z+ijCFijEU8wpHwy9l923E0dP6MfgTbw3oFS
GYQ1i5OiQyeAjl/dgtT+9HRzhRA6src2Y3cDrno+d4JVz4XU8Bd8wHp4U0yZ
KZzkcW0Ny4oGPVOzcPw777ZxjOHZL+LahXowbVH66JgYxpykhgxjZ7yoJUPS
8AwRRrPOv1FKt9ifI31VGxJ0GSDwADNLlmZFMl1jkDhqRCHdK/NKL3nPKPLr
l1bCZxRKMgVceUDx0+G+QdnX471rt3Jo9H3ryUI6UpV4mKhU1gpXX6wwci6e
b99tWCo2IiBPvS+dhBUGHERwlDIfkzWTL3RwGhwbr2jSWbCt5ZtiGLG14Xao
K5iHu7oIYgssClY3Z6D7c3vKDrwaRgf0Ep9NO1iq8hIk3/j8UmnLvjl9wXBt
+6/6NxfiUnNcLQl7oxnR1gPkSUkbHShU0/uOO62S3sbRHZuqRUqu0bbBssXy
HdgKwg172UwECqeL1gemkjqYOxDI1yofaWt9/FIIKIXPPqy5NZVfmIA8reX7
+q7SgbUVO7Fnqv1M1n3igEetmtVcsvX/c/RbiTkKJjH7E3MiyEbiAm/3U+cX
1sLGNNldWkbkXRq41Grlvg29BoCFul7TLcNXeq4BhVf461xTd+XORPRLC9eu
3SJ7Dsi/lNsw3bvBh1UXx+KsyaVwI5sWbhIN2EhkY8GCRRKz7ukFT7kVNINW
3aG0gW+xT4/Bq651rClZijFr5XQzafRu/oBaCPma7h1oU8Yll+DlyK6enaSF
HYbn44fyNuiJVfim53A9lwhkrquksiDSAkkz5NCsfIjRIOJgyHhaE85AgAiq
DRNFCRQGLe1YXoXLWoyBSTWX3xEkfPbFZ8hNlEAUu7EbWLGOUe8LAe8cGwO4
9MdAs/4o9wF1Nga1tuAGFQfoeSeDxCd1JAoLBSI37hzKjDOK4Hq585HgGNI5
43fJEQ/Mfe5L4dE/Reon8OaH9Hk34AKG2Op1p41GnylfI4g5WBIcSXSoWvSi
HSRDW+txUgh7XEx6USxLAcOTWM8fLppl3DS5xEAZ7zAjuttnAkX9ksc7hgYd
UEk13VK9vGI0drcucV1xiVYEPQpEWAez8x0ibTA72DFBcHk/3Hu47RENOPTv
1UQxcvY9vno6lRo8eLqlPMWq11YOMjYb6fK+q83CNn8DBCSklT7jglGjRp6f
l5fk22eEgYWATQwIvXX1qxBx9SAPUdQMJ4J+j1/aP0D/xizKL1ZF3oRL1xWP
MS1VoFCBEhMKZILjEhstUWDHiG5dneoIvbpSx5yCDkDaVIvQSgMmEJL5sZhh
aoguVKA5y21OVjWQwTNZurk4Txu0wXbF9cUkNnGt3qnrPXlD1wFNOvHp30br
25b3ZBncaONsXEUDCDI/gjEG7S2RG0IjnUOz6Ky9DMvWCNPQruo4+zpcB4zF
rZcj9JasH5iV3ZFN3j4TspbGWkAt4tAuB9Savuxubfb8p9rkSlsrzbDQREj5
FQhSASpYTrTWX6KDV4MKK0r6tcsaTwX+y7x0+t74spXDB2r79QEeKO3Lf9Sk
zfNuyzNKajfYg2qOgZ5+hXSg96jg1xbLnPEuX4sEtxlxRfAhcjxb3w6o1wXE
sFftZgs355Oboer8UPDGHjJtTXK2JsSPft9ANyRhOwm89FfmDNJAlkypcO2b
6eYu2w0/mJnXEdEp+Uhrn2wNESa692HVUTR3RLAJU1mfibCGvsRkvPIMdAul
6uhlTb2eUmJOjnhvV57NtZ20YfWFR+rE4ETbEWValdbS28tuvoFcAJu0SxQT
nzuCvQgPgw7SYKVeT+Dmgvfj1bjDkvgDgP9qPTOfDgC4Vh4CC5kZ8OexSDzz
hH6wDTqsOAuUW43onaXohw/j3gLgWYlMoNWtXvsHtqfXayTSLKia3eP6+nBT
KDhyMcSRsO8dlI31Z9aPqNMvxQvKdttvAi8cui9VN20wpAM1XYm6KMK9NSSG
tDWT06zbeQ3ArCnzKiUTmJNDzZayPXODyUSwGWYPgTTkri3Je0g6QXOn4P5K
L2y/57WOk43T41/dUxOuh2U8qVTkPj5Ftm95ZCTg8BptHCUOePQ7k9bTR7Sh
vmViSjXXaePIGbtKblNb8tJ/n7hnmK+8GhIN1rjnRM02+Wof8pZ8OkSs3srf
68iYbqnlgZRXMaSokXOScZemGAsYIOjWpQN7OstCOGJMZHPglMjvqbK+dNKB
EaMvCkNBW2iF5wbsPmYhKEQXFqXuh/GKmkpQEMQWdw5FH3Vpw8s6P2WZiHXd
hiKnLDhKFWIdRNp6dUzP8o5n3uckuFKxZq4ckWdlIY84z3XP1k1zPWysCHcx
Oh5uVZqqT80A/qQ9Po9dSkasF6HqSsbdAjgplGRTt5DXa/Xda69b/tfaYbIh
kXtpDZ3zEBnPTvDu7B+t89T2QUV38VEvWnWnmKFd/lxQlYOusj4+ruBNTfgD
hkWeWuCfIObJRkDpHA4tYJylovx6BdSVfX5lV++uR77/RV7I6YkeADVTUZZB
ACIHKOvuc1hhHFNEHD2Rdb8yWZzb+ONti+3ZzKAhoZG+FtMkh73QX3WkElvn
2IP6xUDC40+XuykpAWCZAMt9B6IdBY6TDQNwUEXQ3sv1TyS+3Nu8ih3CqvaV
FVIh5Bm/WRGF28IEDMM5FAUDCOtNX76nVIk4P6JiXLgd+amHBJHV0K966Y2M
k8uRP2y5SufxdbJ/AX9PhHWncZjj07M+2gv6BrK68HiYkc3wdf4vipwDXs0m
K59yznoan1plxqnvS3kyGKL+bAtWrBITCnq8O97TRp16cNInS9KQCKynSdBi
eafXZSrfEVUCkgWB8Y3TR+AjrFcj06tKB5F0KOZ/aFbffc5t9yXEL+QsYNH3
UeIZCVVvDCZM2nHq9cReJCwxBTCIRpHCwxkin8mc03bCmaVIe5ew1P7ierXF
tRP+JnvvGoOoiJglunpTuhg2RzFLz1f8mheNfHhj0z1H9NHxxPMDTkUj/s9v
XpQsm3RT8HAz95sUCj00OB7Fhjqr2FdUVkBzix8t40ynY26P67aCzj1P3/nv
qJEMh2Ml/JHSlSMAKhEmnp5hhGqgRiO7Os/ds/sh//zPHvHy/RMiNEiCdlzm
FiOIWwYCueyB5yCYLm0BDjrsg9KTql7ty0c83vyDCMWxogMIZSxiRW/nAdLK
BfImKxaw00Wi0OLFcOj5lKGv0geccfshXsNi98kQ85ykv8Eyj3CKn8sLzxTi
MqF6iVzfesV7oyM5sGFNU+TvINfEg4TPMNRHbCbjMSiScWqfKlvKKHA5bDKd
oJ8AXciOWxrel8GifvI8fstUIIk8Kyts+Z3Q2CzfnWpfnYwmQHC1XER+DIYp
KIezcQb5wLfQQ/hdPpPKspDzB9W4P4rloF0BevEvf/nSTXyXuFQhkISdtd9/
yhWoCKWsSwdNawPDDeuCM9rAbvvD32cYZh+4IeiihO7XHe8moh9cKYq/CRpr
g2qs7/qTiaLGEe0mUdXeKCDXfCFVn/QMB+tNkFIjqVvysIw86cyqCEHqxAEG
qPPrI7v2M2lIWOPtdrN5FDrXPOT56HUgGrGqOEpIRRIGzjhhWKDmRsR1v1cH
brQwQosTInGwb/72mNBT3qUtADJsA7uo8EuAx3k1+vzv70sA+kzqQtogUGfL
cE/C6W8kSyJb9SVy+3ZY7pYTtwt0SsLWO8tdkn/iS/AEXu5obH0RpRy/U/7h
H4WUvvBvCxGsLto8tyRJb6UZDLTfyyVTqsVMr2E2HrjWXMvQuET/P4QUju8X
+6MPJVHr94jTPWMX+kl2UP1DmX1hb2MVcgkF7MWoqXRlP7LUsJmq7sO9z86w
QQ+Bi81ZRtbhbTKQDtHgXDkAM7Ig0CvuVI9uDAT34+ucodCp1kiJ7SGvMufk
U2/zkyUY3tUkB/F4DsUpJbVvzEuS3sU/CYibotTjh+ku21uZO9Dl36FBJwRx
XVD2q7Cz+jWaKUQAp7/QXN83o7uIQnyc+hFPtYCsRcm1ZxteEbdHMNCqxJsI
aFXRUmFQNZ3hFyDrIB/CFdg6KsgWeV8MrUpkIuD8rvk7GjsgXm7gQn30Aots
wgpUKlBT62PzCK2WLJ9scViSe+qW5UaUgCoaUXFSCK7QnzWUTl4l8Bk5OZoL
Q1UwBXDs+JdTp7IIrp2ZcxGpvDlvPI8y2i0TslHPD3V+VJgPgfVLOrdlJWwp
eCF4QZIF7Qd3BhpVFloYXXgs9WAZam3tUqjn6laQrb3b8RJgtEicpq6MH1UV
GlayjF706iQiKIqlkvDlXn4IX95zv8lj83msEPJd652jCMtgFYre0ROWSB/B
Y0lBZh6GFw736VIFiKcftlHgP92NyqmQ15blsOclXQWpOJ/us664+vtdr5C+
EHcB+trhM9AftM8xDN53QNliu4KCI3wjDnLvLuyGyJvowttVLqQpGADRaHw7
t8H63UfMNxUJ0o88eGge/1g9ka20eQ672irgGLvWmxrQYpImBFvXQjVunw8+
YLBTBYupJnmWDPdrkE7vcoyRcf7CYfk3zmVwjKu2OUcNwjLzMh9EOZaJXDku
0NZUhL7yM5mEIQQy2QMAQ4tg2W+YOuaQSaIeXfG5zfB9ufOHpf1+EHv4l3y+
Y4ombbIgcP1Z9ffMIEq2WzUXT0V3UiR2RZe/oYSV9oVSe6Rr6xP4ySZpAIA8
qCJUBFMscD7S+R5IADp1+tmGHKlCuWulWw/Bx4+P2BuoZ5XMbqLTPxExp+/V
nbnJc5N4f8FemmKkaf+4wzwhGIfp6qghCGjAS3QVZ/bJ9SERIt4iDfKjJu2R
b39uXYsqOfUqWxukFSyF4eknnoA/dBwLWVSkswQ2f00txBXDqvGHFRHvCr24
xOlo3eHVYAgza5N74RVeSy4yqTbOLGpsFxqBEda34kos4hosKHV3E5eKXzAI
JGWQp7mFlq+e5KkwK3/ZFhs0ygmgs4TzCo9AZi/bxkUhbfSuPZqbixZ76mLx
t1zzGbIlj/95BIfDesxdA3918x3OCoYs1vnA/ajl1itCAYEdoCiHgyuOaVF0
2+bVxhblv9wltxoi+HtmpnTEsqROMehTi3hmJaPbemXLXQKYyyujmNHpMPjK
mhj7h/6YWv1HCGHVMgv4QoddlqxmXbosmAqUvK0aby0x2OHUfCEHbJZ0fTL1
XGMpz37ftEs0F2waNZCmuEoqsrzyYyH3Gr2VsvyXXOJQ99wT1syCMFvQHd15
oIlZDsaXIadcoehuUOHxjvzp2Yrtm1OoQzpDts48ouK0EdItH/gnPAYI8S7F
cN5eyrJZp5Z7OgMaIRfLqSqRntzdXDbFHdIEDnILrholKb0dvdKil191ZaF0
/KsIh2z/anLTpMdep0zGogdY1MPrpgMpIb+qwh0WekeB80/hezBNLSaTL8SA
VPGeTYJfKPNt5SDhA/ud1JzNCClRSyuvQshEaU2sLAeT2rY/D62CPl7WTNTY
b1/1cQ20no9nL4Ek+MRbC5ezA4oWlVAhJWenT7DSTEvYX7Y0u/6RwCcWd4+X
b7YG8ITSPSoLAZbzzFwEUsVjy+IJmKBoqIg84SyJYgGh+lHoD7EtRIiL5m7U
2Iv72/gJH87mDKtHixSKBE0wIZVtfqsusp0iFmVLt2e7RSjnfI7DDkpF7Pz8
sJbAJTyXTumERhlsreTNELvLQhWIxJ0gEzERZHLpQDpffQPN/hy+I6aBD+FF
QzCo0+TaByVBGKQQQULRc2xftW+lx2RXle/ifMZrpGbbhSfBwqNCNyQxRtcK
DvOiDuT22O743/wSfq3DBsbM5eNgU9d3v0eEuENZ+9St4CEDR1gJTzEwdvl+
FO6aBAP5+4YSR0xlJENpmzYy1/qbO3BKu/SB6/gEcC7GeZoUMDJ/cekm9dIp
HdImzjBD6mBe1Vu4TlnCbiC/W6Uu8sRqEAZeCVX9YMs7MtuO42dk1YgJXZFo
f8+XO97krqRwUF+22UPCDZ4GzcKB/Uy7tIKwrYc5piJFJuXINE78jXfbVjeS
9CABYI6xm24uiaRle0WO5sqLeGJA8RJuae6rWb2jBlTP1FbPRMzi+tTnwk3K
RrhyfEoNXGRCEE/4vbED+onxAk1sVWu4+j05xQZER+XRcECWynxmpei/liex
mCNWtfJJ96fwl8M8Kd67zTqdXl276zvpD4719sOALIVXNY5bHYYYkXMLNp4r
Y0ZLss+kAhRwdc4H2kRxoQNgPhtTg3rkYKEgiCLMR53XY8heTJI3ZeBLUeNZ
mMGWl8e+sVbYNztg3zKXmsBI3UqqRUU4JE1ZRJrsEwj5ncc4C4VgJDKDQVZ+
Xe3veYaadwy1UPF/f9obFXzC5fOSgZaXjcD3skNBWI4/17hD/H//SkepcDWz
qtd0BgriZSeT0pgJShJco4bIy2E1NIN7EeN+O1+GEdC2+9r69WbjjcFzmM1S
vlJfyaJYgRqWQcPr18kdOZ8KxIjmDl96Mv5eMU90ZSs0j6Ao7TK95suJZ0Ns
7Gnt++wT3GtnB7GLGPRLUoJ66HGeZlz0iIaPsHlwG90WNG7Af6wb30g1y+TO
8yIaxBZFrQSlHo3HZLnh6Fi+0HQImnErC1YTayjJ8iYhfYHh/+2WoG5VB0dN
aFnytlTibiv7QFrZRDyfDq6URablOiDdMfHdCM3xT8ABkDCJ8Wid3N3ARqdY
bnc76ECUMRPWKYj9DZMOxTjpkfj32gGE7T++c2hF/oWMsCLdW8AtKW3jkYE6
sYO2BJH8apNTpKWw1qL0juIRdURHzcr7WADcN/2YMV08Uoaxj4Q0bHa2DLsM
TwSloZW15gfUdxNMtFeoU8f7dukHrafMTE21UkauVYGY7lhqXS5toBasxrOw
6DHDL3uZJ2QoiL6R8lkDNgW2ospIYpH2uKT+n2TlBzheUzV+tcW9pekVjPEl
gRhYB7Gg1mwJEZrzvHGATZ/zA4rVK7ZmeJaBwLIGrSl4knpHcAsyP/9jiVcD
Iwb+ulYS5rrIn37cMJCCGqAY9v6KhEe3zzLxgWDXVvuUYqLsdgHLP0utEuuX
9Gy10zhGEWQLpbspJf8E7BMGEhqnhftlxBDvbXQyr71z5rzRX43X4TGAqIth
fo9sbFu//wQmj3xde+UbYY/qStrSmB0Dcq1cwtg4wizWtw+GthP9V9CakZjg
Xg4hBCdRnB9Q1ftmhEEGryuBWNCtk/zzxT5RmRgZ+9fXkjkBRK/fGcpOv51F
CeZzR1h5+mNynmtDJ+B7F60R5cAvmd+jKSGeGDcNcDkEBfJa5WUSwkkqvw9b
/51S9phCsspbQ4S4/w26Jr///nGyPB3QTusHqk/90lmLcvaEQYkxq4vt7TVi
vavjODR9/pjXsNUz9nb8tuP75u8bxRxxxB/lWhBdMGKXYbJjKoIxRmko7oFT
j8G+A7+CADtHpjO6EW7XW7yzBh51vF4DvO12ALDysrkp7VY9w7wk1BgKe9LO
lsO0fU1tzqzAop1cXdV0alSISxXeNVP4SBbFGFJ1u6iDhIHeYPZMnE3DMetM
nD4f/whXi5pos49puOkTdU9A29QjdIeqNcxDuwGnR9BU8zhBVTiaCyawCWbC
oDxmrPb+CLWHI5+XFmSnzeI3RJE7fzLgi4tuAxCsMvpnQogaMKMzTx03EAVa
zzIUK9XndRJn5QmZnjAJaTnbgdQRXc4564X3Dx9+SIlNqyLPJFtCm18DUctJ
FmzJiR4S1lo1+fXuPrbYkEp17Iq/P2scOVIaQketFn3na4vmtzRNTV8MSzu7
xFTCWobMAN/rE0LatOOfJxm+Iu4wRMhuGXryeNrwsHy4Xa36+o5reGwS/jos
pO15l3q4XlN08IiBPP7V3T9sjqLpQ0A8t1Q1/QmHbbtKlfFoC0Opkv7mfTjT
RrJabn2C6RTt3X5HMQoFJiw0nsNsheBg2vkE8jaUVKh9eNkzxXosraDDBbL7
xUlzTtAfbHGhmAPwXT5Qqs+hrdKZK6DrWWhMqqSvjBt4iA0898CxfbgTeZRj
k4aJiwPalcE2h3kUNEUI/5kJjZjrLVBVvra+xqveNANKPo4CTwU93Tuqfb/H
WOmAw+50e/fIrECPPN/kSlzywWsMI9A5g0bSEer+I+JcqHqN+Vr3/DYS7CQR
0jTtzTq5jVl5QJZDLIcaPAvSxzpIE33rX/r0w+08A5Uf4wH6NABKoo4rnQia
zGXJX55oaAFCRRmryVrNxK3dPa8MCMIJ/DKhIvaNlM8oEDUjwse3WKwUQhMM
KzdQxn9iz+lg5Am+VtR7F7NGsuQDUZqVyTBqSsgi0PLoFADOxf3dvttnceW4
uOBfn8FQ2+7JEwypM191p/ub3E3fFvkU7bGcmGmOUXUOpdxidUJATWtuc+UY
CCrZljaWudt4pq5w2x8xEUhqX+fXwrtzvl0YgV8hpmjKQAok6qsd8A8ki/wL
1BvfhxP2vucxJRRLBtRoziyym2KbijPY4nr72ousAG1j+gDz+pG0p6eWRbjI
BPa2j+TnijLpK1LBv3z9ZSt9PRJIjdQi3hYMUIMYpqN0nlQMziWpC0urpKRr
mBkMM3BCnVXqC4OttON9by3t5yN6+F1h7MphLJ8JnmwCTarGGzL6QgNkowuO
EOSSSNH6bpC5C/iO1o/PKrPqCXbm/wCmxncLJHkwjt8hCJsAOlz5boT2/LeE
9mEV9ozDZNJgGO4oL/Av7TSc/Hsttld1ffGMAXJmcBOGsU7h3umeXw0L3fPA
2Z37JmVRsI5oZx6OEDZQ74ERSKNF6wKWLesimDs508gc3047whPmNwrHQF0U
ZgJ24sOXS9boBSRiX3+nhJ6MrCiIxU0UrCY9hwbMk0lDubDBVsBRQdDICkaB
Vht+OUgNJvUGZFMucCg1IQSbEJhiymPpPKrW0lYmB8foA44MVI25EKliwJM7
lnpE/4kQw9PQQt8Nfxg4ioOcYkT1zQZrDjj5rVuI5i46eqKWaB3Nhv85ypdR
dGODD5EKR1pNrJZ2k3fRjqcNxd8dGaLSuMsSeFBpwmXkI7XQEABM3KcHkvTu
pMv0dRDoabYaej8aKhwIBDDdnIjBcxdbuCfrW2XDqVzxNaekzFP+ijNSf4bS
PhALaBwxLG2mX/gCxcLvTT4Tb0gDQCKLI/vTkyMWCB/sU0KyqdJKWM5sCw6N
czOOdLw3kSsISVxzmQ6+P5z/Onbp39Gt2BpmIPxWWEvBDEoy03EkfBEiDFn7
4lRCIHPEJKYuGbxSRK1jripngkAX56AO5doRRLaTrJq/Fa/Op7FMvpdtfFwJ
K5FJlHnsILoPwchUaJVAaktRN1hlRxeC9nTpEiH/zvbEHnr3EayUDqMb6Z1u
BMki+PB6BZ8db84DP2LxVgsYqGi47oaXifTMTD3+9j4s1Lm+y/rH66dGjVsf
6cETAOa2S0jAfkgqzMfLiRULXUmhLs/cBnLnFfn+hw02IwYDqCSe8QONi4j+
s1eE16fCFE04QbnLMtLXVZeO8GitF8VGUVlZrrF7ZDZf/0QqXxhS8VtEcpu1
xD+RWscHMBC0KPaDDyfufM4LDExj1toYEEhh+RTCqH/KkeDB9tdQ3KheX604
xQm6DviapfmiiMu5es0DCBN4awyl/boUU9Z+5xOojkivQVQzKTqc6vfEqEW1
AZczgdA3KypmllZsPVyUGeQxTCiQ7ZbRItkHtjbCwrmSzNWdYQf8eiKZq3eK
cKiOX8mGN2jw+q/bJXHabOecu4PeK024+B/kxwoDne5hLRpVrhT5leFe4gvp
4/gFq4Ud6cIKKIMUtM6oDL8wJF7G5MrdOpkAOnhdHmwLLCl+NK+aRbtWwDYh
3Of8ixDTPTiL9tEjO/NPI4NR8szu2UXteVZlF1SW3CydcIdm2ET5iSqVrdKH
Xzw697Oo8MNjug0G7hIEf2O0qEEA97ZqRf0X8BNQSYJz3xqYJ4376tog3gZI
o19j4suGSTnupqg7xCYPtZVfP5KsU48uPOIgVmS1QABA7K1PibDpAjvRnfY5
Rc2kzR+VKutp67gCLw5DtBlS+lC71rBAh7lhnRcFKiJ+NBKrR5CoDiINMeBG
Q1GZnve3D5WJHhPprOSc/nS6NaaCErJLcUEQT88bDwdlfVGlsukpQerbXu9Q
A6GcCkb0a7e6d2DoQ1oTRysQv88ZhbfaLcDsztgqmT5oH+XTDc0uvjRtNCTz
xlF+euZ3pZwzV7Nk/WcCR2RoOPdNvT4Lf4nUWS411panfedhHt/alNuxCJRn
RsZBfmvtINQ4guTZKE99bBNd+ffZxKlYM81E0ptAQjUt4F2XuWkwu3Mn7Qgs
3c48Wo//6gPfK0PA/lcxW8mZ1vwKpfbd2QR6IWtZd/uIRKJ+BvdUM9uIX6Tm
/Io42TkMxagOjhiHgIzH++0vp6zXbwJUEI3XbqyX7MEQOZOwYPNUuB58xCmx
Oj59ylwyPKaKtowBEgPGCEouawaDLRU4XEpiIIv8QYJAcj3Fk0x6FD7XmgTT
Vdo+IJDWDk1VdxabLMXfsc3FJoztKUPQ0U/oFQZGh8V5MpSWWrGMLzuIiXpD
SdkxKsKGgzw/RLBm8AhI9ZWK2n/9o58ENKtScdbs6y+bCoX32QiFjxrRNqo0
ArJXbK3BGKOZ9vMa/OlVjPBnKGqOHMG3a3leAdfJsrfFZcL/m1NptB5LL/dU
Ab1rduV0+lqoIrq/kzEUwjB2sLMiR0iQJvBZicClhlqnZZcNgBIGmNM20pt4
aJyg1cYCjrYgd1QoLEuJo1xxA2q7QbJDO+8YAd7hltChShqEztP+vmoZYvqJ
srw4a7+8VCloEy9k2jRbx/ILuLaiz+bzpPxi3f/koaif+WOeZO+J2Tjir49U
hr3AiYZKVfZikBQ3p3ortx+IJ4/J66s/KghpUj93tD4gmFLueXCzQGdLgK5q
uuG7kcCfJize9djJLP9A3eO2wAT7A8ClWHmy2akqfwBkio/uEENBIV2eSMel
y9P895rWyAcqkqBzTS+waVvrAw3+4p19A7McLW1eHvjzE0aW8AoT7wQQ7tJY
aTKQPWT0xfljsxojxBaFBr8TXFFUz4RfK+rr+D5ReMHLTrEyTxv4y/ta35Do
UOdLJYUfRLXz1OJ5hypFP2gIj+LGeDh1axigs4s4TMNf7alo8BbOzXmADIbI
sboj+lyALfQBdShSgJxz0tEXNGEVKDMImdliceUdnanE2IOInib4p/Mv6vBM
fQZuvuc4r2fZkO3+FTbCT9DP6toGQcdU8ZyhqTG3EIbvwvWBTc6T02B9qtcA
zRyJX43W+riGOpsXHTfVfFwOtFlwqWXOuOrXoykNQS2tdXbTe7bHNVJUMb9J
USbeEN3aCFWokGxbJDwVkFVRdhvjne2LJ/2FsCKu0TU9Rq5IJpLhd+S2M4C+
vk9NvulzglrPOYk5GDgffphWkrytWNRQVPL2unOG792P6Ls/LPc4kYr/yi74
WGqjw7CzVy9Xtz6Tjr3WsWmfqlP+YzOycsy6jpC+e+7iUEjYrU7ZVAtwy7tT
lup+qKXD9lUYQSDwMp7Krn3+hj8tvKCpPeYSOU7Qe0OTINL7t2e3Lf/chIlp
S1gpJGfpB0WjvgdDLK4exc+EkuS81npLGrcVHX1u3Jb9WgoAEarhpDgnVYHi
utF3DLEyyk+aP44nLucJHANIIVXFERNPN65bQD+hjNTgaIqY89Jnw5E5+/NQ
VMClLs6aNHOCeTZZa1KRxh3sdSEOfFjtMEnvM4dlky2CWd9WPJwpXR5lxEd+
fzygc6XC+88audTvgFIGEZlKTBh6QN0DEd4zoDpBO86kOueG48AhyZkUJHga
sFzpjCTMoRoEoLf/qt4nJ2iqOee16f8nfQByHRAKsEvXrgcYuWlVyHgHhskR
N8ZyiycTXOZgdeb83D30gE7/1Sx8Xjy9UzB0cm/zLxxXGHSMZBLI4VVVVQ2y
wCjSYxhnSgLg9blYea+hZe0wiqDxGUk+yhFIuDkFOz/xcoYNlp3RqFnlHjcP
K6hLwpOYoyzpB1tEGAEYHSdyC8Td9A1LbxxD8HHyQbcR7tMQ4Ni4Mj4uNB9u
OK3E3vqBTFf2+jzd4fIxoJLnrncj6b4/+7ZriQ/iltKdcy88YBlQGC5QCf1J
n72iko+hnuZUKzP6KUjVYEwesh24heAJpbU7xNqs7dLxmB3rWGiF8lLOrrTb
iBUwsv1lrk5aiQeXp380gOXkU66B/42YmjAtjdX67Dk03VlRChWM5FfOdAy3
fWWkQgjUvrG013jAP8mV4occFc5bWnbF1ArVSJ5dUvvIkBpPyghaMsp8wOUj
ZRBLb/mYnBmKEQj/BdugP2zG+mZg7Z2e7jKk+hd84YeSGu3XUMb/GUNATeBC
Z13jg93uTkpXmnXr4VQ6ztvm+6/XRvChBvvU7F/tit1cLdSiZH1UZrUonE+b
szY+lFTkJAjQTcS2UcWHJhi5nrS722W70O50/86B3+qabMWCK2FENWtyyKmp
0HI3vOj6kPLDlnFLb2DLeC+AeS1Fz0J4j7u9ZHQUNeS1dKVXVsTKsiwLYFUl
HShRMNtxPXdhbKTe3YxMER3Z0WWeJeaUb1JIgKO+GTji5WVAsJTcfkGvqy3b
feOpPHr/Er8pcQnCAv1T6qvlUMbdd7PKC3dBGNPWbxmp04siEx7OnnUoPVao
qN3N3hD8oUBngTq5+4xVr3SsRRuWNnSPvBzZXdFZiTmFR+i2a5LRoIr6pxlE
pdKcDwdt4vWod5B7TDg/h6P5uOkyvfr0KZBtVdFN80ZWU2cxrg2EUQuQi5Xq
O0pF0g2rsMhSqJGNgqDNv5RCtGdUEKtI/Z1MkHuLUdOh5OPLGkEJ9DFCzzJz
w0yuQevnziAc/8Z8OVHZptkNVAn6q39N7pxXLXYaot7GkQwrDA8+MCPvYsNf
NxQHuL15Xd4eimW+LJy6zhQvGyabm98uqR/t06qdoINRvd80QqrGvr8H4iOp
Tb2cMVtYFDldwNECxxqrxyDJaYNa5dYBH3cjluhwm8WVOZQwc1O/wYPgWIzI
hXkhqoimHYqJBTLS2HsbZE7hHQ9ZzqHWLGBy3o827ZW5GqpyDyrYImUCtybj
Fgb8mAMkMTdt3+y0CGjY3Dc8rZK7urjoasyS+OypbKj5nMM5tIxlwAN1wmmm
rmk4ae0Jug4e4m0Lf4M4XlgmBOih1ImmBTe3KQd0KWyEpxCC7hYfl8jHeXTS
Y0occDnWfIfnBw9rpcqyf/8n5NheIZ0B35i6U4S9V4JQJyYJ0y94ohVe0gwR
tM0cA9K7H6lpncxVhCtewnDn0HS0+SAv41vErjdv3jrNSWLL8CW4wKxm2Ii3
Z2Js4yf3pankyRfww9DaQM9v/PqpExwNF2id/P1PhNz4+nFM1Fj5PgKYQYDL
BNUrtMj056bbSI8vntvd32bkTmUZdNDftGMwAa5gHbYmKWuiiyPgNn+HoHWj
1YkMiDUEMlViGpaKybuOBcdsWYaNWSHF4AV1SbUpAfmyb/vued+wK68bz7PD
F1b+Cxsg+O8nYKJi6e95rd23h33qNr/YWnY1TYpajBmwShKGid2TcKz4eYA8
fyYDQEMfUx1/WynOhe45FtXWWUcUozkgy5YQItr0ScBZIwLB4MjZAx6Y8BJn
TDL/FOgC2z5mnJ6xCY6y/Khb8P7QDUZw2wsEwvQOIkG+OeajbwToc77EEXCF
knU8+NoWjqa6lpcpWPryawUZ8ZgV2WyvXeH8mCwLiIdylJrdXliXs7+NPKrs
pSW+m1qJzO/SMv9iAHy8UwliGSqROqXP1linFBidXH9BvBJ1IrvDdcm6/nv5
xyx9DKeTc+QTR6OwSgqJq+NAT9VbnIOv0VISE9EYemKfo+BWL7PUt5Hry24R
J2Vi+gxnBCX4/2/67eG7IRrJMjrspEwVl4HoA195dFa3EXx4I6Ho3hTdZcjT
qakCNpmY2uOHvpj/WHhNF6OZ/ioqqDSjXdLgYyCfM6oFVhxQgKEP2TfoGX6p
dD7PAic9+sqHNwGmwcJKh/QumQJ/nwNvA6OdwJWzgpyh60HVySBsns7crQu9
Bt8zU46vb4frVj0cMvYOzzWxBcC56+H9lxi4h/BqQA4D6Dj9WImSoK7p+/E4
cnZAkXS7NCFT6nJTJyOH1Gqbv6q5nbc9QDyTM4rQRB/38rSkgTYMnYqr4sG0
oUmArsPA5So2ZoGR8WDmoDTMVFY/pEv4+0defaPtaxdL9jJW1/i9rO7oFZqM
BLliryFh9AzDLEtRQku/ch7OWrW1Y+pXwfxIvzQTfSGY80rwvIX/EQAY8IPb
cAlpibWtycoAN3WYjZorTjSudNANkplizZ3IZRuJxjP1HtCG6zX4ufbW3x4R
Aa8+m57cCyokoElNoot7WLPgHpwvhsurccKfS4g6DgTkJmtr7RGzdVFycdDU
jH4RRpHsfBXkVIOZX0ZiyuKA7VRYPzkAvRoZA9eogvZ1yngPJicFVXc4FIFv
nH6PPmcn/r4bzVl31DQRpes18spBR/Fedxrq/zUi+30GQr5da7zFTGUMaMQ3
Cka5VWGRliTO61EDP4OTS6KFwOFe0MAezxwAU2Lrq0PWvzLHNWJOQpzaZgbK
B1edK/URqH+md1eL81XvZA2gLJrUPc3q3Hl9gVhm+DVS3YgZw2KCGuR7ShL6
069WDAql/lZRe0Tf+ZR3QOmJKNBsjao/rIxUYZzYastYSJLVlTv6QHlJ9xWO
iQYNdDgtdrYlFMEyL0asK3C9T26r1JQixhCkiq0osVLHrz85coQ8RDhRpiF/
D/VkPFyvBR04EXTodyvkt9BK42jqE8iAJCnnbfVIFdVxT4aDwoCUsOOvEzMA
oskiEOdgrHJPTFwhYE2S1E1w7lO1IP/gvH3F4Deq3fQlyvMFdjkZwMTgGEl0
RWN/QBGYTMMBnS1BMbQ1r5WgGg5unLnGxtgXnCnbUeYjGPQGToLCY1qsv9Z8
0HpDlDQ2X9DfZh+2XVvKGXf2CtLiaMWtu9fU0NQ6P26QBWaKqUfLnhtySFqb
n1KBqjx8gwwuRog0jT/w8QuSIV4WZzeBSRSZ19ToWpT52sSGZrpc2EVnsv0O
KOFBImMzgv9tb5LIzOyubJta53IuMttyvNzgBPeoL3Z1nfLP7lofI7wt/z5F
5T+PvzGmv7tMGqGSRdFl5OIUQT3YGH/sfquFzAUnB072cF5mGIz5Wz4foxAY
Teq7QfWViWdwJ+OSYZmSA5ksuWf+BHJ4BqbaRNWPX1Kdf5MGXeqPw9zwFrK3
idth4e2Y3KaYe1ysvTwolxBQ+lZTPICHEuMCbnSpAY0UU9w+h0qG8ESGlY4W
jvJofSJ/gs5ucpIPByGZa/7OfF/fuod81rwx0metdCIUeYwYRuO1e78o6IkP
HgJ4bthzJ7wyvmjZWU1N3lBqSOtbFO1wxpKOhg0bJFrj/Xr7RGI9NDOGsKil
ogVBNm4nmSE5hkbdDjs45tMkmcOUjtXhMIlW071imYrzpbbY34LoPziQLhKL
tJwuwE/SvbKSy7/5mTu2yC8tSWcyPamzhA8fmovuTM4tfS1KUHKG3ZZM+uUX
3Oh4I12NW55Ah0Ayv+PWs8yIV8PqGlVNB7xGmu5BxpnM/8ZHv4O+4WcpQRqy
4EFkSMfKZPGGVjLrbYvr9AleUHrCS72h7Iw3uS9vvs/oiyl5bLA59mctsGbO
q2rFMZH1lpK7g6Xrw9YAUnyuULkQQ+eyL+4euwPt6JudW0Qwx0GA/T8sqWGu
d2A1DPHJHKY9yeSJpSswQ4Bvq46gRBxzTFPRf/b+g/URQWz5by+9F4uaD6CN
+njKrZWxo9hSL9c05Q91Ow2aKjf5z+i4lhwz+u3nRrqtNt2LmGDZUgntf8Ni
15zk8gdKnbYXt8ZUfLw6Zjp7JPyBeuG4RWp6zD6U8wT9ZaInlD0oodQk5MCf
vK67Ee5PPWptHKrWnEPNmDJ1OpWwFPM6urECqKhbuWIqeF3KLHYD7gdE4QH6
8y0maSV5WEgCwP1mXkydjyodjeJnC04B58DGquV5otfUzk6wOPUIpW5wi3Cz
taoW0yBTKKDMO7CbeYWbqgAgNCiJmJhge/nbngWrCr3uteRgUYEaxQ9nzVn7
7fsh/NCD73LEYA6KTiPj976kvdaDLA4VDvUVIg8VHtzcc+A5fXBaihQvmPO8
zKokhxkLIifx7EG4L8HSFoS6I1BIo4Co7hS6DIoDZW+7pVRI7/YXA1Dwxd89
B/nsEIbdUm3fwlliEoUga/4hZ5iXuUAJ+a+ZudNZxSqkD2RRArQ+3oyUtF/V
hSr5mBkkApvwD9h3uohCtB069aIk6q6e6mq4AmMPBbViZISFR1qusd2KacVy
Ig74apMKUOOIpQQayGZxb7rAw/NCzuuxdQ6w3wd7EGovrV1dniRvg8gwCsY/
lbpUfwRa2FtM4okquWwUWh5VkHDex/ssNYELZmXTdNLdv57V5m0n3ZUvr88y
qc2+Zv5HpvhWcRbjU13DoKcgzc+At8bQaZOHwGlB+4amkz03YaWQmer4GQkj
o8NHvEuJkBZrgeMir6c9rgmzJBT2WgqB0Oz/lahZGFeyCvM3IjxXeI2ZtjRq
2mpRPQAnIwizTcFtQAoUTdXVEsu8V7GglEewwMB58Sxs72eFyCK/EvpJ4cXu
3KAx+5haNPZ78woLH7vEUXlsjQEicnmIqRTLiKfQoOIp/IiygsU+ZwuhTHhy
kq6uHNX2XRBIi8J1aQ5H5IrA2VbkS/Ljo/Xb7ezmVAF1BFGmOfOWUf1tVFsH
B3BKp3G+prYIDtOg6ysqFgrAMYx3D9GTu0PgEsN3CBYi1myxs+caIWh+Zdc3
1Cudqegme2w9ffhRoWA842ytaXbbGCv10egpljDSfg1SD5Uy2NEuWks5geE/
fCmohdFL99NwBdgrtSEsGwYCBnYAEopC1CCnUQDsyHajQ4fHMpuUe9qHzkRn
l6T+LoCCUe04agnA3F7Br2RZct2RT9poZecWRZEfQfcq9Ub56Ay7XaxHliQi
Y3ms2h2EUjyQni28NLy0ASG4fryW22cGuRaRvrLSav6m4AkhE0m7kR/B5kf7
3C+yIeqNHQIe3EEMiQT6CdVv6m+dxjvsoh0oWMroTxx+bX3w6Zar96UeITo1
AM80RKKB5sBM7YhS6ZdUKrwSFNVNTua3XCpve9lZnJtmSMZ11ZeiqUxWHlSM
FRBKhmT37ArluWJX6Qg28c0ButQx+OEuCkue0ooWFTCdwgyOAEe7jCWh57nX
mdZ88YpXqoB8j2b9F+5OdwiFOFek3hEbGQLlHbqt2IgDt+t0KWmxOOobXacg
hJCOy7oQjhMDjKRVDjUTdncthCXA/ddDz7BbSQ2r8w1H4J5xKLaImu5z6cgF
miECw0uVMaVEE/05cTfhi+u0JK+zYaN3fP7RT3eQf1Qtmz5yvB40GiqPNClV
vSsX0CSvxmohWo+yZAfokBabdvNzaA0Jk9I1Xjhrs614KkeWScqAh3ziEAAT
JGZzXRtfyZrbxiMPDmMLMlk7xfK1dkG+91K2ST//YyAfOgANork8ToL4U9CR
txHUfXuvlfrxWMqzxbUJnN1SuyYcG60zELtza8ll5ZkKTxAGN9yWYJ2aDcZA
dMMrz3kCfJR6vtnE4Xx9b/dEikdJx1S9+VBfhocY8T/g3AOfYlJZ3ov8lqyB
lFVAAINjYLl8kv6f/HJBi7ABZ0CONwctxwIjChFxdRq3lwpnoccUArQg6EFh
UDrkfBPySdJWsNqsXzvQ5GRpxrj06Aj6w4djkuNIVxdkoF0chdavLvFu8ivm
M4lljKpFnMcRlOttNxt+6vcdtZd4QKswH2SgioVyjcPkwONCJOd56wy3v1yB
YBRSOtDsB914AgOsdtLb05aVA3lfx13lYS4j1SyWfbu13E3ST9UNEFOJjAhN
lJH+XF4Yt+HUMIneqH5P/3+ZY9BsiD21KEmlAqOQPfLehU6JeYhkbCdXP/Ph
BA7vU9yKWsNILxKW49KNeAzFZlI5nfSKwj4t/5YbVtmlTQ4GDY7kS97LNfE9
WzFBFk2foX6U3JwHzeSLjbacdDr+WUThyLtXA1y93vvlwNZYSvUZ4ZQp76uR
/7MdLPpDJrvYruruXTwoVjmn2GaVmAws+2mZZAHYr6UrLz0/siWEC1i3Z5Hc
E0GSiZl81RlnMaJIxndFRAxE0aq7mzAwDgxiUc9nBFpGOkK6zNLBbeaZFZTh
ILUfcAs2XMTQxTjG5Dc1b1kpJcvMO3RzHTBD8Oup/dy4fCRuIgXeyUu3ZJnq
XViwhGngcKht0WSEV+2kz5eLTi6ejJegJ865vdct46Wxc7fxmcyNZVwcsT5l
ZXNgxkzaNaor9hjuuNVt8cHbRIRJgZum9LE/dzCh5BqBlnUbJh71oMMG9lre
aiPX/YQ6dAST9vayN+fgXhpkUKW/pQqtPeUftrCdbh/EGb8zWn/005a+LrPn
flW2lkbbL+OzAhi/7FE340MwxyhLPexlcSDYy1qd/64YEsssDyXipJCO91zv
y4vyUI6cYVg5ylG1JEGzjMBSHupyOKXN6MR0MtArXn3eyaCYqBmYx7SWvG9q
tJVkdErFitl0JSJjjRAcrkA/NOGpyjKd9m+Rr0+4UQV6Rg+bp9J7icnDWdRG
6zpuuu898E6v4zGeyHBG6VyfmblAkmgfyB+CV/qBeG1SjrBQyMjfqb7KtdZb
/P5YxrIxKwuQDMnDwLTgCqchGWFY4UmSC0ZzT8tCxq9ZbAB7tM9gaaws9Lki
DhGfC5qSMD1OYiyO64Bnln6VwBglmi4BvrFRwLKl46NnfEkoGbv4HS9jQ2f4
sPQC+KLfYDUjKwCGldhSkJUK26kKLAE0yW10vMzIARZrL+yLlWUkY0cBlUPw
8zBbGFwgpSPrz6tbMElPwvxWgSb3FvAyfvp/Wm0+XV0S5xbqeyQ/M6UVWew0
8HdzREw0lv+VV/CMh9uqR0YuXOHrACSWAnxlHutfxTri9dmKBNJXLL47O6kf
X7tcJnIoe5QgCns1ZM9TLhHM4SqGg+qIgXeOdyudRac01FYjgIvElzd6fX59
M6/zb8UvkNshN3oSBBH1sKqtvZddyF0aGpTETunWt4Hv92lvGg7HHBzEWv3N
+EiYxco8+VnQ5wSlITRNfQwEbBvMqDGRQRk483vmRKhkaSQJZF0o2rVgnRad
ZKYtQzCVpTDLD7JShIknyL4O8aL9c/IJozc0gOQrdWlzl003JLNhmI2966Gq
y6vPnZfI5rSbNXYM5k9SeH5KXl5P7FSga8+9HqwXg15DFd/SEx5DeJnprhPV
Gfg2PaN1yQmEsmjZnuwtWc+ppLxTjfp0TLd4pmYVkmyQvwMksx8t64Y/UuVy
cholKyawNCvIpLdv6bZI8tyGBCQOulRyrlvQZzef4SMjaNpaJUBezMTIOh4E
Dx3/wxkkhKSJ9vVebjH2PJ0ss9Xj9WE5l3IJwHfZMArSLVR2hDrDYuBI/ZSu
kc9iultuxx2s84gLXsyLbIRjSg66G0EQuu3Tl6yPy/Pzivdb9p37dnb1iytG
pMSRNv/LTKNS0lUQuHDu/yNUG2D52YESZWZu2ICtsIax7q1xcgqo8oHNh2bd
lC8d5DpQKLRqiJH7yoISLEAmnQBeHxD35FePN4tAsbXO0jIrWScHypeVGobI
RL6gGqCmm3h0CQkHmN3wI3dlNxk5+NpYg+PURpoUK7wIx79LaABs5ZTMOG2C
bzGJAGHSmdOBRS9GmDudIi0ClRR+2NmbD9eoRaV8JdPWDOq7u0WixLevHfjY
o0fFAxkC+R9SShqGy0T6De9Ytn2faXUDhuy6sW3jBlviBSdpZ8PmpFxv6Gg0
Ri0314pnsNaHfU6rQOlzMxboUOQcdzTB7wzP8XijVa6YaKm2NB35LjAnq7Ab
f3P8m1h5UgpjK+NT6ZfNYe6EwLnoyQg8g7O6gARdDdGxVJqM/nf1rjqECoZk
COJPRlpyUz232d4O98dPsS80hlxyeut3QtQc3E3fbDX657u4bJEzDZ4xHZGh
3+JYVJwZCaMi1VGqwnIqpXOumVFJV7sGop+oEspC4lQnwUEFRtSYF8cCyN0F
/c1+QNWt4snq4fuYqlsjYX72U0zBH8lzRpJkmiKzzqMmyu2F3zY9HUIb48DS
8TegP9woqVDlabB1MLkVmJGLcIfWXcPUWNrJvdxbRBnCDNKRu9Sohe+qWp4k
aJrSLkfHTolZYvaM7nu13QLuOc5guf6ISSghyMw82m48iFV4BzhtTmpSiPs9
j3C/UdIsdqu2qDiuIM9QM++LnQf4KExLokwX5W4kMjRq4pU9IJECtFwEYK2L
yc2+Y4O/a2W8KNnppzYkNrI6X6fWgprPINvDojexS2HGOknBxmjph1gfC8D1
rHQamE3BlpH2JlNlClxcABd11oqoX2xrygFuIETejT22awoagGJLrKgh4i84
4C9DhwGBOgDdBwde2buRCDsVYON4Ia5JQVA56FopuVyynBciio4vDqj/JODJ
J5kXEzEgqZ1MhCO0SlzWm0XFFygFvIM+3gAYnhg/RlsT6gS3eKfA3nT4i0s0
P69EN7oJaVgjClFgDG8UnqLJAYWy+W5PmgWz67z9+ePdFbpkyUh0x0RiFFWp
5yysRVZ4AYmbLLW9d12J/NKAadTLvyUjyADPo/uFdQBJnvGkUmaMcZ/oYsA3
NT/sUOtrILGA9eGZdatzt1KHxB9PbRsj+9oAjADBzEGEtxk5JXUl/SY/05EQ
SDBFIb+oBljf9WLSFZuFqVfMVjfgy/B/QsdLPQAA0cKZxdyRktZPUP1Ai2t0
8Un8Wsx0WPXNUvACytjXMEn5JC5QT97OcRZ/E4Y4hhAQ4sDzx2Dy98oWLsvK
efFbFz5Pz9kWmhTUDakGH37jiqj9B7UeN9tmQiV2f7thYmlNPe8RAfxAbESh
vKS2hiN65PtDR+WayOtNBrA3CqA2y1ojUhDYXl+NdVSJFQ3JZ73j8ye5n+pO
42M6mb1o/G6KysWmUPcoUVDxDOkpgNBhMHVnq01Vm0aDXAjRxOn5d6Jv3yYl
lmJYFgzUlEMYDVQ7stUzwkk9NJmtlYKUz6JsiAZmnuS3wTzxaJopOYrLGaLn
r7WfWZSVBmQWy1HaP1tnfu9plu7KjpSGDa1KW0Ak9XSSt/+1kuqAQcJLvbCY
GKqHwn1cssDHOplFvp0HZCWM4P4MVBuqsMPT8HiE76BC96afBA7ra/kzmMKY
14Qy/AWqMb+iB6ZRcK2/WvDVaSnjfrlr0p/8rzqUV6WVJpzT73oVAKRVp7FS
UExZxHBRlJLltX8pk2G7qb/8EY+nnev9cA3bhHKgMpxJA/HcQZ2vCwPzEohQ
EjI3KKqpyPlDKQ/UmEZDv2XeQezF2rs7hc3qetn7cfD9clhOziVTcPBQnlK0
o+wvaWn/GEanyXWNT3jsFI7xlnupo0XeR1pMwajLgwhghNBv0Ksftp8SxIy7
OMKShKx/IUgWv3xnZ0yng7WfUQyc6FiY83MUBIEg+W2wpKbiDHdZ/axvFYGX
WmXzgpN4W4yN37jk4T/hQ6O9DZsjim+hNArFPhoo2h2bMOUajQJPI4/mBpWq
s+HslHu1sxhm2aoOcJeODbywEAQW6zwSoRXr+Ee9uAX0+OnSYSyC2jZyY8+Q
AXnTP6bqg2BMT//XQ3565tytFpDZkD/tyLZLQak2C1kvCUVA7q9kYNGdHCIW
k5RClv0jkQfVqUlMuT/nRjMQq8LEJEMHZgrZQE1FKpzVCWtH6KYarNyPR+0B
Rinpb6qKgO4AtKWGghVeyegHqqAUA1TUsyC4Ju9hDxFIvu4EVYWvT06oGFMC
qKbtEDBCijTSR/lSyemJvAuOOzk8+PDWj1EmEjF6Dw+UFdhlhNRVpAR1FOsz
hJepG5HfTgf1c8BwVTGB5/jbrL0qNSVZd6Z7k9ImOQWfpZpzO3+1pKAp+NWJ
c5wJr7/yfY41G5AklYIXPHFy5fJhjStoBiwGqSDQ3F3e6Zt9PymXdQTYws1p
t3B3c+/RgGgtIoSkZNr0jHqkJqbmFN4HRKfeXOEwfCVzyK7OvFsb8jXCWGg3
aK2Sx2gAWvr7+enKGZPhLYd68bJ45BsMKqCK7dG2HCPuDz0iU/5dbiQK+NrR
lvQ3KpM8VL2psDiSuDiCpQfEscw0Y9ysHR1FWCcJ5jFeRhdp7FM1+TZWw/EM
dEpo+vJz7EXUQ3qJC8+tIPBPn1NIzpcDsumR+bbiMF0jAnLUg8tNTBftyLCg
zzEIZxXsKdhax0SWsdajWVBFp9wxDIYzZX5C7xnC2bZwsPry8mot/gmzL4KB
PRma3LXUGFuUoo3rwkaY/ezwJng/DkXbflOkx9MC4+Zhr4NyFiu+C3RN81P7
ivNZkCAOZ3tN2ahMABPTHmyMHML0wTkyMopgsQq7Z+Z57na6GmB2OhiOMDUR
vZ2cP0uD7waaFnFCESOvrokEqr4Sm4Ae+F9kTP+FJRtXXkaN65n2JgJ9tqQm
aSHx+1OJZF+S+9Mizwq83EMmVVaXIGCHKeyJt2Rzu3QqOMXo0+gIqbhXlmH4
AjOX71L471iQtaGULjcN+50ejQ8rRq1I/oTtjgeBs4MjPyK/bVapSelIpbiQ
7wvq813ijlEjFOzgxMABwdizfZfO1xM91BCubQcDmuiJnMQ+8BZbi2i/kgKf
s63Pna32HR2080E0wGZPa+BbF75vvPfNybtEkuoaMminGDl9olzYN7dqEaTH
QVvt9ll/Ekcl38GEDXLdWvuHgKCMhbUqD3r9TYWLjmaE1OuA+DU4CmIaVJGd
EkM8NaRe2+HQyS6UuEJE/qqfEUY9Fp1uz9kaK/G0ic/RiXN2a+JmOk3nneqj
4cT5HJpvD946z1rhuGU2PxHKCLQr/PSPdBXy7Wgm2eJ3j0WQx5qNUctdWJzN
M3SSQJYLxXvwiQQLr6g9u7ClfgbwNKvKYJQSnFcyZ+WLzOu/GJVBCaNN0mBf
SAGyO63fiHJvGWZQ4kXCfjbHn0t6oWQyML3uB8AFRx+n2cNwRoIF9iXgw7Rr
OUmwjMubK01F3Jp1w/5rD+4ZbnGMmbp3YVMQ47vpGFiLT9TbvdhGf/lXvRc8
hUGQT+cPgX4ZOQnZnpMB8eqn9Wb0jgfpltJPIogXrr/ztDxEzLOx1Xdhx6Np
qF+sCe+OP6Q4qx39Qy/W0fE/d8o1jdvV01rTLrCe8i/nhyb/ZHMpmq3/ox5B
PAjNn3Nq+J+yBDIwVaVbWAR1cTUVF9l8sifkIIjAVND8h2uVgmcEupzPOpR/
0+d70hI48xlzWjavmdGzVc91pqS9qeWIJDxyWG2VRZtUe9BhRjzm/2ZISqm/
utewuPXxIz3FctD1t5TH+c24ZozvLvfgxSsPfc46Bl00OTnJ58eqzzVkRfik
UG5hOM7hpRQN1dSX15pFy2UA2rfQRC4ck1XGD9NJDmtHGI+Cy/GFid++g0x8
KgLjc1UIB/qBjMpKUQpX8izhxsZYqV+tJC6hLsRlc42gl8DRZtJ+BOYbqlQC
BZbH7xVAMo7CQ0BpN1XUYYuS/OADY2VSfRR4JbF9dbdWYag8We6QjW/sRCj2
Zg27ityfHDBoEvHRwuK1eGBU/SdvPVhedNMvHcQJLShFFMz/+KSoKAzvfMQ0
WwCPoDD5t0cN+32KfL9hGANQ8GHCqUMvEuFATWjmBibH30uR7uBUtbQRXus5
lKP8uH1hr+Ri+OQ8GnZ0mjJswJ8o/EJPm2w2ADY0uyI7tBxsRQuSE3WPANaN
Wjvo4luO1LVOXSS9jy2N4DIRUgf7GqHHen7pk+oS8XHiy1eIM02VPmg3A31b
4INnjenwwtbXHys2GioU6ZYGEMHe+jNjxjh6DaMFnXfE3l3LKO5ucfFuregg
PBzMMVCOndHpHv3AnYX9Hmr0uFo49nmM4I3cT+b85D998JAkpYtFtdjcuXqE
3zCCVhwar4bH3/k4Ue3pc20p1L7oM+UExGvygJiDpMxCAAGXkLcyz96YLzkI
jbahQMK6nWpv0JlkmPsXwzKRHh8fcHEaYU9ckrA5esVlZ3bAQEruxWL3fYMT
a3oyy4fiMSyYr1iBsRbRrefT137SiYQ45tUR5lzru9q+dRKPwp/0vkc7RTjw
OK5lAymLK5JGotgdsNv/FuP1w8S7LCCLuhxeIaiLe1ujmzoWBzRwKuommJTv
wUl6xvMIpTfa2tf7/WaSjI8kXaAlcshitmReAeBEGC72E4wrU7s4QAtghJG8
m86Kt4BlPKc8Zy1+MhubtRz56ydhRXtycEbuaupnFOd7jaHVFOjMH+S9B2pm
Ijb16daVt5V7TvrVuoLSnI2wnTa4I6BFHyojTGoy/2pCo5kt3sOQ/Z4R8k4W
Fx3+nHsq/Xd5dnliWv9yRmvD7rMT3fmM4XPPev5m+cqiohEzLg/WZFQI9myj
q+8Ketj4fuLIrdfjae7hTjRSch0VOhlriXEUoWrTVa01HimqCobSy+/io4EA
ADXdJ76cX8iTZgTRa62FOSvxb8/h81tpyHvjsdj1xa8Fni5008KWE9/iS9Fu
wVh0agOnAuFeomJkTHi5jEeUPEw9Kh7j+XDrTR2HMVfaOZ1bTesRxC8oAaZg
LhTWKgev+IGCor5P7SSZX5c8wFrthD5ArnYwpLWfHsre7hmjewz1Q3IK0uXa
etQ36Ky6M8JnwPRPGtTyQNRrkV0sxr6KZKQEZRaytDYF0O8Welv4WssMO66k
Nuop7wGgF1JwDhUiPzm1sKc0prFTUpnGmOIUJaAQE1fsLb7GfOkTnKIyR//X
KtVWNnOjZnIAUKUqd+bybnvFQtIYRm5aLKWnrEGvnwvBK5eoo3cRX88+7Km+
HK4t7potgG8pq+yw4t1bn+XvPJY2NkXYDVNfcC82FjOymDzmKtekQtbJ0KZY
wGOg/09INoFcurceMzPheRAO/OcSy9OixECw/XeghfX4i1FfQyEODeCQqtJ1
vpRTtgQMSPwgKOKo6oUGS2O+izAox6ur1RicVy7NLlQhYWFITjCCbeuWaG3X
lFHEjvTgsmU9wYAjMTmYG2KQv3wKU9ES1ln2HPdCE9Rxwuxc45K4+VG9IedD
7HUuE8zRNeoUaBs7PRtNOdLf32ilmXmCWbanKp62A3cXgWsffzO3BCxAGDL1
tXmb72JvqPogELzBGUStsj5CqENyL3IL/aJyVt3GLlBMLxJtVN3Or80XlzVu
tADcRvQkpDTuv1wt1d8KHrgXHS8783QiaE4yRXq0mOxVIKRWrQoQ46Zhvy+H
Qa0irwiVCjJ8reMbkfZSYhcRzwx8MEVT3rjRFroY/G97dsTp9KvNideRsOre
GLYkV2obmJRLw8xYdrXlpf3j+rco88w6rIlRTGu4IZcGaasD3NGhTuMmXL8S
tlA2kcG/ELxKl/1u3B3PtYIqn/EI17xDom51K6Jy1da6r8R6wk/1vOgr5pVH
g/zdRhqtKrYimgBrgpVaVOJnN11V+Hy7CERNaI2yCmpBs4SaCco+9lZ0UFPg
kkLyy4C2WkmJEaJvodtq2PZCwSneNGJIAbP1cJdV/vAuWdvmbMYA08QDnxc/
dOWuzC4Xz7HC1WfQzWYOeSVOzp72Q4YQyULKwGtEE3l7W38Y3RRqN0twuRGq
UJvLZe/bv/HTZiXSccS/fwWACHRHTxd9tKlG9dPLJXNjXBFVIvhPLL4JSwCP
+Zc5A5wOH+mSeIOLLfrIdD8yKpU3gCtbfj1WI4PB2Kc+n3kpVyqNAeCXm4cA
0BlFylXS+s+Yhzu7k7/d8ynVASskYVo22KRLk4XjwbWxEB7nOoSGAtAtdXfw
9Jm6WN2DJHJ74PSXKCZC98WGtb44uZ5EiRDqO10Na2Nl/X93jsz7ReIpaD5o
Mu5sB0JfCk8R49w3pP2Ft80zepNyA2e6Vz8MA/4CEXfpRaGXcyp8FnFbRbbh
odyh1WBGabN9vQVZEp7yIeSPlVdpEPQnGmVAKQmY4BUYgDmKkd0F18KB2KnR
R/Qr4fKnTyzt9eaudfdw+xsNRN4Y6kMWfZf2xWnhrdUmjKrd8mu1d1ovhY4X
yZqzAJ0eooLVq8d5NRhyXRcOQV465QlwfqvER3ZMTrIiWbIequru/YzVFGeS
gDpzvMoiQCvCIfbgbgyFqYWcjRV2ErS47wnN3h49h5jDeK1nwwgHVcRacFPR
2qQc6YU2rpC34PiNSgTMJ1XFgjuCAG4DU5dya0D+LDQig7sYeQIFuKNImvya
543yNR+r7NchLqTUmiWu1ScUN655hZ24UwfXS79vd1A6s6gGWHOLGum5XkMg
oeXYOlbK92KLmNMTrJbl2EBkQ9ZTT8Bm2I0hw+QnsP2qoMFPz/ShtAOVrrK3
a1ef822CbkPbnUWhf/X9elkfDfwTZZnRNQrFy5IwK0KK1HFLwsaV5JgNbKfy
0aof6K9R/EdyHq+pu9CZGGaUcoNY0BX6JsABjarx5vO5KIWCKSPE5+/obIGO
ncq4rJCTWN6EFuNIqf4l56XR86ggNxD8ERXP/tx//pcr9Q0hut/dU4KyrQeL
R4Z8D0Bp4PrKNXkUCywLzYkinK/QJWw/nL7HXmo12S1l3b49oUR6U6SQloCx
tEbquc3/WdfD4tntjwsp9qc9PnBnWrO8MHOYny7dRs+a8Fol6PSlfPnY68S+
5/lxHu+OlZDtLtUer90BTwovm2+aS968LP4LLT4xp+7v+0ehiiUzcCdrlFDx
4awSrbylSo0mGLfbxvHEtFKjvOn1fgDxTaLnInoaXMJF8E8WSImZwV0ksYBW
VJMzS+qjF1/v5tW4gLSfNLmlX8UO1RqO/SDqpm1MGTJ/U5aOUoNu/oELc3ea
gr5BeexmPNW38m2LxMj0cSNHhj92RJAME9fjGZKmOOaapUo9f/HrZkuOwUsK
tZ66AQKA6vQu0dPJvjovFeXV3mkYf9VCQAbBcP+F5xUqjokEkySgk/u6k+fK
HoHabfKCTX5zswxDQSIn4xYVi+0vys0wKPvWaPrSg1Uv+zGTACyfTByW3Ry0
OfLWo2n+a/eXmc3l25EUYqZLUaVtYUeSFJEwHP489g5gvJA19hX7gPYsyj4d
gdsSoxbmdpjOg/6aHG4ntbQ8UBz3KW2v+g3GBnoIlUww+lFwrcogpArSkIss
429Q0iUQuFnsV4WEz6LGIMnV/94gvG3KSBZsCPFA50E4m5KzG/D+aLorUgQW
mmFs4CYFT0kvyerlUDqyfnd+BeUZIt4kthywWzXcVBNCPJYYeytA3EUSdkeN
WANs89ELVnYPy9Y5reMLTJ+KOJfWYuObEdEO0cisB+dIJ3UKe9yuNgGza5cP
g39vBF1qhhK51DUef9xrYTeO3QJ0tfeM1zA2bOIX4YG8nrWz49XmxnqgGFIH
0IVtGWDoHL6/DsG99dZw6HWNcNbW2s0jzT4g18KLFVsUHrXuWrq4Ds05uX0l
a180wmRy4vyUp7YBQUmtTOIUskmJEFX87bpZ3dqBTjxCfePJWLKGNtwbS3Xh
M3g0sgYCXnJqec/u8c/nRKfL2LAzmWKwq0t0jaWwCCNDHKpGg4u2Qc8rgQOY
3+5oOQHz8xuPq1SYe79erRhY4mmx1ySQCD5YzDJQhkfo5BDrLLpoDU39ESRX
i0JMQG2H5UIITAzCYrwAomxh9tTIIsHc0i1ZyxYVvVEMLt2i62FRcoAqjvJx
4wIedMNwvSJ7JyxA10qF5hxAPST+VHLr3geT2aM8hboCgpb5uH7qZGGqwDoL
sYhgE/Cyt+ApTSTMO4VnFkWNg5G4UJ+/RGxlzMyAEXgg4GfpHyB6hgE6+Tiq
q0I66FV5YkwBfv11sOAXWHIEBr/UyYJbdvqbmGIbLNyCZIeSAh9y+P3UQlav
f5iiWKJAMFFJ6E3ApWSWLFF6SHerQ+4mZAglo5AJx9uQAUQ3bVM2u59Y4C33
1Vn3x9fxx/yFRilVEIMlaIbgTcBfRuMtDID8X1wuU8CTypzheHsx1ktg+Jxg
WhuA7Ui9jNo6rk2F41RHtJr5Sq4dMpHAINibGPixGBPOgChnQquCyNrbWOh7
KihtSuN4zyyDgrQbYeBHo7JBRodxwkegspU6laAJ9pT8i+lYZPU8NFC+PzmO
QcCrOiK19ZXAWrt05UlgELAwXmMnrFQe2T8lRHE2IjBgigmOW535NdfUtRhs
3ckgmVLnKJi3pTvjN8NhvT2fNNeWuHxxhq4JDC/xJ46EZS7tBObiY96r+6V6
ViZHQMP0CxjdHD1QWXSuMbuEsfhFELnGUbovvSMqljaZhQeKufMJKZHDFWwq
JWad5r8rR/JQd4pOtLyy2bj+dUCiILD4qbGlSnc/kxyLpdJKnkt023vRudZn
6jOPB9bjpQArL1ii+deSx9JiE28PlH6qHU/szDi73txCWv1EPCWm+LbxMcQD
udFb0eUC+VBABDrkfDMQ+vxSQRk/8D/yLedSBjdd0fdTdxZXoZvQ2JIHHY3F
ZUZP9xVriXxdUnvEF8utKDm6wnIYeQ+yU5SU1uMbmHAW60n1NA2XmZ5m4T8R
VWLnz//s/sUIHAAV7fYozDDckGYfgIP9a7Vvb9c1qeYWX2O8wX0hNFUU7r4U
V8du6UveYgpmQ0E0n358Y1G2FkEpA+2M6nS6qk08z6BpAeJU06rXM9Ar7u6d
s2Pki/6+fmYm85FeTtfwfQECgYwIMIJJp7Ll80pF1W0QyD0Nf2+PGfYidxV/
90HF/CleB+jFUTWvjHWVM/o7rEIotCAowx436eMmuKm3cgHDBi8BEVgHnwvc
igIAYSkLh0EKWU+jCseCLE+nG/JVV7ICVrmmJV8weQ2WY0vvtHQqSzN6rLG7
V26EzKAekVKrbIiePd+r2u5eiHXtttyNWLhwReyD7G8av3RZFO1iLtKlwh0H
sNfPriaCgm577S8B8Y6ITY86LujIkadrdkBzhURyjt+ZwZR97QaeGvE31LWv
7GQA3JiA8+wUgS5r/WC2acbXHel5YAomp+ZCMFNvjT2NFoIazI7hn74XNvCH
JSExGiAf8u8Pcp+MnjTTfVS5GJ16bwWnp4Km6ODEQMFPQbnec22cSWXZoNV7
MqQ2c9SmmX3I+Wo+J7h1R6plRKsd8vshYXZ8CSo+Df1DHinB6fNzgljZbvJT
p+KQMCvMivQ6CQL8NpjpgqZH4RhE17ZAlKNKS+8/2K00OIi6o31ScpoYgT4N
ORTkRQeZvHeLhG4usKD65jXvnsa6dWetyCR6QLtIO4Ah8asQvnBgNw3UFotc
T9wUllhWGVmEyI4WWuodEKmElr2b/5HQgkCsr3/C3d2/SmqP4Sm6yqd5KzZg
aH3tE4tiMZ1OYpInjbQn8ucrmWq25GlU7j6OMWT9j0cor9wlkQwUKWolykrc
SQ/KglYa12LPGObiFJ3fIIoHGqysj7ptfT+ws+2vojDzAvYOWQUazAxeJBCj
2tAOfgHk8oasF7DxvGI0dgj5msi5CKXDmxov0Oi8Th9OTIofMYEggwOU+yhK
lDjJZe1dUb8pL8o3HrlJY2/3/2zjOQJzyCD/RG1WtPby29Vsjk/pLqEn1AUz
qJ8RZanNTW3cJrsk/TGCkjc44ZcMqWcBpqzegQHrx/OvZXxQURJGXCng2jeq
UwXYSxx3XZfOKDZ0K5JRYcXdOfOiwQVSo+f+1ivlTyBII1vx2K6tmBnbTn3f
IAWjpp1KkaOVbMOyFpRwFGIkSA4GAMFtre42mcV+ibKhF5wal5MYLKZaqZyX
4ivyKE/vNSkClc539WeBF/H62BMQ6Kt0sfpdJzu3SDWmFhV16xdB2VFJLMc3
JaJzQxdSChsWxVqoG7D+1JCVjlwjNrPr2mfJ8AfBCydKB/Cev/W7WqU5IQ3v
DYAzXfB4qCyPAh88Jj90eoFxTZtqkvyOw3cWYeh3LA7Yz1kSltKEe5Kw8aY9
sYtn5LwWmMN1gnUjwiwmi1k5YAAdpB7+VA1ZcG2F/HflD8ypxJr4NdUlrm4y
3aNV42yr84lnCJQ5x2IzjMvqgzU+ehomrcVkDx2azuVucDJSZsomw1I9JaV4
mwJSKsJX8VqNqvdyW93vrzbOoroIyHLteZuPWPjlT+gSyteCuk9PbdnkKHtZ
vi2L/p0dPgbquuDWebI5SZAlwvo/GtMWZOGZ391wd7M6S7QQACNeU9UQPBR7
+rNcZPR5LOwlw6IXq62TVN1b0XKgA+KBVkhiW2l/3cWiP1r/5mCymNLu5rcH
ige+q4GACTIKb8Knyqn7vzz9jsB4FacjdTK5psK8mu1dWL082GZjxK5G7vH1
dQwAbbE3DLdH+qyMcjIgVJWlL4g3PqAm2o5dvz2oYEAL4bgzQxfyp3NSa59Q
rcoeFqUYG0xMV79qT0rEe504zgMTT1QRbxkCd2e/pw2oxKVQR236lIRJFeE9
wKr8luKONn/VeVuQus/4z1CnqPFA+cqL9TKyOtjm6eaqqUW42ixfCrE9VE0o
G2psBj5e2SUp/Ck0WnrcKcX+e7dfYNo0DefGb5nyIbQKg74UhWPt1yLyp08B
23w7X5ulSUdhU6tIIgAembl6e6y8l2MoLU7pg1mT0cWsHCz63xHD/yxxhimm
3Z7b6qqzg2IW8kOA6YCvfYOplW0NpkhaaI954EbN8VO3/ojnlTmL+FqdzE2K
aEJbRHimFxQmf1dOIovXUtVM56HOLKf63bQ0VB2q5pD+S4DIx7/HBqwcVA2T
JsIZcd2jOcLnirCDZHGNuO76iLLtQup4Cxgll+uvcYAOEAOtao3erwNFxaRv
o22Kb1Ux1+mdgh8KrLkpGmHaS8YdWv5XAnNq1azSrbH88HhwF44Z6MMcV2Js
Pyvw1R2OSFrX84/Z+epZ7Za/L6IMzJBQfxTgnSJJkw9PZLc8p+OuymVv3xg9
YJuMZN2WaTT2h495f5fluxObqAEk43fwP71XjghBziDwu1LNGRhASOZXTBYK
yy24vKo+VNlRTLqCawYUG1U44QIkKlta8o8/Ga1uSpGd10S4Cwd5rGKm4/a0
DZjHEnSjTBBnyTibVqsnkA063cyDanxVHNdDn0QvAb/0bc8FoSY1DsIjkVjb
zZeawPskuXklWBUAAoVBWaCE+3fA1f3GkOxCxgrGU2zmXVvOYM4mDonKzu1e
bVDot8UsvIV4Z3022ppwJpJdRaSc3OwZZEiNpuP5t3t9qug+5mdcTxW3vlmD
D6+0b5QeY9XxXqH8DZn30S4bdCFrxzZeYBGfnrjtSJ9V+Mqk9A+nmIzJnXvM
mG6+UB5q1M6qFzyekcpgBtYvF6AGjQv8gV1VJ0dJO8StYbVEe2MTgNL3DI7u
Q7bhgjyoScxPeFEKgpnNWKhcT5zsygKyI7LPIRPEtEe72gdCI/spRk5ExTuT
Z3nDEVS2RITjpuJynWF+WmDXDtNCCbQvnz9VMaC+U/5QUUkj3cATkTtocdVw
oPJoBNJkX8nhNXGyZr40slAqp9fC7ml/uXvvpsto9DOv0hXaUMQ+2d2reANl
g8JzkkvEEpSP9JHt9kXVep6ysKZPAxMdbz8YYDAOMImw1QTbtFt3CpqQpXU2
3F4dEJIrZKIfnfRMftCzuPt8DqGAWrRFnzCjlb8L3NoqWwXP2ILOmB9CpJ0r
ySFX8J6P0TgmMkkFjCJscgf8QTG1IyysRtwOdbCNhwhONW+4q8KaLJkP4VY0
IgKUCjHvbxp+Fxg7U+Vgyg2aYRU8k3twsQXyGumawPIjNi6FPEitdO8tVpPs
f/G/4Sci/W3cPT2naS6SvL2OkYfdwLd+lhdKdFKrupuIEN+6ri9CS35NgiiB
EjnnHGKU+PqC9zTZQl8mAs1pS7AkMRbXhNI2bdpRZtCopm2S7jtlU2vyHBoD
YSVDbLwEXuBS5GQbizKyZg4TLwQLUScNDD7gkHBHibooUD6PlWep5WtqHIzO
8ATZpKFnXDCAu8Q07azFB5rVF5mJB8ATCWbBMZHgXNzBSbCL1xa5otfFa+7s
cuMLaIthZu3ckcf/Ul7wDMWsYij+MSfmeiuXhzDsQNbbpuykJotO6QM6Q2uW
/+qQBrK/jmMFIeip3A3A63QMKoPCPP2Veud03P9pfqQLiPu1W8+eFtc+giLj
2Pnyk/c0ZP5lNYE1wae+mQceLxUNTa7CPRovgDKMdvgordMc/ToyVkBcUtNZ
unXoDzdIBrNtDOdA3f1Nn44zHyiwqY6uI6wKbNsU0CBpLAJoMZQ5aorD/+Z/
anODkBMjU3LxI8ar5OEK/bfCW0bqs/ERdGHpga9aAW//AuL7wVH5W/s/YSQ5
6A3zWnXu+8yEzvoPXz4XX+mw1yxmRJ/BmT9vQPY7oRqUlW7gAeIXiwbbi3di
oo4VpCdPNU/VN85vthxQJLO4PqtHfSpW6lvE9KB8oajvHTE+bbEBv/+S2uxd
CFS/2wIOmd+wHc4x/8Nl89tThSDtTEGjLhNy/uZDOT6B6YhEPUD7HcYCMcKA
B7OGASIKo7McRs/KVmgIX5FTakWVCIvEbm2g2YqFHtWxA2CUDAHHU5SYPqUP
fIg2KgXH3ujx8NEV+I6z4EPsnS9SMC/5yto2MNU3LQZADMzcS0+KYe8m3QCF
0Fs33Sa/9Py2aVRG0HnaIBXV1raz+CQUX3ZkKDjE69uzIR1QXSTcRrW4tvTg
mrdFhpCgxitVmOwPyhbmJ4eMJ5lZDH75YWylAWfTeRbsXKwOdCrF3I2BXO9x
PvFuEj+R5Avk2hJMeZxnyq5hU+KAEeiu/HPp0sIjEcxTphb4xDgqp/lBJGsM
vU03Wg9q22A6uR4YQsFN070qK+OrLh9dNrMQajiQw/fId7GO5kTWpEIOTB0Q
IPTiU+A8FFsZJCjQ+6jhcukX/BNJwknAD0jFre+Q2cNftt+H/Pe8nEvoLzKA
J2cGG3L9nsqL0ZwM8v6ZNRNve1pMNwHBXfbBnZK7rNgxC2iHK4ohBeisyhKO
257Nux7b6v/NNdnexqYn7MdmKXhAO+x3wLF8RcDuQxH6Xug6n+oeXBzNYm+Q
sF+ZUuPeoE6EhNdJf3OFzGrfMTHP8Vo0Iu1eJYFMu9Pi0gOAvnpMQ1mmpsPb
AHzvmYBCWEW3CtcJIMf4JiM0m1vmgSALjUNdraDezqsRzdgwX6QQt9X8bUlj
GfLcL61WsihIN6oL8CiG/+XEPh6kte7HqqoekVaiHcNXYJS6zoJ35J7VJISD
HkbBAXl0R4xvaYUAC29B/CQChMblVVDBgtG71f66vpfrhEVmWegiBtyncf37
g+zHz3qoIuXw6u4CF9nF6t2kexRO7uMB8rJJ5npiuHaC4nUYCewawR0rvItr
wpabXGAk53hAZ8ptYDpvZOgeYf72aVjLnri9bvztb1LjHkNCj871t93nabj5
BJLcXWwV8Jh4RcUEk7SWzVqbJg7u1eMkasffOZumetS40PcCz537bcjF8tWV
34vB6zzckzo12ZdbirTxf1q93T+PrzB2UWNlvW/NkxO2pXhrP8i1CpR6WFN+
Vhokdnb0ilkM0QZTpSIqaOKJfsymlYCPJcFcMjOCpQ/K4o2V/q6aGrdL1EBg
NUHboj3wDYzhhsK2o+AhHJoteBrB/VD0Wr0GKAiAWsAX7KiojqGyBYtqsI0r
D3qmDki+CHlh3Kqca0SB7qft6bnV7MPHI/tkox3Pb1PwEgzHvnPwgzP963oY
DTkWf/KpFxdnBxE0kYPmAlTHOu7Pfk6bsFM3cDyvrtu45JPkI8xLbUFqOfm1
GPrnEaSs0tUASXczRQNLXqLw7rM+Q97CECb1aDKF+O9PH6UJHj8i/R+c3H67
7miAmixJ+U1j2b6gN7eP7aZbkzIgiX55npLhywmcllkkXDxQaJdsoZWgVb50
sgfdIGAM2OnDuNjuunzEv5riuQEfnPCq1eIs/Y5Ae66/HqgVnMBkz1MUIufM
u6YO7fSOT2Fsy9T0MpYIBs95mdsiAZ8MrlP0PfRYnLbo6XP5fkTv2DLMBVc4
vnsM3gRazL+j9YuNdkkkFn4tqDNnlUyzVS0gU0V7GeFBTdVbXvmv/QhrmSky
vsYnklNoU26RyDXmhipMtQ5nTdaVTEnMVWvM9DAejc+3s6pJ25T1mrOdS9Rs
MFWjmo4EwdhSx6xyUrHR342Rx3Dbsi4hKzVX+mI8y8I+Rs/xPk86OrAd7PcM
UcY0SXwAACGXaScG1ke9bGluh1Pq49VkdwTqPX+mWXgFRHNVypxZX1V4xjGh
umEbmYrKOKAfIytZDPnY3V9DEqDjBl7IZr8v/tblneMP/l531yWcK6Ukv/OB
RkR3RfxBoO3emIK/1KkqYBITxZsh1VFJtRIWOvJTyEHmtZTLqy159wXIwvWF
m9jTkhIG10uLpF0uYrue47qWaNicLwNyX2Exx0dD7PQ8k8Gcr12/9f6RXy2W
jyZaMNXjS2YfHqhpvpYeO49veQw0dCte7VJj/o93726kfoqk8TeK+qesEgMG
/vmWV+S96JgJmv/pDB89b1Ogoy52JWzqRVchb3b8IlYiakSjdVUBdEsTQxva
PSWNLMp0i5kxWAY9a+9RTyqrWQo8umDRyTN4HJn5fy985mXFAAusEkEQl7Wg
09YWcrIcFEEjkVP7X0ihOrf4rcbHKxDAYXKv3rlkjHXrx+miHfgjGKIi+BTs
CZgAYrL/2g4He1+jfPEq8/khR1gf9HUdbd0gRrjgNhPQXdsmh7B9ImIlfrZx
ZUl/c3LF/DncJAnCldBGaiHidTSksyYTaBMgixL0eEooobkFiv9aNnVdx+a7
pVIjeBYx8gDcSsNPGSVMwpZCKD62MDICD7wxFUGdFmDEg+qgPzoC8ZMYSqrr
LmqYyjrT1l8tGkv9lxusFwB6hmESSWhCquqOBA1EOu9dWmMQwRFtiHab8bQ1
/t22OUrDbOi9XNIPpbTWPjosttdvtG2vmm6rJA/TrcyeL+yXIjHElO3wwveV
FD5PFnCvi1FoJ4MYexF0uTX8R5VWKeGgOO5+BSh8CWHJ80AmLoUy2lzxoZV9
44LFGe5+c14eW60SayNJ6GI0p1FeBZZjpHqsPP2BKwHGIrGdKTgct7++x7T5
ZirogEp6uvwsVCa8XEZvIykQh08vWgltkYR1Y3WYMVq6A5lr9XtWcy0O3x7D
AUylfiNcwhtIp3mJ+dkY7N/wMj/djG1o1lrS0gD7cbJG+Nfy7wqIHQLEu/4O
wOj2R/2pwKR9x+HoS1+Oq8mriN+O73fhdfBl0tNlCeanpaPzxOU/ZUxReB6Z
NHPLhNj+/ZzjGHQL3iFWc1tNxj29WgcHcsg5m4+uanpvyjVWtlUhu2NIfOyT
NvuujgRMJ+PzpWqQ2mOTQIspTHfoPXC3FyKK+OPEtebjP0UP9knWwBDdJfxo
I86i6jcy1XkN2+I4by5ifixw1npMqDB7cr0dU4+gIFUHO/O3fiT8O0CkM1Fk
mAA4BHNfByY5kUrpRKqorcWsx+tylrB2SIdJWqyl44V/O9QITirDsHnElqPO
MPND4snsN0ya5p57eOzlXluYXDhP215P/FVajJkABVARSqlFkqORVbClBhst
rFhXnxrIgablgXXyBWxZq6NxTN2BxHQd6aUx7tyzExPs+qZz2hq682w2dDN2
zQdROJOi7QKbHWPDdE5hOz3pkxcvJAvk1//pqR6GSmX8j9/GbaZw42MBSwBu
3PHtymJK405xUdLbudp4Xe7V+b+EwFo1JHzdHbce0kl0lWECMIfFQqaK1Kq+
bpZ6DlS27jg8Y8VeT2oW5qQPfO3GEUUbgB2cT7sjebS1fN/QKOaSWcogH/v5
QKZ1P69Hrkt2x+2xu1hkKlNYjeegs7Wze8Efd84WCf0tu66fQHO67cemnJL0
eOG0FVUGHsJDBFXlLY2wttIA201edhJwFfuLYsoHnP+YougbBPNTFLWIIusO
l96BDCJfAT2EURUyKS7oEMXSAmjRFPEkY61aR1jy7GZzNANWAOAxPqffwb72
Uh1Xi98C34DBtCjFdZPnQ9gnB362yAQHZAnO/NDlXqVt2ATQxV+DaHRzaygx
LP2rQ/d+gjHQX2xKfKil4rmFLuxg5l51hwUi6YmvY0oBtXtqdN249yidfo4B
BbIyWxB+F7m9Bx2O6OLhk+ThyNlmqVFRMJLR7nRmjrwD5xpj46OIwpDEWbi7
t3/etIuTbCR+Go6pwvkpr4AjtyAfYeHOFaSFLNazx31COZ2MJ8zKwAtxN+Ij
8ZzYjYXPogqw4Cj3yQ9H4zeNa0cYOqNaxTyA63wI3Gzl6A8CtVGOPe5PpjuU
X6krcoXdN81rmKh9AAu9dn0uAQc1o7tsYvJ5z08/RsmvPuqzB8kX/m01obKx
5AXiQQwQJktt4AFHttHOUTXodYJFJrNscbc1u8IFViLcVGTCuXurkdXv9kFE
IefZ3E6n4T1etkier1xB+T78CyWyFkOyk5tO5uYYX0mzvuTn6TOAmRaRroIY
QMd66kAgaVcZo9XLnJDwF1LDaMCbu0yqT1IRemQJ5Bzq8MNT7CbbOuLCKcRP
V+DB9Hhu8lCMINxYIsHn+fva+cWOqkAbr411gWoJd6Y9iXhfDaGrvVtawzjy
rK/q/uiQtCUtEl+T9IJrNUleBsINj/yyZQYBVhi5A54fRYLi8hQoL/J5W7aj
hTPtGzxyuYy/YgHFkqafl8B7Kc2T8JgQEyJxPGLEGdYlep9Zzy7MQMwgef73
Wn1IL2Txn0fQJUbUFiokfno/Lg+u046x4TlV77n5TQqcMQKxhcFXDu1f0m+p
4JaQemZaohPXSlL33zbKxvJ9WMgpDxX52k3M9VolbGfTV14ncckbUn+Z42GW
N+y4LTNnLCfuppYvs4YEq8CjimtLpT8CV4/RFqnbzKtfqdQLKDrXPLrzxf/P
k77N8nh23jk8PC08QWrN4dwmI8uaDko/rDKRzi805VBPxH4ycbzmguYy78n7
AFYVN9vcH9YW0d9VMK4Nh/CJ8OphQeWZm6bcgPcpWNdY4d+vhV+pmEPawccN
Dl7EHe/8W6TbnWXavQU/Ulde/gzi3ou/MYF+oJKNvZe97YWOaX2Vt59DuwvV
ysY3NpFiTGdaeBH44o+DEPoQjcpWSf+h4ZwK6fOI+uwDOiADEskgmNVxZVpf
Wr1DLdN8c8rYiIyBm5lUUb+beLVvKafNjwVb2A/CNwotYQpUqPgD+l5/h0ET
De82g3Rsuga1K+MStf2xPqsyo34uXVdcZ8zmM1qY6UrNH4KsptKT2KbUsdBo
PV3vRqVuAtHQkk+nUMhtxYJB6ioy2+EAj8sib+5IAB2xz7kWbAHBgxFCb/tE
qwxusmkvXtGHEflsHoVRSMRWOJaBl8ApVasbw1aanrRKh1pMDDnfjGH3RmIh
rjNZYwsRkUi3wob84n788vMy+SZlP1jVGgVQyTXC4eh5iwxxaNQzTm0R2E/o
MabY7uE1saJ9K/sgnsU8QxQi6dDWMSNxsORu3BzLbMP40/y6Sx3+A0V6uzlY
98+yAbHobmmnJyz3q8GyjtSuthgmVsd9fPsz6STPfLm9a/hovkQFx+zy6T9V
0yq1jFiKQqmPq43ZdDmXe1P/6Iee9u/cbJ69OcxBuiku+UYEhkwIK/nt3vYe
RW7aMMusIH5+MyzvQJWrBZiEueGdKwjQp7oByac7Cq2VXQA0B2Epr3lq+VFs
MZn0ouUds1OgnNHUt8UCX8V2+99j6Ei7Mmc3IbWmCWbf4uKRsJsGKiadVkSg
e4XMTumFA7STFz/IOP/FTitcMYxwwF9+j3cGo3gbX7xog11MyhQHK4WFuSdF
2Q+e3hWOghqeqeIB2UC588y98LI9xz1EYCfy6V36JTAL7y8FXqF+ygV56SmM
qo++7WOhseRY6mVFGE2U/bYe8GX1W8NNTulkPSKDYt59+7OuxiL91b6S43A5
9sLtKz9Agka80hdSBft4LMUr4tNd755AKv5Eti15e9g3/UvLaMfrhId22WpT
GRcYMzNhaczO85mcVwhfZVXtO+mE+/RM9/DYOS+za1lsC4+ZPnMqORpdvK0S
c9IlFuMAMX3eOGqVO+DFxwtYakJGJ+aY9UhAnEMRuiyTGDdTx6ytleu6V/1s
eU8hVbG/dwFMa1Bay2Fe1MwOPT5jPZH1mxwsvoZO/tO7YzbjotW+Q24aFsKi
HJydIgaMUnPB9SRkrK2L5iXcKkbgVtBYT5pmHATydULi0ErPu3N69WU/S/hn
QeS4XqWN0LjxKs14roUbO8zr5vyzwrkl1NFLBiAf8/DWlu89mASo53LWJEYB
YlTqBMf63/EDYH5BYfY68Ui/wTXgXTKxSkO271zNcFAYLPGoRyD8sZo2mQcS
isP3XOX3R30vvr3wjj8oiQP0KIOZJfYgxarFhDV4zeRWA/uQNFP7YjFQ6JC1
hcNKUHksF9npj6F9wKHnewMwdbfR230TKMSPfIGexVTfn7RbA1R92HL9Cssr
9dgoO6ubaTaqZNZRTc8e/lDNLaFEe/qmBWIWT4lIlgZKkdNFcXDJh6Orzt46
2tJA9OICWjAuS4vmXvDZsQAncjymtDBCkV4l8w5MKDP4EzfMoT0lzvjwduAf
bmG3bVXt/5+r5DCbFdY/E9RZhGbRZI2lzHF1Rong+jRKG33l8Efngkol0Lt0
DEzbUA/MrpEGGIVKgZcfCV01dwLiLHxU+R2zJtHMaI+n0BIyhrKu+iygJy0U
1vjvCRUmjd+HUqKPWExWBYvhGwpGSu6Raqp/gPOFRVp3bwRlbcWM6IfKczW0
m9yxdXyemPQl26cLF6185SVVqI2HCkot5u1oExP8PUKl/dh+8ycnxIUVCvlP
xaKjeBBhHkzt2LJR9kzL8oZd9L+cjKrlrToSd/jIVMGcpI2+6M86Bed8xjWe
MhDOc0+0/Nc31WjzsVpA6kePdLVtbhtK+XKFTXL+fj85z/mLnp3GMQ9gIMC7
V3ggzVFe9YEQNx2JBxG4gyR1T1onmHPjdZITB7Jcu2uSh/E7xkJRFKUbrafr
qYto158UYy+/4IDJykSse+b5mRvcmZfggODFw8znRCH0wDdl4LEn19EXHHdp
2XGr/yCm7DI+SCEk9bG2peXifQxkhHdljZEZimZSJyMKEiAe0XNq4R3dait8
B6N7kmsLruNTvmHZC+Gtvhku1ggwOvTvXi0Mic8A3y/2j/8eTxGtg+Moo9Iv
+Win9jqdcwrYtVA4faoPRLtlpJo+7v3hNf9B1DhB2QpiojgKFQBrQma7U7dR
a6Vrlp/Cl9uEXeCx4TGinOtPGAGFTtx5h1XwJ41TNVv6hhhErA4FnNhhUuaV
rwzyAzEiKyMv10muFUfIOCYORxKpzk0FJquNBH/RXoYdB/09J2Nd6uo0oBly
W9ZB8QniZosHFdjcKw7dHL7+4T3e2sPxve+yt7gzhoSh0qP8zCv1ZAp8Dy4k
mtSe+IhzBwrYZ3O6xqK5kKz8pB1/DWpP1BN01pWeQqejQycu1JE1YD4ZUooD
k4u2vTAuA3HfWHeeseGurXQRY+sUvNXKpiPfEC6Xlhbcjnuf34B16Xvo7WUi
ipnFXKSuATjT0fw7pJytzJpqxxX2zGzKBpRhUsc3Eip7kE+SWOQ5PHaohOEj
3S/rFYlDM8JF0U504Oi2wrSzKVmxumo9Lj7P0OvMTux9y8IauZB0ZwzxTE1t
FdtBZ7ojzfhsNRqjtUxIPPn0SmDiks9zGGA8oPrglBsu5kBEjYZwZ3h22aR5
VUN+QhHO+sSFO5f5ZYFJPcM99FVgfFrk5Lf25i41Gqm+U5CeT5ngk4tlp/2w
1m2Km75RONL3C+ZBPJfDfD1x9cAbyFXHgIk3cvkfTC5gMyhNhWm8mIBz7ajw
WKQvG/wo/UVEHrFj1gD8R8/rebVTGa3fnM1fF4Ihhj1PbJ6xtPT2gQzcME8P
HDfPD4W/uWQaL4gqAEzK5Oq3VusBdJ6Ky1V7DjQimp5OeJjlSVu5Ah+ms6rx
0nskHoAzNChAfu9IyTGRBws+hO1slD83kyDx6FhJTQ1k3UNv87o1ynSjnIsK
DbzHsqxaiZaKBppqV2s1YaHTbyxcVXn1A4xKTBYjw4NQlljUkWLks8q8g/oo
YDmdol1efNUzUh0ox/2e098K3wzVws9XNXsWXcVgM5nAsFpVVejEzII7z8eN
yrlUkBzxO00lpGVrtz3mfdeDzo1N1PUlz9a2sRHFb2QU6uvlJDeREzap18n/
aYlZrEsUc8elL2pX8Wx9rNBt0CA97oMOLw0EKTixVXawHvTRVBJsILwzDH1n
TqZV7pdHYADGr9SPWlv9eT/2Mep2uICjy1ZTxdPENYEX/BUZI+hrPOUqh2F4
lK/e8CW3HRJQVYNy45FkXFKrDcJQCJVGf411Uym/o6Sxg7q1N7qlneptjE15
/6rohnOZV5UuGnW/4B/gCyHggs/kpGzFWfdoPN1aErxCocVRkwjdsM8lTh8s
cOreX+FM9OqJC9KQQjn6VkH/OwdgtjA3ma5eX4YFN9LfLXR9wmB2+WEn3++4
liq74OFc6f2GBapW3gdbtdXG9E2Dd/vrdI8oBBBcoERxJn7s9k+mYkAzfh5p
Reuim5D3ks4vDNVmMvxUVl/gxt7Cg502KjmTZq8IeGiLmDFXUn06n2+hRFP2
qf1pU9bmB9/4VuYf09e5TT5yIdpoXsCzphFxn35YveI3AMEM0ZakZUMsip+f
ildG85AuBNPaVijcoHNPy9VyMCyaO6mHGkQx5ZPnj+xJ+7iYFolyRL7fpuJj
rWvkYmi2iu2yz0Mve+DcGVrMuNX1Sn4j4/3OSAtNNnp09O9z/rltYIvQD/VA
H9ZSc4WeMo8RUUDxlU02IP02KlQjaSRjZCGlJOMHqr3+Km1ux07yoG7s6Jfs
Ybx+vDUqvwInMP2Eht34AnE8zxWFcn0Y0ndjkeODNPnZAwT/c7WkFV5wybdX
VdKQDeNIXghkAFgyY26PUWDRIhbS+sN7JH8zmqcrz43uAr1h9h3/vx3lmCFu
Gg6Ou+GbFc+K3cwjR21j0oiDx5mfsabESWgBfsJGSd/JfJYFY5zvHdjDdTXb
zbVjz+EQVskF1cYnYin3TSShUGla9zi78smDUKObRZKsx0caFn2lcnIX1tdm
BpV0ri9f8ouUU2wlFvIOxi+Hd723W73FxW2D5yhfaURNC9Mqbyih5rAoww+w
mUW+nNGenXexxRQJwAE4SMSGEcGYcD+N6pCZXRGM8uQkMMtT9D9506LJ8TuA
msYYx5of6Ee8Bqguz6hio5ZCIEShB/OIEG9fEaQoX/UgzD8KHZjKEXsE4Fwt
B1PaJnkXQIzs7yu3bcYtMo7nLyxsOevNhi0mcGkORahDpS1px6FkbHvQGZex
2U9/s19it9yVecOGa0hk7nkCFYgJUefpzZ1kTAVGaZXq8bcOyKIqJcHM6xKf
z5wMYrEznYtWgtbiEz0ooyAJptp5TKl/1xf8W7HBsnkWtVZCxg5cmmFNdyxY
exsYZpCrvZZ8VpNX4riif0iLr07+0aO0h52jew74f3B+NUkli7vV24povIze
JU7ZKOX1CNyYnMMXXYD5c4XvkYMxAhRwmbCDWZv0cdWGcE0oQkW7Qn4iuGBg
rPqsFKP4FgdKoFpfQAdCuU60cLoyFMfSknFJLr1tvrZjQasPPcMlbPoA9OHU
4NvK3NNZcEXejVZxQMXBpP1kJ6YNZaTUdaQm+O1lzkVHXBE5e6ImJtS8wRgu
vRy19cGxYBhCNLBIGwTP+phQ+xERjG4PWyYw3MCklWQjNyJu0UcQeNElL+tc
JMvlzKFO5xiJqlgpV5oWsJgTC36PHTIFuTGf6VdR+9dummmE4jvXk2GOWid8
6Ga21rw+Y7MtiGG8w0h4kLRoX1D9e9imbk5ehqCF//3HWAx7cSROef+YBDYr
GLqd34IyBITezJV877zaVabbqbkK5BFUNJoQ8efxEWA+miL9njD/OIExsm64
neOI+eQ2zo98fZRZIMLBDXWA84sLzsYWSe2Kjp4PzJp/wwL7x0NpI26XQQqO
o43SQ37MWr+4YW/5R7PT2xnFvCEH6/NVfs+5lVFF70XbmJPLHnveO3ORtKL2
YV6zmbiAQaPqX4KVuyw/jmYtaaEzTomgeqUOZhMCnoHVSGqibaSlXlxxKLl3
hZE41i6K2lKKqf7LddXzNcsLlStDJV9L55XQk12kVUNCV8wQ2plEUH5QyOd4
nyWjfxtnq45zruSpHOfRRMU/jS0JMgnA9895HzH1QwIZqH4sdP1PUXx00E1E
0AHKMW3WpxSP01Nm8bthHqIUUN5b9LSD/Rp1bzv5m5fyfTTi1/I3j8qfvU/W
jk/hMDBN6/e5zQb7JPSUodcvCBERstVwBcepOWuh7yOPSoYl+hiX3Buva1WW
lP88jdcpYz9wwOWFKsu/gt50tSOdse27JXo5BBT5DY9wPSSufLg8fkqz/dB2
yZknJS9ri/E4uP2ABx0ghE9/9F0O1SlV1SGabTT3Tbd4AckGxgEBKOrA3BJK
loIeEskF2r2kSSVzP7ck9BkT+xnP9my8Ekz5RTEmGIp0EVfKUNF72HjT0njR
hVupNgQzLTKCOk7I90xWIlN4Ab1VSgMRlPNG3L+l95XoykYLubS2biX7CZw9
0Vkz7ECd3M/SHuZFoZo5SxZscz5A/J5H0RkOihzESacQ0mTwNrBgfmD6wd4M
VukTmtvUwQuvBUkRDLomCeP2gJAAnFVI0iced+LX7Dyw8KuwJtLxuPloXyTQ
yuHh1QXmu8zoiNU9DjIiwIX5EXwITA23jXgjAWG0zG2eSRQ7LE8EES7SIY4a
Fxcu1PjGvrs40mfBMRFwLED1i6cOVmou1sxIKzjSsKnAdjeImn9KnUGVBPlR
uTzNWKPFaUqdLO3w85nKhiC7EIxPRWqHhqQbmN9U9EYrxd9uErN7rFAf65yL
OqYtX+hYVX8Gwral/QPQNnMGjPd/pg9gQ4h5cnhwxE0UaV0Jd3AkKqCOK7MU
yUAKrv2pjvezeZG1lzCyZ5q/7R1hciKkrVJkveZLz7muo3VIF9CyW4h1o0iF
aOyfyqwL9xGdP8+gmEmFTeVp4RgV02781ancNQaqj/Thog+GThHcEr9iZHpW
32sPCIt30zQlnVgDoNueJRtAPTnqGTug/3hulPYdErTpFwTDlzVFHcj8DugR
mU12vQ6fkFNLi+yu3JK5+4qOf/MSrKcc+vPNMRvlJh7TTha4kPyYVuCrLQCN
V1fHajRd36WDz7NW72fw9lBLZb2hNWWkzVhPlJZpUHO7y8PsLstT1xYeQ0p6
7DQfagjZqiazwVgJZ8DNyxutSCFhuu5meIba/QrEzkHiBCm5keYi7KMzyznO
lZjVvQC+LEFinyg/jh/T0jQE9z/+hoJWhfuHPF/dLGXEK3EAzRP8yaE9o/RJ
2l9y+ukY6ZVTI+xMkrVo42DpyrX1dRTHUEnbcDbVbEjSfF6Pj7wRaFeseQnO
9BZFToW71xiEsJ4IwqrJJJUcjtntkPaTQpYOn5cC2XgYoydsdff+V6L8l6L/
OCveNeJbfuSZOKSrvLDkUfha916OBpIGztDun5RxAJ9TJ5w/k41yS0DG/Nzz
BXTLKn75DSeWVnvUNE+j/smlzeK9vLa09s8mcj37a3HTQYp9psr65Nj4fqiH
wojOII1fay13y7EX0hUxaM1HebqJHCqxO3FtlEbteYHmviqJtbK77NNgBnnf
XhitbnwGP+/a2gu5GqmbCDsq9fR7LlzpSONpjHP4fDnN83antaIN853CB5Rq
QNFuEbm+TcvCx4t0hjChqfkNcwFBdBahFMYDTn3F+/dRerGg42wTLIVDHAaf
w6mS3hKXuG5c1HMUEV9yiClWbsRVs0x+4QkM4jexV47HtXdK+byrQ3aaYF+X
iQWNsq22o931PTBtVyUES1w6kKsH4AIi1eHXvOY3LMZQ9sfG7I0zNwM7zeOr
92up6zvm7fDOH41J2F/caD2s+BmDi3maJPVyGzMzF4CoqXUy4MadMFi1cglX
/ErXFEvxEPb1bMQp902oB7JvYXer+NWCProkNxsVGauETHcDISkYaSflHzov
WkIq7P/JRn0EhVUU49rCanpreuXfoDLgSpc6jE3Gmwwh1SucW2iFATK5OzDS
cz+9KipMRCCCq3cxc4mih46azUGW2kWxzKLLrqAJVYTZKMU/ZvNdU8sdHwXg
I73lLp3ZrJrK6mWDThw3wSI9TmNo1t0Cf22WTT/mupw/t4jFdUt3VW4aQ7oS
DlWk44i6D6a6muQDjKGehyp1QTywphp12ursGN5bAFgWnzWWgxe6euJv/Y80
O+u5HNd28OJATVneVrySr4cRMmEAIsT4cYMV+UJssISc07xRXQaBTuAOIDCg
hYi2w+CLn5goiL+F0cVnX2dlYGptV8bLJJdYqLADfLEhwCW4FIBNxc3MAKa/
k4y2fB1mLR9yfE/6ZhNTBCJZzxD0okI6oxnmGu17wu7tBTme+2hqGTAErxvc
5TbujoTF1xaRY+rjlmkmkrI2M8zefEdwgRHXVSbb5m85mfBYNrtJxIeBgM81
R7qDWk51ALiQvHEVZJYja412g0ikd50J+nBIqEpP0ilWDhlo4XrjFRyqM+/H
7FEN89JSDv4WoHQ+8DL1cf2XNffipMgtD+af/qpJUFI6YLK/v6Q+DHJoEJ8g
R/srkhPOAWEiyjZL9iT6NRacM1J5D9/jtqqg950MKKeIMs+cecxtvSWy4xZh
5QlBKE5iVEZ6M5SJaoBp1xEzpjjBvL/236PWpT3b0nwBTZr6p5vMDDPwML7J
hkO8kQj7nKYIjck4GWgkAl1hktGhIxwION1ATgEwpTFX3OM99Aej2h8wnZcC
10fIlALBzbmGcIq8/Z3tFgq/Qnwd0T6En1XXs/krd42scGEOBgLRGuKCpTzC
b1Q8zKO0EbOVDEg1a5S4iCkfOiVO7m88HVwv8Ok8IwkC1cVLFzloR1D6F+Cd
7zhhU9FG17vjv/VYWhfZj9SDTRHjjSmC+uVc0X7bgEH3fmLbfYEQPRX0jlrs
lz3JFRRO6MLSgjm4/Asid2CMUe3BJsGLE5+/bQLM0M4lj/ORCETUPK8gaZLM
v2VZjT+Z/vxNehzpUM33X+7IFVTDdbq8YFBJfCKd4jc3cISldZiU/5WRI82t
A8LaTBKiyqfAnT2JsSGUviQj9WHZaf1sVWxhBrdACmB8zaiApdkcUoVuqqAc
uAMfpkExElWAJGNGmnZmHWpc4chjEDUh+CYGDaFcGqbpp8HAtOb0ysN56nuj
aRHrn6yt/vXRF+LbMjn7iCWupm1N+i3w7zakObC6kq8oi71QTeKyz7NOj7i7
XxUSp6OjoanPJvmXDRliRE7yfiSxxsZsBh/cFAK0wN6CSBm6JX2gzIn98qge
zOdF7j4EHf5Tc+mLC6gT3GM4/kY72PtE83/wWXxXfYiaoIKKbLUtD6m9UkmO
CqHwgNm20YK2BnPuBcvYiYG59BqkrlTFyuz2AfXLKVX42Mg3drPgpfZDiClr
vlKAbynKXa02Bjay2J8AGEsEbAjuR7VccUFHRdhLabonEH9/uoGAPlHsPQMh
xQLhc56x/lshEbBkQddvbJstTPS2OiYJ0ZjGaeWCI3tDn7ACAq4RNWIV9AZ0
V+Gf4WNpjf+pSvhXv2PpyN2fc1BjLV7znA0kr93DdQBb1gtocu4D5dLh0fcf
Js3170XpWSxIbfgkW183vsWiSQBqAmD1akY2zZEDOG73viuO1nCtFQoqpxNP
+jl8OVJfrGFdOthrr8IMDxOvV3t3CjDwZ7OqhNVjAhFF0ABESZejmn/9scGu
QZBrlyx6EvJZRQYHonwVCeTz8ThPIRxyBP9Df/CDkufYsMv5qSfGpMy2Xxz4
2GW0TM4wYUJk8LfpUBk14j+QA4nDZYV6B3oQQFSQPhkVTJJwjK1JlLabDwKi
ueicCEE58wBmZRG7DVfHwKMgwA1g/H3kBqIkVkZSY8kK54vrIqqefXgMXbtH
tAIflsBBMwpWVECchMdsqUeyerxTV6o8dw4HI4P+X1b0jGYECsVv7aftWt7h
UxPMpT8lK5Q+elgrAYWJgr3H69JlS1opHLfwDHLBMmIokQ6AI2ODxhZS1UkI
8yL97UdZ2nrFvdtcFbJG3+ke5oyqINn2j6PiVMB7voRs3fMBB+Q5WFJclPfv
CUKBna9PNFJ2cZq2bsaCOnH7RS+kbWp8IeUIxK0+2JtlMR/5BwtBqECpjfAv
rJhrfyU86R9izR3OnlKE5JMcg7Mdx/FNnAq8SdB6wRWN3AaaTzfa8fMxHt/x
55WwjQfBRkwFBwB/HLo0uKG3eKZW0UwFvcpsjmDW8kvwc2Re6233xtsCMx0Z
FK9kwln8L+wCza6tP7oTCxz2CiiDCdr/Q69Mm3Ab5ZNRKnctQb/PERVzngyO
zXWoE6IoIqhBaTehRHLL2Q1Mo3czR+FUHk6CmABfufsVu5p+QIndpsaSe/F1
ajDnmi1TcErnjC+D5zIS06KucghAEt/vAR8cBlKeazsobeBsF6uE1J10lkd5
Uwj5JUcxmv0OrKRqUdiv5o2eO3iPwQ14nGMn7it3b/E00Cxul9DJu1tqUN+G
UFeKX2FJpA+KK6L62LhPlQpb/rkGjl8UJuwlnYpGhEY9HhIaSe5dkhGvAfru
LX/uGVzz5r7w18qg/5Xwjj7QA10Mn5eUw0VZmRdsD+w9YxX5fACPirVcypnL
ycxV/ck3gWYEMp0q0BvHT+UyNOoDRHxqasY8RNrmn9ax0cFjlDtf7I1+6bTK
tnsFrBmWWu3tSPQij516LARd9oTWL2b/O3TiYG8zrq4fogdHfJDVTRWaGhRo
bUKgC3cd4eJg10CbopaZE/tdnsg3XvlDXrbyW/ww0jXP1+C+gjnFe18D7EUH
dcDpPSen1f00E5avRj7dYMZwe3dtjpov/p9DIPOBj78LQHr3CFvzRk38f2AU
SxSTS+wGL3Sz0XTd5T/Kt6AbmsuVmyj56FwD6HClaQiqpwan4ZOMn4Ih7JeE
JSn6tWwoGbWEXfx23z4h2vK6BiH3mjSSXlB880IKjZIY8yVTUcqfQ59hWsYl
kxmRuTwrhjzexcXDNyT+8shVFaXeaf+VkRc2D4mYXBT1iP/hxUs/k+hMW4h9
n0E6Cl3gKcIiCh/K6Q7oG1WTHGT+jV5rRe0RMcUe1OXN3v5nXF9dLZBtYjQT
Mc78Kert8ayQ+eNDJ8jh8gZjQbr65JK5My/SMIrMFI+Mj03VrTIlOuNwn4As
HBkjGAohYnniYuM4Y1iMwNBOjVud6TxqZhRgfTAqwQs/sWI7Etws3kDebj7D
jaGoid+tJUxwdFqjM7lqk1pmEezLqm+sW02KEdN71GESaBh0xA8Yhu0bzb4R
K8iWGOgedzBYBAmSKxf8MLr3j6P0wuvnOEAcH3S7E2wku8vzic23F2Eji26u
sZlpO5yCd7qEBWcfjzS7eRY+wvnC+7726reuw+GqtVm5/eEGSRWpimnC4EQ0
LDXMXTP4b6GN+3SR/VtawC8HNqKsK8FhE+t3AVAo0QiKoTbuNnBbnuvOEM3K
noUWr+9RSvcYdktFOlP6eAeaj2xw5JwDnIHjt11iDJRAfq0cGRg4E/Ztw0nW
QZJtQCTyQAUHWoY4wM56ywFyJQZlr9SsvULGB20Cm0ItFmHy56K2IVyjWWA/
+HN3FYIrXjjV1FLZzlN015L23Oaxch+eXB1GypEK3y0x8IIcMmZtXFVvUP5Z
ePFmKypee8153XKQAhapcm0d/kTCUKxtRCNmBpvO9mBJQajW5gkm4Z6LuQec
wXD4nHG8DYNUeqLG/Yhqle0rzBZFPWyuMkuOn50NGCafM9wX+b84fS3A8lJC
8hRuHmIb/6P63RT7VpkMUZvUvNLMK6Wblpz01lCfVTwsPE+NxVqWfgI3VJyn
Q68BbHGzMoFaeG0RiDA2/sPD1jR1a3AgxSan+I6te0ZuCMc8IDb+6b4o4xHP
CO5xar0LQV78LUlfg0LdXagYQrDXfnbPFmtpSbSMe3hB8sKXmCtQcDGVLOLk
lYtK7Hfai8u+xd5/Ft59tPieWSuBME2Fys1iHBWBszy9MoQk6TEhR2ecimsN
EzciIOQ9P1ij+Fi6/4YGED7vgCgte6AWg8hx2DMWvknST7qCYNOk4sAPiJp1
P2HDsOwkvJ4bGesMpf8GdozaP30jbEqY/FS0eTj8vSaDElUhgp+DFaY+0moW
NV3MGykI723XUbjyjwH8RwBVPxEGO+A3KmSJIbySnfIHUE/zE0Q/qNdhntxW
YXSBDIErKcbvWvroaaqmYYegZpxVvVOhG/ptJd3iH4GvJcL8Ku0N/uw7ynlz
Iua7Ktd/d+rBHAQl0hjk0drOYJwyuw1CXyi/nOXCdrZVNbjJcAESHt9h4lf1
4ATJlGQC/0dVPEpINe1WB/KIf/XhwM7OTqDz+oDWSt8IOoaH0+TfydRCtssJ
DgminQJSo/nuoPSNr/TJUIF/HyATsu6C3cRGc4SMpJU6TpgtZ9KwaJZihQ+u
KDSWsef/3KTh+FXgBsCzGpcbq3tXPHSexrfpRNLKIMTTfUfaVHzWGkd+o3bT
29MCGFWUr7Rdi49v8Hr9wjUglY0fjfgBehKMxOtEI56ZyvlvvA4q+iK25lNy
7EsMk/0XbRXKtrLVlOJd+F4OEu7qod0s6B4tQ18VGdg71B089obRJ5bhccu2
5Xw6EqlNf01JT1h/a4QLM59HUGPOEwCS+VuOjjd1chL3DZuFXaBLpCo2rxgw
OVQvMFxgLNCQoWfCn9ydteZK2zrMEEn929X/zoVcqVHxxxlTmmkljIJc1lDb
URxdiUDO02puvb6nDn1PtW4B1M3MqyKUJv5iTDvnQYIXyHBOeCZ5qnY4td+J
7qpB9q1mo73XzXVVTITAJI6BvLacIAcf0JheZ2QObNcLwEBavET0DHuDZv+v
220dvFTrOdaFQ4NuiOSW/iZN1CVdu33DzJ7FN1VTGyezr4UsH/TSz5zo0qO3
CE+G61Dd9/t03VnRqE75KBtLN7XIV9PIkkTrV/ecso64KQm00csx5m0yo3Dz
t4iQXF+QD9VrIwtr0yP0Gyi75tHm9ZlQZYY8vpP/IzJk4D/fZWAtCMSFnR07
jf3iMq/LOFbB/1L4EYOjGLIN4YDXaKTLjA1FyM85NQkLQt0QLxtkQcW1peqw
ri4am0biD9cIwSggLv5ABlznt70bXX46ZtQ5rL/7vB9NjJ25Y7CCaFbMW1uA
QBZhIp5GW8zi0TPMTG/VTyY4hbKF0Q9WhCrsKk2OdcSEqz74zmltXeIE6SrV
MhJQir0L9OTl4moPt5c2i8GyeWdWwiZzQGItgM90Fo9zXqyKoKZZbXfWTfj3
38oxYOlnNsvVurH4omR+NYaPsRXQ+khCDrQDL83SjL8cBnhWSd/gudZuTC55
axexrYAVreUnqbc6sAh16puiUB/nNqdnVFhBR1cVrEMHU5EkSibwY3hrtveC
QQ5cndHuAApxodPaWPMzsNBUosTeZmuyfGrxFV6gfjxzl4t6T4Gj0DfXWOmn
DSwDZ8aXclpq07531WsgcNFZ8f9IDcKlET6MRTmtvtClg9dGD8slYhxJYgcF
N5gd/x4kHjtsYm8zYF1htvWnqJ1gljvp+4++3zMW1+Cbgx5D9Mq5VTSqtdW0
fG5U/F4OHX9JNDrhz0F0K5vmzldztNHfLA4yOOfFoFxdKTtzjRwxkEvAraFN
Kc2VErkfj483geLR1drHcnsH3IMS+z9TdDKMUT3IxJHqoClP9Uwse/oQFjvP
two35BtzxRkoAIfs+706S5w/OJMe/cpI2iJmXtJvcGR2yNybMbJMhfXgN3rJ
SW2LB1XKSDPe2CHMcADT4zrvpxud07xR+MVi38OxZkgiwygS1r/7GIzUZxKS
uhJA6BzuCmbIxQBUX4Vo5BthVbMQdIJbqv2+DDqGAApCmCufTMZxzXrv5AT2
eTkS/rhhIPjAiCrm9bo0V/qREdacRg7388FvqH2LAFPMnFRNIyqwS/a9ZJNh
zoQRBqRzCXNbmUbSPlH7aj2N4E3L7cLYwwkk3ee0q/dooT2huuINGTNUwy3H
lAd2eWVnLWCXDI/7Pm8j+3+WtiWSqm8Uf44nNEz7gZVYPTScJmc9qp7IrZdQ
mG94f9l8AeaYA4pMlETMXXb8lc6RkpE0N4bGbp7nQBg/7oZ3qBQhv/3DcdXG
X2vWklt5LB+Or1P+xAdVlRr3947XoehDrZEPqQj0GXdxwCzkldmWaNwiGzv6
DP0oxjz6cvSGBg2MzauHIpjdY+8x9rln907YrQd6UaYYIldk9hzSrjOV4h/X
NYyNVTOUMOd2wruAwMr7m/cUKZIBhn6UmuP4DRBzweJcnPp4gLj1G0Q+kZf/
x3LsEqa0Q9MqlWCX0WDNoP8w+i6miE5Pnt/aXOQr74FVk2X4UvdjSrHtNvTH
8vqLXakAYAxALas4Dwx1Sbf+UvpI03noIfcRU9zOrd8j3nc7oTsymOYaomMd
32nrKZ1HGcLYZ9i26fHNG0Jqw9klMG/Qr0p3VPwYdTIB6D9i1e4iPE28JWAQ
aaaABiDQ1X+q+WOUWT+wWuGH4j8LqQFjt3N5W+pDXrocSZnlwk3ykGpGvjl5
GIB5m2q1kagOcXWh2Mut5gM+1xQd5STV+OebekmWrmU5GT33+OSk0hir7H4X
idKwyd/bHdgYLqS//9VGax683KRw/UUDsV34QuZ0p/fbEvFzaxIDPAPSqbbr
UsqydRT08TNlwvnhM4cgd8JJwVC6vdnpOnat8jzmJ7kflZT9G3zHUEIuL2/T
3dq1zN+I4zupZr7XHb5pQj1V77rIB3ZRKPVHsHSvaf0mgWxwuwMhX8igRhhd
LtzC4H048VoiD4Pnthz8KwFLntVP2UCeXlunNW8ZKM4IJ8RU6pjd14cGsQ8k
Z4aAkWqh1Rc7rw1N4uCaNrUO4kour5Z8jphdJMiu8lAUJ0aZSL5vbYhz5V2L
YvYSYQxDkt2gSEhJgBfC7TH7CS1/fAymD5BEYlyI2jRV4saNlZ636HVjgHYB
bkB7FlfgIzhYnt+eSf03hRjS+uSZyDuDPo7CCG0XWrhQniM+o7kngbT93CB7
F2R28YXyjVoLwqF/A+I56JRcdgI1ECcsHUpzFFGwmK+gOMPHvvvSss7SVmlJ
hL9+NIGjVjZBOS/hXKSEydAh8GATXSoFFmOPXd/Qv6SKb1hoqx8IcIYNCrEN
EnVLTqLB4oL6YbHlqi2Xu0QQ36NaPmgdhx+sht3yl8jGPIL3/2C/x+GK+oMr
7EcD5Mrm6ITIgBU7y3Qy0JFxJpkbT46WBtiCN91so9E/bHhn6zH0AfsiUQQW
jOc+y4KvPT9AZAUYhQXCQ6lAkeH3rGmMcFYy85uD+oPH6K7oN25ZXIJzzIpO
JIt+8K3tktFeEBbcTYRRdczOnuK1zwvAvcbT7npck4Gcgk1yVy0FZ3HmqUhN
iTxz0AXCNDA66E9Zm4rKNSpnqmM/EP1EmiFasmZF5OS2fOid9Lz+7m0YsnLD
IAyy9vHlZWbB566hYmNm8e0/U2K9SqDK0sT70jDmY0YVnImOVr9ZKjLxWrad
SrHKnQNv+vqjHt+NnF/exnxxe5j5f6WkxHpjFfD7T4KU+4cKGsNrEASileVV
4Bx4ALr8xQTznpkEx160mMEgP/5UTJYfJM4YMZrk5T+prju8SogMOuzVGEF1
spqF6BCs0mcpv3xH7G5Z6ujfcNrDBJOF8cGHgSyFuEghEbPTMh0Qj/de8x7q
RXNEhXFLgPhDg7yBtHIvK/O6JvMEAOlkb93627ZwVa3N9lcpJfNYxul52J/L
G8MMokfZcYSbwi9SwqE6zjiou699/Geg1PpJoWLT29sotw21d6N9KMO3cgIo
k20Ndw/chXJgeLVr7Yyzkmv4QdDqXROjPDkKivjmyJKyaciAWuupetW9uroR
Y6/joAMd8h0DOemQszvnY5P+LTrn3J5l3UYpWVkwDbS8rXCXpZyxdwTWWJ0g
WWc2Yd+vr9hoMuGHftZRAzfc+2Vxy0jY8ME8qJh1hkzC4Xo06p0EkwB/859t
2Jy88JE02FrthOJWvLKEZARE+fDJxUy/MVOxlUYrx/uVysLaUkBecBhSk2tk
beL/1VmLdhd5Q2GuD3bM0XUGCYfy1BDIAk67wdHjR5czK9tao6qX/a81HEnN
As/nVWKH5yTnpgs4hbJEvoizpdljfcgqS9TC9TttHR0BSstaxpNuZ685jkcp
tuuLTlH430vS1/iamiyI7WnDVHXDOdMPR2eSaJqhftSRhSyKtE/z7JyIhmoi
4ULx8QlcC6GRk7G6TIpQivt24hMpUABAhVGoP/J3jvytxI4qtz3eSlKkNRHY
5Ey/XwPNfe53sOB3/rpExxc1zaBFrThiWxBrnrqJlT16GiL4Bo5w5QgblqXr
MoAOGb4btJm6P18c66ukq2gfKOAcOH3ZRQjNG6nUmgGKXNOS+9+XXm4MHM3x
djQtx/2tRV4e1gnP5tcubuR05F6x+0mbAYM/WLuAqHSov4IcCw5UA0Zs8Fak
Dr+I7hsC9YgaToQlmLL66idf4p1uLk9dr3FVu6jfMlzwnBnBirfbzAEzLiUA
E9IEuSllXjJWHg8JUeyfbjg4HCF1bq5moQ3Sq0Qb+FDFTeRppIVgtfd0V5oA
e5UY7vuNuP+XgKnQsZBEvJSBnDhKew3f3d/EF6Xq9vU6tARZbft6CFWpz7FA
XghHuhWbuOfjsIDsoyvMjAKr/C0ySmLQdVTVcd02ct+0JQraqay6crpor1AW
nE/rk8sB4Waz0S+pMzMDxeyfCFznxgy6ghvEQZqFzB7hd0KjyzlHCFxdppQf
iMheRGQtRHZDIqz+y32mIAb19Plt6kzZQmtNQOmqt2R+gEtbf9N2LhaY6lch
KiRL8RA/Ra2dlGZsc2UH02gxFHFZMpJOW+iF3Z3Y1UdE6tB4ufsXme4QJutP
Qu/RO4FuE59ZsVqYpGzw+gQTxvgMp45HaE3yoRxDq/WsbomESIBtQJhzMRyX
NILWZUmPeculnVHg4NuzXcxn9Knc3+lkAgo5oFD7DZjDaQtfNSIxYsJ+Wbof
R3zJsRudLF9q22WfewQlSjHAAdXihEFT9lWoQ/YDpaAwEnIvDL7qdDad0iK+
VcqIJCTW9XL3pzgcupodRxd2v9cF49/FOWZ6DWoYqTEH1LHdIFADWw3Ab7iH
3FvvqAJre27g1XyRf8YBRsj2GaVpiEqnQJeyw22AHbEk3SGSaBATHtV0VcxS
8n5oRo3tyEmrtBx8AjMjGg/eVsAQRo885AtYyN9KCOf8+dhY40r3+SSlcghA
kQ/vT8VH5ybBJl8JUeT2wVXxn40ICVW5LMgMAoRZF5dzecIyAop7X25UFmuX
MfMYaJSLXJPFulieRnkIZmmEf4L8ItG7A117L/TJsZEjvm27glE27SFc7g5Y
2GRhWuaxMQwlKe/aOWCG3n4SvtEOkvepsngax+L5mmzXiDgHHdnVEmd9YT5c
Eb+oXaYhprBHGGLf3g6+MZkEDMZfSYpCFi4y8KF8HB2HgX4Qj085400O+9uC
JtQ6oWmXnSzG4tlibi532RCColdZJXRdN/YduFUpuomeZJGEUNPwevuu3n4e
41Cq+U3Df1g78lVOqqdrSNSL6+1q0WxRNU9Mnx1ZMyklHzyIncBhs/YbXNNi
FrMtgePwSI4DoN98Uz8gLhHFCSY4/a4D/VETN3gEDX73otUmRfvQ8imfpA5p
stmmQXZo8yYnKBB8QY9ye2PrYQT8v4R6zaYpVoIPWf4HPi45SJEQ8O+JrRga
i+CFrY5AY/J4B36IPzy4zzhkAzf1RKzftwqWeoqwlt+nYPv2ZPyL6ALhjcJb
1uE/EFgXuxWjRNmld0ycdxlh6kam1zVt7n48GIsZaJJ9mzCknKDMWSeClV/+
zgoTExIco3KYSkHY/lhRObk4cPnBMK9MTSnPeS+zd/GR+SO2OvIda2s4/9m7
Zs6mQ1eNTpmuRwizVA9mk1aNBM0GEfgn2o0bOoeG0S9peFtHLyA7rmG/Jiep
rtJaNvavx1USi7/YTAye3yTMtlqOKiukhtMb7TgoJE6JaBfJJCJXXi8dqNqz
a2rob+klF3tySb9BgsoZTFFl251DUDGzja2HDkKIuFJGteCKHDVKuf+DQgZi
/50Cr5hwsjkwkVtluScb/kC2zxSD+/ZyRRAplHzexcs1Ry7cpfAYwlcWr2yV
zVs2pnotK7NYxzzGeSXSni9vkwW0lrcd2/wQbdqiZLjIweTqYDioYaVWExxk
Hdzhk8YoswYp7+zHcfuewV4pvFyr/R6NIE2cSz+Or6Mc3GjjwipHd7Xdi7yq
jLAV0TVULLsbwhTKftSnU0GZ5r+VTy+Bdl2arSi1KIq6YeFb4ECxw0B8eCp/
zGgD8Wu9dHhb6tT0888pEpoGT3L7mIKi6X0DK/nkEq3krQqS30n9wJ6Xq2Vy
LEHV4AAlGJO7oLKQEn8w7DdAwde8QcFjjaZrDuiStcG65gI9I6/EXmNxdNze
zFVzB2w6pC3y2OEHWjSI42bXXlhJR69I43V9oFSHXZ4BxN4fQkzjtsFwq7hZ
fOVM+1u6G/edzDF8+Z5c41deYnes4ymjdZ+vtnfRmwUnU5Rs4qsUs3SpOa5p
WYCoJLDfKXNRwEHlYxRBRHS3swqCDDs2Vvaych0V3RofVioYVeO92Y2XLvsD
qHqGdWyVo1SCoSkvIspj8RiBieqfsKMOlnHdZohDL8wpil1AALOaBc5nctQx
2PBEiOrm7WyqTKb8GR73FiqRn9TvAnMnF1ErG9j2B/tS/WVQ/Hk+ylSqwfOz
12VbD8QM9gd3yreSMpP3ordT1TsKvwXkFq7A4ew/0TerPaCtgjdKKJDLZV8R
j4RMOIFhdYp8fIH7ZAWhWlAu8QRBE+WiDPZHrQlRSqkuVakXiPnkNQv2N7yM
RwzVdox6DJMmv7lCRrkAEso8DfYrFtG6O0ZvHz8OnB4ycl0Vy65fUH2ArGvZ
mAbP3QWHNC+zpKfgrUZ7UW4fSz0cHYWiTp0XvgV4sUSaNk6c9AeebZ2HjuH/
LecFTn22LhQBS9OUUzaGXnTzwunQBPLNEIKfcOqO9+1mpe1gvBg96B+Zdk9k
l0BA/IVYFCV3D4wst4Y1GEKfyNsF62AUNsKduOXeeTDjdWqV2LaZCaa+hAl4
Ou/km18TjVmBMtRYV65yBSMGwCXovg0J54rkwC7PBF+D2+ECPHa5A5TJrBur
QOZ5TbiiVatdKjMA1/UwT6VFBqxNh74oq728Wp6fDggFTb7bt342ALfGTiE5
zDzKoW1d7Nu6t+J0bGKoie/0c7u3rIGRxH4tkzf3hq7g4x6n9LCA2rF6Unr3
POxEDPfejrzd9ZLMOBaZgHJQVS9VkYDjsm9Nt0ZnoxbkhzRggmoHmHR8HtsZ
dfmeVH9NbdUo4N6NhSkdL6lkgx0rJlR8jQpSPt8jEgqNJgZd5HFCrZ9Jc9s/
lNsd+0MrEn/6x7k382lXKBRLYursXpKXlDzWWTxtD1YmdCwayGMDvMY00MV7
10XcVKz9gwZBBXDcxcC3Uy0Wr6LTYylztuqd+a895GN9G1uPFxH4M3wNwicz
aYjG/YwLQGHNOFROexdiIcFD6e+L0zKuyrM5a5VOC9DMko9cp/PpqRb5g3fQ
lLtyDbVSfp5C90EANEbtQ7I7bFN5B3iKpB2clYbzIugXMbqFh4nY3eLqdQun
xYpzByjz1RMfzkML0pd8LTH2M3vyxaP1H358ql4EJ2Trl404zRphdjaxVfBs
fXA4Mz1G1IS+EmMKam7+dPMJuNl7lipB2EUJzJQG7Ewgc1geQh7Roj7DCjc+
jzAjJWYXIrHZ4q1j5kHNNSpz6bnxBr+De7IyoX5+XhwSaAvVpUiy6vn2IGne
Lret0knRsX9QXRIrVtNnMIOilDJwVBOzvKKeR0YwjriO1A5ry0Tn3YRK9dXi
RObMtFvuYMm/wL7SWP8lPytuLb05K0stmNwcBgD6kFpQE5dGg/zZFjozfeHQ
/AEc5UEc6wK+IjupYi9gbB/uCY/EuDC+WTLPwJxRKBe+jxK8Nbp2R3jgVyR+
N8tiQ8L9vjSP/KRTWqZ/K3XeYvVYDftxmnltIvETzSdfabshi6TPNG/6Eoam
xSbwqqVSyWwvRtnrNX2QJ9aTK4MF5gsGNpzP9814sXRjzJewjrATBTiZyviF
sJLxvy9fOoEF1Wp3a1et/q74uV7zcvVHxBlTN4w7uj3i5IXWyUtj4WbsyT0M
1/y2XlKkY8i5RJIbRt9Sm9hcUuW4e/v3Lo/nWBU2jBK0za2USSFxpi5AA4Ls
rn1xYXsFQKv6tXOi711SeN2JprTJN22nTe1lQdfSFy+Nvr1Gc1qHmPA2dkkg
rQwdi9FyXtQBONpghKxVmc1MxbGiYTsj5PUZUbrElN1PG0Jb2+JB+zYViF0q
0Jh+VeltwczYlZDsBV5tEhzLSADpYBUNfe28wQsSj0bemLriJNxrdCnSY1Rb
GtDva2XbHq9uH9eUihbWB1lVPWJzULmng66eO99higiFIwYOjQm1z5Diysoh
ITsr1e5RDuIkJhxGdkybw5Hx+mgRAQ74M9fIayOT7w7w7QCy8cB9YtRXUf/E
eTZo0GvAZn1q6MZMv+ONutaI+RC01yYmtjRX4fRraetwv+IXUueDOu69+U9P
itzlPph9m114cT1t3KzToIy1Vox2v92LKrwFongoWDEgxg4gh2EZBRp/5OcG
N9QK+71qAqIjgHpxgpE2naDAG5kgVWsGsbTdS+OekBD1zIWNf5YLec7Hl0+0
uNRUB+wkCwyQTDrExvy/F4LywKSszdzgCyWcEzTQuQDiD9qr9CrCeM0gl+ZM
T0WCBqWa/OI0wGdiWSV58mTHQ9lq/d4jKSct6jPNpbQZ1BUUgwAdiL7nmYaI
MOdQIUII2b7SM3FM01xSb5m/eA9Go8Ge3pJdetXjcwRsb/ojX7ljv4TCmW2W
47xArgPtEFgEJgxvnyLDrfb0hpESqhaR3BbyvZdXFM/rf1m3cpHhyGW4oqI1
ice70ccleGHC1Lvh0lwpLisSr8Ya0uVcoMHbKBmITGNsDvwvl5q1r5Rsn9Zd
3QT4ciJCC89ApensYs2Ut+4UjWHKohQ0400RnMOCABqFih8k0Yz9+FmYzx/w
PRkqy2ThRMy1QVBh8omeGTfaO3QSmd6PoYJtmUVVNXmAEX4exiX7HwUSofQO
G2pUZGM56cW1BDvTQ2iMpwxXwQTNgXqODBmpz6XrWaZYdZAlgYi4q/nvVGh3
OdiCNk96NYvP1HajJgs5AGeo5Eb79trdJ74vmJyFTCQ7L49nGaosAjuJF73F
Y6G2fh0dlKzNHQfkXgxj2ZGUaJTpMyfdUoNvzwUAFCQfRYKsdOt6Hx4Jd2+F
nnGe++oPZuHrHn2Um6G7MNb6E6oSDZom+ck8cUPXuaJ9w7sl6rcjd/XVUHeM
wGDlGz29/SoCEIOmzpnF9vNncSrA5T6pJfSauiuMyfwsBSfBMagFmcjiwfn/
tf+ZkLWfXMujUJTbNH624P2vh6TbsDFUP40f2KCWOEZy49gNj0Bo3iuXLeTI
TCia6wkWQlsqZ6iRJh3KHalhGtw/UO8ENvmqkkzadTN+8UN3LOHld/EI6dIj
NWxb+kDi+euikp04OEsDNTal6w1iMs8opQZDYKWpVABZzA9cqpMwlU2nR6BL
sihkjvpzlkWvwEosbDFBkFa4Xe5t8amcnlpFZSGPUI9Af3a7xCMcGYBwaPMa
pe3Z4AxpYaE2MSr6WjqV087S8IXrdFMrWDXkQTA2fB4AsBLASj9J8aJjY/Xu
2DSLvjJxUmTN/gy9GGp+UPf7DkRmEiZZ9T02D5CUq9dv/tb840vvooHJpTcW
Jsc29gxELbRUb6vmORjZDcA5RhMVi3YNiQN/9AlpsyTjHrVfI8iZDlzEoyZZ
UkbNPVjV6jHEbpb9+nUPZGFTtn/n5s5TAM5cU+YwWlAocNc5Zre1ls4iBu5g
JV14J5/RRJ+oGfyqpiHVLlkUJecjkBzZRtYEAWzzjDEBIPi5Kwzuo20vw7qj
H8bNMx9hLwgN8Gbdl6lhpdvIfiLRODFW8x3mFUR8zLohWOe4mwiz5WupIIWg
hOtIUthlRAW2eOv7knq9BNFCeTSGS7vHMOzfd5CAUpzLxnwy2wJJvYtIflVi
2ynJTMU+zwUorqte2TX+ZSfsMcFc4luOMG1ZlwmK1JPVi2yI7hWyl6f8MJ7p
5qnZl2drEgbhnDQqCGKwXENHg6Qx96tsQYnhRJLx/qoeVj1vogPB7/rAGg+M
wTAZTcAIZ/XR6HqQaKCKRSq6QUlVTcNDAZN5hbksOGbr+Os5uk1pm711lDFZ
ME4smdRv04UEt7FVHgAJi1yD7YMuFkK0mGSoyh287i9bd+U8LxeHCcOo2ioA
XQUJTVq30pt5SiFlIUQr9L5eIzbbFbZQCRwzG4aH1k7xHW8wUc/hJvGJ1uN/
eoMXrUYr5pMUqa7vrRZt5C5LatbmVOgGemkE1v11jUrjBnTtS6FtewIALn1B
sXpOmPJGaRZ0AO91H0m7Pe/BlMxJ5HiF9AnZ/FZ6CwB91V2UAMp74hctjUXe
R/F0sJ/dgEGShH4ePN2SKr7gnwL86rgjiOtCtsECJCyCkNDIEW6494FXe1VO
bU9Mi6nGl/JVxSfbhRT0jAdYkHsnfip416Rh/1EJ65/72Cpl6HHf8pxnXrM8
OH94gSFkmYhE6qzBkVivWgtGH1f59fl3rRPYrjKlKB7Rf7VQ0dJZmRCexMA7
NGD4FgG9tXyhslDIOcFCftranvUYzRVYyDU0UEgJf8bEj+qzcUAgg0lSye9A
KFCPEcED4Ruo7qR7/XLuI8o/k383v4APW5M/v2fLe/oMyx9IiiaAlaXHGnaG
RjxwNcjxA6k1/C/JOD2C/+P/01w+XCK9IcSaCqT0WZE4CtscWnBvJQupXREe
I3Kmy8L81PknuKoqtRXJDoVHr4UYWsrw+NfempkFp+KPfnXFBrNvS/qh3yDI
jMNjexEni4cHAc2yd+wwieycE69pi+CBmpKsnB5dKliMvBRqkbP23+8X1o5o
ft81Ck9JpqkdbhWQaQOVvyompDatniaar+PqsjxIIlP2uqUfKypjYlD3Xykh
l4u7Sfhu/TxrHNWQ3dVIF0bL3lzVpf/n1K7hTDJv+xDIqb9Sh0uvgPE5uBLV
Q/fvJjuOazu7wDO/liRg0SKAuOPNR96OQP7m3nzTS+uulQDRFR6fti+jP+kX
E2qP9o8KXAA7A6TEO3F5Lysf1M7TyzH3pqC9YtltYbAZLIVS1ekuMdJ53dUN
hWY6zoFpRcMnsqzORIYQfQ9IWwzMGxjM/fdZ0xE5luXfDOdHh3O7ckiSRFak
zCJDit9plEC7VoByvapDAyzdIw2g/iJm4yH+GjZ3FxqJiTCcPCZ6wd5Lp05e
2Hd46gYgJnWxJzQtJwJeH9qd501UzzX8J9BOj/VdUgSjQ2OHnIrMyc9I/+5D
WDb4BE/+AledmVN5l5azcS8xIEuC5aUfLdZ8T/Dc2kjf3eCs95AHNdrSb5Ii
3iDlICdD6zhLk2GCSMjE21u08TrGF6QuNZTsHT6ZtnwGNv+5KVbzPLVwOhGU
zVIlF1kZ3R3FjldUPIYiWOrG9mGb8+KCU5QbA6r1ooUFSnNNTmLCcVKLVOX6
SbRVtJSR8fsycdjj3w1iOXiDpD0OAfqMG0BKw9X8BaJltB7HTU1j1nQbCbF4
f9ltL3y7Dun+ebixFrtaK9bxmqN2Edq32+4AN3GeEtNeItAAlFYJxXsJpJNF
vzieOb0t19l3SdZGf0rT1PTiOnZPLBP5383hYMLfLoDAfTmIuLWhKrQP+NtD
HaAAWa0AEr0nZlMrFxh50lGx4RPfncGyQLQ5lOF8VuXgesgWxpb4zWILHV6h
SstLR8iE7hI8EKwUI04bAt1pvZ6PDQH6Ztu7VCmer4Dkl6PgwnUl0aLB+IBc
rNSsEc1YtFL2W8/D5U8j2x/TU6TuisB56kfF8aIt9Bf/uVaZc7qPIbxN9PUk
2bugxuBTBkep//nVT53hYCS5o3JI4JpKAIdZuiLmhH0bwSLfhJFL6BCSW5VG
Cos3rNSJxlFvvcz/7YqLtch9psZMjD2kk6avD5y8bv4RKEWKnfg0sv28XIYZ
TBV/ARhFfFwVwH+FxWXwHCrm3cT25dMeqQmxrQT+yaKgFMG5M88M7zQsDR6H
DXjIxZd4pqKa+2YZ66asMRqL7yKPeG12F+R2er1B0Wrp3JVQ3tiygE5boolc
zBbGq5XIgUs7h7h0VIMvS5kneGRHZER35OP2Qd8N//QEN4oDoZhQr68teQJB
67rWhms+bgV11B90AB8NQSoOgQ29/zW4wqm7qWSaockv+C+4sUJGnWJDSybH
aRScvQgEYShJP2mPydBzksZZVQdZ78weUFgi5qNgb3WjoRe/X9v3ZIlGSsJ+
5lXsbw0In3tgTnEQgpfHxIFGsmprKwRq9/e30NQfgk/J29Sl/kG7X2x4LMgH
5qtHpy6zHjSX/TNB3S4kFW6C2AN17sF/7NE5au5IyAuZO/akhMzFEXL6CPKS
caxuARsiujX7/Hn4TSjXwGjQ/NY/0o/L3RCGnzX5PXxQf+hcWrFmySJ0LUqP
Vcwqil8CTTkIeT3tMROfA8Iphrx1WzLyGyHwMZ4oV9BEyLMz4uEEtSlT/cEN
Tt2hytUGh4zaqvEhBp7P9rZTUt/+SVPPmdYHCp9ymY/svXwp6U/jn/ohd8cq
Q5LOQuA+d97CxuG3qfDBCaoTj+8mAIPZm7g6b/dTlGD7qrCk7Ha1+kpUbqCh
oprSGRzwlfbp/uU2TD4uAoFtQVasefdcllfFp1lAvOABDEt4aV6qeHyXKY7C
Itf/6bGVvLa7XpFJ+1CwDbZ3y8cPbBrC7C4zCENS4XCQc0Z8+kG1w9Ugrh+y
IRNm5ex8lYkZYP9gSQUAhjIy61q4ZiREBO2Dv0cSyOJ+l4ezvGwsBULXxWRH
RzP1vuoJuwdYhmRGgcBbhEasbNwqFfBwjuRJf7NAFaERe+l+PuYkpr2v7YE8
Wcm0KaEF8m+RMBGrtoQevMtOzNLQ4iSvIyz8O8oKBuZgRXeNFxJbGN1hH66T
pwemJ7DwmycHG5h/HonNzYGJJNpDjnT2QQs5IuQQPQeoIFTfw1BgDWq6agRa
WI5SC8MCUuxbErosQdN2t7fnRvo0YUbbqOQvcy1/jrdVhS4W2W/qdHJ58kqd
WZV3PdV1zNTG2RAAp3tYcCNQ+d5Cit2T5Z8tkuFYlv0lDUMhu+lxxPky+PYe
RleHvsSrLjv+orCpmDMS8Jw57lVbB83SiWaP7+z2FOcw3Bugho7wdReqeHMT
rstAe8yIbQO5UKYrjTak4Fjx2lQsdoj29fvWOVgxlpuLeOEqTG6DwVvX9DBI
bAq3bytY7gr1qy96/czbhKptBYWxTUmHBwtYe7p8Shee+IPn0kER94Fx5itP
qXbtY8T85QMJZ7CkktohfVmGkWc93oVtjUfzacC4WIjIY8BWMfkmMhv2Grn9
42bYu6egGCboOib5VsC0qV0dZ5Oqq1WSS23B3AjYwBSMefGYkJf/GoxZiMEk
E7VSHWWLKc7IYBx9PqpCf0mLABCsw+qoZNxBcauit597W0tffAddiPJXRG5u
KjE1fVZ4P68KnmURqlRYW+gpkwt+EIC5cH0dC/FLCLIdeQwvOyPh7RR9S6uO
wbKzRf7ua3zT1JOCqIlIaLoZrb0Rod1XEJ6KwLMoI0a2NqwagP+RJcjAfbUM
qkJPYSDVwqALO0V1Rxp4zxWmFFwcN4OafjQNx977bX+J8rGTiRddknPDq0AP
HsnNDWJe7S7PdBeYWqDcqNU1K9OdV1Ld7tb+GmohUC5XXyCKe190EnenUwj5
31HouSgKjv22dnD3vqjtdFrnSum0ZstUB2xfV9l6olKyxcREea+lEO+HwsPY
p1kWKymymT7Agg/VLyeZHzNYoFLdIEZ3W26VC7f+nNWmXednLf93RY84FQ4x
6I5lSb8hA4E0yqJr8G09WbMRzfYWrgMzwQJBuMyjXUKoWK6jzEIxhvWzD84G
llK7S3gCRC7vkPXPVzY6OlRK+IorQLaK2RzR8mxZ9owIB6/vBYlX2ckW7kGT
3NO5D39yHrl2LD3wEcJLxCEYC23uwT1CQ3RIElnl7ksDisbzkuE4wP5tAwyX
yJKZK+aLYeczKnXehR75s6+dcsor3S7VJ6q0exxoURE9Gipt49nzh1IoyMje
i+i/NYCKttIMFo2/T6f6oYx/8wo4cJpHjs13zM+gbxbVx1rg8te8iZGRXA+7
sqWe0yDa+zh7BWOLo7fpU0OE+EPlFye4CXcMYknT42UI5bmv7mYfkyfwW8Dm
J1QREuekapd+Tta2tk64ribCgNduSUkBfyxiAoujHtUQUC5PHmKvjw2sADpI
9uRdsb/1ZPXH1Acn//X+z9KyvWSRgrIB0MuQ+ELMXluGspTDRQVFQ9vEFtwJ
+HaCUi2PbZjkbKJGsKkZdsB+9Jrf5MO7K4F3MOy5bqf3+vahC2C66sGWiqQB
E0lKSjP71dkx5wwQlqlCuurSaKYZnVg+HGdPMsaAMOMlHxVLtYqHolZVrGB1
Yx3UxnqucrsGltjbh3St7uRU7ZA3ruOhGvB0HxiAxgZj75GcoljyIFatAMv/
8gy8ABKiDZZts9rdN3YHOGlcUNdoc3n9ldLJUw92Iedl3AxHNhW3QpZ5ghYw
UGmLZu6fEsBXN7Argb1m6JpAtm5rfmXLLaHds1kMFSMrPKcbnxKcaeI01BMI
FuA/TAT/J9QBCowT1+1PXoSj58SHBp2unz1QKKkKTp2KNZtxsX/cR8xTFwpW
yG8WKz0q/bBqr9tfn9lrpAzzX1lmQUKXUoR/LusnuZT10oPF2JUDxPs6vQuv
kvXLB1Xgz5k0qW3b8WIFot73hCe7oD/DHf8Lh6U4el1B+w6jsXFMacxLlTxZ
1adCy7pz0f5+500Cj3Jye1bLUr4D94yAMeE0k/go3GIWjh8li9VQ3h+V7Mhr
yTQG3dQHPZZGJ9KwmrX/gK1vbG1uBOTCDOXi9T4n5h+B2FlNuztb4ZKv5F9i
O5jecUGRrtj4Kb5xFSjcfisQn0xExiTsYrik4XQePccteXzTbqOFgyEWWu9A
cGuSiokXoUxzApSRqIxSPebxsqRivOgB1wSmHNwbt7zkFKOwRV7mXl1sX0z2
zf7mwC97euyPc8/rWpefLRJfXc/Bdv9mIh66HrKn1Q9MxS9LgCQC+UmJWwam
KnA980El3bcGCD4ivpxUCQgDWI1ObrV4hpskL0LSVGXG+lHcDqdI+360WTmA
f44rKN0MUvNnaomVBCh//l+9GQc0xH+GZKVB3b7X6ENyw8k5Ky8OkFi7iahp
mmi8WIZsCmgET+hUYoNo687E/bYtnsBu6POAoPQOf5CzzES7ISk5UGsc3aSw
StdrFJoJcqcCe5iGK9s+NnqxQnmESHhOxW19aQo6ft7McjZO9Swotjcbx1K4
JfU154o8KYp5VUx0h3koNjB21kGP/sEbFOG7EbqRqFBzak1X7jriYcKh5z6s
N7ks4ynpAqs/h4Gu1mxYTSr4k11kRufaZuVwmN8HQxE1N++psi1SGtI6b89l
7psqd/NfN8RrBSw+Dz2Tj2ZDgMOiK8y4ZdwFHrV7OL4dgFD9xQgMWTuUBW03
lysDZmmKUVKCjN1uvLBcBSt1lFigJkSURiiAp6NcvpKWvWS0joyc7i9SkT7G
z+P7lzDXxBZZhniZo+q1YsBYwBdQGtXFl9fc27Um0VKXmYYExejKJfVEjwwn
pHdaHmuTUvODqumK/ZFgWGT8+1fyeXgFeRhoCPm3fpE1SMYpuiOhOM9R8Lg5
EWbDA9G/30jGrubRAfNA8lvoVoYtEn/dOfYAtL0N+ZYMthThzLhRvS/dFG+w
jRDNaJ5m18L1q3OSMx9uh5YK+R5ch5hZSkqFEZqALB4XyQ5dtGvEvZE/qBJl
Nl8W63gwFEFQBGUgkN3xgYUPykAiKMRdE2tsMc8Zt/1PIYUmGyJPgwFQFE6p
6tnSWvxoiqqQFZmJ7o7/vJqUVrsQc8zQgt+KAmMKJaod9NppPTC5y8Ph1Z30
0gLhI+ryI2RUUhuDGLve7KYo65PPEkxZrW/mwzgktcCfwD+B4z0S7PHcKi7w
Zaib0iZrZoik8BhlgI61Gb0wdnRf5qNAZduavbP7jSURjZc4itCBG4n+9aL0
65gykXnw7qolxtwT720UhOPlaaC41f++ulQ3T1ssj49LpiAAb0RCCVeRd99/
hY3ndeIAEPDBpAlYk8j2BxGAR/8eGEf7YLvBsxnHuYFVgqpSOaJbvOLTdaKR
ziov7Z9qUYFdrDdaWVpYD/nNzjMrW2YhFaIgRsuwizktuGBX9BTWvYllJYSa
W1Xs4r0NpJ+kKfEDiyFND3UWzSXuL069bc+R50K6gx33dRcdhYlcM5wvh1U6
zrxplDZs7Z3/Gya0PGlc5aePXVTCmMB0woDX2ocIFMYs/NcT27vWWNPtckbv
2rU0EdBR9FzmTckT06r7zI0IbcepYuqWZxrDr/c4kzguIUcR6FlVamV7b6LU
S7SMbWd3ECArlXIrItbcUDsuwVSprlrjpOAlHZ0BOds29zlz2mPwE15P02Aa
YEIXowrtfRNMWdjtQtwvkg50zvVQ4ac+2TDG5uvVuRr3YcxYytc8iewAkROw
YZMgNSqgMeNJSitOv2HD/FK30i3FS9/vrVdcFswC0PivCER6VahPvWAHnd6X
VmhQcwK6FafU8GhCgG/ucVxi0NuKoaSwB9W0CN63bMSgcpUFKjgM2p+XWHvc
h83iwc0FVmWywPW/7mTLdAw+ZS2c94D/n5Vy1uaFvPO7Tv/jktQViqa/VJad
mjdeXHKPsRoZJBp+vXXkOLCtWP1xR3/2l1IIfch1IqcGSWyCboiTpmG2q2b3
JIupdWIg9X7UNg6VP7q4ra2c6HDtdh4Dv0SGPUtDiU/f0kn5R0b5GU6/AnFP
mI/D9rr48eOAmq7MNdLby0e4O7J2Pdz2jICAqNwH2b8K/zew1TmfWqBU5YSI
Sm8DLF79iVK8Lbq7emAqTCpfN54my4h1QI1e+2TTU5T7u9OOHR9Agu6pdRKP
L9MtrPYHlrO0DuANPmGjHwQkoBLQzSNnhZY8jqgb3BC71PBX0V0hMKL1k4xm
UDgXDO3hpiaIf+5pHyijQzh39evUXURwKwuGFGwFjhNohVgpfxffW5UR0inY
K1X1gWDYsrb1pqPMMWUIekMrteKWbf9iu50mXDIeB0Vu9hCJ/wlV0a+A2sam
2bL+JP3TsKeVlz+U7IKzSUBSEV+k5UGlYyvU6gqcnBf2x3da+YUiD+J4YRCr
YDPj8hakCcuwynrppLhdG9Ybsd1S1lZ2qogA7ClUIa/d94VwjAQXLFPBHm55
kw6Y/pEWl3KVRNknaJGf3nts//n0HyDmotk6FSzsbti40ttQjAvPOinWS3Ti
p2+Y8RTTJwmXm3guJUPgkoJBcn6Jl1zwLPRh0p+R64w9vuQQeKY7ek18n+Yx
mis4e6FaYkZEZxQnQhHUwoQzrB8adRqZGKKPz1ZaGgBnApf44GZvv+cCZujK
ZMfISb5OdDgC/iLp80gHc7tBbpkDPBBq4wtu/sNY+BKTXHR+X9TuWrDmnb0N
As2340d+ZxPP4rF1UWgfFoewZAQMOcOok8TgifVcjbwYDtFeoWD9/TFbBNWE
iF3GADMya+oULO5VJNHsk95/eDhiDPQgrf8K3e1wn99XYppXLmQR+ohqMGHj
DotB13kWdeC63UD2Vb+KFJrdM0cHcnJNuKWI3RV+dSz1CBrbxDmX3xbuqvBo
bqaR5sgmtbCMqHpfC0DwIz3Wb9WCGDnmVb3ZtKPve+a8u/ihqVCcmC3G1xub
YkQh45dfZiIbTLRDubR8qGsTe/XHNYBLnf4P4jBt1i3ALX64JRI+93GX9Q18
GCwm7zwl36SJ5HaUsFYvRkLh21MC+KKW4CSgUpz2INvbReZrxn59xk6FiPnW
q+0jrjaAHycrF+oraLO0whs2QuOnQhexFZbHbiglsxCxv7QUBBWK22JxzAV+
zfWVjHXgScR988HbWEDpUAKhKUx+Pa2Kazos9iuTfRLyZmRrAPZQmkH/H91v
T2AOJhAlT2gvYhcU7hntmdA07BHY1WiL+uFgMmQJH4ip/nVmZLM81FG7ymZj
6uQFHWoh37p0til26MtCLvnjv9B9eJXc84q/sqkLoiXKbTIlnf2k6URpStSb
yxPaketJAkwJa6hHWDx9rCXXujJn/txxduvBgvwVdV1OH57AY9E28a8EkreO
1VhgvFTxg2VMY8KwWpf5aHcrIMS0qplRIChTFGgdIWi71Y3F/vCjHKVrgS2C
zI0MeygK25Sv7bsHvJ58qpVaxpe+OjjSkI185dTRsSYR3DqnnTbuljiRPt/V
CgLq74If2cFTALyrwyZ2hy1seO/vBSa552qUiyPqPaXS1qX41KqrZGaRgnQQ
10ia0ZlXjUMms3BwymoIUKPp61RivGxQE9ah3YLI6iwzd7Hzq2JnkdOqcLT7
nJP1oglmTFyqScKEW9Yrl4/pKf22smwr+8v/brT3BRGB8pIIQdj0z1tn3XvR
/m9SwzaDot+7Q7waMTz99KZ0FG+P6FFeH967miA2wuyABeMHsdqAoqzDlSmn
9j2MdJliVxLkx7JggmPNYjw+zsQSCHhjGpP7df5sXNJrG5VWzwcMfk9kalt0
IG0cAqumPfnPh4UzV5J0M4o4gVNXMz5eatRCR9qQXfHzYrpLJXB2BgqpIDVN
Fo5WsYmsEnPPzy6xyRqyOt4CTrDBOg9OMCP1L2VNH3GMGZNXS9OWH9/8bkXg
TMj79yvLOIpNo0wALK5gA5R9UAExoC4WC6LeZAsUYfXX+4+UAMxdLZzGYvOP
AfduR1yXL2BGww7B5xXtxQWlFsoqd2nUW9rkfxbNLYyTxIoqOovYRI5pHv9G
f4166lTzgxgPzFxvUatfRVvmysPgUbShUkurfkPMsPGN/BygLyOX4+rRYUoV
D6XPZiQqTcBE5zB07ksqkyp6yJWSB0wmEWrspWJo3oCvgBwXm82ovfwP6uCv
f/jFOBUgVLKoFFhdShKQQgAZnREgVeoQ4VhJ+0Ox7Puuyqeim5jQvgtuakN7
FSNdYR+xDbtK/JV7/LmcO+UKfzAxMyODy/mY7p0XnW63w4eKxl+Eri7NSUKh
6XZa9Xbf1f9XC7eyEDM+NfqnzcDnJwtf+LYXdECN4JHcO10XYOFITglQhkxJ
QeKdwPUIJcu1JYhbEUrZ26ro5U5g6KcypU2EJezSVXstZJmXOLiVWfo2lJLm
hlIXLQibFEyRRZ191dA8ROpc0CecXLApx0KfWBqFdGBFXsTQuM8+TOWMNcpr
BvzOs4qCDkPMJ3b3zqKux/B+ne6VdeqxO1hktQgUeaIj/Q5tbWlJQqp36WlL
j4xsCH6ngPT7VRZzlMlYCNU+p9kRwTBO1Cv4jrKtGRfrgcfLJyi7yhcoYIu0
0VZyEacYfJtZd71ZEm0Ku0Es0teWtQlDswr5RU+9JJ8BXwmgFILRy41Pj46z
XCRFBjcVvWNALMnWrXWWrW9TpmJFwFDUZ5mm77BHppWt1WBe9CQhIM2DR8o7
5drVMzZ83BZWVOdURoxK2waOpx5AlWa99j6X00kR4uglFsjBknqxu0yWxAlF
3XLdWFyEXf04Sxzm3gJg8TpFricgp/7wzxbt2TtYTc07LDw02fIKucthphMV
mvuBRb7s6F+vt3dT1bO/xXlfTu0sxgSQo2j9tMbBYWPAuujfgf42C0jMdjbZ
U5iUpqDlfOjWuvAmVBSw4XKGhK9DA1XPEhTXVPdgZc1PO1DFg9VYR7U7F+Nn
whT13r4EPyYU4B6Z48JpUJSExGUZbI2VxwR952Cc8fQtWZ1aKhOOjSsY0mHr
yW7B4JIz7AG12MFnYNnFqNu5Si4wSnKogJ9k7KVTNeQdb0oXcrnEyMvieDjw
AHaFAqIUmc0klP2lrLcJPgIxcaV0fi5H0DUs9ByEpLiZbF5tlLbhrZpNf7iL
GOuD8mtU9NfN6i0iH/BVrdhA6X/GSL5p8yRru9wOepYoFQxEIh0aWY/vJ6Xd
fv6s6odIGFsex1xSWGHYzNl/ry6PVoZ4lRXSTCNX2gHbXCN9xIkPU01mQc3k
6AhsRFTVYKVtbSFNSWt9dlZXG4PwyfQuPymGERkrjMaJpeuUT2DxFxgDXM2i
lIAvVntdugo2OeyI5CCJxLufV3WKcNoN4qgbMQ7OLaHpUWqTQr4QSfR/uTRB
7gtTjYwAAWDzCJ01PRxl7Fbu4z8g9steniTgmcfB4IBoX8ow+eT2DXyBs/eH
2qxCeYFYh2ddBctKKVZahW0sc+Hqks7rCF7ZRcfjxRB3+wY7xBc5x8L0+fAP
T2IZk0VAu/XueY4Qv6xLIrJp8degOKN2ly4q1MK4PoliqGYhZS8NTsSdNwe0
/d7Wz97dj3uG6UUMjhVn2nCbKcvD38C3io1474v166zIaoMNDlvokAUZtzEi
1PIIR9+TmY6+1Y5kDFigmLnoKT2bukrsFhhWVmIFdJOzX8F4IfGPqU9dBe+V
SQHbrMIjbSThLZsYX77SWj/9FcYt2KSoMky/66NwywlUQBpImJEor/nPHeyc
YsCmjVWpgdBCHIVgz7fE4EDi2RbRpB0PkPMM5Ld90Pv+PR38etesmPaCeuc4
EJBjbZ48nmVYFPy+f/37KxmmHcDiMHU6xTSrgq3ne9tYLJaPndHFfhAbO47N
X2LqmNTIsNYlNHKl2UMySyE2Mqv98c9LR5QMcwefcUybrB8/IljdQ/BXRXPd
QsT08rDcxjsDEYGqpcGBwbEt+S1ly3dvs3RH5H+Xe0Hly+TIebyRPcqxYp4f
SwHh2sk6cCllSbLO8u28Oxun0elHhjFbcYbpJQ1VOTYWahaU6qs+MnoPVfOL
TxIvAnRZLiX2kHdH1D57BnCaK78F+Ibr1DiQo9CkrmzeO6eFkMBP/DKepoQO
LUwiywPyhSAr2DoA82QaiBO14xSgAmri36VIkhpd4revxLaabbP27YRmK/3a
YCnwCYFce3z/FWWvQzq4kMIcmA+Bkstf8PXfqgq1uQ9Q4PIleSfMyDl9s6bf
RbNuxAh1IydAMha0z/VJKLNVyLegsUWSoOQ+9W/qmzKyDlw2nQW3crDFTOfp
YjccJcOLQsLyZBb7kSVXh8ynbxTMGe1sfGyrOgf72LIBQXLRgJ9G76c/U4FW
opZr/9ZTw+OizcnHcezHlDt49s/BCPHiAgKp4VGBNPZCaWTxaorlZT3EOPEY
hcJk/FE0jzAn7qDeUkcFjT/3L9S2KrKCgCp/w4z9MD3eNp1ZRWTdsjp0F3eo
en0ZCJRYKaSUAdboohAeE7k0B3kyvHBo6lWI1/37fjWlazPnGkX84ziY093i
oTcbJIhptcqwvuWRhVOwtQt/ZYcdkjR+uH7ocBgzHXKnK4AfxlGKf42DCfXZ
JsjRmDqQKc8018eSSZfH7+tm5txynsQMcB2jWxH0+et7QqSnzqDUk3uSeWi/
6mSFRocbt0zLs3soUZHNlD0T1rR9xo4qpsyTEm7/4hDXSjTSOcGBpjymmw70
ScNXdJHFSJUBlNMm/QHfcGzjcPug3QtPx7IS9wt5cMoryMRMFzoGU6wZlEMY
Qnjs38OztNi6LRELJ9nS6GNZw6wc5LeHLFNt8ufjfezfm4Zt1Ok0xO5+r0ub
JbO98XaErgmTJRcKYEflkqrwSFBgQJ/USAW5rIud4j6HYnzFF+NGGm4sGX8D
N96zOd8zX2EeH0x9Igbt/pnIiu1PGUI2pJP2o4J2bJ9zGMxUmryzc1yqFN+t
Cllh6GqWiMSvS8h8vriVeUHLqlLhIBAYgpKNp6BsMAA0eb1DvuTdIVmPThr1
0MBfGAl6tlS83Smrng7EAASIvIlB7k8QfEvEqMa9nQAPdAgMUco1I90VxWFt
E+MxQDiaZvavnF7KKfsQaqQBLHrRNq16SuXI9ZoJCEohwXr4i1P5qxT7MXVo
gnfdKzSndBx96/b8A/MCJwoPYGl8aegoRou4GjbrYFALGX9RM9tTQ5E7q2zq
Av1ijdXlJgbzGXU6liF0N0q6az6rJrTADIHxUBd1Oi3Vt6ME0jpwkBkDgulE
uL4/c+eh+mRsJAU47r9cs/8PR0zl9WVoA59tNi+R7AkFPzQxYf/1E9KzW52a
M5LqYzv/1DJt2/7ug+RMqVWLuDPZt11w+9lQO3SUxyPZle4RRFSPkYmpIo7h
J7LXiccM4ywdGcpr1LuiTAIFzP+0BErkzK66FEspubc48xLlNypt0LsZgsKx
xw+WmxI9lf4dKsmANgiuoqRdHdjXgpCrGi+4jnD2Zniocibz3V+UuCxusrmn
yN4VTwtfuo2g8K4A3kEO2qWnv6WlSLR7Kvfwy6BPnifntTSPgAOLXCev8s8l
/kUaVBCTJnd7dKWRfJbNstLyY7zLX+RM4Z92vXxj9dQakFlWwsexfOWOs8x1
RPwCed74i8C1ReWcypsgTMh7sj21TbChyz+a4ILCDJDxqvKFuj1vQWHYCrNt
zccjD+baNhrd6iQiCRNBlNwmiGTp9dOpq+PIKbQeWSJf4B/L9XkWRt2wCu2r
hsZ6zjjZmiCuNx9xfCnAi2vaYR9nN/QSltzNLguuFD5MTjAuJzW8gNppZIoH
vJ7svPhcZZhsuBVGiRcRS781AvDKnoea1/Sj2EEeVzKddllWSzL7pshC2CoI
vEqsbluAJ3K95rFFbMtloBiGKeYDHgo9ekc/J8k+DtTID8boGOzPB39x2AwV
KOVw6ddLV3f+gnmP1BZa/GEZgad05HVQD5bd2IvFtlL5aGem77dXlJEKxFvf
+J49HkOvjb+FFYhRkjLizR7IHRii5TsNAFFf6sFCCP3wcEwalzYnH0xN3VPC
TZYYmQH4LqM8nS6s94RmhIzpzzkYrA+SrhIBLtN4T5PTFmhx/hsg12VQAK4r
O18FeVmNQcheiYl2LRIVL7yvuzVkHy/NmVbJndXjfBe+Ep0ixAvO6D4iDUqd
ZLMteuy4gULvqv56svgKbppi7++CuHkUX7bKcVx0JWTwg9muQ5RvWh/lhsLp
DzZK5jabW8M2INGuU7LPC+zsz7l5+SQvNWkVXo1OkLtdteQE03TNykJ752qu
TcbwNs5r1vrL02OXZMENPPtM17naPLvfh+KUx47cK2t3Ynsj5ronpG9WYiNH
YWtOS6eJSN4paGC51gUKEnhIMqlq4l10+CbxttDuCbjS/tkJvYjShAWtPbkd
NWVxRQqXb8AbRUN7vglHzBG5uGObmb6vh3D8zBFYuOimMelK8pTMJVVvfRds
2ONmZNts6XcImY3owAJQLkDKwvNI7J7NWH+UXG2KMlXSedh7hyIz8+3CW2Z8
h+ZFmdwxTtIueH8ZYiS4Qeqjynsa/ognnDUqKVHRime45jwOz8vVhvi5Kjvs
jgFaCm5NrrXSkIrMGeqPjYqgOJV4Id8H4U/U4zmePZi9GzAOg0rEff8yd6Cr
4QWH/eCWtTe0u9HxbGHx2IfRV9d5b6GgHbc/yXUfpgu/HAbEcA/AZgLJ3sXa
v8K5os/UGh+XQnV3WSPoMYZV+AW58qhW8H0kGanl3gfVMjA4SvhwLNOvlQzY
wT4Ed3jy+V/3sUL4VSuXsg0kJ78HRuCafMSMYhC+w083MUwNhVC1H9NtNT32
M9YTrQhleYa/XenPw/StCRXuqHHW20r/5u8Z7raPfApc8r/WlwwPlIMHJsFS
Bgt9wOOo/TcaMFmVU+UM2O/mFE3yftunbudrINR2VyDKuigj04UZpAlZ2Usf
Hd7W20UF9NKXBVzQno9f+sg/3zT/XLN3A0a7sdcaW4XQXoFG3p5yxd4OraTT
dYHnShP5V+OV3n5W7YnZyG7wLSf8CP78BPqvMSkCsto55GULsbsYVti43TcT
vMZ/o140Wdw6FdbiZ5tDRNLBV+VnmDeN9PcW441FAZUriJPoEAjD1+mPFaVx
1XxnAtdDsK8LGN5Una5vURVdc2iRQ9dX8qBFEaSrk+geZ46r14ZWAp8TAgK6
geGds8KMmRlv045BgNNHcvAmVUgLLGbH982JGbvY4LiwaJgWWzrEbfnTADqS
lQIPcKmYYaM/Jmkt4accVQSG/6hALL7I3JDtQ1vPkCYcgLw+jo20dI6oLX1X
6zsNj4XnrwfH8PaVVn/tY+jWFV3HbbBdWMj/0nkrZ+1v6FLHpWAlE/pCFGsT
VsNRFV/O9oxT74RdEcJqR9LtFqtuTyVFCETzThgBhs01XswCzjDuYpZHVpIY
oLU+gAb9Ux4ODrbFc/1/4IHyY/oUTkjwOUtAD3TvARD3y5PDe01GJtwqXFD3
j5+Towp4HC00Et3dbWSnqS2ajPa4MRyNsCe6NtNXt49G+IWTt9FlHKHlKrvf
hz6ztNE2404HiLvIRR59gTelsDjXTrDs/vKCb0clpclhMuuvLeV4eYK9ytSP
xdM/1ojju/4b40uLXqrEF99tuQAXkm5C71PKKurFiE7UNc+LjEKiay/lgQPB
psgBkxEzpqC6kLYaA1EYVxkxQm5Aoz2GfviOa/xHfDz9h5YEj7ouT8jY81L1
r7hAC5PUe0B/122QaDDhayTQDARuVdVY2A+NnfNTtf2vyxx6CP+CYVXH65wk
UCcMJ9xOY1RsxsPElQUT+0OvM29jq3O3f2v2RVX08+O0nOfVLg0SpaDldN/O
xuSykbVPSbXJ4Xr0FoF+Mo++1MiHhgKuemWH4hmJACSeoPG8q1P7JJB+uuPi
qNEpyjYSJbYH0rlo4CT4RRhSaHAxz0A49WrYZdcikQa2u49mdJHsAFSGZDBH
0FbHn9YeXUW6XRBw3x1exF/zCm1c+Dn9fI4fHQOcTsOiNuQcgCMKwQmbQjvb
aN8wKls7WSNtott8owu4+30xxqIie5bFZ0N9nnlR3cqP6/SdeKb7lmpCWH/b
8bNmRMHoUnNROXcWGUfLe8K5fQNaCIgHTDC/Nux5XW5usqhFGSP6F31R8FrZ
ZlH4KX9LdEeBUzdeyfh2shfye8tVWCeSVCSgwF6nR1p/GXiA7282AGSIv7mA
kF9VY0pYfIu9PadETt6EJnyHSP22AI1lBAAdXkRuEcPwE7OxED3UFMF+F7r2
C9wlMk48QDD+X7hunSpTyv1/mTHjKarrlcm89nz/HJEuc0WTALoiUpBCFthP
ekOwVHGcrRcOaSNY89jHStVVZzAqcEW9IzpjUjbZ1pVjgfxEj4NErYYqwMEv
fTuyhTmYRmPkSLueNHYnCIjIhthVXzgkiQhkIP9SrI9sliiGm0ayFo0cQARs
8PVuLWExTQH7dVVY/JJH3J0GNuJgvdAON03OXq1KgAHlhHWz1yDk9ZVHHJ5V
YuyU44Qy7hoTGeRba9Kpva5V86vfaGi0y0b/UkmoLm3t/hvt4HvMUWGk0m9d
8G3zDWFXas67e4Z5husMkDzMX+EGk2oE3x32Y3ZZve/LNE+YBSf36yRHt/Qh
Lpnk9iOojD2eEhsFkGr8h/SpQuIAAO9qEf0rNX4ShsoD6NuLaHePnBffWuEs
CLX4F9oRiCvpR/T2R5VIlHv8TRLycbj8K42gmHDqwwntuy96I9/6Bc7FKeoQ
+ima11FVNPH9QUDjeGk3W3RrvrcGzefQ7nCe/eK8QO6EPbZgOCUZqQH6UGmn
xp+3aXtfddEdhKYn3zLANfIqCi2fcutnXDD2iGKnTlgRP44g7Z2rrh4zWPBg
mCWy+VeM076pXGHYXpThK5UaY3PPu+nl/3Ryw2D0JjP1A4tKt82PzC8GHr0l
FF1LTBach3OH5RatLIMVMnv7DpUh83VgbOrH1xpKV/loV9KRU5zzfIweVLSQ
0fdwy7Dt5a6A3+AMksm8nuZzqSNQLJsgh8n6VzOBm5lWIWRCXskR9OmighCO
LDxOifdCpAI92b7W0cHblHBW34ktOxp+emMobU/zqkcY5slKMHghKCWdtvDL
4dmerd8OsREURx72iGq30S4TrH2h3Qk2fllq4NyPyWBcZmaJJC3tHd8RJCkR
HoJEhnuU7DMugc54ut2uqeU7BNDAwq/uDJ2/DXU3Vbg7KachGOlv/t5NVLj5
0AGYljH5VY/xlNEzdjzqCaxy3YrLsjnZLT0kcY2vqX84NnGLpjKHaqr9HZ//
rEmtILFpvf4Yn/d1/I8nDcBEhgV/kh1+mesFIgwqbTG2yUYdQVAjRc3+uIfR
g387fnMIdgkgTsqjx+ic6G8irhnEmwhVHiCWor0+Y49nDBvYl5mSJVS63M0W
2P7TJObaeEh5K49EB7JRYsKe9ZloLN49DYq9Ecevp4lKzMrhq5Kho1A/Gfmz
RdVDghL0T5A0H+QTePCfG3R0KrbXkFe43e9fSfRqD8xSFYtRAsGCxTB4szdp
J5dY5oUStvOvVKrFnwK4q6DKA62mINZ/V8KIzzqLA99qLR1u//5UxNMb7ktG
ziujikkzhQa5HtpNklk0rs/m0ndBlYl8KqStnMvWmwA6Vnl10vF25NUv4yKm
LRQt/1twuskqa9QvI6Qh2/G7lr1ZCZ976c/PCC0J78Tgmfk7JH3u4639B8Jq
WJr2oBRt1wyGyuNA8NJiSin0QZ1FSuFOp82UocdA3dGLTYlI8mV0y0QHSu4l
pizuLHEiO6mTGuHGkgnAYCR89xWW0wEu6s5AiiRa8DRz41NF/13tni+NMged
PAhaI0zNUoNT6WQS+FZBG66jSgP5ZvJJidvaHnCLtaIzyPRHL7uXwP5zVQy4
+p1d1dVUELLRcEDVTKKjBOte/4P5cmSDMkbYaFX2rYTsCx37gAsaJj3+kY4W
lBq0bC48k75Z9csWgrnZkci++CmQdX554Jz5nqYJKdFnqy7s2jJ/S3d6+XH5
1gmJ6vqVOxaR4IcOHRWp8o1EcUCWdCHI9Wpb1jhQjI6YUkiGKnUgEw8nuPaq
Pm0ly80ooqeddxGZdmGiqg7HN2cVy7Akd4OnyRChKcGithQxfli1mvNb3C0p
d9YHaI0jShhU7OZ1amq7rtT9YzFByPQc0mBSGGmmgLuefXpd0+eAjJhBDiPX
hi2PAFt228r1NIjRKtWS8+XXEXGOZW9+Q4GakrU6AyFvjYqrFUBd4WKCBthk
ufVoJfPEclxNhoL4Wg1f/m2vUGhc4R7xENdNbdDboPII8kYBUebylE4lDNNc
X1GQ65oTwVkEX5LgcGGqi8Zzvp7tCWtWfTVNAZnKrmMLNc/RnoHHonfT5OVz
c1n/thz1jfu5DBhA9VrvUpgqwKN+GpMu4k0QWcWV11JDunWZf4Irbr+wX2cX
WRw/T7E1WO33u5jiwPPIERU7alWvbaV6lla3OfDU8hfxlmgrD0jiftwtmE8T
zduNC9wFmsjcfI+o7C9aIdJjEnQiedZYIpMJlA4PDoOK9VjPoFKTolO/zQ4x
MNWU82qot1ANqA+wKJo2RUzncfZGIce5YcrFAjkNkv6OAMKb58acM4AO3xWx
Eqd0U/WKBAS2HL5DAdK2RKt3/nZqUTP0gxgy8x9CX0vY9KlMtPW0AtH7QOTS
rMgdtBScyfgyFCFf4EBy64x8sjmu15c/LxpdpQ3BUXXeYTvzidolO8kWkD60
0/Ajmk3fFOMqMoCQDML0YSCAJI6ng/xZHITdca0YdFDertkNHQYhqpEek1yZ
rCDmKJv64GFQXTmfr7eu8nzNd2eeP/AlZyEaASLz3elmApxVCTiKJEDdeLqO
uyDe59HppuIquj9ED4ZBKh1CNC5NA8CCBMxNdPYzcUZozJFIrJ9cwGz+kz+z
TRHrGfdAeP0g61gKZpIlWRuJpS236KR5mGSDa0Z1/9bo36HibooMHIdNDNJ0
wpLCs/Ur1BkvzOiUbY/Uq+naKKX+bwLfheAveTxnLjYbtv1uD9+DKx0O9R39
X6Mpr1fBFi0W46MSENkFj+8bzpF2W97IvXowYReF3Hy51kaAq5TseagVwKdj
iTqxGfE5T8WtdY7HFlafCqbC5VBWWFmxfcUyzsmKfRT7LN+n4GZwRW3K0W8r
nsoXZNAjAHFdJ2a8eHlUEI1MYxNzu3N0El6MwNYa0iA/jkOgRPATR5FuTlJd
iIcUK9L326+KGrpmJ3000TdZhkQnoIUvAv58QPTwEmvREuQW342Tdj1n3IWt
+rnxq6T4btwGkBCkmjrb3r22fKuMXjMxof5fn6+myzn0/w1w8215WTWwplVu
c1PiC5czpvKoKGSLt3MtY9IqYB5RsM2ye9MH6NUWWY/p+oisgCP7M4ZillyX
kXbz868rIO1CHgx7eBE/l0UkoIENQug9Gesf8keWZThb8O7aVS5MsZi+JK3o
W3xeBlFBHDhWfSyYcdmo/OWHvr7qGZMuxiqkdsjXPJuQsA86W8ZOIsU5xQ6O
DGskHMa7y+dY5tGUaVBKcPX86U7S3sSkWuZJb/e6loV2qRyMZjLN1WQIjqGw
LBfCKxt3G7Si4OM1CHpE6FpCEiBqalD0vGp5LQkwhC5xCt7eu5ofOVW9mKq0
WSMWVJOSa5AAbnpbKWyiiR37YPi2q8itgNK9LMpEHy674uADzYiNbUqr9aiQ
22RAH3IUPSUDO0oSj5j/BM7+Q1jcD87gYE9zGH4FMUCF8awyIwaEHZJ0xWjI
7LskR1MoP1wyjd3zNojk4t2fWUUjO9SftQSkUniURra2AhM+kxzndRYolxLd
AxriQgPP5qnwhCwmzXIADCdQuc3EBI/K4TU5o7j/gV7P4dKszJ3I6TDYq2qU
p5ZxVAjCNYwIJk75ozwHZhzLQN2i4R9QPvwtRF9A9i1wOsbcDUAurCPeiBdl
aXuC0ooerrKH9aEpHVsFM+IkMEEnE5gRtVj52adnql9WZ65v94KC4lf6BnI4
LAwGx1eR4PvThDGlRuW3Lrq2coYsHb2Dr3W5a7CqWDAHkuUmEnSpLatTQJ2x
PHC3HO0AnMWwPF9pOnDXbaDMJKB5JyHw7KIve78gmufNxsnxrUdtsHedchcw
LpOxElGav/VhGQI8Af0IU9Z2VanoHvULYjYDjLCmc1utLB9WKEE27cSBaNeJ
WcQkXp5TnDX2ABye6XnpCqG9Tzz88FDz9Nz4OA7r0aJw0n6l8dihkXzNilPs
MqQn5x5/6l730Zv83KFdCitC3ds5j5XzUYV95HqN3P5IZziI8fDOWdxrK8k+
ZMlGrE6PgCC51HVERsTo595Oq35u7bJT3nwbz96pQZLpGXD8/rjOjyULFR+B
1tgjZr6IVwORRyE2lgJD8g5+ZMa1fBFOVjMaeS9uCMfKqrjfWOZ8srDnBd7F
drDSq/RBnhfcMp31JaANik/gKfzjXTsTRa5eKYiPt1NDexFtKkoZtav54ds+
mkXuH/lz8nyqJLsbKy5UpyUTwR2pTERrMiX7f3bBp1ioZkOngmPjsNEtwoGc
PAN8Xoh7lDqkeahJQDo1ghrKytJw4yPpTh0o5YUw9Guwhgb87hyeY6sm5t6k
p8pFasSdSUyjt6Yg2YeBngNMoCsLNKhZMy5r+NnIrO/8BNFHhHFyvFiGi0hz
UTILvhERmwngXmcn+FvNlocO9UVhklBeHBUWn5v5rM/JirXXh7t3ySO7PR5s
7JMRybZeOd22TbFSDhuZzQ77UzpQVk2TSD26LTNHCz7MRR37whdoJ1r9GBm2
dXUA6pa7Zb7AHVclJ/F3GMFdtp+3CTnPmDXmJUK8XGZthGYvRtsH7PeSO59m
gQkew8kIWW2hrsWR80gV/iQVH5DPE5zBCyJcCpCTF3pXc/4RozlyqjGIcBaT
xpPVxZbi+8NT3sz0TsB0us9FIzrEGvSYl5ZL1iCVJ4plzijNWvxxnp5/mv0A
/sEVwUNFH+a/kG1p/JPnsW5n3qdtfMCb2Ao+MbxBmHRwIwjN+XPjiH+Mo8EI
mL42Yp5/XHvb2vNCW4XCJZFNGt5XkW3tERk5ERe1qZ0zpL7SJZd8yuXrg3n2
Xay8V54JzQICw0ddexgevpXZMnhnMgQzBmejsfSpUpnKEaNXx/y/VuNOleMW
JkGXnPceldVNYWK6W0MLw52llKkumOnozjKiqbjTAW1XGxwM2A40nGlAFmij
QtSZ8r9GJ+Zwc0PVJ0JrD/C8hglvC85OVnenDrAqLkFR+v28v3r2dJyCjt2m
abko+9H1xOYAq8DX87pe41lj8x20u+NfgJ1P2BRYCKLh7ylZegkKXXFhvya9
3RrclsehwD6Zw2Yu2MertuloA+fV8rLgNguhVQxJPteMyEVCWK0TGWiG8BW9
yjFGf0Osa2PczlauVDeiWl6Ol1CeBeTmWyy/Rqgt+ro2CBWmxiN+oFXnm+vY
EiZni7HCotHCfKtW8OlmYxZ8xWVgsZo2q3uMELptnYs/MTWR03hpkJyIDQh7
q2JgLdv0MiciAOB8qB/GDQS2G1OWVHkbGCEAY2w1E3udz9EqeFkATUEl9+rj
e+IMfTMZ88k+DtPjy7MzSvTEabthzO4zMgRscDXXmx5JSD7doTMewdA6Nq+1
jiVjvwUFq1vNV3VF3aFimXuT5p0C79zrHvv4N+EbJprlaMYzhf5jbsnDv/cm
mLgGPXQPCYHXDhTx262mDaaNoZ0GCFTBskZLrQdfmo1o0PdyqFOMgl0Ex5kd
XUVwR3HZU8MXYdUl4LVt52VAywQToJe5yvohEjox7f/JGid04jNWTt2z+FfJ
ebUEz6yP+bFXYUPHk+ZNb03QOicw5tlVpvQnkl7GyVT9By40hy/WLXGAkIel
1DWK70RDGy06OyiVs4UgOauLbH38q0aHoAKzZq2A/J0WirMRiKlDNN5WNzF3
lm+cojvQUnddrFhgYFe3JsaoGr601K0hzljDlC+tUcXZp6qTbkjP4esNZUQS
w+Ho5uhvdS9j1B/7OcYQUJoplCwbl9/uF6wvHR6Ag1h6hjXCK/b2ZoOzayT4
rfXvYjmci25ec4iMbiAVGi8MA22xOZU8EySB4t/sWRKPd3mFxXX83OLz+Zet
Bpg5vacB2lAf7xmsmO8ZkTJz2xwKoq0ZI9cDysu/cInLD/lOqb6E4A2vQ8Bt
9HrFh7vW8ty+pP94h8KRRADa+zolAJUUAhi3lqbHssxaU1N5dPZo8UJ8hNr+
I3TlK0IUXfyC6ErE9IRlm3guy2a2t27jM233duEOaYaupXJg3GmhZN85qoLT
WUmQRZZlvVCHbvVpzuSWoicDePRa6+Kfj+6OmPGrkzLayXR0TpYEcgpUPKWo
3bAzBW0Ud0NnkPBKWfxMHF8DzMdwolB1hp5p9r8GCd5Udj+NzvyGrw6CrPG0
G+cHOF6VegTxenHjT4QVAMgK/JSrrBsFczbKxjgoWZciDZMNXiGdfE+ibH25
h85zYQ2sGocc0zSdZ1YL2bP0PIHMEdCIqWDbts8DWPS4yo23kKlMoOK5UKtI
O9ssKcgFwvEqwwEiMH8iLc5Dwtk2GBbWzCAuj3s3YBbc6dh02ZB9i57nm1RK
gHTX1ETeenTUlq4mBuQpxrB2ZkSq3B5QyilxYNrc064BxdiS+o8BurYwYi2q
jDvBkiW6rAMWuuDu8XDmRGzk5bv3DaumPFYc/9mccYnaESparH+Ovgsgl262
3gWkOvc5Xj7vrKhkaTBg++XtZzYeJMxU9BVB2nU5nMFtXUcNuWMaetykHhmh
VZut2qckhQ0gY3s5XZN4Xmj0cLUFfqE5lLmo67kGM40AbJPf7QdXjHOKC7v6
+8VNHaGEO25gj/g+J4kgjwf/ZFqpux56aqpqOE0iDYc4rfX7L6Q3Vs9mV+66
g7qfUTv9kDNE83J6NnEsSutIn8sC5WdVzCTUoqLtsU6a60nxoMW2XyXl2hw8
TceCFXPiUTKABNRykOfOaWYlK3smSbjeXMgjRdsKR/nVLZhj9ViwifZ9ni6k
8l7FtfhMb8aUGOXwmqm/lF1rfUII/2TMQxkyiw3kL48cDxGr1xcGFxbEkE8O
wPa/zVCpgQj/GawA+UEMjwKa0IURPTqRWBS1tYyloXeSQRRayN5xGtZfo8Kl
Sl6QtZt4a5Q9kbR2TnOuZ5meJ+YCGWK5nawrPqk3T/9o8h/EuHGvrJa7NMsW
jrHp50SavVt9u79N7NbCqoAacm0QQ7Y5pEVVjzPdT6vFHQgmUydNaKZmM6ro
nn1DZfP/Lf06gQEpjnZzuhDDwVWXd442/Su1ZMguHRNDLTEeyd5drq8x/aON
q9yne1C0l9lfO85yB7jMgzpgPujLeGUSmOyljbWobTjAxfHwqD6/fDK2HbJG
1E0TSiBbD6Ni0B4KUS6xiqLdssFAvdT3YndqulhZD8juqMdiiQmfSXACftam
1Ixq4zmuIiZb8xd2I5y/FyOurV32LK1HO8ICO8Tx+U+Gr29d9g6Q2TX0YUjc
15bjKTY3uv/3CBUVo7prwA4ZNnic92s/l3HMTq/j9om8MFeikY3AaAI+Cirs
XFuXMDu6QV7esDwg8ag7qtuf+6lcGNDUf1LccgEmMValpyt45PJEE406BExq
DB9C1CjJA0M4XSgWgoANTCS3cH1a1j8QQ/pqE8uCsVXH1l41Ly7rbTgWB1Hh
1UHyaqazYgEnBnk70nUOscP/vu/vhaPUrY3NHUHUkKgcfNUfAXMmbn4ZxUlo
db4PAcTKnqStjATp2nniWrcnXuOQABoHtsg89tf66HquuV8OHReY6cBuuWSW
S6rIeiTfkE5wRAFBgVYljAnT89YOEzaYDR6uW41ElqTpBS/8dhZEEoNntlyt
NuSUG40sbJCcOvuM/iRCfjnNYE0rX8GBaXqy2ioMxpdZboyAQwTpcN34SgzY
vPLvEg5hJfyFBtySaRkb3vnAM7BMHmazH4GtV2bdRLgGvoslONr1EaHs9rv7
wIqD9jeS9LU571BpZ/epusm+wLsoHlXmrgKdzA1LA6fQMOsWd+P1fRYRkENv
AmIuUCzAprYd1rMGWDsf4IWpgXKKDgpo6+IjA4NPnEWaWFUFqzGeir/zDTSg
7b47bYCd7SqT67Pn6JOZ1qomP+Z8YXb7quDlv8JxT6qUAfQ4otLTMwBAWK3R
Dq2qMr1X2yEV45doTUQTMPqfQe/MOTZ1e+B/l7Oavoh5pYNt6OD414o10vG8
L6U0RG4Jt8hFnR9XaT/9YMkOr8P7Kxyn4H/eAy933xxRXtHQQJiq3g1uHQG3
v+5jGSI9nlxc/iuzS2BSCDdg5R9q2bd2y9uoJGY2QjL4NnP7U0syYzr1D0xl
QoK3I1sg+hVRI4wKC68nfcwlFRVgZfXDrHKF842bKbDQjzGlN9UA4qJ85Pm7
12QWCzhJ7oGqKuF6OxoRy7wU+GlxjNZX8zDhRyfhtB63TVlhjNE1g5asI7FL
Vo6GFfZ/sJ7AiLGjsUth8VQmki+Voy+mdJRpI09mtEnjSoUShjcgdphlXGhY
R6RPdGOAIGFFS0JZfQ4+P85aRA7FCqQUzk/OoKMv8dssCOaiZbfEA4VXQgXU
t9n2It+kCoMTFFQUJ4q5YJpcSyCGNGIwdv6A4LHUcIRqYKlAoy+BOBeB22sg
YVjAf1Uj26B/Y1GprfX5JUXgMAN8HNkbNH5vmS11SE1Ni81t/6RgehPsoJrq
yn5KiA2gF678ag4PbaybOBN4dPRDWyjdF9l77wUCWwpRodeAZRVMXSXFq5pZ
OPnRQsvHPO5j9bImDyM6e6OdNruo/BuDngqC+EqPCfAKAGQWTxgBDeQ/bkf1
84K65d6COHv+1GHBrOBQ5yZUN2WlYSkUKW/N31rXKp9v/VyAnxOlAAAgZMwO
lXZKHOlP01DIxvsO2moXLmFuDLAFVtnnjRxNplGisE3lJDYRopHGgQ3Lc6Jt
8Ai+qCmI6wkSb8+U2jJmJIY+J0NOq/DvmE0kogJWlF6EBGO4rqz00VmOyIx+
3w5YLzprsqnoVCMdVIABkRvk1rMqKYSFqQKK++u8CXDuFaFLoY/eKvcVfX9d
L8nsQgSgP3SeWRLNpzcSfnBolX0MYYLC2FP5SeLpJh+82WSrNAuc4m6wr8Eu
e00pzsOuUFOVosI468oGIMzvbvpMHOdreLKuqBSGm1rSnJV9voF3sfYZu9PB
5gQwNXSZWj/5aa11+X/iyocPqy+GWWxdUVcK4CgBEKQulSlUD246ZUhJJVnA
yn4T7dJl8W+dJ3t+IJ0Z48RH/vmzFbpWDTQ5Ok+6VEta1ZosKAiV2BgqXQMd
2UdLnKDfvB/Gehp6hf9fzydBpGA8rlf2u1rSpsfQEjRX4f4a+CuxZmJf0Lcs
DgX5uv5k0QHHv3fkSkHdanAuW4tJSpHrld/UpjbZpaaXZdZnOpA8FaMmFuCI
Q1hAAFgnn0u94Ofleeuob/d+Oj56OBJ6EBFYpYojZy9hk3dSC6ojuKY8wLVz
WAVP+y/V8daktuMfjs9iOhJ2wCMdRloMS8rCn1poUESkEL3F85TycYUM7A3o
F3t5DXq/cQq8NqsQm4gomMHf6y2KtKJavZKWesegzVmKxz348RW89x40wh+b
JNSJ0lcM5gDqwP3kR7T+FngcBCq75V2m3uZtGwnBoKhzQhm7ojtdFJrusyTN
Illda+OmryTFOZL0jbgsnrbFd/QiZI2LhBb0bSyEB1cDg+dm+1xKGYCkHwSC
OMXfJmPdyjP+fTM/Tk7W6pwL621HNd7xnW6MbUKztVsZqUb8kBpqcmR3DbJe
ATxDP0azPfTKsPBcJEF/3LWckoNuKaXSVewQ1kHnEUUlgFAKRduW1kaeQc+R
MXHUwOFTYuB66Vh00ytr2pywePZfRHU167waCdCOoo6GysgkGK9tut60YO/r
YqoXtej7MuJrgq2v0s/4rc8wcXdORY6Ml1N4eEyrv30cAzgGddP5iXIxTLtz
CH0QETeaOGBrzPIKK3d1d2VO71NJxonK+03bt6F8nJKS4m84ZBcEI1pOsi+G
kQVqr811aOQsR22GCB268kxnXWo+A0hxz8aVHEYrMP8OfnRWALa+31aLh1R7
E8IGy5sz391bGKMAIypiJB85yuf9BrzTVB7hI29wSB+1xJkJHWZQRGRtVak5
YxJ03nHHasXG7Eto8LAekHhVqJ6Qj+CMM75vMD8Jl3JRFJh7k30T17wxtTLl
2cqx4roA8jQMfIByTjbOfLjNQIBFFdqVsFTVrEdxj4xdNDD3bUuC+5y4dfva
jH76AmYh7uPt2rvK3EmXIO1PeMAw5IZSSQKOAK/qddvNK6udftC08diGs5ZZ
Fu/kZndHsoY42ZNi00aGWv3FZAsF4Fm9K32b8+v8XVbM+k0isjd7QgFcXd7n
2Xmz2H/RfAQNjOQlSJFLgaWhn0qCr9nssNLRoS34hILw7hyAWuL8KuOIq5+v
vLHFosIrwg74rjXNDhmo4BEU3alCdV3i268E5+2qznFV12Y1enYf7gS9M9A4
/EOxTRAFivee/M2w3riLXkuOpPWoyOYuH1+7gZ1H8Eq95Dm7+/N6CLJPBp6A
LZF+NQfkykwwpJXZDGwSAKWouNkLvn/KybI2D8OKc+tfeDxZRENmQy0GMp7u
4+oAMBuXjHRSfQ031VKE2AlEk4DVICsbkRQCdlDyQy99wRbQBCB5el7Urcoa
Q8XkNhwgnJQ24By1I13pwugto8yrzh6ZKmLCnKKRkorEwowuPdlwcH63vfry
Mfd0sdYzAvD1I9vBNuBXA8qrb+c+O4RFfE303bJ/YNp+LIsaMMAWRF6Hpvu/
uBOIdrdT5tYP/gvnF6qTMDp0GGp8nU5Y0ASatHwNP9CHtiSLJEoNXKWVmoPo
QmyQXLBlG0XdaGcrYggocK/+VAEqwkeBj+NJqLEjBgW4wz3Qic3PLe+zUbsQ
MCLeL4zVy94Vwjt3oRa90CMTOttithvH+al5OwDl+2BnlpPL+0npmfC6vtzR
1SgZvEgdSlFNpNrNh+BK+Ap54h6cOkm1UYD0AwOOgFLq6pe2UifM32zNzehm
Y722OcNvNB2PD1+I17HSkBN4QpdDqs1GVUQw7HDXjEq20wW6MgqBbZL+2siY
MxgRg0sWgecM6n5LMYHT5l44pdFEHRxBorv8IqQYm1qcn7YEN5Kk83PgGqvG
3m1bQmkXP4eCYc6+kWF06YEwGVq35zP21xz+tCHDkaM8/PBhnpyYTV1omhqL
ImZhI8V+6tbgIumPfNY9BUjWr40vTj8GWPAVoFf1cnQfixBf6QM0QZPiRQMy
GqCsaey9KIhf79FA+i4bFrPcJ4/OT9lWeTutPD5M/g95Mt/9O7bDPnf3Kidb
+Npu1VLRbYsFTZN//0xqD9p5NiIIQtX/R7MeJOM+UQxDr81AVl28b/NBp6CZ
XHjl58HEH4l1Ub1s8u8bBiLwZ9Eu33XhotFGA+x8TmL9qaRLt9pwDo5ote9d
c3wqRjtQpDhsZkAfYnh200w/5lRvnthBdm4Wsqw4haJ8xyO+Xyiy3cl8zXHj
KEnwiraI01PVIs9D7mmFQenWEV++p8CjVVMjWSiOSqygVmXhf1hnR28yVYsT
TvjOTGdMEdjQkxTrJfPVPhBpyqKntO5yA5qrX2xSwNwU1T2/BS4gsbTB44GB
R04adpWWTXXu0AR7DBdHcky7i3i0hTZqLOBPsasqSpxZotBMxUbWrvHi2bz2
Gw2kFryrA3dYK1chwVQpjfBnMdiOkvbJcrrNUgX1bgElMvGQ0RgfWa4PDzMV
TDZ4PSY8/6YrxF8Jyxc+jv0mHabw/SmV09DuuB08sjmpTsQrP6OS1GJ6s6kt
3rqIjY6LcYbQ1/5p5mO+jBda0xMknl3yUHxh4ZN3kBm1AabF/HERa8slNQmP
PTgIsx/LygWtAgniDTtnX3H/SYOc5glh67gGlAlW6z01z5TbHwiwsAP0Bpat
oFVfsDbzHBGsQpQAkfVB7BCZvNvE92bHiAjI/hH0rEytk6BxlaTpq/Jmeohu
5sqR91aShjNZgqZa9WhYqBFOEcS6nNl2V5nYGN5UY+UFpIYFQ5tpVq9MZ9Dp
kZrAJWzFXmnLajDsLZPSihTeK+7d5g1VUZqKXCp5N2iY8/30jeyzGABVRXpx
KwQ2VQMFICHBPxDqedotZQ17Rv/lrxAKhTd0nhQg01AOuxbUHr03hxxjiKfF
OP0AZH+Un3pWxMaZ2L+JgmFZ/LBQ+2ZCxq/r4EVo8JKE6iP6Fsc35ztyO/W0
8lwFR9gdHs5c9VQJ7lQ2+Ms5TqtNJJmXODGYARmM6ZRoV7h/pxZLTPiboaB2
yPyrWjTQ10Iyzwq6K+EVz/ES58hZfm0+qmG5na60Sdc2PJX0T3Mho3+VIrrC
D/3PKUpINGFPRiTYIedPB6Gt4jIHmAGZtTGlS2YHUw0N/u5An941NuM71Qg8
CvUAckrVvGL+gSAX9lVqkrRgJZ1eu0UeBcDMuWlQLgx13HiSBWk1p1naVBj1
CGZfN+hTpe3/v46p42rrnrt8fpva3GL3WXyxBIzoxlInTTI+onQWQWqZUmBh
vX0Nl2tzjhzknSvCnFQq6olb3qio/MG3f5KpLuwMnLzplS2NAZRqpLs4CXab
Qa6o5LQAbOdhSyEY1ZtYykTKI/q1zGzP1zRY1Osv28VuaHbAUP2sSDoWJK/0
q+Jc98aSx8IxXYVf1qhUUNpkuzBAo6E6uzqpSMTtOtCCOSiL+HtxLhIEnx0u
U1d9wmjInMHYdg8PzF7q0+9ZEEDXbAsv/o+fWCkB7Yv6nUNKuPxHE5ZE2jhz
zXchrKVRqHImGtq6StJcIF3HwQWOgUueMVH2Wz7ZB3Iy6HbaXltYDbRluuRW
MkYbQcPEEk1OuY7solA1K+MJ0I5ABnYKiQRVFekUnnWxu6TFoD9NkcD05eEX
KRcUL1kepq/Hs4l2hYDV57PnyMm/lbEilxH9tLJQMYUQrOXaq7KrTBcOXgxu
4IB/MS1gDEZhQ0zxSN5ITw+RmDvsCOvyIE7bBO4BWu2lk6awxwtmgN326OHv
878y/HR/2tjqsH9d10+T0lQJ3KgAFtc+POJpWRTF2N1OESwl9BHHk3ixyiW8
h845cqxMePyK6YhicSZVbLcJi6CbJ/cAhA8h8uEruToKN5ixS9Ev2JZMyqgC
9zVG12JfUFMUBgjD5WanwMEHUf7LWk+JvA3tlskdqoZ+/umoLXzoMbp2tslH
si2eKg8JjH0Z8sQifNg6/0n+ckfw4Lv2fnQEbGa/A201eam7z5qcKhyJmpH8
0eYq/gf3SCC+iyRRMKksLkSOqYf8LglzptWMjol5ZSwjtHym+NHAx0Bs8Yma
icmaTv8enu/QMwggxcFsWv6wWM6sdgJaaCBrvEwdAEHxT4pIGHhS9YtbWhzE
CvVus38ah9v1zN+Fo1knXZQ867vHpvDM47TXKv3ox3GlTwn/U483bmNCDQky
Rj5ZVBdiA+091jUDEDzJlPG4t/SQEvyxpURO+9BFeIwnWUyl0uRUdWP8Jo89
iXjasb4sZIJxWdx+jeItbNxK8yLbXdJ/MzU0aj58NAroYS3/iXeQcadi7GK/
rKKvZ78W0fdzGplJSRo3dZsCHT2uj3dEYR3aAWc0aevbZSLGU9VeGyQWzwPa
Ba5N4o4+rCM5yLvNMtCqTNqskhVAo5zTzx3FOkg1fqSXARVBrB+jSkGm2mWs
rBdDJvQmSe9ybA5DTchh1B733A2FIDaWUUa6Q437tVaCMURXHmgpQJc/mclL
9Snyg9NvbYy+BZGp0eTMyXC1JtBv4StpBUh3mmbS2ymh+wwsO281L1lsFtr3
SlchRIsrERHaQpQYNl5Z0mxwrJzWg2uKoSSZ6JOyT6BW1yQ6hnn41TgDDwEF
IUJ9uoXIfywSVtPMEVFnnRmOnfjJG/ddiWugZK8CrDPu0kZ2yxJNkgQ6TN4A
CseqKwbAmFxwPJmKvnNtZg339rqnHZVu1J17YiV362V5LbVJXLVcAsCRlu+N
mnZuHl+L7E5F/oc9JvikVlmkc4PUxhkxnUOWhBuOSJPtUVGfHrWpA3fmrZvo
xgPrlhPEsRBf8Pt/FgMDhFoiEi3n4FetnykSVIZaFtj0uRvrHacPsMcgoYjo
VFmGn3SIa17g+3Qlo+uW0C6q7BcWI2JXfboPXCSMKfAkZerQ6IdhHg41Lj/x
f015cKjerUEhAg3Jh33bm6k4psXfz95aBf4RSPFQckHzRc8XBnrI8/QdzECq
ZS9qFpGJoicVhg+RU8b28XR38vn6WhVF+gPDUB7gXOwlNstQo030120CGUGd
vXnQ7mWhCwxkOuC/9RnriwSfQCopr7UmQBs+AOyT2nebW8Rjr1mpuvOzhdMK
8zmxONKVGfnYBIrR18trQeYL+MY6MgNIvN/jBUdbqdgYnvOMjUEaaZ7RJaLq
nT7RFtLJRnH700J0UENeUzWZ5A0pGOCpti9kqG31foM8idqdE0fbIxFcEYem
IYdvvIgO+1BZsUB1blV+MNili64A/njVL+gMTuGPFMVYFYn9maT5frYKdw+a
hEv5HRx4nKWCLaNYdSgGyPiwsxFbeaFh7braFneLuU0auX9eDN7DL8ErUp7p
7y6wToBd69sFIX+0ytoslC45i8N96R2TGPns2h5yeb40AjGpz5w/QBh9HJeG
EcCgtIOKC6gJJ6oD9R0eBdXxgFMwLhKWjpS7njL2EQq0hIVG8/8DMrXPbWVz
04id/IXuGtfQatlaQPj8BzPiYFd4Kf/1oi1wxjqZ7hZmLnvXJ0m1yXwNwleX
KMIrhd1SxzBG8O0sAs5zFI63AuARHw3umt3il8gOVZ1/eb82F8udh6+BA9XS
xnc55v8oQWt5+muH124ZYTQAchDER/dhkDWL3AUNmbsL4vy3Oay3TIE2QquG
0XZIO1qrCoNHDCQyK/XPywfhd01IkXWANYAz3ut37zkH3fMzuv44x4bftjFn
fjOFq2ZcuFMsNYHkgj0tn4iUNmPE5uKTqOQl6bDAmasSJXJ8M9HbpXX3MlKZ
97HGDNfjMTWOwxUsdPGMqhZMSvKNgx89GPJ9SkNb8uD12+g6Ky2AafvMgTT2
cxHRZDDilzNCbx84fUUqCXPUcHCm1VkZeeX0PXnD8IUV8LYnzlSFwLUCzBy0
078xjhfdNFP1sxuukXde4GMQMMNwhOA/t4RA72+l/yUoRbLeU/52qIRqNbdu
RyEuzDSJQzbfPt7E/NHsZRl4z4je9oYkDHdxsR7v4WXEoKPOpSjUAMouTZ4M
yr/zhwpxZMJHesLwI/po/p4jrj5QPD4tTMGx4xNS+6aI9Rcl2HToCJswSmhs
9pfus1frMhSG/3WrsksVu9W/CbkEsn4Qdb95Cm+MWFFi0kONE2q64BfjrhHB
XBZlcCwewRFFmiyBepz0Qw37GyAP81JLsd4ODcxKpeImQpb3jVh/wgz199zZ
dKc0kJscM+e4JGFm7Rf5PTXCqd3RZX3lNOjVXCWoSmGoBSF/ndCmclYXKmkG
0eJIX+hZMTtmbdbK85u6lq8RcD2oq/1tIHhYtSjlPGFhWTK5zuY+NWxXZ0I/
G4QR2VhoNJbWphKPCNHbTCREZ8nAQvrX1PMqadLjBG3I55QuscXHSmREHDqZ
njGsYbRZfbzf4O8TLF5o9qCAMosqty03ZcSsQLi/wwHX+AsNPNJ2ykLq/Yxa
zCZS1bG46CJajpBKXeOQZ0D6T+iWe5CSO5GmX3RMhwJMXPEeYj3gVQc85JbN
plQfUlmCIIiVAnpRWNHXQx7AO1NXtsuq1e7j9BHdf40Vcua8mQk1AT2V99Ci
/EE9Ua+R6aoBZ/kXxKCYv9irEN0UeUHzekPGbXa19PEu+GuMGvsHfiksURuc
py4K0/hF12xRJ7Jkz5oo5A+gamL1vujTkWws+ikE64HmF/4HyNNmzteCeyww
1W9MOCYzS2bFnGCDXiO4oobMJsvI/Y7Ov7t63xehZWHNxl8MzGJh3gLAqk3U
vj7xPslZBEWDWm2p9ZQZKYRQF7HmwSe2o/FzmuNA6X6G/rNwK6p0eFvyZpn6
o7Xp2UWQMudwpcAaep7jVGD9rnkYsRG5ou7fytNAGLf+6gdqp0LtRGbnKaDd
dURmvU6MKxtn4Wf8R+bZG4I5sIUgRIONKTpm3jSW0TYRAiP+5pt+UG3ZmYw6
YJ2RtiJ3cguV37w6a/6RUeVf6A1LnyObpu2Bc6HSIfFBj2+jSNK/SMWu0qvC
qIELNaAGpe7Zd5PToxbLzmRbX/Ssn9ktZ1yg87adyVpZWPZoOPrltvdnNDWH
Q2qchSXx4DuMrU4HrC4k1qVdvNfpZw9W5D2VjfAA+BsxhuYeXTqToxT3QwH7
0qIHO1dof41SX8DiHpAM+q212N3TSus3NqKvaa3wlfQe7nYMeo2oEwUnZAxQ
Ukf4/wCtFKkXMj+qScwbXewxwMD1AWXF3xLM7LCoWa6LfmXTA6GZpMRAypNO
ixcrpuiPueHqfO0tW636/eeOb2LIvlQ8ld2yOg3PPbTCavjGXYVt7zL3d5hL
uydxJyp2MmUFJU09fUxOdXXczXGf2NXKpnydqedeAklHO9eW7wize+C3sRec
TmFSR52xgZRufmUP0vy7uoOuS86Befpetg4/N9TQSZh/jUn1TVn9XzRYZucC
lYOsBMEbtnoLca2hgy4DuN0FjJLa6CglIRjr3Kiccp9edUh7PClQqs31kvlQ
uw4G6iWZQkstA7k5SE5pY5f1F/VUqlHNvmwngQ8UqUcCkLc+Q2FUu4I4aUbi
XEpb3ruqLSYVFXXeJlHc9jBixqyfiGmBEe4C3ypcbhJftjZMjJIIhQUeEc33
71VwceyK9qWv+8CEO3Ry6yfrrobrbkIf430XghXhIwdK8R0uNvsafdQ9Xe0E
ocPQawGkIC7reRJ6EB7IKCwi083JL/z4/GAvOXDb5woZnTxJVhLJ3Xti/bf9
AJNXHnDdmyi4pPUkH5WCaUHgZzMtxz85wCiGoPLMbh3RmRENTS++yfgq/YVL
hsg0907d8pwLCc46LmIkFVyVqZXWQzJlVBvgucVKdi8l3GIT/y+fNH8zCixZ
Xy+Df7Ux/UbetKFTD2nR96V9ZonM2+UETI7gHCmwXxdYdWO+cS64CDjTDIoS
lYJmRpcqRMyNHY1d3drB9iD+k4tCI9eyqw1BoGfiGh0z7T0euJIK1thbIwzH
3CapNB4qjbOn/VtHUYbrFCfSwgXcrK26gl2M7QgXe/2X6zER5Id21iubkCTm
2GKVEGzHb/AYux02ZOWS/gTyddn1nLQgxF98CkkwZ6g3vfIK7A4qYdQTGOhq
cDF8aBIyWoaUIwot/t8Y08K4J0Z8QzbYetA9KwJ06XVsRlm3K8od4M6pnTok
wHI2OJ6eC7Fs6jy4Hg6BNsZnGJSxxz5LWWhGvIFjzluEshQDuh51r/v3vyg8
Nhy3nnxFUO9P0/g3oqKW3lTRiyC6DnhIyeL0FNFWd14MXjq5ooeZZlUyeIVu
g/TbuBD1GoL25W2BsGxKDF9nTAQ98jiMdrUF9EfgqXhJ+44N8+9wXdiL25l6
77yAud3iT0MUBnj6syfS6+2OGhz27Ev/mas5pjqIdNuPuWBuKSxT6fIY+fyK
5+gd6HIFmaojUVSavaXm/KWZoI45faR77WoXsQeuCVkUXzhMMSvXBTFtBCyp
yn1I22riSwWt4WKSRkoUOlpfwwL5KSXul2elt9AYl5JdhCOx82ty/1mI7zvM
nAppPfmZGcBqvhS/XpsmfMqsiLSotpPJSS+2xJQHK4wA/vWWmRsbI3HZJAmv
GcBy6uufdYGThxscnoWrlVti7AYQMDrlMoOwnBo6xQtPZZXDr3erAACPOkua
BQVPdkfQviveMjSsoeq2VoErpUwX/sOYOq43Cdm9YSwWMF9+IoDEqWcg3iAu
2UB+RfsLHd1907B6e6AlkDVYVrJyYT3pmpEbqjlaqqmppDAsCfK0Zu1gjlf+
7TD1bdVyS9gLhCO7dzfATNX6j1yLZa65HvJJ8AOrTv+PRZ8mVxWsyY+PBFj8
39m0zexYDtAUD7wNC1c0gFAwChJc6GB+j6s2vfbXEZjB6LAwaq5kO8RTVEzP
/iwVG/45YkiyF0c3P9sLeUx0P3Z2EDNX6qX8u0yUrQvdOMRQ1OKoyRx+yG0W
jXJINj8va60euR4RRi2ewNnsxAsxdowZKZBJIeC4VLGL0x9rto65keWJ9umj
4eSrY1s2ag9txBWir+Gs/nU9mXvHAwnl3voMlhDK3+udv0zSOlm4o1gd2gPf
IthNLtbKtrobEXMx2AW+1qGPQuCUrvvnt3bavltRIxdQ+N7c7gd+7lhORHmi
HRAoz3aLDTWWT1qVADRw6pZxEnGW+zwD8gDYYsi2VERpZzaLaxkrfccC9+3M
B/JlDiByJJRcjotfw8f8CExokqq9ZCjb0Y5vhDfWSCu7lSuBOfhB64hhEsjf
+ZKpg7teHTutYv0nTRo7jApFAh64X/DQw+RYdw8khHK9eFb0GIgNuuSoeOQn
f9FTEvnM1IVQIqIDyqDtwSVHQRdf9/+J0J4OxOiMSzG7vXDPr5u1APa/7BwV
rPiE+wNaDNfeytBiDlYrq7sAoV0XUHoRINBo9tEFkuaLeAnKqdTlrJjZ0+x7
2SlLhgH3PZCkJKmbZt+lKNVLc3eZ8uvj1r/KRvgQHYfoJo/w6uSlbdwOuYBl
SD5pEFs94SfpPzYnParhA8eApSYCI1Kof3P0RjV+EhewYcdELHYcKqEOCemS
5cFAppyCneLYmkWCVN3WL4uVm0OlcT9PYhb8OOaBAukcgEtRv6Ris9H6cDjp
i1tCF+AnDxw5MZYIJdvquU7pPhUWCJlsXHeXY4WZEP/SCUnIKIt0Kk0POgd3
J/nJe8ZHxYBQMTIKFOTSPCk4lwWVbufmMTjz59qNSBTI/q/R1rf24jOo9oPe
hqmK9gVnBsRmiXz+pG1bNYhhC+Qpp8ijI9g+G0+anb9adLNcGeDxdTRYh3Ot
8iw9Nsq9Cu4fIdjgUM4npawq0nqR8C2NB/tgT/+JHE+QeBvddZx2vHilkciI
sr/yaOpeZNehQa85RatDkZdlJz2vmnFNUOddnRq4MR7QbpVHYRi/DVbjqIvP
n87+5bkMMQoHojYCG+pGdcLWdo7WrMeaPcZwKq6N4uHqn2NzT13Br3BL5CCo
Zti4VOScOGxh2borxdN2Djxc2o+kmL+/HBRDdP3BESYg/APFrL/1BzOCrDVC
16sATHOPhzKDJVD4P1FQ3RqDwSbo44Fj4PqokSqi+mjYfQIDVHQEgxTw+6H6
B/57tKsgtYRrBsUm6eI+kxPYdCKHBhvWxWYzBwsotQCjyO35QfZpGURPkeBe
Cj+ADH33+gEw40V1P0XwwXIzLJCMX+7kz7H0rgY7CGVj7mN3wRZh/6ewyMrz
jqchMyxTFigf4ZaeTbeaw1bboKPcWQ/OsVwQGSSasYV5fVKARXWrWvrBUBeq
11uZl9e9MCrgZg13O4wH759KRf3SDPg8w28z81vjkdZaz8cky8tdetzbBiHG
rwKy3Osy/CsQi5RsL6YfGrunHnZR68bgxeReP009UjCu+WGIgkPheXW69UXD
xV70cGGxd5a6vhJSlkqeJQQ56vSaEwWCpg6IdpNK97ReMSEX1JQnuRBlpN7r
qlmE2GPU8Z6oRLQHkk8zLOzApv+au/MzN1LqVM7tQ9STOJcXq+w9P5fC3S8v
O6WjBRaUJFWlWEeccnl/sSU+uS4z9jK8JD3GPn+Dr+lTx9BUhXje2fVqgYst
VX8tFH3XAPpMoesvP8IMALooqbYAcC2DoVvnHP2V088u5wioh2dSpE4VryAc
W9wQNGdTNVu2MATJ7tMtD5J4waMl1cdY7vp5WayrbD90XoyhWddrHpT4dsd5
db6OKXEZfbXml2umXEDIs6UAbZbrkQOHonXXnJB2c29ICH/pJulp2Z5jrhtu
FFOfkZFnzxZXIypoqcArKkGoAZLPbC3xN7tbZRkdswAM2OS8KTmhrCmDegNP
jsroYDjJBMpCcw+adSN3rcbexA7KuEQv6d0nH9ItxpXBqNULucAOmRxVnv+p
m5xt3sLbBbhD0eW1gr3yszGg/Mm9U4BjdbIds4MYKjt49EnraOLsZOBB3NFB
c8bnaCa+eM3KBR9LnzGWcE9Ai9+E4fu1D5ixgKAtFBPCwzJ8V1YEIzf9unb1
7pnpUO43NPYKTFMboDFwJGGR7wnSxCy0TkClEmsof28igHg8fQwCxJtpVW0Z
3/EWvHQmQJkEmlO6nFwPArAXwXG9ZnLLg5nlnMDGa3jHa3pyhORMqyzkvXG9
xGMPEVk7QUYjoMzFU9dBZzutky4g3PB5LBxHcaXTExlWE4DSxxfCT1HDbEOv
34ztSviJvW7unTfnZikpyDP35V/iy5WpjiINnZKtgexkEp+ZkAkuu9DKnuJ2
M0G2Cb68qwiR4GQgsnf/vN3yBfJEwE5F1Qky/8bukAGl3tmzRSs6nXvPSlxF
MfivTJFKERoFqZ6vOMsUVs5C8IYaXLoFVtez1OR5uQrwnnQKrx0Q5zbtYovv
W1elW3LX4+DcW6UK+aARGZ2L7BKwRKJQE1f/1fMEtMfsF4OX1eCIAy9nd9H+
lu/1o2xDqdiIUMFcYZS+WTYUFct5qGy0rTQR85MUZoLZ0jaW04SJ+oxQ+TC7
j82+cKMvAKb9IOqkAmP0ghYHHtk6JphZ9rdYqyyaC+zc1ZRENMTI7LOI1x6T
H2brwtfIKGbBigQRHp60wGqza9nlmORRbO1LH1WO+1QjpqLKoQFqZtMgAjqa
1K+tSyTLSvimVJmp7l2xFjSRiUqX2+xGG3ICdgE+ND2c1EguysBvunDaUAtB
4M2bNa6zDqUxdkrMmG/0xql38wpdNl4VK1DZ968uB7akEoALJx60TGxfe/qE
3a3hUKEGU3/JdE1l8aL4d+qTP1bCKOk5tb5mM/AmeHrFCBdnnfiJfs/dsJXF
x0aTfik/k/++VJsYMW+ua2HLm9wPTVnoUgfsSUSSmkjxFRPIU3uJ+hiRMiQd
W0d3P1P+ApJq79Szm2UUQ6eIZZE21DQYFYFjeSozThjIyoHoTnhYwZD6G262
ks5QZINoaaxxWuT5Kbuw7LWJECT06iQMjCo4MNKkJDJSsDOeVrJvQR0vYED+
IVP+a9OUGuk5t/7emR0kzZlBiqWlfMVfaok9pu6qYcsAGZHe29PMoIK2mwiL
EDmnTWQpXBEXVJfQUv7C17ua2+BqknYOYzPa28b1zrLzWUVN9m+gIHkiAFcM
1Zf7mRC4HZGlVN/wfBx3/OSPU5FJn5YNgdZhXBW+zIsOU3lZT/DXZn6bjwSn
88jdiosgCymSoE/fgl4jZzWhubbqYZWtWXG/doo6Wit/tvbaVK/q2i8v6GpK
OFmpHJ5ytbmQTBWRAPjbTar2FxIBw9dL/6IDvzccXpNN3S5BY6wOZDMSnknu
j6qBbtmJPYb9lP/g/eroIS5zc6p875VWYxgyt3W/IuxF1Vk8UFPsFpwqrf0r
LmF9Aw0NFZ9RqrC4Qxjz4f9L1yQc///3WMD1DPwUgOE2EC6bEmiJ7seuVs3G
EyOG6fYnMCWPdXSAtV/+b8E5GbCqIVw4THLMXr+A5gQs6X1PqVnFcKJudTYv
hSUo74SS8Zq3sonRRCItmzsdw6pHF1dYFG1FmFT1m3+9yf3Nq1C2lwyX6bUh
u3BHn0ECTUNFSJ6pmx7vMJLrTr7cNjkvjfsYw2Eo39Jz8TuK6xNxF06oE7Lg
QMiQVr/eOWE9mbX69bz0mF99QQimWM/nT2fURDoKRXMkpoNAsUa+eSHkrmaF
RUv1S9EkCuIb5GJbmFSVfekW//gToabCkgsKH2oHGHHnAvxTMLzpyyqLanRQ
uNbY7knGpw+KumoJeplnLO1CPWAvXAvRqd+GseoxArcf96wN4ZdfPq++SZAx
TCMc5v9WUNoHNt4Xs112zOwE2aQG39GzCos4MrAffgmKgUM+81o1IOMZ5GDA
3KgklpLs/WrHlMHi6xDyIBQxQVOPDzS7H9fMUAOmxQCMdubL/fshd/O4QsZT
1zO7QuJxkA6cZeMK0rXtS8mWbayZ2thyv5IBCuwm5Zv4hWzO+ru0Tr948GUH
936cicWqu+NkMG4ziaG7VAIMD11wG8BP21JSFEeNjR1vk/yGWJSPu6k/1++w
fCJ7TeTp5GR4aJxUqAcTmW0ryHGVIV7wTsS1LedbIimSo5INphR0y/L4W1rn
p3GKHNaKhWKB3umgB0YZxSbrRi57koCkdXNTAYrd82rD5v6FuiWitZ6gGpTi
HnwVZXIbwck6XrqQmRa9gvqAVnmptvyHTGCRO/38HtKM17gCKXu6S01oa/Zh
2+ObtGXfS+yJIMjsc39kfus2mTlrLwmUpJOIiPviXWjfDuT0BPreDbAP2dvr
cFxHEgfAMvWMStBCA6sAQijVxxa3yBx06f7j5jjbY2OcOgJLGP57LHZ47iCo
O5AG+OPxbdwXqlA/rxbmIh4noe0kgpWOq0vhBJADVJQzV6rJnKxJH+ikhMHX
G2ZFg+0Mvos/7u5cruEtteSq0tF8jZFvFneHoO1dA+3FLOZPd7r7SWY11Bcd
fzsPeFDbdkDemTu8y+gPK5vn9OalIONH+ZMw+gy2J2Bw5zMNs7/dsIUG3tmw
iilhtDSNg1AaaAkh/42+/mAewZfP6eoFaoQ2P2wRD8A1kfOJ/+VsKxH08lZi
vnZVhvbJQk4kHYWujh5ZOVTx9ceRuXXe086Wbi+2Asgmfi4WNKYmwADNpJNE
b7JolzEDhySU1rM6+l1MyyhULjd0n8DhoKFgTDNYNfJw0Pb5LbvSre+UtNej
NyKWq5WpQpXsOG/NIUb3IqZmPPYEse0Txb5op8DWpTwpcnd9JwDhdVIR9RNo
+rhjfH/apY80ffuySzyXRCEI6BZlfztsEeR/HEf5gsC3wl/xaa8YKm9ce33d
tlfdqZeQ0pHVWOvGTktKXv+Ip44KB3jkOF96qFFKrNJa2ZpNM0b5j0CY/4FV
m0taPpz5AA0ThX2ePMVrIoQLFcTc2t9UfNqpmhHDPcKTz2S/G2UK53LCL2l/
IJlOF8pzKNMlby0+L8VFGBhIlLdzuobnEZ1rZnmiLIxh+KZeaMCA2ic4memt
n7u1KD+a9qyRpW+hGjQg2eVuthrZ+kfGJoAiSZ0OUxBAR4rFTbjTfNM2ACcX
yXSnIV/uSKIAXnHSCK1WjYdnQjXS5/iEsUkVJ4Y3kkt6smKTPNtIUUFgnrzO
ryOBfjSsahVROO6voCK4n2u8Sdl3DrlnQ592nj8KUR44PYHkv0UFiYJmakBH
ffb3NrkpZoNdZIYTY8dMySSI/6dIi4J8eb8uvqZ52BhlLQCi2guNB072Ek1v
1M6ygVCwc2B6k1Wbw1YcV7P91VyeLcbssIO1trOuCGja/9rUW5CQniN5FK1i
LMu+rbDpikLxJB4pTfmVHxrs+xm/z1ZuV+ddvKun9borDOr3wge272N5+mcu
phr/NqVHaTxLbI9N6HdKNiqEaj7+biYFaWs6IQih/ytQb95kDXmZNz/iiAfp
0IGEq4xOG2RWIj/hbr/F3FePYdcq/JafkaHteZ6JvxJ0fED7VPye4Y7YK5zT
WAg7q46k/W3kigwmiskLCNlrfpqCcLB3tWfqwcszF7ldYcIkuOzdCl6MKWnS
nuCnvaaF0jaaC2f4RVplJKHUPia2rBaQhcZGF/j4WZ2Z+0Cyfj6zqaEvwNdZ
sWFrTYD+lUWcw/HRfZV33B/YX+UdnRxrOiOAZMHJTnHXph2Q86x4fSwzwAf6
46HfSz9ePC3JVZ191FzJpMrWV6D1hgLpR0y588MG/8jXjcOTGU5AArpoEAv+
2LDtvgRFOqfwW/Xj77OhTE0Z9btqthYrIXIO+N7S1losp/xT3vwX5kqCpG/c
GhS/eEWPciC1y3jsBPnXoRhHGWgNGDZdUai1KZKeGna7MvRM/D8t1NQLQZTi
/UbMhvZl5Qco1S6XDi7V5MrJ8HI2AvyauOSQucN8hMyWnZvmVJoQ0bTLazSy
WEG7R+2D4lw+hXilhTe84Qh0JLGMUz+wjx5ke3qIg2LfWp3N2s1IP4wLRuNa
kBe8ogl6/QdHDe6M2pqBdnim9+89vxm+43B/kG3OdGFWJC6B98MBKySt3xrR
FB8Z6ULR54wKj+D6mbonUM4KBre/HaujpzL6iVxXnQY1ymrtEDsFMa9MpaIM
UOkz4jyPWdSPqavDP0kBhyi3smSRVU65JsaiPiERRI1G59rizmsXaxCNpM+w
dZBcYjPwEW8ItWBNdOkmRtAXySWdmcJs18x+fZQnI3Bqz7pZMWZ8GzLLadYG
5CUyLzTkVbNaPOHUq4dqAZ7/jg0W75In7QyjUNikxl3GS3ylIcaPd90HSL7R
+mXSRewgtzu/+aogN5ROikyU/moLQWOfrV2awq6USoKdubeN0ICOnGCTNJgc
ZxgZDf+P7ovKj2IaVDf8oZAeoe//zmQ/wuMftOWGVoOZWRNXJ0HLoUJec4EI
1GUhchKusmbNNs1/xqmgKG8tDMTu+VwL5qB/PgOGXOOSXW+pzfN/kivT5nI5
ERLz1aLvWUXsnfR+2iUTAw/ChIyNUQpreRy/VDnRqqChKufgZ8Ztx0YeDN8h
8UobG3zPy4QgwiVl/sTT6S1PLTsUxJ7FD+MaGcTjsaN8MkBoYyI65t/7ZTgu
nMdN1i8QGZWj2QtfsG9KCk0DExS/htQ5edIR3nsbMyOza1KmPgq0JmkRVTjz
Y+RjdhdUFtIIftuP/lrPqcO5Nj2/IuWnjRXByCPtUDrvKVamkltIr8SQzQfO
CVYx5v/PxbuYg0d+1Xj7PkIxbQQlHYxJlXDiywH33GMlsl89kx1bM101V9pE
6DZ+KQSyAjfJI34tqqlCHXIk58cD/h8tblX1j+Eab3oiZW6wkK0bxAWJMfpb
MRiW3cH+uuFLavhosBW1quQoK2vR/H19yNXrq+7GAypQ5WRP6Zh+5OXkrOJR
tdK/r+FAc4yUsXS5nhtLiwYoLurvwPBh2s/RT/uRsGSw8bPj7mn6hBdjhNy0
jeoVTVnu4HUWqD41WLDx9NfZjlCZmVT2YVogITSsGFC+FvZQeXLjpkt1eywp
pFS+9tWZ2TYERg7ft9/jlxJ9QnVOGnLWS9MErGk+NTX78XaxVwUwa7e9l1lx
E8KIOWKIyj+/th2XFteDbuEnGkkgGeKzp7RfFPIryE7bW9zYYwJwIxp/N5Ia
fx5lrfbWyIP4Ycrp4DRNFjOlQYpuh2N8tN3VDgx7eAre3RGBLLpt6s0znRMB
e7Edo8dk8VN6D/axjCqa1EqwipUuqbJITUUggzcI3VC8hv3WRD4DwlAlmvPY
SA1CiHmdD4zTGzfcrxccQirLWhB31MFtCvr9zdEOIVFwTXpu0Uycyv6ROlwr
EhMk3aJqhG9w583T9Z8L+1xvONotYVRyk3fkRUoEPa5TE1w8FggPy7kFEXVQ
REUVhnfdvfZXN92upxtWzMoLTN4XqAh/JNuReu8dsadPpD1e3or2RDdOnmAj
l7CI2i7xdkt9YgGnnATvZGYcNiXT5tvqvSty3w9Y92uty0etxLMn1K2nXZwV
2SaclK2uGkVmhm9K9iaOy9vELVFhVG/KbFKOE/pwlaq312EMn959iffl9bwm
Jyh5mdeRZ2MSmHsU9f+2pdk5Sc+238dI+HdxarArxtcPgYyff587BCYl40qw
ZqCyzCxHxq3nUOYWUG/u/CenrZjFXDrwSYdkFatpLQUnW4Tyn+hfwsxd7qfk
vOCMjGgjdMvfirrSuCGRJ6eQo+j3sOWXunnHUCjqIEZUQHyxzy4rdPVqROd5
Ub8sjGnk0WOoalIfBiMYq53JT0FWhe4JWkk0Emg2hZ8PwiYD/ji39Y8aLT+i
OCcSTbNYB9tN6bhpIf2atYRg1UDEcM8wAHS27HYtbsK9xQVG49R1t7UQEizy
vmBfdjaErzMSdRhuPrSLcr0011I9bI1I1IGzoHF0KSi70I0qHGNURe4MP5a0
VmyFsJrxKxCJILKjXpI99mczBSLTuxPRSQbLnqFGWP9ukdvkVGAhx4XXm+Kg
4xEih+dfYm/Z0CQsHpgknFvOqyrNOdyd2cHMj/IaT7/bQG3Lf35ZkaEnT04i
MbaKuL/JKZjxicd8bDxa2KEiVVwVL5U+Xwun9xjEBlz+eQmKE3VekOMCSg7p
z99lYvufqEepgYRNWxABs3w/bFiHpHimhMbIioOb2Y27vT/5jBVbiG1bF3+B
NRxZ21J50a70dpdR/w93Ms2LYIo33yYC6Sg4Zptf78Wku3MQcgaRvFiojhWX
gUPAj+MOlPZGLYmSrxnr4NqP26i38hW8Y6aNIlgoDfg4jZRQWgY+44emzvVu
OUAxgMR9rBwu+E4IkOxIN7Z4TJMGQWyYiq6psZMhiAeeh1MDvRHUp8AAdJ9X
AOyP1sb4zQ0aKQl9Hwzu5i/VDnF+6j0kM4qid8GX7dZ3w0KghpHbSa5DXVJX
ebv0iTH0ucxEBCpL2FmvJTsm2PqDTpQx1BCN8zMvnDkfnOD9KbtJz5fM+e3i
AMI4PF7TVLSFu8CuyuVS2YdNMz22Y7JJgOGuhXxuIGM5PTtbPjHw1rB5SrvZ
xCOXsTivRzxoYJ2kp+V64K5GaJHUb6kAsRHcSH3mYHLXbUuA40JK1ZC3yIQZ
mFLHmhIhWKo5tYiNwe/2EyWqHD3cz+YAwcJYe+TOg67dUHmaVJakyUzyZGD1
nNoAo89rgVDV+N18JcFDz9NmyFMP3IPQsa1v51zqCp7pli1+cghMLIq83SYG
jofsMvudqqkpPbdMfsE4HLCsMhsPZA33LXjV6VDSGYfUOvatqSEBFbgiGDLs
6raVYSIYutjqs6wDWMEYRqPbAxlBvLQsACoftzW54I674YwcdJnKoZnmUZpD
SxEwiRkFVROiaatYTtj9QxORcQq13OfYy0ugOWnA5/RRW6r+ghZTLyUbv9E9
Z5CE7QHOrojYWEmhJEFDbhjWyM3RQLZR3WYEyt30xp2KAZI5G3Ec5e/r1VI6
YzmTkjMi69iF97jD4NFbWrGndPLTwqVzI0gEXMZ9ExpKHNQ62u8SZbBwoiw3
8krZ8blTCcwSmjcFkg65Rj7x4KJom7EwwsxPfdjaE2m6duyq2EmP81cJhR2F
7vuWZcefHritJiYX2I9BG0ZQvof2QrXeHVdyYl0RzpbmNPJKBo20ylR0k0pc
2r8n7LjGAwGMbWLe6BfiqgxwqBpqL2EOM2Lh/IGyq8L4m7vCE+GlfJgTf5cU
fJ6B8/PDjYofwV9wXdC+GnOej9sLpHbRWt6HibzgaOcK1mqFKROPyNEZkpW2
8DIiBgvs8tDjYOUpuZEyilh476422JPppow4uY6Fij4BbYApfQLwyPmqqTkD
nHV/V2YIdU+/qAhowIH4iFSuG70eSzYhOgkRz+s4NWQmKLWbn/E+pbSmLuFQ
080m1WAFMT4RIpgJaFJPV7+bHI2JPlsDFJjhLcTa6PqnUhdIsP5wl2W0tpp6
MphrPrsq8i5o/9ddNYua/BBuy+3Qq5zayhCAYV5A7kPHLEZFkVV562AEIYhP
oL2+i8xnaRHR5Hq/FWgpvZ0JFaEwQo/5m9FMWdE49DqGkVvIRTN+Q9iSD4KD
LlYStuEdnY3aZvcGvyotu86+opyUoXBhTAUI3IPFxuIh/3qPwsWfZ3zFxklU
27z++pGnU+sbIZvu8Qdc2H2kpGUo2OKLkmn02blgQNkGu2D0zN44FVlIDIjP
xMDHIS2v/315ezoWcm7qAEwSNX3VjzgqDmeGbDYeMJLaPeiV6ou3zJp0WeDK
HFTrjnhS5EPPgsKg0SP8JgPNBOy2J3gtA3hXmuLUrHvq3d5cxS0Tf6lzPMj+
6iNbe3ZdlBnAkVT9iCd9cSShdZrGYnrLchVgAxfLT43MX4irgJEXOEvYED7q
fqcslGBe5YWM1LYVoTD5mq6arQ2WnEf0CiUwhlRpSQvfeAuNifqSy3dRBxh1
XG4/OB5AHrEw9c/jdfCVetdCOTBu8yVR2GfsJTf/iTEMR4JqmdsAEbkhbRRB
HRxDlzwZcTNG0JkIv1jJD8dbm+419/x4ISBMdJij4KkkdYi2u8tVUxG/AmA6
aRDeON6HW3Rpe38Rq9Py5sJ3xD43DRG2oDL+Vq3z0DcuRFKLgCHIUS8wL/CQ
QWmBBwmpddxQ8N8YmYVNeAvURsUeiqZ2xVGOTkGmcpKtyR8kMhS5nTZ8Fx7a
K5Tjyqb/4wlJMakkMM0W2z55qq+zM3HeVeXzlO03leY9/5w6LN6zuj5IQqZ1
8HtWxp0EhTcsCYdnNGYCcsMjC71i8tV3Mlr3fcB4TyDBExzd5NaXsogF1eiM
mPrzkM3QHpuPyeFXudAa7Um3pxpmjlJJecyuYsXhsajHuHl4k/YzDfv1FBGz
Nrl+mFyI8+spVok02MKRO4g8B8pB5yvH1faZCGA4vrSnnViPqtVFO1MZ/XS1
rO/tJazPxGx8pRf0BIvrnKsBQYClXLLlA14NUEK86tNeJDLhdIGHxlw0z9kL
Pw/mZaHiz4UvjQis7jjhjlCs+4Lzug6+YkV/TzBfupRQD0uXFsvtWqgNehzP
Wmc7gFPQGyJmWMvx5rKoEvI0ZS+vnozKyavUUmUfwBbB4VT00b3TH3XjuoQw
DQM3y4GCRBxhD/hdqikGXJ3er/gcaId0whSAFbIZbdJYg3m05C8DOgn2EoWH
p673/JGrN5lchLmzPbKuI4RTqcwrL2/6wTSW6R0j+dY1VhoMj/BN/ozpyc+5
Q52wQeJ2yyEAIpsRbU6j5sV8T6ChQUj2DYpy6kKS8RmNI3AzbvpW1Ui/9DCw
46+Th+xdQzCXYPzPqQvgmu8zwFgIIrPniR4OUtcaJmhlkyLkqwQBp7pG0twL
WAb6pzthK4UGv1DHMVGURoTZP/NWUsi5HXzHtxDP/ssoxP1eVzawhuG0nrs8
TttX2OSYaUu1qXwPn1z2NFGujqwEpTMSvx5Ho2mkibRsyI3NeMbdYCNpshlG
ghstMTdosluPTt950j3KiUU5t8FrKdUwwKgemXeuteaRX9MVFo2xE4BqhCzM
mERt9igESAaX7aOFJrxrMS9hO+hpOcYW1K+W19NEy9qk4/1L7P31cjzaqQlU
hOOLGvtxHVbOh+VcFSHyQ1zRQ2+V8PnRG8gHPa2olNuW2cTiQIGCSGK4w9Ix
Yp1bIHBfJAv3QBouVVf20SDg+3lHrIjHlo7yhis1k+5A4IWDDkV1TJ8af6FB
feM4NleVhQCo/muRdk2pdmjH8En+LxNP2q7Opm2XxCYZjQmNMCLfravkdugg
vGt3Gycx0qk9x0kWGLX/9BZkRe03fePjwLCRiDLlReUrrpPF52doc6QxjgtV
torw+0eeUtEW4N951yr+qEg9HbO6PEategkQi7ovFZdGxUWdboyKVvGMcnCL
AeYkWCLrL7VA1gaUOrsxCaOOFZ1gzWs7octv9/xLkzOcwBppmvtbcKm5S66v
85w9ufEeyQBZu4pll3F/m/y44Rnh86960Sv06tWqfDQuqY5ce5r15ONYDyYh
Egs1lh30lNuvJVHd7YpB1UMstBVc2Qlu8yFy/kHMUx7TPE3CHKPckGuH39NL
Oe0DjwWD+EkqISjP4v+c7xX6l8+mxYsky/MVSLLiQS3BDpqxJdKG4Dv4+x1V
Mqd18SUprdnKKI7QTKiqM7yFUxI5IyM0HUja6vcMT8NXJnf9jHvPGE7E8Ly3
XMhKQIv058axt6WMwHPivnaj0dvDq66beQGaRE8WpVp8UTz+E+rr7kEHK3ch
jA0n4TdhmPJW/rNzUaEPc94EyPlYhZb5JMKqfa07Ia2K5ZcN6NR/1thKFh1z
LIHESJbkEZo/A1OcWRHKfcv8mTXJ81DiV3xNsNXKipZ1NyRskYANOe+7FFfZ
C23neIns2DCq1k6VB0fUCUqjJlU8mx8SJzLz/jHXXSUD/9aJwBnSlPRd+30g
2WnVkEMJwhGOw90d9um+TRaD5M9Nz54PMi1jWrKwohkMJ/4bEa613t+MHs7F
flFZ1XmTc3Nw5yACDr2tzk2SnUWSv6tOsxp3LJibwXt0kOKoL8SepR3IZaJC
A9k3IeNm5lHFEINmpWkvkWZGPxvImrSvKG8hZcpJ1FFVnUTm1sOGhO4DnzFf
uaBQ9jqCLQCnJupQHwH4H8tXff5hwyqyhTY6S+rq5mL4/wykRJLkCSc467QY
kJWgnmT7T0Sdy41Top+ZQHQm375ahb3TjYQR0/Fbd2wozy7cxD8Ozbr676qY
hbLNB6Isq9YWj6D7tAZmaRQCXnbu7QX4DwlaQgjRsATnE1FDIt4BeYTAfeP7
1dgW6JwBldGhbfrdKNwu+pz6Rs8PuRpFg10ydZryEQpyEhsCq1heHLvJ+DLQ
d6ka8J/oApzGHUqQ/i7wBx+yPPaD8bPn7oZdDEI0lBL2ui7dVc2H81auvfaB
U0pXT+66eAbbEP5PlCjO2E7XtU1nwkjSouyosz9WDNTF4GG7qiIjctlLxCt/
RiGwlINERT1E/CnXaQw1Q1Hmd5naKuCb+D4xU7a29IJ+GgSnLS5TxNevwoa8
9XqrIpJVu4w4C9Q/x6iEdzOugqPC/X3sMT/8LEKQQ7YdMMZ1XeRk1sN3/5DA
94mn8+LvX7TUNV/ndlosbhx1Yi5szPNTTcGKjEmPxKOgP4BL6ILLX4GWSTd+
itvbY5nU+XzOAeU5PIUNL3vLrIU9DeITbluuFFN5PoVYwNhDnk7WU1l0anVv
zUPitY05b2GhoJZ00DqXueXX/vK8ehQEy72p6yc8SdjYgJc3kEeqT/Bdou7Z
JwAINoyrBbJ9DwhySWwLJnG291viNd/YDv0W/1eTPqnNvJtYYRoMW9u35OJA
qvylHCmEWCV3IH6FInO6MVFUYO2CrxWZPKZBzbu4bwYvJxB/yu/drusE4Pz3
/Pk+RCVWi76r1RItN5xr5lT6s6gPQa9XRBvX4ucCRUvRU/x9fTL2PnfrYBo+
vIRf58Ffna/gb2yErBR216dRODPkQlyvQVXhRuWLVlzOM3NCHpEO/ktTJW+d
altFG2xwPfBH8/enmWCtJknOnzCUGh7BCfGBUA8ZDzyJPx0tylvmLgLZvfF9
JP5F6K3gw0ssJStlVzvWgpUqfgs7rNWsFpW6E48AU226lMntnQYD+cCwtNbL
v+Uli/EYxnQI1Czr1kDlCz4e1CzyMNXvGJska+iOD3BWV7sTrlpkf1MqOfFf
PptAA36A4BZWKSAfL7dLbt0rfN9mdIMqH1vGt7DCpvUVb5Pu/OS+6r36B7bk
0fOPbyp5GGYmqiPqyAwyVec6YxF55jjxR/3afAObZImbCufX9JlGAI68JNd/
2jrRaXZsWyHGwP/htcg6BKkfuHL9wHdQP8/KRwBx2mLEYWUbZdOJY+e8sb+k
2Ew17wrsIN9ILQ2idIU/4xgrDEw7PVIAll7+A+5Wd+vSSx2H3EgalVr1naOh
50zTPXH4rj7906KR5FW+DQ+uwt4zYsKI1O6J+Bh/FgCHAjlKk7HBZybrpqsd
bil16cytj4U721IM7pOQidPloAm1ieXwRvQDH6vo0denLTVx/oMTMf9PDlCI
mTdh38lyfdS/XEQQ/giyksNfy1j26LKaYbI8Mo30jgfIw4gALXaDpxJ5QPa6
wCsIuw0qkIFwYeLCO67kRT122oFya47/pibfjBYpUTK3xzpR5a9+wRrLSm8N
j1mcbRmLpud4W4trIykPkrzK+crZqf7Yt+km0HyjFBnEnFRbDWWjUtM+WmcR
mw4fzSSEkaDRzdEZrZmG3ub64pl9xhl7HHsFp7UwTdcFD/KYav6ncxcEBw2p
FSkyZSKFvKcV4yPkml61GA6aPOubTVc5HbLn52JGQWykCw7pBwOhIG6e8/7p
f2OJp/dHon1z6xpWSa3r1ypsvOLpYRAP8EbQ6NjsMVSHBstTaA6jTfyf2kl6
qwfYsjV+FERIYmrox76DJRLDlyJ5BJf1MmNK7SzVZRD9+l5T3/eDIUVToQGq
JTykQ2MbaKRMlBMUJSbQ52ZcDhbC3zXiUi+yZTINQq2K2924BsCE6UDNSXtO
ttaGYHfR0o8hWI1Me3oKMgkRTHP5J/2+M4cWieuuehYZPekyUnO4KMXMe5Ge
V9md1zQ0hu8+Iw5QuI/R6GUj0lpmhwTmu3Aylm/WGsDLSM8r9q+EfgOjEBkU
SqJPyrHx1khrIkw8l6RAEliWyWy991ZOcG6xHp6m0YxrcycbTqCoS9Da9R28
is/n04DjZxRUKXmTbttRM097XESRx7AWImCl4UVzc2zpNGJ7UyFSzStN7RfM
uVYen4Ge4ZA38NOd5zMv0LreokUMMZ5y/lmZl6LnIoxFJJNL/iEPl2Br91rY
JCreibk8uPxum7/q51epYAVJEtpdFwfVMqdRHotnqx7kN1BImIfMRW0tYGpQ
FZ/Wwhj6AvoP33e/v3KAA+lQQQEb5f0p1LoK307sjphmrguawIsRH5MXnHCA
GlZ5+Bh/EHjbM2cbUcG/ZaP0wr9WLRuX3hTii3niUpr/5cUxE+LIAULpusZ6
jN5NJX5HTfFHJDixjbNsCz0fz0COPrAfnvoSDlCDbiV9xINnJPh2B6AZdp2Q
JI/wzFHvDDzgY2UqFZIsZ/j6wVEovceUCNSBJ3KcYj23Q6uHjB7dgxT5t+aO
fArJb9Y7uiUr8/IUnhm2riskzIx1N2cLRbIlIv6/fX6mOFDZKJICNIm2pwXa
R0gb/mJuBdIpfs+hN5Yj599OAYcWOrLNBYbxgTK6tTf7d+olx1WLOxeQWvOM
s69SwANtt6780q82kWjpZwWwcd5lHSeVR6sBOPAYtkZfpRXKmu4+vH7thHj7
EK5LwCwswtnUbzdKqk/5QCIbY4SuZcsqTTuBb8U/74oj7cDsTazPGn3ShjjK
M919uyoJCVgCGTwT0hGjmmvBd7uUAYbq/bhXvO/Aq/BOCjsuKtdWwluazev0
FPR6Ofy7F5kwqDEz23Cz7viJ0uLkK5YAzyT2b/X/nBXXa5Tpf/RdyeBz7mmX
Zi96JE++YvFzw7z2jvAfV0jTF0rWOucTT4o4+T/e/Gs2aGSWvMpVf2p5PUkk
LamBo4ZMnEfRP11Zqdn6eqolKCq8lkWjwtmJBScvTgYTUF8WSJGYeKR0Pofu
dp8MqvTVUV7+foNoOMnyBmTZ5oFtaxv0iBd1J6HWPjiclnh99sDyKHx5VNdd
4dMVDgupyISSmd+lTrC2R+v7k7B7bSmeFjpzn5+R6+Q/j3FLj/M5YGV9WpgP
FEI4/XQwcwU08Mk0C20q/94QIQ33LJ69/ofCRgXi1Ru8+Mo2fQib7ae2PFGh
dJ/Lym16/3lQ3mIlKXh6nodWQm+xuL/LkPLmn/mec9JS6slj5Tgra0HBD9F1
2joiCfNpaLaMjw9ibUJFeHofCK0yIeA5ElPgUfHo3Ste6nRWKrdsyluacna7
fttnNvI3fsf3YJvyT706b40KCnzmgHzHTJrK6JIKJCKJCZpGaAcpvlwD8BjC
993TKGU2Ok4adp6WRjOzMKylkKgi3zuhbtRacMuoGDkCecGSeW8MJXMUmijS
VC/se79eVbp58mGXnv45RbDzTr6GLTZYNnCknIdouwHhK/yU+zsTj3LclxCJ
JS2yXOVLnaTd5Z6BEEgcTFZXTwQJYxyT8KB1jP6nuIfB4wllNKS7KQMhnxOz
BKjYuj1wu8Z1UJZbf82nhz96q6uoOhcTuKnIfFUNi9nGGypyOBKkAAxSQKfb
pePhFcNpjasvKzXLzYzm4jZmuAiRQRGhqkkgD3o/72ubgeiqXCkDSg7clR3N
FyalzfApRYrSXzTQ/jC9lc9Z3zx/jKUibJVBJ0YLjtBeoBOQTbdZfqkrpGSQ
QCE5KMUTlVuF2dVhIhWazv0C1NSD+sFMljfby2/08U/SgxqfsgcJqYnQabW9
5jxPjB9sqUrckyJl3iQLKi8P43eFt9hHyI3ItZEbwAIl3/TBVkQH0ElSZ1UD
dYmPmdi49E1bzsq0Z7OsJ+Uy2PqaI6ARQ3GN4X4HDKPadleq2YrbkyMdqfZ2
c8BmtFi8yG6/6d5i00EX0JG6kZJlTH/JM4SfrnZZ+ejH2EPQwmEfj/+FsRct
iSYZHjo4xnGrqAEh1zganzCg5s4o0/nt3sK8Y0kQkV/JKEzG6KEoGD7E8/Jc
uyVosujAhIczfdcCc9ojwDtq12x7nnfqs/TCJimhLu20pnwWYlUhoh40Vei4
c2QQ/0qoj2XhdgjpHxoyUWXauzrE9W7RXNHtOVVE4zHGP120D6WPQgSvRWSc
RWVv53AAJwYCw6QXN2j8U7EiyBFodVJ+J/YimXO99rOtDDSPR7YBru3uin0t
ceNZkudt6zBW4GazDlboPLhh0Mm47KwGq0fVCKBlQMy2EmD4h+AInXNf5z4w
NYThrmNvFUA9EeybsD8z051XM8uMLLlAth8WegOZtTctMoeW9IgvsPE4mEMw
QvNNv6uz7Uq/2oxZSICso1fO7j0eTuwOQhCg1bwl71mPeieNBGgrIJV0Dd2M
3ZxMpKPmpO1mrNkELPfEnSvBz+wxUX6Z7El0mHGMahbaDlLVGAHKvAjmg2TK
bWJmKGlLxibUvQaqNTnurOu2dHL/zinwLuDFjHBTpe4wRlEVIGAmGJj9Skz/
hCMo9mzj56lNAizB4m/F2TRAVSdPsBS6xjEn6McqCePzimjXCLchlVGLcyjX
96+8n/gjcDwOrmFWtaNm+47rrUlZF3V7TygLvxwbA2MBdUvOaI9Mgw+X++J0
PP5TWNKQwdqre+CjOHeIU7Qpn6iwRL7GYBpyrokQPjQdr8X/KSAzkWFkseBa
qDhWOWcCoii0fOR4moxw30ZL4PJ+xMUt17ptGXGpXZidVU60oi+LkijT6iDw
GP13Cb5Qq0dTnXA/okM3zXtaHzTfhv8PZ7ADaCdEMg4zwpHBDjY+TAYiCiVp
2GRXTPeyd55bCVZia3cbx+rmjFcKPsjNAEZHlD8VYwdBXMMgD9OOAJdIC6k+
AA50dIaP+LMif3/joyf+THaYG7+UWhhvXUS9/LePNFl35h1zc3+82gasTdyE
VHQycvwQ5iHrZ/4PPMRGX4XkhKsRA3clmt0udvDSTvcNYqicV6MG3mgJUH6p
gYAxf0pb1vajMFGig3g2q8n7HiBTD22r52G8JPd3NnoXJz79nsm1eFRfhAkR
YtUoA6ssRrBYTp9MqoZP1DLKwTj/grIRN4w4x9ZEeO41WZW1qkzDX6GDGgvn
3gRUW1yAFt2zAjxtGhQpKP56IczhK1SkkL9i08XHdPt12a646AvGrh4qcZ/0
olzVNzO0Uigwnm4BUilwPTLJrnUo7OeQncHqFl9WIDYbjE3a7hxu1rMA2RGI
NFT1RXXpzaRcIOms/OqWoZWOTN8FneA7/rYCYN6bOYzwiAg13VThzyU5QVCv
qhYK+ksl9dUaZ/ca6I4lzKI2zDOf8J5tbpJriYmfCgmQA+XxKhFhvb7G0NhX
MXrLP+VwDu+dVAvD+llPdoe1Sl6u0VYqvHpoYggJO5t+nP01FPo2iElJJmSm
Aeh0cMi3X2djUe14P0dXnPPV52CmoUEm7b0xnUWVJ93S3y5l2f2mvjy9cHXr
MIt0VMVpVSa/XFBHC6nD0V1sRCV4bw4mnK+/ta56AoXlVM8Xw80M194TVgAU
w7yIPSW/qciCnjuLno0GTe97ul7Sn2IiTjzi4nw/L+1xXTJd3RSkn+fBbnZI
pcYkT1/ObowW+26xmJesxmAhYlR/0W+7o/+ZSHTQFHP22XHtGHJLgh4D0u6Q
L1OKnD5/E272fRYcLTlyoo5eGxwdtWow3dlZKNZ+PSik2wFnzPozMrsq4wl6
S+aLwtN4HbPIpzMSigF+L7HLQgBotH/oK4zgtfw9hY3U6v8vRx/rMiHoxP1V
bLkByUgqu2k+EGYMmrixUADgGbsEvolHQ2havHYWnPF3ohm+qEuQyunLVven
B+QIzqNrkPuV5CcTuZzAQQ1bqeCBHcctpbUMMdChBegkrDqmWNtB3rjW0Uth
xZQarSWHQvxSlrQlPg9lE5ZyV4NL4+0twA4rU0iTVOtCMgBzMzBR2/cZXIXa
y50ff6W3mEyx5jWW60YuPxQ0psXR8svy1E+O8u7g9jmcOhYvsihllOZjTPPQ
983dQMXs6hR/tocSTmMw9WpHTnWxLvcOAMiy1G7pFQS9rzmwEwoAOA6mKi+D
ioo0vmm4W+hqEXy7tnbj325n4JkgUfp6RVARELbn1csXu16ZgbOdx4TlY4Zw
2TjXioYgUIPxUdGrjAm6nzMPz3xxpZbmwqqVm5eQ8+EM4emDQ4YgTWrm8Mx2
0QdTTYIMAtb8IrIgYJ25f2ElJKqxKjXQdcOu3Rg1iEnqhAus8fxrU6vmF26+
MPsSw5Q1/3WxI1VO1uG5B1uGXsjsamdY0iqz5YOu8kNh+GNqEb/5oZdxzmJI
bREoKRWrk1yQ4SK6KqsN0Zrf7gFcgJgNCNOSQUI5I9xWSr670VEOBzOMNm2n
eNNJNmpNzaAjkQlDEr8OJZ+SNQFuN5NH56rt/FNyu23igRxtgBoA+E6nFyR0
AQ0lipbYsu8R0UpMv8g8ykD/JAmX9P1qQXnzewQ14FsCh8ZgcrAGwmUG64RN
G7DNJvitJdJhEN0vsL4A4G2JnY+YhANlXDBwL57q7z6Mr+fWqCTtEyhLWhV5
6HWA8qqIdded4mwEfKulLjeJFrGeUCa0TOo0hfcZkc096oZhTfTVh2pDj4ko
qXdRSWCxXwmKqii3za9em/GguGZ1EFmitiA8jOquodeH+bMdoWYc9ovYXNqM
EszSrhO2ZbPurSlSbnPeSD9hrbffbRCKq+K2eCvHz4cG89kKpPHMixTUFyF/
78F/ZWP7pctwG3+Ul7TnftHuHhB2E8tmcb5l9cbwOD6ScTwN+lqdvHqLhLKp
3TGIe15kS4MzstZd2rmbO/09q8iFFmg3fxfca1tf8HkwxlLfNSgEaTT9R/Rh
GLF2Huts0hMtWoIVSygFeZOkCoKUyxhF3zMS300HVrIE9ifpyiwPmON7CFZ/
matzyG2H7GSf3vqVXSI50DccTepVBA6n7/2wbFmWtbf106w21Ukjca237lRt
sd0DuTnru6YONdXfaZZRgywQWts58ngJJ18Mfv1CdqvNtRGHWE7M877HNMuA
ud702xGkBzLfuiPGXLYVGaf1KDAJ8SxfWpsq6KpCzayc7WlIqW12eWNklhh/
rJvWFVJ/qK68UT+C75utiyDEic1rdTT4fYUzAngYhaAjDtmW3VBohtuX6N0Z
jl6rIqeyBsqpWi4xpY4a+pR8xqE04HOO185ORnpN8hlDPd+AJVwVFECalN9h
eW8uoZ+0fSehwcg1fm9q71N6HUZAzdHAhD2Mkd8k7q/Dcg4Pmt6SW122cKZZ
go1SyH7WsX1IM7l/shKNCtfJdo53TixnhUFj7xg1TFCUkhtHyg7wbMmj/wdd
JZ36zRUYmzBaAKTu0VEUhYKYYRvuOlSNSgX4EClFcnhHJRb7Lxgb3kl/qzgP
S/FOegZBmAbrIdP9VWkzPzswcGyWdDcbtvl7vczPSum6JlngwPJlop/hgsUn
NMSrw+5bcQl0ycwZt6VuZDmFJztPvJsIaTm8jSnin46LGpIXSEQPBGiDtUo/
Ape6i1qa/tZDcL09xXYW4CezJEgMMPaUdNnEnQAQTKZk2goQCBuzgCtIDeIw
/7MUFgcsC0yoJxWCiC7zH5+J1/IW3+SBye3v1EhG4Y9mMHJN09WAplmNj0he
79szRgqQq3K+g4XvYnztnseWQrIacVM40ObLnbEHBQonhKIp51MLeDzMcuM2
jXYyHjJRMM/okE2KFngAfNK4inSlt1Zwdw/fluvbuhP3REQsREFoZuygSWmT
6s0mN9zInIXBS2XTlagdlBBwGUTyctmTxX8Xf0Oons4BGoewGbgHJtUf9G0F
a+0A6qmxgqOF90Z/BDBgUzX/67QhKJT0NZ5l7KKz0JA1n9slDNbpcsLL5qee
vKliroVnSGXs+5CGabFANPCVuS31Q0Jn9MW88nBOOyyRT4GJ34xC6HlKcd89
5pHfdbEhJzON9SkqaCWWMb7WEOegpg+ap9PSram3a+E2E7lT/uuTThBWD9g3
z9/vAz5gulCqti5CMUnBuDiHw8Ng0Vh0Rel3XnrB2r8MCsi8pY3EdEC6IHrz
U5T1m5ULGL+hBGsfyyuzYKeVZbBE76UbncIpPiTITJgkHUgtE/5vHr55fQtk
Kqdex4ks1frHCPzgUJhkA+b/tmGKIzLuTB924TyfSqdvVEm+AOo/55IBrFPN
wvRcN8fdo9lcToEz7PG82hPt9n8xLKzwXWvbIoSHkkGyS8PZ30Qz6UPNeLNv
aZQNDMZXH4boDM+1xWE386pCHZN59iDNTpteUFZnv+AGIYbZdIXFIc2qCWk3
L4x+6fxOAI7/IbzCw4++9yiHRv2CFTmPTMKT2ey6O27Keg5WU5CsGEELFXUA
ZbP4Uz5qNskDGVOnP599fT35NsQuOprAyzxuz7bsNj3fs35VLBVc/dQh6P/d
+olVp6SJx/QPqL5czBKc1UUuN8Ut94JeSv++3ukV3OrJZihP2rGdYaedz/VJ
H81iCVkidLekDUHo2KJLorgGhNlh0HqB5Q/eo0s0sRMTFC+TLzUJ4GttMXgh
QZNV+Mf4cKdvrFjsoci8OXZ98xuD7CHoQ/oTQ2EwonYQde9Q8o94rWZ0Q+d3
ydITLJL2R945syIPMhihbHq2p2RtMOknEA17bqnGHKezOG1cl+Fr3aTmwIzf
g8RYIhtk6PYCiddK88/Vy3R3O9H0lFTz+PFohjPS1Xm9moQYi19kOpUsmWZF
w2E3UAUBKUFyucufaD5+3IuDmCus6rxCt3TiI8K85pJMmwNMX1qi4r21dnSP
xtvORRAgxPQYBpiI1FcsZrWhAv6b4GGLjO8oMArf2PoNl/xyxh7gNg+zZnJd
TUV12VFZAGR5mHqa+osQnEad4GrvKS9BQB8rBuIRuNsy+lQxLKCsvsLVhAs6
jAreM0n37M2aYeftRfeyrbkpOy88UEN6GOSyt0oBpIpRnFveZUIZNAxrhzim
fPmYAP+I85w1z7YYR8T+NhWg+pHNkwF5iy0wYvDwQrpqzfOHyZPZ4ZoTf/xN
wFNs35m7Ivpih5lmbPNpjK7SzsAkYcVutPYVDlYW2DlgviR4RehaZ6MOC/Ba
1i+sxvHxXwfBbvvAH8KhJnZHLQbF2gh3MEo11I2GuW/+BV6KaLmJaJCJkzVU
jpOw/uBTUF2J8YLyEfNh0YKbNok0sTeEn7NS59Ds1JNPYxTLABqXdVviw5qM
fbrxcOL3+G3sTvSKgJAB7RGRib3MQMq82tdWfvKQXFLUBHHUZMFER1l3V/Eo
cdPFrmhargzh3DDrJ/ukRJoKUFX5e7qKCJJRKlOcGyPCAJFZN0zz+mGrK/Uh
v+DAd42V4Llr3GDLVDrN+z0AJB8t8J2sUOhhLL6ze0UpLCZfeQUrWhdZ5fjy
vc9YG6zPQ0NZJwa7iTJPPt3rbdIit53OrS+/+o4PhBs7DDCxJPIa6EMPTfzA
CF8O+BZUPa9QcKosepCZC2e3PUAAw5812Veu1fQrREn3FbZc5Zu5HC+Yqk/s
kLCb7AI/qwIxNfcI6pJJLQ4/jnBOW7sd1q3d0Y9LilzRrWGcjHH4ia7Fwuqv
cjDdKCI5WD/Zc5+prp56Drg3VXzAgpEkNOT/aAKCoXFOjydbd5G6D8cdJ7aJ
B1ZXV4ADVXS2GHGgZaII0+6fLkSztzJEtdE2HN9jMdhC3UHgxedS1zLbc4W5
/vsCbuKJ96lkegGIZurF/57Qp1+o7D7xvt2PZWf1heo/joPB1ROuZQYnc9yc
x+TQ1wFR5TGydgLaARJ26q9MMkdDyZmUpXuXIp9MPxxtvJPY160D2lngHWOw
v5pf4skF1hXBwG7t/0jVN4fvdYjC47yP5K73whYPkLnMlRQ1SEl0ZvhNSC0J
fVGY4NLeKks5c+xBUJ6wfsmUOkM82rV6oaUANMe2+dRYPgX+H16PujMnyurK
L6J2yV4uirtZItowiQyAlzvpurxAooSxZDXAh4T6ZH9dJ7J9ZW/HQKhLfP43
li1EUr4WGJUCkAZJuYuzzn+h8gvUYhiRlWvYI2eGSQeMcjElK6rMm39m1C6a
ITngxh4Bfwmed2PuIhbAqg4vnpF1Sajy0EC0Plhv3nDhRqczMFKXvQBwj++s
9CN8IuLLHl7kx1VykEzyLI7uj/nyO2P9NHICYBfWxjyU9XIUeNV39ePsORWn
UGS9b3YWXB0iT9yyGl7JXRW9PS8phTppQdkiMIztesiHrgQWFB6uyP5KXabv
XImOzMqfYk9FI75Axf4RwlHxViGFZLco5YzOVGeqPh6cFJjPkM12bka/GLH5
gsl06UKRQdA5yqcUvVAtN/zG961NOJVuIWmG3/FIEcqMGYiUs0jZ5XCBXt2T
I0vtVyRwASiTC0RWKsT0v11EKpy+p//fjq1GlegijPxMQScazsrPrdRnWXZc
wjgmh4UEH6O343f+p+QyaK3YewqeWKKjd4PKdSaTmQ/FqzFFfSywWwQIYvgT
11/RA8Oo4s1lbQzMROsGebqAID/h21UuAXoLZAX0Qdt81+afQuvYzPRK8z0j
dbQ6snA5ml+HAKTBC3U1NCcNyiCFYk5xkngX1NmeSQrd6oAeAtiTd5Enzgw1
bCksngrHb77eoowfDjKK/0sZAfSGumMBlLCjJfbWml/WgiQN/bQjuWG9Hbde
ZorX9bstSlWeZtgpMAt1gKIiJGGG8yM/kfe/dS/LVPlQl3hstD6aRlYW12Ap
tF2uw6lrc+Wino9qyg3/zcSRbgROdZAZMcH7hU0NAKLs5eVVEwnLh5uKG4bw
vjhEu3zbZPDBalxdaH+eDYdjYOej7kLvOasvCGjlDrXgTNqvVu7l4OhPE4CH
9zqRpb90nbZxzFC1+Z8yhMKspmvOygXjmlw9q+NFBjQDgb39E+DrB5oSDhoe
/Z0p6tokzR6Naj7znaqihCBvIGQ+zGH9WnGcSeY6li77BLxY1E4l1d3d/1LM
L9lKoiT2vTtXjhkISsmiKA7whAUZ2HNQCaGUlvlDJdvNKcekIuLkjnp5io6t
NF2PhWMzzMICSNXVwylQ1zEwv9OV7TQEa9HsgiytaBjF3/su2qE19IOB4tgb
R0+MkikOsSLT57i1t3S7WmKNOodGYzhYavC+ugY/Z0wP/Va890KErxfxomur
AUsZpweWY+VwClLkk7JBAu1VrLbBolSGU2mPhTdfs25AanTmDGmcOuv531Ya
0/s5inLebfZrdvU1lCx+6pz+rOAeF5DnJ2aOUN4KxzApOY1gy6nIGm6QBTf3
wxM4A03m19PqydQgVJxpBK4gN94Xcj73mEN/jMp1/+kJVAAM/E6o9th0L9nb
o1459FLBIDC8OSsQOvBdrjVLhLl/8hZ+rPqjwcDAlCCTTzrA2H3e9i0vfrhP
00BnEZHsgP3ILGCX40UjNHL68XZScOHVPsFweTIP8jyHsc7nZsiQVdbcmTw/
MtRx+SoQT7rwwO+J1xsCRALPj2/VmGKBktUzAwPp55jbf4xfaEY7ZBFsytHE
IvNNAEbmBpgZPHos3lTep9HtizXFyJD8Z5V+lIbYQW3iqfaD6JW2kddA4HJN
ShSapqVv90f16ZXChJCF1uqwYc7mHpE7aQhAc/ppMG12VGvClXQv6mTLe/oc
o26MxDcUJEzGdqruiz2BHrUezK+PmCHKTiISyLLkjV77nAwpui4fmvP1gKWJ
6iaxXNBBr7sEy/IVCRorKmV6JDRt7bS7tCcKs/bUZjl18Afe2CwwM1TM1stt
OcTcrfMy47nzbQxxUjHhp4XDQBDbnRJkJfnEwg0anUTmD5IDrm/oiNZAkETV
J2FFianyZsyaxdi0unv4vcjMmlGeNDH14+YHAOT2A4TmkCuh02QoMvdad0un
Zc4LQkkzPvD7ACHGmo5KcSDSrE9K3QmZDBW9Unu7T6CwTN4PdqQUxx31GEQM
xFRMd4jFuF+AaXyoul59ETJkrVjcOo7VFyGG3BSwoER2J+uF0YAbJJma7dan
RQk/d5AsNquzXE/TK8qw0pIoC+N8uBtm2Uc1V1P8C5NAP00paOF9GRzon/R/
hRBb7LckunulcndpAnoJflrPkLYcex2/D1UZUMnE6W0tGlVZgnUOzzanU6jf
sd3zP44yEdvpjWxx0/ozjIxUggnJSIbmCHZQ++7/k7iFKuo8Iy9hhHgI69tn
5ZiAfQiyR9qd5045NVHS4nFs2a+EOTFgwJUeNfxuIqixtuNIMOFvSxzab+gc
JxtDJyQRNXr265VVDRx2PwQylfRbVLAxzMkWOZJs9HQNSnw1PEiFIYRGQVSJ
k/W9k9ZySSGst/EkouNME58McBq8jPxmqSwelErFGwjjXTE2vFxsyzZav4p4
f89/hki/YNU1jVbQZGi+le/KhqYCwIGB50vU6RbQGNBFfEM7QycUfE9vAiAd
Zb962QCvVSBP93078DGpUEqC74/4cy236L01+c8oMztusOpIRXVaLLe9G6cU
ocInEbQoweDOtnvTiVsLe/iOH1kTzC2GdtkxyK29G7l2rUV0bnOHCuOzftIZ
Gy31rqXvIQhqzg6XlFMtdQkL2ltNEYZ5qF9RfAFp9fQCW9erb7iyWdD14bgK
WVuspFAC0JudEuJL5jE/DmwP0zfFqp/ujOBN+pdd9msi4B8rq/mtx1xebehN
kNM5SQE4ZI+MmwgrnADAlvqyrVsNT/oBeo7m/54g3+LmV+RpE5xxrcCCiTSn
JINjkMTb+SFtbYjnhVCaxHFeE3qgmKKT8nLUHMxF3bnuyg0kbp7d/AhTBysi
8vRWlUd55qcAgn7z/muOkz07IhbkcdlDJ0nE3zxOSm70cMX6wOJ6aVDSDt9p
yBxMMVzzOMTafmiMP11ep4BH8cj+Rd8db/5b98rl6Eavu5oAit+dwZRKXgrg
Igz/tpEN7Xhgb6/kG9+4SLPIN/fDDXikcrldlhZxC0GdumdMVbGNvyKXejYZ
AW15rGMxFQ+zrUhZ+18Mh/2MnoEQUIrxnz05wc4bwZkgAsPifC/3/ddO/KaQ
7eYGnDFnmN3MDy7BGLnI4vL2GogSq2JXZJ+y6O/fWjhDoOhAiXVrcHrbH/gQ
U8khrd3RcQ9Z7lbLix/XCQKJ2upck1SRev32M5J/WVnFYMDpvjkIrI/4TNCn
3Eh8nIRByyZKIvHmBPMF/tEVtcWgAj2aiMoNZJCrqHc1HIWDyaEk4F/AHZyM
uddbk4LZ9GSmbbCA6G4VExQJioeVnfmBhDHpj+sxme51PLYz9VMHe1DpAiv+
wT7suh1Z9hHmhnNVE5Ev3n8QyBq3eF3a+pgfV7dBU+D2jX8ZEQRxvan2sN6l
jxD5pJmoIrKWjsWNY1rtKnkNzEmg65gjtDtoCeb8es/3zBLQOeSnA8Frt7Qd
kxxqYNgrQqoJAGxjXB0+fCbg2wafOg+SZM0Y5DZa9lx2OLqaSihSSSJPC+C8
FyiWGU+4jWmE8u8kbNu1rQqx9Kahy0uC1U2WFRL1vScXYvgBgXz1ohtZPHHy
g6Y7z5SK0XUO+CU3dsL3Moo2+dwMVcLhwinDUD4eh+1eayO8+cJkTxPevZK5
Pd1EAKC3PtN0eLWPOGTsjuxiFlwbjD73z/NBUvz1YoNdZEKfChdi/QQ0Vprb
3zka/EjHRXKnjIV4wowJFvLscsHPoI8QqZxxyp57EfN3LR9oDefWIg1IPZx2
V8UIJrMJ5GhSP8h6PdRSHn8TH6+1pf4Lj9WGUfsHDfDKm+U0MTTDEqmVhbOs
ayax9TttnRrTxOlk3KbGNJYoucRr5qJOSQpCDA+6aN2KO7K8CbXtKyWFVcPw
9pU8KmcqBRXP0qUEqXtQKWR5tQ00gvDI8I7oZ3w5Q13qHfilVzSjAnlbkq+B
0ZMPaZs4zRgPLaLR0rvlXavLyctX7JqfsjjedSOwAiTRVFgiBCAhgrxLUV+S
T8tBDEVgax5Uw/cQa7BJVTYXuWE4rhfqKLOV3cyjom/hC2xDZssCbATNTdd5
wIItjS2Migv81MTOkmp1FymcgLB1pyQguSjtmgdKwwkdF9geWN9f7XMmjGtl
U1syvm+8rZ8kIJkyK0WpPHq6cgJBtt7h3PQlvpG7SjGoF737quXZeIPWwX/i
27LcrwgnWlstwmipg/XyhRgMBMuABodikZ6OkmNnxqZxdGfxgd+k7rIF3MPr
9l6L/I5njNFF4NhQpX35SeP2jzoeVyQTq7469NDCLtEG68aUiWl7OwxAQGBF
NDA9alJEp2T5daEAb+Q/KeCeYGACxSUAmglFhnFTF8QcNPfQh5ftFSN9Duz4
4f4ZaB0EbwJkIb+pqfQVo7jwmZZkjn8Xm5M8mXSeccTmvvNvuzDMd/nUoAGd
meFY77f9PjvIkWNXrYDC3SfyH1uXy3VMtkJLrA7AE5VDKKeEzt1SyjylZD1d
mYtBUIA7Y7UFBh0MPUE+QYNBi0es8hkYGj2kjP8f8ZPum93I5S1NdVEzswsT
BFOI8hnUK3GLPQHx0goNDabtUbDmf4rqeXCK54vomMSR6uwEFQtXEdW2Bm4D
jJre1sliYVuK7z1D/SF+nfon5NH3bMcxjZ1xHMobTIrSLefiYNGXirSMhHMC
hCCjXayhmxe5GI05LwfTuu/cYpbM0fbJw7SOnLs5CBqZAPQ8Np0PQojwn5LU
HCQLrQyUGzASgFbSgMCa7fDU3KOWIwRGc8PZn2HcdAjXKhcCvyESQ6unTYd9
6t6+Zf4tjGvxXlYL32zHfJ8LwP10kL8n0ACzjPvBjMI6GzfaWUWH1YTL+PVW
qxFh61a9fllKVH8BqP1hA7uXAIUpENBCXI5M0Ygs4/onIMaluxFKaetFUceJ
R2o1bwQ14qU2NLwJQUa+q+nYcVj9yFmSqu4ELQCt4z9jZACkdUvd3eCKUfXL
gOgC6PeJpbz4zdmeA0TK1VPlZIsIDZ4AFoLhCB3nU1uaopQUhZbXGf0nYOnK
QFitThHNCl74rAoFfzYr3YA22BG7A0tdBc5AUQ/ThexVX8ZAcbIfJzZ1kaBI
g5p5iIQDzNmuaGgAvGBEA7TUYOWWZykFCcNb/1E6mp5tsS3VO/Z4AMBs+xb2
jgospSw+habwb+VfayrAfZ4GC57UQk9WcQGNvB6VlDIi1usrbmSUQULVBdPm
Kr2t1phu+leKJScwF8FQqouKkIbjIBY72yiXXbvjqUfhKjydZF9X8lYKBzo8
+EELWl9TH4rNCUeFQbHRLPoRUJ+884B22EnQ5T4Aua1enFwhwCD8xzVVgyxQ
o2eIBZ00GGoLf814Enz8hviYlCd6OPX6+Qikuuqw5tM1RvJuxtoZbtCXK3Jn
h/JsQKPtFMJj1jDraYrfxfZfSrNToD9UxOzPQyUSom5anFVT0zM0atHBJxfI
MvQLQvLmvQ5Gr7782+mg4RvRAjNMWU0AySOl3FXZYoaAqFhmzl89t0mV74xa
fGIPcsxHFfDQ4oA/lcOclIIPxkAHiU2g5n8evW8Sjyo/bz916yHuO6pMeSCK
GqKhsnR5wPHuWKzFfVpmHqAUyrHnlyeMgiX5YfkrQRwroAEU2wCj5eeOpnrk
nC6Z2Cu2YkeA3TosVpuOrjo3t0O1GxmwRIR4H/BnqmWOKlyxMA+eiaLLW6VC
UlVKne3fyy5cf8uQyyU42cDURJ8XZGwjalxYceP+nik/tCS/fASubgIOFmJl
qXz8LBMftNQjNNtYEtOcwdeGRFrJ0+03w9IwF0W6zPBW8ySdHy4OzI7idHo7
lseEI2AVcKDqr76X+30gkWTxGCvWYZdlR5HSEVtVVDGc3myzQskUf12QB+4V
WLkoGWGsRVRkLEFGWwPEBv8+EYX/0nAJIevi7dcY7t2zFmy6weroF9z/gqtC
OiYABIJmckgTvPm4S0Gi39B9hlWjI6MUNdy+XnPQWM/rCnwrWnwHY/7U5epp
k34tPfa4SFCUJwWdoKhbu+MPMIS6MsvF2cVyKMqYlrknD83M4WB2a1C21xjA
EcvfwZOBlc7O05GG+GakDd2IBIW5oTZDcV5xlZqxTcZMU4nExzviJhNuxUqp
1yOSkFe7CJxTQhMy4tH/tBu5rThQAS9MHsBz3LNJDBjjBJcwwN24kyBnDpcS
DX530vq7FIRB6tvAUGwkrZSzs6hXR+fSz8lzdoPMLEN+lTDMLRbjheEOKIk3
bHA+W7neewr6O6a1DmS9W1QVsMIFQVrbXGcd0VDw/mY3Fv/FuCReYuRM9EyV
XSFD3loePHkYfsw+tiksW3s57dvmJ8rgi6XFCaUrorCJVapTzOAT4xeVYKpt
FkkiUpPnedx5BTxpBU8StOuicMWuQryndLeMs3qhApTACZ9DYjZ2ks1EAxWc
v4lLfiD90vyvnBn5m97FtmBAlPAEBDAuP3CVKTSlncC4c1sUeAChJMtjuxHz
uohTbGsg5Rm55jjT2UQgxVo5F6RPPAaAPV5r+JB1E7znfNUyO4nGVybdIl3g
uwXebvbKB2SQT8ufw03uCul8w8e+Po+FaQtaxB5gtJ/Vfvm0126vjpjNPn+E
68aafquXi8Kbvv+wZ3izfHN+KimlLkpyllVfgbO6bpnNoCX1fPafM4QEJFTR
i+EcFZYgKtl93r9/t1pXbUUAOt5E9cjYS7H4zunpJYgm+iSwbaWnLAOfwhbL
qSo8m4jZa0fcLhp1PCHSWkgXx1q9F+NU5tIGfod+69YLsodnEjvW4akxbHxs
PrGlkmHexKqfWi4xZyBDurYTtABgG/dMkCtSd5HtLcPrlWiAV6YoiTh0F74p
Jbkp3NeDLrDwGUJ39Bg5y+yk/uq2V+DzD+UV88Ebor8pWrgR+93Gt4zkJYWQ
kyKqKILwkranCyRB3N7IoKI2dgIIDIGSggcHkURU85Qn/MRBPI3YL4g6ALhl
CrpcLoPDg1CiIv8jhj8DX5l1wJVit5fQnV+RP2T/fg0e5Eq6eYKj7CedEPOR
09f7QEy6rbp8Cb2LixKbgZ/g5/Fsmsypc89a7JzZ8tLPD7jcw6te//IoI0k1
Pb7UT+AIe/ye8sw957hS97QIHLDYx7WtxAhEFgqcQE0QmMivtNM6SPujOy2j
sXgzDrSw7o0XmxwRhXQr3gjcvv/EIY/CejwtiGoU3GXFKm43xb6h75y9dyzR
JHayWJokQU/IY7dx4NWaRqjmXPrHcd4nBoCxTWJgQUKH2Gegq4VQCcYEjOyL
Vy5sEumO44qd0tiMDU5Ro+nBVLG+I5yEd2mfSGPEB7FWu322YEjlpD0sgG2r
C85LAw8/h66faG6WRlZ9HKe+yhLIaGMVTTQOXXmOZJJn8QjnF8lcxtk9G6/Q
rR+umKy3B5q/XzFs4YsS1Vap82wQG7unvfJ1pnS184UBVSSJy1hCZs5ZEG1F
SvAHMu2Fd13BfAUwtzbgdlbMqyiUmofnIaEBG/6SOF6y2cZdLrd1gm2jgBam
7Ejw3XtePFVDknz2tM5YdFpppJwmi+FEtXsKeZzPrruMTcjbjzXLFcsWtO1G
jbKMWmcJ+L4lS5qApBd7RqWpiajeXR0CMssQmWFVqu9eujxqrJhyiEAdvngA
5vnhRYOMvN/Xmbv//pIjuHtS2wrFPKKi1PnFHsNvVbM9qelH2TIRka/3JKhR
4fOksCTcAxSLxkEuUa+XgNhBv+XIRnB2a5Hp6Lbfbc/Qfq2DgqXnIffpMIwC
YH36FNq+N9Zq9ak6C27ZbUpSRq3g/4lO7HcAeYxBavaVc24u1//vWNCtmNZo
o/eg/YP45mzB3h87dUA2OEmsrTh4Ed0xZfLmcJiikDXCEVokwQI+EzFWlQo3
jtwCAPt5iEP2yhaXbmXg+JnlCz+lqxdp9WFlcirzDUL68mvfhDCRPiG+RPB9
CzgnibrJ7y3G7YJp2Q7JhpPeM11FaauEGd21Xi/4/1pLEkddwL3QavZ99qY/
Um5fblqrrrR/z2haU+HijlzQUZBuasX39mXLTUGm6RcZsLpjKQ42a+naSAvr
GFD1pro17HGFOJI5AQTw2HGmND/0/KLhGw72enFJyKImOIU6Ppr23URfCTkr
tZIAo8424V9S8aF8cqYKxHzYBYsV9n35jmpoITMWBS2UKawY/4dJRBEUdwlF
G3lR+W1x29Aaz43WR2XCcr/jtkZqhfQIjute6izvlW9p0n9+qujE1otpab8p
c6BqQSypRY2cFO0v1mq9EX7l313ZxNJ2Q0cl446dI8VmSHHsB+WXB/JjCuDC
Fdp/OzIaOvd8ack0y0b3cHXUNUPoBFTonHBPWuBNWs0SrF1MRaitZgCnSIkf
CSb+K3OTw8cdxhY9DibUfFwKTJymUZh7NTvNima6x5U72rgvQGw9oX+KRwdS
MOQn0nK3DN0WPg0p6FIpSmBDlGP3xWvzkk/T9kawY+3ef1qsozMTGtyZopWW
1TjblVkXW/S/Bc8VoUf8FeXcNnxUdc3VcQs8/6AHQg0iKJMuDpssSKLfxZGQ
oogj2hqJfmeZgZMMl7lXaDMhd/J71dBWge/RUHbsaw4f1sovcZ/i301WO/xU
JzgnFqekMiNwBBv/0PBdMmlooreevOpUT0Eec41kzRQrDsonsOo4cArvVrW5
MpkAQXKk0T6bT181FpKmPptLVbllQjm4XDzyxjvw29ioflNIGnwJW2zHXiOW
IVraVC59Oqel6XfBtq8aDC5dP52w3ZRODzhGhkdLAxeEdD/EDOc9LAGjlqeS
nRwgtULvzikUgJG0NLAyLBA6G11ZsM/4K8Uhj2d8waYqTSTWGKCTFoRRem4T
nR2Q2sqwY4+E3DpnETGcT8+T4bRTY3rBBiYrs2jZvdYiaALJVa4VNVDow6z2
OhrklRZP/3R3C6MNfIDiP17b4gPD2JobVzkVbKtbdrP8bF3+veGEzVrpGLrG
NYKUMMZCBiY4XVvgUHCmKbuOz+09cXQeMFOOFTByb1zbL3JpmHX8OB6j3PbI
Px6opTFfZ+1Gm2Ylkj8m25NNzEeYo0oFLp/2BjlCt+EEKG3TUKJNXDLzB9ZS
pD9MZ2IP2eXptTGzU/2wOByGy/LLKsv/XTd5zER6HAslAmp80wQf9FPX4UNK
sk0047azldtTk4UwgvO437oetJgHPE8UHefb0FI5b6pgNJD1/ex4OMUwlHb4
8nb/7B8UFWOOm8HUTOYmLg5Xb9fKQIFJngUHIq8NUrxv3WWZLo2LHnMzlUqG
bun7h3xwSBK3+G5IpM+b3NxQFOjlHxskrX5f1hXwVF+vBQ0HAWNHn20VMztR
evwNxY+m5ab17Sq8UrGJ9pZ9aYt7w3QJYQIM4Lpdf2YzAbQYGidJsaAWJ+wt
HmUSLMcqBXZw8X1sHMB9OvcvZQsrXi+NbabF/og6jXgeAyS4y8y8vP/Glyz1
a59EebyzrZzu4giGBeypoLo4wT9tqCY0xrW9b4GTI75yhp9G4yZz+8u94xvs
95oJxv7NZ4qu9T8rqJa1EG1Uk5GrcaNMeY5n7R/hczsQ0bzew5Q4nzZnPv4H
ACJE2FvjPjdQmz05GmktSeBe4U9jdRpOnkS2czBZbQKD9SZNW3bSGM5J8wjU
sT5CpoFe+m8+RmCzOv7Z5aSV+rLZliAlTA7p6KlM7etZI95SiLqiQocVbB38
6wM+kWiGEZLx/CytI5l6PTsjSfMdAHhzNDZy2fVTtyVP+MKxBed/EmY7yuis
Os6BZpP9FJlU3ajjeIeIV1HU08QMvaDr4UdTt1NtpLRssqY4wTI3fM8U0doA
nV2h+kA5FB/kXCPfJBnIgUMLBGuxdjGPbjnRsnRdXLIiUeMf8VCMMD4DQXfJ
xYQi2MnU5XedZo2VlacEfSx8x3+7QxBfVPez9e7A8RhujBWpKuKxovDIGkcn
mmyK3y8Dg15Nne7WVTARYGsNRAS+u9MLBOtPZ6tp+RFweQkGeKKj8QKM1lHy
LjLdXb7Y/viJZ5UmbEyCF0d6uAg31hk8RN3uGz/OmJuIbleBUcy/XeBU0uMU
ouTvVvOR4WKHUJBP0nwQST/JeLrjP6l/p0TPl4Ze9xmyhyYdVnNVUNK3P0ft
FOGLJOQ8KAHnmQGi0zK7Qbom8DQcs6rFh29/zvHDtbhI1axXOx5GXKK3jk9m
olJb3LPgUGef6VvYaLc/jQIMFiAPwyCU/HvEIgylMFe92GLi956FWIkXm6Ej
bkWQCRuOe9WQid33Nt5OGLuryvs+A89y9/VKsupLo2yCukbSp6qeudkYQ3FR
CT1noWtWL2xdLIvefTBlIswwnhzNf9NfT7ydR7Lxb1N7HDinspax4r8FM0gB
xIqWapMtzq20g9TkJ5WJOfykVEQse7tzE/wYOEw+PuaXQqJkFsjbMli9nbx2
W+X+cz6yTTZggQYF1Cwu1oOQFm8MuWKZD+mFn2iZKgqjmkvCITZnBYFeGx2s
DUULu5LbPw8VeF0IKyzM6ovmXU+bPY05HjQXkT8jkSR+1pxaCNR0iU3BA+Lo
2StSvw8pJZbkLzyCUN6l+iPc2i2jIUbLC49M+UqTD2tb+gy2nBvZEFdX/Y+M
Rtj17YF1NTx9Ses66xNYAlIijT1VyRqK6O2pbHvxNJIcqsUNWAcEeVNOZVnf
1/8dceJf4HrxTnlKAZOrP8U7MSP/HuheWqRPYKKIYUlKxLgxMOsaGu/CWo7u
qEZk55Gdap+B88XoKBHfQJ4t3qtD2t9oIc7HYbP/Sb/VIfNSAySeJQt03rqu
tbjeTavHIfu8oyVLPUUUDwClSl/p9pfa1DIth8/32nnSzeqFqjxvrDoeJjaa
BRosD3wFVX/+QHOQTwH/39eTvFvpzgM2VUwAtRXkv6qtb17lk35jo3pWO1ks
Vz+GJ+lP3x/2SaQLx6EOk4WpsqdFkngoTM2qUyJnj7TfWZUgjRJi9coI+SqU
VsJI3SgTe8dCZQw61ZxhBfqEbtbkfSkWFXzWvGFMTTFMkTwLd4m2J6D8hq0C
ZNcGvYYme9VlxDpBO2VAQCnTaJz182sC/HzA2QCUL6fIxVgeV2iSZFzUFywE
iwgSYi8kfsoYNLe4FepXjNONhQ+GhBHRV1lN442Ni1QhS6rTISiYKUJt1j5L
Nwa9eS1oBjf7ZJ0tdbsOQ3b7LYySo4q9XYwTdKMDFBLvP08n3mpK40witKlG
X7VDEApcgwqwZnLvuQV8t+rrA96Dc53uoTLcO4p91R3y4RQfK/djQPoZrd65
B6HDYLRyYqf3W+Tg2qnBWmGPLbH1/+Yyd7d1dje5Qlmut6bT/D6M8pgx9bW9
w/8x2bwW+gxaDvsbGiLIDvEmQLyxZDXJMQkm9gHucdDY5SgTt2RH+r6WD1QO
nLdRYsLt0ehuXVWx5bJFlc5UHMr4IBhhLTjf0+dqsC3OvMJqwnutKaDQ8ofX
Xi16LqefdLd6uJ5lB0Z3gRFK3zo175XwWsf7q54WslRlSsYfaFQ58xbJBvWJ
bK3JmWcpaQ4vMJLepoMCQtlEKAJ9fJkvioKjpKHz80GU0jY9W94iN245WKrP
yr5M3a3/xWm5FAK7YfX4LqxjxLNxsW5vgQmOImkarJFrK8mwkKsUgqDZgh5z
H+taSPwO+xT7OAR7EcNnYUj8T1vN9xCwiuhzAw8qvbO5S3emuZCf8v2NL5zw
JoeWmLeqMVYcDE0+o1wzVRqxzW6nQYAgy4jSLRzwRPd7j//DByXJ7KiIHSzs
g5ejFaUkyWm3ZWMzz+rWfI/b+hZ54t+vSzakhAixRzrUqXCNaPGEwpgxNm2D
kw9421qXWJav3bdTdqTPANU6NJZZ71gvahASw/q/rZFfDswFrVlGEsq+jUOg
A/Xgmvgt7NCrxcexFqgAEL8vj/VSL0MWPyAlBYeg9dW/I+9z3N3QENgQB98+
/+2oEvhN13LfTOeCdr4R4M/kLLnorGuzuz3cexsx3cyZvuywIftrIxaWZznB
1Ol1++q5FFjcxARZ4BVzWG0AExePzEqR4qJSR4ABtWlBTdXCbfOBgkq8mgf5
0OQllVMmAZzIHvWMZ58czUVtBn/wMD/pfGdwI/AhPAEE/mVA1QyilFlECm/D
IUttsjD3HU/zYUeyqpm4YeWPMwkbQTKK/F+ZpqB6o7lBnVjfD8LLegL/YcHE
MbVcOvVBCncO9NmyMeftdwNSE/7/eID9yBIgsi2OnZlRwqQkVaI3NqYfvCLL
9fPWwWLYY2qiqovTltifoDKL/NDb5JlhYyMPX1JLROgyZpV+7QnR4/txdooz
RD37Ee+rt2AjxgNmwAdRQOaZAmcR/9DXWP96N+ik/O/yZEP0ou6SNKghqstR
VmzcsMtyPpHMhQ3vq3mQEqrqY7WrTFlhBTP8Hp4Kv4phpoVdi2c6nPWM4tI0
Bm0vUYYKSQZIzzu/Z66GydzcEzRHxmf5nG//dA0I8RMsz0Fegf8mdLJPi94y
fMA1dJbmfBAMfXomsrm8V84I7NOCsLj3LxCWHcbgZPIbBapelO49XwHiL1DE
gQr/cyr8PE5GyXsT64JtzI79RwrnVvvkTcGd2SHDZcMMLGy31THO1apMTNC8
LjoNy/D1yLi1JHCZJgrai5Ra9bhIAzmlMsRCD4NYMewoLyI0PuwKfUXGKj0o
YMbVYOucYOkvmJNwzbNq6YbZhzfW0XOZ2LA5YOFA4QRrktG5oCxoDWk02GTp
mU+nRkF2k6QSuTtInL7YJ6WQzgoI1245X/OC8BjZpkCtTJzjJ07rC1Qt50H1
XRz5Qeu8NDaBhQ6Gl0PioUbUjjBo7O96qBM7sGQC+en5Oo5dwSXhMXoauu5l
chgUYKbidiy8wlI1xDUCDS9Jno+JVP4pj2xK+TrtihLVuTaowO4CkYTpsqGi
q/Ex2zeIt7NlK+W8abhznzsVd9up7U3gEcCmy9zAhwdbFF258giOIWF8wwdL
CZRVjtexSCSMyFxKNfk/WTHaV91BjJuMAMY40gTbAjj+KlzsivuBJc7GTNL5
6EfOCX2NtX6k+1QI3ZzhRJXZ2q106vdPel9E3gLDY9nv8zbnTwuWUKW8Kx1/
2f/7UlFeZcmbRSCwAKxy64WsfXcQkcSlbTg0liVESo30oDQ8bKMdvvutyKzC
klYlsKNaRzMHQZur0tFbRD70sUJsBIjQuycJSVVnJbKWiZfPzKmX+jNFBjTn
p4NH8Y9yJZfJYBj13SLnri5B/R1ExO2f8YoKo8fTCBsRKENlWILYM6chpqa8
h8lZwvexo1KQ43CMpopln+LgVNWBUwiRJxlgviwQ5x9tQNvJXSp2P8XTY/sD
k9ABw26KJ9/bvPaNBx3mB0uLh/wDbL2UxNIjf9z8VEhNMGr7S1Uyn6LJulu6
bzQO6CXto7m6BhMw2klUZtLiMaOHFaRGbBjt+1QlM9fFNoqJLM6GBnAV2TkU
B4tH53DuuqwvF31K7z5sCt8tG0VvUOPx8apm0Gf+dd23x4WGRm69pViCMgog
bLSx12J2hz6KqockQdNFUEl476SlofuWAfttG5ZjsV08DhQUWesvPDUw6uOG
W18YuFS3N4U55kYENkosf/uyury+3SzRvsgAL2Z9ee2spgrAJVaujsbf8D45
KgFG5AV1L5Z2mjQ/8aIiNib0+UGolHtMINnjU2cjLWASm8D6YnN6eUUr0n/b
Hao5NIRlUaoCt4sXJ3pS193h6n2pujwRDNoP0HDnQBvkAmEUfETWeuek8UUa
60iHqNwdkz8YNqin+RiDj1MWXTKjChQqy/tpVAPkInKJxCoaSmhazklITm6P
ql3pHKnB4XfAYp04kjavdWoHIIlQiWQm/eClkp1IXoMIzjuIliAT9+5T9cd5
gdJEFuUsvgEC+DQyTXq6JyRxz9FSJs1pW0CYps8lbdm99B99/cXFKLa11e+i
5IsYdl/WZqV4yA56KLb5K9+Na/SNL09pCsx578Dovx3S8p1/EInYBdcPRJOi
QfC2siEcfe2jTGL5QWT60yoP/UL6koFSdrRAi0N526q39jFdfv9hSWtQ2tix
g8/5qsZFJBJmFHb9cIQSlOh8/aiQH+ySLQZCjuwCQAVrhodFGx7WmPHNA6bO
N3qcMLu5HfjO1Z94YHebtZvjC16Wdx9IA4dbC/PINSOIM+2NSpSwLKzrjCmO
w8W412CZ7rVGyXoaI/hlFI8eqBtIt8SCRH/9jzcoRqM3RPmr82gk1pHtRVzY
1+A7WxrTR5uw0du0eNXfHMxOj7sIOHFpn06qKdR5+ZVcIp7m7isOEkiXMYOg
G2YpPUOY3L1lyjI3Gqe9AZ1P/0e+IS/sUIDSlIM+11jfnDhaNmQ1Q/ayuoxr
1o4dxroumgGkI7/6v78L5BnraeLIyRHpYWbYSA5j3PUS+xNx135hW0ws7dyt
2gXickgfjh7ZIw6O3Srk2XAJ/B5j6MzgImQFk1nvjSTyafkhhxCZ6LmLl/t8
5Tpc8Wow2oWid9G6PfCqCdxoaDND/IulE3vZKQxx6A7n5ZPCCarUjksgV+nz
i2NadaINXaSrYJqZS062axbEwdYkcuRWzgwLEZChYCdfFtX247DXiIz84+o/
thx3OMpDtfnqmguxQpVBQKGRtXVM0i5Wh18FI06hvtmFCO4flrUmz/gEyAFe
nNQobGWE4arUGfUAZ7kZrEUde3riUPTxkqpr3KQ9IInSAiILq9vzHbMJaHk6
5mpMg3PeavpKSyqW05OpAvnC4savZM0MvnVt1rGIEWFdcdfzJAnII//BaJIB
jGJ+FahCZrlQx1nxQFfOZffAUMP+oW8C9FNyA7mn6RALtxnYWJWx1jOPmm75
vMhHwzrE4ONsmCxgqJb9wg+TWz/bHCJZlkm0qtu7fGweOFEXa+ztkuu5kmbn
fv9ozYJd8eiZSO6xuNOVuFNtwD27X3VkC0UJeJpC3ScS89oko0GBQc3BIrcp
xIqBTCMZOZy+bsNVdn6gcSUj2XGvScZdXWSbvIF6k2E9FJ3tg5DzExwazztD
V46VfZbOg9D8HqbtnsvGbAnAUbdJfPJ+hKJvTq56gpdSdZWt/jfD11OfWdx8
B4TJEzU87xX5DMDzYx9fKYouXA/ugnUfDGFJEQdaiazVCmA+04smurA6oWd1
fOlIX6zMZ0xqZhMZTYOhGi1F0Ep5gzYTWhgJ3YGxSqONPF/mcgGFw523qMqh
JgHILibWmgfLpjOBKUPqxN39vPd0/T6UTi97nQrkLQKgHsVZqr/vIoFD/r3F
CNq5YfAzyzQxYcnC8AB0C0JnRKklSlEiFJwHjHHX63tPX/Hu0PEGBSI1tar9
nJNfoXUNGFTxN9R/jP0BcDw8HW2Uy8A5YbXJNXw3xyDIpTRGE8UkLWDe+71Y
V2rLe47KeqjyLZi6xk/agndD5P/Zythtc15uojXQALz5TBrveM9zVcBMKjBq
qeT8BsL33XnbkftwUWJyqdEsO9tTqJiobcVb8/YrtmxnFub9NnTuapsvVm7H
ctIBg9JujArOHnOIKp4m3g12MOYUpF0BxVKVoffTFzdQlYUKc/LOQ2plkYPC
YZtRvT4EXsX0TJRKCCPiDiqLte3oGdyxH1QMZdEwWs/U6tIJiCMEkGJDskxr
usahnpmB2abUYcOpH62p2/Z+6VSSPefSIU60TmoT6/NoZjwcBcsjeb5aZvHV
DPg+VS6T1EEB/ahX21EKmxi+OulEn5c8X4Scvo7l+c6yStveKrtmvni/Bou4
BEgXd40jHViQ6gLmZDSanvyHb2FAU6C4B+5G4G8aoC5JAZgWz8MTOvJu7RPy
QeDeayAAZYWu5wCDLfu+tm0hQGaPXVuLRDZGKyZ3sRBDa2tI6lOPZXBRYVQc
O4biBL1GZCy0cbjks2/AfYfC1o6SSyuj/rngYBKDLUvHwN5cutbId6b8m3Pe
54nOcE17XveYJUn4Qx+4pAidfWlQnxl4rIxVKnHhwSkoDb4C6mpdzP/ZanbQ
Uw4BKndWtYqW6g/ftoi/LLBy6I7hmOvhYqXQWVc4nJkB9LuKD10b3tUfEuO4
spZCh2HJxM+jWbMNzMdZBqMuN3MaLm1eCvvEmsxYYlVwOxbr6LfyIwAMeRri
ombEXdyQjqJX8hECtYKj54Dtzg7+C7n7pgCxgydD88RcxH2Y04Oefd3I1GDH
wXbS96ivS6lqWRGqjd/nivBXwkSmgDc66/+pn1HC5fnXSx0TlBDglWH0FDzs
tZcWIyccOyA6tXo8P6ImXJ/bhRjyY8cA0mb9yI7qVnwdnv5161ypGzi944gm
YxBg32nxbih5NxZlfUhg9bdZ074NY1+rX2psElIUpbh1SYbdCuDDKPOwruBp
uF3f59aD/EJs6PoYmQf+gr8khbFOz4gIuQqqVdcm75g6bCLY3JY9yEida42p
+egBc09DCd/sifj4m8bIjHzmPvC0Ije6qglkYbJSVdLMtwa4rEGCmgFEabib
wIYxqTGLMuoYzdP2od2Gqdf7OvWD9j5jXCLvmW27l7jF8VPY3Jgt2DzwebX/
7+ZxA3Pm8HrfXo3GxsP5NxFr/c/YbD98D31fXAxpDS/QLrJUFNZpYxR5BdKZ
Skc/lYQQugBvKm96aEQURAyfM2o3TOpeceH97LcY84pZZSYbyt+R9HzYJwZi
UEh682ZwLLJovSgr5Jvg6RCg6e/pkxSAi+lyf3hibfAbAMy7zn+e2jU/zSQl
aEFah/22+KG9vIjFhmrUYosvHiFe+4dySr/g7eGlulnus+h9AJaCFvTwm0kG
dv17ytsklK0LU0FVpfGCp3wrbX9ki8trXOyweBFIt6+zNr6hx2x9EWvZinIe
JSSZ3lrEv2SjMH9EW74h3SV5SSfrTCgwjcaa212FIaPeMzCdZH0mcY6S8oC4
UovpBur85qg9KaiOYxXnp1p+d49DzWz0zai4J3iS3uiINxAV0F8f2HOVe8rb
NDwMgdyRfvWn6yM/TSsxjOp7lYFGerShxNtGeltoD8cWix5UMg46A/IATcnj
v+YPUtZh8ZMD52vBwHY7JhFdqxtCkM7W6kS2bn/Dsk0x75NgRZl4XqI7PUZ5
X+h4+LtoUN1KB2bsnMR6eaWPaIQWRSRgUynYXV3cyA7q6oOIea+Mo9ct31RA
v4u53G+Ifg+HSDXyqYqB1cY1Wc+ILKzPVmn4DRcvS3UbpA6+miv33b5O08fR
k1TH4fKR1Vu0So9b59GUB9M3sFthjSeSNjSeyZJ4XbgdBfaokJbFLKEXsmJ7
DAg+StNuMuxQRelbVBADnemPKd9NGoyCvwgvYVazY+T3O+MzfxItegyfxh6f
dUwSueGOHwxePYEpO3xI4jvFLZXJVb96kwdnVmOAqBdOhOXytUVFW5FS8/5I
2HCx3EA4Mxi/0HkMUC2EM9yKiA7QGUehHaP2sqIS/UzlUQTk9e8Oiif8hmFB
RBmV969aOqV9CEp7XWBB+DkZ6jqD9xkAeVL2u+AmrrC6Kj65/be0PKXxL6C1
9samhdsocwmCWteu7+C00z9Hu9OeAp6RxwgF/852ey+NpVacpv6bLt8hBR59
qxzeOCWD8bAC4K0cpjEmw8xIswCZoL92Bk5tZSIdr2WWP+1PB/MwYawHsApB
+3O+2f0LHgQA5kV0QdrwyfrVgstarM1JjaLOT05vVfPeJjpsVNNHx3UY+e0G
5lUI4O2+Uenb6NSP6/VthhzejarzGT8tvLdzJL3BWSR2CuO7NLqIZsC1eLJL
JMmz3P7UA0RFZPSohYHSleTN7tYCKLuZUjHDxfAIhn9GULqOaz9YRE8uXU/k
cuvpzAm8SOUh25tby3Bgk6tnNYcrH8kRoNQmjNXajj0q+ySJVuQqFQqQsanb
DyHmBnr5lrRC3eH33rCn22Yg8uVjAL1eSJLUWseWcfm+JQstZgZd7TyrWYxy
XUwTSYjLbx6VJne1oe4PEA8vYi3n4kq4n3NgiIxZaI89+T81oxLFZOWZlMSx
F/P0K1EcR+UhUVxrDpK6Vk6HiB3kJBuP3I86G3yrAveCApAOhYTzEdQUkZwo
FKuDl+pMMZV5Vs/Db3Ds1UlvxKenv39MnkMlp81mNG7dpRR940oGvl27hOQl
vlJq/NJNtVG0mrpUu15fzFt8mzXXynLgFFsY2rjj2ODSNEuDLVPZ634afRd4
+3nZCW9aXEzBHTcMW18VW02QPu8+BdkIsiOHj0H0w3HIN9JwiX/VJvPWsbUY
xr2IhED9A3WH5wL+mlgMhpaVGT09jlHMhuRDLVXGRz1zZv1qYT4I4vm45xJH
hs5Xge9okqm+wW3CvxU6xTnkJnLpHDEld2Rjc93WzoBZoQ7bTxrI3e59wndu
Zb9NUVZ/+ruTn1W9ijV78lvSJAw5wKk6ao/xFrpjpLzRhRv3dStgNsvt6BKh
9NMNPQk8nsuUF8VzTO5uKFcc8V78SBQn2ZJOr+KGJ2BVPmo8u/BOLG4wpJ4y
UtbG795R2xMd2TTkuSiJfD+QXwXPTYbx+Ntc73e4zgmQk9S5RVAbt894WvS4
GthJX2mSL7U21RWJnDa5D8AvS3zL7F5fUn21+eaqwo8jvOH8XmEo2OfITtyd
KbDp1b+8WjVEZxpILiyT2sXpRDN3CCqCpjLGPJCfvAuVpRmxELqHNblZdQe/
05mCA+TQBNlrF9GtBam393h2mitKMl7JVFH0DapV+9HpETKngMphxXdwVSBf
WUF5ZfRDiPyzNHhuHVPoIRC2LusF67NWyvL2LiHYjNDZmeCmia1SpQgSxob+
tSGFdGyBoTRm7VpQS/jypKiK0mdOJmx2llTDMsEPih1prD2t3HHN7rydH4bX
D/sQ2+6A9X3bFOdPXq9354cB2vhK3q8wXcj4npJYyPBAkca/8HVl/v3f1/dN
b1f6tXHrMZySmLbY31/qyY6Bd9n18TAZNJ0983zClnQtdahcGILZQw4F6qBi
98h7ansbf/JJoI3Do4BXgbRwnzH7QV8dtP6VANS7Odr7FqHB2Xheap1iIa59
X3sg8usEhvWX1+/i7sO14VVvNqAOShrgTCbG78BqC80sHJ/eCqqppAzIAB/m
yHLg9xdzRFXGYquEW7mHX7D7vuuE56PQzUflp7UMvqi+3c7NHccqZXgLVKxd
koqMvtIxemq3BwXCnA/bkCyZ0xwZ6NuS1rN5MBYoeY1yYmYamGbBl3g2sMpV
UNqVH81s7um7Hm7b9xvbSD1Rp6r9idGI55J3c9qqXxmp4tpAHXz7lW31i4c/
yMIkyu3hFVCzUuPb2X6qnlMWsnan0bZ5MT1Gw8ycAxNVjp1wo5Jfv/AD0ice
WCT71p0Y8KxPYddHaGxiOujkUWWd0EBwTrmGLpx0XpYBr0INq5SpAqkC7uwE
y/R8EZWcTw48S+ITpM6s9FUnCR9NpAuCav0+h13grOfZ24MsM2K5oj0NQXZP
Ie1U8TgIFeLJJumvkq71T5Ye53Nm8zAm6micHzlZdVH/54Bt+bGIeg2VaDMO
GkNWhBQBL3OFfA7l5HtqJU0GVE3wsoyQjKD8/AmfPICMhdb/apRTj7UH8bai
aaXCd9iiSzbEHtVxusdhEUxM1Jljl9G2xrxKAIzZcCDiZd0blLLxpQZJ+pRq
8dLtzMPa+4jjE2msm5SvxONiFNku6Z8hKN4pyS1rLVHrkPaN6D0tjlyhkP9f
eMpEtb7A7gUFzzkCkFIi5yMim787IA9PqkxgY3KmG3p0BcXvFw8CwJnguoPl
DDBcPnDopd7ZngChiwPjPhQDahBK/4+9ybF6bP4nMK3fxHiyqW9apE8YOJDW
4njJXvaUh+nQGgATZcqJC5hWylp3Kkfgccsw4wlBvfbZjQ4od9bIr1Pji6LV
uZdG8G6fhgttUA5rW8WqYf0iNA3CcndJ0XSy+k0er7M+aML5P5pKi7oWEo/X
hBu/QQG9wQWxAi1S/ETVEnz45F30gBuMNiRgXVUTcsVeHUIqhTiigCPQRBma
Uw83DzLagLuZWnHGObL/1NeqfPIAlV2zXzdz8LpFfo/ZW5OhWjU+ztA/Vwch
c9h2syvW2lRr+c4A7F6YloAlJWgbVeQec5eQ+klDHU4/mmFw+kc4iKIJL9HC
6no2xvZ2WDhsmieJ001XXHL9ewwNgxkDqGTWk9YfaAoLJo66BDu8d3P4nby+
mgFxNIIZTiu+PbDE+TtpPNifz4k8Ou+DMiVjc4dYkl05eRLuLm2GpivGFv2g
1wYpqmBio05HQ0Ul6665vR1vfHv6uoWKDNTiYuU2RGE13ePM5f3enlgCbrLk
Y0X2JYtZw3sd8/U+pY8bQfh4A/eOFcb7IzVY3L0mAoI2skC5PtMoCXJxCMtK
BUd4ujdXLUMk8hHpVVc1YTRVlmkhOAcjXno4/6p0kE93d8seFF+0eB2T1jH/
uJH56KxRG1Ivu01v5sxnVvstJ/u/wdFOCDOncPD9WqC1B3LSDuo1DxeGMTGt
x2zk2bBhtxUaAFGXNJ/2CGcZbluZkMzJweEnFbG08v0yLiBrSlHYCzrlSvL9
wMtXlbizQH7PyetCFVzb3481ymekRB2rAU04dxu4mu4W8zRKNzT1/UZVTlRt
YHfaCjD+pwlviFy+d31GcAV0lhjI5n4WB0PMLx5OvcpYNnZeplDdh4aKHLOl
nlfvrAmY4p4piBVnoT4jim67Hg4SlotWTevlk5HC/JBagZ6A4sfRRQAhL/SZ
UhIYWWxZW7P7WbWjZ3H6abBOy4Dsq/HYE7G43tzPKuVVq6yUow//M97rrQSN
ASJmEu6Nws0jSsriKYZCxwDd3E1S2cthT1CAvDfQq4/ou3/lrJN5SF8/zVN0
bhB3HqCf2n1mAKvY++Ic4VNp0favKC3Xox1/F/vXccIu0KIvXlBuXpmyzycj
fllRivmmjpAVWm806MLwR70k+USWyjGTE3f9jVOMFRg1DUCMia0nOlJUnDnR
THRQBh3bJFvR4u8faekdNfhrjLXqODgif6pDHHhsPUsV3CmLjBC/p3sx2jjH
915fIRpJR8RinPGhNRtacHPy2tGGifWazHzg3vXvIApE5KZzevsbLQtMMn6S
XTIMDDLc1ckPd+1564evp+I6egq/oh23YfE1/vsh/dGi3esBEQKk3vS3T18p
tRJERom5h7JElyWfdzyVah/Buye5SdVIVeDiZi8wplii8+I2oWakGtq/96Ig
hOfRRx49YbF6iWMRbc/lNINeXa+UbuwBcgatikDTIiI6jXuRYyrS5k5vfG9q
g1KdkzyKCuC7NPID+X5uySoiL5zP/nYEEl2uknlQcTlqnz1ciqKr5IfcLOp4
QrKIAbhSl9a5Zq/22Cj/MQmdelmdS17MMeDeIVzKAx8PLu5Zmi2kvTbqiaF/
MrM4rkoxMPFqW6w9S/rcH1I8s1yyK8FzCSCgZ4/6+4qjQRkisPISmfdiRVA7
h3Kc34qSTyXgUOEyTvu0JJwDqe5A15mWA8B5rvMpMO6uVJZvpFQ5+TnCY9K8
DmpjDpVuDP3zcOHHa0oBGYAg+if/1ueBTGwqmsZhNxH37VoOUqGwD1SYyXMr
G4rIxMAh9wsr2TM6lGGK1ftEBfuPM9HwHb6xddrfCs+JjZR5/aYJmeE3Snpo
ttWd5tnPUCyou5S2u3WiYjRLvaDWPveXU12kBzZsLtKtnePogr97cHPdy0UP
fsBq1elzuHf9Yz7IyOi0a23eyDHf62xr5cZPIPN+GpALnE3NbisSbvFNJLfb
3b1+9VLvt8+w3sJ+7Kt/QAZTo2Inj+wXuvYqfoZWpsTOXNn4yDhbk/EZ6O3g
FL5xnwSwYX5zHacszvAImkSE5mDCXXE+rspO8a2+CfFewS6xki1HY0cjEB2o
Nrs+pnyOeQ38g8qnkoPEa/xV2ylRSDhjB4Ou8Vka8siPZTf4UjNcPdqlE9Cx
mtDpNArsgNGlkpsSSdEP54JN5Dtkha+Z73F64S92v8I6uYTKCMvXPp2BK3Lv
RQaExY5dXV9nzQsBKdZiz7uoomNnrhD1V5kGyh7/tfIQW5nA/vGyW7sumo0e
TwGshcA9YmsnQ1yl9uUOeydvWb4szC1owC9VWux1ZVUIok12A7wSOAtcoffn
I5RxExUMLlwwc1r9FO4FneLimQmZKq/dZ5bRaPL+hlLx0MKeyYB+uhpo+rnI
66wdy4mxr/gbHzbNX3k0OpuzV2MqB04hP7Pov/JNTb2HdUnedHpqyoe9so9f
gU9xlZ4FEzmkve+eV5o2Ce4YxmtQdXJcCsh8v7bh2YHX9fk/ESckWgkOsIcv
1sg75FcouUFGiSM7JkpcxyNLkjnvfbjJKJD6zdwzp+uEmQrcJrmEvj3uzn9o
KbAfZwufwLTV1aBstkKol1LwvpHkpftBVlUvrFD2w+JIsp+ZY4RoE4KWcoWf
dSailctJNFVIeuXtHbDxdMV2v+CHU7DtUdnYTN5yKS9pfiwvhPIzDwDeB1N2
vKkf21OeXBB1n7eGDrOHQ0uY2a6zhXhLvaspQk+1l2BSgforGAMVvmznBOly
GsjGZU5idveWjRgwkTgcqNpJX3yV3jncgWGH5QHCejqqP+9sXoGRHqEORdjz
vroABEW1l0a3FMfhDwiNFPjHFtwv3lJYXSo+AWGrNOJ5+wl2rCE0oaz57Eb6
eUQpIp2O3178tznsjN/oTGxC/O7CDGqGp/RvG3mmWksSj9LREar1iMxCx9+G
1QENi7nWzDW3YiG7gDzdbDSyIgEOWWvEWKLCUnJD/lmsJwphgmjJO7YHkUJj
ttnu2DNaKn+H8gVOcKMf8fCc24WSoJXsZkH7xzU3RK3iUZqyI9bi+Gfk60xy
yozagXsS6UA50IFImtdKW/lTDTsVt4L9lmK9EvlzC5gz0yqayfrcPJnE0oIC
8Ggyvfg4UjC2JG2PB/TAwTTjf01psqwRuRCRfvfXrgvDuShZW6QpegTOrLmo
T0hTlH6mXeUiPBEdfY8ZQwNiZxuyRbMn0NoPyXd1BD6QQ2nwFJXOWEmBL0/y
3hxaoWV1lstmOYLSv07jlX3P38n5ad9WdCY+Uh0FhGKKx2huReD/F7ZvI2Tv
rcbKyO6GDFmwplib15uWyI5xgRiQQrwtvEVi5CAplJlPCdTtVBLtgZ5oufS/
RztenOxobmbdrs/94kqwNilMeU+OLwg9BCGjOr+xdSDlzbQwiAqrMnr8jM0V
pB1RKdtNL/VVvJat59PQRwfJB7Yv+WGjbJBNOGYRj+vD02xJD1saJ8g9/ol7
NAg4ykg3mv9/lE7mpawMj6iXr2+USsMC3NhTexVsyYP9gCWnGQJqVDLuV76U
UR7bYk1Hqt7BUzP2p4Lgehamb/evoPQhYsQVDLz/tiYwen0rcPZbTpNEz5Iv
5ZNV8ooTWUzYtjd+4GayMscYDaqhhOT3uDu8R1tpCPTfPfDmhShYUoNH62ce
SJb0BkUio1ZDDrGXCLOCpUid7G6lc+msS6y/rFYJ60L57f14neBldqOW0uMh
vU0UMPXoXRSygIuzXJWWDWYi+oY/hdckmNf4I03v/cOfRJlpsWdP2Tz1nva9
/TJI0aC1fDgF3lxF0dFjnN90z1wQeAKZehkVEtL2RTM00hWPd09CsZD1UXyg
EhPpanVtD+vUk5aJi8iqkF9ngKNpvy0LyeHip5ZSYpDLkaxIwP3cGAlPCOZv
AHBPShCI7qV/z9jZpUnQpsfmzeVhHkyVFmbX7eu/sdKIilTJD5OZI3e1WWvE
WYbLRisBPa37ZYZpHcNagHUE70iWtlg1pUf9/YjY+Jig9oL05+wHyWKaAgez
3ZwbTkngDXHfKpfUTDrE4/ILhSpw6LDRXhOvNw76pjRoPmwFk1QmZXgwBLoJ
06hKnYFLojawdEObGhRLSdsRBLNarFqCc+dQpmiytdQJH5tFWbaQhwc4Yj1x
JIvubPFb+WNPm3y2F+kieMkL5ZQk0L5fXppyTqeVNuftFlI7ulVt8LeLGEco
jBdeZnI7Q4tOACB9QDN6I6TtkvRS7X2hkfvVxHJBypJOHzZzp5kmU9fHgYe7
3c1YRCVcU1Cy5DxLEHc7SYIADzcCvwlQNgSd41ouxX9aVsgvMcEipLTiGI85
hoqyiF/SQzekcrKzAOTTWgXNIJfbzBp9mTycoXQtPrryOKOIeWCLr86zqZDn
yP5AqFsTD8lQ5I364x0WuIJ1CQTVrYePyHrlGAaahj6Aytt/dyg12miKCmWE
hpQs9d1wRYj8zsKhvd/I/ABVfPTpkp4d+1PiA9Zvaper/cvBqhupGfZPCbB/
/aGvobHFwt4v6d7wQDy42v+TaAYHLjhWlLz/aJBjyq/1TH1B4XnEtzK8PbNC
/0rko5S8KcZl3nX54D9SnMk8ZwE8iPW2VGHcIrhJrXKwEw77bf479H8uHhsr
43dpu3oGWui9Xusdgz9dJ59+ZxalLzd5topIHT9nItDIgCm2P1b7iKOKpkUy
okfZ42veKXTGTTRVse9dIeqX/WalH4FPHnNr9iZI/zwl6VLivWEGNaQ06/KL
ht71op/Pc2AzhTK+hAQkSklDGRftkqrirt305J/THO8ReL0idEZkmQOvbe0c
y1aDOrCQA+P5GHYLFzooK3QjjqWnogizOhbjS2uKVGHUk91uX5IoXigGNWmU
rszdwnGvyOD2YA68hgfjiaxLPR4e1S18hEArhFPYlubjm8SdahNkwlqcHxx6
Eaal5mA30kQEBY7niTBo3f13Bvl6+YV3/pl6psuLRh1TLLfye5D9ZAW2Cn0Z
LG2gOLWiaGLHGHaDI5vqTmoedNgRZPQWEhhIKz5z2dW4UoHV9tRuidWI8IAw
oKNGj1XjIWYCuNJy46Lkq417UtQRNVxXJE4nsba8Z917w9MAfBEtZnrav3S0
eqLpQHSyh5tJX6paJsguKz2DJr/s/cp0fzBbKxmXKpIHk1ZB8KopD0tZ5/Cl
jT4dqlWM6TR76BZwbn++7YzEqf+V7u/DVg+/Dd6MrsURxInEKsIMofU5PhOz
hrNp/yNpu6R0joSSQVds+8O3DrZpUhiLJyMgxIsRIhPDYAXSciAj/ZIsYBwQ
JnKXQZBVdhraFwA/PAhjSNq9iNNCX4ttsc2BOLiz6elkB2r/HIhvkgIkrnx6
kHWr0YCQnjy6PSLPcmBD2PhsYakJYrfIx8c284+NjqW8MEKkB7lwdIPkGbcp
YxgPXDhDIPbY3sIRQavtRD191/V+Cisx11IaLfNF58riGllR+lN5GI1AFndN
sFkFQ8acuHfdqMVlrDiTUbatMz3/nm7sr8a7YLgo4iOln9QX5qTAjBpkoglm
NKAZZwe70AXyCK3ewaPcdNx/YzBWIqm7u3ruQLXHs70OI+evF2oaV/lSK3pO
jb2V2ZcP7sZEtNzsTTm5iGvTg3vSkhvob3xritDhVRZ07PwrZFW64+5L7t+3
P2w3zMCxzs223EUw06rmwj7NioAIRCZhNB2XNDeXuSH+9zPKMQHGjRAlmjii
QN0wITwgTTYrYyoHCK7YyWM9nNrXEpEqX5/H4MWkTASO1hrj3X96o0N6VZpb
4crEbGjV2EoiwSNhLEwpY686N9+XS0gsXmU6kbcf9+BwL9B3JSIYbUbOSWSS
uR2eKh/OB+WOl2G29+kIJIraj81F8MN6dre2w0mLsHBp9G71xvVSnrbPW0oI
/mRzL1JszAG/GmfPOFhHSerLCjipCMuM8DGRafALfpcfzFYEswwVJXmJ4gwu
CzZISLj5s605bOYtazHWp5h2k4iAkvIVtQScfak0opauk+FUxBlMi1x8BHyN
8ey7rVKGm9SzSh/NRNRUndu1zemp86RaKZuPP6FidE4SP+67Aeg98/jPMPfb
OFZz3I8DL7EoVR1NUMw477uFx+0aldPOW1+YEeJFaxrEcPFP85OpldtRQP2l
YRIgJkR6SExygU0OkJ2flJ2VBAfjEVIgGJ5cqCWvQNTRA4XDzmTaVfHj/P8m
TrGH7MLVccXrpuoiuQ1GBcxmoKeObiXnLY65jc79DqR9ONMjFek6rjWjN4Yx
wA2zA448LQIASFMeOaaKSr6nqX+rtGRdvbNvDwlKj1L7CGMfa/nfrHItzgLX
uc+uDg5kv7+2AU89Wc6rfnPe2Ij0V1vdqxubc1NMQmc+wSk0W7TIReY+ohlX
FvWN380jvs46FJEgc1u/XOUjPJxJccIUUDARIdc6O/R2zvQHQcRKwGPg16NW
t+UgE5I6lnlRibQqGgpgF7H0BTaphAyxQrkV85F8KuMCMNdK1ZVbKNRv/8wi
EQSZdxrMMsoCyCKtXRVqbm5PfcDRUG/YarrjWncx1oH5Gnf4jfvVUEUCswTw
endFBW8c4xDewr8D7mECvd6pnU32L83XRvMUHKxL9Q1ZD9H9uU72qyiOXbWs
UWKZdkjIcUii9aMpgkLyCq5Wv3ak35JKyOR+RZQ8fzW1cVMCVxNf9zVULvRq
x0jkJeje2XJtgyI+ej9aQ2Uf8guA9RbYhYI57P3d2ATB8kmV8DooezmfbLmT
rwxS0spmBkDuW47Qui3lpZTwvXVUh8dtZUGpOxX7dRbs64bWKnjvMCmurmAu
sdn4XvsBuxp/+DhkB/hvpY+kWpGGihGi2L7KzEbd2X+e/wKQ/PQHvYeMMRCB
QG2lqh6gyAxmYV/gTvLJTb9PcVS6pxjPA9KNNC/f0zE3Ky5MgXJ0FD9eQaHq
QONivfm409W0yGMXPUVobjMGgm/Du5AeIRZCe86CE5pJOVl/bc1gV7HtoAJL
R3sNRMzeumnDnEqUWkMqpD0930mqpBThRBE1iHUywzMgC7b29piQFsKqOOZ+
xQLCFvnQGWsWqbAjqOlKomS35RyVJdJTBYzbdViwVUosMkmuiL+5Nl4+6CSQ
ggG6La6lsr6mu64ckyorF1LNurOHe8HzfFAgHExo8/JZcPCkeSSi0D4i1Njs
9yXEQFGfL/1aw+R7L29JWhpqiVO31jyCrASeiPLce67KeHOEInUb8cqlWwvi
KWdTzGtIMtTCQKlCNPqdo+ByzFSOE4gygSiKPDkoYzUQrzwcrjhBlO8ptHB4
cRhNR5tqM8VwmknfSktZxODAmA+YJMzg7e6gU6xTTJivHEfExf58CD5oPu/8
aWzKZMkNHcBZsJPRV0LZbTCAZjB9KCumrWpfgIl/uIzBub2hpdbZjnrC/tzF
MXEXpphuVQkC2WkzWgg4s0PdWHJBMhkmVt1OT3TT83sfmk4G3wZkLfDnRWLr
EcnfKqqy9LfwLcV2lqyzQLHvy2vo/rqI6qWIcdSEcZcexMkbw5lxpIKnhiBX
x1XdxaytxenoFR1yZKRahQgiQ61rqniDu7XPblOPvzNKC28gNpaQSWsP1Ash
p73kdA2UdkT9C1WN4QOObddjfIN1p9skoCupqHIseo0NbjFPUC+mV/Ll/Pgb
ThqOCSdBPH4JwPmNViQJYe8xIKpNMBaHjFMlc/ymmG21lQR0RwCJt6E5tLRR
TzLZ+qa4TqK/dp0gDHZfryKcXbYaTUPpKY+5D1HRZPyPniXBQsozp8GQ6QmK
S3PcYxobR9pDms91AN9/EIG7vFJWe3Aa2g4XD3Vc2AHmsICMPrjWLN+e1Sfv
VBu+wj/DxLd4e8q4BlW35kOBK7rnk2pA+kAKYLvPfDIACzNAzypm9SJpExqW
ijbUnqy9JV1kWbrKedobgSIU67lR40U6AeCkkiOQq03ufzZnPQGafv7bmlC3
3kTrb+EBJp+e/eMQMV/4h2cgoQchHrNSIfYSIfBUgP/V6pkGY/1p/jB6cwdr
ftdYENGOEwvwpdPjejm0uqfJ1nCGVXsRjwSCZhBwTrHofaYHWZvFBG6+/o1l
Hs67v2k1qxDDbV49dAPg+VzU5k71F5zrWE4k2G4BhF86U8sXqWEy5rdxf/sg
gSoOqyRU8jrax2Gk4XdavY8xAMXGNEpcNdcqL2JkGWGOaDmwfz5JEUJ0k/nd
znlAnkKSm92Tu/X626a1RDoPbYIINkGw3z9WnH1qmlUtn5OGFbkGFNetQRHS
SMl5OI7nDa+tzr+cUTGFphTlDb+sVJeLpN6CVmaEsTXkz4O7GkjfMxmtzE+W
cCevM2dHxwr/6r03z8E+de6X2HBWPRg5RNDBMQLSsJUemphvL5G/qtR8dvSo
OcHuc6HvXMZI5X7WUZH+YCAc8fz5CoVZG8c/zdhPEaFFWW8MByofUDmS4htf
b4GQhUSkZGnf8Lvmo8TC6tAP39MmG/TonOdnRrsFM18+L1uxQ6HEXKPXC8Vp
wNxVOQ32CRyL2F1PauwjAU9pBls422FGM08uyUZ+9bO9W0bWpuV9w317Lj7G
Vl6rgNKHf2HCpu0i3hq7pTaXpOKGzBnc9GoecV2X7MKUbZNDPxi11kG8PxJ6
Ut/e5pScSj4OeQwws7ODphAvLdUbRBbE8eJeRJLfOJn+7/gexA4DpayoZOkM
7aO8mKW+wuAqTwHdx0iPOXDT3hc9AoG+upI6dRbh4Pqx1MDVASx4nl7ejDiW
WBE94eUc00WD0eGjdmky05qaZUqogJMMYxJZjiS2KPvAAxqL3DkvhaaN/iPn
7JsG8pZoOx+xkUq2JGOYPcK9oyKiCc44NA0L76YY4s7+eykuLSDv5E97wuyG
JUGwFG/1XZBsFELgiDkFkZ+3MwNc6NAK4H2HvwXcGioIMJ3ugiiMIHN2Xc4l
+4soZLGtaqtth8NvnLC6UQ9Y2Uc/vrHeVOKgd6TASSS8STY3nEsR13l4vZPY
lLMjOCJAdPyZpQqIkqzG2GgBYR104XOkOHQiKykbUHGZyo5FlOgXFLpq7bVz
zccTF8bZP/GLhQbJEDii9vesHbqgk+X1eq+x9383+VHP2rpMzcGvBFW7+1BL
16Ll29nuhr0/dm+NBnYrz0DoyHRKRHrIHEGK/WOEgRLFPasItw29e1wnLuam
B0pY7RRMMVlVB4K1g+obTAKEK54C4YekCYWYnXPNIrVkzjREqu+MGvOrJfv8
NpLELHmyRasvt7YC2f08+DTivB4fFa0EIJLm9HoAu9EnjkYNExiEcakZRfFj
G5RnVeYw78mwR0PgVT9MMZxht8Nx3b9rKdj6i/is1WMBhiItydCP382YxoLX
V/XF8Dj03yOmoqnT19pfyv53yMdmdF1/JsJHE64sTBK1lVk0NvcvgLZeOsnD
D82qNX/zNDNk1SItjPD69jbqJGHl+uFqrqON0Rqz1T2TEB6EJoFPLOksgMXM
CGHLLXi+CTxxonMyailfhMUTpbGU3u0hu6VBPu1cS85e7UswgVSkRqVB/pCp
XSXxkB20qymX8f+YCUHMjbe4QrHctMOtYV7/oSlFIoTubaldVPSCgsM7c8oO
J2T3fS7BBdvJzZGmi5CKg5vvs/E6cL0bCiUqTMibVB/J1HpzaIxGz+UQIB9w
kHJFtU7FRQRNIKn4UyDqGkQ42Qim89OYZnLTNfG0IRYYD6B7lhEXoWIIWV4Q
Q+G2PIoOfJkkk6VyGBkx+OR4mV4Onthj0W5EuUUGcSLLFKFpxt+kKTS7p3Wh
wPBFl50pECUqzKg1USg2LfFYu3PaQg//dvS1Z7L835Ygg8vwUmRP0UwZbamh
0YM7zOR1/uUt5+gqmM4rrVniL88GDTuwurU2ozGlsk8Az/kRcj6uIN09wNHq
CMn4EVrz/PagXa0iocIZAcUzR1aXEDfp8s4JC3+N5mIXDzzhzZVUou3XFfFC
HwACBIGgJjH80e8FfKpcD3ocomeZoFO6ym7wtPkzV7We9MNi6zS+VrR9zYmG
t8uCnV5yaJMuM8L0/O5saws1iE2ro6o6GTeuIs1UUOnKAn9XsjUJiafSDG9y
3k93Ae8pG6VbR7GgnMp/HfjNFOkRf5h438aspyJZFuYRzNhs+lrBa07nOFTq
olTvgiUCRIMSY26L/qoI/nUj1j7mb1c2Somjz5fMQ8evyv2Dl5qC8+O8fo4R
+kkI56LotQDM8HqBxTNIZDYMdbt37/gWMrfjBgAg+62W2bGHRdHBQ8YPdYjB
iUAZPRsAqw21zLKWQ7fSF3FM9rf5wxgDF4R7zcgmCtcs5BrNOO1itLTRc9HN
Xm4yfry6nQnNOMmL1a0XQB9ZXz1FHVcD4gsSccHTe8pYFCHABBKqJ6oSddCx
1kDLW/HwK0XbgiDd56M2IHWP85HGOW/kGr92PAKRdUe/MkJEpeqtg3bafKvt
/EJRa8yiwd1qxOPF/DtNo5Nq6+TkQA/Mi4vgmNRHqMt1x0hLV2z/hgfa6+jm
Aoj9pJ1F2j0HdXV4UnvuiJzlTPWP/NmkUxDLtdpOztE4+h1aa9J//nYUYKQ/
PshMU7MLN3pp5D6sMtPVJM9/M89DSTr3hitsd3EnSTlfezwavisKh2PO0zYl
HsBJsFR0zCgMWI8Y0qLlkJt/Ybmcda4uY4j22dg6/z9qxyCHhHw2jWJk+/9T
NMgl5/CkEoX8U8tzJC+6fqUp+P/YE15XlnijAgNHpqtxZ5sOoX02Qq0P3c5+
s/Aa9dQtLcmRl1joJjr4m9gH9l9npkn61/fpz8KvEdl6nkhZtWacYoDcM0lD
ReZwjR7qSbzoDBl4UqwLcQE27Mf4YQlwVhp5eOegLqzXf5q9fLfsAT4uHmvT
gHCiPtoNc/C+psw+p2o2qtLBh85tAKrsURyw6uSwrhdg9XsrsUdJoO0KK9fg
rnFvQqQ+MGlZM5fJy/bWn1NDzFQCa7jX4dESIrwbeWIJdGn7zng1TZBHwdrQ
6AXQDzaNItX18HVhdIMKUPqAUoJr2ShYaM1+aUhrU3KEWZgPd2BsZyJunLYu
Q5eICKeCvUwWiEmmECqWfZjAyJixyvAnQ9RwhCYP3Na3WrRRbl4WHz9HnD7t
t6MQ5GRQudEYZH0z9BZmqwVgBxlvxIZXZTqsmtUtqqRzULyjv+DxxetILLjk
dAg2CiV79MkJFP95z/G93HZi2MNj2RyGP2wdhGeK0askHqfVVHT1kD04raRg
tMyKrv8tI7XUk3l+3cdeX4ujnga4FcSLczRNuWrbTN/FVvhPK2RCPvxHsLSe
3sSCZ0Y0XjgF4fQEwzAxp89MqxG2EMr8aYhELt1K/XANJF8aVt5zAFvt8gid
VPGRzIam55uAHS4wNGNmjYOKnerdmgUhliJ5gU+48Efv1ZLZcw6A79L/fMEn
/VkFjEX1/AzziXkC+B7r5xhgJe6wSVNGiUSSXG9T/SagmuXLp73c4suuFoSt
xtFECL7S0GeolU5rzRn8hZ7tGfi8Ctcenz6KuMF4o6Te4A3qHDvy08IXlSUk
RvhZxuaPcY2eevYbVDzj9OW9/MmR2ggrS7O1fbp/yiabtgnQBwTPesq/f/L2
Xm2LVyuRyRV8RWaOwzxVYRZ8ORxXRqll93z09VmyAkvL7oP1Q2yu//Ak0MUv
ZYmyhBnX7OwfFU+e3tFoK1HXiNa38XPKpHGuX3Bwq0Ez8f0hS/b7TdRQYQ7k
aMQQUzXfgVe5DrWfAsUvRC3hBs5jUqRl7LNEEhoT/sKqPq8ms48FQKAnxLGy
gfs3zwLJQrl8mdJHnGYWNfuJFTQ5XCOkh8u9BrZO5CEfVSZ7p7XwvK5jas2I
e0CVfr3njO8d0/Bb6SGBWFbsHAl0B79XjrLyr1WgPLtZwLw7SWtcRXC3Y2Bg
O5KprevjMgvMthyIi1Iu4KaC59kMkmhOAatl+DCmFGjkmhF6yWLM9TdL9DRx
TdsJEXyc7yLmNXwGFSuL2lV/WS5Z3Lsgtw4R8e+GvWOXRu/XLDu5OF1CXC8l
0gIahUKko1sFAdvLjzIm04HGLj4O7KRXx5PmFUGu5rJfNqzCwRszmBmxvVhb
YByZoArccMhRFMf1Pu1AxpF8eqyABuHHNmZAWiUidxwQAGwZsE5L88c2fGn1
7BM/B9irjqkCVokRCOJ2o9K+JwzgYXcp5tOaZ8r9GUAwHu1e8JygBePRs5XG
Sy4ggMMawcK6qFc57JJQVOPS3QVXNj9JwXtfHgavZR0wwiBCcfHv1VXe3lyC
qFnzSrH5cWAtuVKqzEyvz97BmEcBAwuHhV/VykO3r+y8AF3i0PDe6K3z+IfZ
fnThqcjM3Rf5yDLgtLS0NniZKSvfmKv+2KaOBLH41Ta+FpjWfCnAO970Ge+O
UAaDwxJ9wmcxDg26kQ4uEWFUcfz5BUMFy0TWjQ8pO8+nAkfDAJQD406ybw84
rUcC/OYwTyl7VEZY2BA9jBV1Wvvy1DvheiRyLKgI0/t+PdxJHOUGh/DrAcGD
qzpLlfr4IkN6CpEcaR2dFSlMuX9GS6CIeA4HX7U1xbJGngLUyLo2h2lMQ7TL
35y0km17FEERoaloSxs0xTfiatAl6P7PnmO4LPQ4gtAUSv5KjV15NTFG65LD
zuUVx3/noWfGZDCQQtmgGy9Vx2SHcomix7X+oJyL3IKpVBLjAtGqxmKz2WHr
O6m6RFWNu22ft1yYFNzj1o6OwLwbuPlVKLojeX9e392OBjdLRiitMa6XOG6O
/Za+LJr+7pPtFRwH6RZWUHdQD2fAIF2G4ck9C4F+eoGK6onRiPB1673JFUvH
r0bCmXWa8kK3JRp4OW2LguzZ5JcZYiH7q856j3MR56o4h2+ecFr23u3FHK7u
QFukbK8TJamEQtBK4XMmyBOUM0D/jixcM4VThkwrtqR+7JwKpH9dQgXEccak
ennbD2D0zpsbj9BrDRm4NpfWw7cgD62Y0Oig/N07KlAgB8aK4HzwY5esWHwr
xPTXR/lxJ6lwwmICjk2YplF5CQ42rv6IhWxtMH/R5gDYScawYpTzwac7MOcq
PcRj/2039qbUO9yGgy7WwN4ijQBj+NXt1HOxqdDk8njVpAC5KQXh/fI8yzn4
CPnalIvmQcml39bIvR/0iCPu6AK47/MjyJHqHx4u36vVOiyI7r9MeV6DOP3n
uBBbbZcL6u+NwraibHfRpR3DZK197yWxLjLUx/MMgT0KqHBreuHv4pXgeken
bMnusSxkwXfv2VESw1qe58dcZMQm9aQwDn46ICkZtqhluLKM+OtqyrxfRqxV
zvSfwO6SYQG07vLo4SyvaQ2nxymvGPTtIiJfsOS/ocwWMepXdy7xoSxSmJbT
z4Kko1Z/QWKDDZm1/0r8N7BG0oXqIIpRjFEcYh0YW4F0PWRzkbeWC3zAWY7W
PISzjJp6xlx8o/1MNUzFO4QoHFZ7zfmE5ORPaq+yODwIF/bVDgOeQeZ4AOn7
zAIAKecnihB9o9CtbhwXXnGFWvupnj9uQyYt1DPuIc7sfPbED+9AkLQgAfON
xQaJ6cboxvtoUwTjM4+Zudv07LcGExBGKFAFV9vKs6IomzNsoDgO363KCsBf
+GpkUUnuSPHbmCCUsItInqTnP1Ptmqg+iLuCTK5Tz2drOhQYn1JBoFYferO6
JsNRZsU2TylBUGhWavRargDtIlNVASLX58b6t2+FdBJnGtIFYlD2NgS05Cjk
hM8ygTgAOz+6tMAipQ9rat0R5V2SuKWWvp0ukrUu+BGAE1IBDRb9yswCQoC+
fEdSjHuGBYoj50q7NvvFmI/VCHmrMw75Qhw26amKoJJfhQZZxLcy0LHNYfzC
Dt1asK2Trnbo1JJKyJ2MYYjMoaBkiBzcQ7A0knpf5b1wP7RTOZqQnn46Hvgp
c9EmCV1ycMnBMOUcEJal1/1jgVU2x8UM9juBdsIGXWk5KrT7qLYXweiM4NWg
xUcVioLntdcHN9WFoJZ6wRc1PeucZ8iWXJsX5TT2VhZsZ50CI9w2KCX/5rHA
QI/K2q3bR0NgrGDK1Y7C/nLGlyDqQ4kmVXFCGuphQuQpYW52M34HA1cAVIrh
XU6jbsyyp+E2eQzwC9mQEnwe75FkSfRbDmQkCXER4GGrdQIfD2mkmylG/wVu
TY9Bxxj63k/w6LzKV3i54/JuV/vKVbNenfKGndlmF4YzAaP1bkI7LaNw8OIB
d+LmtyPdww67vKAQDMDLttNLJQk5cViFo8kr5FPqhUSk33jUpluy4E2lpdTu
5aizyz+r8Soe0AIBdQU6UvqG8msWfcinWnio2viPRPb6e85udyEhUryAshQp
CAVxs9R+1VEZ/96+eC2ehcLPBJKASqsD0PxFy5xNe8RCaYPSLqfsP7ZvWUjs
guMMbCglTr0gxLZ6aDHQv74mxD4bxwNYWLcB3/6ahXJHlvZJ1LJxQM2qet40
PmQNSHz5Mn/HAHo0x2zMR1ZCbgcul3tpVOCKTgnqlyo4YZ75tFrP7jXRvK2J
XnNXlCNI9xeRmoCOCi9RDK/o1XQRmAAD8vLFHl0g8pbYnRQkt7kecaqplpkF
S2fYsyA4MC5QuwAq6QBScfWPUDPlChZbtLWc/a13CoHEBxt0JIDQf933Uhmc
76qpENWqTNgOI58pYVhFP3hmT5DQabD8aNPnM1wqfa6TzAEBOwwHqxKAYuf2
+Xcg/zGyeSOAKtQH9fWCqOjrYRFnxIDUa2zka+6iFPlJLxEqYUwBq83ntXOF
l2hiVPUOlWO0OSoWCH0jj9UJ07WCnoLYZu1xFm+YZKBgebPt4aPtVLFbK4Ch
bxR3HWKBsWVaxLugPGj5/6gwAflX67/EgKLiY2JIiPO4MeufEsBIKaq2y1X9
HO009YOsh0pxjAY8FPIvDAZr1vkRPqOPkoCJn6ncIbtqfWn3irbhH1oAL7nh
0hK4iP7DCDtvMUAYOPZE4i5xAr69r5CBPLtLnAq+9XLHHYqwWw8bNSCzrzXT
JDc8+2ySXIZNVJsTcIhxutiC5JuGsvstRMy+2AiT39gFHBAwv8p3yfs0+eo8
mJLpeJDmHTsyYo3p7u/kElhg+h7aoJ2rtMeg8BM67UXfOMw+Q/904kGNgjCv
iQlWx5s3/QrQewlAb2TiAgHrNCPF7XTeQX/ln20i7eHvrfz5UP9AMsV+3o2E
08URYyI7H202bzapzV01kwvOt+hSeYLe5ObxSarzN894rY8izs+VCMEt6xcY
py9QzkPzrj4RHH7892w3BBQBwrD+vajunaLctmL0cJUNY2Y7UMQyaUKXoQat
UaZwXf6jo/cIVZzAkTJ0KPhFIWccm6vA7LZehnEZtXIhQhp/ZEdyBTIGS1u1
DIpeMtFsGD4AHJsFbgqlFM4gBAqKMPLRCBnVpRP7bc0tIDseMBlYccG0g0y9
Nw3f5Fl5Ad08t7Um0G21zLgecOB2MnpuVYrQicDQznDodLx0MA6ibHK2TOCJ
y0qJM5i6RNruDW6pPZrW4ieNSJudX9xB8TL+qKfFvfSwQyuaT2swmY2G/dhP
pl3Q/1h/J7hYtgwWlYMJYsVO7NvXylOnDIyLvAniXid2rXCF37KETfqNYHVp
S/f3EREVTM0TLuGKW/W+u705ttKR/yi36wzuI/k3unYIAQMwF+9SyqKPnlsw
GCWxY0A8njQnzaf6ch8WsQQDgtPYtS2Y+GTfaN5piVC4QWwjXXduMqBL+D6k
7E2+7WXAj/KIQs/3saTTrpAPEy4yPEZaTKy0NzXfWO7TIWdMn7iHIKkRK5aH
qcutZxX7hdbGIiLAXcVLj3hvDCdWi9GqfR/grajeqeCR6cKEUVUjmQqBCmB4
BwfZlGXHGGwkKbwkCsVwjfN2UPsB/YIuttkPjk2i3yZnHcBkcrcOzCwZXgB1
rxIbABAR06GoZk55GECf8naMuW3Cojl8O/jl309f+psdIq27LSryRTfmm1FF
3R+xzfTBfx3WtfpLu98Np6bgY86kHpqlunq/0MiQLCykug904ejKmY2cRRWM
IZ9OEkyF/INl+caOFrrwCtn6qqowCNR0dlx+pHPospDuj76mDaS4asgHIG9K
j7+90wDiNCV3BaDHMAZ4W1jGei5tiFIl5nHDvAuKxbOuaCa7fyd21h7lAqJ9
AAkEH9Yx+gfWB68Xlhpn8JwiVGs84GbBi5hSrfW41C3VZCYh7Eky1UUVXhia
zSV/P/Lt0kJg11u9ejsj1+O6CeGjexx7XA2qNuuAy3sMONWIB6eqDCYG/Veh
P09PIlAB8Z1/NpLFxwcbdKvEXx33eBxdf2gNMzHgNfyemMpQHIhcDGLp14hF
E1aLcZ7TYu7+dG57WD+WZRxfJURWhgr9+gOSRl1lrYRYERxzrz/Nrr2AuDgr
pjkO5MsEA8dxOn8DISoFG+xTbxt1Cu49fZ5wWVV/2xYGsh+I+DJNkjDiHPqN
VbLtvpn4A/Xm7gWNrZWnG5Ro+B3XHtvENaPNqpjZKcevVGKbEDX/8WW3Q61J
aEcgmbAGpUtqfao2Kl3GxchdRm/eaVz6X8+vxkORNBEdG3nyciEXAu7LmVSK
wjLE1am/ouQZmqPx2iWmt3Xhbk1BamWXiXVZCljiOJtxEXUJNCfgKjcV0Abg
7AUJRDlv7Rh/IxKKRhuXE450o/hGoOvAKBf7/XqauV43zUYbwP8BU5j0j1ga
Bhm26IezG5Vv7hYc25UjadtQUtxHJOcZFg5qriktdN+RX16ASjxzm0W4jZQE
Y60a77CNNI3BLzi7hl1K9/cheYOrLdMibwyRBsjZmaak3MFtVuslUs496PXs
6qRGuybvy+M6641MXBkWPN3TrqRzTYpJDelCyRFEXWFYwgMXLMrmSph/LYkX
QFYXPP+TtanI0u7iIWmIMPhrRXV0gXDT7M2zenl7zfPY4zlJGrPJjBSXv3or
sjDio04NkXM48NDIOLawLXrXJcXkvLUVzNLTSfDJL5Aql7ksV7JIDxfQpQp0
8omol8J4t64RAPBdGIjqk4hSeSD1Rx92c3hqYkqsTFtACjLw8Zuj8MwM4296
NLaYCODXHI4Qtc//yV5gCOwy5T2/OqjcZdguxinoH9fB39f45qItEDn1vCtt
qViMxinJb7NkodTj3yymVJtf991uIcfRtTqtqFlZijksmlxAQ8jBw+IHSmra
XYub+De3JXm0fYaSGTBfW0kX4clp06KZLqzV3fU/5sZuYXsR7ZKPcUyB6TMo
3OsCmGPf3uKWJF1UU4SpMzc002E5sY69BGvlXczD9AqJwi2p3hxR5/z0v54m
C1vdfRoba9NBoXKx0zSMmvkOHdgDTGTxbc52N1W6X8ySShkFTk5dHdsxrxqN
ff7m3z0tDFrMUQOOf5zSPVYwWjq/3RsKxD1b3YuoFfjchZ8yNdzBVlSOOG5A
QZGMzIMxMpMZ6Zux3m1o0vAKQ517yjbftpb4cTlQRXSWHS8WwDfy+Kavg6YD
vucMOe0O/8/hBKDAMBNoPdfCA4MGy0cDFC2+rFKnZgPIwRoxKN1vBAHCVpz/
OgSQ81/iZb5TDGA+mDxVPf9Angcm7iyL7WB41lVCRYpCw76XKb1sx5oTgMAR
QoIXYS6Fjd/aArQNhDZaVN4+8ksNP+U2vCnO2/iHGjUcNvy6gqdkxEPCEJuG
Vtnfb0YVNqxjsTnA6AJkMVxiHNPqcS5v7r3hGcuedU74ZaMG1+6eaYSYxHnL
LP+Z7XmUgWPQx50VUUgjE7AzyiLwrHJwRQke+Ja4XOrxExOVM6Bzv6l7n5KZ
vAmMWp2Qvs2JUmUKWddz+IXpEYzWJK2RoII51BsC3ay2c2kGy/9rd6xkk1rt
9zHil9MZlKIEWXWs3vpv1x53NUBv35AXcoQifVW/iMUGroz8oUHGlRkMx068
1LRebeoWcNsbHA8WsGX6B5F8h9djsZPGVXtB/pvos0HcXeNJ6L2ut2JWPMsF
3V+xM0BrpD9wLbtTQLiRTYfPcnOIT3T+OKcQ86+oqitj8sy5be79WA+mh5tN
JKWwV6CR+bDLUxjyZieRSMd+JsPgi8NyZDWUGCZUX+6FSy+Oaos7hBI6i6IE
P7ouVY0Yy7XcuppsJWJkgNT0gRtkny9owU5OZ1HXQbLH8Lf8+3A/geTKJqny
mC71Gzbb0LIjUE9IGfxfPXJ11ieT4mQSXgl+ng6lnF7l4G+FMOBVu9tI5fNg
QxHU7wuFjWyV62DVUW9W5gxQGuxbyVkvJ+88Xx/5ks04TdYOWB26ZnG7xCOL
VjaNzVc2kRHNczir6yu5Xrse4X4IKf1ncbxElAYQfRh2AyGkUoShpo+tl0G3
pGC2BqAipsFNEelOLLaC9SF9xqn5sacAZvKHo1jRY9TaMaNPudqDXSlz8+Ne
avZNaV6CRXcSgAB5fR8HrMOIHpguUiaU/HLlNcsvU2gKvfnUOmmZ7xNeDaaF
O9qo5DUjOgp7NUqwWsrbDv+7TYmC5/YZZbpdoAZ8ykn0lrygwkdUVoG9OBPE
rkvQXE8ava9iW2uEWFfI/R41X1BQ1jqDmWF9u8utuTWkRZP9lYsxmsmtnf9T
Oh1sKkmK7LLNhmZJL4/B2BPcven51UEmwUTJmiuIEcET+jZ4pp7BKt8p3Ruq
vXIKVeWEVY4UJpG2pkwJcvzSpINhWy8TGurna2xk59NArXcgFqbKS2QAnUk5
r21kpH2FiG/zVi1Qe7s5pa3LXKvXUz6AgpROFZiW0vkJU1Smi/OGG1Bb/QV2
6tmCJNWsbpKcO4wEE4MbRBLy+qSPH+j+9NRL++HWbvUYebSuuDeydQ3+M3bM
xbb+QuUKewqCpXKgMtZFdkc57fNbRSHK6e1f2PjzUb3tzSdt8fn5pC+xsxcU
wdnuKE7PSDxcylfxQwULkzERrhfDpLKJe/vdnrIOXQvAk4JALzx309RMeJQU
RVpHDXxY5Bjc1K2AxuB6kfCvtnpa2ZIJtk4N5slk3GuYjJ8RlzZ/TK6u8wCe
HebcITw/+pkzyxZo7dqNVMwqMcqNaWGkgouELUg7VvtyU9su8mFTOVMSzOpY
lEammR6O91NPR5nrY2gbfzTKI/fru/lWv4gwJfwq7LQJZkRzXbkp/OkkEfQH
q2jEJVa+8XCHLauq36WBDDgUGEKH3Z5tpkLErAd1LECGLRZcD1UqPTbs+0MK
q+MJLA37m0CwC+deRwydYh6d3z9pyyXX9J6wEnmA7Z+MHx9ecFy35rqzoEtD
vVbL/IZuYRt9rFy9eX/NScV/pYwnddvgWNgrm9+4MiuuN1xy4LNglgpadSZz
4c3yyuVpstcQUjuLZhmOSzp4MRMIo9eZN0tBUxILUK9bUbU9WtoD+/7EeBVW
8w3276GDUuBXYo7kbuzpJUYsFBSKM8BwRIW5/rVb14FNGS3NbYRdk6zeWoGo
je6wUM48uXZQeTP87bqvJDjfi/ZdO4nPRb9L6q4GCImz9KT1iaNtV/1JDL1s
joBNOexH49G0aJiYd2/qmhUB28pindwFilXmIINu7Gy5NF7K/08F3XTQ2UqE
txe3Up1nZ369+pPbhHiIs3qCRoi/0U/rZrXzGdgbLEb/28lOZB1P4Ws/bl7B
AABLvIepe4wLDRQVWfW+7eKHFqE4ukGHijOWetcb5V0orgnkF0lAbgc2hXYs
Orom5zjJIflf9NXiIyyaCbuXXN2RP+tZKvUWFCCQ4Gk0UrlLtuTIWv00w6FB
hB34V2pE5GY3wiWBPKBHiMnx23FAcVbiOhv5dhE4rjdTeqOQgv4ZJreeUBO7
F9oAIQEuAOCp4k3xqOFcQrNiQRROSKdItmyLUb+0+wyjnPWkVjwL9tdCtZ2S
Ja/WiRjyeZLHXEJp388wn0jCB04Tmfa9HBeDoFxy4PhVc0QVQvQki7sfV6g7
FsbYuaZdgmcA/J3Dfp/17iOE9BH6ShlHvzlndZ7L8knKlDP3k981AtlPHUws
eCDSvD1NOIRrqGoPXJpawhPB5zeqc5oIUktUV3nczvav1wbiFEU0ETM6hfz9
rgxd7dsJDRohS8L8arGIv6n+LEKIL1dZKNJG1xVDk0TIGeYqC3nsH4k0hc4f
FuiFYcEKle1seJUDDHbPVECg1sWuK7a3x+PsCg6p6I1yd+VeaAGH048h4EmY
uV9YOuJZX9zfVoC89qpBU7nxOajdNyarM97EdD2wBRb/jZxo8E1zkzUMCiUQ
DI8CICGIb7cBWMNr4my7JH2mIvj3De9LKDppfTayChm0bAjpi/3W2ApajFN6
5KG/F3VQnm5wDRpZZf8g+CR/v967Kf63RUO+0JUsCN/xMg5TgD/9BgoURW/5
gzxW7bKHOWYCP6oty6hv6YKeBGrjR20R/XPnTFmkbkf6IeQ9tMMpuEkWU9h2
9l9KDazRGVJC0Inv6fjGZl4Ir47DIhiELPrgEt8aAi+1LEU8UZ5/QNEyIEgg
cdrckQmksn+18Oh4q9Ol+6UhuH3WB/TqK6GfodUHoDJA4tdnw9WRPnv/mEv9
K8d4QpOtKx0/1TuVYhUTRSBTLRXmXUIpx6t5v7/DwW/nh2crF7OD6giRlRJA
ZzR9iWDngDfztAQ933S1ILLv8n4/oBwEs+YjTledSVs3KxCYwjbMtERALdqR
/HWdrWvhBfrZmmPYxQchN+F5c9+cKBAFC3kQ0iMkcdLScNYTGBR8ZBM2dOlS
V2To+yg4sj0rrQ393XzUkxmEP6cESOhKG/H5CHyizDcWjhu4GrpURGisGVBb
75leIoZGEBk+lIrFw+4ZWRNfVYBh+0vQG5VX7Li8iQ/966ya3VIRMbx/Lo1w
3SAJmkeyNBM6wgwjqAVfOkPbTuQ9lXYyJ19yVJU8SrIql+dGoCYL/odz5YUF
SppBbUDEsz91JasOS+BvBEfA8qo2n1RVWCwgxkCKsT+3SJ75GHMOPhwTttaf
rKqcr0FxF9keK/xS201pqtecnHNJI8nk12K4973xBhzxEYx7YQpQv25dlhVY
ahPhhYmhjjMGzWeigHA0fjEg8KHP/7ipSxAc2meTITMYsJuUzQAm8542yZq6
13cWCf039ghALKSPqm+jL6OX3jXteckblZj2Wp00jN77F6jPNzByEf9nQB38
wmw73xWn6/hP8NjxEjKdxZYCXvx+6urfeo0xdctZvY35txTQU5CIC3iBMo80
PKex0My0QKd8CAj5j0CTWf8RljnEg7iDRVuX3hVvsl4MOepE/PMqy86qVARD
st4KOS/ev5aex/wg2ZMmtyWuC7Q1QatZ3LRqA4A4R463dphl92iHd6EKJ77P
afrvrTBn/PANy/OAR4gkUtrXvw0P7qa0GwgJew8dgF2FiEs38KlFLqFvlNqV
/X2Nqfm33P8gDfWeGL9eCmMNjrkRvp3m3gEDklM71Zq/wSKZKSzkJCARXNGv
joUPzlSA1aMJxsKtRkAHyl5FhPQr7V3cg9viTx+yneiADvA2x/N0eOn7m53B
YzgWzGi0om43QW0/73eaClNEClvVmJrCcOwnDCvy03UC8JdWX3VghKSwl8JG
G13E0Xef+lPS3/OV1hmdp4GAInroYQW8EvhsE3fLjo2/E4g9dr+ZSQjKn7vm
QJwiuxt6w+a/cFXHvqlevsq2pktbXV+BE23DBnBwGKzJ0C7WiheaU1lR3K3d
Nh+pmS21Ce6G6Cu543luRMIns71UTSx1Ns9kRKddXRUnKkvja2mC7lnWKdoD
RSqPZ4EM0bUTIh2XcKLQiNTjcYl1BzvyQxxhtQoN5TYHH1Hj+k3UCnjabdb5
41k+/l6QPLIcNhNIV6Xsvgf3kU0KikHcRn/N32U3KGMzjpv9wtREWQVDjqiW
jiRrct52ejuccfSQmpjxGzXXXQ3oEBaBNoVawqBuLWCXJFnwNVB2E9QQZKVG
fgz7L748eG5hj7yFYdTG1tp5zy8MYNQqOGA/z27MjVMqTEb0zbUSCFcuzLIM
XOv8yfWvPDwjO8fVzKfJsAgvb759hF0Z0WhCPWYaFLBAxTfFGGzw2NZlKC2h
7otl8rzfpwh7zITPxHorPuyR8HOwCntMLB13nXSqzuT3KATy7oQd42fS3+le
E/ssYNOH2vH/UR01E3eRFQ6UDPXM6aI7s+wCMH2ut6iR7z4muwEs6yxVqv6C
6HZCa8tH28Ui3IURfr+Dg6AwJnKE4WY0WbY3F2LpLg2x9gciO/fHYM4fU3yK
p1IdzXap1PlhmXYEN0+ab+PYgmz+v2OeGWlhxOQM5C8c9Pyc21CxvCHBHZXS
n2RZ+U8sHUDUksjeUltMW53/gNLgPyj1lhnM8aZJzINDBZgkSNxZ+wYH086t
f+cV8YGCMOWKHlT/r/rcV4UM5X3ffwkcB0sXw6jd0DDFWj5nljzUPM7VLw7d
vTaBfzbCr/zJ6kx4a941C+r4kHFXkR5J+vOnsMEJzGf7WleFQiaYR5E+IUgb
5FjuiKOOZ6BxpF5+FW3IaUgfmvIfR5rVkkiPsQT1Q4dWlxSI+VM2lOA+8Vxq
tgnDlQFJo1zIYboVAHXYA4RvBJ+mIkiEsYbfwJTlLvwBMPEbz1LaKV/+1mFJ
ssgnnnePa34rX3nZaapCCI0vxW/U9lj6potZjLHuTKhjPcfsCh1nQ30DLhy7
At9aRfjp/I1X4hSBIoM0gl5QgBnkGgdiPI7wQO4MyWe/Pie+mus32iP3jqUN
g7kF6rgrm9DDcllyang2aDj/METKfANt7rBD8wF/QbztH2cNDxK5jep2kWcX
eYfFH+0SXZYQU1n0t+NwF36YJW86xUGT9uzrx1j+rzqxIOZJriu6K1OP5iCD
0fvoeSgaaQbigi+gMIoZbVkMMBT+2b5KReIj9+aPu+41EIVlB5DruS6kwVKx
xarmehIyrfojNqomQNQ6RjuQjinV1lPvVctU1uDMH/bT0UIdJOhGj/wUPgFX
Uu2P95bjiaQoLeo2mJBTv27LIL6JjA2aYS7Ni5tvWRzEKzf3q/vG2Mlpr6mZ
ahtGKfYZLRN4vR+3mUNPk1o6UlUBwbs1qubQF3T9ju9Jzh7mqN1CON6PldKo
CpP1Jgg2Sy389wYaBnSr++UwvQQolMMn7RuH3anw5MI92IsFlvrpFKlSQzp8
iSvJTsbJrmshUUGvn24MBrtHr1E/CjYlb1c5CD36lXTUUSH1hhul3rS8EvjI
o65UIfoCiXAUqvfchnHooAhrjhI93WOrZy+jK59jcKrMNX5+t6FWHZ4/uech
PcUNh5IQtp3g1LX1N0aQB78cYMJLF3ODL7hMXfqwt7MDf4fgPH7lUj5dMcRD
t3XfB29dk9+EjsCvmBd50EvvQ5lANgNtMvK22kjOefTQ8G70mZjg0b1A8rWT
Ilq7LL8NatMSKYCsdSGYiWGdALMyf4AB6dRiHF6Fhm8w9TTV9U3a6PmS6pXm
R/HR/NIYL3+FPlG9qUxrhcKrCCmSsyr1ctmOpfqcEWMgCsJlklmDnXw3OWAE
C+dsW8eCvqFBtpsXVjeQVZ0B59U2581mtvoV9yknYR7gOiuVgpn4UeVbr+ps
32Ya7OkvDj/mu7g1uHrF0CiRbq9m4mhwAJx0FxiqOO8Ry1TdFK3+kn7vk2e6
nl95tJKYMX6e4nFDyAe2hBGMghYaSbBdNMi7igkX1VJNTxRojzfhnEDhcU3t
QWiL09YZzz1vscN6rDWEX49IFFeSq2UON4PjDkkBz7JB0cZfAoE25ltgbOfO
33NLKC+bUR9aUP8w03WLTXZmXDRGAqx5eTtv5FP8NyUGaMlarwi7TyB9sTBU
79ywMKtnE/hgh9nNxt1k7HPcDBvT6/hIG30Da3SSO7lGfKn/K6vZbUoHV/Qd
H8wxRtpXDshkpTZjtYDCz3NRjX5jLY0CqOjV62RCKq8Kff2vIPD1E6fbQpMu
X5Uwil3fu5n2/ilLNfOeA72SgYf3nem8TW3yjJNZ8B3mgG5kKvEgx4uAugqf
WYRCfJSxg7jLGBRuHMI7MxudgVD5nuvzUusVhjMHIiPvTfYzQYNInIn63uX5
zLxOwj3yDmrxSG8e2FU5nYEBNmkqQQ4eWtm/1JHj3KiT/YcSwkflQ0RWcl6l
K3EorihzOC6kYXf3JSg7iZ5/IyTS4ATxMFE6NqmDlOa+UV38hsGJON3c2a7L
UjROL8Ymy5Po8vC9/cOFAbZaFZJrsd2IXmqbS+A1xOnIXAzclTxYYtfGYI5s
W34+SqoapiCKA1GOreZRl57eMz3SD6338sC4ZbsB8Ey0aMcOXpSlwG99QNuQ
1UrLwM11I7JNyB2EgVjJPad4eE5hzsxCBSfEn1MIxnjfyu8WGeZ9IRAVmlFy
tPFDn4O71Fii9htcAz5rAD3H1tL+f6Mzjg3Lm8BcEhhaf4rzBTC0pGA+pvAc
4UlhKnH15faKEteap1gKPTOkVVLcrDQRVTkGrYMgCrGftJ8WlEQJ39dN3BCc
RE5S6D/e6JqmUcVlBIrZQ2sPO2MINKYjmZKHjoZ+P+994Heka5+U4q3RBqEq
xtOE7sVgPnIsvTxJU3P3jFJ3SwR1nqV7Eqfa46F0jYpmhN2XB0EM9S9jJbrJ
bHEgK2XBNg+Y0G6WvQMw+v9surEwoUkrkYgTK67EinKNCgBeAdgjUv1b2UYm
/yifTpPI8ayIU42bGjTJ72OGNjwhbWc4Fqhv98QE9AapZA9qOQgQds9cYWgn
KLusEXYkz+uZz51Jnjedf9BdCl7M2lmwfRkjQytGJW+1//2aTOChcAxP8s50
J4KoMEXcpxlrjGFZSs+DuUDhOMB45uDcAeuKcFY4u1Y0B2WOrKRGv/TkCKNW
VjnOxd0R5nGWLluk8I7g2jB2p1rxbRPgrmEKK6VTT1WgtBZw4bbc41XEr/kN
n2CWCIMiq6/wJS5tN66ydrd2sqMxEkJKfGNBQsvYszyTPa2XLPP2JQ1kE3yn
CvPPNGES8UFaEnjXilYIpWMhUMC6U1717z0cuRAs1OirRUresk30SLV4zOUs
uKuSdytKUMcOlvi4fplSjNMUy4u/9fB1Eu09Z761uqiYS051W18LLIvEtdDv
TdqzQiDr+43odhNRdpF7zJxaEfdZb6TCF52b1rJvbg1/0rYRjkyxHv2IvsjQ
wUEQ8lBBdzSg+tED27LhAtLaJmIFmZmbvFMw/6Y7rJJ+Sgg2fQJhdK4VjsZU
CKhApp3Sq+DUbiQQwKzJFV1ZP22zrrmcs5gm1M+iHKiMYUl/dJjyLcbI/gcv
sTM+NGBPgh42vdhXyEmQp/ahLZGhmgySW6za6aSsUgBqtcl6ZvbRFCaetn1E
9FwQjLtzE01vMoZ4/HuKP6iNUW660lXkbFmh9UkyiAb3Ap+GPwfs6ookJBIQ
xOO/nJ+JQ62tCVHD9hUrGUv5hWfiFK/aTRmjl3yvXwc/E/o49xMxDAgQywg7
D/aWn2kbSUHnh39EC/s0o8L95dgFby7SibO675XVzwKtL3Qduf/sXccFTaD1
2/zOVxjD7gSjlPZ4T13TRYAcFkA6HWCosz4U3nVZoZeJOOSL4hOkXTVNugdv
OyOMzloSqSl5993qH1hQOVmape7LLh9/2FV4wRK2wEkcjmP5IEUy7w7qsx5O
tlAxEZf3jGFYMs9FoDheI7d8bvR4s2u0z9UttJ040vb+FMKnaFdpK+rAAy4e
6Q7gWnJn9A4xsAZhxYXOCjWOKNxfq1d1egJViAcy2c4yc7dnamrALa0iilCk
cYBtyhn/w6177ONGHl14ZidwMzIcQY6fyPJ5+4RNONkv8PV4ZPCT4I571nNt
XnKh0pDvYMVobmsthSdl/MNXPw2aiWJ/qTNkUh+7Zy7SOkAFDWUXlGZa8Ky4
8xHdmO2uQ00KDXpAwthDbk8WfY9ODeuAMqXDgVnOXocNK7oa+nU0rqbhJ+jn
s+B6TdQfMDFR/EDrQ5WM5EsCwyhl5rHFZnMkZv2iPEcInWefw1OSxLH5Pvsu
RfE+Zol45li3l5wB+/KWLG055qAmE1ImcOtGjQ/UAZp30BTQpI+l7K73czli
92IewF+AjwrAIWGQb3jOI/cJSk+WTU6APeW3q0sLhe44UOH1YS1x1N0h7NnJ
pqjwEMSlcyFptJmaKX72w8kfvNAYUD3BPPyYxhRMYtFiGg/FHZHTI2RxjsYB
5+XaOOZi0Poz1WWa4/sSrwyfkTntmD/0mN50gWPObdHBnP1bxIf6MY7j2TCa
FxOufx6fZaynvezQ7OldLSzR5czonFiH7YGBvHFcP9Eoe3FujE1LNFBK5UFR
ImWPp8C1dFEfKx86ytj6dfAXKEOQvQXUKUb6nv6GLQ4Eh81hrQISdfZW+2dE
GHqHLKF2E0c9mNSIBznWUeoGvtKmtnthf0bT5ahlQ+mVdj/JfBfTQss1CCxy
1jRT7zh2K1jzGASTulEZcmLr7/hOeK6urRI2NBqwgK9O1MPRZzCw/1wSvEHv
vxvR/WnrQaNNSDr4caXuM2GwMhu3xgGFPwFNAjBDH2KnAweYyn+9pZcvjYp0
rTneupvjbXT+yRmpGx+w00rnJ+kEoAsfDgmJz7vO16o4FKiS3xI5dGNMalwT
P+wZgCr4YLkZNK3+Dg+tYbQKaxxl38wfQP3v5zL55U0ciyuWJLFynCRn7Qvb
hOEw3AyNPyPztLqjfPrL49lPx6SxAnU3WXjYNhg/P/mdg00npy6MOadfhQY5
uxaNmwgfijWncHBdD+JvdRMA+4JJ+gTzckUb6VVffJQPCO0X2daSLVSV3CvR
JDh/aTFTDJhtC0CoKO5gw4peQ0ctuQYMK6mofOOnzMIY5YCG+l7qfHMhxS+X
waw98O0PFW4PrSAjxQvazkRzcXoF22KaFySRlfEsngN4HbPEncSOglkdy26D
Rihzv6VnIzS0XSq9Zc9KjzIGhzdW/gtEJVQtMUEkfH1H5b5SK16XfTRktyYy
ahEH4n9U+bNio179m3VgtU/lyOOD/IjyBIjsUdsa4Diy/w/8xIEoeMdn7ocC
NqQ5xsXh8TLBuSior9pbhNBxeZ9vfQzIddHF8CiJTsX0RpFNsQtcxTWyyxiP
w6kz8s/4FW0e98QdFzGqRWFyMd5ojt+pD/FGxLn+QiY+oH6m3lXd77j491Qw
RT6aS6A1PgvrS+T9RigLvAlJzxnlkpPPejtn/qlEFPfMLTdlIkkCSLRF4ddV
LJuiqWmneELWoJFAWZW+tSSTW9HJ465TnnkdPCi8Ast1jeMyL7mg68Cfl7Wa
oFV8qR8t9g8dNvKP2q/CVgT+wEdssGv95L3WTyW5GpBZIImlIOZnki5a+wqk
pqdFJ0rYYxyGn6d4+XbKpeWV8Z+x2pehdIPV5XJu4V9a5v5JmpJD4u8IXoIb
pymcHW45noQI9S+em7hjDoOaRGJPqLQWrOaqzTGbThlfwcDHeiW0/SkE17YF
dLd2jlJSnao4lc/wS4ZGaTcqWvK9JrDgFIszWnHdwGFSDEc1ec6sW6oP1iW9
3flZQ20F87PJM8eFKcrLntcn3+XlrQewX6WQ/ER9RmUcXqmxAzm2a8j8Rhvl
m3vkatrucXcSklIzsIxfA/mifije92LRKGqqzr38PuHGjYG5dQBsp4q9IvUc
Yepx0iiv9hVVrnT2iQH41WIfdEBE2iJhV+L3jD9zIutv3/bpUd3vBomCRdb9
4LgHZwP89xeE+suMVWrEn25lWHg0B1bZok9wReJ/Y4DxSPC9lrRoidj8C8P2
8e+1kS1tSbDnx7rHad+6rlnqCAQzPASpkn0Y8CEtUiUFSRK3ZIad+bXaLs64
XvKbvuREgzh8NUzXyL31CaIM2R0/pqljsSBLXm2gCSoUa7QHZ8bJJBqnlCyM
3NQfpcE3raVYCPTAiBjCxTODvF30Gqek8wyC2oVwvLq3AHZE16vqvE694J6U
e1R9v+xObDvDMxAzOcVVWoU43/TeiOvA9JbRtC0jIl44aniPMKYy7DMzwzK2
LXab5JTsh6l905JYmgWZoy/mxLwhhW0fZltg5hMcJDsU3Sp8Pz/oS86l6Xpu
8sWomwkgdYQHpQiUMHRpQNLJ+v30qJXX7XUx6B2s1ouh/Bw2g/yoA8gjOFWe
q7RHIErtDBRdQ8v/oanSkHzrIYo8rPeyEU90l4rCuLBXd5uzrsuwZPaKpj1j
8E/pb8z7My8+yhvwagkunOnsix3M8Nl5oJh6ie590oNFzFQVWfIjlsRlh3Be
ZmMyNhQcER+sr27q7s5r24BHsOkm8/KapCl+wp6PT/yG33zVsVz47dRYQDt7
S+sGnLzEKp+CTB88YXPJlaQA55tlnk4i0EfQrGSqZ4BFJgB4T65WUak4bCZt
i5BUvrpc/cqxvmaiY56SbTIOvWtnmKg+KbmTzP1f/39ljyC2kPebb7nxHsIv
U7/4D+SHENqCevCVJhzIRYGXGOuSGo+6q4oXuy+qT/fIFMvbWGChocIR7bM1
FsP4BQuklBwfKJJi5EXhcpyk3uoZ8/SMg3r5zzln1XxRDdKxAPqdT9APAZ1x
IBs4UdmVTC5A0U+/4fn/QWE+FbD8PKyl419Tl96ZWftOOCupIGWp8TpOd9zA
6Rk4HifpHogyu58dVNyZG2uJUIG2xvL9yNlDhwVQ8G4a6nEbis/XdTxHacz9
ocFMTv+r7sR3g23KlI/gXKigPgtbruVk7kBzsMdvGFBZPbp7GjxvWuDNN+8U
yrwetb3zklc0jGjac2SQKyqr4RVfZXkatjIE7WxTlh2+8g5XACrHZAhZimoC
KUErKUlD+V3L4hpXgNrX267o8FUKYAsL4sF1B/r/f89q4ffzZeXA9lgkBrFa
mxkstz1vZEdgeZFD5DzFjRax5z608UKGLSNUHC6bOWID997aSfuL50+5veH7
YSQlonmrb4l07IgLX0mLL7qZCBnTspQYkZbPIeUoKzx6cjYTYHh4zXAIhnSJ
rDZOAsQuvTIsDBfnfzTq1gu+W+jg8JQGKF/DXnrStlxw1ugmmGjU7fLULenY
5OrMBkCIcUh+RdYEostIqCwZ6gSVGEJ3eEdOF3zOp5P7aT6KoFh5dS3P2Inl
hj4TJepT+xRhQITFFZfvAqYISRLKIRgkAJ5IkRNxc3epl9OM3uwZDK04w+O4
0mv7ds4dC0FWoiaXbGMsOSz7E/E0xeheekBnO8OXpqKTrE0vXlAk2AiPYmWK
eMi67B2OG00NUeEaozCPaEqcBach4HrppmGS1/6yEmObIdy1g8f2z1czbho5
e0PlDxvIVJTsCEJ7GnnvPtOHox3WJKScM09TyHQjSVq8+rL0Jc5ce4LQvWoj
yUY1Pla7s3tkODyBwiyRZQTy4ZMqlR6sa7uw90pGpql0A8DB4CdWWtgEPJGv
0NdWzd3Rp+otjyoGh2JmmgB0uGM2jwuqeX7rfYcVw3rbNcWPSMva0bRk/PLY
Pwwsh8g7f0DrnS7rThYdlYWE0AF0KV0Mb6KfV/Qdi9emE1oeDreuFPxvv6Am
j0sRykA7Duc4QLyvZaBAX7sdXpKyE2Txe6StuBpUn8rPf1dR9lFWxEhINTFD
2kUdacbs/K3xbSfR4MBBgPIP0o1XHdm+CskVRZIST3GXA23QKpCI5Tk4VMYJ
f92MgTRRsGuNH8zQTX3VfSNErrNPc7LZ7B9pQUHgJWGJ9fHIVdSMcB5BP6a8
jTxD1vPMDePuo7DvO3P+JHPdK7p1u+nQqUX75JAdtFQ18n7Ncgtcpj0jseF6
GNUr8NwUvB9K2e+kKzQTyE1xAkNNGwlxV8CA37Y2TAMS5NbfpoR8vtqSj5eR
UuqAajNaERO0qxA7M7E6xw2Do1XPtyFo1nMZLKigw8Ha7K9Wb0jBf42AcM5l
DJH+b27wqdZi4WkO+0wamjAcgFpD9k2uwHlNGnXpHFWQOVSvneByzxlkUAAP
tjzRIXlndZGxT9boJXSZSu5tDKsqIvG6sMpgzGZnNYfXf1mYQBGSe9NCZDsf
cR0sH4Car0ePQNAcTycOSd4//+D9RcHdQOuO/40uBYsd8a2qUCllpsOgYVaJ
v4LJU1Lw9PQVRz+m4ilymIPhGSNNZLWgdrcDOp1sWyFKHk3ZrhMqHgfWf+Jy
8OJUwFkp63HTuJU/fQ/Dry0VkKjmSqBIj4sy9w4uSoMjpcuTGLuzdBEcWC8M
CqGP5Ico6rsMnCvzYfXzTaffXEtHsNOQY+TqwLlOdur/nooK42hG7M2A2pJe
woSerCZJOfz4rhNUIt/nXNXzQGuizhv2Qp0P+Ej7vltHq5jJTSa+Ap37efzz
/J/MCfD6skhWcNLy0XFdkHuzAatDzKLwyUbb6ej4/knFkEKJkzWJw1AxYypJ
GwaSfcxOG5ieJhYaWmqfYuj9/S5FF4LzUkteHSayTCu/Lj7ltUHmr6y3rtBl
kD/U4xM9+SZU8S3WA5YVUKMmDUqmR9Ha5MWSrx9MGBmG1zmxlLJCJNnJorpL
whJkvHP9ADS5josurL8LE2Lt4a1WjaM8dtm1k8hr9bQKDQH/leWHjsxoh2n/
KKnocVR+bZF444z6Lb/2cIz52WPtafoRqfkp+Uj5zApoQlSobDxh7me3H3Zr
kiGK/H9gwZXy/FvqgilJ+Fkc+cy9PtaLy9RqhRy/YMrCr2h7yVN6DDDS2DXF
usU/BEfkM6LYaCrfEZfMwnDnN5PzJStJG7+CnTSmDLNGH6PQG3FpZoCvFaBt
aTz/XSyWS6ZMWRxTn/DOMWJ+S/IZYTqSFkjAyUhb0/Xg+QKamXFs1VMon3Nm
m6cGj/L+jZwqqiKMbJUJUGawGAcPmLSO3eQKmjagHITd0GPJLY2YlcUikcUI
9dq5Vkng72m6gqCRyo9BNpCMwhx5jmanUdooLhKLhc27e3CAPKH90ORUZl6p
vXVBIqhVkJN8Fnw0toB9oMzY/5XbKHcJcz0kXv4OiUmvG8p4fwysZ18Ts8Zh
adXZPBKk+sC/VvzSWINO7KCzRdcWXIm/qjmMyMPP8pzHhnYqVu5IjePPNs6f
jiiGyJ5c4UhM+ahE+aC2AaXp5f4lcJivoVWzH8GpQL+o9wpvYPNlRs+mCM+s
3nEzVgpRiK/R8Nv5nPI544tou0A8tBwF51yY/Ep5qr6/8e9cPqn4r1cF2Mcx
lUc385h8Nt2VWbn8tyrVavPLsnvbNXKpts8I/2Tgg2XjUfA3ZZ3iPDiP/jPZ
J65GFO+u9Wo+rlHdRAf33vFw5jVqg7eUx+xOxymlNIVm0DlIldLWrKvncAv5
2a/40s3B1Y2gM86GT6qwxJgMYQUuf26tml/hYGFLlm65zlbqRZ3MR4IqJdom
hblcxjqMfos57mS3C5ln9go/eFQk7HQ6DDpMObSVMdpBvYntkvg1KMlvmNNI
cR/b+3p0EgMZ3AmuoUBjoXsdV9MiYJpG27GKxKui4wr88eBXqI3UWW+cUXzR
3oLsgF2cEwjJZYrde8t6vXFFcYdbxZ9nNYft+Ow1Rig5NMYXcDRPT0GS7eRA
zEI9Cz19hTrlY05IZ3RrhIihBcXJE+pdpag2NT8QPW4CujRh42dR5qNR/qrZ
aOdveNL6/SWTeIzZSxrY5UV+ckncCdc6pNu29SW+loQAgacTL9sPdssOwo0V
WzBHK3BRrwERhTmhraijFljBvXX8tUy3vJic7jCrayGFR5Qy7Puy2a8j+7np
8uu5gq3uVMk9gIiSO9ik2BEfDezfIwaPT+MBiOqI+Uz2BVg7YeucRlvkbZ6c
rMoDZtTLieSRGt1syDyF7hmb5Rl2bRf+qhCRl1jacZbL3KIJhtvtJpgQTXCL
cJGADHK/YCqH3yvak0Ik3Yu0XVu/a7dvgZgam50q9rJMlV8Mp6UCPrsk0Kit
g8c/mJ4Wq4xLqCOlJpMbUQEaP0gX7R0XnQI1tdYAebppen9fqk6tVyW60Gtb
nzUKwk3OlPIKWu9zE6E2gCZY5NuwaUQJxi4KiaS2PYKTjJODgF9t2WgBbHcP
E7MTVFuRGWMAflyHo3PUNAIRq52U2NTqCrOdtiJ/hCNX//GOo5g2Fey6WO8H
WVIjLM/ISYrYv9vQ3hYAZd7OrsLiogYU/AIZnrnspLBRICbj+gdg+Vc7SdW3
cLhIUcwW7TGoHI34Qx+jMJkFVjghJOhbu9eHOAIZM5N/+k6QqzMBkpoLHkgX
9ALlp4y/AwZAZVwSN11vsuW3sra26NchjyJsrsw1SHtqXa8GtZ2eiLdpKK/U
rVknkEp20w4yW3nptWAOVrdCSeegtKkNDRsybDcDL3Owu8PCVnZt5zTNpYe+
O+Q/wCb6kkiLy2sw2N4a1RlbSzbBw0BcbVD3sdS8+NYsi7+oQiamgDKMIRmx
4shrV5ClXakD4RJWUQnU2Uq4XCBB5iRtxNSWoEjFZaL9X+swm+CTfZHiZjox
mmwYw5N0S7t8oLbunEhIbWWamVUuIYExZgGuUphot+KAQAJFfULR5VMhnva3
IY4+mmOijA+xOdR1r+wY4ljtElEztZSGmB/hTL2dZA23t83Sv6hQc03ek1N7
JMvTGtHXxm0rumBDCMlrH5EncsjrkpRl6xdgojsYO2IKUnpt9P8KizIoL3Ty
fbNm0pKTwzJjZTLR1rLuGJ/GnyUSJr/D5xxQPpg2Z6lw7QoKh1SvDXsNm5vS
0xOS8k5UNvZvQFtHKQ1720kSvZOde60/kfiKXaJnshL0tWhgPX1O25tJK2ys
GKfoSNvwRsjR5VbHxMigETUQITYcuVRbK8OVYP7hfPM3Leyfo+JIR5g4yILX
+BAqtCE9Npzb1vJt5kYOT7Iwe1EoxLXqgltE70aNycEbaXu3nMhZJc8evFdk
DmJwr24dtMVeDr3jEwkweu9Vx1dZ4KH3T3D+mPKrtPWY63nQWT18TZK5QQhH
4AupphNkpN/6HVrjaozz4vzGGUJQnaZHFLARF2FViQz7oQy/Ba9qyAA0ypCy
xbIZ7GSjCRN/d3K4JiZo7EH7caxQYqMgxoPuvn7KcpZJBgXuAPyUAHckqKux
zJqQrFhkh7XVCZ3U5tLm8oX+50s5d8dEbiqaZjRJlv+g1fVwqOV3Pgpf9Vbv
EiB8d1K14lcH6+NovFyySAdzPOfN9rZi39jPUEGfplyKtXFJQeoMrF/zqP7L
n52suumJIRcU9aZq7YKxJ50uznDLhBpkxd5TZnXIwMWlN7+/OBYCCvhxORBX
v6cyk2mopPyuQTo3tb2+T/lZDQkyNnEWLNMyzzKJ9VkXt6nR6n1Y8ik+zeH5
OXMP8/N1F+Imoh0F0iMxCYzYiBgJ21hK8IWNJyr7s1HeHih0v4b4Yr2VaOJ6
M3jF0Vf+pQM8MaBNzbF6ng98IJzP2fFQtPgPINP57+lzVC0ELOuX/3frhaIg
62shzAGQjqNvESDocBu8LJZ5wrGaLiSF9Dd+xJXfp4zfVJUN0uhHDM0K41Sh
NHWFnHe4Ga7F0tbais9fAN+3ZR3aybWjeA9U56gZBM19UyhzckubItdheOE+
+X6EhCi3UbcUmLMBVGmIW4jxP8eBZa/yvJaqEnu2v0bbYyA1Nx0UZpdsG541
+JLtsBnvryRwkhkChIi6R9pc1eAQbpk0gzuSpU8y6TbapeztKuurXIEX69Ol
vU2KrHZkIG+jnOnczhCVMJj1ZZTerrZ9GgnPCnpX+hcdeKp/EBZQ32ydvEDm
e1fjB+MQ2zUJ4oP7FQi6GWYVuf/dmYJndBGCMH78CV7qHMfm1yBtJ2D7wUKN
WdAaxizaYLJ8UJGwb7aKXgPGsBzCz2hv8JkdNGdMOoSiXF5nWukUIhwhSggt
wAROE00mPJOd3FvW2qZvJq15rEKQ2H0cclWvZvtDa4+nrhuRvG45qEdJvF/k
EpvOapX/QRnuKiCa108Kjh2R2Agnpuj7M7IQECxDkbRni68UDFH79euoV/9x
n9FTnHsSoOO7NVkvjiZ3SLr3CjK8JYEAo6Vc01qJ4MOJVNP2Rh0XEW9T5ruV
0Xh0cITAx+gs36+Lvx/FvCEegWLf1cSTo1J8x0RuHUzR9nffvPec/YqtBauP
A2ewm1SKS2K2u1FLupss84RvhLBynAsKoBRD/CkoHKqbq9qB0/sGWVOvVz07
1y6GvHLF0KByHLsEqIbyqmpzbVBTGAMNMgs72wI80i2kcdkCJJPe/sIIlzIy
UPc/xuBc2WfA35mPb2OGpuXUAmFAbsaZVifkr3AYO/UFSLTjkq5G/LSIezcd
Asd80vbQbXHsqSZHEv/AlZq12HAeO2WWkQzoFe+kelJ9+9P+TdoX56hI7sX3
7medtpfEmHqm3DcGMTyklc68gC4Cb2AcnwwRkFrODrS2sagKCTLKtQBFMBJm
BNBnvlKkHVW40vmxAWw9LMKAhii3ajzxOqQ0hik5dPHZZL7O+UZb2kxA3mmB
2uiqnS0KLnobj1EJwkjyDJNzX2klgvzm+1/kJa3t1ZK7ncIooxKlcqH77nWb
wscysd2Ug4x48beL8Y9TdNeeQAUIQjr2dSAohB9tHgIBg71hFYigbdixwxqP
eFJHsZzj8eroH8R4xJ32DzmkJIBIH4XfQ/LheDVVEbb70IMQXlyFET94okBU
7wLmnwEn3l0HsGDIsCd4NqTsR9pxvPl5b3giUg0WC50c6VE7CI9whPpMRLRj
8uLE51PWr2JyDeUwNPFXnl6RDyB8azc2gO2VNbdVMr4bbhM3Px5BIvL0eEsd
cnjobI2jt52sW4wI865vxC2r2dk4beaYFIu4Sz+mAGjTew1yM6xLmUEYfuPD
o7Mm6bGYy/6uT0SVydmsecY6hz7nxBj4LA1pe9UZ9P6WRbstMRi6LmpUyqQ5
rguKHhk095T4CnsDxeClvb78H3FUX93uym9YuwQ8HABAY2K2nsCo3aJNS6dd
J8zBak5tzHP21LhDgfG+ThEXvbkCGEvXaYDSNqgTZv786g+a28dHa1U/K44W
3btSMaUUDtD47mYAu9Idnky86lvktcD6yq19EQltLwpKCF19ISFL5U0DsFbJ
DFtpoaODCGWzsJZiaKoDBabsKXh08tK3s4FLRtW0SoksJNj6+FzjccH0lRwd
tHpjJxQwpEpxB6LKHC29Tveo9Vwb64EMfXN7j10KgCC2EOw7x+LDJwJnscq4
OKCL9FZc1xYuk9NNCu/EOOEEsXxkULkX4K44anZL+Jylg7NrW/rQqANUTUtk
JJ5mv++/1aS4I6k1+1HK7SAqVWQgnhanpUAO59Q6jz09+iCf4th1xltlpJre
3OgseZ9dhvzwtC+/8PnQMsSXRbKYN1VtqSteslEFYq77s0S9tkT8ADlwYupw
zODmrK6v+3c6SMIv3Z+n5pNOTc3MlUE51+pacGekYio4N3hLefrJwCWjsKTO
BRgkcLtGmD45Xn39K/8TRFwIShAgxeIjCDyKbLhTqVMFUJ/stVhqcjEzsVi0
HprEyXvDpO84L4bpmiHihizGG5364sr5lQ4oO9xcx1YKLyg6tcWMl/YQo95d
WWVeGr+MDpdPL3f3MGUvmq+ljp5x1h1ueeIqSqEeSZslZPdQRH+FyRF/rneV
37yDqQyus7RUKO9SUpUECkEIpJTECFWbf7JVU4g7n08zVldxH9Fn298bSfi6
nLn88Na55tanWWSdHbpRQeMR8CS2b/zgD653HfNY0h/KHsfhN1DpcJNchWHv
RAVsMRvXBrDp02o1zDZIL/b0LRufNagWP0a+jomyqI6C93G2BsJQ+GckM5Qx
9Idu/pCNeQTPuSE0u7Nhsq8GGDAyYbN54zPt+yvEiQRbbteuyOqVq588KmG2
9UHNjcOe1gZra9k7SESm8gvFyn6X2qoRYaCDXRG5vXoHKj5Ckwrunc+mkAij
Yu78Y9sS8ZiW1vq+sCrOLX6GQ/NVqjFdN39sNYRMBz2ct7C010ldC7NRsXdL
4z4DCBlKjGzIzEiZ4i30lHq3w/6wB54AfdvtPmSwP6/oOG6Q8NdVox3ITdWA
s3b14YR3vTizkCSOW6RvOEa/67mgpNoOtYTjY98EON2EUOq1qt/SP+E4nonm
+WVe11RL6G/TubPlaSWL3XH3oujAS29XWjzyGFcv6ledFD2pfjjRlBXZLOug
hA3aEv232uN5u7+u4WvaVP2GRJ5U7YWT9Dm/Xr5Z+iA9XREAzrc671MZs0hn
eqNzBQj9n8cNDmVBrVTUy1E/oikVGWmdpyEhGwrbJqS8Yf1E4VDROMipSvti
cVruIKVqesb7mxdfMFq5s6HAbmXq2s9Bdeexzw3GZ5FhBqx8YfjG9XLE+y1i
ygGQcMolRTUkiKdITKrw4nt25rplj6c0r+zvywVIPZuF49BNZ1nXtN/D392m
03zAeNm8QnFiTlAN2ZcmVQt3hLgylSCGAzaRxjuvYkksDMjUL2cgM3ZxFXBZ
ZNGDvMob5PXJjcetc8VW4lNG2dFuTdse6OP0F/g4cuvqmaWh0VZiqmCNhKOi
7SSJewrWms1ypOth6RQfHpQjKnP+EEUvzG+zsXXU0GeGjPBYKvVnhnCXpeEl
fJ3LxNljSCkB3NyZoY07xXkReFMlx/AF7Jo5kJOLJkUzT1RC7M8m++v2W4GI
63AZOunSF3EZZ9y1TnkpIOxCd3LWz/cY2RJ/QEnI4KrdOKANccLH/tzv4MH/
8NNaD5eD7rDgr2/wXXq8F6RkLSrPG5VmFwPuJY9szxMWrIxpzqIVHnjEplQ6
W1cA+ySS3x8+mM3d/175yOtmfRHHdLjKoIhfpSQG2aL+42PCVtx89T5GvwQ0
pt/AJaxcdLoHcdLwMstM+8xA99GqfQvl3KH6xEvAvCiN+GRw9nvw/GUyvSSY
sZfUCQ9l85jqsN8eAbM/iEI7tqhYGVXIBmv7Vw++14GCAkUgW1LGrjAXGRg9
L0XW0y0fB1Rb+xDOVRoCZaKIPm6ec7vFN2PvVkKbnCxIlB4/fGEVwTkR4Ozy
uxsiaGMp0UrP7Vsc5ucX/9gXcbgPyzd4OBqXmWdGe6RE6lH36Ytp5f/ugFM2
qgB8fVxqZ4ED+EQRyFI/bCNy5Afc92AmvJb6fgDOvTNYEXc8LIbIdA+0Q1F7
dVkqonvXxAxwXEyZSGCyoEhYJIKks3kXkNZ6P3KIBaXF5Nqv+emu88ALO9wy
Oy7u4yXDcKWPyyfvCl2qtNoCr/3pYU0LeA+fvtqvy7q0nGfAOMvX/r/KLF3Y
j92102+V+cQrQyQ+eZ98mNuLxzO3XAOnW9GwNwxGOL4InashHyDgAP7YTjC9
aCU/HQhINNr1qVTEDt9V2DEIYp7ppc49AVWWQAuiRi+/9hILa8w9wnSGYCa1
mY08Q0aISOfUnDvWy1vFzThti8nawBL8fBAT/nm4HvDh94RcbUrh+HIedFAT
I01ct/yO/b/nMMUpEMLRWVs8gyMSISQG/7vnRnADJ9KFdJ9zttal6mDA4MxP
wwu2CpDzC2jFu0BpnA0IcQyskm1uVYP6MLvywiyMgYGq9/Ifx8Rc5/+PC8t7
srjuVhsRGSinGnZSA7J6sWA1y+rM41brnDapC4/gNZKEi1ZaAQeNpuEgg5B8
QLp9O8eSSaZOuccMS1TFpLWQ13VsX1XOnXws5LG8+vocSDGXfzsbJUQfha0J
L2hkjngPGDPWyQvP5ovrAVQs9yMS1FASfP5ZdYPJuBM1HACEt9JJfTwxgUPM
4KpM6PLO+IReC0UZVFTsPHlXgT7uEz7gTEHXrj7iz56tM9RrYcKRy2ZchKFU
xqd3xngMzgKJAzGafIyQNzqEgNubHiDbf2UnhkQFSKKfQ+DdfaPFAdd5YORr
ekGGlweSpJr3cwq19J6yDwEpFPC5kQz2CcGSKs+PAAyd2wzQZvEb1tNmnNeY
McOdVNHzSiGDO5NUyV4vIuRi46ZfWycCsRs4bgr8928cVuy9YfHlTxSB4dKl
gx6RKXqE327Rfl6taAvPUtIjl8eD7jOBvYwNH0miOKz2ukKez6bP6SDxli0j
8508chbvszrJyvK1Fz6Eb693St2JyhE3ajs0W9y3Fjums1z0I5it9r3YlPxt
z2TS1vKxV2eq3V15ZiKzAyAO/VfmFW0AL2N8hjYYtgqcrtUq2Zyim+SMVTvh
sMrnah0cEUJpfRO+e6aBAJl66a8PHU9gkIKYrNDSp/1jBm/HJFQU+JlFe+pv
C4bVbPEnkSrZotVHWHwexcvEmrh40gIKG0xWWDH82lIL86xh6CLXUGzVc1NZ
rU3+Qyip/5RHxMwOUIltLEEWMJCm7tAOqFCq45V4j2p8WE1xCce1Hd8eAmwN
aBXn93T+SsLmFHCnrxzmqpTH4O2E1SDpKtBw6NIeUYZ7XRL82r9lDXmRiD0q
5maQlNiJ+ahhXfWlTTvjhFOg9cHlSD9yyaHPWrAIwUdQXxcmR6LzVKOUDhVI
CY2EyPAIvg+eAEUO7nth75xKsYq4VKmCplxV7nKIBeEQwWUbE79d8dwM5LU+
PtoHVZ+g0nqtEk7FLFku/xgg3rDixgKwQ+ZNJYIo/KEawO7Ion+IanNjPD7h
cmytq946D7f6PtzNxOCx9dW2YFYBbZ8hyLCLkcWYq88ReENpRBCit6lnEuse
zJ6l9fxM4nueAlCRHxjkOLUU8UiWiBewXUhTdFN99/ZLSmzhdWKEf62n0Piy
rHALcAcUOrbzGGDRVHacw4tTRYpJSRiKIbW8agsMFkGIM/OI4EbRIEW5TZzn
+aDECbIjOg8sxSeGa4QbFxuCaz4XZljEzJpMU8RKWim7HHQUo+fZB+4LDffY
OaEs4jQoj9ytgodM3peV/5se2yIYkCXNwpCDPTHj+hv3JMDI3647y2xpYdip
8VsnOBNTNrJD9Ksy9iTmCh5Jsq9brdt7YaPvjn1yniWzORG/VdWyhAv8u7ui
aduygdiuUgmTDtFU2rlNRBNP21a4QdrgyE+HvIsbARpO67M3611qBI/JiZXk
YEaW2vnuWovFJCPkoOPbW7CIKUMCWToitYa4PG0QvdXJnAC2IVkKLgQDOMGt
XzFa8HxYo3CIIITsV1UH6kfizqirsh1M9J0H7CzjZj6zKA1MTzrbHgyGcOkn
hNzrCk3JAkDLzszuTOcUKvQgv28eAdpm2CJ2GDR65NH14R/VjAcDFahpIqdR
QSsOnL70MFpZ1HpjXAUynczXTOcbUxszNpHcyVPgpC2z8Z9eGZzcEL44W4h/
gWYIX5pDv/oMz+I/0C0OoSLOFJDK/wTKpa4+8ijq6hSVwMkPlMi02JDlacOt
ZPRfolt+ZIOyPStfr+onkywqCVf6xE33959Yv1DflK9TMNQX0DuMPb274X26
vlfrL/bN9iTwjOMLLvYI4/Yp8VrapwwIdJVnKHrRnAVEm0KQ3jN2A1JBL8Bo
bckMhRtn5qkuaIumXFdTnYOIFhIJE+uhKnShD0O5xlTU6IE+I2e/gvHjrUBY
D3YntTepjt8NLcnqn/FfbJacNNf0EYEIibm0iat0Ido45dCEtrjJ+IPRu4Po
2NiNYUSW5LWevZkxvmiA2KDrAR/pDbDmWxq/lz0poMXTW55TDZoazqqagXXJ
0xC1DN20+Brt6Cb008zIokwhKxLiWnDJjAV2vVyQYXQutHm3EY4QwQFv2scg
mavgu5BeQC9GyiWZJ9z92i6qdg5UxARuGcXf4RsNxugR1NVu4KVxbhiwDHcF
PSA/wWFyJHO//KbJ3/QFaC/qCPjAhK+rnyt3XWmddFmztC2/OLaL+Trl5g7D
YG8kdu4Qe14F1feI1O3XKXr+9XB7vfY3sAXUMCkRcNRjh8K12qZXpxApVZGx
k1ZInJKDA+tIRwecVm2XMSH/ZQA9dvtw5EEyIs9ANvNMU7W6LhQU85Us/3nx
GY2tbaXYMOoKRls4IffRQyW5muvtl4krWYRg000mqq0bTKGXD9OT2puBpm5d
6c6fKAbchO/5XzCCjB/LFxxfsKe+y+X6/ganxTidHLCTigWD3Duv9QVnDW70
vLxwVCnK9fqHezxcoXY4YB4lhOUEy+q596AkdoxjPlBHDbrSehqn+ipz1n62
ZlMtl2UAu2yFOgwoM/1GgPcmKc4PGdPE9iebSZT8TjbfR7aBi/WmqmVSEQdO
vcDQXtWneJTTOwVrSyesO42NOo7tMolLVU2Xm2yN+C30IwPr6mGCb0bo2L/8
1Vxu77rOcAspchky0ZUJMg1lATrewOJFXFVRdFX4A1movdO9U1FYyV2dMQyR
8jODuSsT0n/UiQ4SyctVJXzE3SG762GQXL4xTLYM++wgrMyF+ESZeIRzF8Nl
POtdJ2IN/SzKZ7lMsl4YpD6v47kd+MZaaT5iCAvSrzrqAUr3AubcLQVO/IOk
8S1DN6P6kDJoQgBTQWanIIs+YluFfaamTMl6PYBrlW5HLXECPtK7iRymc42c
MDoIgH/fWe/So7EEMUXhkoglfC6kqs80sj+nlVIX+fh06Cmwz9x3/0w4x05u
vVf7Jufm1sJWv17X4T8mnzei8QRaM5csnxTfecKR1wXw1t65r76Y6J/spdLO
bJWoSmNe2n8t0U0UE+7gJ+22c5//nUEY4bmvxkvzsxRfk/gsShW4/H6o6yIg
0gjoHkJLuVFRbuZIL074sakYQaI92Q70U9UqJhfDOMRsfiOXMF1mwIYu22hL
JjJ+5yTjtbi2wa35WycLnOO7G3sZ6YNhIGkn2wgP2Amq0xfZbBhkcCrRCksL
+RoI/quq0cxsrNCusMEA7qd1ZnvWjY/y9itNfAmxRR7iLaJQ5YKFWRtmJBhl
dsdVdQk0E0AolBa4u28Y1Sj8RAbn75k+nMOoghYskO7Ev2twwgtbK8HLV93G
a+P4xuRQB4BRp6oZpT0jg/8p8uYm2+Yq8G6FOtLB8nX9vGX1Ai0cy2ue2aRp
T2RsKEGZsz8SUY5z6U9KG7LPLCIEZE6s/4DQFWeh80CpWjZrGcbJoj/m+URq
OB/gvVeS4vAyoqTczvThQF7nHl5H3rddALdUMKcYvezcIlQxwJSH2m7YJTqA
+vQiqE+RiSun5sIgDNs8r4T/c1l0AnfFlDi/s/C2Y/nSS/nhnqivQdk/isGa
OtQtDTZlgHWFFS7DLTQCLZduIufCwcpix0/neeKzl5OGaTZWN7KsaeEkoSRc
N0II4jeR3uRs8LLqWEz7GoRQapzMU5wd29vOUlEanc4T50YR2Iv4Ui07t/q/
lN7JpnmSQmiYj2fTUKaj8XID3Pa5sbOS6qnsrbV1ouvK9/pmYkciXNnEhZrj
wCoRTIBTB4K3390uCC9CxvUGz23o6sypatgKuEGExh6M+VtGRsEPXJnNzviu
v7HQI5TlDTU/ZAOUulNuUSyV9gyhbyyBtdEJxDfMmueQWnCGSlHoyf8wMlkv
4lun4HnaNWsd9N+gGzMOsPLRRHjuiW3aIRI0j+ob/iNJMwtbtvLh8qYjqTP+
K3t7ylIt5FZh46RhqlB+ejgcseVzMzuePgAg1rMoxO3vWRwYIxQ5ihk5TJ7b
AzpdZ70Cui5OxnEpkjQcgrjRktEPQQmHC/yDPOuU1yCFYJxNcBAntQNl0/vl
8vARh8bSPwbmN8qWtfNxm4blnnhBuUexEk0azlaVAaRY0MmYpZMuNx8dVrg2
A5EGpNcoFPidZHNDVyXv84CHKBjxtORdjepIFrpIqutcGXL2vLi37I05KbUv
Hwz4vlEbw1S6RScquTYt7WODauB0fMVtexjnRwbI6FjatcJUhN4OPqG3st9P
hclv++SFnNfFaGYllzzSwXBH87foJHNKbUcdAxXeC09b1d/lh6g+uNV3papJ
Hg8WJ+FxI0nma533y4rmvrOapCLfa/krJtLET2M2JwpiEVH5dtf0rTEpS4A7
0EposwCFcpVuaCfJW5H5oefJhOyTlukuxMQXuiupWiOcLw0jo4reOV7K1Raz
939gZuvOChOTeORVQMqudAGbQYkn01uKAL0xBh3rFWaAsVJo38ViLM7pDPA9
X36rdyQe3JpO63YBCVOQrSnTKla/CdJ8neU5JlYnqw2q10MaX7xL9wqI8Rx+
IBJPsyHvy3zNcH0JL/AjjqE7WKL/lDz+HBTtGPg8dUX9oYFrrnik+ZFrhdoD
iIh5LqYx6ZWEqIC6rnLAQTURqJEkjogzFv9fEtOkfbN3QwpmcVa8l/TU7b+J
oet0/hgN7aFls3TPbNu+4d02/VGn9zbk2zHTXHMe0YJGJh5hWnTzIIB/SakC
r7yJqi3LRTMcmeh0sfQU0hTduncOGI6SetS/l128Y5zmQsB0zVTpxrAvH2+R
hkhhftUvLnYd9hUz+O2tYDCzVavDf4KddU9XLgll5Cm/6abhy+8IX52hIfyn
79kCasi7pawWKNVx4/lyiJ3LxqYPeJe5vC/wfeQBC5007vWyzGTHRQjiNpLp
0X4o7e9HC1leSYDDRPDG74azVfBNXVFSaUh3ncOogcEUG53PFwz6BTzsWJwn
BbzYxUTn2fenecT89ShdhePS9mWth8LGaHk6k0zMHypnVCMYhfrg0hWCQKqb
GaUSh76N6iqxrAeAnwGdl405jDWyofDo2gP9PKO2Ke16QhJNvL0eqMJwZQ1c
bbmxNvurQKqMeUkjfiMp5GDWgpnHZ5dsjni55wx1B/1Xi8MrGuCjcoIWa3OA
yW42PtYKh9P0EIjEe6qH5HXDcE8B/pG1smX9lHmzME2s+WmC0XGEWwvckSXQ
ZvXrvZAc1UoaZE/Ai1MsrLHQnsv0vkVTlJmyppnO+jgFarVZMBoZxM2FQFnI
MFMlE3Kl5HBAYjKAzsYeZgI3TkFc8hA2SmHKKQKApNnBtsTwO/FyQUFjkBcI
iyFj4zY2h5wBPdpqAWXbiBltE8C14QQ1odL0oxn8Btj1hTFoIJdfIVHaJoDj
0rgXXAyqjOIJ0p8ZMvwqmIU9LlJLK/7DwuNiEgY05/9LpKjVPHL+GYbjqTm7
SqTylfE1Xv8fAIHHf9rN7dHQWRe/n2wQqDOMNQreqFRWmuV8hrv+2+z7Cnrh
oc/wxKiG7XO9uSaVuHmDcchdC+14W9WHDA9Y9lKSVbDOTt3EagGVOVtxbJCE
JFpbIG5nSi0Drbfs81bgjlu9S4OFham50g9HsS30Oep1qUuVgrdmPcxhk4+q
zfh/UoEzXDMeSp063QrIgix7dlAM0JB14WQhFbmapPNROMlX1a3AmRjcfItR
v0FF1T+u2jnvyBfzvsUA9KkdiaY+K1jVE2Gub2gdYtyBSMzXy3LMmAQgIdgK
KP6pJkPzzq6/aOMvjuPvLxjeaCpOqnD9WsMSwuSbGWTXQghnfYCqPoWhs7iJ
JUqPwMPDXaXRXoyh6OWaNutHLzX4vxgUnJFnNtK+lyZcgecFsFZoheZKFVUD
UoHpl90JEMWmpd59wyPSys5YsnuLYpqtp8KUUPrh5oWtnxynmRq1fstQLs8q
nEMNown118PCIg5ikJGxzr82q/0HFJGq4dltR2aqtU8Rq6xV81AfycEmgnAF
Aki1P+b+QRGvjMQunouFb+TBZxi1u1J+vYCv4U1N/vuP92fWOUVe5nNdKQ8M
cPYMqB4+sz8eSRZjDtrQoAvSF7P8yfyZiKeQv2eRrMwI+MD/FjBSzH+mT4Xo
SUkBaXO0NIvvRg61DJI2FvEX1BklT4I/4UToILFmXPkF/d/fa1FHXuCAqRB9
2zg0TJaIEq8UX8dyk7mboZrhZ2PNs8S9iaKuDnq/2e8GewRkEZton48ktuQx
R4KTEC/giCSwW5HtVeVPx5rte9eIh91R0x7QZw3nqzfsrmqtHHh6izVTWu1a
ITXWTJofXoJJtPzcgHzcxSHVXxLivHhPwJcrmJgtjOP4wmJwg8HGmqPSfm/2
XY1gd8AmGucAZfMP727wYaeY74HkLEAKk+/TKWwxkycYw6AA/SoQjQBVJiiX
zvTRCs/vQz6qVAxI4yrvZt430JO6lSULbOzMSJyB6hFhJNR6qHaIOPGs4zF1
3nSuQSCpV7PXZHGbSkJ3I30AnXHcoFCi55LLepeXFwInzfRVCaK/QMIFYlAJ
hIpUkU1+GQtrNIYOQ8xy8MImOh74ENFtQJH7JdnOgdGkpaOVSNFP19iEe5Bb
MbwDGg73sJJwoC3FJ00frQcaWacPe/xhQuIa95583GEHiRpukmdASw3XREsO
0hv+mWHVxITlMzBs8+6i+B8VZCHbMIwW32h6UFcQnV2b8erGl/zc/0w3tOkM
4QibUHOFjLQF07N69wmPqM3N6o59Y80R8EOH292HvUGfAkpi4+u9X9wdeFMV
Rfuzv+UvEacE9aKsWY9dnTkeuBZOPVdcin5qrbhB7dheyTNMbGBsRi5JKEuI
Dv4WxN1TpeOee/zGCpmqlSJMc9UWiEcNir+LQ3o4QJvcgf/Qt3HIYFe8JBkw
zJposN6oMfwMxKLbzVOYnuUHMdqzuRkRgBk5342k+9cYpT/rg6pLxBv9jjFl
L6VPCUICis0F0CAYpythoBpzRwEekSUD0DnKn1P1XEROTYScBx6Z36VEKSjL
ccD1TINwTOv3ITnaYFajOfbuX0QII/cjztSd7mcGLHG7Lq79VpaXyMBJQU/0
WD0sU/uUU0ROl2wRDyIF8B05ic442CtJUijW66w9IKdWtxjsxGrhT6C2NZu/
fID0o0p1qXIHTasBvhK77Fd7oIxxMMAN5zKcJWWR/4kKUC+BSJV98QXhJquI
pkkDmq2w48IVOwAJKAQgcIloZXj/oFzj4TV49kNKUQZPCLetjPII5UBJfF3O
gMkCIY7Dy6KTNMqLeuTUDCtUhJJuTNe4YXJDyX2l1W3Ebce5z4tjnFW30mHt
Cs6KPLDSTEs/w4Yip9FTttM7+Bwbnn6o1+lWU7Ho5MxxHL1ZgGAyQn4TxgHI
I+txdCaO8/ofUnH9nyjcgmb0ZV3CVD/LkxB3iNTfUACF+App22Q1yeR5InG7
X4Jbc6lh8Pp4JJlMDnxYN/DqotmlVmW5cT4vNEs1kcpohMt5H0EAI8N9fE5J
HVs9HbYkpQeJk088PlX8f4lLa0bbErGMoIIh+Y5fhm+r9+vgtog0cedYCIiV
tXnBlKAhlpHejPuy1REAknVW3ktQCj8NQaEoZaizt231l0Pa7giHTzd+rdAT
t8SezAy/J44MiLtmADMQO64EY6WoX/krTocnv0ZOXPsQcO/yBjzc0+kdooFM
DQfss1tCTlHxnRZ7Pa6QTfTKFGfZ00hkjSNzb/ToGfVuOtMzP1V83ibl+6vm
zh8TB/xnEGZ5ghtafylRQttehXJB4oVNoezksO9DtRbBTwsTZRpViGJYWL8p
ESoEE7aqmMkrenmVca6exmuI+bm7Qfr6oLhKt52FLiU8kwALrwnp99ULHLYw
aVa2mi8Fq+PAk1y2Zu1Nz8+0P/mG92eNx95kcvL9I7bztqKdgGgsFJviUYxr
T+Xnzo/6YeUUaJlEShwpsyhsp4+20aWOuuT35vvnuvcA9CA9B4V8PigF024d
IwTN+VTatBlNYM2ps0qAq7oPBTO2bHX7yxNYMx2MdAa0ssLWImmI5QyR4f+t
OrBAxoF+5PqP35IxcY9gzdUQ9P0EpEJ5gK4KW3uBS1ontkDewAM+KcSZvUe9
xZ+dvg0Rn5XsQUUc8O66ytb6viLpX+iChVWvE6DNxH9nA8n8SrT02y4QuIPq
WkTzb728DUg2UiKFyqcndlxk4F9jZ5nkFciFWrk22060YGQpCdM+GTTC9nqm
Hber38FB7C9V8Ntx4eEiwmMUYyOgMoXvm4IuFmvnqK6S9wo28Rvz7fzuXIhP
HFneyYfM3cu0Hr3m5PuvakJO5iPgbWdCRVwiZFzIsDUDUohzQ6hEZUaNImSw
e+j0yq+FFPPQDRIF96ysAmxy5nRxdajIDetwVp124Fcyk6mkuk4Hq/yw8UvI
bees4ew1C9DV53/eu4dRiguSji+Q6f9ZmpjD9qq+fCLeKjYhvLgvV/2ZWy7G
/uW6Ljl1Y5nVUtzI11C0Wm5iHFL9rTptdkezB0fB/bJB3YwSS4B5VNIUfdwU
pZcs1HNET/B9WjLQMsdAN/FuWRDN4CCiD2fpGzkafpc+ymywsgpa78XSmtb4
VORSmJG1xHbV1JDeh7JsKhJPPfOIPiTL0vJ0aEL8qoUfXb3db5aXVAzgJ+II
kJ8+7h76KbCYFkT6Sl4DbOSY1UHJhWm6V4FwuSPLEJ46dQ32G2S2Y06+isWB
YX2+dzRGe3FX0ev61OSucnKiFvdG9SZcxfudXXpLvm8+sgBlic8TQrskgeuf
XfrNWFNb34dWL1vP025wTtbz4CL/6eO63+GaZwNYrEqU9MhoqwCqaaGuyCsh
NCX7ZF/JmcdbuPmiiMCfqQSEkZ8Ar7NGfnpPccISsna/gRx7Pp+YFe6INDnM
cN3sHapxscQQXN/cB13/61q3Zx5Yb89ZeaBMXnLiS70sQ/zoT/Iuky72CB3J
plAEWBihtLHyGJ7BZD67n3HugN2F8iRe4HQihj88dZb+1C6W7xv4l0BFlLtK
Q0TitAR8AuwE/OTC4U24Fr5IKt93jxjEjGRkJmCQoG/9XMS0si7Zu9e8DRuN
2m2tJorgvSI9Bhw8lrJpfae7/MqyYsDVEYlpWdJ3JQZdX31J8+1z/GFEqczN
dXjoG6rV15NbJZ8NJa/b5HGjArv6flWIQ69A/Tew4Bj3FJN6RXLk1EtQsS4Y
Zc98EwEdxZE8SZyqbejYjfsA8knBQukQW4bD53KWXannyXDM7WqxCav6yJv5
FWuV6xcn521OaN4/oiMXwMlcJZRArM/jmVouLqz75NO/TZNxteO9v9gPSuPn
Qy/IGVCEVLmFiP3o0oDTw/pUZrHmAlq0Em3cL6rwSwxq57GR31Db/kxvQUbs
rbrGwiycgT7xVAFwUQR+DQTAHTB8VB1+DvhHvz5sYeEA4kn0etgZ6jzQc9e+
1BRvVvKfv2NOgEeBSyla53cX8pFmlVVyvOicLDXCavuHTo6MAi+xq/axGaMg
mLvgGgjF4K0bHftXss1eYJEaYzUyAbqd52fMlv7jVSPoLzezE6WpiylD4c3c
jMeteC5IlH8jm5HPQLxkAI5hXMbjJz1qGMvrbdCMiLxUJJlXl9L9F5LEEo6h
NPEHFGEOTM3M56B0HMEo1BKIU6/shc/MMXjc8znKFF05DHtmxXgwTK9ArYUj
8uZsgMlHQDXm/8zlVBECN9hZkV3Wfd08oSjV5ptXY52+di+JKLD5J2ivBKCf
LXd+pf/HuWKa/SxOHOMVJlPpB3Nfs2XLKaQ4+KDNTcHlIA2HQPpKtRs652h/
gC3dgZoruJ4znhit8szceFfMmeHlVRlhRDT+qahs45uXzwbwwQLtiyWS00rD
0MAEhpvlsjdgIjElryfylhziix572BlSYyMdUSpHetXbnlIjM7tO/oQ53SvH
yz8plQRuACk+wJH/l3bufAUii479n7ZrDpbXQ/VzVgFbpzt5pq/vO9/rtlY6
49xnaG2Pl7iBZMxuzLfaWFPW2zk2og340Axav3LyEx3+V99tQp5z1TwIBkBQ
j+fR1pf5JLxMg1+o1IYDCUakDp3TK5fhj70mT4sfkc4DrpxKQcr3yo7rp3RB
Q46YXaS7L5FRhJK3xe8p6Z/Q4ChYks6X/dA3Jbcy5MTaffcRuel3KOelQ9ew
3F5fadtpsF4uFm9424WMsQ8TIO+L6b4oJi2I35ns12a6bCYY1vov45D7J+QT
wR5msGNJdYihXvZAzdHOXC6iGHuLcpBb71AVlDVlzBnWUgZ7RsJw6b4mT0Vy
0bYZwKO7NP59PPrO8VZhiNOh5NTXW07FLvZ4453TKy0cthzt3j8LGNtuEEZ3
9SckPFCAt8aDLatENwtDOILH0r225VkQg77/Pzb2LlpmzwuukD4ib7/xQo8t
kmHdpKSne30sRci5rsD2S7VbStIAZacP5VYb7UXaa49HCLtQSzWUsLHw+AJz
E7kfm9o5gSUuE0Zb6WtYbAsl3aPJ7tPXpmIvYykB5PnWVbVxAVUISdm/qXSo
169U8boLZuuCnKEZ2N4J9R0fpL85tz2t7SaeSA3jOwR+gMuq2extFMXpWKCu
An50u3Q1DCzFd/r+ydKF+EkgRywQgf8WgmXzyF+jtlJ8UN2ylgFpl0KGT4mv
pUmx1xrLvAHLmyQts0dz02qIW9IFKHHbFHUurZQ22niR+plG5RCh9LBUpJ4t
WIXxqnKslB2e+c+sstWdWTUM77Y4DMh6Ij8lDqb9IqvlRk6lmmgvhAQGlWPn
oDjwT59AaBa4pLea+vbAY7rmM8sdHhxFy9PWAwWRtZziODXX2QZFZ1ai1nyY
vS8Cn6VYepusM/wwnCCWTsOOFpr5awrOKrG+Y74PljOUaW6UvNyooxlbc/Bo
+BqQW3HlRtyA1Df+sOkgiAnCGQgvqiMKwb9rleAECnSRcqtY2Q0mRlGdXKW6
4iTmJkFqmm9kZT5Xe5mL504MCbbkN5Vs7q1cXdQRjr0oaQoo8XM+saR103b4
4ne3A/sburV4zkNe4IHhiA3+smn8vkE5/vMsUuFJU3PtGRtPm1bumzBiNj7T
Zs95tDegBWQkseflPKjeZ7zGpChEe/AEcdDT+Od5G7kKLZQjoSlCJyN9I09w
zE5sCQXaMiAtEAplB6wRd9yak/F5hBlu4jQVKhgeWKQI12ce9aWmSpKE1cij
hwtuqTjlPY4IkMZBB6MY6xOoEjLdSOqhnwGXxnA0+Q1Nvj7esrXfbfWrRlu2
ppd0eztN4ESF2kX4RFB5P/tZtV/5ecUbmTanmSdq6mPBapBz+cINGm9nNK1f
hvdP3H01yyhSrPOzmQtaDNcLp4NSB4KNxJfXnit3pjQ19WQmR2CL8V0iVDwK
PUVCTEmaE72BIrdzyW00SZhaoi8z5/1OUYTZ3eLbOv3ecFLf9qnLnipMQDzR
7/8fERhvpRD5c0DE2rijZRZCaUDnBFQ1JGEF0gxDwuEFzI5B+F6vWHmMWKVj
89tQnlyh6IBf203dev6qZHWCmBwGtDgd9eUMAwRd9Q8oB5tX8LXjXAsKR4Xx
oBXb4p9QcI5e6DcyxnuU7kC1NA+HbY6iC46QXIupyHp3sx5vV3ZcLf9m6uq2
aTZEKQl7hOk24i4XMoWhrc1o3RFTXHrKNfnO1Iusi+jwRgec4aL7KmxWhFJI
gNWbQlu4lB/M/6VPqDqjGxRcQYKm5VN/vB25b4pF1NvRFss5w05xbOZO7aeq
44wNQk8pCdmAdYnnQRsN228WmFiTlg2tCgKAoBoYXs2vemQxD5ikqgo/Inlw
mAGzRkHqZfNvWKW/HJNPW8NH30fZSD8zvve1d6jtAMpqGeg9hpe2IiUw5FIu
hb2ajEXa/7QJ1hhK+ECDQbiZG7ijMIpw52L2p5uwIlSLRM0hUEIYRHDHdbaM
DEuZhXMphGD1AbO1L+d/LbM+2vbPrBartKzxI3gCTgrVm5dtgFekR0gGmSJt
aCb1iOertvuISHZ3AXHV9JFExZRKUC3PUl8x9usKypEZ5TtnRvmlnXpgzWdC
qCC9/rRng87chBckWLE6ZBsQltLNatlx8jztYPcCPfoY8V9uas2DSHI162xp
S9dasSvd/FX34urJIzHvJiChX2dYGLRBsBkPoSZqIoB/Qm/bPWFKJTemvyg7
hZrXR2XLr/4nRryu5/6Px2kCUTQvmPjw0xHeRNrRcUbptjETdMXtuSUzCxy6
UzvdS/sg/38YAE//OAXFwYeVO2bIHg1DCELxdRA4duAyRHFKDcVLjYzyW/wH
W+zvGdmT8ce15SK5VYcntGMbxRHnJCP7XF9Oxg+ZT1Tt52m1BnkVXD5f5diP
MNTMmoDtqnE6SJsXBLag7v81d9a2ZlHncROSKhgFgNvM8jTe3YiunOZaUCq7
Bkypd8c4dBLbXgm0wVO5tYNDNNKA8snHOjncRtdjKJhWVIiyg1DA59gC5FlO
BR3ajf32exXupbo7c6RUor7IGqOD1+/lqGUf5DQ/cTSswCZTq12cIL2UHgzE
pj5sPbFTtwSmcZkQjkJECX07uM8s5CwViD0lvO/6//wyVZH4HpvVKrKl/+WA
05kieRed2ludTDzSODyvG0eJIMSyoCbuarI5/A2gssVvzSRcd6IF0XAKLqAQ
QnIpBDHf6JRXBzjVMWlXrG51JThcgr0+k3BL8gDQYgFe9OVcEXWZWpIL/pDW
obSlHVEVxkISOJKUsuV1SbZe3BZZoqpTSLikKNg/aUi2lU0qfMzls3GbeDzy
1//DRFFINgvmle5ktuD2m/BIGF2YxhdAr5h5+lKRNZLnIu1IRYZuVgrE0AX3
6eOi7U8M+ZZU94Kdx+vqRphHKwPEJofA2QKzjG4timYNqzudqup9V/tp4oyE
EATrUWQQLo41mJdsxMmJpwo7ILX0NfsTPzGaPl6fsbsWqNhDMRIOEFp8udIo
l3Mf1cPtzeC3VVHO6dKdEjtuNM1rrSMDJXemTb1pPkz92+LYe+AmtRXxyd0s
Lg8j5gTsQSgX59K5euB748+kZyahBInOEt2YoeEe95R2DEQ++qnwmX/GsVHQ
NDKYuoWW1NHpG5kTSfScvC/joqno3auE0vKbMOoVbbeRDvsp/2M/Pb69pvPp
fl2iVlvOcdJ6rkyMxjEVSGugyI8xMW5KShtxtUsZizDEcmtvr70XvrYZCSNe
IbuAVZOBz/Umo/5o2sYHjP5PePVhTHORsn8GEf/nvH8JEIuwegfAvToch0aK
Jc3whAhYDn2DUS8AcMCqhHPGDmUdnvo/gbbhXUmoDqNsRALJDcsCMRnSfray
qRMhzHfS+0a2cwzuJQTAy2Dc6WHkjVcud35uTx5llpSM/rtIvTPg9YctPNW6
pqTYleCKHrDCVHn0RbRuEfdy4D1HuXaE11SNu+6J+vkUaO0N4eELU00QYCnm
+qKG0XA6DjG72D2gMpkd70iV6TvfJN9uYCuawF6u9JcqgqZuYmF29s/+L11/
cRSZo+8hUWi8sjv+0Dty6zOd+70ZSulbTzwmmhT4XVr5Sy7l2rlGRShI8li8
AawiYDtoi2iJk5xJph4yRGF3di5S0+SEp6lW2a14ZhpBLA1Cf40MqafLmy+W
tomFlJGMs7l/P/qPOf4DFQU3bOWCYT8f3VgHBG7w6YvaoHk021gSG1qd559K
nErQ2bVUUnXIl4UD3e0RL5yfDVTd1JQ/30Mdrr9HcJzw1NofFT+lhvZ9KS7j
f49Cp+0DpFYH9pdvLiuZSQbEm9WrKMyJKixH32ZiV3A1sdE65ai1/S2A8n66
7+UzckEQk+3SGy4ZCLsclFvFbTZi40rniD+utpJSgZY40Ha0s2WB1dyIROcg
MOY+T4YY6KsW7g4FVp2DNwZeq8ZWz4D0DdOdeF6OPPPd6FbuC7J3toQHh/9K
S5I+Vm2wFBAzu9xnUCF+PYI4NacBk6tEk/aUp/xgwOoEXlhMVGIvPWLex9uI
JYCalOW6AVUiOWj68CUZN/3/zvt1DPkwV7UIFIDhGriKwCzjbiusluhtNd5o
nA+7q4GGnkwYu5+UgA11ASS5+2+9JlYksDRUv2ok90QOVSTu/8avqSX11UwX
FBP1nlfu6v9lDl4x/Uxavqf3M81pHW4qkadOFYGcnGoMqu82WKqEaL4cCYtG
y4uiLlRa8G7FnICS+tLqV+rR9fwvgTttjpCLUlZWZbQLYBDMNbgIoxMO6M5A
Wr3BGXt5j4VWhaDuZXwkWbODjYyqrHwna6fZpJQC5/E7D+EWt8boLu8EOXXw
SEgBl27+akDU0LClBlHeJWK0uFzj2dPKQr2AL6iAS8NZ5abq8C3OmXagJt0l
32My8xV9jxmLd70LiOysVqG8GIgOK30tBzll3PEfZUXo/1eT1X0BbF4kuTAF
PBMgLYK22irppJ9c01dXXKsfjLS5T0MRhrAMXgsQQ5hORMZuJLEd15veH5sM
hfFNZIwJxlplDTHLr73fpOo917tWO4E7hRPl6/XLW6MekW7LujXgTxTe3B2R
e6I4xSGSXKol/FAZynoZAK9dIUP8FGXAQ8twLkFSOsQ9e5Ap0cIFRZ5701zA
urlozRY/WQkhWFcYqUZDSRbA7+dg9k4/oyOQffZwa20rfjteRVXce11kPMpH
+m/5cheV2O78+Ne8pgxxDMMApFWl41Y53QMKb5rOZ0QL1iQbr0DMou254Nvj
SEbMLaqLxr9KJiO5Ju67NrWEAlQUOAUTzRrXK7nhF6Kx+NyNh8ALWZyTxT1N
lUDLLTFtNg4dNAFBS/XEvpwAQMj1PgkrVd8R8mjnh5Qshcfy1iIv8TSI8jZH
OUhioJRe2zAHyR/BCPhU9zIjddYiHrXXQCvlWZQB/ldOcgDE5UlUoR03aDfn
R6e0RgtOOG0r+sAW8GHHMDH96pU2m3Pk84kMZPVAFT0YWd7Qoub35zIEHjE+
PhjeX/VSolgzUFCUtxRXzsFXgjJaYQwBvPAgMnYZqj34eepmhs6KAqaAUsQ+
S6eAsBnXsEhV55YUhZk4C2LyJbXE4GeR51NmvrCG+dqmbZ8uCzJT1U+n6VNq
RZyAvO+PtRENmw0LGtrXEzDF0Lf7a/ZC8gyb9omTGO35YCaHVtXLyB0soOto
2OGG3vHGMRb2VziGa49s3vZqH1L20V1IPGqZ9BTU/eE+bL2tm7ouJEgViAM5
VD176bIV6h3kp/nqFSbJTjApG28nQFCqYeasiInHUVi6TYlTY/Ggu3/A324T
9vCsQ9OhVkLt6ZbUwIzIWMvbqE9Ryj5KR0HbtIVqJSykkmN0hb6sWxBI+VYs
7iKt6L2UxJuQwBrotFhwCO9oJ9/r8eC15v/4jcdbdbYVxenxLmRmq0PNDoGe
gnqXpUGjkPBOynV2foFCPqIFQkNSCqP1oJWNPjK+YL/aHi3jAR4m7yyX74NV
KfaIiDURRkH3GHlXCxOfDA0ZW34WTZx7jqUCNwrEY+Vo8J4q2IOyBsb7Q/Yo
U0Tha70mo0nxKIG1VAUyHAbIlvuLRRASEPUB+fYUABF9MDhutpjB6CmguCtn
pKYS9eq6SGdzzVuQf+nEI5P0XFU4Ll80aysdx1lnTkmVLiCdrXyMXVzx0U07
5h9m20LC/ZsiMfdQRxu0B4jvTsNAJ4u2n5HWFoE5IGo9/msXqnUnfbjA7BeY
MiaAN+i7oIyhnzq0eHbp0zYrR2US/jD0vdm2moIgpkanZJ03QkmIL4snlgrz
1Oyu1e/2ILcMUxk/FEICtttfXgq+oyb8kYU0eCFzlZ5LYxF7erDyjao/tje8
ZQag22DpBtWRwg5wj42LX+/ogtlROynYIZPEWbcTWQOQf1DzOmDLFssiI9Oa
jgWpG4f0SbpAqLQx9pxDefsXD3CDhbHl4rnB9ATwhb1NoGYc7xo47WIo3coi
8fDZ5RagR4e3RAQrOehD+pQfV4E+gOvyVuPUXrXWWFgJycJ2QN7gCQwkFdj/
AqcdzEVrcbw9E8a20cPV4+dCWM00MK2Qf49GckU050W7OK35sivNo/2VOXdg
OD7d19USNIbmo2QEcBUIC7JSaECyLIxJtuFwCP7ftdmdiNeofgxnmge9R8lr
U773tF43Wq8Hrz3x/eqp3FVYprzf/AUFypH6SEw5P59ycZ3fhhlVpbWQ9H7w
jQfcxrBGjje9khAmum6PHHKbrYDnvtTbOOUvya/mSrGSEGVlt4M+/+aB0bP0
M3mfaBRaQxC4uV3Vchnt763yB9ZjDRRSLhOxWyQYCJYgiPL0+RaZtLtBAx1f
Rxv/COp2YAewnTySdEJZkJcZUnS7RciDBrZcfOGySsHhKXDcF/t/QNNkS4lh
b9EotFKPpLT8bSjZusmM4Bx4/3IV5ptjfV3gxi+85CnTDzodHxwtcIUohLk3
Trefg39lZDy7CC3VDSDL8EzGq50/CbzcyMrYDwPA0I3h6nT5nJrGHDje4bcQ
zzWLaZHOa9Twa8tE2s1aSC8UMDm5ZUvRse+28iVGPSKYGKTKR747AJ7+8ozc
pKvSSK4RrC4lSiyybL7FFQnA4rX2Z2ddHXObjgDJtZK5Qe/mM+hTgibAJKEE
c3BqJXskdbWNhBdiPIKBiHQ2/WTfpSNw+v2JJEv670C2H8ji+Z3UaVk41xmD
G6uJdIrFpZE/fYcyUJLOaLkmLqIQlGx6/fAWNESjFyFsqF4Wv/9bs3SnbYzf
KC7B7lZy6CLxpRjgcLz/Znsae8mBxAXlWco86BiPIGkpDiuWGJ47ts1XEjwT
YE7Kwzxv2lTPvD1WfFne0zAvx2uGEjY+6bvcn2mDfoVRmE1pb8fHPOi4lLHe
2U2Tz35XLGuVD4MkGOXUqJBzpcF9culgGhCwu55wyYqfd6os48pxggNcg67/
zPzP+YnDiRfvGqJw5eaoPZDTkCtEz2v/0Odt1OlVR0GsvKpkAN6vc87NqJOE
xd+3mHcTLD4i9cTQUljd5o1Xs2bhBAiUwR9Xh/R14qjLvQxVIJXK65bIY2Fz
mLH6xhwLo0hHNghGiTTLZV+JPeMs1D84S+7er0gH78fRmgAssSZ69VFTmUNI
nbdDvBRKIxsaJyRrlawlwyuzZ5QQ2k0fXOXx3xOmZ/OUAioXnpUULWQpsNz3
E0wwbTxaHXt1YtxMuPAIr/aZQ5Xz6HQMOAD6tvja74exrDN/2zABzoNLq0Zz
jykwyZQQ0AfcFCooNoWX8LJ4RtnqMpOl6pztVTkiEkiz92lsvkyYz9A33yi9
zZk//eTVVrcswSRknOKiiyNVcITJ1YnWtWFKkUemFvcVK91rRAqLKPiOwp3e
0sOxOS+DUzAzprxJIfSwFKdfSZlWU93ye+SKjiLRR8CKb7MtqhJJpqtow45/
aXv649BwTp8GB2b6qlDTsiIMEopK32Qy74m47JTnYrJfSDN4FctphUopuyiV
FaZSXBZjDjQH/7Fzn4RqSy+MXIg9f2c069nzMIWz3vvclcT2tcXMbDhS4m2G
+LcB1KO6PunjUJ5gwPJu6asv1AZVaM6pJnNKkSNHVw/caGCZKgGS90UKN3X3
y+Y+xEiWsPoVfkCjpns56A0iNV27b+vuOqIN6B2h8GRSgZpDraxMIzs/pC40
627dviIXoHjeaTJ5/2VnBFd5fQGNIzf/8XLuev+FiGkLfgxR9YBs3Vu1iAai
cSyfpN1eqZ75tz3VPvE1/nCTGC8AOkjg3JSiGR5juUkKxhITgbkr4Prbrh4a
kd9J1uz9vOqPqJ9DiXy1uhLpiZXpTeFtREvQs1AHKPAd0ildjwS1GcIHIZPl
IHVZJuoa3ZtVpft08tQegvZoD25ljKkeKmTFBDEtmtv/62pl6mzW+uzbxpql
bLRVixD+BjP9MwEjGFPQi7K6bR8AiI9cD7rxlycBiQDVaW+9wupqBIlLfqu+
9RMEQXWQFIIZSLRaSedf8jUVNCjSlCEixGkfXUkFoZSZdBc+hy4NSggZ2o13
PVq47W3bJzL6a8QP2zqZuOaxXBO2qIKVrjLw/NF/DIwclBusTXKo5yrZ2kU+
OggihP1UnmL604I2lKEh1AZ7wvuEVuZYnz842gam9TYDa+FFjcKYO77YeK9u
v8Pfbwqoeeb6rsu3/bXISMAMLOeKmDsirYgaIQovku4Yig3X1MUJgkcyI7TF
s2NIwhIxikl8PcZpnz4aBZteYJZecezjhNYku/wKbwsA2QmGHulAIccb0Yqo
nhOY1GiQCabD5+qWOvwj3LL8yRJXAD4t/x+mtRAzHjmgChskRicizhGMdWa3
r+8EOBuX0WaOMEDQA8v4Byq6SangWoi8ip6EVk3ng94kipwEtbjVS5/0IY0f
CI/YOc2WIpprQmI1no8IM1wPyzFStbN9VZTI2gBT3//HJolRhB3tAp16XcrE
UErj41YrOJeYG0mMcU30YimtXhdmZf6eUtGebMg0WbzPc52QZ97BEQDnKNFO
8RmiF2P0IoUeg0mirmt3fLL6gFU5V2SboZFk/BqKy78rDg18lem+jrUwC8Z3
bUJr3Y7lSoRFRkzZ4vP1uT9dE8cGJGZNa8w1EJSohhAPb+Hx0CopoEROcLGu
NkgDYhbeaCiuSC7LBEFDJYillZZzSNpNzrkK2ONe27hWjefhBSNLKHpF+N3E
ERajS9ncNDRDLA5FJRx32epllg+Z5ecVfMp1QLJSkzD8+/hLP4SXUTaj6gM7
teJM4syzinuPCmP460hnTK6JrNdQarxcnmguc6FlRT49Z6b+sVysysFgZWyU
fDQmaYTb0sFtQMezZtK9yd084PHpipUJ7j6/kujQXs2AbnkHXBsxnO/DqS1m
tHQitoyJolsOP3N5B2HwNoIPwT2EMHWPbtx3zL9YSkBtVLv0HXZ8PmJ5+B87
2nROzhIko5zypE+uHI7/o2P9TdBb2scJFNAnnR6OPeQ/P3B1HFMVK9C48ncT
p4yNIZ43zGIRXjwBp+tiUIjOt2hyphEEGTFP5nC+phuS3pOBU4Rt5rh1Ym4K
M7Ad9YZ+wHLNE+dlv/92SY86Yp0ZbQJGGTXjMyWMaNWjyJjbQFXRAPXCQiQu
jRfkQUuDwvTi0Vh8zzpvZLahiGA5Fn5Z6K9rOz6/dD0i21bzOCNSn/NT2i2v
KQwq9XC+JMTMEDbrzVVEIi0UhEuo7rFii9QFMYdT/ReNMMa9UK9vy9vNP9xY
ytC2Og5HAmEBa+lHR6brHPFImgbA/DV35s7UiBDi7/XSlF2QbXJaqLsLclmV
Nq5uIGkU6pR+NbmiJDmqi1AqfzzIFlKp6iv6gUGc3rAlpETBa2OEkhvVuUlh
uNzqPnKZfki5JA8znKne2DSOv8Nfs8Qs4cY6XLaJOJy9VqcGbh34Z+l07AFK
qn6QlG82zi0zuSCShLHTqRs/WGINWNRG6MNt1dlgBInODOtUkqcL6mAdCHYO
CqK2DZl2iJc4NfBP31Gs7zDUtNjRUEQ7dVBoNgqtFCUA7hfaRD6CPrnwBOf0
7a1sMo9Vs/Jd9y/J4DvwBwV5qOn9fQe7H8DWzPTy3ptQCT9mbhpVbQZlw5i/
SZwo4E9oTYPmn8s4sahIuubTsXSeKsdMCiM4bN/JufGPMhoqdMo8uOxpPepB
QtYX8jTnaDajT8JtBMKQJs1NWHrF55b7PaGKgGVZXEIscDgyMAVRtdXEvqHp
G58He4VSV4JZA0CFe6PR64VpgQGYk0BZqwtKneMeFyg0PihsjmP/6yCqujlH
ckzeW9CHVtIbYxx31ZL23iQU9Yz7baaMioeKPFitzId7onDwzNmFr6+/8WDA
ag+S3BdQEJG0mL8KC2MPkNHKO2OZjeLQCRSpimIcjn/PnqJJVByGShAKxQhg
KueFj+7h0fK0sHDlu33hM35JHnHTtBb7IDhgapyM4VI7RkYlnUhFfT3cMMON
3WjGel0XTx2ByFFmbW3uG+4j/tUodJINd0ILt2CWGv08CnCaQfyUYv/M9eus
AACRstlAIa3CWviWiBtNhUuH2USlZhLAYbePj3fj+hY3yCuinumF5Irwi22L
Xrwtqdzayf/F3aadnN3/IY/ivgx/GGMREnoQwrbT1odRA587TZdxBJoqefSg
GkXP1E9eR95ME9SoiJTfYNkPnEbZNTGZ7RRPbdkC+Ttj106hHzrAH4uSKRox
28OoxAs7SP2qrXvSjXmVMzYkYzRZ/ek527WMiVPnQ/ymQpYWPnoVYx+7QYZ/
SWZN4AW7TkI+5xn7Sx60993HfgvdZAMAMsDtLxNveybUR8mTSaQhTh6xlH2u
/TqVKAkPL3OXx1kAjDa6CGlaxULuGizMsoMCvfQrfH+BM7oM9H97m3IVp+DK
LQQAjLQlvW+pFtRE0CEZFkyIgy4ebDguHfqyxEtRT8KfOwDrRDz4NkEp6L8o
YyG7B2SKj1xWMfG66Efzgq5ltSQ+TsZFUZXvjMw8Ow+rSjsdkq1e6favguZE
GB3eXMZaKs7RxoVyG6Ib5gHxNwtypeRpGHs1B3J5KHx4y7h+tvMMbAHEMX1A
a/0Fs1F7imWrjFnx4AjimO4cCxJaDTHZukN8w9rBlgPjQKr4YA9XJiXWbBiY
QOJVf+2EGHop0zKjUS3sTYJW4GOJK5FNlM4/9jmi4rMPalxPH8Nrb7RTheMn
NnTm7FapBKNg2L76BhEhEI5RwOsy/5qqE7xYHmJ24oNtqHoM1UDEJC8PW8wD
HwkVV9BaDzQXXP5h4kR/4RAb/nFoDlLckQY6ZJLvg1q1fBlnKyHyrBF1pB0e
Fr38y0sGkKnQqZIAcQJlXiyWICtf25oBEsXJBDfo3vN4Sfjz1VB+FhEoDXZI
G39IWdlBKw9Bn/CrLS3Bs3OSEG58t2fr57YqLJLXtW6pqXW3I0Cn9KBtsLVo
DhGX7gTc9ZuwKIi6hqoYJBXTEQS/H3b+CoAe5A5vCoYE6AudWZwfwdMsTvy5
zJP0HvbnoM/dCF8Iy0daMVp6mZWRF8RhQpGWIP4JcpPaUDIZCkVCvy8cHQg/
8Mq/c2agwRW9LLJXmuaYAj6wdP1PnbqS5XUCj7GPEfODP+hke3YCO367hzAS
1RelTclcUxOAmjafyWzIaKofflKlaZoMTxVJ0xegDGIX+AAdhoWluf/Qeaey
xH7BXqgYAgu4WBX2JiuJtkh3PW1jprb6ntFWY7YN/SDYnyQEscM/l5cwYv2d
QBliwFLp3nvs82+B2kjyguRKbP591ZjUAL9GyWc23txwNF0STswmad6+KBkS
sFtQM12vlGjnTzrenPGjrRmcvZ1hZyNCmDxXjpef+z209+18chseZe1tMjPx
nhtP7w2MK8iwRfetENSC3HjWfwqvjd/oIR3Q7/VIaG7pn8aS165kEoYMAhIh
pkQMN2oCogxmS+pAUhqMKddLKamMEkGDJqRWb0n4MQEKg7n4yJ+aT4al4FxM
iDYtMh8Ul3v6d6Fj8oN6Y3cyFTQuU/93m2DiHsfG3ZQ5KfZzX4nnV9JpMXmZ
NQDVpNpsQ4H59ZFFX2NQNKaKPmtv0Y48cPUEhqkvhRuvpcQGeXKux9MRPUlv
3jYAdZ8PwAJJNoX0edO5qgyDYuv/HE4nDlh3MSYIJofCAENH/obiu2uOC4Fh
zjOhV6bisNndx10GW9raYxwJqR0QXJg/HknBwU67mJxwIgk/k08TNu8hZC43
kg8cSQYWSbMSCW/pHr3/Zi5ykYjqxY7n1rJOLP4tINYUuc5ew46FeBcAGeFY
abNbOb5sJWNFUd5RHiLgG83IndAC6ZRA0xM5g16GoG75WjdRxR9bjXkKmLAv
ezQuMfnbJwNQ3vEBqyrCgH8n+B0yJ7I2Lvdp/9pShnNoo8J68eDM+R6VB3O7
79XF+usf94taD5OIG0OJMVOZof8Bm7wPOEQze3J8qW8C0Ier9LbFV5a6UmD9
V7yKzBO1+00mzSlvZJ2BdmjUg2F+5gR16i1pIKbccsxAoP7rjyp/D9Tjtgk/
CBRuvAJLo8nPYF1aMyKDLqgYwsDonqBBsEC7X3G2E521mLMm9hoV9mAO3eXv
2Djd17RaAP+RZMvIFCo9ASztf5gVFzNANt31SdP3Z54cH0xZnpvp1uOrQ3lg
+nU9FcZj/cC/XBpAyQxKT39uEmZ24l7rTnltj5xmD5xd1ZxXEVQ7ldIkIfgf
anK7Q+7lcA39H7Ngiphw7pcXz03upbhQ+4OxhZsMDmx6wCIiw7EfGg5weZen
5/kpoKKgkD8m6QHnR7DBtzkCoN41KjSVUAmA29bySGIF2efc+HSHh9kurcAc
WTwh7/yt7YC3n1xTu3s2Lb5O+gEcxnySfzUw6NH+mEjylHziq9pWm/UqWsNo
9qwmxQcS+ehk5GgWWv0MJgGNexetlgmu6VqvGdT6RJUvpDNc8iFmZ0gFkpT0
pvNEJ7b33sRUvcRgxXYGw0+dKIB7zPtXDlOWCGSViKspUvJamC+7FCCX3skt
pF8x24CKs1o38Y1QcC0A9omTHtgOihnM5lFaiUpCSBrZBxUGAI2eW2AjJvfh
OTmHgMVrUKBPfIo2Jg6vkcPgBmIO+B6gSZT6HMZlG+k5NRQ6Yw3oIoBxZ9hJ
wuGQhG5lNP+FNmSBltAjkidIFPSZHabmZsePvR+07RHNn+WZnr/R7BmJlNBy
0o17Z4VlyRbbSC9l65NI1EMQuYMxXC2lQKq9sL1dfqltc1m4K+9DVX8MJ1uG
qvuVfgchiIrzwnKapmihyaPTdCCMdmwA6sgpoygm0zGDKqf3nw5PVc+EXzWB
7TbgEKWOr1lwlPU9KQxDhf3NyRQ09ZwD2wn8r5QX6wcpm4Q1j8+ZspdOur3V
PMwFK50bUVBEZ2RDwPrHFwxCNq3yHPDfNmSt0SAdlQCdR4kQWINdxL6EJrP7
S/T8A2vZN3xzJPuNUBG1yHONym/gVY9IXxFOLz4MQiqRu9zkBAHcIIwbhR1M
4ETOWgMlQXD4EEY3hHOBeg7xp1dJ+FeFD/nB4aqhB5RA7gKvqBiUDi4Ru3I2
mBYh7v2sUJn8LRbdD8rpvi3PAtN0Sso5LV+YvjmrPeKeTLfanTtpEFPybAPL
DC6HZCCKJJ46tQDCotac0kDwjjxCOatBf4m0WnMt7xssw04EfG3QYtz58Tgs
cVZpSHiWml/47lyCqMYmor++JizqjmxEfuO/CeOCgs8EU9e5n9Om54CtJLCO
HUlWMSLzruYEz/gXsefwwO/RoGno2TIfbzUYOUYwPsVFwu5B15cs84Ea/7Fl
gDHrwfsW/MDBuL23lguctt8TjLdT9ncm7f1+3M28fDqRVlr5QLt/vw3/+SOQ
fjWFeYx6zAhz/cQLEnsZdbnBfforvdOYKkZlSRtZa/6g0RvsnHGkEyacjNyE
/TekTxgcTrJ85TcyRvnbxmIT1xKbtjVxYArgoqe99tKG2B3HtSvKzPsbQHuE
c74XUJeGGLXqTgHbjc3LlJRdZ3ajGICc6PVzMSN7MPQjFya1U5/YYZd6IACX
nMC9OwfAbWzL3LL4pugJlTMOkQElZHoeQQrrRLPvhKCbfMNGkhgfvZKI10nl
ONYQoHx/OkaYfYDbNhJhB+bZS5mQD+mpER+isOZRqMHl4kvSIfRm00Y2R0qX
KmPBYepxjKcqaaTwOBRrqXnqDG57Osr0T5TmUEO9l4NIfyqYaVlh25rdWy06
FMbRWbJe/ln9Yjr3rJF3UIIBxgRodoH1/7f4XUJCb2XPGr0FqN6XsbyIKsiD
Di4x4XrUA4PEX88z7xRSaTpCKYvAe6pURcHFF+aaWBburBJLQKbuDrfPuUIN
Zmi3/GxCisNobj6wYVUXuAcdi6oEBnQEmyxASXUDcPSIbgUi3COO7m2UTENx
QrFLs1A0GKr88TFJ/Gi1MNPPtViG2E6VnuwFkhgA8CMIxxVNXVvSnc7wfIG/
DR7ibQX0fSmRQdtMh1vpfGwYO4cfSPucv6iq/rRAew674LOJhsDRGUNFBjlm
vp9E/gzNeJjqORlHHrHUqRzKiYkBBoZW/u2WhiZlc+/eH3MntqC5ufPLKPUj
SOtVEL6b6TYApUABS76MkLqXZh5F0rlOGLt0ShTgD4FamzDH4iW70AeI2CmN
MHkQro1FXAw4wvJX6XFcYGsLkjDhpnv9dwfVGSq8M5Z1mu+ucGIpF0k5722D
dTkWtuN9R9gypHpwRIHdqSWNrWict+2TNMH74pVvHLgtMQH/jfuubReye5tB
XqMxe+2fj3a8yxkVgmZM4jDMoecmG+v4hyb7qdQoYjv4xHjt0BhOGeNpanz/
VJXPH6H2tFuapRK4BPC1q73rs8YxOPPOtswfoXOq6wO7vI9XJXNBYvH/JrFX
8VY+RjaTcUMTeOLRDu0JdkpuCXFyHFlXFuynMv66dy0i7CUPhlVWiTkHoHGP
8G92ISf+co3b1ADxBJxv6+MawZFBTkzjuAtn3B+f1w0IQM0mlSd/GrpKgxDb
AuPGNkhXKhWleuWyB1H2MnvjDbA44VsBjgYpBwA4iQF7eMeppmrrWTLFkqLJ
WHouulRQs+eVSCGtA+AnJ7qN9dQ7139wH/oh3WSMT6/fGkl9xiVmcuJwyK9l
osS7pvteao864DpZVZ6dN6Wf02ffUjFUJf1oVuhZ0EVdinYvm0Cn61AyQlHi
nmxDDOPcAdsk+EPSJvHMATlzr+JhiZhlZWp19/kWSbufKJSEdpGMRCDsUk0p
AwhisNvedAPRDucAN/U4T6ouMVWY6B7dXhXJGe/xw7Y99yRIdttXwbx3TJI2
jzSOLJYWtlgjBqubEabYUtxbbS+Lvkc5BxvuES8Prnsoq1HJY7pwNg/vUZv+
719NV5uDiTPowhokrijO2ouB9xZs2Oj96HOL5/mHUzkdGy+894WSxw1yp/iU
YvE1V12EI4ezRPlKa+yQ5ciyrg0/ddF65edpVq/BqBZj27IXnciU8wqhz89Y
uMs0E+3Ti9t8GEn6S6fxmC01QWJIIrg6nTCsAVcvSMX5LfvxHWuf57s1QrmA
LbkEK6/deCSPgZCJCS5q7nFA8aKAbguVI1J4WdK9u460gGw3XS4kyFMibqZA
v7FVMYTjQh7KExD9Zq4cCvJggKu9apilj++U/shrOqSbv82Y5evIWDNob3dL
EdTVooJqVbJxQPW8vdAaN6ZMFzP5wToaxbyilmt7Q54qOzoz9OzXYfVHw368
ZW/d9TIVo8FdQLbnxDCAI54iCE7uVE3bojdlVtKv1WFbXTjKfDf9l7o7i7gB
BmbMN1J1rCqdspF9COpnS5rxTHE2MlhBKIdEdyAz/VjUynptN9aXOlfMlmD6
1LEmtA0FwwTEzLMPCj3W4cRFV4AqYAwXQiRodqzc91nSsPJC9zhEoSdXJ1ZR
ciD/JKqmM89nkzilZ6Gjc066XLxFxgJxgsYA1gOLO1tHC2v4otvWvRW3dBl0
Qb9O42VdXHgC0t8KPPX7ZSy/Gk9Wm4tXrwwT84a4joNmX4pAzatOpDiEE+4B
XeHPDcu1hcPHBSCbyxNT1xGE+QjRa3eGbS3C30IhfuQSezbBy9dlwGalp3x3
mOyC3xvSJG8E13s8cUL2srIfLucddR4hg3f0jjXJYlpVtSJ4vrw+PdITRp6p
qHIwuqPTUqlMS4OrFrxM0aI7TSVa3PJtRQGi+SemIrAAAGdN6djtjHyljwPu
O9eks29pCYsx+ma7cxUtpW6+y52r7OvnPzT+dPLX0qEJ/IMJvUoT3qkxUMZm
3DNXOzmYyvJ1ggV06W8PH75nA4A4vaQBBDHiMpYfTbRlj6woEjxI31gy3NAV
elJT2IorgX9CWJ1fBq+0ziJSK8Lu17l2fIX34kNhFXf3f3w96JDY5Q9y6bF9
zLxaAktjuJtxTU9JD8Q1qdm9ls5tzFbAXnJj6rF+Jgj9PDTthU68pEbYrhs0
pm1+B61ZqafOsupwLalUGRbbNMGKF0O5ozcpZDlm1rVe/xUEkrH5z6fjl++T
DedyXehGvxk4TuSVZ8OjolQdhwqMrt4y3Ei9tkT8dZQaHbqRq03q2/dDc5+k
iL7ZPsN0vRaWsnjvzm+grcIpKyG2nGyk1j4B/7k4OiY8XpZPHx9o+rGqFIFY
Z7etMC68CPkusnzbOUDO/SHq95MaPxk3wsTcbax+rH5Zy8L+yldPQpL6s9Hy
E70bHkSPFj4ine9wiVOI6wsuddf8EbTsxvsBqnPgOpoBm4e8q1fofpiYanH7
6RKb4KR4lqfJ6a29pG/5IYjlP9lffvCbf6JmbTABozhJb3M5G/tLYN0NErKu
+gHrz92IMTlM1ossiB5BL8/S/LfT/590djAnNHTDvfSsnDj/RuJiz37MstLm
z4XpxpVlZ57AogEbhDOgUQKLmqFy0QoOV8E5lUaPti4qjuplBddH6JLVjnqb
2QvpNmyluRuhZhLGk8rcQMd99hd5iweKnUhBiMW9d83TOGK7O7yXQWdnxJH2
Vf4vkusirjdeZBmDIsUW+HfRR6sA9EVf4WbMviro+T5LCjLotyrhSrNaoPqG
MN4vePdmJgqJ9OCNeK8IhKD2U+TKpWnwgsUkcV+MnkTi+fkE2HSpoNaClof8
CDSj2uUgAWXsb3f3orrJuxDShS3CLfwfgXQa3Pmee/VVrUpjH62FxKHWXcfC
HlvS5uE1+1G8YwWE3mhFaN5GUQ6SNkJ/7jefUihvx6hnYjo+q2BYM+XWI+7L
cf93/AT/rgKujz1JpNPBbMszdbR3sHBS6+r8HBLiX0dKGij6wyHlRSMTNotI
KEn6+S4ZddfZpmy7bSUOE/SYI3OMg+d86jEeTVZfLLRi0AnmbcX77NQDk48T
obpdlRKfIcm6TCfyZVrQv6am7gd1Hlog78LGfbUOFe0wDtqud8YABqWSnty2
71C0fSSu+Ggr0rmFYNMoc03Bx3C4BVLxLdvguPDf/uU6AO7+FJnSnrJbt+/8
j4VUBorj4ChJtVEAsuiTHU98Wgn1YpA61ATmDqkAe9wrcsVR49mO605MeIfd
/fTW9O7lxgNTzkuOcPCRG+IO8dyl+8e/kkRHTWqJ8qPl4cv10Gfo46y64e7o
9eUAfjJtASsen2ry9SCrpTXndxks1261N7l4CM5naHepa9up6lSq2T91EBBz
LganoenHEclTK8g4g2/86OO4pGjtQ4oFDQou3q7/o6x6xzJgmdjVVzQ8EZCg
WsGLaKvseC8rLwHmH+o8tmAXhwYaQkiQ8q0wTv9VCO8BBxauq3JqQ3pg6xM1
3KfyfQ4RR43yKTxz9PoAwW/Q/sTFZ0utufXLZXFa/fUBTFvv+FIbsrxSWT47
MDEQ2+Olmobc5HJORMy7OES3TXEbbJz01kfahZ+J35N/YpdItqC/MChmy7iH
UIvoXW/gzu/ZOPUUx77pOGZx3uwWppd2jf0ZBpERowABZW9w0vQAaLsxTc2m
Y8xQTSh/Lhod7cQJNhxAWt9RXIhKegSzUNFqPvezjlkf+zDEYfSfD80ofcWS
c4tjsI0nzBwONWFtZS+UFbYOeT8g3MvvuFqLDRyyqAhRUwNqfnr0jkSZVR9r
guMahS8DJv2KBpylwkPQKskfwbrHLxxvi5U6Ls/F9p6vc3uMMXbAsxD6WhqG
/YyRhPtjEHhCyxt3UGQCjPh0c3KRaSib8i3Xec/wu1cJLffPKK2WQSDMHpHJ
+Lw8rUAsfJPfjvXo83z01zqW1CcxGT25RH2knsclWtJ9K3p5GllV1LV19Db/
4ys82aqIoVT0retX/WIVDuZzG3JFQ03ja1CR8m1N4VSjbEooXotlrTD3Ay8L
gUOQTCVWztzMq2Dc3GfFiBbSmEw0I9NOrBJrvZFaq8/XnWX+euNiKOlXeK5d
M6iTl9siXYRKEaUmgZj1P7NEG2SquYjkCRoTI5L1TPGZcy4WVK5opBsv7DAT
QVhCTF5g3mywrUCMjmho+MpvMDdtjPshZNiEzCjwjYAJBUgFkXK+oAHSjDr9
IRbgb31RD7YOfsONF/Z6ge6z2ysC0Nv03P1ASJac24f8M7k4CraNc4R1Q4QE
oRKRWtJ4loffQissCHV9C6P61mypUMBnsFwiXc5sgdCqhAw6OJ+jFkmDAY3d
urlsVgmJY6mT7EEazJxrMI+az2h5EzD0k4/+bqzubtgTRAUaBf0CIm3fB8Im
q7JSe5NLYw52usIK8ReVm85mmnUKHZ/ButR3v10MP87aD2VjDIpXtUSx8tdT
ugCRWqfK6cJ2IkcWNWv3yg3U0tDbwcVHd2FfuPSWNpqo4xY2zeMXSHIrXvO3
XfKvX5GbgZM3V4Y5Ft3c+1S+vd7tvAbY6/J//xhgBbjEDYwxubx6vCe5SBn8
8JZDaIu2XUFPcWaNRcofEbugqg/Jry3jEeuLMyek1UGUxdLmOJz8v9hffxra
gnhbPPvL7ssXk6plFh8u5FrWqW/1JaF9h3K67Xu4PudCEFRGGhAfGPSgtm4X
tDfpTdjme8uhyBwxlMVtWwfeKH5REkaBFC05uhp1B+Cv+pprAIp24EiOv1Gd
HSSRp28N8KL1WoZyiEslAEcrZnyO5WplLH6MmEghp59/vXCyF5Gayo8ht8DJ
QG3hxvOFU7BXv/OI6VyAPdWwHe46+loMmAzyYY23DQP0SOpG8cw3E0TiVUEp
Briu8Zpnzdm9Gnh5z0BQPfxJU4wMjFwu8Ojl2jWorJL2bvYHemY4UxvAvhJD
bwMZWoPn9oQsXMRBqWcIiPqGJ9STmYsyQgOd0pE/RlFrDxNE9H17iy2iuHQJ
Ak1Ai4sKvj9OXE+3SR8ueVEb28SJPcHdrjI0H92EqG8PSOIw6r0nsbtPcjTD
9nDT/MZsbUTkoG6LbXwMHJxTFsbGls8tCJk50IfHy7uFQLtRNVLqOhULGKbk
E0kSMZqvuzDPYcEpAQnNOHke5HJVVZiAqFi0/pXWBta/kXQn7Hdr87JBiRfj
kJf170u1yB8jng0ox0khIZgeXb4ECpedAVSC6EunQck34EZclTbaskir8cUn
ldu8n+kjm61+CBpBJx6xwZIRCBetIHY/jexFWlU11zlc+qFj4E4cxvncLWrF
+8jb99GNj+C8MvgU2s9y38922rtXsPqzznV6Ar1qMPskKOjrX3kqyE5ezA8L
E0ppX9p9vdwWb8enu5GzPeuLi66KfWEegh5/G8OIavb1As0rSrZX4KURFCCf
atv+1RwNViIMZpx++JGrjNAYVr12FWrXald6uiNBR4KvHrxEbBiNnrkpHlbq
Np7jHm6UXr/tP+5jVnOwqhMKjU3yEHzMXPTRhYa6E+7FoxndNAH42a/TMIal
wSHR00uae0936O0KBCq36baDxu25KEzsFHthsOILqAP4CNcvEYMEzkwiRGhv
vsnEj6sG9lnplYcR5PJuKjIfaRiH+wBI81rFAUpW4uIAPkGVtH5Qe5LFdKj2
I7GmljjQTZ+Er9Gk2egGpNvPhsdGKVB5APvUulLqOlD0iikDVHvHETsca/2u
XCPk2qjTE1UiUX7r3F8Mh9P6t9HZ3vx73w1lXKLj3eO7m73U/4g88/27lCSA
tkAxnStPsRWj1vUbHyyidK+1D4WkK9xuTKKC1w/B+ThWqApSTocm3VRQJdyE
QN/zVgjEFbsH9ZIShRUojqbFGSNI3QnpSvCCGriYsVP4Dr0WpENz9qkZf4Oj
DDliIlSlGDCHXucqvbZ45pRQmjAq0YayIPlC+b+QVEJ1J2znw7IhHoQMVI3X
vA74ZNNvQqXruhUNatDT6BHixwqETdLgZ9Y9ZoJYd3LA4b1R1UoYftEUak4+
Q2D2+PBqfzFw3slBpY2zmILCBBi3I6vSyFNn4HPDHUrVz3DRrLeEyNICqU4A
Yb1Le9TNFGqrQ2H9io/BmnqYMH+Oifh1a/FU1jTAEmZCq45IWcCjYCT9jmve
iON5ABPWEGS+FbM5YxAnyCd1XnM9C307q32ysfBjrEE++l5EZd+kJEd5HHTP
8CNe0nO6wiVfqnl+rRtxpT7DVX1uIEZe6rXJh76DNfrvemZUG2NS+PaMTi/l
QGea/0mKVEV6BbdgSj4MxoTALlaPXw5l+iGVtYmQ52H7cOGUcFJgHA8ZL7Lz
kPARgSBDoTKdcHQ/TpcR0YFVBMeaP+3uRd2ZHPJ8qeM9k0Q8VGwZA8vf06rY
FMmGfatjUKhVeAvUcuDHH5v9IZoM0XRBda41Ll2oWxIXe1JihbknPRVQtfLP
K+rYqe4vYmgI4+oADOKMmLfgf+hrvWz80JhNolv44pwX0Nk/khjIZIoAKvlZ
yGt/zus9rWbgDY4b30BK1USiamJKaofEGiWkETxgET96kUO2e9zk6T8w2+lF
3JnV/VBys/yU2MJBaW+isQh6vhfxXfAezJcZtr9kaluPJ6WCbe3fMdi6O5mo
cXUxvghCM+QlPPh8eQM6clf77SBVdbNMa6MEoeTjyk601eCemT92mJcuxEZk
4mJKh87asVA/gYJ0gNy+wBATicgH7lOTEJkkTkd98y86VomhLfwQ353tQVmb
PthkcheuxRaK2uBxMn1SdYu2FK7HmAqt7jPx1oBtNv9/tyJmMReNAbXwe6ig
dqCO3BzX8RLxYtCqMKNNXrPZhpvRaRPAwkaj9ix9LZnplz3QtI2AGgMofWAJ
otkFT7JMTnwedUgL4ahICFIA94iCWEGaPsSCxLNc5PbrGYg9Z7pcw/jHGV1m
sseuhQRcYHSONYDnA59gJbRgrAHpGgsFLDmmSKM6AYASKz6vhXWOArgnd/Ss
QjbMwb5fHX4sh3vBIQFHbWQPbDzzRf4vbfrykIMEhOpHdMJLdkLG99zozzXF
3mRhha+c4zKNHobcOjR/QTFAI56c+111vy5Svxup6XwTKAxjV87DDObUwklu
5yDmXcUxYZphbohgZQnuEudCrNgu8PQJSw7HToaPZXRYFyP/TBrLsuUPoGnU
+WQXwdeAqfO2Welskb96r50R0SkeCbkbttwX9v7C9TdcpG8y21UHojikZTb/
KS2/uPNyQC5GTZE0Z+DEC6jbDrwVyBj8lBxQ8SDstSrj34LMP1NHDqi5LyQj
uqN894VE+lTr3X8lpbAHdRyDP5OXUSEcFXqa7QLX9Z6hRKjqnsLvXvI/sQhn
Pud+Z/pt/Z3Iz1pI1seXIvwvCObepo1UI1ZOTRg4paQUlQ9tDd4OBn9L5yWG
slWOsOdDCnuQU0v5WcKrrPb8SqSvxJKTj91Oal97z5pGhpW4OoNLs9wQ1b9R
MFwu/i78/vO+Oz0opVuWwCqkFNuVknd2zP2Vd0LjuAL6MINBh2LBNS+EwQea
bNt07zrOFsTup0FfVBUAUQ0BMnQQjx/ArHtiWg/kOVTrTLOQFlrdbqgXVzQi
irCWhHWkm8RChBBt9DnWbVZ4eK9QY0TTO4qEkekvdksk3YezO/ajZkD7pkIy
ytYJN++echhbepdgKP2r15vRiZy4VvVZa4hMuReb6LEiinyQ009qBkJPhMim
4zCZ4rC21cbFVXQ5DJwg/4Zw+rFkuy17inHAESxWXJEbr3upryQEXMHwZI1s
DkEJi3m3QOYGHlduw7AweTg5M2cHsyM4J1sPGNVr0WlZAI95/U55PhTnGbHL
OBCnv6KFNxOPB6eSYW0GmwZExpqtf9wyn3BMaCxlrh3Z5B/x2snGY1xVsdyb
J7hyBIGW+vjNyX+qrbgCJD0b+uDxECFnBfzKIjRCwn+F9M2XgSWkmY3IiVYm
bDQLzB1ggGlpF0H7/WRXGTJkD9avx4uiBe6Gwd4Dp6CmdEHMUQGnhvW3gAgu
N8SK2Nf3cnlxpY1bFr+ehmnpNhonJIEPkx4S0GyompHefC1F41hdV0CPDtoy
9YvaOUcGZ3k/NBHoCckcy049dAHncfz/WY8yrOxT3u19jX0AkH6dAxJjLlF2
misqpveWiiC9TuGKZzx2gN4lSY9ZomrYgnXj6KSwS4RrPJx6uj3tCluKdpgG
2h6atwiWDhAKTTNgJNU4JxXV4FruKQzLYomn5x4/QIGI3mzhgMSW/ax+/9/7
+qp9n2zYutHBC9tGX2B2tT6N/JCrWRYjbnsK+HDSjOGuvAEbV9k3xNyI/X3+
2tcGd8RlgaJixPeUJ6XqDUTSAcY5ADxgT1vRscUIGrMa6iSNz9Z5dssYzNxw
8lzKAwKpMud+ldSbH9JGeNn+AhI1VPcmqHGmbNW9tUlf56FafuZt1Q4UcT+C
D7GfKctzBm2l2cqmm7UtG75GZjzDey9dO7L3FB4xwcB9tMuqDnuBZx1cOAeE
c1mAYf00/6umk2PQa+Atp6jS1lmLsGm1w/UMAootWlUadZuDK3c+q+I2dTjK
ewDevDvXlhlmBWMzyKWGbvu9E9eKYI65T21V7SsJS2c6tfo6dLMhARIxYFJs
66q4s25cIx7BHXpwtKKLOnNiEMvfd+2nD5C5klMxDz9Qma8C7uOYcAgvCIoT
Q3ViZbMZf/t/zSz3OicjPiycUmLywLqs6oHBTExm97Wq/7goxokJf3FWM1w/
wFS5TEKSPszDwwrXt+du9/4EcZk1tovZM/fkOsayRV3MM8X2BKNbedsuC+g9
J0QsujAaQXANFH/vxFFzn8BnFq5GiFIa3Uj3tC0euIDn1ieCSZG4SFPjv28o
hbGooDDyJpYjZ0AhRYYLN7zqCJJLiqS95XalZteeO8qojHYlEXG8C8bh079H
9gROWqMUR4U8Zpekblm2XHiARt+7kxDiPFp6wp0KSdQ+5nL+Z0IgHhwRic0u
aTPGe3mVj45IfqHou78G7wjdrfkNrZPHI20ZRXm3rkuGMLlizTCIZQAIucCl
dkndKYZ7hu5mEuahB4LsYA9tKdlfb86CbvDGRVkeSh5liBl1hdEVxGSk4nkN
KN6htVc/F6a6MsoV9nJTk6kKOaZaCVXeR7o2gyJVQImgTYBr6fjuaTEEA5EU
Ek7RQALA+H1dacEUWblolYPBo7ng3pWiWRKSGFAYPeEk4CZ5AVtZ3nRDQASd
aAX1ffh2bv2Qog6maYzEIm2HsQAxVwGfyQgEemVmcb4WeaW/ea9/0cQW7gqZ
N5oPJGLLDQBZMxbYfrmdnMdtaadjYsmArVrA5mW5JN+pwvxhuQHS6x7H5HY1
71/qecEGFfTFFT6kg4bdSIYc/awvMa8XU7cj+H9B58qzN5C7RTejBCeJAOv4
IR2YndSzFwpLYy1AvX9gurKE02wAa3Sv4OXZXDzurv4YdzdFUgFv+0RFCGzT
2QGDDCucTrKLLmm1qAAu97kfeUNe9R+gk3d82HtND7li0qooHlcmFudO1GNm
0TZQGe7Iedn/RaCbuScCJ5bLPE/NLQF7Q2Nr8cVY+XFgtSqky/VJM3eFGtqd
idn7JkmXYhMcU/tR9o61IjZ45yRPuKwLhm8St07GTECx+yWR4OkapOItt580
ZXHdvo8yym6LxD2pouzUBGjRiAG35DZjAVOw0w9q9tqsLJs9aArs4iu72Vkz
rHeJSfEBym03z9BxRipPSeLtUwhebb+24H19hiGLXTLO5zqNvZL1/nwDUMqN
+Xehtgb/a6gCJsaQtdJBXMfOU066jyDnuJNNTapwYRf74B2GaRWWn0BMlU+S
Nj20sdYIaicCWHegmHb5lJisyl12RS1g9Gf/i1oIYZ9LzikfOCFhGWO5JyEU
YFdfeUTAK9cR2Ob5Fawm+0J4EL3xeIHCqVRRv1Fxwb5XqluCikTtKaYPncdD
K1NMivIboj/mR/eEHzTMez7HQsSCcmWL4LmdMdXGXibvQktczz/JAdxR/Dcg
YguTirYYnj2z9knL5iVdVgmDC2bOG59cydyGzQ5dhXDmmB1H1i++IF8kjXhG
vxNJ+AIQ1r3CECC3allZa/W/JYCVlEpWjFsiCnnSlNNqRIco+X/Pjnqaa3Cg
mRW+MvglvAandoDnJQh4epkC/nEXkYLsAygUOodIAse8cFd5mlXRNspg/ViL
Hw+2PP+AY6xbiCFLy57Qv3LXQJf2ri6WOARhDMABxFoHvjFcU7LuPwTLGGwX
bdhmFn9M8nY935XoFUdyQX7GK8sphGvETn44wMdoHAxmVUVhpog9gyEl+Fwd
XzyfRMO5N99lk6AMqnYyhzKAJaaFtH8A+2nq98EnkEcrXS03ODf3M3l3QAVp
9jHFVTM/S3yKsVyGJT28MavzO7DyKo0y45cKklv0EFMMF6FeCjguaJfyJLut
Y274AJXPcVHoshgMh4+tOfIGDWs6WQ3wPPhwmLlAO1KnRV4EIrqPkT69nFA4
ceYmGDNLjKZIBhmCUG9TtSYAx2vTZSrysokh11IDJabBdkNbcbPBzZnz+z+9
T6WoXrL4q3JPZn0dFe+c6aO0JsicgEae5WfE4f1RYgmseGcjDciTL9DwxYsj
/+iiiqlOStl8SIiK7KulX8DxW+lpvoYlw+v8cnDG10HJRtNIhg/ulIitZqOL
yYSaUXfZAcUZ9YRu5lY7amtys/iAkVHika4SPQ/ZM0LVmHPEkHuaWYrpu5mR
gsN3KWiP7HmblK9nookdQqKieBs3D+E/GLXgut5+nUn8iHmbTAi2zFNX3rcv
JJtRSMufT+OYhYf41HG6v4SDqYy33T11QF6KqH+zKxDEi46ym0mYobrRUDE3
A/dxYykz3MhzNTBQDbVPBzPCGL5bFD4zy6hJrHMkCg0xwJRmIihc4sLgupKD
TvyHpJav0DZZ8zAq+5IKyvZOl4WjtX9u8matENlfEx4vOWYp5XXdwjnQl8Vl
SqE2EDtQW7uqqrihnimgooqapLDLyR8Vcns3hrMETX43m7BQEcevIA7u9Tx5
ZLSBNAtH9go4m4AR0XGM59l8wB8HN+Tw6X1nzKolDv2W16qip1RSY/+QVQfp
sYRh0plAh8y7KHtf3/oAkXL+HzMIGwZgoG3fkgdHFQXlEaWCnJwmWokcK43d
pngQ2K2AOVADam4z0in0clhcIgkSAcOnVr+E0m7PCiLgD+ePndrLlEMKxDor
m+aI+ZJJXKHmT7TAJES3dtasvc/aQbz2kgIhgtC07bE7/G0RZITobtaOkykd
iCIelu1+YQTDc0HZc1G0tOK8CdwmL5VD0rqRQaN0bqppGxOK/pCR3AThYYMS
POOj1Y2S2OyuD6AUyBWT0EdZMXCZ1SeZY0q3dKrrkNKlAQvGeknyMiY6rQGd
p6ZzVMn+5HQWHUB4L1KujXppt0Y1gCrtmEAB7k6Jq35qyhXNiy0hoMilHGAg
3vQo2dvEg+syz1pl95mjcMFsgQlisIa517nr9UVd8RjjfN7LqXY4KB1ioIS0
Js2Vq/lzn97PZGy5URCkg3tonZxPNMoFk0KemMgM2qznemjKwe34HRjDUt3w
q+1ikax/cdKFQhmYb1zhzAs1fUAIht7cXFdy8w91lODhRw0kx0b2ajBpU5ga
rZkwiawt8JrlyiRWltllbL8WO+3CqB/WW85LaM7awBHQx0eSecRANF5nCRxE
Jm69fu6KyKuk6cUUHtQuOCQG8ODE6r1cCpb0MGTm6xJ3X3yryqFiVMxqNq60
GO0ys5nvyE0xxmjaX+2srx2Vq+/H6JnKoLEIJNF/i9fjf3zHdGMywo3Clpx3
2hDPrfVflsY+WRtqQZBE5fqcoQWHT+pEjNpapm0qn7Ny7ZTJMjPgeEM4bTL/
+cF/W7ogFNoplijx0/wwRsX/w5WF0i5QNduqQlPvY61Kfm1MGqhMnxs8tvsX
mGfEj7frVt4nXMJZZE+1EWOEaJsNR23vydAZvyVVb8Ltxfeesz7HavSQ0YWr
2Og9DGA8P0/XLlbvzpTzaiqiQ3uVURcvQPEbo2KY1hmIhrlnw55t//9dE5Ab
+D/AeF16i1ndxw9NnpPibJeYphXb+yefUD6s8yh0bwBaev0RAdIIbYlYbEih
dF3ktJ/LEV1ozPDJ7IldrNfdIZMR4eHRj9rCC2C2c8wRroTHcKVRZInQaZD2
i3RwpBpEyFpZR02FZr2qMXPlgnk9RwYS72lvqbZgBcoS26b7EbyAJ6eqfswT
2H5UfFvbgwKo23UXfgzc2X+ECIMMe37d2Js8eCGpVbr4FsuBWwrKQB/pOkGn
8teLCEbqm9B2uYB2LuSfjPJEZaSlxegvcvYXEZn49Yc1AwUMUSl2K2oS3Llz
YpxyxE0zaNevO9qiYiUKrr6py3obNbY1Z8WW30m25+oD5SlyKBuKgdHyDU77
oZIaZ3drm1+PzlZz/9fRkNCbmV8ErKyteI5nORAavcvLFpXxQbZELGaHdMNy
KTf2wmdQGgAaMTa2kd5/UaQa7JhQNasmmZ2P24Rm5IgY4LssrEtzcpZ68V5A
6Oe6L2ZVkLZJR/L2vLHTzaZiuDFy/dTVCop5S106K/oa2zHMczgiQGXIUCrO
+xoF7mV4vCeyZBmCEUt4qYMKQNu/i4FEC3ABeZ/L4EwhzEPf10JN2spXLS7g
iSNWOxOwt9Q9IxddopWO1QulhejYeS+JASM625S97WWzccTuOXXHZ7DT31ft
grUY0ag1DjpSvjpgmD3Eh832FlzNMuW+Vu/gf6HmHCyqBb/YPSg41RXFu4OF
OFGzFigCgWec3y8YwNbCHH5YERcXC5VBqIXuh+PkFIBK+6mqkekQjCdgRA4B
2gXv9B4aARzt9n65mlPb4Ati7M4Yvd/S4BKPhf7KyVXs2nJR/MtvnOBYcF4l
lVymPSJkAJscQESBke+QGey5FIaeI+o6nhIijt6+Uw0tjoRj1bTvzxc3TBXQ
l9hUk3r4PZP7YXtSbw5uwvkb4z11HVH5chx+5no5gnY+s7Mp1PkTf66/0r0k
uK4cpEIbaP+xNqU9M7LPqLnrv97CWWJfDAVhDweNoF2lr16EjvRYbdlgQ0CC
757JgMXFlDjb97kj5Op1yR9lEtLsWAGOh7GzzjSMROOWy7QDyx4H17qqCjxB
nve8n0gqp+dpSBPU2AmaRhf6jFLGHvvdgL5pcmcgA/4g65zU9gUMKIeZEcx5
H5ILlaZazJoDqwI9zmK8YvrWk8BmWKQ1HRpX6i/ao6KClrkWROi78AhalA52
0RM5djd6K1K8HAF64VTaQIQwhGyraKX2nPxClBm+qp4J2n6TOqNK+RnYsMtg
ApN/HTfTWEvlcVjT+RHjVu5hw21cCV2UP5Q4EQpfwxbgHfwlAuiR7S6nEYuj
DRTySFDWCTPYJCgBjLBPENbWWDHzh74AtY1ZgPY4vbE6fzFjKEN1xdMlhE60
tdwAQ+bhMau2zD3CnT6W5b9J8FrvcTNkii+5T1wZpgIzHddOl/a2XgYRwAPg
O9zz4lIFdKKB2OIteFYb09UEJzJe3PVyzddRXsEGq6DtsBtlWmWjOtd/13+C
veWcnTmtGct74U2RXKSzkxTiu7b4cjdnW3N7opq4ZSnFzITprzPZ2kPOXmVI
E+ZefsSOfn3xUfWaLFfNWLEDHo59yhErqmXxu1XulA8bFhUZXSvGOGjcEIzP
wPQyjqCE79snQOOwsSi2AvI25ecL7PvK+enKAMQrWKqNY6imOpRNS+eE04OU
pb+8hjtzTYxIQAq/nCEfqOCBJa6DcL1sOI7o+sZDoJRd4WOLsEHNda5uYuqc
qEBbEs0HvugIpASd71EVaqNvQ/WWwCVZ9mI/TqvH9JQkFElBDXDKOypCZkJ4
P0/GBEQ17In0DRuZf0tdgS4eALTTdVyMPRcXfQkUWa/WCpB6bEYEAlGXJfxf
w7sYH2x3dgqW5l0tqXr+S3VsFe3RAMxBJnjn18I32zwcilFxJMXJT0voyA7w
zIfKGtXTKiVOPhg/HjZSnDm8FGUv5D8qTRGcnQObWQ1M9wl7SDdIif0rB0UQ
Z/Z2plj5Hx7UdpEO3iSV3JvaZksRcoMxTVc7x/Nn1Fi1JPvlUxpENcZnze7a
W8CnHcsDrmyoDWRTVyWHaRi7wsb/ZicV3AKIKfAmsq9mG8qLrS8Ja1L9NbGW
YL5s6kxV4ZFt3TkNNQwiZvFCGFEIZcguk7QW8t3xpSrN77+wihtfCvUyKNGR
alA0yJGtRwhsgIzDLxthVf0whT/0CFZX8dQaGDg9sMak6XCVj/bUBc9AyJUn
P32cnw9pikcQDCKoetdchlOXEyA0JcsNjgh53Rxq1+G+M0OKkDmzhvnDWnFz
1CFsOAkOo5uRRsxBd48JC1vSrsUNQLZLgVJp/uCR6PkkXIE/kFi7KHXJxrDX
d6Ldi+Z5N2H/544ZCEQzAvgMLtWmjuQnko5jtShb9cDwOxPwWryGS+d5IpEQ
homy3heDYrkZfRnaZOQ/Tith5ztynb5ri0zHErWrwm87uQ1zLQHP1nkSND3f
XRgn8wRZpzkr/aMRJ+3711HfDs/GUZooyL1j411lCyoncLQSdw3cpbbyNVhL
IAY+s1SzktpL+S+Kf5DzeLGHUScT0sJ32W5J8EUzyxngNu7ojqTqfiCsabXT
srX2MzVrUGrM92MLjf2dURwcW88cvKEiS7+zHTqSCE0vwVg995ZcEFJtriKN
ULUEsH52OaYKIMPCpxFPldvUbsYB9imf2FF4ezyszIb5i9mJAXHFzsTpS0xC
pX3vE3vbPIfqhPMhB8GZxK48ZEmLABKIAQzRLWQDHFD9LvXU9lF0lQWxjG7K
0/DMD/6xlk22S5kIbRCNuax2ihfGCtCyOwTwswHIS2WYD1ZVE4hVUrublEux
sl7uEpLhJ4aKGTa5jZPil04psbCoCn32cpsAdsMYmI74ZcI8zmfkA9NhY5o2
bSVYtriSqhhXM87dUJqnT50vmc4RIBNZESC/tzPzduULCWF4p/am6pOlJJ5D
NLUKdareTcIzuOJaiwA+2vpVXRmc3VxA/LFKTlVfNd0CbFWUYuMloxMXxqQE
/UHRJuL+QlDc05GxkOzUPosuAKjRwNncWY0WmXb/kP5sTpAcKMoyZiWCnJ4i
CeB1YKQ4FS09sDFxxMZzIDTCul3sh9/dhrWGkPLb2J35z9bC4jndW7C/g8JQ
NXjb4Ms7qifyqrXarhXKjdeGWaKUlayczNHLjH3plT6eQTPD6OgNi+qgS1b3
duHP78J/xNpH9FGjWkZlFp8TBKd7lYqaHXFxTeVRwvU8FsAPxytief/Fy7QD
Jip5Uk3K2N+X+bqpe1+uZfJALAKkqO4eN+Af/zCTSuShtqdlK09v5UihuRxJ
XdfBPyfD/BdtDIFWltHLmF/4OeM1EjX7bp/uykRluwGZPPqg2TEGtiF/BeDs
H5Hcf3PBoWTpPkwM/RYQE16anKsbFc9cOVVwsM1vETbKmxrMLW70MGDrdGm6
qkkvaRkh6L3g+B55DtR2rJkwIsJrk2z5KHwHh3mYF9YmGW6flES4C7CG2O3U
rZKgreuexjIVzOidy7XV4FCOQI7xXQnDKpd5DEmgeCufJeYoVWwPnfViSkFO
/mm0CrU08kBvGbUjyKGuC3IWc3Zl4kUckUedygoDLD4HP+IGU3meFKSWFXiC
TdTpZcIjR7uZ9mFRz6NDd1e5yOKhuDBnZFM3tpzgM1Y54omC3RG93ag8vZh1
qkIcokYhwY/fU1nqkR2XewracIdeg1k40eTniAkuxiJV1GDAsSEvPiRD9zuF
T0G3Z9GLxFQHS6SdDwGXkgTpiD/eneVoU0WyYC2STFfTAk42OPJ2djWzhBm1
8glQDORuTBazC9GXZAMNcCWQvtdZThtzG57cbk0ohzJk6PZMKmXrV2tCpVnO
3lyK1JRZmWwbJEuy0mIxbYsYE030ti4P+j80XKd5E7f5PDO1YinGPRUV//aH
zCcSwgqilMdKIfRu3J+Zu4kEx8T3fW37S2jLQWVTsFbEHqE2VCC0EkgTgOIi
+VYq9gWfECCOzNSzeZRsHFq2gbcd4jU+aBftrhydyJWKHkhxbkUiNp6me1FP
WAffotT+8/F26aS1cC4s1VOWuTY85vjVPgIobopRo3jncQwp5UpOFReWVTlk
Hy27kfrZRXATK3pJxIwRBFkRS60YYQcIvn5zEueS4thBxzE67tRopQHp5+6e
QmxM0OdozWV6unWPvVY5OHRV5E3qhXGkGT/vzeQWcDu3zYWwe6o0yPEp0BSx
OYgZ2n6rmctCouU6izUG2QAVUJyCuk07xopmdbDHK6F2C/xIhf9vk53qkhqo
IduT/SHcb0WCBWo3XFOfwyTB02lyjWB8krhXif6HId7yqSN8gAK3FQHgAja3
g+O2Mc6a4zmgXqKxnrcZB2X5lsF3u+uOhLvztf0sQ/tYCC4yroX3m8u+r8jz
zFNr+zmvxD8N4BXvkoLXW295SEwrAd4kMGAbH1q4rBR0yofRukmvWXfrOc5X
HYGecwlrV3kV43Vwc7+shTtu9We4OHC/wmSPZZcVm+WjUJ7LyvO/pTVmh9tR
jYbbdovsGcK0S2Ofo8JruruInjuPLun4NjrHS55l7sTerjRCR79vsqLsyf2m
EB7pzkSj4Vnd9Ra8HuxUC3bb+hWb36fmwiq79vZwY/s8a7ssp5caUnO7QVy2
DaaxjRNd6Yl1/IpJ6x/TcRfY8Diao8VnAVXTQT6YEmPidIWpVFDsT9+cS03x
jQlooH+S88QE54Oc1Mxh+/S97PMha2lAaIFiSlKc2D1/ZeQK15vBYHqsbXa1
5ZfvoWGa0fpjEIFyPtLB02Rh7h9olY0Vqwc80a9LATB6hTT2s/4aKw1A0Si/
tP0J0frjclQEKCoqAfpfAww4N7Id3ESTtb7/lYNrIKEZ43T3uhVfG9F8TcNP
r1PDmh+7IDILZDghNB4R/pieSPSwni0UHwJHpRac9fP1ucz/fpQX0XjjTf0b
sou8gHyAGW02D7a9A4NPpfcuyzU5goAkuSKi3gXm7ZEKEGv2KSBJpGn6YWgz
+5tuxceiLEx8fqNrop7RKBjLDqdFHDfFRVuHkY/R79fsFFOKYdmit0qqX+X5
MhgckyWLqXu6jBN0twHxghCKSAiv2MU+K5IJkaNKV8gBTG2m1/0eTbDHFD2Q
v3nEsnboHFnkUYIGPbEj0eyRaECeSbq9Hli2tN/6/M5ynJd4UDhfxeXZ0PTh
x6ST+XLOFPho9nGdDb8qaFwKdkw79yQqsdKRJZQPY7Xxf//oCBY7Hr9Vpr5z
osMkCAROb/kBDkaeA1knZVTT3V6Yvpa8gbin19tsJ4VVqpJFwwBP1YIeSqpC
+emUpxH7IDjQI/rvibPNKOTcG+D2W24RykTbBh9gg+WolZEH5DBxwrahYQWG
VRIoZqmYBrMJrQkchQK7zdeGNlIYT6j8ZXg/0SgCM0rM7F/YmUF+N/bdcv7M
UXNBMs9DYVek7bu12THgL8pSkbWvt4xIU+/TqNmMVsuYsj3aO+/fP1TogW2j
EwdCvRaUSzL4ICHDqo7Z2KiW+VF6df747FjjD+PCSrWXEfjwp57ZvW+3FPkI
rtKUq8ORxJFdgaS+L2qOOlY+D99/8eMkHkGQVdYhbX18PXuheq80lQet9Qq3
Jneb0Gc0fce2a6U/STROsjTSddh74pm44s760KjxKLAOeHPy7CU6n0l5KFuv
TD+7PtWSOIs/l+4+hEDbDgjcsFbp2Z+WM4oWz+EVZ47/tUi9VWYqTbau2Ot3
1lrhaEm1ccnpVZcnAlWhH2QOpPDbkyMpiT5PQyJ6gCmFQ2NDLJu27SWTBoS8
2LikfVOjhUGouh77eUVLikS6339k56zOo0o6QuTjobPAS8X317Gy2rQ0y0om
Rmx3WdoaKVRD2OvbQoY3mAYJ9RQMG9yiOwYC4/rBf5poH120MGqYk6Xm8Bms
vMlKnlfFuaYnOPnehBT2pyLBcvcjjQbOp/3Svf3Fn1vqZPNv2vqY+3N+MPX1
Kc0YLOGwgIDHPVEgUpcBGtYicOx+9ZpWyIqorLFWUpkkFoBPonImr5baTcG1
8pVzbjln9omw3c6Bchw7yQzuAcUesWQuek3gMC8Dr7vZgEPY/MBmnSJ+uVl5
Bi5bAp3QIXO9nanb0ReefDbNHSszlj9HS/yoNda4VuilFLMZbEftBwyTAM5B
bVzvdGjOsxmg45Qaz55vwKJQDAT8JKM42GX4HPvdXRk/7h7tq5PAj/BrfKX3
M0X3sIoDZiEYmhB79ELIBWhBMN7ejB7+Q70ocdQ52950esh0SwYvRNWiCZTv
DPF/fEvF+b1ijrPtCQM8QnjQ3qRS+iPrh5Cw+A0sKGhLjFD+PlSNgGyAdn7u
zegm62/DWXkSFpZhqoLobOGKmoIPBEBDKtmDDF+LjYLl+xGbPNhteh/eBbyR
pbnbefTCwb3YyazVXS6yLawcCMVNJ8/q4g3gMh5W0Cu7gKi6KRAb5kFrNfEk
evVgdwOV2joH/irphBVYxbHXNANNT6m7mj0/Mn18Px2CmphtKKqrEuyRltbI
9VB0LiUGH32sQGQXO6BoKHg/uU5yFy7fTmmWibImUuR2ef0b/Lkhw8QFxvUx
t5XRTAlUPejVTXTMNMgAlMaQ9WEvqcEKH8aPt6qVQ4uwERvvnSELnhQn7H4R
m1QeK9yuBAL0i9bKdnqqKMloWrTWIFori5lDj3u/cDuHhNeQuBoaKVR0o+7o
MtTLgAd90KZHZBiHd3jpIf9mX7zIPf1WtScr5Tyw0oOzGtZRLdPc7Sr34OPx
Zl2IWjK1CyAZNLWyGRovr/RMo1FoXSYWKVRWNIAvLqZ22ZU2AIKXwNzPz9YM
cU/HFxRDoOeA7W9Orm3Pwc8zBx8dRN/8hZLbGpI0dJO/WaObdla/hr/ZjPiE
aUorNdklZqqkjmjeaFRXYQvo/B5A2t4YUI8Hfg8zC+4PVHLPLjrVJ5dJpQiY
Zukw6z6RvBLPKJ34mkOvdaruvGJnHi6+7o3foBe21Dnfp7qQtotNjoKkzzRW
hNK/t4cDVXBXwoCS6VFDoXbRfEzm3rh5cFf9onPExJRBFlEocEu2rhNDGkYH
IXTLasmheJ/jYeQnwkCO44hA3bXwNcKdfy+d+tYcCBNgR+dhWBR/PR4pw2ue
Tr8S9TRszcobhuwPPW1Lam0Lff3QAdE8E0OMgEbIma6ZzTEueLI7dxF4HyU4
KWLwqZo45y33R1UXOmfwLA+tSLGSrv43ANqajpUc95d7mYpPdH/b7XM5KptU
Vil40yTiCct6xYgdXHsypuW/+Za5Pw8/y3FTRxQBUciz75a+IVC9q15aOewZ
penSL1039r3VA98VCWSgHerS3WE67eRu3JgoOZaDznmWd0kozr/c+Pxv0IKp
vGt++u27lFw4ftFgwelJv/9RS9wwHTuXYC5KC5Uk8E/nu6fWoyS/d/lO7CeQ
+xQGlsqiZYv6kjVNF70TdebdFswk1CtfkvOp975ak/zYlfkdGrK2MgkVRIQC
j43/zEP0gOIatMpGUN5AO8o48jjTUbZr97Pk9iQowqTFL698LWgF0C5XdfXM
d7SWmOKHpocoOtzmn7dMi6KkeEG/loM6+ysKgkkPLM7Vqt1BAv8B6wAbbGkm
e6wo+QR7j4AiEFs3s8J59//04TJGVG/hSWnlQ6CC9XqPX0aRtcn8g+LYLI2k
x0ijzQp5i/AEdewYCWIYqQhyaejHXgRb8MRszyVLnzZ4+LivjXYlH4bkFeaZ
9oXeMZLuD9d6iv3yoAsS/v0dVOl6CONk5PUpg6XExZiXCHQymgr6+0/DC6UP
L/rVK8EDrNIqn6YbjqwZqdgPRNQSxGjtf8WC/JqjM5PvvCPnBfRQAdS+TeoQ
Ex/s99AgPGmtR6LRGCclqeMAYpVTG2FsIMdyHgfCMvAgQtaid+S/VmuQ+/KG
UlD+DgifgDyiSvpTuKHNt2Q1itKNAyvKefLKDX+uVWmvvnTfDN8mwcIYW+qX
t7LNRtM8Amq4ooUgoSRoIIjs3St9k3hG4aCF+CHGArIRPPlEvRqL2oiLFcpG
hlJ7ZUi6IRMYtIQDxDfy1HXWhccNVUiTl7jqi0RxBowVyF4sl9qEtkB+zia4
DgzH+6tzK2xq+KvMWhNirsC2XfkEY5Z/6WMqDr9UFQTq3YR9sIgeUzjEkYGm
1KzLWgUhQgxFPqp4YcbeZLRrlEZLAENIljwkOl43UD5qEbh0J18Tr6JjSUxQ
E5hW5O+mFfvNOjBzC3BlDcjQHbZ5516El/3Jy4Lp0R93MLSRzpL6q6TqLhxX
NxGrbbOJvj1j3ot6rQ7A4iTiQVpe6icwNsQxI9M3htOEaH33wNTDcfFpDPDq
VvEDEKdJ7oczhWZBv2BkAl0iLz23N80PQsNG+Kzqn6t5DtJ0QNwRYedjSkFj
rkH/abgB/MxSYHNQzfOXZ40Q6GSqLqbvNUIbwPuqRnZDJW+9mUfsGeWBFyeP
wD/sjAC7tj8Gciw4MAMihyvMEH5PH6sYNyZh37R8IMt3TXS5QiFl0mDEtmKb
eCCmkhPE/Le04u+LjxQluz6DIPOk4Bfj4PQTRsayo4oibigdzTJa9Ko4/cDZ
A6heH+r9N7P+9XRqkqqGt8ODNCode+2Z1Ok29jH2YbxFPsrJ6yQH+eaQ8zgK
gsFhH0+Nz/dwyfOCP8Eb20pTNLOnTXOlGqIPpMJSec+VvuRuYKsgN9pCKEsi
PkTxIspKqKj3+wLwDJvfKUPOWZwqwqTr2zkVEyQ/wzhJJjxtpZjoWS4xmROM
gbpglKKyM/tL4OexFoVpjl66xUsyWjLl8DSElLFix3XCj2MtNRSiOfBbNCrp
Xteb1pNv+/5h1tNSVrDeG2sQbciI6CWgN5KUnj28+CH3Al97e+PgBIvlUTuZ
43JAuX7rIxPoqIdnm/CsUMAocbtNVednhUL+NI9AO9V6qw8dsQcorK8bIsNm
9bCUPXuNoAIqEGzcQPJeLSccEw6OgvZXY7rb8QWJEZGIfJGZlmjeIGGhl+RQ
kuQoepW6AGD3q/zNYwZkMJqPHRUaqCcBQPAQLGgVovkGWaW99NBNnzNjO4MV
M8VbhM5+ZjUkBGHj2RXz1X0qnMVFUP3/QqZbQs/PGf78JmhexTVZiMisitaY
eec44mbldTyesJiTisCBBA1U5NC1NMZiBzBkagiThMr9JanwTq+Pn/SPYrz0
wCzwaWQie3jCay67NmswlzIzii31OU5sfKqhbOvF/hN0zOI8GHmk+UwIJp9E
dPYYwlpFg/ZV/nm9GwqhMQIMJHp8g7mZL4SvbNoxKEepXmbsXO7MrNDI7LaV
zRyGPn4aQhmz0dWpM4q74b0j0HkV/8z2q0hrNDvAwN+O7UUVJq+wBAdcVWy0
vE1UySiBaTYFS8a1mbikbH4XFfaVP/NTrcln7Kop8r8XDL1fN6xeBMd50GTF
VT4tAmJiJID2o7/xFzZLuqCBfH9oVflZxs10nK2Txfp+gJAUNxUlo+Ab+b89
FEBKyMY+mfV/9rKTxrlo0efSb3WI2nhwqHn+31mtoXHE6ughy5qJB1ryeCh+
JBfu8wbasyEMTc7PzBI5CKH0EoSWz/Iw+tZbMEoOMrXFHKnCg/5T7vZ88Qw2
549+gXrNZ8irIe/Z23AX2f7g8gBFvQqebaSPlXW49nfuLajOd+O+qX53tjD1
AJT2g8or3+WIV0aPxRt/5mZszcX38ZzaIIdi7CiQ1AT7sntu1PzNr66voiE2
wwqBf4pDO3mfwn98jJ/h+QTIk4AEtV1j/tb3S79goo1QBVgadc4swUpWqpnz
DMCsuV3p3jnI/mGLyNBxSLfitgi97irjGgE52wQZL0xe8OQlWjKw8x/jAhk4
2MW4ObE7RMLSsGzKNtSmX+YUDZhZoEucgCW1+J6WUMB8JlTDIaL03O3n+OQK
LVJFTDefMYt7voqjeC15+wGm2hnjKapg8DCk0QyiFABuIkNpYNcorUmw66eb
y9/M/uCuEPOOCFuCBXgu59O7tPCYXlRJqL4nu1sJCt4PlXiFTxEr1mUWM6jW
AgC/c1CObb0R/4DlyS1T6Zp6YFTETSNXZQjEl1HYgc8L5phbPiVv+zJF5Llt
qvOaj9JUvGeso26PhWyt/SkVB3i9F0K59OoG0v/fYtLsosFXuw7XC4uBl+/G
UicJ+4xgvDgQ6i/6YVqXIYnUvBgKm3OI+88QkRuuleTg745lZI7OCBY4cd0K
5wWLE1P+X8O0EjH0D4WVGaWS5+643qI/J5OjnUJsqZqYiNmL0736X58Q+ILG
CwrjuswgK57Iw9iK7Y8lzaHco8WnBIQ+WL/QOIKevRKmyspKcU6yKvUHXdbf
zAxqyknTEsM/2tx4EYgdYHexV2fm5kSm1RlIbZFzr3ZQ7iMWf2GFrp5nfDsn
QQkmGy1RgVs8gf0r50BIye23SjIAU9hDC4RHPQNVCKBSwSDzUXJEo970v2N2
KDBqD9hVQCU9qlJzoAQyzmTdHvT5uyuoXxJNQ9ymTo8TLhpSGN4xRPonbGTn
4OPzpDnwAoIOfiu1jn1TRvj9FDvPWSptc1hMyXo3+lH0QRZTpQX+swcqOg/H
mWLF6s7rQQB2lfm5sHEtpG/xVuQIUg/m0WdjOOGha6E4PG3PVbvaO0p7xSYK
I+QorjlNrKcmbuClNEsdBmtutNupowHtF5dkFhb02VVcK99owhq5lBxJapGG
9j7F4IifS8jfpi5SxVcPqZozF8JWGYkn0qivqtuS0kRmqrw/9v5aEuQgB6vt
hLl5B5wm5JuEJu1bhBm6WimcUkvQNI5zmk/NBFFN5wWjy9fUukaXjrzJWNpp
KDlBq+iqrmVpJpg7z8TEn/mdEtoJQdXDw68V2tMpEVIxqOkfmpcAFPGgm+yr
2T9Y43kUrT5OeMnqDNRWQ+R4UBDN+L4WDE8cvqRRxFVmpGX7mbLf4nuEy3zE
As4xGS51qba4q6PfEtYyr7GQ5fl1Ajx/Yh/za8SOrt9NV7QeR83CCpDgzfLR
V/ih8QGL0bNqVdSzlfWw7WWbpFTLuM/SpncpyWQPgmTN6jTzc7v8KcIOPk+H
dhaRAsx+FuMV2au5dQLoXK1zXueELMDhtoaQw72Np3xO+OI1pLSxTMD0PQ28
lqi4pFjcKvRGaF+6v6r5jYPxv8lkB3Xg43kSfuNvQFaF/7rtwwAiRMcFpUay
Wmrv3DiSvQLEG3U9IAS1JeG2b90aGVLspmCo2flFux8aQN7VgqL2e0tLEYYT
J1P3kxeqNrWaCSS1qL2l1VIAhehGYv4/P7i2UQnMy1Wp9HZROkqYwCT9s4vH
BbqwPN5pE8CNIOTLDAHAdGqKN+iG8liKUBlXDq0ZBQ5CvPfdLJfGFrlpNDYR
vbPrjrAe8nIR1FXIIQcAwcqjd1VxUCBIN7WLf9huGxFLpn7WP3R5UThXti+l
8fA0RodQNw0ajQYHrVSS5xO2C4M/RQhV7MimtTTusJWelBxV0ZBsLhQxmNlt
GKVRYyz5jOYM4JEJsH5YCEakFzXCa1CKKkjDI28ZlsiCuY+R1b6OQMsl9mJA
DJs7Qe3Xfir/fkwYjI4b15xNO2XCBlbe09QYZSqOJbDclAScbD+wNRjrBOis
5OOyxtB0h+iw8/uOiqoiLHPeXxnofDlxqaIyVmqKIODg38oJsmuoDyCHMjWr
DLfNC9apbs75tFAi5T7ALCr2jYEe0S/Aoo6Gh4ov+4NW1O0VExL0/7uAOoOM
XNfqZRryePNA8do6e9g3aUdTZJyXTprZHoOLXWLllKYFBo3tiifJ3jgV8jkf
PMXYe6UzgI5po8R1ukxMqtb79nbrtz7MtuSVhDUn/kntn2Zm78lK6Ycwy3UM
EeOSCdzHqa3kmI99BnIr6JC8S4aO1AxqLcyW9oyrjHC2p3iPY/8A0sqFJk9k
QkSWOn6MivbEJAZx0xL9urnmZW2rCXTlH+2MhTMo8Ctm3I0PN3Pz95Q/HIqK
gP2iVTuOYEWiymApqGodGM9frX+ZIbcDKmgXLi0/8yrD3594dVUUhbgZKnz8
cc6O+Tp37HkJxVfOSoFuJRVLSJk/pGL8KrFiYrkzJNeVNIP2bbTQO1bpMuMr
nlXlbKE6jB4Ks0XQmngidBpGFhsvdU9cKNO4fdP0/3iRXrt1xl2qyMkAUos8
ASPkC/gvSzElAA4w0PhC16KJjzDNIly7lwa6W+IpCY6UfC5fF96HP0bIUIxK
TvHc8nSrJfLPOXPbGFK87FwN+ffRXcU2Nzd1rQARNNVM+tyQrCIdRoLbB1Lb
qhuyHn5xXrbnv/6DjqnhMNbN6aiZ9dAGYQyLjdDoLC55YiTnuvoVREhLqUZ5
ls1XrfJ8bwbQn+P+2xCF8n28NiQ6iu0bzjm7zutS6naf9wVSN+IWTzuVVOTf
MiPriNKOZgTFUh0kMqvLBHFfsktdb94e/a7Yv2fcwqDSZtjBr1jHc8h4djtJ
gsk9ZRvnzB3ILqoPcTg80KvNzI8j5p39YeF9GUs2CddBGU0hu4I7a7tlYfPx
pBMoIAAnwvgWgrJriEHPs2zh3PYF0E8JE3Ymuvg2a4riqk9sJi/VwOQaZ1ld
rs3fCLBb/I3IYxhJc9KQT4UJdcZAV/8LfFnNo5b3iDBYivxRStGOvBaa2yHW
o+WyuJSpkoufezE4MDTaEklfqpdpjNANjOKqL3gQQjPoqdoQxWly0XJmqfOD
AMokA3Kg1zzSZ/8pvLr5Scs3YVUPgeVbXfM+xlZrRY8emc4YOAATu0piEEoU
IGplfVnD/aR1k6rC9YQU7H3Aahou8KSbIq/HaNjpM2vcbj0tEV6W3vB2ETBR
+uch+9V7cV6d2yG9tyiRb9ok5HwL34rTlGPyKz7TOmsGYABIqZ0ZEoPrlOyR
KzYhIqfGsRvo+mKwI4RerZ9am9/2/DTc/BxGvXCU/1LkXNi2rDf/RGuVybnb
PsU9q7mCYCeiubgAGY/30M7NQV6g4QVr5cBpW2Ruo2pwLyqFtyW5X0adFblm
xplwG86bL10ar4gEnegr7tD8g9IZ+uhDd/mxxKQWrnLOpGgCdt/FE36qmBN7
Pa9U/t6tKl9gDj1zS/bAXXqnHeG4L6IQYRd0lIRYrcvvQeyHspM0q3mIpyNU
rgMOdUFNhugjkB+Y8GqRk5VurKKqFqLrTC3yCCR94PVQ/z1rE+shw36gnlrs
ygzen7qFln/PzZB2vihNj1SWHAjJzvVwHELi4/f9RFSyKKtpqAi9G4LPQSlb
78f1neeVBt0GSoDnU4l/bZiONn2z8jA6Kz2HZASDbzsS2AkoWbLwXFZlzOW7
nqgEkGJeO1xt+/HLVY0XPMj3MCw56EavM/4xz0OEDicNr+gRow5dYJstzZGD
vgt3ENV2jWKhicW7QJqTSbz7YJwdcmfAKWFGlJbwE4nPnh0ZXPQCqPm6KaTE
hT2CcC60dmJS+FuYMBa6L7nyEnTtew+9r8kn5dOq/tRfvi0YeWW7F/V7ijzA
3D18O3Sa1DlyWkybS3vrgVuOmCLWB0YnZe7zv9xRbNPVBAjYudlK8iWA65/L
DuMgBH3X9wujd1WIKg0s5PcmjQzslh+wDru+1tsUz4mlMhGK1XjiJag8kIIP
guzqNm0PEnpZtXHUZfLqA/bXCnsZ20FowLPXPsxogqMY/a2rgQ6XfDvIvgpT
iQH+22hI6TV8boeJFBocwANtiVFCOrh8JATH93102EO45RweEI/kbxkjVobk
m3XiHh3fm6tqB6MXYDd8xST5a+uhLJLe/uLrCjy02/JzSzUOlOWkoL4KYStn
gmfSIW1S2XC02nNtkZRa6Iq3BRIqtckxDgn6L+BbqrMoL8AkGXsxQwMI6HBp
CtOg8Ju+NwCh5d+lo+rfXq/kVMjUBVo0BwWDuIEKnic99UyYFDvEw2lZRvIS
pFeI5EUzTtS4cLX8xuMkD5eBTse6CpA29srmjVqvkYJ7i0kb4d7qt9dhZ1Ly
+tE4k1yRlrpIVnndPe2HhzgSj5V3SPpUhFhOOg09whqA0aucaLKS8NKJHlcM
fRbpxnxs+Vsj5AWgmWYiPg/i3sWVJRCYAv/DM19NG+teUPSyj3MuvW2AisKO
CwJVI/gdhcLpOJcz/f+8+pPEhARSLIqJYgTA4XNDiLPcKMXu+R/Vdrplo5Ru
1FKkqrUzqy0c82b6ZAMaC8c9Y9CQVVfjgnMjpDsWA/UPWMYtqFk64IhlDqsL
Q8p6XHrBIiixDDYib6sW5OGkL2hdKGzJ0a2e3BaIieU7YEzTFcdrkr8zXhsQ
T9Wu1rxcRqrz4XPpiZlA62rE8b6X1CU4Z73nfnnmgPCtGg86wdF9io9J59Hv
b5GvHvalJOoLHIFcp6abJNelvOgsOMQ3wB0h6HTFAb7VGq21uF1cf2sK2IB+
ThQyGuXAVV/Z9YLIpofU5g1HaS19J8hZxR6EXn3KlSNh8wFuF1h2CRd+WIAE
7/e9NvS63v7g4XNO5nD6kZcb0DgW4PJz1i5k2HdVMu/pis/Cz7QcBJyIzDOY
YQEh7ZxZP+AZfWEDqvJDS5Lz002WT8iNmHGifzVjVjbhb/bUETVPKNGo/AP9
gF+dc7othMTNAhXm2FNgUQEROGiEXPxHChBFzPytaMFQ+ptzmZzIiy8XUKci
XGfHlGUBvpcrYkIB/KTOCbRrEjbHW1ZWlNlGTZVeDui61xD/fEG8P7cxeuYK
PBZeoli40sDjy7dNvmAUxLOSZtkUF51I5eLo2+hyXIRvux2/JA7PYs5R00sE
PKJi4UIDbBAfna3gfWmTqjhh2SThacgxUUmt+ZwZSLbu6KGWoJHWlCeg5XUz
02smRGlbXP0AfEQh7W30b9vofhx8EMxe9dWY2UWoV8C7l96UegXKqe+bvAil
oTQbHIbEG6a6o3hKVV/CoahnKE00JevQttLuPHWwba/CThfkoEKOQDLoj1tu
IoMrXM2XDX1JQf/UYWftu8YXJavOahGcCwlZAVFT/5aatDdo8FhSVTQUUX8Z
2aZtRoLcyuOrt0Y6y8M5C0kDXEEipYEx3mGPECcIqMt0QY2vwbJvBmeTf/gD
JF2dos+piqBKcrl3CfN2PMlNaNegRPDpR7gs1CCxaw2pPvXK+yA3whSIZwp9
9qettjplkxyKSFWETh0daIaFN9i3UXOe6r+EFrfrh8OXp441bXHMMtmtvKwp
7Tv57f/zoBPHdls07k+0Sni/AgZNuu89HgCEjBPGjMoATJJ36aqPoo8Vhquw
VAvaN8558JlmS5uf/BQZc9Vu2uaPdEZIT/d7Gn/Ty93E7lS4TFNLFPBXGRdf
XV99Bv7UnlUIGxB606KK3e0iJJC7C5kSZ5eVJjdHSoa9VNAU0DJ7MyRIWI8F
XaWXZ/HDbclzBtRu5Wt7coNIeCUmLupg+0GkteY07yDXMJ6fU5XJ0KtmnT0l
AnO9c9v6RFqVSMKmly1EaPcte3b7Ey5mpYXQ3WVfBqjGxAU7Qxx3QtSUFEIJ
YgFNSQ1Mrm9PkAleCsiP/Uz93//0xbftn18OTiuzyXCTBP/fzD20fraqCHNl
L39iePGOlEfEA9unwwOYAXjAR/aEDjHRxgHy4+lGCr9F/Rj+0BB+d6YuFLVE
adRKJZ+0VGVL1XdZI+4haei0pY3VslAr2GgQDdphj5tnp0icVuOC7NWj0ZA0
/zTZXWqK4U4/Xu/15Ai1kdQYtEI3Rb4LwS/z5NW+RFKHtDpMkzA4Af2jviPA
hBoBahWIN3sjpIZFg3S+7N8BIFmgeqUIM2muRzGVLcGIcGXDRVRYLt+s/XMI
9OSVPLTD1lviGo3DPDORLg6hKyHFGN/+o8xOsyjdgigUF0TvuJE5yMeEEL9C
A3AR3PHcg1iqJU/BUcJhk1cMtTDCVoZ5GGSOwKXsDtJUwu4IZabUDnvmTQLu
hlGQUTB1aqxL31Zw8abXSxCn94Q/NiWoMA8j5NEWpydWYLIkLyMW+1Ydv9Uc
+nYXqtjZLDH2y2jhwRBPB7nEWH8ivLcbcAhGXjIDfnOr7QaeFI1PF/pV4VSZ
xmA/UAzInroSg7xS0lJ+Dd+lnE7solhslne+RxuNxdKR/Shnd5M/eu2Oi0kc
v/Cl1b+4joUQa9EoWv4vtAQoA0L56BgHb36XR/HHPcVC38nxjZQ1ZKB2OK6p
2UevdbWmikM3rSOZiq4A1OLGM4xkfiCQVq4f5mhHg7ukp7Kaq2a3KsO1hcdy
R4iQuAGS6py6RVWubpcsXtcoA5ZSwzmmvt2xu405W+xLLEisc91JsNojMxpB
TbsgXSmHc3TAm8JwHXwjOy60zlsyJYSnFich1IEkJUYr4/tjsTZ7t47gG/MW
TUjwIOEersBBhHSbaO7wJ9TzQbT3sD8kXOS3iKikj2oLORucuXUAYc2cjorw
2f2gf9jIJ1eRUG0PIj0TacNOL1Xjtc/PjUrG58S6VGPu3FbZiGhqVUDfS+Qu
YrHFUEuXKJzrvqpITbJ3o2NMeaGnOwfDlRzfKlwfM7+3TAh8DX+vXj/Y5oJA
4Pb9oUF6d5FI600gUAVawDtuFTXdzrCMwsFq/n3mLOtk5XA9Drh4ZcchwydY
EOmZKdqOgSBC2pq+JkGSW+9xZn45xi9GjZypE3F2J9PDsEbFQs2pMAcbW9NX
UfB79RD3IZe0zr/maSNgKvEZTQhxaBKzBIvWOP141IGQ111sroKlFnuSW50Y
9CjPFfk4S0xUwpzNE9I6fkcO9hA2QOIyok1fJ9tI3biyUaMNS6mnXeDuKbhH
+Z4GjBZPFJBC0M1kXCwpX96szUS+371NEM4s/RVqYLPcWtz/UvS2GanADmMW
Kb0lRGnM3X2JzdkGt5ig49yoYEjV8yyt2yWLPNA9711lsjuO9iMLsg3oj9cm
cn8/SMuVuUiUB4+bN893tECRx9uKyhX7AQCZY5VYvGNnecZHm2u3JRwVGOIT
+EDsCvRzH1SXsP8vzhrY75bH9AW42EM0fx87fIbDXt0HmTQSzx/lht42rXrj
vRF8KgmNXR1Ox8DSDkP7s+7vMahzCrXec9RANqR3nE0GY7yHiQSZN+n3Nn1D
+2g7+dlZLtZG5+d7mAThdNaBypuAlYUN2j+LHoU0b5D7TdR+YQaLcRD95iwP
Or27DcG2eSxln+11XDw/Um7Nij7f4kN2grlRrNPOKzP0O7ZWAJxkrZ+Vvmrq
X26ewPU3iYZqrPZR/iEXxaHfDjzncKZR3lBM29NOSmRWZBbHePjT2cUz53Rf
RWDlHQHWZMbSGudb1kJFqIyVs5IqTUmWnfkhStk71+j6KLs81Cty6mSL1Bq9
G3BS5+CQLwaSRCBOESgKb2SApfUcqVhDlvswmAo3ks9+0X9tRQ3zsQFXXMTN
GfrqXG3uNu3UjmrQfs+I5CMQFlHwWLieJF/3GbOhuaEGyAelkfYitefZ+Yy+
v+UnFs4BiCf+U8Z4m/6XOwdXAXSY6lSYBoTmDShvNt2bGmpH7qG3IYx113/a
jFLihWJrd+EJlEmVqNu4LgJmL+gX0u4f7mcPkbFxijNkbpvHiMxs7UKK688J
gbDdeWIeEF5acS5knJm5me+ssRAcEIHcGUmqp8K/58CfdWfK4t8ubQmYF8xU
Uf6MciThf8i9E83sPeVPNYg9UZqKIKqo/y9+1trSsTMi3chFyjR4JvuFvfbS
IxN+s/x/6P/Mgz8mkBT6z4L+2LbWFsWDjML9NPgj2tohz8YjUmHBaXiyW9Yq
AjwGS2G+yChzDvT6O9zuvQd88lLoIyRGYQCFIo5snzoxNcxOB/TnA5WuuK8a
MGd0m0IL9lp+cZOXjcupsoUn9DJzPc5jpjV+DuOEX66cTxUlYGDuUO6SY9IG
+ph/3w/sfZ6tc0JyDPI3l8XYTH+s/3Vk1g88LpPzpAyqNkcoIQUTCVlszMBJ
1Sb2MaFiskyC/mBV7lFAYVTZRXP7n5ArtKNTKxw6j+lD6/iQ9637o2Y32jDQ
iUPVQvF2Og/3/rrLRDU9hrnkNF5gsSO0xbFCVtJ8ybgwlydbP7czPix2JKOq
5bEjhwY1CJPATj8Qy3AWiId+83zbtQlXdXGz+dMgWVQqwSQeH+TTqj/fruJx
UsjS+OFf3QinoX9PHSJ3OZpuyVdmp++lZm5WhBbLJNBKOPS4aQPHymrRo6LN
FUZw7qiLqqLKm0ln8FZm6SddwfOL6OU7db1+R/mTPD4PewPwqbmBUywJ0+tZ
NCMiWf/nmdM3ci52yQImjX9Cs3TkwoNDoMNVNSQ3bNbKK0aP1pRohnb9xLdL
adyXmMY9jj2+JQrCOrs1TsUga8NE+ZMtvNpvoXXp29aWTu6G0pXwTGIR2j9T
DQXehi5yn3wgUILXnW3O8Das3cM9RojeWXbR8UYHyXazPgDnCmznL5aa17Zu
+9sR+zUOCzvZ70sjz9bvAzifzr2CeXklui0Wa2FOWGsGY1prpw/u8Rgn4zL0
UINignIZjnI9+sedgnMEBXkL5/Q1qxYkGP7f1ma3Tms7FgBF9NFcZEg37cyR
Ni0TWi4M/J++GzP5mA3lN0MzyAEX7CoW/VGKZ655oySQy4xtx5iADf+fT6s8
Mk3S6k5Cizm3NN4PN+znAJYdcWohdkYsee08bGioLSFpe/BGv1gsMdInWEBc
TBzeLovG5rj1Qa7YfpFnSrYJ5bt/9+LEweZcYOBSo5gFZRkKK4AdjJpveskz
Q+d8oiW3zWRopS/JsF5MSr+5VYL7YzeIR37IlmSGEgxuyz7GNk03xOT+4PI6
5u6urWQKrOndc8b9XVVwupaWA45lC5lnPD9dn1TTofus2GWBOYdu98FZN95h
bjxI185c3IHopKhA/xY1B4X+bnkHl5KzQ5mTeGI5Ylm6zu/aNbmF6UpKAH5R
WG5JvA9vZP+P3N83ewLERNqVeB11k2My+iaKlm33/KfgOrT5W8/fU5K2NViP
Us+j/i+u60/Gq3+Bid4dLv94F4EbBHRXKhqjQCKcS1rsFi5MaGuWbDNkgjDW
hGvNOstF7dyc638cnuj8snrDq/BQmtGKLvaNJ1b1jHdBCIOulVIfTqyZ0LOZ
IS31opXdaSvW3xKk8rvIlAn9jCYGzJAVR9SsjZFbS5yFU6Sg+HzjTu5Y3FTO
vZmJuVKP1j9zwUdWnvjaGl1JcBoliGFyYNMBOWvLRGq3wfV28cl+smXodMRk
fC6p3n9TspA32pUXY0TlR13hHB8YALSX9WTsgKy5JW82vcCLZG4y0FPKaLSi
ewJs8UKMZPbJg2zLwXTAT6o1bo5tiCDEmzwcMYORNQeGzFJ1LYvgdcWuPxU3
E9/7JLGUE6W0dg6A0aa4sIm4e2g+l6QulkdqJqngHPsVfyKNokARHXnBkmVm
Rh9Rp4dFYOiPgHG+5/5k3oIoTH770KDAU7G1mQezd0+fN6K6SPkV3KvEAtcM
tEVvC3ozr6vRNeXfLa5Vy3hbJzMpllxXho7Qk4gNF9QmlxnhbMnAo+qI4Hjh
wonXMxZLPLW8QeN5f5XujWJodh+J6YRy/Y+tJ2r39B4sHciycmrBntwuEglQ
EbpYEjGJPSHjWJpmayKj0mX5ESPzx65ZeeDyd5jCOJJpLrDb7ZroPxXch/e3
rivIFZJIuDWNz4z9zuQhHjvtdo9ZU467uUTUjKB0pZFMD9xMjJCBHyeay5fF
JFt76bUU1UmdboIEVshKnjp77rWaj0m5ITMzrcMHgQcYcBoQEWBC9tMZZTLk
ig7gXZEC7MV4HFkzCx/iqqbtlGWMzxdsYKgwlcuFJw+y4owEcSH9RthgXrRG
/MIBsBJKApGLI3yHHZwdOOgAp0C41kCvcKvv9C+Hy/MiRQUosn3lVSEuepX6
bbrkfHyZYx8gSaMCRFTXQaLSJIwYbqGFzPKB4lav+n3pnsHCt6/8eTbkvtD6
wM6QYnk6I6ZuPeEm6QNpTFRgjZKcZWKCDCSJwxnvsq+BIxkfzAO42lODmdyp
pY0035VrxjQmyN5LyXbZRzpq7x8ybJRcng8XdLx5KVDMRgyxMe0c23m/yvG7
8gimAavvGAn58nM41914lLWj4Bq3gdqRFDxBjlulIYDsNtdpz0xrW1R+vQP3
d9A+tYbBrcm8rwFZC3B2QwGIburn+EyXYY3z3onQTyowvYb9rV22ZRzm2vU+
yuyZRBkuUQwUJqx68I1PBs9G6LXp/ZJ0PD00F/b2RFefso45bE5s/dakYMk+
sYk8AzpWMO1TyJ/Ewfp77zZiK6DhPQBQ1LmcifyAcyNvORntKz0x3Yj9o4hx
mMNRfD7iduEBsnMS+6nA9Xw1F8h13MR8FIRjMcXhyAxhRse/0m3k7AwGn0md
T30j25VeJ6NE18IsOz99TfkpzlqbGUSkBuikfXUuaX2T5l5Wna71z15iOosb
IhLDk5HW2SDaX1SXMZGEqYQ7TSbK863o9gm9/+JriOPkIWgzFCCUePKy6wJ+
lZCgJ4P55OpCYNlA0mQWMXqBNzxcKnz7y8K22GllJRjw3GCMaq5H9a05TlXI
41WE9DG0rGNm9W+FaWEfcvO+OaGP+cXqFSajWxyuh0Ai/0r2y2w2pQR1OxoI
/+agtEF0IZE9hbC7JtECKtpVwDHbxlIEY4fnplyESxfIzwXJpKlxMCCiXemq
A33qYakZA2tvSr5Ii9hvGTajCOAND2NjccI6vBmt8v3Hz/eXIT8K2c1nJvMh
69idDLiTkwOGh55Mt2z3JrbkFvqqHY9NfRD6sjC5CjTzUMfQRNcp4PsRfA7v
z326GvHQThsx0tR/ETh+3Owab7B4a6DSAFnWckdYjn+1BdrtS+1evoTGk+bD
QTkilGgfvS6qzYDWf92pUD/XAayIIUOc03axYVDwUaZPjJ9Z8p43eETP9Brn
QjWPJdqdGsew0zIpQiUDYCAwAAHmSfOHYhkAntcpHfePbXkjQzFq3qgnpYMs
K2i0yK4RApbvWtzmVIvA1zvfUJyTLcB3X8ibgQA8/e9HTaCwBkkmmkU0LGZQ
N+7N+KLYkuHWp6EnHz0l6i6QTN72/zG8s15ozZFSvH9JFXMPJJh1mW9VVLU1
gjrV7CltBCwnPcpiTvAyUceyMCRVBK22d3ksh9Ml/zsyaIazeALWfGRoN6Tm
c/uUXrjq1ko9jqe1T1pV45MFcJLPjKKBCaZYOETUAZg4mKpJMgwPtI84DRmE
6PuD+hIomfBOVIS2JQvp/XGClA4cWgygKhmLNfRjdjlkxvVB0xPNF4mrYAU/
xwz7uu9AYQBhXmj6kBlHgfDI7QVAvitkGJVofq3JlRc3Ct6xdvTSwFjhQhOZ
3Cd5cBdREoBZPppsPKKge9UkucnNpUDW7flZJfhO+8Z2Pk2/wOv1eTWflI5f
4Px5mLJPeFS9T/2bPIgknZl+JfqYRgW4WD6FRpRTdlY4RPrIxpw9zBhAZ10p
/ropESI2FrIbzzYmcqsfNntN92p3ZjDjchmYonS46eLAME7FwSeBWXzPQmxP
bwRy1uOrGpWJC+kdQ87mZHscsU8etGgBQzMEHecbpe3CaUxCQRremhimzioc
Sd8KEIoCkdomTYnl6VKzye8vq8BncL9Y7bU+d7ETIqfNpxKE9eTIO87H0Vax
wpYXOcll9zjj6MJSIiUAgfzyKutPQNh+Hj54GakfYcU4pI0fM441vY1oSvGs
ibj0FAJSQa4vViLP8jPbS2MV8rtf1nKI8/XAEQqps/GJ8xtggQJ2u5k/Z/pa
iwgug0pwOVyvzgvDg/5VVXdUl4CUMcNRyVscAKuoLxVJ3is+jUPC7ow348MK
d4MowJ4bhut42+aBDFJL+elHemSkxtWrDGUVeU5SClrmZkhxF2TZsaB74Wdk
57NL8p3J2LzaM6S1ldYkZMOM52rlkEArERKIsCEz5Su46FoNiPTOK3WEtL+S
AHXTCGDosLRNJSJWiK6hZTZws5LMhOqrdj3viEfTXVTfZupMjZAnq/zBAOyY
2XEvsE+FhNf8QSzjxslY8MCu6zQ+mkmSv0EHuYpZKJc0KtLFOh9OEwpxNLVU
yLIVS75IsWDIifg7eveOHOrjMnhPysXfmB0Gzz57hz4T/JFxHe8/5DAQOgOR
8dtsJEhOFMzDiltOvDoYdPz6KfOuzcHJVsvKgdzlZD0jKNDZPkW1Pj7rvlGd
xX3YvCZOMlnbk5H9tZ0MPP5TP9CrxDKSDAUMAv4sEH4P61lsPAxcIMk54AYL
3GQjakQH0kcSLWw4VBR6NKvbLk39Mviu5syX2SuOeTERmJu8NDr4GYN23pd/
xewfJlz5XghW3tUG/BfHjbum7fjELgNyTumSnpLllS/0hKyMFAtGk/vdacpG
ZVOPwr9R1nWQL5pOdOurbfEAGvXk00uT1hbg2+lz2lm1DrSazK7sme2C2nXk
uD93wK67y5YlKinas2xyQYU+uddsyBtB3RIgZHxaZlKLT6SwvNaV25m6k6Kd
h61oxNTaXF++7u+m+UZfu8q2rcQJ/t8C+PMz7j2wjH1xsMSfB0h0pGV4lJoS
ctsX2rKrO31CFncXlWuKhcLrShUetEhfN2ZcCjG9JZyTnVbf+Kq6ZsUu8rz9
fNHZ0etGhloBG9k61M46KxyFlRe3w6pOiLHfep8zNzBBX1Za9T/26yG1IBuB
8iJAO61J5PTztNmp1742+9m7aeQYHx9isw3tfA2WswLUMxrzX3YpWrlgj5Hg
BLhSY62QjiXFRF5QZJvzSNLmBj15CpldTXfMPQ7wuewqivxsBPGseXMx51fI
ztIJnDnvMPHz/b5hl4vUvlXrYmN91eqIEG1DJ0Jfmr7chxIogCHhIMBRFv6Q
e0PDa3Hen6mzRBJ3zr7HeWz8d77zBf6svbvNggn06KiwJHEcBH+kzaCQz4Lp
idPB3/+xeN/pg9cLux5mFPz1sGrKXwqygsla0A8+QQCHnMXtM68OLZ5LWZLl
iC1LK5py8d9hvOrzWgpSjbn/rkIfYwxCOj3gupLjnF3aYQRHvK7WPg8p+KJU
RCmUrqXxlci19BcaMuDd0y/pNyBNcjLZ3X1ZG/64UyX3SrOnGf8I0CuXL0Q9
wUmCJKC7WdG/Jhz+hWeFWpQGMb4w8qztN8yO/CH/8g6xF+B6jpcH+GxVWqB2
Ofbe0qxzQckf/Y7Jjy/K/liOZkhj4lCtGQUhAe04Y7am9t6fVNxb74/QL0nj
xyexpu3Vjp+prXQYTTvbGBSGLApkG2AZqBi+bFILTP9O4e5pENv2cQoQjPfr
/ph1KHc1fVLfbfMleBMYP3erU8XZpdlZ8Sp1+CRQCPU4d6FcEWHrw6jijMtF
lE+vH1aLhorh5uSE0CKmRm5zEkyPbAbL95OxNk5akyNqRYYwVEltJDRyr5+A
Y8UneziqMAzuBq/ngZNSf14NgjPl/BjASq3CCnB2z6a59tDWchD/LsL63jeO
EDPXD8MHFwG/Lr0THFHhpyQDzIs5dvoxci9k+QJynzIvr/rLF89XmzV0nh/8
9OO1eJAKPixSUTcZrqyrCrm7KnV8vMmV9V+17v68ir52j1cR/Sd2UnddPQfg
RikJpWVCn47vFNdgEhaBW1x3InC6K8MpJd/wqI3FeyoYeU6G89pRj5ZenxCF
kMgAWUe4pe8IJ6Z98ZPhrTGQCVCia5RX0XzhBHF5/jpExFLoqj2QSEKinZcc
P7wOmW6bSYv1hEJUysHwyzzCA5wew9vI8M9mMDNeyVA6eWlMhXJU8OqNMWs6
0MTEfr4wAZCKnWGj9Rjq31kT0zPSdB2jEXyYgmkSFILkcNopl1GGUhwtODSU
CvGggk83m/JqQSXmPDH/qtS31H6DFOiXrrk/NxAiCxT27K8Fuoa2gMBmIlmn
UbdCV3pwSNpkcZSJ90m8ha8furq1QslnBmBcxzm4Ai+alcAHmINdW5SbcZd2
tsLOyvFylboTTPUKbpHuU51mj7t1lygOw8xF3hYvOLK7a8d6IbJ2RhrJXC1p
2fd8wINpWIT9RZguE3ozKZwHLidOygay01MvCvT3QxuhUsXGHuG7A8Q+6siA
dniM4H31WSo4lam92gtjXwNqbZvBBlJN1OxOCUEYb8iTFg7eFuvcnHcFad5n
Kef3OQbazoI/mkJ5J7BM83f6qSl8cV/ou2j2i3S67N0AHPWqgo4gkMIL+2vS
iXGr4poqCBPAJHW9reluRtOAYvqbZQa+tontwHM3HAPYoK4BSFvZSUUjOKeK
mo9VdfejbDRj9PZ2NPE04k9kEh0QOYbQhNFuDNKRTFoAp/iwXuggWzQ7aUmD
JuVuSgv39yA+WGqYeQWqdLfuhrQEUxTBMNyzWLU0lcBw/Nlb+BAkJRzhzXFI
S8hYlT8AiVhHDlxi36+t1FCY88/Lr9TKJ/YAAn7t9fb4cnKGQjVM2SGtEkas
NdZMpgXd8svETjFwIdGps2Yg0wkcZ8bT4wkj4wdqZ4YxZ5HGkooUcqjvPn/M
cTGgONCh6TK7qtrA4JhWga5AwWo2wL4eY5cvw8frp2FPvhWdlMjojYwPYOO9
crsMdvOnkoP7d85hFkFrCJQirD2JTwZUJWZVKiZueRWK7/2JdwyS7nKeKERN
t1lWpkXqpA/CbS7M4KnpfHFIb01kmKKeMhXMKKBLbfCM1HI1NIAhosvt9tfS
4Kgho0kNlGGY14pYJYiNdRGsHGEVRwEcDk+UB0N49WgFQSYpzCrzUzIzk24F
yq6iwaz4AR9G0IO6CiiYEAQeuDLLHdy3NjyWiKRxFN9zrcM0HxFWtsbxxqJV
vzCGxS4WuWUEoUSqyhMcs8xdjHcK4/o25gzMhvSj+ZXcnVLURqCGsaNf5+Zf
BWa6+FHj5PFQ6mPZZ2d9SfCdJCnhfIiTDGwifKVHf9IX31jDq9TiAcck+bC7
6tg+JF9/P9eWp4KsbzjfVxjY1q7l7bqaRogW/kZyUy9RClmyKA3JmqFOtxmM
jU7az3JDtjIBzpbajNcGO4MX9dV6XMCvJjFIvHbgpyim2SOHuPE63d4Eqjno
RtDchCX5n5QsAIOqMmuJTvERIu27XqMtOmlJVIhM0iV6jaVBQEWPnsDfMfOw
MxToYHDt9wk2yUS2PoUETYnhKwNQ6tZGm8unoTZYCTYEnbNnu8WCRopy14zq
nDc6nRwAfuh/f6RyoN5X1QSLkEGOjzEFByhV8FlhEwq2cVSZEOtjRg8Oa7pp
xCHln4WhivBKSThhw2h3F9+spGzGICLnK/MEVUYYgTfVMyy0KKRjAR3z047x
u6zkfu7AH5CW+ceWZlZlKrMj7/QTMVb7/Yj2ETCKxb7iqJP6x4JbBNGZS+/H
vdasqk6QWRIfGrv5dUt1iTAoqoc5a0CfyIDJjfN14hEL+KrQLPH5HJo/2rgq
vus/myz+jq/50NsG+bYpO7wd2LyXYatrKHT+NZC9SAqPnIm2Y7HEtNgvSeh9
paa7G339fRA18930+5qaKwMb4s1znajiT2Hi+3UNb5DC8DQVeJyUcWK4Xa4m
/Bn/wCAghQAv8JoHJZK74GHLBOwOT6vw5QEsVStmBI8At0BEGRUsXfLtOA6t
qxWouHagNzfYqpUA3AQyibHi5a3nwk9bPzCY61zDgvLzi5zHLu9x5CgulMHn
fMA7bdT9iVpFYf6Zk51VJdEN2xYYkWtyrtWPLF+//wZYbCsVC7DULnsGPXcn
JbYg8fSD8iOFinhTh7dEBvh/7818HV3vaZ3WMkWEI66WSyKCbIODXktBdSOR
1kMUvqZpWgtwC+YDSH9+Pcwt8WFrFntZGvCdnZzw2c7uP6/s8wPMTxMPth6Y
gOtk5ByUmgLV+cDFpt+PiR4dovaTH4L3cjd7qEQWo5IGMid6lasDF7bupq/S
yIjRlEiZdtYEYhS+S8ibPhEXgosI2JkxRynj0VRiZSiKvScsTvhIsOygUcRh
VltiobJ30+i4YTmTP1+ru4pxJ5qg3KwwJl4To5JH5DJhrI1dOGgYGgndYhnb
WpmRXFetZQr/UUwPAUlQTIeoQLnSV3zlRgu2KZ+YVmgtdiIrmTnMjsaL0DV/
UJCtqyEavR5pnCTOyQQmjcq/MBla6Nu/9SrLhv5vVRzbsSYcFogNuDsBDLMW
Lhx4LqTbebgIXG2RdVHTp0YYiFo5flD2RXeVEGeqcVw4cRZJG6l57+Dkn3gv
YKURVYfWvwJe6MfwaIkoiI3kIr3QtzGnhENx0QZG+GUYGe5OnivO9Q0vsQlB
NDdpDRazRvqI7r3StVX7Ffkb0aXpKxZ4McMB+ai65wwDXwbFbR/fD/LJkv4x
jG6wrJ/6V9Lu3z4gL8aK3V27syjYlGRVg9qR5kXJrMzIU7XCFgNj17B6MZWv
myi1pSBD9wK2bvrmzaJmXoDN2SoQBx8RBMLNN/SOfJNtOvMvdqwhkbd7aMri
erZoHI7RfNY4X/vlC3RHMmQ/W9RaQmF4Zbfl8u8JSplhvnK2U07bkreRWnol
cI3wa9tX48Ji/K6n19DjEUx8U2dINRbF+fx3mbeZgDUjA3Br5x3qU2qh4jak
9mCcCFnCbcdhWgyqCz/l4qRiQI5dyDFMN4pryWdOLyffGFDDWork/Wf2u1Z6
vVfTUl6dZd5gYUysI1u4AddfZFSvJZKd2KrVpnkgaryItWe+GETbD9qL1lom
Fqf2GpZB0kYXpnYE3FZTfY4UUgOYp52oCfQM21O+k2AwTkQ7Y4TMv7tvfcS0
LTYLtYug3o6oYL0WpJj5OQtRwVV5/oLDhJkWD6Agjc/SRbjJuRPLPzyhULdb
xe1yoahonMQIYLKF6+5FGQq+sGqJdFmJ286Xv/LH8nQ/tMeirVRs+08RU713
XpWtqVk1ewUsPZMRB0ptLoaKbOvJTPfspHWBy+MVSllcuqYMAWMO8moEd+RM
v2MmwpaIhPMynRIx9/tP8VA4z4yD2TiW5I4uJ34YZzqD8dwTmFtaxqKwD5rI
W8nQmNgnCw3uAtqPiKjIonDfyAA2MkZQo3OtsWGy0WLh5m1Qsx8VBvdulzIv
/VxOtGzxQFPJDZgziRrSgEDF1Zx4EAwPjdqCxObOSKrnd8bavGn0/uJ9zXZP
1UCCb+z2d6P+ORugg4fjlJ66Mn4j9v7+poOcONpUBLtvfsLadPyg4FeYETEP
H3p/pza/6rJIedA+ccAyRgqeoE9ByHS3UiGZDehbpyM/QhMVAjg03FLPK4Pr
TY1oSxyo6ZF1/WF3Iv8OJdWP9jQOUi18aD6PfoPuaSFQHoul5TMMmCdw6zio
9vOGQUIZqyqxbIA7iFNaDVGndeallxVCbxFkRrapsmHfGMQelxg9cnI8Dk49
K5kFEZv8rs4R9rnJkipypJugkHh1qitpdLusFjBMlTH0ZeNQ1KA0A7jMcDOL
V+xS6GFafbQ8dSqYh3FJjWDA85f7jAwK3lcIgaTelRRuEfuQDauo98pRFxwN
6kyEXBN5444v31iovvR/O2Ie9PjUaMP4REUeHpj7GqkP+sXsJkSZrrKQ67/W
UV9KA7Uql301YpQlllF82qtMYDqUAAm7xKI25Mh0mziUswx/y9pSSrJt1Uqd
XDm3EbHgk/TzoGv8AAOdKImSEiwjYmcWW4VsvZihrczqZFs5bNe6RSqf/XCg
+nxbD89eueNovzgpVy9tmlvwwiRfrfAWKhXPedqE6zyYnoyg4oA0xgjmIUu5
woF6LjLmYg2NUmRHjM+PEmB/CQsserD4XWUj2jj/Pg7pr8HLqHhdN5v4iF6B
aTTXNQqn7to0XsNmKF5kdr5OKh/w867Iab3P0ZDj5WHQPUqwOS74jFnBqxv4
Sf6QEQJHKG468avZP0olv8cZPT3U78BP4l5v4E7MK3+vAhzMt+zK9RFFkq7k
BRG1pxlwDJdw9sk5Q4ClfKuPicVpC/nLZ1uzern+UtJB3uZrdyJAwyMcd0gM
L515lr5Bai0qXAXI/5As0ova8Kw8imktnCn77N7o/9sD1b49RTAU03XqUTnt
BonuVZOxzlWsrQZcfaoQ/QzMQOVAwXyzP9yNLOdQvp1ui2bwS/iM2I049Mjm
VXwz86tWs0O+wpSY0SfLdy3kQW/X5jdpyEC/v3ut8TTlWv89FB0lbSro7S/N
O71DyM5wHlClBE25zKX/JpXrVSfP8LK8Wl+CnL3WglLKoI7HZiKoeQHoHYIu
y+t5zF3kM/tJORf5CGPRr4/nKAoxfZWI7UBrAjWRKjIFBeB+4FkmqePsQrgn
BygGvrNkvvM5Q8+Q6h+cdns9/WlSfGp/FdhsgNEI2GiSkk1nNZl5r++PlD9B
xkKj4u96nuz5spIZLtTISSzaVbH1XsSwA3QUNCHEJKsTrCuL2t6AcKHth9YQ
Kw4OUQuivIjodW3L6jbJhBvA7AavK19pX7z7k0pbWENTyhOx3o3d1+pmrxfN
TgAGwaqwmC+Abyy1ExsadrbQcc/auhZ8ZwgtxNdbIG1JfTUD0J9ng/M4nKCp
pYElXF8rOzgGUaagqt2kk2uYhjb4JdYV/eM6r21/UwaLw1Kel47GbZ/IvJ0g
h1Yi5r2ifstPqgg7djkW6adUCMMEjkeT6WbLBr+gtAWCZms1GjucKwlNvbWE
ry/KMIXk+1y6174VOrp2oJqX1RGUDMerLmYoqSHcoDbmGAINqhMAXSl9DyMC
KCPudFvZ3tK14if/f/+T+Pv7Gmg7UKLNznuyAoCz5iyjnmoVt/tGxwP3EWvZ
3MYFnyI5aFL22GBfyzXaZZkCSCpbEgXxmtC6rJ3/Y2+X4YHG0qOqQFglF23+
e5SH+TyPB0s3JvsyfiryfV6Aj9UICL4eqJv3CgCQ/dV/TcWvdnqNVxDTnTif
Kz2Q4hISVSaSj5ThUXj5IRIpdIm0cQReoX2ojDlU73WCG+IRWatm2xoNqH2O
GDeRNncU8YEkUaVh0jhAaOo+F4Gnq3FQsb2u8qT+vz/1/Y+7X8fegdFIgojt
MCrqp+8pVq1yTfzhtt/u/vCjCtnutlrevAinyTNkECsSRi9xGZrpv8D2pWeC
s3CkBD2dATCQ1Ti1qCBxZEpNgX0ridZXv1WvFxYMSlou6b43uu7Gy0vG5ZCZ
CA5eOQf5ZUGuxFWoHissBcVyr3ix5zI5420FHf+/lTodkoFoSXAewpwd4qGQ
kXvY1k893SOLx9P5EARtj8XqA/EanKOACjuQZ9xRCrbAr8qZcMPa05I+HG4E
uf1mYCj3u/bO5tO7Gkw47LOaME6brGcDtv87CvsjSJUVGSW3pUlr7e6SUfjj
CG7+r01/m2KXpqBZVwbBBDtXavO+kuoCOst1UPLxtCmSAIuD3d17bD59Xown
IdfrH1+VazGoYSSVscOs6v6FJY3WIu6nl+6mLwld3M00GSANaTcjjVi3jszf
D1XGwh5Vm+LanPRia6ZzMJocNv9SXogagj9FCjW9ggmiqYnQe9idm6jfk4r1
jSAta+n627LSd7DpVXSlRl4GPGSPzkdbGWMWXS1Sa8fp1JPyDow/76arc+XH
CxKDWKgYemI5mWtlnSr/HMA7ckhyAETkCZTdKK8Y1ULETJOeh5c9g5YTVPSp
aPKiPsR53rvQRwnSSgMRQOvnAtCZY3K4sVsG/XbHvEOD1sz94Lkbob1ryjbX
OC3RlruOL/ORfjXmaGAp8UCJX/s6MUrtZGMH0pQfEK1ODecSeSPotM+aMG4G
I44C4Gz+TCCqGm2mKomW+bWpHfQWHIkhmiYbPCtJjLot5HAYBjqw1aCLzL+6
yFmvmuqQrjgMiVcrtsQiEsJvSAfDAadT3pGlUw8Iz+Ox06g0OQGHWKJQpctZ
hLIze0byOhYiWKSTRTSK23ZNeZRkdxo2suqmhj7NJNz7Ag6JWOwHwfg6LkS4
yq3iVXKgkaSK1ivr4GFd4AVROG+OdelErRN5TkooJxXwBzRsWg779so7LFYU
L5fGVOQFa0NaFhjFvUXasI2Tfx+eQ5NjpX/13VRy/lhXz4d93WldT9SPtvVh
u2HvX+DWwe5ERNIeneWg4R2iS5nf9BH9eO3OBHAJ9Gdfd1m3iDp93UNLlOIp
sEE97ATwfl3+7q/WnnVHhhGb51PJoyIuK0hPmGYdjahlNz860HP65HOT4rJD
dL85IjzkdRSmHoe4k/TrM1Oo3GuqaXanwmDCWDKKQt80BbpTSjH7ZzxFiO/q
YTj7E73gcRU7kMWd6ctBDkPZ8h+kgECWOg2UOhzr1kHbyv21GeBB10cYiOI6
2rWV5KlVuhZv/TToHQ43Ot5MFwFc84Zz0k6/zATFFu24I1zx1Q3X/TZoHGEi
8StrNmlC7g+AIT3Rrqw66BIg1xfpZhil08oxrFCFIe5fhGlHKYRUOy0AYOZD
qR/iSAMaEPETr/iywyN7A5XXeJr9gJNAoGCu8HBg/hsUIn7TW1KvLVa03vUe
T8dx72+7p+iekFrIIHKrl4HDf5JXbghd9DfTsCbY8rEQf5JWpYQdMqM78gL8
9PV8oZIojSEzWkv21XMbNDtrOBIecx1DdnPvVHrAg+vkjiTlZ/SaG+C8vSp5
vB4pNJ1m8Tx5ia302mwXvzOklewCU5OxRG00DuwA8XxFvobdEiS1weA4jqxL
I6uamQZd2iw04LPOPb42OCXsR2FWG1n8LfbqFuneZSkMd+08qTLuZ5IAChsN
hRpKXf82/KeAKRilJ4L+x0yvsbbayjFDyUVdsWKKYGwVKpmS6+8DxuEFOF31
9fVRDerN0N+ZXL/18kVQWNHtRRERqf3RhMRGCCga1T8p7E6w8wX23Hcbblml
vqkiPQ6v5cpevAmZjBx836vUcsb1qv79a8U2sR2cu2f3JaSw6ozJ74IiEu+y
jglyPtfKZB7HnB7Up0dDTdINbm22GXRN9qJTcbzySR1GHErH+bsLmFO8g2zV
0LqGth7EI/H3JJgwLrV/XtOsuFb+jWwMQfimHjLpYJu+0v7BUfLoCMNus+PJ
Kskt+q3yR6+FwexO6Hfxon7NS/fPYpvmuky9gxhRVeT7asyHpPR94hLuvi0M
ekJQRWGeZnTrQTKs6RNI4jLGdiPk18+91yMLB8eoXomeUgvD2KxtHG1+Gvip
1H8iXyNTrC45jyePyIWXXDz+2Uke0QjOzugnE8KEsA9DMJ/Rwzd0x9nsDz8J
SL2qpcIgVGn5wWIeN/Q4LJek+SzdURGPMge9f3kBCrR/U3yzM+/uZn6ndGyK
nOlKb6jxFVDjdUWVDZA65mRd1PSSuFqV4jcsQ/sz1oktrBMywAVeg/knJ/RY
lSZBuMxj1uRpT4Q9j0LA1RAsRPGR782X69P5702HCnbL3KLcFcslStEQOA8B
83eYSxvhvI7MgMM4ChuY0wj+SnCosbdVSRqc/gXMp2/8x5DW+ylfTZWZsOfX
7QKkBOE/VnjZsQn7Lp8JdkRqjjq8XVFhQoL6gXycJ1jMHjElRmfQ5mQw+fk1
KyQ0BC7XNd2tRA3wieiYFrWedvkQIDf61bhs1C7C0wUVgBiQcxtsFLgIyaJF
GLTJRK4TjZDZBWMwPH5kXqUfQ3SOqCj4uwnhScaRL6kEEV2/nZE42/5gE/9/
33i2BsUkRkbLE1c62bXWvG2xivsf4fpg/j2USq1+EPlaWF6N1ASoF5yoIF2s
2ig0LVOBZCDVxyxyy0Zu0MGIhnn91RE3IyTb8vmMBcNIy8xJdPUb/omhE34Z
mb30FVADPwbpwDzrMejimuMK/t9F/BIppS3FuR0ngEKrHbWLpJ6SIkmHOzak
D9igKhpCe+o+oNKzeBXoC5+nuSewaqE4q+MUkuvsctEv75PDR6AJR4wQmLrZ
kGwYJ7h/s4UZkugzubYCyRV5gwPRkrp+yyF5RCsxMJGi/f+iRGHRg5ht03GG
hgz0cxB0okmfwoKM3BRccRoxSzpKYXSPlXXGSLrb1i9kZZd7Jh6PRtnkAE3C
a6fPVEyTqqz7+Mm3JAwnZZiQj0TNy56hgeQL2aTWATsahcg+nW9dtoov6TWM
+tQMrbXQJKy9Co1saKdpzn8m0/6MYLFl5oNUeQcpyjcTNJ/PCh/Vd2sd/vFr
LDyVf/mz7zuHHYZgMvtc3l6HchOVW+pu4URcLcjR09eSZZJkPOHpydZ71r2x
YNdxq+nFlJ9ieBn5KtLX8jwf4OcNSIabxAHR5p7duIHWMm97aieDD+84wJk2
0HybMONIAzF+cy0ioTCXEf8BEf86EykDAynNTVzFUD7OZb2mOeSRMy+NVJrz
CoYLAeSOjXrnf2oXwq4oTVKDAqQyldZKwdGU4WwPCW41dD633lDtZHC7CXhA
qGlHD/MnmSNXF1jEoeAyg1iW1poUnUbDwOyW67AcZsiqHr0Qth3J7uwsKwA9
azWFUGga/rOrESoqbhNKUfbFtgZ8TDNMAJXIbCiun6pU5iuSVmBR5DLNhB6G
/xRnlKhDS8uNIBf2HHAkiCiBm1d1PbMHuhXug42iLgt6p8i7ZneKjvZcY1oM
oT4F7sfTFcgP3FUeWhLHmtNjdYWo9GQarHJ8ARyqws8J5yy/M/CrvcY5wUo4
Ue6hFd53GiQH3/350GxwH9PZuPEgTAhI92v5d6f4Fi4ex+TVW7dzH7MnVFBC
goq6F5kLc+Iintk9sV71B9qg2DF8kGNQzcj08AZpamyCbStwv/GavGK078m1
YQAP8v2QRd59F5POHjTsepZd/O4wQQmikRRiQ7toP20SWgInHDG8zte5tppD
uHwqtFI7orhovGdRrrJ5wiNeePDuI0XoQkoptUi0Y23lWeS6duGl2Zpj28gM
uyfBOuqtP53686CQj5p7RFrb9jkwhw91QOQhdBDRXrdu6+51+uBTaN0tJb3Q
lMKLQQ8z/NCGrwHHdbyUhwzcNoSkpf8QumcTaPnMJJSBKQowgFoVFcYIFo1e
dxuZJBf68pFvqen1HiWN/17trNcatOf9H2ABI0ohxqFbTSbscSSaY33ZUaeh
fs2bH/RoeUr9ZrlH5twls6/buHWN7SZcGIvz1fhmGQLDDw5/LnAmRm3KvbJ9
UTL181OO1giA/1nYKT6Iy+VYPrrApflJkRt+qcGEyQioUJYeEbeVEYeeLVfE
WiRM3C6X4+4oOPhJPHr7btaegriycRkm9wnAiypVNCL0YyciLzcjBJlfJ855
P+T8gYiErVA7VkGO7lD355iGRaO5Dbi4aKrejqWItBVjZ0BjIevNABoTUBZJ
ow7EQyZUH68cG27M2/fcKtGKM7fVMq5Ro083f3VW/ECkoXhhW4ai+mC2U9Wn
ME6pFO56eoNBii+IYcNYYhPor17nZI70ZxfcBFzQE+Z0/sHwzF7PsFWlC+qK
gPNoPPkF36jrqWUcW9XuzWxwV1kAaeBMmOhbAPS5F/ig4lltEogTDf6Iq/rI
rlgyhKd+1UDn/glfRkLyUPmZ3/+gkiztHe+W9trOqXx+rXA5NkIqKUQXwCiK
1qDizfOt/05am8QeM7p+M6jAOP3mIatTmQipWUwtHpZBo5rC3kKsB3FphGDD
hh3bVMaEtkGxFHeB7YtmMDlOFV2Yu+LUAg0c/1G/LaznAVVgnC0qIG0JfqLa
O/L/BCJItb7ConceE+oh1VvxWWUDtkTcp2RQZtH25A2S6gXpHAaip3unTNvF
WciGGl74Z7S6SX9nCt9XEgJiG6RhZqogQJl+4mgFWYxiFE+dTwf4mjw18MzA
uxsv5sKE5oBGbaa+wRzzbL0dtmpIzGLk2y5+HGYDm6BAPVF75oX7y1x3IPig
l+HXAwR3kNVLU0FKx0c905gjKmDK0/sd6gGCVH2W5HC5EVtTT5WQNNDZSras
F71dYAW81Utf5UQSLB5jiUFIo3KZnf+/AjDSDfwmpdssm2APK88HYP5b71tu
C8ywO1AWWsR5zU8jOHFSjlvDAP9Mzn15wGWVXlLLdSYk+WtKGcz7XTHjO+b1
nVbAZi415SJI0mQH5WEQccYOJ1Ni2SvRWEcNA78Dt0PiawWUrJDnLeCefSct
fPtsuVhaHqk1NYh8Gb9WD9T/5xtxM7O0YcF0i1feunCwMENgHjWox3Gktb5/
JF9mxNhiX3BkWQRXb6cU5H2bDknYSotNzU9vGUB7RfGvJTthjT1YcUOSkEKe
EB+Vq57cnJMLIpy+I1+i1PU0iPytBwmO9ClnpK5J6Y5pxCiAf7NPpVl4IKc/
Z+qCwc5Idg8CymDXMELR6DktrtUzvSr7zHkbsmBlGky8TwATdAbNsRshuP/i
RbyOgCIJzb7qKk6COvB4fX8ez98/oT2hWB5qDkLL7WrS+72QF1J70R8rExoa
ZNZQk9iyen2ZfFn15k9P7HaHMlasC8m8BAMZZmCcVAkZLoE3oMCcXl5zaZmh
Z0YmLZQYX8cTOSOFeSi63CY7kzt3BdkMJH2NRo8uPXJwJDoD6pfarjnDmYZW
A3qXq1sptCIo13JfdEQbfX9am9SQh8EMyUS5h2baaRD0dwfhHp/G6AsfG22K
TAfgi8msY6fSvenjOFVTFKD7gZb3pkfQF6OANom4/XWH07jAuhP0KyPghXI8
UWZFivV4xpaYMKhVmYUrzFmFHpx2/l3A4OisqivGUxxEFnxdvJre6ykgFMfZ
uwUaxoV6h7iL4PGrVQCtqtSmokx3vJK3+hplIqDjXGsC+muIwmhn4RsL6G4J
dEXFk9/h4x0aeCSRuvOjuGZKA7mw+eaeyDQthxdo9n2cSlxCrOIimP5gbSGW
hvQXSfhn6Kjwguv5H5Tbd5t/7E3SlgOOCIfkh4Gj/2GHWZ4BlOyCNCC6CMfM
qKUkvDWDDuWUku4yfRldJtxpjVAqB+v0bpVrWRZ/zUzVzCqijatjmrZU8fIi
hp+cdoCHXTp397tBf8uJuSMlsb6W5ZRdOHp7iPGf0uAR5xiP604F4cBf5/6n
OnTivOBqvQeSmlP6ozhPKCpGzCHnpjckFxH2FYGVpOQfq5IrOgPdfsrKKQ01
Kzwc7xfeiqd+bajvbn+C/vYzjHeFZSeScEpCL5oCV1IiLPPf5q4WyGjdLdsF
4XIt+cthP8dX+EPQ01oZXo11qqXN2VXn6Vr9CY98HHVSP7O49e4eNBL6tRRX
5uvxLrhs297bJQL4gNCFEztG2M0cq2Q5O2lEf7s29hw0gsFSZxBVd9cCKbbh
4TGblEI0LD6TDJyQ2ielWK34ysxJnfRSFMsHlGhf2aoOm/l97aTH5VKKNEQS
+1yvUmdHo3zmaKwKu+CrGJAn+CAtIQ8me1AaThLb4YfsXiddVJWhoFTwoMkY
7A3KXsnos3iEfnk++aqJcccQ7b5oGkj7XHEvPzceJwEljnOOoe/w/LdTXsi6
qb/DehJCFJMOGs96QHpp/aN0iPPDmfwewbT6UZPxRGB7F5ZTzCXhJP5C0/Fy
JjXUun1h+V9pOukDEFv6mx90ojmiA575LHBeMipEfHtI4nO4uknJ9hRw1bwu
zpjT13oM6ynNGOi1+PbsWcXWGReajofQ6jeD1q4cdCrtlGB02a0fnBdOI/iI
U3SMtqz2sx9zGzUtU+cIJEdX8/jQOMm0iLt9AXJFFwPM3S8XI3Gk2ovXEERE
ozFrPyo/lkN8l/EkaI7aFfJzym8JH2YwEKc27oIJY1GPlvNPjz5LeEcTAQ3O
kpH807cH6vcZsj3O6BfmS/XkpTvEpvMY0UQ87tYwGhGkQop+Oj1qoiXbL9ee
FqZEz4L3/OUe7vN55rg4efUGfMGxEhQWvOig1dwcMMuG4qYYjjYQg/i9Khjg
2Me8AJhMDZzdCoVshaUeYewq7LS+Dioe7woK3ZuzE+f9G3CpjH5B/pHeP4/a
KB3PLpGwiBqYyFXrjBW/j9zaFYyaZOAYReVu/USp9JO5bGQyM6nYTyunroy0
jeaNFrOkf2wbH7o254tUACUSTBHbyLr7bBWdPgagE71sYFZYvn9hEJON5xjg
hOw9dIGW6ngCpUf4C96ITq6xa3kbIxYJ4Od9p0gNPbdXz4H1ZjCfTIN3IIFi
IPk929fA7pZH1cYPF4o/1a0eWmO5oEXBGLBWjIBErnRhFidrJgUNHeLYkKQ2
cTNfqBYrqy/RlfZLwAUOkSYtnbyYcp07I4tmteKBxFG71LR0NW8Zl1ZaTcKh
yZOuGbY1BdEUNBK11vssr4Dcx+JBgipsEM1hJA0lw1k/TG1a9Udj+efIHoLh
30YxtM+Xy98DUfFVc02ljgo2wiotSCmDjiVynamtmk3GvV85xktPwwQcyJ6P
GOweu+gfxSvJllFJ2DtYh8oiRst9MjtXFPfaiETpGPlI64ewqvLZjxyD1zS/
Z69JEUn1vk9pkbAQVYUZsO0Mbxtj4BsD7bbu/c4N2XSZtmHWCbnT5qiwVsoK
ooD/JCCwLh1LAtodj2UwDqP/QFoXXHQeZj3K+VY7i3gE1ctz3AgBppcJutcM
+yZDpDm/ft+C92+yUbFdFk+vZi3YTlCNwGO5U7I0tVcGh0bmiyEVfj+GkUyS
SZL4eOChzRgYUEDHLO5tXN3dBSLW02c/eO3/CPyyaY9dbrgBFERWdDP995Dn
EUTzc/YEAeGJnAbAVklcBz2Jw8+2LmMa5IGS8WlaPy4zLL42bz5qleJkfh/L
91LKaY+RtnsxjK3qCaIrngH75vMMdy3bZrXVXCWaWeY2S3Pu0ipZg7GzWthP
mchvO1iJNF4CMPnnaP9OWfRy7oO7+8uZ/QvG3svZiLc5uwkWKMPzU6R2nBl3
ikmbo9RoEdlB5BTPNAV0nKWJSOcwlbkD2/0lUSzKSxr3ER5CM+wsWXYh8Xcb
z+t5q4eS2pD7N89jRvbLru4F63caSVC/3izXi80+vrwx5nSqofp9MXdRnYAQ
kHtN0JlIpz9D7Y5HprZ4sqH59WlT14F5BnOF5LQP6fsGc/dJKieVkn9/Xj8z
rutI2vVOiABZT4bPa99/RFEu+QfmxQ9uWqo95InNHRpPj+nRjDlOxTFEWFKH
NvLKUXw0frSsICtpTik2nob50o2feRU7G930Cv2XjCmcPHD72xMYaIYqYyP+
xbpFMYPNRp8mPfuvt09XpHUdBh4vzX9GmrySERvECG3DEOYSS1bl9APUn6Ae
WlFmS27evDTVcEJMzEkF5AcG9r+byZSipkhF2U0q98gkiisPi3MQ6+7FnJWr
2sLUPPbQ+SEl7VFB+41vwIUitezEfB7DgTfIEF7+NXy/72+L0GMN9zP4pV41
+9BYWZBLu1b7cFm9oVEgOX+K8uifmBkupd97aGKd0vKc8IMkCvGDPzYMJfyP
A8dsghQA71tOxSZ5sZ9Q9IY4/W7m9i9JMj2oVrz1n4gGYCracOyiZSdtAURZ
gB7v7KFXrrwshLcrjm0fw2thJPO5Jsu6m4RCagir4xwDHerxNQrxntGZtBHT
35bRMtXm6VnwueTxKTaYWch6DJBbIa8mSNvX3ZB7mY7+I39FMGr5cu2VRRDd
njAhRT3MTGR1VRDF1iIbkzqkjq4RrC6u4ZoP0fU3BTCc0rruXg03UlHZpONa
jmyQpsMJ6Vrh/oi2ZROCdl/3GO4EEAMsQsO5cgLd9n+Yz8b6lFK1ZimGeAgP
Gv1qlphLWvsfbvu3NF/RqA/wsSvf/E/XWEF8jDU9+rXtAKuOiTNEHV4gjBgM
ahK3Yfaje4ou4wlhLsgz3OsnmhGLg1lIUJYdRAotZbyNq3x+mvOc1Wb4Z3jO
Xf8gu/PfLBwG8HJ3Lkcsz1EYKRZH77ZojnmAOcJrycyGXh1dpCj034dZgQRg
NBrz/pH4t45mUe6WoNk/3Y4OC5RrdAC+JuliMFpd4aGPDcisz8a+biaf2bwK
2aBgakPm+S+ttNcW/ciGJmk86P7mapWwgt3Bg+kGNB7v7xL/DAleUQBfqasu
43Gtp8TRmbD5MKLuFBA9oyymQO3pzOgnbDZibV+pyGsCXppSgSO11fURHSi1
HZCpHJpn3sC5ugCd1TW5SO8sIsApcXzuw1F2H3qfA9bA7QoBZFd2Ju8UM3Ig
44IT+MGZlng6KqJwUSZFCRPvBI6Hamo/QAddidWMOMPag59QvMYa9jAne2oh
TtERVizElArozEwJtthlogLq85uxkSLEMQpUhPgW0IefkhJVDx5F6swPnAYT
cIkxJQve/uXzoUm1iBv1VNmcXQ069EfJj194Q3ND5LxUWxVtdQ9zN9zG8fa0
NkIroxODpE3cgtaMI85z7j8ume+jYCl5sUn8VH/V+L0vJPwJK6P3xYu2Ux6v
ceSg5eRwc/lo3mHufCv9seFiBErVBH8ay22fKm27MOYn4WINBu9FEqjZU6PG
wde25XFiVNsHXY8Xf+VagYMAJ/YWwHB3sczRGHtNzvoKsfjolNw93ezX2DGV
ZO6t33T99GEV+5yU3kCZrU+h9f4+Q3/XXUaOn3w/uTk9Fjwjzh/psKXOhRYw
34fjMn9BDDSUbxD+BjCwyKx0iJUW3zbREznZVpuL2nZpqkJR9u6Fpd4CVgSa
YTymoREUJ7rXXBhFrS8SIdC/CPmdawO0ML4KbnCjHCFr+i7Bt5VmFmz/txa5
CWR886ndZrtrEjBPPFu1t032lmku7JmuhpIb3hVJTP6Y0g50J/aV9DavlVGy
mRtC3BicvgbdHZErnxcqWPdwQmVi9zWnNMAUkHbN2+ZmpABYs9taPeIzdD45
Hsj/yinggtkjXKdqmpjaBS04jbKyycK5uQXLT8HtU0Cw/2oMoxghYCdo5N/T
EMHBNnjTxPTKT6WONWMSC+84q+Cca2NnFNI2gsOpyJ/0cluRP0LeDFDE20JN
MYmzQYzx6VfAN6xJwmT369H2+hf5pDBUaarZ4S2jwVOOIcOo6R2RS3kF2x+4
4d+HjJquRmQoBynvic6t/rH72qM/C36OuXQKk6ughiMR6fPUBBKWAfpp/RGE
WdVKPpWOtKC/yw0ykJ+xniz2QtH3V9UHRCo8y0dwgo0mZbzeNqW9piy7hEZm
HJmt8FO95FLS6ywsdecpgY+tor1f1rjvDFUOkj70vo/WD8AhRE7IqeZeB1VK
AuK4H6zCsfW5/pXm1OnVlDT2X7VxsTBvK4HOn/ORzMZ9Tky/3GwO2svMoe5B
nhPGqUQ3M+dzKOSUyaxTcDu7RtfGZ6iQYwzkDgQ+b2jKRpy9gSNWoFnkgP4B
7tI6tBBNo8iFl0Kp71HiYNc3EgnI1tmXQwRQKIKbtBkiT4Rdd5Bfy+fc5osF
SqMN4eDU1IBBJdNcJRArx3Izjd6esQmHYTZjjTIPzs2uo+e0Jms/qKtFzNvw
zdJ0KzBuXIs68yM9+SBT92Tyo8+1/qa1y88KM4uzHNrriozpWQN0TBkhhZLo
11bj6Hl9V9EdAZ4g0ET3cxoZ8TboRnLNSmcEL+LtE775L/jaJe5IigLcSnJX
vD0yPF4hEDw3+LMk7wvs44/FOExv6BdbC+JXD/7OBVUZdJ7JUJgHt8zbS6cI
Pam8xjLqUTTRywRmNPKRsmSYxd8dWo2zsDOKUXusqpoJmSCcPlligG227GIN
Lc0FI41xrsl1KFvOS/PQYPJxXXhhaaqqSHEmHBHH074A6tB2871ZS2WaDQJ4
5EpB6DajnQRrmuPr+7wRiOLvdg2gAX71Cezz0v0qEuduDYFdUB4gmMhE4laB
OQI7SCmMDtFJ3uOBNmbK66IGi5bFVEWObPJkXPNS1ishIQfpAVmhPeJY4Vow
vrYXGUl6RLrpUrRQyJ9qIy/onVlqCfF9BRZ3RdHZZ1utOl6wuY2ZYaw2b5Az
+Ws1CtkvlFGNvu645X8Oen6kjgpnLaw9g1ygHIbXa6ZGayuun1C8xhTsgFNS
F32AEaKseyjTu+VXaHj0e9ltt8gPkpP+oP/dQicEzXM4eJjwQsxsszUZkB1a
JaHjdneTydjPoOqWuqi8dDHiieLLknKRP4WT1oX63DIAAT2j5G2WMxOIuBH0
F4dtBG2X8StPfp8Hfv93bVSvylvRkNAGvXeTiJYG+aGY65HB9NcUOugvuTBa
y1w8YyOXwM1Xu6LDgLl43/NEJMlDSzuvGIvnhPj3wLr96wlcQ4wLwJDlySR1
jGq9jXqsnJlsHvXxUTDrvLeE1YkkGw/WhgY/CTy7gSELQXeybBT9cxONoIza
S/pwV1fmmm5elEEteFK5I3zaL/6P/WatrffXijUNuR/IGuJpdsZFmhkscAj8
BC+dYYtjCm2W1WFmxzl2UaFpP7FLn0OBNj+EyFLXB7gHaJ2S0P6f803Np/ez
qZDph+dGkPxROusnewQBxbPQDFE8vzGMvW/Uez/4zb67EdcUspfWvPXYgbEi
dQWCbFOLuD/9GJsDxfpJpN49UoTlJkxXYc5m15elS05rkfEmQp/5PZazkulj
FpcENN6IOGi95pNbqdngOmYk9+IFSFOfEO1eMtaJvroyQ1HouvFhrEMIbjhJ
MMoYiAA2M88LbU51y6kU3c7jzj1ffD9cNRoUJwLoPM7kMv6iC7gfL9Jun9Tj
dHCpaR/C+TZmhsniY7UyUWzSCCIBZyhdwtjmDTIBW7iXPduKKm5uHsou5kPK
b1GpXoyFkxf7app7hieCYJEeaGPRe/bJxBp6foZFACOb9NJw66mJSUSHo1/s
zxIV6ZeCE2JAkYq3RAsmd3jdJ3TCnWMny2x9zF//cPVnq5Dsb80rUIbcXf3F
HiwLzMefniHiWFVcnJ2F9Q5Nh7cplVaROupJ5GRnukbkNN76IGTNLp14vdft
MNDogAuihEno64ea65Vys0f8fqkZtrfPjVNS2gPRDZ+KjUFrgesimXVEkYGF
2B37LRIwJRwRslUyFh6Fro6IabtLaCAmdKgUW98irC2PMhrPZ/B6P9x0KxXa
0RXr9AjTdiEHQoCqGSBAiZqMVc8gERp8biRSkk1dHdpRC7br4dndeqEDC94n
C59USjGSKecrFTMdGfNMhU27P445I/iT1rMEDRQDQ0dF/2pfakaNM0cZU8z0
hrZ18w5lnSauoFOdxBz+gs5bFyMP7Om9vyvIw8AIfG/AktDliH1w5VYsiD4i
akEftX/V2e/DIIUig1xp+17mCiaWxpJnXByhWAr1hqoTxa9af7zz2NMXQrIM
Q32b6Z2eZziHjoUkZEujm/I7PPAKfRvE4QXmB6W8fNarkff3uTrQUUnY4eKU
Uu0oDZCnh4TJKfyUzP6It6zeeTXbFyb581uWLko7HsDBVDkeLg04LFS8F54u
pt516RO2QYZRXl3Sy0hIB2wBZx/32P8UGxDjwIO2iPAnryRXU8peIZPnKIVr
vBSoWidYbZF9ivozqcH9zw3gAJDKPYXLf91hketJn8tK0rI3GBTxGw+vCtcA
QEWBHSG5rIm5bDtogvyhKYI+CnzJ7URvLC46H2nlExcrscdHE2L7/QIJ5sZ9
sgNyBN/B3UR4DUCUmHyMy7/uEWI6uQ24XYv2KeR6MnwGmkArAbRngbLxd6ej
9dsEVVTJP6nN4T1JSVaaU191nfXHxZiFJGVSmD8I5aZ8CmuMI8y0rW0DKepK
qNKdzqQ6HXo41dvwD90Q4HCfZs6Jb3dU0PqK/LooS4uliRSMTnkGIL6jh5zZ
hzg63PY9nuVHkEuicz4Kg62KkKPS8QsGHp5Ksnef+De8bpjDxenYjXbEkBOX
VI9kY30qlcvfDViidnhxOwarfMQ0REVtGHVSkOPpeknSH+J9JgBdpEzjmroe
jOopgkLEicEx+EzaEQTVwLWONW0fwCxQRollD79Q4z1bvcZjF8xJX6TJnKD0
fTEjJEjdxlkYQz4moba5a48fRsjcvjSsw++9Tc40t/JwXaoLBOAJ78ObAzaD
Uu91QExjYnj7BHTDRf1yAzowBy77QjlCp+k1EC5cEob0MAxUAbMQhXAs3hA2
HzgvUxM0tgHhsfBzXhiblth8KhXMwKtwjxpvR7LjuVmnRACbm8e4mU3ZfJMD
Q+JF86xQ4/+eVuQ0elOlvRwG2MhKo2oCpWd2atCrsow6Bua7d/ral2iBckwx
ZpttjyswtEEIbYj6ZGRgO2tHmT8RNrlEqfYkFNIlxQItg8LCNhUCZn2/Re9c
aVckF3iyPFerWjdUBAVg3gHklIHQ1xc1C4Nb+XZNwpTKrXn2UW8FnHIZRuR1
WH4Kinsw2Zflef56bR3KqQ1Qm/Bp8Qs882VpYDwsFMPegJnepcjzZG+r4PEx
st90T2RZuvNY+7Ag8mriqpCBJViMSVOAE+Ux69w9GYhgepa/sXW6MPmV6tyf
Ejam1t/z1kq63JWmSatwMtn8ZtikyhtLUpV7sHwEvW3Lmprzi3ez31NK2cy7
IzOFYlEEnNQYenV4S3EVxvlyzOcIYagU/6DMBudD94K1yCJv2BNKTIcnhEOd
VgmYzM5eDMNPi1KCoJMjEU7J57W2CqjjeObDG/raCsKJxAZ806leN6uW8Lvd
02KKwDLLOJt7ITrgrH0AywPFbwIkxjL6J8fGpSAK79JcImY4yiYasTUyZnVh
nvditn0abDxWVodqHqkjBLxkwC3GT1izNLtry8ivHMbkVzMlaMbkcPsf0sKv
ocKgSI5jWRlTPI1DDAUoqiIsxhoTIO7yCjOgtRbnMfnAH9XquVMo9li53/cm
RqTiX+10m4y3rBKf5nfVZZB7gxs1DG0VitICsPgXsz9uQZ5mCEq2iFm1J+m0
eyxFjuFCISKQubhbHBTIeeWz3+ky9bXaKQ7YTMLdYufkcsy00AGpougw9tDw
xDxQzk1k7y/RDftDboxDU8JCHjY9wr06ssFYz1fWyWm/HcXHFz6ybaqO5rfm
XS7C+7sv6oBvyyIomaCZ0IEfz7CHBcnm87X2S7H18FRlHq2dFUqRQZtrT/RK
7V0EWaVVkbn7MjAwjDIjzFuaOYimgX0F06Lkaj1QEvDJtnPVyIEwbEJ9UDIm
FUSVa0JiJzLHSG0N5TR1GSurHe4vjFhXhBTe62rx6PvS061WpMimExLiLvlT
HtcoIXo6xuXVH91ph1AwEck9IqnPSu/ewYvHNfcr1pBld1xFBrWVNfvl+HbR
G7HPOOnXOSMqCSG9xpunASwMKvEhVbuw1aWREyzpW4atzzr2a+cMSkLirAgi
2+0AuBRtKGJe258735SxUoCMq4F6opxePJkYr/WdnX5SvSeH8ZMCnhYPnswN
v4GpJMKEW7pyHz+2QgEGI97up8NBYL+IkvpK0Ouw7bHsagnWZwl2NdRFytq9
289Ai6ZSW8HVuGcvHa6rmAL5IKlfVpmpShBPbz85zoAJcpSpd/hqEbLohzo2
54yEltRHHwZkDhIO8DwHXfQ/7PNUTuxMTOtipaM9M/O20pALrRD6BTxe3QeW
Y+ZLfICeqUcaJ6/g8jZmGxkFlP3DF7L9WXbMGDDSCHhWGJKGw/ovwHmB2BSg
LajoMbofPAIWq606F+ytLotrXQHhr7L0As0tTheGZFDCETuCnCFsb0hPZ7y0
MV5utH7YSJV2IuFtD35CxyaTyTpNfUsmfnSWjxL+8zmuqiN5FqCdl2x2mh3P
TY2pC3ce+tzxJpDRiyaVQg3NG+7aSvTFLRc6txr+/3FZgi8e8UIpgNlppq8c
L+cE3V8yx+d+x3vGsvRsKn9weHarEpS2Kes85wKlk2H7cFHKiy7ZE2vCjdYW
kyVyZibESz/ELs5oQgVe4ymL2pvZdWLSfOzUvR19sstfsJeZUbb3NMOT9pks
hmby6mJO8NzbNfTd6nT71d3wcvFYCs8kx009p8MZSEAnsLdMs2PZjO2JwlXx
2f618H0Ij97uQ4Ju6FIpNmU2zJymecoeHQL31qDs3/R5yf3lJrHSbQvKOdzT
MGWINdKnzXslYOd5rvJn768FtDm0q7gHtJ5xynhh8ogtjY3XqwTAfHvxfW7J
z+wEi5BWd0kzEhFP6ogY1Gzj/SJmpMwuDP+JoRz+SekPB6AHbfz7Tuaf2LZr
SQiC0QZxqYqkVWWYta+wbydw16gbjEmEeHh/be1b2rWvFFIfD5cxnqd0AfPK
tRkQ8jkA/obTGl+RR0llrIg6+WlnuTqEh4e+IY0nJvw7ObLuIsu6y6nmYZye
Tjf9l5fefSZwJCf5bh9wr/J6TLqTrz8HgfFs9jr1rVC6RuZphplh7u/yn2Zu
/JbJxeNwCZ4mD/vMe46QHt0OEBdxdMUWXVbC7P3+Pu6xLxu+dTEeGFgztkWM
KyqfYRTEm20di3SRQJz+qpfESqIgIuDTyr/CZkL1hU6IfPtoFWPoG/AhJG/m
6aLZhLHidrXSkGgv4sdR54t1gSW+xF1cHQ9a0HePPqsxD58WOm0KpsRd+AAr
5Oy8Xndu9BFjmmujQA0+DJDkYQ2TDkleZmJ85O4iq+dQD6AOTeZPrZ2jPsaJ
A+z5ihucSW7KejaSew4J3R3LTDTgaSA+ICqkUsEa/3tZJ3s8JUEDlji4LMMt
oLXeOnH4hJUqHsZ+KMWcrVZLHvKmdAv4uu9SSxcj/nkZuTwz7BRX9SldjAGZ
2LyLE95QvF5C5Dz8Ai+1Wc31vpJZh7WvPeYwDYah2rjKmydSmb0mfg3pleOo
EnjKlzVP8Mw3wvQVLi5YgAnq6vZa2E0NoLPSYvPoAqHxB9WrL3RAK7ipRJN4
rf8WCuZfftXVJrfS/Eg8ntd8IQdtD5nxuWiyvyJPNtQGC9yBjW4G8HVaSHeS
9W0udFq+LowyTok3gC12nkmhj5rvqX6HV4q7n8tyKHmbR3Em6aa1QgrD1CIg
/CYyEmmpUz4pLWWtpCwZ4yvYPD9d9pQReJFxDLv3WHERFPQABfTSv+KDnSuR
9mlQIvkcC5b8f5eDuCZgzd+98z4v1A7LwEiNqH8zBNcxZe3bgJXR5pZViogm
WV9VHKrmBJrwNkiQ0DEBPYf7SDtLTMbz0e1ZY0UmPAGiuw6Vv6hya7vBuc8i
lAmCYpDIqVsnBmC7Sy/EycncE9cJv4yee6vQ95SVilk17YsiJBNcBmsYNxdk
fA50I8qr3L6/xeP4BRagwHq3j9XID0rRafs9HwiBP9IJQFSnxtPRwYYgh7nx
aepmmAGkoCnxFMkyTscxyg2IDB+duH4rfzE2LGR0vTNFrSSgPl0PWWJ8tiXt
L5g3/5MEq1qSQGD+4aNGP5lN0PJdyo7xWvoPdgzm606yHMvFL7Kj9vMYHes6
vW0XFMTVrqLCb5p40upvuYUYQXZir69chmnlR2O2+VwgA9SoITLgjxTx9TiH
cEkMXTrdLSUHTj9ToibI/u/XrvX01sgSOGQh+yvMvC4rlxvIV5s00eqrDRa+
8LN++JQzUhbVubFDUOMGc+xNsRhupaNRsN5kQXNeL7A2NJv0yP/TNdXuDXzp
kVALxiqzRQWQCro0EJDSq/bH8h95VwT5sVJn8KHHlhGQkwGmpBcMc0N6uP5n
vn7OV/FpT10bjzV08RZ0mHwmSawB8Z8YfF1+lMKB9aVCHupcXltnOxba8Vqv
9r1EgPgsS22akkLk0EK5286XcuX7cS3Wfvd60T9/TgqmWWtZ13+QM3mdtB34
0rt7d/F95suDaHT7VQjTBkKMMH2ok7vD0Hni1WI8Jdegmu+htg0l+CGbsEmu
RNraqSWZqhDlOa1UljtH9E964bfUye5YX3opSefu4pRCbAj0N0Zl1PyW5mjy
nA75QfubFsh5YOuYyvxvmxT0ARw7T6ZdL3H/xayMEGoI4+6isH5dEg+Iuj+s
tSC1+R+XzGrbmZ9HPgOpOucCKcLEmPBVUQVefQYaB7Of+LkvXdI+bd/kHpcU
MRgx1oppn5VBKj7O43z8d1mMt2eOA8CJh4jrw0a3/fffL1sv6fDSDUWUx/wx
J8Y/9pAMsEPZRAwOkb7fPWHEho4HUMzdl1NOzOVslRgOaTQN1UWU+DCY23VR
Xq7WtHr632zIRgFBaoIXLU41r00gGn63sBTCjKizPBQ9WJwTJBW/LYgu6ChD
ed90YzPlB474hYe+MbxTk+W718PRf2cF3/F/ie56PaDPUydksvqkPQIxq1nJ
+EJ7pXCgfQwtvc+vsY8fX7bDGDPsQoZ7DW0htW4+1jc8h/Hc3TpYjxXt6N5B
5/7HnH5D0RPgsf2HU7se7Dq+mZyGNXqiw++6tG34zYOQtGEFDIVH+2KGE1v5
JTD24mJcvf+PtkgTMV/5PcHKQeWBmwWYBbrKzQpSKD65ZGZeTmfqXX7lfnE0
QClrgadJWA6rIbCp2l1424EO6qAF0bUO5IpsdNlRjHVsGUIg8NaFKlZ2EpSF
WktNBd1P7QJ3/wyq25SZegY3KIoYeqliuJC9prBJGByFzjRWnMa4kh4RGhMI
mFkYO2CXM52ZfvSbp2JAFSqTPEFryMvQy1T5zSwseS/KAEqyl3q+MtA6xrd/
GTzvWyaga06UnqtjOMjydqZb5bpROKStCRLIo8mez+TOOlrWVEHvzG2Nliif
BbwKXTGkEDxiE5YCl3QV4BzXcjGETy4qkuz2EI+MMN0EKr9cvc/cQ0iKOiB0
AAQg0w4vOUCHnuFjgd9MQZgyK4lauHKWp+3b9C59H2SmFJjL2o8Hqr1NTOy3
SoAI0mXHQRHS0/Up9pIJmpAGt2NGwPmhhlhvw3cVv3hhf6IIhyIfXet9Vn11
P5/BrTbsevg9uEZgNFSQhY/QCSYoTzSZsttx86Tk9CaxIETsR3181nIdRysi
DUr7yGTANLridhogqgrZ1YsdQR9295cdEgfqMhXNe8asnizkdbkZ3H6iH7EG
v2RwRBZhgDyNqYLA7WM8f0q5uGGmMyTzS3wawhzzhVGawfprOYZxRcoUFkG3
MHZpBj0Y1ro80mn9ala/nWK15dL3ISv1jTUYOGURPJHJWwjBBsPh+nmnjcnH
yWQ7G3rcAUnF4cNiTf2e9haOhEkD2Uin166ZIBz/3SI6+2bdyt6gPToDI4jz
0CF26K0wS+Whns/4ApWK41tU9uPEVpvp7OiBEnNU5phpPPLIU1gpOosd1hUH
6+CCOM1iVWXQnF+lmHImMIDpyQLHljSvUaIEMO+Es7Wd5YUjDa8/mN1Gu96l
gR04qw52zd/x3zM1A99ohELHiWNTaVjI8h+DwdJnugfO4Yc+xYMOFbqVjNoE
sRiZWUE6ICZrsS2a7Pw3gV48UknxVSW89r1+/hZE7ZqH6iAdxYq5N2RloYS/
qcKG8ARGyTANRT3Ybu6iW+O50M8AhhVP0TvVCRwcVlBGUkGzOZP61hZ3+QBE
4oIvKYDcKps62OjIV3fuEiPXJ/Nc6PhXfpO+1PUjdTP+SrlYpU0iTy0CUHrr
1VB8C3wzufgsc7b4BJ1onipu9q+rhqBhjMF+4R7n7QkWoxCec0VaIewtOUfX
36ZeSoXM61rOh3MB+j1o6ZgEVs1YEKOYx+GFMZf5HaXR3htZoBfarN8gMByj
opTDXgKexV0np0Aa68fQ8DWTubZnUoB3RZ9UKCueo8rubj/8SqPlINt/DVF7
bbH466rMr9ggeEJnEW2xh12yw1eAtNZlgf1THpEXpqqMJBtgHbu58hEaKRFD
fyvoVa+loYP2GrdWzMdXyVCbj22OEnRA+Vcqrh1h2Q8Q6kTueYMETl5J3mAP
3vnTZbX2f/FcbANLMfaE5btPBfyjudlBLrSpp25HGKXCM2WhAFbSb2iiryiC
YqRiyqZF+zU7XieiUkAx3fSGpHRlKLVVTShSc5TsyC+zuCdL2WzgVv3fpWOG
PwTkR/3La59IFIzTVHRSjradg4FBVBE6iYBkpDTig6OKrwyuYxMbvwFF6Pb3
BPOHkmIRyV4/tYy9YdriPek2Skbb0uKL9G96lWuT1fLg3gTK1kSD00ZqJAnf
4TIpHffRwz4CMY9d7iZ7uLOY2ve5B4zdcVmlMTSZ5sVT/oFmYVvvvAPTo8u4
RWqfN2WkB76JKz+Hx2rr+O8gdSkAUC/CACyY8DPUjscuND4gkvYctPMxhmtj
83MlVrHTSYVkyJ9fmRrEcgh69pjl0wqYTIPGuK3h7pZy1qAAz4fXWdM38UZ7
ZstAjP3OZnjLo7A7xzQ3iJd3nN+pQ/mLP1Oh4Bi7YsUhPOfC8PXs+iribz5P
3+cgXDiyKalxxCWIIx+NhcJmj+54x5HNFXIwbAEhE5Vmg1GeX30caqCS8eEN
wRr5GW31o0hkI96FDDoZAIPEygRS8fVJnNttrDF3gd3TfcXBw4DkzXzax8/7
KCEgm1wDeaySP+urbd6XUH3BFs0MckBcJYMl1+GmAA9xh/SwsNn14rxR/Qmr
LWRPDdf2bMAqkF04YotnanRSDD1PrCrAIzgPI0hT8ssAMA5mYz1ZaTCJmn0G
YkAB7Gp+q7jd40t5StsG4shKF2Otgk8WOuwlR74VW0YTupBGQJsO3dhD065e
qOoN2X/p3Hjvs/YulrGmyGhqENh0ox35Hm7mianRT/AZgolM6nWqNKJ/Lq4o
7KjywUqNSq9yr8FQs1oaaxdd+uwZshoueucoh72Nv3vF2k1mWOhBIAMrn0o8
JQhictSqqkFjJVPOqsgz19y5zbIkg+PHgcXvYrd1CZlAW8w9721eHyHE/yTG
EYxOuGx01fEYbnEM3CrdDDqROJwik282KmX2O1V3RxaRHGz+szVWT7qVr6u6
Z16lWeVoDgUATRlragnjVYfMC4ODsFS5BrKpbr9wk1LPmfpybGz9oHgJHLu3
Lsnt9n47Fg0CtcD0ysiYOAYANLuTl1ewnBxce5oPg09rNT/xSAO/wd3tIDM9
Epkveb5CMST2tGqHV7VwPYMi/NRAh/Wxx4Fl0M9e54OCNRz8RKy+dIsVl18D
A1gBwV3gMMBKh96mtnJYzKdRsPDofZIbjiCxvmg9oFHi2/3O5KT8IJ2dQjqH
0f5dehdfV6ZA5Jp4TP5LmBzbwIEN2JFv5wXRsWrVf6t5S8JjEkxVMOH9hnFq
rwA2JLiJbvOaGmFheiNb574C+ILYRbtjHncDl1LBUnsv61o2jz5SNuky/Jky
waGFXbnVX3OmYI5gFkPioD3n3mnDNPUGTsfLmejQc24RhT9O/nQuBix+3gF6
ukMlM8pVJ5Yo4aBuEDKHUiiGV2mUNwidsai7zwAGsVGF03UTqGg2Au2QG48B
+/9O5JLKXrSizAFnbWNK3yE2O8qQuZB+OnVkSpUg9EBeB8B8mbr3aECpOJpd
BmWtwy5xT2+7A8Yah8QEFZIEitE+XwYqu9PsdyW1DLid1HJdGnlFOVXWP+hZ
k0RnZcwK2QG+etY77hCXV+0bGzCKMNKooiddGz2hTvAwjuVfFyGqoZc/GiID
pedK6cvn5sKh1XMOyr6MiAKunKFHCigfHo1GAiQvi+eZCoTzStsVoNeFUdNA
o/iVP67+AoqrDakRb+X7FhwHLkgMXnfcpYTsJZJlR7LjAOgt+Y21I7lWhNMo
EHHWc6In8Pe6wgmgYbZoRJpUzdppJA+g/Hfpp8hqpzvL7+YrJ7aDp4lyhgD7
gTkC9T+CT7Q7D11TEWWBCSTxuEhBIYpqWEixEpCTx5k1IKsfj3AReeNubzz6
YImJJpSb9eR6k6aOzm+mP736jfrLsP88FXe+920MbwV4eD7mm6BLDRTWa6SS
hmy6OGAxEZlVOHOmT82NiiT9cVjzh6Ih4oHzhO/6f5q4TZsuUQvqPf6nv8rH
QT9g0Gqr7UPMBXJETwfWcHv/EESNDlBwTprFCjUq+0Q7f0Y7kqtPiOY5crp6
k6hwtair3fCODssWTpqUmol9zfwhxbjNsONszGI0FCqTKgTvfvA7/7RZN3VK
y6YYe24ULGe1ouwjppiHu1jw62yoteFVwHJ/GlqC+sxM2ES51l0PJCgWQOF2
LLKJMueBGyssBCgKSdpMmZZllaaNJxlj76FhgGk5jAVyfDmkW793ddC10mYj
Zu6k/v9YYcjY+OTKtWVJ8fiOiHxxEBckkExnvRPZVyJReYS93QEig0JZ9OVq
dDuBpnn2JnSJk26tigS7eVmucOVrqICO6DwJ2Ip5opdJoyVXLt+evkRt8PWf
mkKd0WaZiBBYWM//PqOn/+qxnAodi8A84ngCd41jUAP82xLSaieTOfjtaxuq
+fCLebg4N9IBHXj0dH/47kAhY2/iuASWxya7Qsr7uu7moJP3NBj+Wol01Qnq
CtflGk2QN1PCnoJeiODlPzstXpwhMuLi6AUtrV3KFJwsyJiKi5TmKOc3UivC
/MLaCBHHVEGG4gGb4bF2GqJ5YLMXBMp3V+81y09Io3gVbHK56JQCwSQ7Tfzu
tcz8dee89tfcjKoS4XtTcO18yCqKHYvLzxRw76d0gVN2/+D+MutvMNeYIkrV
5y0AbLUM4hx1kNOYkCbonaniLNJCgscjsXlTg4zvwudv+kSgy3bQv2Q/2817
NlFa2YizFrFSPdOvJS0CL/V/6wBuAmDXOadlRxmNlAeoqygw33B7tpZvbsoI
GOdc1EK/tsS3EX91Fi2xD9s55hE8DMZglywCXasgli3a4VIOixbjyW6ASEfN
Wx8kYS7r4AE0QM8+eDgQjkAivhnZgRurOvmVS4iPriBII5Y3m89mVZMcqlis
S9TyqpFTnNYeWPZwgxbl7HkHf+Vc+GnOR80Upg+0EJE67MOcj5a0It3SAiLh
am+ZoaxxSz8ZU8HhpAMw0COlij4AYeQKHXzbXmPTsZxTt97Spz/sTvifP3Vt
A/5j8Y5Vo019SUDieWNciHF7aKUdKg7f1uhE2Lq4iBFXX+i03VlNS+GBj/eD
YRzo8CNNsebuvLsaGMdh8O7FiqDauwY6q8sg7y1ezvSYzS35l5fGzGNIFvcc
lChsvMqn64vyD3Nq//okEwmjzXvIeVvlo3LbHnJzlYR/bTS22Ywqf0x4J+qL
TH8aGtitozaXoBYui81qDBzcgckbuxWviPFfdoVDtr5/OnCOhVfNnqbn+ZbG
KB8q7LC+BXQsnyf3uD7UE4goaQGfCOZTYCqxy4HvK6jXA5LSB/CVjZeXsvKe
sQ7y4dxg2wAz5oVW50D9L3bqW+x7IIjmlLmxE1Wd7eSYD2rFdlouUs+qiBD8
jIsZAjFnFeni5XbsBf0joLYvul5Gzf4fQKX10lw2zsTi4qUmTwWjpGM2mKsq
aPS1BjJObfKzOv0CcR/h6VduUc9kHu3hny6AlJIoRfrxeACwv91T10Ra2IJa
kSh8GsXk4u8bhxHt7wCbyJXeRjd3vs94ghgXWcpzyi+bGCSQe20KdHUhx4es
FftI3js06xpVrc+soiKqmvi48vhWj5bnGykYSA1i/rTn/y+NYZtCacZu3bPD
v7IZcYQsW90ReYtz9XMEqliIP3zOHrIfzamVgcVNjinKGu4aL1IWvgB14u/6
tAFSLyW+5HMR8+8k5ZD9JaiHCfE/kcS6H4PL0h7eN4cpN3QhyTpX1uVKx8I7
QaguyIWUUy1N2FDzJKj8+bG7S5xdMXt1YnJBCCpJpFtRmsqy/wFeZhjYCEh/
Q4KkCFtVOOPUETeiUbMuMr0kLJ9unhCsIzC+0054PljY/e9AFuETor049pWa
vrURHGikNy59wXE3hsYhAAJkV0O91LqSz7nnNnFXsH1/U0qdkzw0ZWJpS739
cYNb+4JuMTWmW5S2QfouGfQQhIYhsh9+mzjQ4e4+WEl99vduLCcJw4FuL6gV
arOY6wdgwIvqZhQDEIJ3ys7JS7xjv9ETTe0Frf+4Ms08YaxIfUT+BH4dwLmj
dldVqSwvxjw4adhbChMgsKr1CvNQo0YBkEuB/Ul3h4u5up7o/xZGzeF7bwiz
19DrCzqtrOY5wQjQYfUDT7yY8Smks2E8teq/Kd4rR4AUmWhhRUK5JQvcPHsR
Iz/HJTuyW6c2tEjqV4On/FKHC9DzGroIdoKjMjeVAm+a9KNZlD4OaBqo1o1I
BviHZ4wG+dt0FEcbbnQd6IRIWhvhK/95g3GqJqxvKCpEWccJavvFs7nvf2ba
OuS1xkf/xmj84YPe+1J4DmlXNMH4twMN7wYumzMJI1Yak3jj9dxVf4agdW/2
blZMbMTkrhYm1O6hUFTW1godmzVRI0OlyR+rIGaG2LCqcHaXcAN65GSQFcuv
MUrOsWEg7nDWvcM3y9Bryeo4sfp3yC18cdaa4byZvJ343kvTiKUAwOLAUxo9
om6EQw4bgHSD6G8l/EfuwqN/SB8SvZ6ahPBXngH/9n1FZ00YFH7u29xf491e
jr0LgbR/5kWAJh5dSG0umlQoJHMzf0DhMvS1cFM6e7KUvN+t3vU/fKBwnjQg
d8Zqw/9O7aKWlkRcJaHzNrtIeJAPxEXSDhAAbRoIOFVQISfZRH2RgtSKRCdy
UB7LP8UpdNam9vrRSEaDQ3b2IBud7hDvte1LiQwsr+HkkHRBvre6bxG8xZgF
7i8UV7AGbfcDFZzffTzg5Y5cDD5M7VC69qdOx/MvcnjbR267BdVkN1oq54xj
hm0vPEUGp+bYhDob5V0aLzwL8M6j9noPn1IHA+pu6H/xj4GoEtPJRSxc59tA
1NHybtjvXQmZ2La3NODqL59OWGuEpMOO9LRh7jht648+9uVMw7lXMKbNV/v/
2VHljeIHOQYkrI6ziSfU68QO7G1SKEDwVWe73m7rNrwWfau2zTPUB3O9Lfol
sjEJHmKZWYCiIdmPFCGbjG5KzOROAeApUbPThsxTJJr6HUFjcKq0QhBwYvBd
94B+TQaXi2cxijj+8RqTTQkJxx8dV5LJr9nXBUBEQSvsu8RzUfktVXoUMijU
YkHcmMmsNfuxEyiVwhOM2hWElOLxS1/IVCr0HbQQ1rPtkk4yRKqpVE1rHNl5
JhIEa7vi4yvHRwCiIyGeeVT8E5ExWrXRQDkcbAXkUF8XI1G/+3Erx6ZjG6Cm
CdKlgQcYaLRqFcxE/YW/cGnNk2jz3bdrKV+dGiLDp+7IPI5y1VA5Z1auRWkV
TUpfrOiQd9tbWSgwGOKgdMNgmKiki/Ms4Bu9JF0eJvyzFy71LvrVlbWdRYkQ
BFwQ4IdQIpsXEELkJX136Rs+NiBJuHCxscw6XYArG/NQTSYyDAwkMNHTckzY
WtZExCK9px3lrs+JXd+M1EAStAc2Havbrk35IVYkKB4BgwzetD1Ye0GTW32H
T1ouQoqTiSFVw3AIrajK1/j0jrBnbtHkPWHqjFSbUzROqK0ibgJD+65hUeul
Syqu/EhhMaDzdHgAXY3Bk4WKLak+McDi2vXY/3Qygb0XhXu90KI5zQJCaq3b
iugAPqXhXkp5y9ShPfQbuGijP3MnYT56WnhKkOCc8vfIkraAwmilzTHieyNh
VqkfqctnFY+HKbYIqDyOure6TiSmM2MhJW1Jy6Ylj7J79LSNK6szyPq+R02/
+9BbbJjYct/OUXsyoovOJcZexZWmFm9w0+6bcIvjCT5gkWk7IbKtwB0g2H2B
tm4gbN+ZoC1MKRFVckv4Xk3erlsKE3+QALflc/5NFR7HOpAnESa6Pxx1VFEp
u1NBKB2oIpFpicPuvJ89eyxysFEz3B5LYmII0SYwC9rc4NXZJXqbwrY5dU2B
J7S0WbSbySpBlaHCTfY3SbIzbBnohXchJ1uFrzhXy8EfK8ShMvti4rcmaFhb
TSpWbhQr9BKNeEm0IyeiuYwybERjoft1t7/zP4IkPm26q84h236tqtwP3iZh
QWPjLFQ0SKAhXFdEdgyy8W1Qk1YFBfV9SuZsHRk5IRk5phZDhMhQYPWz5CTA
jGCslzaiQP22cEHVfkvIsjTOv4fMswBXUg8yOxkKgxBrXmPDHOVlvhVmW7S9
KR9dkk7NLvEvERHt1WEJys0JyUF1ZpT58w998m2WAQJbMrfH8ddV5+eTj4y6
28KiO1xqsGVQhqUULYzvBeaPGnu995TWdU16tHUVXpIhhV9g28WydSeHJP9v
LJz1e8A4u89/TtB3tp1DUUYFyQ99y4dlurvYuS+0xPgL3UpoB4uiUH6IR/14
FDSNwVIwXgbc50qZ3x5vy1wSLEC9fBBMPn18ftynXY8xFZa9Qh4i28j9g1nD
f3a+NRz/I/aLw0mWVcEbgGgiIw7F+Il035cNa44nf0QTKPKiMa7K9GaArfBV
jl8jD6W8XV/JqDCp1dLSFyY/hUd3OYgK71R4yd+M3oklBEe8p6QTaWIMsRDn
8oYkPzyACuZ+ukeFyzdjgh+jyEfbHBzA10VRYQAB+ZmywrpKkb8poHHe0BAo
rSs5kcLBXNQt3fD7jopjJqxOZMcR5MT9rCt0t+HzlUl5b2+m7mX0FXP4w2IY
PRos/+CNqNOjDGLY3fkPCodkNfkgKdA9vq/8lHf7DvmgnIyk9NC1JAPM3OUd
mUMiubgpJ2qZlDEhJmC78975iMe968NeIL69VQkAUh7z6PUEVJqJ6WiwZYTV
ZEC0utj1m19HwVvUYOVdn0GNz3qCXBk8b+YGNEEJLNsyDGgItV41c9cF9qor
8EVZ61E9hkD7aOIhAY8YxI/XZ9tp9laW6xaKbs2C43B50uVO5KB02BkfsKA+
ZpDweT2gvMYMV7EY5VUgwf2+rvxaz7HxFd+WRfNkq4w3V5HachMEkFR0mQ0l
RB00vBbZjhZqVmWX3tjkuCOsla1yTX6SitCfyTmMCQqAOk+N8XzbHbxzu071
1Dz8nDNwPhttpPMAVMhxVVTBuJgYeeF7bQ7kPlDDmdL8zC+bsXi7dyTXuQIM
o+0ogENmu4vY0wz3iOs8qIpvi+R242qYa4yh59SbbYOk13SuJHDYtJgS1X6z
yg/LTkl3bWHtqmZ4dL1hzedqqQ45oCiehOQUY7XvAbULWiUw4R7JUP2/FFWR
L5LorRKtEqQo00PkHQefNK98FHmEkNws3j/qdrHZ5OoeJbFPya68zIEYXNCT
u1gJneoZN1ef4xeyivePEzaNWGuhLejB2KGsqLH9D8ozp0R+0AvveaoYMF7G
bqqdYNCmFfDfPWO1EbJh4+ejcxRqn4PXq+6Yilf5lEhmRNjeDmantcoVpdzi
NtIHaWRTn7JV6ewzdGJQXyU6GeKdCzY91/uYE7Yyu2z05Goba8jg0nxZvhFb
UX64t7nx5p4aYTTuahJPrTsBJpXpBg86YfkqRIBEs1/SUZ1DMbKKyy2fbAj2
b7xM9UYq8YEkwxhn35LVypbQelY8Xuxa3+hlMpaarwP961K5ySCBs3+DuEL5
g/6RSRflucFiUcpyEQU8h75nkTzvny1yfskUTkBcR4Igx1BUXy+xNoblo7bz
bBNAd0Byg28VL5jpGS1K6NGVuzHI49zCTiEcuzAe/ofVoIKdQEDA+aSrSg5H
aKy2eXI1J5jPrkuxPrLfXXpyWP4L+0vMsKTOOkTeVZpWWXRcTeywfoRRdqxf
2cSJlIfh8FpSzytK3makGhKUu77Wvl9soUdec8WhggpnfjOA4m15upOYVGvA
b2A6Ly/lmjfCqeU1UJQnow39C7y2NGDQ+TLXC1XDqjRqE4FyEpcKpO5m04Yc
lPbykeji/MdY/9iQWVUCXWAN4Imw57Et5Z4ejuHoBVHAjoRejwyrUwgCoZOv
64vLvi7tPZiNa2NIYz5GcOg2P+wZwbwym5LfcVIdcSVoxhu9GdXdE5HL89Ci
H9PaxBFQ01J18s5sf5Y3h5+Wn8ExQPeTYGvZtOk6/EPnGRrTr8ht045gwi/0
RvBU1XBdCyIb5kZeun2PBUzO6Fr4oOk9z3P0p4hgbOwhfSe2J5ToDes5df/c
hW6alygye8P5H+UtZxJJxnss1Ds2sJAa7grqEOvEiLf6yQrRGQLb5Q7votcB
uceR6C05OqbnkChItsSGR+vc3wfMgUUooxTtyqo5PxOzTl0xnSvpOp7xPaZ1
nspkBGkYkBcMX3zqd9BxzQhZ1WuWMptEUUJedf09iJJPU6qbxISsGJZQoJIg
f31r/CWjI7IrMG/cxSL/7bapsWQy1VUF/H9oQsFwJBJP+/AoRlKqIMnMhSz1
m74CFlwaR41XCuiV8Lcpmyr0D4Nucox8+hBjWS8dGKkD4QBd3xYY0u3tvbi5
pcRdWQmb/POHTgZaTf8D27RgsdgmQX3HfVFEVyepU/mRqZP0MNE5rFa9qifR
2Btu0q34puog0tT1TnXqjXEfovgf2XcROm3mpEbbZyVht6xiTVTpZ6viupan
hIAcRmVHJbt+8knBQcdtSpW5r2B348dseWE1SnNKKGD+GpLytgDZYvWQ8bUa
TTU09+2Spf8nib9kX/lXdsPvKd029R/2nIA42qChO/riB1gzAQdKTO00X19d
cgcSpOYUNQoE1XZk1PTEjJHDCOvRugu2uyR0lwfk6WMQJMvUuzsZs69RaSEq
SGwDDRi2Byp1SNvK6RYAxlKy9faCzOkdHsmXGR2XaWuSOdTxmHZNggRCQksH
/IkxA8daor/rb+q1lqKZlxFW0t+kDzH6MaGmQcUl9sEY/QlAjIuzZyzviCsZ
RcfABuUxXHNg7K+T/YT+9DApcezQjFwHfEpCdWvDSBhvOn+Yxkzc8HG8B5cB
Qmg+hnL9zGX4QlIsTXtUfkchL93qdSnwjpFLL6jSKgbyeJ2yw287vXSM4M/b
QpxPTT4x7iDersBcznD3Q88RmMLqiZXzrCiQfAnihib4eeKzGG01BEJVlxTh
DhgdsAJ3Rw6CaHxJ/bCVZ28ARjX09jE4Gyf1Zpn+r2JDRvrU8TT0/uVjkb4w
zwOxX/iTKYdUhdBiHql+mKD2qL/q4MiVb/1wPXaxsGEixEYqSO48W8eXh42L
6ldYpNP/A0d3kUJmfumaXEuRk8a4xZD8KDhVn/H2+anZG9pMM6il9j2oHY56
zdS3zpCeOZG0Mp0uUBhouRXkG00ZfoD+XxZaRmHciUkBES/E7mBHmuCmu5vY
mTbJYx+uNirKxvbtN6xu0BOm50MqlpVRZ82dqdMfhHEwjOgRvJLObqmIOzb5
49nw1H0WQRyb6TnL3VQE9ZBODVIgkYQqnqFbnr4U+Gs0kZCHAcOjU3UezeMf
aPuQYktr8TjUNqufVgVK39IjUOQJDTapw7mnXmfA86f1yF3EU/nGqOCocPkc
6FQdJyJA31EmxYBlM5MumQvOMed0YXMqeHQ3Caaj6svQYabZElUdD7JHcqcl
I7DEvNvKNvqWsLG6YU7wOXVKalidla3jj4XyH0pKvtyq+Bh72Od/GZwfX1QK
Y7zc+Xwep+S5p7ut/KMCvRUEbK+x1fSknUXEzsLCzIhGtMHGFAvKpXhfkg7n
GdSEA947WmJBZjSi4mjcUF5LHNUJ2RKMtff4FVniTq8ZXlT2kIXNH/SGgNnO
ZLIGzzuGp/+mgtA9VO2MKu8BJqXqUqvRB0+nru1fCZpcDYFDZYKrZM60DTiw
CJvRFLp4Y2jmLcs7sPWURH5vX9d833lLFEFRrz0HRMfJZZNc1wPQvuiARMAd
DqosWnClFrqcJk6cpvClo65OaCYhqd/PDlDhAKNoBhK5i+w5rvaVPLsBqnzY
6GyTKT/9U9QfmYIoY+/JDK9F7us4k8i7rE2Bn3N/hxV+6MzPCc/zaM/eSmKQ
ZXEnCca7D0SGc2GVZJlspECGE05Akd8+hGInQWLaCRBF14UzNexfrxOZgAC1
K2fcr6b2lxw8GCfiVP/C8qsdvpPzhD2RfpNxJ4/EDke56UbdTa9GWqudxtUS
vVhk+MPj8YoI7hWyS7tgNj3rlvOmBNH9xBMBQdRPCLtcKLwWipmXcEg1XIU4
ceo+eP7j7ODSWhmJmkUvmh2ebI0JwmZsRlEC4YrlnR+SNkza9sq7y4jdYwRl
MFdm15dJVe/UDkopqjrDfY3rTlg6UDL1p1TNHr8qNuhgV3z8h17Qgw80gv09
sN5hyJZk1hFyM3n11zJbkkc7Sfzk9CLPi3+3/ECwOpJFFusCUa10WJd/7vDO
/Ajz/gjN+7VtsyBzCRLjbBlfxLsEsoiVy4A++k4+1HdVuzIkh63of/Cm7QMP
WqOERWms4Uw4OwKklJonj4FZVGxJ/3m2n7gh5pvlcSW1Kdlp7Hg6PM9ca+rJ
y1hDZ+GVRVku4femc1lpU9kfVm4zAOkjFJJheWnTT8ro7TZ/1H/k2kXbbg/k
3+jPtXUKDzVxqOy7hYqONQW5XEGs2y/TdsOeLlvPkPsganPQodU+LxbnNMzC
DkYj+FAmnsjtFNQ7H2Ap6WggZt7gmchmEUfvF9D6u2/D3J5GzIPbxJRYH1kd
tw3jgMsjcbOprRvWRuJCf7LRNH0IE6u/Ln3dNx6Cz6fMIw0OxVmX2CDoUyo3
4OZIO9xbaqAlXBNjJfdNtBONT7XE+A0EnihvKgq/a365Lm1CMKPVrWozUiE9
3BePZCj9V38WpFx/8k7QJBZ8nJZ7SfiMcvBTa4RiN8x9odQgDvceVRxiFLFR
mUKoi3gDMUxEWl2pD2uqI/V4VWxLVpfMt+fri8JkuUZh/rw2LgEo6xQGi0aG
UiQIX7UJ72q5uxhJTfBtUd6m5UgPaaDgtnamvYG4dvDIgv7JQ+UErNZhWu5l
Jira5rEUPYfUZFgoRoE8zTe7M3DdueWKEZaAdb6YkrAYLyJ4/9tBvkzKfNYW
znlg1i8uUhnkK0KxgASsRbl4Dqg1loKOadVzo38uyv4tzPyZnYEhOsXHF7DQ
M+PUhgCSVWg7Zdv+z5CJK8GPd7mOWhcMOosEwtyIOFt2Zl/79/iCQo/eji2C
DS9stQKQugIXCb2+SPRUjOd+41dgvuZrqn+2THsAOmUPoRpWBfAMP2dNgo3g
UaOhgac9wA7hha3FKTTZ8RG/Lsv4WniojB2/bLLeoigYzs87z9VHF/Ur3nbk
tpbZxWKugJYpZ1rdpwjJ6vDb+QI37g+uL2HJj65+4l6XGQAmizHudTNum8y9
yVGw9euad35WwKx8cii4IwWE/PSmYzJqPdQDiscLU9wHWYkN3YoY/JYq4qou
u9yBdEeObmkmiW1PiQVFKGAjn4Iy7O7TknjOp8Mm0+1n2cbNa1Ng72QdE/D+
D1sY8UNXhHm9RW+Q7WosV8k5Fz6YYM3hgpJ1aykLZkf2KmljwDEB8QB6BxvH
7aSsM8wO4MzQpQ/DtVpAUCivXEqs8pOO5cT0yHxH3guLre0bdUSKiDeIvg5u
lhguj5ErJ9EPNEAs8weIiH4g57n0BaAqPaZ8Vmzw2FFxNUyAS7DQ9mrmNgM1
em2JTdM50GLLYEzlx3aZ1T/eNHTDI5cLfH27I8MFWyBulW+8vGcGLCsxW/2i
34VnhRVJDn10CdHHrrXngj2k3IXkPx6YcFC1fqVDsNpgo4yy28QWLw7YgWFY
ivTAyb5rfXJ9lhV4yOlPb1MVSvw5sasZs1MeBIyILKx30KAQDm2lgvrDPixZ
Xnu4iRedNexUl2TTucJQXHIVUim0toJ7LOdl/rHFOeKgCYWAgLRTVyy7lpXN
j2gqOKPNkKxMEeTME/OGgz7iXfCl4+uY6cZZw+txXoxsxXAbzsPyrf1kCJkN
M7GCFiWlxvJapA3GBPnEvBi6vYvHpBNXV+x1YT4nykleMZRdGAX+mWJoJdbm
vzKdE+8cC6diYpWh0H2Lt3kRT5+UicAS0RjgZhvXpaUc9zNzS8aIm1VOJ3fJ
Pg3hW6FmLI5885atwuv+NB0na0jCgZVeLCQQtqYodvXU7+Ntbeq95k7ti4LZ
5WN6F091MavTIj/QnpAsT+NIva3hrkVEwWSWBi9/NxlqrhiiGLycLdC2Fkc/
Hiv7b1AdAX4ZhfnJIqSnbx8q8c8+S16I1WNtRJld+OvdkVirJaT+cD1ubtd+
xobBIQliJsyu/Zi8rbCSr2dpv0J1OzL//hckox0j6BQQDtbomW/PjEpjKx5C
pKijefhB7fdvi58T+A3NqsSqJvH8BhtyNyFsWhF0q9mIws4fT1RYybDZWH+9
HsF6lVKaRyLmxcEw5BtjFQnP3ws9xNDO20RuoWibUI6g5V4O/8I/UxMduqeT
CE0zB1+BGONWcMdRGEpp021ISlNHOOQtRPE6/iW/Rx2kuNwJZHJP+gkud3s4
asVgQfs6gW+taBdCxEF4cqQQy5QlL1uzXGDzYwv35sdXSMGU4qAZcSNtSyMm
cMHGbeQE9zgBUhBcxOD3p5iWWJgFLfXrqO9EfZfRu5hoos9UoLGtsFp9nZKJ
OBeQb1tgQ1/PyCMPz7R06l1X7BcnzD//krb6TnWTycmO2BhX6RyJ0qBLrGaN
yAEVKpCPYp3/S/BybKQFqoQ1reyXw/htx0Gwzti6Mi3drkrNVd2JAAwvpKPZ
ufYjH6xsfPItPGx+V4rHhaYWvUgr3O9PTUIWtWSVCoKjcXieN4NxPXX4fCft
e/2hGsDwrZF2qhi5C5f5N1dIx76lB48te4jF4lc+0uUVpQhg4BvqGXtx8qcj
xJt1SHDgBgsZIopmm1SsOFudqKb+QM2SUhwtvzLzaBBWYd6UoZn6uN8VjAK+
G+UrrytHweM22gWM3F7WlF6VfTSz0SlicSROLMDcqxVCbS+T0V4I819Zp+pm
oL/8V4FtJErX9KrMX95iyOuqaabS607czSfhWfO/JFdGn0vWmvQLdW3AHFqa
58GvKaTaDB5pMtVQxx8WUzELQFcUZf6Rq+wrENW9XDW/0jYh0PKXaT1EJP04
gPqe8Qa/crW04/xHkSeZMk/7ik2MhQYJWPgBngM66eXfe+AO5cyQwLcBXQEa
LLJzAKp2M91Nzaz2TDnWaG5qa8Df4vM9hJDEEw/9IAU9SphN265de2PSTeaL
Zw23ghrWGnI5WHzXZp0Js8LvPxkNIRRp/S9Lw3Kui45YHOncjYHcM2XfOY1f
jWf+yngHwVBpXuw84yiTl6WJfhqAM/cp5AJ7RpIwZBYgF3QJ1CIq2qP1U85Q
TdQXGAspBWyDqoWDhKMM+DdwoFyUPi7SoeayagJuuSkL93lPIMDcGQXBeS0t
VXdYUsgoGoPEcBQNLfcyPpe6NKHry7MnSNjGMd8/WCQZRzsyIQzj7w4N4nIA
TRwOoPJjQTNqMtIOywt1/dxuQQz6traaS2f+x+4lJ063kEjTXoaoiJQxNO55
pfEFL0gU1d7mcZku+j25ZtB4wm6Vid18lAyDBOTDSSIL+2TnSaTD6lqihsXb
tisQK3mvkjAc4+04u3R8AkdJ/CXQ6fjw5bVWea0JWbq9jiICpFbGd9h96SCJ
H6wztxhO6yD47k2TKVT6knKB6DZbxDfGLkZSBR6CQ6rwCpBx0hImCkDG0RQf
r4s453ESQzmiInHyBLxypub54lKyj/scrThzA6CQMU+P4Gq+4OwiMbtLx8Nd
GcBqrS6gVlGZbjn/Iy/7mmr1K5l6QK4sj/SY9uVf2JLYcVGudjs3GQjJYHBr
T4R3ZIcpXNxS26iFoswLfBjJEMZ8BOfyop+k32q9j+12WIWJy7VXN1WggXiY
JZIKREwKjOE4ytyOpAeWu1I0XPKMHfpzEb2OdjPSwn6v4GnM7Dds3Tc4SNd4
KpCKDs/1cXnwmN+EcUxy/oNHhtyx+EjeF2L0G4liR5TvfdqeJDbTVTRzSCZI
+mzISlVNmK33heNyxiPjNnaqfDOedBwv5sZC84mKRPPYrFVJnopHEJk+t+5B
mKXeHCr4mXrCd4sNOXOpl0B8svBtO1XHRNDp7FGJwhpT4fm3jk76DY2euyIg
YK2Ydb99y3sXMn5jXkLLk+xMc61vNa4zkZeVLunwfoWRhfqzMpDuc979EYyp
torLin6hYD3IFHZ9jE1ajCF4rKHDBl+j9IqMyhLl/h3DFrFRSsMGQhwq6tSn
k9lAoHx/NLemEqdzvh1cXhbpJZoi2WQh2hK/7EVbJty1DA9wrEY6FO9HsT5a
nzfeX3P4Q18pBq3xtQcWBtsM3QdIiO7I3RR6ROz2DCR78kmVEeZrzvgvADpm
GjLOqNlKodNvpqaoQmub7G6ZsiwVi1hJzBSmAdpKAIF8IxtrKR5l98bvkcgl
1pK2iPSCk6SH0qHp5xJ7PVXL8ZwekfjQoxEfV7JwMiJTMF16jMVElggW2GsW
N7Aqiq/IrVfGqOTs/I9D6J0LWc5htCkZNHeloE1DV+59hwc/T8gwDdMPKmNR
t831Mf6LnkLuAAGPLCtTTxeqf/PrNU1fhR88Yvq8b8skYD5szeRlqCJU6KRw
qJhPOD+ggBeo+rNFYOKFvmAhk7krAdqdHjnztJwVTcf6Nz7UNaPeS5tTfdD2
b7eqn9824Q+xuWLWD0jPf217tkpkUOitMTJDqCDjeZpa8Zt1PoLs+vg2NSS4
RGlKX2CKtf3L9jtGdb5SUEFIhfuTDEo74IxBSsqoP7XY9lAbUi3KkO2VjP9L
iSye7WgMvlEX6SiVqn7tWAlWwnu+6bOXc5wMP54mGFR+ts9OwIkedigVHNHQ
PLvCkuOMIzIfG/7VefCFBMffKVPqFncqABVIR6OdVimtKVELBJinQbyG5cPl
DGOZaMKoyt0Rsz6JQLKTSZkNf1v0gw/b/5picBgF6UqTbG0QgTc+cEJdlxNk
9qVF/b2bcHT3VtchuxbXZvErImvRBLzpo81ksSQn2AeKhzwyMTJX64aAft1V
OQaDPNR4SdcUiHvg1qz1UBBWzxdn8hygfuhwxwk2QqvnGpK1u0dkemp60FwG
M9lIJxaNiAjujV8DUbXAZ+a6IPuKJEt9zVlkHDcp7ihDlxHJfY9A5mNWfbix
i5p7B5AkfXnUgJW5b9ZZENNcE6/Fts5qr1TT2ndGi8NUUIHODpbPD0cjs0c8
ILr37C7SgtxjAl2kbb5D6u5KYYucjzLXC79F6mctAfG+OIQSrCzADqjCRGcR
0G+hJG+szKl3BRQCtbiVOodPiYvEWnspw1fIJvOq7exHWl3ZsaDVVs9ObPPJ
oTasw2Gc82sBOkZD15DhD4mHnPo+KTgRNGjAEqd5L9LWh257mwydIPSVg0fS
3Mg3LA4CO18sCGh0paiGKIh4cYuEOBP+cxV9QNHni1P6RxEq9zBh3ORkEfdw
L5Qddwy+1y6V/6VYjqNsAJX9ccwQnBBTlhlGXGZHRQYly1bDqzXjKs/VcDtn
b9/K+B02zWwLb82ji105rDGF0Q0OzGWGIxa1oblS1Lh5jZG2jHXmLB0jhLaR
8/dBVaEUXi4vVgRFWo6/Wx39qErLjTI8K8J+5ylnjJx1jJSStVA1eVnH5EPe
WXSJh6gWBw4El55j163le7/X2oxzu2S8wRXPkTwFgqL7Hq+jg0Ipi3CoOEWP
aYgShxm66oqZcBsXCoLlo6KSFsZQADGgelmn3h5pD/3GQvXCVKpArRnyMw5K
UDVMCXYZuTYOAobZOMkdhMObzf9FFFer5hh7lOJemIHhUB7ZImni+Jwkbm9p
IsH9p4YJUEmiwavPK+z5s105wyFB/S4jZoMH8moYBJGrbOIFuI82uDA61P/F
ExhNdApwh0DdFm6fAj4jySqd9eWFdTNh+YovJbjEf0iYpcbrG5XyuNj+xL5o
Fq45+q9RYKOzoPjLEkYxtyvTP8dVw3YhJMYI9DFXwQsbmMQPYGUgTLYmSw91
cWS4YIQj0c2v1aLL9NavS/GRoIswCY7jVON0vpGOdc/8enOIXD+tfWJcpy86
wDEGcUFaILN9IGGo8H72JjX9Gb4ZIebHTQAMIcKAudcwWqG6hhKKhCzx7o93
0JB03Uc8/FgpwyVktpexCVBdR+Q85z0MIL1JiJyaRK9jo3gZFX6wGpaR0s1u
YKFG/Rs1xgw+SPPQLiVSeaAtSmhnmjK1ne1aLMb3CDAYFjvb1U+WxaM8Jf6D
UrxiVQihqvezq6gY1O91Q2PKPWvtveKzFmW82FRBzVAO0F+OAq82LzFewQOV
2K8c1TaCsaCuWLikCOthvyqcskU5tLztyFDzuE35YoIxmTxj9KB3zzkVuibf
L1rWQH0y5q5ypxYyek5YJZwGpt4lqBf4CqcO2MdVPntBv6h6W0oq3z7Vt7/G
9lchVhmtDCSbWUdjQ3XayKIoHLTMxrBevN4cyRJF+XHZ9hUqOEHlCI4S/SIt
NeIUvR3Ykh3Py1x++zhu4LmryXfDjHmjxGBD/jRwpQL7qL5cJlTsic58rzH/
oJY7WJH4+pYCudMLNex6z4xCeO1rdDpIOMJeRrSFOt8Dig2xypHJb01bWShM
GvcoUTfJtXTw/gcQILKU7sTZWUt2LQOCingVLofibfXbs3f49jpgBSYcbrYE
xehPpdZKVLKiFnGo726dB/WSPqPkPOlKN868E42u20rZdacM/boInRXATHd+
ONV3r+51abBqaH10EKcYFFjtrbwwB34VnuVv38L/UoeUhEcqS6bKiaZ8rw1V
oK4WMBHzmTcEFAtS7WL9J8ibo3vPTB/+t5holGHz2zHJ8z3y2bupcDxqMSM6
sp3sv/XmZ34NmqfaI9WA1/4DdhyGE7y+h5vO0qtEfSwmAdvXAOhp5MhAN5cq
OofnyJQbk1JSPyrwNaqoifUHdE6/2i0dQ8IKYQp15ifTAhbplkhhLXzJrgA/
8FAUvGYr9lMseJBMSDi6WTVChaDcllwNPAg6tq9uVEoCK8Ob16V/XRUJ+DYe
Zzex+c3PYjk/0A2HeLHzqGtZt/Q32e1SKD/Qwy/sL6mw9LFhfwuJIFrWiZs5
irWX5y2GV6kWHAk3dk+hqA5B3GyZCr0Cem95PNSLIMNrFmhw8bqgqRAf+4tA
o4jwiL7NrJaaJ+Ly04ByI3M4Gv8NOX3UnSU8enWL+dlPv8n8I9GaYYhxfhTh
sKc/IpkOUnI839sxFlpVAx0vKD8cGqpmg2AXaec7nu2EOy36owXRtS2znucB
GldzNfnnS6lgHVcEBNmo4wYHkaRYxUxDMlBiIRk1nO+gXkdYg7wuFHvMZKVl
Gs0N3+ZBoab1ttstfXyQVDx2eLZ5T7JV7mLvvmA2+0+PFWeHk/F0JKELQh1K
VZPV/8yvdDDyGAb/LyMMFji/0mPrObWBzp/mV0hLHeOgBqddcm8HTN3dN3EC
l02ZysmiqKKoOl9mxc5Kq24FD0lrXonBLo3f53vHOk3qA+2vh4zK9qD02fav
Swrloq+TJLHzXRjq6fSm7QXgMiTTEGLT626WzeE0fd4Y4Fk7HRQUJ95O3DcD
gB4nl+AJPOwUaQLgAkJO118zoWRCm0Y6LdtRpZcbuCb53cK1Q44WPVuDudkJ
GARdzeML3abHLw6+w8oHa/XH7dspolHG0ZAEPiMLtaNJfByr/P2Ntf0paZgE
QnrQsYr60dFtEAJTqtegorrzqyvrO7qRxzSt41z3hAtTY8ji8WRBB6VPPxT3
RtJp7vCckat1lgyBWL1xVrpSQXQNocLNKI2jN47SoebBxoL1hFsRsNyUEd0I
nsaSU+ZsHXRFz/AXCjZoxRsxznWgRBJ13FWZfbSVTZvZHQ6by2WwTZUE7M2H
lsvzZTsExAixxUVET9exreAgrqyWOOlXoJzP12jhuCfTmPiNqOWLLbYnLvdh
11yzm9bONF5tyMMDrYTFGKnvHAd4IMVc6dO4oufHAFv536HBEGOKFP4Az2+r
XWKIFb0ZI8fJlWweN+naJ3IQwe1hNx3wHRn53JCNrJeP180mQ8v8Jl8F6dfX
l38hRy1cne8zGFZ7FkZRx+8BYXc8lLHawl80gDrA+oxOdUjjJlg2ASr0EwmE
BdprkIuDQiNKYs/u7iKOo6GjD3Q60N3YGJZL/bNhp4PrMdVN6lg0I1DC/Zy8
9uF6PGUBg475SxxGweWBR5Sy3ZZZ7Y/yyZ8B2Q8hYndEE1f9hS0bQSgiYiV7
W0Vh+ZiDQvf5hmojw/sES+7TD9V7FIIGmXhPHt2yklFxXWuvVhfXPC9F+4R2
SMDiyzrDWwrqisgJsJ+BFZym1MANXTXjIhmWXlO8w8I9tUbIup5Vz661bc0Q
+zFHi13Ml2BtBxmgfLbmIKyihZjx+4ksm/si+f3Edom6dGDmg94wu0EPDU+d
qiX6xWViNdJUxOE2rIbF6YxgBUssmTclUbjzUB5MSBk5BpdVlc4ucLSTjDXB
aJ4u2U+cSO0bYD+ABQM9tmbNz3xDa9PODurBGiwpmvyc+TbX5Grtjbak48+X
niQNtadk7paOBWOVHbvqp3RRJicjbxH1oDDw92Z5l/w/cp/BxpgG8pYSvqkv
+B6atZz1/RrohV/2LaEvWXjTzWcyYtU8/wF9+3VAPQoLzo78ppxNOduIqsca
mJzIDy/7tSuzoxpTVQC9C7GFdm7b6N2Qa7Et6vgB/3/IZJ0GjQv3C1FFm/xs
XyUl1WP/F8sDlzpb0/4CtFVw9HBmD/SDS85soNbzXCrWyf+AYDq5Z6bgWjPZ
5gQoEwXxajFF9tEkAK7MC4LFGAbI3E0ObP/LkSoV/C1oTo0+699CpRblguW3
oAvR+JxAKpiHObgcuQjm4y/d7hGSIxLLLpmeiQc4C3cTCXd3wgmdacZXWYZe
PN/o2Til8FShSa6XT85aLtzxFWLn9tPWy939T2ksqTi7p4pLN4eXmbrv9vCL
PZJryeq3Rnc7bIka4ryBSzGdW4CAhF7AIT1kyqPHJwhj08sd+6M21bpYhzoi
1PCfBfm7pzIUCZn7c7fYyVT34m5k7uA68YUNxMTopABLLi5zOc9PfS1XFE4U
PyI3Yc5QkJhSYBps65lSJZ5gadRUli6mjGzZgHTQ1vYHLsnukz8guN7BddhD
fvHg0ZFaEo+SyIesXrXmA7wxZ7sh5OQ0+Fy66PmlSEdKCLd/O6DyfurZyQ5m
qCxKI8kULWfzvFjjGme8LMxpA7xWJAr+4impCjrMd8+D5LFpPbi/umu8rsIK
9GNvbzsF4hszaOngpZaqi9KKmakTKPAUY5Q4BXw9XIMJcEkyNVrhagh+8FKa
RdMZhflrOBSkQ65EiNvlRoN5jO+OJofsfPYAl01v0Sr6o3YX0ZIGdbfHg/rY
3P+ie0zPWTLqCeCGAdSYeto5IKUMroNVbYIOf8LoJu1ez/N1wID6EOqtiGIW
ZGC7H3w8nS8n1j4STzy+E2hwJr5ssxMmZvegPIu0qnjG3HjBMiBG3q7WGDNc
fmDsJnLhNuanuSmHusWxKspED4OcZdjG4C5IlBfXiqbf+xS0QD5n4idIyA3V
bDydyszEmFDLSLpKNNuWAq97oV8gM/TpGnY/cUHr6DE3hp6pNYEVYImyLkWA
cPBXZB92msbnO62rn5Y8tMdNTyaXd4x8BNVivQ0uv4igiecLZ4sppMzwZt9z
v/YmHOFs9WDPfTiJgn75lHBtIexYlFXyrBqeyQLMxzocu3F2JIOrmqcfr1Ga
UAAUn2f/P1HHzQ/pM9UOSwCwM5AOwfFJ9dmbJHwjr3/AT1gb0RgWqQUnrxjV
/3pK9+nwbv07Lux/jzmws7Y+LkmKD7HHQaNI5cPkjvjbm3HQz2MRCLBi7hql
3PAbiiLN/0bVHN2DtMPqUF5kRfeGyd1cX4ecIWFrVHGvDXOpBmtcmOt3dNxh
DvxQZoYnX/FItS1HZL49ZhHIXRc/LzD3+5yY1uv5mKXS764iq2rRCi/waHnB
QmTMY5AnCSJ7eFTtqdyabeaqLwn2xxcBn+eBkv72sRDltqzfUxSFYzBvYBda
IlTn9EP6tvuieATpNeGr7+38E1eeeReEEadyBhq2tANGsa0BphHVaWOnX75y
miOUZUB1NXfYSUzjg+aBP227Z+Lz9yhOSSUbfTBlLf0ipYZVxzQw0WqEDFh9
Ry4Y8x5Zp71sOjV0c7GOlSlgq+y2mPX1EygZoHNHQAms4cOPXJOqDV9YkHL/
H2P5RBIO/aBlKBG5EgpPAy3cNupF8iR6P9hzqgl0+MBt0CwdCECSOZwyoLbs
zIpDJZ7c6sh42YScXqqpNjVERslFA9QEPp2IwK2+S8L37rlYg9/UkVp13jVP
rEy5WPIfjDfTgsya74Nib+Y5XD8S2hlTPTyC7s68w/G8OAVVxdmSHJ86wQtZ
eQ7QdX6xxouAgI0Ftyvk60mjBzohZEk+Y4KoGtVs6cX4PA3+RAI5eEOQdmsp
cvjZq2W1RDRANtQJBzIIb5GNI1KcBKAe7mA1r3z/JzvFFg1F3EyNqtJII0B/
jz75BXEgjH6k3+8JfEqaFWwwWpJoF9S3NgrsGcUVvxcSScQJ6PcED7u1KruM
QtIkXaV629FCW/wwFgRvPkKHGAO75NFmUOx0MiAXh/ogwztVdDtzfRo18Cso
sDxq2+LUYwWrHWhjAQeC2jrti8n2j7YSvEPqQqX7lYzinmp18Bya1a/pP3kF
JGn7a+p8WgMo7KlvAayH+ASndxUJzwxfB+A6siG4Pbch2/vb8wm4mqemJshN
R9ZMMtuJfJdQIrGKsAqG5oCm8EYoChD8MA+/GBjRqjxm3TF242OzdjZamHdd
HyrBH0XPTPy8pc9fSEkd7a0TxxA5Huhc9PYaFYKFXg9relytR1SOGl9dd+0I
DRJUAqTCtoqJgYqUmy3Cw3U1LG5RJybV3AE0Yn+r3WkAytd4BTQWSKt0mHKW
zFtBuZcoa6SPLyx7Z/FQ+S13WzUe5JKfl7fE9am2Uky97CZQclThl/QR4o9+
usjIYMaKRQhp6fHyvsfsRFyMijNHfYAKVjGcDPQrQPXIGjJS1+0r+n5gnPH4
ijpe1iYwWoPC6bz66kmFMhShpXesP54lsZaWu7PVBeKevodzcjVcHgJ4opPp
A9CSeU9sPPGNNysJw1lJUAgkiQNoZrSfRqhcaTKxKSKj3MR1SWbUUkdDd5Kx
OlFkE1Rc0iosSaNOBsk7eyNgdled1SsLIqI8Xb3jiSi++JIZAeWYpgG4ZswM
PxhcYupEYOAWFMUz03YNMNluKxPBBYaQ16iiEcG3c+l6Mi1X6F5UjM1MX76H
NLXwQuylhr1x4IQC3KcFUakpt+AVit2RML2LWtKm0UJG5C0g+/ttk77gDmG3
r9ixStcJFzOIS3jY6FBrbI3uNbv5RVzzoQkaIsTwY8Jy8dUzyL1jSOYG1Mj8
ab6ErvFMNlsbSfuDPyOdzj9PhTu1fzj+NtPxB2duidG5npLIdUoJHRx+bt09
cyoW2EtPxLaMoLPh3b/FHyDo8aHdRQFzihP/cIfYFi+OAS2Gi9pHMmAs9dEs
t9yWXdw9fBQTzHSrbolTnseU8TlTsjNVg6PDjvLit2ZcrXaq0dQxctJT51mp
AtbEmNFVHHS+volKnEeT/h9hdVudNO8HyaiAMxFFZxYg7FZGEESf+tIWpRB1
MrVV0W36mQlHY8y4pXg8zliFzpNUW53hHWYTauzNlRKcndOZNgxQmzGxFlZ/
BW3wyFUpZ/Sr6rnSDEeieEz/xdkCDo6ul2uU6y4MrvpOf0GzxJs9zZ5SuVcW
jIU7yEPBNXKgRV2HpsBvXXIVbaMrt8BMMXGNnpKpmBtw7qK1tyvkOncComJa
XiLfgGCbdWhNzWWo9ATuCNPCMYzuuoKlelrm//UDxxcNfLBeI4frH3EZmgYZ
2c6KunmgIos0edUdZuhesOAHr4lwfyW/83NNhHftUkNQFc5dR8hwYP36DHv7
CaBhV5F/mzMYVDgemo8PTturwFbSmKj8a0JDc4mepn3Aa7XVLGix1OeUvRZc
sBE0pQ2IGhq73wztbKvB+DQgqVruQGUazdlUbHvljxfJnFUGJv7RrlttMfXr
WmuyvUPFv0q3lY9f6vKjdbG95Pew7OKANtjYaTbEli9bWfhbL6Kc0rW5EDI1
8UfMhoGEyHU5QlGQ86+MYLpJIgp/GyMOm88iZo4/6CLSxDzuclkfRJ0VkUqV
PJIIc9420acIawyCX/VVMiRimAzhYRlnctxmsXECBYe8+VYkhVvZWOFxsodx
mi28l2hxO4jMkVDA/etXwQo3ct5ZPBUh58e2wUTCSg7EgiaZBsW3FLzULBwm
hJEWgUvsQaQlmj6zNApyXKrSMaMY2562RNbKyhRMIU3B+sfceOoqYvDcCEoy
VeIVCns2bdW6wU93y8VF36utM54cgv/1FwRuiueORaoHuMS6/iXyAOcsmsQf
LLhDFkiDO4bpvKWBsR2kDVU5a7CZrlX2PhnW4vw+iFUgWBKvDwX9siUNfKKt
C7XZtpIKwR7ZnEHdBvDY0gECbUuNI8iRl7zGq3p0Y4FM/gKON3LkrpVVsjb5
TMrKmlKSgKecHIlCyAFGUj4jRtmlpBbRN3X7LQm59UgXoKdxmLZJvnXE7Ik+
jlLUfBvRSfqldZmS+KVjD7bP05Ky8G6rX7bGkNO/mNOkGuQt8Pq8fThFl6H6
rnbaMhvLNpda3fXnpy9lHZgHa4nuXV4Rern1jXWibUip3zYXfIQjfw6QcZGC
BY5SCDqSbEkGwlDA8hkBKLe0IQW2njlE2Jqnzd43Zt8O/2MFADWJn4LWFD0e
nhzl6IF5ATqcG61Jml6n7clEgwzC8YBdL9bDXB9mzQWdu1TVVTqsmo3ve0YG
61762za2ytWSjpPTWv9kjVvVBOC8snF9RFDicmFTWXJ/ap1fDU8QwR4khYMH
7icR+qFbWssBoHQaj24SXK5daMaY0fkezFmqPU/JqEWrXhQ+d+O6N2fWLuRR
W7VJJbYiH4ennzd3py+VG49vU5bSssY0NesrsqhpTuUVmIbcDFy41//tgyCt
WtOxE7A5i3uh3hLyBJhoYdjfKatZDBHKLW3rZ93HIT+jdQ7Yms+n0W/7At2v
fXl7mYRRhGxMYqbNYvPMiTCcnijm87jSjE3Jk8N1pHo0F8IgkjJyxrE0rdeF
iVUs3842ZPKGGKS/QCZ6a+kwGcVBKudp80GnNavSpywXoPM3fCQ0dNDyI4QY
0jw3VKlgNChUDma6LVYASeZXbjKaZME/sR+s5qoPJoXeaDts3HY7ttjBcEug
0QiAL1Yw05EyGPmvtCoNWTm7jGbEeb6POM4jlKAe2V3lJvu8Og9prjSt1A2/
xM9kwE+z3H5wuTIY3t06gXc3BfuWjU1ZbVxjGKdPy2AvbSnAF8Zp24wxFoz0
Dts/paVO+XQFd18/dQ/yWyoAFHT4Tj+Y18HsNya6rgHuxQNMzJdsyhCapuqb
+KnQUO7+Z1vljERcdGseuyuf4YBLY6p+0m2MJjeeCq0fakUjWWbRrr++fOJf
qQqISGLebo+9mlE4bvQK3s+DSmx2Fzlnf1ADQHb/QD3W5Eyja/Z2zrQQ5jKT
oB5ewaFnovERy0m1IcnoYqSlQrRVTfKKSu9fcv+/RJIbpmTVw+skIfKXvGzN
QAjmHSn0xgrkM+/wIz10q7C2w+MmIHd6cw9spuqUeLOZNLhJtoE6Kid5MumQ
FEkjdQUKvq5b8gO47QY+8Zumeq92BeFx/a7rKv6p4kwO+lq4u+4Ag5d7Q0Ow
Q3J3m9RXK1Oh0s9rjk/CZHs0wwvTOw5HacHmAin25qh7flOy6vq3s4nf6tuG
E5wUZ+vsvfu3m9qVeU56pr2U42i0UWdUWRgyhpgPLp0bubpwO0lf3hO4pD8q
KYlnDKlHaNdqVwPlbDu0IoQNP3bEh3hfkXu8ZpFrOsEPcDt5WVWtZMtdnvbe
9xMKV71VcdGwfeTqE5on+w+VsgpPc+iObFmx6cFyO0DuxSr3cyYJ2HuBEnqB
9QTup1wCOXadR8rUJ1R6MovJoKUM5ZsDY52/NWonm9YDZm2n7gekolmzuoXN
pEVIcqiUXQTqbWCBOQTK+6ftLxaZ2q9P528AwP56Wh2gHcDsHIuoETgiLiBd
5T6f6tGguhlYozA9po0gwfYfDfsuVZ2NBVGyEjtDzkdlWrfpdvYgXH7UfzlD
xiPjlBbCgla37YxKvzn2MUHurh6XeVFRb7GDAlV8/FIf7zHTij5LF9bfY91E
uG4YPDpnQ3tMVLBgV80LZAfL+2HkACAmBXsVMDVjoXFknEhIgsTeYF90nytX
Esdg95Pxk+Has2tmpEO8srEwHcBUhM5JKHtBpCyDHcCzAyecSq2NQookExCA
gtI878ZWLj+4HB+st0K21FT/ld+FZhDBnG8uHKS3pKsEtLr9xtuVTRd/WEbI
FkdFgNZH/22fHKkZt9JMqj0H0/y5p7eJ+bWahGPXP8hSRgTSimlN8XfiOWsW
Omxu110c9/bUakfKQgd+/lmn9pQMf3FNaYjb84po+DPi4TrJCHcZACN5gn13
ntyaMbLK+5yF2/xW4dJw1u7I91AcAr1Rnn99zWInzkIlGCLDGCEOG1E9gXaO
AaG2Xaijgb//qI68BIvO8LdGr5fAcnq7r5s6OAdVfuQZhguzscB17nNKMBn/
hU1SjGkqRk/YGaFZSDGtSQa7pcln6KB3u3h7G85oh7V4IohJ+HzHB9mL8Lm5
5ro9YBidro2DeAXMJ6Y6tfSzQrUzr7R4PmceFx8aMlDHwAEux0eueYSXFjWf
xNKaJ/mTKYDskV27bFwM64hLwxaDBwn5++57k/w52wJd5vY6pGq9bVAUXd44
yuSyFajsWjlswifjXx6lF2Y7ed4ZbA6oF1dAaR3BcOdxtaDXPaVib76jfT3E
v68zwMLVYJkhWI6xPe8/uRHAQxnhya1nS22xtxW5mSrUlea4zo355MFCPX2X
EVnlRpLpR98tduri0t1U5XVBmhMEKNkCpq3ovk2ABZBZKpEQF095dleHA86n
Rkl1tHZir76LVqAP0ZTSoOvFX+LEZ6nDrBwxP6Ps2A16O/nneXsRk0TPMKj5
Rp2/nz9B6n2YnGORojPpEArWXcj13uS1kgpJ9wgDIsrPiw3V9AGrYcTiC/W3
AUxOF6AMx6YI5HKuCOWSuf78btD7IafpMAs37NB4kC820Bp8b3LUgPVxKn4e
iMRUsvNo7EFD2hu8275K2grmztmpVyNu25/i16gfEcNKoELiQ/EikXn1ChM9
IZ/m3F18CEl9MV9VCql1XB4Kf+HnFp6hcxn/W4e1RkqFYJOqjOTwN5TXGzrC
wNR3yPBDiV2KxQe0PVdPzYoI2BxVWYGgMSYEegmmwa8lm2TWgJ0Lrxk9MgsZ
SL8LnA1EogLeZ1z/ZKYBBOsmy5c5vsL9QR1+jfhflkKVSc8Q3idivtsVp9Fr
SM/bO2cLXb/pOM+7xPNZGhJp6rPWLGFX/0+tmhYKgWaWg1Z3LZ0Vd0VVt8kN
epneRpjT+yrRJ37TqrEivioMeIbQwvquJthszvhoCgFAaweo5LpWpS+KM2Go
+9CRoBWPZXQXwFSwT4dERY5E+CVTDS/UkCiSbCBZXzPCvSESFgl3dcWOiyvp
D/Efp9Cfygd8CXtePtrMzWtKkNxx0MdLdQxMLKQK7RhZFMY7uClQl672dnKg
cZTacezrtnh4cBHVOhktD7NI0RaKjnTNSDzTkE/4fg6g3rbvrXKA6JotxAlt
fQ8W1b1VRMrMlFKPWZ5+4rTgIAb0nwiGBSsPvLbtajXp3aksDBiAmJMinWVU
pDB0yP8qK3MFXYuyNFkD21gXUWvPEiVy5m5hlpZMjFLWSyJWYIjTsKQAJHuy
XmkoRaaFjIAavlXBMZs7bG66+pAH07+dDp9/a3q8VjHOXzfCUr7iVXFKzSIy
Gm2O8wOZKkgo0VMo+/437feW7/86vIQouwT41BP9M8Se1kNU1uVIeF1jm9TS
P9+nKMq7/DsYvJfuaIgFJIV6j1n5ZDNkDTmUCR3gyg4VjNkFzjSYgAgFJVvy
XseaQpjisxcBGLw6HEd1+RsKwi6PBxnf4YEriyUx8ODJPUGXaPj4uda5Vgy1
ktwV4hRMgOdA412aTKpDDfM2J8x187NqPEe1/wLMm1hwpt2kE1f+FjKGwXIb
B3/LeOr4cIwPOoCArv53Fim8Mn4F03gems0j+xNtsATs29XXdnYeSd3LcBPN
vWnTgRt0lv43ouUUdMh25/M2ag+afQJ2q9ePzk3hnd0SXg9aA0H520ZCe8x6
crgkCV5VVvCfyTIrPsWnfHloA1ZtlYBgko8Y2HTWniF5laJFQq1UFh41cHNO
vidIKPSTeC1xDF6hjR4L1+FCtZ3ARon6cw3tbO2J8Mjah9RIM2Hy+hZdnGn2
7FoaMyo2bJQvZGXdwBL4c3eL9v7C3b4ZbDjwU8WU6OMXJefrXq1FZaixo/oZ
S70GZbm6A/4yHt/u6gZ4BDL4hTRWIVMLvaERD08HmZt5v+/tIKPmAMBN9dWs
e4SrGu4WP65x+HwZBRl9AQToPeRWd6WC5G5d4dGxau8SXDY0+eAPGym4eBE6
B8Wjfunaiaiuu0632m69bN8RE8mceRJj9Th66E9W9GAkkhYPOQlpoXHGhAHM
TqZwB4IStvG56TFYW/WLveBX9rQjYd/c5NtcDFG0HE1U1iMm/Cx13zrXGYC8
EzTKD0kecGlOQaMBq1hBbfWXDpUX8qvt2dbfDy2aGyyck7F4DFVSHk8XPJi2
9YRReOua+xrDys5KVWLY8pl5YfkXA2pq8YEGGv+0wTw4ugq7MxsqcFtHSI5n
ZiqsoWcj3p4am3DM5siaHj9sEIcgFmiZov4ZMZG1nFdR4LNuPmVufuww2Yv3
I6M1kUurQ4HcOJNSTJiMQR1/gelyftm1ITrlCOFYyTKxJHLwv9E/OkPpzZbV
OnUPkb2LvATShFgjp2Drh4PhQi57mij649TCtDk6o09WaYwyn7y3StAthG3R
7UkKgpgIrXsm0w8ryAlVKI7u6q8sxcT3KzVMeln3uqNXve5zXw8xBPvP4aW+
q++HNqkWQGC7utrcfmG+3Fx9u700BaGFTFT+B7sRRDpOZVEnRhhiMAYGpjaD
z+75ZKVF3SfeMxYxL9ZkSn1pC9FYlsoIxa6ujoly8BO6X2ucRUJhXQuEq/nx
kdv5VBK5ULzFnkVljkhKQ3RhiEaxklSn5YXpoGxtkMeE2YMs7ITmdvxCLh3Z
xMqV0h2+51c1STxmeOHjPZgQSVdborwD1okPHaP8w8ItmjH0KWn7Dw9TAvvm
13qSQmF7ixB5CkG/fvSrqCLcOe2ZkOQC6rKP6zUqUnjhicLuTyZU/bD5uAoV
UOrO+MK76pkrgl7GFsGiCNc2JrUPy8H+ZWdw5HYhH5hQ8JkgJqnh1RPPdCFX
eKmF3OKGCoSL4PmZe8+uTY5cc6O9x43N5bNM4DBQUzBtbswX3QRiWAWrGbWt
ylb3pMxtyjYtGv6zFBhM/32eBCri41+2EEsRy2aoTdZifB2I3CnFMIw+ZI+7
aZ5k1Jp+PHFju2SaUkwCVeKv5tIuPLlL40vmiX7gUsIS1SmKWcEwRdrgnbQr
IaabgkF0dZRBDUzTjDqis7FWcKLw8FvBq7t3ihSEHg0HhT9qMbMOXfxh4XW2
wrd72sdtSO4hyxDmM2DtGMtLXB4c24Ul9bg7X7ZN3Kpk5K1oKB0Kx2stjNIc
FQqXUZnImUBFdu3qnpMwQGYfOn4b/IcinW64KSbTI45XVw1fBWjCiWO4+1HI
jNb/ktW8VsPg7LUObxd0LkgUcu93A75Rx0DSv4GnDp1DiQO/z6gANmWsBUDn
yQHZmnxQkUIzk6qyX8cxmLORbwzmlHI/WM9Mpos4DMAv2f85bgMNassysaGf
oc7OavC/ZJEUSIWkB7osNJYTifL3cI/RobYLEA4tELImPX/wgGfHB6HxQOE6
Qu3uPphN9ozK3r7ch90EHrIV+SMo9PD4wp68cLL1R7op7JX4VEa2zt6X0e51
5hc1VUtkQ9hU5LtBRmlDbpFP4eeoFocXvl3gM9FyD9l6qUsTdsL/wJ8cA45V
Qyp5cmu4Ssx10On6g2UYX2FwSVdAernW3JxsifreP0KbvK+3LwtDfVRnPoyl
Vr1Be6y8FEQsLM5G155ms/s2EOqj0KLtIMRZGwYwrbwv3jmwptHBBrfNyxOQ
YE6k0xiB1G+GY+Cs8F5UfV5xxwJTD31t968PZagxgDfyL89uNBPmURU10DRa
+iK15F1wdlomaZKpoaMqUAU+JLpkDsack8v691FYrww13MX45gppSXL8dqwd
JEZ8itCfe4i/FdoLggdxIR9DQuwcgZ27Y/WZKX/vM0ceCtxeXpDsBL20KR/g
G+s9JtjTIyI0gwpftwe6XaJV/prqKgorabKasyQox3zWk3xAas0PUqqdAbCD
9TOIJa8Mn1EtZAnpYTMw+qLkZzUP8gIQwVd+3E5UCEfnPwK5juZAjxZRN0Rw
eVmrKDYCEUukExF1f8LFjO6muDHpX9teywKljBTM8gJVp+Z5CxlOydraNZB2
7VituYiVR1ulrh56MhX/HGWhYKxhgKWI/1Fdb80S48sw1rpXDB8gHKSYjv6e
bdxxVPG8HvMu7Qu+B9pFZcoSFpKQ8tLtv3/eZEZV/R//Gy/ng6BLwjoDD3Jm
0oHZBDmsdxBUeAnzYXxEQr5EklKhSgrziDXqnTGIABJzKNcE5lwZXz0Jf44h
BRCKJonjwilHJVNclNHT2qJ20On24I7Znvd+XZcj59PUo2Lhhgk9hpCPU2mT
NnQkjia9rxKLfcHjdIkegwK/+mpo/0Q+Dldp/XOh3B/OL0lD/JPuGRqCtpB2
XnQ0K0gQgSI4dkFxuQpxNykXUq0+CADuE66NOv+tBC5G4pyD0U49tAhLFNtK
fIaCxmXhTNk54N8XFvpm7TB2w1MClf0WvVhLPTypbjzYnLQWWOI3gWZw7+/J
164tx5e+K70D0MzBiyifgM89G7Do6EcSouSPJGd9eeu0M7ipLXG/pRCjEJzh
mLsUNVQu43kk+hBrycMTmHzOgp9yq2mYZB0K/YRMwyh2p5bzBk6fMhrPnij1
qDSLmj6AsRyPz2taKMHCi7UWvHvrUCLdQK3ISUWebIqQQgY58plnNmJxhGYH
gs1tcF2ori/l409Tt1SV/ZwPoUTbXR/M1x9n2OJBPO8WTUW2MObxb7CVvrsS
eL8r7y1ug/mM8onfMFD46HlTS6T4KFGEj0o9uaP3TRLQvfcKZr9xlEPVGbei
5i+v/3dloNyjd/m3aGAuphsqETy6+FB3oENzyBLIrMMPjcijazyprbJlQulC
6Lm9KW5rd+0EvtgH6U4JoRIdAsZxjMUgcp+UXEztlKVOCkvH1OA0uz9vrSiu
172wEIEPydyWdi0cCnzVcX7ICHSUf0jm5Pk38SaB0hzqiz/UkOWgwioD5Jd0
gOk9Gx2+BE4O7VzeoLbHErq5UWTBu55vSJVFpfsqbdoHqmu9UiLsFr2fj9BM
trCRXP+xFEl8ZKzwNOU4SCo2V0hV0H4jbLkbiWPPaaTTpo3/on8BY+NDQfs6
6JOLBtMuRx4yVkgh0JstKAWJmi/f2ShmUuCnItrBBNJt7SUVnfgEjXuAbrwS
FXJ+mWZI3v+WcHzJfV+GotSA/Ld3GS/+Dv+loGl7Kf13syEsbVydofNBHrIy
LuQPo9QccQEpRpx/1BdzBYd+1dA7jcP56udlZqxzDt3nsLlcsgqpPc5s2FcG
4psWYdCPZgO59a8hzQ6RBhcU3ApsoCV1u22XXA69K+CIebZrl1le9OomI9M+
Ot4U6Tu0OBQ3Cq6O/rRx3ELIac057dG4Y6RiXHPZWCDfdtagaPEc18dCEJj+
SFrJKNJO+SsGKLIVQbFOoT0C8WKRA74tpQjZqDr0W0No/9f1PuJnSe1IM0uF
p/zZo6OBHyYlqpcigi7S2rF2khwM+JKQGdH1TJIKen6hOyc+jH4BFg6vgxQg
FGFLA2Y4wKU0Fe3z4vAWTPGDnP8kvRyuwq7gUmsKXyJa4dDQXqR24NHQsBuH
AQeUwFDc0ILMZskrG8PNfIpr8GdUApe6GBj0MmSOARGoRnzOr0MT6BWSW+k4
lF5DW9lrPMvoKn+tNRQycMmxHaSkDNnU/BAuhimh0OoB5LpgHtb4bHybl4UK
9RoaXy6j3vOSodIT4aTyow+Li2OZEe0V6zZQibWytXTwLSawT7vB+GOd11Ec
7ubpvx4uSUe//UYVn81Us/X1Cyae06L6IzPedO8XIuEt8nIsque89ynUrO95
abbqoTVNlt0mB/fHu60806k/NhiDCQVSmzyTQaz4rETYk+Y1FHMVNrpPRFwV
FuaDqFByiO5Sg3m0YtybbswweOmXnUqEsouUGjYDkbGTe9yL+TwQv6sE6Yd5
Jy8NjnvIZFBgG/eSiPSXXXqGf6DJ8bHVeKzQLDKqp6ECDXC3rxa84P/Mou90
ejm6tGqLevrCU0Sk2B3dcmaCopHZWY7ca0MWQkSpC8GZWxt7otzXBYpmvuzR
3jAvFIYZMkh3ZVuwQMIYI7ocC28ymkD7XYBLnbhuOIP72W/VYt2uCj5rUKZx
cWTICTcF8oN0x+WhHWIX659hggQtchJ+EexujNolwofntaDfms5Zi4NBZETI
XKDfdVzszO0426/6Nrn1Ak/aGbzUcfawsiHHO4wMuEZRGLcu9Sl1szmPfmXG
KEis0HR6j1ST3SV6jUhSfi9HWqdFZQW+rHebTQJUMpaLjpWOUVWpIgnRC9kn
Wq59b5p2AgXn1h1ONIz4pSgHC+Mh2I081NpjftEdrjLAk/EKzs+bPNt3aPYn
xAs338XZOjtbbsM8Jz+42idQCMG5TtspCxHSmaOl6Pg2mOLqj03ea2zelljY
vNJAsW/1lCYtmMSWbwFjDAGeUWPnJz8bKzNSlx4ObP46ZBpYxeWyKX7YoFWN
TnAg/ABpjqWaYvfKqrAPiHGln7Jg6T+LluXGPUK+N7ttaNuiMJDh83Knj3jI
9tJt9Q08+sUYDb+uICD5TeDIm1U44IK+ScW9QH6l62j3ArfLgpmTHsIPeXeU
fD0i23AAC4Ny879A01sjvMOWeEOg0kT+B/VUvo/8OZoZA/bHV/lZtK5LV9bo
UwcM/1wbafDw1vNSRUOE6kLJGl2hSEOhNZxDzo93nSvCX5tBuivaHCH0Bgwd
ab7e4vzgZVSuxHT09xxt/ivpr43TRxpXWdRaJ0/1VeeL3QYCMmKcEi89O9tK
7+yJaspf6Hc7Brfmnu7dgFWJPFF2Gic2cVq/IACsKjFa2fiHjedVup7C4tMZ
hzcE5NuClhmUPenHJMTvfxCvdH9yMjweYSkmrMMv0Rqt0KxaK/K0o/Rq4ONz
jSWQDdWgdKLjDu+UaBmEcAo45EXLoTeF+gg4hlAYVbKBW3Eew+qzQUzch60q
X49T2IbzP2ogBFF2rxzslIeostuKhRrVF1CTwRYgPWpox98hd3Gq0pzGllYJ
4ToEMtsp4HwgXpusZeN/g64KfblCw0PJ1q6EqKnlYBvz4KlzPtlOQXXyYDeL
Ng2r2/UXm4kcITdynpu1HHDTVGJyHP28zuUkR3hDS2tt/OlVP8SRrnDQzJyo
bvD5RBeZbduph6nDnjPJyUacVygcKdD3dSlDb65PLXb6IjtReXYoq/YZ/t2M
PAaGfp/lgLStMRGgJGuY40rgdsd3Qdlrj392W4l4dGE3baOGjEqhUf8FNwLM
C7YhSIMHdvuHwIqkpWF5CnnYQTVW9rV9zhYi7UlBNwDvBA5N8n5nJdh34TUL
iTVWoE32HH1YcMohK2GMIpHEhkLPt/4QYSR1fWLOSfPJ3iw9GGn4ZhLwIjNd
VlxUTCPNLWwpnis2+ylwrCI5utd61aDEUA7qsagK79fjuvHX6FD4zEfiSCki
VNa3frLsZnstkCN+gWRlZ3KoX25O8nTI1r7A7xBbCv70CBX+KCrEj7N3yxXL
Brhy4PXrXdd6Jl9la/mV5Cs+o8SvBnbrsaH0VQFYv7ZDAia9zqVohaC8k+Us
mBDy9MXyJGXSiYiXr67VAf/cKBq8DXibKPWmSJ1ui//Y4rAjeuSpnRXy9Ndf
jjQqwzscqQaOKYJSe9iiz8O3MCwRgpQRvU9LiwbzR8HtAP7x/GDne1PvzplC
mJ3zkybQ/dWCJTVXSCbskXIBhlqmyppaCaX4OYpK5Fjm4GZPXsjytGbFVYPw
C0hA1bC8xnyaA9WuGxISpcQHwJ2ywAzvvq2y/ejpx3rEse3FzojOedpw6lcA
iGhBhh9gJjTXBlvybUjtpGIPTsRFC4NxuTZQLJdAkUDLT/xXEyi6WJKVjTE0
KP3agXkndIRvIx7+8h9Iy4ZUzNTFqZd4LyfeEuM0LGt/PeL0RZv7UpV/M4mj
zTGwJrNhJojrOtcAiARDM+11TtIzj1TTf7ZtmTH+F8kc5JIO4LA1ENDqB9Mi
atmso5nHQUzUZRQDnHzh3igE0hvOhvW3iohCvhjGtDcQ+tHCGV1o1giw2d2y
XEsLrVhCtgWrcPnIWnqECriVBAqDwZwrTBYkpfmRBh48+Y5BQMXlhey9Kxrb
BsVU7T/yqk/reXOtPm/XEWcEunK+ZsHcHATsGY9sbNpiiffUyjh9PLP7PTGi
t1oQ0+Z/pDpomkNrBZohf9k5w4F+rtGjnt5J8a5UCo0TgacxIgVh2JjBU6tZ
X2QAgwl2q4R6WuvRfrleUQBX9kvboha0xDeLVZWKnvrLvu83iQuPS1F8bRrv
z6yLUHNCjB9Q1oeEQB8zARzGFUGCN7OzKoV4MNKXRSkCSFFdQ9D5yHCpoFFk
t8CveIy/GtSzjcJjl6se0w/Rbl6F/CACBVyP9HP6wbol5q7hEwvw6Jzont2h
DUOXDHqxA/HoQi7kNPq1X13k/l9HkgCOhSSyWZJ0A0LoLI2Wx6iImObM5z1f
mJNDh3L2xgoeD/kLccMuArTDMZMyaZOlSZwLqbvQMyURGRSKGLtK9Pi8bTLJ
cb0c2ALL2WewUb3KcnMSMfi/+qSydyCtI+fjaolQQFroA/1l3s0Liv/MDNmY
43DV0xvXq8PSFwOHnXb2NCYu0iyMsUjwQ8EPseDjLOOej/b+QTlrtcWdHG3b
Y/k1w7xKd+dK4EKI/EI52+GwYdgBwowJ47WGLjVK7in4eeZmi1h9twYVUeWj
CSJRHGfFGpilqsj6srogHXVqFywCpPPeirovE/mqinSDGb6KUEMR4+8NVtb8
0BbFS3o+RIYVfAOXIDXHDn8rugcLpEEZxAs3IRqkz1AFRbrHzqKnXPQk8KxM
idGvkcmw1Vpaud5odQFpi9wFdlgXjyavWBB6BHYUAqVAKl/JbYN+hs+ZT/JR
iOhFACF10ErgOetYxqGZe4decTTZmUcts92D+ZA63K1hRE4wAAprmyxqqa04
mjTfyQETd9r5lopvdpe/DPD8ssWfSTOYqdg5zLsH1ud3UowWvf3/ExXbiSl9
ug/fihawFlSxCYYPviMgxyhiCAGCzcFnGC0iBbpfFeVZsL/vaF6T7KU09MTi
thOdILWcWnJz6VXR+bKlEIOZW568PnVZJuF5IRlHSm1DtmGrsd1MtP36z2VG
30skosZgnqCpQRg49fCG2BnXTHmp0bTcl0eHmnyiAlMsAm/Anr9Im6eXT3ID
//8p8Wgq6dvjhqV4laUZPu+78CPw+yeJw7GJekYVzbS6MKY1Xc1XmSJL9AXS
HvVIT/i9WQfMr/rheoPjIW21+9txJcH72PFxu+2kZZHcNV5ssSV20qPs6ylE
1YTHeBacXxE8s+ap5Mf+G+Bg0GlsD5+0kc5vS0pnpS4G6jJ1vYkYt6sUjxO/
E9j64HOI0y6Cv3ksS6IG3kT40z+1EIFOLp8TjEAm4MJPy7Up4ywgJwJmdfQz
hCx58TwDQeriUyHQCuwXrT4MGc03DWLa7ChkHTuefZdu68sG8xVXiPQkYP4j
X9xRQmTaWO+fX+ur3LhnrANn33mdtswDJNMFQYhzFw7vbPmCyxthsA4eRJjF
Lg20aK+m+0snRi13/QhAX+5JHuDwK8glSzYmTU6G2ZES8oIhEeHhAjIXG01f
lUUaEmRF2f8cp+96C9D6+v+ghruq+zaN+YeIu079PYo33eBDvPtNq6Ja8LVn
/2rYbo5aemyUK2IjLr1Bv/7JwOJFXJlrszX7zl2GIO+vYXyG052nDvaa8KEx
cQvPEvOzCNw8DSenE5dHGIgFyelpa8r8sxtui1rZxaQn7L0FA5ZDkbAoXp68
6lkVZTYV6eBlXpM/nJnty1pAhpPdTlKVIakIIDG2g4NhufZ9VrP9NINMhQAD
bqEgurSRvCvTF+2qx/QZ93SAFhrkAR4KkKBPLKbeUOCaT6y2cZCAq5mdCKG4
HWft4ir4MoIyXVDs2m2VOwl0X3y/+9K0xxDdUmaWyhdAitPoFF04abte5lzj
6z3f5Y8Cd8cNjPvQSPCvLdoFW6ieGwZkB+p+UbQVfPiFeogpj+7qmc2GSa1/
8J7ofN6P+uKPho7Z4rNouebJDrUPXgDrSN8hQt2hPT1G+0hjGFWQM7ZtA41b
ZNFGcxUsac1pfELIbTz3/OZLCsZnRKgGG3hRf7OqpFu8WOdiLECm9yTJ3tMu
J6B16h8aWlycYrhhCgNwoBmIGCABLiZe5iQv7Wil/F4iBewGOFmQETrsBrio
bkGr7MxMceBEiyRbAuFWss58c46oA6VV9nBRUXLKSajempLg9c4lsw8o8ENG
4RxMwKqQ+Mj0bOZqe/SkrpwYyaKpR+SRrRrfESHrSeQOKeU3VAndBphx96Eo
Cv3qeW+2a0s3GFzSzgVgRrfcdTwBin1ssuo2poBA+zqxJ1egs5qx7r0ATiMC
I5BLp49+dUM3P9OGw1Z9XlU7+faCxKCEotpQ5ONOLo7o2hAri74a+VXbnI8I
Rp92pL0rmt4zT9gBts5yY0+ZYpvCxxpmuJAPGUcsuSWHCankdI+SajjFSDKX
7Fnf4lfVYj8nAJyVMYLKdHncpvGdBAe4aTDw4nT3Jh5GeouDUJ43uW75lESn
Co9h8DdzrblIf4insI3TYdMXzEH4MFjt99iYRhneVlK72VYlU1ii9SD1RBzK
Q+rxXED0kA4/WL/aSknDFwXDrNK0Ohcu7d6z2tnFUc5mhnohsLXiH60G0l9Z
CMShtbW6HLOpcXOzj2UGpDmohB34NvyC7hIfuDrKWjVE7MJaQElwO8DBnDRZ
oiohIo/UnFgaqqoNMDs9GmD4sWvn9eWUZxLW9QbP3f12KR0eIyWiauQcXaJq
H4jC/3DT25mfRmzocnX41Qj6FQNPUWc6xZndqxhrLBZXoeh4ByAf/30fnBAT
JYWQVB90Js1u93h3SiZQXPqTdc4pXk1vx6QgkcN2j+fXgP7PzfbzeaePQg+v
mYiXU5w4zU4PrSLv9XLerQNN6zlmMzN9hPsw1DwZdwhBdtHfhBD/k5hGe/vU
AjgwqdQ4Thp5oW9VpwktbQR/oV53gBFygP85LjZNlZ6uCAGBf+Xm0PBJI6X/
UTMpYHKCnzicMlSofNxnrixO+pM0krA6ATUM1TnNPGdecUXTH4z1D/ZFma2H
vHa9kzneR698LT/YBlPyi7i2HtAV31u5NcWUCDkfnTyQmjLkK7AjQNWW0w4S
kLPtmMJcd0qKYN9uoaisiwWj2Bdmkt2bxxEE1sa+PfzbjmkieQToSakV6LXs
C89OvR26TtRTa/VyM1ZVx/fKn7c2V90S25hSvSt7DKgHrrscr6RK5ndVm3dc
XCG+a95g546FxxutFTq0/be/YKzgKT6D85h6m3dFmOuOHNXi9vRXBARg5Xi4
JDm2cYIHFvqM/YbkTSOtHMHbkEIZLSNtEL714T0ZNJuxG8u29g+d4G7cOjjU
lIlepa+OqZMGOQpMxjJ7pe+5r/K6TIdfWJ0yTMWFflFELTJkPlWyh/fTszYo
jysTTS6xZc6CzE6vSFn9Ek7CPC2ELTaKZAT77YAA0xiqzYxI/Py4NaO4+sfm
0EOv/SxxutfgfoSTEq6dMj2YdOuPD55Jsi4wjE6b6NimOqN6c0erSOA0Z4Yk
d8GhkQaEUSIswRCK6xiODC0m5AxBa8OJZLR39BjP/6o4M0CM24driLEZ6loc
zKHC+SEhd5e3VX5WKkjyz/0ACGcDiaPPTGLt9X+OO78XEL5bU36VnwWGn6rc
I0fCAiLpaxlVzHjOQtncw3UMvY/OqavQQaRKjsGLJBflPyMZv5yh2/AcswwB
3eAzeLPFkLk1BdpBWPlJaU3cniPZzTs+lwhXvHULM1lVjie2dXUoj/waiv9O
2TyD+ibDbBiQr80X2TENISGqBFqUgI5zXfv+G1L9j/F/HTJu0PbY65jTw7a5
FUsBCAqLBzbsMQHY0l7cX5Ra3Evg+SHiDT7EF4gU7tk4Qiu7vL1G1lu9xlF4
hlZoYEJC0jBP36m27FlbHKRQV9crrldPZL1iTvSIfPP3mYW2SvHQ8HhABGA9
UrrOGw3oTFurrLAYuuZKzjes3/QWsAgORO0SxH8ZD8z44v/ogYnP8D3oBQm3
1RuSwF9piWz+S1U51nqEaFC42DA9ma1VIgJJIOZqB2kjiblkr+GDCusdr+gK
WaA2/r57xZMQTZJKaX72VpU8AabPVt7b/ChXTULZeEYPLKc5BtqmJq6mlU5C
skrUWuWuysreBbkyEbcXll4Tx7SnG/YfgReOPnhDylkkGvvCd/YAmdWNsTLk
uFlZhz3sWc861aAx3Wcz6zyiVFuPQW5u9fGSpwHtg6Yt9i13m93ZI8Usrahz
bmJG8ZW7OueZpJnC0xhlMG8wS9hprMzDJmEXcB21SgXfP3z8NFGhtfUJ3+MJ
Jbe9q+5YIeQ56aUArkyu+MX54rn0JbD7gTPpQJYe9r50H/eCVvxSk5EIhCM7
yGJEb+xmZmFNN+thEgImsFIDuhHKksDc6xqx3IcNeKrj7Bn/CssaZsmhoYEa
0ZQ1ZCZprplt/8nQmAFMj/FSFH5Z0x5h7wD82lVe0ydWUANVmhZcwAIvDDO4
jl3TxSW3RT3kesJApBqlDLhEBhoyYw7exN/m7m69Y0PfIqPFDiQUd8IztiVP
ESCXNFARyNC9mL7aZ/Oii9rS9xDdHdfXh9aDxZNl+m/v0PbvwGca2Fbc7Liy
pGciIwyLT8ezDmilKogYx5Y3y3VovNpv2n61xKA1x1CJ37US0ekV2ZQBf7Fz
X+ttezyLQRt0YHgcgbXodyJWtFMW2+p9J+c6RCDP2shS3dHAmvmleGCPm4Hf
MhljvYzBbHyN+smGz4gFfCTCoeK7AdHLpECYU0W46MGW1bI5QAO8Xqvf2ACq
HDwYEx+hB0KSL4EGKHRNvSA303Mi+mhYtp9kaj/jm4/eBW7X+QaAlUKQ91U7
H1QOw3LyCX6nFgAhhIAWVbjEYvFlH8LNSjqQ2TP/a/NzHaK8VSzxxQyBRfnA
c0zz0LH+UihHJVjin2QYlOYbyVuaTyDfqQcGjg0S2do1XW4ku2Ax/eBaehol
/Rtbg19w0Oz4bjQD6/KG4htRKyf6y4G5YqNsLOA59bqJP8USU2qa0f2gK//G
Na8ApOx4a3ZKQgR9qRZ/Q88onnnPCITce/5Cr6jLHEWHi/DePhEnT2HFOfqI
cSLTIh7IAZudjNWvKJk9bUGhqZvDkvCnPGox/s975Br+db8FfbRwfTKhuQOV
FlHvMTfd2rVNA8VLcRY1RvzUtFpbf4ckRrjWqI2GXW1NfFOxtnXX5QHEGf2h
GlWszLU4uJBrihV/LlkFEctp8crY6KJ8Oda5sN5U8wvcfQPNvwgNOwOX7nEn
MHSvz3Cuu6if8Jwdfi9IeOx5L0m4EdHfJEw6Yhrjvq+ZitY6DRfS4cHY8sNS
htE4k1jh9s0XGiXB+apluV8xXO2mJln3IiZMeWTarpgyYJBnF24KdkfZYyq0
jI6QMpg7u/Q9y0noE95VYjVCQyS95ZSNgVXtBGhFY02D8BH7oVK98U7/jn2E
62X36C7or+3Vrry6D6+QayNqquxuMmaaW6Gm7v0Og1v26SWOPm2dwYE85bGr
x/P6rIlYSXz3z1qKoNrpTvQIg5KPYv7uPLRqf1f7gR68na06wLRwc1gxK0Cq
DKcKH88Fl0yTWXI+J1vNxtdXnqRrKYJZuRcdkIc8Lu3bL473PHdp4TlqBqEV
Q3CBtF5Aj8iiRB/p8a+b/LXTrRwUNurfgw5zsLxsSQdqXlu0xuEPdgXoAd5t
WH87g5SDBfGDTY+p1SwXg5nCyeMH83dzQBNl3M1uw4AjfeHgxB2AV7FJPQOL
BK+g56qy9t6eZcSCLxKcM+9ejFztyQzzjdCqEn8jr1NT1Z+kjn/+wr24Cpkg
acgENMyyhrP6mXVViDdvvMXv73B/Ynyo40Euq0lPFk8rpe2fRxFY/S54vq2x
yJnxTmJu5yPMYfEFElmU5Tuzj5ujtd7nO/UNMz2q3shjmbir54+6rn9Ycpm7
OrvJyn1VNPtqqY3e5PidCU8RWFtGuq1FUTuzDoPKQKoQfvp3ZGNcZSpY7umT
o+4fz7ZgOANRIUI/prAncKZzM6QQwkRnq/w3ZLIB84nYfbmhtlb5Yaurb+QE
vUqj8jCx5QSvF+/QioO90efzJQPvoDof3OHBhEUVId8cGxDPPkDHXK6MHgn6
X/HWQerK6IZEx5f493hhhvhA2Yr7/xkp/VoKvo+xQsZf6tKsiy01HeGDcg8t
w/jBQOTc6aO5MsiTpExV4yaN3tcAoV41TfZbjObeHeT1H92SwF5D2SH93UIU
9mHaGffBOCeLiNk8j76iJfPSp7lBxtSw76Lue83mgvrW+u8rPQZTumPTZlYC
1tf+Hixh/nGGo2QcfBVCWIMiaHjdFzonorO2m0KSIdU+/iyGIgQhr9UIM2Vn
0RksMzNdqBz+NTaN44QD63NCjksRzsOYcuy08RVb5wesCF9z3kzzXM7jlloo
zGY2Z1znr8SAvQne60V+M8P3PnCqfo6M+OBPLamg321iCNW8rhAP0Xt8MEBr
rqS2a5zrez2r4LCX/QAGEwgZDOj6xMKsaG4sPe/QnmxCPZfxegtD+ydN55Rp
Ty4E9wROTF1UcGFjcNgeb9EfbOzaU7Udy8jnttF5wx832CyMYgR5ejwBJm8C
bxBAdJIXySmWSz2QUXxAxHyKha0SmkiD2sqJUfguXiCagKZw0W7LuKWsFemR
QI1JHmMQFdRHMnpHWtkf3J34Zm7HoCXASaWoIvc/+tH8YMxMyknsUALI6r92
LwM5Thjbq1Up8dSyFHZDi4E31CdSbqIigfDXObQEyWVH7zwOkzYFb2lz+I5i
o7jpka4r+msKobffE1cSMMS4FNuZwAgQyoVx1HDzQLD6ylyUUGntsM4zqxb5
HulgUBa674Q6s5RZfu+620rKCgWpl0KNy1la/BtdSO35o+LdjGk4T+kWESo2
DYzgS6yQGzh6esLm8jvMDFhB8QcYFfR032gSSckgP9er8ZdbOzwBreszirg2
HQIRI7Aun4kgG6SFXkUHjnWWY81pCw71K2aDDQtLr+wCXbb/CQvYtjrcC2AT
dVNJUe6AHU2eMDwZkqCQammV+NlrW/MvrsuFCGKt9gwoCNI0gTRmk10hlQ9+
2YmSdGZmv/MpKxQU95AL5H2AdYHOWUsoaFqUxRRDBoC/2PdBooqFkA6OZC+y
4o3gEV9us7u4z4NyTBGHwQ4mLl3tsl9faWhJ+6l7gahvXRSHOaFJsgFD1rxS
x7XJUaM1YeF0qevKkwbq3iOBBPxGSbpHlxGBd6nELNw9AS8sCHHaWd15ett8
T3oP7PHFtOovxuBwvxnwUlQxuFrKx41D/Fr347raekHswizoWSIbDz7vyUgN
Ux1kL2V/eLYB71ITz30bFC6jkDOyF8OFoBy6/VoLopQkNssmsCnpQL5k0m0r
kZ/mZihzSnup2U1Uc3yqE6nHaiYySq61h5lzlAgfFk2JUiCHbRyS35+xqFEI
w1OvyttFtsHAqrq7Z2eBnxUs/+SuFnWc719NRW+Qr1Ezigu+zHnG85r0h0hI
ek5IzqlL6PNZxcpLvXuCKm9u8Q1bFAef9Lr1OkdZVmsklgVliV/gseyaEGQ0
6PHDZ8ESKVH6iiUHw1RUee9IxD7D6RPBnRJCBqkcs2/pZySve/9/jPjWVwJ4
CoSsLfVp6SIJ7tTzbJf76rHGEHlQaod5HoqvmAaanHKlpB72Xq4+ndAoP2vn
MraHu9CAtfjJmKeFjj7SBuPnUlLWtsBcQzar3jlpPQfump/zecrbvGuU5LKs
yClec83RgJm6n4C9+Z1P6qspBBsfPzXVuUM2AupoD3nQeECtPFv2hbTDxYXa
sDxlpkT6eu1s433Tx8Q+pjfeNoCpTEF+zCNMdCCLvahHG8FUVjMQosNllIeM
hLVEMnPzii9pAmHG9c88fR6Wdj8aZ7UO9j5Qso7vDE+pMCrNnO82wAsLKxfJ
34jgc+NQE7EmguG7Qzpy6Jv82ROPIK3hbGFXmGqtbnOMHcxN1Km2rdjyzriS
iQpPofd16Ic/Xu1xrVurIBKojeCAry+e1m1HabrRBXONaZrkyWRwoJw3dRlM
Hn3p+NwVR5NhXMsz1FB3zjNcoqZjQ8DGKHBt6MOr/GSSLVNPgAi4ISD/iMy5
O+dnfAcTYJtES2X2PpImPsc4QqprSJg6wNP3zUG9nIX8F02TlkQztEAzJrM0
THIy0CIsbk3Px5fZ1DwwoB3EtikugVjF69kbpyP2neGm5TR5UMvcqSnYptTH
P8brQf8LrtCAjiTfz4kTcWdFhRbrnCIfFDDTEl4HmgAH7tz1YdU6Y77tX4RV
LGNym3ZY4ZPfkZgysEFoWKUFfaYU3d+X5Rc+mw70YxiL0xFowiOCGEv23XAu
cvjGWSPWWpizhcTzJck0mwFKDrxd3DcDEuhPsLQTgeWZHu3K9UXPJmHCpqNL
kjMqAReUtK8BQdnSbyMo2wHPox2oygFXkBIA+VtlJdnldXGovO5Z+P+/AgkH
5IG0mrYQDcbqIpLkwxJXYKP6tYYIj0ZSER42+Ruo42D5QRkzqPyArnlo6owJ
VXTE56dElMxpy2KTIvhZDy2K68ejrX+606TMragF42d4SsutWRmbww7N+yEv
XRl6zHU9aKUldn6WcU2rZahZ+tfYCAWft6olY289maAzT77NBvWmQg3P89qm
kxvjFpX9KUsP6zSTt+cFFmkvp6VwK0BbnQHPCk5crInA4Ju7oTavUL0wnFVW
cqoFpn6MCdGiaY4pJ98fMuZ4NvwCBnIG0J/ibvvWwaOP1gLKcX4VkZO0SYJj
c5Ybq4wr1znVZx42eCzEPmObHkHzaQXW7ERnHRf7zwnW8xbKch/vTLLe2g7q
ohDIB67fIakvpZaIog0TRhJ5IMffhsRhkCNfqoJcKbWHTJeHiJU7Of8/lD39
NRL2GG+pclZyJ1LvEZQl7bvxiDbK8KBBKJfShcmQP0h1F51f3G5W2StYkD/4
Y2t3kYLN7h1+WImWU0Dor6i08K3GLG6HIPe/pxSAyn8ue+Gu8KXDOGw5gXng
uYlJJGzL9iLpGkSK87mzrcod6XFrK3zIsDIXKRpTXuIlajBWYa92xObxdK5L
G3osoEuNyFDAyhoszLPYTGjo7DUvu0IaiTEpYrXf+onOFogSoPW80TkZAEI7
o63SApjEq3r0pRKnE8sx3J0XYWgimk/Sm79q+TSt9+E6tEAu69eOrYHMOeu9
mmzM6ci01WsmxGEEsg4igU6sTgLWlNkBApGbh6Pz4CSGn4hp+nNTzW95nB2l
Xcwfa3HrsnWsKChQ/7mNcCsqABKxv/HlWEFe7Q9UwiT+LSaQ6biK4/y5yKsr
hbyJ6PQ+h8i5AbP4gt2MnIunj85LXcMi+J6WW0fV3ufFWA2EevPafHPQTaSL
fZA1dGMnAW1pd4mg3/IuhsZjeKI2J/qLjcjhK6Ho0nWHQngLwsvJqI+h5rM9
TWjfSVr749CSXf7IWDn0X/pNVWFFU/DlIzdF+x3jDmjlv1CZ5fRMyOm154Tq
jywmG3xa3sOXNAe2xd2MW9wzQ1YWIQLHbTfVYc2Ghq+qdq075ubLHwlsE4gY
RWrkdq2sonRh9uQ7SqLn732E9iS3oe9Jol7wMo6S0kHeQgx2FfY840rkAel+
o1jMEMo+OyBtpk0QaljU6J32slnzOv8tDKQwTrlyzNf2DMJwFpjxt1BvZb8Q
TB+ismALe3vY8CO+hyW7Wj7MgjRNH03TgB76uGOYfmoSc85xigum4QJAL12p
/dOm1TczrR+d+s+JaxjQuHVgnYR4m7AA9NSTWTA0Tv8lhpIloPyxy68+Vpbg
nQo+mIDglQLj+o2xKlVHBjz5I4BLEonyEmMXuu/fXldD0Vjg7g+pqKSpnYkW
QZCPmGXWt9l/yKCCp/WqAxRJM6LmvCdqAD3+9yOi8Kaz7uTPJKRw++MKL4HK
3dXMZqIsAxVxTMnzfdJc56Ed+sJqNtWxkVaOjAtvpZzLS8luxr/OIy9V4luN
D7exdCaf5I1THA2tcg4LhGefBi4wgruo8N8YECBbtRuuNIuwjvRSsY3PPxt2
MZa5PrSCy1XyjlZheN2cpmdDPBnNqeVnOoCo3RbDZhihHemBTAMx+Z2cu8Vi
NXEg/1KL1zBM2FVGOMDQtmhAWMyLnjiK9nrRyluw6BFC6XXLo8otuU90QP+j
Fx+o1XNcjB2Ff7BfiYJ0HkObhLHDCKxchEydpdY5BRDxYqOP6jgVyK/9HvuH
17LYIJqAtkwcoLRdtj6oSVXfUdgXG8VGWuzmaxlPjRQEwgg6hNewCfN4ZaGi
vIf3KoL+uX665XB6AGAGlfqzMl700A1YIFTZzM5yRVZQgqexXdyns5X6QgeD
GGp0126MRmFUJaKG86DDzNUALIl5uuwe9hKjmnks4rF9xdKAxaWONnknG9zO
LpxWUye6rQuDXApxkiOxF23BHAMqVVdnAk12OonrbxlfU7WNWzZRK5J/vtpw
PeLtHCbqtpRlMo0oKy5qe97U8lsiBwp6DP9dk9l/gBZMuQNiKMbhhy4e2Bv/
Pay3v+UWo5BYiYzma2bs1vDi702hDWk8mUmM11LNWKt08fx7GW476tTfCyqX
UY8yE16eH8/zvElGwC2hjicJbW0RW9Q82EKPckeUEq9lwUSstvaWk8onAQFF
tg7BPXId4BogN+d250IeKNdmLmqPATzdpSYKVX9tA44oevGXL3pEEsrtIRL1
py7Hc1XrC4rjFI4gLTcxYI9p/n5zzBbbXtBODSK0sXVn0+H4mwUAdu3E4MmN
Ku/SPajjpqMZ8lpz1wL/Rc2KBPp3Mw0tTaMXyd+CtcvDWDWy8zvr43g3YmqQ
jSV1XvOJxB85OqVd4xURAIqcHRqLRkG/q7rLIZLC9GRRVUcxQ/7HnbO0/9yQ
lCFvwy/CtA84Ktti/n2vaLvmsKKiOU6lTDLeAq/ydF53lLon33Vn89Ti4OXE
bDfc5c/rVHCysNz5la+KR9y9b4YEG3KxwnkF1f47e7dnjUBjHHnlkbuIBtgm
L8Go7RS/k0DYx7Vy2efypePGWti/WMiOWFp8jUT7DziAlE/9CK9uS5/egcAk
6RTDsghjrAjzHzQ/mNUK9YbGub1ccicS1ewgPKV6R88inJSAuLbdw+MT9Dop
ft46B1nJ2zoSOXpi21UMeczaY0HcMkbjR1XreqeWR9OOW26WEG4BKBhdLWup
lc4dASAA2U4GfFgeZgZgOLVkyXUDKu0MJkOS+Yx30pdDt4vDPsScHcEC4HZy
p1D9E2oFXCAQYR+KPsZpB0ZbaSB8q8/awvLANDy6qRi3Prftveur+WsOEiwL
NZSGEY3TK/96uu89o5zbNiiiuuW9YZ64c2ebx+AyWb3S6OiKRGaNHl27z0/K
KVONm0UkZAJ4jcHvCPmUfWm3QPrmEG7fILzYoABU/mGz7Zc/PRnneJaQvE1A
c6g7UouX5C9sS1+3AgOWtgXuTKp8yS8TJlX8KkKykfVww5G95Y/459AvCe1W
lekl+9RBOBG0P6bQJ9XqItBqs/NEfufx4jbKZZptonjF8IyIXLP7MQRZRPyk
ROx7TwzHPEjoDqiSVr1tmf6wj5NLDtB7jomkL4v4cW8sW2jGiDYrXUo8L4d7
H7bn+USAxu5yhF8r2Zf/rXsTW1hOIxbxj5vPm1Uc/KycRyC909t68tebnwc6
dnXDpluwjxQ5SpuzMoVmkA36SasctYlSXt/zo78nY4/98qXAXXZs4SFhuI7Q
+Llky0EaY/oUIA9tKQod83G3v9umezdVCiywUxZ/Y7Ta3N8bQnxz+ckTOJ47
SoisOYmhSHkgkHPDZlCfNNBgzDxtD6BKCeaSuQb362fepDnp/JiOXdN2gu2O
5Sb1MrzOvIwA4Zn3rDMtbuMB+Mqc902sKLE0I5PfZC+8mQRFlK2hAj8DrIY0
lr4fagQ7wKyk7XoReHQ9yO00Gj8g19EEZSNMu554JTEqZ5pX+3cisCZxfZ2h
zXOvDTvThiIT+FuFNw7L06MdtZ8SrVZkW0/nRk0QeDlxzqRwBwzMFpVkKQ4C
930i50dmdtBPneFQ6tljhD2aIf+SoxFj72yCF9K/xAtLZClQ1DkrGCe+KG4v
UXcRpqKEzfNZQ+fg58xNzIUCPtkvMBlgBKqxjzCKM44/1CYXWB1xVUeamZzg
xSUUECqBaN757O160LVBooogjnhEEmRnWqRXRYwbZC2nEFiXDRWhKjHz6DRs
FtULtCtpr87qWVfY47/1UlM8kezpQqP0SnryGKX5TZFQlGTZ0LHCtpxOgwhT
bHBkRMn/0lXr5+qtzRsYmPX6t/gJ4uln88N+InQ1rdrgFAfeV1I6zFXC4+cE
HsJ5GUR03y6r2cBKXFCmzB89uGisCiwcJ8H0LedaNBgjuqIGoumQB1em41A2
ENTkpSXsDPCdVoLw4S2r36+A4rBbcBge9XySsOCZSrTiAZIpmn34KOJ95uO2
5Fzmt76x5+9oAppxxknzw+IS1Raj77oCsca1cARgaoAjFu4r/9hYxOV492fQ
kThKiswsY7Rl7/BV9NW7VaXoqquPIwfe/DvyKEE/LNwaub6VpxubwU8w4iL6
A0ZCL5ZIDyJ/70DYPzEAGlX9/h5LEhshPY0cimub+WBwZb96bYuxwJTu8kKK
tgiUfxGrIpCouMx9UG8bd+UOu2APL+cvuf8SU6vqhMvMj4rDuGzlrbaWJUYY
QHDfdjzmoMPHCOoOko1tHsHnRSWOjhk4IyEZcRpdafVriOSUIjYBW+sahpft
9M4tpDsvW6qrIjRVzbjWTc1KeQWG7j0OhIF70CVKK7SVUxe03Vxj0aKOoMoI
y3Q3o7CCyiBn30upSEtIsmf8+U/iXMj/fnaK7jIja1lW/Zs1O088vDMT+wLN
EaF6kNct0h2TJ/khe3aVTaXwn/WjNrjSU3P85EFM1WrU8gK1Q1i/qBGuc2iy
dm0wUY6Tgx1+2OaP1CGOE0XWGrwc4JnDPATV57qTVf7GcWOkEEZIwfzApDd4
67IVrxwZkpNmVZnbbapuR4XAgp45JOsHhOrOwGxDirQzhMBjQ3q+BuZseDIM
eA1vxZNUp5FCTaKY6ewP5MqT7LKmywBoGfS41BiOEfJBxQtCeCDlKFKLuBNt
6zLexH6E5NS29uuby2xG/S4pRCM4AFE9i/USzdSvx/FXs+zXJevwutZy7Wnd
7ax9YwRhjP4Wag0AVuYmAuqydQaaiUCHlWmj7gYGvgE2ulPL3LBk6WRooHbJ
gpp/Ylm4fEFYEHrih88FhwVkfXZcphoqRCt86ffXDBnqXQ/Drag6pKYRWmYc
A+0dTQ9aVx25jWDPGa51rTYi5xcRVz7pOMwWm6ZY9+9ehaCffHGMYTwLc9H+
0UMm0DcJeHN+Kr7PbHX9wa8INlkKLFaIhcWeyttd6HhqNK8yi1LSjJ2CB1T+
/pCagVLDGrvw6eEcNdVWhbi1fNIhyKN/19gOu8rxAwv+M3Q696FsNZooK9cG
pWjDv2/e7xRP3hYUu3qNf/Yu3Uto7txriWkFxKBsbZ9MgVB2t1nbrcRHjV29
7fZ/rgvZu++XdPnt3WUDzXwI2qnIfONxOKxmMu7RXTSUnOVvuE/NY/wZA3CA
6U254EWC0hKRPXSbpnX4XOuBGYmLTb4czgux5zozRXV4zErmNRNQxMJBEkwb
ieWbxnyDtoApBKX6gSYOw0ykk1Vrn5pvJzRh+bchwjEDGKifTEHGnnh/hidQ
ty7cjRS9Le8CLgmtjX91OIgWHnI4UBFYHqnrW2ezjey/flT+umSx3V0FgtU+
WeypZScn0NvfiqjCeGqa6vr2kJOVEytzkAsS0CydWb1HDDKC5WABwJRpn5fs
xTjW7NnEdA7lOehm8gr+RVFsqM53Qn5iCTNeGYr1c0OcqI91fQXDfMMMnyyF
rK4lt8hrqtqZeILfHIG2PoG3e+jh2lwuMMUY7/+nnzLlKbrOAxwTRa9StUlH
8E/Uqa4o4Ynryfry+cdBjOXFOsGhq7ADzaUzFypYl1luXYNxPDfIXPea0miG
KsU2N82d/AoIjQBFvi9L8gAlhTnO0E0dZBcQl+OKc9XQLhOqkEZvsdbJMQwI
oG98n9v/1DQU/DysltMfUULXPjhK0jWJn+YnCO7o1i1uszea0y79jExzcsas
mzmS2JpQymsqMVIU0cZFNJ/oKBg/CDL4BmlAHM6qOy3Nw1WU3BA4ucY4Bhxu
cdeGfAxR8FAbWn1o11woOFmUAhTRpPCulPr+U5dqKlTFrF+xTWWhAcSd94l2
dPdU51g+Eo4hS4+tkEnNPM4B18WRibQyzb6bCWGl2jWE54P39+SjZ8P1GmIb
0DBEL2Ah078sbOPbNDdGlNqeX2tIJ86AGpZKQDB+NKxF2n7SMq4nRWkTwhUR
EkGbwOJ2EuV6Bd7Surqk7KmzD2nVcMovt4avdsEA+XDquZKf9p4HlOPOt0iE
nRVJj4aQ32G9LkDCW3bMb2xDC1DtPqgAAMn7hYyDsX8YOOoNgoRbrUeccRG9
B+LOE0PgzTao4FIRd0wuCUc4dAmOP5gBk2HSIaZoVp/aIhoSB5cFHcN0sAXU
ID461piIGivcYmOT0VDYBMN6wQwNGBTPG7s3EVyN1w6GB8Bd1YDDTRjF/OFZ
OfJS58HBSCMDyD++MiMfyu8AzetEjJCxWw5H7VMwyDyZ400Mle2XbxY2CPZr
reBxnPm9bDBPBFSL5Jf89SoCN5owQjuzgYg3Ln+NbYjQIrt9N3VvTb76yvlw
vnOAKq+25AxcMcT1pmr9wBPGSGC5Zj8exTw5+KbmYgWG1iHESTSq3nnE4Cy7
J6ga5hTgsl6uRvlPoHuuw3LkjYOH0ORlg6WPgngS08e2OjoOFx/XYObHvRMw
pCXRm+xSdeZ1581edNAxXn8J8pcAWYZKN5+IkoRzXgUOgBpiOSDuSqasbEgH
mF8xKdFYJdjKPnIZigtkLeTO4YePD0uFT60uuxpT4XhSZLFh/gj7d1Hu8YLh
sZ1akv9sUBTb8/TjsvqpzuBfNcmltWfMHwZKsYcmTaDfifK8Bbgp5saa/gSk
ltvqO1Y5SzM65jqFyTkiPFGIsxNbqJyJo3y728/OWZO9k6jfI1zvUx0rmM8k
7VAOfJdyraWjFCFwY7Fxxyh8d90W2/k6pvllNBeQH3pu8yv9QMqjJK94MXod
Z6HcegtsMNI4avns1KG+WdTu0wkbJxSDzCsgo4RaDqDwryJomc3kwurMyUuU
wM8yitD/TWDsGzO0nzVTgsICDeRZUUMkY+ok9FBpC6pvo4t38a548viDvD04
s54Iy+HNFkUHc0XwNVkZFbTtICZhnEGaWBd1GKoajMcn5YFVq3EHjkeEJBiU
Q+pz6tduohzT0SBvnO7jNFJ42B5KBJ2kxptxbxcO48Ute/+Bw5qkRjCQ2j3n
M88e44rzkk74LH7irEF9BSJwnlVyjsd/orz2+BerVBSljNojPoKNn+QZI8dJ
nLXbj0HSiqB8/hJ2rFI51g7or/260kdN7BjQy05h4bu3L4pt8FX7i7CUWvG1
8mz5zTYGGlmjYx198StDCm2NFhcGXF3SnjZwj/lwa5Z7CNZAdfPv7sOZTnyR
zqfwqzqB17rtAYV4yrfRuyrosSgtHrIyFe0lPwUKEKdBpTX5fRopree5/xXB
M+gFKDIE/9JQBAJ6N6TNjQeT/unU47CxptvTVSNvlhZaPuGY8upieyeROeg4
9hZmlhMo9KfjChttj2/uZ8QIJJQijjGcRwQ4FSqsJPdFa95aCtaBJFxD1Gha
KtFJCQBOEfzpzB7QOXfrsFJfS8CDEFrJWB7TEN4lSFSaE9jNryg+P+sRGk1o
NI4ko3iPe3JFfxYXXujzSvBLJ2LDtlF6V/3SSfPCfgFyWYVI9XWuN1+2Ro7n
i5xS1Q+egrHDmZ3b9mreztHk31ISxNPSO/Zus++nOpUeUUIJdumLEAfW9fAb
7mUV5NYDKUJKVOxgzF7cHNNMB8RTfUrbdWC/Waf12QzjI/rZfxJl5ldZNGhb
MZIeOiOz7cIQ4Pvn+VDjzt2f/HbjrDYHgRs1/wCZbfYO17209DWYtkFPqOjs
et3U8XOmFNb4cX0BD4p3m1YC7ifuIi4I3Sz9IwlgFq2XlTVsWsjkdK7zkecK
OArxsioOmt3mxEMp+leflkZm7xf/U7ZNNIccF6zTsJoqkpM1hZV+J4NEABen
W6j5NuThiPQlKsCc4ZLy+AdkKjqr6agesaihss9rUGQVZ/xsr9wdSEgWR97l
NBMVWJM+xbSuGSyfgf2R+atIaqgdx44heQdqGcgJCMLqfjf11lV9bCLDlstg
5V3xgnvMgyQ4oz/uaaNdgguFzKZX5JCZs/tANaYEbes9MaqON5mzT966H+cp
83pHliVo/T7N7Z1dIIDp6ZH7J2lcTz3chMI7mQ1EEkVuDdIKSmLY4EmdNbnl
KDGnnt41ge1HYNSAB9yDNWlOcoAU104+6wPagmd4dDJNgKIYzHhwd90G8PZx
u+UyZP7mLR2rB4UYZ/VDLPyE+NpUdLApy7lQEi4Ecaa0W2JU6bDjCxSiOIyp
vdJ1VnXMobhzpzBtC3hgIjSmbCX2c0n2Rd5DXgvrGVs58PoogIblSeGT15NH
UJBNlzQxYxFf3jd7vkfkDgqh6ZFrgPoeygcIKEdUT2/beOOJQS7NxISpapBE
nc6iLOcC6YJomu+QkOEinfztQdUkDlVdxw2aTOOxXCyMKw6DOBvGY7uy2c8r
zFYa7cu3Ug7bIydHyLaYOXiCa7SQTWBlJ4UB4NS5Qe+PzKeenzBhmVMiBCTg
gsomZ/xQ8sDr9QlCHgYkoiDeehc21NrIGl1S7snAUS/l9hiH57NF+DUqYsBJ
riIOPVH+61tNMyO0hfVZVuHPRRAakY5K4QLKsO9379aQ+sGl0nkmfD2Vuncz
8gpJPD26R9vvdhvTwqSlaaAuKEQ0LFvz8ejobOu7KNMhl4ddFJQfCvBCaEEm
+LRPBXbs6ZIbKrS5JwCc/QWrOUNshMAbvtnwz8gA4n1+E0MLJYTLyyWgvjkB
Bal2q/NFfCFiCLYSc8CfOwa+BVIPw/PpcBcCYUvYf/qfg6JvG9Sqy1OJYXN/
5pXdaY5pV66L16id4ZH6tHFqxeB6HPXawDBMgWsaOmgdFUDjiuqJixwtqClN
vymsPapN4ry6dE44ZJw/nMX+uYG9j7ceNOTuSCIgo1NNGV87HHj5DB6eO0BO
lbb+ExI7WaRk/EG+jOeDWwCUkYhItVDThWfNqJ47gszfkZQwCIgIKu+hLYua
qC9mOrMzZEzUKyD1yJDxju3t8RVkR/xSxW5+vvCbUifLln9Tj/wi/OzmjZYb
K4chanX+Yrs3VcaIr3a5fcdVn9y4I++g3hfOPw4RgynW84r1WMPoI4QR3GCt
SKwg3mHq/bZyKRmx+1VH+T1Cqbf+NgneBguireXG6tDjRp/Q6YNlTTgX3TLZ
8LZiuP83e8oRQ94jLYjj1akTvyyHaRL7ffH6EkUH1LIRY2f90aYoIh86YqE0
P8cUmhp2YXYcfj2di3HLlFBVUne+m7UYeWcibeSpn7O+Mru6a/HcdPeG3cB3
o+9U0gSAcy6Tq2CM08ampnvZPDfw5DQ7EC5O2m82jZz4cms2HmfgCet1ywfj
tCamoZ0LHya0/EAs/sVY0FsuhfEFIpqsCi96EJzv9buVJiMYFA9J4Lfj+ofZ
CzNDPy2iDeJu116fhBaEqUF+BC7j9CcJZ12KRJFCOxNYi/2bA4Q1tHh6a+Ex
L3T0I6dUSy48K2c7nS0hVl472ZIjhJBIgeDAKdLQvyp2uJz2IokcyC/aJb9w
FvRsTJB+KVrQnYnvEkNPuRuSGubm4211BpwARk+28bmKdF58UlK+FHD+StHM
zuURtgz2FQfwhNeQPD02EtIsSs4ePrC7N9QlVOXfByRCgenHnFN5AJoH5JKD
o2mhIXQij6k7C3NVd6Uy4rzmN/BmGJEnKXFPCediTB0qcGlHpM8AAReWp8Bp
iXIxFwvxwV6/sF6dQIv/3jRsisOXvuFfafq7aYLgXOMCE3V8RX+3S9NOpSfc
CewaTvozBL7BQFHQtiXmC5ZiRnj+mtdLxT/F86TVZpOVPwlJuIhO84JiN6WK
Favm4TFCSB0d0V/dZVR2oy6hF5SXe9IXJhNMEOFtYe2t6jHah25qdIBOj86W
t9sCe7YnzzKqCV/0/zXap6tXhAtaTIsxNarU2UUbmn1gWIESwSD44Op7qMZp
93HjgdwtyMCFtS1/2vge5TfuW5WvgVFAS/+T7twph+mIbnwy30FYL+ssc2pX
PJia0f7zgowRJ+r0G0wQh3L/12BtS6Mh/glURiibBvI8TFgzSe20xPpOdJhP
YIA4m7+qxXujgieHKRns4myVue9za+c+ieE/NJvsUVixDVs6Vr5DZz+14+uQ
I444rXHWBNrugYd+uD9uubs0c4cWDXM0WNekmnSjywbQHo0iTYbtuVPBpi5r
Bi7L1m3FCI/t+aeGSkqnaY6zUgxDmp9vC3b5FrzzSxhSYcBamVUWfUc3QMgU
s6t4z26ZjLGbqOKef7Gy1hCTHnaRCWTWXUnu3eMzyy4WuRmAwfKJoOQPEUcX
gy0Dlo1tH4k95PLa9S3AVQsmd6j98yegfFGj1M3f4g7cSKxxCC1j4CePGxai
/nKnJt/KyUexpGdOO9H4H1MzQThldVmukZ5xz5m3u3BQsl+AOYEn2jSUQF9V
u9WyKA1baJNhLBFu88++EGonQp5ZYQp3t27RjaBVXPf/b6cROHQGrsFTQxPt
d9o2Ziwp/58QV+/hcfD8IPvDROOS5pVUNHEWIhDfEll9n5oArp1SemqIOrps
md9HZTZIsJw82tvv6BiE6Wmxa3Re4quZDB2SteFClmfPmQ2tWlLZMyncQ9X8
DytQfMH4Iss0kmtg7ss9P0B1gsCZfDpBslpwUYL+l4dKiKAW11E2d3MjMrBC
7I+NMLcx1iIOoSaC/0vt4n6T3tMXAsKFq91WlFSF6b+b+0aT98NwTtb7ZBKv
BmGOQQgihtFi2cZ8qQqT0WIO6eHKXrgHAnRJveKzPPDaAquBdh+JzbJBFGXh
5zMGl87NcMCnjbc77TQ8K+uFFR9T8kKUMRhExToSp2rJvDiiMvQKNS5p48Z7
A7gsoQoIZWAMOhuaPqy+ESXm4XU4E8umQg7N2imHbu3CKXr9rlOf3mBtXMdF
RMT0OGMG0P6eMrcTo/vbpF9scCeRu7Zhy+loSKuEx8Riu+A2Sn4GBRyloQhI
2sIK59bFdRXtnAmj8KBTwR/IJ7raFRGethpBx10TzXEN89Fkv2VHVqx15LxH
EheWO6fs3nVsH0KPLz+CaWMHeocSS/NSpX1BauLNwRmAMxKqGBdzlFWVBq3m
MaifmOIGg01Qnx6TT9xNNB6+eCNXTfl5OxamDP+sHvmfMUC68jlJuNGNdi50
AW9YZG8q0Pk8LyZBgDozv2TkC+72m4zZgfsQ0e7UgtVC8FJt5XBc/j66/iGC
zGAD9ekPvPV8bJcLTiYW4Td5zUr6FpvZfF942Q1y+kxC3yDf06apfwkISiqC
Wj0SvhgV3iJc5tzUnRUCT0+JXiVGfUvmmdKxz7IQUSftp8tYybqxX4vUeTvD
mZNzjOf9hAhVZTADOWR3N2khWUx/FuLPasvSMbFR70TbU9M64o05yOOW8ZvV
vzFKhNqhiCzTXvfPAgABVNFrLGiR0C5iAC4voxCcvoMUrq2xw98om1n7Tmst
C+aPEoApioHqbk+O8zo9yBS1RZf1hPsrDDeycjVV2H8JNc2WxKwxjjmBCSwM
XHsfTFxJ7FiHvtSlENVXd+ra3IL6nQBxi2Xiz7u4j8++suwswzJo1lphr4A1
mauAryV3XLwKG221nM6NjxVjmn8vdCqSRTZtfSahzzNrkF+XqI+RllEqbU8p
S3wILrXsED2nnHksYy+TzUlHEq/fqXvrYRXtkmxadtrNvInMkHISNEX2Ek2b
g901M2KuCMpmjRGwWjEaQKi//zbNPxfh/zCB+XPiOSEOihAUBnygGaMy/eWr
b4miK7YfnXxgGfqapDiuXbGHrg+d7uKLiVTTBs41h00DoM+lB5VvBsKuzgX/
FmGq/wQ5yflnWqVbi4PC8qzaqkwXPVwp+lq/qB0GPwu10asxPYNV++eQq2hP
I2mA66JYoETXkUvqQgHq9bqcyC6/XIamJPF3iTklqWb16Tkc9gRPLpw5C/Rt
KbBCcdzAcrc5zK5kDWk2RozLXkWfNHgDRADPYecpr52wTcsfJlx49cVzuZKd
AOYjxm/DXS+BudIVayY4JAZrswg0ljY73SICua5CXQg7k/UPpHsF104qdPpi
gz1xEsEDTHbpI7kpCuh1gkFP16fwL82k9iaHn+7LTI8giGje+ibhjvepDzZ+
QXc/cabw1Kysy9BD8DLfBaWPtmQuh4oaqR4uq4oqP25+UHWe7jLPl489lC6+
iJr5IFj1wEx59S8qqCB9Ib374vpG6sjTiDXDkQoELZzTKNtdK5nGmv6g5Jyo
Kp4SKoqW2Nk9Y70BGLDs64sL+LcJBGmZPgNr5qW7dOGax4toO63sOrj8Mz2b
omoBi5AgHEQGb5DkEI3s5uDM9j8i+flzJJpfWxU60l8gBFN0bhqBq2a3jnhm
RBfWb6SKGaGyZa1RUwMxdXtU+2hA6TRSdRb2L7dEJkSDkJd9XmvFkCzbUUBO
b5vcFKBDMvwn1HK51voZsjo93IHUKuVrWVMnRA0o+lYPVwOdHq18oHBvT4cP
q8iCjO73XOHW0yLdjCnhOWJQmgS10wBDsseJdkyuOeV5nBSErzuFXCHD7fk2
LNM6Sa1oI3IJCUVn9L5+dlEsjNKLj5sHC001vZLVHSymJ6gqSiI8iApFcHuz
PZRWYdYRyE7bLud876K8fS6i3dU3jTTmCukjt8764heY8A7BgZx+uGSiTpyk
r1tPdZHDvfi3uNQyhgvBaTWLQ+85A+YcFhgGrVpJjCFnB9Lss8M3jagNpQ5g
Rg38aJ12wFnxzmtCJN7sUK00XyPOp+Auon6u14z5YZlaGHAXRzImgz/wDw2t
dBa7ckqhJszD3an3prOs8FjOuGm/a4ACbHGakNmWlVoLlEoQdEGtWSLgpLP2
ogl9qHqbh+3issbpRCaMdWKQT5Svzv3yuJsxBmQf4c02oUCPTIna3Eqt+zTG
jSh/htFsIFO7e15UL+25Z5GmEuDz8t4HDLSFWYcUtmex1SbQw7jmXkRpvVZZ
ozekcEXfoYZ2UxFGzjyr7P8LCXWp/CPv+cAkA2+VbAax2I3XRYGSV5w4NklV
2GzouucSbpgzSw0PVeUm7+u+Uffpkl+Rsm2zA/QHH/Clh5S8MoN311zcieLr
cGvxw0AF4hkBI5yV6XcHRf9jme3rvTi8M9bHafMJKjb+7pYrmJdfmmmVmkkx
na4OVVF8u9xtGKAifwYz9fwcjVr9Z34LPOeWATs1BdiUlL8xYB4ZEoKbbH6j
xZ8MzkHu+odT9P20YKrcQ8LH4Kd5bkyYei/hhq7xriW8CtJpvPaMmvTEx3Km
nZjMyksI8ZAl+zgbFygUdrd9jBijKavAdXI8dmfAA1xYnywsVj8uGlljs1iA
KdimmCAqjzLKBwBBmCqTeIWkxcFAqj91W3Yum+TBdObFv/6wGbHisOKaRNqm
N9h2T3wzBX4wrwq7GSRDWempa2uR/+6Xf6EYI2zQEB6p9C5mzN9GZzLAmmQ3
CU6FfTbDjx9qptCL1NlWCZxDV+bmZz4WE2BGgtVIO+f/bcGBRA+nYqrJWTkU
iOaFjbPr6ELi+JSUfw0UOQT761XB5qx4PKjI0cpD0odGqPVM6jGjc/xc8yFD
f/zwshjfd0DhpF3MYY8JiLM3KghslNe5ZCiaw1Jq1UmCQyZ631JiHEFF038L
da93G39MMoQXRKYEutM5sFCtra+JdVLbO49pMaHJEzlere4b3nj0QzER64ah
3LYvFBmvGlNgVcxpLQPgcxv0W2CxyG/WQsf3EDbrx29fW3zSFXXz+pbqcv5k
aGO+aeh+FYSoPEnEetu6ox1sSW4McQKVqh6ejxiU8QPhO1dBuMTNfBxCbFYg
Gi7NzywngF6Z08WpeWTGVGVIgXRabrha9NH694nqIKKkHN995/xfQePK4kfE
XnXTtO8Gu5LmH9ZqpCfoRbeoAAldH5yXb7DOARMdN+dsi2x7+I1SeeCjIUCM
zs7uBwKkKIJEuo8u59IasaPzGugP70GTElalRlcpj72y3VxglU15juK5WN60
uyXoSdfeVlxf/ISPfkMyOWGcADmmV3/yZDKHUhw0UikAdc1fgZ0xnrNDx9Lk
6BzMHefp6Z74y2spV3qXwXc2CDINz7jA9/NK1Zl+WWPNgkbnMynw/8JzUxYu
Z6YPdhkJvJdUrF5cfrCICWDaUg+bjU0uudtaph+VU1YZ1u3V4DJNwNzwt3jI
ML1APV504cQX76m+CywxrsNf3uzbPyJsO/+2IIsIlIlYZ4cVoNtLhVgW901q
/jcHoXX70vUxZfph6wJdnAMSRd2ohjPQOLPHUISg2VITMpe8fwek9d0ygqUx
o2vygJB2ae7bzVL7WAB186zgd+P5QEmD+SqopAGnfEysyAmd3ZS3RONbgyEE
bB4tlrhRxTeNZcd2FOmT7vLpsducIFmlWWkj8toQPnkPC79NKdgEhInJJeiA
CN73Smdu4ELkC9EI/HrpUgrHveH6ey459HtTJhK5stSpW7y3l4OQPsupVnoW
Glj94jqrUHiNjDMx5+KBJgXfC1cEKv8z2k96gUxb+6L5/D+NVYzpDoneaKVd
cpRAY2C255+xweBn3rBA4NmMlU6GxoqP6+N4I1+P3YS5K4gT+wUXll5/wVQs
yF35UhPeMcgcYBeyITedYqcfji6D7C3Xza8cx03YjTw0bq7T6oT0f3TjXZt7
GuLOotPouwgQaXZNSk3eNrZkSNarx7vw8thZpbzhNFY1M5hC5w7cRyFFBrmI
2C/Cqp3HXe4yzU5GgzYqGpWFgynGtzQZ2CXX6sM4x0WrRL8lRPm5uhSI6XJF
aDrynpatmNsC6W6E8H3OVoTT52uROXH+HCFUE9UQCifM1BYEjCFV6549fjoe
Zy0sjDoa/ZpNEPtfEQoyd0Dn1xfdPAdY9e5lTxN+qiTuRv3vFXSaR6HYuwrE
8M5Y8yE1hm6WVt3S31a3fOKDBc2C9CPNjKhjHz+C29ItpRma+CzvCGbhWNhH
0GFSsOfIbH1N+coCxkdWFuQJrKBuWIufJYB2rMaGLXiJQpUjjR7zuGzlMLnO
lzixUMj3xzsYzWZCDuQNcR0b4yrTQkAnUDfHfICpoQ70tinFNZOLPMBygupS
T9qH51IDHzM8u5iTcnipFIX8E13BmRds/6Exf5gJInJqGybk4HER/bU3X6I/
cGR70D4xNT9adu9XuWJwLlOE+o0QSw+mpNv5APLX34MXy20g4OBvMAJwzdu1
9U5MyZqaDW1Q4EqRziTIWYz8Bk+viWpaXzZgd2BrVg6uWozkQRLV0M5xmt9E
tGMbtLa7nrYiwnYL3a8Xl/qNM8L+csnGsffJpmixXgVrG7OG+dETUyKTWM2h
AdpxRu1CT0XwVCJ9bDAbTDwybGe6juJw1hBzJ0M//MeCK+sbGl3bW01MMHEP
JSUQQ40JWd7aYHBJPYlY3UUdiHAXjk3hkvZlYUFgVjW8E7iUJ712yed+nG9d
ZELbjsYOZs6RdViv6mWhafgjqvAApHaQ/VRdh/TufRBwSAKD6TIgkGntWbSz
NEbWHxCOQ8Za+0iUtKlNbIMRmx8yg0Xkip2G31gKKpNVYFV02TOPlv8QtixQ
4rjfZSLolpEkJu+Pyvdzmr68oc+CUursehWG8+XmDdxkm/VpRDuYH3obhFWL
CEuNk4JrQO/u+1L+9bNCm+CH0uuj9oKmBfmHCVlSylaEvO2DiPOOQjvOsdkm
6K5IWEASZ8Q8/kjoYZ9mxm2SO1E7hHfAuWRfLHC/8TGTfS7pt6JDj3gl/f0d
gslz8bj2Db2Cz2lpyRuT9Y0VajD8c3dbMcGdBtZg+IFH1/ia21L18csRrtJD
phez/zNG+a7v01K8gdnXQuljQX/wisPKFf3cd+/hpJzQW9QPHwneCpgk1KtP
IiBimGtAdvoqEuB0pHvKIfBK/AWmDvE3XJMcMdelDgcCnAfGDMKUUc5y8I05
XkyaHTHHtmnHCE9As/8vYiIecU+zqH+UO/ZuxXNyjitsgrnbB4Jo7eJBWCUI
MK0nuyi9Qfkr2pdhEaEtQUg6Pd3+oVxJTw98kcrOKAtRPUO0n8tx1TK7vwbg
HmG2rrdA/r6CWRhIURGZO1EgVebyOFwHxnIujxavhj7LB7WM/sbgp1Xz8gPe
Z/tu+WBXkwZFBd/FAlGoBPyRBBElQQvzO7VdvUenZ133i1gvOTFqhlUGXrQp
Ubej0j2gTD2lHRWrJXD4O6XdNK2XVxd7WYaQLoaXmBjXWK7V3s29YRuAfvWl
UwL1TEHhFu8+utZVJL+1wZE7kxsUbcMM/IBhKaSiupjiIRYRfBTFo107qzcC
S4y5GaEVDkHovf626LZnF44nH1+lYI+29SZyy23aMSo90cKK5klCCvmosTxZ
tm3SELdWVoBlEMs1y2bue2ZPKhLjLCpydlCEuFFUJReSBJVTYnmw/gVLSLC+
hGfFFv9DTgts3csWC++iXwB9vuIOwYg4eb+yK5H13ewDK/U6Ob0gdehu1VWn
5nbLQUcBRY/lms+hMc9IDbkftKxlQyVNjG0NlaRF02MVB9C1EEtdQfX9kVx2
xIfoqENqqpP+r8nA86o0g8CkpcEGit7Ho9vepTb9L2HAik7hILCnyrKQV9Az
AOMX8UBr0MOfuZu7g7gfuy/7OqYHT8bAUQ0QWcOpuRXNzJfH/k99Ybf35Lv1
a63ozxLcsu0DNnza3Se9rWWjJQlUiSvdCZA4D6qQWJJ2IYklM8TihvFlB2ud
t4w/pVEybel2zhozqGBwBoCXkT9rAYQVhk+XP5f5JyQuCD+WXogafmFS2Fly
3RIyr3GTFdc1ODGmDqOI4cDePJQ3Gt8wSEwHCNNyeHoQm/IGruEkKP1G1Dxn
K5nu00ya9MAMhitLbHzQs+42CVwDBlBpHt5RxzKCksFBYPPSjBkQc973VW1x
LMNpW1r0F7iyPqYHpHy7nqajnyl3N789zQwlu6AlKsBTIN2XFw8r9V5z/WhB
sgovMLc8cQcAWGICOLrUf4dfSBnJg0ecGB8KGnoAE6b+bX5yyEVBvEtH8SLv
Xaym0tu7xzXf4g7e7vQyL2xrlFqkjIBZu6MrgFm2pTVoMK2hbP94/LNrKfGf
cZ2B+N0Ij7N0OVm5mikDdAhnHBXvBazw0iNP+j2ZJqNzLiDfzirlV8t6NG7g
cYp4DodBMLlMyz6sORaOXEEqJ2VG4HhrAugoPtrforCMnblGmHRrl7Y8b1ih
GVKHFo/49ME5T/Krc+VO7dBNqb+deyqv1hjLhxRnoetvtH+27oJvM4OMvp+O
6SVtns+NTSelu5XWuKfmhMtKoMw7AHUGUqb+4RtLFq/Uk2+P0wpiMB0pmj1b
fg0RTsrsL2qITG5DjMMTb6oypLYVJwOJkKZfoLlHd+NHX3NCgtx3ri5Q85mO
kMOzJNwTiXIooGJe9fGe/KaeWuQ0T+pkMQpBNjpok5kxGL2XcLBTYaIIqnFA
i7AJcWdpdm8NpY1riBUoXXaD4wE2/UBRQH00vFUm6ciLCE5+HtI8LZ5gZs55
eIFNAZi2cvz8+DH5tQcgz8twK5gGtBxb/Eeb2uAzclH6L35kdUgFILFjKkij
GJJC7eJTt3obswU8X+lYX5L6Ct4hrjeXvFN2Fvsk4o9JH15JORpXGtamJHFu
H4cUnfCRPhDTSF9qAv1Ka/gC8oPMnOP804WV382hyWSlxwsxOsg/Z7wp+/JG
1H4RjBb5U/U4qVp6fo3X4hF7/iWFTs+UGgB3r5+ZV3dNzo6hDtQrDbOHRW3+
yfHEjLUNfqqOCIuR0XpkpBwylk+eR557vXsM4DGaQbqK+V0qMujT09HQ3tMP
SWZz8PDYFmaN4mEdSOmqAADBChMNK4jv/l2YL7k2TbK+TSAPYwgVZ/BlX5fm
/D9Gdlq1p0fhYqAIFGB7xdh572N3+eZHJ0nEbChSGE8NVXVRtEjoPc52s2KO
f7jaTvxbzjGTuqoZy8gb40EwcydTJN37QDLZx30ldqp9Ol38ZLT0vTd/Vlzt
wKfq7W0J3b7e0vNBs1juAieZmRgwaOn8C7qyoGDQlBtuTK5qa4WdaFzEr8jP
gIx1PadPocuTVb/9503k42hiOaOLVrUpI6BnXnqNHnlcXNGt5XP7f00BCrSo
bYv//Lek8Ja5EfoGv5l1go6/hENe2kXkJ4ilh5syAnDZJPmxHuYS0gTHyTWK
T5WGEJuUslR96MX9ArZ453tVQgPkGvLjLxSuvf97j3P0tnJE3CJ+RbY3UtVl
5GJKtQZqjneSVczED3ykMBr0hfSvqn6yB9Y3ulR0xmBIZVTmDMxVCCrqfcJH
eRjisgckprqWS7LbrTacDLS46j1i3bftqq0rdUT28kHvFmkOTvArUXP1fcOw
BK7qsbxsNDwwUFu7oxyhFfNj8ARH4cuXsFenMqxCwQ2fd73TsU3gCX7jNCUm
1YSLQuM7euXGXgSrGfZF79VWHCnvz9GUrX6qSV+TC6V0dLC7NTi7hoboNWeU
9E5Tm0Y3+V21JE7eNh9jOA2TDmiy/bRRc/3iTD5GZjERFdcCmUk+GHfw1aZb
7Rl8CnY4hrzE+KSFMDdcgrEVcxwaHWviQh9CcBmZb5tupgtEWyPv6Na1xVli
IDZGyk/oBERy2lzybJbZwlv67SsnD7IOblUlG2AscShXlLvuA73L5Dp8accg
nhmSVxTxc+pHN4TBm0qDtISmXUL9uISZw4R2Ie4l8hTFDMDCN7E19C3Iljfh
oezk0imkhUMqXE1aC7u9S98RC58iPTxH+Js+f1zEqpRR0MgV+QDe7w5lqg2/
saYXLK6ixAdAMnLNX4tKJ2vH6JKSO9mU1z8TLjZ5b4od6I5ZTedI8E5s6uJ6
g0FCebW8egCsPboBTXW5p9Qx7/sxBnELzamI080jHxkBTv1oFIhHSHZc2UZi
rl3Chojx4ThMrbIpTLWZ7fmjBXGY0BshgLOnuTAU9S+n9oREbZW3JcO+Bd40
JPS9Z1EUkIUZKV5jdqnJm1Dv6YAreBr/aaD0B/KSw/jIEMehmLZU/e10ffW1
LemptEABhgxaK69jXv98SMuhTTtNA6vY95bSVcLoJfw0fTLXK467thB0TyMv
TxhnQ2pkjfIEP+bGhSU1t8QJB0UBU0BcAf6C8vrcSvRhej1GM95sJ0Bt88QV
QC+8VGmEsXWWU7E97xJM4SBdy4E1AYRVJKzlJ4yu9Ew2pj84i0Zj4FFrbafx
og/zIBRnSu2Qo+dbB61bHlFBDzqpzwK4vkQuRMkhAOxuKynyRAvT+ZnH9Yhr
WPMrgpCcpVzWl4QE0t3Dssvag61N7HkusfD30CMQA6SHC7Z6FuBA3VifdSSf
rRfIBf5bYMOWev1RhQlfiTPAmtwOEnmXKXusy1xuAnJ996SlNPjR2GUp5bLO
kXrOUDcFEzfyRxaWMwKUEEwp3D3RXFHLekPDeURRb3nHsBv6UtceTthMto45
caXnZsEIGNJ87p86hCWejv3FYpuYVZ7T3V60AVymgzBYUR5WQ01ztRVSNssu
xcFWz4OwUSn93MxYgl4i7NpSINGjxs7nOCVF66MPd1zfRHGqGAACHszTi6H6
ccs+/hbAis+9gKgCUhv/58LZOnW0dw4EH8Ctpp4wfgPJqC6GQ5mazX2eMwye
CmPfCOJq68URKKo2gPnZwkqgHImQpkzXgTOrcyuFRrfW5HPHCPydCpXT0Tva
nqestIft4hG+9lnreDma1Uq2nnJ43E1N5rIgzog8sAuyqUp7EsIPEM0wQkvQ
Pyzz507IymrfMdNnwc7hoafrHWRVWAOvNWV3CP5Y8LknLvVIjNYNI26dtoQw
WBKyU8/L6nCpJ0TOrBMzOk+t/Lyz/3bnkLc2o6fPYpTthOiLwadkGBjzfdcR
9Z10YrfiPOZ0OmtzffriKZXw1UJ0cUlw35vXaY7v2Dh0FbnFlA4PVBXeHVIt
eGIzEJnCdvppj5uak6Qk/t5vjFUOLKgjBIHqmhV/hQzcphqmKJWsdk3SHpxj
x4u9+HdZzR3RWWw+vujKP9Q87xHj5nVgDAArN4RNNHDE2cntDEBp8vo5RQG/
LGJABcNp810jBLN4yFTBBUX9qT9CJLw0bSPVem4liokDbZ7qy+Q51Y5/veTB
6MCNsWUfiQxfYzZLIHjX56uzAp6y5p8sUP/FwJzuCI+XcIsOzhrCY0Mv26J7
MiK3oeJR5uBWa/FoFfd/MsYPnNSh7G+tZ+WPo9NCqtsJn3Q4RoIjfrA4kN/z
SDei5uI43m+jHD/Sg9tlvmdE6b5D18NoWSXFIDgSTgsp0RvEo8zBpozm4+BI
LUyOp2tTL2u/N8Ohn5YsgdJH/YphjbsggvZOVsOTeJc2nBGHQhyzMoW5szGQ
W3L1vuOT/ahmLQzVVdgxUn9IzJ2QkqyXcqDzt/mJoTte3s+GaC2JqaFbEzcH
zc1kYQ4vaOtp6eViwHbWvCrUqcdjuTWYWp8wpb5axVDga6NrqYtsmYZESx8s
daNEAgmWlMk7IjI/ls59UclFvkKG4yrIeYihGEEfllq+So6SkJh2/q5wBQbB
FYUn9jFc/b+VNfoHOeKv02zDxfQAFu2HTyLLGWR90Huj01gaDq+hJ49HMEtL
Nf2Ia40+MUbTxGWHgHAdNlTWTBQd8oYsh6Co1t3+bi2d7TNrFqsP56FWrKoD
gcx4kI/5FUhE8QRb8cCtuEs1ozp7DXsdbyqe1spxVf2G/y82m+cMk06M2tUZ
YH3zc0uY866Yp8XXMh4wnUXoi9AApwib2G2SueIS9tJ3upRlsqhMRlEbBoqo
i56L/DBVVJzYeGNNbOEYqHDGWDHNTtO7F/WgoDu4wLWpuKRSjYA4Hw88gp0K
uxPG3qjCOLa/60t6SJUuxP2SL+30v15ShJ5pruE6h1t6JAdtR+hTL4WEy8mx
U17gKa6XwDrfi6xIQU2ntH3G71hYP40S2R2kKnKfqlumuxa7gpmTvz39dObs
OcYaDHM5gIAqHyf1z3ShmQ0xd/R7FfpOGmPp7ixodO1n6l+6ny0IjwFHRyRw
HJp+mznuI2W9MdI1AFrC1FI6qnk4D17AkI0rY/oHtotTyd8EUElw43oyAsW3
phafMRc0um1sed3SqDsNYpeq3dDXyBlFRyUHmzY7ayVrs21ziixl4VKS1Nib
GuVUfg8aSiPgsrJzB0Zna2R4HimUTBxym8SH9mgPXqebzMCvWke2AJnvphFK
m7appcSZsb8B+KuodBFRYngkrZ3OCVgBuFmjbW+pQeC0tr6Ck376N79/L4fU
OxQTVtoxNe+fRgC2ag0mcGXPu7+IrdI4PIfSt4pGN1L/6u6UAxJux4eZXnbu
OMXtkFElXaJD2pv9+kR6TDrDVVEy2S/QRtk0S0lvnjRzRyMmuRkR7RZbAskK
2n0D0qyxdFxuO3V3BK505e4CqYMcCNZMk0dX3TGl1SLgejUu1iP2Bqgua9+F
6e4HKRWpUvTgmnKL77AnbMU/L0Ne+1AhcZXvWDVq+hURvimCjzc2aA+AkJC3
L0VhIUYE9U9mJKgXvCZ+kbP+RNrWs19puoPEADOhFuI7K6sQJTfC4ELeiVka
dL53qedkz9MXzmocrd7tkbLOPN4iHdbpUJ4LkEW7VBLGrTMR9Cb4jupfnOx/
57Z9Xsp+9SDz3IEAnQMFSotdRTGKSZ7hZEG4tI/bsW10rarIPVeZLTcuORPL
NnxDC7KoX/IP2QagYhYe+hFzJdkZ2ciJ4qYPx1bPJOT+hJ76gVmf/tGGCGTA
wftKd/0Q6Sb/0rCAKyn5BTkNOWnT5LFDpCqdxXqcbL/wpL4lbOB5lNiFLstS
/ZKfispsHu/onuiRxQOrdwY1Agq+i2CeBXtZgxsxc528vuK5b9taSaGDUIXj
doLekKg/4Dm8R5l94jxN+c1W0o5grzKuQw0KXY6KfOdneUCD3E8eq3TewU6I
yYHNJ2R7qKUaiVsnhVtGjHEWzCzMXZGbtr2rJTl1tHyHaz9IKj6xtMKoSYzs
FOAH0RkjEsAcxxW1KLtK20fz8fXPszbJaXh+5RMQbAY1sRlZHZi3waoZkKfA
la68g2DiOr5Yt7Xgv6Nhe2riB90etEWNihXHBGLbMMChXbCEDI3HDBry4jOM
LQh3JjgmimTkXSzXsNl4zXB5DiFTOMTECNsTTs/uV5/DbhNL+b3KdvtxjWbu
e5AS5eOU2uNQy4xaex4hJPk/3gxtHsrnm8w+0LeNoMYDB2D2HsnTQxVbz/6R
hPPaXzXXLsVvglasgZ6bQToq2FZeZIwq6s++JBCv5RKzyPNiJW+vA3D0/4JA
yAmb7FSOGwmO/LrGpuGyxrPzu+HnmlGugdMDAiJ4nGqnlYOqU+0chuzDVtMJ
YEcSQGsWRuq8ljj7ajSptZvbX2H9GONPG87bXY6JaO4TfPBBkWyLcGQqjCQz
sSaRaNQyzimXHQ9duPXPgvCg+VAR6mb+McNMuzzpbt/ThSPYEhhvz9n9iOdH
ElHIO39UDOpRr6H3hz1tlVWKAuTyFoHkfAwrIQUTnBTXmhpmpOsnAwzbzzk8
Q/0SlZ9O1pBX8c8loftidqTPFhgPJtsgXNf2BKL0jJePiNB8zW+bKDe7s6ak
mCDxFgpqE0JChWrdVpPl8sc7ZYW1ogQ/pd05S7/ZV0FRuX4x6rQbcVEjWOCp
cFSgsKke6jBGWrY1iF15/iv2esxy6mZJLWW8utEVqYgPF6s8oUVO1hFA2rTP
TAisjI+c5t+tGAcMMl4FPicDJblwztVjKGerSQuuk3iVYqLKWDCQh8ujfNPH
FeAZ2B6wNdwwiR/FAnWJVruXKcRV4TM32gnWPmaGTzTcZOwoQt66x+GdTDqF
rRdcDsI1SzouPB+uADOiaTXa1RwSI6McqYQ+VMtyrYhVzXbH8Ybpbyv+wxi7
k1gbwvLu/MwiIMfAHhF8OSehAYODeAappxzDLQnP2WFfvenJ5jwVnFpj3S/D
4Gznzposzj/L5Xutlxaq9t7Hq9uiHUafxD3kna9022BX9tEAUeIL21lidfX0
enZLRBQTUPSHJxrfvCzHUb2LxB1ObMz21iGxdzsGblX92b2EkXjWUyTkN5+j
/65ZX0d/5WBcZ2pKoamBSnreiTq0fd2Lx8IK1O8V34BUhyC37kkREvOGDH1V
Cn437KK+lwfkq8rA7R/pBvYVqnjpHDNaS81aa5b2XZwcfAfGNj8a8cDt8hMA
/FtjMQZ5OgGG6U+5xgvfkhCFGPWDC8y55Q52vCsP2GGG+1vvbi3N+HwOBNW8
19/H0CA3iVW41y9t0OIB3187dr9ZTSmbBdB6YMfswzYs0xJWrg466Rjn+I80
gLlB4an/OcBm2HsJtetVXy0MEfSJsm+0QU4lPOLlZ/GBOSVWuocXXF4qKxzM
/YZGWXYkRZoE/H0RvZSlvo5BMl3uVh+y7YdddLjEjVv6uY5BlwU3782hHuht
E+5DhM1GQziE6gXL04Ob9EPHfV0rS3Mh/qs51ZQHkCYnDGzIwytGICnXXv5P
8lP3tIADHjxmPNLXPbNLFec2jqKXdIPlLuXHTvxQ9QmqCDAmf/+qJXMniCQL
AMmZk8KsAVLhU7bwzl3cDE+Z7Ofc7Tg9zNScBk+JfdD6PxGQdWrBc8HtmWrk
s6wDsnYkkWtDVa9Lc/HDd0Jbs4yAZ4YPeYW+EMv1wpcktMRV4on0txTkQsVK
2FxUm7JbvgeEgQXMQx0xlo76ok5qNE+MJ7Wd9v1/4cZncf8kwCoE3IW40bW1
9Z+AqaoXnHVTO/dp8lugBSiWYypcyMpsV9bvKL+6ofRxjhw7z0Hsw3FHS1wE
Nz2waUS7yXk1npzWmh+MJwTGx5nz6gZ5k3uKeUnvEq8IFTm3VvmCLDPN1FK4
GM3nRwGQ97pNDMxvCmeRqCO2VAIflUZKHWyrxDqTJowDrlNyeuSf5ky0KT5Z
5fsgFu/G6b93zauP8lmYHL6X83v9VQjxLl4dcZEs2h5ADyqavHPOfAjvwpd2
vloAy/Y+Pny/3B1UcP1bl1PcCBqhC5//YaOtuBOwkLMEeHTpXhp62ejIZyyG
VkXlZ3wHWlE/nSEx9elMxMk4cOLPGEMQo37U6dvOUuCxb0XgDtDAf1oCwTMc
+051XSKvwfu0qhASUdiHIiy5eZwehmZXW/PcYCha0SxbcjgmofvXcLSB+lwq
FJdg5+sH3whJ4a4Mlz3gHl6cWHNpHeF6VNbgR2CFG5AqO4Knd6/tcwFTU5f8
OFmb74YycgUnlhU6MW25VvQUVAQ3TH9/krSzcpUtO8fxSkMTirEwywCSNYz2
Oj+GimuCEjySSQCk80kTaQBHT18GmV9Z2Y3381LzeywYxw3RbP3GF08WbRdD
WZNgww30pgSzImgBAigXN53oITtizTSmKVNdLW3gS+wUKzBaVfmmB/xDiTus
WWsYeTn6oTVrt448sowv8kd/7qYuYkNiCjxh1Rz3nktC9CggnwZUOlOntKQM
zGcwl2svnto2zkjtH7WKcmfnyaU+g87C9u5HYg38TJdSu7wyYzhefZLt7OdF
3H7iuBEp8iU9xKSJBpBqgStrAvklvunmvRIxfhUFgEtFuoO7xXUHQE0fVyG/
MN7BFaZEtqwKcL7OMCqG+SEDcLU1iUGixgWXvys72xzk09R8vStk8tvK3xLH
HPLpvulETpNirDv6FLdUWqIefYciBRSxK4kNRQXQJKW24jVsMN0zbq5HDdKr
bLonEOogCKVk8zMdnt3zCMvBxkXRxeFkxWNGTK+lpgCMUkmAS8QK2zbdTRx1
Jlwb7N/wH2S4NbQR/W4DvbVgm39nsEcaAkK2VNnFDsoZD8rGkVgG7/uEAo78
WGUwHLzlktyzxoKfF0cwuYo8w0Bn8YrywHJ+Q520P/bICUddF8cQo/4/Cpp+
BeJfy0Jhomp+VCJv3bEcAh7PriEZoBkkkyUu31XgvmOAXuC62fH/MrtCzT+R
poYLXKbN/KoTNfWO0Nn4HU854E6P+w3pSSB21NJXspetXizwXqG8waVWJxi0
iZYdIxh2Fg03RtKeaOCZOIbarUDNTqClsIKpTH1Xpzdz7RBLACtWixrgf5vO
iMA7pLao0AtI7uW6+voZJeU8DUvd47xFauK7x8I1k4+OrfVDfPHJdp0jMqUU
Jxj3YROhZZB9WHQFN5ZhRfZ0G1fAo/WiXWY25gbhvWQF6mc4Oj1j2iBP1MWx
xd+WvjsOfdz7Uyi+wGWMH4iI474XZ6HNXc4GWgKpHREbLSNa+9XiOG4JvIok
gsHEfS8/joozHlYK7gFh/nAP51CRCwhYoSDQFXNAuB5zq2a09EoSLadKSTtQ
nexS+qVLmf9XKWMts4h1LvUdziiqxKiFq+Nco4zeRw8bB2NTmvYSVCW8l+FK
39CMkxH/GMfStnxK/d7v1X9ZmYmXVDUf6aUCJsDKAokSWqZrdHTbq6s/JzEW
EKUPlU5c2YasxUrQxsRv/W/j6bWJnHdj7GDIP4ROOgWu5PKTzP7My+eDcI1Y
ZgJtaToVADifpUF71CwCzMuC1YwoCzD7jnO0XTZPg0TUSfCYzC7xe5Jk9Lc/
nh47cCzTU7RriAMaUMDvFQmSV2rEmthcnQVHrOYDNKeJiN+qpHHckjBjCvtF
IHHKVexjC0oMjVkGc1wZslUQFg/VoaFP3iedaJ5J0ww7c6Bsj+ZTzwyjDAhp
p/N17lGXDulW7yCQrSskTrkjOMYMU8czgFpfaNdimLpYqp76AmcFt2X401A5
Fm8cDfiGtg194/Mw/K9e6tPcqbTw9Kk0XiQ06vizeOD2/cHVFLiXz22Y6OJG
mjQRvzdMjBHi57JCUyOBL0JIAniZ8CLjOpszskDzZyqTKh82YRM7OlQ2wg87
bK8WARWmzJ3XXPHH9jLkbgKeDeA2rYVcDxKMSWznown6mWYk4Glf6gWSYIXu
rsqZ1VdlyFB6/M5r5KYyrFhYHIh3SZXGoFmPMrewGCWog5F/aHCpuC0a/30l
d19CRomrLn8v8Bw/Fgh4lQbdKGpNNrPVysBF7C2CYcjkY7fL8ZiSQZVbZDE9
wJUtr9kwUclsSj9mOJRA+raaGwKP1FbRRefdnzzMOUNip7j+ympCoCKaIu3H
lR74ocyWp4Fi06KsT4qsDkQZB8a8UnbjoZCeQHKki5jZyfWht88nIxUNt6Yd
PK0CdxxgUOgVkJXHi6/WOAa6bT4et6LOgihSLVi9FJ7jb+eTUXLmRCq2TVl0
YPjH8gHGLvijx3/wOhpd7qUdt34HwhpUPuvpO8gCTU9m+LKQGdZ9i+OArhRc
gwBYj3sAhf9DdDZPKkTvycBc2MZR9423GYCwDPlMED1DMlRr3FrIpAIjWgTB
qZVFXJjeQiTiRsIAgfmymXzNgBWQ1N8eJa1axJHwY7RQtJfPrGd8tyASrxyp
UIES4EATV1X/GpuLz5BCaqQnIdi9PFh+h3qhcQxXzimj0gSSR3GzWU5khQGO
fvPc8ODvYd3fRiNYk/mBg72BZ0C+qQWTA5WX2Hh/JeBInBbaXwmGyROWzljS
2I2y7OihrotiFvNPJJV7mPBsEQIKgpF6PWhWeuD99WCf1Wg2dwgmtqF6JgFO
MAKfRxw2VLf8/YptVc+YSBT3ZBIwl7k8/90h7SBrIegXSPQ5M3qGJULIh/wC
vKzFllhui0Dr4AjMo+vQYZfWJXOKVFaQ2rdahmt1Lo3ry2ZGgHnfuorGAB2R
5mlN/a99FfhoAiSpDn2d0BIHs7QyGaEhEXxcojZw9keWsX+iD7bpzNjIh/NW
45AQaCYTLLA91xJf9MUv5hVno3TAdmgq5LlQhadl2i7UwikVVgXkUzBrPxe5
yREMoPBFg2kiX14Azaqjcdt1GBvuu3y1vXL2ts3Nr095JTOtURxfgASZgL9m
zwzPTM1VY3w2E9BmwZyUsYd5cdDXulYWdiwvYWnDiryFmGcSRSjMr3DO5GuG
Bf67Qb7XOq8ZSC42qsXZmxTM7i9JTs3dgq1r4ZdY+0YXjCjh00aUexrOnBBX
PS8RV9xsUBs6mapKH29ZcELBaS5D2EcqB/i/t1fV60GYwgWodzRx84r+XdIZ
oBaw7YtrNe++vGa63lJEpiJ/sgeNNwoBDn1rKfOSa4iRfk6SkyN8f0LV+Svx
qqeKBFOmGtMNzSYE9cejdx9XjH+UlUWM5CIw0moNDwnAst247Ke12pi66Odm
ZjBcsVsqNIkgU6OhN9+GzXKUUDfdMGNRXMGRECAdCecOC73Tv+nCPwwsXFjl
kNUqImePYfNoq6VPIrpd6cIlhw7L4LgSc3MHLYGu92l1acQ89CMEM/3MIN6V
Aze6z7VUN2+Lxv/OZWYR3VSxwTrUdx/8CGjjYcYVvQpTWwPUrN5fE4kt5Old
AflCvN3hj8pNsJ1OxY9Fjo2fRIrCLrW+0HdzvwPlCbJeMKcLtHilEr+PEEwz
c35IkekVBslt72OfTNkuQxemRsUXovSRj1m0p4U9/J30ryH8wy+Re0h8rs3k
/KRlu/BKIlY7tNyW8fpxR+IuNMiVOzpMYIXBM2b6roAF7NSq6+aYrkUB/+60
leiQ17gEWdqzKMJ8asrkTS5URjM97728PfXHx1ptLxkxzK9mf68vEjHTCXx/
puqtUie9jyalwi10PsEiCm3dwxgVit6se2mJxFVQmuciFPkm2P3tWioZhpY3
fE43gXG6f9Ue1qT8VCPS1EiPG2yfs3mr/p2ExG+ArpRzLxRvFh9+TrGI/x8V
/VpK12rRdFULzJ9e01Gt9NK7U8M5ZcN6loD6u1yRubIl3vxMkHGgLEgYA3cK
68KnrL/A7S1CrQZbqP7qRQCM0UxOo/EOL15aorhMlbGTZb5W1arOc9Z5WpsC
bQR5//MYhck2TES5BF6vxLHCcavSbcr4iSDQapp69kvo8pM0FcvQqNo5+2X0
oSc/42bUAYTIhmX377wDI947RxV45J/DQOlgqA+QwJHAqzqv3EC8HP3Wzz4w
owxnbOHLxQATPumt3B/9JBK4Nz50+AGnFd5CVRqTBteX9qN+CB9SRtfhfo0X
TbeYPTYSnxcVdtVV121/DCL8h40kAO3vFppjXl87tvQlwzhpzhly+V3EWDI3
YASXtZYzajdy65MR7zcNE2bh08Wd+ipDxi8D0XTcwj93QVBzPoejS+0mELBs
GnWTIkpjN6E/cGZs0AsmpeEx25BYqeEKGk9hMdZpn2Sqf8aowuhifCo9DA1g
N9v32FzajPRWGecsadwHzKudn3h8XxhccS7ivdJw3Jtd10t8zuZyDLd1mCNz
GInP/sOpC1u+ahq5rGjT/NDr+SjoIW6sAI8sQYwXjhuYhnuGPT+06TeIvski
dva8paqvb/f3anlTKBhZ+KKUESbF2lldQb/wPIUdjPnSjDPkS0LvlGIieQ7V
WL5jMGdZeHuNpDL4fZ/i4ubbWMEaJg84ookAF0QNOPTktaqs2eQnCyyP5C1j
ht/YNecBs1Xj3Nys1vK3F1oU8+iB2UG0Ou02OjyvwiC3d0hpY15PlVGTZY4F
6C7VcyWYGfTNRTyV2wDwPTezzw3+IOJKXMPSUFVeV/S5TpZ3yXu1Js1GIbSz
lWib8Mwo9pSXsIorfzYBen4lRbC9Qno56h4JMWCOZm1MfZRJAHWKkGBgZUo9
EXz5PiTtRLjFlNOm3/xyR0avcSgVhvRAqQRdkwbnS+4GU8/ht+nrhNpR07m4
XIhWpWdLCmTl1H46OEQ70LzDbZ5+ITRJQ2RIQUitbyXP+gERS61caJPqsT71
J6POsXi+rZN1j0VACGd32rJMpIS6T8L9jd6Bc30MP8gV1YRBSZHu/yUgmVyp
6YjRjGJDXzOFkpcFU9SV71USUJbyKOuml7faYmnd98REyI7N9spt4dNg3xF8
Zi3ZuX0pLjP747crHYKKU7GRkUlVJy2+y0Uzzu6cwwJjkrXXOIyYnqFO75Mq
KhEgDjqKODTdsps/04ajvo91NrzwCiUg0b5yFNu/pGdIO6zt4TNGrJfjtzRw
MXo8wf0yk3l266PpoHB/Er7sv11hxGBlDbf0V1jmbTAwHZ28B+v0McgkN3bY
QpBgcdYtO8VisxZzrSCp8zCd3bcGntsjHZPJLy17cl0VhlkuBevF3pxVrMtM
7sjYJJZXNkVt0i06h/NCaRB/sucTRhyGZPU89D2ndSiqr2cZc9arCnw52i3x
NgQfVTLhQLcUQ4PmA9QxAC1GeiRE3AmZtl7sIAUy60iQWjcC4QrFVB3ROvIa
etgZSC+oU4C/ghm73N9efAXE2O+ffVxXIZ4YWqRtUdSKPEfr9a1AmLokowsC
BY47VeewB9vNQUYoQzcIOtETplzyCV6g/6eEoXUwVChp5mkZ9T1ZMeCFNSgL
1r1QuzTMHEB+lcvvY+CqMbCcvKbczq4f+6Gyx7B+p8ff6KNEilDGTtgPdQKg
8GeEHpH0yAu0hm7C9JGzgkFHKXPZXz9kGRxGpruIwoOvqWZ9cvESgPbIyXpJ
mEzlDz2YZUttIU6fKOUYsoCCB96qGcY3DaepqRLoL2fC7OF0Z5Vmtm0EByPB
AD4yTaA7O56KJn9OCO5xTSBU7cIVm9qJpjZ71fsWe+nHPTf8QD81gYLhF8FQ
pBUWhVLg3XrMoinZxoIdBVIMoCwv7BNn9s0BbISySbG9DXeDWdyMwqTqT/Jz
LQI7aXxMIUnQzJFKOBALF63urvlves2i+w4nKDK1L8fiwDq44YtyTyiQtqEc
uqWgkObC1dalCYbIxehWxmzVBc1T2/zqbBVTPPFD74MVuMeR7hAsj6TYNWBd
yQnfFAr+ajAdecvHzVTGzJwAx5BbGBOApAaYhrZtjEs8LV2bzn7aGSeiVm0c
5oa5AfHgppKqBx3BNEr7X89zFkyI3COKplpDxD/JJSNwxIL1Ego/OGajSr+4
dsS67rIsNiKnBkVRL1BZh8Q8Pe/WNQQAVRKaPgq/l3bkldFS3eEfDzxyCaPo
D2wK24f/XBe4dL4HiA1gMu6ONqnDXlO9WhH6yNOVUCZEvkSxl01Cx/kQqMgH
F1Y8Kfbb6dSz/rtaSuE2LJrtnp8CHCvso6O9rCygKkU+xydYbN4rBjO1+QR4
WidTzPbHPriY/j7/U+EyLkIR53WZSHju09xSSboTe7Qkve55MWtVpNYmTje9
UWtSFpOkuM8ETXrIQAY64hMBY0P7gg+9IFwJZB538P2LYI9VE9G+S/J52PU5
zOlU0bykY9WQ8AgGUrAPKlGm4BZMScRgbzxUYBqVKcyf4Q68DXgSN5E/EQ6f
VSNyI+fhhDf2wI1/WFE20lOoEdjJOJXbtZ8/NaXvgbPI2ExHNsLBEIZgDKuu
EKP+16d93uF3i6EdbUbfsTiMDmLLIHH4r9Ur90VofCUj2xJbC6C7jpsTrA6A
SFORxb16e4f8dddkxWC3WNMtbxYm3TOg4BfFCpzW/v7s/mWMLbJSL/ugZVy7
X9ed3yVKp58Sv2uicjFd1K0lY48pXqaxFlh3GEJWlsB+z8LNw+qlaJiG195g
+OCR9olzItHI053X4rnf9VUvg+T1AOlexwdzuSRuukJzeNCijxIKwwURxEYa
kZpb8EpsRZz3PYIeFkMmkz3HRXf2640f5X1LeOzzqMXN0nDUoi35l1wc0ezR
jOJ3NB6W77K9lvTNOa4sOscHLaeTMepF4Lrnxrz8QiCy4U1M/+RV4QS9xtty
ZkMtA1bISH9irStan6+OfEwFW2EosmukkPEBVYYZf29z0L6+guu8mYOTygDq
oG+Nfh14zjEEIrjPZIOdKqi0I9fBLkuZbXNTcoOvSInU6gBsCoAcU7Pv5SOA
C5BzlPvEE7to6oC8fHiVJI4mvYdPCugefOCuDYPOJuawdSzYs3dZjQ0nVcoL
oi5DBHR+Y/kUkWPF47sJTSELIfdxbie/Cf3a1OaczfKn2AyA780QNnRy4igc
Ul3sK+KHtUelqR5zGywa6rPYBi+OQ4EI3oWZ5caOJ4iZoygVuMpmB+XBNWhL
7tmM+VT67CvDcb7T6iX9K+BO34QkgLU9bldhsbYAMW/4ITgp2kfgpL8kYloY
uTkf5u4jPRqWsgVLlp7wwX1rLIAGoI/tQFEvQNf97aBPc/kSR165vnQkfPE/
Pi1KvlWVT87jQqt/Np3GhFTWZwpGpL+66HfaUjSWCtYDu8wPBDwvy8Q8FUJ7
ZdhrZD6Pjkw/fbzq/4hzeAxPp6yF8furWz81r7VEpkYNqh1BOgPw5x+FlNkD
iGle7gGQV/3VyzxOUlaTOwm/kDihRzorYmgsf1IiW23B/o+ACeT3Ih9IIgRM
wVfgmUqmTvzOWr1AsIrFWH4usO/ur9kBRMhXRpc+SkLHAFyT/sReG9vgDhoH
Qo2UEhH4d5LUHPeX94AvYMP8sRbSFKoEmWh3CDwZ22bZg158vejm+JyxKl0q
j1Af6c0b+WCwoisvhKHNyRQEBRHSXDgy/PIb5DiIObFgz7U0TpCecqi2N04H
d1udhc2hD++nQhlUiikh/20QNoJkgTeOJiJBCZK1VcHxuldHk2iO8NTG9SL4
HQp8z50E5YrhT03bvijBLTT1renAxixsPOwIuL6V2hCH/NH9VFJBwl520A+Z
Mh9CJnTrdZ6rCBq5FXI01th8gBYEzrDMxLR4R+ZrROUTJz6ZeEBJulOvwVVe
aXIQoldwmGQcHq0mbzKTtbFfgaihfL24tr+NO+SR07UHdOYf6aeENTfXQNOU
jc12GvVgPChYv6MoHTlH9YhBKdJBnUEXq/5nAtuvYSjfME5NL+l6Gr9hH84L
18hNss8RK/YjcMxHks31sNYmvHqFGmFl9Pzt74CCvz3MWwLTbtSAD/OmNDOM
paWlaY8Bl0igQZuQjyBZVTbQ3ZoLlIidZyyDcCa8EIIDACKeFpe6EeUXPK/E
XJPAr93RYuMNgoxp4qEe/H7/l13TNkF/H4Nzhmv5lJMyZgbt03bc2LONBeEf
PLm4URdZYI/wIoLKy2CWJ8hLrAQ25B4IZtmWvAEPTSYqiKEzSK1hz7sFj1qa
ypBBrzkNwZdWsWpMjz7YDfG3WfcVeqJLCF8Wt4TEcHth/bPNlamA5FkkKIA0
Cd5fTW5S51bwQYJwzXNrm3fERRUr285RoaFeCmV07sOHNMCgwkCMnMOeRWC6
h1QZPJ+vrXQJidgJAyRosYQhETpXyYFBRxoVFrRZrKRKboNm9EBPVxWFtrk4
ZBasZI3HHj1l1HEzFOVPiu7fA2OuYnsbw7DjE5V/NPSPgBZIV8zcVHdmItXh
Hq3+iKTIoEzg+BpEpi2W0xkDDuIlf8Fr0eOpVmBpp6EhrrXBmypdSNu4vGPh
g6OKVR5sYShN6EUairHKZHP9/ZpOikpYSNg6hfdbV6QAcG/Tva5tZIFW3t/f
3BKT8HyyCzUA9BdQs1h44Cnzol04rQaqtC55AjaPhuK/tP6MScYakNSuUAQe
Gh+fKwlbxVMg/MDhu2BEtNLfv0kCym4W61HVqUkp2KqPiEIt37W+5hanFrTC
cElZaDO84gPTnP6XvuiYe6Axwqtou3xS24ZBrrxuyp22PCjLK0utJf/rc5Ko
iPvZw7mKpWg5Uk9sY+u3uWGiKTcpuinTEObWzIkFGO9zQcNtJ3qJtlZt8ff5
Rakh9KfO5ZhG3X2aC5C+PaJGArF7S991rG/5oJGReJfEeVl9WeqMFZ+dE+Cw
nHtG65IqHwrtGse0HBgC3z3yHReK9jpP8L3eGOqwY/bUkZ6N8E782cWH9Xnm
Qu8gBGBGTljOJAQHfXIbjvS1nBac1Om+cK5JocXPSoyvDpV6ZbSpRkLGH9dT
lNEITUigrafeJhYicG1AN6CUArhIFP+CllN3EC5niVcGu1nDnlwqzb3f586E
RpbxRVdiVgrBNVO40rM57CLAKcNv7pMeQXOB3RRONb+Z83ZW9XMK8DGFOwhH
QZH+wwQ03Iih5pc8nsPpFmSBLM+gt0a092Wbne6LcWYQVB29CCsiI+ccFjCE
hCSes/3PO/aF4c0t1ihnyNmvP22StOFgnqsMVfj//+GiAcLQjy59XYZPIA2T
rKTfUqp+yzCMdysWDbP6FVSbbUS9hEYyjl7M3niD2Lh3wvVJbklEI/GTrkm3
TTgcPWpYZ0pzKjW52aQOA2LWRAOLyb5u4EM2EqcYYC3RuKvG/rl94gFeEIQ7
5spLoJ/YXhXI8K2bF1Ygbj02y75oQ9oX8ReoA+PWAVJSnUcft4WColkOsKXG
2b/JK0LWpMz1g93cbjvAPGCs/qb9czRTs8lDSZ5wFi2EPo7zjZ97J9mzPV89
dNye+n2TaLH6Uv7+JBpqIwcEMJjI3l1Oqg+sPLTLH0Zc5VWQUHxgoiWERJcu
MKalhK6QKccsRq084AYrJYJJj+89elY+M/7ewnf68j8C5JDphGSOJ8Kjd2rz
S7DlM8y43V4r5jFuIonPIqpMAON9NsCLR4uYS1GE7Ig4M/JgmTy0SLGSJU0K
sB/etiJnKHI7Z3aDLJefRYZGD4Z7sBq7CtqPG/vPH2ctEpMwEkifngHOYv5V
f6ctSzeTMf/umZjZakO+YnqVynimstVmSowOH1RiPUkm4Av+gwvLLPNbp3IX
G2JiL0UXIBjsgKTL66UbdvDEV1lf04/HLX07b0WmO3NRNfsn9+h99zcZtEmW
NbSAisg/Uhxbx9/XGMo1G2LKPacbNlW4F2aPf2kkU9a0HGt8YV8Dv/0jIrom
xfINzBhg6dCx+4qgYZ5BQm3BG9GS4/RNpVCmDNfMQsfspgxqdszW6iUCeFon
ZTPRyfy19nM4thIoXZvC3O/j9NIWDLaPubg5tu5I2O94MFgwOqpNKYrU9+9U
/saRUZ2p6YRC22MKy41E90FClamO+rN6bqPjc5qNB4Pdx6XEODWqPoDWyBpX
aufN0RQX++WPCKs6/gm6niMob91pcDdHWLmWWj1786f4rIn9avXgjzZkGbEf
/t28YgzWWNx2dIw5yeZoGwNvKlWDYJIyht9qwq8RbPEHlzWHrvV8jkiFtswL
COrIl8bB6hUmbmdVcoclBRIKfagUUyNcJ2HcuT9Kee1jKiKC7Sb++RhbtqqC
7ZRmJt12UvA9SFFJGt5dA2sKpLuuvgit6/jHdITUY3TIsaAIpjQih0l9I2NT
wgjKBflFqKenS4aXypGVfNvXbF8iz6hvIppU+7Szmmnhx94S3BMa+gZcMMyV
yq352QAfzRtHOrEg6cQV9YqV1RCt1mElMKIJ0TngCukuuvfn1Oc2+hGeorp3
en1KDk4HU6vwpMc7Gv6r6SkHiBgl9ydW23J2HYwZkmkXK1nUueNLUoo0g3zS
83FFeN2fKI8/oMLLDWtCxZ8kyfidPL6dR2RH7LWjkKs/VWnMjTO/3aVr1nUJ
A7D07Lg5BMVA7rYdVRnHUG8C06tMy4cP4RBxpElWsm7GDUuJvpoI1qTAu2CN
S0qCBZZlxhza6pl/ZScvNMeDfnf1oyPXMv1opoSWvlrK+l5qEU47PLoLIbDa
SZXpVfw55Rt1Vsn5PafjdxAk8nU4EGfVP25Tok9lJnVZD3cpbyktm/0VylT5
3vwRxI2nUaAEF3HLwyooa8UYkD1TIHDeuv+gDRhN8YU45GaV3ZkGbe8v2D+p
0JhQwXILd0DMqIZCdH6yDJ8uqZmn+oZ7Rhg182bjbWSyKGDT5l8OWMWQxHPH
FKPSD1/wJxlmiseTWS4hh0/VtH/aSRgEv5fZhVdDJChYOsKiUfkwxBWKJU3N
DuL7mkuTUJqCBU9P8NFnEMSCGgtVwI5FUIwbRG1uUzrxDM3yIYjeN1jn4CCw
+k1BVfuThBlyU9X/aFWpGLMRwHoFJS5jkrTX/Iv/XVL1bqUQA8R/WtSoY4Zu
V2ed5K45VEMH1Ld3CejfLTJKmGB33QSmTgsWC/oBakQwBkxURHpvsR8CGxfB
wJwKXqBwLfZWbYH2sK79+JH2nmsnCyfV0m4Pfwqyxky9L8398LGxAXxo8Gl0
o7IWveR/BwJm1/2mWXoVjY54oS2O/zhgPY+fcF8+gFbmX7iBaSVnqYRy3HVd
PV6eYNipb2mA8l1HWMXwCGEl9Z17LF05y9EV5AxO+1UnuMClnVTj6mpf/fpA
mpxw7G+f2u9+0I/bqgABxM72+aiEEnHt6tkDQjrIKAbgGqQn0zIn1DeGamEw
RKLbb3RLWTjW7a9bT9JmnVZquvJcfUvgIs/Z1nHYuPZEJDmwTs2JMYlAtHYN
RRJfJQXkwqiwm4XzM0Yjk8Qg1WrPhrbQuGFtQTgUD/KJbZ1Jy7E8wMFpfPT8
sZnjUuDyEXTUtj1Jp0/+bNHJDCVIJnbXiUcIMdZnjx3Mi4d/xHuuvxDNRqN8
habhKv9rhT7KZbuihKiOwEfztP7sNYHfnNlcufNdGQhpj4s+ss8BtbkZK8sw
laUBdBHniTaNL/qJSNcqfXifelaERgEMnYGsZ+JPe/Vj63fwLN1tz9xj/2fa
1NA5odA8Roe1/jqTtxCUIWpNg0mh8Em43yHUqXP2e8MboFh4bFro4todRnWj
VA9hFVB3VnS5LQwiHiFE8wxKLRDX3RR1MhqefVr5JXlIrA90x8qhT3pyJiEV
sRM8hHAzFl/4HEQkEs1bRfSqdZrNv6j4jSdQwEvsjSaflQOrQI993XbXqgWQ
lcvrAlwYe3E4rH/aG9FUcFBhQdF1Fy517R8ZZE3Sf6IMGu4tmA4ShqMOYZpw
oPfTtQEs7c1Rs62oOIJWxGbEBYgKWTIxaJyzBGrYJW8d+ZrP86YsAQr1m3OS
c/Fka3eobjeMTwynUAtE3dw/eVnc08HR/384TlTeFjElRiWvmyFlRDqDzJoY
lnw+puPTkxHM0hrRLpKWxbeqjXdNYmLi/46tk/TVl8bbLucXzfkYjVZVsIIN
DM1LOorsz3FOW3/lccCZ9aN5c1hXKofrUkpPqqJz0aX9ue0rFITx8e2FzbpH
0/2owV2VRWIx0/e954ACvlGvNjsnkc/BjYdP3Mr207WlOKaeebx7w2kM2K+w
vhAFa9dbPjLguabzVBj0g9jtp0BuHHEia4aJTuyxf3MJYZ4WL2HoFdKOD+5k
H5pqe8TpZTNnqxBiDu1RlYGuLK671XjbK83IFfl6mOSkqsMC62EAi3I810yo
aMAJv/pR1IRBCnwJ1QuzztGHYnXek+XfXsNKKVfkq0j+xgrQXZa5QmhKXd8N
3Ph3rBD9mHU05T4nELrANvBRgZAdGspdkcIBtbJ6Qt9iQWkb+fIiotkaMR/D
qr9iaFWoGi6UbpDeCitdh3OjBZ30qw/JVdXN16mEeViOy2mP02QxMaX1Cjoj
i8CdVBom1xNlYqGz5qHAY+ZKO0XzPYMjBXY8AEbhSV6kaSWbPc/keBDQsbYd
jxlf4ttjYP+keWpHSVcJcqy/Y/Pv+Cx8J5/tAXvVuo8g2UBzPmyFryZlgNcF
Okywm7PofpAlg3uYCnKpsRCU+1d3IR1LmOYaE7Zf8ukniu3yZV7MEaPsxoAo
xGE0kqqN+QdIDTQrHQtSvDogzB8qpleuC/2vlsat7rErQWIcvWLfKKAl9JLB
6OZh/P4OcvNezWj2XTKtorquxturGx8IWmtXznvlDskkGz6Z1YSJMIp5zIsn
Kf2Gi1u8WeKctDracZxQlEil6WYavhHRLTZzadgSxPIu//OH91p+FkLNqoe1
bA2M4MS2PaSDlzT977fu7ZvELxm1eGxZpmJlP1da/x5Ef4/ImBIwHIBUryv4
hPak7dnItMZWvnL0E0MIYHc/jbULqa3HJzpRcQJfm2cVE5gAGjiJJj53Mez4
bo7r80lpwgXGubWBQEFm4dX54+NwzZgQ73+WR/CEuE/Kn+OxUNWLfiQF7hYW
Z6LsCKsdxeVZfeb7Gf86GV4aNio2/3kaHdXOvMKC2tkuGLjCtsfKjOep4Wu0
7VGQ64noc5y5QVEoBBmMPs9yfGNB92dnuJsWq/GI4CKvl9z7WkjjX4MYuloX
yjJFYRiqa1+f+Yds+5v5BMdElhEo0rWuALqSLBD0LnRJdfq6TAAkm0An/juz
g7AYKZcMtkxhPO+pE0z+FNpXLazh93R7y1SVkps79oCzlbCGBopSMMXt9YKM
pxQ2NKNkEGdJxwK40XfDTmzbdYuPSu4V5GR4vQfCkjo8FI0ypiFVjQV3H9sf
DGXCbk5PGxkTXwtvV62Hvs8yTj14CnWKrB6kyxe1b2+5VKHgxLg/uJF8DecX
ODLgilm2ZpCavO1ntYv7VVysWCNmeXbgCohj8ZNylL9t8JQKONXkTNq9Ys7a
Sj7MvxGEVlBbSZKIDCZYSzKrMrT37LDrTVCVXy4If0WkKvKzvklX0re2CGkq
MsAfYek0uDNl7MeuXxSIjXioxpgigSaPQEwemQKHlVNi60DJ2NtGyb3mAhWA
uOSWkzqq3fnV2Jw3aabeKv99c8Ggf10EQn8liIx2vPl5ds8vvTHXgd3UGIGF
OLtQDmAdGop30+wIHX+N/TkhEQotw3XWJyaXuZkzfmwke8MIkAjoe1h8Iqh1
JdWg8pr9NJdEZN+365GGF+y1/XodZaMRkc4Aoan3f4OLAQR9DhjxCyrqKVp8
tWIT+mM1ChfrcG0LE6nhWmdvFn8hnS+I41Ujz4aG/O7QJO+FcBL8onIV0XMM
6qurGGm38/hQMB+bkqe9rAuEmKaXegy655Qfm+0RZhIczwAhOiBLmRYm5XUu
grtY1uZJBwaWCYAmmYgn0pN7m3DxCDidgraF51uuE570PvEUZc2aHPxGVtKj
BPmWcVdoQQAzLTuNf0rA6l+p/y1zKa17kIsH4XhZasC9bQzDVBBqYoE2Uiyd
ZyTdvor8WeIelHY0XvUBy/OcRJJx07eXxYuR5MifOpGBi1F7m9QD6Pkc+ili
B4Uc3BxXHsImVZrkSdPW5GgD9WB2Bwuzv7RueNm5t0F86+vNqDYDrfHDqoZS
TvwREFqjdYQxIvd3pUze5XfqSiRV38FyHPaIWqrvbZP4M2f7SLmT8NOKGIEF
Qg/i8yALlxxqtJvdXNfESDPSth+R7gQuTMhpasNsSOU7mRKUfopPiOrfDyL/
74gBYorHF88ez9PqiWyT8HZKDCrXlo/kzAyz86BPSts10/uFaEXAfG1NuikS
9htR/xri+PqJUIz4Kbd+HzoTeAfstKtnQNSf/bbp4wBiix2tEhbDCnnHqbwS
oD8fzICAHZw2Km0DvGkL63QCXoe7TFqKGwSfvF16Bg3DIarmAh4067qgzkkB
iqqwk+NzeNXfbwhV9Vk92Ut5Kg0C10R9CEghCRy0LW6eJP2+qNVG2tD8NBbw
QKEY2W0HT4w39gNRQKto4Zm/ciGASazavI4T62+ba3IvCLXwFesieSbCul+A
qIbMVMMwjvQQTdhuWd6Pft5yfs8qnl33IKLkeMC3CqbOr+1snATX66Fy7ekk
lZH3MqR7yvV053/kHlYpWmtICbQJ7klKV+3RvLbdbkURkd/Qs5rNyRpcaaHg
2R6BPRBii1+SGb/vT5U4I24QGLKMb0guV3ZUGc6ZgUP+irX995b5yiB51OHm
HKVQdgUYiXj5qH5OwRitVhTTIUDUYQI20IQM9/uZtbIFzwTiYH6lp/ArlWRX
EZBJZCrewZvBIMDgVs4GevAVGL6pH+dhad8f2/7dtiR3OsyDx6CElVQT0USz
yebKhbmR8S4zHiv53AAIYDptAe3XpUJF7D9RGHMHarFvc0lI/5Aor6BD2AFh
VRHFDIbVynMJZ5sctkD5RmhhFbwYl1Syg8nKRlPPreNTkwfwp4zH50rPN9V0
2vONvZ7NAaryLhknztorgjviz2dnrD67iRVY2UrWsDLy/w87LIL+Ex3u3OSQ
objTlhCmaIlnIFt6MuzpMZXonYHrKBXYRTNQCEeP5TGNA++xPOUOugs02xKt
yJ4GYFvRNOIhCnZVh1x2LS/vOMzi4TO+31d/+beUKtXCwZxXiMQexhUgi71X
5G5d29DulGs+m0D7OnDo/tDEAvC9RW96CgXW/PzpsKt1Znt56sCOKcVioPZG
2BBIO6fh7lMjTJzXYpyjWhkg6aSpRrxokYAePBCTEpLLRU0k20IupLM9+Jdi
AEkgc4Om0wU3W45pSR7m4i5aRHBPaNlAMZm/FF2aLmBPQcXIGtAqEpuOob5c
Pxpjx4AqosaStnBkf3UhrmvhT3lS5Mt1JtiJIXk4pGkWrlhnAIdW9cGWzV5i
NWQ5rVWk7wcmKA0HpC2cdynVFBQRVIHLhZ3OAq+OxUYgZvQoxhu2BvWCWyIo
MotVAtSi3yVs4d7WorzN2S4lFc6dVsaWHV1vKV18tdftIgbOcIWgKKx+flj2
PmNDH920Te8554FfWhoXDoLAAFW54VOasld12MyPviGCaR0qjzLzfF+NZgoj
y50/bzquX7Ais0tPzOTtpVX8xzGkRFnMhRdjyVj/lONpH1a7RgeNUSbflom3
i6/iTxVZDEcZDib9y54tMJ8QakBr2guRTSm3Fbq7FnNZ+JWs9I62T0rMKiJd
NkVqXckdgWFQICsc6m+p+G+vxR1DVQbL/zfdETqubFIs7YbDKsUVd3vH/uox
1lxq/tC2DSeffym4Is/ezs6k0THBxGYCJYZi8zzk0id8VYL02swRqd5bHvJO
rUEjZBPDk4jRnx1S+XF2+71EABW/IB0D7t5DFrmubsVOPyv/ZjFDFbKZ6Bz9
ZvM3opYAK3bBYlbJwHZVyNmP17lcS/S/BA2tIcsUB7dWBXqbxeG7B+WYiVUt
ObJ/R9Vb+N5s7quGY06QXrXg1K42sr5QvDpRJRfRw0rkq3F+8WabinKIjrC8
DCOZHLrbhoCwROHzTEwQLdq4oAdowuKrQTBqEKrsyhNjiTjjVyvtVQCkQJ0z
yz/lgVNKkT2IUQ26Yypha1rhxJQyNGo17TQSiUYwG8Ni+TsPeXQbMvqBme9+
xgNlBfjNmcwiwiI2AuAN05Kd4r5K7bogh0gxwGGLKVh6yRMIls7NnLmqjqnv
3BH42XFBQYmh5X4IUGyecC7fCP5ydNl9cg4efnXB2GaW5gBuo6OzBWhPQQ0v
tAkR89cD6bB+/BZLaHTaI/qGh03b/n7SfRE4e67rwqE2Yzn99ybz/9VRq7ES
owuBkXUmHBJzE/674SRC6/CmK7GsuUgPkwDWCfDSrLkhFm8xGw8YUh5GxiNz
DdzG6Tqe6BQYFpGAPfFfjyqEpIZJ9cUIOGi5bD+f77TPz/ENk7NOD9vak6Hf
FvdM8gCmx3Rn2uz1caoAIx/xeEV+BFsyySCaieX3EvXVRRam/vqxACWlrCQv
Xkl312CsnA1rKOwBhWJTJsm1d4jCZquXuAkYhK695KP3QN0ch+TmVqqrp+eH
5U0OIMtzsbUybNysiuE47KkGAWGcK/0ELYHXiGifRtwP/PmBcHpH0QMCQB5h
+24mcfNzvyzXipHkMtvL2XT6Z3C36HFg6xVWmgQG+p+QGfGXNdASvQwqQDi3
ry6q37iR8YJgKmkZ0oTbvpFOGh9m+4ZoG5dFQn3PHlc/1rrWB0+vORz9EYGt
wxGkB4k3DzcPnHP5gJf4+k9xzhjrdw0vf35qM5b5sgTcsNqiQ6NL21y6xgA8
WPpintlwCuSx9Uv605jEZSqrqjITCx/oJDipKNegBKMTpvMmmVnihxx6VMCU
FhErUb+DFLLvE9XKbuRvC9xcyd+vQrqpBTo+vVTjRrnU48LKqHc7Gm4x9nQM
q7Enn7jGp887mavaCWrFoGvweItP1GpzOgXQA6HR1oxZd/fnvlZv9b5va+7c
cThoKaOFrkwvCsJWTYbPBFwSkhyP66dSSsui2CTdO8YSRJxKA7R4YhJV4kDM
EG0PcdRMqKg7Muy1jdTga50YulJl8JCDyoCbi8+rg1WBzOE/cMWHeBpIMfb7
I5Tq/GoaAG57YAU8aIUab/t7EPLNz7BOLQoEa3YKy6cJJNGakN6/NL1gYcM9
e7/GpXSo6zYjOGJmoD7+PnxT7AKLLiFpFlr3ddRu4dY6p3OjyDU+UkjtguW3
Rw5a35+8L4Exyh56HnL0RNMpNOj4hI4DSmzlczOOA/7CRmgzINsQDUMrMpe+
n1HT2YrozcX72avoViuxQN+8pml+77Ic0yYC2Zee/Mi7cKNT73tcThNWo9L4
O00PKg1VMHqUxbwotOxaV+hNHRUZQIIYQsokq+++YagBB9Jf1tt0XA4//sm/
4jLDRV8zfZQYPt8w0sAsEcAAomuMdT80q2oAj5r0UQlZKYJF6l3jLbmz6gww
j7Fa2v451OiTvxHj6YnEKUXZ487eaA/QK2e6PgF4Lz3oSS6Cjdisrx52qQX2
AoW9qvCE+AtFdWibKqtSjeGMiGPY97+xUdzTR8mCM189EBivZOVsKgTTuToK
mKZ4pKEuyoW93Ncl3Hypl3xrBt8gPdQsAfYtrh5PtXSU6V7yuTj2hvvEZWXo
uABNToO75YdcjgsYIpauNr2Qzn+4CxJoT70LugvbJCHb2D/2l8tWKZbdk5cF
5lUcrzs6dUGBE3XpUuQ8uJOqS4yXGLbl7Z1xTpA35IH31YL2U+XW4Q4Lq/sq
3he3zcZ4YWFmXEdf/GnRFpwlCrEy31xmDeOVN+2Yd/8Kj4Ay6OLWUNFA+dbQ
Ga+ubCDPpZI2Bcaf3EpzDK/QU9VDfC3hbngiI+LdiS3YqovGbM0tPmOfQcJE
s+EAT/lkcDyN9O5x1NHPxTsAIbkrcZnnXrGkoXRYERlvUF3WCmLhY0diHg8R
1070CKatEV9leTuXy/VgskVbgkk2ixSXvcYzvZbsiw/NPcyKsIZNLFOMlqE2
erVCzoQoGmxUDuLAn1jOsKkuJV8Q+SgcKDpIqUIhpeHJBARk0v8Pxkj1wZ4r
UkoQCCZ6V3ZPEix09JP28oCmR7wRca62iD0TQHSDP0BPyBPhlIT9di9i1oDs
AglzXRmDTlXWFuUbw9Sf9Cntsuc1Jq8mOJmYuMnGilzeUy/Wg/RN3nrUHJ31
95T0R8uYQO0yaBYk/HaEgK6u7wk5IEg8UlAgFGUcVYCk0zIqlMVWfhUd0c8U
mHzLL5zkIUD7leCIDtyDWeqWOtnPDsh1v5CF7Pni2H7n7ZN/tt8/BwvdsKA9
EuVanrmeKEnzIQ21D8D1LowuPex3m8Z0UAQF0jp2DQ3dgVUky04iX0N8HSv4
W5mehD7h7ggwePXk+7e04RBHLhiHjcH5PgFdxVKcKtJeffXPYIwn9TKGQyTX
rLANvGML/YbEAqrs/HWgaoN+c8vhzckssn/4GEFyEc9e2Ys+ZgMoCFegL3qY
zCbqJVj2VwGQeieNOM5iwS6UBv1kdCWzzvSUrIZTKyAK3aKDlTt7WuWUHE2p
VMHsctm+0m2olPGdmlxxoMmjPZ+BOkTX+IZy9teBUJUFVC3GGaWL+8KvlvOx
bLlIKGTkPBof8JlxrqikGglm/DI32OlNfhuX1gW2zeFIavWf30T7zQBFDbRP
gUTLqRTInnvVNw7X9Fg7IndSCARAjYogS8nOqqZ5WnJABuSo+9hyanVida1Q
atodBnIbNrH87MKnVctmetQl4EJ2plNtqex8WNSgjuaHfBxYFPqqKyV6hst2
EAc17Hx0ldRFNwypzu2fZxGSZEUBhbsbduROm2ItHRQwaRH48ccNVC6n4zoN
fBsQhJPG/yvXCQMpaR/1fxfwfdkI4aSDu3LN3B3KRudygm0YGvDiqCDHslIh
J6mID6SGCgxgDsh4yb6aEbzyMGO0T9xEQm0prf9NiP7PGSqAC/FpMPLO1W5g
qqxq/vtRNdEh+7U0+4J97VOt6HBWrfHLN/Y98qg/RbDdjMH9hJj58gbE+Wv+
ASMkzYbdOE05WodKdQl+7rt4eXEguW5HHCWxY0kKSvBoALCPJwYhbLFwcEjM
YojTUKP0RUygrv46atQ5e4ZEQ9PT8/RLg7lJW2C5IPT34r0VqZnGHe+q1N6a
0xskGw7OJz6siQlgwgi673Oopab2uTPYvpEJ1XQTfraB3J1TwxSrIU2PMQmx
+9SQn7V9UVeB79iZL7C0CI++vDPd2Fl/++BU4RwynK1IF3TbwRGaZi/WzlVR
A0KPrpyPFzYqmXYERSGNWXiu7k42+53NE9erjYMvRDfoFmDiHgGKLHKTcgeS
QQB0dAb+SomczF/vGVbjwt/7gqfppGLrxn1Fzme5Pw6QVL50F8F+1+jpT3yK
YWuj94pWs2bhCvAfqYr82Y6e2+QztsfyDaJgovinWqDzPSeAHU5vKVr69NX9
cwZqv8+o3BFZ0zdVd864YRvQnRcoCuv2W+ew3jg8v4AAjq4J7kqzzw27j0iV
dQGd6bId+mYg+hq+vNZPWVF026TIOBUl0nvcMjVUS3jYf25DyW0rm9mSVGCX
VP2lztUylt4xKqFaFf1LgVbFoYglwHXD1bpwBRIX7GrgudbNsUufyHACikGt
m53EPZm6cUFHOmlj++tCrxScJbVyqGoTSMc2GTaAZu+ClxHk/SpLc7G9mg6r
fywoSZjnt+Lm6X+gOl1vC62gHZkg6ZrdPLwpajSL58nUbgxZYrg4gm+z8hL+
aQMuUT/jTZmZvs707Dn6mjLfMriH3pHRAr1P+ZHsHu1hbB+JhnAyaAMv8UqG
EytKcUkmjB6t2Ezm5vVu+jaQabzkq/H7AfqvKbL2C7XmmlnH68cnspmdTPju
K21vz2KXhzokHfA8aE7DARPkplqm3iG8Dx+4oTqG1nycb+LF7CTMkW5AKQ8k
HX2wrYkxe6YLDtvtZ6c1Jh1FPBxJQOCiuzess/lnwdnHLFJxy8NEZ+tHLBmG
BQRuNvwh0tucPL4/pjF5H4LUAluYM1f/ROs4JYzPPVlRevCzg4Y/2g6nQKEN
2Dz7t+NRkBfatFD4Ze4vlgWxbP0t9diEmCkxs9kUrHvXx47vQ+fGqFvHZLNv
2QjbEEMpUV+MqNDyEE9Dl0DQxKqRha7vvU0D6JJBr4/ZFPrZHeZfbLClkCcz
uHU9EA5wJNAraBw2TwwRvyEhNX+j1OBzY5tdqRYgBptYqAkm4+uUGPmZ229n
wbIMk92ay0GJx7mS/mYJpK/53kaIVtCPy4MfBgCWcwPq5yPsaA9cJPUWD8cu
17397kCVGcbV/e7j+rphBgmhUdhYZi/o/yqbf2rxI3/6Y+gMAyIWUF5FkUEd
PHqVMhOb2k1+jYtNLpiVMCk8jAzh1SkDh2JcnC6EwsAets8jzHiXXm2zxZLN
SWURKRhRV10IhnACS/QPJfj1XFyyTIcD9aq6855Jiy5T0hz5rpYPnWQMoncD
s465u8Fv+yA8hWV+2sOh43BI03GeJ8U7hx4AkZbSWZk8bGCY2bsC3ZYTDSBf
muxA/gQSZ1HZq+3dXb8TQ+MiLiL48tAYWLq8zsXSnoNv7aokf+bqs6XpyQIE
qQ0x/sqI5RVnoTKUVnfDKnDGSC5oAMIARq3auR0i7xqQdfHHigxNq3spyqWE
6+AeNz/e0ejMBI95pDyrS7Ul2ijoj0JmjvDUt8yi7b4DakYgoxSnzMPBaPNw
F4aOU1lYwDcMrxODIkkrm1c4c1YuprVlY2li0RXdckBmQyopI0Z3OrIXNiAS
j3wqkZ0IBGn6UAPbIYlDI0uIj3gltQkE+9paXOnutRPcCXPyuJOW9cvzCObJ
KyS2N3GsP/wgziFvT219KFlpudQscdw2Wtpyl81sghBlb/xioey3W9SbRFkA
unNar5PUHmiddcgISVbwNylLemNn488lkGs8wGeInthSYVj9Hd5hznKI711G
G4UWPLwR2FIpsvar5rXGM+1ZFRVnmnIsminc8Qp0ZtIHSUY8lfQhefiLKbMa
hb65Shiz2M6jhD7wMYkNGaEoEFcXsOvC1ZcyGfJFOPXTQ05ZtksrHP15CYDY
NQDWRfBo7q7nS4wzCyNqP9zGdL1k5l559IxoPmBuu3WM2Q/doBChAi7KxrEK
RDPN/ekA+lN8YA+kzr4yDssdPNQJ12qoG4kecdyUvgKtAJGACfKNeoQ1vB+M
AXRoraiIwqcXDWkZHbxLuBZbByNKRqw04wB9P4g6D+B3nK1Es8ROoADwE5TZ
LkQWd1zEfaWC2bDAqg0iOkty+IK2BSqi/crNTGAMKVEOMlR7xkLORmF+90Zt
nsKqaGyxk2jMNmffUy7AHgH0SPG6yZJqjunS2znaRACgh8I2Hx1q3NdMamUm
3yQoz260peQmRHeFNZ/NAzqR6iupXr8Iog9M7Naya9oQ0lCzUrAwrkveu5hw
xRpDZWwptDXEN/AdqCOVCNvqHd6auDG6hu85ht+sEn8NFWOJE3IuBD/9wVLj
kCIE6PI5aGSKs3Vyl01gWpi7HaJqirlNggUQKuVramtitl2t0dbg1bCrhzoB
7eTaKSLAHOTl+vtk5/i2d8aB+R7HLgVEbLxDC2n1gQ5oPoxJqETYYuS29djg
Puoxc10og+FwMZFtpwJVbjHZxGYm1crd+5lX3yqgvKu7dA4fgHGAyAK9M11l
nLrRBQ02WJX687APEaG0SqIJaFgvpoVFwKfYwV65TW3Qxj4fax9PnP1wGFuL
4XadddHpvADcO87tqeCNitM2PeZ6evmpvX2KQfJqjxdfbhM+sngcjg5bVtGP
WxJCgfGK8suPgKQKIrPejZFAAnJYtwEWSk6VHDF57OerzzLmp/lusRwXEWiQ
epUE21YIMw8gqr9pcfyl3xaLRKa9Bb5Db+QoBFjptLrokRXmKzGC3JtH7gD+
+wOhEwMOVghzFMkpJmOWoLRbAeLYaR0orVQ+OJgDK+jIxqWoI86waYQEcTW3
DboySFmw7+jOrqrQpbNUygXWTi5wWTaHm7EKJ/bRHmsv9uVMU4vWbhcSQzR4
R0iPaTZ5/OYLtgXiX+7YmcD0FOuoekHstPpaX7n/tgc8MzYYcXKtUygqSFIk
TaV3BpYeUXx7V4Z/YS8OktEmupoOV4e4/iymLeAsClh0KoN1F8vdA8XBHO4Y
oJPp/vQSmLa77dy2Vkh4l7e3W2qi+eEFXARgecphYR2t9hke1VcrfgNxmN0w
M1cJbGv3Yuop5U07tKelYE80BRSLKoYHkzszXRqAzbMacOozrpLXFtldCujI
R+GG2rlve0TsW0/46u/5OQK6D040PBv1ybbHMk8Aae4O5/iOsuinNQrugvQg
NX05bXY45nGNjBro6AQFE7zFFavh+JGLX4/tEaqensChtt8ekqVwjoJQmYa8
A4XJdK58wTh495pOIfaY5B7JGhljBBTJRCKYXqdwfq9Yji3Ss2R07VF0q78C
976obsFV+Yix0VyxXVytAX5cV0aJdgtcY6g08vfKlSLUGHznjcur2OkcyN2n
+T+Me3IOtVTED6kTlgoysQw5ka28/N1V3d5zYXvIyG+6+EPU0FUcDOcBbZZP
IrigN9an5DjHlmRr8oOBqqhVNyUUs/+0rse29l6m2PzXEaLNlxaBJF1bqvZ+
FLQss6mH3qct65TJDjnUZZBEVrJtCEoN39uuFjjJEXUtia7+8ms9lu+R11w2
MBVDyMcCQfkOnOcATL6GlypfoWaXCworgrFIn2wj6epA+0MzGgsVr/YHY6MD
iv/SiP8nM8IaFvU+Im6FRokwzFWq3OONqccE/IJ7ePjkHM4sxIsEwb0YUwih
TFSkjnZkn5SLVZgUG87xaVRhpM4bGxxXHL69dFxZEvyBZgs3KqbWrOzWhoOW
sM3tyipnYVP1/ihsUUdjOCCZjYV5Ctc/rXt6C4ntAnWPvR6qJT8MLEbUIQ6o
hBITh03kRRx/IWqKdmysKuGqvf97tiFMQ5S0ggJkCaOT2cxPjjcdAOiqRkBZ
TlITSSd9NNZx7ywvNxvFqDqAdd3sJT9r/Ell8EDmNc/Wj5sKhoS6vRDSq1L1
TQjczlcgX+lXPYqeXEU+FbW/GSHI4WuK0ZpOMTISvKbxY24etvhctPxly/A7
PMjFhOQhxUJAYX4oMVQNHlGP7iw4PUiKyJEVvXxOAsiLQvkE8nuw4/ahvc9E
u8BiiivqmciV+mAjucEX7YTepBsBcGwHN2jMACc6DzmgUkigVxHyWP9r1f5L
IMguTheVLUNj4gwLPhHRxYWmC0sxk+NR5fYGNbH+HJfXqC1SNdrTMTR3zUHZ
d9zzi+tJsFTw+1vRvYHt1sV96FCjxUG8AP/kAeboGkYgl6oITNtcr4IT56an
Zg/YIML/cvJo6WnakQrUTJ2AExFC6OBK9LdudqhCwTWLTMWC6oaR5gIFxHfJ
PXSXyDIS+wbaEuQb+CX9shlWgZlINGubDHtfmEXvw/By/wgfChic4OEnZX8x
kK06FQm9w3AovJ6fBA4BQYjMI8paalDN1ItJ7AoPpZhMCIyT1n+DNgjaNDtx
oA0uurL8Mt0Zk5142Ue2S1Iz8Y8GUzn2hO+tEIxjABgv745H1z+CfbjJEANy
G/7mGDWfu+rF8JBiKj+4qhF/Rls6radkcqcyn6b/MhulEcabskYdEda6wXrd
8unOVgwzqkplbclHSMZoqDVc/TFlPI16s6CKM6Jtiig+kCExZZWnUD1vHMIg
vkXw0HcGGUFa55fmzTAOd7Us6FqXNeVr0Xj8O1xv+w4pEofImhbdtFS9DYXO
6s/5WOU969zwvLHWHQlPQqALG98KELWGJo3+PN0bjW6a39tNkME/fFH+EQIS
nw11FZAVUG+QAFuYl1I9X8vh/sD3zFqOuy0CU60TXZyYupr9r4ruAxGPTb3s
VE7Tk4+dIaGTmpUmZ8vKPqlili6ydvZPyzZY4pjB/1HGFv6QgBQ0/AoJrvE2
vPxzDSL/D6B+HaUz17Y7eaQ/cmYCbG1+XwwGbKcpC4n/JmDIBTxkdXqwn8L6
wJesYEEnZu/khSX8k0P5rZEEpMLkanaFwfnTUrh9NbceiB31th0y7IQlErS7
tvYhKr5QnOQkJElkpg7CJOauRNPREavc8dAo28+a0dU/93pJqe3/hLN2TvGD
e2WIYXvmIDeBeAPcUnknkW/DBwbcKqfmoZqMtKGTCn79RJ4VLwdMTond00eE
Ik5TslqzwEBRD+8/E1fOof6hXtPKRPXst9sFPTMEUBRq3BAvM8DnUIybKROs
Jl7Y3ncFV2rTJlPUL3kGtb+YqJ36zH78CAs/x+pLIxUd8z+2XqRsuEQFgB9o
kF8c/piDMY6BeqYX3e29WK09QiNB90flWi1Oko/hyF2K6N0bIxrCwWQvtjYc
dfSfmgTIggx03Rn/ks1iy9web/bRKvtGt4Hl8GwvmfXsHtm51cccA2UR/6vc
dSX6Mp5zgZSiSdXZ1ScxXMCei8nTYVq44fEuVSI5jPOE2pWNGOABM2PrJPXC
6ewSCBPAlKIcopS3kY80mAlg4U76fLpmqSHasfeuO99cPBUzCMsCQ/D06tpp
jpCDpw5urwiXxJu3egwEFf4B1DLLE1aiE1iE2cvolqriv+jjAQYIFp/EgaaO
KaJDnqcj43VxeRV4j9iIHejdwZHs4to7zB463irx6N7bbq5/m7frBU673AxP
lJdqWaQxrS++xJ5il0UBl7oZJeExc4+gC7y/zQSTXWe5B1TW7ZacfUm3xBti
IY4GP/rGz4K8gMEPGd5CXnvltjHuixEttgFofb/GCejoqbmnq9SbrVhgwVi5
7kT9xeBOPG5RFQwlVSDmy7Uf61ykNMDMcJsCgndsIeLKybLvRo0Jh/Sx2vbx
b1hrbzwZiLLPxjlsJtrx0LN5SZ/jNvaG4nrD6awCJSRtZW4QEgu7oInl5DWV
jSynHa7K+0Cy9B1tg8Xmffdch92ZsgaF8KXje9BjxFr0pk7gnfIaIF2bakDA
U8mLTf+/mpQq7WCPJ1Y6QfnB2i1CYIrxzFLk45KoI1pU7VMVSMQY49LNkXfM
VvxoEMXpFmUgO1NU85+t9sb9Ximl6IrL+2VEMykK1HJM5qqI3s/DuRg4CwEr
7NLz2DGJPXJrjb4oF/O71EvETXxlWbhY2ba1Bl5OWbNqhWSdJ3bRX0VLFc9c
k7lwzZlI/6ToBhu9Ej3AwX/EmmQE5VJ/ygJWPYv4ybiU8NKDhgrXWXf1eReH
F+TGFEM3RwWV1uNrk2ZAUw6Zzq9EjwZbXlKDx3cG/XpXGRXOsQX54i6fZBhd
2s5ZQGgtIxEZZpZS/Wrla4JPY0SFVD7q1k4ugEIw14oCVOTVbPN7BKK2vUgF
CH25HK96aLALtg7Q5mu/ZFkbK14sgjIIrF7JxGBLe49ycwkYqX4EmFL9Ot0u
mAxzF4sWzW5N9171XrT5drdVXQWIA+G734y3TUMYas67GuNktotbAQBB8ZgW
84N3RtehHCUv+Pxv8rfNVpeNjfyIPGNss93nEyZqbb7J6hGTLXf4i21tFOta
16McXkCqUwyT5FN4qKqn5Jaf2mhxGNdFCqV3GVQZSOOaVPI0UhqdTDwo3Uiq
6IMJDiDJwacJEenBMZjhi2uhT4Iu/0FTo8mn8XV4bosYlYSC+ZvzAQ4rVp3g
TkRL/zYPpIxi7SrREVWUmrdoiakbBmUHeIhgulleyHKpDDhWkMpW7N89DoiA
Hx+WLyu2SG4aHRVktFe1bIdWL8MAkM1eLK9fMncGSIEaCMXoPAZoZoeg6mza
Upw4clxeP8G5OL5xrFagcVthBjbSiQrs25qKFhkYT+YibERsbsn2J24IevOO
w/bfeLME51b3Gm7yXge9glvk73N6m+kbQpLZKnLfxLApDzsvRW3M3p/kL4lO
uNy9wT82pBJpOAM7M56Yd/tPoJKDiUZtF5dKueGeF3t4hB8bCYfKfkMUMYBT
9TTI3Pqcz34+580wwT+76awgJpDzR2b/SnKSU+CjbxJgJfUgAbDqzfKKQe5f
ZsX3gZLiqi83IXxlBECgElv9kSKffxBJ8tW74/ZUU8WxmGEbUjG3T4ABerdx
amWcDvcEhP9YXdQ/khdNvDTtJb/BWnwOfQlCvdO9dkTGCIwArVJigca65fOW
KIRWa7PnJmxbSh1B/8ZbdUhzj2eGEln/vTHk0QDOHyfPJoBYIv7OqaSkI0wc
4hkctr/Euwl8fi7C6Mdn0+LQiowi0ErvHO488UujuGrwAPK6XPnyUiTT71aF
+B4c7gez/80ht3EuJjVXPCowQ8W3QKqvgbQvaMGneXMA/7XzZOAwWpEuo1vp
vK8sa7o9HfeOxIAWrUtFNRnwHFmOPRDb0mRWQJnH2l8LbwpeHnfmfWzeWRKf
hWbpEvab1AL3YHzljKsCI0dxh3fzgzJAV8H3jzhIXjYRdI5CKJZtu4OjSRCD
Gxa0PQ5KZ+wvJBUkZUdc7NFsIQpaWLyq7dR2OLQWOfuQts3i/aHT446fXJaV
XwZmtpYqBoSc3AKZJCur34pN70TGFpzcWHKFeNSgmad7883qTz7T14JROuWt
5E/3gGElRikBWaeBXnAnXk7eFnWya9cJl+6+jyu8Qj25v8N7ltrFe2flZT1q
Fu8Lzb7WC0CIuyG37W0anllvRoPbogb3sJPcpPuhG7mkuxfZ+CsiKDWjBBAO
5T4YMOZYUf//Xb4mJ81aX/aMWO0ZeZTI7Bx6QRniSbD8HdSUE+Lz794dNGbd
Idktec47KOKOVbpkL2JqEU/CKHcsBXY3J+XcKuIeDy2pjdunXWBebzAiU1eX
gAHbv893USG7jwxHt3wjtDQIUxZZUWCOkTZgWyZd2D4yyDSWFgoiH+cGiGQI
DlUEz7UK0hvEuWNwEwcpaZTZgLPHnRIrwj5vzPZBWkjphs3GGfamnfvj4OBH
lPereuyOVqnkDgNPp6VYjlR++RmJkQ5fQLLb6eZybbdOgzF5ocltTV1yv/5U
vRCl5Ap+eVdTQa0HO46Z4sMIWMbcmnZmV3V3laLF/q3jjZl92OLAeK+xPxPq
1TaAuvM8gUoBTa8kJCQpuvAvunEmB0Qw3cWjR4sMQEy1X5IZx4qVjIh105xV
S7XJah5Q9AqIY7vwcpVuiglZ85TPZZViHaqHaB9MTmbe0Lq21nqMhiSv/AQf
hY7E/uKL5DAGMDsQD+rgYGIcyfE1N+OssV7IxJPp4u/eMTFPOQEuaq0HTy5m
YHKCBp+lmQSbjG0WGnFPuNC5KAQEeDUzT6AJUdgBE5IjRQ5iokJjpzcW5eTN
+ijady+KICS95pEkSKx06sJPm9OTdHt9nh+E942QUACDXFohw/B6NEeCG+8T
ND1ZbkUrckJM5RVPDMpFYMnmRbF2hPRLCWvV45K+vqNZQtb4pdwO3+UklJ9L
HJYt2qnuZTSwgX0hFsqIi7yG1v8Hj5BoyflgGslrip127pmLykehVF9KJFzf
t3IN2+plZ2Z4T63SmrX7fcyj//Y+6a5nWkaHbLP960PnDl6DBn4lhgsEatfX
H6Y4rB5rHBbranAn59fY7qbLaMeprcZlvFJ8bgaI4YM6nK3QdiaZKLP2kHsU
HDUN/+tvFdcMWUM/UzkP/hOzAmeiMgEZy6zgiDjRmZrypamwsUzdUwJqTq7C
r1N+l0WtoESMYLr4i1UKXbUDXqivBBb7VxRKDZQywkg/ny/tLGLsCQPPUBIf
JTBNONMpGZ8HHMXJcAH1z9j/Zz7DIkvTDXHlw9nFl4MJbVjaQ8uvpK6D3Q4W
8PkDbC+JWuJ3K72CJTv6tlqyZPUkRP3PdO5BT0eelaJnCudV1FsV6cS5SQZM
DQ3RzDdg46eRXYlYMqwrrcu8aRqx40C1DVz3K8uPxDcqD7nUGbBnzrWIdFen
ZrHG5xaXx7aptS7i23NZVs2WtlPrQqssWlZImhZEv2cSGnosLQtFodfYMDiq
iMVhVGv4d+m9Wn3g5tHeD50dBTsddrmG/OokwYnS3yohQtd/IWFQd9Ds4u9i
PXhjRVgNss+3YgU/TV9xtQPRtuym8l8S5OEk4WiTBZK3joYGuOPCN+SFMupo
Sw50gLJQCdYChsMoJnsj0lsSYT5igO9tJ4P8U0MC8HLtTXRB+3+N7rV4xEmP
i2aJpg9ZNro5LcrW9GgrrZHVcmPf5nQPBFHa9xh9RVQgAoUIdYvQqNGW850c
//JrjBvYp8c0BBvCOKi0FJL/u3Cd/PtpGclZa/hgZCgMKAupRvj+axl64ygu
vIaXj/gmaVmUSoVswTjyyl0r6sE/kveh4+8XZ/uZ0Or0GFVOIGrJMAD9hzf5
YFm9OSFnASL8eaJgod86oHzC6GcBVnAxnBtybk/ZxjGHacHn7fA40kV/Hxk/
NsCRKlgyY6nZbZk3hJaVcmjmYvc72VDSPo5+eEyqlxxtTJnW0AwKFB8geXc7
eInxh86CxvkendaNQREePNJleIDsCOpXobg1h8F89sRLJ/LWHK/wjOkkczBy
88n7MpM0UzJU3dusIsBv2yS/9KjdOslyZQ/Wd0ee0a/T6g0Nq0iwk9b56so6
kih1oM5eG/RV/pXmuIfR0itdSZ8NztWvLEHDFlAF++qwm3/qiuxuP6AwfAjF
ia6qxgTuXaERcaB7LInHXYDTkEYMu1IZ2+oOUL4LrUOXQ/5SxlJreBFKiJzA
j2m/381vhF9HNrK8LAhz2eqje43FWmTHFsvh6dALnhMZ2GiuFOvpuaAuRiDR
DODyCtllr2EkfLeOx7h0FnKSxcM0GfxcWuUcweL7LYZOHiqY0Im8G+ijt0St
GHnkaGHaPVrVnrV6m2S2ECXoxWxhy7ToAHdyypxTpAkVLW4KGTbe7x8YacYO
2aOP6zNW89j2mi2sUJS+6VbTwMtSKSafeFJ5zEb+pN8Jxqlh0r5BVCbw0vUb
ysJX3ZLlyOU7MFfiHH8zyfsbUGgz2sCD2Yq2sPPrqAP6UX44XLweYLP2DE/m
hqmS8lNoP5l6L/ejGsEYuUm5i2RicsnnC4/sOx/uNIv4QYtqYrX1KPWJbmHi
SifNHDufBukwcUONjeLAZFr1rl4fm5ZFKMTtK+I1dTH434m7qkK/h6wlorKt
HWVbAXNFx4azJrTSUXrv1Vm8Li68S2TqQbVP04b9D1K62QfLXdVkNhAK0VKQ
XrwhBjknGCfEnhRdPjAKJWrnW2t1q6iEr8xoYmMkbCCWJTvklKhRzWVkL4IR
+x7bgHb0eucrLF4RgqM4vQSet0Ao3J2gMos6Qo50BE4Fd4SeOIGmMwxcg7Iy
RtnVnRnBnMZMM5TkPGBa3+mUnBxcy/xH6VqesBlWTmGB62/SiHjKlBj7s+X5
r6nwsOcy2PdgSzWsalCheWZi+d5/RLNOl1o+rt5xndKnuP/YaAG41AnN5D9E
bISFKhLx44uONwxrQzDyif5Tgn+KEhglLOvUvwBPJBwvYqEi+qvi0Onq2+2F
BwDXoQjz7SW06EKXn7OL39DQj+y9zFJHxMzLrLmN31EbmUdMu8bxQTozNCKv
wKpdotvHOqwbSJNve0L/+zhIODmbwNN0fBa7iBXxc7azmcg+izqYGS3HNwm1
2FM9YprEG3A5fUtwga9VLWZF9DktZBXPkruLF0FXEQ0os6fSa79bX3CN6gDZ
I/eYIfv+Ejkl8m7EULr71IvxL8HDKGUPFfasTZQ0Gt5GMcypYezZ85N120La
EwagCibP0BKn0RvzHysT3Z4Q7xAZDgCrjUfKb0bQhismW0q2D8CuNGMyi5g/
LPpQ9tintlc31UqG/9iGrvGlS1X6ZSjyywN6b1e2U+E9da5jr0MmbLOYYssE
+bT9GnbNPRNr8sG0uNSre8NUWytQxFy3mbl3RgIWfI4XEf5YeTbD7KPUHS07
/q/E8Rd99l8BLr7zbF9wPwmVcCE2Sh/5K4rm9tmmJM/0fKKXgLkizIUuHiPD
xnIDppcCzBIuHZw3QoBEtIiv6ja6bX8t9p6s5VHwjfVAvwzkQPFwr2aYPxK8
DLX+hMJRspiTKKEGKvHjrhsjhPUyn8YWHGeUgsGO537qFo9m7BjjLYTqPWhQ
IQwkdMXXJCsJVjYnBiDP5tJ3jndIGuif4g5RTwiE1nE9+yTqXosL0Sdas2cj
Qufy5B/IHgS4okXdMo1z6v5U/ZeR3G2VW1uoYm2Fe7NzALInyhCbtShoiy0v
zB3NH/6aoKeptZjR0A8iFD3sUXQiGSpMK/MJMp5eqOqWlCBJdzHfTtrEHK5F
6E76MAECw52l08BTdLLwkL4jBl7VLBJEbuQO8XPBulAhIK5U4ADbWQpBvI7h
e9uzc9e+QHcE2+X6Or8CNWmuTGWn6bx5OkhTDc2zrYb5YmnT3X4bL9IFNS7n
bB8LvhADjTcNs0fdKgenxBL16CKtrOOX6C+emF2yF/wgCD4O2hXl31AK4ZY8
Trjyn2zs2z2vpEpo/NXm32gYoXLnmlLcHflv1LPaf4L0MW1H3nMNkbzzfJvx
vVcc+TtoIOf4tftQjTnhoTJRNT1CopMlpwIBYCrs+okYp6sgOyM2cY5Q3++O
eEEs4xofEcDhj6r63P72VAS/XvntiqOAmoxwEzaN3fR49ASD3lhFuy8zmiQ3
qQ4ydBKwKtLj1zazaQi81Fw0DMIOBy9sBPf7utunosWiAk7Y1/DCgVrJynFt
dcj4I3/q3Tsp+Sqz7RL12AXQap6/5pj5NoBpA94Os5NP53qCTMQpfSCAhjRk
/A1Wrzd3KpbMocBgMpwW3tF/JeQVRS6ad0hhPnP6N1js+ozYxIdvHCAObmdp
StseyCMQDHUUvxVi6TkalJsw/ka+Jq2Oqvsrc4YOMmVb2khXd0ZlM2jF3uxX
e2Z06w0XxXRx+xGP+n96AXfIsqytFH2LnErdeT5warUCWUdm4kqBZImSkqmn
vXJa+F0x9TDKsEFlXBjfqaxcTXf9W7pLePNjLCxcr+PIsuMaP+4awDBa2BWm
nw9LK0UW4a4TSI44Ar4Li2gu3bjbpe25aqdF2wjwI1XsBupJ2xKdNEoROSwo
MAi3rMgih3S5bHZf3/XpN6WCsZPMBmP7iS2AVdHlIj0g+KJXMUpTJ7lMK01m
XRSwLjIfWMfoVWEDryBP6ebECZe4rnHI0UdGqOOi4PqVW3AsjRux1l093Mk0
/qfy/W1UUzHqM5qEXXmHxacaR6DgizVyjW/lXnBiSrZsgz6RTZDVp36q0j/S
xgJuKJtU65yPuIUokhvwQSVAsrb34lZoK4TO3C+NPt5wPRE6F1Ds11UNVMA/
5bWUguGpLUlEQj9d3NMwKOiDecSZdF2wq8yP1gWkB5X+iqb0q/Xm5EihXeWO
K+yld7K2Gv7lzLM7nuURyUl9puc8mFTAWyYzIuKoDoe9wFL2nxlHVNjEgDvt
BjJLjGALxLPT9o1/Gy2+RMiQ+jZM5iNPVvTshZQk4rPkV7eNYJ/VdvsUdF3Q
q4iQwezBhrejopWAId6L8v7KZMkYEi+B6/SpVTPxfluTWmTL1Bxfgjjmbjag
n+xz0zfNqXd11/yG4E9zoXCgTPuVav3Y5yc905dgp2NSZY1l11f6VksSu5go
BeFpd0o+kMBBMDR166bn2dM5cUfV2mdVyGA7TlmnKgvX70qXOjPSEFlwuxHK
5Jp5bTFWc0n0KgDNEgLr2DapQ5w3WX/556LWvSJitRssdskSEdkBpRWxAFEu
y+QLD+Bz3R/03w1OeIBRdtZHLNlClpS/e+68LqFh3hNl3ZkBX8NkUHk5UBCW
Zf2AOyR2PNV/q8/s72XXexrl+uc7IAE+VMV+FK5SH8EaN079YefiK7U3UN+x
FON5QR7eFxOseDUdbQV9+gpDfl0pOaoeBLQoswKAwpxcwGvK4/Tg5umI5xmy
8F7GbhYj2MinGorGAMCPI6mDPG1yETqBel3D4UDbDXD+pv6mkgaERG4+KD3J
SkqZwfowDtUXQobKhoVomzWT78cWbkuGsNpJjqo+kQSG40WW2cFwsHXJWdUE
AanaFRPEYEiU3Y3fpEJsdkes3pU77jdgl5qiK7Q4qhbvfXA/FteOxaJ5lY2J
T5/lJEnMVx39eo55hFDR6rdSdVX0aD4LosmdbeNUZTIZwbMGDsza7myfSz7a
Ak1TybgCYvGV13CaxDz4MXCcgjloqoyPTLTjaWjoU8r2aibnlVj8K1StHG/C
8+F/dM/1Xglk5Gf+VJTOI26d0vKHlnAi0/fiw/55qq1Qa2gL2D5Tthz9eoxL
lszJ0j7NhuCEQxn0MA+IJk+5j5uzp/8/Bl1NUnEJi5Q0CWjx8JpM4PO0ZtXo
YEqnxdZ4b8RaNYOq7ES2ibA6MhT/Pqkb2oDyCTTcve+hD6vuz2iQBBnOTtfg
S0eapaUXn+ZU4HHqAKHja/rgHnq74vy2Hqb/P87JLeN1VDP6BtXmN5zaZE/I
25M+MJ8jdq3VSQgOoQIbrQqn6mRr9vINudwRFcYNNZm7S4ON7G9t5VMX0NHA
weuqp/GY/Ckp11Vu08jggX34kaay4hTFh7b/rpNXT10Rk0OE5aK2cBsGI3DH
9TpRMfZihXl3IeKmN9+97WAXpDxhCqVsgbwv0njxntVr34ilH6Y8Ss9qEJWm
MJAomIAzfSVRUHOM9Th9ihn+wMgWrP6F5WNMNuhcHWItcQhR9H8D2XZW+f1G
n3VxRbEX4dd8h71YTIHPStyAKvfeq0e/Gzm/6n0a9a/E3iGjORjHNZkvfZ/r
tmjhCff+I0tzUhsLxJT/wg+CJM9zgS54wbmqJYsb+GytGnsGAe2soi9T5mnA
MZhPLoVLFUVnpgpkqNvvg8e1REFNJ/IQfRhGCwbXZCAJgkrCF3s4xzdD8fwB
1yC+d9HlQ+neRV34PL1399POujmLT1AseCTXy70GucDcdQi4rkKAsCoPU6z/
IC94GKaRr3DYOT0W7Qp7UVZWUwZBIy+UBt1QXYtAuUVucV84JSAA3u+VgQHY
rnmkgmtgrKmtvXoiiPC4e/zId5H8q5J8cMTgRaN2DV7o+p59txHo9C3eSGd/
XZZJlPUhS3KRyAv/vamqJUk6PFCkx/IXVG9hm/cREuJy4SETIBgUyEzNDqZO
OIe8DYxQIlwZ7KqaESfIFTNRmYIrJojYULBFyV1Z/qTBGPGib8IgDsTqxXQV
SFF+fgv/xC1akwQOIn3oF9CP9uW/xgkSEyeQGXS+jtIA/sbS2AxEHfg3RAgo
oCqs4rlE8tXijvpEiILjhDmyr7z7A69fsuHJ/FnrgtYMK6O/UnyoaHoBGBQn
f+Cq+CCqjnK3uQ/v5YwJkVVfyAgsXTRDS3rMeAV5AM6Ikh63xWelWyWfQqbx
yaEufijXGVlxhNQQbGLOS58+DW91P1l76bFSUGuklbjD7EjUgwG6hWA0VMS6
NW2iHMXJCwGyajj2b62sJ8OqpxTIUAE3CJJOSLMVDQX/vSfkRExEIGfzTTwJ
GGyF6SqlxmFAW52Q304sMvly6a8ktRELMjmH/0aq++rb6AR5iLNMW6NYX/Pi
G5aG0QmnKqIldm2T9sqPYPsazhYN8UvOIQ02uFIpIaWDy8/UPhRMve+wXYCg
LZs/SEiENxsKwEoU6VRxpMmhA5CsGJ1zOK4W3bL8cDYsO/xa8f0WapZpntjG
qCblr2ieaEqbcVdzzm5Ba4foseu8tLK4T6szYvLfh3yNTiUoa3PO5+PSRbNm
fg0BAvaCr1/u55XxjkQaU8TxT/IMjQPI0Bb3E4xyx5tEr6e1zPSrqTSaW5Ur
v4iKNZ3kG1HUOhgPdrq16EfW+zSj+GvN6ETw55arU/5ho+rgTLmdCHr/KRDD
VsTONu+WNS3b6KBhPMt1/N39maYoOrCFzoVJjlcz6lBbPdJfLxEk2oifrkTC
ezjIkgucpwJccyNgTvSHcxIiae8Ik6ANdrnhjDc0IOagXBVQD8wPJ4SpjMki
6JPG8/7gY6eIkX7pre94MkzZwPR0bvfNRH2T18/VImQZYg51xlZyUbWwh6rO
cv5EvKj8SFzY70NcOIaa4+XutckZu4j1fBOXWRM51Oohz5REbU4fPBpDFqt/
Iq3Ny9Uo0nppzZdhs58w/E00BK6JSPPhgcIQhEMj8YUIN+BmmL/xoRcKPETT
YUSuEdIrWouL8bX5cC6agsBfuLm5/9HEiVYhUfy6GhQ4aje6/p8ZvWDlLxBL
cpLndu7GlgJ1CjrwnRJoEn7LhB/YWtfOdzO9f7afcM1Ne4e0VNAhtcURtPI2
8N9N0gDDST3oS8giMy32QOWJWPTLso2YTB6oZPDXEOCbB1CKj26sl0ItdSt6
LbN2spWdrw79R253hB2ERPO6l6KL4KTbqONP92OnIxJx9ecwBRnO2WrEM7r8
SYETgN8u1Xqfn9AKA6mfAzpAXsDH+egZvw6K2OF/e82ggm45RB5LZCOZYLJT
jEH+S2t0+3y9r/3zvkpcem01+t6EGrDt+U0CJhpX2COa98WG6nxTstxUHCm+
CdQhzIVvQGT2ZU5HUFWP17pMCGcKMQ6oThI3mLBqINL7mfl0Fb1GDZtjevlK
a1In7mmkbmEC2nOCRgjLh6pxNPnm1tS0QL6eU5VoNpy82dXuCEaUAfNEvaX8
t3NCS2XzXnN1sbqY6CMzZUuGoQ300L9OdBlWed/5D8ZYEdpPfyHgRUWHlbfQ
72s6/quE+IdN9yExWeIa2G/IYJfR8twRQOtjS4/jEl869Jg/NtKCME/0oAyy
2gOg242uaSD0Z/ts6Pl6YEZY1k5b83gBqEh/mVZjZ2RV7BAMnXrhG3QzJTXA
ThQeO2oEHzEvCLAmJ7q7uEf/f9jM42Nq8QgPGLil5UGGNnM5ryLQ8WD5c8gd
wUd3wj9pO8luSXFtyZvmrzu64178CNOmAxrgyLQBHjRhE8uxAZz5NN66z+sl
xbahfxfevzsOFNc/WMjrcY+hQm48VKzTlCEXbhU3YYblVzGmd0Q53jWKa6TI
yiQtWuE62Zvc/gr0EV472f4wddhFGV7QXeTni/NYp7LS66MdTd0OGuOe47dT
oxuhtPTtrsF5hI0/8DR22h6tSPk85MUVfrpb+rft83K9Mp2ODshVa/jsRCjT
Lmc6zOGqXlkLIqXcpcL4XfPUoBIsk5WlzdjWnKZEc7HbBeGlyyFl8OwgEuvF
/kbqSlui8TdlGoGkzS+Zx1Y7xaqt0AYiaHDForB7wsNsKGSMpBMzwPWXafKp
akkyxCxCuQqAlHVokjFoH3xfYoCPgild/uTV1iJHBKEG0ztLWLI0X+9EcxD0
BtHMGW6HJkZqL6NPLyXqDpOxbYdfyNtfkond2jGRUxP8l/BDJ0EAInpAnpnX
nro5DPcASZH3ISFfCGHK7zpjC4Q7jEsGpYD31hOOj93uajUH6DdIRjPVgOuB
BlmysdZZcLrXRqB5MerbCVc4glcWZxJ31zDwcy2uU1PEssFaaqOxf0bQFdtj
NMLDuY82ep5LgoLAGT8UQacXVULCznIbO9o3slHuaOOyWyCnRQqu9eEUDt4h
6+P5gMwa1wpEca5M+6bxdUO/sZ5gk+Sm21p29jDdN5tupucwO0Sj+YafxyMY
hwj0pT+eekLP6bc3c5JErynfJziG/xW07fD6OX3qkt/VE6kCpxGLdwHZ9JE/
NZlI4fWsyUP4Nr5/JOMAiTBJvu6EiKzNbqLUeaQP7XRZbcfGxVCmZXJ7IZPt
+4Cily+2mlzXqyKaOmsN1vdOnCo2aE3nnjS7K7lLxcy0XaSgAAn6uKWwvLtq
w3/QGjtJKE9UuYVM6U/W/Nxtt1tKhdgVELHM14V4HctZwUJLk8Ps+cqDCyqY
DR583gkIcJZV3Goen/ehChdS7204+KSA/1ixdq3leKY7lQf8ybJZnKPeAgXk
YFjJvnBaDBIbyCRjnLylnD3l/XENNHXgt/iBoKvCiXMXAizRviIM6XQ0obUC
KK869rUtF8KoADihKJ4OeIBvpgENoMORvZQYzIE9Wuw8gP/YIlhn1D4I3Ayt
QjaEAtIgnx0whUkxyK2DOOhcmufbZ2gUM2HVlCVmBiHGBRZfrpVs+ST9mIwJ
/BCeWoweYeWnEUyz99UyihX29lQFnV00p1Uz0LsLYhUDjwdRpfYW0w4iT53z
UlgPhQ+ZO6WGOL3ru1XR+rQ0US/SORsBHWPxi/Zew+z/9j+SqiaCxYUgyFC7
EBLZRPTrENMQVLKksshAZqTzt4qdgavKXHiGRVaJpZKnDrWC1dr7+xN46gAK
iH73yBknz+YtlcoDUY9BjjItSwfetxcCBgtZ6WChgNcFKKf0p3UN63GXzejn
pmN7Yi7cQe99dqSsy8tgFfIR3GvJ6x6StQ5GoLkaKR54JY8CBObWjx8PkyLS
gPFZyIC1f2ZXUHmjjt7eT6FSuJNEWxdG35OTuuTrIEv8VKV1O0h3csKOxaUd
9I0W3mPFI3JEyPD1PXJgTiiTmaZHinVJJjC1KB4i+9N2huUzGxfAhoYyFTJh
o2ddxmenDCWTyoVYG4qiCPlAUasdYXqvY4yzwZRsfju4gIr3Qf3mxBbe+7G9
QkehTSws2cm+bEcJfvvwUDiysi55BrnqAWJMJzha9ZZIm245LmfQiB35Wj2r
f2gJdU5RF4vIqkmSLAV46fx1RIUndTfxgp31pcy26bko0rhzuyukLi35KDyW
qqLwVZMGWpOnOmb0MvFdiaWcbMT7PuVUCNP+uEDVpHSWRHt8zNYGlkJX87io
KyZXh3EvIElwq5PDA73FsHn76c2UEDe3ycfK368ceA1N4jTTdtO2Q9Z4ZOkN
RlkjhsFK43MTjAM221oN6nTRpaVPkkmz+bvYumcxw493nZVMHEfJUDdKweki
H7Dl9NIM1kqKQuvJQBh+6RVyCjiY22jwDDkk9yuVmNL9aXUUgRogg9okdi6E
R43maBGCKBKAcxHCxS8FCBGRNNYJjBpzUxtRjhOd+VJHOq4QG1M/8qWsXBPw
qPZw9MvYMrMVCsQE/k59xJGnqLu9905vDdIa+lmGigWV9ndmA+UIJjsMnYOx
TCLnTMsmtZpXEMWu5Yj+9yQ951raDqkzhSnPTceXhqJbsQm4UB3KJ5kxMulb
5LwXkbC6ijc23/0SmgJ+MZO+Hluk7juUgn1+SBzCYoRC28GnWjaU713TD4/z
g9uj3qe3hZvGptZP0aOuHi+TEPCFEYadLXj/bsy2sTNGPH89VkciQFLNaujL
cKN8+RMq00u1vfm/Nsee5v5sHPpslbQt8dh5ACOgwWmVSbm8LnyvB2UooB2H
KiaH3OkUQ1emyvIyDyZHoXlqE6q8VlXS+2PR62c0kLhJ97E1oKRM2IBXP/7P
ke3GEVIChmmc8ieDIlifWfcFQDwrNDwX1p0Yf6fygL9G1l4J8oO6Pw29jmKW
aUf3SqtQNbmbS7H9C/XvAsJflExFw0XR0QGUBpGfgMU7h3EAZahQFMqESPXi
JDEznHJtEcHh9qXhZFbfSIKBdUuVuar9odXTZj7iP0PBiOlfk0rcCaYxNpPq
Qk9yziemD5q9BEre61E3yiF6beUx5sDPtIKpBFHO90SL3Vk54CrjMSebpcZN
JOiZcLw7ZUS2fywRQESOro3AgoU+mkbvbgQFkIIc/l49RofVme05U42pgRii
aTp1T6cCHxb5fa30vu/p71q4DcbxvU4x55PFyllMBJ8vH9iiRJvjvaDjE/rT
QtysKX5WQGjWDOiCJc2koHEQojz59xL0ZaP3oNmkmUjIiBziHS98h5hjS97W
eiCCXONlD3qhYxkpqEa0G3WCksO5Xh1YmtxYxYziD/mm9vRlx3pI+sxL6yRW
l1bN77VGGkBDmDpwDYKyvuDE1iJiSVvOatwzmLB7g1V2CVtzbvPsehJo3QUi
SQf0KsOkJDM2yeo+Nz7pbQjbAJFPzjra3rV29LGLa5FiFelsf/5dCYavY7FX
fCfaqf0Pi51JtOhbbEAmO6B+fZqoTt+G8ZXgGPZdL0PhCDXHQ0Q6OoLJVUu/
2ryIdrmNDrel54IYRTVFEyvLk8pRlgYWGO26IhVfKgV4lAmF7hXpCVjo1zKD
tDUjC+O9mmzjtAJDc0ar2LW3LXC1k37tC72Ijh3Pexz+CdBOICuel6SuxPaq
JPW+todUX4DO/kSDmEnm5jslWalaSx+sUbBcWQyEewvt2RpaUpyCfyFv9/09
aNNBLTrlp/boaEZQWEif40fLX8CAakR8nMRe5tOSWpEISRBRqhB013FX/VKt
I9Y/yo1JuQFLxk8XCNJkONAOhBZc4BYFljCr4lavL7NyacVYvWhI4AeK3Xrf
WjlMhi7f3pPoGfVXWq44t+xTnORvjRgXBVE+jwFnDUYQGIxHmXgciuy03ZP2
R/BrSvqmTSA8ndsTdKf3RVe3Ae2b+x4biabd+hGIHS1vEyd7VQ97dtV/cNK/
WwXonRVxO04QMW/uxNezalzQEpSJjfhyJ0aWI1ZWabgU+pHU8feEKzHAiNxV
+iAGiYukjfN0qeNTjMD5H2vQAb18d+AElVxfLIJtWVwh6wsQSpdzLASdddgE
ddt5BS9xUAZ8pCCM6edv6L6iZqgsbCQ9P+5CYr+kXJTc2l/71qySMfOF231O
M91ZNtO7w8s4SD5wqpk3Yepds2kBKxVzTuOd5EbDgS31GHMstCsEZKX6FyC2
3Ec12UyVCzhIJBpAFAIW03k6mEPJog0DDLIYvw9L/UOBoQpYlzk/O1brKlJz
463inQtyVqYPudLPX6D2AIRWNulw6thPemxlNgAhjRY3HWxl3LlVeCk+DkHD
SPpqcKAfhD4kbJWY3viTOdbC1R18GAnDSRvIeLk89RpPN64CFy+w3flpIKpm
ZO5FjzFlClqzMKWErGVhIWq/h8PB3tlgDuFeCL9w7QwMzrYb3/BtMK0XrdGT
prK7iMTCKxZ41F6IkMFdx0jlUjkIE4I8NisxtCvTACalFyZXFEb384kr9qfv
zFJq/90GJzeQpkb3cx2rmNW6IV7RZ6bJo1jZqU7w31aCMqRmiXbw2RDLSa8z
Zl9N+ru6BVXUKNFuocJBSYqpI77moqC+RsNRry04KO7HuMFUU6s+aHu3RFtY
4sloMgkjCSpbFeIZY0KK9/cMfjLf8Ycfcmmb3RG99eoGbsBQLlp+tKILeFrN
YZv84ToxU0ZGZL+pinY+/ct3CDskJBWGYdRQxtzszBevioI/UXoFZ+MNiUwe
BIBEn64qAv62xo3OQB5dx7eV1XQnJ4YKqB2nYgJypZxxkoI5pQW/iCMI0J/e
0jhwixMGcEWiPTOo9dkRBYLNZQttdueUiZ77LomXIf+pmOQaRmIAFZbFAHaU
2Goy3zkr7RJ3PrkBNqZirAQPHTJ+FRfe6blkrJMfESZEFsCUuxvKXaE8DAnb
YBKfkrYWZk4CvHa+NLpx/guh6bY01SJNaEzx259bpc2JOxSu6bMeYE6CBDTe
do916tidL6sl1hlWPJ7MIs/SSafSMoY1B+fnE9JS0QOsBwDPAUgP49ULJPab
1JrnmHPk4VJe4CO0UA6ZtdSTepTl902NdDkBsRplXwCkFJfftlo6CHhbXjfP
7+PeVI/l1XzH/ZrKItVC9AJDMxcxL6xGZCYKRYy7XIzyD9L32byScvaYWI5S
7zURjcFzIOhzVv2xzZrShRp4eQFqiaNY7Dps9+sYGyt2bG1vU1QCybG9eg+O
peH61dxJ1g8dfKSZG2e7OCh2TcZDZNulVi0wcW3g+N6oYzRUBg2VTrik8Hn/
wqMhemmuptCbO7gcsTWKsVP31w53+UOFDUiw0H9zcDuAyVJf4rmeykrQUvqe
c24PdMFeMzODJyjNRcuNkjajqVlhY1Sa13e/qFzEV/covKSrEG0p6icNQRBy
F0QUeX6OeH7+7jGEZej3iyvx+t/YQ6I9rOG4gaulHTYDgeq6FDEfY8K5CcSk
P4nKp+n3RIGDPyQO9QXeh+DqmkhX/EPRMYhIivAthtIl8x95cPIys+oAzzaW
oXZLyKN8X1LgGQMEqmpk6JerNk6XWNG0uBHerDwahKsOZ2/nK2gByXJ6tpZv
4XbOqNNM85xsqi9iSq3rei0smONCCU+CwMreBDLMRphI9sAn94tOKqUHpfmw
UL/fxNiFOVL6L+s5FhYCxbmQ4AzHlZ4UTObJ6Devo2/Amo39+4D4EuhRhfyu
9UcbiR6SFBP0/z7Ig/rBxHCIDIoir00h3XY+Pcc/2gK0x3XBOC5uFrdAZ3fb
y6QH52UKwbUtjAGiYL1zyJKw4DCKvlZQZm81VL6+1T+FJzrkfp2IQePfGI/k
CJtlXBvLItX63GuBHnm8CT4I/RdmHNz5VwjEHLQaqHER9rt5N5u8dkDbR7Np
UiCusYF5FAa0VKz9gkR/KTCyqPaPPROuD+dOQ2NY9xnR4m8HNDure8k0XL35
6fxpEz3mYZabJtm7PmH6dIQmfeM3vfqXnTG0bj7SjEiPlTjYvAS28R2yVM3B
GxLiQjbmjlmtjZZ/hNr1HVuVbS43/mvVHWHxGg2cMYjPaXap1FsAmEw3qgVa
wEVChKA04JuDVlZUHQYYLwlFMiFK026NMzSP5rqswnVbMKp9EE0J54v4LvHT
sv3iWwFQ1xGjyoZX78bXVWLTQV+pjzj6en3RxTtHXqg70bJAnA+JjHfqaZxw
pGbXGrjnECXqzlR6tjTeSWzPaoFtk9UH796oGePz+K+MESwv8A0sUiIN0d2u
L6g7TNRKWQMqYsLlmHf3pN/ISYPTs74Q/1D7cWjwLlRNSx7bTJrEr2Yta0Kp
ho1U7LBgFjqqJVoiFhjqAu1rty+RQkkQZe4JrVdd8ZARI0UxeTn/XjeHSTTn
VS4kFNBWgWlTKCvdCi13P51Og3tRKgMvN/1DXDd3S2HDf0DPgzoOohc+CFtA
wqx174Yy173VHowMmsjeVvXlcg0CUqwcBnmACd987zjVdlBSbPERKumuzd5J
l3F20rCGmWtsOTqOUdHbSd/jtLaA3YFR1YtC2CwEfl7EDkjZqtP3eHoLsZFZ
LKT3nt8VYUfyHY2TsgCWS/mQ0+rgRli5h6gA+jfxfN6wsKeCFtlibeIwL8QC
2ukahEWvRRxFCPZaQxwF8pFxDdfLkf9u1BmJSQEAJPprFA1/Ct3OwCZzHE8c
EzwaM71WuOu62nL2XxOkE3wSvY9eEhOpMpAIR3Gcr6wBbfTxddG+N1YU1NVD
0NUGwAhAEdr2DMIMy0n+qmVXg9LggVkvCu0Kz5O819rk8ruPJIqaH/HcaiGr
BZgaZDU6NIGaxiuwGnSVRtAJeE3cRSSusovZun9jRipYbSCbFRrTjU8L3awR
OdCz7eEKAQyAd/U0Wgh4RiwLXadmh1GTEjBXd1FRo9dEalYJFmRgn4hkutgS
qqz01SbYU2Sl/CffHq0nbYDqctvXfYLvg/cpWOPjUWsI7ujdqQwQOuyCBh+8
CPlMMkpxZcCfmShlP13GZ6lcq84AEzwQcE9vZDQqVbg43qocRH9d00k7Hp4a
h5AD6RGLg8CCMGYnFZ+l6Lha9j4SbQEvl9JGn2jermG0fQRngIGcHuzsWiVy
uwa4I5qEdfHaAi0ZO9zqwOSjv5pSKNZralEvZjzWVChToK1ksoYpp7tbLnKx
rdeBptkSYFWcCCI43as5psWDyho28eTIyWZO+gXXNei+ro52V7SxJxXM9pPt
1hYnJRiywcSVuQkBSH6jq5QSvbyccvz6DSkeDMXW++23l6eW83pkZ5eU5Tnc
5XKurWRK5x8oaixYuG4KBopO7jMCOZDuYLEzcNC5heACAvd3i2c1p2emvwM8
v4Sz/KGlqqjEP7qAaf92UfoqNHUURuEBOLpFWh7pqPH00HTUbBeOn/S9cclS
4Mqn1zKqEKw5B5f00SoYJ0xd4YMn3cTahyDh+uq1cRrbm+U23F7NQ+Llmmhq
u7+VcDsn4zC//pYe+3/oSVDQVSx4MhsbTMlM5r1DNSRlH2UF61zyohRir4cA
ufeRdGYOJ2mmOVzQGioy/EpL1OMg0oDVOQSKgPziw6F7BuDl8PoHgtLHRrLx
8fMA6FyfZ+hfiRkfp7ldwRtk3pQVUIvyvoMVTx6TJkwQKQQOLBvVyDRrPWJm
uLy03Zm2yp6Oqdd9ZJ1jVwqb2tVQ10SmeUe0WD9idwGO3mnQrDvStZBDvUAg
qhLuqUQXy6XxWqilCJZ7i2rHi72//o5SYbnvRoaEEVLKJVbS8ZOt3Q+TQJiq
sdnBrQolenomRWejtTVdzx2z5FwLeDTjUuaf6dBs8zTwTh7+PQfqamiR+hQW
HYYEePZXvWM/Ih7QQDWsMScNZvcuDr+F06zVCHhSpXWGDvu9PFV9REAHOc5V
gyg65owUJHOUpw4S2MeqD9pHv19yITAp2vBISd/FzctcFCVUM4HbZo4Si2gj
SyvO/x0T0B/LPgVl8s0/KAJ5NGCgZsuPNfs9X+a0d4ZLu74JDeeM1aKE2p02
7xBMZryi1hT8hmnZGZa20wkr4wYwaZ+LMVNTJ3jbtTqrKhSnG4H0o4749CK5
v8XRUg5Idkr9ko5Tz178oXM7j0vovi+D2Xd3NJqTa5t2Q45Ov+TqQuK8DDK4
TTabNU3j9931lvJBPk/Qd/0Ljzny9N8q7KBQMbzBMEgVCK82ODoLKg/vRHAV
hofiEnE2eAGSCNzevktc4utrPgPWslVQd2x90Wvdc5j3lylO86AxszQndtig
/K8l7YbIoNQaFBcS06lzbHUi6WjQKf5Fg5MM70BjCkipDeWRMEG4HTMcRX4L
XLbqYeeWdVLMJ89SDZFCtBw1NT15wnn41Nt4AuyZ4JA+o1kOLdJI2Gbry0Oo
auyt66O6K44yKPanusPomIYc2Um08vzIZ8zz91xvr5hFVQf0/Hkiiwu5ZUaP
y+S9ME+GEdbLJYguBYLdH8nWx/rxwelQCtZu8aqKsE6DfTR7HGnZQMtFtHTa
H0f6zivbr2Sbfgb/euPXUctMRoUnfA2MzKva61OJasphlPER/TQIn3apDbVj
pKNtt9Acg0LqBoZhLvUUIsANp5WJyClvE+qr0d8PAtzhDLQrJBlAap4lTsBI
T16HO0N9Al3WCtIFcZC2eQHQS95kb9GtnArI3AL7uOjYWlq64pHZsNs+fDvi
58qqR01ZDubdxb9zrnNXiv5Rsfo22C4DKb7U6qjK8tEXtCaYleJ/rtFIJACB
LeKNH7Xsa+EN4m5dCjGxifB9+LwYlS/Yz1+XZ2bxFoSlhKSrKuVoV4pwkDkF
2hryRc+4XDlXPdIY2on7d0glJHI6VEygnfj/+gmoxs8aRcotqmM9QS5gLKk2
1cdpKacmXLc7pp77+0o+vhlqJaqqCT9K2ctUKvHk7eMs8/CRXSEyzI0OAJlt
FdWWH5OcRkVRY6E7f7tT07O4AZsN89eJg4MbZch9GYFsXCuSqsWgeu7JUhjZ
DPxFbBJF4tt5a370Km3C5jT2RRaLiZkFV/E5iAhu18GGYHLhWbnaGHO5UYr8
ioEAmmjRD8x2Ij2fbuu7n9ZM/wPgEwCU+LnuNMoKWqTgaG9FSsVK3zzWGOpA
e+UvYyyzt14Xy7zz3oS9nPz3CxCfYY87ztMKA7OnFck4/wMiHVIDqn6RdxYz
L824/eU9gvK9+A1vXJPlf0JaN+kvBWXTRIoG98DUyBjgJtReVNO1gXYLJFdc
n8FrQRp0ulomnAOLkL4rwdm4B7AwmsnRxuAP4Fc5CMrby1K5+soLEDbwHmBg
l6IhVgrMtKhNrJBswFKBV18xICzxOzYI5AYiwjtHkktW4/5GCIBBnSTHxYwk
UwLIvWLw857Cy3TpHXoo1h8pBLb0UNkt/mI2udipYHCKrLv2l5IAdVj49W5d
0+g0cxLjxNFvliML65AB0nQam40Rur8e8djjnFhrOhcK9akVWz/qIcD1DEn0
U43pswhANJMpWXkVX1HcRQRF4P0IGCi4A9YU3kG38dsyAIsq0Ih0KwNEQCE9
UzNa+g8vfdKD0q/ad68EXVlRbLEbbevRHz8ysG4adw5w6cThPeqDkPJXhy2x
iuubwweIsp0QYJrvBj4zpr6c7MT0sIzYjhCYnf5rhFwEzOTrnApXP8QwuxzS
5jAQWENuCQ9NzFQV78TO2fsYk16D+y6U/Exsj0ojHy64bC7OQZjZ76g6Nzn3
aKYTKRj3Rp/nWUZlk+3Rvz90l0mpwOim6PPeYg/u31EDIpOXOCaKmM4Yjelf
5DSWN0Q7OedPG2ZiH5WpLj6HscdUyZqltqx4P2dQEmCHoOa5ZgKdkt53L0AL
Ae1IuP/mRlcfuWriHI6OcQacwREntZhl0JHVZN8SnYs1+19IpJxll9fDd9XJ
CsPbEN/YPjj31OQvLzcEUHzqz8R63+XAdonymB2hN+c+CGrVfua2U5oXIkAY
WRDV7rnXGAFjtqFqqGIeHQ/KEpiVbts63uE9muzxhpuOl1V678XP4srUQDrg
D9zfVf9bHyc3yyTPBtSnsM8UNbpY4ylJeAqQpq9qQjZjqVKjIIdFhnznY/2x
ViSZnOLSAZwdJkRz4XgckLcR+aCNIjfjxyVujIqdbI7Tww4GrXM6P+AUKgzf
RBbKLvbDNcLsDECnZxmpU18UhjgaIvaVupFGXoeOZhyZ0QNf907lYnP7Ucfo
gZMmbFJ1rX3bkn2/f4EGeqEH6AxTrGCSYJ7WsXp7fEbUJAb6y3U2gXnAjsCw
cM5Un45XvpII7IeuwMexZ346ieVr8RSjAp2NvtNtHHDhG0LqWOZ/GXkP7c3V
zA9Op6ZSfIwI2+t477oKP271WCrJ41SEt2IlQpdPRWpZzsTSe86gjK5Fsa6a
bUPDjNm6IO3/6psavMzuUAMkOQ1xfk8neGWeukYYYoRi3z0TgkYPfHqMS9Gq
7Q1FTOFPEdSi4ZLfaR6h5/EIzXtU7DQjzxNQbUFEFUvXcDY+Mh7JpFxo7vyf
PqkFC9FXUq0Ic40s8LHdOoVMqq0TRVe8A7cv0/5Sf3DknzP+5OmvSy2LRKrM
Sxz5m1RUOoZfOppBTOD/tPfPg2K4VZRmNwnk2ieWOzAGuu51kgRPrkG2ofwo
JqlJv7n0LkyZsHyRzadksuRXZv2HEYCz28uASWdj+hiFrxMwyfnnyhZvRBIu
iqFRIBnCxFmQ0b5pB4yV9EoEJ5MXZxwM8lR+kcCAZLitragKzwvZYbXz+WZ8
c09XIp9hodTSe/cFtdmCrxWTR4sdFlZgVEqxePfB2f1ja6V49lzzWUjgI7hE
lF0Pp+jNBPiqw5f5yUVH00kwtlMud54S3wVXlDN4CcnFMVUmzGjktW/8fpqx
lmur2Hg1DBgNM2mK4e4fONCk22mZ1X2PH/F5pvl1Jw0903KVCWN0N8KXHNP0
qB0kkxSNNBHQhvTORcrQJlfmbx5f5tV/3vusebH7Mn8CvU+JTQarVAmKT4KM
/WOXwGJm5jbXUO3FDtYlpW3/MSHnPydp/r+3J3x2saTzjHGCXIkVV/u6qxNs
zMgwfaErczixQ1MFxvyTOy8+7TtOZ558T3viA6zUGro8b/GCOA+2uYQqO8UH
WUfD5+TzITZ3EC22YC4xoXf2+qCE1oJqD0STacmYfc3pgNB1ntlrKo4ksZIl
LVjdo2PNcwHbYxHNKqsrWVyfIYPrPUBDYe1fIxtpS3ieo00nd5UGMuCz2tT4
zCfwkdkNHK2B5z3L/fl9wsjeTO0bvG3jsdixLlm7vYjQBtK1y6hsdIVg2wZh
jE6o1I4uZL5YnrzeJpSLqpR1ywA0jKUC6bzXYnRMmXLfGYfI6N7EEn0hiA7i
ytkf7DE6NaJ18GDprPqRmCRjdo+8nOjFqj/Ls+BX+TQkLC5JOapVK+1q1X1c
73XGMMwAtvTR9QYgvjCn0I46AJRN0NU1aThQwoIqHpadEpWv1Wnl6woCgXDt
C6dsB76IkByAYw5iacY5vYQPXQu7oYM5Wn93S4tluxtQ70pdo5ORwXjaoQ1x
/1sYjYqmBYrpdenxUJj82UHUmEsWYaiJfYMES0PCgvTN+p4WOVBVmKKoN0ib
Y/M1NyTD3asFjuz6AxOXRRTJKiwwzp3UOnGis6mIND+iamLcb0hgv4GRHkM/
6WQ7czh4lo1SptE8TngtK6hy3rSSewfyuwq9W5PJ/qpG+8NjDvCQJmvfzRPh
vXen6sZ88OCRByuyVaxhagIiBkgTi3MZPR+rSnyS5JztZjR6QJMT9qh25zRA
ExBjbCWRUI4tMvFYKoWyTp/1S5jNg9EQ3vbgUEE/Kp/c79oaROZA3Dg8b+Cp
mZmpC1cW9P1qF2FltX3Gw8TAGokkVz86jf2mDeVXjW2npwzPd7tbXtCTjrup
nIKSq07yvToJVIQWsAd4jdVggEt4+vtPRau3eFtJoAvsqTpBbPqalYe/pc+N
cM94N8Yy5zFRSGMaJZoGt8DjQbxPXi0/Bm27LHongvXXWDUGOcae6dh57sPT
tvm/xEVY4IkYUP/bgpVIr/clGGOwO3RXmX16ojLpz4uKg70MdeLOYw2tMUCj
p86UlLonN1ekPK4H8pcu+7iGYXuJxgiLAWR51MwX8MDY9UHwqzs+BICDujh2
AGKhiR7cdrBSZOFY/MMmIbWLFnTH0EfYeQ28F4X8lnf0QYdLdQQXLm76gdFy
zNxGmhLsg3FzYcyIkqZ9iVUeHwdvge8zZLUAVfUgHwgR4bLeAQtEy38okaPV
GUOtDL8q52E9V65aXG9uFUfU6hCOA/fKTlGhbI7U1Mzg3yEGCUagDcxFRoVY
fToSh9wAwHkrGYtIJWysXOL7tyRqK6+3Bs5unRZX6WDPDI9mhGRnbrxlRm71
TSk+ySsVPG66Y8PtrHZ/qpdNu95Z+QFV+gRsV3OZC1OMvOpPSwkMXdMP4wwI
d7Omg61FcTCoJw6Cy31Fwqk9Q/3Z7qKnHlXbcZwkwg9o8v+0xTfA4rfQYrrf
igmYJ1O5W4fSOBUaucHtU2vwOoOqZ/md06ZBA7AIborGfXVkA2TcAEu95JW3
CAdsc4Gv9OA0YmMhlwJreL6xn6fGfhMzw0HQYftH3R8gmRC7Glh5ajTUePGW
Rg9/TrgiT8Bq7KjD3eDTuy6U7cuRWchz34+GL67hPQvwKeprNIqWHisW+xxX
pUCdi+EIcqZdHehWbtLEYIzqelACUfyGkAmNg00Eyy68/F9qnZcD5Ny2aFfy
ks+D1hEMsp1zlNwcpnaM8OozlYGGz9aolFqfL8VPu8cqX5mX8uVbRyOoX0gh
svvJeDjxEm2lZt2KE0bXWsYTFHCac7GH3VuZHYQ9FmWBWR+d56tSjKyd8Fbj
qk6KV68VjRFIV13UuznSq6aQpc1yihb7d3iMCx+jUzIkRnRchPRxd5X3mYaV
Nz1WlGy8tnqMuiiUriEqFk0lIuO2D86Y0tpaDJPYswrXzp0fuhUOBiEyqp9L
l7b+FyEBUfhfqaRjcn4q6gvg5xbvLgifgW7rfQBJMoz/k5D6Yb6rPi8+mB+s
c3+bqVdsljAbyjqKqWb8sbcm8fPok2S261H4Sj2uqZx7RbZ54xr6xhmhtynZ
WK7iwqQeRMeod5xeCwu+iL/XVA6lg1BVthgSwJXLiGltn9mbVFkOSqewF/OV
Wh0g6PchxuMDJq2SGKjOeVNSLv/CJ5cF9rjbaJaFD304LKmnDBq/HDOw7LmH
vpCig1q9pq4LeJmu9P6NcJUJr3L9Af0RBGOq8EPKfUek37EJVRv2W5Hw05WV
3AsOLbXtVNwbY3EXiV9HJpcuWHL2BmtCHEYHnXr6fRZ3tAZWTOGR2AqnaOtv
nLoD1Fm1r9l2BiiHdbDyj7Saz8u8KsEyZEnbQmSSLgutv3aBSjjtLHMUgC2d
KLMjQD5e85AASfnkzHnaOpnFnp8v44X4Erqdxwa1il8s3DUlYp02uJzZZpjX
MKv4BUQxF5/8zoIUtdJs00gzWhMGf0+UXxTmotr5Nj/RQUy2hnsXwUlPcWd/
WCFs8VBy2WjEkfJ/iT7mPG+bhedwEApDzBp3uPu0GPs34C7ZbaLLRxSYbo5W
pjsp8lKARgwk0fTcvorMxnvKd7cldZz9xzvAYQx3XsROtCsWfG2cu97u8Qjf
cKCoOUSGJBhBdhRZJ7fodqLXounaOrUXThZ8R9E2zKKPjxLpM2S/D/7i9/k9
r1mG6YyoRaZDqs1UZ2FCxe50JPW+hL9HQyaxjfuWyLGa1JVucEMhSQ2Am/Bu
NIYmBCEw6c3NdPX+0GzZqJL7gnzJ2iEzKYTkNNZSOw/JWOTJgOT6cv3ta7GY
gyrHrcmEybZLz3FeDQLreAMyUa9JzOEgvFc81DO2VsLkgEasyyCiCooEHPF9
k+MaaK3htV73u67OrHxDtlAus7j8X0HsSzz5bWpdtcWMGvD6W/FIuGOft8ip
MCyZ+n/3WgbXbuzkbiyr7qmFwPIRkLc/3pHNv2wsljW6h0H0I5XvVMMCZ1Uv
GOsO7RvXJRLbFA3j0qXKwrPQiIh/uJPvqFcTSaDm7o1EH3fcCDXyxsqKLvMn
y3sXaj7iqzG8f8+PbVFhN7PH+PRosLaa54/JbrwwC4y1FIb+3oTjva52dFDW
+neD2zDGx3bTelBErxj038EAizmtKvD1sxAjXoPirR0n0KZ96vX9AyuODZys
jMiQOhgxOaUjqGXqhSvnJPihpLeYNX2MemkYWvFp5bfUNAkNcJUpI9GddEmF
NmXz7m+KSpoQF8CQjoR1E3XqfAJsVjjmyFjLDSyvfPgUxRvGKQI4wcGLw+rr
HJu2PICwrU80mCwdbRHuJ5/Pp+uhYFr5ez9PU0aEap9jkWQapR+mn1QBsyHO
dwCWfiSedXwqxm1px7ppUW3U/M/n14dfxQf8Vzh1Fz5xr7DJYUFPcl8a1YPZ
gz5ih/3IPGEbMb5Rbbj4ybpoJq2fevJ8HHIGHt8FIvIJGwjiP0bmCYR8xz7K
W4PgZwn0XN0JL1r4n9uU584iMMzvvvEiaOgC4F9i6Q2pQ+Z9xoOOC/WzyrEU
WhopjuIatvA6ruUhHqf1KWpHE9GqKBco0m8LLFPDNVmRu5mI6wD26YuQ7bp/
uxRTh+XN6skm5AK5nByKHVu/9MBRgsyHDH8642FMKZk2ln7VbMVibvTvA2xM
pGiBtfeMvrV4x8sddbmlM/bb+IU2l6nkC2pJV/xtOqwSyorLFUyS13u2WZXU
4g1pJJ/GPTiCKuXVLkgjyWvIflT7/UBQRXS8EJ4Kt2RYZVCctqviYCorxxGV
MCTvTbdtOsqAx6X7oPb/heo9x0xW+6is/yabb5t3ge23LXZvOghC5xWAye4v
7/mwQfvwPnHeltwqyYu/vG0rowaicU92x1Do636jsWCuAT/ZqiHmNrqIZv13
WYgXbWXAqxM5EgZFiEcem0fAx75MeYn0JZBo1HL63QqemYF8cKblbyqjzKWI
2IK3qIWOkiczOe08IFTfB0VggNhCkoI/p3c6Z4+YS1WX44SekPfEQU+NgX4T
CohbmIPHAwrm7y1EtuxIpxDZGw6JjV/vgf5vG4+AKSQCrD9AqqKTj8Hj4DF9
J86bkKGmMUAT8z0DJxAlr4RfFkPSj2Nuoi2aserOKYtYEE9OIlHMD+coJORz
UwVRxNvxp318fMF9LUuyweqRoC3ZC3CVJdCdJO2w6uoA6uLI4xm2j16KApyN
1WNv2FijrLKBe8yIgsDGL6FXon7vWrgdlE5RICEOGtjozXL85xN5LMgd/Bf7
xiYo5suGMYmTb3eaPrdkVNX4nwNyRtoMgpQZUmfVJz0gE5nLt38vXH4qSOmH
fb0MyJW3ebXBS+XmKP3UMbG3DruoTNy55OxAfLPyBzPodH7Z6GofvC264HDe
aj8Do/3jO9KnPJ/FMr7JluZnTacRh60wpjfHbkdOAfyB7Gl+Pr1CS5NDhlWp
yjQUGSw0OjkoTLimlNCzGtrQ26oYt4btBzQkxPsl50u9XWTcy6BCGgypFzif
JKhClUokOhkgrI764+x3pdbAttaKn/du3xZIHlGELOx0Cl2IeOOYEm9jno9f
2RFnTvxRsnbHr857IoF6lh9eVfrQnuIpgRfD3NWjtQNlIaFrpU9NXIrW9iAO
Z5lPk4WPiJX36Dzk1AEalfTkZPdLNbaFoSP3grygctcc8CeNnI7DSumdtUt0
Ttzl2U7DEprsF76cYU0mPFs/G5GuKmI2Tr7XTq4B2Uzc04qeHnw9+U0yta5d
n+gjTfVBWtZ8kESZBHGWsc5kpQt9HtSgXv0/EfTdGLmkt2uiLx+SK410EV4D
f+M9y5yTwU298Qq2fHHInSi2MAeIewhrBrYmxSa79MD/oUWIQXCNEjgdX4aI
QWH07G6kCQ8eQyXCtzeGKce7eDxkpSLqdNqDribn0tOraHDOIInSBbthHjMg
UYqcRAEfvoTU0Bswt+CzY9kcy2S+BUoEP1ib4RdwvsBxhLtJpRbb3Ugzxw2Q
ZWHjsVyBDcEyh0H4Jmy5KDcq6s8IenDaUylqc2ceW1KV8wIIj0zXVGrGlhUQ
E7KnmMKaLqePHmWFlv6tZcvu75jB3e+2hbIy0pGxnu08WA64zhkYNxqkpsGu
+WKX5eIbq063mVYnFHTLMLbJ3pzOSNO6CSlAiA/PzDlQLSR+vSnsMN/rL9Ma
UxK6wnpSXDq44dkkI3VxE6y1lUZDn3nbohelUR97WAPPjP5++SsWppAn3y8U
mBDiaXTEtLp9OitPlH8ZvamXHc2xJNVguiy6edIsxcoBGqwEzTHo760Qyeka
nKknNnoQPOCduSSWDBT0aB4da8wNRWN6ZHL/reXAg4+4XouWjLL6b0nbMB1m
iAbEs5VzVTGUI+rm40EH+1rvkhLlF3BekjzM1m/ZacTNAEP7kTHvciDuDEZt
kpAb4c3qvDbg3ImSZGjFujOOe8D9sXOl7y1KDd03Ta1OoTIURDfVhmoqQFMb
1CyCKlRL143oYsZ438hNMXnyIflozIWddYzs2GwiO/2OMKWGzxXN+/F+/xHz
JU1U5DOu3EsDFbz7DXRY9L+hhgjYBHk0Ij2+m3huj1oMTeV74Ezr+VddVQdg
W7ShZllpCF2055DvG0mLBnMC5UzgMIMf6dk8bH1l7fIdX4nj1f8p+dtiERjJ
oJAxumjtMuZ127+maUC2LpUPyzgO50jQjzPHHsw1/7o/2+gIbfkJ8p1b+pXZ
QfWI+cYlkorByQ0TRovpuq2EWLvf65w7yYUG6AoL5ADTGclPFuIrmBeotTSU
wh28Zyw5c7xhaIhV2vyaifXs/tmxwMRu0NXwOsnymWqFeYRu2sPl7zf1ig3z
l1Kr1CsIVvvgSudi1DDhl8Ed1t92k4ADIcAUVVsaQWQTeWH9cH1oix/dcxbf
NQJfqsFSz+HBCmZIqrDL6c17tB3OWwXLIgXqFhSmpqB4f6JtB4oUqV3qEUHQ
gF/L0raSiYcrp1TFA5pw715g1/HNwZyis8CsrpcOavcPkpplClf0uNupPlDv
UDs0nBqGaJ3cVxmKr0mdI329ftSWXhntUky6R1kyD8LAoyDUXMlEKfPBCXJ+
IRcum1NU25vKbEtaTtXCK4wgaDTtsHcsiKXxuFY1VMTVZWkgBcf7vP0KwXHS
rb8wpWLgSnrR5FdcjsbtMN15nqf0lEwx1tVN271/rRLwnpyro4J38LDtE2h4
Bdnhxn0i+mi1+3VAKMCenH+kZzzufhGSQnRALQkwKjdynmR/+heQbq23D6m3
cH03SFXmZv0Imo5uER9edASO25ifGBdYzSBICeRljUaVDm9d3uXUcuJCZeVr
1OqTrkJjTJoWiSQlavriAsqPe47TIT371QcjJ65/qokSWtMBzGIFvaU+5XIZ
ex1bhtqDKhRPvXyT5F9lKrMaz6EFcgacb2LlqEo2RydF/j6XpDh4MX9Q25Cf
Fw0t2Tc2+WPPpBoHCffd8wJ89H+fmYXbgkOPJ5J9n0zt+RkH251tdmLZR/ia
borayMikhoVac1xJRDdG+alN0ZXjgRncQW+DOewYgY9ozXkfTWDtXUrKUWsF
534RMm/Jv2Q8Tf2w6MPtrgrxJsmcdzh62InEpPU+EqDF4wsCOzXa/mYQZZhi
L+o7EUEnmIZ/4p2aSHGFdSf8EYjSg7HgZe27azKeqTjybhoqAhLKsFCnwImZ
luWZU3HwofH/vKk2YmOD/gIeAfAD8leyngXlHeMZBvWDcJwOtt8/v1foV+Jd
3EFhTSW0be9sQgQEjMj7hLLYmV2ADS8hoZuWZSmKz0/+TyHDSSqJ+iRoKZq0
LIYMXv5MhssTUOUiD1xa9d/zWdM03OJshVN0Dn85MCQjz7iF8XXSyTpo1Zz9
psmF/8lkN9Wv95ERJRB+s7W//w9DGVKYGJ0q4B7b//Chzc/+ld64XWeoo5+0
FAAjCZK/KNO/j7zUJupDT8cUm39Gb1qNzL/4XFZ4xFw/dAFqt3FGpW+/LbL4
L2j4o8WHwH8lbSs33HGziz+9+xnHoBJUY14R2pDQbfH6SVkSbYkAn90P3pzl
V6GmDk+ptj8bBebbl/94QoxSXngsze8wAhwO3gXqfkhL93/+KwaLTf9CL2xE
+10mKJhayxcghwdSB4/PNxD/laUuIW4/qSrzk+4jbXjSfOsGeuPCSpD7IzIr
SYRYoE/CliHWOaJvCxBm4oWttwr1I357imhfoGtfye2VOSWOS+ysE7uNIhHA
2VMjNKIvH0mi1FHy/qtdsiXuERuYIEfenSDPZrAxLVwXEbWB3gQknXxCfdI/
HprFrOO2ZgUGg0weh2P9pZnwJBH+ZYyABHTLx5nyq0GEkaRZlFjBbQ8Q3vyt
WF3kyvXzpMq5DEcCziBszNaoHhTVAl4y6g13JKunuxt8GrUoB1YgmBeTukmW
BBFuFWKsQQRgHJLgcDL7C69o4S7MMeSqKeP2VWt5Z6su68aV5Hg/4GigDGgc
n4kabJGoqWmW81WE5g4Pu1X3a2+IWTqexDE7uGbmaf6WmCBMjsbNrJn7JbiY
FmLSAboSQOUhR+JZh9Wv81zX4MLLEi9mxQQRycJV7ySrKJkJo15dpUR/WNJr
d/wi2bRO1O7GHp1bVzyZU4Cs4PQxmwyGfaZKo1sebxSdjI+AwA4bkDxaoJpQ
3fbv0Xfiy9m9dXXKP4W6/ZaTMvIg6RfWejYfF0TFC7yj4r3aXRI/M6Muu6CN
RkHyeSC9yWQDGrvo2puRhVPDo3aLhWrIwptaWSYxqmI8aIPza+ElmrSMaof0
/FvJOtjEJFo0Cs1Mwzh77hKttbL9kxIk/RXIDNOx0p7rQPoNqzlJ+3NZwuWg
vetW7J1Bb7eYi7jpo0dUPSGNm1d0C1+D8n6IHEyiENzBfRU9Ntg1iJS73wL+
Gnz2b2h3gVQfX5zYIAOQKp2PxwbCOpJn0nHCFuAeCP7gyPIIsADa6UdgSGi3
AWFkuYGt+/Udx+uvplTAnxvBmGfKIhGLmJDxQjxuUFUFp3C8W100gt61WwWs
mMP/kQO//Hk+VxQQEYL7N5TylU2LSPyp6eA/tR65hkx8tuWgES7isuyLH8/b
A/YZEO47kbS4pICmRCwpDAGMfu5313j+uFdNPTZW7ccfDX3Vfey0qowchft/
N9dLjg8uQ7wv4rnRvqF+Wg5If4zEzfVP6ipyWMr5/lIxFvzf2XmAMForlrHC
B5/PwT+7L/VLFtvYQLHc2cB6VmUDGNHefvaxEBUNp1w/gjDxaoWgEgwdvNTB
+6FsPr+cUVPeP4cNwtVFlYzybfYXtl6pzoCvFxCLOeQFSQR6Lg8YWxkJC6x4
KolaT3y1FSbdYRIle+C1i+fj1cV8hAt0owh7AKKpfY1+HLOTrY70g7Wjac3p
r/PLICYamLbZBJrGkesOy70O4NVEzGbw3ijht/yXKktTdLTKVeGBwAu1eEQw
d+gSWctliTXWICg8FeuigNA9ChSW4lvSB1wTzAdc/RE1m4v7j1mabr2Q15YF
aMgdGsjnR/rfbu/SXi90b0DLfdAT9UxaJsErWGyOsU+bI/BsXFzq8qHTc5qe
YjiyKta0bGXlI63oURh0BAw+lu883dWGVQhj0ZPjgt4MlyDtOWSgOdzbj2jk
RFPDDAa7oe9LhQ1q/Ra4l09e+Aqp7c9B8K1kLtcusBnt3Yul+nMnQ6pALami
VI1KiOOY6vcrkenCtiOKxh5nPzIxzyY1qutWBXbSr8+cJ2fjnm204j7plFR2
KMDvUrc01OSxfUjEQaLrq1/ujGDR/LFKYscgRnqWzTRJy2nC+oAdgzSAIJV3
ak/NG+gFV5mVdoQ0zJ78qlW1eztxrlDKMyK3n5jaetFWD6w2KNzADyFNtK/D
u1BkmoVmW7Vsc/uc1YPZ/f+zU60ePWXwsljr/aXVo0wVIC8X+UZqxEmSWQ/o
ENGxs0mgvebRwyTyGMSI2x4TOn7voEQrKF3ltf4yPnjc37khPRtz3sMQ4tSS
1/UhfoONgKyX+yWxNYGF0fDYfdYcbByoaiALwyL5BH4BozIa31nyhMdA3VRR
pbGj0idgBMGYkMVUTzagE4jgj0TjeAEg4D5zt96cZ5FVHYJNtEmYgQAXtyQO
jHq2jQ8ZOcAQvQ20FvssPi+JeNoaEzUCsL4PWCDrfjvKu0iCLBwDkBKwmNd9
ZijABYMci4P3m51xKeBGUTBPvm+5Bj2sp8baxeBwylS3kQh4Ygy5bGOwnz7h
LVq/6JNHxvB08r5kjku8e38iq4fRGr4dZvoF8BmNwcJK4WRMDZ8e68paEj9u
iJ2Qo/vX4YFcUIk6Mqd6nJNfC/klBpUeXT35k4oicH6DTDwJ0cE7DnA37peW
cpv9lvdva5SCZsqHZ03/NdRRvNFrarZ0kK+FSXP0hU/n6dp5pQDBJ38Obvbz
gBfefTonMDLcdBB704dZWUHsXWKlYnZ7lxxcZ2YOeC5c44xHp7EVoH3TQmC3
uwip0IJ6EX0w5F268ugG00V5uA4v/Qh2sC1ghY+R0q+lySQGqucbWQU8b8Ds
UNszGKt7fM3198aQJ72NsYVRynXIcwDGaG7D/wWNTl6xm9pNN8PXLtvAoyIs
Ak+w0HcQLstHeKjtTgK+R0yzHq4yY+RpQCKEfWiur7lBMxsPah7n9N7RYYHv
6X17BfrPsNsPRcP/qAL67ujAU30Vk95oCkqdb+GlWe3czfy2WW/1IMh6T8AB
xPNA16frdH2xjZyPFAkEd7DvYstEAFSZVGEsWlNOKGfWPIlV/y3CsEl9c4OK
mQ8slyQitoopLMhY3uamiLqrE0hvNeZhnZ17Mbzr1D+nyTtKDqT8itYjeWjv
j4/cMKsiaYD4j8HAJNgwYvX4q+JWFaY4BFedVGN6tL+RMQBZn00GrJDvWJyT
1wrxQpyf7PXD2S387QkcPk9lF6Q1MhY4DzIgDQVVS2dNn9qZGxCm4M3Q2b9P
jz8E3J712iTTl1OG7siwtIew3dcWptwQlt0/9dvuGoq0m8YZ3/H9TAUNlnmO
bWgElTUJ5XekFTVpIwG0+fhrzCpYQ7yBlj6ZykZ+fDvI1K8MmMHWkFEb+T5d
gNlFP9UbS6gc0PX2jr1lu/TmdfxQG2iGeV6Ed2tZFqjK3gDltBHlPPmtIH8t
ZgTNFiVC/PFEKXsjPGGizrH0Ak553KWQ5Lm3P+Mn9RDBDcPBx8GEkcRybcKE
arNCYsRbfTJWnJIOzVNUzX0T1/1V832ftW0Bqw1SUdO/2QA6oHhG6VakZLNm
/Cz1t4LrWtmPANv61mkibCB67L8tyxYN7xZCs22hda4KK8hH7PMv3vWniH+j
BHUgtq6LQt0ld8VWuXdj4fRLtJS8XmoyY+VrVphp5qcT/aQZ8hu1/yLF4NhL
wMTKd6BShbMcSLcDQxgrK7QXNKJNCKDXrknkvK+yxB5Fa9YBfYr5WhTXWKl2
60+kudbLFLWjnHOFNQynyOc+1p+fxgpMepSezYQRW5BSbAtMnwKkp5A/Fi3o
ZyiqJctUGTVaVo2eULXVkuVFkKww8hw7kQCjuj3ToZbvCxpg52Aa+asqSSZE
RfJzEsRxEGTyoSR4Nr3GqZFycVW/oAYF8/aWsCGXKD9UZPNRapWFVQW7ka29
tA6F2MJ+TZNUu3U5x/sClSFzKE7HJKuMUJEuGc9kxYc7TyTNDi8KhunSjXCH
Lu2mHJQulGPlq6DQLTSji4xWLF1AekMnV2YoPHx+ctUEWPyiqZl19VT9kKzT
uKhABROAcyF0BZVEsDsRgbRKBlL22c9sTxXAj4AZafTKRV7qMwCpy/MYueg1
gLe0WaOLoIYLB4IMyWKUViNbk6HTMfWAMT1yUbD+3wNka/PNuULvyDU6TIaU
AmwNpKX1Osad/w3sWLLUmtv1U/9G8T9B/R3RlWoqCRgihl0lfUqpbzfZnel4
aimbpI1o0Rj/xu8pVOueX4ZTJz9jGIHfKrMcTCW1Ga7xlb6I2aNLzAqKypG8
o0O5VQ2j1sNwp4jXWeXwx86uG8BEG5ydUyrDaJV3an6eUs/9K1hFWZW3wT6c
XGQzF3B8TStE19M1xdV+0nIQKWB9h9gvpa1N0rDivi6G1x6GNl5LWakPTUdp
C1soipmzobkUfo2mhhC8XEY2Ane2yG8b4Kpln+HPzFD/KUNkx620cYhro50P
UWU1iS9xUL2VkSrCxIqDdnD+yOluJFxSu30xgWonmcAiYFrWdp9a6/vWVJpY
FAnS0nHVK65C8v8/IeYZVVRTgQRn0R3hHhgwkYxjk/phEKPBJrfmrO/C15f9
gAqhJMd33zIrKC4P4s/XA+JHP+5ypgq9gn0BrY/D+GN7n9uWIrWtpB+Mxp23
DLUo6K42fIdY1pX68UTJ9tf0L65pH1Wf61QnOzraoneE4GnocMwuYUaptfQb
O9o3wGvCArHTNSislEND0nen2EbjiHkrnxmR7JYGESBc5MPpqqf1LJbYcToB
Zz2TvkNlVtbmdJ18w0+AyWwTzE904ElthjTw6k8vzIqYi7AYePfbgSLYpmuI
MMwYUWISavWYytpoq+m25UNPlv6nAiTbQvqBBMCFEevJlDvoeZWv4axtVGFk
9TMeTMjB6HQV2KX2hntbUNxQqk7RsRGibcODrn8hUMp/MafJav1NhYMdoZBg
llLDB9tSupbWM/MEy4OxNszAwTTrGwBXs/VyJgM+X0r472EFOM0YjRBa5MLV
jvuq6tdyTI7oMd1ANWypZD0BsMt6n3GmJhUo2/tJuxrC+3c68zhI5oqJRT71
czU40uKXAMtAymjV80U5lz/cz/90N6OJIw5dqmRTYhEWPRAkXOuB9Z0Gv33y
zTuenZuhRb4A0TumD4UKK/wYrH+RcnFAI7FBP87QkgfnIGZfNrQaeXaXzsMX
fJck5ipa7UhqNOq3nBbBg3k/DAjAe6Og8dcExZPPGgQ8Hgi/IPRiPTxq0DM3
6kkzy5iLFCUZugBDI/xw21i/ZrSP2Al+wJ7UymLOsY4UEDzhYGZmizMNeNFC
URJetwn1AXNnfJV5l+BPN6+/MBwLST47dYT1qYLc/UNmdC/+eL6c7gscj9vz
5aKYfRuh7BOg7k1LDZ2dyQK89YFPZpXMvRiF5bTEmW9LDJmqZnOoSy7KOyyW
1GAQFowS47mRttiKs3quVfT+w48RMTxs99fmNh8BPVNjAsoW6jpJzcDdwdQd
58sL0Iu544cchHJiqhJp0cOVi4f+JrLdDPa1QVISKLNmBfSKgHR0plLKPEHo
XXzjOVKI1Pj1+SzvQyCyYJQYEsnrZt4ckRzFe2N491HPbBV/zOfzsuKdVZMQ
GxjNKqNYBVAD2qYckX1jAta6IB+1vbYNUi1+YErm9dRTChKgW8sXJbHFzkHL
qY7yHarJ7XDwBPE73CJaX+GDX6HOa0rXZ25bJ3YyZwj4AKgBN33Iqxy+5owH
GLWvWoCCU9R0l0ObINXtD6xhG3cjpPBlzNEYhE9bgGu0AR+yatOG48ULPZhU
BJsZrHZGiY4/a/t2b4YoO8cwzZ+y3stFzYfV4EMeiebhBUCMfROvy/5OhoVe
N+TjkiVKouiRuNKOOz2BrCIAGno94Csd0+aREDNoWi1Fkl1FG+iKf7o9toA0
iwgDgggnsy+tzxK9BiLSyGwkCmU4JmTXYO1YgrkZVVf0cFlC7C5D7F/Rq7aq
NGg47yOaMSPhH1IsGx1xw+UpOovfhcrJnD5VH3t9s5rWp3CdOS+fl5xZiXnS
U7lT2zbQj3JXTopu+VINmAJDWxotesjtTkLTC0VzWZ/2xSTWp1DSDkHz7ZCG
sf+rgFOvXQx1fJIjnpWmVOLaKiyZ2A964t6HMLT1BrekYKgcUPUvCRdF8UIm
UnNo7YtGw4aa45rVNEYAk9O+WUx4W23wEcBgNXfAixSXuWMVbcsPqrepg9tF
HDL0adTm7tpidkulppy5YpLzCSOgJH3f17IoZ+2RuMJUHzDuBFzho5AKo+BP
VUTPTvHR76IHxl8+/Lwkn/CnAKByx011vIVk4lpeYVwnN3lbm5jEots72kC5
mch6qmuOZ9imD8vB3zjp6CGhpUKDIwNNm6xZ54ot3zVF3onPpuXay4n9heVu
S6t3sQslWXwm2haVDbNH80uPEKm2H7W9omBy4L6UMzoAAMMfXmntVPZPF26a
a936xCl/C8+vplmSEcDsApkz1CjLIx6qE61wz6Qk5nkbJy84LPPTyT7pKa8i
3lhzDaaPpHosEv2lJP4ubhSgeq0i4fBF6OLPkrgbu81gyj10w1/t7hQhOgi9
Zsn3i3DF9YmYkILATlYj0+szDmtUWNe7EhDxwwkzA4luVlWdCz0gxDKlm5UK
hSC8c3vT9hPR5bRJFXlo0ZB1TrhYblpdRD8ECXDY2g79gqYRa2W1Og+SwoIg
TZu9t3TOvyGOj5Oc+XLkHowdhS/ohSOft8fpj0gbqmUmHnYIdKR4TFXSM07h
LxdWgAZhPhkKc+BEBJxslCCb6RXOy3ImbIXJQheJsO3ylT4s3nKKMelbBKt2
ssiUmGfIDtsduU8GXNGQN6vK/MXgAY/6hVwcvI3OH4UAJNFe+MocD5o3JW9o
hxoEt345M45MbrhNMugAMoxxEqgZLs4s4Dg1BGiHf+slNMHfpJvWsbgic8Og
Gl8OdYNhCZZSQzVPNqSzDiN+BFuMeKFuBOlc1nmGTkm9YMbG3djhql487zgD
qs2VCimoujjhrxUJhxjv+JE65zLq5IDxyV2+ys+AaU0gX8kIpqvvzBO+3Xpf
mIOc3S2hhI4GUACMi1hD8eLR5YZCuTBIQtTViGJINvZV+t/5SeL/Els526Uw
9WJnC/u6EjJ4xVWfhDRkGGgrcYuSbvVqHEx1j3rj59J2OkaHCULvMcxG2LwW
j1rP2Qy4LkOCb4UiNe9dGmBle/rLeQiwLjLyICKaPQUo4c9cX4sLiofOvlWa
2WzVHDiV9uUyIbG06W5BApBu2XLwysE9h+ekRZIB5xeq97W8cDmBWpCA3jNB
nKyQYMtMJqGglrCgbBi6/2K1e2RXh2ORRCdF5gVXAPUv82kRqnOsRiiZWbQk
HrLNRBB7yJ2QW2zCJX0Y2NO3+0cs9GCoX8t91UScHq8oMDUU2H6hu0INVMIL
n8CBzBGr8KdiYfDHE78FFZvLuMsl7EQI+Ci83OAVtFR6TfyhyD8q351k3BCx
tKMeNvsaA5VffIijId0WdhrkXU+AVNpwhXjIkFP6thco7ca/IsjXsdUgtsJO
301DTwqBryj59jjyVMXYAa5yLiIdA5Uxdz4+BUVy76EgKESUeJtGF5ETVmwk
r0NHcNBFdVhF5ToKoy9UFNrgDDwatUzJD689OWfIDkIN7h0g/wwBHhRrgfJS
2L/1yU5pZj4zl8il6kBtgkihGCJvWVPSaoXU6IKd8FQEu1Z4j4usgNMoTLTr
/Ulky9Ct0KdBHfAiL00RXzSKi0Vp6P66DYROUCADz+u33vXdP7iTf8GjHD4b
GvXNKc/sDKZFTJsGhpqQAynDgtbsimmhIQFLAH+SfHj1LpjiMi8GfgtkEVg+
0QNL5miGC6WEb1A5MZEXmcJczga57oFdC1Gvjb0PuaUJb3OWfvVH767Vn/Y9
Omy0VIVhTXQFrndKf4EKJI1RR+gFufSD1TRE5M/PEXk5Bpk0vcmLf1CDFREP
zOSU764d0pvL77ZRM77sug/Ft3YhB2WBCkDy4RElCz/zA+WGWSWXusUNDTAr
NbQt5Hd7rtsgcxCzhYqfkwLesNw5yt13kQPAmPIZddxseEz8hCnNZJbse1W1
RBzsdC1oP2iBCIXyRXFEKDVZuqpFZl0EMW0niBZXflGxQS0204+UWaMe9mBQ
OPwJFVfcNW77opKo+vNI+Tco3A8PDsayOFJXyzsh/eWhvJYytzzulaRMupFd
28Dm/2Fw/HEm6BcbW6zZ2lZL7i+pRvoBLWR2r2jv3HwEiaWccYB4hn/CR1Rc
+8n0wY7JuaxB19ShzBIebIPPXhRKWfPjQiPStVRjQjB/vSWFdi5lMsASCvpN
DMCOTSw1UqwiSIFDQ5+8irMgDnYSEVC/gkHaln4S99fW+EcvpulyQ7Zqw6F4
2rof2OsboNUuPmkDOpxGNp0WpKt5PRhglhWyXBI0zG/itYSfX/MX5nEXHC2p
P5ZF4gm1wHJryH1WnD0RYWigW96IXh2Old1zYK+CGpcjUFddKCCSScEbdn0J
JWa5nj9qIJ37Sdu+PGjTgEw+M1hpikJFQ92aL7oalwUSjIJRbB7OODhQ6w5k
twyEKzmH6G0SQ/3ZF0b0rWKdSyMFqo0XeM/Y9ueifl+X7hZmXrepp8gPgooi
VBRoIvCGMgV/lyUapVxAVGLR9DeOrMpxdOLFprN9KWKq03Gf9+QK5Uw3kK3d
q/CjGRB7qLJTWeT3N22oGWBAmqvNPz0mpMIgvpMtyCLMo/3Qz7QLJvLkb5G5
Vl937SfzW89i5NrlGDBCo6kFVwWoeyJgmswMi9yZJrJXUPifL+jZYgC4cqFm
mc+/3Zo85WGOFAlxsnuV3dL1nAQKodZ2+3h+ghsH8qsYzw//iR6bZaDYK72k
kBfy2Kai1QWfBjdLrqiJEz14eGW7DrzKDt2SMtilGACEEVZcsa7B+a3j6Aga
coZ2igfzLEKXAHNqIHg6isZr+vc7ZAjJX9kJB8R/bDOQuMMyOO4bPIkvinGD
pk6x+MhPWa78yJoN7F6z95+1QP+fHKCkihX5Nn7zvo1WWnp4HBcohiWfSYlV
I3A05PlbgY8zY3j+wR3o4aFRxTwnq4DhCZ0WOUwSMm2cYBq4HhHFkAm0SycG
FZidnkiv4zRvZG3NTqm5uTFFOi2Ew2E+MDYIGkxd9qvKm4AsefmtPg4wrXxc
hngWX2yoIp+crmw8Nv+Ps6dfVC6VmULgSxIgb8y6ryHKbN2Fne1L418hvtkS
ZUrLovWIWWb51ncO195Ay3E9UL70txoIZ9I7KvgW3br0+5mvENHDc7Wf3lJg
3bLeveshcPFOS1nDCRDFo2v2y3Z8PlKECFTil4X1KSEPZAGQ+0l++b3560jf
jXFQfl1q/f8mAIsfKwwlETBEqn2fTCHpq9TlRJMUfTGZcjsMPsv8yYgeuQxf
jf9XKY8E8XSLC+nip/qCQY/NA4IeLUkVDY5FNNcnjP6xMNfVlVwvmQ6iVRgI
serI4/9X2eI6scGm5Mg1ZZpRn21VCVR8zgFgfVGSainTcXCX9Y6eF4VhWaYY
Ip+FDCs7x04q0EyCwaNyJDFoe6gyhss7JYWMTmLQRa9NHtdhrSwidnzSIQV7
cLWPwByHKcRoYA35bOCupmTYbQAfs10T67OCJOvn510oO/64ndpngrbY0xJu
hkcJJ23omoYYruPiu5nK2JRASZqh7T6JDBIJIEIvZaLcHWTVMPNgliSRNwF9
uGEctFSzkWEEIEXDhOgX2oX5q9nM9FR5AbVIu0aSBc0NPNNvxzfV6nf91XLC
iiI3SOuzbLSpR1WtNjYQ2NHiQv6TJrMP8ttWHDq8jW+qnb5ac+5wVwGDD1Fj
iXRcqHFsU6khHXfgjlPPu1nvD3nHkP5Dac8NAuAB8WzCLWzqCzQ/js5rtWPr
qoXsGywqGZRueoZ0h4EkSdcxs1PqPHcuLO3nisViaVJtPu7hKC+QP2KU1OCA
DKr2Efx7qzD6Zl+mPgeoO9BoxyUMShiL2n1GlmCoGdFL53A9j0TkieC2b15z
wsT0QQrNOPY5hsE8BYdjyeAqVv5dAs3S0kCmSqpbMmRgJZqPNuhpPBlHexRG
342ttp+jpDE2B0zXgrTDIkoauLXYmpMXk43hq8yMzjCPyRhJIS/C7mXNRYRD
CzR1rUKEqWtLsdsSo+NlkxMEctR+dTx1jxih3tgCQ0wcXgwfczSOJp0IqzqH
RWr/bfmsza2xWTAqUDIt3fZrQW6OpOOSU0aT66eQyOsRTvkCCO3GHbub9ihQ
CfLDaBohBB98kD5emh5QvM1iNSND2dejOkco8UOy1eG1Wfx4gXyxGRYlA0B/
k5LR/7ZpzrU2DUL+yXZdjrzfccHsrdLJLilmpSq08hlQ/ZycFvADXgq1laNH
bKmz3dtpERHVn0Yc5t1PsjdvR/XY53iI9kBkzuKzCA79UEgZHLSpwzFwAltp
6JCqzwr1Q1hkTqFHRWYHBwDABFig/aPccPjrtcKmiXS4yyyIZhSWfW2bCgYY
ELQZ3BVi0jYWyjJZBze3M27WyRzfHehN4iSbHbfleWA6uTvbFmIqKiAgWTRL
ef5P4jdzqiE13TCfO/Mja+C1mFz9sPVC/xsQlNXxZLymTD/FlDKRnsYlW9JP
4JB+boDKOScXIwIfS+3Qxvb4QZ/Zrjncn7H0iPa62PUaYi/UZhbVeGMycJov
vgwp8Z9L/ZMX0SS6zcajyY1YE5GkI+m9qvQdYzY52PtESYPkggqTXFQsCu/o
Wj6NCgBcLN8QiyNMpuDTJV7N64ch/JMZW6SDxQpeijQqu1GhYTUMHQY4BbSa
MzOT0++2XnbflFzxoCD9nDX8daehX1FBL9sI6LlY0GVc4ALnNXQQhh7/ZNau
IIXMh2ljaPPV8BOI/+wYkvAsWdUJyvMLwP6elUgZiIZnMU5sIpHI2TFtYYv/
+vib2EIFCipPBRW582ZhlMKMa2WI3zKkfZ7VgqTdBTScn0Jmj34PFGbTiVst
zIyN9yNh8/vYgtx8sahJyCWa0y1BETulXngg8X/392qQmi4o+R77GXOumHw/
y35rCy3wFtlmaPw6NB0mXS9KtPFkhH1sOAojAqgMq3iXPQhFNsGlioVwolFn
DT3uk9fGR7ZK6FRumx3sp4LGmEHaY/OiT4tiyRpG2r+k+CRft4Oiw7xv/13h
RYNVuGG/XdCw5iMIHc9nEee8PsHbDv4yW5DaxTyHqottD1xz7zkuZ0ZPTGfK
uQr8/NUGL/KhiExEq1MTnjSIwFi6Si4fPCx2Lz+oHEtqXkc/c9TKqPSV4WQc
nkOkCsA/2A327QFFVIT+gUXJ06viRSkedGkz8CdvGTsd/WHu4O+ns6O2AGXT
NG3UFZCUx2/B/FH8kpQTA0LUQr4JkptQ+L1MGNTzWtoK1jblc/zEaXwWNdf3
MyzLMXmd4vgVow33Jaj7VyZU/zxJ5Pzy6v4VbB8xFeTARF3kW6HTylmhjpyB
LND/M+jm6XqHMZire1haCNwXwVfCq5QW9ip1pVAtfFz3odecLYIMoGBolxwK
I168v8+K+V8AFwrIY4krWabFPKupD+Q/7TPr1MbneTiPpMVaXq1KBRd8xMeA
ZcftDfYg/d3N605L+TB3/0S4ojtMQd3Ul4SZTZ2WwUVAWs4Hr4FzdWnvT8n3
TypPXQK5afpj+Ew9lSCPptifVrDcwhWqKwV3+pUG69kEAEBlY1XSetyGJKVR
f49QUgJELRh0pWDYfJ9zFrhRfjtQk4CoH5bhEO43p58Vn0Doanan5VG6KT57
3IbOyNox/Po/2/8PMWLWHmbNR9cBMY/PrEd15joa9wA37x/O73pj2jPswZAa
qY1H8Jz/YcFAkxT7BOxffk56bZbITh+4+Mml1x6c/L2xLYEETluKfg1IwuyE
zYqiVtAs7z+HSdJFtsLG9FtWi9Dnnf+Ckjf8iEdeYUHEWxsCCiFgQ7L9F2dX
1Y0P7BERvw14xDu+NSs45CNyKskzB6hi3A7T3qGUEZpMWP4nuTDKQt+T+48O
ZUED9VbT4w3aBtw1LJ+VvI735GmbGam0OBPMLsM/25US96GULwHlyXjpYovX
EaBkdD897gN1/MCAwVnNNqMwiURtswQ6jq10doLv8uUw6m9YIPalASe8/QbZ
pS9z87y57O8xX/t7rtKCgTjlKEIc86WisQmW2nq+3olbRIzzAuNf8b13Zzr/
nXQjDq/YN1ZhqDOCPr5E3jy/nJGvjN04MDQhWM0NlbvuPVTFQfk6kCj0CReM
5if5iVEiNWWcCGe1kBottZhVjOETO7ACgVdNhxua/QBHvfa6F8iUASVKl9U9
msjNaOWbAa/1fOImyxFPfIa2XrwrOIm8Vjboo4vgiorLYrqQW9KRj/61H9YH
2IHXh5JNHdMzwrYqgmZv55Gp8iKdCrq4OUzo4vzJ8CAdCcx6/b6nfSfe0Qnu
vr2InUqAcTeWgHoZ3ZWNt/Hb56xSrsEp0guHvBqCYEqS/7uLyaDVJ65auQb4
d4QfwtkJwD+o/3+51CIOYXFBXqGHP3gB1rCE7tuhBE2kKNDHYwJE0Yspn1T9
9YnDwaPxjv4NbqNoRdZW9HAHu97tbM53mksv3dAGGP9sENsbbQH0ZXhjz/Rk
DJUWxDKIYi4I5mOxjbg6buY++TU0VzrhkmZK2ygFDobWbCs/QQMvfFYWOBiC
fMHhyfvC2/Qq3x1jUvZtIEG/JhYi1h/iPAN23AtYucSCUij4C6cVYuC8f3zO
iBIAjPfH2OTnK2qU+X4JCSjGotG+a3zkmiiRwrHOiJ/T1ai/99oymJu8ruuP
IDcab1JLSuQ2CytC4RbSPEgQYVAXpQ5xiAjgm7hOVGogst2cPActPUyuw7Bq
HHmsWH7epLfkwF0bx5WnC8w7cot+snT+4BWIjxY1UXh6e4khBUSZ3WEFKZ4K
+uaoG3onJypI9A1lmrrMq9rthqw929fm9x2+VOL0TRp5bONAGaCuhgzLEASr
Hp5POyNym4pjTcPDaJ+i3QaK271EVxXIUIZ0XkF0NXbtPVSYtugO6upkDj2f
u/hNony7SeTy6lCCN8kfQ8tfOIpKynaLtgcsqg4dqM6l3xtbXlvNe7BhSYdT
Bb4zU7a6KU1CoqvHSO12OagJl/TiaxoRkzKUz9JYGA0JfxymFHaQiXu9jz0d
mKqobSVGHY+gq6pKrb47mR1q3I6v4sr53frR+od/MTVT1i8C7r/TBdMrGdJw
cWjWq2KItv/1IU+zq+57qO2is0yjFckjtLQDoxVJiwZGnDMosQOG43P4Tbc+
dt/HqULpBbILGhldixTBSGBqP4wzguatCA2qjtLUugnDc5WUl2LNF/nVwgoz
wJb04mVD6FN/Jxx9AbTiPaPJDowYpfLcLROQIwsWZm/DE/Lrb17p9DHd+AG5
GgUJ04T65EylkGPD/QPJyFcAem9D+2KncjlRzFmb9qddOSwG5EXyoKxdUmDn
kVCRdoqfIHB5agkdUzdmgkOEoI41L1x6cHD7+sHT+pJrU3T+cevSwNXfEuvD
FUFAPxjKfL4j0JZHqPPKS7yHsohCb4K2UDJmarKbSCR3OB3vtzSYnBh96hbX
LOQ4Fc8Xs0XoK8fRogel06p3pwHHSxuBXuTt2hJIY0gkGsWw4KNyTNdGUM9P
s5a/MRiTXISLdI19U0N7jN4ja8X77HqnhYBKloXYe77mrk16OTOILErnSw5J
iP4OxKz1wZ+6F/1N72Vx2WuI1uTG9E/WQsosOIa99gR1wz2nQfUm1AoeIMVy
NNK39k5YTc83RmI2sha1EFAt5NiCG5M1Fvkl/bRefRl775gLFQhUJHddmWvp
3XsDRVENjYWU+u2BsGD2sKoh0XjoJGGDAq17moGGCfaj6fVu4gIdPgOAAP9Y
6ASh//j394JghFivFhYOwokJMxsV1Us9cD4cqKao0a+WGAc8hBkIyh3TjC0q
I4ekkW5W1iz8hr7rfe0giEo2FmhD+00AKx1E5p0u+a77sxUIEGasoVdDN444
BHf0auIOkhw8Wx664lJst5tJjPKdu3G0qf4QOSI9KYKjPkJ7kYVaRLMlC/Fr
vqXW1pPgRdDQU8cs/DIEZev0WPChDlAvnMRt3pSdIXo3JxtFMCWxl+h6o2dw
LbUhC8Qxmwb5q4c8GbtJht0dkxDQlSqeUfXEPdo1v8YVvMvP3CX03yGJSM38
K3ZDyuAJ5Cs3xk1UbRsVRQgye+UrAgybHqeQq/PWjk01/D0TXZ990bNBh8ze
DKRxRmFhVRGVrD0+js+YFXU29uvRf+4qmLjDEjSTedk9JCkPYCDow6mlEZrX
nlfBzxymC0l2nKma3whSYF8czgv95S0DDN7u/WKEJOxMNZa0zn219GC6gyME
JR0HXrMspEx1emdAsT0Y7ZNJSH4Hd+GGr/fiQzstfbHnca7UXLZ06QRIxAzY
Ak0NUlrYLc8JmUieYdbKVxSklqmblGt6G1vK4QFfxDtBpAm6RbK1Ol1nDgx3
lQVj0fENupN7bDwXhAIljZYnTSsffKzGIlDvUIahEmyRajHx1+1lq+c6p3Nq
HVs1tW/YAA8rsWPYfVqWK3cac5OYdllFpVJ5H3winO2nwKMhpgYguD9sdW4G
O/R6f0a3zvu6GCyt3nE5aZX6EfuithF6pMw/l83tnSiqUVPEJ/aa8cVgWnni
VdmLYkT1iqilQgbd4eXc2TLtNwlTOtkTIG1xAdsvMT6pSqclwYSP/djIkNr+
BDucRE5akSfghY2d7I0YrWcd4k+fXJzK6hHAf9cqsofyHrW93FWskjM41TVr
8rIaurB609juP8maiwJJzBCOMB8h+329ILhoD9GB7qOvSMzmnOUfnoastxTp
z5hkyaA0H6NJ19Dq4QMcNf2M/Cq0o3cacmIkmZxQYSNbXgLROA7GPWj35LWF
5eoAzRDfvVkkSM9kgmJsZZebHDUUPBZV7q3YOPK7VIvxlNs4khNaWqTxY8UN
g/kXdKjnGEOF+EFkssKhkaFQrZtUWKAhtRQmk48lx61xTI1oCXzeyO4x6xNR
WZmw4liPbMekimPRr3EcXiHTHj3/idPBqLP3XPuKsGB4HOL6ne2PIA/vadG0
32Qf0j21NYpZF8W1/A8wexlm/Nr3Arvf53zC9d7wGXpvnymYe+QL8wz1RhbW
mi8y0Eq9OGF8CTtRyuFjFKYYsgcJ9hX5jb7QRvAkEdpMrsYK0l1vEqia+qEL
romdCWAh4z44Rvl9DzasICPMXLb51sOVi7FtmigA4MezUQ4jUAGf61aZLc4x
FNtAf5diwQvfPAkkHojKGBvnDK3fGjOkXV4CqvuQK2hAndZyVQZLw/RSgxZQ
Y7dA3O3hAzi11WunaQDbb0MoSI1YEPmnH0Sx4LQ70yAzXR4ws8SvDabdVVn3
FjR3kwXmJ/e4eawYfCpVg8gkBejYi7ed7kIv6M9TqQR70CENPtuGv4d1aYWO
ihSGiAvheWMet3N+QYYPeDH5ifAuoZdhkm1dzwHB//3EsX+n0Y4MejMbFIsE
9ImkwC0hs0kcM7rJogxwlPwCmK1WB0qeFAbXyMqENGnhO9ylpzNqK/Lpj7C9
oNWK+CTFP7nAPvnsUoNoQgSwUKW8e4sDyVM8JPdxUlqJXuQgsUhyV2kD/sqp
xRZ9qKZ0jRbXaye1X5j5UaFjRh1iNLGOvUT2q3x7xYdLFM8RRgdkBSQ2qF16
5fZMC7XlDIW1kEGrEOLNSpdofBhsqwyTs6VQ9lDP5/o5plUi0DhgbfkVSP1e
+NZ05+ALv2Rn/w8TaIBUQLicLVGexSXx/v6LSIKqygZQ0GzozjyWsP5++xjJ
q4haictrkov9WqEdNM5izCAHep1ZZ7/ebJpmEuE3US7Mhw6BNNbto9TxSv9W
7nzCsELvSypxNvLvIwCiV/Q7Pj5wtYoW+b0GJKCv+uR6TPZ+LKQ/yNdl/rvs
SYXzumFKRmzTxXb0+ByGc+dwj4vpqBnTT7MspqVBuTM4IBzgPHdHjPBO1e3v
rDO6TFxXUJ7V0bt7A8olXFv5lHlRx+G3HZ0YCRy3shlF+sSPSv2Z18HNjCir
YgXWvXCHEMGdxsRDvLCDw7S/zEteGN8CzklJNJvDP78O3QHI/0sk2ZOYgimo
n5SXPE9RjkhCGvoIvTAbKyQQCZPf/IAChXXZu3MUB+oZjcwXkI0JpQVSpbgH
bEs5Y/DUwPwGUoW28Eblrh6C8VP7fokDN7RyKS6gj+ngUrnrT4U4y3Bakssj
hTFCTQHNPPneQzkv+feO/yfCLynTu/ZQR0mC/ziuIvjWwrH1WvKWdOjpyjSU
2CiNB54aYXnTn5oGpIDsG8lg6aSr7yKKpD+P5JVIBK0e2PmhiDKVuXYG/+3H
uZIb2tXRLSKINVxoDLSSEYasadr8iHKxEN95bw6FQQ31Od0y22q8w17uWscS
nUMgbf2r3u18z8Vqzi/eeR+JjbDw3jMylX2POJ/yDHXjLA6uyB+Crvhr88zS
f2HnJKpD89bGp7kX8y9JdvIR96fDgnGWf3oDlgviYbnRSvW/exiPCGNeOCAQ
Uc2HfJ53l8ksFvHldWVlUo4okrclNrgZe2tSjENwyr8gjGvzh0vQcNxlwT0N
E6H0+u/yk64IlFJ96ziwY1VUy8r3gn7EwpcplLavBPvOQxnt3Zb4r8HXFTKz
fDZJmNWvcY/wF7QZWQmS2VGANT7jY9rBfGwg2b+5kwdV+2G+TI/LCMlvuc4e
biDbi/RrQCuMynTnrTKd8JaEFKbHhXWy2Zka0f6c1exd7TtPXjqQqBAZsGjo
FMDP8yDgaTednS8fTz0pq1hzc0uqB++rgmOhuDgPQOPnMe+REH588kiQbPQx
rFygFtVQwpV11Z7fHC4eV0E7sZZFS5DeM3K0mRO4O9lWCx6zYny7PM8qEpRb
AniCieqUSmdIgPfQMxWtySoyqdYAgUnn1L2J7KU9zITKSPKFJFkDHmaGzAJQ
n6ayS7vSC7a+uuyhoSBpo+8nfSmbsWNxUnnA9kP4JEoWP9qpLmcYPiKLMU7H
FmQa8CFzd+ud27+ttAzSS/QLWiQzI9EvbvdTmNq+oYNQLrfuxJpb7zAiXmrd
DzaKMgu9EjDxyixRVSnWiJbCbeBKw1O7NXAGr0g0UcOIJ3ZA4EAbGN7v+tMo
cQdx0Y2laWsFMQZyJwPfbospo9AE4c3TPB8EVx4R71jeKXgL3CSOh+tpw/jm
kP5bsuLuUf7RhjEoPkmlG5+vZnBjCHMaeFER5f2yDdubNFKJgn8LVuJrG33u
wTBcCy81IJc1cyVRR4ybA0o/p1QoaHdNk/WQwIXBaQdMdXHLPomkO9eUIAEb
h6e1PWz+9WBrjX713obleEd1P56goe4K/nhHpX1tJBT0GLRzG7ZMmzAvYKiT
V9Dvggm6li4uSJgnt38zBXsxDD/TS+j1KaPcHcejF5NOf5enSQKK1CUgRw3g
Gn6bPkwJeZjoaCCEnO5X0vH6Bk6gG2fQp0/jTDmQJhd0xdPz3eXY/yu7qqMc
V+uDjtjdADkE4qR0XIAUljYWhzwDXX/Yw/nt2oW880cW7RkLz9ObApbKIDjU
TmVXsjEMaGy1d3GLHQePgmax6TFA2Z10+t3Bnuir58fOlx5yiDtW24L0w2lT
tDzkAiDPvLG1Tt11Vt/UO/TAiMXQhqLqAdCs/0/SBRqFonM9jxeMtLBNqMGh
BaWgXSdxN3NTDSLZ0pEI/ujsl+CFl13g9hgllD6TE3GmT/vTnkM4DxYO8C/o
5ekEtSmhYul8BErW7VGGNNEPjwdzaWcG4wE+KpKfF7LqO7O1nijP9l7NgM70
uW/6leNw3OGvoGmVbHybN2kHRnLpJV0IEAHkybQasuw/JcXPWN9dtYvkXjrS
GB52FXUz3LE2QYhLBkEEZzDMgcbRQZNnChIWkTPvhwEWZiVI+bVlXr9DS6G4
Xv+ALEzoFCf6ZYQ1IquaiV9VrjWya9yltQi9Rthbe1rn48lyeJw7LT/WZyQ7
UCgiq0fvAH8zPqlLmySjJJGV5319a0LStiNOzN/Rtp6eJjS2JzU76eXyx9pV
6V8h/bOnc7GjPm9Bnqhyy8ibWcQV8k63rT7fTmSRv5g23clWbojNCeoGnSjY
gK7S/MMDrQF9ygPw+9wfobnbJJ4bPs5g7sGYeU32tLFwyEOJxMa0SrYOPUx+
igG4XfpmxWjhaKUOJfBjw5s7Nf+55FYhu5ImypSPqjbbCm0RPNX+Bs6RrBs1
+7FQp04QzxnOWjRrc94ehaTCtroo265w7eJPjRcjgHZWkF208AfEMTx51Sda
w/WS5t70AXa23a16AQEBQZCtLJFKWDQ6NCjjT9A+b4u3vjGX6mDi2gggzBIb
+caeMR9TceaYuKhcapQiDF64oLKFPIcxQ3ZyG1F8pqy83XTd4WNDDAJtcUP0
7cnjlyAzo9mF5qQVgVZ4f79VJA9QuzD0XjiLg306CbOLG1Tkn02dcW6nvXle
3d7iKnQ7E6ymyRB6UznrimsAYUH0x0eDIvnpGi2Mij1/QEYJb9IlCFwjdFzq
SadmCbQbywE9NirMrsjHoE+n4IJTYEZpGfq2AbatE+sgi2bDtpNU00HOXGNc
zj/E2QPeOyCTjky7hokd7oCfnFjA4X3eM1O7rxr0uh9N97r0t3kH07NUXvH/
wzBFod3kdMMw+Wmqft5XQvT5ZtPyEh/uhPT94o1P3U9CrhNSFKfQW5nc2OJ/
JlQMrxYO+ydZI8uPuyhZ45aBGQv/6aGKhTVW2QRF00nF775iUY9rGpbUutIg
kNr13cHAIqz8QYu2Jeg48weY+EhlTBvnQbFikMVZFuFcRc3lNvvTHa1G3vMf
mrBpjIOsr3CWVaZD0ZnWT12c6Pf/Oq9scXzRfNFtZC152PuV9ueX7/1jNz29
c1BHzqsbxC9jBpF1MyPAPIynfT1dYQbugJMf3DF7Pu4VA1EP7C+k+QSZ+Bv+
wXsDlXW0CPOIZIzhc72iTYJRFN7Xg3v7YQfFR7mRJwO3jStv03lXeEn8dG6b
SEqgkKax03Rt04Fs9uXLbmdVhRlbedNzlbXoB1CzIDAvE9YVOB3bvp6zf2Pf
OrjcDxihxEZ2OEZMWNq7TD7mqt1YSRvHhE03TjTvxBh0/fK0noPJwmHZ+0q/
LTARNsTbk1LseT8ZPMs64gSHK372uopJx6jdJ+Ow2906UfubBFyKtusbE2c2
x248Uk+QoLj+GWq8iKrsCowb8q73F8gGOujd6NodNpvutyJVmFAdxR1dZQaN
i7U2Dm0au6TquBZcmbBvwXcvySaB9cTecl612O0C0+8O4VKUTBs1ZD+2z2cL
rM3olaYnK0gyCbtfjoOrzZlbei4TciHzSeC9cPtrNZNhpva7rlVvNcpj1iYF
OFK1cviJKB74wRhDvvNcvC1PmcAYnTWd3QSaSqpw2fYU8kbtu5xc+PxFuTJo
KIFoiLwgmKWVRJ9+IFyL3BJ7PmK/gxPi5he1UzxL5oUCAQT1mFugUzR/8z6j
by7Lg7NGaGae2YZbZZOcf7PJMSMiq8BG5CcZeLFiA0OVK/D0CSamezsCWDEF
n3KoND49EnzbSDd93tG4QnQd8Eh8Meja6OeYMxSlBqfP1lFCQ7mswoz2h3k0
zLgkl2ZRZGHDKTu3CYaQiIeDMC8jzrWoNINgQluSUefzecplwDyXyC+P9Pgi
MtPQBMMAYT2W4CrBNL9S+JUSGcaSdbOxM0wm78jCJWkPV/4HyxdkGUap/sov
JJXJFIMycEPJ8/+Iol5mLkWzhthsx5znsTZ03w52LNXzO1qGVn2daCUPjj+R
CMA6U4CrpDTyxZvdDSGf7DuYrvJ5FWQ64o5AeyGO9xDMGcjXZCMr8XRcmvAO
onFPdOJBibw1gIcessTKsg5Z7bFCrqbUBI9DGEppBYFsfErYXsI2w0oDZNIx
b9MThZxI9dKtXws1tMDGxd9iWduv/9/dGQTkkb/SRQgp73+KwnNtAmVdFi+K
B/my1WhlEwjOq51kBTt3Ey4NKlZRa7UcsjOvz/K2/SNn9WhEFIl22TGoagXS
ELdi0CNWmYDWEjt3fAWM7G+wudA6+pyVJG+Y/POQOuTrN6Nd15n3eGka05x+
PUOex3I6/fS9EiaanJfxpwopRGrmrR2CUEpTIHkFYqu/S6z5zGB/TSOve81q
V158SGeRZckH9DAORRCx1drcqzB3Z6lt90ccA2kBOu1ut3q4d6aJorpLOIXo
2mOiSgMM9ciTh+4sh0YhQgRneTabdFPH9IfXXdQidUOEpybvJGp6Gfjs+kEJ
zkGFzNv9geHQ107+fS53YsjD4vfyYNO/3PbE6r9mQ/74NllJDXDr8i/C/+hg
gUrUJ+GlYxGBmb6OfDlWEEv5kRoH8ZbqfyuUhEgfHtqF3gPOkTDrf9+6ECTI
qZ4mWryygAdb3y6EW6ImMt/xpwpkk9IKqYHzBU8HU7m9+itAWRtxp0CwrPYl
yakXCIuk3t47hU5bNzeZ5PZzIGTXFOHDMNYAjkka5DOSvlg9eebecyvs1pGf
5/5uAFyUoB0uOpuQcNXJf1nNHNjYfIvxsXEugMSWQbBV3ipkAMIJcn3/25Xa
7vK9Z0WCNK9npTta4bNHrHLkdZzNCPkUL853WPNu/MvX7oYdypZqjKIpuGqL
6Ww7YIPV8IDkY5plOO1BS8WxJUi5Nd3IjCCdaV+2HfvnJacpioNrKqkwh4sx
GhmdXElpJ43QpR6aFptkHnjwP1DX24QAudI+oEK1qS9IriU/T2FPwkzjm1jL
tQEK1Tuv5LeXZ0sRXLe0+TKr3TcDeyJmsrJCtcTcoZL5VMRDBePZp5TgyOgr
qRk2y+o8u4zRs5RjMPuLVNghV8+TzW3PVO0PmkH11Zh8OKeaTA6M/2SWp76U
ue+VdPK04UTQgK76KfmS10CpCsiJRidUi9/2tsh3lcohbZjqQ+3tmmJHvns1
YP72jSEGcXwwq0BzIRsz3Fwq14dczNbfUH0k9ah6C8/3+3haz4skWEhT58rB
TY/dgKMyolhEv2lpUPWXTBiyptbdai3y4v5AcqyMGoct8HN+8PGiDd1aQfHd
msBBRYXoiQsql04rc3AoCbqGT4yACjQ0CrIIgwfIPeFiq7V6Vyuwszd7cSQB
J0GJ8JoeZ/O+zTa19iDJDJnpZMkcqhfR19Qu8gOxxv/PBUcMo8JINUaKQ87i
qiqQvMOqHRpYmJJCbQDuooqUskDs5ZnmX5PNWJjUkP/X6YchpTIm3/3XDcWd
SBSOgAvXqLP0foDQ+wCAgUE00/gkty7WTbb7+nAeIaLrsK4W6+P8OYEw5K5K
jdF6My2CdzF0qCSVkrP4IGtUNOx4HiDkoY1fmH8cgcui4mlsjnzU7z8GKy3x
t/k/ECN/RNIqM6v63++At/bmlx5YzBjqebm9E6iLSoO4SdrNu7GEhDlLuMcW
cLlq+ygOlWUvg8+GqAJo7aaTrblhKCtweFJUyQ9uXPgsWheI9PzirKip0R96
5OmFErEgVUJqiPXu92s+nV0fpm4ESKcbsueutTay9wEjC9omfcHhPqKK8v5+
q+ODE523QYiNKmwDvVWOwdxLm/+lhHzadtW3qu/kZnvC3m0Y0VaXMVbMv+C6
gTsgbynb7SCGoNotNVnT9AVTHf06aTafB3HowwZ7LWDFRpPcufOs4bKN3Cxd
N2YcGhkbyMQfitKp6fRjjZsUaHvhn3+gw6CxPtqjciOwIMfV+ZWXJuF+JuyS
l5MvauW5yP2XVLdZWogfWJVMxxe1IEvY+71cAJ8xVU0BP1TLwBV0Oon8EG+u
OHUXnX0aV1fLEWXDq/qWnWEcAXdd9RfTZSEV2xLI9iGL355PiB3A1bQ1210I
L/xuFYB/+U6dDbV49+tKEaQVK/n3OiSieSeFmSnst9hoBRST4sap+LxQDNKV
7Z5PB7h5LeeghgElFVGw0nV00kSmXO9Emm+sehlGssuYySmv+XBi65fOyESK
GY658Y3UXTxpVrErUZdx+HGfeD9VKQcCSDlqv3q0BTeQ3bRVVWuFzqLZSNAh
WgKaH0GUHW9c76OHq4lJcp8sjXVRDQzyyj5i2llOSrrtU6Fg6atv/5xEvU5T
r9p9L3RyTXHYSwPN1D0tbmDv6Ws3KzavwZM2t4qTdmcYzatu6hfaRltjPRB+
uRbIiNieyO3W039rLlz0FpVce6WhLGWSAvjJGXZc3CEmvy6UxaP2doGS+xKM
JJhWI4wMSAHpouiiIoHx3s+wzksisEKpkyPQX6+66ZDLWch+jJZqfxnHztlk
q3YdpZ++Fut8SH1uMCtyWjcjGx/9G8RaJTtIPWtF3ohOiePcDth0dgnDTw2o
fa8bIoBi7/uAwMZB5ErZMZlLj984dJA5NjaT6c61QKF8LwlSkf3TnBQ9Ty7f
RLmpx93F9NSeKfOq8XGt+uHabBNMhiwXi1MTYt0A2NqcEWzpjrCOqnvX+Ybg
tH+TLXC9p5JuiFuZ4UYNXEqzTaeeFDJEWFPEDZJow4dLXeVGYtL0tvEEbZga
rci4cm6Bl8syqRoAi1U9VjR32iEfZ0iFEWa4mjC9/3IiCknUXi5BWjfPxr1I
90GNOlZ27/6jK6nHcUb3jbRny9xWqPX5HDRWKZSb8L93ewqpeCXaM9go6+hU
yj0bWNVizOw7rkalmFANwCDS7G5ygbPWjlYpaZQvuMtY7CxfR2L1sJaIuKgG
altVViHD+vWi0MR56O6igUjIR/wzBoFp25oMf1/LzOXWWubCCU/pSHaQkAhy
oAKHuHu7Vk7/BcdlQemuwtGb0b4vKw5HSvxeP2ddhPOhvhSF5LTf7ub7MhvW
gt0F20SrXXCLDCifTgMdiim3d0iaIJPerHFayIU1lTKWbqBFBFXK2O5XWHLQ
AryS1Gv6pv4VBYNPvbgP+aOfTXF/lQWrPuBKGsoSosZE9YuEEwvzv2Xgbwni
1vco1DMXRH4LNPyu3RSBlwscPjYWGo0yhcAQBKXQoWdz7gFsP4IILdBKocfH
jU5K4wcHtVA3lhFXo2N/qxPSfE6vKQ8i05sonCvTN8GWo5e7xt+KupXOwhhu
RjmnAde+k+GXm/BK41aqAG/rAtHcs3ECBOb8Iv5zY4FK/fvHb9s8pFReHYyT
o26iXvKHt4HC7okWvl+yK8Mxa7BFJih4609jAV+3YcP3Jw7jc/K/N4vLzfDc
qrDwM0vNnzozPqxEipLwpKnuDRnKwbCAnMDaXyRnxsX2/H4WL9WhRrCOGeo/
hQyy2RT+MCBayfF6LPjXTqcSD00vXdm6Bix6p1ASZi6W+jVEnaMNNd1Mgc5x
ch8khV5DuCXh862V4pht5TgLvlcXaKekqesE6+mHoGYBJ6cVaYeF6RkCrpUW
qiTEq0bdo8KbQ4R9RX/Cvc7cK4yukEOa9WvG1g0PwQPhqz0sMDShWs4lMNdx
XilYuVJLfjkOTJIuWm3WjynZkQo1RV/9bsZFJZxBr4h6nltd58UUnILtxIni
dLs9l3Jl5Dn4ED4dzWWaVIHjuVYmMWYF6mnjteho8BvnX8J9H4lpZkNU0IjX
gP4sOj2OeCjgD9M2j0AKBZRYM5FlPhw7EnkPJ4As1sd57wNsKyHyIN70FNqF
sa8rlWenEqagBsVXufxbskBNLEVQU4NDM2e8cBwhsi/bV7goanNZN+abmYbS
5bZ6y6lPnrekki0FTjvQHm8IgvtwLKWFf3KQg9p7/m8byD9BbuWYq8KcAAdv
LQICf21PagCVfTuzwQuKPLK3yDjaaqI8aQXkyl1Y4gImdNJRXl3GvQGWvHtZ
cgPKglrRCTnLk60oLaPlvDrruZamXgKVXTakGqur9eheIA4k0gvR29OJ0KT0
/zXPMl3Z9o1uxepxX4+pC1OfTm2DSH1B0vpZCjrOqqezRMgr22z1Thb1REPq
VDpmwRviQId6GaGMJsO+mtkn1gqVdqjkq+nlFenwJ/BWAGnMxYhbnl/twNtn
La/xHWUZS08ktvDP1yEcJLLXVzGSs3kS2nR7veb+QI2BN1rZ8j7J6daZK0bu
qITVi7kL2+AlZoLdFP6pxrPPc0f9Ij5IguCnoVDEQr1a6JAVXtYw5NcPm2gw
kZ8/q2tCL74G4BobrRR67dajvjKO8lgOX1bm9JyRVeXnDaPvVEzzi+IZ7If2
4dJck1bWcg5U/z7gJS42C0MlWYQqcpmrzZNJ41FVUiU6qe757nZA7S2HuZw+
G1HY2/UG7wX3BqZSjzPRebTDTu1ZMG0mYRTRq8G/RXJJBBBe+vP6XWadl/fQ
WWUJPshhYMcdtIgwHjmZA3uYiDMJzcLZM8hWYZOcLO8IHuTUCb9oekEHMKuD
QkiKnkItv8KPsAGg3ukaXRFA+iypyJ8ZZQgjpWUhtP/1WSGMujlI9QEKP5ij
AP9cNDMPPlv3qxRhAfdDWLvRWCOzPu7K95pA7fJm3zcv2GcCLpjHtVVgH705
/Hbhzf85gAopoApxx08h+KUU+GsOhu6qs9pvZLx2dQv52MoUKEm67aO0hSMJ
3lb5L2zxOdamvAOP5p8QYr4z9YOSigWYjtoWHfsQ/YSgKh8UznGWqRLYWR/K
yQucKJVcQOQGxld3p38JyaiLb497E6tf6xtsuYBqrLGpL0XfIXLadRcppjPE
Ol9Xm223+ohuDlZQBBNS79mogBiHMDJXnW8ewntzWdbIiA0oGgNWSdQho1qs
9wuKilflr31VDOf2KMgya+cKHJZeHMctx7DaTbj9xmqew6N9E95TUZOUm6Cx
MlnybGg/9i2Y2PXn7UKBIR0hgUQhdR5AiyjZJS3TZlc9Hm85+dcU5ACYrbWF
03ibIk/xc0HVyT8oj/N+VZoITAEW8dJmrks9bmJzXlIqGsdYWi7TcRCQ35hG
jnedYtm6DMz6HFU0ouSfzyhmzgi58JjNGzBSLYF8jVWpVPVs5+tsWTK6OMFL
+mCH/nGp9t2YdXgvi2/s97X8dZbgbLIvP1wUMnWq2JX8CgRrfl92J4rRvw8v
Q+jPQJFjX404KkVQeMc1x+sPCpCo7OBY3mNki3dS1L4hVbPjpLxUdvKV+US4
k9SYFamMjO7X/cX5U07YPyDVTWvyUrdvs77j2D9uxb7M9KIfYLQLI3HXDMTQ
G1k3TpucXUETR8vn1DtofnLq5CkrOb2C4boGRO1ZiJpy4/xjPGuc00qfKFKB
j9bh6BKQ1cbae6Zp/mr+F8nGTFPG4ThERoL5abOt7ysK7GxFd5oRiZvn+z10
jKlHrftsJJbmNrzcVRKIDqtr+26XtB6UpgN0I3Ur7GnQqPM1Z+vFmHwqIEk1
ehdNZLNG7XMNYKtrJN/yyTH7yqpt8dsubSF731vf0IXjNlDVQukfyxF7muqD
YEhZNSnMCuxb0CU3AwyY/c7jgG3gRSwMKYz4l88oVkIEu6U3MQjWrExTph7w
hw3JgjUPqrdhvBIcs+rW7zDbA2yI4sJCEu/3Q7Mcr1cGAAfQOv1IxfiPIAts
W/4OIuN/W59vmJTfz4808TTgMb/yjsB/RzSm2YefVXwqCSE4H//qGcc6EnSq
De/8Y4FiJBUQ3bdTRGfnK5ekE+ovEFSsq2x9a44+5o/xFmuuFjn5JEby+qBc
B3XK9yQe6/zy3r9SDyD19djV1QERABFs2fapqWcj8p80Z8Huv8kXn05Fo1SF
yV99jrem6T4aWQ/xBdvql39+66srVEg7FdHxXotO0J48+XBlQ9KVW2SFfYht
fHhRGP0Ca4Qvj+QS6ndqBNASfO1jIq5kI8GAH8+J4LSABNw4EXiMpK/9JjVx
/cGNBYdvAVtsf6pUSGNOmaZcPyZK6Jrl6pekZaZCkPu0huEil+4h64CQYvZo
Q5cGxJJnCcMmArodbUr0mUh9/JxMGOu+CVVPlB9WqnkQT+q+0bNbJ/Zrz8RO
3DJsSvruf+D1nR0RQ768befFHu2DasDOUlmsQ80qOSjotLq85BI1n0vPn/va
L8MeGPS/AfbZdQ/eCjkzT8jRIgeQoRphaCDMvhcfQc+2lwiVRPXymvsYNslC
Y44mPU94G/w/QmvLQalRWB9orn1oiOVDJJKK29qfiL/UnYA81Lq694iaQtiu
xAUKdkqrq7BzyV7xca+XnzlYqmGXTytMn8qmThhoyfpUfMlVRuAcIlqxtWwF
+Da0HmqSgEyPEybPzUf7oOsrS/ztlAXMV4fgMSkUayZB20XIhgywkDDEUxwd
+vDV1ZJJImhpmaUNZO0on6j8LIt7hvE3S4msw9e8S5vawFYNIWymnxeN3kB3
MCNBy0LcQyP8PQpI8d2Fm7wzKwxpSm3AGr4VcpbJsR5ncsZi9zF1NVqz+lTX
a6P4humlZIretzBgiGoPYt3c9iWEOpBoXZHnkhadfhb5d2xU9EdnCg7ThPEr
SL5UVCla4Xu/Nei6VHIWRkINzIb1TtIfmHAJaUYDhYeUjdPfHWYs750hiBwa
9yg0T4sravbNhOw1NKGlO6GZJGseCXj7cDyHkILKIpoZpmla6cPyc6MwbN0v
O9ZUau6CBRl5Lc8J7LMPpZJtNCDzxqqWxmvbVaLJY+9Fo24TLHmG4t4vELcL
DQSxiyp9DpCLTuEKcfxNxx01aMhbUx3IUrd0Lwn75YVULbSNfL1MDI7WTCVc
YvxmbDDaIN85m6y7yhpqZjGeg6KL6AIpyQCOHfk8ymgR1U1p7a9l4jFtPghb
c7+ee+ZQw3trI4FiUIhPJQgHLyJB5sEi1eF2A3wifW6Lf21tqITdVRzEdsi2
T7t5BJYY5xPcBW8PT2APIpw15z4PTz6/VAKcV2aV+nPCWlI1/72+nHS9vgO2
7ODSuCgYoZVzxIlouZOLJeQXBLQsJMmEm1ptdonzWm0XXzO6BunFm3N6u6vy
MC4rhLetjDRUWsLv9q21AItU2b7bDziZoH4z3n11j01TWlcPWys7Zo2JUMx1
LoRH3uFoM1YIECGv2plAMhvZbgHvQxkjvd+yyu7kaY7MNnSzEhvJgW6EJZD0
p8dMm3yWut4GIyR+2v1H1O66NNJgKsHle+JR6wQ2IbJYHX+nXpYVhDdAgPgf
it6EZOry4qSvn/7KBDxcerMYLN0poknaxBe/O+Od2N+Wo/sFYnVLwf8ql+uq
qyS/1qPj1bIXLKTiHEkoig3e4cK3L9Vg5Iwnp3cQWMTZ2nsQAKYrJc12Or6Q
Cio2Yj71KuPa/LO1I32QPxD+Iyga3rNXSl7+rZEHv315WEDNlKoo8i+aztMn
6KwzaP4HvrEs6Q3GMbBP3jbVUPX+xFDpBEOsbIJBpbhfuHT+logQgkLgr8Rq
jooeFAboOIaL4AP6cstZ14SCaBcG1fpg+zmA7woPDXESnU0/i+VEwykh2Drl
ztMn81cr0zXynp4nvvSn2abShKEBCjCPUgu+K2hWFP1HAUq7jjN+PgfRwshP
H8QBcz3L0DsaPwV5wsqomw54ot5BTnq8iccPyiYJo9xZ3ZmHrSij3Wy5Bvis
6d+t/cew2DqG6PJ27eaEsRoG22xx3YC9Dp40s0ZWuxvq/Af3h5X6eLY56ThR
ouWnDbHlOxLKsHgTkXImZNqV//7XIJB+7lXy+p7envy/fl4IcNLD5BGklGUI
nCkcuWFfGeh+Wd7jQFFV06HUJ20h7r4QEaXmoTfhYgzlGhj/ZVW0a/c2l9jz
Twmra6B1L4iOn/7ydlURZVlD8+UwHNoNqs+pjecUfxB8QIWjXH7Q6npOLwf2
uSr0unfX3wsaOcQJY1HZAQhMCFQjAWRMkoRw9wLQML8BJlP6p5UQDeuCQIUg
vSduRjEM7iWo2UE33XQ/2hU9abJjoSzjG4dN1FSUNwMyIOBgpwiBQHIEuggH
yCWdx927/wOhMEmbeL9W9yAR4Q/z+XIbcpGgQ6bkQEjtJiDDtFb9C2POLGMy
E0mS5wsUXLxhOAlRewFEqkOzq/kEaHZideehKDic2JUkws0qEFChk3Ni+r3Q
nKxD/seGhTUTqIEMITWg9wJjgX/SGM1/r/EUn9+lcTFIdTtdz4R4CCEKN+Ao
QrXWGlvllMpPkS+RtcHhoEZ+t26shqNhb7mXQDqo9lAFcAyyEYQp8xT0sGcO
P7oIp8Gcxaj22VBo9MvfZy5fVcwcuvu0iYwewHfLIvCYrE+hjbFd+GVgaA/r
poQCgE9pA5yWDqSemGOgbXE5SEgpvHQ1H/zlzyzygdBLWuV9nB/fpxt/z2jH
vtXYpkrbDEl0HrJ4O+xC7C5zeDOs0HBW/iSmmVOevjPh3tyoCaU4ytpKnwtk
jKpqOd7rUthKZRDtcXT2lmYF6zevFP2qpssUJ7fDOO9WYmU8ylqjpbdm0yY3
Um2SSW7RNtaBHFjXFLVxiF6hl5UsFiuKfA12YzpZXpBZA3erXfACSszQizRf
dIAbLJUfH3Si6HSSlljpltcbDE/yaJDF8R1/mA/6oKKKZBGGDqQvCl1i/sHx
hLJa8vJJEz8K5mJVhMw7kIb9/4PGnbqzXcrZhxzxF7esj47NVvi+Oqw8cYAY
ScmX4DklBLCxrw5nsQpLeeO9fLsocTRgMCVntaZZme2zoGPTTCAicKY6k+Up
zOBsJq7Qyoo0QgL4w7jphOZdI/ei79kPXBZzRNXUgF/bIQcCCrgq6nrR5hRt
ojeb2OhC3jvH+oCA8W+ZZP0NATZaOOpEPryrZKF9WE3evN52h6C7iEO2EcZW
LpqFofNxfYiP26ynYPpN84jmhYMMhMZ5jdG46TLlvQD/YCARiUvvlB5TdBI7
HN+MYnqACYfpQBx9FzwULgbCTe/tICnrTJzaLhs3m07OFuw8GLoVx0DB0q9b
Mbmcy5P1RDr5CE0sgPVoElyudmdqg+bE5rLt3wj3MhkoSW/SveCZySYkiOOp
eXggqRc39Pv2uPuT/4yzz3Q39cYPlP9vBLc5ioWCODZewz7d1moGT33ECTsN
PGsH8KumQPOzStc20vd8GbuVKkpqEWC2W3i2VjfqOp2oWFt9/SK0YNJTBkGX
cF5+Kash2MpnqEmrqS6zuN36c2AG+hbsmKR6Sjo8RS4ao2g2iLTsgB4aGRtL
XYtcO7E2AYrbLUMi/LakDqVinotoOkjX+xmudrN78rQ5XI9/nz3037Wu7P4A
W3UworkkFw+g9/dssQ11CIBHxuu2/vNxeLUqN9ZRXmuag4e0CoLrHgI2GJye
rYfrpGG4Ygnk2oKRoyQEYTe4XrJCOFbxsnU+akbbnSyBRpknUrkKGBdK1tlM
J5+MpLUz1p30JLYC1KvONfD41u9dId8crT1xn3iUsYH6BtpphnELxi/gihNv
2p408r3MwYMgnEpVPf8Wo1dTg7Ca/4L0VoQ8QGvtMTHRLPYx2uJKd5m23YDY
CMl0ilgC6FJakvxfeoq6gFbExnJvrotCLtR+SMdgGgtjPZvFgEgcRMjcQ0nt
2J6BmKgn5MYRLTUsYil0ySOzW7qnMnuxTBveqf0+e/vXsiQVDnDpl86Vajm1
xZSZciiqKF7Dt1VIkhyjIemjup1+4TWvrweoCbnHMuNgrzYkrARtu1i/vkBs
muo9wuW2iAcshzK7oKeRjTax5gqjn8BS10y3+DmMzVzpX05aP1NZDkDUI8MG
G512lMFT/fkgKUnnDvp5DPXTtys7zET9iaEqE/r8EwH7hE5SkF6brYG2+jmN
ssbK9kGKDlZ3lrqpKvRGcqMLAK7WpBxrxF6NG+oErDmpbQOemgC4Qxkgrsl7
nXFoqfjSXZQH0msWCwMAud+tGLaBWLxncC2u6RQKHny60ZtpGrbftQL9cxNv
ceQKHT1od1yv4xD//7G5Z/z8Bh8tphpwuRHFIZZu1jk4khsG/kmgeGe02wkG
PngqleGvxgFtiRDw3MR5vC24Don9sULlkUVzAegvqw2/SqhOet5sMFeDdOgz
xfuM6S+9QvYPYPQUrJePfeSPHMIPiltFLNTL82BjACOjcg2BPDqMjM51aoit
/ONwbUqarnizqg+pcB7+a0OTOcjdNd/nB+yhJeJzT4G4lzdnkcHEkB4zzwu9
jUC4GjUV9qMDStTsfSCLoFpawCuX2S6fbB7g7QZCXSptALUykEIovQNydYfq
676sehMz9+zrQJSi3HPSXyqojAJR0+GtgjaApJpMqzlLmnPnRwlsgpYu7xqG
U2kRxikcnHIOicJsKzZmDTEFloVpLclgrCXBcD6YqjXNHZVWAUcr1vrrhhUD
a3o0GpZc1fhAYFIQsCyhTjd9V7iC1uSEd0h/aCUbNBIkATzF+dt532ZhJVsn
c9FvPlmEssW2u+KoBaJVBf+7XSqBoSISWSlf/xQQZd3nCBlsLyWW7tn6gKLM
Y1kg3ZjFSrWK1KKm4zIL+rFBVV1eU88JwN7hVvr/JecAh7W9f/t3oTLESIHe
WTbujq/ksNqYFVygXAh3xETS/8b70HsG3wDueaEu5LPUVxYsyKbK0JQIhPep
rt0Fd9ydom0ZVcLElMcig6pKwfSQHZ/rO2tydnle/XKd5XtUlAQ3mODfYurT
yzEY76C65dKegjuHa05VQsxc3K+TYyyvPZqFEFvjsSkQw4ZpUHGaAFrNmReP
eVe5vmUw0Up1JkEBWsLGTevPCG/dja/mPWO0F6ec/kq0SOm6VnAQKMFOrDhQ
Va9ZQkvHiLS6wE2nTo+4TvhjgM/QnXVxnCOXH23Z+gAyZcg3oOmv1McdLXy2
dU6HgORXn+w7xbLsyt5nLqBdlUE4g5DFIdKKsKDk4e4Oc765ZOBQvSluy744
eTI1VT0o0KLXfzAooErfpLbBKZ/8qOna1DasI3NCempWMvxs+meNYheqYEbL
3QpqnTEnZ6cZd/HiR5eNU/DSJh50qzFqG06uKmSI8i/0CBM8SHT3ikBhG3cC
IQ8+jc1fwmeYJE38JUCP9dPDb/ryMypIGvlPsQXHTfy5KG1HMUDDhRi+OUGl
g7pFQIUT9vVdr6yVkwYIWhkKOZhCs6raM2EQnrhnN8YrfDFJCsqEkaa8N8dH
IZURDqflqDsvFXhLx1rRjULJTSpfqeTZ1phxzQXFDTr53PYGOA+Cu+N4wJV/
PXUPvMPCP1fW8RMKmyvHV/oiDQepPbD55pPqlK6t9slLxhxgX4DTZfqDaBDo
0//AfrG5KmnO14CSVkFKd9DEc00BGGAqcsFZY4l/sCVa+MnUo8E95MgZ7NtA
mDd9w44NjAA0Wqh0PSHuPO6cwS4czFDRHjv6lL9IzBIZaWzEkc4MqCnZhqwc
l1fWK2Wt8aLkaQvH6aMyoNJBeqzD7cpfz+H0/83xEyRNAP3UONgoAWdRq/Z6
CpUdjafo98KINjJt+YmvWCanXLn9QUvJLsdYppPTmE7DoMp0AQKqxjAc16xi
RpROPOLy/smAESqisDRAdSzQDS5tG9daYYRuKnXol/ZyF0V9WAYrMecfhHZ4
2jiPZcjptqwXsitEcxyxE+OKEVIunmZHBiAWfwt6eqGeDprxobrsWF7HXZuP
paqLRMckEfVGPG/3x0y0I+8bU2eonCxO3OXoLO23CneuLd7+bcwCD0bAv49Y
8gVpmH8ZvY4KB27ll9IGgrves59dc2qn632ASs3FgodpbQ9gEn8O6RnXuaIy
xy5+5ts8jmg5y+N/u8K6mmoLW6AAwO4+936vYVIrlPUdd5ZIePDN+zABTNMj
7a9ZD6oNgkRf81WkMmJwXTFJmEiy4+Wh6mJL9Olqe+EjO168heu4n6rPL8nI
BbZHxFzCRfjTTMaYYojuR9OuNBbT1gGYJ1biDamEMNAhlLxaXSeL9PhWgNA2
NHZy4EJFKZWHV6QS9sw4rSEgbP5TDAfF4uR14TEqy9i95uyXF6gMGTpexQpM
8O9aj2RwupXrJE2ACYmMxvXQunAlx6jcepV6o3MXgS7kEbhu0z1SrHWvh3pb
Cv/YIL2+nHu08avyoXIQlI2M283ZFfcMqw7xRJWeCh7MF8WzMtlGIyn3bEAl
4Y0vdlrkQMI2Mpdhf6SlrQsvc0WD8brkxRZV9XiJjtOnHeQznn/uZui83uwK
BkimgiurSwqNplHwLfJYpucO3hKSq/PYGz9rgkDXfgB2v9CyWMPp3UO7aetJ
Ta16IhCKZMfP/0QVLtH7JNbT0t7V6ZVhp+rVYnRixx9FtNCpkWf3mg2HFzCc
jQkdEpxVU4ThWPXh9cHgdIjOgVKuS/Np1L2BRSZridpSeJ3rQyhRyAybt8xX
ZS/+v3Y6WscsmVr9ZsQ/Qpedoq8EdE2T6ehAFURc/WCYqFQ4qbFxEemjg/IB
pXBz76lO4AU+TK3SC5Uoi2hfPlErVb+olwxvPak1a82OKmhODC5hkYj/jYhs
Ug30GETGRsOYQjmpEY7yKr1Y+zItP0eBn8pdaq+PozBcxW/rscXUsdCu5+by
Sy3PUoppuIO8IhGM+786wImJs01qfhWRHuA32pTcLS6HL1fYZVDBJFXz8+Cy
ZUsmQA6iipg/51dsgUsCPoSES1DWwb0EF82umZRraio23C3dIzF009zrHEz3
wVQyZGbZU1C/+Lgkaeq/iVnCyjCcNmtKhC2edMrHZ5EzkIh1c2foTtqy17yH
Z7TeDJL2LlIGnMD9/9NRzHDLbQjmrsAP4vSiygQ4Fsg5DWArnPMV4ZyE7RtR
ogbOD1gR/RwZ3SclK2HhuPPFvJJRwuJKuqQPxG1AbbywhNul70DRrpEQR+aC
G6l9BRPlyatCCZwSFXX21515R5dvIlK+ojBxTfXa52924QdtlBH80wgv2W9H
SS6EC0XHw53ndG5urD6DH7qDXmktcRuAVCLCvJeOXRTcCi8ihSSFPtwUCNxx
jpRGC7w4ec3Leml0tcWMVthh/JQ6xAqr430BoAgm0oYfRn+RRhVb2uOHYPK/
raeqrA1QZrhH8LItt57s43DiVds15Rp6pEmSUK19uM6W9gsPu8kl7NbNiZad
KMC79UuD5QqEqOze9TEAJLLRiSurZhW7cCUl0uyynMp2+RfxsoNxg2wBKlUB
+J4zko6yeTstYj5gqNz83cj8tR2rRoGilw1Prmjz9GYjZ8CfDvAPBYMRFXiZ
GKZA04i1zgsLJuN5lrR8rZ1nYlKUDeYmW2B2+oN2b2YDxGqNlMX2+cpQbO4r
ZuTLloLLs8Fnv7Jg8jyUzHpbrCRLvUBvwPDwLiPfmVQdydT7Gd3qAxvoKuKH
9kffuPME/xuwlRtOBgg3ZPcYw9fcZgiYkcNWjfvLlYVKr1kBKXa91Qax8Yat
Xk+Tzabuy0VKIoChKU/Jeo1NbAUVSOQHJ8WYhU/HvF6y13iFMSMGGhzopZq9
/q2ypyMiD8u3smh2QleNzTtVDtO2fGgC3OQrR2Tpx2bCzKQrSRJUyaT9SC4x
acrimK7N38+JwJEn8lU+ThW+gc6H9pp6ArLV6BjMmvguEHyouwVczzqgc0rI
mXler5ioKIb+PFMdyX6NIqPSvvQpjOiHFo6l2THXtdKwBaKjQVOGLYlQG2TS
6wovJqeneNpQopNcJfURBZTTMYkt7tVv/l5pV1vNNeP6QbwqNJrZMpg8wlXH
m9for6GqfdXCR4Ietow9zEeYyOgXVEwENKAUnDR/8zXZoaBl9cHO3C2jQ8RO
JNzEeg0VX6FkMphLpA1qNuxQ8VNk/an5wH1Lpe/Ft9hKHZ0g5CISLvMe51N5
64GEZQTeWGJKaEvztZLReT4Uh1lT5HCE924e8Vz9wwdMs5S6jmLjtMM/cqHM
V4ltB6Rg/1aWvJpymK6UKplIkSUKl/MeEf+4ieIyD8AJTDvx3AwFpHvqgkHm
xNxjfG6YoO6GLfiDsL11eR+NxOyXKd9uve26Z9iJmFDX8R7b9jaU3DHUl0vH
nION6xMVikctrQkn592b1WjOuYUEpN5Up7TckiHcsEC4pHwKa6n5+N3dmbdj
GfSe/PCutg3fr7xqwT4FMPGOKTVgHGquVs5Nh0ogdts1TYGCKBX4ydVFH6Pf
tGBvdU229juNMNleoDx+vz2NE9MR8LlEMltq012DDdAZAT7nD6k7HmAQdWbH
3NeMMwT7TS9PQuo28liWCoSJ2wrI/ep2h4iOWiJBuRUTpRMQfvPj6lQjmC3H
PpEgAlfbe6MbdkuwwCUHiaWw+NOV7/LVvk8e/+WQzkXIhvsMj7ELtVKQsCvX
pCq+nC5hr6GNg5MP06eqAarwZqJBP2lKuUXFE2isB5F79rLcmzy8sJPt4hAR
2nc/76QbK3Tqsu4x3wH6hZIFTsNvPUQ8sxJ0DqmfbIboUz4wEgLBLuyhgZtK
AfZ/x2gDoOIRIm+61gbrtn3q7jl55qUzIJ5xO1kGjyVCK9+6xxTtEbuVBb7B
xcgqBYycN0qoZDbyLAY5Uu1pfKNaLLkDWrz5hErcmQzqnSkX+OJ/hr0cmklW
2F/eHyk3Vd1/mw8+bhUAEIjXiHiVSy1X6lbt79JMzs8hRs9V4xgNdQ5VxGau
wuccrfWmt12XtYeGfdG8pyCeNieoQUv+IQca05IPKMWBjIzHJF8IOb0jjZpP
LCL06EBaPjApgcf0fiLBRh6LGMmODT0WrLcqgOy/zKXnVqz+kwo3E+wMTPrx
f8y1dDg3ngvwCzY7SFxbM4hD0KC+nJ1yvY6daQBpfARjZ96l4WJ15BHVhR3C
e62zxPFBr1llH239QqJD2V5sKRv8e/jrAGfuxmQcgrCZ+wrZja+ew3W0o3FA
MchWsqUpbAb9idcvEP2d/8qTIVu5rI+NNyfr3HXeWGEL+Z0YHJ98OepaKjBm
mzHe9CpL3yryQFVDqMihthP1KLyu8GfZF81u/rEzOYQh21hmYVS1FoZc7itn
n3bPSziVkF5wzh25aqLBKXQHxebTcg+H926wB3TcnJpzU8HsQtkpmlqfplDY
MwzlknSLQfbD2FH1C6mfUoWFLpEzGBfhjZqDXLLNqZUNOXFExcBI7/N8lZ60
qUBOT+JV2yJOUWdVv1Vxobsu+F83o6z5Sj2gGZNHWVa1hjz56+wtze5HJB9B
GsIDqVxT8oUuf3Wgy8b3k9dvGmtnYvtNbkj48wdXhA4S6xFmCxKp6pKdRAHI
ra0Js94RcGXgjrubu6YS25daKCpyKk43EZbQEmKAnp1ppspxQhaoa3ykjtQ+
LwbOnEJtxqlK5Qv3mb1AqjNDRQmmcu11vzB2OrzrZg4frB7tngzpkiuTtRbC
7xSqq0jVreoOhvuHiTjWMgKCPRdnKEQZ3i4+HyKRCuoRp5kaf50Zt63/ahPD
zxV49qegsNxC6GFYhE8ZSA1Rnk3+3sjuG05bb28Ii/h0Xac5BT0Jw3EF1gTc
ewrvc2sk6bAjJk7elpAhOD0sPP7erOPial1iG1sePwE3s98vdlk/I2FCJjPr
5GbRH7Ru+qkiF7W6W/N66Ja6jF6W9dY1fg6Ts3WCOU59UxdvkUmnlU2AK+uZ
6xHLGG4Y6AnLfk9bY04vlHWeJO3neXezkzg4tiBK+LT27D6h0lHeZJjw98Gp
q/OMffC4IU17W0pj39eWed2EssxTX4WXz7uIffMSa25+ELeBicinkIzTQ2dp
vxWoNrSlBn7eBHVOXJzYMzPqRP926CLoCkvIgbA0y6cT+sHpIva4luFyon+B
/0Pcdjm1JW38iZO6itLRtSOGINMwgMEKQblr3UFwWIy404bARyeigqrY/FgV
mPAi90HFG9sGxERtC2i+zU+izjOGM2BbyPyI8GCOCw9EAV9byrG3SD5zLp0m
XOHO4w6S7LWqs+8BbztMWQMjoBB4JnWngO+ye/beF0KAch0s7xK9LB4KG9nl
Zzaf8VyJdF1VWRUjnbAKtvU7raH5XPf4ofo9mARE/QxW3ZeIyHmHIqDCXF9t
Nn9pseSe7EgTblFfsdF7X9p7ezpErPKuAOTWMTdDz0qbsBBapjEChWk/mbST
wsj6xa/0dcjKC+x0+y+uxJ2GZ7LWB/3pa6Dh7LJeWp1Yo6cnK1v8wC3FpTXe
IET4BnEYmetfcuLGAyUFN9y3ugKNG/gxD53NSjxjdFIutuIxTM/dgHXSCE01
8oCoFaiZvQ5piET66KDTVYV85cZy8FF2KjaWFnU9xftyILTeDBLC+K4xzcn8
puHOo/rPAYl//94isIXZHi1ubmM5ddHOdcayJb/HPQols5wIFD4Au22yIZdP
LrvmZiH3o1EM8gp0K5PrVwmiDD015fYXDaJMJRMJgP/OVFs3fMtNtipZzLtL
s9jgm1i8C3tYsFFAgJjMKLzbeSFCvjKlFyjnLziyXpEtoLoWgA84Cd7aA1Iy
l4anUr34AkwiwOcc3u23IKB4Poz+qoMAxWRFEn0nhug3pZud+hdUXt3AQ0js
zISKAuRha9HKLaxA+5w9ZTT/fzQtTdiRfTj/QzAJRc+WZcFXVni2ovLoTzQr
smPZbxul9M+1GaOb7HfVxpQMaNB4Co5JROlrqMMNYFKO6JTmTOHh+pMGPdEc
NPNIe2h9A8M0iGswEbii3fTlP7U6v5b74DaUJGhj48lFQEs7lhGutkJqwp8Z
cz2M6GmtiXeyVNZ4GakqSUyBkCQkMjvMKLaGv+FpXTfnsdEHbC7ahScoYswZ
z4jU9gHg/SN7qViYW0/qnlBrcOdkLZkrfFv2zhoSsW+il/fOixX8O/2F4b0C
StdoVSGFYg8k3zUYw/36FYcK798Ss5fin28Kj8pLY9llf9DCWOazXMR9vOoR
oie9iWYCAlUoK4gWgPsrl96iIckEyyqNtxm94x6QWS51P8Oj7Dt2ZSmAmrSh
m7o2I/laPnJzyClFQlCamT1WF5QJVtaiXvzv8mxzzOLB4ukaSLMPGtVEtiQg
txPmwqcmBqnO/X16r87t0uwUcx+ddjDH7jYa6FR+4YCPKHz4Qe1gxvZnn6Ph
/4NM8zS8S1iBnkoZy6XNrLRkHdttaCHUvuLNeEFcuZWUWBbEQqYzt4E1ncDf
7F/OjarLKq1JcF30zGj2rEf/myTzgoDfe5NUpIpkXDFRnRJizgKsiPEn/nSY
6OlYeAbsEO/n8e/A/4wy5g3NilvoYzKZrKxsPdWiIjHMbl0JNnDVtXA2hLHI
W3uV+n8OAzAJZsEgTClnyzFXkNr0lEM01yZDnLDw+wiyf9eVJELgScw6P5gx
UuMihZXH5tHI6GIb6J/o4f81po4farKYwBT3aEw/eOk9tW7bCnCJgAogXHgc
CjfI13/GyZBZcblqh5avUdHYQe1B8rWTFJQlF9vzkpl8UFQ3HaZqd1YLBsSU
ZrXQ9jdHd4vmRDWaAICeVjtXecSVnb1NUV69oVxMYZh5dGyFCyD8yadlcgI5
j7Sf2zzb5LZQF7hnAhebW/5umla3/nYWkb2g6wB0A6QNyDI54uopifcf5oda
fp87o3pRZJpPZ3Hsvr6jTrRTfciLW5vs0n+DJToG7VvOmds2/KLguDwqzAmG
pVvwRNcdLt+QR+cTgRNTNbzDuo15wNuW5RUVP5fEaBHdfyLMypcaOczcWZOm
fl0tU3owdJWVd5gnx6kkKyiZjQfsG8bxFcgqfhG6S/KwOUs9U1uMBFhKTs6I
CWdkVZk3KPDrpNNWp4hcV0gzz6vUzgWee4LnUMUAIGgnFPOpPMeHkAZOKcQt
R3XzHhrvQaEyCxNorklEIGdlQ1C4oTFbTKiZK245NWWd1L995az1wxrWnVRR
ysLpQd5N2TuJKeBdXaEgZqiJWL8/rQWNK5fkkCLGUSv2Uhz3eHN9Y5P1rWTr
K5+Hhe0pTSZTzOz8HOZ+cUWBn3GegBu3jpR1B66EBcziffEFLuG0gWmVTJwC
9s5TVIX+gKW1jpkE7OlG+XRzHITyblasZL4ueGDnqnn05kSQERu25iy3X4pj
kBvTBlfRWMavnXNi5FVTxP4kjrEpOqRdIMCReHZCCf2MCNpm+OaeH6OMl1bQ
8zPKGxK8gGpHrG0Fg6CRTbAOoWo/ptRXbDt0Za9T5jgYBEyJKsSqbK2aDzvB
mgizl0PGRAqJsSqFOa1B9ZP1f3c2oRXc5CTsCQLwIgQ+5+gvcypF2iBGW0gC
9kUwVe1GkESvBL2AILU7akreiio7U9o31XsmPQ5e0y+S0Tut1z3vhFJiVgRl
8Ep+IST1eBtpDzonNyyu9o0FxpjMt48qvprZ9jgTRuha8Z4BE8b1Am8Eu7Fs
F1VdPcshaqU661sN688ryoDAmImOvtMTyGuWrJene6PJsOktKAAGlOJFNBGr
PZL7R1yRd4VvR3rkImYu0VjUsRpA5qkqRZ+sq2oxeI+H+mSYAI/125m2xxN8
/WZjg81jzZfSbI3BYoHn9fQvKPfIDzsMJ3secETHhUkLitbUNJFVpLn9xiLe
RNA4G7UXygqHCRhqi7FMJPfK8WXAZe8gi0dzR1HMRucM2YCm42vHT4WtGRAL
lZ1pMqPDvoMhDRfoTX2u7YDJL8Z/1FSdmhs3dIFKhBSbglthyoGB5qWvqp2r
qk8DbVRvKszfKW3vo2lF735+jA4ERevIeyEn1OA8SwEDlKBrEZKKVZLFmEwx
YUmTRNTznqieQpA3LL5Hzzqo1o4CzPyx3uJutlkEPuaVWuVYUx3rM5yu4Cw9
FqcjOhAAu5ZzQCOigk0F6yFzHX410ttAc+ZuKEyetsF8ckRVWexYtjLgg+MB
ES1DpQG6y4lmNAGx/r18HbF2I6aSB7d9pKdewP0fZfyyz7OUsUn0kREGbcWq
r5CWpAZC1nmfUSIaBzAHKD/iMI72m9RLNyfHE5BOj9fYBi/ZMgtHb8ydc/I9
EAX5GXxF2zPorITJiDJiWDD2zS/MmryEQwuiNO2VKMaZihiCih3eaBZFeFnH
feKnb/WGPcOHiCVmcTYa4BAWGSRWEB8Lv2CTE+MNR7GZQULYkYPWurT/CTrY
c1P4u/NE1MF6eClWAW9c92Cj3WTrlWv6kkHwKSFDIWeUX52cP4azzZCHJyQm
Pp7ASxksZdYEiecJRXBu+aenQjKWxPB772gdCmd9pAu4Xkxb3rcv2fllQlyM
SHH5bCCdkWKaDs72LVQPuxzqeEsVhbhLeTmerTrNkVpSPLlf1M5cYkSb7cmP
1kyuW8+3OXGBmH2p7e/tO1prvgymdTWtvNBIjhSbcrViS1Fcec4h+3atsEBx
Ce2U3s5cYCyhyBNnfylTCrUpS8mF0WbJn3I+RZD3KQOFSYDKD94jnZV6eFt1
ywJMi4pOSkx4l5KJzwUZDvI1EQ++FhOJdgrLE0hRyDH8SIex8NNi/ObqU105
MRTDjNsUfrroB6uuS5NPZEtm1GRkyB1OnS/DMXB99bo2E1yl65qUpCZXjyG6
qYjiZqC/NB6DEI7izfl8jj7ZjH215QC0hpse4X860paAa0WC0WbwuKS0uKV7
NX5f8XyHCDffJZA67+ffY2gpFK+lobu1JW++AsQgXwRAGUg+EcwzDrG7xI/w
jhArARgAs9xyZOyZjUTV6bWD0FC4c9CMkij1Zt0ZW7Oyu2MJbWHizle1s7Vr
kEAU6vEq6q8LgsfVshEVaNS9VfoTWJM7lFwYuYnpcaG383SM+q6AnVy22Fp9
ZyejGd5MTGjxtc0KQfnbeaE1r8TJ9QkMVLzmM1q1ojZu9IeIpQw3p1v3Aq4x
sEZR0+5iGHBsCryzIjKokWmVYImRcG3b4XGu9NyW0X4UXU/3tyhcyxwZzznp
5hSeFP+VHqLSw/uSeUPJQDjsZIqvGcN9OPVcdoxEvyo6TTtEwJoVsxPhR/Co
gIqS+sVvtw0fZP3jJU39BDpCSsZoEqRehnEdZT1ko6PiKKJFVdKpvFLgJhP4
GZX5DuoALPtfXFpHF0rFM/sEFZDoz4nXEJoutObbjHIUzqMBbTjeRSiPr/EF
Lnt8uG5siYiaxX65ECmRnfBkHg78y5xJf0/n1liOPeuUaD4HrJwkZ2dQDZgd
Nol1HNtMNHRfUHaUzrMW3vgW62u5iPmylEvaIVmjRCEbGJrO6ydvYha1+O03
I+u5sua+tPesUqJQXhoqxNanIbteo7CRlb2qEOy96ckQEl1wJ/idI+f/DA9b
psO2bgFR08fgZgS7u1jyk3Q3+lw3sZdyJhlc9tebHwUVoi/nHBL8GbMVKAND
ESwYkJ6voA7MErtZQP1F6EskaMDUZMdnjpazb9YBIGHzJgN6lSRUMAe6zhp4
3kq3X0u5m3UFjFfTziBaq599QQ5Y/j3QXeKsPR+4t07/ot6kR7WfIYxkF1wv
d6IJ9jHxzE+ObmXHiQ5qa2r2bgb+SKj1X4e6IpXC8sWhD+x55Uw9sg0e1SX3
4/JD2hqQ75dGxXPBp0iHPo9XYDb5tNvKMatviiwc3kTkug7MeNz1AVu8V/H6
C8TV0aeyjVQp1dBFq++jlPfdC+iVMZvBMuDH59NUrUg7PMO5FJ3VTeyG+XS3
0dePsIFUYRdT9etjV6Zrj57AHJfAseuN/Xai58irAkxeeSRL6PgyWHX+2FMn
ivUl90w79VEwd1rkkaLZMupZt4/W6oXInDiagUVA7mYLq8ynEn7g+gZxO/SW
WDLrahP++DdD2KQ1ruRdhg7RvGSvSZY91H7BeLFLnRH9a4QTaz2ChBl+Rm8r
kYEMN6is8UPTlAWdRIhLAAOIXzdK31Y8bPQTH60FmFfUy5lZKzJYob0aYS1J
uTq4dmw1WtZD9y5WHl+g+Qq1DZTsywnfhaTzhcf0NKq9YimaNDPmcYS5Y3kv
0qnnIesEb84mRRK+fjVn62RoRQu5+TqZa9snfXIjw6CSYSo5BpZXMxcyAjVp
m0cM7e4vnXhH8WI0LEJAXwq7yWvngSJz1VRulI6urGrnIyD7mkkIvasN6fo2
rXPD9AhhDaghqTlSqMrRLoJIVhcSvzaQnlWRKFe1l3lZ6LCsOzTvwjjE5HH5
n47oIX2DlLhxWe391WYwomj1rVRGLFAe0ArKHw3YNrt8QIX28uWLKRjq+iLB
j4D6mWm8KS+TVd7c8MuzqyTkzntJfhRJkOq2x+basKKLxG+h4H/9pvMm/WVR
EShwEifjp39HcePJCJTkfN0FjtI9qp/ENCEMpWuPIH5gJGcWxgn8ctU/uyJQ
prMp1Ts/8cJSXztLz/lCsB0x58hlepw6ApzrEDS7k/FpN7jSlsegPP6mL9Nh
VTRoRaoB/G0mhLaid9l6eONOPEOqWBohnC/Vkx9t48XBW2MBJDR6boL3Fze9
X55aLJdFzSTSmzG+3NKdcs4B6Il9Jpq5nbIUqy9BYNQo6i3XvX41UifYrdRW
cBuImu/Qt/2tAHTkD/fcMirGVTlMukq70+CaRd4BifemnsQqaSpsc2aEstv+
B7zVKJcNZ0R5Rth1G65RPdsb+9ZVENZK59Sp8KdS05PJ0Td/PKqhfrMMsrpa
YUBdrxqflZ4zDqiITKHBF4b/MApSel3LILA2NRbyBGFd2PysRl0CISyirDB8
8pC79DRAem8h+qqQXOx5MCbSCh654E0esouHB5nczqjC3iZH0LlYzOV6fnGF
zwQRQBimzHCkTBKFZeJmIQpQc+O96RjpS4NH+9tJklXD5gaUdzG1TpoHtbkJ
2ybSwZS4FrqQg2NgyKFzReFvdi5ltOSzbADLpst2fmJd3U2LI85YVcYDMUcv
kh4yIIzrV3v2t3xbQnRy3YvenR/XFSKGTmHzqgpmu56jXWuIzU7bDfqEL2z/
S7FyNR3tbdtcoNjltQ//MqAObENO+TmWOPwg/bNuwlHiswfnZHtVEeUzfP9j
+dKPAapUZU+P3pZzTHc79gnlMhit5K2lWqkAxuqi9Dr0DYKke8p7QdXILHo9
sywb6dkNkLBAdmpOPjILOJqIXfSbLTQ6iBcw1k1icyZE0FKnsYPmWVIxgoYS
rqKp/MeClPkw8O3YO0XQJ81edGZ8NMRmQMh+COAKfhcbqvMDEM+S//WlvfKg
FrwON5c2pJVi9b8z5Noe0ImRlghNrV9jZpFLMhc9t0sErDrped8eYgSDSXnz
G8uofxQ9Z54seNcW2O2aMXPZu2abZA7zxweVAXhe+EPnR0Hq3lwzKS+bkWmn
76JUFmCOiwNKM99cVFsJ2ZXNiqysCRVg0e1KrZIjsVDAc5w9JeQBR6xy3Wgv
VOx0HZygnEH5exswWZ8ZC2ND+Av46/3Lzmj/zo0IPUPqfhoe9I2gTxG7e6G/
62U8Qh6Mo2a9ozbI0L6JbjDWGyohQalfhQEfrOO/DoBmPerrnP9MlrmPA7qt
ORw+6eDjVUqfifKLX8gKIrkvh9VFkBX1nGRLucPfW94GwA9K+ibJS8DU808r
iq5UbffoLi0J1oBWYnZdZAnMHgir6AiAxJLYmvH2OOAUIVpGimrGC7hBHzs6
84TTfY7kR/T7Q4+q8wlmlAbdWSLqPlGPpdXutfXyY3mwPQMtl5H6Ei4Fg7yg
YFxsR8z+AiHyTGYGT+6REsFJpyxVrgcRU46q4YB7ro/gRp+iGu9cltO69fQR
uWv2AWRLuJWn5wkIHKwFv1ukhFKvRMlsjLzkOMcYHTlr0r6eFO0NCODHR0cx
Z6dJBTOF7PfDS/jLboj9DcJjhl08svRLY1M5pzpV89bcLjskl6wxYHHj9X+w
kNasxWPSGzttOjK3QPZiS08mSHlJl2tLej8J40j/9RzroBwL6zQBkstp4hMb
9DUDtTto/ahN6q7DBdUJMI4oAFt5/8SsDYGaEqW/2a+G49RIA7vLvIVx/kId
BOwt716NZ1FGY96HQv1CUQVY5BM5G0ySGFnvKul7qGEI7AOeJu2jbdaVXJNy
kX9NbeX2fyN0to52ro4rXahXFMeZZsZgfDGYGkHjuVf9zgXFvxX5+Ny+4w4d
SyvSZnuYfFJ+U1+nX4k+4l/V23MLV3gWMo2TgEUN990KWVjRQpOtAL+J+IXz
zjXbTH+bwqDZc8sksZ+cRqPSUoRISnPhhFYueebivuE7mSIga8um6BjBolbX
slSIX3ysgvZxCNLytQTQicYm5f2a6zE8nQiQM8jRhzDDdcKRc8B+NruTw2sj
9eypwfYVC9gGlBNionLwrzxuuCu8jzQFNz1aromtxuirf93khzL/TaPu6Z6x
gVZDHpc40iJevTmgRaTreOwdhwvPYBNDZkX3fGWqJmFbFtNJ5+mtfoESBXjY
jEDoy1OxL6gIm5grXCifda3WbDdgXVaFt+43RalzT2EkIdHuypfm1zYAziLA
T4/TC01QAZfjqNHKgt7n7g2vjGBi9mZ4d/Ot9+r0XALdfe5k6VMR0ycsay57
Rwx0Ip3nv/hi24T+zcHrUAVq83q2gB5UE9IkAP5IgHLRAKDuyxokYM6IPRr1
qnrqA3fS4S58SC4/uNcTKymjEEti1+wBuTpSn709pGHfD9OEniiib3TgGc6y
HmIti9T/YtM47GiWL183YtC7PfoOCmS6OZTMCgazdTVxck1TmYGLGIW4pv4e
wR1RlzcElVt7S2BlDEVqr62Ps7iA5S23x99Jd5cj+LksAsf+CmdK2K5r3jrQ
O90GyVmgrbcdLPaXILUdLfsHX+N49dS8L5QqGqvz3LSm1vmtleeNK43QRoEs
hGKvg6PgyN9vXgCVxnBCuztByV6MjkAJPSdm65UyycyLaIfxNuPbFzZfkDXH
zkw+OCwjxbxFZ/7MR8ATjWz73j/E63/8tuJ+Z64sn5bv5t8whYr5tnfIUhRg
2QYtwKX/ed6lRepBR0XMK8qZxw8UbVWy4zeNu05P89HBPSRTZ04KKcVth0xk
z7Bfor5A5AsDVaNe9B6LPeaUkWoj7FwRBdCToG7LhVT6ZYXKZFlt2e7266LJ
H+HTVNDFLz5iBGNht9iYMXkEHBoyzCLrHh6oqXlliorzWQAmy8obcdUEmrM3
Sjdkc8n5vU9/RTx5FQfOqsmiQpxcgpqaJCCyN/9SNU9DGMb8jFC6+wPi19Co
bwRdSKW3I/ZeRB2SCHwGPb/Whmuc7N2nfiV7uiOI6EnRZzRgVbdQqAghpIUQ
SI5teNMXU8Hx1HWMmSVdu7gdUCpedWCQtwGkZ8XRCVGwJlqPdhQ96czIeAzA
pOAEkH0PW4fGIStzwoNYnU1lHExRl5glze+uW9ORDSyTVgkWv+JxnNcP7/+R
DncAKLIPB/IDUWJRpW9x3KApKYWnIx1snsypunFgjAD5CmRLOym3itI6wM7i
aaD3cBxdjTRii72UZ76gQzzeYheVcDwWva77w+hczcecJGvDbu2mkX8RHenH
1Y5Jp0GCfqt7UVoB2+av14Sar6FgLHy0TGDb9SbwJusbihwIfnSFaHuJ8GSE
CBo+m7jLfN0vxgiD8h3laznWQVL1X/CiegN1ijuBGYQMGEHJ22FEXNfnx6iM
u/Hm1h0Qf03zgNBLmRIl/dlr0MIkYdKXs4QSsZ9k01pi5Syr/Ja1Qs+y335g
cDx/YBiSrrudIGi1OmUwfdk3wffL1+xiZlgeb2+n7YKjiiAgcvUs8K9FjbZk
lHrgfoAwyJZ7cZrfAxiL5lqqzI+6CI88RA3Z7JYvMdJgJk7mNH9m2rnNH/nL
BqUwYJy7nDZHQJKa0N+RA6by7e5RSx5h2zU8aWEJG0P0GIrK4YtBQu9yPRO7
VVzKj3xe7GCWfG7mEwSp7qWHEO83rAalubjHPsW8Crp4RQsDC0WaF+uewEc1
drQTLcjBMKm21ANP4FhhTPeZVfnvh3veunEBQaBWhbCBZSBbz2REFk3/mFZ+
NZNE1DhHNx8SU7uEE3bMFOE+odwnVSdgXd/nH+PlKR+zrxFi2oQDLfJNQcEr
G2It19XZYS0J2xxS4i4Rc8NFHIuQjpTzi1Rbz8Sp88HhFOTe8Ihah3Gmfjmi
Ur7Dq7+fkE64g0gUTlsLx1CjqE1dHssnmMU9FhtjBqRvYrZf4R8dtD1P5PRH
OzEElg3x8fbq546/1uqTkAh4r7GEQVV0u4h0xifD2evpGrW3unq/qa+aytw8
c8ofjMvVlTXbNLMINROYUKtbaNPkOO93q23ZDWFmw2TTQBe3szlqFpn95s2y
0ABcynCmrdI3kP6vfNFWe996Y49evhNiUqSG1TUsFSF8A5iBCQhRN+f6sEqQ
jtg6D9mxC8OHJKPLgL/chUQdOcdaOyI85xTR2AfZSV6lJFmWjg7ySIJFpfW4
NnvJ+JnrpdcnYvlr4uPNqlHlzgSt6OIwoK5rncS5JhEMW1Z6bdDg86BL7Dfv
KU8SeS2qHkNq50hmTUPxyc2LSdRvPnWyyq0L8a/DnEUGyFr8FPKTult1s0I/
ZM+KM/CxBgE2icklsipt986uX/Cex2ij/SwXyU2R05tSdxrHXraoqlaTcN/w
cJTZCAf0buqhgbpSinWsuxHCIeYF+z5rugRFycOqwJ5f2ExBca4rt9DJjyeG
S92zdbAzg4Opko4hx6U+kjCC77bDIEg9n+s8NeM3y0yz84hS9zyCT7dVluAT
kTHRKsImSRESk6dbhACUj38FwQL5DmUv61WwvHrEk4MUBu4/EKXw8kcy9zn7
2ixmZtXLUdj84uEoHFDmVGYxHGReZR3UgH6CiJWF2DUMI/gbZxNUYkq1Cv8k
4fmoi3PZzT/7F+RM1ICkGS6+GRptc4dMrY4s3OmtFFg3LI+pAbsuVX6MG4A7
eJ0weIs5EtyUm50QRmx06jm9Fm0AX5V6ha17Xw7NilgE8kuhuww4PBinFpvh
8aIy/LO9RHs+txErRGyAm+E52v/v4qkcLwiVpn2HGA6M4iR8pDmBByig+EQj
i88lKS2EpUvp9nl6QISce7oFzaaz2WIXu2asnWlNIWMStR08FGTv2vT8vMiG
snVDRTPLgP30sw0RgOF7ijh8XXLXpe4yc7WLitmBFzoSP357ZzS8zG51K6sk
ohEu0VfVehACLzEocVFJVved/J0wnexCqEE5XoSxhI6nomqdgIJcCz/Nhwlc
UV4JkvL1f59gAM8/jgZYefEG5IBdwAhP5NJ4i5j8zhMXfe2qUjt9HGEx6FJj
0xdtTwBdK23p+4nVd8kjqp2TfNlcKarkwwdcEbzXFVmqTMtSDJc/CZRulF88
jHHfTUSMvnkJLhQgyKRDpAo69hZrvaA4MkFNvPoZnIGXvXQtheNhivn59P4v
pFKT96kP9y91aHWgzyBqJKTUMFvIwaizo230tyHmq3ZeucU9FuKdimCGCoRf
QcAqVgyvt0UUmVWQEWKUPJTij/fPKLkVerKJSHPkP5B820ilGyEKdc27M2tT
pyX5yKkbhBel1HESVoCn4UyDRBGne21cQpbf/swXSIOedQzdSHT4NTAK3anw
Pm/KE6bn3b5O1AmGsDwOvc92za+JxbNly/+IB6KiWS6uQCUFm8IeYiF8SDCe
I4y39ZprLJv4eHUNSrekk7IFJxDkiVmfjfK8RFD0ALlZJV5V4MDejOzED3yV
9Osbf7qCrys4gwovP7Ckpl2zxCG3HOttX001Z+Ch9+099Ezyz7yo7oxGYefp
EXieAz1n9Ud2aI8NYvVLUVyYMaoNewexkc3r0G5lq24IjcLq52FdPCChHUXd
/pmaQ9jYguqbAobx8R3TMVfZ/RqcHbF7xxgQrYdfnfu2qUKlCwCpjsQqQ+9K
f7xUWfjJmELAdm5Y3eHvCkTFrKPz7yWrIYAFFrrdtoBW39AI6MzFgIlPFenx
u+OGpj+BjNIfM8WhF7CSyCG4LSNMMMnwvWEfqerK3jsEhWcubqwYMwrWY/9g
1pdvcmIkuDpbBm6P21V4NzZa8pzQgYHrQu1HaWtehcmp5GTKSy3VES3oRA/J
d7ybjcKENLjYUkyYRygIuBMESLMBvKAnp7syiciqiT9yXI5GkG2Oq3JqeHQH
bI3v+3bwkNCIMOvaT6JftVjjLz7xH9bpYn0gDzN9NR+vtraNm079i4k9yiRC
nqeeUnY5Fxa0VI5z/vIWCKjoOmpXn3dvza83hBHv+IB4h9tB6pZR2SVAo/dr
49LadrEb9hEVykLbVfTHSejFqGq8yxBt3RPF7BQJCX98PSyVHxq19lM3F6WN
SjGipcmvkdrcCBU2RxAbyAb1nKZzIaymqwFgY3LGbrVNIkYxlQrZ6FLmA8ET
u1DhuSMwNKzLf39X6NV1kH5sF2Lf40dxpe6MSCOvw9auf5JdcfyVbgHP/866
dDd+I43vhUAIFMvzeP9XC2UD4tLTOp3s0baUeajo/V61J4tohL1PDL0a3tMP
DhDBbNhJadkRmcW3MWAOLy/5tSATkgaDI/uG65ig8uvUSDUsYdaRJ1SKyu7u
w5V187AJRoaxTQDB6dK4ww11cdjlti4QNIsXWfyLwCKXVGs766Mg1wEx6vPy
91BsdZAiRuJjQLSiaLsN91YzHKPZyhi11Pp/X1Pzb2nUdObq/OSl2HBjaniS
O7MUTzaqW9G0OqT4dBMzEkpwJlYEbgIVtk6+dbumcYcSZzGMyCmDDYDg0s5u
W50zvmIvO0wo1S56P5VWB67hbVjodVXTI7Feb78PAqykxxxq5ox97XvonFNi
vdBMqzdJIbv8zgtBzSTXVkr1NmfJSLgyx4rxr19DglwkeEg5x4CINg3rnRCf
JDr9lRlqk5o6Flh44s4MxyUpFtjmQyVaX1oIogsj5ZAM2z0v5glWZ37iDcF4
2lEVxshqzUZjkGgI6bEhpNxaDd7oeitHvJ3iQnBJ+r+7ZZY6LGZCec5PazGp
jleOsycCBJ9NM06RZRhH9yQnUUCeNLwdzt9jpXxi68OqPTI0IFh0xMTsMKdn
dnisPSRmHZfs3Plb/cyfzcAERcX07xhZ7H9a4yFhuNQGNqMI28W9JGWGlLk2
4cA0vjizlTJzzBpoKAQQRBE7AUJRnOeybCZ2vB4D1X5PpaltUyFXEkFuupQG
FACq0O0SFnuR7hTHEfxiC0FPComUdxtsHPcANdWbJNcFiFlRo4BY0wxOajDU
5KO1Ew5U+IvXjYtyU1Au+MmZOX4gDiJA2x6Wf0QzJOVzifHvNSSuuzeNHPS3
gBCF6+KY+AgwzTIY1XdDCZ8Uni2QhRS1+Vr7FLELjO2bgGnh4IJDm37EPEAU
ysmfJDUjcqEBCww9V/POYfsWWahvELMe6o98FuEHUZJM5bVWsK5/NRuWGI2u
xSKgYS17Lr+bIQnr0cFdTBH7maf43JEYmo8SKshSQviNgowtzMNj4+Fhevj2
p+BWmP23prS7xpATgJnrJJtu28TvyRunYQfe4ybnTjd0EykR7G+zMcb/WB6z
lKKGXe9/VB8H7CnpXD/E6xDUJMGp0/zBy8wm4o0UIpqecboOQRkh2nj0QEu7
LhfLg0XdxHXISNE7k57Ph3WJWuGhe+YlUEoPDd+ffOEHpo2S3Jc3lhV7/jNN
q17sJ31HKyEM5dRx8C1rP/+2gQnnZuf/cqtFKr8BbyxTyM7NPDDQCg5J7hcU
3srsIYtMeYw1bs7dGVNbFFAX0zqiGXxWIBVGAhuXMSa5zkgvlDq8e/DWHyGU
HTMlwx22q+u0bAXF1uqRjHmSdlITC+MEh3UvDomYp6LT9Nwx6GrnEOrGOgOI
NvOn11OXz7qKZcVno1vrtRO/1z8Fd4BRNazDRMnLQQzPiQHkEzNhVt0KapUi
GgMsI5Zvy6Bio3Brlcsg14Slh28MZQBrmhDupMoSYMu5sjLhVppn350xsLv3
DAO7b7IydmEXYQ0r3PBi4ab/KWRVMv9Gd3Y3MS6E7wb62wQjQ5lhb6yRuqS0
8i2rkhJd+uu+wwnUGeVWvkFtSWL3QyYjZf+elFG2fpqUm6U4ti2bNLNODIOd
KGWCAGwYZAYnny9a+TnpyoBe+U1HC+tsHSGqaV8g2se+sMJFbC+VocqkUYVh
ZPwAZ2ZdkNpukEwJYoBmzrH9wfjBZBiV+5OO1Fp7k//13LkKyngRKQnTceSY
34TMdvcHy/owehcc9aNP/snFSU/N3z7AIWvlhXokPFhcRUsR1FYL+R7rLC1T
FkWBxJEffzSU8WVC660d+iUuo4uNNZPGBDjzB3CpLhx6ukaosPyA/0rTmiT3
YmfTK9DXd42xXtqYdIyI+6lH4rh56EeNBP7akMTI5Y/oac0Prho6GnNnadqG
Ra0PIxzIW3oHofGd7UGSIMQs4Z2Nnji7e0DFFCbDYk6iQ4XRzsmc5yiTDkFg
h4SPMGRZaJS/soVaO77CA3EvHM45+Tl45RT1cv3QJzFzNOgD3vEv7WZSO0+A
5UQUZ8ZLyrNrDJc8uRsiwg+O6nQFrEy/86P47B/VLu49ElLulgfpOUF1g4Jm
SN6wE3LwdNDiAtr5xb62diSHO50WprGlWzO9V61zQNLKEtQIfItCF6uPlFeu
2NGOJD4wwMAUx9rkzjdloEelQMXeXvJl9Hn9tMnSUO2+Emb+JAqwdMa2T/iU
3xaMxclTECKThasq3K5GGp4fD6wqGTdnlMoR6djOYq8rOUEjzQS5LDhMQl2N
HR7IiECP8jN8tOynLwA2LbFe7p8ejHTCngvlJ2HxqIRpOt17dU6/CzFJBKzh
OHuIcNUnPksLq3IOqgL8iQUXYU+TFlOqQfSnAO/yHBGYJA7B2KCCw1bezU2P
po3TEQ+ABl7sU58/9qC53pDjNC498ONtDwwydySs/51JuRf4YMxTc307fxo7
nYy73m3X6KdA8UhDDfyL/KC+33xLZFPedR2WKgg50pANEmOQ+Rxotmm+XOt9
OWCp0jSDwqRi8CmA6jaYJqObHMx2qRohWBg+B9A9ivS4+wq8+M0v9yYX3Xm5
dlPy1s7CX89BSAAD1PtBlJwGZt++z1W5OA95xNcOmCcM96pR8Kw2pWP8snaI
+ixCqFpMp4FhCXOKLAyK8ExANBbdtUn29cBiABYL+2DmGsHgiGYJoVMbSjOm
Oh1u4E0RvbaYJXlwZY13aIRNVJsGZlTGbcqGyb0cK+yRKsOl52HMCoIJVA5i
oTBJMR6IKRde4y6/FuYjIyV3NWWjwpeGiC+mOF7CRuhxM2r6JfTqH4MGqbkZ
8jHCYod/jmqJnmrV5IEy1jP0JCQcXi1dEKk7gXD8ss3b7kH/sFfQxtDNFhnK
1UZcn98A0GSrxrMbQmYjJxsH6pvMbv9tTQhr6Bzs2smOEYcyfoPfEJEAOKAh
edNJ+i+kceCeiDQikhtS4yKYOmwguwwCVzetWQdypuv+5aTaimqoIXvRs86F
MnP6uiCzZZKbL2l/B/lUS46UuEX9cpzIx/+WBT7OV+ILRVM/Q1U0fFWVTukq
5cUIBfE3s6BInNh8lX8WFmhOyr8HTTAaG1jQTDos0wJzLJpN71zRCAo33xEl
Ylo27wK5xceQZvovWO1sbCCd7knvIJ50H89kRZ1IDPZ/jow0hmJoiRwk6FJ+
vVp+dhydqGxSjUAIhCXQ5Pp6hszFHbQqJVRbJoeefoD0wxi5AiHJJ4pWO+VS
jjJ9AV5foWgb94DQxPjnjF6wNUJkLKL28A0hTlIubN8GF1rpV9fm0DXObnRu
rEdv56tdxytE/xXsO+uXHEU+3VEkXkDiJTW+q44JR7blAl6SSDSQNho/AKQY
NJBp76lTqKIcezxGLCOFD2G2ZwoE350lWpzq+coxD87oCpaphSLK3IgXea1X
oteMtVnedJDEbSIoVrVj/+pef7szcezEuIWHJNoLkZekTYIAPXu01GtVuZSC
ckg90wCWgUMWJuqKyKDC35ZwwaDJ+OVUxANNcCfLdFvWacW3ydWVbe/9glKR
o+6DSB8qg27WV3c7umLGlLjqUVkjYXZHDazIoMH6Jjfmo12H29qDjSNARkHv
DE+I4/2TSLOz1i5L6l0GiW4aPUue2yih4+W1bKst5nsgScl6G5dfj2AbyX6M
XqumrqKD0ropkcEaC2wbiuQEZTQo/GGeetdnoWnvPxyM8up4ZHG4VEk/u7aM
ppaVquwYbX5m2WjB+jAahs95uE0oY0Bg0sHpIMV1ul4AlKdANQqIflQSB9BM
6R2oYJIbIx7NF+z9AFT5NsZup1KEO/6tzX/Ls8zBEicEI3B6yklRSKTvifhf
qVkezSyX1xrOrzUs36YOb5w3mVTnCAwR+vFl2dI1VnwWpZIWc3wLy22E/BQp
COEVzESluuM2J8Xt+auD9D6S6npjspFw2PnA0lWVMc6SwAJPywiIdOJTZolC
VBhogL8qQ32VP7CU2jWiK05QwRxK6TYOo/I+Xl4oE+P8A7k5ZHlvSYFQaC+b
ZYZKl/iF7sD5OeX/cQVSqR0l/76BP0iwEzoTtR8zwJ5/xmS0AC3mTcMvHlsD
DNfK7QsSWRh+gsIn14NbX/vKSD7FQuGxFUhxQ68C3nNxne1kT6N8tmEmxoTi
YxwxzLB64hLx0WrEhrlhvun5xfRDzJczXA0bW5U6R1FhklUhMjWWaX5QcFG+
Y1GfMRUyZWw+Jg8HSNfM7OhznkerReLRTQEwREiewM7vbZVGz0RFhUAvLL+H
kHKNyXt+kUMDAuGB0nLIw26Auwlv/LT2txeStPyLh/DtnQ1asxGb47OEklwW
ABJ3+p7ibwJpXoU35nNIA9/IuhMTirT9T7mm/pnVPWN0+vMkuQcMUt/pvhSK
M44wkhLwXNwHtn3my3SqJp3SHvBP8HRU4Uymi2xfNEFn5qAKA4HJTkzZqJIw
fzhAgU4fgOmRwOQpard/g5ES5kTGGgNkdY8PjPk+0FS8+uy+bwtucH+DXWBp
AU+sgJo0x0+VVJ+Xf+LlRW0bNlgcMdYD7q+mCsUtpP8E1Zn2WRIWI4Fil6z1
ThQFgmzH8z9Lzw6iFjHNJfb/PuZTr63BQomMNBRHYKIWMGyuGelM7pJidSxl
r6ew+BKhXxYYSc/vc8mx7w4lO1FGkRayK7aQmQpZxWVBtNzQwROmqGNAdR1Z
k17ikAEisyWMRKKHe2OlZ9xIVnP5usygOW58zZfEu+XFnHV1km6rn8kReXor
ACpngMjduhrBAC3ydNbUdlByquIZh1xpXrjJF3F4RPxk9sFa64q7mDuXrOgB
elksPRni4vWQTRTakn/3ahsLlM/ek9dqcTgDNxNwP5cARjoNArLUST1sIbzP
5bnGbhgNG26dqUXQ7vgFXsEqZuUeUvS1wFJjU6p25EiNVEkbu4U4hqNEyEjR
sjPhF1iWVt/U37cYEXfKam/sTV4OD7JMzHBMDayM9yAcE20nQf+qrB7Dj9CV
unXdsrUVyjjiO/iOzj7oVckCwZgv1eFz3IMn/tqQMxICALfCEkbnqkpuAP4U
QQBgzgCB2ozqCiz/SJGzhZrNa3yG3jiRz0DQp2FjpyaUqyc/1bJm/+7upckQ
sPvzYHlKgSD4KRmZa9ikwiQzGlPS5b1Rlou+8j9YtOsVTnFhIgwhOwQUAULI
xJ7kMoN6jbRgn+QGtMwrW1n2D8MxO1GjcWwSIPUltOoxUCnlQhqsSyX9HnZQ
fF/ULqWrKFic28R2SP2obqleqd85bk0i1nz6629PPdjzzsP5PclNpkg+XAre
9pR8e6/vKW5vcJ0+f4Ytd4DWB6qf0BdavwqJkv4h4jAe3Dp2KwsDFJG+CyA0
SrHJawkFBRlNpcO7u92kY1ebMIzl2itK0LHKPD+HX/IrHQT0gdy0x1NctSq7
iP/krL3+woUDSd/WADWXUFWoRWEW6AAPo9uoO/wNJROj02jEhMRbgs3J280b
e+T7DWZQ3ca21jYReuPkL6M30Z4wZbrvzX3SUMC121xHRyZ1rTu7+43CBYX9
vMelPygCZht+y5RVAjd78gAxRGy8uEkoZL6Ks1zjhgVEC7HRjPWhRBgLCxIg
LY5yjZkWJRJXxTXEDdHlS2OAdgSqxgMzQKP0bVk/UIsvdU8+gzWcEooey6H0
vjI562BAcu8coLnbL3sWe+4l/jKkbeaiZ79D0vD2hxp6ER7CpoLFPmoc0RNC
rUb3FNHkSEqtyu3oxKS9kOdkQH6THOi9/2k93LFqhcgrQgVm0IYwHtE/kA5C
y6/18jETOXhpgl52/dqafnyEJH7GTu0Dym6lneN18R3T5COoFITTZnhnIo5X
GkrUyp8rjC2xZMg+n5hRb54+PMLKZsHtc+LxfbW/gOhyweNBjnOSSXVJKvoC
RR0IT4V6A/4OhdVSUsiwmCtApHNuUWe/7hGf5l2jClfPx7fQrkiLc7e2vnLY
smGPU+yT/QBFtTI39FD03Uo3x/Mbhe4aaa5p4q4wUEfNG/EPWLaPqMIFI/Vi
5QJXIk91oax4gariHeBmAOaBCXMSWaQaTfnok0VHxflYRRlrhwiEz69OUtH2
yrfxTDigar/hly2ZmZPeWUrohjvDWireWaSyVTf2lTdPKkMwXWwNZjinxFho
h3gWNpCEhGjE8nMaF/6udGtBm6TFfaJSeKI43kYROcLndWW5cB9XHsusu/Vl
IG/O1zNbVr8aIHvQGiXCjZVt1SAoeq4vgbSwvnbGRnOfb09ZZBz81lyDfV0N
tFbAryiZZjMABL+1LDYL3SDIkPTahY/yln1L93zOckVU5T2EZFSSInb+KDci
79X7WcOboE6H4bxSo5bos8a9oJ+06Zz1gcrB+lHH4P4nASW9p7Wvl4YNDqo7
+1Qtgl4OCB9qEfb6KT+bgzr6zHQSARSEx55x/dizpIJPcIbCt6nm/PikXMSj
+p6M8ktMBybOsuVPxuPO2uN9lZfPlnFQtARsLEUbsAXhBXPGErAazoCycaRS
Ukg0FPt1NYxmzAHECNFObED9uBTPPbEHkK4y5PtU+RTjGsuNpYlD0JKfTmmq
ps45pK8mmlIBkH8+DgEUpa85EsqXEJ/HF9eFZvraOuUsOeCUptiTbdtrD1mT
7Ua1g26eDrRWunl2ogk0lxnMxUnZKtmf2d8IFPH2ygbQiLrCeiQf+kQB5sbb
O0u44aS1xJ6getPVDMcDI8JsNxG48nhuVWp2lyIkiyX+DGFAgyXXHgfEIzJh
0J4dEkAPQU7jynhbniriyNjTL0K8y3v7hHLl2qc484R8VpzytdqaFwZLGVKJ
FqNZgPL2NTsJfCWs8FEttfuzQN/rQjf1k/isfMh2H8XwQ+LNsPO9En6uYwD5
/5yIM9s5Amw/apyvUW9qQkpM4MZ1AhvEOO9M6Uwr0trl8E9zuec9eHHo+lQb
5e70XWjT5WIeRNtmiYpw5sNbenpXjFIMBmDaOTevMehDjttGABWekzR9s7lj
X0xpk8AjFTXIs0NH8Y5ResaRzwk7UOdImiTLjLapN9uKegSR1IhXcxyDGRAl
2GcXNq4r1oN+7EYm62jTBtwHA4QD8oXYpfhAZtf2tEM8d6EgFF243wIUhu8r
QWoaTvK2KYm/DuMcqBwVDbe83SWrboLHUz4NgDIveQl5Oz0idYNmmlvk0TOW
FRz7O98NlRgWbftBZHQZO/aMuSgq5gf7/8dwwYzi/0e6usJNrWtscPTIgAlp
Ql+kqHJgFOBW/kOAr8eJzmRcgf/nanjFM0+xSmVOIZByLp2bBXRoTgubXmyp
cr5HVRT4uk9GGPA7zNF5tKw0pTLD5+x27SeuinL0TYbZwY98cJsoYGGHfOEm
gs5t4IyUCTsUxNNoDnvbuJi6O5ZJr2paeygNQrdwt8C4XgSIrwu893Ek/ilV
x5v0gE7dzHplOWpE8xcEpBSoLCQqRFgBOn+legSepMLXjQbz5IonEsqEDto1
VMFIrSsL4e0furObR9lb8sX/gdU5+s0B2fc5MgmFXDKXcbpSZSxtYRQ28GKG
Syy9KKy/vVb2AqQHzVH9tHxZirXkuPKJgUK65o1Av+Uu5l8qo7/3KHip3lSh
n8M4MGqPjMOFR+m5WeUEwCSXf35Vy/dp7JMdkboiLkwXNSrxjco4rdCqBl6l
5Pt9HxobeEPx+KSHp3hTqBlgHeU8Oupyx7one5KNZHC4nsSawwHxRjfZvlQV
WZW/qUGn8/DjiDekHqUtEUQMGHWpisfr1LbE2Qqd+V/HP7oJ1tFYgucsXL6g
ZJ7SmPteg67BZsvnctgbwjyXFOEMjZamSoC5d5dt3nNigrCQGqfrfHlMWB0M
dvCPBcym0zPsMs9pH9imlTIruH3j7hURijU9QFycg5myrdTLxcQV9E5buvgL
Ynjqb4sI6rJrtmpZURbgSoEB4ny1N62IQWeCktxLjXgaSZPk3kU4C/0aD551
R7YFFAecwgaOdsEIfoPfYda1FuQKXfqJge+N3VugtUKDroKgokM3Ipp6S+fm
v0HckdAiNOMlNFXPjmHqOnwY5NaxUG6SpKkzkhC5K4bAXAhZ9rNUIk7QZCvK
TxzB8IJuikc0TNWgdBb7bJGWc31WSD6cTXMHpryCzWGbDih606mXAeZgXbgL
AHta8G4aZN2WJS+3cll0+TinO31Q0L++HvH23caHezZNj4Z5sU81xTWCM1+3
MJTlUHAx8ms56nImkER1ZEfNXZ/azJaDGJenDEFg8Bfl5iWPSNIAyCNlZ2uQ
DJnlJ18IqIHmnsT1Npflny6bmFewczZOo+0rhTvrAZRjBJNCknHEND5s/q1P
G1hJtILIbbMeqnzWwQrx4I8VEPrbDTlcHv9zoNiyi3DsusU1vyyhLkl9lSqh
VQh0C2jEQBxNTu8HqCStK8zEgePp9QUmoGeki4z5GMPXBMTdMPwysMuGqeyl
Z5oQ1VE1tBTUnuod/+10Ddz3sJOAQXkXOndYH0m4vmdBYSmDbaqz8HW+TeO0
QL7cIzeSwTqipoGIESpEfz1vA2zNycxC7fekj162tvx/pYVkVHBIMMhOYlV7
xgVB8ItRbZO8eL3GTePPd8t6DBe9dGfgxWAxcpF9juF9Kf5eIZ8UuFbW6LGm
E3LgSbXQFWJVW849Bvyv48f4O+tRlIq4gS+Po44Pxk7V0VhE6kEK3cpcjDzJ
htx96aOVndItnoUm4yQXDPgSFy1oqxb9qIHsOWMNNtTOFv5PrT/NC5ZBKYsf
JQbE9HS2iSLhrmsPVbZ9PckhDTsamsll6iDXI4QBo2Zc56awBkcpmbzCIL3y
Tv15mfl8LR3vI6wbwO13dKlABAFhL7f2d3mSj5Pc4gLEB8UON8ENqBvh2sU9
LihDNXbW+oQBxQySODHeYKO7br8crEWcnCZXl38aGff0oS93v6Jo08lvIW12
RZCjcF5WrXtFU1UiyXq27kfLUEubuPWs2CyMQsJZkimd4KNexB9cbKNzsSiD
uR44jl+VOuTaSJpOwNv+wQ7GCgzkmCRCDjvR+AcO/XS4OahZMYy91TB1qbnU
g9chEOasAqPDgQdRwj5cxu9MFJc9PnnH0j9lC6aFOQSyeRLmeOtmNb/N9rhL
SgjFPtOUnA9m8gHAaGT+dwMJU6WzZMcfrb8uD09fnYo8Anbj6LdD8Y/BVpFQ
+TsZOWV7hWB0ElZHin6iIM21BfDIKQZ4nqM59Tbgb8yFPG5Fo1u8j4WTIol+
yGD7mhbm3BB3oKO77uvZJk05Hs50L2h+e2lVVCihanXssIZy0/G4vdcwgXzH
3PqKIr7SCF96SclJoT6//OGMxggPGUIL7urWChZdRVyef0wQ7k9kONS0E563
Tl2ffYkZVRQlry3J7stWw+MD8C+dMsvm6QSsO0h3ivZO6V8U235Bgd2+5UCJ
WaZEiCgFGBeMi4X+mauzFpzSWVHoc9jkhd/BetrNFESdBPqmh9keLbH+yCT5
2IxZQ7Drxm1dGskgUNecBwOXoxebKF9dJ4MPKeWCBEXdsmbHw2LtEwduxr28
GOCwm/F0+zyCOnwyM8DJqF13VSGTVACGIkzF34wu8MV6pmAfxi7TVxGj6qeg
DoXTnM6ft9exfOrKQnZveaItIisd6gTBKMw2yWhGM5gd4MKv4vk2/HW1M1oj
ykK7g1dKiZQdq6hKAVi1RgqerAxwpdR05JkzvQiNASOTGKldCS2QCcCdPqYH
DeLiR5iVpo+HcKC7zcHqytqbGOTWqqG/s7DuoRchxnZ8nYEJA91Z6XJiZCHg
W1OY0Soi+gDkJUKvcs+C8u0MrRncCbEfLJGy+6ngqVEA5kPx69ulnovMBvzf
MPUA9+B2Cxss7lTvaISbhDPEAE4ktMkXFcuxAb+qfCfQalZJP/aAcwYAIkLV
V7qw2VtiVZbO8xWHF79mCe9BpKDWaov96yyv/v+M1LjrFKyH0FaxvOnkwkEs
5apRW6SSYwcyNtJUeLmmUMetzsrznyj9yy+GAwz3+PPgjocY7sXJCNMAqWTd
iDJ0cPq75+yM0wljY1BbbWGLz84n/UiNRCyRT80/YOHZpTtvVCiYiQVG7o5X
YxdNnceR/ieymMIidigE4bDvJwvOSva8hA4xJIM1DgtP+/dCS56qM8oXiRyG
TWweOckTREs7GUBhWVuuTzTk/r8I1eWW/5ORqpZHDUENeQi+1ZbZdVTYwHss
ePia9Bq3zQR00C6MGKbZkpftso1759Rv9Uj2wRg8ZfC6R3QkNKujCTRUCigU
pCYPvh49aAvTOHFG4AVOq0zlEaPnoamB0YDQAjLtU6lUg1pf/Bt1u/MsLuOm
4oVqd/fNOKkOOlPp0/LOlVV/3Sj9Fhm1etFsGq77d9PD1B3L+Wy8fBvdOcZW
BsrxnXQIFysFKBb5BDXlx5Jn5se37t3C7tJkBQ3CtmDQaXjOjdqKNG7NlZiQ
8x/5JRsEKmvey78drL3f4UfR7GSCZOyHcluaoA12wwF2cO+dKKjuIQxAj1dk
sxbQpn/5njRpGtsqqrOnHoL/FSxQ/r1g7MmhdzGx7a2Ee6372qJsSeZheGSd
gLNif/RAGriuXujNJaXN+W16wzTqCQTq1tLVugkyJjzER57X/zOCl1RZkOXs
FA/Zk7MPSghhuIXuznd/a1w0zdfktCa6XKCuALJ/cwcH3tLkfjuoCVQXwIoM
m2luKIIz+euYsM0rSo2V5EdaqonN2IVkuYffldul/pytyDlLJRc75LCm9zMq
h9gSdSMWLRzPqWMa6fDGGMumGbpJ+cFm6g0aXCNjbNDOUqlc8mKgdv2WesHV
RpxrjeXDk/GVvJMvXdAYcG7jjvCBzng4Nh0O69DOuR51+7EjnNq46nbdS0RJ
hYadMZJe+dj+jBvDaUguL2sIGItyOH0mntkrsjvBK+cu1wnVz8VKrNabosTy
eoLzVDvavxnj/hOHSbHUtdbg2hvhosQ6z9VeABkNRpBdeb1pNt9594Ss39J6
DxY8JaaPmRP8GndpQzaPsT9mV8ZtOmFItNStFy0zqokgpCnqmS1p2/LrMU3s
7u5V4GlE6ByrBE5XAthigu1jD+oTP5p1V18rPiKmI8haHmVrvT5MJtqV1hFM
UBsr7pGAT7X2IsBFtL5gFgFhSQatFJONdyf7hEvPgSyCDo+CZjr28r6/Vy1c
PX6wdbpKNL2uJB9z/PSOalFcbu9+vHAdSnOOGtaGAntqz71khoehu0Bnp6Gr
fvJTUwA6VpZsVCU+BRwzV/r0tvK5MJZJlH/XH1FdGu/QVDVrgxpd/XV2LkEd
o87oVKUI/4POU5XAK2CWALs8TgDTjyi/15ABpJz8wxJxTlUCFdtLl8uxY1ZF
RXm8+82f4qDvoorQMjLewP25RsoM+9067FJYZ9bMpgY4haFepBLjlw2flEXe
nK7lqdJfptjzRMo/9B4+keyfmz9lN03fI+ZKNHi6LEKjMUwTvigl5m72/J4F
1biXvyVDc0eMXt9L5DVkrNW7b3NsZXouWfqJoE1SsRZ/xuKzNBqnfKNhrWqa
f6wNC5RFrpwMZi9x5pTOgOUFUADyFNLMExemBzsVdaYLiCQYNlLCMtkrkDRz
CYrogsJ3Tm1tIPs1SygOW9fYALfkUc6eh5qdiDotUh14CE2VK240XTn60KvX
18nTYDRFLQ9ooDHqJAMAkth3aSR75Po5Ds+3fcnAXQg2LbBlbY0n9s8t/18x
VVOjlw9Ix8CPzMwkm8jBJqQ5/RKFByriB09Oa6wL3t9ZestZXfHcXKxGDbjY
aLLzMaOrrEkvqk69p2UOONjMsjW7LMkfxs6/SdzIlrLd7d++XbQ29ymsYjA6
3cIHbEP6utmkAfJmr/HPfKuvODeZvyZ4J+Ju/k9f1Xqp7gFQTQT4BFrnozaG
e5sVUsT+iIJjSbWNa6Ce6sbJ19IgNvv3k/ZzOFY8GR1XwwsWchO2RrRodLCS
MySDW4zGsFto2VQYYAXhkSsh29IEEW4plPq51cuz60XPRESoc2eXxZB9km4r
b9Es/vxdH8N9kxAvDCwRuPRPWnt11JaPWVU+yXvGelmGVVegH3YilJk/hIL+
Fj/b6GiDySLjINMYvVmhaDbWGm3p7EzEReoYETELRRVKWl+VC83LDC8vd5q5
1IdMKL9BJUUZ9evZ0HzHN8p243nH7IT7xE0SdvOtPNzAhatsTqZTFE86dDga
vgq+xXYM4s9rIqR9beL+LeaqCJ2zF7FRbe2DpM7YKQ7D1G2lp8s6Jd7xFMZz
K8qyZEsMJpVXJfmLqVSCWHkeNDTLvqfJ9JcSycaXWiWhIrFiw9Y5UHiV9YZr
zlztTuXG5ohWiehaKKDG8LulQxeySBe3NTl8S3J1pNcQfhrLkipzo9RAiSEh
IkApWdnX1Mjoe7yQt2YVPydCJMBCv0UPTDo+8ncBqfB3Hj9JIj01/9bTJIfo
cw9MfEUf2w5zLiiv88KIolQxESbLDY1aPpbtD/BooNRBiDzv1m/9edpap2YX
Sr9sftP7oXmUaYGdOjbFCpplvWMIaLDKdWs0z+pqeBfjdrGilRjIbyBom6cb
P2Xrx2zSoMuo+++LKAH/Jt1tnGF5gjTsAn+JhnggtwxBofQJp5WkPKcRw0CS
4OE/tpHTAmfJub7sEgKfNueeHJkKrOhVlc0qwnJNfFnmiKr9kxRjax5PP8xu
ck77VBqBxapU27dJa743IfJXbjLzv0ocDRXf1/NfPWaFFhdcxtbYrWspmkaD
8dw0OFRfHiaxK/VqZo0rP4w1gvKY9/ohrE/ES6/5/hZs0+zWwch1de1eK6XI
dyaR6ZtpOgRb4SQ0Lzsy0ARX20DbOT0Sl04ESshWb22a8ftORP/V/Ik2Vg66
vGswenm815iFs4kXMFd4IELT0H342LxXLUiNaCI5THQEFGrMzfhmnFP19/LW
xC3Ohxly80MhX0N6fF91TK8c3Ppfb68fWSgZpuVR9VrofjfBY1hwwC6FfaPp
k1oDvjcv8dXwG0yAu1oNQWzeFdqIaJK52fcriyirmUVgv9tyaiOoQ5oApdkK
zC/mgq7C1iio057rCpphxt+WDaxvC+KmQhS8SLqvhRTnJCBteLwok9upkLRH
PmwQMD+R2hR+cVu9Fn2l5vYpqz4/+5N2VOZXzvgAOFIKu3ArJ7zmrv1iPEP2
dxA78daBCLnpyCtMqTvcbA2Zyi4dm2MaXB7JLyoJE4XhQTfwnT/8x+cst+HE
VknBBzDnk0z5sAqIUw1dATxOc1D0Yarz3iIp7soHR+HbZCZ4hgblVvylZKBl
ogb9eUiil0O3HE8T/4I6cQ9ypDUyPrePr5pM1OFuDawlcir1iAgJ3TkFeAhF
tvMxh3kaw09UJpT7D7HA8TdHmo5sksoukGQXWTdr4vbF3t+iKbXUD5hwRjQq
J+EuyxLWa9C0VvvWhEZUHsfSNrzWTU34jGUsRJLoPw1+fq0p/FxhZNRJtxAX
pq0+4nzkQdkWL8UQJLghtuo3C6crDqeEXUoZm2qcUGeDkfVwDxMCugPptyBr
wnaI8tWpCB/2QBVS+EcBN+0T4JgcOq9N5+bHp47nYLl/EcdxEo7NeBZcmexT
g4tTwj6noZ/RnuOdtoLIWYwf8GcozFvknA2hzxGMgMgGFha10GfxOBW/G/PD
1lvGHsvZ9232NU1fjHTR+ZabGGT17xDT1b1mJ+L+qZlER9M0/DO91btfkbuT
cGF6fCPo2dagqDpfhN9gp9/XgM8H/mRI3P7ebeTVikiQiaRHfR6IudhoT26M
dRIlqhqnTXBsJittcifslOI5Plsr8K3vrE/jHXeh25zjMLEZ04vawReDgojU
O+NQVxp4L9mxx5mPAbYroU4+Lz4HyHXMpHhJmM/sN1eWhxYRIh7L5QUafdFR
jVnrpv850ipabUPlEUA0jSsirDAA91+3/SKGh6BdAIvp7RhO4PQDNWMtW8El
bPHzlRhaHtLcK2OaqoJ470wLmcOjDIVj6ovMepeiE1PQoj+Qqqejc0Sd+Rpf
ZAIODiTv7IEEPc2b0UsDbEarlcRjxKcRHL4qDkWDM3qQOgqXhdrdPExclzq1
n10lnq8958DXTCuoHJhVuQxk3PAZNPWcjLiw8TcKJP5Uzh2p3SaAcHbxD0Zr
8a2TUIFxl38vLGIe+WFpkOxUSOesAAWHh7W5WQSokYRjhZbqnZ38jDBWAvPR
7/k/W2/QQBjXlhc7GNQ5iZaI3iCXEK2wqk3unTaDL2NnqaLG2G1L44oIuLiV
1CqSunE35vOQb4g4Au4Gr05BAzxDenl6Hz92moPIUb/ZbDYH2/8NGk6IXvrj
WgdLklWObX/PGO7ipwc58oWY4A5runXqZ/Az12OSCxD0yDPqqvoK3TjD0bpO
jMgZry5T1ebg7zy9cyrcQf6ht55mvoHCsq5uK7RxLTy2NHpP6TPIWnU1j4Zt
plExrrNtnCCobSt4pwPVEsKGG+1jC9pCYSlChm9i4PzSYkyQed9rZy7oRDrt
TNH7+gkEJkt7OVyhyIRqBq5z47QCILNHBoskRELEf3OJQbjFe6cql6YOJ+CU
6y8FAMSPYsd2RqA89zhvKz6JV2IJW3oBXgTAw5A+61OMSlZXBupNBl+HhFcD
Jahf23NHVgqgNGjCMw5fzjPOQOxsQ8yx5/DKAM0E9qNOrkiwBrxNvsSHsBUy
JlmqjjaBo6VIeKjN2AvBc5Y8UnlzCOiLoBy99kehSNG+BRZPEgoJ/ZGd2aoa
bZCdaFtf2ie2W/lM6OnijwNcTacHPfkti+JAD6pu6EDaCTPj3VTSl9YP12XX
mIRpfaxlSWW2p5AwMkerUnmqcugpyNENnTHQnk2S65UHyzrZtkguof4xBcZr
tNyf01U8LVl6DXC5yFwZ1rPmFyEPIC5oG0eo1RMc48EPvpltU9VvZJob4zhJ
N0aLnGigoIv+vugd9gRy6MfPi0cL/8M3gDsGB9sIgp/G/aGgD9UaB0rIJHIO
X01iDdcnpYL6LoPu2REWUVgfRfrIiuuetu9JiMDKz5p0gjufq4ff6gJUaLhF
bSwwhYo+ant6am2UDETZzjeZZKpqXFyeyiJ30VA3L9tRIdkfWu68vcDe6upr
zGNH1xvuD94umIWa8+mZuGneXjv1fnJx5Hw9zgfTtlwKBXETIvehs5ixWvMD
A+BaADtz7B31NP+Y2YGnR2YYzr5aPixrHP18MzyCJN7oPshMTNcHbEnBITuD
IqOKyBvL1nQx1tPs5kk5UJnt+zp1iWtwgajp5Zs90lp1Famu/a1fzDzfD/e5
TQRefdiHzwLuQJpemxO3/zsrhNJMUY4hFWXkUbtOAz9SoxqD5woOfDmwZwji
78RFbYF5NjFNQFRGrxPw/9U72H4cw5oulf7/CBjlS4FtjLdcG2uSP2FXDSPv
X1tZnQj3yK75MutrzVDYiSXxXPaferA91eJXnOxB+/nwnGlOmZ9xkMAV1RY+
nQsFzmncuuy88DgQlfKT9dxg2lyn5QcwbBq3w/zQtCdjkYLMz1zJ02ka+29z
LQ6ODgF9DV388fimOIIUu8HuckMmIX7SH0cnr2OlOmIgxAVYd/pi9jGPv5bS
SI+omLDirA1CBBnWjduk5dC7wngkHcDkiiRVrY8y6VD/ouYUIT+Q9hrpqjed
9RarCwY3RNpZNgSs9ezeuHEkgW4O06nVNOO3rkQpTC3W+8bRZJSlOGPR1SRK
CpYDAXsUl5z35sB9FbNyeXlZnOqrvmYyQzaNwQn4XXckKixOBqh18eMZ6m1h
vHjC2Gle9lMvM4KPR2wqztWmVVmMZgauqiCrYDAnf+FVwABYQC2WXnMy7K9l
jgyUfS0JNw5XZhwr3MC340W+RAtse3oMNq70+mLvRDyVCtMFq4lmoFTfpehp
e8g++wZ9wgydXUZtKbRq6QktDlEInkSPftqX8gWK/Kp0GkrbXWcqQg6iU31y
4Y3IEUiUkRw0lce0rN4XxDda7WHwFM2KKmFC9E0F8u7sYJGvnp6jctdMgCg5
XI/pyJgqMHXL/wNNiuELM82R4KhraJ3RgQsFdhhCX7F1nEV272aG72bG26xY
w0u+61mioU3sEnHt78TL6pXqE4yCKqVpIETT6Pj/7CtLMJ+OKoIH7oeV0nzf
I2s38uObMLWoQCpaDr6aE0KJC8lIXoUlZMnoetgt/3zk1bK8CO+dXbawLksE
02344jGlTGxfZXthu/tg+f25d7WnIXiqu5v+jLshGOBdoGhj1bJeLB6lLqrp
BuXJ+OcGWuChxlNovzoHpSaiF/Nd0R/dU9b6x0QXH/XfBsetKMrHpywhyXlO
m3dOsagrqVOgwdOxv2vT0477JUpY4AglipV+EvJ0ouL5beXQemHvsYdN9NU5
Y2BqUt+H5vO/W3+VS039Yc/U/8zmIZBMrTRs0EI3bgdpTY7gAIEcGJ2hhpy/
m/LIAUGBFHl9DcbWM71mxa2qW8bLq/ptfQGMdmhqIn5Ycw6EiVf/a2JQFacI
VOqi4BoYBpw3jocKQCCUTIm1/j/rwxYIz1kloqgWVTVt/JUP7L2uf1/darG1
x8jEsAdJQ+SxS+sGk5KxF3TlC+SN++ZVotyXqD6jnZDvIuXZ57gI0Pxq259K
MjMx9twk/mi7kkB09YFgXBRSB+UuHpb9KmDp33G0bMeyNESXWbUl8EP9Zf93
07qDo2E/R82NU2I5o0oCSoCzRbBfFRs9OSuzLSMl9Ljn1+RBfawxohd84bGO
4W99rv0IoStONERNlHR94bDg5tolRPaBDTmRQSp4CxCmh+ZoSnujuanHwDIg
e7pc/ceJUrfIYcSrhmhgaphXmfsWjVywMJDeqfjQ8Lmtr2UW8atWk9q4xjpG
aAX6r0gF57Lvl3X44sZtjMJatGjR97ygsxATkIRyqG8t1AfejJzmGYeVw8s6
JTxFintcGdirnpq6apJ9NlGYZQ7srVDipvT0Ry/Y8QGPKTFUWQ8dhPsxnRNo
SqKVTC59Au4nodmqzEodursgCiTwMlZ+9EfRkXE4wAF4ik8eSPyhBco+Ti9D
ulS2C9nSEbhM4huX9MIGwbeZ1dose5ubT//pZZeCs8u5E+AjT/if/7W4R0nb
M//YBz56C0bFUK2kp26ihjmRosLChJEFLEH4L9O/glC/LSxfzRNwd8US1iMQ
bKQXXh1Zvj2oRZYfbLI4y0/V/m3pT6oP/9cGBEVMWekNSBJrr1J1tTwrEQFJ
QVPQ2BO5MmjItEQRgL9YB5Y3wwTTMogzP3FzR3N04bM/JgOaMLC8b7f9QbMS
L+HdZh2Vm38WeOY6f72yiFiiDmAEWifJEjxYsAOGC41YWf6ON7zzxTgWwM01
htZB1UU4hFSU2cujTeZE4/U5W9G4Asgts5g3tFAIpF9xpSkmLiqGUgxJ2lYj
1zgv9YFW7ihwc+IAU5q4OMMqt5IostKYidUOPnGDAEi5rr4+JeaqCADWQxnV
Ph7Xha2B1XwKm4/m7GGELs9z0j+J0SUOR7wLTi6ZUF248mgyANP3j+db52g9
P89RCGYETOzs8WDlKw/eb7WVRnpgwBragO1lhxAZskGJp89VK1NZsAw4UJXM
Z1cCkMdQJ+wutL5zoV4zeDqiDRcLxqw3J4p9iyNcPXXFIT/S5yxt+ZYDfD6P
ivJ99NZpushluRHUD9W0btFaHzXBwUOBCTVamQ7LF4YGdc5x9j7C8McCV6f9
8ZweignAMaQ+d/g2ZJjEqI51n00F6FYneII+vxW5hHY1lx1V7UMtMo26X1MZ
yJ5NW+Z794HHoXzAbnJj0dtvncxwF0qd//sHaRNI21TzofutcTvGKDPn6zmS
lpHGZtbwYod8lLygjmZq4pD/nm3xhDUIW8UeQnEqC45x4+VjLUdZJF86ev4L
jVWs4omnLfq0kKp0fToUWLYf4rdqeyc/LJmVA1eYmU1xXrmcbkz27GXlCzt0
k/9RR5YN2ZfwmlQciq63pmLkxmesKiWtVA6IiI2t4t6szINiQ5ICwJRH5oWL
BNIjEO5UCOzhBk2GxlCix7PVUQzqXLRsEOdGS8zAFvNsmfYTj/ShOoOg8UJ7
x1ProkUol0Yx6RwYja45mfsl+FDsklkxQCeSCbcIfmaZdz3sJHJbpnVkhJbP
PkcwvIDDQeL5MjAvSE73eZaUyX5Ujd7ViwtGGB5YVMOK6M7rJZ9vyQPgm8zp
JBLfyKPk/PcjEpHKXJmBIFa9OAWofEkGuX7y1RViVhWAqZYJMY0fqnAqgciN
Ap/lsXMLC6LHcr5s9FTeFqL7UVgJ+ZmYf7/LBszUY6su3o3wFNrc3Fx4TMOT
GDzeLeX9U84BWW9//DsqXkWC0DB2oVaGw/W9cX1NQscVYv6F+mjdoqzcR9u6
dShnZjbkFSmSMF/BG/5fHRULY4h1gx6B2GW2AJqw4MO+7Mren4YL4h9xfKuv
RFoCNtkk4Vy3jPPkg1VCCiiNl4CRAiOrDn2fYRHAK6MfK65lzhX0jn7Yhg3z
bbE+ELEd+zv3rjt8BgkLTo0MhbCFhxoK/BfLZWjVFFiSPhEIwQhxLVc048fd
mycjzTElzl2YCsuEOlEZjhX22xOEzXg7X+rVXrAy7rtlMqG5RrGwaYypwIlQ
wq2GA7V5zsRdZUwF0e7SB+eH5VxwXqMnlItzA5sJcU3uCMOZwyP/Ba2RyYxj
GF1sWN2Q8C89wNkbgKXuj1v/api5QCkwI3ZVo1AVi/FxV/4ZvrP/1j3MKURw
U4M24PMpNjrd6jXVEErg6NmhJ+9jpyUZhC3asjyYOwBIS1Vz4fWuWOwiQwfx
4rGhZBwyItryxJ1I/KV9orpZoMoXZIFxpdHrkqDliZ4lps4gWPZJhg8eb0H9
nZokFa4Evv6X4KOOwloLen6tAifaRKwHMjhqUougYzkmIllUkOXDsAp2R2oh
A88Hsvh9HjVj/ceovGgvLTEuOTYuWr/LJhqu7bqVn9FJg6B8klA0SyW6obqP
mklAuCnmQnnPEXiIg53Diz+I30oFuWzyCf+NNXj/GTsU3lNlnIwuHv3nMddd
S57Q4NsMwD7fk2gl7NkV0EZsyT3fysTMRtNUubsWT4PT4ZNQaAMJBYgs/0Rl
O4JX7bw5N3dhu+o6n9PuQQZe90oalCfT+JFvB8tvdRpqHcOT43n/KLHBnXT+
n2yxtHvZbkxlO82Sqe0iH6JDj3jt/OSUybj97BXMHeYhYGmYEy5Ht6BHL942
l8NP+UB+huTouSPTdQdzhuf5q0uCshPTBY0IDwmmjqK7KLkYDJtEYqbjdhvx
mNtx+4XkkfJT/5CSBH4s3BS2aTdaSaCQfl3qUviZeRIq+g+lN+CygQ2+czfS
rdXfBEfwZ5aWPUx7VRo8ACZngmU7ZNNc2MSkBkKxtNEO6UIUhc5mICbAP23p
jCOfa2u3NVhGIGJHAA13NuwFMB3mfgaEePaLGDVhrRXWs9YF5GeMvfRQN7fM
Zdq8YOtWQCrXDdvJ1WdO8CgNroM7dHvm7crN73ky+amc5NUpGJmpZxoVeL8l
w+2wImxAzLTlCk51Ujbep4RIrTXGCc2MK1cyJb0SFypmj842YmEJtfaLqKDO
fH70qRJcxJ+/WXH8asQ23DyhgVThu58i7pwmRXV5O3W9D3D4sxZ/7jrtvskk
7k4aLqcPFstHv7AU5RxlRt7Zl9g/POnI44K/AlrwAjOPuX2CA38cbL+5rT/n
Lrzbn9BqinjFJhtvosBqEoRYY9dXW96uiwPdQfYuPwJvpQijoorYsKb4u1eq
dEoYt0LZ4PHYp/DJvS76aOE5Gyxy3oSztn3fJ7kpYN3kqBF7ail0/FsNU/7y
5dulH+bLQmbq/md2mdaOMIbzLjoQbu9uR3+xiLyLBC4UA18iS/kksXXPPLxH
un64bYkZU6qB885Bwl1lqqWV2+5YEw/uyOqSEqIEqcPgYJiKWAUBk79xEgxo
jNRX1NJBSmIe5TP9m59DHQUdZewFs5eSlEfmM6dMEsodeiPPnSyumUmGlmNQ
T96wa1Y5YlkCBVPHAHZB0QpeWzmEPdSn+X2zzKmYKKAciZzI4YZ+pLrr7Bwi
pa6/9MhlSmc8rerdEvac9dW0TADoYTshajaO3OmxPGqKh00qRXBwddvssKBx
Am3Hd2tH3CXEtSZbLHhUUfocYNrotV1d81SorCknjUqLE9LCliPO6MMO/5Dg
8Nx4058ozyG//cfvlD7RS7c8x7LzWh6pKQqBp+XDInwRYla9sJgE6MSXm8pf
orDOyFmMGOo+sTIBj6kzqsOijp9fC1sNKSEK+GNHRz+fQ3klXfA+61qtdLFY
DXuYGd+iIwP02DquhLY4x7A+aktJbeqcLYMP3LwNbO7L+MpsITBdZRnW7FiN
/ns7lMBL2qkTxRQ6KHCAmPL/VA2oyD58mIdN0XhVbYCNLkjJiyJW25azqPVa
lfeX9Z1mcJ102qs/Il3LC9U8tZrzq51iNMag8a/oGOZpEZ2qj7CjszTjox49
YWT87J00Cjrd6aBACXaE2F8lwDwf0vN8QVMzx3quE1Dwl68Q/GTvj3u4UVCq
mrUYjGcOhdyYPJAIhb2elLseJ8L/E72Sm9bJJZyxUW+JQnDllImfikn5BBgK
n9y6vh5jkUR8sIJBCDPlOoHDKX+AqLHEwNNwIywNXrmqpkzJOQGtn6QIrdML
CCdCYf1Frb5JUa05o3CNfbGD83njRD38SOnl9TsgqMj3X6moU7u8SfPyccew
alawUmj10erAZIveZnky9xm6RdhL3Z6QbS/UgKU/i/P756J37mm5EPUlD9AH
J+kS8KOV96ma2D2U+NSn5bd3e2U3rSmnOnk9f0xXxWM6nwkAtML/cQ5YQEqW
NkgBsR/qz9oGFc+Fr/LN/uBsLv0ce5dX9MFOu0gCBwidvabfo7d8Q4pbzo1t
h9bX4N5t0zBukd6rsbHOUZ3ciUia2qSegGmdc2OFEEmgmmT/wWuvNlrVl3Th
bSThLRcZ5o8kbOgPWdztDTk9P0pRdLWr4vJahV3KMo2oML8orptiEG2kQAs3
+UfqYMN/8L40qHzX7/r8uCgHAQ1GA5J3go3Jx2ukRL9zGk5sRTJFaKC/OC6N
+YOkAJpwTka+Cmy7XNmCZYkQ2A804L1TntZ5mPViC2rDTamHp9TQNg9OOVvX
yOr9SUDuMBhDEZceEtw9XkhRt4lKeiSmER2yvvmIEM0pepLvJEEiryq8t35N
r1RBUdIsoQjm86dw5neWWHAO3NreKS9nqxyFKsxlGSibo/463v7jFYPBityU
NVAcGVPtlniP+vLRXfa08KmFhoRRb1wPolSHJfuWnED0cs+OCkUExyZYXLFh
F48HQ3jQsjoNbjd/n7Wawtk/6bUtrTD1Tv10k/Vv97L9UX7awdhSn0HozPDK
PFzqEXhneOg44NKfePKyp3xN06FTbkIj1omMtpHZacW4Fe6b83e/z1Oul0PG
sXW7ukOisdH/JovQAbDxpGrM9ySPq4tGPKhGzt3saPjrgcnwj6Ls/L4w+Yo1
Fd7yySK8sXb3YpjTJR9HiatGB8LQmqOP9MJ4RmhKh0dZt5upj8Yvwesaak28
Y4VukR58LmaCF5epv49mSisCky70CYmMk5+WIPeT1r4e7CqUfdhF79zFm2Et
FrXEUPt9aoe6xvcw8vU2bUF1jsyoquNhs/IX5jYJQWnPzVPpuVgQXU75vHmV
wsuzA1jSJTQ+6E9Q/3Z+QZRVfgdKPijZAXE70UanQtnNXCqGpyYKorM5Gl0A
/0GtkjDCw1PfO9Gl9w1k0NFKlHovZLzrKs+jzWZiJsoi5b4UAad1rb0+0GW9
NL6lp4k9I5SVTnzcLXg1Ix4kccnROj8lkVHXeOnP/KaFUlt+616jt2jZA0id
1GecMaCe9r+6N8FLeRaRdaKETWSLKaXHESCvBdBGUH7s72oqTVfHFMH6Vh/y
HUk2pg4ZuNmPoN/ehVD+20mWe3BcpEz7EE1f5dhz8lrKFOquv+KEGTr0nYUK
fNkcxTpClnu+B+8j/JNhm4oNqsbT513/XgWApkwbwHbAF5Ya5l/LXRy0ntFG
WWyg3Se1ZBXwTz0qD/sAZ72wmTkDxj1J5eumUOtgcq+gccqcWPMS1ybXv5kA
3LXpoOXzsiT5cBggcVBRD4S8NueO+WnFPnzFgXpVSnUhmgqdxBXM3aZEdkzP
hxMLMO/5+CiIFWCyUmAreIpSlnbMVijwjCs4ix8ypkPj2qSQNndWSs8VwYNE
2jKlZRT6yeW24uNFxghtQAdPMvfaaljm0X/mfAQkSN52RmmGdVLWiy02kNlR
HavWtfp3HxuKC+iq1UlzA0RhlZJHGP/LVZgJlzRFYrE8/F9snk8PmKtSN1X+
OlKCmDNODAFZ94H2iEFiLSFvISB7AcHT9/+wSMgOusQrmsiWxuuEVFs7bTWn
AsrUGW9wXXEu1BNohsa8PCsAf1s1mi1YVMx1+yO3t0QMSiMLGXFXNd0MXleO
b8P8YarcthL22o+2BXvsl0dpJ6+Civ1SF/A81itx4Q3PJ2Etofoo/Zk4H2Y7
CfahXBhN6nW9ACazALH+hJL8tsnnaMOarJWoAU4cexqebVKUzZMJYtVS1RKW
gaq9Y+gMNKkfL+lBMgUcr0+r3fWE5v9D6LY+0D8LZ/43B0hXjXQ/qOAsmAYT
3C7lZMb9VjGVO+fu0+J6nP4tvnKLM+lR2jW/11T++YfsF7jMz2ZQeUPfgWCf
as+ip8QhBlGQZZcc4jHoLPpCLx20JXpM5b3tgJajy1q3vKiQ+7T3eBaNV5iX
gJE/Po/4iTBpvyxctuzqSD98FzM4agupMs0EvO3+WAWPD0/WD/uXuM0j8Ge/
nbFaS7WwtMuPhEE4D/Q/f1xs2xBe25bN6Gf26y2Nv8xVrZ6tA9s1zlolgiT9
0l220qR6Pf8N6ogK6b0b4R0/7RMOo7M0mTV4LEPmzmqAa59nzAVKudDWW1ts
AlE0+A93y6VOccpvd0svW1ONFntlRlN8mBAq97SNCC7C7xZbn0+04G1ehum5
XVyc3QKNaw156AsmBLY/Zhr26jD4hFuxyNU3L+qE7mrVcMuLP6hf40U5PaW6
UoBzF7PspHnw3+UG1R6jKv1jBD1NSKyI1n8puDkQq4h6TykIE6CXSJhuyTsz
FedLPSk+Lps3LW1IPePJPAdh1VR5my9DUEf4DNwLxodUQVAd3ciNpsGzXeRS
fzz/OKIzEh095rAi0dbEmqiCita5D6CPgmtlnsTsl1UQQCr78oPhzxELfVMv
nfKouhl1yi2XkHI77G6hBXxYk7+4ol7+wtEnDqQYr3n3xLAzz9Ctc/9cu5+O
KZwDnvPTlt2RGzLPxlklIYaFcutn0UHp///JOCE6TV7z8WJgavTtIUIJbBy0
23U4SmlYud3IyKvw1Ndrqb91Ll0qjOy/dApBY+ySCaAzeqjUg6pn6V874D8j
uZkU7BmE+nCaq9RsUzpRIyKSS4SsDnWk0l/32WaMkL8y4406AN5drDaxDrC4
ab1JL5VlTgszlCiJHpe7ih+SYimRxQcaz3/sCBucqz30o/EiT+oqM6NtuyOG
c1pVd2GU1Nk8Qyfmb6xd0hJQjWAZZRCGYBn9hnQ+ETVZ1bbHdSNDKqiawheA
xfHoyd+Q8Nz1BDic8CJ0NOuhLjlMVo6ATMnbeX7QYa9IvsgBgZ885UK/CVUU
9gSZhtazcEXMh61q8t9tEdb3ByzneyIkJ01uflgh4DusRje2/E7bT7NBml9A
pjUZ6d9gDbc/HvC8TnjUApCgkJ4cGMfUI+9UdsPp25kRkC+PSyH2HU4GHcfH
eARNm6M+XvhLydFmvKA2XmNgDmlsQbxkgWWqLLqXf/1UqWoUCRILBBQxj7sk
Qd/Zb6ff7Jk6LsKV33U4itW1WfbF6+KNIpg/svGjjiNbhdBQmVE4V74dAAC1
xJFwe0yCZX5C4x1UpU33eB+JJP/YN9eJFWdwD19X2QJmeJejucsLqLJdTUfo
FxXoHVRuteH3nriyZbNTu7/pM2dFS6rjGATHDfIZ4gvbbhsvm/MuxaOiZL51
3g1ZSOi74wLFBrhVW0pqV/kCexKwHOiFazeqc6CQolp7Ey0h6kVaBkmochgA
YKTdk2MboHwbz7z1tNO7ogIdpklB94nxjitVb1Na6b0KUiKb4qeqwwHFtHDg
lm1QVWK6uhSSnrQ/pC3m0dDelldAVJU/J3zK+XFY3Hp2gc5RhNyiN00A0By2
G290uxxKMxFEtvbtMXllDVs9C/Hejdvls82sCoU5B4JmiF8LSkPbyq8WndMv
B1KKs/wZ94efM3jLWwNnZERsf76iwSZyl9UjX5FprX2LR0oNcQ3uWXTQrjRM
vUvR4bsjJMVBSymLorGWKQMCUj3HsSWBuCSAPt2lTbQ5bboH5hqKqCJYVyX4
0Ln1HEx56JQnu4gR3FIL3t/4NYr2B4dYaQsEtpg2Eabf4y/vRMSkWPe9PWXe
YckwWJpGRYtFy3zq2m0uwSbqQKVmTckXBqIkzoBUHsw2hgGt0s/7NxYWyQQN
TC4LF1gXsmGA3lnDRQ/k7Qu9cmuplHZoQYwimrytjBgKrRxjNC0/hTKGgyTl
eukjdN42Tf+Z2pZJ3Vs7W3hyhwi8BPuUQMNGeqtDSIXyxA3WoP/P0+08kfTY
zIMGX9KtNG9CWAKJhm/PQ62J14+hFmHGiNgnf/sSgMTTdUIZBNrujCItl8IA
+1yzgoRpBXV8n09EaasMvTufmMJeAuWWH7FhE+IED908CpW0oUgJMehknQ96
7CuZSFHgWMyo/aMQgyJqQNr+1YJiNhcPYb/8iap0qQP6uNmPhCpwN5C8RUha
5Uezbp5GCTZGvyS3ESbeQXDw1/tIcb9CrbGfU6RQ9QFwG17tM5rjWQ536gGx
LGoB7YTh2XVwwtx35nvItFJq0hCUr4jdGSHY8JvNUj0iEUC02kxL02vEtPuL
61SAWUbClVu5Uex8hPd4HaQYYu+nVw2CpVyto2hHgZeZ9aLwOg9zOT9Yxqvp
JjO4Fw5wVvh652UXd263trwo8AOTa4kBv52U6B6XNe011YjwbFXyjsTRbxtw
3/mFhlvj59CivA6qj+NJI6IDK7Nbz2iStWyXciQK6drviWseRaVwUgDx/din
zT9D/8pr5r+TjnpZDU3q98PgXznwVf3PNm55m7xCHDPm17zwOt402DJqgfbc
KVeN6vJJUFcirRSdkCok2x4aqj5Do9DEnxiojSxiqFcRtsABGCcorvbRWUz6
Ypn1VnetjzkwFFhSH447/hNXI7NJ5A+xpp6gAWwo29sZm7uA/gNesgGv7f9e
/D2Ug++eGdpLDKbX8+rpzmEbQHSi8A1ki88zn0R+Cls7KDniCfztvzrHVS2r
VVADMiXH/gV1XMAvzocOnYkEFMNrj8M7SgUzTxJzw7EeGLy7umdTovmMMLZk
FjTCtTEHX0Mh1AC/kD5aaK1IvRQHvJI4wVdWjhD15B95on6bVTsBAChtbH3b
mFED/RB9M9Q3NGHoeXb0qKRuBZuwbxWuS9b9KAuqGs12IUQDRzUvSS0Rvm0N
uwHPtzO5E98SJg1j8ZYBT5cVZtDLV8zFFZ3/4kTR7T0FbjJ7X4GunkhPoOoD
gfmBmbfqFxipAoW93CFI1WPGBLsLdQDIpL9aJ16xOJGt/hUXmOFXDk4Q8es2
h1QSz+OriLQTBEq1rCh6ZcqbXEsz4SAPAyhct9oToPdydf46UYmAvRw0OprN
d8OTVjzRtYOgpi6wLZHgxouMYx8ub2YYVx1MVZQOvmO4MdJUqjIg3YVvhbT/
a5Ymyr/g+nkAKg2KshyA0PFqkSDuUOQP7twmOnELllZ9OVC0NF2v1zGuOYig
KfEkRufJtikFbCqvPdKifs28kF/4URB59uix4C8f88cmfhf9k4K4KAfF+Aqg
f3DT2YBi1SgOf1kVSRuNLLkAIDbqK/TzK0SjGVk8IGivDO6IjbAMxmcLIppG
feoaMDv0hJV9zHvqJ7LeFssvycNdKoyoJKfZGSM+Li15IuhB4W6R9NdZFCwb
H23fg/jsccW/cq+/r7eoNu83oK4B/walOoRUR59K2dYEUqdZRhq168iIPOAZ
MfiVOy64vyZWaACX5xMTupmpysrWYpt8Jgv56Vew6aIJMSotD5x04bzz+2DK
44NrbzbLJcDf0MczawQ0yGVgtkNx6l/aS5iM6osSsn0ivM2eo3AFATL62kqZ
EPS/pcentfY1Y9FrLFmZU2/mTRcDpBjMy6yn371t8nj9mpH/aetnIgiK5i+I
ydeho70wDmfzQY6aJE3VgHMKPLCCahxrok+EWdk86/Yha8g5myWixD8q6h/2
IlITc7dNs8prrtYB+LE5aOt9p9WPXwopvjhT/J5O/gZ8H/neY03Tuk2QMsBe
4hGc96UjrBVrzXfwn1pf8oth3fscgWRCl8Ms0OO7cE24v3KxigW7r13CO7w9
Z0VvXULKNdtk2qTCTtz3iOtfVhV5AFFE0h6/Aqb3XhqkQBCKGpUGjg4tllB5
7WjF0EKweMqDgScUt8dx/tPALm491NzMc1Fk2/BYXndy+eQ/GTcaIEHAwjxo
YLPKiC/hp1t+rFe0XJLZ8qaODd4W6XRgZAfLo9OsiEczs888eJtddXbK1Rz9
Q8GIvs02TZcoKFzQJbjFsABFgpmpJgVdT00+qREti94xsMnZvS5dNZIPG/l2
qVNHfuK6n4RYonY1g//29EglTsuuqHOOn5ZtfKns3FU3Ev70VACFLBHMQ2ZH
p1KPIy+414Zp61e03PiEXHLrFKTScATqC8Du9vhJMZ+JbZMbRWJWohc1GGEY
hzL4bmWq5xo0BjrZmfADYwwcc40iYtlHlcoCaSIdI1gpXFI+Gfw5m3xkhp0+
LhHBwz8yq8bUn99gT42f+LZWC0SUCbXxCH4o/D/yxcW28GaPbdFX/P9L+liV
xf5thvW8frC/Ujh5MfCYMBBpt5+a2St3JWXSF7f8v6LhTnd5WdRkW+j5kQXj
3oow7t29wtTv18YoespQvR7R1pIjcbWkkLCSEwQ0RxfnL130ZAjID5TGvvgN
AqWwbtEJrL9wRvTtgTIOOwiY8VMDMQxSH58jfFsJusE0atG6RtQoLEfR+ZIm
dJPtI6Rttnsgp+d+fg7ZVRNIqJHsfOqt8vlj8zQWNHgww4UZ7mGohUp8wEgv
ab4A/sxGX9/jan7QIpxTLZu5EJoukYXwH583y9EIa/A5dcfKepefaUX/pTau
GwJzZOTeqDVY3fjqV+lAk+rZG+oPRE+JKqWWjW1GzQzPVHwhmJiTvcLGxURx
vTK+iIQeKZExv2pYGoBSQV1cXVeQP3CJ8ptTCHRkAzUjOeVfN2q2np7JLJpW
dCesFbWJJdlWUzTr2Q+kZ8h1leG3/6uqCsa5vJBtbB4MC9olY4NomI/go8j7
L6kVnzLr2aybKuglGvDxYgKtUN4bg5YpRuDxX77nxTvOXX8qKGE8RooO10k3
ZXS+Z7YxFjMncMmxPazuFMwZzwi6tOc0IDlze8C1K8NpUxoreDNKn4HhzN2g
hvaoKTclnMPixAFbbq7vioedq4cGzDY6wUn2eYRWJPQ90vSOTa0ou7w77VhD
DdaZlbLAdHlDK1mxh0lRJbuWWz8h90WlePjVpap2yM42BBOcmkw/q2YcqTh5
2cl2q9AQPDD9aymjYHyA380ZKROullYvNPP0MKcYrkvdgaZ5fSe309HgRyVA
wLW0Qth5ooTwJO6SBfyvvKlsHbcLg6YD5qwf2sUdQ3LvYEOXDjscHAq20kgF
Dgezryw4eDlLxRKPodtBCjrFEwqcJhFNooHeVtkKnTKM4DJoCd1biRlFb0re
xI36fvSoNe/xtsmcdWNXXC6wsAqFNIJ0uFXGqNCawU246IcO7kx7w6TGeRqU
JUAtuoCcTtUdfj+SynqmDYCyW7k5d3KcLGJ1S+0BRVGu2cEJ85i+GFLnePvO
cNGYEBNnLNhuOqhCjRc6rDI44lqveY8aMWzJzdB6WRIAyznE0Hbm0HaqeVis
7a3rIODrn0DvMEcpswWhIqkxnUDG+fEsoN3jp4dUJ0+GXKCk2G7/Is+JloLX
g2r3DxlUfYhF+tFRcG1hMmlY5Dl0HI02im4ipEeopOgdxJ/CezY7xT4Be8Kl
+GcGxZkLRG4bJP4NHHfpPBjiokJVyaKsc5am3BVxmTlscflTKWAqi39miS36
x/nKa79Bs+72d2HRefBDjN+TJSVPhrKVRTsLq1RjDvu27S99fDXJEup+6cwO
Zc+Bhh6TqDoRHedKqVhCFf89r0TH8FBgFBe5EarcdGjxqZP9TWct9SyCpxkq
7QrSAL6vdE8sSXwAK28S+el6NDvSTfoMokcim0V0FQf3xwdH1EyqZnHVLEU2
Y0g1YnuJRaoqPYJcf6QLa2da4SKBn0p9FIvGnwcMJBuHwyO+7lVuVW1IZzVi
Tj/Jmk4sQzl/CmU/EL2SESV8TCxUVrzdO4iR9JbW3wCv3GwO8+w/EtOo81q1
ranTOR4oFHDy1vEcn5vJyD0l5kEsXyzoi0MT/Rs94zOaS+cVBxvz6BJXaOUx
AOTrxOL+3aFsxTIPF4FHtU2uEvy7/byIjdobP+lixxfhZm+r72lK3zkofJDf
hYoX/OPZs0Ddw6ulX3vq8RVz7qTrPtfmJThg+Vf0f8XyEw7jSauAdeiOT1Dr
oA4R5ZwoNfqKXnqV/Ajx2/Bq449x/hZONvAWtSaY+r8ag0KlwKMJIiy+ER13
CP81KNgDI2KoO3ZZeOss5gstp5AAoaB/Z3rF7A6wa1ENUJ6fiL6OFtXPWHzd
0if1gZLWJfOYIr70Vps/TWLcuHRKcly5FokyCZ1MIEhfl9HYibKeWFF8Bury
5VfgLhgYXfH8vuopBFNVZ5dEfr6ehhJ4PQGeynpCwzFgNRp629IvO9mP/vMu
NaOxIVmDVs5MerwzNLHqJeETF/anGZQr6N58yGeO9WHeX3b4qfnTKEDnr6JE
ND1ZqqlG7ZK5SCmbs3WNdZj/JVnhaXGStInaXjbaKuLr90R7MjbJlMIjnPIL
+EU6Nq2MBB4K37/BqeX9eobBM597IgYZT1Wo43t6awNjQR8yUnQ6J8jYIuEW
LrxRfvxqBdlx6djdXH9J7RpjFJWcgKxACgU+DDj1U71cC27/85+EL1n9U6Ly
rtPBJjzgzdn0Q+xg4rakBCxHVl9PxEmheZ54JKMbhTVR/YFaBoQzMO8g0Q5Y
R0L9FmIobYS7ILYhRKFTtA90yOmYtBBIE3FeosD61G3oEdbs8zk8vKsZhcm5
UfUJlJDvsDKqlhH/hSNstJP+2KouIGO0DgfXhOyQW7hxvug+NDu6G9zIaJYN
9QJqO7GvErT70gobIXUEPvXkkP6ZIruMVwZeZa0Aq7JYQ7h6GZn2VK9G+sMO
nZshRsdIK1UPiUmydN4moHc0WSEsgCGmifnYDiH0MRltBfqDoTykCsue1/rd
o9odUn5EQp4LCe1+1ABnJgNh3+ZJ1vFsvVewMdNqhsHMJpWInAyZ7nOSM6HS
4Hy+2WF57sgcIoVug0vdHVdWBJCGMbi0hlJJqx/r983S9hvnNyOaJE0VudkI
SIlmy06P79F+yb7hzvqg5uupHQqlMnQ+TgRQtfOg1q3AHVaBvDY96C/Wv6B9
OX/5cFDDp3Bk+lYR7S4a8FDD/v1ozWwe0KKhPuF82cBxTa1CQFnqG2TvazpY
10Xz4cE3eZ7LXzqbwEBzXZUwtjE2ptQ6eLZojhg7SwUdBi7Apzk3OExG7rZ0
MYlck0OTK9oUitONkhRuCcJ6716MHzpuMwDDhTGGxtCzagR2TcO7oTSwQ7C1
nmtGMFMrhR+JgZa9Nhk6E6I+IrNfR5asMBUwQSIYlw5NkDFE3q+tbLR8cA2d
45KnZoJhI2BKzf/YgAoyM8ymp15qeoJT3buXCl5757ruzLviL4VvWfqGYXLR
vQGBXSfAzunL2RLz4W/bqqVRCW7rAHy3CR4j8315dAJtWygUgRmuGy3twk33
+7o3hQkEnTcHDAN18dsTO/3OKIqhArbqlhcQfOrE4sg6pbXLgLASyowqWpGc
dMerxaFyS8Dpo1DGahd7WJI0c/UhcO32Cuco3R84uiYzE0lrzdcEaJ5HhhSa
v1Xicx5EC+mM2rmIY3RUQNBbk6BjSV1AyWdl9yj5NGvlwuvERhx8rqag07r3
57ixrUCXu+nQvF2pDHFE2NUtLI5CWL/IWGSTeWAVISv4LWJ8AcXpRLBqL/qW
MXWZz2d3+ehq2KvQGxrpYEoQiI2M410D41evfPXz/irNXeYaSw7tTMt1jjYV
tNF64n/OIkPLUsd6iQj1hcthKkgZ04vbmCHiWJ4dEBSWl7Kr68b8Pe4l3P0H
/VwnojVjSRqdFb/gmez8YXTqvH4WfhO89tShAk43LTz9Y3lhB3HjqDpJQvl3
5aC1JYkkFCofZSgDEAZ9TKe6J2yidCuHV/NhKE/t7RoxxarQkuC9/8orJJrc
SPIAeK1cdUGhFwUwIDWZ20F5pEhdIXdQbN4sTsxMFCpHDNJAH/ru5jYlY8N0
50v7TI1i8Cwyi7wnv3u3+9Xu/1GbxC1DREHmI1xzT7IjTKgplZY31xZmqM3N
7FsyHoQjSyGBesHE4QLO+W+Lpgp/j41SjEGN7Wx2nnHDuCPgL+E5wGtk87Hf
0jV4/Dl8+UuxB7qTol5ZrQNpq11SWEo08XrJ1c+lB+b1PYuke7OuuX5Yfqo1
0nwHOIaDB1TQACqiI2XJBBNsaAtCgkGqJxJs2IqAdIhlezaxGQQazF2UVuSn
XvQ4yyGzqooYRNawNoeqRSRyUQZGWQUBzcPhmc9+NfVFLD68g7ft2Owi4UxD
38TM48j3fAW4P7WQt34hUXH1ELEKqlJWLIiU29w4wjiLj+L/3y7GG37/VV4i
ACNlJorhKloOwo6+VyYQyFf2YVl88Oza56KT5UwmzFXz0HwZI7vF8gnnmbDg
wt8Pmj/5n8qtcUpTlQPEM7w9tVoTEXEhwKa0P8/BOkuSClQ7ySmDVVzikGF0
Tmn7W3ta9wVVWEPa+/FjLZR1KGG30iqXrquEChXym8TC6IQU67pVwuLPBnVa
HbXLAvV1yi3Pz9+GnUB7HNkpkp9b705YZ5GTiDnUPHUx6nVGzUkztUFUPAV/
SDS3L1EGGOl3Aa2u8wKqwBmS/FsgeBtMmm4vwFnQotqPnrmDDtkLXxVV8sCV
1rJf48keuZhBplb4Kc323TDmThzSpozB/t7Qd35NYg3Q1fscT8IP4/7TAjhe
uu86S4Q0VbhEqJYuaY0sehpuI6q3g3la/NbAY8+8J070F0L5j3rOoPO4RwZ8
Nl5sgQXr5u15n0z8xaoRsYaqmo1GLQQ/EaCrl3Uj/0/DOu5BZWWXbLIDDsak
ZdTdE7PrvQWe0Vz3E3WrGbEjEnK3YFAYSDS7qhMXyJZZiS0ZZAIk4q4YSXXW
eacvKf2XT+QkJSMlpNi8WPpyD4OFqUQRmoc9uBoqAhdlW3D97qIKEoFSuQqd
5/odkkmeGqA15tm222AL2nBme2npsfqONb413Awqbj7k+3MlQAd1738OcWw7
IzWrVFF0bPw9pxk6Km+u6UjCWUPldMaVJzDDEClQApGp9wBeslt9DvWk1Msp
jHUlPTitCcyX5OWc8LdQ5MufYFi5xc5Sox+vhUfIzIW88bQCc36XgVH709pW
f4ZfG3LyUiynMRPSMzrDb7eq5V8VB3hu+KGAJw+Lk12NfEYrYjcbRLUgZcA/
v+jiX2MnikgpNmAz8hykPHTBekE5kQfLL+rA0vOkxlvpSSx+T+nw+O7kKViS
TE0TdN/cyg2cxwU+plqF3bKvpX1CNkyf5zTALMcnihh7GwhqAu3Y39pNMaWk
nL5YjnhvltrHpTQTzCCdeNfmIr14MWRMW4Wa6LFuN7s7bKCD89/mHf2zqVgu
xfP81ZjjbY0CYuYHC/S2/avz8QIlHvWw4bfSXMilUN9C4GWVzMUUVZv6Mtd9
QoSKehCFMEJaO/xTA63UF49/ngGtNpLkSloSgVTAdPFg6LUKGv9SSrbcXBmS
3FtvLq3zLxGuj8j5uz785WTesKrhrNpKlkpk/7uctd7kcY58/XN2yad7zXzZ
9L5H6rqKOjKiMaBjJv3Bcl/vOm2CTBurNdoxMPW2+/Am2rS6rG4d8EWkaK5E
N4AIHyOLYzix7PKH7LK61y038t/sS5UVTnncTTrJnol8T0ozEyig11yddiXd
89lwYfpX3dfBshpkzbdsHxHO3GSvRXWjHm3BuscoCDA9fBzZkxlfz78WHA4N
rSWnLqls9OdarU1WQ7aNDMSyyy/0D9rXFY1dgEswwjNZczXx2RjrBOMlZqtl
Ds5k3SIhRM/wPSun2VFnn3WO0St7+t848sSfcutJgGW3qk4EsfQxLMEFCtCw
JyiVIxY3DPMXZPH3VR1BGqYFsMQfBXGG0rozIj9Kk+ldtzBhn3BKp1HhU/jh
WcJG/yh0Qa03nXFYETBCpGPB9ik76RM4ocvgY8xjWdTLysF4Cc04IcRW/nrk
ThvOauRutmXLejVjQMnEsI4t17bq6WK2pr8gNej25ZsM6OBvHz0mXBkTbSxA
UWAQNtveaRtMgOJWcSocdh6CDiK0tQkuhwtRCIfDwt2Ku0LQgEFx+4XjRTU1
uzwaIuL7jy/QXnY5/dzb11PFnl1jcdR2p2e4ig55WV++/WoLGrtylcaEJhdy
yMjUXkZpo70BXiJcJLl7MimIly+QNBhi1lKCqGLQ75yPUT95cRp5UK5vxQlF
Of5bgnWZbehVQmo/s/i1c0iAxxVREzlVirRJy4Oj7sGYB3pNCDGtmtaI770Z
EGXK/IihuUwQ0fuOxNx+K/RuvMb+ZtC8/9O7+ezWE2uQYbFSQ+JW+Z+44Ml0
Ki35mIi/LJoMNHtS8gJnNAhCdrU/pHBZPkM6p3JTq1ENkINcc+HskTx12d3y
pdu+w8HLbIns+Li4ldS2rrfb/T2Bi3d+qA6UFwrasCBpOVeMqu72t/VLXRFv
AU8wpN6yLvzXklY3crRwYZ91cyaHzE6WaUslN3t0UNykC9/R5XCB8TvqsxY+
oJEO5P1wC80Wo5P+nzQjISYjsNdXFCoaQi+/mASGxckYeGHmng5F+d5dql/r
ov/hYcdqXQYw86d4FUHPBzWz7tgfdHx1xE0GH68H29tfkD4X6KFeXgXAoxyU
xT0kDdmTFomyAK6iXOvTvDLONeSngyxB2pDcLwkqjcLFnyyyoSx6PFdLZ6Yy
u32+JaHA5sPwFBwfoSghy4MtZJvXdSckQlmGnvwgN2qUwb+4FE/tkm5+i9k+
ZXf7tpIF8uhCrCOtekFPxcJv7rEErTLRPtt0ERK5HMgjM4NRgt9zrKteDEBM
2z9hrTkugmu76fyUAOXA9Vz8R1uOkVBCzd8EUjcqF/0XsUwQQNIcbDKg03xZ
OI9JsRqNTbh5r/UHHQ/Jpc3UwhRlBeEc2GNMNu+p15FuBpwceLCDvXFX9ZV+
IHiQUtjIYzrJ7ok4J2ryHc+5h9HQfZzJeNGIRozs2M6t6E5e2FIr0QSrNRx2
JDbWlgPWRp9JkL8RrFJwqFE4gjvflbPkHcldk2VK+Qnx4772APAXb0h/YSMa
0tnfARV9NoPswltyC7xr73qVCjVuVU7xxGbAYEfDj2UeQsXZsYasOg2SOCOG
o+SDLNaHiT0TLaKVMvaNoL3ACu9j2s1g5T+B2rcHiWgw+XNEUp+aMHF7707z
mcCmYJNW2Wv0EbhYGJoylF7P9GS3ZK5VzoN+vXDTOtHM8rYgg1CiO4Etwu7p
+8apVXiUzU6+jABwuLWBxsbjFP2EaMeBwAdocGeVRpyuU93DqYFmFff84sw9
FqFHuiImhIGUfXa6L0lR4IxbYcePLAX3v+UET9/FAVzVmetwjkddGovPOIyt
FMe5PX7LzDMWIxwFif++uXIKMsbihIvo+5ySKriVHjk/K6uFtjZJIjs0cLsr
y7Wf1KbkuX6UrduLVz4NGawlkid2tex0QWCL7Qo2xJmf29vrm/7oDcouAZtn
ZAGeIVSvKd6W7yFM4GtxnQVpUMCADIaeoaAOQ3Lg+5DTjIzAPfkOa3jruWeW
7avwvJMzOW9hJpsjk9IN+VKI7PTE9mZgCj+LbjwjF0+CoUsVwmkxBSfB/vsc
rwucBIodCVRAy78HuKWvHEy16KnRIGodS2dLGUuQ0jaJUaSLiT768ol7klvj
JYxxlmqrSRVVD0X8EM3OZYlP38V4a/O/lswuZBYWyN1ub7DIExnRb7p0MA2f
IE79rLXYYMiLRadYW7s4ZwkChWXgu+rczOzIVERaIjB3ZgW/MKarbrRJ7x9k
RQJcD7EqIfYrp3QQvWrFJg/6JtfzNoGxKb9lytbZ8YVOWdKs4rGiMCrzniDF
k2MmEbQ8bwAgBVVH5DJstD+wuheP/jVLqdgxBfrb2l6LfABPjapS+hPREzud
QDxBdmCLU01AC1zH/in82LvHe/P5vfmyneL4OLUohhwZ5ZtkVhV5ugvjKwOK
zgtHa9z8TiGJwnkwG/P3GuvN/NtfgZG0CeigRidd2yQio0iGGcvAriHxcJgs
j9cNeOqIp/eIj0+PL+rNeO+AOidqc6/GSG/q3St1nsJcJmGmBN/5qFTH0LPo
wi3gUDCXWTkImJMv15WXwq4oNykyP4bGF2q79Wc52wO1SlU02g5dD8Ww4O72
DJWJNZs8lzOr8FYpRR5ZKkzTioKbtRtNU64Z22wvGY3hoLWNDAahytbS4+pY
mGM+o4ea7jZvfy5RxKB5/3H4VD1U0a6rtY31wTxlR4t9Ltp9wyNU7t0dT9cq
ZCfxLakQhFMnmEKCv8Ut9zRRmi3CmBoqGq0BL3Xr11p432GqXVffhyC5afPx
GuOZMY7V2HHyFtXxnI5mArwkqUUlxHfEjqrgfXpl3yEvXOamQ84GXnY7ond4
aFxZge2D/spy+LCvXhrP//1XBmBoB7OcuQkRs/cT369W9/3cXFxagJ0NghhF
rOBl2b9BGrqyo57BdP2009DSqfd2UTa7nwEUnxcVclGOaVhm4jSbWzgoZsq1
XSAiZNnhQ5mFfMfD9jfgAXpMiMKGrdklSim0c58J+K2Q5ZntlIyhGcZ+wF1t
zpT8WdagQHW7vucVKWa9a7/8uOSde40ku260Y7IBXOwSZ9jOqm0JG1oQWzIm
YF6lRrkIeGJ64l+2MRVI0KauhITdjaWe9zXqUDTRYzjSHb2adq1IMTcgKSlH
5JefE5o8nRKjmyPCZCxyJKGnBFAUhSr6VXj1iLYLLR3P06jxh8ddD5dy4lAu
DGNA5FwMQopwkBdL+2xMTHgQCyCTaM5AhEDJALAkUbMVNBPDLsf/J2CU7hkQ
v3BqQ8JWmEMm9X3INyLjBICahdOBPgVJEJA9y4r2hyKpJNms91FMhi21WNyN
CbA6Yp6XKmfmAh7mjSP6cjCAzkP6tP1WBDyjDyPG18KT5vLorWat/FhgLmOP
JJsp48XYz4iLk4qe/rJCRIKd1yGvX+f2QgdcMbLut7/b6I+UDr0o80BENSNF
8DaAY132iS1BAsCCAqBZTlckitVuyaFPdvTKWsmZhfKm/PFjy3u4ErGIG1UV
ZciDlKx/Y/v/6I53L30ImV500icl9+gNrG7rYi1YSqMDCfU/ZOvkz7iHw2u2
6HZR0QbFUiONQtUM/shvEq9ImxLL8i8Poz9LdF7ULqmD5wBPC1JFj4w5guQk
/tyHGV+yClq+2iinohzv7qKLs4eB9bGXKrwPjnmZ+yleS35IU6/XVZXd1tlN
4YFBkIX/8xIuUiLZlcNyMAS6XdxaCNdBLGX+C5scVjX1yjEK6ezUh04VHQA1
rz2OMDSDYDHFxxE1Ccm49R1R3k+mRnM2BV4HnUcByJF+AAFO25XSi0Mm+GWF
Tp5zkahXWvbYsIR20lS7mhq2iacoCMs7LjOXfH96DudNHJQHnM6yq4Rj5eS8
gnWnfQ8FCe75KY/kw24SSXIlhcHo9VFjOAq3d31DA8ZY+C0Crf8GbWwZnVZy
8SiyLPwXY42uzKv23MgjSJPGsitRyp33uxzMUPJ3WEt/YtT1nJEwsBsnVBk4
vnVqaCv4LHqcTXBJGCVp49u8vGJwfQhzlJiUKrpZzfS/1nCRQvLnZn88k/eI
An/dNTACihH7odlkBQBL2EqLchsMrU7xdsLSiI3QYzmSsn+0D9D0TNKZ/J1u
DD0hRydufmQ+KwcI3f3FEFQI9/rVOC+0gqriQPq5qFb8kGJ4Y80Ti+p50UYy
hP7kUE4HQvidNlct+cunKG4Yqgei/GSObvrogpIiKFkfowKmWXr6PuzsHnDB
ZzZSHocbZdvHHbZXYNtJVSe1j4FsSQdopdcfdOzWXeLHf9uM9/GVwfBiEloB
K6bFhIjcCD9CW1ta3uBJOVlIBhNgDZpH5snGKAoIAfcqtt9XM4tKcRpFliT9
HD3Tfm5evgcOIFzf2DRcraVYq9yuokudfncr2bYafgmM8B4fNAvJhnzRvgGj
C2P0dLcNoEnG4qDIBluNIXw4e2jJJlbAAVBrUHCfP+MasGOE8BUflGrrkLn1
TDnBX9TUT5UEeRKL9L/tyyojN2gQWU8CVcyI7BeFvVOBTRB1A/c/hhRPE31H
dV6UyrZDu7iJsLfMkQTfc+zbloFIvizhkm8cTln5fFzt/yPjxLDNfSMi+Yzy
wU63EhQrb1v1FsxjGCkuwC30LVL7NuqV8NUWn4H1TU2bWgklEiOOcIVOxUN8
SN6tIAVhOWPizr3NcZQxMdvvXJL+Cvb2XHyG3iaPw2D6suX3mZsdbtrhpZvI
TftsrpEO1LizgDZ67a+Pqzmp8WflfTinhAqlDNQ65XbE41GgbeVIaAbO46fm
kiclLiedom3f5TgfOGgN9vIiNa4xgog6xTSZNaeRvG2KRXhLU0JY9cam4D0g
Lx1nJ6ev8dNgCJsB5JORIm0MN5PYvRzAMDynEPVjxfg0FgxfFiNDmV0k8QDQ
9w3MaLypBB5i2bKOCMjR1oJ8rxB8bKGVubOHgkmsuGHw8aIZU+lBscTqgIWg
eTZOA9iAG+Oy0cpNSfNHeue6snq2iB/H3BumaduswyomFwfHpa5OEfY/KTqg
1M8KhQvDru2QrLkt4srx0kICGWWhcXm6GoUD/ucBczVP9KtRJ+HuIMP1UUDX
9ySA6TT0bi5xH+XlWghqhb0Ol877G0NrdZOE0e3YNJizMp2oj3GKrV02z8LT
Z2wykYRw7YQw6V5+RJzlhgTINdbZuiEOgXlPVMIcoozKXilfdse+9G63Ip4Q
7w8HKyU0CgzjC5hpMNHPCa/wcQmS9StCE2R1jTxqEsq0PGwEZYOakYp1FVbR
MfCLPdTDs31moqYOZnh52IHSyr3xHmWTx5YAq2mMG9Rq1tKeZ7c7HWGJshNV
1TUO4RRS4BT6QFqNDy7P1h6/ej8n3vAtkJxXMQ+bDw+2hLWm6Z/AZZpPCblO
hZLtiIjWA/4yeXzWzrN8TiAn07/fKKZ3g8sfHODgc79mC5KqFebZ4A8CVadI
7BvJ3M7Kz+A8naGGEDP6TN6pJSOMnZxu9YzDcKvrAueo76di+BrMDglZmQ3y
e9jnawA9susXlEeQTUDgxEbCrIEkrxNmtXWkheQnOEcyO69JdUPuahC2+2Fb
D29KSftLzPwALmTQDKhVf2ReO68PL8HEYFxSxu1a+vtsLDBRhRKa5cimAkqL
ODslmvfKXqZUWF4ObUE1nmA1sw6y1z3X2WsLDd6o++cwEfU8IymgzDXJiG0t
cfYf29f2zW7paTA/9thRfW4P7PWeo2smaXHOu1zauwJ/9ff1CnOo6H1eyxLH
WRdJDnY2eqRAkhYH7P1PAagqDpwzIdSrw7q+uA5mnkXijnFFsxoU7SZHZCq+
DUnsoaP+4g5wjqTJ8KzG6szNfFZa+sukJb9xUxe+wix5rq18vHAOc4uKUJlo
3k61+W2Avx2NzzbfnVuY1dBfo4LTw5bFwV7GFQ9Rv7xvziqi1BmzYSdDs4UP
iueiFb4X1+1vml43oECm3HFZI88wQv+G9468FA+sP2DrqpkoAV+SJc1kRAnO
q9hoiMfqL9aEPJD+g8w9UQHW7XV+Si6WYd2cwmK5c/rmMtb+OFQ++gvNQV54
o1gQUUWnClNRSlcFZgQulnvtrTqfRVlf3symDIrx3FeI4AP1It7NtF/vGCjA
sW3T6UlaCHhM8HQRzbfxc76X4BDnKVDcjSBP0gmlZJUx52ajEVdmabx0jtKr
aayyLBCp17amPZEE1cmNr6lQsEpoZzhU+HrHnxNwBrCRUbjC+lXH9dNNd8dD
7yNJtShcFSJhMAnOPBa5aZFenc6OcDABskvG4wPPk/s0+QFAANIvaTU+L8md
KpDqi6fjwvl2mNjlPx/3ydda1xL6gbjZvYmzXym/uv6r9ONSXi2KEvZ7BPdm
vHUforBb9lQTkJK0kkwH2RKbZup24zSOShwhv6YV328+lABNCr3QoDzpoX0T
IgS//IpPQ0jae/6OwHr8kWb0pz2r1ii7b7f1Zqse36Jm3SG333+C2pqlVKsS
96XMzczVSOvTTru2xdCyOUhjPpTpC0K+P+cNr1kEl30Aiz/IXW8nEHzDln4p
QpgVzl0S4uoQdFqmSnvm0Vg07ytstWg2jjkFJi6vu6CEYFUvJtbGHaz8vI3o
AMBoy2p2AAghL/SSJTz29HSFPfvVqQs+yo1EEIrHuWPQFWwLLnHlEVtq6gCd
SO6H+x/ehLRSolNb4SvqcWH9doSTRWXVayHPXJ0+uOvLowOosYzrDEw+3b7z
67uvq7hrRcqfVBskgiNSnGnSNRFTeq5elUFFC9wF0H3Pbl8ZQRTJkC/USKcd
BiuLArd3QAgOawuFSIhUMYJ1xtkkhIyN2dckeYUesc3wOnzhidzqu8jEg+nh
RQuCIQJi+0i+yc5aBXlAsWNoBlYDhvgnbnK5RtnHwSvQ6joeu1Usmbq7i7tb
DJMYKgF4dRnop1WzCZXlRDTS8M4uKWen0AvICPytDlpmPlTFJCoL3kUZsL4T
GPxKPDk2IUmLh3yI0xDRT8HmsFtjHLHuKcBuOBcegqLbHn/6shHrWnfiTRKo
jw83PagZemUi+Svtl8w106GpsNEcojU17XmdzBY7lGeU2fE65Si1uY020FWc
/1u5TTGnt8HLxdLfq7jXgYh8c7FSkKU58XatCAucH72WMcUcRarkxZOb6c7J
z94/qJPQgRZGGTtbRhccmbO53s1kEFRPpBjxLj4tG3r/19GXUvIvVFh3lqXp
+//uAVY0ga6A8yJZm920HoJkl7QY/hjlnWxbnUD7UyTqYJnsNRXi0uP6TP3d
GrvUkgQBJsbTWTTltK16XClUEN4BtlUNufOiNqOMHdQscwMLLYXtPOJPR+2/
TZ0jYmoM1TFdAvp6ytcpNca1hg6elFFkp3vzO3u2H9PByfe9cj7Ubg0iwIfl
ISuf/7tRF+0EhfF76ENK5dxkJTQ7eoQ6q/f3DR2D9TFHxm/8Bv6Mswbrrk7k
B5XWdAzQoQHYd9Y9cRqmL2bZyb3Cs8JttdpHxUCSfoW/ItO4z3Lv9MJS9AxJ
mPI3P2kgR6somVSuIPDKEl/xy5jgBE4mGn5gf4LflKzeQUImMWnIb0fDRGOI
yEJtMYw/G8nGL4X26knLnE/L95EBYFTL3Ots5SBSVV6vAa2VK77avIRcxW3R
w5UoPlgU7CnrVEeZmK/LrDUhpkTVZFNOoZPZbGS+itx2iy6Xcmz6f3usSPDz
iBwWUs9w7xwaV58ip1noqgQin4nZkDvhXv9OjNqTRyxRIQYHt5i7qnIhdd6b
OvrprCusByslbTsHklA/0u9Fru/S5y1ob02iKSr2Y8cr1Wdp1lxHnNccuuyV
uD7FW57NB64yaQzquoYCR+j+7LgaYUaw54KHgboivdXlV+onohmS4FBslReu
gH7NQ6SgRvWxTx4jn8xDcah/jCGHOUTgztk0u3x5Jq+RpqhayAkjETivkTy1
OPHRObaTALaPMFSGwMJwVOc6UKLjCHHPnZ+f/AFMEfgufn9P1J3h0kCySraB
nMgC43kaowtPz2y3k3m+HFz3e2CYGNjhPyoVoz77rIxgk6isU6Z6WJDXE4Dz
3sggcH+sgUhZDxtv+muIufM0ZR7pyRf6Ol+T/hp1Vb5loMM5GnbPKkVe/dcS
PgU0Fv8Wx7oxV0j77ua/0lDsjZ88HYQM5p3XgUhkhSbHOIbvRaiWM5RARauA
Yrl2tpDNYv2O6CdsM8YuazIjO6q8rjvZ6hGDWF068eikMvXtQR2T+gtI/Hd2
jMjLpVMooetwKLxdlF1ArHPrndduug67FqSz0bQ5g8rcw8b/unKt6tEURpNY
GuJAbyjg0RqqIGFGRGnRbDgESeHMKT6XdzeJEeqLVcjfoVNgyxDHFM8Za6jB
5Sirs9ko0eHMQ6ZAPgig/4yWYVBhmgMtj22RoGwX0R6WAsB+dgoYj2vVGr2z
OtItcE+q4DyRqVsvJstvGHUKb43QfAbEB1+hYd6zau5DjVL4GuSCToLX2gTx
fVHtRk7TV5hOgHIBhnZIxgaRlXHKeIm/yxY1SgWLsinH5C4nESdcgrP2MMwu
KNyp5m+zguZoUYEt4Orn5a8rqpU7zRIFfli4LDWEjclrIhVFGw7JakWkXMmp
XlcZuzZS6Dq0xeSHnk8xQ/TOMqOzQonobsfEEVy1Bb6tXIFazfRAqOfkRDTS
Y/JEqNLsLLMIbCnbtkGpVefRg272mKvbnTKlKZffAR5v34R96M9J02NGzKTQ
AlSpvT4ztYR12wgX73NQ3D3E2Wbn3Z0w5b6XFHIaWWz5HRF8ZLhUioYH/adS
HoyJ2wT0YlWwkTvWbUnsM4LZ23tz33peBnoS2bObA+ykz5GbRSK6TrQ6FUvC
z3YcIGr0Wwua4QU359gekNXba+6weQo4HJAUrQklykwjsV9Mv+MfnIJZSDbh
IwFW0sCjrFSJm0Xuu9tsgbQGXj40TpJUuJfrc8vz+XOdiu7CfC4lL49/6+Jx
pwwOJ2ZIvefVF848zpT6/DwQHVwufMMoo4sWD4sDC6L6L2NfuxnWsw8EHpFH
EO0HiTo/gByh+l26CM6StfUT7bUC/enj9oIcJ15NgjT49fdO6gNRVAMfig2H
50IN1Lo1KeXDKKC0EgsY6ddSB/GvFLbBnkZasKKO9iVJOrqhAPO1/N3qgHtU
20ZcdFOxQjDHTaG4Hz77QWGSui5y5QP+GUbaSa/nMj0CkNSNE6sZY8ngl6c9
RxvNxcpyZkgVVt1BSn168m3eqr44DIZzRLit4Y9TaXPBo+8a/Gcuf0tx45jH
065j4rywWDDx51EKndtW0z081qXSVfP7c3lDo9jNIPRB7eV3IAwd9V2RvLtj
4U8tC+nHcFO6Y7BfrZZOeZY8xxVx7qQHWrYzmN1rtUDt5jAwyp1KXMkqnLVD
Lcz2Chf6xnb8t7Wkij3JUllUry3P9gs/cnirXmA7nF2prnYUA+XEMqNUe9fQ
l3tk8DKmdR6uJx6bNFWzqU9rxlXBvX3lVR9SucUq++moWaRQ/eq/BToLj/Rn
Q291cgSgQG7VgYjSTrSnNls0aTpb9lvrL9qIYuKVU8diTNHmg59i99i53+Iv
T+MYWb0rhbq8BkaildAkbM4/U/L+uTSJIgTGhljz47C/u7QceugMtxFWEz67
KpSlup0XEao/58Ow89IebdzeTEIb6ld23s/wn9M68WY9p/yPxCmOACdF3UNn
Qq2Ps/pfQMdzIzofwyD0pAPNvyvyMw67thlPvEfNWcQuNfekQJ1kDdpYCWji
iWStDE60WlNMCz011e61oUyUalvB+f8xOmssJcSACnRgOlJsb6z29rVsQIkq
ecvQZRblWj2WM6nZ6duVqE/jHduK70NwwHGYbZq6AtwcIT4o0p8+ccn3HKle
/6Hfq9za1wouo6nhppI+1XYWuTEr8d4OqHTWfHNURAk7wMWEkumvcaaK49C9
yWtmZvg6XArDReCH4Cuhh/R2D7WnEt+t5mqPBaZfqDFQNmg95yLhG8xXUT/K
nDPQqPphq6gOj4u1r/N8fWq2ak4SAqn/B2GCwqKW4Sv3L5DpIw6zbyrbtoko
fsOs8AXv6ZOPkYXmG/p9hKhpewpW848Kzq6wXwYTkXQVPyY+2K4hQZjGm6b/
Z8hA8oca3YgplFtR/LW155bfqiWsx/IT/Y7L8gVUrzP7GXrBbpgMah7h5hLA
CmftJtOoWiM87L0eIkH6unShBcb9mZYivgsXvig36ueQFKnD+gV82EbyK1c5
WsozHf5qJwArKPSIe5vORQ2mKVdEK1kYXNhOTp4IhAbFbS1HkIT2XgQnaUM6
auli1LA7u+sdUx0FNS7uTCt1Misg5NUMhkr28lrSx2Uglw2L5L/3NNz2IbMQ
r/Rr4G3XnfylUnHeHvcobmtbIKQefp4qOwuuiPD8ALlYrO3uqWcpf/GbSGIr
qqr3g0nQQHJx/MzVqY8GipQkyIwUZVvYJf/k5cfYPc/FKzrnzOTMotiwahSL
mS8PaUPFPDOenoIBM+T6lV+ZIuSot8wq9UY7QgeXJ6AX9egKfKGbn4VMx0jK
0VjGQvK4cwMt1/uBtJAUfpVZZDI8XvY+qWLBXLxTV2BEtaAo/VnWGEl7QbEU
vVwMOtv+JUg3fBmSdlP6aWYqJmk3lnor8rWqB8dKGmpFAEz+l5klMeQlndtW
D8fzIvGn+Obk5vWnoz38cNvFWjY3ClZ6yAfYpnRr62baMSeDlTcLR+3NuIhl
vGwLtyGBYuZPSq8mLqjjRZGQOtQd0AXPD0I+MdFt6kcS1+IU/zbXd2CyQt3O
gid8xoLHzrgUzSF+tkoRycFW2oY1PzUewqSvCAjRPJ3xOevksAjAC0o/izGc
iTbywXdaklfS845HWdhIycWIykNaP8zlrBk5b6MaDXhMPFyNm1msZ5Asy5kk
5vPMWgk1Hp1o4o200kcDJ1uOvf/gLcBK/7I7Ozajk4/1qfUGDj3orc77Gt6p
Bvm9K8AhWDiMs6c7hZq36l3evUtL5EDUjYBRI0+XVL6FirCGTR5bTKBQYG5M
7ly1xBKTXcwQ3QLQ6XYN2nWjc857nOdlK4FgCzxRGc3M3t8QqR1cOqoonSrq
X1SEfhv2LHM8TcF7TOTzx+Pi/oOWV/5vN3mLUQofqyEW0d1egNIuXHO0eanq
cdf0elD8uICQSt1/FSvGyw4NwhWWwsA9ZZbGITh+tnfq8vBzG0nwizGQmsHF
j3T+pXRf3MsCbFM94nmoDRZ0VOI2MoApupAKMdE/xdR8m77S4ZEn2zfR8oPU
qp+Le0jV/vr/cIrCAgtb/SiaoZW0sQMp/zEea9qU9bNRfVuYwPypGvRRa2a3
IDS3x90nYgL/QEDWikqRW4PymaT5oIIkxfkBYxg9LnFu0tgwIB4RONbJYDcM
c07D/j7F0r9x2cXVEmHOGt66BLIbtWoM9+mXFq/Tgg70uxxzQdNwkGbzkbfu
RzxOea3iZTrKFSboqs+iXqenNyg5RCfVUBFVn9/tGHytCfvkMFh5pDrYORQS
HPowP3iIHWOzA0qidSBAqRcFoM+6Y+dIInEvqtjVUS3bv3UZuzSFQohEw8N5
bMo2ivqISitXeLawnY3PFXQD0T91tAiijby9WVTc1AtupfdeKO7meveKw78W
8adEaeHwhuiRVkxyBbhABobQcv5qDgdYZocgpqYYwinD3Fp8ZIrwejNRKnZK
s5dsSk87eny+7Ck3qyzBNZbpYXAYepjz23podwbkq/OzQ9KISPyO6kZbG35T
v/FOECbsmYK7hUlxPRvAxg0Q++wyfb+LP9Kbl7dFx4audo7zqLrOUlAiRRsZ
rK8ZdcOELd8Z2NdHI/U8Jqqv/RvPsrpL1tgmMErnujVwWiBlLnEBSv8e/vxj
CYiED3oF5mvBIRR0dpy/ANwQnYmBOjVRqvkjyNyJ9Qo6o9J2Cq7dXQECV9ev
zmWZmVIMoIcRh1dfGD7MDXmnLwthBZun+5eusQy41oVxZaboKOzsuz5hgiJE
3sqGkavpb8Q7IBPfaE5Cd2YscOL77RDlolAnVo+zZwVMX/zbUaOEGDqZMXBD
o0/oXNCqD+u8fmMrRhNHZmtsTItXAnxok1+PriaVAUKu15q6hIvMc/OwkZU1
c9MLAZ3Xv4V5Ormd+N96jTwmMTL6X5hhWNeHmdHrTZ/voT7ZoW+NBXLRTZ/A
7Iw6K5WOQtHrPIsY1cI4DKsW3bS+/9WfZjnfshqZWd+6rwNm3zgpAwafSuwY
jdYw++M8CUcvJRdvCXXNPLhH1ol0XuPf0YVDyp4y0sR8jU9rZJxT7mlsdVs4
mCf2Ia4ckiF6jwJqrWbk5F4W3WDODaBhy5ocKp3z6LDVZ8v3OHpDwgWrnGUS
Cc2dAfRb/fyfPZ19u8Qi68Gwthex/WNhlTr/la9KYm/OSqMqKXh6DeyuzYfl
j9n61K4LUiFC0gWC2C8UQ2k3v5019+6pt3s75DQoeSdSKqKo6w00T1wcvfR8
vMfIA8oqOB1dUAky8hT5TZQ0kVtnIDGHqpygJNAPbAWAxUQlGARj7yN+4hNb
PkO9LvTT5X2bnfNgytRyW0j1vknqdl10z/odNMJvZa+0nrUorY19P48npit+
sXPRb+QETAM9LF4+RFcprb7owxWpOmlMxnF7R/4m75vB3t647D7cNfA7OQJi
6YDd0y1iQsDfESO5q0xPirSbS/4rR2PvIYoIT6OsJJM82bWqR5FWn9S9VgVv
T1Kr5aJIYV3pD0b6+ewRAUN9iKxqh5KSaKWtr0N9QwF9pdqGiqM3ljXBpLl5
zEkqq7NE5u46HaVAl6lXJM91LgLAwtQRGND7pIKXn8difxg5oZ0zJwa/Eepv
DRq4O4tgfPP7j6By/Mdg956L/pGqNsbR6c4qIFQ+fW4N9bYZTGbgbMbrY6VE
QoA1gGfFLrJyQquPVAeVQc2/+7kwLBT9r3YfGojURucgz5XyethqavHKeY7D
g8Aj1mli6Jr7vEn9K7zVUKylz7hzj0zlCnoltEdswuF8ROIsd9EeaYxcFXin
wMTNy7aUqfyrB4y7WH6u2y4858Hkd/gHo2vv9Vvs3l36w6jpANh2A1HalOHX
+w1myzSJH7X3ECsBhsmD+caIrDne/o583tJFy96pMUteC8ukIFbPyDMUrCXQ
CNej4tC4woygEUi+QR1dQ89IUXYMTX3qrDHYHLD10P1pheWOVkTW6ENQYE5C
L/DXKq7zGkQAlpqtqWXDP+RYtR7N8LF8NZrTW471z/gJSEDxfa9izDzklrj5
2bKB+frBZp513FeB1cjdtfkxgbG4+Y5TgLeoE3TK3Rn88sF/Vwgdk9sdl7fy
LwjtpMZs+CeDpxsMQ2SOP48D5FRFOhUn4ZfBOU/S6/fiHFYxgylghP9DWELI
WVvMSze0D/4iJaKubn78GVF7LIMRT3hehKDLR5mkoswHFYhIVmknBTVw7wP3
4FROHafrGWQN45H9nmkPDWVPWc068jqutSjJd5/Qs18Nxb9u3OPMVaK3qbkS
C+V+akfmSxEivWmFUGGp69F+Vrw2swNbe6zYFQEPtfSs6i/gkCdJYY7ByKuh
OUHcfnTpGPZUaDJGiNhNoar98uFMWoId3GksSljSzYtkWMLR2gF4bw9ltdgv
Ol2PH9jxGV8U6aXf5k1N49RW+R0SDS+HrrWQhkU4qUC8toG4lxqDOlKdan64
YBzO1GJ45j0j8KJkzC33KeyzRp47sPsbszAQYZ4jOBuA3S/hshpPJQ3dDbjF
goi2DPEm6rQA9LG+RmqGaMJW2dhCsFIV/MwAII9AXi4+tXFERXI2n8UFOjQX
IV7scfZbAOnbqRyS5EUakzFxqbPQYwcd3RCdZVh9PwJejPdNnushdk2agmnE
3oBiTCBkWPq/ouHXw/Kma5vqGU3bF59Ts9OXHAD8uhQNJUm/Qr2C8KiTKz6K
ABV+rNQ6rMy+TavjNn45Q0qXlqVA4D/XDsBQ/mb9/ctt76LWpZgsXkix8x0d
IisrycyPhR7qleNI7AHGWB5DrYlomNLQVstF2C5rKghzPYKzlAT4YJZUTj8O
+uAVUCybtX53UyjU0bUtxT+c0Z7Z3tq6diWf97VvlHth/HykGGTmHB/zxYMh
4uSS54GSnPhcoSGgu06MWuXCo7Rms4zwnuyYiJOEv6V6l6fQdjkgh9zsjoJI
MgxAT1UQjkSExgUz9wv1jpSbrV8DV4VFpNUpRu/bY6PEQPHzD5xkqGSUcFue
iQiZ547pO0BWrgGvH+pfRMZPtKlFInQ6xlvGV/MBh71rT7FS9n8NwSfYwbG4
xqMWR/xG+QKuJFzqPyqaeV1n8llCLl2pvugLtiBqtkHCBs49BnEELWQMUn6O
YFdJ/lQbz9sMU+6uDTQOU0XRSTy4b7x7+PKMmQZrFX4joXB+xzAH9oIBFy85
eWsWCWeDNhfMy8YylU6gtHX8uF7HeiZHSzMSfXSAKRM5RQ54Bt3KrwEv27QY
oo+i80CI2dzaUnlPp2UfUe+3oZfG8G6ra/rFRydp1DfHd4w7knkQ+RrIsLg/
15J8GMyOs7H08iI28J9e6qCloSv3GY5DdtvFqUktG0A2RoSQkT9HH3NYSWSZ
sUFWe94OFj4cfNz/qM1xQVcQ7Ifp+L3SuBsx0LY3Vf/vGow0dBa59u8NmfMi
XMvqJD1M0VHZ2mUKSAe/pDIxaAbbSA8ttLuIehcc6tvwsCazx7N0+4MORlwq
GKO2x0XhIfWxNZ8C0gdzO+jajJb9JNF3q0EzVjd0XszYpOrEIWI6I6uN2qH5
WGINXM8L79OMdmLu5yYCLhh/seeEGPcvL2x5c5B0lS3FP1GqBkQ/0Z8YGK0j
oFEp37lCjtv8NVNIz3VznNt+OKpzXGyffEn9Ipc3zfpuHMzu64sFut09vMdh
Jg4Eco+eubIZCwAVGOxlczgoOeGsAssX88N0/blLJNDB4nzXudjCCT1f9KT/
cHimHiMSHZIt0zz/wFo5tFMpu5rMrvK/MzzQS0Gph9jBhOrehHWhzos56MbH
p/8UQc6MUwTt9IwV5E1ljQqj6/QavCtDuEInSXjB73ZZVFGis7d9ZRPhklYQ
qmhJj7PF+uJOWkna6QWdc9xDyj6mp82RujfHnQ3kxCgEMDcDNBN7HDgr6PRT
ok/BtEe7IlevGAEj5qw9+3anfeBnG3Phv54OlRc1P7ZrDJX7wA8WJhTdGSqd
JPX2tnlHQlexcryThlGSoS6QfstGURZ6yW3qpXkmjoaedodMsnyRWqTYNOE1
cYgmqWtplNmVCOTobjtzHBxABruQpzNs/h2QU1vxOW85rO/ADfMktPhHOEdc
FxHqFuEngCBEiRlteFPckSOTpxoS9Y8dsm0keNKlXzR67TqsbjGePnKNUG9k
UnB3Fnw3EXE25g7dR1L+a/rNgLuVNpRZ3p9HxY3/KqXR6JW0zDQ/UBvujDMh
fhD0SebPs0os3gs1sKJrrFA4gr4Mn+7h40w7uERy9G3h18siEaVVL9eUaL8k
JAaCn3/UZWYvlR3oXoSJEOWm0JOJ1HoLaU741M0aygyMvj2mqLG9d84Rm0G+
uegswMY+adsMciYuQYrZ8jlD5CQ0Zq405Uu3hRbXB0qJfjveBJhKNjNZyRqm
ZwBB4XP3VS220bSNhHeHusS5k5ulFyLm01+x3F8uEjO5js027Co+7Y7HRt2S
mGsk/lU6nikwkBQwf/tF39IuY4BWcO7BJf35noAX+c6zXqWJGCZa5KaDHx2i
Ne8BNx08ykqzGrqUnD/Rxpl38wjgir2X1eBpts0etAP03QlqFCitJF7lJvnn
8HV9R9Kfmul4vD5JqFs23l/jZHqVXZKQK0tk+MYPumO16Mveblu7GuLBTwH6
BtbmV0wXH2vSU8WCIK1kTI+PvWaev4b97YvWLbKiH1hgnVdap5FU1Hxe6PHG
M5w9VpOnssHQj6Qbmo6pZnir04K7PZnxZVNjKXMkeu8ew1yqNoLMIFYMuP4C
WGIc8ZH0azsjZKYAxL7zT0NchkQDLkKncDPOvEsbWUzhxUkrDLv1XrjH0QHK
wvjEC/qVtsS8ZsJnmFjRnQO/4sbxDsyvjohS7DKSxlRGIGb5NNTl8RrXc4uA
nypIaX7mSyVAdr9/7EtqLq3kP23tPeFyFpuVqxTuTrUQtWiooPj9P7RjtG+k
q62TUQK/OtfdO9cN0eQo9McJSegSvf/fpkyUBpS/enaorl8HFDqXJw5xH7j3
bOkofMtxskcWqwkdw7aBzEfGDMHAuCRtNKcB0xY28C2CWidYc0XAvJ2q2Hoc
WEpMCnp6/K9rCM+Bcn0tajK/jcV7HymvtkBavi1Jwhid34SAEmXckCuXpYVR
mbp5ECF0/4ZtqnFypUNPWOPqP96FwbyqaErYYEB5YNGtPhcQTCP98hvjJKSc
ZbTWxkgGSzXTWt5EWjeUKViJo5bosjkfxXcvHUFNt+6G2lQhaiuOgoGEz9cM
ZW3pzb4aVKifhhyiv+oWRmHguwCwNuMSGE7Bd4a8Xr2kgeL1RxFXLAbk1Rwx
adNV2jjvWY/GDr7yDOTuX5kUzjyT+rf58wdO39req/bDr+RdVfqP2X9uBkwy
xsUgqKiOgHEJ1awi79p8DxcAtr4vPPEYN41ACohBavLbt3MrcJ43w+iuhly1
5yhisPSRhwWEbAiLnMN9Hw8adbbsPLMIJy7dRySSDfJzmh+XdkUpS1pPhcHG
SQ9LiWQtmBlBLnjtKvjhR+v2QkmWzxLlYikvXB26D6jnQNyoairyCqL+1fd9
bTm9GsEug9ZaHiBE74WGx5FP6Y3Hp+Zrn6QThNikU/xg7w1DbxLGKTUh5cWM
aLLodTURlvvzKje0TNRAxDHhzQQrK5xj5EMKh9twj9DRBM5RUt7bCUMEZ5ko
ysh/MHJP20QYezAXi7Xd+iWRVb+NoF1qT+9/nOrdrWAY3LVhj78lYJoHQfxo
L3KXsqVqpTxJWP8RhjY1iHdYyfpv1V+qgoBgxNyBfSDDi30j43hJ2s2dSeli
4w61dRFEsBKxzRYxSe4iqdby5uPg2l87jAQ6Avrcar8AR9D5XuAVBSpj4WeD
yy/zXSkyYScajbK+fi4rClO0f1q37NUPNXryKh166ykKf8AkPjCXY5YkeLxq
j+Ag+cfw7bSjSkFxoED448sjpWzZSj/2UEg32e4km3108HqXquMi/yh0LVna
XVkF5ZPdrXg5FPS0OnWgYxDtHsAgjOsyNGgyrenGrkH8QatIUhOtabh9VW+/
9NTZu6UHPa4KooDYN5QeCWnyboxNAytu1g0PDOCM4SbAVh8l+eVTq0rxQLJ3
vD8B4zXc+5A/iLuQ0jXmqu77HDn6zBNbfQHGlor+UvTchdCiDKJpWSV5vAet
lSQK7sLxDFz683yIUk27znWFcODxBew6NdBgBC9Tl8okQsmwkAQxTFnCut/x
fJA0LaeUlGLqlgfNHc/BQt4vnj7bs04XmqtePLe2F03WMmxMVKnPG40I0a+n
E9pb7ONSp3LLxFyB5vaCOv9T4tbQGD2ThM+rxJUJIDPWCRi15VQ24hXxtgcr
+BdWk6TsoRa5MNTv15SGdI3YuTl0u4sikwhUI8fLPa5+6hwaDvuSxBFtX0n8
nCWkL4DBFDDFWm5zmMSTc/O4W/FBErfbrlwLzsEMNxb1iLyu3QQmVW0PGqAo
JbZD5OqG8AhRCLoTiNYvvY5MxNdu9SVhGBwy+QarEqZ3+QFHhbngj5/u1lNe
T1JgollexBPLdKIBr/2H8pRUBRWi/xaABOr6KPLP/vmUrl8xX85H/gI288Z6
g0bdYzDqd7vsupnSF4ekjr50fDFSvpOWLfGEwBVR5UocayYfymvKYwllJ6Sb
Pg739bzTWY+SQ9NQ1vrBM5eajiRNdSzHh8SVe5aG7NSYKh3TxmOatFcIV1VG
G9NjjIE06o8QvxwSc/jj/fYyuYOWQl4yGQnItOd4n8/mCEsscJWJ2Wah9AyM
QFBKTgxSOmHlPEGY5t2TaThFT8Tpi+UL2PyksrLZFh62RU1n4piYcn7wAi/j
IG8FrRE7By8stzKVQAU+s5BbaxD+NPPkhtWLmnmEDPYoYmR+G8sQLDnUWnTP
GMgY2obozr5U5/4JGp6q+GAavIXcT99+sIHKM6N/CMRPSSCsx80V5dhzsOLT
z7WQZ52izBSr/6EE8n1nkEUoW1JD450hT60wzaqFw4Y7DfhgNBF5E/p8uhZr
R5GlCB0p4j3UwHhPYC8/k39q7RqXlFQCCUByUCZIvUd5lxS8YF6fdyHgOv/W
1ig5Hs/X2AmeJ6/hBG3V0pEgoqrbmnwzpiRsVL7No1vo/NGaQskc1RuMR50S
iopyJEbQtKt3JSnB8JlMfBpPXolwwnujYcWL/4Q2FQmMjra9aRPvmGhR1Uxx
yiPADd1JFZgHG4n0vk5C0SIOvsG4ASRVYft0zkklbfITDurFq7QuvtwtujDx
eCz7vzUNQYt/JGnc4NAWaKnXi6oz/2QPxiR+efrWjiq1AYm2MFDreTRxZw9r
tLCzOLnnt5rUvxB2wVr9yAZABqpmAI8MGt9DcbxKEiSbWumrs77zQNvD7ncs
rKNXGTF4bsSy2O13iprJP92DggAc+Act4TjhX5LKnZlzZaRjoKDTunaFKIYN
IOYIY8ucobBn2b7iufZYk5GynwbWNLI48C2sJYJhdFuBW68FfUSDhi2ZwStA
tdcz4vF1mP6Y/Gzf+D5IFZZ7HhS5MZM3AKYXb/RaXE/hiHHmlo8/0kAWrjcT
sZnqN7QZolxqxR2wANj/+oZhiHEFVn2JqS4Nx9gGI8wskM9l4BVjESnOKYb6
6aOCM9DbKM0Nh6p1j9b+pjABSC43eQ5vsPdBwro0gQh3aSr2F4C/9G4j6vAx
qaINUSpfAEctUZgpulEgAeisqiLXZQgNIE1oldDmJGvEQiQh1uYH/C9O2D3M
MbmjWfMrU1AWwnl5joqCPqjbiyPxp3nKfIZvkn1TVS2easH8R0W7YxNhFTjF
jw1ZRah7lZ177nbd4BkouzGc/1Cd23saKBigeAF6FvgAsAoEhhg+hyCAQ2Ko
6zPAblXxiWSuJbjL5WIrKyT2OtAPTawCVP9mXinqiJ0EiZ75G13QRfEmmjR2
yPR6X4fKYhB8mMvwxZeClHKkGtn+KQ0+mIrm+fgSPcVBuofYhGAmvLAfebtC
SlnowjQ1MXIAIYreLyLtIp53apoiDihjyU+AhQZeWgbAwKnYvhTkncCkoUIl
Hm82Qx1OS92EcqNt8RpN0TNsHkglT1wmGo5nqzHP9a+ncbCpRvjxG8V08+1V
VPXZxJgnz+KOu2XD5d+vfE5NakDMsZolcx5YyRA0HmpcP+jewlhapHEXjPTn
cNY1KY3cjrRss7ayVkB95IjYk8DbCkrbENXnCiA7WVZhHOoI0U1b++XqcNm7
MPaCExzHwqzSUbE66x+yYiSrgW3l3Onc8qCYeBfVVaoG5C5BDuj3AJwx5xUf
WRkxSJnQEbfqG+axTh1EwTe5m2huLIMYTcCGVnp3NUze/uppXKj7ROAn2+7l
pHf41g+f4WNv3SVZl8AzXu6cxHocp873KdgYC/iWWvtpHgGiPQDG3Go1mcKC
ws2sl2L6pEfz3Rblp0rLrRATeC+IbI6jIkmHr+QNXeKHVkqtk/yl7A8VLm1/
ruLjMfvEFbCT4vivfjr4Vqn3lV8XL1odT6L5GozTqIWvf7ITgMAP2N5dfTQl
ZbjsLzLJB1XHfHAz4irj4Ka/qmPufF8GO6drrBT6ousA7mOP9FIO4g5RHn+X
8+SA7JmnUi7Z+zNMuVI8MV0JtDaBsm8KTxbwfH2xTwnWvNFS2/pAC/SEhhY8
AmguMRGAsuN4kOKwhawCmpCQ96Bb6dteyh3nTNG6i+2+8WR8Fg8R3UvBGxdc
+aXQxLVBF1zVMyrCc1/tHa5fMFGCs+7GYmTkLe6lC3Krp6CDpA/Y9rdPmVts
fvKIUmvZNrjop5/xYEZqyMazaRcSPg8DPtfr/oyxY1R+T7zLnnjRv4GrODmK
Zr5EgjZHGcOliic1bVcAPpcPD1OYOh6P6mdBP6opA+vsDdEBquR6UH8KRKPd
HF2vzZ2fgDNvNxBjNehzrzq43c50vrpvzMVvq5iHPvowoERieFtnGRAjzGrl
Tb7T1RVNO12nPkeNk3YscXICNmr+xhZf90hBvHpH4woHoyVHVWfmTXjXyEEw
hMbGQvDJChSq31ZMEYPQKIvLkwIzd92JUw97bzEHu16XyJhg/ckiSDs5D/jH
8Wk9S8d17T3g4jcba3YPx6KDJ6IMbfPXugi+ByEsV9aycmZPebqMHwIS03T6
vc1+8Bx0r/61MogWkJstGpyxZWVtLPf/NXYQ0+31ZVtO67ayb2Ks9ww8MqcF
DFysjgrQP0jafX4CnaImXWWiGr0fAWBYbICYdGbViVyUunDFjmo5vQ2ZJiC7
7JYRHLlH9yg4kP7fngT7jFE3WG4oJ552GA7y/s1HcO9jvQYGKq4a+QLY5dSW
ENgmJdE8DFUf6z1ahLASxp/sRieEi50eyTEP5TXhchM8Haw6asl+NrwkqqyX
vUsQFfmn1tbcetjZ4yoeK3etI2tLIy9ccgYVxrug5ljKXdGBpE+Vt7B705lZ
Ecqnz2DBAhI30ogSRvNDfGj8/8DCT8sSEktvqtv9vrDOzkq0ByKzzLD8AZ5E
MMqo2EmJGi07fAmBnxRjL1J230KvLOY7Qx1zl38VT/VM1qsq9jbzAvhLsIpV
u+NHyUOYPj5hXec1qkuG3PZ4s0607VXnxEqQVxa60n38FqBICc/nn817Kh5W
O8mM2U+T94XrQW6RRfr4SWxsxj5s/9NZOiFbOiE+5EMPXlCf68SCgcGGlQmM
VzxYWlsXKBKtIf1q9gxnaQPeQ7sbnnBMgjjV37sKMVamy0MY1pCy7fiHgpqP
X8lCItV1Zql5kMMHzXAry/6BX/myHcL1PkjjHahwep3d1uJb4nlGqMiiU8nT
DBwPFoz2zd/AG2Cov9RS8p96n/Uf5WnoTJTzCHPYV9QLqL9j9gX24ItKhKcd
m0F3nFfvIiJJtz3MWlZWb4KLvC/2MMbyIo635NKUWfDBJgVIukDRTZ4R9+29
ejZ2n/P9tA+nFY4sil6ljg2gvymJxvT26v0JD1hsTs1XbIC3szmZSama4IPP
oyLxPK5tqK61eUpWiDwefnl6ihCXzx9lcB+MpA3qENL3YiFrIUrnTXmCGptf
DKAf7a5c/iYZDIF67VEVqdCW6SMI7uQuysl6kbm62VgKlfZsYBqHYeb8OLix
ZPmgizjYHggydZj2wGoC1FH1RqRKbXPw3yZmTU59n3N2pu8HiwSS1yiaOHM1
y1VPFSjKCX4eI3iDJf8r9wYQTk/elYXEWow32o4kJMB0IH9Qjmjn52qTD+qT
4R6b+VBgq2dhE4ZLwOUXwaz8JPdczsaWE8boPVrxbW+raw1mf3PzvpAG2SmD
0cObHX5Gs2WcyaZRgwkw9AGjhdGwbSTtze2t/rNHPrDEziDkp9UqrGwNdYly
g7hqhUvvpW3vL4Hh9ajT5Lz8Ar3BXPCaHYsg0C/2XOoPa7M2BTiSilA5HxnE
/UMiBtLxiuNRtYr3tFZ+mp+AFmoZeWTQl/hlPYjby67WzQ0W4yPIakLDo6kM
xL2xPXSZUHi7iX5NJ4fvv6JfenenoZeoo3kvSso5XwXDLKf8wAl8eK6MkcSA
BH9H3gVcub8L7aNGv9nL07Z+gSYoQuq4o8xokaayhoSw/qGlGCI1JziTUcQQ
AykoR/wBv47Yw634NX7t8L8t+Fs9JaLz9iHiIqHBaPJkx15TDnVWYUCfbXzH
3uBTwj7qe3/JX57vUjYShPZzqCZIF1/oHXK3xp83G3CdNomObjj6qE4h4ABD
oDiib8N/KetiCsiQr+/EHRd0HVrUwCG0L1Ig2uYlclgOhHBscnk8ukSRTLTo
7CMIJbI/4r73CezPqZ17T+hxdlzH0pfmr0trJiHSmFdDuodb1HxtUckMyi3l
u7cdO/UAxtNVhG4K+LnPngWVjDtlHM/w6w2/eSNfYxUu0D1xhnLwS7pGaADX
eUCEbn+8g8HhJgAvIRiAHlroiLL7H2LJR3nIreV7aEd1gNJ/5D1ainTMDDFg
/xLyLryygS5N9ob+QML29h979lZA0ReuOEmw1EpUto8axrQQ4YMp9R4odqAR
vCdYEzUKgzRkfCnTMcmU33vJ8+x/qhl22OdvFbU6m6R3246hMYJDlSdlrfvs
R6pYptxGlt/8YiNU1w5dmL2xsJKnGflGoJdkgRnmRn68E1oyVWZIc2Qpnozu
3HHA1/0GPXYmtFPd3nQgkMsj2lLBerCIhYZ8I01Of3UmhUQ/se1CRVrtKYCx
caVuQTj0cGHCKgMgu8ClZ2z0Kj1KVkSO+eGpjllT1YlvRKwjz/etN4jzUIVJ
ZEubIzZwns2UBv7rApzrB8H2p3y9+LWy0yb5OqYD2sE4sOIL4k1PljOO6GhU
wpdOvxlK3ClfRNNqjbnpavz+ke0fiAyaHqeGHsv4cL7BtlMiQQ3Ns1WiezVE
TvK798qMIGjnJQScve5kjBNjw4y+l5db/UPeWQOm4+4RTj4FhUt521A/HXs8
J2P0WrZYPE9z0IdMsj1YjGRJujj5qyrgdHspDz/98sZ04m7noIyMkQnyC7G3
Ntuo5pNMbvzGNxjcCEtWmd/eYN6QE99sLuzFfns2YGNIT6gZMCnQ22+rh3L/
pyIk/Fk3ajenWJG56bj7Glxh8Uw6/BQLIpF2dm8h4gW0+UPfYMDPmZPcNq7i
IvPocu4Lhg3//RfGT/W19z6+e4Rko+Dbq8d6d7hLqnIMKzd/CMWcozotPAYY
lVpEvXPuykoM9khj0x2dvhp9ITeJ23GxVZa05h1W4LSXfl+VMraMktn6Oboa
Cbb8HCwAtH7yz+LSBnaOgrJn866X/9uyEwcwOaswv4tK1UbHrzQrAiO+6bAx
GtBcZpk1IqoewI5w/tNyScfKp2lHlAoiJkJ3WWzip0N3CY1fX9RqQv1Qn/Pe
QIHkmqzXxEy0H+ZbLq7uGf8LpfTfAC5oGjxtTT/tBzfv1jjq/6QRSOKzS0Lz
QHk1yQZnU9+54B17gVL8Ujru3o+jXxxBS/flR4c6z2qNc+ogErE3Skt1O5NW
d9V1WnZAgDYj0vIUG0GssYxsAPyv8M0tvg3tKou3R866HEc6RdkJ4QG1rlDg
yQwDGKnvKNcIi64C/bDt0X+aLikoORgg/FMR1qarddU2yUodkq9slDvXd4qm
3TXpwKm3wj4Z61PgpFgw+9+XZJfspAVJjlHmz7altrq/uCbLMIJQBLJByiWj
rKLevYOVpuf9CnbkI9YtVYhwXB2yRXGSfiOjmRiVNGYvJHE3VhVJ65H40tis
mzNExkgu4o7m8zxl3Gw/Yt3uxGM1ySkm9qaBtL8vd6c3UwQQ66N7wS+EaAlR
pH8hspn0155mKVTqu9sGfl6XSiVUMsLtE6BQbWp6xt2ux1LzUf17ZC+bG6Ve
0n7M7pFxZnwLutojGckxD2F5v6dxMSPESfBoVWe8K4wPfeGT4J0KTqf4SwQq
kIOUEt5EcEhEIM0Ho12Dn7j5DgK7KI9/SzmdTpyeLKh/pguxT/jkqcOGN6Me
/ARLjPD6/M6A+lo3J5slVYxfcogkTKXr1Y1l7OKJ0Zet/6yERTL1KK6Ta2+z
0RYCArYDWR1U20m4nWvWi1Wv2hJ28j/ORfgKds+vmVye6UVKvdU9LK/2/kCq
xNO74/rw3Bsqynq7vbuy8+z8bPbQYGrf+VJO4Rvk5U5PfT6H8g8r6goKMyM8
qoIxElZLR2mrjOePCNnZcL+jecy/iL+HUo6VdCKn3p48A+xvo7RIPw40VNqL
zAz9kU8VNKUdvDJK3rlH6mIJDo3ak7eyP+GSIt4UcoD55J1zDhtZkunSTzJl
MJFGzCsV422mj7bc+xSIuZSc9aa0A/KHm12EI3vk1ryyBRvcUyHVZZUQZmjD
O7JNnCm4xGD+mw5Ud+icHk914EwQjuqfFQPTnjUCV+KgyJ5YmBV9gJh2g9OE
oACxMF5PnEMePWWT70BUP//st9dY5JOX670bTnv8uasPp4Xo9hxqbw5mxMfY
q2/dKcaKv0vIUJfM1QplvY/gxMKTh9gr1z109FoiJUEaHGVpMKIO5VSJrNNu
CqhKwrEMObOtAz+yKoy9fvUsU3pRrchen7F61stjCxefiMOKklB1+TVF6L18
JoKpwD2AeIKcW8tmgB3SuFFNbSnOQtVByGNOwsdsTF/ZHRymUp+O0fQfnjiH
d5hZkH1Y/gLMoeKTQEdjrIb93DtJnKSUnukOAryqPutgGHXQAAIw8RAfBG4+
oL+i++UD0PPlUa7XTlIkUBUVeOuvduftfbO4FB/Ok6LDnXa/TukHbHBdpIpX
sEGNODQuk5soj6apW+MWz5Gc+2x0LmU3XAj3f7nPOYPFHqaPjObbHefu/nqL
5j0D+75ZSppas1vGZ5pMQvLr/l2Tz/BapIh8N57OIRuk37YBNcQMny9dSUqd
H1wgAhGlkvE8/x3I0Jr7Mu6CFpbcChrELwUvEtWcuz005RxWu/ZbHz9CcxwQ
kmPbPU35akcrQ+niJmI/FOq0mj0ZzLcvtqxA4yd3NqxgUZUaR1bY9XnEPSzt
JgK04gBZPIfizSuDZ4XAC5VA9UZJWraUI64gNp4txaQ9iLhL9Cuz333YxNAh
16P4rZuD/bW7qcPn1IXZhhPtH22SZoIE9VL983gZphyZET7SWpaUhuy/CFY9
CFEdm5F5f0zwdXiGMwWKdmix9kksBLz8/bJSWoaoK9h9Q/HQgLT+TQOrMUXt
Nu8SuAW0zFnLkbgBbSXnkDSkTRRO3XlJmSL0Wj3sSV4nmNebrBztkHIwcKGN
c9ydBQUc+lf+T18Q/nFHye/zMsbqtc9QenB5Gp7uEKC9G9diqVlkS5jR1pmM
rHhf7iWPzFaHS6lpSw8+f4tdnCfuAgl70x8IrFs/lTe1zHVXlebGfCVMiL+o
yoeF/OPq4vlK6qYMUPncUhDASzsiE7JP/eyLMg49zJqwaJ9aV+dJQMJecz5P
XIEXIAIiqtGF2EBNOS5I4VXe0dQC8Zc09xo6eo7G4vvDIjijaGmG14MOMXC/
9WSuTy2o4l3/WuLzovtzKo861EdbPo1hPK8soCnuATIpsNRBcFLdN27hFpCz
WbFt32sXmuJ/DhgVZLqxhkZkWoIudlzd89yJvJjdHqu77OeX1qbnEIqJvctK
+cMYgt9spuDw/dpik+bvgh2BVyghKkKe0JZpleICFqQJ0Ljv9VrMMJr3Thb7
4RwsiytMsEXlh7EJpguhcvMfbULKxUcT5/R7agfz5+brYOkR6cG8OMGQqJgv
oTwvbuH4FEbONyh4sNeIaxHg5kDOiQjHbtvDmzJK/5/vFpl0Erx3Gp38SimV
aHVhM5p9g0S3FHjro17Yti08300xWeXxg84RaXVTPHB1FMlcaFdZcTfW4fix
EU/u3xF9K/LOe6QKWGcviZssnmfJHFvjaK/vZUfrEpLXeuAXVLGdVjpx6Ff8
IMwPwGdCTfYa9vo9o/F02uQE0k05C2nIalKznsiLkqsU/BIcB399+YmvtkRi
RTWMDk+lZJRLBX1eY9gERweSRWTKt9PE/0pcRSYjiehJfHc7LoXI9knGkPtm
0TetIAommzDCLzMl0YFOpeJ3eNzwCL/XijMZfeY7Dwib0xiBhAU9ikK7rNWR
4j4I4P5BsnuTU2/cyZ5FR3PZcZdHxz9B9u0+FVrwv7h6UGaV1XJ6DlfKvWvg
AYMvd8ZQBy9nR9v3ZBKtzZ3/tEXkLZFojfE/K+mi5w56qBx/SRlHXlfXdWie
iutewEdnpxGxKhGrIJNdcruYbZ0gIWkVgoaMgrpKlhjSUyyqAwnI/7u23iSB
gs09mdyA/e47IhnlcxJ0bgar3oDwgYikauydAv+ufDp6YxudS7BeriR8lsrI
WwaoW8WD8lmTC4KDoPQ78bbPe+gyarnc12YHFPXxbAr1QOGUoiQfRwGCWy6Z
A6lPKaaaEAbWrQxJJXgRWWrKsg1SVR1r9SUVmdXY5n+nkJlYhvfYwOpA4lip
U3JB8ZQg6K8JYzRgCEueDkj3srxlwcdwNqMEnaMuXNBOV5+2ZXzG5E7ZqEoG
XZ9o0KK+G9cstAxz2CrMwfwuktDz5KsPBdVdXGGzaw7jR3gPQzwd8w5f3ujq
1qtVEm0gfg3XkUB40RiIGzNm3qcm6wagCQ19y9LxOrC7mRPjkQV/WPt69Zd+
2VYz6gPHHHhkmTs6zxCtpwtO9241HUh8wU5AofQ3b4tK4CvN6mNA1Z5LdPHI
8ppXLba/IO4fMrumQsfJ51hS0WCf+gDufgY5upOL2OLTWnVkqFMQ1GMrjZvz
hfvoLhT4gNTIZtka8E8J8ASZsYRTMah364OhdgiDfnnN718+vgNwNfXYXRlU
aA5dLQOfxgNHi/QE6yRWlQPHvo2Z0avkimin9elgzdAh+fzrPCviyGnfDOe4
ILLjzaR9yTEJ3gKlCoYiCHxo8L//gUatUz/pQVgQOmwYQ9X50OV71ZThqLX3
HHwkN54wk72k7jEdOYtuFdyWQeJnmg0t0dS66SwtBR90P+LXgpw8vQHCll3U
Hq3F0+z098W6ff4gQRF1XqAHuI2B3rNkacs1ofKIQcXNTzWBUhh8Twnp/1n+
EzPzzuOAQXFa6LsnSzYs2IyM/nUiTQZa0szCuL9kJkxWHHB4sXxnfSsD1Ph3
LwWXQMkyUvxZbisGDp1wKrN1J5VosDAr+ezbydWlcIj/2dN+mhgSlgbgB0An
E/pjOsrYfkttA7xH8+3O1jn/ZaL2d+IGjwYIjt4WmZzBuHyY9gCglhzRK5W5
OjqjUgHNHsyxk8+X8UjowjFRbIYwSxeCB/eYN1S7Zuc9OBjAMwVeeJup5NuJ
qKDdc+JVozOhowE06jbh7gjqHMzLIwNXZ5ofraHTWaDv/rI8ST+WbBc9/OHA
mXjsFkJdszmhhcJsGqkFxDpVo20bIXX4HGn4JAVTJUE9A4hCnryn2vezwHb2
tYN4Ttg2Y+xWuC7LYT8nKUH3RHAXmQR9bljsaN91zGuVHV6YVAAHk3H2xPxw
UaDs0uL48hSCtIRHn48Bh+Me985Xd8Mrnmhlqv+lDLQBHj3S3T2pWbEXwXEv
J6fmnv6VvJKwEaHf5oCGX6QES6eCtlcOGEQuyc44EjZgxsaWREE/keXw/cY2
UbkbgpGVdsa+uAmNkFy54NWiDD9V4IANUkMAl+CJQO4JffBXpgCE/uwyb/rT
b7ATXSfh6bL6GTnculdnTtNEFrhf7ykHVKoBfdb/n8tBogJvwNS2mCO0quWq
6vzkJXjEHUEB1yn1USteXFIvFVmlfXKsNLpIX0ocGe9K6+NWrk1QJu9dYIzU
QsqeL5rA5qTY1to1zY+Hswf/00oXr22qYp9dtNcUMIGpi1hPLAuv6CjehAmq
ulefAGju4NlTCtUmyw3GRr1LiCKLdgz0boq8jxlvxFWYx6gxfx3h5JPkgiBO
qjsIO2Ys1AiHEfGXihm8omfyJj7fJRosSjKw6N/c0ZQr3bcNPPEInW0PaMcd
1rlkKIjwhzdsD5GVL84gnbt1+ogNYuiVTxUYeyPioZD3RispjN3Yg8C6rqIE
UzFc0Y7NTZm5/q1ZIGCBW/G5ujj1Fut6gLaLvxZuQHRrfaYEX5j9tGya6nQe
zvwsU0CafZMfaItawXWH1GjnCBCZTjFYwD6OCFDbntROYRGrBx34yM8sZU/U
XJLrXQ9jAl05un1jIjYjx5CnOsQenkqcv7SVMtFL1oxIepTN5xXwCIW0Qr7+
RDdok7I33k0NFly5tWQpVLdG9iMYLU+Xcu3LgucNryCXxLSlXZJGWiqla8IZ
MpoLFrCGXt0Y1e4iHtRmJpNK6vMy1+mwsrJfc2M/0tlODsumTbVUy2E6wWMh
8LUybnIfXofQKu1YI7B1N2G7Ogq1xV+LKPKgrUUJ1AKSbtMLyBNMXvEiShT3
H2okTwhLeYMExWMQ8zxyCYxEi5G9ptsyhRhVP2RWhLPPInhfU0RM8svIacBS
4sJzl/mOOHZn8A8SX3bZC6F89aDXUWmbrxYwI+ApPC9boOyUj8Arxpr0Ry7G
V0BRluVl5BNZF2zRCDfb4qtzXUjnd1EUVfxY94e80W6es6zk2dfc30n+UCN7
+AattsZflAcpwk21eDZ0iharjtuv4LzulFQOPlnrMDpF8eOpFtsGNjGkg+N3
pkn2NQX0sngLbuaPMLGnMEhB/d0kEKAsNfsTB87Jr2N2STdjvsyCN6rMgGuu
60Er47/CDYDcEtD1Z+lTvm/vwCqXq4k3aByrtd8RMgRp4VAwgtTdKyR5cHy4
UFyBbBl9pHVTtijHRmdFhm8myxP5mLirGwR9DdBjlYcy1pkoLqInw+7oXjeh
sLyXGsXeYJ+Ssrj0QSB4OMM40o71vJ7tsKupVu3aA7mRsS6cfKCPhkOglig1
Vqvelx4WmZnFU04RB9x7kdsNAcXitrplxWC3J3dHO1u4fEgO3ulyJTuQAN+K
L76bzoS6sEv1H2nKqyDEtmxD0NuEIJmnAc4QiDnh3emKSupYlLEsp0CUQfdN
fq90LWkBeNvwWWz7Q4E2s3SLP/KIfHbFFbduCzNpeE8Ts4cOQKEFuiBilpR8
B4BeDlBJzwi5Hqh2fgL+yZZKs9qQS44CbaFH1xZJmgKu+ModQCClU9BA0k9U
ls4jsvrJc1olbmh/pqagJmJwq2EhN8QI2A+2ec4Mp2kTE2GZNHkvy8UZOwde
U73o2swcV3lEq0YdpKHbvGCRr8SXC/CdFM9svkQdCOjgTeTnYyZLUAcsYc+x
I1HX8PZtkVEGXXTOJyMg6qWxw7SRf0AWKItHG2mDRnXrgSGthTUqNoBYp6uh
prls4sCX+2KRs08Gq0ePTywCaQHRLErfg8Y20bRzukGBe5/c9hFotf8Y7Rnh
uxPnYuFxXVRie9j+6bovaBkUa8wJ6Zn911gnwbDZWIRspf54+Ul2hlcFBlGq
jVmwaC7NkdBmrKV/D2tc4cRR4sB75xk1++pAnFtVsOncn6LPo5FNOK/D3Xz8
gruXY+uQcqp81IV/zTT3kHtPdc5ZSFFAMcg79zxO5CuVf2j/2FcBJB+F0BOM
49hemcNpLNuWIpgHuMSHLEREsgXLvfsBNWKLCIBjqdMcZu3J80EJrktazutc
bmHD3412Pib/BWqpmY5io8I5M7+c27iEYK61PU7ZjooT5GYg0oSlry8H5y/H
RK22IOdCroZXpflQNAcWX06ga+PJjj6ruUPEAULgCS25lnVsCDhNY5g1Zses
tuKsEY2NUEyDcQ5JOAIUKKGwMHqXjyqLh/Hv25YPD93QGhHbm8/NgFjuYUCS
9I4J/O/SsAdZmmlNJiFqCQur+tlXazRrp/fuhV0eZPd95SH5qfm4ShuBzijI
Shs6NYczD1+PJNh9BXigXvOhBy5x4YlOHlGEOwUOwzkcZdbgqDHVrhhpV/Lm
/jFsK4/6TCk49EtEDCJQ5d4SAFREWStcpEuxdJDNOiR1oI8LeoUDK/J1vewf
QiWfenLSA1fWqpEFbDvyExv7zc55bN7UKihmPHXQwCUNwBzBaAU1xjLkPQB3
g78CxqjVT2bjed9/oyRWPJmo7F+S1t9FcxHk9X+0UUjrOJVay217pUin9OJ8
o2ITp+VZf50QuxHH5GqJe+K+aFcjyMuBmQPTtsTJa5xgOayJ/YmAMqNb2LZq
kuAd0do442B4Exk+zCkuonaCLg3hn0LPzCUiSjw8R4FgdM6iKs9H00XP6Mui
afKdxZxl1+yzXPs9Sw+WVR6ECNdXZ2n4VnHEt4W8RvN+i1cWk4m4nNzypnDD
WLr+49CAYZFvxco3s3R4KNu26MeEBxj6leXw12ENyeBA2XcmP1vNK6WIk/A+
c73n4Ew/NKM4pIrVRggUGM80Ak7hKMFyNaw+AR1Nj7FuW5jlIa6wPOoM61dx
O8qqD3CaOqlhrzpiIc9PSqDddLwTWKCsxtV8VLlziexvpT7nrC27/zFePoWI
Jyungik8PQAp62GaesgF34ETSkcUgTGo9oOLk0zPcM/IM9VEwc/DhpmmElDq
Rt/thbuGDXTLkhqO0Ryzr8KaYLNoBKmmmvmxOF++QUeLmmRlikUsyqT+wnpl
bzksPVVU3/VDFPSzQx+4rDwbcij0VDhrP+1kIeKZKqdxCEdEXKSMFARIzg+c
YYS+gVbEAjFPHywNblpUTOXZHCk9naQB/heTyzWYkRHzg6pcN1Nnx76WM8Y2
H3OOTilkIrFJO1v+6lns22IFaAVqHp+zxCcKzy/EoZ38O2n1vk0ni8AES9aP
ehJ3FKfzS3cyh2JUxicebc/ONjZhnuJh6aHyZGtpFRftELQbBvaSUbvZlGso
kk2tLN7KOPhNKx8E7IfBgPbsWLDgPI+BXg4TfDqRppmv/e1FUoFWBga94fH3
loeqvT9ug8El7Hm1CQmxWZONmvqlYWwITRJXrKsc0i3O0mgutWjk+sa6pOkV
N7XwhFS9RIiHRsf/f62NdjxVFQwiGXFCKiAcjCy/2S087BpIwjPBx87inFi3
NbgdNbb2MKbc5mwIhzqqUaVsU+xWPv2iCwqT9eB8l2FHC7G4ZhFQ5cn2uGGD
mwfUvimIkmYN53oRlGylvnVk/fTID6o175QyOklCrpUI1uj/1ahEOvpuWT+/
ncThNrtu3baJuAsDV4DhFwDREmMbeXUhQYfNVmuYIE4wXeKDDX3MFbOpEJOb
lu6AWCoJdn91G7bQQyIW5OBd0ba+41noUAnEecmNlZ8QqNw9CnTOK6PT3ZAv
UrWFf8AmjvmpMvCj9hz5o0CUN6jgOnKpL0Sk9Wb35wCwSXpGhzwCifQuXzZT
6cQ82fk6qLGUUzM+nBXlWY41voCB/RVLnklhbbZ2mHmK2QItxgCBHuNkvUsK
SbV4/54S0Sim7MTpV26b+zashMdGbYz/YQpwWI8iWyLoSO4iUyIYwKAsbkCb
GCdR0aGbZrMmm4owOhCK/ZSQnOwDIbDsC4NCPwNnLNnSfx0LEenZFbHWeDjo
qyCL2Ij10N/AtECfqGqxrnZ6y4T0Xifz7y1HKiF0A7e5WK4r9rCieaTeQH6C
BhgC2dWFYrLwscOLbPVUPj2drhEoPhM1OOI+/kZihMIJ1SY+pqAUmyh+xB7y
QeFei1bbbeBzxyjmdCcZUlW0r6D8gVWA0p0udQ13P8ShBDyUr0Vj0uQW0KnM
N9ZCZ08waEFaArRz3n+Efu3YdN8cNaX+xFJnWFs5Qo37Gzh6yaTZ2rlZlKr9
cNX+0bZpc41wXfDJsVC5+46CZid/2mriFwfQ1qwXXCfgtfqZqury8QshvWSs
rJHe1WSahPrBKLx61ywx+zuW6XgZ1M6XyHoRqsHjIR3SL72diKtxWtU/ofdI
bcF2LV3kJK5RC2UVAwhJrV4i3B0OM3utfvNEUSfBnHuNKhfa0N4bi0YAHlva
j7mtUydG25sSE2LUXJFtYS8ajgdOEwcwPPgUQf+95y+t8I1nbEdfQJSgupoX
LF0rm5gBvm4/ZnbfRZ10ka067A+WbyXz0z1BTjv1sXMawO+ORY5b/e98FlQV
Vmq7cj8ZtO4K3T7KtFrE2pfiVBB0AU8mpSa4lsy1emzwcs3ONbCWzWICXLzf
OOyOg4lQlbLcy0kFeN1wzrIZ5A0V9tl9+6hGIZy9iOIHWYthKoI+Txyf3tZF
dhJlJm9KTFuzuHWjmIH4MzaQdDcX4+IqS05vZn6w8XVUl8PQcTmMalHZL9PG
aq06RLNpM7pCtyIokBPUKP27zpI4z3EbEXCJHt5/o8NxIsPFv+JAmcfL7Juu
VjgVL/i1QjXny0CFsD1/cmH+/UElI8MiqmJz14mP1fCYfF+xXGOzLw1FaZ95
+DkPmMkMg0+ltpsuawMZ41zbgm4DjONi84CbYrtiBm1lNCRXmfiwFHCeYqSS
8R2hbarfT1SMNWZbicuyUO3T2XpSxLYr0fOtKepeO9k6uLG36owZpMJQEdHo
0GP2cMe6yuuf899CIV4VghNOkkBem0vP4nzw9uqWBSoR9JjY+2WYELSSqqO5
x9UASenFVT5pCqK8F2MXqcuvr88jSDJWQM4yE1AOrENvwu+9APX/lxRCN0cL
WcKTX1pQgTTjkTIW7RtiP1hR3/VHRH1k5oISyunyF4GXtmar0ZA31T3KLVRx
HGiVw42OgUS9bsv0n80t2Xgatvw3W1ZqJcPfJZwV5zjbi0WBdLq8S/uinaU5
JdQ2bqVaUEJKfit7ddfNRBNs48xKKHCzqSCSfZFHxOYFb27YvCMnmhNZtSUE
Oq8i8slMEEgf8MOtq4sdIpwoSQ1kouhoI6Mz4hUiQ9XoxcgUnc7L7cU66g2c
Qo7TLjggezXAFTsXcRqaDZcF9RGzpZG+Ota9EB3es10prfZeNZyPyQBPc4gI
Xg/GMRRI54pyczbkrqR4GC9HqeOA0AuBpI2zD6VW6KlvkSa1aLbYPEoMln95
IVpaRLT0+ooU0YWpOCrR63W3T1uJdXAbxm3hlZRom/ZuxBo9a13+4cKBu6uY
79jbiIzHrrssmRV58gUmrjNZYEYCFUbsubhxxS4UufW3HdRzzwHuT5sFau/I
IOqbh2sIqph3jWSmYqYZQtty4APBkejY5tg9a247UsJcbFiDoYx7kyYoe4s9
ghVunnxAsdUjTV4fxZMUEq491hgC69NmaM50NK1bWS83ZSqYGg2VAvWeS7hs
/8AuYR/2uduLX+t552rzgpXgt2JAZhut/aRgNXxKnx8d5F3Owz2rts4BiPpo
I9nP0heh2Y76bvS8m1mutSgAO14vhwprLlU7Ur4WSgplAPNnZWoq6Zh7TTeA
LcQOmyGJNvfRf5fa9NU/ayxGy+0G5Zc/fx52siHHwxu61qnnYH6cM+UKC93X
2wh+1Toa/vA9MVegGyxlDppDNXGOPdVgyZOo9INXCBm9ZLl6RGnrgNayr73/
fCaW1mC3yqcRSBDUP+Ba2mRy5kh5ebeTj9iXvRIptGFBeEYi7hdXJYZ3l1uC
FYa9JMtnkg3se9xLcSrG/wFkdwJcTkyNmdy2UkF9uj176z7YcfRR4BThbaOE
gSaiLD0DyN795MCPDlnBTKB/tEXngoxh6I5QOgwubOCQGXt8NbnkKdWlmXgT
1pD4FIDXiUqkquRlHsbCnc9lcpuXtQS5kfJZHfaekAEquBnTv/U2Ks/aGiUj
f4+ac7Nl+MqSQgq+5BRTQzGO3PpoSH62fLg5GeBlAyYpbcWA8whOy9iuqQTh
kcje07WNoNh11LDNlH/sj2sdvieXNxOnmf8HaHfSTU4gd98DZxK6OB+moi4M
xyRo2FdB+uruldCn2QtVwka7v0Xb9JhzOWTeag5nvfwmw/UrqYZRNcIqfxwb
gR0yoccNV8ZXTfGYIlNQ/m6cUwV0S7Bq8Ar6gXlo+JzOVvleMvfvDsB6rurE
lxOPs83DdRMAwL2A/GuBOrIkDLudINlRoq7Q7Nw6FSMdsaTV/SXXl7vvgmNc
Uvpe/ERC9W5USNOkOh1/62YkfJfLhl3+Pk/TyauSHBE33MbbSj/Yb+SmXB1y
CUgrBSHd2S76OBQ4zQTOJxA5EsLLMoYwZVsQc2hGmsvzXrTTAtBBLT+9Uvt9
aUNI/CXJATbfeyTqUxZXcgBPfyMvK1pOSX0ZeCOCly7gaqLTGJITzfrYUbEf
f7YfIBTHUd2WV8r00f4vJzzrW+osyeFCOS4t2FUt/FFshwbxYS2R2n8V6jgj
6JCsoVCX8zmplE+3A/sjPS6xIruZVXG2K5VoEOMYwcyd2owh4cELBYjrzCn1
kOGUHtjkaaqZn9QGcAs+XOCA3Ul3RmJVpYX9HSXhr1fEiY0OkFAGv3oPcpsn
nkzA0po9DuIZxptE3WfQADbCCGa+horAnGxILSPVOC0x0W3WoT9RZsfyPU77
296aEaNnnLqJhvfzVGzaXPX6TeXHCvgjdTxubqeCn5OrvN4cw74YK23AflJc
HPpX3d9MKjuv4JgsgYksmQp5496EUp4akfXmMhqwOdRDr8vVfEJOS/FWlRUJ
ZZIVoA5uuav9Xfq5dll7xe6uReXyZodJTCw3QaucqYSC39V+q+GuZedtGDWA
8VFOI8b9wpf6jgfAD2goVVftUuMOg2r5IjcmeBEjtfz34Co+yfh6ZsRsk9J7
KzhkiM+u+yUWwI5bMSyUkb2XMhlOKW3u06EDmyKOf+YxP1WnqaCp1TycYtwa
cAzmVuhQWOsXYjp9B8bEyP+EaXG92LyHwT5psjYOiD5yH6/2i5x3PDHNp0eJ
nIsXpV5LFeko/yj5GcBhMwRmsu4baTPoOe1riRseGHC4MwqvYSe0tRgJwSfe
ygFTN5kJF7mSYHjPnc5LHG9H1QZB4/nBZaK+E9mxGdxnh2RGLAzyOWM4SQLH
pmUzlfYZSUV1x51IYJNdTquwkV6KM2wkXk27oPsPS2OIOLGqDiIdwAsDDBiI
TnWEmR6ywE1S6ii/8dExCbyvv8/5Po5TJB+U9PNMj7OTyp/K5FSBPlKOQ80N
kbdgE6RyIUoT+f4z7doOHoyCI73C3SkAEPZabPnmcm7GpGfH/3aEOCGWZ5bp
ZprTl05b5XtESdbkDDAFPOO0aJUIx7nbbzZ08xzVQHPRvvNhSWv6dNm2Bgav
t18jsi3+ph3/Gyi05bc0kKK7g34z6wo+AABODTsoSFRBTsmv5y7NGPpvvhPK
1Pt+qiOXXJFAhE3XNgcBoru7ksaSRHlG/nd+ePzhFFjCMua0WEF45fDo93hi
Y7MPMLY14BG2T9YI2WVS1Uv2pnUBmZlTv9HC0euyiT/q6eVKKFDNwKWubERd
iXdc1b3RWLpGrdVtgeVMobh2k+ESgSvqjXGq12GTfhMvKYy7ug9t3FTUCj3a
A978VMsfB9pXRptNbll3m0QEl03Fe89pulBf7taCnth6jF8+no5kaCbjgn8+
LU4JnozvgAmbrccK98rzo0z3cRBAZJT+APvJ9gu1kufy/TJKDFovjxSQSRlM
IR7/pLDTtfylp5WrDBoHBajEmJuBVhV5Aa//H3RG5p47dyFc4+mBSzWidl/7
BI/04GdwZZJL5RpUKdmTAKDN5zyg9cCZhBYShEtV6rRt+5yXQV7JV4On4JUO
rHmGtSBbV00ykn8T0KM8xwiAVuFk77hW/NsumvXAlmKbDh2HRGNdiOY4OObm
SpSPyWTaP0AnFZiqT3b5ygj8/lacZ1KOugIRzUXMAAJn1yLJvuphJUhEqL9f
3DSahVyZ8jezlYF6+VGmRi00WgGfARSJVI37NStZKD7lpgDTpsvxN2kVRZu8
pM78podfuR9rLyjfPkQtXeML0D4+UBS9vFpoX8khEmws+l4XS5cjCvUgiAFh
nNiCdfam8Pthn81TzhVTIUEockDvvOmgPRAVfyVGNwIAmwQzlp1rPqEEYayR
/Vz6O/T2MgoYT1gbs4nwvCZHVQjrszq2kxG5pdaPTQ7Is2otZziDzo6wm8n9
0zHdpvV6MyT5bu3a7iL8FioTgQdddyd+ltu4yNqZxK1//PR6bvDRiQHyZL1X
0JWqWCqzW6X3/ojpofOdsjGU92/S0ilAL8tMD4RfTK4iWCz9n6pF0vccnD4X
Zf4W5NnB75V/yNjBef81wTE3W3TYSG34Wfgkuwui7uQAP/ibqvVTa2IB9LuY
ifrM56LTRHBhikry+ktlL4PyNIdM2KpNZdsX3kJsV8qBMYvQqS/VzZ3D5dCR
tIFD9uv3ixe/y9qH8KcFxUk+K/SW7TXnYueqYvJ6NgEqx/0bWcB/V+f/8UhU
YyC7ktKv0S0TEAHAX9H24YOcMu0J4Oy2X3j1/QLnf+Iadc391tUx3+KtFhoI
AAyw4O5JtNq766kScH7zMej6JoYSYuPgM0icVuV2IYE9ynV30hXuE/FwxcxZ
yFyImz9e5Nplj6zYqwNb7YWM5z1IM6Oi6RbJx284mbl1rYKCqd6luxEOSJ8o
gQ6qDT5NEqSuGAr236JtbNZXarUW6fyg3ohbjcWUVFJKu8IXUy8pHkXvq97b
upnGWoFhekmo9B7iBTOplFm5dASlMJzSqlAuUbq39MIcR4NUkaImeRIR2t6x
TZVRGEikEYWYdiUtwlGR+3e/pQZxGlGjGK2l6PlaGhc83bKZqZaoiw3AXE6x
4DOjH+ExxQaovO0fweAwCUWF9PNf9MMRD9inLQlJ2sit9JcuF1UCMo7/OBE8
qbHs3rHKpVIvmIShVMYVcm8XGwQkiMBONBN4pm2WPIZhy3P3ahuIx0CVQLk6
cqDCt32II0iJMUKjETkwVrocIweR13jQrlWHmRy9rrC6yPivqrF9wqOJdZOp
u2EKwFF05cGXGhqHNlUMwgQMqSz1VZN+rcGP2rvZrRtNb+/Ab85k/yvaRri6
eGeDpJnevn/UcD+ahjhK19GMJtZM1BuYeJmP9CyP1y6hX6hgeTQq8yyuxywb
k0VJ1Joi3bDxLvouP3Iy4ds+MgstpjtTV2d/GzpUnopNUgoqYNWbJ0U5FkAU
LEtOJJrgT+GsRTRvzEOHiNPfAwBcVxeox+2GmKsOdqDd6llMAWv/ClbS6WeZ
Y2YjYGAVxLi4SKD8N5xrbr2qAaIZW/0w/P2T+NuHqIj5RVbahkUFVlS2VFYp
OVobLxQ7B69XrSOw+Pid8jkcOPPRTbOzZTEn+ZeI/A77AtfkkKhFVOuzFg4e
e1InetLB8wRSeD7NA0+DcS5yGyzBO1hSQZ3kSexINBdmdra3d1hsuOZUx7pU
wMh3Gp9Q1ONN6VdeRTCF1uQy1c7Hyx99zSiCMoqXcqo9LiTT7aWgeugAUr/M
Vp00UEhzEJWHuYu3x8RD1QCcJRe5jQUDsK3AHGMqrzcDUhPNpcbTRwgY4Arx
qlvY/GqBr7GzbQc9cfgDpptudjXohwLn7iHPmBkGY11Tr7qlIEoDi17VkKkJ
G8cJ1RPRWr9CrDlByakxfkvIhZM0mfZtfM55rzabi/ZySBXLfks+MbzN2qCW
rLI+7Uac/1oimE8MXwolNUpyzqpTHVHBnLGqVjy69/fA0tVGV8QtcudMXMzp
V0fxcGNnPkvVb70VJknQF3qFApdtm39JK4VDvg2uHRzTOEZDHqcaqfqhxqUO
gsRq6T8tRZ28X4/DFPU5pVy4vOCpY3tTHsJZD2zekOe8qKfSiumd3m5ghxfp
WPZU8KK+d5KLSFW5eTHrLJ2dmTIaFlhkmAAMghyWSRP4BYwVVF3Ji3TlWpPZ
M+nwteBsAFhF6TxQlWHZoDo1pCgTXbIaumvnhxMDcIFxQYXJ2Ugwh38Nwuwi
OsB9tY3+XyPq2WoPxzvvIH5BYvDAgA8F9pTq5UwcC/W6sv7RR173+AKoKPA2
FaiCyoOekMwLISrc3acEI/431BRRebuTtBNxkP5e/0yRyCfN6gsViZP/eqKN
1LQN8tYZ06fE/fsIhriQZUVI/cnIxKn/9VXAB6UmDE3mu+1740ApCwtvK1S8
H80txX3sbztZA0GTLjUybrwsNU++acB9sNTxUQBWThPh+JxDRnqQwx/po0oO
zsMRjUnjgcb3kq35ErER3RiDEgBDvDTCkIkdjVhRPR4stqNlknH8CgAuIWYg
N1UXnGyxs8/GX9t0s20W1MuOjPJ1QtSqldxnqF1+AI0Jg/6VyqyCMKA5daOD
4OTTOv5zo9fcAs1XXCQr5mqEdzwCPrc39I7OJhzX09flemT288A9YZvKw7a4
I8WDICH9Bf0yi8wH62rNRQJ7GZac+UznPOTN3DiBDvN4eHsXQ4xvzalzj9oB
4HNJQRV11njInXrEgIwKOjxR309TdGvTIlNzg66FIQi9aZV8BuVup6UzMaBI
0mDERwuVuMmpSGDB0H/bU87ZYbrNqjPG29UHn2RD86jbktcxWceBhfducTQ5
n1FUSIFtyQkNskOWO04vRAjPHz6qdBrF4yU4NP5oPjnATiq6ylT4FoQQoj5C
orjqMSpG+awrkhkCPRDHHcTPhcjcmLrq/WzCD+pCCeuW21ntX0UeeLoB0fJh
x+iOz1h0/nWHwcqYULdDbhdZoiuO5bF0jKzz6kho1laTCCY8lq/LlGrCAyUh
eGx+7J+jBhZeuxVBIZTLNoBe2OKr66P3hYyk+CZpXesnSUmHsard6etp/1dP
erh36GAC8vj+m8zURzgdgBgoe26f40FH0ycS1RXgNosCv2SO3GN6ug92KE4D
WFciVpZeIqUz4wCHVtvl8p7Wjlf5oV2IbLndnKcACp6viuRGNUBVVwyjetJ+
RXBwvxAsK0MesPo2EHXWfO2Ocy849DEpEHvhRk036pFHisK4PsTFWVVrxN0b
s7izyIEZP1gApznGotya0I/O0M/gkhS3OgErJ6MER3HbWw8rud+TRg50tFsq
uKIHHjjIW+2qdp0lEKJDWr6WXSfn4W1oJPWmfnfiPggmLoH3RqTvp0MDihmN
p/pTnNt1YdzvVc5wqzqgYFcHLp3ubO4MEjOe47VbqrTXN7dKJUzn+ycnlO6B
stF5kb4LJR6uO2yZJK85R+4gvRjFVdyW/CNVjWZFMNh5FKYMI5NnFgHkO76j
/yB3d9OKT8xkFbMuL5qD8zrgIM0udlC7D1W3gyiR4AWQ/zMrrWgReWtwAoyk
gQE7pvGiLOkqc14FTCSk8KNosjXOgmk6cBZ0R7Vd8eFfSZ04qn2ZhOX54WfG
RIy+kcsoLmUoYdgXfct33YiWOSniLRONYATV3M6kcGxLEZoqnPfwUvWh/9Zf
NQxvUB3PLxxMqMotM5ckPuNaBkNWXJOA2UtxUgkaeDeqB3EXFTLKzMOhGRwo
e+Gp6CHfMASPnegft5FsnZiXo4MOCxvem03SstLvcEcDOhk8c0BZG6F8UexQ
L1NH7BBdUsH6Qi5FXnmt3KkhzdAE01tIR6FB/JLthUiizmHAHk5b+3oj72Y6
UcDcbygihoqTP1u8omHKIbwTJFG39qFOyjcnNj8IafpZ0/fSaFQqD+ZIo38B
quI09nh3/WpXJJQ+1eyeWSTpCVEc5lMPMlRs3nSYGCqIMShP+d4uQW16AWto
3hwoxJEBK+xT2dzQX0Ix7sSljf0ozmuqNiXtEFTfp1AKWgycImcGEeQ4YH/Q
QWrMNiyhbBtGeuo8TiAnBTpYTnyUiMLjmfcvcnwUAPUoemxMMSfcIv5k/LJW
4EZW46+nKYaqMqlaubm3GdRjv1Rxgob6waL2FScOrHQqf7Jr/D9vwoXCPLtD
xlzWP0Ef993q05yCrfsxGjDLNhwSyCZnwdyuueJwYdSebwddgP7nQp3M5V5c
j3eSIsWQkvS3Huk0KB5fCN/5eIiatYUo3Q28JOR/Isn9Mkb0c+ps7/X8HEZX
FpzXcITx6AXMf8Q0MZxCD0lfasMEuoty7ykBH24X4kc2KYnlW5zu3HRwsM7/
u3BYaw90THnZlH6vAUswU0uXOccZRzD/WaRhyEwpZlWpnZt6nEcm9vx7JsuL
uFKwvfDFBxsNoMC0N4pOqAEgpd7ThnvGISWOrigOJYE+SpFrmaIdLup7pTCB
OSBxKRZjRUDtNWYYW+ZzeT4YIZYMC7nR3rofFOxTzrQxa5ym4qaI+t/yKOil
pxcqc7iw4TVIlCFfGgVLZW9gtYGTLjqeVYGouhJmND8+vTjaQXZDKxQZpCdZ
rW8/93qLQyOYV6PcfPJ5UABxMZPgN3QILwYiiWU5DILm1qkfpPhSn4zztCq8
Vautik7iH9penaxNhDpa3LMO8uEPByIBxuQv5HJ6hjCBqu6r5WpYnwHE0V1b
t5/QeUl+QYguZtkvErJWV6U/NZkFnCvAVcAh95ZIx0yXfqEfAIq3RtAxdHC8
gVuHgYoHi6Ki9SNAzjXIClgykZdFiv91b/OT/SUNRSUuPYFEhvU/bruQVme9
smsQTzZdGDCqaglHlnDkFV8BPtERrCVD33cYP3ndLUJG8OkXfG1I/s6D9yn9
5LrGn5AE0UOYkEp6IQXn1MifimdFe79KdHnmveqTv93pNJ4ArVOOF57Ibq1k
bUyWL0uhsioEC7ydnxlhCMH9EAAwXonIcT1Ms2aT5WIspCoqHQDHsifYbViw
CfTKusUNcZCag4wzCISqYwI/d1QgKmeGpfgBnHWupRaMjoFDcbL82eHPDhpV
Wao5GOMGKH/h0NuoOFIccs4tKY2k877iDLkZ1M+CJGcNoujIJeTHoAvkgwy3
oCCvCxVgQv+AyK9tWBtSK7eyWGjsxFZRTnRcShOsOcBRxWdO8u44iSoQAcsO
yi3INK3/MOFcXR4FHtxA4UxdI42l1OKYs2fFVBq/WlRI/JfSzvsbal1n0f1X
Lp+GcnsNt8ZXWqNVPTGthlYj1lCQMZq39QTIwKzOEScfzidk+f6VtLOyOJ7B
iTNeSNkjC1EnTz1DeAxpnlIYj2Y9AG5B8TPeFUwKfwZwD/4g09e4oTMBhPM2
1zsqoFUzKVJ8+5+dYHJqm3MuVaRnwrPZbUNwPi7QqNFGHtdAHSrZmO1TKVAg
Qv+xF6l2aY5CoC+go296vIxd53og7lXZz9/Cznxxn6R59/y/eS7iWd3F+Dry
9eUs+rdwvOvjGBf9eTkNuhn/mQmPARGJ2QnIqEF7CM3blEW4S19Jk+Bepd9m
zA82EimtzJfXiP2V1BEJ+bhGQSFoYWsH3EyCJVg4fTzZ7qTQBUlTH8vXV1vI
3u4KGCE1l3utxyxSbmSm/J+AHFAM4VLalzsKOPZIttqBwxiCPKnxGiZYzNAG
+hRjCYsvH+AAgznelkIR92LPA/UxW4lNV37TsGJTKbq5l8kLqGGAvrQyxvD2
yMZdGLSXR9XzTMcd5ZgKizKVY1ezSG+2OaEpaiYIyRHc+IQ8G3iHqewCkHB5
7Pquzl6j0b9DBc3SFaweqM8KtUoFCYLCX11avfi3EhDp4uN0SaVTe0dktI99
uwA3PphEvV8wOLMUiqM1c9S7qpzEsM36a6+B9noqM9jLgQDLzt86fJqgqYML
x3fbOYkzmeaILm6hZqo8sBLrZ8VNAqdbE5lTwJoXtlssT4HIQucpdCMaf1DY
iynZHO7EvffzmT81IJ5iOu2TwtjDgNVVPW5Ux3NgJt/gLQqID5lapI2HVb4X
Se3qi7IerpX7dTZND08+dJ0RVakEMauHaIhK/K2PMoViKxRAGNOZ3jJBaGuu
0KR4MRTGSkwsQz8DSpoaWTRgpxDdoJAurF6wegpM3svjabM01mJH/pzz7m/e
r/8SEK6iCGbLSbG4sdjjAfCfFfLYzh047ip61M6vmAeXpxWrnNswK7Xn4i/H
QnpXo3nod+hC3/lt+yfXizZODhKJL/h0P6E1UXPed3tonyIm1FfoZwjE5a6M
vrhqyrM2jJ0Rj8Zol3ZpXIrNTemGrLv5TXlsgc5fGZ4Jscogt4dEemcUq0bW
T44R9xj4TYX8UVNwoQbaTwFXMIaez43SKHvgkT0ocOb9AYMxqOJUOrRfRHdR
dKsv/DI6cJsuOdZ8pPqGd37f1YDtDTSjRHYci0aeFbWn1BSHVr5AaxJyl8uO
vRGZ2iX/9sYj+tx8hOE1o6nRecDzbkjtUOHWoI39ncrdVYNfLVHVHWBQLop1
oRwht7OetWWl0ulHxJnuOVdfUpmDX2zXSQGZabXgqVO5QIlZPG5du1e5UM3/
6LE+ienvXbDtaKvJXtywm1HPlqvnrq5aJCa0GbQRtIeZuzlicmOzjyCT4fDX
s6HorJ/3ZfX6hsntfX2yfV3VT/Njx93Tg5mBUbF8ONoF06WvA7nQXbOExJ1t
BR/anQCALFi3PTZ6lC7UD7hJ+U/arewUtW+J6l0drFvXkOIAmMSM1Qb4SAn6
SLXVBVbjJGdMdvndllKmxvl62EyrKrTyWk3+GFlWc+e2IFsGpggDg1oT/Hwu
2FyubLQqZu6rtDml7hqqdzpOgt72LZ+o+rCb3HjsJbkbn+dTul+AejnB0krk
iBwuzq0Ji+0EMhV+bPf6WVFxraQ5x5w8ctXmKnX2b/IBwz4CfVccvOMiSmjJ
9kxqQ5zIdBZ4m6QRuGY6JnvJdh/LtueyNylKsJ5ymVAjgWwHkjmT6F/HNuL0
BWA/m2gpNjUY6eEgwgeoPM8eXZJS8tL7EmHecpaerxSzRMs/waanFUfJErTX
fAWW5Ep+ud3mm/uXf9LsA30i1xeeivzd0bamPAKFeTOC0JicrFkcWhTdYo4s
dHASkP/AqbgrOWCJvEitTGn47IXsZ4cJrq5+bH19Rdqm33WLn2tR6ttBDo27
KLPkk0b19c0EkY5sTOeVfgAvAWQ9yDGYnSzb07Mtdzte3G1p33r0hWLdQN/r
1DbQ2bOKqNKabJH/+N64tIO0GEgx7gbqE3NlNfiDtNCz9rRuEDzLEL2oFxtq
w8a1Qbu9amxMBn4ue3x9ZqD7W3rBVao1wL6eHPz0CnDKiayGNqu5NOZsy8Vn
VS8Bptb4sgsmuvl27Evth+FRAHEU34Q9zpmynkPn4MEhp3uAspu8f2kJW82p
LwFmedCFo+MnK76tn6+1wDh1eUNLyRDQmUUJ6OSzWMDXfitDP4QFhL5I5XSG
yCboE/bNP+dBU15OlkiXuyZKKI+F8imA8ef3UvMChmoFcls/8jG05QICeaqy
yNRcomU3kLKJJry0kOHadeBqY72aHj7e18CG41o+EttOdETTaZKtlVMVQkDI
vD/+k6A7z4W4XLnzkFY1H9J0/C98I/PhakQJGTmztbhj8mBOizfIe8DMbMdU
/Ub/0G9+fuOVbJxVQhabDKGUaHqHz1WMSBiZfRvoMKaF4kxr1+eaG08RQIdr
t2BLFyHNORyQ5zM83UtXN5NexLLNeC4a8IriQBA+v+hmcIt66KyacTL7NBeA
F4laZnYsKegJGse6k4u6U0LxVy9M/2P2Tx9jgKSs8fEZh4a1Le2nU5eJPYcL
bXNXLvW2O8f/8+2Ck1Uz5olw7MUQO7J0qV0c18AMPJ6G0g7lKcZpigNHl0kd
Xd1wY8Nm4qJEdj1EMHKczfGn4OUjpAwnRIsqgr44zs8mVAY4+3yJ41bgfPUP
0OXOAkHvVKPjioK4A/a5iON+n/JK5zZomFnR+opqDotBCFKSHFyoRPg5O1p3
EYY5mybCTFzuRmseWE7rHuhNj/jLntTBavs5RjxCbqO66E/QP0NPHPUa5MyB
Qoo8565HFui8VNpaRo6E/pi1od1FDTu3epcyjWjDGUDLLTV68Gi1KN5Z4NNC
ug6N7s0JqBrCbVdNzd753kaM8mQQm67U0WhR9HAbjWpk0L2LJWNWDuAHPexk
MHJsSRevgizVdwVZoETqadNbJj/OT3gfeWokjfH55/jYQ25jwkLcbyirBpV4
0nK9o1z6XWdv1iuC9kf1bSpkDFcMDMzduiYlPJ93m7L+u6159unUlXSqYkMY
0+HOTmVpYCr6P2rGbPiHmHcCTtpqH/pD9MxhZGVe2Ygo3enYEOZZ//H67JOf
mh1+kIUCe7kW6eM5ejFFqwc4D9L+Wv0yhiJ+5/stmJZ3k/IpZON517+j9Xie
6K+EzgfXMrWtf6ABKDe1R5pXSHzgy80wsTZDXrG+t5N5mRQn2mvGla2D4a+6
iklEY6/5ewly8Ns9pa+No3optljpE+Extp+/0ZyQBOayIpjNjz8SbGMzyptK
ih5U/UNsrA/DCoe/qRswD/9p6s+arX1p/SHzuw9RpxZW0BHKTJhB1oj9gYYz
8f2V/nn3/Yue3HCl1lL+VvZOSgqi22WtLpzNTXBbtyEnYxp27fKCqnpbbguJ
rnlJMGzYilngJ7wc20a7zwSMMhw/HxElBNBbj+LFxDg8+8OlDDskP3xBzDpZ
pomY1h36HRPeD3nrYnWq40lJPeiFzq9rVnIKbBpaZNGxeYkVyKmlhVKKPgwm
kg5z/AuDabKlZoHhrIRbJs/zHrou6U2qbFaxUkr/0xFMHak3KOCPIS1tnRsZ
FkOd54BO/rJYcifCQWc8MZjW6hp6M1WxdzP9Y+Wx0m8xpsvMcSJEZFh5xsH7
4cgXwXbrzJXrTKsmSNit4p+guD/9ALEhBbL1PXaHp6AoxY5SN3/bziDMibxP
JQD3xr2APlKn4d9o34vdnCKQ/Gn45PeCGDAC/U6MJdj+FM1h0FHRnobbrtL7
jIuEyj6tBciREj0iknJJGoavMyxMPWveyXt02aMm3o/edEf0LWCLZ3n4Lh42
FA5gGwQnI91cvEsRjUF0vEolb6eZu868zi4ZtuNK5P/nwC3zoOIo2iYRgOty
1WJFi5d7r5YlfttwtigUwfzq2uwtuBYq9ncQhOlds688VuqX17CS2sFkn4fT
LYOn+8vjX448RwI4Xr0rIYsqIZjGZT1mgW5ghDDwIPP4x3iWNH6Cq7yj+vb7
OZxnQbhvyM+YOHIIqQU1qAh6H9hqbcU3IGrV6EcTkwKVo42XwsiHb4+GiiXd
VKb/Lh3UBDJXSrHN1PeWvxUfmFcVG41JRtRzO/xjVMPcatHfasBeLM8F88Ep
bY7B6PYuvTRQ61pz6ZLnvPi4aJKuhHuh2BMMMCpxCzdujncoU3UuFrEYP7IG
2Cj+Jy9RXO+jh3Ilh42erDKtMRZ7khpTvZF28Nm9uai1yADGOp6533TfEVWd
AvXIIwcxPz5fvdhAlJ7peBgZddpOn5btv2QUchkZgAHMRJIhR3sLjy6y40mS
ydphexjjhbJoVLELy9STwGiGz3XXaxWPuv7m5r4xnk0q0lc2lF4zl1b2YQO9
je7xbPWKW2vpzTkCkdZcXqbGj6ru0odlWzrougsCxa7oIdpO9/I7VQmaghiA
h/3qZmAJIJquLHN1AQVmJzRJJx7k2nM6L97ifKnOt+IMPP5+9BOpB7WrOZyP
ugEvhcfZ1rYFBi8RqpnKK2YeKFGN0BtXRbkqg8aWqSA57Z690GXnft4aIfcn
DTAg/BV5ckF+CUa1KYu2eIrXcv5jALqMSrQ+sPJk9QDTsH9dlOOXVjY+aPHg
LHmORqET5KTd73yxSqCP3qIalnX3j+YQE3Ehjny2+kIP9sD/Q4nmDZClK10V
kGL8psUVnGIiynYQ1AAUWPO/wywhiebf0DP4XWLPCKP0K1I4c7WcPx6bR6jz
DypHtumbzVmwW6yVu5XdhRmkd+txXsoBzB6XxoXcfkf14pHPtUdSXysrBWMv
AcEskOzDkJ932Vk+yrMmQy5fe7AWJNA90b9LkNMKKi/0f6Kb83Dbki+nVeqM
IKfwPXrkGAwXmVY7StNLKYtdKRj7DliMhpVLR1NKNkd/LZr6eyVjpNYtPVN5
E/hN72wISXGbq8cJpxqaIMy7DOmfR162yHtIfJowmN771EELsm6/EN40jtrR
TBPZD7hDzNR2qLUMXAoMIJK+p2vMDJFHshXpp9GJHOE7aL8FCbFZXeRyhcjx
J/t+e0YNgEyeRJVwyFBkYTwupJ5YxKRc8UOmnA75WJ5sZ9QWqRlaqLWey62F
Pj7/I9EqPb766FK1V5IJc5uQNxTTJqL9CZR969Eg9SLYsMx5kpOQcIuLPrlG
YRHAxOUTCUmlC70SmsunZHjJeQeWoCCJVSn7JiYYimcuqdzJivnE6NVuq3Nd
vVPC9Eqo/TJ+Qw0EsTHLNh4cQXKGqMApEilUAWhOqZHqx8a72XH9N1F422VH
7ATwY628mEsO8QZKxQzJxpuZuUStYnmnoJLnLix080fehFlzSe2sYbbriAbE
7M7Eo6quVLmFKvaiSWhj9mkZnGRdA90F3UB33ppRbHfR8DwE2hSuWhtCdEgA
ejcHaPETDDeh7141UwiHjvAh+UoP97jFuNooHuSj/vFseKi/UamdIhFQSgpu
86jD/CWjCneMdoQcMIcscRsSUTkKR9jeGkS/EFv4NBZAFqa71YfmHlOYGeP0
j+QymJ7IjxpnOB5+d5HvNcpXG8WSJCG9tyf2A5P0sBlfEbxX5cS5lT1baNiN
zNkKVwz9qaUKy+8PhZ+HAtzuT5NfgXzcQeJyMChF2f5Ipmr+9N9awmZyMXLP
/Xifmol6B2ViJ/17u5IBxu0ShIH2TMwJhoUzbIS36nTf5CZHHCiG8Y7Z3MFg
DnxVHCzPR8WaNe4/EmEq79n6RlY5SKr+SxgT1yV49dyO2Vu8QvjAKGvwfQFJ
1WS22XRJJ9MxM5Xg7sPjA+b8DrmC+7RViPaj7/E8wbX1yONt3XqL3DERptxG
wkELR9IvyoQI8q6YgmcpGtlAL18uhC2TIqDjaq5tSWSx3SQtmCJIhGjtHVl8
r/NxP1Zrxevd4P2xYsnDOUWqvRE5JjLtD7ZAhiOTfukiaetjduWFOZAEe2OQ
PnXaOIb8HJacfdV3/nGetjhvLDY5EwDe4vp1UbTmfoec5rjGCAEvRmef+4kz
bM1vnW+rLeXHetzq1ViYYNebxicROGaU/ZeRimdlJYL5wmzCvWMsD2bIzwuG
oWywos8EsBrSLUA2r9c9vvg+LFpEpHuAP8RyKBuFUauAulDj1hr4rUNJEGdW
Nm0kSAKGS2dOYagYe+bCrhnHgZrbctf0iY2LTQz2/Q0Mf1vb8uKXp9fc8Xoc
A/wx+9zla6O0IZhsgjnpq3z/0JeUM3CTnA3lSy/fhSpbN9SJG29phQXkIyVg
/tjdNMHPjiL6jnDYK4GDfmoFMWA2TzWlJEfyFMKqhIIs/ohXHGOZkSfOI7su
dTHBVnpObhj6coAevbKMW/pufet47PrgNFhMtOwm+hrP9rbRIb7vhvR18zfC
Hj3TIvPbUNiuvLh+q0VTfuRJsu0dIt4aAdCIJ+FWgsgwIe3HuzO+3fn+drMm
psGnQRmUGq5I3CxCShOJB/jMMBV7ZhfjujvevjHtiY5l8IVZSjd9pbu711t3
7MeL2Ud/4IjqUbRuCwwACqspWfOFisEqfEQ9w3STiuzkuQfJHpcs60a9e+s3
vk7WeN8dt+stnPhHRWFqsPa1+QrYX3rH3ZhAnIUVHUNNjJFiGwGM3ItpEA5j
FnPR83j2ggTS6cr1wsXvFJttaxfOTYNiZ6lmO3miegb4z6NDpMIRAQvStyci
fCnu2e/1oCpymSPXxxbmATwirhR+WNA0WZBYQFC+G/enIh0yZP1ilzqvB+Nw
QhPob0uHt0T6XcVZ3hsQrT+FhIp+XCdlPlK6KBwTOJdlsaiPu5Ca3Ut5/iLE
hpbIoW4FsbEgZfsvN++OV2UzUnHbqW2Kyau3LZ7hSu5rs5Oo8wVMw5EY3Jvy
gjOHnnDM5ZxvcvWYM3sHOBYsxdnplufl0vBxjF0YZZn/rPIsoJn5M+Ltnwzq
wzFoCZDkd3dalBqsgpBK3KeUbMC6KYVD13ZduJgPIn+E7oGpIU8KTiuOlots
NR1myRn80LVbQRHu8pzel9YsskOg+Vwu1a5iFBKwa8+6xAcPi0j6IFkdcZRn
lsch+Oqa1fOi7UoQWaOFz+/j52BNAS8jvBLc9L/Gx12aiWNNjIdsBNSm8u44
xC1lS7cHKEyuQGCBm16J3JKe5QwIQpufTnFpAc8Iu4RarhY+k4MbHuJ+Bm46
riUDanFMEWFaCgyq7Q3ecYYzZYVHCmqwMM0t3zpiu2r3MQw0187C0w3OrPrI
eGiPoEyloW4v4Wn36q7qmZ5CYZllEm5/nGrsqJrF4RHjFqfVix+0zEV1Xfv0
8o82sS1LpbYkpAueyh5GD5bguW6812Qeb6fCvbWdGKKJgwgn/cdZbfnxQqma
AaAxM4ghkePiTkInm3ZvPijrLWrFfzleUzgmBzyAaRM2memOZyI5EBP0naFV
97GeUq28octYva8RfIkovtnfDWbRZ904PhrWPMpnBRXEDXRWUzrfH7hzUdF+
WFcVW29xnjoPfpGWgd2DrjpdE/FXHkfyme/2Y5IpfR5/7J/rJfdg+e3ZNM4q
YUqWWaKAHRcMslszllhrx448acnqH9tUcC3a04yYJV9rd8f7e81S16+IWzUl
U4qQB3O+muq+dXIp9VoBmI8wdUpCDQcLPKuUaCtA63to3wQXXZOHbX7LlEds
rC31VAXrVT8MeZHaNAXNpiDSzq/8FFXMf3XwQzx+93673cEB9qko1HsVJjtw
N0gltHg6JwplFPoArBEgKuDWbPHlNgk9bO2pMlJFr4PpV3o6VN5f7qHebDcF
93NY03UaxtY1RhKPugTIpATtBovezphZDvj3u6mJgtsxBkczFXI8vpTkCGnB
dfdZ7XGYJsfqg7eLp/kLBNOMWbAlNdYM/mp6qSwbJkNxSEIGGUlr7VQrJO3y
3OXmCKpRa9gp0DpVmBhvYt1EjnBuUnrG3YqNLq8BI77qji0Qr1UGxjiMUiii
63T2TIume5DCuGe+2usN85kKgMqQp01aTciQ3vmC1ES0QKeSxgcEzBDnHFk5
tOAXVD3U8oczBZJmCIu/0/DFuSe7dm62BUgi0m6L9GeznGyTKTT9B8e0jF1b
tEaP6T+5V+kyTINuFJlIfzgcAuoLfUAncD/oDbn2u8+TXpGyNCm7f3MuLVVu
hH3Bw95VfEKDh8I34Gdsr5tRPJ5gWhxwJgwKKGP74agVL1TBOJZKZ7RjtWPG
Pz/jdKKOuDPlKIGYAn+SFHbX2jy2d8ZtbEBbzjK7FwmYywCc8CECZIqMkm4k
yoezcYUVBYsj/gwPMZu+GtqUprKZWDXsALPo0DS/dmoYv2o74Tmv1X+8l5Ax
OvohjY0T53Jabx3Fh/WylT9KSFWLHb19r/btxYhiBZU/7NErTq20fuiGF7rM
o9Mdb1w6waektUgRsgnjAzDD4jGeEP/v0YHaLeHSyD02CkkvucjPma50xKzS
Q7kVK/IFqH12GEgG86kQmOjH25GFk4gjn5Vxz3/tvb7hsl90c2XXFL+WQujy
HZWRmSuYdYBtN44p6Sz5pBsgPeNElwhddfR1oDeJoEXReDwI29x8Fk/zdYMe
Ht14Cg24smqTjaq91puj/LSKyNFQ0KaW/KFgRmze68/D6MXceyY/FrYxL13d
RIyzk0BMu5s3zoJbaY8BQ8tUWgHjOG+AZvMK6U2/KzWMZ7X8TfYbQGZwI2zL
dgDMuH3kHSDj2/+9l7rg+QlBnkOo2TCrPwdChzhiCSRcrabWrS74HnyWVLER
WKxM4zaZ3JKDG7oXYQluIdayyMywQUrISls+l1tX/BU2nV9dvz/j+73iVBe1
WhYyVBlJv2z2oRot5nTM9auZR4bfOtiq1LZ4e3JhQk5qAjloLORaLOUr6fmH
Nlv3aw6zihmhKLrXyHtJkm3b7aGjTuDZFSQDuD01W6Q1VAesMd9OzkTGwC7k
cy3/3GY1d2Zlf1fU1CUljUlf/zQfA4WUkByeqfgni4Phr8OwdSyLVCjY6Fcv
yOK4jc5qqSxrJG7viZDDN6iQp/U9TY5YX0T3fa8yw3iC9t80bkF2XxjGa4zp
OplPVkYj4JUYocU75KVOq7UnFKTulFyKN2dXgWyukEV23ggKaCo9gnxqclBT
+D5v67E4n+57CVWlUojpsSAIy7TCz6HbRdh0X8B9ngLSu94HNwo2Q0i8XCu5
K3Sz/Ej2CUWHy5reXLpTcNphFTkbVoRL+vrF0qzaqiSvvdXe7YvhbAhX289E
Jpl2pPmUCMp/8U+hMZrK2TqFg4bzHv/eFZJE1k8WS4klequX/igm+YEJIU+n
TzHEO/Z4b0SKFI+Yw4yRfQ0Kg8xd+chg2PybsTU3YxX5IQqn94RlUayeM13R
BMd9ykDfrMJcG99OsUl1iFsPVxyVJRBXKVx9jtqVPAxGzCv6hh/5QxIkXnM3
Y+85CZ4sUpEStj3ZqPoq8CI4l12o0Vh2nw5uYJENHY8IKLpzopNlliUJmx8J
U0bRRoIDEYxqOvxIrgLHjkRYmZyofeWIiAf/lVBS5jBUk62b+hxqUXvzVKAw
/QflJkFU0o2Whe4hjVJIaN/cBELjdsPCwEZtRa6nBOGAP+z1yVikcmoqZf7h
S+YkH3TLGNyqp3l3hRRtS+rcCCrx85Ie1FfFQ50nUKtsNu1jFEX6gjcBEcWQ
7yV1A1aFHpPJchgjbZs8CTNxeeaZPvineef/5v0Rd6oRV93WUiRYLbFiV6Wj
ETi2nfShnoyCbWVmj8NYnHbuQN+kiSVMA4VlWXN+hZlzQIZl3RLw0mM3eaAY
I6dNxJMmFGeUcx9qNXX4zOn2Q+WcKO+voNkUqVPHYXLQSHUs4p7uC49Gp9tu
LiH8nFH6+sPtDQe2HGlhqkKYNYbQH32v7WUlwf95/D0n+cBA2Vg/gqlJPDkL
PI+z7KY1RIB/cIS8QVQqcYK9u6HDY0l+WNFH50iheggRMB1M+BqRq1uoO/rf
oEYtqOIfHfvYv2sMASc5dBVtY4zWkEphv5LjQve/zK09LIPZPXcmydskfOLF
dRuE9OGnNF7fgnEMNLu7lLlm7xSAKQ9RIX1boJKUyvzZdlgziLwZDI/qV15g
DjQ3fm98MeCz/IEhe19bpycCBQ8Lbh3JiJWJDyBKLuRXVE27DpBpqwozfoTx
V/sa36gCo2a3Rv9UOApieAZJCBGqds2YORP/Tg6GYMmVNVtBJdrTZmOYcoCH
8kDxT6ELoq0JXfjlaKEOZ63DV/mhhjuAExTDk1Ox+rVYgSzmuXQn6n4NwTub
ATe82lzjF+sPzbiARZoemAI8YhnGPsJGt1NAJhr+m5nXqGFlVPsxppjSL9TV
Tax3ZdkntETK0On3TapKDzXkfwcNYrNDLgZp9jp6dnudF61zGMEan6gfziJ1
4moPaVhmypj+Kn+/ug/USL7nUsaw1Vu7Ho+UrWP8nOp6d70tCTT+G2j1FDhN
LY3wGfnki7nZKdDpuNtC4ToUpDuiX3WYSEIfaxDPuAOkNiN6/58j0L4+3C0O
1ysM0PdU12quu0s8W7vvV3Q3W1+IHzouch8IJhVGHIfPAEV6cIudgr6Ai0Dt
c4h4hjn/+23l4VtWzgUwzQWmNoPie+shXER1oN2wrsR5P8gss6xsyZotuPNB
/Gp9+HLb3dOQ+Y4ybtaTPSr+wMTbKdkuT1cm+6bsDGrOtKd1LmHmK+zAUVJr
6ptXeMoLwCkBLLj0t330dziogmZ+TOm+y1ZDiMHITi1yQYTNAA+kUCbzHT2r
OoF6DHHrIiQq/7hlp/A++/tU/8MQOi4I7FT7w2f1L6URR3azCNuE1coPs1F/
ftP0kwy1gV0mGHMHjpCE4sGWmcrlattBP19FvPlCvR0wCNjxCUICAAHcJOly
7oCPDub0SCXIYc0N8jhPLC7VHCd+9udHSgnb+yTDSGixxDq8fPujiMwALsGI
BClo43+hebzIXJIK9HNinnSTGqLR/xbS7z60W4r53iJkKKPX6BQ+q0W7n/kQ
RjhP5aBrqg47IOZo4zJRNQBOj+HMUzhGHxuv5/DQ+IMXUhMJ4v6X0S5gFAl4
1vvQQWxAtilN+A2ByE5qQJsFLSWnwBHtK5dNnoFi88Ic45Or9yuOmvJFX7W2
90PtZxJiiY+kacgGuqdGbkGsJrtssSZ9zHOlZYNlWpt6pSxMu6jxg1g3z9XJ
JigQq+zfe9jYH5lIYC/8BQUpuDxzpC7GrK2H6fuJLg+CqpRHIYAcPacyYEyX
igPePvAYI9sonsQkmcVGL3y4TRt0A7qSsaII04q301gTEkhOjHOXfNL1Dubc
qg8tevo9BOUrglfnqYvcynbFUS0AsmsIsIOWOoHqTWV9Rod4LDVPALw0tdJZ
BhrYSyNzgDt+MulHsghhgwKuVcr4T0fiOhAypPpdNXvz0UyzFvrmTpUHw0yg
1XCIi9QyecFqoEh7leoYjNBvk00G6dr+kKaH6ZsyVw6PJ68sgqah5uHjNR8U
2k3xZR8aEkT/NA8E7zxk28tIg/ryjVf5osUQbfyu3GtxJSyvzj74YnqLHEtO
uQ1ODKmKlHQkRPWHnJjTQnxZbiEBCcnMX7yg6tq81Sh4mg5wEn3YnNysq1+o
b3devmL0MAWHa9BbQJm67Jp2jLDCidNSZapFeyyhdSTO8kykzr/sU4rTlBUg
VVlGfyumIFehKfbo2+vbnF1J2LMGe3KHNhG5zKhEvZkmIMb4lfk21YKjvxSv
N8XEcEihi5UFkQ9ognHTjRg8Li8EQg+H1D6AzSbcja5cDcl8z/JtkYsvQsvd
dntDwweV4pOQ4JsM58VMOBiVKlQWQHS885+XRKEFAHRudmOeYV03AQ5YYsDa
NC/5q7HQ4n0N6N3/Tow9QcfZ/uysjAs4QEJpwxRZdrDHi0JUji5XLnk20G9g
rIzaA1Z0sMGjUAvWLCcOYBqauruW1EnJ1VHMBtNE7fqlf6mU1hwSuR8lPiUY
YcPm3l3iXu/l4fNkDe1T72x0STrzAU9jZvyGqduVvz2xgqMTSk/d7aCbrEYa
bqiGk2Qc0ZqKMt+82O/N981B/WOJ1XlaLjTNA6CqJ9aBNYoxf5nf2OTjFSyY
WR09gtWYDyswCRMcFIMIbbyWz5nuX503gjHm8t0ihH0bTGud4vYS2WMAHAa+
ryRW6W3fpTIzXPDiwx2F/C2V/ZNyOdfc+B3xQrVEVVjMC+v3DKH27dZ8bO15
joljLMYEUErW7RqZBExt6AZH/daGOgrmqrQAT/U2z+O1CjTJJn9++MW3tkJ0
yS40VTvWuyYh5bWmIEcnbGKXmAIuewZ1DwXX9NoeOCmWLy5fj3r8MIlc40nR
CTFtN/QeyUhHztIALYT8hPunNeYvUiB1d5l3YHwegDh4zkGVRNniGxpcY0I0
hrhQWvHnszwbnORHLISWjSD+FKKEqmnCEGC1JZb/GWzh5I7lPUAuVSmiI/y9
iQmh5BDyk0ueO7cQKTYWuoyXOhtFVGbDy0rznCm4ahJKfiYcG/xHBfqe2py/
cXKd+iKHcIcDT6QQtBvh/xz2mGGYl8hIfkbnTyddo41W8zn6NbWH6pvv75aV
VC/kGG3rL7mGa9NLs4CMyDJOndz3xE6sxizbA24JlXjymXsHmrXWH4xOczLL
18ybNGr5jGAb2rWmjdoRskAUtmOmL4xhU8UPJw+3FX/zZRgwJFEEtyYJsXDw
6/P15bfDx8ArCEVY/x6zGuumnGalFkgenxgSsBwU/cyqCEVfgHy/+O4RbgYO
AJqJSC5twi1hQ2ZGyMkKWpZsJrtbQi8boJ5Lwoic6s5puehRiNlSCTzH6WCd
J11Shnr1mz+F4vRn2BcXXkXEwRTJSn7O20vcF9oyRdexcRs2Ulw/aB25dh5Z
19TnT7NzsqATARAv04xDTqxWfkAlUY1HViv6BN8NquJ25wnHiXBCzhnik7/G
3HYkO+Vin/SPyJXj5A6UprOJqCRzuqEvKG0MsGtKDOQcrdMxdbkUAIuvL2v1
ocrPhVIDS7a/2DX2Qp+eWXXhkH3odhwpD7sEtfXGqBQX5GAIQ9pMnaphX4T1
VInByhgeiIJEufjTrzuXld5yXh/B+ylA9zhH6TfGqMdE7GbFqvDSmqDvOsiI
N2pDL/IHHJcYxmOZn5oHMXBwkwM68ei081ORC9d6LA8p6Bn/Jlh+E/yfyPDK
9eloLNF0ULqvGE1kVM1CG35ZqdeFBqurKlW/f6v842wDcc5bS9NQ93JWYlQi
ugfqpi+iDZBiwgj7UAWkuwGGsbF547UkQVXC83KzVOp9qzHW9FNaoBnIJXMk
W9BJoAie+/9qW5p5EnN3oE3zelFTB8gAItUI5ZQE/srdBFFrzM9Kqsm3J3e/
VXtdffuRLptljVdCYCz4u7VLbEESbGwq/h+kCugg0BtYdVqb9S82Uly7MNJE
eZcRCOT5w7dA+wlCGgpkX+YUQD6fhhUnqZzKz+tdg9ugvSbVRXEc321DvlSr
UwkdwTZrAQ2btkbVEb0zGN/tK8Q11Oldfds1gWyzXk02wr3t6hEwXeWzWoXV
aGvCofgNIU5BqgsvvKS42yFQXMnCxpVkL0XwzdsVdfuUMfqs2OexUR4ynDgA
vlCmvLvcJy+ZJe78s4mg5FpplQ2cCY+cNvMkA+fM2E1NhHByhiQSMM1oKMX5
PAZHONPbYeF0I4OWjjBAzaA5vZckFOww0SZVcUeAFFVXMWbsxIbpPhZPcmaQ
7HTHI9EPqQbgGRGzeQqDUdV0ANOku7c4yWdSO0AtNG55mBaIWnaw4WtzHTOC
gimOK9Yv5WS6B5oCLSHEeazxgt2/BnOTfxBsA16T+yoxQcVr1HTwoc++YbtX
sl/uCAaUVZHfVORRQUs5L6o1LdNKO1x8d1F/wliaz+JIhfC1jEfocE7/SAEG
RZ3UZbfzdCjrQZ1KfsaDP6XzbC8AorefWzBwOR/qJjMLDnlarjIOghTj+Ys5
uST0Wd1qkya8IhLZf8AnovetyAvv6vCeSqIRt96mxLKgNLGbKaE4hgPn2reB
Y1t3x43THQoOj92i7Kv1N0dq20DRPyOIkWDILRYojJKNt+43GzH+OQERoERh
u9h4aTCqWvvMqWNCCHsAzv9bcttHDBTEWTfLSvhXti0LGSKHiyq+qRn8F6c/
zFZep1W7VoBImpCpppdH9t2AdXE+I1U7ZnyL11wj1Hv5bRI/w7b9lN16d9XU
pvmqXrEtIYPolMkNn/YavZd5K3l45vID+fVVz6i46CdxcuJeb4IgIbfc0eL+
yebILVI2JyrMtw3oKIsW8RoHjOEh4hJpoeEHySSLKtB3H8cqkewr9G9TnWtY
uNX8pskLD4Xl++DcdbJ0WvWyw1konXNJdnJ8PeTx+3HaQjLkNsPaLmOnobOP
J+GzFTbWGNHC0XgZgFvPMdRPq+iBwaPa7Cg9QRjbyVS+glddWiramU1ZlqWf
caoRCuqWeSUgYVKTawBZtV3TVKkR1dHpMyfABd6FnOV9+FskU017wsus9i9A
NqGqJeBwAUtW0bq25kFW4P4c+TtYYqPbZTnWk/eC0SsVOSDPpbQfynGdcTz7
7FZWXHjVpAWQ1ESvavhMF2pt+uNX01sepFwR/NYRWLbHMQ3jSq5ZVIExqB92
sGPnKUfsY08ee6m5XmHz/Lbg/s6T/ylnKxmPRsxUZOxG8KtaxSIf01jKBIhx
nQkuc2hGz4vLCA12JmDmFvZYbsYpPZoug7Yun/uyBp1JsNR06YBslnw+erUI
zPolMNCd1Hd9mx+P43z1L7MmMRSdghIOH5voN3RlOxJIvUBvINpJhV1i5fpZ
VUSEl/VrZ0ltBSYve61CEc/PGoJnXSHaE4CtX5rk2gPwvZ5I4SZXrpD/gmtv
c5XrXKV4fiUD5z4Sct2XDsGerekcve48Kuo42HvSZCvEcf33EadmqAVgBA/1
awG35Z6A65NBLTi95AcuwYMwun8LcizmOuUIe3h8iyJWSo+HPo9g4PcD1N7O
P5CYz3qjOnWcTcL1xWU7bD+CO+5mDFh1JnulOBiRFxROhc0hNSZiesHoPtDI
YKfKBJW0rcdH3szgtz6DKsN4S+OhQBMiHzPwJNyUfoUVrP6CzQIvl0Ymy98j
GJlgpl56qmfp4cGLh0E0OLynf82wti8CotlMGVgwQOlKf+XPHFgk0lDn9307
GSHDt84Uf0akh37/WOURWc4q6iYJ0uKK2AnhT6TGMMV0zq8hXdw2Hvs9hmfn
pQBAyiSLERBGb+QXKaWVZFGh7abUhs3DVLIs7FZYokcPJCrfp+DFF6M2TIDW
4BzU0JbYwa21iNryJ/Q+u3JBJXm5iJfp6np1fbSaczR3bN8ewpp4GbFR51q1
NOPWszAepujjYlXRwQ9KqgarCGyt+ArgcEsHTI2l3W8oIGmJ1WMUuIbDCgly
30hpkyxYU58IxQOJkEcu4wVmU47+kReJSMwF+cYmRffYY+Q6QbUPhsn37RcK
BuBidDVX1+JzcxKaubEtt0pspTON7sWbZrS5n+DGcYypgYi/tsJM+SrXHhqS
WLv9Ki4Of/x0G7lD7IA+fdrleWKPxDCh8uned68c6n6M8FaD40oPFaapjIYJ
GoOkAHq1P/KdfVUBOJg4zTQlyb2pXbp6JuSNYSQkN//BqBfDT+PKxGCJR8rk
a/SE0D3llEsZ9zPVHjO6cjAz4t9zvsNtqobDpkvxT89PyQBqmE8NgF23k0uT
wN0PYwZSgW/X/BJ5uhgA164f2y9lZhYGZGXPBqqiL+VSexWJU+UGndiwPy67
oB3lLfZIiRedbJGaN+1qqrG3QFNJr7KS59xbrSpYhmER9TzP0AI0vXS7XQ7c
cwZskGtjeYO4GjJbNetfJpcJnfammy1iAnVN/gYDSGsmZGCjVSQ++m6eH5Gx
L2vtEw5szx/2UxgzsP103SMKjNcnYioVKs7cv5BupWNTlPgPt1+auyCdcfry
JXisEB2bKhcB7tJMObPRCqyIS1YWEHHdS6XD7CNErqriXmtEBUUi0mz2+Rva
uEa00NWOSm7ck8SD+lhFxb83gr9P6/Dhvretz2apz1luVaHXD8ZbJUC4pUya
sTVmn6wg/iOZl9mWmg6WojP2UGBxxgLIAQCcDcFvsBJrGWtjGL9edzBO9RHU
m9isnZYPmwSfeOx2mbtiA4vIuIJ7wXZx9GmjTx171TCmsix3ohxd6jFkjFv/
tmXVR0UV2hm7x4NpVpHK3F3NYJdctKP1mQ8CM9vrmDq0tnTITN0ptzlC9XsB
4Z7gF7ZIPiQL7zB/mXNwnYlbZNZrX31G++5dQDzEdzj7vXs+JUH4kV/LgTym
pSE2ZgASvVomS8QA/PVBL7JNdPZCV5pm0gnzjAC+fss32GqTWrJyrDWbROeh
RjA9VsSs46hzypTrF0UNzHWJX5Uc/m8FnxcIUose7vGXqX8Q5JVaOqZmUukg
aC/lTIrU3hKUAPJ9u9EZFspGv+kAI/2FTTHoLydSuUcHiGYQ8gGg6pdBRZLx
Il88ssGAtKUZKcVRFIKygYcvVKJspG580si+LjyMQlAlJNHl6iJ+GUAAPKeB
Er7OTrBvTdXvje3djuTHo0sdYlP1JtqxyFu4JwVqjgvA/6VhSObGaHEusC5Y
Y31eDJghH73B+2h1RNdovvD9ykPw6yPOPHels0W0i5LzeGzoqahljT/UFPz7
VsJOvBKYm3yr7fzpnQ9PPCsDcTEeJGSXzWvmEc6wFTVU+SPJ1ayPPuH+IWIx
bX7S7G5MQy2nkrhjUnXNnAznLf+ul9nRd8R1qzqvzk9JH2eMlag/RrhOkVAj
mlKtJqgwYmA81PjVyOTOEYzIBbw8BP3o8kvKTcP59JvoHkMeBJYudQlGo9QM
bqwRo3w5Z5LV6opPAxmU3IeKjuT5ys3YBZmQv/d3G6QpWxChh6oyYOS3sT85
qIwQ5cl1uIJYV3siVOlLDrjRSbLT4BzAXMNSUEU2yHBts/FjC0luvxjRReDU
OKMMv/4yrtNzEmW45/d1D9Lcu7N13NZzp4+qNdnG+T4Gj/Aha6DlEdqKST/U
lEVL/Uq5J5K+zG3uJuFSb26q3iLIm6SgYWluPc2cYVMXs4Se9n2yQXAIq42D
5pzd5TC3siNomxWXn8AgQ6vp1nMZNsX692/hWoqT86VuTsY6dvu436ws3qjV
OU5CW1CZNYZ/OuzEmhYPMCs+8qfSF+vRC+ueXrrxOoFi3njx6mENZaO5eCXK
4a4kYVEAOXAhOHKUNjmCecf3egR9PQdZBJKnQcEVzhc8pG1sle7rVd39u5OH
ipmwv7E8KktELXf47TGFr/mfROr5GHNXyaKGSLn9XjVDOcZnVDlK04YJaZk1
RqNgURgpFay4LJLTcdPpyMKOzQ8becilKsJRr8rtx30O+FTzJW6928OCXj5X
Vg3dy4hjTJcTKOHwGIpESxjHrgDzFSoG5cXQ+E1pFHf83e0zw63870rtngSs
OV9NQPf5qJurnYLGTq2bMcjh8K3IqYHueVHbkCnnzPOSlkn81+0GKIbjJqgF
5A43W2X61/Bso7HQ9bFnDbkYkCxK1xx6e94eecXxMYWTvzk5YBPGMYU9FKah
CdnkUR0zNt7wqf2qN1U/MPDHtkmHmcV94/JS+bHEBv8twS7mYjjqdB/Hj/zt
rKJxUihb6E8uohG7QgDJgwrFP8x2ey2z1RIK2HYajuUnqDtxiHMR8GeNiS63
rB5VF0l9gAOJQDKmXWVW7RqsZ88UMkKJr85PB+FzEaNNaertkBVWL3Px7+Ko
MabvEDra08XOfjdtj/bHQ9Eq29/wkbD0nReRW+WWZC0bxSIZY1xPEtpuXTMF
RGYBjMO8JUGQYW8gOTEE5PLUycyEK0apqCwEp6qNxQBVcX4NhjpOXiUIVtnX
ZN+3N0XyQAL1UERYxQEqldbxe0vBV0lJ4BWWOab18cQ9p9ZGlO0iVDDjbn5L
vthHbKl3FPLJocpWYxFKFzUHTkG2LUnkrsD9bRtIvkrSAqiuCJmUGaGjG6xc
vans3orad7mxUEtcgyInEXlU8YMOJbpcGv3rH5VrNC7iiuM04nFT2+ELGQhP
UDEWYyPjBnfOp0uBLOTAIbRBXp8JIwYrUU5Swv98A2WBm2mgL5FagDtEuvS9
c620Sn/aWS3RNqu0O+V3LVoRx5EVOUNFIj7ZTt1DzQp7SW5gJ49vTrk8v+yW
MFwnI1SH3IcNJCfQvPH84C4zE4jB5z6FHYqHiB8pQrV1jbz9GsKUu5mz90Sr
sY409nFLPpTzCgui6X7/urBxVvkuzvu6hd6WoeaE5spVftf7/O4YwDlMbCf7
BcuCEHuYJ7uiI4exWEispDY7zHG/X/l/iKPWJCyFYPkTqjYvuoQtreuYKrKR
19E4XJgBKpCpWY7ewTTpJZ+UMLBAbVi0RUOhyVkaJRn4nepifAVhpUZIc+Wi
NT+aP+9AloWraQpDrETZk5Ewhben7ZGnX+f9n14nkX9ys00zEtVh5Rt/IfvO
keLmJ1bCH0Akq6ZmTOHvcj92B4mzDt5VizSc9WJp5L8G1SF0QPIe7G6feuKc
UlKrCDzD2kcTzSGbF6Ecs6hs9mKzPvG1VWyFSfJpOuu+fp3hxlMiqVSfkxw9
EtnaTfwiqJgeCiZ91lTjnS5JBfGBK2HIz7HfeR2czQFSVISb95Ps1YgEL8di
IIk1W4PXsa1v3AuixPkD3d+yJEnZ75OwElepodQP2Vy/gpK5mDuaDPP2BJvP
OsnVMxhM3cOaltJLR5/z3Rv/hIMiSMFHnTmYhQo+J9W+bABn0gYnhfmMo2Ew
Ai4BxB4/Mm6i7SqrW6tvAWisc2KmrqpDCRpiRNjsSIc7D9vHrj+SaYWFaXo2
dkvakFfzAzZyTOM8PU3Px2bl87110IRDHybM7XJTUTYcWVixHet4GAqDPWny
PH2RvVsTMVhoqIcBA8y38E50qF7wy1QMxlSQiugbS77BxWmMfDKRXWMLgDXp
TI3wbrV2HUJfEFsPnD+EpGa5E6aKnXGFB/VAEsuR5MkyqkUQqw7eR+0xWyjq
5urxp6n+8F6kzzw1CoaFa6tjqBLCLIkcT4wqfWIiBQg9GMywd/wuu6rvhDuR
RQatl/Gig85gmv515bgBTSHYDPTmMawxFeAYuRZi+R+s0e4fuI/VaVRpcEIB
I8sWaWFQx74DFhQ1MNE9SgiE2151uJDTZNK6dnmkK1H1ykSZFLwnbxYWFEbC
PRxZzu/3zG+dE8j50h2HVgAXBRVZ3euUpQcRjcjOrACXyjF2n9PZnnxA3Knl
aOFoT0LzYWuRnbNICjxMCx1Gb2k/Oqf+ahZGDKuayqAnlHzn3sq8zmarv40h
t0GGlu/Bp1nb7q5JbYgeiMmstGX6rJ+DVgf2UFwaDXV/WNbnRQfVmO+pnPv5
azgW9tVjwfE/q0mXA8V1VXL2ZsqLn9ppA24wp6raxI1DcVS+acnUCKJdU2WC
quUjhak56ROuRodBXLk+C05zcW1a91C9I5cdypB6/LES4pwtEi1zpZXA6COD
hwz4pJ2Q02C7attkRLuGR5TOPRRzcrd2BFsMGA16T6y4a0ayNp+UqI70UaVR
FVRF/kQXYulybrHWUtaC2t4KCE94UqXk5pUBlKxXL6l9VWQs8RCznN61oJaD
ZTjutM+qgW2zBfMGZnTWZ8dnHUx1st8qVYcPVR0MdssAdsI4bT6/jOJCmTYR
9GVCcrJzrAoYVTxIwy3ErOXMeoaHmJwXQSYDnJ6TfpvFltCUVQWxohaQQCeZ
KOwnRx4C35ZaQAeNVxqjNRHWJAKXUN0cb4W6W6iVgAytVr/zQU+VfI1rfLT/
Myk3fxZyExF39Mvb4MVxrTQ+SbUq7hKY4YPa9vZyybolw4Iu0I+nfdoBVCuV
YYNN43uy//dlabG92YTD12pecib/jfvSeVP+vHfnakzYrI2oeiwX4u+johNR
7Lvx0nuRReaOf7id/yIRp53zUDxwUSOmdSD58hOsEj+tnLmQbOSOiX3Q2G0J
On+WPcqMPgV1qJMSv64nxO5s489KzCQidEBAItsvv51BXS/sLGw/tlHb9RVH
dVdZarIVc9Jcazd5WgRcSZKv8hJYeh8aMwNDjfQnQXvvbIDW/79oJ4Rt3J+Y
GXaBz3fD7jBz60xh8wpDwCteicfMC2oDgrPkNjPFo7M2F/yOTvNwqlSQOuj7
u+eAFRQXxZpsQOrgThsZgWOeAGmyYlDFL/VLu9SaFxq0s9HAdhoklVwhZuBL
tDBqGOsGxsGeOk9tjSl2IRsKTmAY/G5vfACA1+Berr93xHRLDbyxVQQ3xv4G
k+zGsr+f1T5MXgJW3vtGyHHkngUq2rXXvvEvvlYsETzkMFQg3NnfEQx/W+Gg
wAcO4elupabwzAbcQLDT6THxe+nO7u6Y8rM31X/ZLvIXlFoJt4O/VzVgBoJ7
Y7VXvvJgwOWOixcT45PZzEzxMHAoJUm48PHAS7XbPqJraITZkc57QkhOn1Rk
1w4hUlpiKTVK4ER/txFKWgZKGnTswzhaIa1F+ImmHWRZTXU6a/uy0T/LlPst
qaGnuQv4scY4HBpGsj3jI0oZcBZCCCqtUCLAdj1+kwekYOwhQt58dIXnfexw
s7cftDlJ1FNEsLCu4niLHj9VI6iE6ve99RTe6PFTAAJkhtZu4MNqrPurpxET
+xr1Bpq2vqE5snehskhvuLhL8PXvE7yg3VcL1xoLMJy1XUuwN0K+mCSVL3t9
BmrkIhr/A1fcIVQrwCLHbxm4Pgnqp5QpoUf75tELqGpBZUnx95O3JswDBlif
AZpxiFgVG5sAE33K9IC2+qoG6vUqQdJh9jXzmDfdexaGgfZR3mBXBeOacMyN
15pO7wUh1AaAOWnzyjWZb0rPxrQykQBmui/4xYNixGpqQOUzofeQivbDutV0
NkCfSPjmA+supuMwMc83ON1VM6hKJkaBfMzWAQbnLmxlpVMLxJAavvJlbUD2
YHafl1uaRxpqvDYpKKoqnZdswf86BDl1BhJ+3JuFxUY4NsqpTw4Qk4hqK5ow
bAM5Bs6emGPUpvfoofXdUXqiLLKSzha3Kq5fqXmRL/EFB5FV6jvxPPUV0hro
JTjciiM85FkTxhRSjwYV74zZIgwkGnghySJYAr/IsP+AiU2IFtxdEw8wN9jk
OWf8LH4Q95+RCXjdXC7gnudiRVGuP4Lyz3k9dK9sm2JJFmWVh3I/hGi3AKCQ
wIYPCB5d5iQ3HN5qemsznPAynsY/rQgEaSbYclNGlb6STTVne11DcWZiy4kM
v4NEhomNDTSE/2KQjNFST4wX1gCDIGoOzEsljpu3s6vmNxUdy8iTZFv8E/jl
e7wK4eXFlXhiAu1sgDvaNo3BakRJSsl1Pbvkji6/kvdyt6gDupg8NKTC3yxn
c2LS4NpvcORQlbZ2zjY1t599LYCnXFryaGw1HEfwRIF48Tm/JoIkbCZ5ZWto
KiOJydUmEQdptDhr62BlO4FE9X0sLHi6QQZtlKphHS/SszdVm053k9OG1EOh
4vSbgPlc8H7tIHMp05l0eHFGoiPDmYPusLAPsuNTUgpu9wLnhmgu3FtuSipC
MzKh0coDrNccIcmFCMxLoxUkzcAavLuPl7vv74nucuF05rqi0DpxBc1wxe/m
tbQyK6MUQ8gEcDS0Yn2JdO8RI5UZxcIsv5YRKbfZs/Z02EKXHCmOaOj/Bbcz
pqN2mVFpOmVGIHTukWvt/TF6D/srY6xMi7AQt+7ICKEUqeQLrTT1CnbxDfSm
jE/cJY24APu6S2H/gtEyu3hGvMpYLldeguLmrkLAGDXK+wkYIx5RwRNjg/Mo
fHAyNC1OO5Je2+N7+Q3687RxN777M8KKUDfG7vOCJA6VYiFu9ZCDqtUjN3uU
9/Baj3L9cD+/GnX2uzYwpSfZA1SlNAx8JOPpmc4i4fWxCVYC6CfH8uvoZiq4
VVAs3ThBz8Q+NS1XOpudVScLrMXrHZ5b2n2sqUU4bbYCJFE4o22jlq7xlmhc
9P5bXZq8i7RzPFEwgzLOvjeXYMOuNqQhW4xVfiLwpINohfz3VFJQ3LzCcvbm
I4ZBmxBulH+k7FWmKujyfp7Tk3OwXHwvrLr0SGMsRUvHiEu3SWlMGk3S9cZy
/SnxdWcnjp9CVMlxKer/JZtUDW09484ndvA/RKn6o9cQAOS6QGhVxy8vceMh
efMR4g7ji6f7xPlcnvsN67ajeCpiN3etRx5bW9dZvGkSnW/Y+hePQga7NZI4
HcbeVE1H1tcli6nm41d+raN+Slnrqef2ppEcAKDjoS6z1Fd4LrYlXotG1o4N
RcAtw8dAFkdQb7KuvNUtUSYqeK/EwHIrmvkArGy7q2t/KZyMZ54+KkVi+Wd2
ZnKoce+T6Er7RGGYKJMFK4NsWXJKYlEhnIH9qK9ad4ZTl/IEEufBgWLwWK3U
CxE8+TRngQWtJsTNsGYW/5sJf6fouhWaeGWIGiNF1L8+M09uqLHV6h195DMW
FaM/B3dP364Jl3gGVHi9ZDD6w27+NxAErv/ehlmVW5uNZd+x0gCWQLFnBUHl
WxwQwPDaejzEymW/QUht4c1attBdGbpxe7WXn2RjX9/ruGGiP7SUW6gBltTJ
kC5xxDAGdt/GQR+160qUOgoROHT6/aSEfXEsSvsvd90F9mrXg4yeVC1CAYFH
gr1qnfv2qwp1vuG8GdhDTPvxu/j92h+sTW8Rq9gR8UUZ4rm+9N/zL2Fw+5H+
fMb80I4VAnYXVM4AlZI8+qyyI+q/teVX/7gWZlR2IzhIOWrC+5ej8bRAKzI/
S8C1J11BkpNstNu6/MA/sSzrIDDVUAqLaGV1NMJYi/CO/iuf1h6cn+s5hOyL
CUHihJrU/v9KiPefmZtsCaoCMgMt5OF7kRov3Mi467nH3HkvuxWG+gSpR7Dr
GocLf8PjlqZ7v1R1PcyYrssiNavsdflG31iZcFjbr3BkYUi6ebuYbRDBgThu
CqmVsMrnRT1ocQqhCvcAuDVBw94POwz51p6ZXGyHrDLrG78wRnuzJ/9dDvEJ
ol0VuhLDpMX3BaTouKTM6AFOyI+O7jfFeZ8es2CultwnH86AZkCSv2beJEfy
9WzNZVaPxvBuarzFHiL8xpv4TmDo0vHajpPAnMrJWKAv+VZcw1ioEv67BWYu
J4r2+yhf5bRucOzAZRbUhIvLOHUSspB16Vhc/MCM6JKSN9ImsYnpJdEA6AGY
Sr2+Ac1l9XFmjSF7N49/foK0+iuNJTz9K1jwueOQHLOcwUCKVjyRsHyuijnF
0m1OOv5SlTRPTX7DqMCrdeH7NGnzU380rP2JXPNxihY/FgY7UPhIB0TVlr3h
RMzp8RahXz+OGAoUuqOOO0MNJitoQileGAWE1lJga4nGGjw9ojtsg8ACV8zF
daW7DVnVT0jb5Hc5ugYnFyWyxUxRoSbA+lXnbDIjB0Pemr+cqJMvtC3BxaDe
ZPdLlNfkTbiwScbsN7ozDPS5HS0XMXULYb0AgEEWVTTUbcANnNOyW9iGMJG8
WpodCkS3SwVnxZEJla4hsG5Gye4ko+WfvdeII2hsniJ4pdOoVQ/xm2u2bQC+
fZk/fUO7M/6Fx3lznuW4LyRXD1o2jbJJOMOSc2qkkj19gVtYK+tPWANdrtIA
rj2sMxzVEteliNx0nEtHP7GRPI4TXVuniSAEoz+kYhR/CdGIUwvYqd/qvvjB
nMxgLvfIg8eQ+zYrA5JOHdNLgSOa6s2ajnn6Tnqjx5Rwf75ktTJz3fPP59dc
E2aE5rGAJxO0zM53jJsbdQlZD22eEqASQ186r8YmKy0UY/hq13agLs72r5jM
pl7bHBW5977Iydb3fvdXeKOg4b+OeXJM/ZCLlU6vtAw52oVR/fh5pGzCJ5Yi
blrCxjw/ikxL3cXSLvLs3+otmcSV+V9oPjR69PVH1VRTkpoJINkDL4r4Ef9S
isQZ/eHWH1qaT3iES7xKoV3Nkx/J30je3Be2/f3NR4i5mXkdjnid/Dm+x1uF
NwliHj9F8YfP5TdDSTeDlGT4ozASvH4UlvKci9YnuQAMQ65wuKcAlu16UY2p
rXBkASggQigZRLPqV8TJwUbdnNJNN+LndOYcr8b0SvRurNKSWCwEAm5h6FIV
p+UaTZB0cSi6zzgfsrF5f5FBGTEIJmOcJczIrgnJacRWtRgk1sb5rIiZo9qB
5MIcoOl0uQg1KwvXBGiz3L4E0jBFePUKtHAK9QKGTKMWxaTwtvXbB15r7ufo
Jl3HWUIrtccyFjXs4o2T7b76u7rX7H+I1s9l8JykADmlot1ociKL1qkgnhs5
FSBGvNDHsyfDvu+MTcLysLiuO7tFiFctRAo9+yvOHXTd5dOGIP3AgAdAD9qd
Cx5lMNIzsro5ep4VYwkk/PjcuIJsS1tK2LBxC1w5y4cFilJ7C7OHjYOHIVl9
Y/P1QprrMcfNFqwJgk7lPmSPBrKFvofFzWcFfPowFAd2gY0EmKxkku2zxO8z
a2I6F9LG3oIFtn9+2tcihNosl2wDS+f4GGCWCGjXMqDrodvXa48m6Lke/tlh
GGwV1eCwVNJlSDPG7F5t86oyYFGXNcHcX7LoTH4X1QselpL1VIW0qnXlu5Vy
igbGkY2I4X+hIfSRI+09cYRWhPbhHhriMWpr6b4ZveJyy9yFh26zlErg5u9D
CdturyNLEfXPUAoOETViqwOD8hpR9zm8bj2ceEzjzPRvbBlyVXJTap26CaxO
PV2yzLGke5IcJmVgcEgHZ8/8lj73FgXnidcxeqiuZpWpKKIbD4LKcwfU8Ekc
ncHYGimZAY7up/cfi7Z9kr5akqwlZljiRa3GuamX4EIyo84hD+lxUzyh229Z
1wJb+iLqwD5T8eCkyXYG/5v5wNYSW+tEuX21H0i5Mt1TWd9+/VB2JWinjVzW
wAriyggJSc8H0ICPL5Fh3wOMNvCu/3Ip7UZw0HAMCyHKrisx7gjDs2IHvYG+
NgvU9R7KLB3gsb5ZbiYICbAhXIhVkvR/0v/OWUVheSocMEBbWhVUWFLSO6Ad
z3mdq1Ovg3rnR+nd49hRxOr+VCi6KLwiMGUgkufHOZ9SsudCuqxWeXwQugrx
uooJVNV/9MqfFdTGX4PXMxfbt2iq2S/m9epjZ0byzlzUAfJ3NcaKRRIOMpiW
B3r0y8k+6ivOEr+3be2cmo2W91PGfOYS8hMjI54Q/LrJ/CQeMLwM26SV0diC
oi39GMPJd/84KCmjJdL372777/qH5OZiGLJUbcMpk/F94iJ8pfaavhgoy5nN
abgzIAAZt54jLO1R/nWSgKhkcz4QT2EIK8juCzkn2HOlROIchn9yLDsUNiwj
Ge96JPigqeH9pkQb1+xjcPbUnyoJVK8A3qtey5L2svQsjiVyohHGFjsX2VJ6
Z5CwXQ08fCLrLKQorV8oRxpsOag6Krs8Zp04bQBUScWIglhBhz0cUSzrxbNG
Stqb7PQiyz/HnaeCyJQZJww+ES60qCuhEDXx0NB3vZgMZZs7YjkLHOScMCZR
UxzKs8OizyFUeUVMljJynB7NMDH9G8mVIbTPfjQl17EoXHZYBo110wqQuHIy
MLqlO1PHSpCIkHiZ4ilKjna5D1/4KULq1tUS4uDydoF4x0bgq47NWzjisPTV
VsINj62NOeEW7ft7QxwSd5gIIZvlxnQqVrPOBskVbVBKL+qBMvNKlEfc6hGk
aVCR0W7Sad79NVG71lXTxDnJ3LkdgEquCzzIuypbk1AJ9euW6kS4Ac8GmgrZ
bm6h05fOwrKzj/nWFeE93fwoMQdd38Q5IxyKuMfORfi/GqxLK5fST2N0qfXU
PrOpMNACVoFc+VfJiPk2kiGxzHEGxJHGQH5EIr+AbroSXfQrQ9MNg/TcLu9G
r0yFGp3ZAC3EwehLGeLJUEA1X368mWi3xQ8ixPGjsl62Gj2YEsMKFWu/x/de
NBsdMzI4TiywEnRZGjR3c6UQMXEdv8FcmDsgMxMA4WhXXOQorkcXfjU1unPK
4YeRAgWfFiUZD0JgQoEGmnmDWBVM8hmX6q5iekApR04U/2CdjerMEVSVmUo2
3Qwzd4rb2JIIWHjs0wkGRN+8epKAV0gWKb1jNh9aKhiyweIXRAwMqvITPnxB
jqhqOGFAxnNa7veM78qHxI8qZewbbHGGfMdzUezbbRon9Q67pzlC+/2Gxj+L
dPohqPs86cF3hpIGd121og8fy6L80cLLOhwHqIGgfHxvzKl3vxM1VTU1Nnk/
yU1mAf1+gFFBKbgPSp+pRjDy+niI6mtT1pVGaYQSm8O0R+qbaNEOC4R45xGR
LdqYMQzGmVTlkPXUxnljHEdu0X6MzAHTGTqR6+9ZuUBbu2k/5FICsf9WKTDD
GRCS8CrTQuspaK0P4nvuRGbQnN0nY1N9ZlsNaxSSW2ivGYQ6Njlc5GSiMXZL
tTxa1Yiqd8FaAfIwBmLQLslIJ7mS39QL+ukU4BV08asdaaJFsNcxq+6w4IdC
bZ6ccRllfUCTQENIPHLCX4sSvPCtss0tK6Fz5qUEExFhfrxAP6H1dPvEgFat
Me9ybbpOTyn4Mvaqjs0SMlJAV+GPqmPngHOON/eBP6RYedzrkTh5yAHfbKj7
CUjFQeJFjc8dkBCLwmHHRY+YZwRhWqWUSo0CnUcBgTnwNoXAFDVvKVw4iaZs
NSboekx7s2JZ+5KD3nchkTHOpSTWvuR4WOiewGfHMnAZO+Tj8/Ph8v7JljtH
kb2S1Co/zdY7TfIavfddHOtBFIAPWCtjHohG+EW8dy3FAF2v3QIOvnJEaler
D9Xc92n8ZuXgReCi8HoeMw86a75ZwJawlnK8Y4wn2wcOEnHvj6rMH50cx0QB
RXM0JDp2vtGOxv0SJ9H5VcZ9qAY1dEPeY6zeNSYpdukZuTVCcPF8/uH/6STO
a0xrpMMoXGpY8+hwymH5mkViuKh3DfAVVqzFdecXJLvjwIJ6xgZKbUPHzp9Y
OxL7O2D1EMvQbCkFIx0VCRbx/CwNYh1FYCyvX484POCTJhNqYw12hbDR8VTB
/z7o9yMfPgt/k+mcqL0SinjWkJsHJpv4YmRdLSem9dyfYS4+00kIN+QjPlpf
dSvmuyIXIicYE3FbzngxUysHIfOwuxjoOlLXUoF7gT1a4QKdiRRb5Uy1AKMv
1aLQ3F67NOiKzdRbRy18LEQ734x0mtUJNP6D9n0fRC7ITxCj/LKrc5ZD3fXf
Qotu/nsTr6FKzlSrkMWUrbe7lML0pUPqPgj6NVRUMqDiioMWzhZNGvX6PsaF
bNNnt2kw3BsEFRRqi9QJFJFtk5/1q1sj3TT8joGa/nKCkDdeklnEcIAZmMPP
PLzmpopdrkdyslDOREygj5OXNy1YehTJcvQ+sXOzG/oUTA1BjvP9HVieNcJq
wygCHoKV0KDvj2wxFmU8fMIC/yKn/ex0mFuvN9Tq4evpm7CockxVYwVPz56+
Z9gE/iD3LMWHGO3xDAhiHAuuMws0AG9sXHr/y3MahWobg7DtUxOALFds99AJ
NrzqFhkFp5AwFmHO4v14oaq2gj36dcXhjjlVj+XwprWr2JxW8jYovAvrKEKR
iw9AjHIhGQ1cWm5TpkZnAR9H7pE3Q3jAlSZ6/FwNudZMuGHGVRJaBFJ7Phno
Z8Fnm8n1UzXNkqoI3mexjX+Cou8NXWcA7vc7i9qvjzBnOga3TNq+hQ6qrwRE
V2BzKfKUhuPQ84iqaI3mWmkHhAc2G+7TFc9Gzla/fPLzHJK13oHBcTTLZheh
CMs61SF0y3ZpWDSBuPC1Pr/JRZKBHro098T2aOHb1c2wJ2MwBJwcaN4gAJHZ
P/hY8fDWTswGR0/3V16zyNRpBOakgqZSVnD3mX6+6RlqzOW4tI434h7bkoWW
pfy/O1ZQS52hQbubAPON7kd14UglKZRID49adpTsQme/tWaB8QbO8lpJ/45w
3N3SSM6HiJWdOC4LDpMnUGb8TUqL/tBcufGY6wxZ8U4Juo4zsxK04xwQPca1
kznt9qPVnr8tI70mQH15cf2xDTFvuXGvHvvzpOUh2Z5N4BKXdS4KpJlp8uB/
4EF669cqjRTO0twDjvI1fe3r1DCmMoO9zban3OpdqISwoTCHatFudTLyuCJn
aLNyFbAJ46d973sBFzmkZwEr8nCNUyLa0GWul53W37CCOAocrG+W0Yjhf2Js
8xc6YkVv/TnGmhvPu0MwudPlwQMHeLlEjjd1PKcZI8GgPs7LkZh6t5BeYcQr
8F98jH5JNRf1vS+/bTcuPW80ZbNlQyWSYvciNco2HsRAT+83YdIYxgqH9Did
Yb3Jpz0JEb/VuJE5w6OTy9AtGfNiTWCxczshlZH2pepQVCO9K2P1Pb3IZ6zP
NgP9Co0yxW9aT99/4piuxzhVslYsa2XUO6i62HiMKK77J4rioHP/bGp/Oj7k
cZg9dPY3TWPETEiXooqusx3AEbK4cfKvb3AG5yQyJbuBfdAp743MmwN4y4ZW
2Z88x+kc2MiCbn2N89a3uiM/RYuzWjRUot9XY47yEtB3J3ErmBxX+q0w46ik
XeHCogIhWQ1rj7gzcVDYbppx7HANxjqHyR58Qodfgw5n84DsAHD9r83XZ+mW
QR6gSVtNAhXr4VzZIqc6ItDF2ZZRigR5O2f6Q2AAtBawNNpee0bVdzIlWm3+
KM4Yp2QeZPFOk1i5xAwjhJ9RsLTT6tz7ntfVAz9TJlBsRxeqvS7ESMtGsf/p
Ec9rwHO7jliHLTAcWuYrDxj3LKPXX1WXCeHUoFIlQykOnGyY767DYX8dz8Tc
odeRxZhpayJYZ+YNd8xLWS0tLVSxjKC9/t0lxvN6Pd48xOSwRgBP+wjn34le
8AeyZSQWTDMhf5sEHy5GSvUwFd7JUL4h+wt5fdhqTe5tbL1RPBBxL+vpuMgS
pCW8tgUsDO7VgXykE7wEt+JBmXeU7bwDuBWTmccM8FvVCVEnqPi/0FpPSosd
ZHqZxzSq0pKYuFIfK2GxJ64VCBDcUe/PLbx5sM5T5T4DPicWd+64BjXVcL70
qFxNzaicpNqNcN0UC0GaY0oAv4tvCwVyj5InWhmuya2f7mzh0pvAuUuX+eSI
qY+XfHauUy2eBNpLUF9fFEKVEuvLDCUC6munHiN4BONNxEjODWHaE0aWZv77
htyUAjM2pTU12doC0kKg6wT9T5EI9OUaRJlyWBraDkcJe9VpW/1du4yoQrQr
kty21Hq2ouJqor4m5FGsm0hkxU8Sjfl7IRf0ybS0baux2j/9T6gRd3mZpIgg
KDfkM9MpvkUXZUKv2tpGC0t4HJfUjA/ihmIoN52IIUlWGOSqc/0Ba6NCWL1e
sKDtRnbrpqbKKt+nh/7yr7EZirWioHHN66piXlIta+Hdn8UiteHGXFx7THdk
RaDFQckZjncB7QwMHWqXHUSiYAxRMwQWtPHvPGmJcWYRzvtgPSzoJ7oIsJqS
X4kJsf1pXa1q3jT7NH/JAygk6TETvtHzXSHPDm0REepzkzkKY3QnL5X8ASie
+xdjLs1wMTOyN6shSRtMb0fQujK1Lpf9xrwug/pRGfle6PATsMYDkvMRAMfm
SgJUhZDyogjrYa6uG2KdZiPWr6myJqW1xtlCZEft+82djjTtmcJZ2p202Ln3
7+KqBlNTA+tq2BuThkDpgpbipn5uJgctLw5flpH1uLstiT6AxyfldGXYa3lz
rkS6+hqmRnfPjGJepgRhi5ezdrZS+lWR2baZ2aB4YmEp/flZUf75eNWt2+nO
lOyaHKq++cXeTYUX9n0e4sv1RbmQmfIPZ5HeIRuTXgp0vl9ff1/DHbkp8Y0u
OQ6Wy/SAZZwCm3MbQCPiExg5oB8aTURJSqd51hXdo4sKuaGnfaQ4vLa9ECQS
gUTGkvU6PfLdfdnodlOfe16eF/LBCN1arx+0OoKDKHu+G5pNYfxt0/EC/NEw
F3+kCIarsX7LKTSAa/WujegL0wDrj3EZLJC5h3Vpu/hU20OdRtBg0Er+HGno
NbboK1xstDP2E6VFvPe61ElL69GrSOgARbj8nVqkbC64dRm14NcXC9zmgkti
eKcYGXnLiOLdn4mTbkC6Z+v6T/G/Z2aTCKf+CaT7rPxpKIpLHv1+voDgXJF4
g9M9/YjTjrXFecl94PsPWq1JCiv0rgmWwDEOgf2+xI1E26vMlNyhBWj42sTx
pBinF1JpPDm9GvBKEeqaFu9vTLxjcMZ0TIgCrlKZSdwq/ROQBBfcQ0v2E+ig
Fbo5S9JtEOgc4oGoBdEuwpYMH3moMXwAm/rEniTI9tEFlTxZgfjFnFw3a8dP
u5EOIQ4dmyx9wPeLKNMtiMSoa+SJzv436eZWuWQlc+RKlkLUYH27edfViVxM
UJlAw2kHl6fhopytKJw33OA+fDBXgERqGYRErR7XfLJkgPbXPLrafe8UWcvX
1LUC5K5FNPaYeXAC8M3ng4qb5SSQ4IPPQXGUGzqIFlGe9hdjSw7YLTP/nv2C
bUHvCKcR94tXb4YMgEYnivejBz6bamuA7taZbVMSGMmQFd7lNjAp7QtlHu7X
aC/6zdhxsxlm74BadVh2CEEym+OHfOmYE6SPX/LMfnkg9TlcPQnO5K017hMq
zWVtJ9CoKnHio7Ook+HCou+4Jom8oxrtMvgfzGaDO1J9CyCjgpuDK1n3igXY
FImjqL2uR3tItmRxbu2/DE+mfeP15n3iCrB7Wve42QmZzlxl5+L3+iIdN6IW
8ATdck/zGrhmlL63Eb849+Ilz0KMLMn2EQqFd2h7HXg411BeBVWHi5ffLex7
EgCGOZ4nGjI1fUgvbMC25sQpDV8ZO8md1+hojdwvRgaC4+wgxID6aT6TNYnI
ZcETW3ya9mV1fO7dvMLbwzcBoqPBUvp1/fPC2EP1Pg4GI5JluFXKUht7ABtK
AVSirwaUezV9AyJYyNY7ocFgxwHTZe0mUxWk5BwXum8TRa4K9e8LTDeLqzIK
RekMk4GBjiErKG7UckxONihYKtUd7LLk7mDoqcWcCnqbK0Si5wjHOjSH2Z1r
vtixsP9MjG6By1SbETpbwQmgtpcV73WTRuaxyc989Ot0kthY5KbKAjTcwuZZ
ke7yucb1r1suduMwdqY+tlQ+6LwNqpMizq0w6H6zF5RWZiA1NBjKDvya8P95
FCp/jo1wXr7mdioZ/3THddMI6H0oT1ej05Vlq9BOYzE47+3ZerqJELf/f+qx
FZHsTyhIIOKflxAVONs70W6gUFuj3XEHQMABaxPmiYRNFyJUmJz6Qvs8pCw5
N8j6vVhhg9MrPAGlQ+w6ZLAINZUlWYjurghDs5QLtnOh4ebNTqcPeivvY+S1
+1kK7cBr1On8V1E4C0agH/XmOQ8Hg0wqOgYpM5Gs1SyoWJ7dxITjLDQeE0s4
gurkXxiVMcTfzj32SxUqNX/uFHOF27DgBrRdy+6BlExtrAY+qpbub3Dkkh4F
cYCT8tCIbNqbPhYNNM3fjc99xXWokWrjvCgVtR5fUIQwfLaWzKsKsXYEo/XA
G5nhkWdz+6tg0uTj222DR3Y/c3a8rF7u06kxgUPV14537wQAwKLYCbHHYSgd
Fbmh3gb+/iEb9VXFzjKEHrSGHW1AGESBPHZ0gOT8816a/IA70suMtfB7qEey
AjHsnm/FZ803urfnMQTbB5ssZcWcvX8gYTzp9OKVgOUOybx73t+m41LiEnLz
ltdBj8echibUMfqv9tsQ9+KtIYSHA/u8qbUkD3eGFbolo6gXJygSW89zuV4a
5TKbDiZdOfvitiu7NejZ3wgBiP1FaT+DrUVf6m6unVKuG6nsf5EKmgmFsx/p
w6ug1pQgwMiJpZW55uDmUSVFYrSSRGNy6cHpp18Uw07SBYu+G+TW5UcPWWRA
z+8fAliaDgOIeX4kRtllfJR5IRckvNXOzZzdxLbl60ZB2O6rwijwlzMqaFYG
Vgbs7G2y8KXFbHZntMvs4wGAGCXe8PjfMXMp/GuNyJ5HB9PrMtA0fe9NScGT
qKvTFQgGv+Nv0DLS6+rqfbH7G2jWdkrnKZHb8oogUtnFdoeVM/DiRLxqUUAU
qEC+VndWImyiPgKAT1+UGpNTU1A3P6isUKPMQEz1W9+YozR6FwjNXl+wEzEJ
Wr/kqEltcfx097wtvf/qW7iiICRSI3D3uz1zlOuhYkSff4qhI8ITHnMraQFf
n0miXU5fJDokt6enGPS71DDW42gxuOHsvoiRA7LbIhZI013n6DUK5rivzlkn
7F74x2KegvFdjxwK+uOVu4tPlNZDNSXcRZj7r5uHvY0EeaihdrsHmU/jLnmo
nvWCbx8lQwwPJVzCzBZOhvFb8tkSEeZ9yy4vFGq3IEJrXS4nBBZUIF8Khxe0
Ebp/xKdUXkIMejTyjoa8qMlVzKHJ3zZBz4KfqlIi09OSq5Zey8MvHsoDLz5E
w+FVQ3czmF09k0Zt0fyLTd0cFmW7KEfD/xP148Hl6UmkrTOdK4Y+1lJ9kAR0
MObn7U2TlDu9xCqfiWYLQ3gyuCHuo/NcC2S9SdwuCn4lBWwEP4JzMo8vumD8
bcqXFuPKLOneqiJfR9ta1mHlLTjRv+dbwuw6ryrXh7yOTJZCaoeF3Z6uZH8I
6TN4NBNoOi2q2bbMYj7lJML1pE54ACfPh9UosOy2hnTHHFLsE4vOUHcMJUKC
DpJPsTWd3ftV6sBTIK+sAtSSS7AtDm5o+dM+6CLALQeLxsNUB2yo+9CVrY5w
3wj8Hj6rgTdf2vL8Qff6/7k6uieqwVzy2BpcoBWQaoIEPvPDiCs+0Uf6MbUu
H3mHwYG2MpuGOv+6GvQ27cD4Vh19Iflj5zN2oZnpeh8O4vaKQoolnjqss9rk
BFR/lyqYuATAskyotIEGS8vXR6xgxaFzQWpC+P2P2tfVoRRA/qso61riHBXe
b2xmbKFmA18RtpHqD0ykzbXV72h8MOj7z8nZE1sy0LhGHH+e88sEBvbqzNhQ
pOJcf4l0AT5lUQ2ZodBAeEpVsvv9mfCiMpMONZmQQaKpion7hR6o//e3Gf+Y
XMzIpecbGdVuMO0w+ptlkgYsswf6rorWUCOUBurh8bLfYL4Y7z1bogmIesEx
fmf20+iE/7KhnQBmPwIB5n4oO1whcgq/Vw+AUOg+NOkm46Dnv6DYK5ovdiqU
KwBOi92InS56R38cNZ/xDTvWKcK/IYDpvxfF2wRXVpOeg71Aoy5QI+DACZOn
0DtpfsyGqLXcCuOI02k0j+24BULOlBg5rcVAixbkdio+MzzJnx2QZjYMJDa7
cLowDgq/TP0KScSvrwDryh8DvUBiSNkbJUAugOE6xeFBut3xFXzviwI9Hid4
sB4j8fDMplBOh667YvJR3yYksV1kJtVxTgKbQ0AN8Ihn6iiuipVpR/ibFFRF
CCgM5+jGqDcpf9L2PGZU3OXWdgEwf7FBvHPUPGNaPVUhezZH9eWnEoaS1aEX
XK6I+YuCIItyySAKPUldxdJbJ5RnMC6nNwWibazhEdWB5jykQH2uV1PLysF3
ALlDzADvZPKuDwMQJZ+SnZfXiZnXi6Jkn8ApiJkGL5RIpNp8PHTHoktpSVNv
8lZhq2ozQomB1nwOE2UYOAUKRnRkrpr31NruEoRmQlRzUbzNEfaBKWtE2oO5
UOSWPKvdHV4+TbEN7YhIJZgNc3kc9+E+NzoQZ/qF4Xvxk8JIctjCQRxjWMHM
mLb6URING+XxiKbpdt8CrArt7tBSca0XYQQ8JIT+RbJdsbPpY2zW1qNadaDq
kW5+ZX7tB5s9R4AAE4OdBFKs6dgfX8GTsq83F4vellg66QRqTvDf4vlbW7gZ
XyworJ/la+DNNBsqAS70ASD+DAz32lZcVCmL3ZXPoHl0nsDUr7UaiNI1FSiz
Ze0rsJqYfg+82aaMr23q04/WxSR00xZp5/E68Rl+9RCr7W9MDTlFSB6tpRvP
sKZsMi7onjEzKxM+CcqkhKhNsaRYAh8J64fs0sUF6pKT507GK1R07wvu98i4
Y3i10Ll7j7t3OE62umPRxCixO83lXHa5PVV37e+boRYJBUfAG+yAETyOTW/b
GQ1dOSZsnTv7TA5+5d0JeImvrLhHpST5Lo2g9yPQtMcUEjH/q0FDHCf9u5wu
l+s/Rax0m31Ka+ORaxKB1+sKa1RIZDSGYltrXdXg/KHvVT3gR/t6QecBVbnN
91SxDO61p2Vd3R/D2eRwlpYpONIc8bP0BqeJjLKmLlMQXH1/rMRphUHqAT6q
p01Du6IrTsq6SXGPQqvPh0lPrw1UIN35uJ0lEUZpmixTs7IEXuzpqg95qAa7
2Xim4dWvSFeFatdsjMJhTCLZRZFTHkXjFCD3R9LZ/JT1QGkE3Ww2ahDCemlk
aGF/W4QWormsKqv2MIdIoobEdsoxEAvK+XO5TeSXUUXTrwapXaCmbfST7oPu
Oshp/cqlHnYv9YJ23xcDaDi+43X7I152BNfgFHs9JgWzP4Zb1jwSlF4r0bxr
n3zZbXPVf1ZYKJA94hWdvEj6ujKkCb4mv5Z0+7/rg40lA38aH9RelZhKj7a6
8IPGl6aNyUam3ouoVshPc0Vc19uOfOwGS2vHEjgC1Wjmabr+rR/uC9fxHKRv
KGtY/RGBFWLJjWzH3HX+NkV12PhDLaL7BHGnMOc1AB7XZmg4P1v4PwkCBWC1
6Wcq74PZZyzoCg7dQWTD8Qpdao2VfMUMESbfm+FcDWg+BiEb+aph5mh720+Q
DcqaFQ28oLObukxF8qNCyImKySXyz1yIL1Ksb3o2WYvG3sktxlBOuYFItOeI
L3XHVUL7uAGHYh5uamWtDcy0d9owejTeNwforzpZ6Cwrfb6Xyk6UF8DVN4ZF
WKXsytXypv6P5eE4MlceweS1oISJQLzZgzYIgm9kuQyAYo85YAsi4DO/Ekbw
IRyNWaaOqdaEAyzaZcsklvRWchkOCPjN9JgdtXtWpu96DbuNXlF4R5Ye91kL
DadUgPl+XEiYwL1WiqTNqREoLtxAarVqM9eOq9wVdcpTi2IplXEj0yhN4BCf
wDBKpIJS8O964YY+Mxf9tlZkMyEMozVSAUQ8+XK5AQ862QklNCcTseJaPfrA
UbyWMBiIUSginnmSq3gML+HcAxQdehcxUeWMAR8sDbPztun56Tt/R9N4JfJ7
jQ1r71uP2KvDOZs=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EyygBvFLLv6gYpLW5iPXFhg+q134eBWYGmGVxFPIafvBSKWjIdb4soAajJs3QfUrDSgMJuuF1aRe7tAi0sWy4aFlG6XCkxrERSkVCMCC1REowLVYXDxfNle62Wvm7FE1Olen25QYPP4PYucn7Rgq9EhUW7JZQd4rttGj3yjero+rrlO8zQxY8+mx9Jz10170RN3dLdbk+4qqM1EhySPlxYkCOb0npgvNk3bac+bxn4eURdcUQimFN8e3e2B0N4gTWdD1bOOL2k70vs1a7zI32QDZZSdf4FU6LvXZ/t5iaKRdobWEOPBGcbTlb6WNTcLurP57SSLBtIRfXF1ai4rl6Nw2VogtapcI+ZTVvVTMEudLTWk93+jTlN750HaLez2+ziXgPAIN3nsAPI4CXiwl77yTaj4o1nU0plVZj4q5vG9ZUhc56cK+oI2T8sLZMcPYAgupjo67qi8F12Ix2DZ7RS8qSBvER7cawatlcLdRb7wkfjAp0+ClqzUwRhYtE1YGmSCx6YwaCeX1LZ6uxCGk9uZbqt8QEeJBNJBpmDYLOX7854UsfTszGh0RjeOjwypvrS2xVVadf2v/Hr8tQu6vL4kyIyI9v6Y+xaRF6rD1ylHZEZtViqwSPEBMogCG7uAkm35/oe92rPbGRqcwTBPQpDe/1+UniB2j0J55sJgiZNUElVjOBaOhIe64YpDYfqSp0yvhuQsP1bMQfBzKtRTzQjqEiMy/tXuaKYbo2Y0l2spMIGD+LxZgcuikcxBLu6Y2h7F0thrW+uEXOIk0AYWFE2t"
`endif