// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
io4rAdnM/P0I6w+4YCTh999FmE1OxjRon+FWMDjtemGIm8Vj0PwH49T3qrnO
7MvLV5ec72hpBon71hR9fPaM55XUxoYYkx6vJeJ7SvPqmx94iP17Hxgb8qZ8
rEH3iJIrNNfy0djzDX5RMRrhvLUBXrm7bOGESanM0B9P1RklPRtfUG6p+woX
zoxRmd/r7FI4krwlqFnu9Wh+lydEFUPuMZ4RvqCEoR6425qwArgUQEBYwsd9
kbYcs173b8U8f+uH8L8oW0BzuEPj7v6DSyhG6z534fzXMlpBKm5ornGI8crC
YiqCEpjwSZg9b/tMi0ogj3s+zOJcKmaKKxLE3VHnQQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nMqfnreEHsJdxmrx/u7Tp7FiH1n3ZWKsRHrK2Hlyhx3mt/ZDjwLg0z0tryH3
9gN5wb5jCNPIA3BFOlQnyudO1odeQSzS24AT19PYEjgUQg5TuLKaxj9QOZ6L
d+5Sgys0wKM6iQrc8WPlf1yC2akyHAl/bNqmzV+5VFoXlEUuUFvqoIuswmlb
7/nFllvs1awaEi9NQhZtoMOi3RWLJG016ux5VVr5aDPO3GP3GB5V5H15CKLQ
BuhP++T7le5D+LyZ1tqGtmZhMNuBzGS14VvL1UJxQHIivNzdWfdl+4FZI42R
rJoNM9a+zd2BpSKaGMqlmjvFfO4e8z1cOYhuR1M77w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hBwkPo5Tvk3tifiT7HhbBbYk82ohwTgBpSUifJM9RBdFyHBpVDcOdn2AERl6
oN9hJ3YNu3+uGI2thv/Lw6TeKoDwgWgrIguPb19TL2rGEREpJMZxtRWHK4eF
5TvfNz2j2gvgoYh3so8dpT2gKm8gvqrk2AxBom4B8mYFg0MtovHaTgATcXU7
5PqvqhnW6tCn8CdCDhAGh0ST/NpXsdpWpjdH9mNa1XqIfDXjXw3QYAIyBMuR
2Sq5hUtb0vBjzykJxJw+f4m0b2JM+eoTzhPQMnvMc5/5+q3jZhuty7+RNmjV
nb2lxELDRDFyNpYtu+Ui5q7A5WHEMJRmFoYQZ2OxTA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S6lw/WMfrrTeY3mQEMZLc2V3Wh12ztbVCEn7XrHH12Bhru4AOxUXTpD0e4Ac
CsMoVVtVUKfwW/bAuOke45pxfoVhGR2IS1tj4dkOZ3pTX7GSBOlQtFuNhc9c
zpyaVFB5t4mi9bwXjEOoFn9LDlMwO94lXMHf2rIy96JTsPWi+AXZei3kUN+P
1kJq6OP4GMIZ8NW7Rcsp2IvXJPHAfECZcnNeRA2KBW4002ls6umanA2H4KE9
8HFMo9E2Q5omrkuF3lu8h1jAosaead7viNv0drPOuepPtWLvpUpTQWkTbzkk
9XEWjpgsMtxtkNY78d3ryJbO5i9Kzsk4NquduXArVw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aZ4kZaH9Y4xEMkCH9yUi16uyXlUJLBqMdiJAIX0lQSkfP77Y1UqHJg3UI/5a
aozvOUG9VBRdxQB9nRd5lARNL3jaHpmZQNsR/vgCL6ddh3HNoMWGPiDClTCW
y7A6/twySHBWNaoC1PLOuau57O7onYIUTVfmUta/JGuUEAFk/hw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ljfsfrc8bfKLgFd1rIMYQH0djESyvPO59jkWWDw08pJhHeHDsv2YyBLU+LQS
6JoNbWXgf+3Chi7zeacbPQTjLRw3z+RyPLiYB6T98WmveLJTNLaQQdeCVZno
UeC1TmNUVNA0tBFEStreYgLNJSv4pBvvShLfgRvzVOzLQq1UCrdMksZzAJUB
p1MAIEhqpw4gT0Oze9h7C64pLNfvw1IrsDW1oq267SrBtwDt+pzKKIvQu8BQ
if7q7NRP8oFZ0V/G+SDBtkwTcX9GZhr2umKNBwa9omScId/JxM3w4RavPADl
aa1YmjarnVUkdF3LLuTVizxgPIvoZmAUE0WoZWe0pY3WYwFvDqLF8uvKlfrE
SF2WktuDI4LTnb3Wx87Jozsy9p9rgphMl2eMELCUSAMrio48iKOSYyxBR/nJ
po2ThHkxiyZGJsN38ih4RRICdmPeOs3Y3ypF8Vbuk6F/6KqYSIHz//GmVgzU
iBernSZpRnGiAyO0yS093RxJvHaxUqOc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RNVjCBoTO3hZUtqKHg8y0DnyugugPH3RELwZ3YeD+M9Jji6HqPUs5UP/vtNs
UU/NeEcek10SK6hKyGT7mljrvN2LnmDOrFs117LSEDg4P5LYTjHdZsdXs/Xr
0gkDSWfoHsRCB2NwRdS0DAS1DUw9kzCRNRE2zz9uHM1D7tD9GTk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B6u6tB+AnwjAMCm2jZV1A3jVi8n861xHG0LAZ1pxU3x7RwfBA+l9vH9hGFAr
lJsOceoo5xwiVeguuvTh517pUZ9NTiNxxSBSkVQgpMX+m0wmvCTqI72HxWTo
fHGJQVXsIDKZ7zlosoR3nhQ7O9aqWYBxzf6LBIctyWm25OxYl54=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21856)
`pragma protect data_block
wmbiimS7/bs+5fOcdwVjofhR7Ha8+zu8bo41vy/FTuXX+VF0UuBkj8ZqzLT3
ptRjoiRBBEVDsk+aq9c8VcNOXHs7f7fW9lE9H02AHibgTGPqAnyrgbtVABkG
RInZwI3pFo7mVEFMluPaQqsPKj/Wz1NpxkQaSMp6rrZKJTc0mnvjiNlNPTKF
6NsUW7m721XaYTMfzW9kbkPp8lWnbCmwjzBUFaxeaDWr0mNfvfGXZ7NBDJfX
/MRwqHfeUWugnS+QDnWn7sR9FTJAOidweqq7CzkzHwYkQh+0id2i9VrqVTj/
oQ6snaiglEoteGY+JSV7k5/zPjhy2UIx7AjOc8F0acYq25oB2+Xih/Nu6gCa
QYowcTrGkSFPuctfadXRr63P0pyrBBAOZZ7s1FRYmzpzZxjT+32YfMXNOy4p
yO3UAiAjbwefCLMyj/IfkXIV6MCfLcfXqcrX/Z11+9svC3uv89ohx7kJ/d+t
yDKPh0LSquIXxTWpc4pNrYRM+YkI3GoTLe+SeDdNygs5ZUkQEKsMNk2aY+Us
ODRoJXj+5i3Xt8B8CCBRfQB0wv2+kD9n1wdkwtrKKrhvTM53cR4fBwBnt0Xk
wY/MJJOP1aCUQ0/oZVECfDhFRaf7P67o8AeZLonZ6RA46i3qGs2WVaotdGOq
8TE7leDjSRH/lDR1+r8s9nOCc7ElCQVA/ibDRRICpOwcenoX3fMkcQs9eZMA
8FGhiwDXMLPl7Pd/0/jRWq36ffJ+72KM0if/GuejOj4u+JSuy7mIqP2hcVyW
3C2SnzJqxYuzXoUIIYKCoOrOXbCc1yv8WiTZx7tzMS/f4Eu1+phToi67bXl0
midrHrl12NIv5KXNKH0CoEy7+lQP+9ssE1xXoqiBd0z41GmH/VKrN7WNCh4/
msN4ow/G77X43uFzNWufbxRbVoYUXDSRYMXWPSSFyqoVjDiGXgOcl2cWYMea
AsmPwN3ULf9380AWB1dst68u8mPUzX4iWGKu20Z9GiREllkOmxtTdW/YjvZq
ihBc4IjbLAa3ShPCz42yzPfsE1ffKa8fy3+NHuCIFAked2kIWJD7gVZ36RLt
KZxkZbm7wqVTpJtZqBqzWgXuHQ0oXeudj2b/PbxmQTRTEjO8490Ldn4AFU0d
P95T7Aayd7rvOjpohcrnt8uvCA32p/rqLzrYLo5lLvqCxxGXzLnzqW+tZRHa
ifdQF6CP1fbvqoCu9bBkt6OgzvONTwEHmQ3SLm1zKm45OOhil9k+SwVgv3JL
DUiHro3qoHkKU9JJKDIOmNexaD9T0PuFOEqkdmfXoly9AlKomQe4I5Bb3GJw
jVpabB2KYcdPniRzS5uz2DCL/v7tUVWCzvlEut/0xU2RzstarnhKvQo2/7Kd
r1ifD9WfU7FK52oF3QK3Kvo8kbVZxUzduERvv9RFpZ2JuMz+aoFK05upfyfi
u+JsCHYyNWTeUwiK9KnyXvDI5G0QB4Ai/QjmTKfksGnacHgfkxDF1PxcyAcg
Dli/6bNMj2IBfG9e1nuSQNMCYAfR53FoouApLiCLUn0Nos7QnQ9/wc3/isK/
1h84mXN/5EYVOSrDuRSm3hUYOdS81sWAgo7lM/TS3Rvv9IOcXHMH1qOayaV3
WPS3X/Zv73++itqzBLenS2Yrs0f4A95Q9vijfRoA+4Z9nbff2DD++tzYt8RI
Ds7pRTUjFOXSJFloXalTFNulQdUcDhWoHaljuubpfzkcAv7LRZog/GKmuFmt
2TLo37t8F1SlNX2nVGTSALCyXqR+m4aIuWoxGIaEUZzi5VsrYJmn32q1OngA
+vmnWeR+BRni21n9sdoGftk7pr/xChEaXRD3rT7XjwwJHfcLregH1zYtkgj0
YoLWljCtg9MLdOt+EMdHqMx2hwvfQGhaDo8YrjTFbnRH7waxdUM5clUcxfn+
SWfwkJrmPXBqgGCK4IZPPNNKrwVimuXs0xd708zDIkQyIrG/OzANxM5ncd1s
p3MBuzaohKm9+gU4gJ/py9LYvg+vTQ4MfacFcsNisAyuabJXZFEzmMsPvUf6
Gh/DqV+pt+0++L+t0906Ia4aC9oukvLazCIcXFAT1fSYUJngrpANtj8yZzZU
U5APjGnL0Pf08P+vNSTk9rHuLq+aPrUTRV74odxxgWln6I9a9nJLkbSpGvsN
eQWxB+EG9BjRmGp2jOxyi5cjg0gHqb7xV2EhBC6n2nBrMKFpJY1x/uzee281
FBX6154EeBpazVHARrRGp23HdkSgKOrftOjgIP0KXwXfsY2db5fl3JBpYERU
Ois3ROj6zItlFIHkhIroPEyXrpUMUrhP/aCnm1ZdFPg5vff4EKhw1subu7Po
WuYNsWg5UDtFGA0P2h4bxBLMbJ+GuJr1532Z8N+gIiZh5kHoeso2sWT7VJoE
8aW/qe+Hhs6PT0rPfuA/6d111Mo8XwSuU7Lr3sKzDsiswoWIvpvenK8EkEp+
gzpzFBVMA5D8XQcGsO4Cq2aXzNfGjdSmmYGThRwi6ALVfLRmkZCzjcicOoM5
pt7LKqpB18FUEVxB/QzcaSyZ9jZiTQB03aeL6qksNilzjjnnnMYvt12UJQ4O
1mJIPFeY73VuChpDxOcLIyU41i1d0ZxkBbpNjX/MP7cvk6R3MN1VM8vGkJnH
LF3Hb7ExZHcGj7VqxfCOdam52VW2tuo4DQiRDahf2wa+388/+k+i2QZ0xyxK
8pMBB0pm0Jy5XNVhPeA+BHsAS8D/CN6taNjJgMW+Ymhb+MBqKfqjicclrRzt
hRAf1UTOD3mk0fWgUNIWj1YxanXtHFOs5H/eDKNgIZ+GIEMb8UC4np+Qy9v5
jInTe6j9zk1C+CSU5GXxflUjhksqsuoViTgZlGeCvqI6LC/OQURq+JXWSptM
t0P3zp+rHwdMI/1xDCLB1agk/KKm/H+spQRYUzuiwj5r4y0bC5dIL+eXRmHi
SPgGWrsitLpQh6rwUI/cuG1Sr+qR6r2WjkIL1GKlZGyFmo0/5/ZVVnJSTTgC
0ahjWxARLtv3Va+2SH3/FVi5MhMKc/8YBeY5Jxz5KKxwkFGOpvmj8Eoax4/j
Kkt/hDeIipCbyEvPlxe4zjz8uTStSefiZiAJMaYBFkAH3ltQU8jEKu5xPeYZ
Qsk0IgDSIM7ij5rUaG2dp8xHdkhxg9a+NWuCSWsdMMeucrdFMuXXYrhD2S1K
ng0BM+HIlbQx+AkYEBQBnpcXiaUWs2Mq7GUoI4vziYPx8TxiB5OlYorXXER7
UitZP8Nc26NcVp5xY2uG4GNR2+IccLcYqb29jXYYHFNznVXLU+HKAYgOQUT3
UjHNa+4lC0j+hORq7sk+KFTlt1gkhXdYUbg/SR001RIBNjB7zDQyPxiSd9BZ
fpitqaYf3/K3OvyeUsYQHFfcr1+Js+3dvRCsS1cNzEEowcDxPeoTCT1jDd0V
Xhk4yEKhdiXGactAxb0jg3/4Fjif1Omez8F7dAI+m/00mbcKkz4OxQcdJNLC
ssWDISQU52581B+wByqLOFN70uGuO0iTr44+dDOYw67Tdw6Xk7JeA1WVCc7A
+qaM9h3Qufi/QDBI/ZQT49oPuHvyuoUzIMZ+5AunkpHk3FkbiZIHygYS0Xqe
3sxIswjSrmpcmTQrPOs5oOuKg3It9COh93g/2IfrI1UW3fBCoQpJw26VSDsn
jotP5Of/E9ceGOZfomhfbL18Kt9M5pcDhl7hZxPAUz3GHrksvDtOIgduxCb1
1z4PJ589Jd/7/XtEX+X2+qWC2hzEKBfyk7jwsoGCpm+5NH9r2ecBizguqYdG
ADYYUZq9OCrS1f6+E3tg8jWNFRjKBcLPiW/LPKDaCqn29Jptxj64ixUUmsH6
3JS1o4sTrYI+pJHkr4x891djRWivTjgUYhDwRi5iLpaEtUE0JrwKwC9vOfbJ
Tv0xWx5LMdEWaoMlnghVpBvJv/896tjrqwFwPay/Jx+BxyreCnzkUzETNfcU
CTWAUCb2l36yuB05DpR8oi9egm3Id2ZIEy/ZxKr5nWZbpBvW7IZkAwaTA+nr
XppdFFlmJS10ql9KczyJ01d6dGvwgTsxyyyFNoZvwIG3q6zrLAcF0DRKXtkx
XZmp9+KevpD9vB5difjARoAaamYhqoINCzavvVNJSr9ZTJQG4hZauERPHzKa
qLhkulDEIv1s8BbkftA4q49o3EoQ2/9cPTNhrxuhrvlm5xZWO3HRdqYNkh+p
myxMmdyrvJTnn9IGhKk9rC0nmOP04SUoYJ9IVr9dFuW24He4O3AtMQtLXoJj
3YpH8auoCsjQru71b6iYXCAVnGrYyBzo16ukqEuxQtv/Zx8c6ql0mnQgQ2gm
85Y00iAUrqVIS4X9vIuRxCa/4Fg6q6vCzpHB4CUxWhCu6eeZmej1FgzXHHc3
sit0FBSVNdcVd82th7PokObMd/7rzd49oegbL+3Hc3/de/MFjinvXT6OS0hr
skeqLZ44J0snCkiXgdzRul/o+wyHjeyTJc7pFNa3t4skiWpjJ+2NnZjsiJn8
j5nLnj4oLxECMqxmODmQFpD0Ws8BpHOO7Y68YwBvymisCZwhVjFspCzhsF5d
zGT/tyjlf8+7gjKTrZFubhBSikQvbGuHV8Srbyrm0g4B+qzEHF9lcga+BKo/
EAWaEm4PBbo2AISCnHHTxYNDOtESgeoj8vJr99WZDgsbuSSOJV5pgbVuaYbt
KSBQnFV31N5xChMVejW2X4sSiFsag5pH8ijvINSoJdkADfLR98TxpAYR44Xv
lc+emAvl04e3wDAJFTsT+QQpin8evP/RumAeA/7tBj2bwktyQ3Fj0/ixFZM6
S/xaTat49dJaakJrUHTgYSKFvHbVhoUUS+adpJsmmTYrAScNBNckYYGWn3QE
1lYCAWt9We9SEkji2ao/hmV1aucI7IudUwNuttv+FgqVYvcm0Vv0iYlWHEDl
08ov0DmZKnYPN+GDPz+vAsIfpyjbzTrXE8kxbEgW3hlYi94AlcV1p1X4dQ7N
q+ZV87xEcIuitvYg4f9DMfJkfJiedllmBflbZH3X6w1kdQZjEsq/3S4EFU3Y
JGEM+GkTpWGO9YBmcrLhKYI9SDkVT2s47s2vwvgiUA9iog6m7MfGqaI+j4eV
XcmKcgY9uWE+EkblsdT3o/dCM7lsrUEwoS6DcJH1RJgXI4nENhviIZM7j12p
+9FKE2xU/NWxlOBiF4EMSD3wrXbkiSXoCL6wj9ImIWuBF7xk0nPJQJuvYCrk
mGXIMxDQ5CTz4kJwA12HJPHFSRypFihF2X8zf7EFjJ3iIcrSOZAb81ll6yw8
W6oOy/WQjVHNpximSfZX3K08hAhfv6UBMkeEOo+QAGtGaSj/iAMKQkxLaaX6
bR89zNiatvLFFuPxl6icgT7qN8wy5Ja23JlIqoIFvIKeU+9Ob2nWK2WUCAqX
uaKVo9O2E8VDY5tFcrgLKp5vApB3fs2rGDIRTD5MPXmapIQ4qrZlqyB1PH45
NnbcVHiaiDJ3OXr2m94oqzJ8TP/q8AF+TzN4y8xtpviiVz7Zx5H/rFZTyp+s
GCSW3e98m+v70s8e+3z9fBSJFqu6Ki14oFHb1JgV3xMYK0gsPTxm2AfTFowN
mtSPLFpIFWRRQs8SJl+f/hN0LUnekZvLh3dlHjX8YrFFKJXXuvaPPAXW5S+o
00akJCdoKG4g8z1FZrkHo6NI8U4P8DkQgLp2Bq6SmSbHmnwrlkIikRumOHe0
rwysRBDD1Fpbz08BGEbZJVHHaZQr5YTb/nC0AJERPT4u4lZvuORijHTQCrCO
0f1UoeG37pjYBeS/nuq7XDWRtVLbqGDT+HdUcjGVlyM5i7LC8iwHGy2lOAHu
zAl1PPTLVFbkKcwHQ4PvSHypFTiyZRBl+uqgy4Ra4ZmUcXAotU/0WFbyfKcN
GoedQ/WtOrmeT/hUG2Dug4hzFEFPp06fZqZI6TdCbPWHtSmIYLFebQ7bQBum
UCuWLsygYYmRZ+UVXaRsPFVSb+l1cE/KJ/kSz7mdwW69GnvsYjZ3kZEd/hxN
qRrS+QZBq5sRvctUJTt+sozZr7o55790C4UFbXBGWUW2Iw/PNWjGJafPG5yc
fGW1BGcGNJdL6xIE09xKAbm3+fAAHHzla1OvZlu7eJGpHfdVm076bv/8YwWO
T1MX2NbzOtKDPxMfzdvMrNTvR1hIL1OcAej6yTwazz64mf1wz0Vxwwu9ydrB
8kj096FERUfgwXYAHO3+4FtgD/CvopqWbz19w3iEKn6SJ5KPo5YiOnt2JB49
rzt1RBJMAzC3ecAPkYc2ND8Jo87tHS9KOPKcdRsnsrmOwOwl6kLmGHVNAk5p
tT12HZS9uLvPubYDJhu6SE42qsSzDrECLCbsvzqlje20OTXjF48v0PUReP/O
Fe/BYeE0hnvxbjP/tsmDc2Yl1gFzIFrVjJBrPApnRaB4yYfh/2uCreL76mDZ
Lx56k29owrMswaUKButh4LKsUvFRKpFUXB0js2o9N39v3OuqE03j4m+JXk5y
K8G6kssE50aj3P8BmE49Qh2HC4RS8WovbbpNf0m14x3VRVxmZjc4qBgmoSAX
YTkzZriOKy5dpagKDHTmwzzSwycxTI33b7EPYY98WNjHYZE2P2NN67dZvLMJ
DjRiaKdLMmlIQ/QjbtRnypIM9CEgIII47ofMPu4hjQo5hZKnxKNH4dCKAeEy
qCurmsaJCl+jVesehauDJMMsuoPi0g3CFKZ9+fGdx/5suyOO616STDBq0eU6
6GKekaX/k0nbU31hO/x9AxpnytkmwbNXEPjtgfzl8XHE9vgro83o9MDqLECE
OEo/MiQ+4euuvsNROiJyBJ7flQvvCAZVqqq1icXDrXTufEf+KpO656sii3UC
kD/sHkRF4bAlNNM3agRQRsI4ke+7rjDkM1QhLYB+bW5Ax3z/uyt62u+Xwy92
hjxGL+H2QXph9+oaZi9ZhSUiytoeK2t0G/KsBJEYGu7PtG6j4Dx5w8u4hZNX
O+gEaq9hBAkQ9/eszaVf7YmI2kpQSKwnbCsLoBvUfQrUDJhGJlcuA07KWUEf
ltSF3V5Lzk9YyO88np4PUaj8ZFg45mYu88Uz7PGCVsR6U2jYkxOyCCEtosy/
67rbKYAiKd72vukC20IxCK2VQSBAawSATRPzXJHMR6RuOORS/VBCCZ6udn7L
1K77JNvmlvtIJfrpCi4rSgaBia7aVXTXQyWgx3MHVk47BzvXMjo+P8oW4m1v
DfxSUXajT6YZ1hCO98Rlm8zkZOJQQ4AJDCinB8VTLkfnWcQQWICaVsYGw3gI
ADQ4JU3c5w+b5TXP2EhK59VkX5KFT5Q/rU4AZo4TnYKddw79l/d57KQsluX1
4LGU+ivnW2wZHJhz4n6hwMmHIPn2He5J6B/yq8NJQeZ4E7rQgNBGUJTHvLzq
22PBLnKR2wCzAQNNLzPkixd150/yjvq5G1+6Ot+IXr/rvDfoyw1qkfve29Ey
09y4zOJtepu4KrUlLNKMGYUIUTjy9QQY/7LSHJcMSZsGZUAzfFk6aq4KwcFP
jjyPqRw6v1kPV/3/FNdTefTMt/bCuOzSsPGvtY9f+BnxMv06V3ve9tfQWt0t
wg+tjuC/hQycR+vEIDDhl9e9Nm70if+nBGjpP/ipM5h08QuBHtjmi/BbWswC
swe2H8PL6XN/QmRR/ddCdTovXxPw/O/uG1Sr75tb+q2t87UoFXNKNI8DVMbX
djy57WEUv4KeYsYZOlkS7/6TuMeBb8QBQsDDvvVew/1P9W8ii5mSQ12t3M7K
7UmS6D7Fy7enRJOYPAe6rUgyT8zMBZQvr9Lx9YWVPO6+AyfZK0fI2s/QQu2E
VbWlYXC+WUDKn6KHlni+fUkXqhv5rgs4ncBcjdXQ2/O3N210IlBFHI+HwgPi
TxmRhIGTK2Iiyw5MW8zAOUraUWbkTJ+4aR0RddpyuTbAaqLSzMKUVpZIwchp
shsGXwUSBi69+bi8Aydui6xA/0yVHg5u3YJ3fbDDZiuNzXHuA+fUugCVO9qq
jjnGEVzpwhDaLTjFqCjAY/80CQCUTABgjw8C1F6CZO336GgQ775m7qk+wBs3
myLM9GlJx37LmdBPqz0v3bdWSqzrjkrj/BfDTanpLgg1Dl1kdrJvdltGZ8Ej
/GtRAkUCPyuWt58tnFTx2/zD6ZubWxyUZ0s9K03UW2fZaB1SoaQ6XiOfYT/G
ZHAPgYwC8hhLpBmleun1ple95Ok1VZlO+JZFFcYUrqamwRrStkmbKecyh6Ke
+WQ9ekK4l+u3WrLNND0fsfjKp+DUdZdVGYf/eHANA1VG2QVM4EnKv51jiKto
0n6r9XAguNxi8bFUT6K1tjBnY+u79/3jIwcSL2Thb/5S9SlglIv9BBHXtswQ
1fBe1704l8SK/oo/GfufYrLJ/NuEK+wEikN3oNn7mOBeCph6bS5FX04K+mSt
XamuJSPFFp6hy3rbf78mIqLOVbzPvkzHm4p6q4EzIaEeCdwPYcare45hxjeP
HUZfNrZadpDrykHoV7nQWTfDC7UPHXig4u77FSJgQie4ZciK73OdjCyNh3w1
QjpuzhhVjOcwA3h+KZG5g2gR/nEPswA4M03mJYYVsX42+O1Bm+8h/OijInAF
P1gY54XGiwXSar83ylcVIhPlIYpV7BOgshWHKXQxwWUg2lzyfTaPMOKWZtvj
KePqslyxe92NI6abQMksJGCKQqqkXf1sJ2vHfdEXxoBkyoAjuVJZhqt1ZD6H
BUM3hPHTpGVAENChw0He3UCMP+B44jeAtEXAdiLGL/ienQhsjhEOVelZ6lP/
arpVPWXu1DB3kdPEJv6kj+d/QY02hTtXQcyhwhbez3UyXg2fZrvZCvlyoWAD
uWTdvHbv956sxXThCU+hksO8085Flls2+YbD2Iya4ZraXKCx812vP3njbHvM
rlZVdn0ZA78LW1ZaeMj8rY0anOGshp4H/1TzpYEUixwp0I8Zqm+MVx2ofD0l
f75H/Oy/C+zzAg49ZzbXAfVRuOh/LhdwsmR/FKFuMdudSfi9lpaSDDI6cxsD
mlI/5G6rnNNUiaHqSaPAtlff3OxTChHhialHa4sbGHzkLSm2OLZNhyjh3I/t
NOLpezMYjDHto1hNw3nmpdc2w0Q3IqbpKvfzuP2B/+jLIR/C2qi+ceGA8J7X
zbp479dAa7aEhYCcgkOdOnXqVa2bFajmykcgOKfKxJaYlDzgE1ct3TUs5cVX
dEi80F2m1mQ77AKwq+9NZe/M3P2+w0U2rU9Kaf7LlFYUA+lHarud1XNXhhpi
s9bwwanFFsQKkQoUMb0gaEIxulZsdg4nk6kQzSA4tb9iBMuZZ+nxiuTSgi0J
YlmAUDwsz6DWXhkqyRLtc6oxAanRjZlgOHqOzf8ySIXJ6OCbhrN8JBdnNvv+
yxKMkndRCgAmr7D+XOdTI/9uwoZH153//JnVSOpyyaOowDhWVPFrdBTI7I4+
vCrJcZYWR3bW76ce67pUKLyLNOYepQJL4YFzvbDZyC+VR4WmynrPxzqVRJYz
AP37VieVzT18kNMTJ1uMOMCqd46zhWFcUxKFF/XQ2C1Sj1Mvfre8inObLR9Q
nMP8H7Fdo2Z1vGRkoelmkfqgKzy6yzkb01mIxIUoJdTZt+8ZGInpiGX655JS
bRtk1rneCp/ccmkwzmoJVbLaIzXmjcTRdlWR1OKbKJfdo7m9QvoZn4KliIui
THv7PQ5qEjj4GivEdwB2bXI/T4AH/YQ4lM4isrdQ74KcEcPVF+sNf0i8yObv
5sEyNhB2dm7FEM/GTVakddqcFjRuB102ohJlAgZHOI01B94ptteETVmbd5cS
qBKwnmymwjrIvtvNwDU1IsaotHG/K9SsWTe+wgbBfWHv0JjfV38zYabDYpcn
Pd/eyMw/MTfHJ8z1lt7pcySXNNofmOETNoF0STYlSsS/A3netIMLm6XPLyE0
S2o9vkTYtRNVh0muQWQmGzEBp3bX3bUzRxre46Qo2emMEHtedL1f6V7Hr9zq
USaSCiHpANFc+kc/mhW8AfoAcHDs0/ZsPPld3tBqGc7RQyWdsiIk91E00AWf
93WbqP9Tgw1qtWPkxVezbjxY0MnylfprZLT5l5Uru4W6lzysqkWkXjwoIytG
3aiHnhTLMrdIubrGriD6XHKWW/2e/ofQYnDc7/5zzHYK/NWVbBmO+ALo+uxg
xHNF9u2s3Kx+imdWYM0STeOE7ntv8dqFudQG3Qh9JvqldXBHL1KcIMizAg8c
vQ87YXGVvBmt1BJ+gqQiXa91+oYoIFu/PM8UiFKDN9kjaOXzCX6GWMCRWzLP
+j29Ufndm1Q/7JfPECgh35ofoaGLHmv4s9F6YbWwUDWbxpqdrV22vW16e3Wj
tiLH4jeKT7+HDM8HWCsP30E7h/3cLkWPgzu5bUl2/8WX4I7e/efK9TAcaDDw
Z8zNm7GdSOR9cLFHQ9fDWXgBdsRsgHEj5++6vMbVCmPIi7n5CMHMk241LME4
2exX8NZ95tUOUh/T5VooNxFeg83yaGYWHVn5657dmUhxaBsj0u3TmQAF3Vf1
MUIHt42Z+8cRJ3sICB9R+Lxzuf1955E5nHmQZ+gnQFsWUgCG40TXR9UkFCrs
FSQtuQxw895f5Zk8uV7AkFexay7XSI/EwqgEs11H5RhD9qEdGMgpUN79lvBY
LSU/bHpZI6bW03Ky63hOSgW1WJ/W56afg5e3dLD9GmqXk1KmazkU23hA6uEL
nrROLMjHD1MT8gj/7Wg2i24gmasBEQB02FCjeoD6Ko3JlSHWE2cgGRfoj6EO
hhnjaK6OUXPEKd8b8H0zMheBegU98F7PU2l786Z1FctJcgv7D9W8Va9UMrl1
LZMSrkiQXgSeYTSJceYRMGJDMrvgMhSbaky3UIHqauvo4bRlAEquSfDonWbD
jHiRzIjFYARhMh1gMdqp8klHN9EKUe4y1nBNHtU+29sv3KdRgbUBz9wBFhHB
Kwv7PIGZ5jw/Y8XL1pYGHFVztjDOvcrhfZd9yZTzzfpbiOuT8N1ZaKBQ2Lj8
iXRSXvFCTsVW3BSLEiIAl04lVDtSaq/ETY6TZD6QBHRZTwCTR4WEKe+z61mC
myOcBranLL9Nbvhu5qVytDc/kcOXJM8qUnoPnT8nyV1q9JKSFq725JnkeX4e
o8h0qgM7Yk1mb7ww/fDPJJ00eFPLQnR0OLGrFbxyigk9LYI2mF0VO9T+WVl0
jDspqTSDueNWs3KbDN82HlG3nmSDy4qlCMia+2dT/Zb7C+ZeywPlhoLTZ6ap
4nrP9yXB2fTfy6NpgtC06b1yi7dpfufHdHL+chZOn+MBYPrMf7MY9Ti1qzgi
Mfm1QZc6mcH86OhsBjJ348cUMXH1q9GjfmPBHi5mrLmu3aKX/5q/LkIz1jbv
2RlHE8hSK2wfyT4t0UTsTmsn88Sj7SZ7PVl9mMwQXag4mXKHgeA6LQJ8SOTP
Tm9cpb7K2TvC7PdopwZ/oPVj9sjvU5Q+hTEY3j4zvdCd0DqZFs0r7Lq64teL
f23K0SeyobbyEbXQrgysjHK0JQULuUPZXSvK2nb7vy1C1gS1BbuWOWu/MYaM
3Dij96RFOYyO8KmkOzE0R0s/VmhwYk3sXgdXaqt2NATwJ0sS8ubcFe1X9Pso
oHmkgkiQ2Qw5/5XpuZmDERpwu39udTC53uIu1hvvPL+Y5HSzjj3XnVmPUt8E
Hph0kHE6qQgURjpDsnkrooKGJaDrYXnB4SZR0Cl++qVu9TITzth3TB/q+tr9
LF8oqKMaDulfUulqQlSJ+TklA5SZ97CCcJndAD6swG/3C9GrerGdHvL6Bbph
I6m6BHpVkmqQk7MtD966shaBSyQkhNw2lcYMAB/7TyiMcIYx4as5MtTIz/uP
AMpL2SsXPbXwVELcrjCUJGNs88x8fmf9g7q1wGOq1ZsFnduf2ilxpFx8hzkW
5duflZKPmzLhkfe7uA6Zl/73W8sTbEArW8O/hBFn12G0w2tzkVDnsgDDm1RS
Axrg2VF2wq9/+hhDRgyoaUlF3vYPhzUhD++fVbbQbxqwRNopqCyozP3cMOjC
mxNVGSGx3rDbNJ+TG1J/MyfEXy75OeMo9LSN2GOWVp7igraRb+iWoG3PoKZL
3RLzU4ctIxn6EXcsE5vZhPIZIsijpbAllCfgwCKUcHt3GcBvVqsGv/nDbV+I
8QLsXmyFZequPMuOuAPLFHARzc16WUaZkPR7cA0I9Q/ZjSyYnB3lyq/aJe8f
1IbLZlQK3CyT+Ktr+UXRf+yxz0mzTPjQszyC2nptOJx767kXAeUqZMXzdG9h
X75Xm0yiXY1eTIe1QfpoVgdtLEQp5k+mAKfUjg3AjHFJpT1xyMFLEn6Ea3GS
vCmUcoY/xIwPNfIl8xF1xSsnI1S4khB2viSZyMiiyUbMbTlYPLNWZF0pIPvh
EFnU3v2yz+EdlTgTu9SBnWctziwJoVvxG1FHowpdrg2L/7mwet2O8YgfEcec
KMdHhsmudlE3A7qv7LwslB7iEDNYxiXG+kZyjN2Xj8Vx3KapM7Maot6aMOIH
yZ7tr+4GK1Z1PYzF4S+Qrm3GslS1OAk6yMeUwFyVbXvZGY5m1LTZSgz1Ekz8
mategQ/RLoyDla/ZapdeZSpdTpJ5M/nU3bDWG1uIe/g/J5Uwqb7ZcY3gG97U
eIBEwtA3tLRfCd3svKzT4V4nXJkSqEs7CnHYefNe6YbGqDeY+N/TKtrae1Rb
qee/yrB6XDmwQjlwEZ+1K6XPU0JX1I6IsJTOZbqkU3ioT4j1US2agUvH24aI
Eb64F7pKNwKe1iQ0vsqHEDQ/6T+hIPaFS48SuaDMsPz3LIyM2FsTR3kmK+Zp
GcCrA0pFZpyVJ56FncRCJ8fbKbBuwBq+kVNXcoQ26TIep2FLY1C+hFHjIDEL
LKG7x01zELf5dYIHz+SNpw3xKwh868uiZG1gRxBEMmQceNdmcK650FKTA80i
nRoOxE/YQQhOh69Pl2WYZhoSPSLhz268GFDLJawB8PQCxJ5hH9sWxSOKiFPu
AVRpCjJhc4S4XSqAM/R8IgYPC0OCsNv8NBudTqmreDA18ijSwto+AE9Lm4SX
jWBRRm4AiPqYY+aWZRZcC5O2bx7KR47OLScoDOcjJk8bF74EIorX3WpYwdTb
dRSKANIY4u4dE6Kh/aK3kmIXgDMYbx2f7yxXgBqbFSU06Uczgmx7nBC7q9Du
Kwp/n0ULA/nzM0pdREF8hy+MOOg92TdsktT3Z1Ar1t5XViW0jd1IV059+6xM
sbAKrOdnz2Cs2zLCaExTGE9FsF3Zs51ZnHQ0NMEfle9NU9Uoh5KBZ7xzVeg2
MdqH0JXll2nBnLvSKsQetNXC2IpsswUl9NCqvtO13YwwhO1wuHFmgAsmGRI4
aL0w8G1+4IaO5BH6rWPnVNWaXmQ/+Xz45/Q32xFgAQUXnMlmFAnHeVWl3q15
RkufFXy1RQ463gNBOU3vSf+JFN2Y5bpzWo5SeQlGOq6JeTgyNvWJIl6aPdcy
EHJJACIXTraXDXOAgG4aNWM2P69jnG0B7/MDPPLJAjS61b00+qBjA/xmmM1J
lPJaSeBMsb/HuMiuCIsSoMIfFNwki6NbHroJn+8fkBnapsfWWoTflwsED2OC
1e5aBgjl3Z2fBCafMuXUgUmVBfX2upmbtl4voWjov5jtZZeOCvQEMKhAu32C
haJ+NK7LfDdv+Sw2nCQ6x9ieK0aYsu9iVaywjNLfTiG0H8DyIDqFXxjXkMb0
B1gf/S56FSdqIw9DUzjxBYI5eW+RG/0UQZbigSaLhYJgWpPEQFQ5CA5vrG7o
bkoQODdqBEhrEQgVet9+a+AwnLDVSuTfB+0oBiQi1CKNek3WrlmzYDXdyTWN
Flb4aPoFSDoDBAaZG0TMi8uiYJqOm6NKiq2GF9VrdTo8zMVh7azrAhk+5Ns0
RazQt9/w/g40mQM83PMMgPi1XnD+zFlyAZLqHkkXk6qJ8DkBjFfV2psADVm6
ukeyxsV1vt0Nqg7MGb8rECsB1Dg4/PDBSFDcufvWr14c1S1YtCffF51B1PfH
Rljce6uL+o12NSBg9FTbN/y00egGDo8TmLTvcEgcXHN5Pu+aImyCru0X90N0
rk602kVWj1lAb3CXP532BtXryOGsKkav8z9UwqeptzdpHb630sYuo42i2EsH
2hm3dXhjN2n2OtUP5FRG9/iH1hQw1H18qGfBWWPzLfS6QzkgYLGAIM4vfJ+9
jdwOOmBQiD9cOukcFT93eD5szT6eIommN/1UaIDmLmVx1tWGO6Nd7qxw7Goa
B3TWm0UOGqhgoJAKKxTbdqQTEOqMh9F444fRlrXKBa2od/ifhoQRWKdHQGya
fAM2BXDdFoS1wxdLW/78/T8f0CU1tJv6+7HWHaws1NO2iE8WSCT4Eek7AmrM
YKFC02IkvneON4pgqDfah2loqv0zteRZwQSkaJCQs57l/joVfOvbzQN3ODLc
frerhKV3JPadwl8xtxju/MmGkQPBWy/zkoFnTTDMsYuf3CMX7hRf0DAJ6rD7
ggpwe7TRezbTHoXXec8iJ80mmInuXAUMIdOCdrAUWpi/0NgJweeEjvWdEUhQ
9UCVl/L5FDjrWV/mcvQnZvKKVZfu12vVUV175a5Gv7f7SkAh/AOF3w4Ghznt
RVNENm89UwXdsDvbe7IGTC06EHHe4e9z0952QcmDCc7A/5NfmmK+DFY5EZOG
NtAdWMjn+iiQ6F1mI0IPZme2myDnKcsPD1+7/gWG4NKVl6ncoQ/k1pmIjh5+
PexSUGpLPWndN1DUI7RozfPUFIDDZJgwbyUKRqB5BUgur7QfKlkl7mtaeGe1
gdLm3poMw+7mGhibApjCtEYL0twt//kGa5cJysAP12gPku91lw18kWKSRNUF
JQ7ruk/hzE6WRyTcdwyuP6SIo0hryyp0VJlUWUFsZ9DgxTtq6Far12JgWXMB
BdWQoBlxuhy3InsaU6rw8BmrTpRxZ+LQlTN5Ta/HyE8rKNjB8jsaYw6sTdB0
WehOg+yMTyKv4NiTK0J8IrI2Rk+2RM9uA6T+lW+AZVkjrPSzImnZnMJqMpt4
OgZ9D2+BbuqW/4LRlL2vL9mteAG/N6eaHlJwJcBKMY5Vqr8+3UTF06LC4CW4
TMC9xMUSd3wPc6+YC5nkwvmSWDurv83gOS5OCF9Fn89VjUzveqwIJZYu3Mp6
JBuUsBmMXJdBBr+vkcxH5CwGSW0Gn3ouZKjfd0Bf35ez2dQbqC5akC1UACFd
XIit4d4tn2nE4HTe3tojt2lL3C1DuW2GvVJbsRFJYx1hq0UIpCdGMIEnmeHw
NPZAqZ2VisEDS/SsIobY8kQxFtaQ6Q7M8aocGt9MoJtNxeyoWrGSBfY1ED0Y
8ZbmD+f4r2rt4LlaCjjJ9lRZNYUeoKUSf70lP0TiEfeTQFSuDYev+uIeGBPs
Wd+V3XOQJiSkqdGA8koLrTahypX92ChQzj2xle1GhLFVqbJw5BLMgGLjK0km
+CpfK5EA3bpl5hxSoignp5QwVvQYGAnrO0L3XCm/pPyOh+l4GPc7ELliYpi6
2v+CCAVdGjeUakaeNzlicvhW+7a2S5f9EeNpGCwjs1pWM7tTiCFXUfyGEq3Y
iKOI1YihGnWvs9qyqS05l8fMX7sb9FhDepHRx7W9y0vcqtZfBNvdUFErmNWh
n8tB13cxsyyFy0Dq6nIPM0Ylbuv28Vp+lJo3ngfiBbAEf7eIKrx9GaP3i0Wp
DxsFe9yiWAGIZ6xCVbYRDmygFKUBRZfm1ix1YYS96n4bIUHZxCKzRScY0xI6
iXR+Y0EBeNyt/gNpqFsGkIA/6/T472xi0dWov3uIskKZDYFeNY/AG1x8/AQ1
Wv/6hrhOcpEew27Ziic0hIBALRqtUZlc1JRroTvQ+xtsO2D/wnJNqjWRrAwz
DxAdZIDNZDzp+Muf67/QCBpC24z+uW+wzeD1oZieo1oKDstsJjhHEsabK4KC
Xw1okx+dDmxDgcn7oyOU1vTlW5NOZ6CezRg5bnzQGYQysfEPBC/LKSUS0fgn
hStPfp2+bEImKaDrmMqk2JwLAdMcA9y+9sWir8G3HqrSMktAYjSFDSjEyri1
cwWNGBtdLRgcHOgYCUQsHw7v6MZsTpcwnEDXcNZ43y8PkVOlszap1aUvlu2a
cOfmLCOVAzQtQzw62507PZSqgbQi7Wjrot/xHrd4xHC0r2uf+vaNYDg2wMxn
l/lz8H3GWSG2ULnJCv4xo3wi/POEK7JHj/Af53B7ZEIMVZOrlHak4TYwhlRl
BvswwB1t2UNHzLURl6fofFUmtuD1gaNjEh5465HsKtPeA3PwFbst9NIYc0yJ
4pb0HQ72T/jbD2xXRsPoLB8UKhmTjFGnm1oMwRhP5xMsTb3wWyZSyl6RTw9r
JD/B2XCagqKCt8vRnWSZUg0zfDgmNLxHLQTA+vUFa9Ho2EJhIkhM8ReMNqdv
+pyTbcbHyFkAf1pR4oltOTRsp1ZSilHoZzTYf5s3ZwPk24a/bQVdq/CQ0iVy
VIKoXqHaWd2H5JZ7mjvJiJGRz1CjJQ9L6xStguFoHWD8yl9mohu7wJzWOJnk
8r90VO279H6AfhUJKzRMPimbt0o3LK6WTXM18Zi1eADqyWbeYTJK/zRgRGPZ
ECiAwNE3QppL7jXiK/Sdw8nNZXp05vXLZIatSREjOE+R+L7wcon6HlSNqjm5
VdYB/RS3JRMgtwdY6jnE6jtHTedzJtXfbTRtZw7WbH1tShBfNk91CowAxykL
Bw+arWPMej1c0LRDEM7EhT/IecI17Be9F3O/+cbP1lGqEt+dpxIIwJpE12jY
V7oAS+EWSZHdUzlaDh4ytbMi4o3hGxsdxFLY9Ne+XqL/JG2SiWsOJZUgKI3L
nurjH1oKmThM2MBJU8g0Kt+HYmMeRCcOCP0mEU24eiDxMXAP1yHg/Azvvsna
k8CIxWSupmwx5pSTgHUOOFUbDcAWzRW5+pBLLwAA8bkcCzrw1K4mKby2sp/q
z40KI0SekzunSUNhiyJbF4Nmn5u2eoTVLMJB0QMQEg1FuZ9eQU9Vi1NqNcki
ClLrGWyWL5GUdr7Z7OQjLk/1l8q6fpjb4Dxoc+m/uJYW/qLfuiHDoPjC26JQ
A1ySDTEk6g8KwJsnQZKxC92nWucPFWJE2SRu3OUDTNxenTenU6qNB0xwVfEn
DmclmT4pzXwBrAdbImq+4Rpxe67QYNSJ/A/ikvgY7DjhmOwXxa9CXoUlUv2x
nUqO9xWWPEzTJKjMeT1xp0VeI3NC+S3UsqJ5LDV7qTAHo8uL8OCTO+IvfT3U
484Yi8dZCBRYpOIF/Tz+ufothNmYUS1e2H+9L2c/9DwqR3CAfpEPhvxuh6SC
AbBaKOTBuepLeOfj2+J+TNIzyIw8Zes412KaGIdECUAIR0+XkjFvhsjGj8DX
DjbFbQVv6pQyIe9YgL9Xw318Fqgu4IdnvyNz22nl+W+yvX0Vj7z5n/2Tb/3w
2VpA7O4unPSxMd2ZDb5jrYIoH88F5nPLNIUTU3phRNDywEDtXhCYD70b5/NJ
/A5UOfyJmSYtmH9Irf+aZECxjwO4muWILHJtIBEJNRYvfKMhUFxjGti0tHsX
xk2hNVnGD9YLIXBYJSWihXVGw23+Nd+6capNp7P8EWZrlrpyTeRGGlKNgEkZ
XlRSqp1GvfbbrZHPGq23qkCJzxrMqXJ1FBT53VktXEQ1LULU0Q6NcaXrmylL
trIejGeiYGZxIuXjAc274EUAxIT0nwtTC/zFxVX702wWL+6Z9JIzyFoizvhy
9q/pPG1skDa49CG16TOKTy/lZkzn6zgq3x6a/FQGfS8JaiHUFH8rN7tiIdVC
yTuIcvAWUE07PQk5NMPhNO4tT0smS6nmL5vVD9DA0vfPZUlXb3w+BnbeKJ7V
dUvmyJbGGc9GR7Ua8K3eA9MPDEy9zQbSGD3vHoJxOveSpoH5rPdT1MqsV9b/
UmZXAh0IQimV7NYoQ8OlTMmsfckrFOsef3XZ9f+KPnSoK6xqeCP8FqvuuTtq
iK/TRViQTNKeZjNCxAelySVODq/2ER2OQcf7Yl4gSd1/p2pNrLlpgyz6Nz2O
PiDAO76jEmRCaBCmb6Ib05jexS7mFkzsDULyBRsAznhYRsuI/u2nty60KGgL
pPFSbWsV2a09TiH/nxAiO/fKJb+BboCYOzGMApGJdERUTdZjffY+3T/pIBLg
0Wi920xxmjD5cqyZCHrM7dK318vGPz0QlVQXlqL4oq7MQB+0xJFmd7TqBP76
b62hPM4AZkW1B6GYeb2WR5podTEGtQ8UDPAs7YOtRHIKesSJFqPxxePba923
VYyZnsL9GVjyM1CsQoksIkMZJFfOAYOfCkJ3oJ3C2+A1xAEq16i57t7Sl2AV
gpiOb555dRbm/N3ewIfYl7moS0i1UpEdrbFNTQAjQK3FkufImjAcwvS+ZuV+
iWfNPW1ZUPHRAH7O2SPs+HMopN5lGT4nMzQmj4RVIpEFKOAZQuzOTRx7w1WH
h4rKXZI9fFVaBQVqB8ZStSkC+p7Tv/Wb4W4cFkirK2gCpR1N28mu42tfNJ7E
nOUkv42y0Ck1W+KRJHx147Amb6BHTqMA9zUIO0u3Xrj6yCB+f45w7EsL2pCc
v8Yo7fyeMq0iqlPPQVy0ffRSM5JEUBKFpYQnoAhCP5Apq7MONJESvYnxn+6f
/aZZw+ktUvFeIqBZ6Ewlq+n+5K+jAgvHCHC1dMg12EYx/kUF6vU63VDB8pqn
Pp9wViNXYXR6fpzaNrSjm5WQMxdD8FgM2POg2cxh9xkaE8xbohVwjbjkXbU6
Vbi6faLIKl/e6MsiFl5Dp9yCceqYR6PWicsd/RTCEL1O6mKnNJXVr/b0W+L/
ATLciasDVA4DyuwVladciPs6r2XEOwiMdlFOqfAnaq71pMEFiXU+7aVgsCJn
QtBmMkNhVIcm8o4x6sD54tB+9TjEIlszxua2fTRDG6nAtBfyl2t12ptvXvQV
4jL6x3KB2VdLYgJTIswf5sbztyKa6+Mab0qqPRUke2+3ob5VrVxV6MQ3+47G
vcDQJJ+/zvCFWEvUp3I+RKVa3/jx3WhOqQQ+CigXvKKCU4cMrp2goNyxb+lV
ZuvagF2z6g68UKiRScB3/b9vuFbenL13PVWRUkfHbTRvzbSAd3XU3m9vpY3W
2qjL8DOlxmc+K8YOUpncaPIksFgAERkFWEjAaOzyTxUFVRXGHeWDC5SLMHHh
N7AGpocTvxPG5rlG1pGB6l1qH+ACFwkncm3Vq+v+yivU++r7sV2gIKhazbBR
UKHhQCVPYzokhLisf8FMVCqcdYt4kA/cl901HxcRAUlP/mrLa+s9LDgr1m73
Lt6XcK1nrJOSBPbDwKvjgb8aDzIhUsskqYc0HUaqHjXcz8V8gxDQEcOXQ2cM
9prXmGSQHpSU+XcVJg81+rcVqwj3KqKHUzM4qxxOX3u1Ncsgiwm0NE+ahWjT
uswYaQJIgMlIPHOiIaFdaj9NyFnd9ddmmB0GfZymJaomVO8eTwwiwDBXUxDq
653zNp8929RMEOsePGeoOoETUKMbI9l6oqcPAVrVaNQSvi8fluvsmy7weLCa
P8q1yFDdlqjeoKnhfBZdundr5lRNWsLzxyKZoGJjOhpMRKnxUtCWatZSflis
nGNvvrMgoQSBTa+6opUbH0ILsPR4eELh+f2BNIEJyljW+g2svxVNVndoZc6v
woOnR23ZCZjzgePoiZQ2NwSHRbL6Y383GEfbltaQ2xZBDqTwMbm0l1x6OQeo
kuvdKNh+dZgDeJiPqvf3mpAPlvkUHSWulHAm03udH10X/vDAljEehnJ1wd7E
5oq3A/7yXJPzec/FLCAERFGwzftxl1sbAEmMxi7puSVLrEpPnk82UwUKt0SI
qVoT83DXKJJvxSJUhV2shJmEsdfVdAc+TNy0su2yAEzBI1RwGRZfIYRCCkkQ
3RY5VcW+VSXOBIXUFq/YDRaKP9K+Q4+W6jun9puPK6NIY5PsR+fKFhvYwJBz
EnvvX1OVoFIVGgty+gjyddB9L6S2myFd4WU5BxKGWDymQqn3e4D/qg4K7Vz8
aXhcZDNT4FXmK2xtMz047VNDpnxLbZwfqiLLatbIbrBek2sT14C5UYRVk4Xa
bq0CflXsdKyUQm6UXLis6Tm9xiSqZmbjVAV1t1Ru462IXzyYr4h3pSl0V8tj
kcAacxdJhfYdRhB5X+5F7jdYXS48vmjlsnCZjKku9VVp2iVPApGOrhw+Gw6n
tG4xrfDs7ib007vqwqCerfRDOd85t0lrzg8seqZKnQjP2q07hIr0CrSDH8lB
DSg39Ex+7aRAdm9pbSm5LNa9IUWiG84WkERNlgy3ihMXRb3ztdz2x6a5SD7P
ZRICFCLTtUQj9ph19ZlPqZF4s673+TgR0MGsEQFqWHq4V0UwIXNPgYNP5oZh
1HAORwSQwxQU5KK3AZfk7+cPd9qhoTT2o1ZbLmbDLCLab4JvzaUHUjou8nJx
LOtU51nOQDgWWxmNREyBeWm4Vy8D2iSZHcUka5VjU9vT494/ffN/J6IN+T24
N3/1SF5Cq2bMVE/xsuUBtMPPsYkaLm9Gt1rSBgaNj3IboEj0I98EaXb+bmN7
VBPD0WPq4rZiKtOQXr0p+4Ejf1b0a56RWBadBz1k07GVWxXUuPJQSfXD0Xmi
d9k+o2An7EVrldLvCy8pebHhQA6Zd6NMT6gTv28+CYMWLUiSpKb9XKSXIYDt
cSTnfV0pLMRbDhyTgvQ/kFDpIW/cnZk8wVD/4/PQhGBqt+5laKM4oDsC9heT
BS62fUXGH0kyodGuemt4Koub4al27AkgQtS+w70CDvD9ezFv3pEJ1RRXGjr1
6wsRqxzUzCSMKZfVdkd6sIBCCMU1AwQpqd3tu+zwEfghUTPk3n5UK4sQkknU
Rw35ogl770N8ok3sQe9e5b4RRn1BeGAE7vsewvDZMYUxPCstkRA1Hu5HNGAJ
u0ydmeWzru5xiew869aFhZRKqGky2pix5JeVz66pNGHNJVwJtAnH3xpjhuJz
lOJJQSbKYL/Us6Nr6ZVdwL4nxz0UpTcbK9nD15Xavo52m9/IQ4eobM5kQSho
H0BjZBrCxE99yeTbWfEJGycPJwDpa+zvXfI0ewIlW6gz9esArpjvCZ9yOBFC
0XK8lOO2239CsnqU1HNwJZTnSgXaBXmtp4seTeYCutycYpJAlg0T2mT/RiXz
1sB0zYfFDc2XcszstIDdWHgoLwjbKIt45nhASUP83331lGwf6Wln1g3d2Yf+
W0rW9mRjspeMpbNYdOzpmET/YGPBk/s907BXSwArqv9RUqIe1dcLHQUx+7UQ
2/aQLYtbW1rWOOQpU7rG/H1q43l1XNO/iXdWAtd/gbt9nYq12U5Xf95DR52t
o8PtKlKvAQ7ICnQtY360VCANy9gmnG0EG0N13Jq7UlMO0bXt1HaDk8jGOTqV
lQHonhua4YtqYb0yQUw+DjRRH1EMznyw4l/YjxuE64AqVXN3KubR90DJImJr
+61SYl4VcqJ5fYOWtV97BKq17vILs8fBzmiqs1e9ciAfr0VaAo6UZYXv6K1h
Kmw1YKp6VitQ6xQlOvqjYK18Yyfgqifv5wCKD1P++L1so8NgpOKB41ffvx6/
lVsyLXXFubbxALI/bLoj9CwrxRK5mSscsCuxQ4vjvlcU8jS2SfHAH67/RWdB
mE8XlmCQTU6HV8P4rBmhW7O0sUC0XMKAgvjAEDuzQbroi3lVpMmANAAIHYG3
dHJyA4odzbIIPPkTNFcJqpLkvfnnVAwSuZfVX3c9PpxVSC1XdDOC5RZLoghF
SrLcFiIIpeHnJV0BofkcBox784CtL+TfXuvQltCPoU4O2FMqn6sTHpFVlBaK
syB4lj3aA3XqyX68ycN7EVj0OLu+prXGrXGWbwgW/9SPjNKtpippoZmM3ZaX
8PtiSsz2Q+ESuIJN9T3aFMUQK4EI21rpBM7/W2roKVt+mqkLVkDIdt/Canct
jB7jNzd9n2EnKRs3UzVWND2ImVLwYFrxDAynYhXfBh3XUE5dzsSLT7wHvDxA
rbNMNoiC8WIdcmifD3VgkeZB6W93t7W9nexrR0E7aRYM8RSYQnwHeihSfqBw
hHUxGvaskj2Okj4HAUkjsUB0SZPZw0Xly/Yg7Xj52HgMauLw7dyCE18mqktI
xTcT3HJcWMdX+rtiGB5X5SdI4GUY84d2a3zQCXVRVT5LfAt8hHYRoyX4Abqo
dnqfS+r6fq9GZ1/0gPnuItAAOLpZmn+xIUXfDSDWAUKHlJ52Z/uJAY7/4jBj
DDHwjFx7ltRwdoHUNcn0pTufHveL25G9V/zO7oDJb4nEhktOJvp9+ItvMupa
pfCZ6MmLuD+58l8FJu26vxJ2Ciz0OSnneMXQ+TOY0mpbVgWO03iRnlrrlMQb
b7d7tvhDgW9U17JSw3Q/7dZDQmw3ssgq4iZbTjEyVJyXbhd6+6mlwFByaJwm
UVES3Gg/eElOojHg8fQJ8uV6n2TFWPWahccmpzCJ/pOQf5vC2trWW7sS7260
kQ/PdH4zdAiREk/t5CioSvoPUiVQyZatbPOtN0Hv/yBC7II6PRvQPP/T18h8
Oom+uc/EelgHtldO+EavtLCzHSVCoVz0/PwJp7TjjBrzIS61HRRnPr8MU+BM
kjY63EqhgjDGt2QsDihVHMwjy1l2okOT976rsrFUUTVX7bGjXN7WVlo1xvyr
Mza2CSSDrLvm1FhL27HkzP0GFebcfy7PLG1qB9N4VVQ+rwRCRdtkPA4xQFrK
qlIXRzgPNc9rYcgTxLooJc2+2/lMD/8TCXx7jO4kQaqM6XNUkm4BqjoPeSxe
66I9VX5Gkgt1eOvUH+BsH5FrMyVe+oMEg+GIFBpZ7vv8cfkyP2GM/nSYMUhr
esImQqITXLTkf0Te38pv0ps3dj06wWpePnoN6hkw36GpqRV35lAjmcecznpF
jt8VMe6JLSptSgKeLdFvPFbzsmFKb0zvlnLN7LdjsEiLGXXOawstH6iSGjYh
XBvoRJXd+H/O+HkPoI66cpXExtlTLPtZ+zXymFaj3VpFqxbHIuyA67VY2L0m
PbDQruBl0ynKYF+w1XBX8vhJyy/oCPVsP8jxZ8YS7xiKUjyn3e2uIKL2VBtX
QOF5/4QgIVmjm8iBSI27M2tG1ErxebA9JTjFrlpBrjUSzD7zfOsu9v4cZP9d
vLT2RbivQp48MQYLe9ybQ2rnPpx6pKgE66sgI65Hu9Tt6efbdXGyGe4PSGx8
6+bgspWANNErLhXb57e7G7YnYQuD53pvZntArShBYVJw9T3yiofXozCnQPwl
uOwPk41sg4h/PtALXMRJTZ3JC5+E3w/Hl8hJjgEyG0BlRT46rByQEhlAx/e6
HhvIxE8ZLY/TRcVAOLUCyO05iAUg+9atKty4BWxCK3v+HmXfUg5BBspUx9a+
VKwo4XXKg88PzHxqljFl/Cyum2S2zpmQYPowbMzpI2egjkfHW1WsmhcQ8L8b
Cl88BhwSHpOURDt/D+kjYr0swzIPD5+Y9w58JX0ApopNFt/7KxaHKhhn+QCx
VkCtIU4XtWF4zczV/S++9ArsHB2BhUS4O5jRXpL0Otm+exIoFct4Qu7t3Xs+
zPbakMCeUfnTrh+WkQreubtcP+c+8K3iRHpgmdQHzMDkrFavA8Mg79x3C/Iw
CkKuicS7lkOuAP0DcSLy2l6K30yHFkrUGXyVRa3smCRjUJ0RlgBSWTyDWoPG
JijIUHRAFRdYuFk6mdY7euLoeeaCgdh3pzk4rVbOgMw6Vkyn4Dtg3ZBWmXCE
E34CvsdWseq/etn4pnqsCZc6uftAPhCzFBR/2Znw5fm92DiXjoNlGhXVPlma
XmhZUDWBPF80zGJZyH4y50h9dbRRgG1IVA4EE9q23nfeqxQUZVdhDgySacNx
VgL0ZqokR9aEhQqn1qsMKWqcutiA4Xruc/KG/MssVOiD0INWeT5n7GfSfGaA
0iLUZubh8KdhDsAnthfVLRlKvce0W5qJb5OTMfp++2uym65d0ppwbawdSFRS
By3jMKbdyjdmhVvgTsS6K1zYZxjBpYdUzUVMwkvaBesEIa+whRgE9k1U7hbQ
bq7g3ylkeA3JqORgjxEqst1HwqZQL9Xz1oz+r7QKcS9wmdU9rCiGQuI2zv0w
SrR/5rQzc4WFBIVXci8mk18mz4kW/qYnYJe01v2/2ISpUjvL7pz4hV7rdbxS
Xj0wNqgURSquNH5/KpNjga4SJrnZZINKRgrdnahLyhZ59Pp6Ca94yNoHurx1
VrOMvfS89qCXUuzLVM1FBoYBbJ4Kgng1uM/QaikdSPVHk4lwWtTUoQjvFG8E
fZVOz4NZHVSWqNFATlQ6ByopyiRxu5Fk5SsQ/bs3aapYmpewoPasgaMltZwi
n4YxIkkRr9sJKNPXgQAvmc2+Ajgpj2jXVO6UlRwR3Zn8RyibTotY0l9slHzY
utoH6CkZGfVvVR2FujM0LnSenrpPzug39cuJQUs4IB2wPEWpNBQeBOsWOq8K
PQXx1aX0BMKoqSnmiOlTkiKCI4qncv895levYyCGhDeHhrniBl1kuO33EJA2
nHy4fnkBygZG4Pgn9GkHHAxFkmZwS0QM/Kl9uHajvzttnmCXDXkLqLo+yomm
tXG478l/WJ7GkIOk8JNuSfUMdWSjpqczBXUe5OPrF50vt/94E/Z5K7XxgL9T
5ULHqUbzNNHLXR9UIsliODHTaccoHlDVYyJypq6x9OxqPq7/+It1Oo1KtDUk
yhMVyFmQzvjFYpC9gGG8HuDCPBcNIlItkBZ8gKZyE4rCqFA87VxzFLg06HlC
OzOqp2IBA0JlfMkK/scaYRWksZ7FfbS2q5SZmaqIt6irN0U6qqZ/coI1VA5O
ozUOisQ46TQba61RvflD8hjHQYSeGToAcB7g1fNg77aRnGsyWv9ZJS3Lej1L
+i8G5SYa8DIwYahb/8xtLYc7kmggiQ/s3JNZ8gOPtC0KIEucg+84j4DXHN4l
+zbOSJqRUaNRGi1kvto8tncDhOa4P6HKlIrDWzFcDtI//VmerLG6PJ/PSGws
SwkS8Df3UTVmAN3BXNXijmJTxyYiPrvWC06KlpYIB6Ct3R5b0bu6+UDIEZyh
zZDCNrijoR6JBtaaRyfrkOIXgD0p4vSBPg5VxN1If+kTKTNJUfsiQ9fV1lRD
4RVGd4u7SsLW3M2NHgLhNvOuCQutwNlvFCiFOM4nsaIJwqfc/F5s5IaskzXO
VRWlY85SyG9jZTZjqtdO0SsiRJtD7a4StIGrVYlNEFDpCVresFr3VThGUKjX
JpsRJ59BXHJK1z+cMu0VO8ZgNWenbJv7A1nMlL2mIFaQ/I6sqigsW73qOD4b
mtFBvfo8tNbuvLMT5pswhbxLrNuLepAVZqWQvhGMkkwSoKvOnC2S3lbJpcbS
ohP4F/4hBHz4Yq8iFkSoxHQdB/aeenYR8XiXnhpTu4JNHlYPLcYY/WUfTdHo
xvPVmIUkadCjc0Au4Etm6sQVH8HWI11suYcH6WylzS9+Q5Ja7EHS0doKo58A
zHMMWz4QqGhbDe/5kvFcdpnYAlNM9nyRcnN89lrXMeYTwydNEJDZGlQI18gB
iJYZhnOJVwKJqrs8TQR/0us086It65WiD3kSwyuCib4wUGfOpCrtQPPS4usP
GgzyXzsdg2k0jO7ebBHyqBO7QQLp8cT5FgFi2G2D192pRL74n/RQ/BY7FP4x
i2Cei0rWfCxKFWTfnYzgOI3gUaBN6xxKNq5f5RYxSnxzCtqNnYQ8IaVUTHSu
k3MRxSbpgk5VHZQaswjN6hTRSSfYJtqRjU7fey4wiTaDcllKCCSqsAd2lYbe
K2GIE7q0BeAQQT4mjIPZwMkqmyoOI/o1lssAFLP01hoNyuUMSciAPyJt0Pzl
QaieJLTjX3TwEFBKavCjhWOZE0VZWqNLf/wrwq+xz4ggAR8MydPvHzKOfIqr
cJwLMS+l6qV9F+H4Sgq30hZqMvOODRB/By+grSKycSdb50HTHQbQScIaH8Qo
afRwyv6Fy5Dr7Elt+rMrfNfCKgCDF8GO68mCdo1+s/UqOGpU8BcgT4Zvfw+z
TGt3o4MAXYq6wKcmvV1Ozso1rwkvCumIP9tPup8j6Kd3pkLq43fEOrpa+h4b
swV9VXK9FCF23UJc2TuzEEONF+DeHJCbwP8Sjo462CExA40drclLGOxHL4x0
FwgZORi00R/B5HSLHyS+Bp8de6UzckfWNoHtBfv64ZIE87X5xz/sk0XdYemN
RvaUXiktb+Goe0O+/GzPpsNsXgHrAzmGjnJ8wwR9qfzeQVo87rsDGuedp90P
paR1QnPTUf2D41L+Eth4ANdEqtcCIOkQgBZ9RvR5KwP5XqIjeLSFUTftkVfu
l7FzHF2xvl8Nc82ZsIC7B6iAAXLBu2kJCtsjPv+dHdMmIwnNhNFDatJPnYg2
0xqIlA+siZeV0GtSNJPXBxn2QT3J/1xSDtuPwoB1w1ZX0huo1GkZ6kxkgMQr
kLRFFv02lWDV+wHYXZIwZWUkg3Kyu+OXc6NxY4iTxNfN83wXwHsiFHjCR3ac
RZ3kxPM8zWA3bftnM7eiMFayVsx8ow4hBbDkoKjSbKD5TE4oVSBrPJCaeScU
M7aEYWuZZsg3WhPsdgR6zOFKrGNUfxM5KcxEU8P/V+S6PymdBMvjw+k0s/hg
85pg5GnAGhzHwyvb7OQppEWZdsiQSStem28XmsVCtyYXVs4fnn6sZlzCCcva
qjlqHl2GReUN/xydimj06DL0TR9LI/C+16H4Gk9QaCFPL9MA5M1srfvXRK7D
lekiaIkSHtnuRjApB3zVd9nsegaGj7+dS0ewWYuM7m+dIlsU4Jzp3OnZNREb
lxkLuG1DXd9tmtgotW7ewrpORzfHzFhZH4nQHu3eS7GqyGfin0EaPgzLILoa
e8ElAzmL/6MsLqp0P9JN0yzJymRkDIHjuCfar1Er4tjeC0tKBLsKSvh9IPU4
MKmP7LMYhQJ58Bk2fXrMX3icABW/AkmMjeu10MA320VXF6ono46lTCV7BNb4
vZaSf75SLQ4DQ8dFhtdv4us1dfDYrK/PiuLkxulyCFvyvHxqM/9mZG00PPWt
1Vkl4IOCHCTusiE364Brp7rmtODT+S4gOSvRU7etgI2AlvyuB+jtj25Bt95O
QUl4+KPnv4mAmxefov5VN2fW4xXgIt1P0A0dH+ShTD88nAc3JaE2oY3fmptN
EBv8S2H7sXl060oyNF0Kigv+ZQFTAPHgBuWrOWWkO0IrTD9HMhcMKwrYc4JM
kSSPRNOWQoB1zY7kTuDbv6/2ceKRiVIgA3CIl4J6ojJWVm5iAE3nB+tEfeoC
A2VzxU9mTTtggNah+NmVtI+WYGbjeiwPuDhC++VSaauwY7TZgShvBNk9BxWv
axCKkfi+9yR53UE3lLZCfJ5IhBY+wKTpw36LAozUdOX3hql7LWRMXtAVwf4T
MbcWlS4AesEtkVaQ6BbJ8KxRWtPA4mWEDXZGGJ2b2QwIuTJLoraahBjLr95j
ZDH+HU5bjhUJwB60BqzPTVheRB7tmLwqXQgW96MsgQSci/YfiFKaily8rrtk
5575peTfAuRr0A+74i65bv11gxoWeU5nXu/O+4LXojuB4GsEFzvNnMh2Epw0
Sa/QGVmCzug3sesIhmRhnh8XboNr6DM626a7OEc/9H+8LQFq0u0wyrGYuydG
AqqY9drb3fJA8va7bUwJHvJhAPAgHB0zQpjvCugP9Y5RpTikVGtQ/U8qi1Gz
uYYuvWBN/2x3Iae6b0C2klwa0kDDqbuF6BL5anjUtYOSdIuQ+ThWHSJIUOD9
bXp9RPwDSiBQ6Nmwc7vx+bPaL01EeMLx/oyjHliUsUZMLd+b4Z163BFXEI7n
FYwsvbzQ+ibQgVaPMXbfwqDneYWbjfs3V1CwF/5mOiNe4cSQdVhkXqeoI4LC
LLgR224R4Gw0++/TgXUbLmwi1cZxYYBw8fdm1aR0NtUQMolI+/qfjFicwtpI
qlzqh3V7LP7fb5LhQAd9sAxvL2g0RvTnhY7guuhkIh89cMzVObYMwiYHgWpp
ss0SoDGG4B8Skqy1Qf+eToSPI38+37/WztMK1029+adNRd7uEuJ5s1jcBy02
A44BlvwtFhii3U17PL5eU6Zh4Dadb2/0zGJCRqVMV8oADSaDp2LajBp3zg8G
Kve5IVJMkXFvoAJCroXfSPRVxily+tyqry4drFmMMiTl9wQEVOhzNUOEUmHp
3gZPdl8G7JTBIRUYrz8LAqlM3NPy/0AhKyqXtCRuc8Sa5VzXdUqxtbuftHSc
/l4pLBEi6q+ZpeFcAuVzviQ15GjgoL52gJUIPRjWvlwj/wWtcqfallylw98w
Md3O7TnXtshLJQvPQTNYybfn3qoOii+t/FbFVF8F0o7pMr/G6xsC7y4T1otW
6oG7YiVXjCOyE+49db3g2R18Zm7ERDnEArfwlMl5MrHP4Oxuf0T4r0jik9o3
BuuIxtvVUOs0GjYhrRZoHaOXi2NH5BYr3yv+5V2yEohakMqusxsVziBpk/v/
nrMGZt4LseKt+Y0MH1iBCeFcRdWYANpW1wawBBAmY3EQCCWAFrbomW82XJBi
IKuHWgqmi5q4u5Rw080PWKE4fxLsX54bI9EkJ1d2NlK9f3t1aJZFrVehhV2h
ru8f7AofWOWGmkR5lUDfwjd/mz4O5NvxrpKJIukb9Y9/rpsB0wbCbnY3zNt/
R6bUQmPrjXcl9OtsnHby4xfnTaOdUZyeaa+V5Bds2E8hRF0L6yNWBCA0CxmE
W8DPJmQ8IW87o8uVMWPtflFUdQhxBXQhE7JMiNCEumWBh3hCWQDC5bEofDm0
qPn0yR00rTMDRZFaGUDea8l3CRdD6xqxYyZzcYhxlGp5OpG/DqMfd0cplDMH
3asLtiDGc+kw9nKu2KCoGvijqsozxftg8EHDFO+zNbNCGdv0S9qb6lcmGyyO
chr8JSYm7c3eXlhfLotNckH+YrgYVtGYDxtkj5CWbTG//76RsnwFUC+OX5/1
MyrkWb+c7Lc6c/CDK3GfIY+unhxjJjLQPGgL16+l1VsYBHlZpJi++wMxRrCa
8LLRizC1WK5wogjH4SKNL6hRosiUIFC2wNmtaza+z0m6VfPNyTI7IKXg52+Y
Q1sKZy5Vm3SL/ZedX3AlKck4psrfGDw7TjR+K6558lVi+bsqFsocIwAO/kH7
nHNUqfvfhuso/EsLNJVdaPJj/QqLBAss4VNkSXjz0Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErL8wOibl5c00LZ/tOrPY9pGyvFs9pyfKBS/903K7mCInTHgU0eQ/WLoUzYO5OGUmDEJGU2Ajp33j5witTyX+mN/7QYKzy3EQjxQlJwmOezTo+zmunM5Gl83qXIMhHKEaFWhBL/EH/MIs1+8vjCZuNkaQyDOUSqUrDHWpxe5e/66T/qRAUqmJtjFTM7T/hnsAoQ5b/Wi4O3ZsyfjKf+fIjs+GISEejKiqKYAUinsGGpv7VOkp/xRmktCeKd2bQTcQ0xtjTueVc9OEyTgs88jorvYFHHFpvfKuLShZ/PJ6hHbcP5qQfIQ1pZ3z7MCIWPVWcooKGinnkVRrt6w3iH3TUtN4RpDdYK4HSgLVts82KGrmuTeBtmavQLdV/X5bXIBky81jF2otNF68uaeWtiVFORTX4issTs6ZlE8DGhdGzu9OCsToSvsjMdfmEPhjveFV4la3/mZTku/iNABmyk/jNuP//Ar+pIx6HxiFnUImd9j14wt8PXHcE2r8+GWKEOI7gI3N/ydtRvJGvbhjEL70x4cnkFyQNWAwNegJXQ7Jw3trHoBkPWdaeUjLxCaaN5I6N6FKtcWqIL+RloSDvTFv0zK3AdPKDkkiUEeA7bQXmZpEta29qM/8KI7cCfAmCbQ/jxHXDvc10Qe9OCSDsYadpn4PKx20rT0d87WNENfv+ENLdM3XzeV/BELgpxlkpG8kH0lSWQ+J5/cjuy1Uw76Jcinsc6qevI/kPm2MSs80e+6lfc+foyKM5lVrg2RONqnIjfF5wiAq/PA/CIZrMdeJnn"
`endif