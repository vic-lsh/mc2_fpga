// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
li3YFCPzFyYCmn3DLXxrq/XHxCCIoUVMCAKGr/QaqdYN0XTM5Wh7S9bVN5ex
ORtSEjJFveicsFHxwE2+9jtg6k2P+FK77QWUTQikBpeZsI2lqmF3W0U6Lw0f
20T+FX4Gea7FGcRwQ279izA1IFhGH17Ylou9CVYxmSoBv3aac5scxZbitONX
cDIIh/GGhs0rSmXsPj7QDGB3x/aLnuy2yDCt9O22C1RgeQ8ABopoqD5N8+Q0
XT/J9JFF7aEEmH+IBREPrZiKyf3LMjcgVde88dq+UsQ0O2hD1sEYg+HFuV4e
1fKEVACJRs61++C/1GswFEnE91PgXMqm+M8mXrSRFg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
inW/mnrxp59GrTejAQ8PlCOakohff6gdCAhrTCak4QPgDQpf0cjdMnvVUPSi
AENOWRz/J52rNjPeGpYQVRNa3WAbrN/APAS3WqpnJowlEq+wGe6g3ectHHL0
E9fLqhppAJ+6rstLgumH6qy0Tun1FISDa6Wdsnh2MPxRB/YJvB/4zQY3fumn
MUM7doIlb2CAm41jvlF8rzVPDs2NRyxSaI+sTWTwE1+IW4Wm0S4DJHsFxH2W
RvKKDVHu7eZtvMeisg1cEaf78FO3H9esXyTigiodVawqIjhT07XaTfN9lvk0
ApnLFeTuNUi684hy9kBSfVFSmtw9loGf84L14d+Lqw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YgicY5arX2zp4iY2vupBNFlxkDmA9/NyOlh9Mha+xtLRkZ/H1eG7/4NU8Nze
Br1KEIpcLTs9ANv2bgQsIBNquG7ksUQxsW/bZu0LnLgr/7w9+575rslVF4Qi
sYQuB8BWLWQInYzBhBex3yTmDQGs9atNOQVRKtJJmXG3cFWjIYEsOcwtuOAa
pI+W7Ybh6m2468F43MddE8psWe4ZSIEVaprqEiCFUBLD6QI1R0+9asP9gp3Z
2MgiMIomSDeO8+GhMbyEWcsv8oISA4cyBmsD5fTfEe1GrKFtSRzkvm5x6OLa
x2NvFm+34BNddL81X4n3re/AVBbpy8OXKCABPuowXA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GenxRCSH685MfkFv1+fsfZZDWTJkgq/lHGlCN1b7UMp8AShfsYIwrlGi/h3H
sfKyT0gBAXuocKitjeWZeYaDGj75qfcgHhjIPZhRU879lxns9q/5vdkySY+D
i1rSBzShrJAw73gM+vAnzQOFk0Tq2m/f+NYLNlmWGofb/yF8LJUwIUlhyhXm
oV6F5UmSLL+Jn1o2PuQWgBVOqLpNY1wtu6LYbzau5AemnHG42wGkmaTnKO06
1IUtl1+lN/CTf9rI86MHlnb3qOvroXSw8nnZ8N2pSi6iZvbedjLi+BFpM8pF
PvV+odPKT6uSxNuH1hZMknmGp7DwbSvF2HQgmHV4NQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cOm4gmgx2P/0+4MYnJfGibNZ0wvGYXC4w+j89zsloS4BNywjiGvxwV+ASE5e
Nzusl2FmcH/942nQstf5JjTqkWJXLvlJshj2SYNPhM+WX23ot3znsywY0x2J
XcY7q9YmQJT6GakL6ESndHAqXTpnvy5XNIZiTaeeocT+DY7+v1k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lPJ+o34y1BVaJnykomiKxm3ZwDzID58tRoShkiHjlEhwcylsC+bDm8LQpOq5
S7bMnOf7CGtXBwMt6ZIOxJvCzpwVW0wLAdwL0XrqUTzTh6f2AveR6Z/GqOlq
ZtfczHYpSyrOptGIUkqFKgHSbBJ5ndkWSf3iKfktsV27bZGUSFCbOnIZhMbf
r74KxGPXUf4nc24xbr1x4hahrt0qGwR67q0MKSxRsJRggh4+s1m8HYFUuCdI
qezcg1kjjWa2E6zeHDpq9SpCu6OqaWchvqHDMu9vG+d4oMpTwLTDqv38H8n3
nZ+TYdxUOo9Tfe/oT+OhKR3/FoqXk8S6dlve2crprP7AHMohnm18zb6mADWy
li4kX1UT/lg33FM73PjkKHYcBRmDHNueEWFsxEDgUuHUkqKxDhrT+NTfBT8p
pbhErV5bldZhcN7ad49h/xL5fUvDsYRgnjA69mCWKh8a7ThwQ+27hVIgzGJ7
MjvnyeB+6WwbDMR5FBz3UjBfNIEmDTMx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KL2uUpezZvUdeg06oXLYkLUFTgR8+aIkdJKCAhoeut5y6aXlkQQKpYzMBhrD
IHUEWHl2y6aF4hEdL8W9v7CApAD+usK4Kpda9SRym8gVsUdxITgFi87t0as6
3vmxIYfZk7zV5kwn/cM94G0DJffrEkqcBUucfRwda6WjJon7ibQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AN1o/WLrsTQ1f5UTH8xaByu8gGA4mvokxnRdQyCMSD9C9K/NIVSe1LIc9gCK
2/4b7Q5Bw1Eo3j/KUE9wQYqDqAeIwGg5D/e7nprWXChcSkAbssk3vKWdXmlE
GKNJU0UITNB1WB/NMsvXR4HOcjbtTdvPjkNJpEchHIK9K+1j9Ls=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9200)
`pragma protect data_block
wSZoAjTZR9UR3QgaJ2UirC4MDZUi66lIUzMD6xom7oqxYuTOD3WpZiqMxSFF
PP11/5x78ao34bE2hyV/gITz7SJffXzdhj8kchxKbboxHg5ZGSvyGLPe5I26
cAdGUwIui1yfrP3EGUN6+/Fpjql0gj1jpXMijQ1OUQPfk6Kvel/d2ib1ZkV5
8nA+4CInmOPbTcsW+BbKGhPnbeyP/dskMTOEAFe+ce0/jZO1OHnN1x+OkQC4
h55byQQ7PnSxs9G5cK23ZvtUOE75nKgUwiIfSCk0Vaf55XxfnQLZABlnc40v
4ub1T8o6htmo/ug/0777az+9uucttc1f0lDvlOY3YlIz4iTesPL/P7bUep3F
gRql+sX2d080WVRGgHtieVD4/l1vVyzzfS4a2vtWGZK3drPlkD5pT9ZLE+uj
LtaGkyTkURJ4yL6RF/ZJurBDYcPcTXUg5g5qzxnP2sSenMl3Y8ZaX8SHyTKi
5tf5IivQly4MdFfu/N1hK1VDpKHHvOaMeTRVm5vKm+BdmBcoTIEPdr1mpblq
+Zof2Qb0GUD5BJ69mRMjxhuq9lfbf5kRNiFaXcfKZOi61Dan28B6+YKkNTqJ
ag8IjUAWhCPMxackBmRlO0eMQm1u5SCMps+/tym8A14V3RKSdkzmxWTqdQQl
1KZVp22hgYdOvHGP2gu+k9QA9VpoEAzrJdsEx3nHro1ho80m3nHlgyrSxe4w
uSTzPXlIV6bL1aL2AB7iMKe2Hxs0hpWhy9vIcSZB/AKS2t6Is5mwLrDU2ldJ
ei6lBCGSi4boiHHDnTPIBM+MDnCkDIsjyTznj6PQmiWTs4iu7MkOThCrcvBQ
LKLFrwbjPlnL1QxMryPQ+LzXyE9Y4i7WgjxxKwJh4OAfpzFCIYAFl3Suf4FZ
erAvr20Bd1VLTG2KU5oxM3q+x1qAMS6EpcbtC1nJ97exHCHEtjZ61KsnSzBC
owvB1Z+ldtIAmMifPzHKDuo1NpfwRAptHIjDs/khkVR0EwDVrcqrKRPfiaHz
htsMy+vwiwE/Euki9N/UI0tSESStT5CndwKGoKEZiRv6fMEcZqalUpWbyiFF
+l/Vi0gSzTCHnFmKYinFKFrBLB1DQ2QOvrk2yNVqoZdsWVQBJSYGmoCKH2rf
eNnzhxzKn0676p38W7MbMqUGYVHSiviweZuk0XWXjFPgsMY92JnG69yfhDwg
05FCAVyu3TqOsypUdeqi4PMrXqhAnllKXBky6+9xsk++t3QI8yFgSFbneFro
Ry4rIfWtioebfkTeNCkOD2YTYVumAk/lkIkc4NObYMLviKIrXC2QlMK42Luf
mZa4OVuJmYhqvEDcNZHm9Z2QEkSWuZqJA8hUBDAJTu0jmNl9Gf0kaveivx6/
Xxd0gD0RDDCCSLI3RuI9kTnit/AR+ojjN4jT4+tmC1v+U04TKAbFLSX0jvf4
9LnJufXdh5tpOQhaOlg1nQsJKHZSXD79hHItAespFvxW3RW2SzJyrLz9dc0j
c6eE0HNKDrYR1hvLhLVT39EpZw/8lLAWmSAykyIw1QL2CF/hq2I036Tak4Cc
Z3s5i6YqG55ZqXUve6ItjYSJHQ5joia2b/L4uk+yeeJkuZlwNxhJB75sRI5t
eiBHZ7VeafGnjLhEITMu8wz1P2/Ur4U5B3Bkq8yIZDG17jk4GilM2HhmbiVP
ww4IVuPxFvJOjvx4DaEBzZKrnDtGP6NbDBxtB5s3KMdryIlllCBiDuh89h8Q
2/rJjyO42hy8Qq00a86yNa6JzI0E5cdMo+jejXUCky2oqhx7lBTHzrBTnwPp
lfPWu2EITC1n2nmVDt8Gz6Pvjj4FvzxaAtYsGb68foOAAuRG+r/1VXuvPUAj
zyV5wx/hAfB62xgWCZ/QM+EbEpWXZAI5TC7j/LWLwn/Phw0GPd9mZFFUll9J
aevu2DarDvGzoh31EicpC3u3PGekbL+gj2HVvu4VFV/VKhlNl09jAG5cau9w
YkA60ErKoOiC1TebCGKGk0gNTcNawrt3kIGJmKjxLsAbipcWUj0XmB1illfi
IRfjwB5mbQh3CIBSC6u4DiFhprijUfwdIyy/LHpq46cdXKyertKAJ1QpD5kZ
cCGPuIW64NcDz+NznBf/8VDgfwiGJHmSq2Vt5xNH01HR/QSIlJ89gEATjW3L
uErymU2ZQOh2FiZj8I29gGcZOgZFbJsihVjXBzDsq/1idOGpego6CBcOPxGA
iWhqHrMtsqc2U8niCgYJvDOviIAZhuOP2aL4f2IFhtl5vKy292fB0jNsnT3D
Tsux0xKLTESgyYe0i/93mccWF0bj8w0qY8GwAXfAeGlmRChbcYy3VsNFLKkW
eIqW9xQs6qK9UUS9yatN0Pg6cu8uuEXU390ql6lic4v7wRt/jkp0VGfrzkXH
rZOQsGJX9S3QPY1GvfAaC6/5LgclSSlnMA1gb6J4FOAm/JGH99Wr4tGf0c7o
i++lhYesADFqtPrKLm4pZ0IZDv5f9xWp3QJGj61NCqfo4i/nT4rgNc+ixEA/
j0V2+3BJd/ZHvRs8/sidG5wsDMBiAxzDBrpN8d1KDPVAE4bp59au5Cxzeo7q
8crbYC6tko7N471v2B+Q9u33CPxWBu9MzzZJI5UCoC3iB0oUNcT2TJ+6ywtJ
SMo+rlHJtoESDHDiA121B3tu+8ozsGAs1g4+VIABG56LMROS02sDgTMAfG3c
p8sEXx9L7W7dPnL6cv+h5jhptrESYGDnOBVfZ0RzZcrydOYcM5LZC1ylQRm5
EawgvLinbKoDRTxrB4atUFl9EWvqH/mFjSZ/rCh4l3/Q0xQ4HY62SxoetSwp
h8xtZtGq+JrwKyK079cQYLn553SiM4ryzvmZAqO59hDxqQYWEzJKGl4mB+zy
fTWGpdqeut42PNV+gm8lmj9EZuhOy4/eUI3yg7fHSZ46Gq8X2zxysktSerki
40UBmxXThYyT1f2DXMw3u09tL/V2bugytfi/ymL6PnNUcasi5tES3DDfLGGA
rzi2gZRNsthQqEuOUatSFDVSFqM11YFAMz4yfDT8wYH09w/ptp+ZPSwm52sP
5pf6IX8B2BqNzsH8mABlS+2Ypkrz97zJxzVQU5uIUXXIdZoNIvtFQh3sFnks
BS7iHHSV3pfiTkCLIr7AYFuTtckAcQG9xq+H+7c/uVc9U8iERzeHsOkh4CXc
vqC9O1a0qyPAH7lMQjoSBubiYN5OUic93VcrcKWHh1j7Jhsv4fRSF5e813I/
nOFjDZXiKnub7iW1PvTGGBTfLBYJ9G0s9RZUZ7dQqfSrG4pk4ClZytzjslbC
OjBv4sxCDEoq/sAYoqx6BXziI0rg9FbdmbveeWznA1qgCXTjYwXzg1mHUNkS
s4+RuA7IvSbktZcMHpXnzJGITImnk2u1DGrBvbOha36iZpCf92RIlbVZK3lw
rsfa80hT7Uij2H9UlvaUY0lVYtypBflxeLBXrzM7v5ogOmHHAPAyeoIU4gqw
U4BDT0P3eTJPbBX63mF3wRTNGJ033x8IwGwYcLeuSEDW/Y0dRYtvGdH3u9TZ
BLmCg8oIeUGkQH8/Fw14eE7A8i5dDHbtwXNLQm9WO+EYFFraUl9FwXpDbXGN
9NB3SvSIDnhTn4U4xNKPxhwAyFjs5ag/JY1QbIEwEueKgkS1M6YW2TLEtdCu
ra0pzIwmTrFp/EbfkxP/JkvIqs0BVkStcSnqhVLM+cRre5tjBgJ0H8loW9Z7
hDszZ6Ojg9mOvQdowLfjoJPLFjXCBdpQHUhmW1DoOb5Iy/Pf1urxJq39OfTc
PEWBqj+2MizXvBRVuKEmid+kL6XpDJtD4Frb0wHjvI9KpXICrg/AiCCWk/Yb
FyBDb0URaxpUtWWy7KBRBcFdaaloQKy9CJcYb17IC+4vKYQob7IPUHxYcOUj
L96aLdSkkPYv9eFciYg+lCv3UE7SewiXu/9VFBDMi9Ws3Hi+AN3Y64suEVPG
TU3ODNrIdkpBOA+CzULM14mCcbAALHczTuTPWsEVmZwS+dP/qJwO5P0qsUNp
vPXApRkhoL37037Ng5xJBFNqQfBtGtu0VVsyrTeLVxk4bGT2/CfMeqibx+5B
USMtGBzKM1mPl0I1sFCH8PBC7MQMFalt5uqvinGLBf4lrLhsQrChVFJxHYZT
uTZ9+iY7v+coiwtMdqsmKJPKPo7sbrU9M/th6Wm/bd7JU+Jokt0KdE0PZfL2
X0JSkbsCgnMXzkb2Boewg3maYYNB/19d7CTC0aJgCRif6kHQtxVlRI29eMAY
6Wt7og4u3/Wx5o5eXw0Fq3pb/m/ZftjPfm5pIM3X3HQbvXtVc640+lpY7hY1
+lua87h4cwmLUDri+rvSLxd1NrBkHYf8l2xgSwHPqbXHv1H2ZGw75+vLPwF0
tEDMNldCb3kTae233qbsOZyWZQB+gn3V3bGPCyX4Hce4XWX3Rk+bFtTJkNF9
FXo9MZzH62kti6BwJPvUBiaCnaFKyFJLabSG1CVR022IdYIBJ8SEpGItKXzC
aIN6tKzuPtTdQ9iFKag8rtqlbmPjCIGdceabvMJKGsGtZjjIVGE9zaia1ZTn
4QSe0lT1HcS4juA/cs4uJRdEP4CIOZIFlrZgic+y/mWq2agotr/MQVobf6wj
Q9+FSDjzVz+/OK/z+vdAkvrjXUFaD4lys3OaPZ9vjSz3ojcBm3eCAVGfCOO1
wEGkoF6DkCwjy13Q6nFCfm3C8wyjBzQ4SD90bEFG91MXTBeF1PoNWD/nWaXZ
ERDF8CIgcTs5EwOdsceUOdX2WU8ZXy7YkytmbxIi8k2ZOGZ2mXwn6rMU/7pC
jRsaBwZzNmuW/11R+2aRs23lPEIlpvs6OEJ825iQNy4t/ubkJaX/8kN+mndI
upyM16Y4ZIOR8gIuBLW+2TzqNNa6BW4RWyUnhZaS9DXVMNQcXEAZD71TnJW5
EETH0uEv+0dMBB/TZb/s7uObWvkJFFGzlcEIcJW5M8yE/lSmvkF4rA3uKTH8
zr85wO2m+WY341+Rw6O9OQhttpqvpYmsUP/w4JG6cFAH6JpxPD+KMa/9+NPc
31MvnPon3U04ABdppKDJjIExdGC0u4OX/xm+gHTyaOsyixEIVcdGJAdrvYnf
psk5xbODG0wQuSfm4Mg1xu4eJEsK9Jxu4Bmq6+4XwutOW0f2egesSPRWq0Rr
dKpzGbbbuOnh02DbmD9H1ZFo5GnlZIwyeBW3gNEfb1BesuvOnb1vbYikhmv0
Z3LYl6lMy63v3PSUbej7XSE4Q8rpt7sKFpXddguJJ7BhCdS8v2OOr0/lym8a
uBbGDXG9av6l4XLFgoyV88X83oDOl9w2aCxF+1QR43iCHuQ/NZ2cKZaRFukr
j+epSMflD2JXD+jIYLLlnmptKOs+kqzFPiR6KweSUL5Of14KdmY0DrlsJSE3
Zng+PGfxzd0CxMZr0pTqSaz74rdaO3R+uOFolmaYDJch1YzZDmiOrRHQua6P
0+FurFELb385fUSfEz46MFNgIFALrXpS69iwsgxYf6E6xItj7kc2YHkV+3xS
UoqrMrUf3B4jxlCxLyOUCN37QzCfjnHugRaF1OtVBOUDFJ/hPBD9p2gosqER
NYqitD1DxYtM/EGGtkfRniU2kUdlm8NT3LY56FaCchyt2UobVefSjgMXG7fF
Rq7HUzVxHkyIIMSIiQeVSUMQPRwQr9Bsn4mqzpALrUO55t8j/20aSGEMPESL
/aOpO7iSKAL+C+/LRhMHSp1WEuQPIGD4fMTl2A1hL5CS5MylGrYvCG/KJTFi
SHN2FBVjcDhOR/AWZsVoRfct/ME46k29SpGfeDzru+zhyB8fYQ4xDLq4iAxb
d6b1R+5gkk+11e2Ze+D4E6mryx+JQnFJgm5a88du7AuFYEkqwk2HUMe/5GTK
kmUvhoib4rXmgs+vXUgAVgnEVdwq25Vj8yG3cs7gZBklPvv86fS4HdRHYVdO
zRVaHLJQWOOB3A+VgAAeBGt0iqLUdI+y7wPI1I6m6WoUaSr7rTNEyROEcl+I
UAc9ZYHbUm2mXtLKSxFtrj3LIujI9RBAEXIruMDiaQzakV83badNiOsfk/pN
7g6TlQB/wZz500rNwIzNJ1ywyHHAbd9x5z1zSe6Ijv2XzyEa3w2Yvw/uhy1d
DjZeIw9x1xaqgqQH48Uo29WHNU179+Id0jsM3J4NBw9nhA5725Cw7cYGs5bo
BRTEyFV0CiXrAiVYQxEtgTBcemVsbENuLJP39YkYXKrHNzb7+qCvL0oP+bx1
OBUpb7aMIYlcR9N3XHjSbJkH2lcg/gVFEPHlnhMc2LjFx2Ti1RKKOpQ7IZEW
S5TWNcRus+Xm1tynEO4+YUCM9YfLTWVksgFwdxPQH6tYJgH8dFPyNUgTa5ZJ
BOtj3DJwbyIEFcSRYiYWtOKUPxg1tVm3B0aeHs0mFjFYcb7U9gedq07ed1ri
s/l3s/rt53y7hfhaI6uHoKb6ULPap41LpcuMLNta1gWzfCtqqT0zBSvWQPTp
v/qX6v3ZEcDdk+aj7QM9mEm4VASDfGBus/M1AzkMLrd5Y7PuBk8ZMZt2tzLm
HBMxsqrNtSkWApD2CU/s4Y4+JJVmNWwMNq2Tq+0XabtVO6ewXteoFKpoHrvd
tarNfyShImzWyKHV9zxcxy53qGITWpe3KzFEf5BLvAm6s1bX/mxxRFFiCFOI
Db8/uq5rd6UhHQyfr55xa/bFG/YVG4zNH26w87t3wrueIDi+KvJgmUYdA7bB
vebadVriatUPB5nWR3Ae3+rweTz8xgoEAEyt2OPUKg7gGc1D9EGcD3ypwtEg
veUgTZbD0hKlvdThl13xwIiFNEJAe3DChP2+7XpIZd6v3QPLNLt6DZ8DpwyZ
Vam0dtzR6ca4wzWcTvWZA86RhvFUFihmehzcvr3l+qX9URSLeHIc+8O/Th2g
6ileFP00V+b32eIszjPC6zK1djocvFGziyWdJE6FMgr5Vg0kVTDOr5PIroCN
M8KVGL08v5uLw0cgM+4FD075GVSBQ3It3/VRy1CwmZlNWnBcohj6wYNn6i9s
vxZEu8irOir03axgMxj5X0EhDVOnnVj4ag0VYft7o19GWh93zXmwgwKPVyYU
NNOf6o1JcFvLQbEKbgtmTFlQQxI7Nlz0nMQQ1dbUv5PCD7bHqHqIc8B/MCS7
95K93ra0o2KAMHEMgtDM0YOsbaSMNrid2J3T0XNzie+rSilMjxz/On0Pn6Jx
bPJp3J4BeHbenXGKBG9zYShzzgalKTrxjUhaytznYJB4MwmBv1+ihThSjpP1
oFcadCHGDe5IullwhegE0Jivfc4oLUQxXvmw1yf7XmiqpiJwBsRVr7po1kEo
BxGUEX8NhrOp866wee8wS3RVqz9eTVA2bQPjsLjrhPmFgVi5vsP32ElOdznp
7RP1OX0tWinkjUfxV4/MBpsHdXmZuIdVgXLHffgZ6+HRYEm6J11tOowTpDn1
WGLM/nwMOeTyCvsFbcejEo7PSYr2ok1VHUCMoU9EwC0B3SNWJv5+oCm32dgR
zdyYqO6KGJ0MJh8pL80COfW+lBT/u4KLzXzGddduraQUQfxgPl4VjFcfvdnq
nMqFsI6jqRJggilYbRu7ufdF+OONc4OtRjkEKXPFdAjbYvd1Zn4dMYJA0ILg
llnTNP2QnYPWLcHQp9bep8Tpuq+9OtAZ2eEE05wI8qYX4T2fYqbPpfRKtYKe
6+EFdoMZZVNwHJZ8UD1g29z+2OsjKm5eEwhW/0kUEuF8qj8BA7mnbaZJATe0
UoHPL7Q1gmphFjqSInVyxQ0DfySwdTjXn8ZA6a7FOHEq/92x2B+ijvfIB/6w
+J1UTzQzZOoUS4WNtHc87JlrgyPb1OxEZ+ega1Ny0eDzkZChrlx5yf9+mW1D
OaR4cwQPC5F2sApq5Yt+2tgpRP02VI2kFlGSgVevp68LctImVq6OBnzWegie
9rpvnK1ocSQ/JoeLwgKPwQq8Ph21ecC0BnLBm5wPCKBrxsQfKCxkvn8BvuTF
kOnRxRXBQTkeEVfPiO3TLvb0z/deSCka3ckZ5ccmRjM1yCQpyuUxreSLzJm7
NQiIReB1ZmX1PHU8hFtGqDNqNxc0tZoN2CE28MeKTyyvDIg90SSDR0iDIdT0
bTmYVfF8KWRLfuwxwdQFd7gaXRNo5DUuuf16ywI38ByVJFjk8ofJBYRGwuaQ
9w3WXL59/Mnk0L4Hgq5ogVxm77t/tXBl5foDcVZ8yKSxqzh55AoSQzrac04N
raJKm7dPLzTw4Bkrujsb28ebkUtPHksxSbQW5CQtFryN9vTNXxxTSzIasfdg
ZRTb+48q0hsFEG3KDd/QxJXoQibu5Wrv9LruDlgTZYpUckuj7rZ8HrAOaM43
7Ak/OkiUmAgHXLc/mTQDkv+5gHmWNTPTzrMBT168yh1XLdv4CaTxghXpzniN
cVrTFiax370gfBkVCKqwEsNoNbV/5weKG71Q75e3d1BfT0QBex1iZfyrf2cf
n2XjjvsEe4e8b0xoEc15Ul62Z34zdBdr6oggP71piTVjRjlKBsydMt96qnG4
igY5GHOiuVuQOeTOYFoC4OjzHkKJAcIVRRBi/N5qcdoIIaq7FekP5cakP5NI
lAwwwR6UZdQb/MV+jcAu46/TwJxWhCM4lByU3Pcx9rOOmOvl0wITeFNdUIQY
R5zj1Tjiglq5+/smtjC/2sskT4jvFSjiZwpOL2ynJ2zxT+zWRQbyj1CXOS1t
yPu/95XXx17z+BVr5uVZtIQd8537vAZ+yGJOA3B6PqOwFpWoVovalGTUs8bV
2tmcWKW2gMwc8UO4rPsbZQ8WS8Bn4EE17HpUEF/GUGandSP98tFGVxrj12RJ
UFSpmzH29uhzTEPeTtL+e7bRERNsS2U+5CLe7G5rU37Pd30FeP+IfsokiMqU
phXrxFYIcFKth7NU2SsXqTjbSx+G8x724LRFm05qnpiUrzYaMXpGX7OzdWsL
y14+vs7i34Inr1AjYhN8XonD9d/cbzVeu8CEoRF6mxx3W/w/XvJL7YAPV2rh
4nZHLmWef0bLvyQnZYqreBvukS46602LlRlOhkGHGesjHXM7p08PkAA0AxWe
VBpf1XQeOeKZSMCOmfZ3DzD9HfYDpr1mhFc8fs5gLNX2rq3PBEz2ssjTq41U
/eSt3hNszZX9JfBLQQKPiJpD1VV0B5CaWgZgIwsYBr3jEPxGAP7Uqc2Wtw74
nh93RjvY2BxPAughlMiNZW+D+taal/WvSE6MJxnj7Ozi8dybdU8zhW3XI9yo
lLVHM5z6lVxdwAD4fWHMi3F7o0268h1GEvPTGdUlCMrSyE37I7Zs5etW/f/5
IcwuDhf3t5HYLXSrxpZsIxjIxnZevVJkIT8WNC3tK8eez+LmJB7QGFXoUgIW
fnTa9cAMz0d5k+fPr08C/unHna/aS/k44urX7MOJlLUj6fjAjbJP1wMsECRk
iXhAUk29YG7hrI6UfrzsFhO2WSHXaL2icLWHKmhY+9ni1f8eTQ7ip6KGmt3o
xXN88tlC/Q3Ogn1uQpchsCwVbb64Ly18IiYTfsvlwVr1WQRLiielXgqt4myk
B6JSLFHbTO/8fBaNUBKt20+nmjNcwYdGeBxbvOu/PaU0xL/t+BmCGLh0XAY/
taIccddlJz+tq+pHb3ik/Ay/PGbLtChZRAn3at5efs/hFL60mS9tAU8vyjcw
c1dbKl0rbApl1OEnrQineBAbTrMp4IM4UKxKi27XQ0v7ZrGqpFsqzhikmvWr
jKSF1QfOjZECPzaPhei4Lrm83iZz4Zog6505e1/iXraBsnMJrJrJmSRIWirP
9kF15BhIdYxE2eCRNeIqtU4wllr0lTMKcQTyAc4neiQZSoT/We+dXY4IKw+P
EisMvNIrTN125vnqXjosfUXs1e3jTTQNyZaab627xVe6YArXup0kHhADfhkt
cO7aKsOZ1bvY8dv8jUo2+NLiKeAB3Bc4BI0EzCveeKgOlksnCmV5j34jTbem
AEYTULqJWucWVP6+tUu+4fGJQyqXHFq8TPAHaKoMJ4chKMeQGJc88wPFy6MY
NSiViDs48GAqzEOfZ7LgkdHY7A0aM7Y/OUW18W7FPt2FcKtrBw+nEHPw2TAQ
D4HP83z0ij0uK796jY+pwkBhZHGyx6iFeFcMU9rAJvhIY9Jw5A3bGa7GPv8p
rrc9VX1lPQBN3Yp1Xly2fqotaMCD0bV1z+EGayrwATCQYTl7zGoCurvKid5v
fCcFPqi+LSuPuPD0DfDD++ogxLNgeWErntxSqY7Jwlrewgj0YjNJ+tr6DQdj
0+BN5Ywqg+YiCFcgUgLfEW12NGOCKFz0s8sJSh/Z2J6Jkbly7CCNlVCUIRJ2
YWmIGjj3T9aYHKFufJSaZ6fxKr75f+aBwb/d1RwvjpfwiGiu5PMz1Yyt5Ev8
t2GgUa7Aq/FoMKCDem8+4xk0o1/b/gTk02JolW3La5CeHYp+TRn8E1itgj0h
gMUi8hE+nlqA+2ix1maCCtUUa4f6eMSW88ez18gOYg/uAKy2ICTM9caU2vGb
/7RWWM4/3DYl9AdKp3YrNhfTfUmO1oYRrgvvdHyCjU0nNsgEKWHFc/HnNz2v
wcF0orT8qCXXeuP2qPEJfIIpF4PQ0VFihDx+gVM42tD9tdXXJCdgnVdVDKt4
1GGQ1kxBY51/hpiK0V3/XHqKtcNTLfuZEOa+JrSuWJYprp0k90i0P147uPtc
f06eJZaz5ec8U07tcpB6+ObiqK2oY7cc+VuSHzn6lS+T3DLXNCFBeVyZhZCq
wJorncIMksGh5S3mlyDIkkX7kheMkBJC8s56qN4VHH3yxPYfefmVsUOgLe4F
UkDFXoF0DWhFpKOxyNho1UVXOsWv5Fqe++6yel1BCDobPwb0/8RjZUSt6TqZ
43lCGS50cf4FZqW+4SK1ibifTtyd9r23KaYWzAzGFo9nXzW5Wc0Tol2yiKX8
kGTMWM4rj6MZFqJINDqF6z8bkv3PAraPhHokafdAZjZYGScsAXsG8NlLQetk
FzXA006Ze3wxfHQ1W6lyDcLwlGmv4NmxvxAiMOfdNMsFsFMmXSqJBFGQATbo
7YXkiJEflpiA5SX7qY2UB+SgW7SBRa/pVLltNUnMuYfXsLS2zj5On9W69ACI
HeQWpK71/3Sejd+34yhJLgoPQjWkDk2JjZX/s/ZYYZxhA1S3bce3zbXD+IkE
tGmigjsucEgFVVKTQoPd+CzQnIskAEM+RrGQUPBylAJ5HyOHS8LO8rdq8BG4
9860ZEWhRQhu3kTOnvClf04pVmNCuMYrEdyyl/tbZyFUR5mutgNCbw0ADOaY
BquDDGizskqKZpyjUjNUJaZhygoZWDvr3waHtx7ZGjRlaSWC1I6mm7dB3Y0X
6RflsNnp+sm4ZzToiKTAy1UQWiakREsQx1W35f9utYXjYs2Paq+9kMWbe0mo
5m15lqQ+gwlr0+RN/WEZr0KSj9DRCAeqZ4ffYZ/JlJJ1KMyQipoeQWFOmjhk
mpLVIRrhEv9ptfYW9xUJinuDiYrfQ+qtqybuvR4alSB0CihYat2RPDMUo70S
lZGIpM58htQA5aS9dZybVJ6mn1dQC5TNqKKc8RP01ZFHPXKHE5Wbo/EWCBXl
EdI1bqT1HQnRJRkiwyFCp3mkcal2IvfJ2zjRr1qE73OOUEUstekrxoTcr6GD
7GJ65FATH0sr1hYDfK/rxJHtnk3cn6S+ti1oAJHtEN+mu1Osbk7zjyF5Dzz/
nDJ/GrGgmsIxoT09b8ScecaRXN3ZYdNZTyFBRRs47tn1Dw4atOozlMfwArLy
v6Q/fQ4gXL95ZxMImUd0cvNqGpAZIvjJynB8TY2f90G1fORrN5MEM0Bu4BUi
L8M3eblpKlBnQXFFZt4IcR4ShsVEVx6IDZE41URgNT8mX5IEvCnwsaszsyCo
KtNpE9Rt8S17mFe2SlrRuWiBh14RrRyPvfec/8uKySyY5FbfNuTR3NYOVvT3
2GtUfZAi4sw7JlPuqkUM5XgEGgXam9RoGjXT2NEBw2Wi1HINGmAiW2OVccjy
13s2w85dE7D8qkl4kKIsJKAAv3vQyuuwsiUkgQWzgjlxIwhE5B2gLVn5hD5B
gisQXuaq1uoPJmFji1W4mzEUdDDj7DOtEHBPMf3mvvxJ5B1YoOuz6zQD5pS1
Hz1kBI7kORojHZ2PbUQWOSvVdUGzkfWDz4qZ5kTSB/EUsmgO3OPCZlNeBvV8
EfaM/ARplIbOtfc9GmbCo4ucnEsacerR5na4HpIkvHMwFlMSlGkRY2b9y+st
EO4GrXIfduNb/2Hhq5RQywa1+Ms=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegBO2BNc2kmzb2laVLvZHowDgETeqZvZOuwnksHvMG72spvG5Uit48PG91T60a+Du9CpYuKAT4bLDGcvbWPKzeXkKPV5ZE1+kQcJ+7DJ6LynirJjLUjlm2rRXdKf5PC85rnTrzOrdYJqsvd4tosRGsUebaX9Vur0lP9GVjlC2jiWo4AkU5Glu5Dl5gaQ3jg55pNNKVUsofhaTthdIwboD/fiBf6xTFW9sSpnhwITrzwTssN88lqAAzcOeEdcp2DDM5bqo5sExmZwGdC9JtKzOtS73firFUn6e6vS62pGZwW0JXtDPJ/EDPq+RVMPsNF3r+GnAG/YJ1h5XNxfHFMjlRa7jwj8EqQsCoV00hy2rkfAhLT6Typt+U5lnAz7YTu7S7v8D6mIFRoL68lnGSTzo1gxlO2rvmml0t7/Qxea9cn1htMhPbkiEj/bG+fCGaAE2nbbyVdunDM4M+GnCY0QFP6z/pA+rcV1ZMZMbIreH42x39ODEAydCZVb7rMnETXCZUlFWXQekLW/L+8DjRkEeOuGOD45oV3AJ9CGjLNUH2Glx6MDqSaNO4rEzVZDqi3mvz3DEsILXzEwNT5y8wVqykR2rFWVSdnKMUQG5bmDq+RytVRqztWZ03gn5CRQy4kWDkcEVjD5c2TiEGGzzkBhPZsQYOSD6LOk7IhSoXoRrPJcX/KHNH769PqhKNRmCuGMkv1+4UJrjnWXbKcHxmH/wIilI5Bon93IoOqv1CMqvyENUFIHA2qFvnYy2NpeIj2/mSFmPg/x4mqOfuHqyIKaLxF"
`endif