// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uNcMqOtc9yOhO4pjYSFGZ91GaBKFKw8vEVESP8xKI010p4ihCX1Pn2s8dK3o
yZ2+kHJK9Dikx2DN0K0iEej2UP9buYBT3KC8Wi09O9sLPlN3it3q9rFtExJd
e0sL8PoW0LxQghzfJLZmzj3P1L7xq2wSyJr5fec8tD/IPnaKSMUuFqRNNB0U
0OvtdkQgeW8goPdJHiKbdPhBNGsmRcxfvaENTDd+kh1qjoxw/Cur579PvaJ4
DyVDmvRi0eSIBs5ZjWQhBQavM2Tx+VGI8baY8AXyn9/H1OSQO8XDIs/QDTDK
vlYs6IauIaXHdyW3f00n9aLHwveyb9PgNcgcPUZmIA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KJkoZM3Q4S/cVYbCpkT66eYCgeNyQJBm0tmhW/JHSwc3XbQIVQ8iBCGKq4iQ
rBSKVX1Sk348m2/rCC6AfYTpnOnd8ztKxG5M493J1biGMWckGOdh60vGBi/9
pFtWTgzKYsZ6+wYEsfVYqAqLgD+I7ga/J61o6VpRkBSMyrGhH0JZyK9vW54u
ucC380OOPxFcTA0R6o3btIUymZ+rxmQcrOSbadrKWXL0FMa2MmXDU/dzSS4Z
QKuL0tZl39wv2xbbT/BfhwzPgcWKeVeo4MWjKogw7hpJECtT1Rkdn60oTbYW
sWLGxufJ1WaXSoONVb9I0LNkaknZST4frL8R+xYCzQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
roYAoS5pab7tXzGEwlmojYhQ1kKOjHJgrKxZy1xrkeqjk1jpsBINIkUIHk1R
JCLesIHfYxCzzwG4X62Jjk2JUnzseZ9/aBH4XKzAwb80YsBadKjJPkwoZ1KH
GzSG1AZVd9BRiKGqLNETEt6DohpAGx/nxfLZQhlJL+T+xdbOCRDPA3FASdYJ
qy1hv9atmW2rnfnZm+NT4hZdmg5kjGUOaHixrr6mPB8aBX/vSmh9d7DQe+Zx
dXuwhQEqS38ncskASnuz380/AhgkUiKmZXMomXiVSHhITr8DZ1f6SEn5z7Ro
IuDSNJAirFwIxOSFgpLOmemSQL/NPiTl6oQ3l/GhqA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HzEwrYjZMGTzPhvjDuIwddolDI1jdZePSwMY4TCipL9nqNDXfFgbh3Ha97Tc
Wx7H9Z4NOuqxyOX/f7Ycpm74NiGVwvCUITv3pCL4RgPc19BpoGKjpMlt4Rsr
cyVQuy55105J3VH1ldoggiYxEeyBIySnP4Z3qzz0DfTQhSDwpaQh0g/b3r8V
TNu/dtjwoIKHK+Myp5ZIivVCZjvAujqjGus+k4fCw/yTL2mGKw0Auh0ULH5g
es+F7TBtQeLQuxQbQ+TGyTiuvTnnFRHtXgQgwuHJp0HXh/ZhbDs9NKquYwV+
fIN3bhD9sQruFCMzToZVM/z+jU4qcWkauj7v/P1cHw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZAkZip9ZCCIpcZDldED+hbEYM/ilJoAWoBk/7OIyjg9yHFynw/ecjVLnwRjW
i/8mLHt4oBAKd4cQuHfRI/U1OhJiKOjzhh+epA28zK4Z+l/yePg1AtiV3CRU
vQv232ciHzSqm+JJy+y53KPqWfwLUPlCDFQ9Ftd8VrAZv5uXGno=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KBJy3Oh5V24oNrQsu5hgyTKRwv4N3ya45FKFt7Gw1TZocUsfdVTIRSy1/lG6
yhoZfgfh3H3QE8Rm8NU6kDKDtPCaw92144yD2EFO+Mqsek+uBiuAKqX8P9y6
Sny60rpczzS9xhyPmnnx6t+7cKyFUTZc/otdGgfOEDB0HtxRBZfkdUku7GAn
lxraph7GVKSRtUQU81VPZ//HqLbrP4Ka+4XQc674qQhZVEccUZYGNDZB7q4j
JtWKvlGV/5/8pSrkNBTG5OfetU2aZGXXE7sfO82K8PAxV5AQkLFkkzHFSnRk
39g5lI/dho4zy0Rba0ckKuyC6EwEeOSoyPjQN1oo7BwPnv/fQ/u+RQLL2CMy
+NWih+o14qgrSSYxzpahs1qC5s4o0eu967q/X9uQQfxxX0orpR/EPpuSBRCG
xp6xWZcsT7X/OQQVA6l8io5WOB6/dEQrynusOHT3XHP2m3SwQ7stBjv293C5
WfA3dXWu4Oq2fRE6ruQzTS8aGy+v5SX6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TthNfdsqoU60Tll6Fma4LbbW7K45gSz4RogZQuPzm+XXTTWuLWN8MpK6X8/s
Xvrn1IhVgYdi2xevbE950wybWiqoqvRA0eh8b11+yQWgzRTQnTw3qe4oQ6pr
7PgNPjekdBTseC1YLZgZT94hqasV/h8UKY1c4aZp0pRZ44cmvT0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RiT1gZbMJOo0AfpdAxNckiEbVDtdJbGHd2sm+GgCG8qK4Fcz3iFVq+Atqk0h
2qUyVr5csQ0ZnisVSsoCZwfJ0TEl88wMOgBjfwsAS7R/WALhqPXa/95WZF6t
YCCcUQsoXAa+B/UFDD5x80aGGTbk3XnS9h1et5anWdGnIGDM7kY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9392)
`pragma protect data_block
jGGJx+zKRf+Sk26boz44VfrjgFECoh5qTCzBSfXEuouXyUYlhBoSXI6dMUtl
e6vXUx/6hkdeYFRTMpKikWqsBTDKKvlS7WrEb3cFYfzU+rEjnw69llpxEbIV
FKYfhnmSz3lUtiHXX7tlcXUGpVX1iwAuj6QNFyaTrRhPjER3GcdbWCSyMW8u
PUT5e1Z22MhPX5OQMh8fvIjzwbSjwCOQsCw0jC5jy2qHhZVy7qZJRCie3UZz
7HEkTT3pgPGNWQYzENR+gXKG4Q4pXEnwJ3cqb9SGTOeK3egvHwcpjfDCYxk+
BRsf21kblyvCwtvQoLC5FPEUFGPcgR7vfQrDRZ7PfSebPBxRcyhMynxj8Em5
mTHnBLvOBw3l6GGsiLW0TNHpH+YwV4kdzjQg4Slv4u2CSZasDO+LoVvpxRmA
MM0nNIag4YXTUCVtlB3AteXdQzsNg9In+k2CL3R3NJUgiXfLHWxyrEgjmcc9
aJEjBe4QyM/pAqFISJ2Gt+bEfwwgpmq9zYPK1z01uX1hon89gGTywjMxFj3y
XW4qaRDFabMd7MBxPZECRzL09EJ+CifydXz3iakhlT2r7cRM+ILkVr2kC4EE
4rblVmyvzSwUzNo+Ey/G+dxDUQn9lfrZzlb+gHKDsUruMDv4HfJ8ipFGBynk
SO3Hq/kfeHgDMCl+ilqXMR5FGJTsjRa00ydVEYUVrWOAbJ9R2suH7aUlBlfg
7FurpSx27z26M1BOD79ck8SuKPf5Ul2ywQ6cuG173Dj0mkI3LyHl3b7etiF/
H7lURD1VBhHTfZpFW25gvPAMnGwrc7TaMSBCI2st5SzgwBaRdyctb02q0dkq
nnuGUpD92N91CxpQHlbiZVEAyLf6TvTrco9NBScyS03cVZFiqQrN28a4ksty
CViZ5+ylNZ1aHUj5m4Wrw07LLASAoWcsv3CqoQRRj7izzJWF9h43CvuS0mXd
a6U1TPjSp8DFHmTET/Uhrmq7O03OyksHPUWVVy30s0pu02qUyGaUbQVavBMp
asLVQ4kzQEUYkQS31UMm2icgoesTL/XinJlhLTqLlz+xzYhvWt/ZE5+TShdT
yDGmnuyHOyFUogFSQYDHyRazXvL+q16eKbZOHCoFot5g6sou/zhTezgsoV0i
86DuNJYI6L0XwLw8tedtB67/I9z7Bref2GEHhLefclvbdbXoj5VYOdbRQq4b
tS1qcgiVNf9CaapWMHl/qGhEZi5N9ZTWrKY1w5OyBdaH/xwHrSH3H7q10yMm
ai/PyZo/pPsuh72neLSjjV0ekiwoLO16ZsTsqCNrehdgcxLnVF7mrRSZL1po
lKgf8ikVRriJU4jEPgd06Hyi+NkiVJ6+owXmyzM2owGYPBz+D2xclMdM6mYA
+4moR8Lg7NsidN3VdUj11BIBNdKO62/wYGoKh/BdLUX0DevOvbPBie6bsQ+E
p46Pf0PurUfJVn62n/EpksHECmr7amKInwt/pFxxtDw0bWwQOwkM9+2hiIma
pfmS+neiWZfr6/xY9KTmQJPhi09CcqSLj/ty4huC2MwtVe8x4xAtUNMP/i+s
7q2U3VlNSsd3u8ySBa4M+5LOs8bKIDWGRdOYbqu4c2sYRxlhEPT8KbQ+gbcE
Bs0/T2/Bk2RVHema92RN4PeNEwlWifvLOMpw/ZCGEqAHQtLsaqM/uiXPdaHn
HHXeL/45o+g/sfaFNK3PWcLnJF6pFQhAm+633lnMRBTnJwEl2Cq3rHOMirK0
hen2MUEkbC+CYnFQq+eRpGRTpzq33D545PkhGHGJ+82sb17gG8Xnz6TV7Pdv
ezSguHnf537L/tT1DsNt6FFSFGzH8Fhm27mPYwCXehddWHeMUC91BvaJMD3Z
MzL40XJdZ1tMHYbsrwn/2nmmXwpcox+YrFD9svLyBgxIOivnWxF7a6kD7fqy
nQMEnE4qfobhpU7AUCdZDf2ESCD220zPQ3/l78W0/tNXpUY7SeBAag5PKrc4
qvlWx30q+qwOInobJiaytkzK6X+3qqza40dFeqOE9h8Hw+7S48LDUyc1+AwP
U00d9TKKhgK46ZyN2ZZ/Od1b0x9qIBkTf+Xdk7yEJRPQbmPirOJfi88y3L19
NBNQoP3sKLG3e+SKVIGub5uyRXSU4mNLmC+31DoTT+Tm/d1OOX0IarG6uB4m
fRUN2W/apt75R8pOnJMMGiHPIXZYw3NqRVO17xtCXm4pWNuJXXqkwOBlKOjp
RAwRlUcedKDcHHl0qzlwnaM4emfSkhNk5Xy+sVKiHdKMGW0xvCzahjlmXg2J
UzHzSokRHGTMthIysmY002pIEI50s7an10NJ/A88JNuPatcwRj3ZH6c4av79
WqaW3HtgjITSgf33vZoNwPa+pHM0D7wLcplC4jPkFc/4W66HG/4onLnic3Ci
DNSnmKwUrtFrl2p5qhFlQ3gJVbDuCJCe+M/YX0mNFZQ7TVzydsIUET+9bgD2
yfOeiVjmgC6ltnUo9utbYo3Xn5Eb23jDMXAvZa9vKSaSZ9QWhOpuYaJNFMUK
1u3wSTL7d8xbBckb8HOCe5Zh2bN+HoEem631TgObBu1A5kSbZ3c9kKKoiZ2w
r9B6P8F6Gn9bOkZh38V7qjXpzEAix2O+ScyTqGLURIFgqIucRlm4EDJuom74
9A5RYKVi1N3Ha5F1sbcZm3PxNv0us5Uy+47YpuaM5fetkyl2Fws55Dlsbd5r
PaCL/t0vCysqKfFtZNmA2gOWqE8HYD81cc0GrUhfzFiPPiFyZX2M7QOW002n
QorBUu6mFturaEMPyeiBhSeYMzmy14hsCZX4rDc7fYJJr76Jn8fk/6LsTYV0
WvDxUc8+Tm5CyjK8TIk30e+vR65VH5YbNNbp2KWywVAZYXU+4qCS9xMAZKGS
sSFyTYb7OoypFM6Mfnzr3amrf9jGFSI1W/ejzsJf53fcRBkDuxgkZAd7U4AT
C9CfCvVw0j28jMTeMkxA+nNP0wk6pBvtBv/1H4mcjBQ6ra/aXkCK2Y67mNbD
VzyzVx8Ho72IdPfQGbv5AwogNOmipaeZ3EOq60BF9Dyv14PidHL4PLp7WVF1
ekrY37VNkekQzESJc6fIvYX6XpJSVb+NoHvfWwvqjbb04lwKbturqhksh78j
8H8StR/XOA4Ey6Kf4nLO3aDVI9383XiSdCDY34n8goz+PeEF7sr5ftSDobgf
QPizRcE1kaV4NKz6I20r1ARZFgcNVW8rhIKx4yHa50x0WfkMURM+vZo01ypA
p5Td60IsacZAkdmPwWXgDvedA/mzppAMAkNco7BE/7MRYdtPFWYQOsxwiZTt
fyocXL2E4qm8atWxSa1w7DqJ1SH9vX/WDPHCOwQTjDK0N9sRIRO0jZMeSyEx
QZ3ys/cTl5lTs5SB8Ak65jlyybAqqDF2C8uuPYvy3I9BykrI3YvPijyFC/a3
+5m6sDinmCLa1RvYHVubEVZYRJBZwwkOJJ4qBjjqbUMbn7l8qOJ4BBjfmAeu
Pvfyf6/6Usb8BrTFMY8OvMxHc0E4CZ2Qxe7FMePe4/o25BfiZDCQ9fKZ0qnB
QQ8OK/e8j1Vhf82L8iu6/Sl/aQ6Udgf9HbpOq32KBHsAkrPjDDY5Syb9FFVm
Xx9Xl8PQsSFOJtF45DVaf6DT6ipCof5/0i6xpIS24LTsBAjpJYMEF2QDSySb
SrcOFnFe6W9RMfHH2ZVQfuACVAAArM7ZB+/gavTqpty89PvG6Gm3Zn2dm+eQ
wlC9Y/dYBsTFqUwg04J8dvmc4mjbNo+LZ2/cIpuIxVMwANxaHcK0OTTxlZFt
eShkZYyYwuSz0CuIgyEjJxb7xapMCtwsgt9DDuqBLlB/UzoBKfgqq4NgjGt0
G23KYksMh/9mFpR3Lj/PrpEK29iMCmZf/Cpq5aaDWaDknhKIegEFIg3whhOU
bVxiKck+Pxle39R7Gzcv5+LgcCCUH3OCQVJI7NdkCYX9v0IOk0eJw2L1dxha
3Q6H+NVb0e2M/S99oD6w4X5Fpk/Zpvc38VJjKsch/2AoNTHCbuJHL5DIERd+
42moZEhijONH89oK2azOlagBN8eE/AGjSPnNbL5ZCxzRNv/v3DQHngIVJR7z
f9hNYMPzcJyfv0VLykLGrxRZIOUG/sHmxf4vLnmFXbxH0Zmt9e4qHiFIj1LO
HcxUqEx6AT1ejvJxpTRVhM/dyOeUMglxvf6tbt/TZk+SvsJbLpNt+Hfw+C2U
56NZos8Y4mHQDub5DVtKTPMrY/GBNJiCc4o2OwiG0G+/CgNmNVVzDe5E9M2E
RNdZ81e7P8zUxNQsxV/vbet4a8FFyYU0i4PUj/OFRulxHnL2lm0vnOFOslDd
U//KayLoub9yq+057Tbj52gD0DfvBINsxdYkCUpXwZ3kE2AaFy0UcoBMB7sA
lL4TGZKJaNaagkAuEPHlORplo/jSgYZEbITiySaxXFzBOOFf2iSzW4Lfz0rk
tcjx4yF1f6Sy7fjqaSNeuR7qBOqvi+DNiz5d3lWNtCZBHZurtwb+rg+ydOBN
afORH7FqqAKaSEo0z/HCSf2aP57FAB+PMJJT5KQakJ0vI+8kakP5Jc/prBzg
w5NBVbW5wOh/uuBJCN0o/Ql/JSngbsRQvFJ0yMbf1LWJvbluGQjEYTcpBJQn
dPZCiwZSlz50buncBpQufkaYxUVRBH0u4Krfh23+oxbTFtdDscWHRtMPOlR+
K52q6pnTQYaencACe8oZNjpZzHcy1hV0zc9GZbY/WjVTi07raewDhE39XVoe
sYNMuD93PCE/qxLAN7S9Iij9w4NROp6uKqfFtga3DYIOq1MD1znjtFdgKBhU
T7lRBd1vEQzooOBu4feTBBl+gRKx9zUnYf18qRNTdZ7iYNpGKSkVp4yGGTFh
2gCDiOmoHCH7x5PpxgxNQh+kcfw/BMAcOw7nSeKK3wVn5ZFXoiVxjSmKmRz7
+KrMkrknEsoGBZ8Icw5YZv63cAwb+LxcQuFD3ZxxbhFT4ugehUeigTpD0WrM
o0XDQeQmLjMyRH2m4/wbGRRT5FYOqzV8kiGtCoraYunYnr7h/CqMh7k46Xw6
Cmh4ffQ+ya1OUnB2RkH7IG57JdJ9XBxq4W1S+HN476p7bIVhoc1t10XFPTkx
LBNKULLqEng+F+39gYc0LJ9zyGF+9xOQxqbMJZfonX9u5cnBNlAc5+A617VU
NSjKkWHwz3jZ6epr0K86sXSd0cbPwPomZaFjg2TLBxS5IHazwJzx1qDbkd25
1k/2EvYxc3Dh/RNVYoRba67qL6o4yW9pSdmBIMiKQdPm0F4pDNWOE698z33O
rCibNvl1YcFnqCUm/RPm3CJguznrntvm7bVCL4ouIjhiSuDoawrj5KQz1Tbe
EhRdOt2vOc5S2v9jbNf+oo1ytW+/WA48Mf50UQjIlkagpSRoM/AKlHfe16J+
NqvefHu28+r5ACuz/m8KfOEA4EbelDgksAHGIt0z5pD2nkgP/CKAH4uJ77UD
WqwIRDsUo5Ksi9bM9X+7w6GjfmTodHxDRPAIAxdDfItdo/fhuNbU5337lKoU
WNO/UoiL9N0UWKVTAcUvTmb8QO2cRhnTJEJ+ZUANO7tIEJ7/+czsFV6Uhz5Y
tDegZ33HQj8JDBKS+oXFLZ1Quhxmc/NzwGcmn+liIaDVGAN03veuL1SzIV05
nKFxaTLu6OTlwNvuiHL1gXQ/Jn9+7te564QYCmsDFAj1qeJdqZ0/7FVeaHCy
39R9z7xiKIdPbJYyU1YVQQ9DdN7S6/ADK30AYMux5keDgcrLkL2LhdARHQma
W7VPT0+OclkA5SaTEm9HVizdSK+7TbSaMoKFwnnPoUH9a4+unyMkEg6TeU5t
9Mqe1i6gHqIkIHFo4ttL2RqIi7FhwCsHvv0hsVTMIC3OoFy8QfHwUROK5HrS
rjPez+lQmsYODG/cflAQH0IROGSFKjlhCLl/3fmXe8XN2ApO2RyGI8JDHKpt
D7Ct+C5WAKDP+cXf21K8iB4GIHEt1vd6g4G5EceJfI969z24oTPtZnwHgfP5
B+kyNpOGpcdkZp8qfNl8ofdXFUr9OgiRQS0foGe2c8OU1RhinTAFtEcuY8xn
qgXiqnKAQESHErQbMxpgfhe2/B1pQQroGFtWu8WJ/5mE2QQrK9hnEWNyLsb3
pJ0a8HtRDJZN/p39ZppJW5d7d8L9Nz8l+tzZavSmUvbiRS0DYQRZD5mtTAma
tn7LzsFoGQat6TRtZuGIIh8GZLVCn3qohE2oea3gfZ2vX/7Ii+DERQvRl/q6
ZADr0mWVvKxw0pJFMnUc3B8JiczP7QwSq9GweCfvKXKvBq0QG0U+1weLSQJZ
2bFo7XTs7UtYstd+v8el34gEsqbih11f9CchEro8HQkPsRhn+H2hzTkXDxzi
kSzgZAs7eiJaon+oyssFWHWysdJ0OXy7wpNB4WKAYZuC60onafPcTHGX2sfM
lkHYJ0SaLUrVrrPivGAroA9hWo2fpYSe5msC+/0umiXyNLDOD9hWYHuX514j
hlPiKj133D2X/E3rsqKb6l4ySAYQcUHEhMUisc/5GYhlHopAoHZ/FBau1J9G
qgh3L6ubC0tu6d2WTkYq1t4bdEOgvvfcTiuRVGQciSjnno8Jh02f2xeItWw9
YN1/lShB7KaBSsnVI6uWSIf3XEJcvraie7CQKQ9FjaD1Bv8IIgekdcwMAXmW
+Dju4cAOSVIXB/mslMBWmoMtvY3l6P6iMGtFByiw6r4GBig62zAbuoIyfpmv
nhggKpx21HYH9Q0yz+lmqXeItCCTrbHodUUNZVxK5IrI+1imgXtSmaOv+513
KetKCdrmklPr/OdQEP53Qd+TjRjay+uHGJIEY2TVFRihG7lqqS2a+NOHwSbM
H/gqc84VHK1zIsQm/Zr7x+5vJos9I3crDQHHvYiaNwUdCECcY6eslXq966pX
blR2waOEVonrY8IWjgfil6YDnMV1PDPR+0jfolNISWIMeZKOew9DgBHF+Jw7
K4zSMOans9YULw0gwmFZtCwAXprXkEAPlllGesfdGO++8z/wy7qAQwmyl0Ax
4LbAv09BBl69MuRqy0xQ9bsFdw0iGXZkb1iQ+tPxDFWRU1UhbqmMIhJrV28O
I2IYf27BPpq1P84USDS5+HhUsW5suYjyAz8/roej0anJi0CzR6V/xe4ITvx7
OwweOn1ccH9FQqQrGyMv4q2a34ZR08ke2YLmD3MeANBFnYxZVC9ab0a4cMWr
Po1e7gefXmz4MKulC/NR7hzJtrXU9iuFBDAihYZyZendKJNO1QW5fCXEOEff
efylFJAFvKkbYGEd3WW4u+KI5k/YJdor0SUIaCnthJtkjciU7jrAkOIuWEmX
5wU0vgGdlYV9dknxjJgBRKpkWYosRVG9J7XDf9HSSR6LpbzQUWL4RyG2d2JC
+nktihTZRc2ScNUXWjz8My1jV4J9836Dy3gpf3xerts0Aqgep0cXRNC9ky0I
EodUR2PCjdoAQOyNowRT30O9VXi5ecyg9Ilp2uc//hafQAnEtv3NWSBOxOtW
0YT37mr3+fItJns1NDekfRSY9AQ9c19tMxhA0gkEOXfIFkaWEfMv/UO8naMv
72pQXSmUblnECaG1YFXsFkQxcyE9xHVoovtfP43C9zBXoa1MnGjHkcFeIdPf
95wNJdGN/ulSFdzGka0yun6pTT6p+XmPd+hBz6wQuuivCQEO4TqRaASN0GZI
2ToNKHOHlAq1cezaFD5IHW+oGrvRgL8ai2DmcbgsGEYcmKK22E+X9Vxmbhvn
s4W3Cra1UTpmwfR0zq8IB1u+vmo5uWHS9QF6neNu73aa/q9Rd8ZuVMVRj08+
7cbhXWyuAmLFLbYy+qGpRz5jjqkQArlTw8ow6AVg2QEdBzg84wlYF0mUNoEV
zTGJLZ4YFd3pdFTznRADGjZN/DgWxnJGnmpIUl++YA0tctdDbVB1MqR4ZY28
sNJL3aT5UQaV5bOAP43Cr60FYZ9+E88A6OfCPLt3qD98Gm0DT/2wvGD4zgh9
egCQh3r5nkp/DOYLNMnYGewPjR6iZCfxIzPVWP9Go6TwpQL1dKona2FgoN9O
1gAtxmSdEie4uiHFpIsfIB8FvoEoQve/wb0YyfqxSlJjjUIEDA1emejr5teB
ikKMwvGjz3seuxHvXP/w0zWyVADFuhv6ILEuV3zymsbxKMIE4IVhInMHG0FE
Bh1YUt2TmI5yLnOK4V5/gTUFZzbivUyDtSd+XF+xOAZDKtgi+8Pbj2mamXMo
iAVSJaefvDZwf43PCyp5clIfjjKpDY4Ut8DSjHI2+mEot1b4Eo0+9gIL+RYE
kPfx8UrMfV7w5xlgSVyU5eMmna0L0+uLV6gGk49Bmuzopq7lK3QIqcysp5cQ
IOMUdTlwnYgL6LjgvO7tgj8dM1ebUBTxFE/0I5HCXFG9b77M0DGFfmtpmGTf
eeZbWelZsllhNS2f4okwwM+wupTKtzx3TwaO8SABgp+RY1ntYnzcBQQ5M1Ro
0KXVAIWpZfdeFLeQIDTbEhW7GMvz2Y/p3xn6KCxr67F2MtmV+qY1U0ZzhnjL
UmD4yhsJ5OxlbZHqz5YGyo2rK2ovipNZbO1+9ChvT/tBvKlxo94a6qYaJk1f
G16UauuJj+8rPHN3atTucaHL71TcRGd/07ZlDq1F/6TFwlZr4KPpA6iY7/QU
ILE5zrTX3MNFIeyA8tlh5KWGN/WhF6fCg9kQyh3iEp678QV15TxVLHVUzmXL
oQ7pP4pXcROF3DVWrY+YsFdDaVx74PmtX7sO6YtgcDY2XYNyZztgbQgIaWug
sLMVMkKRr3lBK3WKMh3wPvL3x3mFMqQQ6l1zd5JWq4n4SDO8LUKq1l80Atyy
/cdI5RONZkJIoDJbUAdp+saYwv2zdM3rvFBQFBotP3F6zvaBihZNl5EogFqz
1Kv78HkXWoX9VJLo+GtPyly8EYusn00lvqqbm+KH9WWUJr1uO8rcVOTq3o3P
OYr7YQihVCgJUmd/KU5AonmiEjRbskZ5Lte1/9+juwNbZrWbJP5piyC2iez9
WMPfKWcQUoU21bAi9XE/pzeTRzBSbWdpJTVsIg3DQ8na/mNLR4fdX9qLTsRn
4VcjZYuF3QD7LlCKFs2bJ7TxTtHTYkNYUUwGcbMPJolvLm3jt3Hg1LZd8X/N
faOnz6PeAQxhXb2hM5XG0YGSMpJMSVRZic9UPwSi9UESGGweodOhpOuXlaU3
2oo/iuG76Q861nvP3GwsRBMJ0Rz84cR5Lle2BGayem/bpdh9O7IPkyc/6J+H
vFFScMMh2G/Dgw5aGkoaMwhr5rvNUi7dOsvssDJi8Rf5XzidKyw9Wr0Aprcy
wTMs+Kn7y4GhuQD2V6qABIo5iFgKdszUfy4PSeUJ9clJZ+B6KjhWJ8N1TOp8
vrzILC9Abz80u84Xkmn1u6ag0BUWN8R43CxTF2OPKhmmannq3E5mxzJMqnZZ
u5863LdWEFIuqSGqG7jpkQzH3CHDMLPEfddIf+XfIkeMNo/11yjQr38ouE/w
gKl80CuqCnP8H6WX2gehd09nsFhujQsviLfvdv1bqVIGH4hznRHmeRzOdUPO
SVwwefGabQXL3d+VhrWx112ZgMw+fmhrkPboM/QWCwZgU7Vp+Bf86trO9njQ
Pc9GUQgKGBU4tC+uhFBvqqQWPwttNYSIM7xr2txOWLX2YCXz3uu1wxZASkTH
UVeuL9Pol3BLmaxHZZTdqWSEKO1V9cvDHGFEBxdAjWRbL8jRGg3QPUi0gsMB
zK02iuLDoiE72R//s7apv60lf3Ar46kke0UdwFmX23cwmaTXbUYysYCJxs30
cxWQeueG2pkgTwyC1bkfVkDSsDWeThpmsckORXLxj7g/K5v71fbsBCIaV/vT
yn+wgszpCVS5sysiERxMKjUb44uWQ9UWK2O6sMU2fAQ9mpzy8a+Zm//mcacP
WINRlYsRDRzruae25WcKcvAhUwTTfHuRR3XBl3ntM3cA2nC8UMoqmE2Sfez8
mz6K/ti7O8NeSyPt876aKs7Uj6hHogjbkQTLEMIgjohzoLVWjsjUn3fOYyUU
6VabvOwWRUXxnD4+gWw8T3J2lw+9We99QFlAAvCdTRIt4VFxXToncDqaaCv1
3aaIUd471AGvMJZOyWBowa+NXXsjJDnXflJyipDYjZ2JkKJxvNOLX185e9cX
IBIhPYBUt2B3INmpo64qZlxK9AqBDuIfjmTHtiH9gXyey8OJ61M6c18tL+IE
TFAbHjCj3Ojm47nL289PCH0zPokrnS5QVG8+G8UV7NPkaw8mtEcr7jZ3CgCL
Z9p+/ZBO/LDmNy/ISTFZCvc4HCYBqNhjAWnNZIAyQNZNFM05XCYbglZwi+yb
MRIucKiGruNa14rfPa0jJgaQcaNd6XVlqTCffDRVlA/Jjn/45b9pw0zlrQDl
NYSJIM0EOvcZ3ziCJIN9rJFYfJb0rrKhqO0G9MTjA92DA9sq2UY/A8TKx2Nv
43jDxJjMmNHsyS4OAcYAzS6rT8U7LLMczzPiY/EqBLpo/KQzjfG/IPIMHs/S
mIu/q3htcEJv8bKQ1N4XRt9r8ta1waflzicVXE07j46ZvNjPiygtXuKj56XM
PDC1312kYxlvSKhsxiXP6wJFxjNRbBWvc7ffJjGAE5KGdthsUvYmNfzht36E
DBDA9iSrki1HxXtLRRC1ol4s7Pp9zufRIqQB1PRNIhV8hUxBJ80UUK9orB4C
ZTA9M3WiCNyprqBSV8fIT5tXdsK8DdLRFYGrHJuoDorewUjClzKefRyNJBwk
8aPviGrehhR7o5ernOGOA455eDSIehyoWwsBfD7deNDdlqcyxPchZT/VZ0rx
8LTpTvwOHcGJMK4MQRXmsMvvs/Bu/YPdoju5W8B/3hDmC0Mstrsx4snqoV73
a33Ue8khYfnI+fTt5qEyOzKdUw1W3FD6SMdxzUgUXdVWVBFWgDTEfvoqL4SV
0O5cxXl176TYem++JUhlx6k8UDKtVF5iRUW05LbVfmWFuHDJA6Ole8b7gxee
OGE9TORdhjnVnay4RMMIhdtArDIesUXtOosNrDl6dybmqf3B4/ycfA1p1Cka
ztvqz/mRg0g2MsadPEjDnG6VuIipx5lV8VRViLfSgBk4pBaTw+fzY/5QOK+b
6bd0/cpuf+Est8vcH6mVHHrQAJT6AFtcFQOr43v63rijhU4gocsfv9G10f3r
QmDZ5E8PU5DvvsNqA47v0ECGIb1d1AhAxLGFn9GXJCBrvlomOTeIvn4+7Cvb
9SGd90pPRlyIvcQPM8zL7GVPtSBdNIIuIeecfKIyyXgbxepXIugnqpnXUn+b
ZAMNMS0J9cAVe4E5x4HDWrAaFG56eMykaQt4i2yXnUqlApJlTD4CmFJ2oM45
MbYKskzMCGp+1aPKdbO2arjVal6P11nfbmQEVA5dqtb9C9fBJJAbocTXHx+2
uQLVVQPR/ZEgpFrauYOAS0IUncgizc3KvnJaapJ0RXONzEU1DoL2ra0GOdRb
EPqBp964+HUJRZ8fU3ckjbOA408495nFW9hdKwFodwh3dwxEllgQXkXYRmOB
xNsswiai+6U/Mi0VLyb2E/+AEx5UkHi7o0bSsuI3Rb1NDozJjSiwYmtdPL2f
0UhdlkIRcONpkIjwjb/LPo/cKBtCIgxeSEkSS985CpF0U3ad7bsrna0trrf9
MYAT8FJBBI51tuTCqlvJI5yJNDujQq2KEz+DM/QiWFtjvXGdfoKkvy0eG34S
RvK704dS28xZ3QbqUkvSK42PGd4yiqkbzNl+J80y0a30FuHNrddI8OGlFdRz
3rGWwZuLndux6l2iveOlL01CpzfPomhUUlW4hGxRic64wAZfauiHINxtal6I
ApG1kUSN6UiSbeTCRjed8yRGwoadoSTUUMUBQjjxzDDsH1YYa+ZQEMKgM0it
dt/prRasSSvHYsrpgtDY8owFP1QZa3H2ZxjWeAOKLHADVm+IfEYVA7e853jn
lo2tmvd6gGZSJh8BESgBfplsS2b4WynJ9P8IQHkgH293JeO7J/UDSuubRWXw
m0ikD0N9mk8+5b6wXgLMfWiV4DgTJRWgCwCG00kQ+sGHF9T58HVyaCGmxtWd
O5Y5R9Ez1Fh0NvYVqJQTahssGNhvSZAXSj8EKci+6nG3myq+m9RxpJG3RImc
W7yp5NkvpW+kzGSPwhmTk/4WVQG7VOfm7OGMqRXTPRjDs7p9s4rtAGyrysZ4
zALrHvRNOAnDKdAd1kM/cvPZiwQ/vjD49jpHVfiTTp/Rb5k1vzVQ6vmTULRT
JGGWdwV5Be1Eq9Q4x1PomZFe4cHMaDKmo4aKUxLvYAP7feO37YQUNRl9XV6z
HKe3feq3YkzTU78VYMqnckM7nVshnwQnVLDpcY8leDuvUuPajeFC5G6l8FQh
ekR9YqGKo1g8aDVBlNkb09hQV8nWtNtyz9O3g30JHZItFKRa3efLEoBa2XGE
Z0Qhh7Xzu/6BnkYoCFMcDR6bfKWgBeqEnABOMRrx4TP3OkBDQVNtaz11BVko
RHbBTsPI4llJO9lnUkSIxv/tuDEQFPKSyGJEjHIeshw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EyNQRoe2+uX+DwiCq/oXOLiQKfZB/1P7E2CioouUh1mJYj23lQYUDTewJbeboHTagbNYFPvOMqZtmoDF5/YaWnMk5GM1+YW9S8BM35iJkArKo79uWbSPVUWIAkb/+Evd5GcDyCyG9ZHULCvGrQW/LwGoUUZ59bd2rAofCJW4nHoqVznG/Ov3b9yd7UweRxfRgy7LKjaHJOHLQWjXXJnJ1fvbCevRxOi36ohsfw5nFpy7XJxNPKHemFduL9faGpjaKBLwonDE7yQewIfzukzDPfjrWWLLJuuvpDupwZaBGo8X6VKzMhS8NcD4oh9qHgJ9128NHrvCqGMROaFCQwSb0ylLeJUmi/T37yNFqYGH4H3iZndBvXev/3wCcbLti6EWcp80gnRHhamnPxWRsxdtshVTQcdxWu4arHuJpwTWKBXqmWVIRJmLijNfA0bB4oJ8aW+xmmDer++4mtoq9RoK0O6/L3J7t+zX1VlO2iZL3MuNG+U+Z9afSVP4mabzMaPzWGHXRn4EJIoC3WbkkAshA15981Ckmi4f5NwVPvTjGA9Qxkpc2E2iA4T837wF5q/oHbtrc74xQ+aftyLtbKhwVIRALpu8XuAMh9lu5BE0/USNGossAtNoVUaMgvhIYp3uFpYV2CpQd9QqzgbFk+eslKZXTjklwg6Flp3yLeVL3pd5oS1ErxVsdg1f13A1HnRUi6Z2/sg8pX5WMnfd4g24EUPo0NNPFmebDT6Pb3pX9FbamoMemSI00a+aliC8QYNrnkXR9jrEMszNLhMLMlmQvsx"
`endif