// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fgHRA6CXnJtI0KWPlBq8G62WIz4MOBEoQWhPk6Tm/BQBYZoN5A2c1Y2vZZy/
SJzjxHUs7nlF7xnUpu7buWw2bZcjcp+a1FMuOUqJEqEbUXTVxDZlAQDrxs8S
TJiVqIZfu9dSLyxcVLCQqDmDpHII+MObqb7awvJySek2f16GS31yRT/PQn6+
SvR9DRGdoUIvYeHB7oLeo0fvE1kvfCvmkNS4TLJ37msS1VRTi5z5HKFusV6v
wLFtVTBC6oX4TuVzGYRz3tbMiZA6YrtQQDpCODU+QL/LThNQJF7UzBcS/k9K
IYnY/rIZvFy/mMRyP1GUzV1KClksfWKROHh9VyUdUQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fp7lrbJI3CquvHLMNZNqZGg/9P+KrjBG6FLF+/HWWiP98Th/r0GEhqkKl7m1
+1WTSlBF4Fvsk2yYDd8Hv4YUf7aHuo+V2Ip1ntjaFs7icuZ/jVWdJD+HtzuF
IcC9pRD9ER/q9BJO/5PwK8ONBrsvSQQ5evAL3hXMFdikgQOWB+CJytHgwZFf
otZHwOtmHSocA9FGGgWo153dIdULj/VPDszOEjywbnOQQaHP6vL7PDFm+O4r
SM9JRJdOJ7cNyXDqjydz8AsKq1OWlKcY0nX6Hn861vYvvmzko1RzwQYlARPW
Ghu3H8w69PorB75gFmXXt6FLg5CbzzxYeQ9u75/Eqw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qJ+in1kU1NQ4erqYbgkNt2Q0lREtPS/q0RJ1XKmPwpk9Wm2nGPS2PZ65TK8y
ynY9pnz/9pyty/4AdgTGgSWEHd8DaCqkTvjioPy1ACxAYN/txufI98wyUJ24
jFlGGDbXBagM03RC/ZacAPF4uOYxANoIiSYEePoE4LzDGnM7zHipep3bXYTY
NMhSpI4Uxfsb929yudgXnnKXM3Bu/E0npYJ584tWkkzPlsPt9gZSM06t3CFv
kJppn845N+UEa1NoC1R5VZlV7XR0NUC9dZH33zykP6vHiThiSAJ1Aygfb/na
7zQv2jXk0DTPO60Jf8Bn47TkZg+AMYJhPLGGtss2Uw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KHhBDM+EmkRdd10Z6l1HkwRpplNNZhqkMf5o0ThRAwbgeyrsSV/S8+j5jxjz
xXYpYtKkuxunkWcpxjM18ztl9AeqUCaJqLF4rvye7Rn49k5xLGrTMZl5Pzhi
AcwUlGIiyRzO4mHXXpzOYILXDt96/RWLaV9+W40vNTMPvFROLXsPgzSAI7kZ
GZPcYeHFP52834gk9KAQEsZ64HnoMxpl3J15kIpTdvyhouRUjlWb0DqED0Zp
anyN6sUdKk3Ahqz+sQ9ocTf6Zsen+jTcF3HXP5JS0Vn1noaR/j9NLAo/BRHv
oz2Lkm3ElySRbq20CNWwCoAN3t4PHH2c9WpxwV8yoA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PIzFtzDXk8pzbYwrtQF15d1cJRFjFTxsiVheYG5TWNPvu46U/aSq5p3F/Gic
Ien0YexhBFZofW5u+of1P1ToPP1bkZEK86+fXlZsk6MAJlV2qNZG+/YaBeyp
H3poOlEcSFZL7oAJYqDyi085FYicwGHQ5G+G4DMGO051H4u/YU8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nzr3FciarUox3dnpi+OKu/WJifL1LstD9rWW0YshV8iy5RpKWicF8Zqqwobo
085fmAe4zyTStgbFfiJ9eMwdywkReSURj6OIrkMTPKHG1xqb0VOl1jz2MUGd
oswz1ncJRUJE9WwVqoI0oV/KJ6vZ4mQDbp7OlfyMM6paHUilRrJvLsRztaN2
y6yxUCb1RCIh2euP3N3IOhf3hzP8Ka4om5Qk7D+yhCPC1cRPBm1a+V7SJYdC
SJwmVNmOdQUQdH5a1ntHcBCIIjHxirPfuA7bgiWjWFrTG+MaxfPTNT7+ns/U
n1JCVp4LHOjp5qoAVXr9ZvSKPnfbLt+ljbKa1PKd5s5lWNYR/4fUs7PwmCxi
QNEnp8xdOZ5qYlR/lYw0kJ4vjGUZKxUzNxfE/fGguuhUFKvq8AHfykjPHVR7
0pl4H1txezXQOpYXSO2bkjEedi0JMm2+JB6+mO1rNzEkApgmPbqzLq9BfDoi
YrkKRCphtCnlKbxRRXqY5h7kYQlOdfbO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oBsMFn/PDrZ/3+gthfkD4riZTDiZ4P6IBLNWqR1dWDgwTDwRdBkoI2xQg2Yl
Oa4PHbgtHZ/yHuSRWYcpInTfalH570QUYOtMorRvRLRKjjq3lN4U6yEXU2nc
MoKfCB0FE41vkm9D5mgjRCX6rj0KZYRqsVcx5prj21KjI6Ga3xg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
leIjuVzGIUyN66J1nYwvODZK0B+Me9OCmIODmXKmA4X837apmZQeWsw8baPd
sX2uZoC/uTYBRPJYxdP9dfoO5gUoBclxtnQuav8lPpdVYXEMvdhJpSQjyme+
UqjZ5tzZ/74jImJwL2b1ugEIAR1QBXEKKw3rtI5yVLBsThvpCcQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1344)
`pragma protect data_block
8HjnfY9JSpTr4hPbOXIK6XaE7RywxSSBCRkmTGftGDAZAUwh24NdwpagKSUz
ffvwgFN7OJzEMKJpe4MP/C8GOHRdqe/FtMmuIhYNz7xuNniy1ncNgpuyGpgK
2KR6HJ9gxAA4Qw61Scp3cZjFoA6czr39tnRceV5nDbMCdzYyEoDKxFVMQuib
lBjzz1Lq8PEAGHn2R0zCGEiaga0eGXI0u3lOVG/ir40NzOoLtkS/MomGc7cs
/AO/TIGVfeBjBxx0WoNT6ilhME/5D+UGMdhEu99JwODdUsM0kPAfXlW3IzYn
l3ee1rXzQxUtgabK2CUCS2XvTgbY2RAAakZTFZ0HV22upajxcdA7kmJtwHnY
dVqyBnGBajig/KM5dwiZAckS+25fMvX+JAjgnN3OahoZzwiZlktjxEGW1BAo
MLBpKXiQGiVA1SUCRw75IJO0H/7SgC8Fhz/u1S4sFkvrZfE1HzJXuSqL4Is9
pOGuFC2Owy8gla3Byqx1OBUw1qSfQAHHyzgc3JXS484Fyd4vSQBGWq3phj97
EMIBAxiBAhe2KNFTDcuRAHL/GmHCKpRDdO6N6IOw0UMmiUaZvftPIzy0CaZP
QItCftTXgD/W1P90xWQgqKV1fwu19p6EXK3CBeEQkHQw6YawHjgIUdCjfm1D
uKPKPqBxLwuTtgyMMfxKEf0ZJ+pG3Yk3dfPMgGd7cmFskpmcDzPviViFuf3H
cuJfqKXoLTpzS0gTNAZ3KbWc2u08BBR+Y2IQ/p+V60V39byKaENJsEalcUSd
mVwmBYoNWIi6w1JOuxibJZ5Sk2RESV4pcZkgP5bKs0F1Lh99wNZ4vYhwiuOa
RH6uLNcIp1+B9ArUk0szWKG9EpqPvLISztIkpXif07hv9OVX4KgphIGrFEBL
xnFZnFPAFH7i9tEmuHte5DaGq++OCLeJD8S6t05wGcIwwABvdzM09O4xwmWG
o3ug+8VL49ccw8iSxbOG5JBa4Oe91B38bAUwuS3SCMW5ETPOhwXZhKPh2p/4
MT+KqgYXPj+i0gwELQrycOvGmgq1Jh289cweyPXyGhh9qlnkDq5C2KCJURFi
t0KC6xUYHW0CkbPFpxm2MaimhenueWQld4bjI+Xzd0oEm3dF0cUgQMGZdmEW
ykDmdHoEzcpl2+1Ov3/qMa0i9wpB372yx/MjePvBddCnW7HsJjtyfNi7RzHK
23Irk/Pe9f94nJneh67u+/ylcrEGH4YU+HjwK93nLuKkF/Jn5WpPK9yGrY36
FqMEr0HkroHt/PWGg1EIIXCCnHOV6d0pmsYdVI//eNiK3GVeAX1lSsHoa7Tv
RrqWc6xtG2MeDEmAcU1/WnyYF9xGJ8mlB/Uc3v8xTe/TepfDOLvUCaz5aUZC
V7NmlKc7hQ1RxOCNcplZaN9VCze0bJtApMWRa6KBWH+9FRnohkMS+rAb1yes
qzboSlhc7E4AU9KZrdC7kddRpyCIXhTOwCQZMQRBNemJSvaPft4jAYdYFNvs
NePF8SDYRuWA0bH+TTyCszU2VsTIaqbtVZ/Lhddhw7cQQgFlRkcf2DzDB1YE
mfndyGbegwB5W3z1+QA/6k/E84KV2vGBbqkdWnQvJ2+5JSpr7yWjOhQ7U0T3
/7OQRdzGFmhtk0/Xtz4gaikk2/i6epia3hoE5erhLujrj7hDRuTwzbmYzHS/
g7trkgQTrQoyl0MxmyoGDSCyThTB2lilBNDeu9wrFRvxVVw1jc6mbM2UknjH
dz5eVZn1iQxd6Ta8pq0Whg5OKw5p20C7TXVB3XKVIgJ962YhJF9k

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qSIhiVymWchVPUjCmpBObCrqaepx8xTv2h2qleBFj0f0+MiRmGaaer4/KeXxo03vMbvRUIydeB6iFTxJjRLVLR5k35WAv4w9GKSBJAp+/aenutmLFO5Ksm0pnGR0a3eqbfUOty2PkKaBvaR51ttojUMoyoQMhrlz/bVqO7fJt6AlunfCY+jdRbNsUDinEI/MueunUVRTH5PWIYGLRmqFBWV69FwOCnSWdQqZ6ruRUjZsa1GqCOJwCD0T9BHo1aCdntgLMYh3hPf9EuRtfDuQwoxv6MvRjtSdJkzbit0wABym6W+RxxuE6PkolGAWWyZxtWhViXYx+mMzO8vBtbxeAnk4UeyzY7Gys3uFW13+U8ljMb++LcB1Au6oakQRWeD3x/lgeCKvGegIXM6OabrLiYuJ/XxGCFZRqxejxs44MGnsO5ZblDcawW/WSJPSTzLg4088YCr2KhEQKVPftlxwdst3OhPhgsmWAIngq4I4RMsRmXSxGAZitjypYatOgW9aDuxJFSv3dr9LOlmAhgnB4lAGlLPh9p7wtaByKpM6t7PMzME6RJbTe2UDfQwKaQEVicAxLKrHRZBSZk0VK1+HRfzukh7tusBvINf8PuiHZTW/qMfGth9/AkwGmT8dwhuM82yg3fwP7MEtqefyW0QZvRcaDF5gHmsv1J3efvNUk6eoaNQsgduQtT3FdxYr4UyvseekP0GFCzR7walm3CraJTU91jKhBOGA3xg/k2RZk+ZH4jqg5ke26EGj6nWkfnu4o3NueTyhS/zSWoHeBJgdTJg"
`endif