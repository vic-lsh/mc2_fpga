// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OsqSBQyU7h3bD0HYNblNa38mBfkSGTSvZTkBXuNx0cxBs4hMGTKJ+sWiLgEc
yRAqRl0zxdJPojAf3aO1aoFvzsMq69dku+UbND6Bu3wxTYf22JGCniLpp2rj
SyccPEfoJ5YUgsR2ZdwirSBg8VTTIKQ0H4KW2jlRlWFuCLRaroUZT0wm/ry6
LchhpB0c7YWg9FANrpaLTOUIWoq3qUJ5oTr+gn7Cjul+ot7WGYrVf5cjvXen
0MXHeFLSvPjO1XgaoelyuULly9qdZxzYxLK0ycDRdVYkqWn2yY37BnQHtbxB
BhBn6p8NBIrm8wb31+AJ4SMq74OBbtY5KU3j/FKSeg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SCerKiuxZwrIJTVZYo6zgwmAkXjAV/M8qSOKPF5yiQ2NBTmI4NYyKR+SkjEg
UqjB42Ol09z2MGQkfKkSt367yqMkatUqkMtf1SfxG+g0fjgxG48yo5fn0fSF
cfKXqIVbee+ACjj4rHaVJ1Zbqo7qzJJtXCoze6JFBoDT62X3F+uPn5OtJJE7
TzcrLVdogE0mN1alnbYHxrolauot+mUbCgjuPqck4IrWRUAKKhulSnvnuSv9
7LfIwscYU/rjQg22WoH1Q87YopfidTlpUAY69e9vyvrd2ruuy+FVGg/jx9Rb
Zr6pt+Jda8UNozPdDGYXpjjoGa7nKA1Xw5VY9QcV+Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PGlWe5ENVAVQj0ordQfidpcsuaaPkBng4dMOK02Bdj7X3KsSR6mAtiJo92W5
R2azTzs4E5Nxt4b7gLJ82lsUCnUVCe+/LB3p7UbQCeGOjIwmYcKrNXU9gf0q
E+VtfVFDrZ2ZHvtMH0UG8nE3Q+OnInP3eWpqQQx6p3oxC1aAvAxXhvh3vvw4
2SCumC/xP0tjiwzpXCUjqtxz7fYYvA88nY+LxqhGKobcPEnCiHR+pN6E19BT
2kC1wcGa6wJaqw7gjPPzBYFiX1y8N1nENpZX8eTNf3+uxjvThJLxM+Nn5fgM
43tCGje4111zcN6jKNtA0yPWw6X2i6P7uhtfdWjXPA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EtjaXIdhXFvcHWJfaWaU2IY+8WM+0yo0sAlcICAHO/F4c8AZkfuTSX4wMVba
1EE81Qi6tMTPP6juqBQ6q2WMEKjUAgA+w7SS+XzRqHJymPs7/+3NAHuIfw2F
NWGkoOg89Bvd2RSVkbZMLaTRC4sV5ipzLhpqOfHlMlb8wZxF2UbHr3jKkEGZ
tutaFkce0IR8J/Sn0bu022LtWgLywB9eWjav9kpjvRS4melINf1DOjpUa6n+
j3JdaWuKLEp/Me+70T1soFS8ZXevUYpL0FUKqVPDL9WHTy5v8Byij9/YrtxB
Wdhfc6IUJNbT/O+IC05hdTBUpVDpcppS5fI9468M2g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Om+DzAobJxztSfy1IBWo2M+Uamm/C4QsN7plgm9FZUjb+URQ9iziedSa8fhE
ixmqxyOyGFF/9ynAaFo+FjuZHIotSPJUW/Nge8fUrSSTZk0YhSnTm/6QQyLj
hPoYoUoFzla+m5FnjTMdmccz8EF+qafrlBf/BrZrYc7RIGy5sjo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Q9TP8f6b3vc4BV4uG9LxufCY6xFgdgysmKgscltlLmgGB9pWCUkRlIapKUUX
pr+HIxpdtelGdzHHiiENw23ZzM3gX5JbGDD2s8FvdJDNLofzPptnF9V436HU
NUhlPJxs8iFoMs4rqiuTjzbkCIBkHCKVo1wOMfISPzWdmC58l9DjXR9LCdU7
sCcbGL1BVxA+x3rbJvWH9jC/A+22uSvkvNq3V/ai/pMTP/nPA/vUYosiK63I
et77zM7ZyVAGhp3Ovh0tZwt8nAAXN/x74xuJn74o8m+Utp+/7MO3igwfL90c
8+0+mCdhoxWlVkt8JsSsp/TCEel1ApogkrC/ziryOiHQbN2jMYAdQwL8PmZ5
WyEORq7/e66vBjB0+7v07VQaRGTItUYJ5lL1hv0ZlEXrhe5IwmLMIaq9Gt2y
/JtgZGA0d9LBOu09q8b143a2MzgQ4lzI1RPskrWm58Ns3GRWN5AubPx9vr/m
u8YxmlZrthrtozqczUOV5/qWYrj3QjZ+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ILMbHz3fM6JgeejgpkO5QaQ9W8bTTAez23yC7q34vGbU1uM2c6h6+PJsVIGH
+RJH7ZU7THIbAnuhsIwWnhc9f2+/Vp+NCjjVm+s+JDF0dfoBXuGv8xbSGl+L
il9JaqtyMIMyWQFR0ovozJgpSrig+Z0cKfgZoFthi10D/skDm0E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VCBB7HVO+PwTwJkyjzBB+X9+YMT0kgBsGRXFIArhJnz1TaptAvOt8LLk+2K5
CMeKUuNkhlrdyuL1rr5CoS3w1LhOsc4FPWVV8Kj2pHYmwG+WitWK6EVJOkOg
AWhua8cmyXLsD9zOjBjCUY9jaUezK8YQusyFs+yXVLqq4Op9+Bs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14240)
`pragma protect data_block
NwzuU321QjYZtUq91C06QLNEcDuY0uG8g8sJdlAPWiJqZgDrpGeuuBmKHCk0
jrc99u3aGXEUOT+QD/tP+PehbJY5txMaPkZcIxg82lT6RezI3/van906M3l5
YYgP6MtCPehU5XxSs26Z8n7EWEaEUITSFK4HzYyXgD7y2zx2ShZjp/IM0ar9
wC24FhYlbSkUs1nWs7SdKyLfEJ+FhI+7VF1suDuSKsgOx3Ha7xAmKzVwtqJq
q7RTAFOn8fkH8Ur+1et1L7EqEEoJ3fKyc2UegaUn9FTs/5SlcfQ3BMdOObM3
+MqgA8266IdT8MOn7fwhNdJIDe8TeecsuN2Ax03zYfEkEwZfu/hAYF+n8ky9
q9gh8qvsUmH7HQA7bsZ6wBYsuaXznZFwclhoKRkyGC2pOXaonaW1v1Zuh1jN
VVdftNEVDEQgr4S1UE5/RyJjNBGlKKpKQ0uVBPa3N+HHsLsRI8USULkfO6M9
vIN3TDLoW4k0ltjX03MuyOKEkmwRgc2w78ckiguftPqaxlTaYf8PS6k7tDhN
WXNJ2Nr0+J0Vqq0jHJTm6CMfjgv0SQz7ZlHqVn1pBdwnd3mYJCtWCAeQ/f9e
/RzK25tNeR6GI0tKjRyTgd1jmybZjl9IexoakdeuKsr7JEiKFT9DpDNm+rJ3
lCyJWF1B+4994TD3x8jwDgnAIAcZ0gpt73Gxl4jo/pLSI5gXxpnSBztFpUiy
90vsmx4Jl2CmMdPUvHlDVkT66Q08IrruJQ5wxIcZX7pHzb8rqYfBeeXaY/Tq
PllOHPumQuxm6ASoRE4tEpcYZnDqrh1tOqk3It3PQUXAoDWVLJfghMHFgU+h
R0yUh3caZEKg/V0UKvSk7gTG9Ax2/sTDIy0sEfTpLmluLjnYxNKupZdxIXPj
QAea8FKdDgO+6jkUF2CkbHm2dXiqpKDLmX76dNqaAfBwOlwRl8AUFYFau7ML
bfrvSsYA9Gq0xCWm4e303FEZ3jHTKadC4xy3D3n09825lkZfaRa1SsjWnK1T
NCVzgmnSQiD0QrdIh2xc+jmXzTl/iJFHRxbCBWjm71BH01ne0K5RADc/uG6N
TrZjMKA9of5x2wL8ty5iPFMeNORZdllrSJZXXGdNWZug2w9OzPKvSJldg4Sj
eGtXNqWrUwbXIh52nZBErQnhNZ6UZztcCAIq6MKToW3MQ8IhL4QzCVJmOEC2
BF0N9Xxmol0KZKJfy68xtEKj17ogdT7gjzYlzmqrROGfybMDChmJy+nTZ7Ru
dlnxM5QpLudml8EidKXVVVXuruiH6uiveyJTWrsBxhhKWrJJi+jXhARUgFQt
heLcEIU+jzEaDF7ubhTcnkUKxt/fs/S2JBmXLn7klU7vRTA8L0I4wK2mWjIl
yCa8RhZPN9BmffvnnpZPwcm1TQvi9WDi7I/o/PXTIz0LH6UCk4JToapfgPfA
m9tHiMxdhJ6uA4Krf9QKEpTBjNPMKbFzZkCk1StnWr8nJMeNduGIOj/ktlvY
q8KmiNwTcsSjjfhGS3Vu5fprrl7JpRR3A5Dcpy4J6y3aus7CSj9rUN/3k9tf
uwU99kOuA8sR+VuISZPnftxYZ/jXz2+VWejC0Y9M9mdCaZsPkAr5IfIUBJmw
AKibR7flzzKJYqV0ebDHliRjXP2uc9BX6SGCtuk1ptzqGinnyDT+kk68SBBT
U36b290Oi1gfEdUX7a97k7xQzROyNE3qQvqneI7c0WO1t8bjItvRK3aoKB9v
anPci7/vaZsYu0+zxqfNsYy8mwxymMovyu5RQGx+MFvDi2geb4RFZa+Mq4Mp
Ay2/UwGmXp/PgAWSNFTUmUGfF6HOOQdy8Lialk1jCBMdsm22WNA+5EoYyeFq
1NH0c4lU6LBXBiY9sqcjksAZy7soePJkJXqMjUfdwfCbjahQdLdAXuGDPJv6
o6OOusfSygQDhKeg6XeQahVhPk5WCoAVR3z+92tY6jmWcZME0aZClAoB0bt1
14YVUGYSoS5IgHvCgWYFp+wT+M9klUxkRTn7G4vg2iQ/5b9o81EVi2hHskuQ
1oGIADqoSU1Eaad0Bvk6aBbSURDYWJTJPBqXqg48tKZw0C0SOtOsXm/yrlq6
CkRIrcE7BxWSFExPNXlee0EA76shQ8XcNC+VxAuWnGhz6jIYkjH4x/bhb4ER
qV2j9eB/InDY/AdL7MTozABVYfj3IKdhcvPt8eejmAdazEaeCVUlL6Y8mhr4
cAzx9W0FSTkCmtYKqsRgBfuT3xziAkR+IWMuU7XpvumzQKoyH5vapjWLvv5d
hiTICuu78ZqKJt8PUBUQOc10pWKvX/FHCBRwnZ66t5Ncqv6NYIcLHupfSu7a
JapXNE4CiYHQX5qt9fF7gj51TsOF5PwQ4qmw8ZN/9ZGhMG60KPwkbS/bL/6z
gpnXXH9idOOaQbLz1C07QGiklwQMO8ERsC9SeIiroM42a3bB1AFI7t5lhvQe
FVKA/wh3+JT3WKg6cXeAntI39GCNP1l6dyN6QJn8CNAMIXfQAM/1JvA5PmqI
BRbyDdp8b8VP3Pvcf6F0iEzEWYRAPWUnLyAPzFlc8048jqgb1Q6vnBOOm9kl
QQoCAit9o8nzUERXtVzkPJuX/QmsJ9ZjmidrvdeO7WawDrd1nHaZKUX+QjLO
jm86RowjulFIb9MhMpeu3CIl+/AKS4OFB87lCgZpvH/Gc+tOreByW/w2dqyW
Z80ro4UqUMBqRCGojCJG1mcx8xqZNlcrwfCskS87Yh2tqnlbVI59Ot6q1TQb
upiCbZDgrmWkZ2NeuQ/pcdKAdh+YDN2fdKrjNkLdieZ0lYoeNS5tMe4HYKgF
6t3gnM2mlj/xsmdiPvhNbrkL3vuUFIRe+U/49zE9eMKl5uoXosM0w2Jn+fFl
1xjiFmP6YVmQsOPWNdW4+stkYjX/rMoLI9apmVeqWoiYjFig0w2SX/+brBQx
Y24mnnxKVtb9XwWir40AhQqOXhsK4AKPq3WV35dMMk2oVbd0svN35EgToGXT
02q2MgcrBn/Rwb+xVV6v8sjCSic35vtqBTWuOEgB9ViFY7Rm0r4w4AetlkNo
rINXsoUL+vi1MOfp4yhyLisIaA6/Krw1+25vJlnbN53ZalbHhVzRoMFiUbaN
KTJvz+RV/uzlXirlCIMLCBNFdzQhfGK324dz6M55vkvJu4pSwkQaoPNmaMnw
UjmYLmdrGjN8K7EOlI+qHw0QIjWiEwnqXT6wMmDiNiMGTXASB5bkegkj4UEN
Acm9qhsGpfhRZjg8yUlzFTD9A0IMFCxV+NuNHgZJXpitYeCTB493z24TOSFo
4OSYMVaP4j2VFCEtJ830R4nBaY7G/Ks5nn57N0P0s1l22Dfj5uQiU5w+iC8h
YIL2j9LbGRfU8v/NVSngLg+mfRNyMzoVtESBnJAxD7wWpEYStAWQ4YCvtRH3
FSpve246seoFrQ4h1bD0tUJJhcT/RSK2gH+/zj79K3GJe/QQt+s3j3tHHgRU
12vef8oeRBl1cTMamLsWETlsxcTZW7oSQ6n/5NmEvkxcrIGylBlMFThbrZ4O
BarhC/SOdIAGWTCmtkYABSC4RPRWb7vddJn6VrbhfiaUOK4TsycPDF9oFVTH
J19C19o4CobmdlNO9Ii93fqH9C2jcEiXNcAu18Lg5HKrhz+dd3ZfVkxrLKpT
lV6r36U9hcSPs2Eh85RNf+5vbbZ0yEknlEoY3UJtB0T3LTP4iX17jVuL7L5I
P5u6Eh2gBfkW6J7NRMQNiLKBxX4V97GFA3fEBZsmARE6Uehm7jnLGY5q5lSs
kTveeMvnnyHdgllR4dz1FVkAvsnVarElDLx44JdgkV7yz/EWxU7fj+a4TNii
vVlBH7IEzbLSOKaeLs3LXJHgpFbycBVS+sTWyzb2CrGYcoP8lEdvXR4cjGar
fPmMO6SqIZ0Gi6kAl0wn8Upx/NiZJalV3KoLjnHMFZ51hNhLHugaipdJDPcd
zzvNcC7Dbn9vD8Wk/ky0DktKiFT7QYaNu/QSBvsffpItvhlFd6ft9dX44HQP
SjxMj3wtu3aXuwHpfKreVNdMDWgh/4OGL5H3Um7gu6vdpqFuaPFfok6LC+oW
GwenE7+wqvjNi7KwAQhLMgI2QvexzBT78NiOucNI67z31xDg2byYOEOhWQ1c
PYsD6NcwE6CmjRgDUuuBVbmXokECC99vZ+djBWevrlHBmFP7FhJ4yM3j7VKx
pg9PPZ9ZAyWfhZ2HA0HADBX6f+Wj8gm7q/uzDuVNtJC4vOw9lKLIV/7GLx+6
8Mu+s8+37OFByksEmyFepB1O7UZwcUOxfvAIbnsKdrYLsI2pp4PIvFb7dmJV
FZqXI4qIlswl00yb16H4o1w9FEkpKu172gTdt3J09SEzuaVf5WuhEMlCxg0D
jgq0YZpljlMIrmoX9WbVCtufYm1XtqxnYbxkvgdq5G+9yh4DVAqvD34ebnQj
XlNJ+a2O4qA5UZ/UIzeEb6m/vz/o/twISoV9JcD+ykETxv2WqfctF7nPn05x
IV0NLULE9fPJCetEtx4JqVRvSnrdZ+yACM+FPiP3vf3e/R24aB3zXkwiE/XQ
Iy2SwFvG1CRf2pIDFSoZdsqUR9lzxrsYhyiYGB2HRMupKjBk5ng6BVBYenOk
Jc0KHTtdomTif06KJut8igX1+cb1XL4R71lcbKJTZIBC22FrPjEciPjPzoQy
a0Vmsoq2h800F226lbgusuYO4JPyWUS3gT0l/3bjLwoZd2/ZRqWcHhji51Sf
XppeaVX58VPRnyFhSk598D/th9pzPpVwjlZebvvMNq/BH+i+2Cb5Ow5U/SGg
5xlAmUuUDfNCd+2mxRzb7IZ+2slZS4B9OrEhi9cJgAuGzn6no6HLjKEFSUH8
MSTYlm/Q/GXNv7vhN0YfJscda+9XrpqyV8/hjnAE9bkA5jq4BQQYw8mVRiqb
9QTGf6iXKwNSvnl16Q+FRMQsNEYfySvUD45Mi54ER4gX71/vJNrLYxBYTxp2
p+jNTTrwYVflilF0nRgABgfUs+okp6s3RBrq38Ax8Xn+korMzFcK9XC8dsv7
sK2/X9UwSwcY4msc99UlHUtWrSIIX/ihINaxLvS+LaBR0sXoH17RJVFRRpvD
DoBIOcV5xaiKj+vqhtd3EM8X8rZpJufjzefE6E8weYNeuNVyCh+UMCOEiCSl
yRKNhB9lOxnbnOUeMRhSL0nE8ieJiJiAkblqeELK+ki0Yey9lcn5XaXiG7dd
716nzYQdHwRgfCAI9JM+j1n9blO4Oeip3EBOV+tGxtpvjRBbm0Pvnm9KpKQm
PiOWW2rlpg/RP+fbMsLXz3aoUZ3r2saUBiJZ7In+d7R7CVrd9YoDjf3bS6B9
RmaZWBuvOlsSaiTgZk0EfTQbsiuu2qs0fw44sh8BihkbsOEiiWcz+TLjzl3C
ionG9d8P8UOCKuDKtZxRSIbsV8q77EEUnx7qorRg542EQfy5QBo8EoHSP5c0
oUSXEJCfTygUwdZ4wOPfhZ4Vzap7pGh/kFSqpmoIzApw8PdySaIRr4sWoku8
7wXHBUz9H9lUYCyvm2Fn/5ZfLlOceUXyCSqhdKWCepxmaWSlTV3Lnu2tkJG9
hTuSnNV1CyVn9jmoxpia28vWoMEzkoNm3WbMexzD9d07kCK5Cw9Xig2TRr8d
YRsRSv6JL9YhwQOZK59aPPcstgcho84OS33tW1+k278ayDhh+dQvb4TX1Zx/
EQKoKdyEn+gIo7F65jHyxn/4CTbvMV/nGqj4mrpvzRl/7wzyztkABHFt8RC0
/DUrhJfRRvy7Qh658bu844n5NOiXBBxdFSOJV2ETTJjgZJr6eQ6RPJHJIQ4C
j7RPS8tbRFr+SLwliT3wVY2kDefa7x0XXSWlmfGBkn/sxw/po+HkF6W1Ky55
eGMnOhziRq8xBLxaamXtPDmtiSw52M3NLiMIMzmagkwQXC0Qg3HtpiTYjHzw
WQdvJGvGd0erMZ2Amn0mqbSG2Oj6IpG8k/RXGCrUmqLWfq3sdwCDJvJrkPop
dkiDNq/SA03ekLrmis8GNzGoKUPjhYh5dQKJo8IUf5oY+UEm5r5dWtfOIWlX
jApECdcPmYC3ei+fjtR2gByW2qDdb6xdRDa4OQd3jVbE6NC/uU+0XF69AdsU
g4rwV0+0mVKMNWyhzYMr+OlmiQuOPgx/5PnI2yRNAKqf0/CuaC8FRMN2k0Cy
/yILQHAltifRdxVLjJuyC/W2DzT7jWJPqimctvQ1MGElwK7jqYSoqkxEA4rf
Ehf7SnLVAweWRFGOeBjxpfuE69eKAB7LygihE5M2CrX0WeBbXjf5dddYS5kz
faswveXOVgNOaLDBEH/jfirMIAl6OFjyrhna7HEGmRJZfByGgNMZ5VN/pBph
1OJJHd1Yr79UnldOlmxwoAoTEoHjSU00Hgh9O83EsFlAz1dgoMAzH3T0BaOC
vqZUzvAtjk3uCjuu/RwuYCarTetvxPusBVoNIc5+vo0ld1Qdsyz2sffG2yv+
hyzfdPXW53kW0bkGqUBErSywB4lK1XoV/rO2XeVhyjDlIuzlU8qiBDHpAgMG
h6DnACgI4zL9GDoaWw4lG5nIp+Xr3fWgOAspVE8RvrV7aDY1cksql50Yfylk
EDiZyczw6ls/m6XhvLqUGU9VCTMSVNJ8xWuj2xbo+PqWBF09LjTdqYSlUUBI
Df9OtvaEbouSUihg81QLFMbpC8lz4SVY2qCQI0od+lrZAR+pQdAF0/IBV3bG
eBBl16Xch9qz7xypm+WGCq2UGKTyJtQCI3bR5Hz4uUd18jSnEecU4ghx7x95
CncI0m33thQSEFlyTj6pqBNDV2Ie+hBJV/j1A7+ZINvRy2psLTF6tVFs0OWL
76g8BMMfQG+plHWUA3mmEwJMqHysUOJtzn8gLgVCmHy8MKwfv+jtcSka+4R9
Y0gQ4cum72f77a9lETiaxpDwWNoCn1s+rpqIMHHpYnI+kfX9qJ/+ju4KczTl
vUemNvJN8fiEqtIp30Xxm+KUmQBEi6dZ735Q1NBmNpTbMDbAPRrRY0XAIN6q
rYaaQCP6WQylNUyY1E/aXbPI/TVSWJ7YaPTU4j6xvZ3yX4u5sCRNf157HDzI
kt82WMOyuWLkioNid77zHKYSMQy6YAm+UUsUIHazFthlQ45l6c1lN52IPy4y
YAVTkPqU2kSgJdg9xSp5CJKWQqdiMR24z3weElatMSFRzCrRj1c3xlTtpu6Z
WMR4YARA/UUsid/ntWU9lZZU4JzxGtS7sZ0+Wg9Xau1JEADLytRIvYwK5O9w
VGEpNRr/HFUpIU6l2MY/Aqjp/Zc0+S1BtC21mo49hlCfvesoirIlYaXEW7hA
08OiTV71phlRY58+uoxC19ubLJmiPBBeBJFJjcB53P0nF7YDSyTh0hGCJIqt
YUebWXDiYfZL+EEhwhqXt6eWAGPO4n4GGcZShOM2qoapvkSH2BUfdV4gaurY
jKXvbDz5Pqu1W1QzBkDVjH8NK7VqHJm7TKdtdmGNTj27bBv4C8gQePFuz68S
Tj70nxF/GjG4pEVSn7Wi0wzedxdurDCi2LodOHnjkkLEgRR5L62Qi5cRIDRj
p9YxlQDkP1PP0P9yAJ/BYoz1xqhqtmn7pl8BZAoPFYCs00nxH5zJMH/LkulO
Ws3YKWHNK+UGKUf0qcuBVkHq8uOT5OcnLfFaYNIB3mS+V9ogLrsaR28Ve29j
Tp7DPN89tzsTz0a+niW+LJupjB/GVsjijuTNK8DTMh/k/v3ZdEbZPdxigaYB
iI3jFYtJV8MZdnZIpEJlNpQfkR8AWl1WMln/I0qelHFcqao0NPjVClqemDgf
IKRzKtGPvwzyr77eoy2w47b/c1vOO1zCjuyomIrUTzA90KFLbYl+7su4HmrY
1Nb8bcQxBt+J7ba4iX8Vhuz8bzCXf8Adr8yCDVlCSJPskehY/kcoYqoJJwuO
OVQyu0++m2ewaDIrAUnMVCPbXpaJ5MQW5ux4qXpoEa9QbZ/KRBux/6JGl98i
3uw3XfpxZLBWkugU0bgpUn/VQtqHRlXXtOYVzTFG9Ia/kVb6GOBLlyG9vntD
iPK5gNr546gxP8XqBb2vKuLQRxb+XZ49GwoN0APqqcIc8qqMRV/mTCVKA95Z
iRWhNamgOq8G/44fw1+LC4nepeuZww/h5+Ysf+C9vz7MhEmN+nuz9S/l2UG2
fkjM/3xbXB7ib9wB3NopkGKxxOLDT1jajfG2DXU2VIzBtuaJe1i0DmKbJYj4
+r+IMsHXMZe/xBrwLxeqorI9/zZbk1MUoAH41WjqtLq+0sCQcwFFb82l973Q
AhQKnlccZgBd4lgRpORHGaoDK9T3M1ikups4BNxeiVc7ihF7KgdjSz4LukJQ
ntZ4G+MK/hXkPrUPjJa8rFlijYR5jTW9g58El1hMWTMlo17FjwESpIR6N2e6
CkgSoHsAaUEF0lKXC/sHcPnVwbjwA13GnvyDiPiWeoKGe18jOydDfRzYofzd
nawifwGidzLQyy5trHcoGwz9BzsvfsACYcEgexRKw9JDcEQPiiCnWelp7Npy
cVXkVZRFUnMz2kv+vjtTIEMmuUsAO1MCmaYLhe/E0O28+xJOrQilw7NoDoYu
SLrHQeFCurXacCrntaaRYspiP87ANdz25Xu40aFxqY+FHa/6xVCw1lqc3pKH
bOH5qPrpiE6VIsl3LNYvMGwd2AzYu3IQx1jJa+wLdUvUYNIdl9hox4npQd7L
Op89cHCz8OBoErJ3SsH8PMxosaE4vmj+UTnsxC93Eikb+T3qFMIX9BmO8spz
sIyqnm1B6zA/IoMl7WHVIYoNf3HuIBz6blOqUySaJWG3ug8hCatcoBx6Vazf
HjmK4mrVE7wWkU4TGtoOFKQt340+8J6D2w573qjiWqPHccL24pOr20AbKfeC
Iru8fuZPpREqjCQ9ySJs79yc2FpEWvqvN6SRhOdKKIJAB79Lt89BUSA2s2Yi
JgajbTYEgvlarSoHqequy20U4K42L/A3l1a4t9Q3tHUOV7sYlLYs/GWnHjKQ
YxkcSv94XvqUQmYYkqnMOXMtPJsuMP0q0GFlL0bl2XX9E8pWYfDKgZ3SIfY3
ldl7I6rGSNXLQgQ+mgaf4PC1hkLNFer3qAnBs/V6qe7RDgAfVJWvOPmEB7kj
fmCok6KAKHDI7j95JFAx0FkAVJ1cbZp/tLU2PNHY40EClmR/NSXjtTwFwaJH
2UH5hPqZvPJVuCjV5gS3X5IXhHsFWQrYhMuNNNoGjwywcvqACZRSObhvb41+
yTE+cXhDY60zuqE/HMXshWkgwYyIa9eBRAWKyatJ7tcSaUe/gQxKDP3R/H8K
ZoNE2d4971vHwJdjTIvyJp3NJTowvZusgojb6oR+TYvaQnQuAbNdnnMA5a6a
Nsb7b+1SGRw+ZaGfwCg/jJToQNiDirDiAs6gJMje+N4ykmnBV5QXsYxh6zGN
Sl89tZsD8K1ccf/VvA9uM5D9OCwIdQitKQCttRu2DfW6njyxNAbogKi+c95c
1P6UepVcGIYt6RDxniloZflM2CF/eGUgi3mnOhohNuaEitEGBLtnhKsVoATl
tCPSCV213YBSa6vZMLq65R/t6NBjUbOtcOgu2Y3+Dm7AvXH+U39NXfw2HI/d
NQqqGodeGgQu0lg9+kBe6nguNrcVNExUGyBqt0aO4D7hDurP8oPJq8VQkS7e
0xyM3gEF/AnE6L3GNNuAdVKTuDOHowGs2su0WcQb6gseHg7YrZzNL7qjHmN+
gCN9FgPWetrhcZROqFlbX+pYIy6tEJAC9gpmMWwlEEu5k1G6gR0bbW2iWzno
JVpdhDN16zBL1ONaYBB9nRVEVFhLp9ZfwhOLfNBow/O5KbS+SVVrDpvXNFLt
yjie55i+TpZIJJX4iMSFP7sZxMmdy6hgKo3Z0mZVYyqsDMb6lTcLgaDB7ZPH
6VrHHBOzTNxIGs2+4iEpAwsCzY92qzyO15XBOEMEXgRscLTAYrsvJx45Sl8l
lxx0BrUJyAaVTWsLRCKJKz2HiQ0ZhRgAuNzeciOM3ePh2tbM615fIPrwGA9T
q1hZkwJkEfis08Z5uBv5urfXuzV6rOepBtrR9a6QaRGEjy9ghJ8Dj4pZI1Zn
GIR75BTWBo1iayWwDT/01CmEPdBrrlz0bqybXPFdOHbgCdd4McNZhc1n9a3+
DzrhkILvZlZXHznHinSs+bftwPoSxb3k8gpie00p/opVZNBqtdGdt2WQzMwz
r8xFzXBeX4Hrx+dKnajWg74Om+Nf15e3jimW8Uj/oZGnD6NSVHV7Eo6nnPub
5LfTbCYDCh2uQk0gdfb9NJa2kqSd9hDIjbrfAMYfgLbGM20442+Jzsy0dkg0
8JXNVlALivz2uxRb/BG+UUNTGYjJs9w2agP4Pk23d5pRoae8xtHBQKYcjB6W
spk6q/8FYnYHB68n8SVKW68yqz8QWcxFKLm0dl9vHjh0gS2l4tTIIbAGangj
UW+thUV5zi0zyiC9xPdbUTN62eL519D8WQn54Ls2iO9UrizBBp6mkuOtXUye
SBS/GX/Ud8n+IU8Xys+L+dIxo5YzQTMrgRDPrddxVYUVy8gM6W5nRD6/EiMk
gOSbm9GlwqWIdliIPqA/UNwF0r766D/Ke8aXgxXST1vCxt87pQKlfdekl07O
mvlnQWgqLA06E2Viya42vc45YRui3GeKgNIcu93zBTgKBRtsIEabSjPwsDBT
KHcpw4BvkksW8n/+4tDt01dFBxE0YVcqZS0OwW+zkQwa2QbHJFUlm9U4RfJD
t7vsfRH5DvR8iJEKAt+L3deua8qQLkFJxOgerOAd24/dIyjiMxXwLBa2rhI1
H0C56j2y12+qTTvQ8ZubwstFi7o/FU00CZGd9xaBdBAudqRoEaOURP8OTKZ+
c76AxkTowSJeOKdvAj5atKFfg7nWZXy9y3Q64rWif2B0O81m8AyBPH1ccM5T
m66vTgmu3qyR9FRRKo+2P0FuK6osFoQVzsH9cQzIlI+YCFSmBOe76qZVkRYb
vh8+yDuvlJWx428CQGP7Te7w+7RieXm/VJdt5W50v0m5yz9jZ95AffPM0pCn
jOLfL9HKaUfbD0dOko3Q8kKmH+FeqjyyUBjUTG7cVSpA8alakR66rujCIPe6
7F5sEBOan8ph+fdgYMx76I8BpTPoNAaJvDk4AIoeXDR8TM/n2idGttUBoLtr
DK/dbQCLQq87RLg/ahBrnUSSoT8B2yzHjx++8HvOn+PlUc7HmLbkh5CHYDWO
mOo5FXgxM9fywdZLSxqXRJyu+QYWt1Rlhff3maAS7lR3ZmHUjNptqf8g5ItC
zridT5oCVWgbf/2lessHMkTpU7YqQzX7n47f+u36AXML9lPcxOOk8eOphJvE
ipVBtr2gxdNKN0cZ5O49Z0szdiOUnf8k6zJOKvuohAlp9WVnXqQQlmFuESzZ
H+nlRQOZPrPx+k42yi+4iheExMAySaEj/fH7fPzfdql1cw/k6kj67STWwaYB
/daWbBYHIguZD31ndc3Oy9IenufJ5xGUP6O8MkxeauNner1VYg30UsXl/Cb1
EbK1GhtqPAQU/pKyKRBxp9BADqXIgMwJ1WSz9cMXG/LJ9roIIEnnYdpzH4YH
yXR3r8bsAPUzTKXGNEFEdZ+lN9Ufzl9p2m4+3ZQ/5ZZrnn0x4NOhVVR6ZxBh
XBksT/iH1E2dkiYL7SZL3XAtqYdOl7xSTg6uZxINrCHeVPbKaGBRVWpdSicU
V+CwCAOQoqXqYEEWjDZY4pLDyh+ylGUsA5nKcKocve98p8Y1RFmihyz7/gLj
VSTZAsN0C1yHFTYRS0KvcHd1T7iYr8eJHA8WQJYfG4wT5HYPFMyqpJg2kC4G
NiHYeIF5kLOjGwq9oHkfPyjmRpo86YiWY/9iIwtM+Bycse9BN3EXiEVOq0TW
UYblivPc94DX+FkJ5skXBiByCDTswy5DA8pckrtPzQTmL7RgBNejhQWR/DNb
suSUjIUvVPH/Ksglq9lCKzywASiEa2N/WPuCpwHPUNPlpxr94fo0gosDa+lQ
ZEXBYequ2h3yniDV9Ok8xhf2fkhKP0u77qK28fRAOW+7BzmwZUKuL3jgIQFs
h10wo/EXExtdYGvmB7X34xhbZjeV1forPaya5I2uhCUyhwABMX7BAizCFimY
Yvt5O+QEcrwhJNDFJXf1qBWj0KQddV/GjpDZZHKA23VatBVH8uLHkEX9yCmU
YUQfSbNTSVZ0PFY5HIZ+feR/l6Sgf78gt6xghblQ27T5jrjRKXkXqFdX37RB
7YYcQ2BBAFuKWr6wgjwlMRONqL0lLUpBMNPK7EvbaSq7OkL8SU0RR4QMXYoS
xISWfsW3w9WhnwqR3FD8qwrXcQGUXYnJrrFOqA+tLec181RsNHiNvFkrh9Kl
DQPENLC6k6Ov/AeyyO4yOvIZAMxzdyAL/I6DhQu96NOHiG7ORm+sM2LrPDTq
zEiLf40tvvqTJslTQwfeZwR8bGR40y/BR7y/FlVbQCEChC4ZOR3+b3gjlooj
6fWjAdRL8dDwHYC/hktA/opqmiKJTvkyddJd1HDYECGmpnXt3W/EJHWHoSi8
7D1xBM+zPnF0lDWzSBvXplh/PI+apqT3K3njyGdXSFqK7javDVuI5vn1yq/A
RUcvEl9xaMu98lWldEwLPZhz6DRJ7wYSGUk/rQLqiXWZPq7XBKex6VbDxqLc
vG2vC+zKkFt2Kw886tfYL4yLa50d+0qmJJAOEf2pTCwaxC6oirk24nEXhjye
cdWm0RkaGd7pcUVInkivJiPb0Shuw0b+a82h1o3oeqzCAGznbn9oasakZq8j
Cfub6+44ixDpU/VUlgPvPouCaYlu35TQhRIeJw6q4jWUE0yNQYiKuHoopWN/
Q3cDZSHvj0+NJFyP+UCKfK7S7V6dCm1H4QlolrfyRYORpuXwjlihtT1uPkRi
HNxmJWUHa3YjYQMc9dZhR2QozR4D3AjB/H9b6K+xk0RNrlBPE6h/LkjhVfij
5wgvHHFi3vA6xP5w3jZuOv8U+Ge3ikPyBhcy5bU3iUw4gPu4E5raIvxXXvoD
dQ9U+IKFQmWY5XK8LpuWbIYyYd+23n+gBqSsJgjwXEd6ZQX5xm9OH12PgAE3
z+X8a5DnXmjsYIdwhMJAjVD/kSI3ozdunLZ/uIls4Z9G0EzsKFCasNHc04mj
4ROsswxyuL0AAVl2azoXm9RW71kcbSz9narvDpISPyz1w8/Tk+l+ZSMQ/FOh
KOcDqMjhILcov11IZXAK0q8e5T1JNakyeMf+ueI/RIY20GAzdD6zDsDeEEbM
KmMqFJ/4CrU5bbhu2zair33cIHRX5xW2EsjZ1Vkj38+KSzGt70fExHqYVeT5
eJ6WOkClQnbYAlSLFUKSfOnDRmOyK7RFZOXHWBRtrbSHLdi+0pNAoH1vOrSQ
rKh5eaJiw6v0VFqlxdgOVqh2MIGz4FC84us6JU/KdWT4xM2f5ToelXCVqPdl
fxQG9z3zsH0IHnukMCQrbW+24ff6ME6U9waMKQ1MLYoUspRIhiAWwFmHn5Hg
WxGgOpUS6Yyl1JfIaPyqmLLhEQ4QNUdjBiIFfYDe028gT5HiQurGZ4TVioYs
qx7c/Pl+g9QjQ5SWWARmuhre8VwTZIOrgRMkF4r+R8UvKjEW0NwosIAtVExD
hTD0rLpTFEd1jXNZmtziNy46+rQ2u40HrbQnY/9yTxFsJG4WKaYqPaAKRNIl
ipSoHqz09XWu+fyYAi7fmPP1kf5rOHS77E4fhzniMTOCKD5MBbYqVpfeLMsf
q1G7P7VB7pPl9tE1SdfzEtdyH9jk0kN9iwRcUOjYWR7B8kcxcFnll7b+VIgd
jm3wSwuWRXdXe03FtbvIUDRKsewn9Z8wgkKRoBqGmcs0g6lpvfatlXz9RAqq
joIhxHHY79pbLrynoeFfqhjwyUXTIr/uVRsKE2nVZ9fw9ZJkMANCtcYdvV9s
RtXbpAvVZFt+7qyCPgjHouYiSgRPi0oxhEgPO7ZXK3m5sc9UBm4z7BUOIroa
sW5hPapnJlgY0vvXFUd75ZFP1T845Z3B3ECGdWRV+VSPYJOWbGyk05Z8Nfns
mKkKCY9qFGuMeoDQC3Jri6qb8IuF+7xG+pypFgY5dsbLLhBl244atvXnKvg5
X2YkgB+yJWqLIQI63sNBwUTSGlq9+pwSIohp7htFUgBnj1bKnXTBbPe03zhC
pGQptmyYBRKTRCXTDlhYSzJ242I6aXSORuJSZHD+IeKsIXLewBgd7P7fdov5
HBorPofgDfCmETIfUywf+jdTGyAb2B7ZZ55ODD7djTsmVMcAIW5clVtZsdP1
fpv6rN67pXVrYhlrgajdUdsbOQWXmE4g06PS/xMfL2buHFiMog9mgEtWLkmc
SOECfA/UniwFvqXsRzaTVXaC4FMz8Y0ZMPUbNn9uNpGt0oRyaZyI+a9gvNmo
kZCS7F4X2UNAQ3KdyuRyAnF6+331fUR6NbeAnFEsucfa+vWe5ybPzqCfmLRT
tSVl0nuyC2qCoWUV7wmjoxlU/bzstc6HytHW+MZe/9z65SuSqo88zrZQ7Hh8
CZ08+wfZfZ8THuFH5kXp2VfBVNYUQI/7oLHc4oiZGKk9WOXWfDyrBUSNh1+a
omZj1yx3VuNpMJ/6J+IrcXuVmLm/YpwLNN9aJdzk6DMwZa5X4sO8vMZm7wSB
bbNHMfY8dzrYxJxQ7VJ3esqBQcRwf1y+x7hsyhs2efgL2kkOFtfZDEp9dZ0S
/TMDU3mW2+QghhZ27pvtG5HbmZV3h0n2CNR4F0NojnTwXGPEbXBkqr44U0dm
hDZQCE4joasdeBtSRYpj2ymlhuA4yPPUihAU9xRZrei6XMv0VTPypB0bxZua
BINmjteREW/OU6Fyv9m08wawPjwvB90y14ZF8YGHUVHy539YfDSevLFEwClM
C9U4rlADnMDs+opbSfVpoWzDNqKbA3NElIjYe3Gvo7MgYP+Sh9UkNcpdX6+k
Nyg/JqcSD2I/p4FFy5AJ6zppSD1Vday2e7M8xIM2VhrqYptOSm52o0Wl1J4X
IYKZ6PKrzrwQ3poOw7g6Wmpu6eS6Q2txwxG2cVds5yvSbsGsU5swABAjlqtL
RN1ztveIgemakK7XTiT1tz0fc6atcTPMvo1PG59/JVhV162z18oYz2yA27It
LBk+38a9JcFQpcdNjZQPmHf/mMqexNAk9TqRnZJ3FW+WqQjMddMsHzG/78dL
ZS8CIfwt6rSGBe9K2+CeJ7k1b2BfVqzYgY749NHZHunpPOyW/pheSwzKsw6e
hYL4hkhHm0fK78zL2fscVF1UXsfGoTPyMr95oYRARxuy3u3v+OloTjE4iuTv
eI+ToZQBZEw+WArrymfewnBVYsEjTYd41wphaVBgkYqj1gOrhRdJDDk+oCRI
tSGulayJOB40QkN7sa+hFX54s6C92TKBN2fS+WFXP2+u+6tRdzGSzO300GDS
oHyzJ86snMA0P9yjfELy5QpDeHYHxh+Xkk4zVLOU86v/A90YxFZkvpymmXtw
ttpojlKim6QeQCp4+XtnD7jO8MD0uYqmfhQUGkVil38fIsW1nHzkwiSHdTp+
Jk51rWRDgJCXwbZZ7hwDTmqS3LtJ4gYE+FpJDChjrlbATcb0BMhX42Elf0eM
IO8VoNHuOYS/WypuB/AYVlGVgamzAhlZVeSY2H4l/r8wfDaB99twDYzsQgRC
mH8vsaxFGlzD2n3fMMbXggAk4T945njUW2ELs13NYPaDu+Dx1VJ+3C/VKw3p
d/vij6RrB0V25e0Om678s8wb13RfSOoeZEqE5l1t49txchJ7J7g2sVBB+Ufj
ROXMvFu8ld8uV1ycwfBe/OZppWE1dPQf6ugTxw0FowrN2KlZhzBAyflB6LfM
CDJweMEAKSaClcgUYGax+dqgomfsT7O3tVBlivkYvSnfTnfSiiqH2Jd2Zy63
dPLh7ZM9cg3Srj7Sq5+NzxIfI0iFrn+mr18cCz1o0iTeBWJd5Uo8kxMcoXJ1
be46VpZ7o5V5xiPvIdOnZhsq+QYO1cYMlAsBpGJODaVRMbnZVz4LCZw8Jd5E
Of6az2Leq78xub0q5zNPSECN1OJJeYc4m1zs9OxB/82Gmw+oSxuGz0TgXzhK
LE1CeWQFDk6j8KasFe/Ped7dHtmiieCmImV41xsxhP8DEJLmD330rlp48QHJ
p3FFPgYh4W6NodfCcLwTdVQjDcJ+AvexKojF6znWAcaA7NAg4pMXult42VzX
IPeMLjQGt6/KixbMQWiFijuv/D/YDEKvFOyriJtoWdB1ne6MkYm4pbTTQrOW
V52CLir4k4DD9U9DaD9/mufRVkvHRCDjD2o2EOvYIUsWCmhA3EryQUvRGq1i
nHfHBJbp9gPHN5PYJtet43kqAVRdx5tXU7S4HuBMjwPaGJjN8G8zHOmWJ2yH
o08qAmRZ4TcZRM3i6u30h38kKDPkwRwkBTg/YtTc5ZAouXlS3PxVcj6WfqeC
kEqXnb51Jq+479r0fPqw9dre6DamR5QYuSJ3tAJbqebw3z/pS0MC/l7lOPTS
h68wHErzPm9vwqahxl5ByKGBmdPWccgBgYEFxijwvjI2nuXaC8Dwyf0S552e
td1fXFyFHErhrrbdtgaCusu30QQoI5MWc48nw5TnTuJzSiyaZTCnnzzFxDuK
N2o8eSzlf+JUSjVWH+omaQE7IEkF6u1OQCNNC29adAUlIhaZZM68P0sNKBvb
RBq4zdrOO4sH6Ny/9c9zTWHrz9y6py6FCWt+MOrXHGpc0xrfLxJf/M/yk0sM
50iWUmYTpsd9HNdaA9+J6MzQoCGE/QMEEU8mxRm1up/kwHYDnEFlpaAoTC9N
/Ju/1YcpryhfhOY3tETaEDWIhdKOLb+YRlNLtxivQJoksFjyuNXO5XPSr/YG
xVA742sKFTR/lKHQYx002RfNQMLO9ah5LMXEo0dp8Izy1USAvyuOS25+M2J4
4e+1WSYdbdz1+Gbxuq3maC7z/JN2XN863ZH/bMaf9782HsiSioKhnYbPqxqX
H1oR1j4LyVZVfNFcrPtYd6iZEJpa91L9Wh7I8cIhbZVL3wRWpGxp7r5Fd5rG
3OYxw70uMTKUILBCqK2kuRIj5wXUhWzxK4blWsFOVSJAsoNgVVZ2YFQeKAJQ
Hq/kSxqnARIj8S79VO8tqNKfEzZoVCMJ4RKv8lvLsYEdfn149SUMeCnN8f5x
A6YIzwF3t2ny5QR/vnfS57MSQlO/eOoXM2BlF7tutf7vNloLwQLsQh9XN+yd
Tb1zTiG+gz9bEgRRZa4PWecBg2oYpGLJYpI8p3uEk5V3J5VO7nyISs64Kdcs
TGrp1wiLaPKL9vz7IlYFFuQBRgKsvYkDLgOU/p8WJbYoxQldQWYVKyCvr1SW
FAR7++A+A+NtwlQzEK+2KebvDhhn3t46nX6zQUB2DsWp+6vq7k7i4dcmRzG4
H44b4URU/I9PQJc/rR0+6REs/XQ5Z3yd4/HDQZXDe5nuDbp6nL6AgpZistZC
2E+deZ6MHW2W3iN3Ozz2cgWqA63prEYBq8XrYLduvGiblulzpg0Qs6pUcAUp
XrJXDah0gkaymOD78daU4pp046hmJgIlpKT92CVzGL4pBeFCHRr1ALhYb62q
alpdvJQQqRNwaUin4cvzIoWBEPcemKTrgFrJOuPsbwe3l+U949m7le7nGsTL
w88VKAmX+MovNj5oGAizucQ0DvMVruRzHZ/zAYRw7oUx+LMTGhr/DgPyzfIL
4sosU61ZaCLt3IEkpT2sfqaNQKMNJB8KhCKoIMgP3vQ+rQ5x3mIyPl8i1oNl
ZWgebYmzT1aXQEiA73xuNGss5Cmp/EZqzw7L4z+1RtIL1KG+4/TbrA9hXilZ
d/avy8PQOz1/l2cdshQMTPzOO8RPi2T9+iNBiPVZJc+WcC/f3qhb/fXsnk1D
FtCUmb7GmwnfnLqnKlJk5wiW0WPXn/JPT1/IuAkGR31G4ssk9soiEdTMiqV0
z/O9vaJQ6OBo+DJSy7P8BC3p+8mkMdMf/P8HxVxQCjgcAuGi9BuUOcSG2mT+
OwIwvoWLTLKjdDQzSE07eeisoUPOu/fjFrSrLBoIRsBUOPQQz0piU8kNN8HM
/f9q00rZu6rlGPilKZc10rLt7rg3FFBUArM8bS+jdnYXYBxicDx2+jflCjGV
WFQjLvrG5/7Jswvxc5oHYz7Xsj9paYJmPP/zSjVWanrELjAdHOcE5b4+iNc3
E1uwe/0SIeuSVG5l2h2QFi4KmW9Yg4tWdEsahRjbYkJkB9qUfFTtAuJ2ONSa
TkNSgEwkbPlzLTz1iyxnQu1U2i1tj4QEPFnKRPfbC9aGmtGpZptG0YRPGhum
0AdwOoTctQH4++zdThfv3RD7s5waLMIVp5RA80hCvAxKozuaVdPzcHK1yLy0
Ya1Y+XQlEqxLzkYnMDGkfGUWALPBjDJDProVs3T/JRtBQTIMpZfntwurOb8Z
rmWDwM0ATRC02SWzrL2h2c2xgdxR3991isyxvas+m+HLIOCi4Ebsytfy1xIP
1jFyGawFProQEqovF+QPVnT3n54K8gIzOaYnZtyPc3WPB90a8s0p8CXFpQjI
osZXWdMkAcbmeEX+H6oDjPK/zLpooIdSfsFWl9Tvkfm/Kkl9M9073ZNURe+S
YvC4+hRcZoPmESBvT7Yk/wS9MxkqLOE4KJMerOE+6auzIZxDvVvoWjgr99sV
9bG2ZADVFY684Z+clTi2zKpZCxh1mOlD8shfX15nh37Nf2m0K00akeo8HZDL
3aE/3qRqv4VHDhuWjown38PKo4nng6KOAC3Tp5wBpBo6S2vG0BgE+FSq4rW/
Hcknqzof3r21zTJb7/eD1NjqmS3VjH5QasDenjJcwf/e4cF9r1uNwT1bOPmH
pVoIHPZSikm5ERWj9i3IIKf2iDygrWtIGRF2LNfIiKiUhm5vGUW0dj7lq3NZ
rM0NTqEH+jrViIybvM3fQjEcnOnx/5UuNfQ42zuPtzG+IU8WoXFUEFEuzRxX
oUfOHrkMMWUFAheMaen4tQrMvhY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KSvMUSaIivcQZwztNws1Eck+zT8GN/dRNmNm1fZRBhapUs62v/Zn9RIWZWxiMlpIBrsnfoXgTGJj13OtOqeKYEWbUTRLV0sOFVlgOctjGhb1qNe2WA5EdjgyNypH68sc9HqjJWR3PZY/KvwKsus7EF7kWtCyd98GwXyuBdaDoiXfKlqTlgJMjOwsWQZRRRmoDqMf4stYiRzsued0Pv5ue3OaajvmDUynZsbWhvVBdBbQE4d6uJ1nWr/OaVQQEcPVsXx7vZ+1f6hPN6/yOCSgOVzDWHuqd43FNW8LUoKLEhi/uGSVxHFSMRJNsxSFaPyx1NDZC129pX29KCdyre4WdbSlOXmQL6qR7p0bEfAfkIEYCRRHnpdMhh96KbE2GuAdrqFQN5+zkHyp2AYHMsoJWhNjqTpz0N7odq8IRJgz9g98b/8+tuJYbXDiSU1O6YbJjaMeSW8hw2jXC2BuMyDkFIHV7jX5bVSbsp40pUSk3ZEGbTOWSZCKQXo0GSE5qKEng6z5Hg6nyhN2Srn/5RSMw87SCJ6oBuhUXGNsnY2MxU9bGvQSeDAzNCN+BRnjTiP/VNlVT72IncH+gAFBTeqiFQmDP8ux9ERlm0fv6b7ropooe3TzF0psU+yTzl2KU3mLewYHgjgrTVBwssiymdU9iih0Q7Tf3j0Lb61P6bs8tMPWJNYM0M96PJII31gLSvKuegvjyYWRhiWpj02g6MCF0Ax3mBVFtJvL/fs8q6voefkd/3M1+GaQ0JeVp1bkzBzkKRw0uXec/MICbrpqKKZgdl"
`endif