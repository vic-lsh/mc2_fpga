// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jCtcM6BHWLeBYLselojI2YyjdnCZe/EhAcl5vZZIAAEb8bzz7JGs7T9RrLLS
bkQfvZD9rICOSHg6bRF8pNRrJC6KGTLFxDVS9NjTpwQhoiVaFqhIdUDl05C9
DY0fBQxXFzWZ5BYyjhMTgR2SGGnrMzmtmKZJb79oRbHMPklEPzLyBZK+Zgzs
NXAyU/MZh375cyyuNVG4J3HIJmmBxhTjv8JHF7wW8UbTv9SZsaKNWB+MQyZi
mDal2J5BYoaQHhTmpC8lPud+QCxln382oaWz4rJVYgVLhUpVYSmCHLydnl0f
L4PZxTsSeX+CN1shyf5S3xDhFuF6OWldXzk5yfgCxQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OrWTMPhTMqbJ7LK+mJJzqpOV692W0Ay3WOMx/7qpKYd0tPcDIzHNLjSHngR+
yeC1W4oJFfi7ToXE/OIeoIawDyJ5VXwFPt/5RkwpPRBZ6aPbGLteAf4V+AyP
UqMOMAKO3nLifzH0gsIGDduF+/zVBQqoYGNqmGqpvGK2KH3O7MfoFmQ9ThSo
KXWQBBewgOYOyD5VCz4sXtaCVL9mv3Zt3yyYsuKF9RHmxoGe3undKOKm9pIN
HozJSGTt1TS03LtgT1H7FgxtajoY9JhfbGd7UlkZrUu0v8zgIpn4kE63BPjJ
U/zRY53NV0O0kJUogut2oLHknk0KcthBhw/2MrajwA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Wcpw2VFxgqqR5+OZ82Ed96/AiIWEzqsKIgkA/aF2JAgWo4AOuXZ8+amOHj1H
L+8FBBryuQvFHceNUmgwyb8zG6sohezUBFxt+96/LEJi/7ZQSkd+6s6011wK
3Invqd4fFkmMNYun3DCT0NFdxeZO0OsxeFkco34Zo7NHkLiYuA8+IhsBxUCg
QOTdgEqHo70tG73gymKczEpgcVd4uKp2w+S2uzr8Gy99O6VdigdfwsregI6N
yKCxShugEFRiFiO3opPlx+RgAkN/B2f+EYMrtcZzK4Uuyc7QOiTfRZdN7FhI
1xBR/CIVrilU6ry6cfXSlyor8WJ+Z7E6ZOHh9PB96g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WZCxdxOAEzaffIhZ4bg2hApKrRBuP0c4xNY9Raecefub8630CIG2aPOMG1wh
mpHC+Tw/CL9CtumiOrrtfsHnDQpRfLV0XUUZbLNffwHLTO1LowcsvmbJG8fo
gg17cUAx9wRaW1bsG46g0x3sv+xLgOIEA2NeB2Gv4EHjZ9bx5D7+HIIiofqt
ZMgPqww6DQYm2kR/W4Lopx8V+jUCTFUcuVBx4Rdh/3ti1/i66XugsWSFDKzF
5KWWG0pTZD2AWXfnsCODUWa1PDY02glOJxER/NePvXdcUXAG2p+OQWTYrGrL
OB6intQVf5G5xW666stazsTcqYMaWEY6QvnHJvagiA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gk9QlxSY41ff0rILcVMeS2B6h+py0EMl3+dipDIa7Gc7menmnBKsfHo1DOJh
wqu3SzNB4PLo14W74j5MVHSO6nQniBRQwraWOjcFymJ0WbCfooEGcEmN3JGT
RLhkgUYatoe90suyKi3kTbZ2EgnaCLKE+QoCD+9J05ZP7AYPusU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ihBJfV97P8xy5ePjqOT+MsDQJDdXnRCr7GSm1IXAZ4C5czoIsIAkK2bWdl5T
39OMcZCtZV/0MnsZUtse3JMLpMPmOFUL3kqP/m20YduVSm+0G6DrnminbXFW
KvQju8r7AVsu82z8drM40XFqqovbAfHFVdEMULF78asBS7hMISQCjw/oUeHA
XP/mz6m7jpBO8YATqe9Dx8zGN1KhYda+lVwUsVPvJcTpym8zTuR7F8Yqo5r0
HidKPGR6u0fo8Px8nmEp2JR1+YokVEtezTEXEAZ003+CzsJV0xgq0nnIlHoI
92ICpN891gut3gOZNXMiSS6H3k5z7ZuhYlKjva7F3DKDsdVOcFr/+khUniGP
2euK44HCPz//exBW7npin2LE3KPbYU7mFnbJWxGTjB1jOzcNp/s7RNmtUFm/
3+H1cXN05RFCRrvPkYrGdGu2SxpP418uif+r4vYFGRYWqmnseTsjOOa//5ac
Gx5mLG9gVUgha6JemOJYgY82eclFgP48


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Wzh3ZhH9rvwIWGiQMFN3lxyRukwH3XNR7gW5zogG4JhfI42XlaZ4Om3RPGUw
I74O61QfZaMzt84L2kUu6QazubsQ9U+r/q1XUSu3kh83I1EH8lg1B9nR0Ad0
XwILB+tLbt/2jhKxPdqqkG3xByCTMyfZhBsA1mlOh/teMNzngX0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YIyCVt1O0iy2h+a3mYMm02S6WwE1hlMn6stMrHlAXNt0EK3Fl+xjiJGN5V26
C2pWKbxZWRQrMlfSDc7YYhHsVBrUOYWgvd9jii4M1tT8/R4WuwKQzrb7ndWe
8awcd9zJJc7B5njQGp+P5jpMwQ7BGd6W22MxQJ5ejVOy3isIafM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26592)
`pragma protect data_block
UL3gaDheskKo5ct6S7MS3EzSfOdacHWG27Uylf39RKpkDY5f1lpa4DxgSM6h
U8WQ+93/0SvUwsLgfJ4cbxawX50ZqVY7U1AaMTbVAp3kQDHqoF7LV9P9QA5d
7nPt3pQ6yAPyp6b3beUQpP2b0IuS/S0N1oyNbQzp16++BDComNgBEZuIR+He
Xyg4Lboe7/W7+AG1gqGC5aiDxk45J5CfFFEXuNvj/smrsaXaufgKC5qbGlYl
1/nrx1VQ4nDmLAl8vv4opGOmXhw805hq00ZbY8PLNs5TpnnLa51Bwoci5sg8
j8AiNu5O0MXhF/H0SiGIWaNCp1zJyuH01SFvpWD3M5a8Q76hBYJ9t6p0ZQU/
Fy6/XXktO2/UN5nLQhjx6vpcOpBZde8F9+nLNBetafOSELKd0/a4p5Vr+Jyx
XXxPI9ijKoQpm1GakKx+T6y54/2u9F+3i66nDfgL72zj+DT39JVdteeFJJXG
iO4NcCA1a92YNBXvBvhQVf312gHBgKgf1Mz4ESM94JzhkJHdNqQp6zfxmTas
aNPMB3SmX58XM5IbGUs4dVUzXYy5SlIzMhUP50ylGlvaOSLpC8AJYPrwd2Bo
rKhZU/q1zqlTPR1RZl/G2Qs1F+yRqv5QwSuF0IXfzNOVG65gUty1T7FcCsbI
sVv7rDu+4wnciDt8fjb3+cK+8zs+iE5zMy59Rsu8X4bRva0iLx0YJjrVhbh8
msijW8zyfPBh9i5WD4Urjy3kx7H34vU+CzG9Pew4nKpT/PVarZ+INSt3V+Wq
+H5vU2d2hWd4/drJSJT2SRhMZmTEoHnSyuxI2k4VKGtr07aZoDcyP1jOwMN6
a+LWV2AiT6ppGXTC7OjUvlNEy+XGYOZDmUVG/EC7LafgluNSx3ZCAkRaSQ+Z
yiHonBes0gtl8SgU6OQgBt/mfyupB/nCccs82UEmmJtmXhSWCcviRTAWHJ1L
CUA8SUFU2lbg+kpWXYN5PeXt+BS8ETsmG90VRE/+W73TiP5ZsbvU8xevC+8d
bs5/7lOHtois4pyzdwaFlG3sABOmyMdGd0JDeTc2cKusRuYIxwMyphk1mTQh
bTFdvRdw2ZcFppj4Qi6QwGQONPMeZlD9JmVE7dz+RcA2oNArRH+7YgwJEMfl
dQDyLrrrdy61URkG+SUk3DHO8ejmhk+iCc2+rvFc29DywttFGjQD0cXTS1Hm
2y50Zy0cu1F5TdbeukXpiXH5ARXLFnOdo29ajD70NpIB0QYAJhv0JzGzkGtH
B7InvOhivo7Gh2l6l9cDL/OTFV8bd0eMVpVN54vYSw2C+R5MEAip+PGFIHK7
JJYHNAGofk2mpdSu/1X5vAyc4wr/9M+64KGdFWowPmB4c4sdgHKMdXjZ6BTY
7Nsd2VJZ/sa6+l6Zrk6oN91WvSReCnpibUTdEBT/jl9GW1mc0JjhnWUCVIMU
zUe+lyUrcDamesLueKf4lCzZozlewFTWYS7BGHFQ8KIpA7XKuFTkmAgijH5r
aGSZftgIFmmWMFiYPjbqtdQrKkol5CtIjkpKoKgjfyCJGRbcyYJV0CmjCSL+
eiJxjeULRdw7PdPBknNo6lwTDPa/WpIGGdN+asngeuPDDNGu03IgEQwl65B+
rx4kAcuHSUbQknPZrBcmZEg3sdWwZvC9DYVD59PE6iTKo9ALzUgRHHxcJ3+m
vTvKjB+OaP+yBY9ELkvaCdKJfb3qgCiotd7mU7qgT03iZiEWjStgYx/x9ky2
dJVbwFpQ4M9tCBIOCisEpDVBkQlaExuDPI2eRAtUergJ7K22VXxMBrs5r0n6
U1NmxCua4x9zwbRqdoWWBj88x3PMtCL2x31nBlGEsZQAT2aGBBFxjRf9XP0r
/iCzWrI1WdNMohrXOox5DQPR3XOwwH4RdRxLkl81n6QNXAfCEulSHjGBv+zB
Hn3syaV6yrkJfG47YrNAyICqR2CEcmM0Ehg7CVZ/KdFigKFNIlwC7AKhcbVr
Y5aHd2OqLSb/6KeqTLANcaIGOZbAFf8GqMPEi84cwDy95fFAVIYYbeW72KiF
3gqobqMJbkBlIkRP39wtTxDkE+xuObBHzreNzzmolJfeeVth1EKmeIFf99/J
kTtqW9r8sZT4PRwJYsdC2qlt/ITOKmG2j5PSt6/mYN6aBXuWzpsMhQkMv/HR
kPVVlSl86y8qXs6gRafDBsFk5fnJFJ92TyM6PvwPo9c2qZmrHZuxWfdu+pOF
3lvmLpf9O4hES1NHWxQkPc6AP48Zw4Qjnas565Sgfa9IKVRUBdV0y6zOkT0W
hgf7C9Oj9t9HK66pnm6CL+XK19M3YbenPCHtl+9DEXo6EPyBvH9z1mHYZSdC
MDx7ma9RyL8hLWHRhn35EqKhcFsVmjFEOQON0qTfkODtFlODVq/19PSCRC71
b+9ZyrNFQ+9ndoRkWh1dHB/R3AYuoRuh2iUgodSJfPyt43thR0oMRT4UCvUB
ERoeLVA5DHfh5x8jc1fdFzRSk4tCK5GNX0Wr3XK0qamemhQV2vp+sVDeoZRz
Cd97mVEyN9JlVf7aMKSiEBvieAH1idXgvF62JuEkZhYBpf/nnA1NSbyLvhxg
v1izyNEmLvcEBMMPmPSFB8CNm2BP1Focdf4QxbNsUKZ8oBeaZ8uUwbtNw6/N
pmiucntbZzv0o0vGDH9eQprxvHWlrn94udCoEOorfZSdFQajJRmy+9M3Pqgv
mJYiiS4gxHfGTGpNCrTiGYXbCYdklqAruHy/u+ba02i2fY4uChA79QY5Rbky
tDg7JL4iFwBGsHzF5vIcMezVBIwmF8MvFCfnxwgcrZXR9NyQxsGRyO7kea13
wyzKHfeFkqvMhUF5htAl14syF/PPVQ+++65+YzKWidCKBWQmQGe6zbIFB+sq
C2MoIg40o+YAkl12xVZpao4qqW2qlVFVG870NFhR/Im3AEFoAXglYUD2zfEE
Up229rRYLuMZCsLihEuAkLpEFg0RMO8ANqtaiLinDNVT9dCL1fYnUda02I20
Rotcto0jGklWueonBn503sO96VwGeIJRczGyw2vqvZfQ6K7m8J3tYwYO6izb
mA7+1rh1IC4cqsZjyz5TZI6WborKKbUmpQsluDioxzi65vib/+Y+wYXvdN7R
eM127EfH0kM8uL8uEvlyAIvxcPcY2CoCTZ8bwgCnFDGBH9MiUmhURHQIqz2p
aV+uyLHNdc+MqOWmPBes6TG2YMHvZu5Nt5s7iDGW5SWcVrDQJLeq9Apu8NTK
aWmrm6F8n2qVEerXR2mmJzlqkSw1bHgv8IP9UPBe32KBwy29qtiIilBR3hOq
49/gcJy8lqiSc+DRHr9oCMPXCDAtGpfWEK8LWgEn+NjlPEHIrD1sBpCiM6j6
VEUs98KmhfvYxp7NPC4jFEoR0NMGdhni/oHKjoNvBPSw3fxrZqqtFsnDvFls
sQbIrZihK6FEi89bSukc13lsOcfGsXBHFaEWtx2u7wRdp/ezmyv3hRJI/W3c
WQCIz8qVwrIL9FWdePtL20Hv9uxn5h9CzTnwZ4tXvkeHv0JWde9MWIl7RXd6
PFdbOcQXKxIG2aTG7H0eRBO92aiXU/1XDEdg7cmBMKWjTAPVIrILjTkDd5Lz
kmema+sB7gN429KpljN7CXB3x5xbTytcsbmJiVdMDD3tNJyOyPW1vD6axQA5
n3Z3Lwf/jg2osQaW2yUnFDSxI2UKJ1lV1ZT+WjuJH7mnb6oHfvWR6QczoPaJ
oEZqligh0ajJbHASPX/mPSZwPw1M/QOWbTH1ONk91+By36hSiJoxd92Jfk6p
4VhBblGMywRLiWgHXanPe/BEykS3OmX7/uMHJAafvjNE7snep77MQamjjCnF
93E69RDiVJj0Iub1t5cp2WbPRwPbQjkCP3aMRkkoq5JjsCga83H/bWwRXPeM
o8XvxAX6KlpYKLgReRuFq0CSAImtqotZ7PhLPCnmuAF/5eBUfNOxShPxkSlX
awiPoRj9Dzs8VGoa8CAaccpneN+KbjMDPuKWc8pdq5s0x75jg6NZ8jkSbLy+
9qRkPs/kxubBVeJmBhFVdfNc4Y013XAmVHjLcHNs9CYvBoNciuv3i4jIapbF
0anDHd2nNq0l1CGRzxk9wWDoZPpqeltQhjAtqh506kZb6YWFH20RSnlOmj0D
sKJJeo4GvvL3p17LiQV1mfQabUniM+F4EZySYSJUK5e6SVIlakYP9erDEw57
kIuCjF3hPXDezsz/FlTaNASxsAlN5t9HSlKFPqTmiK4rq19InYAdaMpjx3R3
058XUqdMrSD0GQUJtbEAHZqu9grgungi/XUXG62CsWRGP7RpdHlR6u2aQ4A4
5s7qDtoZV8ZTMHzmL03+s1bD3bJeatRgcmVfY5ecr0YM/aG6e2RjP24DghnW
dDkW4GPMJk7rf06zrTh/MV8fg+Fe9h0Xf4RdEzMjzUEZBsBn0xbwzcM4pzP0
YZ3mptYnscTs639OdPOi+lJyJzIdQq5AAaofZSGVRzTjUSXtn8OqMSMhFCq8
wB1c+6tVItFJOykF6kQkpL0gViDj2VGVof3Xje5VwBhUsZi+vPmG/6MXX+IW
fKshu6hs/dE+IfDhBfnr+WHOcxEjTuUHydpRB00/uXfs1uhzUTrODv4luAYF
MzR2OOa/dQI3FN3E5yynErwWaRLDOGpOCkRNfqy8kKI2x5ElL19yqwcWfweM
qV08oCpqP4QXK399KnRVFbIsoY6CycZixsyxma5ryWDxSZ4JX0opC/k6Mgil
7PxMA+OWf0HNNCaXpeKwBZfnqQ1msTEufr2ZDJqc73QmsG02c2WO5zT6Q+Hg
K9gq/jdvDH8qi9nLNt7aX+F7He6revHxjq/4wIxy9OAjhpMYKVc1WGWrz4o5
zM4Y7QOVAhnfwZKd4kaoej3cMFANAiJJT/WIfkbgQ0IjD1Vl8mmeJ7rosCvp
vXVY22KExhN8NpBe60C7FbgFrRiW7QLRt0hu+HqdQcJFcdBXXhnB7eysoU1a
rZFt+6iPGWp63kN12PLoARkXVdmQErCHC8XUUQA6bk6trPbhogPmXDA2rjl/
RfC4667k0gV/3KnqQEiGVR3EI8TqWEASZXapUSqIMSE5XFIwnMXNW6KBV6vS
U5pOR5wsuoN1ZUzcVKIKSurUpcbLiyNjfrlwWHenmTIGhT8UA0dOWmyrI8r0
TQf71e4mUX3FIn/sMs7QOhdilIggr5PyqzZczZJOYx+VMMePviXn5AxIzUZq
1UwfjYpevpIlg6NnGRmeb2Tu5OUq0AB2sr/dYKsNBRQc1IZpQnI3r9UC4F2N
9NKQPISzScJSzU7SU+7mwKEphFftqe2t47mhpK7FOWLVf+myCcntryh54OsE
utCFHYSbG/hcTzfv/CgAeBF+4cys0VTgq/Wv9evsqTHkfVAfMRdWtXaWHTsT
ta6/Pyvb2SkJVPhQJP502AyJDKjvh273U9gxZe1P8yrG+G90wL/kYC2E+Vb2
mTFdsjT49PHuqzFSBW/2X3BEwWP5/1Bv4wGh/BRHwOyq1LxvSl03ATvXPwZR
cFv7ARahSuLsYdXdRU8OYiosw+ffV8Ez4OfaeRGq8vXqRxi09D7Zk/GIzB6T
Dgj5cEvXOHzirNBCWKjF0IwrJjndiRe1YFz+RmzleXu3SqYJ59H4ze4RFWLZ
jy5TVKre2+fj5BofzCQDrqB2+oSPMiwUotQwhWFpAH8o/SZmlXYi545nHBLb
kbj0RqCRbATyWfSsLHxQybOSnqFC7MWf5ic9iHQ+UZ17DH0bNOpVhKcsIyWU
JPf3WD58Ar9byzjR5BAP0wBdkJsnCEwUXH7pXGv8o9/rAJy+4cgqdghUKGd5
4CWCxcJBTSz7mOKJaDcdZHdmlwtVCUfyz/1Ya2A7lHsCkgzdsTuv3yDCN/gU
NFv8+vJnxF0OMzDvxE9VwZlodTpPgTcM/ydCTvyYOsxHwhnkn6neebIy/5gG
sMkVe/RYEIiQjFqSmR0T6NBkIQIHzVkQcxHeJq9+mp9OgMBvlIt4QRAHmWlC
TcE1I4QPD9VGXpfm0iIGblSn3xdePYLvgSBzWVo4zwaDefZDr6XnHfsVpoCI
ptzy5SuANh4c1lokxcpLed5zqvdL9cSEx4bzoauxGjILjcGKlcnWbqQwUdqw
vtDNvsLN//QisVk1xkOfZeYnJ8ru/gxm3vzM35s5A/gsBbiIOwe0dukY4M6H
WHwAsZSdD50ROS2us4rOLUeLt7w4h1y1UrzqUHZH0g+PKIVE76RuOzyxO57C
d3+gEArG+f1HgDgiGy9MbmuYkmtkSqyWGMWjbyLnvbGKl8gDAEt3wwynS18P
S5xlVW/Q9yLATtp47UEhWFzlxrHktA3mK6s5VPZNZ/I8lSiyTW3gaNf3UzwL
VnIqRj0Wmecj1F02m7x7y41Ow+QAE/QZNzvoaWSAiOuIMiOJHXnDeX+akllo
fZwazxsvf/HLokJK+8jQUu+LYvRcH5aENFGduaFuyDeQgWbUqxzoVXU8o205
QsZVWTCv+9Gl/VLYSYxB1GbWcCJXng985Z5jFlnWEuKTxZl+ijLr+65uD+ZN
Dz/Q9bwAFvO4cHZdg/Vp6MTVXecKKMQfrSNZXwhnMMkRn+lbNp3OeK9pNDL6
JkI/BYOqS/2+ahkJOzVA/4xevdWzbvk6L4h2qmhTCX7BlauEJPPYwoH021bz
oz68vRbZZoXtUATsM0HfQzHtFIK0qNuM2ykGx1a/8uEsgci6cbrX8IpM2bBD
OsB4q/q/yVoLNn1a8tZo3EaR0SnUeCqgCdFVjS5V6Y+2mI4CFpbjaAbApMNy
QqUh4l22QXXwtwqpduPVJgeUwOOBjsUrihjFgAzcMO7In0WIRmb10J6Z+e8p
Rj0+hM52fkGB1P11kwqAW3sY2qIVssZt9Zv2vWLi7afOn5RkaJ0iGogb53mx
Vy+02KX9+VbqEq33Dkbux03Me+N9O4H5tiZeMtLYVoDHPuXfBvZWz1pYD570
k2ThmezDUiyJbLd9WVZLqGecE0EKsROpZtetTljoqmofbJKU3hxJgTiDaSLm
j5DyqbW9gWJEMusbYCaEgp4WyTdyZ6d7fB2fXwCJu1AvJTxFJ/fmVk4iVUPS
pt4bQh3QuOVeHdmmSuhHtnPrFFs3E0ug06bVvh5JnGvZ/uA12bgP78SPCezt
kr40Gbr10gEaEAyP+5tUANK3MLRpwxsRKy00S8esM9vyAO3XhsglIEa0fjs3
OXcLeL3qNdgqifL8hwlhVn1qgMNmK+yCUKynsfSOCQPhxkFwuKXOB6VpyW/I
0ImhdS5ugKeD8KZU70UU66qzd4hMoSGUZ+Q9u3/DnrVFWdhgck6lpBXsY6io
01lz0jBRcWDJhC7oFIqaOGLCXzunJPtb9TeeK2GPSSzxgk9tC2JMu0GAW8gj
vqfJyyPcYG28vx//NNSp64lxD10LzgqMfWOmmrFCFcNEwnq6SqRn5Cj/uHNy
zsztkQraQ4/lWnAnNP5QftTVILKQon9Ze4b+L6znob2bY9OZOIKP8lnoq+Nr
z+rpkO4ovAiuwx2qVQamwAJ8F1yEeD7hgRY62zyfiUORS+Ip2BEthpU/bQVU
jPS04B5+5vvoBjo7S2ZoY2mrLUzFTDz/Uo1RL3tSXYnRmw0Ss+6a7eaN/BlZ
/O5SKzZJ5MVi3G3UItieg2eMkGarGEpRPEZkBy/aqgwU/kaqQ+JNWFm/tQS0
YdEDy9mtleO5j1NgkFjuiOtyscH9Qbn8zLQ1GpGJf5GhSkrgy/9LVjVHMy8B
A5fOGbqOFTxQCJoMviRarCJ/n49XzG64DT3AMUmCjPUBp7pnmwv+wAiqtQ4b
g+w/hqESiL9Cn8TA41rUCIhHtG1aNLb1YwIldwuUN1d6QIYgcfSo/MpHCeSR
AooieGVHx5t1UyiLN7jFmiEe4r6HfMCLicdFbhph8Cb7/6el+OpEpcM9zWpu
Fquhfmxv1XKFgleIHK+tWvItXn10JAzdeKT73BJhNOER4g/t8ckwP0tbMsLo
nNByUg1vmQKq5bNhw9JUzLCs/XKvJQEGdoNim54bKggJd0x+BoHpYBmU//Wk
/VTidqQ5w71bIrw6qo0CT5g26SR5wGe3sVreNpr5eYdTVm+CGJ9nUlpGx3rW
5z4IMPFKMLH+FUzbuVeJBcJgHWBaMlJNL7uWv1eYXtXGRb6s8T/qvlIBSlno
nd7Cj07wc2xYgVbJpawtJ1jzCFIsupCBZ5YDKNM40fNE17NFvgO/M+lqxaf+
ENIkSqPBUFEpsNAsp0c54Jy8v3nNONFSvBQQYnL6RMhI8CS8Sj2LySlik2DC
TnfjvqrbD48S38OSD0byAZu5k0I3AQjWuCb0OH05RL91yEsplP1JYIWlXqLe
CHu1jCzKNJddD4TjiEpjz0jDOyIzVgykR357NlIUd379h68aOiAK+nF22jLi
GsgoLbnjQ0KOP+LwomajX2wp7wJPqLdxIhwbpWQYglF75u3KWpMWDXnmkR9z
967br7Qg5hXgDmJinEzP55CDhwyt75VuEFxbc1ZCcLwl4x99MAdqmGgPGIeb
tsV0H/uyqxso9t/2UXiOYMt+HHmz+urfIfxXDZ/jLubUHLxZrexDaZySsI3y
7gmRslvzcZmUTovOCDvkhbbzxvvA1jZtvT66EkivVmN4MaFua9u8/DIXeR4b
vO7N4oIkwudrusLrx/wfGpZDU64qstMe6SDhiyz9xy8s9nJUKa5b+6rrKp42
o2mccIUWNxJkCgM9Y2aelDNLp6RrH9oWS6V3TSpo/RRMdozz4L4qZYkF/hzN
e+7RvR8XOIX02Qdwfr5ypoecsTqedKznSWY9heWafBUz9UG4QpL9v5M3suDZ
Mah1I5GNi4VWcZwl8IqoJIK8j1TjyblZM/kQ5RUOWwYLEoQ6h6IXVtFvXQNd
tq432l+YczG+Xui1Q+EjIJsx4ax8Rh8GVc3vZB38jJaWVhC/SobRjsdeeu+n
OVSn5pl2GGn/0XxfSywZf/zEgVCQSsRRNY34TR1LpDO179mHjgUV392Puu7N
FBic0A5fqmt90L095qruawZ3CBV3JLDWPNWHKTJQqC2tg0dHIAlJ2XVFgZmz
avoZZFBXdAueFkprRRupiZhGda0gz1sRlSzap0iwTb+c2mFpVkGeq27jM6SV
t0uoaD0knhUs//0FDLuKFSu6h3bylW6g309VTMvTuv6w7N9SIQ0Xo64A1+4P
ojyIu6KOby5Ha3rzTj9SeYjwLRU8HLJqCUkhvvxDSj7qrKWQ09SAcP90sHHR
1xqq5UZ1HfEv3M7y12tjY6w1+zqiyvX9jWYisnzhl1rDnRaFVOK9KkloOaUs
q8hJNY0GydeLqq2ByNBc7rRzkQHKovZ8iTIQtyQj6k3RAEpiXwV+zSvTUw8H
M+0YXXqHd1ch3uYaGUMk4sIOzsMXpIo8reK50Q0Y8IrBFckb7wdI3p/IyHza
QTVyMxEhOaGEjFCbL6aoUSwQuufGv9saHPiahw8vqcijRa3QahBidKLaJJw5
/bxZh8U/QER2BJa2N07Qd+LthwdppgIU+qjj0ggeWRQmXbRjwUbmnwVXj+O8
sSCFWtF3ApzpdDUW/6pebPHuHndBTZ4Z0Vn17a4dBE75TZ2yt0FtagOMU0JL
x0TvkH8anXVi5kJhrUxwI6E95TFHQMJRT6l/s0u/pJHkCP5+krCNsHivVw61
vR5njzSRnCCtfnfJfz6OCu/TJonvPrKzjZFfPWrf0mTjPn2UHC4eAXLNtT/Z
2MQ0m8sV+a/FYnriCy7N35YNBOBfm6Qkfk219wdRunACA9PaL976+e+vCPKR
j0l9Qs9DbN5zleeZq95P0qW5+IDcot4MozNgjbP5tUSQ5V9aV3/X0M/A2aeC
QCqeDr300QTkuWLvug0poa1xVqxB+3W0Ywmpc2I+oNNNx2z8VfrkyVHo+2iM
HrepN670ivW2TQ4W0/BxtVquJgxHQ97nhWYIN59CZRPTSxINSr9HlWKUMns5
I/x5a79Fy5oOWgzjRpF5OZElkBbcfa/JHJtD4JGYrkLXnjLcgBq1Msk08JGd
AmBPArRhneZt//vQGnT4NRpPENKNWhux3WyzEkpLric6WFZofYD0jhl09ET7
xnRmVgWoyy+UCXXvBkbnV3DJqQ3FrAgOhw5sP9v+By2PBXrm8lBT0tCykVxS
6kzF2SiRAf2z7hwiQTEzWwdpYEJTTQGM/rvS3k90g+h/KLa80hOLnetgueY0
mqq2PORIjUA3NCoIEEcIggASHsdXn/6qLoUeeWNo6ReHgurk9KYldvEaYwzU
42xa7SN4pA7HAN8HxRpEJvtWTXLTWcARzi9Su9lUkQuP6L0ShdD42r7qUTG7
KjSO+RedxHBe/JNS59u73LzyZb+PpcT5pq8h40ejbY9EzSyQ6Zm1Slklwhbq
vRGyj/zicZ8+RcBm9eDFZm16uHS4hok2Tw0anCRJWL6bpVUOKHb+Sq4iriIo
OuO+dqRCR0tB/moqJFUgLn1K8nwGzEILsTF4WfNb/o5XJ/ERsWl+fPzrLc90
zGuYIokdAMMAunNu8MwQjTfQ0pRdcSpHN9gDobqyAW91h7QKzN8DuzZhIZfP
55S+ypa5Q7xdZBQF6WMXlhlT0SGt+mZhlnWwJm0gdxcM/63WUGcsUuh2uUPa
4QLR1ZOMDaaZRy50lQ1UVND3c7ZGIS5BYL730c9H/Veg+OXwaGI1X12vjRLY
N/tV5cv1+/BeQXYnYvxBT9S9/bT7ztSt/Qh+y/uZKi1oXGz5vkSc9x66mLMm
c2hGvbspOsjgleBX/CSqpMtPmiRzSWgtCcKFH/ZSDDaGBEZoJFA7rMKrqU+A
8qHsIYaSmd0yMI0ccenuDmedS72N+Hmt29Q//UDWa7h+H0vtJEAuSR8BVfAr
AXAPfxNTSz1XlKBowJ1Wh9C1eEPh3vcEWx3Ku8n1tCisFs6L/6FY6Uc/vptY
SIwLfJd2zLL3szyNEfjBfIsN5UcEg970vMhyVxGRgbQq1ZlPxVPPbgc7xFbo
ZA7NDJaFTRlJp2Q8n2u3vgkV92QudWJrrcboMTgCepVHtORgMIqT9Nk7SVXR
gG0SacKhQDvuDDY9J0hqstIs4ZAwpUeU0QbQnq98yPbiCIAb/Zf60nlkFuIv
HripBfP24/AYx440LmCEX32+GCHgvKbX/SVY1HbOdw2EqjY80ZT2WsLfu/8V
cCzJM6pWVBHJ6hjDB5Rdpk3Y9fK+bx7QZ4IX7/nC24La156ET3oQ97DAiwBm
DXqctMRzm5XMQT+oN3OTRSDLczWECqPlPIgerkIK+9To3zlhP+SRTR2cw/+6
uKnprIgqD1E3YXAXJD9zx6Mvb2oiPQd/Ly5j/fXnkuC0+wIFVrJJHoIMV8Wt
9n3VqaWahYUSLO/E7LOE8UVkrBtt0YXzdvB90x12viJbrOc9vWOPLFnk7VHC
h6AfP9LSHGjDv/hLK9D+KokpWPtHphsU6fHK5qZpCckeXOLALTgL1KUpCy2p
wRrmS9VPHHNXsSGvVFXtKddjNyOnqYwcoiQJHjGcApCAaBtSp5IE1i86ipJt
47pPhASYHWv6sZNd5poaf7KfXzaOeUyLXe4/F6eRvWRSl730JSFlB1AMMq8/
SP4oxAnuPcjeKOeJqe4VT2e7omOWU5oKVH8Y/v3U+TQVDbn0sQK5hFbfLAlk
d8gj4cFEjulISx8rdpcKcIBzbbJOklp2GcX6nc/sP+EQ82J+Gr3pnfHFp8hn
MJGpqv08JXX1yvCLXT/5iIvAtE9KznRo2wT95u+WmxZ8o2Ge71nbVkh5/fjk
krbbX3ciJhtrBihjxjH/EjzOFHgVZBIvgH+1wK0YPlpL/S9yJslWU2+tN/5p
vpfldzc+teOgxoyLl3bve3VuvVXIEqiRzwX8FUf68P+9iGbh7fUeKPnMa6Y3
GOUtaYyRThYLiALXf/Pw+AIiVKJCGdTrMMJKlOJY44yuWHJt5Y3JscPv8ACc
gOuPCZuLiBbgmQIqEp5aaCRl4Xr8IxPxapnTWdN30z2JrnOxkMwc6Zzk8MKq
1zWvmmjmhiBK7uA452grXoysa4eGoNKo5lPb3Ato7vh9iU/vRJPYggQ94m8R
D/jYww0oV9TDJRTf78dpUjKVv8Yv4TD5dLc4CDSsBLJNJsUEkWvgdbl6DFT9
LR8LIwSCyccPllDPxOP8sIxgp+RAkYACEulwxzvdqyBVeLin3XfN4iuB1wwz
0AoF3skpdCATAMLLg1fL6weDLWWpiQE5LI6izrgGdk49sv5nvBhKHA6cMTTj
IVNcyfpHt+I81ShMUJ5H2WQS9fhxgDrpSDspX05ycgAm3GnsdvfziGYCc7AY
73EtnmTtKWKeA1nAnpQy+Re2SsmGx3ZYkJYilP9N3SC6iaxhOjrK6JOJ5i94
ouwyRE82FuceNP4fq7j57gikXYind87yoOkuwiWx7GNnM6bjRjjo7a3Y4YRB
jZcedkrNzqDFKf1UuvBYTBbPp4Ymx5hg3xiQcy6nbbLb/rsi5AwWSd2TEW9n
KC8xaJW5Qe8Szs6AjKMu/v2/gTHDRJKOQ4JzYaNpRgomgtVq2whGOMkovH52
z+IAq8ozDVqWv3/HOBqp8UeWUSAADNLMTKlltgsvWZWfHF9g227/elVVAuxD
ozBmyZfqC0TrHG6tsSEO6ffO3eRSI3ERZ3xFgOcJfXu4A8KFz9D8D/BFz5S7
vTKQwY2BrB51OmkU1TXARxEKmf3WnaRc4EUtWDhPT/xZLGqgc3qGDr3X5dBh
R+K0nnOgb0bXNHsyAYOoQQ4v6k33iv3zAktp3y88hc+GXe0rOseS52fepDSi
bazIdnCYTcmGRprFt55pwWVS2WuzR9XwWSjB/eei2AccVeknZmv+A8aK/RoP
7kTyR7Krj5dr/mt0Y/pudp4kEBijQsFgED1LNMfhBwHe2+zWZeP2f6HPKZ32
cwUpR6SUFxj0lfm1snnhAvQZMaMS3Lwqv6LAo/jQqJh6TURcZyximOyaIHnq
OTSVN+Nnzb0l3eszS2WerDD7zAhGdMnKZmAjqExgfDMoQRpFrzuPAPl+d3Ye
6AakSKlGLSBpG53iqUXiy4pEYZwtGRjWVMuqhsu26YvJh1K+HotIczj8KYJ4
DyOGK+qtGdlCTiuDD07UwaL4qCU2CLlTkr5yIWuhUl5hOTFfRBbG6P7n06Fk
1x+jSvl0RfL/dnpNcsR1I3WxIssKcbXnfThMRqo46/6mMvvzIQCcAL39Oi/5
6AODS2mMuvT3xt0eeWKFAMpk9sVydUwDfD4GaKSC6ikP3bU2PV+X7zFIkcjb
qjWQKW+psCeGRxIlYqpS+XW4phCRBUzSvrjd3bKZR6Av8nZvkYfGtwII8AS3
ZFbQlAhJcRenGKdgP99hbbP6YtwC4BwqH7haaRXiADpHCBKTFrvbFbZq6U99
Fp/gSKXq/lEp1c44jCtsUI5yNgCo82GLgag75ro69uqc5mJBombyQXhUpyT9
HbxjLbGfjE8LnVHJWWhAfKDUrr67zLiks9MfOoVTgv/oOdwZt9EH5DpItliO
BiiUUyWCZGTkCu3sd+xTIfCn4OYdNKrDoVGi1B8r8mlnSnMAEIN2hCjNMlFi
nOISFncpondBOc0vRpj2/IOeCf2ucQiZlhCvnP+Mncq6giylJBm3r4fMthid
5RLtwIOFymwKp8H7HfjoluU7+9WytLo1NsVOXuHMhsuGzkV5lOKKw1zAqZBa
0bwobe2Pw6qPZJXQX2wzdi6Wj28LqYTBhlG3UYV2ibWa22ECCqCN8D4dCtAS
1hw5v9HB9gGI576d2c+Vvw2PtynGoZvogYA9kbPEV54qeBHiTLO+6h+Jw8Xu
l6B30hNxOHuLv5dkJsormxVSJ0i+UZJj+eASHqX0NETeRDZ26uPJvuK9NfVP
u8zyIxi1GHyLVQH/98SwRCb/GpRatW7EZJvskAC3V56qVqguGeZ6KADZbyX3
M+UaRRYMZwckZbYftxKnI/KJ49d4gpe0R5aFNrs03aF315k7+HRGg5sYKJU8
aHTm79lj/PVrWLKfQIGzcU8+sIlWYFhyXx2gYR/V0XqOxHcg6FmXrasWkbaD
lQpOFYVI5UhUfrMcYiPzGC/EU0wtP/KzAJp4j22EnLvD3nfVxdF8GWrrIMZ4
P/tp6m1EYKUyDZOAbot9L4AGn29b0F5sj5KocCRCkE03XAiS5MyvgcQQoTJB
A9rgMjiafqO/Hfj+O4ryq3fHxmXSyG44aaim6iaHKs0ar3oxfkQSZawUj5Km
WqB8XheRy0vTGJr8O0/Yi9VWiV0c68KYNaO3kJZF1hAuAGSe6gw3/N/jX4hX
4oaSV41XENoUvXzC2ZLkMmwc3IojAU3gpY68y6sHfKtEhlOgumHaVXHbMbXr
OhTVn41X2fLcd/pEgvdxnXZoYDV+qH1ZVCrtK3bZsbFzgUQJGap33d/k6AA2
ckK+Bv+ZXBsRoIgR9+JGPDdbi0+8cEzlp9S89s2yqNncGxLS28bnanVpPAhA
hmfHMwxueMpDObagYKRdvuNBliiwiiKWPgE5FFdhwXxUFdHnDjC8QozbHlmb
4FwPyi1xs3jaYUUTPaUoV3NGWEFNLgN0bssAJCF4sj1eE1ZK47UQCSEIstF+
ULZsSFZe71j8TPnRUi1H/B5qv6pondimBiZwiqZt9/f9etx+2UjUK4lZeKl1
wk2IWoWWQqXJGmJ/nwFcnHDtV/iQ2RQ112ZTxV7PsSszkOKoN8BQpsX/WIQL
DLAiB4h7poslNJlMszTqtXSJfjSd7Wvu/Rfqf5GrDbF7exjJxwwV+jExJ+FQ
VXpEuUDmKEBgeIz78wk0nxHLemgnfL/ASRyJH3yhvJadN22DuQt1udXDJzIT
KNOjfJ1VFsWsEgKA7LxaP445q6eWv2Wz6AvJ8PPqMEXKbYowOir2rS9/5kOc
afHgxyYlcLpCiYXunde0SrNP0oX5ViZagQGjRKtSvHHMP0h4pXLQ6B0MLdVc
BIL+Bf11/G4Ijr5HYh3T/+ncox7yWOG4/MOOZ5a3R9N7tktIFBqxHyxe2gWH
WIelx4GVZjd8LLj6H6y31RKZullsXKMz+ctAEm7+xXWUCobr3H6VHIKQozlN
bfxkknEONhg3zGCQlryNNTrjinhngSseNgLX1ok+A/PBIBrIZEIUTtldEm6R
O/zGpudlj1iQDrkBfcUO+EoaAy6BdU2gQZSIgxO+3rKbfgZLAaDOCsAzBrVi
vkzS6PRkPkFwQDY+36hq174na9hnGG/dgDM7hMrgrLqIyjyxbWp4Olgnqc3A
KJEn+0UgVcW4y7AcJp20KHEEj70On4uBhEVBXINnIgViYqXC7pkT7iDIhtMj
GNRZvjU02wewQaYAfYvR2BxRsyBXf5Zhdx+YQxeVy5o/Ki6+pmd5pzj8/qMi
U11500Gi3LOJqQCSf+wkGSelGCksbfb9h9C2+QbhW/z1cyOpMkpjk5FhrdqU
xUrp/MGoPJs6OOTJzXzokojcGLmUz3FghYSEkBywLkgoQbHDV4aWDWe8ae9r
IlJSLDlBLhSyeJGCuVTWaOcJKp79funGGClSbW96hAHaGuDwodYt0eHM2Dnt
qHU6WuWP/mvH3i4rih0fw85R1SWshblzuTB39SYXmxTm8ITXKeBKBhQeXbHN
w7H2k1Z28La/DUGTLfBjMSsuoGP4CgbNHDSv4oAVqQh+tD2A3wGrxu7ZYAOp
J4jZlVJCSgXAcyN0E5V+Zqh1+I9tocDS+5c+GICfyaqFBLeMg9yPEP6v8ekh
8WbQI7aNu/1Z4DWwiIi5OkXn6ahsoUtZisPT6Jbm7MKVziKBfZcAXgwPAwoj
uGaE7fiiqgTcf3SEGr9zdFxTyie5vyiVIMLHXNZnwheh8TD1RuY/sxMYPYl6
fB8Dy0MFOl0GLMtDLa2kKD6D6ZDutXoNx5IGN5eGGuK/tHjs2TyO02wFdMko
Yi71ejAkjnge4jNay8GC9zK6escf6A1AATYjjF0r5H7wWaVItv1mdHGgL8t5
7YP07ZOAUiGlOUSwbNtKGZNRVard4CYL3hjmDvCryrdB9oo12cavfrPfOkI8
hTVbFCSpZB5BOz74IDHXhU93MttZuM3nBCuKv1JVN7eG3mopfUgM7kAvPET1
ND+CSJ0DPxgwplOU1CfD4mluTSk3WK/4givZSQUvAxBwTv35DWNM3E+3frkh
E24QqOtr/6SUqxkSWyT1piRTmYLugzLrNGl5+jj8gc9KUnrLIvyT0wCByGVw
9AaIhu0ug+AOuRkzXtrni3YGsamWQwhWc1wrL/QkPUIa7f2iEjUgkGnzAeeR
tl+AW1CSLPXcnZWzXNZYDOAE7dmO9UVnRFoqj5SwwsTDaL7Um1EDZB/qyclt
lPPpPFv5C+mVohNf1ZmBcxxOfGMu+CW53qY+pRvk0S/nRsdBSoysN4UOA09c
lhvbdurWHs46BZR67Q2BlAmBbQLpkg2OG+guDNVOkj9884ba6nMN1i0I8Cje
SLuwTNXh/XkmLiVwV8TWfvmYlSKiZs87UvzIhCpuBtRSaADQLRMqwM4U3Jf7
k6PlkoaRdeBh1dzyjKKQA6zAKUmNd9LRLVbsO4yKW2FSR/3c5+4Fi49DGS1L
h9Fl9BGN8EYoF41y1nJQR0IwkHnuUD7j+69gjDWjA+4Cfa0UVPXinJM/dhpT
Xaxj3giATAGqoDUXINqiy8ZO7rLfHz2lEJetSKJgNNC/T2rZXaCq4Q2yDk5y
WPjq7rvi4orSBS9GEP8BDU47tbPNv1BI8Ok7oPfCHRtPYSU725i6JV3KHmGk
cCJK3aY+9Lug+AK5DizPllYoLjKEMzHbSSaQdXCFZOjujxvWuG2tA0+bBME6
JPP5lguAFH7ShN9JjI1JjDVhgpmVZPS9GChVFUCVGq3os1l2g0ilFnY1bshW
eLR9VbxK1TaDicFVk8iajCAhClrh6iENkDxNC6SpDB7e/avHe3k6yNY961vD
hjSHGnI64q95BZ8V+nnWpM9wW6Pmj/75V4iaQH/Np0PrGBbIqpX5yiBAeLh9
FfPX8TWAS/q8BIvKCq+ZH0b6O0ors60IJIXDi6eQiIa0hvjZ0kEIBKvknxOM
AM9yBprCKWF/ZZWT/kbIDSUkJbDXGhCAnUZng25Nm4DDITSUULJXxNT77kj/
3csno/ssFUUWulSu87EROE+1TbWSI+rBuNSM0R1qjkJy3WjYfrsASn7//Ft8
0+dCvWzvXzks6xabPQR/oj98KNQTC6vFMfNfEJWBwrFGKmQMZu3nhb9YU6+W
477f+5m7jq/gspORokK2KCRoZOVfy9zt8O6kYlbPgErv/GZqYab/DNgEH++c
5qiFRF1j3zuL4WUbAVFiOW+aREFLsHgnlO4GvbMzZNGxRSe539FH8Droq4Pj
NSIO7zCEbnMIeNuxYLfDGiHqECr2e6kxsklfV8kp9ccdRVjGy4x4Cw/2k+Uo
iOHWZIrBElVXvdEHZqgEQfkc+Z+5SUAR+C4npgDbC3/b6lfl2CxvwDx+IbU5
4aMCFKUpqWYlT+gbhR9ekV1/NoRDztlmEroJFa3imAu37IN+IRiJaJHzfUYy
NZSW4srqC3jSCxYi6/F/rYf2C9PSKarh7Tj63iytoG7yCo6VW+lNfHAsv0xG
Ux1SHEsF4W3Sw1fwL7Fje0tPzfSfREbn5Jxxi9l43Fk6CZSsgJU7ghVoFUI0
yeg3Kh7yfUj244ZC2WjxmpPhIJY4XqZBdAqbhmdXKsIqmPuNEf7mfYF4L2k/
+Fgu6+3tNfTfBS4VeV3QG/BViKfrx2XhACRASAq2Jj+KVQoGkbwJ0D2StS3R
L2WLKUYPfga+4een4But3yuQxynuOrs48RiQ7cRAfp+qbIp+G3iT9b8hQWeD
OZhFPjtXTYoneL40mL8xKkIz7HprcVOBMxcbl/rV/W0Pjk6LEQVDajTM3XET
KGE64+J//Zuz3IcIfd5hhGcyiAnYB+Ul3zGDA0m5sB3C2idN18TlZzwlU90c
e1Ats3lbwsMH5SUnG425liAElzT2BKJDtgdEUmEzrZQ+ol/252OLaxYVS11l
LJ6z8BqJd/HjfeQd34XdRgEbyjZ4rMl4v1ijCgI1m8UPi3IFV4SwajCwAirr
dgwYMYvXh7I+g2KcCQ/aRMyHNfsCF3Bvs1liutDGbdXV9v+pteUPxfardjK9
pvHlFxMBUG/666rjs95qYNEgcp1ckJTs6od90JuiJ+HguTp6U47ZMmZsCEhq
mAnVuJMt7UNp7sXVkdhT2b/2TdpfvzqqU6kEJEsU9p9+Jms2m0uzJRD9uymp
eQb7nPxCtx/hRVUohW6KLWRXshFv4o6S5Ev0oA8m13F5kx7NwiqyUiW/tgf4
NCxnKWwcthJBWOxlatmHyP1miaqMe+M0YjZXuLAUpbbxSRY/NsV1ST2rZ2pq
RxM9S+dfq1dZ5yph8q+FtKHphvUIeD2wvFHvKjZ6jM6hOTZ8iHx/0Koth6G4
L7fWfLQaGwr5xd2cRvitro+A9FrlgwdtOwj7V8G/uligMmFG3uJXf9ClczSY
XcTmAujQ3e/fZWipYX0k3LUm1c27Fl3o37loXegKjBsvZCkAUlVBVcC/4xhS
aaejSjNFiz8h+OVixF/jFSxa52LLzR5xEhOLW4MTGDSj/dYhBg5fL23z4chT
5gIjqX1rfShZXzRu+Kdbpx32pKIety1SpB9xMVNYIluoVmS70OX88TCXujSr
P1WiQBi6ZjQjWN03AVaJHlfzsmxbpLZTADNPq3vseyArCnqFEXhZBwqBoBV9
QzMZxfrYZCzWN0x5E/LSZPHZwt0OMD0aGHsiA+824MYpo0tXQm+SVf09VYJW
RVjfumj019eLq4gNy6PqjRlSQ6cWlGznNsHGWTMghsM37hBEhgkL1Rh6vhPh
BlO26sBBhXr+HZ/1uNvWfwnnSymyGK3nGEL7j2xq3QVJejDEb23z3Rgu/pnM
ERsarwC1DO2L+cTHvht/XFxBzUqVuojmCNq8AbN/3DcBakL46HSdvkafGtOQ
wD/bdjq32w9SGpkI/nCyImMry1p9nPQaCrYPijMzsV0q4Qr5/czSlgS11DY7
LLurLikjXFudb3vxVm3XAmHhmd7lTX9SM/yldjW0yn3PbOPIl65N+/Nh7Dco
0vVUUfwNHE5buW9E51sRbC+9N7T+wH8otpIwqJsiTqSOjdPgH0GrLTUXqRg9
lMMIK9Fhi4hwT3RpxtzMnr/91SpMkAplGqjvutBwGiik+Zn4v5YWzzsbHe+y
ICGtrtESfzhslcNOpl0DNcNkB3+vHpvbDGvxbOVfkbN7iYgLnoaU9vx+71QE
G5q2snMGMMbPw+olzVhAv1/9fjT9ECNNgx3vOa7m4U1WDM87KaSRBcahWYXr
ZIo9oES/Cvcfq6qSSLP/IIC4DS0RBfrLxMxiQ2UdaRC9fgdOKAvtKTSgmM17
9lfdYlrXuQpMgiMgMfkbOCokRW62F5D5iG4PoJSK1gwHLWAhChx5PIyadgPY
ZQ2yw4eunhliJIJzfRXU6IfcrBv2v8KTIqhhfKhHM5fxvFwH+mo0otxI3kps
5d4BM16ZOJZaZmI0R/tPLk13DWzkxn9H/jbhSOeUMyb7/9hwQQBB5pf7fQ01
/K5H135D2Bymfuocpkr+7BwVzDwHzj/Z4XQ2yHJGEpjoVTQYkyucKBcEICef
GrozmSs9bQHrFIcDFEpeTt+y8u6Uh1IL6Dm3HLG4PsiGUmdd9ROK48wYTIXX
xR11XBR6+pFyc+5ppahDuma9lK9954sXUlxXgxQyxmrnbqaBh9W1mSUiFwpF
a9JtbzILecKKrOumkUVEJVCVAoc032FFIBJxKNzC5+qQP8RXcS7Xjkt9wkl1
UQXieO+O+VQ9DdEWMGD39lkubuNr2nMuJB0nRAOceQHhtg4nsQLlZZRc8tZ+
8ka7ppzxH6iesjM+oL9AUz7Xz3SFu0/ehswcKOTVEeHkzlR8PSLvY1qRC48h
4xDQ/syuj9GNVJhX+YTup0oTTRsJOXx9SFl0fgKaoQkt6/2NzSDKByc8+orU
oNlvrM9vC7h0pJt6R/4SIsOGaKkDYcIMJlD0iotWoWVq6cNqF7DXW/5BHx3H
okpvjqdSXcFTN3W+oHzexb9o/C4zBgtUrTsIYHam+X5Pzhf/Hgl7IFkAeTG8
Lepb4KrNKz2OV4kqry/tEpQwN4G12cEhBKIe+OkSSY5wHOvSFZwMgsVvbCON
cD2jBoBEYSeI8ZC+G5fu8YX/AjUJWDilT7PZdGXm/8KZx7RowmINZf6Nco8B
iB+KMSucLF31RSeecqW6298SO2SsrjlbSGAIT/NpaA/4jzNtKFHH50eRX4ns
7EN/KGIdOK2fMkcoroe35+cKGqfgl08m7HGtpweZNZxA+xQ+U9m5oG0pi5Ak
A4tELR2i4aS96AZ/jeZLJb6S+N+pgrmYPeVZmnquLrVfilrfZl8ypQPbpxp7
Sne1T+NSBcOlMJiMpVVZ+0zJph8OXqf34RjHYzttkxo4CK6SBKlSljwRucmN
4u7I9qJHwNW4Mk/dLkCH11/HhaOoUtMspAEdkJoNstZ5n7eiaAYKNLQLTYxU
4eneFpUYkp7IxAOW2ViBkyVrmfuXJrqq7bhNwIUMIUFMOrLPVBpoLCkxvXTy
k/BeSGFsf6HYlH5uOhZJ3p7/sMneZeCVlQyZa9lJg2C+vaOIJvM7T+ekQTcZ
H9e7ec4XNlof4LUjiJkb5y8c9vjOSAFUcG8rN9lrVxBUyCN1m3UfztgPQa9T
WSo+HQxNqiFitX/4SoHmU6DiwMf28R5aydmz5C8lqgbQWhZ9RC+PUOeHSKZG
24VZS+/g7gcwvEzcsAx8TKJ6t8FvQxuFPhxRodH39FRMdGxQlVLfrOtApm8b
str17wp8FkdpVe5FNgs6vZW+kUgLpHOxrT8hC11+3CkJMJ4JQjAgUqPLvs83
Q8srZuueiWIUomVXV7/7ktfWD6kQ+nd8Hk7nmrM8oT+jAnSkZDJYzb067fB3
wCLv8RaHhIuHubl/dxndSbKmVRVLOhgSbrZ8Jl/EBeYeGQHc7GAA8oG3x17w
nuvTQ7GcKC9/QIV/XuLS5OVOnyMxhjIsmhC0TRbU2poFZS7gdC6Q5lHfK6w6
jVbpg223U3a15Hweb4JZsz1Z0VhGWRd23sfbTxQRTW5Nts4y/Ks7gvKR1f1f
YMf7P7KwL6htPBunhr3EwrlbLz4druVr+EkHMmX1feD2Y34E+OAXstZWlJG+
NO1VGoSOnCrxHbtXOi6XJxBrC4Mw7Z5m5/usL20KxqpLLk4IbdIBHH29KOI2
5W5InuakBqUfSH9XHSEFr+8tFH/z5zZ0NeoZQeRgZS/1ppcJBwsyiTOOV0iX
cK05ZFWWUEQrJIvequY6zjiCdbGphRUNfpEJyXFjZukMH+f0ZaNJz/QchGvB
dOXbNKp1QBI82z2jQisUrZ7mrO2ZsqlNmhClexCYb5TePIk1JvbBorHTOwvS
vzzzGwuN9oaBgpVt1W9J7KaA5wTSwZwVAVyJk9jgbyf963GvtAJNKLtQsSfI
3cmm0m88G9unxUIuWWBcBR67X62qu3VJuMh/e+xxC1yx4TM9AbfbIBJwxJdb
8qzs8hYGwMxU8yNgMlOajTv0rWMVY0fCGY5yADwkCVNg0S70Jl7BhPk3DFj6
hn1PklFiN7N4ttAjKOEkGgucQBFVBl2aSTtSriG1MFgJQlSSDqgchEfW/7tS
/UIgKeJwXg6Ilo5BjPGGhzmPqpgEadcu6x/wHT6lweFuzjzZTUWvDl10KDxb
WzMAjutLYcGK1AIEB0Rkd/hWMLeHXNaUlx0uINuI9zdp6fVCw1hcj2ZAkGcG
PfLeDehuxWeB6suOxqbIMAc7GaNw71ZManbIwUNhs4pAiJLWFYqbK2UoZb9e
d1n9GLnT9p9Vil17pbdeKWhTubZrikFWmqcaLnyExH2TIVnDQm4vXve1bQ2j
ltWz/uzutNYStQM4GSUf0K5KzNEZsWPS1ZpLuDFvEBEHjBWLSMFVcM1i+Iyn
tNyI0KWdmqInrH+LuL4a7P/rcyvdIqlaMGIoLv2iYEKI3M1NaRPuTTfbUaUs
pU1rHMt9UbOAFsC+tOPyLCIAmj3Z6qBekrobwSyV2uxCZuHtq2G3rlVoARxR
vCKpvCgCFKNjI8JLbuPLqkPpubUk11TPlQzNsBO0tCaoSm25vYc+gCSSobAF
gCmtEPKv8wFCDslfFlnvpCkZojPOM4knGVuZk8omCVf/ZxwY5IYhogZv5yLQ
SPr/TqgFcy52ter4nW25iFYSFr4phMnOwssbarRl35DeMfDml3k1PokPzZcO
RjsFWefJVkjvB3Q0MZnCm9pFzs4A+TONyigfyEwrJLKfaj8rdpGNpMkANcL9
69xMTbRbVcLgb7uW8WtdvOWdun8Z+nJ+AQn1xpxSbJc4Yy/SgGRQ0rMwalA7
6VW2X5EqFqlJxZOEvjbXgeyuh4dvUBYMh2liASTG6ozOXRiAHaeBcURXIbO8
Z6OtxlrveLiLzQkfyXI+isi/vOrO/rozf8/MnCxK849nBmZGJ08QKK5OHmef
vAoR+IxVH88PpO+DGGBT1/vxglVPrqPZzpsgaK8uH9kaaaPjuwuWiK2eQWgY
DXNbM56nJL7s7YbXvKRIaIpG3si4BIxjvwuiajqK5MNwt++WkQMrCc/Trzlk
zCZmgTQ5/Yitt4Wp70OLUhjL6c/9u+JXQg3JVzP5pBkSBVtMrUlhQtsPwaX3
qVTPSijGMh+/Gp2W/u6JIzGL//oOIY0GZrh1MPvHnoUOy2qPIrQ3IVoyWRYl
xEb2pC2/kAjmo0qqEXw/p8bH1Qceby+P/VP3dSQGyITHvvlYZ22dxNsjqUjW
SHGWR1pGFsmytnlUvR8J6gsGBraDSX039ME1eX6C6+TEcXBSAk9CZ6jOPoEt
knta5NiF6mFs7hyOxKiqqThxj32p8Ijg8rC//UsZeSQHtx/Vi7xZb2H9VYGi
YgF9KkKITZIIdCWtwoGpO1GK2AtJTflBNMqlNmhnoJfczruEWVlnFgZnSaz9
rmZ7SKrvx8SOYpn9VFfzHPOgbMybY8KY033KqjctT4DAIn0tUF6zkD8Y3lsL
v5wFcE+g+33k9JDYJHKgSRIULyqKX30nrMolQfUZgwutkLcJAGxH4rwwWIFc
hSHMjQ6zMk/MOoEAM247+m66dLmwXt5RJEb4OzoDMS2gWKCYKbaBOzFnGsww
zbkZ0tTDqFSHl8hvCJZ9/XTLgqyfFEc6CDt4PvjbBl/H7JVxFmeKRiLImMDz
CCvKL5ntIGHwOaRSK++KiUkQuXw9CViYahEopYnfxBVLvIXugT6isOZ4NZvP
g+gzyDzFJhrSSpV9C8Us94ERDnRVH9N4XPn16hMSAdETvRGWK/DqNmXc5772
BR5D6kKkxahUEDosWQNb2NLr4GjK0P+ahLSd6vkF/gpMmZRXLHVvuQWY58j+
VmopVpxd9c8uQm62usgV7WTpVRagcv6D2Kij/Abj9/iTUKK4iIv0506so31n
dSs6zfTgnsNbCnu9WObR8s+2d0B0FeSLrzBhYP9xsnlfEqn90OkVsUAuTipe
97cTN1L2rDnzZ2FX3fLmxHzH0YXfI+kOXdSXVBV+QN1xT+1KtN7+wAklKVdD
8f90oAury4HDf9/iy72ekGvP7ECP9s9cTlvs1SI2zhkn9AvVJqllxcKAMoTG
CODvJCAuVWqtQDG3StSNkJdmaKp6+7N947/zOXWTJZ3Z5sgNv/LPewQV3Zl2
sZQ7/p4Mk/z1XKnXwYgcXodM15cjq1fIkyvL4ef+5CiZIxuEIFZT2lt0JDCg
ib4owb0ycYsJZ1xnmb27WpWtT+WoXRj/tMiDkEb6yR0R/zCw7xMKX2UL5erI
ulyMey9srkj+N2NYcZpSo/mczk9KEfbzl/ne79l2JhDnkwof3osHxZKGQH8u
MDQAMIZUj70flC1IuEnq87mWP+4eo5A591Pp1PJLWeAbwb2xsmEsqHHtK9hw
Lr0V4MMwkDeuhawjwoNdv6bJyzCjItRJkRBAChabJG+pUHl/VYEnzK4AHCaZ
mmODkuv7asFDPnVpfnDUYBy+//YsN/feo9j0AuAlY3McXWnpkXzDEGW4KPsr
RN35AoJErVgubiCEuQEyzh4C/jXpZPWcmXOYFs/40K7t6yrWxhYcAbxMlAK7
G8x1I/FECdZMhK9ftwX9OxV24d+pcqbFDMoNcld3H6SUwg0ffE7XVQfSa7gD
47TQ0zoF9GKDT6jw2ru0TjFI0RcFbf74Pf9krAI4lNB8fxIXfM9NDuxgWr+1
rnJOZnaDVVpiqOGgtdtplsCTVh+iU9DcphgCkdl5I5ForBNfFbmsrvxbvTqv
W+SwCb+cYqv/eAZFxeDwC1CJ/PBusgvAWg9gfle4yemyAtuF+9ChKqmox0rQ
kGwCjOaj0R5rcmLNz181cOye5g/Ts2DWrj+MMHI/zSbphjWrWKXgegEMaw5j
Bvl6swhxaXssdMH6MVl3wUfvl5+qpaVMK3ldCqO7td/Ls4OSqZRsms4YyeOH
i6DkhzgixJYCGbdSHGs3y459VyWguxVbGl3N8wwyzsDgKibxIbcd0jY7hNTb
g9HzKot2gDdNn4NirgYSasRzddDDFqVoaHOwXJhA4BTolt04KDnydJL0d4mN
+WwXPgRR7kqIO84fgzKz3CYXoIKx+PSDEAH8P7jiuewxRCmDWPoXDgmG6rrG
URDfM3BtnfpkKDJlK4zT6R6qRvQHNhXDi8rclNLJFI2at95PuAa1sj20QjAt
cZW2MtFo3HdA65hVErwqCsuqpBNyvTLFBCu9FpJpgn5mCDsAnNJWCpX4cueH
CPSAarDN5qv7oRQk5fvB///Ps8fIw0eGU4gkoN+U/h7rhrd8SSWO499VDhaf
sDCc3AvdbwHnN4mApe5shYV7/rcEgLvMJaYPxdih4/HJa2qGtDiyfQ0tsOnw
fIqp/cREbV8GSo4Jry4O+5Lx4AM09hRouAi3iMyUILfhgUOe9u3SIzYHqunR
R26z9rccs86uoYsUbqccrSEJambY/UE5ZIj1mOKF+Bz/2BSpHGqEx43waaAs
lMRNi7YcIRAqn8Nq4EO2uM47/sL2LdgdWEuYj+GljajTTun9dCPL69yw816P
xZWH1mhKkPtbTwX1Tpb0FpvyRCFTgE7frmOSGEda7oNwb+rpHpIAmF79Y6VP
ndHn1qHQWI+j25tKrpBqUVPaWjUtJ2IDaldlUSBXJJI4HjFvWLOPwYnqGZjm
LmGwWbMHD2PRRJYB6M6Vnz3Ft7uxDENn+nDiY59jCp7hGu/33noBTI+P2k7I
5AZ31ob+6kjOtqDMsCtKGTLEW4uYy4pow9kjztnciuoPtiWOnWfTIiyoVry/
m4NQYqATm1yyHjQa+eU7nmS7Iholmo8HmXDwLuiE1ORcXvK9ViM9+HzzU5OI
LpIe0r+wdxb50x3TGBXfson4L41PRUNka4cOzLwE4b/Ne/Nx7f0EeiWSvKK/
eP3r3O9vhxYI444+nKjH53W3325a2x1HVDktW6dPc55nLxIa74JW7xsaYjmv
VK99+7w8dC8uMGyf7ZdtbfS0AEjIfTPgiP/MmiT195Mat6AmeNduhBxJUBod
hVwCHC7q2rWn/ItmKy2zNj1JmgEkYCR83d88ocxNjqxg12gphd++3N1qwl4D
f9qpJ6id/n9Z14ULkseSCsjkfLh+cmI6TaWMlcuScve7n67jfs3W37+YM/cw
rwZJuFN4f075kuobTlPnN24TCJx+pV3GIge/hW1YLyxc83CzMnVGe+4KTgo6
NbbGfYVFPwRhAYQ0zAL/bmzMA9gWbGTqVkH2DlVyzlSE/+ISJ1gfjAONqOKv
5C7F8TTLPlsC0Fd633pfo04itiIvRIgMU9xDnCZfr5VFefHhaDgP2akG5vck
km8gw1lwACJiRcc4vj4mHcvDhoRiS3h8HmZDo76hB1yk0DuVAE3cX7dEKOd2
8yLLCmzzFS8NRcPh97y23mexnLZKsazyfkf/1XQLFrYBlbu+eb+A9x3HIpo/
QJaeQtbFNNJ0ZfhPvMDUfGBbR3WSnvjhatLTuNeaotZ+GHxfoL2Yx/SnCHMf
hreyvvN6HHNTkORlEOPwBobDj5V/IUROl/OrAHePfcGauGOkqKKt7lMFjzEd
D21pQOjpTZpX64WtqouRy+bNVEi6dyjqiLEVj7i7MW3TpsCSzJkdHbKoPKvZ
fJn76m8ly59FDweXziniijiF1cC8T46eN4r3M4jQmlBI8hx2Bf07zFVN98po
E62dR1bFpipewGtzrWw4Ofxj9j02OGJlG+pf3EJ3tutGsiuDG9i6/u+B6u+a
ORljDa0sZwXMlirX0jDY4s3mfqOp6rwcm7/z/0l+544plm7EYXK36PuksZ+Y
gsa5euYPsOiko8+Gwa7MDwnqIAAbbGf7fcXL/JOLseYyjYcZD85ylPxBfJk+
zHCWhPpiSj45ZthfehzgkF6D3JDicyAnw6etTCvQFkTdlVphGtChMfY0WXBK
naCruIqaBYffG8xMsLinAbXcJfRkGb/6hJ+NIr5a5ylUstlB0suMcWDy8Har
l4lysJYizczZyYPP6uPhArmcmhhgr61Qd5UGjr1T1ExmJuxySCbgrCslyadi
+25mrkQCQ4MlxR+4lcHi77iXA6n5RVe+9lXR80h/wxbru3X5uJ+fwNfjzezB
zMwke4JTzUJIiNB9OeBHY85x+wSyLkFF11EscfA6jxYu8D4fn9exBtfa6euX
h9CuhNvXBi7mgfd78zahJAFodAlSEmRwYa/38JZNI+eMM+w6euJ96mzSTRVb
KAmcYoqHl80DWmm+mp9o134RxM6yS+oqzW4r+vfuNncxvGr8NBRw2a76crgA
g2z4ZIPq4IvidO3DTwLdj+dmMoTYTW0wLA1LGxXd1ZvAqJbNKxQcMk88eecO
l27NiH5WIzhj+26lMsLCtlx8XbbKurrz+j+eGJ3knwi3nLOH/xpCEfXJj+ju
FnfBMzmKu7d1LpyWrz1kLKPxCzrNecPz7Y3QQIo8vKuVeeNnkhEF9+G+L1hy
M1rHmHjOgSy02sr9Dx/9SmwI3lKeEH364UWs1KopMeLTicJiPEn5iSFtxOSY
RrVjz8GMbT94eaMHLT4Lme14uZlj5/mYOqhArwNWQ2aaUyWhMCSMDpX7LSwA
W8hzoI/Y2oJOF/5eiOBWGj+9OHzd9cx4LSRgXk6NHwquKjMwSLQUwzeMX2u9
ITCnZSQH7hQLl/+yQp8XsQACCk//4XVgMQTaHYDHS6A3+x5dZ542kRDeRElE
Et1maK1HnXZp5Q3AgLlh9Bni5n54FrRbiohmC+9tzFGvvuOcnw5Mt8Qq0ZZU
xgZCEKzLQyoyzoYj85bNc0kR4Rcoe2ikhnKQpUOUSmaP+zfA5VCKRoAwAvpo
fNUwj9Y2V/CODtJe+UMg7UGpPyW1HnvUwSmg4gpmNVSnmwNIjMkDeDQqrBO4
YT+zKZNCmrYGtmKjKpFoe6GxD+YjEsSv9xjcX9TNNgPJv1F2ut5TKuqhuWYu
Q7y4xnFagn2NOqysTe/pv+Neov3kdSOsFJr+3gOiHEOXdskPQ1gO0grD6Fdr
+1IXaJ5cbXY9k1Uimf/J1aH3B6UcMi6ZbXB8NE16UaeDzkcMxJ0aqG8+WfBg
X79lHytDlyI3YOkBjLjvHq2Fc6uMAnLWk5Xetk+7yVT2EvY6uORFDj4xzYnH
80EeQnlW4nXwnhhgq7IeWhNm8usKuX0tKwr9PFDKt0H2FJypA9msJNnmumdP
+AMDtIQ5f+SFpZbtu+XkegbHEoxVUcKgMFfbmc5A05q3t5li4L6GP5HwqwBW
LJoSy4ddEzIQeSSi6sWSOfcPqXS9jp7IyPjNwHBNhtBhNt88Mwd/jaXu6tPg
k1Eb1PgdXhngstgbXathAQ/AN0LdJTWdnWDBW3+WlhbZc1LzCKa6rYiU9WlU
m2H/FQoMxDvVj/IF8/l7e3/0mPmTl+oMnlsuz0E5hH5UclYUvUjStyJYI4UK
maFg0qeEGod72SmTvFSrAlWPyHdw/FepC+zcRYaS0GH7Lo9KsIWe//z8dtbC
1crYS1O/EIpkkiwJohhQcBV+1MmDBQ4L6DTED+X9k88H8wgz7xgnlVGxkn11
Ek1giv1uMiAYDhNHvHqoFHq+2S8/Jt/CljQBEY2yE4WNHbY/0eS/J6gn5XsQ
nvh0X7qtXgeEHzZA++69aUNQXiDHFyO2IrSGpuujAiRFEV4naJnz4tGNbzV3
S422UhhCS/uBxON6NG40/5uwxBiDVOCYHwznFOZ9YOcj3QP8Tbq1XxJrNjiO
ZQS45HhZSK93v4gEdtdSvNDrxRNa3yOT4WzeebzuG186XJtc05Kd+0Txty1u
8GSAXEw1kv1gsVey427xqWiukj++TGslNuqYc5EMrB6hpTAOEDsdtW6gMyWH
zO3gnyAwCYdDZWs8LJDj3pqHx6Jp9w9iu+nE0Fr6VAbViCwZEsWc6jdEz8Xg
bubhmTDT2bPVne6VP20C/YN8AiW6RVFN6LAY2gRPwffheDhrPvKoxrIEY+pO
1sVmtRLEL6ojKRc3kg+B5GHoBodNgoDg2vEwNep45p10qhwDDaCK4H5M+Wy6
qJACybZi/IRkjdCgDPkO1y+QZA2q5KSWKt1U35nX1NQ2GGpQ3kXWjpj00RRN
QH4b388nQDkwuuHEbizCaKNSwYQ8n4zu+er/M3Ebxn2vlMVBrqYVvM3LRiZd
3mk8URrugGC6QzDw6h6c88tiurZehzb8Jf4y754JkROcBxvMUPpD3njDeTAL
HtwQbWhVzU1NvV0226w4BDH3Zf6R3WY9brqMvoVaOdQ+ch/uHrM/fPwos0BT
o4G6j0AX133gLOwIJhILUaFqwqduJw7vrx1zUW0TegpWmdg48aCxAyIwT7Vz
KQ0L9hGFAe36TbSGBggUHkc3I8z3C4Mb9qnn2iu1xxW7HmXP1sdvooIdlGls
9AOoGiQIXLK919UWGL14wZv1TX8oaU0BIA4S53B37fabFjIOLZWTIVBw70Dh
PYqXpezFsbxhamX6LL9cB178x2OU/JSSO82VZTf4urPMTNXuUVnUsO5vgIF8
SJWHyji6VwZA4HFy2YEB3UU2N1BCDQdeovS8LH6ldnYgctvXzFvSa2einhPh
LFSp8rK1WwmtvUkUJXC3gtdJaqcDCSZCmd2X2EpNZpq2dM3H5bDdHBoFVo7V
gwmcy7HAHEres3+g4m5DF4PMTP8lU4RcGsSiPL2GO5stiZmKMLXhSQiQWZ6N
JCQ2p+2WEVyNAReNEyPjOtEL4jwxlgXybM8IvqLxGdJHn9XCWD7reKUKIrJx
reXdz+swW/7MX4C4y7gpPz0RDCzkaR5EAcBEcO2fodgSPvCdMjUklfzdgUWp
+NvygtjUcyc7kKUbforCfqTqYVLdQVh2I62ClR2kQLQTWdcb/vxYpKMOzsnn
jAoBeg48/JmYUpo6MzpvMvqHcd1/zQJceHydxMeB7gZbLKoMBxCp50M3T0rN
AZ9qcbv1WzuRp+u3k+Yu0AM5e94ujl4W2mkeJxQo0ACVJ0Y6IKCp/+KjNoVj
ryfKyEJnDDkiU3O4SZQflw11c05vW8ScoBIrpVCHk98Tmbcc7WGFN1Y6z7cs
Tbucm+b2N9nnfM5D37yoFfAB1wnbV7WCA7Yzk9htVgtMYqyB9ySUDuU+qtY5
4yvQ3Gc1ZNwgF6Vf/Mfmw34/ILEBvpwiIHgWwQJjUDrt2XyJSnlwdfxpmuwC
Xh3UgMhohvI7uVbc4JJUyyrY0FS9Ng8FXNbbNt86eld3OlDyx+7ofvNeHKS0
31OpoXAYLetEZC7ooa1+2a+RXKMg3D5Pp+mvK4EDy4qS8pTsB25sP3BOLs8c
9iqQMh7kJizWVN7ne0sQEmmnynmDfn5nsukm6RnRjGxNNtCJiThf2BBbEBQg
nO2BT2/xS2p4xLX7XKxGKjSLTJg5dWQHa/lqGGerIpbG5Dcm7lXEZM1wRheX
5QtYFZlk5A+KMmRILmmYtk11nn4blr8KJavpDIbb8e1pi1Ru5+V13WmwTzrp
3vbpmXxT8OlwL/MMxdWRXSqusw+oJD0K3bUl9taLvfV+sqq6qJttnCMVrjvl
TrxU0BrZLg6BXalhitsVnNlkvO4c4JFa1Qtfxfra0QaB4t96xRh4EGapn+PK
B0LwTUylyECWN5FTBvEXE9QUj9goxe/ObWegfCg6uNIs/iIpUnM7WnB9MFQ4
mccawr3Gi8bEo3K+qHqUEVuaaVQcVtDaM3dU5q20teyG9LptO5NcGCdI4zO2
t4+3RjxES9VaK5xMPXw89AURg3zQGo4l4ujY9+Vb1SfaJg4EhX991Fr6uqL3
rVl2v7b4xBsqAB3Apj3rbt6BzgIeMoKXdxndkytN4AwkFRs+a5wYjFxS9oXD
6+7DdIbLUz2pkiGhhr+XQdlmQLF76N/Jn13vPr64iq6Erj4ZRn5h7WXw0TYU
C7ow69pmZ3EIm4NbUQlwBUEIsP0oSvZaj73tiOmAzUK7yIZ5ft2RoMpVGBjq
JA3dsDv+a4/QTdqTyvAkoG6Ii7RS2tfbCLTgO7PTBOKF1U6Wm8DoH3aigdG4
nP3+UoEUAE/lIGjEVXr7lGdnJyrlM1JT/up4X7X+EZXlHWIQYWxyS1/Og0dI
WqfYiZgkziyuqIq9Vde/28ly6JLc8pOkD7IK85abOQNr6aHOBJYk95lfTVJr
WoIWfgHPJ5Btqr9WSjj1UhNrjbcKJn8Q3YUNON25j9YBV1hBVqaSEgQHy7mA
zC1d8oIms42IMJYgeJu/rJ9/TOrqMqdTJnTa2x6rINaBG1cys3RdaqldvgIZ
KRflNpbt0P4UOrhQGOZTGC5OqeNotmrJooa4bxyeEErBOUC1w9QK6iIQMrbB
djb0g7HpAy8JBlzR32Hd6vXgYVVqDM+zo1grtAh2pTZW+AabCM1SaROWe5Q+
w15QjUzujJLbyY1+4PAJLosuXGelA9al/OGKWZrWExJWtcB9X+Q7oWNuF7MJ
13eIViXfqAIMdC2B6qIjHAo2eScV/9bN7VQpoyPWKFHN9z+Gcn7GvzCrbAUB
kOYU0VRn4n7yJ4CHjlCd3F9KYT94VHf39gwpDVjedkOj/Rg9C7TMOPgtZxqu
x6FtNco5JvxQoCr/ixpRT/3E6fchnA3UuWyFbBPx95QoUwUojP4EbfGfj4ul
c1Iho7PkFjQkN7pj9E9PlRPcAcT8N2I81Oj4Vv5JjOXZSJBDkhA+poQ8zekU
1ESNdsTo7AYeTcETSMhcd51PjRTMZAb8S8JR0FGnZXKKyB6KnqOX3Eo/251E
FMSwH+A1lwNQw16hwm+tnaBRQ7s5MxrqdlHiaI8nxGJMuasWT22e0PdNzUfV
I8vIzww8Tw0rep0cLkhyJwMEeNAmOwC4KOA+S1e0U7aSDqiKKXDh/mEdIMD5
bAPZ6OEZ7yxuiuvX665TwP6eBgPKyCptSuwXq9TkdCgCRZ/9P1piQTgYZkph
v2DijP0immU3SBevSpRlySlpHrXaMYOvzCrttvFC/AfpH4Qh0rXdfKx+ePNZ
iUQzf/WxSk9P8ZKBXkfdEFTbpYOofJjGblcULZsUQxAJ0VXENtHktbdx9zrU
en/WBEpOD4Wrbj9xB160zEALb6MjIXzPq/kzTEAzLhZniacAQIvnj5LbvqC5
5XR9EceIZfGxi8Rr7K9lythKyJi2mtm6At+qB3p8hwABpHhQbIQYvuUxVv3u
aJON9g0lsUFsLHJPneBT6+gVpnjYgcwTxz9nnDxR7CQ79oZqXbut8y8WQZtE
3agVZgHf3XJvbkvckqVDOW9aZqwrXp7OS6Dooj5bGdjYwpTbjtuwK4D9f2h2
0wiSi40BkqLSP5sxDhm3nnzMUZ/y1JVKB/oBcwtZnrVVhxFjlfum1fDeg+8S
lGkjWRjkD9fDgfqElJNZKx4E86hdutLb1knnMmpEz9NsvqnhH9pn0CLwPWCC
q+0eRBN5zCy04vmc1Bqsxpj7cJm+C52vbF29ZuS4U4HyOBRX4Rx9f2ZeVQMh
tbLYDhvuWUbr997km4b+lZsHyBjHC0pghpE7EluBHzneT7BleDXxPvNYN+ck
cHPcSAregYu6BY2V9Q04Qo6hZFHZe9VFKyZyqmKA5mZ2RCqd8vjwBIYKtvip
1tyRqJ5/jWC8V8n67Z1roDs3Ak2rEoXGbssN4c30hzzAyiYG+SZ2yj9HM0oO
e2qh/zM+ceYUfkcGvrbB7R/ghPhTIalDRyUiuYyeYuk8w1UsWdE+8rqnDQT7
uHCFNO7jY7wFlcqGe0Js4256oEVzmsKyFJwgwtK452jLMrMTAgmEPg4YA3XC
6ZaO0UX0WZp2Nwqg7nu1uT4K/JDBT2u8FyyOCy6asp6cWaNzWL2WFx+0GgAU
SapSxi1HM9jzIaHvOXCt0NSb0btezIMiRoqoIoQvQvGtHdGt/1e9m30cPVmX
AO2U1EyDAvMFbAhHBVQiMzF6R/4WfSpTMKZMhSJ76vkZPeQa78wb9aP2jtXg
G90SIuhQe4mrVSuNWXQGPCUONLrRjkwGRnVJ8GQZf5sjLCyrxRxAdoutyFz3
xjYY6mMwCgBM6Hq+yze+ty6ghH2ZPiGSKdb5iwPxeAAr/xf+0C8hbWY8gsrF
T3YqPiCdNu4ybL7fn2qmvab7FLX6VADTcdFNAWzPYsNOjE2zub5kZYfMcQXU
faBlgydhSexv9goJRVIyDYhyB38n+JpBpdbFUufqZEwmZhNKlGzzbQg4JjFL
BIQcpaLew1hHUJxKqcWhQ97OTlL9qYfkypVXuMqlulCyz0kAm4guvKwUTLnw
g9im3IfOf7xchNtXbtaKnB7NEr1ZJaKZ5ZJfSbMUHEdxlnKfCvbjA5lGiadP
DsLRL20VuoIFcL4JoifeF9hWMhSaCrDIOBJsb9faUeJYCIfaAoG/8Dmdyg0F
gWrNfdwhkCDRmSxGCajo49C2TdBly0bhQyC8lAp6sXaMMbOfZLjEUb4NZAtU
n0To3Atj+Q04bxkC3Wj+0kHjBTTFWusoO0HbMIosyspj1rokl+2+WQGvNbjV
b1FRENL7V5swY10WtJEi0yozKXUkqNfNaGhlkTl1bjIx5CxM7lwqQ2PE3yaC
o32IrlT3ayLV8Bg37CPjWw2UiXC+5Tpdw71SNCR7ntQfJ43EGZeAyezs/8zI
21Oxo2Ab8DqEotgs31B/3g6eAi8Fm12fbB/Waa9KI5NsWGmAFQTogBQFhp0l
uKsriHtRJoZ9PgjcwHTowD9p4hSm+rQx1bC47ZzZg7zXlz3N9oXl4/RAC/EM
F2DuOv63dZa4bTlzgeBFoQ+nAMBskoyT4YkfUkzJZUJHuu7BE7FjM5VAY7Gt
+JiDbxhshdMgMy7SjRcLy7pnCrG4llmn/S5BaOhnG31Tl1QHBbujDYm/6t4C
Qfw7/GUvPy/SP3laYHKqoAbphTyah/bozIzsPm3Lguh4OQWUDC9QEJSzORgP
/zqzXKGMPg+8J+QyNvYymoShpcnzEsgQpBUDpHoBnO8evRlAtrsHGo7Lk5Eo
MEBhsoyTsJip0jncqfDjHDYUI17CiZzsKEHWIBUVB2HKKgv8c2CyVDmSEFz2
EA8dQf/b6NPaoDNKfH5gRH+BLGcl42f9kDwR90UjkDqi87ASBDjJ6yXA3q+K
THQO6ecZRGlQfGzoH9e6v97b4Xtlqizxu5RBU8cpN0Rykv4P9yERG3telNVR
jimhIjarEvJf3i8SMnwylHGQYWKeeH8+RUF0JK2UKSbpbYEXkcp7fovtLRzg
fW8jr5Y2YLGLNL2FyNYxHTlWVPLfU/d8COTZ1FTnxq+tUuCf0LZOMo+HmQl8
bhkvgb92VeLGJmUsoWAzoFLL8uHAOFikDgvImt5pC+f05/D0sGkS+aCVb0gz
D3m55TPawOtpobt3kxT7i97QNgvRlzwgBUwNPNwBJdrEGfXag9c4flqCB+N7
sHsCzWNM5eJrb2VrqjBmNHF/h4lciEsrnEOWiGG4suww7l6231n14rWiZhdy
m+x21aIh7I6U9sNxLPy+4V8V3JKNEGj7oi7mqoepUqsL+GHNKE+inzyErBVU
DtkovbknvwvDTmu1Z6KDLUdIPBZUTSr65JtImUXLpfj7Zbsn17awtNGBvlhG
6+fKCNjY4BkYHHZx9Vhv4mqcUmwuYK1xoxWwpMb/ysY+IDNKDqRxcFip5fse
azDBGYUlj4J8jrq48Zpt3SYY0LisX3u50sdpm23uEFqCr7P1zf/EBZrmrfbK
8+yeyOpaodBWzxnKlDC0i5aRb3wvAJA/paxFMY4IILimvuBq8Chvy0nxqzZh
Ff6TliOOfnb5z4ScUGBqVvBq0joPycGDMP80iMixF/8lCa5wcxRmFbPbMUeg
SFm0oOxHPXMIOkwhXPwqoyGmcxQeSiuhIuE/piuZVm3+LW1R1vSNSK1GVU/D
bRI2yVkIYO6maHo5/FmP/as7avtGVnKqEN7XCgsW2s9mppbD0BlsSoJsk46r
/tceo/YdQOt65U9hc8qP57JGvFFabqrSvVGQIBB0le9gRW0Xv5PNgAuxUZpY
k+Y4aYirOnl9SGQcxEwVl6SPwmtH+ZUJiRCd7pl+z0kadKawbYEzsBdkq0rK
qDCHdQsJ+TawLiZcLZ+NVmmJVTXDRck3zM3dJvX5eTpVywfzWIELoB577b9I
QnauurKZMcOaWGLKIX4PCQ5fbmxOlUQZyEFcx+RFaW9CLsSwgIsjZPxvrT8z
bnISNiGabwy3Q1RbfvwSw6PhCkcXVxODHnMQpJodokT7txZ/yc7ovkfd5V8s
pkjqgEz29NCexJ6e/4XnDsk4zRTY22+3XlG6D8vHeC9FOdyNN/KzZMz1vMhN
3XHCx1eMH5vLOesrNLVgaODzZFvGxznumRonVZABZRuy5IPnQjJMD2L52nW3
/eStCpyH8QVe61Hy7XlAHcsZdHNYVnS9JksrFEn33Knd128sEFQS0HrcQHvu
qhoVjeoBWT3pupJVo804qBdzY3R+LZhm0+38oFN9C05sfqC4SWDrlOj8CxhQ
b2bkTRrhVe+lzbsB/gXyZkdbPCZyeZqgCV7EU7Q2unel/R1yl/fsi42QdIPK
Jm/cQWGaf8PkdUAoG/LVQBG40LUOLjs+8p5CascGZoId1MzBuU8huLqSrLZ9
JkLnh8HSXYEhcFJnmZrT8qTH4+Twk6xwUeGxuVaLOcIpJhFhdmvhRpVor2jc
FWJYSLHylJz7Ps8EK6pT7lxmWpRuAFOZGm6gyIij712uuoTHauQdD9pe0nmS
uljsdutCqC7t8LF9uef+TQrE4TtPtvk2irJFzipDahAy0spjzUz5vwSKCQbu
Bi6cEnWxanNc8bEgbzw9vM7Wq9W3YaheMcNTG4dCVL1yWAnEZmxlyHJ5fJHW
C9kovUHpK0RdnCsgcp1yWpDqrWyByglvYow3qE2NgLrkXcIZ/vehsh3w989/
q/bU0UlzaaFZi4TYFOBgtAtI565Skz3fzdXRHV2gmuUqhxcHawhUDQ62

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qT994K5GIMtoa7mHNTPOq3penu9FOpq1EOp+Og4MKztgJMS8lTmJsNA5dGz0csTNQfyIj5R6442EJ9F2RDNVU0yc9qtJVIRBJsxT762XzvGWUUaXt/V1ww4hGKimYRPKe4PdCJQL8wSmjhoSm1cAu5hhL8y59Hh+9LoOGwNU/rafhjaOTatAgZqd0wL5H1fQU9/XJPEob59qYAtipc8NzYfRNrvlecDKO4lVNLSekIuc331dJXAWqTt/MoouiiEvLXA1C/MrHbnxmJjFzW8VMSAjuveq3iDuF1n9HSLwgE+C+micFcptTsoxQq7CKtqJ7c7Lg/R2tzOlgC0V7VlkbpdTj9AQRcI5KaaVwT7DjNz31vsZh+j2Cfm/opl1X8qzaIa0dQwMETe5dIgHnILAkPE3R7REopq+wlsiOxx/YJhhzrOCfrqSeGL4PP3A9EUFY0wlsqsx3dfaK1Y/L9ngKu1Vo0Sdm+cRBc+7lTFHKq2N23qAPVUkKUfRStrZNHTNpj9AIq8HSrLaYss9RDZP9DLn6EyM2IuB795m75Ncd21sm+KTeToqdsluGsgkvorFX6FDshW+hD8ntS4V1BMrZfH1Jy/uDfpOjfWTNkWBZ4BBDfm3SKqlJMf9lVWjHIH1uoOTnsJZqLA0M/wMzHQqZrZhC9Qy+NU1LQEHoUs3pBh7J086L9R3xl6099LBU3KywvlSyHASeCCq8HOC+Tj/QSqP8M6UI73bt4/xcvHZrT8QVsx6coSxEzPbsiwWFDTXkiCfK74gFptzD9oJ7EPbKsJ"
`endif