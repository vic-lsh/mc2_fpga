// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0yx34jGfGVzDItu2o+36zPIRk8rLV8jaJmPWSGQLt2EUtARNc8mdOOl+MwUQ
Ilg0+xP08AUDygVSsItoImeJZFtH1DcJH0ZCYyKCI5sytwaZHkL0jin9HDAU
bBPKCKx6WbTpzrL6GgyYvfcXz1d7U/CrWEkReOkMAQ5yKobCGcT7cIFlfP/Z
iYfXk6Mdj6MmlflM2iPv0yWZavjwGuYtuXuwU1sZNUxSLw6n06UPmHPI7EmB
BHhoIrh03EdJdZ6hjG+8GJn8Wx93/djsHT2bve+DTbfYrIGDbmQ3ILenE5ZY
+TGlZrnT448AHzbYi6cWNwXPeCUwsXoKxUZAq0g6oA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JV/x9UgmsfwarHWkSS0RdAPRfCeVzvKKAw/Wx/bEBagaSFiX8v8gGFbAJPBt
ybOS7GhYlR6jyquGcLby41IYc8bpwvkTv+rO+0XrARqRK5dXR40egW97+7mM
9fy0cTUudhVN61fiBrqZGw2b0no7CDbiD2f83krkZuR6ASTJ8mmNqCL8zrg9
PagfNAVD5IrAryUYpp2rhdjLDdL59wpxYqTPCaloODMrfkU5b84ch3YAm0C2
xP0hLAY8ZI+s7lCzAtPlQZCtSvCVsfI08Hk1CZbtTghIlvCvqJ85V39dIXYL
vW5gVgWjJ6DOrYkDG/GH3L4xDXplev66jmRRZ6fwEw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cEbun1hy/5oDpiaHalmgwXmlvupmi6aApJW/UwPXAA5MTRpTOwBoT32vXlDU
G0qgl9fZHsT5ogQpUpALijT8Mc7H0o9YCXtbBtxLGTvBiq+hicnSVLgaGvOr
8GKl7l/oBEj9er4CLK2po7CZVsOe1p533Uvo0UiFHO1V6nR14tJ7OvjtUu6r
3wwhmxpTSmog+m/2osM3HsR4XjMrq2ODTsOhUCmWmE44FtarOE2hnU2Qnf/3
fzA9zweM69CUpxv7dC9/UGSqt1UPkgUZMBH3u7FAKhihn1cY8FXfbiZPljoa
OYtk01ThqGm4KNcfgLPX32uEgOGaL29gkkqXXUyPrQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kHzcoHT4BTM6LNiFLogJ5mwzcXapJa6XIBr7ianRomW6+1febTAeUXocXjV7
jW7f+8evvcWgeYhn20l1dpG/vCN/PIT6fM4MV/xC9J04QjisbPcNOT8kw277
PQ6SSIH09AWiSAKPcpBIh0rAzMQfg2Lwa1FFoELp/gEceObjujijbrKR5FwT
NCy7CRn+6Bhn1XwHxCH4jhu7Gzm4X5Kz7kPaiYG+sJdVV/eGQqVqUH1sLdpS
OMTmM95ZmgY+SL56uVFzUaudn/fOJzxZU25LyWvChRHDZDJKdeh/shynO71S
Jd0H6LZm35t9np2kJ6hBnFfF0dGWvfhm3UovieMnBw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nOZql7cezpocB/yylYyucRrgC6JKJ52jBvU7SF5mcH2rhPLR/8s9n3jQfg6B
MIfm6+eyqEwqGfK4SXqlT2M2mS8qcQX2UpcpZT/tZ01uP5YhutJJJAHWtxoU
gkZ5Gr8g4oryBs5F3MBxfyUnZ+vQj5fwUBSkM7Ke8aPb7BFj4H8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Vk7fnLhGAIAkWi8IfYvHaW2QxyeBkFGvLsfaVydZoSurdMn+hjkNfLweUk1J
QVm7x+GsgffpHwp255m+enInhS2SNauSe2bIniYsZsAnG0DeTfbRzKEnWgiF
uD4qIjHxW3fD8gjPu5Qd94vnwBJ+1quUEpuOuCv6zBQdWdxjMOuQJRk/0zuz
0f0nhRyHxnrkYkIw98JEHB60LwTpesmbVHKfO/S+mvJb8oB9awrlZqi6PXuN
5ELs6ewutV5uT0Xja/FXq+Y7l3MX5JC5mzUee08qBny24hd70ZYC5sGmUGXX
gk0kokWaWvOAJ2IEfb2FUbPXmY/2CFd07KFMMH3ukr6oI2CAKWwq5NbrXKvW
zuuLpljzcwvFezCdykSqVVrWG9xpP6lrvjzNi9vslW+bkqeG14aXxjac1/RA
OocMGvF+ESVCg7Tq1XpHcJm6YbkkUeilShrQ7d42debD6lHu1BiA1MwU2cx6
tbFoS1GVfxyrIo/nPcNt9CreLedTtndZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ib3H+/xwtZOU+kVXjoA3uxoa7iq98KHaj4Q1BDBaMDDHj5gUJfyRvGfx8Bm8
zumKGMOmuWfVVpcmtYhBAkw3kZZmk28O1d5ThMh0bekNAgpzjeaTQN3ZTR29
ax1LDQE666TxRaiAF0kkMsDLSkbeOLeNG65UoGfC/23EaPVWBVs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HTRuE1YmU++qZ0KnA6OleTu5EZK+mJvnADmGEiRO+t4mrJhIobRjxKBs6s+h
B4Czx3e4OSbjnnVLaH975jz7DN7W2OEkPJAmxB+wMjgtVIvpU5tm6t3jA32D
aSOkx//ezH5nCvdf3wuT0dw+SD0flGUT7/tLQElPwfY2wvBdm68=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9808)
`pragma protect data_block
qep0caZzPqAXm6paYe+lR+fnkm0yk4LnK9FGNegiNF3T98Xlze+X9WeZITIr
MYO/hvp2rQiXPRs7aAw+W97Al3O/mc+0lx/GFdA6vQdW8eGAlccA/S6dicds
mLRFO+ndXE5qtFkgysbyOOVR9TOi5fIMmgCaryfGeHYiac5y6rDp5V7CRCwp
y1Rqcky3I+FxcjM3gPoub8KP6mYWdWof71Gby5qsOX7/AZfDHTkxwQnANUc7
hGV4zcbcW6I3+Bz5qfOEgUUxYrRR5tf1yg1RO9wZQYBkmDtDePiP34GfNFHF
3vtN61kcQfju0wUdRYOA8Kty4JKYwkiOKe+HjagQUu7C/eq2OZyBlVOxTUPb
jOjRPyPZsawErbJqBS5hXgCljd6YQVg4xwY92W4zMiIiqoteimzvDapdiLtH
dodPzolCacok7g7qb8rZgAXVSxb19jvVfF4blqjJDS6u4PfUu5DTZwV2M+2f
WNWqW9B5jgfHL362ufIaieaLvgF6Lj1ojHUpQGEH+tEt1LU5+Wi39IMOpqaA
nSwrKdYPaMPW26L7Vdnxmlim6qliUoUVjwhChFnmn4CBCEgzOl6GqRMTMgQl
tLlw5cIgWeHwbXETF9v2ZgZf9NqydXHfi0CReTtTsxK1bSD27B3jv+a6lK+Y
1eSScvp5RN9Di96sLcab4aeCsNirWnV2DMsFCUI8cvdMNkOR4wvg5IrlT4NJ
KtT9Pf0Wfay5KSIlYXza2d6BOF5IuRlmHbxjLQ2DBbfejWB2qykFt4WuWlrx
DScbZUExnrceJGLQUXS/zKCnl24voYfF1f4VCaYxFcsmnc7T64TuiPvb1CYK
thuP8HAMrWMjM8wmIiRa/XbiZMsQ5AzUM8856fALC/pgpciC8lF9XFvcs2Vs
izOe6eLBojPN0aNg69Yqe1xONZbVO5oU6s5vTPAnyTWjVUAVBQh+8FerJIud
BP/lpm9ZtisIvI6gVa+og9i917FfMzal9Vzw0MqEwWu39CjYL3CdI4SDCKQR
J7BE7mnT6Z1CEq48BIwWG8+SCt87QVobinxvy87dSxHTEw9nt2mKeK0V00y9
UTj9xG4j3n+P3RnOXBwSlD133zG6Qc5fdcMRKALfqBQr6hgFaf/fKLcvY3ap
dPH5UcLDF7sox3OfDyYlV+rw6S0QTds8mkBYby5lR8qap/9r6mcgW9vQHkDH
FeOIlmBh+MafbpZrJ/V1//dt0os5I4j7Pzu/+3MYf50Xo4erowxMzKIN0sPG
s+ewSFWSJ35xyrU0kmbisWkhigZYECUO7T56QlWF4S5XsiMBY0DqszxYcI5w
bJnxTU+E6Yflm6BwBTdc2TWbb3tJj6ReO/MOWOwIgPOV+o53XO4IrlWoehf1
bTOE05zudEcAxT/YVdOqQxnVpubMh5XqDTaFGfq3aq0Z2RvQXDevkrW2u7Ay
Ryzmu9lYnu78xNFHMMlBP9wRsLTJcNDgfKQ63hTHz2vaBrFFfQO8qAk2Aw2F
ZUA/wivszUN8mdztHsMDnOHk59Y56ujxBleNbqxu8hgRlwrS3uvAckgPuaJB
uPEt3RmZwx3yUiNAo1ht5MCpJa8VwCRNDDiblyoUdHgvdkpbdgBlwK0AoBQp
KLYq5uCx50DZ72+q8CeAaOX1kYTY6TakguKemsQmDwEsPvR7CMeZ5y0z+2wA
EQbAP7BslkBDCbWvakyUnsvqNn5zDrgyNcQT3ZCMHAp4DLgi/ZYhaxc+SUWf
BmHms+qdQAAroqqWKwizvpp3G1tRJEO4irJxNJi541IaOWsa80nuvsEj3B36
y6UiTa+lnePuTo3b+wTG+qG7tGSslTuCeSL3uMvn3dBQmT6WIKJSReF0w+y4
ioY0H0ZF3Lc/gJM8swimFNNcgy2qG1pjq8/Wxx7HjIVz3fC4t6RNRKjkmBNF
WqffBf2nO51dLutP1FVl6qXY6TF/6xmXVUNDg/zqMK8uVF79oRFLlTY1gjIW
s3CFYYfoy6HrKt1lwOc8h5W0JmBBBlMtonpnZuOznsdQauOJnUyh28S7MGpJ
nCCeyhg/xLr9uWvl/K0Qjjw+yO3dRGqIuZ2Gto2fsONd4VjdgbG2ny0OtMuk
a8xBSCv2HWBiR9tavHjKb94CbKQYrWdKsiEw+KInhWY1DYttD38r4zOoOtcc
d9fHZQ+73k2vrbl8TXKFFFRx54PzVhyETG8l5nf/VxJAfk8eKICqS+8mh7sW
p991plYTLhGbODi86MeV2Sma8N+1z91FfiguXjnhg2lJ3j4ykNBAUCLaORZo
Ap4kIiwfae82r5YfAdepjqK4rmF8Kvnoj5a8+Mti4xjmvXjfHQdxbA2zHPPl
f/9AP5K/DxM42KvZIjScc4YPtCqUpunIN7HS8HDugGAvfDOc5oHUjj1WWBfT
0lfNGHQ3J6sQuvDBnHqfKBAkm36nETT9QGCVW38z2sXPK3nIl1irQdBQZfKn
wPJBRCeAu8EyMxBMWv0ZBcsvIuiBXpSw2jghXoZkuxIfY4/ccQhMKumyDaCB
PO7JR5kf0Mkn6MPyyBaWrkKFEKogKxl/0ie+nYYehrqlw4DMWcdaefFOtS07
75nGiSQCGXAzzTbv0J3aQcYR7+2i5HV16NKt0YyQmq5JKcy00VERNKBUsalK
Jh7psNIYKQAWiuA5JoOz88jHKucRth7bUQOZJf7p0YoEKsOzgVNuFsOq50Jd
PAHWjeVgTeF/NOyF0xm97VOQ/5S6/Wmkiz5ECoI9KzteKMlaJW6Vf2nO6sH/
354q4ovdDomQXgZq9SUDuPECYwUwuLUuHbZjVBo8h09TNApsdrc1Zuyoufyj
T0OvGepfwm8mYUnoydj2ocDKl03L+7Mw5o3WfRpvVWISPA1OA3eBVHY/pXyM
aTinVI6GlW57xo+3Hr+c+4cBk1apqxCHTDe1SgCcYIAZYY2YlKtN6b3l80rW
ZWUKtdtlppVw9SMFR5/4v3jFUpqdKJBcQzOjaGjWSrfGJ9jH+IF5nxNZgKsu
lZGwYJON4yGB7bU98xhHUhxDByzGDHktvxGblF9S1xZFhAC5tYSgkteQEvqZ
TOiCxXNf4sWWV7cxznEyKE38vQhU1Od7Lb7IfqfP5sirU2kUnjuacXzxZkU8
momxWLeTy1H4AFXof7b1etzTZLwhT9F6pir6mFS+PKuV/okVu9qO+gC4jP7I
TgFVG9qVBib/0BQfodMh+IqVpYlCuGMf4bAijGyI9Arqdc7NdVeVVb1z3D+y
DghAk8DanOn7QeHzhlwh6ZcWQlMz5LSoIajmm3/AumfqG2wIlBqaM2IoNQIh
fGGcLcsXrIrh4D0SnlhJSi5W7SsA0miQmBL+oTaCn9bkDrPdKV12ybIVfOIQ
XYXHlj1mEId6WHfwE9yWgs5ZBT2YHOmYglUTFoHG+wRmKVz7b2tq5FtLf4Fk
MCayRHDzpPwnKjmSrb7i8F9CDz6rwJFWtStnpm9eIkTa6OxIZKPoXgAC0r7O
TR4QqgJcPAqNn5UtyvzLZuRN1o2DPgnzRcM5+xamET9D+sDjevY/08jEhC1F
6MBEOLUv8f+CgnXrDyTKvZC/gkoJxwpMJdhUcsI4HVT3YqkNz6uEO8IH6ABu
RxFdturrsqOsVAn3As//dLN9j+kzfqxVfq81hekcdTghlhbWsfjt/kyLhLbK
AhVXxKwbeETKioUB6obHB0+IJeNvQTUclfL5WBwIK7vJzGYr4rq5KT8vqpSr
RuGkTPwnBzSZd4E6LjZ1LHjL13RI5mw2DaqIOB3i0HHiGrqvq1+P/9szf49X
DAeR6qsqIAGcFBlSNgYXAvUk43TPvsG04GiKR8jQmUHDzeWVcs/TOBcdhAcq
MdxMGIfWhEJe464ybv77LASxlgNaTBF//vG3kb58vd+yfaL/8fFSZX0tzJkh
cjr+pb7Ugr84TQJFzP39N4L5uzg51Hg1u11OokvXUGkrzfNbraVKWfTmvhVN
6fvZIEN8JDgzlwaWxT2TzrEPfXXfsULYWLeFJf2R5BJ/yVzPO7irxFH9iTkE
2E3emMoKSqpIb9d2NqemQ1MwzeSQ4U4njNl2JNuwPK5r3KDGwefMT3dUnlcg
k1jmEpzOi/DrDJlrBMs0pxEsQoaSrrZhmpAYdFcz+yRWY148bcVc8OScDrHC
qZ+wskOVYue5+24JFdiCx1CsgoI2Vy801w/9c+3NDtY8tCHjzi/qsi5NjwhB
DZBgovCqaJ92Bh/FuITx0GgsFG0KZtpUCJErHFbayDg+cyY+6XaRIXxpIDpB
bm01vZU4aJ42S5CFm/VyQhPATCBTL5gUFncAYAfuOGYVvNtUY0EvbcVeaU8d
f8uoLNFiHRosfHZv4i6Gmkf+5hrcEfWxxtIigm1I33y0VApMVhYb0KixX6uM
wTcPb1eRiLDzuEPM8MIXdbSs1lZAD1DGf0/aCDjXOJR0DppFMCISU7o5D6kh
WkWZ/UG3+N4tzuRzBRtsj4a1rsTViofYBuIhTM2X42BnUN+7XswjJOEpGbGw
HWw99Qrp/eCQ+ixhrZB+R+F+z+IVoWLlwiEzwRso/fH/6mWIGOwcicPCNtoW
6y88ig9qYFDFUAYIuUANSyjUVpY11GN1NMCwIbV9KWT0xbGVl84gZb8ArJkc
XJKdqxuszLJCjt/KbV1bWCzwA7vHbOvHEJAHhXgmHLAKxL+c/ubOdd39y46/
2SmFg1YZzIFRoDMhFHh6RjfgA8kdenqSjT7sXzXLvcUHIZb3OslZncfdJeAJ
RVT1YRXziUe6BFhLDIrOHyiHX8AvbVQnHqE4ApNvaCiml9TM0TAz9Pa3qyaY
jTaTi/rnbxLPIXWu9wELBdrluB3qHI7DZztu7kVtAH/Pn/cmRge3QiAkGQeB
exNEujw8dUbj6TdsWgiwG5JpP4RG3rrqagEMjW0bjNrtx9gG3W20Eanhnsrc
H0WJt/OJK0WrSBbl4zphnXrIuTv8Yd05yf6zKhjBCOlxWM6w84XWNgYbZrm8
UoZm20qQQa6/8wEaUrLYFgr8eqfJsX2qcfEQkZeTqveXOdSU5X7MatViZKlz
2xJ4MnN6z8haS9HZMkO4bn8bP1MI2/ga6mURDjSxkozxu1Zq/1EUbF+Q9bMK
kYbR+gK5NLSkidK8q3brbeJlPKgMZHOBgKecMFytMXcsGPE/yt1h+Cw2MN1A
zp2lzrQNOyD5bSHY2OV6vMxXGXO89SDCe+GFb3qta3MuvU7ScqCDvkYLn0ff
wBkhYE/xn1VMJerG6NFqJmdhWDHjRTKstu/mlQDorJehJqmT05UrAbRCGeek
y+pjghKgRcWu7cBZ0WxKQ65wmfKJAhXwHpUeajwE5dALhwrcDh6ufQeykJdl
Yyo89i3U6JFkO0hkgDBedphyl8PfrlEvYTH+xmVCAxiIl/HxvRV4XVCiEPiM
mo82pWqcPkuETjPYlx2fko4BAlqO07+0nThd+S+J6gjB+KZkKN+tIiPvOP7i
uKGA5/pGQfv4haWimScbT3XyfoORBixX+4LO1VKGztrBOKzJ9TXeTqbgEqYS
xAXKSZYOMKlBPo7ZkZRk6nLrBE+nZgOxJzjUF5NbGR4aWkoD6kxZPbKy2n/1
937v5ndFplbMxla+O3m0sk5bIT1tk4SjPVd92dZKfewWANTLYdIvSZnr0nkt
Yo+YZNMnCuhc0OBWKO7PmY9akjgVUyWeNMHJIQcKNKPAWNgjG6pxJuB7kddm
anhvyWD5TzorGs8CAYusKLiQlRMXASTzKRdfrTWERkfeMZQ0BfyWfDVGinP2
/QMgHbJ1BXSpCEdArlcfdvzID1dEnUlJUcdikQUteAGZUtCUtfP34D6u+wf1
/nej5SQcfNI+S2wglkrxpnrLUqamZ4uak4B2FYpVHMgMvYkFpTzz+atXz5Nu
OBXCwZvbmgJIY9Gk52GKd2casUYSa5bUIIA+3u2ZBp6UI2p7OMY83H7YJjnp
SXDsp5fqPzrkdzdDWzQ9A1gO045jrjSUbKFTwvi+UIBLXlRXuHvXjqFZu/uc
DbS9khljWvYjm+kKQMBiUAJxTHbH1GHfkjUQsVzRQaaKGA7/L9DIYd9fIABW
Fy26bzSNWcrK4rwlNcTv8wD4WYWUgcmrzTM+aSy8qUUPa6G5X3pY64VhbQMi
ziFiRQtH1MV/9ynVV2XD8ScMbvgYa36ezP+ZVaxbJKrMTofkNKKSvKtWbeIA
fXIyVQPWQjWIAK5t4FJcPHVen/47PTp/8ouEUToqV9Hm1zvZ0A7AOaBSdQOW
ka1PiPA4wloeIUTbuSCPFBPQrVMO40cY7/zOmah24e3AdzzvYLbD7ZkCziRb
cQsYq44Z3rVxJq9qr44I1jAckMvCmwjc9GHOjnvw8m2LczOXOjH4WDLCNskw
8OUuvXKnXpQM5LhtzSeLyLM9ungawWiNZKbW3E1VlHhFKrqc5TW4FEfoIJ9N
WeZF2FYkISn60+ELJZ9H8vGcJohzkQov9VPe5+Rl7U80wHST1Zd8Ft8wLAtS
4EpkUYmxJ4sFGuM5o6mlNUpW2/um4cwuGbvaDZZwSGeOSMyaq4m6kU2OuPZR
Poz+vnenDkqEuxEElTWnMQzxSyRiOHE7hvuX647VVHBHjB58EJkczrPBjE/E
Egp2tul4XT0p+VHgqmRx4rIO9PXepGm7lGCBwNr8bTvUL7513z41OKb/iBaY
ZCGA+JqltuoETmFn7lx6fydS3yBQ88jvjqQCWKvHn6zFWd3xlkFzk4TAyLqe
/2Tq3COPhqR/4Uz2z5ThDJySAcwHO6Bvuh7rRCW57QP7Xse0pm9gt8nKyleU
POMrRefoJHJOWVgqQTsxRX7qkODRhT8QrHXqqYegOrXkcK5xzQsnDbJD5fEu
D74WPKpgPpf7AGvNL014nowo+DSUrO0nsN/aJBtcNoCpJxrzokPAZB+WUzaY
QCQJGrS3mJHHwfmX5h/JfpIVhgEOkbFTekiYZ2cnO1nLAqP1s/RHtxUV1XII
e5CsaXpbANi3dQpED/WEA1EgsR6GV/o/l+4Qa95yPFfWcr1oRE/pSXORchDw
Oz52sxnMY1QEF5FQEQUM1Ty4UC5zRWmSSkMjpUDC2P0+vfkOOJrpglsp04JR
IKRmFshouy8vuJapQ9Raj6KSKeHrG88hS97Qrv9mddxv3IAIxrp1tMDWUSJz
QQc9WW8/ir/md0eqgeoqif/ErgVHYozIVhvKCJBrwsDdOhJGYXs4UXTcuNqy
kyjadgmiaOSrEEfHsrq4rsGYjAZRcZ1pL0oTqKC+7PK0ZMeSNGWqDqb59WJg
Bm/HH/36mwgCEaxYvujirY2Nk9d8TzlOffS4MOEQS39+ZvLDXvwqkb1/BxYC
AyrxiPfN/SkPsWc+WMOGBkuk8xuy1/+sm/IPSATt2FzZvxksjqYQ0VW5sIBe
MTQm/qzLedr9Md/cpLGbA6NcASN60jo8/GEr/yItLKbQvQI8BPnCtHGy2INh
e29Hg1ug5Mcbk5ULbua3FZMkxasrV0Xbxfpl9uchYaaryTOxWRWjG7ZuQpER
WjF5xJbMjnS+utOxUVtuSxXzdyZO6ptHWxFWhiAjbrtnBKHutf78b2lES7Gv
V88A1KYcR3TnRK3/IsTQ1umabNCVnRb+BopvmT3qPR3yfWGCZn+LRcsg9soW
soastsQglusYQLfwzii/cuWQGPanNVLdoeEfu610FEku4L0UnwNjec0xzxZf
XF6XcKW4KezY7u4Lli6ZhdoNaKqqDAweBTCqRZVA07n3Sl5mL4PlkOB8UKEq
JyMiIAqZf1SH3C8Yibd+ydo6HAejHT3D1XCLt2HAS4qYnvwKGSqi/qmNmT1f
EoUxZXrcWnmY1uEbkIVfwDwUUuaEPoUEUUWFULiZjFI6mET28EZ/96MmFCGL
FLzwAeCOq8DG6oGbgav4CNv4osMv3LvnBVFdyrr4a5y2nY2XVbcNEOOVE5p9
jwgrbAkfkoFkO/CoeqWRxkhY4MvlIflg+O4CQqn2KZ7VetiyIwLLPE17M352
odN3039rR08uvWRELsLoi8dK3KrR8BsJ8fgl/UZhC2Vw2V5+mf/c4rk8+ZS6
nT+YiUMHHFHwi2wQMu8I/7u9LQdSqyo83u5H2kQElD8IxDrpMpjD0O9r4+nJ
nXLrcOo96AXZ1Bu9U0X6L02vyuFaSIh2LUQVQ25FHDApl0YsT0t0TLCx3+sO
nyzUXrQmQa2IuX3IJzm0blyaC4cXWL0+qfOVqf0owMs8Pb+IiixiAgtnGhIM
b03CMm76LW641XLyPSnCYsIlhUo8WmxdCpiRmUXOiuo3w+hoshuWlCfsvyYF
e+9BtYIgxjVvODJtlPuGW6em3vXSt+8KM57wOfYKNuAJ0A1KI77fi657GAn1
pCk1QPOZ2xzj9+YLiaD45sM90QtF6UnqJkQwAqbG2r5eiNzdVkqvpnxLva4P
bimA9zEw7iPkD0d0nYgYDRHPycQhgMvtNUkQOEdBUJ7qAZJcuFg6vsO5RzPg
NtQ++2BJIGGxhCoHskISLZ/JtRO69B37Etk9WaLMFYE6dIemm7LsQM3XWrGR
yhJ2o14UbutmOvv+9Dogh4mfYBbLjWMIx/GDWzGATwUuXhbdHIP2cYfxHYM1
ggLbkvBtk4Nrdjd8vFCDQaddcNT2PnQKGv4KPuaZVJt5KrkfjxNfYU6xSRun
1nCVmTcDDg4aC1745kdzPf6uFLUCCzdXLpqMJvidKAJyw1d0lK0G1xcyCuZg
1VLpQoakhiBwzFJGSroqM/Y2+LsnrKS9qrHp6exiFwOthFIyWhCyoGxqoeGq
MbvuAYSYE93Pj9UHBY+PzP66mytU8H1b2aA5WdN1vkA3Z4xCFVgS6lpG0L1G
IwUvj7pfJP8xLOAlL+7Ick50DB2mun64Iql3kF3KgriGI22qFfOghGd1Yb0O
ALrmxAQyHOUUY0paxgItLCjIXTYT4iWLWUe9RXdLd9hyf89BIQmrE+Yjy5zq
ep/LRKgwMTZbPvZdzOrDuHgSDjM6op7BeCLIfeXL3fhFPkrl9vu1DqQ9twb5
5p+LyzQvuMMf1ghF02o+As7sFnn7VFr3Dh2wUqU6pN3gIL7GafTlx1KOYF5B
MBtVNmYLtoFFa9Lhebd8wr5AWOT+3efp/vaUOIv/qrDmQSbYu7GyvxRgrY3A
ssZUDyoi2e5/KMT8I6FWZMgLkvy0LO7aoqiTeueemkQXF0PrqEGu/qBH83Gp
MWxGkWgmYERnGJWatzlIYdDru3/XGszYdCV9RwoSwSCsxZxlxZuDM6j8MqS8
Mu5dLSin6JoN1DSJ2ggODFCKoEJmsaFcUnRBn1yo0k0y0ZXJjXL1HlxO90kV
84ccJbbIh+BduKxjvyCt9gbwkbkda+ZUdZn21EKBYsKTcHsdoxvYSL9Xc6OB
m9Bd/mNXPRYOjQbepA0C1OsWMqnWoGYD8XL28kyIzNbE0Lyao6k36JUxPs/l
4h2ATFXAUslHYb1yxcu0fHodDcz7uMB48v4kjUmWkZ2XGIJ9lJXAu697PvwM
p8n3yeUrBo2b19leX8ebJpZtEHOVQT2aQYj1X4bjtLPxFcy3E7Pek76Qa+Y7
J29PowW/3MBwKkXUKDGQBWGxt/ZLhgL0Og6sAXBIwnj/k80o9pEHOqd7TEZl
eZrO0y48Y0ofWtfmy4czri1xj+nEKh+Fvg9EFyOsiQ2y8dNR1YsCdAA3VfhV
uAf3Sh+O+TiaKzWe4xoXe81ZyFcSW7+k+hzyLqY5PxeevtIOK1DacCvKuRnO
/a8YHu04TdYE5fZ4is+PMM0jzLk3vV/vRtksMa8l7YYmHoyVxE26w03LenmQ
7tMGW2SNADJ61WrnlMv7O1/lS4roLXrGYaGeR7Qrqr7pbDM0fhvCm8FaHrwZ
qcrOlGrMk/qGEi53Xscl079v78KC6A30tYHmuoV2vAfdfsFsEm1fWPbL7YCv
KhY1NWfR+GK4t4glBdfYekPaNDog+oHfOv9hheMSn8e3JtZDCMBLbpenjnE+
TXaRn1NIowXh70GayBYc74pRN15JE/7tn3YGcgYdsvm0oaXwryqTWb7+13Ml
orELTcXyT1OTOG7NU4vsuLgmydcQXRApYGSaIKxqyUYrG5lAwcTWnWXRzhcj
EsypdGs24qvdwlOHMxDLS1925RgQqi/cfu93tJlqw+89TfbAf9qgkHIGulh4
1bkZ/qfGwg7G+GNp0mQYxOZofdj5mczdD1HYDkQxrsgVKcsBS8foc6k9edUM
NbyzDwAOJZwn0XoevAr89S+OTCBnTt3xRghu72hPnuz7/WzKfi3DuM88d1oX
nWf6qy5qX1GHB0/xzcuA2eO6uvpA4dHlf73atqnWieO2TUv0tHTfkpva2j8h
+2yZEqJWBjgxW2JXQAbjXQTj457HGbvQ6Wnl5jTznQwFKo++4evVK0KATDO7
/IfCK7bXIyoZRzCy02AgXGzECkKD+Ln5ljPOJfkbxG1qmL4ZpfAA3KoRDnAy
Ml8ZxlFddHezLSbRkSn92xnyF+V+qASJ1745VS0/Z0fP8SDL23iIi/FuLWjB
oE9E++PNORjoARiUDsLXkBbVVAPC0sfE5YB7sFSPHu71O/qAAeLz4aDoo8VP
Ldf0GZuq1uUeJ/eIUwFlEEgcoQlaxtARpJzkieDcChQ9KHVNhGF8sZ9ncPH1
UotfdjB0OjDADQVeaSzA414UxvOoUe8e9DhyvKLL1cLd9XMm06GavHN1Wdqk
jfQ7Gi3mWPcJwo1sRRyZY1GjayP0+6Bu2qi2mJzWwLlDv6ZSFQ/rHj9RpxkE
DKqlv14p9aywQ0VSdykX5BiAA3/2FNgC9vlEdiPnWDfwweIHaVqZtOavTJqH
Q90sdYIVW/daKtjHuhYiNqdvn1cMGpGzavBZNIQTOUsk/Hir7oCD3XeN8CBx
jPKnyUH14xjuwRKjA/cyREmaDjh2zzzLAT6q6nWT27pGJEgvwD7fL/YFv5Y8
pDBTxxUQnVBBgQ4s4UiUO4XJUxImj93773xC9x2wSnGoETo9IngLpTzE8V5X
wAcnvqn/s876aAN81tOAG6pCLPY12HgSs7tsRyZSZC1Wcbfr++wHVIFTDO1b
lJKwaCXPhP6bQC4JPoBv9bkcmbJ+AUCA7FQ4pfFaca8Scl/C+jQqp/ZQUr7l
cNdmrTCvGM33nSa2D+AHjPhY86SkkO9+B6/o2Mt1YqSoJSR7t35/NcADqHXs
ReS3nFfeWiSCuOVqxicbKcf69OWDtRMs76D+MqwaBNeKdZJ6IGUzjSN3U6Ir
2khKWa19gOTCqVhviSw5/TsUpU3uWSlhzD1LyZbUAOiHTlGfX4Iz8z6b/Nkv
U87jrOSOIazQ90Wk8NiDnPJOIwqPjd+Q9i7XAWpTtXpJznsDH+OvR0iWkxbh
KnHkcDVIwsuQPTYNTMty3oZMDn2BAojSMk7n3gkoJ3AMjzBxg4DnPKmjx8/0
cVOSruO9WcWY/TgBeJrB5qDKPAau+3ayY62m4nfatjJ984pcdVZbKGtZx9Nt
aG9uG2aCXqDsZnVvznhPpBhXPclAi+tbnhIC//Vusnfj/tUUBa7gVB/f7QyR
2MDBPmpc2q4bxwBgyvDSv8lo6ynMCZQM7LRdab8QF375qgAivMkqiaJ73Fho
82VtWqmx0wpMvoeabxV+xoe1mn3DGX8/5NDIpUjx1hu9Wka/jWP0CuYLMiMz
fGi3I+siyIfbQpqwzr3llZPdv2xBT6b1uFIWAZPNy6rrl4Kv5a7bAu6Vhhqs
dxuRcmWZbpBuGWYKmdm4fu7Ug0YUEnrLmDGXN4JZro+umGrcKTqGVuepZ3sg
EX3fl2LlK46wyA2AH5NsmIhBuXI2b1bwGhQmTzp2XkEK+4HV7bLBcWOlKY1v
ou4RDZVuoqjwG001kzFsVdCTfVzXKFtGKDrrvH6KAplYKLbeO6VIc/WeZIzB
DqHrlNybhpT07wPAsXC+7auPko2bQ/wm66W5o8wmSwmkP/FvgPiWSVO5i9KA
mrpIuvMTGawOmW9TQveJAvePiTlGV7+2gsO7RqwRV63Vsbacf+NL0/X7Bb3R
R6xC+a7mLw1wF4NHY3FjyIgXKL21+e72jH9/E0FNvtq7XZpkcRUEUBJbw224
pNlDAvw7sHSlC7wm4WdRSBKEa2MKLoYxQJz77bizIHrsf4Hk6ERPYMjMvnY8
iIjMmajcK0H8CdHKwu2Hw6xPiIh21KsgRpuDRI3lZgQUm/y0afXU0fzWWImZ
hnW4V/S1urrVIodI8hK7Ge/u+F3lIJQQD27Wpvtcp+dvlePlkv0lfBAGAq0n
2MBa35rxpE2e0f/aSUzLuzOxRJqV7nPp6P6i5PPuzCqmN/CCpD68TB/730sa
qUev4CXiEHMc0sfLpVNSrBdo0Fo1jggUL6UbFFYNUNHoBRMeDiruSsTsEF8u
+mYcG0DLJiBWT7UxoPJeHzCIfL4TRRUmV7WL0KCRXJRCp/+4OAApOAPoFY7n
Q8nVG9IzDGLtUD55LfZNP9Jw9+ssUR0TeYbzLCMfCmbyb2u2KSoThkJ0LfVG
lX8jpTgwXSYOcS7/3tYbRIdwLb8KvoTrD81FwD167dO8AyVX1wwxF1DRgwW/
RhYZyNUElm7lCjKsPYmGotq0s12a+YPE9z079K4WgVyeQmXYEzblz8TxA3Pe
YIBjo3SP5PZ7J2zQnmlckFDAEmPNSyWiIyHnYSaNDebTjPku1A2u8MPOS9kM
5pIq2cS17j8kj0sM6fEykOzUYsW1gvvXgKMrK2JvTzfuh9iXd/M2W8yTMrdn
SiOdJHVy0r3MkbgqO5ahH8j0tw6jGDoxV68NyWqw+/S7TxMYCv2a6eJKK4DD
CX7OPEipILtEKhJ+k2ATvCb7kI7Ts1/F3kYEimnybZtFazj0mYtnkkQ5MDfn
QkGaG2tbHenFLyaxk26aD0Y/nkdud6E1FtAawBllwk6LMjCM1L7b64rwRUsp
SRlQn8WeWX9J2l50iVyc9bsZQ6HE6Oe8g9Q/hGa2f6GWCo9q6Ku+XppAnL/0
m6GV004FeOPQ21rtnjMNizUEL18bo7H8Tqesx+BK3RJ/0I3jcXtTvo0NH8vY
u3EhkYVzvhTdWNb1cPMCXKbCOxe4zN/kin4fvg26jQ21rCo926mtfuhWuQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpej7iYrjgNRSSh27fpzBDMn00ZcR0kw9kgBQZXKbqaK2CdFZa9cVNrt7FeCQk4ELa6b5rQ6MMOSLkmV3n1PQ4D7Zf8wqEhGazv/eX3ju4I9Om/pHTmGw3hkIIiI0IaxAe9hkQfYK26qR9IWDJdWrZ1xSHr5dDS1BfBONFt15+d19631JgU1+3zEq8PJncj4m1VAxSDtyFGwVMIZW/3Ba/FFHWxM1GgtAdSRf9PgltOrib0ND4w+6Z6IJ0aUK8Yk4+//LHMhW34ofiNOPBeo7FW4WrKg/PK5ijlpp0RNzoMAw/G8Qp74oQq0Vjh1r8DzKW7ff4uSxKwvK9Hyo7StJ9aIt65QLYZCGMHXARhoO8TT/Uk0ElodtEPzEGzlBNnIE1ulNIyLQuwJ14F8xkfuy2FoEWAhuj0Ztcc8kNHsTqnpydTnOwuQCNTtemTIo63s/lLb+/jT+DAwt7nx9hroC65NhzBQTAnpChpgX/WspAS6DHkFPX9oMVSnQKJKcZO41zRi1X2TX+PgKaOQacfe8V45/uKOKKTV1qmiaom2xtuY09raexKs7CYXGGoodC4fD3O/97++dPPDUKxRwSvc6cmHulDdNwppx1njPCX5bxnmv04GJ+FCUUogFHMZkgVpFq2U7J+hWtL3Z5xczNzlcTXTfNAJqFshumJ1bYjHpgZDvY9o63mP7x1AKuAfTYNvM8O+IThaxIBkiqGXIUEWcPSEgFPhE5qa5LK5UjChWvsntqCRZ7sZegCT4IJIBBYe2aBQ99LH1+t7SpVHPASx9NPxM"
`endif