// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kArNnVzLYCIwoTm0NBZUBbNvz58fhIhvSE8RRRcZD/JLBpZHAfk4I3oFy45E
Q/kiQqcm9XucDKw5d+u4NAwUmFthIhA9r3wyNwDJU4SNwlw14u63p4RVTJnv
lYBzKE3RKtIw8g4/3JKxoFJd+yXVx2QHCYpfcphsN2wXbUaObQ+Ek6I61HVO
Zojbu8vkpeyERp/I27+sMClzzGfKFlCy5Gb/C6j+7PBiOpi2M9ffa0kOtzM7
HvJK68yizraWb6TeUsvyTWgTH1QM3u33wT1QAHAk0A1wMOOw2nLTatRx1nlr
ZlNuQGdLe7GxV06JWjslcuHuYBotRthHs4XLa5Sssg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bpy6bAKWhefLenBGzcedlIPs7uUwSxG+/JaONqvhZhZkTdhjiO/51KuuikoG
r/IGOS0iw6JlEHsoaAu8ehGfpsECCiuks5xaDEJhz/FIG2wqKz1KEc+mcoQR
y+wvu6+5zuZOOxTpc0UUgUVbyF05uHeQ2YbGguuzzPLZxbkjh7vkEO2nwy6h
oUwFQEf8NaBm4mUZ1DTemVZ4CNWtnymKmFjNPVBrlTqGdgJC47jHIgXcmYBJ
soPvF5/7VyG5TDTQ86d+ktZeFUo1MXhqr76oDxCue7gr6BicKTBBpdwPVBgl
DO47pwqDSxrAJ2w+Cy3LEcvYaeOidr1Em3NRs/8D3A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
drT8KYKzjVy/tLPE5/t1W3yzcqD0qSthMq8CGyIOOTRjMP+tHqdxONjTIgYT
XgWOwHp5s+3xGZ+z3JgrjU0Qc9Jb81J/J6EbbjraCEoJRsnynp5oh+MPShHK
onpelUjBvieqippxuZEODqepB/OsRVP07NLxXetlHrcUhByr4pt6/EnNGPMG
9ZWTbPlPk4Yu6QEFFtO5168FT+JhxKKQWS6qGYesrckdmz2i5NNluGTeC/9G
OwpycBftQm25c3n4ppfA689xEIvtdKT95xty9O3KwK8oacfWb2SFeaC8ebsW
kAxgBipwwgwQf2ary9b9vg54y3DX1EJOqijYsR72cg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qUP0rLlPlvjaV5eVuIalAnaKTY2QpeVLcXZzYglNqDewwdnED9YW0eUZn4JB
WRM/R1RjoiCJpgpgGmIGf6zn/2rDdo93SSewjLekILUccyMx5Gt1uPyIVVhH
WlKWg7alKgXS7CQdD3o+z/Jy4guC1bMi/+5VS66h7OCIiiZr5kVwsRuQevxc
KCoZgLAnV1POq7lMMsnHyNjETFejIXoVehFJJpldEILjH8pikrAXBGXwizis
LwKaACdwrSkSHZ3D9i0qsl1sDFaxsgjYswTAKh2wCopsPwkS6cvtOGIEzOom
z/Hsjc09M2UWNssX2VHiBQfN2T5Wu/ffxqpaq0BQXA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TlPxYrBIzkDSMvFr8dHm8CaQl+56cgnBqf4DAk0JYxa7MSCjKwkYhzlKzkWY
uSOdO2xu9pL6DkrQWrLqZ/giRXZiGFOByDWbPrj/kpdfN3GwH8ikeu9rdFf6
pXVNQWfwRftrSSJM9DWIeyFXOTmniVJKf02X8XNWY6LqgRpc75w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
q4sI5JdlP3hqdtDRngie+8mvvrVLNVI987888OAdzLOFPw5K39hgvVRaCbci
grA0MRCvdTG095UTJXTb61YsvpLbhWfHgg4BhlMvHjExC/ewp/m/cjLgabxf
/Vz4cV2P0yyYokZX7YU4v7h+/QJHSsTbe5QDw7Lstlx0zMC4aMKPc3/ogZbp
HFG59oUekaDtRAbUpocyfb2rTNVqlrocHGl+GDzjSH8bXJ7jC2RjCMzmWIt7
MbhreBEnEXrF5BHyNwl4+Zgt/umE9Mwb9j/K0YeCiZzeZEFIvNc57s9c5Rfj
JZ+PjUI+xlbBrKb8gsvaVyT2WHp0w8UmKwvF2f3xNS71FKXAXJJ+2aZNp9TH
myZJ3DVcMTWOFGzALI2HX0K0HJnrsx+UfK/DJne8/05zezbhlKoHEEq40UfY
qRZNktJn80FYpgfSWSQKQgRDMXchOySDwcUnGYay/dvICBoo2uSCcCvvuoA4
uPYXOQ5R7g59FUpW1OEJt1BJ9qiHtuzw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BQykhutobv9oM1Oe7PzTLOYMIo3TrX5a0oBvooxTqASiInthG3q1ffaoVEo7
OoAAcHULh0Nm2ezA+oI1bItAOzzzNYUI46ENHraeHQOXt2AGqftkUN1YjCsO
+ZyJwBwVP00sWOXZKV2PkDrNkgedB3hxeAfHKwwgo/X+4IeBClU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YJFmF2p3nMRfvCY89B7zsMcD0ZEJWtg3nv2Wohdi87X5l3lgosO650XHp4jM
//bXKS9BkfHy5McElb2na5CWWJZ2QTPmnw5jignoaO4g3wUzu1VC54ld5BG0
zQzwwrHNxfg7bLyowbdO3FtqB57jWgVQzentqojyZZfmuYQizfA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4560)
`pragma protect data_block
J4ZfjDsL+bRmiTUzb69cArU4bfITpm9FnZfQy0iWso4nouz/T4qlMAS3vgQH
JDTBmxpEo21U/EAwqJKrtpOX1KdAqL17zsRGl/KomH8Ju6NYKgN4oqopLFH+
P4GivBJE4N2ZPKGrfU/f8HfPjJelkdp4VktqctsHZfV/OPZ2tjpGBrFPdsPR
iNo+Za8HeYA0mc8E6vS6fXx45JZRdF1LHul6Tb40aXsqHJv1kX9GdGdRuV2c
CqnSf+LW8uDHX3VF9l6nWh0DI7ZrNGwXUdCbS4ZLkSPWuccerBl54wFqtAHs
LpPNwyS/hdKHWITNnY0+3ujXQy+DJa88V3pBlDGvnJQCBIGmAL/6V6xPRBd8
tS8OLAR30yrjsGw1i3G0UM+Bgcf2l6v4LrbbcgHW1BArY3LvXzXXGheh46+n
zErIeC+J499Z9Peljg0Zn1ZV1yEQO1e8z9hgZf8Dn1/mBQGCDLxWyLLhizVr
Pqt/R0GYE1Gz4AvMuWSf95lj9MO8V3uE5UL/+1ZW7QR7j9tkdnnAFJOLDPBW
MHAAegkIYRy/yeSTQClWuvHBIlwdRllNk4lmA9aDtwCogBWZ1yEAaqoQ04xx
+y9cGio1riUIJoqao4P3UnBBBCBykSwqxIMB4Bx5emsJkBqM658I80n4k/rH
1ek8mUKVV5ElYW96C0ET7UoVRxtRk76eUzpvvWuyJPDpW56x735ZaWIum5TZ
u0YNlnlJpXaNLfloyoMN1vB8aH/UvbqhLwcdfxqE7bTC9f4SZfyA4ZMDyJsV
THEhZ1xdBeXzlgVzPCbTNPIqklh4EcOa+D2iJo6YXCHxaWcthybFagoW/jS4
bnO1xogM+odVEdsGU2382MQ7Klz2R0gyxSX+b6bR6v6ykoUdJ3YKYZQa/tco
g2pi31i0HIIe8F7ATJHw9Me9vaQFRm7yvwaoZT8fZU6COC7qXJrJSjVhI4RX
S9fwAqFMlUF+0wu/F5MPCLPqxYRRjKiwNXXuG5EM60Kewuc6DEfutt5k2PBk
cSLRc5Y2+O7OYpK4UZLZ5TodYfIpMHXSM7GxLro3mS9ViCPMEPhJeMlyNTJz
/hR55EAQp6RKcPcE+KFS8PHuOcshvdfRotcROjLeV1p/Q+GS48r/zk6WlYWx
+Fv5Q5ZgxETMp2sS/0HJcBew2LNatAv7sox7jUagGpcbZQfIR7X7nhduJJOk
LoXXJ78ef2v4HMrQ8FzHH1Hsa697rvSYBpuRaDxMKGWeX5Y3DXLqRqtcbzYM
RzwpjEjiBObR+/zrm/kEQDBHOQy2ml75v9IzYHrUevUvyFCxz+ccHTnESHt7
nP71BB08N7B9Kp1Zv60nda26oaZDVnAp3quyYy4t21dmyBtik+L24Vsj6aon
AMn98feWJNijIX8yEVmfyOFJ4o8N3PlcrVtanCdJ3654Ne/CIWsbl1vz6xSD
YEVHgsc38CVfRmGiPASxqFNFQlGuVLVjTMuE+ZUcdFUp81Bm/CEop9exuzDg
4+oIl45aOZ9n+qV0ExCgAB44SnAdl+KBfMnCr6QBBt1avOtSM+soh0X1rmCY
WdbnMwuy6cR0Q2JfQo6FWiBhvgqoOP/27t30i1cn1nZn+jfZwOsjwSfq35X3
V+w2cIcpTxHI9XyJ5eCnIdmc9xXc1QY1mCXn9Hmf2InJ49LWCwHpL4PCKQFN
IPDYN40MZ6cfIerqveDd8VnYIImuBHVDsrBwKtmXoWp+1J74X94iMX+WS0NC
L55BEgxAUDmzECouLkg5hd7pZ7PiZ+7fxAWV9HGkJGyeWn893SZABKcsYaEK
CzXhtIqqtMbysOQoYxIRvNY4rvn2q3UBtCBm+fCeUqtWWdwEeltHsZBhj7B9
c55w3eLsBEsuwtU9KP1NxNWHmhCjY/8rk3P8gYupusJoQG4WCpFvIA4351ud
SpAIpYH2DVh4rJXsFRIc4rhZ9coOAgC4e75J4ueXswuAYME6sDMQX+1Jq0ru
FOKezdNt6AFDxV/hdEjROIIHyKNoNzUUA14hgxgkcWKzc6WJ+y31m7lccBX5
PRRUjSPi+gy41xwAWLLwloMWAhTAZzYA2cH46C/ppTI2HMWCedqTeH2nS/YW
wqKusb8RU0ARtJEdRYvpYWIvN9B4ph0L5MY2La3QO36q5S8B9MWSdSJ7cp7f
743fgDtoaXs1o+QXfzDxmObl9lFCPkvOZ6xnU+Yd5sO2fG7AHXnVNPGPVt3g
0YVKDM50fdDnXAIfVngYmDehNBrhO5gn6v9k2+d+7lfdhCXW8mzdDLnhcDLg
7qFbtczT+Hkzd9Wi2vHsAcaZFb4iU8y991hBt/wertQcVmyMNwr+FigU/X8R
ij6Gqy9QZXAAhrINUzfIu9UiEn+0mXjq7fsrs+d+ent2JIZY6i9AeW7tQ52+
rNdFTpeRfgxMjgFBrwwQIMwu39g04mLD1NQmxAbn1Y9h8Hujtt8f36RU7hSm
BdnXu9vPBh2a2S+5NSfEyzl/jq19NJFSU95AjY0dMQgBPBl6Yc5cjADGwD7x
cQsEnBVDTo10oEtXxcrU5fKy0TH8B7gsFw7aNT59Ag0SFiuEy23DsiGRl4Eb
7hggONRA+ronQTAqdtU1+u3odVS9eYC4OuXO6e1sAmMhrZZH9BZYznbhIKTE
4zWVYNy+EIUoBiB0Rr0zhWsDFegA3UEnKFeeuctORLjtyY73trlaClZbB6Z6
Jw31mjo9l8FcJUyzEkm0Wga82594jarWlVy3EfIdAJQ3Iqnz9CCcXkHXdFzb
aMKdzTX2KzhvjrS+WMXAX98LT3MQhUWDzz94fDMKr791CbsS/rgLeyASRrAl
bJEpPOjRBdwSGsIbfTaexwmy8jsBFnKKYMjjnZvbe2fsOIc35KyNWnR9f1w4
FkWULwUxBZtrzdGM2FYfmjGQqXS6GXz/zT4y69NivySZ2nVXyHJTVstZ7DlF
0aY/FBr1jBQpKQ1Z9iy5U8LTh5BRdWqN58dm3OGKeel4eSrNK4gddiOn4MRY
7CwG1LJkkkVc0Z2/4EmfiIDk88H6GIGFFhgZrlewVCAnO0G+/2+Qfowaykq9
wcX+gazwtBHfRg3uXr+J1ocmtir+86GPirlmnWu06hPwHdUvNDva8EpoPnvV
mxq6lLk+p+eFg4/tgv2a+deSzvyfvnyrKRcG2RGG1mcUkCUxego7nnBhvilE
KkHjB1a9NZnMmU0CC1alMUcJ/C6KMNHHhREkBFkbMx90PZzqu/tQyWdMqATg
Gk/NVMVfQIcKOrLYhagFHS52uC86FRgcKr8cebWtHfLfj40oli6RRMWGNHtG
LuUeqjjYzZoJvJ00Hdqb2T1R3mJM6fZOIZSDRyXSGazfoua9kSZhvIagK6TX
FG4OwYcgDECDM/hL4EBfnKowY47i0WKzp328ZuQLpn56jSmLi7YOb4WRajsI
qX9Ur0dMfsxo5+MtNcCS+xHmBcLYKjpdH8Jfi/+XbsXXJdTwPfr/CH1KKjnL
7lw5VtnTd9qsC+sVc/jDF6Qi2r8P5AsSe1TA6cNKh2k34cFvP8oX0EUOnGCY
hmtOtpn3QXJViT2yJH36Crc1N+b7GwkTEjjZS3c3hbfOXNRnEctIKSwrfAFK
6xsl2rr3MXg7n0PAGmKPTClH8vcTkSoM+6DOhmAZYj/cgqrTU/IUu6eIqas9
Kqgg8me9F/1vOhNKKMKsnZ8O0YCH2+tfLJHZcrs4YnO6XYDxfPwpaGoMLmAS
GarCaWcq5ZLcSDd88Greo9cgzr8d5tenlsQ+YbhCLlNwLQcgBZobad5+m+iN
elyNEuMqfwVDwN42C+vsDFxMG5lJ36EBsM8RQNtF7N/3NRtEl1Y/kagaFGkX
lgvkGmQuYHYOcWSWQFK//LnczxZXdf50b+IvkvJso4RE9EsMaqF9TjFcNsZr
AWzo/xQaBRIjwsSUXumdL/nwjCIhUBVk/SqmTKEuAHJVbxTkmaJ7E1sN4Mdn
amkgRJPt2XFhzzemTblN6/A+ERkXElZ1wbHN8bg2sMP+6DlRLBPGZh0Qly6X
B7CavRaamBfGpbZhGcjDykN2dWBktuKze8PTPW0Wcqh6CSB9gLDIWWaHstvA
SqCeDEEuYogOCcw56tBRO4c0Jayti/3JBGHhLi4n0u5GuUyf/paJb69cz9tU
lEjtnXsPtiFTvlPewVhPA7yp31YqYYGp80pe1HSTzQ1nNP+pRA3ct7BnhHGd
cRo7h8QeARr3T/mm1Ynmh/967ZxQbI5hKh2wQ0iv0CYhqekE3K+TNQk0uJfE
Knf9h4H+z0TeMJL1VJA8Qnw2vyXYdqY46pfgAHC0rjGYvqtSU/ftQxyk/g7B
oP+rDC+Em4gZu3zpf9d2drE7lXncd5DO5h267XqQWbj8YUMBTFzgmmA+lC+T
ScohKyZ3wbs26T8VuMr/w6TwtutOcBK68CpfPv9tOPQi/IFAbT1blofuWm+F
uWpKbf7HrtiTUMyAZLW4ZXxxkMcDB7ARGxaxTTs+CwtXjNv6Qq/HEaiMz7xQ
OHJK6LLKIfxmPT5/x1x774jG1T4iMbr6jGxPkuMscvSWjnx2vEc+ETRkTpMV
EgcJhx13ceeQN+eee8/E0cdYTpTn/C7jhnTxSp9edf49emywiJSY+FY4C9w7
B6G44ms0QD5EdvzoVGlyoRe9YFQKV0zZvvxLNWEvR6UQ4gis7O9bHae2gRqj
hsvZ/vYg4w5dg6SGfl22hoQVhpMYXx9CVXTKPK5KXgWlSxqwDbIy3+kUUXUg
zY2kF+Z9ClhX7DQ5qbGmiSRmLLekgNUEeUP0/ZZVLAAoGuzbAhygSBMYTpL2
u1FuPd9ft9kkPT+K90N+Nw+dwsNIiQmAX0iWJwBNpRzNBOE1HIJk1IrLB/v+
NEoZaO542vmAMH1cFcHZjW3ACCYEOHjG6H3n1GWeOWGw85Ct1o2j7DWPzCZo
1mlVhvzf3OVYcvMTGd4tYHKmCpoO9y7alZBdWx2aoB8gsPc/vnxMJ5J2mEYs
VQxwKacM4w5otans0k+G66vWCoca3IgNG/4J5Rx9aTeghbHDV1k3bU/2NQ5v
HCIafVe/8c7k2tDyUU1mWagBp+Bm8RZ3xvNonQ6+t/9kn6tmSx+r2DWsmIxi
rq+khOw80B0FoHi1dI4BwDaj76d7bb42EIHA8WQnPlp+y2CnhaAv5JQMtZ7i
8c6el8V+nFDVUZQ+XrxISq8f+H9UX1Quuy0YhWzHojSQWvGyEv8YegkLpEMZ
IQ/NxyR0wf5kiVoDr3Eot4aNcZ2rSfCoRSCFjDqFrdT0WLB4DpKurzRW8caO
zvgYZ7hkxzjAsvB38+2pc6Qi8JAIKeMrRybGRexiUPj3MwrDtl0JGCRunDut
60tGjRr4fw61s/bptmcoDEE7/ndZKPkLOqm/8tP3vfzaak8PqrkMHndqvpNc
1fMuBi+sfnuPvHIcr8dmRB6byla8dabHwegmGiq2774gUah3Vy/vjojZH+6g
qcbK8LWrIZc/7bv5nJaer4Ay3P7aeMK+z14S4FrRaJXUd4v9Lzl76Og99F9B
cXJ8faexQa9Ql6WKXdAx0rTvhbtetKwc7RlZnk3TaaE82CsfZqBQXo7VfYI4
zA2/sb4QbfuSKbguUSrRIYYbZ+klrhgy75CL1X4vb7DYi0vo+yy8iYE3Zp1H
xUSJcSFd16BthXDHcR5a37ZnzOqxMl7q1rAuk6Z6vC8bg19z5Tp/QtnNBKK6
0/MHjt0C/37FQd/xMAU36kSaryutiAsKYf1A6ZzGjSSic8izFEWzGxwXnxmS
lFL7WBGg7i20R9BgqCVeYC82c2yrto9IvKBKRG8ZRMrKG2fNp+OXr6tYOz0S
9DezY7ySO+TAj9PoycQI0yc/cerZ2ZbYhLRaJblHEuUav+hilSQWDYXx2Mwt
4zqv473S7bUvvFtHqRg+31WWg/x4t3Pxt1QGWzfl46fmYpalEoal9hAnQSC5
NW/dsr2Tnoxt72hyCiYAP8B+olWM9DeqtPbRx1G53TyVlMKmhFGsupWAlSg9
PQOq4eB5t0+qOHIWTHat5fW6X7zx2JhIRm47dZrkLOP86yUtj6sxMN2x1s+Z
ymYEKXcJSkfi4LCupolZ

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1IlxzlwAPBUL+wFHonHU5HOj3SmQ/A6ZkQ561YMp0rxV4JFluS65AhMEMB/SItpnBzt59BNQgPRsklsWfl/WXQomXqWwv3S2lfSxBibVJESBhV4CDZ2wbNyJCo/KsrTHggNkKkL+AHVAmcp/szk+Ga6lldK5c54QbUnzPm1Du+67qrI+n1N1wKA/+tbawD1jvUHdLctJN/AfsjtjGaHmRw2pEC8+XrQmxH/kIkB7XpiElAewKD/4Y1ysHCV0ZXbD2f1zWnqVbV9e1YjW5y2C6pXt9E/ZEBbkxTZculbFB9JdnngGxOD8TeP6zDHL0FPo1EOpz/knFW5HbfnG9RJ+u0ZxAsl5SgPFfFjgxnJ/5PXYE3rK32+aGduTNrkHIzDA6neW+WM6aQ2Uddv+095f8eDwHBIgpYN2p6bnseuBCaOYOuiIi9ufDTSEk02deqnt10LbqyMO2twRfd/pyeWnO0DReEZx5CznWyypPa7ZO6prv2EpfZi1u2zGK5CKFz26MZZbMU8Su+Api2BybcnIMDW0/zarbWTTt17nMbU965C/kpa2K0dHYMYznIDRpf4ir2ne5TdCS3mYrlbaO5FBTlXs5orm0ZiWTeOkIq99ukcC5CmGa1Jg7i/l0KYEhIcCyBsDQsvq/h0h8IQzo/l1rCvenWkFnJ1H4BZAeP92UPuEIInnudJqtg7HK8AY0fGQ2efPrk8anf+7F2f61VT65sDbq71eVnZDEl1dyqK9kLjsZe0Mlf6KfXgEseptQ84Y8tGmxaveOgzUVCRSQXWQn2l"
`endif