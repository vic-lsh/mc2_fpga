// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EED80hCH19XApfhzqDdOmm8o76v//6uPLQQPzDcjHKJeGrKmsT3h81eXQlp5
s5heBItafW1dOQ6Vz0HEpgFE4JrI6BLXsUXyEeD9eRrS/tFVsDC2bcNEwb29
2YIx00JaTgJZKkOhz3I4gupM7p6XMXRn3sXFtwwcJLIV31YGqbSF2E1L775U
LhdTlBKAZk28Tl6DCWwmVdrz4VJmIHsZ255bs8X4mlxQrRbe8s3gtFT5AWSP
6oEVVYZRZKoswcC1/HgVDPXqbXYQvhDTREJdxvmlw80YLrgKUIl0VVvg78wX
4XpqrNrsfwSJgK0PuKXZvNsUFtOIKF6O48FHFtSrdw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cOYqZd63Gt/d3c9meOnfMHRBFKsba8qstuUe96zLNN2BmtankqvHK0q3kgc5
kf+c5Sejm2Ox6mwN750qHpFGZU1s9EVhKrHaRB+DBibU3m5RS5PTiXTBHa+z
BmDsI/H0XOpBt7XbWhgKx93UCqhq0/TPp/hkxSDbT4dqQapyUnUtZn3wXuBd
TsynzD6d99wUomi7lrV6/zB92EJ5TfqW3k0rMuPMs3+NcgzGQiClxe7hWxRp
2ZOMqa9fmlDKXMIAxJe8947RByMfdp7kGNii/fpBZUxTBVaVaQvVuaAr6vBE
S55LLu1a/Y1G5On6hfx1UOWnKAWbwZV57xXF8SwdQA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZWZRJu9tGtV60cCiBxGRGGkTRVjY3Z4TN3gxyfWLINoqXZNbBcAuGnMronyG
QRSI3VyFamz+TCCD+zYUT4PyhsM5WCvZaZbJgyeRd0dKz0azLncP+O2LYdRa
d9oco2iVPsXcUPQ7AceTqk6tqfIe1i4t5sR0lsBT0Ne1JWzroMl0ET1f7pKB
9z1lcdJWCD2bHkzx7dJaFpmk+SLwNMjMtN+YgCBiIr4NZOtnuZgSGNwwvKS7
rEsCf1hkDpb9RjQ2vHwlFfLeKw7FBCjumrVzcEc6mdNNiigjMWld40FaT+M5
76sqWOkU+Bs+npYQNiRQRIRqPcEDZbjfkzoGTB7s3g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ewIKhBcLMLaM0JHBum9NGexdqbLHWCB4AYzg/EEQzRVP6Alrt8MU8vv48UM7
AaK0UAK2pxZXUdwxDkifovYDDRD2SXRqXRZo6wZtTbgF3a7l3NBr/iIeyBBO
iF8NVVrcQ6p4XSb2KCD2IKt+U4KfJTj5O3O+E5pA2p4G8eQv4NAREnML/xRu
ION0ZT1lDRaNFPgdbu0RlbC0s7GhfZiG1v5nLz3S8wfN09hDNLZnqEn7pbKk
C+UxPb2MhkB+IifIzTgBPfvEygIsDhSJpYlPVmWAkUE9oF42fN2umH2/GRT0
EmkAKnRetgVhGoaB7ElzZvtPiPDaIPENHxRf4e8aug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DmBvS+TmLK0t2msL9UZ1fEvXyjViVA+Bt3iZb0bnvXjNiwaXEjUoV3Hno93y
ONy4i0fdkfZbEAbUt7O6GrWvkMmdB3Q6JTB7pmNm52cfF26AGkhSN7sYEr1k
vLJgvrxSuZHie2fmV3K3isnlcUXuo1s+3XeOb01KXEinO6JXkTA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YCAPXYh6QtSyWZ3LHOq+AjbtroOSeBpX3tIzOX8reY+glv5WoJM/2w9RngCA
wCCAjo00OtbXOEkhXshjO+nKZMJyqczSKWG+k+k0AuFo2CKTuyPFLT3Jax/H
kOCGMzJtUBMHw0OPM6oWj1Fa58eGdap8gr9zrZLw+xTPOxciKUK7faxLj3a5
M0EYXhiSfPcz4xz86mhUVhxEur1ZWuvU2HcCvwJYi0mN+mLKUEtoFGEKLTTZ
T+Yo7G8k4EA5f4WWWoB2N5KA0BoKXMZfw+401UA0zRjnnT325MK4dfLN0bAl
bvR0QrG3cSUxL3l0swEBFtQRn8lyn/216uO2nUrrfE9S9YzwmwY53Y12G2Kw
XVnGXNKVWuiY543LDGOtoB2NZRQZLwhhpoH62MZY3o8+6axmB+u+apK5uBUt
Llo+5LVGwhWpN9+MXQqjnxpmIaPonozONk8BgV7af5kQMOT/VzoK7QNkawsc
AUnlyti0kVxPQqR/sSbRuZWWzmlLRqXg


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B54EZIVUT/xVNT2CO1PLt+k23H+BQk0fosMhBnCS8KseiL99HHFT8EyiGLW+
dASTuG4jFtRDN8tuTXlrLpVhvvJD8XbxaxEkjJUCaRURL56KaIx/3zRiqrMb
RdlBz0IZgheECBz0Woj9Bn7UusZToTME9kI5e7pE1dFWfbqWh9k=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HHU4m5TG1djQog+BP4I8v6PXbJeRKgUzn3Pwk1zeu7c/yKjCouhi8imuaMNW
12L+0mccBbeQEkNZP15aAEIvYeF+qva6BFgxCbgSYDYiRyyAhYEUhRabzL2H
7YX8g1R+fnChmDEXB8XyaL5rhgkz8MYc6OKB1K12LLbe3SNwEMs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11136)
`pragma protect data_block
EdhbDfe3mKvygg9R+KjGv4uimliE0nXvhQXd9J0p+uh745hfPtfHr+latMmK
SWyG0Ne3taZODCxyz1r0WdUsk1E7jorcJxezwXOP7p5jCKTqepBBMHS/YGT+
cYeQgbgPMZyYJBg4/m4MtKMZhmtNHICPssp/ZzPaK/rTPruOqq5z5vRb5muu
Rjqxo1mbsnHEndICx9VEer/9j4PJ0l6KErTklW+7ggCnKmdqt6vGeyq1Up5P
k6ZJazna61XxUB7XsI/AiN9b3qO67Ik0aHrM9VmsanGGUf02gLPcyid9iIOk
BxVCqYuvSMIehTbIXd2S05xLlJHRyZRmS/aVD1RKltWlVKD4kjvACsgoDWpN
33t/UOYLMME7yW+xTAXJ15r6LSGireTOvk8JkpCGEdb9NATrrYppcsvr8z7P
7yZM58IWb8CSENpMb3sUssnPdrHCGwx7//RdLjTQDe6mjGZ8sageMqaPASgC
9ShDfZr9D1AFF0YOUVM82ElgUkazkCt8OOGZ/i84lcXKymPUG5KKycX16sY/
LKstphM0oeMVBNMZ+AGDdHayj9M/6D3NxY8Kq5aU1XgtzLfvhF0pZYaxT1F1
eIzIbYypYPxdaNWECVixLQ+dCi5B/ifzGhHGOdDd/QnIDhASffSZzQTPUfWX
47qyQIAJ0YZH/eJcGX8NAAxg9yJ3lhezshZWhg5eJnLaWOy6I2Ji5keYgUcl
FIxCYbfFm5vS3phkUhfp6SzjkKeWsnU7ne2yAEZ1TEPBhh5QnBX4ZfAVWibl
brbxZaV7GqIxoB9fCrHni5s80oPAPa7s5JUBXOb4WrvKzG6CxaC6IF5/yPHI
B8colLUAKHXR8AjxTpx4Ad0nVBZN8spSF24rxp1c+X0BQg/r6MpW0sOYjahz
bWZt+d9idVs1MBVKXHWVi10u6V25LAO5DNr2AKMkl+z42gSbWO7oH6Z98hT1
tbMKymSYK6AUc52mkiU2V/kMhuFZyoXoAEc2iKBw+TbbViysaT0VGJUt0Mv1
9JXZBWEPqiEwtWE+5jbgARlZnjq5fvBpKMD924GscPC/u9w98JEyXR73QU1A
dcz33HqexLVD0XoLejGgGa1v1xcQknLuWMU+5gzW26+Nxrgl6QrcDCg4Vq/X
+JAYzFIXf5D96FYojuN+ldY0COAanJ/oyLjEauAFronv/vTQbHWM+ZYzTX8s
ZXGt+933emeg4HdCwOVcR1CjJSvkAUCNyDseBPKBmdbcjJAhf9/ltgbzdWTR
ESEGVdLiE8/fPRJor9aoN1G8VR2jK+yyfuV7C5kKXXT6rFLMCpmR5z1S9qZC
YfnUnFjxeurgcq6CzvskB/AX0w46jNCzQZudTjHnAtNZVoe7C+8sVCBPZZ17
/8a/Jgsv55NThg7/yJYMZc+/eb3dxNQ11BZkAOi4U9AfM75U6RdJZI8ac4eV
1H7rNx37mS+WcHVBR+QAIN0/GTxEgpMLYHtGhhLEgBVT71KdbV5tKoRjvePk
gx2RiBVS/MF85FqTZhIZQwnqZ3683wyepY7elHOcwf5FV7FxiAbSk4+Bfrls
7Y5Ck0Q/ZxUIXBHj4PUriE5b+Z6UQN/6Ek3NeaJFt1tyLGqTln1Nv3cBrSfq
w58hgAC248Znz1lAEh0zAxVQy4uBS4eYeiQWoa32n/cbUx1PCH9qwSknMinp
oX8tUs+MJr6SIc1u2/5S6ngWG+cNc57wnAZeyaa1/5M7tUKJ9BDBIExdHebW
NtRK2c/qK7qlwe9ycGSR9HrJ/zMaXPoY8dv4BuKvO3uthnHb6Z/0JfUBeQBZ
nG1Eggm3LxvcIHp+7XISVhxPxA4WbB6NagoMto5dVhcgwadHirqkpwdVDOH3
RoSMMGxP44J00/sWTDBYiYX29WyGkIrBni9F8JKkRtAepZ5Q8NABXpXC56FO
7fEC1Toy5MteRXSCFID8PaFp7IgIjrTEW+fTJKNG5HpLV9B1DpKWRD2NxBLv
fmbgzxGFeppiAuHUEUKhcpXywlYRUb/yqXLTH4B2GlcGwqsgo9fwBnrTP2se
4hidaU1gUjB9ZprvnXh1XqqMIsWmC8/Ua2JfjdVdJ9QrdXu+vbkjUNvxV8S+
YWpcVZfvRtQdpE33rhzKil77j4WzXcowwwRVKHOHoDZVl1k/sS2ZurTDxOp2
c5ArvBlJYeprxNEnl5OK/Vj+Zz7QkC+ai27JGktgOSbfArH1woMPNWNlfer9
V6QHIpdDMr/enxENgPTEF6b9mV1ew72baKZ+nXCybt0BZOfBFV8y4RrCNW2n
2XJWiviKZwvywGJlQ8FEw+akseryEhuU9zu6FnPlZRfNlYtg5e2jSHj5GVs6
QrVcJo6gE9VaJbd+DOtuCuY1KkfPfkOg8/Wqw0XOGpAU68sFHpSVn5L/9965
ijhn7HXa2MBA4FqnKCdtIK1SOVJd0NCS1I3+izW/ay6XaEAUplngrrdGKxjf
QCz0/XiVaAUvj6HShh/PSEGWm9sCGwvIhlR7kI+jfl9pLagFi5TmeXzmBlpF
rVD+BRfQnKTguwYSZldeRnX62Yx7oP+M+3nc1Tkv3bU8kd+U2pSnURbJBlUx
GfM9bwGHiReaSJ1+VprMkg/dIBgCUceNZhVf8OSeRktDX8XJJkXKgCrciQL/
DtQRUuclUdnZf/pxmcei3QYS3LC7bFcIqp2agFOMGe6IhgJypookGRsyuE8J
C1Tx2Mg5O9y36SbmzJfleIe3ijEYGZh/cnB/lMOlKc2sGij0fw5kwFv+lsEy
ZywKmGhPW2FZqCoOPG8CIYLXZMeMLISBlCPiPJBdWH7Kzav3ZCxjDGTCJDoE
Fkv946zSJF5AGpN+g0vzn/x5y/eezVq+pGS66A7rsZ+CyKK4WX9Ahr8I73BZ
C/gLRBGsCn7HeYKENezl+QgEOjHh9EK+ZiQ0sKASnJ+Gc+ZEXp/nShylWQ2w
sQNpdA7Ii5OTTywIT+ePpa5BzoEMbiDK4Wp+7HZO+pROgydIQOHK7fHmqKAr
BDafOmw7ymi1dKnjSSQUz/BrWMzQ1OmkhwnUgzJfNSkHYcyeI27yvpIx8Fdj
CeZ1ClNZ3EanVXCFYj/Cv28iTWAaMMy2ivNII7jwQ7gx4Ujbyk4FD9ZCthwD
1jMhtfbDhavfJmMXKfDEje39PQTuhO07O2rtFEndKRy3SQxr6YBLiu/vKZIp
As0O3l3KBaDeEIoTj38oikMFGwwrAvD8MvvG2nemMr11KuMzGcjVeU48qo7P
Dmi6Z+wk7QiyvvL3Ph6nOy15QnN9/paRnsi2G8HS3Y/Q3MSRB4MS2w5M90Gt
hZ50BI6NwHiWVVbmXmAR99/sZDISg7yuLp/APDo0qUwhTqTd/WJsExxU8u6o
AE4Sg14TMwbjoBnv0fFVy8h5wi9TCVaKVb9MtlBiMdJRBu0LwHB4gQ8orOag
2JBpE2umomOPanSPMfv8GeFhrtWxsLUlMrkkkdoNIzqwJ3jb4ayhOYUB/IDg
uPTqgQYdEohCnLvUH1iGiPJ70Q5o48x6MKgG27BcKG3NMkf7vl1HkGta3pPD
CAyrKZQ7mt4VClUsU0atEAzUJmt6Br7EFmlWBvbxfrIWZ2JmXgH3imzfVnRa
XIUZNBQip5Bv9qJyZItIAoQLbqhB3FD7r6SDDHw+mts2R4w/dVKaHkw2JVQE
FiR49Ikp+/LQq+1LmH3ZOZx4+epHg7OufMlAWewJLzo+9/3+dLyfDQxZAdGb
FgNNwYA2N6MJB3t0UTgNL783FDJNramhEardaxOPKHGLFnuxTjSZV6SfJXXS
FCOtLaCMbIJ81e3YQnCWwZnJPgccgn00yfD2CxJH/Cx2OSNJWtjw2j3p36yb
WWiCRRCTr0pYwiNPmAqVIYkcq0rwgnm4n8jRqAcqPdhDssguBhkZkj7U49zR
D2VkWFuS1GJTr6OzsLWBRAi8zb3Xus3PXdDxb4rbO50FJdaL3dSRK/sS5LKc
xihJGSfshOFamb/TneZu1ai1cf/kBl75ayuwemCq72qnoAERxMJ3axEvwp+W
v+pCyMYEBH43WTlir1msbPLSTJeFJJmthJoJ/5Pf3qp74smkZkk2OjgriBXa
TkRpzGZiyfXWZ3TuT7yXBjMewCmaFQy1nSMzWEsecZ7VpAiKs4PQfLbRmGa+
OBhYJ9k0NdmohiF4qLhntLuezGI1tMJw2XlRHDbyMB8T451/mfvpazzMUeqZ
o/+bhrkS6uyN1ZlMdCIdgwgqipI8oCQxShvREySytYgbKACDnFiLWyirOP2u
LvsQp60OO9PoWYWvTCTWdtEairS4eP2gwP8/44Qs50o1IQF6NIV/PTaCFFHH
VSloLB97PwC36yHUgY4C/Zfm8M0CU2khSzy9WTsxcVP80vfKe2zM4XxnB/nG
30Hd0YbCh5+aKK7xR4LKgRnrjWhl7IXnuZeQ6RSmZ+r3bpXBLj7mCoIpWeR+
srbYsAuNUUZZMJutokEmXIyhG07P7PxvaLBwM9Nzj9NTzPID3kZkkKpTcgqE
hG95Yld9LwfFMU2vnnQ8iLZ8MESoxDhFKOpbwo97srGxPyv5stqp0wKNfunL
q69ixjYx0+66sLv+BghWBbNHxaio1eVfTXEdZnYH9itAQHibYL920Lh4bwDW
36p9hssWSz2jOLHXIcLcsFEwjDn2DhRuyTr46LTp1ZehWMyYkR2jxeBmCFI1
gEYS++cw1LRz/UjY/gY22A0+M/WC6x8z0K1EpeODx9dbLD3cyn9UT5v5rOQk
IzrPG/j6AktR/u3DGMcNkCTXErNlpH4PDBfjtz8rdOEgH/cy29X/mhcBKX5v
1l8jkLhSh24Q4T9yve3sIQSiuXmvTWpzG37Hgje2bXOSGzmvx0QHsZ8ojtda
P5FZqxCHcPbYFKmWUlL230Odcgqxeuf9SH/B95f7w2xCS0F37crRyq1+9K8v
qS+Y67WicVjHUlxjIOrlnmO9KVAQPQHzlBPmdrkKRCvYwOBa5mPGdTHdXjaj
nY5fxUYeNO+pUwBP/C8MIP+wiwJ+MUepn3FJEa86YV1AzhZrA+u51KrgUpM5
5myy4NqPjWunQOBR2bqhc3uk/weTPNAxBKYNbCwermPXmTnXpBIELlhGrB+v
U+ZeLDx9a0c23OlJhwi6eb/kRJSgvAZu1mX/BiwGdhHR1iMZVREEJfr8QLYb
qmvI9lKdSHgEaTaa/O6gVXM9dLTROuukJ5NpPa0f4C7PPDJ51emYiGpL+HTR
/mAbdZ4mXnWMEjDm0d6j0fwVJWeGqAfb6rlaPcsuVoeLob0Gaa/tckZrG2TA
sye+rfkjWMllLTUfg42Z0j4lk14Smi4YNBeKaWprbL/a5GPxpeX2Jp71u1f6
iYdeWaapvP8pYMjybyw3ytotPZRQa3+lL/dwTLYN7S/viMeJQk3nJey6mcBv
b2X8xWeuCoVah8kHR/jU/dV1AiDGL3wg+JMJvXgHqp1rzuZVe7HccpNUem9I
6wRZNmwq5K6BMlTzLcVDkNaJuOkEO4zZKOoBh4vv9MRPNS19F6q5Y8MJlFz9
JctR/+3lE5mnP+6yeb2ZuWbK4VJ+p8c5dwT2tgmo64m48oYWn6mVMKPxB1sV
75m4iZJmCSDx9549jJ1ytNuo8uIj124ywuvOyQqpCIB7VRxuReKzOyhsEJsx
IMfnBrJMf1upUT5MJ3BJsNyWbpSvHJYNrgpD4TQc9c2MeKBTlKDA8DDAGI8w
pzyc4hRumcenpCcQt+eQU9UQCld5UV7CzrhFRymailwDwWEuM3XaGOVPNcrC
XLazETXRy6/RRVhwfC/iaomzuphcBdoVbklown9pYkX39yEghszQTaaWZ5kB
ErGtCfj1+3mEEtcjgalcYq6BmJHooQJw2nRznNCDs8knKjibyz9/zsNoJmKg
8OuhpOdut6BBYWXZVotBeCGjGxsM2sb+TDxqOFotvnKBa5jgYriwtrb1vopb
suMwJ7rQu1v/Ffj9GKJHZbF3QV2WZA7K5E+NDynMgW2CjM5pOQ2J9ktGKKBO
oGIWT9E1xr7FhraKjUGOz7muio9EuJU3M7JjGI9BDSu0PIaOd6BiWT9cKTCR
Oz6lwnEsXS+gD1O3fSBn4eqoeRMOeJBfV7oBsdLctMWVzgA6GAP+gMuQfVww
RgTTvb6int38ROF6E7gZuLKkLEO1f33FI2FZ+YqR9G4CvleMsFwLLkp1c6oc
2XOPxhT7nUDZPTPe1E+4mGGDRRr8ZG1jVxYNQcRswokykochJh/k8qgWZ6g+
cBa+cRUD45b0jRwMNcdAfj2/Vlw1esyCf25hR7mCYU51UuHQvDceG/nNR1mP
A2Yw9W8xk2aJKvfSRSTzcYm0zo4xwAUxBqb2uQ5OZ2PtxNHfG2fEjpdg1B5V
ZmKld2DCmA7Eu+llkEeVqv7KhsJlM1MxbyX9zjaZfwOa0gf7nmHGlcNbIRLl
K+l+GAW0K+5+KoYQIkUIk9qfQivDl7I66RgDDy00njZCKVX0eISjfRlZpRES
YqmhBvRKHJSFi15MIzHJk2ydsgnotEDLgvEL5O8EnGWwJzo6UzE6OGp2cvGP
dp5/pv/KLlPXmKO35q+w1KDIJI/sHfrvMq6rLwO++/qu/ny1Itns/Qicy0Am
tn28Q96C9L+B3auiDSX+y4NKyf5inXvAxBBtUGWIa8Xf5TFxd2t66m3vSZbo
BU7KRStl0oUkDz4FiTmUHaaPWuR1ztK3B/GgrZdF5oRiKxOzWtSF1s+iLv+T
w2qnY1SCvBEdp+7DrzizNuLx6Vp9HppvD6rIFRZ2Ih6wW67Rf8xSoBvtbFbB
kzlpKbqRuKkpIY1ZcHrBqT5gutvzeREsl/jb29rItd47VRoLbi385IQ/j9sH
gsI9Mq7Y/hcdQBFv4MVUvuedSofY9k1wIDZTe0khDZXkMqSL8G0LfveeBqIi
FAcGu00S18bADPSloYpukL0wDEPUP0wPhRbNtbwqT2Z0UKwJvVzgwWiQt8+s
yK+8+fRy371NG3D3Y+CNEifJDiAd3NZvGPi1zoWU3HKkwt6r6Lnv1L8TOSI6
7JyNBqSvqn39dxkYdK9i/1McT/4fDZCdhtlzTjeKXoeDXdFuwxPN8ljTXLOu
1YEW5VAJt870Bn+62+7x0w5NFS56UauOXyeQ6BqcLLjA7GozaPMlUDRl0zpE
k6A/m3gW9vdw++QjrtTXh8UzPJvM5XaWMOYleKMhSvTKrRP0J0eVcnohpxhC
LXifpi6f0ksBYIYnaRRZyp6OielFQafBbkJyLN3w6cbxrAjoMqfWPJ/oQ+qg
NN6CSLXYttEl+dRjsCsZM4uz3plp7mPr+QmDr8KHYiQMfPIZ8/UyNMEGIZVs
CF/1cEfemhul2DSAOpNJyA3Zzv4DTNmWex2bfi6ipG3SZaDLVGMVSYQ6iHpI
vdAqBz/d2/K4DlET3OClk6sCWc2p+TgljzYcJnG9cj+z0MLdvx1yUKEYuXQK
cw9RtEkrJ+oNeHZ0Z8tXcaCj25CJEEjmOwOFifgkragkSE8fix+HMPWb4jFD
6vsJagfI9sZeEFyS0I+Vdh0MepdwaYK9e83cYV0F3NvbLfBsBlrXE1empjbC
WqyKGQevR9UkdLVbduxlapdXFSOgrSj5OCEFbBk2E3a1TApTzfi0zdfb1OIN
Wk8F9m7L6blLk92zunXmAfUEYay0U6kDUgLnc7A5y3Inbc+mlfqPVOKEAGc5
BQ91pHreBsU+zwYbk6b0nMdI7DUiO/FM8IHh8BJVmzRELmGCqtHhgsnxwC2J
ERYcue0b0p9c9YyXLRwdWrqhNOAE1OF0bR59AFP25OoSXl9jzfvSAMSVvy3V
jitwYvNM83HQ5dBuEaWxuInyzCZBT5UaFPDYxQ2ZNl173+TLMQ2h5q4Ffwpl
/anIE8E808Pdls0L0VHA9n0x/wKfov5TEycvfycENWR1UdFHVtRvYqnbWlWz
msF2BlWUypC9/UKELtTyR1/SqwfJEJ+RLkJkAGv1soGLY5JmN6MX9rEMNEz7
0pe2if9NlQYdwQfqGIU2isYqJ2D7RHUCtG2Rq2X85nAh9F5fpOL2hqHiZzZG
6/6AJfRa8Fs9b32PSyzxur+dPBwjyC5u764O0fMqY+QFXoYZVN0f0kEG8Mch
njvDUl8RwpwBTNhxJ95COyNbxt/7gNfKRc+f1H+tXrvqUNV0JfNlXStmDKxU
a0ZNpR5UpMKv5egnfOH5vx9O6gcH0srIh1Vc/PVsXdjEzby50/PFMf8L2mme
MOqrpMxCuoYgimdlMILM2wgMDUahl2CkN/PDrr5KoibqPSyJdzHFS737NmNR
5PEU81cFegX9OqF1mjpswEH/jVbPgbPjzPsWwejf0M8URHh4y6+Gt5HYQxtI
lT/duImGAPJqzLUYba/MPEbOOMeuCJyCMAo3LAFXQoZPmleRD/LwrLTnHIye
lIql6Ic8wox/idf8Vs0guOaoBx59zr2KLToco3tnLL1cVlT2YtyEshPI8l2S
UwM0YYeE2sLyotc+oJHB3XjAzJCH0ZsEXRlmn6rqcHxD3pMHU6jp8j4egxmq
+IRXTcan2D7hQMmZ48R7eXwt8LC6pvbFR+YywDJtUEBkX4IZkncKFZIoVF0S
qvgLA9ekP25Exq8OgsA4QHyawy5nJF6FEs2hKnJGtJtWWwPwWJrxE6TJgCJL
XsK40w/9d4WFaSfDh6QBAk3EOL9lBSuxxq35EXAsgLQ7NS9UXuICQoctfBOm
2PbZXxbjaOyoj03ot9GQX+iREhihsLlA3e96hU6imEM8Qof68tIzE+5R7rEb
rYvqlONim/8qikBphTZXOjUcmFERlarnmDB9OsWtHTWdYukCXYcKJOIi32kI
deiEoNWAfUr2qlp+j3MRWuOXCY5BpcPuPjfz8iqnWAe5Au9k+rO7620HbM28
FE8SgAciDit+nEvD9MgtSLuM9RaB7d/nKeRpr4ZVnH5TiRQ5ENZzmrPVYf3B
RHAmC5CH+2h3CuP17h+n6Wa67gW73eSBEkcjDwbvFMSVNZ5AioIVZPTFJoO6
sK0Ke5t40oNGJkI4UAUSSLnmT2HYgPpMcMkNVRHs94Gm4r818QMKgSw6sIrd
5gw74WXgrfphjT79DWXDy7q7tQ0zT+pFGB9esTaILwmqAcvmq5JdnrhBCfHu
ZHyKAwWOxe4ww88BZihCWSi6PfBsyj9Lvs3zzdUu5m0HnnRs6ScfwQBpFwTQ
HnDYec7TSmaFNYkF5tCYaavdjE5lK7o8jQKq2zdePC57k/c6DII+SpPnETl+
9Wm4Htqrh4PAleBUwvnKpqClr79lpni0MygXFjB7m8kZWK0PS7UakAchZrAF
aFL3kX3gNlpocOuySCuiHIpYuNxt6qnk0j2jsHEBCYOWOujhwIcCGfQ583j6
kSRGaoJqyT8p6fgDW/9KZELiIuNXnmSgK8ierkFQ3/1yvllD3ZgKdOOHYRCe
OYgHLfETWyBPocNTIsoOtc+7SOnkLndmDyQaPxqSXdrn/ysA077zWbKCk0R0
opdzbrBKhc9gsNWN6R4axEXUUS9Vk1dLs3TQnwC+IC/ni3zt1Hb3wpH530dU
M+DWjSvUGs5dEDIfE/A6J7QqduEf0BCO/jeMe20f0EUbUaEGvSi/EJvFTqSd
bzu27med/1dqumb8HTlEy6C0j26FL8krbrDPnzBJ8HfHBkdYlFm1cJE0QfQj
/1wZnXA1/eXd1VsuY2FXcHL32Yg5ti4P6l6eK9LbtsiVThFLigVf6/7T2biY
5pGkfnn2KfBaeb6KIwiMCmlW4OntiCsgruuwAD59KpMPADb1aa/ISqdZL3Pg
6HYBQMIooBsNH3k7rgxFZLJcUDzqQRqdYPl+VU/qgtukCaYvXwcc02A4gURc
Su+pKhcZ10MvFH5ODJTzXmxK941xncaANytuLXhBc+CRutQ2S+Zwrdbwhbod
C9fmGaeCbSwErg8pj6JIfUNMs5pFxEMUF7xp0lpxej5Q1D7FtmqzZh+OYqqv
ptGQGMGIW/lANbvFyZwN70AMvTx7oKSsiD3LwWkV6rZzXOuyJsj4Oix2UZPN
fLr74EC27mm22B68IR5EAKfFN6TTWJDzGYQAnzn2M/dNQQbw5+vsyVBkzx6i
htAiENmEQ+GRtzHNmPfJI5bRaxNl1k3Tywx4g8FdsZeGayoams2IOCkzScEm
CgF/VDypxho5uSUyEp8NFW/ujBkiNBT7arbZEf9Mr+ybe4ompdRRfK1Njh9r
aa2DOL/8hZ1enbesHpH4W3PgJmGUGtfad9pCOVoB2fKRNdCFRPc/isKpg+uo
gVgLRQbcN4ijxd5eKohImeOYAdhH/pM8Rhybgw37lm3HO5LyNXGpcTGVjxWh
Ihjjyu/CUsW5JgDjj4JkDgdY6nrSI3lvPhW13vR59zErlXvyVG+XYqkpa36i
zbG2zWix1pognYbUWPMV3/ZWszSMxrn0gW4CB8NAZ4Ogs48j5mP4aQOd0Wf7
sluhC5lQZri6xcRRo1AczFCUexMVRQa83qxBPsjnexrAB/Q+wfC1BS9vZs9D
W9unzkOg/p6Jw5Ym0OJYD8QinjS6dNnTaUvGeMVq2NuKkRXLxLZjpDZVmugQ
UfKYM8wZg6KC74MemNgVxSM6qS44MqhW/Yjv5F7gBP+V/cSLkAGj2xLdJu1X
y7pY2gXGdDApu8MAYb3p58bdprEP1zx5ZTlIosMvFPGTUqmGX26hikicxxmq
km0nmymZTwUuO+2NtaJNE5Tf5MfBw3NHJwIrFbiRKQth65dAKj/bHzjsPJd9
RSeHyIJ3PoBsp0fV1pkh5VtIZ7Q4BKapT+qkM4sb6Zc5m85YuwtnS5h+k95u
LTUlMOBfyIuw/5CmsIISDvAUjmsY8LzhcxpLxFByGv4M9b05Ci+C4oMX//oo
5Z4zqQ09U6rmOaKa8rF3QSPgIY0Ge3giFQtyY8ljGl4yfI0ZvUCOec7FHR46
n/vKKBXcfdsGgJ3aCdrDWa+oOmWH16G40tE8zHWxycF+FBn3HbkOOhb9WUZf
86RAAtNXVMJoCvRezfaIIqHs3Tm4ruBLLfjR2ewlPZ7D7zoGNp9u6uxbvZN4
AQFYL+RSlc4ay8A4bXxcQnw+bAXZOxSVDWqbmwe8uGE0H7oe45rxmH3yCWzq
FrSdF5QRArtpch0eVym7MnC2EUmlutWzUZ1Qd7BEnz5ql4h6af6MmPq9aKO7
OrI69RrHEpXIDg5ou6JLikCJGw0qdOn6kHq1PBmg/UdCoxL/E0BmHNEQC321
HHMdNOdSln7WztebzjKDpgmEpAWXhK85JMvy7o/Kcc0jGa/JeyoO38mZieEx
Nm3WCi19GNQxBsAGAV2INQVPeN1F+1AFyOkL7Zs/H7fCIfkugWgA/zYlCBvp
j2QLjS9MygTMVeDMd3Mr/eufwpQM7xO6z4GcNsMJvvCaygfmbzZzbVsS/4gG
3QkZf/Qvbz8+nkVFkb5JPKX/JRmmatlkW17JQepnkAUXj9cOff9qeSAgTSkL
mGtuR10qZY9EYkgCNodkrD5Wjjwywr/g2gVKXZWM0meYNMuvM0KxYegjlbQY
S6uhiRjCjfrI1D15hFC3x9FGRWXxvrmicEu6tSUFGEMgp5wtD+X8ka9TadMK
3tGPpZUJKmZvM5dlBFFZuhA3LTuLQ2HVL8C4WtcpJkv7c8M9h1LHGR+SFfXQ
+zL6RHYGEbv2T282+fHxz3iALm+//L8ao0tO/McHhcMTw9lo7EMmuzamK4yM
SX7GLUF3yql1IWBzlxM929sFZC4iNfz5wHOsvkOtPoiusj6cZ+42YWhAE3sg
WNbngchR5J303N0NUqztAtQp/OggC7iCvtwISwLqephLtYjbaApKsrA9dN/u
Vy+NRJM/YJsUoZ+spDXuttGc4ps+Dm5ogWDLi90TKVOSzzUJMG4UII+xooKT
f/Qe2FfeRh5ry58mVl9BhVkrZ38MooRITLXsZWDlGH022xi61Nr6GKDkeP9I
nVxN1jgKM7J+6iK0QnJ/yYrnyy91L1u8JAhTfzkKOxxB9G5iilcGtYouWfTp
mGwl8UzyA/v/yChZ1GaEYpiIeOmGh5E7KLSlgchePsvmTK9T5P7JQaI2aHyA
phS7S8hNHOyC+TmA7FOHZiBhAPn4AJM6SY8u3RG0ka4Mr51qu2RC5KEgpGIL
Q9CuoJRVBXqj36BSt7nPlxTfC/3Wzb0J/Dfb8f00YZiOEXtZ4F4gxxLfJ8Eo
pe9+Cjst4WB8oYzblyhjDLE9yw2hjyowb+671PnMN9AqBYZ6CyVacfMa0rc7
ccGeVl9Mro4tFqCFp9ehe0fa74Q1zxQWlHCLdkExBGbgAZQ7valjs5+i+pEr
D1V+zTt9pGniNV8Ua4olqYvG4Uk20GS24CGMQO8hD0cFSiBYKWPyRTPC6dzH
pbIXfThxtyq1EykyZjLzrGDdaIBZNyDhKCwDIah2Z3in1C6kYsD2L+EsZVwr
iSRIHQUz+Lt99vOH5BADhHOfvie0D1WzFYnWFkMwzdJaSCt1oLyAx9n584g3
/jBhjExP7DuK0JMJG6ZCJqnGPSwBsIflzi6szKLMvmUG4BFz2ZsLzMUJZaQB
uROH+yv7oF7R8YH1LQsfLLTFhgqbyepZNfqcrfm9imq2NWbpyw5djQ91lVCv
ZiiqaO7cBZAheRMTeu0G33DkgTegCpvL5X5i6bJ5DIfPE0erBSEnYy6i5n0j
rZOE1/xeMrOvrBpbRtv0Bwnpk3QUkupV2+WKYXoed8nAQHlFKKnX0BREqZxA
yO+IwmmnLuMf591joXMQI/xiRFnoTOHCIHA2tyLzZBABnpYK2UNcxWMOahZS
ynj8VPwPE22IRnVlA7g6FB2sgxLx2JbETEoRUsJeluEPGZM+tHy0aeCahk/9
UbvrIVZo2kSMAmhqHUi8d70mbtI2z3/1iUNPGoIYA5d/hKb6tkbiqJs5rXow
1zvrslnXkUbHLZ8Ra7gRHgJFbKYNvGeHhsNMcwI9krbEqtsXwvAwMRprlYEG
QnvEM3XrUFvX8TF2hxYfzxuLkRYIWrFD6QB9fKLBU8IaqyQVWI8oVWtEiLVo
W3+U6JtZYoYomHusIdaCk/B7QNT2AF/6eRCttegfKPATJsEHcLjJnsW1m9G2
zLXpOp3FRc6DTY4/HCPtJHmIuJ0ppHMlN9R/ThL3PAejXgDdrzwVGBB/uyAa
FF25N0WyAA1kU/0OtMIjeoseZcYFLxorVMT+Y/09sbcqCYnAr9BWM+q/T7KX
aqAIvR9t2fYbrUOZhi6goJYuN4SITUDYF560I7QOJlcXkuJmi1i+o1v/bpg4
FOrjAdXMrixawTj/QRAjT5EsvyBeRRUnGh1xyBwwIamkECJJRvbSeOpLujvQ
6EbUD8ybJAL5582Wz+ApLmZJAQQMFVHNqrFiLfdJBj2XDJax8gpJKq5oyVhn
Gunz3NkytMC81Mw1+hqrGbCDcdabjPwibbRZiBrNefNmfAMR0PvzdzWb8TBD
DjUCbGH37cRvaFmKn0Cq/yuUmrk1Zu6MVoEUP38cBJxJeq6+JLA5/4P5JZxz
KR3tWObfZGiTHLBrsoIJpts1cdwH3v7A7J2mHePdNYpbZZs3o7MY1H79w3iV
y73kPM1tOXCAQkhW3PvACxCj+gdmwnlJGqNiUfEfvTdp3CRiwL/bSzYVvEH4
0P3xtiKaprpCq2xvR3RIeX83URC6bNeyaQEk6l9Ztf7sWd3jsgSX9DCVWBfl
7HjGnPP+FrWjOhelvHQvYtb+VRhHfCTBzneaVx902DgBsJjUAw/zoqGSEa7y
13AeIm2wEBGtuIwwC/iO2+ioPi3r52/sTjv/OJyjigZX3FYcm/yjO+pB6NDW
NPaTtGRR/ceb1PavtDqeVwn2AW16n9nJbXIy9yLnD9jToMJ6/UOA2Md7eL8H
UGQaWfsqFWgCyYfFNzQv7gorqODz9CvCUypYzmYXc2f1aJK1KkNYbvYbS1cw
l2lo85++ws6t380LBmxyOLvXNVO/npVE6+S5NmSW/LcAHSQjc4kVsUHC5bfJ
uOfOqiguRUBX6wLPmMidK+3au4yW2SIQ2FAHbfL6smJIWtJfqyXfh1FY4wEL
OgASXrTdtMPJdw7aQt/rO8JQJgPsJ/rd55KtqwIgKEyA6Tkd9sPSD0aNHtcj
PLqXhoMvjCr/FHG6ExwJ1M0x3R8NhJuXOT5Ei/LMngVhl4bph0HQ2oM1QC0w
Z2JOVv8wQEqql7beTvXa3E7IKo7WqnEE3xEwZ7rpnu2Y9GvBlU2bF2dQWJmu
7GiyDK04NZIMdswcEuVEITr1iyuveDeUOWzWfc8ltdyL0NcbBnXpTSL9CFhX
TqLNSDkbeJJFUxfUJMiBwTHdoHx1Egf0wAekYPNgOc4GrFGKrmXecn3p4kDG
za9CkSz+P3Izz1dNs/xcPcWrxTbuUskuN6aZRmi+PpJGO5LO37eKeqxq6Mvu
w5Mf7qftL0L7MzrimW/bUvikqTPpGhUjTXWZl0KrxMA//brHeAjnOItXH6EV
8+laGo2eDJCgLNNdR6YuW6FPKuBI9F9ZYl2mcMLM4ZRqoq5t5U1sDHeX7teD
fQ6AuDKEEgbDgos1h/zBClLeCCLBvSWaGDQr0KOLa1jtpQSmPRWVhYNVdt9Y
KbNTHgNUAi4Jo9qc0sQSFzDJFVOEwvcLW8Rw7nfa+Lopjh+2gmibOwyTEOok
1rs1rxVf1K/wctn5l+mxcegksuwCzTpN9Zv3igUFhOB5MK0XThH7+ZwnC4Jf
jee+SXxFEkqOaqrCb1HDiwB+e32SRAbMhPFtfunGLLOeXJ+iGerrzH5Amh2J
qncQQf/GSA3zyLaovBd0Ya8OiLnUEtWT4Rqi2LMMZVeZSjt9ot7Dj5WA+ySO
qMhyy8i873DEX1vALrFQ0dUeaPLg

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRze+kJY2cZEcQQW8y8SZB9TOi669QHGMb4Ts8gkwOqrtOAYcLZF77Ipe6QpM8PEX6pzly690XueKpj84vDbiuEeGp2T5M6E4nStC2REwVCoQU5k0eatc2AbxpPu7+ri2X1RyKePgbHS91ScaPx8sCd7FuXlNA7UO6+WwTRZvV357y8JqlBoorfJ77Gr2BC8irtzKhDCw/5JXTzV8cIewltMnHr/SOhW/xWKxgUyrHdO2jp1e50Xx2/11IMZ462fg0dqVp3n91d05m7j9TnyS8ezvr39Prq817YQq/dTjZ1CoPlpnrldLN1mupX/8E5YKmozPsSxcx7xhSAP2HBnfIC7V2a2Y+eM9ryE5yyEJElc/p9o9r05h0RwluRE13yDs3sUzeuXsYV1N+5Qv0BcZi09UQHgzkuV58Q8k7n3yP6Q1tudqV9MTOeD693iw0wsPEvY9SVIIhOc6maIj2bu8a3OESAF4Nu3CDBaby/BLEGJ0cWJpsUMakmu88ESCj8CGIrLfSX8qZPJv0MkpvRNCetxpbt/Nic8DIBOGmRKkTJ+kZlldyoG1PWm9rGWySWzgXthKp9RXjZTQhOVMBgk31OqvHGuNr9XQqArXTQAAUS6M4cRhvehNJu/iOy+ssnhGpfTVuy3gTstwu+r7hjFxFUC7tJrGgpnSr9x+mFK5eJDqJLXEok0jOJR79MBeGC9l4vkzrhOf0XH7nWxz55gen76Z3JxsLHrYRJnYM1c+MK7r2c98VsKDyGW7H+toSUP/zyFgFrp83a/s64vo5/BFD7nV"
`endif