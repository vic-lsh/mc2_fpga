// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VnsimmeEbRElLys86d+r4Gaj/MDkZO+A/JdOK9VzRfNAvWHGALFg26nJYC/A
BEyp6DAPs3ia1BMl+mlcbGVfFuNnmU2ZCXA1sgzkmeiAv35O7imaCokQ40xp
1r3ZQxo55E5sbEXeJEF98pDsjRQuDfcinewbtlpXu+LKGTfkhMZrTUcjRziy
EGve0G/VNy6l/i8zJeciFWheLFZTOzGWlqJxNe78fMU9da5dPwk8WUBpI0YB
hkXIP1KnJ7uCtJ2OieAubWYr12r6oej7rPdRmxAxUoIEOOI2M6O9Rv7FzybC
F3zQGpUGlsBBsZ5dWn7qnqhV34oKHQGYqBeZhdHaXg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
j7QhCvFZVZOxR76U23J/3OXXaU9eH3Ly1SwOpXHPfgs68NGfQP4ZfqXgZRGg
li/J9pa8rgc8FwziVtpO99JagYkpN82kHHgvxLd8JuigC8TX7H+IJsE+0A9E
dhaUqda5EgcGLmNlBmm1ha/l9szbuOqyTRVULjtmdeRF/gH7U7KUiXcN92Un
y+XGkavFBQIsp0ViBQCicEAZ65gnKnUiU8Qe2pkh3v/+V7kdIAtBEVxLA2su
QzHP2WxZAqwsfLbejUwCFEPGLJXMT+yqEH1B/juRjyaDxxFkngRmQYCD5gmo
QoOfSfFmnXzI4qFIpsdoa1ij6wbzmKO5LuZAgTCBqA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
evJ6PK7XpqnvDEMtqbSNflM/KpMFz3KCk2M0GGzAUmAbJXETrkEdqiK3xwKH
J5HhGi7FSpbkbTfl2YgoQ+CoTQb83uMcGohGmSzWlXhCdbpK7YxBqHyBR5+o
4ylAHmZrcLLoSBuVohZWSX8puLrR9jhpwTHEet/O4XiGQ6LC7MZfC/RfuaPK
6BXqxFK2B08jp5SzUMGNNBDxWvrbdIAT3KfqXASzaN3Mm+9AWV05cGbWtLMI
FedMcdrfFMCfDh1EB+G5UhKWfVVkxoMBe01x+VdphtFYBj0u9Cf8Cp6jrHfS
aPBepvwmov46UeMdEVodNCoJuwqEEorkc6Kz+uiqFg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JW4n4YttD/TqNmpAJ3zTyzSBk0NvL9k07L4g6mo4AaO9u8INxzHSsylkFMk4
PkHQYufSEyRQl/sFWvsVBlXACZwn4KRvaOaGrOtnLpd0UKdnAnH9hFQ/pZmX
cT96RBxHyP6eo1MvQxnIUsckQRnEAxxlB61mix8ovcXMOBm+G/AvcemZbTrE
gxsL2nIBo3KtsoYx6ZoHClIsDlsIqLJsu5L1LbmGk3BpxqI7dg11/I5GFr29
9aDDWEaoeKBqUDaJyVtstAfHPJBWu2vZK4flY88No5hra4Kh4xTdHkF41cRU
FXKeCL7L+qlWkALYxBPcmabqSASssi9jO+v2RSPPWA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KIiFnKgs9oYVIQnwVkEVZMq7696DfoXZ+oViNS48NjCxrwJHRmDy31CyWJcc
tietzhcb+YrCQUrX/Y+Nzs7JNLAsqfHvndt04rlLBZmTYZbCbkirpJy1Lxq+
XF2ToZjvyh37E0AgB8SwFgMAP81F/vqUbwDqO45hSBpzzUh5fUQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
af92d+jK9bs2695SEjF4lmX+Y5HEcRMGmyHn2F5xKtaBCyHZCes3g763d8GD
Go2yoopsmaSMEluBRsKO5Xq3nfrrOEdlGKkyAQCDXLA0ePcomS8MluXNF82z
SG3XW7JsDoogTZPbh96B/WdGdh5FYota+ZxQxMlHZm3CLijLQf2GReqdZmtp
8BDkMIOwyYZCsaXFhhC4jtOi5FqCgydRjGvxiV0W+ZQsP+MPJ5RpxZOtQhj+
Fo4IZ55BJ7nnUXcySZI4VrGhumpb42PMhksh8VvNFdJZCzvHbba33fs4MLQf
H9AL9p7X3Ijq1GONLnUJ/h7nISTQMobgxtM/SB2S3K/UhLdRUiF/m3Z88ZAB
u7PsDX/iTl0A4UQ6kI20BJ/x/7SOBcta96BPEokFwj2Dkc922tHDmBf/YIzH
GMgxAkWIDweNnhgVmHGa1CmZV1zN5SUI3rCmr0R6eQXgFPRrKZdoe1mf8yWp
DBoHo6CZKnjUITaiTwr/zijZYKnuCM5m


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MY0YOFBcmcliTkOF4oBBQh9N7MefJnj2/JfMzdtELSdiDPPVz9nRpfKHHAOx
ke2IsJL9iOrL90pzmVrxKcQYAEQgaL2TcL5NPFhx4znnDXf4v+PXlFI2tcAh
xTbpfNj0QKXrdHP1ITHap7qDg/c9QDJOTJhXdD/TvMcs4/rd6dU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gzud+Fkbq6erFODWCKK1CYp1UdlFVUYTk6ONUi6+62iiGoDEMXmQk3lje4yV
A0dhMCJZPAi3Bgr83UMi2APth6tGgtF01jAPTTlCIM6xF4g5Iyuwyikje2hG
4VPErRnHXfJSTJWZuxeiHFD93iOarOTb4xwoovcBaK5mGh7MW30=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12272)
`pragma protect data_block
AzMc2aoDHRhI8ElVydn1f46FN7lnp4gmQ8fusvatmdayAtKIjFPW1MtDGHTc
nBs3veAqYjxMO1hFExa5xmvSxKQg8VN31AVkInwgxU3tDfbZauYSqXTOi3NZ
mnwS0+l3PFb/c0oSM5f0q56GH1s2zU1OG44mKyAgm+01JorPzX9VmYu0oYPh
h6LXNyZUVjng0U8stDnQJdXDAbUzd0hb3w3AoqLfJVBlLz1YXeV+tY6K/OHJ
qf4q+RITT1mSE6NBUUKWT8xg0SH9RUtl2QSTxu5bFrGs6sXmg48lbFfTALCy
8rIYnJW/T0BpWxnZYyHmFphg9Us/UStsd+ryRAACSzENbK30EyAYdCBdV7cM
YXnmVIuXOR7sMoZnwNTXVmP+o1Nz04hBTPXejds/ZpPJ9L7O0JN/ANnRrZ7y
Jd5uu7TxXlyRZg8Vhkjn3F1uc7ylbXg9b6kK813aNb/unjpBiiwXDAbLmtct
+In/esAyzkovTkn3gNQ34tGQpyHlvyvsSwwDKKf3ueodrF+ccW3iLoQKe930
BWrQqg2C8G1we8v6BlwoZ/BmPZBuoUBkK+pB14thracW04pZ5tN3JEhrAJRQ
63rhnRpicQIJxlG/WXFEdw9WTVzugba8xFYzOJNTzL943S9Ljla2HBnPEFvL
CLm2OgrTtJVYs+D9WEVlBre+/hiKqBvDCFYbS29hOXFJ7KwloDijyq1d4Uin
EaCY7HE+qo0P5boc0UX3h58nIrhrWmtNJyobl7Yb/3z6Zlz7mlYkdu6I3hkU
gGWwO8FxbxrRJSANLQwVRpglKHdXxVDF7+vialLhiSz7ctnXRgrbLKM9mIPw
G7I/AKfthWIUcVIw9dZGWXUiJecNjMGTDsdKgFTDDGGZMsA8lBVgRlrSkL3z
yjr7EbAelSPlH4uQ4UGjMhOfpu0Rt1UGWrAdJ1KVWNhR86RCeH6j+AksFjfW
di32W2rFqKEasK42JeUs3+KngSQK8T0HVLY1NQ+RmBjah23H2/pQDequntIU
DzTEZVqUkBHJfWaSGuhxGnVk6fFrCFy5Mx5cwhtCsFzupCoPNF04lromjUeG
emdqB/k4xL7/zExszAxg5ma9zuUnXVGS8IJexuvhKGGR1nocTB+YDlX9misk
ME9Ax6mYVlTllP9W7h7Kp52BtUmJ+JLh/0lE8HYeK4Wh9ZqzUrn/3/DcbK3k
hF3yqCK2Au93syQtmidKWYDzV/iMEc0f1HHzhCHcgpiyZ48PC37Qf4/PiV5l
TLvTWDo91nzGpbsFrc/6YTCVPgx/q4tDMQRUvr0C6hDyEfb5XTV6CNzljqFm
83P+64+g6GXAVJFmxq61lvEgqJPxcR3hEJA/PtwcL/P1MjYbMNx/kIMHsFAg
9uFO/R0m9ylv9a3ywBEqEMPJdsoMpIr4b45ZvuRRVYVLDkQFt+do0v940+UC
90oqDf9hKaAcAehLF6KBqx88bnTpzmEQ98AdvXHWZDDWvmqTV5Qs2eS+D1E6
0FllAwvXVvL3rinRwzhmOKYPStzZ8i3UheX9QDE4K6zXdA8KAxyNeXCCM1Wo
BY09jPIlvdRtBOYFomRhkF+NFMlmZWpHCwuAL1Uwo69Xwm9+aeXl3FVl0YZ9
y/cHcU+oi/zviLhMz2Jp5zn6cS7S3KgaS/F9QVSNeSUJbui5mQnlBBNrIdq3
I97PonpnriI0EfJZJN4le3kTo9ucSRzwsELA9DLS76rWY/3z9+YPqrnDt+TT
FlrurgB834Kz90KApOZMIspLTuyh8ep6RvCTfUkt82Rf0V15Fsw2QnKlwgOX
5co8zDQZSmly0WBoEHtsDrjiaplIATavJ8/uXCFuQ/05kQTWHn1WOwNCE/ZU
f/2yak/xdMXzMupiPBAohyK0c2e3n5VJD2N0r1Cmd93YV0BvEAV2KDDWEdrc
k1QePcjqq2zCcWUia/ww4qLUs0UuRtfO10BDVcifhBI3d3L9cSGuY9YRYRKL
FGZrc5QVwNGuR12Tl4mEmawQ8x4TMcuuoByslMdqRzwye1kaxcG3XQzUiz+D
nhZJ4HrYnF4GbJi7m8iMeyPrQQqF4vy64pjqINxvrASuaFOTMIO5FhnDtHfy
XQcg4e5C/ydQ5OGYkPcB8F4lfDvo7f9UZO294nd7YZpDvlF+IGRogtnvlDWr
La0bGobSjwqxtFBsoABemlP92lvRoHUGqygAR98vEhufqqCIfQH5tASrRXKW
NCZhZaqrSMRREXvylMS9mYKNKQ4Na4sKB8M6N67vVH1MNEo4mrZdmuuN5BEp
F0P65xAYVP8WS06d/Fid37jAy3Git2l2xfrGFv+4ddK61zcmQDBDm2+GxNdR
0Ep3Rw5fQfBmE5INc83FAJ1X6DfYpO/3S8/a/J9wuL0mGqdm5w8pgPq9t9Ky
OaUMvd0uPavwStFLFe8ezLZMJUwP4nqSYqzpEu+Bucwumpr9e7AnYrhZN6aI
xfCQVk7KFUB7kJqYMYwJpzI9cSPYHFw6utS33jMapJ06KX4vgwpOhKJ0mV5t
EI3FdHck1PXMVkEFKEtikfp6ImL1DpxYggOl8T5ZVrvxFxYScX20sJujZmTX
JqByLuFkMpzxafWXl4TR+T59s755fF6vhCk8ftTDdBG9FKqBfsoepJABEY4/
lbNbd1Hcz4e7hCFAOpuDqIDmsJpsFkPbKBblO57rB5qtBLIZvtzrbZysNOX/
1aKY1H0Xpa6w0Kt3Ur4PWr6oG6zMpshA1IlDD59N3Fmjjp2EG2TK61gMhBph
rasu4JQVA3pIbg9JFSN+J32Cw9Y4Bl5L8aJIlYpnl6kvuXRgUUMWs+YsWAaF
WcYgTQDpR5TsFAQbqAWyJLVr1tK4YvwF665yvmJZoDU+/zPLEeq4PO/vMiLD
LPzXgCYrMvnFtY0zk4Yok6ltIDXOWy/7J9TbKEJA3Q9T21vJN0s1P8bxDn4f
c73Bnbv2kk73Roar6p7wUAk6IfHqjNmYjsx9noXgJYKZdTN91vHm6j2B0XOc
bD+IjY1ojMcpZx+/B/5BSOvc4WWhKL2NU/Pk4Jb19NMmjpFuittL9HakqsO2
l4bB+wHYhawWgqsSmvVqytWHiLnS4LY6zTePZI2Rxhihz9A+pOtwWTtwIjCw
/RnTVP141wXUrLJgFVpttiCyqM2mA33uugkh2laPyvjwX/s/msfABzuGbv3w
Ps7tbIJB3voCyIovxY+vY+ic88OptHlTlsrL04RGS/G6hh4DW7iPw6nSev+h
uN7zNO5pgHMbH+jz+FNpBYp9BzdAgT6cjHbpNPNV9hb0o1+n9e2fw6MUPfjm
MpkZCKUe4aJJR128YkysAd7wPUuJHTo9eiSr7b4TkbDNQUyoU678PXW9wbbc
B4AXoGwh8aLGwxLvFBhtpIRZgJeekjmPHxU+Duvc46RuLOZZiyk12u+E6EBr
NgeUtigN4wkN0/cuhITZuujDOe4S0SfSwKqudbr71T7NTsGmrtihhlCYj65K
kV7gopimbc+gv0+NY/vxMxgqIfc+i+ZHCw8E3TihfiuCA5h9Wa0vFlTHvvgz
oiXdcKym8Fcdym/7sWtZv8CnFqFLnn7e6sdlIdwxn0jfwFu3RXRcSax+kzxU
c9Zzb6+rk7ZxCPrXQTiPGO6Qg4urEz3ElBmx2CtijWo1C8i7lZOPBwEbtQI7
ZyqLBG1WAal+RUX1ZnTynSoK3hqvAlXuxmXBW4DgDyRWIs0+3Sfv/yEc45Zm
/XRuPSI1Seo7ma3m3G39U110kXGE4NTPsZzoALNdbbytyjocAbPw+DZu25Ov
WIVsE4a6FX/hWip6EtwH8BrfczwUhnzbYk7vXrE6Z5xphARSsl0Rvv6P3+qN
AiMA67bwPtPhU6N5IMeGMWExoJBh770vyie8ItXgiIulRGtkhk8JENA8uFdW
jGyY/wI9hiVtspAPgzJ/7ZgVAxIfalUMrum9YcY/ieUqhoiXbDsZUDYWkHb+
+Jz8zGJ6M/b/zaPvsEc9YUrEtUkAKzcFjwVYVBA58Xaaa8bkEU1aN8lLvJMG
h57x1S/wZDBd0hjnMzDfuu06Q82PzKX5v+1rB7XYOfOP1rX1CyD0R3wNNGbZ
sZUcx9LQGCID+bNwxpqt1oYbMvIEz/u2fjt3JBchf/pfMU+TslZMV9dmvHMO
++z82Lts/23d83OxGagY0c/VAOCFI61qRl+WQkZ2xUdzYiGigqr3pXeka97H
0iNlXhTqq7d5japPNc1uy2Uj6n93YyKhf5GF2h+nf1i8ELZ+9J9r78npZ+R7
XLxCbzs8SHEtdyehdjgbT3k9ZyBtTU4ctrmbuBqs7jIVOBbcVi1Z03kCfgFT
hOVqRHC5CfzQIPq08iRVjwqWAgUJOODMxEJAI3tB2acgiEG7kdyC4RIg7qPW
wrmy1+OtmC5IOYhH5vOV/JKpbdKV2hOXTTCTd1xivZ4QUZtQ/zPh/a4aWXYA
ImzmhOwMrf1HRPFT6WskHxj0je+yWLbigMEX1GxkgVg1HuOiZvAKiDOxM5Ya
5102D2nvEqZkgJ7mChl65eTqRqifua9j1kYVbxj6+GMnr6RBWtg/bbZEYLCY
T2vQI9MnW5+6c2Jn251UW0jYhcU9lNe2Bu5ElrPVTwZPhp1XO4enZnxaonmN
4MzPYOWudMGEAuEAVEyQezDRbJfl6mQNuPijuUnZ+ZBhp0+yPu3nyXnNy34t
OGQgItm5wsC92lLNB9O8hCD7PyWhsnW/UQ0uQX5T8bIwRxJKmm5RfBIRBAwZ
Au97Iw2au8dv1QnyoM+gZ31SpN3agFyoHAXMB4dvBQX/BWRMzNGvPpJ8C4Bl
cyrT5o2Wboc7iAhlXV9J87WSJn0+7LnjgNU/erFMoLGc+ukL7Of7cTl+rCQE
yNkSTQmyWlyb1S/6MIRss9CkVcF6AdA5N6NB2FM/sBXQVd1aOOOffhdj4z58
C99nTDHU8BOlsFbKzgbuxo9vE3T+uTpnsURZGNfnYF2YYYxJSVPgvKhlNC09
kxmL4cpWhHswGaxcA5fvw5sJGRiU4Tlk4rLgiTdgvzjFGVOSuuIsW3KztCKa
FZV69F7c+9HX+UFMxDxvfFFZB5j0MfIk6ERwpC+hi32ym8R00S/DOJHmloJa
bgzu8F6zNAGCRM9c0At8gfjfEwSXKFra4aIRyw0ihVZmDLYysD0oQl3z9C4B
8KMRFLBje5pV3pHtLDnX7E5Lu1odiHNQltWe6lseq9RdToDjA1sxVlaz+P3i
i3VzrpSKNrURTY/34Rt7/xtuoOreX/pKJcxutXVhhgEAXpZaAAAAsfDVzWFf
0TzfLIOMLeGTFrrtfC9neBeOQv+W1jpUfnF9hUigHADJqpgDhGmJTqTdjRtO
DeKrDEZhQm2rgG7wtJIWdFj6vFsnxZRW++UAt+vuwHRP+3fflFUScUs5SVhp
tdtrZxjViK0IUmLK+mNJ47UY7sBv3pzXPSuQzBAHf7BwUGK15jnbd9s19uoV
8YBcwwoQz8rCHZGXmNUqxrdQOmSTXOX/w+fgro9R7B0deec8FhHWY6RM1JXf
1sLyb718DUYrBgcS7qIfOLQ/1ODbt79Jnv30GcJGudSQGi1o+Y4LEBFPPdY2
xpppLtHo4oacJVHBfFherstgOWGGarw1ivXBccUtwcdWVMXgamzWQMiEn3D7
LD32G4pXy1dlWVSxVgYmVdzSZybHALfSUgtRps7wh02p9GMkExAnks3fSuIC
eDswYQGgnqFom/v1p4QPEqpX4WT8u/xSVQbFrY2jLai8kRDcFpTT6uv1y6V+
mG5BIJrVbyY0G65TzaskdMGTFxn8XClF71i81eKGU5uGVTCeqGdpNjnR6LlF
oEajWm0Ho6pznuqJu/Syu2Q+ctd4+CVTKrHiIldgUhjAm4ZXJyoaN/Z5XsYB
QqPBhpQMsyjDO3mNUZtnedTk3oCGTGU+XP1hLXGDBiY9Gro/n80rljwZuT2m
3psDZUi3QE15zHzDRFLFJX2OwyVLrE3U41LMrxpNVvJfwjQ6BrwhkF2kZtlo
aSJY+oJAi6HGZSDwsmtt9p5ygC2x0pmV8UoatGzFSKzZl5hGBzdmZ9XRDIkw
3hE+T8+82MVn1x5hoZnsPomeNz7UauujKb5WSfud4YtIWKNFIp1a3LNpAUJz
+iYN2T01juNma4bXG+Q2O1DmuBlwUrgegak9BrAC8G37YuCSPHUYAC1MexvC
C2dces5O8Ae7cAVasKuc+n3HFRFoe5YqqM95MU13aMzeO64GBkknlUevCGP2
KSwthGwf3vDhmzEgS24KmcuBhcIPqwnOGeuyBvISZKHQqsW5tg0a90wkeiPw
3DNwBtSTmk2CFdc1+mu1hH2RZXuUMwfXmviWzbA8ig1q2BiuCO8VMy5LaO8z
gz5yn0PX4nYQ9Cq2tCQZvPD5MUyn4klYrsaEJkSbcwZErQgIyx5lc+wf+lSl
fUHnj6XTsX8ZHc9rdOvmGgOnisti22xl1vzk0rOrerjOiAJ2KTFteS2QzttG
Umj0xjjweCGaHaWAExm/RGc/3P3G+b0tutdkscdvhcJwBDh57ibUfhc6PU+B
vnbeLsBKH2hx5HMI1Psyp6UclQfCnPGYsSa8NJP8FpshhPUq1cdTNofz3007
rw34XAQ24nyzvfcFizl/9r4xVLkBoFU3mdqzxgFeyYnrh5I01ZNaDdwMb5IU
MacD744uvJ9/R7X+S+Mz9KsS9bhEtf+scjII1aQyyg3cNZZ/MnVeRE2MFk7f
hpmM0HsCJ2qTx0/V2Js1Fclt/SW5rwhHQzztp6TGlj5WS9Mi5PLaehE4niQH
TUXp0G4NdiM6uiyz4/WxHGGpR0N4NAVWZsaWL5wbMu02Ke/4I2m7hkk9iFdH
ryWdyneaX76SDJ4CLuF4p4BgISN6RHGYb4PcsP8WKyiKeRcWw8pSiwIiXtkb
YW4Ct0dr4gFd2e+t5NRXUbtljLjOIsmogY+bf63tv5c/fg41rEUR4muCqmBy
MPHuYxeLhz+7J+hVMalXz7ySHEGvZLQoqe5Mg3XS3AaYYCkVzcswglntotiQ
fsmhdVJurm+2vmwln7JAP+QmuExCy61/4EOCuY+3RygnXOg7En6IJrtRh4Ym
S3h6I3XimDg3LS1t58A2PNxRUm/tYRxIzug0pomM0F17ru2VE1mJnm5Se3Xe
CK15STsN56SY+hhy+Xvx1m04XVKGeinSuV5mT1g+AUXf3GN60eniSd2gm8Yc
/KttdLdhOD6ELxKMeJeqjs0u84/JbIslIKoJhOpKoCqiNak5z9bHQx39b+Vz
fAIJab3O+KZFseCvhqdgcDIkvF6q2DOt8vya2mYG6khIaobtWi7sqULOA8pI
Xl5u97DTlq+3OELDP5eTnxjNyiby2H9gXr3Q8Cr6odWZhzmgp5zLHBThFYBT
MMp9HgqtwRwDjK7MLD86Fk4QX98nQNfiPKYQkzQ5fLbxm9a5QTWJYei8B1dv
jUCd3G7tUVlNtrXgjickSEBQqUorzX5tUItC1hoNX2BdIRpXm2GnhZTulV5a
/9q7cHwtdIOsye50f9lz4Y5NfhqTSu5tL6Lweg/SQxzyVHIONToSzczvfTKy
Hl10MEQQ2UmNbPSyElG84GUjTkGUeU1JI+c9506cdXRGFC5otstgxwFGeioY
V9/ie4xuPviQinD4MtI7wfSehH21LByDvc2HrAsgNbp898tN16/gua8NrLRD
N0chvSWXcHMUWXAZAXWIWh48IxlINVgsL2+UiSFqOVGkinuAZOZXlRV0Olwn
KE7ht9fQhFbiiIfCawuDNW5bljWXvH1ytdOKBkVUecaC/Nv8rNC6jLuQB/Hc
IrWSGZA+f+6HKH0Rnnrpw1s1bxyuwZYqFWwpSj5/FowYCr34keIm2xqRhoJv
+59PqFdOlHo6uareDi/88hpAF8NWm/ayBjaT4K0qyWo+ILNlc71fYYsJb4K0
ySVtxVhUVlOgJg9P0yZxc/2+kAP0mzxKyaJLQ7rDt7qWjLCDjJB0hcpJvno3
tXGAABdZrBcCJ3oC2eJkDVAC2oz/vnZLwl9/IlowQ+c6dkvOphCuBB1tXnSf
3DOyBd8T6/Kf0K9BLRnpa/8k1mAHjLFZJH1o+XDerAZEwzCrIBhHEwBexVN4
njyBZrMyR3KvRvkJ6z6bXG0XWiRtkG/Xb6pRrA1pVOQp2lcYDkb1gecIxuFw
clV4PKsrlAVr6B3J0KKH+pVF1/t5thaw8Eq2znihr7G/xtwSelsHNA2xQtr8
pWnQGbfcompbV09DlI9ryjBCN5BU3EidDXHyS942zzAolhmW0w96lgMazAHP
unFNpNgrohisndMthPcsciQ3KaiYkOhAkCH52gW7S9NX0BnXO45G010161Hp
YqYrhZSjllaVinIryzJqCtvKzqlYiN+65W3+WsfsAnRkrOoBIJFgIAM3y+lW
fDbULdUX10u0U2pnvxieIois6btVrnDbuqX8b8ggyHQNFLuGm3bGY/d0AAOQ
u/Sp6zz3OoEzGjk3LJhlb0zm3ueSzrcRhgbZcnUirR6UfFP+vKRyFBk4rVUn
ogVMvGhnHptncLZHiBeVNO/VrWf/yBmdN8gMuurQHR8pBAT8Ru/efKihq8O3
aIBmj/RyAYOmXjSplS+KbtI8WAcuBInhavCWp4y1Dwf1eg0e6z0JtYPwOMoM
r8OuGdtSb7/EuDbNdtR8tNqaaE0eyQCmujFo4NVQNrCmXEjsbHxxi+8E3Cw1
o+mm8wZMe4aty7vJVdWS060pZK+U04qB8E5cZ3zCYf6eExJKyVqXE7z2BVnt
Is090YvXfs9f90RxgnyI0uPVaLqOui/Jjz1XIWkZUsEhcU9fazTndzfZu222
pxt5G6xVX+fnOwfTWw/phEsGdwUfKYMqpaY4PT6H7pxCX/mcb5l/NBtTvE8k
UxQqeE1ZKx/QDBxy3J4MgGMjpRuJc7fZvq+bFkFPNHs4X1BFSRow5c7cdSGm
N5aZxBvPeNj2y83GOJ/zmASzHEy2J8brMiSWLNhHx7OF9wHTRFwv+51op4T6
4PGMlA69W7qRZDO3SJYGEqZayH3KGWOQ84BSV4WmlrMenLFs2dGeCMt/Tj+3
XGV+MjOWrZO8FnogI71EGhzel6guXL2BFSTY8nEAjTvEKRlzzUzYyO35u/DG
5rlvQhlWQWMgFs34hwTy+6kwgoaUx1SxjvYwatSV3AgvKDqcnlSEdDEwX8Jp
kXu0BSgi4475qCSSyd3eha1HrNKtTg4baY43RvsJRIhMZZK6LzLNmHRgDFOW
mRLqzkrsVMsUnaJcEgYZvs+YsYvBudIQU2L7bMficsdlLtJ5IuKyl5Msb/Lg
zeCxSNPQdEzyPfWM6hXFIiITIqoTglpRK9EBD1UTa+arnwNDkkdIIUG9LbjG
4nbtBFKf1/ynaa6JWMjB9IGGCX1ZubZQyQQMmZS7UjytKzV4uWfz+qy7rKf5
khyQGa9jimsFLGtIq+orCQ4SYQUD2cka/VFzwCnXoyNdEvx4p1/sW+5N9AMV
2TI8Ef0opiX1JTKQKjjrdVlbkkOqwQa3/uOGyHGH4+WWlJrkg1tmIZ10UnJ3
08JdJh5ytQJVrYaNYbpmg3aYxL5OpEGXvqOW4in77lwdI2ZNlaHGsZrUVF8c
PeidtTkQEle3uoWUHnT4JFW6QBAiLPkvVRunJ6TvblEOnd9Q+7CTwXsX/KGe
WSQuqXZr98NMizo3tyK/4oKPh8tM6P04SbHYDgsQ7vxed/qH3Vh22tXxOMLM
xauvt8FNdFZGv7Z85IkMflj13mdqOo2LMeS5qwlwDHD5xIikB3TxK7YsfuM0
orsJlELBnuCTOSO2pVoOPEMBYQ/hxx8EKHvW3wm89OvTB3zCnarfea0w7fYc
m8Py5tud8p225bluuTPTjSBmxnJR23TBGVBvIFmdqNpd4Zcy7favH3p2GBz4
l0226sic2Hd3tD88F2Q+tnaog/AiRoeq6AdMFxAihNfunZFUTrF7/WFmknZA
69YKo5c54myBzDQytEzpOxE5MvopOrdPxsWHM3rdbtGi9sEuIlOLN1Ly4kMi
RSpmc+C3ko5dhGFEuT2CK2ZkovCuNQ4bih0fQMuWQQpcRJZ44FmL1X9qjatB
ONS4pap6sISmYbK6CLpS75jeawTbifrXT/n6riDXrITKiC66PioEjnAV9Dg6
h5EogfkyuxL3CkNtz+skt61melnL8NQTigI81mOoXR3GhB7UWbelOAhUMOPV
NQkDsaaE32qx8/URHkrwpkTRS4ndwaQbIyxcRAITSnnTjsmOOHnZM9UyrmOE
jYgrGWj/gP+V6dPPVRLeLl61h5c2qjWVKU0xycYVHxMj3Jl0o3ClhmBBEY2v
iLaiboHD2Y8WWmE4/gulK3VTN8S+w+gKeX7nrv+iGeGqaA13lORjBcQqx4lh
4pnyJM2VZr3cVJSSwpNs/aw7Vo/ZA4XWCzrRGYVzTBuPbEC+r42suO54sfId
bVR/91dps2i5Ug7Cwgezu32o/ImZtf5kyS+dhW1TjjxAYrUzvuUYRKcV+WL0
2IT3QaTMj68Tte2DiEg+IyytIwF6QFRaqU5DKeipx6y4O8RZx3LJ5NX+i+6Y
dlBIvTx+dQrmdZAs1hEVMhDH3DEUDgsZy2tImeCq2uwA497DvcymeH8ye+Ur
Q+i5pIKkbPYDCclxhwU1OCRCKFu05RZogl9D5PesgpQMJaE85pD7aONVAaUd
3MOeGqN7TlSsWc0KBj6L4LBraA+LvgyjMy+YJjex2HEcZaysW7cI4HJon3lc
eU0koGMDiIVnC6zQg24tZ/4RxIVEVkGw3DEgK0eQiqZpzVpK8xELItQpQ1mg
8mrw0oilKddRSTQ4/kXZSDlg3dOUM5tMriFH3H5IIWkZGHXy749T9D+XU7DD
R0xkYLszHSOCE3TYKnHiAVgYml27QubV0YrjdmJqqDoLBrYmuoWaJUp2aWga
I3EMmq/Xv+gdHfVw8RSFufLGnOVknCpcZtogjFFh0nwyIVEAP3i6M08JB2WA
nl3hkT4/0geUOE/0wkwu6TfR9O8j1KcTuvnIJlty2so0Oli1QTX+AlXNJEAJ
apOUHNp8WNUgFXHQZkFFQT9zPgun20RD3IKIeu9Xlnhuwc2E8ywdOZbs+rSV
ZvDfPIquJ5LYiUxnqjZWcoGI1ySIW+o1HJgrm29ea2X646lxJ1jHeniLgaY0
a+X9UqFvszO19Xcp2CywQrmyIFtljTenm8YlJlVzhynAfQtRkXRO1MHdKHJv
VinisiYtu9q+iGuIspopQa7cuZEJszcG4GzJ+nalr6D/pI8dwUG2olYdBesY
oQM9A0OEQ14awU0c7t69RgZ/T+omxjsWgz0A9O+BUdijRRbKgwA1RctjL+JO
tArVo+yhbEIVLgGIifKWkqp++bX9rEWi3mY2ieQ+4YTPs0FIdC/Dljx14Yog
smxOPv0Kk3N4LVNZZeC/cDxAM97OzRc3CcltK7irWjO3w5tD8veDw3rSL6+e
kAisVdC5rfR379mXrpphalfw9Kt4ZvXHY/lIrbcpCXGCRdC+HQM2i26n+dqf
bIyr+2GNgeFGlxni437dqfyhcwulTmYivG7PIoquS2WYfY7f67caUtaTERQF
eZJukJzBJbCC/GvQ2LgOVfqKfvbjbEMqk6Wz8ie9tDSuWPVXCYtoJ2DlCKiG
CcQhy/Shye028fwdon5WeDV3WWOpnQzNG7y0fOQ93FhOKwpf0W+WVn1GpuAz
9NZpZdwI+i/nVtiBPqHK2MJrnczl/syjFw3zrS8n5L56UM8ddM2OfPyXt50x
eYWbPGgkFBHI4q2blWFrpzt3FgTPQCd8Y7GpoF0JFN81iaxM38WTDKLfPhSE
ItS0Y1UwfgjblwiKKp0hc1l5tHMkea8ZjXoiWMXu6QHQhxneb911qIA3enze
tnarHHYlZMhjuhyMYnIUBsCgbQmTrb/lFcGkKC8jHLs7UFrpkePfGJlzhmm8
NO5D9CRYN5PW+/blVnHUYua0RNMKKjGI4etfjRsjmFg0lQsMDQQ30S5fvWpI
WlQuueJHtF4036VGyUpv/Uc9nLmcMzpQiyCEyOk6ZZ+IxBPw13cy+KIgec4k
ssBI5ATOZ95IX7KX0QAZxdxLnxPyi7xKchTEAEmtF7mUcZYYfGseG3sMOgt8
KJerXJWkf1c82yT2+8539nPgIlKdzL/PfNn2O8Pu0xXet6pe0rOeiq/Gg3Kf
oDPjFMRUoYO+vEgY1Rg4iLDZ7buQX2wYYrBrOvbjBxTHL7/1gs+ULqektX9f
FwWfSEzjORfw7K8ZnDmMkUES8P2N/KmNWK2xWg3gHtwlm2qz1HskVlz3xdZG
Z3jG6QeC6wdCoB6+fymaJpty+4/Gp/GgAotGfLPcgg65E8m52emgtnXcBKtp
Pv1mn1WEL9qKYO+SBbaQyeNJtHtTY1QCmydd8oCxGyUsdouU9TCY/4mUWE18
7N35npu/Lczy8dA5LCQv+Mrun4Y0B0wuiFGKCm1/YMagzx4mQrOfXYF+ojOA
lmyj9PtSBwBKZHLPCIxK3gdmUpJhTBrTQLXt5osHzWC61VUDiT+jHHu/DUNt
9+pzonQgwxezAlgfEoE72qgLpVKB9UyapfcR4Z+dgqrv2Pqg1vPJpzMgINX3
aW6hoOv5yz7MmMFJZeN87x7RGgxqNs0HY6GTbCSqAEMSas+t1huAYbb6dNMe
xYEecvMosJb+3TnVi29DXvOWRAHktOpVQ84T3Ckh2OJv/wKxjvUkbYhfzL2E
qcIwXp8W+pHW+yZ0raXx/BkYGCtiJI6OaR2zYkLGTfACkRkuFehnn0yaGGXs
Y9PiVmTVcht2KDRKS8xzfkT1Z/JltTutRU6mdiJPHfIDXPJzX4eDgOTSKQn7
LfPT/57GO7si6OwoclxpeWR8Y8kZhjq4sDaFKSyMPEhcc71kd6uhigDgXCLC
JCdGswEAYtgvVIGBn3ZEFNPcShlg7lBYP3F7MHQ/NvwL0Rqb/L6/RQceGOQK
CuVD6aIsVb1rCIpj2DaxTRYmrVIrLfaw9RQTmNNZrSXnc6qYOjDjA+3ZtI/V
LK2RiD9a+s3UMqFsB4q0ICLpYItBbcEJepJxTKHIc8M83QzGt0mZxAQrSh1Y
A+1RKsFyaaT5jhvx6Fh5s2TaLyNrnOsLRpDeh8Ldrk1b7LCNRNTo33M1k4JH
L1y9MVNqeENfPn0zanuzQ8sneLaoF3k7K6z0B87Q4mYYrEeWJAEqEmpb61ja
xRi90Q+/P0SLljzqYzscIhbxnX/FWLwdtgxn6Ro4XqRRUl/6V9206ZBlicYu
gs6r7OsIBSbrBOnGJkW79bzLpKM5agd5QkkJZ24ilHge2pFoZI+4d1bE3uZ9
1Sk1xAq9XE8yUbUqKEBAESeQ962WLRB7hqpi8dShGPeft4t2sooHuXWT/3i1
3kXOL0JdkT/y2/UYnW3GfSQIrCJOPh6DshnECKPwffH9FYauv2qmbVD/2LpR
pddTw7qneaO1TyjNkMoP8UKn76XvFifyqPunIjz7U+sAYZin070b3LGDiTxU
F5vbJj8892d5AkNpfmTSc4DBXDEAyxBh4xBNNfoGprEZWbY4RTBdleNxJFsd
6yDdbpc+sYrx0OhdRWk+Y8cEDx92OnXt0Z9tCfIasFRnT4Q6W2WXZbk0iyt5
JePg8zNmpGOfKs8T6kkibH/zw9XRgJWuw3FIsoI/l3sDW9eWXkB00M4O5Bb3
USitZ61OzhzDi5F57FkQUPQussblQDwKfCvApfprsnxBHscM1Sv0GgtSbc1E
GGyjUiX9uHGHXidRNoULF4WeboAol7lSfsTcCzGQI20HH7aWG8lacUuxtOu0
1owYTv0ib/ptQ2CFGDmMihPz4y2wp7FajIwFO5Gm2QfALx84C1voKIiHurT2
b0KxmR9uWth9xEhmns2m4N0FTNInDXbuAyPVFZVrYJVXW4e/vTxF8l+D9wSa
NjPK4icavB+Jykf9d9coDhM7/YTrmqaMQGLjunYWjnYo8m24wYyFAOCtbvI7
waDy6K1Ny32eDZNM9MyD6ff97hlfC1QWMgjgiPHsuWnWum34Gy7CSlZbOYHQ
p6mdPvti3sRz9JgWnNzC/bM+HYiOvj90AZTFYvMNp278oIxOdPSPfCV+79HP
IAqZbwIQcZRouNfitUaViVVjeF08wi2hYrewDi0gNvvdiMFSNDLA9Q/IeB2n
41f/TrbwUnMnbwqiE5OaDjLornzLE2CYVko3Kpw/TEB77muTcrdKRMD5vryT
60kCqLvX36IcEXfmIpNlhWRoBQny3mKG03e033sal0bt2+tixwq5jG/PE2u1
J1Eto5BSYbzm0fJGhzzp89qRnDhj8mJoVjKKTPDjk2lNErw0ajptv0rSZVPS
hJn8YlRPmrvfjcX7udLCCGjd5c71sTUTV5JGYqGcOaSnwMqDcpfUJ7akJxWv
IO7fO+PgGXLPiUHAQra0VHRQXEbiyS7nVy8GizuGtgt/WrX52vyZ4ciCKssD
DeJo5qvQ2gLhQ5biFzshO0oIfcCv9EpA+Gzfq+CekNFItedNSlQVxXXPHuRI
9zrRkSxP8RL5KLkvTejN5JU7VbVJQjBjK6DmSOllxwL/XcZq/rdAPYahWXDh
+jffPIgA9GR5Sy04QaOtfPbuBkTAqJPoQqfEcVO5MbrPQSoP13hMg76AwdXT
24xM9aeZGwgR/U1VqVZ96OcRNObHl69NKZfZJLSV7m0+JFugQ9r4QrAeSJt2
ZVUwZ0gxUhOfT0jzU9GI645iiA/FEv1mXJtE82CnIME/BonygTekc+BNFuau
H0sKJhJkGFNMOju0lS4y/CBlRBTRhlZx4YT2FMzHUS9oNMxDof1/QutXW+oT
neTZGt4p4sToYJM6pxixY44D/PWmQoaVbCUPCnhgEeBtJRDjydN3Adx1XTwu
IY+PBYcBLVtNrkJqKDBftZHmWFGLl5yCgeLsbTPqEhpjdxsJfoKupB3dO0yx
osxUgN36C0c7bEEoh3Cs8il/dPUDrs03lB7soG3rRCVXCXj1qViYyY58uI23
ZqWIbvvp5GWvexNAF3JBD1ExRNqUmMG6+P025yw/Ul3KQUsiDF9+OBBm8CoG
XXamhQiSret08ZQ5W0xFk36Ld28VQcChKSBtFZChr2dpn+Uxg/fRxV0/eGoG
yRxaRAYvxOwlr3Z2Zm41l6ijsW0z8ipRgLe8FMf/fOflfMTRucDnW5hQ8cne
RGB9HeX49wMVOMY02QJpCyN5OXqfoqNcQ9bzEeI+LOUZ8z/3A0qSFpiX1KCj
SGWSKf+/c+JDFZkxRld6cHNUi0Zn+9freFIbV4OpGgGMRk6YeIvP2mj69ZqU
yQZRONEtbND5B/fTKLDaiFFPfHPFKjfMHxO3VqhQZ+kNH6SV1ug/9dL7Bj2w
WnGPz2sC2JRkf3pUAZc0HIujOrUGIpkGRfhG1zb6UgNVIV0ZJY6I5OiWLnND
ysa8K2HxF/vzzadW5wiCiOKb8dSISzFMVXmIpi2CoRC1pJyCpm2ODx6Im/IF
i+MZWMTSjDK8c6dXuibCB26y79ytiZ8eR4y5Htzww0w3Qlt7rK/eTIai/nQi
GhjfyHkAuWalcH7WPNSPWPBLrdlLObK82V0iCmKluNynVPy899UobwSO2ov1
xTMYiPZ5AdI163WYPOkCgIe2pvtn5vw4bopcsAuDDYFEQuC3iCK1eO+9dAsv
swlvDwqNnkcODErwhEnqYsTQUlXe1tBIVTL4NDhFtN1UJRNz8ub65d1yqmoE
eaEfVBbOcgNXniWnch0lvuyeOQ4UztR3uMbLW+Wm8b3kRS7GR/IS06LxwYLQ
IuO+RL0YrXmqcD0969X6XV+j/YA1dRnpvfltOU2NcqRzK0GCnKLR2g+2PM1Z
VbpaH9ZbsnEvpMNXfPrTeh6JEnoN7DzVsZv6eBbahPM071H4v9kC6KMMHo1F
00sFv1UBB1eroa9gSqtQDXkHYk7Ncr7RrjNZcSGNXP0VdRR6huhDWS6kRhpR
DZswwcD/RtBbObd+nmY1sWL1xWEG2Q9mc8UO/KAeUBWLTw0h3V9slIR873h1
T6xKtguNiuMD4Nd6i6Ws3PbEFCvQPL/X/+nVpVeSoMp/Nq70HLGtjFcDfeWX
6uRmh+lOWS6MRHUiYEv4HLAOm+OS+hSZwErd60ZZ/iJw0YRCShORY2GEh7zJ
E4CwCEUVoYgWgbbLeFJvZhse76iCnESMTAAk8qFxXUpPJkIXYq3I6d19MPXB
0TXwDf+m3c+JgrjSFvo+ObIJrRsNL+kzrYdMF9V5sMR8/V1hSC7G0VPdBGEI
71AP+n6O4v9Dhin/KhQXhjtAv6NVqqkoLjwnntRWbBg4iLhIH1LVA+PTD1TZ
8sHzoGiif84J3kjPy24HHsviNqcV8U7Iht5m1ue3OKQ=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyL3ymWMkavX1/KjfaPZmbNlRDeoCTsd4nlJx4oV63Hv4ncfA4Iu0mGDJabVut/JGSuyakm04FSljztlvggIIFkT8P8cnJHoBlTg1JXxIyyxBcyysTdaNmDgmiEZW2xv4hhi4S3hHM7yTTLXE2hbLGnWFuv9nNYFoYMoS9XlFqh/wRL5ReTuWc1IpoandFUj9YsJiWwLQnyUHwVEJPxXlPcvvwV3OEJfC0W+8W9j9XXBSsj+5DhzpbwsGPfB6PtKdfRVxjVBR8PmOL3RFIiiLsSUSvLjWtYrl3K7vRbQlRoJHtSksAoAurOz/UI58FsG0NnvSjoKebD0zHg7BkdYboNgiDkJjp3nV2ADKNBWxi7n2mugaNQUQ1lMjQAU2liiEClj6Immjktij1JMIgin2RK+k/r/IccrjqMNYO2pvDJIKMiFDMloK6ivAVS6J5hoTR7x/hfaaVlRF1SRu8wur8Cvw0nIttqGwvn5/mQFYJ30BtbkRzE/tOqk/yAqKQz24LdyaN0cNmtfXgnw0S7ZraExwhn7Sxdm5W8PM14rZMShzAGoNhbgeq9w2YG7A+ZsnmmG7jePvWWXmycIkVsePaQVfG3ZsMno+OzSU+LaBgYJQjJuGiPF8+GEajrPumWCFjtqenBppdghTh0m04/mJseZti+OOjOE9JmKSu4ZclVY5oVIhzq0AE68y3g9KHnYH9QFgWNMYwjHdxNVWEBTz0BMhz23waUuJ32FrJS/Y0qTXsJHVEqN3AZ8+k7fJkNphMJvAN6skxW0O/LBb94RKrEk"
`endif