// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b2Y/CirkZsndL2ThfijEQ3hduNsFGjWR8sH9ckYkBbT67nLRM5UBcpeE/AZC
HX+WwITxxsS6koHoez1orv0C7sd21o/6oBdc5xyZg5iLLSUESqbQUUkHfkQZ
LA9otihJfh8NOIax46wt5hntl/FaYQeq4qfn8Glq0mFMQVNHF879x8JTvzXP
YNmYcFSS+YsrMq1vVp+NWwbAS9bd3KhEfs72IfvWaSTf6TbZntTpjslaxcc2
gTfyIb6AZlPsmo90V/Lg6eq4yH8QR7AYsDcZhmXHgP0yywIfCpP/Q+Fz4vyA
tcHQb2U734aLCWN/WJF6S3nvpl0UOzzX4/nHl1YeHA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n3ynBBsykX1t0GQ5fjyFOU5LmRjGVf0FUhoPbYi0r+neymysvPCbJ6YZqS2z
zh7xip+UipJ4IWEv7uyHD5AR14omPWOsvKSw2fkbyV2RZqMHs8aFZoPK1Gts
g7g3XmpVJVaFJEvIy/HOyE4fRC6dtbdUqMDOQjGU8Q1FBhdsK99NrMLALIkL
vA8VRlkypbP0anwixFr459WALQkIFe1TZm9gn/cnlkImWTIFPiFKt7VMvALH
qaFhOKl46T2piwB+U2e4aGwo74NaD9+6z4S8qj2siAbG7VWtqvpBlqbkDLSJ
SV0vpmFN1KEGpZhHQkNb6UnAYuAkC26f2A56KqarSg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GNG2N2oNZmXZ913IiVlYq1lB6jJVaqQQ/9iJ+SpWoLIEguMKapeA3gxhE3vs
+Vexg19o/n5HRPiHpjKQ9YVl1muCxQnhTFG5KxCIIiJIoYO7v3xn93ufaQzg
HIU7k2uyBZjtsQZt1RC4M8sr4OTU70LIMhGEcfTobyEPDacs0IwXMFJ6dLs/
XDbNVolWLjf2Wn9TCJNmegxRGDHjW1sSe2tweKFwFUOlKKAv6SU8PPLLEucV
pm23Py0J/c+9VQBA9q2O4eEn4gF7mR3dTeFskExHIBY55CoUocybD5uMCL6g
awzBbtA0bUZ6wx6mdimXmVbUWq3h6oQgB2TAv7zhPA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VjUhKO7WbYo51QmkW4N39xRzZTbEi7qiK6+Jv3Rk7CKnDM+CUhAKBFUiIudL
Q+z587Or+TE+CQSHFH/YQ9GTvXtRVGmn9TF6KE+pgF4Brid42kj7/2jXmze5
VasImTvFasl2rgrV6dOR7iLwCbryi2jGRrHwXXj/OLoViIuZ8tBn0JHivcZ0
xzPDai9yglGygn6TLCPJ4/BgGaMsycoDscXsHe9JaBAwyVBSvZ7WAOtq/Rb1
k+yUZJntm9jplFiRfLHrAUbw9D6r3NqPUHyN6XCv+QMDgfP1y7bFa3JNsZtM
f3eyGAX6i6BshLHAbDOaf/UE+7J1pmVmL45abZT4Vw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
X68Bt02aXNo9QPS/eTi53R6oARKq725lLxIlYiNcWkCpnQGPxwGwS1OHwCxR
6iiAozYjWqgABI2YkK7F805llE+x6kIUx+L9GMQ03kPW4w4GS65j+G6KMuSZ
1oO70X5p11fW8ONAyFCU66zKUDYo3ehp9+hs5MCMclE4zSE723M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wrb3rTWt/U1jFH2CyVOBbC0CsYyYEv2Jv0GcM2WCx5A5rbqWr8DQ48jMcjXS
cJ9ulQJ2DGj8ZgFdwyHt4VwlUPtFU9T4+WTFx6FQ6UC5eCUZOK44W1lIM0wZ
fuGd5/0SCZOaIqI/fPpxQMCwHk7ZxovsQYgFq4+JjwwUisnvmrrAKAbTHRJZ
xc+sYxu4UWTFXjXwqC+rAMPIPM+GMyCiwENPMWhmHD9MM8X4s0F8YYMtFR95
vrJZ1ofNsy7AfeGi+0gJYk9f7t9h/jCZcqH4SYmSdDOGOQNRIhv3GgFNYNmt
9plnH+IZarMZMFlFB3WXcviVXI6r0ErhDvlYaGQYEbghyTKW9mleVpVCFWno
url0QevC/iVKWTU1H5cctYGlAVtxW+aCZnY99vm7F2y1ObDa5wkOEgNlwLqZ
sXbohLnW4IbL12yb8CAoE+Fmbxa6A8X3dwj063tRlDUmXnBp68YAmr2corR3
SdN8xXAFP1ayQhyO1bUm/C679Ytdk1Z2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s1eGZvw21L/WYrXIjmRZNNc+JQz7/nxNI5IKkPPcFn3YhLeCjAHSg6gJyCrM
redakjzim2+/9DTLfWlysfiQPgCSf4INCHpy/bHIHm658mw6RgAdgzEfWpvV
Gru/CzJQ2pk+auKjwbWKoLgkO9ObjvntNDGP6XI76z3QXMH7pcU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m7Isnkv+7ItFRp7zP5iB9ORCIuJg8KOuyV4oZLUeXxKyTG9SNLN4XF4BrAe8
gz5MEAg+2ouW1as9K+gSqB4tIRSUhnmaX4R++n1EYppBg8m8k5TKAs1/6FBW
FvJ3So/7x+Mvl++JhHo5nfmuX5KdajquynZLtGXJo3qYLqdCvtM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 76128)
`pragma protect data_block
k8ymS4D2R0frccrS52FC2tG4RU4blnTDULgbzCLrEWUJdl9GnXsTaaDISJrY
PECK8c28d6EPwbG/DorrcoA61wYrKkvslZQkuwGO6rISnW3+5RFIwAXt3dLX
N1kn5DAjieQILXSj846rfr1xmt4h3n+OhRKTX3zl/11mtkC2AJhuCedeF3Ym
uk+r9+5WVpMVo6QKiFRlOV9Q+xZ4s3ZrHl9GTKTNmu4N8zUdr/KHx6h0Vjiz
w0bNhw3bbFhfXurj1t6xASzPrHi4JncR6tqK7+wvOc0WAS3o0Jpfk34RYo6I
KKXDMO8JLgDIg8jwrzylcbq1lis4V1YQs4hB9DwkSISkgsnHgt9aWz0gN4Sy
r1dg+IcHbRHZWDY92V45kFhmLq/3aFMdQc4IQgqLnAqpTxIrfEXNfpP2ttpu
oWUgr1IEQvQ3hjZYbFoYMn3yM3ToHmZAWej6HmxfvTEgawZQcAt2sX/Svmbt
MlyBPr7bVp6iMvAsJSgWO3RMBR4I9zIgP3HRomUh6ClEuP0AMBuImTRTcRPn
l9Ow+1xYNJ5D08ER6B+t5kpG/GHqtLbH8zjpdc3Apyyd603YYALcYQhDKxi6
yOj4XRbaVicpA6s0sf8cX/w+QPLruHYvq3yj8U/dal8Ql5BBWyQkIOc8+wDY
Kv3vo021D7d495RELigjRTQIZiqTiSHpZrWHTBOQSGGFW3cRNtiLBhedZTFh
m7C8RIF2dza3D2y/Rk7phT2YeqOmS+In13V9NGxD7PlGAJL2P6Sfq9cOne53
ibXKZPNO6cP3oUDIi8eUgYDSfQQ4yav3D8oiFfKYKHYQJkon/QtbLTfrhbG8
vj38lVYvpPFU68DLRHoeuk9aKRD+IWbBgueCrhlyLpFIxEdSN1zddo+8GJ2p
LxUG2nCr4S2emT/HKimMSBJGVVUzL26v3eK+tV7XAPsRphZ7Dw3pjfkMGsxF
bILnT+e+0Vj+g6vERSvGjB0tA9uj8/GV4Bnv2E4ElyLtzpj81g52AHgl5iAX
8TBhvLTE4jWuhQBbvY3oSbrER/9eiqbjQ2QtXMyBPB4d4Ulqie+BrFmeB4oo
5rvhuWYEGHdAM0iB0dqUCndcG3aQuBEHSggU67S0FjnAQv8E8VKQUbESBCrv
i+WvhIdYgxSnwrwZ5wWIPCbVYt2kepiv0/H88xhPHSPWaAW/SGFsGTJsTNkk
nSaZAlLg+RfqWCZhL3Dsm51DSEEYTp/ImJdp5Y/MALEhERlMH2rzMzKw2R+x
Whj6s6UBoT/ID2zU/cujyY1TS71f4J9MfggEzHJnlWHyo8vURyOYXhXa9uo+
VlLTNlR+rG6O1qVMpwxP8PmtgYoRwizbrSHVapY4usdjTdd5JAefkwQrjlv1
HDsywOI/fibbCMr0nJ+s3q+7wgDK/ysu86fH3PI+E8tGpjMLTIJMZHB4/NuX
91fK7izkzgSCZ/3J7BFBE5YBidtyjMMPSDxrB6ej27BEtKi3/+AyhFMr5PlP
J9/Po7tu/iDrEwV6tNaegPyp0qgrYyDB3Nw1dq1DN9tBS1A16u2x9wfq//6l
OxR/IjyEAK/rRwveiIlEd2l38hymgYMm3/r4dalVexF36835uzqVID/53pN+
BRXzAt5Rjr6UjWpo8eEHJOJDRVcqHw62O4o2Vn3XjrRBeXgbC5pL4Avei83o
ZfIHm6jUSf0VVs4itatkbv5vrNV9O0ueDYDiZspnm2qhWOMjf5U06drlb2Qn
LMfQ47Q1XCHI1kFSwZPkbkSJRppXev6C587ya2CvOShY2qY4oe1ioJQhUjhk
lKwIELTl+z0Qaut4IQir+Gj5lvMql4J/6Ldg/evRORNuUtS1P4NqVBjuIOQj
OrAgrhSmXPyiiUhpLXRCjWSX48FH56phQrL0+XXnhydKlVq1VlpJPaZzm3Ow
A+88Uifgra6RAtFux4Zf38msnSmzALCAhUBEW1/dIe/+bPX6i180WaoVtIhl
KtAjjMxInBV6iRDVFdkOtbQMOKVln64wCUjqnsug8o7QDlut9EzKvFaHT1WX
oGGG56V3f2ijEdVrI8C3GiMmhomb5lV3MrSa6yZHbVRQoMJWy59mmMzczXp+
ptYOD0t1uQB2drZ/eSsCmKRSx8N2RwPqrjJkP3n52hKvDcD02GsX2icuV9MJ
LRUhOqFZMaCVvxZrEalLydRzGo62OenWZwJZFGkep65CWWKG8wIUgfGmq+b9
ZOKTfZP5ovtKjcrTKxVktF2s7CnykHUocmd/ZjjcQNPS7My0ljqvILhkW0Nm
Gj9SP17LP1h+19BZSjs+tjVqNOHoRhpZQ1a8BjfrmV+AlIj2xQeC8flxVG+I
2aONuaJmC5NZgMWK4SZtvyRFDXs80hfhpbaqQLKr5JgpfbsGbIkvqmeNOzO9
u6LYlOemX/TIrVak2JcLyB3YqMjCsW257zaRiSdNcPaV8rH18QYxz2x6rzNG
x8qZO81v2iYF15tvswDicCXrZT94VY1WbuQp/7CdUnAY+3H1QPGkzD0y1xt4
ktj1VPTn0rIr0SC5MT7YW2UerFtnUg0OYdNC9mZ/3VoF9NeWt0kcnlJV3egj
hRXr+H9inhk/5JQVUdIsy8J4cpgBj8GrEvqtvC0RZinuOpCIrEx1OGVNWd03
hDPggPgLEkxIPOoiDjDx1Q+xS8dtGLMYIvo94U53xruRnFmq2QrbU2y6Qssp
F1gl65eLtVBKZuBi3xw+6cpsTgbYx59m8DS+OmDClIywl5JinNk4EAQ13DvU
XaE3TRIcr9DJuKgZQjGpk8u4yiX3GcbdzCd1rYtdY2W1r00kcGaX0K4matB6
cjWYxAhjIk3LXtpSIqE5i4qrDytHq9THfhbjvi2lE7kvYj3gBiHtPNwDML/Z
TZIenzfJqVC6pojz1d17qdIXkyOwB4WQBz5f29xCT0bnpliz3akxIX/z2g9F
cbURNBiAZgbn8mbejafBPtAasdB1vCc7dioa7Aa3TXB1ZcuRJl11Z+nQla4c
L6n7YEqKczMARUUn10Giub9fYPED1WL+Sm5pMR5I2pNreepqWpM+NsM3aY67
y4SbfM6cdeKOVJEtJAEVOe0Q7AQ7ii5Sme7pKhGzzDwWsXfvLpyfAY4mmrt6
NxSQMjey7ONwNQdivUWUWtrpwi9S1u2DhsqBUFBZ889IxguhzB+o0or/Wwns
INagR8hU2sXHzQfV14Hy3ryeGw1cNIlRxD/KEXRet/ls2oGDcK9NeBpGzegL
gCIFMUg3/LoNdAY9B6tSf8DkHd9uOK6zF8KAC3E/3SbHvRWc7iuwCiXB0h9u
CXztSkX6DtGTRCzae+UOgluv1AkMkHHLaPUSzZ9DnDAmLCjbOb7uG0vwTfVo
WqnpZtw/qOC2mWP+DD94YU0mjrNOeptCo5nMCFLjUauZ8GLu4TK/WlF1/ICH
7W15r2k9lfLtfYAcijXK89kgQ2XXTF5qAZsMaNiPyAKyAceVMka22550ejpp
2Co6Y9k9mPKHlZgcJo236X/USAHrAIwQsKqnw6gNwJRtk9crf7jCvzKio+8x
dvF98JuEsWhFD6ScdPf5XNkr5fkuanAeqPejXfx0v6yFs6zEU7elsNmtGFcM
1FVBpcAycGHnlA779o6HXs/XnkUIHWn2ET7vzkN8+tzn1jOaMpIEMWczeCrs
/BkVxZPTPGU6f50y4fJgU78KhdxtDlOAKd9dn2z9WiI9x4fz0XWFh1UZv7M9
kXMuodW74lvpAv2t5Z1ai9svd6/oKG7f8OF9KIYwvUl61ST+O1AIa1d5XLUR
UrfPmZLB0q2RJ58Wcder94bPrUum6ujT0P9Ya0hSY2aZZqnSoeA50F12CuMj
AToovwR4QpVDGYwEbhoyC7cd3W/deV9LAwISNkLC/woGHC1fWghveulYbvk0
9vgaHEr4XUjDsWQGAh9oSZaUnWk4TsWIhOL5Mwe8Xreq3be7btKr+AGqGJ+l
NF4XCKKRFrPrpxRvmyJCmLP9wELqhzzowaXOc4IAMYIVIooJmpbrzRhZzFGv
o0aAWpQ4G7jDxikv/ibYGcUico82jX7kGVHdAzxMFsMydOXekxcydeiZZ9MP
sIaRvgBMiIx/nSUS2gSqKAf8kLtxRWn/NC3opXoGSS3g1SnMqOBPdOVAd64p
OUBn5NVeroGFJfZJqhABXh8uJL6ILGuDPYRzKoCZ74X+o1LMkBd69l5mVD0p
4qp3Ck0JDS1WkDXAz7dEjHKd9HoHtDYRQuO+FbzPT+mQlFynhAJgycLHwAAH
Eio/46OeEVyn6E+9BzmTrKu5ru5hApINdBcu95pBxoYwdYR/qLIfTO0nUAo6
61zGXJ8BlYZs+1aYsoOXnbcEL37ZKkIYwtNTe7AdL5ks4baiEVMwr9Q3AIXL
VvGLUhwWBrM31OCCWeGfCZO2ftHUquFhBpkey9uQZqGIruLhY6088tuAWTKU
S5o+iBnUuqsm32Nt26G3W21/366n6m9OqpKu6YoVZQT/EkOGo5FIqzM50PjS
itrbCn3ds3mE756scSN+XVrvU8R9dTTa7rnxms5BlsoUqwY0RC5p0nB4986L
T8LpM5Cm+U399q+2A+FA/wXUIh7t5UizybNPfriOSy4VSdOUPyAPa/vCzKSd
g48zlwrSzhEpUpbByojWm2QhHRM70+ZQg74Eo3TPS2Yioan9tgKsIW8MfEai
njtXXOOsz48s3dU/4mEWuUzv1EaEkqtQ/Ve87Lw6Bukoy7p/uJZbof/Fr4To
DrmRx7qKUebfJ2QEBXrFiBb2YAb9iBAQ2IyyLuXWxjdpZW/Nli4f74KbVlwe
7Oszsz+249ci8yw+xvo/2FktcGuNVl57AaKTfxOzCod8GZu75aYOEfPEUTZ9
rMQ/ygL6g9QyyM+WXHyQSpIC8OIDzam7hgNfFc7sAO+RCewYKw9+GesM4p5D
ToLtcyy6T/ICQ0VtCHK1jNo+qeN2c67oVtJEcEte3fVXk0IUE5LHF87qPt4z
NqmFP0MtK2Dt/00wRQXiuwwK//VWO7GZWkWwW4cipJYIGXTkj1SWxUkSucnn
Ze2YNjBrieg3AOtbwK15zneQmT5REc5NqcLTFYRBeiY+AEy6EAF/8LdPmYQ4
ShC0+Vk97sPxxORva1Mf6MBVau38f8NeowCx92dvoazVEFcYU/gl8a1EKxwD
xMO/PMkNkzTzCttVMUFsQelFbf9LX8ncnQ+1vxhbWb39d0PcbHkuxnbhmvJB
kNwXL22QaXtxHAQRJOq8KQX8XAAXWEdz1zer2qZ1eUJnW4vaELCxYeysyFK/
go6vf+6OxzgLHaIQhSX2nJi9BGQmc2xtDyOFzAx9nezhISoFCqpDb6hp/N69
a1oZAfMO9/zrEnGmWGKDaoY8pfmnGqgGtgaDHYp9atuWsc2TVwoO8hUTdESl
xQMw07ecGYuapZfHyrrqbO7kQbE7qlIwxJRp0868bzARN6Z4H2MZjQUQYXan
8vYIEsasPGZ4dvp8aPTX81020uDTBqSQFtJ8fg7ljovdLYcFOukyd13vyGt2
LwQ5XftZUPrl7nKG2GeoupaaujliK56CzssaysKbAh9iweB2k9T/IK49taGf
qd/UgKsSoQzVJ2vGCgtTOHgX/nNC6Wf4WpnByKk6ou/5BPbZBshR+qdpy6vQ
5aFYWoX5UWdCgRDdRouPp8QzZUP9pySJ4fr142a220s317JRz7PDVIeRZJmC
XeVRdvvCeaerxtwU5P8vkCEzf9NdWotxIJ6VJ1NYlQOSUTlSKDAMiKv2sX0N
lEiJoGlTWy5O83V5Oit2bhDkhvpYv8cTJCsCmNS9WemMDdcLOLKf5kArEZGY
FfoQbKxMVaTXGdQhpmorMOft5BxfdG7qFE+/Advrd7uGQFV3wJNRSa+eJybT
8F6yU2Dx8+fGE6PEY+IXaTw/TatZhHA58cQYwpsgwsYWdgEsRxUC94rimfgA
+gZrMCblXwC4Dcnk0vdOYsNq4DOfNVdhsJazcsN5SPTOXoETvyBURICPREnr
J7M4WAYlzIUnQh9hGOmFlfn0ijIGyKYkjYdS2CrpsB8lpRhZwjuE1p8359Kv
88ikpr2Z54K7QDq7ItxvVemLH80OpG21xqF1BuMd5EsSxPZoJtvjaD2P0gn9
74VoQY+TADrnIqCUeHcn3urhBDEQkcPlJV+eCnsvD1w0TZL3gX6jJGBnEbj+
qj7TmI8ynf6YrCJ2dogR7ycs7ylUjON+WRoyBTbP6+bwsNqZaEVDGbHCIzIF
wWSNC2U5hSca6zMeyTjPqNyfQKgiuiVmyfHQc3kVvJaeaVyf0Y0GiYNJ6cWc
mvZzZgIH/OnS8AykBocIEo6WS2WHxDJuTwqutK0Gq5L48w4lHjx6yB4PbIB9
CtNcec+JG8H7dGE07EOzg9c/AQVHULIWBJcAHqnD81Qp5C03ejAPUU29kOOh
0elPyZJQLCCiepCqXaOuCez8vyOam5MbwzCkr2XvqxlZri74cO5Q2l7OJAb0
ZYHXx6MAXhlp3lFzf5byd9UNb9TCqYpxp9xzGUELzLIEhl3Cyi4pvjRcufec
klOJzJgfxPztZJZMEnRnMQ2EeUtks/e4dET09u86r0tiZoc/ecSeE+7trVmo
2314Jb3pNTWWT4bHV3sbD9AX+bne1ELdwstPi5BtRMMN5znil1NHIHEY3+PV
1sJhCjLszNOKOrGaacVjRhlPni72P03JItAy8VcbjPjyG8o4gR+k/SCXWS7T
8Krscl8hsAJgh1WLflCi3frGV5etN6Tt5/DJ8DDpYWoyH6DBJkrbJmFhwIhp
8m7YIaqqIVZD5OP9Vt+QJKsmUs9Tx4TeNU9qKVs7btP10RkgcfBe+8R1buVj
lRbe+PTND1JkmAklgHbZWU7w41d4Pj6L+74rmx/DESONVQba8ou6bYHgWSbS
GCdoz2sP5R8rf5DChOO0qjt1MFCwvl+ip51ZIoBKhJYhhqeDr/YR2MJoI+7Z
fA72mJhXWgMSGKCxzFo6EjgJs74TwHYWWYQqqrzf8/SlcUoV+VINQCLab7Qh
YmxWurcOOZXesC9YM+tio1MwIRMcJ86LmUVfEhMZNYtizToAmEsD0JIP+IrT
3VlOMmg+XEByXy1VZKygf692OxLbfMppF8SbOqIBr7ucT7XkNe81hX8/mea0
EgQtLJCpvemOUpJZdcHJwTWB3z6D8ZNPN2cDwnPBBjAYB8Thpb3846mDYQnv
fIrdTNgkkO7IVTH8GatyVnifSo/oadHplHxR5/1PMVGzUsqd/947EYBzvPsX
nP3rwYBdWvbDYRHq6cojz1rxG9oeX5sL5qauHuPPaLg+C42jawsrPgJdY1Tq
o75etO4i3A1WXNCSagj0DG+bXpqV051NduNJd+6lQGtBprUJ8aBCq3EoooSc
GyOsm2s/W+UF/myrP99tM7swaa2qnwESgB59SW5KMvcWgQJQSDKqY9M9GVou
Cc9JZBsL2GCLBxXrBxE2hjzGLPHWaMqoGpTuJAq08hIH1zetcTJrs7rTZazo
/2oQYhTvY4sDgnBaGqxINUoG9GWp1qHzEV38n7Qo5oPh29n5HsQJO+RcnK4M
3nbyfaPy2bhlvcdfxlc+86s8veoiY0Ei+eiRkVvucA7ckvnRXPtqEXNYuSSi
L4OWur/j8wue5RFkbuXmSqvA99lnuILv1G6SSxVaLkE5GwIwxIyGx2Q3q4vN
1MisQqfBu+TqDM3U52WdKUdwc6fddYv/NnWMIrYHYzAaRgwCicAFf/FIVLpq
tbH00vUa8/zws84zi3IIl7+U9TIr0EL6UJCFkBpd5Ce0+zBYcJziz0Iuk2tw
2+ml1hnRw7GPSS7ZX/y5UsMWx4ivn0qMS8wwMzG/JvGcUoEg6GJIhCE6XQCa
UsRBCFugHz4YJk9MKarRGhAyTxQz8fU0mfbAOjOWN9h5SMbwFQ16mTD3ArZn
Qxqv3p/AFN/8Hcb94kA3JErH3yguTdTX/r9fdwEWqNUllUUHkeqglxmrykj0
u1i5PJYHrYE9Z+eZh7DeUmdzQa+8F+4ImLNCYKrrjKKupnmVoWLHmqWVYy0W
7J1lBjMC/EEB4LLq2ShMYGderHYSd+u+g306LMiQUs5muPXXdynT3Y6SiIn4
BOJBqORN/rs5VNBjwhdWm/IP+eIxdxPWwhHqQt6cvXtfxfWzyJntz4LzMMAl
bJkMbEA3rwuA/COT+mNJf5mejhySo+hf0piWl8epj02na41QxQPCpp6pEIoT
jcaTUmD7SRc0luJk6hpfvhiRsT+AYKuvqad7Mb1EJfZqA6D8+TW8kRIxnUQs
jsOstCehXiwkDjKv5Jd8aIyHP9tRNzuenGKtXoQ7uZnMcmvhJqMzekh6B++p
1R7XrTtHsFQn2P3ws/42uxsVdccaOh8YdCqrSz7EGjLADSe3JcMGtFculWhN
5w0CfUz1PneOXs//XyayiLKiZe1GMRv4CF1rfyo5nKLLg9uucKfDn1fjsAYt
YVGs1Bqf9Eg63/y6z/ZNIN1wlRNMrWjqeCmTnpabynRN0i2q1gCXeMZ0VzWS
gz7A8eknYyjOwunbnxqZasbqxCXoY7XUWTFF0fUgrsoxaCEl79AVL5vbDANQ
H7nZ1uCEFBDJa6Mju3YoxnKuOHWPq64TxyukVZT7SYELzyzjsq7WkW+7JLo6
c0c9wB92uQh8sb4R79bx7o3nGj0mef2+Wr/QC4Vxopp5irqlY4g9ZvkCX8+a
LH2S3LMUk7Cts220apgvXHHFQv+/gH+Ay7mcMTo/ZsR1fswGR7H6Mc8HDswT
rW/RmLujqhhP+yEfa6vpZiHjohjyaw0YfcM4Sd23Fzpevyd91gV+DGn0zdk2
YdhVHHzfTWLs+NkFOrnfRLeyzHol27TfkPC3Owl0O2AlKbi+EkLo8J0G72et
QIygKxP8AxPmP5nAmdFDNcYhzPpUAncX+vN6AA61lySliCJxSEqwiiVI6p1B
lrqD+NzEuo513HYGpo4hI3Qq+MlsQEeKnIFyw9gYhwVNDvrsTlsMS7SueGOv
v1hWGMs5qhd0DlFBL1tvcY9G3/HyOE3uc/NAsag0PBzetZA/Raye7sfcYJZN
G5sHp2Jq+0gMLFS/FhxAi/lmUbSw0z2eVC3BCG/Wf3bDCbxA1AZwug7DLOV5
a3RMw+/urDaPPifkOSeCMBMZZtpzXa9wa5r+GMi4EbI43LO3d5wxqQZFmWUq
jfI7OsilzI9cx2OZ1ETprl1Kq6PKuJbgizFI4xpsXn89VNz8dvtcpNfoEJ0h
waQpitaZppjLiWSZjlGgEVZRKDniJTARB7mMmUC8CPbmyqFTGlXnIaCVHsD4
jRvzHMnyPIw3fzuE/boUal21demBz8PF+7sIKI4+LV6J9fXxrPUheaLjORHq
Qk6h5SF33NBGtDPBG+aQB6oUNbzFpoxvkAGuK3A9PdOFi+5UA6ZQCfVBl2bi
wmQToRHsJbC9cjwrzhRyRHME2EiBT/1j4x+uDJ5yz+/kYTraxxe7WGD/tZ6O
imSb883VPT4mwPvAHgYnC7Bx4Y08sxHTl8qM9kJ2Vm1P8o5oONK4+hW+/i71
4cIe418ZNy2SNmdufryBSt1MXYzXIV9uoSkLnTibsgFZlj2LtlpdSGIz0ycJ
A+xBAr9MR9o2GZdIfIEkzfngYgMiBj0DUWPlcZJInnWtU6EfssOuaroBa+BO
reIc6fyg9Y0ruNLHu9AQ2pi+GhEiQUa1JxL4RoPuENehchX9LpHhcYNTsUZ/
5vTYz237IUu6qIZHXnVHPahiKmLbkXjpkia/I2JfeTHag20eY4YvpJzy6zKx
9QYRph3FumuvkDQjnShS5gQSOjiBElgU7yERWa7nIQ0LwvRq42Ka0IxENN0y
XDrqogAZV0E4JZvBdo8n6sxihogYSKaIAs1sunXNlpaq2Q/jjtZZOPAMHPSe
lL3ZpVn5/sxiW5NPcrtTd2b/215BQpboiU1q3Ypk37GkRQcdoAxWO97QGCQc
LUm0KVRaBVZHxS+11ydnKksXMw+ERoi1TDn9hBy8c/tfReLVQ8v0z7MKj9fv
DA02Dp1J2LLlLl5DlMsY9f1SGwd9GrWWWcIsQ9qgLN6PWrZlNZSjJOmhgC6W
C9yGzjdg0O4KnyXuCi/AnqLMuelXpQ0g7BRn6xtY+AWt+kAqrw0mT0HpNTo+
a0SH7nCn+lF6rnRXv6cJi+rxzSqiI31epiA4RXRs4s0y73IqDuIG2a8+uZhv
Y3PlkTb9IcUpSkyb88JStK0zb4c6bxxSaGHI6tV2Y+bJedcHXkEOrRbA4eaH
8mGdh4hYGx12AGR910Lj8je3H7Rfio9gGcIZNwlqm3uM6izy2OBnaN+3H5Ha
Sxx/ulN4DWJ84eH8kdrGOsqmPA8uPF3nLgGtbQLzsxsGyWLDl+PbEjgp9rlx
Gmc7MZfjre3JMs+AlUi3m/1XvunXshuTEZeo1GIl84VRVdx1LA29rZFIuwHN
G4zhlM5flts6P6UTVZd4mLLklbTyYJfEZH/mIJ2Uw98+EcCeiqgb1cThqNBI
iOcuWKHBFxLOu9ww+SnXZoV0ZNUfEXuAoD+ft1zPoTBEW9rQUnNsBdZxw8J1
ZMhrtGT5LBBFvVatmvJ/8izs5kSxdIY3eq1OgUHUVH40GfIlO/wYSrTcyzDp
7uGQ8l22F+sTQzpsZ+/RKU7oyF1o1lfwOgu030JyQT9qTT8Fs9V7vDoSOPWF
IRM7BdshszprrqYbaWPOkouBty4q2MSaVpG9Ae6xxkPZKh8td9qoiZ0G88or
Sb1Fo2qU+BXMLqlh+VuTfOpxDZqt47HUcT/3mg1lNRsc2z75PdLxijbMBPmk
3P5ueFV1v1GPuRNOoj/rlW8UoFu7VszK8bUABg25JtXchn59SZ8tyhtwcoiA
dyuoYbgd5MWnkHu4/FC4QZg3N8KOPmhB05mZkf6FY/wRI+osb1Jn6BzKVnq8
RMVARG3wcF78Ev90ne8cYFknM308X9CKLqZfFuzK4n3gYyfYWS0uJ/IULp15
Z/wogZIceFZVr+17JyldshoOhirXyLiWXh9fj3bUdiuoarfJnY/2FdBbXSuk
fo7D1IslgVr9feQ5OfX3p6VnoUvLSpizYDB2Dt1DdUbBeMhusbroQpMEaExa
eOtLAKv2lZHpvY2V94ylGdxnEcGngudFP39UZU9u68DFEi3HW25RdRAf+ALV
/rmpijUwrFwoaTv3VqwlCiOcalYJsOCbpyxSRbqQRr11d7fFXmMi1srFsCbI
BYNraw/F0RKFlq4R34Y8tR/fuMkRYiv5txaIqxPoDCEHnJYcd3Y6Btcd7W5d
d+Y6QNuMZyV+Ou8D4+FKk7QqARoPUufZ4zZex5cwvfP8ZRU6E1tL/GPtanhx
u3E/LE4RvLi1z0RppMIf4lBZV1+8CZj0+LSMqAMPYcKkJ9L/OPACX4+nyifZ
BN4hbyNFwY9eMOa2d8PeShEmf4Q7o3ZyoFDIhmrIZjxoODGu1WOm1LG01HSP
ddSYt+JcCKzheK2IO0koVL+Am72O6bUoHFpwsT1hPn2SVZATFmwlXwzkAzVx
so8kJECiKBulyjRnSQkewfPG2h6Vrot+CZUONIXlDSNP1LFL284Vl93we3Pa
bgT0bNqzgN1QVyycrBpHwhiHb0VI1ZWF8IdXt8tuwCO62nrInQSlGUvvMKr7
mQeNeWQqX7ObuU04nDNCw7tZ2FOG/BNR3HlhCfzmCHmkULpuEPrzb5oU52l4
b/V+XygiX6pqDTa1FuwIP+L/1oeSFo8huIRJGAl2C1ua1DsDkP9pUA50lNF7
cZigedc0c7YEPIb0/IzmMgPqXtiGv1ndmjum449XkEjupl8TvX0k9we7fyv8
oc90mnO3EPwENDAN5AHzC/nQ6AKui1PqqVhLO78kgyXiYiBOmjAAez2ALMgV
Mb1vYGOzX3UBZPL/F2NiScD1p5+rcTIQQWIHmVXnVgy9kimsYKAoLW2rIcJw
ZLD73Y0vaO0R87Qx/TMNKgn9yiestmPy8CoFjXXVmJf72dJiyXOmhLplh3XQ
DXLPnnr9J3onJlhfEPVhiGUcHg9UAcfN2oZ9pqhmQPdkpLKX7vKfBXsH5eH/
WibxZ2N/iYgHPdxNtN4cgpcR7yYsgS1hvEfN8moxfSMBH4v+9/ilm8GYufQf
ree7HWOBRpOV8ZziItwTbl7reqVc9g3LYQvAsj/dhkPL0Z1aIf8t7kHRWf91
kEk10clvVik5zHXOojTh67bZCP7a8VruyKunfFGdIPtD5VabHW59hN3IVNf+
K/DyDHUYKAYrlfn4TOYvbwHe4IqEbyrZeCbcNtaXh9iu3eM5C7wDnnKOgXhb
tAZ8n0V2Iu4XmI7kdzGfF3wap/wLL9LLyFKgASGfpX5TWlX+G/Pzr/uY8s2l
Dbj6RcTo9t4TDFy98tZURvgyWE734HyKMFsbl2r/TBHmnVAzL6btH+rY+L7c
+bfqxFDu80ro53xXxeyk6Szd3dxJlcXRykXhrpYBjX28eDaXnRRbu4AtWiyb
gcxlckCx9lNiGXuDCxamQEXXo1NifR+QBYfJGd8jyAKVw/WIYHqi11eHBPhF
lGe2lRdlLsrcAZjcfC5yIbPHVmxzfajGZigO46E9TYw1njfb9akS2HVdNOTQ
gGlVlwB2neEf5BA3HjSonwRUjgtacv5eUWyK9ko3jDcEDbqh/44xElb+zSQO
l8LvnfUbSmmrtAfWT3pWVuUUO7QwEr1xe7co9cvfko/RmN2Rh56nzgkqgcZJ
CnK1ZUSZ9g8Y7saS0P0H+ytgd3STF5+iKmxg3loRmgGQBg14JHznjd6Aj6qm
pnGZneoJWUXT7+ANgOdurwSrtZH5jC57N2mu0AG23ZEKFKnlogbu1cSjsD75
cK27R4VsU4v8W/0F9v+F1u7g7uwdZvCPHJn2BXUH6Zo7GlXa8bht/suN2Fvv
Z1Tqon4NLMrLUyueYOhx2PKpb6zhY3+/jPRhFRxNrXjdTXOhl0L/1kT+mutc
zFYcSbiZG+THu/QC5ZSP5JLRCF/n3ek+m1CUWzdFim8RRQM/r70rGA2cQm1e
a2qnnAPyhh1dJFml9rV7DgEY5lkqN4juvbfF+o902FQPgY1QQcu40GNQvT0V
CStmxm+85kvvQ+yvVgR2TLJVMy41+nKgky2nbUm/H+g8GZ0nDIcyfzNg1yCq
fvwTy0ysDg3SqnRPN5fsxt9kERLYp8U+ciCr7tEpzMAm7AtKsjdHgqYQzclE
u92HIiNAPpyFJhez0l0o3fdg7lVHCLJPk6s+SJgAO6rc3wXqI2lJB2rPNQmI
rwza8Akzk/OTILv4aeGm7DOc9duGILcVKuwn/46glLI/132AVZUveN73Cvr9
LXj28B3O/xISqPVoLisb1dCXmPn8MU7A5T0DJsxR6jcFYdkl0QlX3IjWbAIa
lNjo1WwhCdl3kCnj79x048F72H4NXFtIWq8DvgphxkoZSw35yOKoWlhv6fcw
0+WUyNlkWUTCLpRyM3JbBgZXyVIgAFYnITr/jVI1zU4GmtWPExREy+kJXLnb
LgHp8FYq2yob6sV8TVPEoV78i7W09+pGBNktMAoLMRJT+wS1zRwhTUpFmq4D
+qrh3vNQuqB0ksE2kz8UD0oLD3mqg4JQ1yQsmOLehFoTO+FbDnwYQBWHXZw9
En/WUhyeiMjp/UzsLCJPe4t78roBbhLigvRd5Qx11r+jNGscHE/Axlg9KILF
e1cu2Pc2J1ewgRbO9Yj1jdHiekabPJCRF5hjjb88gHmOeTklUVAk8YMopnPa
LGIo6mVHu+jtrELRp68HKMOMP0Y/eqxWeYChi77+f1HGlMp7K9QtZtOhO7x8
gmQTvJ2baTpSTClz9+/6Nqx4uJOIVIGZi4aX2MZH/ecrfmAJx8hTVB1e2oWk
YX7waIoeT3K9t13UE+CI3zrpiNB4ORs5M068ii84EkVO0Qn8Df9HJFD25nfP
s05AQf56PuAlXyac1QiBs8lXTj8zF6Ylf8aSICSC1Nt3h+cFYePQbEgJEQfO
MqVqCdrIJHwgCD1WRTAjS/Bp1fvFI4bCx2ekwKi3bvBRzi/AKwxQh8LKSzAc
d0Kkzil4Gio4R4TsvEhE9sETpjCxXnUJhFCCH33B3pFu2wugnzuLJbJVUUZv
wB4kFiNNmejOuAYza9yMN2T+iC+nanrdMxSvz1ETcTmG3bCpGQBohnDcpsqb
w25yAzznuLvV07oT1Ngt/+1HG8/vfeS7r8LbLZS7mHit8wsy/0EWx1VyVu+r
J1CYR11+0iMaL8GS9s/eer/l46ZN1RLRRnOSNzv07VpLxMU3EudK4CInEOBB
0a8nM6sXBswKNg8H276Mpr2mxHsmbyz2LM9ePJQ8lnvsjtSJBIe3f1+mzpks
0eqfg67UK28DB3SA5q9yMZ6Nat6+TomnVdff7PVPk/Xn7Mq/rHdbHTsnGGzE
w7cUbqGPtrjuWSb3q7DIJnmM7ovU7fcfCN4NTkeY5YyHiWYIu+HLzcJ9jAMf
UBOAs8BwOtNmzvAJo8F/yvugv63rO6Qys0ChwxZer6yP4h3spsdetendPO4/
7MpRvoh72fMJiBBleFpLW4cBEWbkSY8K+/Yduy0027Gc+hSUFZntbLStYx9v
zce/JbIHwz3pQqs69EouG9NNUrbKJMPPon9txRRvxCXZAWe9XOfktcqiXSco
l6QbsoYolPlkmGxUySudI0L5oyv7yyQdv/bWUQnfXR7V8p9bB6RGF2a65Ix4
O8HHQRXKsEK2PwC18HTU1ChHZi/1qvFpLaT3X1J3ioX7LDftjDw6gUqVhodV
C+r0QluPDqvGu2Okf8srhoe8qBDnnigPUkWO9o3UUTRHHZnNc+5okMt7+fcf
8ltfXSyW53G35UzlZshp8Tk5glR+0JenzgroQCI0vUwpgP0lc2bi/vILUWOQ
5V7tbHLKgQJKyREnyL/5CjrIwGIGjR3dUjHjpBrmhLNrX38BcrevpqXGp6Nf
6rt/S9fTND8F7kP+ZTPG7mZgvMBqdLDzMsuzlt4ssDcKwXYwKs9ZNeWY7IXK
uJKSc27s48GpBl9A7vRfTche2QlBfLQH6V7x+OgNYgm1ji9+d6uYfnqVQ5Lp
wUxfH9UWx4SdHDFI9yk3ThPI9lJMhJxMqVqk+qNwTfGj8HxVsbNIaqNXj9Hl
ha9jQcKfOK217QoxF71nhLb1qJnkhxiJ4ysdHkvs3H7IitE5V9eqvLCIUYaI
gsGixFvAvWWnxdcAiN595bgfhCQUh+aHSDYq9AwLt18L7kaqPpIq7s7RBuyL
CBQZPAvVjAhe2IE3WudgytJbLldDrEgv9kp/NGEkZIPmb6motuzj+jFsZr0i
eNkdKqB1pIqcyIrBpOuvWTDlKm0zEePomfX8Ca8Grd1r6zh0ZXAegQG5Nc9g
xYUmnvtpzmlmbKF5Vg7iCWVJrh0uLvI+/U6MHyl+JSdQRmn3luWBUiwjtVXd
b2G4e+IQXv+AjyR0l8OeDShQZamjslpH/2crqKZnmyef2TeWMbWOyEi4FYCS
d0srV3ECwmjYrdc/rwbKGLv4BoD1bfnZl4AHmNvSzgpYWnWGT4ij8G9AuRr0
ziU5o1gH9agzKrXCvZiVkjIwN6FFexGMnXdDkX7i9D6/Ejguo4Z94msoFtMH
4JuN9chm5Trw0mFtcnAs839xsjz7ki7JtKTjihLwfu5vn8fFvTGVZrSXpcv/
SWHBoFq3ih8WMMqjr+n2yV9Kox+//XKZZLmHOtgetOxuJd9lXHr5J1lQM4e7
iOgAX11dkSthN/Zg0htVlx1ZHXG+QC8bUw4IMn04QPJ1U7tBGBMKFew+SbuG
B62CvtqPDcDgsf7JXdHcUZwnyGIfJT1aKoEW61xK6czOAHn+pDHgG8nFkyQ/
iiNdXWu07Y/DMiNztXJ/VULFt1KgPS55WY6aAj9pGX0Zam8FoGSb4hcV/Llk
Zs3WMU4wMWstXAz3E1OtkaRcofGu4gkx6myjUg27mrZ4lBoLJznmnjGQFhEl
O3losPlKzE+gJzlUF9vTtUTLZvWuIKsuV0IHqHxXXnagHKm6ROj/QgK3xxx/
SXd8o7A2zXeCrztAsrnj/c+D8skDG9IsQumM07Ykujuzq27U8JHerufDLu1r
rrYh2gbIhI2KWKhogITuFAqpa6aBLX6rPQeO56y8Mg2TN6nOZfMdOZdjzpWb
7cOjof4roqtv7R3/0phu0K5mh8lKxjoBYcda3uedfGMq9D18n8eHFyG64A5d
hETBwALO5paQ9GmWCP+oYfsmikn47TqFrWeWdigcI2F9fsw+o3oIKOULHM6G
dJAOuRL0wvpDzS9IJRHk5gqCtZ2RfB/fUtk2AmuLI0AGlWxJQoFpOhRQ5lIP
7A+HfNW/rtXEfjp1UGqdtVg4nX/bwBLt+zhQSrPPJLuXtnaLkip6sprin1fV
TFr1tDvOkQP3KZE44etOR6owuUHt0TdL0B8/vr3F+JsNaNo3forxQGmEzJfM
RjPKucmuvotvr+etPZisHQHiVwrARsZ6cWyb0ENb79mqjdZ/YkPgoYHzSt+Y
A4ObWVWbHE3xLbyRxW3XBGYLqhLeLmJAm/U07Bh+ai1iVcvor7Ctf3GKFTme
D92PmN/oIcHjv1lcXi5WZCS5exMHvYO2sCzYqLRWBSJjxTikrMaarTUHdLkZ
X6UMu0ZWVh9JWgxgUSvd4RhYgsAQIbNd6STr3OkOfqBZbKhOitIMgZYk6xM3
vv0FWe+gSt+er3FoNYSz5RINVlj5TiP2Dn4zZKsyLHMnJvuR1fTxIUXL6gIK
ksC0TX0FxfTwy2mEtUQs1BECw9x4l3rqfIonwfE51J4M6j8UuQSm8yoyMJBJ
bynTblAj7CIs6XDERDwRHPKwxtQWp0sWJjb4fzm6P4TtJ8n0Vtnj8P6iXgfR
ArASlZqrMxiLVm4SiBeN9izPdq3yw3Q48w5HaZB8bpecZTrmr+HdRZglqTr2
geUp+xSgag1mXsgNw9NP8PAzxKWJVfODuM1/QC4XXGdNka/FZ62Qw7xwaGYX
5K1nIj9LnQ+hVRl2Qbq66lD2G2Hxur5/gD92QpV8/ycOPGJRUolc7tJvbApL
E4yixiyuC7FuowbIIATcBKrImrMqtRk0K6J3bwHwPyB4BpDTvlj0JGNlBJcC
kvNdO0k2QJE423Q6tOEf9BiuAFa3yHGgHU38X0jVYXvz87jJ4kULuhhEBdp+
p13TKipV1apCxSTChVpRLX4KK2000SwoozWhrE57+SHvg6m0uaGCEOx/LctB
l+OaK/r4uD6tQxx4YpRiwhR+eqvK0OGzGbns2lTGoOg9HgbosQpDwxS48B5h
flueKWSCfH2H4LqBvyRed/I3m1ctXhWoUSo2uPFdj8iP9skfhkTQuO98f5QI
xPiBsMTTV499YqPtUW2ig5lQ1ZKvOO6b5GvGf1suwOZ2WDqyYA1s+RDDezw1
StYeqtgKfJ9TVo4D0iTLOIYmUWFIfo4jcjiU3+JRp8vfhDHcWaf9CwnRsr6G
XgKtN/DFvxO2PDvthObb1TjyFp5ISMxOQjmrmvdYDbCGy5pspbZ6y1dqNcrz
cJ8iBgSe8aT4pykn4xg1QTd3KV+Lzw2KfMiJpKvmhMzngAZfKVOp/YJ5hUd2
NQtG1DaWpvOpZrMXVqVMrtXSFFgGYf4hBPfG3Woq01eL8d1zgIVuNzK5chNV
RKPZiBPrFMAOCNjhHuz2B7oB9LGBcoPvQPF1d//17oDie4KpPIcC+9PfgXVg
KLZLSOUv3U0n+5BTbpzMPVkQ4tL/M8EXXHQULJXgxY+zbLICZfLH89doGi9J
JOPn2TG9oLkfTzvSDxomRL9Q5iYUmKhnArKciRL3MJODGHop8/Nfa5SQG2YB
dsAlgl4Sbk8wGlWB+OVQwuXe3ph9aNYFSCz29+ux/gHk3jPfUvttTbkk4oaW
1DAu+nwJsBrSYRzGUxZCPevIfX0c5rdZY+W2XIds/H6bFzKHzpBdSE4mbypn
DGBLiDAdzHelKrBSr/tMcvIC3RwRdGkOVviHJdRdd6G4GYJlHmABxorIp74w
ztBgAMs0JKwjYEw0P0uhu5JRa9pF/W+tge1By4VI2dA36zZ797hSEDukVMW1
Xyewqsu2esoE9RrjKzA8ATHCCAwMWxAVcVnXLY9k9A9x0PztWdhcmelMXjp0
qJ6xqzgJdLN5A71B1fkGy5EJCDBqO4vNqTHWfDWN0J71njKcBfCYLUI9DIaK
BpFnpAb/ucAqDw74tOu5kniFXuTQ7QrxDRN2yOiK4FLj7uY1xe6MOHuhFzcN
R3eKoF9jSGg7nFNB/7F/MK1Ihs/VF/39dP/sMmaRSCOmFoWOjxgzREJH7xPk
bK4eGcLQCJkhtbj3bBcEMA+ck5fBJx0tV9SrhHW++zxvvKMb/Hlfcp4YZUMi
y6cn2txWLw+pKO4SW7AFkZNr0iaYvgshjJ94xXdhYVYZS5gvSPfs9A/NsUgf
M56d61akNZZyvbDN8SyczoeYXhsw25mEqtRl8WShs7TBRpkT6acJSRjpunrn
O9yrdpSCiz4ADhGN6W6TrWodQVmRRhE6iD/K9GW3iwm7oc2h9SFW26he2q6G
i1FSITNL+OGcWKIcwyCFENMYyl4xjwMA0XOpusesycOq6DsFWPGl3yipCUzf
xZzqJuzhnxi4HfGnAVniql7SqE/bViBnlXHpW+EFpp7Tbk6weoSuKXsdt1ay
Fr1+xa/v1w1KgJOMdqQDbsbpBFYxgBzI+VEGMH0tJslzEqMwcFVICQgHRi1Z
J5Mu9opLi7U4CRN0yZonj8BbvCWT9aITZLCWMaobiD+TzwIOVcgTl4DIadF3
VB/Fm/bDZSPHL70Hc6o+oJ8xzQFWamBMt4lMfF1YSZbCRi6beeClvBwjtgG7
O0dUgSLmWaMyJ5VK8PFAxJC/x/jSNeW2TgB1j24Fd6488pdlKy8i3sTtFKLp
md6j/yYU62CABFz8ip/HTlV0fa/s2SCdA6AdaoD5wpsv2H98FSjTBZiR3+c/
SAgMdFEWeoo2AmaGCWPMA54aOA/jTFV2SYaAbX7WUpFl4TPoYf7P+UIDiNK4
s8hE/oD25srdiirBebGTbnemumJwwyuF0OUU8Ii0D6724F9STr+jMJpC6kR3
6lxHK7qya01FcnkOEIEu1zMmJrU0SefboPbB9ByXd6iqu/XRi9cKCTcmQQdU
T+Z2+SbV1MoppQZlpMaACgNKkgDlxzCqqWjIkHDIP/bmEM3cCJjGjnPPeY1D
XqISaRHQp4Qp2+84i0gG4+XD2j/Kz5Rt54l7dZ4BK1YDpI7q6qZnbLpaREPu
k44J3MkerbfAnnc5PywDMoUcQnBFWqu4n5ypOmRffcut/tkNQvl4KoxdxFdZ
9X3EL1Kw4ut/xhdTOXG47BObHA4Lwuj2OuM9OLyH5G6xR+GVXGb7at09i7Qq
G0uZtUtJlDUGC/uMzobfzglY8P6nqLaSjC9twKX+0pI6b+B3s2Xe6pq1f4/z
ZecY/y8yypFItSOeMk8rr4yTKh/bRZAIEgykvfhXtOasRO2gAjHg7/VBUVAr
wVxYR8WFkLWFos0+NBRW4e0QArzA49l/RxAwdcc26lQiOEGeoG88kA40zoBj
9XW1IE1gAFKZO5ccrjZvQDymtYDvN/04gVQTaJxddEb7tgcnhT9p/z7VtklP
jaZsPkJ618UsIFCwm9Wb4JGh3bElNls5Igdi0ipn3GvMEOylD2oYGVqKuMSh
DiNTbMl62kfJ5Frty+NT/FPLmxksykjQl5QM466Wzv0Xm2cU0vdZpGns3TlY
n2dMgAPyzJ3QgFKCFVtIych7k35TspjSKL7vv+T9BVhYoarDz+nfdKkZM/pw
Q5xhSnpJr4skVuyHqrmm8hJOEfFsB7+d8dsF1FCEZ3bXqXvyvZNj62dm6d2n
TkndgcORKCISrXtdgElkaxLfwKsxltkzY8I4R5B6di78mUpK8h7wdWKfLeup
IAykuwto0LORAZ8lzmIemW2lQ8nivq9EuU67aq4PQ+l07wwqId7x/bfGojZQ
OYXCJoZTRaCwNrO1G9ps4yjUgKRXchihEOJ9Olsoc+T++P462vbPj45pw/oT
TPgAAEgTlITKDy7xjgrw/aptCwVRd0KVIzsEN2blpwIYLxhL/aOnA//jsESu
rmDi713xg5MrFS4YGDug7jE45OWK9+cn/u6XDrVvnCVYau6XVrVLbcRLT3Js
kX/TsrxegVb+IpT0+Kicz2sHLkSTtD5cXtLzhot/tq+WiJqT5cWg82m9FKJ4
Otvc90swqr8TOaxuW0YP4w8D2sV2IlzMYyw8/PNrPFt1td7K8tqCKGZvbKoN
mbfD4WimxOUHT4VEgGIv+96I3CbTHkDb8YcPbg+uP7ug/QNAZphSWYrXfggX
g+6rvErCagmiu1Bvxp6xS90JNSKVzzuJ/GcYt8BG21ZHTm7HVUVIYuVld/NR
0QNqwCjfQs+WBx4Ams6m6ZFw5aHFFIsFblg1JPQGXixyxhNrPCwMrAvjY08N
3xwpE47mesBuBMZRo3s+K/KCMWFouU4yTAJp94DGeD6PimOs63KoodjngYKL
HkFKJRDlzxFttcbJynqRVssto9NupXXehsLoAIXCsz+FirxLLsKAliuaZmqd
ek4+5S1mBpOu2eGep2o3srQAnpT8RqpQGyCtMR0vi+QZIgtHnBFzrDtZaMEX
RvZJDqyEiWioJMDmmC7vRL9rOl6cVmovEjnxhqFZkITdGERdIb2h8PZhycH3
TsbulzHwGzY3goD0vCCFt4UYwAjCwTMWR/gCOZBNf1iv3r4+52tVTcFtCXfg
Hk6wFVUrHczpFRB6gjAYvbbPPcOg9e7dLThqgPx5mtWZfYvpZ0jZx/Hu5pz2
WBjLWnSAwzTqbPYClh5ghH1Z/QM4GmIt1ZoJw6GGbDgfwy0qXQqdPy827LM0
t46XRu0we2S1nKoeC2cuTzxrAr8/1/7vIU2iZA1YDvKtxqYOKvBvspmmcnKL
wbuz4L1KhZJN+HusM89zzoJcRqmGPSqN3MQlVeRRpUb3/ULVXoGakniDyXck
7TbpJ7hFdGsiVOlrE/9FZq7jlDivpmY697kocVksZdP3MpiWYeQRZRjD1z50
8z1veORJEToOZrdWke1L+xYCiBq9viKjf4g4FkI54SvRcjW2y6jUEVeNtQO7
jVIF2md8zHdLaVMzZWOLGFgOHfxogIIYtakGcxmXIKCSrwZtxDFOvXgJxhQS
/i9xqRGYHVJ/HvR5Evt907f20e+TrvGr6pyqEv7KULXQosAsfCzUOnRhggOh
M8MIwa6PrXNGtxx/OxSnBpb/po5qDV9+B9fGDd3TmjbdsP4Q68z+iz55f+u5
1r5w4Jb8Jl7Uamvux5nKLQwd95v8kC/3q0oYE1AsV4rtiptOcG6TWWvDYGFo
T/o5wFc+5xw8UPb9SI8ZqUBrbCGalBG5cq8xXjs0Z1lSGHJ7J8NWvUN8gn4A
/HScNJcCerHTIhrjM1H1OD41NKnKjxfTjHlBfaVOLlMyoO07FLNLcbp8F0eq
HzvchO989AQyKqB3Wn4cxP1LnF2rLkXLnXKX95xQwGvptiU+2Is2EmosChAh
keMpX8eX0hzhJM61KIRztAycon1yYCrM5OWyY84KUFT1kDT2wvBUpKedWHp7
SpnnnFVJbKVFjZuiIrWZNxlALQFKmEpw8X2dJV305SEtLG5D7SSObEbjtTSF
rkuF5BnKlrHqND4xwzFKaX/PkwmKc/2UydSFg7QHN9Cdx8qr/T3/MqdOzI0h
9On73wy7/PG9e8JSkaecVum7JhD8y6kCfv2fm7CwGVrPudV+9kJ14gCLb2T/
NJXArOBqUD+dtKKAzSrk4LJsHoi+n0CYx4Q639cX423P4LvkkqVO7DvrqeeE
YfSk9fBCOFzX3J1sEugR3Kagk/37AZQxJYmHmL4U9itvIHrHLYx/MB2XmeFr
TrRCFg5wymtQqxKO4mhHykE+JgTTu8mSSRwRtV6il1k7AsPDrWq5Zxusd0Dx
jdAWvr7mi34tUqW8a6dYqkWapwA8lOKyz1D2s+/RbYrhQmbM6pE/XraVmr3L
1pmzNxCDu9nj+3+qyyWH2Ll4yJTO1qj+V3vnYyUp67F5Y+VohXm/pduux394
C6aMzBs8O7vpS1Z+u4UVj6KaFIIYINpA5nNNm/tmTldBzAMRAlIFhKtUVOg4
RhH8V6/VaQf7o2IMHh4eCjYy/dXL4FWLBUvOM7lwGCL0vG5XLmw1lbscZ8G0
4sXnt1zPHVBvD2+UEPI3/NCAPW2Pa7QMiUimgsWnbTqSWU37+GBk4LEVdjCU
eDa7BkC6Q5nzziMEXwhrxAhRhrnpPza/BS800allX3WfayeIK64G8iDpW9id
e/bu33OvpNgsDgBE+RvY+1m7UkYc9XNRJaVXaCfWEuz3WLsATcti41i55aUJ
5dMAe2zgWLzrlqOorjXrGC/GdLgXYFYyOTbJLCjRHN64eXrsHnkTH6qEw3ze
hdNkkJ9lTYzez8giXCp47tmmoq/Zp0ilRXqCLLwSzgSmjPFOe+LILAQ7Vm16
qS3a6dicVR23OGVQx8jJxBa0MgJkEBAMPsBqdP6sE14xhI6NNw1ZrqLlGGmZ
LcqjhUMj2a27BHcICr5d9DFZAqOjt9gTzyD7nIArS4wk7roCgIdKu9zRCpxm
j/2tQnMTurmrNnQX1epHIIYl+sQ9dUgJb5EA9ER1JuEYLNnyhVuzX4KeDRXn
3yQYXNx8l+K0yefxDSaSlirYmhxiq5D0EoxAsop48rhv/SihN/cZ6/n0bj8X
nNjmbzU/c4VqsGQFLV7vnYyUsGbZS2cxV1Z6no4dRAifnmnLiiHsK3FPUB49
yaieTXBXdUDrmhi/1RK7mmS0nBCBxm7EvBiJKTnMOu5Yh3DGAHRk+/iRxvLn
j6C91WC1K0P8kWvvoc3RAtJ+oFpL5+hUXw4q4gwjUj/3/0/m+QfJ7cDsOLRx
ZBrwcBRfBLydYYjXMuKLiv+iLWuC+hHxL1JSpHN3AymWCyhQA1tgHvUmxJfV
AiqAPyfIc1V+poBmBPTM1uj7ahMSAVbyqa/9u871W0YB6e9I01LrcwPkniol
U51KQeFkTzLh+8nVhL+bPHO9RxAs74oPhZ6gAMWjvV1opPmuX4sKS6ePduQb
YWPA94XL/L2HIDcMj2W0h1MhcRJXtErPyTYhjveirL7J0+lAnpYXhXfjlKWi
cLZnxs2B4rpVRiSv7fU0G3zx09ol5bHLgrAxOcSUymd550BjwoXxjxILH1ZP
yhd28YlI8Wm+9ivAsksgUUPkRvyFsMvUifpikw2GXOzRmMAz0AMlFgZLgBCL
lwOhUNtpPWWvuEPlJ6H2dOqznIyuoD3tmuoTKYsPVRT4sHU1giBGtVgPaWeK
+0gGZndCsT+yMHZTeO6lBVbyDmLVespEui2mLW45C/t24bMh+soFei+VPmen
7vQvx/fPaYL9CsH9szQVRR0+LxAtbcxIenTV8tbXNUjNRx2nM0QNGSIn7AQw
K+hrAcTHm2NLYqLVUvKXC+EVEv4oMRhxZM6vGi3ddj21wIqngKF0qmt9CMJc
csX5nv3C3hkLh/W1hi9jXEtaZ1Er1bFHTlQaLIFXRMWSR1y0XREu2AMxPf3c
UieX0gVjiytzi9RWcty+ysPNBI5bRLPQ4ftzWXSA7RGqi8i6KO+24BtPb1G5
v/H8Q+uvzf51KVikZFDsI7wiLjzuWcQ72/8Tq9w4VR2l7cYgpx9m3sE9rNFG
rubjJW7aGYcasqEbfEpmkQYoOKfXDRKYV23yYtw0kdo0GmVaTZyMiFNlFii3
8CrPbtQtpXV40KTxTV2d58DQ94wdQLgXH6lg9pV9qY34asvcBZmQlzoHWsj3
Y0RshN+F9oNSoxMiwxj+2VsmaQDMaq64hhG3henq22ThHsWRdl6jALZRzFWu
VWQIyqkxdc+vvuq9CYaOPt/Aydkdpne4irPZp/PL9MRJj7wAfDq/RyC+jb1B
Ti7wU/h6JS/0iv+8ZFzzgUr7IOlnflQ/Qr7lKkLn88INjX3ZTjmJcVByD6AV
IiMuipAXyeMX/PMXQNZNDXBuHiKdXhiqbzoHddK/dnoVQdR51iewsQqJnB1Y
+lbfNGqZR2PK3ZWawfdtNP9N7tsG0NASGfDEPkx4YMyJQNRpymOGPYVvb5n5
HmYdm+mgLvNr9y4R5imwERNM7KzxNW96YiqtRSWeamD/NQ78FQPeWoCpZ2Rm
VNz70R6Xbmziy0OY+TgnGjtU7oiuCw3QSgEkw9MRXvfbp+PqIR5uLMhIC7Xs
yJplJ+5+tNpmW4IYs4WSiCqIRz72IblKsCIsh/MtqoF3ej44jqpR92D31MeY
RhslmpzkDWU1+DtzXaW8LwuJ4VVi8AWrDqpZYdUZSh381nUYbKEYIGrRV3So
ym8MIAVu8liayv/FfMcA4Ag1rOxSwnM0uGjRJMazqScEeOg4ZLt23z0YH3L4
R/pQHqmbyDz2iVsTAlVAxpTUaahVznD+FDClQwdkuv8lMxrhfSc8uq221ZiW
atPhqRwHnZtiq+lbQ37YhWbR3fz8DA4Ug0XIPCgN7XZOtY4eXSpTsd3AOThD
QWI4SltmnBTSSlO5IRLTRZ3HAvRXDAXlpvI1oluKDpVkzzBQXgT9TInBknJJ
YztnCRdbCTtwOfvHizTzTIFWqJIzas3zM9BU128yc0qCrve5BfyEflyr/X/+
N7li6B6ZJzqp7u/ZWrnNgl/6DL7WrgWRDZyvuzGkOeM9BlDONZc6UPD4NAEg
Ng7T4mMHvbxN8xaw16SRvjHjUIUq5RXCJ508mRmtMITiPnrs6C5JsC4loor+
5nAGinrSHJO0YXhIuy0rWS3ehQ9lhkzJUy5r5abKs2snIku0EpqJ2SdK5Z45
OEWLYq/gtDUhUsouFz1ohZXrWlIJfQ+DG3zFWPTiDi1JcWIThSjn3vgRreAA
FG3UoqSePrZA6TBTAluhiQBMqwFo38dg3+bUQ1B1r02uAQGjWjs7G6NewtMb
Fsx+/mJils+VR1x0fAQhJlnhwv9PmtchAGCYXfjjckd9tydMMW0rddLdC6lw
vcLRQ9IRHFEtfJKtpTEtnqPO/7cqmpUfL76vN7lOSJXZ7KMz8fKIgvgLrE2E
SJvKne7zfJ0NIGf7CNKXSwx11S7IHiy2l2qE9jhrUczoEc10n9LGC8mhcSLt
4MixGWdqhqgUWNBOQzFyOtWDFsPB0aStIJXBPq7/nb9cDgd5e+4YBeoFZpZC
k2lZtpYBWGyhQOlU107U8m634JZ+qfXmyjtYMuPrF7UZC+/Hqpk0nqEdG8sW
iXUeN8q0OMvyw20lszdcDXHZpE50AFqNFV1RyPFn1FJjiLWVMrAF6DSP0EAM
rNM+S+jcOa+F3hb8RSml139DRdMGhIF8xAmk+h+37pFNiHSUvnI8TkfbibcM
/G3x9/6cShABaXBx2rahXDBjBmWCge4VGHChtSNLjSuhRcjt39XAnKOaMJh7
NagK5sESXOk+E44V8uR4aVwjZF2FaOHwh1DAUYuVk/p5GhNPW23ykPlgAndq
8CJqUrAvFOi4mpwmseHKZuzmhvUY23OdO8Asnb5FCpZk8WOEPVU5WT7ftKqV
Pnpudkz6YVCR9MmlSQRfmKaZaV2++q4fsrvOso3NIOHAjfacjNSAZcVktoSB
WQXMjw5u/IKNSLMXHgbPu+d71+1GUinQZBnN3KHcoxaRntRbYDlENfN849la
2fmXo/ue08Wq364OfeNw3uXrT7wilR70Kj9NwR4wDwSkZiWRgR0mbUQ9o994
JPsMXBPNRyND+39vA67CzPTCB8ptB9bFdVf9BH5+k9yV8UyF9WfhXFhJRwI8
Mc9IUD2vcPhlNClJf6I7r1HsSCOchl/9OFdOt4etzBALHs3H5JOV6G0jdMNQ
Eojk6ifGUyCWDm7TvuhP19Vb/ppcuIeYH6ZLk8apcs7escxOBWEG+rNCKLrl
/oI/lsUjvUjqj6GD2k3ko//qqbClJ82KU+xL+S/wgweB1sXVCimDjDIpZEtt
g6LtAlf3LU6GuTQiw/kKJxicIUenZaiAYqDbiADI8Ywm05G4iZvrafz3vkxL
8DfYBbemILGKla7kKO1A/bUxKlSzsexb5He1OreIBgQ4jsNTmkMnAGCWt9ob
BT7Y63BqX/D0396n2IDfvnkgHHK8ITAvWQp9zFkqHXS+RJCsaw0lbtUOwWMx
pElnYVhtVGyIi2pNCOK45PUXdnSigzhVx/PCkSkSM6uwu/RchwwiS7pKobBy
3G8HqYD1Oxf77giTsADV4Hq8x1g6LAHGOqDUJrYXDAf/tN+++AigwzsdzE1t
5hiGFAwzqqGVPVCH0d5l6pqdXy2CDio6LnuYZaQ30GJeUrimNT6Mvk6qwSkI
lyY8rhp8Tdm1Gz4YENHBUikp4pxeZ6N/FnPQ+c0K9li/SWyjSwFTnYkbo7KU
1axmh7WN48+1zognRD5t+k3HXevSGvJOx9eOX7esyox7B3PxUdiJMPxzdgw2
IH6nuAlbeO60P3krqKD3jISzcKLwC+zM3zfPhLQRLmNFVcGhGzthOtESTNQ5
ftTus7UXR3Xj7exPj5WuasWdez6v/q7Wki6Ct0x4eMlLV3es+bepQNDYnAWp
TzAaf/PnyEXhdiLKqCnHjex/vrlnQ79JazjITPktIvuugIRarILqS3bKF0l8
tAnyePjMaMNUnX/ysDdvbvYNHPiL8r598YrzKrMlbNjKXhekxlCZD2cAsieu
4KxLHdu85hlXHj+fWOEYU5yt/VYfJK0r8J1TPPUZkTrjn7GfJ6a4IShRhaF7
JhHqPAEgSVslmYq4xhfcOtgj2I5c+0UZhU8a7AYWceyGC4EnNpYjlf6dItLb
EMRHHuObFS0Df+/ca23KbGHZwJcg5iJLLOWX79j4T736k3R8ibFeid8RZqlD
vpnKPyo7z65FLr2Afk3volkZ4NSSVcK3ZINOr6NcEXQE/NZOv5ebA6DeSHc6
AzFPw7jDOJ3lJDNmk8VqK1o8Fi8UrwIC3bt0PWhrw6hPHhA0fR+ruakVR/1+
JCnPh+uBUI9WKbjpVDsMdvD4me+zz1550xNyFC9qAxPI/mrUGEiEc0w94Eub
TWcjM3QBy4UGzZRCecJNvIglQfJHm99j7bgLz+8IBJkKnFQKe7aMHXpePB/j
CvmwSKw+hY0b+iwtWWhPuV/z8zcr0xuk3upS+A4inIrFs68+utTweRZ7ZW3E
2TTrIgdXgt6M8h8fWZN8dxCUI+w1iyzuV03GY0oqzMsIbaNPMrw9wfGcxiT+
aHSpaWWwYnIsUwyIx7BHi5l9Nd6rWuWUrgZPBJk599c7S7EXb/RUCWHeN6yt
HjSiEuGz3bn1I/IduTXkjiRggj9DrFAohtec8hQ2A8wUw579KGTqNeqNl+iQ
VooZ++Lb91+FfAZbPhAvBkY0C54a3qMilXqd4XnZMmOrcaTCxskUSIuMYSSx
iYIhCP58A95KQ9ALuAH4WPIcTqobF2tJ9LYU00ZBvP8UOh9C95q9QuX33yve
uVaqNeJeYG3i6rVdPcCb+9z7X/bpf3EiMzmRbKFly6X9pAetTBiVm+4/IYte
n81cD51uv4pp+cmdKAvIbwolpUx+uuWFtwqoEmv5TvW/seud4R4kNj1pOS9h
BZqBhQqo8n8Wm6BKdKiH/mqR0NPMDN7ThJt0NtJwET9IhPNBIWJPFbRo3fVk
2dFikGCMxh1vq8kFqw2nrm5HQASLo6vO6YBRgRPL003u/97YEpv3mfaNxrvi
BeWg/QDFYWD288iB2pZlip2TjLdHDvzOcgoJVQpDgQisnDrUbqHR5kbSsbbq
h1bRbsi1cMVBnk1me5nq9eb2fS6b0d5QHiiJIpWkc4wSIP7EWEVjGtY+oc1H
D7UzZeFDx1FEQLebVmT/jsWc0cCeDdWNLUKgOxhf/99jmxB+pdKCDmZVVmqF
98NGixgocpGioe+D05qw585uCrtd+DM73OBPy+yDGX+drDqOQl98VVcGUeFZ
J/OZGk2z7HdLgaLVT8KWqdDj6L5+i6HEcoHL8v9rQRR/uUjpWIGzqMXtG876
p4Wc3jw5Kc6oqq0m/PmeHBXw4oql7fQORWdQbgXHVOAMmEmJWEvE+C81Ex17
GEE261L9XQsckNjIHGnu+hv7kpZ8AoudcWRm6o5vpUwC7bY5VkbaDjZDoWzO
NaDUFHQ1AwX01AdanrjVPQxtC6zvt8Lw5VRv/NPDjGqxaXtHi7zYYHUxAFQL
dgcrHWG8vm6VLgyMG4zCSE/blDab/q1xzmqrSXoHqlhL6ABg27rv2HcdHWe1
PTRELgGQk8b055XS/VI1faxfV+1xkhVYk6x8ISVvZkzK4NRFN4rLW8gcpmrT
ek1IicKSY3tZmfHGwRFqsQZR4IRiGvkBrA1umbhgvSxH4HbZmlyE2b77kPtz
4jBMm+7Y9DEFheopWxt4MoIiK9Fbaeh2Fst/21aLfSRxaFxdM3bQJ8Lj/m3v
bx+vcGEtfxVlfG61ggP9FpyFQ7O6QrF7wla2F2sLky6d3fEqbPvchmEHtoyi
Mwa4whID9/Ze4q5FfurJBjbq4ihvW8f11hVXIoPiCYetjWxzabxZGnzKYFpf
p8kQE8+S0qlRuUDt5YNRMGV4llQX2nXc7MkYjWVP1Zq+CmzpZp6yCPRQXwyo
jXtQQmIBuQXfUh3V/bFI5fAwxcNIcyDkO0rJQbVgB8RfhTAYcexxBp5mOpd7
ze5FeSePn7DiKZGInK/r31Gpj0n4qmTGhKhDW8/FmFJK8ve+n/PxNfG5zDXn
TtzXd6zkb5H2MvqVS7E0hTDtne2nTHRD9vLz36ob+EaaSIMHmnm2k+ClQahW
Hh7sgHoT2z+YjrmEyD3QhBYmtdujPydAgqlTPWl+S4C7ovmuWlK4673djNYf
xkDjnhtpRsfXjTCQzU4gXobAjFVaDTMbNWvPdZSBEsJstX4LCzGT5dPF3mTH
pptibadxx9SDteVt7/1/wtUoEqlajL9MFcHn+Wkd/5ZH1PlJhLEKtkZA+aQv
2iu3IW336bqfjnluX4jmHtFgP5IV3rndxA1l2CmDaQVxD0lUXxyGhTsJnwPj
yiOxX57Bc5v4oN+rk76UffoqjR3MQ043YGTHE9CgT6sOPpsgcrZFQf2Dulaz
CHVOgxKi70aeYyL77W313ImbUKMZma8Crz6MSJBrwE+BwXOwaKBLGz0yjA9M
XMwZW9Q3bIIu7gi2PmThybZBsHcIMa5xf/13B2YensVjQBop07g4gR9gJTCh
uLAqBwkTu0r90MrXNkNPiW0LORS15qQ0IEeJxe31q4zy/+nelEgPkG9QI0pP
Owe3C6MaSmnhJWEjoPl+NoBJ3xim0sIqMFTvgsmdHRtTZIQTu6ua39PF/4Ef
9lYLkL/TQam3PbJqHwHVK9BwXgn/PhjvpCPIZxQCDmFaVY8UbrTMnHVyDiT2
rYPij3buSd3kSSxLZWZafQA45km15HIAMtptYH6VF7bY3UWF8ewKr//apXFn
xZwW9lY2J4zJBH6/DK81OZDTS9d9njq7jbxhQpdnSTo8AnpucVObpUFi3NLo
Sxog6XLtWkVenTtDFrT4hrdv9Ze2ge804rr1vNoYfYajLbLRJR0Q+fuQ45/q
e3msB6Mll7jfCB2L+yA33n61zN34pF63Z6ovuIT95kGlPPhHdo0F0gqr3Baf
6Y1DL3klybxF0pjHaAStl5MJ2IUXfNtZ766+iggMbHGwCbldRYWX/LiFla0O
VecqrJTMMaogLxGHe1gh4llqnUvRQ4SCFgvVTYNp/FoGHorU7rXKyliZWBNh
QlEbtIFuXbIxGfLluG3ux99DKtnwf9HG8/YbU5V6K7an7BV3B8ng3JkUm2By
Rf/AkUaYgdrwfrOc5zWdq6hdqWrEnjJrtal7lmVbkfdiZO1S0Ju/Nyw8Fu1y
mBnl+NOs327hoYxVdovxjtiFMd80hrTJ8DtZTZ37PeRTexDuvR5pQ2CnZLf+
L0w1nioAxOkTe7RjBNDKuytEieVLNCcCdLSEZngqghkWLqfMWlzcw1zDJRON
KoU6TAuAE3pl6QMIJm3LPQO7E6M5D1tKvbMyhUIVf4SSBWjVVBkrg/T8X/ll
avnSyvcoOBvA+BybTJjRiFD3d1lOMgJDJwvrvOJqvFks0q1rnbdKASUXYXE+
y4e0n7yXcnEkphv+VuqPpJneCLHF15K6gXaYiNa3ikBaYXczdxlS5f2VxXw8
Di5vphhlH6qyL8jkNX+9olBaIA8cQR/AIY1eEMSLUyNb5/JslK9Y0yVNbR5T
X0lgbkpmNsYx2dFncKljGIMcGuadU5d92Z+vN7L3Cm9l6CeyerZ4T3vVQL8d
g6aztYLi77GDmOeFqsPVSbvxop49aleZo8lJu9o2+WSMQYvHkshP+ZztYh3j
jRqPyU3mrV7+mbRpp9qKDqxKQZyfxwKXJUbjhHe9xG/RtpyArMv1vTpx452z
q6BXKi2bJZscKZF5PNCROtS8dQb1ea6iZIyrL57uHmCO7juA06Cjv+01Q66U
BemWvHspbXfC13NggYKssXy1ad3bIrIKajmHKZaVKpiFFlQe8EDXUERCBzcb
LypgRlbEMXMjJDh/ivaK5gsb4/wUVi1ULtPbiggfUNZpED/POAUuxdlrRJCG
F2PSAavUXu+V1XY3nUlP/k4o1O15tMs73F7KP39SofzftnNaHbD/9AH2vC7Y
DNoo0FdVdbULHVtmqLteQS1d0xpqZo2zrRtiqwQC25IrLBCHlpSKSp6hw2LW
gYLWhTkLg2Gs+1fBcPUjL3llbZSLLvCic+aZeNr3Wo52AUKg49NqnN7olNyv
2bUDNzYnusZvm3B5ndC3gJUzxC5jvvwOHC45h1+wxqXjzfEDvIRoOEaS6fbI
Ciy9i7S7ivstCYdh9V1dpOD+yXHiqaHzXtTnb/S8rFJROYiNlVqeanR1KWe1
BixpRRJUCAaWYyFUU/JuuSjc4ok8I16hoxi9S+iLPwdFH+YoCLFNlJ1T4a0D
BlOqR5wMSyhQZEKoXUHOkrvAu4a7ururQ8sgNVpqrnqQpzZBySidGgQBaZA+
G4ids0SGEPkzgJ00waghVC3Gfl+GOCKdfNt6GrOlEgyD9btx/QfvjbDjA44v
/RrIDlb2omxTNMStZ1H5OeR006oPzhoQh1L6g1s1tJU9y7jhy82C+quSb7qG
r1xbCaXeXGdW9ynvjx3w57OTpReFO5vk7hRTHrIozghA5llDMzR6Wo4dxAR3
zvO5d1e/tjo0q2YkhuY49U3VzQhn+JSIEBTpfDR3xJ523t+icuOEffMaGim4
FdbNMYh0zOv/wNTQ5oa+5J43dImAwrk2vNi0lrIqsY5UcsJLPAmjSF2XM4Vk
Vby69V66AeHyBs421zSN3txN7GvOn65X5krdzBF1T+Y0VH6myMYRr50nlrSG
SePNJ240A8NLXIOMSu6jhvVLpC676Db2+mAZXa0OXhJvfFYgnFo7T4jp00rn
r66v28QxD3PUiuHuyoO3G+EBfT5mpfXfOMSKQ8yusQoKLHooSrV2NGlRe645
YZc/5t4brUTPpdwe7bw93f6VIPQNJElv+XNWMlv7Ns0xbhMZXJ/T7wLcif+x
OjNOmoLsE2kia69BlLAe7wiABI/wOEABMN45+R+k2GewYl42Oipa9xXsktu2
3mqwFWIdy15k5P2g6Bkw+7rJJFCSJLeNwJTSdB86OfQeImnN03l0BDif3lU4
oVsYievoEzmQaYrdESD+/0+5N5Q1ZFlTWbIdc7c+BiFcYrdOaij2d5+P32h8
s+fEGL3yvq97MDzSlg7Tg+OnbUwB3tq9PGk4gol049+i5mel4nIXfVhE4BWp
0bEQKJSIYNJvQYICSU6K7xDWNd6st03Gzd7G2QSjqWM9j5BjdwXwyUbz6tsI
IoPbKjcrhNom/h0S0YPtt6TSgSpCpheqTizBDQFEW95XuGFmtdhhdGs87bZa
RAhXJ3/EPHYTtYpKYMaPlP25yBk+bAtdEwZR8pVQ8/KwKnJtQerXRAAEnpwg
+5wLv8J511IwS6QDWCLVS+SMcBDLGETbXUX1GaX1Ta/xrhV8MneIFL/9bSSy
i+mH1vBmtnSAyYSw1kzoaxkDeTeKhVzT1GApTZQSNlFkSB/vZvbfOgvfGFqq
XoaenLGTG4MdSe1w2MqM3b8hYrMSGcuwXJOG/0xYVhoLklKQk0mqBowJiwB0
AxKRvpEQpTQPpQTCWYMX489yCPezhQJ1BPVwEqVuhvCoK5oFMcjLT7IVVY2B
sCnixf4nMa3TA9s1lSkexjjvBZBRgJ/6SQ7BxI/HKsd38nuwY8x8vx7hRfGE
oEePPih6OhinWoKDPmskujRWkK6+kjkZREVDJcICj6SVL+nLM6xh7czrB8SC
a377fVS4Obpks7kiiML4I9Y/1xtakgYkYluw+r5cDErgwTjuexqDwjUj5sJx
Ut5nMkNR71f7eSOOMgvhP8rTkDPkopPO3OaQIeCuS638tXVEEmTfr8K01fqW
7hMEgqqBD9T0WivZXiW+Hzzg5sYqAgcm9B7j+aIxugmEa8sCxOsj/T4ylNck
i6vibnTYZiR4aCeJr76/rTRgYntIX1ZG/Yq4x69zdh6OFIfdGRojEJddAHQB
DHwJ2n8xzWhJuldrTqbJLgmiHLhRG/IPOhtdmHOe2aDCNVYwph14LvM+jyA+
LCx7BQlhSH6S7TDxYeW0xZ8LnYtK9E/Zp5a0fSjQ2rgQaHXUriqb4BWt9wOn
TEDRct80i9qeMnceXMdBj9bryLe6pdPEgn5fNUZuevtoM52At60ttf1pzShX
xrt8QOxYUVxgJ76jJuD/VrehR+kIOgE5aEgOz2hon3F7rPsadbZzMtSwb/ni
YWhpV+wDhTvudmTAYnC8ZMQA1LnZ018PSiuWf1qh5sXC6fyC46mW4bawDX39
KSw97tZcEyA+yRNlTnZyvdmNFbbkBhE8kgAsA6+T+qGXHmMl1BMr+6GqddGv
cGTgn33mDaQ+OUKpXRxCiSyoUt5ppS4TSB05M0HjudOR21saeAf+SCwgqsIq
a5alZIa/UTkZYKIMZmIBUiS8wdE2/tjIKbWOB07hV+j/bD4GtcmWRVcOqXNS
RLOI+hoQZUoeUQHFk8CnB4irS0uvQ4SJ4KKkClDlBejNaKe9LwyOFOMnWnCF
osPErFFTB+L3gcmqYfU6p20YldGKqA8cBgHNyeytjmvZqKfijF3hToyg0xYc
4szH9CuxyiBcYIl7GAxisOinHBNXM/93MjMsd6SsEZzpSB2JOkvHJQrSGHBN
RAMI473r7ZlLwsyGmqjD4ZczGDpH4GdnSd+NMd49TCRYgnezhhIDqnDtmEjI
46pgy1SytQsnIgBCPOtf/ZBwdM/lsiN88/f2kXCTKrvjw81V09jq23VS5/j8
Y5pQruDaLBE4VIIj8NRZ7vvezTiFzCFJdoJFzlGlSK5ZAavufqbmpD4WB2NM
AT3EgqvbYG8+qynEo3HN69+I9Qu6prs0sol1DV1YFmDrU/PNuaOiuoTi8TeK
KUfOzzbvKoOg8buUMmLZrl7v2XZ3M8RliuOO86Na+iWtg25DtqRm2l1NpevZ
5pFCM+b5ijCtQIQEUx5kXMTcN93vEDiS8Ree2CTNrwhegrYJueTeuDZApkSJ
Jo8xv8BVAEh0KUbyDd+LjGiNX93PSi3akvKpuAYQlbPxGx3baS+eOle5Lzbh
4Yx+myax8vSCXI6yvlSNnJa/SnzpholJk6zYu+O0w1yaPbtgwQuol48YxZtL
c9xxy4nvcgUh3jCeAZl483+Wfjhr1xEaXnvdjTJbAHxTlgJwgFgMk5Qz0rVV
Y4FKJ3YUamTG7UcZP8z0LXptzfbtAizN8CAm4uFtt+LcRF1WN8tt8moSNrpW
8n8525aulFkij2a7Ta//3l90QVWt61UE9kfq/xmYJGKlx5XScMcadwLvt58L
kEpn0sPiFeuUvuVZoHWLjYd9i38iva5gLTiTym1mhzl/g4XDWHntAyN0qomK
q04+pHZxh/4d7h71Hmjn+3ROUxo1/3b7MfDPn+WMK9hLQJcSJoberbj2uapP
86HLsW534GqICud1q42wGXfbajd+7pGtuFng8KK5VZwH3OCr0pylrlWxZgSd
6vIJCmwJYglzWOxE5J62A+g32KtQ1d/HOTacobI1Ci5u3CQqCc49on2A2+4H
chqiL7TMt1Dr+CI7taiq4mdYi4+MTaX4XrX+zlKy/o55a9KT8mXxc9Uk2nHv
uzhqwTuBNXKG70fqTM36A1qdFAfKdfhn8SpYzvLaRzVwtQgs6mk4jHYa4ti2
7af20gfjICqcmQVcJxjcisLT1goAPAj4q15X0eObOLe+/0sIQ+0bae4DfytM
N/G7xS9lbgm2Qxd2iMxpkU05ESNgu4REM8S2tN6gRemUtWSFHzCLiu5h824z
tW+IbYrKTgJanhoKI2Fp2iNsqWTUyTnITsYVkkhoBEpdCTQWv6whB4Cy9cgO
FeXWr5kLnUjztTOEBRe+4N+z3G+S6l5I5lEV7rjnQsExQPSugHuuWXIzpg0W
Ce+fQLPrUYeSedpdzA4EVWaV5HWqgxGjwSzzSHLl+/rjOq+Nd2tQ6U0HIUFE
PwDCeGSfj2H+zpQdYyeN/zSw4g7gWpYtDZrVS6lxwI+REsPhX4ttZELLzuIK
8nyxPFncZKJrStsbhNX0jMY96/w2wwoF/CzzTNOyZbLO69oHcX72H3XdxX7N
qB6kpXpwd8NCgv1ZuIVrHR5/ZDwayVTqSduRCK4tmBGK5RDCXh+e/KLv/sWI
3enTdzYGteAqS/BeLlNe5VerUxd/oovBdKJrRMJ2LXS7iROBXRWiFfkbCyhr
QLuMTB6dEgphkGCUAJjX/vC+ntV0ZQxa7Wqm98vR7yWAKM21yfyW2lgyibfS
xW8Oh0SLL3g0gaO5zA6r8ma5S2syEhLFeJCYl9uOnhv86zf5TtVk9jHy9yEk
jGKBBre23ZPnX5zXIB6hEk1c/h/6ss0rVfGr7Aae9C1FpgtTj+f9NJNVdtM2
+EFIX6muhir4Tmim36/4riX+ZGwp35GTb6DktvpI+pMJcOQgnHevgpbDYeAj
BXkAt6FkaUF1gwvW7RGu//fG1yWExzYTombQBf3RshERtI6YFstFdqAQ0/hE
p7JiIx9FmPzuckkIZ1LIy9HMMTDbEtp+7rxSxdURH+bDtWat7oxc2XFWlfRP
eZGHHJ5e/fwW6XjW7dZbNci3WFzgI8Ha8Mn+Z1m46o9BozcsnIFVFd9YDB6W
jUJvvRC0tBoP1K8mGzOJUf454jErDf/r1VzXh9zNBD3/ED1AOOhzEg0GGyY/
aXjo+MXETJkKiu7ufEGG9LoF0fVtkqkLsAofqXrkJ74mEsTYFN/6QMfLnsN0
booDvlEdgNgNPISt7+RolRt+ODjhq/yX6tMw68CyS0cV4hlr1pOFx3iDTXgI
KKXy5PJ2GDHypDtlfmSgHWZt8PcRmzsjOsNDq8XAovibs3FN09cEl1vFepj+
ya+chLVEdHtjLdm81BhlAKcQFfVQsjaUh36B5JWncIPcEaLYVD50asRiCRSA
zOnnDT7+0vjpeeFGyhXLj6gK/wbH36xpeub0+FfUSiqm44zfTGcj36gDoMaX
9MYffd6ayJyI84mxzoQH+xwmSN4zf4tkNNG+oAqQw7BxB6dnQA/SNp+/9ZtW
W1g/FnT14yJur2e746GxCi0XKDG2aaeI5t8OnngrYAdCJYrfXifT0UiPYDHA
vwoWgx1iawBp2+BdXrlMANTvttPYtHwZlTB5jT9uivncgvzEZa76+sG4bzmA
jZbP/BF2FgHw1Odoy44On1y05tAUkn93BADOi3yjL3Wolrltgetm6I9hLrut
yxs5WGBhZcPCpp2aEGmG0jMF/n3IbtVPOPhfNK+xchBSvyJplMRptZ8ZVFZb
V1hLyTK3ZAQ5RAZVRA+QlPX5meVXdvB5hM83mfBY1sdMAFKoy8gIT5yiXFp1
bbqCxHxwz5pDClGKU27Kgpci9hZ5m6szbelEtKmYruZP1tKK/ivllkHqw3Q/
x9Vti0eiNcBnxatclYFhMV8EbgrfFyK6eFPcQXX8iPojeL7NoCIeGJRT7tPC
QOEo0Ljs1ZIOa6hHje/UjX5jp/r/JhEUuwmZTCBUydhIo2KIr+oHOfX2ur8Z
CN4nlAyVbIUbLI95iHnm/+Y+a67Frgf1QFRQ7FwIuW/CpwlCly2XbEojgHV6
BHwwtSTluGyqxz5sMyq6sd3ph+VavIiSoxfPQDTnlcNVy5yc9QOSAZ0DAqEg
OuJ75tc3c7MRRCowikaWBjyvW7cq7oEZlKxUoo51c7H/Ijjfup463QruKTyK
EynVGlIFgjNCmJBrZXyPBcWq46jlYi7f2VmDPABtRa8ZgDDQw3FAzq0WvdBD
kwBXzUw4tqL4QDZppy8i3Liek0RAAllA//JTVvjVXURWswNEbVfqFW+Dv9uW
MyIC7ITYeugoV+iUfgIQ4Vz6DleuBJuT4PEyXSmSWuQMUHAOJTpJLSOWpDVm
Ei/UoeGlLnA8oNYa9SdZNVyusGOmhyunXCySGDxrj+YtYlgSM5ao3eBat2U+
TmLneuonE5YB2IfU4uTR5dBv/9LQITIkzi6Ks4zUoYnnCu8KxnFLtvRu54Ai
p3ilN/z4U7CoySt/5NUHVHP5aQ33A8gffdN/N466GFYzx1Bg0qY35vfooGnv
7buy3Jz6DVjQAEyTpWZuB+ndKtGbB7IenbamgxgychMlXPQZvRvWxggqo7vQ
PaMlLOzCdZvQJZV6I7psCduyA0bR7UDuWaRCWMZDsJjDF1VlA746+P2DA7Lm
qmydOc58eRc9gcg30TixaShxPO57Bw3i1mVJ0acg3l8POQRCeNq7iCtjyQ0x
mXQbOl6bnRSs6sPFVNyC9NXtH5dSoNIaVLl9ty1sSQw05fSVbyR3Mo2aTqTc
w+A//bKTCD4nPlKJYZJEqacI6pWO+m2aVlUrx726UgSTc7zsWaF731FtxawV
zeRSWyPb2ggbMsHjg1dcvSLRWCFtpFer1ulrtdmMKcJHp31P2OqxJRhCCVer
r6qEKbFuTOP+RthO6juVpyJUznmPy/4sj+R5i6PnTvzYG9XzsLjchaNq0WwG
3KvImSikU/SXiMgMNFOJoVutVx5RYqCPVlEBbCBYG+va+01Jx8+siAgEW17S
En7XvHCvNSGAp1BQNBwH2fpCz+1eqjXe6mkcTYF8R70zQQyVFIYixgIMdZVx
x79wlrYF5mpb2vrbU+9Nzm/xSyf/Qx+gCrCtVNayOBDcxGs5wTDQ82v2yTig
HvaRZLOh0/R5tOuVunQo16IVjgGjCkLgzrkjPcVDmEYn+sql5bUcOo1LkJ0S
OqeEStBTdtQpsjb/ZlpvOsZvLRaKwkcKxnL2is+GsNS9gfhfFfZ14T0swpou
lbo8VWyFRjIgfxht9RJA+u/Dxkjh/03ARjlXHe/w7tg9afK2K59sREUwFeqY
tz2ITVPvnfbpE0vw8Ajw9ma1GteFUHDIBfLpn6sV8UsSc/TguoPWYSXlfpJd
LJD7nHWu+xSLx+sFQWfoEx+it5ErLIe3aDUzNPFwx/buGO/42ZZKEv1LvNRN
3ZdDvlOxtYNF6nUFvCzer72oSID1ipLb6NNUGYxSOieqXVPagkoyj1vnWv2y
smIsPVJTueyRxyZyu5hDtqinw6lnZ6hlrq+7/bfi5ppVKgfsQVUqgl+y9aFg
CAXaIDVsFW0pHAGx2hj8n2iwV8lr2JsJQvBw1eCKpeNGHFADrtN67AyYTt7W
707bvW0mmPTzF25eB3YjEByE6bhXnqMnhQA3ecvErnkdRc34QV+HG64EhAun
f8UjEDXRsjJ4YD6V+wVeEnoe89676icJtX3ph2HXHXIwRsvJM2QsMDkQ50Yj
gi41u03pvUlaUCugavgzRhdbNYJec/cHvXGhTN9flePDxjkdZAas8jTV/W31
N7FIoxJYQZ3dXmKbAqvXefk0QtQRE6EN2xsEOhKg629hUZaqeZ5FakLndSBT
Pc+P1VVYggjlZkLzrOvJmXE43e6TWxqnp+OiWSAB1WyknZ3M08gV9d7g6Yra
efzINxCEqrcRfoCHtCFUQdzG/4JiWSnRjwny3HlLOwSnCji1e0ka2kQBysxI
SvzYBzy2mG44qe84lkUgIREm2R2CPoz5DRqK3cpoNA3XBDX6N/h6vIOycf+e
CSnspGVH8hK10P9yQx9quQZjZ0diCfmuNF1CqgvGHQMOArS5nWgG5wE4G+aM
xolo7g9r3vUQ9t6j1+yVyXqbkp7zEUN/OxAAuUPtFJJuUV4I8H1qOnoIgi1S
sCgy9ZG40Gq0gJMcEDLu0iNdj22HTyX9M3oK6ygWBiLH3homLl4R9AAafmuB
rf7mIlNywxBKxODRfKd5llspceT9CTVJT7+2MDggFH4QgbYclDCBDZ+O4z/H
tF/ij62YYRs1gHymxEZ/kHun9bJperB6qIRrfkGjGwkDn0e/FvUKcqJvUmPQ
2Wol2P8F6UovflfAjdS6H3aOTY+pOI8DbnB+dG+2Dia5bFppV3ilOgIVgYYT
g62GY1e4ef246E+T26/CrbNIPraV27PDTsSZwId0OaUnoAks5s2WI0zoqQ9/
GM09gxRWWgTUHaDfqHlnkWrojGJK2qMk5hAvBATLzC6AMmBZxTffmzeRBCYE
edq1ep2esugNXmAPh8oPf5HfjaVuSqktjF4pszF0cuTQbYA3Pm13aTaSNcP+
4GnYAeTQDbvwdmZ0sroFVZEM8zhs7MenUPQVYDC+mMb3qRDFw7+Ia6boI1/E
Mk0VBONyNVFEJdPXRpHOFLB+FvK/KgUlKf8ncgLoH+2fJcOP0RBTlkw0V0mG
lhsFaK7A7h/gHRRtK2OkDxrVZqmFeWvYC1Jc1QHkIuZC1mEBYQYWCUBStL9F
THjG7nJ4EpYp/Lkz9JVsxWl3GkGQRmPuik0qAnaaitFwoTRsxo9QuhtAy2I8
7b7vq2g3PFr3HW2l/zPxpSZYEHCgoARTh6feG5Vns+Oqlx4li042RyKCXALH
rRilhPTUSTH/CfUbNeSboE260P/qfZI4dNEWa1d+GQwGwt5veO4JbrpFQnlw
auNdZYULO7z57mcFBBFK7GbSgzg5qHFNag2LWa4KPrRUG7lyWyX3IS/wn7GV
iN8ulqqouONEQvMJP3DJHJpSxyLYatRUsHeGizLddLfKDLV1BTDJauhEVqnq
G2YWqcbH9hLIVBo1CSNSFO5KtLjFU7Crya+XDwmJhyqmqrcv/g3aHtykoLY0
8GlM8X40uz7BX2OUggm2HqyOgy8q9NZ3O4sXdE325r5EKvp6CC7D7AXgetn/
P+hsg3OoeukxDS4AZdtV04b7N7+jHd6abZSxWv0Hi76Lnjl2Q9IG8+89uQIz
u63lJEDi/nJbwgnlDAhRUe02pLJRrDkWF06eHyHrGbyG95GEI3K26dwMwPrb
3ySwFoO3K5veHnPZy9/OR/m9HyIr0mK9UNClOcE+5hLoFUrfRwTy7N6F3vMN
pjvQoZSxlKgmMrEcU38d7WLOF5QXOwoR7CK3sOKIHzoLwiq6CZBqtckfsoCy
FgNseGFQt9ApLuYG0dFBGTD/FmBG7ty4pqToaeo2D+9wXSj5UoDS3jpxowK/
tXO2c9/0d6b3yzvkAkR3Amxufc6yTHeGE8xvQ1/c/EeNZcyRBrNbQ1Bgwz4h
rIQYX57fXb8L98DMZ81vy7b0ntJdl+haYMRN5T3Ug3FX5d8RTvwR4yRSfjTx
7UIDrAa5c5tqyFk1AN0t+zqdP3JWfHEZ84onkeX0oR/6g4umh11PXUv5t7e4
Nfq1Cmw/LeL30bNSOuTF78EV//0KlSEPWsAiOdBZddUwjNCP6buR74Mh2s+U
ViGeZQThbBikRh8u5cWXhBMaQgwCrwENbDpyKYr3J+uA9x1UVIkf4NyMYsp3
iSzrNy/ZvgdKSj8rXcGAv57daJ9jQE+64td6FLzigq9dt4XjBYPi9ujR8Im/
P42hI5ShHOa4aO9fRkI9Jx/ORNh9A1eJfriNkP4aiDOP3YvRgV9Tgkj0mx/w
3FS5Axy1Wnv+s5z7Z+0dwZv13+U+yegU5IKgmRoixHmDEmDgXq38swZN36AP
xFziaoSa63GVvJ7LGLB7X0FqUvTsZTDCjz/gg2qsWAE7fuGVMKU3RFNQ6oej
eXc6UsbTykH+SMPoYIDb7dETtRdUDmtaldLcBW6+f1klC6ICXfQ0rhbWQOHQ
4abt+N+INnGmF4voL1fFq+F9HlWU+uJ6SviYoywxH/ZZZiNOtNqPWfORJGP8
E8xvgBhH/jU0lo02HwijkWS0eo6y+W0uu7UznNjg1GtPHPdLyzpMC4916L3t
CuCPEWmDYT7t0vCfmOPNGbEujFQTQGF+MhKQHlW6Pbz0wWfc81dS5iQAtFil
syTus3YOlE0YKs6qOfZTF/vBUAadWw9o7HxuAWr6A3ltgEmtXhy/58aW4WdC
PZ4J5SzKVLshy1Lf0ofeWNP4p+EnT+nJTKp8YeioL9v6P6UVKaSm6m+GTafj
As3Tl4KnWBKlpRORF9uaZEykjtW46KHk+z9CXrzV03BCwJ3Hfd7tJ//oHSqH
t2tv/DPAZ13U4ltF3baJu5cLjIDz8IYttBwUDsHdlJLXdBMQSGrPE4cYtO9R
qpQROCwMKoQ4qD5jbYwp+Qbp2n812p7ILMOt4/YLvmPrra+4I9avm43mgi7D
ZfoFN4mSwNqlis8VTa9/71JM9rFe1Aj56sTinJ23Z2ATbfjDZgjltpoyeqHj
3UDFNT9t/kAxcpkE5rdHafBXVPDW8MjTx9EOJeFFK3OaNwATTFJXhbOvI6/V
IR4eI/XGaUSMQkDxDl2E/kD0nzn/yWwV9w9E5K2P+oR/M2Zc4XelgqsYudR8
KNoZfR2o38/nSMXR+XcXb7NVzI13NVD3IehDXRUp9b7Pg5xmp8yoEBmIOjbw
Fg2gHBITgsxEKTBPSzoa4/rC2OBGynehTpnCdZZSuaKIqUgMQ5zjeWk2GTbF
2FbZ2gKgOnR+ANHa790eDHOet35KRbaUNhj1Zy4bhmpmIgpqEfdB6LlUgFTU
GkHyK7dpj/Ndjg6aKZZApPZwmL2MQtTRBwl3cEgr24lqX2ono5VnAszMGVrH
GGJbe+b9LAJODGLVp8Bd7SH55Zq5Xke19SPRva/O3wiZ78fCF+moX6ao+sSD
7fgMTTr0dq2xdJGyJCIrkQ0nwKAMr6CUzWjfprT0YDP3rb6sSjMV372tF3Oa
e1PspJxrcI60uOGDvIC1AQ6A/PkwKuAputCWen6dmXAMXODo7ieVm2YeqsU0
8OY4iwuoD/T/CUnvBQg0hG7MGcqL9zFX6zbU2v86jPno6faokHrNxi39kTEE
ElUrU1y9lmAbemjfqAi680D9Yvg5y0n8Lgt6S9MN+adQKHNC/2OApW97Wqji
3CsGjFqspuTmKtR7pSFuZGBV5JY4EtFv3V59F77FsVESuYXDv4LFuvgximYs
t4Y/g3i9WnmdXEtg6fQTX3OUq4ae4FEG+8+pWzAayx8JXvIbm013CkoW9Kti
+i/kLjPUp3x973o4rFkdqizHlzNOitho2GcTELwP0QhVunrK+UsVH01PbC0F
MQOD/1ZRwu0xrvnlxMuueUqP83m6+qgNGnHCuT4rrFwsG5LYk+JzVM4n+n/Q
ab76b7Vj5qh6nxLU5WYXmE+ZFJ131y1Txa/R7jse6TrFIjQ35voMybwykqMe
lQBEB2RKr8ULsUE0nj9V8+eq7Y4+oORbsuzP5OxKCPsL0wCHiPr2pOxMJC9l
Zuq1UAv8F6jK+xjSLmEzBmLXsx6iJQXL1Bw87ubNdDIKnebWoeHNAZboIe27
hZmc/WWNjGRqRXlej3cNEb4cL0+/L2Gju/Bq0eba/X0uwXE3dcEPUDfLllj1
36BkJKS+fqbbuHzNSAZsOc1pGUBpnXeA4y1/sSZfI45Mn3lFMVWSWTtnzHan
4GjC9gU9bxuZoJcGXKm7SCtvlgrQiHdVmsKHdZv23rDMqNomrRb5VyRe6qa4
nwL99CInP3HMyMf0p0++JN8pFBgeMjRqeS+YgJsl5/H1KQtsZc1D06s38fND
yIF2/1bUTvQJtwtq1i+ZRShefaTTB1E4sEhaNimD1i1kstmTLEmDPxiQuNn2
fuFE2btAV2CcqSQbLCTwlPaqx6usCr4Gvt0MiS0Vx5ZUmnZgfkbqgyz1pKCI
JTCnpP4vxi4kfAr44LZTYmlDnj+bePOdflUmS/zsFXvP+Of7vNlOmxVmjkqT
13CD8quyJRgDsYuhIh0HctkwfpUhhknwT1Vfk+UJIlSAIflkJqjG6f84JGyD
/4ToECSTHWaSINIeTMMwCNpxhy9ZGjrCXh9FzwsXzamtSBvfM7o9QlRLY4Fz
7oeC4ISGuf+BwzLR/KL14MmgYHkYpQ2XQOa7ihIzpHEnCJK+YILL40liu6v5
h/HfP8Pf+tniCSUm0SNiA09jgonJXLRjOBHj6UJj1U11Cr051vK9gqbVe0Vj
hmxzFu8+0GfV6BEykWC/yKT/HznmFj9jnaO7KaomktK4gRMiTCILFxBX4eSY
vZFhkeh3ah9taO6ojYkn5C9/tjPPqep2CZpkG6ZIYU6WXW0060otdfPaxQft
JUQEqKmDqb8/1V40/ZxgP64k5xyTRf8feFOVOitINgt8N0ZsoCrPtLXd+79y
J68q+hjC98wDJ6BV8JJioiYOBqbxlry8zBw7X8aQJC8CCs9ihWzb9oB29/Bt
4jeSHsWL6uIWPkAx+YXt1/8lcNYaZTggWEyfMYPhDgzuc37vq0SEamwNvzdH
uX1yCYEe806lhZM47RDQ3olNU94eogpgwECEi3nO5r1nBGgpfC9iIXrbwmuT
pS952JXsisyEoKL06HxST/c54rjpTxeXwxtSwvjKY/EO7chG4tqtdKgqmcKK
pK4MTgExebWoG1MQVdZCrRRE+INPcy57FrK0U8Mgoaw3kej1FmD3SdFCXLLs
kqtpEbKcdaVmQ/CljFunzyWMk94zu/BoJXuSckuFAbRSRIr4i1VMlIAkvgUD
rvQYkeijRnIQZGGBQLzgX3XAstIY/vjpouy+mLaFqza+M47zZ8U+9pzXbb27
CY63V6vn8j96WRxGqscm0psSXbeL3c6oT1Wwg3JEc4ZyvHQhrCsX2I7xIxw+
V3n7c4/EJNZ3gkn3GIkbEQ2gsJiuvPeMsmywCF8b3qw5Zui60QeYS7EdLqLO
YxXRicZ9A+3dMWNYUacHqR2vwgBMW4pzXxD1Ztgx8HF5nkwtI2E7s74rxsqC
+xlWVplAp5obeUiCr/vujZhVb0tO9/IFJqJ5IC/dd8eKAySwHqdqcrS9nc8v
Zl/LP5mSqVVreRPG1vTrhIXFWEONMcZFhRJhgd4NjV1prrdk0uIsuVbXTcIN
gLyp6vwhRB21Dh92m7IPPOGE/7aUlr7ly8e2qQiMeGNc1lcuntA+69udwzij
WA5QNGWHOnttT4XoD1trrNTwej2Whv0bC5DeZcuX+GMX8EmFQsGipME7qajD
kUW4e1ryY3gxxmdNqqviBevPjnHL4KKdxGNdN7muF0ZxF+f4WPpLg1mFcxsy
ZqaRVnmTMPg3o/khBu1XYDfYo3IiJmLNHatYTu/aZtOkzZx0j7QV246g5f/k
nKNOfHCC0dyLF74IgjVGd7Tk3w+PQ7t9+OFR/aZlL/nubjQD7C36XoFB+tnS
mLxwoiDiYFdgy/D+im5VmfHzev4EOEPJPlJ7WyFQ2h6sfZ6T5jG0Xl+93Sek
hs3bGU9fVYQWv38RR3mXB/6nGPftR2UaQv3R2orEKYveAprd7I7rOFvC0Iev
iLuzO6udYXdInQQSuvwCJWeD9s9BN2/yDMu2e3PJvAKQVP2NziZqt+LOw8sQ
Abjhet8sqA2tlBDTgqhLJpaQdMrsgV7L3IH1ockVVytRgIDX7FrN3gRSgvY8
FbJjbTA88qe5ixFhEgxhQNw/rUQb/GKUlwxMPaLKLbo2GUcOkFhjiinBupOT
tC3w3S2uGuP+rPaCtkdpdqrlk3mue2F7GVQPTtWDm18h3x5uLmTk1skax726
PdclPqi3dnoZ/3g7v6hNoMa+11hs61UWeZp6iVSAnBizx52VwsMJ2530q32f
FLVgbniQliIFCVVeuXDfDGi6RMaHCUk0riPcappxOys0Aw5t4tSEg8FspNT7
AqMg+a9Wa29Ai0tazcbDR8YLhTuF9OZqjvKWHLH0I/gdOZf2s3KJy9zs4VqS
+mZFambDy4GP9/RYLWlXwjQmTkyLPuITv6CGwqnaUA44jACXWuM3x5+aLYpb
ftwYe972Us4GecxR5CbODBhHfQWxwRq6e1viam2Fjnq3a2RhxyiXt0lPYeUF
GcTTxnO6RVr3IfzuloDkuJ9zUsPvHPH5AGwJXyWbgFYpJQu2fQWy8zyO+rn2
fmXtzHBRXrg/Hke123bw+kTwWmEOD2HOkcD+gbDndNBDiCNU6TphPdIwi6hH
Nb/LPgptGNl6XYbmL0nfTKKomkUcRLyEBrTEuDeOcsyj3yA562/i1w+RhCRF
M6wE9VlEsAGj1s6tY3PDw9K5M1cMxJJnw1xhcG8BeR9AeRoFXm21r8lvXr53
jdyB0c44S+c6R38fBQZyme5Rv818xyfhqtM+AQuxvOJSFMCsYI3PLNft1Rrz
kKzwgns2w9YNJIoHAa4Z67vEt6DzawMU3MVT8VQEtZAhKcrsLrFyjfsatSDj
KctEZDk61H69Pvh1SgjcX6TRViPjABCloZdXZ20GlImBoDHN0mvs0OBYxb9C
Z0H4injOmP2LNSpIUgrTLErDuSWG9QodaLxAkzwIvEP6f5X0p80BslwW8y2T
iSf8+mNQV6d+8otRx16lBUrBbDeCWBGXGdjZyQi5n4cbJkksF3HcPS3qUDwn
wXga04WZKBGd0POk53q7WjqGCtXTKSpZbYvTqRrdnCCJB63K57zJLNsCyrnd
uqYWXuPequTG/p3txEfruoxMXZC2EQbWcOE3mmHzpCP5Rctr5DbkGD5UZHls
G6z8KdXmB2x7nBb//48EDlapoG1IGAHjxB9WsA26HAfeCWosxLwTFHoYL9Eb
MzVZRhz6p+Jis8lzqr/HhG475Uql1NsR/WQvZC+TbSe9v1X5WaHqy2dbK18T
hheTQ8C6y9tiIfdN9vauw93x5e4aVCAFWn/FHkeeRKWVzfjtKBvZ1havw71h
0PNpGuMT/75fUUYqQwXuaBVMmpWoIDsBv3FlBMtc0Qutr3VCvUncqYn2cLG2
EqrUutkrBs3rzL7GSbLH/xH3BGK71ntMy8Bc97ErI63W9K1KsBlECSduTFfp
biMlSepE3ZoWDTA9qvEMdb6vW+UYJf6sMP2uALiiqCN9qzhL5Y7cbSeWntLt
9P0h7LFC1xSqL5x6JITwmnOcGiUBpVy5RMerVI0WVgADYywraRugVtHdxuq0
AsW3zI8rzuBBd0skp/v3feZTXr/mu5lP8inRQmRW9VnDQPZuiTAW9sqlMdYb
9CFLADCXQxND//QHiimJO2kRFHu+US/ylpOXFOaEVwIyEvhDrYEQnR4grmvZ
+7EnERBeheixto987qywWOy8KYSJIG6Zb1N0ZWIDcK2/Dl+KJha9ade1woT5
GwGYJQbzmuP6DRlDOEQOzqHwoLgb/x4348VC4DMvtR1r+v3Qg1bX/ZOyiKXh
2eqvHqWQOr8h9veDsy6Obj35jFxBOR/7ii/Ziufha/CbAaEOq95fDbqi63Xa
io3Dnn75w6B941kaTXZvZxCij/gH5lfaaM4y2eoLNtQBefXmqA6QBRGn17I9
8TdtRmTRD2ibiClkLZJiTcMR2B/XBubTOfO76bRlfP/8FOg0168MfWxS76o3
pI/YsoVgEMbR6kdiYhuk89Mqx+x57rMTi0iEiRq9QDpISV+df4Jxrpf5ppF9
VjAcnlwCtUFDs1t9lJDu53uHq5R7Mp7XRYHQUGsv2FZcsjx3x9D8lLS9XquS
ig3OW5R+8EAAZGQ7pjW04oylkpDL9kbX3n2wgc2yz/T4VWJeHj/vqqqKc+A8
rLMi1ZjPy44QvUi/OupTd9/sQ55At35jPuvPQ6IaK36ppL3jTHmA69xof8J1
V/kJ30EmuJM8bgaS8vPX+aqahieht0msdb+M8vXulQqO+ebZdbhl3GrpRscK
lnoKjvJwtBwh5kxybGV3RlPlqCgAcHXGeNpc2TanuWmmP/9/Bkxs5w6lDsrQ
K3pvyb+RgSTUyNGeiQfOg0bw9At+8e2lHK3HHC/da6BG1Uf/kPhob+S+SmfP
69cSCtepudJKI2mgXwjPJZ0BzsrW2ZUYErxakt6+vUWtzllUUPoQDfazky7a
/z+unn8l7YfLGH0q3v2yiKPGn1yth2ajMcUliUhSpZkZVwl/ovZxujbpAh1o
EKeD436S8z8EdXJGHl7tVT2Cke6GthoZcKodWF2KnpOIYIvLXdzxt2nU9GBI
cX5Vkf2N1p/jxMRqdU03rvzZDDmwFPTkSoO3BwvMwXePdC8P0iFeSUO7EDaT
hiCB9VyVbptb4Ds6FE4Ad5uuVf/3L/4SLRG0uTeHz0xydYV4iyvce2o90ozU
NgvfUXcJpZn5yViQGu8I3lA5pmT9yfbl3ODXET1qCqMB1B+bR2OOu48XpvMb
NNzGXjtjtLgMPBsLj+tLvidy067dIw2uETRNd/pobiJqqkDTZzK0WpzReLET
Zf+2zJqopGQMSSvzvOJ0/aWnVk1BFXZWrz37UJhd5JTCvHfWbPYJCqQ5pPuX
jMdmUqsX1GTQ0qIrGT2pARaeHCJiZiSRKopv97Jk17PKelJjZ1An8Xs9/x9S
fXgN3C1NXQ24ZOQqqKwyzZ7GTU8LYxuHf5SoLNcBGmmzmSq9KqzrhAyMgMfh
Q66i4JzBRlNyz5LsHLXwr54DbAb8fRYaaB05zgtxgci1qrZABaWwLCLBkcC4
qU7urFJWf9COKAX/lpAgCEA6Vv6OwxzuUgCAs8zW2HWxXpuBwujNXKYb99Xt
XTZe46eqas5TdWsxy7hXpPcasLZ3CfOS8grnFq03lyKyrDT+X8oPMRH21mZ8
w8XWemdBBzeeMhg7ObgWJG1mJ7aYOh7sMTVzb8Y90pXSiJ/oCjKVO0i97qtC
1bD+U7/Nlaaj/z58/SIHDpU+494w0t8PJT9HHWWegRMUI8qSkGsY8tgkqLct
k6aMQ5qFnUQ6cQRe8XGWEutYzIVdkWQKLALdoWIqhsk2wN4YoutUPTxPQdIe
4I8Im4Eyi3VX7XoYphWnRUu2F95xATR1avvDi3nsMJ4pul12wYXohS0v/U3d
+petMQHUsExZeZexPmD7DREEwI+C1pu3wiRsctEnCOgxcfwD+O9fTzIATFzg
ZP+A+RvuROVmT55c2jiw5whj/hOdYH7TWbpaCReEIKUzYf6UHwX+/+wRuY5F
C2xW/3+b/doe/0lk2+j+a2pAB/4ELplXtX8GYMu7a3eAJwIga137dnxSl/3K
RNxg67UeJuz7ACHJq+C/QF8e2PtiKs7JgIRza5dvqd7o/oBmrc9XmzPXDRrY
b0gDC3C0T/IxnrT02wsEQVxKHF3tkfBxcDv56h/LUrYet266RVpBFL52mvqt
EqXAJeTIwEQYv2HOo/RTU50rnF8EiCHX/V5K7nQQiTNQYJD9sgTe8ZsmMXtz
rc/HwDzcpp8iAJfAe1GOqMtVGPp9nEplAATAscOQFJ598lA2YnPvHq6v4xus
s/gmbDvteBsMkdvnf/5eZFKLDUf4XMmzoI9Y5nfjkAYUdy6fIT8tCtocNTX6
krGCXpQtdYRg7JbpZDqS+DUgeK3E28Ndp0wCq2DI/l5Kbb7UM2X7lbNnoEN0
e1wJdREd/c6fXY2npPxI+BQEaDwVnrnKXzXIIDX0a8SsG0jIhP4NPXVqkHWz
Y8eYUqmZhlntWZZHCtuDlnHz7Kq6f+yylLXPSrh8CwKwlNPh/KI5rpIbGWlO
efF28DEp/3D8PXTrPkKME30ye7A0hHODGbxzw5d5ykexdxAn4jm9q6ZM+o4d
KorDrFsPc2zMsoWNQ8brQQ0H2yWA/nd22rF74HXzpzUOPRF/nLamyPVyyvXl
U4K1nBpoMmJ8CL5016Czaf8S5IKBjrPKJz6Q2DuaPgqVa8EHNhHseFP6P5I0
l8cCOJnwn6Sdymf9YkM7XfhkBnSVbfsN9GwIw59LCH8mW2hXO7d0RfciybIV
XW8QoDsQt9P5vI4lqmgYTPQtL17qcvz84SOCCmXd5TXBSYbVZ8Dqs4Ms6b0q
fYTvsbAicGYs6qnanPZyWo1bsf6q5hDXGNR3guk5Cj+YPIZeAi8hiSfHGY9R
BqaPOn4sJ+KQrIgHm82t/OFEycxFa6dlfcIm5SS57RbFK+kW8uYPEYTvfebn
GwuBKfJYiAayUsX8nCVvtWhwFsfPJDYOrya/Y5S0NnyLPpTJs2t4Rf6SAfDu
q1sAibesYQZlCYJBOx9OxDixtSuKeweeL11pehiks5D4I7zo+CWOHyeV162o
uQjbDOZbc0XFcgOzb7xnvyBbIUWoSnw1BoTmN3TGIFKcxujKhy0l4cXmG0Vl
XL/pTqxuPSwBBy6LWSRpHI7wCNBNOVTNsxGW17K2QhaRUVgE+LejVqAgG5e7
sK63ZY3LNUd7rDKZ+MBvGM+r4QNKg6UbmZJhxslefhOWnlhJtvF7Q1y1UBqu
DAOG1FBNz2IU+7F5Gw9tJARaOLY0Yq1BPBn1DKOQNx38e0LCcvX4+Q8jenDX
dsHRcp8NP2sSBGZmuNrANkVV5tW7Prd6tQWvvlww5SbU+rBjHb6ARRWMD4bP
Wu5V+D7gWkJqn3g/sjRcIL2emTN0rVVj49KCELHaBpe34DOq718C2GfRSa5V
iT9s/OnwAUA9SCa0d7VRSFhRP6ur+vukSYbs12AIBuVZZmf68HCRBWWU1MUs
DdgGWUiie2eF5d5XNzWnzwXRnXqSRuaDJTdMCsYgBVjDP46FdC4W4PELk6Ly
47T1tSNrV/mChXXj4w6EhJE0INGqbpcSwyGBc1e3v+1xADVF+HQyaOybnIY7
QCH/vgCddI2aju0TC8do0n/dRlsWkNCOKS61VhJ2ARdFwhjSgaDOOmwOmeHg
TsT3x+B2jzFWRbpfOXTbpu612Ih3eb5Z4OM5XMzB4ZTKG84i6dthVx50Z1xB
LzkDG5c6mo9KI6Y9BAMpDJvnDjJMg1zzgGoZ27uCL+X0NunRQ7ngI5/Tnosg
8/v0AnEFejUT8BwOwjWNbLBw0MzM4tDAjErJTrnNlHJmp2uvcfjBiY7rPAG6
8HxG13muqpw2Fm4vPwRV5ZekqyJBTRxw0C9CAWTvzBzibjnsO3vJgfGxHlrq
/J0kuB2K/rPtjcZLsCnmypyQZ/K2fV7phq3taMRuTdUc4+g3cog6v26jQD5j
drqvj4c8BN+Yc+BaL7s0pphkNFOoaZFMR5+RGoGfIRms4nYQHlaCmXPEEg93
PKIMgrt/Vs5ej4xKnMmU8rHUtrV2dRJfcGaFN9WLFkTzcYF0l3EbdEhysTpC
tbDRaIDufQog8PL60NdCGqa2tI/fF+1zkqr9+ygv9iOx3eubF10OXDDGNxKm
f9T8QRx9wgQ8EZI8j4F0/+64ab/iliXt2XUBqc4AG7Dcv5VfOgXMKJ7CYV8N
CLtmcq4RozcdJXMv3JH16qM7T0pzP0IZLAF9g0MvVBrLM9nlVFAKMjFdcaUd
L5Mvp2abxkPSOE9Q2gcXqaRpIQMOz7Yno0eABYW2Ci152jKKyriNwBoYZx7Y
RVaPbyvB4CSgGLt+8szdqzWeaJKDJsAtBLUMZhV3UFLm+VyPG7yacsg/NdlL
A8Mniw4xzvdAlhnWrj119vpvSgQn70m40MitOyOR9WpjHdv6lREPYYhelGwo
ARDUI3e8B//lZjPEsebJNHcmM4PVm7Xg8eN2XjAt/SiL9R5ODXeiKSbhwMKe
T0LqF551FuMOSvbh9MtXyEYdvvijIZxksnPbo8peMmjls40Z9JTh+0tXY0m3
DLt759tj6l8VcYGqdiNMeVStYhjdFvgpRToy2SnQSgcsBV63IHgh/c0lyeUf
G9FHKmj8vv1qTrpvPgZRSYaby11y4cGpmxJsUGQfkglYiLqAwTkDlwB5GJzo
liL4GmnnDkEjkDEU1sDZUBsoyKZFkoHu5wUIgGkM487kMYC3Cbuq+t+WRp4S
jo70pA8HPXlhLpagMxKtMtZOXQah4SBjVLrhpMVXorY73l/aJWr6djbbpBV+
4musdpP2C7v+IWOG91jTtY7+PfSZCHxapdFw1Llj16LpgFSLJineE74cFBHf
qepUCtMpThSZTQduQTSIFCepDpLlN4z+aj7YfmiLZbZ1PAydMfBwgr+sHyBx
fxyKYs5M5Hlban8XqKHTrwbvX/7ipHRr8CC4upzKvXZZduAQMGy5Sx/YLOqo
7GluIqrjFWMj5SftYtFsNtNGOzkzK28wIGspChn8LXPAdUAOBJbZK7SB8l+I
0ffDZvux3Y/93n5eIv9jv7IL/DSjbm5vjWHrfJjymbGivaixNsr0N0qZs8RB
zv24HvFwC42qEiHkmrx/9XZwlmv2pvMMoPq6wZXo7BUX+eKHA4dlLX1qdNhH
Wg66EOkDIRaSvpFGa74hJVlUtFJ4BHE0G/dVnv5138mIjIXP/XAjb1XYMx5l
YJzeViXW0dLG3wPbLdq2zC0lznO4UP+rNfXkZCGKS87XFWM+tmlTn540w9BS
RDVxwew+ljmb58h4wLvC9Ls/mkNhYsq/DlCI2KEXQN1T4xi/u7fiSAIuhB4F
C72BuohpFUKdWcNYfeTTJcCJnIkFWmsWEDdiHl38Jub95wC4peBDZOQKIwx8
lG/2aaQwZkliGEDPaGpNo/bDcvEjMkR53Z6s8I2fi/lLF0JehdIDGSAyh3p2
Y/2kzEowWiGbKfTkaqGO+hFhyokRwGQOwuOxbfQiE7rFF35pcFWCuNG2Nndr
zXAYI64fyeS635+rU77JDD1YPCpeLZXtSwY1Xu/GLhxfl+sXB3Oj0tF+gQkp
IlWs7M7JlCvxUO5GDa+9DHKksnnTm9xGH02iyGwOWXGgVE3tS+2y/hMUl9Mu
EZSxKjiLOUX9Gi9PK3lsvwrd9FcYliOHtfzknx6vDHNYEt/M+xCJSgxQbTQX
fLyAB4XuQ/NjxxHyCPt0/jVWO3qTkeCC3l0NR6mC/RXvUMGP/NmUUOwWLOwv
koeBHmFTAxPVzhJCip5rri5OmBoVEQSSRZdGRhf0p9uN8mNI/PFhNJHJcMDE
vAeA4a+QwW2D/AvKYY3gSd2NhVt2fnALtj+fyIfAq5mPpi0qMBzMgFww5faZ
7A1rP/3omRFcLm89QYVBeesT5iXGC4SBOygjRz/C90CVK93t2C8DaLrjvcZi
xo+DQSl1K/43lW3kGMPAeYdfd1vEKwbJliBojQyj8o+jOqoC8aZF9wDVH/Js
sEbQalZOgYr4Cib+jjDPy4JfUSddBnPeeYh1OIer/3pdwq1cLTpw+mAY1j4i
h6p/VFzmcc+bjFFXVtIC8EFQOHqA0+c47xsjoEPrMAZufsHVtX04CFW3BXbt
Z84pbWAy658KC2lGrtbuZFRwSNQGaJ1Pjh3gak77F1zOEJVaBBIlqRo3V0OW
zyVvqFiIvJSalDkp4atywSysoEuDkMIQgopmi9plwtoZ57fQr2ipn+Yon4qF
Y5kqrZlATs8iQapBU5dIOvUtoGEy8hUAlxVdVY8qbXgz1AzeYL4VYIeWEFeS
eGhwhTJlwtNxWWQ4A+04IRX8K764iQJUDItur+JaMVO413tnSuhbRDgH6UYA
OCzg5osrLAih6zba+FiHgRD0FFn+Jd0Zi5h+vPY2tSvCyQm5a46cwHfRtCHf
wYL1BxyMohWMv8tGiDpDBL7s/M+CmJCLUl3aPNXELARKnUG6N8aYxiErP7zg
1u+T5I+nme08QrfISOKqps4wSs/y063VLLR0AEvGWjyuVGpk/nd53q1klqkp
qbsfzySNqK/8xXEERi1rw5OWFXzH5t4GKV+LXvCHyHO+5a1ic+a8lvlDXILc
JK42ZwiAiPjZwxvIEeX/RaMG1c2KaEBGQOhQCKXalS4ZEEj3NNtKLE+tqvk/
O3UuSf5+8MSS9SGFzRS6yBFC7toKCHQOYXE9xqvlZIr9TkVlfM1P5SYC4aDd
grsNvzEGAIUx2TgvdPHr7VracEbG7GE3fW9t/l81M3fCE1pawv4uBhma7/Ig
Af93RFsprlh6Oo/Rvuv93r1H9vl/UmXFOPgN3kvLVL5l4UIOwI3OyrTZQyos
C7xrRT8UV1D7Q42qlYQKUrovbC4XxNdCIRScfqAcjWasfd6PkJkF+0xkohq8
2DZRYGeQ7mGK+ZDnRtiG7PyR6NmS6gKRcjowxOKYvGg4W8N3oJCyFZZ6tPmi
pPejeMFlAyqXJXuMTb6xIFS+9G6Vi68DuL7trL9LLEPBPJpm050VaQgKsakg
Td5opYhmAUl/PBceZwDWsN8VsZRcCNoUOcJostuGSPoOhmOET4g6EjibkTO7
p3j74XxPSr2mfDVl4NqIIWoHKs6hFTEIGmhT7lHnOGq03QU3UyhRgVkwuvWk
4hKm7G/EluQIApdi5u07E4DLTBj4oQn6CqwyxtYeET1cs0A4ueR12p3HN0Ub
tlpj4wL8QGTU0KmngOgqvLfU3Cc/oa7A53gH5SvIHOEjG6Z3ZvfN0RIZyMca
IDxHpKD+G3HFerzNVsmfmlwvWI+n+BOXQmVOyOBJOcfrKrs1DExC/LgalOcx
6x6vaDVWU261OQ/SgYk4qKcq3z+WMAU1HTomImuqXoWbXsfmq4v4E+RnQbBO
DoGhXqgJD+b23z0TfBs3jI1P/nlFtAXPST43pWPniUnjePralwE05P3hOBuO
qH5aW6b8jWUptI9ZF5JAdVnF4UDSaVs5+pRPR4bC0eMlgqQ9G0d7hQoaIR6D
u/wFSVn9axEDjC+3GvJUPhc0tofsBCbJIiZEZQkBZHgIdabuoaawjB7F7SPK
Tlk9vE/oRqWPw/05RO4CrlkYhCnbjUOlEV7VEAbg4mAGYvv2Y2z1fpC4ZuU6
0QyhfM5fTVeKs/3Z6zKF6i048Sc/92VLT5FA3ys4GFncr4h68pm5soKVdQIQ
r3WHggnYja8zHvLnCjQZAvh6iwxAiOiyunYBV4h2oO++kh9UiV1U5bv5/lvU
PYXhdQZN5pPvwIBcWG1MDJkRZqCJgA3MMuUN7Ita68fKotMmFwOJFXIqzKfx
nxMkwsTUByBpTfNH9vG/aMv0+nv/GpI3eNW8SkwZq5dnouAwT2HEqbMxbHNt
pK3MwbzpiJOQ15nCk4K4dFyi/9v+/TC2UQ94mkq8fZvdCNOVeBWtgrjvhUzs
+afYtTWG7GCjwEGGVSdnjGOYzArFYoHvGTchAxSIPy+AolCCOSfKctgISAYN
/K6ol9s2fJ/OZ+uZ7wMvdYBNjaKHzpBriVUlWtb3is9Vm2QZLPKzcpjInCVu
Nerv58uoGXhSjPVCHmkVoqwJfpelzFXzQaTETK15nsHBSk6XDF+7siLlQNAA
fKlp1rO34tRBzQokrZIym1gmeae4hz3pqO2p1Bb49OfnLNLEromgpVI8/apJ
VpGRzjWKalucCrwFrHEhE/txiEFyCnDsq7Bb2jwAdd60u9uD8cofSelDLLnA
6WcF9Aaa9QXt5/KgsIebzNK+GRH3haRqS8jtbdeCGLVlnLfAMFRJ+Xbk3gwO
Cujy5R8x3TUY57n4SywTVXShUDQso5ac/VsxViVf2mbpP0cINmdCC8smVEM5
3MPt4dodHSdtUOVf87Zt1NbA6d9CXsTkWRbxZA61jAMwMxqSLKz9mT8RMFuM
1KLNDmcZX3U4jTFvxPP0wN3bBYlsBBub7JDz3BPQik1mt/MMIiwSYPC8GmSQ
d1vYl3HmRsX44D5hh0ZUYy8jW/fCQmV4/QWwiJLb3aCLMYeKYJ7mM/LdJyWB
Zp3vN+Tb4HXFJWyzcQxlmPEHDh/45+dAyBWqLiPDzBU+RzSq7GH5VzoxO3a9
OwKI16s16zwDSqKIPidnPBM+Rs+eqqy7V1jHvbzhnUbPBLPGF8t82xUzUsVQ
Va/r9zGZ6QGhxJTZMvxoSSFD7FLTiePHbmQezbzBhLAfIIpZkLnPpGYNxRiv
6EVbAxoTFAKQzoW+KWAIQPfvs3oEK1fMedX6M5Hcr3ovdq+bCmWWZDGmtapk
VxASRx8EJkekuqMnsHLt/5nnkqE4TklkAVozHRVamHkpXfUMxpzQVUt3lLrL
TWrCt0oTObG0zVe013SGeuhVY2wFjCsj9XYpeI+XJbA2Iu6srqjinMhBZqNl
5/xdWN/PM9rXk36MdWSABgu0+M+cOKkdcQl/sbzRIT16Vf9TKaAXT7khXsRH
BwUuUNbAag6I57iqszqd8sQr+p9ZwBsMtLtYfRRUopGeg7nASYnvCslAY1JW
07mYEjB37n5tvt8thFtEh4eRCipqxjKoYCcPC90BBf+1Fg7Vg0jv8qo3LiYQ
AeKpkGG7NBYwQ90Furdxc/R5grh1/41tDT0YnTlkDEHVMaUSlkyNULv1Kz58
wb0hRTuhKi+K+wol/P5JjKgSqgUhHLXtjTsz19ogjdz/8bGehGQv2JgDFbFV
GsSO/FNmdfmot3JY7HmGG/D5sqt/JVLTK+Va6vYcmWOyTbAkwKv+QQcEeOX1
ZIMC/C43ABxgcVrfaJeZjzlR4OzScEiZys9d+XD8IayfyGFH1ONENPxCj4Gx
/sVrg4XHcJUOqHyF8sZQoyncgcpTJfVyplctYoRR3ZVftxCIIuAudq320Sd9
Pc1FIwCVRj3Lw13j4U60kpoK5F4u9fY1oDNFGVqxqq+r5JwawLm2lSMryed3
/a6uFEj2ersrpk342dILdpd+n/6nvBJzWtPng+GqkJ5iIbKiWLkxLZ5DXMps
kfp5TntQH+u2LntxKxdPIaDzqBsn4Rz2xctcdCHU/q4DAr6X/Il/wghc4yE7
pz/tN89Pkjk3QJa/JilN5zdsxlb/7pTuGzaOTfnGMLucsYkoxQ3kX0+mCwZg
jMI9C48QWWqKRpUbMBpU8dHr3/+73EOLFY2ViMbaj4JfRPUKcUtWxZeZegee
VGcXUhYgztdyFJOldtZ87Iqk//FQm0EYNpL4tym6bzm/t7/Yj4w6LYV0QiLa
OK6aM81SokuaiEUy0aWFSoEu6K9Wx+pIaSak+gdFV1v5JZ/tnEW2BkMkYONa
FEb7PDwsAA889C7zVZY61geiy2G3F16xHH1QyO+kIL78XrRxB6iRejUbYWOm
nJ9sdMRgQxwAML2LmMn3JyC890O56te9DvWr0OH86ss6+OduSjWN7QNtYIx9
h46p4py5nn9iDBvsXYX64aLYlp1eGsZgfwkpFeQdft3PEWAhvUmwi7xvoE5h
0bFp0XQLpLnSK+7bzuJnRdtFwVqfvZlMH0mevV8ApdZehjEkI8Fp95bpqA7n
ZkcMUhg3bR+UAh+LFMrSHnYizAi5bq3XkpzcT/2maxNxis7i7X5OQhpuNn0x
xshBiBDnQWxst0Dayz9O0+YKxwcL5bnoWSBTUJGvNHl1xFvJEuF0EKk/Shpn
Tt12YTMWQnzaxJL9ey7NQReitsKGMcUpRxzum80gKHt50nTfcWvWqEA9P+5i
cumGBfpKpQdWPKhFYEyg1dFKBe/W1syISCCRqDG73qnCDS/4Ii4BeJd+t6Y7
qio0/8eEzhKei2k9ymIsp/f8jjmZdEs07IZQetlpB9Nm4L+4ssT2cNnFAsyQ
zKFXzUtOFHEefD52OfD++m7wJpNmjfWwzhQ6fjaE6d9ILiHe9aEuFBZ49eM8
4/Z7iBWSUzWyXlijBN5fw4Tux6U27ppBs9tQ6HPLsd/TnQgOibeR6X/wFzXP
Dkwt3EoYqCYpV2qPpFXlWf4uit+hMOCdA3+o1mzsrHKAh571z6g+cNrB5cSS
xu/prO+hMmPuE2OrR4Over6xvPBNE2hndxzquwkeZEn26jkPCG9BG4hSSU6W
a6AV+Vzw4fA4GBFYWpvaA5j8SH5DhI7uha2o/51Z4BFpTx4nlTwJkZJRDUSu
T3CFVP248xjzyiWzntVGuBjdNMDuxjkvFw1ctkgrdQNLQpactmY3XSaVDtWW
A77PXD6BbWFfUAzzKlXngar1OWYJVahTo6WIRghGtgS136DgjcX4Bt5dsLtv
JwyAZ9XmTk/vn7U614eT+N/IanVyNY44PwuhwXwhYgOkUJhLa67aI/mM05fE
rcUO7W6t374OR99h34CBUAV4qY2IqvxGgwnFX63sQNyiZQ/uqPuIgp5TstrU
rSvZBb/QbihHZNoD1FimaaeqLum0f0aMzk6CRTA7lKBlm50kszcMWkl0CRiR
YDcJWgeinGSe1zSAGg7jE61dthAFJxOh7MEZvMwnLUQG5qkFOO2PtYvDOZUj
iIkPPNGr8HuZ/um6/jm/23mGzFPR0S+T6XxktKm5S70zahw+8Yr81Vg9IAKI
+2FOTbegA3M/wxgm51JJz77E4EGVc1z+37HF4Uq+FLcVv4Wdy06CilBea6cb
11uWH0UiwKDIUdhwPObxbDvhscNLIKNm9Hj5qgkjIcPd963Vb/lz7yB9h2xm
kBMK273b/+F8aTbBrMIp9yh5fyzX4mbKLEqXuoP+o+Fi24I53zf1mQb8yEpG
W6zonKNTkuC/0zn6jakuPG0OH3D4HOoh9XBNG3o1l3RInhlU0Ht4gR5uiHKY
QBFQK8Rlv7vSd9c7d4xyZxelBA9Mv+0OaCs9F5gK53AAh/92h9NtHYgqGHVD
b9fQltoTdYc3IgqbSZP8xCb/IEVcHSYOgp6ujPpph992WDdhYExlSWrVVZ/b
qubqErnHCc+ui0E102UT3tczW8JUvlZP0zdngBk7GXP/8O9iCJr1cphcyNLZ
CDBzTpz2CwJit4I844Io60AJEMfbUGBMhcFrVUBjzRxc4dHoSlUf7HWWZozE
N3r6JZaVcqweFvofp1S9S/fYfQYju3h3zg5NVmG3Rf+ROgYQXgwuor9216kR
CHLxC/djeW/yZ4uNsrkI4z3FvX0oFmususmPKB5g8CyPK2E6zuu8osIQch8e
G8r4nCfTuGCI/g6zZC+xvyUTWiYBZPWJJgy3EA0h8h3v9mmAfjrDbBS4e8C8
irpQeuaseiF7pqbPO9m2a9ZYBnlxAm7/gApfKq87Rwi3M5rs8sRGe9s+xYmm
S6uvB/5UYYNZfzHqy94vXjgLjDXx9hs7g6yXyjtSMwj2tzZFkCsr/IuZRe9l
t+sweDb6QvB0ytZ1c+QhiT1iM1lltqFRA5Z3RPdEnSnasOeXqNpbCAduqJKc
neoGX0ETSYES1pFlkJDliRohfVK7OPLdRyIR2HYHLgfsU0qxj2bV7PQMLHRG
YrpVc/628g72DDB3F9GVnWGDtN7hFCRJ7P2Q3TGiThnGj2m6aYY0BcOMwpS7
5Kr9cflVJZ2Br0WOya64v0UHVKQLjFGlnOf+c+lzr9U94Nlk/TnN2DEMWoEv
0Z8RuOe2YoL5i2i1dq8tqY4kU2LIVifY6S9LB+Sx83t/ttgwfbVA4X6FYQ4r
13fJMgE+lEfr71d83zQw9Gn+eaWFKMwB7JaqJfKTqOTXRd1sTV0+u0NSitDn
cooyToJXvCtFCXgSKqDro27mEMTg1M7Q2c9BOkAsfupR5TR9rxfoWUwT8kHi
/a2UaLHjnbJ8pxGOy1bBoR3rxuErCtR3x8ahlcmVN+S87JOqxVv43qOXJ+EZ
giIo+P11S8ZM604+pAzcP8ADUvK0yVVc7MPgILUlPtQ/xhSuV+ja3CPH7QFu
E/GPbU6/UtZZ2GsGKlrPOLYYkayF7oaLi+dIzSlFHZNDWV0oBavGT84V6OgF
Gm6IFMD87WgaXOkleJacMzcifg53+QYe2k+p8bvjAsxjgE580VAm/usZV6wx
yXMA72cilBbYG0GMCEGg1zgqFZP4pLMQC1vxZnRGyC2DN6g+p88yELzSzwB+
iGPJs+HAQUwaOJVRFXPkZYyLiHj5pOqMRGhsOA/S9xC8EvuLvmhvZ8XZGT0w
0td5Ra9g9fkPWPp6LTYyQvquVSNWC9ug3p5LCvlC2qsLMrCO95GlZP02A0cm
GsBTxQqBM6Fu4RufIDhdPx1Z1EeoTrpiKVQBbZ9G7yFnLtOD9W783FAm8veV
5yRFnWqu/6wIN12RpiK2qzRT0LpcQwGuUTstrzmRYBAv9oJxvj33oxogHp4a
tVBVd1TlF1HXwi6FcVgZirSoBWIQqyoTIBtCFqSnNzsUNNYe2s68BGfwyNeO
NzbV0O4Py1jgExnWCo5EES0H1Re7y123PBgEE99gHWa9yzg5lK6gYBRp3BHZ
lIMWDADJ5tCZRoog4H2Rp+gjsaSFplogebILAGQWtCXWF/+0Bl7vISjQUh8i
1NATbWspeLpSsiDl9kTT8zXY2a2iul4/GCOYs4FCOfKDOGrbOBebk6Hvnoq6
QyHSyzhRXRZVmTcN08fmoN59lm1nJjQ4jo/C/k/Ixz7VmtmzyFapuFc+T0hB
h/iOtrHW22rODMod+U/dhad1GfeiaDoKfWKqPhPcgkVpYbn9IiW92mYZw9KT
P8RGEgZK8HBE74kShdyC2Sr/kbZRwLZKCZezMjyxBb6+JIVK69Lbynt0+ez5
F7RNRjnSE06AU25YPP0NQx5ni6bRrM3qcaBtr97jFUUg3jQq5w9eqAsCpBVV
mEKCgM9Ys5CC4wPBIJgAZT2YQ41JMCqT7IsONhpU620ofcpV9YW+rx9M5Jkg
tiaQwk83g0NqQ34JCsSLwN+TOAJOJun4Oxflvo5iDggXRwI399pqBP9joWIe
P00lp10nPXM6eUEcDffWLxeMNAgF9CrrDnRGQEDFCMtr0OC1qsLtk91kGo6E
ToweoooAf66erXBEehgbTfjGOLpiTYy/JVMDDms4nOXwC9e67yOD0nUz09aX
SS8rQmxQ2BpGGlyOAW2VzmWcgx9hHyf6MHxQH4xMjMD5vHq6qA+EOt/Y88vS
57UbsEOPHS81aE4beIwR9R5UNrCxO6fAwTIcB9Pr50IoSM52iKckOP4/MNC4
DDeeYc1iVMkcZ0CeEgKJQKJwtcYn4dxD2UdsG3aR5TkHOgOlgO9sH2fa+ZAu
WxHiIldM/MaTrBjwKjrQk++MvQd2fbMTYRDP3AQL2gLHWLOP+pUHZu0fczJD
Yzb1JxXdO8lpthX+BNCcu15JBB7a6KYtAHKVcGF52JtLPCh/dowyN2WKmlhJ
da02hR0GPd9JXsZs1NoZ7rzA/aEpVHyGJEPPWlk23FtH+x5myJhUTHOhyh2Z
DeujgsxfP9lTO+Ll5geUOukCz7Nht/BckSBeLQ95mLmIMlGGJFZBIaAufXdo
Zwi64BRslfMyfTxg6fxP9aaG5tjts6lFWCd0myFwE4WOiWFLJdgEgLHT2uJn
Hd4VJAFtQF6t2lzBsigalq4rSLXkIgQaXiUx8wjfvh81Yt6i/ldquWMmTmaY
rZCesx3fIz9Ja+c98ZCaDySjnXzVTHY5vO0evb6Q+jNh/zfr1XpZy0nzjmwP
OpzcqGMW2OY7u15s5GXlhuCD5iO+pp8Ia6BkFhmSpBeywIXnBCuzYsFU1hsz
2LdLt7u/KLjc0T1KzpTVLbz0UoacWd7NkSYx4eaZlqyD2+juZWy1G4AV/+2T
0/CP1DmEMfMYFpqitlUrZ1AZfaMQxiEt0uW+gWM0pLraeBAPQic4Le1KUGMC
fWky0jIkOLVXxEmBkTwV8qfmpXfn4t161SlFGKsihUHmBFKyoNfOpN2wcQW3
cPqjtwJ7dU/IMk6AwTYGSeD4tY300I6Rxc4b9uUoG8AiqGHWQwpB42X8c4c0
g2yvFtEp72HDwMXOS6vTMUv7dzZFvzVCS+IqanRNc6ZX6URmeVkH/vEgKtPn
YhqKf4e4QvMCi/s2hEnh/cghU5Jl/f6csxRjqYU3okHiqjHMwguvMolP3cuV
QFiLwvgDr78099LPMBNpGj5JvqThmcUwjvZWqdDMTfEiiQ37092q/SNIdjgK
ev/+s/zJvOl0Y87sMBkdLcL602UTe5WWVKV8C9LS1J/FhDFz0Exz7Qbhha5N
msvQL2xFsZnMk3vniva2O005/AoElT/x+RWwkjBpKXegkZQ+G6/pgG7d89l2
SuIAbxOdWdxeYQKNuctlIOvASTal2Nmwqp954AjeRUKU+ftwPo3GjqJ3HVZl
E4KR/48LDLyMUG4//P5fURaWeQ+aJ6LFXw4V9p8VVWI7G6XCE0YlhpxoPr7w
eCRYPVyMUsjcYfaYvFB163ePbt/UgSyUY0lNIDwxca3yqLShuIt6WzdnL2pj
LyvnKAKSqa6Drzsw+iqvtnPA80TYxDcEaZrKBUOuByUvTwL79P3Lc+8Ct+GO
Ba+G5YYQC69ij/Sb3Sx3RFBXLA8QLPrvPhgmFndSwQa0l7LvnARCzs5YxAAI
DhY41x6Xo9FMTI5CJ/Lz+UcfDlYc/lb6kQwmWGh/I87MYat6P2gwMm01V+EK
Y6mPIuD2+RCwYGZsXxaiuFSG9/HaSfwttaevf6vRvxbVtZEkzt2MdyYwnRIL
BDCTdTtZzGV6u5bdM2g2wPbaBbUbbeyGROekaHzhE+XHuLq5T0bUMuVQF4Ee
lh5eBAvO8TpAvrO5P0eTgYke2YMs8h3at/1VPhglVHCyl0oiJZlJ+IgGt7zL
7ujkww5yIWdAJqMFCR/iThq3icQFDf8t2FgmQe7lTButYqHEMJCphTgxSjcc
/g/3/zS/uwjTKoopePAYoAmlQeT1sdr7xF8HwbHTh/zaVsnQJuedUHc6Xzse
ltLrWNYM98qvRXAPZhXzg4BT4Q0szZC+QzXBR1715l7axZ3GEW2aou7hWdlN
bJgfIWw2zog2f7F1Gc8W+WolLaCzSK41ZYXd7Sd8ODOOY8xcZ3eW+r+YiuKy
u0l0osIXvYrQQnEkKseV8w4rVzJSaYrNU0suuMpgt8B8V0PxGb1o05AvWt+0
2154l14kvyIa3Rxwyb9CQEAuB1TxvPWtXBl6HhsfuilUy68zT6u80cu0p5Y/
biMWvLlTbrJthm1SyrpVeuN1ibFzF1G8THaKzWHate29tYwv4bVZBxTekFes
L1hqpFPKg0I/R2fbyq6pn5uczxw67XVo8U0JB0jDPPqb/gVU8h+tLGnjnxLh
GuX4cYtV0PwxB8Xiej1VVU87VioitQTOBbw/x6ZKw7FodaJoAWzrAJj+x5CX
xh9ABM3ekQWmRNWT9abmTEPFy1Vyzto8P/M07Vi1Y7j9/jxMGAIT+kXqz3VK
+Iey+ruAIpPjROei+yx+pihxT7nLGMHmm4ZdPtsh8tQcF5FgL/lzxFeb85iD
TnMKvijdLGwbtYl3wTklIgfqaEYd0eyS1z8EZEkNnDBZO+34v6tjyx6jDIG2
LChIzDQWO9K+LEzcG49Aw0UfBYLvakT6viBEozu3Lfr/a1JQRS9MQVucTW36
dE7Dx/PHuiW6hoOuX0gbf7abbiKCIayZbtii/gZR98fWkM6GlAcLy1XcSNoz
tHc/VOeCW+5/VMpEFE9YBKvQAoThavPoRoC9jnE7qSBhjeTAKQa106aSO2QI
/85q8JVks3oS0JAMlqErEFU3eSTUUKiVRZ5mgHeUay/s2CCUjGlMgg0tJlji
hgGu4GPpZ4VJ8T3+lw9+/6g/B8JktNPNLlpm3g/Q5Qq1EkMI2IYBIvNx81zL
ITM4CG7H2df06OdgkLZXdoOc21T6fdVOP42ybu5UfFg3bFSVVe9SmD4w6d2J
2ntkPEiHp15WMS1lNsnN8y36anSMKuOYkCZekUvqnB3UfxF9iRoMFSWy02yl
rcCZ5F/7ooTrLIqcVPXUblpamqkxJ3ms0qclTCi9hMxDFc61HDJvd06Th2tE
AFFqHoIMo31yNEoZGIH64KGqBYzOVXNVOKNVf+kZXdgE78zySNO4mVPpAyLA
j3SuHBAvfd8rFgfTQdr8/eDj49+WlRWl4kEl6MN41bxZmLhUSmzR2WE/6Xhr
ZoxWwAOo2OOAP2wRUhhBvXqUXnfNM3HLONPA6xVTJcRU58NpT54ua88dqYCA
QvM1gnyRMnJ7oHXgFyC4OTtPNnxBlJmhL4QmAa2hX+dWgjiCiTNBxMp2OCm+
o5FKWaMPZ43fI5IXR3sSaiS5PlFc/mQjVr61xUyEASZk3onQ9EgAYCdun4xw
2f7ts10Gpl7q362f0fJD+vQ8Xm7uFVS7EZkG8XOKAjRrNPKcLP/s1wS29A+4
l5ELzfk9spQq1r6NMvotFc9NC8QxPAyKm+dKoByDwWdQS4fzJNOhyX43cv+r
X7BY8pkPcTB3asdeJzoGaaV1tmkN4RZDkIDQwel0ml7IIRkVRBvWSxVx8Pe8
D+dUn7bNHO8JqxmG49qhmpC4avkPDqms64ogYNw0F3mhlQeEeQwRZ/weKADK
rvy4An7t+pxoaxynSq6lfE3FvzI+yeexpfUfVyGp/AfV9hF4fENiKGq6rtml
VKvHdO36vz4Jrc7mpjR4Z9O8XwUwZLMPVIDObwh9rfL1nlmrw+v78fbWSEVp
s3D+27J4sgRrZ4v0T0cfMViH4gDc4opvOcabCoUpq4CpGdBUA9w30kabGk8F
hCZ2BIZ+JXB2J4jYYymMyDbw5dt+SWajKg9jig/YS5zCp8za3sr0dHzPXowQ
KaavOGphYlx4fBqoXtQYmaVGzf1yvK69XPLbKhy+pPMARqUi/iFJmGOoM2Mf
4nQ185BGeB/WbtClSUdJ1xMF8tDajfKVYYXlw6ATo0WmKwBP19wALdbjhdYC
43PEfzrwZp1mtb9LrWcQGDe+2FZKypHdsuRCcaXYMDvik8ocbyLH1MGotdC7
iaiUqTcPQpTw1M4MQbJqy6R+ERQ3A1jAqEteBfNoJrjByIX0vo6x2tAWMh0s
HwSDWf5xakFe8hKqHcR3GgtCgeMb1gx/auzp2tI83F8tqhennWYgkytKncH6
q2pip9n9Wu4XiJKEuH8LefIOjg/fq9ohpQ0a4vFgrFqfFSIEhw/DG6azFjgS
YSV/URsTWaDMXFl0kclIg01gUt2TuBC1+QuI+Nv7630yFWtw7rosF8eRt4+f
MSIfV4toFaVfUsvAdz64ja1eIvzIDk+FAiS/pZyJXNcRQ2C5PopIl4qt/awj
jpj3vwnpuAd+Xdun6ogtgIqzbwUinpg+jvvPj0s1m3nCOQ1tJapoCkvr8gaQ
efyM5nqXidj41pXWLIsBf+TSFLBsxsDn+s8reA3klG+Km9HamsAc4yOyK1Ku
hIeoxg2YKVSo3zGEbbeYO5g7NwTQ3ZrstSVacddWdOityRER6dzV0pOkeDJr
3vsS9tCSPt3qEC4yp6OwLvuZoqexVw7Xk4pQnD7kUjXmkCGlL/OvQ6nIcYEX
/FsbWnkEgnkp+jV5sLaxUY+qqQ6h/OL5ouWo7sZfopn3zNjNwIcnnLdsvSrU
ZoWe3xQhwxp5JjvtYEuJYrGZxojv4V6kq7R4qKeoIMFJBrvbr+41GmPWkPvK
z7a8djdkrejGd6Pe9SyOlCR+Jnlm81htBwS0+JNlrqB/8G5ADUnv1ad9L7PI
ZgnrZUjQ8pFIjKewNep8YNNODYZuItYuXYJq6XbHR7r13VKsrC9FcENsh0du
JDHqo6M/fGNVbcpiBPgXBsNIjg0ayFeFMlR9gJJScS3mrsXpNY7uKfSaXvdq
BFxKUxrrydOdl7bLPnvwMySTeFUfX72CpCBk/0KAUz0S+qEO9A9YCr8PRFa2
Wmq8/TJYoKHPDD0CJrUEcaZAWhorvf17CTT5vLOn73VLA8oPELyvK4FKZ05G
512g9o/L1GCdHOXQCfHnSjp1n0Muql1DoZa3s83ryMY5jI07aJHkZDAwCddh
4WDZzuyHS8JYsRtLV1AmpCIjEzxB5/AbHWk2GXJWb2Yhp1HsdS07C8kfkkUD
tvwGuss4rLJR1wMdrB44l0SPnEf3kfCxNmL4K4Lte/hfbhhm+yBicFoQh8k3
FUAmvRjBPRF941ZApT/LdwRbdvoY3CgHhI+2Hp+8QsK7XiIlAn2h1Fo5wbQO
aTRKEhPLDtIcSnxVq5fqwBYYvntffFcnU15mPq7Ea0j3oublcZg1tiwSoUpr
gLtyBwepcL2b5SjNpBWd3dxVXLw7C0SnF4vEKHwAojk7dYVg/1GLCokdy2wS
B89aql7uIzV7IpHZIlXAvADqp4WU+61dXtOx3vdwDM8z3E10u76HQN6m5YID
ldHxLbt5DLnxhzBq2fr1mGxDvk26hFKnFsHxnoVIFwqTZkvIOFz4xdbA2z+t
hGgXlFC/fQjQ7Usleml6tJUa4hlRK6otewccHH30+IscSIveTaKQ36xw4iQ5
/+YQ+Btb2TTzJ04a6YxNIQlndoY2Wd8djGKTNTUebYaC/S+e0FfJHHC4uRsZ
Hs4P2Epy6/8nrSRnleHgDd5ma8q8ihvzhXzjuMsGeVFa+dGTmgzNekzNfefV
fAaD1KvS+jcf2EbecyFu0zsV/HImDh7NVR76eK/xYRx7bIglLn2aYbi9oYuH
KAW4d1WLEo+vkhv0bYXVz63Z7GFHUXzyj+ubRZ5NIsVczzQrRpOXVYHoSEIB
gYi/x9py3czDcpxtZ5l/6QYXvMeAG7etHoFfkcbl/PeB8Rm6VUnnrWHhj2lu
srTqbJslKtaX1peScMuCjjHkbQ5YJmag4myOWAvnRQwAfwigSMeHNorKE08s
QKvRL0xF5LPYpqDRWFvCVseV6JXUgozJus4k6VJyPyIOB00Jx27kK+UJoM63
VkwhUm2C8ImrWeDhipch69Sa7Wfuliz7P3H869R1VDXyqANDMcO2xvQfgW2w
vPoG5zwquhldRQuV4NKNJtcqfCi5nO5IPZqLoC6yv5uhlDEBQVNgR+hq9ehL
1fRcMpiqHgQLHpPAOkVSXt5slgZuikZD1184Ryzv8Fv6fO7A5w7YEgt0bco5
4atFLEgy8LLQiE/6oX5r0yjra6l95jWFRWj4hs6SbynSGlxgbjVxS0gOzQE3
wC3Vc6rGowHZM3N1XX5Hf0wrBqfPiCM3HhLIP21+x/vdWPYS3d37C6zVoSDG
bg555qbp7RZEBRv6qiWLzwtHOlxBZ/K51qgjW9Ys8hI1vY1Xj0JfE8FPBs2t
CeM/ePFOtlw8xwTtuu9Z4CDchaXO10Ee4/y/cbK3d2rxB2R94J+O0NcyEBCJ
eU9gW8852j9iSdmxLddTSN+Kl7J3c1zuHhYv8ociHmfyFQ9Y9INws2EuLCJB
c6K9fHMCM6MXBhaRWNoGDWFHKO8TwOvB8IGQ0GAiRqYRYrHVDAU6RIUfCWSU
lKV8CMoYzXlzRcKWwAT10GN1XiJHXDm+H+UqYPit18bi1b0lTW86vxqkSXoC
RzBTmf5TbBtvAZrR4z4lDwervnm9zrD+E4S9kVSKYOghNf99QGLlLfTk6gNJ
ZWtsjti74MAJqMXmzhtw8ulZUSIS+zXh7ECtUmHw+fZMeksLpqmYozhFCXmo
Kcxfr0gGDkTmmPpt1kNUZX9EzjG8zcdGYhJdh8PBcy6sY4tpg4FwDEJQ7nZx
hdaYboTftxr1sy2bXMvwOTdkwszVrEvOQBh9jZUBm+m+GQWw6f+mcCnAIqil
0djozexsjI8i4KjcIRh0PhB2jKsYkOXslMAmIfMux4IdPKkc+4rd0iJ06cHt
RToVKzawm7haG1Piv6RpjsYTwAsDshJB7/nZYndjG+RFc9oVJgZL/qtztd8M
uyI+RsYzBEL9sHEifUtrGyoZsdnF6c4eZI09Msv/skLnfX88G22l6ZcuBspR
m8Om1ToT3JqiciU9Su/FvznzczhcmW8BYZBhnJ/gQuyRjngBpY1Fgkgzh/Vb
c0GyvFONRQey5t9/xD6tWxC9W7IUJGO/z9eCHI4ZcYJ/ig1Ayv65I5lHAPvk
9K+Tt5aXv2ygPPbIgqolJQPOZrAwvAaO8MdIjo5OE7p9FpzbMmYDFuWwp4r3
yDNynzqZBSZ0qWStI9YuO0lPdwRKXZb77Ny6iq+kgzg/8/lMGPzrr5zegnlO
p4hcJi9kU3xEE3QRotPG9Thun5bdOIkrOgqJtzYYcZluGsZbfe057sL6X9ME
fa0vNglDEKO6/+lOPcNA3ItS93REgu/+deLjPlhIgj6CqVZIih0hhcajaGM8
Ws5fK9Y3HrWRI9Dbecza29nbnOTbpz7g1xkote0mpO4vtfCjJ9OlYFZDn50R
JgDxJBAtksnwLxMX2FgvBl3ieb6yKFM9BMrrr9+4IXwC6dzy+9V60H4j8Jgo
Tc0K7CfCap/D0VDT7WAnajaALz+rTDPCt2glFGcQVo2s2BY4MkfL5ImI8H8z
LVnVZs1Icf/klihY3MBm4Fy5cDuZvNP/YLagLYQgMQWQS+I45+HsjHrY+fjp
9xkxayYXdJgAM0xfzyx35EAiJNSTQya5/0e6NI7PbQXprzR77/qT/mBHsRuh
SF4FuWdOrwbxtWsn5Flc9FLc+XfBK+pKt/hiTWAgVDF4SSHRWTJH5OqXBYAX
i5Acg2GuR8iz+4kqGzBkA+8XJ9B2sGtX4AztUz7WQMtxvNdxhV2f4fT001qO
f81BgzUFGc8YasySJTe14MjoCGilnszgmJC8FtH6LPsrglc9ibmkl2fh8dp4
0hXHl1V20mvY8yJqxd/Zmteh3pQHkwCvpEk0ANXvzxvPQMc8Ung0n6oIhKkj
qWfqKTUemdR7EZ9YQhXydPxLNpCBK64MOYfWIm7qUGbBAsDBglSmz3X/PVbN
URn5F8IOWi5JXWGCsJiMLYeQfnh+Z65agD2Ga6P5NhKDVyzvqz14BHnIFhrv
kZ/9+8iKq4IX2yWvThjaTFSvY/3894VLNFIrcEiMJ+hk89+qFtGRFJ8RyHyN
c9LQR4+WAXDIsV3BvlD0n/R6PNcCTwmThGeSHlBYSltfFKGzkfhBUjt/s6S6
foLOM+r9tMw+RGiFvwKCdOXqcznCq8P4gUj8dKsFFaDSw/XnL+AyD/QtgaNz
CXc8MnLHynaFP/0gPBhJNCf1d9Ldom4AfF3SNMbsA6nPnCjWc7foRwfW+VWO
p+1CM8oguoHnYdeHYsBldKt2KR77wn2XKOugR/12YIhvQm8eyLneh1lVxk0k
LfKvdabKoqeMp2Oc/2/GOhvAC5kUJNeIv8rovq1B6pKNQ86nrq/UY/tOVfNW
2OeMOgh/tHi0EU6MSZs2ulEiZ2wYFN/4aHHWYJCryeiNaht0jtCR7bT7ZIgs
LbjhSzqJ8OiIgbAzgQJOvabhbsnjsFVTLOsyNcxoFvTwj3at1hA5RszjDZVW
Vief/zuDZ2xIKOYvayOcmYosIo37a6oNKsRf5MRw5MtQh9xc0zApW2UiKv81
ygFvPuENCiOIe+qV5evS2uIfROWLMJSeHz5RA0GpICOV1qPTmt0WGL3tXn8y
QK5e5D82YIvps4IE/AikgpexHYmFBPIjcoEm0lP+hFjK/KbIFhcnepvmSc9O
B+vDTeT5Mb43LNFj0jJteG0YhkafA68NayBSQ0rwebLEcWnsrx8Ncm+G5yeg
9i2Xmu9GILWDq9Kpj+hqAeVT0M9JqcdHYzrgL3NBo1zGCpAbsymW2Ercxgme
wbGk+rDy93A0j5TH0V2oDdK9ixlTZz3yMKqBak9s7Kdi9G/x8+ysDjJBMVMX
+18nAm5Qwr3ftFXUoftY/11zi3xGXjnP6uLdYrT4J+WN26YJrvz5cJTpROH/
4VsBk0f6JBH/YR/EMC1mCCTIZStiM8Oh747ieQg1sdMZ/dwKPqpLXKpDNZWa
fRxRymafgoL4uSiyh+WbRRBkuD48Db8yNxXGJcPnFOPpsuRaKACnj5gPVcOb
3bd3vvRrw8IuxPbWLf1c2f11d/nHobjR8Jseh76GqUSvPDnk7C/WmRnNqiAh
OwvDpH2myPPNpRXuRfbTB+PRJtLvlTg6YqWlY48vomyXdjHXj6ltjgfAzYM4
6UFN9guzDZsygXIHgJrgzS0YX6vll5uUB+W4DLH9wPlpu6TZVcBXt33Z7alJ
Qmt+uQEBDVR0RUxVaMBq8PPtP+jHasiSiWlPU9ujBCmJxyspmFgjC4/P7eM0
d9GivBmVr0GoF83Vv4DRDFcq2TL399ph+Xav+034/osJbhcRTkIqw9YK4BID
UiT/ncpeQg70k2MdyL4wHVJQkAisezSZQ14cG84L0LWfO8uwJdboDYhnyajs
K2DSyyFlJxw2tbDCvJnwW1/qJsOO+jiPmdBJyNqW4HexFADSyNKW+keMHasy
4QwVaCbyINzb93SzvIUp3xdWuQtdrxyq16Jk4guDffv2nQPfB5XNvm4dkAbL
bqSr0q/GlbN3yhGlGjBIr8TMnBb7Y9jiuA2xqyzTv+D7FEHkhFNbpqQZwVHh
3UnO2AU8kPYZPPSb3Q8dBjTnd/myubINSFTTQuOb7BjyEJVt176QWSEhM0aI
sBP80rvPQVrwuS6Zfrh4onEZAmQ+moG1JYa3lK+yz5DnIvjjWaby0ARuiFWK
6hWREknApnf3OTzhLVJupQ3NZYYo1U5Ac61waM6vkLr24KbYpQWfzAyuSm1D
rSQretrzx6BeJEHN0sLEMs8JAyuiO195SGV1bPiCK7BWF9Txk7Ys43B9UZjf
Ct7uouTNE3QoQ+FjB11US3uSXw/P2ixxE4Ve1nvNR8hyAAlyLR5qVNYkKe8O
UCSqb8Jnco4bdutSPHt4y7VD62Fu3SfFww/5X/tCkIbB1289F36dLkGbXh3B
Lbq7AtYX6rpegbg6t9HsPDLgRcv6CmYMxrkihvHIsmDEN4NpA5dctWF2FUmx
PIIIOfeLitJm26lr4ynjamg7G7kpspIbP3RseWR1bvcRIXPX4Fwxv9m4WOuT
S4JOYIpRbFRHi040iJfbWtX8/5uALKF6H7KyVDrWXFcGKpICMlAjdsexON7H
IzURZw/IUROSKrMDtBtUJ1M7y9iBGT+fEqVsrofGGUN97Q0Vq5aqH7x2GGlD
M6W8tZxcXyyz1DM55gybVgTECuk7MHfXAKoLihkYMi0rSwfAb4kAqTQs75SH
5rCBYFkqmUPqYwfuX0SntHfUIlUPmwl5X0s/CWbMGtdfKFk8/ch+I1KjVqoh
J8biHilyIgeHBNAMZXP7tI1m8wNP7iFJDGXQiBgypLtP/mEBi3qVM3b4pjHi
Tt4aGNMNatwV677dZ/8ze2GWqI8qmILJDtx6rWhxp/sTTkfEArzS7WMhJHUW
dVhMb4ol52yWWKDwNgH9i45x748PTgbl5Dve2FOmI95PVoydk1ZP7gAkJBZT
gD1WM4fym/omjp3bkvvu0nKCBLWKIOBvSg+rjePwxdNu0VHGydVjasbXIcYG
bdJMHPQmCbcWnDLnlMFuhAJfZz8bdkDb0ZmzVjFlV9oM7qL0XpDeT2e1j54Q
08BZWrLrmEdsN0C66pzVCcwd43vd6mJX5MjFjrZ9VOtfDjULslTWiLF5U242
OWEM239bUL7QFNuZcwaanhD1S8nI1+Ocjhvgihby1dN5OV+7u2x1LZpLhaVW
p5LZMD5LQy9kcJ/Avfrc1eYzsUr+D1m97CTnwzYqqLgOhV63hVd0/sZwMTrP
HMl0ZHz+lGx3FLWyOK2csh0+c96Gj6F9n6YRTcTNNfIubj4Alq0cYkBw21et
0BQBOit95hF/iiNR3Hqb9o1+AhKUEQHDsZj2s6o4cd9CZW3jWqFtkzjUXYoa
SzJYPnWD1AX+W7+6B0elsEXk4DKU8OA4VkPwm9GgiQGZzchIXOasa806/jvf
qB3W9sFxouzS1YX3dRMPAj+ENYsAV/SCY29ihUlhpxwauYyTNkq4OODayKn2
W3DttByLRhXz8A+uix2SuW3k1KrQjL/8ey/vVNYe1TYUl4Ur2t8nXPL1mISK
MoLRk8ugZsgE4nn+C9MaDUC5+vLgj5Ng3wVav0EqO8zje9CK0TZfA/tnq+jH
nsgGjvSKfKwWcC0m3WPNvk4FxbPflRxRWnF1u/JvK7Lh8Pu/TSxkEgziyZay
JkvHtB8y5E8RHZV2vDuUVaFBHofnKLPndFlCza7rOrtSSd6iZfw8SIl/E49j
fnLzuIewsIpy/ToE5JtgFlhiMqXu2jbx4igzPTXqjxl6MpTS1S3zdHWTkute
G1mXXmjUgEIuEo3UHHmZiHhBJennsrNL+ju1BAzhNod+eQP5yJjw+xoGaNOO
BKrj5vxp3xajxhw/6CMwM2bwUIwAiPsAtKjlr70pL/8rTvChR+Q5FgvATtlP
9DLtJtnjeSmQ9iQmisxx/lYDoNLp0fS3OvaacMBPZHaE8JzBizMeGpBKQtzv
B5I3sbJCAfG7Am/5NK/qtr+YsoMbAQCUUk6kxe6Wpbz1mi7VqJKNL12JBulu
f7uobCXxQgS/PNXad4htS5rL9rwNaNYGY6hFnAeUQIyA2AWFtjwg6i2IQFhQ
vhT2zAy4B/ZFMrzGVAyw0ct3D6TeOXAmXqpy40KHVC9eaoicC3WE+kHebDuD
NbZHrll7kqozzzV7HbRmfBOiRpWakvc/2HUMNqZbxNBtrXQ3vma+BFioPF/p
puvjhXkd5KaCgdS2yBWHQiQcuORUAbNxB9EpTe8tLh6W6V2cN9u1M9x4cODv
Vqzsq5sQQbhZUawtu3xqMO9Ni1Ke+th0MehO8RlS2y1goUGprx6NvFYX0bPA
9ySHDeVQBEwp/LRLQEurjhFvVVpwPKMu7aWcYbVIkPCx1cMMh76+28oLdItH
756XHcmIUkcjD4b5wFJagtU9rUzksbPQBWGFgPVASAYS/Fbt9XMzY/J7ND1b
CZdXltc/TUxi6rarUwXDCpRfK1ih7Pvb8txjZP1HpubZyUW9cReZpm3wqftf
6fqihKd0ecOatVId5vDW4mtqswf2nPe4RIfqEd1L6DvznTcciWFA7U8NF4F3
7AKZ0b9qmYX0vuaZCFpWvnpf5FJl04LRL+ocHgAdS5NiRQ2TiwvS1LXLC3rd
5zredxNl2EjzhCStjSf5DlEbJ07VNO25k4vyxF4qPDkGKaunvRJ620O2syTH
9o++dyM+lE6ZK0PDNBwBDUJl9xZ31gdm5vvfjYeAWANaJ22k0MY5ov+LJvMR
j/eqHE9H858QbMOAuVmji60SzMBXTgnDq8SUcz5s0QC0Mqs1iBh2wPGJm/H+
rJ52kgtB8/1kgZHMi/yHcvVsnFIesV6D1ecdu7WKPQXTcGwyoOZKy2rwe754
3O06D09oBrECb5AnsCzkvQVXBpGhcJexhrfy95660kH8YsP7q3TCfyMp4f8F
+g2DoaX8Y6QyUyACBsuxUxo5nw/ao2+I8BoH3xFfsLGWjLVJQJOxRmSuQ8ei
wjRfDjrBctItWSPmGuwD5BJlgkp5GO2rQbbdqICaCM6PDwQGIFOaTI185g49
FtlDQBaOdyiyNXsN04aOzJOy/2R0Cc20hSuTrqaH0q1GHtm/oQisa6o/KAZe
R966CqhwsYeJNpRf7VqLKO3lpMaQbn5Qs+iHusWlYvzdpDIqelQGTFoOFINo
HEzD+jEjKuptsq7mbjwOtk+Tq7qGi+BIBHE8ebbRNIhUAIt1cXKBsLh1ksra
N0cWuhSR8im1rq+kcy7at3AlgSTH07hhLEsFg7jqNjxgIysvaG14GcSAvwWs
No0+5+0JDL/1Mq7BPRDt8xgk3xuS13lELBbXsziziMGcRgaBNXpvIzKV1uua
ac9yEq2HWD+iUVx/MoZw5q5TGdNB5LqigNC5hifpC+DTGU7YEU+32ZhC6/m/
+Wx5FWFk7+loudpFqk27lV591uBNdXYkMeV7AYUOxdKypoy3zLv9JCc47wXl
odXw2fooyaX3wSJlA25XZxacuTGlR0PPoFeYYgd7ThSqoaaeqSQGKRwgUOI8
SSISzSG8cI765bUZW6ZOpF3RJl3Uyvp2DfUWMwZIRP8VbPTwCMGLIBBHorxN
IkuY03fw6I6MUjykVzS0Zw9z2qw5lHf1gxXuAd2XqoD9JWQ5RRYhiW+QUBnv
ZRfjpr4jJVjx/3Je85TF8DGOW6d9HNMyqNwHzP6v6J9T1/x578fjiapLwukx
Zs8wX2hl++1PYEsyTQ8zJQsXt3hP07QBaD2K7B4BT0eSir1uaUnFb2uQUFvf
8zDLX/EKWBHpIqnFJa30czvLxDHaiqTWMH2Gf3zRJRNJCPYbRS9wLkhHb1Xa
ZtcoZ37S4r3ISP6LMLMZcxyoIwbR5XC17abDEnYi0W6sFb6gLT6VDXy92IPZ
cCYp5Iq+sNDpOx+srmTaIHuILi8+ZKx61sYAt0A6GOCJOjw7mDgiHb9EGyIW
hiiIbD883tG6DwFiU2zi9PykvZrq1JGTstVgxAwcIivEKdxeC+WY5OthJrB6
yQGI6vkcsFUfLFTck6qUuUHwYXroVCor/KKORm2h4SMKktrt/aqN0LtI669o
IfRz6g/l4jCpPfDBNlsAp2JrFdrGSGKZ1B5mjTHRjgSbGP3FEkxLiJdeWx2N
tV/D+dpVbN2+YWppzlNIHtZk+PiieObZawl+6cmN3AXKq8tZ/lK0HgbYPEj2
/GJs0mszflxf/ZAzSvsnlMk7typgjhYCgtwrxO+EEx/RZQ9RF+aqBRH7iOpy
gwGvulxjsTNo+/5u7gbrmCWleduW77Rq3DFngqac5tThPyjNmxMr5ZIQUmXQ
Lj6FAFg+VGBOW08zB2p6145uomwTTZfm6HabhcB74aCCrZwEADNAigAsZZUi
g0MHIPyh3HyJD2/wHrTZP5JsJOvBCCGH51BKZjZ7ea4uPw7LzxxeswJSj9Qi
fEypeaLxo/4+SH4o1vU30MiDMmn6bbmgfV7ZOQ3vRljk3tMNG9uKGn13r+s8
RIX47ekDMZXaZejWehqZbPp4nJ8Qw1G4sZwTfRcWMnIHN2CfhbjE5oF6UCWS
a35+qJ1KPx0xX84lLvRKP2bGhuzvG0XiOq/CxoB4d1oqfvRaeRYlVTPZnTy2
D8nEXgQtWhuPBkunuXgkQz5E3BSpLDn8aiZ/FwpCBg+VBJd5mI+BTdOOjkyC
XsSgCRRyygfm2yNk8Rdw+yYPPD0D/vAw1xGvH6dCCjAvJ7hlZ2JeutY0Bn7x
Cvki/7nejIqPytNNO3TGvoo5p/ZZ84bSSEQ7Xszlxy+H8i+Zk2oLB2vUN722
s4nbsfI5kkTsNTtsSHaVHMcwFeWZbrRg/4elIbJobJR67srHwE5hhjvWxWCi
Ir2f1GT1Jl9wblrKzd4riIPbz5r6Q9J/8len0LIb2CBl5KJYjsvbCiZzvaKd
AgEzJDZ/KPEErVN8q3C3fOvhdHOca3o8tJyj6/Hu0nINxsEk1at9sAiR2J2W
QGia2jnuvqRb6Ya0/N0lK8DGFG/UeKdgOQv6iV2bLGHEuF0lIFzNEyflkGJX
wsRksAfcaSZO2c6TeCybNs2Y1YB4ZiZ9KSA5Eu9aQUBu3NZuImBfGe6IKATz
JiVars5ITuWx/QlpH7VCF5Bimw63n7lgk7Twy6nJU5D/dMutP4jyPN/PVK9w
qduFa8+KCGyVZruFXQ3xtSipVA4SxF/F5jLdcBo8YyUJfazZmEfqq8TCm81F
lKZSG1VUu+9ElLR0V6W4X1vRnrhzz7uzwiac7EPIZoHrKbB33TOIX0gsHOiR
UTQDfhzqDy7PylPUWHKu8dkSaLhVoq/IFU+azlIivvHv3vw5CymDSaIhdBEr
vR7n/W3a5rXFx26dof5ONHqt16Jf0BHPEfY+vrr5bNLmogi1COgqGtNl7Abj
lv0P6vv1lBe5ujtIVMWK2aryzHEZyTIOAGsKv6Axmdl5dX/3Y5F2gE+FNQUP
IiiZMNapHHFJ/DGlPjbwuQgw8ANz32Cdjv0pYt8TdqCirxqWXHGGYAZOXH9x
lBP8UprXVpJRzGKGYWW1dWhMspRt8JLqeuTnRbf2Z09WIAWYBRmeax9Ihj1F
SX2RY6uLcmxVSTSjLn3xlVMlkBtgBgsL3JnFPhDggAafBkiZyEKyD3UDIsd+
IyRyG8DWnc00KmmlQp149UfZGUHKgx5kFqiF4COmDaMPSP3v4aVtKWvUukpf
Ig0L97PRXuprVQazuur0jHwyAYmMBX7XzPAHTxYU2JMbw76SLTTXCDNlYNj3
8Rt5ShTMWC5RL6o0xQc6rRNNFAlt0hsOuYAbvK2eJ3ORAjbt65+Sb/2Ib6Rl
9L/IfezRNmNZVa2ByCKNm4IaAQXYQrkwm7lGp9YbEhwWjH7ilZH8Kjae4m9x
V7/ELbDxtBM2s6KUkqJ9PMj2Cmh57BGZvuP8mX02gUllFBkbw8JexUwu7HkM
DKqsBY7FhWHg9aqj1xqDXRlQOJJa5ZJ6ldb19HDCu/YGDkA0gbMkki00eomX
w/CDVN/Sz68QaY3uaUBy2wVI0ASzJ7whYCRMjpBA9u6GeN7xGce3Oujgj7RF
xk313FehoH7A28TtoJ9tFyxJdEiqGW3N51JSnIym45cUVAzVIBOAnMyq0vLS
Xn88YQmsAggOeF259no6jcXuzjTRsXCigBeEBrM6L2xvUp1QgEHoLxbtZdRQ
w6nlWomuNabBmTG+bSFG1wzaat+Ij0TBzJZqB/Q4C3Ih4EFsB7gjWNEYAZsD
rYTybCXYrHemQj6qud4u2o7YzZgfqCCvOkKnocDGxeCbkgOE82gwhlWAZmBX
Vc5tc4Q0NDyTY+o1MJVmdgyaT0xwXCG1e2qzte/uEDxNzIr6cxLQ5i7+cRap
E+d5pa+FeJLgacdHq4/yEJH2vyX8ExUxC2NcBbSMfBzoZZzn0+OuIblSpBuf
R4NGJRQX+mxreR3FO6EPhPdiAVW0c0LnanAcXFYRXvgrgIwTltsw72H13O2j
t7JdJN/5nTI9OAiGv8nhJHUVA5hbpJyw/gGFo8K4/BKpZBr+5eASfuaGLdtz
EzBs8aljSezirm71anqJVun6FZ88Fdj1tGuU2/lZn/TKueAmrjN1uCa+8Vsj
lU/2tpa5FkjrdNjIkppAgEL6ondKlehJKur1ortHVAxQjTNPCIdPiN6o1S2F
GepCdV4aK/j493stds/G0CNJ2enKfMQ6wfhVqzzLq+Xuwb82cHvHg4rBZEjn
8icu2kcnPXWfFpM3afMisdw5HzW1ncRu7PbdSv6Aq3UG4nI7orLqR+J7zDvo
G4Nj3ZgdgWLkQ2P14UejBbN5MrRhONK1r7m+4/wUph78HMbaJHsWIuZJHoBh
4ncX4hCl9obRTBrVaS7XF5pCvFT7wiagFzXBXyKn4xdsqSAHxZPgTDyUk5Tg
MOXaOIPy43ZMR4U+4AwEv4AdDKK2Gz18dy5C04S85Hjk9hFPrq3Tt8K0Y64F
GXBBdUWsSvPEqU1XD1Iu2LQ7Rl3xnd61Ngb0M9kfRtI4z7ZyNBMTZsA+9CQN
Am8oKRSN8PnvFH2LN1Que2WZGagYVLXbRBg9YPsShEuPNUQYmN3lzafo+lbF
DEZZ2P8gvZSeSIHN2n1DVxcqnEmIaSHu6FQfgrgu9hS6mUhRguxHVeTli0KC
HknfRBFcpwGNuYCY/lm1Q8h1e8Emu4zZfhp8d+gNYhBt1jf8ZA03GLIexEMk
IXcuqcJySiqhZbFiFz/ClRRp9KmG3vV8mRH74x8OwDPtSImnuZ9WWrk0BwnP
TP+e5aKdzNkxooxkx1t8/tPu6HgadOqG7XuGa4GDSWkxkkBrnUV2KoeII3Wg
n7OQPfEg0MSVZgosEnSEb4aEMtoj0iXatCaPIO7+76JREqwpW7bj4EU1Cjbm
v6qYxbKNuQS7JgZ/DDQgXvWb/eZKHibUX7noNQ2UPGHWkkPsVY9PG4A0vSvc
BpneRD6k+wZAlRy3t0cR8Z3QND6noAkTumIN7f+IJs3P2nn5NAUUATt/7yRS
RFbkuklunvuO1/LDimVnWvpiJxiHac9f5hHDuxM+ss8sr/WCx50c9pVXf7BA
fuo3D83BVhEMTjZX0jlS2LuiGKY7JkKlSIUNs9FywM6qyV09zR2mapzdAkuc
83h06qq5pHG2IcQuQT/r9WgcHmqtP1lu2AjM9ajCSIiYtF+KsNdTGMqNtQ1+
f/XTBtqqMMSHSIyArW2r3L7eiXkPdPj87+g9V1LNpc9owfh3g1Rq/BdQRbuu
DYhgZsZNEZfOd2MDcDEW86Q8v7Cg0p+SwiHkqNnSFhslHfWWqtZTHFPagE94
s9x3bEm+9vE1FB8ETT64kGoXHEF6hr+bY6x/Stub28zyFlBd4AOf53NJjrWV
RQ1r24dwhA2cMW9q5cm+NRbx/e5/4KCHJBLYDh6T5B+j8y1qi8Ml1ihmAdPB
BvpKv2EACCPio+DpPt5ovyxVNE7RHEFGqW5S58mghkzv7T0/ByDEciHI1E6e
83kW4YLPQ6RWHdNYOoorapyOmRLqTn2sZSAlzzVPKGT4UhlS+kMkXZBmsGI6
JXker+fRDStg12fw8ED/XT795hnJvSdRKkaAKgvQeEykE4jOMb2P0B0F+CdJ
XPuSDKWwScP5zTv+U8Xtj910MvFELvyEFi4RBkL9sxB6+RGMkblGq4eGvM2z
VdCKdVaUj9I3ZF/NkMsOM+5T2nvK6u2AcNOfDdUfAmZvD4Nkdecm7tpo17Ur
MwxUzDRye1zFcI3eWsWFJ/e9x7PB8i1sDCw01BTwdS2A4ZhrSZYjZju6KwyQ
p/1ycIbFfSyM3/zXmMX85jz0dZsnNclChcgYlvvd01erBWNfDEUWo287eUuL
iFa6ECn/xXEye3zoEGRme2QlksYBbpkj+bc45TpzB0Z6Kyqb6a+HTZo9rVod
tRjaltSNCO3jvt9Qv+b2/nmES2gcBxhOWXuSYNYwdFLDIURAPAmW6tmpkRrw
UKqSREwiawIgIXjBqHyuMJ6WTjlybg35RQ+1Hb3r/d1fNjC/RkAjNxZrArPL
et4eLj+bg3gUg8iQxPyi9sxw6iBqNw5OdCIaJvJOkN+P2zuNpV3htkqhO8SN
OF6bScu9fi0zYBJZVZQ6p8Dj1dVXL8AWG8ruPygI/AJU8lJbIMI5pcnea0GH
0H+OrXLAIrRLMal5zSNKZhFYyTfrvn6MMrR79uGUvR1FoRYFMkC6vDMG6NQZ
mVqeSXr2+xZ5W5sOyhBbG0ct+6hvNL/GsCluAoCfHoC89+IrzGCmTX0elfar
vPj79wxKloW0NYaZLY+APkHzVs+UU1MY5lCzP68IfdAqD5uW694UHsF+MmZ6
Wd7eTvSvlnpp5Ii025xR4/PHdETvsVCuOrXSVZLKkOr5DMwnBYvqdK0GRUID
mHsz3M9je3pdS9c3u7yNCOV9cwAvHTXfeIyL4NJAt61pCaKhbqjK1qwJ+wXz
apSc5wUQPNPsiHRHR3dZMgCz7lnMx6kW9/SYgDAUJ41mFBEe4wxKXhkBZAct
CsJbQuA+mdxnV6kEHOJ/tNaMjqN9kvZDGnMEA2gl+5XFDGcgvnNId/CA74Yx
NXeJLlzbtP2eSHAIFjH/oOBJg0qMEDxreHmhv1dlm20vC/RkQIkT2dxtmoWv
njcFemaM5lny8//mFquMyfAFBD/05hSIyhXxuaiEVjyj3aDTomX5ve3B0I/y
miJhgJpSvhw2i/90Kq6pwAYVb2DS6kRDdIMk9vX4ZQXu/Spo/UWTIJxGM6xo
/2npmv/MlgQ15z1ed6vtICdgpzxshuFO9kFDt0vWQN6EfnMOyoYYmxtgi/Yp
XOsLqredX+fXszI3amMU2WIn2wYDYOB9cYr7Ec2VntAAoKq2Dm/AcsjLYYjS
ski/OcTlrSJse0sbH9nprIlq29xpo46lnmzasue55+1AnYHL36CuNdP8cck1
qMStOywrzuuiYIaZE26xm4o++5udy8cz0oNX/mJ5ZiJyBa90hZ2XbDZ8w8cA
lef3YTfgqexYICo3OxY8/UsXznNmnWK+51NWIU9kdJmsjzKmtw3c66Cx5WYW
hywrtYGVrRY0K4U27LcXOyneWyYyAT+Akw/3FY7wZlLEfhI94oCnuBTG/HBm
Q6rrHNiY1H7Asn94sXf1eYjzQ9Cydl7Hsujdpwb7FGZHBTpO5vahJ9heWDRP
Yq+1SqDCg3ITMBzqzduAhSDq3WwdOMIPJwaHgP6snChTVX4GYGDs5u1bglX7
5T24dsguta//C3zRum8ZLh1XY5pWs2Dv+PxilnEmxa8Z37g5iCiDkUVPt06X
FVifHwa0JGtgoK+Cb3+kml+7isTPBtcQKoqycSyN1i/WI/KefTOWTxZ+cOxW
gfU0dMyYvGokKkqkNdMKTj6aZeiVhiU8Pvzj+UW728Yv2UD7Xsjyk7pbq146
dc9vkPxP93txzbv0FVWjQrlrLKwD013WmyH6rLKC+VoO2LHZQphdsTB+dkFp
QWw7/OhDhzOGeeUzsXFprPbZxxQpJqusXnEQ4fvfI7jVp4p56gQCpoYWLb4h
gUrNes5IQVApyOyV+gpIlcUn5LJN1iBQJ1dNT4tOJOH71euhOpf6TurUoOoX
ZVchQYWWvAcTGL1oxPUrJYlxLGNPUcvPbObICs6wE4NZkf+q0+svmVoHupS1
PSauvfEIGnaH/RplrVeys/eMKZ674tKRz11bTnLp4yJkPB94a+ed3V97e6XY
c8K/RUZkwItZbXEG+bLfLiTf6eCgE1ll8ixP0oaiejZlHq1tCpwOkT2w2N8g
FE3AVdVh69ZsWGfMCV8lRcQ14hvB5M840azVH1t0VoAKaJ06k79E267icvMY
gg3GREn5P2AoJ5V8TohGZeaeGUJ4ESQNJEVg617US+zMRYu4isdbnzO3Ofo3
TDqyWLT1z4osWTvr4VA1hb5ynvQ9piUnPkDM+OBxEC1m3/O2ARLx1mjdIbxW
s/YuP+x6wexOUb8MVp8ABd/Eu9ACSpswjxJy1e8e8VTDhER+W1bQoIvwze2P
M1k9d6XlF2QkcQkGEQK3Bp/i4o4I5Esrhq7K52dUbKepB1a25fg/e79ABofv
Ge/gCq7TLHZ1N1H5auNtwElVJU7cqq9kK/HrN4PE9C8YR+ee4WmfHDsoyjlM
xwDty6y9YszXSfm5QCwqUXF2+Z4mKeFt/nxjbgX6+g6os6RIkP6lUrW0UtjL
xgpYOOFr/QMD8+UL0X5wJn15PQi8TGm/Vc3W1Cy1LsTdQmxn1GMLWLV/BwKr
PRfHK3NR605N63nly7ORm5tEkuQ/4cfyqG58aO0t3qd09YKZG7JfWdDnhQFO
euPLsk0BbbIqO95bZy4bhpDH7GiS8q6QUZYN6y3yGmuQsJVblQudoy7eBAsT
/MDaEQiJxTtGuJWu5a0F8sV+9LWufzd6NdM9GX4EpbRYnVGo3PzDERKjI6ER
b/mkXfdf6RPRFsD7dsDBPlj6BARCE8dEQ1RA4esuFlmnOxmN04/IKrm9rweW
pEjFoEmcvkcTjUPpwQ1KIfcIZJUOkqUKMCj7jOCVWUd3VMpTi7e7Urx5e+cC
buY0LAW1NSd5tFaaWq8SdU3sNlLc3OMAkKh5JQRDblnDHBjdYUCAsyXSHSrD
iJCIOj8fmk4CqnOxql+QPeIMPsN0jniVB8raE3QmKTbByPoTr/9MFFcqmWi0
S5ZnvmQwLQiaTVuu/LtCh8V8WWdUmHUBXhJ0MxfztpDLXxY9AxsFayL3Y9p5
QCoMPmhBUGvLTQcYhRYPEFZuzhLVmvLijwGsmucwH3F4wuqW7DxhKg+fOwE2
MAh0aT+maeTstPYqRxD4vH5+xBog0uP+WnIUySN6zjZLzXg5YKRqJSCMDMm7
CrKWhc10yu8d0Ms30ERA8OnAEBu8k1i1kdOppEuz+tPcZ9hefSQCHLDFNMfN
W8IPrb1+1M2t3uXcMyi1M1SHzLGK7Pc1rjA2G7yoVDWLc6tmZK+8/MAgaWqb
2U6ADrWb5Fhj6EC5Eosuxv0A14CtJm9TbosKKSxvdqqICRu9VFmAsT5JWTt+
ujh4hD3Y6eHbTrI0BP/q3VGeNd1U084N07VzMI1WU8suoo7OtdxkJZWQNmk3
dyDu+BVpv9v6HI8Qdu/xZHi4Y7P7hilR/+9/CYjRZxkeaIM/46Qgz46zxJul
+FwmQOWAcaq6n7wAnrY0oUsMgQ+uqSri69VD/IvbFr/hdSThY7/RM6qLsEWr
hqm8tl91FJtu26r488uoSREGmYfjmI1gvOSkQqnSWwAq7EmwBfc+ZbTh8FIK
OBko+V9DLm0fAm6MMhCINuVMtRMybHKHlUJbi63kw3G6aQfb1jTZUzTcM2c4
VuSTEV32rC41HYiBVXFgzcwImJk8j9AMvEP2ARjgSGLqCqjC+alEg6LmLn82
H90F28KjGwozAVnJIBDwsA+7mZqDo2c87RmWedy0WWmWKlxDbIkRcOGDo81d
YV0oGNKKJPvkO7cm90hJLL+wgONVTs/dN0IPaLvefi7snvEE2fWq+i7Gzfv2
kL6VAouRO3SPo5NGo8g3KEhm390XAoVeM9LRAMrgmsTKOqGtvLIvaoBiIQx3
s9CtnmRl6izAgB5xS+s3MbifDZyUPyHmw3qL0ycdbWq4hTz8Q0orebWIWVZQ
II5itaAyp+6kYOMsEgyGyVMubdMc7RpMIbQ3uk5H7REihES67pPyfbxAdLYg
EHyQ9PusEk9esnOS0L/QE0fyrNaZgMH9CCLCb07IAwLMBpZYl9KSA3L2rTb1
97yRUMinbfKuHR0fvl+cfpTRLH70CI5Rm8PmM0Wn3xuGgsAHg12noej0CpFZ
KVnjV46anXc8l7KX1UdEJnVRQ6iC1vYe0j6hrXJZ9KQUqZYLSIUxyBx9jJm0
JDt41J43wJIH7T2d991nZvnxzkaW4/+kVT4j2D2FJxsfpGN9piBf9chwMPuo
1GmX2LMbn9fY5nBRI6KwpBu0lxoKaJLSlA06TBnTNNKsut0dziUmN+8mkzVD
iZmSGcjNwlKTW6STd+E+8c3CH+35TjzWxwpNECrsJ1NhkoxQydqlFynDCUIO
QKV2qzD9ZQxcnr++FxUAZQlvcA13FJWk3cHl1bU8f+hG3wwyG7LTMEsYh8Gb
Eh0H+N9Y8HQIlgg3zLVyqd8iavjdToMsGHl+yH7u0iMHbud47oD8sypcRqCA
/535JQCAUjxXiYNvBqfH+YrwUPLZP7wgn3Dc1q4mmevTa67UNq8ZIFTAHue2
vvBtcIltwhnoUC9PcdVobM29R4qV4c3LmBGYqKyB0Mo3HLLMAVsSxf9g0Mnt
5mY9GKn0i5yrKse0Z/1GS5qIJeco0LRuDW3POHEzguzxQ6KIJnyk/wLoU4YN
p2v0IxtLANPOz0EUK0eU8WMxEC3Rks7v18QY3t1qhHLjndti8GceXVlTS1l7
/WB/xeVIPid/nN5ASDG/LPxpwwrLjYDfLrENR9l40qhTHVz5EkpZN2SHrKtn
Y9N07TRcyWJun4D5ZYgcmmVQ7UIcV0fRsTrsZAdNuGRZvcG1P0lt+9yXcvE2
JVG3YvW+ZJyD8NqF91vK6AEYCF1Q2CEmWX7iFOMZvT/ESsa7j0SFarWONGaS
UXFMDMS8cx8xRpKksWvrzovQICF1Rt5z7pa+jFlUqhsVikg9ybhVc8gYd+qr
ChBqAwcXNkMXXm9T+7TWodtewUTiehmEXd+StfQjd4iSWFKCd5TCZUjko1wS
Kw2ttjtZEtxxDUvfIzrdHx5xy4ZBN7u4ed9YBuyX8ArLT5aCq/0o5RWJWYyO
LqYFUPBPs9xnCZ9xg+NZ1kEVywNPdSoZi3OdffBiUbqUqkpH40wM4NTmKduU
3VizSBRJ66UzMP5F0aFsP7mWV16pt+aNCi7LWg7VSngJkVoHVWUEzKPWaXSu
rL49XRP4qZFKlj2BLpFq/iH0jY4INRjMf3Dtn7GGL1Tesi8MPV1aoiCle0NM
3TiCalrE35g6tL3E1WM7KebBDpwvoi9d2vtlauLq2Uj0lvJgaDF7+R1zYZ4E
mfoo5A2es1hJxrAyyq0B9UKOX/KNHKsH+otHH57cwjF2oFlrepJ753BZPYhO
PYtlBV4D2XVnP2Wes5w2MSTIbov2pPbCe12fgZfFpefhbWoWb5NPX7wjBQbx
mXQN7HO/N3MOJ+Ey20XQvKcX9Fwy7Dc2HkFDdFIA+eC6Wn03D6RkeAW+kHxW
lhRNNOkLvQwbTWLFGu8idUZKbVJ4P4SBFNqfHRChFnYL38EKhIrW2ozW1dAn
1miqAvfT7mtsv+L9rhz5aAi73UDvVq4VcEqh+KARURwqgVZkOvnGDu4Q7yqu
YDmOr1oCIeHPpooa6h+66y+meC+pGQelVeBtWLq6SG9rEtl+l91HmnC6wOuz
LxfpdPUKPBFdsyDxDuizaNRDEZGcg98xw3Fl3CpcUI//SbCkbI8MYgDFM92H
Jns+1Wj9Z8GtRf9JFQPvYsdRdtVoJzKNadDw5hxObacZumxEAKRaCXwS11fz
+tU3gB9l2Zgn647Dq8PSnxiKHTZk7Uk2rbZjM/NT8mR/1Kn+0kDG3zPXhOHr
0o7Ma8cJdA0VFYwuz55TFdHZAkWA0dmO6BK4PHABt4pchMjPtafWpLVSh1NC
Y7K9cuoRDjOQUTdlsip1okcDNWjr6vRInmmPb8xQxUyNvpVLIxYpckdrK/fA
09J6TkBXqGS4GPBUdtDJbXVF0ZF79az9FsgewJc5LcoHOgVEQhzpDLFq/MOS
9CR4nNO3UtHxVHUJGSP4wBCAybS96PFBqaih/zwNoepWKfZeePTbkLnvg6mo
cXQRevQB2vttClJVcGhO+x4jzSbVZDhgIbZMCQevNqYtaXYGlIzUkbc6fr0G
aoTRC3dZzTsEbJUrCSctKzvJIg5X82wtiodF2vRVFbM/wl56qjUcuQC0iety
QfhoHGEHp0dWNbe5DWvJoN1AIXjiOUQ4XavHRclb+STqBambW+LTthKBibel
b0gJNQ2gVKIHgktnhq0gtRxI5DPBO6uUjZN8QiWK+w/3Ysju4koZwf3fYI8w
wHCOCJ6hfkOOw65ItM+lBECbY/SiW4cl6wNjDgBCWLH/OyZCLMBoIt5oEeBy
eTf2/monldDJst9bIcB/kXrfba522osuzam7s0pk2k7mtx7kRx1YMmsysk/6
ZQqkWODpl4vStPOlTDi1nApCgeSSe+lhGGsrIAvkCrkiPWddvEmvDwWxMBri
5q0YSf9KU7EcnZZtAP0aw91XBzzf2NIsHJtDbw2PE4A4/pe4Um+p21jA4ihC
rh0PTWGrH6bUYrVbszntKr0J4El9yctDlSOnKCxr9GPd1hyBXIEZXPBRJ5BN
xvUUdzigIgaJq96haUmbdLgOvq5IWGBMQ2MHZrjVEcTT828XFDqWuBl3lJ0G
k12di6mHTzqII/7qeQ29a0vTtxrPuuI2LZ8NVIShWHqbgOrkNkoWWbVELTgU
8s+mnc735qkmFrERtUj2/JTIfKLVY8Iz82TaAbJDWNdtTaXyETXcib555hiX
dxYbz/HslgVIL71N33WWLk30av+nK970/quuXXuT1LOfyoxC2mSN5up9KMGP
Ta6jyMEnAYaIxkg/wnZaBYXipBMxFS+cYrDczj4MoUV8ZdBmbNINT55GRtSv
XFPtAPYpl7hCEgMBOhp3qWKeZMcXVXEGuLv6h+QUXVUwZBytGcEqV7SxIT/2
D30LVS3vpPQEtP+TDEF52VyiUA97HJOBfg2uM6C0of70G6Oo8ND7803m3XtN
MjBTUHwNBSOfmvW6ytxycGgDd52uLejsennCPxYHPgBG6F1RU67NejAyB5FW
zHGdpJCatXiTlkxufUp/Lh4jJiPuUzwV7MVNoxrk7FBn+TB0CiZxpjoy/EEY
Q2GApRh6uov25p4a1PcyZEzIxqg8jI3Mh6oAlJ9gXdhANLTwusJdt+UzFWJm
xxhMY8VcxELaRodsMOQlW0mAaODD/+i/zuiRwhz4IN5Ve0j1EVYBD1x19M8o
0Uva6d0+XAemMw5aSeNXAM4vSY+2BOzLxnXDvi/W3s4att4oXq6HMGIPdcdG
LCBqqdddjsCbay8VCsV4fBXbu8FQs0HXLQOzALaTGdqQwFNuS9Z7vPHriCfQ
MhABeBOn0Sgvoyvpik7hgm/BoCK8zlttpCgDt8ExI+9tsQQyudxUXWfEplsO
L9vagb39DslJIjRynqYGrdcClT3KCBWm+q+5L8J8CavpdljjpmX06fgCyx3n
Mb5xMjvju7HSpWwh9GRbR2gb7F2wxCATS/8MriFRiU1kvUAOpUo+Jpl7eReR
7+ve7ebH9IuPtsQZmDtFGCX8Hmpz30WlcGLl4wSaZnNtHRRoRTAfZ9pI8k2k
X6sPX54s2wFocf4rSYVAlaWPY2IFZ2/B9gLvMt2M062FPW0awx+6FTEU4lvM
EOSTLqwGgq99XI9JzdOsTqk+6WRFnBmmvyh8xsmgeLncKKs6oHS9uJjK+M1f
nSEXW3K8BDIy7tfEou38i9lyR5LDhpJgYuMYjNCzArICxjooRvmhs2eJNlE4
aZSBZYU9tKa9QUxKwj/pesijctK/WuNa85W0wtRivVPAoCj/RRCJy1+3bh2t
/Go9jPS78H8Ku55pMmupxeSZGAPpf4E6IG9+wnXBrwJ95CQN4OMv7h+so6kD
k8LYqz3JsGZLRkIAG9nDMDdn6tolE113lSnbl0+UYhXlK6H00u9U5skIGvUe
uYdH41pv0phrPabfOezhjoDoWMiwB9Q/DGHCHsrPISvV1D6/pgfZAH/rVOxs
12zs1oltxceR+6JF9arK5e5KcfG14YiAUSy1fa/AM3nbhuP53voRCFP6iQPL
68/wWeC0464K5pZxFGSxdgs5ZshDKi9qXMDNlGrl1JuHdQBc6kAT9N3QuAT8
i1EEEZNw1bKU0iHEeGBwna8r9ZCblnCAGOr+iJk+viug6o95Zit7K8U+tDCo
Y2Mb8Cb/KAiHjeVTzUX1D9hp3eOIRqye38BQxLxE/PPk88Z8qkoaoaeY0C9e
IU8syQBTxmKRoPeKo3Z7gXbMFbgVo/AXtSS8mWDZCIOGP9VF930EZciDevde
ar+51EKJycqHdxpmUT4IyafTKzw+SYHitamJNIRdpSmLdeb4+ep72jPtBbGb
ikNWSoKUSTDKybUGMPr9AMAxdEbrWzH37SKy+UknsEq6u+Lc/SYECUeyvVu9
X4qmpfnLD5fVw1c6QaVaVdEeHd185Fx32zHlaYPNNUQPFv2UlKGCl2jw3okh
gjOQfaWWtXwo82p60yBKj7SjM6IswlzDpCm3mr9AvWe/zT6F6P6DR8Sx1fDy
4AVwlLiNIaw07ZBVJJYd1ZPzBgUM6oCIM4I7SWM5vQP8X3OcB6QXw23pvXhK
rzAj/i887XN74/JLQPlu90UHwdWzVpE4bGuLP3FPKhG3bKngc2g5gOUh3CTm
ZHrefz1N8HtXHhoDXuGnauvS3FhZvwq8OL4/YkBD6+pQddhkEUTGGa67uSUe
LWv22i/Uj1v3cmjZCf+veiOcepm0LiaPcY37UNnySPiWd/oqxsXwZu9funwZ
qxKh408nmpRF6Hc4byzST1FLtxB69Frym+Ywx8lNXScW0zLX35K+fFhlNzFu
qu3OlX/s3VIXzY3RZJosQSg8Pcvz9/mkd5DsBEtOJi4CdELXanUYSmytBwOJ
ATPKQL/a90FaNpJPkSf2s+e1mzKTgJE2ZtQA16ab8a9DLYaG2TTqv5gZ/iPe
HIY33QuE9mceWsLRh27nLweGWbM9BH36W2Aeey6VoRMMgPUB4Bt59XFRildH
stgFtgDDlZ9oC4BT3/D3qVJngadPD3kCWYnKkPJ15ri5dZK2HvpprQDk1Q0z
/dIHpOlImyjMxFBQO5x5UyDjlenSskUI7iQCAAKPGovkQF5VOg4fDgU4hNHY
5NP+id97tmFFkG5MvWUzB8jCu8/jE2vz+saDBZa4+csinitiB0DYtRxCIXdB
EyTAXxUE9GHsrLNMnGvJoR4eikPoerpEJlc95kLVY7PPR4/6Xlr4CzDokatD
Q7p3YZPArOTGUspY3UVwylLU4GXXtAZxeZolEdFmU10MwMcR9zenmkGJYUPg
5ozrUx/65dYQWOIsYm2yfOE6H/ilfbJBnvN5Je+hwV7Gaj9TfendmUt8CNDj
+xbcsHrvb9S6tz4FcLgBooMR+WMshyrTVxFtbwNSa3zMRy5F11lW/oY+bEMl
H4f7VWTNj1TygzC83m6bUWwtXX3N1y5+9w+RmwBtNALWI3HTdmyWf3mXG6Mt
QoPgthgVxM4s01Ee/1Qx5FEksIB46Swi3k7TS8djWU+0vxLI0f/X/DYaghZQ
Cb0ZlsUlFpTXawbBdjND0hO6qdWvw9Yn6eO2tWq2i27vv3TkQot8etoZopjZ
u+TIg/ulnjYDKqrjN8Fxjrq4AdwSihzcnNTFq15hpwl8Pbo359yN+YG9ADbA
3T1AUGmFgnok5rl5rVpUgj1r4iXfOTJRLw+OxqkwlfTtMCXlb+C0SOYngXNj
ebZJ7sr6p4rwUsXWc6+LMtXs7DVAr2gj/ZKfQnRbOIeDtFSrmsPRAOUdPyJY
a34zIIKNXFrfSN5rfcbsX4onRXhvaZGZX4zIxs76PhI0d1Z+PoOKam359f+h
sm7CK5PSbIOQr2GaLYjJBg9uDuKM8lBiD1xS8D2iXtKgzjBw2LJLGzJwOHJM
OudIA70cbG8TDbcAgK384z5MwJfuOquExfw2FgQjOiCM/pn8dHuaTl0Cvqs2
gB2IAiEeX1MCFYIKldb1VKfggZ4HX0QHIfgl9Q+zgtUyIffnxAUcNsfElfvH
JLrIOP7XiZK2BTG9G23CezL6KEQkqt5xkOMnCTtXYjGoN71nHPpOPWPXj+hu
kZcTtlmnq8uZ0RaBSNfoL1Ztu8Zmim8qkgMkrNJ/R5GIXw9QZCsXMQPunF3W
8Bef1ktkXtBDW1ZK+56C2Mg1JZRhLrY45y94SIFDAytZTgNy5xcSJeOS2U+V
OgvmKhM5Yp+2at/OxogV1OHCGu2jBI150h+ZhJsvIcavu7kcgdmuYWAJeNiH
X+GwYu12KDiJI3nEoxYnXg0mADnQX75Dme6KaMjSfFLin+S0HsqPQXgzmnBG
WZTFqrvrJIJ6kHKwm7eNbmX8dA59EAC1s+PIGPA99z7t4FZNrZDzRhTgcCao
ln83Koxbx3lGt2IAOrzkCaA6twmMgjmnLct0+CZCQuElVKISbFvtX24wHYaU
ClzEUjU6M/aR34tSshY2nSkkBxJNXywQBnP3bbMMBgWmtsUgEW2RiA61rOCk
iSpAhEpc39kBpa1zGpyJmaF3hK4gRp06bCgrR2wJeigGbfSZPVaGj2eCMcPy
zp+YPYU7jViNVYj7czywb0aL/I/ST+rlRJSJbA1RXjVigMJISVv0rZEwlLBf
bUMWVN8pmNLXNH/1Yzfv3V2i+SsLsls2ReSK6llCqaos4tbuHC9LDWu1d1wS
6evqT7JVhDDyMPQR80d9cFtXdZ+ptnH/W7pydd6sEMR5HNGPmyrqgG83/MpS
1u7CkEUDahbr8PyQA7rwp0nmIMIHcD7jqjRa9mGWEJhmYGp1C7RvRgcvtmxz
0oFIpXIl9dfG+bQ7dpc8ezLQYuhwpbYAKYyipGzgeqG0Ahj7xZFlCqRt2Xkp
RkYLwBWxJ0Cj+sC6E4KbQCJ05Y1d0AtzS48foeUb+6BBwR/iN5anYpdWh3bK
4vu2ndWIaYXTdIJS2hdIaNphnDf/zpR2Vz8MRDNKABBMlbz2nesJD004jmj4
6Gsmsw7IMEcJayRgvEDyjgS9bDQSBWftORciUCtDqZ9FI+fyQiW8p/G1YR+G
UpfhviWQoligaErLbPm/686sqAv+594uUZiUChCRaUoCBXz77CTeeysRYBXr
+73aidZVYFLP6OveNdrDhwcKJAgFHX2rN5uzzXFhfD69gqply5dUH8/2Wsig
+L7lAs5joSgvj+FFObmABurdolbXVGqqrI5ElP0I9RGPqQWbaZFXJnAdyYKp
C31pI3SxxEGXxP4QW/zx5yGVRhR2Ok6vwQX56ZLLg0KZb4QVjZpLL1KUKs+u
HfpRc0ELkRGq7HRPRZmqVHoCvmUrytYSBKlx6Do47A9oo2btetTbw4hz0SQZ
uoZee1/lFuDp6NWkL3w9UL23E8SGdKmJGgu0yDE1+d0zzeSXTeD86XMPL++p
2CAL1G+vS8vew+2pdJn+ojxe6gYdNOa7dWeniy01jrDWnprL87tTakd6GcOQ
+MVep6fLbEeifS/1bXTgJ7H8X2siqn5tltBZA9sJHtUb0R9dJdglEyOKoopw
l2X9MMpbfx0kAZgf/Jm6F1y1TCPyxV0YVus/iKUxTXu8EnVA29UmH2qwAmzV
RQhYOic+6RGhG6nBg8Mlt/aETq7tMy9lgVcwcVmbpmAsrRdtD5ki/Z69caUe
2USNL/nYKlPRTk8ebVJDTAtf0CzHjzJHC6XOFRsRHWUiQr/oSQTZ7LlrRUbL
2JPPGNudsyWDi5yji4vFXdGYfsCkIIKSuvFaVxdJV+1kybIA+kOQAyuEpO0t
RzrvRA/0lA2E/zTxdMyoQiFJxnasxThnmz5Rp2ygd2ABFIxsNBTxd6Ac3h+N
AdRE61qWGlmVfCHKKtVImwkQe5sKnTy2bLDvFkhG5poougrffeiVcjsHHvZX
IDHOtvP5iN1GbRMWsvX4T3bXpgKw+9yDuiqXc7r+F2rmPm6S07Hi/uvoY5fu
5FYZtsvKHhDp2F7hTFuKy7CnaOSg2sx/OcjEDOnRRqmu65uBHqN2GDfXHw5t
ZLh2nu47mSXTWKLQDZGF9UKripuKr3fV07sXwJvymH1vQuDfPt+bUlC7W63Y
Ieg/t3uoSnP0bsiaG7l9OwPA7inlOLOo5btpKrDudEEwVOZtL8bU/qtuCNYO
XWa+Qs4GtrJVbGV2ReZm9hs+kVuJcUdrrZP/6vP8FN3pWHpfTyn1n+ajpzbW
KH5owUr/hAQ+MeVgq912y2itXNQgbYmnBb0FMHHYTd5jybmbOppebPZ8z/nU
BoKkPKBdngeD3GQwyn7LKhetRHdh09Ryxlm2f/tfOgf6Dt1CzPp9Ge9S6Hmf
Gb2+cmuod7cw5Fb//02Ix/MSoKshT5mvTgzkAkmMxcdnM0jrqtoZkSG5MJHg
wkWLQXVIWXBvFBGdAxvgBuSSLUoGe3vYxkGXkdEQZkswaLaBzc2RBDxswjvJ
uY7xGUV7kjJdCPULvFhPITn9nIVkJVfYam0SjRIOezRk3XSjOh1BvpiUm8iM
9R20MoEbtA8SJufePuRFtL/vOXVSJzgRh+NrH/uT8GDgdzDR7D4yAZb3khU4
UJ8R0COO573GlzfS9xmqPi4cforX6lH67eIT7Gie8m5IGF6yduW24eisKAcN
0N94F1WXfSH5q++lbclyol+nPz2TJ6FDN4FZUjsfVqV43gv9aOC6JhcTr73L
DFkQ43tR0xjXwE3Vfx2UXs96wrDRFQzK3JQAFMIlJiomjWlVg9ANAFlgbuh3
SWYJJTlUNnjO8rMRFEfQsepxCOBGM9N+bUohrz5N8Rr+i5PbTk3mfTmqKPmD
y3DuefL79iaDzKjSMfZKwL+J+bD2tLL7U6095MAOgqsI8pnBvsUjteSeK6L3
Hu4bsZCmR1Cncq2tfYl59dLgFaoOSK+gHP3GnfoajWJr0AFNtlyN0tiFcW90
8IWPhxxBstsnCsAws+mHf8eYgLPEuy6BDl2v+gW0ILirDuqLrR/ID4blZOUF
tEMUqlUZvFLUp5zGabXA3pNj35KFzGml8KQyXTOHvrCwaSiYzPPu/tN8WsJ6
qLkKX77G11IcdY12FB53hGx8hoYt6WYdiveE32nVHdjqeoqaTkwwlQctVacF
CE549KCMy4LW23x+d7O6J4+szAKzBngG301sUeNI4T0OpoYRax0aSBqv9kD2
K7QOLc275g9DbfkKbNReGek9dbVyn95NPL3iGjso1Z4lYhJdsTPddA5D+yD9
oVjbc21UYv4rz68pF+++nByTzo+tUQ/+T31hildtbKczyN9FuiCxHxkTQkrG
S8+7pA/32kqR3VfR9iM0kuXRhBFKzyPpv/bXAooSwfULDObcZu2nEPwquOC1
dI0PfmGQPOtOTKJ35yLa9kyE+QkbPODRDS7j8fl8uSx9+DebZzgY+TqjjMwm
N0VKVOQaOSroja8OIxJx5lGORcqUsXvC35YIRDzymZf2fqvfs4hGybzJ5mAH
qEJUNZ035mg1cdlG72uhUxD4rSdsPEPP6bBezL1Kes16XWDx7LjWxE6ZacfT
xdKl8O6AifuhVWEM7MUQb0YTurgwMjRvaCGmySbVKEwOo47f7nEJgJSrZF3S
7NDjPPLvRP/flgXqJ5AiGHkgi5oCPiCBOm4aNlOB26RrBePQhx8OzTMvnT3m
Hc7T60+iC+KqUJaZkEHsKQ04XyQ0zyV0UQ8Gr10HNEz5/ZFdr3ceeV8y5eHn
ms67J1qV0JpehjddpOQkDnXg/nXWOa7bjBqCI97NTSJNmbqYSS1ZJQflFjCE
319KuqZi3dj4MlYDFG2v1VRylBfMR8tNtHR13roGwZgoBEcJL3Ol7oDXVery
T/hjmg2vHtwzvCkONJOiwVtsC0zd4kHNdwoWFEGGkvwJ1fNMGs2kb43lPpO+
etSA/8/8h1GlwL4alD6xx5p1IImSZxNoRSvYUe+L89H1bMlpE0Led2cPMqd7
AJtCvljXPsPO0JsL2vI9wqarzOJ2Zn8xwsdHjoSrBxC7EuO0k8Wkr1cqVzYC
P1GMwY/QdchgVb6idR5If6N4xf9fTKg5IxaU6IY4pE4V3H7RIwq0QjhGAvRF
sv/oRC+WBJncurr/uh3yVQAwEsIxOr18tJDHQ/ojj4MDYChchA0RZnZPyoFy
rVWO7tBiUZ/vBRgG4iiwVP2Lji7cSpQjAVpvkCyNawHfs6/SN+dosJkR15/v
7OdGHikFSqqyZnkWLqwAScR5tOJT2jhZoU2QI+87cvk17RJB0g9jR/Poev9H
M5xkGBHw9w9mpnZ51BFiMGvHIWUs60EYhKmmK2OG2EaYGx54PONiK8PKBxsN
/3DiZ31GMbyMgSvZwE1fTluB6MautiQ62YjR+nOaIddD2beG0cvzEJ7Iz0y4
3MzkrGDFXVlk8h6kFHrEQicUXC8nGTbRNBR1swXAGpdHHL51979CrYjGB7Aj
ehYK75wSl60e13irGuEfO9z1qWM6kKz0bk+k0DYTBnLtHdIQz5jvw9ETeZZ1
E9DVDUjHJjzrO8jkt5hrfZ1WKothcR+QNy8Paqfj1rB8SY+x5kgvS4NWCslk
SkNy0mJGvNks4GIM0VxVC8shkcBR638GTdjvbclqIb8MWiYGw9Bv/feHCREI
3i9ILkRimHdeExKUJahxRllTZvSy54HjVDDX5z8UptYJASYvMK9q0AkpgvMt
0sgXyi/cMMti1XQaQ3QsJnHlnRJEHoZeQIWEMplbJ5qP4SascGR9p2tDpNgf
cfkUxIy/EQBU1Fg1IKLdJ34h/6k8/hEwL1hsa8S7Uzwk7ilGyOmTt+oPnJMU
2H4NhyhRM2pw657sF5kKF2PO/kUwgZ5cA+2D9TK6Rh7E3K6tVIPep/o0XSWo
RJRR8DWIT6MG9g9y7wWoNmnbXyKluNV6UbjttXI7X1v8czNvoT5kJ6yc3bZc
KeyG5ZrVod5lFBzfiX4d13FgxpJTSBlJZBVPgG14B+IJih5A6Y1U4HLCqFsD
5rSjGndWAcCaKLaIvxfGkhOiw6GACTDnqq5oC4ehDnIB88soe7oM1A75moBo
H3Hj0gQdR+7uU7YOD9s/+oydp9RCV6hfU/ezqOZ17nFXNByBGue4Yhd8YCmD
TWeSMcshAY2fMNTcGkz+OkSoEGVtSVFPBBGW+fFZpNX1N84i+taF4myyPUqj
1Ml/Xu1UbevVGuhQR6J2nzKrd/zu49+qKzujH0mbZn5YK8zlRBDwdi4rv0nw
JzR3WacTEL4jpwQlhw5Z1JJmfaNeoPD+RQkQxNAR7uzgu6nQTq+vBkGETu9k
PiRXdzOdEEWBNt8hs4XTfmVIZms76rkvzMo1P74X0Cz18oQ1J14xtzMUMQ3V
20NUY3xQuxP93Bqj1cCabr0GX1tWFfMNoE6TRZQBUBmzoSbPswv4cqacqkeQ
2P1NIR6zpkBiBPoUiZeJmz+OYvSro18Cys5GllXchxXRT10QgMYlInS6HLJe
hCrNalSj/1SIQSWQmhkHHmRKn4xJKG1HFQQI8eUz4p+4NUvhmIU7UUBLBLvi
sL4FaORC+ObVwCZf+9TmQVu//xR1Rz24lBCUuwzZAgYDIflTh1W44jwYIRde
4yEAKwW7uHU1DL4aDvt10ueep8KbjXvFD10KGQmmoUyf5sQ9ZdrC91sSuyZ6
ZxYE+oJkDjISgN1axweG+UHdoI6OWXXW0ARqeVdViqVweAf53ZwMIQoobRHq
oY/iOq0gYk3U+dVWgKKek96w3M4HzCWLVhOxkx4njAunSg7AhGPMGkjcSLmj
H9r+VmYi01OvLRwW07aSQaTKYnPasnDCwIL7YBlXCRoGTcDxkOyzuR56KUg7
IHWxVkutlRXB+UAHZOzFA57gZMHoriZdiwmF7oBI4QLkS6sWATqvcY6RelqM
cpmBb95DIM1tFlF4XqUNl+rDdxLIUu3GS/dhgyN8aEDyjG1ISZPI2zywysPe
Uhkfyt9rWXaCChfjQhYf+eIPp+WxM0wyhQ8YbNBt0SZgIBoD5PX/5r8IXR1K
dM6yI25JT0D1ape64N8eEkVJE/o/pHXkudhjgqWNMhah+Nkg6LS2meL6bSGx
6jOyCp/M2DPXxG5piIP2e56zZuUeg/Uw1KgLFPCjk95kbZjImegjzYHZDMOv
3ZtiFXHASI/oatqyyQMxKGTsvKwRuWE1griReISPAMzFRx+R46DGhpgWqM8P
HdFbct+rW5LvNHY2Fd8IhQjIhXtbWrGtIA74mVdk2KOQLXnsoevCV6ajoZOL
FrxzhxqBO13cvTn0CxJQF/BFhpGtM6TD+nP1qITDbW6Ryyovny7aGISfRsfb
42bNlcoqSiXQgOCkyRqnmiF4wOfsvgQawdHem4NRI9QEE/0GWsyyVoULB4u3
BFGwWwXkOVU1XiKoL5jxjQfCVwTJZ30pdN+V9tyTNb+n7hl8GdzhOmQmBYog
fvoymEwWLeXwp4CDFNq8vDp2T3CejAYoimS902PDGPytN5NWs5W3WpRWEJ6y
1ed87OE962ZkyWRoUgwld+aqrV9fwqm5WEicdOYbnMt8ZUcCQ+mLdeBphqCX
d1Y94ep1mM7XA6254ay+x9jzOGRY294F1djQbLFF551jF6JD4yH+mNUWuvb9
d4wR5n/YkPaMeAAPmE1EdrGgxpQYuvXtxK0dnsPAw5sSObOVLXv+JoCYG6x2
6Mh0Oi7Kafur+8jm84LXjo8fla6n5kz1M/4t1+lR3CTBcijOPqifX6Fzievm
QTaBwGiN0OIAoDKpODz5Hl3lONGqNIIlnOZQZLcGeGqhSI+5efbx+pBah4hV
QUJ1K+3vZ6w4O/Kgj5MoMZmhyvNTZWrxlf0dctqvziLJ146mNpZKY+1cRIfC
akT6gW3soolHL+GkMDFdz6BCw0/dTbMs8Yqiu1Qn7ddv1qkFjdaJDKj77onq
xBm+Bwjn6ZHwznCmmbaE4iqio1Py/lI9dqQk6BQDhyJxx6qno5DaGPpryfRP
SbkPbMu8yP/XDBb26GIfFH7SvFbI5GeJ7WrZ8nRNclb9sT0pcbM6qNY3M5C2
8wbdOGt2g5DEZCNef9xblJbtZH+5HsTrPj7a/7F8/74kmXO8jXCL3mp2TucK
G6wPlJlULb7Cb36Jcxjp5QAzLtJ3nfV+HTXGTJylzcP6C1YR5X6e2yLD17Vj
0PiiCOIrbp7eDSmoXw0Tcl84sJ8owq7H/cnxEZGWUQERhPvvsqj1tO6HoLFI
0J9GoLceze+uAGZIqFSWHZ51zBh4yMh1/bAFJ41fELXSsNAybPwtzwBmuypo
/Ul/ofipQv00q2bfPfoAwxd/E34rN8t5zcRt0NLW+/C9Jjov9ZuMVIIgzKgN
BEDyaVDPv+X4+Mem6eU9vqmaRA293gzuJ1kY7bcxeE4pDnrTVSkoRbkvglWn
gbN3TCjrZWjKaumQD3TccRa/B0fxoO7wCPL64hxw8McIkPydpJOXBu4m2tRA
4dDcbTnJ5qZB6FRWIGrld+JRqKjUXlhC1aqwqwCt+a6nbQvxGI5AtZaHz/Ut
S2FmSxvE9u0dxH6pDX/njFvtZ3SwZOIeqe4xUUcagIOidjbHhv9tGCha7He9
VYF/RSmE6vXWxxxhD1Q1buKG5f4uqsaurpMNhIR1nkPTef/ws6dujCcR+YQ4
axlV+FfOelN4lQQ6pgiwklzjDUgZ2+39eOrT+FeiZN8fEGHrEUxMM+gHNLL3
/nmfrqHqN8UA17hFOUISPyBxQM5zQ5lz+jsImgQBwdITW5PElIsns5nen5g7
vj3LbuCUgFykS979JPxsppJIByn+4tzuc7f5qk1LDCUGtgiaDH1oy5tMI0OL
W8OW93kqI81rM90LhSLz9xypqZYW2teH8Ub8rlQWKvkaJPe/mCRRVhncUgDG
RQBK8J9hf+AKblVJSfztD5cLTgjJJo8vdjfdZC3D3fg6nmSG3TC2eMAhzO+m
ckbxmYQtwhJlLtuapbqm+Q6zMoPxfffNT8nbzj4ozcwZFle4h5mzXhMyO2NI
hkEP0+vllTF/weUngHCllRLAD148r5enDgO7SRr22FL1E5aDrPwbggP1/doi
6iIrv/6tedSsZGbR2ywl69fE7l2qCpDLpN7a1RC+sRmSOgu/qVawtrpkVrOP
M6HSWVqcoSkp3AzD94NFuqaKcGbmmGsqSLYaNe+F0/gE9uH7546MLy5XKjRB
/FHHVdqrCmNDAiB5PGcrHQh8vWtA84d98MLV635UT15oE1K3q+7FedInUILe
tSGPqta4SujLJaWQNSp0FVr8yAjVZ82nx9FVEAcrFVRMStA4t9M2RygGMVZt
t8St8VwQeYHKU7sN/9cTwepg51Rk2N1Oy1DH5b94j2Uz5Mmhp1g8uZsPV10U
caPsoWw+ll7cHXVhOx8y1r7Qzo34MPqhvw8y/vwFQzTdC/ab8JFIYcOQpqwQ
WCta1tLbBwMVlXEAs6E9iEINgooUg9By/iPVAbt/NUES8m9Rj2ihvkgtlYCM
0w9PsYCsNzLzw4/ClknEfUVUDW/8cg8EEO5VH9Ki2pIppjPHUQbNkZXeCsfR
TC75iHufzcT+cbFvZAUv7fyQlrSfvFS1qwMlqQDfyEIDXq8Yg/rA3vTwmAIU
dgrzID89xz1h/QnK2SzJ2c7RsY2i3vdmO+2SVHfGD/gn/2MD8EuALNBkfH4H
8n1cGJjn6W1EzaWQGv7YUtSDqRVv70U6XSp5W4JbhpaTEbTBEa9uAeYnzqDj
Jc9GC/HjWEPlE1BVwp47F5Kw9wsEMzWqd1yei9hn2UZ4zJMgPRTif3jcDG7k
HQztNneWbl6mMfx5fyrRTyBoXpwj2w5FiLFJODWD9kNm3w5BY4EouQtOH08p
wsjT02kUrcZFdTeZ18Sd77tuo9Vi/7Gld1Oww1mm1H7tUZcTfV6h+FoqMgPU
iYLK2R6JJj3YAK3eYPgeXEl8GrC1WCImpQY23Tz5efudxLmdaUgECeHrI1db
WvXDBGm1uFzOdU76sHNHRYtYEve+FBzyjUU74zRcvBuFXWlkC8HnZHmlGfcf
ax4ntyHe09VN+zpbQcnLJOWJjWY3FSa8CG8iE5bdq3TCQ73ZG5xfO0syyoAv
ltAaOf2j96ENd9rAhqegjJWlxecHMu2th8dbmoqWxdoBicH3hO52sVoSlrjJ
Myeub/tVfNSJKO93pMIfzUeczuKkd80m7vZc37kqmLRoqhggNx01F54/AX1q
j2cItGL9oaLGJXAgk1pHydpZf+KeMfPuTnWoufK5STFDlix+9oBoueHUf+go
VwOeQRyAS6UlkHoet/YwknmsYCMeSy5DoUcOIyLNiW5B96fNiKd7nfisNDUo
tKT+v4q5uuqjIOXS0r1tMwxHfsOQaIcDw2R/H9+rTtBjv3tC0dk0FlcZu/VI
IAiOJRa3BpZH4+6YihJHmuY1M/GDs5evc5tmxWLs9pmIdmzIP2kg2KFAGQsT
w7JEORv1NnFgnwyCJO84Cr5UbR1QI4isPOfBL0iNBOqPYYaeoiVhwI10QJrH
VW//lBnCtPhTW+ysci2NyEBos6YDkQ21Xy/oYeenDZue71s0dtEBPkl2o8n7
XrXWRaYIcoHDEvLDD5L7tf3/8Iv9Ck5bxxtO5QlvRFj3Hx+tPOoJPUxrXsHl
+dy6FbnKTiRIxuero1ce/BcGuO0/PdnlBx7WCDbPb6+wPZ2OIIxbTVDgU7Fa
yTIwegSed+WQi9jGIxP8nsyvpmALqKuJku+7Vy7iQWmX0dlu5IcG5q/yiCFb
7ryItMhZRg0DHZgNYk6XnN+ellQBRpb07GfQDkBnFbIHPBFT+xgpT3caXlFZ
j3Ul5O22k49TnNmAv7LPpVOpkmThH0wFOrAppX3n0Xia/vCOamTbI7tCeOGq
wp0WAevG08WFoSXp3Wh/en6nMdsRw8kOhQBLa50oRrsOM5lzng8+bcE3HDIp
DjHYfpIbLO/n+XKGt0kdZQvk3tpjzcWYUQKqRlGFqCCzCV0HpUzl+qlL0qF6
d/OMnrXX3Llc4RWbBhfuApfNDSKlWF8ybwytE+ui9u+9h4sxzQ6bRZ+Ea2LH
KUvVOnChlasVzIFWEO/BGGTKVBfPrl3nxGnK520BNbxQN568svMABD/8TXqP
cxjrRPu/Pb1SYtBj+FZURnmbOLNYGD8dJAY6LjyHptURfyKB/30wklJSU9PZ
UroK9t9+FCDawa6f6vzdoXk6g5SS2Yv9ccGFqk1kArIha4IzvQ+iwxJ5nGZA
QGJQU3HMGs0l4LiX0iTP0aaTUR09SyXCFMfcRh6Y/Cx6R88r+2UN2nsd98KZ
aHVte5cnExEQyG0Dz2rEDXY23Wh4TaLTaX/nuZrjYKEEzYzsCPdvLpbdHNA/
T6wv9EUfRWF7N/JCuoYOTw4eP4XSq2CEypxBRDO3QGM8QbDNi0vgyxXwFkx4
ak5on5F+DjBCOwSWGRUMkKsAy99jeKyFuTs4FTcmonabF+O+vfXK8mPsKhvw
NTbE8sFLZweO36NLWN5NDYzFZ2hk3ugpuNK1UxDV7d92X6ZlWpv33bRI3Emb
nF25MIry9ErL1yY8VLGl73mVAx+DyVfcVrQ4imVTw5VPMpIyL173Jgght0pm
dIWTV4NAKXbSS9Q42nP94pv8l/xoQs5vfjFfSsVpWO8TY+TWimHkhPev1cms
EKz6BdCA9BCv2c39lwlC9hsgEtHHV4KZvVArq9g9PMWqfmun7xLqghy2Y3jP
6/ewlpDlPj2DSfcLxVLINd0iNlpLO/7uw7ymcuWoN8Lfs06bvFCnDHHiv63e
C21JTdBUWuilGVg7KpP1iVbkddWzMQadhA+Eb7jtdAngoso2xLXCHu/QsC6d
vi7HHVm/1ibDsAOLqxchQu/Cv5LWhOP40F2RRxmG8cj0WXILysicQz41CN6L
HC+KpFhFNj32iyCVz/XghOEqNduEQ/pMKHVEdOORCBOCcK2ttcHXjn0TyN7+
3Yoe4hIeP9ayDHlqb0PwS7ml+2TbT8l35jXscR4VjN8gwwFfmm03NsY5H4Pw
ancfkSEpZV53k3nUsZLBxNW96rdYas6ikDeHfxg66wCMVaKeDRASzqpkoJdb
ofg5Ic5irrpy7BWem4LCOjD/ONntSo2sVBAcIYw56izyXwOd2fLFCTjBJIXY
eetxOPCvrYcF6PhsB69ykTVvetRIHwxUIwa7B6CU+JlLhn4r45ZD3utFJHFU
0T4tmN1kioZzoJsh6FdoeiENt84j8qKgJKzA4CiMR8K5DBLdW6az9XzGVaVn
iH3IopGYR6fJcjkMcFWq9H/lxNQDq+DdP3SAoMzjJwq7Q7fBK6DSnBiTssvG
Tb0eB5Sk5XulMT8Ua5RvgiITdIjIEpZACufZiMP/YLJlIkzaMD2tXAq5uO/4
mCA0umBqcxTpGC611pWoSZX1lN1s+wsvRJchMmhC6/6YUdxQE9ndjTazx1Ea
VYT+wzOpP9r2Yu+UDmvOfFmqfDecmPsuKJJbcHUnhFGWYjR4AQ/OZmq8w+u3
oDvltexddbID8KXsHfr15VSNlNqg/BBMtKmU7/FE/fsKSNKoURdR257Jc53B
r4WuEFE1y6Lv8iPOtv7bUvhikHDJ4AIjlBQgBCUBwD0qIEUYPTEz+E9/cobU
9TlulqFrlZyiGqjSoNYikA/P65QSU05hLTsIrPer2zM5zUrZeTfWvHQ+yyFw
uCJ5HEcUo2P45xQGRTxv6H3Xr8wL6vkfrnrz+iiirHNiLw5Ju+FXMBIMDVGV
1leIQf4B0jveneSG/jtnJ9ky6uoU4IxSRxiGG/I8uYwO1coR0i9Mn4sRRWZr
DaA0F2To1KKP3a2A90mQGwzHXSxNM6xCL09QMzT8dXOKnOKDbNBxetZtHRVl
+5b7hC8k4jF6pLTnQ7Jt4wFxMjTPz2DsaSRhlSuNGe6Cjaft8PzXW1pjq0LT
2XIVYNCIt8sErHTCrKhxo20R19YbosiqZ0m4zLYjn8WCWAtjWEmBdMbuDuyH
ohWSWqtDvetx2W/RaQ/+y4ftnoS9o6TrOK8PRL11/NnLPiB0Aluih4+QB2x9
5JQxAFaiA8uqupQOkNqTpXn0H+moFTVByyaDxXFf39DITK7nCtqhmbZJ3amq
xFjBBs/iF0CUdP//7KdMAOVVU0JkSuZxrtaqao9n8U4+rYodoYl0LAAbY89H
2ZuwSzefX0LXY2RNmNk5D1y3gBHqua9MO98o6XlvooK7iClvGvzjInmoC3vd
vbJm4SWgCiKxWwnXuRR4dG01HbZtAFXvsoDDneJMEdGDJCAY1r3cxH66g4L5
cdol+V4Sx0f7F62xbya5hWATiSVCRtjsAkKzIDydojILVQ1SZOlPqWrL5H87
L+vMcLrbygfQwxbm2h/TQGCyz9cxr6ZGZ0sbDXfDqM3xduJO/3cPl2b0ENIf
985KPi/AD3N8UeRd+2bkT12Matm1pYrMwvCz1HcBd6TyG5IbT5YauzrikBPw
WpTYirkrUuUVc7yJP5SWWKDbvrMRM31LsPQ9aNJ1bNjJp93kCM84Q6HQ7pS9
SD/ZdYr52RhRzhEDUB4QBhkzNEFGkpLN0I+CiwQ5mG211kQwCk6w1QcKJkM3
3u+kZGV5bdbSL5QCrHpAE0Lj/QYz7EWkvMvHccrc5Li4lHRHaGJWW7I/8pWG
JMBnI8SXRUCHWSGCD2/SDFsO0PKY3NDHOblCmg8YitBJsYh0LxNqlkqXlJO/
TsQaBRlPvnKdxqkbOk0umEWW7Yf9WqDKi5vh7bFuxmEcVcs5qoaG+QpSoq+T
efgrMOld/mQtLDv+5ulcLaD52rO1ash3ivGTS37xv/T96bgXxE+siDDYS6qA
XcY4lHc49FfY67v/7jC18UYnC8ZORkorsJh/o651HgTrSwrQqEFmclzRjW+H
Xgm3u4DR0HvI+IB2u7bjuKGA/f1ZOZDtzhpdwhxPOfNW3iHzI8bEGy3w58o8
i8fNylymkq9nZv3j4l1pOZKUl3ubPiVfnH1UeTH4u0NtLC7+N3soeDNex9tC
m2Etxp60clC51TromBbs/ZuoqIlHRF8E8AIgfshxM8FwaDAadSyHERLf47C0
zsHN97DQjlCmWbTErB9cGVQ92d1iFQ+zCpPlkU1i3NSuhtjWOldwyG5y3ewN
YbgcGDOCwgg/as/pdU33p6W/pQIgfBCO4YUnhWxK/DrewCZr3szR04wjeUMJ
CCRM/QM+HLtquZftIA/OS+k9pMdw9Q726q99zyGBfAzesUAF4/huPQYaVatk
vXkxrw0cHH6yn83k8UE19FLMr6vpmrUGxJxUf5ZGRqP4A0Ni2E8446rrbTG9
gjvOpuKVjJPmP9afUpvZMr7n1DnB08EscahMqHQ1bDYegC3P+fEZIBRf3q9z
T3kUsjhgYkLQg1NS3c7us2XHeSvFg3sBjIuVTHySjl/DXX99H1zY9Oz8NV8H
0zOE1kyBCZnPLKTtz0hZ1/4Zozuqw79vYsT4C9RW4x3XfTaiXSeawNM934S+
0Xsn+B+vzv217KzXyfZ9I8Wyj/lMakSRl6zC0OByrJZ25AmvDGRqX/hhqHhz
CTI9gzEEBWxICNpb0PLhZSOJvvRoREQw7XJ8TgKXs2ymzmIOMJTmkZeohvnF
mWX7kf9BXLHSohC75kuga85jRSTPY2Y30+Xaz1wOBL+0xmtBDnTGZ7SPBjmq
funFsIz2QDUgq9R9YLwj3/Np0LHiGiWKBdj/x37C2+Zkw6tClkiQ+Qxh7Bgz
cXy5Jf7MCgPB/0TrgP1pCYRnmAYRh7Yc9SWbH5h1vM1Ulndkp0CZgzJY+XSd
U1zn4heJ7FewLZVEEdFwDXAPSXEcSOYd3+l5J06Ap+D0MkELfhFzL1R3/gjD
nRs5VIavIN/UK/LiQU9aEWRcN8tC/a1XeX0HoOqFGOwwAVVayDXUJrokXBR0
yOG+OZEvlCKfQaba0AX6Hc/qk44wClG2E+p2CV9T0Kmmg+M7AZRC4CZ3ujF7
HoifZZ+i7DI2HXeUQf5f0zKMouneBBV2L9a18x1tfMmu5LQhEPu2s/TV7vO9
pP4qrBnz+Bu5cLsevh50QTpwjj90rktOYMyc6FyXoYSS774GvIYeIiqzzEP5
p84WxKh6vnDMiiH4qZBwmCVeArFucXjcOQbYIa0IkqnSSplkmTshpCylb0bE
ubvp46PjgBZoI0F8MZ4SVPQUA97tiPp7fqmIRitB/wV30LzKrSviIB3WYlwT
iMD9kOY+A48qNeGAiTrvIh4lmBvziFgl3y63Gv/UNbb3SdFI14dYu/iSN6Yr
rXpQjZonvvwjrCbtTC2uOJ+WIYaK8bCLi1WReFCF2JsPzOtWMvo/uzuByB9W
F+kECXlSRJ5LxFM+MszvtEsQhMG32LFB8+Xu9v3WJsJFbDkOx6Bc2IIXnXLo
S+Uw1lPeH9LCTUXeCjgiDEU7S6/yGJ47gKVt81UgTgcI+c51IISm2HlmRosR
PrPNS6e+1899nSMBpvwveouptrlI4RqmcVqAMeTp23gI+7sokvPkwjrPrVst
WcRKFkKHxD5uWO5BSEsRFJY4eLS5Mo0O52AetIO/ezUgdY14BPhDCzrgJ6Iz
tK3DNMdATjVfAM9Pj+rlFrgiBUcL7UDNT3ADhZi+KxbKVJ/IkIUlJLbTcvTW
iRzi3AQ31c3f261g7JjhYaJq98e542u2fDKWM3uPaC3pFnLzcnxUypQSaPO3
rKKa9zpBM1UFN17YMDPyvgAcM3ijyAcNYHkp9XCDqEq9hqUteYSJnfkLZzk8
TPlgQlESM8Mv23mLe+nfogYUoDvOLwrRJ2XQBZWGm2M39/r+1NcmPY7S9w/o
VxXEjaiLSyzaRwSl+aim21bYVOCjR2n8PGd6dOKJOx5TBJI0WpOwFdDXQo0k
8L1pXK5s2Kx+llB3Kbfy0NHMqkTZfUohKXK4Ij3Hc0ZSzN0KXHyI8aTI2fcP
a+Raz/YtHkp3zQBVY1CzYUOWZx8y1ZE9ngW1Pa2PdohxcIahECS78vn5ySR6
AJSEJCKY6CPwYaDzsm5noQhPertoaWqRWKChg9Pwxcu0

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpehRPNiBn02/+oHdYFxb5wJYWjl9h92X4ffNo21XWZz0tGd7mkNA10oYkNiCldYIkbZFoszuOyg0ecrgts82o2YVv1zIUyTUyGZyr2z5Wv36lPfAOYnbBb9GmmiQEOkNrRK0KMyVRD1YedTOS9O71cv7aNBdUw2HY9ylUGxSPZLA1kZL613wFsvYndD4xGaJSeRCswL7grcYWHj4NZZjWpAXc7h0/cxdRJU0yJEwym/egI+kk3Z6Hqcfbrj7Odctquqy6FRIMUUeazxJb/B1CWuyDZf4jdDSwv5jDRXoznQ+f4bymQ5mMmtXh9UTm94rxPctiLqiC6rlh8i2N6T+/HcXfxpd5p9pRJVMa9ykduzE4heh9qGXae51WWsS2DGxEgS93l4W/wYEASpGSopIM4nvgfBNVkZFi/EdJ2jYsKR22iIboPzKW6t+M73RbSQRNlmyNr/5DCsL9fOM20D3tswv8fI2AYQd9CN4YST62kjPYYE6bmo7VzKaFmYYBfvU4oe/HBf3EBSM2MyJEuLtsFsMT3izLxSaBjefjkwmtFIoccXMOmBs41GTxqkO6ND/50WybmlXrtWwN2/kgo3Jpzer+1Tf9S+9WV0tapZhh5k7M7Pn2zhMqqRhhzcb0PwRLM1w7Xvv7iO9hyDysbs9QI/nJ89w0ibN4OTK41BsPt+dOjgzVqvipoU5HfRAWfnXpoThEfXpOqnOJlU2XQK/1XyEwkXUSZtM6r5RCxVQoOl81/ZuUoIPXp/fbi4a4DXXX6jzmrZ0KTjZmiKhuoUJlyW6"
`endif