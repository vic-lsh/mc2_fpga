// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MNvsCY957FCgr/sT2G6D5BKOcNUrWd/9EQSnR3TQNu9QtHA6VJc+Wv+4McwX
DMox624FdGXr4Nv9HujeALC4kqIBvEn059Tl+BLzIGC0f3p53355NKeiEyw8
ne1KtS8Tedvm6/83nkqHWpHTJ1Bi4YpS67t5mXU8BPmoHP4CqfRf+xDq7WaD
bPkFOhzyDoFYCLlxscIg7KLzUUebDa8KMdMxBL3R74eDoiW8LAFZpOuzleJj
yF3/8RCPo66K1JDwzMm/ZWG81lZx84YdCk8xRhLwHccL5ewEMYHQZkvEgMsc
Dzhml4CQKh21yo8fqy1JhNEUghJxUf1e51uteMU6xg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BSTBmhJIzJ8B+ueLhIFECDPfz70uDdz189VU5Sc6hKIW7xLI95B3yF1kGrS/
ED69Gf9X/FqXKTrMoJkLnS5hQafJH0ROdQnZPBJVeapb1jMVkICHG0WDVRc2
b+EOGGpGo49kVrqvWRxwkBFZVsbV11KjL9AS+uni1TTaHqh04O7Bpy1Pd2nJ
UlQJ1D1KeLpcZaJsIDYr3Kw/d/gsTIj174qAVA73XLsHJhO9YZpVDIkWqJVX
L5tLMhJ6lmOmN19YVCTtw6oOtmmwtHSOND+98C8wfBvd1z46E1bg1DqTuyFH
ie9OTzKuypAFmHrxFAMRKPs/u6glXhd+XTrL/7kBIg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XItwM3a3N4OaXOfEdAj+GXCEoKiKsfkekxBH8HvgYTTOhfCpzRA9UjWre6H+
EugWNXepamw7NxdRpyI/fTy1xnH+4FRyr4VB6QCDlrZ/Bnh1LmPHuqozwXY5
Dj5pPo05iPRUuSDPcPBxfL2BnKcaUVVH8vAOfsBzLnTnWL3XrhfHJkIn0wL0
0gsfYiLQ+v2q7UX0oT7LbZ8V4b/HTKyAK6y5ejuxdZI42K3Ghl/L55PGhR94
vSaFrKRNopOWBBVAj8aD9yFKLZcStEcGPS/tGjE9E/emOHKa//8vIW+XqrqH
97mDChK3BoMqvfsxYAv+HJq1DN85wSPvRJc0YfQrzg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g+FxdxAnID1X7KvwE/phj90jQZlGrW6v7tql3LQBPE8HQ9MaqdZ6y7u/6Y7g
IqI2s15BvvoX3O1F88ZbsuGMUY5oaivDtMyRyD/8eGRQDy9OF1kC/ahSCA5W
sAQ+EKA7PhnZZQYZ6L/xCfErond4ILlk9XiPxW6X64JxAsu/Ng4qWgZym7bm
m2fE+byOcxBXYG9WCYA3BHpPv319RQfzI7/Nt57dLdWMFeqXz4/eU85LPXCm
ZfseHRnRH2LE2ptZ+4friHrrMuWpJk/iaEIz9TD1bEh9xRFFmxm8ZK3B6zoP
6sheOd9QBGpzQ5Nw198MIJt3NlfutCo7+tv24luNwA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MeJNeW0TkQMi39l+FIg6/+YgagjclUgPJR5JYkWe8l3M5X55uqOLLhc94b+f
cfGTsHUBHVCcIFT3Bxs+U6tWwRzq4hrBzkgGnTzprnwXGC/gAndIwsRAc137
GZEeYQxB1IApW34TmE+xBOEpi63aplhnWhU2J4pU6uDn9IbpGLo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oHcqAhdqMwWtzg7igYz6CHPuSTTA+VqBkNH+IFgjnP3NLKMUXyczF/54PUkE
wf4DePHF2bRO0CQtvkVXO6oE74uCd2pZc568ewR6Q4BLfhHYChaHv8Z9qCNe
Tqo1ErsryaSY/DGEiL9dx/5MqLGIr/ixks1W519/lT0y88Yg03sjDPWlC8AE
VF0zE1ROoVH/LqYnFmw4lJ4YqcdQcXOa9IZzvITKuQlL8W9mqZGie28HGNM5
DsmygVCjBNf2P+kdn9LdeZwJmAlC3ZpQmZnlr0S6OSFWRFKx0Jrif/6vu7Jb
jfsFJzIwCsWQasV7U+ROAV7Q0aJjJO1vQZML9EeBG7+CgVYqzjA+CpFpqA1X
j0lyJKbL8VLLJ3ngkfQcaW8XYRpqNmuVjbHXUNv4UUh/mVLjHHc4baMMvhZZ
wzxLqkD5TqhclsXzDrVfyGmhBJ+WZ4SC17CSe65zjR1YSPHfABnvvfsqmukq
VN9e7P3hhkVRI1/CeA6zWl56868GU9mn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hmjjfpl0Ths/tjIw0yRJkCwaCHJnCaHS+PETIOno4DyDYT1Dy0v+ZqKyLiqf
uaJp89plqV/eqk/UidWhG4pEe0/F9Law6rr/2ngAhJk8BPXh6sdzS85b09Jh
s/F8QZKc71cYiMOLsvIvka8ZDK7/HVnNc+z7z6stEw1mxclr3+8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
INI4OxDh7IjEjnCmub/u+i4+GBrUniqm9WWgc1EKE/n99HMtGmZ3hCuYL2OU
Tbk7Y2/DKGzlsx0vHrgVDv+/FH5V5Mh4uuW1oAw5zUChG5ub7M4h7l0Z3kfh
c9BD5mSpX9TRSV168y+2QdfOTC55n8n4AEBktEo4kCHjXMVvnUQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10016)
`pragma protect data_block
qtuU5Py9SBXUCiX+bzITYhugVWcdRpIZzwW4HDC9o6wPOEJJo2m4SNBOX7mb
AdFbP7fAZSEF8Q94UqFLP6/2mkdAQSxUie0q5Ktg69F9k7ftQ3OLYp9TpHUl
41bK7XXikBqGMD9RWQH9RiNXTz1N00D92mKrsyORRUDU1KklZ63uGM6dgVaD
iXdzsS7gLyyMOVJyLBlK1dtZID8TiL+4roPuw+OqGKDPsttyc4cRYxI3qony
Qg46ODombWtb04lUA3z6FCATnun89I5jkZVujsSyxIcna3Vpdh2R5PxBkS2x
p8ofO60kuPUyLiEeawL+yn7URtpHykLDU5tnhXJAEdh3ZsHa2KI8LDDtKTFQ
aQJZR14k10hv20JnetEh7uRryrCt+Z9JPnT2scKgNeweksJgIqXDPIIjY2yk
g91qgbRWIgtLfanX2ERgFbT/o3YgVdBhj7AZ9jfz1kSN8hW04lT55LZh36CX
Sv7V1ERCgSIC8DyeD5Ygp5h93lv1QHdVxTvv+/7BqCWVW1duXj4Qc9dJssSh
HETqunGy7Zn5zfhCyPRK9267G/y+jayU5rqhInwc3nVpemxBxLHz2NdQT/Sy
PIUTobe/V69fxnQ/W+YYZ1bAqeVMBpDJDTYxTjifVxMij86gmIX+xAPmxtkQ
UCde8j4HfT00C6dR7Xm8Ie1rCBP7bSsYw5GVTfZVMPZeRny/i1DQeEsTYg1q
IPEMoq/HAWl0AY3SXQf2vtDYyOsG1sRksSbhzrVQ2fcB7Lu4zk8okGHbJhe9
QGEVheBJA/+HBr8rLd1ycSbOWoITR+udD0BOwM/rKa8HRmNfqh3KcsfSXK5Y
B7wrldAwaD+VCvWhKHei0blQ4WHVr1LOiwCQo3KJnoJTViqxyK7SGif9pwA1
0Y3ghxZcovalvoRVW+YCUskHBCZ3moxYMB5GSxbHYBk9HIuKV23BINk29D17
Y4esfzLMpNDiE76A1ztMIM4nvfz8t5ycBYrKnpGnnBCTD9VIhfY16LbD+DLA
RioCQlIJonYncDkvxNuuj1eE7AiJrJYlRqojChx8mezPTrm5ogCf8TG+Uh0t
hko6HyN4i+vGOxImwIDwMPJbbkzuBFZqfbV43Edbf550UfoANlg3tuOC/Qru
bfYgmk+cXOT/k4rDx8Dh0GkLnZd5vUcWrl5pr7c5U7urJb4hxxpmWegf4ocn
qXiRjQF7lEa5Zhu1413hQFy0f/v0dmLB53V+xCpXEGyKE7FL4Um9lSrh9nju
7Eur8Te+3W3JaMzPbkwVktRUZwJdQcUAg9Si+CGMVtrTqhsdMwrYVxDwVV+J
RWbGnxSIDoFJdWVCwnPtEeEo3uOiKF9Z7NitoklCi71AV3J0TXOYjFrIdnNY
lV6B7C8tr04DpaNT5o5HgS88eYjLp5EWfGNiPRZN2FJzijWm5uRk8sLwUTUM
rpu8eAb6xvE0i/FpiLPYc3RpITDNfqkM4yVjxf4hfbNEe7pCzwD/5vnr7vo2
KpSzC/xBqnEWPuqFGsNCryCzuHqyyrNLbwCuRnwhd1X9RGHE7lCeQkjRHObn
d9sZK21XbHXV0LboBg1LTYpHjktffBy+rqXXtsjYP2J+zXqmnu8pT3RSVPkq
vbB4kHMWEqjwcy3HM22fmvNmOVGRkT5/o1rTOIKE+5jxhTw8zFg7eXGKyv02
Kpcao6oNPcBpSveCEEAJr8FCqMl8Q7+s9nHRZXSVOtDfiWZBD0VK5ugJn0o1
OVgx1vFT6vGuZRG6tRk/YvATnKwbrEbPkCtsbF5K9/975FfDXkSytS/t3Gvl
FhQO1z4h8yydGz6ShT6o1P8uzUAtBuiMgFExWiRivSdSupPsy5hKUhLK7cfj
s1J9C8MGcxm9sfhnOO6I7fCof71Lx49g4Glow0mQXfZRSQJdak3E0cDnTCNr
oFLcfbf0BfHhUenJmBcpzGZCIHS0+TncQIObqucoEc7m+efLy2gcIxlpwgFY
DDFvwVtFwKR/FmUDOSGEErK5ToaRtCb8ln4Xj6jc5LdWZLWCUtlOupXDP6yU
Urvwp1F0OC/2vLhfxylWgz+KioXehxMSKZH0/dSDnjnwg+s3hKfjNZ1qxfWz
NGs7NpOXL27ZKQem3J6Hvkp17hX7F7JFj5qbDjZBqMhRc6o+28eFKbNH26WX
xUNqJUjy930Tyb0t9hpVrIlCIYMna57FbzYZXHNir6kYFCPW/ZNFLCuUh5nW
eGHDISFp+cn09HKr3fe4VNP7NoLa7F9SW5iNyg7XuMx4zCYeTbatIH7dZl8E
o05awURmXJ4SdhCicLRozNv7pQyu423D5zZ7HGobZ194gfxZD7IdCyCV/+Ru
CK8TMSWf4TaMc0l1jiYGSVvh1Cb7kAzsHnsO/jJncRgyyI+WeL0pyRdv4c0X
o8rTvUX1Ca7i1OnVT0AShz3JObAvTegT+L56eu9a/doxCc+/LF7JQDZXUZEs
76i3R9z37NeuRCTpsM02U5MM4soVXBidKnXfN4KBcDtinE8mKyDjjBd7GZxQ
AZfDHAdlEcFE6tdQhAK81colex3ox8sEnH+rFHvIPQUKk2p1nDh5wCvb4SV8
c0aX4UxT2cPOW/SxbnTTgow/KgtlAt3e5hdJRxdL5yF6H5RUKvmw3o6qnIoh
xqvj/H1+vexAwviiBeu8AlUbxt7s55M1qlyGZnW+7YsW8sZMv9AfWqUypr3T
IhStrQzPy6HEpc+xbjpqMbHTeVhgCKFzcwvOsB5/u6CUSXg2HV8mvQXS6Tj1
gqWeTivdelzkGKWs7fgNSxKfdi+kpoj0kbdt4MEsOeXHRkp3quPvtbgqtLR1
FtAllZ1JarzITqxRsUirzeZiAVnx6X+pbtdEO17Kb3QuOmJsUfXuzmhixBGX
GVckO1/UuE4mfqLuHW+VstB5vm8ycqzQ9mX1EA/tiJqFdKJ0N7qVTmzmR+aX
2T4+otuBGJ6McJQ4VMbJUmJ8bEr0W+24Xp8eiaVdutD+1gHfnehTX9lUJ9Xz
XHHZiuJxPOx9ZBNsG/s6Q09AuwN65XFLtHnQHtuG1RltJoTIQhY7Ba7NchD7
5rVKLcpDRvrjVhMbhyPbMEFk+LNfx8ejQfeIRlyJe9Y/8eUvzkOSFkCZwXgW
hUzwNLf+wsDFsY5irPclQqajs8xg+oYrFWW5TSWd+So56ZICMhehrMp07S5i
kev/IGUR94NYWlJR3nEm6AougkhZo9znOJ+v9Q6DGCddGlWabVYfv/9AsS+5
7gk28Jo+KFsE8JGTFuHVo6n0lx83hr5/CcPSOoOJIkQSeEiefjisw1A3jCwb
SV122e2nfxyO1OP1p2hBb56JFadLsdAbPgRMiVs/zUM0PGHNJbH8Yr3Xv5O2
twZKC//VO0aCkWdRsqDKZKcFnYtApx6n0mXDuhkDj+lWaWMeLY75Q2UEVY+k
cGPMK/G3d5cXbugxiC4Q4Sn8LalsGmKLrmUDAq8PYTl2oU/hxmCL0g6ixFaX
TuNc/dmLY+Y3KvlXn0LQCSGtwW3eRvLXJe8gpVthfytPbwzrMeFCSPeQhMZ1
cYopeMO1Zj3ftFQfViGjluhNBH+q7LnAmQM1fbAbVDt104iWVsk9jCynX9/U
0gD7pqgJQZnVX6Bq0XJ0Rwbg1P4TmmeYXFdvCWQYAXdOqQwKKr3RUNoACFPJ
SoZYIkyj10vLsoS4jD4N5hA63YALxsP4OaKQZHfYfbAucYgmdTU3qCUwA5c9
fYj4Vdi8SKErhoec44+K5n+bYBBQXBZXf0MM3SPKKguaTmMpkqCQf7JERfpN
P7xppoi+1n/OtYoxaeTCyMgETrkM5GI+6s/abv1/XRhktYzE4Gg+6hujeyjz
+zqS6AT6h5DhQ1ElXjO8QZoDFLXjWPTLvrS0k0kKfA6og9i7t26NSSl+q8eR
5+7tEnVNUyO3ZI9x22TOT4Sd8PPTFO/3Y6P4pkppQGBWK63EgvCgXo4q39ZG
DyCrfQiIx80CluCozmOyBi0dDnM+iVfnEgQmsY+UpYNZMd6JpJUu8P7Bftbu
+q0hrWD6b4Tm0bnB3jh656q+oTsTe4216PnTDP2Hw8gNI9NCVHXODoPb/VH2
oOkzuS0uF4HP9zxs1I8IT5zuA8SdoSH4QlsNZB6ll57+D0hAj+c+JAMid2Wh
xIp6h8ZyUCdDAPUWFSRCvVdSA0W4IkQTkBqVvO1JAZhrOzy2XPT0Kh6IL91c
URECcmvKxzw7X1UfFxiZqdKzoh7kYeEzlPZtrqH4VxIoVvb8FR/DEBykdqgR
SG5vQtaCd1ub+vpwmVTKI0WtE6IaA5aoFaiP/fr2nzUOYWrCSGbKpfRS13c/
HJqcKW0noiE/k+RmavJzsUt1aMUC4SOEqDpI3VeaXVehPP4KoJ8NoA1OTYrs
2RSFlf2E4+e+kLqU5BrQlWhKjQ6bhxwvpJepkp+iOKfvcjPBUyuNavxVOyks
ZK4DHIfCXTzvKvqJhvSEGQ9mi/IH9JAvsznJbQ1nHkXr0HXny1XbljXuTWSL
NNRHTe6wLPRv/gXD29V+9XeCBRHVWzch9K/OLvuM8/XjM9e+It/v78FOMlFU
E14jztDPBwvqjSVlpd88zpWJ3E0RN0FQ9pbO2a7kgeQkuGfbKypCk3QDBVQS
ZR/ztxJX/Bzr2IZtWO9cC+NbEwNWkgGKIDLqOtwznv/YYXC6YBJ0eHOGeUKI
UYY8Vyxd2oJMK2Pyi6D0Gb4qA4tUgFgvZ5drqr+QzOaEBc/6WEbJJLEkLdv8
iXmA2qEABeEHfChB23qpg3+jKUrSzQDPvVujTml22lCeIYmcWdLJCsbumotM
kx/p0000YrYd4dJNmh+v/57uqVvhkIrgAeglwZvsgqzvepoPUgl9Ll7bXkwf
8dZ2/9Zg2Q4ByyFwKyEGmB6/3ZQiP4pftXcrOG/wLJTxi0R4Si1vaZdWLmjb
O8ougcsgawMgKE8OHZmTNp2rCWfcK83fzKxZwuAX0V4s0SG+/b/4Etrlmo3b
77gpY7+TLtM7ajIUDdC9xA7ZhExwolWMEEdklPQ9yE/RLn7h9xnGPnybHH4s
M10HEMpKzTGABAkEYjttX3G0i0MYVO0x9OYPRDtYqTzkRwtXnYAjGpHon9yd
6X0hDAVy9pHbcGrRonTm9IEXmm5Uslzw9i3uXl6yLTzm4ygh0oqIraTrw4uQ
9p4878BDICPS2EDehHm5ONUfvpwBIGeU7njGSKqJLMOmk9FRM7T7GM9Ds/3W
0iREK540jDBBiF3jJ75jvfuG7TOUNdosHioe12DP0R9FxouFPnbIM44tjcV6
lBJ0YqEiPgQABUbpsmwqbCkIsI+g6/8d2x5TyRKkTjAFCbPdZ84IDs1kicaN
vQH5pkW3Y7c/LTZFI3affy6u3UILtGlsRDgk9fLKfZiQz6/BUxMdJ7rCvv+y
0HwtphJ/Wd4JSu7Sb5U8yTB7WWc2v3JN+pBli5UYb6yww/l2VbUjRK7Mx9sE
8TcWpktejj2BcyYZZy/KlBI07ebD0IG6y3DZW8Ewcl22zXUJY5ebZyjt2rUi
2Ema/BQMzsgmg0pOjZ4uV4Vf44dKkAyNnr/4cTTMfVHYd1PoWYpYyKmKQN5c
F7BLW8zu3ueylQZPn/YgUhT17drX/jlcmVaUlHUQwWaRP9xCrkbAwZmPoisg
SCO/bK2hMfgyDEmfk1wdR6n4JVcMuTTnHWeMLDtLMj9nL5pARAVcqoFAHZq9
A1IZO7RIoUrIJpx0a78fLtm7jEx2gTpGahJnE3mUMGwHuj3tHIeh1UJ1FXG5
BVak4099mE4M8GAt7KDUKeOoTJJoXJ1HS/lN8WJNPZCrg2d41Ml1x6w+hKlt
3JUhTkCekwuMsnF4F0RPvqi0dgv7q54DjvR+U2pLAvlsMYN5YENYsW2Cg1CS
zmPT+UdFlToqM5Ksp5+fCZC9rcap/kvt3EODAAHPy7crHj0578wXuohiBjFQ
nVqWQLV3K1ppWwlo3jDBAcdEkU4IXQcssDbTuDYYSQ/dv99NfRyu/b4AGUCw
GL2Be5N/IvJPFjJRoTqQ2Y6dvLq+eOTaVUVn0y9qdtT0wMPqDuT9PR+xFBah
KaMAZ6QXqlpi0YVGWHugULW/qkQmxViikid5oNel/tDhcMZc1h1W/POaaL1B
YSShIkDsN46D4gLchDIJZTDz5CRpXKiF1z7Uj7MThqHE503xDoVp19FGDqUL
95Jzt36xFat75ubFjfI7j9M3A+d8qL0DEpQ376Cu5nCWoCoCTcWhLj7t0Rch
8ltSkEb9tfxqkYBMAW5LMKRpq5352gdZLi1pTiVI588UqtIRhYNfcX2vu/yb
8gwNfC80Pj+NzuANQd9xaG26tN9jn079ZF/cTc+DjccnfhRELVyjvV1D8hNB
UcFcGSZdKaqV9s4s1GNOogsa+zSiKGyG5BjJ2UHsy45yOwhxEkq6xbxe8Duv
fPiAubba8Fv+bLPCqK9KRsORoh/acAIQppFkCkQ422V/tJSG1R7aoNoydMiv
lORd1a8wZK3b9t3lNEeA6+Px/pJ1cKA87wACQxGQLVAuImNP6O5uSVTazNyU
oYbiICXAIT+0lQyr55zBBlL7tCU+Re9yFGLB6xKlNnrl9ozb6nyZJBLkrY35
IVMvz4/QZ8QHuvpUzrxx5Kf/AU3jjbaWqkpClEguYM7f1NojPwtcfFawca3o
/SMmBzWJkSPP6Yw68eMZtV55LirK9IUqp5bE/Y7oRkZEJYNQxmHLQojhvMAe
OeGYkNvuNJDi9kbbLzYvP1oKGHBwHaQgcwVm0+wMGnsPOLNZnuqURjeyD1ta
htwVfy72tAF2zM6mYQXTV5Q6+gKuObKx2ezXalsXkkPbBr2xEU4+BSoWRKHd
O89/ei9J4sHlcwuJDN5QrIOvdnJ9rsmF3MZn1FbYk5RMa2xdNn92PoAHcF+Q
JTkF7ZuN5yGWn8ZGSYXzZ9cTkkZKpX2QoT6YGyq/BLgEqkJOqCBtZK5iPwF3
amsgJ6JyFJAxu3nkLlpIKU/N52uV5iSc6YR6+qQFXoVL03znqMAB9CVMXt4F
Ll8qDz7x7mmszBap1T5qvXZVuxOFPL9aPacp+K3gn90CHk0DrcoKh9djET2V
gY7AE7nCcsSbpz/+rRwOAzDccMWkWMWeu+LjAq6/pmZ7VMzqZMSTTxFY2LUw
D0D/Nurq2iJ6qOfOhsb2F6JapOVqQPUtSlUnf1H5g2nC+fsEFBo6tO7s5enP
PCnsVFxF208v3FzOJ3NCz7GYMYIEb1Q1KITNb4RtowJuDEgkIxAj5TP2whAr
UqbddgkEun72cGd22UdRtvqMSkUTox6UbnhjRo4TmCHFvfkU2TX0mE+/w/sm
R2QlU5xQBmQTHBmlvX1PGSJSzd823CXI6ZC8NhO7F1a6+/vNXjfC4zK2QTuR
8V6pupqFpyDnNl90du9L0zPzZhaLduy5V+5QqX9YON9HiJ3gHxNA5jJZbk5Y
CKbohrvJvoKbxAMnxSoFKX+BSVVAY5ddK5TjTeKF0TisWBhtgUTGXLnLSIMR
vQjbkN48INkfTib4O7Mn+g/whyF/Oa9MKNaGjWWXu1vHa8sOIZem/OsMyn7q
EOy6FUKVVZTZeqqFuuUf/jV7SpMYz9GG5x6eJsPULwz9yCIhupQfvjZTgXmD
UEEHIYd79Ao9jNX+Cji9qz88rFmAY5cVNjt/oyuJwSpU38O7XupjEMGqiZv3
lOPJuf6mEKYsBCuuJo+cNb6NVU2SH2u049gISyG06Zb5Zh46eyJ6GVOBCh9L
9iB+BRmFg0FA9lZDn+qN5ZLbwlHalgGMFVdeiEXjZtEy+Fh56tm6rjdmgjZ0
iobJ32+XtU1BJObg+k9/Nson/4hUO7iCkEmb+XgzmnH9DPpxUsCHyEA4aYRy
eGLXH9/SZ/Wq0qyGC8iVtKdM6Ll7BeyGWnCCFNaFHlZQhFh/MqHIPGKQYPPk
7DSSwG7cFQG5Mqr749+XEQE/jxr4jg4d9gdtQ3nC6dokpYPPItfGSms94l0S
Kp65O5Umlsa4jck3VCIXIvED6ZCeCty8ped1EDV+yTugLMmSxbM/MI/q13iQ
K7uXl6NF4yhZvx9eoaR43cQAZjL2umaW8WlX/fJKgxagpyj+x2pEy1462lYO
ZQiVl/muJcKO3DZjbKhQSIDN5R44jrDmSeTW4+f47kslExynlJNUWU6noykB
2ZhQRgEf6sRAGmknYVzZn0t494pjeMKQtH/+3/xAFIFS1K1buxKy+G7jTmKT
76bcTr4lcEt2mNPLt4Qt4/4JPeMousq3Xx/O91cL8urJiOG/I6XafEpbuCBX
sysNxI+z451me8FSCGk2eDla4ZAEOme4ZAnvhGlF5WicXnwLIn3b/LCtPVmM
vhSe8a6eBenynW4sSX0fOwQ4QsEHpVRrxMzjy5u+ZXDRnxmXL1qv+WcBsZ17
a58lRVmUXuohHZKV/ieUemb1GBhNmc7ajsupdkts63xNLsKTTRNKtOYtTINf
8ax6AvI4w9FDeo2P7nVBj0VvV/p3pNnaWGklTBsXKx+EQhukb26qF7k4sgJ+
lewDe9T51rSz5cuVzqZ+5ZrMvJRiFWoKURljzbpvv0rgPo9DkFDLIjfx1Nbn
elnUSLl63hSOh3SSgsRz2c7epgfi4ZvteNrDs9Gex9l+LNxYtFFU9XHrOp/V
MH0TIgIQZmQOjbHOGCtLrFhsAtS6biGfpn7haPFI3cCwDkv/rpx9fy7dvwYq
8Bw7PmQksu0M9TfKQJsLFCGTW1B68wkZCpORvCogrqGEIPe4GHhUhOXNo8jz
yflpt/WMsaiiQedl98qekWpvxhpsbXCO9iLHRYMUlAfOGori/9lbtpviswMX
6XxbGcytAs+0YZwFeQP+hyk3H6Fai6E0gkSwyTYO09Q0K2NNEW0VEfUWXn65
aLnQvxgEVqPOF88SNAJnhctHu2kpzs4IP0N+VMmHVMFQpqChnt3zWdGrM9pA
D7fgjbbkg6oLmk7O0SAjPuSemjQM8Ivum+fyz09HCFbnzKjiEIGgcUo68wws
digmz6+2bUkaCxffQemCweP6If8XaBxBJ7Atc+xkYsQRxE8GBRt7OuwnqX2K
ro07DqwmWD47sBvM6v1kek3wTt6kYvshewys42YnacAM2e2Y57QRXsKPyqyM
R8TK58oTKRoLIvh+mhjSy81qPyMpHJrfMV/90eIOQsXortajRyT3rARtuIna
YUbNDXHoTiXciyGlmxUNdWwoa9zUwYeC8vZOPWOI1HEza1sGtzWPQi5FkuDi
jNNk9LJVbAiJVuXNMrAKAQwbdOqZgAgHO9NIGAiqPRPwCzZpkd2FGn0Ew1GX
mnxqPoNMQ+tKrg7xL9CxcPpn+vOb+6mbHMuTKrVsCe6Ug3jBhFlyxe8AoWbh
6slEvsCD/guJOIsqQU+BOqgnyyu0qbJau1pXq7PEJdrG8lZGMcrnukgtg2eh
1JHcRI9WbTnUQdEfyhiIi8sF4JHZ59nzHB76BV3rYP3PMl47wKddzsM/zbTb
sqnrh3lEioyQxhY3qkzpdZbhmzi9NRrEFprORjo8LngFmDwd/GUJJyLNMtsC
jRiksi86Xfh+BZFlIj4j/XNAv7dQ8U1Uhgc6rXhDQzPGL+dqtpXUNQfGNjC8
cyk1RG2yhXZmcNILUv9JkdzhnvfC6rWRFUSmwrmm3FcsNgKS0NOVw7gVUpoI
+kGL1JNIC0wKlWVzw3cTInuhl6ar0SBEQSl9vE+jBS8MF59FUNwMQENH9nku
pEWLjNNygs5e7t+3vBMRXMp1pXCMHvI++Ju7vgW7i79HOQWHB5cB4EZmM2iU
CFGAI8lpzbfU9xF7BYBJI5WYDKXtm/IxJOzfmOe0L5Ip3p/JGfVpfHcC+YRm
UmD6LcOnYBu2531weMTzc16oep6cnoY1G+o3VQjm7e/66p2cWruRxh3l9MEs
bNSVk3hlmArHh89Fw6+hIsvNtiJRAbCyPAyEmlKvu80/Eb2dD5RLXO+CP99W
NGo4SJNZm+a65zIZEpcUWKvfzky1+ehTXBNippUUAgQ13S5rUpBN1+Gh/CJc
hKxW69vElfJQFj8itiQpuG6r/1HXr7aCYKHklvTX80cFXq97MN+uY0wM+64D
rKb7AMM7fKd/foI9g+RH+RLsdqK0QFTyQ7JnKeiuCt2vcoTC4dDoEgSV7+qI
eKIAl0tci+0uROPBIRv/7iRX5sowIqNXG2YpC4Nte0guEHF9xlGuiW9dBofy
7b/HdIC4b2aQk40u1VTJwx0fh0vCMyexMkifEkc0ZbqgWDmbeJ3kIald5dJQ
/SE1NQK0uIigIt+CJK1e98u9HXTk4KuRL2rv4xaPp+pXsp7nEZ3RTHMFdXRy
nROECTfWnp3VwtrspwMvLf4BlpfM816xkmIGfqQ8qpXPog7ZpBCH1Z4Rb3p5
YpdO2gw8o6kSKWZZ/PQ2FG+ZoVnL0mT6zTawTo4UsvXyVb8zt2oC4IcrRKyH
2z1uxkPro9f4aBQwZKE8ZGPjP+JUedSd3do+0Dy3BXyZsDEQ/Yk7U6CuiYR9
IDcpFSv7Dema1i5+tAA1c8Em1nMVE8ALY+7MjwHQicmSLxlkW+Cc/IFTTuYB
iAkPiqmmJp95z8eMze5SzPk7eVaUU2wM3BuILRxAI854THR91FDGZxENrObK
5DaNbIOu4FGYtCoLVB6uLkrOdpeUEeAgTOJVSlR76ASAAYNb0DScdD4lDonr
MSn1GCa0ry+Zj3qovJQg9c1laWnV6WRnAbVb+7D1n72eoZe07wZuqIniAlDy
vl9WUZahAAHcY9Mb0XEGvkpQtniQYlk1SbuVkX+lmX2zwKwVqAL3XUBT2GzI
uIhJiL2QtH97KOXxcmvh+J/GW6FNPkeIWSYomKqP2i06tzNXlJDBizncwG7s
CJZgCFSkjh22ZPuGgUPRzpGDNudkjqG9WyLOmtsFphMgHJYM1/mA9rXagtOy
UApvMiLB+DCjMeqqe45ykObbRoDOrVgmR+e4aHXNlenRwfjeaDZ6+BbuJwRS
KAso2f/dT80En9sLPoN/kIxwFIohBIpX2eZfFlcqq+iLvwpYAkG+SdC/jLfv
hK+0LkJacNaKF1i9aUnJ4DyYZfk+94c4ehv+YZ8E9LNMPv/z+/MwE5goESMD
FJDF3YpqgJ3dfjTFBqe7U/gFna5ffOpu9kgRwqIhfoMdAeTVqPUsV3op5zzP
RnwYgNGGbCs+0MX+OnKXcb9e9OPkVXfZfbhBLGgPcC5TP2Npm7dYK0M7JeOg
0dIsSlJL45SCBfEaTDiSixWj/h+9frIg5jg2EYzTwUBYUaxnQ1uV2GoZyLjb
fnpoqf7EPxWEZGy/OVi2QH+dXuvmdBjhFOVWsdM3kpoPWgMYspXrgT3kz5jl
aSnIqQs1HdGhsJ8TFZDV1uM7qkasX0gYx1RS4aa6sAqr+ECvU7QEqkzacX5N
Dkk6c8nZPLxSpEhligSmASpvwYBm1QF4tdOs59SqjlrWhgoV2Nm9XF42RUTl
BD2s9lKT6lJbGLCQpfBUB9kea8FFibl1+UFuaLVBYrM+uhxR6bKOD89fWISz
NC0sv4H/ky+LacltRutThz7JE4uab4Cr6s0ncGqieU78UBOonnZ657tBd05F
Ien3RNlZbK+tu7F67tKOQjNXX+5SWp6Kn8UaBACvq78XbUS5FYFRIYesMIzA
/jvkL3sl5W5FhEp1tDe1FIdDaELq0fsJAZz+RJNufy1s5rRINIZ4QzPOReCx
EYh6Soac82t8/p1DaGjEyznrDWGclIqOFVcDzbcQdOIAoLWkls3RBnsKyhW7
OlLRDWqwEU58hzKGcnoccvzyjm0GBgowa3CSZJ/lQDWk3Kzab1wSVPV8NW0N
rn80oCFE+2l+SCjpZujNHRYxxYMrmJGApty2AJ9Bt3Qbfx1c08x75TdfkaWI
YEmSvaDblI4gRCS9/PoROdXdHcsrlFCpv4X4gn//ErupIavLauciZYtJgsud
pnMXP4NCIcXRoFrwOXz1nWWLWX3nMQxv38kLdFI1vfomHylDX6I3sJeyGSka
6ClS93iuJJUEIW8VpacvGtQRTrfEryQNAWXMefXIyG/44SpXNgzfebbMwnXd
Q4WrSuE+nR1Hz0ZAlZMOTzw8DgKsGK+DSm8xZO4YSwICqxqP14g8os2iLwxW
Gw9DoNRYirpdwj6Aj4XPobk4DdUImyH2imRaGcv2wXy4qLNRTOb/v9QF2ADP
/3cJDOnRgH5JqCAXkLvoMyvwZcDUVN4ysumxvOfYM5HUATrQ+FI0odaJELyM
M6X8N6bdyGcSrKRfj14ZCHUXptMwKAzKTGOcwNlbgdc6vIAeyIKcoOEf2R0/
LkGoFvLdp2RUTFC1hfd8NJHRSLIpGl4UCNcsKxzPAJhAkf+i7jQzAGdRFaQs
LO97uFPfLKWBoYQNB9fiayudfeyZCDKR3wTsQ6Nr7lgxqM3TEdpacEUh4rXb
vyXkX5i/ZbbnwQtfWKiU6cFLOQz6l8PWYWg79qhiwYs9x4iIOgwDAIzteqeH
iGT105eQMec11S34yq7klUGK2S1k7IwNCk2w0Panbtd3vQoYWrqix1X/njDx
Tb8b8Mhyex52rVDM/7e6RpTOon39QN3WiEDckgrZfu+DG5hnkDFmWG1iZ2j+
cWXZ8M6ou9a1EQxqs6cNHE4N22AruiPHrxpuivkHDeiWiQTO2UWdwyEQV2fX
2GqAfbxiZiLaPphtz7otXW50ap8gNdIyZmHcmZFkLzRzvyyrxTj91zy2I/AL
DWRyLCzUJAjgrqwKdMaEZFTZ6AzNt3YVC8hsnwD8OXYtcCP9qmn7qmDy8r9b
2/UGugoij9biDXHFDJVGQd7rUkHz9Mrr1xgLrnnS+BEJElp9HnLOuWdl+Dfi
2mTOJhP3w5FCS5lEyMMITBVOwYx+gsdf73FD8uPH4tmiFpTfTtkdxmntyztD
T7K6izG/XMhcdJ5eLwdQQRXQ6Z7EiSrh+d03GdTIu+8i0PSWvWQ3yzsTz8cz
/BJzu5yt77NaqmKR/rc/om6Qo4HMNwruqihyFc5eHvZsn32mmD2ygkPE+qqw
ja2S0kH3cvFDjoUPa8q+6+wq8oEST6sWBo8bmVhgacktlf+OAiAJ2oOguW6G
6j+tMOdJDo2C3JaFgJT3MTVEZHOMKLc0u/BVgWvdmiESWBsS8jtQ2SRhcle1
OdzbuDjzWY1u95Vz5/u3yLNgsu3K6PV7SbZVGTILcdiXNXReVZ1L4UGYXrjH
HNmn6mObrvnxIu6oPUYvjY61sGG0pTGUIf49yyOmjxxw74aM5Z6ZeVCp+R7+
/1yka2wPqT2qOrzFBtKpaUeL4ZSLU4IpUD28Mq55daGmU8zviTItSj6YAbmv
vLg5RY5LxvX3rqanVjd3eABw3qss2AqG+qo=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGN/U5bAoIiu9g2EU+rplkupeJ8FKFQ7qYul9Jut1HrG8KYcClCaowV0xqzhdPy7nvlERCXCDQTmWuUAuej8M81N5/O6g43hhFBIorB7dqQQW8xhOoJ7ZbB45xdnFE8qZP1nsy2yJ49ouDO+T6dBsEavBBmPzYnTo+rqAEqRVR3PaHkboFPNqUhhNHDMs8emBFpdbSr8uPs2ID7z0uEGmHZKOtbf5oaKe26q/45pNXikESMMxUWN28hEDHRA+osL+o3mgsquCOjjOU6OujJ2BMYSCqtVs4fbkjuXd/lv6DDJfEISOniV2TUjlSyzJooUulstpmGLVk4v+ZfXi4t0MIZnUJwYHE+Y13p4Dbj8AVVCUNDIaZFFJdDitQl5U9boPv49IJLJyPrNn1dHcDVvH7nTTdHfqy5go2lCkrs70XgBIA8vPrv8P/5WrTXjhf/G3/bO8GfGU/VtCc1+cXD7DpB5ot/vDMtBlPgVrZ2J2XFwA0d5kNBUgOov9xXJOuuVpg1YjY7dv9OcImkpuSiSjOgXn7HOM5175P9hLE9IhPzz7Dw833kF32Zw0LYvMvphjADalvRpYlXPRMjbKANiohJonOaQ0puwctVVfjPIRMgVvFXcWy9yHONY55F/12qdNk33c9WFiXWb7muGUAz0MtfQ3Ap4+R/uLMjSjJZ3RfiZ+AvaKYEXYxbllehpkur7dIrhVRTFSvH8XtQdu+A4IikqlWrBGzaXbgQyJzS3DG8fF1qrzDUoZNFjfWG9edGqX1xRddG0TaVTrE6JM1ojfCKa"
`endif