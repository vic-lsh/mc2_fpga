// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PVoCYoUxPV4eRCH3b+VKgMM4YkH/3ILWJxBRD7c+gwQ/fT4DZzGH/L3xYC2c
nrNlc+GCGqw2i43ht/biXAJKUzxsvxXDY7xW4s9TMll/GM6Kev/4+mBrf1NQ
ZdBy3cKzeweq64jE+7WLN5opEP/eA00EaNdbQi5xLusO6k/pWO4qyBim6NiO
t8OQ5AGI7xUuui1q+vZwZp0e26Nzc0Rbjek785tGcetK59+Dihdu+V5UNmX0
4SdIP+04X8LKUzfPI/5RvmIOh8FjAPXj2lN5gMT7OOO8DHMArrn79tjGODHA
wGmA/6VntsGQYNM0g3iZ6cLIIknfdElO3acLFM64kA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bqVzcD340J4oZZjBakXzlMxXd5fQzfIovPjs/wKGak0TxK/NOwbJvBtODhjG
LiWlrI54wgXUQ/u9snFCGi389puexH8LfGKxS9wU6qSIKOM2ydqtTToYcAts
SZuiB92/GhS8+gQEcfqb1tlHaKV86KN4WDgaK1rG3ktaXCZrqU49aeF9JVcQ
Iu7zyYksmNdOez8cHQVjU+ZbEmqQRqOjWjTa7+dUhHdKM+apGuIJWzS4g1Q5
X0UYL2LVicCk7Su/HAo95AGmT991yyI4ZFqBkPg4pjuHxxMfWC+/e4X3dpUs
QbsOE0sRnjqwcHSxsl5g8se+CIs0+G2lEHQFtQi1PQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IFqCki8ITcKk2Mptn7ewXEHckczNWgT/geexF3B+h/QMcRmdVL4j7jKevb2o
QnX1ikZVZAVVSO8traQ2JRmzDrEE9iQyTZjAb9/mLoPxRfyFMwp/PcQk0ShA
J3HJpKofxsvahfYLGwvpyX4GxIxKLdOCdsKOazRw2V1IdaEG+pdTE1fhNz1S
jMPyvvh3F0lzrRkkiwNuP2sC+Mdp+jkhVcDEcq8WGxtIwksWKrdE+52w/tT1
jK9MvhVu1bTyMeM04Ruyv3Ggv+Dydmub9ghnRtC+TEo8h9y1MfL9+NtfzYqd
u62jO8U2inztYYdRJ9dfa7DgcWTI34dUL8nDKt0ZGA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qeR+NLkyn3hHnjeJ7g11oBBaUj2UAY9gWi9Yok3EayhGQdWSu8l8Ms4TSdyx
cZBeIcdCwA//qolOQsWqTplKJeAFzBv2rtB5BlP9GOVquLM6Ydjg15hkUSfJ
vPdZ0o1wSAulMql1EjKwaQvfnNX1zvX+4PTyWPrARW6S375VH5Hr3ASyPkUH
crZ6+502dXRRjCeHzbh9Q44I2owgHre3ppIjpyABZ9i9VXEnZ246IwG2ZRly
6sCMGL9cWyJbliVrzhW9TtPVwTb5FU4Lg3X7IySOOCUZ/Xtojn8T9nyBo+wz
BqasdArr3TV5irupTyouVIrWLRdbQsA7ZHE6g16EcQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WdBCGUfZaJkF267LGjKTOY9Fx3aI0J9VEJR+NmNejjF92hLnjgpvD+GWqzJV
FW69pZ+8UyDxGSBQaUD65caECwNUFIcD7EyjJAOzLXNH50D4KRPCO4m1PWRU
v60v4FsTI+/qXGDEaAIJVXMS4yDK28OyVvK3eQCsxRpFVd0umkY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G+Y22PHQXVzpp2fynmz+ZCG+cC8Yt2XBPSTzV+y9UwW1HsiFXicq3UwMYyBm
7YUwyceUDSPG4pVWXbWqJzT4WmkGVGemrtyLke+n1pRxLaX4CIsncHL6eCA5
TGebnZPHKAaB7RckVfopeVMa52Q4Gv0+6VFEFmNLm7olPKoUeIzHSaAuoww6
DXn80hoK8itCerFKYYViEhGKRxREL/7Xq6SRuNaJ1bbi7/r90iQI5mJAtDom
yCVO8wde8k1/qqK3AkmLq2MqwuEQX4TQabWWKRqH2ibHvRXoWoQ+FDFLcUFG
Mq1vXZkon7Qjl/xSoB5FI4Jrs5MDtmKLFihui4r2Fy+0qjNRKiDPEiWHjHkR
ZUwOF9IEJ+WJxRGNn4SPS7HxRkfP+0+j4un7LcLADCEhI6bV+rkEfF65eNrg
naypr+bwUqz2AXS5jwQ2bKqJC2RNohny4rWCTMVFLX7FhIij2orq3z7aLsCW
hnQ82in31P7TEOzj8pnEc7rp2wW90SPa


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K3y5v3GLtAfR2FwZ37xJcfCjs5ibQKieI6qF9ydcGcJ2tXwAMPqqw9NYMgtQ
DgB8Onc66TRDYBhT/bnjmqSzZokuI8Bw9/J6zgnw5KrSWCDkCudcf6x6SMzv
vnQ+DG/W4o3ox7E8JoviyJ0G34T2tKrXNDdmGPxgqesnrNeq8w0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OtS7lc21wZcxE/x7Lml4ck+Lr2HUHJdajUHs1cBi/BdIWD1JIzjhofBMm8Nc
h4kUjNFJPz0Yicu6jPVFKGkXex3ayzuctxPGdJGxB+o2xTwEZn1U2IdFoXrj
pkXpcDyy7mK6CVkUhOBAHjQltyjseUnU8NJjcocwQ2EXzGL5+o0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91936)
`pragma protect data_block
zZvLzXFhlyuRRHgvMvRVqIxlYufozQNdKiNxSAGpTKaJYMaPZ7gcd7B8VUW3
DjSfqVaK8lMvB/S2Q4FlOKg7mWR2GFG7u0y+DB5xSsPOXgo1gqlbAGhZvYUz
iK1p0beE5BMSgxe3i4esdlgEEIL9I79yVlem0QXFcY/GxfT/vIVx26TAq5xk
HHYJme/XNiwjlCoQ4J1jnjgqrtWvTDt8GPvYjShK1Ke7r5kLNHfojuYi6otp
12VcCg46WSKWf1kxbKTWUIHrUV4LQeJyMd4mAVUa2HIYlWgkl3EEPyzvrsC8
D+aVAfQ2nNsU07TUHhxItTelbyAK89ScnN9ZZAMEZLSq0kZJcIoOWEfJtwoT
VqG9xglVMRWHgaoe7vLccicMWYNX6tJeCvPZEs04EIOQ3iZhS2cwHYfVeUzC
vHVD7/rMAJqdRaXSBKsvFjC4nN0KiuR3v+KE6VonsaTTqK+wlHGq+/Jia3v7
V8Bl39Ld/MmB8WNLB7q+4jrp5zgBozsXpZMMapSK0UKxhxN/7NA8h9937jTD
PkYLZt3Uq4aGnzAeBuh3Ew53+CxTDLfZXfDY9P8C1iuXfkLm2nr1c959SL6h
JUJy6KhtDuxOkflB09ReF7NvPd3h2qWeU18tv7ut/uRHFGoyzrlkkC/jymBV
ZtmtqjFIky1/2qPZUwNCjRANLgqeBBl20Goxyh8tPm4rWqGEQnDkUwozwYpg
4CV32YMoEQF6pqo0IVyvX8sL4oyBxdTzTno3O5gtF/aCUWYgVHHRLpBML6Qh
EYC1oOB9peqlVxcUOY9OEylRghQifGK46O8o7iwvaZEG8pIz+L64wrXCBjLs
YW5kg/Anp4cTnOmJt8LR/yp54zRgGkApxKZgNkuqmpGJ5oYj8hwQnWvwF0Lw
tTNYaIZ8iwqhRLjpbbYcKNKgKHBqkx9SX94kK/eKF+QJSj0H0R6Fx1MD6Rf/
RARrCEy9R+X9hYvPoT1ySnlw4tGNxr+wWQ+3z/wev/hOnp419vTpv1JarWOR
z8Jn9kpDRzXKfRcdw5PP5jKNHbhiKT7rnsqpl4/R42XGmHlhxgFZN3dzSBsE
oosDH+wqcQCelFOKFhLwH4OVp99Z44eQYgmVVbrsmjHLXxg9UORQpH4EhnQx
MjIOzn0h+NSP8lbgMI0LMvgL27LHtLSya0fi4LkmbbM2IhWEGTsLkDDkTIXE
DSF18Lt/22tz84Ahr9vdOvGsSnewMy2yRJpyxMlZThwgxD9HzkHR9RVsuCT/
hjBvFz5pAuSjSDGp4pamfxcOzalcIsGZNGEG48z5KLQT5C51px+wd3+tNLOp
2wIenEWK56ahhiBemh2FeRmhn6gJajmYIcFexWSTyr9U2RGZnFH2LlFlIikU
NoAkKPavb2KbmLS29mOfJpy8bv/RYLyBGTIYZuQf1N4oYnBYfqXKCAx3eRW8
IxxHNTxir1MCAAlPy0qg8zwnjefOZwG+SAEvp3sTlNWO+/2DLgxpBZJk5+wG
K98PX5waE/rAOPtR7AAZQOT2tuykSUsQ23QU0EQlMZimfkdBOpvmwIvDnZOh
xoAbG6vgLLAXJme46mwyDnBsAurbrwosC6YR5PUQrOnxYAJCn64HMrxAdzFJ
NVCfFyii6gjx0AuY0ZeUFPuOVkl/mQ288J9hjvgGU2x5/Hq+CKc0GFsj4C5w
Ke8mlknxXmbnGwc8IKI521xohlnA6FN41wEzRSa0XF+9yDI+MMAz6Q9Q9F/u
L4xqzJdI0Kp4BSL4B7O/J6XUJaWtLZiKS12Ld/rT1tWQUqXyiaZuxLkSs463
WNt8wJHs9I2cJQd9fXBb+kJaMs619mlu4JmD7/aWrZnYvjF8RZqguDqMV0Ng
yZT1GwbZZAKgAcungrelmEJzJjhSW0W6jMO03Nw3NaxtDChr7ODQDbkDlNRS
ZAgdcgASe7HVSsEDYe0qt4wd7iAuhI7ypuwvBlf59Bgvauxc/sTZgoJYtl3v
uoRYDEPQ4DmUb0HBmml7BtS7dee4N1XlljQ9TjtD03vuAKBgzjdDFn44YiX+
7E8P5fqY4pu6+bUe64FLqm63KoQzsi37oi4pVFfMoKPw59/JrH+n6LRdalgl
rdxB8Z6YoGV7yRIHVCUarsQlqKXm3WER5EgXkv9Z4yXbjeOntuLQkIoN9aD/
XNShB032r9Ftkj6q9EGzjU3FtErytEWBSBeSlSN4f8TkzbiLSr2rxETsVpGR
3eZ30fTcTV/KhGddWvw7zsmKupf2WcFaxRvYWpxcyXK4GZNdWUfyPKvoT95t
c/oD3NccO0fvWOh5+UgpMsBl6hs7eRA3n55syHFtACGH+VVjh5PdGSebEEU8
jIJzJdyZgMnK6pC8nOyb8lSbwn2izBFJc0JjwyN4nuxM+IvnPIcSgTVTglxN
x3PJrXno51Fn3fcllJLkp83sanjfRiwk7nUwjBbs+ffEdnJxda4NOjSr4yGb
pkb0fH7sHtnh+ixu0RutWx29m1HO5jz6qz3i2DeCG52Tka8D8O5o0sslaN0Y
SO7lhOjX6pPMf7NweErO5M/zvr2k30qBkKLA3/AEfwWwRM7MacghhgGP2MJJ
MVomCw9iyJHDf9//8hbPFcS5mS9rhSVyRwqnJMVQx0G2K5wfcWBCME3du10F
fzodO+NtQEevYB22vKDJEZ8xKYqhaWvpGddm36JmwIADxoxfx9su/7Pq0k/n
Wc42mfAfNk90NUEn4YjcZQBRrhXhYwfmJXayPtEM67CRsWewu4NL7qZItYRb
tzfkrk+BTma6QJMwAzVwTQTKH6JTiN9/G+FOTiwfgBzAiZTrpM9fy6+jFpqU
f0G66xJRuVzNZIKG5hfoTLAmegAzRWamRUuq55Ve+HbkkfGsiEH5k4YwJc4B
gNrGltPzE5zcWuooWAguQC2LOcZWaYaQoG/fCbjel3hZXLcoA/RZtVhsKIpI
Jc8jxjiTajY+H22wWMZYtYcnlGIt8au7ypswdx2vNsLLPAS11bR51RGeQ9T2
jiuzYkClOuGR7+ZyUEoQnDsDxIbzA4ndyLRSrWyyweb6fmRETetpjhkAgfac
J0CcEtlLgX8lquksJGz2dS9dhh0Luo0rAyIgLVt4PnPBOrfr0rimA7t4Wjfi
rg1arK0CzS01ku+A5pUSD6f9bTHEjjdwbwsRHf0cbVhAOu99laBSY899DwAD
GYf67i8gXTZgMkGAXigG26gMr1Q1vXTB2NITZNmoWbJCc5cxmBZkfSwasLoV
neQGcyDurfODN1sC0fqvS1DEr2V3b0pIZ/DP1N5C3LpANkn6yoy/+5JtR7D6
9UT+Yj71AbjvINYtCGNHF4qarYdw1JdZ+3b7NAA9zknpZAx74XkGjeufuzsu
cunfJoUaYVprH9p43naUV0ve/0Sdfvc8TVUYvTL2W4kj0ftXg6mqlBAhSKlY
TvsMMdBAbF5+pWPuMnekNLHUSLym+3nKTnqWsSit4CuMKr9jOCrDl1SO51go
3I+RWhMgqvKkzcV0TY3U6pcbYvycZXUJpfBBULwhEwgV2m/wIOS2Er3aV7JB
Mcf+hrG8ManPDUnqG0ZEuj9KivZ6Ir9vRWJ6lQbxdftB3laN9BtClOsTxfFN
iyPfKsrKZx0xJtBpQ0BbIU7GJ114tk0CAbB9Mn+U8fHgPYJ3VvWObUBpCco0
9sl59mklN1Jb8f2TzlaPoARo1tNEOfJoYAz8WztXPrcLwfB8VgUcK+Ymrw+m
UBIEPmYU32dSoEaMsbsxaqeBpuy9io3Cyt11NUfp53b0eX9trLmI4ngXWREp
czwNVvGa6g97G4rHJ371yIjH7OQ3joju4tDgteUijfH3GsEetwtsvvWP7xXY
GY6KhvLjyIkrHyhAnfiSN343nB+tMSyQwBZ8GYS8m+DsKC8IpiCeKn7cdOXz
xXOmia2DfrHHRfmwFDba6sg8byHSWnB9XOTDBM997eJ7TyiEsHIGVkDRMcyH
dwSQhEZR39HFYhR7ss11narPFZI9n7MaCJC/Eq6TKIRm0mQkptiE6O6/52dt
pGTn2pfmhPyE1pWR+fEZUiQr/mPwsEA7iEkixLEtcneJvtCiGTmzQrvE1UhJ
2ylMA0XjPl1u9KvaVTK0OTfr0A+2eqnQB76W4Zdnj5UocECCiDbkdiRBxTWi
P7Fv6w7NxMDEyCIthg0wzUhDxuBk5I6naBiItRPE9lyaC1sHInSb76M7bpWg
iem2Kj1sXST+9qNouV/9sfqpo+8Er+jxBafGm/y3DWGJxk9O45SqgCMjmNU9
xrgCbdu4kXBVtuS8YC3QlxhfiqKfAtgMCK9lKnuRqpQbBOkCrDoFpvqdpjyI
v3z2RYO6VEpRYRMpB2SKcQF2DdGszdGizYR32d2xhLfJ896QqHsTYve3NZKr
hlPkBrmGpG4NDAYLB8zq0ajr36NWb1NW4NtQ4vWMnyghs3khm2S4VHLG3m6I
BBk8pnU7oR9HeI5Ruo57iyFg6C2Z2p4+8NMuN+x4rlQ/dWIwMCZnLmnKT0SQ
JHRAL/w6BldU2wLAqCsP80CLcxbl2yUKu3mWuT4Bemxs+rXT9gUIW+EQoIpB
o/1T8swv+QE73teBpmAl9BiYg3B3P/+OjHRxdOxNVocSZC0kP4X8OC3aHr5i
FjLT1wdigY2xV3wssOl5vO5nHRhagS3yi2eeUZSqp1TO5rp3mPhRls4PUZ79
VIndHIUlnEg1uTSo7wwsT6nGhiKaVnjGkYuElru2MRF5xq4PdWPFGfokOob+
bshcO24N05QnPH3upnCkJnJs7e3HdjncGyT86JF7ObvsjYn1ke+CXpLkb9Ec
csZwp5/L07IEd7X3+HzD2QhKrUJSTWCvVbnRe8Dsy0kYe3DbCN9SI2l0peED
mGvrjp65BLGoCGdPp6xx+ovVny8ayef8AAcNsStH1akypupghBwWu0viM5Jn
abo+zsATFEv653iLGSZKlVcI11ss0qvTPc9Yf1AjJgXl/SpQISqOvUuBXsOZ
0IJMmfhiqX47sxvDDQlB+bl63BHg/U6H9cU86US757AsZgKCA5MoU6oxLsYE
IXVCJDvUBfIFvpfsYBwN6PlEpGPLLRit/8DVtvJ6fDrh1ayDMr+s8ZGibZGP
2bwQh7A4+NJs9Mu67CH9s/wCXwbP4+2UI+/fpPkdvvUOCGCaZ9jmazM+nLPz
oF1kqyt4KWc5lb2k1Xdh4AZZqFNZglyjnK5NJsXpvFcBoaSrzEGLhLF8LTZn
ikKq45gE3A9KG5svPqv9N8fTL0NIpGODvyQKWKr0r9PWQMM9dJRR7gm9/2bF
OM+wIR31oYgeHP4BZXhvHeFc6ojKoeLja+6807Bi1+MEuPUxPdDPaWuOlbP+
OaYm8fVBiR0/ZozshaR0mfhVTp5vEI3eC4HwFumoYeVWp3uvuq8xJqmiZBR4
UFLH6FnlzcTl0uwmMirB/MYll0/BHpP8qeHXCK/2Qq5/pfFtaVcXTSZrJuwU
38HSIw7EctAdMeYrU0nJuF/fQy3FzxwQceGje9CtcDt9GN/9v5O33HpOJGBm
6+ap2RBnI/utr8lM8JnhNLBlFetzfVIRfUMtmnHGWqXiprHIKydNxSFGZQ41
OVg93IQcg1yFqTO/aOjeFjWG1V1CBXdW1Y6ot5O7YAz1oCgMmubZ5uuI7/yA
trR8ipWclbol+xC9MyZ5zasAb5+5ZSjE4ZfQlD4GPiudqTxMc6S1sY6su+af
hIqdPFjWNyeswm2EUOucDO6oTbgUDhI5mScQ0YzI8jch9HSpwwKC0ICWUSUQ
7aYCm0HYl0kUK2PzoCTEUFUSYZ1NBAPb2Xbu4kGDb8ywZCwrSo5bZAZMHqTT
Bwor99P2NAdPRoh4tKtTGXMZZ+kZmFxl8sZeoYHh4Gu63vZmXnZnpl6C2p5s
uMvMznFZfsm7lag7OcGW8WpvB3mKBPKwnHFlfV96BIEdOxar4GzI6XpAK5sO
BFYK3AFhdUFdjQ+zhhnqyzwbqog+4SzkdHgwAUBIZQuzFInWsXh+Lc5Rl7L8
ASKJucpCbdlwYM95HrpgoQ0m5xkhTPMHRNy+dSLJRdC39jHDkn6/1lMcAjzM
HAGGajNirSpl+eN8NU9+6GEsImY+zYT7SFB8av08DPxOSkkPAWzAMH0/8wZV
mk71d0Wtxx+pgBpku/b/JmV8sKUNzezxaO9TTMH62dcoiSkYUbaRemrkClR3
9pmwfFKhP9OAVhGwDwXLdIq5Z5UODWD9LMrqSYEjtm8nY5v1q2uNrB7FdOaG
S+jcFlFq5xA7zRx8mtpGuy1qzW+VUvi0eghg4WJ7BAg876xw/duqHC2qv0kA
Pkt8P5C2Qwf3tsRw+s8ATvzbC3EKJr9wljBZ7oLzdBcdCs3wClOk4NjYCWRb
tNljokZ45umQl0lp4KL9WO59x67QHocRzYW6fgx2HpKyJG7sVN48Zbw+fYvM
vu9tzHOgDI/BDK+lyD4t8RcjMmpXktXoxIpoGPMfabV4Tyvtms505ceD8Oy/
iJYlvGpdBrY9Up889e6YOU7VB15ZSMdEuUMomb+gkaeWyMjIhba/hxLHV/SV
FkHskb4zGaMB4aRCMOZQc9WiT8//+PLOBeAU0yeW9WiggnTYVJDOzsPHOSUp
V8xsDVOaR6IL6Qlpj2kijDFzLT6RsfCA9F/tCHopCCRJBiTGkNTiIJ70ehjE
langapQjG6CfUGvh8LWb+lE4xOSFWPQ+ZyQHXesrA1425pdQ0djrX9bwRdcL
An88r2xTtH0jFgFOAXhKOBjmPj4Dac1svjb98e0avxzcxzEd+QMR6UvRMHxb
rI4EVyl/g0nABszQr7pDLLE09iJjP++BJD0jeKHGEEJ0vPn5Eh78vz92lx9R
5yxmZN4HpDmgEuB0kS6odpmg864wFOV29M9lDJKbU/07X+q7yNIHI6BjSb7n
I8zvIGZ22z4YbiXm1rDfZ+D9IOllqtg/b5RMxsCsXMJw1tm9sHFXyMB5fQBy
zLvLTCbMtIrjfmiWTAQLF7G3thfAB9ckaFuiYXIRSvPCXb9gZepvk3l2jdkx
ICe+qrs4ZnIHmA2uqPfrAS/BVe3YfMD08Vlf/geYrFUFKD0JTUzouiylXr1J
Xni0SY1RKr34bnik1CvOEtROCVF2HqoP78HdzzKQY0RJD+llaL/S40zALt25
mMEtB9p99DOf4MnfKY2RtuiIu+Xn0v77lWT+w4oUStPmtmrP0wbpva/JtODd
LE6dpZBHPyBLsSlrqLhkh/sm6qO39NiiMSUMr0CGQcljJ11iDZsa+gFSSKTF
E+aCmV+8NCUV/N3Hz5C60k0LyhAGdxqPW6z6cmdA7f/MIwxamIFr5pGRN+9g
Du5PVQFrAE6g7o7j45KJAkw07X1dy2PjBKbi+0ir6khOzrJ86Jj8LFHJRR6e
rnOnSxT6XQ4K5n98dkfPKmmFjD4+av4aw6YbPmwGcpvD5OK/8e8QA7w9k9MP
M/N2qEp4P9rW82rqFYWZh4QF4NejlxsSsrcKFUPragepfZC8dzawvRzIe7MP
m10P5M8o8+aCpcCSxdbmFdfr6gBBa+AxW7Ev1f75snB7RtmktNZG4WmX4ydH
7aKKKYWrdJu1A6TufWJwPcOCtf4MLcVZn75GqGiR5D3eUAORo4UMD0ZD/Oqz
DVf8+wwewtrmc9K1SS1LhH2pDocQAmM2divc0O1ORpVJBO+vsZOzRK1N/8xj
y17H6Z7qZjw+27su4mRrc4303FawyFcbAP60ESFh9KhiYm8pCGqJBpwnona9
6KSvdceIbi9uzEwpQxuxBF1MFb3dKKD4OaqlEpwlsQSnya3OCAcUtcNijOh6
FULd1LmpKDK9wguHzqQqilUn6PWB9QgCeoiOG0E3qKXoxnpwmcZc1d/Yxd4W
Fyka3pboUvI0ulE+Gl5RuoKx9R9FZv62Ut1A3dTVj2eaA5ncatcSwacFPNuC
OTKCFBrczU3/r+u51OOy8XA7xT/Lc8FPhlZsPLtZNV2fBRh7ze/YrpdL8lZx
a9mnoYGBv/7j5iwSOY8dXmq+rciR7Gi8xVFSjjGFi7Va5sM8qwGZcTURa/cV
uT7nAfXZBnIWGakywhvJm03GaYT6wqgxlaV/pkgaEhOAtK2awBNYzxlNaZ/A
ELRC4HR+oY427yFEgDFwqCXjV+c1M2hFN9D/wAUqATy2wJzm8OyJxQmoLOXm
i4cbR7H7nxkov1+DuWI1nsRUcA3LLvu+fkBBswKcFpFlmGTC5PmsoJKhnSTo
sTflYu5Bq5uvh1pyhrGBXvkoo999+hR43h5UC/hYV+qCGHFNd2HOe9Rc4CAI
sYui/PRdB1H/dO05Uk3PmuJzam00vU8jLZoMW7eRjgm7YJDLEHTZxizuEov6
vlakHZK7IwB6Ldx7CyY+s8tdCYlcnQTPOLiD35MGjU4Si6MBlg4vtObMLCyS
1YtYb83v1nsXsVbkP3Ihl+mAxFkN88cfJICaynyhd4/Th4Gp8peAFMwrHQEB
HCzUCTcjkQTzvnlK62blEoykYTPXlRVGU4r5j9coxt5ztY0LMvdZCrzWcj9w
JpZF7yNRnbGH9QYLsS6hRxaiIAMC7ZsojH4gGJyyo1VwJ5dNkPWwBPxnkmFP
++8b8oYkqUxfjL2keGxdcxENG5W3PzW/4SuKqmgw0GOv6eZUe+3AoN+PyrLa
dO+0UyCQ5arPE2//+KjaYQt7GyI25l4sILkHkbipgRiacv5K7PMPrpukw5Yb
2kCuaR0WSa8AtvPzMx0Y0QbFagq1v1RjlS9NCLmAaKBtKuj7lExtdKAZDbMv
l4/oHuxiBUgWzrpaps5Sn02xASBNvN9z9KFtQV7lma7IlTu4bYHVhzzd8UPZ
N6C4QlCRMq1kSiBIJJesCxNT/WghueK8rf2JJ9AL8jS+nnOfEqglO/wa/9Co
7pxY6lDVd+sdwN8KrsHiNCp8zUHYNyC++9R24CABxs9+DoW1r/6dSD1w1OYt
LWE9BnOKQFsz8OXyHy65010dcX2jAbcgOkhwJ0WKTWUbKaZqvSwrnreRyawk
4DvatqLy1Deu6w38voxuxBaRkU/YZupR8TgqcxL7nNfP7V/oknj7vmWo4te2
BEI0kKgI1liJ+2ZH3/GZ3HisWTWrutJUwpW90doO/5//+ozTFZUd5QHo2Ick
w0yRlcVCx80EZcl+1VfNFFqC5koOqWj4/qbOejbGqBlXsI/ZcxsLAaa16Lph
tOXlVComnGnxhYTxplW0H+4qx4TKHliG9kKmLzEJx3ob1FJM+ZDHw7W0t/9g
/lSOebjiHPsr3y0na8qvg2uLgz1qq2FwpDFUNyIGCbnknkRWkBPCVTVSz2Q3
hHW/pCpPwBdGeZAbMzCkYGS+AcREqFS86n0ujc6GOM1fD3WW7g24VP27VEV6
+CwGNvxCbYKIIiGr1asZRq/xp4XrZUTgXbbJCIN0xCU2km8JpWvsX94wfSTz
i8XWUF6GME+2vV6sHfmkVkkcooEhY7pKsHn7ZKX2SWgjhA6N6bt2e+sO93ho
XONNCM15ZWOSFLgql33f5J3XwDPkOcgL+b6yB4GenmZ6DZacPav448cDEVlu
p7Kiq3cOe4Jdq9MI5RMsccjPfLKTPsqJjggCR9YjRPk4yqJ3/5x8RnQj0Qlr
mNqiBdIfbT6cCNoInG7jxURTeNZ9qifYv0Vo7NoT9/x1Q7UkFoP3ZYpekjx7
1KP79VVbLIKSyZjdW1seRHxg74qOuQnNhLC9/bKLVddPS16Vfl04pbrdMXFF
nzO80H0Tc7RaQOlhLRFi+SI/dDcldGzC4lAUYwPE1f0zRC14NzCuftL0Luno
jCF0EBpymm+kZTB1tXsUipJHlRqHJ7Nm6bPMyCv9fv8wuruMGDYfqvuXtElc
TeSTxGHcJ7VNwu6wUXbl/ioEDR7P7Gnw9lp+1VwHuyuL8BEfcqlr/D44l/Ph
Vol+2m0AphVZtDLnwg08q/Yqa3Y15xGADA8cqlGppyixxeGx/HZdUumB9ZiD
0srjdgk/QeL+p5WB4GkqTCKtfPEg4C7e7JfMyg42Ypprfy2dVoUTQgMebgUZ
dKS5+0ojR1j748wKYwMd49b1IjCzYVAkuV+iHflOBBNXBhXFu72YUqqDAWpa
lKYZLdZM5ZHKdhK5AcZINd8qr1nPfkeegPh+uyI4ZPLCrntuo83GI8srlVST
iwF/rxGIuJZOXh0DJwo8AMgzPMBiFlpmo8bFbEhUOd/kG2TVGYn9ZnXtDbA/
06KW18YjuGSFSI/4CnSIOVWGGts36r7KsUB2o5Yz5y2NkhGdMJha51ZT8Wgm
yEoXzpEslT4Tfb86RJ/2GkEcZobFCjX5x7LFhydUBtdVrFvnSyCjWbmLTS0C
MXEZStzVFDmaznMr6/6qjLnW9+h03CD1Emyj0hxuv/6rw9RRS6gMDXcUd0D0
YmYiNBbok+2Snek/jc3FY3KCfnf7RPN3ho7dVUhSVACtD+BBuCYHqlPKxaem
bGRN9zqtpEkNag46E9ebnt9d33u/3dxYzoUnnevh7ENFVkpiwEHPmDsWlP5C
uALufD7FGcMI5ie7rvOF/YdSV3ZfcMWRHWDzSzDlHtpfTxWCJSCCChwyYlMW
QZX7ErAtzLN01dGsbV1KF1KbBn4mnUwmdo30whjqcYo+NuNXAYEghg6E/h9b
HJ8zWbBLMjuo5rm0o3VYm0bQKM5zo0t6L2jipQCIfRgO8F2Ca3wKdqRO3X2p
4lExms5k6T0VklI13fzlxu0sS3JgwasxXxhBqGgoPuWEpOQe+jRBm5MHsIQu
xHW7I3Alwqn9iJmyxLkUlcxWvd71QHt+CRFPW7c1cuJh/T85LQLYqxvJnnqb
G8eOZuXOpzD6bn5HIiP5qV5PAKZgB6abWjz03vzLELWSRF2U056qejoMALR8
Hz9U4VDcWW8jFK4mqA4sxgT1wDxFIOZO0jekBx+93+vV8v3G07j+4S864zGE
/DlacyUULwK0pO5Z2p2Waf/ARxcmBctNSgjUWrOsW2DbvruexD0Opm0+9MWW
1ourjETjATPq4iZ2k89WYwF6Sssdy1JhOIcX/Jaev2hq4KsGhmsW8lVKFV4r
5K7CQ+ZfkzpWhAOM+PabEJxCK77o2B43KHEnvgAt6XRLlxK52Zzr9U1ifxx5
vly/2x+641mR1f9oJxLMAwcmBxS+JeOQOKlka6LdexuDijBNAuBHvvQslB04
vbrHr+/+t5TJIq9ojxoJPoBoBli8t/rrvmogSzqj4Jo+0B8tD8rzCHzVEN4n
slovGjnlZH2NSTieAStrIlrkBNWumRj4Yk1ujV20CF0MTsJPt/ceCeGmUCKY
32ELqhj3NbYdA1CP2YTCGIEw4bSRlqdgDcww0yrUpzTpEwtpecN8rwrIV7q9
rByujbUxLAmfHyLU0AjDUl2gjLrVlhPUaI2KtwkBMiRMtQLWY+fbWoXlaMje
ysctxDX/1u7XX+ZTpItL+AyXbjL3ogSqDhM/eiOzL6pOVwRPTb+Jhrv+MovL
xHGM+HA3b/D6iGzdiMYpPWpqkKqYQZeiYBkUIxpLfz13o4E++iotOhQcVSJn
lbb87qIzeiZmL3y6uu8hQ/fFmy6nC8SPgTX8q59Co1rLe5CYRH68M8Qudij9
0HeSw4+ckSulSh8cAzZyr2Zm6J5GZKb56zYiaa73ZKAOcduIzl+rVPEmUo7K
j2KYnjSyZlPsryZF9wR+4cAWHMQGbX6snArwu8kPTWa2jcpSBedsrOUhmF6E
PEekY8w8tSYoLE8HdLjyUDFhXCO+4YqNWPboBafjt9uGP/hriewZCJN/pCUT
6mNPywG0kAuqdTIlUcICAk7q/lFQbXqoMpOyU+pprxx4zvnVfFhicXi9fsNH
enrlfTTMXStyCmk1PYEIkyI1m6X4TfXb3ZQJViV3qaeqjMFDPgaJimghmc0h
kKvu2nxCjReiEAAFg77B8yY+fZWUDi8vOgyxgpHP91lajeiPS2bqqRE0S6IE
OOFeAJNdCQD627oas51xRQ5WXW7EXQds8i10VVxER9fGDBHwxDs+lk1ybMwU
LD9l0hnZ5JHa5pRARIYeE8Xh6JuRRwY3leR9Li1j62XZ+Ebhfaf1E7A3Y7W7
o/8R9lL8rkROPZ4yNPogfOsdEF98JBccAHmj8Vg1KISSBs0No8oEAvRB9cvq
jWULsdCCuU9dIqszVyAWMVYyZ4DOVWj/c+sh7HGQlcRgmSOjgjBMDozSJFDe
jgMIBGI2Z6prE2SuhdqYDM45aqDIYO683YRM5kwfXCbLgh7erDJV59rDopqD
si+teysOz5BmvzRPLVkP78SDUJmTBZC+QDGa8c1TFLUZ1lMCJEB1CFnsZ9Al
xtsZ95nhqG9sgLjlDMdTChc9hd41Zfd+w/KSShd/U3Ob62whFC4nyo6b6aCV
4pMD8qw2FEHORHr6M1WFcUEhe47JSJUQv6Y9GUoFXbeFxXvLjVJqXZWFgPSq
oqoffVLKQ/7J2l7WXMmVaypGshCFtu/NxFSh1timAe+UXbO0ebqD47vwCVy2
ZYtsg2QPDaOANcuoyUfoFAEi+NqJbxS7O1rvr8lIU4RnC+w8hLigc5ytUB1c
3G4NgE2flUmvB7RT2d1im7r/9GsaAKmc3aOqlYkkisJmg+FbCVbqqB1kelqr
tP3d94DzAx1lyWkcbdpPW0YSUVFMD32bu3pK79qIRngJ5y6PC9Ir/9UJUG/Y
wt18Qx3nO+F88Yj8QQU4n4zR2nOwYkgAm4Wf6VGJVYPxgLdEzQgz5862rIjQ
OIkU62IlisrRgpzUJui6JWoa0zd6WGNSls/AFhB/uIyVQkFnHUfK3EgalOd9
rJXV3oFOiQUHwL6QDZA+GtfsXKiRKAA9jQwm8PFfc8ZMyI0bKPKOv133S2lo
0Gjvzq7s82KzS0YgLzm+gXVfyy9fokqgU/1qIxXTLCfXwSPm2HM/BeIOKScJ
31IHNnn0g+8n3ohV16+F7WGQLePObZLxThrSEctJCD1ForJ2+WghNxQ+KvgR
ZYwkGVuJxTtq3jiwe2PvPaQOOVpgUHw3+dQsNZTTW8n6Ru0cLb3e/eqoguEK
Fmrj5SL6u8URGEb5xPyMikFfPsASZH139yp19LYTo3d1a9wc9oObBv/Iflhv
CeKWG+S8eHfrtETxpOjErrkamv6k7G3zZCAHVA6d8E4mI8UlP5YsiggPHAPr
Xo2V8Hi6HpaBlGGxyyw9mqm36z4E6Ho8Eis562o+b8cNl9loxD+Vki+G9z7r
CsV61ZakFpy/O5VtE3hhMQ88dAMfSaONOi4WQjjSHPTSPhXbpcOQND9ppImw
djwQyUwpHWi5VZJwP+cQs2g2nGOjWo0lFaayF1JZ7u4vZbm7Alfz1Cc+QTvO
r+cVHRsziPGoW03T3mAkg5HMn+K4CiheyqxVRKzJeJj5DQwleV41U0oGE72I
9JW1SVEitT7WRYexs1lTjSmGYtV89TYlL0aSAkm88PJl8FJZO5AWRZIsF3cF
yRP+nDHISDQh/d3ojFl1R36ON8pPAFNeBGxnyzGco1sp4czdIfRMpfKLPe+N
ulJ7Nrm2jjmk/Hmwd4KPD5RBL5YZdySA/yYdkQUJ+vOgu/misr0E9fAsy4UW
nFtYmMQMztuffxpqcS1rEwRyVPESTVBMUJIjii7jeve2OnjUKv0ldV62yeOb
/zX3p1d4NzN3gl6p6khzKwDoyKboDMzGks4E4fFxQG/T3cWfXdeLRJihQPYA
ncqeVZqA8QgrUiasrptcdpTpgq+6F7aHzhAs7lpqlSZKgJ+nSxygn5gK7Zlt
W7fhFbthVHK306c9/AZgwq5rcxsuVTgBHlgIDuIzZlbDNrFQ1L3IJI3uvsEh
AxBh2IyRh/GmnhaOV2h7vZE8HdGNj5UDqhZfhSkuJf1xGFXQcqd76V7jkkv5
9OLtIGMK2EXPXR0Q0hVoSnf95otulbb9jbxRHqVGcoVyPDHtndrWuRmQWLx4
F0eLzWdfaHY1sf9gfLNaMzM2rh4zOAjN+2B0jZv8MiVRehPs1P3Tkk0YD9Jk
xmwlzNxSCLkQK7/f4JpIF3BHc2j2J7K36mMD4o0KClfgt8BgjxHgHMCUF5nE
cPx562z6vBanKToZzWQS16U9uNuGnhyrColZtd5qIw+tDsAMfXETiR+PsyB7
7T/CZtZsi9IXn7RfpAixMewV3oFbcKWPmIsgGUyWmkscRwPXo66nJ/UdjkgM
h8nnl8tWiIglap3VqYfCUGDokNee9osKSBMdGLIFtkA7QJdRYXpFYsH/W65g
3QRnZl+eub0Fao7asXBWpAAJjMgzbwTP/YQTbzJy8+0RPptewG+Hi0DgPvDJ
BZsDBkTP+KRNkO9s/N9f2FA9YoyIcz3HYjpMxhzb+YuciUK9fJN0INxGDoQx
bytInpXVtE3zspahKYKqcP9iQ3kHSmm6cKoWbG0WjOsOIBQEjAbB4hJv88/b
O15hOrvs5uUIwWcOWUxg5vniSqVcMDXa+kUfnHFqXhAeP2lNZfGAO/LakdqS
uuJCPIaX7yLKYWEByOgggZHZAhq/oB+asEREFWvifLH3KOhl/1Bsj8MOyjvc
kKOziyRJ07uDXu0ZawbJWL8gIjhySTfOpXOpKYxu2/2W1oAVgnyEnz+FlAJD
/iKqYANUDkpETKBoSMR2UxA+HUlHnx8GWxc9VEdGV/7Ltpxze6MXbRFDCT5G
KEkIn5h5GCZTCZot1EHBR0FlDpkOa7LV2DEzxgJtIMzdmyvxcEIsiCSc5LFa
XSzCyzwRLw2EXPK5izqR26DNnRJ7GlYL2tlcHanMsyjgfyd3sHUOXDM3HVvI
/BPZ+S+o9rzKVl4zsOZ8SnxJuoFJ0UbZRUWl07BdmAUsK1SzEr33d/VWP7Pa
WkdlUj21VnInlSdAcyS/hcUN8d21H7fmlPnVcOMWPiyCYZRjH26rUD0/kKMS
9GNCIZ+pd94LWAcKmIVqQBkDZoBcGdoKfFpMWyXVFk35KxsfNFVE9kXfJn5a
c8Cfbmiw69MNy0rN5VnRbHhOXVQHKfUlgXB+i3p6N56D3LVxDmUzY7iLf52C
VOF2TvnVX1m7xbzAVrxNheEqod6CGSZTIv+ljxOdCujKNJ6Fid3nx5M8txaE
3dBjzJhgNUddRp+qNinj2k5yf779F6NAqAQ1dky9uleE3UevlU+EVZnhL6/8
utUbKylFRldULi2HxgzDDcZ3UVantZ+WSlGOQMh29Tn4xSfMThYaKFR6jhOx
yJ9dXPe0YCqZahLYWhVuSn/qT4Cwcu8igK4m1O/BIEATzzn7E5HXkxQLprIt
VfIuuTFHW1CbDQrEwuqQyzmw8O1zc4VdMS0t9Pl80cmCO/ymfBm0ufkjdJHn
2vMyYZK26o4JAX7dAAVv8NIYowL6iIF5gcHnfliAnTQ+dGjk3xqlBex37kVJ
XDKAe/49MISoMwixwK55ZHnvnbsZMRSVvIOs7zu74JsPqxfIrwH3hA/yTljY
+p5E/MzJo9ZdZ1tvxS/tmJnj0CNflpW3eDgy0xohskZvCuPJc3bimfZFQaCj
iEAwsL6dvkNw6m4UuVqsvcR3IHX+v2KO+7gCN2eDtWF++4zk3P2EbAEyCRji
4UCUd/glpDpKsnnWs7GEJjAGMicIynFJSkAdDLvIVy3mRQicYAxp8rf7f34W
Dw4up4HFnoUeoQarW+BVzUkFl21mZ3x62CEPOMIdbO6m1erwQ4IE9hFqcanv
Hc9TYfQLW2kfCGjwqC7xJcIBuahXsPc60/XK7mSjUIdy338tua8+vEFirxXp
xyOQLdNOQ5AH+nnso36OoAMRD+P9UbsJrW/q5Su3n1liCNtDF5jSl7IxD2YW
Ot432bhjwZfUdGVjiWFLWNwCKVtfXfCVD15UdAzjx5Rr71KIauZMPxH9c1c4
5KtyHspYrs4UPhEquH+nJxaCc09Qsmrj71GXYINyjKi3cWefwuMKGCfaacrz
242iebx97EXYjURTDbPO8MIIvbi0iiz0n6DosHVgiKWZMc7dmtL9WLRi+7mz
3LY1uSYSxOpSXL9shc3H2ggELcO2XAR9uAkAgGQhXLP2JTFyWShuh047pYsN
ACKQg9fQmVPuI+6+u8U0Vc/qGmXumRRX++bgvKWBPVtes10rJZm6aopJUK2s
i1/n1BN7cNsNDr3wvfwz4rvE6QF1psVvZPG/n9nOU21C7Vg6lP8bx7m2XuPn
5USLEln2Rwt+chEvW0D0sypW1+4PitRsXbUvR1zxMo3RhL290j8dJlGxahU9
z49FnHZEl44ZlzjxVGWoWcj0FOimfrY6e4Q0Q84ahDEVLidmxcEWjaXJ/JiX
hKVaGVm2TqYGzxOXBtDoGPXceO3yZMgkBmIS5EQu7U9YpKcwFrcG+ntevfa9
Y+5ZX9zpCXrDLgvYGA2xgs8N+wvm5aQKUPivbpYzCfPbIU16VWcDrvohB6+D
mphn+ukVxq6XYv14epCDsjkuQk1uJJqzlD8HL1et1foaxYKmcs+MLV9e3ALw
zucvMMbOEpnVDdy9jbJEWDjmWxe1uwSzF6w8eLGQNYk+9/4E0qC6WvKrXrB2
WQFHhESPPBevz9VX1h9vOKVLut+w5gwicb7QSz3dUjpPWKzQ47OkPj6oNuBW
Y6AycIyEx2LucXjLutUhlOyKmkR1X3hYFeze53t/faaD9/Y4jwgB5eYGPJ7f
UmdTEtKuB2kmLt1aSD26rfsqO9TjCad4nlxAwqebZQA7/n4RA/mbvjDjo2VL
Qd2zEpo9uMbBHBY1yK5dnwx5nOy8yo7DQLbrwFzIg+cR6LGVz7NwX1+IHSZv
0UPszbxHpXKu9icz0/TiyruA1K4bvE+E7cVy6ZtCNK+7JRJUiud5aB27fKGE
ju3b4jSUjBg/ZfCFRvB09VXIWMrps+ItPSDFaA4opplH7dChs05q2ssoMyA2
lx620Fxo/r0joDSoV9mXRx35lcaQNlU9oF9tKfiBn/8YSlspOsgjzhKAOLWX
i2UIR4ptcyP7tJa3znRaYnfQ384bAZR9jY/yrXFn4n732v1X32TxWjkdHvmw
9RpUTU2pv/vPB4OrITJhKeKjs7qEETIYhGo9/3LkwPemJthJjvdHmPPjQf5g
rn30mOfwtjF19HRJwertzmuTsG0uooxXRCe25jc5zhWSMD2f8jJvOAsw/yey
fwDhcS330oCcPbCkvfEtIMeLD744yXzdcCdvRxgk0p/AeZ7DASlllh3Lr9uO
K7ezQySQ8zgSEHE03qUFb51Uxu9g4GdYxTkh8z8toxe3WJcaugk/MMHmHdqr
uDNUF0ox1rCpCpQ/GopDc08JefxYMRoraTYu9EKPB+PCyUeObWcSJpuylBnt
vjrG22OUJ9TQD5W5jmXrhimgrFAS31Gcj6fW1pLiHwro9VvCq2j815MniRFs
m4bof7xbyXPOzgisfnNlV8UmfWqFhiG9HSoJjz7AAdMFjtxmY6o3kccoE69E
ZppmxFolZbASRCFQvLEKI16QU1tCrKCZsv2foBsCnSCjlcpubNX97j+iUHKs
SVZ7fRyqHxrSjaLDQ4uf3cx0cYmef/wEmDRa86Rx+bX0FbMmByZhopZrqkbE
bL9EQJ4O4fOLh6f0FUQl3w1EvRQT6HkiK0GJIk9mrwOMJs6YbkLvUl4yhp6q
PrGn3Ep4eKuEZMbQCStX7VSQWVBqXHrM0OrBoVpQZFdwyQQCJr1J9DaIpH+c
32Sl0IMmRig3p36ntB1lZVMGofpTk2Dw7PykWcIbcm2lelrR1Gk8JRROL8om
hNrCLxy8rEOQmLC5vx5Zm+gSPniDwVe2aUiBYviq6OPPjyJJ19KM2/Wu2Ncn
0f6kXuCBQoGIyxHMcctdqqj2Thtbl67bmnC1AOp9NfV6LI96K0VcZy7dk5TJ
mxKIM0q0ckoba1XADHWgD0Mn4BX8sImZHVihPMi2opct+UFWBdUtsI9rxopq
Szl41Q3lIyTZpO5AFNc2dgfbFQ7lzMIUQGLBEYa5CiCYTcYBIDMr+ztN+Noc
LqgNnjoVvCK64EM8iZa24sBTxj9t3fkLyj6KNBQh9HOiJmhZn5VUYz/QC14e
MzpReirKkxK4owANu4ksB/PLFiLHETLugHZBpfedVPd13ZmBYlRRprxbgCA8
+4dgdTNrNcmU+dhti9j8ZDGivlf+L6qEr0JnhuDjXv7vWe1+w4B0fPtKLYi2
IB2A6b0vkvfL8g0yqD480IuxoHphku4IPo2xjQUsj+oda0wfkQTiHHkv9VVR
Cc75fBUcfpaEPqsT4FHGColDoFBSO6Ld+VBAFBHZkxwiMViIdSh26NrqhO4p
lZj/4/FuulgJGM31CMmxwuMwc/sn48GrY/E3eMfNKvsANFX6fReWP8KpMrHK
kCBq3YhixQa5QccnzjVk1LzjtFcnLtVowxEnYoCVOYaF+Z+PLFE2hPvkQH9X
c8EJVVCbGETDWWxevwEqKGtaGKqszETdU1ERUOkC2tluimyJncFFWRfmfCy0
Y4lUFmTnS78EEVMvLnlpIoBlQc6Dhrw0uOqwlM0+yOj+U+MX8Jt9qjgEDj50
/BheSmtq0X1iFir90V3LeCwIfHqLhC56YkLrp5njRKP73eZJZ+vtVhtPiq+j
fpq2WR2asIdmkZQyRPSTb8jIyWfbrVCA0JsxspVG7d61HLDYuMmLrphyZMxM
JMWqvq1nbuXNmjxm4GRuPnlHGFe2lr6JU/NlIC8hcnDVZPJu3zJOPGim0gKD
1x/cbSidFRRL0zQxZL/ges5tNhW+HRhrreLvLNxNnLfhWssl411kSyyZsYco
oE4/FpNN4aXxZiHuo121xGav0GoisQHqIllI/PC+BnV7Sx8yp7cHXcbiArGb
T/1/L5jpwndIVl5GfBx8FmdzS3fALTBC29MtOkJPiS1KePdtqh02yS8s15cn
0v62UqxJmXFozQz3P3sFEp/5bV8rkQu+YEYPPlf/bueum466LSq4PNA3g2As
eDZDjp0TkTzhnkqcObdIniGRZNCS1aOxRx8HkgKGgBdNwxTl0bYmtbjwLeq6
t1/HvmIWTCVoiv9kN6fLDuirStf9/iAriJW7fWBlY6hAtQgE01ZXX/SxAyKT
l+xfqSmXhzxuVXoGm42s0uy30c7zI1BM2pME1iZrSX5NyOo69wrqzlpqE5wu
iL7xVBPQER+W2vBGAaReM72Hz4+m5A89786yTk2w1E+Op4kl+1o+bfBIOVkm
O1vfkYGD71i1/EbP8j8D1f1Kp0XAxUTCoOWlMLNjA+k+lcOgpluZazO5e+Gz
DLQMkmzrZTtylq43nr96ajeN7HV/rbBXT/VlLmKNolo2WS6h4ZSJbBnUJwNH
8uAJK/F2bUqrBcsYjkGFGvUy2hAwegr5ntK55EMF4RADvjIXJtKzCY0D4cdF
X5aLiffjSjWhQLoSKPKFexFvETXShV0fyPGw2MXnLIZ/aS2AB4LORl1hs8B6
KlsXZKrvTzinolbSO1X7kSnOPO0PYys3NmzyND7cQYbPfagyaoOWfRmvTmTt
aUqOl3bv+wsxhsc6U/5R+25DgyEPwWcCwa9ejklG6xvqIHtAHI0RKwWVMgY0
lG4f2ImQjVMW0EhhZAa/M69UoG8st8HNPgFUCVeQIhTOuYWnhkQhEk2Tanlt
0x6b05pmjK9raw/DZTSXLt3okaXBKzAVcA8kSaFjBL700LPvDejGCj0I0Dar
fMyXemh5g+whKdQxnoJwoMGVT8wnAxW85MQAaZaH8LeK+20l3X1RMzrCxpjx
s9GzxCn+FCwri0NlKwfs74i/ywKwHDYcI7og5ntuDrT0wBPF+sZPy/h16KVL
9PmxJVbPCg3ICcO48fM1Iozf8Mey0c8amZSxHYS/HPWOJmnNrog56BhwezPo
PmBa923M2s+iWCDf8GsHI6ZO4n4VrbhmVasV3HeOzBgnmY09fe7KFpagsiby
3I2rvDjVr/QWLXCUwk0j/zSImsrfvGF80TilukXe5/U9bGN1RsQHK4ffdMEz
0Wuqyfq2MKChTYQXEWZObNIKqlyEtAIx8wT0iAlYVkgK126nnGltAiU2DXOI
761XsZtXz4zCPC1n2m3COJUvicvaviXXnte0YxkqsmwTdfO50J2AVFTaZH2o
sS6DOWnDB5cJZaLR3lIcuRQvTBSXoNlTxYRSfkekjnfylMHyTKS8MEorZ4tT
b077fnbuBrDI249of2i/lNTQusxSfT58QN3qaV+WqLL6L4TbkxHBRjJ7MEdf
nAoO/dHTur/kbBPs5jSeNvL/GLipev01kA7e5VqQHV9+xBzxfO7qOkorffnI
qYu8xkFWCzJqpq0VzgFRTkwHtVjwl0GtUyrgzATq9hwEfWdsquNxU/2UgB56
oDD0k6wzEEtGcPUvdUpEvaZbHjfKoDedLG1hdqfUgCxxp+AgrwXHUfmu1/8z
qL5qZYFIbP52c0Z+4hWyoRKGavW7OZDAHhaaOWkSznt9KkABkdCB6qND/Zkq
kGyMqrNgT51M6FFbgmkF+VZ/67rpmKgj9Rp1x8DQd/37dNhXkJvGu2vv2Bnn
3DkWd2ME2RQ+2B+43lukdW25BC/JhaUnv+dyMedh1qrFSBIWwQwJ1mv0sKAm
e5S7m8tVwnS4eMApckPlXsnr/mUxkKk/SrDZgPiJyf6KXIdSqwSBdwH9xce5
50LGa/83mMAWCvQpENI/0YTk8i7QkwXdDnfZ1FI1Ca7EsS27o98in9dJyZyh
0DAfxhKodticEECjaKxvgPpK/gQ2HlGrJtrso/KW9D5Ji6b3sLEPi0bySCob
D5tYXWs9fvkAy2Bo4txH6/JCVXubRJGr8zi5kfQbsZOQDpUsvwdsEhf2pn6Y
dXo5C7okZgoY46qepTYz2KPiYogk45gY3wieLbDB5tuJlJFzSUAnRalLE1Lx
Sy0W6vOAbiLOXpLdmYeuUd+w+bfw07jY0X7197UPlqf/smP5NK8he4Tf6iJQ
e62aaX31wG/70llM4G9zJRxTD7EAID5Qm3ZPwsqU1/+6xpYqFfj+/iCv69iz
ix+kZQWF4GHKNx6DhJig4zl2Ghqv873x9jyUelB0TNxC5pEfHjXZVfhfmKTG
o8GQA2ewlOIuIsOCETqDRPPW0hb2o+ED987HqlxAPwHxAqjvfXcJOcw82keu
tderR2fiohsErGsm+v8Az2mXFToqCPmExSijf746eNwnGT4PCguPEEVIxC8x
g3xuKxWJnbjKCU+eJE1g5fnJCHLFj6RORP9aIOXcIHg20/7Pydfc2ScG2KVV
6Ha8pZVavsTcl1jczwDZ1bpUPIvqO5V+QdBfFuStpelsZH5PubjdYYojNq4j
wVr1f6NRsH5K9RKhHmmNvb0Rkf4JlVihZV/KzMX6ccP/7J3hGMkaL2fsyd8Q
19mn9z7xGQeypjqTcfaCUBtLFI6JEfbEsaYrCVvw/8Tk+ufRWzVKf7FusCsj
okWKZrw7MdZkidg3XlHjE75zs/j7rN7C9ZDEUDcIof+Gurqv7PU9ZIXHsUqi
CmLG941q4DF/SAcHZD+imjVijBTpf1qKIZ5PNs4ncW80kiRFbvhsOwJk0iGm
PPfZB+zljk35PzrqBy8Yao3asV9ziEgvTRPQw9cyYpfQXYQFoiVP9Hc/EOBf
QwH/oheCRaBOi/fHXEVa86tJcO5ZOjGcRBon4xgj85wI1eTH0PSfYyCQz5Rh
Hx266yew++CNpDIRBJe4FcrVMOm3/b2gcUDaOmHC567xsbbZq66NkkRH21o7
tcTw9LMtoTJ8BLKjkZ6ywNxqBDofvcEATQGWuUadTtAJMt8FFbGUzWBetyzj
6Ov056Hz8o3uNFbvh3eCe13frM9wQuDjVW4XnMAsv+sEh3tT2H1CLvy+dgwe
7agmmf7nItfeluz158rSlRnv3WBRRCprb/8a4sPH5RrDlpgnAFuj34L6OM5+
gb3NBq1+qDWSjlaucaUjQMsxgZbTr4ckYY2rfdIzkeJioFlUITR4B6MQTnfA
2wKGiG7SUBgh8WDjrG9gDinL1ZwoALC89A9ISKCUedTAGUW0gF7VBj9WK4RF
i3yujUTxUFpryp0sqVFF+8MPXIIiU/W2QqAKo59wiAShVElwFx3guhvM7pDP
VFGkvWoxqoOhBQwFITw73cheGeFBvvR4YI9KqLvWXNrAqRZcXkuVPSSGcGgX
PfmjyezXG8BI+BKMvUPPuJE64h6zniGe4bxDO01Rxvkm8GL28F5DpFjfKMT0
YGJPCpSS3MG36EvjnIy9QqPDKxZytFxuJhYWa2VcosleGfL0ep/XNbfoElON
oAq/qpHGv6dOAEzdi/pLrdkUEYUdPNkn7bJCdbOF3gkzKCcFkKg85ukWOcTS
ATdWDOoivp4CWNw/t7vWyKf4o069rWiB8PvC3FdtaQyd6QBddT5Skfl9OrT8
huZVrMAG/uBd7SlcweBtWbA/VK+6OIyHjxeSuLf/k4QJgv4rKmfBxafxUc/M
sFy+sV+n49p3ARsIH7qezE2Ho/C+sW3QJmcJdV0MitIZ06IkwA5x/Xd2i608
fQF8pdMaLBc9EGDEeyufmdE7e+TkL7n5+6UlCo55WF/NfuUyBKHPnFU6+V3D
SAOzTDz1vJzA3Sx6aRvqWaJDspQf4o7jyoqQisDuZjcMS2Y3uiZVp9YDY0Hj
OyLC1Rcg0NOcC7Btv+F2eD4b5mzyE5eHlT8ElGBkpSZexkwoVHrt2lK03OBE
tv8l0emOq7phrlu0ee0+Mlq82jbrirX5dcy0Ya562J9mcPkcBaLAkFZGL7gK
+D03tB9q35Gf32B1nJ+qLPwFjHGDIr7iwuRj74F0Dm7gnNoknjMwQ3Vx1qf1
/GQGK2PGIVxh3oj0MCNRVAJWw1IFbD/LY20uixLwAuwhCi19Fr39JxbIxdgM
O4F11FCTe1jsJnCMUuEyIHEv8LTz3uiGTl3gme7o6ugXMGFEALjJrRWLRhhd
9ReKViDjFmLz+chh97zDHjjRlldR1XSOwXtLdnSFKtdA+UTp+ZB1iRzoOiGf
h6NapYsl9ca1pu/JTTNZA0p2tz05YoJuhzTW0n+zFl99n+XHlMYN48IeOCSv
hu9bLaoC9xim/YbV+fWI1dKbW/u3l86UXyUqiTryb6YwNiept0GzUJ+B625l
vD7CuY9lUZDUZmwUZuTEm0QtiVa+JtmDX/PwZ0H7q+SG5QYOeua/DgA2C5ON
b3Ibc9XuJQNxYP+JCeKSbkYu6L8a+mfAiV0Y6hhplW+ENZe4K+kE17sk4fdY
ChyyerqDQQGWDdModlyVwXjVzb+3wU9ouX6T8Ht24pGWqz5RGdMLTSxhyBgo
1RwMXHr5t2F4KFcfhVxRg0lR8XKGj424HI/7kNd+tBcX6ZxFTyNH4eEKpe+2
oyHMOJ7vHmtKFS1JoDZmNZ2LMuHqBs7NSyXGSpv0wouEM4KZLCeJgN/u1MZ6
ZuHQB6b1ZMVY/JaQivnGJBJ3QaaWQlh3n14mWodaPQPccHkSS61fA6ZCMdS+
77v0aGPLjb8a8sPOEKEZgruUqU1AX6R6KVTlfXkUX9HRM2IkQg+F9kuunpui
juHhmVZoOx9wAjLAAsPsHGZ9nW1YzVgvzXI3Q2auEo9gInrN+eIy0wggLh7Y
g4N2VzNpsufN7RTCq2FYIigpAXw6Hd2wi6WNmw97bqpJBoTD5WE1/k6Pe5YY
MiembT5EPjyAQlaceXZSohdBzUjF75NGxrsJDZEAhvQ8/W/JKyuqU2BRo+62
+kDiTgcgj92zmaLLMC+YWOCwrlCLu5QJRj0R1PKUP2PJnIIcqjkU5om/dnl8
swj4Zbwz62bbSjJ/10M6xgebPfGRimoGz4vnISKXGztT2dM98tB9WGOcUiUh
8PciYIiYehwxjabVlpcVlV7vb9ZTk6XRPhmFZCiAj7+ODa8wTtzkwoAPyCLl
mbCGAgg60btGEQjIbP4sxmd/xffeZd4sYO+BB5PD7wM2MSlyLPAEMTsEjReF
3Awltkq/q6+4EzXuwOWYyhjbMo0Tv0H+8ikubIo1eQqEOlb2tcAjAtxpzHYO
yFL9Z2p/QB4yOG8f7eC29JhKxw/W1o2/4mqPnmyYS8K3SYKahBngHAQ2m0De
j/Qf5FVIqRb1zMPUUzqRnMDgmv+QOkKcAXza4fFEWd5LI4za9inBHHZhkY3E
vt2J5M+1ojxGj9wgzvA7DeercdzbNBiKnB1pvJYpmiM6WdiEPTErzMkbM7Z6
jjquikX2Jt+QNpu2XONqXKpzKGWVSdHI01aYO45JspE0QC3yElRqCXoQ2sll
bsJcRpv/dTMuuSTyEj4ZSK9/36KBoNt7Gjf9xXrFCtZ5gWY2XuwAja3pImkH
Tx1HO9A1SxlZ8vja6oHHmP+7BqErpJIRQbOFsNsOl4boKfS11VC2vdhigY3C
uRaq9uJ9RYdVf4mMX64ThRucU1OoRCTEyfDH9O5BBtNQAN4eSC+yJnQTGk0B
TFw68yLLYTMS0R/0T5EHLcn8Je3Y8hXbBOPX5kmQkZNPebz6PEPultiPBr4A
bXz3C3vAhUVV4a0pBzF6kWQ4gTvRq0jUFuCkNpNCYhS3BAWebt7MUI/17diA
sgue8ZbJ8mvSOFLCHoUOu3Hs6+zjYvIa2/83SY6V5cOuPMAyD7pcFLuAaCr6
qheu8ws2wHboIEyMRi7simMOKxIbIl7Qd++RB60C0+OplI2ZdjGcuGmp6nur
hc2INdpQ/4L0psDfjYcRU+mmIKsODaq9Y3+jkm/n4njRmVX9XjXI9jYrZNfj
dfm/z3CYN0Mp1bUdk8JWNAJWFkvkWBFnUY1WAD2kFgWEAu4gzfxZbD94MqDM
DxPHzh3dv5cGRnK3vpi8QOThRUtgpIey13CA+bEXuU3bvKezHiFo/awWnRJP
gYM5EVnM4pGXHyVc0u2GElARWKFS8pftNqNSjgtvKR4fiWboaMrIaDzIG0q7
gkvdizpSFHaPIpDb6xON6eF5iJdNqE2diSua6C4xeYbwOlxzn1LCAx2dyN6X
gU6/pVBcNVUgswoMouVbpSN1xerF6eXwU3niyb8CGuZSLt0T6zxQKIUpGTRw
jPA+HL5PhsQX/XS8jeoe/lBTaZhiH/lYkBg5JgEM2Ldv7IzX0nTIV7LDnO1Z
uOHFtz94blZD3xp4dmGcC+bqgniBuF2mf2nMorI0q3KZfmsAvlEEzlcYihzd
1WnXwWxuzkKfYE6OfQKdSN1I2/Gb3p0SM0KtS+DjIIM8DdZhCxVE/Q5EJ7nq
mXcs71BzFC5OjD0RdHg0jNM7UXNgW8/Dm9Ph6iymyxjeERiT1epMkCbicGy7
efe7XZ+qEff1VmxFiUFhY/xneWvprZISg+GsuSQXXMWxAMecFqOHlM36BAhC
JB1pFzJEugOMtD5dmBugDvEjGjQSSwjGLTyXuNrBup70HbVkTi98qKXSyY3v
7ufo2cjP1RH6OANZ+rcdMcuszrEd2ERPMCPeIrFIzBWYPwiiOS8WsF6CZBgr
VYSbsDyy7HuoESnTTR2mG39rizjZbOdL+1+c2lzU1lQrHOSVCiVL9sA+ro0o
0gbie57/0TGz/XqPlat851Te2mA1sS14heb17RVZLM23slOvdEyRZ5MWgzMw
kVa3muU3is7VY4wmH+x5xVgaVTM+nv6cHi35sQPV5AM7Ajys/ekudQZ+bqpf
7vl5brhE4EFLX0ij0SjTpjRW+JFHVUmjEElN/Rr/ZhWYb+iNthKjuBuusTys
3+LC45Sw8YZqWhDCwklpcTfkJ1OwXxLhkYeMEbnNOxRgBcUxui8wA+wkJ53Z
WU4AoURLa4i3zVnCXgQR84D0pEvi4gmiP6SzICZNGGmmkTzhHppuBkJjejqD
x+J/inb0dbW768tBtPN8iLd0TKOGWFvVCDzWlQL0MKft8d4nAQWxfBGF2lM0
gcLcnVNf4iQm9Gap1v8bNUbh3VqANZYiOYYJWebW9LW8UcA9lyBmT98pJwXW
y4k0DqjaUGZNyzlUHbhH0tcrbab5Kp4+I0Fs9x5idwwFcA2aSyONuoIzX9X+
TULHqyiLZmq3wWNc7WrwILbHMGczLUtTBtWs0F/IV9rLwNv572OobIjKqmvf
6J6B15VJs0pwemsxd0yIUN5U08l1a8YoSx1IXfu9eZ5VhKUnBU2ol1Y0Gvfw
u5dAl67h5oPky3v5WXDUgTRjolRNv56cq7RY+cQvG8iWYI8uaCFrA9ya+2/F
LusNXJ2Zzns9Mji/+gTkSbHNsplaTN3NVHmuVE7nrzmhVTguTxUf9f65EpmZ
ysb+Qw8Ev5FXwBSZI7maSfYpabdETuJoYXGbyomxfJr6he3JrAG7LDT3hmiM
22nw9Hsd1yLxf2ae2RBFCW1Z7ZS+lSLZvdhPruU409OKziB76sl8XTgBKMKL
W+0EcKRYx2UhoYpI17SkZnd5whgSr0nFyNS+35qL4+c+T0cRjj+yhdjtMsLs
jf35nub11DeH6EL3YQ/1fEMI9rhMrpYFn51zSeaw8RwlUG2wm6z1Tid4uOOA
uYY19fi3lLwyliQC8CTOaQdiANK1/ohV5RXhKbs1TYfp7I7ZcbIX1LsHbtwA
LMoRMcY5iTwuVhoAfEj8fOUCBHvHfsGuUlLexlCL8FQQvdhAVxeiyouiN2+3
TzAtL+hPvKoFnY+kf0EQQdewJUw2A+SkYHXZ8bbiVayP7FLzhj6O8eXum5h9
Bf01Pap+lNV2IfbG+UHKaQ/Sgj0lihw94QUOr/WllO0IWAFXctLUJ0YKj0Td
9H7FVCgvfBdtO6xxrVSOdWMzHuM+pwUcpLFUB+au0+Yr6Vo4U5U3IJpchUh3
3s2c2PXMnJyQFbWsUATcT+0RCCmUShFm9hHcTwSOlAiuZvptTC/Uuci8b/1N
lax0AtGQty4clepu9+/JwaQ0bI8wtkATEAcaaSsilTGLpt/rbUNmm1E4Fw1b
1jU43Ip9Tfzwn/yRwK8BmrtAMy6Q30dTRW9/Hi82CqjqSYQnAd+9U4zcgiVn
Y6RFi+/mvhq6b0FcxIjnWUIKqqnOSGF2h/P6wrsWQfFLa0q81rKFoG/nv1NY
37noFDnO7wXyJEvvlzRH4XecpMtZ2AByrja58HQavzlNR9icrCRdRCiAJb5z
fT2dX+9G1ZSc2rvhfc9Qeuv1Ds1fDIqTs66pQZFxcwKYmoSLjrs5PdGD+vyc
f1BH681KHuLN3IBqcpxb3+DOggwLvfQEubcszS4Qzp1YaQsuzKWe+qzM9xSq
XA6bRGeyY9dyf3McaUaKT2BU0Y1T9xBpGCfh73iQh4Ijx2gR3OFhPpX37pa7
74C01xID3a/zmmN7tab+5EwEEGbX0rbv7qNDxIIcGphWkXTeTpP2KD8jvpVd
iX9lNM6xVxWxJNjtoFPa9OEfqUIGSQNuQ4R+7DAh8/g//MX4E1r6It/awoZ+
/n7LyM2SjsuDkjitwUfPSjluo4QAPH+1X2dGh9fWk8Olz9iyyrxHNqOkPwlv
XZZTs9p99Wb05yfPMXH0rQN5wC+8ecY+1kpAizKDLheyIOrhH85qleMVVLpL
PqmKa5BLbIRsspN3y6MDv7pBE8EJ2rpIBEE9atptiWKXKEPEwpySlgND9FqK
2OldApHBCTjbdVEmLUGV72YYdz8VbEMIOoh4r+0HFaBiucFZvzN+61bOqLaB
yBbfga3928FTVlB51rHMQJkOIdV+WHOGANaeghCjyRBGMzCRnLN33JTsoc8C
yxF7TVG7Jpr8olkfDLlJyjhBkyUaRcrWp2PVMgBaqnlEv5zWmUeoGTUlrIPS
Cc4+54hxdHi5pfFkX7ul5hyOFudXMsdRU8mSyvka83+jDxdsQvDTmMidzBq2
0+CBIH5w48MTm/GR6HF5LcV7FcWuaySlLGVdgplWsBZX1cSsg20ahZ9pSLDh
Lt0Pz8hApv3gYUK4/Qa4K8wPBE3htW+FUR4KhZBzaGz3A/0bpyuLsS5bsdBO
Su1nQOfYPnh9YzMtWpVSiPs6qkFkvcS3lUqQ1M8e59Z2Ujg+C4/oXC5cUMt6
m3HyYLheYkDzu8Ot57165bKzzZQmmCh7KFcUa3KtxJGnurqyMgGxuxcm/Jb5
uO9pxLIRgcFQT0Wrg3UGhqBqvqb/DA+TmYewXGYyta7CiKNNlJjfCdcv/2aN
YD4CdeXUttX0VhwQtrvaPncgRiQ74zoZsnCCWkStffawPhbjXA7/ft8WQQgB
R97lb6d2/VoVFhgRYxRI8og1epA39i36l2WdKnNSaPY7XQsJVeLKzEJzjexY
8xxQhmPONI3pPGy1/PA5r6sG6i7OSlIct+smSGUHxoGuGrc7fCQEjYkFBaQK
5vUvg1Li+4Li8+6ZxCGmuI8ZzHOCZt0xm/+Y+yPht6bjIskVY7/8VPg8JTS8
Pk2+SfDbIAWNJovvfY6OMKVdrDmHYr55ciUkxhsy8XWztDekqRirasL6vD91
48hB71Fq6nNnclVzVA57pl/iY5jiKqooZbN/sqN95Ttw35UMjPYvaoLGcZ0W
qexR3zyZ8EEXk70LcEdkW76UowAHbm6+ZHHc2hThP4S0NnICvmIyAKShdxXw
ykqmYadwji+ZIfximam/YFRWL2cJfHDnmbcywTinsreJw4eQWeX4sxD6BcJk
dE3Kj7fMn/YgreVO57beOl5rJeskJniHgEGdGNonNcuh1ZzJOAP9Peed8/Xk
Vui51ZDgTMlyd80JozhcPDi1Qrc9JukKrc0aurIiWxTjuCguBaW+5fsczGub
BaoXmERRHas8D8aJcS+IIypf1bUF2CkWbp2WstdRxQUA8H1T4W+t2O/WrHIU
qIe6vPTjDZVdJMpL4n2+Su84ovBQGl8dLeY/KiYGBdAMZ6m1M2rLcdoX7m8e
SQa3McMJZVv0k6E5LW3LrTCmMtn6j8qwVjLcZJFlAm9Sb4BJUjKkws1pUy1M
oZAfCQwskhtG7KtYUNdc5Omz3joT5Mjnr0yXjm/KwdydUms0pXodDm5oyERr
ZbA3D8U40kDNIDw7lzTFt76kS7+05yLKKRaZnicWGF8qOLiG5/yRf/0RXr+F
0yEYwkEJ6FrCtR3IU8kHZE0HBd2pg2nkY+JT6zdQMAho8ejwJkjkAN9xfdIi
zTyxE7/y8YMmGvcfnBU9GKVyIW/SBSa0yTPzG1MEq60o7kifPzhvr6Xse9at
bZ8GhAfQrVOj0lLG+oqbnFL0OgNfwktkAr0PenyYmUBH0A5DbSgz26cYUckh
f6XrHNEEMCKRmEJQxDkLRHg3k8dhhaP+QZuaFTuX9zYGNzUbJpxoncDrGnpK
FBpX8d04/qLLStZhFBpZAtseY/8snyde2/ISWKvvK68HRGKoLCTxoFfPKOpg
AiEl7uPJSU0LXp9eLcRZEB5VK+oHPjTMTFdCC5ZzyztodfsFWD0EsjHua40d
IPbMDZDsX/usv6JPWvAoR/qIBlU+X1ZGCZkZGiVGWlgJwZScDg1fo76rtOYc
yfeLDitYCz9QRQkpbXaeV88VpPYUu5/Gs9WtM9QBRk5CZG3CBV27pIg0Jgyw
1yZfJrZKoWMaiYwD7991Cp8cXjprZRKlipGzz70bwI0Cqs0x4E/X9ztAO9Tw
3EO6X4gTVKeZKvQ3KzQ4VjPSoXXyYdojVBwd5sbDsTKF5AHXPsXxy3IBGB2B
RiTrjSb3kO3RQZCZ2YiiTdLSfz9mFK2/9KBrYuYA0mfwW3Qqhwz7Kems5yoB
5a9/f3vDg+Pr/7ElWpBgvTH4GCzd5GXawhHUUpk6mumHnCgglMlcICND/FCZ
m1EAN0jDKBRy/NpTaUYT9/V6apVVANw8hzVostk2oh5EA09rHJdo99paVKIo
o6CqOIHQV9DG4BzXUl6SgcMwta+nVz7B+YwoZKChjQbJf+NhdP4/89Zlumuf
HYpOzLq2Y0u1BhgjE25bN6Zy3He32Z33QXQC+oqRIPiQjZz66QTqmdnsSL/r
QHkDuqvKu/2GyV5GJ9JNT9hUkDO3djhszHUa7EyUuOx4XfJVXOKXP8NQ7Gdb
pqnYIUKu7n7r8wl3prkxK6ZKN2ww25NWENIYyuD5aYKFGCVzTDgDGu8yleZo
fcT6eVTZreg7PTd3PdzOv7zJxNQ6+eB2aRuchxzy4SRiH9D8/Q6DSfB4/6bq
DGH2ZCS6ZHxp7bS2l0O2Feg59endXLQDHgg4Es6O9UYckHU/4Sd+FehLVJ+2
D91pN/I4QshLPOlNhUnliI9EOaw9aZxamERmHwcEXdzcuADo4xueDJGik4jS
RAwoVXnxhqgUX4xhfPaH81XCwLrQhUzBd0SuxQa7j/PLqSR7QWn5UrwhD/sF
WbE6VqHqZEhPcO2laH2RaNqWiIKKfSkYNlhv6rgm6o9jwEMca8UUqcISG02j
5zayEoH0kgV6EPDPeZrS1Tz+gMEJNF+oaNUjzufMFaroMVGzV9FVFBcCZelQ
sBThQ2hsoNUV0GJe/IQkwquoZ7riu9a0dY71o+2FVyjAaq5rcrDw+cWl9/Ay
1zHZ7FOoy8V62JvpqElK/gQhsTZWIQrrtmYJl7xOjlj1IhcKfbW5V5qtxJYC
XtU1JoMFoVWPx865rAx4tpaW7Xo1bJ2tzcqvfzojOMD+6IwZErlNiInfJQad
rzKQSyhzFP34/oaYQf+EZBe3Pqq2r7eBj3btkyGlcxWUAFE7984By4KBhwxM
NVzLHbfgxP7CPJCkS7JEydjN5ZhyWBONFUqs2JV0CHm9qlfOoGDAWdhFcoED
KieEL6NMJKARfPrNOAofQjFGe88pscNrXrA7+F/sCAWNLWOaVwrtm8YnEQeI
txjGQkfQsWLoi3sU8Y0xYH+WPqmCj8HWbDazS12s5ZORUAfqPeKeRzTTOQyk
dhOFJ6SoEPkGJGYdz9f3Odaf6jUYvBwrUDrPxYRaLy49V56IMJbEMq4s1FzD
YX2fHW9lPdk6Ctul9dRCgy/fvNP9zMDBP+yK9t8vLj9hpJtQCCD7hb0Rlkmi
hpWrrwiLEkTJ1YIHGVSGqQo7cSlC50F56Zf0WgMyXmWWcH5JXCxc+f+y3Plr
pDCPmEYTa2rw9HCLaQ/zeoiz+ECH+QEoJNc0Q/spH5vPSJKAgh4oYVjeIokL
Q5eKMiO+lR4NFbhuY248B/UtilHrxZFogB51Oc/bN2DYAlN4ezbsHwVJAnOP
x25w1t5ZibBMkWWHWTvRTLVmYEW1IrHp07XzgLNnC24VS+YwvI7XlGubdJ+N
4/iou2avyUEbQlZDHZdR9x4StBJS5veMic45X5ItV4eXQHpfPkHzkkBmjjif
zvFPpuXZ4MSeQSURSFtau8fTHx5wBPargUWkjcP0J4Px53Ps8YXL2XuW8Al5
qbe6WmA44+mmn0jPxvTUjju9/1IAUItbaVzhafInOJ0aoQqqTZgXHgA/EIUY
zr0gnM57jhhgUPFKhGYfPnR0GTeQONkSV1ZfWKfqOShj2xrhCyAIW+EzorS3
ZjHQm4u5M317O30vxpZeBtZDFR8YBpM6hkN5S7FYMxSVy2/I2uuwnH0fPYfL
zG4WmW1IlpVxLmJklFfNj6phRMCuTT5Wl9NOcG28Arkh98rTfSPrAb15atMR
sptKid/T3ZktukGpFYmmkcug4xZreeo7PwNdaP00XEMzdBtMWOE7MA/79zAu
AIbZqWrlcK5roOoj6zY4LYwXODM/cBhDCglkye8vssnCDcl/bVzWdcQIv5o9
AjCJDiyaNsMhjf8WILSVPLB76nfcTkhKYfbLpfFQUK5NWoh4K1d9JO1LcnU8
DE/5k/UqbbYwdiJDlNK1870Cfv5f31QU3Gwj/CsRH2qOTNeRQrhUSK6+ucgZ
IJ3xQbg6v4CNBtTJ5ZIOVDh+HET0VWEm9YEYtrM0hpqfgGKUCz9F/G+GdQ5R
T97TEWjXqBIla83FXCotewPVnlrxZMsSp+ULlifsMSFqOKY4Q2LAznkRmTbB
6uNSRhMQAgsvQIxzF/FiQQS/Dj7IDtViTWjsjo37OiD+Ei4n1WEGONPnrnDs
A1LGsEr3u+yCLhK58iTS1ybOLnkONh1aT5mHYzQoBGXb8sVsvXm46B/FpSUi
gaV8HJcnY1rdbHJAoLFwn14E/034apI/dfhj0ohTSwMYj6mlJWJntHO26B1r
YTjc1Rb5iz4Qap75BxkWCdSDMLoxoJEvJPnLJL+es/2QeUZo/+A8vWmEmu89
k4tejGH0jAVuPFyyAZ9yO2X2DYSxHDXEX8Bbp6nBwWN65JLog8kuCEKKuL90
FEvBMEvCUv9vhnoLUdEI3k74l7wJ8oznXmzLihjWhjLeIrBikpYSBlSF101q
52o2EcRF6LFDiyzP2Affjf3cdpqeOuLQmQiQnohjho4+vWegA8rQo6F4/Hy0
Wl57vSiGDCjR0mZPxslpbwo42DJ/g+vPcfzqhiVbBO5RbaAcplOPmhZiOGbW
TOgWKJ0YljA3HOniT7wF+blJnpL2VM/lg+2Vzv6hMAvEFb5hb8vtrU5P+glv
nMhhxZZVjg1hI+1S5BBvo4d0/ivmJZ5+4m8uGuY4DmgLb7ahIdlOjqc4ek9w
jp/nz0/plri0uOq+y/gmjQRx7pVoG819E4Z96W2+14OpPu+XW1Y8jweAofkc
m7sm9Dauu/yBYVDbkobgeNg/gnNa7al0DNaipIBrdOURPlTDhKkki4lSAXMW
JVcWVyi7LLGPInvwpvBjEtbpsK1vgZdX3TCjzyUWWtv5LPPHJgsh+xfL+D7H
TYEXhvavlCp7tZLj3WJj0j6Rp2jrPeLrOQ6lNxCpO/QK6JyyICo3GUVUtTfr
lC2rWwYgaA4lDAy9LOQJuGKDKQFMz3uPl2GllhJwR230d//OtCbdjFX4VqIw
u/H3bXCXQQRu97j1pdDJ+Gzru3SaBKsk4uRwjjoAByk2n5mRb9dTn3Bag5Ed
a5T5R7pg7o/91lgiKC81icAOzumX1fjvAUQyNOJl3htpTOBcOdGf3v5e8e04
an2A+K4rimmyIz/wb/5l3Qwjo7XN8yA0yE8DAOZgBWZxcrZ0sXDZW6+hoM8w
aBNTNdl+KTAnbXzYC6qQPGplzNFutZr115ghoqNbJQHGA1HGtfX0S+Rm04Zv
2JSg84lIsySqfEC0ffTIK6rzO/NdCsBiqQ3hxrZCMG9O94buu0Xb8YVNWbFa
nnEND792KfnCuTrissSTE5/sUvNojuvhIwgqDfatof1e4vv/z6pysEYTJEXl
RV+58/mArGMAoCiYj8aeg+KY0W4GpRB+B2hO7SyqufYKZW+TFy1ueUmZN2d2
Fek7aWAGGOdc4AjGqkyDkE1KCD2xgg1qoLNZfeAuowWDL+7sryggiFTHRu7O
GCx8eUPNFbyulwHibbuJY3jeu99Mc2y/DH9BOG5riEJa76i2c7X6XA1L10kI
u8gK2UdAcvCS8zckZQt5EpfMdZ7kLoEYeTGmcT1jzAt6haDop0Qfqj4Hf2pT
8bnFSP2H7yjhW+Si5zF0H8tqDPBjBO6RN5Fh6Mg8yVQUp+FtpDXZ/bhqyCcq
Cr0rzB4GlLQgZKO0J9B08SpXqNaKd9FLO+O2D9zPHC8jpKiRxHKibvADb8ug
HiHqRM8WcmFsqTxy13Qjr/l7Htu4fBGw1ANsqTlyGkGxrY+cnFrd+tE0Rnqj
TGbM9Azs7qx0Nrcrz//IpgxNG67i73zvc5eHZTUQox7FFdmClAVUg4Z4MPQh
r7f+2Lav3V+T70O9VQQ0OskqQQjfswRPe9ZdXr9EDZKwQsA5t9HWXapDYpD9
HmP7JdYRGiALIasC+yesquWJdDtx0TRoAi1u4nXEra91cLAB86DZ7WRss973
ypv3LQDhVaqbhtLHe71+wiUzfbt3/brxMURaLzPx/lwM6qRQpSRIDgTTZikd
k8pmFVXVG49u/ge03NR3lVPHa7CKVJIH9ZcD9/34i+qX/Ojjk9GGuSmunhiL
fGM3UC1aJgXlc7Qq/fCxLyqAlPZNOjW8MpMKaDHyFsE2C5hNLKq180abPCX1
7gHJ5XG4OSDvWzsoRGl0oFbIxz90n3XgsRgFrpckQekxcEpISrs2YIIS/HtH
gr/ynbWrKLobDogv2RmWD14zlwgFGnnij+c5r/bbMpVwDil3f+294WXFLAka
n5jKyVtn7OuROAyoLBZlSymwqpMoI60vNNNaHqn6X30VRxXblL0ymdJ8c529
NlWCQkz57l/4vP9deAvmuf8LTvN2d1X5IPyE3DD5DmLzXNJ5GbRaUmq0e+av
B1QPKi/sKZ2Cd6yLVuNews+nDlkDU3/2nes4Dy+cDk67NKGvlM16w5AZlFFu
djTIc5/EsmmG4KvxqvsDrlD6jBmJQvT8OMVO1fHeo5KjtQNmf8AapiKMjZi4
HyfjOKF8z2zr6jYE2pAwKYiXq0I6XbiRyXK7VRyaHZoSUo/zr7B8UP5Ra2f3
LaqfI6kbN+/AIJBs5oKrHKObJgA208kwh1lv5Mmhjs//7uF9Xw+tb/Saqfek
wiJIhyMys+UcIeanpKh7TbORtkC3x+7dUAyxI23JVgakkJnEV9Yl9QWJDQGM
XVb4JAdmALiFC98/s7agfmcfe+kVUe9261yWNFojxx3pycbujEliVttRID5n
UapuG4K66+JwdH9LPn+r0Jd5ETC6qG6/3GyOYHnQ28bLWWZP5mrU3z83Zmt+
CtKFXPDKgQVPMeSIP3N29vhqApQuCXPAtpH4PV6jVbvQuOB98AWQA1bevLti
0fvicZ5L+0UlKJ+jpyon+kQw8K2D0MwceTO0Hf2m0rmmpdlQ/ZOr2VJ7BKJX
buHQVApwEQG4HltmCJ2+COZZdr+bkDAdVLpUJygAjFjkyAF0W8Mv248KOD03
WT1uVf+52t8TG9dvFXW/jUE1jcHcfGRAfwppjZzcmGD5eQaKqmqmsoiARnUj
4LIlRtleiGfalu6cErJdn45KNBlKUWfrNMPYY5cP38phqcua8SNwZiF2wfXg
76zKdUFUb+87EOnJw49IJATe1mgbGQZs81rOZGD/tjFiT4g87Wq/za6UlrRh
h0ZhjYclqIxwOAAIQjD0A20yPswPuvcNU1r9gUWZxbj4HzT1oIPfqSAGlmDE
RhuDYEr10l/DOQikz0f9dAHo/zNXTMCHSzj5DyamFQmY5Fl1OvS99Rga4Job
Fu2WKigJxmjuUTUwa9/anYJxVYxmlv5o72roaCSMAd5dSyYGqtzcf/EJd7VP
25c5rWoB5Tx8O/NqP//W2ZspRk7a/qfjOmVuD66Bf5yI4u4eGPhhqFc9LFE9
pqbCJVPFuY15F1N1Vdnre9olUmRV3IiXAsG6HbhP8bs4++VHQXMlrIRj5Sxi
GdtvrPL7RwCr+8gg4WlyePqxj7+WM+HJVJmbwzbabUqB12Xvt2l/2wOlh8st
oQPT6Y5YeyUiQzneknS4iU7BgiKz+EexTWPgvdkCkR/KA0sV48OuDr7DF/3v
DKbYzympkd6rp95WrHiLw8osJriYBIJC36KqpR3XDk9/lCvOYTt77+hus82p
BfkwQKQycdnp8trBJ9ehoDzAFKEPw7wwWDWykXSOVRJUGUam9eC0tXKBYgCN
r41ot3K2LJwMKQCxrTeweaOFDnFDJIIck4szCjPt4vvr+QnVOl5urmMNYsCX
KMEV8ZU+Iq4phW8FWT9gWP2qnxsygVeCPt0KNefLZ4hyrAqBkUs6DueV3hKG
idONDFq07Qh1b78nSpMCrA9Ve7jqEM/21xdX1e/l05dTHgYdXEgHM9z68wUn
AXlDFBXo/kdclPPuZdblDKETPty7bgg2WTMuZJdpGRO64ZMKvpLHdBk+lqGa
ranrYePwwpi8L/42aauynjKGBDaykNkZQrHrsZnvjg5JXY7Emu5tqoSJZvZ7
n1dAwkWGZTy+yQZ+lNNr87rnNp4UjE96TyOFUYqH9NpGdqAfsP3Vtkmb6+0g
VIieoUQ8Eqm1XSBmP3hjaEwMdNVXIwj1dmAKkAnDP+abiemxGxVAUe7mpZSY
mILEDE6YAUGd6EoOU18k7Zt16U1/cAcoT1FjZ3Axe8kGedSbqV30A6X60FF1
FqtjQUHiOT8Pt2oGi9vcgpkBGGbCFE4eiZYP1g+rDXh2988sEy+EJE2o00ow
VE9gIh9ht33YBCh+9TOVv/jwCGfMkBvPnAZMOzAuNeJdIzlTWTkjYl0o+55f
lSEfZP+aVLc/3eP+VYeUOLJ2A8fJ5HOOlIIuwiwUtvSui+A7oMJpTxReE1a3
3APgit3EOMSUS+1P9GM+BEWCKF2dVmzHbcETXHCNf+dNiEtu1VKPH5Jw3JyP
BtgnzVWUdOvzUQnYxMUovJf5uNRmyFrvl6JqTArXHUdID6VIuVUsiR0tVu++
HgvR7ZYZZXVXnOzhNejNy26C5weCCbFT6Y3l7cKac8y5tqIeuUwdVxvAtuAN
8nqkBGoRGE6PKH/4HCBEUUe1SFcRADe1jrgLXw/hnj5lG37NbrvoDSQzm+zY
B40tEK9T1vrsrSXyo6njQVYApFnRt6rYwHzJ+e4eMNUntOqjayxS1ZA3oA5w
XBo8L+aJYpWMKpSIq28zLtNrPIjR40VoPwUEuZ3Xac6pEeJIql9pUQhIkwh0
tej9JPludIX0H+okhMKFJLfbQJVm8/0K3DWSAkJF78KJWPCGFR2EPGTYo1hA
h4n10Y8ceWeQibbCgwpoLxd/ooVfvkyZNTrToz7GvO/iUVZRg45PxYDQM1mz
zy5WjPIkDnWvzD4v7VhUwAh7VbM74MMWqUhoPWWhpxc9jdZe+PR4Rw6yjl9m
vyZklImQxqku4kUuxNtLqcOU1WpbLSBnO5BnZeK3vHfMVoTM1jhoMyLC4MWQ
iTPJN31Wr362VmPOyh5Jmv1z1ov7Cuqve4KB8SWqIYOk+i4ufpBNff3W6p9m
MlWJhmgrp5ffFj8OG0E+0uXZu0zweSwSVXnnnNatV5ZLKYZUD2SywS8ggEjZ
IPWMPBQuLf3WgQAXM6CDav+q3B22hTsNXY9gC4vCHCR5UyEl05jg0dFUkyme
ilJYWd+9yVfLgd59bISH5RkFXv/rbO0D2FroWrdVTPEk1uq6J4kPpGA5UfBq
dQV3+rpl3kpZHE5kDMxQsnI9eVdbp2Rb7jAjEjKlt3l3pg3ysGgwz45lKBlW
G0C+iQ3iXj0A80Y16tVmOWi6iRsrKy8ofxk5yLkx7yFT73Ec5rMBUqgjziTh
L+E+c4BmYVBqsNruEJIv4Z62UC96aJgQ0gA2AlqM0qowNBcOi4x3qBEUYxph
B8JHqzJRBoPRo0McHqR7IYmUUass1MN99bKYkBZU2TX8joDqeePGJJVS2dJT
dHKcwMnEKQ7zE56q5FRrYc2qSs4Z270WDtXigieHCH3i9prteEzLPq4Cfm4y
2+0lqSuLL2ci0BiqYNTvLZkGCQ8gMP+e/uofClI4CtbBt2+HOHpsQjSlTyx5
Q3FZM42W52jLYUw6cr0R0EJAkVCqIE6XuCQ6cdcy0jun6x1PKfrK7lZK1Tf6
79GLhK0n9lY/+lDL0sMXAwclQ6drQhBwzlt5HKP/ZQBqQTkYiaOMNVngXy4T
tm13z0aP+8e0AR5RkfGp1o2LPtIEMtJEKd9G+EL2yyaOT9mMedy5zx/ud0M1
Ni7x1+NY8wPFxsUNe/6ZmNjzucSJFrBrNAL7mrYL//lSsSsRDf8xT3keL7mE
GcwOUPah7pQPMJzNafB02jKRwmFSBuHRq9GEJ1EMsXBBPbc2onz4cFDSsmhF
XEWp1zKwNepPf+T0WdF2LY7Gb3xwp7pzndoIBxnLoZ6CFJEZz3T+8HPp+xmq
WuUIHnPyedAnkx1q05EWbpvLZd+6saNYgVg99dP1qmxFdwdVTRB/OJA/nntz
ST2MaAm+ELJotwV7E0N89tyOSpZXPVBSSBj4FiQ+fr9VVBFxte94ONkbWjZ5
f/s3RA/9IUgpfu5QxAZVOMhkbDgLv0eOPkulRaeCLg4o39YejfLtqV5C9Y75
QFtwRyCdnJBm65QROdoM9o0iJ7xgknk5ugieBGoNOnda4ivvB55YX1OXodAt
4ClgtTrnviSl5qHr3xwMko8s4XBE2GW4B4taOYgXv8Gbm3+E1M67VSE9EQdB
qaASHJcl6j5LsRQVAfXVTosqDcL7QKzX05arW+L5FNlTM1afWilThhHeW2T8
4yhJbEBvN9MxqLcc9BAYMSXCPRC24rzJr+hrnjrySqRedYezhcu8CeDm3sfi
DmufTRsvZIV83k+IOGPTOBcFU1ui60pTMyq7pQDYawRVfORHNMicthau6PaF
z6baEOunTSuF1rOrD3+p7FSWW0TqBtWa1BErTA44kiFVnxUrAKxrqAONG8Ol
mPHaHF85I5gr6FR/c8YEfjNrgBqXdROqSm7PfJByMmxqlqP1QK4s56KJcXQ8
ZqanaimLbAMoxqkuDTFAtIr99qeXHJ2yZKhcmpgmcLKeYPwKU/rrP4ZoQSY2
2Zvr4rSTVpDniSPvcxtEBW9MHOCtRczjH3/W26kbRGE0aauNyThOl7M2D5KJ
QB5gwMMOJ1ouXrXjecCP6sOq5to2tPcu7eGQ0Ry0TAZPjHYEpiFyWa2ncQha
J3i+p0Qdw63usT4BF1WsYqEkjysHvFx8kezlpy1GVvG44INnjjXcfO7s/Ah0
oztzRBLkNM6jwdmoXtKk+FcFW6yz62M9QevIeeCFdhOIhG080vJdotUV5hsX
5Aecvbqyf81S7Qk4ZIklBiU9f2I9ROFUSh9yXT7hZv6iJT0eTykodp3hn5W6
oZueRcwv6Pe2vRQ6OXr9qRAyTNKdDIvvPFeX9IS62xdYWMmdosXYJBOXFGa5
pAJLECZpc9yuGIOc++oGoSJa6c4qxn0BVIBXFMlXlSqOLZWOpAITv0L6idn3
f2xfUxlo/JkDkYL7Faz4yXsbgu4qo1/TaLpj9I+LEor/hxqM+CCem9fXbtHS
q0OlXSJaf/5hLrUwOxJODaklvWlHHR7C7amrqo/dUA5mCrV9gCmu1yFMZIn+
wwTZiV0q0ISGqSguySj5Pj0Gaxyt7VRm4ptWG8SnTX1EqcyknfBQJD36RyPJ
klmVgA7RO0NmBRhABEXJg1555fuTmtLjKMayOjh1LP51ukMHZHdqQ570H/71
bOSBTOR5eet6JtPq8tfeld+CJAhc2IlTPmIa/bYdtL+m2x6j20XuEBfOMg/q
Xa/K5850UTCu5slw2FKnCG5JGk9BELiZ64eyEX4Hzh4QcekQ9XTCWN0xu07b
M+y3YVf9tMJ2K9v8WWWGE6qS+JfkFQvlW7kXlRpPh+TcijffOkc0YcQhsd1u
+uze3pCaIHxFjw4CPwHYml6ox9i+fo4cTuX5FdlA9npxRebYok8mVOq7ieXJ
wgTa4CDu1u4Pt/ou9qOC1BtvWqTuxkC4uAGL/jPNri7paZmrpA6aUI384+nO
/tzslSlOl0bZuaKMXlK94xx+ButSYxxfUeiobcXqe/bHXKiNwJUGtJ56zQGE
0WSks+ulPDAMb+PV1Gtrm1CT2njJZQRYLqgnKdtciSUS5PlmRxsNrBqFT8CR
6fIxez0FuM7kk7W78GSR0cumb0BsNJbzJUquharnbRw9fKqq4BdzJ/EeJ9j7
D+gvvy/U+700gpddNrDow92JHjEDC2LT7e+KxLV1n8bIh1WxlkbKvIBxATsJ
UoV6T3CrDvTPMD3NDv1oO0cZ8RqrdsL6HFARi3nr3RfikzdCX9lIpTiSdmtF
BtSRjW59VDVsy1aZUpMfY9hZDqR90Tpu75B8at4JWgq9mTZBBrhE7vzRZ3AV
jodYpAyOYRIyAxkykvxECtLgl//lDJwNqAo5XGMnJAgDD7vp/gdKuOo6S8U8
L3NpkoXAW/vfACXLgE2DvLBAVdPvZQpaYd3j2lKmWKhnCct5TNohXAr1nmgZ
NCI7UjvGeh0f3QtdKa0zw+0tlwnytzYd6YV+yUvTap8nUGEn+30nnySEkns5
T3jwmIBXU9Y0F9l9U98mOiZIQS7wuRK8F3Lk1qVYyMVmThANUpJXQn+Py2Ge
1beo7Zj/TYoAEn/7Hp2irAZEuUO9Pk65iffohApPdx3N2k0Hx1x9FbrhQoq0
cG0qYgZ5iORJUa00WaSGPKxdxG6hOsSundRW8kEe+6UntjT1raRUyCiRo8eE
aJX28MSR3CMyWMf/qheq0XIVy8eq847bTdEuvPUhzmAN90+4+J+WmwuR7NOS
xpaUPl8cV2NGwMJ+UklCE34kj+i+4FpbKs/dwHCnCOtTPO2MK1u0PnN88X0n
xnqI7gFt1IntlOj2MyXGmY2THtxoaZLF60yGuIPNGZa59F03DSGaiiR8lUSI
/W6IDhNAhHHy23qYvdbt+6iFeNMmo06rH9zEQePrLcmIxrNw71b+jsTPA69g
xu+0fgPZ0RauB19BK/mNdPy2Uzsg4W1u2Is3DnuawNsSFzDhcaXw310k6wfj
h549ECWQgst5jmcEFm3OEnn5iWsyWP4ukCSMTa3zZveoWF/0sS/jWvaaeEer
MOOBbiF5DACPjveTHqCKYJYMStEF1To63mSwIpJR9dE+kXlCREToIs+PZGM5
WgMxes0rL2Y15f1gDviOl60yJ2D30DxoWAJvltFxX9Wp5Z2ES+HetpDEgvuA
TjhWnVtmrk7B+z/sYnDVmCr91aJv6WGBMP2XiUJUkBuhSPF/oEIk1IvGMygJ
m+RUkXA9juEA0C+eHd5nyuikPCVNrLHk0SO4Pc3vbt/pc6UbkI5U+t3ZbgWI
bZ215XJGHUZYp8BW2rnDXd9dHym+51sj/cY4QEMem8+eLLl22bRvn7PMXFNs
aIzBrqVlWXWeVhPlhBQZDM8S2Gjr7a3lckdjk/oS3kZdiBvKoOJwukrExpav
Akw5+MFSLegqTKtU2FnvP5KhFckLMVmrLa30S8WtkG3DnUeJTBKMr08cnlUv
VtKq8Hup2cXPDEShb35AZhyZaKo5ItjvNNe1eb7SadqPTSqkV2hXoNmFhfQs
tYcpADozjZ05T1ERXmvnc7NU9CwaNqFQrq2ULrKUcoz2erOnQ3MB2tDEOvkc
n1UK4ne2jI+hzFt/Gi9EaiTgH2166WeErYCf7MIuXWh8iixFqTIQNAY/WW0I
fbAcEUTBgpy8OMA+4tdXLgJQSw6TFfXcedm39SI9Atlr5ZHQryySFuQhs/5m
/36tfGBtBacV0tJZXVEgvYQ9hZUdwDvlVre0St1oBgTcG0e/d0DO0IDfTRRe
eX5XWBm0lGVwgqOjKlUTXMeMSXRlCGsUy3V3U2cVuQn9qW+PKlruV0WzmOym
1E3mYHPifv0lcvsxXpHcx3Acce3UYpmxA/2/GUIIPcloBwyyhnMMDMAExwbs
gLyiFLSGBlBQTmCxYSqH5Ct3jRzWTkTXwuRgGeYVy1E567ZEMqUfTVKoUP5r
n0QN0XB7U5ZucsPc/ajBfiL39q45TOmAIhXn00VSqQFYG3c+NFQfCiPwF1TF
54K2iJ4vBS984fvOFNYsIbKS9xbOz1LyQ919c+k5He8wohRdsCJvTcBaDVfp
FXW5PoZRuuro6OrGCBgWzMAsi79qgL6Vo7+riMcbLR86L00iqcxBefRjuN5S
oxDCIYhLre57BnJ1ne/i6zeXgK2/SycklXwBIegsmnAyyMG2/KKC/haXbew2
YHWpjYLvrkWqMBmlkpWJnbFOvLNWskFWHde7fL9E5cEFhA9w0Twdk0tOZ5AT
yEQVaNj0EECCfS6lfqa0a1kqiOiE9/tyUfutZxu2q68vgArCg6RRArAwTaYA
PS9szqWyQBL6MHIMii5J0SFJIsBG+u6QGRawJ52n7Az7l2Wg1pM3goRtDcaQ
HcKm0Pl11O4iS8btf/XDzTdgugvFzOMH0ci+diWWBK1CSjAiL6IWJ3UUqwiN
X9+SJuHbsLVUHpgBHsgxKY7xbK+ugm4MC+bnHd4ui8LL1k5EmbARVFJYlccf
ejoTzq9OS9hozZlF8nEGgBPxRL8SkNjyFrx8/Rt21UDe3uvMt+shYfs3W/co
Qkh38aRZyk82b4oqScAOAolmIuq68V9G8kSFVHaYks8+Yas1BG2V0XG91vdU
SkkfVkLAUxSUOaF/MyhW8GKdS7Ud0zHS0iJ21SbM/FhwXGFOMybtQZwUw0kI
YMGL/iZKmJ+E3niMsqW2d2to22LO572+9LGF2aSD2LaXgDyiaJ9HnRNDc9Pz
d5HjowXP7uum4c/4WgDtYyBVC6i590K6Tb4PaQVkCf/yMrFxaWCZ+Wz53bdK
I0aPqtTzPEBv8Eb9G1/1kz/cHSGjAKCIxRaTWaI4frxM53v6bSEYcEeTfJ+D
zPQdpsIzNXGA8DHZPUldyTmMJhuJxYzx9jMdifZ62oGTYaqQlTO52IzxKHgw
mOBh870LpCBUqC7fkmgLnFiJWhrZSw/LeGEg2O7z03ofp2HEn0vnGWb/vwqY
PrzQOR30Zimi3jSvpFxh4CcGkcHTVyYO0RMZIGpV+Vf5806q2ypbGNX0j+fU
oaFl+FI7OKQmfUXggSVGTo0YhmMX47pJv3zuBw6KGphC6Ud5qLItn4PfxUyS
N6xhUmDkORauIdgFMtKhVUD3jrbEyK0WEXk1oq84L4Ff7au7C6wVs0fQCPJB
JlX0iAXmPpzb66ujVXqLWwmVCtQ4RLClxs6CVA9rRAL5MOXDw0P6J5ySEfMA
et+hApQZur5qJXbY16LCJig8bajwni5YybEY5fGqFu7ZvICf3suBM6JGlSGv
fD62im+uuGrv/TYtqVfTxGUjgUa+rZ2lshnTOVehJPcHuueFYCa8UP1qjZQf
sv2uUfd6anRBp4+syZ/I0Q68tB/T9NHkrYsv53QGL1/JxzQA8VS6Coc75FVf
DJpdoIxUniig6IpzCUgy5Degrq7V4m1NTYnrv/K2g4w+Wwt1Q4dsxG0zlHsf
a5kQjhg973dGyclbeDgCEvITaaBgEtTBUIf+/aFKhm1CknVR3X3xc0k2wTq5
mwpOi6zcMYADsztjJ8u/OQLL/PzOrovpAJf3j9HdIUBRSY5l+PXbKZDd1XqQ
AXJadMjN9ftyo/9Wd4hjY9MugR6yDl+O5NV6PlJ6i0w1M7SVzRo4S/RtRDGO
zb/AuAyRUJTNdNnlE59iRuBuXOKdJ2tDsCPJnn2k19KfKhjZ/5k7Ps/4PS5s
fk6qdqooSJS1t3s0pFS91WrVFw0etWrnZIGOQfEIaMwOTV667TfR4aY6fFn1
ZyqecIgRcBXLE/15PvgAc6tq6Q1+YaHFggsXlj7qnZedLoxBIthrD1xPNww2
rKia7wD0ck/P6EAvjBCvgSN1GlfjKDrwoNF+3D6guKNRPBrf3d8VStzD6SZU
LNnTqBfyVCM3bXlyccqjGdPD4N7TFgAh+9b/slXc6SO5ogEt2dP4iXAZf50q
fXcsst0tnH72PwP9mSQFM+vdiBfy3BuV2yUyYjZbkrz5j0SIxViSRWH3Y0JU
tgdouQ08Wanz3v2uaMFC+LI6HvgbSuJ++EqlIXBAumJMpIS7TozBAF9UQqyz
KzXpge7YUJ848CH2NxTp9usj3+LUXyWDQybKt5I4z8sn0dZ5BkPCnM0vyDcK
o1dTqwTYzV6/hMVdiiQWh1R3ypSod5eYuFq5RXuA+K7yk4ezL6m5qLm1btCv
3bIL0QUQrce5eWPov3wtF2qfRWm4d3l2v6PAB6tzxY1/ZX2tpMwGh76UzuGK
j9ijyzrj7oy3GB1YSARCyTEAsBiL2vmZoIVnH0JneQzPzbQ1CCu6z3+D7J4j
M3G8QUyYfkwXrkEhd+osIqwtKeRAsJSNJBHft2jo7XJeRhtRyro+QhSY2pB7
NXHkG5MecRpuiiH2lXnEvlALtVGysZyZR3YjeOwnNMsgu69/XQfnUGnDVOyn
2ywLg0yDBxmv/W4nLO0oHI3htGwrzhOsZIUaCQR5z7TJWSbexjVdDsixH/xW
lEdxxa7SSt3WeisB//pMNDvfMPElbP8p/wWAuD9yCnNF4UZ2SmCIgIl2A8k/
rWHCo7w/fkFd3yc+xwJnhc2bfAVDsaPBGItlIlpuRMR9iB9i8fgj+iZI8d8v
SRpvv02QxyEHBva2vFh2PA8vwI+7TmZCh6JCm4/vt1xbIpIHJzOdrIwVQJRV
fFvTQjRkck44y0pzxnPHFNOqAoJczg2nKyYzxzCikkpaZAal6GiiMEJTbBfs
OINkXys8cvCsTHjuBTA0678nAxVpt6pMZ/00xOI6SuUi3sUkq9Isn/uPByKm
d2BbZGhmK0SHOkBhaiEld11zIOe9x1Kl80nUi7EVIvC7gomQ2qjaGfFZHwLX
SxAyDvTvz92sqbwOhGWB0YF8zryg/or6/7PV7IQMREm7OswBhuyrwIUxRzaU
Hajj2zMvutaM5fNfFn/G7PyZVqU7OB9j3I28DtHd2lT9zuOfqPPhOMmnr2KB
5RdIRodQHoitRwsp+a2PmiIJdoxG/hBB7fDiMGFRAHbPwYRzwDyyBprHXEzS
ZAUrIJAAiYZB7wEcD1YPb+4yiGJz0Esli0n2kVYdKT0jQFoe4v9uuNa0RWDE
NjA2Z9fn8WtAWrpx2oOLIR7tP+22P+7nyBvrLhX3fG6EbqtO/LbbmWpzJKiC
oHiEwJTkTa1ef6y4ikv/13pAP/PyOmqo5IVP/eUkoRVY60TuYm65rT9HQI2F
VtS7HbkpdLjsIzen2Si+4qDAVAeANxVpIOYFPcGA9wSH4+IZtj3GYJBm0xcn
WjYzR44pnBiag2GTIGppppsWWsm+axQdpFNTUBarSTgJRYu/WIWZfmk+TP+s
hYA5lKh3/azArhNyTfg63ZtyJpAsFezPOQEX4DzeLkxRgwgTKve8nhS6Q+oA
xhLQhmw4pndzzgklqKqczO33kBL76XY+bU7IgXM/G38HUmHh1uORfWjNq41r
0UUhErAzQ+aNyTphzRucypUPCa7c2c5yb9ZIWk48+8wnAv5JpAbjTxvvpRbq
TVOlbRLo/neUKDhVpwIwcBVN3tJKw4SEIx81PVH/fGv4Ebq+BPZKDZACymmT
LC2Eslt1dbmncXFe/RkEM1zr8wmB4KbnqfOI2mpDoW4K7zm7TkQvevuc5aNu
LpZzN0H3W6vi8Sn+cDK2blCUrDOqmE9zFNCrcHJ4C3wSOBHOzVghSYnhAA1U
AqoOdu9b+vuCZFxGKvM/KIhn0WiMGIWsy1vkj3LfwkkOXWuWXOsh6TDtqI2W
ParRwPyNq81+7vBX2QLZ2ihgTOnDKMSm8hXF/Wckk8v+TwPEz6GZu1KVOu9J
qgmD6BDmrc5JmlAEnvZH14/Y/Wz0NaWmm1SP4suRZ9oOjrIx/SuyCF1YubGi
HuFH/B8vFYKfw5yzdJcmone3WdXiht6YgGgRwQgxpWwG+EO/9LrgszBIYHI5
igaIWCa0jKS+eO7YGuPRoLBIzzSA9PAJ6/MXXRWSct3yUejGe6qOWtdnP7je
vN2ZBilBHRIjsrtZqJ7lRWMECTSweBIc8BAv1NYZh4Ql5HKHMj/9nTHXst9F
N3V10ScxNKXnfHU3kE/o+saDcCYi12xfoYz/KrEP3v2WwZ10dCY1F9g+RAYx
whp6bIVEd1qb/yG/RO148ube8w18OSzoBipG9e8eTpx3zE62QJ/qrdwSGEh2
8K9PKUqMPCC/32b7DF1bbXdGiPkWkN/FRnGHjYj3qvbI2GQxhf2RKiBY6si/
qE2IbmNOQht1BvK+XsWZStv4ii6pUtWMeBiDvP2JNwRm7yKmgbzSRVR1lB3T
bu5cHim7bkidrDOT2l4/oyAh5zArVJ/6bRiMS/AwzbiXEsGMI6EfrkaGyYWY
T1hISjQ9Ih5nqoo2NWoKj57L1dFfLwbfSAAxUTB3/h2zJMcBLpwnDQgj1rtd
FIlB6js6rmWyFOF+hp6cpJTAmxIyJbTxtDFacoCOEX5lJRlOpGPBPSqlan+z
iJJZjFONh3GqlgEOF5Tycfvc33JMVplsrZkEnJ32gkRuDh+s77Gg8S79Rmd4
OIgM6e+sFc+Rqh0Z/rFouN/kKBRrx0X/gGsmbWyUX65kgbW3D7EUxmlFoaXp
TVIx3dw/XYt6avcnrJFL3W1IFpngjXL8QezGEeugb7ThR/s6BwZA+ZspQjBY
r/urBdjkA5wvKlTn+zYM7OYxOagDTAo28cwF1i97oEZdNbnOHUZc1iJYESy9
F2UIxUfOd2dUTHmEUOcE+M8VkX3/yjqQdj22qaegd/Edagum4gvvri4+wKVp
5k0cIrR84WXXWLFuh7LwgcVL3axisHK5WMD7H/DHiP7rKHY21CnEZb16/ll7
aV5Ln2kU5a3SHsO9O36/WvJoWXsXJshm6+xBco2GV947tsfXTKtdqUhdcehe
5BnEeR0jMUjEy4XHIDXohP8z4F9lnkxoOa4BxEj3Zke8Dme7+65r2CM3P2Id
YCk7mwD0D8juJB3C+E1lE6Pj+DfMkMtAc4ZWcOHieCFlqCWePG7H3Krs23vV
C+RroGjHo5TwCN2avbYpKuPBlT/WAUu1sh5hcLC2qRWysnGY6AtiEYvytLCf
Jxs9s8qp7/R8i/GyLWJ2rdRokTpJZ1d7dvCKyrUFjVI5zhKVlrd9HA31VgWX
M39tQanev7BZFDCS03QHVURsq6vTgCaQyZorO7mQkuX4glx6lU3/ZRuE0FKV
83zXX7kMhS2KBndlxj4AkH+3sCt+MbrNNLCHQQeQeZIEEidZZbcu02TwkMkz
PG/YCIjCPkx2qzUTRRG0dCndrj670yyKzdDG4stCZdbutbu44iIqFbaXE87l
W6o5tBlE7GufLbnF+VoLABZe6rBlGQH36LkRH2j0AMb6DIwfpnt1eoQO+0oS
bFJASWyYCcTjgoTBW5zgOMfQpqJ5+yLmSiXus7dXGLei+bbqqk9lZOz31JUE
bni3I4Dbat1pQKiHxboBqH8JPTsHdXfCcqFzOx+U0e7YUYkZnfyChN/SCOpa
woxUAURoixn/0JRoS9StXvTGrlwF9/AzTxyRD2ymkZTYYrx4CjrASRR4RxKm
57qpOxVwfo+Frb9Lvv7u5t782w8JM6slqUUuaeNNlblqoMm5cBwOd9pAShNb
RMhibCmAU+uvhU3/8UTUCa6lOpH8voYV7DT1AZ+qNFW0PDAFOW/SssW55wJs
8RZ0sEmV4M4qtYbUM8AS3IwXcHI6UbZ+OC1LjynkFfXEbZ35KPFYshJo1D1d
JKEDup4NiYbcQjap56EyGZK1LpiFwT17+eU4+/YGy9wKR77mJbX6d4cMye2O
fUHHYof+x6/4OBeOMhZMzM4ZxwLTpAvYrNDRM5VrEAIrLh6Wo5OtDBtzhvYt
feUZ/LIxJabU5aYRhCxTB0eOEukerQn2Pf7ytfbDDPVmh7LjKisftJloCfGd
LMAj8W4uaPvG3BrrrKFd9Yolc08W5CdhZontNmh1826g4b5+obZUY1uROM81
GhvInUmXc7BdavQ5ZY53C6r4Wfc1KJd+U6i2AfU5BzdSv0JZV9ttc2pDaspX
UDfYUSq2iAiMY+fSrVU51Ae8BBFGoxw44LIJ+htRqbziVK5zXD7AUxtYtGtv
ChMmTo/XV3tCeEqgzxE1Wyq9VzeEoShWsLXQkFXukbvPboZjPYBJ9YnLz4CO
GoJYaVDugSehcEF2RCeAojriJFznbiP0PFf08Lo9sm60bodk+IdMvpHFtzCp
ohNLJQw4jLUdvY8C8jAx9HaEEcpE1juRDztgEGWROCSzeXmOqOndt5BQS+wt
82g75Beekk9i+QYcORJ1FVd89PCeFsW4Xe9yRsSimQQgYwwJKeZfOJBvDZe2
mIogB93lXSlW/Y9cE/VaqUYLAgOIAu4gWVTRtQhTMUF5M4dOUIocK5gFTsco
x/P9ZPAvHOZW/XXsaSVKmM/7TJEgBZFQRfY4HocgnkfG3slV/8le9qJs1H4j
RnzO7/v5hhWzOYnBTgYUOzgEU6h+INqLkk2jnULMyuS6KzqQvLq8sz8lxPi0
EOmA7npaJjPAQP4PTDLW+pSGQIpd55+9a4IUhfuVKVItpfZx1kznsfoe/fIK
5GpxJVdWZZLKfoaU1ET+ESQwW3oDVCl3HCRFqDe8HlgbZdICLdW3sqIZageO
DTqRhFRlzk96Ght0rkZcAnzrfi+rFbOTiaC5wb8xJxpFyN1e4mW+iVs0c5G5
dgTDxTHtth1Hcz1y3kuDgiNrg+76p8OgEAu/QztO1cdx90fjK2bFhuQux4Xh
+DafTQuLB5Wb0WsMkXJcIKyHDw5tjq9wvxkdpZJEFPGkr+Wnvz2GSuH4xzQe
uvQcBjU3zrMcX/D9qmhJWwS8Iy07MS4zEYtWD+W1kEJ9Ck85lf9U9Tqgg7QU
cxTcgjUM74r7RSi47Cih4ILo7fASVOoOKhNfm9QbUvl4Jj0GuKuH4pSfrqBY
qnAGRUKXJ5ImYCBvi7K4n50LUjBQXP4tlKxStSQhHJ1g9ZFxrk41VYZHDZy3
gvqAOSnneaqHWIFIyiM3x29Xa+iDA3flrGEt4nbnLmW5PsfH7Kjnew6MF+W2
1p4B7D+II6s9ZwShu3kCCP84IhKd3UWSl05+ncxD10IXSbLrWiaUaAuPGMbQ
rGSRDSd/OjbA99ok4GXWl1375LnPgtcJN3pdbFGKyNJGBSVkbphtlYLPbkdX
v5kzzrUT8FwjV4qOaQNKUOKU9+lh7N+xf1StZhHUBOSC4bEG7lqTDcVu6Fg4
sLozdERK3FKTc/TwH1PoRKPXOUD7hj8tAVH3TCbUvP+rW61zLMSa4lRffG2y
pwCb/nCiOaGZE3ZsHImubXiAFv76Bm0XFnbImjXQQyIaoYezNCk516JCu7zU
3VJqTPrH11beUZ663e1r0ZhMA1G3IlpoFStWschTHdJal9xfflG3r2OIHsN0
8krZwa7WLZh0H21+uDzqYcQ83c6eU0WqTC8v8KX6uDn1TRXKwVBcz69b5fI+
3ZIWm+vbpmMoo9hStMhzoeigDDtIJQwDY9jW99cQc6mHU4v2EeEbsXgss5us
EZVmblkcO3rHlmoPC7EbUFWvttQ5D5BrdnSOKt5Knb/6RzZDL+7ZiHYuv1GB
AE/AoupKXtdtk3dAj6Mt8F11aTXdc7MSRkoNakxOcPHsEl3PDk2MSoZ0b4S4
0cYWDFwC0JGzyWp3WuCIHGpYNtH5hPyWTh6L2EjDRiR/kOFtSeoyGEUACzIa
m/Ohra7/Nh1lBqtNfXYMLdbeaY8yONndmglFm1CqOreQ8330fswnTnKGn0O+
9ruRgTUCdTkhknKX0gvEHVwa4IOYDCr9Fg5MvG74/E6s6/m3pacfjhQQmR9b
dlnswo7X2PjXyUi/Hunui63Nz2d/XrUzZ3vF/mO4RhuSRII5wtZne2vuMYxT
/sV0S8r6hOX85ICvRex9ahKpphN73oEiXMASZFq9et96JMiEAMP5OUFRI7Fs
NiP2OgoWZz446kBqCN2OILYmOaYW9vM01nPT/g7uED7x9GRPKu8KBtScKqBV
sKRwRgCzsqfV/R/TKXOSP/DhDmJMMySl41EY443D8OjfC/jL9LYvfBK8drO9
rwCQdtMlpHj25jmwnQsMGqLIFcf0VJRd4VpwMgkF2jmCNVKLWOBI2BydHubf
a108R4hJut7bcQyoOk65jpzoGJiu0ZPhB8OYAdzWUhL+CRSfXUIcjh+uJenk
y9wz8O7zSaH7IH5p9cr5TxLaDoQtFamQdw6LPadr0n8+SfMLniPaa3dGjrYl
c2x/i3hUVE/q7Wh/ccdOR7CIPXk3Uwt2ZVVK7q+z0LwbDzSSPiFdWXiNb6ly
1dyUzSsxKJKOL7r7jB+5C3nqdDVl6Nw/70QSmEHK/4aFlpg/e23kbIXRiIrG
M5j1ie8k1vrzRaUssC2nzir25gEOF9K7cG3Qr6D6lo9J/xDEUp93wYygyBPa
dua8k9tIq7oszt7ESrrq8wbRj0P87gyb+wvFjLCH+kntxuERLD9EPxEFPKcg
Gv7W8j2ib71QSUEiA32//KToOCABab7iT6AnCRjOQkUZHILHNH+CVrJwiQKz
UMA50tBLI3tPJzFOojIvKwr/8BeuZmy5tXl3jUJ8+nDJw6CzOtO9SW8bacYC
sK0n/2ao6FjRlaOKVtLBOWnLSNAouy+NthMutuIJ8LMb2io76Zwz2C9aGVVD
IzaD/i85Wl1WSiHDUE3EH8oizBLAVEtSHztGR1GZgOCkQydB9Q+9+H2H3ixO
bfx1KZp4PwuZXWucgXTcJ6+cy1GxLIfiMNN4brFt3jU3451j/BNZIUcuPJte
1qmTAjY35d0nSf4et3AzU2iXSHaLZMiqIYbeblneitFn3j+c8w/UAuF3KS09
hLg8DIaoBl5W3iSICV8BIuqcgflMi2b4PL+cs162B8wBP3LUSt1KLNwBHJVz
PhWm8Z9QhBiPN3WkcYXGqy/LA30u032WJc/PLCxLOpbO8P0CHMDuMGYfBqYU
vrYDwD9gWCCGuVVtK3mx53VLWrLNb6+8bdXV7rkUhvmsE2Vfm2UssHcxGKc8
noJki+GXErp7QdSSLNAp0MMdmAJXUMcGYA4GWlQpYHMQn4eF4zXM+x8fby+L
5IDtMqblpPkyVIBUDYTLkHSv2FdF/+bG9FI1owtc+pAphoIORpjttzjLeLd1
C9tLnWwM125sEcqiPsWAAxJw/sCHkXmr1qskLSPXO/JchdpCvAERviMUdRpz
dNf2dYDd1788/9nC4Ii3ODzqH/xPiM8GDvYCMTgpLbJlN+SbUMtA9WID4Hrs
P/VbLfNVPFg5lwNp2X9e2xDXUk+zRZGWb+7GEdAwy0onsfS+a4yd7Ro1fkdr
JFYVhUACVv59sSc7pnOtiTfrxJeEdajrQ1vVQzD3VZvPQIc2QtQ8RPgH/32j
KrZWXhwMoT0aVzLvhkXOBUAdv405W87WPdij86t99hcyndSmeWgK0wK9NN7h
xjct8fUf+0noNdXbK7ngo4YATqZiPTV12hKIIqPS9L230qlqWegV+eA8+8CI
lJ9NfoNDVRWLlMOPdgM4VMUZvA3+KAxoryZ9R4u5lYwzW11xewUr4t6cKrCc
18b/HTPNju4DYbXBafiDNFGQsLzoRBEYoY/F45x6MNNmLamm460ohOvdM9pf
/5i2KYxV0sHVoFS3xgR3G8D6NUmu0N8Apr1YR7I3sX8kQljLyaBxAQZDJ6n6
/oXjsEtPBjLryYnOMcZvJzPrYopW1oAQ7xQ6QAg2gpkl4xqmzZNr6XIA5vZC
IvsC2rTY2xIDMQmg45+dexbEyP8YO1tEaJjr4iKDl1MeRGCiJOJ4yqnWIbOi
q12difgsz4uPBociZ6Tux/qcUxnTgdsp20XjlcrGl83wdqX5mW/YmyorR+2O
RmveWzloroM+SCPecNHf5rFSdACQ8S6RTCPJkOOfjAImN8HuK2NIbQio5sf/
desXFmqurPD4RzZIAVqzSdGBw81WaFAO2bQFzDCUCwVAhn354X222Ojo1wEx
Q9yrnWcQtjD+TM+jo3V+YbJ1jJ1I7nM8lv5RRprjA4oXHli66saC5Mlh9uV6
78yPHEeivswp9Y9X3X/NDasyXlDusMY/KIowuwVvTy17YdaYaSpgjBWl68xZ
o6DcKmnhamXMEsd16oszunvjNOgRFD8bjAmx/elAzrCbups4BjQC2ixhsC1I
KrkuqSRGZtqBWY1Iw9ZUZ19i6MNdtScqvT6Z/WEMtw84rvqD/NgOn4yz7BuZ
+j5sBZNrh3BTbkK18kX5p19cCKrptuGTRu6IcnqYGZRYTixy/5qXs54llSsr
NSQw71zMpq2U6uflZJUuZmnNHChAJGGzEE/3ABHV/QXbuKNA9p2zIQuUCy+0
GZYAPUTOBex8R+dK25aMMquoWzQRfGwlGSdBtRvovIwPEjDaoK0idaCwADVb
bJdAfhg9324Mpr/Y9X+/eXfzEDKOhwP4nNZ+94znzGws1oSn22NKias1fFaH
1i7hPhydODlYMvT3U5dlq/Cow4IqDUqlHMV+0MCms1fxNqUhJHEpfm8sLsXY
UwCkehWJ1LxGR+uXL2b/y0gIg9r1hTYOLR6jF6MWYb4jLikITQAnrZcQ8pD1
qMPc0d+YvP3JJyplNqSCuXxo+Ga7YuhtNYWCj+DZmkDhFqlITTTLSFqD+gwp
hJ3X/30o8klvMhMVFFwt/dwfQWdHcUzfEcJ5geCseqT70aMw1CMYbX+F2ydT
A4fJTel2L5ub7EOKvE96bA3uvtG1v11XWfgbeTJfoTEOTf5mt1BWFcGlnRFr
rAwn4UWZ5J8ONKo62sTHf9HK2aYqkakk33tndIT7KqHBNFMDpmMwJkzLFy4F
f4acJmD+Mnv/85PJHgMflJD989TsPotofHMOy66wZbnZhdF+hiXfttoOm8Am
7+fN3iedYhNo9svADLAbqCmh8rjEbnzaBoJ1H7rlr3bBoBtFPqLosra48NOa
ctt38MjzOBUcRr5HZusFffawfGGch7KrdLU6X5bqvn7gFXzEemdf6HjLqowk
eKMHZ6erzuqLl8It3XDEF7Mxe7CswQrOhS9IOQiyuzrsYdDpw/QTCaOjbY9X
Lz7QTtDXySXWmrcwxPqHkmKTxGIYCmbNHwm9oe5/72KtaS+oATc5aJcJMUs0
yRaASznQ0q6nKf7yLoeUfJ8L72qdP6MeV134hvs7fi1XUG4lOSVdXGanYmbe
YoBXLdLcbl8GfHXFkxJ9Q9j8P/6KJ6sj08h4aj5AuZtutsD0d9Lmb1KdY0VG
C8sccZ480MCE0NE32C9Hytgxhr4jzfWNesupmSUGdjeldAj39Tm6LTINkcOI
QngMBQr1+fjo5OS4n0Vog92CSX+h1EUFGSx0xdwtM2R3vO7wGhb6LNb3k2Wm
tYww3ZRAUAxF0NcsvCNEj7rK6S0mFhTCQYtoNyAYj8LT8QphH8fEdzbuY3Sg
ox5ZfA3ZTylnHWw8PLVSA4bFAkkK15kL1BEajYiaqOIc5YRBZsEesXqhcrN9
Qm6fRyPZ2zvQINGnstwvkR5UPH71DQVbYp7Dl5cmNYp0ieCq/cP5NN0hyaTc
vQtcFUTzwcKWjq5h3USjxy12b4ZDQiZobDABjwjKM9Hwe7ffpn6v59x8ETEk
bHQYea0EtAMbFSIR1bk6tJ3AkwGkPJGkDemYQ/XeOd5B1IuszHXwFou2Tp5a
3/d8Pc4HaPK/n3YtSrFVlPhr28o1/AG7KxYSahREmQEh3s6i8quUBmzHizCN
yV+CZV4WbjcHXzz0hqedq3gNPIk4N2wRapuBXRdLCx0pKwkpE0Wura1Q2/yS
b9ExqrMy+1CVIk3JPJsqhARg9Px9gwYPd6L5pUnhRmzheY9bgBXZjz2KZQ3u
uDQSA7fWuakgVWOUVD10sr0wVHC07TthFiT696mcgQdWWfdrK+aHiU25txmJ
1hL4STS+ZsZkREvOPC7q+kkAPsVemk6WeWiqqZM74BtRYTb1jtq1GUn4BJC+
Qo2LHezLuKtID3TMKIaxRyZDf8eb9bUbhPT3FZ8Ym4WkonALyDIEbm+JM8es
VMjUZw7d2z+/lA9Mr+tZFHttS1uIslM/rRKnfTlBPlQC6O9HQsn6+C+bIjkG
9o6FR6+HYLBR9616Tio5QN4pzNaQrvY8YN0X/H2XLYRo9sNrnf3fLYBPOhk5
eAWCRu9a3nuBiU3HSb98lh5Md86YAIB+Z92oh2nkx9920jaX3bAQVY2ok/q1
D17Xwej6WCstLGRsaLwQnlLBG4twjyqzlDdI5V9n8pAJIaxVOYzq+rSwMl3D
0BVcua+2WqYSr4pQuE1dZhkDyQV3Qa8YzsOU3j43of6iPvlyhoOHoqMYtNYa
BOOl1s8c3SN2TjriKQF5vFkxlqdvxaWDLtLhUud+XoujC96LkWrLQYxjiIi5
cGUmD8TJ7SH2XDyPpwNDXmEyxTmfLlbDjicSeZnhZwyt9nzYRUCmTbyeVh/A
OmY0CY60H/YpEXZrR/vAmXxRhXLkqW693HcaXkSbEUQMY8ZMIa/4Ro3TV8od
nGy062ro/DT6SvzIkEmoniTw4ZxMG/QwjVgo9of4QpWT2l81EH3TOWMYrgd0
z+B6IL+5/sdiReN/Z2ufHMzopRnCCBz/zg4eRie+WYaYnGVX9bBtzgFzF31L
A71ZqiEIXneCBkJ4v7H++u/0A/F9m4H+WkkC8N6PMPJSU53HvuIVY6ZPrJOY
qaGMXD4uZ/hcWmO2IkEnDHojj7fik/aSRsiBZITs0HVHuxUexvecAEAOUPk7
skkCotmwaew3ST/rSHShzwdNd2PpvOuowLsYTwo2qObJVBpT3SB23SC3br7r
01znHBI7ai2fNrpyv246lELaGKcZiAXwcY2kPDvaTPP18xCdu6jqTwM+i/BW
1gz1T/J0q4Vu0EhpXhlKBAL8yej30GAjh40wSKQvKm4RUtI2AegFODlZwPdX
aTe5mRn+/XFpJsjy1MQssQY4pzSuw5q/eMT/T7IAeHaRHV2VEwpLLpFpvplA
3gBMOU5X7SdUQ2fomWIcXsFtiEarEZptnyJirJW76wzqGZGqKOcyVRYYXosB
fJs6Wlk62B5eJBFe6OmvecwVryGpG8vAQFEZYWbVpBoTTFWCQnFB5pSPuSc2
PlAhag8AgsOfd+oSxH06wOlOqWm1gq8DB95V03OfqswMrwh0Mor1JenXxDrI
mOvLi51qQpiYY0EQ4by6oKmiDboExr5aErbmuaQec0g7RE95Rss7n6EZpLQe
0pA7Vm+UyQpsyiTq/8+4IHjjPdMqHk6DIF5R4XH4uxzHEIOfyx2m+91R4JaZ
nmrjfWhv9WHD47t9sWjnG+OhGRQ6awK7QS9VbEW0J3i0oXsNHkoSWjYO5NJT
fyAjEouiihUvY5D8VqfZa88UHokfallyGcSDVHJZecXec/Dv0q+ww2nwvYsJ
FeJTu6emJDEA3ppg1c2GfJc6uUjCjxUe2RTB9TjJG2d2WxjYHB6kVGmbKk48
KvpGROoPMmV008wi4pkH+7mZ1ErMVYtCs5OzSBDCK5vh8H/b7qV7mnxLew0D
sDYIXs80UDIu7nWdZW45yC6f0OPbvdX4c9feA167Hj5r3TjJfeX0PheQ8iJn
Zw6hSjZhxdNt4uPkpDadvgKsGbvQ4jdvUssxRf8Vw5cOiBh2gzhRGCTKfCej
cFk62N/bAWzpfP/XP+zR/55Tp/W3YGHm/zkHtJlRfIBx6w9pMNY6lTJgy3bL
eYdM2dYtSFz50eTTop2TXJRCSxs/jiDI81oCL+SnCPClmXVuzRIqZu/OLRNU
NjOTwe94AHK6npPsjv5Af0LnOfdCJfrO/Gy9kVkMUVzhL4zBWQylfXdlZldy
rqhu1wvZKPoDvbhtrzhvXL4JKxyANA53iCPQhRv1+ya33P3DqYqjo80LbTCv
8N08QKR57qPQYw2ceRjiVbv6n7Kdx8tuJ19gZSQba1Sd17qJ3mjv9LG3inNf
+/X3eaDRKbAP2kx2Cf5E0X+QMNkSdEGD5fRbd5nVaKNGSLO9Xwt/G3f8K3He
hllgZMmQ8HgXtWua8wxWyqCgZ9PkazIsKtivYzrCkGTd8SukuT81pKlUq71x
NDb1/mO3GfLRpGV+prjF2Z7fm1pPtu6Qor9eqUe+Q0zRcsXtJPNoquOm5GdY
JiAdOWUB+jILpkYXWIM+xHOL6yUZb8W3dlSsX3A4c/m2s7nrOuSwG6aXP+Lh
xoNZL8PXy8xTxfXk53wHzGrmt+Or+Vo3BlphHHNObKUO2s72gzMlDcmZC1Kr
MQIsZJ4C2kchiN8p5zGjIwqOsG5gurcQLD0L31OOWq4+mXBgcY9IP3eDpYHC
78sJtGlrNG6n3ps9iH9Kpsj6YRZy+6FCa6IwXjqh++ZR9VwkPMqdBPqtyVhC
bioV54VeYZLq8YzhkzqTHe3r5Pki0Dls35u9zRqk1vmayNBq4jvYWYcCQPIR
fyQvxdsSPwKHOnrFr/00fP/ZJD8V89Matf+rVqUYOxMyBIi0L/hby+lFt+rh
2nKr4BS07NXZcIptoj1xAIw5P6OL0o08A8H7VhPUWfiO/gXK0U84qzq0HTRn
5OoSG/VJ0eK/ymkACNYccQvJq+5a8k4w6qepwAa309FyP5SI6O3DiONjrnvJ
jxFQDfAETuoRAarhYbv/BIWh7vDs7Q8WnIuyepPFH6WvrAyB+V4nKh7UlmyJ
sd2Yl7Qlr1Hkdi58DNnPTGakS/ZOhdWWQbT/Dj3l8LtJvgw+B2YCGynbbFUX
6OTxdCckmdphsCEIKGtgiusZHxB12q24ZSx8LkSbAy6R6CWfOMe8ksFgDB/V
QhvveMlJNZxZQgYyMAGNx+Y3TvQzCQ3q5cHtz0K6s9pOEMrHzXMnc3f//i1j
htf1FGBQMhxe+fh6i4ieEfz6cAiC5GAL6hRCOzKu82ZgjUkdgX6wPo4BwUzw
4wTL+0tPgQJ2dyuLrC1lp89RRAXA5XiV0SujMke5zAjWnvcZLVCxfo4Jnu0+
oalT36kKxz0rHNTitB/RwNqG5+6F2RvYNg2qT9M994FZScmHn+Qg1jARuKt1
4u7IBOqTyR7HoH3KKwgT0mvLwNFIisI89K1WqnietfAktVn6Mser8WBV0PF6
112g2Lu0TFF+gFUnLcwfmyaJB1cLmy39kUiFhdzoMaGQfl+vUTWJo7RAhWPu
dF6RGkTl5y+NR7YCkyyYYTfTBpaGdUZ1x9h9l7tdPdB0/K0ULYS1KhrUUm4Y
Tl6xDgMW4u9Svupp7rVRP7QPAya+PDu3rgSMLcTm8BNcdNQxJHeEsEptLjem
ta0nSsYO8NDxAbdD63I4crc8EoiDG5ABhI1ssFilpP/wY3phpcRqn9hKYfSI
Vft+2R6f2uLNi8UkVdqPlYSn6M2M+F5PrmjWdhAoVeeoceWCZHJjfduMjkQw
v+N0VcqsflRB5kAkADl7qO/71872DyriVVosXRK8QmX7TQ1wVBNUsa1FZXxm
K/bCjOoYT3gFc1MVPUEY7TVe6tl1bGcLfsTotqZhltjqfXR0Ta3mlyjCzBv1
+4VUwEVpEsnF18TPaMq74A6CIgGQU+yn3B/75pRROPC+ohrUAtIPr85GqH12
SrQRYsJIPPdnyAQXsXBt12z63BaPAYdu7EfuDRXuAOOCkp/MUVMdjIC4/b/P
ZehwAjlEm2UNgioM1lWyCeTFmGaCUvcwIkanJDJuLc2rk56tSDgh22zGjR8o
2lMNXh8OpLdUFzc2947wjFBjg5hSkOUQCtUBH9uLLPtJWUxZj54i65NiGUw2
T/TamwyEx488GrklniO7AWTeltAS6rGGQzJc8nwkZ1yFUvJcqTGm0OjcYi3l
j4nHumcWl7siwGod26U/1PvVIMsnCjyqm7mxr1xD4EiWRoh5wkYbJEkE9npl
QtuMpQ4LkrL+wvnkxo9+9CW4D7OXKdZs4lcK805kkh2xbYSXq2wiy1KUL6PR
Ev9iR4ZAb3DaFpgNfcK9e5kNhTi7EpZSDN4p10LhCyFPG8mJLFFVq35hCCT1
YoohrKyAAIXULxr8ZOOcArcPii5mNH+DEBIzrERSKmsVLnmkzxktgSv8HUMB
TGMsB7N5IRZ1C4Y8fOn2aA1u/9fBU3uoOvdu2OBpE82PwQmDHTcCwYsalfrc
55dxdrkhWW02ArsK0ToQi7qe9jNWHeI4ctZKUMznOKno8IyNlnXAvQdgL+3V
nh7APycaPFZA59r8mwduX8N+/kAQq8k9xgOvVRDsPHV464YsQu3fwFwXvuRj
6dlhTe6JbE5nc/BGoyR1Ha9pnG5XmVzWe9i5Dy1QwO08prbhqIdMBlOMfZee
Ri2m0Zf92XRnBOcRDcrK3psm19gmAa94bRnOlgTvgKkEGOAsZUcZ2vYPi59V
lwnwhtH2W+SBldE8EcID+bLPERSwQm1f/mHKpZvCPURkunMg8z2KBzuITJys
QKZKQ8RlAyFR2XZKueJ1fUy1/+He42nrVRm6EWlpI0F33FF1pLxFVhU/jVkp
j/l+CAvu+0pSQ6F4XIw8g1M1bqGdUexsJBa57LafbQJy2v3DkCKRcrq5pHM6
jJTBRxHT/NxxZyO/0v5qLm9L52YEXGwbRv/OYqZ8U1lewq9Ks5/S+Q3q+qTN
ubVMEX4GpnAGYkbwjvk4Xe4cKQ9tKWn9f4sFUK4yL4FgxiB19cekO+6ne9kY
JltFQhv4UnHOzOCM8fHPcno+No6XP92S/9ALapEW08cn1BZAGPa9rSMvSWzP
B98uWgLaW1/QhN5Jg1HKXb6HBVfzllSv1mI1EW3kr3Uszk5blYn28Z4wKN02
0x7hzp7vvitLyGK03z5d2KInJN3K9Gl17Q0697Rpv3NfkAQ41FHzsTi/aJXs
zIUQ5Dyz3+yvM11cshf+39v2tTcN8wx/aVx2yLf/vwJzFlmW6UQbDfJejfB8
hcb1MW3LfZrZr3WRCPElEBggMbWiyGnlSB9Ka5v4HxAnEFGN6J6FioYxj+gJ
0uY7oXR+UO9ZW6C7ayM9el/Dxeln6kRjZbbgWxQ6Gw9UtAaFv9S7Y4IGtyvC
W+CdfIoGteXS3ci7DlJCxieE0cvGK86Ls5iG9Yxbx7vKvn08eytBGwk97FDT
fXlGvwaptErFAS6MqleLGsSyylZhQiVlpXId5LTYuiP1XLgMZKU7yxxmMFIC
FGUb8MTisLb3W6zGeDT3Hy3eDG26twytdJoKJnX7VfZxasd/E6NOPOBET4Nj
xiZ1fJ3fWiDBg3YULnKAlM0ut1SM0GzhLxEWp+AWD/6DWMDEtrvWiH/aXCOm
hvSf0oqh/fv+l3na/ABW5109SmubrDs38LKfebNY8PjOUM/2FWOYvrhgtQA8
hSBZwNk6btpm+LuzNuc8PEHI7iNvtlJCkfArwGaWLp5BU362NtHcbuLE/81l
LT7awtFeAMAAGesa9G7I/DwxxNugomVeE5XA8ccxrSjw/ip24ITF3NCdAKvN
shrVMuUTj2JEV8dmSCLthp82fG8g2FJ1+st9baA0mmA/dFmCwqrXL4PRi+CT
7FQgaUWwcPXdHd5cXpOwvQcjHE/8G1E5Gxl+1u7pwx+MtqOi+tjeNFMh+0Sc
EAY0fn/QXtlaGVtKkzWgqKFh6yy93wZ95nFzN0BJxggRh25uJTsLOw7R0oI6
wV8KsG45HWGpoV07r/Bzx+fFlo3zCKxEqMROxSdjCF1sfBK5j0jClQiAFCxz
GY5Hy6Ycf59QyfnAq6Ivy9JkhqW1xL57v5XTD1L+ujcfFgpN/1dJK3immeJh
ly2qNeMvYhgFthRRWYuz798mI4Px8wqPZJxT/CHk0OrFPErZzpO5MOoyqaNp
M9zitXihE6g6MPTjnH8+siUQdzJyZnSCeohk07APB58W5+Xgd+Jdyq0g54CG
7OqRqAxcs9TJS3Y6+xQopr60P7xpe/nPLq3UWhF1EXIeNMpun3isPz7yFH4t
mFnG3owiUsOCB8ISjfFzCt0rxJ8kBp/70LIEEpXJqdHlAeUd8x/QQiPwSDVX
5Mrx2WgA+amvL9+moiKX/OR+MzZB9b4PRVKu2+4Itln/cLzZMxsRhaFcpft5
ggh1WKlWwxemkWt8p5oSE65L7OoMsAftS7Qjm+/IX9s/OorTTLR/jaxQY9h7
ooX62pkaUe/YnoHG926NBhlsNBlZLOGYoGmUNpd7u49l5ryxQlPCI5o84Vz+
v0nxFHrbzyo3v+ssq5Y7v6IBvAxcW5d6omMstglQDns74b7lQh0RXRZJ5AYq
fYbTKwEb/XzPA1ME9be+KEnRqnZ5tnvtDHg0EPvE7GNHN55/P/BvC3hz18PB
8kehTDMbbdEq3QiNqprtcMfIybZvNyxSEDkmSsEANkivkQ8Y1GTcIdE5ebfS
8B5HeGFkSmJPb08iM0TvtiMfPwVGtfctJ1PUZp7fyw25ZXG5yCcX5N5ipwh4
jYdH5p4gEQf/fl9GF4mbCT4kiW/URkl/v5O744PQMOeB3Mr86hFq884d7o3h
9IoqKbdq5xBabpw3e8DYlDP2YxFtH0vSTOQgdzRkhJAlE38lLxRl82YRdX/w
1T0otP5RPr04ZUsJQ8ENXLmNmNRrgRFU0JwHwneHO74RsbpsHLXuJWX+72Pr
Rk4+KMnUj2BHkRkczhbX38ZkEc77nAgCEDvQmQxCPamwQmCpnmy+jc/GLD12
PMFIyrBkeQxejs6ifX1AN7jl2iWSITC0VDVdQRJexwWwHTbjcK6WYfSXfFYF
NOLVgjT0mz8rNGVV539iJpetU26Lxy2ecvCg9P+v/NgG+aqQOkeHRgyMPNmo
PG5P9Jd4f3DPtYxGiQs17CR4KP7PDFUSJKtQ9O8UFVTh+1lcIy4N6tJ9Cmmt
1KFgJaHuYGIOFB5cJo/R1CCUlcCT6CAX6ci/snlPm+lMnbjNUH3HDy8HrRzs
ump6eLs8T+3fJyTM0Z1jyejpFljNv0yM+w+dUAzvHYp2xBuW66yG6/dd+4r+
sJ3s0vc8U8N+XzTP8ftSBorSQMgMhfJ0JL/I/4EaIC42JqczUJhcogVoB2K9
QFYs+by+1nX306w+iDd7rzApyf1YR9MGmPn6c51euMU1L9jfybEV+RNJh1Se
r5hM0KRv5SQmWRbE8xfXO3K7WlHGJHGyKgAjQmInBY4rAYPfyL+Mtc1KJApg
XlCp+XD7HpWuTglXF1otYjmmTeKR6PAqZMN6tp+khTRNpfCHdglFtFrD6a9H
srqHUQ4mNRidSOIEyscEv+Pd/je/ymZ5lVFk3s6Q/jJwTZmBIKL0q1wCAwu6
QYBS3rZ+1t+KIYYHE+MrcsOnWCX4XYLSbD8MGDGC4qmpl+SXDhlwmmx5gh0C
EZpAGovZKXyNpeendImMT58OuoxSmUHsrG/Zbl9ovE101HoBY4H/ighXqKT0
pX00O7pWtSCSIt0Xt4s/YrvkM1VJ/vngPkWtMsfLY3nW67NxD2WkruP5rq+S
YIody26MPFxk9gIYmMyVi8PaKDlHqMQ86QORr3l3Ejd1y63JNG0NYS6PubCR
EahSHHnHMC8gxoMkAZj9WTK4vBVNsWEE1JIVsRNqpkwPdLCT7Y/5Vb4OM2AJ
tomveHyxKwC+HETsTfWIVaRCT5XFGkD2P0yOJYFAHF3g2+TVYp7wN4jlqBpn
M/XMwixiRjEHS3JxuDAk43HXJweLWyXFJDpRNFOJpxrHc4tX3aEcCnyOTpXx
mVJ3R+zj8FICpFfcNnpCF1FXUlo9NcSRaRPjT1Ewbi56kQa9CWsOlk9xGDsA
7Vhue+WU7b0Rnot7CnQ4LTi7vSG0BlQGEa8qI25mug4lMW6ZKri+gdxnno1W
Kl7/3desyyZkA7BOlCO/J2q8DLIpdUtGs40nn2xQUBNWTyj6+NE2hVhv03zz
nLL/tyB8itqOaOAXCDaa8ZpHrxKUF11C7WYsbAZZG312HKjzf8zpEZdZaLV0
FSzKzi8o5vfc0C8R0ykOoXSgxtt44oF5nnuOIYJw1P9hqa3bCkB5SglpXtab
Ob/v7Wtr3FsrRLqnaPYfHnGjuLQUQbqfgnX//vMBZEqj+AAdCv+wFPHOMN5s
jXzuQKeHY2pIf/zyIsK9OHPjE0M9LKFnN0FSpZkwo0mkleFgWgLmWbjzPrT1
TApaG148KYq/qtST0FwkGQd08H/CmrajjeeWO81fDxgzceLz+zUszI/iVb23
KQ4KU4fkqEQI7+DCcPCzp4Qmf0cFeNOwa0Zivr8QGKatp8WkK2WhHew/Ps1f
H89micV7msDERvwSYSEI6120SGhurC+jI6AZe5obj0fhBNvWumyrq2t9C1GS
nOR3igoFNgKX3/V/EDkF92BqDACsCJJuY0gCdoDJ9YP9hTE3F0FyGwzBhgFD
LIH0MOyQ4ybaqiYYcfZyqQtV/PUSsNyZsMtDbFhu1uxL19btJP4+MYmQpdWw
jYTN+jXcD3rR/s83V8hIFz/WcECNb0V0K3dGrCTJmd2dzzmfSjysVLcH+L9m
ArNfi6njSG8+OWATNSU8bqox1OkSGap4r2aIRBANmWtGmsRhZgd5SyAbCXa0
xb7Psmy3D3+bx33a24sIecQJ1W+v2HivZ9nnhvGUrVgWS3xl4vye1MQGL5xs
3da69m7wIISF3KkgULpe0cYpJZCbVZIlvnBc8n+0Z5FGuMP/nDubZ5f75jI5
XsoMXCbrPZkrK3/4Sxw/QNSaCWJRx07hYWeyMMOTqaoB6OXMZtBohGen7Ijl
O2DHb8hNNCPmF/VA/qplH3PY/+eySmBtShCpNBh3l1Ct/ZbWJpi/clNwmpu8
wh2FRDufN34vlyVVUhyvCtZtxS7P9htc+6fl2Keet7XVdc8MEzFGG7KgpACV
8NV/d7CqB/vzWOtgY1S3cVa3LUCIEJXCPwEggL0cg8QJBU72uInlc/aYLy/I
6MM3JBKeTfGVJAPb8lZu8+xhk/7/JAUH9zeBqiizzzAeM3r5ptnJjyCn3hgV
+hPxTdNm70czImbA32rPG7gPp6UN2SXPKU8XQwo1JMrSRxztIRpqS6EvHMdZ
zSTplDxJZhuzUr9jsRfLNTUbJBMNk/n+n/VTBoHcgiiZ1tq5U4IfR7WoYQV3
60DTnSVe2+m+ldg8fPx4/O8BIzh5ILpUSHiSWsaoxwj1LLNGUyhLgktoTh69
7vlEzMbXwsNleeG0gNKp0V1LAGAF8OzA7Nl620zZxpiSZ93WpWh4JTQoh4Sz
vsXrQaDDQ1V3jPPi11F7FcD0i6Gqs+W7Xopewj9aaOWy0d7rIo8pgn0AkAH1
TRNpT5Ak25ZqWxb7t3lBbtPrzWKBhSahnsIWTsI4OCdsVODc4Bu6yGs4NkKf
E4ULvhnz1VZdCh/SVwGOXZQ7zqHb6ddo9pCY94QtKtgdUs/3Lrd1LtvZnFnb
rdAuy8foVOQpQ6nswnqVae4dJHtXtX69zZeJbj4WsRB8m46BOAhArhuUf8F8
aE494SVIyCSuJPBEy3Z0rVXaMCcV05mikv8ZRZk6mx7hBEtqTMePVrA8Ro4u
xlWWHmDU/F6bbk3KItlOzyli7uzIOqrCafAhfkyWiGt2uZ7RoYTupql5WH8Y
Jr4lwTa8/UypdjxiUlwN6g/VVqfcrSwXOciyemgjiYFVscvJkDots/dMWeLh
U6SYlvXZea49cM7Qb0astwahn3fu8DKsKL/9ALpKZnEIWplmz1l9x1xpmRUO
C5bDi4wzlVdSic1RS5lXMShwVdsP/jAWu7xxArTeNvoZQThYNftDEpciEZOV
XSaOeiXuCg/MEfwE40VXNw0IpBRP31GAn7ZMMO49PyIB2da9uJ5qAtba3755
EDTTzvH7AK58VHhbNuZ7V4VFlw0aA6AtNdQ7qFxBcqiQG1mymDYOlhqS2t/y
QemXqLBN6SSPwfXINad0HuF+hFjgDKgsHjw4WClyIiLKpfwmfZPThhWg2bYS
VUYtgnHNX+iv+3w46wrrjpsxk5vqMV0LE50tm9dE0vNGggjFQ/BLuKMPA4as
dL5f5RGU48G3QHolDti9+MHylsf5qd3Lhp6ZaXGds3fY+gpMpHI1kQkoP8E3
oDqbWbShS8d8qg/Phmpmr4g174y8INvycdREn/5vb9lWazrlCQ3U2WMhxhCi
gHcnCMnhNyI11OqBpdknT0VU8zjtnjmxD4Rl3sumNtG4XpRvbANTzWsnNldk
1rBY2gRFpjjzmWXIAL3iZEWI3VtDJyZFr6XvpHxQyH+dEZ2f/Y8ke6h62oZp
KqchcL0Dv7Ug3bqOS/cVrWk/0L49yqCUGgNt4EDBkC/6HnvIDjGhG1d4BxIE
P/LPqJD3Zy+RYa3le60yIpDMoTIthYB1jIz/Ch8GSFM7M09PJ5jVSmFVQt7o
tl/gHpCPnJfBXV6FUEkqhJ9hKT66juuPWvr/f3KjXI5Wri+iH4NkcRL57TVy
7GTigMmVjxHk2S4q+WXNk3NbZCCq4eB2vLMq1vMeAWd2AyO0S+Ajf2KCuHmx
mSiZNSFDWIBjiSZCFiR13DD+KC6hsrna1P1mNZSFAc4Bg8kR2TvvHXS+pJdo
4qPhrWUGICceI3AHH69GdVSau9rVfZWu1CX4bwcMPDKAeTSZMYJWXEBcmnQe
+gFKrjCLGCHI3BNCOn4lE9rmGUETlOqpIxJubvUKBAx0Gv7GV8llSLl5LaV/
XlE0vsc+YwHHL2sBPTkhTq9gcZBBMH6InvvUN5NT6v5XnqUn7W0pikGd6M7C
pahfolQS/k2XTsLM+3J8dRZk6BwWZ5JKEV3Rr0mExqd1MjdaYch0WQiiUECn
IPW+NKd3ZnsJjTotSqZrRc3xADj1JHKQDOpNxQqiEcF9HtCt2fVyunpP+uiU
CNtYxBOYwRVyzkNW2XZfw0V6V5H8255uXGPPTmpoRmHOjCTQjTMNpMUQBsHK
1DzpEPxC1z1A7rqMGuhgq9U0d88CQSK/9tigUVQWHx9kUqTbSpfwL3Ecrzwd
Jk7u5OiQqGrvuktTE/NLZkDjS+23H+7pI9CQiYDpmg9Np9GznpEwrYPXyGDW
QUyjmPpsaU1pzB3bo8lKufzuulxE4tmf4pArxs9ktDnxViEO81MEeHe/8otw
yK4c/51mwCUn+gHOisSuoutmc09FbYMwkMtMVLbxIPEBTZjIX0WUX8xTgyNi
UasNsrN+BQwA2/yOtulQlOVZ2pWqDlIgYlEoWZAnQ4MasJcLUDUXy9hMap2z
lXWXEpmHhhNRcLzCgTkkpERbrl1t8qgQUEoINY0reeGyvdqslQwfDB4CkpeL
3X8ev587pboUFPg3ScIpAC//f1uP7kWSTNaSJAslzo9PLQBnYRPB/Dp0AAEZ
PzSy1dkR5I4Chz+1lT9SdqetbnZJr9ijn7kMkAy5sU9gYKcrbaH5J42jFZ9S
tHE/55JxefjHi+1PD8VRMPHnQj0iL0364MCaYqCCRDGIxUM42+D/pl4wajXZ
3eCWNYow5i+ugQtQB02qXu1dOd+OgxUUum3nLfERx1NbLeC4nmqBQj8j/8Yc
3cx0DsGB2S4SqroGLTOZn1RsP43pvP+8TZonuAflPwLMu7ZAh660pJ+8lioq
7UGLxrbJG2SAdlKWU5ol/WWWh39nSeQJC1F5rTccm++PWp+Mm65MLCI+3RDm
75LPPmYeOfFloLLIZLSLnW9GOLmRWCzP+BA0GtsxOCuB2x1g0vscSdI9Zw83
Ce2/Zs757zAQSGkGy4BiIymwbdbnNidBiJLus2bIyBpNccPtSliUWwxw5fPH
Kqh8zxBEESPWMl7hI2pv/0OQYUgR78F0S2nxSSFRQ1b6Sodebj1kA764ooze
Ji8Sju66METMGcHLiOdVyPD9UinQ/7+aOynSIHx8CKSYYn5FQMlu37QQwWtM
VVlK+4gIobD3AuoxsIcXfi2sCXhDm7yJxhXl6/cTll9vIbfbj+oFbNGKk1rJ
8yhnpy4zdUBqV33Nqm5ijilXmWnYTBnU0ypR2qEAMUCgpTeQvz3Td47HHYxH
iq4aNd5QrZagDP7pCjWL4E1XMKDXmT7aFMRNkE4QRLdw9Kj708XQagLmj78I
ahFqnLtZNlvyE75MhXk/MyQpMx1Gg4AmahTaLfto2bVJOHGY0INiINe+empq
ne/CECbgXUPvFTZZboZoLglaPSG6abWzBQot89UAi9rWZ7eRTjQ4o8Ie0H/w
btC4g5djtlX3g9VahX0ofSPmXhL99pnJ0o1YKbumVx/Q9Zi1bgnCdlYckZy3
9uWFGKI7MPf1wP15AWOuQxwMo30TRFmo6vw35aEaGI8zwl/MoDYYll2Ek1Rr
gjyNX9iwc2oLS/Ek4NOrohyNq18GZ62kkeZtOoDNn/GQ13HvvnrkHTC39O0S
yf/dBEuJXFOOyo/Kcmc+Y4WJEk85Ukqw71XJIL84/faDGPeyqXzjOthCqAD6
e9oO3FQaQAwchrlb+tqNYLwbHk6dWvPYm63863GnXd3735IY1QvcXicgF9D7
47ofsFL5xGiZHeRtc7vjbUiYH0LemN99DvaSJ92l3pwCn3pMJljwz8pHiAOq
yRfJUH2GHWTrWtzk+67bNAwqmBGIHT6sCN1IphmC+LsF799OBlbKaXiVFC7o
yYJqDWMQdQrJOU0QAhvIbDB0dvl/ibSHC6boqFCffRWe06j2Jt32egUeccNB
lPnrPz1nlBXq4Tksre2NPbDVYdb4n5kSk7CGWBnES0NJFCAL9rIzCxq5WSGk
oJMWBbm/3k16hZEGqKd+KqLQV0Pjzdn94cdSJT1+3NhtlmggvePi2M/nIhFI
GK7eCOE45pjOkKjfqzbxFzJlKvBSu3S/5KLVqKdzmN6gIi3AGjDtHlaBnBN5
3UaDtT/DaYIMQAPpHJN1T1qTbdTZM6AYH6ioKxMsmqGzZZjZMDfQJ/u4qFNB
/MXMc9VBjp8eSKPhzjNjvwoh8UA0ujs9xuSY5tzfuFuPCsVgMrqdwagHugmn
8hO9r2077i4uFpG1urnxkd3xLSKwCxeBOROc6nlOUfve4hb5axsUD24+F+Ft
mEMYewItEKfmSsEOT4Pqg5bd/3n1ei8Q1q7ELayCXUANnJ70J9/XNrqiBxK1
saV3AVycu6cJlrrrnbjOSzHSDZLm7SW2HZ+Y2jgJy8mdDdS8FNzYJR/Af5H1
zNlGQnF1+10jLBtCnrXca0LAEfCDn7x186KBimjDks3pycNu+gO+94sAg404
vpzaC6H/l3El94QQREmTOES4z5dKLw+4v3yrnQO4dHGTz8aL2SPQbm9Zx8sX
v5qJZaIE+2fXQmV7xW0sLMDJGcCHxv09Y4AFhzw/YpLuOa3kwRI4GiSqj9hp
X3e13hrF+qG+kZEhnkOL4r4XAumYfxYpWhxbngrIxaCKJZnGNFY7X/fhwPLO
jJ9Dh+5Nfq7kYiKssOrQEWXlRpq0yF3GRT+S3AzacpsDPr6Sd43v3xhJ9a02
5UksJSFdn6dlxYK9IRmYGGkUwymCMX2CFhYPsVzjTG+io0ZXbEn2K/kEYPX7
f7x5kcYladUliBSpp6yon3yFZ9ZOHmZ5fMQh/gMdiLQvXP1Kad67cOWMI7yP
ChKdy+ULTV7RIrzXRZv2baaGHog7iASJWasHwtMqPoI7WE4o9L86wixf/YEB
Ve8H+U+zYo7ntSBEFPDWXFIqA+Q3TZw4IzhS2K99eYMlvTvlnbcedRwOYTK9
0M1QDArlmbs6pg37Kep3rCX3iiZerDtidvvvH+E8ppiInSRymbWBVYAAG05I
XWIT3HDzKiVeGmTIpbJwyO+8Z5LZ9SjvMZiXtLSrGdGOiFk68pNw2/v9ckuv
yF7Wa1DFmaQKemKqvVyTS5TxDmbtmFvibIw1HhWARSlPZVS/ex3w7YnAOYOS
SI8yUmiaFrGTBvmmCaFq0pYxziNWAVanNd199JH6/wvz/QMafuJ/slxGkIXR
bxTjs3O0aIVxQEMO7GaaX388y2taFLRcJjPxmLoz649kMhKVbnwiKEUw+sxu
UHn9g9UZseUrZkWyDciafTN/UzovuSQMN1ueKnE0/VfSG7OBXCqs94fH6faN
/nxzRDu+DKCXm0xptfGY+JhLOjx56SIcRYx9F5W75G66t+g+hU42/zyLhnRv
OXfx+xMP7axvJ2aBgVXErqoXFWusMdC0f65/ifOsTOruf0GfIvwYhHhmgZqc
TZFbfTxl7hZfg9mjUDoIeSPoUq5ADiIyOAK37exSEvi5zkFLU4g4UeporYwO
oUCgDaNx0sEtt+cfCxfL547WRDY+Gfyzsu0jwH8Ax8FL5MVRfyF70ZXmjarB
lphswnB2wfOv14qAN5KT3ZqKr09DuwAGwg6u9+K4MOmUWxETvCwFZf6hJr/c
7TmR3z3/PPrdG1kjoZi58BBMg0ZGZDEaZFgKEnC9vTjx5V11gdsOQp+xYRLx
RPya5T9dzX9zhdGlF331kviXmqHscWMmQjJgkdGuKqF9v1buLDxmbIuHzoAQ
gDp9UO92rZPDmYf4x5TdRUAL/6yB4qrrj6FDkqgPfRnT5Kf88KhZLTBKbNU5
fhqDrOne28wwgxDonQQTDdUsEs2dNDOYVhc8DhizWuxbpk+znzvHN04izSio
P//ac8ZHZmbU4gEwyArcA/N7xzgoJsrK5K9Qkm/X3hfom8ZZSvE0I2JM2YC+
MZPdU/cJDqp+vrznB7hG12z0gChvnZpnI6FWCSN5X4ddqicKxk6LL0kkDU7U
7jpEyY/ONAB6QkoHG3EMVLmT8eugz78i9Lagx01Cmp5WhqIJS6QXtllRCrMI
+aNrLh9JQkPPItY526uhjMHZJWiOmXgRm4PndFN6dvyQDirC+QASySv6JuRb
Z3y8Nd9zoaxFzXSknjpK4XBY3AYtIdw/Nokb8wnePGimqHhK1i/qN5T3lg+i
OWfxnbOzOlOu+sXIC3EKeJ2Xv7cnnraXxwKNtHu5qU+uc72slE15qAflk7Og
kdaZ6PJrMnm1DCr/iTlD50IbhunC2fK61/hhCJwB9Fa/GBqFPYNTh+2JDyl4
ygqOWAWL8bwhs3DjU8qvCDUvJGw8GsQn7LBbH/aPo+jO5kLB1YgmcCU9GvaU
FdQszNTVyAEhomOBvQNhTIcW7Gh9D0vTxS9zEiQVHDb6L5sJDkz8MKDKvHE5
rQbSF5bZ1CwTIPKb96p+eggEUJUwhhN27NSJGmDMP+l9msP7qBwUvcW3siVY
PdUjIC2Lefv1J3TF2oED2z+224xK5qL+Py248mExs78D1kDBxtGcZREm3tjb
w7O8KwqFVF9rPNC+ZJsqa2LpEWPD7rqNhDtzA+OjBKLDMyzC6sdeYczALsm1
tk9PrTdAgoaQUAQ9cFAukSfG+jYnZTXyu1CPNjeo7EG6XUYjZbPblx47ub5t
EQb3BxRkafTKZ4EKBqmfd48Bdp20TSgM3ar+pTXm9WCgMMeaaBIJaLhgCD1k
8wvkDANxOiF2YVIip1hdWM/1EFyGZyghaapL81/yy5JY09b13z9aghg9snep
mXB9tgRxDl+xok/FYkXGW1/QZNFAQSc/3yRvLleXQVZybK+suFGPencmPXi7
YQlJ4FD2cV4606nfotmvCDA7ZXC1OiNS1uCy8XNzKLbrd02NoaxjflI+10nu
xH+LkQrBKUHIdYlSuvCIi2O4nAXHpbjZU6FnvN58/HEN+HqirbUcgdJqtQxm
iari4wIhTcaDQ/bndR8qdATtoVm6KAEj16+DxZ7fUKPu+DCjG9bdc4XeOxM6
ChcTfnujWjRba0gwmesk/X0zYOh7vhuV5gk3lmwkEwc3OK5O1+gOzbNgTN/i
I2KFS5Vw40SYId5GwF9MCGRudUnI/DCkUJ2UUwLJ5aFmjhE+GeWunRbvK3u8
VYdNV3HE7lpsBJjKywvBolUj9MaUJD9dQViZeYHF4WPBslrp+ileUi3Rrzuz
rQmldZgjpM04NMrci/psJsWKrU1Zd+CN8oZXmFsfLifdHCKg3OZZSIjcThED
yC0CUu2xZTAsO+9rCsgzw4KanDJCqnXVHMqK5nkd0tvLBHdNcdIusRKN0mkB
RAhIuz94ZkRK2v7D0FbWP7B2EKHNH4q5IchhDxOUHr/6Q4knmGuxHwTgQ3J/
oH/L7O4Bk7ldMyRSHFRMyPdRkCMsT0WuOoqTOsSi8Z1+wBqV+I/2eMzVCo4d
x/eA1iPBSMd6h4xo/xZx8IAKya4r79dk7QX6bj9lT3bKd5eOaYcnN8p2VyNj
Hjq8+dvsjgud45phErwemhx4RgJYPcTN/HS+129DvqPRnqQUqGgqnxZx2MyI
QEUqNMJM3jsh7AV2txYE1wYD6cFYHL12+9d6O61AYNDPIx4sPlEVrna4d9Py
k3wOGU+MJ6QrfMeFhYs8VVGnCaO9Zkt9AZuQHH9IMX3KhlJxE1ygPDMDLy5A
VwpQtxHQM9szRLVK0oi64am5muOMCprkocOY9vdgtQ8QeF4d11aJdU3jlHOI
Py793SRZAoPHgEOSoo945xzI7zfAv97BErCbJ5DG+aqL8th1zRHdHrS7tGH5
Flt73veNFv6Gy4MEC7oMk/2rDOSl85EwzFntXye4sGE6W/tCzDah04WhZiSq
kGkr5boD78WZ6u482zmIfGo4qkerrL69Z4+2JjnzzjDsuYY80Tw7a4HctNyd
gzhBpEkLsAnZrK8eHrJGXHnhoaSQVoTUFPugW2uWM3lQrYMyVRcA7Ll5SmwY
OuFbqt3rsoTjCvclAX/8Bj57CBku2p6jW7C/Ri1TejbWhV0uHo6si7FoLRrc
cYMXPBbs+daemRCCgflUmevaYmes1rX2gDFpJSmzfrrIi6/t2SWVq/mvHFnQ
qe5cIqNMxpfcIVrRsUjGuy9/vHnpvAtD/H3xHmFlP5xmcib9QZhOR929+PW/
1eTrnEgAwezJAO3hvtSxjYSW3Ia9Pp4EAQXXR2U4zsCyrvYESr62SQpNiJKg
QPzP/k8Vls131HynCBmH8JI2QuejJNvjBjdnbjBMjzHsp1VHQZpXFMpOKAqn
z/45rVHuKR9QvSQSo2rrheLjTVerjy6gCh4nOIQsslxmZ2JjPMixwD30Z2E+
cW/1ZAEC06BieS/U08zb8byNdNc+JsqNZMqsxB6SpR7l4SR5ig4e3ip2CSn3
+352lB5DA7d3hwNsRI2o1mUGLROjNJyF5mvKG3Nygsg/DkZTY3iMBwigEx3G
zwPR+NE5lsaVIAN4BpWHtTSY/UpDoAXBA3ehUChYxjPCXmSAQcduuxsEDnje
sZW02pG9W2xCvvXfU0DpU23egfWh46+vkLXt7MuNwBrg+yjERTgpWSD4acfP
xe/kjt8j79QlGM5yBFDQHgU9dlITY5En5G1eT0JpV8W6Jf6MkPM32ZQ69TT/
TIBsrqF7dHzd6JOz6jBIKEl9Bd9M/tUXme1apCtZdi4EqXf/nsRGpTvS87Ek
3cGtZb2KjGnj52XLKKfb5Xtg5KrYrsTFQouhohGB2aQo+ipavatSqFwTAfdt
5pkZOdODWUvks3o+HnSyOwpnOk3p8WsJMJAnxiNkbeV5kafHVnIN6Uugyo2x
XUaGyIDwvihylw5tbJcmpjmu7i6vxsXjcLTE0o/6F2mL3uCALFSsL5btvo3b
ZifBnDA6L7dpb7CwiVrrYa/3v1g3OxTMvaxt2fWgoNHbJcimyZZQGF+UyWeB
jv902bFblle+1BCOimOm6sutyogLCwEagk3tqBCvDrPm4YnGXH2W4wnVVz5p
5RgWP7SzpJqG9f/1d+dNme2Gf8oDhwmZXVFfhBdoIkkycvNTve3DxaYXa9RK
pC0W16Iq++cyJ52fA74Hcd3jSuZ0/hTSfIzLouK6ixH9ryuoL+WwTO8FfpT7
FeAVTabY22DEeHREmofMYOP7e6rkYA9wr8EE9Q4al/Nscm0U84MrJiYEX8id
yeGV1rZwe4/i4IeRmgLxVH4SM+zVd2ARHH0zusrKPRaM9BJKIk5/bgOtUdI+
B0rbj5Hd9PMJguOhhvGWtCKhI6CFBsLCkjB1vcJg1Qnts27tvdRaNIk7kJki
+Bf7wt2SJa+zGLaYoZbMFATmuY9oxR0s77Kw2KH8yKa+nCTZ+lwcqGyXxmw0
KucpGJkJxH+fC1AmcRI3Hsec9DuzqLQYv3OKW21+qfgCZaCYTOWxqXWPewiY
nB1PvwPNxCrd+y197QYqJlRUzQVhXFR40nJ38u8nakIw6AFeG2ygAo/NgtOz
/vImWHZzKxVi+cwdtN1uVhGcSKTGp9zRBis2bXt6SJBsnLV4THnOydU0R87H
RAaIn90QvUfhgEW8JmoQN694DvMwKDHp6Z1TnIt5Lq2Vf39z6uhizlKmPg7j
i4DSgLQicaGdnZMlsxIyAoLuzeJg4z6r82D0OFj56nKOd3D0hnQCVfb9nfJN
buMi9pUjw8kup1sXjvkDlopGPN0M0EbA2VxoYd7p3q1ZRjQaK/DBPei/1jWn
xrnRYXvt13euWMKG4l0oeZ0uPg0bLkJiMWkkc0Fu+slSL9rcvuWhoI66pVdn
Kr7LhVoFpELbWxJnJIALtKIDum48T1Sr5xACzzmUd5iDGn14V488yGstLTMc
iot7IyBDFwp+OwcKkpVCTBr5+Nt6dnVIDJu/A+Kg0j2U3SGWh31Wq7mYtR33
0sD45nZs2ZBjFM6e3y7yBtV2ZK1hCVtHD5gvKSvHyg8tt1LluwLofUnDIqdY
9G4cAoo3i62v6eXi9d0tnSGyzKlAO0BncY7FxwfleHi6OTqPLXeqSvalMYor
ql7kKVwzjd/AhuOKUjX7Y6+chsk8cVIWgEoOwveYd8iCjeOnDWf0Cynt8Lbr
NIKjRQJVeBz3slwyBDdKIBpYgietzRuEWk6yivaqUA0RCNeSxnoIRKmQVH5C
kx/ZOv6p+ikY3r5jqwhvXChHpCqmOnmkdcrJ3Bw0Gg8Vsdb8m6zMS/yA5J90
hjeFuHP3DnmuwSlI4vjmvUk8mbXQEvVN3UqbxawUzoRL0QkfyIMiYbihMGl+
DxYb03TlPg/zboFLCdKRrIvTrm05wZmHsH17xKx25qxuQjhpNGxUQlFEIDmF
l0O+zBqGRM0vt1lLArUd/yu6Vmkzc3neJ7lO2HogDD2wBxa/D71QcHKaGZ6I
N/xjWeOBx+cxe0kS0kKdqbxEbRnJuUj4Soricrt+llXPKMdKUo3skEBRljp8
K3MAWkyFrfZnVXN5Ms4f1GPZf2MCgRKPwvNm3Ss4VKs6oA6qP+txvaTdoKdK
m2AYHiMu4eqgpHm+V8d5tgqSf3ZcqwGabm8GwpzQZRjeS09aSyv48hvtSrJm
jeFUbml2gyJtD8Ydc6YhXJkoPz6O6OpP5lxNG+UFkM+9ucmxVuDlG0QPVg+R
gSwBqPryoEA81jTqhOcOEzx1ru3z+swmt9OBw9ntt7NfgDqjb9a9ozWG5Doa
5r2mqJa+K4s4XQXSnGTmZG5qt3lSVfArkSVqkR7tRv/BVDEZEPfJixRsAB97
zozvGT+kQvxTHdUxjP3pnqaqdOExXdUGFHiGPO3cCRKUlmH36tiaH7QWe/M6
xiwZrbExYrv1fZoU+GnKJMgyWG+RiQgcB6HL9QAAMCoSBZDcfu+K+8YKSQTe
UAJ1Vseam2206v8IW0LnyLTP+TPVZmA2YiXwfsGsthacz1hkLwiUH/Y2t4Mg
TpEETxR6xgEguL+VR/DQEir3E2bwWDrTiqlfWkXCgK8uP+VN2neiE1573Zv8
Jcgo9KJSGswXUebIdJjm8AehAon81eCE8lxY139/qPMA7GiBFCJ6rmQiOKDR
X0QMPbvE54+LI7SUE2i9lJIIRXMBvuS0Gpn2uGV4h3uFs/xqT9TEmPGHafCW
PTCh51z02VE8JGqkJUVPfUIVZ/X3O+nDAnoEsdhVkmcyC0VT/k8+KuQAYrHY
oJ3lCOlSpa9+wGNafYwVnOvbk/Dq2VisdOCpRpEIxL336O5Yln6sYB71vzYL
LzCu1DAPTtGo4KkmAW/vouzvrVHaPuZF8KA7LZl98V0UeecazeWdozQD/r1W
19L6GF76l+TSGhoNzkZXofx6nsJvEU1qYLST6UEOLHLMwxey6fa3k2+ePyk/
8XnNkXMym1Z+UhxE/JVRNyrRlq4uuHiSnQR9OI9AB0i0vz7vosi7eUx/Q2Zr
g5WGcoch9mxcJs+OWhKhvEJ5UTA6NAFEdRhvmb+Nas1DUCJO/RMSPw0vW/8r
BNAVO7aRrGtWV9TKmTY31H9DnJmq/06sbyn8Q4gW0RKi2zGkGhJTHPqLS6uG
9Arpx1H7FDoGgt29HvrwVgDNxAaIY/qzvsELheyyqrDhWOMLbrG9xy4dKBNz
S/gwO1RIpaOilztif57RXpv0lDniLD9irGFDHwg6JG9EUcED7gEySwtD9UdN
DeOlqakXOVqBS0EOPY1tx6jWx8LJgXbufdt2kmy2tzckNPtK+/9GH3yemjV/
1P0ZZKbm5Gwgsx+PVKfm1oKlY8aq/Yn7IXyoZB0M1k2fuMcYda7d48WMCJWU
I/QX6HPxv820+cJ6SGub4ppDeAJPSor4dQhZKZbM/P9uyv2wv+T7HpDMHnC0
iJ8s8bUpC7FHZak2gPRS2/ZJqEPJ8SWv3dIDJ3AxYsSkHhFqc5Q0kzPdINF6
hROP0S0rhi7usc+RNfZTH3bWg/+04LNZFnAOUZKdKTGytlVpdBAzloyyc6qj
h0JKNJKkB6HmHdr0UCLj0Wcsm7AwhMtTF0+0jCNquzQ9hfHd7jTvBVkJqKhS
JVOtvYx7s+xGMcgmQAx/uH2LAkriwK79LJcmbgUjpGIhQTbkEigpukOLBily
mCG8+v8ibizEtO+k+5AlFC0iAO+3nu5dGUzIFEZ2mn+1ljoCGcWKCyauTTPe
e26zJYLEpQKuu9f6EyB4eZe493Ya9pkb3lCB90N96zla0mkoctewiktxoNif
KWihg2wtrhmDp65GUd3ydUn0NSj1kYBMfaxkiwSpSJ6rzlCiCTnm6PAvo2NW
/Dwf27F+479xnQcYh1DuTITnLN/ZZb+0ieN6fjEhUOIg2faEgVhnzKeDicFq
RTxmnhYujzBu9g3vSh1zXUecs7Ukhsbs1PKI33GAlQbl9vQ4akoVDrXB8Qgf
MoP0dZgoCvOg77DYmUEqv9FCq/jUloL6zQTFcqxxkDwVwVQcttHY2rk4d23s
19QJ4Q44zg8zT0/7bkxFjakWmutqIWB7o9liLWbLWCch3KZY3JuCUz6bGtq2
bQQF+vqPi255zl9hEi3B2mU5MRyb6OorWRCEvBSdml9vjZbii61ntkUM8yia
VPDifnE4VhFPADxHet8HGdqH2/dCnqsSjSFmCao4jFKi+n1+TAyYxiPo9/pz
+BsBKKDuhzPEtPWtG6NvnnYUNwsysGpxhqi4hX8niuR06Fuhd6UuaORuzld4
2nj1TF/Plf6sVHAPYeYHGCjptRJ2sHIArZfdyj03LtcleUZbY36xfN5BbRlx
tphZ5Y5va+ezbm5gdJ7MaTH+EkTsryxWxTTmMzrXLRh/CdKrrPf2vREYbQAe
67rKaobM4YhmjP4G7R9DHwEAYMt5kZ7it5XM61FE9U0soitcAmZNWkE4BUmV
eS1w1LR1AnRbbXvwHab18M8Ms1IyyLvKYpRmL+qGwL1N6xuTGBvchhLpxv+t
H1e8BI6EGCtCvGc7rx8EkPlygdjA0ncnhdhG+mDldwmpmTF6r3JgFeuGZdDF
mpo51gtpJ2XQkv8qT4E7/uTjO63rJJxxZD7VG5/nmDNMokWo9yEHPQ78LOda
JrMK95xNJ4/L7kDsDfe2rGaunzNKYOaiMLH4oVVkA4R1XvoTFoYuKzuUKqoj
DkbxVNKBBhlz7/g6K/uYSzWGDUAZG7bi+nwBp5sUZyZSDe89VfJPwacjJR0E
Ezr7mQicdS+mLginSeC0x8t9HvDFRErLLw277dtX42pNB38XSPWBmj0Xi84T
ihmsCoX9YdtIkYrsAomI9bBPejveSOubdqbJGuky3sCxEf6A4evwEmqYI4F9
OfAUoj9pw1+aWciav5mB43lAYLFxqUWjLE49xSiOyAuVUhEQFF9okAUAzHOw
cuIMFCuMUfnsrZ28Jpqejzu/kbEs2jo0Os1KRslEaB//nn9Xv9sGNxSq1uMI
DNrlJXNWde+qJBNuMSLRJplF8WFWkcB4g1czFFxAwI5KjGvhyqPlfa+R1Qkm
YpFcT3p7eH5j8Cx4Q4MuETIQ0zBJ0XDkEyQgbcxMHOAtljpB060FO+XdXneB
f0q71/fQi4nBrKSJe05UIHBpdPh+RioiCC8ty6JRBnvyPppk6GOGC8GBqI20
ho1I/hU/g7LLVuNFKeqgdZc16lkMjvJ3uelepqdY4Q3xZIVBwd+dZrOzUkNS
KOI237wlf/HLKZlLP7gva5Ruy1BbdaTjsffnjC6+FMa/uZGZprdRpKMeu2rT
RbUFR92xev5zUKKdAx7i0sathFh/1K7S+dj1X+rxBeVLNArQFfS9kC6CDz2N
9xMlNl6PR4tRLgBll584ZPFhz2rETBcNVsyi8dzOpcZpqW/zOfLTDiOCH35R
WFch7bd6+in1otorOP+QuV8NpQcI7GnKqUS7eiW0/TCVvjpSnD06bxMn8l1E
qQW9Yu4vL6jrDts9F/yQPLfDWtZtFCTBY938Vx8oaaVkJo6xoHohMeY1p/4/
LYmSfWq/5BTk/UIPhFwOeExOenhqWkd+9nOCE3U1FEXqhFh696ULzNvi8pyr
Sdfrej9AMaDmb5U3kbuTRuFelOkUyK+iO3GSOSufNzwpkIAHMmWx+Hp5GAcJ
zioknatS+pS2LrOQa+PP61mZ7s9c868CGhive6pJJcU97WlCw50L2RbeJFip
UyxeMC+4+h0I9PHPgVo1bksiqocpW52KK+YjzIB8BBKk558w5hX2aEZTKtpa
0/GGaBDlSVt1WR8U6aAYKmjH49pN+ZB/V5EaCKjk7WDz+0x73F6oYzoX2p1d
CdovlyDdW+/oMUulpj0AuHbQ5np1M6U7FHthsVowB+tcTIxxQyDxREL7sW3x
n0e7X0u2kGv/k6hpI2yagQnsAOO/Ssrx07IrOiaVUVptmqxuN+nosqAjDygp
BHop6SWqRb3x9a3VlYHcZWY54C+bExQ3T2YZOtIJ6Jfl99CxIog5jVzqX+Pi
YGD/Qo6y8d0Foj0ThEsgU6tvvfB3dfOgmSAj96be4EN3VgXDncbD7+OFdilq
dev63R4+De3ljImGIeKq5o8oXnmh4BrIWUj40rqx0Ou5q2TXVjdqQpZpwsMp
XdOk+rgHaVsjOHTz7+K3R9/6hd4weFivkF7ErhWjl0qXdtb0V1yDvcYM17GS
C6mFgKqBEGGvvRm5zHnig8bYq6DiykfytlzXOzxmq9Ozxqbjt8e2FFQzFJfk
H7XcZHJPt4WRPaqQw5e+3gcZflwDoDltcyGXCg7u0IkdmqDhD6GjAOcYyAKC
MoW9ShIKIHOZj7MZQXLW0LvkyFtlb/IsCxpiG/73zcZYVod9cQ1S6y3GDeLf
pM8zRrHo0uCYYbWFtcgIIeu+Zdro3Dznz8Ni21bx0A4IMetug1ScA1LbHtwf
cX45ouepiqkxNxL41YrphMR2cQvXx8/YCE7e3uw55rLiBMZYAPFabEQDuRlp
zNfd1l670sGZlzsd4bbjmjmsSvlkVqoYlijD7Ei2ao13a6/dbJ8/NlmrR8Xf
PMAFhpvDAmExsKfYT0comnSSBoXdcZkmY4pzFLMKLfzhux4F/TYzYKpX/Uo+
06hTi3bxg79X6/zxEMMIvoBWouwvyeup+NMp7ADMud6lXv8EhjjvOIwmlGVK
zbAC0i/FwneeDyjMC1AAOtPODw2jgTFyiCQiChXbuTxgxSzjX4r3YEiqLLL2
kl1L/BNjsimgQ+8z+L0vk+uhI2omnA4sOApAthb4XBQ7rMjtpsNRRAvvahjv
ozwwM5cU/KmmC0QFV9bZywkXbKTGzbXDWCYwm2JR+2mWXFbWM/J/i3SiA12R
b6ezbzSqSpRGVd+/5hC038sAQCl+7dC+cg/EGQ2TNg4oJmc6VhpxxrGGkhDb
7cp3JJpymhZM06o6bjiATZb5/n6j8ZimaLUR1DIZU8EKMoYickYWEkMk4I0Z
938D0b81SoeKlHRS8OVfQQYJ8xPGJ7xWtWgCUxVCYBv4YjgBngpIqyAkgmRn
Y6nZtlIfobtK35cqlW3rx1KxGYpCGJeICpoW3Vl9h4OyttRnS4YAswhEKxsx
hg6LkHQ7+Cfhr83RORafR1jcJJT7FelTu/iTmxAYI3otzJe1ldqOPXTUjjyk
txko5QvAEzTWEVmgpf3DdJ8IHI+zyYpPqPqV555yAPZEuC4yqtGJdfKClyxr
3Z3o7fdmtdiyIXmXh6BeAksm9rJ0MdHq6SJd7hW0xftAdMvuTm+95sd+nELr
km+dnvPnMVFH2ynTlJUgqzybYH4LmLDZeBApMh5Kow3qw+1wa+YIjU99XZA4
gYaUlWTk+67Ga/GAbC1uiEjZHBwlhDZSCa9L//8h5s7QcExNAw2ZG3YL9gD+
cPsFbdioMaM1LtAJEudhuD1fX3jNY9CIkRi4ukMb28hFP++jmpSrA6K5lNAw
+R5SfpgQ5miGeU/kQhgEx9sKEE8eempAMds7CWICwgeV5H8+vOXizt38QY1V
lXdg88/+CYoglg3uy8s7MLEaRndWWHjmvfXpYrU29I2/DPOuNhwc22j83Vce
FwNLxmagLP0He1o4sY1iMfKXXqxf7pmVHeoSG+Xi/6LAmnEa2th4u2Lrw0mZ
BrnDnGxoyawTiIGhQ0r0yGR4JXOT9VDSC7i0s6LB/Hs1MA2tI7EeXPTLN0et
qODctqMRA5H27ihI1/hBqiIEXD+yJbJVugcBHrIqoh18Y5jTWMwjmGZdNoiS
qke5RIdb2XIw1piWM43pahAG715vkwW/cU0uhCfhwNqZm5oW7/hGPLGNyaYl
qNeJ2qB5SLMS0mune63BAioVpdr/tE19vaNryA1Kv6+hpCLAFjlsEqJ2RR2F
fKcFaIgYBNIChZKN9PyzkW9x4MwAoJVeVrSasyMqcnivLnIhDlj4tCJIF5SE
OItRWSU/fntO3RYdx88mG8fMc4PPNoyF/D30RZRFlz6WRvlagGSEcKeUOCC9
+2kgryiu8IG0UdTi/pAIMkXaYMUrtGmj5hTH261moUKlv4FzVBn3+y8UN7uK
up8L+WXI/qpLOyqvLtwMvKjxPH/rsEtB8HeKxlMr6cg8fM+/EgGybRtHNTlT
kp1qLJtXKUcU+flgRNOANIDchboWwjslFZUQkZOaEFHYsp3uC4cuqwnS0gD1
tZdayQ29R1TBCXzGN7ro4FVZs88fyy1/YLnN1tZRMsbkPRxPqhxCME4/zz35
WbL2kPX2NrZHUxwBlmbMfiFS5A5Gb9rs8Yi+D24Gl8GmzGlT/6B6plYZsvyk
s0rFpqTYGoPNUch635A6IQOI9xMbz5gW+yG7JL4+ahAOQJtQsKRP8KOolutl
daDtu4iSxIcb4gT3SJhI49h9MOiYZ8iEbIRCdu1DAagxHVYsI3POTon92RVo
Uz3vomP5xgt1atRvFyakjY49eUe1USOG+f0+1Rsei8lOllsZFRANrpHbcw8b
jfeWD4nQLZ2V87KEhpbIHulTiLI6wgvDpM15kGVAuhNu25yZCq6GKw+PEGb1
saXvgxDx+6GBPyTCC2jZkJTojibEuceYTugjT8Y1AbM0YdSQI4lMTEsmUpnS
u3HN6xTuPjPOWWsHxRRQQ9EPxM6I5Q+TgahpQj1+Cfg9B/L4Tlq1ugVhg8SY
XjByFpcAQEL/4xX0cmqxOyk+G60KtVK39zGNkO2N4Bzbxkcrs4BoA8aUDeP/
epuyl2ZpbuQJ2VlEuavmorX2d4VC5s6fCqPbpSxAH92CvVjgVLx2u8eshErX
VUW4iZTjRoi6DoIQHSiVShNtaPuMg69wMOhryPKV7rmER+NJegFX2h06NXBA
/uOSOjK+IDAtLd2BxAe8rYltITkRiNI0x5oRD5UjlR6fjGbbFSCy/aErLfOx
uxtxm0pv4tmyCXnnel39h8+LCH8drdrkwjt5wh2S4haRqMrHb9X6jOxS5548
pViEPPUltlKDZC2MNi9VOow8QwzWHD9GrZdjQvPqn7oJ8s457o4r5JgWpFRJ
uYRzNjyhWS/CCd3zYIpl00YXTenxsCkAvjsaRlGW0TKT/YcOrrDC1syXsODv
lY/IWTYRCl70R3haaiQuDobaEv3vxsYkJQFZnUl6S99BfO1CK4ZKDaqGt5Id
NYLZSSmFjeMs6yczkqpoFel742lvB8tNeedA6/WK7Tb5z11Xkd3LJnZ8jfFf
FTtb4jk4y8nvSRFK2NGAYyeVOAL0Mpym7BwEwFsVWebR2aZkYGDTrgEApWKV
1aoNb4HsaWDHtYkjI+otucj7y0EDp4CC7nzjv13BSnTEwN9sCzbdZegdVw1r
L/suSo0Gh6ZU68Ea1SJGXPVqvw0Ekb5b39aokVdS1pJPv5os2djxqrvIXHAC
OobgV2wd0DNdQ2qjDseHkWtRJHViTP2HpY9ndexl4r20LHquJnPjIpqBgyqi
2Mo9y1NjslDCNEtm/H0k4QIZk0/YsLWRYOCfQpcnLnOFyx8E9qUWRO1jTo3O
k9pUyl4SJPZWy5giO3sCVQqHLsIpFkJ45LBuZKqYhIS5FbmIbrqSINQwp/vU
eknLCNhBrEQtxdbTG8W55nQJPj9hiqXxb1bi5NVdoehLRwv2DhgxYzLuMhj5
5SBYay/YVecZQaM3qtQsrHYh2ZpARGNzz506bu9g+LT7fD40xPJrnvqykO9O
INATxWUxudkJyZI5UtDkm9b/t3hIeCZCcWjRGQt82bDEzEkgIox9ags4TlJe
7sW28KmG1gEEABwNWnntcmZUsHocH7ahR1jjuIFNTQj9miACSuf6/Eln7xIQ
5Jea4Yo0mYeUXTutvAhQDwT3mYjJGEGnCr2jFryu76SSSZ0bqXOszo2jcv2w
dGzuXYTiRxoVkghTDJPqwWKSS1mCyEtkVQe1eVwBDc2iGVLIyUm4LHHk34Ug
286W+cDe7Mh0t9uyicrNTBtKKVj1rTG/9BCHGsWjDO3LpKuqfpbtzdIDuDiE
Az4ZWn6FYyHoLq3DCinzSEjNsr4zGqOnHyzqSTMBjarnn0WP4FTeOv1MxjHp
3edcTaeMz7rIomD93Xt2oXLtxcV0XMNYazAQz4UKRNpLOrbAE0cwURR6mZvc
dK2ltmcRmuNisP9amRrrIgzuAmp0y+uIBFJ0Q+QfcyqZK4jXPlWtDcBPWtk4
4cB34nYrjfNPeSXMUL5SmgW+RJGQwX6FBHgrIMulehXzR41zqL9hpupwndZj
JWKNTCsujMuupR7MKhgARRA9eKY/pGPRGY16eyct1q4r/n3MKK2dl/znkqbZ
BoGxoQxMA93e3VCiTNXiJ3J5rKdrH3AUvyA7wkiWKdv7Z7YBDuLaEJl4Fn4B
Gnwiv/KMQFwMrsDdwQKmBYd+2qRH3gX2urbh+/++Dk6XFRrT9OPhNBQNfvWd
il9ZrBZtWYCxSuF/D+J2cMlMAuxuO5cNiEADSer+2zrlmEqmELXEiTNGeQLn
LMsZnwHTPumCxmx64pA8cJQE3LGMkS1wpGMtnSCY1WxXsQ2I9MTtPezULY4H
KiGtp+/puP0MnRsC6SxCisexu/N0lyEaAkfA1Y5bKf7fvjjqXyObaTjMRbFp
tlB7ZTuYYwj2US2ixoRmdXmrTtjx3YWYB+wmJgaeuwgYfxUSIjxcO4WdOyvN
AuDuzGhS+yuYMLjfLP06PEiQ5quQVYZVRQUj+1LK+h+WDcTBQTnEpWp2yc7R
9DMNgx1P5xxZetRZS7W4aCpxP/pmj+edFgebDCBs1pY/B5FigLwIqTjJCpRh
TfjlPDYOuKlTo0pVT5YP3vNm9Oe6w6pWMXerCR5KiJo9R1ipu7jLFc6D2oXg
Bfs4RB1AHSdkgbQ7Oo2y0r6j3Q4oAAlQzFudSLv+0jTFpG6OpURi4pewT5+s
gH8GUkyXyf5GdkMv9vyM55RYSDugX4iKpq8Drz0qTotW8JmIz7xNNSHCQ+en
W4vT431aThS9LMzZin1p+juDKljwvRv/YD8r6MA3mnBQxgPrGL9wB9ZdkE5c
TUYMHcLR3n8ZBXJCA3eQcBoOM5SbKC8+ll61T58bPBvCVJEKWjFXn6ISFSmN
qj9SeQ9PahxgatDvbSHZY5XYDpH4pkhE5U+uwahXP5vRNo1hW0cHz6VJszvN
4lRAW23ZmrAL+suIpjfPutJQHHG42tNaB5STqHAOX/wj4/jswG4egHKOQThx
6vTSacXQr6svdoVFZTYcVO4MBZSk2Raz8LIdkLIdvgJIFt7nznOhsHgvbGIE
8SGuR+7DjWXFVZxEU7wtaVKZHLUvucD7DWv4WV0ZgZLfzj0k52QUwWtB+Kq0
A44DsjeO6ctQc9DFQiqLORmNI1VrDnFyd3Oz78ITgHXHEslxZtLlJRp9Ol94
lt85dnwhPwwgVMfMpLPCcJ2TffWDxAeLkyw9iuzb9qBV52ok13mu36YWHQsh
0Df/XzTozbISJqE0qoDM0dve2sHsenEnjKEBSKG6lIF+/aT2Bfur3d1D9IuU
84XcUIYPWam1y3s4OCitEvYWtsd93KkPgFo+AuCPqGF7FTBwfOnHjJj2811B
ZkENKqzX8IVCGKYGyhWkCqKqBQd1FmNGo2zGH7XP9zgbszG0e7QaYApQFecF
y3+xDSEgNjkssMvOI6rXnSImGg0mthsquNh2Ceh4wjqYTZGxHCTKWjUOmnc7
85fK9hP3fGSS66OXjCA48QhTVL+Y4exky3oAxKFAbXmLrWUjsrTjeSnRX/M9
MgHt9cs0rYdIeBfWtzp6FlL67nFTKy8WDkFMjojzspzNAn4yONrH4HCe57Qu
zD8Bb/YHJXfCVz+INSSFcDh1gbRoukX1uFX7/viWtSEOvejR5C/TlYYsbuWV
dPGVwlDZuEK7OfRAnCsFrU67ld504CMYR8p0NJrgxbitOV+fhgSvCcgLLbmx
MSLti/NdijgPNWli1AxybAIIQdy/eZ68mwuimN1JrGQgvEGQhQAr/BhgVlLH
W0QvWxPyGTgeJ5kh+9uDUiwmj/ZAtWGdoSQ9i2BbppqbJv2Y9SI0HeQADGvM
2Wb+BGjCaNyO3vUSfM6uQGrRsfP4LT2cSfBXCLHqQDliu/FkiBMvHLRlVW74
jJLRWDpr7jY/JRhtGMyKaPX0cJfYzcXRc9nx8CnWJU2+hQB9SFrOQoJRqySa
ndMk8YSXnFje3I64/RjSJEWodNOKIA9QwjEbijSlQErSsDvFaqk49RRP4q8f
+EXz/N+NmSPLjwew6DVwmlmHmzoYwdDZO7wLBs5F5wQ4cms8cOUtD7I7k9wY
R4Eyn1qJDfvFFTA9I+ElWkWhsxHCczYOvJxw8rJGjTxlBN7AljvBn2PxOGZ4
hp9COJEEZHfhTn5Ci0zhBb4Qa5kPEbmAJwR5XBVKjGM0vMDD26bAKk+wo6es
wt9ej9YA6ZLD5xryNwfzvVOieM2FySZiLdkTra8B0dzqO33BDf2g3rniZXhl
Dp3MRYHW2GgxHXSE5uOd/HfBJdcQbSPIJL7OJZLiMRJo3yEUbgPQkd0qUq6j
aUrOTtgZ4Jkz7ZTRsN8GfFbN670o0eKxnsV+XcAF1Q7ycNisxQQBBxq+eUvI
X9WQnJuDtSHl+cANsDo8tGkQU4poIw68sq7/l2M6Uk65DiCIKPr7zSglM4yc
7swd3KnA1aT8EURi8Pwm/V6oGsG822CiyZhp+HtXy2XYleH76Am6xNJkdkHq
cowoJclWFBbizmFs99914Z0e3+5YCl1LIEMj/5dh2oj1ceZjmIg9lwEwJ3/Y
WMhU70IIOc5wqpVP5RgV8Xz67RFbb7flkWt7lAomvkldl+i5aZAY2XlwCT4G
mkG6RFta4uqp+Wpjoo+JnNpHle21foR6/y3kEjWNCEID1X4C9RzLtC1i1IQt
p3nZAYrN+mKctiRMuc4bidp+S+0IGHOLC30NNGQ1F3naODD1fj5PUsLR17XJ
2QZ3z5WfaesAF6JF9v41HQ5Nwo2xtKppJlh0DB9ehb/krRiRkl7IotwDqwKn
VZ2KTKzNbvZFzmo9O2pjlY/ba180hOsBOi2UgTOkM0Wi51qBB7Tf4PrKb8iT
CANm3VacQ3v89ArDa6Iscq8Ks7ndVbrcQfdRUYYM0bnJ/l6vq1cMfSIuxCi8
t5B/nOJr46RV96T5lRgQHSpd+DwkSMNuhHqR0s5GZ3JrG4uHMmFpYe4SI3/S
p5+3oI1leRnffgS62s6oGcs7Vemai5TMI8g+b4ojstKKJGHHTSgZ0ww8AfBy
rTxnb2Q42jvpy0l3cpTMhRXbWO9yW/LS1oQzU/1qWuBrhAgxaTGPu2vQq6UI
OFjnDh8p3LCcv4j8vOC15j9ZqfvAljmmAoaqZZfR4p9cUWSLOU4VdxhpKNOA
qVzrjPpuQT9Buq+/ievapa2c2UNfbgLHN1iR0YPLCq9I8KXeRXnKsjJB7QHi
ddEIJSfrvJuwpjhDao0vwenjXP/E4OUnHuZUx1UXiSogm/6Ig2kjUAwfg6A2
8KO8p/wkVzdI5g+7lQgZHlS1BiXI8W1ZGYs6kUkmBMkccAjvw7idBFRXp1Kt
KOcb+bTM/tzGN1GH7mOrL127jgTO8yvRvuGOaPfHpYGMmmYkMADgS6WQZlMx
Uj/J2asHANFqib7+4EcPYPuAcX7BTEJ0iWyu15PNVzhXC0giABn8fyJ72RUL
PMY2vcbemoOWzlLnjFHjfopImUQhv84DijNPGmI7GvGJeRAEf7gfGUHfb0Zt
wVFtdxorPtiajAmBr9C+ZW/iBx9SDTezYXqMkvwnozlnPwiMDHpnZXhlkMZ/
H2WSsPC7Qb4r8cNBwL/RhZ1GkEZM2ktVps4iACSVnNm8tf6toYNVyOLF36c2
NXMmetYbcKTtah/AWxjm9/NBRNq3wXkqy1h+JpdyjZtNPiXYjJa456CNN/xN
tc61bFjaFR/vUXvUvLINNMyCvaZw4PE1KEbLlvkroJODarXBzI7KBgADgr2f
8AlutcDmMcBpHOMEV17+TGry5aR6nOF3+6sI5TCTepzcgo++4RE2EhKil6em
zn12J4APSC/ac/8Zv1PafkXkMxidkop1I1j3R+XI8ynG2/Mzc1iigT8CRbf9
adtrmAbM+iQgluJh8pmsmNMiXfzPMD6cEhMccMwO0/R1B5zSdAiSsXoaT7xh
+gMFlUYNBe7It/RYM/RbGRbEDGIYsArL2lOqWIijgmeHM7dNmtxFCXN+hpFx
qC3NY2WGgsjNEK/FsUxV/kRoN5cGkEDEcZ+oSyE3mQOErDZ0cSxNtYYAEaJv
+YxezVpwc8lt4uluOPoL7EC8E3J1RJViASA2Bam6685UMpjGnVSJhKYaIS7S
4fswiE8prkkN3A00M/rvCHuKE3BHDP8Vpy2GOo+4qP4+ROpJcrXpposcEM47
MCg2YRKlZSGmz47glkRg7TNNBDmldM2XMY2VhM4Llo5NFityO5vGqqM8MJLC
6hwuOH1s8UoZ6kqueRcik9xxdeMxlyikoZzswSLfc3i8LSwPCNvPCowCc8ZG
tboXHyL/A1LhzUfz1RDmtQIRHESng9v/4C+Uc1AU0niAtqVjKbHamcRhKtND
MVIScKhhoaOD5gSkMSxGC+PRkJ1yyL2bpKTRRa+13satiop/Yk2J7ifqYT1o
8mNMOR40tpFHGX1SN9XkaRYOufDB4BjscUUDyGkWJeIeWxCXrdXZqyXJURpQ
SV6fUWEdFUSwxeddEOKg8CMws+4QGqUP8cawZi7F8bDbl3atk6mZQXV2JwfZ
7ccvlr1eqjy0pUnq/l1GrNwCs/hWn+0WQ9hqvPRT5bE6yvHQZC99ZdADx5QE
G0mU5ecwTXGd+G3AYOw4tr0sI75ZgDRw0Hz0llZVtwo7XJmkiCdgNuR01+aL
SzVpyMwxx/lwmoh00yK39nlTYj9ZxERd+LIDr/yPoGoZGf+j21yUkmOSOFce
G0wx5ESz9LGRTuNA7uUXWop4aZLV5h1yqT2nWXCqGSULCkQ0izUkbyef+27y
7YdFfaKFt83+0GYnK6RQEeufkGhYW9mutVnwiYUq4fCXfChcJG4n9elBLZfv
0DTPjhj9d7UsRxDKI6939/wdT1rTL8MRIittjEuQnK69odCyrHHRHKcALFhV
RzLs+4iSbQ1jhd076xqXwNS84zNlnIWqAAo/ad97Xee/64y9XTztLtvtJAk0
4Vq0qiskV02EavNDlPEFpcYMZYXU4rySlp8GRmqFCGZ24UgiHWRWhRhv5LjM
uD9pVZYNXkYljBtwSQAvHb+w4lghGpJi+i0TkHZdZMe0ZHt0W4uTFvw5u5Xw
8V/Sv80Lxvynhs7XB77lLiOvzbG58beNSV6MM7tfzeWShuDF4tWlFFDOQ6Og
1vbxpQLzP0KqBu891gWVDbAgF6vZT7Vq6TLVJZVDvahmKnvH5ZDynIZjq+QC
KY1VGq7KrnEyd+fYMjpa0U+qwB8Ap0UETXDQbvAY91OY4gIn7EXmsDe9dYrm
+/lQL0vJgDTsC6tdKd2FlLeH7W9m88WC3zEDtnsVsR722Kq45bg/tLI8hzyP
3A7dm8J43bxPjVULHjvrXxGJnSi/6Lu+m/G48ng5Kxqp6Whb9adde7OA6WRs
7QQRErfkMI1xrkJFxRu6JkyDM/g8vf6AJ7Nqd8o7oyvxLqCvwz7uQx0QLXv2
uOaX0wyL+0yIbc1TU9wNCx1dU3jBb8HuUyUGOh515G93juDenJor9lfovGlC
ZYM9zm2XmHYje0+b/zBnZ3leyIsi2VOVEXv7MnIi8kEwH8/+4Av0qcXuLLvQ
4yHDuK+kFr7W+6NEeq7LsnzlCT5UQ7V+1TgqT5jcH6Y0GX7K/3GaLv078XfY
cGCRyWFMWc06OEcrGkg9n/Fy4f4fafJ56qFsLxy22qFRlYX49iG89S3XAb/h
NAvuVdluDY/mld7q4Rn2eNKRXaj9CsmVoB/8fWKi88OlGK1i2iz5vcl9cLKd
BM34GC/iOt3bDQKEjUv0Ix5kOyu2q+7mA8v9CgrdrHZFEtd4aHvC6601WwSZ
yQXvqQIKTA6U1BCGbOj9KRXYxcVua6Bl273oWK2Q60Q5hbFW5dqnLXNtfL3W
HiupbpnjcxKpngAFBNoKKMwRFSwKg1X3IydXf086yFicZN22E0lQwcHiTR8v
isU31lun4U1hYv2G1/vXYnptMeyVJmtcssC1Oosio57GVe5ab3bkgbVvrHnC
pI0sB3JGymiBuLPCd/I2v0ivO8M48cbXMKh57Jw8o2blhK5wiRvSwyEGPr+d
r5RhZpO4fIr1Nzk3VhMJraFyCtRYwYOLdu4dJaQZhooddf6Q++75zaBKajb+
NikmyFcatzsnFq+aeMVKWPJ1qqByhuR0Bkk+sG59QWmKpCDsUyE2/xPAXsnH
T14Se5htkt010S80RDNfrVcIu6Rb9HMKjWL1x9O767/hmVaqrNWFtEP0yF3I
qtMiGw7o9vsYVgvw42zIFL85nnBXINlkUmHT2rxY4MP+hlpzStsQio3CJBIa
c6k7pdCjq0nR5RX61bfpA6NExg0RQj426Fl5nCDYNO7E140WAI5zBMfKBWyJ
BZYyADx93G6POyEMpmEwdGw0glVqa2KPWJUf1mjYNbaYnS41newDKGyNsQcJ
q4oJtgnvx2RngzdPAoC2wN8nmLEM6fZyPic+kRNrBqtsUWmJPGqaEt4WGfur
WOQ6VAkJoN+zaPYJ8IuI2O4/dR981kW/wt2G7jijFbkObtHDVYo1jXSeO3up
ZGrM4hqepK/s5+OkeCqF9TkgaTtVJ9ZbKGXkdX8IGyrBNGNPIY46pBrMhMBP
zYKd9hG0VpJ3v4R4jOCgIsPrM3KaJlJzVtKSaIuEmHJDbJp55r5rDjuhwpjx
ro0t+FV7Cpxp9g1nPcH7CDtejCphPDfUkT5EvUoUeMnNoV+k9ew0ATEq76hs
CJe0tgsVv4vYncgdXgqOp403O+YCiB8Zm0CueLkwuzRUMqTmhFqn/eJafSRc
vBoIOlAHY9VJb1Z+q/YvAksj1ZJlVPau6Pzl5AdDMA7/1YZQg8aGl57OY3lC
TYwj9/6ru00gmCMIMbtEshCaS3lSzhIVOt71Z4UC2/OMafiOrMA6HlccmPQ/
72wtxnhA6Z9ckUEWu8YvcLIonZHbJLM8IRrgghm5Uvl1ompnogfUozYdQKgB
PjhZufENZMkPkrU/qENEFajqyE8Rj3O9bWi+F90Tq+xI41+o+bKgTDZMi4ke
qd8fhRhfHUIVbsgsa5+mYIxceMmzMvTDTPpagMInLY31G7poklcZ4ik2Zsxu
jVG+gxeKpUX0jmI08/4ss+ipb73Yp1EvVIHlaamUe7uaFRJY9NNDJET1AlK1
fVpPcyDP2ffsTaNrj1qGp3/87OCelHjomSU1VX9bDEmhlZXSUEGpBePBJTXE
wNi74tw5Bs6A/jmDDLRj1gboH9m23VKYrPhj0OB6WCFeUISM3zJsgqp+RlB5
nUCNlEd5xo4AIt5EROGWEqfXnifC1xDU2XKswt3b6R9h+ItJ/Y8DHP30t5rc
41eEGPUlV9vE9VrQiNw2aQ7umGXDcCX+wJXaOQjVl7MFRKjt0eYm2hZHaRgz
dy5x9krLId2wXhsNRDb4NIQ78hxggmEAenQ45Kp6okFOAV0xciMlHPKOu3Zo
yNkLjJO8ZkngiMTQKYP29JIU46qvlZFf6/SpdpxhBvE0noF2phkigYnZTDDu
v7sYVqIa1bWCT0jL+2zV+tml6y8Ev8ZYNbJgEotE6/TA3EPFXldZMLUe0AA5
9Kfdh0Dr3a0rnAXvJ6OD3oj8qGdZbVvyFN3KiEUcTNU0qE4uyKrBFIbLRB8j
wYOcSufo5Yn/BtsvmTlOHm4ylAT/8RnZgbEqFTfZP5VUAnNRmqhkJ1vo8FrV
/YymBbtKaVgvbaos+9L6TKCz3/Je2lmsEg7A8leM+IVAt3B9yhjD2r5twZvT
RjlQM0vwY/AtnfpDD2AmvubwsQBnPAUk1oklcWq4175n8Vl1fGSLQls8iQtC
0xEHCAD0lRQXLCzBkH7XEM5HPLGyf9/ynDPTDDi6bFTefRgtV7ONK3PSNnER
vShGDXzLLGXXdoFdxJDGC1aw3x6srFsR2GJ1Ng1i+tbq+Hg4FPltbTsIDaSM
4S3kOL2clbnSYHlwo+XWICwIBbKxQ2jj26C4EoPSHmgzX+UJxxSyUTWSASwE
PbocyUetSGJXU9fKHJixQXW6+/1Jp2LvaOoQ/2TYdJg16H3sSNybDETWRXoW
z2Y+4KH7+LhMrSK5O0RStZY8bIuhce7QCLR6fELIw8f8aZVmp5DROCJQnE3I
Ww0XCFxvFr+So7J2KPaawEjsCFb/9XWo53UNryIbsh/s3G8hLol0c63VBnBK
P7yD2FyF0mgcriwbuaoAdv5PMAWDnC4Ui6WnHmqVvE4ymrXlwEC2oa7lX0c4
FNhCzdvGCj7xDeCnr1zXSIjJ0iI98Wk0uNfiUUBCqRWE+ukMH2zY8dU7cpiC
ltmz34V3Zd1U3cuk3rW6S5ESsPdraRVmRMi0KbTtMD1hhuzlFtKHGQqxSVId
vND0nYfMgq+tq/OKr1QWIthR2Cb0ULrLd8cl+a1wupuZ+dPO0lH2DCw+8fTo
TiIPlsVTh5hO4kbxCrLufYqpZxquX/1tsGH18LibSYklz/tiSDTF1Z/HJ1Hd
+hvy7yD3yqo+JEbvXZbafRC7bI5Ct4YCZTPkpoVi7gMY4KKbUK0KwKYxaprs
gju6U1g72GVO8892kZZJpOUlWI0QDtF3F2TjjshTLTPFw8JXrh1fVBZkPfrJ
gB1yse4NpoGAbgiMF9JYvcW7pQ6ojgkYjg7VICQzaVIvik1Q0N63M0uJM29f
IBo1QGILgZ6cofgbgKzmMs1yOzXwEK4BD3tWGFwSkNAhhLVOskwnU6WyrFou
j3Ggm6GlR1iRPKMbJQNsSVxoeN4xcrAbhOyWeYBGsT/6Vbrv8AplLsoouZwM
mK+Cm7PqyXFCvOfElPG4ABwqPeU9aPphEZHr+zcOufxHHwTMT97Xx222dwtS
IN4Gj5QVk9tPCoMcC+VL4K46KZANMYbl7ZWKncEjnxfX9Z6qrI+TrQZgoFg6
Gd6NRXmCwGct0oMjK23CvJI5BjHXK4adMHvDxlbOK4ML+8EE3bxA5lx/08NG
u5RW+vwRRcLaPhz6TYDFuRjr4LUx/RKZY3DDnkX8lhxQ1akVI56hbB4c9s6u
h3ZaqQrLOyuKb+ILidbAVJBuSRsPmXRAum719SspLKMrw/XKBFC2vy0isdXR
JaPMd2d9fUFCqNs1mlF+of0CKzZ4tJcxPD52xeoPDsmWg8fyCGKnGKJFhQGR
kkqSpZgS2AHKwTd3sWjufgs9ZzbeVzVGystSwKVD5b0xB8j03T/8s7b4yWW6
qVt35gOGAu6eZ3h9DYD1JWoTHhpnRRLVOzUDyfnRd9YL7N0I8uMSFzDB8SxK
zo7SxFZNvkI7ARpM6U+Ndr57/XmYnId+pjo4MY1d9BXBZC2rU1OsjbB+z23o
WaL/GleifAdOB+6wkKFl7DHbjzAJvyr5sGWEhzWvu3zCK84kVAowBb2Fmi93
QIf1dvHbgMxngntZ2sbvcAE4vWxjhDxtfc9gsBDcHiBIcxUBtBt+PyMDyocj
JFqAjUAr2DDaw+LyvX7PaNl1ur1dpPJWduUVhPSe0Owjqkz+0YIPtjbpgp2V
yvZey7Wqjxxcw5Pi8rNHslEUmhkNwedkkwUUbhRHwmZZwp+muoJUdWeErpdE
xmrCC2m9itYHVjeSZVbyeQr6HAzrVSbcmOo+UEw6aMov0eSveIx81zsN0PRU
n1730GaqPzGN4LgxwjgGG4fdXIRf9mTB8Qol9/m/BrCCwVQr7mxb6SeSv2ta
3x0UMTNYcDClhlQtFBuEriGrR9jpQRgNkcgqVgdWeRmcLGlVhkeY7k+aEvIp
d14lgj9oVF9kcxp3RHwbpWEJrm+47VXo0oyTf/dD6XbT6uD1jhj2r25HjfNG
/0JnYPWECu65vDBCFEbLZi0HXL9XUaGq+KF125X0HGkbqF9+2APsQ+4B3dOR
HF7Y9qkxJPsOkcaPK5u+Bs7xP0x3VIpTN3r7Le/GYR/tpK+mX2P6Nc9ZXYmt
cDsMqy4QLQxBL+9joMrQSDlPehh0KRRfZqKRTmPAJF04bjVEQXCNmcisL4jt
GNP6SS8LwZ8psZRu3NqXopG7bEOwgnRssSw9r8ITYTuncniAKz8MIJKYWm0g
BOXt6Xvg3jjg+pxvro83x+WJarsJpgHuKqKczP/CmvO3p4G2V5m7biO/hCGY
Topsv6Z/9SrpJ3Dk2bEygbn814PVj+5JmqBxmWFbELh+l9kJ5V7HKEBjShDZ
Nu3On7nLuYAUeb4eAV3HPkoF1fE6fBei1F+hIzoxViOhz1siPS7Nb1pt6d7k
FozuWJuj7KYDqEvNaeabvV21ZOmBeLh9pBm4N854wuYDhKX5NcNF42MCEsLz
H27YY2Dd/NwTuFaYt1+J4olIIEPb73Q/9s9z2JpixEyhL66JI/1g3lQifkF1
+tzpzCcaZGUdfQbPsUd77T5PMjpruM293qHkHuB0AMWUyaAxaZVAKE4sC3oa
C/GobRMbDt/XeB3K+wPjTXHm7vDYd7nRhLUtawUaYOs42D9jDCIhb/pmk5su
rm6kYUYU/PhFIs0rS8xIlIwBRgGu2AtNVLoPKuICM6lr1192d331kWTLkbcM
tYaGDV/DCAcj6yxIfAhiJS+QAWnTsQp3mEE2koYmW3EYDELTtzPQdt5NjN51
3gb/Tazxqvd8G0Gh41IvDrQACS9ImdPWkTvkwp6mBwURq3B4DNKvj8Z/cI9p
vNfkHODithGYSPGbDZCsVt+J00dCEQJIEfjJfT/Pp4uULMCShndasvB7oMy9
0jjLu4CQrRndH8NDqBXQuWjKsiyrd3FcWsluZ7/OynK3OkxecyyDgG+/updU
LOKs2dmPV76LgVZiClc49lewLLheTGcQAiifc3e33Rf+qSVuBdDpURQgOcw1
ob6TaBmQJpY+NZcQ+NGX/GcqfIc3pEFKxwgQ5mU4q3GpIXYcSuAPYkZDXVJj
gNn8TutZC3WsI11eGo0BdkbL6TOHCOg+ZF0NxnLcbSYmJmkapYItKNj0/fId
fRHiAxATdE3sRJkoshziY6nNXl+Fd645bLNYXAtWSHLTxKCrvSLytbpXHQYj
l4kHmlg4y2HwBEk/dwF8hhwS8g6rE0YzFnwG/THpIWtoQq+bJVqRNNzUCoOB
1/+KE4f9IT+0GTyv0wC2ZqKtLZ9NxMdZkJ+rLD1Q9Q+XQz8S6y0zSDaWgtZc
B+cP8D1TysePPgar6lMF2lT7KqMpC3XC69KDjJAKJNkZA1TKgZBV/NGJTGCQ
SA9az6hBSfs5+UcmY7tL9Ij4kMBQryZ1nx0JP7WVOc+IY3QSoQxN1mO7/QBg
F/9UjsFjKxbFq9YTFtmI2LAH/kODP7AQ2ew863mGvhWqhz+liKW3w87bz4wr
DI7fWaRu2ptYROFRxzt9xqUlDnPFtZRdnDu2CDd14uz9ltPo75bOyTSdJLtj
x+LuyiwW7gK/QD1RzYElS71RFRlogkTzkiZDlyYtbulRyJGNKB0bVhIhySbN
To6OCtX3qLSTo7QqWvfSRl06HF6iKdnumyiC7tdXOPOE4ZnyQ31O52AuJEJ5
84prp9gY5vBfDjqqyt2O7WOs9T/WCHD4Agyn8aSBUZ8Uwi+j4iGtkJPEt1ZA
kb5yhAHqOM7sTHO5uebvzHVj641WUCEUJXGK7BeJB3IUDwtaom4PqBUmGNkM
L5ygBC2V/hb/dsLJ1K8ztf+ODvV7oBUuRpKY7Yg3LvuzKbPqRU4MUUJC9dUo
jid61okJEI2tql+jSPg8GnkPuNbPnKny82OpmZdE0sfAr9DsWp7AAU4T0bfl
r4JhNV+J+7d11genN5A68H/iWt7ndk0IfSiD/rCUiiebo3Ne6wL3SsOxVKEq
yh7tZL58jt3IZAWBQ47C9FYFTIUP/xWL6cjPjqO9TOTGjIzC9PrIbOf6l7KT
M8/fYLd1tE7NsrPRNf34W/oAWgF8UhaP22N7/EZmziCSeCobQiwNDKT1q6an
nb99fX9DZpNI8S+W9cn6shVCIkfJukE/7ac3B6gtnjr/Ru2OLa7/cY8B34C0
ZAfXeKUUQIIVtq3vxo+HS+bkBCT+wIFF+htIqG26JGFRIu/waeSBbbbJJPok
knTWxN/d73U9450avpi2tanX4doM2LIHB7Yw6ac/C1SwCiHmS3WHL6wF0+Tx
bJTVN5YCU6FU0Js3Y24U2RJgCoa+bOSHbNM6ApHBsvO2dlyC+gPmXK9H3uUz
Ric+caL3GyhMztsLoKIyZAkP2ovJmzRV6OdA3Yivv4Z+GgDdAmi5zdLriLo9
FQam9DCn50plSZbRCHVIYQRrspNLfQLGdo7aqpClp4qM4jDo0AhDLSk0LNwP
Tu6xfU3elx+m4AhfEBB4jBit9ASK6jMoanKMwUxfsGJjvHhd34g+tcEagPo9
gsZFrlfNOqvjkCwDCUJUpZal93h3HKLBOM6BuSlZHMHvIgFvr5P8t/JCuz8T
Z32grC2mnJNEksFqhZ1MfXPwPcu5lonC/KRXtsYpM/TvOkz54mWfDDdTFySE
afM4lWR6DDjwQGKs9GCbkzwN+69wdI3N/y3WZ6PilGOCNthT9G3JMoiiNPpj
PaEmrpHF8lJm7MT63ViFnIKFRFmiCjJFoL2HWmVqmpswhVAorunbkvs674zb
SUQkpOc658dd9HqRZOMWMSzpOl5Tat5TvAqlWcPJf6d1oqfJ9StfkGxpCMnN
FybOz91orz7WXBf94FAAcmB2vY+vtAB+yczpSb1ey0oTbkA4f88SEkSbxtu9
wBvoyDnf4vGnOiR+kOu2GAayTXWZbAJ3nX1x0QYYmTa1aJBZEfyFJxqhI2aB
UH7Q9dqk3uKVVVh0UYycBrsOZyfWTKvNefvN9chd2hY/V7kSjKUel3oSw0BL
jI/kTzUkDnYaduWwcX8w0RsLHoryOS+F3a3/oMXWHPDN7SirklbhVBv51O8g
INJYph60dwozU0bl32KbAGwyjfGLZAZXLrpeu1ISTtYIOJzdSNx/PqOma6Hv
I95oFnL6cR5cveognCdRsAIUTxmPkfL7VxC/pL2lK6AeUXSRykCZBhCLk+1C
yDe+HUoY2/deCKHBKra4w+b75jmBs0Zwbr7sRBj4QqPaYmjKeMTKDIt/azug
RXcbF0OGeufVZ9FjyVm6irms2xH5QQ7KPCejqw11L00hV0hJnLrYExrxj9Aj
uRs5OCF8N2JEyyDkm7LZ3bcxEbl1aZXug58p9XjocbsZb6/SsJIl6gFD4QgA
OJWMaVfF53MDIJ+VJrzfQrvAyh8fwrY8/JzjHMafS9cLQ8VaWKp6HDc7ZuJp
0a75Tj1e0QXy7drE2KKKSGWV9OJZzE3VPf+G4lATIABeMolpANkGPDPkrsag
Llt5+hkmR58j/Z/nhz7ZSoXab1ipg9Htxoe2tJW/Gp2u8a4Zafy0nlodH1ca
m2wM5zCt4A08MB7eq/dcn/i2JQziNNCI18Hyaeu3yUEds1eTxyFXI6b7MHVJ
/HZ8JXcXoHocOlCkTBWDV0g8qPgo8+37QmgVBpMfNEJqiVL6kZDfvGGrodyq
39+d8ibNmA8D0CmkNeFrjr8LAiL41Xq61A44+vaxUdzVTe4prKpBC+2vcsfJ
kw+PyAc8jFKJqyGYWBybYSzRIJMs8eT3A83j8yIC97CHb+O1JY1k4gaDiWUf
ILIuyK8WrhWXUR/84iI3zF6Pqfdud/h27fkWWcOfPRi0o+WO4SL/a0xqyBOz
t7UK7Y03xO6ItjEAPe0sZV36AAJ236p+r9z8BibKgb4vEQqcjLwuex71lV6f
vzRooigpBc98dVRyoqx+sbTBwZma2bHDv4n/C9AmGXUCovh+M+JbuUhuOnkY
DBLYL9sCl3flE1Rxc+jV7ipY8AsjZGjz/yTv8BVX6+gXZKTrw+GQNxJPJyYg
jJI7UjbFSZwjTrr+f0WhgEn/HQK2W6GSR23ZQmQlhmNc4lDv54q7E8OBYFN8
h/e4RDXtxw3y3/R2LxV69rLyFu9HEuA3285mJHxPdwKHLqIrGoxaEFw3oELW
C1EsBYsDKty0Jwa1yX/r6+36BxelH0ep4P/bte34kjQTHoMuzVLXdACoC8DD
XniKkBAOU1Gjs59s6yCT2Zl6+bMxmoUvMm8Gj+QXOOkniWGceezbjbsbuLTM
gYvvZLj2J2qSEWAfYOVDpDQEMBQWhvWPF2jEuz81xCcDC1o9ndhJ46u620pC
9hlhPKYoS00PsMP9b89RcHNS1STbzECzSHBCbyjxUDMK+Xtq52S7nW/N19Ge
suTei8vThj4ocKuPBNzrZRTHm46OCiLqAiBlR2WQ2YWyCMJu1Bplzk5U1uyD
FDQKhquf0zzv/wYeG9l+XUOU12DO8VQ+YMmcC4Xr54W9bFRMLw1xFDn1M0K4
QIiHJk9yL+oaDddR2kwd/19i1wyUgJoAPvoGc94Mb/uO0MjDEcgrHi75begv
2v9CixauSaP3slpg2Puz5dG0XvTpxBtRIfV8lNp4Limo1UjG8WVmJfpO08zJ
k9E4ynDc8ET1RfzXG+8610DexNPMzj0OqU+NvjMZ4MW0I1kR8Ri5wr2zNs2o
heUnGgS7ntpCQIPVx6n/yy8xEkP1tnVbG1j2vthqULf/t83z9yaTGhWcroZC
FTK6Xwbl5oWWBKZqttrMN7oB6j4LYYsbGFVDUtwzElVd9yhmkl72y+Ui9QbM
2G7k4jLr+bqkL/zlBAwlOntGrFqrqo3TEXSdxDQEw2jZlNQognsEa9U8M9yC
/PYvY33bmY6Rrlx7FLqR1ChHkhWp7DrVbG4bzH/ln2yIIGSPRrWHvnNoa/5n
xYt3QzO2Zzu3pBqWxG+NZ0l8ZP7GKPsKXIvNbZq1D6byLQ2L92WYiAZl5GC6
Yfp1jOWeWbG6ahvxygT13//y/1f06XZZ8Pl3TjG+Nt2QnBCVY66oFUBxsvp2
8fPjuooN1cT7wMa7phtO8rfhX0g3XxQCZh5bT5Sozlw5mKtCLJjAJeAQnx9N
M5UwBiRFQDJNpMmVWupRDi2CBReljURlP60N6XJ+lWssOzkMMmL+MSaHkwhQ
aorOWyjeDuO+40MFrYsVBScnJa78+vW8txTnhP2ov9liYAeHzYzGaZSu01of
CX7CKlqYFwr86Kt79Y/utStPM8uMBnzsiDc+b798BgTiNJMtuzqsmvzubgiP
pgNaQJgi1H/PMO6P+4NQu6RFwfsLV0CH5kPhyCJzT3PmpYJSDe9ttOmVNnfT
gpOoQBMBdwNaDTrB7FaK1Glbs/n9khm2wnUoLT6r9dMUp6PkORdCAEKz2gfZ
wpUXVC3hqhyZPCIlA7n0YaN+n6NYXgpwTHDH4euke0dXfLramwh1ZjTbuRxs
EV1/ztdRNOFl3vIZ7LRQUhnzla67DjJJTcEjUaJAtXfpwl5dg05OSfbnlHf6
Ap0K2vilR6Mbs9DiRP8SWbl/n8Y1/iiXDtP/3ima86xZk8/oghfr792AVgbZ
ecjSCyfOhrydf9Tf2Tvu8PfowU5z3nWZi1EaxDI85zSi8UTBqEy7jdXBCERs
FLtv8wMUmM1qlI9O/zmFmfgtVK4ofsJ8LeaGoNiN3uPaC1MERh5P60WKDIAD
ZnesBsuUdbRoAsGnXd2Yk/sofYthXQbDsuCMHJ6HRjzw5kgxTZvH8uOkHAdM
KUAZfOj54gkxrjr+qAID5iU+nONRIzyOUB64cQIWqDCHQHe5OJIg5VK2N9/G
Sg0MOq7PlJsIAdpYQg79xfUkZ27l3ncO9AupvUjNvgSyWcCy5zrvrjCGZ5Xb
YJlMi7XmQ84kk8098CnD6siZwmrUs1rynRqe/Ntoc38KAORRPSP/7F8Os9uw
VdG45yx7F6JTPABbGDHzJs0Fvi2PC7BXNLY6+UbbsMcV75QNlKqmiIP6bJly
TfVqgVgEEtWkcPRIfEfi/HevPBa5q3dlBTLFn83jrxNyVKVMCUkHhN/2+15k
9eefmrnf/PLuDSsQFtrivitu/GRuv3asnzfupFEGb5U99A0BMzGYJtcQfXoF
KTjSopGvQ8PVpRW4rzdK003FIbUSDKjULUuKYKsB5+If9Fzd2ceTWK/ZYvEa
uBig54N0o9KaRgPaeVOaK7nQcp0BKR6wrByIhKcYANBxlj+pLlqLN5MUi3AZ
YWZ2VFj36CMCMnJXzj0kj2XLDFK+ZBI9qEI9JY54Mmini13/3Uo0EbocDBAj
hRbxFxdI0lvLDOsIyv+tlThe+HcaMmEdYI9PGXW8euIdOxSOY0QxUIRoZrgf
/gouiEC+nMbDoDSF8lCfYsjyyBd25tQTNJNdmjiGP4ygM6D/IRDfx0aeNqYf
AsXY4PQ67cDS5Mp1lvp3k/I1uOvMQ4tdTxL2ylQnT9myc8bgPyIwK2dZ0xMo
DFV+czRwT+yvSILZszJUEMD/oLdPnZQnqUz8QLi9WJ+oBA85HZWZbM6nYhXr
LXnHskv9NjB4xTr8HBdIyOa7Ao3i7/hGRlmFWxuDHoFRGffPnXFwKcapH2xw
lrduoPq7cCJDnjfbHvSo8EQpDO8bKBLhQdM3DwDI76HFXVn52GeCKngvuMHO
NIXd7rk3o+lYM3Y/T2euyKXEDeEF7krj2rY8SGEe8kskikRi9ZxnLpFeod3O
VAYR251zHcX8jATLN9cPU/c+ZWPpkCfAixH6/Jlh6Zk7eKKevFFCzEBF3mRF
rThw/eJFD+KERVvPreiuhLDlYnQ0DpqMnGXNA5NZHUpAq7+UvM/Mx2F+YeQU
uVTXPSJt3ANCcwBeg9oV67+bESn+hpwFO0Xtwq7GxTidhy4Rr8OviR5yyszz
HAKD0wgIhyVZ4ObxBsmvdDSl7RqbedR8C+xCvLVk7Jfub2F2HXb5A46m/+L5
nFv7Zv1o/e+ULsJn6VSnafow10wwLANd24NeZ5GbK/NUgcq4MUmRc8/7z6eo
CdXO4QWru7f5mkTS6mok67W7mV46hUf3XdD5CIUNMTG+C9vbRIRTPTd1oSZu
f/9xtRKdDxmeCao+7nEtmOXLyKwF+u8ce15AU89LfaGoJFiMkkMewRGcyzLZ
B5UVR84nH/5WKam4K+sXaW6MLZ7yShA7EFxYSMpNr0Wq8vdMV8Dymf8ENQyg
fQvFJwoDQl+Vc0qplPLJFHjaax1cPTsPDFQneQgG65gJKzjuQ588em8JZtCR
dnpZjSDLVyJSlxVTp2vtU2KDTdbrK0hjXbTaEYCHSXP33ZTyidJf+FZ2Ml+o
SCKQM7TCLreyPznLrJ7bQb96iucib8BVBWnVPRL465S8qL8U8tuDqUj8BT+R
vYVmqw11OjQHhyCq0F7Cujb8Sqnb24mV5WUCh8xIlRwUEG44gYcSAsg7knaS
kSjG0hHIoAqpE9v2eQiwXHoLKFJNPhoLZvGRG80nzipEfw6+Wy9O6c4yjlSr
El0exsW7DEgvuKtsMrCcv5KttNJDFhSPHy+orAL3PPhPNmx1f5tuhiFx9gxP
feTXgDyHnSxzQ7c/HN6OLF+YXhNVJbD8KQY+cLIjdp+ENUHn66dI9JzlruS2
IYWyNN5VRUIiYAhjqNHaHcDH8nfDYYtQaw5xN9Fp26cOFX43EDF+ET0VLZp6
axmMIBgzy9mTfELbfSA6H2kzPaF1EpiCnPCw6jLbFLCEPUGuVWsDhhw1Pddt
4jnE8crH64Jy7Rfhqo+SUm1i2TVzrTkDMn8j9sH7octUjWLW8Gt5qosY6l1w
LN7mndo6TT1YEEEGLrcwanzKit7wjLtpDn2MCJzy9VR9FPMv97qWYy0XbpEJ
WGPkD8M4deGJOwOogbzgYQ2QeR+4ewEBQM2gZ1xejlYVI3Gcm+484Q7lD+z0
1DEeyPNQrhB4TRZ8nlFdHaptftcCVPoIuZYB3Copu89eeQpa2ectj49RaeCr
rTKcG2SVqaowq6b8waVO/Yv4ZLQlsDV0dr3n+uT2Ugjc/aZ/aaSjNE452y1q
WqdiglTXk54TttLbXWxTxJr7VX/AzW8JkQEKhkQV8ZjBF9rVK1XqfW5RzEn9
zZeRijOnwyOsUrn+kJk0fIq6xHhn+/GL9F2zhu0wvum5J62ob8tm51nA9CMO
iQlEU9M9XxYgAuo9K5iismMvW8X7IxlKb40iFYULdlPXDgfqz1MnVjTBgf7g
lF6hBqXvFk8HhusHZIFG7TaATYxg/i3UmTOSlCNo7f2IAGf1d5StPyF5s3ld
cDtk84ov2xEIaQ6e97JcQ1UGNXW2FNUwm3RgMhvAEnYP3ZcvolDJtoCSMqCJ
m7D6zvVkJ/90xoUB/LfRGZt4uq4ejLJU5mJ9Bf3ozvWQ5MvsM2KzCdMCgaPf
lLRVkv94dfYbLoMPWQo/5fzc+3B3X0twzu1UeJzSJUGznuSgChTRdPRVRYYQ
SMZSf44SIeahA9HHNlKe5kiAGf+Kr5G5yeq49ItpUiYUZxNBXb9rOH2HLysy
BGor9AvjD0q0ObSuFCvTdR5zqyqMQGnkt9AUk3wJioUeETWKMHl2nlT8Gp5X
q8sCunMtFyyUkte6W87XbHIfv5lCGnKKtb7uTxwHgGkCA4skOJUdvquaNriO
YWI0/u8CcwkRnq9TVK95wHFjQ0McPPNQtchSgR8MHpeAxiCWLkX45uJIFOhG
j6xLkWNd+T0LP+k+ftdiDuch8fRV+RCjFw9ZTelshQM7xMtFWaA4qhbRXOwq
K5V50bK/22JZv0mcK/8mlC4NfQgIkltlqKXu4bgx92cprJIvo8xF2G5J0+EZ
ru+QqZxyMPDK3aVy5TasP6zMj8NKxDqaVS8puQqdDmYvapjNp5Dgg1W96dD8
NNSq4KObZgRzk8kRCmkak1xjshl0T9j7VJSYr/HdpmFjss6e6M76Cic5s/HM
sj1FoDWRZlm95lszHDiXN1dvfh6zYoMrL2K+lIpnz4vn6FshZoQDtaAiuVl8
+BPW+Z+RZjK59A9xH93IGo4DQymJ3pQYGUHYCnxhZLNKREWgqrP4m6Qs05co
QBzdo90wXWrwzW1fUDHClTMMYhLepREe3I/nSMjKcBZmnoH5NR77I2mop9MR
/JliqmGBnyW46nX7/IJGu8AjUK+NxFHapZSwfwN4ZXo5jjI9b721kJISzNoQ
T4HEYqTV2BA2NlSNZjiiLBFnqxhPPghUxt1vi2DFR07EPwxn0kVVUIMFxtKi
a/UX1wndjkDHic1ASNN/AQLk1HZC/DiNgkL1cTYHz9yAXSdWYdx1VQbAa+VY
49wg+ORAWYeoLoroes9VvRI5OshbSMuyESfvFYwpUL5oAx/chP6E3MKqgD/o
a9WsX8zk2CVO+5ORsbDQC/vNPpbrcFxdQap68SlOt/1od0zorVgk8QielF/b
PbYFieMEp3RE+90gHCFQDMgEG5du7z0dyetkazkObrBXU61E929gKkmqibP7
+uL1/JFgj8sKrLTykDu22soVdElTWdVYJlvAb+9/mbWzBN7dtmQlpuQ1ivoT
K9MAmywN3GCxznGDqnTcHxzam37nkbrcSnvKywLuWB7P2lqc3ihE79sX8K19
U5QTaydYfO7l4yAjN4S5KwXweUUgeweQdqIqwmOKB6kRROcvLLh+Ttv9aOUA
k0MBV5jqSY2+KHHwxM+qCB0l/BMDS1uHvqu0Mw6BQ13PVhuaDunMndncZkrA
skzflGg/NocZhbPnUWawbeeXvve7Iru3KpYR7M0HHiZCxs4IUEyWoi0O2sMO
ls8Pq3bdFf1SvwmjCFfIYvFK23MRF28tEvrZIRbmtw8f2vDcoR73U7d5Xzay
LOa5oHSwJ3hU52dlMlQE2BF5ZpLHe+gj09LjfrjMOJeKzCO2Rr8IEYnLXS63
T1ATuOgCnXz3ik3609r0XPg7VW9pXshQITA1NATMJXK6IiEuPnJstLVhr5g+
BKa71hiqNoXylxyVdLSLBk5rot85ldNQlUIphibMC7jrG0z5UW9nI5NX8cwm
AbnbG7mdFySWsOmsm35v8cygq7dyYUcUe2G1NJ8OPloUVlCxZjfDKRyN2wfO
vpWyyODYlYdj03YugHY94nsPX16alVaU+MpYT43FIrm6iVVQXVbdkyKVSPEq
hk1rtVPnJ76SdVUKDJVxO5bviPB2qaDOOvwZwGY4C1vJHlzkPv90oRildnrJ
+4qCNoUtqmO2m6Zs2iw8VIKHU9EHmUkwcpWRTRSSLmfzvj7dcc7TW7EjuZLT
BwH+2S4twYV9Oc9nj0jUa0+CmrlM8/rfc3dZvxShu1IJ/pCWAev9g0UYtIkR
/nEXUgnyKoEPzMPGHzkPwDwzr7FMeRAcLVCgtyQxibFKYW3IhCH2vQUBZBxe
0hPbwiLzcEZq0gGtFZ2Mv8cqcZ5zR5H8OaTRRN5C7AbXl06IGhuLiyyl+imq
T7TQEKGhfdYYgtrK5Axm6RUGz2AFx6xEV7HXJao21nH0ZQV2Hr6pM9P4eFnh
rvcyeSKrRW/8LFBq642dwQFLoXA65WxmhtFY3pW7AOgbtZdoSON1MdVfI6j2
/pxjl+5RDDrG/fB0bLv9FGVO5ZTHL6oZc37UdN1p+b8Wm8zkAY/D9vCaquxE
t1f2SgmhPnrgnpMsPjWlAlAmRadVyWDDN3EVWpWrnGVpD/3NUVsuKP512jhu
kEvB49LOXMrkmTZAzC+Wv/RVI9hlKDvEfMNy912jNwrsv6hevZSOMcyCuva1
dI+MZIhiiY+4UddAeY2zRSs/VSQtgsWa1XWkiT8tXuwOSctmHuAVpoWYBZTX
JXlyVtG6YNVEa285mhFfHaG+RcVvZKsTdW/SZCz/A1MWN0ufbS0OPbYRkb4n
uMgjsGwzaLVMI5k72ZlU90Ia5yKdK4WPFmlMpMomSEkGrMWfAwolbUPJLttU
LDzZ486sOIynmi7dzVasQHWJrYG46qIPmuyJUjOswHQd5JBjxWzmYf+yoED/
BwyaPy0TP9m/QQMwWalukM+ZLvHqKQP8Rqf09aqalRnUFHp2dWWV/0nk59Cf
Oj/9+2kq/Wh7ZJiwMJc/ZugPRhXxiqmSB2p/JyLWKW7g7LVTb/0OUPV8GNvw
zrmBFT5f5qZ8G00IMqbOq6b4xUeG6K2THVfffCK2MSKyI8BaxB8upfeGqquY
rhYM3zZcSlxFjmMPF7sbd00YLDuflDNqX/nNgz/BR+uvGiIQUelO7InSegIl
z53Q9l0r8oXpTvBfQxKcqTNH8S8XiFs7bei1+rhG18iX0ZwzccgyFdB3Vvy7
FoZwGQfyvr7nE9Wk3fg3sQnqDWEcRAYmYemrXJHl3fAgVpTe6yuVCc+hJHCg
rr8eLLt0eDOXMwE73yt560zlyuq1NqMXtTb6vRBMH0qsEOZQ2bCougCWsZCP
6j9v/QhEKoTwdTHEfCZkLakrKBm4Wotsqx9aOtm5EYTSsDYIQauBpQapNxzg
62GBPGZZ9iqRjHjjRVboitsC847oZA+d5fMtJdcPZvLxKdU0LPGplzusNUO6
K+uZjlQ4yesIU+r8jkN3GrZA1N2LLgF48Te7xZCYm0yVmQo/XXziq8NQNUnI
16nQT3u5s7ixMA67xqcdJY7hSzt6EdCep8OTggLCVRmUVHxMqd23OeOw8sm2
mHQPehPmOun8gB/G7GVUvnEhheOAT8eE1kGGRcXMP0lAGYE2xeueHBfsFOf8
e0JAlEVAY7ctGNORXz+jBXD5WKGZGnWAXzZHYgvAwp4VgpuCaS4o7akgJGcy
NzspvZ0Mkn4v6dhwUPNsO5pKFb6d/BfV9w+VgvDrLyFXfYB8+TUTRBlu4Iwx
8tTyxhNcIDMPj3lMY+G4QxyKft+T2zWB9+arH6nj0YiKrX7FKSdkcf+sGVA/
2OJd6qmOvXhONyuFucWZZpIsR0j7mqzY75kkmw/IwiJfWMJSiFrbpu8W2JWm
Wh+Uu1eh5iY7XcC0/WIP2h1oCAr+N1pOYkVksGeyNGG/VWdPSlD7Ed3N8JPj
uTVMP7JbY/wY8BVJ/X4y5ic0Dc9a/938HHLNIp/7KVdJwPBmdX6ufj7IHv8S
yl/pc2W9wEZt3ULrwcmw6mtJ2srKIXMxJVDeEAxmtHIP8YC95vPUO9esIgqI
IX45jOaPDzyh08wVR+9wzvqH02HLWgqVVVQwhC1a5aDMGccyyyjVfvNajUkw
MYhI7tCLjUEv1KO8d5VDCxqNXHQOqpfCxhygtfDCUFEZRlGC2RcbQQxKRKk3
DNldBsIy8pBkoueohOXfbr/laa2Le3gjcoEtVOXVVnQhepoRPLPtpGqxH/lW
a7EcWfoESKrFnHBsUDRbfzUpbfp4aaNqZ67l9bjdmEO3FUpX/iHwiVuKBwZ/
94bUcBQP7C5rN28ZqmXVE+VId5jpB5G/OKvPYz8645L+173Q5P88YexEDIwM
YgOTSzVdyddCVbIbbjm+0z5OsjU3RMCnNqhUkf+rcgDK3n0C5sDUitIt/omd
6Bfosq0QFR/Ya91xqg5pFsTV41RbS9kQ3JnCjUafStgbRp7b0tmJjkxlqpOD
j6B5Sn1B02B6/DoiorFfG9uf6bStDokAzBsst66/2SkS9C75KwFobG93iZwF
j3sKxS9eYSrSrK3Re+POYbFbFo4tc7gAvH+OGEyZcC8AR5NC2u6RVRr59wbe
GmxJfCWaTZ1lQdc0zhyOfdrH9KHmXYP2Kr468MdVkOPCYTnKZM7Q6RudprxZ
KZudFZTj2xQH6rnOsVCP61j/F4RVz0bT9vDie9pULhN4NJ+ndKmBlgd7I9N3
epbsexkVQoj9xXqmAXsgB6Jz3vlLRCuOU7HHvZFHGbZwM5KJnGbGZOf+igVU
WQGzuTNzFt6vOij2AS9ilu0gHqu/OsWCInAiT9+ggLpkmINuR1MtkYXf39wL
/Q/6/K9Kb1a18xvOKPy3I3cDzHgxcAMrU9ZC/7U99hyJjKtu1zWaDcVRdtL9
ocXf6q00Lmj5eRHzSFOGwrls40dIY8llXMVZN/rJUGzyWMokoKsmOHASysYl
2e3sH+ssD2Rsai5OZP78+ps674/TkHwBrVZO0DvPWZQGmEiRSGlFqpz8xjNs
yvX/dPBKpIlzD6GFPC/2Mr6RhPLlUY8Xvj23CIe70KrLzx2oC6E3NgpZUlC8
aW/nR7vOrkFqV+/kZ5WT0T4ZUTmA1C1htkxzp5JzE3raI0JEq7vMio4O9p0Y
+T3qqqGV8n075HkspZjFJMOnRz3zGvOBWPfX+CxHylfvvENnziFQg0EcpE+h
ZPd7Ia74fLjzUucOg7I0yb+yGShjkyd8xSi0p0GsfR3934/R/He7iuV4iMeF
WigQG4AmveadbiTpz6I9bShNNBs2dB8+Bb4OW6UdfXP8Ngv7WyZdGj2dh6fA
4hiMasp4DcettrFRJAx1F1ngGZcjuW/SWFOLLji3uorMaKwQvcFdPxzKBI1n
pbXr6Jf1C9Pnx9cY1/lOs4RyV4zvdwIcapzDs4oouiBJda06mXRmEe4XjFYd
saZb2b3vV1/I9NmyBROMUhAbqkC1zALk6DafUQ9fbOk0fjWvZQkVVakM9B9i
y3MJg0csASjlkkl72efOG0eOsTWKUxqdsIQUkkeiR40E9XwQkcJ3yVDkfbW3
3GvrFlhKqKa9/rVtWxkx7jmQqK5pl3iuqckWMZXbYk5LW4R+X3Y5+JlJQGqu
j8xr3EyQGGynsAG/A0Rnt/mlNLvi6WPg69f/qof3Sx0VNx4jr8EX3rpr9CmM
MGfQsj3dMHxISMgjcd6ETidvSqvfjvhLu2AQl3sivdJOaJnKuI+TQnFr4+sz
MT1r5aDnZR15IJqc0m+ibXI45Bw/ArI10n9E1RyEoe+Ouz6fleX346I7IqM5
sVC4dHb0/6zm43s2Q1QRu9x+ocKsZ/0NBTbfP56D91qqLCo82NN8eTwngarh
GeuS73S6xkTVbQhV375yQ0W5axexDhvnkpP8oT/GlUC1eE3BXSvlIGLOY2I9
9QXIm+12WAnnrhRBCppKxBYGzCrYCAzKeL4EHM32idePjbyrWMiyfIEQSDQI
9Hl0Ch1m8G44OtCameXE1UIKu+bIgv4L34lilmwyFj0KGtuFYoku51sGO/Wl
KyEkek0kyLvN0vq5tjZDgXscX0p4EwF1L+ptB8PZPnvFb7FgTzydzImahPS+
6nxUCixbP4ztFE6KR1KpovuYFHLThLV7ZBTIZMntDfVFaQQZvTdsDUqmFgHV
+C2rjy8sxjn8ojmWDFW4vVgMlTq6q9yY2xBsl8kDRaOWpWMPPN8BXSEstLz/
tKuI8orKa6PirFtPm2b2nLgmaLpL7DZkJh0vjXNoJ4fPm4LLMefXYCPk9uRK
1l7bPQOLjFuKQZqkAaATYZZ8JO6REYlanZJvzeZXXNjelhrHUHNy3nm7/Svt
RH1mpEIyKe3JfcfiJg82lFPsx3tmASyNv5uK6Zc/Xp7coVD4OMiPyVdAI2l8
MsJNlKQSWoffab4DoFgfdCTK3Fhq2qozWIchG8HwcczFJ0IZxzl2Q3KsYuoe
5W/g2WkJx4BKW2C2R4caK3PCi/YMf/p0Kv00k/PT3rJBKS+U+AoNyuDbWXZI
Ylm0eX2jlSRL1krDsG6JJVVJm5OTb50wdOLxx2QAyYfDTSGAFZjdmoXTdXlF
4/AAbk0XeAAX9SEoFRNNxui6Tar2FPnndhRlFpaJA8kftv5AJRSt8yCWTjB+
KcJjLdiRhKRgJr6cUjxCnpBwClIBW8wW71nW9nw7X8jN5L8AMv3uAEY5ZvUE
8lPs/9XpXHEaexInyJ98pfircYqmsEpZnPNAwqSJaS6YXvF39ZbjLkqhw/OK
jnQ5FWwE+3luer+cOr27S0yOP8ErtTm+MiDLGkYH2xSb2VNYl4+eLqUZVejX
GaUlyGXVw7PBWIM7Ax/GEGmZj1JYBiYWKyTEBoPZy/96fO2wZ93mcijLptog
iPFOCBeHtNylaIraeGXgj51u7AFEBxPRXrLjA97K72yozVlNBnKN0hLXR6/C
lmHBZUXXEw2/cElWn2ei3IVDz3sKF5HhqG/d8Z/kIAvOTxK1WV2qz5EIMMjn
1V/5fgt8umqED6hQVhqsibmi4M2H1vVA61CWqvf989JSfif9+LIppmdir/B7
+XDo8cKNk/PR6kC+Mj5PgQ5F50FGLgi5JQGwwqWJyfLpStoaUtTaeqUE4+IE
GRxeLa2L5RCE0dSqErozXEm5+Q6Cp83W/ZR4ia0n0prhYu4mtpJiV+FTnAQd
8vGLKbIiKdQt/jvo04JEbYh/DLbRYIXvCDqOTsFVA/DpO00K1BR98oGEUgZL
fZFAqBwWyRU75HbwIzcfsf5M910EYiGldI8AtTjfQAKMqM6DAHBN968/a9vz
UbLaPKe+dF6bxWETMJEBxfX5FMTtTAfJrnMIPdCYkXnhRfJ3uP92hB8OpNyt
86WshOk7emK6x+T9cCMf1CXPhcijqPoiv2Dgq12ltefyZVGomYJkecemwBGA
TXh54TcfBQkDf3BEU5ldJPqWUgS++3eayFLsKoZZ1vrWCNVF8JVdPFM2fI4h
wZ7MAV5V31tJNBNPvPoT3X1vrxIRoHArIKiuTtWAZe+4LQLzAQQmf+ubHqWG
C8yxTj7xHs9IK3Ov4jcydYhjo3ez+PtQ51lX/ef57jDjwhfVJd1bLy7YU+1p
7fghWverds8LOND6gDuNd2lzyPJ70W8QntxVUw6TitMiOr3bM5IjpKmAYWJ0
d2RTRgjL/nD5dKenPNUdrqqb+5ml25jCu2MiKT2XlbvGVrNc01/Xd+YS4I5B
4D//Obtr0c4JzCNkvEPZ2Rb8nQvOQkEoIoG3XG8nuFCoLZu6x8oG5QxIitYp
fckHEDAnqUYchdG/yYpYRNA1wbroRDNGWO/BEy8raPb5ITkHpObozXHdne8r
JNz2y+Ng/aebOdXvUMZuUdOy5qbE1JiwJpsEpkLanZPgVmF3GHmIpvw0ruwj
a0T4Xx+3QXFBc0rHGq0nMU/7Kt0fTUz+5bNVgayPXLH//SFT4Y5ztRGtwSHC
dBlcB66ojELkSUnVor0K2rUJftXRCVcHVXIgv4tifvsVJW8MvKGNbGf8s5xe
zCmsQ0xD4o3+aBzufX+6s53VOWQkptHoelQB9xcahLY2wEOgJq5f41CvUT3x
1Mnhra6gG1q/C/BE6sqqsSTo/EsywItiBmPrd1jyBw9pdm1HpVTdDC4v9R1V
d8NWCg9ahT9QBs0eRs1cOKDxqxlqJjXVSah3YrzaHTYJcoCJliACunnUGcRk
6epSKiR8LU1rC8P7PNTXUJb2uTCA255eFcILz86hnWXNa7ySmQsfJ4/LkUpm
XRyeCaJ6HjLLaB6ZVrKStix1NR4nYyve80015d8URaqk5JFOyNJBDD5dR7z5
xKMyBWHkfSPhOZvNv4AfBBYt/PZwFTB76w/JyIi0gHl5pcbFgFfbIpPIV+r6
iJ8Yqym/JeTJQIw38jdLrPXKmurwF1EQnQXY3bbY9plrAkbBpU5TZ6CniXsU
+1f2Yd624Fpw0rW2zWkuJfCfaz/0fOAV1PGE+iROJsCBIwWIWmSP4uwMk4D8
Ped8AlNNN8I2dMdd97fZsgxtTDhAcEyXCWqqD/0x2ltcZ+3l3RYINi9jQZdR
+IsM+tSj60+tgqRSj0Lr0wlqqKQzY773Bb1JeLCjBxh3sBjZy8q5LZGJZbn+
ZAa5SsBFB6m7EN0wdIqFR9s1Oz0esymFlyP5+GBRSkIdFlwE7UrH55PtWT+e
D51ztotlIYfnp7Z6gC7hDvIVYpatFPAdFvdLK5omCmBvDoyZ92dsMV9h2SZT
QI2IHuix9+3iX2NR/SJWYewjhggU5A3bCSG/1u4XfrV3acwL6Ya6ibczxh5i
SeZpcrz8oIDtsJjmRdcceHXzMQsAN/jnRUiKWBSNEw4upbF8Ps7XEu6E4zMC
CEH0cli21NuV+24LHIYXIY0I/4ViBfUdV1yrN86kR5EkVMlk6HJnK6M8Th+0
6/l822OKSXlhuKS1UU6XmtLlGQ0fr2dFsXeLmA76RXLjXczvS/jzOIWJwrkC
yBVq72o1i3E/UOBKSNFxUooL99YUatD6E+B+5wxqw2U4zXVbfBscA9rsqIZ5
hGdASLBo6iXj94YJO9TDSw8vltWAi4G/Fl1HiYWzGNIAMYKSjP6w3z8ozdK4
qg6wAO876CIKiH9698xJYuAm+Jmhc5KWlHncGngreRjVwQK+qjvVOOKuDlHE
s2avxZPYdddIb7K7CxKU5iKhS9ZErPARe4S3iSmn4k5arnRBBi31cqy/9nE8
/GlSTYkLcrIrKH9Vnme6IiSgfnqdCRzhEg+i/siMb8IyEKy+erRVXVoY0kZO
LVH7n2PdhKIDvbYaHAc/GHxlbWvrM6K3ln2/wkb/RETyd2XJJonoY1BrI6EW
pmhv5A6YmqqNAK0+UiH+DauYOshW/ID0xCwHe65Tzf4zL5B7ltvbm8HMMdAG
iICiqouYvF0p34pHzvElrIIOYZcZsEQFaGw0YhQb7lvr241qEGh+kUYHHcvd
Of5ktAEnKKKOdwwaUigXl6GPHH55uPP4wQEVjhCQn0vwgYKdaCYAopFdkBZ4
0SJ48jwFWWNUq1O2ApUmUuWhwLP4VSFwY1FLRKLJN/wsalqQVCJq+CxSysio
DDX20sOr9bz5Dg3uOcm65L/KIdMa3MzLluClEeCetgevUzaYsRo2VwM/jSjG
MPD7tnK8GlsmXgw9dV7XisdeRBDtH7mtKehb1qHuhbzvHgxKoAgkO3+NrwmT
U8Cx+cnVMs5KVsN1hN4cPkdYXlYZIBObMOKxpPVUHqJmQnRvALFJAORiygeG
k3xwhah7nvTta1aks8Z2o72FGDCww7nox9PENFzaOB6xu3r1g7BA+J/ex1eg
3zGG5Skmlz6PhUYIUlxTCVJ/3u5PVrxiV4ZcwpIilR+cw67Y0BbNGHGHbw8x
bzJUT/0FkabW68UIPrndmTLzDPJdHNBGKdoHS2Z37rBkTd8b5ZWN/7Uh7W/8
l41IKpaK5fdoSu2zdriXTRo095hrtieFl0EUMCIHfmq3jDT9mkkk8OYP4AGU
VQWfFvCwG6nWCL3WqVlvHjY9MjhrqHY4rh28RdHMsXQZcpS/eYiJU7ouJsvp
fcwwlZpZyyESN3O5w3EPpXH44PNC9y/O/xU45F/We8It6YGUMiGi3100XvDH
VHSIQH/wrwEApm03BIx/JprhOA0x7XJ/Fk1RsoIJzkVGXljGdveoWC/f+QYn
dOmdhnA+6AujP/AQrcgUuBhhyoxQOf7iM6oMd7T3rB57NkYnEGdnCzrc1yzq
PAFa9+ZkQ5lRJlCmLavPnAoX44T3gaSto+n3rlgR03s2gA3cbINHo1+oZpWt
00xtItgmhuhOuAkil+RO+C9Lz1AmyjpcM/WzCFz5XgWxge8FIh35tITQh125
3423o6ZGEra7sdZc9qJPK8DmO7HHQ/Ho2omcIjjpX1OJizUJJba2Fy2MdTos
FlvkUisXwlQgoETkaPYROJvReeQxrcuMNNuh786onJFXCMEXV6OI+vwEEvt8
XmurcpQnqsGVAk6IHzZvkUvGo38XIXWA1487nTXvzBwvQcLosNhL+k6XgRy9
FnaJty7yXFN7brhW2B5oaeFP96xZKEsfSsh1QXFOFofAsJUC37+629h6ufL8
bwVFKBsev4fWW0yzecyCay2pdmKB7gWvtwaWwWOH861uWbHrjHwtCYmkSIv6
S1AYL0F6N1Tydm7MrBf8MNuBAvaZQ+EhHN5xGUp83kAJ5hDjRBNzCGDPq8hi
A4kz51unj5THdxqwJdRXnGmh/im/Pj/znIjxJCppkIX+8Bp6XTmaL+IcAowk
yZRmsWA8HaETkZKLb99YGuGp7qByW4o9sx3+O9+KoocIvrJC9ionSmOI1Ajy
JgyHVYO5+aZCl0CZtmbijH7BF0zbJmcvrvdkE0acZz4wcxQ7TNqrACHizTTZ
yxNG5XDFQ8/sf2yFGZfKKsslSZ3k1ySzCdUnBlGpIdGKacS1rriGIX7b3/uI
9grrpjJM2W5QcUMKx5WCrCvdi+AQXs6f8dCtOSFXiTEtZIx47EPGpeTEKd7n
T5aCOw4QVj7K9oQnXQYMqGIG0A3A9tMIKfZJLD1GboGz7zvNnU1w1uEV7xXU
bregQpf5PgkXKW6r/9paJmEcBEIqnG9F+OY2iQEk/FLiUbVn/IL81Im51QH+
IVualuCZKvJ50Srlfqu9djcze0czCo11o1eYigxuSL1fG1qmPbVOMUnN9eb3
hUIeRPFYQ1kXUh41aC9ztMEu6jBSc42nXCbFAyp+5pKdBbIKvIQAR0h6BGiw
M3NT4Hxs9Gslcdr8YObyq4h86IpbTafVoDvrq0WCzXe8EUX+wAnDl5Nbm/ok
1BnTL15EcR66GORqEmozUQs7yYG/HWMmF9HH1649FHBLmD0aJARBxp7cxTH/
OTcxxypMnzg8cSezy+cccECuSHU/EqWLmuusDROZtMPnZXIyWsgum5yQDans
AXmASn+UD5oAscs9t29LpAfiUxwLyHZUY7SlLr9POM1+saz9z14EXw/fI2xZ
IIt8Bleb2AvgqgHWLwDvL6eKQ0oczxeWBqMdNkOAopWUme5myzAQFdsl2VUD
/wVhytxiujhUDDcaJfrL2yFbh94nNK+s/0nbrPOdo+5j1/NYq6pC/zclWtzc
Oud6fJNNVTg1gU9472Te2FO1oZXxXvaNcLUoLw+82pW7lzl+inxxeLcTQhDf
yMVhK7jnHhN43GV6wyEjuTZEx39MipkKUgdh3YW3uU4fsMexPJhIIrDZbElD
5Oy6w5mKj6+MkKAFbePEcnNxZkL+ZObHVWUWII5oSoPLDMQP2YpWWfrXFjVd
SFTv+etMOtoFKywwebAuCASzCHsccXDCzVvhB/u5nyVDwmAUeiRnoGHuN4am
mOo6rYcI2pzSamk3fUyFurzUMjKzAz3pNQ/Qio/14hHMwLGFsDQwhOeCyBfO
TCFy9EniUf3kxOJk08VubfwK4XdQ3bvbesy5ikRR8sS4OJuuYRjbcLUINo93
Kuwpq+bM3ZQp3Ng8O4C0gfjUhU4462Z3Df202z62bN8nmEK3XwJqiC+XSNg8
JHVsdAecby94diAzkVG4M2AeuNWeqrRX0wka56kC4yUNPOgjHLB9nkxZy5Q5
cgh6N20GpknS1Uth2DvmycmHAXE9pCyD0FkEyMnedy8z2VdBZEPZzzI6Tv7c
s5F5t9tfhZWhMXefzEgBBKwUnTZMXekqgbzIdoLYVWc+uwKFyvGdgPcoczuA
iqtCC6l2uMryfObLPHu1W72s56rlxJJykWNP6bE4VGqaTGn96UNl0CzRGaRb
v8VdiVkQMtYuDU02hk9Q0nl/UkEkxtGI5VyaEyTFvO9wAfUTnpHyATYVMzrT
TYYaEdbLNvzVrmRdDUR4murj8wN33LmOW0cPP4hMJdGdUiJ/rUKdkcyJpp/y
lgwXp+cEJL+1dqdZ7Q/rfim6YXzxi/OEsSZrXwY3TF8eVBotCbkohDFxmnbD
ytVUxNAyHT/i6Dwiu0eBhPYoAEW6W937DJgScKzCfTuBiID7Ql22GlAKGkvY
CG3anemykqpl3ebfFYtCfpS5FD02/y2hr8yeJy2U5KYFcWbhepcm2EExGSPc
aI8UCs+ex06Kg45xA1Qqc5eKQNdfawsv8m4VbcPKo3BvU6PbOR8wioXlg1iT
76klvgSqh8IxUZoFlOFPxJheURZpOj0vFv8tq1ngi+g0hfCmXA+qoNpTWT36
Ir7RQi8ZbOCQcnBuHieaP7dKL/1PUWjX6lktbykbFmfMjhFiSzUbxAYvQRaO
XBKtfS4C9MyVR21HyO9bs1oc0SMcEZMyzncFqcFj5+DH7JRfM26YOqJBF1jr
bX0s/5g1bGLvx/na1thgGuAHwB66RuWbuXxpqfnHGkYPeW4yldesOGcFK/ew
L4bdAFWVEB4ORs7FnGhMPW9XpbY6q1BOBWjfgiyfTluFW1lYqRSRZKcAu+WP
UwHjdBOZm0P0Zt/Fr+a6gxoTKhqJSnBCZv7x4Vhrn7wyZwRQpUJH2LS8OxWA
v3aqtXxq7K86JI+qz9XTbmI7/g/aRVt208IaBz5+4JSpoRVqcR47wvKPKVYD
GYB7rvENo0hGEwSNTYi3eZg+dnyRi9eDppRJ+cjudDALnqoHFyLer7t5l93b
IZ+Jd0TpiJGTWuqqsHmjqikO7au2mle6I0adlzNRgv3Wt7vR1wcaEc5VuyBQ
X8rE6upxEy+VtV7b3N5N4H+apOthTDu6dw1G8YflY0vJDsKdnQXI5Jp4+R14
NMpPNlkp3kboYA2aEgx+DskBQZ7ZbRjNf8f9MKJMCQdCzM9lo2gbLoW4WMJ/
z8VzNUCnvyr7HSGOPNQLAXy3nmWqcbJMxeVCVBV6bRt1y9xoE2rbdg2t1wVY
CTXuweY6gGVWJVnaROmAjf2ayl8i1/sF2nNDCHUEO6wf3yC5LCni6eUf/XoB
+WMpnUk6EgHZ0XeKY//IQol7fCJ0hSU3KZuHjw7RqaEREDm1K6u7kTkEKLE+
en06E0OYDJolJiu9sjIqW+v+wqPV1UvI73gcSmGAG1aR5HADBptLcGryvm5M
GJR8g1QeFNyJdYpZwLKRvJ4EDwoB9If6bf40R20W8HYeqw4WujhqMpOdTnkK
IyTIM7gTOVVBiXsOdaNk+IQuFSciqnZh/WBpHXRuoNGyDjhBSojvVFFon5LB
prdxhNBjdJeAxx69NQ+49i4R5ksitta7O937FHPOQcG/HBmF/++lhigHZD08
UxA4SaWWg/AH5VSdPycyv2Do31KIdM+Y2EsNs0HfQ7Vm513Ndzml5SmYZxab
jfn+WXAMcd2r+YZnsF5yWq8oDD5PQXoRErJSfoFEO3MXLrCFLxXtyOkXF/9X
XjvADjy5vfwUxKrmpG3FaGXslClxWDrnRIN8QmJxWTNMSQ2f0xY5IoXsWhfQ
tXuTulxluszQ6UCAeNNYmmOHawm/TllI3mgOfebJZddTTBFrJDj0tkcADBHg
bThsZdkj5Ja3VEbJoTwrKPCRIjxkV416QcP8mVPoTFFKMjgY5Z41mO14VFfp
N7Ht9Fzig71CkKoUFsPLohbsdwSjH0hb8hUO7lCQ7zdvwhWyuNzOUVJHrBjd
EY8bBZ7/5LLgJ0feZ8Aor03EjnO+TGDTarCRPKWnstWhTr1By/RDj///PLhX
s/rQj6p7S9IMyvkgAVsGF7v62sIk/Rcn63Kkdoz33D31iI3GqOJIRmYMY2B+
ZRvGsTTdORuD3UmvjRZ1Y1kLVuVTfhw1MvvTWIGRC3EDkG2O6VqDrtdbDg1h
ybVmXQxcrcITmk8zt6KF0uB0gzjAu1pss4rFuT2+VC/WfjXwnzVPibqqs22d
m7vV1eUb+1Vs31CUlk2CmdanLBnN80Kf5tZnArSRalZiFxz0tY0cmEdX1UYv
W7befEfNI+8s82R/QG37mqD/rEZjU0d9yTPkZPVx6jn7DXrv/CuzvljnvMfS
aX5uhhrp8N5nsYJLfBCygY3EhQsuRLtV4wEr8ebTAayFzE5kBuJLhooYOqKR
chztOb7Xn7/9Yu/RekdTo97ggoBqby34QQzU7gg9EAa3oTJ+tt18P1A1dujC
C59qPLsSMwXaDDKXNI3BGO+0ZfYs8U0W8f6IpjpUJE+OokSr+70PKOvenuls
RTmOGvc6f52XpQtkhFKkTZpAO5Bpe1dthYYlZ6zIXXzdBoLbqCmCbZ+AYt/8
1bZHbZ1MiC+I7XcHDKJitC8bx6BrvL7T2KrzydjS2WT+9xv+P7gY99jhpQr8
LUA0bJqXHdDY+gRGs7JM9ahJCRONr8aeDr8alcRksmU4AU0DIb8Sj32AcODT
Ira2KH2kTnIyMpt8mRKslaYtrcPuz0YkUj4Xa43lqOb3+Isin5cwtHBOPINI
pSB9jufw0lyivlY9OvSK7Dk3ro8mItuyLxnyaDm0dnYeQQTHiXQ657AQnYSb
WaReEmIs+uNV1zvZqIY4NT/gah4/G/ZYjdiUUR92keQEqTxoahV7NMbFHJxQ
Kgh4cRxrG1Kd6apwwlrtVtLm8yNZXXVV5JoZtUkSL68pnQHvrWeQApZOK99Q
qY6V7/b8z5OndZlv2Zv3abGYefEYv0pqsZxaYpQ2SmrcyRAQxPfdEnOYL8ep
PZp9QiZqcyK0YZlfMyxCmnp43Kvn1p//FzJaILcJrkoBz8CZIuCQuvDDilRg
b6fd+gJsyIAT8eQrxTomqwB4LaG2XV3b3guZjdL/H/FxZU0OZQg2RAnq5jWg
+7wUpxDFG3GJ4Q/f++7mbskPCxC1PF0fWCj7oxaI3g9DKAPmb1c71dqkHu05
hYszC1drXsAN8dCXv+vLLw6ZMgrAd37U8RXTr4IcbVsCFn0Ayh+rIXfnbKGv
aNjKaILa3hu6w9+lXRXkf99bufzPn0X78cI6/B57npX7mELKPBmEFmt5gHHo
WZz3babZg2gyRYXgbdrNUbKYCf1SsRfAgSN3Oxstzddn4hCgEmDwlhKTOk9w
xLdnpCx5w0nsAPeh7XtrX+hlFzehNqZz89OFVEUD96NQATPgNgBhn4a1kZbU
qA41se+2sxTw+FulqZxgC0e5Eg97Y5hgGhYWt00Ph8LHTfaI5dHP6GEYkK4S
Stf3FZ6Fc3fvVb8HtVDwCSlQs1H6+dJCpJo8Qsd5yOeJ3wcjcBFkNxn1az9G
C6ig5tp37OigRr95tjj2lWrZIpLc5+uYax2OVoHPKFLTKy8dU9plLJT9lr+d
W9ESXRSsbd3od69Kji7da3JqfOxPaveGi8nhiZa4zdfrUleRYwSfmYWbZoaS
0BN8MxYfXoCn24WALYvJz4qIwzNRtUe8SGzcJxBE2AtMe7Ld9b/Arqtm/3RG
NSPyX+olRxpAkQSbFLV8uDKb8hEaKYrqbTJaNlL56PYfcE8EOxQxPqasE6ro
QQaGf2h1AMgw1eCOpEESU+BoSdiJyGa1Q3NFO5p8hi42sHSk6mQL5o9Cr1H0
Rhs3R1fr+O3j/kWqoxZvma9MEMlt4K/EVgt6Tx7z+Fd8UveSTMoYWLVEF+GT
xFlyL4dYvZv7KJ3lILEJbdAZwGUpEBgBu5zNIuHEPMI5iendy9bal/k1/3AO
xGSceR6b1+6+IAl8/Yiouwnw4zK4q3XRV6Pvhs7Kwbr67ikPGSlMxweau13G
lpoKBToWaIWBdIMwdUI3kdftrHJyhi1lysqrDGsTICbQX63xm25tgk8kE4lI
6bkGluirIkQ0H459Z7Q6h9y3ZaBwb4im/1zwkw0F7SXUdiIZnqon7GjLPJX6
2AMwBvAJ5uASoDY03vOsFGUJ3tNU17lciACZeUiYfQZObzhl+4dSa82ObNIb
WEeCiisGdqtqYa6J9uthMVScw9uJk511T9e3jAZC3zp8H8dydTL8lC8XmFuH
uuiyn5EJzwhCzuwigte+C2PUW8/yYPmATeBA0tZkgoZ9XIMB0Z8DshG7754q
5IxOwdEEonH1rfzGc43Dd5P7k6smNgd62XSNEKkTpG5cL3eyzzW1MYs8XV7L
QPwXClHb8djJ2HcY3b8j9KfXHF6/+ebZLNWtpIJoNrP0JrqO899CvlTrtlC+
qconTwsV5kILY0yfyf7bQyLOdr1Kx+wW4Xxj/5ZRGPb52mbPGkaqzX+8oTq4
6reFdM9ClpZOx87+7LXJCwBU6W/pJwM4imt5EBUMbYU3j3mUvVOSaeIiUEMC
uBXiUkh4naXRjE5eH3sS/mivXOgEuWvUL1P+xwYo3b8t3crnf/9r8/b2PI28
uqcBgYBCBQS3VU77eBo7XDY0nNnySeyIOZRBpzwBVc/B9srnYkSFBKe9AyS1
oWATWd3FRYncDE4ytUrnNludvuNOfMcp3pitT1aVkpuHH9rLpcaGGKQCBuGy
j2/TET3sVgkq0YSrN0EYOdn/0ry7ww+bsJjTvD9NjuziDE/VZ1j3pkASdMHg
rEA2WybXf1+VBmNaWJD1BCWr6j1vHPOaxcxowgRWf4Irl5fGE2g+6t3aI3mq
dV28upl+68Ik8s/xo3Pt9pxhHT4j7z24ZY8UK6kMmMffvLJ+XWp4Tg1FvuFh
tZzZKruwlzj2631EKEiMVM1ZF6qIG7j3jkS3xu0jEqWQykaLp34T49yPpUVQ
jGRu0eVkGT3HeBVzA5kHAuUnGsN/Exn3aPkXTbf/YsU5hd/8RU4/3MezxHOp
/jJSbEonf56wDTfni6x4qg6OGpILeSZ22CbWpfIX82Ta1nJsQrjwb1w/PAwH
AhDki9Eur5xX8XVAvp7ewmWJSjCAFFEzNZCh8COriXz5/J4fKbcDaVCuZ5lP
L5XeB04yf2YjUoMU81GM96d6dSAVhh3GaUzUxJvlNP/RVsvXo0vZDMfGXdfd
l8udTefKqKWXabe0jWopc0Xm9SLHrlb5BSEhsOv8i+3VIzLboYUNxjXyc2qb
pzbiFl9QcbYGzpI4p/FMdW78hwGSf3mVRm74sufwi7xmv1Z58R67DCeulOUz
YwBfIKDOL4jT6p6nO0E3TqOMpM3Vq4CGT+vK3W7UBQdvUHWcqTB9c52YxG5m
pI0Liy6MvfORNv71dFOVGYEhbpEK5UQXwzwXaOB36pQx6t0rdg1fqx/V4nwB
ldHjIn5a/IZ2Bb/BAm/LeGfmWtkGS/FoMPN6cRmdLQrn6dJTcp/3VpvSCAMn
2mobZ/59NTMcZNsy8HziyENw5iDPxz9pOiahjlTlg76GJfCE0XlQOEnE953l
GapTxvdT4QUIYXSe9MLYIO4fMa+lqI8RRkSSoXQJLqKd8/UwBb0wmKK+lMpx
2hAv2EyHdYPhcDDEwxbtH0W72efzJ9iGj9SLgb8kyLOnhWtmGe+PVyRD21Mb
GZbiI8X/MScxUO6m8/GXq1GY6bfQy2j7XCKL9WO12w7RA/+OmGSScGCR0neB
spLZ3yfAGnl10HWEvwcUu3UOXHyGB5r6QlFeto4Jn2TbWeV/mWrX63S3tCJ1
vPsv0NqwqPU91S9sAIBKlaebMrOGFd5wz9IMbtcH0HBaAdCN4ALvhXcWpEBQ
bu+1zU9Y7ZN3Hhy+9aqN0MryP4DeCHQDdmKpRtI1DRSrmvXaXJgIZFZisWr1
WT+PG4oQ1T3wSSt3akQn52OU0DUM0kS+CgipHOJPZhG6RESwEPv+TIKG1f9O
/vYfaM2SaAd0i/ZEP7ytSGCOu0+hpeXQnzC+LhTvgpoHf5Y+A8aV4M0zrUle
dLXBJrTyZudKgLFiIbHKk7agHTI8t5tEB7NXkg6tSga52+bz56goZYhUvSd1
qh/lnclVhUK+l9wfmzK8pcuQJgXGkSAM+HNxOAK4DzBj5q3F9C9KO0bEe8kp
fqeM1uRzF33XKWjZxRieqg+I/jgwuKiAWHydLTIX6ffzw1VHk/xZ8+Tzam0r
VCOUkxNONjVEYkoTDJul2BzDSE5N0TDNf0tsFgSB5Vg2hK5lex6NNAvD146w
BzjAITzMvMcy4FPVo29hnpepVEr/ek84DLWEHG0yokZTt1eLrB5/rQE5wFF5
x5RzCb/rVjByMAnRrWAmqYjqIpxxNPa0OP9Hcfsj0MMIvAx5zLg1l4mZF3G7
b+58sSjLpuDGe8CM9U2db8k8+PTZ/KRu5bHn2eenu1z7QzfPor8gZf+rVZho
SlN5ammfjeeOUTr5WBuSJUltsfD2K5f5BDn2mVGlRI4N91jNcQj+eBl8i3o8
GFUa70UtVvCFTK7Rki3KhzjhCBfS+cqZjo/TdYc2B4uLh47IISbjJLk2l4aX
V1XTQlWdo87HReUDOnVeUilMs+bxhiKvRC8fTa6C2dF47sKJffOAP1nmJ4iB
SmwF4HFHLraEHYJIoabloclIuQQt7WuOGQAEOHVbzzIyOBXmewNBRSDxt3hc
lvvzWV3BcZrrSqnwDvlNrkVqweOrmIMlBzZVjAOkTo+ngGbL+QeNCc0w8ZyU
Z5U6oZzZug91pkkmVEA5lUt/PxuGxd5Xwtds36mhR11uuacXrSmIgw6HWVyJ
s0nQMuq1bioQ5EHcs6G+qrC6Sys3YRJMu5lUEW3/cFxPGi+zy4C4gIIgzg9X
olLf6groAYLYpgf0Y0avPL9AvgUxJ+NVa2Aga7m2DaA2QIqu0+ctEyYBH4m3
hI/Dsyr5KdMZHG0gFagt3Eh6s/ffiTjDUqlLr2ZxfAKjBtSnPGbFJ036wJPW
meuPCyBgdUOaoTcIVWokwJNvsCqYiIXhpcSrt/lJmpHXWrEixlOlWzDQXKQF
C/vXgJtoxh0G9EcyidyHIzkji4Bys2RDtSPjPQ6pRHjiVNiNjDaUSKveFfu5
HAtk8xI/KaBmipcRXXdHJsbHLmATlBE58+rtKJ5iqWyNgKfN/NzL7xuCGen9
baO+DRp7BCFCV30PotuPIVkZLjHhFwfJPnVl1Ra8C44dds69/CE0mw3CLnXG
B5vpgM98cF99kkAGT1IZnmxGu+PfhCrS+Q0oflgAzXJPybrVAwsOh5dOFX7D
S66/SOwoQrojkq0LOqWGJbldUWfz0mLT5REmorL+A4WrSoR1rTcgVN54AzzL
51L9ebsp4gBoN25/t2jMSoI/BSFivAVuTekAb44PXNZIwN7whekMfDLyZ9jT
/Ced31McSjWa1WkS5B2AejJi8KNVdEti0G+7j/UfjAOCd2eFZDjLze8b0WWQ
tcFaLYNZ2IcgQungELS7yNC+32983+SmcqbN9PhX4kitf2ywNuzZsHr4o4b1
6jWdDDms23yYWkqkM3glWgv+qBaDVqosWvxiVFAY4+J2Mb6iitP4kngRIhJx
jtgIgAvgWMjKJCCf5GLVML2BOzJHOm2Qf48ayMJAhbTyBuqXIzEZ+2z85EYf
Pppt4qB7kRq3l49Hao2XBVLXr4+CG9rjhoYdS6f5nZ5PsZ3PwFHhtiF2jazQ
0X3e6DGuuyouH4ALVBoK4OeMZK/nh6QpasBTBPjhvNYUqPsAMKoJzAExnC94
luIzaMqNbmjxFg350TNREHsb3Dh4vufQCjcVLC2+1y38KbT0LpWtSGTJWySY
Q5i8Zj77hLapMhDP2h//WgvGcy29ehqYrtqYJ7rvHi2Dmfzk40bJF+Apt35z
BqvYyUgxutSzbIYRQIhpiiITnXz7GAtZrrP25F7ZYURrgJ6UdBb5k7zuJOM2
vwEBvqc4eqan7U429BSOy9ARNhAB2FJV1zcy+vv4P5RWG4xANXtT9wwfxI0x
PVfHIvW+338ssakx1GnmFGP3Erj4NzuyBFE7So88X4H0X6n7UlRQ+4SncmSj
pc2xFbB+DeXiW0EyhzJIpL6G+hO3vqcghcGKpLKqtsGC9vDSMzYy9D/ujNJv
t1X6oIW7SP4LyN6z1KTp0xp4Uq5bf/TV2A7lG9kUVQ9Y58eXfH5cyVbO3vDs
Fh5pI4QL0xpcFQP/3PJdGmIx2YSx230wciU3PoAoDfIWx/clxcwAsaNumEK/
S79FRSihjFMMsuqYHQdoqgdWDEg93nQfg6zYSBsJRStnqy33Tl+n7PWx18Pu
SuQQ0av8ZuxQYgzDTAogmP/8oehraVCk1rq+EA6CD6F8LVlmjkG6JCVMjrue
A+5FO72owj6vOvz2HrJ12vljqez5irFXKpXD5KB3188DhDtS2H9Rmz3bXs2r
NDK8FbklOIrfY56FP3obwex/w2GpgIdphqk0vKMXfclxpdc95LPTspggFOlu
SiI1qf8kc9WtwqGr7P1IyO1Wlx+LMtashm7LJY0yHxiGLsV/AHSqn7xWRiQp
4cKjQyk88aBSltdDWv/SXfDH8PhfuEmtc3hyMdF5shwfCFrIwvrTw7CCkfSb
7xwQ4RKi/QZuGXgX4IPCMcHwfcoGs8R8nbhzgJ2rIT8Bij1qlkLH5/jCV2WM
f5kHOGmx4pi0bHjvNyTP2UTDre6uJ2mSeuM7SaKImqHT+eGSjw7UFdJmo4lK
6WNx2aThAUZWsPW22gRuo8mRKKnqo/SVuUqWjj7IBFrE9/PXbMzeJAYNaWfp
+OO99virFwCrrTS8ROEpcO92a8lO2A099D5B3kaLGA0nkdsWVmjNQcfu9uvw
fUCsFeYRn16BXeEXVecJPga4bPT4c6V+gweKVF9xNhDFGH6pd8v+hAr/ypWN
4XLl46ABg29V3Y2MEjkI/ODgy8LTlUJJrMkvKjfqw8Ymwjwh//VRDY+h+NSn
9uiiIs3cD1vwSbjFFskkMRqEtTHhiYroTarPuw3Hwx5b4ANf/GC+j3t0nMz+
onXzEdqAiGrrJoGvWb3jxjW/Oa4afKIFo7TvEhw/RdpnGjv0R+MryYWveGxA
5mIoiasqRh4GWGidvT+2LOq94rvNEv1qb1o89EneCrbOSGgx2aqYldEW8MaM
kPercT3x3mg1oqhZ1mEyh8HM2LC6R2v4pv9uam0MtMQAOivsL+vKQXbEMll/
B0YRWf44fYRueVqSZbrLOnc7sQk/6l9RI94cS2v55NDSHu3GF8LhGY2E5TYw
o8P5TM7GfymdS546I7bvCpXMUJUBJeslv6a7hYnXyLOb+VV3XsBkynHJbQyx
Trs2jtEFZzQ/kKBQzCrihIt8ZeBCQmKNU3YnChJMrKGmjQ1+rzirYT9hpoIw
tEiDxbwDli97uCBnaXw/aJ5xOY9IMxl2F6pz18qogvMAYQs895dzMqahwoN/
XYUZrwaJV+uRTJ8LNmnc6erYB4Ik+oaAFOAKKSTV38X9Uz15PVJE91PRIefj
USkXgL6mIO518wtduMUConQGy3k4eKbFDtGSXzKAbxadIKQX3h0ZnKhNttnT
Q1ws4gEdM38oRtuWR4qYzd7gYKuVPZWMxwdAJSKXRo4dt0ozQIoL3qL82bMB
5EpKlt0N41/jRb4KE9J8qXqSC11R+shsoWL1WLH6Ky99Ye14yYmzJfj6IYqT
Sh6X0YbZieDZkbX2qIL2lRbEX2TcqGJ8flXTESAWePxgDpSIjf086Bd06iAP
fpyi/KHR1y/3/h4W09MzhSQdtmCSTODLXNt6Kg6mPmbePorD4ZWhqpgQe0ru
WF+DFH8mu5hf3Tlg0fFnp1mG+08QA//TcfIvhQ0A5P4/noSB1CgkH3HbZVNz
6eIBZKQDZNKhZZIsFRerXGar3EIJBk73fa7CgQy0QO5A/Bv+kSlGIXLFMaZS
X3my1p9jHJFZ6oTzR10fdIxbWEgijjqSWraWh1JqOak3ymcWoqos4QllRu47
OfWmQqKEOH8dThUARItGWI+d2ykMbNinBiCOwoGQa4Q7ZCwT6RE3UZ4xR7CW
f9J+3FOmgukAbXL4OZnyVhR6qgeNCYRReaamOqaGad2QSb3lWCnRj+jaXqsH
+qwUn5DVxx8PNn3efvzZ/dI7Lil9af0i5PwQkNqbovX04gsX/nvsmU4IIiUI
f0efPCCX91jUwzXmTsjdoG+yhinZL+tIa454w0HAiDO9FDPF74M7daQz5rP6
+cQXyhKPaIqO65srCqJC1gn+iv9CSPD6BKrW3EKsrY9aSMFd5f4FcGPFUU7+
ejhpfFdJ9SCarPlCyjefbroFsHwOPsgqXtIVU7kmI1CE4qAvH34XaWv5N3ki
QpGxqoSWDeOa85WNj6RUzWjcRzIgTXGzwdpRV0TlfSepKEH32Q/bc6WhdyCE
9XZqAKBC00MgMoQQrf5QxVq1xbHsXwpwYblEVU1f7fPHnkWdewkxB1KtHvUi
dTpl7M1RgynnVSWIHq2HNS61FGWaqFGe77TCx102qWWieFYCmpH9xRJh+DdB
z0Z74nRExN3AthXBEeD+pK5b29fPuRcxt54TLrBV+8AvZwwsAfajL2kQgx7i
CggOwotFXZecspZgbJsTEvkcWy1mwC/qw0WFUygTsGxvgwcCQ38kXDLufH1r
fGzFt2J8DAAztwzYZn21SmUhdtOkHGi9vX2WbqOeLiFO+0Jg4uzy5+rR0K0g
gYjusU/ELF5aSuHl6fHkGUJDVxqUIG/tXS90dDGToorUyayYDYvQ0XQ8YhOd
nX6H1GvoAg2lhh9ex5gKYXrUdPYSOmxNGewQPQ/m2VYt0/xM8ta6jrd+ihuv
sSty3vYCPP33ACtYq8QfBT6PGIOVMs5mywT6e2UoEePEIshMQOmIz4Grvbgi
z/YVptBML9NboFM5M3JoMFyJI7klqYuYQY2FDMzX4TPIzshlehsF4dKfYSHi
5bk5e5ZyMpKbrbBx76oDhWBJExqwc5N171QLJDJ0Qlz+LqtwunxvZi6gQjjl
LEE+FERqIe111VuiNqST0YlX5gMIrUwq5haTXdrb7/ge9/efuk0m/0Es5su9
RQwh5z1EmqWFbqF2g3h9bSM1ghDzA9pnnHO3/xIfq/S5mzkabHBGMRL5AvI0
3L9EzrqVO/DV/yO95ils+EO0IHe8jNyszg5We/ehkmbnUWQj/pv5n5y4wGMW
rWl31aFy+yXNdoOKpka3WD4Na7s1tJ+Ok9nIG6anWhfzln0k5T/sq5OLGjXK
I1KKQ3XsdO86ZwKez+NqQzVlqV7FpLmaUbSx3+ay5boaWCAbJfh1ExaN1xBC
EpAeXTyvfM0UFbcUtnr8RngcOdQ79a7jUZjqPdwGyphrvuvGn3+fIbCFWiJl
U1RkF3Xvqay/25QPQJIk5/CEIVlPwYqkzuVWKUphGe/jJTuROJXWYlW0gv+d
231WDudWBZCioynqbutRq9JIvzkiDR/UJymHUPM1nKNoGEQ6hU6gRP1SRkZ6
YmFEG9Xh2jtz1AwKq9lbfzwbnsU2hWtpxRviMaQNFeih3R47FtQCsf66qHwY
84KWPRoDZDLdStTUaJE8Wi8skCaiC4eEyWXtjDFsFQ/3C7tJA5zGRSf7nAMB
VlW9rdgehPboqHrrlMNfvuZwXEJfqMKa24SADC/lVy4JPpSuF+cyfTtbE7B+
ZJPCjEolftaGCFHshS0f8HTwnIEEioDWOFPxtr5Dh3Ebkgbx+dLRfpZ8A8uy
XTFG9M0LlClg2R9X/53ZPMD/l+/rFOO1q+E2YbgnXJDKmI0LeY4UZAluSeZA
ARn5tTymjEAJAIeeYmfqvDTJ3hn5qckxd4iRaOVb5af3lbirFKFAz4T5nCKa
/BFIdBzwKKmm3ZwQlktvqtF06dg/eZYJGvWkSEqr6UB99bIg1CBl6u7ozTO/
qY6F3xUmj5oD0rN4QsWJvhGJ9zFMpXqwD3SuoCPbmPn0cfUO6AUHhL48JNSk
xZNqM776GU6I+1+IGTrQ7lnkXuK/kKq70fucOZyZpw8dDrD+mqX1htjfW9eT
GjMy+EP62s89S3bgSwZlgQ0eoxfqgp8HwFgLbRzMtEhhIxhhQDq82pNZylCL
QNlu2xYjQ8SltKEUU/2a+E5z/Qc4WqROljuWbWRJvz1l7bVcsOYhNh85IMkK
PTHgoMZMiLVxTA6doHRMAuo2/+YA8sg+lUmZ6xekUs7WWVim/ZKZHit0fKjn
FA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Z1kxvUZ6A6pwKaxOdYs07NFMnLFQMgt2NVR5MKR5RKdJ8c9hslnSwQz63pqgbJulNL2IsMQbF1Uj0IhqVuqvHik8GKPJT0wra1hxuKAB80yrxPtVbyBlDdvuZxuBjXIgzc5B2XcslaeodZFtBeyMeUYfEN78Sx7u3lzsX2A4IXzLnEWV5U6gYlyO2tGw+1I67OKRfL/w6Pxg+cNr2D1Y/t3pkMof+6e8VFnEeyhkMUTcMzrB3RxvvjfgHb7Slw17/Ki7PjPE5vdHlztG4vxRFcAvuUjZa9lpbbOGG/Nb//QFOjjIxkt6c/dU9ktKLp5DGv4o6K0P/TcQxDCfdjsqiJgJLgbvvun0MbejATT9X+B3L1scKisgwPCYYwp4Wk5vuUmmRhZ2MMs9MkHpJmi+Ap1jyVRGWALOLO+9kF/7Hd8MKFNUSF+FPRTWPyhTd392UGtNIWSZQAqmgNCCya64FDgZq+FZN7B9VNcfpsIHghN9msyeu2JKIwfGywFQRwFXfjMeuX1MaeijMCLvbBGbyRwVHfuZljnGqyXjfCm5h2GFEuYGBOBcKsHcBCzknCNi6DBhFR/mHaGJFNsQnMi3dD5s0aRj9U/7WnZEM98UoKbwRwlLC4JgRqX0mBO0CPAySaYA/xBoDZqA6MBDRBOpBXZQdtbjnOgM8+/vabj9jcktOGnP0aHVpVMML0EjSfh7RMXuZML1i2zzrG4s2+ZggVaeVgirSszIubdyI6w41RIkvAlvJD4usGiokZhQJQ3BtmSsxtdBgMRqdKgUbEf8v7ceXXANq0njF/sbLogOdRgWNcqudyy4I3bniypvbyVoO0K1XEAj7T5MwrI0WK8+K2e/HR7xbWtZtaOTbe985Czf2Q1h71QOkOpncXtzKv5DXN2S8uBF336yeoXNfQA1Hm4t6/64wwS9IhcvcucGoOQpvaENuAb7nR7x/i7begaem3ivLr9Ep7Mlxrw7SY5/Rven1byFm9XHfXWOd6zdL1OKgS4CPJ1DUGibOVw8D+Id"
`endif