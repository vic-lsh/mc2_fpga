// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
umr3VYGtszGHj7AKTgQMkJxW/iPLwcl9lJ4OHn8r8E10aRLUoUTRVSvKtHNY
y/NOQYn3uVYPMKq4AwfUglYsHepByruUNevk67ryMExn5zfxxn43f9gxLsLR
GRNBg97BW0FnEsT6V18U4EU7QErRGBOt3ItpRbfnPC5R1yC/1u34aHvoovzm
DArLC9xELhVsBVsgRjZmKi5CAifLIAYaAng54wC5zVe7ietQx2dn+NLjiiao
7bIwCVByq+Vy00lQnHPLahowh2dmL+2lLQBciNOrbyYErhLHzpMFviiixR8K
OIN8/DzvHQPqOOUDl+u2L5XVf+olZalKxiUSbydA0g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kEWA0VOMQRc/idwfq0IWOPXNGlz4WgR4EpiiIINRxW4nfXaNX5DD5RoxXlS4
bkoSwfouEDJsGQq6DxSa1RdfYVyAFbXlI6r5ph3AUxiNa64FlYkZiJZmfF7j
QBF8JfNdSuDOKQKlP8z+D/nt/Z7ELQdf/bK7pvM5fVMwCG5LdbdzWX9zHKcd
HZsT0r4XXsB4mGOgwC8opyurYnf2JBqFifYeSyURVLa3rxxXyaHkkFGHSk3f
mxaYtLRq6ybjjdXLWHGuZ3w1ZJrorpI3jZOcozUD2Tim70w8biZyFtdDQkOd
z9rgD7A3HFoeSTRJ83e/pAa+IXq7nkQIB/SJpGlTLw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AYlAxkbnaOJW4XkCMRCIZeqS+jZ9JeOBbnHYEEJzmwy9vl7QzZgKqpxlvZrG
HHvGw3Qm+O91EwpP4p70V//uopFPt25QpHL64hYrctmsTD+i/qW9oE9k6MYk
U1NoG2tfD5IoFjVYOD9lBDcxTRZZCJqpF/kb9GgJqDxMxAW/ipul/ISFbIra
ITqHdZOAgzF5e3//PwxuAFxEIsevq6DNjuyFZEfC8tz17t3acrAs3e+841Wh
kYB8AdS0L3CbTJyzDQFKofUD+H6ODbsTkrgDa2sBGrgLymYasFCPtSLRAwEV
iJl8FJCYNpUeRc+pMonh5SnExmMHanSUWhkCtaLXcw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i1pLfAd3fHUqjsmg6TBRJuvldL+auN0j4Y0fQSaeO/66UPywx4KMefSh9akq
/oLKP+7z2Yd38t9WQ1tPLJsjEP7gw4xOF9hyJJAswA3it6zeV81o4pYsCdxY
5jprnFlI6Gh7jA4YGSStiu8dUxERK782XSitBLaaGNga28p2X1iwsRvBqLDB
VyWHChCNZ71fRcQFiv4eAe1uwSZrVhrq/c/ZeLbrB7JfTPyCBxMiASClMV9S
lymLXwor7PpQx8s7Z8sl6MkKVDV9mPo49Vsvpw9ueBmnRVjFLJ8MNGACmCJZ
ahLJ2N7W15/I6HKHVPjasiCw1WaXI39L8B5gyI99RQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LDUZYjoTtZUjEXfmhQz7MTCBrd+iB8BDLnisrBi5F80ZM7xDPKGEvCZmCjj6
ErqEVblSvDBUDE2fWC5mM5ojbhezu5t6JnX2gavIQsXWLnYoksRIvrPmDK9l
YFvksd7rOGJ+3I/iSyqFkQRKOUjyTXkzZ4iYzI/kRehKmC9DfSM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HWxpQXB0se9vop/LJrCviVA4Fj46guMbi2oxsn6O3DPxNIUjvMs8DlUU0qEy
KMIAZTGS/0JTcbX4mqfelWcOyHLE2PRobteob1PMZeKHCt2ThaeVBYHCN/2M
foIxWgxbswzYQSSqeVaG4R3jX1SoEI8eQ7ntZZyDNwHkqvFliBgliqQrvYI+
0JVQsQd2HluaLMFHjV5Y3cdK9aT27wu+JhZkkMOs4lOX7BiPP6ObZ/29cET8
Ev7hNFDhFDND+dRClTCDyIx2A0epZv7wutFsBUupjLDurdZLe6VsbTOlkMWx
/+yGrnhjEWGBzrk8SjUxl9M+zzy/UxGaOwv5Kr7HZWJljJlAXWgbHygN+12a
+jYetVPtZD8LsVXA4GoPXPtRq5SY2Pg6mScyrKeZL0LnJBqdVSUqe0WXfTCC
ns4xQL+kdD6G6XeAjFI/P4dTAHoasppX7OSrzsK/3gxl2xrZmz/T6XF/NT5h
1sVBLTLiTqD3creyk5DvGzyvA/YZKuTK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jmMtHAPCSlq4QTdfIUfjcf1/Fg0hq+XLDlBUHadFs/rDGKefpirPqKAOsHhP
rtPoW+1IUYs8Cjq3gnEzySUs8krhh1DQd0uwYOHFuq+De+H0Eg/HdYofP6lW
dyLQlyJ4lt8WyJqej8arK0nQMGZtoTzpD3ZeiJudPJ44vjWkju4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pWL4/L5gUbaebT02pzkssYLG6t+LRegOavi6RcYVIKgyTwZAReG22iBYmG3t
1bD3uKUu1tnE1vutpxyacHa55HUQ+z/tMIet2alunyzfUDcbcfRZJpsa3PoB
b/4CYv85p5eoaLypr9SoRX2eDKRVxZoZiUSI6W1LnQ0BzTD7RlA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 65472)
`pragma protect data_block
79r+lyvOWTdfyUQZMN+Tv5cDu2KDZ/VEsRZ7B5xkPDG6W6JEDFydiBRxrqRg
9Z/wWurhSMhzmifTFb+iDzw7mwTanK+hzB5HpSk7I7oH3wHP+rPr/ux0m6e1
xS25M3FaqzElliUjOsvITzhcJA1W7LWVYM1Nf/yKtoCAN56tlUyxGiIcz3jP
ueBoTQ+ENmVnMg/PQzBklyT382YGgrOZgDngRQtYoBBnNBEU+kwQe1+1JHhy
eCiTPa8uUalZwuiN2jio73VFLWLftPqaNTIWldVS5J/P9BZmIbcjyIRc5NFO
SgwcJe2jXrhB90m8jEX4PnsYHQ84LtJl5lpnAXfzcgigfk3s+h52Kn+KXz0C
BmO49fmI6vGZJqxOXK1N2gMmqmnPBfrpnxwrrlQo74prg6GxTrVb7ztAOw6T
FDMbJpMpqboWiv/eOpR19Mq8QpNrMD2Aw4Bk5bfVqbXS2bqDt5BmuX2C5sZa
Ipq0PePmIKASnTvTkA5jbn1yjUh1AoVQo3sUNM+bTaDZ+wuGa3tW0VgGDaHB
jpGmD1veiHuXyO5yHLQxvJQHbpsPg3NAhndeVp4MIyvnux4r1oSIH38SKzrD
PTrNpYqdfKvBM2QkD017g2k2g870k3yklN/SxCSg5YUi5lQB0Etf0B1Qq+Np
ueEw76JJau0jvUHDmjrLZgMpvy0kYuXRKHAPZZP4x4tBHlD5D1bF4WRD4vy8
XUx6X2mYIh+nBj0ic7nEnG71uQV0o34UsolrQEjtMaOoWQlG9l9Ev4Lkp/TS
2PDxF6IzjrrpQ7Of4QCpbUtzrsLC2Da9dt+buDoR8ra8CmnQ3BkcbFusUWVd
bSAHFWYcKI/mljgINmXUanCxfdnpuxam8BItZEIdnyvCTG324Ej+VNAIx436
oXP/xqkVaWJd5sewe+m8Ug+zOCAgzmQjutfrRDso2tIuBFtTOAiLFSMI+497
rDOh0XZiwqLoePtBbSHpLj3J93LktEpaEkS64Fv0UOqvDiFi+iRptK8htX0P
ghs6UALNA2iMlcwVDm0LjNEr3PEj/iRETbax48XTQXtmNYJecfAxPCpCYNS6
bFcmsjBU/bocaGjvfODL8lEmyKqJZzsk6sTTRskRqUFgyakqdgOPLOJf4OSi
xg2ZckVYWRYDsl9iWarQVBha9siAyVMZ0ITKtjKLzDSuPlYCawSS34xtj4Pi
lYY6T2QNdgROs3v8Idq+QhXn3oO6j6VPgRZzBxJGCyqfjR5t4kEoROPYmQgQ
sAumRCBlXm6PoLO1z+mpi1pGV8lUj8F3+hEwQ8OaYMuki8OUzd7MjYggGmMa
yiC3Uo7DHeft6NRNcKyLMrK3D8sR99WFT7LqKahpjsbrVPCKh5lY8OlogC3f
2DWBJv4cHKWF9GR+PupApVKX83LtS9kLlixRqMtziz5SL8rNXvi22C92QsaF
pBWsol1ozLIOB0kQOHRrWihusOfL7UcgLffh4kH2CE8Aum5Gj3prRBn2S0+h
HL3DU3ZrnaPRzxywwqndBs9B073guivpxU0Lf5e3EkYxH5I4RhM62GL4UuiY
I8zAD4Zf2XrEny/LfqOleM24iS1YShtxJdtWGcmerS2JxKNQ6YCGOq8SvYDe
a2cyPw/mgVoUbpGqAicwqTDSS5XHTf/qvF7Dax+JYXgTwymKneI43gB5EIh4
8+ES4sfYcT+fluzx2QhAQ0h1zcoDlI8HFOfJI/9hRaY3Bd2V3qKGPo4n1s7u
+26PDkEBbXfNN5490CilZLtjuvX6cFfkwZhxlacUIIuq+ZxEfCaP6YSdgP/2
XMSd4ddGVbyghfDTfDNbnwXnrCJo9coTl/ryG/yAWWS/3FoHjQTqdQU3ni0J
Z4/wtrpaSKkGvb6ptX6N2q5clbzIT+L7skft+dcJchsfwVebQYOtsXrgwMHg
+zE6dEKsgXuCsvfEYk9xRIIgmiikyj/QXLxU57LlrmRLcOVNhRJfBYqR1J1R
tCKD3InZCvhDMoppvFgN20iQolCRYEl8+bdWeAw/1qnJoUm/SdYfZuqdOmRZ
OHtkk5puUMUTqw1Iizg4ZCRKBb3hX32TTCZZdlVjR0Os32zmItd5YnksGj/x
atSoxLODH7BTP6JZ9GFXAwEFQyAQMN0GLJRig5outZXxiK+f7c1wn9apIPT0
C5p/yOErnuBGoUMMd9ruUtCYPJQQVlK2tJ3nJbZkxcnik9aqNzbtHRfDNLwy
559prcozfWrLOOiG6iFmMITqKMGZ4kqb9sPeAUpkuWCmvcIEg/8aLm1nlGpd
qztgy2hmD3G7OwXcWLWRsQzm44X4y3TtHfep4MJcKZ+tLFlxtm0fFz+zDLqO
YQtcLG5SY9QS5BvrjZiij/BGKJfRTQW3bJpxb37hS4DhzzwVlSQ/DBmg+Yx9
zLxEgLNzDmEq0o8tZ+Y/IcWsHTeOSqsh9ECj8ua5rA2iW8q98s/O8T/DfR8I
x2jU+Mcy3l/e+1fCYifroavdN0vN+H47FQBFlNOsbslAl0E4lvPJJnj6jdek
MY1BVMugvTs54ECA3SsqtoT4zAKrWbfmNPWGCbCaPifqeU4iKDLL1+5joBS3
IaoUo7Gt/1oPdOViRWMJs9uY89yBG7pT1w8hb5dv86RwXBC3wvktSC98IM6Y
aEVSOb5GK99c5K/gCbm0scFbGYMdzFEez2fVfShxa9jUTXT3L5JYDfnOzanF
F9ZXqNJ18NN+3lGTU7wW19RDasWcOhsr9yvIz0UywEY4OBPap9rL7TLmcCdb
80elwN7NUv04cpcG6f143ZkrjcGNEoUL3i/MZn08OrKWf2WvXUN6ESE3NZvR
1Hwl8QRSdoZPTsJy9enCE2oQ743VVmSADqQZ3LWGQD02rW4mpIHg2SPtcVB+
9MpiH2/8wFyKT9DU/mT1Iy318ExHN/JLW5RU7fS/mwJCEBmUYtIfyQEHCWMM
ZgkNRFSit6Yi2Ih/oASCCBV8rckSrwg+8JOQNz/f3Rlni1ewBCeyUscD1r8z
2nGBuF+ii4pFziBsEP42aUbA9zaJ+OEez2lbbV26vq1eDByRqe7aIK8xZYkI
GAUGqyKUcSWin3mTG+Ka8KxtdRSjasidlaabOrRb5D8zfe2pEbuy1JS6aqD0
I9lH021AKEkGCwdZBOzFEWVcTDTDCcZHHxq/oRpYZKo1y6/lPlmldip1DJJO
u749CyN7fIJcXpb8MFaMM/bq2lUCA97ZLflBjxEEoQC1DSrAKjIOyup/MuG6
20FcamgLaE7Vn4iJXnKTHDlOTJwwnQmhPug5xT/t4WQ6M8YWLYZ/EmrLFaPZ
5kL09u5m3RTqszkxZPN4E+W6z/atRUBcOm5+l6eKtxIg03IMNG/AbmCbB/gL
TWc6l3gsibw+fN+KTnfmBOFBTkSOFBhwel2ESGxr5N/a9lKBolAszErZWjfJ
neUkU9cAsvyvy4Y/TBrsZtNImBZImrUlhPJGfZHqSaVZw9cgHoD/pn4xQFER
HcOc2MCy/C1A8EnmE1m/DLVJheXlkdq+V6wbgazIm3kPaVlKJKwhF+WptV3Z
dfcA0c8xHyhTlEqtxr6mE4wvP+xi7MM2euK04OihKtoD6bOFuy9eUdXdhvBO
hIeeOv5NFjUylNOBIBeDQQQVtm8cNg2Wg8PE6t6bKg/RxnDMjL0WoskqFSS+
b0Lfj61JGm/xM5aDENrQW6ZN/kczzv8IqYii3JaLFjfUsa9k9mRzVgWTOQ2/
dPjEyVE+7ObnbTGWK9Kxxmhxf/pSxMCWp3dbPvrZVCOeWLs88DceZeEZmMV+
Pv5Vjwhhgmr6pqiI5ihMHVEdtfr/XN+6pk4H9D77pWHlEwrSuIPIMdhRBzNG
DEh/XfQhyE3URjzgQQg5skKcSgPU44S+YgPgPhX6NFzQrLC5puVlvV3OH+Rf
hv2oflq93JJUOog6IU2Ry+OyoDO91wFmADq6/FCaim/llbVSzgVvX8BxFKrf
OE9zAWwrqh0CF3y4b3rqRbli6/pGjux8iwnhfvS1m7dZQzE48XA+4+g7es5h
l8fY8fmoFvD2u8fnj8hlNBGMyl/KwWgC+QQ+KH+V08H6eSGgm5X27mVNIrzU
J8p4lamkHmL4rAoskfEPm+ks8xlrD2PeqfA1nkGLo4/ZoR01DhzoDrHvi9sv
4b/qGvcjWiLi+mUdx31AEV3Ks74QVX9JTUkTuT73aUKbGw0dsAUViNVoBrgC
Mnmv6GOrLLhJaPzb3xUxini3Moc5E/IScSXyMc0ARj1jOYzMJKhJ8PxYKokC
gGO9Pi9IsYUizqwzWcjP6Ma6MhFxqciGBoAjF5TlKkkWmlkJCZsEGnl3oON+
k7jesAPiLc5U1/iyCk4W3aCDc0FrOoBDw4rqfLLfYqvxZEZwh7x0bb/n/dzv
hV5Gl45dx0urui1LSewodt7+4Vrz89RFQEb+7jBOm8lw+KKgBr4Iy74STsPT
6DjP93irZvL43YcM6GLzfdwiWTQKk8CB0zdEgc7ylYzlu/t5MUVLbxHvOwwT
LND9LH3HxEBMY9qO7ghgC3pKJUh8Pbz1GbSiqsGB5QL6REozvmAGJNbtaVgb
Im9fYRB6QCr0bul0dq33ESK+LJn6tKnfywUBR2q7rOvJgewTyTTdt/fSXEV7
a9sIKmeogk9MwADp/cGQI+M5BgUtYPlneViq4OoRcb48o8OerZyx3X74b+0k
zAFcNsWJmVQKYnxq497XM2t20pTvrp/9vk90h9n6hiKl40cTXG+H/Z4qr52r
OzrPDrwA1Nr6u0LgQKW5bmhovQ2JXHfckTxXhB15FFLUlIPqrgEJrSQ6Vg4R
uSyZr3iFxpTD6Jez3dchONyigJhXUWARM7Go167z4NevjTloV2ia6DvrHuiA
QL0UTZJ/T1nmjg54k45fVxnqds4Er0QYUiVjyS/QZ4TnrMO9seQLYnaDAbJX
dJabL9asoCS6mnaZPBWQe4bJ/X1yrLcJF7Gq80vUSwtyLbh0pHITWSSQbRKI
kV0aEruwrLgVUTbGppdP6A1F9C6bFhuDJo5O7aU8kCPDHuti88KArNo5Qge1
ost+yj9iZaIEkoUM1lpd1TIwMLI3PWyfsHnXkz480/2QHE2SbrOldIg+sTvf
RQRpbxhofbksz++4tmE/0eBpjI1zewx4np+aRbqzapIyzEb4k+X5DJw4n2au
UGLzy1NFgOcm4S1uSOg0Ok/nt/7y5kEPQmLZ4IrxF+zh+UeJNSqO81YJuz/E
0wafByPQ//HawlQBQdQ3lcmOrkxwCHZEyAn0cUaAxQBkzj0mCjAyzQQf9Tbj
7zfoZwNY26+AmZoZncylWrCQEcyHMU1aKPPAZaptf3CacdMVfvrg2ytDv9dN
QYZDX6g3IOjnKqFLEhZQkpeVQ6Pm/n1tfNAbFIbJC6cuHGUl5Oq50FYI+UGw
cZjFUGxZBqr5naIsTijDwoChOxavBJp8jbeelWON/T29HbXsSqE6xbHGlluR
2dSYHjSRR8rRX2RfH8e8kg+6BJB+Jk1q+D5IhMbtxWaTkpPKrtWrrmN289cs
LC97vQ8AM+gPmrWBT8hG/nlEgzs49rHJhpyJNYNufgQq6pll2JJ4likzXrnN
LA9MPu1vJo6nTv3nPOjN8/tyg6j+U33CUNBIs+cqzBtKZUTS5pwPmARnp5u0
HG/4HSpHYqW+jE6KMyMKCvfTKMlV6r6okJT10/osWUbhBHAPEOeokDQ4q8PI
AEmUxlADS+W5SAvifQ6fGzd6VO3Vp26dVLx4fQOyJPJ8wh/QEqpZZFMR/G7p
tW0GVNaFh9yQ1di9E1TptjzXaCwNzaX6ADATpMMSDanlqIxJROMClM/byWvQ
qD7L7M16BPIfLFi7chji4B+h+IdszVWd53Z7UuBtGef+wmacBpb1fo8KfXZV
vD0G13eMtf/VT1oHLY35P72CJCtXoyW4UvlCu+nnZiBm63+/lctR5ePjh43N
AQ/BG+EWO7Xvv52I83gyi5Oj8lgiWQ6c/BSsNNamWaWo4CCD8yZtTBraAKuI
zTokQTP64NycRluJwL6JPjmh/Ty20SU+Lv+IxMQpUu0Ymt4DivsX1H3dbRW3
27fZ1jtY3G5wqtFVrT3AV2G7nUNDZB2wi1+KR5Yow/Be66kRpMvUc0DIdsnM
Y/3GBYQ8pOUU6TxCwUNQiNRcO8kexPXxpS5TDHFNQfieA9u1P+u9wSAMWgQx
cTT/CzXETMOsBP8GO/GW7TDBsLLLDyQajmQUYnjQgfpo7ld++fsKibNq76RK
pS2ci0mMLKvhKvUWc0R5cM1za6OjJW++Igti8bLjHgsaeTKbrBoVU2bmAfdU
ZH49OR79gmbyWTcMtkONPZi5Rtzu41OhEF8ue5WMuhXPtyYEGzg7qNc82g2i
0UHKeBW/fOsF91uiHAurKU3b5BS6Lii8hIBwHjGMl/YEEPQIZHV7xgF+Pmaz
rCg32qMcpahhWf4NVHQD3hmuEbycjUkPpt485UodDi8Lny7k6BPBMXLacNrf
2l1Vz+8h2cLf/NpLMUDljIpJYouK1YpZCOTxPd2Bu19ce9UeYw1CQyYQ0eRl
/FBVK82rik+CXf4qMvntFodviXbi3sgx9eMUl2WmZ1MXeP8YerWn/QjnvU8Z
AbqpFVk5RYuin/FK8kDgKsqWfJiRejCp5l7GamURMzWZU7UxWmsQhv/SiKlg
8585wPI/tmnhyTZxs976me+lwtSR9XIsP7xPfYMunIxADc7utCEYTcWFytJt
AJGyK05UTwt19aj1Y93jPZU15orAiR492leQA5LkX44i0gllXxdtCwJRVoBs
6FAo9UszUL2GJGkGTx3UONXgch7qznhAw9p2QEOVxPEow18iGwmvTl94qdWf
wFiI+7qjdZXid3uIKRk8uioRYJVuEB9Dzr53uapw20+7vC1P3anAiwwhfCWd
8DKdRXZniZP+UjNpthciIbhmJfXD3ru0JeDtm1IKiHPkSwiMwCrh02TsYFi/
X4mB2sMtnsjEbSSMTWA1nYU3YR6MXkz81NY3DYn9U0l5S8o63J6OscMfO28l
7qh+Hx4cn8rwUFeUKC1D1DdUOOBpDm//SB9cIu577Uw9EVM5l2nhDfFvi88X
12dzEVeP9wdF6yQLr7JQdqk07PiweZQxWiWOt82lwlaWcInLc9A0ArLY/FXK
F/BxVUHBHqZ8jMa/318khXJb3rNcgMygCMCNqwQXzyYZzdVv6UjwvY1vg1zv
JZNstJ4cfuGQoAp6FQZZzqXxfnVv2v40zpyZpi6k387ShN37NCPX1ADZXe8Y
GJ/FHdamCM9xWyXcjXkinJWgrXhpea2dKEJwh2WgV/qGyI4/8uVpPndssLNv
6nZMQV0LVafQ9UKc+0Dx58kZ4Fn2+S5O7eVUFdLN6yZZuuCBbZXLIDcz7wi5
swoE7N+wx2KfVknD10de/M9pezjWRB0+BsUZ6VRQly9fKH4tFhxRstuBiHWO
vHJ+OcKprsYnEK5yBv9PAo9siCgaIyvAoZqoh8V0VfxkxuM0XSf3Y5365GHE
IoX+QFG7tHDtPiVrjdS8rrPD+8if4uhPtMlG/+TIhmX8rO4CELouW5TEqj0E
mBTIYNz7FuCJIbghZL/JVouV6BRvNKNNM+4RfXM4JPb/MFvk/JNOCFCma6fO
QO4DNefSgvCjBGX3XGCELu7P6lznFMzWXrJBebbNkxgRbgsMmkZtvnK5gKgG
PvTRsJf4t2lqUfBztALMnE7EUtarnRFR5d6Cz972XVoLQkG62n3H71/t59S4
Kvnjzyb1u6b+44za6o1+8RqvwgDWbjtZrOYl4jNyJrH7tMHOWKy101m8qWvR
L16djA1pgH1eZyzs9OfmaJZg2zhDuuC44tpsG7d1vrE7kq0K+QTxD7zF90OI
PlaKgXARvd05tZ/Jg7+BXF2aQNRPtdb0i7V1eyJciBcuoanUADn62+RwoO+T
EJkkC1CjOcobtmZqjxs0SYibJFLPb6XyWxhBg8tkGXhwSHWMoIMGUHURBCYK
KzyMRW6I33PSdDJKarKcLqX7pKZ74ycnmaa1VQSjoQL/PL3DmmVdosISQUoY
Oe1yftz7XXRF88YHMsrAtyasZvg5w5Ka1TMcggdqP6BTP3vP92I62FmRONZB
OzgW2vNcHbQx8bSNaVLggCprW62p80XhvTr7+TRKB4X4ta5bsDKdNFWtsEK7
Obih+en62eavLbi0AhXTYMDRvbjVdPaEfMjfibowzKNvgvXPOZllbNpd0kw3
IlrSDYfn6JhEa3/rJH55Tms3pu297ddWVEJNdg6D2u1yQ1qykNBAVnoWUt3G
Be/+tDsNFDP8evzMVJfW7fgyQxFTZjKl40ND9Ii7Takld5E/ReeybW4TezfV
uXcb34apyObDVWJU94h0iMqBi0WEAIpu2JCa0MqmClJ7VucMhbiEoUQyUCu/
t7qjXt7XBkRoBxapwWJAPmzkI1Pnh7yTyMFSWLZoGuERucKH60Q4sHfEqSIP
pO3iFWh7MfnAg0VDaMGI6UixP2Fev1hpZ55eBauzLxhkY1VvWGI9IDB0hWi5
rRxmmJwJ3rISdoGNitWWVHEpOIHhTzzVdUQFQAAaLrCi5K2rIUl+F9RgTV05
i+NwaBkoYrDPdRoqdjQcwKhwMpmCVN3f6HrdldJMMxChVy4TAiabR8kJKEB6
gvicbc5BcBAZQknWLRRid3KV5TjnqUya+GHJlBuj4Ezb9OFlx5zn4z3FbBg5
6HmE9U0XywGWpB2R68ZIyu36dbRFu/dQKKH+wtTaeDe7+AW5TRX3Wb6ljLKU
5b+J8NAiWLcGA93ukJJNX1YJqsdcrJGZdqAFzlsoFRS3IQc4Qh7drQIIoWU+
chQ2PFu3ERUN4eC2OeqVUkxHhW8eFn9fE/LV1mR0CPI8dfUD/MXxmCJX161V
/QHUlVTLA4+cUazdc+QT6jhqCQNnbMFDk5SrQs4VfKdmkGVLrkgdE+ZTpLk5
3jv23EwKGOTgj6q7r0EciqvK0DsX9lsnAvGMWMoYAMsqPQtCryZPLRB0TTVt
wZ1cvQmuyVfeAW+vgApKJZPqdY/YggK6erh81CUCV9svtJhSg8TiXb+IlvN2
k3u+7u7XZUg+SzSVYjcDWahc80hUcVKSCgWljste8ByJtVCs7JluEZQzWD1Y
FZTR8fjsBdaqtQbr0jqOfPvG+BwCdTZcYozjmDPMoGzSsQRG7vsIO1soA6lA
Pa1b3vKXPu//es11FVV+6gHwSF/Q0LGgzejLoYkMWOKoG2snTJodSmNyTyKu
uGCSMbuOlwjAqAknDct3QbD55cagoK1xUf3xpK3E4scmxxnKXxzOP9eAakMU
KXsdpXxibWOqOkLLJYK6rSpn+FrRUF3l0BC+hwO4z8NDiylOXlZSVv3Oyzaz
cdU4C9poSHMzlZvZC3RKRbjVwP6SDiGInv6w0zIfR8Q+wCwx3qYo5EMdbpr7
pmlJLER+VZXYve/u6IvNPteLSyM7RgkaeeM+WUOC7gBLOy/esjD5mTjBDKI/
Tn6rK/ErykLPMArs02HdVIQYQBL9MRZouYswEvQKl2oBGv2t02MP/D5Grsn1
JE5ShXCJOQevBOuJGC6/unisHXEtKGKyU1hwKOCiDUKjOIBcUGZQl8pJgi85
iRQmpGGCUSfyafzvoMaQXyIFKhBlMJqGiZt/ubkRZObfzozqWIMj2A2XvURA
tpzu7GlpU3s0Dz4fIQBEX3ZqksQL1GkcMi7OZywHH/1Hss8pLoD+WVMCPJDT
t4Fxel8cQ2umE7aStf42S8RIARHEyM4kLpOyrLGZgOUCNLvJWgtNvoWambKU
mazyrxzBYItQ1JOJHasfVowKlDJFZo880IFz/3j5tKq3Ci6Dx50n+7Z65QmE
xTMacpJOH+w4tprvUxkun2mOL4Os84NxuVFSg7/fl1+EyDaGowgOcpno95YB
Pz++VBqVa+9vxoZeZ4YcgofyblidksENmUQrUsPg0qyMBj//Ndtk0CoRQ9bu
kw/COu20ntDqqGJ1kfVOnBZl6Taf+fOyKE0ht36XtKBfaI9KZKf1bWaYV3Hv
SQHPAjrXzerLKYDFu91G+sAk1vOFLXIMKPcb6gwCUyQoAekasfxIkzUHoeaV
fcQetwlqzg9pOnmjp8qqo4n1ky+czhoNnfJWYbmCkGt1BgRPzWalXuL7WtR3
1PSqAKDlj8gYiGOl+RQBOT2PNjPpC7qxBg9qahV5VP+L+lcvcbbOP8f6hNjS
49m5kRkD3CC7CZddVJheaU2kAp1dyJAPZqIbcDQYvcZgvvEmU1B71QtI0t96
c/snfl8KtQlNd0wMG09GnpTz7JY1cMH7DkvHPEKeN/HifUpH05qJefUWwvKh
szQGn9PoueBnz3tZUlfnstTaVkGMyJ4sx5qLpvQzuLglU3wfkC/qMI+l1Mtb
quaq7rKjqrtR3CrMiCT+y81FltOEUUujWt90UKFNBFzQFrhuwvxNkJGwSQ+e
dFpQcbnaDHNiXcLeM7QqzDoOVcPQXJjPjCNkpZGP6WfxeOm5vSZG4Pphd+PG
37jEFzHsanLdyWOCTnadve7w1DbEeKsmBrG4Zl4R3gK4X9qJ3ZOr/t+gJyQd
dO8NmhDkkmIfSKZ8UOzStZokqV3fv+ZKNtEaZy+CkSsnf2RzWutGRPzGPG1w
cEnV4mOHhBdbRYuAZdn0aRTewyiobqUgZvZ+PLF+l8Obo+T3HDXwpE96e3Kc
R7B72+7V0fEaor7axaB2xHoaaOxUGVdHfPsxm97rwdxluSyR8QH0rQXdlr25
GVr0dbUgS2N3KO4up+iQ9iOIx/msE+gyEQg/E2cjUlOhYn94zhqCIkn5qcOP
tynzg+9vQgURBS8R9RaSDHetr5+pVevshkSIZT0Eyhp7+8dcEEy2UGiosR3z
opqQ/BxyYKwAHtHLdrybQ9CGcDng428gqEkMMMdEZ2Pn+D04/hQqEL7/LQUa
hnCQQgju5FNy68PfBuOFxoDMv/6DN9uMcQu6Wb+qxrSSYDqoJp+8ioD6Usi7
UBZe0MpFwkWwPm50oZ8BpW66UQkjc/+la3q+v/TJUws85iWrao+v1KLfAVS6
SEqo6fQTJ/rmHD7uUC4zLd5j35GJphWRD7jARictlrXalahZyfcPFc6L2+p3
iMKpeYIxxFj0547NQ2rmRGmo6lyrSrdEQmq3TuhnRI0QDOYqVirfF01a3xzF
QX8/eCaQFtPw9NrPUbj7VPgiQKgn0ZN4XV4zrrb2Y2Uoi2wrgn/b1W1aOOCP
Vjx+wncBajbw36aOGRj0+CW94yGHgnv704GJ1M4FuKS1m/EqoiGBkUFOmTEf
ncfm761irOA4YqPvYDBqwgPzBrfWnGg3k26ccKcHIZHGr2fNx0Tk3LcxyJy9
yQ/lHfSEInnrhRp06N+if3445okXllPlbZJ/6fhfaHUWZBU3G6MJWLsctk5j
YnCNDoZfVF4P1IzBcdo6JfWuK9mpr7d4muVfudgJNdFLCc9Q4VYEQ+icTNkX
V2NP4V/L/1UTsJl5tqosl+uTwkBbrkBW7L3jT3/7eDnPWRB+h9rcoiWaynxt
uPalAlpVmggM4BpwNXQB6JAB/mylCkxbFgs1TKu0z9uwT/1nvHHYC+Tam/qF
+HUyBC7XOHJbzGehrKxHQHH77Syk5Mpt0EFnRgMZqv2TUMB84qfi28FVxyqB
bSlWo3O0hgw/IXus8DUTfqjYLN3jH6LdBrdjcuX8jKaODNKGbRijUdb5Nxfc
0r5g4kkBuTvBIHBgtt5F3XgZ639iIGU9HjfPGb6SZ9mVtLJbqfJ5LlWEKqM6
V3/gsBoYXjvpSnURIYrnPdcliTcog6nzHUOZQFkxBdFyBKUPxZ7MC0wOXgR+
2EPMs1ITpAY4BREOCBv+BkXRiPSZkJd6z3wpzydxVh/aZAVvmaBThHyYL6SL
UYjax2RMyohvgad8h+8s9qeM9w6yDGMK9j2Ts8nOcIeq+VwdJB15dRKj9QE+
gUPhyI3cpXXP6ecElLht2YJxSpXxjlF86LZ1+gJrmtiVRUgPk1bIxYaxw2CV
tNUjUnLHcD99cnfIANjWyWuvaXLBljvZOQWvPcPqiZe1yHKkpgafu8GMjpXn
5E905f7JZ7Wezs2NOqCo7z7hg/c1aRWbiPU8dH3cCFWGzpi5U6wR1p9obzla
JgP8SzoyoQiHwvXR4V9TIqOFh7p59KRUwwZGkQ4r2CQmmU/I6nuu7HdZbMZU
7c4ESO2dCGO+yZ/PdTZJ6IqGqa6NQ3EXnATjd/xklYs3zaT4+DY1Z6lRjgOx
+a5Un+UX77esSpQInc/CoF9irJKSuslU6uKVZVAibS6bFDdY5A1n0FBDRNwL
lZLFsOAV3NB5N8dhuTebjN4Cl/AcMysrVdA69T9cl7fpX3xanq1qcAAiUnzC
Ey07NuMae2n2WeKL+dEFzub4Y0P4IFywPZycBdz4UmVqnus4c42hbDmQMoY8
6q26fLiNOVdlorWFjMWp5aXZN6oEnyO/h9uD8y3bbLPGg9eB9ygtsNBCOkSy
fSkmyowhKisYsnwLfs0GU5gWu6qOsSJMrKp/YwKLdNpb7s06N8uXXcDZeNK3
8n4pmyUGIWcTetYbJyUkHYAHymtJoGdQz77uhBGmh63VUP3l7Let3HfnMGnS
NIEaETfSMppN95bhd85rUXOtWolgtjUHVyXOIBLGum9DeqXTit6WDQS5zFxk
tVjmQLlJkfWF881U6Ow1Ib6OlsLUOkuaP8/T6w7h2DFhkn52YGjY/CPnoxny
fGAt7GUuYrLumhzLOoVfyIsjON37qDYDryMKb/TYYphRVk0+wutxLBjaGL+B
YAW8ZaN9GcZ594Z5ZOl12kV2s+AZkVKezPsVN3+rLqRlbFzqDXUGG9UEKKMS
UbbtVvo+8J5t5nrco4Fn6cX+jdmsvb1SliM/PQ5bXBM4biU/ndA1tCvemBCR
JuhjhjCtaICHpa2PInSdUWW6xY1ITKfkwHzQSjojg2fv6yPnyTDLdNkbf+/w
O/tzoiaG/xrbl9VtX/sNv6XoJGmBaFuSsAkcpecditmQyvc2PuFyziffGxPs
D1vavIgO0mjjHbSsB0pW3XxJzpfpP9GqP3m4dMpnGdoNbfZxSdGxaPdhVV++
F50nfQ+JS0zAOARt9ghEEAxgmkmzYjk1HVUiLbTQS/0b8WtX1uemj2BGtqb4
GA789wpzo9luwfHpAAuTfOM9OcYsuBLCLPoRreJTIbRjEbAWUOFC7gTNBVAW
/NJ662cf7RONgsC9D9gYiTbDW96co1MEDtTqwWDfnV4Yl8pQ/JnXqiPhEKK9
90KOie6pfWS2rwmmCV4XX9gXxetI/LQx8vOBj2SMLDtHoqLNemZ4WFYmumPk
jH0bJr9cSNtp/vGqlc4PKGoiwaJsqbwz1fRiWYKgHXNaRdMc3cByheJ2VKLb
qSBeB7XpD93wUtic7u8uaydlY/iFV4y7h93nMBMHdc7zmAUYGVlWQCuAB5Y+
QSCXAwdFRHGDzERFN+BWJOUkgfq1gawK0sypb+yigGyOj847csdA/yTiyK4I
DUcmJymZ/4avdq2xYOBzmOC8WTZ4GZLeQPIwcFsgv2msn0iJJDa7CAEg83Ed
QCk34n47doFBQ9kvcLXqfLaifWuPtDyLTXG1i3UsJtLNnjtOV+qoIf8fbQMU
8zPT6b6OIAz2jqSEeI4mP4XrdsVskkuITVO1/B4cLabzyHTagcnvLEd1Catx
9kY7Q9vA4CZc8KLZXNZCWOPv21RshG7k9yd277vkxaRIezib3jhuhlF1jVpB
BcNJ0QR+Np7gncr1ZNaM9HHkTsa0r/lWLLc83t/XikQ9M2Gj42rW+0nI4B7Y
mrXhEszZv9hc8KkUVmFz6zFO0y6KCmVDJ5pI9OZkQ4c34De9jJsGuFcB8wGX
laKWIrfCoPa+4pJK6CW66R5G5mnosbC2Wyge67AmHnfZMa1DwoCojfmaPiUv
/XSh4ttniTfwlhihPlujQ1MavLsjEnV7cE9jsMRIpua/JuuVpc21q7wUFs4o
ZTwx2wP2Ifj+RcCr+3tfRab95keltCAOHrDzl0X5xUeVpcjPUj3/JTx30JkA
qDpd3qq04aTpAtsqYk9wXrvWZAy0vDMFn1uogoPuBWqFox6fk3KaZ+G4/muP
J5RSOBgEAk9dZ2xGZSqRBKWL7tcW8b9BwXOwDTXasEF/6zD1nKYM1veQWGEb
q06KnBHGN3D/R7IhIAe8iEUCvulfHhsbRhgrq6Ty10nDWfiJ1rMfWVFMiFM1
58vFrjNO6lxtwLl16/KzHGvsN57knjRsZ9a8s7qF6E+UVg7hQ9LCIgFGjhZd
4ce+JZJ4Myt6QQ7OnOVUaL/x/adjGpj/XBskGnJVGArYFAcCd92PoIfS4LX+
42U2dFJkHt7KM+GfvkgnFNErwuPS0wCqfQ2QVV/b++7VVCjs+RPmRF23DmeO
Gfyz0M2keoxCS/1Mjr34Rd+w//vHHEIXNRvj39IAf4n1sZ/P78D8lOpptmWN
FD99dZVQXC9n/8uXrfW0V3vgWiuqcNWNhz0d9V3EcFgfGh7C96d57a/BcFRb
q1DPG/2ZM1eh/1Y8EEFOnK0HneKYkt4MdnPOXn98JrIKtBm0ufkUKqfIVDCG
bSj2x7DpvHjInpZUqHgVfl+YRg2H6Hzrnd1XhHNIv40belfYV2PwkX6ee5Ty
SS9dsKD8WBxOLAX2C5mH9UJZJ6VWUbLdRmzXthJuxuYCY5fV1ocdrOXGXKg7
tlJ+NSQsxGqWZuFPqHiflj3foJVzShDeafMc5Xi4bBiSlTpkqQqKhbL5wPnt
vmg7jztkhX4PPzPNYv0/w35nEmLGxPbzZaOC/pmnAf4p0ExQCYpn8DSTXoyP
TOfHzzZBDqhVQGC3dLNXJpTl+soeOmRntKfCAeJ67p3MJTtUVFliYeeqMRRf
/N1C6G75VShBUCcfFBac4XxLaR5EohuynDfKyOGQvlEOV8xyS+pAQMd/uzi1
52chie8dx/T/0VRt5HDfXq2Vk3R8Yox19jZRZD2Tu73q+C9W9G/S7cLQRb0y
9tIpGLJ89jDkSK8gOeBXGqkRv4EHegGjuqtfdJm0OxWpYCNV/6Ywssscikiy
TVmex621UeSXZJlYai8lfoIJ/pYKEflBtz6890SKXZkyZcOqvt6G5m5JE1UI
X/pzhTaLL9+t1kpvFmby7iDCQSjKrZ3lDWb7f+a6w1zrlTAPOd/Ev1woYgPz
5ZU/BRCTKTvkMU23ga/dhc4Pfyz0bbGELkLaGtTFWPozHa0pkf0fwhH9/rme
1Tand1r7OnfHyTYne2b5MBqRSqdMHWldlTBcIkJPodKr5sHyaVLFeZAPHCEA
zm8PyWx7vIOzbsaPt+S1b3MTl4oQf+U/rgOioasbXcHjmRPjHIvJIjRC3lZg
ddXmSB+iDFap7bp8XVerS5zEgw9FgL91cxnck00ugD7bqUls74P/3BOUXpfW
g3VHf1FWOXz91mZTIXZvHQcP8uxn5oVhHSYbujBfXHlx6D3x9jYypn4qtsLM
H4OMzrh/Hpqx+IlmGNFkTakZ33SFpu8gn28HpQdE5pI/5fwyIH3y4F6a6gdO
KLHQc1QkFcHIHLIKxE6hGH5ImQGYcN1nPbyNxnIPjkX2gQ6yHokLsgSgX4Rx
sEZJtA1A4MuybSc5UOk/hGhlSyto4+oIBSNARem2STKsIRiy9OQ9J6+/e6AY
HXnwLdh2F4isWbxOnB8zVduLDQlD9beMIu9K9/sfRsZ0bg3MURXS8y7VeyNf
U6sRsKJahOSAyhwtWCATonTjR/dVqbjeGLAGbUjEi9gmT9iL6UF4kd6IOdFd
/6Rp4sXqCRQdh4kU6fI1HNpAr8BBC+HP+Llhn4Jeq84vxw1yFdObB6U40mFd
x82OlEm3NLLMqFRqNxZgw4ImH5KgDUHXVsfR323dchYpHkERx93OBIKB5Xi3
ogY52NbmNdhyXrImioV5QEwzk36vf5gTf2OlyAQnQaciny/zkVeWSde7hWmt
wmIyRK1iEUg4fEoUGNHanSlDwaFjFvFsh64ofX2pc6Oafya9x5tNI/bSCxgF
GsIib3C5luttc/Swehk0wQLVjZafpnqaKPOTsd1g3AVse9urYJxkIUiwt19U
70wsGnsnNUF8el/b9Ex3f3/0LPAUkf0rrbnz+jUGeOjuk0EhmybQZL2MjbEp
jx2W2koSL+utS7gC+wygBvMKIQFxmj/dnDYKNIBrfYN8/e2aqGBeyI+0nQeW
Zm3KXZeLW6liQjgT8Yrh3cgp5YGZSpjWwQ8z5b7TfPFGu6jrgPntEPfvnyai
iNYXJHUgQt1wEHs+1kDyjwP0gvW6KGL1vQt/4D3qKkuH3vDALJQv+pYnYc/T
kwWFOkgUkvUkeJ7/sdFXmKF5m5pZI8LXEExmlZSrJzYwuXKZfHfDm8ejsdRB
4UERaNsh2WMOtTItj2UodknnvBugpdcZagor9rkEouGuPF2quRinioAfTvI4
UQ4IhjCPkJ/aTOyomWFZ3DgGsCIpz16FigEBmt/JoMILjFQcHCWKGgfkIY1S
i7iWECFtS0YxbDumitbX+xs+ytWlwzT/4I2v0gM8muVX4VFdU5NXJBWmJViU
L2CaRRA/POKa7kx8Y/Ch6XnCM9rSPJPUdiZ8Vdf4W/A6Atb0qPRgcvrx8Upx
nX6ZrIJM32So3nNOnpwVGVJsxiNbhXGpBmIsAXTWQbUOTHDoaplHekQwKOlr
HHsggUX1v7D0umDWWhiOSVzsfnN8halVnHYYHjz5Vil9FEBqH7Sn4cW5dpG6
fC84fNZ64LFFMWTdt5IGQ/AYD+ElFkpPLLPO/xusG+Y8v5RWgwyJA5qouOui
BjFhfylBeWmAf7sn41XAg7jIXr9ciUoYVCFj1pcZUFSihhp7c5L8Lx89gOFv
zLt8XozEBc5/mQRYyNUiQyZkOgR5TdPHhI1+FY8OmFpMCRt+9bxnN3Qhg24c
unSP2wVFs76w9/u3hQpkj+NaxCqjZCr4R6lvNV4p8TGkKTTsZfVRXbWFUoiu
nVOceUbiWGE6AeeeQ/HSLxKjO+Neyy/RbLrfwt7W30m7nh4uvSOIsZ0h1noo
j1f5xyCpNf1jP5oHkAFG41Lkp9yPZyFEZzOOO3dnWwZiQbiNwxOioBdF4ukq
kCXQ4glKqvfQmuxNq+CbTmMQWn/kOCECNKRpEOZrMzze2Iy3lMKahUKZvEku
DHejc0Cv/OsdomsAzD/rxbLBgA9CTeLFYnwpNBadTNd+6mwFviJUGQJ5wSWv
M6xUE66pJjq5JVRBd/2634JtPbtFCF0G5HJSEZlyCwYXUec7IYPwrOX2zMsR
yPO05dfe9t+vWc8Ov5afENPZh9H2LaiCEMOHH50bcmIf1PHOTQoNI0NAcDSc
/Y8eBuYiyzIpumlMyswI10fEmrTlPEn/otb6EF8KlizA/e6vjgejhBJba0Os
KWSouviAmyHFda9wD7zRt75bwWqOqX+wbCIARtFoB/yazJloShCQebfG0LiY
E3BK5fHoMoCC+VDtCqrYnUJy354sVmVjgLLqLBzYUZSAc6Mobe9zI8kGals/
fcxxi8P2LcakEG5vQD8XFxrk4eyN/IYaeqC02/qYGqlRlkxyyXEyQ1Bzbivi
e2o0QLMGkKS5SqmGoT1EAbEN4KrLOzj3yohvozMemcDPId7PAAuE3PJ82+85
0GTVIfdA4SHYilyhunqT9Utqau0JdDsVOpj1cHACpdCVvktoCqJ0yX5OJqZn
24Kh/zkDsACVS8ZJbHR8hLyS/6O/TYQllbyI/FJjnJCKbBhap9WLS0jq5EsX
hEcrXf/j5V9a9QtnzQsbQG6hkIgdWLpaga5YGz8HuQRRFaqtj5prdgVAbfQE
HK2jhEWfIFbkoQ0pqXje+U2EuTEjb17oxyDa7Z52QKeYPtnjMJlNj1Qzmzb6
EdxD1Zk5BrP+LLtyC02iiJXjpOC80DnfLv4nLqwPMKn3dkCSLHu6q3+k0gbQ
r/ddpu+sLXdPYjXnznmwiwPq1nrU+wE0gAYeTO+oFrw0qgvGTy6wXEpsAnD1
23OxP+MHIrO7VA9DVSHcuTaPdqdGeRGW7gGkUNsiYue6oDp2MImezbG0dPa8
KPcqq6mB8mdxDgOvkzHtQ0QaPo5f5yoddoSslyinSi6eOyZUcg2jkBIo71hj
I3pVzIomtMTzp5gywwrMMwVikg7afLjuKnsYLnz0z+yQEvZSSGv05wARBxsP
sbs4wFDPWIWbarSU/hLstQqYsfjZX9ujbmHZqwK9lGscl/W0nuEV7nN7ST/X
VXYXUVvAbzECGtwpelaklJJwXQUD/bg4Gw52msaRRSU4VzqgSn5sIoWAwC2y
my+1FtADIeXBkfTzcQxLTeZB6Wkf5dOC5D4kDefhT12iEPgPoDV2JSdA0ldP
V00du2vCgRtHXinllNi0u/RZ/i6nSmYuOu9uLJqcNwTN0Fj21NA4wpHV7Whw
XKd/3T+uSsJ1dvJ5YkPEm4S9UhM0KNZNm5osrM10m208RL/8GLWH4F9rA3G/
+aPiIEvVTstibF8aTLx6Izg7N9VQBfZnO7+ZHy35zn6TTZSehJZtwUzN9No4
gORj9/Qc34GWwiR5hyyK0eTY9N5rYzwTc7VEutaH3YWeG6Exs0PvvD6azRDZ
oRyfyhaLWr6mrHdd1YNfcnSDCEvITfBQR28Qz6ZApVedhz+2Ue8PJrYY2WF3
ZvsF0W5+IrjZsS1a7eG0ffzUURTJ01VCeWt5mNsDNQjrHsu0eaZGdnYRu1cy
PNiF2QX6yi+7HjLRmfDedO5W84ysHNv2V5kYT1VUE3bEsH/4ew7FvpD1wGma
pA4s4BVrgwZ+JaN7tLjR0DKaRrtDTW7Ax2TZJdDU/kD3TCc/CKkt9OO4B0ld
u3b1vxjxGnO7VR1valjZTr56H8KkHDoAXjjVbXUgLpi+x9aU51XT25LRrNI4
Ot2BDRPalJLuQX4zeNtR3B4DLaKowJISzCcKhF2UvfGXFSrj0VYj+MbZIA6l
D+414Ka1yUYRDbDS0z+VaudQOlfPrQ7SqfsgEwiR7njWQNlA7OLA5IsxLdTj
ePcOcvqic0xiApvq5PBxWTHu5oSfVFqABUKaTydkSQaLGVg677EystwiB9ZC
1ZQoi6W0JGtBH9L32UOHGlxMBoJJUcqEXvs1TBcIgQuEBaGV226DUdxLptre
FoPcgdlwKWXQ23CMP2emll9TrJtjaraUlHO1DlOVrtkhpNqiJbK3mEAtsmQD
vbcBhVH85WMU8iJKBgP68OPcWAqR5Sm4qSkyJzqAsClbIfXTUIShVtRz3LL9
S/CHawQeP3uy7mHE4OYVt3u/dXqYJxUA5kvIpNFRav9yMU9seAOO43dtQiDG
X/F9lNpm1hTYfuXIiv1rReVdiAcisDArRjlN+TOuMPLCgIavz+avrnXkY6T7
sb2z7Djkwx1NGfookinv2kBTjhxOL520QGk8Uvq1YFHZAWjwtMt1LNkeuiU9
prfah9AOCYS6o+6hBFD1W6D14QQbLavXp3F1dtSJzdnJX5v/SeZ2m9AzKeZN
H5O767gRc7miC1offChMn14BmCbqUn5tXJ5yrNcAqq9RZGBY0zo6C4Auc/CC
ZelgaS+6YH8COjZH+zQVb+prYN0jd7e3sVq76IwBTSjAeRMLSqwund3nAGp/
1uze6oOZ274vWyg2E6HoN1zF911UzXcPixMobe7VVpxnedXv4fGppdhWAGMi
04xzV4icNWXol5PVdp6kaWCGOqlPKXVutpFRuonNxD9g5sq6y0nz7haS3cvq
B6yYA1CghV76YmsH2ASsD/OKcf/Mr0/sWi+jQODef79PUGZ5fHR0WqcnrUP7
lC553BvKRDST4OkcvOGvOG/tpfmIfrxEgf46AIH5syNlKcTAcUMFAvpGTv/C
BPvdcoEdAxRf5HFlAjznoytG/ZgW+fBOUKkK0B7HyUdbbSlLWMlwSVwUKIAt
3qEHobryZO5pRE756nv3yhPS/To8OEr7eVtHoiitrMGLRBU/XRLPttxB23BE
NZOuNSA20A4XMlAK30hWRwlMEIPR9pkw9BtsW7fCTS6VTURZYWYaKAzv+cDY
BgLZrmg+vsSww1WYx/4rj7Mk9r/NbgKVKWHNbD809jzC4cZMgWHuM/uTXfgZ
kh7P+E1SlRoDbRaMGeYaeqDXAXBhppcISnprC74TMIZcmNUlpQeJPxItaxbO
iF8Q8dW94LTVKKM/UveOzO4VssfnNcqgYXATWGeq0T8QduPu10oD15mcLg90
uRpYd27V/fZDsyGPSBxpHg8FIn2an9UOIv99HQgbf26OgG0cRPnIVz6lBP00
0gCVcd+goLkazWZRncsgNvAdE4HDpsZR7hf25MHYmD9PIkV1Ktt1JRlmhVuL
ULQq+svZCbgp6LLWPc6iJTGkKBB+ftb3YuOklgKjDvwxwXvsZ53kDCi1HD4o
v+EwqWDcakb24ghvw1UVQGgFJyCJ2I71KyyHJKdbIP0NGYWCU6VuCPFt/5RX
ZlI80xgTNrcH2HuAGmupELpH8876FmkVpYPiOWseN+FeIdNhf2FZ6xEjqhB6
Ms06kPEHwBxKOK8OiSxhwsIoYzIMlXbAFFmH4exXosG8EogF9yjzDY1VbBa9
2vi4D3MD9VAvJMAbt4OUsE2kqjh7W1kCNC+mvGrGrcJ09F5Jh1CrYWc4hjwq
PGWn16Pe+RazwenmmgfHA2C/qTo2azUbnX+ORFdyi2UPzx/7XJEN2F4Fane+
qq1BDTpHmz4xcHOruqKu6uKav7g7ymiAGWBfIWT0ZMZY09TukSsvRz2292B3
CToLwdXhjvW/piLR0FPBkyBecH1v7lcaBT/glaULjKcBBV6nJZBpuOcsr5mK
jvsNIU3LYJP1k5bDXVpazZr1BKfjHSTdRulT5UsyFtbY+CYWr+ilnFqR3FIW
hK6MAvJN06g49pwe0W0lsd+CmyT/9gtV3tkau2lOWoW5lhnXmngt8DPXIKkS
ljpM+wd/Px8QPAZt4KCpFK/y9QjawcQzHtMWMbWyiVJrYGEhzfI/Lsazmyov
RRYCkNXJW4Jie19pY9yeMwALZ8ok38AhaPfuLDrUZMMkxVGfNbWWSLvEczmB
sx2kPkxYTsfEcawoYBvrzgVDxxLnua5VdjSVAOFpPY1INe2A0kTk55ZAeNf7
u7HUVcrc8rTktbH2GNEubeEm0s3lz0nluSWcwIyfYBdKLo9Ch31PnYWgZhg1
ZZhQ6qV1LObwQS4Nh8sdhuHBAH3lYR9H2DTSbDu77Ys+eV5PpsIOwuAIUQAl
4pIPxcYx5FnfnrW/Xp50TUc/mtkpj37EdnwRVjmwnqzkuGgywa3qJiN+SH2y
lUtJnHuSDz6bUgTcQDPG/v0tiVDOSJeqWEqN4uUHJhvSnob0nVQOHF44og8L
h4wrU1yEtC3h8LtdYou1pqC5pBOUZbvOS/Gg6AjVFZkXUl2sLJJPlFjBxr4r
XGRURsXiOp43VVINoG3GrHzZ0ZjX7aiVxd4ARZCAQ7q4dQ+V7l8tvRI9xyKK
B8SO3kIRsS8upa7SlTON7aRUPYEeqxSMvjxnjrzH0OMtSzc5emu+xrEjL97A
z7NzfEk8gslvSPVGrmk+hPt5XSV7mKMEP3h+nNG7mtH6l4Rwc4xDj5CJNKON
0ay8ZJdkUo7fIcSoLWNmD7D1+6x/0FdcQeBNu0aYOAvCnNQQbaafRFmHuSY8
ayIf8Eho6UqdDzRKNdAYDNmbU6OiFts2SUAc9zdbqlpvyfikp2sPh5/K4cTL
7rQRdzoBDYdZVblJp6TkgVFq8Qg8W43XnhU5C345dd539wvYA1jN5DBJtoCt
PDZvkRgVGRD9zxTMwIwpCvIb+uyv/ieRyzn8w7+PHNrZLR4y3DmQm6mByOGl
cl9JKQrvgI5ehsEnWCkWnR6iRskSm+71UDeyXBtGXMB0KKCcRBf3YNFW4kFi
CKen6xIailReJhQsjv45CKKeFGIFIY5SCAzytK0SMuFTTohj4JCVx722qR0f
qljy+xyjtAaNO8ui416NLjVPF/Xuvsno9y8Q45JHpyArQjqFpuD/iMkCdYIb
hEci38dovjQP+NHm8SWv77hBVSg4IvNMl+7qv0tjRBi3e28mottbGRES1+Eo
RUA4wYcjpmHTAMnYISylNDA4jB0j9VCfr9INT30PqFzHSK35YtPIhnAiDxPc
qdIOorQWqpJtnt3UnW617G8FnrzWBG2kwO3Bt4cHHpuRwhTRv1XU2Fs4ZAeJ
TS+5Fv376wdnT3+yvu53xfgbkV+5jOdixabUiidX/bFFh8qsy+teIjlG4RGs
x99wBCn45Bp1azxSGjLilolMlt6xJL0gthUcVjhorGuw/btpwjVjjCr/jPLc
SDPrnEnyQ2Dbw57L8hIyWRCoK90wyyOI/KCqHeKLfFVDO+5ht5He+VxfBhwN
WZShqBbJw/Y6ouhH4X4cQ6O1oNfBhyeKDPhJZkd/LeIxjiwp8q4R6nyXxtYU
en7MAmsB/GqBYN9Rq2STT5JcO8teZX7KK4lpKSs0DsM5heL9O4604P1i96lt
8hZuwXu1yZR2smt76yBaP3liXfSA4y8PT5bcf35ZnFTYTDuAIaGyAUNYWw5E
w4BpUTDIaGhyOg2VAC8CNKOnNSyRaGL/giR2ox60O76L0xODOUWRiYi6IDE/
wb3dD6J7GCyeD2PPkRAJeZQophw+g21xDoiMAe6mjUUKe2Th0yJjMhP0rJvj
Maodbnii7XSUaNbkKIg1xkhpQL68SCraEM+3t9Pip3/KvMY+2thXQeLa8YjL
CBThLZS+oiLZ/zgM4i49uxTAfP+D6U0dQWXXXfbh39cBfMM9rxdVb6x5yZOT
6spRska5528beNUXmHHyTC8m2FsmZbc5aAKy15zYr0lRPa7vhN1EnFrWMbJy
f3aZPa8rkFBu3RyL+cgXKPQ9KXmoDDtZNGJmpKA911TXm7u9V39+N3JHMxgu
RgT0JawFPVKzjeq13XopqxAVxo2O/IF9wpdVGXdRmfMW7JqX9GziWm9C+bkB
BGc1PWJ3nbZGMNMklmATYsJx0uoteGJwbG5g9R/UccFSrfwFehjeHuu/+0sh
iY6ZCSG6P7MbzIgBstqcPQyERcjFLvhI6HzFYeU2MszvfaujRPGKaPhmlBEe
6znGoWhQS5SCQ9dGHXjKsLe3ltIZiW7zTdpfOinKNuQ3ZxFRU822RAikyx1H
Yl+pdSMAcLTC/d9yn8u4MiVNQXz1D8oQ5U6s63WlkKA9OJUcFoTdel8+hXa/
7ozL//Nbfuj7loSBYlnXz2TG3En6mB1k79+ht3bRgMEAQfICr1ADqvZBnoP0
j+dXmZsSt2MC1dPwOhj4+YXC7R12CRAH3tO+4tC6qtBxLoWVcKAXIf2cUV+s
CGu1ZlRu2uO7iySskWtDpo+fYhhY0mTA1aJuRJWjnRIoG0aLD3A9BpRCKrgZ
yKX0v6Nbg85xktsZJqcWv+NI4iOf7tKkSG7ghMtn6AoMDxB58w/iJNSq9OYb
S2wB8UpiaRbBBoeUiFuh6YGzvAkgx6AzB1ecmZaQQg9l/De6llAtaJVaqMBx
TjCdTUdJyFoeA+EzhWSq+Z3tvT9/Zq9ISpR9GXtvR/olEQVkZZ6lDHIIBhvR
HH6jI+gROqZPnoK3u1fHyLey1S9UxgcUdvhNdg1A7dPOtI+sE3Cpe9beJKm2
VjFqmtGvpyF42tdJ5BPpEGFLWCW8x8VCxTQL5+AlKwCFZLkWnxDV7keD4keE
tFU1y7rIZJGkBgueykRAeIXjPisK7uloVkZ9Du7AaA/qp6EbcGSTBW8hlQJY
HZH1VU4DRTA+bQZWefYXPHvXh9GB21DhoWJ3VtZQUoK9iLUs4WDg5SpnnyyL
+sC0VtiP11zZus6O1FAOYP3cGedXLuABh4Jc48HfOQYrvVtVvnk41FfaBF10
MnmbzUf1PueQJQqatDkZsj2aZr3UHs7Yu302Ma3hxdDgLzpq3sFkaAi5D2rN
V9iHzvPnzQOLglKiLCoi/tkxQ/VUD7Sqn91/2f4y+0Lf3OSCazhybzKZvjMH
se62VOylZAEeaZZoPkF7u3Z26x9mmCc0+a+mGkV/84JEqkL9Dv9yk9zHbnUe
o5+Sh5zPegNh3IMsz0w/Sifx1zKEImA3DwTQ+2x8cK8JpG+fJbxgB/bS4pMJ
f/nNihNlVG7fhoBGINbiTztUU+Y0eAE3CWBOLsesPmCge+jNYl0WGZp7A6UE
GyiGSqUfAkUiYpxPFcyWkrOLncWCNWdrQL9wHtT3MRFgIViCmv4rvTICvKip
ygDAYQpOp73TPKc8CXu/sZ2WFWmGZ1UGEqWw/na5zaO6H5MURN8ofL3t4i44
9PxVIj6HpbbfneZTZqn0J+nOFqy1emH6i+xhPt4hIXFDYbfKxxQkg9SqI9KA
L5ln/aNI4q7ApCN6A2AJIH4qUwZK8yCiKWzGQ50BusXC8TkiFeM+nKKBA8pM
VxhVVv4WX8jGzHD74G64tRm6axENcAcor18BtSiri9W+HGyCZaDPfKZaea4p
fk50NoAoqzocedIvW5iVRwsgQMLnK6JeoWYDFy0/UfEo30tUTR/jgcJOe41N
oDhAThSFu2T+RkYnOvDc65Eod4L6U31dN/Q3bcFCH4TlkN6Tf+4q8Syi1GHG
MII1UAK5X1nKMLdaaWxwjyuc5uinGNo6twvZaCqQBgqnfEVT5nlEH3TRSdL8
f3puEIWSPapCrhOZru/vnQXiBafWprCatTEXOVA4GZ0MiLDXGTaZGA4omn46
/1yk86ahJyA3Tv8CSV5IMPYMWc2uAlRGpeNeSGVshHMWmk21Fa8wFS2aFrVm
kdjTKqqfU4ZvxLCXgKEtzTdDyu5gcNxZ6bKqinoGKYFzI/wRHcB0wgIieKa5
nVP1VFjyfAQUoj6Fx6yWjTlcwknylNvj0jFSlxDuxCXV40zXFVsHwHKmeoXJ
Ho+iDzF+zZztx8hO6p556XJ3MAAp4jEE2mp6JsKMkrIKX+zHTaeHsXw23Aa7
HpWA3uhaRa6NRFGmc9K/97LkQ6SgIWNASagLU9xzkjlAI4pQWq6KOkbQJcba
12PkUF/k9E8PW7ET/I1O4mPx6IIOPjLWW/YSY2XKFcgTzsUAps01b+TOjTHB
YMOynTUB/Wwxd9Hlp09HIZE44NerCNG7BMBCzz2SFrpBF54bBGXSAQW67cFA
XZIIsPQhg4QNwejyr2acStQ+SmAl+Mo1DcOr9ORG6O1NqFjDZwd2fjjBH55Y
bDjxlEW08STunx2hMjz+M4YD1zj1edcuMLEDnk31f5CTPeNZfrBxu6gFNWnJ
jjHd2MDYVU2aBzUWF5GfV3oq4mTHYVpHgCMO8TQXN91ZJo1em8u/QjTMN55S
O2Lwq+53Iis9VauI6arrZe1vS0hgIoNeh/b11lTAlxQM6VggZKyy5fhz+eq2
ujHwnloe1xUXq/6cI9Oc2RGLc54B6O2SDo5azx1LEPPDM36L9URK+vAhIaAg
RgE6uo8MwTNFDYSz0a1ZnW0t6JoJKRz53ijDtIV8lBX9Z1FnlAkDu5DYHYEA
21y482R4hjMrKDgCDPiMl/pB/swUxDoD94ZDom90KqtSOY1Fv77YirfyX9cI
JpHzug1Rcq8RBPXVWrZtIl8a+7S/Qm3NaxvEeISDqqRnNO103eToI6uGLX6G
fJu0kVzMoqFMDWe682O81UfJqz9vzdG9PTr4otTeMt2DVVCWVHUxg21QFKvH
gX0x45qlInfZCL6pIxqKeF1IabGizjn3fMMe9CHORPL93eaYAlQdqp4tA6TG
poZdlBSuO0gAWnQQ0zmq7MxpgNFiMlI6FOoJ6RKDkBvoToQOuyWdYzqsVzkh
9unKtnquOo4FhOfaEPCAfoJS6Yi6D3DbG0dfmpuEDZZOR4KsT3GfZRwMQ7t+
mtbMfWSPsc5e4TMw+QpyvL6Yluf/eLWi1rPdc4Oqf5wC+v6rrPPASiYn9wwV
XTOEQbRO4VHeDztFcOLvAtyqf3VUOOEhM+uYjK8jew/PIGULIWLHWs+HyYKk
Pk0h0zeWyKzqp++b19Hn/IuACBs71fGvhvBoryUzcA21XavjYC3p8Go4jpiY
p9bRgsniq6CBUqU8DEf/6P5vbOOTwATZAGCcvRYgHRa4MZhHjsRhO0sHrvC2
NHFJOO3npiXdJ0Jq+6NKEF8W4ewsk8ltIT69JMDtjddQrg+eGsiFghL+9SLw
3eNBUc3P+1v0vPFiM+AxROQ+dHkeMdBIHLQoUNF86QxTB4qZOULjSoAXj5Cy
wrSXT9ANRE1t8XTuS8K4iBO/DyR6mzzK1d8TUwHIBZazCdjdwLfedeuhKg6I
0JXj/UN6oK7VWtDbPPg2r1VO9TFzy4sjNHFo4prRqWqxtTyFEmGLHzPk0iRc
7rZnz94zjsXxSmW4EGoUoyTx5ypnkKQYvryBbHuk3Ulhu5lODtYXC3Zkhov7
4ws3202KoLo1dWNKZDhN3ASxKmeKvAxSnYaQaEF4pwMVZ8bd2A0lGt+VsU+n
Pt3bHZCDsyjLEqZc8NiYvq0qp/qCAIIgSvdijh38bfftHSokzeBuZf+RkpJj
+y3n0CWb0luzoEZPc1BTyUhUR4P0th9OD84Nrs+hZ5KcozdQDCjO6Ue56Cs+
iquMJN9Lz6+G5GDN6aNSh72/oG6QyZj4ImyA+vEtPbF8cAWgDA78pI5q+mRs
COcSQRELCA/tu6oa23tkFhyvcMjQgaMn+klNrtmTgLpjBRftUYmGOIVWxIGX
R/yGJy/dGJaK2KUbreZUdiiVdwN8ncVXHnVGGrxi4FSKpvyt9uYLYt/+uAzN
Pbnx/QBtTvvDgNDVPH771vKoVfouQXeDEi7Q2gtdCKCSHJ6ggYRJrIHBRuz0
CIIskxkrrjDINETeWiuceAD59W30Z4suo55YDHBTOimPlFwI6uUSh77IpXTk
P7xaj76JIdTWOCXWwvzprTvz5PlbXXr/6CQ2aXIOIUqywUsv9ByO1dddp05Z
m1ddhwAkyxg3n2j/JP9afHutZ2nEHFKCmymH6Joa7P4JXapyYoJIc3UHbLxU
4bMGTURJ4XYG1AzoFe3ESLRzrpBGmyBOXPQVry+ziiLBsy+20WvVmwL93ZXM
tx8N6qL/tfcXP7UVGq811X2zsUurF38BVnMoOv5sE1b6HjgF4CgRL8sO/KCS
oY9cJeZ7jj7+BTWsmn0jBxkRsHg7rxUSP10idVnoka/iY2gyhztF7n0sHpa4
fBGnZHdNqcJkuNbkx1R0WrLCKII3r3o2NIFxZ2sqFmJOY6F1ARKwXxFMsjrZ
357pVLvH3OcnpRECGQlpT4jTkJvXCsDJiNRdNNDm7BW70YCSFdQ5Fnb4diOm
+lVkc4SCLC7V4J+5aTSDtura6vt4kKDK89KM8qlqZKX54YA0OrT1i75keuJ7
0T6GSeaBVWvBy8DpcpUzP19GtRncfE3/QIClZwJ01Z33s8PEaooRvWFikUTX
RKDPiA3Zt57U3GJbz9XM5Iex3JPcj1WaprB7lysdAP6cTLIQtixnZsxZQn9+
dTwO3YjYPQrD0U1YH2pdtIkNpBPD+FmkKROb0zpeLAFUAnjGp0wAVi1fW8xv
yPsxe08DnSNrwLa7Nl5pz1HS7Fzuz8zIHm5DRd9DWlINW5qGIJ58wIJVvQuv
UsGtZ5qZmSNtWVwnijzcKPsspfu8/z54RjwDxX5m3CGnvPT14r5zCmg1L7U8
GPCSiPmz+1kbwNFfUDbhiFuqZAC3FCFYvfRIk15ffF4s0+OxCkdlXpSiBdZp
LsMzklBAjLFzEC2VT+RmTJsyju4/YB1JbNYbYQkgBZ214eF0cKCiqcfy0EjQ
qNv37jWWh0/ZCeN5CIV/GJJOxxU3wRBy9dnqPLv6L2YDCWAYx0cYR4tIlBft
CGjkOur71S2ft0mJn4Orojz/57kAyns8lxB+Byc8ZBpocaO5pa28/82LTudg
Vk+A1fF5hYZMsOVFgxJvAHK9pKVgJSY8vB6fDUPsydHgmW+HwdO5cm+WdOtG
0L3ihKI9vkwt5jNr1E9XdhC73KuGH5TKTQDJbLchWoPXQ3NelqdGe6eCwXzk
pKkHWCCBwzJZsybWZNpDEDwmB+lJLWwaewJw8wM4/FKDfSox4E/mHjYiVHSo
LzntZhgjSD4353xeatZhAiG31lIl7vYPXgX0Z3v3tYXhT0EDvaJdNgNEVxCi
mz9/QeaJMpKXTJlRAXnRnX4iJy6Gt+IfOGXmbhrCoJIRZLSr6kfr0JPS2Tl6
Lr5JLR/OhpS3mG01a8TPQp+ZRpaFa0z7imKgG9FAnI7P8hD1yoJU54p8UuLv
fPmpckeKJ4Y1mcePUOD3rCQ6NFrZK/oSSqEgBp8sen1UKaVGexVCq3/Ny7YM
OEzaRT0IJ0y4oBu4lcAhxMTIaSMKh25ntUC5CDgaty2Zf2q5YKphvjYth2M+
ayAW7y3vuSjzQq7Nw2PGVLLAKFTq0/DzRmyEqu49VQsOeL+nZmmB4r9KWCVl
I0bbrMM6kY8NTn1k2miQK1cRF2AdNBSCm7V0W6hRTeWUVFRnxYrEYqFAysSt
5JThtwO7NrKCqUGmrOGlGD9KVOZjfoUIJkNFVTEF158Wu8QsuYEja4f1QBWm
+6h+72o/3Rcc7uuBSWFg0li3gLgPtLVKGjU5GxBJPkAwnmsCaPgWIZ6SOB08
dwZNpV5UhJ/1NnZOF5gNi0DXTxTL6Z1IVJqLxc2OzXRg/TP4WGRutptZp6u7
WkUpRWv27V220HsYMi5+YGGDi+yK9WkMPuPUcJiYqsrMJZ56agU4UydP1fAR
cNJ8dvpPt47YCMr38Vfa5PSpeppv5MCayYwo0LIF7CwDMj0MHAtqDTkfScLO
bMq1Ng4egMSmF6edzZYV9arIKAIMEyWkBCAIG8ZSbOYtN/vG8p0beJBRPtz/
P7lDQenNTT95JMMV/GjLX4FiNsoHepB0xsMqwKrIm50pQG+JLcUrdFiokvxT
w5lKrMr+3VV8md0aYypVmL13JtCEP+nRe1ZyxMbL4kyQvU8xnvRTQrmLmBUG
iFzlM3MmMa09mtq96QoDovIMhfvxTunL/SrtTk84VTd7d15cAdLDHYOlxcoQ
+MAOT1LZizwYR2oD//KLUk9Yk42Def9TDYoz51qkucc+/LXzYzcGwQmnFNaG
NRjfMqZUcKI7nUhBneaxYKNcto9xPJRQxY2gCT4L7pLZXmNok5K7+QsRxGQb
WPlr5klcQ2N9BuW/XieOBxrBGrcYL/mQsNk8WJrZIPveJS+7iTeSW1ybUNNw
K6whcV85AgTriw6nfCDmBz8QR89le1LT6d6x1NA1nuwBqTeauPtmxDMqE1L2
OWSOqXwVwbrM/YgLQFulIjtVEPMvU42mDMiT2Uj0adQoGRVu/oYg/UsBJSRt
wpbSHpAPWaJkarLFdy99x5oKIR+GERZGgCjn5fIiNwsR6Qk9bE/LMagMRMVw
gUlf+Q4FaxSomurb55D2Fj+Fr9H41akSzklLO6oUNv4HqPCIIvA7tbJ21coQ
wA/zHCjH0Rp2nbAMyhO4/dOGvyiazTzVwS/KFk0DjW9KbXzbUHXpXso6Ajsv
s72ylhe/itP9D8WcGbgc6rviugbpje916Ygo5jUHbTlr1hC/j8HdykBAWbUW
f8iVnYV3z03nk9vjCoOYHYsSUPD5PyAZhg8r4PmXGW3HT27cDjEAi+FQaQD/
EtHznQGzUXvFjq6f8oR237huv/kjP1TJsu3N70xMh0wxJrHaril/RniOzFZp
ymHcB411q4PedVKXDoMMZ60Sm0dd62mN1d1Eg0Ipuqgenn0gfI59dC9S5XK7
Sr3afrlQH43imSWz1Xdtz4ACoDBVMjYDQ2NZxTFp9V0duGW91Wl1GOQRFO86
cLfRN9ppSV1LBJhg8pxZHAO/u9vDoJ8DQLp5MmpaCggUXCjNe3lWnSZJcdfb
J1On7ZkjzOSzmL/MHl4gNEIlCuMfSuripHJAHVj18IXp5AfWqpHWGuv4PgUV
MRzF75RVwXwv/K2vSuT1Nkgi7UUf4Pswo1M669mqF8l/K1DjI/mJDOQUueFb
zx+kfCYydsaUrULqco05Nwu02zkF1Sy3MTMl/mGk6LS0wHH+Dn+ozY0ixe+N
lJALJQCZComZA2TGeayf/iTvtev21m/haYhLvmx7T5whBBwk3PTLNxQN1Tuv
VvqOPzrYaNNJlSPggXMXgNcx2uIsT/ZTsN8dl98SwSaptb8FDWjHb2/vkcha
4KzVVnPZwzmm8KMxiXD5M9XAJ73hT3MQQnIdIxhIWpHHFddGzjIDT2F3AGky
c8/RB9n52m1kGYB/w072489P+/0+dh8I2W2Jysi2hXTPA2D4ECBe7A9wlBTK
g4rGpwBIQ376e0q6E5Acrch+lkcrmWtRWPigPel8XNPARyWglXpig2RmWHcr
kEJqwNdzSVeAx3MJ1Hyqup3zbdrTRjC2EAgaehSnTp5IyEvCn/4yK3C7f6/D
l/vIAUo+AbKrTdI6srIXrZy3w3X2Bc3ryXSv19v5t11ZAz0l7gjj/AV4q96X
juyVFvyti4lD+oKZ2qga+3EoH6BDmZ0FGN310B163kKisXxGw9hVlpvxsXim
oEYNrbzcETWvORViGAMEkq9AY17WhgMDNknT27OG0yXaTmQqqkal5l1RFxMq
SeBMzo/CX0pEE7z9rrhRbmi1uKinuYJcGQ90Tnp1XvoIl++exa7p0joOoYIo
Lk2i7s9So5N+x+DFoGGwuUC7bqw4aSbYFRrH2TRwby5nTNuoisFjeRVgcBlR
xq2WGSGESCG2YBo/RjJvqwjQLdh0/CUxDmT7PiNilF/ForQm7d9rqZeLqsvF
leNRu5dq3exs34qzgPFr6drX8Ktks1KMeJi0KQ0DGq2OiJMfWPyU/ixV6gVk
0B0CgdUwVooW+lMEm3+j6+SeiLXA0CHw70fXoeUQNXUqRxNdHA+CSkVOJO0M
KpMFJiyqzh4OnB8+ma7Km5zNmeBAXHq6JPtnRXFi5d3PYPJECGqi8bpcNJiv
kEa93XVyyObj3R6URekAOa/io8Sj2hj5IaA/WjPX1uXHqc/46LJ/G0phofRk
EeJdEl80DQ7GW+/Hsb4o9Lq3WmSf8T0C0ryUH7RyBUvBhNwrrRZnfrk27D1G
MG16Xpp0tUKbwDNL/SRO+kodwuV54RtwGdnlpq1oYy8L5oHanovFcrKTROSe
bDbgRwONfzDKMPsV/Udm3habXrDeJecdbMvCIXSfveZOiLf0JfN+jGLvKJmC
1bLd33//W081YL4hqw7DRVKjIqztzyRS1hWIZGsQmPPVdKCV7iIj2KBxMvZh
CY7bKRZFEVSR0C5YpnGI4fqsDp3nzWB6WielkhUsh2UiWlPs3byQAQ9+Beyf
bauP5E9kehrHDahYYUg9vkT1Rz8uygkYYfq+Q2erNkSbS5ScCPiHHbwvbgpz
PqpFM5+NYEDM81T0S8uFnA38POQKioOOdRB8bYFRdUdFay89wOxfXzG5fMnU
uSoivLKL7/nUNm8mDAhUlq5HoM13Whn/wVMqf2G9d6ZgbFgZXVniJFx46TV7
lmH/wt8iEVyhlEX6vBc24XhmTUO8j0fowc4L8zKS5ddV6HejfpBCpL2CAIa3
XrYPISHGFkzHNdrADhe4dtkfZlLS7u1saZdgpdu1a+GOTHY6d/3g2CUYUw1C
telcWAzBZhgkxXtzF1XelJ4RCgxMfwEHLdcdq63j3cLQh1gCCFtvfzo0bFf/
nAjOoPUVc1rE4MGcmMpd3tIumTMjtBn/xLdtO5TRsGYbhXYlLorr2bHupEjL
nwCftryO7SBdpYl5Zf3aDdiR4XN1ktK1RJWAkDCLP194idy1sIiF7IRsiWLk
oRVjewEVDoJ5R9LNIwdNpmlxKxac6dxWU4Szn9LbVeFW6LgrLPCSYQzyhIlu
9lHZIR0drfbuQYsntZTUd50gTBervoYfkhCXOaQQsdhMfQ9+a/KzUUo9Ks7Y
YxCuSais0VkRVG8y74UrFZpALCPaHBPuuCOr3WS5E56QvA8BgXhINta1/Yt4
nAG6oU6fEkA2CmfKes3yWhDf6i952BxhIvdsYZh13GLx/TkSIa8oqGKMV6pB
VSUHjxgX6uhgo9DVv7tbn1gVg4bArnb/nDuLMHJSAKiA9XO+P78BYSjNcXrP
+WvhCGPdAw5kOYm1pwLhJNy8ZWDYC9oUMw4QJhv2n6Wqu/6wVeMwC+55DLFX
DbSKEtvNVunv3dW/8j/00xsgSZpgxIsbGdJRIZux8OGZK3fp07++TXGCDzHS
czuhunmxLtUFXv1knYm/mDpf7Q7mcpyiG07UtaEZVNyBeCtXpdxQXdn7Uun1
KQSuHCoKx8fG79rk9jb1yJh3Oc5574MhTOaogw7jQQS22tyX/K1x4i0YV8OH
zUm2WtQqudtwovEENuAC8PAQwETbW3s/Fpryj+wjIieeUJJdKKNmy7WuQ/JP
0jPadPV1/o8VgmHvAUD9OeCSVWaBmZI8LD1L1dvr2rN0zsgK4+43qLa5eqwL
sOGD2sOBFzj4FHNy1sxo2pswxVeO8/hdxYCCj1/ZGmEumW7AaeI0m0PRsNci
jjWmNc4vMupHwfAOp0v+fDnSL1i1lYr0gfuhQh+Z0gVxF57SaQydnTE2T6pK
I+Bb3vE8evHITlIXRIypUm4o+fSIoiFaWIhs5JJqnURwDUMX7kQMfI1eZV8Q
18JAdOtDQLaFnP/qqMtKrKXBU97mZN15lzcdCLMrL4STTqRJZUf6buw+KZkw
q024ld0JrCEFyhz4mJg6IUSyqYYGq9N7hrDI2o6QNgSXq0U0RhC7z8IVdXhy
luxRcSjG4M3mRqwqS5YaHP1BlaR+p/xhwlp+Pi8gWkGFcDNERFV+8tKs2EFD
TJm7TPBMrp75VDqLGuClmdaNDMA5LRX4JFNdojpzpmX7T3s6+Ypu2EuBV+eG
G7qweWU8827Q7qDLAlisUY0stgF7w0N215S1AGWtL4Q2Mt7eJtj3ejCSM9ql
gl03M2qf/tKak0OmaOm9Xl9jZ2QtvwRHmgveHZayw5ldTRHa3lkvL/G+QSZZ
D7ATSd6kflMIeHBEewxRxdsL6503pFZmd1vYCJ0PrqKg1zr6DUxVRLrJDKZB
+Gxy45nq7nrxZfalaBElwrQ+pGJ5hVi6/gl8RqAGpYKHiKH8EiBB+BAhLYum
AhXAO1H7KmNTq2p31BgTgxR5v3ubwwvh6fzVDJp/HFXChNU6bIzUHMesK15n
TWTLxzNpwgqIMfmP5Vv7GS/rY+nav+lSHlC4mxgtcM7HGJgENB7V+hf2kNN9
nJqF2tY9vtPf2tdb9SJNuNte8CzN5dtU1BqZBSwQzOWURSSNg+497/BmQvVk
n8rW2Evqvc8G9GYGP4QmixyWFmmloptbarbqx7EluMEwJ2lX/jFpsPkP6oBv
+BEFrb/Cs4Cz/AQAHodPjglt5A/QU9nwNIEvDFXW8SjhTO/iEr6pLJthUjAf
v3p9C9Ex6iVavckWhNDETRnbFcglQy9g/aMrI1wAFovS8KxHjfiPtQv294ZN
jGPrky5exV3+MrD29HMpVzY721LfHSGk6MrMjpt8FTgsPle8dfO4mxZui/7q
hYWTxGsgpWZKvs7uad78LyZVydjMY6XpOkNp2ReB/ZgUVuphg/uAmpn6Xa7x
yXynJy2kXQ5gqA+erZ2+N1Aik1hvU2AJNXABZA1oD5EE9IiW/9su4pmVdOq2
ycDspJ+fGSbK0YPQJCCT4B10GlnhPrEzFlwTV3ZBO1qAcToRTyB3Rro0gwRy
mxvfg88KxCa1/3EmdMLY+SizWf+IyqsoUdY+jxoH8kJVTv1b5zp2/IL/onVl
s7E+av1S6S8oLUw3eonG3jCFPa8K7GLVrZymupaME8lgUp2RryJncWhlAF9O
33TLnHL+bKZOBlyu+N/LFiDWmHVoiEs88HaTnG3IiW9GGkaqmBWgdelKkkyh
m47mpSTPsnkA3OmG8iEiDp7WwLeq4VJRKW6kn+Rx+tldCEjZcitldR+XRdqU
9wbgbHjnUEHU6URBACtKWFlAwBoxTzxY722wnXgHUmGqF82M4o3Ha/BNRhLP
g07X1/bX06t3nx6tfBrC3RG2PI36d/03qI7dpvIIPmlcAvT2Mx7ea8Z5ppdH
9C98WaT5pPogxHk0O7abUZIpLO2kVw4EVd5/Vu3NNZipj2j7HF1iDRZDyyEA
IpjGf8f9ZC7jYS9MxUz6uHTo2qxyMe3q3yquvPapRfkXMtoaujsIZitVuscQ
8KZZU2fTrq8kYOmhC4aUNKVA7aZK7ewOhKFtO3xtwFYlEJKP8hEamLJTv9Vp
XYhem8doEPPA6EC+y8qvDNCToVD/ntA5l3Wdha2PTcH7mPCarYBOJGzTnlut
SO2LAksM0x/LWsfy3+lSiWk7GtqViJjkm4y1BMTwVUY5u7G4h6tVWcuiVdtm
bQNJQuzbQjx2yGvHevtC1l1QaAtXeIkIudTXpa8jb2yhha5Z0oTnz6kFco6Y
dNQiIV+OoBoLyvwAqYh7vv9bpDTggG1a1kfitZATQzhWKIXSCEge7PDUXf4o
f4VuA7OKMKBpru3wA7XUe1YPEUIw1nHb1JGVhJgg3Rc5v6LEcuJwsNKewcPJ
bifgkJQzAOJICq7zv/PnhejwSXUzonIe7pBZyunv9bp6voaha7E1FwWtCyq+
pDSiNmF8JurqtBqcKSGlCxVwoMHShno4+BiKD/6mcF6OZXIJntVrfm4uu+j7
kgIdFYQJBoWOZL0SsqBmhpxLizAINUqZDbOBlc42M85JsT0sAxOEchCej1qa
0tmh1E/Noi9edpV0/7YrG7TgRX5GbcldWbMNg1ILxD12uZWtWv0SzMuzjclH
wUQg2WZ3P5qC09j2ax0J6VRxTTgCL3zw4ZwKYJyT7o6ze41Cm1eIcKX5YumK
EpAMiBuLde2XMg9KFVXYz9ajBlc7shP733EWN1sDpPVdQqLcaM5tiBcvgtDW
rxn89ViSxPB3R9rhootDYjnh1OvKUtkqF6R16Mi1rrp+NpjGc90SPKEx5M6y
jfCIHXWvVbIuarJ8agjTLqPoD6IXzEJWM+z+Ke7eeDJAoYsjJFBFPPK/KiXt
sDIO0aBjC75kDJI7JCpGzxNYghE10OQn0C8f1ZMvzdx0WeaJeZW2ilE0kfJm
JmNRlrp9xOXgtoUVb/z7unuVosHbq03kaGl63HeSNItYmPEjDA0S3ZL9DiTI
bE29k+iwow5wP0osUkEN08VOhinSJbssHH2hy/ShGttNtHYWRXxDKGLe/UKc
wqyhHk+cbwoYYiMpbZYz9pFQa+2z1UoE+1KA6950Ip412rcfJE1Ls1ZUvdaN
S3UKO9wJa5JkyaS+kfJPN73dvM7qjv5Im64bcDKo6NLA1b+6gcYg2qGV9cs8
DljXwMKYAv5VCwaaOvI/ocnyuRYAJrynjTXnJt05DPzcEm6gsq30/nt6LD+P
vfICzLbXWqOuYIzxIFRqqTZpB2un3vcejy+kguhwkZu8OOmYDj8v8Tb2wY+4
b8rOW97N68SjFtdSFCBiiWmN5ck6N5BVdoxoUqsLqhWB9pXvRIPbtOLpXoa7
O0qkQ+qM2jjCoGTW/e2jZM1o7zq5XqUafM13TdIMhSz/tNGCHnAmqtElFWjn
/ZT3v/c2WwMhIWJ/b64+6iP69QF3TZTC2lt1cGVjiBp73zDCO1ZeBiDJk069
6M9Ks2GBIhaTp/sfxg0FCjM1AlEjkd8m0Zg5/rbKm+7Yc4WUf5gcAFChi+VU
nBgaNY5cAjQmD9HOe23UFkBmw3fbC4N/geunoL8O7JUDylxXnAZXKN6Slg3Y
4jeKZKmFfYCqtRd6xWHktEZoHaRVSCbOghadQlrAan0sJSH307QPxvmxjD3U
p/1XHbHQG3AjNKi+W58O3U80BX4h7O8RUBXkAyUW5Z62CfCHH/8vclQ/fzUT
jcVUb1JAh6/ZN17Tl3lmEb/UK+U0ARiTwzr27oBxHPmjMbtpmEKzFUe++inA
Y02Wb8zRoGig2fs3U1XMCMfpCavMMe/sdPSuaKqoUOFKIGTTKJq9n4MaAJ9g
H651Bp8voejm+XccSlDCLjUqsZBlZoJkXlSo9163BPxGWvWlx46w/gsMTrmA
0F6EgUgyybzT+JDv6azwy+renkD6wrcVOt8KXqzrtOsLE6IXrLIbJQgOCOW0
lAV0XBmVyRrtGAgNj1+TQhIWhVIido2VPz8Wevuc/OU9B02sYT1V/KcFJo7W
RdKc78h08HICNWpjDHxrSNaZaMK9Zvo6Ug5/stJ9zblLPVpYPjLWDY0EDFER
Gw0SoY+xq+7ACXhBnZqJ4AsgK0z559NJdwemlWN09VLMefL/9o94ra8VDoMX
1Co71p+OBQOlIv2k58b9e6r3ytxe+h8tnFipc9AUMeyqe4YoYY7VWKT+obVT
PTz+lkIda4vTx0YdYXWxCxKtxbEwKKo7wNWq7HjZ83/3rs4AUvXsLtaa02Dh
TCSO4VKzpFvz0q9YDncKHV8sKbPkXDMx7R2G1QnGQtgxKMcQE2mwiIUz1iLO
onkI40S3SJAggypHVfqSvQwby6l+FVJQ0Y9WSzpAnOjsLVJn144nkOSu5Uyf
Aybf5wGsohjSshUoLv8GM86+EpHuYJJ7YzcabIuAHoPkA69ZiLZiJvlSKGKm
MHy03t1XFNXisV7kV3xM9YOgWafNMEWJfYNNa5NR0RkayrkMbN7BLae+1vY8
TGxI1p54RhPuOaXg1V8SwlbjBB3JzGoGpbNLu279DhQ7Rh+OgujO9Epwtlw9
WThJ9RTgIB6P4KCG7PpZjN/fbwRx5muFVSQmRX5uz9v2j3AJA9Zspj1ifxOr
dhiwe2QdTxWsgBtP0BrDLCjh42Q52RYkavgtAnuKTKVng9iS0aM6fqedrZwB
uc2VZsSBNU/thOn5y3vIbY8b6IPEjA2azi/LqyZNM6REC+zpMsmV3advCPgJ
beP2K0QmdyE7yoqHJt5xkllzZRZvu5z67vGRSbUAiltOyksH5IuIe5E3jzDt
w0SIdsjn7x9LDOL7YbyLMLBaeAiubz9933+8uyPEP6FGfMKafcV6dKIwV2JX
impli3r7hYZr8Evhbs9Sw9bY9VjW6PyUEieMkDwW0cQNepR4DVRDWcG3rb+J
JGT5Qb9OUskpDwhBvK9Tqb2bf7taE8AI5+WLVbKfDGOEmNiZdOJzYe/g0C1C
GwDy2Ftkj3NZ4kixJYjXns5Vt+WvQYyRpZE1gT+92qUpKBp51eVi6n0t+qjF
sCFCGcPOsP19ukBwUQHPzvmdrFWQXeblT90Z3EGPlXr6Uu4eIV4CR/CgcnTJ
YM0LAar6zh+3P7Htip2+RZyMzf8kn10yn/A9mPDx4wkVTD7R/Gql2RBwG0Et
Oa31axh3lugCpFOAHRYYdJzFXjgjSVslGdYED+FNq6bU3D5n+EYgl0PD4hSe
7gxzGTVLcvrKQpKp4bT5aNCzceD0yGs4htzMVpyQXybqavC0jBFKCnvRV/vH
Y0CbPDRsomyhs5AAu6Z30orjeahUOqO8uITITwW0IIXp/T0kdDOvRiG6juO5
riYsnyE1MnaU+7n8jgXrdR2qlJ0cvuzGvpVR9rGlnvILDalsq+qxNewC5S3X
nsGEl4Ua1ExBfuWoADxvn2xSw4/9Dsmh6yn3uUt9b0vnwhuU7bX0RAGNvkc+
52l6AUH6tRB3KjRQLxEi2JHagMjRHlk4q9LX14nA7PdRESsS6EcpkNTwPX8m
sH1gJdvWBaSX3bQIaKI9rbCpULH6au1FEpU2EibQV+hGycvEe39jP90VhZxy
1h9CnZBThufl/Ds1hSuzLL0NVPvhy9naO+efuRZnPWEHjbNdaeR/reDhwUb9
qcxMrRlByY4ZVY2XuFL97XVmmwYCe6neT+BuXwazgCDCnhNif0nr5x1ML88a
qjpIlnlr6GX6SXJNGp7hiTL5Y3hpgXKsnwfzoxhkF68g7bdtJg/fpmrlJWfN
OwHJE0BIXt9mXRwIFvij/zxaOa6BQ8H1dHe/Necw1xc7s7ZXjuPoZhOlDw/2
fKfZR2bWDQc97SK4vw8pzv5cC9rybiWCld4UXTIonFIZEV/oi4/5UkhuOKr6
hLC3qt3pW1m8Q2PtI554WzcF0BS9KJeZ16/fqabgEx+ldLM+WWq3L0/0xjMQ
/NTjbnHk9cvZnjOy6qiV+4R8K/t4Y9/q0ulD18B0eMTtS6i+wdmvkLUCDDuW
gPzQ8e1h7Yk3wUhUgM8CkeAgB1o4MxSWPhpSF9o2Ry0Vcf5VOwtrFHnjBdwj
3srXS2/vHFvKULKrszrH8X/wuXfGjTZk3hLFFPECTkEBI2nLggAvqLljLUEl
pHdXUHFcsQ/Fsk2RvC1Fv4ke4jHeiD3yHmIMoLCzgvgqdMnOsAle5z16YPcs
TuGN9wKpPYRNP/pIPU310MaMOKvhEd6ymUKdp/HrUBeEatZyszu2W6cVXqGA
4irMgLZjAPk8US0f27sN9qQ3/xZiivXgA+AImb0fcVcJ1v78l+xzR1MNOj7g
tZpRG2Y6UM85utXmvwNYy6N/NctD8LQVg6tdF+L/pQO6wUXXxAXJJ6e/uJwU
cPAPST+h4UBlSA4Lh9ATzpEErWVgA3cd/ocbihgncuTjG0NkgOFb1N/yLMqk
nEDPpJei5L2mli2XfFXWGKMG96kdF+ntw62xLTGsBnKW0x++dNlNNgL6bl5e
RvCzGRp8SOe87NFpPG6L2fVdqvBJTvliZqfGPBvpJ8FWMDbA0ebz0ZPVJD+M
oVkz/E73A1J+EAuMJ2oAisuQzIVuDHLS6T3ucdq1ptGXjlQXDpfSq+IwQgPI
lK0ddG6PrZYebtaDJcq2jBf4FB94cmnUTb/7cAfVLIF5Mw7lvzb5TkRm3AJj
ItcbWUxQXgOfGnDLcY/pPQuOVZg2EF8KZ7nOXTJc7fDS4AtfAc2lRJoj7AQK
WXatnt/LaJXoraL0PKcR0b7tOKM1/NzVprwBThwU22BQREaLrSBAb4AeYWbB
8c80zQ77qE/6+oBlKnTzTgJQsHnoKyW+rl7PwhW5z+4fFwwktuXN8VuKOljW
ix8Ee9S64f4eQTjUi0vhuyVXBaMs7BGQzzhN7qbfCv3lDolUf8rI0oehWZzX
2NRBgibamzBkphHf3ZTVOEQagqvID3MWs0mTaYZTRntwlSTg3MLI1tOdtmWH
4WjWCDv29tgnXPP96DLeV4601kbjm/wsyfKb1z8AmVnV5fNFabL/j+5VewEo
LUJrs9eNdEEO+t+CN4vCO1h9PfvUcZBAbmp6UZ5mUJXCXgRjJ/XYeXggruiL
L3dxLBR1yUX8n8Fa6Exerivkira3vYtGoBTAArEvfQy3QD4P8MMSNemppaYz
Pofcd1dyrj75v65W9zUCgulkxcapDmYXNn4MMRW1qOP+oWN/juaUWoz63DjE
7S3GgK6ALGfajJGF/4G9TMxK9wEAqGBhr8le/fsmMWrEipp5/r2/GbZbpeFd
vCnDAlRamV9GvqMF0cWZyy3aBszcJVzj0/k4PohMjRShkF7RmfeVjpiXqW/c
zFSKpKpbN5Jeve3NoQNw8I/I7VoRwc8gKUhB8eEKIf1Q9YjrsQmVJyxfBbWu
wHVG6ZYkRY/efQw0Mt/AXPgWbkB3m6Px9ODgLhCD93TcUmc5+m07JkTP0CPJ
ZDLbSIJ+q28deWiaYFcYElsaiZ0qTaOH9iTsT99SQw0m7P0eDSwPwjJOmAql
PGxkPwK19xnCb4Rexc/TFFZKiN4W4LvVbO1shWTfbnxJPgA+MojfJnemuqqW
KsZpoN8rGEL7Won/SmUgyQB3vH2EnFxBdgY919+XGJ7Q9wy91y3GHDBHBaZU
oUDQRjdxrhEd0XePb3CgMzYMvVAJm+V/8Gle9YrPCQ0TAogwLODdrtaDkGUU
aNiphJRBSkxO7n7GIqSB7MtuFBFHtXuS15M/q5lEvwUr58AJNATN97tsIEXI
xvCriQO0qzGAARvYR/4sDfxcGwyia1cbLE4hprWLyBGGJuWV58Bp64l3plLh
gHObPTbISk44N3DpwIzplodRqCj4tyiO4+cHHFi48lJIv/JaKEtI4CV0+V8X
k7+J6AWG3N31P0S9o9gSv4gbh1bmOuIBbNLjyEKgOZt3gvO8Pg3JXjhmHo8b
q8ZIR4w3e53ssk45jIea0i3P4DoELZYp7Ipnjf3Zl2uMYsBvcqVJqltwf6yA
ujvSUGsq1aETHrPX/8NOD/TppZILNmPolsUb4FCU0qLA0XHTUhOCtGscrnV/
fpZr/j00pTJASj9tBX0PhebmW1JkZSFAoR7vsADPEeZkvAcAHidSARYnIeaK
okAizcH9TlZtE9EwnsNcX+ssLaJs8VZH0s2uKzkOKH+p841PtHL3rOYxcaRa
KsrX+jHhPyejvg3J0qxqbyThuOpdw4hpTy2a8IivQEhc0sQaxJbWLY851OYD
pmV3u30kmR/GIVjKSXt7ZojllOc9axbosGFavM++/Th0y6z9+LcdvCok1qEk
45nRl4VFMMMtiFh/nfPd9EiKUz3w9BWZGQrrji8K9sTyp3icuPuxgpPIjO22
RLmyDw2X4Puu2J4uMAHlQtlHYRYyQrk2qcdlnUE0cHSK7Nx+t8IG8rDN4vpo
HvVPHiXYg5H+LViAqgRMu8le/YflmYhAaLCMihmkOsCxi9TK4q/z3iS4Gc7G
HLf4jIYZYMIILWaQ89e4tHT1t4e2TdEO/aywnbEubfcLgtG5okBPqe9mWJmw
sAbc4mNw/pLOCrHgtnZeWqNDgZc3bplxydBpNHFORzzBmTY2vFMz7/aiLBhL
sYXh540LlT4dgpJqMvyRlujfTO+EOaoDBBm0iXXtFYvfveq6eNwXqJjTU4vm
AzCXG9WdH9TUmc8W11oGYf+ix7dItT6BYxuWZJSYa/+OC0XQB4OOvq9BHCiS
AoyoD9iVwtmf/xQ3dPXtMDGWK1D2vbZySGknZISR8hmvWiSLbzmb7y6uPM/l
9Big/ASqv7dHG6UxMzMFY4spvqCPFKuQM+58qtOmBcVuQfSyerDl8Ouw4OnD
Qo8bHt3OGo/W0ZMR99ecoA1eY2QaeXVkA3iq0yrkDVQeLgsij8ufa+1TX7to
RBUG1UtchuZwyKsfGSadD5iF74QTxMoMmNpaxOiSXxYTAY9o0Bn77rLlr66k
AG82SBcj+1Qe6Xqt5nC8mIUbZOu0F7fr9eop3zv1Jyj5hwYbloqNxg6LDccf
MyR3DqgviBAHfd8qRJtqPx4cVVLE92+WxxwTSniqc0XIUpart5vAmc0WfwN3
wkMNkz2g/LXpbp+55iuCIJiuH/jfeUDua6TyABThiK2aIIzerxv3dDMbfVwZ
mVyLI984cZKzGeCh8M1Nj+NoH2vnBBpxRYXEbluiXC4E1iAw2qmw5mjpV+fk
wBtKPlo8pA5YBiuj8IjVWnAaNRg0ivAbE9EY4TSZFnFsQvKF5PG8g54g9WVn
SOiuiwFimhkZA7v3dGJQnIRWP9igy5cf03/hq24thVlmvT48m24PcZ54LdUc
K4WkwqiDdWtB1UQNKovnRi73muPQLIR8RG8niPSLb92A3uGVNI7ZMobEHdvX
AeOtF0h2lYOVzwEFIpxFnzDKV5sPph2ZuXxlbM3v317Y4fFOJ6G/ZHP0+Kg6
+MuNJwWQttfbBESlo655/dlQ04i1umzK3uuVr1gfrg23agwJwRoQLHR6stKP
gKsjGeB+9uCb7QA7qi17Gt6xdcyPAWQgC2mYBtRMx21ke46oTCLWbzizcwPv
I0lZheiL38yqJ6u1orlQBUugMqvGV2pUF4XNERsl0jkB9gY36Cn4D8F84GZf
GnUaYDuXaxYSIm+vzMm4GzAF8XUoAkwRKa5VCB+eqYCINiCOZo+JakxJIsD+
vvOL6u9TaHam6gY47F6feeE9bujypW+AorCdXFQta4N87jZkFWsyBQKV9OB9
ecHE6poGFPhI9++D1dwPpde+9hKsWuBX660iJhx+wOtWY6aqwJ0qRVn6LHe6
boWL3C3/YHS0b8L1PVRS9t5SJMKYe3dwZVFTAuTTT/iEQu3ZxYC1zMrS2BYU
rETNf5zgLjz3NV+YXr4ysqqmGQQuXFUR5HyzOXxUcXsV++4YNFXJOlEYYg/J
51P8cqMcbQGdIUWg7ziqAelIlh+XHkQ2+I44epAnaPfqofqXNDo/9mldmKv/
JRtrsACCamo6BhiHidl/mQPehJgIgOIFwLTAGep+zwkDndyZt7wPYQVxSuKr
acn/bRCvb9T5CMsOgfFfusUqPZ3ayHj7tnN97mRrtFX2EZ6GaTjxJPU/UhsT
V6i5xomeAkDBSEOSb/s+qBt75U5Xz0mGj0LifXxAx75xD7cVo8Z+xCTqS6FS
n6rdr5SI2mO15Ga6XRUphGR4RmaeUig9fLJyySmgCEhouQW23glZiGXtfFvW
rY+YCG4Cx0xPayT/RrPOABCXRzsAqmepiCdcAWyKUZeIJ+envDKvBYSYBq+C
xYrTK4xO6eNOeDUmVkcw2RjrQcPJPfnSe4l/P+stIg+Em3b7TFf2jMNmCSqQ
I0gpE646PypxLTLbKJ6kpaa+fjfQwj2NKlHX9whN4I2Y9+ldtAUZ0Ig2SiFj
IWngKIYy3bsIXAF1PazqAK5T0qg+lYsUr+XyTMtiwtkNB+n+D9BkdRcuUTJ0
Bu3YoL6VETBzV+Y+8T6X4DVgxFwwLvfeOk4UkY9S22g93n7oT0+uSjNlIP/m
OLW6zgcq+vFnbpy8U+Yb9IyWNs5+/ih9nFn3RiG4G9yY72D3ImXIRZ84dP4T
B24PdDO2CNJDiA81A9C7BBGO5fZB7/aL+x/LtKINjHnZTC984mdyTuWmPGXq
bw5AIPOoDPaFnUf//Qx+4q2+enJlLkvuszCJtVcr9ZfV4hw93AhBFnbenCE1
+gTBe42eSRw7aSTSU30Twwv7Oo1FXa3zDjR9zesj66Vun3ix0BuW98xbp5kb
iUmR9Us5Cwmb1trkTVSEiJkWcsd+drFervhzzvrYvbn3fBBDDDA3dYPeXPYG
1L31EI1d/Axs714537/3GDlUyO7M3uYU0a1cnCVMzAqSd1EGmT1xwrLQlpIP
u/BKSjdkq6sZRz51YkAKVhS2FVd1sVQsWuNbrGC/Dq1U2rCMKmw5+aNTnkFk
0yl/H8W/b19sXrlBog7cbGGZ/qv9Ylvl9iZFcdPO1o1Ur9M3taMaogjp+/mi
jHDnmAZVDoHEM4CtLkE5f52ThhetyKRD2T8CjNMLsgMDZylLl1zqurzERY8s
mv5vXbbLjialNrJzerSD5xh5KUPl4M/XGsHpWumAUu1xWQAiL+x6y8Dj6duY
ksr7nlSbUg0f1rfMe0uZ4f4vUhrjy+oFBQ55ouUALAdBDHILsKwYJGdmkHTf
MdMYYEFdu4pOKX0G6zq7U4asAVj/iVfjwlJg/DaT6u4COL7/blzUjitXIXBR
qrq5lWmaOFcBF6RooFXn1Wjhc8dHrfb5YepHoblJdhaPNdP5zkFzuzjSlVm4
lacxxU1c+ZA8lnXwtJrcar8F/89Ccxsr7hujDZ/0vl3IorejOwcr4OIDHDX3
vh7MSOf3C18FpoidZA0Nh48xIMNV+O8A77ki1TaF+gD0Ndm2MUaet9z0rGg1
lRemfpFSA7JIt4wvfWI3i6UqaMz4utyWz3G0WqfkZl1Kun6fUYiK1nzVPfVi
f4PDD3srD7bt7lwGyuFI4/XOJToWenXz/pFlwrRhtJnq9VpxVt7nU33Bst7s
zwSRu4J9/pPdTrBnUIc1xwMhsEwXOQlHplUUR5PPIQyIsd5XW5d5DwZT2hmr
iEgaGZRHz7oNaHRyDtqpXtguhSbOBvPJ5DfuK7IXwFxb38PfVRLVCnE6byWZ
RmEYwj6h/a1bL4xFCguzxWJ2/N07vlcYkZPppzt/tERjqSHN97O7E9JJUlhx
FT2X2ckUBrgwD9+gjd6AO5+iImW8eAvlXbzLIItigi8NguUH+MPH+tIzV3vN
AJ6EQxbIwwDS1BVpUG5VLvivPeyZIUqrJghokrWzxQkkaHQTDVdp+NGtWf5l
fHED3gWipGWZS7CL3+NB0nn8gt4T0gK1pCWAFfEksGzc3SKuSPMKlz2TpQEA
Zk6A2sfdgsDLjl5+uAjtU3+lejBPFdIvBdTv4B7SvCSFFQ2y4Ojjjsh1UyL7
6w8j34Tezfv7IHkzzc6dyxVLWwtqBilDJdjJi+pfP0eJ772ZNd7Tw9J2oF/k
eYlylziZrpEqyS5ctOQ3UhI7w3aXJLrIbkBIYrbQ8WbTFdVIDEqJPuO5RoMv
VWjhwYJfFNmholoDslQOq6JHfxp+dkv4S1RyeW76By8wE3auCvwU62qbGIT6
913AMTs4JnnsZSABJmUSeag9aiateTQHmK57Kp4hzw2c+kPs7ZqI5jbG0b0G
9NvvWiLIfxhEu1/wSBUArnLoVzbdTMbAqFJtjEuu2MnhsQuAhNDsVVK9AD+E
TzV5xcgSlaumh3nA0AwU6oAleu3nUQhMIBiNepqiUSNGEQpJYrCdSSVLffQc
QMxqka2283xbDH9+avbNa3EnMcLexfiO3E4mu3zwnONVzgxIf70up0VJvuTX
C2txucf5Gc9CRMTsZff8nQEOJk0cJyLbqhDo6gESgPYjhYbWfLxE6CqZvxkX
OEd1VqQ04xjALVSPvLIH+3Njop1dsfQnBPJQDrJCEHiD3/QV0dfVnsz3zyD6
fqIg98I6I64wYwz9Fc2m4IO9pq9uASogMlBbmah6bpCTUpWXWoki/N2Z3H2H
o6R53blGrw2UipX+SmYP8+EuEl3R19rU37UlRX9RpauvGvMzdEypNWaZZPuk
7zIoK90Jxxjby7dVpOYvZsgWkOUxxvKb6qPv/gN+NZ/wjvz/3gCGa547G6lA
w9VCJKTm2JZdUWXs7yjNnzXjmaWzyGYVal2mFkmE2pRL92uxG0S32PfcnkFl
ZtWTmSfVdAraRY0Zvtki/VrV7qeEWIrq8JgZtoYXZv/QZOqJWJ2xDYAajvui
f0WI5Akb+6lI2R2rx2s2Hxkh6jiSFahyjyAFxkti15xxfvYMy40+b/PLNQWs
ZXi3pHBZ0AKMDsUMaiTWCrgg0Lo1LXn081rqrSzBFb+Dz/z0Bxjocv4veIqH
8WxgnrWVQmbxWAfm305DrQh0mhWkPrtGWNcAZzame4cZ5LOM8E0CMUU9TVdb
4Fk+B/8LY2gWv9hF9XgqCejeFEnQV9y+adNFfHxrtUQ+8TQnlEnmdf+VfUbZ
H/JaPQR9lPF+XbVtLK5ybYCddQkqJnhAHNOXzCqK07ZJH84hOHdWndseG47t
uMH6oB95fQ7mLsVb0Impw4X080sq+5UXq8NZqR3nsrubV0E34N39xIInVY69
kxRiG0bztUXWBGAEjx4VajrKcV8b85vEUAxiPZkj8OlYNoCBKN9KvuvdIcW7
sL+uu8ZHA57QbnpywvCo1k4ZuYiwcSo2VLZb+++E6sGCdzYHJrgDbHnEj14N
4mAIHH8m72ZDBPdl2QfDvvckBwRxpgcW4TdamiIrKTPnrCyyQeGS7AQckGan
dCnbQyAFV6MABw5JXjzm2yU0gC1L6WCK6YAw14H7GoGHdZaUxT+qzwO7dVhk
23M+D63OYKnUJO4ZBt+pkuYiUyB2VScZ1VKsbqaKiYHX3rlCADFiFZXyp+0A
Jtu5WMPGLEIpkvVCaRbvsOz+OZfY3vWIPFyLd4mIhaVX5Zkgaqa5q+uAKthO
9Q+QB2qHwMr1VFD10QslB4LxH4TmjluVD3nih28e3eK7EEq3oz2TEcSp5mLH
JR32HQbFKq09nNCovGs5jUd/8HjonKUcE+OjsFsm5ZA1YqzU8ujelV3m+4s5
9xXznbl/ND2vt6QZaDwKoBR4AJ1Y71+eYJitGDlaTCyMVyV9ojtzNOgy2Q4x
dNtdZ/LbmgEMxUIVu1znH+gN48WTnD9TVBBhJmqvmg24/AUM1/93ToZgWBIp
ULQs1lbV3hgb3TdIdvE9+55N2qHZDkXoeUL2MCu5omqjekkQlQU37y/Q9TyB
KKVzCjUay+xzpOT0ZlmE5psxcVAdFxsSOoXpheXXAR1UOUQAW5XRRhSe3LdS
MyuslmMQvJFzD5cbsPMdUyV9MGgmaQSr9HCdidhuyYvkYw99Jd2D3dpAbMs5
+0oYoohAiO+xITMfv6iztMP+1F+/ZrwBibLOv/HfN3QXWqF1jJGmC3R1vxTv
OZtPbNnsye4AVXoKI6wSxtFgUhOto+DufvYFfVEYIbwT+QZJo4eLBRRbdt2j
e5F8JJrpCe0MisDM2EqKXvjK7E8Jhjdrx8lWnatMw60b1k9Z7MZ+0N3lt5B8
hZLuX0Np7kP8MtHBh1s0r+ChwB5k7lsVG1q2d/6+DA+OOa1iO831GBmNMARk
Kv4KJzfc8pRAvlvK885SnuRRspCOltownKFchQz9vIfugnpchGigPdtjzG2J
pMBr2uNlSy+SfX1rkHSh7QT1OqgKoYZLYNzCl/Brmk4lty8tffa0I7UPCXNQ
MHO79b7V2F9832lNoGnh5ZVwh52Sp1JnsIQbFcgTOJjypqYJszTM7p20Wu19
gQUYgk3la3oDv7++SHfOpsjBEnkXyNSYH7YQM74GBWyY3/aaBhSeJhALf079
jIyCC1zeWO1Lrx+8dEsHznLvHg3s7IkywIjAAxuzc6FMtnALsI+YYnJQ87ir
y0T0YR+rbT0cWbaihJiZRp0WVRphDf8zvHHliXW3+eRxpDdJnjHDP+PcF5En
yBUDXIbB1Z+cVnvghsDA6Y4tJotrRn/hmAbwnbzfscgkBj65tGZ8D7d064hh
E4jW7vRlAnNwSJ1+nytXBQaMfdXyDBnLZLPBSWqE67u9oOYQc40sdYylSBez
hbwp51BMBCWmJ1jc1QLlFWUET1MtI8HW6tjWL8AKlamZXF2Mnkibvr3qdw9B
pLPn0uYX9RZqnADb8zMikg92jH50FBd3Ab2tyOZcWe23No7tcaYb11UQZ9Kr
KAHM5fLRTwDCGgGTKDj3vDUlEVLSV1/aCCe6RFdcitr2mYrZ16XDWxjh1BE4
9OyJ9KpNktUgKX9ohlmiCL2zKRs4/OqeForzKDAiNAg/F78ju4rZ3w0DpX67
4H5TDWi1AsK32IjxLHqH6HVPFKM5UXfNyei+9w57ZNYEZySPAxlehy1La73y
jfC8PvAnpnXu/Acaqj2x5D3s5aR6pJESNLPs9RYIe+Nae0M/r4aJXWBcabnG
bSi7LkpSCCTOnc9dQl0St0qUE486ECX3muTBEwK6NFeHOZCu6CFowPhzWe0F
hmscuHZTVwBnlQ31V1I/mo7iCEqco0xRkIop1Hcwqze2eSLUvfkvsk2paCGT
3Tm6r7P8SWk8kDZqnfkLeFPcAuEUJd3/WDaXuWkJKhdIZTUpcrY+gmsgKO44
SfSzLftcYN4PHcgo+bV0EGrT5qfzwyyPigpeBeKQSgjQ5LFgsEHgjKhwQCoZ
G58SAv6AdtlqwZ0iZZepjhAcUZ3wSUfd/FC0LN3Wl5y5DIuGau/4+LNjhZ33
5+8j9AoOh7eJT7ENazagj3R/Rq7ZhEorSBJDJvv+rH7Pe5aTgeZ7sUdGKVhL
F1C+9FDlG4J3DrvHpK5w9Rkbi1Qr7S0bTyqUe7mdwQHxvGmNBskBOl4PKMIW
M7+JgFXLtagMXObsuZJ1usP31FWFzk0K8ZuDwTpkojzCZqjBrXlp4ck6F8jI
Z9i16fTr0uGYzpweO7ecevlQGudD9uRGFDk/jUa74LicJEXLwoYj2/sA5S/V
reTLKhkGrVTCREPadeNRH+76yJ8AELPhsW/N/p4i4q+0OiZ3M2hnw9TPB0GV
n4wxAsPotvr+2y+es6zu5yNPPzgIQTENgwYdte7OVhmt4IeBl0AmpWzKRSlp
p3YkuDLm6G8E1HcjNYbR5BXIF4/Er483irD9KQXtqW1VvJ19qaB1OJx9GQae
Gd2gclzx7Okbx0Fq1E+KWGOPnVo1mGXGIpIIEujpZ8yLOFkua31h7vSjM1I3
75iob1ioQ+6npeqS1a39skHeqrsMu1itee6d2Ajfp2Ur/NVUeD++Y5lgprfo
O28dAzm/Q++0+dnwmZnxCSo2N2DX8seUMr3+LrF71zB+awml2zZ3JL0NW5Lt
+eNWgmmOf6uImGiEyMx/2nGUr/J6REeQaSR0DL/Vj7X/an+lCkHyIXDL9Bth
SBUTlzoBmwvAmO5/CLh6jXD2D2G4XWklHf1YNsft0Spyg5xi6ca1Zcp8dMdJ
xJFXrMI1Yx8REfb31nOUFfpg3gIyM7O/3zjzyjLjFRLS8AaM+ShJrOr100q8
po3GOwKBXOSfBoB7hID8gb8v3HNJyd9fj6S7+Gm4vGDT2ZS4ji6JFJZB7Me2
MlGQTtk6aBLBQUKwFi6UMRpbxVHVTv+Aj+iT7t1dEmCfQUKg+ez7EKwVm4Ya
RBez+q1oc+jBUJ5r0oguga6ps+hB7He4xPgBCWjFBGbUD1mHnhEfH94/qxCB
dpZ0dd8EOOhF0HXvbRropwarIQaaSVjUR7PZzdsns1p9GzbGWQNSZ44br65w
2KLkCiy/vjogZEdi0L+1Bl+ROztJjB/qxC7BFEv+vrK3iyws2PkIi+Cz3P6A
ofB9Qsl9AHURqu0bc0hncgHrLfH1pz1uUUrp6VDo0Tza1Unx6XYc4ajCVf5Q
Ll4oZJkgtlin/cWlqi3NRiDRfhaODY77LMNUbNQ3IjutyaiWdm/gqPzBkv5z
sU8WRISYU22yotMyzWlZL/AbxfsCjGr3Ubzf49LnwmQNtuoKGfEw2Tep+Jso
o6fZCLyWaWcovYmeMNAM6V6mofovx0TLgWvU37f7d7yZkGPevQtojTzb4ScF
D+o1srzFvsdxI6JFaAxvU6m5qsufO2pRGKuaBQ1JiVTtZMWfE/1vJ4hipbwF
RvZRqSn7TTZf6yuVK4pDTJUIgSvpCvojucPErd1Po3Q0QKvl6qJyHE5XaBRh
Ug8hl0MgkR3b2E4kWJ4nkEk9sWuHFijkGUF945QehjsYZI/fzhNaJSrBckTH
jV3eaV+VxVHsPPjUG2xHXkBQr8droDKDsEsx5MVjL2RNm2FrgpPZjP3UF5Nl
f21Nud+vrMbdC6Q78lJ2Yqi3QqHD8RMBB2E2Cn16v16jpm7ZxrS0KHw3XlI+
p1oMT7a03/NwK+e5GU+vMjaLdmesCticM2B5LjQYHTis41TKB4HsUnfIi2Mw
JlZCew7uVaZlTKt6zwm1IxJhlVf4N4Q3Xno4ULqizWBgAquc/Y5tSgksMHVo
lDulZlHrl8dx0K7bV7m87v1CC/dbdrf3gpas582V4ol3NMBTq7G0KpN/Df+/
hwrmmbJQnqQeitxPbbL6765X497Nv8GIxKsBhwbfrKkjzZFEbSYQj7sCNDWX
CBPDnOTHOAZUkCkX67EmbGkvMct1qhvx8aMTn2YNkyDBRL6aLIdWr0W5VGK3
tQmtNY0d+lE+QFzk/iRyqHzSdiqTe/4illGheT5DSmrVCh6zBvczr/EfmPAZ
j03wuksUD5VPhpY/P895awTU2/0mfQRUEb7TWtX0Efe7HfEITyluiyEZcYIq
olhBzxYl0YioaftzxfSkpZYTVDJMsF49oCBfqh9OaqmoxS19rT8JgnSsZj9S
MDdBF0gBXXKAI0uuUE1Q5pplOMDsIS0BmmZAQA7oVyS2QGGKoDWVfRkCcjup
3AvzO5TCDyEh6VoPb3gh7p11zY+MRmLa+i1ztKS0RmrZzQL7c2Lwst4KPjG9
lEPZF9l8NlL3wrd192YI9255mBCHRycUtHQRXAzMDSemv4GR6zp0WgybDE3N
dxryev57DTD/qhNy0EcHqOXNujceVwSGZBAksdSxQPF7a/TsKMbqylSTNHJG
r4ZMbF4AfU/YIL1NUhYetcEEAjoxt0GWUxC3GPZ5/r/rYFkwIUy4VguCnQhQ
9+QoDdh3M0BsFL0HItthRfruMUzVbXVmD5jjOpUvb3hWuourz0AD1V56Jc1U
WOmgWGaQmco24GZpzrVY8iDrgvW9VTaQwOCvnkI94HvRUa48g9Usaq9rsGX4
Raxe/aiVywRbHqJ5Mv96ge9zRpAGStQiFbI18G1gvUpAGziLuUizBxkfKn//
Hq/aIFv/lu9v0UTtYlhTt4/XH2Zpb8yLj43ELl0q1uFvutvOq7IxTT8l17IV
kvZ1dKo/p1OyIcrcBInAiR3L/1YmpXSxrGlhDRjzftSZXOrv8plI1Hyg1Z9O
amrZIsTKg8eh0fnmwN0p8vWrqV1/ty4Zqm9C2r4hk7KUWuKPMM3CtKP3IWP3
eSGelcWLJQfDpLO6Mp+L+Td+AS0wlGXVtVfrwYL62X+9Lgq8BFWwDKY9wDJW
PrGp7RGvt8hi/vdj2XGR4nTnBBSm/BcduODqX668n4g/pRem+0UY1dg+rfE/
NSkxlp2B73ESiqs/z7BHa42S4Vjhd1Ev2sLEbKs+X3+5T1COfi45ml90k3Ak
GkqbYFYQ5siFwpc2BvbVFhkvwnIwJNBEQfDqQA6SfpF39tcwwCcoXqVjDly0
JtPACkNBPHY+uw5U2w5EqUlEh027v3ahOLMRQw3+SzpzGEN9x8yiWa1JD4sh
kIQNNR9oXD6S+wwyIuKpXTWqaWS90zC4RPKwc1CCRSvWu0cMn9crHMep7ATU
eH6lg5GDCW5JC4R6gKa/ltFaSsOoHN59NO13h/HB6iMJq4OVO9BGQ6UX9Q3q
Q18u9JNLVmIPQqhAjE8G3cjH2yjPHudbMy8rppN8Wos5Fnmz1q2OTZkURo6J
jtEpuDzq/Yyp6oFU5WHN46iGX/6XaycGl8GC+RyBBR5QS0NBaE3fQjWALTLQ
B7m419OWFxl+6IuYnrwDNv/KagBNf8fLB4Tc3xc5Nec18Il523rNHrZSZUBs
u9ivFqdy58Ho93oLfM1+3Jyyvd4bCm3Oxleev7HHKsxAT4Cwidi2QK5i/9ph
qLzFeihBTz8zVD9aOhJsQf9tq3EbECx2vb/3gdtyz5J5Ii/OWce1woa5VxwU
6v3Y/xVx4mflA00jwWfO089agqUI20oekhp84DhlOhIf5ZBF05zcg9IQ7LAO
efSw2xm0Y3YM7TPS6Fn4eQdpWJq2UC/oZZInUei7sKv7W4ruYH5rJxZqcTlo
Osnz74YmAuZrDvZAP+3suKLinBfdsOAHW3K0dTHieu2w0nUj8jwGgSjfl22l
Kb8/Z1lng00DWp1kZqan+dXioDZ4h04Y/4/yEumZITYEgA0AElKao6xdXYNd
CdXRGOOg+PWOGrxMTqi3wXeaS3cd449tjjLSbgBTWq3Sm/F/+BDHHtSRpeNk
WqRBoJmfsDkKbOCJE/g3vsXXsu3W9a/isvv32rgMQ9EquZLQPjwcF4gSeKag
c5KWQ4l/H1cGxwvi3tIem8qZxjE2KPGBOP0DBL0B48E0MD3mPpyU7OpaNjDM
Qqv2lS7OKpcZMx1RS7vXNeEpKwMIhat+RuX8NvByTj/MXZA7nguuGUiFrlBm
KnCcloCJ+TyoNf4sIkW/sKEDvscOE4pYcNnyWh8tAVJsEQqn0JR2SLxTUarc
tBxbjIBz0fj6N1P9DP+LLu58bCpu4J1LhUVrzp5zkEtvNXL8QvYk9uaXIIXZ
eomB1+F7/j34ezM9EWLoSuEiAt83L9TIcKXP5tjMaSxQIEyg3WTqui7/7VIc
weZsL5ipmHezU+L9oICJxCNiqVhff0K/OyFfZ7iqLA3lAtzCYAbN0j2683VS
Y9gaCeUQlc3Hsm38GqS3jgA3dtmRLSRj1SNS6Dm87vMhSuP3ntthrh2uLMHd
KNx1H34XGYHYswYkNIesErh4OEG1UJVvWB9nvzd6Bf4sRWiif6QjFB+ZZ/4y
T+A1LDz1iz0DvI37K8uOaMvSOWr3H0RViNPKqsSCxqmiaQC9os2qjiXzTbrM
VLBfl3HpVHwStRRDIBwQCzNrpTYXkqfUVbzhWCIySpSAwASshJLxXPSqxYuW
D3IZ4rh0sapTLaCV7vdYkiKqHiSOA/3Hf/Vdoh7jGurh70+5rW93wGqxlnOa
MN++PnJgLDsx+xhhtwqYgTbyDvp3ixVmUbPCkzzpIaIibWNuJ/kKsJdejNkN
/CUshRhee6QJDriXH1OwiQsjArsZsEVqmQS6x5HPE3UoP942OyhUJgcVik0q
6lilU0Vd8CdTKm2X4dWE/oVizZoNn502D9XluhbtmZJ2z8nIfLk7JfW8oS6a
4zQnrj0ceswdVUxj5cFN72NyqEhqRiWQFix3jepRvtl5cq36v1pCbwSY/NVz
ql4lXJiqWv6itcqBOeIQl9aV2UAQ0wblzmpESBy87m5SHc+Ns79T0eluSMb9
fL0qO4JrP/fEFxFgiXCu4ETocywy6lgi6qxqWRdfd7wNZOuAdKlWcgB5Flov
6F1jN+OgeAk92BqpkfXld6wz+lktTex3cLUAt6hKmH+ufgKsZ1B/Djkx4+oO
X7Zx6kRPP2lxpkwrIGs0haPBze+iJS1EG3OQ9yGXfGRwZtA3I0+BzJX5VxzO
xnY6DflpCtM7Ln8brPsgW62xaYfh2XhLYcrYd587laWrhxHy9q3veB8/gHcn
yVu+AgU25fsEFy+rXbUZJ6KMQ2Fk6/5ephM9GhSw1KIIZkDLyGHcuTlvTX7K
i729OQoavFcGlepGbMsfSUe1R+oBtfixYy2imKMG9fYVGhQNnDq3510MjBYF
Ybv1oqZvuIGrI1163ubQ1eR5IYYCpUiL+STnIKYoCsveSb49A5QSpqYE0xVh
TDf5dwvyg/d1AvRj/TgClenFTa90YFVUD1h5c5FIMogLma+Cmp59pBBRhVJj
lMth1RJB57zcoKY0brHJiQBpHT9GgGhSLpjrTLwaiAlJxHXgABrznXzvhby4
AGwbKsksBaoocPjzr//+npKNoz9BTfLy0AUcBlhxjXE5eX5FWqF/BXYtVjmw
r2Gvr3shrP/gs8IuW32Z6C/t10hgMe7fgyYr9DWFIglTdnGuBjePAhvY1zCM
TdN6lwLnNlZ6tNUvEtUdrMgn/XGwKun8aI5g2SDAQ3WOa+j4RrwmuYJm9ldY
5Nxj6lFdVNY4U6dYk60rxm8nUkRvFHZLXSGYlSdI2XXaMRv6tDbTcvUXokVm
XPiyZ1hGFSt0cBZeFlS5yIGjNKUrSsXHUjzjeJniP55nKMkEmwOCQVSaj3Ia
z5GVGVDcMPca8IYX4rf5H0DtX5WP5t70JHZ5Snx9gFssg03+lt+CRFIrZ+yy
qE3L1pNEmtrntmMAYznita7rjTMsqMamysYu+HSuc2hIlXGDE573XZ3Oulf+
AUG/j49ga2gNC5C4Mxg1yY8O+FZhchrn3FtDb65YZfAQO0+6JNv4Mk0cfF8g
Rv2q6XaTFn2m5vi+rMwtj+pBLVNi6FGfQclQnXToNc+qIIF6WjJIU/xp5P9U
bn3Iy/RkbmiIgzcOm97zoyvFkmOn7hOLZbyJD9dmk7aSrPjGVzd5lUJjrinx
ayBey1mUAUTVy8cPXGnroJEqVqSWZycTTI7IMLvEl6Ls8DZozdz+QXMgf73j
KhCKWvgm38WQSeMmTUjvAFUnKeiGoiyvfultW1GazhRIPYBVGrUAWWlC7X+8
pwgRWJPjFAgGrpq1THsSqLyR0pXMGKLc2FZbhGzyPFz5OrVC9JwPNMjIXjuB
eHS5Md13k5MnHMrhISuyOAs+w8SHda3LEhZf3Z3UWLUsNQhEJ05oiD600HGT
g+comTGhIJW58/N4EHsaz/V7puklpxuv8OmQvP23YaXymqJxY2ZgQGcJ0k3C
Z5SPhuw4/1VnRT7417KPavAUIMtczpbi8bFNIs/7X1emrKnNYkyVCysp8SDH
CtUabpAgNG0YopcCw/p1y4+5b3TECuXdFd9jBK7pa8UNNh9HRQGmXQ1GURhf
ORqsuwJb31Pa3ooU2wqLOkjGPjwOGLdset22vQFnkMy2DnLaYj7yYHyfeNQy
82tuu0sJMsGneNhuYdGxBxzXE7/Om+zlCNkHLwS5x9LPM1uDkWVHh3YBHXAU
hNZq8Y/KgnzpKRAWkci4HdOoHS3cGKD/keYoxJVRe1j1+rlVZlkgrQB6uEXB
oxFcXFuwQRtG9xWE140kES+oDiGHru16zqj/gM3ENwM1BJIMfNIgsSkOPgIz
4dxT/QlJGc1tLhKWMdz4Ksnn3roXu0q6m15UAVAKDPkfJwm+Tzi8yM1eJxxt
y/GKb3lfvY2As3jrX43j+knTjJdJmqlpy4nNLIDEtMnb7z6Pz/q6lFNIyofN
+M/KMPODKENgcXyOf/XZThMYrdjIvVUZ3N7pXCcb87kVbsVZ3s6q7rtbDAhV
y6Z1DRv00dWHvSItWZuJJJiol3q/III5+MMD8Vt64bIDXjzLpkdricFMyCkD
Eo7jw9ChTmIgiGDCeBIxbMiWGB+F8LRHZnc70Bu9J30IhCmqJmbZyNu4xAZe
LsRCbdfIrtjTL4BZ0t2Ph/96KSSRsHkkVLAV71Wq3Rjq0C4awdqdKsNYuS+g
JVjd1VlcLcRD3OiC1au4C57P1ALBjdB0RjIiZDr8XJvlD80JH710g5U/ZXnu
W42k5Fw8MKbMtl1x2z09HrBmtxKHTdk+F1kJAZ57qcsZO6YiGtmofYQXk7pK
aaMR0ITRd97Xdc2a1iYOve3oPLrqdbn2EgeLjUw4vsAPknnbSykAMIqMuGQb
hLYEIgwiy1v0QvtQ1b1RaIfySZTQ/J3fbAjR155VctNZpSong7manqjrthwP
gLPM+rJIHSoGyPq8HLA9jJYrh5hV6jv+Zt7VzcwJtGS0Muw8svW/drjpIbHB
rtuy2+R0o+KSaNQP4YdXiyhPjrkWZL4J4VriaotK6RXYCDDOejTGwRkvG57t
D/70aQ/uclJ7TrsMyo+/8QECZhau6lxodXXYlZs2NGwpp9C1jKcOhKVIBb4Y
JLgqVb4l6qR5PxCGZJ2WOkebRBygOZ6tweuS9658gzJ5tJycgZqVTjEcWapw
rL89HjseF5q7Dc+yuKmnw8w0QBbp9FS5S+LzHoJm+hIc76/9yDyTVFqiuPws
X7uG7GpFTwI/9cKRKmXsN2pBj2dQZy++YTPn9sP2gplzf7WK59f0xYWTAHnM
L/c6eNg99YZmAnrLf67m92UBRsa30BTauF4pj85T8OurHhgFw57/XrT1wQFp
OyXWS+0NAl/wJjaYXS4XJCc1jBo3WhAaoFUwt2FaIZtbnMknjlhx0t3+2vTU
E2876FiZPmA2pAcGMGRd52zNhTMxYQjyB8l6aPudeo2GFZgBLxKwBt03U3sV
medV2tsofavaYk+hjaCu+2A0HY147KSjBL5bGFtqQrSql0Dmu6RQifhE7C2w
7NAeV8+v6i4M+ptWJBNI0QFL2zYzVcAo2UPkjceDxU1BHvU9S1pNCy//w9pD
9b7efrmuxuNgftBU9I2Mf+YX3Byf0JCmKONuC+SYEjsZyxSH47Su43KQ4kKu
CrQkBE0Jd7WZxRG69UzxuKcPWgx+BUIzCf26ak3z4qwysyw1aGDFZEQdmFLW
aPeh/Pnk+HBW73JNZ4mc7LOPWPKvvVnIZtHqd1IN8v40DvKYbHa1/GyIYDUR
HRuice1lePSt77Rz6JIFcbKadjcmIvDwTop2nosiObQK9JaTUvJp2H2LIGFY
tzflClLUGNLTQeJO6DviRLBJDZxzRCXbu/mygREKw36LIRJUXDFZvsKVzQ08
TC96xy9pCh3MywKkPfaJH+IgJqjXtqWJNU1LkbplI2DB5Jiin77C6AEJW28S
c/hTYyVemd6KnO3PxxMRQW35rgFU8sb/3AG/WJpNpceSfYCqUhD+IxsMkS6D
NCZws4BQEIVnW2g3ArMZdQK1vwHXAiZ6Yon7MJgLmGIwwfoEmoNTPtL37FXS
d8TfsutMJ1malzEseTuTTG32Vc0aFsTXLTGQZxBkTRjKcZyGwUbRwWc4BnVh
HfDwe+qCBGovA9OMmsdGfLnsvUuPQf0zjQCLrJ5VvpUaPUHwLwgRe+NxIKEg
YrlDR7KW+SfrD0W439+kvf4V3KB1JFP97tyS+FLvZ470Pnrh+ixB2RfPIpGD
gbYxCr8deFvJWawPsmWEa/GvkbfVG688FTg7g0hDiamtX5lKw6USDPNKqVmh
pM7e73nhtXLTWAs98raBm1jcNCMRZW93C4fauIw/LJOmVfzUL2JzeAN80HqH
mVuYF67psp8bfrL+92ZiKIVK9R/T+yaLAtC09UWx9s1MDp/Cikh6W/lnVUzR
r1BYPT+NO0Ow2uD8NZn7mvw8ErbIU6+73dNFYAr8fXR9Ckf6UbhlGb/5ISFs
DrMS5YKzoVbcywlrCrsjf2rxRFLjgIsJh04vXshompooriESC+dODayTE57O
u3cdmotv3kQwkO3Tr07tSJIytrk1m5aKGn0fAGh+0+4RCBbVtFmryRz2ojd8
V0YtFJDcZSpwVRcGD5EWY2EnpfDnTmPFxcWdg6loBSM2ZbvZbZHnRP9X7Wc0
eHKP4e/OTYNWiIa8Ds+iJsLaKZIgQDwKrw3xgzn9wXxORVOmJ/y8/XpR0lHp
qP4ayCyAwi0xggRYTyJCK/Iv3UUrZKQGQ4JGdLt/oaMfyYH5vt1EECECLH1Z
9o93gHtr+o4z/DSeZLM0FC4BWGYp0JVdCeYlR89q/qSZsCwmMZvEKCvGEGWL
cHAydh2koQfY6RWvHbd2ae6aV4bUjWq/v2Iz3Zl1M7Pvm8Tbah6FB61tW5cy
esrblsHVJqjGIfByuNB2EPsgx05VVIAnrlCfmMQSj6bWrI8P1q2AT69ecbSA
cGNe1C6Jgql3xa6rR52XsUUcIPAvGZQtF1K/flNPILyTzjqGg/Y80u+yI1Nu
230rH4dBPl3nMP2GIhbD6PI9qhd4DDaQdMz4QNR4y0/fdgAxqq7oT1r9v1Cs
tdkgl52pasHNHdK6ljZfIlQgo8LaX40xzthOVc+E6iSkM2WAqYWZlwUan0JO
TCLAXm/E79rIzm9FpQm21mi5ssEHaMVwaeHZNQ/3E4UaOviOtZnPpaNs52cC
Ymm8YPPcCHanRy8lQUcDw+LU47NuyA+yVpqoD28vQ2VAq8ZbzLFZZgND5sq0
D20rOGwOfuc3xaF4uuoeIabf0wBduoVitqEcLVpfm88x1a2REIbBiRo0S3ZU
CUSbIuMihdPfrytxYSpqR/EE+Tyx8T9Lyc7RShf30+PSP0YUdTjYh0sqteCY
4yofyRNktzmhr27ARARwXZS8/P2yd9H2pYQ/MHnE/omT+dYSGK1eAqSkYIGL
Z9ehC5O2TtbDS90ePsNEKjRF9Q4LBpK1R9rLqj2gPfjw/cht13LusrlNzrix
0eUGoO18x7WtciyePbpguROmiJuqbPermGqwjcm4q32HWs+exDRLBPUzNKAs
hABR2UxLr4OH9aMXUc/wKHH0GhMntQqBcCSHDzcYAgfSWBVyEIxAY1X4kt21
x8BmPNjDiFF8HqtT3iADGRnl6PHnucoRod4aiB982vCuWlUPsVeesZQ1Ne0f
fCc762Avfvmd09ciOEcVLAh2URYnDCDVvJYAr0xGPTrCRCA+9loq1ZQClnIZ
t7T11cBDwTiK/sy3IF8zNSMjEaCHWmRg1FXY3dDDewwk4DXp821DKC1EHp5a
qS3k+/Tcxx7sS9XhbChwz08f/TBJ+TFB3yx95xU0bPVBom/mejEfPnHWO5MP
+1B8veruYMvLymyy5MwZ7BuGWac8uPpskAIST0MsJsAo3dhO8/LWtJN5CQlg
tzN3dfdtUVdBNnx/LnlkrmVlNbssC1kFs57LR84+bn+yBQAGWAznliEeZbJ1
homjIkrsHvhq3AXqmfbk0zTt6d8gU9ARhBY9PoJ65CSorJGH67TQMa5u82S0
BzKHwaWTspQChuwoXzTM3ORkNOWfMD3WmQT+UKjrHourhr4FzPz63YkuESf/
DbFXwyWzQvij/phuf1bePfuSncoavsH2J0ht0T5c46458iNj2B7D88PhydDI
x0BcDXPALHdOVOf4ushkoa559aiU49cWYpvSQRfNMpOwTwhFcICOnj9eU7O0
bkBrrKEyB7aRSfrDUp3qNOWNBDz8nRPUjqbAhfujuckT6nDm+IZF8pLmbwzv
vfjHGaSYXIiBT7y9aY6LIOKC7FG/RIbxBwCGTTXDHU1kgN5LQABPAduCsNQL
Wvw1qXQHCK8ojxoMsmhepLNcEAdQl6ClBSZM8bnLHi37qh5PJ0ICr9x2BI5F
NqhOAipZQtvlzzEgx0WXF4xm5Jm2m7V1/7wCVutlCTpuCJs4Np2aTdw7AAew
LsCRCesGd4rbzOjkDK9X4aC1bxO9+dBeTeOwzbbs/CGJZkhWIXRvbQ0RHJ4M
FP2bkMi9/SfSinTcuYIdqPt+kSHKU5XhmqGAOUxzESjVQ9CXzp4Ph69jXIaj
6tmV4Ass3sNbv5sKwtcBo1+IAShpyLlbCLQwEZSdk8OeNsgw2O4Z4vS6jwLM
9znotlMMdfOs+zErC6skR+KNd1AEi9J97+FbYgUJZJYdaZ/7Nmg1oZVTz9kE
hBBruvc3lxgQL+4tJORRCR8pKbMzWU8EKXtPylPwR9fzHIZ012MOiaKAO+dd
WXv0WDIhQqkOb/qQDOozwcBdjdY77PFMBQghqrAcbuDd9o1AZcnBJvkjrccU
MrGYztOlsYNo+sjRpbdg77/ThOIt9e6ReXDW4bZht5uChFm7Ab9JKx9GkCHB
39+Ek7+HA+ArfFl/7KgMP2GZaw0nqVmjUyxMWBt0viOIfs2NM6JbczWytC9a
rsAog1QPkN20MewIh9Aj6tEPyfGRgtcOTKo0bLlg9JFVI0ViVlNu0F9RqWSh
Pt7Erw7dXeK45IDgB3Q0yS0uosEcwQub5uwx8X0CvQh/4fuwFbTP1qtuqcpv
GmPk7bH1iYgBkVaD5s/IzP8/am2mnVF4msdIKGDzaWG/FAXLp6JefxZwBebm
STpy/HvASvm7pHhfD8bdUkdBsDZZDngS4rTOkQsBjKTtLxVNoraAILaviwQO
XmD89EnZUPzyCbpZb7a4M3UptclurcLdRQir8nF0jcq/+XKDXTNvarTeiePZ
z0UaXZwz4++EaArehHh9YUJyPMYbLd8csAG5kLzHynW5/dblQ/QGYxcVpwf4
lcjT4qSnyyAY8qc9KLwUIQVAwGvovooB8ryPCwmNan5D5jKAa+Tod5+h/O0g
aHNlgwE/ljYJ7OGqTRSTKi+Swqz/hh2Tgbs/wH+czaExWkAWUQAl8h7f6rtO
oCsd2CziI/vjvZ716oK4FkgC9o6TP1P13jvffOvntBGGxWa5T4c1RoouZZuW
2/tCNP9XFl+YETrKLx7dsNtc32h6XXvAvBZPLlA4XUuCp0G4KeYIAoCZ/9Ij
vJtwjj309/Wh1GbA5mnlKzoTP2GMBUTAVu2L/H+8ekW53+rYrjcpPPReMGdY
uK3/DOHwz2owbY8owjIfBZDQEkwBUGVJb5XJVOMYorbE6vX/pCcoqzfREMk8
tPaPqMIVn59WYj4OugIvC1bx2EZSjFp+bQxvO5W+w29DpSgu35kgjYX40vhH
t4q8S6rGTWbJkUEc0tfVU8Ygc9K3qvy1wCrGJ7LcHhsA0HTSjFbDYm38xiKy
3RRb8BoBb+vkzSqn1nkYViBtFR38r+SW6yW6UHlKZ7zOr+h2kPjWLN6OI88/
6UjjAu2WwcFNYegXXrN6Q6UenXYtndXTWeYk33EjxsVGIU3n7mnFO/Q8B/yi
7XLofiLDpTrC5fIySolAl4MoGB189JeBtALBOux5rQZ5/awIJVWfYZl023KN
bscyf2Yi3ZcD/dRaLM8xdloB8gW/addOdT6yisWinwqUteUpaFCOZ2TtuexG
zcMOQh8lxeWiZa7UV4c6rv/RPhn+RQuxAxSDZjCwtkDoHlywt3X2dpcmM8YX
jJuAV1DLZpN2FCCe0iw+Yctg3LxKcAnkyy3vp1qimPmWSceaA0LoKPpgvifw
mRYRjG737GpPkvClYf8yTNF6IGfDjeenRYUHhkRV0+xer25zT+FoyrEjfKQ5
0t2b4kWgmH3QFcKRn+WdDfSpYZlvY8jredV8pM9xwnvV5xYvhcloNMYNUsHk
US3dEbEi45RQVnogBIk+vCrEq1w8mmb34SUIcL3ykv4SFNM9LCzMFqR4NtoS
u20p3P3o5eDJwn8dM8HqwbgzVUCm4GyYHlOrICB6Rgm1nJ7uGQTBBCxdBrly
q9x40c0cmlfmKXe2MX4gHvZxZnFqiE8j9Ea1X6xYjwk545dzDw/tFgwfaN3m
wOPrxhSBGI5r4g/iLFxAJMcJ4TYKw7Gn26ssTklpr1qqTL75oYBXKh4g6RE+
fd5YwzH/39u2UE6rYmtUIvREvblSLNh2ZyqjiFIpfNDIks0TPyjp0/tq9Fx6
ZoSx/KVOliC8PosX8eJqH1K96N5G+N6qNK8QJbnoLaoYuHf1BbhgP7CtElVj
ukj1KIC+2PjOT/drh2Lm9inUaMe+GZEl6jl941tZohhG4X7Ht3H4as24yopb
mcAoIiTOLW6DsBHRB7cDFoLwBaFYyWVTRQJktS2ocgXnmzWOXS3RGPVlSPa+
YXxcK9Y+6HJqEfHZmmzG2jfX3nPXAjhme4gq1Ti8/ysD0PPoDaT4btbtOMmK
E1P0zpf2LzHw++NKxfvutmlWsoB8IaIlBv5wWo39H7joC8Kcz9VXqCBTbXFY
fePbkHLHy0RBKCeSvPh5eKtlaDLK2abi1ApjOyjTeubhLAmgC6AAA35dBX0Z
R5+RB/hNr+dcQnoxbLH5EUtDBrCvBiUJas1LXQCWuG28GDYL8khADHME1/Hd
QcT3wZjsKFI3KfZ7g3EbYcT7k3KzQQomjrsyHhHpIF2VQvWu5E/4H0jbqBPb
syMUjudby+21k+NZQYRsgSjsarabj7cKb8hpca9gkThpFOVu+gpYRx1cAHZI
sjxtoN0YhsyVnQQNAOI6VdjfYmqwHKPIcoA8he3mDFzI3dfggT67JpOv8VBj
BwhZHvW1d/OINBhLRrdh91eegOjiaPWSFsDbLwa5exKxTU/+K/P3BnmtW77h
VJ+O19F3PoeXA+Sana7uHbvE/anRIY4Z58P3B5hjCpGl63ZsgMrDuPyzs+xC
fl4X0iXLMoUhAjpMB+L6QITdI5NHQNAPx3TSYv6I+91VVRg4wEhlaJo+DVK/
I7UyCsH0nLg71zbi9+V4hiXGbPIVWlPXu2e4bP1F7rcbWYVSmFaMqpNnCFGI
OKMmvGOJU+X+EEvtaUPJobw+FTlDednAWz7zVGU/ex3/3IjHroN4Zwka7kAm
NUNX0+TYj74oIITXjL/IV23bOCmP6KgBb0l5cRnJPt3uR4sNra8KFmVhkxhc
+SU4XOP3Zf8rp9mCS+IRRFgTUBOS2Gxru+ec642LDeFtpljhbifoAx24vB3L
xOS+WoebRTOGrfpKYQrOlp2OY9R8rta3jKnwDl+JdsK3Zu2rAMA1QAyi5ZeU
swMiDvXQuwPJ5RARU0RdDx2uH6HDbHN6TEEH0+8vheiAzYXotZawtqnfKsQe
7kfjqL7CzBl6Bj0+qFIvCMwdywy2HctK0uXC76HcmHQ932kP+271IF2UdjLt
2oQEZpgRQVBO8N0Rk7xYrCPTMAx7eFjpdw+skxJQl0Dwe1KsLJ3nyxKJVd6F
w0pcm02O2yZG0p08ymTwAcKDL9Apele6YVuW4wgNXDQNocsE29gm/pxECepK
A4HYvVd1pSogTo/wR3aai992WFR/Glz0AlVPmRIZMAAHEEVpHAeBe2BR9N7V
Gq/tXnkXdekVfUnPQWJ+Aqg8KsnM0p15qzNy1if4bqeuU+HsfmZ8lFf8GxiE
o8ZiIL9rZ9d+jBVRNnmfcrOZshfDDVl0yzdN+UO2NqmNsnGzs21DgMZcW3vN
4zNWA+D7yAEsNmi5bS5vodFE3j/C9VZshg2N784bY0h/L2d9HwHCFIo+fNPI
p1gs1nJqEZtz4NIBxmLab9uONk55xIyPUtLvdbsEF40ir87tSXgY73nCJHmp
0USRP/od5P8QT1hiH1j+yzBhsK710ZoZJcX1U5/kMZAflTYc4WKKXKkCFKU5
WWjRDPHDgzTT9hYb1RNWIs/ENW6yFJ3DgFjroYwc5zv2eFeFC3vSSmc+RM+V
ntdi3D3NptjegnRWw7aPZpDeSk3i0pW2dxZ0eJm4M7dLOPWJxGGsUXDHqc2V
2IigUsPldQcQIahBu3MzrSDsRmEjFhsuckpyt5iw6C/sFE5J79J67yrWtnO0
QWhMXQbHNnNZM0pZcrgHdgkj5TtPkit470+Xo+mC61MPCETlxPSsrO09uhII
3/DkVSI4MqVH0O7+aJWn6sSjC25PcC9OM/FeMgEG3WQqP+0PRj8E3hYnNflv
+fdURRyq55b/pwO4RLm2113yTHqM2TiN/jCocVcoxn/Pipx4AHoZ+bYBqXDR
pOKOq7Lnj2Q28Py9M/Ci3DiPk6NRROR0e/y/PuYp3ucLpFVfj0pM+EN+Gg8p
rAuBSRnGq5GYiCUYPzWvRApMLKQWkf8h/+8Qe4DIIkLPNbs1Lc+9ss2e5hDB
jQSQBWtKTKf0LXQkfHjR9Caii1sgb8uHLDYhdx6tFzKvocNko1geOmjFSIHw
c1LkTtGeW8rUx0X3sFhFZGg0H6lA5En+tPWV2r5X2shuqTH6y0pa7lbrIEhw
gkNgOOzj2nHq2F5MFqJqRcQcW7pLpy1BFqVrIV28GHNxFi6HodqZ1utTlMO1
g+Plv+/zLLT0+ULsVmlZ2RttOjdujid/rAweJClWeErLgVnsbVI9aSOTfZXl
/IjLhcH2WbDeqnTvx8BlegdDt/G2Fhx8EcwgMI8inxYygkzkDvDLOp7Nev/s
6FIaSzLSv3Gapu+ELD9LPR73nrYWSqkCTSFqo9YRxuBHNqoF9gWb1Oc/FQaO
Dg2UCv+a5Vfy5bGeQD4K5ssOtO9nRsAeCaoqtXjrutFJOW6T+j7h0sgmxE9s
kxsegucJCvCdX8Xk3fpJsCsnOv+YbyJSRh7J3SlESG3TIqkoNyCjUu1KtLJh
EWGwiBnfa89QV+XTgUq1SHlhqYGHQcQi+BjRW/GQ+4Z+nFA13zBOOgYpZYUH
c4GXL1IGfyl2lZJyLiWgruwUx9ZeZ+6H9arave8kZ15QKEBZyugGz0VamUCJ
a+2ydVY6BY0LP2fCXlvl4WxkvYn1iQja4A7Wg+mg6Qa+698mY9y1kW7DCU1q
MycggVptm74TyxSLg7wB3a7BcyqtstuUwLqaV4vO6849sEOP4YfzqK4kQ2Us
j3mD9mgQljYAdDmE/TSX/ZSlp71xbSoVfmS3iHJ4b0YOctO7H+ZyFglZXEqF
pR0Ml9JDSpdAhZIco8+0GEglUihDE6J7cNxRV40eh6o19Rl0CwMEGusT2mIN
aVweVK+CPpkL1+HECevejEPHLvGoUaH3UH7QpN+M8QE2uJB33NkQPyTsyCyQ
yVQKCzD5BU4jtEwoFDQ2hHVGL+eyO+bKVhPZUeUCq6lefTjChrrwEdiqGoI1
f7xJ2Uwz2WdzNR6pYM0Ok4Qw8mUAVNK5Pp0wucJHkeVQMKOMh6A0TUO1P5CI
Fk+1BIUGiLVoCtGepNfXiSRVVt+QKOKh2GVpZ1Pt0Tw9k2rbPbKUwI6cHc7o
tZe+rZf2eTuXqhtaxDbp+0eVfj2KnqIJ6PJQudREh3vs34/2tFE837jLdOkA
5gS51MyuQIT3nMf1cR/nWLIx+QUfvafT0NEhqJ1TrECxX86c/Anr2STX/bRk
rrUSYrXzUcX/urEeOhlU6ULF6HpMyDrAO/PzRVKRiC8PSThwwu3JSgwjdIwO
t1zI5yLBYmmZuqE7MAny90U8E5wrBBUZjq5bb09L8s+2xyW6J2+Od0pApcsG
8a87YrZRNPqhFB8AD160dfmZZG/FnhtXj1sZlZZdzEjM93peYWOt7e1IfrmF
DR4qNfNBloKbi7JJAVpp5OIOHFPrJd3jjkoO/2zCVq6vLTLh3D3pHEQkuFz6
DN6CnhHdL52eOoU5Nwh6RDOd0w8pQc4e3DX7AIAISxo/MqFRQbDvW7unhN1C
MGvqZA1LCHKmssuWfoxnB5lDVCxRkTDzouLzrWz476aTh8dwaG4GHfpCquZE
mpmHre/3g83n6Z5KLYLUZmiDmi4b29zGUyppoQuS+NarUiIze+zDDsqHbyc7
4+xFE/9JyNSFFu4DuLxIijmBNizwwbSSMX3S7ZcqQsZg/zKH5Ks8NEz9r4UN
pIhU0mVPdo8C5BdaIos5plLVzPkPgSIITPD/3WNwPBCjLR46piHwJtMcgCqA
OY/tHczUawlQi5OdNWDFJcw7g8EKNtPYInNuCo/Qhrn9HqHMjF2un4TNYPoa
/QYzffm/KBmXGh2RycroPNl22ryktw2LLE9gHZW5Y4xYzEXI8d6COdeiXFCp
Tyzpi6ZM4pIwvZ/7bYfizMJae6KhVd78/s/7WunwYzxQp36fsNj92X2TWKOM
MsBrIUcnUjcG3FOjsev0C3zd/wcksvDwWZ7UnI5WMnFHB08i9vK6BasRk1Ai
RCij0TbOSRNeqHvBWoZe87EkZSOuea0ZiM6XzBBh1lv6y42V3RsEsndG5tZg
c796ajPk1dnrCjcu7F/tL7qYiO3Y1Z8pZjOopVTmuuXnq0klyWHEilJforAg
hiNL7irUF2kLvb34PsNzv3bR88UTiD/UWiTXLLTWECHGZHedurRh6JeDiN15
9lApvF2sBAX96/2xbj5F0+ccT5vTgNq8qthHdDJp9mhm1oloTfnBw9//XJzA
SWZ3Yliys7Ao/IoHA0oH/PuMqiP3+SP57NzJSA1+4k0sDC7OTzGBdjgqkBB2
hV+EKM2/fGXRTq/oG9PvBhmdaf/0lCw2ES/fCwkkgIgfmaKNEvs/vWUOmeGK
2ir36FPMQ7Jl4GVNRMUtLJW65Fikdr119w0lDjqSRsEFts525as1nKqKh/0J
CvFscDhSgnGc8Uf7e9yykU8OOuxC10/7Tf3p7cTTCfZoqRZDuq4fHv29Z+1l
HstNJvCaHUENDt176pw+HdrkAHquERPCJLyo7lkVpWAFdwCUlUJurC8Nd/Qd
RiL1/vnZyUW446XO2SVr+48t8SPn+Jlj7Wj3jpHkDOba9d/ojE8e/QBarJLG
w5FmBgrDkSvyWMSX7q4uHnb0tbtg1LZxdLlZCWiiV2IQmRyZ1aIytKk7nAJx
J7c5tn9XPGfOkEaSNeUQGm55X2EFA4O4iI8WSdicl1oUyGB6KaXKMr1zRP5I
GevZSYF5B9HoWCkHQTXxG90goIfWmyZlAO3HrNgGfgN9/Wi+mlogVIJOfhCt
qJ6TdaiZrQ0aA5CesdrprfGCbv7bRWs0Bk4FmznzN7JQP+kACSpJK3REIO/y
eReNVUwp4mtYXOMgGVphak5F5a5kB9F5x3j5RqFo3bQNVBCj/YifCUZvi9yd
mx4n5B1yM22bFx7rlN1WsFaAQ2w5q9gznQ+or3LV/wiuEgiNbIizJ7WxfHyD
Ucgne0IVt1dUiYygPtfPQAoGLS4bdtzGKHoC+SNTNK1h4kACRL9oggxWibeQ
DDvWpkfMbsRE+17uisvDEqUEfZAIX/RPocIDT2jM6RHN5YKd1TA/ir+DXd5C
Kslmpgw5gmpdnekgxr57fsJ+39r533/1rjasT61b2FC0QKialbPaI1NGihXB
HUpS8ll+qwinR6nOrdNR5QgSVGRHusBTkz1QvmnZgCOP4A2ELHVwEoIvorcb
OCXxiGR+QXgpYWxRZy/Zs0QbXgDc4O07nKXT5FPsivEbLeJ1z5hkQNoyILZ+
uJG0i2497NyyjCTMg5HoLhy13Y/BhUuVPlZv6ff539VLGZRuTMsEpZomAFjX
ZqWuQo0bHdizizdMfOF9rLSmmi9ZkRDwH0N3MZG4w5KXSZGSsPOeYuTMmz8Y
j2zikPIEdQ2oMmJN7KJhJLqTxlUqjkTW/xcIhJKRfQn6xIOTQo2h01MwJovO
4mm+ZsTsRT64T/83Y8Asw63VReLQG9fGIc9u5+nqfRheBwcbSQxyKT5y6vDb
fJqhYPgrQTW0MVjYwemFw2wF0KDp+XZavEgmefKegLfMxg3V0Ufpa5L2otMj
AUUcSZNKQfwtE8Q0o+P7Jh43MEHu7sSVDyDRWs2pWHjLvmm+57FPSrHm05BM
mzZKsms745WLREsEa9CKlH1OJG54hvwwnakl4xoK1yfSs9WdCMGmmSfIhdFN
0Txak7SN9sQz2L8EIFZXeHEa4WPd6eHW5TGyfHPGBjjsms62fK6yS5AEplZZ
DQechAKnZS0UpQ2CIwBCldRaBQRmOAfvAztjy7RnJpLaQq1O0C/yna8zFyBQ
MK3iMf0pCZdcStqr+q7YUhD2OSbiQD0Eq8su/GqxAhQV34urKzJ1Sgez1vtd
nlWiNl1nSG3DcCgSOmUH75AyxqUbG4D8bCq6Cck8x2g49Y4vlSQGWAgLr1sb
K5BL+AGa7HtkjyCv7BtWuvSkrxivi8D5SymgGocahGCbSziwzhL02vv9bWzv
f9zHXPD/GUoRlK9w//oBQxGXIMC8NKSLfYWfIaQqEftmnHQ3kp46O/F9zdWL
B2KkC2CczaRRBn+e+oBXmzhbeFgvOVSnbE/xxyvMU1uJ4nlriLBEcwtOXPQm
GoCjMuY0R4W8mWW5HeC7WKqFjGK5516nhWewz5mZmVf59Eb4STGiP3/dlojp
KX7r9nVUE/Ndw4TUMKT1TFNgIC8u8iSPhryY/YmnjcSyqGGlSq4YeM3eUXR1
QbyJM8dUGShnkA81V2FW59JfpLwPQ/8cdJUV3PtSMtDzXiYUJUfdD3HcixmF
FRgjwYIwBUvEKlmUNRijs+m+XxzMoahAopdr7StSLIPTkZbjnI5Yfk0I8QN+
atWC3Pt8bRKY7CBKBjN280/hiiAo/M/BBYCD5mGbmfbjBjJb0rkEVuZ4pL1L
AscIgmnWFv1kWgnyzNkP/oIwQl5GDWlOkbSRv5NfYaa8pgmC1CBQq+xRyqNo
vBh1XqTUNXU0qQD3OncZnmelnHLLypB3uEnu8WgENCOAM9tiuAC5Yn0qeF2z
rBXV9xh0wAg/9NGpcJtN6raXGzC1C7PTYur8v1YeMqvZSSQ7Tt0U1QirioTd
UAdz34Hsn+WCMKSM7/PKLhih7wsLjQM3eiy27PWT73fwdlckthxcMjL1ufky
pHGaaMoha5PTLUUJ+R3JQ02QAxS7uUH9lrS7R9JoSIPFyrfwP1sxNZmbtYYk
+enHdow5VVsPYDl3B9Ad5WATTQGwrUHlJySTp0lV72L7Ui7crULjPkn2M8d6
HPmi07OMAn1sWBC5YvNneiNHuhW15a4mZsofkuSolBGIdhC1C1wPWPud/wu3
YcNfnqyfHWILxR+nnZCTAoHVC9u/Mzclbjav9TouTGFkd8Fh9uhMzZTt5bgL
Fqm3NSPpz2z+dKX8agldmeafNvJvh1jVPIKfuu3I8dvFAvSJ+Zo6/By/LKs9
ag6KfYVjdxiBUctiSJYi8PsnOKxnW8FVVdrDLZwpnjVyPU0QyU9cqLWQmtsQ
jTWfVS9rneP14KIMMhJ6cOu9nGnH7Xnl1pUurS0lRbd5GnfX1aqkOa642tj5
MJG7GnhX7OkHcIrDb7rfp/eMMlp3MqGV2dVJIbvUcxc87vQTrTrkqYDjYH6m
cvP3OuzhhCxZl1sTZJOHu7lCiiU1OELFpr0d9kxVmUuvkKk2F4iEwuKNfhl7
l0xxTtFxung/16QUd5EgmmsgGaif1pV7PjpDR4Mz6Kk7c9sejbREKSK9PsJe
EsV3m1A40Hi5eXNrsjaSkMiKC8Ks2v3BryMY2e1bp5M0I5wpqPys0k/QRJsB
5ZOwxRSp7TMS07TgrCzAwVqHdyOirtM0sJKDvxk+TpE+Jd/EhsQ+F4qokBIz
4N54Fr8Yrlg+s6m/6PtvlvdOTX42MRAmcHSSOfq8US3D65o5EITkUTiCEW/2
4ZSP1ukYVGoVL+oxnPG3EnJqil0ss7CRli2iQpVWcFvMiriicNGUstKvglgj
o5pUNW+VHViutTgU33gpaP3j6cEYMRcAt425IORZCj3ntBHgLn5G3t7imczr
DTQddU+ruA5LRl83a0mnpPewwHb1590PQeed32KO3EDovlRjZ1w20phKFMTf
DtFd0EkItawMj+Wc5I3RpucFZX/VSs0n55sEmO8RwkoV+pz9rowl/9I2UaMu
fM0wvDoiHvM5JzMdR2OfFZUJuTb65ROusziFu2wGIHZ5UojRE8ZH4g2Abrkf
d6b+V02gGGvG2ww/H/CH8tjouy5ZgXNrolGgooc8Y71518KkNWMBofiQMwnt
8yCzv2LJxG/LlW9KD5Ew0wBYKyEwhmMgbe+B74llh4oE6GxKJGSlpHP9alwh
afMQeEqB6HGVFKVOpXRe8P0nengQ847vrNhNXmY/+e7tIImNv7dJgZAnvlYO
Pqlfj2j67mfUqoIRi3iPY5ME+NsBOCoXpjfhaiJtKyefrvheVJkjF3HRNFCx
G1QrpEq51vFeGJyRjJuXO3YfDyTjr7FuTaXkTljcN6mMfF8jVyDo5GXIP1aF
Pc5dg6Mo/rbjeK5QJE72yovI/ya5tk37uWAkasezCOBBSBnbn4eCpRlrV0YX
XFzW0Khud9C65+9Nh/wcedfcvaHryTwz6K/Eh3M6nNX3odEwvfS6jwMYg4lq
jshoA0tgsn4VvTExPVfBCti4Pl3NZRNqhsimD12AKSpisTPQRHzvdDPl9Ij9
T+cC+Y4A1HffS7f9UsKIXsajoVOtmYFUaLJS+qc3WXE/LIluq3WjLDbxpGc0
ZzhVV/9au1bb0gzelp6PgmZxBDYsQxqSv9J3ym4isPCOFD+1UoUd9Ni4h1tU
MidajfHsuvUCkVXcAq3P0I1e8WVKxC8YbIy51TOFsl8LDJMd1EZRmZ1p+3Qx
VVLv2OAysBeXKDBqMVNCWMtL7xgD3SMFp5mF6CqIdywrwR+cUZwXEv1PQKgm
tRLuwsBnWU9ekmg8qSt+00toKoi/KFbGDd6fnXdRamDvQNiZxVkg3X77nkYo
H2L69UQkz5i9OExMg66W9HoxjI2jx/LGSJj/Hb/ztrgWlDg3AMcOLFBpiHZe
gvhEyA9bpSM/Y3xYnoM7TbOI38F2qQZwIwS5BZJASqMOdAbbF/+A/XdYOvC3
nOmRyDRZ8waM3gfg+Nl4PjQ4aoKbejNFmLY9ow3nGJLccgj/UydM2RIy0i4X
H0XhzdUm9qDf05dGS+02lScXRhHcjQiQobdh5VOfQ01v8ESohW8QODFSuzPP
r8C2bBDu1d5CEVgo7hEzHHXhR5hxuzvgBwkDOLnrQsTZemvS0Dz36BBb0/Ry
xq9shnrGQoBi4SeFpZ7rVqOR7SS5RncTXU/+8fR16RAkJ5styNfAKtZaKJRO
rZrZvovxdQxHB3Yvkc7gEiCecNoPCQYzovgrcJ2/nwmGZKs+uv6XUSj8odsI
aRt8oJKO3J8p/xYjbaX7nUyeCY5lOhCQ5RHs4PzfvEaorFOMi70GJ6M5WrO3
nyF537WRIJXnppT8skImjEOlkfwcgIw4WwtdKpiEx0D7YBn0vUNTVFLofBO3
tAX0EoWuNV2j+wOBAEcUYaTL075i90vNuqbxvoKKguJwU9c6ZY1lPieFKyY5
JNIexE643AXP6BNz7Tsi+l29LsQQgV0oWVsvPFB+rE9QsK0Y5TCAnYSqrWcp
sA0gO7oRQTN1aqtmEHqCNbdo866O9z8jMgbrjuy2tY7/ro13AaU1Sjzht4hA
hPPKzkq0a86cV8BmSaF1aK8TtK/n9IxPnGsocGmW0L+RjO+JRKDwnyVfZFdi
SvrNzcTqxZkVaKHax8JKzgOdmLI0/RHICH23qsaJL4s8JXd0Yj+EVWA37oNg
IlEWutvB+LWHc+/YwQhO5UQjUrIDrF8Dx+w/YcwUEFwwZ+Z7QvHYm05GyoN2
+jI+bc0RkMvHQqZ+t8qaksp9uH5XwB3wZTPmf8iLK+lYe9Sbm+j4PvU/bF5y
pVLgSN+5HpkJncC9laP1lsQkOJz43N6T38wQ8IO8sut8VOE3WWRipLkAqz6z
Uh0+uQLK3vE3BSKdgHTQNsuzQW8yPJIZLMZEyBcWihq8YYo6+Unw/RcKNK5e
4lRnUKZBANDZA9RbunwHv3QLigY+0G87BeQgqAo6sacRoEB6BGvsRmoIf9YA
X20QvMGFJNJwX44XEDW8olMP4JQmy2/sjmXrZLHiITcox1J+RkmtPAysAWoa
iwi/Q7bGbT0GxKiazYQ4iKRNYaEaqU4IFSKc2WIEG2DO8o+wBlFimf+Y6awI
9dIsBXWpp/3awDQ3ldtAJ7qBqA/pcQ7gs7UynFsn+5Pfj/wmlSi4cdYcINr6
tsb53GJSqxtt1MQ0LudWKCJQj/KBFNL1OKH4jAAvWoEfJGF1M6/NgVk5+vhV
KB+hSUH65p0Qlt0CwrArr6KhyHq0aGFgkHAh6CzPN5+gNo9MIs/ttszuMmjo
dteurAYwmpVBqWPoSm13eq2ltJ+WdXxiUlLnENqg6a1N8vCmHm4yXxpnZWie
+woUxWfaZvUC69rcW9Z8wwNNkp5KZGa46mJbdIf7rAssWURKXX8McZ/GTRo4
vbK2askObj0mvNUkDpmeh3Bj2g+cNkvoMVIg/Db+1P7Im3BqqksktSwDbpWr
YoF1sP5Mu0BgZAH3mkoujWv9WykcAjNKCPIbeVBeJMXFIYSG1XjUUYbsTd60
4woqR7ukr13tgmVtpVJuZk2v8Wkpjh3fy/nHpITirf6nWyWPcVpyEkAllxU8
seShnlFgvxy4sy09IK7JdvgeR0O8zypXiNu+ICVevAA1Xdj1ovxiKOUhYJOR
b4gjCaC9lsfqWByFj1HpRfG+3H/wQrCkTmm0DyyH/W/hcQ8tOXUquZDRD97K
lBgNL3yl9Pr8o7kep86Typt+XqYuYll5VjEoDHSXW2E31+idMI6cV0R4v3hC
pzeY7etmPInE8+3AcHs5ACSKLuM2/Z2Q+DSwBCFTxtq3EIqfshkr0I5nzdhu
sjYyZXde01UMfMuFsnpnsRlBVKgkuNegxcmorzDeYlZJVqaIenKxOhamrech
fuUf8Hr5kjEt9oAvFQA84/zzYu22dNX4ewzoCFO4WqFMJcNlMieeelXT1sVj
vFG4pAt7qD7Cp2WWgA07jvQwhPmawcoSJzf80YKwEX257VJIUT2C2nTn8Xbc
tUjT72fD1d7r4AXty2naS7T1p4/Axa72q38RcBWx9VBs7dVzOyhfl3BeVJ7D
qW3ZimooPqQ4kh39y+YA0vPqOerwlwFgXmhYpc2LguB8lEYJa3gJnSccWAoi
EglWwdSyZ5aS1XcRXJHJb3vubHrcPOOMid6ogUWreWhR1cBC4nGFgSMtA1s3
Fqv7ze3Kc4dNgMoGlultJifvilXv6juydCn52Xzs3wCvgktsv5enHln2Ta7C
uk2tcBfB//pnKtdnudB92DlPAtSqhMBHrGz5onmMZQbmJ6nzFMwnyKunvAMO
Qr7QqUECukqAQf2SRCtJuIH7AWuMcl+m3hlyPV1w2iZ09K5YWMNNrqbSWWvz
8VmypAFnMrUe3qgAYFZm2YHzq1aAshQBthrfXvwMI8b1C53/yAxR4GFiI1PF
gj8ywUYoMSiQe0jFdUE5o5DHIvHYzW4X6UNaF73GyTxLzlLImvzsIvV6hUNq
e/se0UjIdpFFzeIkMldn8FY6RD78BTXo9CjO5w1F1Q+BIKym0q3kKypSm2JW
dQEYMxjT1fFqif0/t2VNXnLayMjmmOmih+vnOLD0ey4STXlwZmqsZMdjTFqQ
AIL3dRv+sHxDYfnp5mWyB2WbZyAh0m2QACaVFd8La2arpuSLjrsFoCK/gFEa
qomMUKf6t2RqYPUy3YYOvZAifh/uvxmt6u1XoAeKCQUlhABTPJwFLvActyUq
xDGV20OKK1Nt+QKiGNU0G8JoJObtoQZXtJCtuk2SkmULHGg+1BjJhIK1B+Yz
2zC4wOYHlCH9NAzm16U4qCSR88o9dg7LJFz3ZK9K5k8X95FiY0e/mDu6zrf5
j7p45ll36Eqpx6tOJjD/VxU0QoqwzAlRMcmozenMMdWWP1nW+3bzCCQsFAuW
aGTCqqai8t1cCZ1+/+xM2dROymzM5W/Ys6mQrUgE87IGIdmzzmpZHrxdUJNc
bx+xdRUDMkpU6J7uDAVWlMHtbcfNv7waSXit6HFa3JTTBERtaMt05gx6sgzz
BjZ1JLfE9X4AtydOa0WsJxkS493kQ+Fma6q9peOgFRyPlJmFyhkyzA9DeVnV
AzqE78CIZDPlf1P0/OFXGkWNM+oLNgpOLaFFduY3FlT9T29OBpsQPwB0SqZu
QY+vfTWJN6/ez2vov74tdew4kiOKC7nwK0xKJyPyFi69wHSCPgNTMkWfEmAC
iu3kP5l5yYYokQmnxMDmKHzEAEPLpQZqlck1AjIZPZnsJ1kAoIk+hH7GTA1D
SJZrju7zI/kUf8030eDk/mtrO2A1ybFg1vdLA9MrPu97DJ6xTwEPygRyV6Z4
5ljtgUWFbHUgFjkWPsKPJvEWprsetb2VOMndH3C5JO4kl8hqOqoujx35RVRK
vXFROqjaNdTSVmptl4RBjP2pvvaJXwoILofA6v5La/a35sVzgLTwDOCQ/ULA
fsMjRyd81avuTcNUupLWnstgCiK3rWGMExlVTs38qXI4zvVAyYn00yVdPAXN
NJNVxW0MSgcp9qXzg4WVaalw2cwTq/DCGdNFPqOYrg3NCajnyeF5j1vspSJR
r09F13NhhELbhmHyYsHiWjNq/CMPF4GQNiwQYksV8aZfkob3Fpku3dH730xk
zMLl5P0n3oyooIadonI8hcyMr7CnrLKG9iTDsr2P5g6qUowAcYGgzGFS6rXU
CF2sm3Mtos7wYevgec5Va6wa3Q05+yhRd6mrvezxAVscMO//HhFS3yAdDRbG
Xky4mgL0xDPR+eMbiYUCOoYSJ9RQkH/+cj991D/ESp+TrAVvglC3yyQWFFTy
PAc8Azf8Ua5aLIrNJfad8o43Bz4ByhKEHNHWVhDY4rK8jyvYae+HtO74GBW8
lQ/Ku2MHtwe2LFRzekFFtOYOUCDNinvs+cV7OrHjghLXcVNCHRF1v7WV00GW
Ky14PIdhO2RUUk9hfAiB6jb7sA/ma/mNRefGN4OAlgFtu5PJ0vJWPBAM4LCs
diIplYvA+9cr+3nvtg4DnKMIUM9tzy2cFpu7+JbrsXKCnxFbNSt9JpfxGqy4
h6wbpCFVb+qX8X9nVUOSWGSxSDzj8ZahGsQnzcyaWIA8a3Xs7e7Ws2sNiPM2
Pd5jiRyAwahaXimxSnj0NVYdf5yxxEuPxvsGvgc3zCpnoxCfKdJRrAp4fHuy
+TM2oSm250F6ZqiChZh0yz51QlpXFloiY6Covsblc8ENHHhwOlAb1IfrlAmR
whDdYN56/3TH5LGXSe3DMNhITCAkApuB5fVb6lPqecVDNnMGfha4F3ORmlbW
jEos+VKJ+rkastYMzzizbVNh+ZdTPgT5WiGUdq6jUb0PgkeQW1+ur7leFcxK
i9BY6jzulK1v5UpiSeT+OcNDV0QWmJPM+d7+YgL8Gx+RviVEEh2Iog7byYoN
zmiZ4aaVsJ+NaL7PVu4Nx/q/Jj90AopRh1sFArc6xd57l6CcnT6ItOl9KLlg
1yiJpwIuYtvP2pySQaKn/PclKY0/2MboXe8ILvs8kdJ+NIkSf4gupyibNdeP
r1sojTQYy6YW3sFvHroVQcsp1DqdPB0E09hCuSvN9kVh3ZjJEw9Ym1hopApJ
1TGRJSHDV3Om9v4RdKXJvUR/0G1Tag2hY34sOnr3gP/IbzLY7fOvFRmhbgaQ
qKD1OgbqiOsNrqWix47JiVpJ/FlDHfZEwMYWPjzk77Cx7r2re59DhdBhnYG1
QSbIEfibeZQ/Z1xtTV+TGJI0GngLXWK20GUC9yfKh1PfrYqWiZJUNwR7julb
XKG15x4lMFyaiyLXKK49q6oNG6YRO/qBQGVHmUHBfXKeLQX0uMhCH2hAdxjR
tmnHeni3IQ5K6ys6cPw/gCNaU0xPCUzRd2Nu2U3f8/clCn5LjOVZadjdgAIu
nj+4RNInQ2CRp1KG6K1JBoqRhoifwfz7enbFrtRM7kDdDvqlX2Ji5LOtN6Hn
NvOqCG4kYZkT3YA8UCqtU+1/N8kRBXYYWTAn26w/i2NwVRx489rW5YilbMfW
7dNVxtudMuQjP7nbmoQr+GmTXbI5P63eZT1noOI9Sn/GHwiaWdGG011mLbny
4covz4PzqvpL8BQoK9EOVWuhx03J96qvl22zMKC8nI6rXrcDS1N53Mi+3/xw
vgGff7wcTB9yQatVdksiv6tTdyzzc83fFIUkpYjK1cO109Cb4vwHG8nz4ETE
J1uiUbO2Lu1sfielFM6CvCoqzyZbFgqjv+bnKxGQZWg3xbmRqzkYP3yHOVu5
J0KiKarua+6n430I6XGZnu2yYLt6SG91ziN8ii+IBdUlXRd4u7qJBNzIdUQv
NHHFcBM1NTYkKIVndLbcjS+xvf2dnkM9ZZEXQB9zRR7yiDV22V26hqUfZDsk
lW59Jn46/Lie3EoGyL0MgM3jF5OYS9aq59BgslxqadsdCZFLOwrXj8nA7ToQ
su+GatZdiRNiK3sEfH9e/IqkbPLJMZe3TuftW5lBBFC+8ty8Z/jLOB1tkQzw
y9KnN5gBJTVPE6+5aDGSOEbkJG2Iv43OOHrkEYNWsfvmKJRSapw2VhwpE8cY
rauiEuHihL6iL68pQofxa01IQgm/cgs0hefMugWwB2yXb37vRGG1pJo0GvSf
iEYy1LgNPEMMC/r7C3Ry9STFsOZFXz5JFzJGsCQ3MPatO43HQdG+82MfLVo2
sMwARK2h+lAdIGjZljDpYjT4ijlSdh6D1NjCYYCtdM1kZesur4EcNywjjDqi
XGSry5YWJrF7LQG+Ne3HQqcqd0XT5nbfHhG8FsGpSVJ7hDcxoy7a3C4qJhzE
6l/s3asIZ3saOBS9N8a2Pf0w+/8jRJC3Fw+oj7cUHAjnNMGKFYC7aHkJ1/Zh
IA4VcDHosIz9pkIE6V7lZ3as7hOOzGyCKZg1kCV1O4dcCLYpGqrVVyf+6P7x
725T318CFf1CJ+0bJMDKqn8ARZlguKArSbEKXGOZEW4BUru+tVZySUep6F9W
lkvODhtB8rEPT4n/MKjhRWrwlNNnhuwJcIHZ43/W17aR5tpJNPMvB5hWm+vG
ya9W44tLxKINL0y5VxVgFvlZq3qY9KXa7aTAd+58kB20nhNjWhFhm5z1QFqC
ggwX7qvcCT8pk6ZeefpIcAXa5f2bu2Ipqmf/vPCrcPue/aQ3leIn5PvREKY6
pM1AP3yQG/EhPdcVzF05xIPA6W9u7lH8DEToBwVVTJVfl4i/7/ZZMVgHrnaA
I3yeqO8UNdQ95f+s7ljguec8x1sIGx8vs8MfuR7yFazyISyY4iUPnvMjCyx9
T6oW1PVVZDWpuGSiPcEGxQ/oeqRyZFIMWb3wGT3C/inTuCVQjrv8q8RI12EQ
CoPJpofDXd67BFqWYBHoFYo629aDhugsCZ0TDNvlqYIRE+JKuuOyfOFNkqif
pt8jtZslDFm4J2Pj2WyvJX7wQ+cD+gEjbbtneDd/EK0Bnf2B0istRzd4lPyJ
GcLtKcLy1mBiMBVmvspikcl7Ju+PBSciiGcSJBhOglzg3/7uLnq853G0XR0i
b7cHOXDcSBgndgzcbee7UcBfnPfQEiSaTj4LnnM7ZGM9IFaMNS4EHowViNCj
K6UZYlC9np5SbV+dop6sp9D2p4qWTtCWHnR8Z04vSNOyxvB21jyVbFlGecc8
zZ748GKiM0lmfsJKejE8x9FDD2HeXtfm/qwQvfou0PbkKKBO7o3sQZ3QkHYi
pZl6pMyk6WVkjRrE239cOwgg5/7kD2AkY4kqMMwYfs7rOir16+xeTezNw5oE
yv4nH8XlhY7hJREKs93cnWu4bvz+0BtFj/dxIYkPWr2oDEk6QU9rPGT/ETIR
8q6DkDZF9ydT0LUXuku/vxYDhHAIhGVs6qcXpjD+5LRCGxqtxTZX5InIqYG4
LpNs8ZfkbP/WcitCnpuci956s6xp5gPMVW//O71MgqQJooPsGJW/ArQhPi9i
8wpSu2X3/6Y8TaizY1X8VI+BEbpbuUTevGiB5V5+NEMcCcd1ksXfsnR8O60p
OTCVYuGr0nEfNo05dAQeLhtHYz/k06xFZgaGgBESfP10mjfHa3vKGHOp9jR7
QBfH2m1dwDRvL/yBj616QhWemUETUzJeSRuNs9HkpVHYa870IdKf6VdXhT42
x5qL4K3VD57SAdPL9sDcAdol580pG9C5vt4P1c2y8vSXoLQ7+pOBBsfkWRAg
/Y/5D8lP38j0k4o/vIcSmzo/qsTx3zSwsbi0wGGh9RivO/Bht/zBDyprUvt2
pZ9Dtw5mHI9AReL5avedmFbKd9bQqIuNJ0EWZqNwzWkC3SHxp2Pw2J4dez/u
eK3UVcPHpcb6gO/9kxED3FQls/SjQ/UWO/hZAHLpMKXpFOW6qjzsVYJkVQQv
RCP9yenbcmUz5xUpFp1wy3R3WfQ+zUQ3H3pj6b4ZCXJ0inoX1J4ZuJeTquLV
B3B9OsV2RfFtrK24LYgtScdaeihL8KML1WIxOPAi1zQxO7BEIBjVUcKkSVPy
JjdM4Qu40rhWc6Dcw5fh5Ctgc0xgaOiSD7X7ZvurLJnq7kxN20NZA4hTzmDP
CUShQHCJfPTBmGVbvaMtm7l+BiXkUuP4sFCHtR5TOTHNOKd+BNH31cvyFHbV
F+Umms0Reb71S0/BShJpCD1mdYw0cn2CIP3IwT8tgTdz/Q1VVgZHrEkc13kt
lBuxdD/QgebYMFeEw4aluL3svmx85HidORiVbUmeHOz/sgBkNR8fgv2OlAgH
iadCsjhHUbfrJGPNqFF3zhIzNQ+VK/sP5Bi12E/QZeYz0RhEOXethHRSGTcd
QiT81NzRMyFLhIqJFQaczD0FBMDWIzWhDOiYO3xaFcdWKXvNDMoVebCfU+qF
UuRjoI3NY2m7982CrYpUHQbaomjYjiCVefWo03YSgBDjWLDKHx/c1XM6GAyQ
qeYitRTVXZ06NpHgYQM4dirAsiYHDTxe2CWqSRwWibGiB+6L9PFBat3TQavl
yojVv9jZJIoddPIWpNKwqu0jI9T9sKA+vKqMMb4dOyqiZul3IG26diiNzLeH
kFCqig/6RJD5CCMt4bB4JBjTPOYPz4VOvZsP6GERPmkdU3VQD6hglfrsi+Ye
nS2qA4cfmVqO7mWTfrsO0eU1KQ504FHAL8/zV0cokYrorXkicPw7CszipUCP
S6oLkJo7WmcBDaTXIjWWV2wO9zINUa+GGCefGkHpIT7ZmyqMDiCfJevLuNa+
7jK//1reD1tZ6gpEYz4irs6CbS5uwCG8vS9ChoYSgLhEst5MJBqN1BkPxkep
1K8dO5pwGN6NxYcwGIgTBsO36xBr2fB+YiliLE+mgR19wM/NT3v2pSmXK00/
VXJFrUgAh2RkT9vRfXRT8wWPv3BekWoYUjGledDuDChL1lYJgm70ZVEvGoig
Saj1wdlnwmJ/60X9mY3ZNop1E25cWMgG2T36OZSQ26z5bXftToaNRYRbmWmg
VQ446vk9gcyNSN3lv8pZekbu3W2dHrnTn4xzKJc7tppAoV9zH/kQNTv19FSI
Z/3bB2+M6/O5S6M6pwnjK8wZqfLwhinZ53kFqjeIsgq/CseiNuglyRb32AiT
+rRcVWsaijWlZmsYgfF9KZTFNjZfUtwg9B/k4pnlRgsv6BGG5wEhQmGyPlk7
asBSrGMNJFgqXiYu07P32UO/jmkIOA9uwGuBqe9mDXJ/iK76eDNHnMymup8y
GNRAL0wdGFwxF91mE47hPpE5sYLzQFs1uWuXA/mxfRwmaGqXxTczcgOiUdV5
wxLrHo69nDadN0oqG+0okZMnet3apSAFa+Zi0FEZkwOBBjTUaLjPNbajNPFW
fNajZXKGYuHT15osVEgVN/yZc4x1dtSTefnMdCn/Plfg42wbLeNiCiHdtAHp
B7C2gfn//11KeidVstXaIXYBC4LRSOzr0lTzlhk4Naaig6N8ICH7OKlPhJMN
hMu8jlG7ySXtzvcpEfVR4b49c8NaIGkkse/cSFAc8tohrZT5KPJ1ZKp09Vdo
JRQTqpEZdKAnfQ+GhS5RRl9h4o5thtwIy3qQ05LGuju0efshzb7qTcdTZ6Kb
QDiGoVIMMRyutyTZOcR/n/VUgTStmQ6cNnsSXuW/s4xSAZdfVwFn4G1mXojx
LFNICSrMUAyNWbptdkBEYBBswQD8XQsx2hzpMeV6Hg+MxVpXV2v0tpNCsiHC
o6vwuzmTKIBzDeScOrRf8EnjryAK++5CG+/K6bLvjioBAJPkSKDXfRDXXqCw
gMcgSMKUfGLJ5544SXY9280DYiTI2vl1SeClS/3YaTTv3FYEq7TyoH1d1rgH
r1khg5HqMR6lBpyhnGo8rNagXPxk9xbekBO8jKERfvsrqeSBC7k8vrknO7Ja
dU4F8j5xR6ramYENaX3RX2qLg+w+2B7PTQuipPEIbR3OIwdGg4IVcjW8QuaW
FrgQ3M/9TVGNxsGI+STMWCEcBNhbUF9g8Ed6nbYFLHfodxlsY6KTOxfVs7kY
R55cfx283+noHdFtuZmmTh026mYbVcJtRfJfow2madp0zOO/lHaLKOtRxfFq
KkiVEPRalNxNvcBalvTexPA/g7VuE9xyRiCd3fdAYPTo4W7OHf/SN4lV7zLg
c61M3GgsqPfqkPz4O2G15iCZ6JPtm1i0Y2yNJRxolRWI7BScgwGXODOwM0IB
86xW/o5GVPNSXigcqM22S4ZSzSvZc/3C0Vvkip2VEvXS+OQlp3lCQNcF+c3s
rYuuZp8Jd2IcAhrZgIT0yJIjlzg7ibZ0fQ1FOS9Ud4x+kikoNQ/sUGVRPaX0
cFYCS+K09QRl4WTOW//nuy2yHO4EcZ0DH8KYWpAT2oI03g7P0R3K0Q5OqrvF
mt/PDF0mpDlpy/o6Ez+8Gn8tnoUlSsNEyOoIaaNh4Or+BIXx3N7QoMNSqQy7
dI8z6N80KsZmaYf0nt+80fmKI/+kND0a2O611a+QbbQglBsZOUCct9SCf8kQ
og5j5gZCqgCus8T3N8g0ttuwbFqm89sRe8B39D13QlK2T5TmQsyFlUNFdO+W
STNSb2H4TAJ1uqr6DMcIfty+pEFc/dYfSmspOgfe3MW4WI9YjzxVs9TjQNxn
nTGOKbVs/L2CEsJ9W/gAUDkBxVd9hDCc8EscxcwQ313r/VjDwOOFhobshKOa
B+l4Fu2q3ruvGnyPUVrhAxGe/jt6S/6tGzS7Rna3m9wSglJtPCP4JO6wcT4q
UDuVB0JYni+A+zXcQAuvSRDiZEGwirRdhAImEK0TwkPQyBXJOfjZGqEbqjsA
YY6ZRny/+wnH61N2MCz1C2MVHBK4+ztJZnUrbsOr6tk7pObF0gXnnelO1LRS
66zzglG9qJiAWx0X5Uqw+8Y8z8o43R52AzR0+Q6QIPVF+BjjteJii2H7XPVV
2zCOwPoUrRA1cOA+7z8iTbpX60rm+vdfBq61YLRHHxlVMUYa0MiRjU7L69Lf
Jg2kVKoiZtEbEhC4T43M37SvVc4grMwMXsGUvFxmITknxuZVs/kdrnBQVHt6
7BCFl6CdHy03fOydD9hSWBf09Qk0p4lE8Y9KTUxG1QZs/sqLZwew7AgzGcJq
K1DjXURBx6URHVVEjJBczYK3N7x6RnTBPpsvf8kqdUiQkZ5TBR3dHLWrsUyN
xOpmSLDMuHoh8hmA69XZ7JTWxHPEEUDbFmunZ10lizmP/5Wqet7Mv5J1MILY
3XmL6RTFkLo14Ofxbg2Ls6aFGZlp7TKy4ZtQArOhnumXCY7o1i5T4/4GoV+6
I231+7r8Ha5xZdcrFWZ9IqGo555kiiQSlGsMihjkdRCQF/JV+5JBOVOXdc76
PQ5COCn4+Q+UemJw5YG54jC33zZqPKxuv1lNODg+n7+ZNdLuFT63Haqq7SmZ
KeLSMqHyDFPFGZXwmYsz7cpDAGC7Ct+Z5BxQ1b9EwKTpUE4ukCQ6cYnkkAh1
euB1l9RG4Gwf21r5OOg/s6dpnpxlp/bfZAq/R0XjTXldCS1Vm/pTWAa3tPCC
+Mnyd/TXdye2ljfYUXaX5NucVXncwXzn7oOx5Xi/DWmlev54ntcjhU5Puo/E
Z0TEjutgz/iwa+rAVBwt5j8NFttMbCTfY1J7KiZiYuOPH67hgoOl5cv/PN3G
mlxsJq+9frlIHpGUeWdsMrSkdl9oJfXyEio9FMoM4ECTPlx5TfjtbAp8dDVS
gNNO5hYGbaaBxwHTrLYnwqMhvUCiob8BKgjiO1DjRWNzmtofJV8DYHQa4Hhp
y4Nx6FSYKYWqPECXeM+8Lnb75346/1lTUw/RTBZU5g+OnicS4E24zJ5f7w7u
xg/88toIsV0HnnlXBTf6oycuXy+++weoznAtnBlpD7StCuzzWMjLVs1BN9UW
YoIpyFNe1SzVlwwr4TZ/Sw+SvM1SB1G5jKUwBCAbvD1p/JvVuIl1WzSevLii
EYOg9JBDTRLlniCDP1NWZ5wvHgN6H0HJYademHnJ/VcnIDm30RpdXad73AG2
bc8ii3npjgDJ39iwWQpt1hjr4yUv5YqIju+9exTfWk/la2ssjdrEvotizPwQ
LU3XUPwxpbE3g4Eg+1VD6F3yVLkBbblNFcxsApiDztruqNzuuYjyoSEgxVll
fEazB0khfIzTbot73ANT4KLMdSQ8hYhjfU4fK7MiCdRR+16fjZQvpnxah9mO
eFtkLeEZ8w6fNSVvtU9wgyygdAd425fkNbxBWJ/fjjVDHmP6NFEwEf967p7T
8PMxP9X5WfX2ZQXxVMecutTuW7ElTtQpkyMS58FuvDZOqu+fY1A2TAipRDQ2
d8pahtEtJD23NXct7cMOHVGDoVHjnpl3mqthar4WThksC1a2h9QB6naveBgG
zLhU4ntf0YE/zuKMR+R5lviwqLkRNjrH7ZbtIvKTMrIzWCrcRHUQUHqyTDZP
8CBl4J8d7BssEMN++zrvqGgr5FmnFpl5O/gtR84LmKJFtJp8Rkul0PNtcRdE
F++CuzB/dfjxTRFAD+zWuSm75qLCgeuXjkDrF2GeVHOxZbXUsqIoVU1EauYj
9WEqjfY57oSX5cgDNUUKc3m7IMKKChUpk7bgRbFN+AWekGJ3becjluZ5Tk96
3So4q7TFP/hiqB/unKr6z6X+riP+GE6TIsGxfucmfYr9Sdbmrb4Hm42Ak5Au
pONP9Z2fS/MEHQS61/rBWYuKtAH7T2bREXb7rLHugB/J6TI7y1C4hA/JHkab
cl2g7JE9CmhqjPRrS0kUfAcaKgJaDikHIXFCKR80tmeePFm47EpEh62zQJs+
Z5XzR+XzThnH7wuV3zQPemBnuFtJ/4XC3yL0eqy6XDMafx9LTcx3TcKLwYdI
jk5RkOcr3xEnyhDjhiiqgGsQArKjBAUvfB3NKjCwIshw4pY5h6Ee1gOfwBR9
m3fHE7q4S5s6ENDHqUFM5sAk27qLsMj+hurvqm5kRf8WufVAwqkV5s+rFc0w
kd0CpLiJewh7c8CjkfS/hQf4m3I2Ewqr7ipwCpxz3Ng0RyMBQoPMcjCwMXeT
6PigdrHnerY2PNpFKyQVux3i+mIqkb9HB5nyCDGGrmDnHTnlI8ooWOKno2/f
gqbyoDuMqM6/qbORxiwo/h3Ccym9eQEC915VbEiyXlQqI9hrTN/WWdzacbEx
gKavuR+F+LfyYYQfw55quAmcXoZsxTsYmNyL37k9hAofrIWFWcYwDuzJq4UN
Hj8Xg3qyP6wyA+uPDkBvp0F+272eb6wWU11C52/2ngr9mOISsVE6+RquFE3C
hBb0NYgs1FxMS19cs68wNSl4YRx78RwhrX3I7UKufpPoUGPRqw1p98UFNEhv
qvkojI9NbecniBgZD57SiSJYHeVbdF2OUIuksiWQFqku3oiiePEXNylEw7tv
L3dZBcBrWV6Cq1wX4XdAdPoej/kcrqbO5OQHAG7DcnvMlvYFJSogl/4nLN2W
hieLHjLXp7dVeOtIWwsMKRq5ktfmu2t7E4iz5touT8DYC7ZIwZSsfW+iJJE9
/B6C6aedUFZbZ47u4J4qonHJdd2xJomxogqhpVXxik75zLplOZthEkgjvDVj
WbawbdQ/NLbNd1n9bCtdc2mhJwPGGn98WOcJOLro9Ja2f00hCah3tEoImbs0
chBZMdb6/m2eokYL0wNQzC/AN7rqUmd+tH3dPhFxmDbhyDmH13K5wcATDQbO
MRHlepiPqDgP/iKG3YwQIOCfzMdLqCdyXjgH3pXgUAmAMKWxVtAtiD5wP44w
eheqMCeZRwDJv9y0CQwzZB5LNqHU6+SrrDy0VwCl6m+yXg3meOutNBhUJGkW
jP8DXqbHPjTQ55KaFE3W6ygwpbQq1w9bgq6lhTyDcgc0RY+o3b6qEKt4/+cg
QPZqqd3boMLvUuRqmmfvKaB09539DWyVAM4+nC4LJPJZb8CgAwRgtNMJgS19
fXi/T57piTx2VpaaslK7Bvj4T4yRBesse5ly44+ZMg7ZirXngqhOdahwuoqG
MalDJ4koc+s0U+YALO8ohqD/rmWDFnPwuAx8KiIDFTFCsFsM9Dp0/MkuhpGE
vXs05FyZkcB9TQdeUZ+TWNh0PD4MZui3/VMTvbO16WTA+v9811QQGuEE/SJL
tU6UTkJeRKch58qet9xvWopBs+2Y96Acv1U14LKtKBzBTo2xizMPlRctDrHc
FNJa+uD3/zHXb/WOnuomuW0fZH2uLvogcncyYD24i/E1Ig67ACvalh4ucT1D
i1iNE85Pj/NHO0mRsipI5zZwcQNJmg+ZPUGU7fqKz+09g4UZhdSfwqj7W2Yq
KCzeUqwhQ/yIX1aF9btk560k4SnekEOQ3NiTXLIVVvWa+2fqbWNeK1Em9+YS
1t5gf3af/J9qtWFghmNXxKs5gUtkLtbQwfsV1nwrroMfcpXFR0SI69nL+76L
TqE/WGLR6gzTWS+M8vn5dJ1iCP9Lf21WhZZu6Sj2RaGG0NewvPKGjjGEXIzt
NXx3IJtAyqTfrAfMX5QwCwMx6+HCzuDKeDFp/Ao/qV8zrSvT0b2sVfmcRZsk
19FwDYe8RtsiePuVYanCGxo1A/LZbKGiPlOnx7JmX8wjnI1sPLCPgSurKDVy
mxD0vInCV2FXoFKQzY3SEYhWkFImIQLMEbDFf8MRyYuzO8iHDi4Gh8BsJrtg
W/Ya/qaApEeokh0hSy0wbFRRwZCeIN2xID2sWFz/yQ+spa9F/p1cNI8mwdHG
9qKFU+DlDbPvfBVlTpy5+n46aUg6KtsFgFNSku8fKnOo/uLAxwg9nbm/bESW
h2n8obxvT9ctelGStJycSxnbVQx+aw0DszjM21/xNSeuNHy+BQuiKhUZpML1
9JJbyos9SAb1Yo6X+R5lLJQIoG+F4a8q1feUw/ENYHXvqRnYXywU7V0q6wUa
aUUcYVreIm9kf0C9KW/kFxU5z4a0geYilRUl7Tsab+nd0oSXturPj1+6JZXr
mbckwHqQmJrgnU5/Bb4rOaDnT1oZLQ86UxYZ+Fti5Wbl7IqVRtkpSPUwo4EU
Y1JldU2mh9F9UYPFRn1GvRZ96/GzNUPabL/SxYCl0VTZ9TePqocxrcnrpvmt
BM6WQYDO+02cs6vAPVuBUAS3mIN5HNMiVOR8q3uVMFhD1ITFym2Dy+1vQHU9
CpF2gIDK+JoRH69OHAvN0Ldwpw0kf48hnkaqSmD/Bh0g5iJyCumSlPhWaLTk
dJrkp/M05tiSVx+GxhtRnXUoZn3xuE2wQkTAU1We9RKWNf0Xyl72OxH3CDKU
73XnMTm5NPr/LadPb2GdhPttbna/pofy7q1KJDDPfTpA7L80AF4BuU7qSCPC
PsHiAyN6o2YWcXWiVpYNFOSb2/y4BBRdLIYNftuGnT2JA5nv5P1tBLT372oh
xQO9QoNAriP7RMKWGE1VsCjW40nFR0bzRqu64A6zhalRnu3ZVmAoJmGfRpXw
xiAIk+Icve9cupPyXdy6hDOu7te+4ZGtjbsJXNI/0UAgRZdYcXny+GPS9g6h
IXKbeaQmsGnsyCOrcR52hY7UkyWgHtt/+xyylnT9/g2oASzJBKzeg2dddso0
koAhGxRc7EQhTQPijdXV8NnPGA6+rWvCs/78zVDJOu/385d5z8oXNJYLUJyC
kP6l2luM9LCrUl8T+rEY5WV8d/LJ7k+XbseVYVaaDn9fm38sZnGDPAjmBKsJ
lgwKt6klPbjPVT/viImVtemSAc41zgiACsg4O0zzK+L17mihY0hYHEZc/m+6
2F5qsfVwxtB5eIqcwpnINyYfZR7LNIP8yD8WjQwq3YfZAskn5Bp0CE0Vfxxl
Bq+kUMk/27EneYf65z1JQ0xCMhHc9AftPwfLo4mdHz6+oDoxEj6O9CDkQ1Ox
j6oXwx4yCwmlXNlSppppkAa4Dq/BHK5VM9UIfa/YYzEjBn5Qvw1K6DQd2WKX
ucauwsXziCev44GNWOZ030TgV+ngj+ikfrB7xWlBrr06ktGpcatXeKw0CIQD
16Vr2oHhpUb2dEnThw6GYE3pkUStS7+CHyD3X3wWRYAR6TGwgYngI+rD0WVU
vdTCBVJUjnsIOcJ0jGiD9AkJ3UX31ScCpqclUlg7fB++j+Ra4wCtogNWNXhd
c6EdlbQ9j2ZDwUw534H70rfVZhYr1o4bUN1iv/48W5hm3rCem2+APmGzywGV
7kB+tOw3ECFU9+gpeM2bgB/eZ8Pguv6l/ZaCy31yBrTt4tdeenueeN9q2Wqc
LpMwZOIXOYRky6pCbf+Jq6IxioG2oxZv1AfdN4NVwKMsv+DZ5cyde1QjcOmv
5XAeLThU77r4D8Ispqu25CnZgL+B5qEg/5D/H3Q0ZlC/fO41LUNzaw6I2wpO
XF7vIxZtaQm3Wdpwa7FYCFEuSMKyvclj5BBSavLEgaUXB/QaJxQj8SVcbVyk
7xn+Y4W3ofYdeZVGGMsg0q3shw24pKF9hCQ04kJgykKz14GcAXcGIDWZBB4T
wYvuk2WYwjiZivaQntIFwWx2Dbx1M6JML1tUzWsbWw+kF/qx4SnLCV9zg4UX
H63eJlsOf8YZOsXmJz1U1fWI/pwcPjk9pISgelR6b6jXn85G80Zbp9KKEY9a
VdKIlvqLs51OCPAXCmVR1H87UucTKqwHp3jBbi33zaxDPjpjdlt+z6N2Ign/
S5UAHZ68/Z0WWdle/Hd8A4GYUhRFvs9xVJaq7jP364JTF7VOD8rA1ccwxHqb
D0Vq4VXl9DMnQH1Tut6JDWhHxUce7w3cG6hexaV2qnMGPv1IGABRpxdlFmdQ
TvupgBZblxd7Jxx5IGadT2zeq5AeOmW3GfLabsIqtJdrDJGl4sHXj/rUFeyf
eMj7LpKN29UyMkBqr5iD86B92Ejo6plOy6gNr9sYnUHlTppGZsRR2Wr2jIMb
V0qwIDF6UCV1r2zbM0Fd8tJ4qORN9HbybXcTd4qskaHzWLz+s1Wpm0RYh9TJ
wsZjd2g8SYfQ6iQ0Vm3POaEr29rSL7IdolkrpQARFD6putle6S3gylMA/ozX
/Zaig3PknCQ907QgqkP7pLVRrHgPjIejXPgpx3hGL4rFUHtOfsysl1VRX+7Z
E7ZlkNArAERwqNNJf3jimLTMLPDStEHzr7XPz4K3hxSy/3b3iNazAEngJZSf
WnaJ36HrdqoEZv+SZajqrKmjnHuV4BZEnxiOLX3u14wXJwieklketjLc/UFG
h9NC78Huq9yeGozL4wJQxQspeZFIj59kiRF8yX0/7QnRQ/oVM8lEaWmD4L7a
/6k15XT/wepqNYM8MLH2Ke0QabN6n4aVXTnc53MZCCPRgpXVQRudbzhs+/Nw
ywOE73ZRkLwy5yE+5qlrSA0JSSkJN1m0Vm7aJ87btifDme2q2LylVoD1oTov
5Fw9y4IuY8HhF4e0PlSHQO+kf8XuNC6EsBrm0v2Ebly8gEbd5m0Z4rcktc2B
ori2UfAaI/0S4Ev0JEiH1a8voHkKIEEB6jD8E6sh4qwDEjbCu5De8RzHcqQi
/qqzYTuEfwAeGKbqN5ZF7ro4TqXK2NcR4GfHLn6ecnDOo2lcPkEyPnscJPXg
6WKAs5Nd8M7eSZPRu99UmC+bvs3SEbH3Vgzickw+Uk2N6wA85Okuok5z6PRy
R8UljCzTzpmSNRIafRytwM4rGv3QhZfIYV0hDHChy6fc5N5AiC1TsyEVxJo8
PWj3s2WqUkJ7G3aAO7JlCI7juuJWcdIsILw6G05P4nMc7pslzezVPFQWPWYx
LNEdu1w43IA2NZpUS7w49cWk9YoxT3JYywdGC7Pxf9fyGmfcUwvVYWZCK2Ao
RdvEwWqblz0vXs8JXw+wPTLMonlGM8588Ac0nBg2CbQjS94vQKnHzNt9fOaM
B1amFbTl4ys6gall38VV3HmuVzbb7kBobX+ijOVJF0LhSgRdtq2kO2hd9kto
+hL9vIWIKj8Bd0WMhsQDx5mdNnpP562bEJTCNk3zq/BdGINXSQ364UHEbTrL
p+Ra0pxZXh00FrqbDWNX9SL8U7yye6k8wL8rWTJDLVzQkN3K7HDFWjzfK3qG
cBGtY/YH5+wPjzPbjxHhj+52EnIBm9yGjyab5ad4hqQ7PLyAWX6CmnQS5Yra
ACEmYVwW+pivvkc1MLyffobc4j9LwS51p2V2GIsaFPuPqatWl1l6fPqoP8c8
rFYCvUUtwVzr/FTWTkBXUUyAC6CYxazF8ySfUBS+7Oob0tIRPyxmlfy1/6Tu
WWQub1Jm6KTZGGvEG6Djaot9dCSDjv8UfRx5ZEISzu/HKvKJeNbuln/eKo6T
VSYDzQtFWMBARj6mCg9zml1boK9n6PAKtdxte1B8+SxK35GpywXIIfYZjQf5
jhTan/hXnchr4GQNtk7Q+ZCx0TCf1RTsd/1Q8Uy/GSw+Yt+f8mZxaloJ3/9Z
IquHUDRXI3p4yip/a/Fjcf0ENVpeRul/It8ACpKqhT+J14fVQnXu3g5x2Q8u
BBPhhakOnOgRjHSQ+q97d0L1lJ0Bm1oslyG1GfKKvMvNFn8k4barOIgDICpl
x3hkoLCHZSLK5jYnco4GDapMrthrZj8gxJ9vcPNq4F7+vMrWajcH9DlLLDoS
dG+aeJMavkdTWEnFbnD1b+5Nm/n+kNjhHoV/5jYNMvUuXxdrJb3ACX+3WsHL
ZXaCQ5GH8J4GkqnEEzTuPLTEckAaVoI8gECOT9yt0F1c+BanR8K+sa8+FblO
vwRRRVsHEKJvFaT1/WSxhqbN5YTovnX/KqG2fav/IH/c0GWVjCszfqsyU4S9
w2AeSBxm5tZArfle0cMHRO90fsGfm9C7Mr1r46gMMxGrA4WpxE2Gj64m

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Z1kxvUZ6A6pwKaxOdYs07NFMnLFQMgt2NVR5MKR5RKdJ8c9hslnSwQz63pqgbJulNL2IsMQbF1Uj0IhqVuqvHik8GKPJT0wra1hxuKAB80yrxPtVbyBlDdvuZxuBjXIgzc5B2XcslaeodZFtBeyMeUYfEN78Sx7u3lzsX2A4IXzLnEWV5U6gYlyO2tGw+1I67OKRfL/w6Pxg+cNr2D1Y/t3pkMof+6e8VFnEeyhkMUR2h7Ab+Vr/ojPxCzfqsll0zdm38L879UvnZICV+aIH6fawd23ZteNNULLemeUnAhs5DfrpruG0KQqfTk/j1X8yZogb1jCdtYdsyz6PfT6/ud/LYm03wqpkYpYWz810+o9BX4N6bo+G31wdz6z82iIb3t1YDk2I8B7cExms1jj5bUOBTnCQYHZ8YkyIPwHo3JOXu6ivC8EPTS2u3uenUsQf91XvUslN45B5N8WnowPmv/wJfdQu2ISa2gk8OpDnULwV7colAMpzPDg6wu+LrBAcN6vv+6/IwTzM6b9u3alNyh9dVBLok5wRJQgu43ekzW+DTEhk12fnN7XrB9i1+1W8Twhx2/DrH/dfBNm4STatL11J3hKOh8Jf8gEqYxyqx1RdG1JJH3lBJTAaJ0+6wyQjAs4L/yyffFFoGQjv7lOkSlVACaKk4JinlOQDpNZHkCznCaLg3Eltz/bMTV/tU9CSEB6LhYj3p3c4kxattHGjF+5OvdEf18pSr3zEfeC2W7xh9IJYkAM9UzoWdsTP7Sfl5nLwdzSZhBGL9eH2KYE0B+cEtEa1lnnzXImPrAeBlafwIS+RxcipsvKQQyMX8L6cTnA73pc/C03Z3hSsUa14IpAwucKxhs0hV4nKHVfUSGiZb38ngv4O4yYmbxqSEIXNE6ljUXNbLGX2zau2d81OIA+cTxkQC4wkEdwl7wDAKDdZzHas3GQ4bFw82jgY0M7bhGERVPbQLf1eCRKo6jZ/Zhem7QY6C+4EUuSDLMzzPLPp45xmyva8VriBJguw4X/h"
`endif