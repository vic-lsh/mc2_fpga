// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Nz5CX6Ux5VewJ5lDS4d8NwKNdsrzEActUj1s4OluVJdGNrc/EPwtmLpbqLJb
RxxG9UF0hyq6iVnGFvWfFsc7rjVfyUqE5cK1gX44OS+okRhQJr8vt6auYDi3
iHDcebjpdXE9FdqR74FOH0hEnr3asY0bBeTghZ6USF+9nXl0VQ3XAVMLqDKh
rbt35dZY/Eo6jvLglLDAZow+0z5cndpxvpS6vgHztnqyI1FYMB7UY+ETPdwE
Qqq/CugIprDjsBlY4y24gQhiWHjPe2vt7OJ1rnZgKNFqwYO0HYn1RXLwrE2y
OZv596eCw5fRGFjClHnc356WP1WeQqgtJqwqWp75Kg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iAVzLWotbxorFwGTvUPtNb4Zqavj9KxF/sxvLigGjK5IZHvOov5VuMKqhPmx
405iASTw2AaKxDbiIIPszYTnpNLDf09L8EfXYPgc4YebYM3uJJEoluuEnCCT
HZ63cZo+K455BdSHKC8jgFI6cticGBbD6kUvZtR63iXnjuo9ywjd6yMSfvD6
A2IYk0B3QRlYy2sKeherr4CqI7cp8kSLWd6RnOVhl1guZf7ZoTsw5cttTztx
taBL0fnPTB0NUI0RCCnbtBScWFYDSoZuC4YsPTCcAymAQNghFwUCntbhxUcq
yRMPBGarE0xj5B/9xAEVmipkGVseNcvUt5B9FiEexA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lNkXsrO4dZJobe133Qu4D/uFPp+yfdYAEMRjb8N0YIqqwqSEr7Kt5p74Y7Pa
8PU4m7DWYbkRpd39W8BIadCx3wJIH/BJDlcmU4NXFtp8r4J1e6FJuTUpRSUk
Akc/WTXFUreShTLdmrM/iKviE4V5c3/IH/kLC2sbMg3a+pGJL6v5fGs/ZSFu
g8+0XkiooFEWhU+zg86YO+qUyJvKTNT2GYTOKHZpZGpT3cSmLpM+wDcfw+q9
J0Ft+XHJcnLJchhyL3grN8Cb/YmFrnTaCZj5sSGbQ0/+gZAFQZygFqCnfjA4
jbxZr8IfcfuFTKFxOJPgNONcm203M8DJaiGaEA/z1Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BNWtCXmrDJXa8nts2GyZf0m3G6DSlQ1bhPozDU/U+Brew8Ev70jm4YUA0y5g
dRW/VqX7oTj2VWl0vxaV6lNpwoxuJHestgsmNjDakFsLKNHNZxn54RrcnRh9
YUfIixFuoQY6uXZUOSB7KdjAIQ0VY1krzsBP+VlZVS0ZgbzsGkbx0S7OKrpP
sg497uLiNdsCqRqTjckpxZFbl9JnfreDLdafWsoqNz5GX2+25+YzeQcnp9vS
t9+iAMvTBBt6G1GwKMKrA++tmZaM5m0LUrPXmd6y/n4dccH8pp7wXgm8qfLt
1JwLDjxzv8+cK48rROqY0scKs84cIitwSvFUmf44bA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lcoslfBBu3DjQ40qrbzd3/1hDWHy3QNsZQC/U7DT4/udmnsMfgSPw0Bsldeq
zdYmSzNfY9oiHoX/PDyblAG6XDz5opb1lJ8XcSbB7EWBLroBq7C2b64N5QA2
IP07AWr4ih5+K3WZ3LjX5BmXxsWVxeHhLQLJWyu+Xvky5VpReKw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UM5y+dwSK5x2NGpaRxAkga1VPzkVSHousNB0QiizEcGZ0kD1alVVIkg0dWFI
biB/C8ZhUPqJFh5fvryqjNqmCKC0Ot5q/LJqfyM57GrVxdjQoCYYJ0ipzgKR
Dcdu4m1FYC0yP4ojrWpwq3/mRPEjCDZoPGcy4RjN/2ZLBYnqp77IDyo9NGW8
49HtxO0e5VrX3SFpONd++bl/OaCFOVR3xXblzmfaEDnSZSY8h1rsq5kBlASZ
1T8MeC9fQM/W1rICeVPrrxiScT4+MkxxH1RLEGl3U4F6aa+1ZFpFedK6PQLY
N6aNCk9A4Zq395r6fpa9FUuu3gYNUVyIy44CUSU0SQQlrJ6YzYTl8qilEQN8
2Pmf6SbPpFmYQCO1/cur/xlO3iAaELgE5ipiwc9quA6CjEq0+kjndUY6lJXo
0g7WU/jWusCb4mNv6CV2CRzl4pSQkpRggMgzseS7F08u9FUS5NxrI2a6sgL0
VoDy/mJOzn7oVFVK0DzSOObYYnV0OxLj


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ATeemWh0qvBUZ3bM9pz9/ZizymhG0/mxbePtnZGZCAHMcmBSRqynPa5W8nIa
EPx95MCvz69RDl7a73i6t/L/c4v1aKAzaVmQDXw/1B0Hb7yAoo4B8vuTzMPP
E77w/Igmvv1M3PmNoPpgmnGzwVd7FU3AbeXZ/V1b2GwAESRR4X4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mEzOH/gOei+VzcYOzvooKjnmis7lR4zENrrNXYjMMq1Fz88vW+dOISA3nGeE
vhRXiIhspSxayPwhjbKRoxasZqpwXaxfAIIGFpCl2C6v82nPkKz7fPxK/dYO
wAXtpWHF48RxBSNRpbrsjibiVniDxcIPojKT81zG2rSMVUJir1Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1008)
`pragma protect data_block
nazLuNH/Hpks+L67TRU8E0D3Np0ZIKmJzfkoOdsBEPNC0VI/3qyJxCRGZ/E7
lqpVkVVWDQJ/r3iV5PbUkqYSDh0/FNNySiF1VmB8CXVJHQfB4e1SEAJI4ArL
JYaLvYrSNEJ4t400yv+WKW/YMtv8/qDLM/Fzw6lw/MKCde3PE4IxAosrMyts
9amrQVyI6MJlxD3xQ6hnQK18rHiysomQOA0dRmuN8RHZ1flZePpFBgoOtU6O
5xxabAbc8x3LYODbaq+zd0chW904VFtluomhbN1FkFti7VCYN+agdK2XMFzl
mrn2ZWUzOvVNIBsCXBBELTqT4lmqNhWePqzMs7yyQ1xQ0TVM8zocHm2pXTZx
yXqG8X0Mf/6akZFu2FkL2UzAtN3LD+PwwXfS71gtjh3q8nBg6E66lZ4gsqQ1
SQsPOUl9Pf29KoyGCq2Uv4xgoPGrbZpmg9EBBGfB5AxPmnkGMlNOrx2UoYCO
PZVQo8js7gM0aQmGdojs6v7uARxUGBve2tCvv/DRLN51avoYbJ+5996S6xmR
ynd8DN8/CoaUMEh/9ZEMNJrDb0JRsoG13Um7C8G5ZnMe0KM8yqju6kYeML1x
aRHz2+JxtSfknODK7rwQm4cTcB7ROokNyek31eLPmkce6x9g0SubXkIt5v55
G0mcRW/Tg0u/iExl16r67afzLW64H+kLAI0/HFbx/Pe3jpyDBJx8lU+iyjFH
9GtITsIJN56dcaC0FSx8PCkNr6h/oG5C6UNySRua0cU9eGF8z5Rn4xK86MCz
bgeDeWu9lhsv/0hgmH/vDaZR/KogDLfqkSITYq3jR+eBeuQyAzueHlX9Scar
CO7N7uJP4FT9AfeGjaBw7TDHJ5g5Damka0cWVrv0KwW9iwBTUDih0Tc+3JCG
5S4RNRF2W7q91jDMifx/714nRy1gD4guZTqHcEGxsrBHNbwWkS2vr2U3GVRW
cnqJYrjq+vp+1UnnEg/P4dvNGW+ir67a5ROBNJwGsDpVKj8AzazDqraW1Ngc
ceWrBD71zj6tz29ql/hfrk717PhD4W+69uhGtBqFrXyMzxjZdq/JybdyUgc1
DWLu8XXqbAebF+Pf6hKblUzJf9uiefO66IETScDeRi08MX/kSpFwxXtATtls
b4cAcfs21AYBpW/QAVJ4AcxWgZKmyqGH9Q6kCJ+OqxhdVRJ7reOQbVppDcm9
GilLlFeGC1R3caioiX4lRAPD0K1vJB6sl6Xz8+hBwFZLbON01D9toGngLMpC
PcQSSbVHAMcktTwhci7eDGOaY/d65U+Dnim6ZB51LDULbsb8oJ0IKBdkH+28
oVkhV+KuSOT4tKfB7rmqZNdx

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoxXEEVS4sdK7ShRCQlGJTpdAD8znyWXs+ojwFg1m5oXepYnaXrcobKzMVDMcH0UJbozpaEiqNurMGz815esbuNTidQj+ucXZlKjPxLpp1h9X2hOjRYworxEheb9Dss1rY3492b0IXItgSKBkraxJwzzrvtJWqfkM6mcMuM/hpGtHi2FGUkmccgpw465y3ojj2ddt5Swa6F5A3PoeYD47Kf8VDWCrrI0757Gy5Zbuw4QGF8+kx53YRpgriY1luQzCTuJ20hpZDgC/G4i+aEc1ulBmYFbcHy0eumPX2d2oM74btbsa58+w2uZlqqyidC7F5jC2C1IStTzbzm8DWloOdN6K/lyRQ+TfSbV8v2gb0+fulGSq0J23FY0lmc+SaDRjaU+b2B2USjDmdTlP+gvroic4Lck4cANBHO4yyLs3t0jNyijZ1zJylYJy3a1zKX9qeLCvKGpmDZTsqm1ZB6oaTWcihwxbtk15AKeXqUqWUo6HhV3JCkrLaluYwN+mK/LZSN3py5zybl+Ab4pXmF62/o8Es1pCIqhhQDFgZi7z35U5Z+oww3nh499plLOMLQckn8z38k6Sw6soBq55PI7A8iwqlZhgqqhF1q/IWahc9Yr852nAEtn0HuWFoPweemI6ubM+qcVx1KjKjbNDX00D7xNPdbKq3x/K6oMl880iTg7DRXivfpvhYaXXr356G1w1E64kvbS1szdga8kJ3NFDPcfhsL2n8V/4hXy2vnsNc1Sw+S2MGupD7a++W3CDd/E51tDI/Kh+sAYKsf6V8rFdERF"
`endif