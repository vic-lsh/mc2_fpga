// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
T2VDO5bgtP/wlD6YM7ivOOIqorRDFtlKA5nZ2vWjHjGMwAIX2e85GcZfm1gX
u6cHeXXT4WUbYzp0pa3fU5ubuF36yHF0pRwCDEpE2VKzXuwyMlsY2Kw2ItqW
TXi214wb6IAf1HXWcwL+IW7LswkLEMOM9w4EzkMJ53tasH2AWAuIKBoCnEae
WgYzK2xhqFnKT6A1oeLixvoxuxoTw0hdsfCl30D92CXxw+KAASsDzd0DRYpn
lr/VveAa33w77xnL4GYGLmWql79Bc4LS2UI4MrUU2+MqKVr6zyxX6HAjlGXl
q6YQ9VCxUiqSnzw6QctS8IpK8n4dmZ2itdNc+RNGmA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZRwo++GaekwAu3gLDVAgUhOEBYy/QY15Ck0sP2PgLlTk1XgLPsuERJmhuoQM
Swg1McuL8is+2Qle9sCQe7aq0vHWebgqGbIk2aRJA8G6u7dw8N9WcgybUFkR
j+2yPLtXZoNbkISXtpjxYasrIZE8dYe+WYGv6jKOJVMLj0ihtTI9f5xCZ1K8
/Ga4Q4DbUDAIlLp1WQZPT3iZtJ77im+gnyppnPIm/JTTvlnzdpzOaR3DQGl8
TUEb0CXUOlbJ2L56R0Go81s/RStZmN/q7+KlRvYiTLbYXAxBShEz5iHt+ARc
qMppRN45ahdR1a8uhalVneOfp7M08d9SozMzqo/USA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PclK5GavuE/+sScVIGo3sxAzBLa/lEubeTOW4g8REaxyrfM6y0PVOnPDIl+/
m7sgecTChOVln3jt7m8cg9xw3i0pH0bDInaOELR66ezM7IA1b7+8GYREaEME
gzHhZZoNLmQrdKbw7y7fuXlzsaYH83FpxGQixD1W/GrL8LRXBmVGVKSx376P
ricvXYss7RPBzcaSaaYrzZ9Kz7mrPmr92ulKdvR7lOKbY8M6DklgwD8Lx56D
/ktcOALvFzDDGl8LsZ34WB8zyXNl8yeKVR99WQAAr5n5kG35Ou/4yPvoHVeb
1ZYrVqKi0miG7zsDdnVwOEo1W8AvqB4ouB354MWkqA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dpW6NcXLUO8NI2OWjlLhmT64hmfu77XJ6GIYNAfeFhQB0TgMTOYdPlEO9YAj
jIe6BTtMYXOIv9NFUVBF0aTHJMQPD/NAEbVdaexhZG4JFnGkg+mDtMJFVfl4
2251G5jQeSaMe10bPC1KLg+FdxOfUZBFs1jzL+mQldLfCq5tihXXXmV0rVM4
MbMerbAKIOgJ8bE+0Rasl02mje0158UBTYvtyk0PuQg4Siv59S2u5KACOOq+
HHaQpN440Fq/+CooGief6z+2QcGw0HxC65JXtbrz+Mq1Qwqi9N1LIu+e5xnb
nno4B56PvWCtaAHStH/dxGAd4yylp7GbimGvhR3fnA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cjac5GTernMGVGM+uxqQmAhfpAWqAJQ7+CgWjcalzpwxqcn5cLqeaxKMrHTQ
WHDYBSfzhT+twYTPl1tv51nvfAEeoiUc9fOdS0jouu5l6IcI1J0ijTL08ek4
G6t7PI5+BfV8pnbSjeMnbFjWPo7C5BjNSTmo6IbGSunryXc/z04=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
utbByVEHkk6amXRE1JwmfLW3gWDDIQHaPSjvl3q9Iu7J/7C+J2Kdy9cebip3
dmWAm+1hmtoJxCtPztf1sbZPJti4sl41x19wf6QwNhtfyBbBXTVflF+60od0
BzuO2O2thf3p/S1GST8SrxqS8FG8dldjp3gG3GPPJqBC2CNmiv9VtBCB+BPD
BtGWPH1DkLp9EdW1v3b72/W+ONN2DvX8qhDTS7Dye47DENbZEzXRngARMeuy
3bkZ4aAXwuJdwY9XxkUAzljNYfv6eB0DX2l8oMEgC4qbn1xrbt75hHodtH8f
xjvi5zL+0mTtBY3WhErFoujjIwanU2J0K2d27n5frxLmSmZ+EeW7/9HlXgx8
Ds984pkXW9V0CjxL/StRg8eXHQFwYfFAgrkpfIT3c5nc3G/ulO/9xFiBrC52
UybtSGJbgieHHVADFkwi3vdGf1TMEHz0+r5hFUFPzh6Ynn/+vvAPcM7zV+m9
R2LJN0PwTTySyZOfaV0RgQD6TgwdIuWf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dl5V3UJEEi1+tMWwytJbA15RnBmM4oNeypGSVl9hx+NU9Q8bbkSTz5ajoykl
IEckbjU+dY5F7FOMoIT9fDBFOltOK7CzqMok+sLXFYOewSXo5LatJHaAQad0
IWtWAnzvi4dsyYdoGPxTZgWm2JSYOQKxm19tcd8vhOQsrWs7LBY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TZ2ysolu4hEDuTtcc6vzAxNbY0+0FH9UZW7etS9Bh1H1FIEy68f5UOP/LvV+
dCEq+RTvG+PWvbvJ07bMbp2sX340OFrnaPJ+nVcqFwlOf7wRTM5I+ynfl9Zi
l42JRimbGuWTAze2wpx+iOUNy4CpueimYBmbmpTcmHnk8RkTN4Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 269872)
`pragma protect data_block
d2XmR58rndAjUvIGhZh3crLcMz/DNR7gjZxZ/qoGY5P4zZ/OpmFowWfhcHGA
L/2eLWoyDL8RAvFwNrogZVd/u35/VbpBDhqmxu2Mrld5DqWUslfWUYcIVOaN
NvF5GqNGIYGD0eGzhwxtwAMjym6LyVqG6CRB2I6GLH/Zy281FLHNWLLFzySi
nIF14UvSRMjkE+fUVTnVowh53cxIKymNenXZuru3UzJfs04ngWtJhpB+yN6e
6HrkvoV+cETBZEnvG213+rmwDqlMsw+ZDVIRa9pzBhUarr7noU8/8AnST+cJ
zTsiWY+cIpWtHbwvjX148yYc/kAVvn/jCMMNupN7BQDbbL0iSENpTpGeL5zX
ns8y5gHTx2XN5zbJNMO1kLBEKMFSiwAwtaedSxeTvtBlKXX3CyAWPBz1wifI
0g0wIgLpfqesijDaat9w2MQvpjs8zWS4Xr/+iwu4Fb7B/G1SmFapuZciTDHj
jO6mtvfsATnTt7LDzfH555oZsi+uQ+Pm2zEAp1UuBhexbrnDii8wm5DfUR/h
SDbernKJxBhTsFDMvz/KPTUjojudZJnPgPaZCuZsZqX7zjcDYZBI+MD9PFAk
hxF7HQTGkOZEwPm3VTSTGc+bTThR4udeck1d/EmM5NjdNnlX4ZSJl9GySFlv
CxgU4TxFmFUKRo8mNh9HwVCce9Czo19X0lHF9McWr4EqXvRBhEPdJIPFIE8X
cv5o68CkUR+J077+6WitwUCCxX6Hd6+6156nJ9MLOy1MJGgBW65oLAuR3XMW
xN8UboRdySviUVCr4yuGJTgqqqUoJcZuKZo/NKRpyvrDoKnDLmUHMcjArTJp
ekOad3OhjlMGCyuHajkKXpNk5k3QQ/ZwfjnP3DUUJVhwyjgIHJ1nJzlT207u
KCKcz9FeAZdZQGBW9nKr/5tHFgPEC2Qp3IjhoQxpdJtLi0VUCd03B/SMObh3
8ZjKs1MDjJF5VGi0Qcy4z05uPsq+eRrWPbU03byd6bauFe47JOauhMri9TRO
3YW/ukiDC5A20EhKLxWKibUIkxYhqhClowu63cFZqfSY1kDrqDj+AnfChV4+
FR59DE+dfja68TWTNdhGkIfoPNGXcs6z4PGCC0unEleczRu1zQrwBSMUSpZN
Nx4f9Cidqf7Qeb1xbI1VSavW65tWhGBLOhQryHvtljYGfwNEi/LEryVgSEF8
+QS/CnP8MAEwSLRZBu7bhiph45ADhVA19qMTDIquNvzU6Gow8QeNbL5owaUd
+2NfIzoW5V1RD9z4o3MYl+W/OIaNYvEk7DBbT3+fH5TtknUwfcCSCTxQVNXO
0DjFuiQMq5VTzGwQRcrkiTP8FPfc3J2eFPJeRdpMjjKSMYdrec8yM1/r5h1y
kv15UiS5+joDyc4UEXvMg7EMBzELcBUk50bI8TGm1mrazhzeqXChLvv9BlcM
OgQu80E5NdI5+VMwDqWdfpHag3lVvrCUAnOxeMJukFqbnPL+H4TFfHy3c2y2
kVutLrgApMWRMFrbazjrTfJRM/gZ6FxPdN27k5Wljf9xpQuVQEIFj1phSYvQ
kC5nwqCIA7Gpzur3bYEOnS7mQR4VyM9XkK2GEnil7+ZnekVAsWmTltBOTXiT
bknmTeYk9LKKZwdbZomvJ1iW+Ce01Bnqbp+kfn84a6p3DFg3nmO4cuCXiPWQ
ziVmaKppgOOt9MJL42OaxvcR4zj8EJ+Pr1oYR8P+eDBfh32DLrRUP1cvjiQc
f+r9g7ueUSP3739FMfQ3ZJge0CGHvcGcoU3ZmtY71YzvHEmZA6eU2MSku99S
w/Z8tM6e0GCGzvoR4UY+DzCsQOj7j3GyJHKwr511ebHkSo4icVKGyRawxDyD
gtRAbm1eq4JIVMr1I2K6IfA5jGbd1y0MD51b9gmgnArFirygOEN6MwtTI7DJ
mZMTSB6fP4FIsM9uwojcJ4PDwETiferXMBpdKUtxy9Uc3duO9syGPoHMpB3q
n4/RMezZToHaILmailMj2eEJQCzTaKLkAaYehsiIfYiGKDFr3c8sWYD845rg
HT8k7b9s/bVPM1BMuZjY5Qbxu9x/DxHNFVGxMv5zAeWZSSNUyGhJHR1r3Wa3
A1+fMgeVCDnOwpAyqh/TP7seu30kcIbw3zXNLzEFvApW9NuVNJzlfJYlbgCT
oIGa5yAHRXaaCH4i7dgJ4hwpa32R6mYH+kscq4t0qGJBagAwMK9keUQV7zm+
DnAL4V3GL+EZlke1uhuYCkE/ymH0QHwbyyis6uGGrDLdfvA01gfwyaqCOU9Y
QWe7dr47WIQugSCTAK21sx0wXQKI+hV8i+wPRjbjF2Z+Ebn33bF0pNvx4uza
m0HOT00TQDESCK7I4pvPSm6Ti8M70ywo5t9UjphCP8oYykl2qJm/VxdxXwAs
Z2jd1Vxo6LqkGILSWluaX3rnTWZINeYbugeW+Kmg4g0n02+a9VF3ooAknOs/
4xtfdFHHAXINn0KVXbauAcsGZTdTjKOpBz+6oO+aJgFoPP/IfzSxZyx4vfkz
vgMUiaJGDhxOhSWl642BRcTaqnkvE8DE+SYgLfpdoBPeAwQeWowoLandCcro
/MTypOSva9IxPOmN/z86CwXv9FA/H8WbY13NaXKF37ObkbWtF2ZxJ1U7cNyB
oocQiM9tGMFg8bxSdoVBPluOPpqj5fPsYNK3z4VVPmKg0gVS+q3o9HIu8uWs
3mvnl1GObo+WIaEVLOXv8/vUAOxDKaWKg82d92fYXuaBiU5V7RfZGgZX4lmN
vbfaUASAh8P7VX9u4ZTGyH8b3bSFX5Nel5twVvuIzNeNkt8HqmGWPt83cc2+
tM7QqVahNGozrwU/AYr8e7YitETH55gVmfm5Yje5Q15npmN7p75j8B0AIOko
WQbNpzYclSLGhJwfShm3/4KUW20v1tPqa3Rsmg7zKjoclMx+XiqBS5+hjPx5
fetk4FsjU2cuHpKBHeSr6qRyeUYg1JOaqI660fuEuvX3AArvbYVRFxxq0SCK
kos0nia+BaYS4GEJDsiRyKAygdQa+5C8utJfOVJ+LdUplmZInA/5ZrIB3aBg
SNP/nxV7QKY0vIsrOD+w9kPgTWeuTCHZNkNRtLRNu7VzHqLcZN/AKqygt9rR
cqiHf5gJt8YWLPBrrvQSE1vzt273ySsPnQoFnpXgjEbmESBIIdfivkAw+zQc
bv0htB5l1z6XbCj5Y/Gpkiif6hwdWWbJycXVs8sGuJCgYty1vXSSkHmBNV2X
PxpGefNsTxJ9ZXSZwxw3y9RDMYa13An9yMyA+GgWSCZFGq3UsBnoHEx5/yWB
IwJBwF6DAO//nEtWN8iHgzYUYP244HHwXAtoeZw37y19Oa3Cbm3KaKHohrcU
6+4qrsZJcN+U4t+YmxYjNbfs3PQd5Tte1+4s8Qp9JNA2WQuFu4aDrn5TE9zr
Ba8RutX9DisrC5BTfAn7p74I+svZsd8dKC7vkxNzZ6bDnUfkDmlLY2BzA6Kq
4bwIsvGvk6e3ZNUzRcJTuF+Qn1to4eXzQoKA4VwDSjA9czoqRZREof7nWWRu
PW3yvxhQjM3ECF8WJJIf3RXtHkfAHsdNBnZ3osBgqoTvU+6MMyRnhwsYxhx4
o3CfveaV5yBVSc+6DYOSJ0lBJv0cg7Y92prtXHLw/PfWNsngH2kYukHgCB8I
IEz+A6HCyhIVIWaVRrs4zjV7fbakM3oaDjbKd1FJOq+Tswe8I+3QF+fdwQnG
vhp03xzfAZRsOGv9Furn9MZggP9AXUWsdmphHUP1JSEYA8IpZo+MsGa1AeKb
Vb5mF/lFa6gcZFcVvQAQhwidvc9q2nPUfyeErg3oxdBm3qvoO5BYtZ1vsYdZ
6NJy9ckwsbMgGSfXrOhqLqMmAIdIXHpV7j7FSYBiZA7Z2czxITpFgTgd5z/e
OLSywSoL7GJXV4EqIGbNW0xkmaqvGbzj36/8xsUau6JD0xnNARBeYBaRcpjf
MZAXnCUylOq/tchdXDECs1GsRPihQxzhIsHuQ/1WEYwg7EYCyfC9y7HTO43y
7MVV//qhPOittyJ5TRQHJL4MVcyW7XuN39LYpHa+zsNprFuA+LeNk3YfM7og
zTlsLhgJ2oT3ax6cf+9HaDitdfr719bYd8x3UFmWuL+7xbPgcElgLA8jMZBy
67OknWF1varmIHyCD+S6doSMsp1HExMaii5p5vg/6cpycv0sWVH2AiBYO9Xo
EFMSQzf+an0PhLFcc5V620eIticrQv8V+HMIHPKqUoVb6InItDw42LmtTEs1
w7X+9XPcIAihU2vOmdrdSXUXR4+tKjt44GofJYAgdgMjHZUuJSOxPa9EXkPG
ULrC/UhCNjljEnnDbVdC1SGwqzPTx1tkfYzPYB+AQLkg4duw80WEebs9m8Op
s5WmJ7amSJkkpbAANhZrAHkipNSK8M2fW4oAUzbYpLynC9kviSHO+npv0xKK
4h4MV3rP6bNh9lhbFyjnD2AYy6iBsThBYDW8/Qx7ByVrZnDquQirNOxcpXer
nKhB/XXe84Juh5w88H4vmRlQdLPmgwF/9cizwx1nWW8ctWp0KSXrcqxKie1u
vZUHKPC82TWQVKsEMY+IHtgyuqjI4U/d0hIyMdubXbtOyHcrTcdqWnakQQ1W
QWezrSOt6shoyGGvGJrAPU80jP+X5luA8aWW3Y19K7iKGQ3dQFMmrIW4dmO2
YGTMMi38ya+yZy37G70jfjzWAkb73cpPiHipmwxDR9jExxzVj2mxiaQssIEn
gVI+zajT+0+4ZpJFB7XCD/y+4EmXDhGtoiWkYGXGgh6SdHjFMZe/TOb0ptmj
0PupsQSahMOO/A60iojtuq+J4hWIQYoXvb3j8MIApTxKjaViMdLBui8PoJLC
79KBWdUEM2JdEdmDw2L4CWpcOonYpuFu6EZAe0UH8cLC9tO9t2RlcAsNyTwL
No7sCDMlGvFNcWEALDT9UfK/ISZ3qrhZxdcvtfrsYDo9qinpkPnARXbAL792
1mVSmgFp5rt1N+z1OA8W0/tgEo4qOERCGBmwZqxjqH/40FaunC3E4nxZEPkp
30dBXilmSAqGzseRbiFJ1GA9p/JBaXw03mYVAgPllWSASVswyOvrdApp285i
raBOMh1NgEWvOHVASFqsSPf8i01M0B7AvPAi94QNJ2Rwebi5Go7Pb3XV4jgR
VVUmzCkjkhZ6HcLArokA+TE79/kj51WEDxSAZfWPbLZAxqiF8iKpvwdXHY7h
Sx3dM76AFO7j1Ch6H/RDisxMuOBbQnVsEJAWSt40pn2hTlVagnIuTh3qkRiU
mYBbDbym5+rTB26FnDDBUOmxtI6dhJUbx6wALwp3YBrY+nb03EUQHpMnSh5C
h1tem1CGNXUyNfKP84grlKyg2Dd0fhX2pyd693ug7lFLO4Uxk1G8OfF9QNbv
0Qj6Lnqe0t/HczTKlFj+fvNXD2JOar4GObuI9PIIIC23u7gW7uvEteCMRXCo
gZVB7BLhHKoPWAHAfSXlrKZcngS9Z2dhnkjBaGdYrn3wKg6dDcevF3BOwxij
kPp36QkaT9LjKhhLPqIz+ty9xqUZSkNBkbR5fItPWTeq/VODGrg1emqMYqQ0
LVwVk0XXNYsrKzMZXfwVvdB1NePdCW7F9QsRsDyK3cwNueGBR4obtO7yadd5
7sKfk7V5NNb+P1A+JDvanp5fdnkphwrTI6tvS5eumM9xgKVR8+XS90cdwk2Y
dF9arXV7Mx28rHg5kBfpJCncqzhyo8vhSOiS3ivTD/Sy7w4+LCAtN6S5n8Sb
svsFsASe1YNJjA8CbKc7As7r0/IObDV3QF+OIIz3GKs+cSYFGIyR5hafM1o0
nyfNaxySwY/kJROTNOvM3XfL/T6wDKI4/wDucHnzMA/WwwTkAvUHizB6LhUW
3AZcXIakO97wYfS8Qlm4IhJVK4lu29wv6lT4T9TnI6cZSxXHXsosh6+XcZ5U
S2exAf5a7u2AN+n3VjlDyuUwfRBDR+l/Qm9AUdfnMk524l77Rua2M7jTzg8m
YyMShuyKNM9zpwaIoOn/9Boy2PgTIM6N4rk6phMwYVKe9erdTzQS3B3KzXax
kImuOkMkHHb2B//2m0oDEGhKI6NFhpbCSKMaRP/bL/+M9RQXLUNfyP4yAbD9
M99dJnlC5kEsLiwhn1jJwx/tfi6ydwDiXNX0OX2fTrtg1Quc1a05EgnEweyU
0inQ/Ptp7cxZkEFEpSTCbEJwrSNOz9GzUPlaOKsid2XoLta75kjzNaXtMPU6
FCljLW8inZw2DwFHapuirrY9oGmkuCknsJKKq6GkgEaZ7bvPoF70+tMFZzrI
z2k4LgMqVXA0vv+el1+RDS2wXh19wR76hBd0rzc+YERO7yDLFK+ahOi0q7t1
NgwyCPqKr2mI0Ma4wGyvnc+T4za6gJ+iaycFkIjGJexwtlJVf+rgZ76P3W0T
dE5Lx2UWMBLcZXZxB4GVTRc179NlbAn3FY3xn++QQOQQKP7iKDdmeef8/cPN
khOLPW6TSpRXuNvI89pAJ+BmiSQLP/1dQT735Y6DVdwaOV6RTXGlSq5R9kaX
7etgWW4cMxpE4gyicSJBbnpFTCNoIDJItST8U6ykH6tRzE9ddopzdJ4e9ouC
qB4pA1NaRSq403TPhA8e542ezOg6My5MBWTaUnVlVTcbbC0cjD/UliSlkY8r
sbEYm9qFRUDlpSFi8rY+AjW1EUvPI5kSTxSLklo/p8nPdVJTnoj1uiF4Xuzf
uV9ViZB4p8iQKzA5UNiHTmQgW0daiqUHF0/BqpPksMqJkR45gZmnSNrwkm+3
OqbGdGWnOBioacaRaEKAogd4ohol8Fpv7Pls790amswqmo2uWvKs77Fdem3P
cCFqLTZOYLiT2T5VEunIOeQNZL3DihQXIQuGJmcL93/5K5pGWzDveVFz+UV5
khcJ7Wsr9RxfxnbPIXqdcaeONnMLz/HKopRU2xWiy6HA5OOaV8tGq2DU2vBJ
876wCfJVdor+VHCkoLtbaTahCv11USZmQwjQ9SwZ6ovK6003HyFuwCa2hC1z
7KLP6XmAup4kSFrsRz5minbM6PtwUd1gSwYXbirjQWIz+nal6rIyBvl94n7Q
e5EFeO/fQhu8IJ+Lpebl5BCfyB2GM/iK0mED3BKnpCQDMGNn/2MdcYmHst+j
slYJ+llUia9ccHkRR+RIFEElRBxJwnlul1B7JVYGgMcXgEjmvKIIuNGGTJDX
5NTvOD9uoNpl+Q8Q7Vw1ULCET3rD776NYNuggGJe4JfhTpifFQ5q3AhD5orc
78C6f3TMTJ4hVXxnjvp6o4bwMgR1SUqhAN+vRS+FR2E+8Qf9VYM9/oUH8Zy/
qln5rGPSCVWxjhprTNaagnVmHcUV2CIwaZPKmP5gCVzhfdWBqhupkwfqdJvp
4pT8Ns593CTR2ryYKnIjXlD2ZpZspVTO74kMcdZlNC8t0bULP2l04ZUXww3n
VU+7JzhWXabCOmeFIs7broY5FNiFOKcvbsqKuTU0s+LYMdy7ECnh/7VoBW2r
vmdvUIudSlZzjqoBvBKYVK/CBiPE5PoSQztF7Un4JdJZLMHfA3M2tfxmqfH+
XX3PIz5b626ntF9nL+KBH7EKA9EYVlqpSO782wozHhbtk6Edxwsqq7IYORqW
UgGgR9wqtARGVoWKdiuZY4nhOHe75T6hXRPNyItAom/rrsI+6IsZEXuVMKaI
PfNNjqnoHhF/haYgFA4tcChYQ7GAqpNIRMPGZlQd9lJnOR54KYO39XmJ/4Wu
8siNGT+oq8m9dbQT3IA1OT7q5gC3gx9wdjVbYrsfd3plZbEi1RkgujgLbf5d
qBsxoGGPoQoCsVZn+491A05esdCSQNy1V1d2oUIq+VG6DkLwzlx+R03twF8u
9NqQQxpd+ZnNKODvnHnlWrX5SV4yVFv91U88jKJ0qJCE5lKJeG/W0usyBWdQ
YxIbpqWx72uzKI6MUMFvdxlilYrRPzOA10YRj/gqRuK19PT424m8l0doXr82
Ad3SrTOcR/bRoEXG7fe0+f1hXDV9SEqUci/WT6FuwbhvJQ8wFRYozxOEJ2Xt
wb+U5DpB1ZZ34bVa4w2ImXY9XQhpAJkXiVxiSF+h8VSS1/sbtpKGj8cRflWz
/+yeXeQLldJfVRIr5Y19P1b478ajxHJedn1FM1vu0W3uEI/sZqacieLbSjRb
u5QQxNkTS8bv+pFP/R3EQb21Z9JL7n7r/sYUF/6L6NuyLvx17PZfy2oE3RuL
vXQq7sYD2Kx3hCX64KXnPAudR+5aoc0aTT1ysXt+iRyQ2MnDomuPnT1MbxN2
Md1WaRKp6kRubcEpORICdQegWX5wOu5qQJAsE4CiuDSBGhbLO3MHN94rCUtd
HBfzkWznqWb+mhcTqNOxVYMt0d+fXIQrTXGYPeUJ7vkC/27f5kzd0Y9EGb6t
TK+oRviokjqA2CHcC/pqXkPiOUcu4t0WuNSGbWaDAsF2PJyR6FEHZbmuRmSn
PGcleWTMMcOuTcT7/YPIwTOd3BPNKWQlfxR3Gw+tux9s1sEJZ2cXFtqfd3k9
krBvqWdJTNAmERb4TQM/+ZVYPK6mPI6lbfBqmdS55llr5VU1TfozFf9jQcM4
5/GfeGqyEQlDDDPEEVk4yji2hIMkXtdkQGHyONkG6uECYnoMtQvdy0mZ+SeY
EnKuIWL6BdpBAHpWJAjHGAYwGFa2iK+uDwX8SkFnHqmoOHbsdvs2E+Lg9e9f
5ZLwDqETjZOtuEgNbEq2YX2NTMB8OaDQMQrdyq9LluKDhtnbzOnG5Zo9/HUR
oeAehWFmgJCGDaVC+rX77Mo+tXnGsvOfVe/unk16ACpxQNJ0TyklJn/LUoQq
UkB+ke2MX/iUofVK0ZuooiNC8SsJ/LSP0U6D9twdZJp148oQ3asYHUSnDlt7
2rLsvx6MWqWzNIp46GLAG9E4r13xMnhkwOL/cDnctWQ9msSK8RpEmsbjdDrO
PIiZAApezrKB3qvZNT98YxewHLWR3KNIT+eZ5gV1q6hM6LSj1/xMxfAabZ/s
v+u+U5fS5DWDfsSCJh1u0VcVMZfHO6Sz89h3SEdWQsdLtswIwLCQOlAky057
aTO9TCLj4SuC6GsDvHQwilNwshedOYPrjie1dAmGDIamob+D2f+6CAWsTtCf
NqAJE99jAtZ/UoZ3+9jgYpw8lJKCCoBCWOLeX5n/yHhjUjjXRt2iEz4SWJeN
55i1EJrY/JQRBAWeN42F8BcLG+I2NF6xdr6ovTnkB6T/eDrJLN6SKM2wgPke
tKhHpjOXR0Pm4nBwFuovFJUA1xRFUhVqjXLaNvXA7mtj2bdfX/YAdfI1Bitn
6Gpw+PuqP2lPi6LYz0+clWC2qm/xBC+m50ntrQNDzpNCvZzLMLI5W5goIxJk
2/AC9hn4vm4nmp2ZRSTBkc1MvfpdPOpZQYnDmS8k71VwfUY7fZ9PnYJyrYyR
g+D12Anwqn5QuLWC3CKGHqOJz4JtXoqvhDNF/vyW3FKpW1Zs6QMZyR6MHYJw
5c1aEAKusF2ZX1T80sipg8bDrVdXi3I686mwKLTV+PqGzBnimqFLeXYyb44Z
8iRd46ZcEgue40F71U1yJ91TTWAdtOuqb/xLTrSLpMZFT0AYrySf9AktkIH4
L4VaHGHI5ZVzqMtsV8uRB9dmVS7M+A5l+MJjJYIFdtdk/XN6oRmzxrR4tgxN
twRtXaqWM8sDXS65czvsVcTyF9yWkh54MKBr3UTIVMUpAE0TxLJfJs670mj9
zhLv470Z1RzUgXd7mpVgn3QXOYuPLNyAlvG9HDOlglKhNi2PugPwY+ff2/tw
sKl61MJh6fuhTYyoZHdyHs/cMLhllYZIN4Aa8qEd0dmDN61UqKklZx+1y3R/
Qo6vNJh6OZlCpsC0vs5wDaMivIHEE4LAHwqgtJeZ75CWvCCnorh4mkMIMbi+
QW3oj5lLhgB4N/wLa4pHWaEvqY4fKIrpp9k9uhkgS9MnQQZeIpVzfwSBMuIY
l5hz9X9UKxz5/yT6oAEgtInaXyBI9HS25iBlx1EcN+10JIBk7OnRxOAL/nLU
OSJJftxIlf4VR6d8hFqc6gknNrlajCVBAgwdiU35ac3++JS+QU1Uk4Q5AyCq
c3rl4Lxk8u5A1oEJiRr8gdGAXTG5inyyKbtBviXKf+jRf596fi2gPcFbP6Sk
A7xK+/xLbwxIySLT0/oPkq5f/vSP/eTuSm6DsTpXW7zs7+zMKWdLsO3FTQPX
RntFBjiKi/zKwbI/Y6Bx0pdYrHjKESvgj/l+/hdMe7APWreLH+nVPJzSedCh
bViqDzNYCqDr4KeborgPm75PA0oa6qWzUKjRoAmX+RvQ9BSCvDxx/RdungrZ
jBiahA7cXHDSfI+4Im2LcQVZtGB0N0FxC1LNA0weVqz0/Qty5mnXF83q2ENl
HiHZDU62uopri3kRNul2E3qPMMYoJTq+E6yi5qqIPDVL02Zvrdzh8LGX67xi
a48XX6Go16yUfy+0u7OcsqosUEqwoAfIGPa79BXczSOXvjEVUpE+KNh5ADlK
CQcQg6RQfdAcdlfgUX9deV3BTT+MUlosepqlVqFPKUDbA8UP42+Xu8lPcJls
WcuQVc7JgxfwVK8oKr5O49A7cLpqCj7A4A1J5IVNbvYlT9UGHtrn4Wm7rEAh
IFNxLYrSKrInAOMaThojJkhFrPYXFsW4JWi+mOK7r9WXQVlV9nBMMnJ+AFl+
62ng6Ts7jidiz/VsTmwM7kU7UXGpqlBDeaOQwGYPLTpbicF+RmYNWQMzEK4G
HtBJ/F5pWWGKqCtPthQ787Kqlf6QhARclnhHL0a76NMX6XHFdxtT9ZKlSlNY
3tKvXl4bL5VO4gl7Ry2qTvxn76SjOjw3S8dih6cvp4xvpoglUVJCO3ESbvYy
pOwO4SSOvchSPYR98mcTgW+hu9OkqzQuY9qnGgEwoRnD7Lj9uLKfOeu5ss/Z
BrbhffNti7coubcWxqxzGOojv6hx6/YougFivsHVI5o5a3gfiqLiKGTLJJIx
pXHdIOLLp2uRvP/x9ZyomKo9XS1VKCLyRy+oAB2QNI+l2+E+PK3jcB7QGp21
dim2+ZUslydbc5NusLVmGU1g31TE3cTD2yve2GdESEL1cDSEn41h1rx95jX5
6yGSixi+j8VV4VEpdKIdWhduxKf0udszMeu9L+08ecUcQKf1UgAm7fS3jKUu
vfq/WfLV3Tpe38E4riMv68GsOzlyfU59jvAvuorLx9/B8emDcF98BHSaMQ4P
MyF0G2MvCui+Zm5hBvxabhZ4eKTWRehwt/96TxhanpPKlkplm4CO2dmH1+Ue
im8wo8oBmwJzokZanHOzK0fXp7TzKrkm+vpGVknaHbu6BD7tynDy0tcHqgbW
3iWCjmbMe3HTEonpur45dqvdCg2tvxd1A10UBSbQQCWLMjBAQaVBKksyQvWO
2RkmSrxycsw5Vj70hiL50nPbLQBQ5UGUCP8qaecoMAHBv6GzSYrOeCfUTCeU
Y8RIuJzmelsakmTzXqpTsnIazZ2yE6buTCbJsskxmVYtmGP5SAIzLwak2vm7
AwxqCeJmm3zIFF6BAEwhAlTaxB79/QmYlYjmTK9zKqVrk5TtDMKXM718RBx4
6VYvOcF2DIP4V1pHHvi2VNAS+sEl4IiHXmTFf6NiV+3pMZMgeG05qssp0zyA
i7BLRPi9k/DF+1oSZYZUpBOPH5TTksRjIhQumBCs4FCLadVPG/wu645wIIz9
N9FwlYqYhWFPHCm4QAFLXcTmSPpOw4f6lVUGjvwwGKj4aSyHxyv8/qq1rtwv
tkUvzoKJ6mHdI2S0o2hWCUxQjVVW3sx5VGBOq6OaayoVagnN1rAWAPxCDfZe
NOlgYgeNR1GvrlRPa3aAN5kkyrHEJDCsuV1PU7/4/iPtJIDOm43r/Nt6cxKr
CtEhk+PVLWepoE4f3xa8jqHesOogwhbq9nrlwFIeAkRgMtMxErLhzcJsP+dR
TtpKB6+oyTYs7IsiDOSSLWbw3d2nRhCeCBKvOc0pmt8b8aWbilvpZGMcLpHq
5SDGE/ab9k7zYx4q7foJuXI5uj29NFQ9fif/MWbInem136xhk1XlRVX/t9sx
HA1RWCHAyL29ML6QhoiRmtlCudF7l22V+fyiXiFoqNvgfr0MPkio00w/1kU2
vvcR5eHEeMYWqzNFfv54k9MjbVK9rELSWifd9uiKwljPXpcF44y0m++Gz6I0
4Es8dNjtDJ1BkacXGI1KG7WSl0q5gYs6G69R1LPJ7vMUnBvFaHbDOE8qqLtr
cnB2u2C+I7LCWd0HeGmi95DEH7ZkXHybpmTi1E3fF3AnjvU2flJ3ra3YlBwo
we+ETQNTYD1Cb+KIFDvr4BE5xFlyqZ+qYcLPARkdbgFT2OUSgClzBxlu/I9N
xfRjzSelwzgdEPaRqAuegipD4TOTogCkfpKWT+V8bxympeP9Yf1lgqDfXBFA
6i3ksNVA5rq0Kb3ORp69jAaOD09kVKUr1rIn+NllmG0szx2YDRGh+MLcyIe0
xAJyhaHbBIiQF1jUS4XUswGZR/UgVimHvrKfIbrzODw6EsZKBDvkHsAFNiL1
Y9BdpnFqN9TyE/Kh4CWNpC6/7OHz/CCw7XT583rVCcDxwS2xNMzCyC5P8NIb
QA5j2Y8ifnfzv9fYACnvKpYhdfwFSNr9ys+e9KGAnQAn5uJDgGv10Ddxs2B0
JqSvlMdEnapUP398jLqvV7Uof1PIJWNIxY8vu/d4uKTrGOeo/pUeyFyZku00
FSdRKHqS2uPtYElilMq4o8hoXpfrJuRM/cdNqBER3TllYHgPswczbeBqNGOJ
DFy0Zt8EnGDoTpf+WMHtwqBwz76AZJnNofFHisQyRiLV2dVdLGBc1OVdgld5
jF/tvzUjkAnF2eQDOhO8MijOO5kvP95f4hmQoM8ntkcvRRuGtPHqCjFT6X0b
04mPR4Z+5RUbNTrXJZGrot1AKZZGN1LAbgTR+/S81hVCRJtSl5ATABUTGjwT
xKVYPk4lKISIiHl+NrY+Arxg+8IaC0aMlQCpT5bCyTjUCN0ltPgSL6S8a4ed
hWW24eNWsSiw9ZLLVN1+RgEw012dlPzrqf/eZ4ugYNuUIQVrMpElPI333wxs
/g64Flsk11ovJ3kG20mIdAKgvfFidtBSEKQupsJvMJ1xhAKFvV+UeYbLuiiB
jC44j9Mf8Rb/sc4xgz5Mz630ExpB9VtKexs/UUFpNrDzxKv3M1f8MwSwKkYp
q55fHAS24ebc8DIrAIOXft4MchCD3zB2IaA7n6qpwAnQIoAPlT0Kblsj84OK
rg/x2GTBg+iUW3dfkRlPmJ8JzNInT0lkFtM6GIkpM18AfJ3uUIxihT3tUyK+
ElgDuTk1aQ/di4hfqmBqpFGIfyAlpZIHAIu7I2wkA/fkhAMwgZcuhOo94HY3
SQEW4GvkFNFtgn6DLhP9mDhpfvUFTeffGKPJADdf+sL5bAnNbVVo5pbUB1n9
47EBdsVeRDTBLKzGevwGBQXX1HrLWeGz0jBV7EUj34Ywj8DszY0JrcN/TePQ
wXcIyE3LdcJ/keM8em9DsIDf7rD6BRfJTyRSDdtETex+ieUnXEtAoY3hF7Df
L7v7deV5YZba+0NpV2PTf9bP3v417c/sK3FBMTTniRfVtmTf7J7VV8Fs7DCW
Ivw2YX1jUMwRLOTYimT/pwXgSLTWFRd1AVM+NGsVGQ9o94VUqGPaYjDtz7yT
FjAl7GzGQxGL0BZxNcsI8ikG8zoIQ+mWcYtKHf2E0Lmh0Se6qqYrYl91Tg7I
7TJ7JkgBvdmlLL604M+26LFqfxM+R6cch4GZVUZ4iHxls297RoVEWwLGZx/l
NyfLVU8DVEBrQDfUIjaF354HjJc1YQ9R94FaspDiKcfl60LSztTzYqwCNUtL
Q9q2H13fg2zIVTIjEaKlP54ncgJzxcL0JHEkx6Y9jlEWoOFq450rZlUrsAli
fRe3hOq3i0gyTJ6JvqGagwL1rvv0FEJG6CwGoToWqwbq8b9OtYCOnZAkp4ms
XdO6+yXz/ePxg4U20bXrRqHky/ps3JoXkdQQRifouN8JiKgjxgmTjP/9gNcP
8mS3hwfACSybpS5fPZ0iw42p48h56a3A3nd1Z/EvKC+8UjzF00bA2k7uJHe+
NHkSPqOHaNspnPGgU98uwzqAiifborJZDPpGQNH1G09JeYZ9eZ6g9A8Rq1Tz
1SjucZvcyNPc88b7sU3BWMdusOF5iEXD9OaS4dJ6S53iBe/U8yME/MDPLwoc
hlPp0uNapS3tUz+dOISeWKvjTaRwbIovrBe6/icsylnWSrCagLuIbueoXS+8
oFExPEPVO20MZAWdryBRmFUnN5jS9LuSi6yDGS0B7/Sxp28Ww7Sii/55IyLz
E5IXVWGafTrhwxy6WxLzqethfpa/GB58jlgUEJf5kXKzUQkdEGR9GmfkfgUX
/0J0+W8PRA+yrRBxB0eRCKbrU1q3AcnemJWjsc2tZIQdmAxXejQY3GgrewKL
8+EoMr4/9YXU1eZdNarEpS+ZonS8/dBBOLPFn1FdUmsi6giAM2bFPecy+sSJ
O/6ZLokQel+Bda6hcjamZUic5NYXmwdrrNA4CuajO8G9lsU3FHL55ilwbxA2
jhUY8o137X5DYRch0CO9CV3gSVbdIJ4d5oSbJtWCxKmFPQtkHY0b7EZTpT/I
LQq/t7/SwVVdC+KZgSpAEWsMDrVOx10Od2c8ly5N8SVuak+NkKU9dKx5W5oD
Ew863m//5MN0JaGEGrNhdihvyLOw/5Gy6KF29e6A4m4no4Xy427J4bAAmeCF
9sl0z4TuKxVWUqyfRHpewLINw8Itk4/LS/xG1BlqtXplp3JWlW+3EfUejNSZ
/xzwnNYPMQLvKW4g3QBF6d3DbGOwgycy+R7GCE61vFBq2OXgjy5oSAy9T93C
V4vnImnQ0xMiYXDTIaSxvCQxhNGeQAsT86fc8oeLFEgmP74PGLySNIxrLcxv
akO+h3Un+rotcqQLNUFGRMpJOK5U/rw2XwnjLLoSs1hOXolf8pif47a5IE00
l8wc+FOJ7/wuNboLke4QRY+gI2dPYC09XuiD9BvWZzo5YDairVPMkIpeZnAi
jDBLRHg0Ki0ulvDzqEYVTThvKGY/DMukb4phX1+KthWQ/ussZzKcPOkyZDua
CDUiizcoEquu1J6mmgApDR6lkGuLEnaOPjYLuFwND9Y6/bH7KEE7gzxZHpeK
G1p21r8blZDPbMY4BDXt/1nc1R+vfRITK4qMvzXzWFq+mMKPk92U+pCkdUei
mnpVWEgSA192025CdaU91T1rYUTWgVxP2K1rP54UR+8Csfw/3rqKV36QpAVD
MewWANHDyz3JeUYdMgxWmeJUDk21wikDNS3Xr/EkJVfs2xJXGQVZ4Q0kA06d
WmGXh/k+ZIsLSmCaz1/ulmNPiz3GkydcoHtC48aCpvHm6yctWP+JnsGSEvfS
T1MLoJ6pssywRaI7SxUnNbK20sYnrP4WQNQ7kG/D5QjgkTKm5w22fEBkvohJ
WQDmS7xpyecBAMd42EmhEWxodZfPOmaiwBbx8Bas3b/PaLFeU/xxIgCcDeS8
Lm+b8HqUdqVq8dlY4/VtHnVHMlV6FCwrsDDY7wrcuGD86w2twz0/vX5ROx25
sQeiIVd2IiLjubUuSG5+FXiVkVUqy/7N8DAokL5O9qs571p1S7LTLz4rDDQi
0Oy2dnPqJ0h+klUM9J2wKOSzK5bhuf6BKjKt5WwDsUWFIkRxsXjdsQOwUYlp
tetbNfWIjoayETGNy5evjoWqPVRu5RHT8MHvm0EVbpowlYlIbeqNvhtqnHef
dOg7+y3o2PaBaSXZR0bWaeKYLY4oHp0RPhoLLf39vpoM6QZ7J++ohbEMwKFQ
fVzCC7v9qVyLeTkSXg4mCor5rkgcfoLRW9jZciSD70DYpXNFqVrZarV2vpD3
E0t1/XvlsaD2yS46OLzZCl5wnFhRUA5252cWpHrTtuRnASVaRqFPl3EEWYZN
VJk1CNaOHqXlGEVWINWHTVf8LvNK39J5B/AFX86uKJbm3ZyzSSsFJ/XSR1li
5VAmLAysa+5DsrTt15GM1XyQPq0MQ2SVwxHJiEPgshE/gkCdXcJWyh5h+QKm
Digdb2hahwZL725d9Qu+iRg8eoXXa4FJjgE26IZlUsaxBgn3S7n4CyLyxhOF
CD0R2sfW+reWYDCmvZ0BiQwpjUXXkGtJu08ZPaCUKk6CwO8eb6aeEWbA9Ydk
dWyILzfQ1llWMJ1Ju2guVvsR8N7vr1YADxaM1oAVidqe5FeD5dlF2NzFL4Fk
qEcpZssaFMnf+MeS9MqzOccX0PW3gUVVCK8twFpCUSNt+SgFRkZDflPDC6UJ
oCN8tIwHtcasVBKBf+P7gTLjTTx56WriSMl8KuWp/FxAmnDDJlXIo8xbMNmr
KTK6fz4XEgXbDnIwsb0Gde7pkFV48JdsYraUoSR7EZxrIkks9J+8J5ODCZZB
SMvvJfNF5yPczhgnsq5jU75JTGwOsYjjUHW9n0yBVYPe/gjziEpTBh6La3Oa
U2s3ObqRbUafieI2rn9gmv+WWVK7h8GRdq+dCraztqSOW7tTQiTSC7S84SnD
jh7cNJ6UIc8BWggi9gBYLNcixNCwcF5v133iaqy+/lEZeGF4lc+L6gmNNXNC
0W5DU46/hoop12/0GVop3c4f8IJ/A27EevJPynBBWK5Ys24+4L+a56jpW678
YgqPVhV38waNGsomkg4Tm+52rCAr3W8MpqTMfAXm7P9W0Jt2D6NqMtjlMR8r
ZjnbaEy9AnFjhKOHV+3nHqfNBrusTIszNCI3QRUxZEaKu87xDC2toQGBKjzI
MG9pWrfVKRC9XR+raN8nB9RwqePdG5KSrUkYGduSAojwq7BxGSzN2wPjfpVO
HDyK0M2MQsuzXYf28yAHhZ5z6vpACB/BEVprqStJ3XWQeNZYsxSWbBp0/Mo9
f9rz2afxTHv84JIcnibG4JtILE0GLAps/cLWFms7KlBZwpcJbbO15vlfMpwo
14MKzLL2ORaW/tsDSBvLLMChopgzw21TIVJP2HC3MMi2e5rUymCMPMMNWee1
2v7cKgwulaD+6rM5HaqP44mnCArZoPcW5oukJqTx8UmNuz5wsDFLQnxVdjex
Gq/bDgqRQfJzsCfhTV8bUrQNlakH98oJuCZZdoaIh5BYXpN+HKqJZPhrlVyS
azAwzO9lI2skkxRJNwQ3OhIiZItq6ehzJaHD8vls+UftPFFnhjwcakaKF8B8
NKzjfyJXyAZt1a5AkH6p+fggW3ASZJFU76tPmM6w5SImHEqeNyJ4rC3m3Tqa
m92iUWoRcy0t0xcNLYmiMqr3OD+71nHKCBKT1T31n1aBTcxLK1fSZUZg+wcc
Gyw0BoqGa/VHQiAzPEpwFEK6/TQp3lC2g0V1OQzUcJ1atptItJR9fqMJm01K
lmRiJ4uh3iRzk/LuAq6YpwtM+RjNMfwAyuGmYzI33RNGZqBXgj+OY9mggu5Z
hPAChLYgSmjea0mlcZOqI8NTlajPveS5yFD43YUrEoVR7Jjrobo0Tmqs5mgo
mldGkk/2Z36XmflgxRZ8uc2UkD/wW1iQ64x4sOGjJsnTgp6IAvjjeh1R5G4n
Y3d/glv0vkBkHzSzAPNEFXWaNWEURCmHRP8cQA0TrJC189mGrpr0oxzgevHT
6C6DtehjGnV1g+NC7DYdY7qFT3TcKR8D6QXAht5fOd/B0DWpJaxwJWroHipt
vYvbokl+o6AKzseb2ISIaGxccIj8xx7vq2t9EPcgf+zUrnL0hO06d1TJicqO
dvuOzmhSUtWezFNIvxoF47odddLZ3nWl9Iwn2URCf1zkeMz7uOm8MTxmlg8t
gbV37RcOg/OVD/lquphLpu8sEu0WaPdK2TTxUm+6L/UM8163AUyXxuMqIaol
xizV7bGeKAfMdNtDDLRXnS6o8TdbL/E31pOfd+WkBY8CTL2dTwKo+OYuHEh6
r7DFhxzPF/35Vp+ZhYPW99u3rlTq51R/LgnO5DldmDrXei639MACp364ANW7
92ajyBsOKPE9eoBuEGGjoczip1DiiiQHVCyFvrOCFq8V2mYwoRB2jm8T5NpI
LQ1qV+w4ouka+1YdPQLYqyIDoSStxckvvFrj+lDAWlGeyXyfMM2qErEWAj/m
bomFyHNadsu6dqaNAc25jqrIa1Bj//mJ0M8usDalhtwr54QBICAnXMHdw7wT
92GN5EDHZ31r8sb0f+jTY6FrSVSjw0eMcyt2olUHlyJBGIkhsjDVrJ24twXA
LNkFWWNfVrCr55h4oFgNUaMbgNCLHy8NtBvp2KVDBqBtORKKRGFw+sklUQkx
/2YA/4fYkbM+0wOli4zkq9kI7/2kNJFAzrIR496jrFTTaQx9QYmwk9K+6qYM
yOjBgZXuKG9GgYSj0tDJ7y5gzclUWv0rRi98lFiF7+eZV6yv4yI8EPMGeHH4
PTeG93Uzmb+ZR+qOISzLK9QJXnttxZwpJfrz90mOj5JZMApmVYfAFvjPA5BY
d7RLhkm6/lcZPMZKYXC/rr1k2aeDjriGiGLtgzW/agT/V/Lf97xXbqcctVLa
F52841CDx27mIKZKSDvpdPavGpADVEQDVhwuHSQ3u2KRE+Teg8Jc2QOEeKGc
ESO46g3mmKvxMumZUEJiGoLNd/0jkxdk5RRzNEUuUI57HE4UdEgr3mpX4Wr6
9TpnKSFsX0FDanSluFdmpcoXqGN0zx3e6VyWW+SZ5UTNCV40z7sh9C91bqt3
srqXZkz5JAq3H4iVGvrSbCHSD+pCTKRIuH2Wc21cfNH66IRXHCYG2T+qw9+A
lD6EE6jk/LvIQkdL3Rq+ra1Ypu5Swn9It7ANKj8WwqcU6pdnRaoFgigeVXS6
A31SAJikzn+TrRCBiW7vxQPpwewiewbYXFVyKUdJ6V4j267wlv9RUYKJSS/7
Vg1IvgjF+iJYWhH8JaWluPpN5+XIg9qt3LuZo/AN29sknnn6QQ/xWnQdMhwq
ZzIgKMCXFgmq1Jp2mc/9FVSK567eilP3L9ju3ALv0GZgU9Ll832nd4K2+pjM
s27H6OhlFm/GyDgB/8lx8BkNBGoxH7YzYKHWXPLYrL8Q8QEny93J7qPmI5dN
Jz/sxxe0eWMzL5SsisEDkf4DUSrAnEa1VU3vR8vJzPfTs9uN5KUmt0HgY9IU
dT1cNWdMkR24NGu1zKR5QKBiQGF3OEtQ+hE27YeLZy91LrVe+yjiS79MqENk
/l2Yd/VE4chV1MB1ioO6qgx5fCGT04JAbINgOVLJfetkfD7okFiZJX9esQns
WW3ifJFo/a/yNsL+8C41aHJgEm8n+XMHkdZvfxtVQCuORW0+8tnVBJDRGZrN
pvxeu88UddOn9S6OqRRLRBlbiWJVfPtoiE0Wo4a/O3wdtAHswYzfGWvD3Q/s
IikOaFRQerWdiHM2ueLwsU0XI9Ws1atu3cBacJ8mmUI3XZBfmy2akAzWBSER
bGUkUheb/1wmNPUHDVXwKVrS5DnVLBC6Sq5WEDaNIT1OJruRvgFNDqQcBYkO
ttp4/J9JFIT5u0pfvEyNI/YSV8++/tXeNu6v9Nmx1VcZC70YKH7+4SJeAzIt
9QefNE8s5fN2mQlGV8fvCS6h/RxDVizWtIS6fIFQfSTf17sTatdCiYQEJJ1o
zKIEMV4pikf9/mewlBDE3FIA3elcruiwEEDCunNXgwZq0OT/9QaEJsxEQNHd
2aQXmBU9/NeFuMpokXD5GKoQeEKvz2f5+FpQ6vy4Caxt11K2tJ0gpwRXjP56
MKwq7pdEw6NBkHEoSVSZgamCqZOW9ks+e7RDxzLKIhmNS0O97owFNldUL81R
axfxQSm98JMej1ODRsimqIok0y1ix4RhG2g2cUCHtmbAFGyBxVRGn9FGoSdG
4J5aPCn6Bo8/509TNxIZzdVYmrndqTVaHtELlNSQ6IH9pbXnXZBxBlLN0mRh
dXnchFrpz3wdubE6kYM3ll++fopdgk61sZ+c5edXjy3w97z0QQ5WClv27DIE
QRnUdlwoVIva7yks83CMCvxhysUKc6JMzrGNcTA7Vvs8iBegYy7LNqyj4aqz
DNQFU/SPTETVDbzBjN7MjqBcswqZ0ecysWyU/7TfJu0vwUpzcMfeO0ceAquP
Q5TBxGG5WIMnP91/K/jPvZ63n/pyeSV5PYBhjvNrUDUOx3dkb84u2w5RYwW8
9R+z3GnBZnE9EVktFlAoCh99GknWNz5qLexfgrozi7XIrjUo4zF9VEInky11
tzH488TKuFcGNhAqxNNuV3e2AeCKDzxk3e3SM0gYBbbjxiVn+UrXL/JQkOxT
+n9f1P/4QJIq93FCB7Ohotexs0ruH+b4dIN156F76fbqcxVwnR9Lc11P2Rft
HOuLDWDz6VscSbXgBOCVxEPxUStLfr7WcEog2GQKRpAb9RFemuCPTnskbDeR
Uhvl6w8loxbj/EqqzCj4hbDXbVqxKKWpy7it8DhTWriCmlgYlXMdPY11KeU1
RH9xrTF/nqup1GP1+xOJyxtG4X9WtJv1advjkuVPNRg0D2ASZEFiv9laBKBP
STyWgx3iL/1Qvt+OygGTaV3bjBQfw9w06+AdAj7FTRsXyMNATD3SQin/otJV
/EwsSd0TRO45FkhrvTCDkUgYrRcHYdJ4LOhh0m98t2Ekp8y5BRTMjmbbhFE3
GbFpBAkEsjRs6Avb9khHFHw0gKrZBieuRnRCCiiQ24RH+vI8zs8OREV6yjIJ
1WxLoqs/sTqabxekNlmDMMBw9saWST3qMfbRlGTVEBQBPSBo6VurGJED+2Cg
80s6eA9qOJiqf/zbWtGuEu9w59wiko1TUKV0eMlKnQjJvn8JgYdV3/3vNhws
bWNrq/E8UHHQQ8urbwUrT1wvmTC8bVz5rbcAp5o2DAhKBOA9IxGAT5EaW4p9
oDmGfOzvpKWY7A4LPe6JszmeXg8jX5h0IyOJuXHf1k07PkNJ78DNJ4J/ukLt
fBkkMfltexMY/TEND9n9+29d3eCeO017ToUw+ocKvvuyUngD6Pi4TsPvOX4j
Yay+R8fPl6b2vHGO3+3BTr2ECbHdj1Rje82xR6otNShCBp+IqGk5zH51yHh4
npdjburc/RfttOAiKVjp1uM2GAkHksYyIwMCsuWs74D1TeuuEPoW37NxzR5X
ZO44ViZfvGkohpg/xvgdEtaiWNTT+H2KcmNCzDv/jg7sL88a1d61LoIimBCX
/PvJvh2kzLpHBEoz4NLRxudiJx84FxlMBzMgXmc/QRll8iRNdw0hqwNccH11
G556sXR+gsw5l4/OWYAKcFqDq5KFgWXguv4NLguOK4mxwj+5+qQfaT+7WRMB
FBpVZ/8dCYAIVJ1Zfg8TjG5jzUYot6r01aPNdQffPPNr7pyQ1FSlYuUzi8/q
KlYQacdmUQzF7S7mGUJ8bjidzRS8+z5c4Cgt7Euu9TVH1kb5x9YNSgB36vdZ
PHHOff2dDaJlEHkw1IRKta5YE0A1RntqS0hNPGxLMFD0MlWRRinLioVURY36
nhv0UhrlY8Y3KuCrGI2M/ciE4FLhGJziteFIBnMnSi58WqIXtm8cEskOe1B6
ZawbNYLJLeJKp4suEG5T1D6BLzl6iLZRkABYDNkx/nXFDl4rIX9fOsysid7D
YLB9hx6kB9OLCXqjOAxVtlpShz5hjUCZk7pAFZvwXy8Aw3ind3jXNu5azJ8k
g7fw/K2iAQso2LJdHshmGJxnV08bwCaMCnKc8HBZV++aQ9VUSvFJd4XYLsMo
EtNe5MrbRPbL6BrI7jbkK7yirj0S3gBgVOOA6iNJiOkgYgXlZbe0bAmBmmb2
NC6nre3jNUSQ4Y/Qz33pjsuDtFrGul6+xsQCHZlrzi/DcvHAhbaugzctWS6e
dlbXW951NfI9MGB1kF8Rp40DhrqQ4rE5heSXpIYhw+l7NRgUjOG8wJ2uVUHc
MKTKbzU7ucAerSqfycp5+4CRS5gvEzwEg1JeT4Umyy9jUmoqoQOKxgaEO9i+
T3Z9CHKFiwOfcdZMz4azxCglXhz/BqyNsonIyKt5yuC4wjUAtv8tonPThsli
MPO1BcjSnKmstyonkexJ7w1bBFYDB25zcGHTzvb3KKEtvon3dk74ITXZre9T
2EjJV6O39SBIWOnFM9KYJ1JE6+stBKBW9LvIMjsxRS29Vxu5nVCWVkSNIaik
U5s1rUU91TqpLnNoqj3ImprKTBKjh+JWOFBszt+Jr7Z6vm2iYQgivMXjK8Jw
G8E5YWPJiPMf2pBjTsvTcwFSoFNTNFL9wTnO/Mh8hvqgHwJfFsZHjV2UOWSC
btRgJrJ0e9BOTB+Qd2iESkhh2KmbOKUVTaKhJNQ3eICZIG3OHKfNoAK2znJB
wbvo5Z50q2UXnS59jAyiUsVA4hDukXMq+u5aZjNHninY7IsIVBFp9dEVaDpw
G1M4aW/Uzt1OllHvIP0jR2nx1Tvx2q2EO5nkgw9XJUTmcOguQdPCy0DUraK/
vIGdOrHpryDyWUzF+5WcPbjVjvv4tvx6lPhJ2K6Mt9479tRYGwOTbfXmgtAw
8wdwT0qVyvApl1E4g5VuZPPjDfhpM1/LyAEwMKK+mQCshPHFbMkqIcbSIZTa
0QIvFwGeXzCRDByhRN1bwxOo8l5emobqXNpB9G/0ZYARzsHE1W5aRRVBtxQY
N5YJmVbZqyINMadMvbc+TLpJNtDsEohbqi+U3Sjh0LOxUZKZ+J2Nc17NpVQE
T0hv38DWiXRNCnodJuExxun7fDLX/80vyCwq8Q9lUDmJAEW4bvOxWoSsgzRM
NeKGZ/K1a2nQK2PZYuBSntz1XE9LYybBQ+56X8ir0UoiZ+aA9vtMO3Vea2XJ
y9CrtlX7gaChsZXc3DVQKZVW4QUgevfeVP2YCssI5yjJHjUs/29/KTZhDH4b
6HYqsvKGqY2CrlRbjZhSvaru81LJRaUSuOA3zw09s3cj3vCo7G4Ay+HrVmc4
f/YZnf324bZYSc1GFo7LQvogIo3+F5J2Gc2YzaqRp0l9NLHtA8qyfr2gvKMe
ljT209g3ImY8IG/p1YS59rFXAPLnxwNSqeInFf3DozyxDwcfiGXINZfc0AsX
iKQNa9+2BGR0qgBFAO6r+XFG+H2TZ9AeEuiAxbAng7ldeCyl+JQFRTAZcnvA
naCHdkvx0dkisddDCNWGTkQbMG7eJ1ugjNonZ1q/0DlENndccqP58odmWe3U
ncub1jTJrEJ7FWPd0qqyZTSRRPq/g+LdAtp0QPl1uIhNIcrryTgo41KWmy4n
SCBOXcQGm0+TzFl7AK/KvDS2/wLJ7uveGugS7j7fMKFVHjzMZK1hQP3c7Run
dwzgwz2rWCm96Sm8MWoUPiY481yRFYN/vwATbRlS8CwVSRapH2H/fB6nvJOf
YwfdY+7+cQprhqHmSekFxXVdecLMPNXXEk8Dvgpj5FmVdixhdcNL0aqQAdKK
WtyVvxMBUaBBsnuVKZL3HEqVYIYFEnnyn1lrDqwGXCe1WaD6ant6+dLxPHMs
IDAY9I+B2qftoqSsoHTNbNZ6NjcOkBO/ryh4tyUv7WvAsKNDvdJN+J1XSaah
Ry6HA9u7L0m+oP0Zgy3UPcLxlJsl0/BmDKEfW5WpRWGPjxw6QzqXh/lTfBxo
CzL8s6TtH9iK6tbrsrXa3wS1tyc/vGL4ObiexPxNJYmJHfWH+wMfh2vdBPOO
9B/afbeJKjWgWi1DYXkMAvny79vEKQpIx0k1ZSkJ5foviVEqHMwXHZpHkZe9
8+mSncn13G5pMvDq4zturedq7yjSDt7Lpyy1BAFHf4nfPX+VWQSWZlofMD2D
T+2m59yrKZcvNYEJ5I85CioT7Ve35DLrOou11vXVD2ouNtvimhKJQi+0lQ9H
4NWMfEdurL+5RfwI81lLqGVZX065MY5wnlfpEaqLkDQE7Z7Hu/0mqQTQByM0
GOLj2L9e5HnhdQwZhh9k09wr+19BkNzV2pwUdkBIvWARKS70wReDYbYR6yZ7
RuBbssMvZ/xUciU1sNTGeaWZIsjPBfZfTclkJmNyEupq0SJWYALiB9nQ2mUG
oc4XYGssi8fp68cVQQtxCsABpC9RMDDspeWajhKaJtPlAs6hOPiDLYWiM/G4
WRpF2fkhET4cG0FxY0izva0CYEauzutMq/+va720BkmTUc2e5JEgnKNkvJXh
vjOWpsikHbT3U0ewlGAO0CqxLpsioeOFHpxlFNDWQAWyNroHyIu3a7tHQwbG
WQMUD5+m5eDqDJscjR3+WC0dH5nWP/q52ODPmUdWBwNHIcezV6DGB8RC/Y2f
+ozPkWMDud3Ldyys2ra32bi2ch2yym5RXXglLL7qJyh2i+QkyQAeaKvcEXUq
v2zogJVw8fDeOL57pHWtQcYzAbr7OudNjGctAnlGGdIgB2XTdh8XCZ9oQUxk
sFUvDxG9L8JtduYuE9Z/TmWzEVIaRBqBGc9wdCeFeIPfEKESfUcPEWaGBoq3
YV04KOTYfqX+9nDRHnt6ZLgmTZnevlpZtbSpMIsQur07strcrUjbup31dZhf
uxTwJeeJB7YBpJW63BdumatbhzJ0oZnHKJ9I5iuVaufgH38KaujXN5132e35
TLvZBOEqoFSnNECkTNMNdmEDJ1WiLqEQQQ2u/KiZTLWXXUAcyFGYJkwBIzjS
jCjPar7PW4l4uSuuS4cpiN7eByRyQD6rd9xZ6KDPkMDjLj5QhYR29y4n/bX8
0pPT8b1Q+BrcCznNzp4pf7bkV7YRvWEcGNMLBg6lGZv+CEgY4W7XKykpih1k
asH8eETXQENYuSxj3nRqd3pxjAbqhgjsIT8jSMtJWygtnUS+uWgIu4pYlpa6
KTQVjxxkzJGy426xgyibcMlojPIius8oPv9958pHXLd4Ja9AbfdQyVi5MbED
6wu7PmOX+M2kub9cOm18AEcRUkyFUaH7Sgobsc46WTxCxa34KHne00clemM5
7V+z9+xmLlkXqcspksrqDMTzQP8HVQl0sPZTiBcnHBfeQsZwBNLWy/+OE1hU
hzB44RkxvLN7roqTO/tpHDfCBe3ykVumGOV2lZed0tN9PzeFGiF3RiHTCrB8
1YngXMvd9a7d8BVEVGj17Pe8wVBJxyWszYCU4aBkQ4f9iiN1iWvknXLL/UDr
/8tIsF7B7Y1GWsKv6ELQTbKDxNv9VgiKLFvIqnOcScCST/KIWxFYx3v6cUl/
/gEQ3cELecrDYW5eAkZXkf5Wg9twE5EQIMPR8m2JnU0W1+zb8INKk78wjhw8
tor0CMeAjlsR1HVOZPMZN9EL87Nzgltwjwh+dIxZae80NdFVlOWGPN4kBfnF
9SdMheRZN3YJ0004tMD44Guoz3yZQYvst8nW2B7NaNPURiGn6SPCvFJvRTDB
VvZNbjmZUDOC+FXgIDznmjkY4A+XxzCCd+7el0avsYH4ixoFlTmcbYAnB6Zw
d3uZGIZk8ZTsDOHYcqqP1dVlQ0pcumLqwXwy8kAgEexxzzH+GF9uJfFX3C8K
A4svhJr61td7AIXHN4MV36YTw9tfzTo2//SOw0wREUrAezbJNURNebzE1PYt
Cv1OBRoBEJc7hivW/Sy+6gRIV0yNccMU9cYXYEb3pPdaIx5kLajZlrYQEFD8
CS7es3q0dFoXjUEI0TGdWY88gOKXB02mE6Y1xEo9ae10eUNwMC+s0utDVGL7
CyeEz4UwhT+IeA3s5IvTZOR9qz0qgUlTCDgUUI9nJBD+1TKTdWtr0/LovqUi
el46a+Pj/1K7/loTm52qPxp7rWpuSVb9j9TspUyq0yTu5+5PaUO+ydmTgzNv
+aSR2X+O+telFJ8owqFPJJtCBIQaIoi34iKj6hmgyWLubC09iEe+4P4Zy0Tb
8GuGNKm7o3yTNNG2VQtEoqpbDvwoyisMu+RCwe9nhIZ/DDriXvmp5IlVbsQ0
pxcbF1V4dcKHZ/V7lXGtYplnkix8C6rRjlyiizV4A908ly2gY/Mnf3jGu2Zj
VCCORZtVLlP/LBJai4OjocAPCpM8bSiJbQ1K1z/LixIwSTcXLWXl+9/8mgiA
BgQVaozU0kOGa3EzZyUbkpIxFgI+Dl9Kz/Tf6VIhwMfDZTmEeGhK1qb5PWBu
D/oZBqSm/LyfjEY3gFFE9NAACTbhNLXgjXZlJJgHpVO5T9RqoAFSUG/UuBfy
RsONwz8xLWqk76jIjQiB5lm5lRDzNuasA3HPCXKLOttkiKpMOY3ICeCtIjrx
e5zZTJjqVct7UO65NYm0ThHH4dfJSx6Eo02YT8PFx3B/HeSLT4TKiOX0VqAX
tL0uN9yXe3CZXc1hDGcDB2PI1O27Ip+Ii7DRAmNg+P8dQCj1v8j2Rfcng0V8
xY23gJ/bt3IzD7xDln6KuhKDKUoQz86b8qiSwY2pHyEWmSIUnDkaQXDW7hdm
OYxd5SGe+nSonsdBWzxwxjnqG36OU2wtXjyZwnJ+HzVPVtzQsxXSt7/SJ+pq
Q969KnROvW8D/mOaZl0lN4mvRPqbUYnbhoxmLFScNOm9xR1tMejIhzj1Fdib
KBxeVSFJ6N1X5L9WAL+brmPboIcaEATUJtsfTvR/a9NqKpciHqOZxkUuHJom
csL7ZEf6M7TpIOzJYgUtbJ0HyKyF6vAArHYy1Qbbf/vfMPlOJ05+2ICOjZi3
KwR2eL4MEJGPhFXNpQaiRDhJ8QGErztC3oY5P1htDHGf3vmUEHoJaw9j9yVe
0h91s/QK0Ab50/ZpTNm0Z5X39p+wBlPXZ6KmCshdXmIDw4sMeukKMW6d2nfE
/A7nJ1uY2i+uPu+2DjqwXwj7wpx7t2gzHWnmmSo8zWZk3tSuK7fuo0XD6CHB
awhHl7X6VkWNj2Iv1EwJ7bBGSP6DSHUDCYY4x7PS9T2OH18bBVGEKRYkqnEv
NB35fFPHeRWRY70qSsqDQGaBQJpvsVn8tLJTXM9Wok93o15s3PMiqAOrQoJS
np6ovtXrOym4JoEQwN32hphLiwE+T7nGDRcdBxjI43Sc/kA0wZhD3f2qbowK
yu+h1fwd2eHxY3c8Bsry2pr5xXQBecDuzUBtff+lnrHbG7niep8L51v/mWxc
Fg54QdcNjs6Kt3WJxf3w2rghIBpviReQ7TDg0zCUqrg+MYRoY0vk6OrxTri7
lEQFjCszPkoKhTmsmwd7fzUV/vzWYfP1xlxb80zAjxVLq7aB9SttS5ZSW5U5
E1tZwatnL21ryialH8u/hgbszr9pWh0ypa731BerJCqo9eZyGivcRMq2uvy+
uCVCB2+IjddeadVJ/WgzplrzTfJRiGV6GNn2vY1GpKT8/fKrjczZDGKWNWGM
SE6IOMrWMH9+UEee8jJ+RIATLi2nkacBF8m+zMAzmCpFP8X2C8KD1+vgIdn5
M2gg3M+XlB1UCvTeUSOtCC4hIFo5/lXLyVwuguWTuNJ8Xuu1OCDgbuFR7E6U
++cAlJCZKpfUI2fAztyrrWH40KUjhAGwX/AKq5qLE2D59MzGFPm918B50mS9
e3zPyL1xhg0ypsC7P39v7lX8rQVHwLKd+wgPKpS6QKrGKyu20nf163lBkGoM
61uwhAEK7uQTcfalEAsQnegwCkJHsljwhIC9gf4caTBmmYx7sTYQxBXQbShA
lsqrC/dqcGoSy//+ct4aNVsXJGD5xLVydS8KnMLHHaWirub6RTTh+u/KgAHZ
eGfs3+ou3WmnkS2E/Baa9mSNWHu6DV24ovc8B6tlmrESf0ORC34wKQ886uKq
UP3fYQSFqzynZ3rRWpKEOJoitX3xQ5PoeL0AX4kJtxbIoCfRHdREgojK6wV/
skQJXBmWvlkJAqQ3y/2hzZg0VXfVwr4yNu3SCMuW7gxRaav2pYZJKv0KFCTe
T/beE58d3EqtQCbCgkm/uvPx5LOUJ6S/ihfRTyn+JtAh2dT/xZceAwoOy5cm
C/qpm2mmhFJ+weSXGSaBOuSGLB/NfMBz/EX0KB5+Fz/SnRYliTYYdGRMSCxu
hjbGJk48idDNJtZg0Y5/kvBQXT+FU6I4YNrDzir6ERENXjqOvHh0Wty9lzKh
/EkFpD5A7AiJVbyzzmKr3jUIvp1LTlP4EB2ifx7FX5k7rhdmmhXN3Psd1lHX
QbhryQ4vymRfF8KRQCRh+j3mcCGL1MhKnP1sLn6ZRskohi0bjbEjmcyaQOyg
28gupCWeHyy3p/Q4GUaUV5AGPtiNN8lrw0pvFQ9Xwzk6B8UfgfYgWmMkJHUX
Rr613FqN/lYH92h6Z7x8k23Tfagn2S/L7wqMVL9uiAOoA3qLha7iBsD3HMC7
ieVZ7GhJz/CkeJRIOuuCOhXtr8FOfLxHeQj1OlFasUjYOWfwODnwo+xys+Np
BzeaaKWXeOTR2Nyh4FDfYirSqVmjTU1u9lNRWDQq3+0u342K4aIW+uUsJYu5
bxkJYSHCkbfzoR/Avao/xqwdea+erI790lmopRlzVw9hshOjVKpBnjcZf+Pk
J7IQ6YxKtDcX6j39WWHIUidLIhlPGlfQsFOJxWKt3nKMSq7oGdtNAWfe2ieZ
ZtKlUimxhoZzE+7ipV8/Cha1QyFJ/mx6F4E4NJmbuY6Cnb73KVVI0adXVsik
hT5wi4ooVU4R43RBiBWomkn1bGneuMG8uno7qfqyhsZskNM/XNwCU2oOUcWd
Nnyojer3NJqAiktHUMBZZmntmP+n6MVI46pGvfulfUTTsUSy+CerHYAgMUmy
53JPcNfqweXzZwYS/pLzEFSb9D/CxC9DenskySyhJYgP7MjPn0NVn5i/qqsU
Ha6PyPFEvXz6cDDAH2R5br7R9pShY0Ix1WX0Q3f/7LO3T6nN9pzmvXwzi0Gt
z8K8+tr1pENEUd+dkczsv8Cn/xhxGDPGu3mK3ylxTynQf8NuNBSKr5EKyh7q
HNeZDSA0Fojsd5r3NnQS4lFP00bbWbcLROV1wAgHqK2Ts1Wz041mnc7LEaSJ
76/QwPLgdVdtywh3t6+fzBvNQA5PNkQueWbd9RHeWwmX9oq0+jFAjVSsjWTK
S09/Qx3GuermjfF9lTw5+wSEyXi0k0YtlRtwVNLekjVOdQ3yBzdRXr3WTOKo
NAZpfgvJsTS58CTlwbuUm0aRyd8+c91jLE08dz9NjoJUoALKDk0CPDvv5RFx
Hw3brDhmof8DJXeC6UEcgLYcB3iOXqMCgJvAmLLthLkjUVncxCkukp59ryMS
B4ray6C8db/T3AliPndau+ebUkeaKIh3V/4IeSuRyjHQ+LhJzldyY5hokgeN
G7KLmbWJSOhR+MY1692ZyvnCIAWwCYKcu/s2CQTfM8Hv/MS5vL+geB219z6q
kDnnnoKz/RjOnTzD8O3LS+bzer/DJJVdH7h1cs4Rxj44ps2hwpCJByK3ZQMO
WUkBeG8g6vG/vm00Ld7bhoIBTzvSeDLM0enfVqLEgKSWWrbddK1EtyD1MOnk
iB/NZ4d1fmSiC3bFhiCtsM84mGP/J0cERJz33XHfmaHEUI8EkxUApaZJNj6w
3E0QrAYYC83ykGffWpmKZ6E3BlF4qhymBiZKy+QxcgeVErOheGOfouPEal2D
05t+lSZzKCLs5dVzZzaRtZ0krA5nm9Z7OZ/fLYqBCfW+MsZJikTm3Z+9nOmt
mR0+Xe5V6LmCad93fc6BZ6SHyiDx6vu6VqEM63BGPwe4Tewf6PT3fpFFC3UB
WGaVRoEO0LQMuqcY7oYM/KFMEbfAZjnJaeDeUPKfwF3ixUYWehqkNDwxiJna
YBcr4UqzzqAZ3QUTjJ6AAb/OlMhAHEEBTnrVpyUf8r7sBzcT9BbMfB1PrrsL
xygu2IMF6YQpuDEUm0YURS0ToYZO91RhypKf6Scfn/rdVW47GxRKLk8aMLbZ
cVjMCklS0ckpzbW1WkwlbzF8Z9quYAL2Yo93XqcSB7a9iAmdU2X3G+Maxtxm
SJE3jEKZnuehbMykMDRO708kYvTaepM701GpVKNpWPPRBYm7tLiQC2SG1+lh
MAI9YM2aSnL5GZoMCRzsSWSL5P0Z2QMPU9WbKhqPYqqU8BS/3FYmfw820vYL
UnIr7i8SRv+3KcXCfD/vaZaYtk32+Fys3jDYc1NdZCre7E4WGm/jIYoncwaF
FuqFPGejlSlJpRFlpRhCTlTvidW/iSZaJo16wNCeYMde55f1q2nZlunT+HCJ
c9antONc7BVxNWo2/XENqe5jh5penkLi8jgGiDbjKQfoDJ+KdZ7tW2aZ/ZrT
BDk84DyYOA1oA/xpMnA+oxjtIjdROby4ndNHbQplNqFEgfhfc2DKflxg0vv3
pKK9Qb9Jpj0wog0ItVAjPJPq0EbKHN9+1QZRcWKMZPWCJug3SoUFkvzYpHsa
8zpHl4VOEA4Fh1K1IfL407Dm4Pd+A4p8JukeISPHCENZ4oIU7gUNXH7BHsK4
5iXuBrFIPZb3+RiOGfqm8lFnsNRAgGYGbk7kYOj6eqOIAXVgWNOJ/VzwxXJA
4qnFhoyURi3fkiB7Qw/3rqsMRdlW5gC+MC46baY1F9kcmx0tL/ifmq8p7bTB
MLuho5bE6Eq+8UMytj1QwIWm4wwy96S3S9Y/B8l4bnvd8KkBYmuFCNI9Ey6m
h9kb8umbyZsj0RXlnXj2A08yCbvYQB5IZ0TK+CrbieoDjTn0N2vwTQVy6HIA
F7ZwLb+Bdq54mYXYp+Jxwmcv4+BL8rr5B5QIxON2x//fkF7HGzMBAxY7DRNq
I1HKqpgUPxPpp2dGm3fNZxTZI5M0xnhOSUA2CMpgWxVCYcLzl8N/Z7UY/7i/
lkVlRyqMNLhwLuPGWLj9yDNEnpnzrHTNePFP8thePB71bpQOIJEtsV9+BrcY
oDoX65gqAeu7QmIUk9mP7sR64h8JABE/8r0l+fpISyVuVCvI0UKWZpkqvUP2
POLjKBeZ3hcywwIDCbo3FQgTcjsxV6fAaC7cXh5OG+/boufOnw1yM6wq43AR
jJWH4D+ZdRh4IS/D2F1pjh3Qj0cYGy6iONfwbU9wzwQSWwJGvbo9RGQWiAHb
4RExCsV/V1sq4NiV0JDuBLqbRZf8BcppZjFTtlkPRYwM5OEppf/QS7Ct6wlB
jxDQY+ciR6vbFm3VDhzfjD2Uh+2/zAkOxngo8rTlbt6jBtfSf1/uutNbq2hR
s2T7qsVGLo3dxSq7qxcX1/DGacQxy+PcmNAd9bIRidXUfOPPuQ83uYv3L2I5
GBMqPcxdy35dny7n+x8CEJWGG2SjoEwibWwSKe4lMrm4Q/HmVnlOO7z3rEaH
pm/Qm3jp+vJXCRZzaG6fJJIs5LmqO9nVaWPzUVAUi0HAj8OhGk86uR6GnCRi
dC6c6vWa/kG6vbB7KUC7Fl67UMdBqXFSQw9Mh966d9Gq9aWKJURSSyhmD5kn
JhW/HcBGecwJI2jQQXMip+8ETsoYjpJnov9dUdrFMoJDhuKuRAGOi7v5fG5r
gm97BzgwQhm4gTgXrYeibIYwzb8NliXOfwrrSVBxOtDDeqiosYuWp5KSYJ6w
MlUwSbEil8tbPd8xazfgIHipSeLZJUTSi3Z/cw/ste8N87dqIEF9HGB6SURZ
z4PeEI/543Z1+UEYAYjE/jSYYwg1XWNSErFGk/KhHgs9sZ73wDK+lyWN3W05
dWRXLwkXrWYOpw5x1lvGUmZZ/2PEp+jLku52juhpHAxzoFrfNhZ8zRd0ueWI
St+/kK5uXlDOy/xNhY8Ufq3/w1TSvFbIqK05obDT58EhKxbFGISoycJedgDo
CjGDzuorcNf7PyqXD5vioNXknsC2xpcNLtmsfNI+jA2bkfcSr1IaLkVWaM49
RQpU6Y+sf2VUu6Z8QphElkw/P0EyyK9B9XP70u8r59Wfpprc7wJtn5P1N603
a8a2cQ/1XqsFcpB7evHSBXIZmyhEPEPprj9y4Yq5oaY2J2/x1uhA4fRByN6X
TiZ5B4lLF5Vkgn0MOaHY7DWNWRbOjLwhgoeqrEJqXH0GeFvjQzt7Owzo7FzF
6gOSShHQDMmPS4L8xsA52NzxjFHJt4IvPIt8XCpHGxzwSqMw+oBn0LaiiQav
gvPLykLSIhRlF1KUWpUDswqR+J2wolhu49kyHOrJSQwq/eYCTldfHIub6iPa
3UxxZYFfvS6YUigb/tczxd0IZ22dK65i1ASS0i1DeW5NBjLhtLBZlZPbaQcn
KUozSG43PR7QFd7ZzfuOppXg3+NLb2Rcly/cbIBSPOzTAAd/kf4GtULFB2ZQ
UGxYqfKuxTCt4Zti3i8Qh4ND3Su/ow8B5hxK2cpen9EDFhJ5w60OYYBTvgV4
ORJY516fzoLwo9LN0NV4zLUeYJk8qeLt6PbmIseOc6+I8WqtDc2nZmcNYJcx
kkPSpN8ZLXl28cGV1xhMX2yEehecfbuMuElOcEv811A+K6BnPvCJPvIv0m4w
woGwTpBSIhKOh2hDoK6G3u0//wPxxNkwk3y7Fk7NRSXISjTkctRyR5Vsvo1z
1CcbAtDp9Ej9EZB/Ida/xFwS78aKjsPq6EDpkMi4g+R6Q05mu4yz4ELaxhXP
ImID77q0pJzo6WZra3kMwF5wlBK9PkOFYmUxVDaXB9XNqCaj6a/3TYZzrLrt
3CTdr03nSNVgAV5zIwJpw2ZhTtauFbUDWV9mWd0vRoXNHJM1d+sJiBUZXwTt
mNveFLY0AM/mN0zgKHJPgbBAoqEMYo1VNBOOnIK9/ChSFWXOXfd0VLnkLu0l
Jj9cyNZGWmW4TTionmf3MiQX3jPBuUzhIZ+ajJoeT9mzdA4OlqkwcPNgcpTw
50BHZkMl3K6Dph9KrvKlxPRQ7mag5rynUf36zZhJGg3nulPZc0FanJKdjXtJ
CmM60nSwDMSsaR/vcbD2/3xpS68pnsMnf3SuiBaSOFZXvkaHfrzeEqTM2Fc4
NbUNh/8tdFWFPOaW9Ns8nfXy6TbQVS3UZJIGp6C5A4aQLgbid+A0Xfo/oCoG
j8msnKE7ISinzSopDJQHnbJaLQXJ+PYXJ8iXRiuBrQFyXq3JOAQNiH8F/T1W
a4voGkXp93oO/tkeA+NIPN4Qn2lYqA0O1/yIYkdFFCLQ5qQdPDcZ4AzY9R7Z
Mh6BBM81Lr7/MsrbQks9jFCw0Ib3yH48tyhWGX+tBUHeYEJCeWdpqpe39Wfn
cP+0/yM5j8ifCWIpx8y/L3KBQxVfEOqzA+gAiSXQBVhH33abJo/Io8kx3q7I
FMNgXb4TqfggL+mv5Cb3sRCfrQ4Ta5pvHr+UkPjb/yXq5OxooH50K79cHrbK
xiGDLzN5l+VKan302GMxsLEzQNKpDoXFApkpjsZjgo52lym9u6AGWuvphIw3
pzczvK9IJUILzmGY6xug7OJWD6BKsm7RhWgE2ZTcV0mMMACgR/KPPiTkP8bk
NcTb1fJ6EEeFQleZtLg9bG8dTZ52slYvntdOb1jgv+vjQXtdVQEkDiLPBjLA
rMPz9sy3AmuS3k+iOvTPivwFPLVc5+zytns/E8BvRfNx0UWwuof3j2xulKwV
mgNP4NIoeG5/DsLa/Rl19lyRFMs+4LwqRFHbb/fzcjDAHZQ9+/G40jB8VMzg
PIwCfCb+bzLL2W3I42OdmNEMYZNGlDKAzFyoFED33qmdUHCEXfLgtB++14VA
R6WY7+lDtSv/CAjKpvRl+SQqB3XMQ4WmPVGpQXCkd8jy2Patgl83/Cu91fxa
3UvmBhy/D7MNOB6Tm/RGOKMw8JUsbbZVCyTisgyjjjbEYNRAXp72oM+Am2eL
JB5fBwK68j/kdYcgmaKYKwTwqfEhsVjOdZozHNXEM5FGHO10eaWo1QkuRZBL
gm1e9Ko7LeMjaZesHK8gn0zYQTzkv/wfdNc0NCvnIBbQycxp5TFcwwVgGqs9
twoC0JnL42MQriG5IE4VG/jpYCtdwYRe6IKyREoRpozC/JWZ9wzE31XIZVhE
BsznnZJXjYiYLUgow1yMn77dcGz7eNvQ2EIPyhuM+6sYEdZYh26koZvqcVPk
UqrYg/mcmYDE8HXTVEdTvNBUSrtcbHGRRzGo9xK5LiH37KyXnbDAvr8x4TA9
elGipWykIFtp3OMfo8heWN8HPWdRl/sTxgKuS/g5K0vYsv4dHWbK8/79yXxq
rAx5PmIiG9QXZOjbDLZdJZqI64z2MYnSd7QbcQ7XGUL/2bTSXvU15PjdrDfL
2F/8b6oz3E8IWrCm6grF1zWCxtRehTyfZE3okeVUAV1iDSK2tNW+sqSoB0z0
bAOenf0NQ6cYeSzNdljyxIDBltlsXMM4bzMTRWPlk75PCo9dpVY8NE/Fkg5W
nPuztuy4ksK1BkXBoiirlgA5Ktd2QtxOV/edDD2lr+0e2Zne5q9IwUYxTcD0
NvYOITuDZ51Hwmm4sIW2dwfjp4RY970NHuDvsQOsWHryVwLjzVLAHz2GwtFw
cEaH/jvebrgU1IwN95xSk+bK5RlFXDxfehLWk7FeF+z7JSV28QGjDOBIQ7LA
em6Ou4vp7BV3udx8NlTGd2wF8N20G3jQISEAaoSIZueaGviFI1KsMfkKT3eL
8nwfO9XeqUBE8cntRrb2vIcQaEtLXAl3ffxv2hEQM0qQsj/hgxe9YRUMXhEJ
0X1ybMAvBtbKm+iewQHoa1eO99UoFPi70cBhL8vFAh2Yng4eAvg4elWckUyw
px6k5Mqck2fep5Pr7ts5MaaSLHaSwFoUQXevYXOh472zimz19a9TvALyvzt+
CqEjmQ7x83vCByuDTAQieHaCFXwaj89H29dn8p7IEUlPftoPbZl2w2jOjaFG
eVNOlfB8FvQ8gj6Evc8Sn71YIYRIAe5JAk2vX02rwMcfEYX7Ja1TM1+N/qUB
XcpUoVQHhkSexofyPucC2sOyY5X3smCzStOiXAZ4w1n+OIlMQxXCOT6L4mE9
7X+2YvZ6EXa1m5vqSO86bTj/Z/ksURxOLchvk8nn+HgEGVDilbjhvmEvBo9F
PhvUNXfj8xE15HezGQUoMfcEopMJ6H6s1T3x/gaWMVqtEL+hgPCqkKgUXVsF
YLkr34lSsUuAIZCStGdvio1vkmgDaINLtdFq2o7HkMro6VcbG9wc6lj8SF8C
hsaCbFHqOqzwoT+4upm5CEkdM3lQAgTnPv2wwqv/zt+ot7PALA7MdVUyVpkp
TDHdywNpqPMEhuI/8nwBBF862NeX/dbnymCtTVKKrbDXayEBeLVGR0+s04X0
4UBFqRKTrf258yK7KqAjn9NE/tfQKZvgqdrDPKQ5cnUiIRQw5JfrIhslT0jr
FKXe+nEFrAi2H0AkQWqgzhqbixuQH3Y8DsKtlPMprqF9f0n0JyoROGHd5CP1
xIL45ZvH1lWfvSZ3rIevXe5TrHZ4oIR3yh3+JmJ3QxyW3K+vsI4n21SYrHXO
7P2x5h4MIFeRUHTgm0SjuYkpL32ldaU1FoH/+/7Pdqf4oacxJ+1r6Ul5frxt
LB3q5dbDfkipORhOx7Fh9IH9G609SJdE5EKP0whze2PHig6rPwAqcTwDpntx
f8s8gI1CtxZVHSnSSbsEaQ0a1az0mcvplkUPqOfOySb/qYTgEWpwQ1kH/ntJ
2EtqISeLYpbjYyA7oH2fZu+fDca5LJp0yXz+pnmBueOe+WS/8EfJQdpTmjRA
dGtXmAwemcdKOo4B99nkkQe8p7+vWgDZ1EuOhHUXDQ+LWmXkzMgCffEsDnHe
ZK+IzRgiLh+ghj06nNIzPK02/Vvdy+NA2YQsZvF4pvnh6bq4AaSXR8CNp/oD
UNgzWmG2cYoAT70L5MGt8UTtA+uBivbrsi3GiOg1v+VHZrHlgho+757nMoVk
nsT2wCvfN7r8GmCbKBDLQXbRfas0WhTTLF6tmeIUx+1sCGaGentTUZNzZpxF
8Ni1oW+mp8Fcl/TorIGDCMl6SkZgjhVxImfJCdiZhaxJHI1tA5YAD3yopOZd
wrb4A3ThI9ddkbOnLVW5xROV2atgQQuEGyzGw547j53tuCm2YVfpUjUa0ViE
oLjqDatmh7Y1qgvKLAwRp3Myhb8mN6mt7b/3fwh4S9TF1QIVtfuhz8jOXmvQ
Qlo+MBHbHSlLFNrtt/v7e2FVAWDO3vUg2FksQd+PvtjjAtSqYh4G7Cq+q6pN
FL/Nh1hdfpWjhFp0Dw5QglPFEidGFposr4pe/Ohgq9nghPowTpxF/nP2LVdG
xXrNY4/sIioGN6g889wJV0H65JfYioxZ+tQsIzsEKer7P98gyhROkGGxGEpX
27/3PyPM+FdnsuyJkJnsotER+qm5mcchLOaAZG1JZ6c+9RZ3aphq6Bkw9eC/
FZSq/G/1jO+jFNoMyPpZt+xklGeD1SPi5rQpWm24THzPgi6j4bpyYqOpAkNB
z18tHj+2pInM6LyWBUc7kuiLL9BlVQGCOHrGegX6KlPZBSpXCWHwHfGinTq4
YRV9ouuSbBKxMdfhOGyn/p1uDyHoV5qEV/7WjxEGSk1bnbbnrkGqNSfyEKKT
6vwTxvGIDOzWjW3VaRujcYm/utUlB+eglcY3zvXoWZikdAdsPzeyZcLdXCgg
Wmml2tdQacsELeHzI4vP1IusXtagafoeSDyXk+ihf8zcTBisaK9alC8B9jvS
qK18vkJtcIiqZD4fAx+RGhnn/YeomVcJxCyXOaXyhXU0gaKqql2sWGowWMJj
ELvHo3FoGAUGeTqMiryXECXUd/5W2syzOP4rOnVE5Rawk43QIDcqpeCyKHle
UDy43ucJ+GZchiNSUV2QFskCoSz5w3tFae0RVmL82aIkkx3HehdO/c5x4kSg
U35sB4OU51dfthTzN7WdwtErpNgXZbQZMTVDU4EIep/am7pvBAR50c9/SbHF
5fNwIXkeR1TsJz7GNhiXNQN6YymVvHDGC9wZczoEzrw3TuaNFM4mNJwSryn6
+SeSEw47hFk28Xj+9Fe8qvcMTUFboC+KFHWtRUX1K9oMYd/85CHmDUUNUarI
RiGkyi07N/OfgNo5QJdTEDo4sIP8yCg++zJulkVDrGQgsqBcftLTUWBOLdcW
p1xvC7Xm/UWtZV5+f6FhuS/nsjXrq44qaUTGPjuIgFfkSWUzrd6WZIpUWmwl
6mERsXtmZAbGrcJ6uZTV6VjKgLpsWVbTXpV8OzIIDNVhUaEWl2GJmDx9wAmi
KSoXsppYTbvoSS+54OBN9zyuYnKINxgkZH80IV9NTIsy0mqdWaU2LKCPRxGj
SwR97Hn5ZdvhW7JBo11uRhQeHsPPprej3OFeulw4q9Xa6iUOHYHokkLtL8Bp
E7i/aXtkqHe9lWOvVKKThLQYIVFsbDEaJNRBM7l4BvEicO4GSvhXW77CZWSW
mtcOayIjZrguMS5oA0ksT8NWDyPtq1S0wZYepdgIR9dMgP3qwIaa9R9BhxDw
Xe20sTkKDQaK87Gj8jaiEhENivBAmmtNRmDOTipVVfFwBm8wGu2ebjxRMCca
ozy2G9vCkhJ9ufUy3y6zWC40KHmmMvelp1UD384JUm0TCqj+XKdA6hMQESET
Z/T0oPkdfE/mkMZgsHKeSGNK9Rp4DIDbvT6MeeUCkTvbnn75u7TtdXtCqu74
CViYKb626jwWFhH4gyvGCrYnSfzO5ubyAYRw8kTmReUM+mm0cRl22u9DDm9W
6NWvrJMGCXiuLb4gpmxydE1pz33Qlza1UukbhHJ1F1jG7RvCHOGIBUIlJe5X
g48fFxT2N5Pi290XnuAPumUT5ENM1VHlK1Lsgj4c0ZrA21vIjisad8FYjIMR
SIwsshHx+zFbKRgXlkZIC4RoYdpq+WFvM+0V4U9fCrJF6NCFD6EMRjUxwDAX
VOaBcFXDn0wC0GthciFdH9en7V4JWG67O2eQMk0ZYP2J6rJNsa+MrxfoKoxB
9rwpy2TtKW8PW9wzlK4lTqVUPijuBCFdfQ77hGAPbC7QXLblxC2nscbtgX1F
tMcD2VEAtsYjhHd+IB1eNd26vWU2TMSw/ZozuvnGsYg4aBCdTITmHwNiMpE8
wMR1QNl+9MAiH9ZOi4MfpsIcmH4sSwzQGTWUrurfbcWTXdeZhj3ngjm1u0Cj
wOZrJMf0n6d2NxU/av3SCVLUPXKBPvi7WgTBnNqzhm0afFYqNCXheENyhBLJ
5gd+oGCBS7xqjCOdqcRkmKQZpmhs97HtuYR/qf83S7QAM6KaDXapDOXYx1u9
8Sj+OEUNceBdbqZUy1Ygl++JE4LkoFhuNBRJwi4lxp2CHPhGMcMB9IEkOEsr
7xN9ThUFJhovUmEFUb3Wk6XQylGOiOe4CGLzvlHJoKUFdQ9i4ejTjPUogAMD
HK6e5jj/52PZQnTeNIiHiJmPvS9+wZ3sL2c1tXCWVlu6Zfre2o3wMDSYjENN
gnXmumcKNYHRacS9+omHGzT7kmcB71mn/yVL9LtVZEzsQYpWTz3ZjMQAspOY
ngPN6JDFd7hXWy1/RzL+jdrsl9T2mCI7YtAf14FR8xamKw/rlBELXeVLbA1C
cUEU8sZOQfY5VLE80ZFTHZ2VUMGBov50kdF13dpyjBxLOZxixR1UJY/WkB5R
hpQG5kbc0rQ+54oHVXDisEUno8/fAC/EknBiB+5htNbeKEyR/MbTgKbvn1lA
+7r3n3a4urAd+uicbdBy1L9n6Mv8Fm33+25UvMZHyes9zBtsLzLl6kasKM3M
ttpSpzqn/JnK0+K5qsuLPzzy79pP+98v1HyzEb+kKmwbuS2RwjkRQg/MKtIx
LgLFT84lmwk1gjXC0391CvR1Go10961glOhb53kScZPEOosk01ym8acHXFM0
e6HbzTAJV2JRYv0jrNnqnFOSwbwUN5WS9ZgfXgYzWw8XiEeTaLlNwPz5+lqj
CZDYb7Frq7wgnBmlk9+0k1F5yvjWQ9jbqm8eWbZNevyfhZA/pJ4cuYKjrWwJ
VKtMi09GmwGuTYdEYrSh05F5nz+uvso7Sq2qIilhNid7yRSayy4WkgFLpMUZ
sY9f8vjpNo1cZEB7wiHzZhcp2j2r0LeaqXukU6dgWIk8x5dMlsJmoJYNXQe/
SBWgP//3a2gxO7BhgPd4Ee0lnOeMerKbtuTJVAxxRGjMpxLTj93PJ5VtucDC
Q7a2nzM+L2sEBJ9h0v27ucfaCVI2I9RA5H93UMlVBjOcvIw741IvcrFOzugl
N2N9h1J/RYiW05KMWRt1n8uHkSh29GJGtRD4poX08ExP25UC9+CQbwYiORjE
Z7z+CIU8VxOw10u1G8yD0tpUh7u0N6oR/dunSqrDxf+lTiVZTgSw+sbvDPgB
WlDA1E08ZVzwRfPTQnbtdnbVWLa41nD8hw8bcQ88GLkvHB9zwkBcpWDpYlI0
PzjCtoADRmOH9D5wUdq8d6FFFxVsjbUNfrPJHdYo+iYhlQPEhZc8D2YhQjZk
n/WkfEYAWL9t3rwBrnyVgsmU8xjet21URm1y5fHYSTC/3dwS1igH/ughym9T
eb+b0WEZpDKfKpk6vjPVzPfkm2lgJe9WcSkiCLSq8dEpCpCFaCRMsK8YVCYn
zegpOJgGC7ZV0fP3zzqzLl+EwKrVFtWJUvT6aOX0AdR3CvFQf4wuP4PRZWeJ
7M+u1JRx8P27dmqzwpoE5loxb0Ya6e8eqtCC81kZ9/E7UDV15wHveukJiSW/
VFaDybYnmxUy7+8dqfkIaV7aQU0EsdUH8KuQkBXEDPVjVsO+b+Vuki5lR67s
SIiIRaf4RwmaCp4KT1BO42rvodLNOrTQflKylMeA/g/a8B0+KUDPN/3q+c2v
jE/Iq3zqxwgHYodikaTJ0+UbtrZfm9AAUHrm/coBM5YU5a/DbLkd7ZVygelw
IsPxb7mlHlLtAZjhisZrUcV2c9xOZG9t6bemj+CDd48HMmQN9fjrMyVwHj86
od99uRA74DeyHnJe2JN2qISwvGdT0PTaVBCXArXd97PcBZg4cCxqQ4jTZKnV
2vYn5rx8JUkCE7eVaG4L6/h3dHkbQKdxQpyioTXFUMDaTB7CosAcexLgfNKb
WAxQyw1q9sOabKC9Le7JP/TPUpfwdkVO3W1+LNLRHBMyH5CXmxmCnymPD9Cd
yDgH4cTKI2qvt0V0fgqR7RnRvL1EZwIE47oaIbl0fNPAbv+D5sbIcmKDma4C
e0bC/CaocwQULobeyWBoPGYLRmQKuSymLST0cN1jcOrXU5dgwwdmnXR9quiD
/k2pZIAKDUWpYFRGihU6ZukUP49ogNl93C/BVDANmTCGcKM7rz9wgHOuRB19
vSPkJ1DImLXFsF4e6542R4pwsBTE3fzvJbiD82f2S+i1VEn7MlIjCKUL4KW3
hcLd6nipNxz7HtpP3M0n50DvsB4tXcRIrDKkKPZ1SENz9sohgaMhdmdqmDzA
HsfeX8tqshAYNLyFEw8CUlThlYhuGLaYMpCbFkZFI8H3XgDJLsDycp1LZSIo
y1C07zgLQsEqwOjtJFlswM82U67sXJqw7XgjKhvHmI+8nAnI7pr5xqQ0N1Ev
3teQa4XJRLIVbYPRBRH7QfXwUuCc8beF2PmbM5Vvbhap0CV09qMdoRl140e5
6Itiq8Un6GBRrjJmdDTOz8dSCnyGCt5m33B2W4Tj9eZ3X7STZt7J8fFToMPI
Fw/AF+J2C7rNVYF8fyAlnN1bhMRJ/dFa7vSX0UG5qHUs1KP2mYIrDkxVwk1q
co/g69i9jYl+vb65pI9MnbEJ7gWQt/IjRi7Hh2J18YVzjxfiiLw4i7gWTPP2
eLHBHqnhJ9bJDop76td9+ohM66VcX0mLq8+SxJMmaXreidpPcIRp3m0ooeF+
xMV7wQYanipJgfmrctfNTaZDdgplqhQ8SpTV6I0kG3E8Fk41a+hxIp0A5JKB
gsFzEEMSpNtDcElhYli0fT9qc6j95zixI8M+UCuza2ATgMgzuak4AjvKrb9f
bap8kNHHowisHuF7y3LWzOK9yvTSy18MdgUNlH3DlNIcVq86dCGm2/n/AdE/
izDElna2+efp5qCbGEBxfvBBaq+M5jTFxLJNRT2K8l9j6CWvMMrZpk2cxHOA
mJR7sdrmHYZnU3raKJA9qgQd14cHn2huRF6Sx+ym3nDN92+U8o7ZJdl0tlzO
z6P3gRKA0I8wb6wbpBTKyUkHUW0bKLyQRhFMs0vsIbwOMW6IUM1+eqXGQP1+
QmZjX9EKQfHiYNsr8vYB5KUjT+b7eJ/IEmXpdDJeeAaTQihEOBBuA6DzOlUp
2cEuOWMar0fdUWyaT3MEN2TSmdpdDhRkfPoc3znljF3uoCmYWAeoaafcbwT9
qvameaGWGtYeyOwoBlzO79l+xqfr3N2P/uYV6eFLVD8Jyi960O1dSl840+01
7ql3yKpeUoQcIBMt5wtWoAYPq4XR8Jmi+4zVALZcxaYmURZjUctSGteqoHdz
lK1mS6dwQGs37LNk64gCcTKstkxJlmGzCnFDAqrbYZJ1RNNl68DAmybLgMLK
4HJSr3h6WvCPOgj8c2zJxSlJxAYS2ucxIrr08q7ne27uHoZNDhHwrVNHVLxf
rWhAsjEcRcuYydNyXDnTG42mv8UoOF4gIc5A0LVCvbovZ+ZEpDms6d3lWtUK
8Zp71mlA6Y020/+xEqB9TkN6dqZsKfYu62oCa5iAlrN8AO4dSp6H8CLZMH5F
zcDtyD++BQvTGLvT87XMx5AjG1BXtqv7bX3yZ5aJihUBvcx3FUnK2vEsXBAI
UavJxbTiXI2kWjHw3gUpN2GmzSpst/+HcHuggJOzGIcMvX/8nkQpyxFPqo2R
NN+e9lC8tT0sMDxCS2lI1hOM/bk+Q+fRHj4s7gGrgsbycImxbJ5aQA1AkCgt
T+OmO09VH9AFwCrkQXbIIuVB6nZINam6vvQpR/LfwUOwqMgYUfg8I4YkF3DO
nJ3TEVhUHQkKzg9eiX8jkfMpXBw5YXUdyV7jb2/tP7oYvIR2sxrcTFyh3+l/
j9m056o6Q7sHnDHDm2p8W6WG9+Olt9zRTik/0lNRjLfXkCLodLIOGRB8QuBm
yxj1fZHtfgWriFKBixMj5i1o2lyPn6ojUc8rZ7GZE6mIBIpZVdtbabUFWvPy
N5LUn5LebhJdzOAKiBSaHAFgiIEP1AXCc9dbap3iY8Zn2bvqQSU0ai9oU61Y
44qxBw23Mq4zsfS41f8vO/k6T8HF5HdC7aXTT4qdKTrtVvqALI/9WHBWsuwx
n3S88Jweo9jFBtNzf+0Vexs+IbykANWmTEEm9CYQx8is3FVENIcfoULkfDa4
6/y/19AU8uFUEhmnqKu2JWZ/RW5h+8OI17of9BBFSBsP/X59Mxdhp+ocSOnP
sduWeXwJWwJD3r5zh1eSSEtOYVfRWtvV9kKULZITTvNG5beMeZSSKtYyyMc5
G6KpDEFHzK8czudSzoOdpZZhjafk5P77qq9RWoHq6fHSCGDd0xIhWOEgHT9J
dgjoiLetkOavTPuzn/ORouQy3WsHHn6aX5Gb2Qk19HaqbVWLkGKYtBwAmfwH
BaEszUwTgA7MWZkSEuLUNO2gaTMM6PnxEBqts58FDvIUT4CIUfsUEdfOMSi8
jVXw9aNXvdtuXPampQWPKkuxqZbb+G4BxaUNutb1oIu/PjfmHESfQMumpLxK
F8GhN7nnKjaSjC+tSbNYImGJF6FpIi5RXmHORywl1uaUMoT8PgqCVDxbKgt0
7RO+dsQEUvbEERpbPDaMgOQmr88o/Qv5cLhGER3T1vtVutJHoKRK9YfOjSlM
wPZ+MNbxPT0QKhOSiqlnO93YSO1ptMYyunv74eEYbWZbcz19PfPgDr2l1OTw
R1a+ra1RzBWg7mC3XYzJdzF7SatUgnGiv3Gb8d1GD6wrWTPGdwTsr1rY2ofL
hfAE/Rb3xiD8BPhhlk9BCijQUJxZArS6GLuAPQGPYzqW4o9/pmpq9gUh8U+v
AaTLN6ikB96CL8ZUbT6OSP3gkGtyQ3BWuakf3S5tuNsglPqRaITylc4l4p7U
r0U/AglR7H5rD/7M5l5B9VnDvtm55sqN/HVTfdHRWA03ST9Nf8ZiGXW+6oaR
J/cNZT8TZzkeXVacvpYWVep5TaosvFv48RJE/9vA3dbC3IainlVmHM3F5+gk
f679rNrZ9cwvWUgXBhOSHzon0hGPcAAbYUUSSCGS2qIyTv6kZq1IHjunELzY
3sMFD8TzbPOaziR0mhkU4cFB/r+UPjvkmeRUe3+5oGKDLt/O2Tu8Vw+znGFl
2Gw+1xxG3yvABDEcW0v1BxEwCwl365vmY6oNyUmih9fd6wmd2AHifySWTrJx
5DY9u4hQ7UBNHT095wE3gpyG/n4OHQeuBtsJ4W4x/QVKo0PqUjkBAvZEryCb
HngENsfUQIsXo+bt3hfxNUFNX4m1LkngvQOELAltNIIM1N1VzJXRnPfx8MRG
YtjQdSMngEgFjuszQWlzr6EtSlobvmvIcr6gnU3js2PT3JL8DAPvHr2wMTkL
xO6hjqZEauchCDnHyMw0JxV8wsaSNTw1nOls1E1Wj8Zu/q4A8fwL4RbQC0de
i9tzMnF8YBaF5yFvAxrjvPjX+xL2hnPVN7KtekFHTvYlIPJBetrrJryyKOZW
j/T3WdidgqB6pde8lHT0HcVUnW2E5XkqJ8SphIZ9oh0Lu5Gpbbq5CEfAPmb2
cZnxyIhUEe1deh56KszW/GC7RawE5Wgcc//Hsc7qGzkzbfSwIWTjMBW6QKFc
Zrz9O/TNx1ZxfWjaB9fbmqawkijXavNy3cVXoceWx+er7NKPxpr9W/aH3U+P
iCTFdthZ9DnSxY9HwOvZp+K2PgwCp0BqU2pNovJBEt8G8R0H9lgIi0sNx001
90qh6OtYs5EQyOXkq9uG9mkRSIQ9H5XHbyZE4oewsIuBTSp35BXQpGiMNTku
3hzIkq483sCyBMopAdCdK0NJidCVchLix8uhC6xCcJ16X6DVZi1lFPyY/1LV
ChxpX46hvwvRa5gqDGx7qpyWRSXiQl4EpSRDkUod9gB2u675RZDUVvBQhWFB
sSOEp1ruEwrocwTfjKEgad5p9QllbL+WNU1w0svGlcU4pGWaBIxR4V4sWIx3
ioStfzMO1blTeW9tTfCZbGXs2bWh3h2wtKls30aIitZh0Zxc59AbOrorcE4v
+9+NchC9oF2OTO4M74hX6SyxL9/SX3Di/u6Z9bT6zdFpRZFc8itvBa1zSr55
xekK4YEvpXQpoHiWCrnx3ihHwWZPPCtkWOyWK2GV9leuf6V9mHwwGX+w16cU
Bznrjzovkc4X5lpJCFgY0mzx7PhjSB/k5MgWODeYlQHOXJVLgU9RHpTqEDmX
mhTNbrzukFElD6hzU4SFYetS0MuTLyGt/+/KOvzMHo49qELj+9KSRlBCnk4w
pZlLZTUyECyme9Tn84K2BckIEUFXhlqkcyVN18jVBkiRhaXu1MEq4Hrp3L3P
thQIQ78Tqs08qR26+nHiRW1Gxf1uxVsJwx1HDXCs0O0PbgDUv6xzP6D+auc3
OV3Hex2mblrUPrbA6hrlltccY0TSVXGTsjgvN0H6NT4XPxbSTga2xG0V0Bgv
DmrEUacHXH07kPAjy5TA5wRr221Yz3GDap19jrNVBQ68gMx54w94MH1WIdLm
JmrDB2pmkDFpO0Ztms7e63uYLfQf9La6Cq2kTyLDekY2vuinqpP2fgpiRQ7k
4oY8xod+17cbR21drZVdJ1k8F6C+Dg3MLxagN43jb+bDe20OxP779PSDxi1e
/6rMA8VeQn4EqF6xDJ5m8IYSRew4HHDR8J5xdNmnhR/suxMtIgxgx2nkSZ9M
HolCTk8VFc5EfuXAp7RoCkr1A2OGFLsEyJ+3H0jTQWgFnuZQ4qgoyj0gtDJ+
NSjStA6XD8pvLNJ6+xZkyNRJlNWN3dn26h7Ip7AmwEsBt2FwLDZpJKvZBAu+
MN7F/oWY7jrgG6HzOIMqiRlSyAYnyZjOL9BtqMg+d08NlZipB8OyWZmtNCno
aY2ss+WCqdwpYaPd3dFDziJE170PhKlwfhjkDYPMjGl81HuRPanoErVH7Gzu
yhJvo2xvRPhoVfi+nv64suqcBZnh2KfPpKxvOY3u9GvMnI+a5S6df+xE2Laq
NBxiD2QkLQ6nsrCyj2Ukshek2k/dNglZL11l6qqmWOKRpxD5sAwV7muNExq2
ZXVmDmx5PkxK3i5VGNQQ2evpGPN9w0IhRQ/0yasw0Q4OUcmNHN7jsjshld1Z
CrclI92JCJ+1Tz6c9B93zD1zC/2iuMBUC3XJccudIpFRpIEu+yEe2fsS5VZn
ZPw6c1e/SGjlad2aMiOKOCcpt8yPVxE91C9WZnNcR7tl6EZH32mBnUHmbSG8
EP2ozRSO05ixLNvogTeEPnd8kJ4akpZ0j9YmkdGXFNST99Pt2AhnnaHCiFsD
OLCHcYTYlm+QLJuyzLYTEUhKI4jh5BNc7nLasw66yJCxY2j9UBmvTwdYB2RL
qRaNcLbRiLT7JMvkI1mXAhUzUH2pSUghVKaHG3hf4WCOFCNcamn9+i0YedVS
BREHICZCFtuhlHWgmV0Cv7BO7AxbmB1yI0WXOWhL5NydedfflwJzGSRuLnzl
BxxlMcx0F9hgaaF6ohn/gAc9Bia/SRtZQfp1+1IKHwz0BbY0MN0pkLuVY5EM
UORE3TLtu4Ymf66Prl7wNmAdxi21Srs3tJBgbci9rPbN3U9F79rTUzv/Gqbk
I0Xzu4xeAJaaRSfF/QqUETPRHVOTX0k5AU6fjZ+XGfu1KM4u8Gh/p6Edz49g
SyArBEPNsnslKZs0O/DXr3kQufhqm1obBQfma42ctqXTOaa+dYr/BZLEKBNi
qg5ELiELqVCkZLdcfkXCCrROY9mNke+zw5giEVQJxNqR46QQAJ0VtTRDgNs2
loyAJp1YdJO3Tu7+Bn7J1OTrHjHrrk+9RIZJL/B9SntUbBgzIZRcb0NkMSaV
iokH6Hl9ONNFFIgW8juumdzBav5eOggzEAcoIseFUzOFeFJKAc19w45Veb6p
5kGiIlJiSjMR/LGcssDbGRM0iOWP4lpHqiYwXXZP0+wuUh8WFd44SI/vOxFN
p9PHRhogubJrsQCe8fCz5oq1Isg1K559SO45Au3bP1aJRXAPqibsSOvJ/ECm
g7SwTSk1XJLUcEKPZ2x0q1ASWSkCwOGnMVfX5aWwLOlBDt/B0aKnMNbY7yY8
CDkZ5Vp0Zq7esFLzg9KVKX7QGjSZ2vN7HjEOXsTq1D0s5PBy/rLRf7Lj4o46
8IIH0QdZbyyP3AKSNSxX87V7NY2XSLM75AWR9I64zYJqhjHLhHg84PCn9kix
OGTBAUei5A9jy96mJxCScFfOQry7GEPoaf8iVtqI+7cEpVPWD53cr2R1VOPZ
j5wV+6m2Z28bY5pYrP/D5+Ja2QRcOrMpuEZslmEOWPlY45Zl71ORHGf4SN0f
wCNTQOaKEvIpC5iKsyxvtS8YHW+WHijq5DL4wRhmh80//CqOI1MoEOqgvXbj
m6MSXZ9M8b04WLdnnqZvYK7xlTlRAyIbKk/kYMIgw3YRDDHgQ66jZRBGBTE+
a+/y8CxOWOQ7p3HxblNNdiQj9ftvLEIWIacEI2p074Cn9T2QKXKXzOulxlta
xNE+0mUP2iLgRr1S1cTR6pDevMb/v8Ji1mmtZpELqFjAduWI7jqNi6te3W49
eBmXvEaCk/gv7LGtDZpXXyXAA0g8aw5+4cM9Lee0I3BiBDZOcUHQU45YrISc
vhlP/zL4Qwnj+rqRXKkBLnoEWxpGx+qTaEbCxFR9/+WGN4rV3PHQ8GKWDhXV
XRav4kE4tgHsKl54GlbTSywFQwG+TSjyNYJ4xug9cHuVtUnz4KtKMcMIbrvX
ZxKaSZjZlUJZrMEFeYR6OldTOa5+7EmMLCnicDfE1huTR/+D8eQANjLIXQZT
5JwS1ATFIbYwrv3YAJCz2TjJ9DI2ucUYVX+GMsAUkNKsLsZwXnFM8pmv0TZm
cfeWShPbCRLkpm3sv4tJZS6e4k3fg/pLiVJkSjxZPRVsqAITlCiJHHbXaPUf
F8DjfYMB7hyQafL5jnhtXPEMr7PlJkCB+eIBfBGw+fIMzE2PYurHgs+8V2xW
mNdNbJnrq5SJGrBCW/tOkI54W8TanOyPEcaZdaX1xv5vzzG7dZSL1+QQVrid
3AiKiKsjkWZWy/S1ry6viOCAxl0FulNeq1wnXZrvRd3qi8qxLbVq2HWn8STE
fL3lWqeo8AuQ0cz8d8xkCLqApKd3mcymc7vsNdtja+YUtNrfCu8E8v5RzBGK
zthEOEAV5eQwjsCOD6Se/6ew3MikBLNvs2DrXbviDyzbk1cbpo3mjtwYZEO3
GguTaB0waCZo1faKYknyLugWg6HyhrvMM8mDJMcW00EiHm3bwM1gWHlEtJ+x
prwP9s8DbFSJTo5bOb+yph6bxj47G2A1BsIo7s0tLTWhegA94nWsHltx6FSj
ogz+kK+YAIg5FpPOS1HdLY+BAs45zCiBIpNcBtAk0oC2zzbgJDd2+bhpm92i
DW47ZpxKR09/elVSsEd4/OHy2ZZe7MVKaIKEC9zhvu9qTFjk68AASdXzUDJe
x/HIQE5pGxJHFYm7IpyAOiOOWfQZsOeT5qcCtRbEVJ9vuvmzgQRtrz7jyKys
NdlEXmpPwXO2AXp/yI9dWnlKM5laLiK1g/8gNr0EvctbCwdsRzk0vzGgUQoh
1qt9DCJzJcLPY0iNE9B3wfmXqZOgvaF0EVjuU7vsPU7X0DT00IqIbnwmtH3T
CiH3GLufCVnFwGGgWO+ewwmoU4dBPZpG2vCf4ssh4tIvQUbxYIl9E10tG+W4
Mzbdk6T0jX/s//IluyMRkkw3++fKRHrpAOs8HA598jBuME9reeze+M0lje28
f0cimd3iHpvsrua2sQBANICsN2UyAKEpOZ3/q4nDrjKJpBNEhIYTiEt6Epa2
nVekmZfjY0QccaW2+Ucp/XUG/A+NilT9681w4h6za6XjyZlwLb494lnSnLSJ
QjajxooqJjUrkEWOhJf8Tl6/nKzyh+SKHUMV4lJN52BJxPKdsWIfvYdt9Ivt
7LAKBlOGFHvZt+cl1/IEo7lO74HC9hDgyK9CLOpYjcoX9fNy1Tv46IfuzVhs
gA7DDDey9WhAEcOs5WLXy66ByH4VLE9Ma7XuDihZt8wyDCsYskSzML2AGOxs
ANKZuWVJ6ZlRsw5Tnhm0Kb6YSJc4NuS/R2rfhKqn2t+dz8XcATM9S0HPuid1
nkILjHsgcIOvaGhgmUIDCXTR9fXwpQVPvYaye1DRqg90EQn702mXBwV0ARiO
GW73igE88n9PcOOmFe8XiT8y97YYxdBfWXi2dbPsISfK/xgNeMHozCXJ/pCO
qHbd/5r75Jrfr0GzWDwbKpC/ACL0ahpKY/QdukP8M+q+PMRDcF7DJt6NMNNm
VCkZU9oXuxQTXfwUdx5576PmrbY7pFufVAMl/8iQNAh2whdy4EqstfDG1ZoH
NWQc95yRV/ie2KJzZbF0Qlm7JXrg6WBlFK0FKJ8igQzoROtDBUGbO8T6QM8i
tcgDrQOIazn42n2uTPCsC4sIwZnuCtipOeznUYuqpxqOmLp4sv7Bczlgi53h
p9Vpmx0a6X0Rn50M72kPIPzVnmDy3nVw299RIQm3S8i21+eGBusnhJOcPY39
V7VCHVjIAVGulwsJjyWHNmqhF9DmFsZ225dAgZIkbEjp8Z3NEWJ6Xtuuu2pN
2bMZxCBwqjTmO08ZGSgNOCBgXhku6Mn8rbS2BhMQ1R0uiB5CcB6Echp6tBDx
v/e74eIHH34ClO3fKHtaNhZqhmxsBTDrBv1XUUQfHhlaWf3dx1ruty+jzzWW
r2NweCDtKgJSEPYHLuL78/BMWq2qQQ9Qxl3AVxs4kvP7mAn6bWhj6Yry86CH
K+bE2Ptl70PgCv/HGCF5HhKYkQy0X2QZ2wpEzFxR8us4xlciIEMWD86BdyKc
nN9SYNZXqgZFdye9GBAqmnB9856S3mdter0Vk/UVSGHiciRO3Aeb0x0WUona
GM1rUqXOoU01Nv7BwEFBNUgnVDCS6HdwacDybXfmBR5Xm6rjnFAe6R7Ufu73
175InyXzBWPJ3Fp1x9suVTJw/gS31AYtCraKhavgMW7E3l/5W7jOY58QQghH
1T+Ms+bYKtgtPdOud/eNL+NQ14Xx8fbF7R9jF7216LcvaMAWrwlj3yegYcuu
MH7oAlRSxN5ZJjRd6OcxmeOCgxhEf2fTWtwB9gCUdwG8HKywLpLwFQci9OYv
/2vUEsWJRULlwDXWqoUC3nFa58DRkaEx3pbzO4BCEa1/KqzmkLkVlzuvEJzY
lUbqw+RKHGWhDkAOB6+x6mbb5c8csriliz9fbaezlw6iV3b2+CV7BLoYZBt4
C3wq8Zo4XA4HptbAvWAkOYnJ4JwTaR24zOob5OC8BzEF+HsKlfW/cT++q82P
PrbbO3Y5sxFydmMMWiHVdnq77v1Ok27WqWxScYowZYcsc13HGzjDZ3j74oNO
MQcA93O9wRJ1geksSBdK8ZWvKO3Ndo1aw5CMBAQypt+cdvobCxALCeNmOTEi
mywMUGCqJYvT1lb3bkSgtk7RQhthWach4g8A6r5xIW8fa8B/0wB8AqPxMbp7
KsIV2ymNAShH+yc1FWDQrQZXPs9qZOqWzE2RenaAJDZSKNk7Xg0/oXPrK4FW
cXDXtiCf1AzDsYM5ki32lYHddxuLLmGSI8EWDjophzpGJynwDX0wB/pbvwV/
1sWusei5SZPiqs47nriTQprMKNIXfF8+kADuY22svwkoHllEE/x+Zr2zGjFG
KJH/MFzPjIEEeO5mJ/XjaRV3bC1jamqzFTJ4+be1ghq3/IIEzWLFaWhOe27v
0J/VPBY2ITEP4oW7qQ4mPlOjj2jwUmMQM8HFhBXn83bq8//62W2Apww8Le0N
Bsu9m4OH4y3FPZhK6dne+KTfPbSdnnpcbeVbON8Ojze++KvFNo9hY9oLDCgu
DYoCA2rnUw0SQn383eUITgvujQlrG4x8GQj83q4Xds2uNkYO+YfD6LY/I/Cv
lKeqEOhMXVn0YbklYOGIaLtK4J+b34r8eN1r2qHvgWWRsOlC+gK7KdJXQ0R+
iW5a7ogi2GvzNhThAGspsJxBDgTjrhxYo4y+286QhTBQwuBgnPmkXdzDob99
nC8+a2Gz8Z/FsJDCkNSB8bkzadWBAAcLRwKT0Lw0NYB9JbgsgcjNh1j8grGP
IJnD2FFLhli5O/uRlt6aP7vioGs72ykxfsvDfUitRvZM7fYJgdU0dVsU+yAa
qbNGrfKiHwMGXaxi916BYDxkoT30Vr0L3wHlBi82wJ263/ZqJEO3apjimzT7
GzaipeutKk1tTu0FqIZM4otO3MaHUykcKVd+iw2qrcR1JaEoE1p7/FUIVSWk
nRCMQ2O+VcldO4bD/NKd46D3Iaoa/Tv7rSDiVbBagla43ccygfWIcJE39xvO
Df8BZgD/s+uKtNDpKG1fppQGP7wNbDrlQwTDWgxaZZeTpj7mje0T171xRx+1
TpxO3Clv9my9qqINKFOFxvHIX6kE1G0F6uJws4tqDsRHm/qTHlGSnDadWXQu
gn+fU5E2gg+O6vv2EQb4OlCA2eBd2IaDEJFprhxahMdecQ3dmulBr7PehPfB
4PGGMbkH2YQltlyK2vQ/pH1HnES6Ljjza0bmKtyCmyGFElu3JhUJ8y+zA6HK
8W2RHyR7kauhxViH+Kddt4C8bkI/J6Lol81PRedWYDhsZdg+prjRdqSETnNn
LLMViQs+kN87Ub+mMXsHSl8JIe7fogmOjG6wis/T6TaHMG2dl1Xa8vl8+18+
1jjYsb0j7dPZZkACitOVYXIPhtB1IkKcqUqiBYj6ydKM48TaCUpymcybFHFw
fwm+xQFHH+DgPojyox3ppf9OW11j36EdqBfa4XPhncECowj2sYQDqv+/q3/B
gmCtE9akQX0h6MPaTRBS0SAgv0JapCwY+XuuioYTGyiRcAJjKVrFzN4bbGaU
mfWgCihOcJofnusRvIo+aE6SJCkEI1r3vUbz/y6BKyYeXJ62eY5Bcbi+9lKy
dei19dm9eYvFsJRHWhifFyHgiQNmNIuUT1vHp0Zd3NqUyfu1qcMjb2XEGNlm
LyBOv5Ugpim1EUFPKi9wZ2V3IWHd7p7/L2UkoZd5fduItMqHjTR1iO8vzAex
RHSQHPhu9Pj4oq3aFWlAhDXjErvJn4XFZ0w+BZOuLjbALFoom1sCVMgRc0p5
baCt7KZLWOSxcN2qIRo9tiq59rPmRwVroaV4hJ857MUsCNhhW4S90C23HY4p
RcW77uf0PWXzdiF/quF8MNPJFjrWYFI7tJG8ECldusU2oluRkTAApFNtTr+G
pz7Do7ejHSZ3e2y5zwtLvFnYvfu384rDtexDwZP/DLIq2+iV0DPAtmhu+rdZ
BR5/+LhRwOi8Huz6hKD5pgvrpuRwzFpyEcjf11DN1gro0p4jZDV34kCTldsp
ELF3MIpJXdy5xo35qpvTt84gORRtOMT1KzO5SyS2WWiQBi5cqdH6CdoJQcaC
hbwk6wqwK3vzlCGGcFzYgjFmnxUw41w8kq9y43+MWika5nPox8AmjLL0jb2/
yFFZwkryN6qeoUXRC19JCqOyhp7iju1+qlnpO+qGZIVkh/ToTMzTKklK5pIF
eiHvcHFbIpPzAhILCbQJrlUv6GpesjyGf2KR7R1zArbp1xyTVn/A8QoFYU/i
XVR0L2UydoiVsd3DSgC8A7WFT0qxfNNiVZVjXVI1JIOMp93TerzLofni3q7Q
5wJSMGYeyV5WsVcK/hFW9vdbprrjqiBPRmndbNL1RJilWbTx8qFLiprPkM5+
hf856E/gOsnpuE8wzykA5GktT40pH871ZKylh249sqw7zv14UCk8InzHmaev
MSDxkEfySSNrzenhws25SXyIEYArXQMpbnJubPHNpO7RkY6NQK4vepOhRuhv
gkmIWzBJZKWTZqs8JWaG4okCl2sxRcKNEN5sv+3JP4EoA098y38zoYQd893V
MlwVY62OTtvUxwUgZnBP1X7acU8RG9DfInwWxy9kOuFhpLUtdlRwPTxme2Ya
6OSY7zjLduj6TADedtnT9yhorBscgVnPGSaqkszEbwvTap9/dGRbs8Loy4kG
OFCYWwdOp4tmCwMEl9SM3U9/d361jZzRciiSxfu3tZiUhTz0e251tZpM5kuD
8UmffbDVykIWcpYdw6K+Aufh9L+5PGH6d8FIJFrvWM9IOOCJsQpdaLGQKTmS
14u4NQuEIc29nDQL+vbATWa+szKFaIb+tv1F8ejBBDwlpSNyHaTJjJih+iYs
J4H7PNcv6DhcMiTWdLvcQe7wXvLQ/xcKyVQO7y/Hpc9U52jG7or/lgAMDLWW
w2DXMd9sKDq/FxpBu7XeGCK9OF2GZf6Dj4RQQyeNcEAElOCfmxb+Xxw19fNT
A9MiFo3HtMGpb69MoqYyy5EfTwPvHZkzg8n5USHwHqUZR9Q8WY9leeiomKCv
e9TqqV3HGHuujmSAl227aHlTh8vGCkjf55Z+zUhTmA88NUzhYeR6cpP3KjHI
FsuhAbC52sTmHN02c9eLDNmo0ZbWs32GCj1i3srDnz7htvmD3E/7+DoTYeUm
k3MXpAFlKNOsux1SHi6jfsxuXHegYTCIN1A4KWD7rvQS9P58GpPtgBbok2qL
gbDt9vI49n61+rL52Xh2HIgmxPXQsexOTVCNPL634+/Yo3H6NSUjb+xOased
nwrK+vtZ967JImnXWzucs2SrEOfeHrko2rBv1eutY2DE3FFibRmTae08MnAl
CW7nOQGcuCnMZf31WaTAQ9AEXU8uEObke6I3BTvkvq52rmM/VJe9ZZs8aeJA
L8kXrVRL8E2DUxlluQ+lCZFWxlnQbiC9WDgiVtSxilCL5XkhYkJuww9lLrIO
LK7Oa9Q/m9yQ2TJ3XvaMe3U3+X+/kXNyG8e8smbSOgNxuYaUlq25wyYawtBf
2jhgyOgGqqtrW794CnDczLIIyp0z6wg3kz1gdBmgYxrBPe+0jd2ButjsHaB3
iQOdd+v1JLJcX5TEivVqha7jbtP6PwP16hmo9UBME3K75OtocION2Iff4jGj
adqNzCWAR+PFwMEX5S+9kxFZQ1Diz6rNQXijDTFWj90GRMCGl7CbWWjIPndd
nxhqv2Q4vBlcPzyGXs2fl2zxggGfRnL6GwhTUEmhrKiL3TQgsyvxV0AvInrZ
jBn+xpz/SgXBnBsQqs/dP+d1va5u86chWkBnpWkRbhCWgoFy7RLiyeXK/Iqe
MFBC7ySso9eTcQ0jguoPaMuq7tPTWv6JzbUmRjxNZwZjuanWzCGDCGe4giej
S193qPVsSKU5KJJLhQRZd08Pqpcyef9MK8geaP2PsqN1JHQvQzCcjCqmPjsJ
Eq26h++9SUpfiTASkvqMAm3BDLRk+02ARlD7GLEyeYfKbPjgJHkScqQx5+/t
7tKxyX4rGltN6ROSZb5bQydo93BdZ/RPfHMqilxzGSzDrEw4ZBAN3YLGiG8i
VRxbfAVtey7mjvQsdgYtIhRekZqngHuZXpVs99fFU+78vQ2J/nEHkiEUhSy7
zagFq+BIHFYFpB8XYT3eu2zj46uVV64Hq9eaCwVEX8M5Isj9uAYVX5zlb4Ag
SV2Zg80EwUPMchA5sIrx2gmAxMRVNwKs7sWOzs5th6xw+raQpahUzK2qGJoA
ZhtiiOfyYj0q2qvfHncKFQFZ+wU5tKEm2w4NdF5IjQaTQ4bafejeY5E3RTjy
KBlpsLPwBiosaDoT2BPzPOaW1bABKofaqd+NntAeDDM7ww6oHaFho+cNhajt
s3u6u932c0kWEvYyvaYYqItX3O+ZYbpdAF+xXlFWgBO2Ugn49oyCVwhKueJE
lbDwuTvTxVyZ1OL+m0fUQRoOvn3m6R26m6qxNamvv5rDkPOxbU5uEvWGfgWw
y5Z15y8P2yuamrlkMOuD+UbKm5jAXcdrJZ0b5qBuJf1o2u4rN+fYqeIlmYek
ns+pPe4N89ZJZNdt3wJPjEK7xix42xJr23RN3pgeX4SPuTkUcGCICuIQJ2db
2hQNOTWYbGYpeh+5LpUyMC2Iu5hPoKSbClbwQMHMNZBtFcJq4y2N17RVq//E
CFvE5Pcx9adTxv6HfIQQ9cV6g5ayrYky7NmKzjOtHanhkjsUJ0d8HDGCpZPR
0D4eccfYIxJ1bK2LIcTdDAF0yYAhhQs0RK32rEG0EkGRuNlqk9ibuoavekWY
Z//iJTzqsgiXa24vtAO4eEgsy2wqaXwedo2jMXxleGT/n3xx/7f5huNwyW9t
Tcj3NRhHJ97I8kpsslVwkMFpeknM2jFP0CR1CadTuZ58EFH0Wfgnq/BvON98
ZmWQkO/i6ZzsUL6DqpBAatANeaFr2EY7ONzbaDxrShzGdqmhMj1AjZ2pgXta
fG7W/09BxEoCpARr3POeT2hquo1M9q8Q+lsA6pq/Jva/8O3old+0S3OB3h6R
ILO2X+IYYziW8LS8O3NPwIQ/obp7dECzzux/zMQXv4cleTVA/BAcwY0wL8Yq
IOYiVSzr4TPXTvMOimpEwnQwmxq2zLwJk4thbQXozp/Fsbm9VwANrm1gdo3J
8vlVC06N9wchSDhaus6Hgizl7jGygx7g9Y84ryTv4DUVllr3V7AznKTKfsia
2JY2UUbH//1SHbyR22P/FrLKHePw23FTlfxuUYs+gdXQvUb52g0PtRZ7kBYY
j0J0M2QXB8GVkXUvFccZu2lZ1CPHGY1h4mNA3FWp788kuGYdpoNyvpJfqtHS
wYQ9rfGD2celgqZNypCx8ud1vPk2tg3bpkaztuwYu7n5lo2Q4EXYWb+0Md6k
cKijLnzlPFj356EgVuafplAYIy5xEmmCL2pcUpMD/4FGy4+Fxb8awrDOnFfr
N3iA62QlgfR53rfhHL1luFGrIFuQYxSDbU/MY3ywh6dYdlvvl3u3/F6R9lIy
zABcaPAhF1geFbOYXhpXtar/W6KwvRlWYa5tESOJseH6jH4xipZHw/jXUZ+q
8syWCTjd5dCF+3jdb19BKtIZ2ZLVaWInZgE19RJpsCgIfIsRreZcL0adIiOv
EVA97JrzpHH3uUztnqZfDjUf747qvwvthlZZdHKtmAIsLTkjj5EJPiyMWQEc
KfRQ+KbOnpzn0rQjdnWUvzGc3Wpc+MJoOqJzKAxcRRZnZBAH7Rd7AvhGWKla
xRw5xwof6um1UM5EMD+o1/vBuq3VzEQYdHVxhKw8V01GEGgCyrg6izuXSBIs
0lPmGW+xHxivKwi4pxk+77stfaO1xyajUzDyyZGCBppI19/0EVz0V6bpVR7x
4ELTl7Dc17vG079uGjGFyMKrePSv4MR+J47SSQ1NxKhUbQB2KhoS6sxonOYH
4COCXrBn9kYdt+R49k3n/rvUoZNXiwTa2lIKPGquQ23erFJZGGhc6ZPonA2m
DSlw3m6ngK/uL/0ZZMZR3jyQE/lvTmtnyEWIuhjWLZNPWFaW+lA4go0oVn1t
Z4L5SK3Sgst9ZyHnzJ2lATzoNoOqWbNx+SOfFA9mfOKMe095yMT7JMJ3XK4m
gsxYZv58BPWdbV1g52hQNJ9qZ5IlzLFnKuWfTVpfW4H26vkWow1NgiE7ER8p
usfrxYHjxLQ2K4zKPFOBRFkS5UY0FMsonsc7T7+Y5g6H0HUdZFKGF/u43o38
WkM4lZmFvMg77W/4wqAR8och/zJcnasHzOBdjtD5H+p8j7bvK7G5zC8YkXWd
twsAyEHfwEXtNgM1ryjSyRqWJP59FP/4rAwlJDtQdhcagIk2AJ50KfubKUB9
s5CdCqz/mpSUjKSthNWeirJOoqMqg+dblc0jZ17CFoYcxHhTRUquHAmDNVDX
d493vhASEknD6eRAhoUXK0PZSYFOu74KylDN3cVJw65nKLsZqTIqDdXv6NaR
DR5A8xYGpj6MUGZ7ug1LmTwxrWsiMxTlPcbbpcNh52D7OTcM/35o1II5PziJ
LL9YsbgT0lsCFWBoIF1x6xRPblJRBd5NwCUPlNvqsjQqkOXi6My/Bilkguhc
1chyrKOPQMjYmzksqCcjWXeU5w9l8vkPngKwdVBTSzv1npOEZ9j9lxULPI9Z
Cf1NYVfIpOLIpDQhYY6STyxGVymOw1kWOldmMv/OLVGp/WGAeWxALHqdWrwE
Zm+lur4y1PKxO/IEYYwN9NrERLdIZ1IS/+eQu3dJB1yZRz9wbOMnevRA+KMk
sCj8e/iNDLM/GzsVXZJwyEQEIRkc7Z/DswzSGqHazI8nc11RSMmNfM1EZA2S
Kxx1spZ9jBn3OcFE6h0vrPVGBlQ+Jm+MlsYsAwZBxX8smg6TRmQcm2uxNi52
66rYaLwP6zojEtynwToFL6DqgKfsqO+IIefwVX5TJSCWWl1jBiH3X/0KVXLJ
lEfy2Cd6GcRwWvEBjXn8wU9q+J1YQkbkqnd9YziD2R91tKUO1a6AHIUr+kyB
rNYPV75d04Wpcg/WwyLc/5jUPoKUDGurP2fJfWncLeoVWs29kLS4rfal+YuD
E3FlWuaAM5ijogGAz1Q/BaxmdnNXGZ3bhU21tEVywQzRIyUbKu6KMe3dM1aI
AvULe+e/fxXhS+gUfQ5pk/NoNtLfucqbISVMF7SXb0ErpeREUMXbYSadCuYz
69aj4K/oTbWJvQG8gtSpptPvypFjPNT1OR3Vt4jMLatL5DJ6csaB8Bbokbgt
UCrEeUyEWdLDzSHrWflJJFVAaDCQAx6Y5DkKmHhixC8CHF69MGY2D6HcgjmY
Kj6li7f+dnck9ooZ7BVFDIn5+5+KpnASSeZffLMoXroH+BfwTmTgEdhqhsjO
Ln682HPEAxGs7wWLYmJFub94Tlh9oezzkeNZ3sdByYKgHqY6GLgz7jc6/5rV
doj2DOe6bqaHLA82T5p5J8rnvUeIH2lqcrQRABlPOUzx/yL36PaVq+lyjlQ1
19WhWMbYaFZx+RGFsQc6Z+01VOtJrUc4Sy3ErXqzb/65shts9kIPljcWzuI/
x620hKmHrxnVPTsjU8O5w3wiT203NlrKwBVzyJnyluSwb05yP7VCJW7vou2o
UwNvGsqKECgtV+69BnA2BjM3bLl/VdijKYLtmWUOmUSJUByzw9BNuzlDScD0
lcd7oh8HsqOg5PmJZPPcDdfRPaD1YMEvVXqhp+A5xHxIQVfSxOm07rwVYlGB
3iMCGo2f5nPUlcJKexVd3vsfnNw4DP4mTGFWtYpx/FXl3dHiIM8GnyVaO2a1
795TXz1mBUE4U1Dr+kAbIFsyNNSPKz4QGoDME0GszUTm9XFk7EfysVUInsgT
iRGBPuUojIuY7t+xUES8De6LZ+48NyMbJ0yN1xQzQHGC63BAkCbvKZn6ReK7
HqNlNOuvR9EZYuGVafTV43oHNKcB0koapWOBmxvCPKMseeLJhM8XwMjQDDt1
NRr6wdnvZMwEc8UMRaWdpm2ABPJOeoB5LntogvDrS/9HY+OIdheeupK2XCbs
6gYUeAsjJx5lKR1NpKHZS9phxY9rsSdGBn+oh6iwrhLE6HGRdVAyEzw1cb47
4VOkkMPn16+fG/PfbkMAqUI7IhCHhvC0mpqcNGsvL1gLiDVNSJvV9UAtrkku
GS4aQj/ThBq492920yXSx+P6UgE4r+CfvLDzIggngdNNY1uGMaJapxUAuh8b
IRE00X11tp6zNlWq/J2UD8P3l1xSGF7etM4eK5kpMolwW0FrmaPlJZPHHENl
2AoVLiO6Sl8pTnuFfw/9jMMDTwozkXNQu4PV8a2l3kx9G4gtLR8O2dNPol2C
ZcsEhk6op3/KQS5n9g+A9nc4Hj/JqZByKH5P6ZY37wu1Pjn2kBhqCrcaITO/
HGz10Z7O2AMmd9io0ANh3TXznpPVUWABPXwXbLgmRV7C8EnoXYN7tdqTAPVr
TvE5RG84s8gg3qbwfAnma64Edcd5z7zIuXHmZaWclLUMKGeYD0iZSrYd7XAH
whPUwCVuT9bUTFXZm2RSNbPRNlsGyYCpFuyp5yDcO7nfaMmz9gZp5xvtsexP
8DbwSEbB17bgW0mRJUkJhuB30UwbKyDsAfuhqlt92pLYTULJ0NpfiUNxHJzn
ihn1f4LMCdWRU3K46i4VMqdYlXET6ntWph+SGP8XVJminImSUSVRUrfiyoYJ
Ob3DgcGdn5r6LiVQgYRbv1xpyp19IRZuMnRTZLS8OUwwxOduQRRmTHZncRX6
BXpIc1gafui374qYRQoUL1awNhzWyjBC+NCtl5dIYPtCYJo83Jei5VcNT0He
lJT8wq30GUs+EROUkIKWOiQK1xgb1HgFQP3tFYmUWPLjVIQZi14vcVKnlOyf
HkYG87tUgu4rqGUPZF89Ib/mChmS02OVQ7V2xT8gIN1Vbl7TTFCJToq3NjuE
wDIiH9C8iTFoyBt7AWGwc5Ro3tkoIzglDI3+McKMMqsR9GTi4SX76bsmfeiu
YoTmZGHr8GVYxJNp69ykX/ueKcgn3mdAi0uwCDOSOhOGkfpCQb57YB+8aMra
sDAYpt+uCXA4p9GDcNe+x9fDdbkpyXhrlkirmd3JjRVf/3KxEbryhcBOZEKs
gh+Hv9p7W83fFdB9I+IW2gb8N0usmQPJo8VwshuaP2PE/m6m7nHPHPMNDQIh
EQD5AlnEsVsYiqR9+o8F0F2csx365AsI1rdHxNJR0clv5j35un3QYcm5KMel
HRJuhn7O2YY7lgAcVGIK5P6AuF9eiojr8AyFpD93wIh2il4wzO15kOd1D/rc
RRQ8KVHZylvY4h/PQmu9EXKqhV3dhwov21tL8BZhWeGLe3jypjcMUKRo4Aqd
8w6Y6iq77KeeVy+yhkFRJ43ZFdW6057TQzycTN1UvuwOGvY/mFGhr0S3Vz4s
T5vTBWkbwjHPCOi7+TcSgj7i5qjB1d8inUalQ6iCxMdXEbQSJD74LPE0rixt
qY6JmTRs9OMydL/Fqbm/xeHiYfek+QapR9kmobf9qO1SCBn/gEKeTsYci/Od
vWafzMXAMf9bh3aaPZO6YPKR03Xlsj4qiE90QvceadG/KffISnOT6p7XevEq
VZ1iuEpUDO3rkVCyP+bWQjIZzQ1l8ORN3uoDoHoOJAFhfJSK6LjqP/9vB+F8
TvE01FitEeG/AIfzoctyrryQ6OqYCQ658JdB/WuuX//71sXCbTq2FHoR7td4
a8Nk0d5/3ajiTnYXy6Ay+MnxKYmTyfVBra0Rcq9iIMQrWQGYicWwajMYhJlO
DNQqnEYRQYNv4djJAzSWW4ZFN0SaXJzaG1KdfxqcWZ3chIKESABh+Zqj4Zg1
8FK1L+D9Hd0GPpBD972+RAKaT6xL3dxQNtcydrEJHkvsMhM3dCABNWHJFWDk
QMRkWMt/s+vqvreudP0RSuWlsluvkz4hj7pKdtWvZeYAaiY7USGd98WAgYSc
/+5SYvV3uhri3fayYe4B8LOiMT0acBYopx3MQvIjOCJ1O83Tbh+HWePJQfAo
zRcIfnxoSJmT+5aT7TppzboQcAMiHFf83sHPjqUy/gsHBPqT0yeK1keSwqnc
No2dlU2NXuQLJV4dz5jfDGu6GH4bdJB9WqtDYqu/U9IQuIUUgi1rOeYDJmIf
/6DahL28bfuIBeT6vAY5GeCqrgCS1uBZRJIMKHRkPpncWZyu+q9x8Y56oCgj
tUAPsgrOqelOW5XGAKFjafk/ey8r2we8PUIuCHJ9yo75nyR9bIqkJGVQHiqN
Xoq9Q0VqwqWrslynj9XlF3FCkdGDygSwW1UjfzB0VKq9EG14QUNUWmgRw9TU
wjpU+spUidFCJeeKd5uk0hdHG8aYdQJ1JyNcqbtBIm3p+W0AcG7Juc331XTn
8d+K4JJj2iTjES3jBkqgoWp7hIZlp58Nt3oQE4KCWsC4McMcXWAWkn96JxM5
8q4JMMIrfEaCqNWjBlXqTuY/Med8pKJm4WfirAx4ok9ygBdA6VffQhaMoQNj
yL4qLtEuCn46TFNo5ifruTE1s43hPXO1SFBr/SPqmah5n9ex07FsAdGD1MCe
mRWzffNdLqlMjLl4VlnClzzcqtX7/OihQM5o1/HsvF8Fqvad8bPJ+KJ3Rqj8
luHz264dHh9QfQowMVYs2dMrgi5aniMhujfhjO/kYthriBYXMmQmvMnFbYe/
Rhh17F5ixoVnCeeevKoXtOdWxbUKBm+/R/QJWxTKZhuNVd3OQT1qE7tpayJh
/Ylwg2GjtoTjmPz95DnKPVIIIBhqScs5dJgXA3W4MnznlcuAtVDC57nROLvO
15ULPnwmFPOe3CCscrRyrVQzNHdS68Mfe1Xfo0BtRH4JTkNhpZ+n/O0lUxk7
qY44sr0IkiM1qV3sBm0Sm8lRKjvHttSOUZHT7616k5ackQn4AstA3kBIphLX
tq78sR88BiDbcSn3feAgMVlHhO3dLkGzG4PvCvLyftFYvagPKk3WlDoMT44x
tTHxVIL7nNVAzWb/OFCw3npuZ1klrjEIDg6GZbQVINlQYxXf+j3Ols5Nr/3S
MRJ2x9T3DsKaVDKMulBG/XK2W2kp1nmIROSnnyEdt6D4RjFez/5IuvWnAnkU
kOawsPr+iPOcN9/haKfKw3RG2DXgLCVFDTPjVScjZXTqEum9JTb1OvgC77L0
0hQIhEClZFJ2yzz2ClDY4GPgiMJouC8Tm24tBT44zutq16mlkcjDTCnhhaZ0
JcVZFWk/rZOh8tlItlOQ9PgIrPlKlQIWE/hHrPXSzEZi8vR8NQXLHskUQGIC
mDbV1slRKpz/Jp3Ga9VAnZWVWp3Bx4Y0AFLI4aXVYQiEYa0u7ZcP/l5mlWqW
0mUp2FiPr0tUym4vhYApBoe9oi5chbhhNG9sSXQEmbbxa39ndeOo2txoD6GF
sbOuT5nOs5cE+X9P+PeujdDNu+W4ca2uMomKgm2g6+1geBodz6puzJblOnD5
2CGZhgbBPQLLtxFnvEodTNEimqvz3AKGmLdu2fl+uLWDXdrQWSM4cQsrYLIW
maZR1OGH1iSyQnqFoABaIB9YBN8I5cLxdiJF8/VPkm05k38dBFsYFfYA+OjO
Q4JOYcZYk+XpOh3ELWc36cxWuLG5tOsBHfu8FTBAjioJNvJighcFgQOVfoCF
2UuRZhwHf1oOwhVIgdDTLsOVJk6/X4bLWMRFWN73j0jsMlLNkpF8/n48Yfo/
us+X+Hv9MyKSb3oTp2UiiudXgtwgXmgZN+B/aFVV3EUbJB6jvbJeVS6BdyKj
XHbtjIJNkjXZpFbiKC4wPqAEPVksHoktEp9SJT3SSn9p6yGNWL8BVfCsdITa
PA8Apjnp0rnkLJpXsiHUtxj8UfcwAgPk/avwvz1JZS0IMbJw10EutGeWkPNu
ScpESMDqs+R613xlF9Ri2Ql60Z167O3L3EtnB0eu49SDL3rTf8uFbQBnsxGK
Qk4rHoJDp0CcHZ+Nl61Jt1Mu/uYqbHFmcGe1LBfsLNjhqtIr1JDcjhQUjkk7
3z0sNk7nq9E4ewobhSbGSe1yMIpO6W1SvY0qrQd94miO3fnNmny22jaJLPme
RyvhsgK14Yoxc/LcOr0TamiwL7WqgDZoCy3R+naI4C2cVdYkcxGakBOQohmL
ENQDEv/FnOwuoaKoLdAfED0Lthn1gUhz68WZeWMUFEA0B/U7UxjaaKEFT87y
Y+WlEsJQsx+VijB3LBnkYAyZxiZuBdzMPbv6GqDHUb1J7v75xrUdM2c9NKGq
R4vtU5vTiDTmVPB1B7mr6q1TEoaPTyIh5Uo34XtdGtiuST84ZIo1EnjEUtyP
23hX4WHkhgAB6vKZruZ91S6oTZaxnqTGeA1UrLNeMNQP+Qv/0lIqAUoIYDxh
86UGh2/E5hys21wZW+h/ViNlaENKtAMGK5LUOj1n8BbiyoxeoF7iIculhWF0
0maz2D4IRKlW7HUx0TbhAveWCw4swVQQiIwQWprTZObRUcN1XPM2k9vDf9yW
BRq4q+f/zMO/K/+WA581kf+AleTNPbklfQY8oz+x9A3JNxpF0BZXf1a+pjXn
JTHN6kdjMpeslyB/ORLDeRhBB4iPrJXaKEj47ru6xxTGCWeVfhEPts6S51kl
F6X/O0OEcfmiJGROIwpp8hLB1p5slprKz5FwXatxWIS50zst7EQtVTDDWUGD
SstR9GN1YFcA/coJtp9jY4pvrKzCjJtZfddpD3DCGHOWyH4Jygm/X8fE7EKN
TG8+ngaphuokIBlBz6NNjmrX4QmKRUUsiD81bNKA0vAG3LLqvDrpgXYgB2jw
E3jLDD6aRX3qE54Lcqy2rsrvnPxyU9H5AnJb2fsn+oJ8qRgg+st7HfZyjGOR
dUWj/tglvFDSlUNe/xfacX7MzXGUAiO1Kw2YwpA/I6k+d5QQkjFKUq3U4E3G
OTEe+pm55I6VnkfFRucwPsld10XpV5HI3Zeyj/DkmD0g1JLPJmJ1EV6dQVFG
2psbpthyw77moxf5hRGD5V2MHEJmmHht/kmyKoLH2v21jh3cFDKU3W6/rtwk
mTJG2yBsz57e63ARzqZ3zX/IOObPud3MWPIAjCKYzPl4Nd4BO4cmVQiVqRqw
oa8yBxUUkvCxkR27GorxVGVgJ9ANYTk41QSyOYSCAoZQgnKUMdI2fGiX+147
ToVVtU5hCccYs9PfXTqz22WjYihqvqoQ8bLlLTS6H7Vi0KrX2EaYb8PTwfH9
lGL0inIb3proCaRGHVi/3gG+4lxQqcwY7OwhshpGSs0wvKPLx+by61k4nM3s
fCXbLvXa2XYVDNyBGh40hufYH4YMvKyHBKdnKjHuTGEKbtOqg8Da/o+BTCfj
QMZkQ9KM7zGWrj1+OyMW1kDBJgEgaNB6QvT/53WIX2t+qcT4e7Frji/0MW39
ApPkCtTHQ1+4THB9EPU5cgL2xA0r9aPm+l30Ot59pMJAWCVUgJ4hddvkVwXt
WTB3NPhxiLk2p//2B28/eVJx0Ojcxpid7V/5amvscZfEqT/dzhNwVa4hzOEy
uaeb9lVoTrCMcz5LT9HHVuLxQTPb/1AjTS1QwCD85h+BerbM3EhUcWQktqsS
sSqmq2guM5dgk+T8z3ZOy01D6ouHKWy/BTBJARtw/zIrcHa3MvAblt0AEbFs
ZwddPv5DEbHESkqIC6DGRKmWDNa+JwwfOitXyrr0DQ7o5e4t+tFPpZLgdCZe
JK3z6JnYnmvLQmmbWMNdZeWkR9fx7cUVu/tvEHAFn/zWjSQOKjmkeBzTN8rf
qF0Tt2qEbf+MdUeSzZZiNEP8C/JdgwQljdxQrLa4hnoVt1g9Wf+el4tXZ/gX
DxMN4mCJZWT5PpNa7Cm7EUlZrVMsyTX1pk1E3GsObJCuosSOpFdRhIW3+5BY
qOklR+qt4ubjXyP3SSIP2PTZZgsxXEw5LLBGSJdBpFQpCmBzMFn15NVAGxPh
gSM3tRQNGJ/+4hn28MgNlxqeb+leW90e7Uv1G8zWaHSYhDBn8Zo5G5SWSykM
WXru4cSqSkjja0XMmTJobMD21KsDb2y5+9Xu7tLQhdBXVAyb/KxaZkXzZl5t
8kkUZxEJOSsdY19gfP/txpXZJdytPhm5wY0oToe65CLS6ApVRTwwJ9d/yRa5
QM19LCOl/+Qdm3XAt66BCiZM8joz/8S6uHOuIDtDXggYpHXeg6Z10ey1jRzr
NrdF5nnIoFFlAG6eMLXP9iwQN1n3cPNeQtGP5mYJEC/6cpEAhtrLHlNj/HzG
ePYUPTslljR0Vta7I7OXlutiEO6wQGJklrlCHUifpafLdh7G5ULL2mLCe+k8
ie/RBNCpNAdO9SSxKahW63CNFoRboAsefm9RtDaatrcsrnPJ+PevwV89xUAV
AFEdh4kc6EqXxKm6at93CZPoMqstqeGSgVjpWEBAQSXcWLfpi04A6g6OtIjt
T5EOAVvHqvMW3Y4nlBJIpxwa0w2azSn86OwbIQtTkwiCu/cyCthFosZK45BN
aLroK438sphi06oarektoJorYhrcIQyIOMYWEQU78H+bLNiUvtMD7dB36Dul
9K3TR97dW+ePlnk6cWE7nA7TbQV/3EFegpcbMELi+5ztY3BVxhE6tr6RVZu0
5zgAU0fOJ9epEgJrHwrSUFQ7rUrlDfd2RqsAt10axpay/DDiLtQeMzKAS6DT
8utRdyUoz6Q/hs0hCk5sIOdCeKMLWj8CI3qsW51vLxltCmHnSb9UQvknOxRK
JF8c907lIEH+zqYWLSUlpBtdzrg09yrwI8ZX0A+QZ+VOJSwwD0i7rxhaVVTN
ck7CPBVQY8dpnbLvOCi5pgeTrJXfzj+F/vdz0ArptrdZpbrBinwHaLOH8JT4
zbTusQGwxswxPWoe6XXSfiHvkL/3tZ+YrItZbTmE3ACoOq7oQiKU9jLHKTcN
WmiMFXu1ulHZ+lD2Ikb/ubpSRBCsnDT4nPS6Wxtfj1J9s5uw51hQ5B8BbgvF
DLftpgdUpGcLqjtzcAZ26ZI3VnxvwE1uar/JenWFzKb6ua354k7KS1r4zcC8
RLhki3mS+hCTXxihYpHPq9oyvp6UcQASjPNGVjqtHmHlYUwkB2lqz7BipzNl
XYQDb/0qeD4oKD4Egw6eeNwyckMjO5kl+F2rqF+W3E7Yi6t8rQfLW47iOdxH
ScON4aDr0BbK/SUvXykPj8I8IDlAGN68KE+utRzYWJ0UUg1gG9glj0z9G3Fi
rCBOIrQ5+6kefgEuDlteZDKqt9sCPJH+7tndAajBzJXd8EqPwUPnGUX1jQAK
leA8DQeqDxTh3CR2ySFSm5epDn+DE+xvEK8opK6GHVYlevffjwIpS+UosYEX
LD+lusEMqbTZg2VLSogSxpJyvuq0ceWxx5elbOqB5prbhstmVoCea8alk6tJ
pJ5FlYCOwTXi368sPczPfFy7irxVawTlu3qwAdX2PWT/N9DLVGOfFQF4Rewo
9KTvLvC9oJ1LLpYiPPs/DnU5iqt4ikkJTc9E0Fa2vgfs2cbi/qBf07BYAzkt
9hGOfMcze4yd7l33OcYdkQ02DNztX0YXzNLiFxBI8fCM9fpFpRsy1edO32NT
9UDW8UhqTra8Wog2e7fI3DAebnqmO9skvegLtFef+BMTrbqm5CUaUINriEeN
yFaNSnoWpwHmuA0BJKUb2JZe50WectOp3EaZR0rUSUeI2ctQTGSP7TpQSuI7
eqgNayAqzkMpxp+yTKqfFZ+GgC086nz6Y6lHFoyL8KV3eNXp+UwKVBeh4q4x
tdUxSJRNrKtfijcZTkmeWjPoN2eqd4mplqGL1tUREbMFyAvnepU2mxZ8Rx8H
jAk2BGrur4kPv/lGfBEvFnwPggr9n6EHwI1I7AzUSEB4NvrH5kxSFjOJ+jFB
eT74t0Dl+k16vBOTzK/o+wNzwRYYt3YsKpT5bwdW1LXCSuSPBu9izqvOTFmC
duwXzvuKdQhuDTLh9v7TMKdjZ+shOjw5bZnVSiOOt+RMYcIiV2aY6YuqTpJ3
Q+gexFMlkdLhnOtTLJqg9QdtVSS0dXduyjnb6PBCKdrVjkR2aqYmSySfgxX8
Sk8NpBCAqZ8AW5hkdw2ooJ8Zv70SVlJMvh2ClYvFFaxV4B/kpdrp+8mMQDZ5
jpAY/W4CkLXtocO7Qq/pAoJswwl8X+8By/dkxpyx5Zx450PCGp5b+cps8rEL
nKn4xVhhNk586p/tdib+ReYDygQ9+MluiDKmBYhqGnVS7f/EOoUmshrxEhqQ
7/kVAbagUati9BW9PrFCdXaJFHEV//7TspgrOxpjHNqVdy4bL9jOIduYHPWA
D0BFc+iMf3BYLA6xhh14t6QZFoFSXxoYXNAN10zO61/RaGi6gJ8afAhpI3tX
qrGxYIU/8GP/Q2W3tCvPYT/eIArFaGrJ3DCt60NykSeVHoFPpSdWfYyCh+h9
+J69GKSDoyZo3/s81wMAABdSXTzMAyMEyjLLKwGcxh3jBQoiXAsPxGei35uL
Gi1FsKXCxslOKY1PJk5oiDxzCTy0iPm/I6obtx9ANjYFUQuA3CI53tF+r6Fc
t2tGqzzL/YHNxstPJ+01Xa+yq9BYJGvoJlmC8cxWAmWx+DzBJSqENZ1wGwRs
yYKK7KJxSxMMQdXMV/1EcIQgiuEdc53rLjAyxhPgeZPMN8tC2QJ5qImVGplc
1+0bz0Wzd3c7infoa3XYvljToN0SrJVirNFQ9/t2JyY6enMapvdw2l+2Dkq9
bDBIC5MwbihOc9Fbt/gzyfzx+RJh8Lkw9IwMXOLJOJc9e0c3H8zTTp81vUQ9
52xG2j4ZG/SOsJiNjVFtwGYZjUgpCK6FCCIwRA8tcCi7C6Nd116gVn6RvZpZ
A/jlsKxLgy+kE0ZN0N8mwFxvkz7JLBjktiKhlmaiziVJBZA+6iir/c2FVfd4
wgIJ2nj2KEnLi0e1DAjE/n9kmraWyfnXqYdQwfvNLCH3wXRZeR64MnEef/Tf
56+C3Zemixc5eF/Pws9H1bAeKmoH5G2JpkZOINq9uj/UNGCIyNBa8XOnHXUk
DK8tip5Ked4e488qeQLBAMsYnBwa9SRpJ4z7h1ADIFWVdt0Khuga/t1STo/z
/M4JriipWMEOz9LNsnKArx1RrKNxErzk9DVNZjsDZboVk9+dtYDiHcQW7bhn
Y8c/Q/j6UoVVh36LP6yTJasau4/u57G/uQeD87oT5nIyO0JsILsUCgimAFN7
LN6ZwkbFLEPsSXDDhO6LSphAlp/Re28T1Vng8ZL22X2qbqVIhIVht2E5vjM7
Bl9anW5HlSAFenHKotjRSmqzW09lC2U7qSvawCxiFk50Xn7cY4jMNlNm13tO
gwmI3Kox5dpkuQYb1F/3dT5VMoMMCu6wcRkKHKjdBuvdHSh4DAyzzyXDXBA8
rA+Z6noiDFqnDy8ddysSrZHADYgRQiMpckB/7g6HSd+ifMP1vaCajafARxoi
M4kC8NSSfNUGImBJPvQgQFXdwcYIVCVTjCU0TJ9kIpD5QW8uIdYqUTIBnl0b
Du4ZfjQKDaUTYx9GOb9/ih2xPn2/iATXeCDobYn0uRD77RsZylZgbpuPC0uX
bWF9lb7Q4hMQ9URiIOXG6Dk2LEqfU3rFTv02ZzZ6YPyrBinh1j9FEVmf/miE
DztunpS1xjZvGH4jW3UYTkw4A1lrdoRiV3YMiDBYZ5s8ilHrnKRgfvtYnO6Z
N8MaQz4OX18anYnQy5FahotEdZK3CGBR3b0RVolCRCulU9Jpi4RurZGauMHN
ZrFZ+/u7IB4FD0ajLtR03qWW8POKvlzqbtv7yhYLnBHGyL07eNrMP/+226Un
yBfOSqZmGaxnGuUajke151u2/aNrOUkb1HCpQQedFr0cS9RbrYvbCjQfcmlh
CDqTORWrzG3MmGAEqmt4qE56vMpPIUZL01WbBBlqGis/YWVO3Ef8mrmwFjQg
DArPqjsFPW7OmjKobK56PmQMSeMUPaQr5hIZTkmeV6EiSVQSo8ctMKl2zoeg
xxhzV0KfoLyIAOqv4w0Yl6M+4jfAjY7vmZj+wCYeh8A5lWAJ7+x5kaVl7Ewi
YFNBUabJlIAbmSEuaKG5vSKOfbVlC2Zvmy7kdzTqNLL3Zq2XJnSuSkrah+Pm
WHjcKwQLa/rn8S7E7HWLMT3zWTVex8Vp71hi3l+/FEGyeOJiWDGPpFpoKfFQ
xEZ3wsRC25GZIB0ZrZucdEwbGQJM7sSn3UXMxfUB0CDI8evOFJZ4q1uUU77r
XHLlwoLvbITr/kftRLwSScts2sQ+OaUJHoZ3LK26q/cAnEzw992pOgyZr9Bn
AtvqvKt55uWJn7E9MeiF0CV3O8cdjNiobWQwXFQR2EvhrggZshxnl/vEDQ4a
U5W4U/sTvxfuUapNVA+ZhQzanXnd7TYK6AHN4CAyhBOqcdhYgeX1hqqd09CQ
/x36LvVbvw95c1Xplt1RKNW3KKHvo1HILuWNNRJVCSJbNAXioDX81zkkYViH
7a7FgsAQrgkV4slA08hA27aqhbsq8AUP9oe03/n9C6aIzVFSbdS0f6Zwmeth
pYtw3A6Kyf7PCYw85Ey9FLpbljkRu28QuS9HovmEye9T6G9vxI1FAJYBS+e9
g770fXX6XOLdLgFcj+wOAdZ4TUUH2AtSM0MhQJEo0FEXA8YOHwoFuO1bAgKs
3t79A0U/KrWCuFNcrOwHa79sm0QjCaKc97pF8o9uwD9LmAqIZ41/33pJUumP
HkHDQUHUvikvPwblcSy7rErVEMarOvsi/Bgw4I8QyoqH/UlUPfaY0r0zwywu
73v5khlSY0UMEk/0jT2mYvs77z0nrVPj1tp+MxijGxVnTN5OUsQ8y5gmDojY
CaKrKtUR3eCpYtwii2FYFRHg/e5n3Bxc3CaSyjcVMI/zn+O4barxPFu/ThjR
O4ROdXbJgA7WhIVsnbesAdl6yf1q24pClznCllV/rkr7NSFaSyfhwg9mpYul
BE4uuX5b3T6eNvlaPbh9C0umRO2wgRnTcwUBVQ4sbEbDLtWFLQZKRou6m97i
e0eLUrjhscYAlJCk4PEAL79welQFYjqW4QrpsY+jN8n80kns4+QkVl40DiUy
4bPKQaWjfju4bPvU20EBU5T78diImuXg+v06XazcWzwSNJanQtIKzebuAcpw
5jw/xeqI4GlfELSjt6h16c+znlHbWVOIbD1ZMqs7jpWgqHxdKejYgB3ypL7I
A1IdvCwV63gQ6oXsRIctXGLlzrIpr6ZbgG1mwVVwZm5fQfBQVdg1zAkhaBcf
r7O8hw3RmPxZHDvo2CFAxLhGtET7XQfddPykbShC3vdctsOxhVzXBJyIZSDT
HpCP+3Uyw4PT4earemWJzpgHLwnjSkGxRtbUXni716mVDJ64ORmOiRFuJOVc
Xh8h/Hw7mRVAB6TuRXHEgG9AKJmiBu01aAbppnyyFhLIVOgBkPTFkuuegkFi
S5pFUXSJFa9AHSwzp073zzSNznkY5E04vPfl+0mXalzfCKvyOj9ckqbSOTdd
gOYT6jQFstaLo010TsT4LjeGBBGW2CLMm8O6D67sybpgY2D9HsAzMJ3HgyBO
5i2m/35fAgJKjZdQYmYp9/kFXPta9R9R7t6Gp8hzqxQJSJZmeKftZ/nEUndQ
n5ZZbIhRdu6ehNtCo6tQisuWgKadELafIYtfN7Di4mbkYs8wDuYQ/aFxcP4a
njwOI9xB5euLAhyOnja+p8drD12OlaxOhk1NuRdLbFx8dUn09l8YNcP3sfb9
g0bS9aIAth9XOmRgUTj10vRNfE8ARHlOCsOz4Uj3zNqaDRGXtDumQG+JjWzt
t1Yc1vApVmRaYh7a6s26lhHrkrSq3Yh8Wl48jMUmC+8hja5mBkg8EjEtUsTt
kEvGMNzzfByHJQFikT8I1/54jVBMJsW6mxmH76ca5IL7rLuQFXUDlsp83XrM
3htYiz3pstREXCBHC7zbYYAfutDE/z8QJ5nv2bxEt05DUfiVUAzuSrMiUSNy
P40QYWYF9kfkRmdQTU2onJYee9l/03gNVUYXJQyYmoCPDhG/ZvFQI/n25Jxe
XyZYrIq5IE9AFgM03NhQ1tc/eGa2gETLj3fu46ZMUTz7DzP1d2sOO5LEC4Ql
fKyTbb0MyXJzXsTXhWZ0twU+BC9qXlGmC1fD3iCi4sp7rRrrNDYo5jYbmCdK
UVrXPOp5gsIKOJrzyd47laaWRiJzRnyVDcFMmRqWtdpGfPr/VBiiPmZ1WIwF
TM+kuV1iTiCB6gtvykBnzJSiBvx+9+h3wG11DYf1XdCKjMD8MPXevu1sOw7j
31eBhrAaKVZ4kiTdTBLBC6M39G2NmtxCDHyCGGiwT3Npwse96ivASITgqsP4
YTdnqRn2UcF3E57a195paNx8J/rwIcdA2jjVjFBcpQEOpst/5sJWvoaxany0
pX1W1gV6/wP4v/YU5+SH3xvYHb+7yn53ejqbVPTjrp5eV338zdkm7U2R5GY8
+GlIf6pcWChuvP7gukuwTr8FZPHOVMOO0OL5gKqX1+YflocneAu+PNbdYQ0I
mgPnAi4JEpCnzgjZpHzbaColVg2Vlz1Zp+rTtEWxcf0OszwvsvPco4jQHekV
SNxbcWJWCJ5jGDmJNaO2wp42ubW6w4kFD3Wy0DEv66yN7pWoJxcprXyJ1jZ+
kN7QSBu6euFimU0SsNlptqmy1AaNkYwe+KNlT1nCTLiQZIg/SEK86jj+OE63
pKlpRDKtgtha0zNV9uwQyCKj8XD9BY8iey8xGrM+xj7Yr9o3Y+A1oaoO2kou
4k3uonlyhx+uqulNQTTSLBuvKYBwqLv49YMcwp4G+hlqiZI412vmO5JYbN41
qDtejH65p2m+e+y89r6OZM1Aa+oIuV/eqz139rgTDeeqsqPoi3yGr9ydhhfJ
2P3hxdlUmpdNA53mJtLv38HmYDarbIaF89XMDYTbrHrTcGXbKssmMyaD8ZlZ
uh9bLZf1yQogrbHPmPp/hbWA3leZLqHvqY2AOKa6AWgQM2pq4ZNc7svFbzRZ
kQf804NPzDKObjC1TzRyOze0GgW0jkOB/GjoYlBhp5gu3AWF1W5ra1K9yvA6
ee1PBKYodYaG3IRX1GFbinYlv3s/jjkS+N1FgtZWBGhfXD7nvftw5l3IxlOK
AAXiI+KBLXadrH4TTk6wHYvUVitHlMhGOkeUI9SNDKq7DWXIXUw0jMRdCRFa
8mrpsKjSkVxGzW0lQi918OROjZVfgCKfWT7jhc/HcoK0mMbqU/5nGXh+irlu
yRJTVrMA+WpxjTmaD8tucPOZrIkZ5gAOkRTvuzfQGnFU3GjNv7GMt27WC/CR
iG5PKlRGtBErYe6pKkuVSAw7XKJ+oyLcPjAEUR/hcJ5kUCtw0zFjBgUN1iPZ
wmmgtJl7ibHkxoizvdzpxTWjNGOD6xnED13xq4dD5MarhZ80kKXb1eIPIiLV
e6Q8tNhv5VvyGOigTMDeH8xxovLbbm6NEBjRdbhH2Vkt2Ru+werH1kp1xpUz
Tb1n29w8gXCLAWazTpXXuUvYvILhhLj3/9C4GxFfLxsqX+CZsmQeDSjcJzV6
GJR3Xnh8zT1mqaOmMGUTdUeRZYcH/fDPLTI3AxPsN8b+hncj1HIxfiHrDp50
GyKe+Ll99miRrwcJng2GkwGoZZpVCxnfsSbNp/q0izCRuvS/PaVL9sg18H6r
kNtYOyNDdshAQ8DTTE5lpL0a738pFRC1kOTbya+Dnb60tEMQBHVTrWL5x56L
JICnSeDJw/zy7sGYR9jZVo00s6lQr1Xqj1m3jjvEEhjmnu9o/Tcl+4kZAbFc
LPUqbB90VOzT8kjPHHbuCC+nDu+XMj8u/TUWAwSuCwASiuaKosvmaqOURhr2
KKbX72qje4QPF/Z0kvD2ojaSiQkdutjfSKpuIipToDeGm2u0f3NZDOUhzmt8
OiZwIkHoN58r9Fjuy0I4rPblfXKwp8OwoF9hlSvLXbZFP6BZBVfuEK80yMsX
KjOrcJ66rankK72u04Su9+m2vkEO1LMA2bMZzTR8Mf6IUcnaoMBI62XQsdDw
MZPSwh9PQHkTsuUJQaD9sR1AkWpYAUxM7lPS/HQX1Zp5Dm9SYR1zKcOBaPJP
iZFPjXUVtYWRCxvlTg6p7haZzUBBtqEO8ybonWUSZ+FyIT8qJ/6ZOA0T8GS1
uPsQYtSddrg4dd0mxyXHLQEmsfjBb4wQxSgHYuA8fUYYH62eSHwB3g7AX98v
naNjND3CdyAFCrI2onJNkFIJn0Ql9hd1LF5BPfBg+1vRTU5RvkE3OIswRn3C
3LD+cHldqiq+zRxznNgqyefzC0fBMfeT49S9N+Utbr/mFdE23bYR9KjmGYBe
/3Q3VS8LHBMoHlB+lPs0/hbnzfOO+ifiQJuwnG1okZioDBuCMoecgw7k0+MB
zrN6Dcd3dAmpEkfAlGRzeu6WFjhdBsft1VReQHzZI99WZsHE3Ti8zJersIBM
8FIFLzIRjY/USF00rjFL3ZsVtwkK+zv26QiMJMiu5dYMO3SImjw2kTSj/SSj
PQdB+XKr+HlWxXBS8+6YOdMHKrljs16QOYBiqqUIPz8WOKdFBO0evcuXNlN+
m5QSCxW4I7+i3rgWfInWBgXJK1VxJZq/HQ4R2h0OsVnGvWI3z+je/nfoxWqv
McF/XZd+qEwFjNvjrCBrj2v63vSTVOVqYDgryG9FQ74mFctaXrvlw+CNmUVX
/HQQanR1aVMOUH3ziScSnDdnxjteWFja0mTt5zsDdEk6f2ZEzXABpOJi5HgV
7dhpabA5fOSQl/ucBPYXyBYRmjLG20RPG8PorZZxj1X8tGQDzdoET8q5zSy8
WfvOjoH+8wBvC9b1A4xo6NZ+n6fIBYJ1wY/5fzuABJwBFwkVW7HaKiLOV5aS
9RMUrkUXPEipfRfda33BORzityq6ILkl6Eo+pTxwNhZejEwRa4Kg6fgYVIyO
vdThN7FPhCZnq8NcKyj7ddV+/O153wlwiHjqtfm4bbhV2Z7joMzru1nES2P8
WsQJWu2zbO4UxdFWLhwx+NrhHGJJ1ngqdTVfdlgnCaStawFvwU3H3wMkp9wT
vzeCqeEH52KFBTvVt6xOlR/1yQzhKAQEjRK9mVQ26cRZHFgJO/toTxkJa5hl
cvgxtgyia3eaakncjUfviwKviFtxW1ocowzIk5uZKiYB9dbFER7AqFY/g1CP
RrI1aeYoRz/j2Na/GRvx9lxbmV+8RJDkQTAxHBCxXA2zg7EGxKqfXZYXnJQT
bOiyS59x8YplOj8irZ9608O4bMHUUs8rO62kuFip2+NuYDCOhqoVogDY6uvt
qLsSyDvpb2JT682T5ndnkdB/v2syZIn+BRdDjIvmhchnE4MzeN6NZLJVaVyt
qwccW0suVJAYvANTgNcy6pX3rjeMM7kS5aQ50BEdpz98Cb5xeM+tYHK9pu8+
a4ZY+zFZgcBV7Vo0Jg402h3dlJgXt3JVeFv9uYJBWoJ38g/dxfRrhJ4hEpvb
LDU21Bpd7a3gUDyJ7Nhn2SHlofH+nj+LErXjzgUv6OftCb+w7RTWSCYG9EK+
ciXwNtEV289L6bZHuf8wqJg/KDS4kFc6wc0eMNYV1mFGbLbDDEK6ad2xP9aI
VgF+czkvxwudsMtHDuR4S6iMdvnVaIResLxw5LLVxuOLmhXI21XGzPZoxduy
QXPgRufzGStYNIw4yUFJ/KDhN1yPasp7RxLvYW7vSqc9RjEIVBzfjj0E+UG3
/AePEzX3Pa+J/3oqoyB0VsV0W5omCSlkSLSRCL/eZ0oeZeHzkALEbdItq2Vs
aYtQNyOD/UHNkwRuJkTx7sZF7/nEjqSrRDvgFc/VIorA2OHooznPGSCJ/HS+
ETZ8tqREaF4Ps1SarXC33Tg45mGygEpb9xyp3r6ywLZ18K5IsCBNXlCDA4mL
LH+lq06MrLIOZjkUfxvv3lTbnl643GcNIUspN7JHbAV3yc3eVp0ll5Pr/k3K
T5Az6s+3CDpQkoQFz3yxYU/LPmJ1wGnrx4Hr+XdqqQl4c2Zyl5e+9yIW1mKN
ft2hjJHwYZnq/+HMm/BpSkvoJ3FOCkcsVFTETUJMD+mTX6qsyeINEtadLuyh
9oxYZllluH+TDa/g2obUFonYED4uNyJ2+jx2FKBnMZs0xpnhrKP41cTlgSWD
VouhaO2S/DZwgoqvhVrAF/RjNKMkoB8h0UJyJ+XabIJ2nr4vc2yP07i7cZRI
ALbbHdhMRwD94vR4eyAIKLI6LqfH+S/1KWq4H4+SiD5Mxsnh53tL0gh0uZvQ
rmpgJEzuSfZVY307fXJU0v5Jr0eN3G6P9XmomMHYDWO+YnKOkL3DFOVmLPOO
bVXfogiKVyWJ/r1XpNNeSEse/uii2tM21FB7+416J5JlWhkCO47sPZXfRFIf
8U0hpzgyS+kG2k0bjJBuSmeI38COIeYyBwL9hUCXuEl+fldxQAbIdYu27nY+
VGcXv8TEORqsY404ftfagJEMEJrpUamDxejlK7Ckq0/kmM6pBswpRQBKsepS
XfdKhVPYM2/RHca/jY/OFr4lvsDE0hFoKJ0l3YREtT0XuLiijNwLQRu8lFm8
24TR3K/bsjQ1DFslssMdXK4L6F4pvbxGcEJjsHsRXgAxZpJWzYlJePY7IZ2B
PgqJu4aGoh+M1GhcOpRoXaUcnMB0oDz3C6XTHeTXfBsCtlfAnJsPQ08PTym9
UA4oDsjo5DmWwXWZXRYjuiw+CMtlXqssMza6FjVxcmSvckrxUlntWIYuaTxR
409fCn/zeZ2Y9YCh0gm9EKt7GpFVpLcQGPKRxVGZDGWOQ0Auqaez2mhInQAR
re56/Myc5e9QtmYL6NdW6Df1Yw9nB+lPeg2Hh+unsVySojjfXkKp0xIqkfSp
XCOp3IRwS30oFcbh14R14eA8ufNhNHQtWeDLIMoscjeTD4ZaP7j4Bx1Ei/oN
n3JhO56uW8wL/y6cIxflt9jDp+4MUxScq1L7xUaCxjk9eRTFub5RN98o+O49
EEFuSLutF8Acy/lZdRULw6bkBe55Ks+8f8eoYm2tZ9KCM3yZWTQKiT1kLfDD
G9DvWHeOFZpc5v16Fe6mEvJQpkpUDP0B7N5jtSiPY9bWFa3EaIgX3c6i1wUv
YHxeM79ct2+RcQTHVN2c6uqPnDIn2qr+bZOToIqqkDsO1iM3WpvVRNmti0Nz
yPT5EnIDw8/W2ho5E32Jx4Mnxq6Ijb52dqq9b/cztIG4/tLO/nBzpZoA2xKP
gPUFzgGOH1b9D8m24zHUeu82Wyf3tuXCjt3ckARh2jj65B8DjRjJkdfvtZxh
nK+k5J8UwdTJntEO9khcGAzwj/vxvJB7fx67W+w5hsJHH38oQ+0WtRcMrKck
sMSp6zjEtZ+HQRj3CITkxlz1n/p6x4esrCNn2mk0lUM0+ZHEHCm2+78+8/UQ
/+vQSv8O+FmtaS8QFIiuJkGgV3SM9LAOAcPxS5ZHC9RX/KcCB4nvhP7MWUO2
LW6c8PatXFvxgQqEmU3ujLmeQWQhkNDTfqdFf7lyeq38U6ffSKHOhZgVTGWW
Simdv4U7e4SFWbU6ELt1Tw+yNGiZKL4PuyuQJBJAgR26rMRcuQaWhSTCVo+k
JLHJQ2hTjN7hdG2ekpte8uyzQD5Ha1xb5ZEMjHjW5D56yQYUpJlaAMz3+GGK
xo4SbnB47PlczSfUiMszpGqhw+D+8VYFeP1QJmAiYd3V5Ofkxhlcid3bjXy+
fPn3HtSeFs89P1aiaW7SOGoJW3N1YKB77ZcIQy0wZ7kRdDOYg1RsP7/AdEj8
pOng2gYUizR9dj5K4mCc+yWrH2zMQOQTU+zZp91KyG/KcdsM1sUW3R1zF3nM
O0yDdegMAXoztHGYmZ/vY83IN77h3APRVNcTGBEb1ifh+jfxFGgYZzlv/mDV
+rHiNihizBwXCAJ/eShKsiLkAFhPKElz754Qfa8XJIZgAu6JkkD6dIJ8iwdp
GpY2c0NlzSaSCW0fwfUc5o+0iUb/59MJb8X6J8IRIiQ4z9RUENc/OY3UD0qM
B+CE0L3ppTor4wnBFNzQ8NKyTTboiuxz3sj1659dVbqoxo5L8ZQuLhUeiVM0
/IlICWAQiuIv9lKKRKxnIbnUytyJ/TQaPkHoYnd+XDENDL5NE1fctLVfY0qk
wuz56Tv3iJoPjDchhu8EdS649ilCoP6N0oLMLQGA4c2lVA/KTRN1MOXB1jKL
+cmIm8Zw4jaZ+00IiPJtDCyxku7A2hlIxZnpoM0aXtglA9OacJPd39ukZAzx
q5ieEJrCiOfTp5eftQBo2D0vnlUDZEjqYRaico2QOZa2FOzZzMGRSQLwggDy
J1rI5Eowes8c6BiPfQkL5FsKGW0oPO7ZGeabCiAwRUE4EF9k2aSr52NPa/D6
sYL/94IxZidjSUv6lxvErryqSarAZZO+Ov3m5jVdmVD2pCymQMhTsMLtAFb5
DBjIA3HakajscGPsUf+4ySjKn0TjZl/3OpIzFcbnTxuWQg/Au82SCQUL9vXd
MC3g0dbaWd/3BhXVRDK5l25IOGIo6nMwqWMaUt/noTKgM6rkdl89hCEJ1xgv
CDSudjJjkiuCBitTLeTmN0HtMxxCPEelihK/YMwY/UVBF4HKm/Y14PNYrn2W
W9HxdCvO6ltD1EQMMN1ZHySox+ochgktgEeh35ugP51FlmFr0AN0ifOGmqfa
FFwi0Dj7CT2YA1EyLPC77t3rMsR0XteS+MbO3ysT9uNhN5J3FfKvAG+aAKdD
v/nSFaoDdd8JrTqMM8CvKr7yuuw4yz9jPFv7SrviImY0a3Q2nMB8O3X/5lYe
SFYHOgy7knVfTG357djLFcTHpabP/Bv0KIvmEH5PfxjDtDjS19YG9kqXXUBZ
Df1FyeXJ8K6x+Y1LaSxRSVL7lO3/KivLvrhXx//Wm/2esrltRRLqKA7HMhN1
6v9GarMxNNlNiigijSmd7wt4xRfp2/lrdiAVxqBSK6cZ9lByzP7WF0Qmzb+P
oPUjtQKlUf7CbR5jlAxIsfvUdiXp255fA7lzg1TsVciYF2WYVTdMRv6Wgxzf
5duETQzd9usvTWi0nPQbHHSJ3blxVjMM+j0rBMRxYO9Yrt22lthl2ZgvmIiO
HYFeoon81iVNb+MMwsu9aA60zM1/O9sVpS3a8DTAZHxIpyuNOsaTecnJiw/2
ZswujJPUftlAy/vS1GJ2D5y90b3120+nZyLUQC8T/reDatHyP1PlG3LMSSfA
5FWZxPd/j9nkepMEQykkju5wEPOaL1ex0v8kCy8wPkNEqLAo7FNxXHrJbCmm
jNXWXi9gVDDdPNWyytyi/zvoIoUCPFMWZXI1AagZggIk43X5He2o7nmVKNhH
ShpCAXvRIFl8APdG7y1fYiv+pifSaTEjIwdfmS0OzXtDVLql4S7kW+xujqCD
MGKgd2Saz+E19ggK35P1hGVdwbrzfd5C9WrrMo7IfW00Zy1IuGRSfym+SCqp
FOTTX+mlretgKOBTxMamFwfj4azPm1xJwO4FRNba92M+l+6oPZcWct3XIjEn
U11IX3qTJBE8FQnQnEKfYXbvdVjBex3DzIYL89roMdO9dE+GQKAIRMgf6ZPS
/bfXcQ/mUNPgRQ08Yx5NLzZuqSbDTTRpKeGIxANr2BFz++mnQ07UhJH4s057
6zLchP17UEFaEUgpQe0tNr55KjA62CNuXT41js9AgtOHkmnW3vuY5DFN1Whf
NbPGRHgi+0aQOP+3eEfln8Tch8G4jseKTG6F24oBXE/H1f6kC04wKjmNgAFN
Y5TOhgbWeACpd4Ta87eB/Shr0W2wgAvyU4EN3iTJ9H/2o6fFDMdONrvHbTT9
787P5Ttzvg8+fq0Z/Q0NdTZfex0h1xtA6UARfxDc5cj10ToyMLLkCg6ufIsO
h5pPI22A+1vs4IKUvajf+3MKORqVZS+L+9cPywB7zTSMtOqOhYkqpCmbyUT9
LyvhLnC6krGBpKl9Q3YVAwHhvNQKV41gXRYO0Cl05+UbEholC8OfRaVcbZPn
TOZ/XTfS2XwV+gTY49l3yPzxauEtv/GB89a27ftKkqtTUkT9CFgUdzez4OmH
H+ur3mwMjMpAq1SvGd4CIA+d93uHQA4zttYdqRfqQE+HuQhcgzIFdn/HPp/T
GOqf5O0uUl7Orbs/+NGTw01/LFpVlnfR2NapVOkJGsiXkPLWiKWufsGqQ+qU
m4Cb1L2sdNRF+kltA/EiSwQ49i6hx8ukGs2wngzThh883xg35eHyWSI/yzYO
oBC2OjJ5S9ANyIT4fLruXa4rN60DaRPZfdb4g3vg79CDJBifQ6O7lBicNBLg
1S4hCSdkwurmadpUXJIKWfZwso0lA+V2yukGe9TfaYJR4hauKNmz5OkbmQ9J
WXr7cbHw/YCIC+vHIt/SGJQQ0aW8p4wthoYKYA4Ih6V0i8BXyg9JOeo/ytCR
XwzfC3+lGfrIm5AxBbYhB13jZZJipnIzQ2fw45Kwqfauizt2LlT2dIXySepI
itQdOHXcpjssmgU731WIDXCpN0qH1/x15vivXIh0kRX6YrIGuoMSZbWIqD9g
d5pZ8XrrhmaOT4uzHLtDo3norDewMOeax7DlwDVnzkfoZrOvKcJyBv+lqlsn
iPSeVdm7egkHMFOPYLoG+ZiLz2uTX9PUVLJEQjlcaWOgXxKqFKzVJHxhDxuQ
GwME5pxOkba/QFgukSFEFGZVd7IIURZJFAXvMY1AQxQUwC/zNhdsXoOjCQ2j
XC48YobcB03mSDxvjN9wgRtKM+AmdehAMgR+ihr73mnvFKksyCITHkQatHX9
ukv6QQgoDBi+LnKGr/ZEvPLg+EM53YE8+3P5P5GtD8rq8Y1xDrIARJ6ArTVj
9zn2fBY1ua6WQ2o7QMrSATQPz8KN2+ksru5DwQeVfP6vh87ZzLEyx5PaBnu0
9X/Cp56DOCFwxgTo1Zr85KuAjbcxz3O2Y/VhCXOn9Tsd9Y9+LqYzDhdmitY+
oa/0jmCrtYoiayNuAHI9gi1o6zZhULfOsky+E6qJPttZVLisdpD37/A2WfPX
6B5JOKQu4Mbpi8LUZi1IyDTpwp3VeOcfakv92vS8XrmIiefzXGBsdBmSmuB8
02okw/jp5hyiWS1CVjuNQXSKe6WvoVE7cpw50+yQQo2Gn6KNQ3MeEZKDXUYT
FTIJl+v8Je6nyXS1U9JNXuhx4jPJRXRI8VQTkYF7WRgF8tEmyHdNZLXM5V4F
nvI6P1CMHmdU95vaZw/mGDtUnKaHsymKAWi76BaUpF2QQYSdp2giUhs13LGz
/6zlwyF8aqSFBl5kWAtojWWbe4995j9nA+/py2NKmObZP9RAndL0DNCRT2Ek
JZ28n/4YbvVft444756O7zShwnuzZKUdyoHurA1jv0sryWU+HA8G/C1IMbI5
m9pq/5B/zZrv6GyTc84xuSGbFBDWi2LUznpLjipQO2dTuhPCLg+MX1hYbY3S
sUPmhiXC1+Dv6ellyQcnIOihtjeeDf4vgjbDH3QdwlAae6AUtvbqfFYgo6ml
XXF3+U0i4thJhKTLEK0aWFuR8bFn8WAdLdRdJy/z5lRxSD5LrF4uZTkNS92y
SNSiRkK9wyYeYGJxZ2Kw2bpxoOuA+U7Jv1lc8R46/MqPHAEeevItUcWpCrso
O7HP9TNJSvFIslqLravRPujxWxEZsI3JJhLkNqPSTF1CyF6LPymXldH3JAAb
yFwAhTLbznYQuFlpI0Kk2X2XlYXBJEiqqzVrfAO2DaE7jM9UuurgjSRiJGqs
m9qmLODY3F7E7MJdTiogeGctGMKnsnPvERjYujPpxikyGYa053FfWFcXw1dW
+axQpe5fmNNU1pBXyub4xPEsnVgYtF1UUGXnoT8DEvlBNqzZd4FTesjdOEOD
c0gRyoZw5/N7wtt/ESpBMIdCwnMBkM1utbP0eNlTuog3BHPJVWZgSAq2mqRc
GucA912M//tuq7rr67NjSjgsw0wuEYH2w5H0xOdJWPN7DluF29o0IAP2MEe8
tWeDO4YOaSz5lMgK9t5dmTYnr5xHYAc+AUmmrgnOEkDLId+tLrUAWrn+qeid
HXi8wpLKTxlV5PJhXZp0od1wLB+eH25O87Kh9PobtGt4NXbr+O9bcpgWwhgD
iRGNDfCyUdleGzWo5tcBzWObNhfnzQvG4spx3eqVujYqHSCnfWF3NEI/Viw9
XRnPwGFzu1vRSjpw2qBdUTwgGC+wBGgw1TSrzveRljztxfy8jmaoLF2BT+bM
/0qe7I/Hpcb4D9G3eGPmR89Md1qKeJ9+22p4qIFxLb5XAOhQf4s/T8OzY5hi
ubhS8dC3WYXbqqCFmZd/2VvOqQp6d0CSlE5x5iADiMxLnL4d97mzXjG6Nq2S
n9LZRVfH3UTzvAMYFQAhd7O0QrTvY0MA27YwU9YU9QjMdATtCP+eqVRl/LtZ
EBurz/Jl4ZtTCpWwJx8fCzqVGWO11Xom29v9tdzBvDOsCm96wbl7tMcRyHMq
pRg9CzOWCt2p06fLRyhYXqnYGh+lYc9VpqlUyuuGcuGYmroto13BqldJJUgd
ycCZKZuttNqj9/0FMBhFJJt4F8rcSZsmpsUDmhLFAzhii6nJzL06xWiggGTf
frKHdg8LnxdY1HHeWjnwyigeZjl5pV+UmeEFCZdvWJRjdzKLb7tB526Q6nCi
6DuTt8BLLoJg7Y76wKU+w9Jfvazx6aSmOY2stlegHeleXFVl+JzpNbeDb1pc
vM34Gntb3YeaOt2DQoOtHXD/zjxVJmAoICAv3GJNdcVsrfMootJdTU6CN13/
QznPjm4J5LzVXUmkD9guX/EZSzzEJ8v+NCOExdwVWihEw3rGkm+9PzW1Bkum
XemhBHYE45P//rSTnywenL+aMPSqY45SlSsNOlL1F6Dhi1Rvr05O1TjkHMyp
TLYmoC75lNTp+ulCbnZwvy45xxpUivm+e7igxVjCVnKEwi9eIPUQxhV3ITKE
mbQAlL703LORBE8cwHq2R7Rr8+gLCj+cg9kgdDjUSlPmZYopn/fu5MtKNK+I
cHcwVjkyQRU1lbLeM1ZFeEGyujLzYkjpVRk5i/YlroH1fHGGc61m2xPLYPat
k0SUhoA2vEU/AYlRWwUcjMW9pPwQonrXw7YouGOFrm0k9Wjj43iWyPHuIIzO
CLj0X6aEx/u2w/VVwyT/cf634yuhQhfirPx10vl4H19nbVN8JLogQ92FbsUo
WaszVpVuE6q565srImX0pItKW06pE5XipJnvu6VbEXWRhkHLvlIl3skT8NaL
SmobCnownWD+LdwfM0WuWzeClX+mxFo42wXS6CqVNzacnHbm51T4IKPW5VFE
TPigxxiDNNCQsTN7/14w6Qqpz+nJ2JgSCJuEWt/W6K3wtveoKs2084Qmsbgg
jFdj9n8+9UEZx7KZKqkXA6M0ErlEylkiZyS+yVyDatqYrM7AIDlOjkjczvv3
MieUZkaPiiRhq8IuqjP2IsZW+4PlWBanINSw2jpwTtCz0HiLKbjccd6pBcj0
iRCnozN8y5bsjXXMTkV4pGuzgw8Tnq36MlZA8cGz4qbYywxIkTAC1y1e2U/T
KcPa1g6bkwxcI727s8Cq4GqprGfq6yTX+aF4SR2+qhsh7XD5Irv/Khu2E/yd
bCuUKdFpl9QKIODBEBUujh3GaO8B9Z30c/OVNUATe3EYnZctPBNNCQWDZ477
FpmrZT9N3AwHkd5UlHum3tkSZGVi04+xZHI76u7PHXDRnCirudqgiNJx4kme
Re1gsNb6W+OPWNIaqk7e0D95IXV+Ab0HbrnQMY3ZCJvh4esfPTurqOCUaer5
ZguVbWipBpeuwmG3y16t4jJ/d2CWXGdpSiYiGovBv2pzBf1yWIgUZEWYInrq
W5sKnP3Ackmsrha0NdAsdb3TytQS6M9I2vl/I/XtzmHBlJmHwdZtcGvNrvjV
waRZdsr4zsb3wjBNjJ+9TZK141EH9u8+zMG0iqRHTKHpVWmjiyBu1Xrni5Tw
q/9A9dTmw3NRFxqUOHiiQuJEd0PnzT3aaeFodzN6/EsAUCWwQHqCdZXCgbny
hSsDI5KlMVsBEXtFqLIEIslWGuTDj8bYFQLFQZJjxfbueusNLO3U++ieQCtO
mHQxoaJNXFgUPOBnSiwLH6Romq8k2WFTEIaHyzt7fmicMru+27MxoKInmdAE
2r2GGbKXnThMH5Pb2ypcP14zgEoBD7OodzL+7R+ajezVGrWO0me0/JubwpdO
hHUSjVoN7eE+r7SUqkSPetNIychZoMh5HNdRjgGHD9p2jczSEi31oshOVMXM
7RZVsuaGs6uNCzzZ0a6lqyaM6WDqLezb07azv4W9rSVlgYhdtWfKod3AUOa9
+HBEGt/vmYGth0lJeUt8z+xNIrFkAveL22v7WZgZt3Zq/EEfZVZJcenr8deN
VjS1dBMFkFkSdWr7/xMKVDLxw/U0b8TFxPkI3UJquVa2b+9MEDE5vOJWd4C5
69LK+Zxkl5ZRelBP6WW9UIxt+4bh97crt4ePBCpp+anYqOBGoYCfOcSUJSGH
dt9U76SlbX4wNuuhOSFtbIxPkHPgx/G0ZSuXQlxenXD1eux/piuyILkWQ/VZ
EDwaKbzoLLAmbYAqSzUSC2xwCru9fKx/OJ0FUMyNezWcJXx1o3ZZ3qp2yhmJ
kvEgf2qg5FQbZXwTsXfVKwARHy9KOUwSmct+RGmDNQPXw48TvbEHf76fdwI/
gPQVua4dU+u4cGAYvfIGbdbY8umauOLed0PAJLY2o/GwdN+w+Pf4159sfWM7
AEEmE9RuOpAW5mdVfTU22JPuODLKWJksFONOXWZsDOHEUouRatSEKz6g3Oh6
ZQPI4GrSWqcL/afOlcmgHrMnM7+xOATX8qLiSMWD27tt8P2Ns2GGc8HVSRUj
B8Os7HdxanjQgRD/H2sbjbXrTA0H9sRM61gv4c4fo8Omv8R3+nHUyJqIhODJ
0H6e6TvEU9LP8cBdnTkPO5Mmi06wQYmYH8tbqY+q3ehZqZPdVJIlbAODC8j7
W6p3ZeMuWgQiV7WE57qSTiZx1XitSCSnPxh/0Ypu5A/4ucLAHgDh+mX8u0eP
bzst6YBoQL+Kg3eJQPN7T6oi2KpZpYVqYD9MIe3wV935AMcsZjnDn9NR7MOx
dTXxV1vZZRVfuRBsS5uOd5o9aSvM/FPq1y0hgK2gq2GUCCJpv2S4SKzCyVyY
jkmoux9NEB1m5aMgcZZnD3/36FP0Gdkfq03JeYVGnYrG6aG5/6eIHilemH9j
DTQCS5dnZcdECNAVlllEkScv5Tyxz4dEtwLfnd2LUiR11etpiUQNRGfln/h7
HU+9R+o94aNrO5eQHQ6C4fybid9c8rmMagaRco/ti5UdcbrXo7LDPkDsIr4G
rkvudQFx9CjqQLvWtizaRXwaGJItApUDHWdrM+SVrvxofm2lLMnag4FopKu7
CGFUJ7ILNM/e1IHO8Vxn4f2MIiwgvzroZk2LKJiaPzTcS4/GfJAFmtJeHE9u
XJcwmVKEin3vnb3eZDcWaKjuZNCT1T135cZwZLKCp+BUP+xs5LtRnlLbmltH
qy42hcyg0ZDR7M+Sc4d6PaIm+xgeelDHq81r9+YQzklYiWNiAag/D3LtEY0U
UkPvf4duZUop7JeZKbWV7k76YG5T480ZPVdEtZtLlhqOX2bMT7xKWrL51lXb
0tqvpf6ssihtdDen//4ZIqLwOG15f6bar2NLdNTEm31OI3T0fBVtyKLi9vMD
0wQGeGSj0Cxv7C9zRcs9maX0Bj8cnVGq/pXau7uuFxgTfXs13Sx3HJa8vXAj
g09t2xo5vltvB+tfsEs+gdZxPC9WeZy8WddF0c6H/MXirTIO1evl+8kkzt51
a864GY6zGL5N47ARTQ5iIQGBiSpveiKGPenDm0hfngD4iw7MdhVy6uFWVBvs
KJRoxz0Lig67Wm/j7gItY3M3bDDCyAps8h8n0aWX4WF9F/cJ7PZB1gZzsA4F
qJJ/cY0TtcnACve932vX4TTPHu0h62nsOXJNZbFCQx7rsi68To7RDnyDVCCn
tPFGnBte9yEx4bj7ETNkeIuA4dO0s05yZpRjIx3QLY/EjqtdQnxi/OjCL0Gx
BNESIUhL7Fi/P//OfaR4SMyA3qx74MNQY8OK94SIbLLtvLRaFNl+gOwMW9t8
/Q04fl3dyw1FqHeemOUWQWYIaFMrOoL8sUfjd3e3CJuGPXxd5Z30FSM5BV58
QXaXrR1KzJ/eCKjwHtKQjb5BJuVvf0rPZPc0ylbpZf2exbZTgjJW/AAFvThK
/+8A8u9e5hnAtz8KxOCwxSwix+QRLjh3Q8Q6rESIUSlWglsGu1eTyK3UZPh4
ZVcos8r3P8qTUwEuNBpAHv3Yj+gAv1n7E2AwlpZCdrKYeI9H2iBya/+OmdFV
SqIjGY/NPavuF1XIZ7lDAs/26QI464hbxxpEFCENK0BLdiN64T8d0fwp2mMO
gjTm886JI14oZDT9M+KUaDrojQfiu5+348idESNaSKtrTLsFDmL5dnQZKhp1
d4ZyUpDArS2T3znK14M9rhXM9TsSznzyvMMGo3Nu7ADmlfyil9+ivT962mxj
0BG43619Zn3AIXw5r3MFTJTR8xkGEKcKw21x5/Ail4GE5+M0YqMFJCgyR8JE
1GrT00sStVPFby5OmPVp4oC0cfVCi+OgHbYPhF704k9ax5kC8tFOaeE1K1RZ
QVhYsJxRYct6Zgv1K99EyFOe0/11vTY1pE8X5RXjKJDTLMlu06b6LpBMTPQi
DD38THHd8/SuZrX4wDtr9JOv/K9wXOgTKsQQfjt1g2aw0kSyLMHsOsaIdgyH
iIVvDy0MCJPNvpN2g87T6x8RRh3uilLeeik+EyPiUrlQ9jsgzoCpJFQnEdQC
9/BdNL69Mc0tW8+zW231o2pcNP1jJ/8H8BwKphC6tOnmcZ8huSNrp4k67DGO
dZQkrWm1ux87erePJW/zulVKR1whFqCG3viQ7f6JooT6DZZ5WPXhgxsvbWwE
gjcI3frRIXxNtk1AK88ngHcsLMa/iRH/YlJYQVmjm6sblIfF9tK1Zal3K4Dn
k7vy61D2fsEiGQ9BRh7GTdHhQAC2oZBWLgcROfCfZTLQQ805PkYAtPyZXrYD
kGIuWOlXW3lUjMs0kVgTcH6kcqRLlb5beEKO4I+RuFnz8AEtVqPqLBfLotBb
YkzkoZrdtoLlAE5E1vbyqPvZSNThAc0fFjbMaFN2AKKQ9Z2rY7u1FmM9q5xP
pwGjcV41QCScubc0Ixb5q4S/NTTITFFAS1s1Lmh7Vb0h1hZID3NbxI9Rx6w9
wJ+y7zS7VVnRFQgdGKlWN7N/HfH5JSDEUoK1MAAYwPD5UBbkCMsYKVwnwq4Y
EB5rHPjLsgeqv5B/rRv6uLctswWvFVYw+eoIQRnVgY1ryXPunGj00BKaIGxS
I3T0gALpXKr/CAQoaejG27P9fFQJyoLLm5vQW6BZRtssUY9t6DIlMOjVbO9O
COqII7IfVQG28MCyCRJK4RLhw6jXng85xyePzAmyX1o76JdbRHx+MpgkVhc6
vcIXfrR9vEFVA1j/AKSVZJsPV7GjHX67aAbR33PMEblNa647LCuGt1MPye2f
ho5O1lS9oO554uXJbrmwWzqUJgNRNp/D9PBYZGH2zjMX5XF0m/SznRw4ZcCJ
0CK5j5ZfJ8iJvY076lVkbSYQtOlFh8aYgYCbDMBYGUPleEpUx/pmXS42peI8
eebv5KC52t3Rh1Ky3o4yBV1qct74QPNoAwfwvsMWonaUkUiDHbx2GFr3GfvU
agrt59fvkIhwznM7bnrsMi1QaYFPVxNH382+9RxZL5fCBGDaIS+Rw+JLptZf
YYZg38T5QRikU6RvNpXEQM/CHlS5XrBHMezTH/GVFI9CTdmjzYOCUAqOw3Ht
l7OxWK1/bJ0ePVslrh7PM1jtN5ePWCbfpVLk9XGD3aCV+uJ+5WPXvzyC9J/S
HYSKPTooZTtFPnhv79RWwHQI/tHR3CaEcGTsLBTm792360edmpRsIEBo2vUf
VvxKjGrKYWBKPXLtWi/EN4qe36D9gTz0mWPW+7X/UaBLiscxPDROTthD7VLD
R7Vk+Qikrrym/7hoxl++cDCl56FlkFoh5hTgSQ8scDPjqVz/MuTfroIHM4SB
+nAqiAhL1lugrlR42leSPJRLlz7qiXIFiEAvCpqmaeNLt+zYgydUIkqt7rzr
Y+qV2v+E9gY1UwdV1q9YBgGr0wf9Je/KqE4qPvmpVddoahqn9rrnobakkfxY
KzVgfhcub8nVJEDQVdEpQDBcWwJvfVyBcW66PNbwaHoLxztwjeZ3pe4V/+by
rrrAUR0xh3yoDO0KesMajVYr0yM2VfdrIArrbhL7eygy754Q+jUxmg6biKs9
r7ehoIpP5gXRNmKCcosjEabF4LFgcoXYTnvZdvrDoACfUHqe1KXA+T+kddi9
ZleK4YzAzaVpwDd+JnjksMh2xLD40lYmyrbvk8AXXH++gEFZyrEh7sxL7Mxn
Gez/LT+wnkR8OMzpA8r61aAXzfDtDfTBZ460nxzxL8bL5SqAW0rRQvhVc1z9
gD0SzyCYzjHQTrGr2ay+bLRxuHaDPmsMuAEFoAJuUVqDGYVV58EBrrsML3YJ
J8Ac898A6Bh30PZXG4dWA3bYko0+MM2/AdqVjm24FRmPliDvZ6bWQTiK5cro
O8+wYJCtMLi+aBRnTMSIKjRyV/pKSIVT1CHueym1t+EWNkbG8NuyOdmTVCZO
S8XFx6ok88TKndJfLkfclVgV5omp0LbYp3gFG3nMjZPe/2O1e5rPR0Hd7dTN
ReC81K1OE3NRZb1fN7EZUhYupuVMhbO7ALns6gC7McT95qSL0L0v1MOZxbZ4
Wt99SnFL8HPPyOfgNdCW4fIvXLWqmTesQmlASwN7+wW2iIkWY/BiLUxINT2E
mdGbEgJa97KYj+rV4ley8g/z0GiltP7H8J0FiLttp2SVQ8Xqruc144YPVyck
DY2Jjs/rrS0h5YDeMvdXjBc3wqoYw9mP+AG7oByagmH8JFUzu59s5iO+qY1H
y/XSjKpZiC0tLgFAi+ELphMI511f4u6ZVHn09YR+ApxhCMrMqhmfLJ6ZNxbN
zGbTQ7vVtKF4qG9rO133vuKlXSqt1AWeFUDM/hn0V2ndfUoBvGLy65anBxRf
hlvl9b6gls+/2VanxgqnK3kpaQx1GZkVf+ILgRTxlVPfjCMBus6WiQFOu8Pa
1zXeXZKn0dqmpQukyzppK1/JEB7NM2z/iJA1YHoFCuC3csuES6YgJaV0y/1V
jQFUnnKLZFbhdlBZK72jqBUOH+lokzodKE4gzdSwzuFJUA2zqO6PNtZYuE30
cbtaBili++L9KAAbA9NKfWnwkimv05iU0RizcPowX1QnplMNwibt/x9lhdQ+
U+dOkEGy8kJ0RHPEHBA58coVW75x3fF9nVC4FZGbtbspZBMYn4CWBiN/AF8x
zv9J4wlIUCj6n2p32zdq3PgFLOutDtUGefMvdNmLrrVjGIO9uCBEOjIHw74S
zSfs6VttLRrhylBgWSDG9cChJtU6+YlCR0GQqx6xiO9jBnIs67J3f3dmFOsM
wmDwp//tmSJQyxJPrCTAVSYaFStocB9q223+msphB4acK7M0T7OEX3WTtvUs
xDBqMTyvPdQgKxNg2KiDQBwixsZvrC8f6pmNF+RS5WlfnoQ4G2jC6HBIX14C
5StqBJDMMZhixuXM5q/LlhLGE1a/tWLW86ynorYTKGc8I/STYBX4QowIMWLW
jdra5/svXCMyj8SukSE3gK8eYCiYW8jk+H/xZ1HSFyta+s9V/CmQdu1IvDpC
ORL0OzA9vjMIGUcHF0j87AKqbbzTuoou7dUnt5S+hymvB4WOzhoqbRgEaNp5
uS3XFVAJjgvAu2oXYPPmFJEgABQ02vQmfIOalAqIu40CWN7q/jdI99l9eEB/
1usfUnmTK3MI2jR+srWSkLbx5wryT4nJDnN3LU5ZKOtqzFw5s/A9fXpZLXd1
MyyneM1QH7THP5JjqoO/hwrEsrPZKrTbZR50hNd88eaqEkW4NdSC8Ysf8EzE
BnfVjvz9OMSdSL/rjwPX4pl5uRGtffLDXs12lB6YrlNHuUKpLOITalRs5/aS
0ZIn1NVrLyvpTnjZ97kYxTssfmXrWJashozuE5eFqsnOXF4WWKt/v1wg3bb1
eWUdImBQJHEZNysW7zAmn6Q9PB2avEx2AZ4kVqqQjZsU40VdmgEdvbKNtiYL
mYAma7LkeaMU5d4/qdSJJvGBgFdfvv/li0eTWVM0NtCJxyuPvh5f1CcEgU9C
SKtpR+t+wkGWSeK700lP1InRm8DpqvucV7FjwAdFDNcwdz6CzsTyDjYN2vxp
+fwX0wUzUErAV1Fyr232t2eTV9rwILvjxPc0dgWARxjlo+lYaBIuXGv9CBJ5
+J+0U1JMtXmvCY2/SvaSs56+YNoezItK+16XIGlTTsFH4Cn0O3j698Mb1IIx
KfNSS/CAS9PXQpd7QARZ7NV57BkV4SGrkD2GVYb2NMVJWPXBnsXA45DufF0L
mRSfogxBLEO686BTCNQAUt5yqrPgHPBGvBzsbQ2aUH9R3MAEnG8R4aG3ecVS
Lv/R6glcFghOxQ+mAufvtPaHqU5VnW8EEvFN33qu393g6Ec1d4ig/SirtKdw
VkAyeW2M6d4Efy1V8WA160PobgY2CtKxF6d6LTHZfFdtH16YXIIoEmAnTKxS
b13FuK4IEoTU2yuxl5t6Jeego8jZKIlWEg1iQqWgBHP9IvP6e//sIGOyzllY
g7KXNCYNGlcnlXvs7selhQPNXB+GAcbASZGXRs7M/vjcMyNmJSfLGW7RN7np
+rAT0EWMtSiwIC79p+xWjLg1VkXw46hQbsaggKAV2qOE4z0YPTrgmJ00t/aL
PuOv6ZSaEQ2sbmx4wCL7XiAt2mvRXs+nTCSmgGnwCL1W9yVukBI6JO5pVpry
eI9RdETb6W/cW0gazV8c0wWDUEPenSIvj+jLtj/Z+J4WRUUmLwdmlA0uJW8x
PHKhcUC09pMqOrqJnIxNsIuhnwXT7CbtrckNh8EROCqgIdY8HrEqfWXT2PFO
9X6MIVhkWormTNPcUPrRv4NxLgU4KCSJqKNS5UjneSXETRbfpWUcQCDozUaD
rs5JJSvAuhcrV66I4jdQ5Xtqa/8W8ai1pdVrdFC3V9sKJ6DbWoB/8OIW3VeG
cKr1N3EAOfp031IhJvi0hSydvRuq51TWF0l5miOzGYO/AHwZnKBo/70HxLle
4fFzCXa+if2VSDzIwweQTHjQIlFsJUhE7v05ZbVcIbM5+JOdivZdMExMiQWJ
W8BUPaUjdvvkA5QXjv//wgt24TucdF4yHvL5/FjLoRsQ9ICfw9qg1gt8VuwQ
PGGqLa6CG5uL5hih1bbakkkjALzUomPqbSRwH+aGIBJIkLmwmggyFDL06BYJ
GbL53SK1XvrP8QOSqzLbkfZjKfL57McMhNQFiFjPo8V68n4eVu5Jo8LlzVP0
qLIsTbeHwlfmm9hOsSx5O8fGYR/7PLuQRAnJcCxq3x5kw2R0fHqtIs+qUGSy
HOymkfjPiD1tyEHQpRJzQGyp24ePmKMQXr69FppNaA7wTu4jZBFwJcWeAKdp
4slYrBXhXq7e6DnKbXcJgYe/aSjhT+T3+MDKwKz0Y6YKqgAJ0hiG+TuzoPad
3enF/bBmQLk8QQN0zelRXry2tkI/b3ydV6NQF4I0tqVc3fSE0aUSUw7BOYR9
o67+DJOyf/JGrFggm4U46+8eEcOU3jI26bZmwxShPjUkV8J8EzLvSDstIknd
ErABi2GhU0PNknJllhq7/pfqM/4u5BF7QQCpVrrFcZMss+n3CAo3IwsWZXob
dQPEXFvPko8YsB/+T6AbKcyxdzDlYFsNdLDUpm/jgyShvz05/NdKdd7+8DcP
6elFv/W0f2/l0Agq09wj5NRF0C+LASFopTXdvtl0kKu8vw43iCq/V4A/wpSa
6Jp1Au9Zo0jnPp32+AcJhV1rEzaqFsyuBFkRyBRUfz4HL6Me/iTigle7N/Eh
t7moL6t4PMGh0GnkUsRnUtMzvda2zIKqz3q97hex44WPMxWx3ASw1UO2x45R
uNeLPOTeJs90p9d7qeR7Yw7TQsA8ubcW5N8Ew9fwSZxKyKLu0p+R2om8iE75
u4HuAbIlKAnMGh6/S1ZPv1+/EG8XtXhfrIr5izV7e7gOtV35p1jXUQG4P9nO
ut9uCdvwMLM5mhkVVT+Bm90OM6W8kOuUn1ejBIs8weGXzb9hHp1cGQeQsuqr
jHzqcrCJBRAVvC2bs0qTDqHgDhAXoMcWr545JSVmDhZb3nIbhTFehk6pPFsH
9ld51vx+UZ8N6qXIuCaeSXxK9tYZX9ADxaiywBx+TQOC6lLOVJ2p9GixBeOh
nbaSnowx1m0j/C/uZUWrM6U41etdxAS+ysmf+hTKSN7kO0ZuprEwTdjjLWeZ
vrr8uPxDQwe+UVk0dtx3VJ9pgH34jNlfiFdy8l4N7cwuctGU5VJhOg3j7gse
PNoynQE31MI7Gx6HHepd2rSbHiTGMcvXq0bdgdPB+j4MxeuaaycU53iSlUyj
v56EeWHkzUyAbwsXUvEBQVsufc1jx1PuRy2J5J3NfftD/CuqV0hnhoX68e0D
tyt/++tMP+Aese3+9kFo8ycstESen8fIEQcZ2Xm+ZN2PPcj0VyqX0m49gzQs
VWV1UdVkFVzZZ36b80A/D9abisy8n7U/rulFLau7RE62/HgQ2qa16jKIzhyB
BNNGz96uvKsHf7kpubpsg4QYev/JY9IklZzxMiWgkJFh+m98h3wUCmXsWtn8
07JWgB58engHoPmMN9JukIqS6EFriw7u6nIQs34JPjYBKlfoylpMmbjgc4+7
0188rA75MG2IR7RrvQASe/RChDXI7gjE8lrUSJSST7GKBp02GtJgj4hMuXPH
sdUMpd2VtX7rJV+6p/juoprn+wtYptoYekfigXr+AHSi0bwk4KqrAZBtwAVo
ixDJOXVT6Ukah+WNkLnc/Z/s057IahNXn9NVJntqq82AMQuxByVlpCynsMKF
zJOFVbqKcsPYi8KJVBdftPzt3E05sThckc7L75H+oOn4oJjkVSngcx0ZBB6g
QOGOZglojP/tZqrN3i0Uhe3QlbWx0kHmkuKEUCAcMPKauR4TWpVxKvM4q+AX
nKTD5mQhmR2vGuCnUfuOkAf/ZYsXlpX3assY8snUa7D3yWrnY8+vgp+4aK3p
rKfmQkv3q3IgTHv+KSNQRKazFMvUvsASdX7DhhG4SvXuZxiMG6WIeDw/cP+u
oo5XqdkEfCwGMnulUBt7Jp8mDyJd/2cTtg1L65LvNy7991HIEgdZCc3JTufq
zLuKlFXCzcQ7HuhX0ZrlSyIbPVaF/RwVNhWr2V9Avti4lO8LVtrqFHGQS8qJ
l91wvonMGm4YzgWuU9THxz0qK0HxJhmqReJ33WOx8d35//a8vLtx4DZt+ynI
lt1KvX+MsNRSUS/Yn5xumduwsfzsioHg4P3zJgn4YWCJiBZqHpBeadaRPVUo
ICsFxAm902s1t1YbK7Sp1fJCM/f7lfexQyjRsW4IHv1QgWzSLIzy9wFuqe8n
cQKG1fgrvLV5UmdneIAn2YQsD42FXvTQbwLsD+pObKeXL50Eswk4n1HpyvYM
sxy10AJ9l+wl/p2ROMWsXzlkT11rwpz/JJmZy1Ypyu+Y32G+XFq+gnZcpcha
9M9z1pNBgXbxX648s85Nh+QiL+i0HK2kHj1hHMFXbN9z/YzCUyKfu/go89Ht
M04tvWP0gev6z7z8CzJTY8n2FWna6RoK2fUO8ujXYg8hC4Htl3klH3ly+MVF
M44EK3Od/onWgXuwKfzqFkM5XHmihEGS1VyYN3+5qLFRktAdMjY6I/5bfdTb
IYZzBlSS6TKn3YLItxv49mGPmoyhXZ7gwOhm1p3ynwiKd+8zp+9RS7AAsZ44
mJ207xa1y78fj0mO/HjrG1GhHFneqZtbQAdy5733neFWKfWjQ/tSwdO375Wn
GsuTsPPe9wZMXO/7Dp7fhL7K+9tVunOgoQOQjrGHs8Nb7z95tK2K77VUVc5g
oThoAA202spGQgHtDzPCquMcmd5NSU1ulUmU8OjO21y0NlhCHkm20d+wHeLX
xaN5gHQyAROEpvFObJS/4YbnoktJ4D0pMjzqVAffrVy2cN9Zn6SZZz07Preo
bH96mPCKw7ZIEB5SGLSNhDG/j0gxLEhKcwerhBd6GBxBeiALKhsei6NhjDvn
5YQKhQSyNaK6TM1XZ1u/E8dJaiYlW9BDM3OZzRBu9W1YU7sUmQTiXyOdFkSt
mEeuBlWVhHsqiiORXMMWrpEq6eNxzGYB8KxGxBAseXx9pe+10w1GbS+oXkp2
kHoO+41zvjJxFYEnURyi28narkhjN4WpQmgfLQcQVlfCwgfikZzugQUSWFEl
mqH/mKpXmooyhvSutKfiDsXBJu8Enh4TyzBkMn7mt26gOSn3dKa012G/jKgx
k802N+AmNstydReEyGv9ruibLeXSnwLdaviliO86k5w2QEI7NH3ZIgFiG/r2
XpJ8Cmj3dL0qgKY6xyyay63sZJxTuyAaNANXOJ0L1PTPl/hKWp916MRI2Ti3
0ELuFnZ+N5lWOlJQSoIGCW/JyqjHq/XKi5Wm6+TH7Ll1rDjJSPUmCVRZssUi
tn+vo3O84FyuUHHzoDro6oj9homw7XLTzP2DURL+a3PIizajSv8IQqir3aT2
57LH4SLrZl9PupAgUUtJK6yQVg7CTuH4M9oupf+6E7oTAGX1Ku7Rfw21eNnm
k1k1r6uXobYbot4TX+yI3dgAe7lYNvGiTSWl6QkjDdsQX2+/PP73uCM+VW3X
/N3NCmBd6rvT7XJyDT9MSlhVd+VwrEcEtxFPayPRBi7v1R3gvXx+ZGNIue/9
KcSP7Q5n7KOq3HalVxqBp3jPWaW7e9aoPGWnrICUaRAaH9fiWVvfyvR2vE9j
zMpow+tPlKzdwVpne6j4lH2RC2dOUHhjZM/TXVEgyIoGh6eJB3TBgONgwX40
1Tf5q/y9FUeghbyaMhke02Nq3tCiWxuvHr16nOy6RPklafcR3fJsNrHoJGzw
ZEHXs3vtqeIzp5ZHdfZroPfUqA0bZ04Qy7HGyhiao4n720ZZHyJA/QwATa40
7av2rqgbnAhKMDLtXHYSlNpmhwbe9FHVQBhkrSyTLJ1mL0v0/OL+1q/Qbcpg
BQGhduTHVyBjwy5fmTT/aJcbPynMOSLJr8Y3miraGXQzpeJV2yF7vb3/HUKq
sBoWuq7rXOrCFa0r5Qe96mM/xwrmHPIcSSwW/kvtXJeo0R+SkjGl6v3Rv/fw
j9iikbytkHi3RDdG9d+dX9TRtlKQ8GKkdWm+dpkgLAjtoOGrIAfkqlwzOqIw
TU2z6/BCB7o8+jQXpJbOm0/gXaEa+8ACjkjw/xKArU3Su2qEYsG7gbVHEBGK
FkM3LDp5sMCEshOAZSuZqD0w1GZ460vuZR12UdY5XHiK1THkQvw0CUWj9Tcu
elAcjEl1/SIWVAvCx53HNXlqpFZumrFpRGZKQGY7oj7360b0RILBF+dROnYR
IZvmCvz9TakDvFoP9FGfTao6T1bluRCBPzPxDwMTjzGzGKqRJgnDqc95Ws03
6oZr8TvDdZH7UCKmyYcRn1ZZuzT4HVjUkLqaGIX8nb5Ll7i/vMiNX3DuLr90
hRqNtJlSGEhOVRSikVhNwKKvX0vLUbzIpWjkgENKiT84FAtFwuphuA7YQ81q
Ugk0tYQxL51QjLT2Ku+rG+aA5TsbjToNCVld5R3jh+dAHZ+w3PtcIfCp8ZvD
ORaUJAYzVAFowo1E3x1btUFph+BhoJxxcgs/6y7QcMwYlQ3HfFqkFeaGSXAa
RZsY2hDvY8QQzZH/3S4EXtMJh58Ni7ZXK+C7YRYNbQGirU8XkENSwLIIXgtR
Tpb6sWepOtpQRYFOT6ezRmKP9OlOW0DFvRJ3+r7Ci6Jqj47XrN0e6pVmwwhS
CklrgOcOV+9aSsqoyC5tppWGTmIyIuUm11IhQHQfg63DV+CtL0XKrZbe/n8T
QZJyTKkBEQowjy4Isci7ODHcC3IYqB/i/dCaW+93k+Sx7aUKgPxqP4LJdd+J
QUD4vdCpkFlfQV2SrCYY0G24MPgFVTOlvNnHmuo/gYO3CI6UKO+uDt8xp1/z
wy/g7nGfJyanH5XwlsEV6BF1bUQWJ7rKv6JpGKy4aemOva6TUfjiv45XdGqr
xrcTtiMyJHHdSiNKnfEHory/e3nsNXDfcgC3RsSNjKjk8NmA8VBkJGXfLLNM
AlS68Ry6TedTn44TlzGmrzJqe7G+5HjxdbNCHdCwMZ1wkdJg6YueIntNr2U+
enhj1PIYKFPUp5/ULEIMsCeO+Rqazd8HNVsacGqsQaJXFYVrgRSVVukbFQXH
mxthGT33Hc2M7sFTuNHsbkxfjcVIhqQu4WAlyZCsLq6NbJzYFC2ZQMCvjfVP
jk/Tf44htbZNMCyanhe28GCk1zwR2QOK0ugheqKaeuVAeXlcAy1bopHRt8wa
Kb3vKucZ+Yc/gP4smMDExcNNii9VoLe7hBQuVM7yKuGZKmKWag7l7pTTkeJr
qPa1ZiajMYlttyL+q++2PBjKkG8c9Xip7CW8BbweOP8KLhvCjm5xWgy6mggi
TI8SzE4vyaOhVyLWmQDd8cVxKgBv9Pv85nXQqwDwbjTDWa5Aqpge11SoUNng
DUuQcLIOqi4ILo1FfUt2K6rhLR50+/461CWiKRfav767lQMCPo2nhNXR0ooC
TdKcvgBCS296XtYqUdkOzTEQeR0WoGzsHMJxBTeNRGShg/j4mW4MQ5clj7mX
JVh4+sBRVNnYJPnZPtcJ2Jv6HeYM097DAZgDz28MC4hqre3zWHice/dT6lI8
aBuAMAN9CI77IBInaU6QXLspt14Nq+ha2yCsnCBC2L3TtOWl35SQzCtKQmIt
7sZovh8plKlVfmbLluaXuR1U2z9umAURftIB/Ox4elty5/RYWqUAFdVuSj59
2bY1cuZSIPV+Ahw2jFxC1G+AvC+an9iBQyGFAvnmHdv/0J1B8EOMa3M4FjJ8
khmzbXnwU20ZLBjVjBBMZYyS1hv+UJLrjmEy8+CLTpB3V1a/GpcMw/KHgZTJ
0T8uJJGIH8CB6+LxwnOkDI8z+9tuqJWAy+42dmW1zwAJpTk03UaKu5WvAYld
vlSXPONgAq4Z0iEKbjAtC8KJdia5mBdbfwlRgVxx4oAIclEtStLmtOE3Vv7t
P758ONvfg31FaoPn40an/iN6yY5M0pOTt+GWspUwBnDQqSpwyB/yafJD1ayZ
bOtXPId1YROwNpZ+Ba/jgvEj8ZW1wnBp3vDsWvCAKihE2dli3l3Dq0O64E0p
Npg+TzqCKOafb8QsO/5Yn0Ud6lf4EGxGEBYkmLxX5ch3PHVeiCZkt/6qg67r
sQvl/CenjSpbvf/qa3mAzBaMplVpcqv4GLb8fLbs7Aadr3aDlnC4fnCvX7Aw
KSecHuXhZUNx/V+xmgoiAGIHWH1PS1X0bufc9+O6XhDL735S92+tKNV06goZ
LdTQU1qogTWa9CNFwHo2H+W8q2aMhO2FvyztZs0/ZwKiA+lF4o6/dQPRc9+5
pK/9aLVSGTRekSGmDCc79D3m2Yk9iQSWbRzd0+eSQTlH+YphgKtHZ/UkVhUZ
v8HfK/i2eaVMxjG1avJA8iG/IVTyZB1Px6hUebaKEjxR93B5iRGXEUw1iPzX
RD/ih9pdKJ1gzGiUIYEf61vEy5x+iAzp/LOYOp8fgQdVBUqcZ0O6w1M3wiNI
k5houqQo/dYQgYjmrXRVklZ5xDe2Btw7iC2d3oWyPaLWuArdYDYtzysGioyS
u2SY6Icdgol0lH8+29waUDWoZb3LwTgEowsQz8UbYfhjw1tH8HPUg11AvP02
iB8Wrq1n5vJ3UQie0DQYrwkMP1ViyTb3RnDiS7s7akbweCCzyuXQKar9MBz2
Sz8yhQkhZsBsRJ55Lfz30fuy5xBiBlvOLxB/OlBeYvRMP9gtT4N7FKpasI7f
h9AAB4f2CVXCaw1Era8MZF//AiVqrKk/FpF8DBWuzSbTG/MVDAzwkbyPqxFk
IF/H9t+NZk+Rq7slulrvM75BY9LErCTWOMXsSvb4AZgj+xXRHwHf+MEEZo3u
8EXcV5lnbHR/Mq9MTsYOuBhgkcevBlzHLU+x/aSThy4bMm2YLiVZayTB9Ul8
+MGtcS161JSGOm6x3u8cbCRqFpG1SNlBwD6e2Ar+JRSOJWmo3Pl7GlbpLcSm
UZvBVKfXKbcZKW7gwRy0oSqXymZrwWwWkbBgJHrVtWjBjxSmtnOjUghkMiwx
BywDwoKPAun9vB7ggfxjj3oVFPCnn9dOnwAQPR/mWm58oT2Cez1KUTtfXUkN
HMO2sKB3HupB9+DRvnETHj7WW8kkpAPvNJlL9W/VSFZROheCe/Pr04js9vCc
tzDFv4EafDhkBjpadZmN2qLTAV0Nh1X0soW8Xtiiqveu+d2N//vnXSSUL/6h
PFbjgUVH4lcs99Eci11X6P88xbUGoEc7NZ1Dw7vUByBERlSchw4wjzXF9lux
lbCxiMA/7VXYrbQigrLVJWU/TPce2PSaNFqCjrl7Jyz/HjRpbkVWadmjKZDk
TRrDBXa/Duf3t7FCw1BOKFe8lMQxnNws79vTetEc1vQyUNdGxttNcVbmt3C8
ydjmm5mQgm5hq0ZZfDCyCyogOJxnxObO8Ze3oiCcOzuhRp/OlOMbPjYmm1m2
NBX6RqSGVz1RMqLRvoWJaqhrawbZhReWJp9HZ9qxtFzuibSET5VoBqN2LdRv
EJfCx5I9F9dpfEMAtZUO53UVOFQzpz73McSVGAuUGiMyYyC/AnJj8C4NF3Gb
v0GE1UGdSLIXexURT1BZu/SxdaVfZPCem3a4Uot706QBZYJtn4VGGpPH8QR5
qqETsfkWrNwQYRbLBwQ6npPSfCTuZ3zYeKHdZHU59j8FORwxfR0SET5wTD4s
4IiwBdG1J05tHgaQ6sS5H8EZFSxF5Dn6vWtCasEk4sAf0WCL51zAjs0Qcmi2
8HNhcQlhEuDZUs9xiO0T0Y2WjzHiWKePvyg3WNwSUMgPHbDptla9XtwLakUr
bUS6MQYg01M2pdVVTvl/pmRAQb9pjBxAosNLtAQorlpvidBXD1CmSDmkDjBE
2FNetCApnIJULJ5cVmfX/vwZZYWLJqZyF732Uf+jzm8wztGpUsQiYVXCBnJa
dTepXU1lMW+TVGxGIVZiFZtZaWsJRcUpAIFwFuY9e7PNE/bYlL5e4YA7goNk
l4Ym0qaOii5JNrjVEPf/Q2zvdwto1VvLPYJjnAyqY2q/ytAWnqPMi6W8RfVf
2Tv+N8tVVd+P0jfs2XjWP+cnrIpsnFKYzgweNy41k42kZWGOlF7dTA2dwgGS
dWWG480Z6963m/YEQWQ0DCF5GRiDLg3FB/0ehKyPgALxzc7VFYMf5GeXrPgN
3rz4ChrRof4eRBfMd5U5tag4Evvp64WA3K8xZ5yFt+1lgeGu1mIwK4kwGF05
hda8R8cYj5HL9YFW6dutq4KFC+AV1zmK9EDvtWOJvYLteZXkn61HrV9IVsoQ
mzklgy3UwV3RhbF2cfvXSchD2kO4P/KDYs/l/QdMqQwNWFd7LcacCtbOin4C
mVwP9kyW1MNq9xCC6zcz0kIk0U2lzJJmpycwZRSkTg6NhPVRPxuP7rscBawf
wnh1YQ/pGEhmLYmuqJgsVoEb/TJSxLRxX0612m2vCi9WTtgMRXOyfABi8TPH
+aSwQ2mPhZ6GwY+gZzuzmb0j20qmoy9Gi2mDCVLSVBOhxD7qrDLyswKs/pKx
aU450t6t2xkZMjWSTEpikYM/YySx40QNqxt5eF7A2recFE3aGqGVrLjxgUmR
UM6R915XG5/Jz9Ex9m/RWBEyVyDf3VIrU6JSQ4KSOwKyCXB5nmwFuR78Qvma
TVWDrPgUj+sGyOxIZ6XQuUyj/TcYdBBnOuTMrOHo1ywrnLDf5IHBYDqIzm1V
c4lQnDsve114OZp/nY2LjCaAeHuLO28jexk0Jy1c1kCtMeznMe9DMjpTnz32
T9G7aAeTkgqKO2gwj1Zdb1s4Vb63BLUB/sni7faY+XNTCbT+T8eeqtxixtn8
NNAaUnR1rdn17q4MF/94dRJyn7voG3kIAyr4R7uxS2ksREGkAdXL3E8oIG1e
za3T1OYjJEkK6EBeMCJlmVzSnZ3Z7cPT1yBKl5Ra7ONJNERFjSm27MTb3Kqd
ZCZX/POCGsUHdy85ieV2cSggmO+TkdNH2ZO5lHW8XwkTWymBbzhZ57S/aI5k
/KoA7pHkgSEgLtGwsBymctEOsFd537dIchZnIDmEnOO2qS0VnNkPobWnVTKg
jHqgNGiaQRFFBUH61Nmdqf8uRLmrMCPoxTxyH8q1bQCacCYsGfG1jiJBhMfo
WjempQD/UTPpIdNdtDLaKrP7mtZ+IkvL8PKR9DEpxTDG5dEbj7pYPQ0P/oaC
tUAvwZ9wt8ywgF5KjvfZzJMC39K849OD4oqv8sDkFBpKOmvqeymbbKLMIz2P
tFGijsZzhjFJlezGrraP7kasBNTgOL8QthCyZeiTwBq+yzVqH7PCQZoY6207
BIt3cmFCgtOXaMW5q0XpG/+ecQKtxTVP47A/JL9goyahqa7xmt0o+Gd0Pgs6
MrPS95OS8s7Of7Ib970QPACJ2ICk46M6PLGD4NqHT3ySqhJT/Cjcw3VTuZpv
9sBhkouhmRZ9QZs0AIuIBuIOlzyq6TjAJ34gL77uLBaT16zP9Ofz6clh6qnA
AIr6u6qbHU+GurWO4o2nn94CVCfNguONztjOT8KzdXFlg7iuTygXqp+zxYqs
spmTXwgm0gbpc1KaUBpqLVjfQaOdH3sXsAJXphOFVcLIK0wwESyVmUG4218A
Oe8gg5HyYCTES2EEO6zCsgKQtKgNTzrRVgjTx9BjHtczpnx9WUWDmyzFAR0r
Dt22YKT+sDzIGXgWmN6BXqfNtqUgovJWCcyNCN3RT1FaDUH9MUAEeX3XvMvM
Bh5CG3tP83JqeeMxhRnvdHtLwA5jd9qNlfF2cFhmRPU8ML+0TueiV+QzammM
LxRgOP+9rPvKLSLnGW8XouQE6R6JfY+ysB3vqB4wWSzRuKBfQjKMwT/QVK7z
QYXLnSyGW7YDImbh1zs9dS40g3jRSACJIZ/+ekUJ29BXmptb1XkSADdYEg6s
sNiGwQKhsfX9oqn48i47U39RP3iyiBAwAxTwVlDdhQqqqshNIJET1aQ6VuYD
3mS9Fg4mR7a5IDXjDKwFWB0WG/5bDV+E0y9nNsvy9zRR608M1EO9zLFYDjo4
dgQr2V8Ld19YdXQkS0/E2LdpMFJpJ7Ah0j5NjZtlFcjZA71Kj9gNibpjeEFg
mxk8+phfMON/HVPg6Y0mqa2CCcsMxMW9giIUYpQ72OSFb6tfrsm8gEaxcmql
Unp33zVKix2/RGMROkqYJOAMtbdWtOUiKg8KglNhFzyuhQJJQdYG+4rkr67b
gv8TtTkgqeTQXRofhhK2DecZOVvm/dECGVNBW93ieZqqGfvpsVw7X0YUwpVT
Uk5R/nlwVM2RmTqfHV0P5tuJhUPYCX9bBmuOvUgoThFa9u2wkNtk3rsXPhWi
Je9i8FWuoTkaMryzmURFZavYyyP8KEfmiQeFpjugJ0Rw7pdedFMFWhOWliO3
9YQT26Vno6uyo2Usf4pACZyBR7jqvmSdgCKNsbmnuuZsSBJRhPJdJ0PwrGhp
lGpf6Ny6f7vUAy0qzrPOEFQAbrcynlEfB+Unn0xERAwVOSpEre43Zpv0oRrf
t+x2KosbrsvHPwDMXxUWUsi/8KBOEMVobXtRr3Mf2T2PNrncdmpd2cssBlt9
vonCIbs2YZVAHTv9fU3eilwUDXYDdpZq7oKjqXUojn5lH0nqOtwqp16H81zt
Rpe0cR4C6SjocZQnLnXTUC37cduy6qoveGHVyo1CiRVoo67S0cmgVdxzY5p3
ImgaDFKSnKZMb63p1pZDHFgOcdF6g71NylYNWOwnzb6lnP6KOHOBAYdIi1QZ
rbfapLRAa9QXVhpjcgIpiAR9Hx7wQLb9qlv/7g5/39UqKOsE40o+B+GgU2vB
hhRRtPzGgki5kb7SmbmwbZ5iSXqmEcww6XqshL/xqDZ13q3f8UcrnLZNaOUP
5i3WtzrP17LPHOt36mPtkbdEvVprxiVOtYFeq8As9+6wtSa8HY8a6aPN28+s
Lvxnbv/Nt4V1BS3KsJ29J+n4s+YdHVI+gug/RYDSvOtB2byr2UtetXkszeKA
g1RtnYBab0sKzIqQsAIOAPgPg/2Q/wvfP+eIN+QLoGwWsqg1wjGemkhUR+f5
+YcOIUMLwWUnDD9bEzTajmeYSR2rEP9uufWDN1qKGl1gl7JqNwl0Dv4kkrew
64YMhvsteG70uDo1gE/FmDzXvAmBLrjgV7eMi3dMjkNkgOWcTJYeb7JjgHFs
hVUhUndHSxfMoIzewSfwUwGyXf8CKFGEpTvEy0AUQNkcyB6mAJhNMUa4SB+7
RJrpS/a8y7dlz93H57lwhEH6XqYOo8RMAInUKRDQVvgoAjeV12zNaeixJJsL
9pfmX4l9/3BpQw+AfulMW0fB1gf6WYnq33FCCvc7kAr7MbkVokGWqTJxOxNC
Ljy/IuHf4b3pZfPfM5hDCdi7mfcno6sbH8Lf5wP6NJ5A+qABdYyeZGzWgXCe
p08wZMDKpVp/S6wUD2MovXOxp7O1iyDDhKMkE7+c5y5ts1ibMugU811PGUk/
Z7ku49oF8Ivo0EjbKtTC+Wbi1963iA0KJ1aJC11KksvQoA2u/Ph5BBFLJ3u8
Mf4BYRD9V3KE+/WITXnb95SAXv89py5ehi0cRCDZlSh05q4hhqMhyHT3GhLi
tZrqLkMqmQ5+jAERVTBtOiCbOWIwKUkg0gkH+utYyqSsROy9ENOaQ6w4yDYn
8pkpTTFkErT7dwwykretIE0Lzy6FcaR6zj4ls5MsO5o6WsdO3pY+EDQJRq4l
ApkOVAGScZyxsa11zMoEt9ZiEHkYTMqEhnJgXWCtYdMxZVIYMwVa3mqfpwMm
wyZy+nBf+yub+AZwo6OpWqwNdxEwk7AIwwY6VEEeIGCD/YkVHE1u4xH1ylbC
DNnNOugNmwuaLyEkU97m3ZF+UGy+0XRLJMQXXBP6m7S9d2F5X+Zo+mKQtOE9
Moa4N7iIT/7BMMWKbKYzpy3gmO+SKNngNZEZZY6bHgpudNwZVpqdBipCi+P2
GT/hCdNdMb6TwcnlLCkujzHWzyge8qO9oc/U/QLPEYcTuAKewfss4lMj236l
gw/yP8UmtpsnNrBUUEGBKauhvbi4FMSMJq9ZoUwNxVp8QhTSNy8rnVtqaWj4
XTT53nmKGHfaArrD0eF+tO1eFj1uz588X3VQgr6FIhhO2aQFTadrOSE8ev2Q
uyHslCrLXFilA8aFof/OUi5xdWqRpOxyqGNaiZ84b5qemkw2hzE0K7PNkoQv
URobbnR/BmVQRI7LDYC3L2tTs49+ACeZQyFSw6En4D55SOt+JPBpIY1r1X2y
s2FGX7C6kH0h9GVV/WdCh8/XGcEQPL53mYmvWRcBObkt+L3G16jTcInJhUHf
utDos8b7GkIbEvuhK74KoV+D3yJ+ZCriN59o9TJnVgqpOUPAC1cdQ9in/+HP
j99p+tdUaKvpb510m2Knkf0/4Yn5BDRNXxMa2xCXyMdxwpJ2cThiOBylidgn
dvy0Ygrp7xw8PopE6vQvD1lApOoqlrFvfK9Z4nODrSoojsULB6LceBIuHoYI
iQgMN0nAzBw7VUbyeh4VImW+auyg9x7JscWbeiSs5u2DZaSw8J9nydT6wWHr
pL7+0ckuZiY935dBU0KCiLGSq9BOAAZ7L0852u1knXZ+1enwh6DIby35k13B
7bR3nbg7Qck6L/w0bcg6t+F+9LK+7P04utJoOL9YfR/NXVtFWgbhtE/DTd9e
5lCmoZUzoSl7NmSN9McMS2kuCM4dIsc19Sypwj/dHq22nWblWhuGNylmEmQA
+R7HwPqpDRbdiV4b8hCztdZ6Ag7R25wiS/QIZ4r8Vt21MGPygBpG8Q8jzk6L
t8WxJSfec/a2m2UUJz9ZBUcQxTEl7hRXaOuLC0Xp7xdRH9keIaqZEzN4yrES
S2K27JMcnBSRn+tZQ5Q/NBdFeACWYAB9DzpOnkNMR7B00Qm96YlORjbaEIQN
9GHoR+GYobXhZJqHwjjR49Y08VRuHDab+hzdEXfoHoqsHzXKVu+71X6F6YxT
q0iju6RGhczCMMn18xLCNU+VquBLNNSH92ekptLfjiWR+MxhxPQ79lLElWP3
ffooAEHwER8Ui9ckEmO0GbqdKsU+TySYTvJerCXR7K0IDjk/CejZm0IXRb8W
w+VYrSzWenbWW08+L2S2t/bLkuLPBV3U07cSm3KaAgyzw0fYwRWRoJ1Vront
Wbz0aNgAQ8/g5ZvOh42igPt7/u4X03jGc6Lbp6bnIDuTMwneWhipLkTM27PS
TSGAt4ud2vLmf2Apz+qPsHUTwWVeHZPMgFzdKRvmE+5kEkQMYh25SMmm/18L
14x+LxzaJMvPacfBIZpESSGpnIilM0zj3Or/nI4QzqqaYjQeB3Dfk4PKXZxV
BcK6BIz2bVZCtccktY8PLHMs44SEh3EE/GTiq4J2Hspie8PfWKz/r0lQHwvM
Gn3uPiMRRAR+2Hb5kMqC8ojgtpnp5P+N41Hn3CmeiMqdMqd+VUUrJKXZnUrI
EV4HZfkacMakfdY/tJRAgb1sAg9TZgMP7GU2nGUl+d1ARXbIJThHC2b87X7M
GohhUwE1z5O38VvVTk8Ckuhz674eN2kJQlf7CNh3N2JvWGtSB0+aRbYyw8Zm
wdFzLVD0XHTxeRK3uf0R1J2J9fjv7KQEzv2faTizYzcNgrkGGoUDO1Yww4R8
MpnzQ3YPkFGc9bLs/YfDQtaMDYBbjhZwCzIASpZ6+D+nTCCHAYD9KusD1jmj
cO6EedyxdHup+CmMhsAp6vi5J4u7ljqXXAvhLbTChqDwcQrbjdAK8PYRRcuS
hBOwNOu1PPvwk961pqwllvO6PW5cp+5Vo14GT40eJhXyvDikMZ0Yl4o16mf9
+tepGCre5gnDe0oz816oKqus64zf3QOiJjE5yRE8LZdiP/EBOWkACJCir8Zw
Pwj6cD2h3CFIKxhYlLQSo4ArtPvZeEXNh/0axfrPEcTlYyqV8Uismzd98c8o
XWaj6kYsHxi6zAUGJK8YRzN/KANilvwnLxQbxggxmB7IZDFNIDV/+8uCalg9
fE9x2RcmSdj3uMwGjZrI9855CrWoQskrRF3bQc3KSW2cjDT2ZWDgNKfcxyG7
HkC0IT+n5pTMQFVwCo7suWFWnGCe5w6rwcwLBcIVKYqexoo2TjcNnE5TsQhP
0XAzj0gdSpMT2AguxIX+whsiew2W2TmxcTPciHyU0ixRXDA5RBJ5JDeQa0vW
nWhlHhqW4evrRfOZptUjy20IZo0wg8hZ/xiKMXHW5EmkiIVQuA8XvFU5mu+s
X4zz7KRGeU5BF8r6f5SX7XrZyUXlM7UYVwqs8i2c5ipiL3r8/7hSwcjbzcGR
1cBN0CMsA2qeyTFSphQbCFI3ubQeB0kTNTI/dsCH0CtdJ0tjgXITNMvOhzAw
JIazGUXyUOLWgYXBKvf+GyRtUAP5w4f2Tmr+ngUf4Oh3zo3AGkViUG9QlV8m
oWQBA0TDMKqm1RZqQPlIgm2IcA2niLy+2re67l3rQ863LtGgyWgDW6lV4DBi
c1hK679F153Guw44+q5lD0M/+VkaLAxrI8hlEEanEfmOvyWpGXjP+SDbVgIr
Zi7+cxk7eqWIjM/drPiwiqZRF/55ZW25VGfheTTZCwMhSeenx3u3kUq9ywHw
6VJ9NNF9AEXDr0dAW2fLY6H8ad/4uIPBLn9uhtwIpH/nLU1TVtP/dJuTcqTJ
yS28NphXI8T3W4Ek6wEas2fCkxiGAB0V6iq9AtSyHftq8duD0ILLho2e6Dku
Et1CZnNZ4m/ooe7n5QLuuq1pI/li3meTnRlJxhR9y1wcMzBCD9Idn1Ljts+a
HhTDhXR/H0LJ8AG8eqXdUz+2eVxguhpLG2P9Q3RecUoNZW9cEHMgXfGfjZZh
X/QXzWrXrR7h4S9IFNQI0VuQLe+3pD4x3kPjAleB8gAekQNyrHACGLwhBn4T
GDRbYQgzCwy//Mi3enroUieUOR1Ac/ehB++e5PwkllvE5Y5VezorAwyewO/g
iVgn/Qiaz6cpPM7cXyMNYiM+LKdv9KKoX01pH6j4ArbA9SCXl7R3W6qsgQ2L
HyFg1NclMCSJz3aHvm5JLJyBDsdDtxUGfeIojph+HoHMfSgkY5ADDmJtwOqI
ad8xUwxxQ3/F5NuOG8CSUH3cJV2EE2qGH+bQEFsviO4BzMcWKOsYmzJfrQ0G
lpkNenjBlH6J6u93v8YpFhp95LUBAgPAVQ93+GwMovc1DE3WEP8G+0EGyqfX
8U48NHEPIgfWHBU99XerJ7Ujp0RCLI68V/jBAGNtaqf+UUqYLAnC/J1+zhiE
ZLaWAyHJPI7V4ogB0Nf8X1bp0TuH8+yuo9o1sQC54MPtXeeTr7JiWqIlQph6
1RxtgTqD9jcL1JW8m25bNjotbVoEX5/ioedPguQpxuzWs049aiDsbZ+jPlpU
MGg7lI7s9tB5E+rJNa3Ye5VBnAOtsOBukiSCdmbFylawjpTFSOHr0ke6ZC8Q
RbYUF8ae+6TFphesLfHSvQeafIF9cNNE5yPFVSxJX3xIMTbwJO9QnLgdbqH/
kNRK5hZTEWXCAgJBOM1RdaYdyVs0+vROZa+EiYIp5IwqTJsWcrnyxaQmAGcA
RgyELYPwzMv9ZTcHUC/BLyTo6f5BTi8OtZ+jIw8rOme6jyhE8XLaTDJnZQX3
cJ7MSMGPFJHhoZTz7Lf1eDcY1bkSf5sW1+bLiwZwv8iY9zyidm4GsFokZyrp
iHEbILQTpnyuQQ1vCC71gLp1N1UlumABeCT1RpI0jWJ6OKNraj2+3xOdDfYF
tLRAo6WQUNvNocL6mP0BGSSkr5SZT+I2+yJn/6SHq27yuQf/t0w63JENwyCQ
PeqBoi359vxIMB3NhuObhPSN80Y5gM+pi4wzi5cWrXO8fTi3eTSAHuN0/vyJ
qHWIfBdnREtk82v1eZbkJom7DinR1wXp4d5TvDz4b8trBKtBNakNfN/nzKS/
Z/tn6/+4ZR9b2+eMZUEtzChbmz3RAnG2JG3olWk6lKRF0bs6LKo/GtZgcbax
E5eL8rp8i9Y6eDaGlqyfRTZXHTh/g1Ix//mUUl7y7F2YqcfQ8ty6bzJbgDjH
uNR4FzK2Sv0VYM2OUznTqzxOAOpgaHTXLX7IHmg81S6vz1IObFC2mW1tNAxg
jruv2iIoh/8/VWPZMLv7rYQ3IL94CZYf+yHDnFRTi7LEV2mTNabGyEQrGwSt
OLQCQBBy2Stdparh5ockGLQvA6NqoSuYm2bkSPhfHm6DBmOht9C4SjSdFPvi
hv3GjPHy/sr6asAinD7ozkIum+NExVz/FA4hSpnZZryx/cDKsC4o9wbWS4Sh
Fy/yCGjpOZ5ih4Ct7/mHQTqeZJdcQk6sYIn2CekrNJ7ARd+pHUwv5eal0bUi
4w2T31ndVpmgV/obyL0fbje7UOlOuPuRwr3Fz/WxYFP7jD6ZwfASjPHL5iYj
GV0C51cRW3KfqvBsXRoEdJ/yHlh6xwczGuCkZa3IczGrrnUsF1GWSDLwpX7N
WhcZBZM0qpY3Km9pz4q6l3cm+exHbKJLYtmedPBUmDjQk0w5FSL+1UGy3XAU
RLnuujqHYXW+jKCNnOa8If2K00tVBrwQPWhnWS0uniJwwrj4iUwfkmNQxWuo
Qck4R8jpYeJqA8OpupCXVwQ4HcMhQy8M3RySmevzFJizoRLHHOBNx2L69F/D
K9Fv6/VjHlEd2rvxd0Z3hKYS0/HoMFSoGtzRMebF2P8h6grT7nYd51fLEYAH
PCVnBaNYmV0C6C2/ZJQoYCiE9yZL06JyOazR3kbNcPmJIvGt4JyXm9kaB8yP
u3VUf8vc7rT8O6v9LW8r/UvY89T8fVIY2/QHnpbZDd0MrijRVw4T4D/JgB8C
Nv6QXrsJBptTgC5hmUt4mZZypJP2THRZiQGCvxFHLLMDD3JBhAiPg6+lSy1F
KtKCOCl7Pf+TI2WFcTVaPjSsm4i7vTXnh+pSLkK3ZCUl7axUlyMGwU7uMtUD
CRo6eAns7QxF37SfKtQAoVj0DsjGsUCeW8F4gELL+NgN9Vt22SQjR34NLRZ+
NAtJyuSZ415jjXxA7SKQ0l5Uow1vW4p2G3zvNfFSdTJpRiUDO+GLp9sAw9vA
GXnXoXwOoZGMuwhgLC3gdfzKf0pGMbvNOTs5JuOn6MaAzqpwGDVfMELC9ZgK
5RV/sayh24Ar3nEywLScy3Hb1QxUv61dNCxuzbtMA1gZOJcHZCWzDPIYXHB2
1SJL8b24xh8fPdn+Z8yJLiJWwKW34vH9ONz25nlaa1F2I75k4Z+HWzFu8gn3
TdhX/7YStKvpwbwYcNN31k52jQOWV1Yg/6CIJjddSG/3YxEaLCAGNSB9/T0U
0Guz55mkoUiPytLuMHYjkK/nyvD4t/er6mcZTo56JwTp+KHOM1UgzzJvTf4O
RF3U9qXQxonVjawwRpNeMV8T9ZKSobWz1cMx38/Nsxpf2aAKabRSK+lQaFju
r69EC6Y3wsJrdSTyXL+7yhERht2WItItkMvgaOM7bLM0XpAxwY0bens0LR0A
3Z1qP4J7JcWeP65DiEVJofMnHnEkyQO4+W4reYwKLPZDIB5AUl94kCwJ6oop
FfhAe3iP9ZWnrEJRCPT5OSxdm/CTweWn7lCm2FrW8hCS4MjLKhOaCsk99EQ/
wu2krAcl2mSf6N+BHvZiO7FvVG/MgKL+ux+JjGI6R7QSi5p5yW28fAp4gRhS
HHKzRdGjImR2s3RJ8g1K6nhB9nosJmmiAiONfnah47wWO20VwTxsPhvdkTza
vvAzo+kXSl4/suAw+R5CojVTPr/Py3hsMSmiZgAh4jg2l7iRYnxQ/9YFH7Zf
IkAS9vHQ1sXXFifRN5EKh0wBb1XnyFuOhVgEcZ7D5P0nAXCEcvdXeQIa3WNJ
YLCq+4XNH3ioznD7OhuA8iPOFdMkHMVbtW0psl/xDoCSIzd+iuh3BUUxn3ql
ue6cL6v8+h01VkxwyJWuR/RQl5ESKiTom6G2n8ry1SHwiryxtR+s5h7Fr/Qb
RCwRfYCqk9/UUDdLuFw+aVH0PunhtZ1q8vOg2urjyBk38lb2X+etP3tBB1Xs
qFm6fRpcA351EweC3USQf33/Gg3vPgX1jdKHcgRSgKw21Syl0an1PcY90s0D
oPgY0mk8S4zxWgTI4filpU4rccbCfDOxXg67ui7odK4dWEc9+loQPElvDL+A
9Al7WrfMv2oBruCZnU8k6iCpYSWNlOzi7gDNxNe7Ll1MPLUhInveeZ9DPsrx
/+RIaHetQSyXACN5CKD+r3axG0G75W2YkmHo6Ts641xF+JhLg2/TEZzZVl0r
EOgBe9JOC/Fz10FYsiXxYZxHm4yHYxtqLgypWbwhLckyWWSeJn9ANB0MVkdZ
SaScaYOI4usNIyfdEdvIBvIMS2WyAA8Y6wffHxiQvkU5oVdXkLCFQI7eYjEH
TuQK3kZVGidc48W/8iWtqjsxgiSAUw3rZfe9nuTuX0lCUeEZGpZTBnNsCNjI
rzCP2YDwlrn0g9rD8nMaksgtfZir/Xuw0g1VzCoFOMqGwZmcdeABE4uUSLUM
wbpqnPnJbKfpa4G80L37s3VKnV3e+Jl/NsltKBr9XvyYhVuWQEwLuUPtiQzT
ayN9Y/Kl+i0ls4+JcsnjBljNfcm/c4gYIZMVXwpqQTrzXHNvh3xvUKXaV+pj
PiTiFp4Qb6kuqVK/vIrC0J9SqUyIl6w6lpz6CVo9MYNs5nj7eUh8mcgili6A
Nn21QYfzkrCRuJYbuVw2IUqiojbL+QF4kWjbO0j9leDCHa0SVvpBHqpJYQmn
A3IQJSpeNTrZotH97pO7MuKxqkJZGqktdiagZNcL7ro0gDBsiebnPIiot7eQ
ghhNJsR3JdvatVeRst7AfShLMciY9Wl995eJ9EGkv/Dgs9bGJa7rJrnXqZCj
tzkpYOG0W2QfMoF592Le/LpDti3iPFiNIlaBMzv3Z8Era0jfT9H+4PAsccvI
gt0blCs1BA/9NcwJLiS7Tc8Xjc18gw8pm4Odb2kvtDMN/b+WOtyXgTUjYgDw
GLVzyNxtMHkt8AXQtNOES/xoutw1AF1p2GY4YE4/g2vMoqtopmtCGyTxHQHH
xjnY5pteyJoDM8Fg0OUQuHvzOs7XpdTNtT2IzY4t2VMEztwOMmflA27F9MqO
aa/Q3cNSQVSMfqXxmAfc1wf8SvgBTwnhMYRhIZddxCdYVXkm6rTrTtp1tUSn
1k616xQ/3Q8syqv9LVQZlpLOdidILIuYZb+rHisvGMuudv3axNntbDLlxrs6
xMP/fEkxkzh5x14HbZE7yMzI5SFVok9FlkXzaVJ38zxdkLcqMTnoDUpCdZIN
9+/DCd/HzXUuzAzLUsRrnZbsRqNl6yPpdEYb3FXSo8l/D6Y/VwnyPuQW2Vjz
FFRRt/+fSMZnj+hzbY/eOlz7ktJi+1uynRUGypjPcE5mDETYpt1xvMM+daNv
psLMM9P+91/EbXi76TgVKLCfTFUflyR2M8VjRKI/2KuLvSaY/IzDSEbwJh+H
funHtcvhVo2BKWaA2g4MpPlfrY+97Sjck/Y4yajt2qcz6qjfmoVqUjoUeKfZ
ysQtJhVpJiLo/Pvv+Xlha/9PqShYqfSSPCFTNjQvWY/3yOQH9saJgMVrK56m
eRzt8GKWp0HNL8lwEhKP0wtU3uwJGus4uIZBeu732cIpQ66N5GTGkZhhNieL
HLpTMSsb+4fLy+E4JMjujmawknrRUrMGbtEUXErhAaoy7h6MsLd5fEs4WygN
P+SdCTrh7DqO1ebKNHUb/Kxoq/UA3PEena7Bjhh/ycybUaGtD89iAVC1Hf+e
Ijg8Oi7V59fGYx8MfGB0UR5Sj1Bs33Q4/Wf8Hcu+n5sp04LIIAfQmuEoewbc
L0t58TnKyaJChVObtHGc1CDGpm8Gp/NwGz2tZKYIdeW9KR56N1HtUYIYijwt
axgSYnXx46m5lUXNwT3UfUYgg43PW1Qq71Socpbt+0SehpaVKctdWdq6hj1c
l3ooSS1n9vhW5DIbUA7kIGmkHE6l17K5FqlUJDbvvywqWOyXbSUPYecLaRJz
aiiOG3BsyixGZehS+NDQHig1zBdMnryJu8cJuIB7pW0HPIeyDqmz7nhI+zz/
/tgl/EHiyvx1VxLXdPdSluI82Cguza8IefhYnes2nvXBArLE2VbU5GAOM6xn
xhz309HHvUKtn9CrxVx8kSjvubIhNB+qEOzx23OyVp2934lFyqZ0Lyf60/iS
1vQhfBjnNGJF4HvV3LhvgEf6nK2OcAeQc0AkRfyFcI1ZDAsOQU5aud9fSTHR
F5pSR7mHUIw9mmpExuxlmWaW6wtJdaaGmA5PzRrbsYZu/ymjQxfh/62ommJ1
EsRGnki2LjyHE0VqB9+ZiigO9GqtbABXbltcx6q3onA1F5FlspCZ5EB0VCiU
qO/cP/tSH+1UISoLeFUgfzGYcPpAQZRqropcUFqbYZ2r1xIemJN8BkJcCtQJ
c3P1YZ5JDaCQRryPS+l3dqk1nj0jr/2Q6S4IHPm4DmpJoBvyEDVRFYXrqIsW
x1srz2/gGPSFoZrDJxFW8XvjtSgAt6WQI1dWG/36WfuwwfitVUXPFHrlqs+g
3PdyhN4X9xeCQnmoem9gxLlphVXKh5MjXYM/zRekUXbrGHKdnAa6fjWea9MC
D+veS9Pc/HgHZKAF/m53lnp7G6Y7lZoCHwI1w+H5lhzKSkcbforQZc7o2e43
FhjaBm/A0GRAzhG3wDBqp9wprIaqnCyH+n4laJz5ySCP8mamjYX6WqSuyUIS
CFeF9X8YB+5/IGdonTZWLaUbiudDiBagcS/IlrU0IV6mLPy55tL81O5+FTuH
ddBHpNOeUUv6cocChCUJePBB96pMY7Lfl6rVmeOlr+sNkPpC+Xo7ORSzcWFG
ZAo7qgQygVCLEHLx6DqPpOoFGWGRJQG/wj5WZO8MwOfPB1faNxlLn1BYcfH0
S8Li1djQhmZth+TxcNM/W/uJtqejfIarYQWLP3bzwsv+3REu1zOX6L3fCyGv
4OZpQFg4js/0YFA+ptcmPsNX8XvFwhE+ceCToOkDKY3l8/cKrstQ6G1LuJ5A
QuOSXNdTde4p1zFoBM9xRgytPuxzp1EvtIml8Ve6JfmO0ryFq7L0FlF2gBKE
rdf6C92A04QkjiutW7kJjctEurmFoT0m7jxwIEPsdo9Lg1LRVrsBicrjnqpb
z21mrI2wh1etl6LIq8DBkUtFmS7a8mQfqZf+5WivGvFk3a5S3s234PYuOi5+
ib9Sx0JGUEdFsj+7pw/CKSMMd9fKO/mIdDc+631uqI4JH2zl5FgEHN76Ru17
nLu5l27DuJwbDJlAPTqtpT2KFR+JhPhjeWPQeZk2LTQN5If/kaoMEH567HCq
RtyR6i6yDfRGeKo/gC5atfIgVgVEFmSC9jmvlLe8oOzvJHMVNONrY5BE5uuT
CSnKP2ySeoyJOfdsn4Gr//+xxgKhxSE/NNV2aJ8vaqqP41vrbS6JeB+dBM58
F4TqAMAVnqOzeAw+ePasQ5vOn2BdFKSxFqcJlC9SBCtK+F3adVqaJpwNr4YE
ocSsNfASCJHVdMgYAb7tBgiL+XWmUKVAlOeyrPMdn707dfHJF6181J1LiZyn
i4Y6IpZgYp3CCqmhRv6nk3xv5WuBT9ZZKfyR2IR+qlvbGXYMeideFneknTl6
UUik4XV/BOvyOnq7cnkH3mh1V2gYUzRPiTJuZR3Xu4qONqhjtTR5eoN/S7mC
qEyqJnslOUSX05+H0pYV6Y/xLX5oAgoVYnBtgZAtL7V65jqizaZycL8n8EzN
FlapjKD/oDSyyA1ZVmyIIHMS5xZlkgFeOJi1uBHMbVpEOb8mkJjJi5eVOWAf
ikBBM2Wc6LOKGtv150akZLGJ/hFLyJJGEqvB5w4slKQjT/sEEpMrq0qOU5ab
CykloWKq24ExlFEzPy7ODlLmBgK9cl6teuJXM8LwlbDQfJksqK6ifLebjO09
jC3NB0NjTsJoQWL2jyaccXHLQuV+J1rpdO4RjLjH3j9oH4bazs3EpwmDw4vB
UHqnuSWFc0PGqUuEtajIg016pJPY8ov6F5ci+xEeN3JY17HwPRYAW153F/Hg
XwBx5y6CmGokqkxnV9VBkrflLzGwMa0q5krDu4cNzxY2JhuerjnGkvI/QfaU
0EsfWwaKC2WCybzcQxC7yf0Y1vQrUOlyxtstYPBjGcC8W2A7+wuIE28Wj1rM
YH5Z2xO6dbbKs1td9fQal6kE4vL0EdGpTwJ8RdOBQRUiFPo2DmLvg0jj/KdO
xtzljz+/D64Cv+TDxzEApqm564wi5He3m62YOn+cKVHpz8BcE8+9ohICOlNO
o2hJlCeD0S6uzUBuOBZZJ/B7hLdYJvOMAT+qnEX+A93Pc+aaP8VgU9IpiFXR
SDcpxPvwzAtfFAESDB/Q92wtJdQWVDYKsWS4sK2r9l5gjhmbAuDT/vnYF3Mg
iiXMjX5TJFAcHgLRubdh6oydwgoUf2HPy+HorQNT8/+9MluobS6g359hbAx+
OyZRfRnOa0Wfik3L7E62QPsfFBEt6WuHhRu0Aw5EAUyXGWH1CLzwODlXuLIN
i6WFu+XmzLN24GZLRjKs/19VIpnNs0q4j5hPI/1ziZe+TBBbJaLkEjSOofZg
q52dAfvrJPWK3uanwEx6+RkYaij4U/GNqhLvT9xVmb5089i7J4IZe63yi8cr
6yrwt/GNiG3gKHLe1Pr5mmGZuPs/TENu2R8yttQdtAQTxH5lpqf1Lb8G9wFI
Z6Go0h5R9ptMGG5wtOpF/fHaepodTvG5DQvQ0T39tW9gsqatquK45u6M9HoG
M1Rr5j+f8X8dWGZc9HwDSw/XuOnOOHoJGeF15i8zVhQ0ggqr/lZudXCxjjVo
lKtktVBBCR1xa87tLJpzP92p4OGh5DuLNRWCgEPx8P1JFQc+cY1omP+0eoDb
OUHlcFlv/poSHZWHu3Jht9nKFHRU2JsunTJRXvZSro83EfZgEbdz15zeVOBQ
pTgsDNnt/psZhDcX4tQDZ846DR92F8mdti+DQ5i51zvQdeR+sc9Z1vkH+nsx
NzIExYh/df2ZyaAqZuFJNvuJ0CH4LUaMMrokQZ799WOrTzxpGzYXfRcAbx3t
Ok4daNZir0UBBHzDL4YtP/qWsJd6kmHVED9FvTtrWqChmUn1ofc8sQXo3sjS
u32qnWFNtYoJNC0MC+Cz9nI3O3fib5tit43Y8SM0+xV7h+ZljmUUFdRLs0EY
bDq/gVOoEZzRG1b7TSuVciyVYwHFfczZQ4ZzsQrg7+P/eB2cjDrS5+UnA7eH
MPQh476r29g6qzCLiNEyiV6a3woUzyVfhP9sAPa74T9xpJxPbRiuUSikUMVj
pJNvbrUF9KCPVvKGeWQBNGFF15qEd1IHsp3pKtSTBkQHDqC9u99xaqRQy3FO
dhPjUWMDi6XYtGY467G+k/2a+/0otoOxLr65EUQq3N/9a8yP97ON5N0WPMNA
mlaEJUUIJiegTKCOIgseAxGI+ci40f3SAQ5KfNcM4KAPu/87zslAZPfKsJDa
Z+XceZ8Q80NdYT1M1GySA9QgRSXbOWlIFEkC7ziSHmcYT1/oE7qQ0YOVnqk2
oJrMmJ3NhgKqn+YYx6SMZQhRsbet/9HGJe2anBcR91a0RihbdxngzyZlfro5
fILwRACJS9ACxIxuWYwa3deAkK70PH+gEHHIBeLPaus6pCTos2svLx2gRuvY
pzJyJ+vKcN/rMVvTRU7lIz0i2qBLgHqWYqYyiW6ipQYhxLH9/OBYU32lGtpu
Nc2J0Iz1i2b0W/bSlE4uaUo09rZJXdJc+nxi82JpG3c7tVUHfvbjZNZ3k26S
oEg3BVp1C5kpLmnRyCQXFxp4JdaiYo4QM4mULKXiqDLGefsoT1xFG5UMtB7h
HuqzEVzUUk4bZUw8zBn6DLWCRfBuxHFxk6F8vs4EhOwMN5Jl6FWpq4JwPpa3
j6uUCjHxP2IpUzja/GJJ6svnj8iQHcjbsWv+VGpX+LUXgrQffnXjPLE/LqgR
bzlwW7+v2krMhtV0ytZd98Sh+4qT20Jo63rHkWmkDXZj188P2duv1PhfBhDb
D9yzZOUx7gKKb/kPvODydtXFNUqjS/7pYJolw1W39YAznG1YSSnprXHQFUHT
9GXj31yHlP4PD1VfPowNwNO/ERiD/8BO2JeeL9CjzF9kzxao4EXzihRwGX5G
7WL1cTxqPqg2kYGNMrd7hpvOxk23I05/q4QJERfHS+HvJXS9GsMHP2vXbPTM
wtN7CG76AFOJoKRY3HbMfFsyswsATdBVPn3/V98iqf9OmFsiT1e+wD/36ElJ
QSLUoH1t+9FA3P0ReDDb48ZqNS9n7Mua5TiZhYukQdZfzfvCwcmeCBaTao9h
9XtKXZ/pmxCKVIxNjpFVrfUeFfZ4iuZoqC9F1+Yz9fSoJMcHi73PCUTEvhJv
IsHuQEN0gfIKyRdn1D6GGSN0XakIJWmLa8dcHj13gYS31th1rHPVlEwcePUy
W/I4409QS/Xljb4x/FLTkTlXvLKvj5xWpbd6RC9EKT7YASOsV67pBq1IQ7ra
J57ZsgKcbehxOeasLv84Kepafd3Qx+gVizn+lRt0/o8fTPSNoKb/dqCDevdG
F0zJglyjLVA4gS9onuxpeqwUyZTCFiYraHiqhsp0aZdvzlCksbJp+U3QkuzI
HSVQbpNsvWTi9PPvHDwu6BhVfQy6pTWXQNsXWEEbfFdKPcmJtTZQk1O/6/zk
ubbeYfVY2sj9JTimcM0zd27ytDYPTWAu5INXMjSTxJJTwyzKzIKvByK7NaQY
2Kze8GX0EIuwCfgJd4GDFRc0WhYUwvPEtTC6WuLsPu6GapEZzfI3PZ+qVO75
9tZ7RDS+k4Cpt3IPC2wcjz9JeUIHk26xDhE4VlhVoFOe8RE56fD0ZR5wADdk
DhIalvy1i4qZw/BtfuIPQbSohSUExgHprn4jD3IRYoUfb+HvtuBM0fWoVmv4
8QaC83cc6emg8AWXhdXpXjh/ucgFfCzvgee9SvD6v9T85ERUZfNu8aT+SlGo
RkGl30URnYo631og+03zKLASMpdyoWOjeIUfOEz02ds+hkwHKar84gVpHiZo
e+RMUsz/QV64gCHnG1ueFMqaaROy7lXz/iRq2SDnfJbQnQLLUJUkCYje+pYi
xby3Q9UfMRc7GhMb8eC1G/z7d8s4ViOZw9YT1P1vl/HEg794HZeHVA3tgCJH
WwzXaDfFJtsPPIdh4iIeDnby/hnzuCy+unK1DiLyyOBMznhNWHW0D9367uYq
xGoPiRHbJ5KM0w1RnnKB/SGQtuvpu0+e5V0hS8GvffL9wPszfVCdw7G2ce2/
+waHT6C+K1+AetP1oFSiBkVa0oPQ06pxwdHb9+7TlAgWVflZc1R1TFv8zXsw
/+keFnEYBXW+P1ULUdiIk1fqaqh0V+fWob5YYMh/tNuYc/0+Pl3uR+NwGanz
N/I6jLz3sWrju96tLRYkcfXgU5WA1mXoSMRgbfRsXdTdxKZZusLG1iugVdkN
+y7M5UEeWix7/lNx2prC5Ildh+dfYWQ9W8J+/kiADG2hd1TqbEncdDYX8UFl
zZWumfGkaaIJOFW+wRs1LUnlXGlMoWRn34G8otdDaaJTCufTyR0lprlaGq1G
xTO29MtSo02MEnI60CNnJXscR3hFL3Q1fLxdxG/MhDqsuoc6Q0cW/yzpmcSb
UIqzt1A8+2ahqLZ7TfWlIB7aiZGqUiaBQKE5gHTLNFTUGA2XcF9U0/qEeS3t
QREqSewr2UMJFeWPGHx6Nh+ZOH7SqmAKgjtIixMGVx7d0zs1HpxR5GJxn5G2
XSl5FYqrNzsnBbqhdoBs2HY68CtS8G8jaRLtgmV0bFGUjUniSvlUO9UX5k1u
DdO7/YKWnT50+7g0MbY8lxbmLeWspJCh/VJF04nJSf/yKid/wUBUB8LpLWpJ
9jDQPIxptL4n7YbtKSVwdddEC63FEKZ1zFEyy2wXOFWiCtPcK521ZM2biddH
uUfIprstxhBBcbgJt3XWxivW1vvPXS0Ca8CeC6Dt7fBLxNenQCUqfffXVxem
9I99y/JwxBNHcjUDXCqkQCEL4p4z+hQarTqviywqizS3TF7n0lZ+QZR5AE5M
QQIFvyvykPcFIFkDEYfc4oyV0u5W0PWe1oZKEi8Fu53LfGzPZ8iG5l1znsTm
bHeW6hjfob4S2pkhMi8nXVdlROQFyPYTyeA3odReb6yBB2xmE8ryq+boOwGa
x2l6VJvVA8yNCpF0acHBsMfCBv6wy75HccJCNH8azEydG1k9OncRLvgbFAYV
6OYBKJEfz4I1JImIsWOsAGRk2v5Q7ITUt46KzHHorcXyj1n8qCoRPFFEBi+s
1W7Luh3pd8N20sTdi6YaHxggTaNgl9P1VEOHFdbjirh5apVpI0iCQ7Dqwpym
cviIvdSgW+8aDIATD5867R0ndDBfHIJy3Asi+FDGmq5WqZbVB7no3f2EU0n2
yyJ4vFS0JB9ZcEYRRtAfGdzY6JIeaayFLvtwhwQbfNVC1WIpXRd0xvzuyfW4
FsyJQqXLjADkFp6V3oRF8KweJG6V9tlPiUZxk4xQKLWNFNIiq9eApWOl1A4D
ZtKoUknV+5VGz0zUgWzlMduSUyF3C9q0Zel17rujfT6X3sncy1MgNFisQjk3
xU9wQXGBEFm79PJXZvXA53IPlrZv4SY3ZdtGvLcIFYqd2bId7XA0V6HczH48
Bo7XAAIvrgd1wG97pwJv0oYe/K0G2YiCjozlOc0otsZOKmmJ8pPnnhag1HOd
cPG2Y0WJWJ+L2SDab3T5GfsIk9yAiydn6Bh7H33++5eauGOqyLJY0QR6mjhY
q1tOPZAW0rzLmy55iqyUOZCw0UId5ECXOpt4AUxrNglLyvKap6HV+RcY1A3U
YiCwdd2CMIkK7hMH7EjNwArBAwIfKVqZA27ENclUf4lmRU/hEBHPv0fwPFR5
/LW3SLpEPXFOSzhIauQRyxpTHr3JEzELgrQvyjEcdPxnW7cdmKfOQymQPoKp
m4XmmK7jtM6cTRrGib1FVmzTL+jHGlzdK2umIQYmNw5GnPuH1ZK1GG1y9QQW
bypxKxxNGw5Rg7FArrJU6SKhwqYb/XfWlRo1fp+W+f58ATFDNDWKOxHUUxpH
p3Cda45WhZH/0vizcCJfeyGwlUeEwRm9ltzHEyoicK4LQ5jPorda88POOYUr
IdTsX6/r7FyD00cUFYFclCe2tLnpZa+cp2eF+pQ1U9kiexFoIUD1Tc71oF+Q
b8k3gJOG7LevxYJRxpvdOZNbxPGOAbP6Sz77vONAJmCQIVmDqM+Sq+3AoQh6
t+hJDPYn6rRhXk+YbcPpJnPmnMaWRwCjJPS4TprDN1NLJafeULe/WxBPdcuV
2gDFDpOqRNVPB/0CkfLa59BOUWPWuDMI1+GhP+caeq7cZucw76zz1NyHExpY
MUiPwMwemGzpEAm1FWd4nIfyfGhxd0POsIrcat17eEKN4d8t8lJmzRlj7YpG
bUu0N6sOfGafBo/nA1eM6L8INcuTnejJVggwLIbE5GadV1ui29H/clwd9tSJ
zPES9xIQyQ9sd5T6w++lGlL6GAPhJsZD+SW2OaUzZiOFqnw5QbCfIBC4DLwD
egMiqaX7laNNOxOB3vMt9Y6i+kaKTn8W0KBj8vaZditVaWydnYKqzsW+WYZZ
XmCmMYm/tEqH4G3HgyNQyy1TlK+N5fACZUo1bNxnWONrRXfRBGVNs2S7z2QM
O3wOsb0m+0LxNQP6II2mVSHs6f5g7fIPiGrsvlsDZO9VXClwHn3jL91SuQOs
fj/DOh24SjdToUDPIaGiFPcxGAiEH+ZNhT0unM66oXkFV978+lp3o6m0uv4P
4+3ObYYgXGtyPgRwQZxylTWHLNjt3Jhvpgn9xNdxmORL78ASlTiprvJgLT0l
GEV2vN0j76h3b50Z5o3N/EYlD2RXbDY9PliSJX+eNhm3NsusvWT3a/26qsl7
Tm6GAvJdVQU8qqbVVLOxwQmpwSPJYaGHo1weT/laleW0QFCqKUZ9bk2ybryM
7QIA53ltQgZPeyZr6JOGaDBCCChmHfP9e64PNq0bcJ2fWilHUYVBJ7H1zZYZ
eSdIYEksw1LKKfX1i5rPtSCe6VZDB6wgFI8Rbzvf6lA1Ia/QmYbj3YUB9BZG
YhzFVSUiy+9cd81MJwhqeSy8lr/31OXWV4xN1VGnjCV0oyY1D/ohGzQ9n3tR
lcnHvNSC7PfLZAgaZzGz640OfqIQOhePri8A1hVgCHgu+fgH97VoGd64NXTg
hMwQ1I+xu3uH7nHVv5z8aLjIXrYJsxptRh+vBd8a5aonsLc4XEk/iqEN2/kS
V6ckn94cEV80L0C/38RO4he8ASsmxSBuVbCeRL2oGDHSllbJPnZgMY1HpBj+
4oM43g2oCGXNCirFlgSLI9Xi5+CWzx/09L1weKFOQMej9hzr+K4aF7yu4fma
geNEbBuXrE3m1mIZi6ywJPwyPcxZhHASd+NfYcglS5ZpdUaDvSnLhpe8q6DY
9cC63V3n7+ISJb3Yy0wM4z33Be6dKISjp+7GuNm8xTmZHJEY4B72B6oUknvc
u5agxlLCf8h/Jx4RFmHqcqRv48XuahYzaSlR1soooE2FdccXYWwNsUht47Q3
MGfBC3+LFU4msqCVVeBOLE1E5eP9g4wfXxsVTXJjaNndy2LXPs0yuOC3cHqM
V9Kc6T/ybTG5s6voeZabgbMsfw3cexsw3DsN24GW94PBa/KNW3lDgVsBqg32
1oPq8ch5zer2kGEfwjWzGHSIRpVY1C6azs19Hbh3cr28EglYpzjusu28LGd8
vInmlWAcahmmfANIV8kxWf6pR7jq89k8aZ+8LEd6+TNHsFOxWJPTkTf1YYML
vgWvLh3Lzs0QGutme90wh3mDHQT/BQSwgpzGvQ+ws8EsQeHy9Fh+gt8GDDWA
+zgMbdCpgL8OzwJzCSNpQLfQhHxHZgBzFBtgt9xR/M7Tvt/ASWp9A/BOU1VM
4D7KJJDC0pfBgbTY64figAHpeJd4qDDP1ixsOVhVkJ1+OmHioT60FnC19xBW
3bJJLPvuyBT19PqxTLJSo74ZtqxVtq+j2r+c+e7nVzhkE23TFtvfM4jxv9lP
MYJ8lCPnPgFze7w8bHkq/Wmw9nZ3XDn3jzGbhwp7g4XW8I+vOuiL3VRf6egq
DuqqKvwVkOHAN2fQPh+W6h+jDiPfLSaj0Z5zKVXWKIeh2PhNGuZ51yBrYoq2
Jh5AFcy6GwMDq6CjIJERHC15yds5vP4lKuifx0qehEvTJMLq/lU+vXiQ9baQ
kLkAk3pirfXKs4W09YoJnQ3jJHpQ5AZke3Vq33Dwm+e0ZL++WQj/jWWLO6W8
asXiPTAzEK9iLu1dhmx/67co7eS05lbh4tS8fHcE0ktC2yUgnSWx43WUZg3x
kBzJ0DllCPvcymILnBJYPaD5bIo38kI3pWrwR5DP6FfnorR6kS6dR42Bx8kR
OvQP/5D72naZxqljMS6SFMDa7Z4q9g3e1/4xdrMHCtfJF5oDOg2klD3RT8jf
cpaQ9tFexQE51ZLeZYXBliELWndLfYPXc9Erujy2GHd0GVrfdWcjcU1zAjSi
FfvLH8YG/h3yEvdOJwgPtcWZqqFXX8tFP+AImP8QWxaD113b/O6G9W6Qu6ID
zKabes2e6hXkwz59CUjtbdaNuzJmIW5SPT36qhgtT9MQ6YqV2Ofwolq3IZlP
nge1UfZVdUUTstoHTfrecK+G5yL20kd6APKREJ5jKJV/6RzDd/4R9ceoYXy6
dSSLsTTarOC7Xy/cv9ziR2cquX9RMdymupJFYhAbonKwGdonLAiUwNWKZIl8
lW6ftVgj0rnD7nbjhXxp52kqKLi19oL9hto6dECLyZDvHAzN6aAt5mqyEZkQ
o0PihG2Aa3KZkSnUva/GkypumJV1GYBl2Ah6+PCXL5U0b9NEXLFgF9hLaVcu
eg6u4GuprZWpsR3TmKZThOLOY/7LYXE/K73m6dRq9Kn5q+Uxd1YVO/8x+ht1
F1n3lxsj3nuVfURbqpUmUKEJmidWqodyzf+Px4ATdLfbTFKBC6eopDcnKFj5
6RX4eGryfnxGvl78Tsb1gA1wwa5mgYIjSGY1ufJ163YUF8pz6YayjxolE5mw
bsi8xjzUXJvBLGHrPtDrwZfmvDzQzkz/5Bn/zHUaPEXyHt+tMvLBu07i3vpp
1CcWUqLxkTnHRut3r5u+tpUbJmEo5JN/05pf0qzsrTxZEkH9+ikMht/gNDKZ
IMrN2bKqfD4zb+BtkDFm+iXIYcQS3YTtZ+g5+X7xyNFBURfKkYo8060iNZ3t
maWGBTD01NNi2uYVWcrNRiyS+qV/yTJhAhFlR9NJa6JVHjD+8LLm3cJj80Dt
xEf7ZZjjXKtuvm7ahh9vJ6MFuwkOOl6tBDw4xQUx76nYhTJR0xdeuegnXWgu
3mShQkXKpF7tmAFxE6xuG/t13AZ5qPB5MT8hCfYGJsUzFGYXadbSGgNV/FAc
cq2eau4u8zO4CAt6d4zQUPrbs/h0rsQVximxkKYAYyYOv4Clkt2thnap76k0
d8fhbs83Bke70DS/gFP5+4irR4mQR4T/OoPeGgiEQo5TYlgcWy3xEy30F9+S
y0t7fHNeN6U8aEi9rWZK7KwXejvUQcdP13AHCDS4/3g3vrSr68+PoPo2FFU4
USfeECn4aQ0IeFk2S+dKmxqpOJlAAJdDtOc0gLyBJ3s/hyIxtTyf20Ubg6Wi
R4C78hKhQvJrAyEOccvKUjDeSer+3ZLjcPVHYp405lf44j5nXJFFiFXb27/A
uh6Yy0GUna6+A552+b6fiMdcVV850mT2QhVQEK/Vms8x22D1mmMVVuVE+n19
ptflOunLv7MFtPprOdXs3YXEW5N3JLtcFodAg9eMvnR5pDvHMuAKM2arSelD
VU865i8R7Ym0Bhc7LOFdfJq977ZX2rs3w9BGsWsO8nhXO//tTypE5XIRUJh5
UY9Oo3kUAXIQm2083LRzGilpHs4PhcGowSEtFt2EZp7ezpjjIn7vOJnaQzCc
aQYwRLdheGPIT3HTFi9UG0iV07QEi9vhItpXQAlAnsJhMWIabkNWj/GCuYpd
qn8swhjLIjm6+7qK4xWeSk5bUqT0oJDaEi3TzTRNN/d22KUpq5W5ZbMKIIop
leHu3YxSA8TJiEgEWFMymym1yLZcf1riecby6aEOdmbkRdgnBfRVr8Gl/94r
weU0vJCu8e0EZFvTGUl+zYNd6lj1dIING+mr0+w/fbhJL18ZBdNn8nNEAVSo
W4hchrmQkDoMSMZ5WP5FijnCX3pUT14/S7i0zekE7Zl/bEHyIN/5oucEBRvI
Ll1DZhMtckkm153ul2k45FDMicfUfy1lDBi06Rba2iO/FG9kl95mgqmiQ27N
J9CtvAhjGsYlRs9KOhoT39FVF+lZHjHe2vGrEmo7FXJHnhPo8yfaHY7/hZ1m
F/WOc2KF6Jb0e9dx7X53c8K6/z7yC3Acng6qaCTyiy3LPH/PqzMnkwN1vLkf
CwG0cd3CNbrudxbyMqanaxESLnfNLI/zz8T92OsRVWEp/8vsfnYPYe8PczS1
7XcMqtwDp3LUh26Bj5yjVnacbFIlzOmOWdmG57NumEfSauXpdhunK/3SDnq4
tiZOV5ftTJUXUzAGl5bNvNgERX162hP0RP5lIBNDmaqFcwgV2am1HpXPRta/
Jk2RYuKD/SEnA8Em0Q6DO2m24Tp/MthMEvrLowLqlPUN6uGL4rqy0RKRo+lE
KBmo9DWu/gnshWtXv/TSp/aSm8Mb0c80LXgoUNSWrMbezuNFhXM3lTKqCez8
3Xgplc2Uj67lEj1KF4Me92ZOTDmqs67YuFUr4vXad+UwNNkSF8128y0IsZUe
IDXGw1F+bi20MPvQytUWyImUSpUo2AK9JtYjkUuXsPApEMRHfESWsa1KNmW1
vIP3QupE9ZlB4CVq8jUIKjdxWnRpkqoP0XotAUIQCeHpkBvr3qlZe8DDxhaX
QqR+Y1u8EwJUG+UzezifW2mqnd3ngvm14GzsZVVAyIP9YnhDR26DbNUZnL+k
1bRKDXEnzYJwpilOVcpZdsDgxYx7xQvDeWpZMmm58DbKP4O0/k9uZA5czTE8
fkMoHv7finhVEoicbz1MF0TRk99NZ+NbTGaZr7AmNu35M7JVe+03m9XJVFlJ
I49UG7e8rhBiMDAN9jZlQhR7B2aOjGXaiXgXrTyXJXyByIVcytaabh5uE5Ul
yO4fm/WN3DcgInEUucy7gEmik/B8K4gfSoGVmbREXlX0WsHg6MEJn7ny+eeY
vtN0Lfh42jlbyBaVTLhFXmRY7mkXt2J+0mhJiWhib+Tz/HG07Q2AR6QMbbwt
gSTUrn+MXbb+z56H75K220tDMlNKMt2j0NVMbWKEMf2rYi/HhNNXL8WnrlxR
Lud43Fx6RwqK8CXZd+IS6aEqAXNawh4WMzZPpbV6hmcsZcMFOACR6zJfI6Z7
jHx48UoWQsUP8RAtihe6KFHX45xjE35cBOvCtFMstUzVLrhlqeQYFARpRbHf
FNkDTsvZ/1fbKww5TakYO7LXNoQbCru5rGs2WuAR9aEzgx+2KfcJyFBcEqnV
LbZdPGDrCKSuEGlSZ4a9GhfR6t3G8P7dbKqVymy7b9/RvdZVhtkZVQWzFkl4
PSZVtfpYyhoaXVZvvoOzawQ2Dy6HQbYC9KzR9PE2B6RBRT7VqXpkk1OfAgj1
AW5KbPpASadyw9a5hcWygi+/FCV8kDIJGI7VTvhDuUec2qOW9yK1ulpb/tY+
an3b9w/bOELjLGdLgUmutcpyifhI/8VozI4HN+AjwOdw9fvmX41BRgJIB6gn
dt78AtunENr4njcozsqbk8QA4CHJhZcdXPpJd7Mkw55vkG+J3CXq4e5VOm0H
IE6+Up5oUSKlQ/4QWBK8SxrtDEh/bZVQhGf7pE+uWkLODGm3cttQwxkjIHiW
58SQmPnkjBkQbDhsqqyVjBGDYfkv2qeI2jR8jqSZbJEAe2si1EfEzSWZnncL
iWoqdY7EiDWhPHxJQeAx8tLn5/77TtBjVtzpfMHCvhbWpHs8Pdr/oYLJMfb8
/+6FatD6OQdUB7XnNGB+dFy0BgutUR1yyYl5mMexYPx1FWVYyVaFMYbX1L2h
EHO8ubL7agQCbufRIPfY/7Yj8TWLCzuJJ3X0eA5wLDT4RQdN2oQzFw1V4Prz
kvDrzCr06LBtPsuyOgJ6CMMKoaZC0rh1J6TxXKiAeTrEfoyUcOCQu9fTvJI0
g/GC+CsjjY+8OMWTuf02q+J0OS4EmjBzFn0CGbTIoxjodpPOwnTd/AR9Gps6
qb4qy9sTVqI+nCO+fDujev7McIeLAIsaPDMJrylQMmu/Nkb0Kx8vDglbu04V
pzJJAnVOu6bRv41GDTV5plntr3KlaL6spwwqyEJ6SbIYYLm3t9MeMnwb50Ue
VbLhOdIfaQ1YR6JLJ6K6Y1Vw8w7Wg6i8iJH0AMWBcLA5E2bqy3QgItS8SOhv
BL20+rYUHECgx5PYazH0KzAVRTGWJ/BPVM5ZuTsyXKqqCMj/aaW7YB9RcwBG
3B8uofnf/qJ3zMc6F64ithlsJ+I1vheZvmL5AnQoGYHm5bWJLWoIT4HbRIDQ
DGiJxjAENHlTZtWNMF9dzgdhO8HAOYLEYESWIkFsvgBzmRkVmNoT42kygPOw
3+3JC01zL8NKc8hp4+JPyq4JwGrIZ6mnHp8Ccp0PCE5arY5KZTcGCCrs61KH
EFaGQmF6zS0XJxAV9dNwJI+MCCG2+PmIIurRkBhwYFsxdMWd2NOgry53PA34
VbTNu608Akyj8NEF9G6wpiHHQwyBbmx2VqMNjU39G5+aoupBN8pa/rZY9Xcc
kORtvGjjn7s7AYoTe+IjH3Ai/a5oN2shgCOI0Cpz+OVGpq3wRBR/BzmHsaa/
B1uenFUBEf09TF5qLnos6yNpR4knd/SodGselyPTEOYGP7OthHFfMnFBUJjX
3QkaTqUlhO56lFzXL971LdMj0y+3LXV7/fNFvE+iUkHZddC8bu0K7BlQij06
7K+usrOBWIgVj8Bft9olNbJf8glti1YLo0JJTo7rpaTSykTdTrP1UlNde+mi
xDxDDwB9OU8Q8rGWmyhTGIkA+WGhs8Cqvz4WZkvTxxQ2BXRwrr0kUDkNCzfy
JHFJnsgmqVn47JxCzwBMdQMp/flITDN10d7+JUPhWwX6ve0/WNAzvTzJ5YK5
gQe4mNEFjAFxUtd30d+VAkFNgkk0sJVaktllOYHFQe13JhAOhwKYSx8pgsZ5
6ZqrpWyHbNMLMcjZLc6x6IT4tt5Fy8nvu+J8WMIalVMO+5nXh2/t3ZMbiT9x
5HltpVUS6/E6Eud+joNhpkHWyM8Y4C0f5RtIdolBC+o1kW9AlLCV1L0P3Zwq
6IkRQS1r86KkMo1+wtvtKEWB18x82sJfFYZ93X1/Bb+B/o13j9eMPCRaEFA8
+aqwKpIDGOfI5giUHBY5HC7FWhAPZHyqmJBbIx0lWknFMfCDmn87hnm5Klvc
DUT6IUi3SVO4Jp5U5WClbCMKLa/9g05xOlZ1L3d6fGgSAC0HQxrM0MBxCdNP
YnxFRObjxbxjudG1wRovna0iEBbktGSc0w04QuZcp3GgIzQbTcvDol6en2EB
/K7D+LFW3OhI/L1BA1KKlmZhgAhbNVGLmCFyUS8A8FfvQ5H3iAvWfKa0TrKl
KAc4p9AT5Cg32JVvEDirJ6r+qM3lm2OG9op96fo5x3wHILyH1XjWd+rE6WU+
gnyy/iiXB+5zciP62B+i2vlvcpJZCTiA8QcEYgOjI4JbEoGmboWqeTDnQ/E3
Jhf4MCHF43No/zy/pcUIKIfzSl8sZuEb7piVh2Kks51Z55TCCW3Wc57/MmFV
+aNwwnBJNNYu/Yo5z6PhmBw+3DPu2147Wz9bxkrZMKwhrJ7Uhqxzy9NA4ux8
SHi5xLEv06G6fsSrmHgEzUixzvd2bWS8A9FtJ7JoBBNiW046SA6LZ1jEImsL
vcSs2//kDJxYd1HLDsLoOf8fkQVDnBY5fGJchrvObzh7T6EENbYWGLp+R94u
lOtqGc3c7G47EHS/PdcbKaEx2/DOobaVgDEewx8YwIyrvKn0MgoV7L4p5dNU
GhspaYIq54+Og2XPGNcZOw7a1cEAdEQSsOvKGJsShcvkyuOvi+2P9/j2w3Sa
bzZMEaVNpDjn5Q7+XZP4qXuaw5OhflMRlXzdKwyVjcxC5AgqJ087eBJQLpby
TjULRYRs2pi+dd0GnlsB1zQ3mCDP6arI9A1+Cwh/VH9NnDoOCBUaKS5X0iHJ
a885P8ECCTo9prwbFQTPQC2VzsiPFmp67EvGmrBvAQt6DPzD2ioqIWHOScMn
cYurDY5ATW35fW+nCJ6mb9+kCB5lw/ZNwnA1oPb6EfZYZ/fZ8r3ydAvWgs+y
Sqds0PnbMgLbaCskum4+7xFmw58P1Wi7Iwn4Vi9bkYzpiKQ4uIjMA6S6zUa3
HQaPiYHxVExkvfUP8ldaffS+P3olUJc70GI9hUOxCof/CVm0z5SS36W5oQHx
johsId2REd52wRxttYRjs8PDA1TdJuMwxbfaITydP8qhAIWelIx0jPNNEcce
3kw2YkPTPfDLfpA8M5SrdX9tvSslikElGznxKRAyQyesSgcrWkHE2G1MQO+J
TxrZCqoNQ1SsW7Qbv8dfdt7yUkpMi74WdXaxk6N1N3Xm8gEpvdrNARKJMhnW
r59O4yR7kAT+qOgx0BDYMyJzIrE5gHEqQ7ZNpQ3u0EtVLk0y9hXRcvXXVCV9
PEFupdtCIYnBxJ5/S//Pi2ZYkSUnP0i8sV8IEE2feJRvCPqFoCKIhBhmtGjb
JTNaT925kdgITfmvZQWvgVbfCriffnaxQP4aBw5ZHShYVUSqhCX8G6pc/DFu
EnMt+q3zsK6KqqC5UtV/il/OouYg9r7vgEeE+jzWv/kVet7Q9OW0SdIZpgSa
yzKaV/SxOkCVJkldsgClF0Z/1QoIls4WaG9z7VTrYULaviIrKWOiRLcWaH9P
YznI2lmiAgopsBNvOEU5SS/69Hl7cIuGM0bRz8UScrTNg8HSPVE7iEy67XKy
RSuDSlIfDbzPjPrBnN3Wk8Jj/kfUvcNMOOIhztOSsp1xFqT+rk+ulL6NWDc5
EdPzaovucCZPDStYif4WXX+BC1iO+tJZhaTBWf+PC9fi3ZKcy8OYolMJlQ/M
n4QvgSpKnGkns62I6bwVBgnyqUfnXcZbwqpQ7BGC4vfoiKQJkfvw9aQzNADV
G8dtW7SuKUs8IqsJmxh0fz3wROb3mSHN0lrNxuQbKGyI736sY+/LbEop1gso
sBC31PwZJ1rXGbjjEh6FDGAn1B6YoTTXB6nvQzT0KyYAzPiFKX1HGSzkL8UP
nXNkVGKdUyWRW3h0Twmj4cTr1R83qIX55oX+Tp2XeRuUF1hLoxBuAXRL+V/P
09S4RSmZbi0KmCc5dOpnqzCZkHoeZemRj6lvWM0h6LNDD+N0OUnEYOokJS/a
wVCquvYaDCxOAjmIQMO/omq0Ze/YwjwYqfa4wEn46Lw/+HKF7kINuX9Pn95q
VeyRlp8+0FRiVnwKZvZyFGfSf003aLCJLPY6rWIlZesQPKluAQYv/aMGB3ga
eZne6VPImnOsmTg29tPdPNFTuhAzPjzn+6e80/N3j9OyD41zhxG9UMapK8T7
8iUoaJyskJU4eh1XiXcwuPuWCE4gczzsV9ZXZz0h6C7XJk6st/twvAmmgT2P
o0HHrEnplC27nRaF2G20iIzRYJmyxuzHWZsCAo3iILmIHY4ZKcU6FebAstZP
QunbCko/r4nFSuviHxZxQhWxquhqul4ePi/NqwFHHYv+yOrwg7OIddm81fMH
TbwUHiP/el4DD6cHAiiK8WXvRDU1Fg/Il4ZUidh1o1IJUoRrjzOlzH7GBLB4
TCxJ1FpnYSOL4qju5ASMxll7BxSbu+OiQ+JxQ4BIscCUQ1z0bx4dmzOPNBoJ
fHl2XDwNN+9IXp5NMAaZUNPJZyYsVOML8HT8njKe7R175u2I6zUbE5q4UjqB
pHHy2WGJqjxbpTEBxgZ4iV6bmtWxbo8qtjuTcih7hbQbRGp0NNJ8o99I3gzM
/aM/FpYFgpiFseysS5FaadLpvcbjtoBIAcb3tzfqRsSv5/Xd9o0aU9YpmkyR
R+xWxp/1DqJ3DUjYsfk4ZVxpNa8/0MzjjnIx/xwtfYvF/zr/TN8H5ma+bF7U
BpI4+ErYyKR6lnNn0SJs5qB2qJjAMTjViMZzIbudlwNGac96T4hY2YG28RH7
sybF3ICiaQV8sEt/neoRqajL3ON4b5Vs5rWkkN/pOgdClY5cSKfehu+XogkJ
lLiafmJPhSsBl+U6g5b3dnGPOANd20K45V7nwN+cRV0KCUHyrGC3rg4qqr4t
6WndXs2UpfkgapbnlhDzbanxWwsWfgf5+SxUp5+QxAIK0N1fN7ISpOsXarzI
5rkrEZjNB68aey0b42ClC5TWb/25oFF92Z7c1yDrHvaZhj4Wz3S8ZajjhFRC
zIuj1OzaFwMeVRDRtmq/lH6qbzR9oiRjRBNsTw7fvMby2+BcFCxpa13dJZLD
FI9Qb+Iovb5G/Suy4EfAURpiYFGpkA1iXxRlRFlRim6KqOZevKN9NXC1w6M7
9aZstJ8kwfYm3Ag+sOqJyte8qD76/5mBy9vzFoeCzczz7ZnJkQNYFUG6/1v7
CK0IarMo0J2zGxP8+Q4LPQPXirKJOxGXu59fZpv4y9PpAXHMV1mIPtP+2Do0
mQkYLXvOFt/yDSy4kH38HMKqMUyW9WO1XTkGbpHL0j5PON6iHcrOSSKlCd0V
/pHin7h8eMAWnTNtwbLmpLj4tMRNQGNTp+gsK1ELsvWKDWV3B5bKndGdiVX3
08JGMe2Zf9eQuwuskDruFrajUoRZKF3xhMX9SbMF+/5Wkxj8YFmtl1OmbQam
TBB8x06upnBlqOeAOlE/x3nCfOJhrt0PPrv0yzbKxgBdbxZwmrmc27iu/pty
RhjEhMldNw9V2xh21fzIl4cb0F0x3xqm5IBRzgQJl+xPqYJ44bWSoAAAmPX6
FM1ja7tevArCUOZ+bOuvdcZCRateTguxSh8x8sdB5wTC+MUc27Zdv12aOE0f
OC4iukDkbj2TpEQPE0MljN+henfbqUr28glT611svm75f+7rS7aOD+O7Hcxf
xJFV7J9wLcndQD9Hv7LsoU8/EsbTK8DMeYXpfRosEeIjVEgVl+rZ13NIaTb/
r6KjiX70CaUD3Nt5PSKszHd/48OQYqR3aoEXdOgDmHSbjqrzejCHfQKLMxcR
Lsm4GLih4eHtrF5K8ZH3Wk2oCpoP1d3Ite9Et4UZnKOkCp4yztCyYQDrY0T6
o3+C3fxQIm+sElHOnBlwHJe0I4Ihxj6P4CdFlVXYKlMWaXhHMQHLcVrV7DSH
Hy/j2Iree7PS2QL5aDTk/7h4KySpV8hF/a5RmjWAcXIzW/r9mBjRKaKpq6RW
KjorI2+RGyzB53CPoILfNqcr/+yrvjI03W4wILe78g32KReuz1X9UL17Fgf/
S+OPjl2bQ83lN1GSSEQKC0/NWQ6sNUNoJrlnZadNveJ4L/0SCnhw/Q73973P
/o3Ixb3gk2gnk2FS/GKYNKByu8YyHLOTpcf024htNzr9wcF/BUbtlZxEBV4A
N40tZg4TVytMGokzSREguJHJT0fTah77jgs2Q7R/lsAOBj1mJRzsFuNpWthe
K6ioYlYjpkL/x2v35ZtrIyB3F1QNHQUY2ErvfqyguugSRAEtfy2prAgfCyI4
fymPB2OQTbPheg3O0n4g4k/0BexFCVhMzb+Q4w1+05xyC4SUy48zJ7fv7ZXS
nt7FFmKoLJVkvrJwyJ5MbAP1Ubjp/AdW5oDSBGYriVPCPXVE5p69FytOc+sD
CFFVqFNVLlbUjpLIOoAznMdeojI48m45uGzfSNvmGXOe4OMURFxDSl33kniz
4g4vIIIf07uIJVoAn1hu8aR74QiI4uGPW6aBEPsyUYc+/0HsXx4UDhLYqQq8
E8wyew+WnmcscF3oj6Kxd1mJ1zNag2FGGiSVVs/sqC4svo7/Cear0t+5GhbM
WzAATFy5oDeRDsEN057L8BQqUdTfHzKCHskZ9vkc2q1R0gwo6plKjD8i2ixM
Ij59Lk4bUQzg+UClODHA7mB0vzIxoJZ1P7UrbagYgTm9euqiFSnckQwVZOwi
SOlNhJP2Z5WC4Vag6GSC2mUtRVS6qlKux+bQABUCc62XLttiKJw5vO3S3vNa
3piCYdHm0squvvHKFGffB1OByT0ci1UQE/wrUi0zJEWqn3w9+ydvJUS4Xl18
qATT5BTrvTxkoH17abED/SNvoreOayvVbVa1ZS+BGWhEHL+szWEMcRF0FOeX
hdl0fTkv5lVrNZQIgM84cQQYwja1+H+iUVchc0EPy0A3D75cwVc+qRHvU7kW
lSIxRBOG8MAhaYqzPU4G/1SHAEDmmqz7KZAtQtuOWGKDB/XxFpZNGVj4uMxo
07BTDYrwG33PCy1OuLotMk85TfEH4GfMaqYQC8n7iriofzXa3iXNnCg833bh
iPPZeAf2yho9e++OWI40FqJo7K2QUwMwNBEQjSBVM2sE5zW1ga9pZFM4Tp95
J1JVCJPUMXvFi2HzLkiS7nHOjLptxoxiwavaw6qY5wzsnk0QdaIc2llpiqcD
cT+1CcVqprIdXxFuT604o0GxqkaGCPyjY02xvzHLXLti22LhDcqF10sbT9nJ
KIY9tzSoWw87DLo9DOuGVnziOpWaRJmMLCYnQtzN/iea1AtbpzXuqhlzqZY3
7eCBuDjSN5bWrU/Unx+qjQECoyEaK9O9QDGmMLH8Nf568tK+gFNzLgTdJm/K
/c5DfxlqiYdolAmETrr5pypVt/c573yB9hw0PGyri4BkVN+uwENNDupM2lk6
IvT4brnhtN+nQgLhSZQ9nprs9p7B1JOt/HjRD0P2110bd1mmQvfgA24ZAncs
p0T1LkYPvcj9Crxc9bu+rlVy+sV6cwSkk0DrHmur0lNYPUBg4Y2n0+BxCm72
peaS4N58vM3XpUf27+k3Z8+YZDLXtN1v9y6ef9Qp87XS03Xl1ruyxTeE6kYI
asOyraWmAlcoBy2W8Raay+6tCwyroUFpEnWiggdoz2G1rgrjCNVpiU6+UmKt
jS6qMGvsnCCIJHuqAVN9P+y33AGCFkV6C+ffPuNCLswYgAzkOYGQTKfm55Fb
+BPqj3LaVKOZx0P6gEPqO5ciL+f2iuEAwrjsxT3QpgBPUuNoBQUbU4lBG9ML
aP7Ku8OqJl76BY47oQ8L/AIh1j6fyz2z1Docf6t8itfCg68Qrr3UM85SMuQW
k/Z6pHXI2by/nQl+UsqDd5pKK58D5y/+ryYcH4wCTpAUzAR4p5gNGY4y1Qdt
OfthjaGpCDYmcn0TlkwMvEUDmSumyxSa43aBozBpPEXJvCwX8c08DDWFKgHQ
/+rtpgmUOoxa1r6yqWA0YYbUmx4A38dDZ412X3L0BOJd4SoiLK1gBAgbNjoY
PhvXkesa/8SKBJwBpseqWuQ20tIUCm51F1qKMG52GfACx8lbruWSe3v4t9r2
uUVrSClzArUxP68px6Kzyj15wADyvyRVIaj1i5lyqYDpA05kpJO5NtC6hj2X
L0YA+aX5LWQ4lEnZreryqRjzu5UjB3oBaqqQXwGPhyM15eog04NYF/k9apTE
DSlQu05O5mgOjwEHNN3v/uzLS5VuBq4Qgyr7rYTY+QyZNz5lDCFDYw+id4o2
r2sAoCGoY49wgXmfh5izSyQsdokMqsuyxXWyXsgjdgcgai9Wf+jfbYXuaO83
5jdxSvyysFV8Ss2Kp7LXli/hwOPUzs1WokZeAaIAxAtLRCV4oLhmOxSllms4
QAZzvkMZntd4MamCLO0soVFGTv+qFDv0PEA8GbKNYZgMq9nxiw7aPAgrFj4Q
zjOwL50Nc5dpNWLwa6sfvGE95WkO6T1XijU3XxP5KyFnCYBmXk8xZhng4lsA
WmzFZlxJ7wIPQKWUBJTmAnFeUu1sDGV4NvW1cevWQ9sqqoNW6MkxtflB4FOX
61upFTkT5JudeVtFA+CMvmKrxe+1toBkn0vDPk5huddEBKgF1A3fKHXHQo6I
G/oIBRGu7Ru/071iKsQb9qlkAssthJnicv8Smvax6iDzy4JaC+Xq8H0F32dI
bMKno6HnPFWA2hDc1kd1OMOw2DpXyvwHoeThlwnVHw9Ws2EVOdKso04/A/st
9i+Vfp4xPwNL7zUU25nx2quuG6CsJQeGo8u0Wo/zCYWhY0yYIp6rgwD8y8ef
omiPcIAnne6tu3H5ZHW17YvvzRZQ8fBw8voBAmP3/qSBtViOpV4bGtQtCNPV
SsfiHitbk9mN/wVsFgagDbkSesfSO+b+rvcnEzC/BIu0owL82ulhSyD+6tpq
JpTzhpGFV7CUPRo7H4ysG+DpYpTXezMO3heVcpS8FiD0npxu7WvZ5ERuIQTa
BdLH59t75ISZYKAJ05SWafBArIrPXYcdqA1pln3lzJlY8qgexziF6KmFSd2i
ddScaIX0eqztiScFCogNAzTdpMmdxL/aLbOF/D8ADkIZAcsBaxgl/3UC+nJf
g1U2YF84uUwX2u8BmLDZ84fYDw8UTf8vehipwijuIm0NVV4LmAMfLj4IGwBU
RsgPIi+jLblCxKRzwO7Yq8ILRb+MuvBf49/Nttq9NZQIeOnQ9RQ3KosaGVdk
6CzVPFjo6YvLjiv6bWWX9CWGyzFMRFqGyKS+NjH7afbpHxMPjytSn3Zf5iuN
dbAlCM8uiGSCRxsyEK3zGyYSG3QFMsiontFhLd/fowQ7ENVntuxG4Qsm6usf
gY7N8xfehxbjoyg9jD72Z3iMBdwKd4tDIGCRb/FtLZF6BKYk5aGAjJveElZN
W/jPVHTLdm5LBbmdwB40H9xf5ZGXzFclsfF433fL3C5hPhFsM34pu6B35bS0
/nJX0YmXYDhtcKs9wlbQYoHeSu5D12hgc4UWVAVVofdHJ8jyRriwhAmTvnk0
z5bsu/jbSM4sKART5nk+y0Q6Gz2Xezmw1o7zPV+lPYeXGLqw5G2ciy7DJ36G
kyKB/+qcRgqmHCyptWO6S0wasgsHLXHIrky4RGFhecwEfGcjqnnaBDjCOiC4
BTfkzoyc7Dv0sGW/6D0S02qXaEsdYUq+smeT15RmcV6StvWZWPptmoZNrtbJ
+WLDv1KY4mCN6y9lcJNSzxUu53e1fT3jqzz6EesVN/dKeR8quPk9gnpK1W39
lLbEaeMVxwFXz+iKYAld9zatkmJhexv/GrQDDq4aGqZmk7U/i7i0zFQan5LT
tsa/5j8iBvtHYRKHFjcuBMk3PAZQ8ze2SN2TV4fWnz9F/8c1PX20ou4CmBr1
IOfosS1lw5rl9Bxxi7oX8q2cghDTrh/wqesQ7/tWqISD9eT3ssnhcgu7z234
t8SIzzH7LTlzbOjEkWkvugUn29hpdIBQmfCL03xYRWVz9NziWWcNJDu+hK5y
OrVYaADc5ObrBJGGT6vlT2oJ7INJqreWfYQfOmrsNTyzfWpF5KMXNNDQncn8
gEpw0PRGaIMgUVgpAoLeI1wipCeOQjXrM3XnoHfSgppv3fFTPCtoNctKjaYG
zK6qmzKs7Zs4JzbRvf2Tb79z90PUwW2R0HNleoGx/83fE0bOUhKfOSQP89/C
X3Gx+VA1/7yLpNjcEm+KmFgPDY/RXvjbC/eJOlm0FQ+wHGdf22SNBPKxm6Mn
uC3+6+1GJkrm1PGrOMXJzy1hNtD8bRhf/DhacbpK+kh2jMVoX069C4JyNdqf
LXFtqzr4JwYqPSh+ZadBYQTHrO60893KiVYqSkronnFPigCqRUe+j2xSFihO
y0+fr0baj+4Lq8nwDIH7PLPi2gAOKLPx2asEQg5aQWaGZJTiHb2oKmFowqW+
mtXndVuG9UFZdNBkb4vYrORtMBKKM9zmZHHRgeLCgv8LRIh/GCKDya1nwK1r
E2pQ6vbAfBBm4c8cla1l4BIeVoie6M+NuUk9Qdrwm13SXIphUqByhzRZvemD
T1rP0999wC01TNp4ySEbDxH2hlyvHpzWv53r/CnnWiZdbyns75TI38Zsx+T4
1GtXmtBn2SbB+P694Xjl6WUU9A2La8WfHsqpkTn3twMbmoigsifZ3ZQpeKKe
0d3J4UM0AAnBOapgvTOq96Yh5ZvHwfEhRJVgvWhdG5e+wEaZDQWqxXeGEeD1
d07j1lG5LJ+U2eD/eA5TAOOLhiKAPT9BlDP2fy9UIn52lp/E3svcpUPsVjPN
98Ty0hEU3NYHCQaLjZiVK2Wg0ORamN0mK0c04k7VyQsMA+jEN0RJAH0W6ilF
GKSaWu7GsB1o0rynN5yEGS5usQw5R2/yvyAdNJbDD3vmJezkwqAfHSgdT/ZH
JbnDGgeWofMjz/lxlpZ8Koc5fEu7PFZdCtyZetwKak2Z7Sjxs0/dOkPCvdR2
gny85bMY/LZxd/bpxnhv2U9ExicW8wpFlh6+4a6+GL6SBLrL4yQpkpmc1uYi
DSVob4wMOF8HZl48rj77mcbiz5ni+le7bSy5PACXstyObZ3ieRLzp0ylVyr1
vS4FHuv34qXbOtGLfyp0gLMt7ok7e/nwjJ8e5lWc9lLbp5L5GUGzNyD3dYuk
k/dtdcYkLHJQblWLIvZbPVsesD6eFCIhSQdr2dldOdOCdImnBS763KiyG3XW
QOFwmlHU9Ji1R0C81oSsRVtek2JE4+q6FNVyaXtyCKtjvlvpBDRMI50BIWph
k8XZz387ccWLSRzQyOfFLaelQXaqHqZwuuW5sdZSW1tL8p1ljhep69pBUBS7
FodP3Xc5B1SFMy33+DmAUvCGLZDkomHW8817BW1HdstHrirLSk+mLgqMGCne
xkcGBs6DvZr4WZWIkrZBaBNhZeeEUPJGBsksCjq4/5ddEeqN4tNKhS1AG52i
LJsIEomRteWCeDNhtLpq2K3d5VJM4unaLIWRw3Lrpocv37o2uB7pJIOxafJy
VbqoxSY0wg3DCQojuBrO0oSmPAtHEDOlvO7iipiXHuqi6oVek6apX+/MmS58
ALYjF6Q6y87AkoyqtyWCIW4AX+PSL8ljLlOVAeZtPMiDhHlQZypZof8pk7di
znw5dfO8BAeRKYFwQ3Z4WNacd+hIpj38fakCHf21EeussEKPOZ0DgYcIGtTC
TSKc63roHtPugCxJ9jvBDpmvoC0mnl+g4nPwQb3BtDNvh+pbOuzNRW0DtVxY
OzgqCS7J6hX62WQyeZ7fOGsZH+4yISem/RLiTymTeuZMgeFdfss6fTscRLyY
5+YyD3vLGEkd/BZw659jr+bXTEuA1eeGkaL+Kk3Q+5A/kEO7suhqOTEfu2HA
qNIaj8wvPmSJ2YsWYXrVErdOPXah+GqK123Eeax0RDrcWRozxCA4mKoKXzWI
dkF2Oy+9VMZVaOWiht166y46rV+m4a4+fCaKMy1I+k1zZ7uoIg0bnROka9xv
7VPXIlRBQHcqe1+XMFXKadqrO8EveJy1TR5N97MFaG8Gr9BO0HxKXCsxAfXa
RIjCvclXPPHSfV7T4ykGBaE1YsmLF6TkoQp5wx10E7/2af/QKkF8YDUTbfPd
zXp2ARYTDVL63B1UZOl868g/qyHDM6QIZmxYwdfaAXFj60QJytFku0e0Pltz
3buVAZv82rlV/gQxNehXbrTA5CiwPC0Z6LqWhjDvLk7FRwC9eF+vm1wQUYl4
91cJIY20cHbnfaOLjAEK9gBybGRbXDxBqJHJM1czBkSQ0ozeEBUIHlvug6rv
1xKKjm8fhvMSBfmQbZ/zdHZYrmZXZx3JOYXKf62r85VGe+2hA1S8vowoT3r8
64vjunvCHZB4RcoTgDG6keTQ5JT3vXV2adtyjQ3nPmnmuO4PQaBkMJMSpuGO
FB17GQgYUt9vGJisihLYi7MO/SK4s5ejYwiuCBLpA37PVc6PhUa+tQ5pBdSI
OuodOjECh4gcoS5dFmBd2dQZMD/j1VJYkoghvIobqCZbvsK5ggLI+eHU6lJ+
6nec/BGPo0UiXah9VHsNgKiUK3YO85+GHsD5DJK/mmfiBVi07E8ZGf78ZcfP
ky5r63d093anRmz+7aW6KncuwmDFOEmrUwjA3QoQeRXlBWAXPsOMXZmPQrz7
TzRyfvyuhWCm3VGmEapFE/afS/hLFzHT4rO0M9Dtui3IT4Amx/gcdQNSb+I1
ie3nw3KOZJojgBMvVeY4kmkFSNtz/E8HOzEfrKJTWgOHG5Q2nM+sfdUY/JQN
By04rAAFLSFmY3Oat6PR0I8lYO5O9nyDRR5fU4giJ8TNSuczzDIevBFRsCir
Em8y4KnCqjrNVyaAbwhhRJeSSanhntlmAIvRUBM3V0b0qP8bdmeEkLCZyO8X
xnYw67eAnrxXiWYAP7lpYDk9Owk07SprQWCSOyhfRcJqDT4yyIE3AdNYbsxj
XqeR24+9OM4Jm8X2LdXJNYCqoPf9OCWzpvssBzkfThEPn7tyAadfMLHfa6FM
cZ0ie6sGYd0Izg//a5lQv5hvhtffZrEtKrk2zlPI6vFJfAz821P+0kS0s5r6
3j0jRMc5kST86z0fP8p+zro0BasuoN/zYgEjf2XE2RO55O7c04twQ3CfHIkx
E4kOJJ+l5Y0LK6R4sfuscuPv9ZQA/f+AbLli+wVH7DuNeG1rBAhmsdA+JdAU
HbEr5SD/NtSuvmd0pCxTd2HbTX4xxbpJzPThUlqnXmvsKzJsECuOl7Fj7Brt
e1lrCPZM+hJtjSzr/dvU1exnj0qlsxE0X5QwjZ0wfIMmg0M60TY05LGeD6am
TpIhrAR4kpDGaegfk3ZSmGH3uKGRGt45T9KLk4oqNkj50uNE3ccN9VMgL3bX
nhIfIGFXOhoTDtCxeugFhilWQsgj5rjIW03omhVlSjiV2c8BBVlMMQ3eY3aC
2qaquHgLn6HfnJflvCJ0UOikne2EM29obb7kkC2Uf1JK0l0YjgMi9tFRApGT
5TPSsM/ddkeedvr1TPO7FD5u8nCz+wJG6FZtujE1iRlrMhF9bTtuj6GhQfj/
Mvgt/DmfqvfcyVIsVM6/ftLI9QyafvMnsu4O8iXE05xGjU7f67vTktTgg9vk
s0sL7E0xtKTsJUMgTAj/mRAHEaqfX91Cmq3WhOmBMt7NZupEZm12xkJ7Fp2M
5Dea3TI3B79I/OHGJL5lrsl3nqwkwt2zeuVvBm7wqHzZVoZxp1jTbmlShgMP
QZ4bKQKHWP7TyjbfqfInlNNLdsGlUigHmdq6VSGL8MVSB2NV/kTmgJcUzYYc
p27u9BabA3ocjC8LeosDWfji/rMYQ+ySpX0j41J5u1EfiuFwHJETaMLRFTwO
JYtZEHdFhyggjLPObvY4HyDsT6tT1ytr8bUsDq2IBTTtzVEeAAgtce0nfqun
fsqePSxZck+V/fu6I/zwk43j5/G1PPLQ4BgEsHTL/PpoMUzMimSe5Zr7aF8L
Oz9eti8pPtc3oDAhCCVkrxE7tYlM9s1J3TavDCGDO20M7Az+Q3/btyCU1TdV
taeEma12jy3VZln//WZhNttWxhe/X85eXC4j5qifAVlS50OVAf/Z80V4rD8S
Pj3JJ7F9gns40H0Z5b33mS8IH3Dz8bPDdQ2QKjYXAWbe3ebXBcv26JXpMh1B
s9vt0aGqIHsZMJQL05o2gqBh/Ex5AjI2Cwyajp00Fzi7F0PO0GQe8Jfhr06R
Laeq1DphJKzqSzUnmLkc9WsuRE5qu7B9Pkvg/PLP6LZLX+SubgmM0YFII4/u
+yY0YxNR7LusBncJtLyeqxEAWwNPGAFSybVR2AZfs9geVUARLurmgFeSGrw2
zd869VXhgVVWHlZokbzO3lNzRrcuIeWhJk+AE2uzLXE6GET5XkryFp193st8
iG9ydwFJmu3Uh11joyaa2WESXqSjv33W0q9Hs/QkufQucvZs/zNZ2zkmITZG
t0+yAq8028ig+rXrRWvJrYAuZ5nKenuCe6sfaHvYrURjdGJy6+y0yAelotyQ
xGlsXEH2Nyq0AEMUAlyPqUnH7+GKCbjdqnpcFmIvFBiCJOwq3c3Q6NQUzHV3
zTp0TZQFj5YNQVjO7SgKTWfh90cOH97zsgmJpmdjGERYg1Soj8iwlF3RNdUW
lxYBkTYa/NitLGIXN7fZtZo0SG1QR9uuDJrGHYoSX8RjO2m+995DmNi7bRUw
YK1vyyLpQmIdVSBvmisWS4tFDFy9xP9b2i7ra3XoylN/H9BbGPASLqB5GeDj
4Loe3KneVCwCNVSp7lSBhdQHylcDhvLpAQhIWLycUuw0B9cZyfi/l4lO+WtM
XD3iejPC4kc2lHMYkxV3lPxLwKQ+jSNSfctqJkZWDObpqt+OzNWA0d3mjVhP
xACDnlqHlmhMx9ZMHWK431+NQANSiywxCJk1VNaz2RF3Ewv/ETlfKXPEDh81
nidVs1Y0WwketX0iIEU5A06tEh5RIoiaF+ElXa3u74BEvaKH08I8fVjEKez6
QoDvuWOcdnI5RF7httJy9h3b4C4XNY5lL9IkneOBnraUtiClZSQ49BMYJfsz
mfSIYK9JzBRaYCwkpOp2CoUL/BoAW+5MhzvBALWi/3SsylG9UzCyN0/CDTQ5
8DwSOp2wFJ7ovu54rROXze077/u2CKqpn7nWAMoZRDfqvwDM8j+qSWdDOhcx
AMRYiUuuF+FJYXp4jgX/oooOgpKPnycAZnd0a/WAjVRRvcaS1Fx3DCc2ER7q
9Utvg7sQ3zgI/CAs5oEBiFlMpvdptv+xlKZIssbV2y7SOYVGpVhY9CztU4ez
gewamgXoxRA5zaQQs9/K2R7YUQPO9m4uSTaa80zICenk71xtIQi5jnYUon0y
anRrsoSVXurLUebb8upjN6UObEDdMIYipZTdinkaTgtuzGHyj5tLljtYW2Po
bHX754Ph7NAI6H2i+4AyKHOxomHhxMCHXSYH1ZrMwOXv6PoRLdYXs+TRhIis
slbfQtkuVJ6NgXQAZfIQZTYhhx64kA+vKV7ngbSqryBhO42+u6l1ZZz38eMg
jca5F9nHG9+Jk7B3c2VATsYae3MKeOkIh14rYO6sNajpQTwAqWDmYIJKtva5
qAJk6MDCCdkY4iEP7ccydb+sEWl7TI2W8Jd+rp4F6BwHDqAtRiXsSP4uP4i9
6xNwxWody1iEVcR08m4Fs6wQ8dvm3cNVBalnItAlBONRQAB184ns0ZpQIHs4
OpOXUOZB0GBOyWr1ZM3Ex1c1efTKMBrl4nutrkHsCq3ZAUighLTJP0jpkK4k
ev/BuNqU6+bN8baHFFTpd7GLFOi+ZpnLmbNsWPjN6WEew+CSm9lJKetTs2bi
/LF/uPKv/aswiTRbzDJETUBgFvOkldVCCXzvB2OCMb6FOfMCZZtxOhd1zoIk
COHNcSIfqLqoNcxPI3UR+faC0Egi4pZjjcXp2UlrFN7uhFXxjUaTGTHawP0A
hP8SIhyKln+YcsApb5Cj5IZOuCF5jmrMVNi4hbBR4zAcYD+wyGnoz4JxV4m4
zN0Lnwfjpxu/98qcUZYvOxfUdXSDJfi5Hx9j4LV1yGuCHMcKl/VYr7PzSqCm
vdtAVPnan5XiQ0pF7HnuM98oOpuh3S2eNloxdew9RgQd5vuXMGM1AIWbGESH
nlZdXI24Kq/m041QbnxZ0fBu2/y9vWzrTHBhkPWPYOyEuRTDqEv6sM9FemDf
pNz+X5ULi9fSu8Lm3mMfGJatDDPSz2yQvpM8tb25dThkx1Z4d3dhGHTVCSph
t73SwUj19gLFeyqwestTmnZIe7GHkAf1Aj7ARFvfaZC4NyA2i3HWP++8DZKs
0Q7/5JcicZoatjKWXBnb/kvQ9GnzDCYMPwyfzfya5i4w7YQ8uGEFs7nN2WLI
RWS8X/vPvR3cjDcQ3MMJYo0WwrnWvEh033ZlzXjODWxUftyfs5Jw2adIdWqQ
+PPwsKI1QIekocIAyI2w2Cqplqnc06Gp9ptS4mqw+fHYO8fVQnNr/IyZwvvB
bRKhN+CNWMVHHdKTKlJKMJnVH9BC1WjCKk54W3L8Hlpo6hWV2CIqVrJtHFcc
ezBFjajy5pmjaCbqv+WN1qxIrYbHyrDSaZC6uYG4WlwxOSF2k9j1nWW9FwB4
IRWMeRlBd41ARrDVn74G2ESFwDgSoLzL08XMRhNTdwIvusHreVGGcDGrZNCV
E0m0xVn2z4E52AMc/GDYnBf/ixy2mArVSgBdMzBo11Dm+AqcmekZyj6fB7zr
CWxR+PhPNmt2zNDkGY1ebw/7zJObRtyhntzKxP9WXR0Av9b0pjo0btkPE74D
FrKcwvN22Jw4cBzlHFC/w5+BRRbmO0OkENXuq40CsisFznHAR5FJCOnVr2Jz
QA6MYTTLUrXO0zvQI7Ryvog9fSBHMBPMrb1knKnG0s0xXUVvnYBCDVaqBA7Q
tlyo6IQaBhQ4bu8Pprs9a3C8+R4alJ6b/vcWolbJX7lN4GyYpZqwaSzJK6LU
erQkus+bp07xKMPePvlBORJ2ACJnrpsl9jEH7VgPhxVvsWaP7eeG450sJqXd
tqx6SAu9XGI0Nm7nP0sUH4Hv+qS1xJ9YXHZH9MzU8RUhodR8joiCZOwjd5tp
G7JSg05e5PIXNyf+GFCkPjHJzHvIygGKEBDB1a4GqtsOV8HTfampy7nE944M
+pbDPFbWdtMKlUhNMIFwlKTDWVy+TYUXnDTojLnWdDQxKKRS2krfjrcAdP/g
Rc5mz1u+v0UrTDp5iTo0iYtq7tMvP+xO6AOoGTo/yuyjgns8KQG4WD3rE7ue
RJPlicYB1v5HK+eZxT3DA9GwNp5bG+paMZQUTMbcukHKZtL7lcEGBQsLTgv1
KflcOSeFrTcyCJFbLs6JgnOxVeeHqhW/U2DsCAACjnB4cXsx3p1i0MXRZAOD
RGJqjKGAzxhwqebaI+5rxiCIlE+NkUEDHZmd3memPwHrXCXasbJpv92WQgAN
B1ZrvCr92N/Wln1IkgWLDhcvVBPod+o4Rn7XkI2L9FNRo4cM1Gp1XSWRMUE3
Kjo6KEACpKinvfDjlBB4VYpT3AWxpe8uZiDy4GCmNMBSW4D6GvZpyfGhkY1r
LlT/c4ij/J73XLBrdzIMudxbyxAv3E+R6TdUtse6ZZSVZJ7ffUPrWKVRTZfx
+5gXzg6gaRRuQP9hH28M8GNcOfES9C/crsyptuGYNTNweH8eoL0ksicwR/yi
A/pdnMPaDHl1uLWlAx9dcOa6Xp75PB0wLdiOBiKPDLpQrsQj44tDHDH4EZll
OH6slEAM0/RB07W1H02PjGvIJZN9GR80Ta0YACf1XugQZlzINKAaiyIUIkZt
lbjlMGHlMav/mqULH6MAWMUXRPPR/iI2ZLncs33ijyKPR0+hpM3IDtNDUmpI
dMY39XAy0waHiHMgZR6/8Ki7zG4sAr6rbiX4FXxhlw/JvqYLApBO5ClgK2nZ
yn+/1PludowjNg00pB8N/ZJzRAOSawnsaUlryyU98mX7PVRJpmxOFjaVWASA
P9nt9hmpTYMXTGaCiflFn8kiB9urOZVG5LRNwZXV+FFuoF++O/KqLEKwGREY
BxBsEywZlSObQpbQVf0R1uRHxBXmJ+gDwTxVBYBuX16PKZplVhNeJ4q9rzU2
83XupmBsiP5VmXJRcDJ8E6VtAsPGbtZ6d2amPNhIKdRlO6Oadbqdtn/rGyoI
PIYPaD6pKfD+1d97SqqEjr112vUsh7SLkr0Kyk/7sS9Tqql6eEE6lcP11lz4
U5GXNJrjsu2XuTTlhKGqxQplXCyaqC2b+6040UdngWDhf0ZijpyopTIfSrFN
Af8z9ZFKu0UxSu280AWKvA+xdA7X7cHj9lGjP2BDttobK1/DH5OqOThr5vZP
NTxF1BYAxOcTMSWubydCWWgeUF/nChBc4kXhVNPlzos78AjuhAeUaNaQIeT4
08oT7SEaIzlJSge5wAmW1z2nPSi7u8ktW52VqE+bkZBK3qAMuWdr6w28QqDD
nuns0V0DU44pFRX0eYKkxVGUMMUziB+tfa8mGQHQD6/jI+kEI5orOwdXC/Pe
/+6S91B4AX1Fb6qDkGVZiyL9NaNpyxMG7+7HzFEErWcoFHSCTxZlwJKaD7fh
/iV7b8cu2Hq2cDt0x433/V+yW7wYf2E70/1EJ9bQHJ79G+JTc5y/cR60uU8C
6qL7gP+kvjQ3rBAbRgWhnj7DLM800yQ8qM5x5klYE7GGF1WsNx1oXraVR7G7
3HKDuFt04i2E+YfVi4NrKhgvc8hQnjTERblErhmvIXOXIMzrRFwuLgRuoAzr
DJ1ejlYAHWO9wb+tCmkmhMhV0ifOYKMpvy/zxUW6M2sqF9fvBVh/fF/LtrGF
JIUEgjRDFFOfVUdWknll85prkBqAShkerQ36CK0u7iMpgbr2EdUP+Ln7OLw1
zn5jxHwj0WAP7TtlSgRMCgxsyyzHBJmtyNtuI0BqcH6kz5qBXS+dEBPV813B
lub7fgf4u4935UZz/+iqtTU2X5Pn0y0BlTFuYevKU9u3mLDHNxDnnnSYJlKx
ChAhLbfteq/Z344IuAp9+q5ZT7xV6X393X/raHdltUXwNDvM9ZmwEDnqFotk
xMkLsaoO7zfodIpLBCzgBlBwO/ydXg2KD+k/U32pBSiCqHUstn1HQWjUD6lG
iMtQOqur4evvdSSLzowuzVZZWryjHhgRcmaGMufuZ7/3bj7s28DPA2LEk+8K
MoM99CWr5Th8Pez2ipUN54mY8zfkeJ8oyq+PC32uVlCku9HWDjj1dTrMpxUP
f2H+IyhUwc/zpN0NvNMWQnoL49uSRk3Li0dxhZHFa8Mwe0JwsCNqjP597Zbe
MmP0FINZIivIiQjFJ2awD41EP+KTHKlKROfseaOlmtoYuYxJzBZHjxaGLt2F
m8AZN+TAGga5FthR4Oua+UJ6B0ZxJJyaa0FBOfUmNMpbMuAK0ezx2NEpqtQn
6W+4YFKut89hNknaxGKgjMhKJkQiKpEyGhcJ0Cy/ylVlo1yeQ+udLbGMeCwK
U1ENSu98H7K2e0TORsytU7SHCRKsOEttVXLBMIvm3C9GcIarHypt202MSiV6
u3EdmT/gb9iA7wtTzmXVwQCjlm0UO3aeGyN31aiYURNTOjozHnlmy5X0CXsk
g8AM207rjhd5lS8weM1JEJ5/YWOKZgvTAe8bBK80ioIPPqRHdBFj1kKaw9hV
dNfFGWzfn3TwvCCsGOVDg/pS47tK0R0oigusaoNHIJOhTylo3Fi0BsutJbTq
IFX8daVN+EYUkuOd0sxihJLiO943F0aOM/onr9YPmEJ4N/AXYM+P/s5XD2AK
qpKcRiiPLPum2Z3KSZf/NY5Y8LLTyw4PENbgkN8kp0NPe6k0mNniz+v2kRmM
UvNJMC6BVKPFdW9rWhP/1CnC2XMcHbLeK+hRYcp4gdndw6eCxQEowU+JTtKe
B20HYIprw5Klo2RVj7AVeuWisIkFmZNBGjvCm6mgAqepxciBWlXdCDuHS81W
d7ZWFOyT8ozpl/N3KfexoNL4i3VqPwb9OAFh63GG/jEFXNHaLcpVy77Vk7Ui
p7OAo4R7eAJXzxMkcWLsbeYyye2aLztk7tqg3rloz+HxoQnfhbuUpzmSPqO7
scKgGAPr1ro65sfgsoHz6eWHF55Qa+uNaomNk2QNBInLc02DpUAMoCO77eyv
gtxn0GZO1FeHWulTFRQUNWSZcipKpmmkjjt3wReRsam2eAe6cYpWYHMhNd+n
Mf97oYcYbOEFZJCmtN4xdudE+ucWp/Tw2/zy7L58c6IQRVCczzLnDmFHw3iV
aoyy8TcfD1s8jY/1HB0624V+hveSCJ6HjRUIq1mDhYYjTml9DlvUnz+i9N90
IndB3tHEG/ZfWF5tdwwrJKEekgLih+IklZ1Fry2VAYWERYeskUQHcs4GlFEY
uyZv+gGM+imALn6Cd4/djl2hPQVoJ2xJmPE3Autqp8/X12OHw0/2lZ7voJc0
i6rjh8rPdbMjZF40a48eRY98qObxIDWkkT5myNyKSF3xepU+fLu6dLxYP6c6
aq0H7lB1TW3qgQynYTs29kCj0+D4HEVyg6cO/sBOuK3QfsuIA/rk02i8dRp3
8Q08a79BOMjpd2PAreqLiYPdioIXTZzIEdpHwbT9YPya8umjmhgUjpH+g49I
uuZVdRYyWrD8szudAjnkgZPokYlvhvSBvQS3WXt2Zntp6hhaUGCm3zupnGfS
m5BcjAOMzVkRdU24ui9aMNNUkZbXORAIsQqtE+l1Rtzow9dlLcu7nS3G+hgn
Kdl4JuGiFO/f8Q8NkRWhJ2JJsdccQlrHDDah8dGbORclawU+luYDkDzBV2Bq
n65JYXWW3KFroSohRkf7a+QIzMlTkO1q6vVeY3e1FcGbP1N9dKRQ/Ftk9YgX
vAcYmoPYZ+L5843LnnjnSo0zfgZTZ7cKV/Deqo/SyYaijFOtPz+GNz5gIBej
7GNMRRF1xnsM6spDM+hMbm8TYVuw1Yxh5JjlkXIbIyB3b0KsYEnJrEwfDLFB
4squgP+PHADQ+fA1RhShLY4wNkVPB1LRhsQ/9sGaSw9o1AAWiT7P179iv37i
kUj+KiiWJYChdVtR0H0hurI5y4zJH7/PP/aPct/p5NDqiWxLDuMT49SgooTE
/ShReJ8iT2vpovzP82ZDyf+lGF4ygC+e6l+5RlTw37ulisCeew07TUUzbDkH
Dp95e0XimGJNsnN8y9sGENiZamgNDIez2muakKnvHz5tMosfgyHmAH1tMRox
X0cCvUe4TwvnawEoNjuQcCnVjwWcZYNx71nc1gWuctY3RrL28WbVXePRC+Do
aynW5VPcD1rk4QMthW4oDS9ux/s7WJBRDvE/Egkcc3AsdXygIv4qRfydV5yz
aPNczSxFB9toEem+9WtSICsv5S1W/nJYRQHHdTw5N3PWhITfuBcqluGXewFO
GrvSQAhblKt41aJCTk37oQzCYczRJwPrNz2uCeHDD7UI1EqYWV2X/kjXi3b2
/4Xr8zNj6z1IAATLzT/yYBRukzDFPhMCv5wsbh+TgoDPE42jHIosRHKdxMEu
VKS9ICgj1YB2wBiqvY2sVkHnuAs3vQ8haFS+F9XSfqx+5EvJDqQPWC8JhpNf
C4DLgJGwEvlv5H3pkwmx6o+epaDpxUQWpjV9Mwf/DP3fgBkzBGjXWiDmAujc
+ZE+RRQFmIgRe4LQlXkfIhoYViHX+Pol9YqixLWAjMm65MmfsJXZp+zDY7It
nylRgT8CINRYiid8QP2Hi57LZ6I9SRnK0cLtEbOkKLwfqCUZ2cqn3ceXBpmX
L1AMD7A/7IUvmQAUTrqhfJCSu2AXUZ38zdwKwhUguas7RTj2/NIuY/mejTzl
MrVc0ffu9/04Lv/mM/UUbmwk0pa6xDt419F2VXaPZt5Eg+X/+iAS1RlZsC0c
+O4YKFqUgta4A7sCktGlFTV4Sqlfiuv+z8RQe10Zg7s/L+nipebhPAHMX1oK
OQtI3X/+Z2pe+NjG14PFs39zmuE+6aYmT8XSKJyv64M3DNK/AVXgWa+Bm/N/
WhFYjnJtjlwFSeLMPvTkOXJAHZWYpdPv4C5pZDivys8x7uESxg0fS6F9vfrQ
8XbgauNqxmBEjKUzNOCOect3NRjCEnNrpWQy5oy0vxEX40o14etXeOh1bSEs
nIrhrsGS7TSc1wbHYCjr86rSOUSqwZ/cYKMmrrRmZNu4p/oytNGwfBGJDodI
zdous6gfj8p3Xx95YP1FRgQIPRJE/Z+qLd0QxdWgFw3F+fwOOkKrubk6PMEh
rZ6xaERdOVduKaRuJK43LonNMFodc4lBfhBkUb3iFZ7Lt/vjMhEHVsrSclgY
A2edV+fSaynyj+eWwjcPT39MnjbbLOJRGMztFMK96qnYbYvFBPnkoztOYxsX
aEmnxSj2LqVNBoNrwPtkzaPwQUiqTpZx2/JrHd3bh/vXe1NbPcGeEjLxJAKN
BQfo1APBNDJjL3/kJrp9Mc/HqWG9Pi4zzYHZWs8QJp9g0RfcF0GX55xZkU8+
fNfrdsClqckoAPH3neV14VnIqgToz9L+mRt7ZYXXVQa8450VF7CrV+zsumGl
eiaVu6h8PSzr+TwKTuvyyxEuG7B7GNxWpBIWUofJzCbsn/fok9vK9GMubFBj
eijswknYraI9I4afeaAu93tbFcs0CarZp6UCNVbZUuiW8QycsStk0Oq3lgWD
MZbosHOrO/4Vubyi0HoRIXYxgAlh1lbk9WXnnEnP+QqHOV6g3MtFumTVdG+8
OWd8JDYE9Wx/enqaoektYhbu7pS/L5nfHNMrXovA2GylVRvZZncZW7m2SMcE
Jgz+ITXiiYh7U/oDsyvMamRDKrgCBSHEBz4oSkKe48cKhEBeIuhhCOHpNU3J
6OwPg+3s/974KUbERhKp7UVr90SB4kCaBpxEYH0s+3sqr7qnVqiVzoAy3YjN
jsJsM6SY7w7zfDqWGX3y4Ak6LX+HnHZYhXhhJHkpEwf2ibOKr9bJOnPbcJVQ
hP7lPVi337pB/Nbjh+6czEJMEfJOELvhYHsZ3FdCgtPzDYg0USSIM2YR9sUb
Cphm1SOS4aQOf40ijDZqjQxflA4qI9NLBlnz5YTwfQEoap3t0bLdujRvAfqQ
rYYyfbEXv0YMX8/RxSAUSPW8km5sXQ7aJIAMqWgiBBRi9ftcbdVxbkPRI9gB
7uvjGt9yQKs4aXyWGnsmHd+Ee1zE9M/Lu7LLwaIZJqIDbXRjamMZqcJJUJBy
DXnt5J2I6rQqhLVYe7oN7L3NCvBr4lR4gx36SFn6aSnObNW6p8HtznSpxxT7
daaokkOSR0OqlwvUAcfkOK2NFq4bophyNN6IjxLNzNAaqiF6om/bl9k6NU+7
yDCw60xlTTloSH5V62UFgmDtdaN02stpZXBxCmV+So/uvG8052guC30ffX43
MRRvawlGPjKcz1h3r6In5PlzMypWdgr23EHvaLeVaaidb6b6M32U2osycoku
rRpfXb32+T3yluLcgeI2r7hBdDoSPFY4R6dVuuWs991yAtezcR2IN9I8Z2DX
oonqJl3WlEFLSxnCO9bVa83AKXuKpgZzKP9nhbtNAIsKV1q24PZ2cxAc91LI
vMRigQWnRpTUbq+jeBH8g4UQBs18FxZ7yPZ0qYGWzpEwv64BosqKBju/gOnW
LxS70vkQ7FdWV3ZD9jUnI4qtm8/1G31k5l1xKF0Bu84t1I9PX9X8z2cXk998
+eOraRhUKsiojZjo2brISZyg0iX8kYPvv84F9ZADQR0cqGY9OjtmXagPQwQX
5a6RxB+yAroIL9IBrbJ75wAGt7hVs78KJREtZiiXvx6Fqr6LbZhE8cobp9QF
A+JxD/6P30LijKn8tnX9nRQ0tUWigCFT8n+v9tQGcdWBNLmvdR3lSIk6g/49
KJme/XBM0xZ5ALvx/Cpu/S2mQozFNDpOGjH/L//FNW4uGlxQxLsVGulOlsDC
8EVM5byBayk3qbs6f9kwTNdxiwcSAR9NMUrb8HEqV9ZiNcSEismMeU/Hnb9k
AkNWXt3P6NSH6MVeik+3qzJIEshX54KMy7oateGg+rIcKB81606jxg/pavLP
nRzzEnPrttu9xS+jGBIVEcZjfAVxUE8iBTrIh6zfNQci2MC9JzjjR8wW+XEv
pU5+BBkCXELWFmoWbPfvNXopIedYkRWMTU2zL+1Bi6X9jeG9a4X44HPqOjLU
9XWcTJQXDayo5uI55/8Yom7e5hJAJGSpRguWWB8Ku3GJbXulT+u90IuFCApY
nmEJVbfali6EAA0mv0g9WDWqU0MeMziI+wKyoVa4Gs7i/OYrCxY736ukEWKA
oALu+Ez32P/saoqaZxPmQVnyl1WWMC84LGklwmicRFjjZoHdQy2IZ1q05gOz
QaOHhzt1ahw5s02fcDnRj+6TrBTApu94BH1EX9pANOGkD+emPbMUg29Pb63J
NYOF9QJKlSY537DhL07ofRPqjDNpFW5NGRkQvHluADH7px42KaeF3OK2TU78
w+/7JLAtnPMMTrLm6UCZlxyOTUhc7fllrkLwdJvNxP44VdDrqaM2aspbR/Pz
gDXz3m2ukHtzWQ1pgBvf/wlnTZTI/3lpenJGKwv8GqNbUk+AJZju2Go8uaT4
NB+DLU1ePAC6I43Ca5oIdi+4X+uP6th2hOxdAGyEevVzuCUL/EeKl5C4Bc6L
ec1E7P/bQV50a2MMgVO74ATA3eFziG24/dn5J9o4BRAbbvbObIRUo97OeJx6
0fP9TsFioxgChVPoo4ZEwXst94L4swrvELJyS06adRDTWFuV8B6Me4BkzQxx
FpW0ThOM3mrpsRmnyTuAQnkDsZz139O+HHFdOMb+f0xg6QQByqni/6/0dqid
Lod7DRCCBdzdi6MC7bC9ca5TqZUAUAaAPxsv5Dl9GOyZRVIeQlf0k1X1pWfM
/SwHyG5FpDCytUuSFPyVxjyzCaWzeyA8jGWaeIYCsIWxQDRYCQ9X49J9PbwW
W2vCkcbuICR+Cv58zVHSSBL/XY2ial6TsGvxwiTr07TSy8KoBcKu70pBxgWn
13LBS1bHVlXU6kxxa/jnurVn3ysjdHDe/+c5KTnTutZ8IKi5+5TxKmLV772D
DZ31AquH+ru6p8nnUTJf+yl32ZcOifNT4xArkFVyOq1BdOzYqiKHJX6HZhYd
dvm0RvoN0zAyxMhSEPmYr4MG8cxlh8T/B4+Ge3AQj50QEKe7VJYI1LpmZhoD
ByD368BAvGY2RIhCIqxRjBz8BNe2Q5Zln3/h7y0JZZgTayIhVeS3j9fu8Wi1
ps5imcusGUi/Lp5ojgwpMtSX+HkMtRGwseAjOyZUw9tfzfPzPci7CIXSk58N
sqtPUyFhbrTiVQ9FoB+gtoCOY/8+S5IAca1n3TB8hYF7XP6Kaao4CzFqSsPf
rkklP+jyD8bNtEXeYgx918CXqqDiXtNj1BBcdT2bG1HQwPExv5oodYZ3ozhX
ZKl1QRL+RP1WXHeRdne8oaiV4Ykg5LD/Jk/fysVEpls/oqscJFLPU+SUz9qy
2mY0BwgyKmS2W3HtY9qJAj2t40ePMogVa7T4PCBjsFITNRXvGWXQWq7KcHuv
OtVc0vJJRQWYd+WrjxPrIbgpmAZF/TfqrHh1RjCWGJnl2J5zGaG7BSPfy54o
qmJsio5CrDMkeRY7z2S6TxbIWrMatk4l0ImmerOrbNfvVH5MmgMpzj2N+KH8
YDGC7grDC0DDi+npQdeYXifbXARKi+ItMb3DON8a6hgTB3j7zu7zJ/zj7Yol
ZGyMp3IHjgX1/bQmG+vTASlW6Ebm+o3uv1alrTUY19/ualjmcgDRYERW7QrM
HmtFmEl0YDJfPlQ9h/PCsuVNFnDPLxbnrvtpeoY5Ql7/1deb1Wk+0eGnbkjF
bVTndaUadhuEFXNd0kILAzWirfQoyycz2UgpMaiTdzB+EUe87rO/4ivpq4x/
NGtyxhEAcYFzJ1pnljRWBVM8hWxvpxUHvkqezJuA5YAEHBO+FZbF9/Jjczyb
hvDKB09sNWbrcFtXI75D6YQixVEfXCHimJhLsdBrUWHWe604MtEm3m4QLhFJ
Deumctvt7DUM65RP3ZcaGpjwFmafEuIVgHCCQTmwJRFR6+VUi61DRBzaCYF7
NPycgavi/OtWIBsdZ8E4uOJVgf47rJBmMZZInL+ZggiAYe+euM9nCS8HcYAe
HPiOwwIUyYR3nZQP7tfQxqaT0aLLpwXO+aRXbTFTiW78j+TS4E3jNgaonw/I
3eMYoKO/6eIvVGCwfo9+5MNF79AZiMNaTpe3W5D+A587deiCNhSdLHd8fZ/J
9ctOvbULpplGvIYWF/a94IRbBHLah/MHAbZ2we5Ibgx/DLCTMF6wOHDpeI7+
Vbakcg7J50lolj8ATqJfrYY4Yq+cSMBjrT/n/CTnh411BsVw/OTlt8lhvpDX
ExxUAv3ZueAAP0UFs9+lKNOCp/uanUPjVl8ArAKJz3CPNFtB9Z/2AzFkHgYb
BdrSbcp22ZqJuzswHOGTZcGEd1ibXMBc5inj1W+wq3sCgU6CeXSuykp7EooB
payok3GRtC3ylPOL97tRRqzGup0+znZfs0OEpii/9kii/bgK9Xao7cf7OnOk
ThLCp9zDuUoX4iLKhflPspSSU9Aus2Dony3sDkMVcPFqcskCej0ColFH274g
ocoSXINXmz1WbdZhmV5Kx0q0nn4rwMYgUH8JHXUlmgwhE7m6ZfRaMLlOtQuY
g4kUuhonIe8aWrYV6XcZrDfxlYUHaO8I8lT9t/kV/2iAVSB8RzkJJxeheBrl
IE//2MUZrSk3FGzmwpDx3mQpWRMpagZo4jEpwGL4RzCCo5Zv+ZTw0S7w9opG
+pyqcoPrzbGNBjg/WWQOMSTGrMKv21WmWV5MsY9TSW2cJv0xYvnafcL1mo6G
N083Ve8APdOq3T2THdNpqRfM4i83x8bbWyf9yZ+LNZfo8UtLhVSiLK4nLkrC
3Y1C2pdtKyKLTjvp0X+vQT2u2J4KSH/eDHE6Zo8aVKzzv8HvfyG5QjdkRqsa
H330lqSwMA9DIkkH9Vx2E4CmbU8GZ5iQ/fE+7zhMlv+y28d8HhrMG+pAr/HH
RmnAGp5VFHKcNaQj8xOiUW/1IHdNq4Cgj2mUQ9V550/H2iy9B8QcIONNSnEq
HZRoM9F2HCTjbQiHtl4oCAngfNwqaYy5q2CzfNlVHDXhW/U3i+QUXReiAdoe
3RUzbVHpSuBrDeDDD5hl/LX02Mw2iRmcCFiZYHdyQaS+uazs2/Qir4n1AUni
AEYNmtqc+Q2MSisTeJYh/dZzEeAZ3e73IqshCA6QVYpkVyk+ZXIebFyMjcXI
9Vwm3835j2w0mnKOtT/ZW/cNg+EwaXyD+02YJbll5WXD5Nic+XKDeLqCIWi0
SasaX7ryzw0s05BjwKIjN67tl4G8JJMTQ+yX6G3pWy8ST2erFeRmRXUPDBQU
4EMhMZ0yug/AcONLiCXoymO8n+b2hBE6tMZjvjAjGU4L0vRgIhibhKPtqh/b
SawYBjN14fLXqIhkHfH4JbYDLqFNG4l8oGft3/bGZI2YhZ8g477J15oD+25J
fLyyqjXjFWxyTeJ8DEQHjVWau5b8lzn6ftJoXXKy+YRTHHiYDfUITKlByZNf
EDU5aMLunHfLOxH1RROiT5FDGSj2oWdos4g9Txf1kyytCKewhozcWyAVlldo
4g/+YIJi7KZJ5XMoeS/ZONp4JI0apJEtFjGsVpXinFmOlQKEJkdHoUWR8GQ4
0iCjcWrCe0HatIp1Pm5+/WO7OJi/gVABPqvmyWo7DMFJxI5uWHYx6BMIr9S5
49QO6Ky8aGrICKOgyGFx3y1deSU60WTLSFCELSvi5RaR1LFL+aHEMvuocdMv
EvELF9pfIofsEQkOvXgfkFfatgTGgEQOwz0JN5lx1BvmRfoThYnUy0JU/Mbk
PFB3vETLJJvwYzBDnu0ZtBD4RGZyVw2FCAqJYK0KG+JNmTHOAME6AA0Eo+Xm
FiwTKn08GWBTt21ZRcxpSAfdgnmpwpf3KO5ZVcGaY0aoAu97nP4xr7KRLk/A
G8HlCnn/piR+octhpPjj3qNZZrzmkR/dPIfy/RmfpUy1bnCTiXlJcCNVxnSQ
lmB+EYEnChl5/mJwNYdiontLJL6bf49KW9LHO6mMTwSJEJOoBykE24s204jh
tjiBNh6HdFwhW2HX6ToUI2zBPtA/UJzFS40Fda6lm/C+MHKUvpiIwI+2e8Vw
aL8b9Iu7+b+Oqy3yMK+IthTHsoRwLztuI3iR+TvQ68I70LO4KMMQFkzfuSUo
R4mSBFaVTQyqzPYyQ0XkgvKuhnih0nI8pNnxn0vVS8EHuDn/t6Qa2Dau/xyz
loEBqfPzpW0nvIsci7NbGc5DqABJaqquXu1n6DVTD17q3EW48jkswPKHgqH7
ehkyJ6c2XCs85ng/cQKsJ2P++35lysLI4aqET3DpZ63AxQ2bvnorQl9yydFL
M7S+sg8inROPRQxoqYaokjP/GlzQHYzS5J3Bvnz3XcoXI01NjDP/roWuDUds
m3oO+FukuD7DXYxOyl2bdEZSUuDykw8olacX6BhNS4U5sIFLXJfyQ0cwCBfk
98CwxsrXKdIVGQnyv7bOp11N19UI1H5skR3KXmSTH6FmvpbKCAbE4Org5u4/
9Cbrn7ioroaez2G/ASkcI+jdia7A9PdPeGxinpdDItdyByFecwdNOpPI123r
1IoPDgDCL5sbWGk2vi7+w4XF8ZeEg58iiIo61lKzgD6CEIfTjBUwzbJCh8P8
qKcHI8huz/EvR7zxEeKLazu6cS0GiM3rRtVx1SO7OZIpvEOqJMS0PbqSHMk6
0TV3Cqq0TemWKHxczkG3Wt1CzDk0KVtmjjY187JEwmP4GyRZqRfLj7rBq2wE
6qDheaPuRpi0yt5mj2KoSvaMoB6GyDQXtV8LZtBl8g0AxLdwA2mB0lGCKkTm
WJR4prtS87zbcObbtMgb8mphUHKknq41PYQTYkb7h4hF9Z5Tq+wjZ6QSZtEN
Ewb90Mb9ELGcbZYpXnQm1T24WvrCS4HQKZKCYpryJT/a1n/TC9KdHqxSwyKt
iwOvIuEy5fUQwXKEVEbR6VkrAlzWyrj8ThmSdynKIw5gF/Sybrj/yMWK/21O
ziJ0ZgnwDQhShY10AZuNk3PZ/EOl1cAdufngrcnNn+SmIVXGu/d2Q+T9mdWi
UC1g468o2HNGgsDRo+AgSSeh4/N7TsTFFUy4Z2gzgUpa7zas5z8r8S+aFvU2
P3AHzO7+UjyIFcpfzPOr9NkF5HjrNeD3TYeSnJvDklPm/JP1QR49asGsCCX6
fowh40SMqmsQO/+EKJ1nHzFn3EoHpQqfI+jvgCXO/0XaXaua0wZty2ZG4KTV
IbDmw+X04McajmEhcI8n2Dsj27jjR3N0/PsU/9+PmEbZxTW0+d4LA7EsCcwr
JYh9WDu4+u1lApz8MGaeAO/ISLHolNGnT/VMyn3S8+ED3j6K33Q1jD1oSr65
5NmgpOJri5V29Q+j6syoYEk23G/HixPzVHA4DEv/qOZYCKgjX1x/svIJnHcd
68aqGc4ZttE0PON7z/rpFSe5BQ+m+9+Uuol3IPnQyhaGe3Ez442TMRnmXLOx
/0ZrwQRvHi6ZgdICON2U0UZY8wA8CzwoJPxVwhDCEs7quWOSxqxdpH4ZuCUI
6ehLFkFm+4UWEd8imZ1Npr3PwOFf1omutK/AVpepSwdlvzL8kmXujY5ojlFq
eTBVZKRqS7sn99hTGxzUVAo7LX0nh5cuQiZAAL6JD8fucsyElZe56hrm+D64
u5hUiOrKi8FWiStu4YO86lCu6po+aaN/sWscdCskmFKujqo5aBMgx+MoknLA
tItssWrRMXcJEmqvEEGo7Kxq19eOo/sq8PFnpO7xSbsEup4J3/iCukY72xv6
+rrwOvVt6hU8SaXWCKdwvefQc0DFj9HbyZmypUx6L6ijJMg3z96K844d4XDG
UrpR6wVptJ0uCEutRxoB461Rd6ATfDn3unxUxJMkvgfCewvDVw5elShfhvmo
UdmRw4ynpwLpYUjU0LvM4YpuxHa9Skwn3uMkCU3iXGsFV/LdIVRQWlYfaSRn
+MmtOclvbVVjnlK6XefYJUdRZ+C3TILW34E6wez4x9gw/VLTS4BHhusLwFVS
zutCxW6r3JUxz0aBPrRVci32OtTPhNF+4jMuofHVixoWo1OQhGXZB1zfor4X
FeI1tmHQPm5rlE7yxNHkon/2vYKKLTZeEK4Yjjw5xNOyNJ/9f60eoeU9mosl
Tbrs/Ybwr+AKOpo2XcpyJTydYeiudKfZj72DrDlze+3Zqvb8BGekHxSoky4l
tEyRuU0+bUXe+OY8JTXjIa/Micha2ePtJ1Rfx2rTZUVKr/YWdj/sqsMW2VpS
iH3ZWIvQp1ChEw49mQ+CjAskivkY9vISw4imdrDH3x4kapFsOvjFcbAc9kka
mf0HxiphKaAQuoXpcTigNq22XX7YR+22RUz5cPO9ZZ4FgN4aEFl13s4jfTvF
TBtbB5fSYYtq++wsrZDTbBbdMRzf19jA6qN7u7zMzIAd9nGF4QVORvuzic6j
G4OjrnA7JF/idShGEH9QyYLKXqdn/V9EshYps4rQBG2IhemnrPNCe+Ybq6t8
BVsxDizBBivWmCrv/JuO0W/OTbJdEtELXfC9qWQIY2sMFf7VKc4JEQlzKgV1
U2lAbK+IynEnGNU+4UlPC+90K1B6B41zx6gl0uM3L4aocFV3NoaIL7HHRAs4
2sVS/dn9ooNtLEZEgAK4+dT70uLTLlkxOluoRFh8dYArLSCF3qrBq6f0P3/J
Yl048en6g5N6bC4hc3/dlHwgpML1KpP8GZsVVTH+V8+WzWvnYdd2/yalsd/c
GeDLoQaa6oV26/j/ktSAHGOJvRumC1m/6aV4Z6p/lk/DZULcIf75GCIYYPHe
Fr4XKDfJYFEz9uK181Kzy56HQ/pmnFbOJFEv/E5+Iumv2nYHfOREQq4vu24j
vcvukfmbNm0ELdGuwkilQqPNmRmnoAUH9S/H/YCLr9MawQc7dh+z/DmrcNwQ
C1uduMGNHYb8br7PHI+hdvM00M1Y4MoQmDtE29E3UblFR/KQium9H+ZxUbvU
JmH9J/fKU3SOBFFRCRQVh63Ao3VmfUonJ/wKKGkGPEJECYPhAnzCEIW8gVMK
R2wcR3KQYbckq3D2XpqJ3wLYQt2977hjGQTjTxPnx5ZVRk+RPrCts989nrLd
+rYtuYIGLRlNCQqioMc9y5R4nmejsI3zNoJ5wdfd4xDWG7m5o/Svnx+IxIGE
3eff5aQngTCwok4QHX+lVjKOnlhrLWBW/IcJFgCeb4Jk6M2f6SYyTvIJtbfd
SJ+v1dC091bAYnZcg8gOM/LEJnjfmo/NKJxCeJzFK4JmBR0xQuh+H+eG3Cja
ZSKzUvBB03EBGiXeqtlj1auVjh/YsZCctXrZgwGyGlCwiROWitU2tbH8756h
2BtGrOAP+6pRj5u9skVcr6IAwS5O/vXvE2IB3djhVQjshoQf9+z8bqucKLwi
YQtAfHW59f1GLRdpKoj5SJruWKxNmyxuzMEZpDfFFrgV3lmEEv/3zu9wN5rW
fSqjj994vyFioJIsTED0+m6nsELGG37PPm8VhdmaHUTF/chYfMc6+xrsgiO5
Tx2cI7LMzBrqUMa6Q7CLnt816AfKFNX7slubirRVER4uTTldAN9BMD3IfK0O
KWfHj3RxjJxymfle9CqxDRvj3DxFfDqcTusq++ZT2L+oxb8LAvQaySVSqK5O
fKREgrWRUye2N+xpxvuinAgBYEman/2J+KEDV7YEHTW9FGcDVDpuXr2W9myj
o+9QEtmMoQSRUzqZMHyJ53VB0XTqRzUCTYXGZ6+//lluPf/uGv5VmXqd+IFB
TlZnCtxa4Bj5C/Dn2K1ruQyYh2FelCUhSlip4xZndZdxDxjECeUGuPRhdaDJ
97S21acH/RnZ/rznj7//Kvn25c9m54hWQcMTOUoh2QlUfB/smVri7+Uw7P3A
QL+auMI7zNrsQcZub0gnYeV7Mk3uN/bu6PbhyL9JAdgwZqLILTRVQb9ap/l7
uf8xTaoMcW0WtcwqdBWx0pe34epj0HKBPLvJpoZzgG18O+1Ry7RT6Al9WvAU
GzN9xh/Uuc0MU9/PtbZh5rDBhtZyQpL0Zi3NaJArZOohjGN4WzgtbWZKzHax
V/uE8U2tDDvkH/6ODQnOKrET7k4zhezMxmQGiawSr4w57VHY5Y3Vxzran0qj
jV6hkLTS0A3W2Xt6zJueqFMfEgJElXhwWFApoyEn5594d538O2H7piEpcLf/
AdD6VApcTktmXosPmt+bowKdj13xpFxvBT69EpKnZNzYXVJAe49GRIhlA+vQ
+uFB44rJ01bEkAz2kpPJ22FAeqZyDWNwcuRVvsBVO+ViVqkdzUASItaRMEIr
HUpEkiIVWyO6qr/ewJMXm/PnMfrZ8S5jAONtNY6ixvj7yiBtsOuMNwBexhIP
FD4i99gdtStHkfO3woMNS/xhvA+Lf0vCntRscvjSyrnvGniB0xjFXv1nZ70B
gjdfFUPaxU+1q1HyzuqAmuDJKu0NYTaj5nT3yKARijY3XZGZmQ4JfIxhD24J
j4yGBdctfOCpI1xmXT18qJ9vVD3H3VY5qGeoJfSCaEeVIy3xmEHLAipDmkSY
KzhpJVnc8ze7j/wtnOpSBnxpaP3v6Tz1/3pQ6qdualx8bA1bBnPtVE/6XaBc
Sn71kF3jmXIgnsYCIEoUFmOULmv6FWVHaK/Cns0ZzuqQv4rhNc4OT8xV5oS5
m5yS+zw2KWxaAIG82WqPkWR2BQbaRMRpox77bHclw9FBhpNXfk8VOniniv0P
ZiKI91bBh3PUOuD8yQdS94VdsQFOegDImGlqVheGG2EX3+tCv+Kz0EaXipiQ
QTcvt+mBJfWyyG1qesgIBGsYIr0uwWBo0sRXq/fvZhuoImcvDzwsNsMgLc52
Dx5Fi6JpPYGtU6L6eyxtq0NH/et8qSlbRKPR6F4jezEq0Xx8qV5C5r38VutE
/NCgQr3PegL9CkoDX6kBbCNg//6pZ+prSTdHg5KpgC2DrQZStqTIpOiN+lHv
bDsxJ+uKnf58ITa6gNFwCaGuyjaiMY8UGcsvC8wSHifeNDa0aUQC2D2d2HfC
TDygPT7//gaHRrmI6h6mA3inRgDUADROy49OYcLFZZ0IIGGrVvo/f5WIlKAu
LzuTMdfEs41NpGigrRBLjhRtVycllkhQwG/one+9Lw7FYgfvajrx6V1VxKRQ
E1jFQtgF9QDPelfwPaIribULXHAGPntM3n0lJGUSHITf5eeHZhVMTzAIhLMb
JNRGghNd4W2K392k8m+SWIMOBcl1SMJy4zNiY8TovD+KMewkYueQ8aHM94B2
1/r4KnldpvT4JOwEKjeD5M1Q2e/ynOKTtOVsqxOPa+knys0chsomHSC+Wx5+
Bb1kCyjlFUM/t6/OrHVDI5wll1fe53ScSkfzgbSmDiWrWCQG4Kfb4Y8ETGwj
6iyOg4SX93bmOFSwSMtKVltP4ljxxVtuKvreKs7+u7VPRNdRxCV1kqTlD3cs
NJr3CqgrEgul0kijB9K5XWXww8meZq7JBfru8VJQF9Z8bu5RAlpcDLz2vHyW
ButnTj0yAejoGHP2R/BGh4pKz4PLse0t25CCbapmRQw9dUi48+Eos5hOgkkG
0wfCoBo2TFYVBuU0Sm6gAMa/fAi/ZcTACkfEx9r9tzvImXGi4lcl2HP8NNof
HhAwoXjGnpPhBdcNGsMq7tcEYTuoYJafn3A2bM9JCyTKMNbcscyoXn77GaFE
Cw+EDlpU8pGeeTrB2HWKuCK33WOMujEG+1jZDsXdSGMkJ0H72b8OdA7GBBpN
jSD6N+tCglxf7TH+IXh9tnJWGDFersPdGhUkm0a8ZiWvKtgQkxIksuihLCff
xmyfOIfimOTYO3w+4WIXHi8gMwlwgcYF5ULH7WKW9gRSygOaOBB8XpYn9nzY
lHM6BNi0dAjJSh0FlEKPoHATBwF/iKB2JeOBNpXr+CA5JP7XqUqAhyeBNQQX
f6pGFBYCaeXzAJ0XVL0gY1VPiL0g8pzf7Iz/zAAjG1h7xEsYQmKuuk/J6Tbt
wUxMNLETwC6wrMTbBD0mN1VXGPJhHRDO+7+vOQTEED0ZSbMIFf6XEqskQODV
VlnbofhNVPol+n+euREpZPzDZF2+YY6cUWZjiF8g7JXaB/+qoTblk/0Y3K7y
HngfMdfWdfirDR0Tz4yGe+fu2zMoG7Hxtdfs3uu/Z5V1tMTUO18gl1apDvt3
fVqg5cB2Q/yhs+tBbw8AgjXn3aTJhYf5zv9pSI+/nGjvb1OWyI2qnTAJzWuJ
EYNZperzdLrrH1o12kxAujT0sSd7u6Mo/gniF3JBVwICPGPJzfawdmN9HVlL
9aw7o0WoY9sMTTumliq5pki1joBw5F/Lr1y/J5FUJtKI69cQWgBlWQCB/asA
52W3BUPeYNEsKe6SYg981TD3bBQ6ALn0b5VuvrNzySu3QNNtPb3fx68mEiwR
ufh5GVkjoeFwo9r+cPVfgPcop8XsHoi6nHHRl2mxOF52o+iD6GKmdz0Jx236
9GUzXNSTTMyx15YkD8rFqgKNkgQRDgbhCacROoLMR+MisBk9IVg/QLSpCBp7
MOXwRnGcCH0N5qrkFdoX1/BPdB/MKWbLzt2TQ6KMtjjA/WtpRXwyT3fqCSsp
TqAKYttV6pUF5D7WgxGppCo8nxJ8k2PGSoLqoNLlCpKXWkSyo2J7uaE3ly6O
PUoWx/URJzZGTkUe/+gpIbTWhTuR7CxDMR2+BzXAh+81PX/eWEoSzU9tDCFV
qqUTWT7DThle5VMcpBUetoqzFbjMX9ql1g30/GLjzeO7ebQROm+TYrykiWDe
hm5VurzZYw7VVhVCu5IJ2GjJoSPaHdeIvcb/wi4ouueaV2QnlOwy020hMZCs
K2HaoEmrq+nnMrJGPTMmMJ7ZwrR7640geg2CBGyqUFJYrCmgk1NNnAzLIAXi
xJS04vL+UGpUwkVYY7a/ifHlydLz1J+VO6/QBFUVrV60t/p69xiV4gjTVCT4
EyLf1EBPy9k+qYoApuRN/WAStqvN1I/d6A86vLMLqKA7xXiCYMpiuqm+SHXH
dCB4sqJVtyxq8xPQru+TlEzdeHVvWmMCgtJdWXo3qVgRXeg4Eo1ZdYPdY1Ni
HYz84DI7+ecdFzmnGEqncHAcRIfgqFpNYx0/9Z0iDRWOcbyyjlF6XaFZk3XY
+t1QCQ5dh1F93eleFbrnKBB5O75/ipcWhUrslXhXOPblr3z64oxTJp3rMewN
x62RNxu5MUsvqmc2AYpBwuesJCgTPfk5nS/m/WeTHmvkSLrrQXgrdO/p/fxM
AU6pwGfVBA3VMasi0+FQstuo1m3q8cQ2BJAZs0220hk50Y3Cz5IWMtnrWsxH
0qKOB0FgthhgXe4t2VAAOra6DZaPMsm0ys4XlFdF9h/gbOHZa+SX7pdth7aY
+7ZB9+Z8dMND5QaA0upKjlzX81QDSCyI8Xwz4auAaL9l0wRr4J8jvSD8CTOo
KAeNte1ksQMDy5Gh8xx0KL/q4C70aluPEWVNp+O5i1mFC4qJft8d1mTKs1cK
LMHS4Sc5NbJW7iFP9whe2RTsgAFzM/Ssvqx7SmfVzUX/Of9GUvmhiK6MCiGT
OBRH0RTzdICHABX+uRg4qe6CBiXMO4epCQ3MhWpzEZCBA0VZKop/poQDFR5r
HxBvA9/wLn9l/5MH+aeRaYy01Dhu/PNZTqNulkpQoMece3n3KTOaHo+WMSvJ
HzjhBD+3Gc9K9JrtWJ2wFXJRx9WoYqE/bs3vEs5eTpL6Fyc5+fkJ6ly9jp63
z9VjdgkJb2PveweRF69BWbpzdWBLZu+Ipiq2En13sWeTndb5Lq7bFQBtmS/h
8lAA/DpzjlzE9rzkq3Pnhb2SW2VUcpQLaOcANFvYdjXlQsI6RqmlVQiU1o+P
qVRGI8dU6GzORDDRIAE0jv9eg8NC/sdgDfx1J1Dr6+FBEZ6FP4eOZOpth8tS
FAj2qE3ZwzCXflj6jUXDl979ETWMdvDwQE1a3gTPSfSu7Pg/SHhZBU2CE8PW
CEVoVbPLduk5ruGuhGVK67NWZLW31Stg6/PES4H5DVyrMdxoWsP3uckKI+Fv
WsjO12E27+GMesvaIISl1nuJwYNStncsA6LbuhlhiaShYrqMsctFncj3wXNJ
k3ttqc6wXSiNUpGKKzLz6yrkxSiGLjicSSN3BIOHzjA8oevbcFjY9NQPLEp8
aJZHTf+wSiMsTlVeaKCB3awmWDgqDhk1sgBWpcXidW1yteXpPOzaYKQ0vnq5
SXqHPTTWZL44UlTfY36aPFC4RD2vI1qwZXX4ugnRDVJC03n/+UH+h2fnQ7XC
VsUmQBkQE4pq5T+15+gLUTm/EF2KPYVk9fvp49FeQnJOlSeoMDQ4E34Pj8V0
M5UN4dZGVAmqMZ81gIqBFDSPTY9ktsutc6gWHtd2TxKTSLMAmwGABYQKClHR
tVxwTKCCW3cYSCb77pBuy6qgvjPXDafNQ2doXPKUvJOxwap7X+mwqwp1ENTu
Bfe0hdXQWyoLSNc05nA+1iKUfpCyW1WVyfvX+0tyR1zYyFMFGsJQ2IeuWbg5
iMRa3Zdak7LOw4D96hfuorotmYx2jwIfrdCMeIeA8/+QyH6pb7gesBvac44j
lUQumOeM86JMl6nb2ZajnBpug6XJvCmcMQgicVVW4XrVirq01JKQYErNFNSZ
ALYgLh3lt5wm/8ovE0HulUEgTdU7TAYhyD4jD5eZObsMOnF61s9U8NM2OQJw
/RY6DNX3ADI59w9VmJngPyH9lxbzPQXGN6BWAZkMkEaR9yfJC5i+AJka6r2j
aEM+R+gSnF0K5FcJEaw3W2orDiASBo22xFSG+SD0UQI4MmtX41hJB9Bto5m7
RiylQz6HVtvmXSp61OWrWvh0OhwIXUZecPKMllPGNr3EvGOTmUMj/jMHNhEa
kF43RGRinZjcZg5JrnT75SsDdi8YdjHDFKX2fpPmKJaFox9m6N8CZGTtRop8
9iH0MsdZqs5Zl4cXjOErpgcoakF8Ajd4yL29+x+lxoNbxVsOABdJuYmVOPqs
HyZijecP8eC66UR1y7hqWtSPxQKGyW2SqfHKL40cbqI9hb4PSMjlYE/s1OmJ
51Yazjz8bXfjaVrWldF2ooHOzUWvo13zVrRQ0eRYZN4dUR5j9m8lKwX628b0
tnHzH1MMAdL3mByzKxzSvgyOoc0UtFDBrwvpJ7Y7j+fpiu+450tgPCH/+NUk
TwIZXz96fuiesqh4WOL6GSVDjXFkOkae4mK/pO4yUl+i+MIpWltCUlR/DbTd
ckALKg8FjRITSyAZ0Q9KHz+ZfnzfFCZYJCR8jg9XRLIuBkkV+fAKm71Cvbpn
lq3j7FlQbd+CTpCteXOvjDK/gPWBGunwSdx0qX12orYHocHRMfaQMxvzPlPH
y58xiTu1jZUKTHXkhilhKHA4+WoXw7bUppT4ZTpC0aEgFeHqPQ6dDaSwtJVI
b7z4H8h9V4CgNjkSDccgMpRqO/Qk+tVHzXBkGaVpFTXDWVDUoAHFXSZlgYsD
/BnhniJH4FiJpZMsNpXrCoP5/5QRaqj38o8//5nyyrme3M/Rpw/VNnBd7XpO
BLc3EZpPwMfimPx+PvnyUbUL1fvzfnl2+e87TfJT2CdXOKfxDxM3Iw7JkZGx
i2i3ci7MjwfzK+HH31ruUT2QKo7vwqtF9zCsb3tENAbhHsPUqMg22qpBVvCA
G1pR+0GAc3X/6pjP29lC/Fr1/q145qzRmE9es778NRJlB4EU5VWjteJXRdXj
46m4zW34otK8Iy5KOR1cNxxx3V9zd6aJqeXbnwz5udc+XwN3/s7dLmir8RGJ
6zfWARMixf8NLNGiGf6GELQpb3YKYsTnqfbEylagEaYsY2ERpo5yDkQL6B4w
dNJNObTXopuXM5sRHmzMoUFbmPTgtJYlGc1VrDdPlaeVoAK/VIEsEsizmlaW
QSOnD+LRp/8J5wZtpD9ZDtYmVXfQ4AN84g/r8JY7uO2fnfbJ2KLbxxn9rHyM
t9tPnWjoQBDbe+pDL9IA3OuF0q9pk/4BBRZzJHawLaCr6OzzUUUMCk3CBj1r
21s6Hl4DiE6rC8Nsbbscenv6otbKBr9MoYBtC9POjSlHdwU/oq1Xs4z4cc+q
5bFfFTMlGiy5ATvR3yH/rV06c2WwGf28jDPzlGn1b7e6+gXWfAdLOEvuZRvl
tLcc2QxaROPNRAb8CcZJBGUjd3CpHg6emEQYMpcUqWu+NvDqVpfrhKE/JWAg
f3go+s8640oOrnpqkeb5Bn0M1mXLZtvdzFNAbfdfxxf+d/VYcLfAKcjtZ7Pk
S1eDG1Ea4Mv9Jzwxx2+0qPlv/HjKzSbioZGU7KUJYg7mSQMYeBBDamYrt9jd
LtLe5Vohe3VXZmOW1WbAtJSj6eqKz/wR36rODkW8/7yZac86hzXuOX7an3JL
ALxtG49x4F4gjpj3oDgWg9QUO0hwsQmy5XSd46Fs7sNtqs2jYQJjftyf5PL2
+p1srVxA2+edM1XXvwb4PdgYuKGfGBQH5hUAJ9zbEVigIAUStGhrq6htBb5A
rbCzlfPfdz5p878sYf47KP4tGg0bvQgO2rC+M/3ESTLbxSZks+9ygqj0zVbe
FTpsIcjOZ5cGqRExIww+KRhcowCSvKQ5yKGa/AdQCEYsRnle+19cPvmCdP/q
QKUbhfBf98wq113mRT3js0J1tsrEpo1j4XmBJ6mJN+nh0/RON4QKzEz4VXnP
4ELVJTm4YjXyOWM98OLcGUnp4j/82vmN1VKSTnS8gfz40MAimVCVIaNnynBh
3O2pZ/hiMQ8JNHEw3dzHGB1xh0JnPo0vPDIR5YQqJtjA0cj1OEGW4cI0sCK4
vP9KusXym/lEbNaI+Gx4SiXO86sMxgs5CN5MfG0+Mg+cY6FmGPieJB04BErs
jsUmuruo3xe6SmZ3UK1Tvik/e5j90ZbiWG9Xebmgk0po829TeJ2KO06i+UGn
mmjtkO2I35DVo9ZHv+7OUsNMwjFHDk3+abkpX9Dl1IrJDpMRLbgKbv2j7rNH
rwyolDojstz+zydUcaw10ujmZbvoSfDa/QURV7OHbGRQpCpsaA9G8HTRc/WV
ZZr/ihU2566tGi6Jt/XYK+wkY5Uxdmr6AWBjCd94EqWLNBz6KCHpMGVL+xkV
IDY6olUZdyfOMoCIAdcIgstu80JRGs0AaQodx6Rs/E9Bo+43Upqlc1H0HltV
ZYbHzbM1edETsDYrqOLuSKd/Go5PDCoBj0U3AHi4KB/qQTVmgc+rMTxIwVxs
kU3wt86VQ/n8f9O2h1ouSAVw/NY3M0EiaUJQkEbjBmWaJTd6TCHPUOR1aGXN
hQS+dx1NtgtaRgdyKBbEl/ps0EbHN/Fhk9W+3mLDO0k0Nz/1HQgA/EpZJ9+i
IFEBsCi6Je/ihIpE7C9lk1K5Ipp79y1xPSt+7IClfBLGqGQ4KTd0UcJ9q8pY
L97WqTbfnnfDErtz22mWMZZkWRiJCGvER/2VttOVIqbBFPxXSt76i6ljOJ1T
OpAuBOdpz9WM+0BWxez6jPO4Y9wDUeImPdTj8yxr/qWmdX/wR59J6U8MkkyZ
TfkEvYD8eYPAmKjSxMV2Z2JT0C5zdfVGtkq5NiNEo0jt8w9Xep09aBC+bErV
HkOqbAVfBUnDA8wNJ4aIloMx6d2kxStl5FBuscV1QaP4HYSjedGuxfNMXgVL
Nvmr8QapPnr3WVylqWud87JJqQUwqT84n39d6s+43V9dBf0MrLcu02n4OYJU
NwcpiiuvoqRzh1tKNPSa778spwY4oLdXVIEYUdT3HZ0x88JaAdFSuRL0hCRs
3E+zn6WcxPJrm8ZL69OVzm7O+QlmTL6qllazHjaVZnmnFSBZRgVudHVz6fqg
iNruq/MCylKkH29y6NRsoXJXPKEBRH42TOocei13mVNupqCRQjIudrCjfNto
UyM9+0+utxyvb4MQOcTY7MEmMkjGMtIFWl1XB2LzWoFT6MigAKweXgrsbxOT
MRUYl/4U19fbYmHekGxnxghBBOj0SZ9twP3q3cPOLiFK9KMyri+rcs4tPS2C
DGViUEGrY6FhgwIBVNxLms7gniobMbBQjVz5FipBkf6ylh41Pn5/HBD1RHXH
P5FoyxbhXKCmE7vR0WVtUCyJ91FG/ABqoOd4AnojQdR0Oj2h8zt7aPteAcNy
FMsRcSdvo5fzrLlfrwzw2L/IdzrHS1SbVFIT9W2sp3YtCkrIeaEVi6292xz2
Rzv8gUp5Ew5/DVrxsVDpgIIzFYnBud/A30MOMgmhlLyd2bgKuxMSdhiEaiI+
nNoUF5Jzijcnv3DmuJ3fUf9eK8lU0jV8WR5VhZ+PnfYgIzRpj8Uf3tlzKbZl
BVE4Y5zikMFOWdG6tVUyA6tYLkjUzZ/ovsKPgk8bGL4kjMGQ3YliDta1DrxK
oJfTZjwW0mrynKtdSdk7Iu4H62aENA6uJiZyPUXGyZjIWSLhNk+lRsgScPJx
NrxXtr85V6YRKJRSTGtdVVk1Ec9R70ChoYJoNFMJt0FhvwNJGlIQIyxqaMFB
+a5EURUaXp6Sz6KJQLLqssv3HorrDgASxpAtw9dHtXYukU44xFADeFIKKS+d
knxxQ+OlM7seyBrdtXk9tLl5WggMGL/TbKiDgDIkQvDI/WNlHWAIkJyiROkq
JK7IxfnYafABXcyunbFLlCm/CfvE/onHollGsbDlRS7oFZYfvHDnj9iQ34HV
TW+KrZBgZe+MdoQKKN3gqsvQSkwsYM2qQ3d3n5UowFRK01FyYTIZ7n/mWj51
SW2sKGFNs164mLhUp88o4u5GrHxjAdi6Pzlz3mcFhDFl7mI7kQ6SjFGwyfAv
yPGa1OBLL0GxzvoG5LGc37B2jDCpEUM8UJF4baoky0SuSb43Acq6TRMXgI0U
rXLG8w80kDfBbwAmqXDuCjhI6DaYpvsW1C8X6ZJliRhEww0xhZ2gywD4RVgG
hIm2TrifkFyQD1mrXRDqvx2JaTrMHb69UPRJsM+KfJh8AbMnHXRyFAky2XGl
N9itGVCAxedaZ9iyrL3nYz/UqD9DOR/++YA+b7vtNvI26KtF4GuG6r+oyWgS
w04YZXbhmyTaO5I/J81DQxVvCDrqeWoh/EYzPCFrnyMXlHiD/nQDpXtoUuy/
pSn/t2U1W9aNxLeviIJvQxndoGuEK2DmPco+QryWle/nWOtYtsAxzfFyqnCk
1IsK+YlIHFMhQCOBvRjotYp871GEWmDUWrOaespiq9VgOj+77+FB9RAstdXF
TWuXFLLQohWIyu6lFpn70iyWj3znb2LqmZpBxcxgok1sJg9kul8mJMozZAnS
Fmeup6iaR501b7wgL86s8qetcNmz0APgvS2sfuueh+ZUbwoFcRLjMoJnYX/6
7jf98/kkN1/I3Q85jvks+p7N76hfC+h6a6nywC6H6jSHAmYQ0dToZr37cY9I
jmnIS9DK6ttgOgT1JZJcDOss7LbGE8q1y6h5O6xpo9Y5c6KC063pijw500eV
Kg2xdVZcxmlfRY/sOh+zvSgunDBTPAFeCZuNgDfNttvDfIs+SUCdFdC1V6RV
nPrE9v0OzKfYXoSOFqKyO5q0VQfcCwouw6ngzLngaGqD9tpozl6pvVfM0O7t
VJQDr+WFgc9KZgoRidZ9qPmRsGNs15y4hQvFsIJe8LyH2gcp6ta9Ji4Q1xMk
MRLsM14ClKaIvvSWEtI+NVjSOzb3U6UW51MKB20X3ypJQX3YprCDJ3LuBITj
DKCuzQ7tpca+yCfW2fv/7lkkg3F+snHCp9njl9oUG+QxN13UXkJzEDJG3RCq
uKxp1uVio+nSo32iOdlAzwJGmBC6PrAt82+r4Jmf6v/GJQu8sNOelTJl8W8V
rj/ENje1tA4WdnGInXXjAIj1i3Mh5kH2dfCxFx1ctrdwjbqyy4Qnp2G67BCu
ZSJkTuLD2v2pkbmhT5hhUqm+YKvDnwoynM6O6OaTNx+4KGvNSyjiDXvJQV0m
jg8vhLy9Duq4uTVo3kKHDXHX0vmn9mP0W+Hfhm6LcOOYyjAZc+91OrjIRi4H
R46elH8DFmpxzHdt9Af31SgYKTgfmfJRRNS2sXzRQqhfn9kut/Rjrb0FxGMg
z17jwxu5KUL1zmw7ZL4N1oyBHvGyVFJwmgwSfnHZNlicPdcjBGCvjKJ9oh3V
InlnTTI6fqNFtRT4ovNYTUyHn/Jij1XvbQheDTjxpUfI0EwxaFEp7uUirUUh
13D+CC6QdK0VaJhmI/y1O+P44OS4m+6zCVN9ge72VBQRZPqgsxEE5F6jFSNv
5BcdhOwLrDnc5WMWMv8mHW3ABrgHdiEVAlQDpXf2u0M88lJ13QHOEDj95qIg
u4rOhu600tOeTkxXso/wUimmbTcmbSukOjF9u+gduRI6Fc0gDhH89NRETQPe
UtW/r14KlRie6IWc37PDJd9k8+d0JZsbpCZPkVc6K6so7eHx2CU2eKKlS0oP
dccAEeoSRgcn+VL+cLhTTElSPMG5PbwB+K9+JkxWLpERmtI/Y99NKn+JEius
YxeyyRzRjXPZluiLZbi3oyIKxMT33RykJjvJbOHno5Y9/iex+2xsO2xW9fAu
8DHAjk9fW46UUjW+vP+SPl5ZwsPXnjXFvCVx/x9YAGwrxM0jVpE8FFDWn0CY
I+YCZPOn2ihxXaDMneEAARkzElCwAvq1+EOqGrYNkZahaHLwN51Tv63zvUsT
V1nDc+0mLAG9zbZFxAcDaW+S9c48kiKEv7QltAf1yFkAhGo6+AcweDRlV6iV
YJ+5KNMwxhEz0ymTzfmcu57qgfXVD21W1USoz+25lzLjxMg1lTob9zETt/FE
0emkerkXvGkh31fWuJliqYdawUAkxzxqb/ao98acHWoEpPkxEr5adynFQ5mH
MKM83g1jo8h7kmuzmdgaIy3UGM8bXIL575YF173fqMD1yZ+3dNWmHrD1uGmo
Z9aY3hTse3pdZD/v43bukw7bGsnRu0RGeP+YVv40DkGILqxI6qpn/bh5kcHS
0ztz+NmKItizW8GUtkQejW096uB0H4vRFNZsPjnVrZMEgUaB7UMPtSqNbCsK
ddbaP6TTO5A4BXFpo2Hmc+WfqX+xw2kROLBM7eBECPO3kKY9QxtYFaIQ1WfK
Bx8BluoUfUIcpgP8VDJEPhzv1VKStR3xHRe9j5E9wtJMrbdgh67YB5+PPZ44
RmIeM2QTpktMvawn/4PiPAAtYMviS+6OY/AnB6mbo/yrA95NCODVvQrJEET7
Dgu9hWarTsT3HITfqZJx1L9j732eu0VAruXxR6dcHN+cZM0zbtzoMrEFwtbS
ejsKmHGmNW7TPK6DW/I2AykdzVVgnPhoEn184sHWt77asCSujwtw0hZL+8m9
Ic+5GGkpCtKkzUP2gRpJ6V2pS4NDZp5o8+1DCaXCOYEwyBH+JPu04trq0xeV
oq1wWcL7+a+8nKhI2Ta2FzJXfe39+B11iXgD3hQe/RQL5ihSTCbKjQ0d7Ac1
Cmaxh+A+P3OtqNK1mJGNKEiWK+VvSCuk04s0gor6QM+UVSLScszjaOynVpE4
0zr4sUMMQozPB30V5rmB7Zuh0LmL8R7McrPVBXFCh0H4+WjPDSPSrMwmb02W
y5sB3gZ3J7IDFpGBZX54ANC/m5/JvJEyuHUGC+f63FkxrUMau4aGFqQX4ay3
fv/T9aC0p5toIakAed5gjzPWo1Qop0qr0Qp4kDV3awTCWfr222pwNXx3KVDZ
mjrvZxP2BGCMu+PGTCl+ePJ3TIc4Ld5uAZ1fdjeCrvzBBeTf5RT4iux0bw6y
baS45pYqYMihtDB2fF3Gv8BJCIpEA9qR5R4rTHfe8ElGXxDDT0oqftzEtj1L
0HvY2HraBPTzaPmszNmwHQRvLSrpsTOVshgTq92D/gno9m+pCSAosDvKgTjf
gT4RB9lvDisyRpCOMmK43VTcE7EhE78PBH5+y5agIFPl/lVIl0JOWKy/VILc
IAjM03cAx6PnONEDEJrBsNk0sLtM+c8XQvIj/Y/2Ln/yyZhENOb+TNPRseUH
IoeCxAqB5GNuwh75ID+WucfLtyd4/f/TG7JE9jCls3zyBSWpOlM7M5oe7uow
AK44MBEKh8nqJeOq0Vacru7r0Age0WegUwSbLf7fl1zJs6292fNPGgYVhduz
YpTBPfTxpY8GlhIkJdNXynR1WDCeNJZELL7aMQ+5E6GOpd3pwh/BVIdzxy6A
NNduFOmdTu0f1ALMtfBTZ6U+PbDGZ7LkI/1EHuBx/4DuA5u+HvpnobnHWoN4
MmrXOI5YVcijnS8AMjh9QJi+xuaxOOqjez8/NdtbfCO04tJkHEk2fFjhOFHc
Yt9KUskH5m1WbcaBP/FPnD5/ZpWiooUtfFOXXzsa1vHjDivv2MTzDFQVNFjQ
44VqoboiTZwaOYGfLOEgmq8+pPjRHpdPtEwaL+Hn4GIMPK3lfOzgPFApXdkq
ERHAg/VyqHk4ha47+RXGcQ/MDzDbAaVx+evX0NEGNtsvMMXD5UWsUbSnlcAc
5p0xg6bu1G7i2teGjjwe3DmvKKvVWWE/s4SF+FpiXCEkwmrP3meo0BcIG3mS
3pLoo/bc+SySsD3Mpk0yNwPgpH7rrGF96CCWAu+LcQqjdi5ifZdEXshIfXL9
Dh9VDSUqEITjzwi0nuBZMjGWnMb6uJU4Wt41OYbIFOlGUxaMPcEQJX31C6Jf
nXlY3xSxp28CBtdSucZxxQaJjTvKy4Nz1g2jPU6sz8QM8jeICwn4vghfUryC
uCy2bBOpkdpDKzXSSTThExPcmzGoMovjaycp4UqcYTLq8tWxirb6+JxID517
4VB5fqLX86oKXfzf3MLKpmrpvvu5Cb2hDEzyFc/0wQec+UZGLEKEgH94i+FD
OLQUBW1sucEgOOVWPEeKijfDcpIEd+Y8TQ5VpKEhzyM65y3N96aNLFNlEjiK
Hmsttyq5eZ/5Pl17NL3rZHmu0w+FkoMhdAJQPdLtRxbmq7DFpvTO1YNrWlWr
fRODHORt8OS4AvqcPiBDjOZwXHSbOqNP87LuKQlCGYzWogrpl9ksPPeEhMIT
Y6DWD46JGvtEnNZpn8eDwgDzVJrp7Zck4F8to9SI0biV7kBxVR7id8XJ5roD
EXmXfi5kC7FGYkKIw20xIYRPs5toJa6lkbr1pxh+UEmTJqiRDt6cW1FoemYq
ZeTlxE6etjK2f5ixZKjl+EMQR87sl7qYvziQWdM+sKS9/IAT+MiXv+CB2/VE
wfnLlWvAZnzdTDbqgHDwZNtxmmBquf2sM29hOVOReOgmOK0oPL2e/J3QvLdP
t/dfOPEt+ZRXHNHQHNcthjg+ONbSFP85S6u5590diN2CNsonql+Rxtb6HGYq
JHPouA3g+ueWuR5oVl3emyYooY2LWYQWeyhZ/RZiNsfwiz8QXP2r4aFqKxDs
RNSS2GAXgIyGzl6ikUBEkErm8cUiZFXe2+o12rawqqSJ5mfzdzztdvi4+TPt
XCMyvV0IT/kouUAFumzo4ryYsj5hn/3DQ4UpZKy9eDEq4bxFa7NKuejoLXwQ
A0YMwFG94tFojIE9lpll4BICe4o6pG63qnrLcL+yn7OsGrwAvpOBlOAOr/4P
KmxBC1AwMEik9qaasV4wPQsg9Qsjey4EV/WRbGe02h5u/b373iFPdqScuYpY
WYlegEkCed2Q+dI9b/2sbRUaSiD4Ac99/MbUZKRROstrwWARgGQubmm5zAZQ
D6Jm2WFScW89CZ6A4D4cOyeXRSQh+qNhT/BlbfTG289IsOvAlTOHfDNXCpOV
KJN2vOHKyoUSoZijUm9/YqMkn8FPf3Wu7fO+aXZF/nHuKA/x/pNvKzBM9C0E
qusIDPdMoEo77eQ3AvXZ64lbrCvF0m3VVHKMOsUMPX631/aRpVmukGZ/+G+C
Ar8z1xu5nvOGsEHQEEBNNfhBcZt4+NlygJZxeq1ZVldgKW06v9jIxiSES7yC
OfGGv0AG1peix2GyL57ohYqXDTZSSEkG+4ZFUYOrHgN7V5+L3ZIUpyMkzQP1
apyeOhIvC4MWaILPRw2ajFfc6e5gGMWRICJVsNMcFphsFpscmyQAx+R620KZ
zPYNh4n/Rap3yn22jTDJmFnw2T8B0Q3gKXGy95jatQmDeV1gK8tdb/X4s9wD
CDrPu2y/gMjteYwpZfDQvUstyalip5kAp0he4+AyAVca0gV/+vLTnntTDOAS
Zx9I948S7AHSqlLLyZH+l0RLM7TbA+NppSidijV13RJ91gz+R7pn6qBD017A
5I2ogPj/Ayi47XEwBMiSX677s71Bw+vbU5uZFTcrchGaGo0LmxbM2ovHYwP2
abu+rfTYQ9H+S5kW8ZFaXcheXLZxSyyb9ShN42+o/skvHVPnnAd8xqNCMC7a
wfOAWy7KUAo5QqPO2nidmtMAwRVaayKlrBoab1qBDmgDP0U5+N6xbaOXiIth
Nx/wj5G3PvGYrVlAfxjSUU7ITQsGieYWHIxxwmmbKxrOVoQ1+IAYXZqoCTiT
iDu1UWXem7i7eITF9jPHE6Y0UoDQwYnv3usxjvSTTM+zr8FoFhuDYDCHZdTA
vYFGfIpQLAMjSUwIDdOyijMsCRyJhGqQRVgYG8vTUfWhD98oZw76Su5Fwfmw
gi0EvG/wRf0eWnA+Kfsxzdpv54UAu8IPW99V9YLxXvZKgj5Z2h2XVXATl0mC
wBt9dQuFE+P1bRaUa2XSXj3M0GclP9DLLaMUHVnkc5aTZpKyKYGFIfjDGu4T
12Vn1fh3a+6E+6bvoFvXNUWrDRWfy+GpSJ8FfS4sq8AVpRpHXHFt1aP4q8XY
EoDvD28R3dncGLX3iDkYKHCmDaDxCFyeKbdq4vmF2hiMyQvUWVe1rGc2Tgx+
tJYa9OJ3p5ens2H9IUaj1uJm+p6PRjzoXjv6TiMNPqniAdb8DL5m9HxwioDA
PDD3OLBhkGawzFNAG6rA6eCAzXfcuYIydk7XNfM1+Jbmi5ua/17HKW0xuJY6
a1NME/4eN933qvt0g42r2H0XbDw+X+m251/sdJweFtjqey5mdCmyUERR9WZH
am0Aued8kMNlVubdTSN3NC99PExBhpOlurnCHVtWttbIYedjzn9E6P4dLqVN
w3WIQf1BGdMb7uKRfDBAONsybGr6zoWeUm8658NCewi1NJfOHF/axUD20/Kj
ZQGw95s0/Q2KJ7qObWvrO0JZmvJVKcuQhsLFNDwMQzTWRqRUbiMiGgBfer22
PfDNxQ3FL5vzLoHbMD7T1Vsx7hSZh5oCZlexE9hh4N4VEXS3XGIZeYX9fEWE
ZBQFlcgVhc+zjxTJjWb7Pb44E9L0UxqA0OatLihJdtqpzwn7DNm6Idop8hkS
wx5KsYYbSCZCcNAEU33tshz9nz62mmnmxS8k6rxqDmqVzMdCcCumrB40HB+F
GHPe4sKjQuuQeh6WVzel5iGnGAHH9B/bUzb3Yg/VXbHlw0roLjeAm2ipj4YF
5qHy8c/8GUffICHRSvoXzegqbAjC/8yG3PUjWHhONLJ3LGN9t1XEkUelBqrE
7KGLYy4aCzv+q4XL8qAHMcI4EaC+jBQVGDcXwtVa4horkmjrvzDXF1dGEPgH
pNTsZ+cG5TxT9qxXGJxxId89xnIE4hp7x3x+L9ceKuP4UvizQrHKNQOjp7o+
bMlJwaLO+uv/hK8TtcewGlKmwWdGlaxl+qykmm6hLeOqTuuXVG/ItvpyhJxe
21mtrVp5cr6KxO48ryAOe+z14r3hMKWLdgIfbEA/UYKVbLLP1ATgocqIXH1Z
AZ9nWzQ7kbCffd0CijP/kyi7eMUkoqd0YxUcDDEChgiR/Wf5/ObzEL2PbsrO
ecNv/EhHWy+ggRNF4bfHQra5nhEVmE9o/3Hedv40SpfzlnSM/YNfAk4JfOF+
uQWL//RE5ujAqXyL2/4K+eDmBbHG3Njhr13OsL+ImXCM1m2QdFyMVyCHC/M2
nX+NxjlsBkhUUdKiS04lJI0SCeEJy2lGq6VZ1nV6YBSg/LhIwkW3Ma8ySfqw
rAv08yr0czfaz9hc0MhuDyJyRj0HZXXxZIGQVtTPCSj2Ps0X0a+hzjmd01GZ
9f5SBHxxzdLBJeLchbY5g+SmD+X4ZEuDaLxt5C5wYw+5Ga5OPBY1g6n914jm
G6A0OHqcqFg1swHXQt68pRijZOqLD8Qo3zBwvITOCWQFAaRrISQNw8qFTxvl
wipPMcHxCiLfgxEgsib3eaX+AaumaMea3f7i1Aey9PR7ZDPJO44vZct749wA
y5YC5nENlR+GFVLwh+h/53OPzacO0xB0wI+oFmhPgbNDius5TWlFK0yJ/Ycb
YmVDC8sAB/93L9IxherhGCpBnG3vlR3wiEKLM8e4VCmy1icfkFtdMUFnrXAb
rT0Mg2oOSJQHCYZq/Ca+t0oDf6xDSXZSbQBy/jAgD5oZiAsQk0qzsqa0IOVH
5EUMWLatJstgghUOswm1K1B33FYhthfZyE9GY3vycbkgIGKEvUv5XFfXn5RS
98gq8prBIQWAjo9T/C/i0geKYIuQnOvdkvvce/bJgrQBgG1Kt4Ts34dndKW7
94f4gf2aC4+VkcRX6NkxepnOuiRuRGkO0Ah0npSjZ/NmPa3txEk+XBuUjUty
kB0275wvQauP8Q/sFK7NxIrejvgImnr/b0fiE0qTXpySs9lDkXa/Z9wGcp7Z
AI+/4gvXfZAUpBhmeNyVvbhyzyTY7hXEtvyx4x+mPf2oAIQcHJwZshzgaOmR
qvniW3THlguMCBNiyW6l7en+1iwd8r+cc/Mqr2QVsiK0AzHW0xT45EuYRHKT
UEh6lFu8e2mvfquj2ryrXmwaVttP/JAx8EGszYc17FXOa5OvgKgkMN4fa5nB
QHNw+lfyQ1H92D7I02Q/Cxmma38PDsDvHQSLP3BWGxp0yw2avslLUcHsdFNc
/kxp4T/Kt7jnVKj+8AVy8r+728rinxsK01zv5bl5amVh0O+3/VjOxUcFNQ9D
oKXQ0qWhI1mV7Eu9uMihrzKLUOiSwPYGE3YHshyXAWqofAWjNBH/wgjYZk0f
WNnSEqHin6iI9jDUH5HbVGBYj4lH4I7gOyujmM3dKqvSmkP/G0XneZra8J2q
/qrsvOzFQi26ZEk6gB5t5h/WV9s0r/JtIaDWz8bcT/ZNKrnCzTCW40MJDokG
RuLVirElGRLRQMJUgui8sqP3/6aBLSET9EqJcTNwY51/SXw8Vs8z58sy/a6l
Lf/PoBjYN++wsJh/BIhvk5iMQ7miCWEfkooo744Z3AfDmDepTKj8BLCnmj1n
wTX/QjFObqyBW1CaP5bNt8uLpBRGS8jDDGO40ppDZG9tRTK5nF+TPrXUMf3R
2eGm8e/uQtEs1ZgBaLlNFxBnXAJMUHENFzgXsak4oV/BgnoQLxiX/FFwIoZI
+W6y2Er+v83xRhyF0BDOTzNYX8W9dc4bvVpIgZPQdQ/1UpcF9QFaiX1FYw5l
VAxBEm2SYd29jgW5R1OfBhfm1vjlcLsrcbej+rHKxucvDo/Dm0hfKCSjkfu7
1VlfoMkRnz7ASWoqL9+UPdKMgSGL2J7NYuPO74AKU5ypqntHAn1TYKD6SnA2
8YaEeox5qVz6MXvLxyGsu3dP5rUJ95HDpPDaJni509CF4Wzku18O6U5BLKtr
+z2b0VjwR7PY2eIezeIg/7q4E0McP9d17BXJRsT1+nTY3qutso7DAzxE76mP
/fZBL2psaXTdNYsODpghMpkUzy6vEZ2w7gHOObXVPrk6OSInTRI1ouIoQgVS
NXEKB+qCrhsa6b7iXefs6RXusK4BIS3BvQ3DBNYfMu3JbhMy9JFFVSy8N6x0
LfaD/qxAPMWS6gKbNLY16laVKT7b6t8omSKHsIdo+B17nPrroXnHat2gjUHi
EoHFDWJxT8cBHXsFUsfN5bGOEwThkErDXtlZRavTCRsu2cg6CoM4rr9ZrDiX
R/q+Luxeqm9jJ/WbgLzuKTWuU0Qv5ecS2nz5CreSb9dRYaeqBZfz0odGhTJg
nhwH7JU7OpMxakZ6fCxGA6LhVDMMe0Fp7J6i+yH5Fs0FxO4mjyeuqNQ64baJ
qtTihfPhLgr3FdP7Dn99/2LWt0oQNYm/B+qPFLRukRcXmPapgPLiNHRzxU0y
6fCnfNS6ce5UunjaHSxqj5Vz/8doBHKJ4ZGRd8HC1u44BA3kuUL3VRu4YmLW
fZ/+KIOPVc3fj8LPAq0MXMPQxdSivBWlQVMpq7z8+VkALBuy5MxwFi24Z88n
wY0JRcmmqtes9Dta1fzDGcfwgmgsMwQAbzzwHcLXw9AdytBmEDabGdF1Q9QR
O8wJy/mMKnzJyEIJ2wYyUY9jqbF113HO5B9xHSuOh61hkoHGf+7JyBTZE6/D
GPIBTqYl2+5mF+OyV/THozMBN5ori5PYgMSTRKKGn+OiVIzxkeOLodZy1N1w
cJZrWO8qn78T0c+//reO3oxct/wHi0Rirz9HhSvfKp1ouJJywj02t8bWEDZQ
77w+bes+8QVop4BV1dCRU3ohjw6QNo2dLILLUaFfeBZIOpGDeTvyPTiD1F4h
a1dLU/p/vRNaxE/nVswH3cPc12HJJmrBXY2NYVTo6lxt1d4pjnUZPspydDkC
b4HUC1SGV9V4bupWz+54Yb8LkCkuXfMBq8pR77b49Wf+q+RA/XdvdZ8y5XqB
7q9MiHoUG2nMIJpbSl+p80vuoCzRjjGkYnYY3kynwNPD5Tg3FdCOKYO0+4bY
G8hOqKymJRiAOu1RU5stafdlmXxoZj/tT3Khb8EPj91rNozhcD4Z5iYTN0Ly
8IeRFsWuAFKvtVeU3uADZf99hVYFiDZCcB8XkoBOW6LJhLfAyxhqs3tY8Z4b
DgNOfwAnyy/FdO3/1iHDeyw5MjWsiknzUP3YkCWitFfa/wDUk7UEJx0RTIKW
SNIkb9qSkcJrDfGWysiGn/NaA+KTcYGFHRLyWk9UKkz+4nLR6ljP5eF0jtMD
Zz8imITzTR+hjlSoiQD+FyUcVOC2hlaX8SNEfQNR6G7LoxYlov1py3QafwRq
R7lY9dc9NkvNntUDUuOt4FoIJ2YLvedbf1kLa2NZUizmE9AtuhYY2x1PODp4
9kNACsM+3qWeVfK8Gs+2tVD3XwnGs4Ws6PJcxpprdgm4gq/sFGCFkq/Uz4Kp
8gqUI9e+KJOtuKQhHsVolnKJT9l8aBT8wOeW/AVmfmdwiyjXFRwVTfaKHeR/
EpuJECdTpL/DZgOtZ72CUINvm1D5bLl9tTb9qQ+GUsiVvhcZ2Y8wmnc7zuMR
iATD5xMi2+1te0iUiSq+ZEi01lbPxebwheHDiP1XZNGkTE1webVkR20x+Lu2
ifrwtS9d7PmneLmv+/A0FJ7Vmh7E360IsHqJyqR4/b5HH9fP660Yc06s1ULr
99G6y/qwpyWa9vgmtlJ0stkiPG03dnGdjerjqh2IEwtL7Y9BIF0gdVeh/0Oe
8r1VIU8gIs5VuJEZyKJk6ojCDuUKL4/dhr+Lt61B8edh2TCs37Ax+m+4wo2c
YyDBa6/zyhSJ5qx6MIvAHwQTmTaBUu6si2a3/4jUBsMOBLCvnZPCBd1bPuaO
+OrX4cOUTuC3cF8YP6mR8S6t67FlhJqPDs0sHF+aYmo6RziOvcJfuJr8ZNqU
rLgTlvGIgKTIEs53gHQfxvMXNTtZ0J6IFb6y2egh4E/87WUxoaxp227LpKfz
WYysFeqHtb5NB7pDeew7BiYGKRWMgI4vY/JAcvzYqLlnLoMzCD0dsjogCDL1
+rxW/ttglzuIJGIQMLIkU0BdSDwSipFAHcgm72CAmJuzyog8dyA6WgLHFCPp
XOM9WocPjlLTUWyymtwIzGW4Sm6PWLpR9xdbGes/Gq0YJ6vwrlDuwq7YPzgG
HMPoLe7My4fecPPYACb/Q6ew2O6tyshPeocKOvmVOi7IZ+WJhznX6M/ywCzi
A1iiTEpfk/LA4Ni+Z3syC40i0JpQsIPU6k5vJbYy0dTW53llvs706nA1xtcV
NAKs9ix8Cj+kVwJ2krC3N4BH6mEQALMp68WJa/HGo/w6NUYqV1elPoWCCckv
HPrcOhwJ6zhFTdaGq9NrM+d21pmm3q6d/Ed8yRWA7ZxvgZiJ8TkmozffyEBR
nNS9wW4VeZoNB7Ne92U+1eBbEk2QmuJ0NtTXsjHz+t/rZjfermZHyyuqKUvM
znqJsKWLc9J+1a6DbA/EWzkUfD5x0ExeleY1pLOw0c/fenXsFZJ108XYwJD/
F9OLm2+866MDyMuSFikof7BnFQgv5xs95DAxx+WuWXa4w52kDedybiS+3pjO
JqfywnzMm6E+BFt6o5w8CPO9RkfFz9Iu6rdzHi0lrUWQp4ManIuqNM+yjYQC
Hta4Zp3F+UEJ9927C9FRR0iq3ov7tbgTaLBleyau0GfvcrmsN9V/DXby3rMU
KvZRQxxmcb5PJ6UUK3atU6GPqRwvFdkWvxYvRJ8DK8jj6kqm/K3gIMXv7R4U
WCS1kL2zgnmFpusI1+HFbOk85ug5tuoil4AInV0yxEZjmEk2xA0i08GK4Hyh
5iAGPlrJwe37ApnadVwPelglgCW1CquRBVvjc1yuBXdZOSrqzofxby86HX1f
oHG6kmiwZv1jGRbJRRByMZRMdg8SqtQoyJrU3zlR+WQktoSs0Q6zDTe3OY/g
RnWoTD5gcNKusR8HfeJ80pVClbLGl4hswfYKUkv9KkfyEq6UGSEVO/JPJuIH
Uq4htTITdC/S8/hQP9nJ7mFVS+kJuf9+xDMbwBdmcKkMbyTrFFGSUltJx1LF
hiqrAAPoZ5YHuwi5fZz7T55awYlbIEoVeI+R0hF7zsdjOlOZie/57L2m+peO
ontlAgP7dVGoX5Fxdjgpk9J4vLiSzyDIdLipKPe11/kVUUISWJDogv1OxZgG
HR7q6yF6K43rItlK52HGSCtwBoYwD9gcVBJfY87eHa+WgmFaVrdJcATwo76k
dLP8V6jWvI8fif4I2kcJX87xkDvbaEFGsr+TvkA+raaxo0Ob9+Ar0h3XWSMP
0wHrabjCU7vjdzoEzHfM6TV7LuQw1vXYOkh9ixQ7OGMLYW15ybz+/XJGHlrG
QLQpp7xJzS09yUBMXxIElZOa6ROgB7GQRkQiGr1dCBKMur9yPtdqWrWI9Yda
V1qvz1yn5iWaWfv/v+nE7CkNpcb3Foml0lFc1Z4fnqqbRiDe2LPayPtvfA6u
WjPyxujkNrXUgqBZtv5dI6dCjj02crU5o1KhTCcfoYeMUHH8wtjygRqo8Ziv
EriK4gAQ4Y9ECT4N1sg36nPRYBn7EEfMMtAslcpH3eNiLhE7bfLR6EBEU4YN
bUemwRvnctaThTY+WryjpF+0vjUPBZ6CC7EWZD7ZlOicAnYtxEJs5zWpWb87
edzx8VWjaywXbMrEjaAfSmR8p8KoF0oqp/xj9wgioNm1EYYjHer8wtf7VuTS
M1azXSPHdnlX4ybX1S8TXxY0rINsbHEVVgZn9bR358yIjwYNHxdG6fKra4XH
wnKJjK3NTIgBOncfFdb2LqIaM8thZP3Zdpm33jUNJS/cGL1MmkMi03On4JEI
Zv37J95Yjv5PzBu+YJwQPgIxFHJdSjLEdDAcM4UKFhsh0UU3zD39oFg+8Kfv
qsjKa29fHv/FSsl+xXwoNJKsfLobLo8bbox0MiCF8Lr4a9zdpD4ClLcMuidT
p3sOFbiMi1FaMK6jzKlQ9wkc1QUXWXqU1iPbytrjig0jVa9h0FOqv0Svaiji
hSB/DOGtUfDFkqvurO0cdFhw89eWy9Tdf9+yuEW0c97BwBdw9Fk/t2uaQHnw
nxyM2RthD3Fxsy19JwaOisi5GHPlmmQ/iSFxt67hwUBI1dHALpczsKVAT6t6
6kmN2IlFWIR448bts6uZiwzulhtDkbUQUj2ZLJo9tij012uqqe1wSNDLc6us
WPQirPd184OPqfDeTUPPhg7qTtqmNtXarH87Q0dILdMfr76/vYtvMCPLgrHP
1tE8mDOBbbH5jKoc/HA7oN/NELZLPcdbuM+AoTQSwBJEiMoCv0Ezw26wAiOL
li0TiL3T44ua6CpTmfvOxXUfVs3S1KQ9FSb+9OCrmqtdROJkZBp7M9Lpefzw
fYg2wGwpJnGdkBdtxEcQG6Ar0yKlvoe3Tq1m0wNL88ZsktIpYiidZ6z4BXzs
Ke3fczsmyBIZlLrP+L7wmnhozZu5QXaxqi9TmWWkWKs8hIKPT53nM8/skg3B
mQiBSJYOSRYZcoyajX9wTtmu8k5LHMsI+/M1lFFMIZXAlF34afF4CnXztDq1
+k5CFzYq1wGaoIMd6GwnJCmjRUYqCihUqasQZ8XrreDHLFwyUKOQhJrWERNf
bNs7d3crk1hLY9q4/qmLYli+ZqBGbJyF63s8/xnXM8yR04wZnfayxKyrrZlg
MsrHGU00co99G3ObUshMMMMGD1a8nWbrI9weW6urzp3DhZYsg3Zv7gVgwq5I
7LJPFsJYsOuuMSKnCoRYbE/ZlL35LMkD6i2h9FCS9PBwuzjuCovRaMT1pQjf
klOK3mbMPL+Lus1ClCAZ4ZAKn+oy6yYEL6qLz3WDuHM+oQOvXwh0nBwcpvL8
pX3MXWQMum595TxzTuPHS2BZTrtjdAfiZVdMa7ebJ9tBhbP3Rg9AdE4UbsAW
b81WparGRM5moCGqsYH3wJo+8wlPyPmfkSdkWTuT/Bb0FbBeQEDV+y3Nvxv4
ruo7alkWMaOe/XZFQCNQ+Wd16GjkomPE3lsovl8horBDbcTAYeIAXfFgqehV
pqu8ibR/PE5iTgs2xiMZnuzlAG4whpxgBL7zI2d1NllMvjoaYZFdgQUYScWn
jOlG0wpFyjskPPJrsVn/BQ7+hX9sQtb5WiwtMG13l3xcC1BtJG1AfUVAn9h7
l/3hthCwUgRcEWOHt4K3VLUxIivGPxn4FBVPI0j+SxaTnCq7n1GtoMpUt11x
tAdOjsTCYLEj2Ex1hUAesnVw/KfTGfupWfnZvEMEYoH6ZHCEjQ/nYEHbxwGz
hrp0KIcVAbPIrAnrdP3SOtHDkaDCsXB1toM7kwO2EjsgaEx48W6fo5+UxR+2
WGSg6fQ+M6z9ugZnTJi53LRdNtJTODLJdDkBUSKaXOBGqFwukH3E9Bs659NP
ZylJzOFhqWc1UBwt0Gp7ofgljxvC5NYS0OPp6Q90Z0vTl0qWfRPr2Yv+V+Nj
iDhO2UU1YvG2H1yBT1toyYpgiBUMqEKO4HAjSZWfzCvBZzes8GMS4tTepSvC
ms2S1J1xIP+MGj4dvbLQnBgI6gTd293J+38x2vtNLk3BGrVnCTDg/ekydTEm
tn2CR0lqG4MHL6tomkGiCRL/3a7qLoU9F8WEJG5bhe3njrP7iib9tUoQke9r
PQHugBpYZ57MgaE51QOeMsSxP9aJxTvVbFyL7ujH151OgA4apEDSOUq3rxb8
KTOxcwuodF9de870tCzZ58ghGfATtAWSI8HVssM+j+xEILFFD/PrLBc/ftQ3
zHx8PAkvctGW1UIiAY29hU87xoSl3+6YkxA1fdNxxZxOXFb2/63qG3S9QhG6
9z/ZPYVQ5srj2/Yx8EhEnPosNXUh7gSUsO7AXRn9ylf+umTLzGUR7JR4597n
thWG0mFOiE5ZiguFOHSCNXpumWSewTb0BzrSnHeXQx2IV7sjk2a4otoZ+qj0
PIwXKr6EwiFXJKV1XnUDjp9C7Np+4HOjs8MH9WAXMALOwLM3R+DF85R76ZRv
lO0sGChROX8oa05nz5ryajnrBHEdPEqRCw6Pxli88rEirE0h9bwyC3RfMgCq
x6YiTUhmxkUVxKq1d75HehFiy1ZmtobybRmM+3EHdqvUZTJpzgLz+1XV9imp
dlrbDYpR7XPY07/vVwBbNRCWlWCy8p/daJ/ebs25X1QfYMUd+AY2ZJUx4KBn
MN5bHbS8rg7YmfTDsjtiYexXKN21FcmaBDqRFWhxsqKTGF0YjWDnwU0kDLC+
TuPaRNfcHMilvY4r9WwgwZIVPTm4sda7R/T6A0ylaufTFe0dRQ8pu8VNJHdA
kXd09hy07hZcQAMD/5NLhQpyoVA7YRrDOMVIKS2AsqmReBE8X0/8SFzDbkRt
t38tgu7/kcodtTKeq47TAXvcg/HVO5Y4f/cdL3lm03yUOI5P5BAzxS1ldTOW
GrcTAn6ozxsuQSMt13SYe99WwFMbpmmu2WIxTlA10MTGON0Dt5ctWOwutvzB
3qLvrKh4l2t+RSy/4Rw5eVVJ69W2aRce7p46ILBlpAVZyyLc55Q1X7ayc13l
V3G+5gGcLJz79zTWOYHJzmevbCjTFmeEIxG+gcAl0o+eE1xSGMAhbG4tyf6P
uuUXhNY6eGQhWLAz/iUlX88CfRoO3hqdq6C13huccd1B3q57MJfjbuAHqB8z
gqfRc6kv0dq2wolbo2FsoNTVcMjaAUtuLgjvdElKKm9GoG1eujkZR6CI2PK2
36h8uua7qcWwbeyk5mePLnn3e2kHBq3QHdhU9XWDbcrLXsq5ukn8wYhOvZv7
DByP8A/W2b/V2BIl1nv11Y9VdKKEZ48D1x+LqGDiZS/R5TrGpYHV4iY9RCJr
LcpK5jA+SKubUa2fOva3bJeUwr9+ej+Q9RbNxGUY69iPSqFd9K1p+4VAt3oq
LTDu8Bm32EsyzmvnLldospUgLG8s5fP6PhB9aX88bl0lZx2sYkEQs7GzxTyU
1zk+kLJCCx+PUX8roAqH32kKZS8RewHNiaLkfqidlAgvDbxLy1iqk9HS3CtX
9wRUkrwvaFPAKhLlfA0zNEn/UQjeJGEEDge/15hwjuiUmdIEkTFNBmDGV74A
Z0y0GQn4GgbtRCWqAiUHl2NH951u/T3Ik4tN2S1l9WFrq40AgoB8hzr/ketD
qt6wKTOf7r5H9IsNM9o7VEFMxhhaAfE97t5mm92Iryw4bJs6Mw3Din6lf9+t
zzghVJKJNeyCN6NQyDqlyqk0AkfwzXNcIwYScykplSd1wMTVe8Al2iEZ9n6S
K9aODBsy/LJQjHfr3gNPZuyugl5xPdsAIvMx0OJT7dz2ZKdoLKBBH2DajtlM
UvKB3S3GH2xkN3ZFdiIOF6lV8oblIgzUSaCT4w+b1+fB5IuFx2M7PXywm58c
RS165I7sXhdWoppVfkdFVQ0FNq7szRTtmad505lQTR/2HWJUNm3Z8PDMu1GF
gQxpKsN28XSuYqsZMUbx0lK7LGk6LWXD0lIxMH9zCWOv1S7efBCFYjEDcObU
NWarNKxPk4+qIFEcf/GIB1YqnxvJb81sP0lpOWRT+aTUVRU3IOHtgK4i5lfZ
v+ZJVNH6F0vPIgQDJcivfnr4PiD2E+npV+/qShM6AjkLZzCcShqmGKC+fGHg
uCou+MmRftCw+5bkuVb/rq9FbldNRfTq3kEHY/FAnjxu+QM3ykCZg+XsPN4G
D2OMskJcJoVS7gPS8HugGbmP5q92A4T9gx4dzqWcGLXHxqztgF1HO8hLPOHx
C8focdyF1JUNlPty4cqiojwKjEVF+iEk55ejDMC2X2c/lpPoXK0aaAy28Fzn
hQFm4yzH1xtQGo2IxfZg/CQIiQcz0KoQ+lk+878pKWs+oz8+ZVZoAJOPjE91
Q4dWbGfU4vzLr1veKx8JcB+QaR0G3LSeyVPQJwFrj4YVnlDA8aVWqqvCc/e8
SJ1kTAgn+qlq0318NjMdHs3ikBaNYWZX+LINeRdVnXH6LNbfYscA8fPxH4nZ
B6DGump7scXZn8poDWD1cZrix9DvIPzf/agTZs1A0TAZ9izmTIVr3k15M0k+
c8aSYy3TkbH2Hr/fwD9rXpbEykymK5Q1jwvdVdXpQnrhnXFYGpRWoBvfHLxj
oJ9aRelaXXKbNcDLMWvXjPrCY+Ljr4F46lLML7khbwyxOxt+WlTSgx326pGe
ZA7fNO+F6X8ki5S8cf7lzrxyYVXFjjm7aUf16elFm0nFlfc6/Wjl8++hMxRi
8Oj5lCg8SpEK3FL5QHKD76UmFOdWl+DXVnzTwV8Nz+OfqGGqNHWRfxs2oF4B
CYAGHhC+t9f6sS3guqDI40RjtmTnRQC7Oo2frABGoobb2ds1UbZDCuJyiwFx
tvTBm5QXFxCF91AeNcHoWjLkYLwHdXDK5odiAvUhJ7quO9brmTOFU1ifuJud
H+vVhesQ7auoQ/GxNhHQXTTS8rF715jPPjuyeqPwTK7uWdj7DvlnA3W+DJcs
i6WbGdKcGtdVYIOyJ5DE9vMWnnBudM1h+vjgARBTXquh1V9fe9Y8tL7xB17F
9XxpIXOKJnNe31Dfg+ixnSm92GAFSPxIHVTrvRreMOscMXEu99FDXSD5iDU3
+9YM9vc2bJ5tU0bJAJ60gPEeyzeBIMbaJhVDRPy+lABdiYBGhRz/N53cAVZt
GoQFuNyxYTpu+saaMibLxNDvJKMFgMw/VasTtVAUECDUznTku9+r8k7TxI9P
83y4nvHzKHb5bxWAH60wvHzwmDRNFmdj+A89yOUfijGaU/2Z2e1ooVAno+ct
uQS+T/SvCp1hEk9LJZE5ILR60z+u6+u+t8fSTNReywBXecFUMo/4MViNEiex
a45zRjWgRZj0k1xGPkllbCZP4jbSZ9ZrsBAWXYBGjWJYwK9xviNPFfxF/Uog
FLeaE+Ux6R7yJtct5twPenLXVMkS3dUzDmsZOW5bkgVmchACGvYyRJJmBTSy
KUH5VCaffmjBsxlteyATgYrVwB9kxVmk2AMx5q/pELKFA4hJN++gMxAwldfm
WSlJUfXm3zkLbhEUjBCasaoRnR8aXv2DlCl17uhtYyzH3tnmQ1HOX9RxdzYz
pJx3wQdGWuTUXTj8wEvDNkyJoBQCGo1p4qjBFPIWyRl5IV5GnSXdf/tPNONd
1ZLtQO6g5es1O2g6IWEeU48O09cR+UIkmLrrODmKOPuCJkk7hoDLAOwRqSyC
ckB96gcgZG7RX0COviFtWqDnodRRy8np27ritngPTEY5h5lC6svvlnWvEJA2
TQbAm1PEOnZMB3KJgaE7OQpKQ7/uTjtANSoHVJALWtdJe5uvZkasVPkFbYNp
o1DQC+R2zUVudkV5xVpcf85C3ab6O1ZUn3PVuuv5zWfOKLR1WRfbfi3Kl8nf
7LMRhfN6AcY30Z6coC7yN4WxU7RAWGze2i2JibM7Vqt+sWO1oeBG3i4rz5oB
GAF6v688Mvxso2JfhD4WSqKeO3Zo8n0VwAFIk7oJx+Gjz461wPasOhd38uwg
D2JsHfTPhxUZzNT3w1zHhMoZOt8RLSKihMIrFWm5RFnmNydvd5FSCKs5ui0V
ihIPSxO6GLrYFDPsTCppLrSA6Uv5dYAXTVJkAdTpU7edLx0mT67mpgQ1nA8m
ZTCGulLQn7letZGibjFfFd9hiOiNEw53yjcLzPLjDhjWDFoFaWN94Jxm9lu5
Gy9jYZgOHkUFIlNqFduQYUq9snC5LLHHcQdAhDzvqLaF5hA9bKZkxmt6sBwF
AOrinPKHWOwg4hiMhEgH7Wq0Xp68DttBg4FlnE/cuaPjXWnmKyiLE13JNbcU
jkcR2bjvvhUlnL3i6oVR0eoQE0JNBEDKXK53Ve9w9d8JEFL9Pef2yUL4OlCQ
FszccaJPKxPSiDfXowy4G1NKRR7Ipi78t8jkre6uRm17OUVF9lZ4LUl0QQ41
5ChYuDVrb70d7kx2nqht+uKmfr9LMzsA6W/BeugkRUQGHUwbuXxwTojeS8yL
oHsmweApdooLM5fpPLI0W6dI3UogTtUmP4mbZ2V67eXAOWqmSDiHIgbKS/tf
kr81R2bwJ7m6XAgmVc3XZfPFxh+hBn2xBY6Wsdcy6rTLvZ8aEHtLqP3gZk/2
qnhuyDjoba7PAmBjnJLfIlDfyeurFN8+FRyU0rZ3vPYx+60oy+ijpf61jH0/
mNizv5ws+IdyYvJcnM4lrmqxxze9QclXYFvuR9KxJyJNQ7xcJcTln9sjxzvj
10MhQcE8KNYCF0sqq/vd3Vzu+jz4bcdMwxpZ/yXf5XNimVJCtzdq2PaNI7fy
ZNSp3J2eg1Cd5Cqp5FnGbLMx+zNWNW/fMC6P8cHXfYcuH6qu84h2RVi6EK8m
3ebs3dwu0vhQaYvkXUEy1z+vmS9mADYownvrddVtfeFu2joUPPyryQW0Ph9D
xeIxUPaQXTaowyFYNM47Ci61ZrNLvS8/7qvg5kdhLDY0Ri4VwKcgBiHWUyqP
NYpbPfzUAarTlWGFIC46bj4Nn7D9xx/wbRTTKhpjb5yI6ixVnvqCbW/0k+C4
0AOvSDgL5eSCR/Sjh8tDKZpWPSV0zs9IBy/R7VGuDnybYHbWIFz7/lGEo91+
lEdzCglz2p4jOSqz6Rs1rnJINAFkrZA3DZ61bjYP2bsmAaPMTFUcpb3YS/PO
Wb1paHMiR3sop3MMGstNdqQAkwfv/Qlp7LctRV84riwBAvibpP/W28GYnMqg
aCCtRVlE9ggD9ChgN8dJ8co2iqUvguzMZpsm0ydB8ZYTW2xO1ZbeYcz8KdQ1
nHbE0qsN8WvsainPjfDZkW8VW+ULU3E72uhDvUrtFo/vsf1oZXT2lXpaHtAZ
zboB4S5spUv0gCnJ+ILrEyCwZoPTIqW1cizgcHDnEWIY+EiVCDdoiYzJP6MA
WIiEtBEfwCI7TGx+B4UP3WiLGHaUr9AA0wvXGeOYYetbCTIJk2CsY090RvQP
yEWLg7MyA7gtL58nMlh7txbGhVIWccgpgClf0r03/meLd+RWDMQaY8RKcIND
h0yknbp70D2BzFHmrNqa1BRIFIgNCPzCK/dhsF53faekiwJ4UPYfdzPNh+pf
cPtXP0lDDQ+9rwXnmHmSRJOumG7o6ZJcY4I2JbWQ/VzsxL8sHbyPMTZVTlDp
s9jOK5BRqjk0g/pU7XV0UOSqrWEHVINGDM4Pu7Rs6ZLKxI37UQUxA7qBM036
Lc4D4ZntTJafoibGu9GgPORiH6ZxiYzYyG+3XLQChYFDoxBzuFvgXIwt6v6p
Wx9Gt9FNS0kUX/r5OK5RHHwLAb2IzzsnhGwiXAqqKvUbjSkS3JW5PGHDxVFL
/a/fj6BEsHYYMmAVd47TucQ1dwlGnPJJ6aWtyxIAmReXYwkXzwhrOW490THJ
3VR7Q6d2kvdSzf/r8hJSidCworp6BBndmlJKY5ZtUDXvwUmSto67hNugpB0Z
Tj1D6STExDOnpvOBfUlFzlLKRO8iiJ67aBvtYZfs80pM2ocZ6COwnRj0/dpB
I4zERbMdswmxrV1QnlVHI5P0PyJPuXhOipGa0jbrJ/tCc7LaEuFAs9yZl6mo
D+AeHhfIir5uJ118K8I1L0ijC6cMGfwgGdo1NL22kKjdfP5v9MVbyX0xAB+K
iITo4RGHrXW7A1nKhoAZCkzwkzzyR9u6FyYVBpcsdbEr+DClQ6gmXdyYDowO
QkJAu7Aod8LGXpRc7vfdhesj1IqC6o2iXSb75SCI8XMrrIitCifMyqvOQSpL
IAiEUXwDJRbZGE49mdzkHAd4sJxf17t3VfIqh7OPOhEIUTqZSrOsiu/KmluA
4m6GJMfFAe6rpCRM4ZQkOZ5dwAmebMh4aaQNtAb+r0i4gFvjCcc4dFhxsnDs
R7lASQ8EDVwQiusPYeu8VN+1sm9tdrH2OlGqZZ6D7KEw2TsLhyqCV2hFRu0b
VjOAgyHTHuklcXYdiRRseYZN4IRuJorE52ELgN1hAs4r28QvtUOc1Zo7S4It
IQkVHXFksfrUbN5VefuPSreTIFjOYXGP2koQHoJ/3CuAZVFi0527RZr9RQ6Z
32R0d3B6QVH5rU18EWtCYXXUL98LJyqC7ndaYgTRWBChEnl6VquJ5XgtFKjO
npa7lPmL8Oxf5Ra040uLApU24ozsRdH1flXQoNIjvv+Z2IwXtlbunRo7Cz1o
Eq+kGNHaCqqBjgaFV4C37Gf2yDKEmDYJOsDtxnGg40UKj2l3zzHWIRbX/4IM
svMZooZ34Dt3beBJC+BMSVtyuxIv8Sd/PjFJzvWcfsAB8/foAoP6rjJKGxmm
UCf7Jy/J9i6JZs5kTt5IYTOKOUinCCszHGtAvGTCxiL54T7ks8omcJ6pr31l
X8PZcAoZ3Ri0bNhyi3HMUNQ1EPU1Bp1Kwulna6hKb5xHVDHkgyylvttg3pOD
rMwc+UlsK7haoH+Y6PZYvMkWUCNMEHfbYlvqwQymZvbyG6XNBGQyILZr8qq9
ZSbm1pMSp2JqXvruJcalxo/IzhE0IB5/yTzK/gd2hIB1zki8z1xkdl5HYZuS
hqQmZ+c8Kt/1/9ncSilJ2qcWUShOTtbdEvxJ8jMEiI387Zcxdx4NlxbSxjBa
DzhxaHzGEMvt0v4Uh1g0HndVeXWiofdUOAQUui0yFncr15ajk8TURKxcc7Xs
QiSaUaU0HiNts0j5k+r5FFwKzflSIMgm1usiekrzTnUbDUrs1XpH3npJSVdz
/B6+G2DQb5OSs4ERoHkkhDCCl3793Rz8vbEdlDoIxvjP40nyUgNQJz5dDJpD
Uy0qN4NLb63MjdAohNAw0S07jNNlVg07sbaoGb7CAVyrmKaZOJ43FdaB3oaE
w9u2zrDZSaukg0WISrEJll3njrE2Wdl8SuGPONIUBZU0/tRogQCgBlu4vOUU
9RYzHUqx1ghkmFeahXw7iz2yTwkL1PzazBqtk1rQDlaZCMIkfZYyc6ySNgpn
Z+KNXgHLQ89P7LcH4Q2g27eVjXETADJPN79ZPWtRvvncCbAUx2g3ldbKjR+g
8qac9E1AwZV0LDO5+gw6+pAcQZylMllTESd/LHSdxj5+zo7TxtJMCooB8/5v
T1+/DRdbKCj07NiveAsxDlbKsOVJ5Mv+wvqQTBoaI6WIaE2cRWsCm/Wq5tOA
qfG+YNdn9fWRdpLR8Yw+U/kAME/wsaSSOuEgNY1ZSTmwsM/n/GJ+d77il+j4
wULEZgD8EgdkFF/+M40itv1N1FRt14aW6IszbLTYpGxaBgpC8sGuSVlqimUK
8mvmhNNe+FOXm7929cJbd/6q79d33mZoP1M5ihFMbutdLmDoACGsQyFWs+oA
Ax6cUm6Oye7D+fApwh93GdlDDhbRboeTtw2bkV7Y520ynrCbV4jW4f2B7cVv
aydgNn+Hvt8n/qPLwdj3GviAHfQyUYQQJm4n8SNbUp4qjdMVDoXM6JuUo5aV
6kJ2l/oTEhPbCrHEnfxh7cIxOFDGjEj3BXo9nE0Lg0qgqHevjfyfoig/Ip1l
maSMCAIw2MoUkaCVLcVuEiSTKU7zayRgXoSF26m00LyVmhDS9F4976E6QTlG
UZULhdj3sUCgPd0CbvYYjN7U3kbJgSgrAL6p/Mm1XkKzTWKS8sBz5idTQ48A
TLehOB/hZf904Q5AUMLgejEoCRQR5i1frJNNk3nKBHGRRqV6s1nWr4iSzjDR
aC9IA2o/G9NBvfPP/KFXptRxHCp1WLK44vC0CkZ7FTxMahbgaWUj+fhbvAXk
lZIG6geTaaxxu8JjVF+2jmTOUhYs62nzLPHxEdizM+wxM2qVUQLuLCRFODPv
E65xFAc5YtoVT/tBHTjhnKJAJEaS74OfKIx/kkviPD/5CVVbtaXbHuHUxBpX
kKlRrWZsrb++6uBsO40ZV7CI1ovTPHM+lH+UkLkWry1gvsjwV34qoTLT+4Ql
9Ourh0uTTybIRRa3YVxvIsgh+iOsYc7o/gMqgVWhwBhxoReyv0k5aP7N0H0e
IgbVyJewlqAEfDMfh3OFAavgS4cNUwCYhk+f+THrA7LKTKKA/je2pHXcZWeH
Mc+AtXy2uGl/2p/2Sa5RwE6VQSCcVjWbK21QDvxl7GJSCjFpHMKd6/eVCvst
bjX/Py84CYXKcYRw+K6G28V+VDudKAR57mkGXw4nF0fvdJaOPeWXt4Uqxrg+
JfuQANygyPTbLetHvq9zYRxaukkeQBpp4WD0yD0LOIB4Rgd0PDRzkPjOCSyM
ZoFzGuZNWuumWvpPqmiYAEuGve4DqcmUWxCIC8RkbkXfEa0o9ubiiJboiIat
h+Lg7FJSg+sd0Cx9qmUtyudzNzi3z/ZDuTWUoQJL+5IqCifcffMU30SaypVj
Mxp9GwDVdsvoJEDre2n/LAwMZkcCK/s7BWuJDou46AubbTX7vrUXVW0dZq+e
Y/xysafrRHIrjWr4XLfxq/FZ+Q0ffq6Kac5wbFI6KtQp8SCRpX6WqrXxm8ua
R3E3y0GKa7gD5vp5I5zjS+w4UchkCKBSVl6RSO/dOnPRb+cN2KFBLDC5YSms
61BtEVj4ZW1ovOwstexATMbDBCwy+N4V5OimmbjJvNNXHS0Yen6l1bAxXM88
rOXa4TrSrDtl8+iX4RvFXXDQRaw8WeiWU7gbflVfQ1Lds/IxLSixNsZeGbj+
5/r/wYBPeRTHlTUjpOUKTTPUH87KLxUKdTkYIJVKshGV1/MS5w7LNYbLBIlw
GEYYTc3kRfhCrCrszlXUuJUeELAGdigChOndz9ea3PQmQ1dLHj35EgKzokZ7
PN804gx9vfLNWw/pupi7bQOaKjzG5PAozjMe3wzh5rTPiaZ2bOAzReNUcsyK
+h63PCkqMKQFHCso28AYfjqjYpBToygWtuIbxHuF8ipcyholbkd4OZZoHbf0
qBMCVJrdKzT72aov5O6XLnmyAr2g+36598is2WMqo9ZNbSkzvWAJ+kg59Os0
ZAD/f1ARgkDLbnUirBCjmx3De642W/a9CJeeUVxKMpVY8prrw5ysYcp0Xtto
ZHn3egH0ms7lZjyVZdMYs7g+HB4ddX/9v483S4tF/wDEDDB+p9MfjWB70STT
alevNmVADZx7U7NYJbOfji4ZX6pfvVchnK4yYymZSj0itcizedzNCl75EdGz
GOT+DwBch/PB7sZPbkkK2/1HIKYtbDusGXKylnnIPOoMFfVMDBzfJYL5sLo3
ISexJGqcnDz67i3qB3C7dXZx0VC4FHZ1gbG69ysMzA/H1SKwXFvf3c6ZcUHZ
oO9+aDSkQD2AwGCL8bs9Yemqw1mau5izpZ5RSSyDakdzIvI5ZcGzCjZPlrA2
EKNRulCZ3rE7ic8Lm3MkZBdDN5FzIU45vczTjwmABC47Qo+mlKSFryUUZiWm
aWH8HcDW3WGWPkTEXjLSMJuWhIG2//GBCoikTmAgzcj6NGFZ5a0O+kU0+sAH
/lTOv5yuQV00Q6OW0Ozwee4xCS82AZk64zEXvDFewMkjob4qk2h89+vpcljI
NAxyaGK3sT+b51IANUELSViS7Q1IW2zWBvbRBC6cKDWVPZ62dCKav5CBqM6d
dhsEO6eHlpX0PriEH5z88iy0IxOu7n7yTeL7ngHamS4yfg5kxQgswCMDfbu4
wi/tI8tl4cp5/HfMmq8UFdW5LIADzGGkWK0OoF7l3RRhtT0D2EBJl9BZ7ACS
UNCNNfS7Jf+6eQVGIuycdx2tkl+RWV0fORqRNd7NccN5WoZpRZTi8NsjnmYD
uR0Ub02KOLccFvaXr4b62Toiu88Y8ORL2t8bgU3av8Xl+yBwTAFT+bvJ62j5
zkR+ffMhcj7LBl/IGfEwTYDV4KDbB0ZXPoA9xZ/cKxrIzjJvmLw1hFOCsjsp
N01M3jRS8LYFzjOoGa+F/XG64ZqjjkPWkmTBfbyB8tGHx+YHUK8y2Alv0Uwc
iW91dVA1P1v392X2QaUFcRdfMgsCZEUi6+wsKWI6n0KoqXMB8sSPv1b/0Evo
uYkcUntSikdt23rrSS0mkLz7YukLOU3p9HdBj+BhHZQqvD+6dKZ4Ud4l5K8H
nMEdP7KIIVPqeUArIdEEL45N6hrSDhMIO9wgyN0FVdv3X6/26jA7rUEIT5ep
a86lKV95WI8DaLoYlOlfQXhd5GmAsNL2haYuSeOiL8trRDC/idymasnF4iIV
47EBybOKQl18VJaDeRd5oUnXFzz8d/7PnJsjORonmmQWzNzRTOgbCYl3IsXl
t4umjnHsoAerDYEAG6gmwKQ+i78I4AZuZ6jNo9SZZvcfXDVyqP7tDuf++fwL
Hfd466nTpqCgPGeNOSnIB+7089QZRa2Pe13JM45g2nyMEdrrCjMRBebBNezO
wWUSGwk23K1WtdM0zls1ythhYGHi7itJyzJbgiytsnhr5cRqyk/0hL8yjujM
kFtmdQMVUq0L5bi9QZzKSQo8g06nAn2v0x3xsjjSbzlXTGBlDd1Y2az1k8fT
v7OR3Jp8XXEC2ktQHTIs28xyivO7di4cYDENAuoAgSOH8MEbMNEuebslX5GI
ptRWbT+5yKTsripoIltTkkynLsnb9nV2H3rXUPzRumLIEOPNUgNMu1jWvXcp
lpz0YGpiBiQSFlnSpYhE1L6fmsScIEwJVX72uSES0RVceaRAFMoNxee2f4qq
3VN+UjCTnYYyT3wwBc86gLbVEr6e3RV8nQmeolsKVztpHekRZzWWvZjRACNQ
T3bnD0/0i5CJp5M2Yb8UHcrRhpd3MVq6oIAXT3HSuBLK8PHl5AvMRtgOuA0U
sXNv7YoX2ubd7TK5Q18qwtvoJL8AEiTVOdA8NLqjMbZD9RDaidFMieC4HwWs
YRmpIYsoLcgnhCX31l54eFp/3XgbKTiZW0Ux5pRyh//DKERCJQO+lJ2rGL+F
m81sNxZbpOjtoPEps2ounv1F7qSYbE4Voe0HhMylGN71ElTMt1oohQ4Xa6c3
8iEFlyKa4/0xn59mFvaEdCnzCsihL/Mij36mjeZpgGmUuo7Rsn1T8ZdJ2a61
r3uI3CcInwGPzeUxo0O59T1K20F5WrEanQeAm6eKivsvG1qYH51YdaNdKVky
UL+mRIrcY+eHz5Nr3ZlsLy3Y3dLehx3qbrUQ8ff1Gq/kOt6EgJGR4tn3+k7r
LnDsMaXtMwzcHYqiV4KSK4QYUjmZC2ya6i8DFAHQaALMoGXcA7rlsM9QRyFy
W700y1AIzR6wPC+O+vP+/CFSVlQdjEMhkr6DdT5UF4863tqNTjZtwiB0sA+y
M5D1t8wuLdIwuU+VGnyq8SCzQB+7hKoMjbUsHTn8113ND8y3NREVftoRfB5R
k1IjkB4Xvu+8TBVzEMDp0Uusuoz70DCUJMdM+WZ7nN1Z6Y2EopNhFQB1JCSf
SOJUBQdPn3yiSb4DaxUMp7IkxO6mOj41cs9tsZ/bCIcrjvwriZZGacT2L85F
cxHwVOPmq+k2bTRZMFpZtHquoZp5A5TmH96xPYNCBOtUHBhPgpfekb1YrOnJ
ETZted3ElFdsj1f7XHGeq/d4o6DOyMEdIGqWFj3EXZuFx8GoHCzz2RJkowPG
8vPWR3qERoGzKpgwciTrALJlKI2EPSWe/84L4cYuT72SO1tJhamaQ4SFm2y6
1fKqMKu+NGvM1f7QESk7CljddqzNs3a+UyHKprDtAatchDkf/0GaqbqV6UJV
lxcCseUDPK1s5Dfu7WXEHI9gccwM/PIuQixXaIW5xIwQhnJWOzcRRrgMDL+w
bZhdXC1JcMtOgRQAgiyEWMfjTsC/UfkcglMn6xpwtCy4vP+Tht5DlfubBHwt
PwpDhzhjrc5kywh+OyQevLhw7MsStCnGLacP5IPRzi0TDzh1Z6U7K4Y9OpAH
VSE0cU3et3nUeSCpNRUxetzvhfvCN07u4BAOgXRK5vfaODshY+6AlKwHQH/f
uVl+fNqOtocdGqy3rqkP3atK5lGQSXdUxEAILulOA2qV0KozRVvkmTmcri9T
NFrFQHtzqLIrhlMDW7tNzw+Gqu7Gq+ULKyaa02we+xCz1Ab0pnRlAZ0G8+TW
jf9aJ6e+hoDSryEKPf0ze9ilVklmHSoTZ0xAypCrK0gQZDpI/U0IWS1UGijI
WYd6dkGZ5e/6hnNQhNLRZKNW5Wo6rmA6qGYeYzbOUg6gDbdNaBbnlmJvK8CG
R7DzCDDvg7xDEuJFhR7nchPH27eKfZgJ7s2oI+T083GPh8IBXWEkZRYlmRK6
cQtujMhRDf5AzQYQPOZajZDA0C0q3pO2UJJcnPP/7Zglfe5Tw0U/raSO58pb
MqarCKvNIcwLa+V4FgUnQW2tbaxLaiQ3fwV401qKTIofl5p4NH+Io9fYbR55
tFEHh4DqwUizN4eYeSfiwjFuAMXEDiSz1DX79hCVqiqtbmbAF56kgXKWedje
jlNJSaGmGMagxc2UE4fdZRzt7oHDZxD3qnHl42tPVxFw2SYLhVUUlXNlYgI9
SelN8DGbOZJ3ql/MhjA0PjHkIdWwVuz9zmGrpQ4UMgSlylVYLTS1S1Jnhe85
L07CQihpXhzzOfKseHRtgiEWk9hLQCAf5EhXfF6lPMCS61FdP9StZy61Bom/
7kJWHencoQzUkl3+Y5MAJYng2kRSJ+HVJRXtOMD4qCxDqvyMIqqeoGHtPLhg
tRkE6hOuQtkvgKcCPPvMPYUw4Zgo5HC3yQ9orN8aXdD/0P7qqTl8Q7A3tEAG
tmALOKzyZeTuDga8pZe/h0Mog47rqkRFEp7L6ci+gDa8fuA9XpGzoHIaLb8j
sQCxN1mR6jmdaY7O9CAlh8RzwDxB7bwhLsfYlevQAkuABV7a3FQZMV30/i7M
eHGjPgIATboQlct2pBzMFfjgnE0fupw8MJa6j3s0spVC4CeglAOOsZXyRVN7
mGgBDXwaAM3tzJ9usBYNnY3Lhx4XD1//k/vRyFeaPvbjvADYbz2VsNwI60aG
kdr52f1UXCHeNia4NB+gdy+nhVP74fyPJ7p/q/jwjyl0Z2B7+5OCBkfnB+w6
vAfd2GMEDm+s+aBfBKU4W8fOIX9v8ZhoTxWSjcHkNByryOo3/oyvfiPVe/DV
J5K0cZ0le1ocOlbHCmXfxdjv5iYcLEn2nLYzg984wlIGBanshu7PQvZXdiIF
PPIbGelD+jYWtol83Kh0pxSlO1XWhjdB63ZFFlPDF8OgrTUhME2bB+6PjSsO
p+gpyYO/At+SMCgJDwSFFCkg/zIjF2hidckeIjpabvZySmmzu5lnRKY9ByJh
qEfd0qxknxgQe2nqpnVl9htaxEwDgYs+l6NHcQ8fU9HnrYiH1pgCqyvIOppc
c2iRJgkkdOk0djqGuZAmldu77Re+yVjZEva6CR+tFbl1DTzKcHlkX3tTIg4m
5nTaUlUEW6KS5m5Ywit4N+UnTlD6IhpMTOsv3oHLigiMGEFfvEWMlcq5pXLv
NeA1PWhHyJE1Ilk2yDk2knR+ggCQ+vL4hL3O/RQEslAWKbiU22NleKfo6Zmn
PKUlhpVU5hS2AoS2FgGwPH3t7rcJouq8t7hkLVIS1jLi5Jh3IRR2V91J+Q87
7zRJw+GafvFTg73bgdUxwfxS1yq867E1EM0oSa7CDDPG1ngwCj6AO9CcszA/
gAbNrQ1Cg2fRAfiLHrjPNkR7jxZiHdmNw9CKHwbqxBTEGf24U7k0FnTRsiGI
K/WLIIRpQU7nKUixLn7hZZ1i7zGqkfNIhe9u4Z2EdITjvObBrJKilsRELUNH
L7ID7x1mLxH5G48a/Vahs4dXg/Bze7YwCaknrsmTY+6XMCszRCCktsyQJicl
CGJr4DCWLg6pgHZIicoCxVyx6clMaMG88uHem6EWwAnNWKMl3mZhGjXuFOIW
cW3iZDbqtboWnftRbmOP01yMpi0VAaSxgd01gC3HxQhLOPotQlUOiEo0qf2O
Woc7L+8PUoIup4ZmjRSa5oopdTa3RkX0WavLSbn7fbO9Cu6LhNebudTEGQxw
El9fz7XCpo9uowUNQ6lCn/11NQ6du5by3w0/bG4YkESl2mo+s6NiOyrVH5UV
OXY03WeqxY2bib/GeT7SjdEMzv5ND40ciYscosSyDsJhHAGNP+mhN1Y0/VdG
W2YK6cYimymhVUo3GcEEocmAYa/9zFrmpjn3IdnWBoYdl2ispFebgHNLDv6f
LjbxwY7N09jjhF+Hn66cSf+Vd0MCTYBwAbcuY71g1yzaNXHJckPzLUrqEIZa
i3XXA/jLx67aY25/DFP4jGT9l82llVkhtb2/GTHJJyvLLyu0seT5XEvLFyRW
/2MYnGxYeKE3z2QEJ/0qQalYrLycN2iGxl6342M8C6BB1iwieWYuZgtdgzjK
or0JTCr1wR4GGokqoefc/UgnRswrAK7HRaMNG7R18zkStfQpzioKX4lG8b5E
WvDvElJCkN4ksfvvt5vpkmjNtARSa1+Ss31Hw5PlPaS1zVVFR1jS7GMiTeQE
mei9WYBmsnIs/z802VjIRVXYdVBBMG2DMdiK3S8TImOrMZnJ92+vlxeOYZLH
AcMzSjCUWJHz5mQv95hpVUQaHEf+OARqi7AkbbFl1TVOJPbKKbPaZ2FmE8WG
nzR8Ud/EvCIasmBBJf2c4jE6CAlBjKCkZ3mPniceH9ltlTgCxFZcfReH38XG
wXfSUehQSJVWthCqQ7CL62R5D0bc6pWjVtybT+lgtUmrCM68IqM7mK3+Tocc
UpDVI9/mFPBUYVVoc1v6na3Pil/5j5DJUga9HSroohlcmzGK4PB8fKtpVr+k
EUZTanEsm0MC6XN1GrFscap87yJDgKJU9RIPpqQ4Ri69OlJyE/Rrc+DoT50N
480Xt1PZ3g6f8cTl2eF+hgk14whVyFwFubjL/9FjmRdVudOE/moHxe1MaWs7
m46g4eJrRjpEnFAmcYZwkht/1R0XPci2fTV6kMJ88behnOVBFjMelP1SKBCQ
/9pB6P/VAl33turUYiPo+IebZYYcHi/hvgc/+L0z/ovn+LJRP+S8ldxF5DEG
ASnQm2MxzRhrXbO9RL0yFoXPOPOtW+qYWBV+IDM6uEIEztToP9kttWS+MlUY
kqm7jYZjF3H8I0/B10jufzL2PKFYhdxY8OOJjnakNkUkyDwRck4iKTaKhBbd
fn043KYvimVEMuc8dwbMZF4DvsZvsKf39rSLBtNnYp5tAMXC23zwDvD9yuuc
h2Eo5dAdJvuGFC5c5TUwKHlvAfDxpHmsUx+OAzDI80Ef9y0z/cqPeUGSxoEb
CEoj2DE9hTluMYvPba0F+XLGF7tz41m1tL5NXQ9hxX/EtiExCokvBG7wNRYe
SSml7qA1gSNXnjof8sG/jlBWgrdju79xPHxaGTjRk3Cbi0uMJp6/rBq/EzoZ
S6YBk5JMVb6irB9WJXtOdbfNC08/9nY4mzxkmDQv1TlHpg1uTlp73jsVg1qA
VmRIdVGjHo6w1ipQTc+RVIDt2MPIhEl1WgAKiEJ3LkRpjrfnP9YmyHIiH2oK
vjPaZD/It31VxidlJWHFQzxvPaxIp/lu9i1ge8gySNuJl9G5HsOVLonAGBoR
84z62Z4bREIip63LNTi39VtR4h8JUM5PAsv4FUP+b/e2raQim0FF3fiB4Tld
tOHZPT04/gYDQuLdhtcyVhF1U7N22xUIVEb9WxEvMMoEyckfLEFqbJ4OOOiR
DTmTvP+RcU5dQONhf5oFclR+Gf8wjcNqdYAhMPWA0p4eV4+btQTc2nLql93e
CktjH7UFuEZ2BiiQ1EnvJFawZw1oI+hnqeE0qr3fjF7KW9ydtAxxH6h3I6mx
QZbwNjWeJ6/TFD3YcYLKda29JyheB/xQ/RsWw93JkoYZ+wljnuLN1Sbxwpxw
mekkisVqf94D2kv6W6K/D+gGKgJPVz7qg0p2/JmMbenOdiU8w1HuIPjoP56O
Oglb6h4839dUSbUZ0uqQPzQPrS7SxT0IZAQrdRsgu2W8GK8gTe/SVaBAtsTr
K+58ibIlnxBAey9mhff1oI4DdZEhxQ7XuprVul/n+e08LAmFmTTt6kRSzfvF
r9wn8xib5Vqw/yHewgRrUDXbzZC501GC/WKv1HYo5890qIf7ORFUhuNvws1L
HErHCM5cN5RFPlu/D1l034fo0pPYhh/uy3ftw7HYXnywAPLKX1zGLtJj4N1M
qpiUUgkfqVhqXa8HDuiqhvucmXy2Q5rRcEA1kYQHD3GxMsw7GlKeSOCjQ7FC
EK8GHeZUhFywzAQz0Dj8rrgsdBv4foSE0ELLlUkTh4tmJYz3soZk7MnlH3A2
NRmsZUiF9bNQNN1veKq7B7EYq08Xf6PwNkmzV+i70KsDg4UCT3R9LKc1Jizs
ZCxMzQytpPKzvTrDIvyRk+xvda7saUmgXYTNvlMBb14UPkliTf1FWotKqzXG
tjT609jNsD9RRTnFFBxksSWr2sOlnVVftLvhNxzYYbeDLUJDRM/YWqEc65eD
5w2OGanu6UdK3JINCIBy/5GY5YZuy69UwXgZdoBWRxMP7v2E+2rwgXNfaBvZ
6OPOssYXRCJWnysPWa4Mxw6+F20GFR2TsGbQGwbTRD6EYjBUDZr46bJmwtAT
tbRvLhIWGPB9o/Y/1BzxdBF7Y0ajLpfzX5Mu4syHVd8wJRLNp7E2eZG8Ihlw
K+koYqMMO18T/bHHX6clYTYgHIIDxjKo083Vf4ebg6Hxuyf39s03lb9EWPt0
R5es1QJGFgGfXcTk1s6Pf/CDhFLnL0Kbi2G4inhGteDzyxnIM829I2P+nnUw
fGd6mDZycdUrQ1Pa7ZnNLwAfkKDrQwGtYTjO+cIiwv/FoI+Kylr6rBXZ1wQ+
ke/CBe3+VTsdZQHeCJJpVcXzCGcKKNYJLGlJhKvSjWGLKmDXQUoZ1olpNnjq
XNo4/YIe/Z4/xqiq1jH4sKgs3Wfe3bH25pH785VQXjeOrxt1SM1SgzRBX/8c
cldESrPlD92CVJMazZZE0U7yGKNqh4c1gX6iWQ4pB8uuX7CNIf2QHDxcilt5
YNNRK6u/jlIqE+fAuCfN/2ho4o1UOVrrL48X3lmUDi8oYYtmAh7qjLhOsH7b
I89+vBpx7B5i5Wns7ECNkIPaqo5SkDxMa4S94S8dpXaqBeZAfFoPgZtRL4lG
0I//gu127LKwQi3XNGYeEbXPw+1PYLsP4Et192bPp1oOp1PP5liNMfYuytHM
6mARxBHKRCV9jXZfVz2JDo/QrDeONWnTpK0Si1A849yf1v++9RSzxxSrfXfd
CIa5IYsEYgwZMFAeqfNZrbmgkZ5vHGtAde8OjwYpJg02YIsM+v9xlhckXjHW
xGdfdU8890aPwng5/T5KXuGV4ST4Nqc+Nxrfl6I36HqGnNCT9u1e9KXqUJDS
+gNwRxXNhnLtrT5aXFsFXkhMI8Gz3d3jgRwLTTQJ+SbKWrQlTm4ZT4yBybjx
Zr7aLJ5X0WgLqzwGJuOn4iLVaLkneDXE7YF5Crl4/SOVY5TeSp3db02206zy
51PJzISc9mU8roGJ9rigKXiK76oDGgAJO3wu1y3LI96eHfSHnzTY8f4C0e1O
i2t8psxH5bdnZ68xsjULJ3ep6LpZaBnrHtP5TF+JaqwBEgcwtapCwwog5SPJ
3bDl4SINOhrsQqQROHruUv3909u3sUIf22LKEJymD/LLZvHAffVr6N5tU4oa
OLklyHhAeXY/Yn0I32WLSJxPKmVQALeKfDzpWOQbDekQjwJ3AIQcwpeUs7ql
9k9gfQzrvM7xWjQ71S7Zpsa0wjCO2SeTb9tinnDR2vIdLm8Gdk5gkCpVJS2v
elgZxgofEukQu7i42n5hIsYC6+ot0ybI4k0Od3oXJJ1/oAXc2CJxVaC6BaEl
kYP3XXDiVInruMxzVsX/8fHjVsyCJd9n7qHiGtW+GvzDYuZSZAbTPWU4MOgB
ecG8qcXy/ICg0v9qCUex1GPNS5NRrrYPVIinAfiIkCb0EMxBCpTd8HOnb0Xk
sxeVDioeNAaPssBmBM0ln0DJ1CEgF6s+7kmAgbYirF/E0G1Aputbv7zXoU7w
pWnY4oxyrIw8EUiyTuLbflnQZ1VCE9LkJrsuJ0tP7Mem+0EkOt8T1wGyfiRa
DWC0kHglH7LW4+qBa2Jg7jmrXcvLU1CKcC60/6RJx2ynMzeELBCqI1yL96UY
g19bqTDoNhGbfVOE3rprjhrXAEpHEp3T2Hx5beckGRh5fZetlyElgBs6kf4m
1PFhj1fU23lFgTJnqaQjIJu2fsz0C5l3o/JrCASjmFzJ/8eXjBTAjB+vcq5g
DhheAT+2QlDnKDIVoJd982RHlYUCgTor7TKz6QV3QidyhO0PWBnXUE39ntgz
322fD83KC8ewZ39ZqMt+ssJ8N2iqEiy/vcCyJrLy0I1f3/pOQF4DlbiuT7e/
IpSwtersKkpNuZq2Sq6oGOIYSs0GgqlBtiTpMoerY5Na/jBQR3MiE7oULpD8
Gi3sIzxIUj3Cuzi9YbpWcWB61vyLbf5NOKi5Kzl732BkNbuV0M5wq1VSl6tW
tbxEd7MLTSda9KPKF5uMsGJvhNTvlUfGkrnS0e//5lZ3Jvq8ayoFu9Qlrfkg
Fg0rUdcyu/FU9iNeKcPJJoHcDB93F1+wvfCuhdwZcdjfrwf8LnAU6v+mtHNF
W0Gr7FBVhmqEOa5imsqAuc+pNssedPD9rAlFtG4h7t7p6T8uaXf4SIEHN8E9
Khr6dX8eP/nLepkdBHbeXTNKGRyifGbsMl+jA07em76xP52Z/+SLt1e7DIP5
gmCGUtqQpMIfBfnK4LsfMqXnR+8BCE5GP75TGy9HqhClS1+JN1EKumAQgl6I
wd2a7YuoODycCKtEDII/vb62TphxThiSG5O5UoDeVjdrA/PtXsRlbHdCTHLP
LvS1hFomguZCjPIhelh3x2s6OFAd+RCw4z+u5Zfky1RTVNMINkXELA8M8EcH
EmEh/sM+5v04TwjMTPd+tQar6+Z+v1pD4KZPf3IC8Y857MC3J2H/TZCot5Oy
dSzZTaQvHu0TQRuweFjN8OOQ2hM4BzbB7fk3YU6TJ8jDeFPZg318vybDIkCc
6IMeFv4UDeDylckKrpMq6UBeZ5W3YxIic5nJIk72D9hCnh7ADQWdOxaXipG7
uFoErBycij7H1pH7sbwiuYVMDK6xA3dbcRru29yhCIVIynEWiMIzVGx0SO1C
D5rpER9fok1/FHx9XWqFFhy5bplpADPfLTfWofdgNf/QGEL3Z6ev6nfe/Xzu
4/NyCGWnUZTl9l+j6HwjJqiAmk/7PqsIHW1+u/uKACBaEJD1co1LmFAt5Kj7
heloizZHvOGZtXm+tPj5Y1JBGUb37/HpsYgRlh2rbXrL9YPF8gpHCt6Dmie9
3T9LkwCu2pp8mHAPQdbMeYv2DzM5PPi8CdC8SSJvXKkOJmJpOlVsTO9BOZu4
chktjDtr8LaHgHMmatavdJcI5vOqyCW/fqngSluFgj3/vjuJDQHFk3++y5Ac
FHcZnM2nButQA1d0PARoWk1TVsf4UGE34MHHD0ZAzxbnf6W/KVqQMxQ5fQ6U
6Vd0MLcP5T7MQLja+WOUhXtFCQdL32BZBSsk1aOzEovSPQvOMerJ93AgsldB
etcd6QKAUiT4/8BR73Z+XKUycHMVN+pRJZE/uFsF16d4KYiSnrbHFRohDOlw
iySSFo7LSrrYWAgbxWxV2bG4xHSXxv95hP+g0jz91dpiLPksq0I41Z1AvchJ
Z4/BaRAosZd3GCNpYmJiSebDZmT9FhLE4ZGUVPFCxlK5kn+dxfxSK0R3+GbA
eLtgo1O0UfX0ZRUJMxzdNBN9tttjssivHwKE0bJfbZQEy+yvBpesqmarHC8K
dtnKPwEqFiKs/I9FcCsgwmirSbUG1awAM1NdiT0ElckL4Ea6qicYZqu+aI3t
Omcx4NtPb0Tp8bJ2hScfjM1nZoyjODMkcu+QuYZauRoSkSonWKjes1dOdEiG
ZfRw3adetaRL+SynzOemTDGXiDL0pUOV2ZhVvT+/osiZvOsA2NtB0vLzhpTN
vojfhFpVUF/7JmoPEch1QRr8KJZmxTVvhV7OkWRbsrCf5yJiQwnpkRBYFD1S
Fnz/bvw30JwfKkgSAc2JyCrbTePvsRv1lv6Z7XtNZVlCz5ptj4nMa9i6+Yyi
rH61lJyiMXR0ZdZqCQ+FDQ6dRcASAZIQGH3yjFn1rEI7/MQXGcbvxwOlPh9F
X3yoUCrl9s0IEiYYiNwbINYnzj5sAX3KiQJrSQiMa6Q8c5dJ1N7THd1kiwaZ
ur4ngKLNlh2zqNGdj6aCqjkPAy4TUir3gTnoTLCXcZmg35LOV80wA3zoKyKk
Zryskva9XsHBZKh1YnHZaWxJudpZstlAYdpbfWU5oLDYDPTleDd6emddk+gB
igD/nUNc1bW5UPAPoNgbQjPsqdJBWOUrYJT1W9Mu0O2ccPZnICSgNoC2+Hl9
tQKv61eFXsjDcu5AJYlii6J2GRlekOcLx66I/uZaNjvz2t+kFZI3HOLnRnZK
b49Tkjxp9y1HLYJvgN3s2Rf70No8X3me4x1uIq/HqcFr4evWRtwoF8Nac85g
LQPM3gD+1xoWzQ+HYW/iH7CtoF84VnUpGa4OHBpYluvrJYdiFfKsqn07hMZo
15/S4T488Efyt+LrS404QmtKi91Kp7Qn5FHFj49P6dgP8CE0IPHM1xlI+Fzs
hskC3lE3oybSKGTCLcUM44OdBYlL5Znbxd0ZPbVinpI5mIW9LALY6AD5ij7M
nXhBuolP2tS5Afik9FhK5uCz3N/z8FeOgsYdEWNE1lhwASsfBKeMSFQ1+p5O
rgg8dv2L93XM+vb1MrFgN22CTS0AVxg1wcaRbfq3BpdZnkKnpecLCMiEdYDE
5G0+NTpbQoIXXmgwz1dJnnhtWz9dvj189s23JVqXPzaRPRihEjOmC5bEqxjr
OeUCNROqgjRp0YrIehPHilNz6R1tHKqykfbndFUq97sGO8hRWcqcjBYfpXYZ
yvoEDD/7v91mMcAxE9lAKbPe/WRms5h53/mmFdIEU1GdLAhlmflx7je1nf6f
e5c+9TFem5wiQOzGFaJ156mGz++V3PYFiTkMdjjmwgxBa8BVOqSuEzT3U6fr
zwW+24bHucFhBj4RGZ5ZdmVPwwHKim2AdoURy0odFHazCxthHHMsYYw54dqu
200qSiWpDPxZjIqigClP906UWJq0whzncJdZ1GeWJ/2uxxmciwzxvxoY6h7N
tTkhHTqtPmnkz4g5sUWXlQLVl4nABeDQkLjbGAqLlAwjmOegLEb5aftT6GRn
e6MRRjQHN+oi6NjqfgNes3nHUqCXCuN1ty9cp7NmN0Zct3Rcy9X9HX64cXu1
IDetOpFpA+XjbjIsM/qe8XtQv1st7kH7hwTVxCpVSVLE3gCK+NxFE5PrZJEj
s8+UTN4qM6uBWgeViDWyGLXybHSEboUYiBkpHVAs1MWCyzConimOAqpg4LBB
7xvVN61LSSHTuPD5QPfTPHImjvqH0e5+jhMBfp4k5Tpl+Jbe4U0Xh6nonzMS
H7cFYbBmWLDM8fCjuqcxhFYxHMhyh7u5Ux1zqdjKkF95gkS8ejojdD2RawDx
JGIe/tgVaend18g8A1RGtM/Xf+JHobL9BnA7AvkOHUIqCXgymLu32Qj93lKa
FYc+61jjaUjVexqCNahllDggWsS7th6Klms+ReoNuIlJaPKyWNUybBEVLmam
EkuQze8/QNqEgQSd0gefrLwQToQ0wVuwZn/ta5fCyK0+eWxcMyehWM5+FP9/
k7qJL+w/MF8FRp6xtaGJzWpKt9k2AKpefwmYGkdC1fxGLRje4OtwIzbCgp2I
xRvVcbNUOAcEifC0s/aMZc3XMnVhrc/IKYJcFBtwhZnsekC6R0LXid+wy06L
0e3fj1gT0ieuXg3vhXslP+e6KACj09wFzbI0xGDvgUfTpxIDSkNwT6efzK6d
NEGCn+WGyEFT+58Qzu2EGu7nZG06veAKR7nPvq6KwiFSxfb1OXKH6RxK8nwG
Vvvq+U+pTM/T3BOWM5lgDTtI0jQVSq/Ejq2ehEmZelZ6cdRmhJOzL2RkjFdK
qstMpmnJMP8kRYtY6mUa1cUHdBb6m57jxIOcdsg3Z5b39xb4c4aToSKuZbhb
HRmibk3sQ5B8CCt9lUhlnaZub/jUt1s8kZUMMJpMwj+kRLWBt6lvQpltNMjw
wQk3Y92lFctsfkUn+xPkPqlqHT/ksc4Q2wTt49p2QvjjADTuJHWw9ujTXDA0
xkGnxFnS/X6KO+l8jNaMCmBtgt3JaUfiSEPnthiY9b1csT2UJqve6B29UmO7
0hXGfDVy/IxCmZCcvJOer8MuTsRC6bk1E8T4W3aZnnKSocX1Dnzvm4IoTxOI
DIv5eo938zxdPFYVN7JyoWSfJtadgtXguRYVOAxh2sbijERfxtGiot9FanQY
plubrSJxcyhmpu6DJaB65TGZW+a2WAnxaove2aHcMD24viUNaK2QqHlsmpR2
A11NvUap3Y6WQghwHJRoWi7uc7jv/Fe+zVVQMgasLauXRZYFSJpQV39a96ww
GlBDjDYamINaU/tIlJ0KFFVs8EEqs4h9Oht1RteH3j9a4wLtgjYxhBrq7QRL
R2C/ROXu816DSWMSe1yooBdC+E64n0L8GRedHnTzXf/QPqwwNM4Ta2ilbiof
JuXKiLf65ssKsXdgFVgaWeRE3D0PTYILnK2MNayrqsskdrDim7f9kSg+KjJV
uwRouR66zuQ0TfJXOZlCVgQK+DAsHCy/C5A/SDMQAybHke8wVBG4ZQOL9CfT
Oiox7LhmyV9EqyWMhPkEG0E0OhjBHBjBbn/Dt7QMGa/Klc/3TFhcyGdgCFfL
23FoTMQhWtLWGsLw88x9ugDYhHrtxCJCDPGweMEk/VrcKPhai9RCNmnj5NTV
LwKc7JMcZkk+W0LggMSq4IfFI8Fx59CmeQ5cTJXWpn+/gD63VMbVoIt4AwQv
E7//z0xNr4wbk0lBgj14lyYVSocDPVQaGwW7IAwOelFTPwjdaltJKQu+hgAO
Ze9d+EUos9bz9CtYWiVjzxpk8Y4QGbD863N77dO5gXySqOLZ1zNQRKP6O5YF
LZeY9fri0L6+VzTcc88CnIE7pH8aBptJfNnDrbR8ROprxcRVGJ4j7nZDmCBb
yivYdZzXqqZ2QxddpKzFcjEgn9ScSbYY2/h6JwyxmMs2c2KmqI6Fg+bjVzjX
19PUU7ixHqFnJG6pPx39h/4aYcrYOzSlex6ABTZjaDqse6ZHTSAI8DJ39yjg
eWjW4ZxPWO3+8x+r7LAtzCdVFYJhoXwsd0+8d+sgumjgvGthxYT9FLJH01d1
PYEFONCpDvxnTqVN/5YMnWT3vH5fon2VgQrFOahoBzuaduhENGXvwEd0auQy
WN096Ga6LHxRytuGsfqhQNRjSEjNxqRyhFWfIZP0p1uMU5fRX5vemltBR6Qo
aXnZHPSrk4cLvLThGU32wE7lyKXL5AZMo6DMOsjwrlfCpAG+JXib6IIO5Rt/
br6Av+4nOmUeIzyd4OrZOuBxFUca4o8uF8JkxXOqkiSz4po2F6KfDJhVDrib
e9deYqQXW5BsTiwMXJ1LJ3i4CknqjrLibsPxwUgLRyYSjpoD/n0+hu1Xrddw
mMqhpHlANIOrKjJrH4aXvbs/pBO03lUv7Y6Eaiidon6qgpLb+DSz33NyNnDo
6EdvdNlxEcjY21Dxui6ae50bHQPBSbPttwNsDlv4Auh5tS2QTBoJEzAwlWYk
BhCNOUbLBy/E03yvYKiHA/Xi+2R41JAjAAM0Xr+leVS+4kINPnpiPkhgpP2a
3l+A7eFBiioLY7eMzcDmbGYA35faSrMEKLNrIdFMaYMiGV9wBXUoIWlApVIm
J/6ht7S/ysfSBs0jrf+ThNAvV/4Ki/VzcIlnRavxZWqrJeWK4gLDpxvwid3M
REQ2u2UJbmzFNeaXk+SfXd9X7Dpsw6YHocvdj9b9jYYlkKa1ez2miERa2V98
RqMAest/+vhiw2ThB84IQ4QsBcGG+PUIWz5xjdejidZ9L14ImVnMIEm9aVuE
fbTX2rrqFRH44k5XftnhukOY8Fk9QqGMTwHf6VO1yefiM/DD5OZFdMP99BJh
uJOQ9O4gicjvHdRToTrp7zzeJfZS1jx/crfPZXVO2w3uaXXkgEC/9bZNjQSR
VMfROFOYnUeGJTMdB1uvRtEgeJgEvFRCdpEdoykbXuEhPQr+3BFR9msur1Cr
Z+7hGFEQwJw/3H1mt5RfIezHii5M1J+66auZuG/pDXA4SD2ECFIm0hjK+uKs
WtCUYJ3XRDcRQUauEZ5CtveH+QZs3zaAXRVVhChlEVBdR4TduPyIyEq0q7MH
ftXY0e05MJYIGwSlVcifkU2buNgI/WcH8eZvk4FksPl6UeESeW8YwDfNyHK0
L1nyIbnRrw0LvE6ubU3Bm5a6FF8tA957UsJeeBtOeYgfTvLBQ38NkD7frMoJ
D5SI+d6r0GEsBO1sfMOJ9LJ7M8LilBg+SlAvfp4BIq2KHBbx7bt/u3ndgvUa
CLgKcwDg0p3ytXbEVdmilnl0mGrNz494fTwiMDEseiAKn9YgpbcYBToe6UHp
CNK4UCQIdxqxpgm4damF5F1XfqTrNaL/xsa5OnyXNqUSD1IL2NeAJxIB3/Rd
7AOzxCvQhaWQ+AevYhMwWOkkGmATxWgy3C2uxees+mGtgChj8Zu1JL4WadHE
21XGdnqtur16nsIbVgjFYO7kh8huza07qer0QnP5ovsDC3N0os+BLbQI51cy
jBKWVknqapkOWhL55mdPMbljY9XW5Xr3ujGHB7L8QbPmnBAQUXDnF0HQ4dzP
0GyWT17WUr7lVVjzbVk12lHwnv97bu6dk+ulH6DcjQEhmL5I0QR4GYDP0km0
dmqUrdA4EFqSN1ORY1ByyzwE5k7LLC/EzmU/NjcS/nDvZjDoBdrlu6efSIaT
x/snuje9uz6nZ8uKcanHh+eqL+RPKH3dcoWsfzof/3h0GFdDl2JrUNvEf50D
m0NJ5VqmEqAViWMIRf/dNiq6wsxJ6tOQzBanlefOAJVBzZyu3J3+ZlIt/j2I
mCsbOcKFmSdxmUUJuDPW5RSKgwX85+TByhSYsagGaflDjSiOSAUDoQQIwv5t
l0zNcRftv82czH2DJBNnh/al2t3qG/6kyRqSXDimT17nEgIJryKocx25hiJp
60c6iiCrnIldG2QRCGsQTW6hAJuFSqzhHcKGUcyduVzpQl0/je5pCvb/69+2
0aAYI1MHYFiiCs3SgfDdQ140GTWgHyOhWODj9WRQIjXDOxF2SrzR/CVTimkl
3k/BMK4fwrKVRHoAMl5Gi3HbGB+BLKu8EVlwfk9WLOc9x78g481HwPFUnNxH
EKm56N/emrWNW3OPs/iHB0aTBD/6cY6pGJ9+iblNLcOJBhXgIKseYqUg6Hhg
LRlODHNWTfT81pufDoXUiCQ9y21eUZnoHF1fGl/G5LTagWNRlgDV+7zCFMZ7
3Lgdt+YN3zAyKwVXMH+06hIFEeKhrWPJf/djiVHAo1Se0W3tnx9edfNTbTjB
PSdQlhU9VxZEz40ZswRc841wNQO+9xunaTGb/asgFJF2qxX63QXw9ffLMc73
bAnTTdrZelhde2DHz6mKtik6W/ajSDGOVR/t/mTMIRNKijvIz5SIso1ATypn
XC0juJ9RKOFnclbS6JBRnYEaMJ1tV8ND5u3PRYmOlpFKZy+oxP7jbirWl+jq
NY/rDwpZGT8vJj09DCLntdEviMLPujGiwZdj6YPOuJ3m/VTce7JMXOKk4nfS
gViQuB+V94Ma7igqhzZe/moLH1oW/ygvnTje7jyqC61IiWhGa8eayd/pUWmL
Jdq2ActwZBqJEMLXpHh7JWH3VCRHgozSGRwPdnrFk6/c+uhaNZ8QzsX2gWCE
Fuhxe/OFBV3o9RJz8AM6qrEwrUxbkcB64avJFGNhn3oAum/6ge2K59PekgHD
zhe/GuMaZ65FfOcwxGtEJmx9KkC+Ke8VKCtPAoaL6Df4gU9gkHpoHTMp3mkk
1aztMuk9t/XnTHmCJ6c5vICXqh0VbihK6fUrha9kDxSP4sTqTllDi6/zV1Vr
bk4jE6TzBIKhEssVM5oQefBiO7jAQXJRkeM7gBL2cYSYmxhem8ralrZkqF/x
S/ElcQVGk9z1SY3T9u6BfeAx0J2soEGT9tCyWUkxeJhuJVijY8ukuKbdi5+S
G7h7rgSRu70nCQkc3TdVy590ZbmxME0ApEYHuC0uQX+0FdPFZWYZ9RF6ehh0
DKvLM9zKBBwXmzI8VWR4t0vEklGSuCXOf0j6DHRiwP5FyTwm2TIH/UFp5asT
NiC7UiG9+lCGVvxbOns1i+6WGD3DwFU3+wG8Gte/p/pW44X+5ZTbuwVnUnQR
0xOIdUYyPSDkZHQ0jigCYWAO36CPwkOFnE9e9de/GeZKaGTZYeDl9wKBDwrC
YavTbcBUFyT8mGcwxNk3X7q2lNNA1M0PAQ9lmVhngCS1nhBKvdlJvK1/ODEt
UDOgW/0aC0QfeOGoqZ2FeAqP/6NCE3f+B6eheLbUv9bUy63xA9bFB+C4K2kJ
Iw+JuQfpDlaV+pfX2NtOi6UG9cYg8mcApJcTF20vdz1L3/dgbv+5U27SyVR1
hWbKD5vtZnP+WrJl/ZZRlHrLSYsX4cfMhu1v12wnDaD/kg6c6OlBRS0b+dZd
qGokBBvFzLLVbl11jy9WjmI+fnnnAoNZO83kHxSv3FVSOessIEMOEea7kV0c
SaEdVryxUG19P4jkJuL9B+BTA++lMxK70eS/IaRKbN4BoTT3bNUKoezmChW+
tGgV2MgewKKSU70mj2QySPCq4U3pG4ZSiMkqaCQ1RDVIK1pJRGSBEyy/9D7p
vGmKCLqP2Qxlg5xu6Ly8iPrJ+G3WXi1m3Y8dEo0tIXi5mNctxsUO2QLY8vY1
Qu23q2OQqrphjEj7CrA/bUIJVexFzwCk+GyJiktqh90lL1OdSotTZ11qtK3q
iKrSjPOnXInQZH3B1hF7WOP/DrXKRTvvxITYr4I5M75LC/TxEFtMgmxtBRJo
jsaov/Ax5wt39xm2W2QFgqgBbbBE9ZCDBdKWclZ5LaqH2JYqmg8AKIZAuM2+
iOkVMVFe2ZoA8HsoevMlD63J+w1uEFMld1qXarsw5vPPOB25/aOyXIuB69fI
XJaVe3O64WCcd96fKb/9GLpNVhgBZUKQKoK/YdNtsgWHw/iL70HO7CqPYL8A
x6gGbqtdd/8+h/xholEhFDXiBuhXyuHGe2vEyG6a++ApAYw19VWx6/0DvVhV
H6BcoWXwAZDlamGrRPTvFcZ5y0nLT4HswZPZbogewFPpNUdix4w+EEscUQUQ
kf9yvD8Vn62jcq7h4uPUTW+gVaFu356yMwvAC4pprRAhDLb0NVpQcDktNry6
7bI4JtwmtGgHfw7e/73raXA6PYmhgp3HOYVaDPGHyWmXl6xwcol0MVVRU7TM
LW0FVTOLL2LBOpkYBA53p6tTZuZFuGEj8Jvn2MRCOGBD9eweNPoKXaXuAssd
fHjnojFk3HxN9gJefd/32/tRJx073dDrXsvNAbJDazO30eJQT1gPqoJgjwSv
fJzu06bWUCPfBYUX3x3Y+Gu55YYBsnGFX/flWZ5YUe0dfyzSyit6TCixw2RZ
CYhZJVVPGlMmtfTVyYG27YwVNuehJCYJ49k/aBgOdx5ZRyMerVhERE4zwxgk
q6lbn+qPSduLchQ37pSHjMIPO29pVuFd+2Lk1nIZsUYa+vqGTAi9KFPFxYWF
mJuKxaVIbbqKQXO6EFW/AANX2vsIspEAadOF9UQT031fkxh6ioMHIPi9uOzF
CiexHGcDSOYgpBA4DezMslS4Lhv97JL0pdVAOtb+U7k/t7KBQZwQCowEBGwu
WxYSm6zoRzufTG7924pBEZkQu8BXFC0bfFBSNJK3rhIDTPWTRLj68S3x6zDU
MFrXuC1pUaDGi2MShPuExO+MOl2A7Ri+c8ocenKurwfaOJaOrvAn+B4Z88PI
koRSf6sv4FOE97kBmZKqzDrrJPy6ZMEmSXsoHWnvcjkGKYbN/3qUWG6CbGri
qvbOP65KnRmuokec1h98N3X3HyfRNsOyZJmDBdllJ0FHQ/aQ30JazQ02Ai41
XhRUEtx6t1oUX6gtzZSfmJxb73ymkcmitWbxvSpFbesYn69cq3Zzj4g5s7RU
IoO9vtH+vxXadL7YSNT4o8CmjuEqH/Ra0SaPEYXrWIJopl9Y4PvYTi+7MgrQ
+i96HY8GGd9bswKljx3nKq8p6mmlmsN3mxr0LpOLBmZFTdthys4j4OjewYCm
Px8244UTKvglu7hEHEjXz0MRsftSW74hh9M/zMuBDjVC6pl/FlCnCZkkAFs3
iYd7c7q7mydMJv9HpicF/fcTnXViEinNM1DL5EJP0YGzrRpPBruAMWDXEdLn
NU5ysrDwXy5OY04dMJ9IRizpre6Ly5+NlgkSfMm2/FIbmrlHjELpKuN7rCxy
ER6nFev407rVGPeT/yNFq5n9cokio06c/TcMcb68NtfVBrDwMVA3rmfPBOf+
nAdfjMsHMeBjCAn1Op3mZsZOfv/ulEhhAmqozxAPK0Ra3hSVqYtricc9ssMu
A+qt2/p6ju0xu2KbRgdIHZa1BJLungDD3fcw2XizVh+GZSec5R6rrJ/RRp6k
R0j+LfjQnaVhFONYR3ba9Ph7VEuAcslklt2wm6jxmht1O47fr6ejyB2YK+DQ
BAcfe3O29qHPzdqFbxObvaIjGc0MM0WA79kVh6W20wES7RXJ7l6vrM3WWC6K
jKYydJtEYDJ3oxU7oMIooH+oUufkxTvsiqFzo8a/f5ma+7RfIVB3B58txnQC
5ywe04czJOtJAQWWs7bKHyW4/+5z2/PXmHyCnxHg7ahNTjafjgh1o0vPlNWS
DmMi+etCF5AYdWgSJ3TCr7eYiyq42JOcyfXeaGEmAB0l8trSm1c7ICweJ2VR
1Xu6pX2DQunpY40+Wtk2/9yR/zz6Btort6WRxCPZt7SHBZAydByrOLVAeC5R
SkyibOjHP/NEx5UhhTXRnfwNDeF0HpcHrqDnzX6d9LzqNLaYOa6bemBDxuxA
1nN5HnB/tx/knxepVnBpQy1lbDn7cNlJ62/YkvpDmzM2SYI6/AEAEUPfNG+k
4boVw+VOTnmRDUFnt33MVO7tXR9sHjnIMPyN7vaARJCF/WrDIicTPKis8Zyf
4vq2FqUtehFqz2jwaaH/eUcZWk5sRrjuOW0CZQZ1d00PAeUjorSCTY80uOQ5
GGFGJMLHr+AILDyvXzo5/NdpCuNUTXE2NpvYVCHCHYiki8THnse0W3kKCfRB
pXJ8lHhey76Jx3PkVDLBTtfZCYRE0Lq11NcGNdRepMZQmPoBg7BKYgkv+/mj
6demfpbTzwwcjssWrDmOly1OT7Tlph5tk25vxMRL9pz5oys8uYkupzgAvdhS
Bs2isqm/d6zPHDw42s5kkvLArB148M9p4zhC8qn1KFKd4C4gdnDRPKFKIJA1
poO0Ozv6ArkZ3muXVGrVGRIIW5UeCnfep7I6SHMX8zT3F4nBey5buTmm00RO
euHORyHU1D39BID2ebT09hBqgD24gIIltCoE2h4zO59M7uSdrvZgnoJsB3gf
xEUFIlpyN0SRtEhTrKLdWwZyT/5EnXvu4/EKK25b7ETEwwrupbp2SbLhsxsa
WcwldAyC0ZpfKtM2T9bw3wSZ3bIMVWZeEKCjvhmkz0OF/a9xtbl5Cyi2b+Cu
5zsHZ+XbM0oWRTzRXSVBL7ZMdxUan4tENCCFCiQQc+jU9VD54iREKBd7hJK3
W6z3Bj2VL8qppqurZk4Xq5rRxIwjak/JFBxXdos9YXlKpl+xrBkqnhYXP8ji
pbXID01MjGF0Np5qUTAyPGPJ2zA/qbwa/SXNEiyrJxnmhdogE9mp3BcGkdQW
IhzYepKWo71Tamn30HjCYrqqBDEB/szG22YhdpGfwfDNKJMKvcBaAJLCTNdR
tcNJDTQkx21e+Up7nUz7zy0iIXlikL1jBlCSUv00qWc8qva294EB7MNAdIWt
ZmHrepEw5dq+pRtf37sJ36uU6JCBUZgd+XrC1O33mOO/mlmXrB4QJ5E1Yup+
OYMj0iPF89u7WEotyYyDhuYZ8TDK4AJFYFI14O2oYK0nVUsvH4YertD/ghpQ
Kon5pY4OiVlmlEBCtDDvup5UkYtBuy5akb7guJHUMSxnolVMvOKALF6l4puT
oUcnfIcR1D0BxQkHtfAk6N7TsSGGD/I0QhrL6BVnCOih/CbVvR/FDVjZz1eY
cx0Ms5Y6kubr4rLE9XrLhMoK7O9Bd2cgou8pg/3/B0tOHly9yaPz5/zrrqh0
TCIKK/EQWQcNOIJolR3TI5Ra3hFqp1ioLWJXLJ4b6I92elQAYWyaTf9b22x2
FirnXNc6Mhc5w/63zGrPdQEFcWpyVl9ZExntMT83exjCf+aqCGRmJF85CBys
ggSbVxyWV3niRmlKPOMrPe01DsqxK1UF81ojmeINOoMd2LB01h291i12Ztp6
FM036jSjRSnmV4m2DRmPmM+nTqScZMQqWHy15OpqMFJuL5vuM4mq6w5eWffY
z8qyIbGiktfBV6flNc5Sxb9+5vBAt3Ihy4eOTvFLOgdCaKNMbVli6aE9p67d
tJa8f4Z21+K7RgjdEuqN50AcB7KWvT1KGIo1Q4h+DFLiaW9rXFsge6+SMt3r
to0se269g1Nz0gURv1Vhux6b0SJxCxK//ZeYLj5NopFT/NjJVLhwE5OQJ870
aUzEhiE+Tm12x7jNJr3/5wmuXVYtycjWVMolmyRsGKX3YTDw7Ks78fJbPJwy
OD6MHyzglPVQrhwjjzDt1tPwYlx21tQAYjZnyvOJJtZOpNOlQWoVJAF5NZGC
O+E9gWAdi23/b1G0qH7uOI6xiAewzqVqFuRvDmALRFTi2z9sKAKMVztKitfd
WhHvE0uDtTq+smmEGgIItZ0QULmFF02jDbn7Ig4UXW/p3HFLwDVtsD1bpvl4
45lp3UevcexOBkm36MjRjFLNYdtSg/K8PwS9iYE3dU5LD5OgHI8F3XJmvYQ5
+2SlyWS3WHxm1TzYa1Z0fyfkCFZy0T1KRzHKQZ5f9nNgdNgSLJcNqzzGejKx
OrkSUN9GdvCa98FB8gubWq24v8fNG5oaPaKk1hM3y35oFyg1YeBKwRsC54Fn
MCG4CUwWGggHU0VgPls4hmAT1S6vPgZREP72pRyHHu/uxL9gTPqn/ModaOlt
wbhnXNsg/orChTtVEKkAs7T00EvpNEvXsdR5XboWyzGXTXLMIa6db0bv9b0n
ALeiyEF1aC5iH8UyGrUIpgHytK2IrNDZl7rudEN9TQHd7vGyksc0H1vgTG45
+MC01ktOWtX41qs9XJRMuNfR9J0tWzxZhWjRrVYM0i0gBPySYLF3eZ3jTjU4
QfR+UzouM0ZfWOovdUFQoPBer3oxo6o3KQJDcnp7MuWx8Uyj42ZsKX4Y+LBe
1K9czoBouQcVl+4XyE4CS/C3Wh2rWFKAJ1mV8g+h74GUyzAd3sBBMYEdyEbv
q7M3TP4GHFUG3jBRQxDsY9xy7FHYfissz82tlfqvCt8ZUtD4tul8fbFNX0R0
S5zTP59bcTHtoi4q8Im/d6IdeONcFLoigbGTnKQ0G3xD3AYNAIJhD2R3nmyA
Q4RNzMEZbx2Nz1X2RNh+FqeZM1QChQQN3lb+E0olBSwqdb2zjYbuZARgO1zq
lKiLIImW4Vx92FeBcuRjy2Ka1bDIgPDGda+8xY6bzHV/kWLlG0NyjeUl7SBc
O23WX5HgTes/UcW9pgJSVqW6HS/wM4HEkElsb02muYp6XQonpD1hvPYt1vpp
7oKgU+xVKalbvAMH/rlGSQIBdypoPsxOpTjql3MxMLSZbVcq4IFtATzLLz/+
Kwby2EAa5JQjpfU+hbUxT39cceiy339XviliW0KVS0EY/LdCC4WPCXxxdVpU
X6SrvtrSpajlUFnX6UeDf2qvya9u3xQysuCrY5ia7+AIArw0hZVcUgoQ2OXd
sQIFlDvlnHMBtk9vJCnjKD/CKjZQEkLcj74PSaSpthKLEHSr6olRW90WKAny
8Lpcu97Eviht+LaERUxV4HrHbpWGFrSBERTaR94tkKNJCG/qR8FxDhSN6bAT
E+GVo3f+sjbiNkxtb4DW0zeVZuMePHvU/Xc+M8OtKfz8hWz/dC4j6xC7Lbg8
U1ZAk9CFFwPo8rIy5UaZ+1xT57M/34CIsIxsbhuldQeK6Ob+dP2OyvCriYsv
vfXJCx0AMUZCw+VjmLIu0BkU1sqR9761p8P04zSVxj3UUxlZnpsolaMEVDpS
JuMjtuTuU4BczwWgG2ZYmjiZRAQBurC48xtPyWr96G63IU2GotzTxKNj+Yov
rt+PIyb4/EBauNsb5g31ktJ/z6GwHiHGSz+MwQ7Rlaz8MUu+0pFTo1by43uX
/d9mn60Mq/VNEWNYUEOTv6NrjxfPrJykP41SkW33FDRD9ixhexD5rGH5fiss
uPvCaGxGodcNSbgL42QYL8oaAqOZXX9p4BGjdghyj7dL/fSOuOHcaf5aFk6N
3uhhE+smm1+QVz61ngH+MgVCr3cwwJFqGxYlMRtmMwVKaEhDXYJe5PXeQqYU
lmh3s+26ZKi7oygag17x/veOlM4elgjhdi14hBfFYOjV6uDUrEjqL4Jdys9o
hCCXKvL1ZTWwhhcIybqTERolQ0MIca+6Hr2LtR7Q6uXOHNJHlpsyXg0vzU0C
TsFzWrxM7c7ROFEk/uuPL0XmxXsn9uVxSYxULv3vK7WO9xpgdIwZ6npLbdYW
PTdGGoB8CaGqoAb4tuQky/eUW2PjM9mtIHot7ycF6Lck7220Ut+1rw8A44Px
clrdTDvojzdfweEjwYpkAB9I/5dVSvPb65loPeD3Y0q0E6GsksucAbdXs8Qu
DhpYbyBswof4oJKwLohZJcM+VVbYp4D8BGqYZ0KIW7sw6yxAetAoszov4Owi
uRhkeSojkdUP9xn1a+CVGzpSjktpS8LsKNE2M51st8RdEdQhDWrOx+GfA/sK
RY/CkG5HNxnG35+6WOwnHE0JCYIVsBOekM5+y94mtW4xUFEUTsNFWMvwMAww
684AJ5prMKbqIH8dMApQe/fe/u9Xag2cYWV479WzY/w9giNN9vKywQc0B2Bi
UW/rJ3sy9AWy2ffymnX5otzsHRmC/ANeiQlRFvpc6QrgGGbki9mJktfdGvYG
1lJEDSVzES/k/JcMj0Kyl1lMuem6ki96Zw0BjcsMQAyEOHUBf1ZJs5vr/biR
OMLULN/UKbJSSvWclLmneafVPTdaZpe6Y8C8OdPcETcePLuw4XQGUEN0kikF
2ALw5LpZLaoYIiWZ2xJSk07eRFvCuJNltawFlaAtPZrnanPt1XkUhpIGvU/P
YtKLUkB10AXUtWtIwNddWZ9ZZafFAqO3FBbw0vVrm5JNc0/n+vtkZuo3jC7Z
Iog53cjXEpLQCj73E8ajOwPvNE+N+C4xaOPJJ+RHmCBDjdejhy/zD3IGCaXz
xyxXiKsMfp9lYcQzKvFIqHp3VuOPbZcTKg2Ddl/2sNXVCE7EOHEl6Pd2RTPa
kf0sAfqI60LvtZlt02lkoRearURH/3qca6oi2ZZeuUsgddZ7l2Ycqo8mjkIJ
z9rOmvYq2v3ayH4OhrZzP2QWP3lGhYuJQMUjZhe5u1DKpvhPyCCLcY6eeZ39
6yDW8nMkZ9mtZcUoPgyeYR+5MjgECRG0bQTMUOpTcvLx2p8Hj0U3q6wTta15
jmKa4nfwqmeJzo7VQnCQlh0B3GmBxSHqL/+utFvajRbmpZ7s2q6XZYS80mV1
vFUPOD8e+vxMqV5qJzmzESxKODtonzSpafbzOXfSqFBKSgCD2SR5jhrcNV4p
tBnm0IlZGh7n1xFESPVrVmaxLXhEzjRwoY3F8lY8MykCJO5k7QGt57c/oqqT
DgmxYC4gh8Cqs6AJ1I0hxKvl1fS5eVU5LswZ4+XtUqjLJC8zI8fYuh1shPS2
WWuhyE45TzCGCVfyN4a/gljpNU53+vuT7utJ7nR1m/AxT5ANZTcUlSlyhJpV
XOx20C5OFll0nP+SRVNEzBzzk8O2aWOWeldcoiUQ8DmQetBtnGro56RFIlP3
Rdx37+qaMyu5EiaZ7SqSxcJMw7tYkDzkSdQRlEdnIMyZY020GXye1BjTXXdx
jYB9DkLPGW5hPu1ngK/76pi4VgPAaDsoeEabT2YkjCpiFZ5XMVw1kxqqUi2Q
tlCp3hlhxEBRfXD1fCnG8sh+a1MZnnv7er+0CbmxW7JC3LBaFiOqQA1CXZ1m
+aOSdiYRWcHL/5edY+kNry5ZFEaDzShjTpubT5wyh7hIviruXFlsgpsGBJ4K
aE0CwQ0FYda7tEDZOiCy5rboWKvxny2DTfcxMGt5Cl4219WadnNWWDOAbrHC
DYuqRwdA64dFVUrdxB04/oRlZjnFTvOoTvKu7imIr1W6BwrVZfQJzlO9xSn5
A8oUByIjV/SPmbak374SMYi1tlXVmtoNyE/kZ2vcL720teRNIhH6aicGG6/N
Q5nMDsXaFCe288K6SvjWkGmkedbnNUKuS2YRbWGP3IEL5FuiAihnjpRlJT7r
PUO0ejWOCkaBkLqBw70BAjpVbTLgvvrBerV1K2BIfLr5R9YofpNgQOy/iTD5
vjhxYUNUJiSWbZhX/F24QpBq2ZKdpCeZ1SoV6dxvi1S3YZy19G7d+bitioax
VU5m3jszWxFZf6aVaBZL7hZZhyFnI40h+e7Gkd82VUyAtYrwfgT6nGo6bN9T
rJieiImi2hNEaeZyKUVWG8SuVMUdCNiqfHeT7kKb3iNqjN4sdHotn+w3DNKV
G95p8P6sQN55+07QuQxZfGB77vVKitC/HsR2F2D5ijWtTLs0wFOBH5oFRwQy
HCwR8MiaSQaA46mbhV6nFg5e542CETkIphBBaGJ2IJpDze0BniU2KxAXMKvT
ruq2ic875KdPAETGiA8h5SoTpKScc+EdWdMTT3LC8jIN8Z289Vqc52hVTwAN
rTspdQb+Cdh3ZCz0taVKYCPuk1KP9UmI+rcWHzGYwXp8ZRVmJOf7uFzyRNMN
yVRyahxWVQatJusI4KlaaR9NZ242DwnSn75PpRxAfszO7UytT0qqzVjzVlHL
BthMZ4x2OZZdtHK5SPeIzFNKZPmHIPl0e4HZl57nHohgzfifwL8roBJEAVoc
iYasluH+07rXuoX/e102LVRxnulde0U+MPD2jm/I3kGrNbHOgqEeBuwBiU3M
KwiRxTz4YHh3e3/7Srq3xjPK4/DhYvdb/vc3/UwN8dbNERg8TkbA8g0Px5Yl
aZBMjNmq2nF7o6j74GBEX+cFBCKVZCBfCQSVcOzpchCR7ZfmvWYXJs3/nQtr
+UcFhfrDmncneS/AT93TI8dU8j9xGQdZ1yoFUHyw7lXPm1PnKiO7dmXdQA5Y
+8IFfO2dCkInhz2OFKdqAD8iwC2L5pbk3lbh3D8T7fwf7EKp75PqCJVj0rps
rcwcGb/BkEJjgW5WBNf55ys36Q7MHRF7LXCQlQtPwtQjKgf+/WMKlspeniFm
jSXdoc9+VADlRtuFiUxO3ZtiW4zDs0a1XdC+Ybrh16xsZ7aZPWXOxiVegWa2
LEg+X6yJjyP4PX2lSdecLlKU8x3VYwkzjz2BpoxD+Vs6L0hy19JCD/j21iIf
X5EEe3BlL0xoQ2fwwATJSz30Gkm+7+4w8GHlATot58EEzG1Rxvsj9SXO/NqH
+5Hj25OxWylhUYzJWNdHImNnhDYoGD8I94vHEty3k6I6TzTRxHnTZclqUTUm
aTrpW3gC7jbV7g7g5rsSdMUCkbexCwaSwDwoP8ZgAxDLvrnI6jxVVPFsihtW
E8f5R2v/f4Ag3Gr1d1QDVgs7UghlCqkGD5ZnM6pogWhqnjB9+k84UmxG35S1
knRnTcRDcpc9qitMjNEqZV207O27FDUOUk11sHgpibuRTBEQcEtByLUsPmYH
V4E9asqpd/J+OO3DySubgvxO+7eb2gYWH4IimeY/9UBaUukSyK/TLV2Uil5b
GcLVHViqdfalu2c20YbE5QkLcrSprBogO/T1RrPgAtBhdLYmjv+BBuZ/SWuQ
awH9aAUrKFw8mzzQwouTnzxxqq0CBNTLa7aSnijQc4n+OEAnMHukNME9GDNN
s7jQnxwYrtk3eWnpqwaDPOVQExuj+ExnocfpUOwbXsDkjxqMFWkK/eFoy7I8
eAJVvoAh9ehZOjUNlHIg3C7WWhanmWjUZylZVTB4yvvoyUFajGxqeqlFu6Me
bTAoUPhbFsP+5l6F0d9BdFQHuKmw/2yHOpnxS3fV4RFz5Q3nX6+e0p0k7c4W
axeOYJSIAziKv7c9cXafsagWgC3xmn3q9/YmI4xTwJAcuPrseTaXFir6oBYC
JFf5AYQ45OstyTiioc1HgfkmhumesDlPcOlevWNNWqckRXL0F66khQ5QVStH
fp2qZ8y4ctXwiPlKvTdTvRpu0yuFm07wLH0qFGbBkITFRqVI7/rWzDkPsPcz
bSxkqKY6Oi9QAXkBJb7yLIZD7rCuU+o9+prfTOpTmkZohc+yOKhCuOYA9pPX
num1R2oOJq0d+VaeP7W3uceD3EGU1728J8y1wIOXJHkmAjjU8NraOFlhhUhI
J4FQsRt3RAIWTC7kwvCMhjeOSyJROqULIcKcVBQ0vAVD/49Qfo0t+xrWIztk
ZPieQiUTrrbeulvWUzENmVuD5Z9rTyYU0Lx0p9R0aPeRWGzj9hJ55YHN3wmY
catCR9mqfvNcdSyqfKZSpGys0sp/0tyv0Git/Cz+6Wqbsa2L1fSWwF+IPC/e
MU1x7HxNwUQCvMTQDmfGm1vjq5/QFHtr8apqwcT9OVHgnYrowq9xMHx7ZI4u
XkL1SQtVwXtqjP37V/h/PwKqlddNVWvaEP6EC39A/V1QH3d116cDh38kfEPH
+Q4KHmHzQ5gt0d+umTvq8kjnx64BUeY4DKdPFG1VKElIR075OfSzfKoYwX7h
hHm0icqK5vARIIu1jyW323nXLOzZRcn+x13I7IHENxXMOnAhw8C7OhiAzXJ2
yTytyQOWQ1x+XXcpBw6nAAqvon3TVOyNCO7I2qzsqFdnqXSb/YW8l8ztIXFr
KJwIePLTekXXI+MtUm4lid5Z6OxBue4VsRJV8sKKaFcGzt9+88hPcKiRv6J7
uaO+QnfIckZxofAII1fx01tXC4fkAj53rMFk44Pse6ZwRiJ8K3D9j6mVjPv8
aAh0Ib2uM/22mDHpSOBl57zMzjXBr+xaXZJQ+N1NC7QePGlnI1DpneHE/3HN
4RyqnXHpWuf+U+8pC+LDBd+gtwgn1n0KEuwCXIea2Oc2RNf62MEfIe4yQWhw
D565v0E0md/kHULoYuRRN7yGzimznM/kNwv7e71vDZr/nfmmrLiixpD1K9wy
vIDrnYwqfL1UQuckz4QUxWEdvsf3q0Wpael8pfkZFa5QPlVXG82JhStEsejn
cEBXtvO3rPiAPR2U1RpGeXhECoHwkP8pLSfYYiHb31VhUb0XGAdoCy6oyc1H
ZzOZeXv6t/ZfOUA1/sOuGNBnebBGZF4rA4UYQ0ih85TLXQXEPXk/IxIzBWu7
nEvhVqDo9TGVDUadZhemPnuVMGkbBLZh13itozFrXQqh9qql11qqFcyfOMjZ
24EsaeqjF+NFkME6srfgNOE+vuxRgQ6DUoTbd+V7kbIVIi7xCQKxIsUnHPCz
fWhKtEuV4tvucF/ZgYqixrQAN3ETXOc+EFMBBRzw7BCi/zEkrLETyVGIChOc
oF9BRrVlQaf9WUpKmas4H3KB2JhFO4l3HlFUGhrYRKZEqb5F1YhIrbV1BAp5
jrdyLIrGFar13EyLiaPdD3W7MMMT+xgSpI8VotMdCT5cOT+YNBFaCaRnLumr
fCgJMflpc7NiXQH0rTLz7AdKHUCQWRT4O3KBMe27MwV/uNth8ZF+6qb+EAPT
NbVG6bEMB9EQsM+PGVlyCmG6YoK4nEjB39J80tB1h6IzyWZ2WkDeiFwu6cqK
YDjnXazNyFOw669oxb71K7xuoF9CTF3eXIUksiHxmIo8pEnwO3JE0dzNWoXO
sXw5ZSE42cleeOGmxxBfv7r1G8ifrlNfG6Z6n0yD8j6TB2pdYvrS2QyOInAb
TE6UXoKd6y5RHffIDPmIv4+mUhhUFZ1p30rSoZJY5fTpQTFBOrfdglN0qQwc
BzzvcMVBxAa+C8MCAYpjUnZ6PFEn6wcmAredeNaTrK6PmjWJHW1kLta/uX+l
wxr0MugI32Qw5ahCbWQhA5NuxhCfXddP86r5CzSRCnUbhylpQe3LJmfp1MCN
FDaHqUZLERZybwxuOV6GnO+b4DXZjxgVrJGA8Qm8jSuAvAtMxPsFvRqaiU5n
x/0PXC4K5i8ab8OEXhC6jpaJtjJAJ0zbBIl9cgtd70frkSAyAx/2tggQi5+h
zTwSPk0P02jaSV+SQY5gWL5DE7mf9VE4D+Yy70qKWsvrVgN6Mt+FTs1Bcsgs
Ce8659wX7rd77xWco7ke4uEsM8zlkGWOmlzZNIsMtuKZ3pvqhu6LZwg51Wj9
7kQUPX1BhfD1WK7zxvRyvqSjUPUpNsOUBWMzKX9gq+5dlBUu31pzflJaPKYg
Gu+3hnFfOkOIycKF7tPnNseDKJjwZJ74YQT1HZW3XY90wpTiN/lR0GoUVdPQ
HrMLvKVl5qFdm8sXfXDq76qGZqQfKZwkc8fhew9x8XhpzHIPe1Fles3fbMXE
FkpLT8OFpISxxZXJejELgKQGWvHBqVM12HQzzYKCGPQG9RbW21GMZUqWFU7s
cO9I1vXw3asfjyfo9pH7UKHY3/NyYWUvxmo7P7a9yXj8xE4TPpgYfm+2spQ3
z3xA/BZcTQFDP3p9C7w5bYykfO6fymP3UEjvqKsb5cCb9yYEmXmjssd5ojx9
l8d4WWDbcnrb5VLIsWmhn75qvZZLWicjXY2ZnnJ/gDdxsIOOGti0fEO9atFi
jPUurMmN75u1R5qTE1V4p1XFaFsokFsgqdEbxPXxZB8lhyQW+TwBWo9ZO0br
uxwpPDfmlaA6zikENkhAXcNLW1mivGL3k1xd173EBhtVxfvwhnz7+trHpXNr
AvE+okF5vhhDpgeOEr4FyFhKAE8TweFSSypjmQ0lpjME1hZdb4nhy1A5KW+C
prS1daTgyjZSqfbcBlvX5JzWqRsHoB23IUtFmAsxITupAXpNUlRayremOk2E
lCV2MAkv6YwPN374mv41JJP1Bl6pTlHQDcPNuTDJ1lqZKGajFlKXCMB85k4+
/ueK8cvNLTr4214Xp5ywBWNdy7GUDwfB/EhZCeGwiQY0WRzqEuVouCXQ0a8D
m7pmLHxdMRPzW2q7OiEdUqz3AqSG0UByqM5YRa27jxVNRF+lAdcyYAs/ponc
RezV34AEUaSsC2C2lXb1BrniQAtQVXnaioO9xk9wjNFfRw7PBcwwwNUqe8WU
Yug1uqleHx9bf9Ep8KEp1oIyKdmbVTlM6gyRMkDcbKdegK0mmKQEv4TpEqhi
t4SJGKoKMMNJtuU8jNjBIX+MNJrgUUV76a57mLOTtRmWLCuJcwJrgtUQW6jd
oiWZJJkq7znD2/klM8E+n7Lk4UsvG+/vodtM8SJq38y6luAhz20LRaVwEZC7
DeoYXREYuCwYb78W+zDZa6jPM0MkN868mfnhIErTqZt6slipcjkzoCQI16D1
tMF592pVWxfe46XYB8y2kM7ufnQiWS6UzhdfjnU/paN7RgmrrWkXi698dX4A
T7pqw0fx148TUQsHU7dzWTQo6oomzkkS0QaCLfGBWc16Me5anwrOz0tRp6/M
RpNckUWJqW9Ym9w71khDCj7EP/pnv2HXIUNYVpJ/FyT5SxM9XMttAXtbhm3u
WiU4EQJHRo66nEqGv5yNs2M6jN1xT9gE44EQPcL28NqymZmOXwUWtHGW5uvz
pOA5ZOGRbl3X9AlP712AVtCWvqxlShvAV/WZtkR1TsSFOrd/V614nS0xH61e
1wa2g/qF7gttnrBTVj2PNU9/69BTufkqOxGd0DBgj+GGHonD99cTy1BDDP0c
/hPCZr1jQEkhiQsvAUZ1n2mPfsaBKQkNAZFyqy/+vI3SxO/yv5Vi1iZpM7JE
ljqzvzB883HS1Se8wirmqK8Wlg3tuoyiOFN/aOoQ73vqLNF6TngOFMa/XcGt
pYoKGGLrxi4rWN/f9/ct1ktzWs+NeWWV0udiXYx58zL7cQHl4wb9OXyKZL56
zo5K4DNydk9jE2Ycpgi4XugZzVEN+qTOvKiwMdzUqPkCmdTiyjgefnonLxRy
u5u5ZQveuMCbKBuhiAztLuzJK19niON+fDNnO+i5wX7wMWDZluyiUP6Fz9O0
6OArQe8prSAfTEPFYML6Ppf6qAiZmQXTAcRvaljfhi3tR8VxcmBdr3ppABuz
ZIACJpdDjG1L3Mt7qF+7+TMNWOs2aiZWGYmTuyah/APT3DL3DZU8D1ifsN2L
8gR+4BgUltZmXwVM9QO5cKq4Raj+cqNQkSKmsNKaSWZmNdh+FAWTEzV6Ts3v
A4paDcF80TnAKW4Fw7z8TSyydb7g0cJdJ8J/456jnd/ROfkXUUjLwu3zV0eW
jnawk9tikcTDMQH4Abikq8p897msvEz+J++obfnzbriYVWuI0jNtlgrhZCT/
7x23S4kdqiae3DVa84diF2xp4+PskfFypLJgG1q1+sscJTRfq/h5S4imOVcp
m9byeklGFT0uL26SXRsw5U+qu/PXY9429oVOX/ewEguXCq5VmeWil67D1B9Z
LHoj1DP6Dx1RZ9RJnzdX/FsBWr/5w1Nvom6hlt2OlKpqEwsdJWr9LkjqVkGH
AawK3FX68IGS36XiTw+wMt4+VY4bOn9x3+bUv1ajKl8wzvWUoUkCAqHXNsRs
cBjjO/OLFBKOmtOLryz2r4u3r72UhQfuHMAAbkvqfjKkRvEiXECts70Bg2Hj
0kmI+OVufweJYUQBufivRW/VBo2j8GYTrci6Vg3XfHd/fO+m5MowG4MGewaJ
MXiPJTNPXbU9TRRN/gDq71N2Vr6mC3Xbp75kH7qaAilamw8lchwysb+TZ4IU
egxJ5W/yr2BNesxnH/Rs0az1fb5Mh4+jDEK7BV7Am0bBVDDO5XoqlK8Jssme
1C192yxL9PoE37eN8ZzvVU3cCRhjPtkiyIGPgAnbux0/myPp2UfJoZDrNMBB
8zf09Zf55LdSRNWLwgu6UE/9g1PJGNPBxxctkB6n8dzSAds4fzXv1+UK7i6P
TsgEndkmr3rBHesANCsXEdHMOIQJgGxtS6cLhPZUCTNeTycp9ANohmQs2r+7
r/bz/FDO1AQwRBck+DIJqDSTyqbMU6LAcNo9KW9O5WveUySOdTyEFU5nBuUg
l39s3RLQW0fYUN5GJYQt9MmwKMLhERn2JkC5mFDjXbudnjgfgfQlezZbm+cE
a8nagvisJvu2Fkd3YdWQUDJB+SY/PkTp/KArqfO0nNZB5/0iWwhwJyv6gwUb
4TYedcrL8YpkOGPM/W+MTCB2/n15ZxpPEIraTYASZQsHL+FrLHwpTl24YAB4
Q8V/zfYCHkZ5Vaa0nNWCuuuMUNvX0CS+13opTJYTGRrwtnKioryzoSCMSUHb
BMgcGeKcx+PE176Ia6AqZ92DiEv8oO712oW8+adoRfUuxPrfLg7ezLjf/ycf
GRFoKRyaMuKIwg+Oju1jQLqNOYyFBoOxByZRa8uG656przipxZG4laL8+52j
2Uzb2rx4bkSyiqfADRBhW3fVf6BM2Q4AIBSadIJROvu5c+xyF3xIb8ibRHWs
ICRJcRytUArpkiZi4sf+L0N2I1fqHfE9dQQaHyC/RKQl6/z9QkoYzM8laNf3
n+2I4f21t2rVWyAuw0tg0ZP9mxWZHHJGXJgKbDbelYJ0cc8mCF6i5+Iqr+Uc
25vr0EhrRP/qgiKVC2uibpq1Ns75ZWVTTy6Jid+bfbjnaiUuOvFx7uXZO/09
F4nllTfrP2Urn1DePsvwZDTmaRCvCD8E86NOPFvFBdT+il61ihQg2dnT4uOF
ktJfMD33XmwsW3hDOxXS2dWBGvqjFYMq8r8zoP/snfg9WwwXcSGeygFqAb0o
jCgR73ZKzkd+/hbkHLQMePBF3sV3gsje+DwgST6Fwtd1yAA67mThuX82oM6m
Z9MYmd7STm4RFLvncaDMETU0zmQUZVUSTY5Jq+pZ5l/i2new3Gih06qBTcVc
2qiPT31iAUqmTRbQLxKlepENXWICS6BzSpfQSvqw1jKfDeEeSBJhPeKrUjl/
U1/d3/NABbpGsIHSgVW9KFz1odgvdYGCQYeTLhJLqwKYedjL0HR9XVrcBkEt
u7lMChuNwcz0O/PAj2iu6YwMxsuqpZ9Jl3doLryJUhSuhCGi+kSqfqmoxBJK
6vxTq+ouVEsk9Sq0mVYWj/1J2OI0YkaRmeqdeCc+KNfWHDlv8dkBSbB8bMev
eeqlMBjyS4LhYCXO0zyqUAV/J0B0WbRp6EVcQLkoBTc2KSJZ0iN06rAtMABK
nCWWWhGPn4jqR2OTV3f+k7NCFlEmNcGvbS4PMHiyvZtVx2Ub3QquYYM9xTVz
nHV9L/T2q9WZr4EPFxAE51uiedw3WbMdFvsPWQK5EPAEEAwn8mZaDTc2o7ZX
mTrZ+bZ72Tk+1exBaASgluHm43DdP+3Kuzay/ANmDPDkAtfNmGGLCEKGY85g
rSiA7yzhssekmSH6yIBhToCEF+TlAcrTDDL11tsBVB0b3n7xIZGqt7vBoWXU
5TtUY9eZ8cB3C6qHmnqL9xeRMvgz5V5TgnVZE0Pc0ssr5whs9bXcSeiqjVdZ
CR/sI/nEBOrf1mBgNO1IghHfhFsxjXYZS9R/orDo5gHf5WDv5Uyq64ZLR+ac
bl/jn3HkMsjgP0V/do22KIBUGUsJN1fwhaqGNWCO4OuurcfP/9KWpAAsvW4u
bUzefBUATyRWotzegoeXKbs0tj1fPFWYVlSlfMKyrOPOt0YWjEfFdArgSnOh
JE6UTclkve4j6sA4l/bXfeWdp2/HMU8uxX+LUHVxLp4BD4SN7nZXQ/oNUwoA
oFURC42K00OHruDEuYCl+bwFnIxh9vU9CKz/scyde4isI4rq2uY01smHm/lZ
gOdYQfnK6T40cbLNjrAMzQGM+X38Eb5jdd4HvQFxGDfSovwug+O/JLp7Apu0
TNt3kjtcHZqDDoOyX3kpa1s3nk5PJWV0RRMWulr8p0kFomayJ5vm8hbdD+QS
uGT8plbOoqnoNJbvATVi4/shJVL1Pk3+IjQ2OBZe6Ju40XOO9xKl4/ecqOyd
eVmlWfCA0e26VjnBgMjJyCpoqnG0rFbB4ES6OaurkVgJYOqU6DKzIginysVK
iTii75i5iKzR0nTXBZIRP3tdyREdIn/v1GK0T7f5cXiqtTOfURDE8IQayORj
P9u5+nW0287jBw3101pd7pRt5Y7ZR7FQhh61T8fxFDfn/v5E7DJ/ISNn5mNQ
7uuMirllxDE2dQbrprAGK9ZsfFFhKTmM/Ovy+MusM9bdte3ZRFuWSjobl49/
tNh68ALy6LF6cAHIIydRkiJ2uOUGyE73De4VY5rF3IH5LsTsra1YZopIp6IH
NrZ76S3IlbNG+E0M/fkPFkg5lVmE+iAfi0md3ZcWJd3alPgdHz8RJNo2iW8i
TqbWnJ4JGhC3FbdqBmZxDFcJ9kVQbfSgg797/BHJhlV/EP9hzeZ3Ifq3Pyzp
9BfbAOpp0a5kr/ZpJhG64GiVfwLhWR5WxEu0i6fHUGArS3yzyVmk/j0lPP0g
MZtbFqzokMk/20gNVQZDId+WNVaRq0hX7wd0SD5AyLpE3CxunJG0d2xgyDHh
DGTfLhzMJ1sBE5ZsI29HSGo7KK3W+USAYEm8BIyeOYENfJeKS86juiSnpHkg
KTs6iXUFjSSxTXWAubZ7my6b//rRVZhWSsaaIHxYeQx8pr9F9Mpp5KKKuGAI
OUjALtiW4Bdvp4nUrF6Le0B9+J3R+TpKCNGoeCAqQwbxGylxNuHu0uXDibo6
yZuKVEFagVkVy+VSgAqG2k4oTORurf6w9oCaSUepB9iVMRHH7TJsDwQfrKjc
3aLcEZZ8JbNCDVPwotmLJT23J9+eXsoRMyVHQT9h6P5nFIPfT6/F/e1O6X0p
DhrUFeb8oI0IL5Fnn22Y5V9KYK7dCeAcyZQ1e4MJzRs8dw76/65PBcgOgpCa
5FrqkNGlBmdfLFeIVYiaE+AgfwtxuF+BGLHu6pI33sGX+VsW35+0CBohwHki
R7sMQPCwg04cTAkUyUqPcXxmKZQOCwjr5Fuews2aVMbspWHSKmqfe28M3/LJ
PnRRa+Y7BfUcqlCxlDnEVfqQh+YeIJekr2Z4BOjM0nnK60Wpm8rbO6cm1Sl+
eFZ5LwhQ0DGFqFfJ/uu/YmkXrQrzoW98xyVwfW4IL6DNQzx5+qcj64BSMby3
T/qO9FoMh4K1/lCisie31ZfQs3qdpSF0UdyJUl0pXSLPstbQs1fD4HwlmRte
eFYjzLwkBXgYESGOurcWMIrhVJ9Sgu1zPBWH6XPZoIyHa3lJxCaF1UZPTyye
7SJoR6nzfsH1b22Hb7s3UErqWmVyLamxU69SLsh8DB/xT9dlQZzZfZodejaR
lMwFDbZWyVUd4onPOMxNT4sckstCHa4xjs88qyWwybeeh+JTnHQx4BAUi1rp
h9fzLDAICQNN4OP+cgXjvmL1vygSmfmE5aHX/5r9U0d3TiHmqcAeG0C9qqtP
t6uTZz/CbIQfyW5mDjioFdokbstn9RvIvxa2Hl6q6/0U9/LoxkrZkJffXibe
aDJtRIzPSKLFsejMr/RXdm3h3RQAIZVnRJIEnsDd1Dnz6cmlp7qDO8AHbgY2
OVYRyhVoOAW4O+RbvSdRMDNXHUYzgWoKfQtzfo7K+1qypttRHczAkPmDsJTM
q/Xc9ueAPj9NGIOzJrk0BgpzvwRAp+LyDOOIqkFpwyepJgAguvhWY9G74R4B
Wdj1lbmidSqXAbFkAuhohJdL6rJhYX6zO6Ix+OeTWmvNub8j6v27/YqxeSch
ITMiv75UBNvtRB6u0mdfYBBhXegiaNfcH2PO7Fkr3nBiWEsZXCbf4Dd56Fiz
TLOKlLxfxyfEvn+BEHNCNLO/alKWlVrdD1QCD7njpZzt4GguSR9P0uItFBDm
ZRX6eOSWmkQ9W3zPJ8SaLJClbsRWjCh20MzJtUeeGIE1hxPbiC2/KDhchVw2
W95vPn02/riYDG1NN4csMCuB8dqMZBjkB+/xXzFXwCmh8iBNuu9knJChBKc0
XYOO75Ewv1g7C64JEwtC6HsiQJJWajfH7Ed/FODZiq50GtQZlbK+b8b4NVri
90YTlbpUfV2oZjgWdc772Q24NELtA2GnmhY8zyXjDA6DDcWdrLPDU1p8DRkB
krOTI02yL5QNdFh4RWJ67kjIMlId1MukdbHtly6cz5DP3PyL3Vr0F95dTgqZ
o5E02enA1SZiD4YgYl8cwhLfXHuCaxs602HxgvTW/JRKA8IQ5z+4+ECEKjcj
RkkK9TneK4wHHT6Wug58pr92V5s3zWCM33E8AqP9qH+sVrVyGg9PY8ZYFVB0
fa7HSYcrzphqKvKYLx4wBQbmgmnKgAxFE8hgF9ebcqw0EhzBMGIr6f5vDD92
blpTvpN0YmwJ5pHH6L6Op8zAf6QLZHMMFV3LALa5uxLuj/WZ9U99kJFjWklG
HI7crhPzZ2URAnMFco7hCQvV1pO41yEE5LZQqUCepa6POH6IYW/m5N068akG
QqaBWZs2d0h4GjroHSrFEqcQHG3fIIBlaKpC01PuATEE7GeJgOgsPivJQk9Z
j/VvKwymjNtOsnTzdim96BVghqhDwSYqpuT27wJJnSWIVzti7RRtXGRe+B4B
dwj+ZBpxbKLayR4l5/xb61seTkxfaRQbljXO5o3dmE7dmo9HYMTDgCNSxC/X
sNEQG4Kq/H+jPrNV49IexclGFzU7sJeoEjZo5G2nznB4cDbKiFOjqRbGBRdR
Oav0ssTArwFxadfciqh6ZBOpXjXxbaEt8wcuXsmXp62PfmQTFHYyo4B4uUu2
ziyitFoJIcjhPoyJwTmRzJ0E5e95XI1S7xy9PHRE7/6573VN2XxzV5n09NwH
9dlU88n+qRIqO1sNiDHxUDw91ZQ3trgUUE3B0P3rYdCO73GlWad0jJajx0mf
NCxc0PjmfInbroUpniAU3M0hE4+LWwObnBlQBumnp87wE7VQ79DXRINg1czm
z07OqRGhMQNx97EkPek6XDBQt2LhAzClc8JqX2CeLLPJzzHcuVsgHxRY2uMP
Sm5YLqByrNo8yAzkat8P3Ddue6AoIfrgAnReuZ40+J3Ev3xVh5X0zSEhO5Hd
XXOyvsl2wMUULHy1ZIca8iC3ajUuSrwepE8cf8eib+EUx7hfBXab+O28Y1qp
h20iDdxG07WMwTK0tNW5MRj3bR9ZUDws+L9zNNDVwMU2BEE0AUxc2ht/DTQN
eqzXmlb48RjKqNc2pPVqauI4jkpKMX0XDYy8ytupfVGF3gSHy5XIFGuejIfP
bw9qQK78I5PS6zvQYWWmy7EnkIguVfE/14GR/BJS0SGkE162LzxuHPISXijU
9qKeP6eIdaZ6CpHHrREfyF+UWTgG+/g2g9B9dFWVfy+vuNatGy7jFP1bOFm6
tdWYHtcmRF6b+iF1Ew9Y5nL3FbjC7Is48lRloQK0+08qtCyTyX4VjUnYA/Uc
vwUccEdkc+EQihTFTbNNhER66IC1+LDi5Whc8v8yla0ik5AFcinFdY8F4u5D
Dq8s8ip1n1N3yKvFY9FfCUsonPnxNiwLLyrjZtoQUwm42Q2/8bkxjapokw8t
ygAG+Y5QRXXZm5piC9kOFN7EOMVtCtHjviFgu9WQICoRDiW3IfS806xPKwKL
MqnlToDlv0/DDu/CUidxcyl8+wxIKp8ePHTDNpmdZwmJuTRc5+4/FulI8IuV
rCg3VWKMfy0H5kinZ25bfUc8Bn1yiDi3CTWUaly7pk9Bono9UOZbeaalfzFg
Kd0ZjIz5PynY8SIrWR0+eD+N3sjPiNb8RR9vBklyxx5+qH2S9l5CKiGv+O2O
AdLhZixd3+xKx13hGIEqWckTBHfpb0qv1aRSsT+W6Fe2WXe15p4FfnMh0aCH
pFV2CKntzCxi9cK3aP+GfV7Dpm5/z2aVgJrt9+3D0GZoAmbycY6MG+1FohGF
M7sUDqFMGPJyxgvQmgAPDhRKONkYdq4OIJKaW9QyLQf/ZPFbRTo46XYUgddr
Nn/zSRZgSUnUnetGr++3jPOXFXlVmDv9V04QBOaQZbFQHBq71dYWOtkyCEvP
Yrhd4vpu/T9Tz+hYvm00YA2FgHV3d2CSv8QEta3OTFDuELJD/TL0epJpivmV
8NGCWhSM/KB2LnyqPcz7tyAsK2zV4DM1eqNGHUdXY3xiJmqQdGM4PRgiyhY9
IpSt4Qv/4LOVYFWYD3G/fUdJBi/0MhtthPImgah86abc+tRS+y7PgiQEmHec
x/Tim9VhkX6BnhzRtvepRj269op8jQ35Ye1c88LQRcOKs7EdY/Et2S4Qab9h
8WvCHqYUzO3GnJVkbsr/6MTE8omgY5JM9xg02/k2JirBFyt4dwqSK27I6b0g
s3pOoe05T4QqIP+lokeE6GL7Xb0QSyTar7xhG8V7YsEZL/L/6TcFmnQMMk67
oJahE8+yr0khfrNH1ZaZUxf2/17yJLf0hh13mW3Rht+TBE9imwzqhVGA2fFw
F6pLg9zxH6Fxw+Ya6S5EAZKALhB4yVJ+sdSQSaOLh8z5e16Y9JFdnH4opuli
/l0qkIqxwnOtvs+8iDq+5vjkXA/wrMlwPZzMXc41JkcmAbYo5+cCri24lVWt
XC8lynSwOH64QGGDAqORvdPAcvKREbuGfaM8Qk5Jlx+8TrMFhjHqOiV7OEtp
g9N+gT2TQrhpvrHWm85fsNpz/vZ2xU94m7YaB4qioNQcffUQwRlb4ynujDEC
jm3GwPdRfxlGPDaAfOIg/8qn1KPN4ZZfgDajuqCFtK5T+u/ijlATeV73Z25R
GFG6PPwt/MR5bN6GkAZQ/pJ81HNJZavGhwSzaMIKNI3HWqGX15CANMEAST3e
og+QMcv2PibBuvlHhzcAGIfDeRHbrAarcym8h+Y9LxEFyO7yOW6jPNnC/XcP
1A8cWjmkxrvBAQeMFnrK0S5PE+57GqGi0xYWp/OnhxPciVSxkmPAKuY8J44d
f2HjKTmVUkvIdgvdy7EyhKOSnN8bUZyyMj3hQqWjgszACm5rGJUsc2LTVCc7
ANSleIRhj86h9hEHSKHzo6UpRzo+rE0VZlAUa0pcWYe06tBuY45Mugy+Sc1g
xOaxSUdSxEjxiaAszPid//h+E9Z/3YwAjr2dlkIgA8Eke4N6Pi5bxFUgvuGo
Cn4l09bX1g8x4FFfZq0uLJeO6sBQswVBPABD5VyxMfWKHqWmq+1+0smKp+yj
kcBDn4dhotBtOb1JcLitTNmzTbW56kg7/IG2nngCbh5EVPQLmqnQgk7FauNu
5JKvYVMc53lgHAPrn2rx6usIJZQQA4RwaIUvUnitvU494OKWkusr0HQhM6Jr
n2fsuGgVBVs6jQAZRnleTvpfO+KyIdPPPUGgGQXYdM2V8db+dxT3nxs6ty4C
aS6MWpX2IBvN1rwx0VMJAAn0FmxvsI1E72YlpvlMzf8vFb9tbS7j4lEzD1p7
X99j0+/WepYnn+4II8NpJo1Ix78YkResEXSa/Fd3xhjeEekt+i/xkXidChnB
a0BroC63xJZoMk8EgJA/xSUbQGb7nMCWqib28aonETt7OOtQMkZauopbOXlJ
EnxyPCdPVvyC7LCQ4BLzbANbWyq9LzDz9VY+VCA91KQj9iJzXs/VPPrNK6Yz
ocvY2oXQg5Qx08uTvhRTELEKfchL3dUP1Of/k6Hh5/dBHDsGg2j5CzcQEWAJ
14JWUVHQNk6TgNt+ADX1rb4SDIcSVTuwIrR9nnqwEgz3SJ0mLTILVvJ/4PRQ
EQv3wXgItjoHVUI/i2ZZJ5m8+baPsatmT4q+r9sOmLu8BZwIwTnRbS5AQ8bH
jSNktsMgmGM4HvjyMjtNsf4PgvKIJVRxUoKX+0xaoZAOuTbBZxq0scMajcPW
pstn8NpZdFeCci1WV+3zfgHuvZo5e2i6BbR7A8e7LciJCGHkd67n/bZwpU0g
1DTq3wgkywAAUYP0KNgGEzx1b1aHWvDlgfCB8ngTiREkX6afvzWzfXSplEMP
ircNm0I6uYP8ng0WzTUSgJwLwTRLV6BVL7VY9/AoH2vjnrsLvRUT6XA5IcKh
O15q0ouVYjus9IjTDg55YsCzprv2l2fJPjBRHWb+nmATGTWCuIVCXkxXLGCG
i0ebsssxU6LwCPn3C/4lApMwUwVBtFoSvNaVYBGIcWSc21U37gsP5XHoUC/f
1cR3wStGmcDNrm0VoFsuJg5O0umEQ6hyqFjf1C4Zd0hrIn7tZV0aKPLLuay6
6CdgaFVMIZHgUD/rQyOO+R6KQRWfuRdmasf11UJYV7p4wet06OgmghFJFCii
R3wdy6bKxeoYvMp3TZIf/wvmrDYPn602swrjBZ4o39dJ3rao5UeA6PM270Rq
+qvZL/E4XWiQ1eEY5rTbfB6f1JcnSJUpHCuGjDQAHZNiLRJCguIQ+lvROvON
LP9ChbWtcrDmi9dkpJeVYhscxYuIi7OIUxmyfOc6BHQYgS5GmDA3+PDQdEaI
rJ/6DLoBRaaPsLsMQWOQ0zuQVLQ4qSkfNH6uKSJeZAw5CDJeVH8Suey4CsfW
UWIUVjV3nKlSrWG/ikk+dm7ZAIGfxAv4vZ+NsOOJi/NUEcPhVcErAJwtcjru
wJTje0AiKBMmwyiDDXCsYQPBpRuu8XOQG4tpnxPXPDcmfFfLJWGuewr7BzSg
FUbMnqiKgmUFqFLdcEBg3FGRfTysGbF1RvmWgWQJd2ewsT5KvLB6zxJNrtAy
Yx2loFI364Io4VmtfoUYuOvXEB6qFVZSVPg2W8i1UIOPRttA5zNKfC2doDLg
cQAxhjPrKbzdoxZrBuBsp9tL/K0ZfMxJZV13zVAUjD/UImslJ8m4gxl/kQ17
kYFedMuO20zvyauSN8DsPrQKHleNkghJ/rOJBdJN8J0uvUedwXSx2nlKa58+
V/NrhFJvuq4LJH81XXiMZMERdXZPiKRvHWJdM24L76BJr9gVcrNF8Vuvsi3I
uAUzTITe0bfQf4bBtfMoMSaSpBp5iHzO7ovg0u+rtdaIAF2PTE81rvpdk5nv
CoPPIrpRSTbffwvUYeAylfTuw31mYdbHGLccyHJVo0ca87F/K6/XfgYZ1RsL
CMJ85Wd0CKrViajMMQRbG/CsVB1FkPEEDwhi9LnURrHD7Ofte/ZbP9RdLFGz
TEWbNwgXlpIW9hJiUpZlN/TBhCkKojdE7Aka9XBx3XSPWb1QNrb0u4/Q5j4x
55OjrTe2VHN0i9HtlA5KFzrwhUr8yyucPO4oYT5KxYvzAHIX1lhZ1QoD2iLh
uSkL7MghiELNZb4N/Ouq32PyDLbbvkm7S0exkhyIiZSXCxkv7Wzy/hHzAwrI
MtDMLtcorAAMN9BZKpDeyKLTgFVTTrMg7zRt+rI5x1e9mWKVb63hiIcEK9yS
zIGIYGv+6HFN4t6IkFRT3vNXozR/s/k0M4Hpk9k/nLsKX5FlIV/Wo+sOsmMj
Yzxt7Jy1+oIgs1DIwPkW9LT7qfUabm1vpC2rKwbMZAXHSAaVFvKdfqxrYvRO
Lf0UVdPETQBaMFVRING77zYQjPtvuxbDflAdUqdzHOAB8gMH/pw1oeD75fDS
ycT2P6GfOO7hDODfP9zt8RVZyIUPGk5tTu894GpiUTA8ATUwgzA4uqiCdTmp
J9hcQlGVKfcJdfGwzd+f+FsXp16vUzGqvJlaZ4sDHV+JBujfYdKw0u/i3ht6
lNKTQKcVbMN7xJBlfnE3OwvapH3zdPyORpyCxm+oCFsuoaL4iZOeKrq/9O2Q
sd5J05i0e2wjaA5vM4pbxWdbw0RsyHxYmejz6OI8Ivp29Yybt2/yqTpIb1MA
r4FBpCgc57eoIB8ThqRLmte5na9tnQC6sVqmDrKqT3a00Il/+G3WHSjNaerp
f62tNTOZ6+Z5oZJGg/UV2bTy1S7BaiuGAOmAArupW65atbRjyo1IWj3TIoRl
54GtN3U4Pj8yYd15BgNCnxO5brcnPlDIuJVjzELzJuFpqjeocFx0fkHhPl28
j1ycwvVwRwC02GwLJRt9fmrTXqFCDoWiWX3dg2PzJMT3oVUDQBhYmivbnTMX
KsXhM7A4/ed9YqVpN1WW5wWy/7cwbcwHcrZBzburoJL2xFGP6lPGAkPZgcib
4pTHV1dPxabge9jZ/rtsTjpSGz5E7s1RWAs+S+mLreC9v8dUf/WNNl7OxtVG
EI2XO8ui13wirVfBJJWFosrATig3OldDibvv7MWGz56IB0+iXu+zSsiFcXwo
aDfuxjDa5jOglDnlKHWKQNssA3nFoiRCaPSWb/hQSUm/z9mJdklNZzjp+kpU
bfaP9qn9tz8qWCjTuGq8fXMkwl8MaHQ3atlrwUe+8Ty+ZsvcsoSnn1O5rU8C
/+lb/9ZgdS4FtLo73VFZ25fS206tcp4NaM4ZeL3maJKuEAdeMQq3JMdHEb5j
T5PPGXO09FjlGtPmSmgJGxrizNZvVjrBSCSj4b2r5l/n/LMeTE9JPHp9f7J+
Li6vtzpHcjwUzP7shlwLN1nlpA9PNZPeZyG4kcdbiXngcPn09z6XR++CrYI/
tOKzAMMguC0HEaOmpbagcqxTjZBeB0QCtsdCrRb/8/FgsIicU3NABBxhimhj
I3WyEvmRoWOb8hY+keolFHDLAHutKMd7LjkAGRNc7k3rY5EhrFGCRUrGgD4O
gmQV3FvQdIwxyTbqk9FMeKbsCm9MsVlN9PcRztRpMPbiTfNZ6sjZs+WLopbx
f+o97h8tOYuvDZCjUaK8+BGXrzIQEptYrJ9lDoMYiOluwFcysWJUe2bPO2jS
ehdeT2OdkJpiXlfy957pfORbCZeVoTevZOcOh510Yx95nf34o+s/rE7xRJI4
om55gFfeXBHjbXyn1efXYug7W2WTEyqfShKZkv95avBAb/acHnSDyFppnpmE
60XIDgayqKalapu3UaOtCjXM8gQL9947HmQ9Maw7bCNJW8Q//1LrL3bTzYs3
t82Hivz4PP+ke0/c9H1LiyUb1xzh9KGHzl8JtkxRbbWtG3ZmnEuk4VxoMZAV
/ksVeYukmoVePOSQrvxrvNyVC6vs7KckhNOj1VRTdzHmn/JRgGTnQdn6lStf
gM17NKJMw3WgckoWSAGXNiIBXX1CKnRL8MhYw5XPv3L7G4ScvZbJFKGHxwQ4
37WWeB18uNc2zvEe9g6oQMBHLHjUrxyKdu18Tt6h/lYAHFrn3QhezfAc8eJO
xE7IliwM5sA5kieC7ilo7ZSfTLvOi75VMoWlzleD6v5fjiRs2Au8iAflha8F
xQuq/M5CKRoys2piY4FZbbdGi7hIje9EGToHcmgl8VL5gtJd3lMiLBxIjJ+w
puWGzJ6csg6/RdcuSXNY+ZsPwyTdNhWwUOLfEqD9zaMkaBlg0D41kedt6HPC
lGZjUfePQwzmNuj1Ezw7TitYMhLH25SYnnHuVzyTMkHDqsQyTiuRgcuJE/PI
NI8pGQtwUOPrRWj6q6GzdUrVywNnW5Ih8cdRt7+BgAypgWfhqwQ25/7hYapZ
rgYQc1ipwAXDZ1fmLdtIFlt+j5ysl6NZLJwUcvuh6iIlWdEft7vtC02tPAB6
AEItYNVTCHSfNJV5MxCWoJEOQJx2sDwdGC1bWJRQEY5UZJsUhFWu4S8bPYi3
TcNEQikNH1sxioKgxkg/3n+4mF5GQaoHGNMRopT+c6wlkMCKsrNPse1J8fE3
aQS90NaUOmnYhCCl4vDjfD/EZF8pIVP4cSyQiVzs2WYoelMT0axBVNvJmkEP
8/4cd4uVJ5ppxNxvmq19AkEa8kFE5VVxWq6+NH3zmRmbXzAgzpak4EmX5Xv0
8doO8Fikl03SVILDty+/gs8tKQc5Ua3hAAGw2J6ThbBA2LBkbsE4K67QGmQx
TOWovXbPTW5byXU3y8j1Tj9Ivuo7aAJFlm/SUYZa/tsz0ETXHCU1her9Xm5f
Kljr+id8OtuAVrxF9+qu3Eh6LeZ3sLGl9BgLT6l9wERtTOk0YbL+BDkV4iRR
6lfeOtv2oSBewNmn4omZOAKQz51DYaqCKGQelJbAtil2D5V6Bo020Gko/xAE
n71FuzShKxuGFCv4bP/BJsxpFXloUz8wbwqZs4/yzNoRk9gqzN2X9fq/Ye+q
7PMZDPasly6OcUNDG5dQTlp9XVgM0EVdHmEF10lV/L8YD5r0mCuCBraENiPk
XN1ZbpSTzJSOGrfgwOc/YJKDleZka2L+U7oyLIuOvPvu7B/0TE4s92O9eFEz
WdiAVGGbI8OJyDQlpETBD0BCQFrdp0OardPe9IrOrv1FbwdRLCNPTTTYZCEY
bVa97ImCrKRJOPilPvOZ1J9P9voSC5vmqy6Pl1JM2BMDFwrFHRP0d92aFW1K
+hZ8LzstzQGz+3znbL/Rp2QOWY0eP2LwawbrMjLU2T/gLd6nC2+rvTUY+qAG
4aOV4VZTirkS+4RpKoQ/m2ET8Zup3RBslV8KlEWvrmwG055iMHI5Lp72VDB1
eV3jd/wn1tYiEJObyhD1PrptlSh8fZdNdELXhK26dJzndWBxC6Sp6468tzr3
Z3CctZuyRkNKFkFKVajzJx4cdjaujD1Ji0tcFwWdYEPRTMmJK/79wVG/AgU+
emn2v0kRhIEKJG7MB9V5MitkqdH8LY6bW2rPJG2LM4oUIMc13JtI2LRYH8N8
7QFM1AkSVgrdn12Rys2CClbIefIiWrJXxzYzuEfAc5bhI20iprP89mxsVE0Z
K3uT9zgtEQNgf/1qFqCNTCiCCMk9Ae0FUvD55GXb+yMTnmBJZDXZCd04/QxO
5d3owmtZdOV+6Qu24LegbmvwFH10+fHaJegH9b+bovs80QtEVjMt6Ht/Lyx/
NJ5R9UrQv6zLBGjoYNdBQHjrhThudbFvlxSyJiVu5V5JO2K/rXpHGZcMQfps
yk9Vrw0ZAsIKpkdQW8UlpfSkEW6GOXI1QZm9KKe34g9mKS1XvWJT/SD3DFCa
YHCIUbJlflv8lRVySXzISQl+XBtcvCPLdjHz5u44sAtXBZSOi6ogQuQQEBgM
GpvHZdMu4bSddncoIraVQqKBK8cdB7hWtvHrLfAae6iJrFgVuRSKN1qEsquQ
nI6+EGKy0AEiG9ezZjzBMhc61fLqQfF+RIQBn/6RAWptiJE2L7XjtmuMe8HY
wIfEKeWHAt3JnrKiVkp3ICs97yHws5zNGsBTukeqcLK5KPmOsckRLZsIzvuI
rRElSrjP6cDRdLYK8c1E9hrrB23fc53CcJa/MWBPFfQ/4Ip0h2K6lA3BGs+O
bg+lVe6gNRUR1RaPLjawi9X9WqiB85K8PyJvPLT9+ISBa6SeesR013EDvjOt
MRpxFtOj5OTIXpJ2ebf8NHIbNRMzyi71UvJCkx2V5+PSE6xKAgfc7gZ3ag+w
juhFe8StH14AUNZ9j3423nVbTW4o3y1nDxxalmcLKevxM7Gv9K+t9EnlMltb
WuvhuXk66e6BX+AX65sexl/bNYk3esybur701rL//xeqHN8IoOoJQ4v/7kBo
mKd1jAUWnJLQAYFFas407czKjuzXn7hyyj4Mwb2MrvPcHX9fbgPygfNbo8BZ
k7JQcL+r6O7VpEzZRElnpc6VK8MwNELZTrRsHhX9m2IHMREcMYY9NYVzCUSR
DGHEXaBj4saVC6Ama2Sv3ULG3NH1+SR+XfAkp1bDSPD5T3HKgCHbPLBLFhwi
wIUDQo+xlUcm8ubLgAn5zzNVNg0Ex7dALS53T02tEeVDaQDbz9HsvwkpKGSk
mwdKyEw9ha+3L/lvZs6y5KagZm2BSIo5mkGe0p8NSQWBlRRPOYjX9qzpJJGe
s1HypvYgSRhFucbclfyAcfEPi9S4Zq80Yh8A9eMHEXLngfsjh+W4R6p5FvUO
Rkb/iASQsm2rqadIrEgOfhkamBmd8JiAS2hQDpgBGjYj/N0IRq7XQTPLA46M
pBRbl5JZ5iBfyEuu0s2MWGYWShPdVqG3+yjg7xG/VhPghx/TNCOw7TL3rBZz
I3LuaW59kN9d4WT/sR+2l9OVQtPK4gWwYj/faT5MSgucgutcInbGwG62/HbX
lEAw9DmEhYTW6vqhyssMmofF4E8brUCcLNs4mV9nYsOeF5gNUr7zSNpjRKI2
smX7tM4X/pibPvDF3sZ5Be7ICbnAoCgQcgBZG+1Zt84ZAZpKkN/4dWg/Xg3y
ugoGPI5vQpm4K6CqLlCtbEt/+X8qq7zgeuk3UoVOYPljTVSIsUNk/7elHHV8
mAZDeN2Xftw2IH2O4gNgkxX2jml5RXTmPm5qeLUgaFP0XYz6dk6WjGnM2I0h
Tf5fdTof3Y4DbXye3yEHbkrRF6a/RRoovMOjJAFI4NfG5DAuy+iUTLOBR2zm
w0aG91HizLe6NqxiOXFHi5Pg3qk7zWe9ODIq4iotpnJqSLm4U61c2OJnBLhj
xvogvVZxeqJIWTfj/iu8KFIm+7rYn3FsCsq506uSEZnxfYtt9wb6JcIHORdb
tu8yxW4rtmf9ViBWiXd9YHXNpKbK9ewhlyWypaTnUmPzKzDHM13NB0pYZUFV
aPXbAQPpVc/JhpjdICQZ62+N69sMxQOU88UxOaMeYyjdRsAsFhmNe/L6YJ9l
L1HEnDeb3m315MGv29D1xKPKINdt1MSycyChfC/VpBe5ed1Bm+2oo1ROFBID
VLfrj00iKWGLrFIe8O+c/jCHYaPF92bzguzF6eYXEAEzNVotYQ0SdMZTxICZ
SsPBxAMdg4iUd+PFV9ZJh1L2DwKbzGncqVv54mMCkEmSCV6chQ4fw7aQGLWW
IOclO6ZLQgEfy4M786FGLSHNrTOQj7NvBTinaD2T+Cv6yaeQekHx9/LeTwVS
LHl4+pGYlLthLMwTMH+7qr85bhkW2pNYmEm6oxBQf9UJ5miKEIcT8MZkjZh9
g7jb2SQl8nPTH3UoPWzNYDUXMN17grhB7S3nPZE6ClE6sNLWvNHqy4gHNHu1
WAmUyauo6VZwcYXUXdyLoKOSCjyZNtdGE4C/AQdzaR7O8ZSenoUPkgoLRp8j
ZvVJVD/fr6sTuyj8Fwvgxvoxw6hWLXOYuQfSgZ6ZOgHznZaITjCXDsYfa2xp
JIZU78lhBDYO6J24F2dNVeZ5wPr7MnH/3/FCt9ZMJRi9yE2FSYWKdhz6VLKm
ZX8TczW2loav7cAgkouT/ttW/+t1TTT1923b/lhmUWgNmcQyoI/axpcL1J4N
A5gTmu5+nwxaQSKjOZ7h1BRgWSwXpbr0f2Lj8BYMIxtyo19Bjyezywcz+tIP
x41dcPRRZGxOJRAaDei5+8EgMuSwE4neiBKWfmOoW9nvEKMPmU/yHihmFs6d
nl5d1Baarl2SWkmNOhfLmqX00KKNq/WFqqX7CRVW2ZozEtPhZC1++uTl5SNb
Ty7kSFwnfCKJ8xM/j9DitvEao66Ov9KaT5cXqCyq0xzHqQXol5GjL0fDKM0a
WEvfG+p0wD+TgWDzEqW8/UoG2eyMRIgWSOyid8Pf+FbtUKVH4SbcZEm1WLuX
UNHpDBHzbOC2yGDTmdSlZ6Xn+AVJY39JofsThaJyMmSy9xZwUoItGJSVSd9j
x0vZmXxCAwdZwWGtTRBcay4tcwHMC1zR8+UA0YJ4Gc8dsHCaXHzKzyosHqYY
YYzuONHbFHAvvTUXbGJE4oSVrZnan7m93OmRAI0kZAiVvea+0MYfT2Vba+I8
sKTkTZebO8SdXCNhgzcAyTUSDVeKqfxB0kqZ6MvWVPKV+SmsS3AzCBoEuN6t
vkftd5L08X7IKe9bYfnF5vZTTaUzfyFvaZCODg23K8qIBgFcmK2HRhuXqxll
CtpDwKVwQfEUTKwzn0KQcTvYHh/HibvmVZcfhYk8qU9sVYABUVGasfyxusP7
5MoY4nRU3C5jkqHNoLOneuq32Sah3u3ihpQVQcj9kOQuEdo0CvOSkhaBy894
HljUKhek0eVyVtz+E8exRjx3dXmGH6kt1zoCmHi+l/Dy/jE4SEYFV2XFR4Ak
RFeizsktbInhCYQ1o6WTepGcBUHCKZ5EGrF179S3pe+Ut+WHc/+Zr0cJJqL1
6q+x+aZylCFbob279cr4Vdh7UFhnMRL2lUoezcgCVqI6T/fU5+1Lcz9gfe4a
SyE7YwnxLstP0VIaABnQdQ3IA7HdD5IEQ4qj4r5rjM/JzjmiRVsv9DUHe/0e
JIAPTl7DQSrOJK+ewCOQ/IyaMNgDLoVBHHiFeKIG9XPLhJOwbzvIzK8Y7lfe
mSul0qQmOjA9K6p6D77Qwc/AJE4Ml8NeMZWjWFG5LBj5JtDvmXfA4JeSSB+Q
VjQFb4Hy8FJz8R4a1LjEOxkV4JlWewJHaB0r2rrdtpomJYYyPsnvOPJI8lJf
qHRoZFVn8a2Mg8ekAt0Lp/4z7UaWzFnQ3C7hwCqiX9723IfQ222IBo+oK+Kh
NOGh2+UKMtMFaprhWgp9Uopbh9sZe9oMKomAc1Q/mpXNx86Nt8pKoZrYwXDR
GS1bMXYn36tpxtOGkIJpim/R8L0HvsfbFa9FFP5ux/lhcFke7kHpbLyVIx6M
m3yClaPEKf1jI/reDzobEYi9EpIHaKLra95CamNUIHaIDUDbIW8uLZkTSQ9H
xzergp51n24JDIg9PsyedgEIbSPTIB6Pl4JGak0LIf0pouX8AXx0+nj/C1bp
N6HprVPOwEHr6xHE2M3Rtv9pGWKefw8QE5FhU+97NxiJzvZAPi7Nvb7FGSfb
XPrEuEfhkeUBV/lRlhIXxm8pOzFKXZvNmY7RuBAim0ya2J7gDAI4kMXmgY1N
kIW2CYc7UOkVaOXeHOIIXmF8G8Smy9KXWEWlVbMo1fAAeh44qSgZHBZxuQdm
6yAkRdSvChjUUNtoICcB7uYtNCYI6Y4Ys3ZU8ODdvD8pmxRQHPVPlLO63ExJ
26SLeGjG+p/c57fRkjBR8fNzcEqBPtj2kqvxpY1sPwa1wqZcoJIK5/W/bBkg
khXB4cpnrYsgW5bg8tb+UdxaV15K7SY9xQER2dQjebLx/auWBuVozx2K18wu
jqnSuf0O2BJlSUR6sNZ8RbwRw/9Y7WZJcQxqpsKE9012hpvf8CaaYs5DMkaa
tOs9Zfm9xhv8bb2ayvviD7hvPGmOGW1JtrB1nq0pn8OCOk/zxJZbDpJJTe4L
ramx9tXfpPTeK+LvbvfsKEuRj7t9PIGJ/3SUaHjcwL2qTRiZJiXClqUKN+kv
3L1CfJGwnVX8V0AQzOcvXfT3KDzdO8Syj2nsjBwowaRg8ucvzr2MOZ+2UQnP
pNk6r9lLdYoCJRLgz9OTAQTDPkykH/pPr2TNLJh70+M4O1hgo88lt/fIA1l3
GLCMomtldpzq0xQ593r+JUXepQYsyOIJxtWNq+5Tcv2oImPHmKvCXqPOquJX
qnRxDfqpsONxRI0h/FY95HG99SF9LgsJrf2uZ2qROi/G5DVobKgccAr7Pewe
+KeYfdQr8wxvyisubuYQ9NBMm9fqaekBK2RUdxloJu452TPcj8dF7zOMoQWG
K55oRVxMXkSUemgM4GnblS4L33I4FzcnGSyAPyxajJlwn1C9wvrAFomK/KcI
1gAQ6JGSp5l8nAvnVE+3+KUYMq0iytcw1II+bQBJ2HzDJXfPoDtup3wtcxtu
vyRUXpYsD0KojaAlvns2mSy9fHYR//CeC/ednQ6LlvppBX1/5rRqXQr2ue9m
DeQ52hnKzJLpaPX7zttzFkyth8BAJde9KZyHeAIddRioV8Y6F4qdHpdmrLE7
rK6sL8tVfoifi9o6IuqyxtM97H3t/pimWxojcOCv6RqU6g3bKTiEOLOVqPEu
yHLLVi5E34aSHPmmx3WuC8lM8nS5sZuDN2zgbPNBx5L/J4i55KIvOrATg10m
yGWIOnR+GQDBFf0l3WfKhKkXK0ZLuheoyJr2YmVMYU1UeYfCTbbQHSCiQFkM
Qp6LtBTzb43ZeQbTKT8tObXdfsmgo2Y6XvDfn3S9weIZ0toR8RpPrpXccZtq
6UAgO5aGwgbM4zw/xxxLvefHumVij564bRw43kn3uNGZAl2BQ02IdNipKpS0
AeoK6BAMCR7uPWIHNlI6kVVhBWHJv1LYtJ/fpRqYxYQNB73TnLfeMtQG+Au5
lQVxPvnL5Fcf5l4KEEj9VrQD7az6LmH8gwXaePYz42BoIqL/zsjQQIa8QPQ+
aVynVKW2ha34e1uyca/kIf0gPyw8yyQoHqas9PmvlDatAZU3+1CYHDb9JqH/
E9Jq/UpDwki8epETT7xx550iRKwaHLBRd2htn3FxL8Ihn0rZ7jKtG0RsOU72
dHiooyubOwyydncd7uKWtjR/naUAB+xWi+32gMZX5D3ZZ8nAxTSGFVs2VEKX
irA2domHGhvRVNzOugTvuAPpg4Jk4pYeM9otU8D9GV6IktOkGYK6Bn4js4yS
neFDGV8xvjHYeqn/31p0kORzhyhIurH5xof0os1qajAfjnTetKVryyOX7qTf
SK0iimkdDTkG9WQ7IZ1X/hbdSaeFW+tjt4DWluTvNwtyegoFaBQzEkkvIa8Z
OROZ9QpWE71v3PYLSIQxlZwJwSwocyESN13Xx1ehGnM9wVVaEKgNw7qEtV4r
6Yf/ogGKzX+0jYeY4thUl90gTgkc/3mqumvvJV0hr2JOq/KeyxYwUJySyh50
AZDJNrT8PoHKehH3Ab1GYQZQNptRkbosV7cocjP4pwTDwqoyxqy0Ld+xwyJ5
u2Di5ZuspKoYLCzXRVOp7en22zyl+dYBDU7oihub7ujaEa3exVRpBtoPHZ1u
rkVol2DChe0BbFhqGhJLSW06dOWz2lIkCgvo0HBDYYY2gh37peCYw0am5IhZ
dJ6j4wfHPIk7YpbD4o/7yxSH24QgKQlTsAkhXrQ3S00De/AIDHxg56edgc6X
ROzTY9Z/90LYM9crxjuyU2Qop563si6B9fXD3JjjrG+SwTQXK3O/nHKIPEYB
7LMeMX0En+wxGmmIEELd1n/qwo1xaKbWVboGh+Vt8+obE38PXnTqFPHOB0/y
7zUcEoEA/5qHcQxyyPb0tpijjCjiiOuGSNdVHuBSXEPKJ2wcjJXRNfLrd0hh
Do09mVYTKjcdZ1k437BV0Z50NXf96GvaznFAmnjSrjM38DreKxlObNRLSK4u
GSbUbLwFngHvoq4/dnQFKHCBpjJrBpQq7u8PzMFfd0zBoqgv0szfl7R90Kt3
1Uc73g0VDsozN44nbIvH8V09fWOODwmyrudCEPGA48AoUz0o1anxS1H/jhDZ
E+Xbp/kH44QclBFiQ05OGgMdK7OfHAJGTT/K3DsIbRekm2pEJdCK+p9ERogD
bhK3nJwapE0GRHBuOHnFFgzI7vJbovXIqvw3CK2Wu774WWQm1dk/gBjTGI0F
lAE4PRwxAMGE2hjF/GJGUkgDulUHQ8r+RKmOaJqq1OSSIUbt8LjNxFpHZFTT
oShftQqzL3Sk4BPuV1t3IRLcxjc87FBgQrHhrN+wMVacvuyIBMY9OQ3wcUOT
0XxixJRgjYyZieV7VukCgeJOhNBYrSN9KAhBYJkEyKRwgJZkexOha2e3sbu0
kV89RC53w/1sFwMtuAm69eeK45Ry8FQqT7gaQlrX7Ybegz3vbe0qP3KUekua
mT6qUUrL0AV/tQ0hiP0nE3agKnCuDLVNMHvS7kQdRKW4zMFZqwMr4B7JDX8X
OHL6iVRvzzRbYaiGOIv0M8KWTvyhTmFbk6W+9jZg8E1sjk/b915yIfe2wldR
VItPLopy2s0pHMv6aGLBwxJN+OwNTVWSSDJlC9Bbx81FPae7K+xHVgB+i1PN
MDd1WZecBMx0esjVEqQAh9WAmEi2/7lkrKkfns2Sks/o78aGTrWmZz+dND44
v1adWjTn2WVKdbj65saoGdvaHfLtrvfVyy/uMcyGMNCpAshxNoEV/y8rhCbR
GY7ccW5nP2XsVk4X5XQBFny6cd07FPF646giqxWuruoHBmfPJpu6WxxstSYK
miRmcXz7A102i2D4VN8xoGjBcDib/lnMfDc4SaHyc4ZgmwmAZhRKQ5WzbQ6f
ObIPyR6gRlFLzToOAF0rzQ6g2KXCxoWgtxgsw6mXgyOl1KZP21bdIdcXyMaL
t6Xd/eG3W/3BnAULDVdtzUJJa7TiwiMVTAwcgd2WG7zN1MwT7gO9QD1f2LeZ
5Z8nsaKlUh5GIvImEdQYlhCMJn3qYroaO0t9nlJO9QW+BJks8+XLacaw1Ir0
0pWkL3JBjLLpy2N6A+VLbdQwtQSGI6DANswQstosbMmxO5dIIkTodIQcdAxz
dT+QRCJktjn2HXNEj5HVjg4Lzn4+BUDmw3ameBd8bquLWbORtBKfCHAKJegt
viyExjzLyeAVieF8XYu6uPXG6WqcjPI2YyPE5niMmn1JnI5t2b82JIzJd0fJ
Hr0PUHCxb8y9ppBt1cwrMKagPZxx+eD4Atj46opW8jmVfR/hd2zrgfKSxTiL
MsZDtI24o3cLKI4jqI0BuRvjgVg8T1sxIhR7R+7tkK1MGrjNpOKP+zXFn312
2Y1Vj3GZLNrKx/uNaG7sjIaGeRyJVjIPqHugJmUJDMV6jS2GL2WlRgmB5rr0
eBMedv3hhOtdeHh5z4dQSw4eRkf1iHao/i/3UE+Rtm5FwLBBGQttvACF7Qi2
SncM2xp7P29PB6UTM/+IiJ34A76k7uPn7TRPj/aljWu0orzwKoCf8377xvfM
jJyiA/AfKQmo8kd4kao0MsPcmGchJ6Kis025LA/j4IwSy/YIIrsmqaw7DR2K
nWI7VGiPeeOCVFzJmCHtLd+D8/5QhTOG/eSfgCx6osiFcm6qL9fJoICYMSzj
Wo6GStDgef3s8FzWayyt7SRrM/EvrRsjAVEbXR6kdSeRYysm3XnE03TcppiH
bHoE3DX9nmrLYxhjHkK2MsPbI6Bqx5XhSR5wF9k9d4+L3rseT3r4LzXcLHd+
KBn//xp1adl2ZB2ki3FiDAuZ+FD+5jx6FFGZlU3XkMCienrJgt9zCd05eMwW
YGKTaQ55/W/28WwY04g8gPvzANNvhODydWuWte6ljBYJ+SIL+yM8wArnVe8Q
sULGbuJJNPWnixfN7WF/lQzHC8OeXQQ1vJKuxaIqDn3X+DyozSm1rjL30oj6
Ly34wXmWlTROjvjPP3joN8tSh3RsGu80sHu/4v5iDLpXhWAIGA9zr6D3lY2V
cyX7OZtwOt2rRosl8nC3hOXAiqkQf7foAu1RkHJ8m0PiXvMCa5msOmYGGfhx
o3dGvyrmMOnHnszkuO4BwzlF5oQ1KZoVrZP0fBamGw2woyTLAfV1ARLjSMnM
hdgPb0ht2fsJu7XgZcUUQO5SomkSPP/nhZyCurQkEcZvEkyWYts/+B5EF0cR
c8jysG1DIZ3wVkTUPaeBOuJsBBrkUwW8+CriYYgR8wCbwBfq6hjdHVAB1BLF
WrK+MGzc8ob1b2sIDsiH68b2ldt/bFG1pqERfP3D1AqYwBE9MoOY8xP67Jx2
vmrFtR+9+VKyu1mpY613QLDDIfCYWoqPYTMfTimk9qeIuskxHfYmJM72iLsr
AjqV8jOV8CcbFgXpesprTj3Bek5pZHS+26r+9G4XtccoSaMM0KGdpFgf4t2s
b251Y1fKR+Yb8HVemhK8ebGT4Dk84u25lnE+BMs8mvmZPtnigq3rLy0y3IkM
VLLMvDeHqeSaLDDCnFFyEeAbQYwvu5pe+DplGktiL7K7v/RzRQpNqminLn/N
eCBG57HVC2FGUXG/NgpTYvCaGQQtFJcVmcelahc65+waidkQxdt8N/02hAhV
wqG0CkqswUb1sXpg8rtMC8Kpom1OD1ux8EAS0PbeRJBJE62vYS4qg34B2X3L
oMp5eUjMRMzpW/pHou6tFU6AjrbIN4MSU2NhQX9GJUQGnd6eVs/9BjpRX2VL
FJPgNPm9vy58XUxSQt0lGUtw9eYggUAjKFvMbDH1uCisxpbBIRJwf4nzlV/s
aZaWgbm9poTwueSwxpGZK9q3sMk6bmAn2UzbXnFm92q+1NREPpj0ePQH6Z0K
NCwDRfyiUEWASPBsSOPhyYwQAb0B+19Pyiq9IGYSqjYuZ7jbu+Q3ZxIwQGRr
4uQ3u+Ykn/QCLT9j3Wu+jcDzNPHvGC+0IeXGcuiadEAMb0Dhy7CGU8ykOdw6
jl33zAc8A+KD/T7lghvKMWIQcs9xtC8r0XIDog0s9fOjCpc7lYDfI5FpHe9K
EaJQg0tGjDeMhvquJLC6O0EyMq2Usjb6DPQLWPMCJoMe9HJUWHBwRUeSUmpF
Qo9bwA+XzcknwYpSox469VRCak/WNoCTqBZ1a4lYIuhXvhkrSqU82cTysUUH
0FHEOdTFBR4AfAIb/H/enVUXYMU8mjqwx7Ul9hq+yo31RLv4N32d0Xecg5Cr
CBdHTmm6aORTldITOwqaAKDmo7w6kN13YVRrn1EC9aXTD8w+XWOdrepPB6XH
QnLyx9AU8C1n0z7AdC9xd0RkgXEGNSckSENGeLT55QbL7ftQNJqVO+8V7KEt
iyF6km3z3ohlhEh/8hwXEJnF0keupMqV2K+vmIiDdXQ1xBW+IycEcJ1nNI3I
OdIP6uzKfyfiktmZHjlzU9qZdDnmM9wkw7N2a1BBGgv68oejBKjMVAEDJxjg
ZdO90TG7Ij9+r9ZbkgofKOuzas6QjDvN8vn4rKhY8Nzfep9YDLKUmTNV3CR7
eF5KhGtuffS35oDKAquqbBRtx5mfy4nY9bjbL+l0oQEswEexQ0/NFBNR1jSs
7MoReUG/Q2Vur3ys73Eim0AvdTZpG0ITrCNwD60VvmACnloTE0hsNiyEpRp+
tU7chHGTFGRzOk9tuiPYRI8Ik4Km3AUeyCzvzN2FGSMfm10AICyLDHHMOaoW
yJNSeen9PVECsPtIe7UTgmAvV33gEkNK6qRRLZDtKvfZsQnvbsbr8cBp37A5
uiNyj10RTokdKgzqSYC95Mts0d4F7ZZ8xTE6j70k1SxvX0k7RXpxc2zkCsjL
LvMVrbRTCoUk6GQ4tNJmTXAs0mdxtQlSUqkcXRGYQOSXXm717X0/9HhoowMG
j5dTRrVJAt0z47E04gwoeugFDPvaKleD8BusBRBqZyafq2E47fCdshR31VZw
t8OaW7TdnSwS2N3j/Ou/ZotZ/kp9TBZwg5GjU18vOH6pe05V28j3eBFRBWqM
zVlgRlBRnO3ie32hiBnwynHCvDobzabIYXIrNF9qOGP1tAJ8lXAHzfwf/tDr
jatnQXOu7vrMaEQNR+tJ49S0GTiHGYEMX5GfB0c00nhMlSau+a5V/eO2yGzF
bFtluss6SeaOOjr+cfmRTswRn/UINveGasQnYvWNWb7NcrRRUmvKchWPefK0
0Rl/HtYXHuSbY1M3Ez1OWLUsZsXDMdoeDZ8zRZBF7AZwudoziLnA9uPQYl8c
o0TSlyaoedkA1h6Bc08dGw3gVoxEgQwA4P2SWCyVLbSrF/zDPXuOtBOsD5dF
Gr4slARc88Tk2xEHCCnABI8ULgmQV538C9UW/iwSd5++14/2Jk3Vop9P7pg1
6XX4Z9pWKGVuLc5H1nb9wTeLFpP8BekldlOnP9S0g+o3c5WWwYTEUxBd5GUY
Y/1x67MZ+uqAH2oFNbZPI62HETtXKTSqW2DZyca7fR14KFW/0tWRBGV4VJDN
n+/t7ENT9NlfZAchGzkBNMKHlTdC+U4YppEva+z/aiCXUzNxImetKXRidgPx
YUb1tQ1sd0nk33V4Gmz0DCUb9XiQ5E9Rb468LYRHXVetPEKtVccZGBqgJXql
zzvY9hJ67GryEv1ErynSO8Pt2CPhPZj97HFchpxVIbOHTR8XQmGqobBzRnoK
XKW1xTegjIhNcooDCDwNMiQIHCX61uG9hstxzoKbb1XCufOHsRXMac6MOeXV
leOTJM3pikNejtkpq8Eaah9mnaS9rBh3AqHnhV2bgYUBc1yMBKNzfXA2yY4q
U1gzbv+VXzh4Z9TCn8swTibg5l9ntjn/5UMo+mefIA6vd35WfiqK2Kphx8zS
TJF3Ccy3UQIaefqULL4A65K1wG66bkFqV4hiRpq8OJJslaZV3pXz7V4IGJ/1
WZ/M9x3+4yqiUXvy/nOlYLGGa1ULsmY7uA2cRinkAsgQDp8unOIje39aBsjU
We84OqDkn2JYdzoRS7v+Ijg0kh09Qxvrp++hE0q4MpwzuT1qB0PCn04qv28X
DEuPv2VLMNUXXrLtJtRSGKw2Vh5YbZUS5gOWizuQfMDlRgO0qti984xLExxp
eTh/ySGA01ln468EpFCdqeB0utpMN3je2m45+ro5CJwM/5hwyzXATYMtlY6w
BB9VaCt0FJibuWE2x/zejMRKdmF9EdEFnLPVt6kU9Nah6zOupLLik5Rh70ET
1PrbWuqSHqrQRKCuuAsOEEZuRRd2SxUnjs/3gXKzNopgjPkjy1u3vwBEXEaf
suQYRqxksoIQVnWmxTJViRzp1zdTfd24BoiO+3ZhBiWMqfLnPBYsQ29rHMYP
jV7mQDAGLYE5RDmivUjnOTFGuuyEw+7mudmyXnNnXgxJHy5xRk54GvTZjPoF
faSxSmCBFi5ngYDsHQlJHclqwsibXPNL/ssRWah8IeLhqh5KUocA6/Jbwq0P
jDVXLStyTQlK7++J+Q1RSQ+SFsaxP2zvbsIDm4Ja9HhUJnaPF1kpFuLehrmy
jNP8hlgyx4Mr8BECKOvO+zF4m1ULFIo2IHS+dt3MASdo1Xb0GmhjuvNKPa4F
rz9tAE9qFbPVTqEcc/fioqwTDDsuYLEwIsun8rlIy+gAJoixemAmTB3udR1e
l1D5jVm1wT3m101Kv6+ESuv96jGNLavmZx+f8xNAIob1JZgHoLPloyAn8Wnp
2ymBPgkPxh8q+9YsaJRkFltAE0+UU9xEILddvMHA/wZ6Mncv0zRBrVdxEXf4
NJ4MpyGA9a7IYUqEyix8W3mRZWSNSh+bCb03h0jHrFFehnzqfH+yFxVChDbm
JNDG6Srn/mHgdoEB1kVilNoINc3DYiLbySzch/qLn0nGSBr+JkFM70bfWMNm
x3l/aZXFB8zRqLxYqcywiZdXa7JdypUp/ywf9Z+d0JSGcivLa3DWnJ0v/orL
ntLBL6PTKGidQ+Il3evXx2IIvWsp5g1uJw5ZHs3fMfyXYTwc1y6z8t8e/nJ7
OIuOq8lugtk+S2lP7J/w//7W4QNQM8oYzO5wAATmcTPrYFBtwfpjeHu89gHP
hrm44HpCi0WR+j9ieap5S+7XenkGtr+dejcLau0pO1HLYX8jAGQ5m81b2Osc
At/wReTnjEohPm7jmaVXuKp1HYBtxLqksaFCUctZ8kV338u5ejtTrfj8VW6t
owGIBQO0sui0I4tLaFy2veConaR/k3DVvnyKD9dzhAUs1LqQYuysJ6UtbKXa
sKhg5pHLLGXkQTEt+pSsXkSaLN+i+eSHb4e68raLNYvzQAD8U9GWq2+AEyC2
+4pbKy7YVLRhL5UIiXeC7kHscHyS3fCEfLUds1sB9nNuaeNMMDIaFIcn2fy5
sEyogTLXypNnfVSvAuu3yIInPfUi10/wojs6Iwe4phw6q02PrLFiSj5RZcbo
/d0dXrRIm6bpoUNsjYIXClPQ3c5hd61hDFUOekjhlIv7zIkBtmEfWEBOflV7
jM7ccl+cjKz89Izr9gOGLzMn4x0p+cuKWrqSnWiYUbuAup4dbRou5KLtsdXz
uO5Mgyd1sCV9sBVeTFB6bZOsPK4IomHGni0zzca2e+6s8zHNphjuCc8JnshD
z1PCa7OxH8a50YqY3K8+CPiCAADYd+1U3VNZGNb5jFROkUWq1+hnRbwRZBTs
ziK8PRQ1ACM5CZbp4zrXUUP+d8G0tn32I/AoKAVi1IEiA0KrSc70E66h2V6Z
5zkS6RnBgWK26Tr2ZEW0XI3Vosz/Y+zm7UF3HsUUAT3erVerFL26HceVPLgd
cYl2ISPotXNgenJd0HeTwzY7IZcwRCk4kfx+f4gxDK623aVOkBGH3VhzXPSr
jXNo82HAo2rIQ6rYEKKh5Qw3FcRggBGajcxOGYQGeU8p20PUGC8vIp/4n5xv
ebvjlW7FRG82l+aQBwHJABjqurG9jvW2ZpAMJ/2k33PlmiIpzh8tvtXYD3+T
N/SBHKo1lGUsbrg35vrwsFRlY2cTVbVzYiyrPIybcbB0/NwVlzAJQownT8zy
WyK6OxP2oASTqkfrkIldsnjIQU7Tt5ExmKuT5+GAFApTcJQObb1p2rXQDGLF
OCjt+TNZc9NeH9ETVrULsoQrCK4aJyoSb7vl2KPA3HnUrQ+D//V3vl7X2UxT
zDfP/f6axGrxt23JnyKJHxux4CpqfSGwNbtZNIU0QMeaIBXQrepdS4dF3rZM
qTk0Hc/Dwl01aQ7DzmtS5UmP0PeAdghNlZoK1IgOBeddrBXU/d/qMhqAKmEg
L+I/63WIfgB5PXL49iRmS51Lrx2mQ1IucltaJ5KBwhh0hUji1LlTsvPXnI9M
XdQu7GH4u/KyPHUQWdbjO/ofYViQl83ti+CmjG/ShwOWrrcFNvgv8Wlt6F+K
AnoZaTJb8AVRZKBR/vHFZ/KbT6kvgo989NX1y2sNktnXcz4agTpEnc4tBR7V
5Ax44TMSmTTjMvWq6GkO8FcEQhpNTqGiufq3WQRxTGpLNhBJ/cftFDHKv/g1
311Lq4rsa4w/nJ7amDd0ZshAFoVEGvt+EltA9pBtVuGpjtWmUOXo7qEl2Wmp
DiMqwrqKd3KFsbEiIAmMmhozn5sBfy1jVbXwKyA9hh3LO09QfdCh3rwjGRK8
NH/WPEuz9bmesKvbVhfxP/i3FEO3zkiwCZQnE6GzQt63eQC4w0g68ni5HHPv
YjuCA0d2+XraUb8jHFnzkBA178q9E+jPXf385Qa18c/T5Y6oKaj7cpgBIgTk
YFMn2xtE5WoqI4DM4OPSBnrxZZsPD6Pqtoemul8vbEOcISyjubSjAKWXUrhZ
MMf2h9OZnX1JDbSIU+pFDOm158TKloV+O782Bad5ROzYe8XqyM5JK0ByRpMZ
R52ZayTbdJ/jB7yUw/jnWDDqpG8S8kB7/ANv1uqN1wm4TfoFNJaMyMkHk7Cm
WQ7q9Oh/s4gZDB0+5Ms4wwc3c7UE0PiEDlA+2ZSCstmKBcdD9YF0RXY4Csn9
st2PH98GDwvbQ1m4i33snHLETTfCT7vgSO+utckg03O20a1Nk49sICJCT8Mf
bypGp2SiMotV4c/Nad4mRtaF2ArS31p/58VtyalMJzkFXHqZ64NufhmpI08y
IIUQtGjqFpLWQi7cbXjmpGW3+KiEjnEixuryEiB+xLJIXu0vwA6HhEBmZgdT
Md9+Ztf7gHReNWA3UtmnhDYHtxRgpHIviqGBL54h4r75DMpO5/cdtg0XUR6B
v0zjMcWR3RUg5+Tr7xNg0vl3J/TtAwYGnYKHxudF8ONFEXmT0mgyWW+Pt/m9
3PdxIJM1RZ5cWk7tjH2n3jC0sbv3RfBUnXq8cfy5FrTPBCwO6te857dzqWFY
jiFk102/eTKgjoIZ4VZOBJCISesiZy1Q9i2qR71aXmu+9GzMskYzsPcxo/WF
eEYfEtzGkn9Sw9FbuJcoxUcSHG3DkNXemg/7+mOVm5zdegXmEv19Bqz4wpah
OJTDIHIaPZ7226DyUtFPx+LMmpILwlT+ekgh+xgzLbpuj60HqEWRBNu3Mkgl
FQVjF49QqYxZK8X7u2CKbP3/ubipW6WCt9gpKW7F/gflky9U7w+sITpSOmLU
Ihki338u2sg/yjBvlf5viMgOWz+ClOV5CAJHfr9ETucK0/0G0x6zbfkxtPoe
5lqooQtTxVFee5JZH2VBp4sGMKtrNrasZoGc7osKq2L09/I8d4zQe8ij1PwB
m7g26mQ3aT4qm8h01GKkTyshhoNw+HmCvdErRn1xu45jU4pr2p1t2M88hHCJ
ZliPtJB9QjLuKsG6wIY5XgUeWpOaZPKmy01cleztG7RMYkPp5KQDkyBa6gpz
m+c1GoUyX5PZCT1iNAEOb2+7cjw7KkHzFvwoAjzhapYpGJHcL8pdAd2rGwi8
ePNk8dTluwVp98GsjACkGr3osbt4POhTTgdDBlKZWbsAtHY4P3o2fjt6p4uo
PGYA5/9ITAaOV8GAGgST10GLi8RbH3XKmqQTvdVXSD9lm9oYpYFTd1kkFrQn
LaIaa4qKW9FP28+V+0yD+sil18OBPA8PINMjNe6ot65yqIrHPQD2DwV1vNiI
wOkcFyIK7G0Q0ndE0fOfqizr15nRM0yE6Lo6MdFFWqws5Q/0NJNsmQcyFjkr
yh6Nl6Zfr021X1qqTXgqUUeHttse8nqG4GWpxCABcOt2SGk6+ddsywrwTY8P
JxLSjL1o+Kj8Jt8bIcj90UP9nOOjJ1QucfMHKDCRJVhhrPY0v3Sal527nWuk
4RVA844Y5OM8wOkOhQ/SaVvrc5yTZc9x0ggadTtQCFkTB2VNnwSiF5di5igw
rSjUGAHd8k+oxqMJnNlBRs9urd8Ec1ufXbhhWKHkoBUTJHvbSaoaO1HzE92A
5yVfEKP0CTeY7olrkdAszG0aRbwL4kCHiEigGZJx7zL6SPMMlZXcRI//oWZZ
XmbiQaNK9EUj4CNMl9Rzp1sh7+ZS9ek8hIqz+8pFpeHfD7fqMEmGOybWugHw
M4djgrVvvarxgEIOzyNzjU/of6LBmQJZPzCeVk1sz6L+ena2Q7FT5oPomaPJ
BnRelRQcpY+7tUxJl7LM+sZqtaD8nQ8V5eWrF8P5X7b3PkcCPsZp+DMo4vBj
3mI7M4BWMllEUogsKbWyQPiMKbjhjn5FkihbD5t4rP5HJHCGt0Lz+WmTQkkK
SFGyavby7btlp+8+C62JJrAlNDwi7M+cFyCPp7wrq5XH9aCEdYRGVJQgpdeO
j1EIpqNjOVJDmP9IAcbuN1rVIY4bUUVCX7Gt28Hf86gFoSMGquBvmJszAAT5
v8pbFfp1om+s9QhqmENWTvka2SLtY5RzfQqmmxrp8L91SK2PzCfo3R+HEaA2
xiBcsTpDWf8T0XEkJe/mSR1BQKXJF/3s5PfiX67PGO6DD8hvH6UWGv1W3Ay3
jajFdWADng8qoVzT3mrYKPKL8bqnlELwWvX2zCArp2ioF5LkLgkCjp5UuVN4
SOFSaQUcxAzogPZEyv8E6U2xn+BdQGczT7JS6ChWN2JaRBgoFZo0JZQgIQWc
uuWiiwUCPreM9hC+mGXanlziPZsNXULskus8HUx+p6TzD37C9I2ev7dWJLNc
amI+LGkbs0AaxeLa2F/nksFKL10Ncb3RDA9N8R759Jl7of2IMrr79Wpmz48z
LsxyVE0i4/adwKyiXhA+a6VY7YzmKJf4gsijPCOj/6w82mIhEgLayJhtAB6S
ffFW+sUWXRLYMZodzYS5DDCYnSRucXm8L32Fq+4tIktiEAN5cZdL9QdSIayO
+dWf9lcSbYsd7ASaweAe75DMzmDOTWlFwmThb6D6rtas+7wsE9Q1SHuOnzCs
XZunCexM8ZijAuOqfSASWao71qlbORcUsZvwm+/kJ4cM8q1vyEFRIovxluzb
n/5qDfGcBI+IctSyLSpYWnUnRDRmnYWb0qsjjVZtEx3FtOmDtvvIbSy1rJfr
QBHq8jmJ5Xxyq5sVtXYDOcce4OnBlsgu0X75FSAdtmhTPynqwWTT28hPDVDM
r+ZX96BYP3cjf5NldQbH386HDtFfknJqhptSmaZ5w0MWB/SnyUT80BWdlS0n
cmXG/TEQJQaKnnUPQr/8qk8AKg30XXt0BqMgv2JxcNoqwLsPJiom4vRCRh0N
O7/k0wnO6kuraGVWIs6/aN9nSnWa94ET18w+Wr1LFICydxPyZgVggLcYP3Mt
PX3YLudX4l6mlm08O+JRt5h26Uw8obtiWiI5HyEhbTgnwxFTQcwwA1XKy+J4
ibBThbpt32iMXUlxv+CnZ3XboaD1CPjs6aEqxJpD8e65qx7Iz+81oClY+CNK
J4HWAr6eK/U4nxSJONgF3J+6xX/Z1v6HRfLoZTo7H+DU1g15gcgNI+JR05P3
O20qaNf2RHkAciiIrNTv7jfZCamMyXHr2si/72n8TDWthcSMO3Vo+pNR80Re
SBmZwkTS1N0iVmwIkXKPWwrjjgbeoLV67l3oEvtziEMqRopSaltuFQo3ecmv
Kc7glgupNbycDSA6J6dnPTnzFIDmvCN8VdxeqP4GLyFJeI+4+/jLB1qFVjzR
ORcHab3VxOlBA2WmGZnAAzar0okXK7PUiLTB5U11ayI7JH7fRPLiuH4pdXfa
pfXL4Dhaa4Mw2nJbg6ydq4JQxr0tCtGxgwZKtuOz8VjMV4wQK3o+4nUkqQDX
pMrKBxZxlzbyXzLb2iBGf3DgZyyvJtuHp5SrsKKBdOnO6oywKRE+EegIzeSm
TaWdq5huevO3kvlY4LCjUdQPfDNadMctiVLXNIfpj1am7igq1XSXwjYeW2hV
yVktdB7SRdRharW28myNsuuUjfhzfJ7rlvTfYFZ7rNLoI/1mqMcNOY6OtU+e
if121Gq9ie/+Gs821MDYBxS+yiTXFTRbUfTnEQjj1kpCTSFyRL2kgoYSnbbt
b4u2yKvs1b8aXp2hBoUB0ksWyr/A2Rj4oL9Qj4sAzT9EpG9BT0ThGrYj66RS
BX2bc/ZrueqKln/pof80dGXOCz+8aEisXevCPJ6clo+FC+H/XnQ8aO+DOieL
EJnPK7GNebfR0IVgyNmjumpf1d6iFSYCDBOBarFurYV8kXo/UkPXfuw1IL0l
3DJ2pYh/ptkGHd55IRQziz/6w8RlJvw1TBv07yFEIwiY8gKwQ3JZueXEW1/W
FR8+Q9bF9CQwHKjFQB2ljIvp6gwMyXkSCu/aSgrF5rhkXmsgxavm9E0Q8R+6
PMbUR3yF9BSxLJGQijAEZCqbH879NZaSVcPi51mUsqWixtfBB/ejX2Gn94Io
2XvPz9top+xV165bYOnZUDxHMeYQYxPZeNM9gEnfpXCwLZ+qI+j6Tj/U9PJ1
4q50lX0yzQ6TuMSzegH4IXcrToAY3xs6mDi65Zu8zazZ+/GOVn1OZi6e+EoU
YzCEiOvIAq6AJIv3FhTrNZuvw7h/zYj05nJzT0n5CDJO1ZsKI+fB2QcIbFvs
5U0SBl8Sx30yAYBuWM4RlxiCBwtYwP4BXW+OGUPe2Mf0zok9mXuzSQoTGBll
uq/zo3FBvCslWJDPIih935IcaFuETudEFrAyDyWAigunY4jQ5PRShtLHltbV
5Gnvul4SyXtnX44a0yu2lJS0y+1A12n1sAKpKrya2tHRnXqwItZ4TwJog8VK
s6CrtDFRSc66UN4CU3lr2fHVVsQLtkEG1Mjg0JnPyiRA2IitinAJBkHVMxH0
hTIjD1l07jA3fJ6XNF8GH0u7lu7uRsGUPGz1hZq79HTtW/bN5U5kK/737eNT
sjVFzreAOZpP+r9GtmXCEokxn7RMbUFXlvWZy7lQ/6bY40E5GIjrsflqd820
VT84M6oygtrBhOnfQ3y/Gf/oz5DnglyXtFruBz7a9fID5AeowkeBaP3c+4ES
hWYqeXaCKmzWNS/Awi5fHTpkIWXBJBsk12Lj8OSalK32znVcswMBtozXCOY6
RqOPmOcMcICYTp46wdHy/MTDR7gOLFSpcH8SUUjMTLULHar40ccaRBbBDns2
n37CfX/cUr1AmvI5EJk9Eh7FNtsd1/vmDIwte8nKMfJRCVcqXYjWVCCuEKD1
hK5AV6NVycOpa59V+SRXnE/geFCMH/uwY3kbqoKZuSXsEgh+5zrpv0ftFR6O
I81AuZ6+/V85TsFBvjGQ5bJBZhBLjTPqFvbwPDSMhpJEMxHtCShccSnFrYKs
hrnJ7ibTv6TDIC7uqGHxumLqpKiDYMH4HOHsPk4o6BJyg/rmuttlv2IWw7Ym
hE5JtLew8h5G9Vte6bsV/rdrNjNFGdQKttARSMZBZYsLtGOHj13urbFi+cba
9KdGix5P4Z3GVx2od1DDoyXtB1zlEuVctjNul8LBJcEJNXzpDIyxPFw+K9V7
gJkZi/hYB9fQ4adaq9yqrq7meABvThMzyZJ5ss7F1u9wy1D4yxyganEnw5VT
JqpgCXdPV5GJl5RVKBznHH6cbfDA2vLe7YPqR8fcZuB0GX2svqhD1uu4xqUo
pDJD38liQp2gkog/N4xShuOMviz3nHiD5bmKmxmT2FlOxCfip9pgVDvdUe8M
gsoDIqtjhF6arglcBz4Km0apm7Lca7ZzxbcpWa6Iu2SDl0b8tV8usTMME2bB
EFdn/TC3f48NoRLvK2jhpmRAIzPktApK5dieuVA8dVFn9KeE6sagMJbHFuF9
+OVF28ARrkRVvIffnedTWbvmXAtYrPoDzKgwPsBOf5A1U/iqCDZ7ubzwwUtS
pOIRMSF6q45Yqk+SVh9tOGhh1vLRFRlZdQ2aQrpG2G1VjLvJBpnzVoLuyouf
c+OSpwNS/S1zQC+bkXj7Y6IZdR92RIzaniPHHb7ExsKCGVTjn2mwfXXt43jZ
ulR1AIhJvBTuGJcgbgLYH8SnjqYf/47qgdchZ9GQ+D0CqqcQFJuj0oilQu7n
GpD/bOiPxpsn5FdgpsIU9J3qk76rGOas/C3m6+SoB1Fg+PyryWuJIMQrRKOb
jP+qEvGAL33i2jlWos4VWSGeuhOXaBPwI6HEuB6weKytCNf01T5FcE9aM14H
O0gIr2EGXvI9KJgqS55jDqm8yFWysHX09xUYbFg4Zi4k2GbQ1l8wzV8wv8JZ
RcKauAFWL89///xyn0fR1FUp/lP4JusIRPA7cUYPO6QNbtpk9yRjv4Xf65sW
5H5RhxzuoEjOaSOV5f7ZIKNYmwqO6JnbW6El8Ev+YIMU/JOVGXoiU5e211GO
V02XxKL8ic0gcFoe74OaFX/od5Jl3dmx3eCS2YC0ydo5yhPX4nYzbL3eLGto
4qi7uwfHU6ET9tQ57QVJIWuVQ0cugyXysrYbm/yg2b/Rr5ukxq6m+9vfobPe
T1fjaGIZk/BFrIi9/X30FOgehxdn0lOGY3PhAecmcuc9v1wneR2hX6Lo0sAE
0LQlMj2GbG2lpKd83qSE6FKxW/ESdrBjENwoSG2FL1ojmGfT5MEN/kRAn6nf
Dh1B4hgNCvJmUz8JTJtyNIeXLg1wHGyei5QuDJyfvby2jS4AMqFO3uIhKkKy
Z7HB3zTluR7aOB6ypDxJTwEXJQDu/aIdTtDYm6OUg6Wyktu/kWJRuajOTKPf
YJF0GQrexKlrw/OoOO5Ar4xWGaf2zWQcvqXn4uqMPeW1ukJV9PTC55D3x9Zq
XmZG2igFYcOTqYIb4aQDGr3Ux7cHGWagrtbyw5Y4Vo0f/oHbNNqu+v/IaqIs
gBoZ/500jy0JxZvYSvp4Wt9ZLBGHbBjfa2QV6jEeZzwlq7d56jfUZjrBnUuK
DJnrYlTICy+4wcyDEqoSs8PEzFlTJ3pOkemHHa9WANjZt4P9VZfwXgcqhgD8
n7YlQ3dKWhhl8k7y2hiFwDfwqItUtgUFZUKWcO0ALJBng8rEKxODcSnvm4Vx
Cq8ThfdJjsZ2y92DnsAEtfxBrm6D6CdbSNUztaj7KmHhS2VSskLxol/A5lKz
D+NtgLtWVitL1tcP3AhhWOvh+D7wXZy+3Fp1OqsUImLwSwW7Sdiwf4agm4xi
MakoWw61Ml9jDr0/583KC2FtCSr2q/JifhIAWL1JsOsy7c9zJv5zjAX3foq/
krleOO4lvQyaXnw751T+eB8rt891lERNhQnZ/QaOJVkmd1OVHXP2QUGJlmgF
kVcRDL7ULTa9+ffx1D/wOG+DIcGivKRNfAlepUf0BuWtHxvu/aApME2poUCT
Xdy3B0zDgneLJyGVxwbeR95qqcs11kbO6HnELHq2EjICEx1BfZpHSpNBndo+
Bn1AIZQkoCZai0+PaSltdNt5rldHuiUhf59I1H518ZnWBJlJmKrIKrD1SFWA
AOojl/rcxnI3sKkhawLynk4f1IsfSc2tLsVGl+rIEP3LzXIKnndaFjIuQ0RW
Kwotlr/J635yI2hcj14IrChrjmFvME2Vm/nQ4OfPw0xQ4dMVIkXgeUr8m8UN
B52CQRfAH9s9ajeezsn2DmM9fzp2R2iIAyNCDD4R7OOmaaC2W7RKMWdT7r9M
PZAF0W9XtnbY7zXtRo5Wv1AsGYq/r+R3SjnX0xPlmjn5eu0vPBG9iokGVFQF
fDodwMQdhfWy+mNd1+QKLqCubSrvv4GXYUF7DTDxFVSBVoSse2DYHLRhd3s+
TI+yx9k2Bg87hZFEQvMIUu9Kw2IlYrXout1vdXm0brB46NPcIH7wk4z6/2cb
/9MzIoGf9Gu96ce7z27SLcVTadaNwKcUmJc3fGjCSoXql9FNMLBcXBxoxhFc
nBNN/i+VK0B4CZnzYMquKoZFZCQPGYiE6Wwq6W8BVJLPVyjfrzXcaH/xdoXr
c0TRQx+ngKnttTiAeZjRBuvVNjZqbFTPki2Flt6rk4kKSxtcbQDONAAvQglA
FcKvU+MMvQH3V1rRduu2TNjilYh3m54MpnB9JKmaYUWAiB4tjuqWRkajrNsw
tbANV346aqJq/C0MoHF54+bxDh0xGqP3Sd81bZ78J0WnzJMQE1l456I3kl3N
zbx6rLZJ171laxi9zR9YsNO5uZRbowKAPpxWjbhJ+u7OJO3lujfqtLwoAz+z
2eWod5CWfhg2AWsa/+DK8pnASnW2HenMtWQEB092LZchyR7TLStSXUcnaloC
Vp3CJAY9OVU2HtXmVLKRi6L2OWR7rb9AjGF5Qda8Q364z2w4RczCs+dBqbgs
YrVfYkhva/78WETZ5qUr0lxRsj2LfNCXJXFGxHS/GoYW06jwYaTuHWfiQ3Jl
nVueg/uTvQ/wvWU46yHcMMUACHxQnEDPByJt4Q8Rl8Lty4b+GaJR+FAUeLtf
Bt6spQzwKM+OIEZQB3nTf4ob/vTkxfdk5rKIzqsiKYpufYYYOYQ8kcT+pCAF
iTo/PiL3FctYDJ8DWYnb/8K/2S0Y56DoDhctDBJ95aS/bxQ5CO4cL6rpqmQo
6i3AUbzJVYt6xivp43HuZdxa9QF7uv7YVg8/1rG9AHiMxttFjz5RDL1WZ1Xv
PYzSkPfDKuXA0ihC5UYK4X/V7NkM7v5I2ae8ZttmKDolYaTUyvlkasNlOmoe
hJDBerqd3SxbH+Iz5mW1vCEdZjlZ5IvpKF4LOyVAmCv6xzH1rulSW0+WZHS1
t5vp6/nGjFEaRc6QDTY1OvElUq4/sdW9PrB2kyi2i+9VJvgLH4OaZ2QG5oRB
qyRSLQyYheLPIDAQGLeMfo9BT9G2x9F4XBMEv5SJ1Yf407DTmC5YBpMxQr20
vBcRkoAMYNNkQMcBn8OVPE5i2k8i9hDsnAbkmWW3lQkLvR3RrrBHZAFGZcVD
/BT0kC7AIrrShIeMwY4qlDZa3K2INv0kvrnXiUnnGW2GhVLofmdti2o1z5ZR
f43yWSqno8+pO1emE8YdRBcbDlGJ4EQJvLYEND4TvcKUn+ahbURwrk+rpnVW
QoRbaMZm3L9vqO1w+hCGjTvoJVCCLFvfhaByyYCJD0CyXtQD0vkucilQPNJB
0Di3bsXc6UY3DePQ2P49CpwseGDsjjIgECKw4MevoSgGnPb7UVAqu89hXCGO
6xA2hIoWvCRC6QHMzfmq9qAynFDIJUKx0n4ajAqFbnJaYgC0HcCMlpj/Yqg3
GbAfedg7blO5CAUgVYiUOUVXrJ6dEItQVsZxWsxQCrZF5D2pGQkhAtaecq8O
XlwgdidO8ClJn2c0SaFbh+FyA9jBPtlvYHpy5BySJ1eC3K/ZYpyMAEPyJKeY
ZVYWV0IWerHo+8I82OhyfEnejJEjmU19tMyuOu9cKWRtCSGjj5tv3eSz2UjF
wlM3IwxudFXHR84c6bF0S0yBsFBzXHFDVf6j7Am5PwnDw0nEG+fmgmJuT0/F
K1eatjrYejzbBFa2qVt5ZdDwDaDvLkXXOWQPrCnHctdvU/pMVeMN75ZVHKu2
2/mm0UAR1wiUlU2v3eddnYNgkb91a+hVkgpvPAQS3SSUWMa9l3RwnD+Z1p7U
yrkjw97AP2q/rFVxUnjOnzUcLSgBpH0LGJXflPBBG15ZgnrmV9RQ4nLqdU8k
NwMByTZ64Vukc7HNcST6f6PyapKEpZ6BOddesBVUWV68WUp5E/9uisu5ylI1
nBPpvVQce/NE2qFz6aMadsAD+w/qOQQZHuaP6SBfz8rEPGSRkHOEfenzpBVx
LeUhsuqHCakelQYv3HUYrsV3NGzkzXNJp6n6VGfPuIfXS8fEKate+fNKffF2
sxcDczNuAqUcn3QgtNFXKUD66UvUj+ONKBhKHeibiyJige3qwEcmUjI4/GGH
5z5VCV9T03CKkR5cnLwKbiLLk6o5KQDhfOv4HCPvJZ5mc9Uv3TIYsHGrGDkw
JbqiYMpLvF99Xd7ofuG8jRuqO769zIo9Oys3Th6NpFsabhm92z6uwsZ7bpwc
wmFw66EH7eJfK8FUfWh4QIjiq/x+BmMOBppntMl3tHZ5iPqWOvB4+2LGH3S5
u8Os+SKeSbHT6Lp5UNNb/Hr6a7ZTMkDos7aj7KL2QkHo0Wo9CgDUiSDVScA4
rcVKua+8908Nk/FMXXAjv6nhZ7eTq5euMBswh8VQyOLXkC73elq3Ttv86PZ3
XjvppEogXaqStsr3o+iSqFAQu90I1px39EDsulHcCrgx3y18/Y0l2udIoXY5
/Un2uW9L74KpMml8krhkKT/IOSJF3o+6SyZG9MaygmLD0mDGoRE0cdXLbtLX
MjexzdiprTv0+A7CnjBXklp/CMMmPXDE0xPqfuq67yzjSGg55rbxQ3bCVmSF
QLvsejRDMDDIIxh2uY4tZYDdiW2Vmp9YkyH1IrYsJcr7I2FsN91YMVfx8fHQ
8L5O2In9uLdVIIgJARWVeMFmO44n1e6fvatn9CAHn0Bu9FZA/yIXltOigvEa
7pwzGfuxfP3kYxcAXvcmGyZFp6maKbaY4RPmdZv+bM668H709eKA7Hi/d95R
5thrsew5rmcO4hK5flAJ2norG51waNvcAhDe67msLCwXstxX8GtBKTf5TCUp
y6FOgQPH07PQQKhTnBTage4u4lbsUCE9XVs+Zq1g6JK+J/fiIpc8GAJyJF5q
9YTzXtGIfKcfkzsQMFtw17Zn6UoTRXaMAf4WRL2KbdAmjXorlVG8BYOVuwy2
7Wrt78rIAcihFKUNrZn7tGj0gurnUVBh00Vhcs4TXiTT9KWU5a08FjYYXzda
zHqfRBqhROIJzu7/6+E+avRy32hYaYAv1w8WSK8Lr3160S8LqF5BUYxX77Sl
tDzzq2U2W8Eso9NDyBQ/QsxX6dhQxKD73uuBi++aI3/MJ0iNZYAaozGa6pzb
ksVk2LKVg3AECeO1YB/VlXJWVdtzM7kjSHCP2I6/WbH4uq3fpqtBByZIFQQe
pPAzmFKUuTwWspUPlhu6f5W+4PlZadvWJOtqfU7qKcP5ApSN1FjmYaGamgC6
nLNj68yTr/as0Wz4pqPV9v0pRuw38SGKF4C7taut3KWqy/5+ELI1YjDxBlVf
TZpjtKwpZUClziGz2PVZOm1CjKn4gL4nfG4erB6l2gIB5GjHcIV8BC5sFgEE
mY1dY13UEv8WyoMO6z4oKYTln5Qy7DjcTVAU9r2yZf/PtztLrDIcZgH+ja9D
BtMsvAxrfZCnmzwDNi1Kaj/n6m8Snqgt0r96qFo1s24uo1F8Iej8ve+jNrUE
fOT0oPhTBtqx0U8NgYQtq53g7/s/W4KvKsnHFv5PTEfZ4p9HvlyqRuY3XDWY
xCAAmJKhJqj/XtZBcHWipVRhh6d1wYmb8oZ+LRNrzAlFHRqh0YSfA6Y+1azr
u/Et2AfRv7+WqcbT3RsHF3t3QzjsAIAB6ENCyM5BuqemrZnhnPT/6MsUtXOQ
jTpExex4z2Xt2xlOIbxdA/2476CVBXlfzs61bytb7MqiCe8h+vpyty/fLSzc
3IgNnkADblEDQmEEbJkDfAEJUxck0zCXgGSjF4vh6wmJ50wCIW6Pg4NnGq1s
m4VAhaheV8zFe+b80LblF7DSGyLQzLn8Kl8OP73YaEWNrhJ9N0d77BOI49s1
rJffu0EhRXB+4ZcP1gZDJqwBve3ARrNhhx+dhOevJckWVLqni4ABoj2U+KfW
YEOovlccRh6SPZP0k3JC2P1SzIL+/zD9IUGE9OmgSwGPpzeKNqVaricHBOQK
p4TqG4hnbTZYX72V9MoiGsVumlk3PEBBL3VUPfKYtRqNVi02RM2yhc9p7vVl
lACyuLpY4q5xxBixnOTRXb1Tcq41S3A1ktcmArpEE4FDILelFRN/ikXGqH3u
yKjy4W368rSsfeEF6xsjEGQoKxxzSrAvP/vVTonfzus2i8fzj7B1BZQ1BOGN
fd4Vtu+70k1zPhc+RcSOIwZgaJZF7IUCUkt/W+2r+x/Kn3w24jrMl0BjHIuw
mXKIxcF9VXGReadt3RXqy/CrUA8b5EG7zeI3AnbObdZiKVuTjYZsgenBVdC3
/61KkSD/cvPb5ev2mz66nuXkgsGfigTzpkCuY4yF3jFN5tRDBm1q63wIVPmG
DvS4BtYp4uL+ReX688JkFcsmbBQlMSbxeebKsXhvQaM9bfMFYmFZU5tE8v/J
vFFlZltm6Wl9x4zjFgxDM62A7neN5CzVtzk7hMjAOO+2m7ZApmGRIqal1I2F
+2L0btPXAO3cAvur9YtW7XyzVr9GUGZ7mOBrAtCGd5gM1ggj6sIxE7wZMvvC
m5nyPAWj+d9CjZ6ZM/iQYaGeoZTUC7Vub8cCsM0Yh8s/N2YfvaEvEwC+GNna
0uJCsdeEExo4ZlxFjfP+XLxbe+6vBwXl0YeCMFAEc7gYGCk9bW81gvTC3kTo
Xc3HhRUk3egVqMsTLr/rvL4DMOWoKXtXSk9enTeraLYYUYDxInMAVEQg7/gs
s0kD9tnVvLqTOz8AR6lhL4lzNarECTQPhstZq20eG0H7MDI6Uf6ShThHXLpg
Chph4H2yX2DSWLGcQR0yQ+qhNd0M9VVYusLIGLVGha9MZ84Dkw8gBgoZ9cTF
GmhlTfpR/WRiPWfbn+IZe0B08g2KRnKmqfiEopYeQBPH8mJWs6dqcSZrPxt0
gtq4zTdAtjtH5JYVoTY0Gy3cUmMaBbKpJG1hCGOXZ3Yy7p0j2iu6pTtFkwHa
Zn7bz24aR4ouA99xTIAHjg9sburn1ePeihV3QJEOp//h2+T7f/MBLjRII9jE
mOEzAL2u6qekPY6jPD1gjDvGPQMZZR9MucziXqDoPPCiueF3N6Dq+R5xxVs9
4z1NhF7Q8lGGWg2LRFu/deiHvFuEUgdhtQECOd0jkLYbCT9ifjfnt7t2ESnw
i+LECamU7yb0DcyWNc68Zwj+gSr4kCpFElymyd8FAQSL9tUvWxAJZPcEprIy
eVAFSNZt3FJzqirXoAZjUaFRkhQtumSmFVXkO9Y6pTJtEcrjX6vbF+mObUGe
dgmx4ZxqpRrlT47LPBlJhgFAI+pWbjxCMubycyPinXnTO75D9QgiONINtZTu
4F9HT+2E6XnSlI2SecXowLTgI9n3l7bpAvKmqtRN32OqCrQ4Cw9p2DYX+JpH
noiHZ7TH0vDv7k7nPip+ZbXvfa7UzKSOLfxh+cmdDCrB3A/vpVygN4MYpMnL
xgL2jifQNZDSi7yl7/mWecTGiIBkI3daXaJJwNPNZK09umgEmunYCXLhSQ9l
pu52oWu9vUyLdMPmvf95dMsAsDkwcOindMVWUO9p/NTQLDa/Q/eLT5SKMCXq
UWJQ2DS09nIHK6xzXjX2TI9qliuQykgXsaJLPY5sJKyTxvIDhTqiMXG0yiXw
RpvEtLI787Zk33DVPhkAxerXc7JUsTyBIApkf4kBRRbBp+QeHIZgzvFHc+ro
/nwMEmg4GepFXASsLEv1Qhq7LfZXkP+uPbf4I6pTZdyWfnv/h3hZxBNnn3fG
FI9A15TQK+FemW9CT9ahrBVETx9WD6R9J6oh7BfhRbKWTuSpToU6pEGk3e64
FbMwPINvWgeXM8736+7tzq2C38InqIqY6C38qtpbVDoeiqYHKN8f2yPO3GVI
NA3VZ7MZjLNQqHKvU4DkzKY4LTOLymcWg0IW7QgKWL9lieOpSGchwiUfNFAK
wb7cZx8qhfF9QhcQ5hzJIyhRGcabTn9C83Pi9rhJderZ7oAhu3HTRRw9bRMC
LYIwoTCdN55i+WaOeVCP9h4GJa9567Uzw4EEGEmY7gmrpznx/IiKraLjFCFp
kz+uOzEck7NR3o6ylKKIcb8JkGpWePCpZCtKKaiiS6KUF2qRQaMDkgsgiaiR
1xsdlaNqlyU9/O5r9O7n19OcePcs9cGAlPErjDj4g0zIUhwCx4t2jqxrEmZX
yFwJ2zdxVkDvUbPgjEU+Xg3hQYEg53zzRLKc7mATeUEj/keaq8fYh3sy9COz
z4uHM17fCUN07/vGjuZYwVQGk4NrFg7kgBnPvUc2LT2ttQFTHJwKwo0E5eQU
TYXSX2HLc/5IQFCGSfLPF/mEG/YeTdoQj1H2bPzwDBZYqqqXeS2sloqfjLMz
g1F5Zq65Gz4da/SVtyj+nTfrSPuKr3U2jEkD9UhuDt5iphMBj6zY+UvtAA3H
fDKtEL9wZWT3UkwMzk7G+UdFi6KoSgjMs0Q56Nadzn2HfZ3Kz4N5L57oZNVW
vdCpzUGgG/BevCF5Rechaippy00aJcJTvL7nZoq4bpuCAI6i+RoNCFWXVv0s
qoEbmxGN8mlleNovJBhfPa3c6UZjyGd2p0L2pKqIlUMyD5EacAPl+0GTXY13
+18kdGJp8dRsm5Y9bF63yG73GhmlB3L9Ol+0WWRj6H6iOmhHl7xCIjjQWCjU
ZkzU5FnHUMTqaAnHzXrwJQqbT2UjEkEfMDSe4vCJA/jS7gWTkDPYknZqdAZ/
RnfA8HhufFsB6tN3LvkFyc6OD8EICK149eGjyNx/X1OnRZKDYD/HyGNHvZfG
PCVM7BJb48V6YihBg7JhgYl3gIdK3Ozag+eJXA13t4iXSAT+FeEwau1yg0TN
u+1hHbIEdSu26Dgxj5sf15MoH98hia4xjEZizDRH5TtwbWmGbZoiEfsK4/fw
IgqFSf2lNvpUIfE/h61zN72N+nGbkHF+dJ07hrTe4z5BsyPyS1ggroOMvwua
nYEm4lNWB7KCn1pKr1j1mm4I2TwHbOnAAE9+t595Py+/U2em/uYQ3gycnfzj
F4n1UNX7A8boQXLEJmJuYMYaFTESm3rTz6XsLIrK3iDuwJV8Rn7GKn68w7HJ
NsiEjwi4gP02chXu0kQqZMqvOWJ94WzaBFDpmp82OODVDFyni62DNX4pC3fT
0SpV8EpJ+/4JG7pNCEi6uXFSsVFMdduoaGjh7lFVikjFicrDYjNhdhlNdD6a
ZymMtc3yvmSXUCo5V60QAzhdWAYKpTuIq4BcUZt+uEEGlY8YoMgP2MbTJyH1
6mrCkR3/YYg+oj4VU6n6xIaGkH3vw43/vlCYuIakJLlRAD8j4mJbVUdTJXXw
6sG/WC7+VAkFqBfBE+OGK/mnMtD8cFyty/Sr3RHxmsnpQGz2XSKnIU3VktH3
wMCI/9I1gue6c7SbAOU02JMH4cpzS4S95kKB7PYRn2nGH7/EZzLxezLe6/8+
gjjLi27s6HIjunVaDm+MelHWvpysqoJltXFxl2UFGNZs1C6kENAzSD/cf2ea
zRcEhJV3c1L9IjBTTumOn0AeRnFfkzSGd0vbmzE/a9v34MJ5+S0zj4nN56cU
wiHKrSqJAi5uPX5wfraXoe3hFC9+6cgtkszI6wm+Cw+gNO7ArC3mwR1LusIi
2bkR2EbXhmPnQQpNkQlp0Ehn77lt2AkAg3cVKgRMXbh5xpmSYEU+jgXutexL
wbYcANaB86j2biKO0SyACG9VXKbq10frh0Rn6+YWfs9xGsDo/xgy7jKrw21f
PZTPFTOpmgLK3UaH/h/dVdmJYuAF1/b5pnwCXlvuUEbpsXKjuxexIy/kEC1K
nuBpkTlh/PZIrXKqF4YUztHpchGKLEwIx01bZdrNumFgqPBK9zgoXzGCqdqX
foHglxTLOLGuSCWrWHgKeYeTYNMrRESsRIq9VgsfybtS05uLWpzdPHSKVRUZ
cpM/HLM7Ui+cxuXnYJn5DhKm04tcK9D0BW7ttI3lSc6WPU1im1uV7xlmHjwL
fD6+UHnkhkNF/LnPupALmlhE2tKoZ76AuglobYpxi8wtrF983DdMeVDd80+R
061XD/l6b2UaEFhtfe9h/XDfLo40Bx/dQgPMKxxgnQg7VeP5pS8yo9zSSpb7
oIIyyLnkf9yHDgnRbCjy16LTKt5ekYTlxfoz6RIqe3VEgr/pNgz3Mh4yt2pC
qklynkfOwDCmt3bVqJig8vpBc2MAxc4Ca1F8hjy+xonvIU0+RYMU03CZSZ/0
pD1IzHn88Or9oUjK+Cg6Ek/YCv2IkgCFX6lvKbFUe4SnbXeETa1VAyAccH/K
Spz9NeFzW0VlcMvZ3I9p5BikpEXf0iEXHxrVlXCtqE3AqllDAmIL8Ho9ZzCW
D0BeyWO8eQ9TS6Rz+5d/sPy0twdcH9x1ZgR4SlosPy2Mjglxo0U982VM1WBu
blIa6yHZPeMx8ORZ4uxaC4bRkir6nwQIbNcW9C5FnlecTCU913MotKoYdBfO
jpfLX7wVAQiMQ6qHH0HiR5nXOZokl6fkcXvfCU3etGA2oVWTTvui1h37e+OK
VGActOgLuxn3Mr1U2gDmdfzuBgamK9495rjltOQPIhOePoCJAyATjo3tZBdk
3vsRSoiYKqsWgZWrNqaXaaH+chr79sh6IRuYtqIGdM7xk7oNMiriubmaisb0
vCN9QzeYfhoZgCH1BtUon1JiWUQXo1tbSfpJmTpoRAjP+TYNysP+1s9z+ipk
JQsb/UolqQRWcSYJwweKncBtbHbjVR/Zn0ZLMKykCY6kOh/I7Rp7C+pyxeFT
KKDMEgDesLUiARsbWngkZSDdMoDHH6jeb8Kqxmfw0zPpThXqHUHBYR2nIsV3
lHOdJG4PfmL9aotuJnVfGj/TBSIs8016EsDfUkaN3rfvqW3+6XjQkDvv0O//
wN0bTaehEJT0ayC0q2MibxEBi9tet54T8JRY6Z7mC6AXeihOc2Ljf6b62OZa
Svf2mh1R9yFxtddPjPjgX7tzyl2xosfjoPZHYTviBtLdIdBWiMNMsyGk97Mz
l/LPapuW3wYfrBNxuBSPneYYzYKd/CPfN1Q7JwAPUDuqJtOGOJTrfI6R6EEt
roTxyVOLbvxk6OPFJwFjpdOGlJTjFl/K3fwD2TxU+4waguck178vfq44VtkE
oRn7dLhxrKiQjGo/H0YmlQ8YGPu7xuq8a7RfDN1G3rBIMlIBd4fb1vGttvT7
358kAyPc4ky81SajlRN+db8j6GOnUU04sYbTUi/DkVGO1AyeX1XWeMBXyuHh
KXRQV3FeGA0qR2paHpaPil6TE2wkTmYquHZBuN1o6R49E5T4MMpIuuHUbNcm
TU5b6FM1evELoMrDOg5y9BJpFo+wm6i5VboWkWAmuUFU0NPfMB1QMMDujpBw
5M7gD3qwr41Eg5arPKo9dV52IVP4UU3gsK433W01kgZCmuN3uEz6YzFqtLdB
L3oTah8Ef6w7kJcWpAiBAwFGAvfp9qE0rCa7NB6UE5FXPAWIf3qKEd04ek3O
k+bp0w4/ByjRHAWPvpU1MzQIthhJJ2pD/16g/MyecN+BEm1SkiqjMkLzUnCd
Dwrb36Z8zTq68csuQ3C2Hz3O6IWvguHWlvdQFoYEDgSvoKAa6fx+tjckNmRn
HQXYh7zDzvZNuw0Psv7CalICgngIE5K98ecdasndOmFLdjsmPxDSdn7vTZ37
aePWVyCgfO4OGz3URVOwvou7t5JPlHC64R2UOzFjiOdXJi7uQfNOQaTAs3kp
+mZ8/cJ7n0u+yGkkl4ErO/grQKv+eB1tn43SQCCWSRPdZwbb2gbW5zn3bWwu
/WU2Awcjb8FqwB7scH+/szR8iDs8SxcL7V3NQ1Iqu/Og3vMEc/O2pnXkyR1y
h+ScksJ11oL7CGMK9hPjbmQ0eB2hmx0HAagjscCm+Mcx7RBPQIO96mnLZ7GV
1LvTYqxu0JRKe/Nr/c4dfGqMOq8avYGDm0qasZR3x/cYw+gBvpQXNUXQoJAk
HL5OyfNxx6jDBJsW12ZMah2WAULOfrDFtpg8ox4m3fVXKWGBkG42kwpXvEO2
HE6Eq8tr1rI/3ajx7M0t5s7MUboKXPy2jjoWbPNIECmukL8lkNbasaem6rbC
7bOERRVDbB8uRfzePDoIAb6jRhYSgEwdVoya4ChfZFXGQyihdeI94+i2BtyH
HskVuA+/VNtZKn9D972AT1U6vi8S61SD5acw+yVc3/VJvmoa6BnXi16Z6InM
AwvKZO2nhPZvE52GYmDwu3IIiDyiYpMvCutMQEzr8K7rnNZZRQYU6E34/cay
hTKXiE+HBRiFFRpYpzsbq/XIyVZMftrS9IGr4PTHqfYqfeV55WAa1fGjG2bc
vJ92RxTWCBHtYtVxJwG77e8AGQ2DV/kFUhUjf7CRlWgCdBmpbkrlxJkWbTUv
3crGL4T9xoDQYgUGBsk2ntCJbuf6pWM3fCVGm1xeSa+SuH/UCwD3ieDTrfgK
NKUbw/34EJh0/2nJ1sSXpLccsA1KPQrWKWqCz68lov+8ic3AjDvzgfvMc6UD
xa43AeyIc4vC2d7nInrjOfL/Aq23B4i/WMWMt8C2Jy6Ka4ThkK/Cw9QDwAjV
pNn63ZjRX8GdgfgsFsGn8kwtdX4X6z2i8y6Y3EDDU6GfCyO9OjcYxTVwh13Q
RitiVmIWojV9c3wKbUg8qOPdcJ5GIZlSpqHLezFFGvJ+pYr9hBuKFeKHSfrC
puxw0gShs2FfCktN8gXUireyJ4W8WmcisV8a7RRIH+IPMuOav8257QZN965U
vucxY5sLnbXtohXEHNnFWHZsJssovLokOj568WuhfyYqDnMkH2FYBigojPz5
zroheExv1lcyR6OVdS04C6dlJfysh82MbQK+Tf37kr4Q2/AgORAE2cbxRewr
WCnSrOMSwtb04AznKqBFY/MqSL04/swJXlCjek/k3jBsjfTsj1QonrDgaQyk
RvXbRSDQdui0Hg9wsR8U8fkKSms+xf/Dd+4p9ohp0NyE9sikFBORIITNzyYi
fuujNubxUwEzvz+vd0pLtmYcgOrdWA4w9Hdi4MwxRZFv0TVKz+4TVCJ2/ptY
uBTynEeIw5sy5egBVtC7H2bi9fRyfA8ph6I7Vfnt0EW2No/muZpxetBOOneb
Ttu2Rht3LgHli3q0LYAqMPHxGse9p9Z3LeY8QjptM4gzv81SDK3K/KsmMBam
3CHuEGyJGJCYHpxk+x/1ITI7gb7jB4Thyzi07sLxBh56as/YEXcLd71WGCSz
dCnjMHpXqWXcJRCXujLmjI7IaG4elWQmOSa0hDfItNcvJvTlgv/nmeBTXtT/
Vv50tKGmDz/giZ67fKZj+gaDttKg7Euw8EpNd4JNqSm9eaiU8sVFXBSC/V7R
gNs0hAohSg7f9L2sNDROwYwQrZoTZ21UjxrcnY3EqgZcnZAhoC5Z88LB/m6+
BuQBsf8FVCjq57rGDi2PcD1/IebRzJPuQBzR4oQHkw1ZFhOV2ES6vaKCHatn
ZUMZ0hrZrAYgV4cs1EFra2DrGo9sUxNByj313oMLzd4Lb06rvBPJn1B1S4hh
/jVEFH8eEkaeYDCAG4P3VRKTxEzxYBajL1+pLYeq3s7v5HZKZJTYkVVugYmb
s34fLJzJK/DcTF8Kfr6ir5I6Y2a+2GJTh1OIipOJY5Qs2hiadMYfKbTU08Mm
q841PIOSxFmrURJ6A/2QfKOLoyELR/jzS+igiQGa34IRRy1ryDVNJRkDqGbJ
UkBh2k1cFdYMAOj9hAVsMJEMqxmkQOv/n6LHY/FCE/IMkRcMrGMJe2qkvLGR
KW4mk7EXqm5s1tfwLvLoHoFO31VquKRje3wk4GAbDNe8FA+r004z9Z4iELpg
okLDH0Y09RzEc3Jg8gSOYMZS0gDCIjtR67jxTIYyOXwo2tebv/+IvVYvgeRT
hpOzxCrP08Q1iv9TDsF0wNkKDLzXN4ehFufuX6zC0oyCVUt4L7tJ/kGGkQt/
zTIIUAP7MrYWjvkeVmDYDW6zZimswDHKCSKCFb5KrXTbYOI1S7n4B0CzHs98
FXv3ARCdzKyNoyiMrMktsA6OrMrtFiS51iOw8uWVtbN5lM5Z77JA5+XywYLy
DZZRZFaUKE6Qhq2tLoqMbaQSJ13YLztliEyzo/KYV54fDbJ/5beiSoyflDQK
qpv8n+6UFdKsNOrOnHtc36dZ4W7ub+3gyv0PRnUg/dfHoY7Rz22lobeF3dl9
ZQD2Aop13371JZkxfg0JR1xBoKG01oUYzv0O3UdygS5+2CtoDiMvUfGp9BVs
p16YWA6AU+UrAHEcmB9Al4wBHEOW+yn7XeASncXBgWp04yAo3RtzQZ3nD4HN
GxnDMdlUFtit5+nHhooDpB0dJiabpOV7fLtwCH7PDw2tI+MSKIBEhBJ91nJ9
DRfSC6f9sALFx1TeFEp8isy534lfgrmPfORGjwhIkcrCpk6jfaaz7JGV9euV
ci+Zzi99PKwlGqOS7Ysa4cFEAucdWmWceNa+013skA3YzZfwz0v6o+lfs/hx
F06UDJB8OsSJREC1C5Nf/Vge7BD9YvCFZJOj1PKCm89ru3p56rTJ0rtdHF84
/dA6T3aQYVfVpES5+Aedicx59O4WGcV5Cltm+1QN3vtf204z+Uy+6tFI4d9e
4WcVGF03gZ2lJscW2gFxh6veYeXOPNVDRJm5rn6gjzwhIsWl2D88h34Hon7X
fEm3A6Z92NUI/Iz0E6xB0Mfrkd1/ptmhQ+gKgHCyJlz5dT5Og4wwHp4q5byQ
3wkBXxUCkgdxt1FxNQO9hF7aJr3Z5cue8sbgkxCgq/V8lAiAxHFhk4r2o92Y
Z5c1I4OSQeuCmeNBqMA0JNufm4O2UCShmbDKV5PZ4aU3PW7BGJ78HMsBd2UR
az1+5vB1NysYNKqn5UVutgZQyHRtDY7B9EL+pBY+TW9sSEbD0nAVFYnE6QQS
X91bsU4vi5hiO73TpAABwsC1kTxwKzJwbw94Jtw4p3qPIQQ0QuCnfgaqrSD2
7p/gqJrw+2hXReorh2OOkb7KWCn/9POrwGCdaGWBzENCs15WN2VMlqKRkimu
BH5qjEKhkE+EH2YceuNJXNPq4geKK97qlKYtwJjQejFwQmRhAmOR7sCUuSjz
LvS6C6HsuLYLaKPYobm1X2RcvhoMdlg7gogeXoFQZDmSjbfBCDxGm/HIvypX
wCF6YJY7d7RLeHv0mTMNNxGx3+McEPRLiNbtxlaOLQqLNuqJ981q/+aITG3I
vr5iEHaB0wAiMwpJfW74OK/q8B9Bd3Gs+nQiWAFzCHkfvLNchUd1uyGe3wte
0ABQ9Bpx43ZxmLZ44TTIJmSktaPyvQtWj2FQgh61EAFYYh7tzFDYGNCISpU3
FR7N1PEdb8LQwOZ5HBJ2dcWw1MuVS7BDT5Y/54jz/rzCqCExuiTUadlpHFCs
xApHhL5Vxuee9sqItIdPLbIuIbjt7i5EU5kh9Ae/0pXSrhzhV3av7YhuyJEC
Fg9W/ZgsMS9hYFrkFXZat9FsLczZHw72iRkpnzP+yhruwWNnvoGddSgMbaoQ
rUqA8qKkTW1V7HEuid6qvF68C1MPk27z8RX9wpMXcvTQMgKHN1tDkVd08PlK
K5/s56UuJDdchB3hbBSuZBQhl7m5wg7Yr137otL8alxr9wJh0TNKTbV61ICl
6iN0K7gDv+DcUYK1MmmPA8pYO5D1qgmfHekdKs3EzWr5N891nGSN6C//6QjY
RB7jguhi++BwYi8i5A0a9Y0JlW2utshWMm/XwNAj30QjIxZU28zLJbhh8ORD
OrthjHmGK2g2THB0iMPbqt/68EBx55f+o7SvJicDLcHMboJ7J9RMr8Sa61zn
iTrtU1CRfmJ7/YEFqyrYBObXpQlbOjbnU6VecyqrsIOpFPuHtoA7czC7vCbw
oJL0KRBUpRQ1fSyrsXptV6p+MF66MVbDdaR7G0xFT21tl+mOVoBOzpsQ+5uo
4CjZ//R7T2muC3BphJ4s9IXnP72d5xjIxArYOSnNbjQdpxXeNdueZPe3/tfz
9JxkRIYLKIsvnavTu0bBM1LhA1LrkrwMvW/uZ+cPuT1K9tkIjlu0YLcHbX0m
STU+ZtxW4iuU9h3AXWvcW3DT0n/zNBrxzmrNZ37vwC16SYm+JbVjpLSLeBmm
9WbrV7HaVm5yr4Kt3AQXTTlO4E8BGezNvaZWpq7rzBE3eoVEMlF6lpboPwLm
abLmCee+LGBaQs8il7hUPxqz+8kVqXIKU4xjBQhxzhEZtMGLziSI1XrBOLn8
rlYpV39lTobxfifgG+ACvFkOzTBa8LoTigocWXhLgfq7OH3o/2ftutjmRG05
PwcyYqqbQDOh4KBqLD7iDEfwbDyU7vfSruZzqyO/AOfFgHsdT1Pfj2/AMecD
DlAhiLEVZVmr+yJVGU1ZDc0Hw1Exhv60A1PPaXT0A9+TNIC9Gr/4fniYX+xH
1CT4za3wVhT87JDz08ZbnpWn1iUteNHHZcxoL//aIszKevKVFxPYzMJgKtel
56R16x21QwGlUs3bI7myRfLg1qCEHukNn/B/JmcIJs72q+kYWVQ1Uf6WDbkm
vFtuKKInBYHTd7h8qR6LMf0bHYHnU7G0ifinvgN+fqJx/n4L5N3QMt72vFSI
JTIiqW1wl5bs1CgcM9NMG8eEb/7aOtrLkuEOlSTrQTLyxFnUOj3PtoDGhdXs
clQD2KuE5Ho3eleXYU6nZXFq+VSZuB6uH5b/c+xiPn22vUAVgCscPot2F8vL
a6aA7JH3K4ZSvoSBDDRFb4LiKGLZhUilyPLxSoAus9jTRFqNQf1mny2FC+42
ws7NxC8hnq+8ayWcU6nC5yioZebVACL4/+3pqLCKeiBGGnnztjAfKHsRnG/u
Vr16OV5IskClIFAHhly3RJVrdocvDva/ZShAjtunq0ijhimCImf5P+Q4Uq0d
Fg6fiz1TacLG12J0wAlss/TOIHa9YIgzzSJ2JBnzYudqpf5kj+1ca6GtNZit
ftlRNeiuWt2O7YXKIgauuR/ZFIT/LLAXEoniAR5oFJnvUEVBOz9ycmPodaJz
jRm4hVthvEvqd7YQjOEa1MdHV6iiTWNsMjhUqm5CNe65UMrcj/N67vwLwPel
q89kbKg0NW+VfxwWljukXD+mczgGcNwUSFPxiP9rlXrHPG5VTRb/eCXRiZzP
JSMMFBqns5tGCiJiKOBR2CdKqiA6vycKfVLf6OKoxSsMhvB1nILXBWBDw1q5
xzcNaLR+1AIBmeFAeKlAP5lmZPzK/jEAXV7X8I1Jh+v8nw8/oQG0apAtdSSo
IrTX7opuJS1V4/w1LM9kcos5j/PgZn7bdslJuipxaNMCLQz890R6+XFPAYaM
Q7Wq4GZoGJp7aur1Qr3o+m+XyHC6KiidwbF3jV262RadY+WfTSXXbMIfI+Qp
4L/dQ7bo8JXz0w+rvEB71ps6Uvm+F9ZQEi31LkwjX66dR9KmQ6IatqLkNe7n
8kg5c6nIXlDipsL3BrrneZHdYFIWrvRkX4xlGsO8MPA7P9sXdIf1NXStrJQV
gwK+toB7KNGoC/AMciZP9HGxYG5/D31WH3qprdHD7j32jgNUcXFrgqFY1pyJ
JIhNar6FCnydSzPlWyMNwZBJIHw9q6b0axcsTqW+WmJo1NHQUpJU5lcUknTL
b+leTMxc0dcRupUQ9NvOdMMUh6ythVAOj3jLImFjw7SZJRgiEQtfAerSmrcD
pmilkVyjhvKui7bZ7yL/huHtW9FbPcxgl++P5wjlxhLNnaveBrP6YtFy/pg1
NSkeygo+PWkXsRnyS9dYImWhraw/e8iQV/WxlprbI+kk8txgCn+0Pcyc2QJr
tpDUhzicvo0N7aW7YzGfQEIQzeImLFMcrgWgdetTMe4jrtudSZiIiQbBlgdG
OXEXBKSCc+80+Y5HtJPwELi6vquxb9GD5s434ysvydlrV9PNgWiAGwm7gduY
ebi2AshoBYUn9B+jYmm3UQA7K6GozkVwZDc8uDKpnmU+fSqS/Y/fisyoA214
VuyIaa89RQ02ijVdQgp69irtyOa/Qbeq9VspTx+gx8bBXrAPrPg5ayZStvkC
wE5rVhv2ITSZ8K5qzSVg2Z2Fkj2K3b9PE7kTQfegfIWka4zhOA0SYwepIYgS
HM420tMVfaxU3cA5issT9Cu+Pq9WHnF0V2ELivm1rP2DNwqhiFQwg7PAdP6L
+4D8aEd0Zz/sV5fXTuj0+NzG9m/1c9Fkn0ILclyvX+rk9nSlK0bYj1tOTrfA
bArsOI0F/WPVHeRcWSTmdjd0YGY/+j8p+2OwbSIwE24Igh2Q1BsgG6/aw3KW
1lYfqmtokc9v4GHPmgYe0rsNUtUoWJZ2nl2k1PYaA9QQpnBi+gro8dTAocrv
LjcVbrB74FsgAxBe+KvNfrSQTsafSFLSq1JXS1GmbTRXYphdIKmpskw04t6X
BbkqSijaU/HpG5dDzqkWZ5Vv+WirLqTuSqZLxrLyNch/aB3mB6u19CmHv9ek
C4W2e42hGHfHBTdIT+7V8bxba1zxGTqDu6aLUau9sfNmJ8F/Ke/BCCMtxf/m
1okScfRWDR2hjQMKy3m3a6JYA3i6iI9tApVrVqarX4lqOwJfCcVqrkWUhkUW
uws5wQoOxLevc5fug9OkSCbCWglMF1bIoTSBVphGW2EwPgcugsWRx6JIhC+S
k1tFSFpopuwZJdeT/pAYh+IDp9Ni4KJ1iaLed1dNktjT/4eFnaYLHLgcPHGX
O+3ClIpezojzDeTzfvzHmzz3iX3UscPD2vqwxmBU3C62P1j1AAVQEWM7wLQz
uMvds09dePZT6zTeK4bRDVhSCCAAptDxFmTkJRvlM1mDiEXWfrMWsczIKaL8
nrcOPIR9vmY/YVZ2YsXdwQKzdgWSQpHCEwGNfNhZ+Uy5iLnqloe1qVNljvlp
wOLJfCrKCvlds5GIYlXDfNcEkjrwmNAKD7GvpK23LYuhAyBFvYf3qlbqGDzN
TwRkmPNHjSfxpuy9vFoLuEIMDsQC2AzJupmb5ECCDv3Pxc8LAUwTt/66HOg1
lo37XW+5huCdBenu0NnI7KGLLWKuNHuaHtnMImvj4EAFOCYry2LGNNsAmQRD
l/cZaLmSBqPgfKZ0Bizh1knOEpEdXMUXfg7lW8JNJMgzskMQDh5VBhi4qH/f
cHyOOQrx/L18C+kVVZxRET5l+dq0JnCgzUyqGhsb7EbulWYEofAf/2oA541d
JM4va8Fj7zh6PL669DcGjA/lDclOU14RzPw9qkFidaBnbRE0odHo9DJOEHQP
YqeRzPPJa6opq8k3JRcYunhWACHI3pgeRK2T+p3mQXRYLrreLVa9+6Q503Pg
k35HJqA+l1XEzTPNL29nJBaSg2xCw26qXCh21kD3Q88/DrQcX2HOJ09gfLZA
zag9m3CObL5j/2+AXrEZxCO5YODcnWRqp9EnqulgMMIpwCvG+lKRl0WNMZqy
Wy9nXylChEhzUTto8BfWB1I2YBHn/IMXGiuZtynt9+JO8EgLUFP3M78w/doX
kfetXlEIIzE5wQBQmwKuI/mgA//nSvtJGUGo7dxBnbkVqwPN1AJ/rI5i7/Zi
QN46OmjgUkcLFtvV+IJFf4NweyhUKvF+XEp4AWbRKL0HLJhcrEyr7cAcugfr
1zYSNukFiqytlo3iHeBupg7bDspczRXDLLTmLopFw0/+F9eJ0tIcoLCihWWD
dmqRh+ODvjsxnK4BNe75P6kV4C5BvUjFFaOaqSEwocBv4a1l65VoIFUHrXT2
7Ea2MofVfxhW7IebTvGUuVNRUYJ/sZl0PifIqYTpikFZSWA3eNsDWHfsYXL8
KFMhrTOf8jG+ECYFK8LdjY8nMsIrJeynp/rvxBNYvp8kNo5y2EFAZgORbUJm
s9h8yJEJiyeJ+x2XMPRmfyhD2Bg5G6RgM5QjmWTO5PrAfdnhGVzRKzCT6yUk
L/UjArhUesjEq+Z1foak5dU2JS1kiHyDrFCOdKRdJ1Txe8w2BcQ5GHqNnGFr
ROyjj7RnJzFYHpdnMSu5ao9CU/bFSWvI0jXRpHidq81SnLs3d7n2ZN+VqXCy
2NxJH3GO0uAlN3E8VwAWFZFM6XDmU2bwA+kU6ERcUidpDqgAZYK/FtU9g+mm
eMaZezciXb1HSrQZMV18gUrBLtnO4J59WJ9dc9TydwNiUbwz1DYtmxxbAtLe
6LPKKi9cVgplno/DVBGPYoCtAkmqIsrnqyql2AsS0Xdb6FqbHkI5jIGZAgSx
XoQOEjgfz5ZWSCyILAvZ1uBg/msDdZabv02u8U13j2MouYpaQrCJpRyBrqpw
sO9YUlq4v3TrW2nfGbc+hvxsqca3QuaRV9Z+N98MlhUtGvYLPW8/IBxki7pO
elo/ubgI0pNfOkBAnQoHsch+2SCqSGlSfOGB3WACpnNwg/7xjcIyVYlJDNfv
oHM3LQQjWa4AJ/cGqVAVdBgM8J0kyvX1ArrgIdGcVYoXqpAbtTtX9CkfmcJN
8uT6BosOh2H0dN77hj1a25VQavMnTyiPNOpB3aMdSROaJ+crNAOLMmEHGYxk
SA6z2ir0TkJatUax+1KtzxjZ+OVRND41QYIi05V3/2v2rNVig0QIVbZ1Iqel
qodNzQqhSfzP+ohgEKcvE1JXWtJ6qM5FUCMQDdkqYtwgwBb0t119HVWQXHuZ
bNGBwArd0+KbZ6IL5tyy12ce6t1PsVnimJucvzAr9FmX+S46Dl/I8LOI1p0z
rz4o8MtBxQbmTkADpMZCOvrg3Covt+Mc674gsV6O7V/lAfrIcdmD9rWcayvR
5k1mcdEMrgyUOQXAy2khse0SHeV04byLX9uGSALB90lO+Fh7Ro1j73/TK1q2
WM4ZX/pQBxDKqgyZmmtBWL4zxDts8jEoxf4gMYigJ4813JDzAhZ414gD7Eqh
s9PW/XIresA82lx32QREYLvjGt6zWKFLoclgUxNZb1JlPkzggjjTPOs2HqQ0
ST9/0flrmA+oK9tAqAbkBM9FZvHaVIwmNKcqu6gXMlnYZHSdTG4r1mpdbwS8
6mzeyfY8qd7QCzKlAutBLRLySyot44suujSTvvB88/H577Y1VZcsWy/VrVyc
L6GOonpY7wGCau9mf4qzehjY/noBgJKbHHHNf6MLJZl2u3c1mFj5SwcM0MDj
aK7r4jgQfRkpv5tg4GsriD2E5RaqcKvblB4U5fF8zKtdteBKv+mKcXO+25Aw
to4PH8Cs6i/M1pkpuaxgfg58pCfFo1BrT6RDRwpw69+9+tWeovOvUC2TAXyG
rWlsciT4aYclVz/mYDMRQOD7vUAB7VXme2SPcctILNu+sNJIRFRang1K4Mgp
V9rculHd6HIs8RETQ79IcpxxhP4UrWktayBgQlS80meGGUarPC5FZEw2Vlqy
udwFPkP3SODE5RPNPRU6AYdUX0Kz0iAV2d1tmS92zbbe9/LnBY9rotlUbGXH
QLJXMTsecOeMmw2E9Zt7dKp/GbiqK893Blq8HM66kaO5ZjwcXFHq8yiWML7h
z4d5dpIkJFVUHw+rEMkQ5oPwywK4rraSRpkYP0eYxjNWAqCOi/v7ArF0UEiC
U6/oAeymipiejpCrW2rpuf1al4ngm/nZyrC3PG7xrj38kxjcfDGdnJPDiXXi
ZyJscqc2Maf5qk1nV62FNQVMVYwnERsv4wDuXfKrMZmpNmBNGGzM3Xm0qVU1
vmE2TBQzbwZ3xho8NT95HAY7dQfpnm1cT4wOl2CFC0YEDX8YwKmElxHJN1Be
TDMGOz5RumBR8Lk657MuMP75CQHsN5zQwGw82FO9VIja45Ng3RZxJ1WXGRMY
WWjL4fvEUlxlXoAD7ljCJVKvwvn6RBkFWdsoT7icTJS+NDNAcjwuKfE5J8sQ
NalWJAqkYaJ60r0pSFnYocgAa7FDiXptVzkqXwieZOuGW8wV8e84uZy/v75X
Fq7Ey0vsA5aY/9xpWdYC8pbMJDUZAHkTUDne76fRSrOy0J4H+/zx6ypcrKuc
jNQXDJw0WObFU5EzK+rRnzf6YKAZ+32Op3jAouWChHlcN83N2q+sgGe8Evy8
8dfwKEVz/pY3B9QD2mUdB7AVwIYu+HvXxsoeWly/RSf4vb2E5CX3DEqmha8C
tIrONaMg9aE+r0vXOf7HoyeCmzUKEBQBSPbrR2ztrEIwjIlUk8eNan2fyHNM
IHS7JDwCFSAPjvNMmCFgID8GxflGjYhu6wZNvyUpLb1lQBzfAeoNxwEPOb5o
cKeOj+pnWTu/sqiaK4VxBCYT0nlex3OzilX6FKbv9emG8NTNOmA2HtKrGH8j
BwyITa4r8IvofqWXubR7ZN+Ams0d5uxW4PtBQsq2m82nsRsIk3dtg6kkllcz
hcqv5yD/UKklVRAGwgTrbhohg4/AsF6bgYheV4ZeBaeoPVlngjBta16CW08r
L3n8wvfvnJ8U5YF3axatKSPBfYse4lj/gIokEPJa+hin/8vCL++Qg7DFlaO6
poMcaXD+iwDmieL1oHFZFeT5ynEQ2JrkutUp4lvzxxjvfV9EBe1NDEzlTm2j
kXj0HuyPZynIGUA3e6wDFqLo9qNprl44TqtbQ+9uG4qf/SZ5h5fDlcLcy/Me
rlWlyxt59YAY88d7z52M8Oji6bueE5Y6ay4jve0g7qZ8CHiYTig7kRZv1Ifq
Msg82FFYYEGL2TNZ9trzdm81i76LF9avbfmOC+3dgI4BMonS/qM6ixRvd2c3
Zhbk+8S11wSIMVGGwISU/HjSQoEJi42W4Flu/JQozCNKP5AT5qUvDzTWssTO
7xB7SNGLAR/5c1W7wLxGg3W/+MMJueH/+rkBZSIGtpxnc6eg094Sha3bD7Zi
9th87Psyh1ApTJRUQlIfej89cogR/zAorcUOoy8t0Aau4pYpntHErQVUmsah
N9LhWXVVkoQkHC2kDGZ2Mvl2JebwMyhqsH+4OWIKFdFliFnxsqQpbZRW7B1q
9Dl/mEDILBvOZBQw49e1V4irbM/qPjWPU7Us44X0mMqR1ICIezhBepXOXYlR
s0l2arNnasS38Ah7oAm34nUSG+wvoyL1tZPgXhwCTbX8OKAP3s2bX3d7XFXM
KlwG3IRzw+PORU18ccI05PSFRoqPB2sQU0lrQszMK5qmRKUq3mk+MhH91jHV
CnZQCrLZJiCbGMXxHk/2yB4Yd87M6bH0Odp51SJcbZdnj2XsvHfshVwuidE5
wzgLIkvkEEQvqyrlpiRlCvrqAaPLkdLvjs5mopL2PSJrockllNvGBRflligl
HMtWX1gJj/PhoN6G+rTdVloy390Dzr1FXe9tvcqtXlwLZ/EWhxZ9LK0W/2Gq
JyNa7bRTP4A+OXlHiyrkdVuxXqUyAVbjxComKan05VIDvw0DH84c8FL0AwD+
XPn5B5L01CS9wIx3tevisZCveruGjTJ3KW6ruFV5wO0Xf/vKoIBNJuUIU6dl
F9LfuGIR9G90PJsjyTead8pSdXodVJkhrRfNKF1kUbXyS+jaerO721RBpLyM
RFU5dMe0jaTKTsu9ejYg46RYXHYXcVPEMX981bPt/lneZb5v2DdCjgyhCz1E
RVnfz1OQ9CBwbJ2uR2/zz+2ryM69Tq7qmMUlpG5FzGUoOR9dbYOJ+Js6I5tf
eycA9N932VIkutT/goDFuNkkFY34rxcOCqyxmlil0lPsTq9hY1gBQvbR7VaB
XpnOkuVhZqeOJRBLERPXx2rI4Jq9WVbST3m3g/lk1Lo75JNXq/Pt8U8NB6bl
NQGI3fSXrhhrHZ53HOBzIu2ldZjWJmJNjAccneTBlZrvEsg7kXnT9DEVS1JU
TW5KPnxfZTD9FIy2rpMh6NI3xocKJAPk9kXRAwqBwKrP6ph13YBuuwjAABHy
2+/Ii1KyjVtOSNAxrd5ncQiaEyX+y/YyJhCgdnfr2RdOOewzyXwAKkNz2/6w
MxeWoAe2QnkOxuwkZiKER7heuBSnJ6P+/oe45o1zjffcmXH7J6t1FL+bVgIM
aO/fgITl8sGHjme3ifqPfTIi9WW0ZEcc0TgpfUafy+BgVn4rhbgaqtvHMJNz
pR8CClvjTPpzV1t82wbbIl8VBUKJ745J5YvnbJfqDy/ihga1r5WnEN9jNlZS
WvrL0OiNP8r0TsRMq8eSpObm5rDfleCLpo7D8yHMDmA5ZvF3iNQ4x/IXLYWw
he+tU4VIXlPOL6cixr1PYrUPXt15d5Nj+0zHDsnAWf0E3g3tMvPJfnd8g4ZI
NJHLGuChpaTVoIGUOgB0aebS+sK7mKwN7gaQxD2UF/R/2Au5tE8C/yGJlglu
Cmc46Q8Lbn9IIvRNSw1GkaN93d5oWEFll4p1L9zlyU5tWQKIyrIfGjYK+W46
Vi2nZKbOm51ih1+U1PGTkeWw7ry41EJCpqjLNi1jRqgAEjIdT4GU7FjcYC/U
sU6D96Kebw4bL3FfaAG84oKxgIPW/P/yWvvN7+ISYQozD6+YYOzO3duOVO5X
p48oPQTTgrsaeizKgI1aHEyxPYmfOrjd8lrz3UVRm/FDzZCBGOzgzrwXrA7H
TumITPK2tayyek55sAE9YuQcU+CvxdQUkTb3O+Rw94vBs5K2aHLAt7a4NJOG
H1s/n71gGHZbiN6YbatfMVt3wz+CBQtoM7UZkgUOpU0r3zgWkf8NrXI7D+x+
/1NaZHmCy1vGU/H+Y066+RFXuD/9TcRhsw0pau+vWKqowG/avLb4Dzw1HvaQ
lnqhQ1HHTzJIfOzK7gYzzTdEpM1DXRevr0p+P/FUXD6LJpmpvpi9DrATexKj
V5uskjsvg4YXgl23oOXv0ZkVKsPKZH8G7MesVUKS443R/ONTu2443ZYuBkpt
LCf2FNfwbZWtd7C3SNluqVlZpCBsNADYwicEC7nkUHk0euzPFiWL4Mpl4Ho6
X+XfocQHgZ91y41qNcYQidzS5J4OOeHl14Ot+Uk8IG8tqPDtVOVI5gFiiKOA
yZjxM4YJ+3ull6HkROqrrhOdud8BHSmzmsge+BsMBa04OaHhyssmuidolwwl
iohF6avSgk2gwtiO87NndkCuKynfhMr99oJJwVJ+GKXJ6UY4S2AlgEK+GjaP
hfdOFwowIlSYp5nmjkCPHgb6VKfk5NZ0aC+VjC3C4IhNPOyKhz2lLgRzDfVP
bXv7/MHvgbgEnDT306Fw681FC2s48Z1c/+waSN4I8vXQCjTIRWjjHaw83T1R
4WqE3gt1qMQkOguc+8tXI1Ma3Zf8m3A1DVRHqIBWBmpTpW5FmyyWnebfxkRL
pemNGqhZYilWg52i21tq2skWCJLOyS2o6EdNjLQeF9Ak+1J3pnmLfDXiJm/b
+w0g6XmDj1VPnVLBdLewNs/M9qZOIHBVW0cwocJpCw9lccuKQVs1afbKorJs
u6DaztfGJK/Q/ZQEFaMIUsE3YOUx4Bv/nBUV4OXjV6wjUmvMiHPA5QgCPnd8
EbF7XuGnbVGiYQJU73u/PbLLIhWSrtqVi9GJVGpvU0X3CMouL0Msco7j3Ahp
8XHVVryz/oYe0v4n2hgmGlBQm+ysBA0nJAv8Q822Ns2k+azA1JnOPgOh4utx
diP4RPkmSRhVMJrltgcqbpmXRc4EcPUWIjbWywJVZU6Krd9P4AFpS7XT1jDn
+2q0cScV7+V4RzswMVY4de1iwazGrClWQEUF33OgTDsAVHe+LvwTvgrAsFyY
3y8cGZut7V1s1CNCdAWXiOT3i7UMAejCi1frvtvWCgCxBIjWKZWElu0m8C0B
0LT5O9jXyOAEI/TEAA+Y1cG0qJnx0svH6ToncloGcNfZqmVeeQ0QNRIRYEr+
aORzL1vyMzVL2X4eKwslI2nRqcSmi7c1PgIQvWXsD37piQJZdo4WvwjP1eYr
42Vh4uuxQKPWlbhcJ8qtWKDF3vs2dOKOQfusqXO31Ic4Y4UeJxLe5LxEkvl3
usxTrTw1tBUFyPC3o3P4d2CZAD2HJFVi3C9gBdsBYcXTRJqjn5WbVbufM34E
oyRz/4htL5M0LlpfFVgQ9UgB+b5sRfMYqsxzCGpLsf451Hq/xFcI49u6FkKe
Xr5xVE8Nje8j7+IbXN5dy3/AM81sL68+h+xpYfqubfv7cLD1Gzf1LKCK2yi5
ya8Dno+iucpfzr5nI0PCw3JAKmTosV4d0W+ajVIXiijJXaldUwIiK1WHPcVJ
c6O4fW9VmKyXbSjxabl0h+x1HkuDCCLOOjppuWNXHnGPHwIJVruXoOj1Epoi
PmhBE+bK4yxwfALIuawevUNQ+LQtj4IscYuQutJORE7ARVb+WavfwhfvubJp
/5ALgkzTO38Smer61XTdQE/+hNWELfL/1ApmDkcPVvOSJfWwpCRKdKiYjCBl
wqexMxVY2Ycea7KnzS0V03eVJAtFFZDe1Iy1stMDWuT+ne1dnpvTC6DIXwWG
S2qPafwvQs/Ih/QGqtyAmbmVyTEUSO+iIUhXjDZoluIIdNhQyiHTxNPwFfW0
lcs3QDmWy7fKCRk1AnQYwgpn7KTibJW4HeJopYlUkO65qXUiHIK1blwbk3NO
U42qZmPPY17OnyW/gW++bMguJ2HAu5EU4ViHbbtABr72IJTXHnn4hd+CkLnH
zJqZEOFa820PENUeHPK6D6atBLbidtYw6835wfFFpNeqt+MtIbFH92lMupcn
tuWTrQ+8MW1dbEZx7DJbojvwfztR/BjZWh6gqg7s+OHxPCgjNbKCPciej2VH
FkgMD/MSVnbmhIrD3xTjc09jNep+wJ+F1TSAJvWRhx64O//m0KlpXu9ahgQA
eTjtPOCH9r1d3WVHMHlEr3D5xrx5lyt1OfH7imU2U1NkZNOztq8pKNtwC4ZJ
dW8227gMQlMYxHZzs+4mCSNB8u1v0FAq+mBVdYk+XJYPgYK1qlxp3yx2S7KP
9/02CnuqY8EkTkPYGgL4i3jgVpGixE8TievxxWl76QhpmcNIG7PZCeLOJEYN
UJFLZwitcCV1LpMg7O22aeWY8xoF1MCTMPzlEn5OT9XEZ4vBycU9AOp/O4wJ
ATzV46PNxRciK7D+S0OQVr8Vxitb+a+gEA38CWj1zylaViUFk7TzBuMYtWp8
zOHOeJyFY+ByoHT6yaiue7jRvLIF5dOOepv9WBvesF+xgZMCEwARbhb210Ng
UY1v60jZcb2F+LVBvVhk8encRxpRq7h7lv/BfrxqsOmjpKua3fQIZaOjkdJe
Spnn1QFjsNOUcgCm5XvvT45kbYBW0jjoADUKBoxR35Fpi2M6LmivD2Z4nH+0
z7qVVroH7KOFAKB2AlntEb75NtDRwtUELFXsplWyfjJYWMPYZvLCdjkV2h0o
hhffIWzM/oiQTa05rhTNDB+3/IecoUxJ92m0HG4S5UPGNjxg/8kn0xx/w80t
H221p4UYoakdmT9EXEm0GpD9MwDSzv7lq0ecuyBLfrjdSl986omV8n/Um7GQ
200+lFX/fzl/026WzFyxuT3EAbxnv3JMjd+dlcbuyiR+w8xla4SdwKjJfPaV
yDG2Hhq5jlHNGvy3oL+PqBKydZVjpHIs7QX08jav8jGnpDNG4NXhg1e43689
PySB3hErUVNPLSMzimiyWLj4xfq70g99Q4OtTbRy8/5zj3Co5icUIYsCrwCf
w6qo7wQGysB4U0kp6Q4u2lWPzi8ctw0GlzQxmi7tkcNklaVZ24iLMJDXFK0P
X/yx1KT3wtRg1j/Qynnh5V9R2UMJfpPOJ7xw9LOq36X3LhUysR1919wJu7NU
CmDZ2aHr6ak2FpvEWCCOm2qJ2Y6qmKrSieAo9K4S9hymblDylEFIQq9hLhTA
HyyyJQ2Sq2meckBDXLJMZELiV+ghmLXH4nSf96pD02l0HXWfKx1k1a66tQfL
CvCpd0c32jDmTTc2MlUEVmU7OdwhjIttcNRwZTWVSTRGmljAY6ky0DLH2b2d
PGxzkBe4E8mO9Wi1m+53OB/I+yuoIsp1BSeTHbvSnhjFgAZC8LeKgLLDZkjP
dxFpan8ccG74injTSPSU1o4PSFZXucr8gAopvcynvrgDSv7m1FOqV+dWejnQ
C7aIJ2r0dWpd+YyJjHKD2BXwRl2ex+o4ahkD2gDj72AzvUCx42tgc80tjrDY
7AC+BRAw0YW9ZLLYpRYsmv5YY7+jXMj4jk0OGP/r32IRjY1RSC3JQVUSJWKM
xYNB5I5veQqkDd4BvG0cwqs5nnUjW4O5hChie+hB2fOppRibarekvKTXsgOb
OED56ASHnJ8q8c+aiTDJFxa0lC/FFMDdqUt7dW1GA9dixEDiryyVe8mDn+ut
uSRAJiRkgtRtOikq7+bcTu0nznfdafDnUwTGA+5scG+nmdax6qsf2iDjRy4A
beKMD3W3V1ahcSDw68V7saJgHWkHroY67ML1+O+wR9rzzkqIYW9ioxZX4Ljj
wHu//Y/zw1+E4OuSUwBpZ3FZqbvyJfP8Oi3wiQtUKYPRb75XchQzmUdzPfiO
F33i+IXiV0asjUJl6Du/rzvCqMVJC0kGuaglUr/Eqih5nZISVIOjdLDDRwu6
RCDDfSNuWVY5DUw5cvqPeIin5e0+WFwO/5jXwdIJ6sZ8RA1kIWzL60DaB4tp
7k0cUFW8dQbQaj/iPXm3nrwxjCTkvFmtdLq851cCA+naES5A6ZfujU7X1JwM
ftPSnVkFYQps1K656b3bX8y4xhrWHGiuUgy+pLO91YQ+uOBkKXyIipIBPZZt
uAE2e9rm53R1yslh9IZ5qy+SbvA9kf14Z59d062HD717d14UEIcScjzFn7qL
bD2IQiAIasQ5HInlsV81PzfshT5hh5xmGXpvEWi/YF4M6Z4XEdzuaGU75tF7
5W1eQBsUxAz+hJcmPHoaKbeusZt7wXwhoYTUb2UZILXRIg7woJOyY0S0ZHBx
3BtRncy6exTOBefvTWpamjli5V9z0mdDx77FFme067ixq+dXWU4J/olCplWr
lhHwo+gabMAimPi1+fozqpErQkd0f+7gBoLepp1XwNdELLoAGYMuaQ0w+pP8
KWM3Fxx7z79+mqIuEDEv6dyW0ijEwteSQl1KnPDyJ0yvoLX6hHAndyLbekYB
GEUNb4yYTT3fFcW/iA44UmjUQoLXwvbZRCVigpA54xV5dlj667xtpAXKDv18
hXh+RVeIr3UjZeaViJu9HpHupcID85aWJtRtf/QiJ0zr6eaKPvbR93Dihf7u
eDSEhQKE/MwbLhSKmsL51Mi65H5vuOGGisoH4fjdVWoqAtZwHermkd5phsL7
JHvvMFwqmkAXMD/l8mfkyjcErYOCI1kgfOzWwOi24dB6XSOFTzilTG6sgwt3
HXozgkCSHETmbC+WUjoIydLABJwbr55B9vm2NvF0XZ20XLqshb3xcOOM7x/n
pCFZ5eP9NVTKZ4I43jANgjWeypJN4erJ12bQoppAe4LFcaTI9ECs1Qs6jUm+
jKfJs01e513zmpUgR+v2XQ99cRRLpN0UtA7kHlvRNffL6lIL6Zdf5LVsFQR1
y4QMLQmr/eKx3S6Z1sYkkvIrW1+f6mvpkkDmTmdFvpw7UqNNK7EhbQVllbkB
L3azN+7BzySTmQgDKnXSBulpgLNH8i+IQ6+M5agonS3QRJWR7SK2ubFRWZ59
5KIOzn+1sXEc8/E8RpGVCqHne0gma+BIQrKno96PeSKtfEok+TawuzcQ+2uH
yabGPBNg52qmheW2AXbRDWoPH7tZsEpjxkUhNRujaEPXObZAAkO6tOVtwWQE
56dFYe7Mnh+MqZktAINOkXjePSGBrvytBeaFZm6C3m9nnmsKq2Nopdq2TDWj
8aN6ZqqPgJMHSqH8lsNeQee0U5zpo7FfUAgUF2Z7mdxPq5pPl9akisLMeSpr
cm6EZoP2G+4wdkY18iJBG8vHuLbmHQouXwKed23CKRrOz1Z/vGJxE3hofjx3
QS/pIQ8TOYRgGWtK9MuTZXa1AebTZ/eTBgPEAUwoBen0sSI8w2rhBDLBBUFZ
VywJ16rL+AwAgtu+i5TNmYWPBundzXfWXeJ2pniJ9ssGcZm7KyqVg13nSpWe
lR7z2F2GVoDxXbyPy9qPhslkyXMTauIIfIa17bBgyDkJWXRwwScFiGJPFdgg
EPnJdDW8EksSeA75WfrWzN5WE5ByWtLlAM/MGSko1OKatNWgCY7TpU4MpG9X
o2vN9mKdzM2lLfdUEDP8efpqnS6ipO6UAZbbAY+ayWja72YjBqkMMqg1RP2J
/sEpVPPpax+GJHdTB2jWPhtmATkrGyAWrd1d6R8+U8IuG/ltVEjtphGwGnAg
H2UJxg1OOwyc0fdYgZ9abxWT+PNLoSVile9z39hkIcDak6v0CB2tob0LbQsN
nJJbmOmpavae1Mp/lM0jfgJN57TPupfKpxHWihIAb6/oJhB/l3CcpQ2OizaM
bV46ONbQs9PzPjJwTycV70pTfmCFsSWm96IbtgwcfZv1bHeBh9jojeunD7qc
CtqBPb04o2kLYihwRwr+fQzxEmUv5zHdIiWbmYXIbyR7XjviNwI1L7kNacTa
ET3x1iACAor464dAiL3/Z/wnbyoMidhD3lQ/9msuvGhQulFHarYqcXMIlrDG
s1MuZ6u15cfpFXcBdsyu/fWFZVh/PaLWccsUKX0WSpzErWe9JuvRPjC0wKZX
Eh/EC+QAyZGEYtYxmBJ+4LvnyU7T4h2iOe50u3vjDcUQv+hVp7r2aScjDJsx
Idig8qrzcIOFH42g94JbMTvuVRRlBRo252rl27gzPOcJ03xo/mN2KC9qJzKF
HYcNhNZM3S4KJnDKrnYOFURk2TcbHEFxG+ZPFauEC233MDSyX/BH5cE5pOsg
6Wzpvd7/JlCZAYaeqP9Jb+U7dR3pfSj9WatOl0/KP6PR7aTiBsfxHDVXjPr9
/EP6d0quU62zkZoO/JyvcrcOP3RU0fe7ekgYWB88MemZlLMCLvIAbaVFg617
k9Nbs/iu9crfIsFG0KvsJYlNgkREYofT/7epC3rIlQydKklQVbh5KqgO48Tk
3xH/KBbsdSms1tK0ZN78Adkg7P+1V5DPRfqyNrcdIIIQJf6wqUyPksbqWuEt
FRYERZdPC3bcmmWmTIPZ/M2aRCfyqazdnGzCS8sN5gGHX9Ae3YJQ5SBtLcPk
fZv8NcRSeFs/KfohawtdsqN0hCY0MyrZkXcNSvhJJGSNGV1abwqr92IkszgQ
b+HmgHoa23DrboZ7Y0fQq8XR8GvEI3nF6JV2e5nvqmC2kWYRV1pzRejkT3j+
6Ea5akCVSsNpMfuqoPHOSUM2SWk8a1i73+55xVWgs9+90xmx1WgyRHviknV5
JtXjjWGX/QrbsOsiGE/1xpB5EE1nywdmafoKWxxv+fuKUPBpUi0JFSdGnbUO
capDleQQ2DwDMNfwg61s0EW2myFV8UW/Gft6YR9J2u56wq7vMNzPMMfpXBIr
fBKM1SLuX3+UhJJvnhOsPQf0QgC7HIvAtLTxGek+P8dDlPjkw+VoMPn9ljgW
zFs22Rf04xbC367dpCISqQH6fxWg1ld45rOoqcz1rUM9dRR+bXkRQcThTohK
Uwk8Na3IleLGaQir3iWdCnb/6doNRDJkqvuNlnYMHRv52GR7jjmgsInezoP5
Nj6DJOd6ocAw9YZ5lZn5Tp4TWISRHXgug94D6VB+qJjM5Tef6CjdMM4kVYZW
YlI6285gdLzj3blWto8R0oEsMmp2RXdwoglbpRVt2m476xrjZQtOEDDvvuyA
C/xJgHuthBHAW6vYvPZXvhfeQ2k6uwjoKjzqB3GDjTFD64NBrHnvPBPWdRJ+
leTw6rlEj7S7oI4R6s+n3A9xmSt0mHDWLRi0ui4NqGmpjf3eMyVqjGcprqpf
9Qf8zNNx9HwuegRwVIxzUaTiceEQpeYvvBVqO+AotclrmWVm3ci6PUemA4HY
FWKSMG/6rjPbou2bT/DDELc7HnvEPUfjuXHspm6/5L9tnYW6l5xo/idVHYi+
3NEVSb9XpeqM7hJ5qe5NakvfhXlK4UTac3DczoDNIbpg/yOlmrlQLhH1v0c6
qRGn75iGXh0A3dMWXEU29bCcqbUj32wXzBLQaIDlsFGn9eQZPdOH/E55kwox
wrMThuqfLSw8ZxTplXMo10AcYxKEn99RLVQ+KzjK01yCFBwZ5YoCUsNIJ4mz
/clPYnioArLtoQJKW503nSHVQcpTrbHK47Jjj1I0m8Ouz63VA+XcNTjQ3fgR
+i/j7OJ32MrOr1tztw/i70Oj1GqsaGs/aQTgk7rv13JpaDH6MP7GIcajh6IZ
PtKtBzt8IvuKgidPOEOOPSaOV9lxSHDu5+rDnXVcFY/iUMBYjQn9TolhkUdg
bU14aQQx9Hp5+eRv+vZ8i3Imyi046CZT7w6ErNA20Ie15gaz1NnMi/dy7AfN
nnubzIrUe6yh+ghDMlf6c5JXYhrx6xQY8B1xOoW7CeSpsBxZaMgBI3VNVoS3
9ZHWAAnsAhc3im9UVbDBXE6YDPQ0Ba7swT6gajtXegN0jAY5zfOPHwWCHYeN
9Fm/6XF9Hw+CT9IXx/0ayu+G+amgAmI4btFP3oTDRhReLqAxn5Nsgbe5Q6V3
fPJ2tuhzmQQEKWslWKcdDTkUS/hDTeq190SZFCYsAdHYeUdBSqjxCnt+RNne
6kvdy31UsNDywViJ9ZNqbYubgLoL1purtMeZFoled7bF/kVMcq+XpEpOEPNG
0p9Os/c7/27A9CpLpH804LpY//hj4NiKE+TMaht7LwUHeTHZsJQBPn637E6l
iCpeMs5ycHAxj2d4n1Z7S4G13xsuNmxllZ7jlRi6VNjQZCQALlHfBKnwgmTS
5xXQ8V+RNbUKp70HvP8Oi3FoRArNONcPfqtRcjQFHmjnnpF5HOfz1wpeSUZk
Cu+lIXPF2++AYiOfm4uFBsCUB/l8hTNXz+rA1l5C71Dy0JegIImb9h25s7pK
gnvFhBZlGP+CZhkuMYU2cYRceHu1IJbOYyytVRWwN/6PC4jZ8ecu6EtWkxG9
1a5wIQT04W6w8uftum0JPOfi+ZxGmLL8p5JJjfMe9tkBA8+b9GWS5YK/d+co
vcJakIRITTcoJw0lvOQnghYeSMZPyAO7GO2UGAmllCry+Lj6X0YBLzi/x7Y7
j4HyIKyV+uosCQqr+wSO+4j1TATQU24kLd4Mjl8Iih+/UiF/Vnthl7V2cebf
kwGearUnsvo6+WKpY6za5/JSub15bu0UWnUR+ILDjBAf2fY3hZCIeIEIwLXw
9eUglV8Qrj0CIeC364yOtyrTjasQ2/Az9Kj9KS3k+kMvGz407Mpc91fW/gLe
DK/G2baOKf/l3pR7AjV+sTEZcRTYvOFLyyTo3EB94YJaWoRewMHqitsms1Jz
y1yw/d+GX5HZ+3hgFerezkwNQxmaX27tQOUa3riYDXFXWG0At4xX5Q02f0xA
KgagsTf1VBqYkFJQfVj7IleEMVGE9rEaW8cy3d2QzXtygz7ncRee+vWqtg8R
baB5DAzTFz2XgerSkmvgCWE/3DkWKRMhjwXbOK1H8g8Z1vreVFmV1/EWAhyF
9pb1GMYFcsZjKzcusI/+OKFz/ITHmGtFQDxgUDJfifONHLnwCWjMJbePbUg4
gonVFLhCkv9xfmRXna7zmiRY2yT+LGcJPK5sXL22oy/f/j1s/Ll6Z8ZK8IiY
UBjdi0rT6IVY+e6Ql0rxsApFfK9FsB1Gwlui0clfLTBeQU8WtE3dFz3K41wD
OFdOAhEWoFVCedtyRo3MS83fbKIk7ye0EFSSVe++DmYz3wIBTwFH69UoWYVs
Lx+CDf/yVHhuJaBukSxvMoAPmkVb/ESTUKWIkH4evD/rUywchrhNtFIL1Mbr
5xHPU/NMmxWnuzvRACrSRJKTGKnEv6DHdewJ3lnOxbYgzFey6sgLFizh2OKd
C1YvyYoF39+v+d2BOYUxgchS9oG5hN7xhYNl3M9x6TdBejn13VanmUmc4RuE
BJaRotW3udDRQt5pCZcls2tuN6xJ29+rNBXnyanF2eQZZFp/6hXVbRv4p/iF
+iV8iKqIWDGVNYyQ0syFWpZ0374P583Fot4CGSFKwxA86sKvpuwsSNGHIFT3
lrqHk7c1/qDH0kGreZk28GioVvnSpxDh/aD1/kSZzRNmYkc5m8kgsSjIZ6Yg
opPG0G8016ngaLUhC0OImIJA+JYQLz3NfOqglVhdOfMAOJs8+LbRIxOkeUej
bKTmDPKMDXx1ZXAq9Zb8aFR0ld4zqxCRMW6AlbhgF5darP4puSn5TlCpJKKP
f69hiu1urpAbCvTO+/N2RMibGmVLqBc50ioBww4EgDxrxrMr+Ey07Q2nrrvk
8hYrrgP9W1HqAZibeV5rl+qn/0NF5U9hfC0NxlDCYgDvneGwzieTzlcb6eQ8
z3nXAPR4vQrJKEU0WVYmZ0zuJkaIrhx/ZG8DpXixazaG4W0Umqu809gP7fAv
FXahGzPVFoeNT6r+KHeCKM2KMIm7dCdL7tdx+S3uvixMuYOSoHEciHpyNPAd
DP6j7j+TTYkDqwsE9stUwsc3d7McYvoQ6DMPn2Vs7DKkktyUhCLmxiY334kX
rwcimX1jIRIahaI40L9D52O6npRj1JhmkZnBrnW/o/WD/WlQyELy8r9+Xecg
HqX+e5nm+1vQKv+m2MOAR4mce0elai2OqfTxTQCzghe/faFbyV0ssPyK0UMz
rsx1CA26N7twGuUIQS5rpExWdz+ngJIEohT+ggvNnJ1Gc407NNZkFlLWHA+z
oezjlMgjDNk02sC22GT7WkF8NtneGNlLC0/B4pnkQQFTscUX45OA8ZjrhB/G
XSpRRPeryALkyFojdcmhXHEcC3tFuFZWdqILBRCtha2Ra9/49Es0tAoQCKAD
/Xr6O1H2rOcTB20vTJs2vxltdMic0wWwJffByYNv/lN9AflCyMte8j1SWT4t
lqf0cjwsWo4pfbEzODW4NhAqUIneFlZ9PNbjDKraav9tuPlXBn1hzCK/Jj+p
6EoxGj4kk7L2Je66Aa9sLR2VcnhtJoJaQCGlvFtI3rLx8zs7brniDegCsKrp
BtoP/tctaUFtBrw67sK5goKLfxzEU/G/FsgkWpDnkQ2dF0uJxfg5dwLKLm7S
PAscUdahmxP3+Pw3uDPjNMiFF8VC+G4qTsCW6otjCnFe4tv0jKiPVAXlABIO
LZi70NlRvb3+i3FP97kF+Hm5VsC30ZYH1RAQgKByl76fTWGo54UqpgevJoUs
uA94NglAIYuFXw/keV4twNo3YUpVFLy36WK9dgk6ZxNjZ9HOpfUlDm2+AicX
NAyRsx1LHajFdd3VIFUYSGEAZQFdy2h7nFiqyZv6DSgwGkQOMbnd0efsJIYd
sZ+PN5Qi1igt8C16sogPxL8gxyAS+9ShJCircf5jq82eI5h9QxqIIz/Xf+I1
MqiXnuslx/nANRvc1aASzQxKP1bLA1LCOHH6dBjM0NCi3amZRgKgSnpcJl6Y
PRBgu21eULE7CzKOq7vJHmv3sxIV8LyZzSWPhX1m29IwJYoD0MkECSVscwI5
VcUmBK6/gl+sr/R/McDeon+O86HgJji0zj3N3OzBeUy2JzybWcJnCFAj/0Js
oQljN02bF0kDSbXWJy+szya026ZU1bSDaDqGEdWNYUhfssU+aajr5icshl06
AVMqJdUv3C0qp/Jr8EMQvKXkixxfE45GHHAu28Ch3HPSmVftbcAF2sopjRdI
H2U0LHsVLQMsw0SN2mRE0mXKG4Jud4OQ+jLrYD6gTaUsXlqNmGJxJPD5T17n
ScpQ0vL6dMNVH/BQjPjxLuMj+JRMVJPuRUDJaxvJCVNIVU0IiwW685sudKdb
d4HPoRqqsZYDm33PYQ14SdNDftJ/lUPPDNX10CrtvDzGgvqGfcb+bAqyFaxO
xBA3ul8nkaOft7L2iE7A8sdtIAUsoW7ylS2Zszf1K1OOm/0k3++Sdri+RUX9
8hcXwYnHdT1jGt4vw6tSMLbAZpkESZDgR77ZOhJTjpca3qpFsvWOqgfA1Byi
IEamk2eNdzLz4+T3r82CVxc3iHBwhlYqjc1+Kv18SNpxgk6QzQKhPrHSFObe
yIOG3Xys2MqcpZaUJOyCHxBTM/RkzTSbnFhc7lC1oMb7mUZeuJkULfAU3RcY
JBMTOP7NgBO6ZptkquuEU0p5nT9qrdU7Bm+56Q/CxNsEaqK1ROyCCRUssZ/T
6Xe2KLXwpNfFErE7eTQ9BikZs6BON1Wj0tia37knvNlKngQdi+sFJjf8IZK1
4hAk+2zwDFZz88gc1vBs45dhRRLzjA19h3Gqok+Qz4XcC7SIdbIim7O+dm50
oyhMPVZdF9YXow6UZDahbsNprrI0OghRBnh3NCSUoAN8aJ4E9raccHKFr7Ae
VnvsEYUkCx3l2ce0g1J3zDOxQILIwV7IAYyQBkoxWuBP/vJS0ZQHr8EL4WRE
aoQgNn0i6Vvam7RaokLsuYCkkfyi6uphEm4HbygHnjd3Egva2z+rAwfMqvlo
4NeA/Z+Aiq2DNZSbQ9vfnnsZ1fUrM8fKxnxKT09CjsoEYzyY5rKV1tPnNo/l
MF6rfxycnqdGjJguZjKfelzz6++OYMGOwmy1oab4kcfZzr8Z4uUvJA9CRKZ9
B4dVqqi8yD3oLectkTAMMPdoVADb9ObYMmUWgFAPg4pZHx5MFQcc6M+Yy82B
lu4cYySAJQSAr4nxpwI4KRPdGDw9Ft3ZUCvIHhSZI6BEZQoJ7qvA0ifr3Bc2
1zAlPh8HxIyl/Y+LOWjCiISHJen9H3xeDTiO1XfxkrBDX4zzgQwDaIgSbtEd
02Xfn+XDqiuDHps2vshmCuymGEBJ6iNFYrN+PsHbNXaf+lFqtWu4KW53EKdL
HZFailh3f6ksEtWcPt9YORBxL4yIlqL0QpipW8TNGGuh+4MRyAMljPPddTIj
SMPYvsa83lIBtRY1H3QoKwG+IRuJgYDmSm5QSfghKDw8g2dqoY5aYlX+tCdq
yktTrSyjKdpP4qiuiaiRK1fdI2pP/zWyTvBHJYDKkfr8er3Wry4sojVcMgd1
BedVUESXiROrwFms5UDDKSXuBvg8zErefnVZ+/uwjgKiWxng+dUeVRZJ/YT3
4EjxWzrVi5Ugh6t0RSgkJh2VaIv9WK4pDXco5YlY9wiA4l38dF0MGQxUbO9y
85T547A6OfkjAVIPt44MUr1I311w7FaQFqSdGjGYupgE2AfNs0cD9/HtBhhC
SCzxUJhA4ooFGtwiLBNl7YfOx0lUdNqAMQSTHo/0x9pOQ29wZ0tnquagEqGP
Waw0kuHCsIpmfAfhDMsiRIOfJlDQaxEfF7sQ3fcz9oeaZPNatwu2/q7UA8rP
p1itI10TGRj97HX7VNwWcN1Ou8qWL8ZCIR6zJCxytGFGz+esSmyOfyyWIWbs
TudhRhglwKcuzPSBE9F2uM2knvJn3rPD8BdpygKkC7WgzcdAmfgRYeu1olqE
YGZhtmf7fCl1+PJH+REm+hAnnfQC8lSPfKJM8pcIoeiqZY2TqfGpjBWfgDn2
Ch+3JtmZiEv2mL+ogQoBQL2lOe5svOXvxJKsdBmcPzauFjMVVCIRgMYhI5oy
ju+SHDJyBBqbHvZDZxSQMQXz10TL+P7zREVVfOgdIjf2/jRSKtjq7o/2CiTr
sx0c7Pfi70QoZjVZ/mxg+AfzK5IFCcwZs4jmQ3o0C3sbUyhxPMlmoD923+WQ
8ykv5acBK1/V18B/ZOW0t3kr+HuwXQ6u3xdT+2sy2ZXORQ+UY23NFIKxW65G
qWEGRrPNhhs+xc+Nmmdboe3gi3zAg7v1VNofz73zy/Cyr5GX/G6liODhR7eg
v4nBGCUqq+SGzUETwGXyYcforjeuHgi1mxJXZNnOJBKvFiyFgAolIjmS1U+g
+JkG1vqVZUJBkBVOwriiqbwj0rBVAVCwVBfMZtabaavhYRn1YKBAEjoXGzIl
+RnvSvCPIf61kc/wLJw3cDDkCjIhJ+oogiyGD1Ym8pSv/XXUbb6qBAdxUdbp
VVrq6fIP0b83YqANfq12QS7+q9qJdStgFH7RmAXP+DGgD+4RUXujYaR5KLqn
exXVd2QL5hFeDJgqZfRTIrypzvmZU5wmdLOEVwcVYBVGNJd61yRHd+yNP7QZ
Eq+hamVKYNWIYWXQaXayzrbrXgRlRJLxddH5+f1kW79eeXVPgPzykH2urEq0
vFEJhN2/lZrCvu5N0ynkKW403Sh+0XhwrhxoYw2BpAArJJLdCf92w3qopGmG
JTBkZxLLbw1wz8ujFgs8hglNrzcoMCeEUDkNBfZxyUnYQ4tSGMd1ZW4yM5Mm
PjnrcZkLewE8T1UGKeprPqHdQmF5o2Db6N2MKaY9QqF0S8urEiLbLmmaQvrW
FVTmAzQ1lx7CeygXolkz1UPalCGz2W5pBI/o69Zsm459azeMZUbiHu0to/J/
E1Vkvgd7RAvyFPQD3RAA1cZ0yMJH0GMJOcw4yfUlZ1UDhAOHx37w7MdniZAq
i1KzRS4WRHjGATDlpdqbnUsh9nG5Vg/La312hQ55lYjt5nuFJXoQBIhwHzNQ
tdJsVa/Fdmh0wJZjOwyVwUr9FlU2WS/1S21Lf4od5BdNGVsdAjvqWEJmOzEs
SFOwyuzk506nI0i4+zDF9H/t5orckkJE+RKktGY6618VGLsYkFRntrvm554x
rtBO1xHtPrTNBlS6VnlnhaU/+ljMsUq4pqWUHbr7lbhXlfToAT0ApcQcgMjw
hqZYHG1ohQ38TMs1V3FbtAPeZawCcfIrMe24xmaDbPvLuAFja3DHRLPwJWPP
KvtashOoqpi5EBOKfQkfXtgrB7r8pxo0SK6R9PRROxQQEY1QFMfcs2HGEnr8
RmQU8WLceN+tx8lodNbyODFOBHEzx+7ez/fXlcA28UZmj/B3lgMFae2oAnzv
xpNTOO7jFfSIiw8V+eFVDdOd6SyFUKh6CokQjB88wCU/ibkMGjh3m1kSxTME
K/kKjoY3oHiQEHFhq+u51OclOtlAb7KXGdxfntLgBExQdGIc86W4SyCKtbPO
GT+YW6Isn+H6hrcIi4FnVCoXbnPv/sCPY2lE8amSi6DpFigjXuO46lk4pHTn
94yPnqee20oCbjLIRDVvitrRsXohJwmPwPZvcIz34BulyGZno0tLgx/JSlv+
8eJce7UiUuzrrQmebtUDiCAPZzsY7qBjU9BfEPB78f1E0cpuqHTbdmbCtvWa
9qlPL4HXe3s99b9CnFW+gbUTYqP6/fiqjerPRFXV86y7M19tPM9v0NvceTNw
oZ0WChhngG83D8PdMaxINkeYlJcvqR3meqnWuMrOCPZthX+Dv5jA2vF2E3ir
UkKdOVV6E/vDNvtRYq44x4ZYW80F+5hbETapnTQUmDrJV1lgLOoZZMPq808c
25vg8Uc6v3MK1OtvBv+qhSeDzTD8KxNuu2WBcQHdU/goLWkXJUnuNF/edN1p
/7zb9hTurNxip47hAqHJTfUciOyt1VEKXb9iNmZR2eFKW+Zp1sw/NiegriiM
JnbLYeKD4Jdmg5ExcnvKYWyTX1P/Yh+lJrHVYWBeMe+lSyJVbsPynpT33t4e
2tkAr7tHueMv3Ef3umRBfc8OlOnITLc87HTXEt9rW/mnaFteUazVtQU3RJnJ
f26/0Slll9jdaBmpAJVHOlmIrRkrcp/65Zt3T8QQs+apZ0TmH08PjtCZrhbW
cjfaytmF7FFJqgbQYCpLIYfRX8okPNUaAg4W4K38rhw7UBHItYBD0jtYnyXq
yFdn8gXa4U/luOJeT0z3ZTil+hP4XLvkUz1juCkmy82NqB12BbaKn0sOGT4o
G4BBVzJrF6wyEoI+ksQPFPWwsDzNtbdIFz5y+9taW/u+acvNqENrhV3NUqJ7
ex7LyP0chM0RjfygLWk8kfu8WPS78XTGwEGiO5y6vZqs5zOHQkVdSHeObUz1
xCEqC4ukAxLZkAgsWVJ1IOa9AcrMAoEeKjkAsJSO5nc7uVUZ8OjOfqD2MPtd
KL3dYc9q+UPbwTZqVLwn8dyNtYrwpYyff9hodpJP88qAZaRz+cqk69AUOCCS
F4vJJIJI9HBqij4v2nxPuWlF0xkB6/d38L4BzE0avYZVQ6zqfwnytlSf96Ob
ty450cpbnKSijuZcfRViJ1gHPXgWoy7/6sqb7g/1/Q0xIVSfw3k/2lGxUg35
7YriQWJb3E/vGUSzIqoysJui882EQiqcT1wMMLVc1ZhrBvdwTk9mnWFNDrZl
yC9KldexVCgQYxFu9xISuA7QAghIDqpE2uO04VnWTKsrMRCMrJcnoHaGr0HJ
lj1EA8OceUtmpggZYmXm/LuPs6vaLKgQ7yPga9ynjqhLbPzBzqQYmG/c93zB
ZC/e91JpLNgDHbsGkZpT/OiJZbA/1XwyiUkunBKd2E7Zo3O9XtZKtzwet0Zj
R/PREdJ2rczgct9m1e2Rr2Odsu65g2OddS8ai2RMJJmkNEcWhnnajBsrVmgV
CER4bCDLTA3xlYsIc2YIck3KmC2zbiy7eg9TFlrfqZ1uzIclzxBD+4pgtC7d
AiaOUw4HM1h16BcUVKsV94ZKTKykTghM7uKKNyMRGn0YNNgZThc9G8fFIJD0
HGH0VCwgvhNRiZ9ystgp0KWqlnxefTi4bsnBy6EKxDmXkBxLrD8RgeigPwKb
oACpKkBDB8cs0MFgU1zKOfYlNbr9PLcwDDFivN674rmRphHXSFgwN5d3xX5a
nqkeu+mhDitvrOzLKRfZA1YmOu4MO08LggjVL+SAWs5wMjJ3kgQ6jnXcTD3t
hmQAFjt+u9EgPhf+Ek5XKWJxsQYcae9+hvGb7LSkZBUUsx51Tp/iJ83oDWE2
EymmJlLSbdyYul57KQDxPmN5bmUbteZVCNWI+TZX6ul81a++BpTJa6Lf4Iyp
c9QBO0FENSmkeeoWky9jB0aAF7Biwo79MPKarz43z627PiXbp8gPvGNZAcRe
8eBGj2FguBBeg+Nav6GopiMpQnWlaldrC0REU2NIeiRoe9G6hcfmUddWRyGm
msI3qRbMWVF8ALM3LR+7iOZiWz0paswqsYpum+9DmuUbTekOdaKbWfJhcO3f
s0Fenq1O4DxzdB4WRLvUMe0Kj2YNg4FhOngk+kOKawgiiZ7mAW65//B1N/aH
JIIMImdHvvaPNlxLN9pfw/eney2q3rqGSd/S2kiu2BoYxhTxGudiNFZFfPDC
JGzw2YbAWFVs/Hr6soKbz/3UEZADo5TOwLZZaw+4oMmn1RylPt4vlCkRg6Hf
+ckd3irqV1nvjz+A9L27yTz7BbMKnBeByCWnAAWCkwzPDTVok7VDv0D05StM
YbcZ3nvEKbCbu5342/Sw9KztzjmCz6VbX4v6rA5287DlZR/u0CjFUrzJ2nXE
K01p370jcY/thd+QEO/bGn1cVgM7s6bn9f0ne4hCMUgia1AqO0OtZeGvihB5
tQEwX9tmaWXGaf8hclIULuABKLoIWZ7e65f1Y8p1R1O/JgZui8qxI0coUzOU
DKSr7KAwLJRRsH87H7Hqrs1GrBM2px0TZIghgQ/gE4sNObXcDeq0TvrjptQe
mJVVzh6zWObwoFkh1vrwauQKX2FFtMZ8K1JiXn0eHGpPWygD0AakU6woewl6
X/tnG3WFUk/8SkMmz/tNg7MK/Ia9tRvoonXmfMQreXkDNokkEyzH3A3RV3aa
vLUZ9//CFre1OOZB8QquPtdU+Ne2vgOvh9CubCOeD/0UT5FO8myLJ044hx+7
uaJLotxfup2ry2harOfYIzW9zCBSb2rPUWA3s7eARCB8k5nJyFXoIaXGFSzt
DFB70aiOi4Rpt5S+73BQLbadpzeDCtWeCEMa0KRZQ+Ux2rOtKybEqOIZ7DL1
R50/4f0PsAfTYBRCs3LC/+ND7RH6tZTH44h4O/gQUnu1p3+N03cof1IwEvUy
vo+q/StKdz7zi2utItcseOemkPcdymwOoCrdvUip9HK9TjhHrKYKf4UddYAj
5kXhYnRgNH+HMRyNM3FZXEtcG4dHPTQcW8LRz+6HeO5Ha7YJnDFqNiaRF2La
cQieMw+gt+Vk9oeMRj/IxJT6Q4MKE0vMMS1AXlaT5zZULcU+50hxbr7TfgJN
TbQfs2FBsaw80lIXkovdPQ/+t7rp1p70oega2j1PmI5glYz6Rs8GJsOECGDR
6jGiOrcG4PKgtOAx/ZLDhY1l++wcsB/6lusCD2IvtbuKGGPrEBo6/c+Ka595
Z9oto4unAHZZxFsBKTRrlZqXopdxXOkIIcS+AThVztPqBJaCpRKqWd/93WZ/
cKcFzvv/sFb7FEKSR6cw6DcPg8eyHQdFFHrz7PwZ4BpC4vTzb9aRjUxI/LVV
Y5ohLAdrZpfSoEfcx+gKk3BFNW4tPH7IDLLTgwylU/+4rMw2aBvVHO+Oim5C
zjUm1HgUuE9KYrE/VcwEnhDWcB93RTsHGc/LCWRB/1uuumxjhoR/U+VkoolV
WiPS4UW/qFvzk8wKYKRM7nMnB9vq3yyWbjCzdtsDqwuKWEy6b+3Rr/tgm0u2
toG5jHonGPd1naMJF4RCJ7eVGh0xhEAc5oT9Vgn3R5Tr7DuecGC8Bc5hO8Eb
fQMmQZZ6J293CC3DSQIDqYs+tCY2PRk7OEb7DOgcDRjF0mYPv3IdLj0e016o
Nt2CzVFEvP81ajfuZJG4llFaDluJZuLLLtIKa8OpwydsCEg3NydGzr/XxiUp
jy0DPtXSTzPsGI8p6N4Xtic/OOu0mnbDHt66adka/y951lRHLgoSE6G1qxKF
c25Vhq6+2tyzvzVISg3v4DO6TAz6DLjdgiTsoDyktnorxIZTRoBUp6kdXw4Z
5blsgH35+d8Q8WjQss/kMJsv+kHmOv0msihbl1dGFi8CREb0BTb8bQ3DkX/8
OE+fkhxFrZLqXjTJcRb3j1SyFtPJgtv6n19+P7D6G5q3mdWxxvvI3rviX0N/
w46bcI5WvXOf1DIP4WR9PK1i9E87cSo+s7y4rL5AUCAjsQ6rKdMgEZXahNkC
j1mlVXZTqKaYihm/8/bqCoaQa776RnZpnF5mNLomc7k5JTgJxFQJWAFj/RW+
IZjBRZW6Xe2/P9JiJVAtKpxRbaViMb8q1Pavm45UvS+TUeNkzZW70AiHof3O
lRtJpQMby21vqRUucL1XZao6nLMNM9twd49r0Fw3xPzWewlZ8uiGh8KzhcL1
DdtTyqVRmYLU1vAFul1B/Msv3Axx+DbstvYOFv3/WRhT89QcpHfW1bakcyKD
3lqgGdQtzRpr6IOzt9ZjHF/fQ0+3FQjSgDQ1NDysxa93GxiNyyZDWpziPLP+
/9VbuZVOTvUZoogbJLhCJxrduLRuZDfGMs+OzkJs1JFFRV35ie5t9ZgRnJSn
64h3tRc2KA+N6HzhBrKafWJk3x6JePAT0D5au8jQKcGVAtuyagc+Fxh87YgD
tA2RivSRsPuECQjlOQCd46yFSwjCCmF97Io22Nc25PIiuiaD/pLDOhLeppxq
NdzjjnfSb1CT5meyq0DfMwdaBcOSagQJEqEUFbrfBTuWPNfQevncWKP/FcdY
3+NxX7mPECxYW6PLfB6rka/0SH5EV2GkgO402TYsEEpxM5AWftg3kyftatCY
LdEsv+yVtdM5QhOHg4paDE3nJoMTmOj10QWoZOuhmP0ErPveoIfpxbiU17Xm
cQ+jPLhmZVZIlEuxnaJlQ2m8jY28vaKXDJ63LnkTueUURrH36HkYtejYTGhN
R/6WHCX1Y53dV89HYVP/uqxW8z+DpTaKVRzzN1M6zn+S2dW6yKXw7DQGYQfr
dOjEsemmYIk/zT0LPvA2OPI0mRPQrLcz0ZBijoTYTP6bo1JraxGftF6ugNIA
RBcJAajtoHTZPQby6PqbKjgpi0deahwU98WARfnEFFUzepCMzR+F8cKvNY4K
R2ghWpYEn93lk+n9F0xvjOHhjKr/R/TixeZ5SCvalqvxx0xTqhf2pGT0a+FC
RgT6D5ubOZ77tXfOnoTO2yuTQ77fFCkhIYY33P8blMiV/q04WWc/xDfZ+MhS
/on2AtnSOH0ntLUk2nGXrHTMRWZQYWQNSh5gO/ibEibFE3fal/fSvWbc5KkA
ZhXnD6YvgivlorZdRNcfeC/i4ISELPteTEi1Ueaq+SN6MH+v8nnEDsbkp/U8
P9Uwm1fl+1vu9SJXG/GPSBgYCUhsqAaOZWgHjGIlWcBM6Ofy6AUHQDJaFCPh
zDcDLn6Rfk/7PW7fZS3RbwF0BI+G3fRfakzVZs7Q1+oFEvUp9YGlVBLvFk0j
vNhruEV5wSJn8X7l9FjOVjyI2CzuYBs/vqdCTaWaIBjyUfVRxa2JmX9sDIie
3pFmtj3SEENIHpvztqRPBoD3lJzRipxgcmiEgKw/pUC2SHUxRrc89s42xKIX
/e3NiGwB6uxp8lb8hrZ44bmYremtM0Zh+VwRAuKfTAjHlvXA5PRNEzGi8nhj
syqKx1RV1oUOZ/rXuNRgblkbssQdpE8cO+bzGSKdM8ciR2Qc+86JEyaZu23z
Zp1ga8hFfOsYse3ljCaUwl1ivyn562/dHeJ69wq4zydxYvkQPbV/bhkAnTWT
R7hCk1/YGREOGSKVTG47ypdf6EHeRJ/TxoV3RBgN9UtCmOWoLt3sV1+zf6TU
V/tLKfuXYD/3NyGsNuRWzCqqAX2QFr+9sR2zrajIiPcJa6FYPDyg2hGc2dCT
CbDOZNKTyDO/fEf6fAUnQFYbp+LICsfbgnDztMjxvRaiTOpNRw6ehUzogdWI
sx0aNVqdEjgt+Kbf+AULhhH+VnknBW/YAbJqu7ia0GPkzEx4h3qMYke+lQH7
llNExuoOuLVi4e8jbthX3IPbZM8OwZYqu9+mU+QZ7I8J7RW6ztyay7+WEYdi
puK+D6dcpE8s8WmvzKd2BDF/OPRUrFw9EWQeV94AvIDVtc0i+kzz7j4wWdYF
5u44s4H74HeWtXZ8wKlo8p5/rD6mV+Y62gMgaDhn0wXOxv84MjA0he1dYeM6
3WFskqLlBLZ0QNam2Gxv1gnGCeoQzIuHytN/fZJBJ3MGfHCd58xnw+1tQ65g
YoEoejIXNjU+sijVeZTtxUf9vMw5UNyTIeRNiG9BsgtqmgVbC2uIYWHnN2/y
slaSewfzSmytvKU6vezAm2toXkL9ygSFoT5CcLI5tK4ApjR9wYgLr85Rrqwj
l/FA+2fAyNutyi+KJ6N80P1IeIgkPaIIoQFZqFVYf3tzGczJbTA4tBysqIdr
nvVboEK38AQ77DIPNF/8DXgwOGH8d/gp657ufT628LoiWWYuAqCF+yrM6H0+
B12Wrb4Pl/zhRb8Kg3M7r/dpj7k3vzw1T6tGJCr7FfjfQEXLGvuC/BA8tbPX
1WAXZxrGf2Q+0+x5hpHr2o3poHM25Y7KX4ZJqmVpyGx1h9tbZqNnhBcIWZ7a
kjgy9RjoprUggW2j73VvYUqI9JtlDQDHsq/MIusf2P2VeBvCRN/tucShIsHs
tEw8A5fVYR5ev+RjPqnVgVIr4VmaF6XxeoXY2C/YBXAJ9zQEsteq3Ud5ZCjz
dCZ7peeyiGt19EKQ6Q3SNusWP+C1voW3oCQ94p1jbJOKzkRPN2ahvB4VP4ZA
DcN2UW9+qzu8awCcmvHiew2W0ZUWYSN0knK5MZht7qamZPtqFvuLU0XDmWng
DAK5o0yA0l+zGKrqZ0TY32S8u+NjvsmVuAVtLTLwCO83j/Z9L127Z+iYRSW/
csjfsmt4OtJzuFZ/Qr80r4Jczxjbyf4RNsuRoJ+9pD0/PQL9tThgb57XF4wi
GstLPJtjI1y91MAfkTfy5XyM510SPB59IWA+XvqMqctj1DlzleTlVzTedZ59
YVLPgGmjl1Ou/pXmbgVxmRE1piIVEzetfYuF1FO/0s3B+CVEkfYa9sjstADO
r+qVJAqH3WCjEX/rDdL8OB32rZb0t0s6OLT3e5p7wg0MitHiW7X3Q37y0A6M
9rxLdSQbPtaMBD+nbVEqpEJLrwS79nfbL73TsYckHec5D+Y2rL9A20FFuwm1
5vDjcjPKOcFp/vyYOlReZbRYcmWAtOlJraQYe1Dqw9c5x6Ufo3Zzypg5RMmT
ior9QQARHcWt84phh1Se6co9X0l0uAM0b6lSTFwQq/XPdE9dwa68m+QBSx3g
DXW1C30lzVB7D5MZ93hp3bs1kT/z2haASi9apW0E0eo0fr3Vo1cSkum2npq3
gxKecAQtbHylVQ5tFzJ0gmpW+F9GPSjZ09QOg5oc9jezC463IQmNZQ+3OX0+
B0kYyuA641Aq3ToolaU0qC1Ve4eCGT13cgdNRIBW+Nv5nc089GLlSfJbTED/
nGwHgXTioFDruoB2FErKd0AheGPmuU9Mr84IEZAxjGrosPAs0Ud9Q09gfgP4
5vFuoofb+YxR/HUY4eQirmIdDK5whAck6a5gID5D4K9398n/qSJCKWNQqWgF
xOiMYAazHxaqwHtwWsd3VOCRwbfEVJuUZLZ6JFdpVjrI9MrYmBudvK9gZI9y
kIQMemVBhxSeXnaeTpJ+/Ta4BTxHBCErUZWOnPpxN9F2BoJGJhooNZkohJrB
d9+P7mcy7SlXPF2GI4AxGY7BTypgTO36FVnJDxhtxfegng1XEqiSEhh23DPC
ctr7amWVFKwkfdleOP6HqXZFvVRlQdMmQP1LLneaw2iHPbfUCIigmiNwxz1R
Gex3DGrTRuSFSLMKfOguPGFBRO/pmp9MUGNBKnYch8mlSFg+F0uD7AUnhB6m
sudhejOZRoY+d2EYDwbwWANdWGvbmZKuShZ5P2i5UsQ8FZtzkVfChNJ8lPfd
rJWjzi6qVWtipD6Q42vQUk1zImZHU3r3yarqVbInVy3uV6VsgcJyuXdz+EYs
UvCV/ZA8AfcrgFcoCVY35z8XeR/0SmDGo9mU/4TSoD8ZDdmW0X8kwovBBOJy
M1Axy+BC+sLVan4X+0tahQxCmqA/rFXunWqTM8vVZ1D8IqYSm+uB+tThw8mu
uSkyA5hWzdhcMJx5gIqK6osiYy+aHvH/jp/iiF7BStix69C3bw4ejVy0Ur1U
JVWgDk/OjWVTB8aPQgVX5buggp+uccAKtvAhaAxVgxv+/a3PO/NhmvQpNK2C
oIHYE5fDltqX9OA8P8NGrFNPg8gwxnybX4cX6sH22uTLvDHD3j/V3dHHK3h0
Xb0NK0XUFLc4EOUIZusHcf61lwgA4FuUrgzdC8sMY10MCvYyX5YVNilMXI4N
/oWTlXYJxzgDZyHtZ9FHaAUKwdjJ8vq3rFFRFWZ9KiUQRzJjFf39HNLwPSnH
/9Jly6KnHkf7vwAxmRFHOR9kTcMKD6YvO8fL4YQATOIzFKGp/Fjpya3goKsr
r9cp5LYHVvhKueQu6/Jj6WUl6sOOwHPiy6Y8ahlDfTTvobIaKgAcmJgHZB1O
171uduzcGOmvkVc4VEdCnFVXxIkFzwkZo/dAHR1aoNf8WEbq3knJGL7PJtlr
sCpDlmNhW+rYVasiSuLpsPQv3OE7gkuoo3bm1XHhxZqQbHVs4KjYd5xvpawG
0mIa1C6Cp+WsqPQ9SHsWDEwm5QeQu+8v6caZeDk5hrzplh3Y01ADjM8etT3/
Eq8usKDb0t8VSBijKbUHaHLFqLrj3jTACq2YlYiab2znG3EXuMVwcHeu0+el
ThLPknCyDLp7ev9ynxbAv8NWR+kC3EhP8OFzPu+SLzMEpXXlAmrNN6jRABM4
jpa8r6hzeEgGttmzh3tEj4xBB6Hi10Eokw+6A3X4KnqlfURtb59ykGjYEvI4
jYLbSVMv0AhxHq0CqTh/fYuNs+JRPD8r/EuL826U8/ZzDd72NDSk9ZUiUpWW
AtDCpO1iwUdsrUMRlaz2E2kxAB5N1ub1RvS+c2kLKQurJ7c5/zhzyEzvIvyI
5O6iIxWd/iKTLdMj6HWAgiUpPxACSKmdnwFmQwI3BeCnzEW0FGfRe0rz2tp1
HEEpx6RP30c/BDaFA2H863CGXj8HYcKYVPMEyky0nS9QRE2+YR/Hy8UhmMdW
wkA4dOy0f4UWHQ3y77YK7EyzuFGCQ9FDKnSQf6XjbLb+rr50dKMr7FbIlgNq
g88EyRDEZaITBtgIo7qdW7+keHPC7el9frw1+2MRGqN/daeZqpFWkwUYvwne
9SsAlmYyNVhEvFD5Lm5yfS1Ek8FHtDvpwjpfh/kmxrxRwNEzYsVsVjrmGJtX
8F5os8aJNG8Z233OynIEn7c6Rns3FnSep+OX+18b2p8ncDhAkP+qW1io1Lca
n+/63U1EvgAOWdeInFZWc0QY9Tv1SK3zQ1cpLkTs6lmpMAIpvJRkjt7ZKNk7
00nNNrMr2cjlcMoL3tpJ1Mu0opl8kNrVOrSdYCZ7pStolPtr4zHeQ4ijKw5q
LLJ1UbEZE4IDVFViY7FjSVyF1uZtTYb497gYLbNpVuSEl3E820EpEamgVk13
Luufw42keOmXhH2HXRbgIn5oXYh4aHg6uiPDCHE+SCWS3YHzzzal8i85XDVM
H+sbCZ0jDQevucAaznn4pZDz6xGi4noXdrKqbvF8Eqf7yfNfDef2Fl2gDKiE
GU9jY0w+4iRRAtPPZ3+8uSu6UPOI6HrADLONs5VY7BO/EN6YZqyWPIfCnyGm
8q2BjWYlUmlFdIdeRv/JZ/cUzsM10vnhP10bXktOizB+nUHzZ9lrz7pmMejw
FQpNNj+wEmVUDiXrRQv21A2iawd3+ScvjgnX37xlKvRLeyaLtDzDPJ8qvkTn
mopKw9wwAzollqT5Ey8sPejxv2hDolgZ2KPBKg/mPwRuM9m2lnFJ5OddqnsF
Ycv1WbesvLO5xPZFbv0MpXYIuyZ6/6EP2zcu6KxF4hdiF/mbM1fTeMV2uXlh
GVpvjkyU+fSN+vtZgiL+fD2FbdHHs71QaXmOG0Oui23aMJ8LadgQ8BdzN5R7
i7uBJapv712xA9e+vLoAh4JMT7IxGjOR4s0YL/V1CollD56ZneiK2wklQLJA
pRtT4Iv4h1gWjhHwm9YHbLVbDNfZ9L7amhuKW2zDxZAmqJy4kZuE4PpU67ep
8j9/o3hhoURmPq7a6a4DhzTyohDZgJADubyx6RxF0F1ahN/Ktz3ai81lTLj3
kDqxZO05px2/2Z3kdcN/JZoHgNdSTa9Z5zEb5kVCK2EYKfTqlqAsehG3w0A9
j77/wmZXxk2ol/IY8o/Zkpqd6/pKo3uqg9SEKlX00bulnvqec1wTxF75mziD
a/kG++gOCyzDQ/Pdp1pcrBQF4mtP1oR83qvhivWhgBuoM0oW8kOm48SWNSTz
dJUfOy2o/y1WPIIrqG0S4SS/KZTBKCN5fmJGkKOKSo26DOKzVaeMHJDFcRnN
FoRlM5c0SgSYjplydIUTmnusv9LuBgjAUYbusAF/7Bqsj0GezW0hEo/Y2e7d
RpCiCEiobZ67qOjIwUWmtf/3fl0t6YfBWQL6tkpuRXDXM4n7QxOBN6UVDixr
Yp8lAKd4vv3TKDjkOHQ/xWXRpu8j+1Wi3Kb0sjYmiK9r14+idjKg7gPiV6c5
0Yc3wp8bNfeo2HR/F2dOyf63OQ9amfDkmYSj6YorrUCDyS8NKWV1R3B8XKh/
bbxTZOKfiX3np+jPLZVs47TNRH5t5ezSy+AhKCMwiCaey1HRd01hS/Rc7Lb5
stvWhtzZQvRCscsyR2quL2cXmxpdg55LYXcG3+d1gK2GbC7YUCkmiTqnWkZj
z31YRSAfdH4t+lCLE9wyuX1Lt/nI2MlrbZ6yGyZuNV/L5bd3qCx/s8Ey17+m
L8YgXvpF1urp0Iqe6zzJv5cKQ9QasJLRwIwlvA4spucMr8QjeSn3ErgfnEfC
UNPe/5J7VZJ1lJd2tTms2GIgOP4iNcS5v3evF2WFmMyhtcxifKiZURSvEHDr
P1udYgHMvP/fhQ3075jo2zYnT7dGOegGFaglpBFD0kwkn2/2mCQ2IYbWLDlT
PdycaFx2+F8acb9pYU54hdWMnP2J4z/ldp4uElyPKOzMIH2zrP8/DvpB76d1
M+4lrw0+QEVW8b2JnS5brDiAoW7ca5TZttvxdjvRaTZOTE9IcPjyJunA4G37
aQzkkIs5cw8JvWlT5FmDyTgRENlQTD5Mi5kbT9dBpjSJi9tgP2edgM0jII+j
2b3Vpp//lbTKSNwV0TkL2iHpr+bka/gR9sb2PJnpYoGF1MDoblcYnUVlqCMN
GA0Mx0uYNCyxqq4TEDDI1sUCD4mKDzKDkdIK5WgxcJVxIE2sh900b++asy9/
ktlPUMe4M2f20pfxCHDLn0A9a+s0bOweDG60MKdeFKsazuXyIVCuRJxO+TDF
fKGHPyaxB+mJvjZYFfAHL1vzr/ONFOiXSXKuR0fxe3mJzmgz2dGsBR6j3qIF
QTLlHSHGTqKEf8GqKsKCG6fxFXUyQP+bcP4Mo4mlhl8NZJiHbG/nx8yj19Ow
MFW+036QK2EYPyXK9qvAVKdE0w3ZC+xMj7RniSSSdVX1vGPBWspHsKibRr/D
2JU4gQt7RNuklCDRyLAiip/S5+fznOmz7AutRh0TyaWOHx5bhG/uAXIfsnGP
cJBHV+5F5MwHo3knCXEww/qWi3bqPXolrYB2ZFTeP9CczQAALRMFZ1LZ4aXo
vHdZcuROm+5Qfr6fCf/dmrP2rX5D1tTyUVWg/RxniRzayoM4qbnCIXO4tFKg
hn0+CZimct3TGOe0/R2zXIIypVEOHdICA4Naqeg2LuJi3NLbq2wwQcE8h1yR
A44Boei009zCamEDiImcraa/5uqdNSiEqR7GqmK2RQdLwvYfHG6XZMoSxy3z
WxaBFNrid8cJ8/weO+OadXNa1Bphza3zAX0kZ8El8Ve37zsS2NRmepin3Gau
eaNaEnXWHs0oOfP8h3r1dHEYXegBjpCZu5TGLVKQdzMt4DCADZv2DakiNrzE
KKH5X4WSXeKiA+BAuKSHeGLyreqCvdgLpXq36M7Ocwe0m3u7M9enBL0CDw5F
v9dHoONRi3frfpq/RZz0ncbr43hF8QrWh5dosWACHxuSEeL+y7VJ5sd8JL7A
F9nwcleG+Qp8HcbDk8vnocCzxeLbxqqVi3RU1kcZsdIhRAhh1Mm6l7xnWi38
ZHrk17hk27cr5IeZmCY8rRg1R54x2z6O0D+TYATl8tF3m7D9YwnswVrXGYzE
rXzB1uLn7d07WxMhq21g5kfEIUXQnlY0omN15VEUk8vuNuwi/of+KuWSwA43
EJckWlG+8VcfthmUH+AzqU2zV7GOVrbn1v+gzXfp5JciidKkCGtGnzq9AcRO
e1V6/WUxPuxmYRH1ZYZmjZmAtYszs59enTsSPwRE76WUhtUNsqTC3qaX+1ob
y+MpG83ljfgGkDo2+g3gAK7fOVDSOAzrmPsWCFMbkRFI3uMuIaYt5c7ro7Cj
q2MngyYyicFuh/laNBUp5yo4iPhBEmA+9hKl3xy9rPVD8HxQW5cnXQK10RW+
adKBFY4E0q9zv9SBx2ft9JpBm7a2pqlsbhi4oyhlS9OEmBKXEWcRc1P5tBGk
CdZpqJTkSi1WCJJZHWpF9Duo32G+p1z+qS55FAdVUmFbxnPweCkajEgz2IaD
+qZQ9D+BtBar/t5G9obumZNRFRFxwPMVS90I8VL0WezJNPY0E0RsbTP16JFA
et9tYfhs8QPKNp19RYe76nUieI2QFxD1Vzb0Pvq4+EfzNvkh78vGf+2rAZKT
60CDYmUyF+Bgm0TleHheO/ic8SzHucKBatEbXvXm0mCa7mSBgRe9wGYSvOhQ
QTQPk1yXEuICuVSoVTQ11pJqgdxElURAvdnALz4v3TMepZoxCkDz8bQ9JZWz
DQfja1HUV3bRJF04N/HwERKjrOZUCuh6S2pT61dMruqoT07NWOpvyxxUQool
KSRmyW/JTzZ32GzbUKhAQNm1BD2/fnyRlBkOuaJnto1GN9npv6mPPOfcEKal
BZ1V23pnB2Hn9jiYcW3iaD9DkRgEDF+v1GXeHDcvT8ZleSkmyCjfgb7j8UlP
5Al9fChhYW87qOaaWN++dT9k+T2yFMtEvw/S4ui+OHux7TfU2BB96QrW9Los
FGA+XfNFv+VBaW0rQktXZxUIg3iADnJM15NVkxZfYIwXzR98H8PXeBqqrvnf
5dZzI1Ufg8aZyCY78fRgxCJ8A6sIhsvyVcWbGmkhPs1uLW6IUP7PDy6cggCQ
28OG4/IjHXNAYR5yaRT4vkJ2UGzfNZif/i7mWgdQFxA/W1z8KEFsMfWTbD+T
6Z0nL0GFv6v3WD4TGf9D+jbupPMTtvGx0r5RS2+gBYH1ihBTlGMog5RLhdsI
oQ/lJY/UZGz3IG1kwd40ssi0awh6SHnsdwXwZKQziIh9ufsgaG3ntVWhK/cF
YaxOBiVrR+XoyiMWRTzl0Ko2pY9Lcu8S8/fRWooh4ono673mN3nLGYhoW5we
+q8LH2PATm/r4DsmpuMGoq1nBVT993M9qhFwKiDBZoVpUENjv3eQDENc/s7D
Z9vVIZQmANxyqoNyEhn2pN1TILRgOrjsOEmqApW1z5kPXgWcXA1HrV64EIt9
zGT6jWmyqgC2seFOIJF8AcGJ2xmBLrzLXYhmjBH76Q0WQe4kWbzOAuGXB1eJ
g+Jje+gzcCprkRp0YUmicDzWVJtgRETyK1Wvdho2tewZiyGnlr/bg59hoRPt
JsME1HCZo66qJG4EIViqx7XvRjhx6AaBCBsOO48VRkyTBfMjapTgenkJWya7
zZHRuTvgrDR2QmMG8L1/tua8W8D+zZ76DqQXRTWefVZep2E8CSch/ZCi5FGL
9/TiFrhkgHkpDzoCfQ2zH1zza71QnZKg5ZnIenpHqLpK+TbNMCwDofmc1aWO
5Zt7zVGpBgxODIstFB4jPferUpdYJEreCstQn4RrD4Le7nKRqevzE46Kyi7i
yvIwFssvZfSJ5RHOWbs3Yk0JZdFzc74vVQh20mpYNs73U47tP52txCbMDLUk
Y+ryOK+9FxLlNCXwimR3t0IJLSsU9rrvFxQdfPrf3CCxEWWyRaxR6bCXUPj9
2VlqzeSIaUFhjsepKBvYvAwcYg5sYd/IM4p7WMftBazRZstNvVjmy6pQKM6V
yiL6uu69CP/DgI4M+w2pdh11ThSXHFTBy+H/QqjwdMnd/QZiKa73uSZi5JmJ
DFC3hjbX0LiJqSIoRNIbA2Elve8Y3cwHR5r5TzkyuPIcpxLCgm7wU+m3yX75
RYcWdSUR5Iq+yelL86GFS3sfik6ewFKE5rWKRP8feyoH2sYzelv7IYBa0uZK
j9qTNs2VNFeSus04IG/2v3G0Z9pyMcVGW2hdi3iW4Bww67uNfcoBoOPryue6
RgYgX+aNMwaxNoJUHVhrPmjBuEH+SvDo95UfXR4ZsA5IIcUbraS9SJBROCLh
ZC5QUe2v3JitONMAN437XGq2+F2xwtoKiduY454rDFB8dhLVNI6WCaARSVhN
XBwFuBkCTMY31LYLvfLf1+K1zgTuRrvopQm0SjuPw+EesVPPfhj+k/Fbv8GE
dQLawg4pNpFB732uFIVM7xXiNQDzcRDQDdmvqIgLaQ6lVDDhBMVJ8gIo0Mb8
+JuDT+T0QzkS6w9wF7RAuuMEegEOnSYTgNplnoLGmwSFhNcjOh0ltAH8J9o9
yDj1Pni8V/QAx+dvjn5QF01NlTgS1Y0XkcjpSgthjtlZAv9Rco3azPx0plJL
rfKM0fk6pJWxhIRD+LOKspu5kP58qqB5x6bDdv+nlLAISTFUrahbDk+IFt16
ZnpBlYrddVGzwjPW9jnb9iUl4RJAwS1ubjX9/fZuKkP++DqbnCtNlpQ6rSAm
F4vck15//U8kFk65LGBgGlqi91Kd9t6ximBrBcU0Hc+fq2tvWEoUBqAUKbpD
fB1WAbodB9416SLjz/8jNglGFivbTw/Z6NVrTB0bGwDUfY2afclgiHgzZDW0
BH2oLqEr4KxEhoH2pr7I2dz+jQP00mdMWAwlcItu/jsF0XvH7Mz78dfZN+V0
MqVJbv5nMocU0EXEZ2H8AieXI9jSMTG4US9yASejRxaXM1q8dmn2CdvRtnXS
BjD9lGWg0zF8RB7aX6lHDfN87Trp+CviR52DAeQgubTzeX2OPhFBd8p/5lTG
5oLkqYH23jeD5tC1gtgrWyYQ6G9+B+M/tVLZ3zdWa7xqSSA1HEwqBrsMzR/c
/g9F7i+cfn95Hcw50IYugcPQiVQmLnwEcdEjzEnwdp162Q+et3KP2qGLyBJ3
vBAWtIlA9VNc4Y8v++pT2q3XN/egDXvdnzO6oRD5z+BNf8Ee5i44jUrmloTg
SiAdRDRSiHynZwkRiphq9s02MF0NKJvMOqPB/8ca1RkIqgqrz3JbrIXwMNvN
yDrW9MwTqnXz1DKP7lWVRkrvXJza9iEETizVLAdXov+/5FVgl+eB0gGbiLXb
YjNSGEQ8E6C3VsWZWynBYjDwCfBTVyYT00b7vJWSje3NhdQFpXQqumYcbnR/
rSk1exbIVgZsIiGY9S1GZRt28unBZoFeYH1Hn0KzIZiheO4NiaS5pdYEX/Rn
06YKMICz1QUs0ppJ6Dov+bFOZr9jW7Jep+ldkvi7Fd9rCheQ76c6FcxukcvC
T757zER15RvjdJDrjrqRzFnqvAugvNB9DoMj6Y3+DjEeXvEw8TLnHrRvqD8T
5LEU6BZG1aWjtuedUaX2tpJgKfp/wALh1pLsODbTH+4y8CfX/yqyMp4l0XsE
9SUYqoXJqgnzzj1FAZd6fE5OCWI+xY5eObko5xoCYSxT4WK/wNJ8wz6lAY/j
Ou6nSqSNpyCaJ225htuW81HAqs26Mm5wroE0EUvUSIFPBhaV6eT11hTQsM9B
jAAq8Fd6xiD8C5pyFQo5w/I79c2XKKwOKDNUZ6rxUDovCpIFvegYV7YKFaTf
nPDFFGWIH1p9F81AMfv5Ff+l32XhfRFh7b978cGaJl2iqxtlo3mu1TB+auvw
g8eNR2ygcStHIKgdFQz4kC5Bs3zcHfLEVbi6xGerEePIF5FuSQype8HAjF1z
RhxswugZ1Hw9gc8fFaMGpjbs2H6wJ+PKplSjsqjiHYHshlTefxUfkx17zy2S
EmTCT6LYXa/VrsvHFFkA3is867K/eax6fDSwr85qlTso6DPlQxQ4/EiOQ3iZ
fxPwh/HLtZCrpU2xxnx+1guArlm4Jh+eZPN8bnAHm5oiFqGYIThMDY7IhudY
wUfgCzwol4fCHf9R6ZO3APSZdkUH059fLoz2rqCR4SonyicecIKcuzi1pNeG
Ho1XaacLOjJ+OAgDZzgmPlN5ASst/3pRdSlyeyIqc6OzqJ2KpIKpeY9Fn/L4
Cm0t9F/0ORYPxTcLUJ20Npe7+V52YFTCND1a+mmAPgqYhmqVP5NI5Mcso3S4
4//lFUUj3/0leX0pr6NF9ducYvsnPOzA9z4yL472Ww7GYnBZa/7WyzMYdsL8
MHspYeB07e5Y3mSASlz5SghP82okkPb051YsW+J17VqegwGpPW4D6OMyUCP2
JXKPDL9+0o5XVpgf0iuwDawaLnaY5F9M+yMTmajKr5AXJ1PUgHQgy/LWcKpJ
PZ/wQBoJMQrjxBYp7IlGlXm/P7t4EcK3tzOXIEqNAiMY1z52nWKcWkv7WtyN
YyC1yMzoF9lusp7c342CbkulBw0bUpWDs1Mhu5x1N3tnMQiCqOJvMQczpbXu
56DQ7f8VLdXw/lVcPq562V2vi3RCyCYONeBvHW+FA3tL41NBXQLJqzz7nikU
owHTx/fQmUpcGwH1aIHMoPZ67LMfd4XcAacK/9kKefUpCpQzhG94xvw3jqv6
y3qbvedOEC2UqSf9kriKW5ePfnPVe2zVqBes0YT5w3qhNYUwSzoVZWE9ItHF
8nmcNMvVRqvinQ2QCkOkaA/bTvHiV6L94Rgpyyawouz4gMZ/heni+jDTFnQI
rMWREt77PKYr63ZdBszcue6jd7SNYgYBxHVvBo1vBm+GD2h2NS7wb4xnbsJu
wiQH/cbLQ4+5FvU/s6miENRiEHsYXEF6/Rw3vZn9ALff1uJFW3XKQeN4K0K0
6fU8cTuYWdjTN1+G/eyLv9NbqDlEAxkWHGlWQ584wd5E1x6vugC7OBAylyvt
nO5FpLW1lbfjdnJ4b/P9HMIlk722F2OXHSTmzwcB9SGdgrbe8jq7/TIzmHVu
GRzj8AYMCIHhn8tx00I9KJJmDJci/Cua+MZQ5OtfnEhM4Sf2YixZmYkSPPVg
7kPmS/PiovNlelqo7KzCuUAxN/c+5immbMgwIpZlEkSQd5BP+nnNdSOeR/8A
oDufg3+IzT32OkrnaDun4y2ADqDM6+755gbpC+FHq9JT1HI456402xosyIVB
HQinpNiZS4kyXXs1AgnTPgPPPdVjHtmOb2xX0x+jXUQ/QqJ1XIObj/qOWK3b
7I2TmX4iR8OWA41D5yLuVVAEiKrL6yFKHWfmiL+RcKeJJ8RrxdOAFJWP7BJK
XkE1UWPkyO0WAbOYUGsqbXx6Ya+cXvbiPycBKC3woPuthjRPfNDXeKtu7T18
JQqpUQyBdjoMnf7U48qCC3QP8CJeHx4mVCdNcDT32qkZ3MBQvRPnFMQtJSwJ
GW5RBn9FlQUqOlARDSk7px8+dV83e/AJNTUmWNp57kAm+ME/bQEqu8bzN/2D
pe+kaC0v1w1M99dn2eZ42jC3V73Rf/6KORNu2s1l5a7364UollBQluNH5uFu
B797TtKJ92cmH5pd3crsVThNP8YcP1+HCyWqVPvZcbGOjNS2huXMVrnV4SSD
t20Rp9hdgw7mAiU/1XA3blm250w2S3j1kCYoM8rtCyF62rgLZKdiODtb5BTl
7he6Zk7KZALqpMRMpUkD/LET90Dav/9H4Ixr1GxLtY5ojLfeWv7acWLziEQN
wUaR9ULsGqSnUVfgGPhOqIQZAwmx6G2dR5NPwfw4WjfENzz+3ckz7Nk4dvDN
KRk0q6d1luhArH/QJVBKoA669z4j8vKkcyTtt/+XeLp225Qc7Tl4s+rmIzmo
yoB63MUmqXi8EUZqI4vfLda9zm5EQs2Bevt7ln+ioYpp+8UTE/f3umUFma29
GPaIzgDxJfK4wmW425It35vUZWaF/N5dlZs8n8zKQnvDGBih0ljAk5nl4rdw
7LztJ38xO4kBORfEQf9lOVsu1qccyX/w9iqu+Ep/PqjPmkupRdUa2mwxULnz
sEaSj4d4Ee+bV8CkzwW30YH1FQXoXjM+xg6MmPSnM7OVGTVyG++sOBjiJuDW
wDw1UdHsKSnkI9JEZQdaACHJrtbdAtxEkinkEEfmvMaoGaOjpPJFgdF5Dxyo
ZrWEh3OaGHvPTj6HTTy3c58pr2ociGWjaq2xNRLPtAK5dmnaUhL2qF0b43Yj
KD1UKUTqWRkd6DheeonkfylvL7qNCjgyzE0RxJYz/fDih2/U7o3n+7naf2Q9
BUV4woifAranphG54kCC98bqjH9g8n/o8tAS+IPXtRpAWQRLaert3I+hoL2f
phT4PEBB29q06g/nVbXsHqmXHIGLkkcl+Al7lk8Ci+AhcESsWQ0eiGlwmk0g
CqfJIYCh/1JX03D7evOG0CTIWI5F80nkpXYZur6w38w4wBpcN+DqTeSAW27U
eH5vVdVWfxIHguhltoweaatVgbGPqW6a/TLhRdYpdSzPwWX8RiiAFqQecuOf
ocmJrqxjwvX6A4NeDGuvx/4oSQk3Cj1x6r7BVEyTXezfXJfdDgxWWTxKERwT
d2ztvJ2cwa1waHQ0denMhqgrFIMo/0oYxE/+eYLZ4vpDF57fh402jHvVg9Cx
4+oxN/j+aoD7osCEwN7z9q+vTlSkqdE6r7ux4xCgmg+jLyPWUX6dZOgTBsRK
zF3fvte+4dt7sizyb+eJGuim6gR5aJrPkCD1gQNJNwLd3KI0n+UXCE0F74kz
Jf/t7kw4vRg7RmCvg0+kZMBYAI/vZkav0UyDIBc1+ShfkN/b0Lj5a3GT5A7j
TmIO+UO8ecvNOO80YHTyf/GSGFNoPNdY29qNdAbSX7hwmqzm1/EdFbNk+ehU
DeXR+FK2jweH/WyqKJNPoDSMvkQzm+5eL8sQFxtoj0zqhzXkjh+oqFliM7ep
66svxPJVkVz48R0kJMdzQ5QQdIzsfD1FKzQ9Cy1Z5JQOPXsKjV4L3Q9Vsxth
9xUmFXVBOZEm7j7dtx+7G7dRpKkHNHTh0ViqmM9Hqc4/EUuvLAphZcXr8XdU
Y1ioAJ2w3WX1rK7Jm3pDhck1N0fbFVlAgbsk/DGCZJwBiw70uLIc7pF1DqgP
ZJm2Y+7y34TEJ2nXVz6Oxt5qy716ax4kzRx26SA7HpsxlySiE1IYWe76CVok
uH5bonxn7VEr6YUo6h0LAjDWO221vavS6YgHjX28ppBa0F755AD1em1llzMy
mZEM6lQ8Jam5DQ40Cv+jhaLSBsbLt8fcG8EQCiku5WjxDFFRhdAdqCZQor4T
JYbyGm2b5pl/ahERs6fsBqPg4w8cHW1svltAjGkmyr+t/KN/ZJWkIVg6jQd2
Um14SVtXShNlveE8tLnj8WGN0yH3gqOhrb/bcx09+ZyXyjm/lvlIIPXsBHoG
KR1mXE6Hn42wZ+GBY098Yn6AKUG/aKVvvsAMOU8z+d+prl+uFCTdyyJb/eF7
PaWAlfIeCTnHJH8ehy9F9z+mopx4gfIS5QDoKdBcGqxxrhmj69G/7wZ3eMQA
KUonvFSE4hh+LY1/x6LWztz7GZTRvRwzuLLNzOTVxDrDSiqs43V9hos0n114
7Y9YxKTVylnNO9jm+DqiVaUHfVKsb6Fpk2TNmeLWIW4gVUQRbbfKGjikcxrt
/kpdDHZUHgMAenfUY7S1U2jNoLa9gzTR5dqf/szv2t55b7EqSZH4eV3Wu1zh
fWB0qD1g/ts2wIpiUNvtcZI6kNy/V867PrxKb03duRM1mbFz9NIMDfIrtgdp
yPiopKgbl9UfEIjlvYk0J6OFmnI+gumDUoaodXRRn3ytKW44zl2vcv+XX4eF
yD/CHpmEdlBFzJeYjn+rfcoyLGEIrMTnQ+v5Zdxoh8ytEUy8BC99SNN9OHqu
xt7e/iEUO1+bO0n4TzUmKouBvV7E3sH0yqB3t+6AVTQw2yteXanqsiwftrj5
LiHr5zQNsYm3YGg5qE9ix4YoGjGcAheV4dLoWp5xblOf8FHLEdFMq3Wk7gua
dTO0PIk5uzQ4xZrbD51bCqCjLlQ/w/d0/Z7i6nZneAKyyjh8QlVwm8mxG3Da
/GMp7E378hUKAdzJ2R4Cs66ZOg7EOtX06F6P5U2fuOL3gPOVSvaa0Hbgos73
nm++Z9wtoWn2yS4/5eC2+uVVTi3AM8HznTm/HIl31UjZf/gDnX8gVXwdxvnH
1qNl0kI6WkXjoxhPyAPiFlhjxAr0fL+RK+8ka3ZQ/HTbmgv4xR2iep3QUZaT
XmuNs1Tbq4UgpCwLWQA0mRRyOpgod2crwGFt9/m3eb5od08CoRj5RM4KpbwA
DrcvYIgaE7lmXKFayN1LKAN9CYBMP0KOgS9yueGMvQX91tDot/fltPvyEeLO
ijoAWXRo7SF7OKqCJLEkBNOsGhhj8PNyl7+ROonrefN24ZJX8plxRzp6MyI5
vGQdCQiRzoNEZXpnCvBiSNt5l57/deBhv/h0Pjx9xG6yl3AtDRQSQHK/OTyY
8NQzr4BYQioMk3Fwo3Grcmm0zZzjpqSd4fcH0dbifs5BgoIKu28QzsvCZT+i
u0ospTo3RsH9J+1cvCfIFZYF/UvGxGZQX/1zq6azP8YuWc2dpKf7LB/xxU3M
E2bpyI5YJEh9LqqYeHZmgP/UkMuk2P1j1jQjgMmTqHp/eCNlcKY8uUVyBgLH
GWWKF7w3jf/ME71tezLFGsGVILerLB5EhLtFjZBfzzSR9dV2fP16wEVYHv2B
XGQ4Zvp7PGgZxV1KghRun3r/reSBq1vp3dyTKdAlRbe0MHHNDqVl+xnBx5jS
FvfWTqGEw9Rj7WgQjNs8sFWjH11vYt9P4l0bpkyT3HY58o6bYp7Hio7EtTQg
Vpae1BlC8vYQVrX+IUAtnI0aiw6J+LuWRrxHxeD+gvZifauvKya8/taG1NTN
KtOR4EupGUXmECjXKAwcwq3zjVCkEP7AKsrm2WADlKCaxDGV3pSbUB6c+Isj
4czilaipULQgCdY6jsKVHFf6MV2+ovRB7ZCIs+/+jKxK6XDDyHMbCUGo7irC
u4qidaFSrNtqofHrKVti2I90DC1+7r2H3vNlrIBNYjLW/1I3PDFfKsa9MCOK
656Yg5SPLcgcVXZumQUOKDTmc8hD4hRp8DlDrMvNlt4TmgYyI3rk6tWG8JU4
FyhQ/M/+4poGR0gzIZyD9pYPEjoqaXzEx3tvOPvkY7zr5qLmvdMn51mjLwUl
PWOTaTetcGZPQW4kfppQLBjCw1niNMmtOHotoEgorB81PtAIRuQ07gAz1cQj
BmiNlgC20BZGcGsXINWrUrCzG4BJly52Z5UNmn6o8L8ElJnMKYXwDhluTxEp
5A4fGpvJmahOXBTSX7JSOksquZSKRHb5aMMmuowfkx7rA5FP+Qe4EfkqyUXK
5g3MzmmqGSrAv9YxxdWJRnCAk8NfY/X2Ft6Q/XSnQcvvYyIALhdmtjWW5xt0
XviiWU9TNmwZIPqkIKVaay+y34Yacu5Dm7OaZ2aN20oZkPuDs2roiPfjeS6l
GddwiNxvdc0+dtxpgg0OuQ0/JslgWYN3xLscy2pNysPZiKYEsZ72us/z+DLR
eZ8UblLTeu9ofsn/8t6vsYpQwVyBq/tQWUKrGvb13nIEuxAVpkiWMl5pd1HB
tgPDKgCjybHasxGQftf0CFkikuG8CKzNLEbk6ZIxTP7q3/irLFcsBHQpIdli
F332KqKhjtN/a0oHj1wb0VTtpksl2npdQthZGjr0Rn3MwMm4XRl5o0BP6Xzv
c11xvGDSWcpAyDoP7GbjdtdlQLlXNjembzTNXld+gXLzRvu7W6cC4yfz8mY+
yfBq/sS6skPQ8eoI2PAOh90KwFGGb5oKj2YRJYFGAAdth3pdhUuDFa3BsKUw
fFsdojMixiQv98MJHwlNM7SmVjTTxj197tqSCEjnrDMmBX+5trYqpZFtUPD0
xcee7kmM5/PxyYA4t+9mGf17xwN7Id2DzOK5VErtB5GCrMCE5FjgcziDM9wE
B3fSJGqM+2vXlMnA3b2Q0SbNPJXaDTJF3A5l5NYTAQlvyenB0av9wRV7FBPp
20rUI9hdeg1hBvRTcnh9EVCEIT+513+/blWXKLd003AtDHbv9c+WFYpmxI2a
ANdItgpmhASmS5qZXCN8u1VSuoA+TVeyQfShROfCJ4KwB4saWTJoBrcOtSNn
x8MW4H8vUaiOy5xQan4J/5O6YbceZDd4H5PAheNciJJCqgLMGMEmyayJbbIx
LHxOiZodWQoxjj1TfOZOA2eDlMxNGiaTB5n+MmO2xroqbALDZvt8U6wZ+d9R
H5bTrruhulnAVK/PAw4NyPGV+8e4epdaES02coModdkYnI9QVZ1B55hDMODr
xIrFDrgcBC/dhRLiYw1qHRzWyudgpFskZVVKd75jcHp9ejjjmTE0zlJl//eH
HJHyyG6jn/Pv3P3LRB89299aWK48cGIhJc7Ii82VyQbcwcA9TZx6vHouC36I
9QWpDaFa4MTkPdy/KKFmwJAfsvjrTRNAlHtGu92Q6WmlynWzSysGXrjD3YTL
OVBSFNPm/IQJBoE9UvOUHrjKDxK7QtGjaiNaY/hwkM9jN26aQMuyAF79l0j7
l2w0vSBEClLpRmb81sN5ByYotJv/3ma6P8DEYV6LGl4VVH6qlRSkkpfTE44v
AxBFOIpLjVBUctllRLbf7NwFIRH5UJcaE6hoB9GTGtyH4tT1jZaKpm94n+3x
904R+XrAIMWs/TxDFiWPA8eupfF0ZaqwsId60jS2UqvTbGl42VS2BT8mQ0Nw
zMBJPAVKjVcgyBDQEqQ/TRgsFV0YqvBhXrpu2BEn9Kk6+JY3L/Qpd1JEo273
oayj2V8fSQRPTkdfIZzKWwQ0rL56Bj+1JqxOwG4bBeWDR7KK9la9ICyhomLk
yfenojfRxifsT+m5nF1MQhtKFRT5o6TVId8zKLeHmn2x2Pz8RnORxk/o1HTq
AhmhwZ4wPLE8rICIo6MQWo2/UA5K7C1cWJMW2yj43eFU4kYFr0YLJVqE/6AM
7E1xMMdraIY82PpQe/30Cv0zH6JqIyXmwngDVplvGVZ3//i0hmvZ2eVH7C5E
3Ja+s28TphOhwXEgMGE6aPL9dj2MT24HaFSl2yFRLrps8xuO/G2h7XFLwfWT
bfvTGsQywmFR4JUtZWHBZts3gmn1eu7HpVEHuN7bu3aoegBSmgA2RlQYZLae
ShPR/G+9f2RlJNmXu3bfu+7c3DiJ5R2EbNlvRZEl+I+UT7OuH1iRb+a8F6R1
XzPRQ3EpBg8exGbbwAh7as5V3R8fGw6qVH4iuwmYaDQX3djCzjDQh/Org00J
4U++/bQ7fjvsUs4h7Qsay9dinmsdET5UkfZD5ZXNI2da53PR3QIbiEQlbeFM
tN1yJyaG0P+j3JKtuwhUNr1toaukVtCyC77yse4clVqIRGFCsfiTYvF6yseR
KibwHiK7tWNCoLc785Vz3fK3Cok1tGZZdqvi5FaE6f73IRNhLC81rC3h23Ku
BiQXR2gNHUu72h4QMvTleqry6ocRV6mUv3/T9ZBCWGxctT9xpdQwfVtE+Eeb
TO0qscGM0EuqSwIUEYnqAYOjJ79iwIEP1cN577kWiKP6t3Mf/s9WhSnXa4sx
s8qoXyQUOf706flYOR4esSVC6jH8atpz0fArilQ244kMlKy+Sm5kqhPDvZNc
yR4zMOcfXXRN0VPIR/9WfZOPuiMya0LYBo2JjxlhrnJwPrxvHxnhzY1is46O
HQ3GHYBn61Flzk5kXh6SANo280UsT+QoYqOly8PdTCDovcekJON+mBpo+y4e
350WAHEQBbfpkQUQpZC5qj4SABo82529CeuZjLdgAldYkab0DWeXnrdbeqC2
XDXuX1GBCxSGmZme0X3SCPQf5gON2wOC5S4uyaHilcQqPns6hWmOX/fMWepr
lN51sf0CR3tYK2hEO00u+I8FTj/TcnF7RMnCnFI9y/1e9EryU+qkUBGQn/f0
DyOXv5f1zHrjQjzC2JmoYovQqRi3uQoWsUmQYixfh0j3En/dkCk4dsGNSDsn
9LiBBCU49ooeP97FXtyvljlsgYIZQanCpIYJ21IuUPfBeddsI6HUikw/tBvL
29t6aw7L02WwJ0EOFz/aJfzKMzcI/CQ56iveZuLmSCTD/vRmPM1xkptisz2C
8qLqAzcT5mn7mAij951loUhU9sSsbqqM5l4mCh/igt+QPZWbyBavFL7AG2Z7
3infZGqrZdoxyPWZNl4jeFJCMr8DD2H5rTjQKEfeOyOu2IcQofm1pAIKyivR
FZi3ua2PvaKewGiX0pYtdMmV6aQPzDKKd6ZxnMkY1T4U/O8CFB0vTSgfsSyh
DW0802YUP12Gd7Vbm+TX9fuycFee38LlrFpiKvFLl2LCyG6mod3c9wH4U5L4
hMa4WgQKXAHr83Y1eiu3FVCqstlDQgkZsBM3nYgAz4WceFf2cZ4v+4lLKAi6
ndMFfwd/jE5963wfE/pN9z74Ds4cG2d0Ge9IT8mniZmttPa9TAdmAzCZIItD
hoEG7oOYFtrSE91epOAhQkIRuSqC/ZXQHD+/EymVQ96j35LZnQEK/QDJ+dQU
8jh6g2NhqzXWUhzXAWfH4OOGfQKhE8KMHCNeWvusrlMXa9/rUvWT483J70Bq
v05jGSbMZubwEqGfqaK/+OgzgWCj/G6RDkgN3nGUjSYTr+KtbzKLhCu7nFo7
KeMHmZ4hbAKY+1+27n1IDJIz4xSYbXHi8TOoRnd8tUdGt0yMT0A4jFwlqLBw
9qWtoIuay0NlSah8PzsVHoQakN7n8HE6K7yloP5jKfOhCcuE5iLJX3Hlusm+
pzY5gvjbicrQ+6hDmMhFq9h65+DY4nySHq+zWwhCU5SoCdQ4qgXbKo66YfN5
c0R7o8JztZhqdxb47DRqPGVQoSo1VUKG47n0dSek6gx8S+gGmHrOAjS2Jnrp
uK9/tZ9YWsVkyv9ZdfJdm45klzmbjS/Os+S4ME0rDk4o3hKTIUxezGe/s4RX
8jGgU0SCv2SOjaQFYWj+YzdwA0yKoNLDAnHO9ZnqPigddayeX4e3j7AEkC6C
FK/twlzmf0Dm+xHc4GIy7nsCiS/O1BRqFO+ervyoymwhkVHLxhSdfejZ/hjw
il2ruflQfrkMqFI9TveQIUpjEBYnOJATA7ove5CArQ9AmXIMdRsehee46at1
EmQmupOg0pu5YW1Jxy1TbuLYBuUddvTiMHjz6YFSkDs0ueenBKeHz70K0u5i
+qtM1x600CMm4YL0UD2FtAebvllasfpZrFAaN5/PPEnziswQ2JKlOp0zSK6v
V3Py0iMYvotsY8oYgId+oB/Ak8aMZ++8n+HmFeHlwTSE6Njq0+dGtuWGGq6v
ob2C9h/9mfErL757sRhXIpEjckcV6+OgZ/mn7GdpvUpHBYQ6Ms/xtk0+7nsI
7hEmwLDR6GQdbaVuX07a1XlO3SEoyfPkdw+oYLRZ0oA72K+Cj4zCf0TMkGfA
57XmKW2uvEfLU4dyehtuxAEUf2uKjQEcxZkuFfewaFwOi5LNAs9JlQxbtX57
FQKc7kS3iyGG6QxCgCshG+pg0njf7zL4pOF9j+gO/ZrH9PBtjCUvtfPFVkLv
KfIHuMuivleKSaUaPrWUfu3D+EXfhT5ZamOHrXPnIMwBkFi/3S9eoZVxZDVQ
FHsSIgPLOxsnOpTLWHRkmrRo7e5YC1NSP1k6V/euch2S5rZaYc9In05GJ9Mr
WH8Qacyqqe4l9NwOkq+BRpsZTXMmS37NrQidqD8059k8hyuuT9808MkHdB7m
TCX2oGY+vKCAqsS9pRVBSz5aNs82UrShU8DoJi/TdQ1lqHFEyXAnSdjKY8jh
oO6OpyySKo+9/oXFQrp++e3XZfznwNAnuCrM2twJB26fQ0oZQ0mpFOMBE70c
k2aWWTg73ZJzWTvJ7ndOQyBGyjP+iWmtCxd0gXaCZjuK2E7BuBL+iBRC2/UG
u66Ygxg+ziG5m6eHPtZWNjwA9yy9X9IRhrB1VjDZL6wcRuFcONhexjyotNs1
tthclmzH5Snh6R7Age3UJCnRly6eJP0QvuvSBEtVbCXVcBjgRYye5bLEatA3
3szGiV/6bFQN+jkLBXPhZxU5+JACBsMf/GRFeKyYSHNtTiB9QZvmc8gZaelz
BoXf7zGy7Pqa631CwYpDcA6zAXx9JBZOIIe9RctNUwtW/uqKvEhooAOfqsXl
vTIsk4Naowhh5xNnky5KsTexyRNfIqckXB4p0OIZ9cfry3zMeXNSego3saVK
LPwF3R3njZotKrWQWHdnQ9ixilnI55I0BdWdJwqhQDuGw27WBnFZ80dvU8po
jwe2z6mlPc5/UdGDAMRNcg+mQ1c1qPzRZJmD2eIxDuNYdO1dBq5j7Vank7RR
RjLuQoPW+C0sil5R1ehFkRNxv6VTtusRH7iwv7ecKSuoVSvT9Y5W70/N7MXy
kmmVrPj7UKKEqfGH0t37qJfnASv7y7FkNj0N8QEgT+iOn3KQtcyCG6wfu/qV
P4GzJlLu6xHboIrUnKWXIldLjj1vZEHDGEG0x0+58n4/aB3PA6qGWRQTHern
TOZqNRYcQifqrC9yLlkgnoH4B8L9PtnsS879XleU5209kHw7pb+izBD/UCVH
CxujiuWgL7poRyMaeq7pZz6lahDghOHjlpIYdJIHtgrpX3+7uEDA9ecFC3DI
sMolHzdemnl8oAynRzXaILtnP/yzhT+kUzTWPm6gwGkcVRajXStRv33PSCuG
TOIvLg+59QTlUWgaJpSk+OtiPxS9tY+K3BMyjNXUxVDsPomryYkGbe3r5Hyx
hj2+ghq45kUIgU22qZImIINsw8esu1X8MwXhkLoKArzHo1wOq8oLCTswu4Ri
+B+N5iqNEpP3f97bGsAazbjRRujpPcD+WpQFhHLE7meCHIq6CalZ8r4PJXOa
A0mcTU8OWeJ3dInVHOcbW9WotPEb4vSb/eugNeX4TMjhLsGByOi58rckMkON
jmIHsci02wt2LZNBoMmWqabxUsPdhTYaXgDim4Z8CS2TAS0GCSk8WqG44Pmk
4RalmBIzhGCVkc+H9mdVPtA25RQVhtjVMTT3gdE6YDu9F2nAlAfUivpTrhcN
eS6VxljvwKE3uC5vPCTnk9C2dYwFdX2h1Ez2LIvpi10ZoWXsdsG6dVwz3LUX
/voNFDr0wzVLBvQ1aUFe9VWXwVa3FLKEoO4YyJTkeslwZLh/RFf2Hp8IqNax
kFtXL2cgZVNhoefhBhpoaZQEjWgPMpE0ccY1LjAxIjzB72f9byRm8uzMekSS
MnbE+QdLrvY79KaLCckbAn+N3jbu9yIGx3VL01aHH40hW0JFQQwMpIS7HTHk
m1eSxv5wsTvSzjq4b+r70zTkUJQ/iusSvv/1Z2i2/S1MooVNpy+NYOgrT5gQ
OIGR3YTiFTLiEL5IIJNyPsCTnAiAXcj6/RKC/HQue3Ow+2Dr0pWj6DNL3h+j
6LiXd4NogpbI2HpauLEgwta998duJ4BaeoyAEzFVeYRGWfGbQUwY7udG1UZt
DmG/qgfqJ5FCbHLDo1ZF3SgC4YKA5BihlzYUQyThSuO9IG3vCDG81kiftXYq
dXiI/kM1dFWWSGpWH3Gg+oXePvA131wNm2okj7QUqt5rR2rgFGr+udKcfOzD
TOoN8yZH6fp1rnaeWkods7DncA2xRNkmK4bdCvsDOFIUsMiq6UNg2h1iBqoc
+7HRiUhpGzZ+ocQY+sUFSRnGsvrZrMmkBLdcvH5413BBhOaR2VNejj8DVCvf
hlBButm7WlLFMwY6Z6pun3oDdppLv/2g4j3DazWTz9MSXytJ08Z1j0zMy4uc
1If2nkenny7FnMRv5hK+efh5elrQz7XOndKSJk/LZaTgk9kyi7pUzOM3f3S+
B1mC+K02et2dN3qdmu2AWdIuwf3//uRS5LYx+EzdzwidD75mgIMmvrALWpJN
DaS5ij7r4T9rHwRBn6GPVdpGoI4C5u0oJxQYu3OnKv00C+0ZYtUCNQ1lzQy4
VxSypEQcXrClcg64fT4iX57tjzWUZ3n8YqUjIj+d0dR5Idr1GmBgsVVlln+F
yfqKeqxJ5Dyl2xscKR+AVy4ZjuQ1354K6mURm9ToOOOlz8496Rb34MGUJoIV
Hjc1ALYOwfSGCjheiKd0/3fhPmZpZ6b4pFZt5X7N25GfETmGvYpoMvyh10p0
bU6dezAzRQhc0atEYJp8DXFEU/BQ1yuz3Mzkt6UhYguRcMlUd/0bWpuXYiJX
hgKyroRaAzWEm6A76JbcPRB7/Dw3SOqoXRn5PcXndagU1Km0x89Yx/MtrdWf
YlrXwV0V8DXKggZaScNb+/cpxE14+3vtoQOtPrBRRxn5ut71ZEw8oDcSi0gq
roWn/hqmJNkOAamgL/xFfgc/d/ev/KfeYkdMkOk5dbzAKLrl1AtFjS0JEOGh
JxvrfvIGmscM2vidUy6OdFNl4ECPYHDUjhkNXD/cdGRK79OwH0JdLW8UjzcB
nElxKLgZEZmfeXIUdp1hKwHjNyOE3r90lZveWkiT6YKiSC8TVApDflvEF5yO
HDAteDsy5fFjBl0rPlAll0Suc/98E4sEJ0NOw4w0Xue6O+j4oxBFToeQpCIv
MRlVuTCoSxzXmsCQPwRd9MeMBARu8Gt+ctPk8ypbxRqDmqibXlFTylO4GPd9
qKBf/+iL3I+xiplHCeYGiZR+w86CVYxL47fJGWuvu96n+hcs57RCsG0pc4E0
Z/a0JBTMq3J58ntZgMlt+KB+UtiQ6bYCFmZHR1/Rcgq6db/X1oo+9oZN8FYC
khnJ1skM3t2irZs1QsTOmMj5XVSDQeJU7CFZf3RAwtTHnLNiKS8FpymHGuuV
CZPRoZ9lUqfFhya+GSwEirMt+dYbncmsTus1qBhWXQ17vA/JPJ/RQTad7qu1
6j1V9cBcXNiiTTF4p7rpJbwCaSv0AszQ/k3PAHjcNFLODUn2T2kypeEOlEeG
uH0cljZ4i/sG6pDmgC8DNGOfNPMSYw9eNsHrM70jPh1CF9YppoN3Mea7ASL7
BiQik+VUQPQfamKXoSwey+NSqlkND19YA7z8l5iifmsHoMJxHWAE5mnxK8cT
a8FmIOfgVNuGiysKRNtKcOdR9GJyyBx1x/3z8ByQCbddI3jfW/SbhteTvDgA
B8dx07JTDIG9O9W2aia5lHGvcWDIm3BwW0gTZ3YcX11W9SoAFSkE+eZF5qGb
o555IUV1JkmwZo4/Bvjxrz5WBHJZX7Nhttme2bwNzxMzzk8QrtNv4ET2Mlzh
nFPQIXUDVJNIQeitPmCHSyj7+mV5IMzqfVxFVzsY/DeRryGJXyAHVgBSRdAV
LXqLoRuUbBkYnuQjFl2zgC71aCgRyRlruI6TELLEAr2uH6kM6x2y0VfWcrG/
sXJgcgcvMiTqcrbmQDZF9E+CSnT7BupnNVvonNHQ7mWqCY+G3KVf1JzBVmUC
VHzXD1bdeLIZyMVfstWC+Mjzl2sGVa5wIb9gHleJfVdqWFNmZi8OnKH2j01H
yd567rdtGZi+jB+IirahhQWhgTq8QSV785raBXI6zbXmO8crR650RHmjNWYt
7zMxj+x3FpjIQabc5KQfvbalMM2kow5ylDSgexZMqz4Aw6zBaJakKbKFJKE+
hjc6uO3G8tbNZ+T+9zzI2j9rYljJYRyaasM3u4Q3Yw9ml5sRUvV7NIizYYM3
wxg/Uz1leg082JAVtK113IgPN8by0DYIJnp2MJwDGKeAP7gjtyOe9GEENrB9
/KT2Qy8m0tKGAwiEgidSQ1AlHKGvd55TV6Wsu0AebAwf9iHcKCEQWeQ4o4lQ
UGvX9aBPbLUm37HxV7Df0+Hl/Mz9ve23YZSc3LxUUip3BdKU02Ofmx2CeLA5
lk02/1uAvchNTXLxP/rEZq4ldd43Kogr+kW7TOyWImrTH9gUq3ZlMradHSkg
mL75BD1L6iQK/eW5nxyrxj/75KAlUql0VAVMVv+VrfazW7Q3Ys2dJOJKPCVi
Up7URJMG2KHRlqYsc1J/2jg6JO1p/SoKqpdePdNuk1LOm/POgk8Ml/R592ze
tPk+vUM1tNHVgJpKDV7XAXWtFYOdLFKQrM/+9rkysvU0HQqkmNeRkFAt0rSB
S1QkJ679kx8a/sKq+fT8t5qt2d2c6O03eYw7vLwrY+YhF59imRuFY+FHdNOQ
yTx3ADACclAo1CtLO1Tf9rvvHzygLcArpsMC/J6Dq3jnaJUxbAqFn80F+kaB
pfjeS1w21tO/OrCXFUpc4DPnQzsBOHdtBlOIn0SPkzgPie+V2x5Hx1LmURmK
qRqvnI5JFVtrWiQrezxkdXRpgPkUDDHh5zYa0nyMyt+VMQTFSQZrERUCdgDD
sD5spUfAIZih0scZRAxbwP2LUsRzhV/07fpfJnd52JjZK25WX9eZYjfxsnhi
oPh2WbSvG1tKjpIH/9yL5CxhFbb7KuOhFx1vXJkGyaQ4ZmwVX03U3hdjxb7J
eqiD0G1tVtn3hmTUWiCpL0haUeluyk+9cfRFESgN8Z2S3cB4alN8fKDd3yFp
xJSQ9CoAlb5a6OM+yViF+oCCh6pavHHMX4E5AWG9NfU7HDafuJQEEoMtU09v
BXTOdolYQeKtQYl30ZGjK7JyHLiAET/80jpNurzH6jsCfiBeKoQ0lGzmZO4a
nSeFns4EYHXivxa5v5QmQNPl1C9PVprD95/hqs11tKoigVpPC/NDHes4lkkN
yjbN3Qi3EMPjReVxceMbMcwtGBOP8DK64aL0CD5J3eUx7xzTi5FwScDzskeD
HFK4o8l2E5/35DkCnFxZzklRKkhfJ5NOM71PQS0apihNN4uXtQ5ArHVs+Jjy
5X/6BPTEogju5RbbCRLUCbZ/Q1XD06EV/Qnyivsfj3j2CSW9S7KHr5VnXgAL
g6Wwc04Gnd6KnkpRJ414r88ZG12AWhypFJ7JvjaVTtPJeDMxo0tdW8snRfcr
ENn9EFuvthoa6aRb7xfILLCj6oX1FJ7XmLjOcMewqyI9DggfXy1qy3/TgVxW
6wRUPoIa+S4aQLYjyUypwoRmp+BZfzMfoTjwK39BN04E3dvQ0DyKruugzjTs
lHTSaK0uoOSPHzBmF9TXwxT4Qez95cV0xaRjnZ6wAXhDl18xXFz03xYAgqIo
NJ279pY7NE3hDr9X7B8LduZAKSuGgzL3401t7lmOB/oHDGfZ6GD+o13jxYVI
pseVmqO9DUnZN3Neh6sL0+sYNIgNF135RYXTs1d5J+pF6M0iQvaZeX8Zgzld
OqLtTy6VI+pB0y4qGwjxlGE9kue6VFBAcD/3ll0lDP0L0wDsz2BVTuVD9Fn5
cU4pkXTVUglHjuQFZV4A+FJzUfPXKpvODLj1QTMHhBQJX47IuqEL7OUr3PBJ
hJDm6+x46dP2c/zwCeqdQlrj72srkDH0YFvxrzrHHJhdHIGLfYIKuL4lLtWO
CAaS622tIo591mWfOSZweuANmiHmM++O19agyIkvigSLh7eonWN5kCPYRSQ9
tCJpEEPCNmjsvbEf/f6JnBOfaZKANFiwPSYA+ipCi6apBVseh6FyONnP65K2
j/WLvx5G7zi/oB4HZ4YaOy6484pDIJ1GfpnAwlxwR/T8V2gp0aMr5wLOA/T+
Xi8kLWU/RcCkjZa+M8Ol2VgeXJWKfSL9Ky7WAtk4aQlctndOk44SJGgJggNn
hK/iJ6YgplqvhIyOCVLt/5YrtYSNk15cyIrtjZ4RLvvTGLOhMA0U4lwNuqXK
zvQIMAhx+7iqspOqVHM6hlEQ5GQCUbWOy53rn2CibQtg85RqMWo1TbhSysM1
H6gkhxtZpeItcyZUqDfqMONH4M58EuvhdO+5f9uZGlEkNAEjG0l2zErTrAeP
JYn8Qskwp1yiLT5Gds5DEzwcCOT2sciRR3iMcN48xOlTofeABpJq0SkwYBlR
S4NGH3ysEqZCDuRYJq2DCCobZZECRCUVtbqgBLdDCYcPKpPI5nt8hJQyewdW
7yECKsHZUBQFQOAqwfxeEx5eenBZAZ55tPrjPzoNtKQqj27NEkY/BO0LGNe1
SeNcNeqZhuUDq4pkhSJ5K1O/NGhj74sOXfrvAZBrM43oKwwt+GJB6yeJY2pf
AMtYU3EaqskIW9fQKFB8K3u38XWjzzHasOmlsuG8LRvnOTp71z9McKc6WpMF
wKC76MT1sgFF+pkPX1ZNE+ODJzx1QLGUo+5lTpgdYh9iA4Y26ABruXWNNqwd
dL2BvpIML1JK9LYw+zCyQzVa4p85l3G9nM7rj0o6vB2CjJToliCR+HAT7Gh+
aZr9SM1WI4dtzpsAsa8PGDiHCwrW5SqUdDLMuR2RFJLYHpxCWzzftcKIuhys
S1Za7QeanoN8Cr6hIkTjQL+Tl1+dKQxH5g0XLEi4NS9woU0QNJofgia2PL5g
Y8Z7bF8QYt3cIe2T+nx8snDY+kvy18EyPab964y/WHK5sf3z/Ces5mzowqNe
fdh4LFIG+RNzoHYEpZXENAM+JbWi4UnXCm++BDTfbEB65E45w8piL4N4JX5B
TO80utAb4VYeHGcJ8sDIDKM2ET2HCfYtHoEhDfW5R44jYrv8Jxav3MEPXvvw
1006oVJ/OnlNMwGUoUrvPC1/aejRe11d5h2pvyNhv2yHcc1j7f1JQoCp8MpH
n7ozXPwJBniOpZmXsn3pR4Sf2dnDNR1brgq3k8j3pT9QxkHVZ7k0WTZsG5lh
WYXa4Yud8D+vYzjubUvzhklD3b1nqDjHeI0L9a54G2iEFGkfBL9isfXUi2va
1i3r08iW0Sqbx6JeQ1TOdmeXgTGpVlH/ViOKBhpY7hg2HIrIt4jWNzNwX2rs
ZiRqqxfyhgmZVcsLB5N3kLYpEzCI9vbwdH7c2iThntTktEf6Ha/aoH/cIV/s
FCxnk2Tp2wi3dkKDfNh58jVBLYZCWUVYEzEQA0YCvGwVPeEUeN+HeTsMWlC5
/7etufRn6lXT70T1c02Gc/1otrrBbPD7lOE0uFSxbdzyppomJZnmMZw/MCop
Kf5AV5IDnjPU+7C7AEVu0HOmL/P9mrs+JO1opPYvOEzavdweqyJi/C3fMtcp
uU2sNfOpYHxuduCuQy9Oh7bU4ZZOgrbWkVQbzl7TLwSMLlF3VgfkEE+ya0vd
fZI3ron1rmrVie8hbkgO9Jvm2DTbqsfdofF24CGY0vzg5N/CZxv/hCnz+NaY
6y+/005ySHC8JnP+QfEyOqw6usF9a6Tjs4cLFaBabX0qQrPrbsCqzI6K8b4J
ZMvaOr6OXLfatAcIk6hZHPN7+ofx1E1il3WDkjZOaMwazCWtjzOiDT+Rb5FT
yjEweU9MNjGivZEg5k94hUa/+FVB11CdLBFo2tMh4nBoiiE6Apa6nUb+RfKr
bMpp7M7dm2yyFSYKC8WTWhiur+KSdPFUoSWC5JgJ3+4H0Gl/vp1m78pTt6jQ
OrBGd64JWx89+Q9e+3AKaHLhHP0mZV0YaIr2odVyC9UZIiQufYRUAPhAPqR7
IsOwsrL07N1t8UhOrrCbWCWwOkYGCyIyioOOvfg59Yv2DyWyT74QES1FURtp
vsXBnOA7Gk3GoS5z1yGyqW0rf6FFBXJ1Hwo34cmb0/c+elUL2PUc4JcMbe/c
zPL0zOQZyhasKPw8//6t5ENzfXGobIab+0kFo4OmmnTtcq9R3lcNIcc1ZQ2s
7vkd/wKowjQG/w5degd/DiIHSGDuPvI1TdcRlZZpPwTYxL4AaGf1lHI6pdxf
TjH4baIHHIK7D66vtb/a57WYW1gUmkXTmDkcOm/9SEr1vnMZFdPVCQ4Jc+zX
QQKi82i6yZEcNwwXetXcWZy10u0zknhojF77Gr1lQQjv9zdU7B930foM8Uq8
4trwuL/sENUM9K5aPGX8CikrNTBNq/P48K3CYT3EaqIv/j/HJea7zmEa4nm5
dDJzaoKKEJkXIm3sGg1Hnv8jDiQAnKL4YeVVcXdEs47ZpwYw1d3kyQvNGmwU
dwCwzCja/0lEsQ/56pV5xmIUHoG0X71A56+bokF15awqquQCqqZF4vVQAGtx
ZlUqCK480m5g3gKRwF6PWMsd8C24rYIFO3JHNddt3cH98wdofltwSHUY4jlE
77QoNyFyfNGyH6O00W2i+235ZhZ+SGsPOvo3tVcJLpw+pOuv3UWrb8GiUotY
Yzt0rVLvrisXJczc19Vf6OF5+k0ZJGc8GjCwA/iB002z/8mPzj3uybhKtCpT
Vic2nGL4HaIue4bF2c7Olga/zKmEvdzSjc9ISPrtqRhDEF3JhLqOOJnXgpKK
LGX6+dqUo9RhPuj4swgVY7tYbaFU88y12rzAlquh2UQ1ypSuIOIRVtI+Cpu9
rX9B9GMnEsXVS915lt2V6hllfrMoL8Kgf1yXUpGa6/6hdy5e13wHoqbBBG3g
GOI49fpFzPuuq7ju2HbPMNW5k3uIMCCImeibfhO0uCM/zEnWBDaBJ3QwJ9bP
ywIWuLryWrDgtNaMff/4J5wgv9TFW4D6YN0Vu/J1AD0/IhoF/2f26QDVCwJX
zPW5mDLLBz7zLmpapXOflzskkVOdw7c5eE1ivBZTHOuYz5wQq9hqhjmVbx5w
FUMv5yHr/RQiOg7oa8JWYzfl759K40vvPRD7va4LGPjuS+S4I9Td71VsIaw9
B3T2IfUruSNeTzRBYVBHa+Vb/yCm1aA4mn6WwWfYc1VNdjM0Nxl2rJNoI6fc
TnztK9dNlvP3tdyd6Q1E5o94GubaoxY0Q4fqLYulaQ5884DsriNN5g+5IIAu
vUWEYWLpQ4+QyntJd2BYepykdiELWDM8VFQtOgXAwRjzF/3gPUj2BrXxGvr0
4Yvm4qpKHoHaGuwoRB/owCYLTH/DaqsJmGI79oMhoMTUZp/gtVtXSSEvqhcZ
d2ypiPqWdqH1plGZeqITyYNg0cv7PdFQwkQiiRMymeQkNzeoIvRJfJDkfYrl
BqYDPnvkZgBHRZkGYNbVjGC9gokADkJoYhsg0jxrBk9E2YlFmnrFCM2JUkpO
C6QQ+wcl8BAvs2mweqWKXp/ZwdOSYhdvWFMbPmJCREd2eTB12/KPNfe79P0b
mIXJ6DDPedhD9suRAYzRI37ywtp876iucp3N1ZZa7dsqlP2Is1Q+Ownj+t7x
8m8sXsMcq0RYSt4Dr7LsQ1qqcFe8KOh5XvKhwzfCwnS/LYSlsz6i8gc2HJfD
FI9hc12Mpb4bW6qCrb/dXRG2pq/UOdy8e+PyGcrFrKr2NgQyGp+tQptE//XZ
AkPE159k95D+As/z8XxhsRKFKbC5yGByW+XOg46wnKSvPzQ0pVzMGhJVpwzq
+mPm6oN5hm0Yc2eOoxROs0Pwsh5/0ltPNgvvs09GlKxwEVKKSE4w2prpV84f
+w8o3C+7hR67zh0q8bLt4gkY0XHpAWUOsungspS2/EpU9cYXihSYTanm+F6b
b9/rq+4bcazw5L8RfTEKGbvvBGA9j8gNL+ai9QtJE9G+Jf5I8AkEAVq2bpdR
q/JpCjSUNAH+L6yCi7vdNRdck3j73vFFQPifMci0BrW34GJgn93UP2EB2WUO
ppUXkozsIQoM1pXXAdaw1PSNRxByq3dDIclfVgexyzWoQgrHr/GbjxE8w9xN
YOLwK8RmKWgLLTGd11f48sdEoY0pDfP2RdJ3RhZxGbaN4xYBohy7ObQClKCV
yCYtDNxE3BpDSUk/5Q7+YirHEqeWW96LDyWUSlttrJQzBshhavKNTIdeT3Tz
0OSmu/nB7pPOIfltKxRv3rRRvPzimSHgPRcr2wXqrpBTiDfjmCeepwiF2LDa
lHgeliFBvc4BycaxHYvtuAW3KN/OnNQt2M9MyOqLcsfvHioqAHaGgwMpZ/7w
Lgn34ERj0cHIl2la3vHekyZpvzk82vglPdE+jc34femXOqaBarlStDP4aejJ
Q2jAVukgqx6ezYI55LEkLJqnKUo3YqxDON7Ok0YtOg1SIGAohh/i8UWndQ7K
aFS4WzGvtBwSo31rNFuU9TFu4fqf/Di1VSGteP7pL7GkGTR7+6JE5MK8aHr9
56OqOxPUXZrToFZRWTRrndhWfqcfF/7mk0j9iIFPpuoSD4SK6zEfOyfQLUCM
jMEtv70zrnVqmLi12U4asLEEdXSXs/kMvy+gj7r0JcP4V9FT7La1Pr98XHuM
Az35nV1bSh074I9PrjQEYv24dUTMJ0sI8k7zCJjP2yIycbSW89jzxcYYeabG
9Q/GYi7jR0M+1Y3iLG6BszVe5H2FrXZmcc50dcIZfMAJBMLv/6ZUxpj5Q7s4
DD8CDKcLYmINYGlBgHkiYoklDFon2Vc5dwsAFVfyL1QfDKmd1dMnMkoE7aSk
UZBpDJiFiHNNKuV8i8OosDMjwfdahKgPIuiPN1uG3k2FNcYF4g1XM+9n4ufU
r2q5eeGW7KJ17e/hv78Hwkg0PZoWNyj3tLv4OFDLdxrCv6iXaYbMaAfMJAFw
czrgi7WCZK/NZgp2G7w2EFUnUmZA/rZ9snLswqZ2sRwGiDwRd9Ba1GMUi/sK
HtLwBHMlbVj5j9lMqezqLWqtfgkWfLNVbZbHHrQo2fFTzZmXnL40U6NDP0zC
7PX/2clcop85mFL1fWA8qaaK4WlrCTc7FNQ4Ddc1pZRMIpGaHlPqbwoeoZIj
94s8JxwvzVSudX8ZS6sYkrbgZQ1MySUfFxMBR6HZbAHJZkC7pq8PPMtRd6GF
pg7esyyDPBf05pKrfWdMuU9xXArt1rKdq1a9G6d0suMdancPTojnL8kXfzeM
c5dC/4qNppU+Q0FWrgXOaw0yfcQ9p3hNiYHnnrp01cAQyRcV/w7Y+DtBKZ/9
h6O6Wq4ANuUUp+AySgif/2Mphk3hobbuVxD4jg8LG8SbW9oNycrj7ikGXjC1
Kh5TYMeKJR1L18A0DUqUkNddSYbrWNk6HhOIzwE7rIAZZfiuLcC/kLRUPUlJ
MBAOv9BMBDdcKRlp5sI4wufvBx1XvdCQ1GA79XURH5rd77iI6uUSp61IRhKK
ne2WUWJM9v28QwI0w+OdYBUa7fn9T5Xdx20xbKSCpT+eXjMu3dgY47pD/D3E
Arf6/k3Y/IjPypa/9jktVyO8lqitLWD9u/TuauXDNTPWlB13skCRTwIZecrT
/RB5n1JaIz18zb5q8guC+HD///qTCa6KuDxv0b9wuhnaxlJUfboJZKYqldfO
sbET/jTY0I1vJ4X+apYtGgX8KkypgOLLhcFE1zT/y7xoV1as3Eq8qbnYKyMb
iYraktcpXf1CAW+l5i0gjLQQQugVEhMczQ8y+vNNH6cpJdybuIxZjs/unT5I
JPayEqJPcYks9+97MCKxqi/9MxuldpJ2BQcaEm2KH/4XKpdCuLXSnxAgyi9j
eLkr4aHmRNuY2hlr2Bxqj/fySRLrF4CDDK5DIA2Kp64gv/3wDrCWVmNdlgZf
HsvqdEasoHxcB4TWSsibWXZctmnmutTc7L8seoJ/E6RQRjCUsA+Mue8fi2TF
/COsgSdOk/6lq6znEjopifHlnaqznz/oLFYl8J5dzLxww17XadGebnXfoitO
YrjjOkn0sWzkAYne9Iok1HkUa1vpT6XXx4VL61QMJruxDLhVXZuFHxFWN6pl
PYvbNc0Ikdm16DdGJJYu/+zDWS7mhVQZgdDiwPakf5PjDXDg+1dFtG6713QH
P8pecqePKudk7cdSAW/xq5iwbxO4cXKjBW0kaJ4U69Uj96aNCKGJ3weUpPFu
q+NR2iei5r8RlvVi3ZJrEHfPPfLWcXi4q2F5SQDeHt/x8Ro+CZY7Tlyrg8J8
sUxWmVzBU1L6KyZYKOe6/QNBYM6ZVFAH6k5yVAlV41cxu7L7Jja06W4MejoS
Udmc+aDEMJXwq/LoptQbsAzU/j88lCnqHTQrti/QT7FCK0+ku7aVej/6yzkP
qypWkv9NCPG99BiZLYG9qAVbo9hHOOzoPM1dn/xwmMwizQoBsWCaecNvsbgn
yZ7TQowju0aVGDY1WRx/wCbotFuqELg6OCuffeUU8vrl7LJzOZiLPFnzY+g+
YIvj4N592UQ6vBT1H5LOFGG8mj2GaqHGI954UtWkeuaBaRl8BXhGqS6vbtx1
tt8NDXniri1gfb8BaqG3EtPPv/NtO0I5iyYvDhqsDfPZqTP8RHToxy9ZUsNs
CiRBNMyUsy1ntl8kA9d9GhyXyHf7WsYatE05rtu/0on3FYYRVQHqbKQiMeIu
zkQLhgHwWo9BMH3EUExphvbhnAWj2npyf1Fx6vS3s1y1eIWR+clGDIZvxc9V
yHOQI9JbY9zthTs0L8bjXcfZ+A2EuCiCRAPbhcA7kpV3SDCEAONbTznnSAFX
CTQpfTrOaFktGPuJkGI1parD0FwSksxB/G1ecuy8eC2aO83MTPux9nk263Lk
jLN0OBPK8zhYi2xirQEZ0ibOWNJbaXyZCH4htFkBqmo4yV/YGYXO8XJinBn6
LIGxYO7vYNcDtsdbTwKhpqpHaQjHJPVph6LqUIw/oF3h7QZZcL1WjKuIL0Gq
aVTIQx+ujj2BMgkgEXeDDdVTZJzu91sl47reTBQcpU7yOYPlUIPT2q/8AAUB
YzWy/OFEFwABkmtxiYa1YUSd5dgeXzolqwdxk24vREnMX/QPA+AGOA8TYySY
3mJ/TS3a26yQ6M2JiwfteAzDfS54QxkFRs984QJaFPOi4XOusQ4nRGwISPj5
PeNXO9TDLHJyIg8jQqbHJW6J/YOjipjEVRByVFphqinwBtf7eiL9FmPJ3/kb
7CS6hCi4EO/WCcHztUum3TEn43CNmBIKV6L0/lXMKxFJiI2k7z0nT0EOgXwi
JQkU36VKboIEAlqtwBjdY4zOhhJKdBblzF47B1hilczMSKrVIv84H5kBguVg
NtCuiNrXXSAbbNqo90gouA0wgIgm/Pc3aW7i126wOZb/UPKYQvjKSymbc0S9
GdwvRwi/RtFvmCGTjXfQIc6kbLtrKLWTsK1Y7k3HwhI82x0l5qfiq8eTJPhC
RglIQ0VLV3Gm6urxajBjOwlBob3tzudT0iUuZSBACfZix7QQvTUgWL2J71IE
88KVUFq0UNQFFk4H4VphqFHz2pqE27dvhAnGLZawnWFkACNSojKmBqpHGMJr
1jcBWXzB9j2jFYW6GaJjaqJyPwhpIPLcSCIaLlrBzmalpEsIjuaE0BaIeB9e
g7S9pzHAy3wCrL2Es7H9ifmoGJVaclYW30aDFQ03jE7yPElVJvVdbAiAQ5I6
90zJtvfEuQh63qvq2gEXFtUq3e1r9kgxzeTgfOnv9mx+mhGrwcv7Jg6SLnsw
n2rhFJ54k55ffK3qD+BIlz2kxeQWaxY6IZqdTLNB+vu2XjRzpD59RzuDIsy5
PZhHxoH0nPyqjRLyju6wGJ5w19Pa4lCDNsIhfmlW79tKoAPMRaUd+KHne+aB
gJ1Ibar5TqE14lETWun1xK/YO5B0WI5eoH5ey07V5X0THt6OjwmIzJ5tHW/p
xZbISAcAutFBdrLs90uKb97vnOHTWgl7lFdvG7sRkJmZeYQLWDzHJspdDOr2
N3y41nlW1m3exqK4emCYs7PfLSXNLxjtkWPI0gpk2XLXotX3jInezEWwpYXQ
klvTXbdFq8GlJCghgzp0GbPN7QI/Ki00IVA0SUqmlcDfzXyYG3RXaRl1uOP5
uy43X7OEVUPTy0+1li0APBIJmSizz+qIjldF/jRc934lVeD4uB+Foswu+xt9
E+S3wNiDCKp9PviqDlYRa7CfeGeuSorJDvCjDDsyOUxmnNczJs+YtmXB9cY/
PGM1k6a6czLFVTkBYi9MoiJAj2GqWuQGfvNK4dWCYWIv0MMB4UjIFGucV78E
WsFF0ZYUQK25gMPQZMr+ZQ8dtELQmeVR9Ubfif2xZ5u4bnvMoNc1ECD+53WT
U4mWzP2Axyn7ZnyQpl4GATanFDzKyaz6OWX/WWAzI3haj1sco1mjYUdA8mP4
CjhBdwr/VT1YOoZ4ihp33fnKAzznwnzu44uKtjb0GzApm4+IYTDX88j/RH/m
InTxwikY7OsR2cTKzXdP2Q3qUm58i0LJGMwkJffRIcUvfG/uLG5GGqicV6A4
ttkqu2X7GwVqhqbz0gGPcLBoyjVC7EKex0F8d+0kCVIcEWxuC143KDEKlIcW
TOPYbUhObH/hr71aLjhxfUqGKFNdvpZXHiF8BPTkmlv94q0aQLMKtm7y6URD
mF/WsrRAVDSeRjjNcIoOLigJS4XSnly9gIg3MSdVxetFm+nzsBjT1M68hZhZ
HfJx2IfwYLl5ZGueUR3v4RQLg2NYkTatLClTDMIOOyt8BuF8yUcDAGftUoKq
EdUSaRvdqZlI0qa85n9oDFOy39fol/XeDUCwyzkcRPapXWyZoEnqK2O06Gjf
HltbaIeQhLm2LFtxRRcSjzyZ3uqBnBjlTg9C3E6JqO9GOKiQFHpHJ0QzuH96
+RLOfsnVIoFv5czizXwfzKp8A1hDXP3odFGktAcldm9Z4zv9jOnVohwiUeqZ
QglX3a6zCRNQ36SXHQC5sdbTBGATF9V9t7P+lFuO4fjpWyWS5YMzu1bPrtV8
TkNh18ahr63p+wKMmuWInCi1PaDBc+QrIvS67MkajJlYNHQf1a6YbwCQhEU5
UXRGZRzey7MUwDR3ugeyfVflyz/gWPIxsYBQV8jspHyIpomkEA+i39WgZTn+
0Jht3inKa/atSonMV+/v5PusuGAM4/AzDb752EbK+1nYObOSXD09dIV4v1nR
C2HWVLkhepjkhduIwUljJFfjQpOwdGXjPmeRxFIJEBdgDaK+RMgdVjaSBpC4
Y5p8P1E+IAPvnBZ1sDXUXPGMk5yH0G+26iDMN7PaZLwCRMnnMVS52ReizRar
N2dqO2R4JG9ydBIg5XEz1YPuOXF+okdrF+qO5xXo4ATyLVzdBlUQwy3tsPZc
5HwGCTatUS1Qigq0pK5mGG1JZEKGj/nb9UkItEQFwY2TePvhuJsWdz/vyllV
mt/Z69grYVpy95swYQCgv39glTe88LxqT+OWjUVZ4vvKMS12milLFHEJxZNb
ge3OXrA5Wr1w5WvyWWdNJBq/OajfPd+6RNteVRQ+SZ1L73TEwhPBNk3eY71T
U8NqMgjQkmh4moY0OqBUKvXAenm0akogi1TKFCtv/q3RN0pDJ/TFw4yYrHXO
qHw4xiDyEbKZnm+G7ZrftkxzycWBuXyDgyufiU+HP+guKnamAe/oTG6xsH9g
jq561T594MYF7L8thnIih8AGibG2cLRDDfvhApw48IT4U5AnDN/RJQrXv1Hx
zOh7M7D0eULEpsHLUPOL1QO5MOhIjjc7w30RfhavwVxmSBH1vl9ln8tAXOdv
u64ioQDguLSUL9x+VAW0FEydx4d1elmQgAStRVJ5iP2etmN+NVByMNhThzTh
5BoaIgZ7uHX+yjCvDVWECBMrQwdFHsQ9/tFjudzdQthYBRUb36Unx8LOgUgK
46WXd/b0Xi1Telx6TDKsocxdUB0Xq2+pQbus7QDi6svQdVwouMInphJCi17r
xrP1l1tiM5Q5mUi6Nu+OdBwkaTIz5x2jdQIbYdKaV8XdTVtN2yfTDRfwNmCk
7nEhohRFvXzH2X9sgBgtaIHzOVhhno4mOBIJcdRz0saDG3gRYk3mniMkMi2t
gB+hAqEWAapMKsLuoBPiG2zISUlZgLXkjHFm3qVLIIgpHmJ3q8sqjQ/kxe4H
5UPSntSo/AwxzNaU348XSKnXUsmpq07OSCZTGyFD5gwSS6QP48tnq48MkIH4
hbdno7V0WrsoAeispwEyg59+GdVfIyYaR9vnOjQ8eJlTgdllUOirgxoatFYL
B7fwVmqJXtimS1BR2TzAb5eucRkKQGrukGM7GqXZhOeLjBviEcH2g3hFllWk
w7u7HXf7O9hykzJStVmoUB8MZYw+9qe47vwx/GhpcLgXcsN9yk9cwjO6thBb
OEmweVlEDOhPRoGLuUSe8vsOFgg616BjoJrYIUAZJZqWroYhRjAAs6iZlJGE
HJBiy1gbNG3EaqhgFOd7U3OWLDbyp5okyrWI640kWYY4XWK8DV3Q1ZFHSy8p
f+ZTJy2rWXYp9MyExw1GgocEJxZwJDsfY9xfEP7j40jDrVQ9nbg30ccAxr8p
fbcZ9EaJQ0vEN+LGCc0YU1+kVCMQ6lSxAI8VNElPxIgUb44p5GZ56qF1dzLT
xs9bsza3s2P91UgR/EdVx6zWPpea2SVMHZbGrGal6oTBivfNi59B73IrRO2D
MAhEuamUGlQo9coZUXwbE/NPe2tWMjkn7lkWYy+iGwvlUxsibhFeb1A5xMga
92rGuViflwrVHL7CCw9uDKMk0Xguy4Vt8xxYvwREQwdLBJqq8Y1mWAogBDNH
okmRTZOp6AgyztNNFC4mthwFFZI9PXtjpDAH3iXQoVNzVTO1zclnzqtTHTVD
mT+CSok9UQYE3ki2E6Itic1mzFFWvNuvmuQK4HVQqHem+q0A6d3fXR+AG1kn
h/GCzQDQEr6f+c8DDpYAoeMeYXmR1zmqlo/64mXHDgDrrGcn7iSrROeeBZi8
WOyY8CqbHiB2UtLbFI5P+EL8cQt+DFSX0RCZz4SxeHjGvbyuQwoJzisXh/Sm
MGIk8MOyPz6wvUDIcLvHm/dS9H/1AxCVg+Qrlj3lfb0dlcOZ0zJ92zqcg4bg
dgasnBbTY5APh6xin+TNjAU2HcU8Xaz1zMzOvojtzxl82Wb6YAB9n8juuk7h
Q3RJepzjFqz+wQ6UsQSxVKgrkhVLXeIW0j3d+Qwvm57LDLgR2BYhQcHGl6h2
rITbM5d0U5cgHgSwDfj38rpDe+LXwnQBJUXKj3rU0mikogzvDWzU1OSb8FPG
X1CFHNW9e+G6ARvhOx15O5MnLO1BViLZyBbC8rQQ4SrGIu0LB3B9SG/sOd6F
q7kLCQrU9Uo/HloVNdgsDWf89xkhiBx9tl9n/2MczL0iMmEOdYJSo9bRvbnu
cgDCg4UDpOCpGvsYePQ+iinYqlUx4MjVMpQnrTVhukjRDJBTBrHX4J6PlxUq
7glgFB+tgC52QgDoRDmi7Z+fPH7plEXGKD3udPYo1Eax1jmcut+fEO000N+d
lT5VsDS0PMmRD72yVH2fOtv1K5f4YDI7QJnlHTBkIcnRon5yNIKov0xICA+g
LbAYWAPx7FLV/17uTys3gW7Bpyq36iXrz7dQK244X5VChssXFY8XD37GUWry
CYXurQ4I2JYa+8d6lQIdNkR02e1w7cBBLQucjhRGa24T5ZXmKeowfPPLBfZh
vYHH3fokkJE7NikOSidYX1r1cPVe6VP2HkjK7spZ1ASkTPQaDOCuZbS5oWRa
1XiNoaDCllTY5ZFl8pF6RR4cfby7oPOE9g3SsUepkZHHVZROX2Vua8MU9rki
x+uwvWUj52F0bJXSLtuStQWuoZ6PQjoY/kAbas/hkOR+uBVFfXlJoZIaZmLV
kK4FEih/ywvoutuGR/VfD6W8GdR+UFTvX7euuoyouvuNoBDnj0iYfrYN0oqB
83qPgQ4qvUhnzZLUNaRUOzLJcZHxGOK3Dyagsxo7krQh/vqgOQWDIGPizL/O
/jDPY7nMlGHRR84XabJ9veQCkEKflBT73LjjvGpcbI+xKj1ESuyfZ/Jmw4ua
qz1+3g+CF2Xq6wI2EcvKgt01a8ea4O42q1Mwjy4EadnzW4pWgI4Pa7nWRzNs
5Nlg3kKL5wJRZEupvkg9bLNw5TuzomCY0XSsqkS7LaXCuXVcC+h3Fh/S2VmV
E0TNCtt4HCWyPZ1UMZnk+MI6mYASmy6hmZzM6ntCThoeA1gpwngJX9fHB/eS
IEfbKDqA6AZyEU5JwXBw8b5uKWrYu47Ciyi1+iX5XVhkeSEWppKcL+Ku2Lsv
hJdu5JRD4155W3wOjcQ7EBxlRBWJknBp9iHzmnessbEUhSHmOVRrXJ7XBPY8
2qGET1pxRxiaPP8wae/GQF7QYabcIhPu8vH7xp0jZxj4j339fzz9WJ0spIQO
JhSZ1akxul1bO/NmrfjfIsJiDgXoMI3sAiy+0CpNQ0qr6qhl7ZNNhI3enZ71
tcVUHFHM7q+IEjQiiZ6Om/5l9Z1Vl/12+e1vdUYaB7+ebGzq/bm23n8ycB0D
/rqOGggOb2eOXVENoXP6RTv9UfwHWQL4Yx972U1Me1NAeg10G0fZ0cBc6qoL
dePmvH3+FfRhlz8zx3Aoy5yXj/5CgMBzlaj2cWHxUK/1DGIqmsRODp78QTST
I9F+AmdTnF7ECCXUNtbSo9FVylhDnR/ncxm6PK3tPNzv6wknTH/PbcFBLz1q
v8JtHyCmefa1DH76WLWkux1gji0qM/U1erTLpZ8iz+D6UVl7mgDARv2ywUDY
XP6SIZcGW2rnCfPj02+XbXNiCEv7+jlxnpto8OfzVtxKAu3pWZZa5cqjXd4S
NOnQTDUPPAA6Lnu+kSnvXp8Dxh4X3qfE440xOKM9uz5DJgahXdyP3PAGspfg
hKsyJRH6k33CiuB9krU935w0l7jKGus60Uyy2BvG49oM1jzoqlnGUSRRUtqy
pxmp0xXd6teqRnr8xhheq9zPQJtkmZcTaQ/wgJBp21Nwrz5f6lVP60Q5J/iI
g2BX+jeaV+8RysczgS+7rfw0j1lhocwzi8pXLfIRaHtNc1pXDr3yoX3d/HGe
654wHpjoUIF8fSN8J1gzs35v3ojlKyPCrZTFzClXpLcWlwSWhZrWY74xos4y
dsd6ufbryqlaOaNNfof+7mvNtS5fzAE/3WbSW+DNiuOkwZeFYwKxG2KeRqE8
S+lxkN34/4lXSvZvxAlqsP11cT5+qyVi7LCGm3ChqpTN2MFgEV9JJtgHyeiV
8dj5Gc7y0GhhWKBSvxsMJhjFLMsCggAR3c+RntVvolSdN7KViCC2kN+vj41D
o2ORD7sdVU/a2JPiu5awZoVqEJoLXVEz/hpjqOMraNPKk9psbX+JllnObKPA
PnYMBTjRgOPe/CvmToleBst5sJklLWTDZ3rFuFoI/00wW4kFvtwIjIauck1o
A/XbD0jRE20cs+gVLeNL0hd07WkGy70gqMZ3e/glx/6x4Gp3fdsM0YhdhXbW
PHT/7wRids+xs4kN2881ShRTLyKBFxL95jjtMwDHBWUQM/7WwP3MzdR0z46W
OlsN/PalXkz+UXGcEXb8TxDTYgPU800AexHybSV6gWqN6ktROrmzWkmH8i2S
xtJyBBnInMoG4bLivI10xFsuZEgnWe2XkwdIUA4paph5OHoZa5famMI+ZTcr
/jdzJrbPaoL50kpce0DCz3khZVgvu4zgPSmmOyLumcWtD0FPzpUe0ENJ1Sec
FgdSFj4CJXjlKzkVyDAElMeaoIiORJTWrsF8Q1QrvFHnTofubKrD8GxU7ud1
CaMpFOVvE/eaARkA0tf5x1EXMibN1sCs1KWazOUQQdEualIN38b+d3lkch4H
uZQOkim6ceb/YBDYC45/Ek+rxeq2DWycm+B80EYhDkDkvfChtPvnjiIN0gFf
wztVMOfOMmHsM/EqrmtyYbP7RKbH1EX6FUP4i+W8LZylL9cQlbLtU2J6UB5S
6Y+pieeKqnt5SrrMRccTxeqvitnxThR7771zxZ14CCG59vBWVAGMZcRCD/CY
DeV60MvW0hDUwPT+4xMZNH9dJsXuV9z+p/c3mwEXt6HQgOcKsNnqeGKU/BRI
/iKnjMsQ2cJStXmXGX/blLHo1XzLU6SkJ1R7E4qfidU8Df31i8zAUWzG7tNE
hW9690Aeop0TFD/onZzoZ8YUkVKHscvbrMulQ/zL5YRmoRtyQXsXghCoGHRX
m0QaYdxPMAxMMuaztGitUBm3ONKjCDsPC4AVW376fA2gYwvWSDuOVT0NnOnc
NPacPVX2SqfTJc17LkOjmdRVOFJasohQ2lWoyr1zQunRZ4MUe063KP30qjAD
GEwjtXSwBcvw+298qi9dIquW/64Siqg6j0lfYCHsb+k5Y5gvRYwEFFmd1M37
dnc21JFg4+CIukqDaA5M3xDLfPuV8CVk/3ysASRYNKY+3hNDNs7r33W7itMO
cJ5my890VbQojb4jKJj/lTGXfjfxgko48bcbafShGE/Y9KE94b22KjEWVkDt
YbLBlDJRw442og2i4LlKdCUPlGSyDdOz0OOzvWAQ4nPgzrBjEVNDFWEWwTgv
3dpIqGiIre68nuukH9kw0PTu1XgB5Uy8YWKM7sNB+OhQXNLkdu03fh+lpd8W
PFNARu2nFjFdPHNeS1toqq343sfcfsZ5ETo1nTS8DF57A4GrrZMSMax9VEC4
iSxYf49LVSUqW4C1xdxB6fxrkhdMHOrBTBuz7r91Rxnh+8Fl4S3byEiByvY9
kh0V3PSraxslBls5VuuA+qg+KIVcu6aOkvU9ed4Fi1b5Z01Z25Lhb0n2Az6T
CGlt7HveJ/BwF5CUi7aN7f8n2JGOo6bH6++lAYwzDHcVQFvR3B8Svwsf0nQ/
mRZDvMqWbLpGIKjxV60rKwkMHB6oPwI76iraqurWEbB4or2vFEjU3i63gieT
cLd3+jP4RB6J52GNtjmH712fUobawxP4/Lvu6dQF6PnOSf2Cyptd3e4YNw4X
RPO62gfgZdajqTaIf0iFAQbAxVXoYqhm48ETgdzFV8qMlxTimVMLJA9WgVzS
ox44TTKavOt/Sf1mAiAcxznFV9mg9r0w6pNFUL+vJU5K88XUiKIVwxXt1b5X
9TALnuS9AuNXB9Z4q8vVxP7sjanm30tHj6h6p+dnrD28WYTPDyuv6zWVVcQY
b/6KKm7Tm62BXpz1hCj2HtzAKAgrqdxjT5zd/Dnia6gF5xt5a/aNdPiAOHVy
FfK9kAQFLKZG33tmBMRdoWWlnBKPwTDwprAwlxiRW7vCQEwCWLGTUjS0cKVE
iBBP9d6EruTVEfmO21yIvEQa1ZM5GFOD7Rjg/do7Z9geAivkdbkHCpUDTwKY
91yCIGvVM5SkJc7dLDcy2mwgxq5OxlSfnXFUgE+K/S6C9p5YAdQ3N5eoJlWR
jNDs+18sVTg4/EX0V91gmviPcFWvceBCa1GZ/P0x/aQ/nl2cQrRbc4zLGykQ
z2pV3N3p8V+aYVmjvtek7puXo8DAg1qbU3kH2i9Kv5h2sOuR536/4n5rw399
yrHOJ5Oqy0u8oIn6g7H1o2xI2kh24yAWIwxyUc/NTSbLbGeaMaBfFg/SmV2t
YGsEPknS2FSSDcgeseXGzQZUM0f862UDtUESHYjE0ZJqIkelFF/txp2nIgwY
FaVFg3zozzF86bp6ey5jbWu8lQFWinkPlkvQsHGnHlW1V9Fq9dkqxCmVtfnt
YiYsnh4pPjEqirkI1UHDp/AZHaTI86/qa9StG5Wd21G0nqtAyXA8e6CfO0p2
ErRyE8gcW7hrhSUJdctGI9RRDDqAE9NdCPHoWLVEvUFu1+nLc5ar1+s0e8ys
6T6jhyZ2GzwnOeQjuVNtAgV1qdVMD7OyiP4NZGcnYSE+T3763or8E5Q3En/L
TjXTMzUbsOWtBQtP3KxIcJwl9r1RuaywAZaB6r7ykizyD1mDF2wxL5e+S+ut
+F/6OclpQvJ2DyZZK80XG9mcrvKECNahst6i5+9s3eflbotqHCBJdRC023Yz
2xhvD7S5LTHiUgEJW7FAUbfSHK4Wjv2Ld5XFI2tZiSxvFVIBqIlv+Dv+guES
DV0NRf4vX6iHjXFwgsnxOjgwz7vGFiXgYbLFtA8lIY/9yii9oSGDKj88Ot2X
W5saYwSRlTtOy59XdYrI9SsVff/u3wh5ASFenI4ayhGw/INW2eQLjvBWslxA
2jxunZe27O9rlqya2SI7jIeest4x7VP4+NwQfbKM5p792bq933x9G+nWbcgM
7lnNjkNZMMFzgS6z8ICoXA4nU4jMG1zL5z3F/os7pPm1Lt5udUOuwbxDdACw
YpKYm9IBDRz3lCQeDRHLJh+LpxX+LM5s0Qjz1KiQKCEY3KQnAPT51O9rVO2s
7oXHTujT4a+xfcQHmsog0iVIkKzq09zQOYrppTbftfPHz5wZs+a0Eifa3dLl
HNJ9q09WoS1UAXcuERPL4GttfHRC/d2KLcrCdjQrdpUTP1uCNt6aytwnTjzT
CYvrS/YwWjAFQueBDSnSUDr/Ca0No1Gq7/pq5CfaL3aQh7iqoboCGHpvQ/ZD
rwI6nVDF9tuujxGnN9Zmq2W6nDFInek/PuFfxpoJCSNjUsX/QO3RcOZ4Pkb8
FwZvpb8V2ai2jkq4CsXcA8BCKqB+qX03nHY7zP07rlNNf/1I0fpgLt1ZuS5C
9G/KBVvz6Vo6MEQsOvxV0KZViFcRdYmblTYN932YirCU4T/9peNMfu7FXt1G
ppVYBCdRyxB27Lu6olHgrPQZ4AdD6iR1FF2euKmcJRzmSdgYv0yF6P+QT5io
/o7mi/ckCMdSTO6IuC9ujDuMQe49/krASPSBSsvdXImvEXcBA/Ny+OniIj3g
NUpRZkEb2+RJjCMg0+BFBUd1kzendrE45l02I8VyM5TymC0f2RkaEMj4A9wc
+mBJzlSLbZfmfTRuPDOvWVMcyjFOZa40zMlgnS8VDJiwC+DGmQXDPcWCxvxd
5SNB6i8y0SS4fIwVGy4zirxyDLw4slJasJfAqZFMcRjJt8lG+9fvjMrU6jys
02Ub4hd2ssiqnBFujtM6ELpAwYXbZdlMgJIhs+kP5hS3e1fEvkw2nYCrooTs
GR659o2iaOQ6jeUCLLxtjqHiu1/TukzmoROpivZ6yNT+SwmhhFSSyVh3bpyw
5MWDPaZipq8ooncmocAUECCtqH9ygqt3ZC/mzhlaTWMFNReS+DiYtt1fVQ8q
2TkNbU065u/UvEUChlYp2IcHWdOaC0EpEcMnxqXKNHpIBx9Gcnwqo+wPFg5c
u2sv4kaEp6FpMt6pzTrFqmZD0st0Crh0G3lfPlnRfWIowP8/3ErNNeHdt3Yo
v1Oc+BdTQ6hbyYtKJswM8Pe6vfFjBC7rPi+y3ZqVqVPwxG2ZMcZyP8UVe2ne
4ic6Ybk2naST3ZNMlsujkjjIbhsqs97Xe4LzjJ6cIQVOfQINU3SI/Fp2Dp7p
iD4Y0b7NqRrI22OgkocvYNjyaVSCs626XA4kAHixLFIJE0YN9NfsmYXO5n7k
eLydAV70uN3+Zzj27KfdjN5mQBVP2GZZxpSEZ+AcIhkss+7jsbqll7u1wRah
JAzbtovBhBMLKCL+8RxpWbmGvN9waQjBTRMiTPDxYEfXFz2TewaqBRtZtCyF
q2BdCqecjlxKclSy/rfJISn1UKLSKEBPQKb1aym87+oRt8Wpd69yRMqQDpF1
9A6ggaEr7BoFo7BB/2f9F2AWEWB5OFxKDZCbSPLfendLFy3FEzTVT+ny3r27
2WT+9tzkJCrGtS0Re4Y43ORjaDyWeWO6qKJGPBZn/M0sVn+tvzx/MpKnkdM4
C/Wn2e7JhXewkPQekU8QHU+wcggt6tztTvS5fTeYQSnxxKFmlJ2cc//tpLNA
+Zlz0Rms+45HLV86N3/LZWU46fEmvdN4iMW1k+a3LojmaWMWp2CVNPWn+1qI
D6R/Yt1j1Oyn+96X1/DUcVQUtgg0gHq1qRUr+rVluNJKI0Z4+ic56wcixQ8t
LESnLy5ZfVu+9GV5fbhYreg1/rfAIOCojWP+Y7NVcXGi0GDlmWAZQL5bVaGT
VX493ygWDjUpIgwu27OOdKBIbH51TRcERTjCsh6JwWxdSplCpoyQrYmYOexq
OktBQJrl3huEfmJtNIiK6kvbF9fFNgfgR6E8pyJdabmlhFUiIPPGMz1jDS7w
rxsSgfNNBf6zQ/708XDArgQkQrYDJYuDIho1VVoLcAV71tdc4Aimok8r9c/x
qDPmmgk/bC9KOMG2aplS6fY+zZgMWwlN4ludXcZEhaWZjdwSQ6K3RXDcmtoJ
VV+kRnT+SehnLGIjwfekU/lkf453msM3fMDxd1pF/eWLxkb5oet8qExZGKzf
cGz8FI+IVcGVlw2rq9VuGnRnZ5SgG34jXH709Y91Jt+pXtKIYNd5QSoaMJbK
nQ1VdR2LvVqJDD0SeStf7M64sY8EszQa0SmS9fDji1+tO+aQBOFMG0vEFPBH
cRSFLYEy32/CfQCD3Kcr6/fnhY0XjWslpoiFjRGxo/kudFbgDSAUoygs7adQ
P5koS6k2LjDV9F+zhf/VwWFLihY9DgDmE4khiAEigPDr88xGOGwzI3gPNxfT
wWxlaEP8jTu6DD1M3BPkV6rOoQOCuY+IuVtQXDzXHy2y54G7ztzQCtrTLV5L
G/LX9Al3k0370XcKiS+yN7CPVSLZzvoXuxo8N+wLgPfNy+d+s1i2zXJWgGGJ
kP1aCwUIMVLFKgTerWpzGmuVTzpqQvCfPiPXrlhtan+2U2vP49B+pNsm91Qm
jdAOjzDJtOdi7bkE6jUrzccaOPGoUyamMsGmNV0I6tKZ0+lpMmAnGDi3OTSB
bWegLooPoVJsREc5snaDQeyNbrcmoGYF2TrsZ87oCrO2D89SW1z5HEOpidLw
/Jmcm/twNFh6Lfuck3qr+vK+pH/1k64Egj3Y/csqay8GeyBK24x358iHgi8l
k+IWemKZ+wKywS48foN3tzHAMLGg9b1awRaZNWJIUzNkPBDUWrcxhLcAOWOz
NN7ACExNMFlupVlpu9dtF3NuZvc8IPR1C67ZSKOC/FJY0OiaY3Zn269eVjGw
qJkGKlTVjDf8oz0a7n7fyGwf9z0Hg8VSCWTaTCu/8BlbtySJPw+wBbkqR4wO
a28kKCbr64DU3mq0L2HvcfMdxQkoe6EMkRno+wi3+UxM+1YaiaQw5WBjq5fF
kAjf+0guDaLPeOG4tCqDUPNI/+yfYAAwt+iw7q02IhPSC4NtXtsNO+XcNVgf
PucOI5WT5tN9RhRfcSZ8rymwPlDwnnnhasNTo2hVY43PFQQ4rm1SkBzq85LR
EOPAcJUEZYantjNGOjSS8IjRS5wZdqwESyiU6RgNSR0LEvAW69qUtW0NZ6iz
bzjwSQci9Gg+fzr4jL0w5HproHTzIyw37cCAQWV1Rz4pzjJhs5G3iWF0xFkH
QBYTtBvgb86MEDS5AqBa2homHHGgYF8eSYsSUQAHzU7M9oKBKml5NRB75Me5
T5a9lGlHQNk4BY1fLqETq2atsL5BsEqosRSzQOS4ro0TUoVdJTheknjxbEJ5
EesshAfAIxYh83heIbsVxWazczmVCZriQzY4hU77R27y1+M9Q0QiTxmFxBCU
XpnpIduq6/SR6knWOlB8kaZu3BfpLU8W59iaZ4exx/s2M2qKcu07pT+6hBg9
+sVQHc3Ud8A+calB0Ju5gVB0DK6v8bvA/vmbe7gfPu3bucZuZoTAopVsXV/i
ixuDKsyUsT/BqIvDCLN0PY6Eg2dKcKPNUr2VbKVhUU81yqvXAh6D6KeRPbhh
KF8GK9DNe75QVqVAXIHpNyogMTIB9Q+oscGtrWNs1CENaaK6n5ZSH+Km4q1R
RvZR9+bA9P7ymwl1yOmqYttEzvuypiHzE1xYUEs/nSH8OfZCspYrGin+bA7u
FOaRmvfIgeCtPRhlaTkL84O+gYY5kURld/LcaT4Nwdz7Yr7fqK0zmLOe43nD
bIHKKlL76qD6Gm3DRlxlHU7L2/5HBcTGFERy9OzyI8fZdSHQzSHwRSIuy+M9
DdyjnmEsDlgKjJakHbna1xSkMC3AyW+FPbOUsmwakR6aYwrWyGJDwnr5UD1a
9iQeACpZzog0LvMrkIXORvTlReZn0+on62ZefgMBYX8uiCxVdQuZtbkixEMs
It6YtoplVdo9G7Mm92hHPRIDxDXAyXx9MZGahi0BFJE6lHUpfqbyDT+rXFSX
0bgYRwnxDa5jLgg4ewfN7wMVi81Wc/aGxnFdSS7GUzBsU0yC/7Aue/OFAS7e
v/iGZL2wPP8+lpby2SMdXFCqVzk/5mNDOVYitr4LQxeBuzmPCGk7gSX6h7MJ
LpoyzRte90SY1s/pnn23bezfFCcwFCxagrseIPreEeVSpxtcw1vbqcEljZNy
Mt5gBFz1JwCQbYtNY+Fb7ZKwRhDfLWjpyfEuryyAUET+N6ZDvuQIkZRm9ZN3
J/YFmtApsDOg5RxnuSdzl6cp/b8NwvVAs4FEVaFG/H3Vt6XuUbtP2O97l10w
iGLTof8QWo+KiCLYYAOsd59VoEuUWpyW3A4yg3GYKqY8oT6qKRvLozMxYTDd
x0DlA6+q23K6IAo7YCPo/0GMd5viv0Nfkn7AjZkU/LaDG7pgiYawJ9bLrnba
YvGB9ilSJkAQLOoK2WpL+xy8olgrZSzBOfgAiMTJkp6nxYnsNgcb+yQzM7OZ
y0P5Roy3PTfaQ+I345WBiBGMwAtW1L4fAFt8VGpvfrl2xne8AsMVWUDNoTx3
fjaiesYkzVobLxifxzbWRqvHnIn6QqgzUkit85jnSJ6URGY7aEJkD8Xt5ZaJ
usLX+ljylgQS3Dwgdkd2wlTBL8J2nTSpnfvFoitbc8iSTYaIObssyUbMc0Ln
H+kUdjSIN3MrjYQiOCt8GgIw3oWuGf8rYqz3NNq/D7tyRRmoS3tajN68jxCb
lqU3XlfPqTdmzRHq8GzCkyd6zucgFlxlE5L2Usx6IzN/Ef2XN5nR9iYBUZv2
LZfUSWbIdcHYWRDW6ExI8kXAENKXbyDjIj3TL8PahqHC1Wt2vuOMCcrI0R22
KUtuQTVzoAi3pY7gX42MM1/kWU63CcJZG3JU3odzju7t41Cf9A8fhdHlLpjO
HqcFWSMJKoawSMSDTEibBfOtE/Mx1tJhseqI9imkZE/jrxEuarvF32kL5N9P
zp8THfuD6UHo9KGPDduiqeNWJYySForQpjShGgThD3jf4qJLDXVyZgCubBCy
lCntuFhGOV5NBwTze5EGcmqKlspGwgJhGOlq37IaQHK3zCSXWFtZ15Jway9D
Trcnm6cUZcIuGKBvrp3TvaEW+hq1ANDpJvLGFH308DrVwtQs4Wv7uB3Xspj+
29lDcUKox6gViO+cWgTb/3vXn2MUPOj+2d/dwf1RmH1sz65ihorlQS0arOvc
ZcmkGM6UACuCHdBXW7SiU7/TENGcNceeLWnDkDFE7mkduvUJZvc78h88MrR+
mGsSaqOx7iUq1i0CfsBEpWzNZfjDHEF2rePfVGzdH4Hl9nsyiHaa+fKE1XWl
CdF5VLmsEc2fepquRdZ+G5U01iCyUjkPrG86XyVR8ttwf1tStrtcImr+OKl0
1wpT5NuXjFSFrMmuJwu7jnSG6eQDY3lIXx9kBRvvRdNkrqntjCGWyxjt0Y1R
qsCvDoyCZKFlnY+aXcNkkyDUv8aERfvZsHUY6UxBneodqTRP5FWtkp6cRxy5
rv4bUW0HNpTl3BnHw9zS3isJJmQY1kKDOnFKmOiwXT6pqzTKQYjdduTuwwGm
CAJRHex0G1X5Ew2DNuLWbYbDijakqYNU0UnNaVtjZYhi0BiiHuPVs2AzFsLh
R5vRhVKmc26MneDg1ej58t7YylrWsQ3pOqfX2/uFz+qp/QCqWraznSkLIm+w
XPeq6li+g6OgbFfXAZpOei/1nyMfQy786HdPD4gxaGT/kpAFwL8b5GanuuH+
0+yZLiqCa+0F2hSlqDoWG1DYZw+I6HTFx6LIHs73Wrhov8Pjr92jW7+D1VAY
z8SkU7ibWd6tdAyKwf12T+CTY6dvM2/bMKsJuzT7AAcsLs/J1YKSymyq78kD
lDihDixRsTZ7U/S0JYitQn3hLHoJCtL7rYq0eWRhEM5f3QjqJvQ8cFOONAq6
G8LZxlc6Ksj0PTQ8fVmzK+F7P2vyGdBU43t9F4nhsGZkB1ORr/o+acduggKY
+eZI5rYglErBqZsm3To+6CGBTvtbeSllcjhoD6np8M9T1rfYN8AG/3+C3gdn
KutNzj/2fUuR47BaOSepgG1r913vkaRaM1SwPdwpF26QpzcbjSRKAw3+DnbH
K5Dx9ikx/luyPfqud7IzXRzZ+4K+KPBYUw/7tU5ckTYad7FSbwkqGh5Z1dDF
bmIKwbFpGva9kG5ga3h9tLz9Bi9gevufdnIXyF7rZRdTXtR4iPsoKWm+1vEg
zqbAQRHnCAt09HxPN6HYUK4Kzu6KeTffZr3FhZ+mQipFlZCLlFfRlUwLPb7L
DnkQivWiOQ/hODfL3Whd461Ngi7QROLt6BkPhQMaqtTeprPbW72rpQV6w7CG
cSoUGT9wmPW9CxuKSuWbOIdubAHoW8BM8CdAPlIA4XWWxLRxriKKjHO9tmQG
jIW3GoPS5IKWhaQSptfVNn37dZknamLb+IimMznbnOOo4dADJRusJOnecIHK
SY4Cln7AnAzPZUPGSJv3B9udK3do2/gVwVpX0ZBu65+7gbeGJwmYzesLyxTh
xTZC1hI7V6wWnfRWfqab0NxcFR4XgS+FrhCozXesZVeZumomsTWRjMYqH3Nc
UpJBB264q+tQZsxNbXTwK2Y/stPpUv/JBWrp28slmeRTtEAejav80geO5V5k
hMP9RcfmEN+2XqgZ90Q0sg9VrHDxGtPK9ief5xww7OKraoREf3DyhZdgZmp9
khX21zboGlDKq11L7093nANnXTktgK2nnSBA2M/r1/rDJjwYicxDova7hmAC
CPpFJDj5mA4ne1PkJMMGMxjBpsiUMvdlK4eKnUflS3tWjaQid56NCoXoN8+h
nRl+/U1Ey5sePnlvpkGFbJyYHwfatKyUM2O7CPfWInd1Z2VlwyK6GJLx4qWh
X7lqr/g5vZmySkattd9p57SlHP9KlgmgFCkrGftd6HhB6unIXMAdqC7w8x+S
Hl04aml3buGIpMIdgSIpGGhJxrGXG1qCYyC01/ZIuZTA2VliWM7gC4dZYNQH
ajU/A6o7NRRN+S2aBJ1J+vN3RFCMj1SpZZkuEYWs79DfhH3XwIgudEAagSoA
VFVRuN3/uMin0mDONbJ+TFxKUSBYS7AwH8Y5q8ScLHPRiUdlBE4MYQ0J45e3
sBaFhaUA57XKRBu7JvYE5HijHTAFNAlLUXxxpzHSEkiUpJcR2MG+yDADqGQl
+hDeORbYSWkkNRr8zoVdQRoXa+1jsc7D3c2FfGnZpb8UNZiqSwHH6jmHWZuH
bZNnh6rUsP6BNtOlXxKi6tM5epEQiticdE+m3vsWnvVXk/NeMf5p6XNn+Iep
X83L9Abv+RHW9q11vDfzmYELb70skGKq/y5AR9sNSAywY8Rx0LJMmO0uSy/W
lpy7zmc84EWhuUdEsQ3FecmJiO6ypYT3qH0l6UGtv04ZcTIj2odcKRx01yW3
bOY2hMkpvEQoIKxogXua3DpupXB2SJUDVtLkw6xkFo+xTzGeDSE8gJ2XupzI
cGlVTknWlntgfgKCcb9KmyK4aVuV8cs6yHhsW3qcbLVKZH33l6JuaJPPy4Ab
PSVPeXpZ6oR0Ty2Yg1MroA7LEmurxhFpBYCStkS9c204xHwgyF69VLVDIzRj
Lso/Jd722CPP2cdHLfF+MlsTwjaxlESvBCvg1X7yPBthuBxS+U92jqn5GCkD
3S2A6yRjGmeNp0Me0N+xMVkrJS5evDU7nKonVKRCZhV5dfygjsc1ACHQ2CNQ
7Smq4abSNjl4Fhzn5OO5kv2yJV7KQmZknO/cTr6QI+vVfizYsKs11i6xetSt
LDRhgYM4Wfgkb0+43oKNxl5ZO1s/Iu//0S4uOCTxrCmBJ5xS8d5ZdES11WSl
t1Tkdl8Fp4p5Jji0Vf3tKL+7edZRZBfP4nyOTKsZC8QMDLIBOOEk5A0vbnxN
r9nLVUY2B3AZV8UtsOIpQFAzcZ8sk9zFS7+2vEm7UE9YETR4M0mZYUaGvQaR
gQsZLgqdxvmJeZE0zKISdB7kdzZvj/D/hbklU2cqrX7VLl1L6x9JpNX4xoh5
Yy/hUrf4+9KU4UT54q/A/vV7hO9OfiiU9pYJMWhyCFKeKMZq41F5DqH5rIY0
wLUdNrxnU+k6nDL67kfzSUtj0Egsu9jX/uzxW8jkmdUVOf1W/FXg2JvOpkxr
WUDcPD6bWW3T/g2boEhxxC8PyVEYFwJ2rNhSj49lXY3BRWSgsBcF+o1P2Shx
wa5nN+CQrB6LBN7fIsmj/j4ymKX8ZkSOVRt+XXzsN6s+dxpolVJbV8+JOG59
w/t+cRJABAkWXOuR/+tUKqAdvISC1DbLBaS9X+Iztqto+yNdCOWHif6DBxfG
Ld6cIrEvlJHkg8Abi8mRoNWk6tVTroSWzAR63Ou3E5GKsrrrquzj3onxHbOQ
ePqcy12Beca9UfBYvhV9Zjx0SFN85wtt/bkiidIYgLpOVZSz/Bd2sXvE9BjH
0SsKS4YpEpTJf1awxLiir0Qwv9DE57wfXKAOe24plGvl7qcTCFxzxc5jVJmu
4CocKkzOWRMB/Z0byMOt0bIR3UDY9S8GV2nO1YqPEgn7gCjxHQ65VfWmaS5k
79i/f7YLuXz4OPXzrY6NamgTnCETuS2+i9k1getWLOLMMCNUIWK+RLXNHpcB
7CXGwoPrSleNMT8huf/4NH51NY3nMmfg1D2Y+4qBWuu+HV/eL36XARNytdMT
FQPUrZl1dHq3PvCLIJd6Q0/dQc16vyeB+gRYBauOlS8okuOPCfE9u1UljIsM
M4TCkvjwkAB7dFEIaChTD1DKDqDZ2PAGmsyTf0IvlrwlW0WZSA8ajjd1oNyA
jt6Sr5ZiM4XEsNtqOYZjzH4IE7tsKHioxwyC1UwU7FcEFxF8sFPRZGds5z5o
k4/pciyIo4YUK5cQJ0HatNG2kT9agjjtgeZyMMGmjdwObNFVrAHICFUTXWN8
03+sXfHFILV90iliKSFIsQqIPdcOAx1Jz5Jw5V4ykLpITT2XBNTi4IOYvg/V
gM/QE1kZ611ea0FQtAcYy/boMXHfHHDXrAqlMU15RlBNjGvJNZC1eOgRLEiU
7o4r/nKKqIPcd1iAbsw774Gqt2QiBqefxTBsDXxDLhGZfoZFhMCCc+iHp12q
oDwpNAb+Z65xDpYQC8SOFVilxYChW9ohu5VLB8a/8KmFR0C77AnsPYpE0Qn4
xaJlXWgkH77L80JRqXFqtwxtRL4X/b+HtlXSWBebzsSDbj81sj8yJIGHdOa+
P/iUUCuwAPjRUymF46IcycZAJCcZAJofFyTP0yklbFoEkLMzgXN9b/HtP4Kq
GzGPO0AyLIZ2T8zpjtJfkEYBIgrQXlukfdYQGYz39MLpQLQS+MMfdzi77TI9
IC+2jZvyrnWXOhOoWIky7NZP7xVKczm1GkZipV2/2LoGDxGNDE7E+bt0K7HN
vOlnE8dklTQ5VRmQgNKIf+JmQQw8cqJoIvZhBKL0ERaI8OZk6qleWyWdWKPV
rzzMj+W2+yXdFe/FQNQUdM+PAdfRo4f6+keb2dcnBC7wunT5nKSwtlF01SXJ
31yr8zdwni4wGjssbpoKpCkmSDaZ3AyrRDCHV+VOgXhC8ckA0KLjE4tzoR+v
GRwnKDpf1gpCfKgKqlH3oEdLAAtD3vd29tDsRuA4vAATqbKQCb4mn5eOwP4W
wxvPpi7zWgHNTzXxp5z+vY0wwBlSlW21TV/nWvP3ZY3XdwxnDcbLYjIO7xv7
V0atvzMykgBuDWK1A9+gpWSqqF3YpzK+d5DdXTzrlyqW3dq/mvk9NKUnAUeU
NiO7jCUkg1REgHw4Z+Rj1n6dI6mVne6s3MSZCUOVpOhwfQoo9Ra1JCa5yg5+
+SAFKKYt5cn0fxOc8jC8s+9+aWGrEApm4cR6nWUpfeVGVcesN1uHjbLtRy5x
q1JCoyuqVQWrglFlEy7EUa5jedUmSFX5NvUAoin2cjG+ObHo/bNg/QH93H7Q
ln6iKKDfngRZsflMvOu4M3cBK4/rl/wYJlFJTwB0qAbXtk6gDkycOQBumubD
nb8T7Ik7mN0ZTyQ1bvDqPOGIVpP+CQol7T/yNgCXryR3X3jcNzgjjTxan1wp
yLD4QVJlYrZJdO6t1fESCRQBnhN4NokYzN5pWr8GFWbDGfrsFtST9SisO3fK
3XYfWbJTfOgKjpExc4hbqyNbkWFJzU96veQPU5BP15sQeJzj+H/CpJGuHz+O
wQOAJZ2VIMa4+8XzRHiI39OGXIYM/J/Wkl4nLjDE1xXSp8bKltBsu/wq/0eM
fl4WDXtGNysrqPpzVysT2yFhtg2zcG6ZFkUa7rO/w7TPhGI4UY8wZAAVN0bO
lWloGf1zQ6u0apetOcVSTcD5h53EAEqZLER0E1ItHrxTVYb4mDGkqQFYGcfP
zsLEqLNrA08gFr99oyWv6x8toAUFIyWpuVc7EAizIIOAsRR7Qcw4dxLZLqUm
o3I2KFeGjzHn9SxV4JcRs9Mq1wHwb3VdWjcHTaPLhxjyUjAxAhGI/iSmn3sc
S1CKUOdzw/gfKlcaQPHVuDr8wmbs8jp2P/nGMXPtVyKVwPKGWzluLvBoGEEL
UPlmpb4rxYp0lCtM5ZJ+WFl2j39/c1aPK4hRUo7S4W+R2+9XXN9L1AOgLDiE
PK5LQ2Lxntodd3bMB+t4Ca4LisYJwMIC4pAaPxDDXkUf9J5wliDKbmKxCT3p
eOfu6cksTPg9bKFNiykSyipgt3sc4hMTxLC9MRcwxF4rbaQEL8H9+mXTQLLa
wOl2n+p6iPy/6+K4LkicDTxJOTc+w5DfRyolWUHZhLjld4IRHqk5eNgfXUk8
fS8od3Rs2B6SoqRnG82culsQvrVizKkSLl6/it7szCdmaK53x7b3/sNIgr3W
q0IdEuwKbwaZpRozfJAsfuh6G9f01cBLQVU2v0FpJp7DQyslGOUcAxZHJP9y
VJwDli26QUZlYUsLZEXja8OxeH3VDX2Bh5nYWGklfInJOw7D958netwhqfun
oOQzeRBjYGmUEWK2fynTdDQaENOov7+4XspAsI4qS+/96xRSS5IsoVcaYAwG
AUa2D/7y8etntvwR2tKEGIlpBSezQqlPK+cpd8AwBlMIqSGNmgooeDjMzAmw
IGCw3o9mCPeYcMTNIeXIoS/HkXlyz6KJ2+bpLf4xy0eNBhG4Xw1grqUdoTc0
H4j9kONZyb9b5BAXhDvRsRWS5KdsjGXEdU5Fx+Ez7vHCuIHabbmsECS2+ily
J2HdH035db1yhcXhiKfoUStHpAEfckrxV5oMR+v8xhKTfgnH9SnLzLVXQb0e
O+UtLzpHwwpcY3V2cLwUbDJQEzdD2goHPtO9aztiEJZMMqzVHZxE1kOoJ77l
zxU3TOh4E2UcIughkeEIBZv8QkqabHk9bXhDnPqcr16ofv93npEeLbpbx6s9
gnXEhicg9URzRIrqOVFkVh+peajVmd1yeik9CkXxBWd4waCkLURYBE7Ip++a
Rs10HMyrOWtsiQY5QTfOrnsTh7oehST0QGmeWyn9bEIkkQ7Yzp7oreKFCY8H
dGeB/jAOfyGX6E8Wk7B5N33ElEIQ2F7XB9ksajMlYq0g9Ts+SDuDtovmllWj
ayhNElEPPR2H5U04apAlGb+0IMyr8v3dk2dY6O/hmh62kjwxe7wYGnqvcldA
sIUoC1lLtrwm8+MBEYY3hwuQynz4/91JwIY5loy0oJHg9jXFvpEqm+cKidhS
mC9kll+ksMTjTRm5HXRUwjknbjxkou5rniuNq+YaErGSU3CTvA94yeaX7IGL
uBvW/bsgCdy7jVuOnPiJneCSXQqkLaQ3z5rUbMNh4P6hBXjqbuuULdD3Txht
Nwl9ZhK985hHoeVI5XDrSGqrwgsUbsUp/jld3aXBDmQdnFHU1mEHvz+imjfh
JDqpGNtSvN8zzO4iGiI+3k6ewBL1iBbj/NRI0dri76fteqadtYSeU6zhAD+Z
vsMgJg20jYsS4oZjIFz93n2yaIZY/tMQ4V1tgpvW2i+0dI6sHifkzORBS8fn
iTFYfx68WeTb/zgZOo+Exdl3rixN/+wvLEm4GBVO9Tf8uxgImKis+8zKozoS
MJkSLLpdQpkxEVaJuMW5aW9pquZInnzSXL42J9SP4gWZSN5soH5VF9uxYBAJ
iZokaZH7Hne8jX4xlLshr1MIoSv0sq3D7o7vaJShRNK+IU1VJLc16B6ir169
WiWWuBZBi7OAg/S08YtkpwKI9tvxKUpM0yeb5H/1+X3qBsGVt5ZbQDtZzxTc
i+YjYP63xf4l3wCLthhh88BcQdG12it4rA4jegHlEb6o+CVAK+Z5NtuPDPHp
HlawHLU1zZTQFz4ftnkQJr1egbzFis0sXJzJb9TEIYNpvaKE1eiv2o8onyts
6zUwfGMc6kDdvmQdPInV0qnmZFrw+zq36600svwOewKVNKfCs24CL8FLKWzL
JzMW4UOegI83ZJ1A83WHjXLj+h3D4D9c/JRGZD3oCYzP1WvKnSHI20ovRc2M
YrWJ0IzpHCol1QXhNR+HhG5BXpwQ0ZDeBCY4409tqeR4c97VR/y5hmfWnH4o
i22nkTe1d5rt5Ywl1FyVULOwmsPJ7ya387MGc7PfM7frxqF//hYOHQij69jS
gVQ3c2piYge+CcEmS/iJBjIew/mYKVzUvWxltwf5ctydTxCHnWZ3PpoFw0Td
TJe60YhZT5j95aNkMM/xMxXah97NFsSBtClsTug69nOUc1kFY/0h/NJ3pIGt
SsUFkTv3nkegcshgmF6Vnh07Saw7p/6qkbZBUyFXhvgjLMM2d95zgdUT8GTj
miDOHOSdZY46aKv8G2ErmBbeq6EUkv4kOaFXmzV7mSXt4AkT/x7Lo1kb7/rP
MqAfMf0lNK4ApThmUQJRcuje3WvvVR2IC+Ot+UsiVlu31Yzh2y6aYFwX0UzM
GuKpHPQD2Um1A1BQuqvkwO8QPqrMcGvyzCzy4s9PscNMRAZqTe20b4BuQizE
NFKErWQsZl9h3Iph/QnWKxslBZjkfOx3CwVbjq+JLAIOFzLsQp6drOoYlC/7
k6bPLGiLUMfHCdnSXKDVv7mUgJas2tla2LvNCSZKM0ng6meYCITtMNVlVX7R
Su+7QLaQE90uY0FdsZgn3ffSJVYByCo0tIA+CcGr+0sQu8OPt+k/7CZetUi2
FgUu8A6L0WzMYmAb+Oxc3pSUihhhsrP0w6QzAUBXnoIxszicHdlacFihiGbw
mqpH5OJFRthRsr9AtFO0FxJfPP8vyOWUaPr7xjmCZjGNsKeSV/EukCj0uGnM
/6ZujH51+GzJ2uE6wpee4U+ydYRxVzo7j8GtROjljiEEdaveUXpTdKlyU4pb
hwa1oKgZ1Rr/zOKvwZjsW8C0/PNz/cfjXtfIjfv8aleE4fowiR4XQmuDRO/i
Iln9fl4ygAPIAhxUiyFMa9bypMTkd3vZ9a28B1qLtIszKpjV6+keQxn7c3eQ
3HnfK4j114B1tXyeYYkA05ktePiUKCMf6snHeKYtFFiG2WOmCfF38Fn2GhQi
I3A6C+QV1X6O+TAbk0dSKSapXub0S4ZQjzllR1WWx56L8XAyorhg3F7N7Di0
XYoOrpGpgbkUom4R17Lz/jd4xTgaqRhf7vC2lgEs8yYC9QzCP1tCG64YPep+
JLwcuaZmqDKCWbWzML7SHnircrJXeYlPYZH+fv/tua4Rlqyab/lTGRVS7joR
yUchtNzDpVEzAXDyKjwZmN2z17FbcylGlV39v1onA96ahqd1GDO/QzU0gTNS
4rRwN9bh2tP8MsvBAipgCrMeSkNjJ1O5BVh26J8d8dt60IIvWeSkQJmQQM6n
i+rL46nwHysyJqBaJ4oN5gNYJqMYR6oTGSgJXZnIArrR6QFHxEHuTPbvQpe8
j1Ifk2rHQsteBqHAWWd0LfWQxcYcg5maYN3/VdYlw1WV/cuRviRlqg+s+AHM
EvB2F7MufCEEayNC1uWJwVj8FcCX6FYs6GAK0yFnKz5pTtLSsep3Xj3JnJvA
8aNA+hyf+IJzhlm6xVTZpEaHVg9hrQLmCMEg9MhlJrFio6FRL6C2M5BQ8Jbu
/TaDqM+y4dg1hubJ3Jihsuywu8P3EJWDO4Oph4ywdpe7kXucrCCuV3QU8GUy
Ttr3Duo+n0X94erS06Ddmnt09P4KnOzslnYSygUuem+U5Dl/Yj7Btv/eAHxX
8uQvIY7IveLlpx5bsz2GtlfwMQWYfuD3yIP9TpLJhHiAcpvAhU0Q16HHbdjD
wre4ez9WBbI7vvVgEb7MUVQd/bJvY2ciCh6N+rsCq8MOidWWbtYBNwajoXTy
5bL9Ic9xcpg8VOOmk4MhGSQtTyfuMMACe7jV1+J94Fnz1NIsSSsz0NSpPVOv
6WPvzxNCqtQOaQ3hc4+qFkuBzpp3R6BNFkzev4C1b9QE1MmVXNqVFjTpXnxh
PMojhYHMDYKavPtC7AFWoJT86fWgsMn1GkFOW3CysfgjyavvWoksPufxfjax
DmNRlZ74MAQfwaXkDnwhYEozii+6CCPbXlszh/oUdmoyt1q6L/FAr8EEP9bC
JcDIjMreSPXI+gmftCql/B9P/0lxXjAdR6RWGb8TQBPB18VW9z43G34xJKXj
9IPKtGWR1z9aW1mP7yPzhec9bjBDZUIClEDm2sEeRt8mdem/c9JHlE0NpHzH
nJ5j8W57eeFVWSJ6ydS1KPRB3+1nba9a6ul9dOzw5Ks8IjrhnZv4o3S02GtO
L+7s4lM0pqJKEvheLNenRtKtk2Go6yjqXZrVr0h1DfW3Q8qQd7KxAxVQlGj/
BlDafihD5nHhRWe9rTBWXtiuCbZJmP9E2BVPSGZ5mpYV59qTQpjB/aDEylGH
m+45eWOrlTJrgjwX8i3n0TZ/7k28wSq3Rw7XRg1bFMjU0k7RaqgNbIk6oPiI
+faBK3mM87RQiCbit1zlY9jtGcMZ8mPEslTTx4vz2hRikOqr/nEOqx60MlF4
0yO4bK1HAXrqqWN/4UofZWkSqF69XfsVYWqa6EodZmXA99ZUfAXYmPAAAsZy
EArSQ7BpcgC+HbLEroMriamn2vmXkSsency6gZdGpL+nxvAzQcgNsAFqM/4n
WFR3HyDl+nlzUT+TLUJqfj7H8tWfOX6GV1YjEM+7zXyO+A1/dZKTTAWzhieo
5X+GYCuedlBgh8xRTJMJqMPjNSAu+ADAkEeSLNhrO4clWpyf5UUJ354BleWC
PHUs4BX42I4DMkll90Y/s4Ihn4e7ZX/6IhMZ+++9lHoa1C98hjTzJ3BuN5+R
76XPPefIS0B5Sk9V+wnK26wWZPBjqdxcgq295j4rfS/ORwxQQZPgDWQ8DKcO
mUtnrPyA3c2Q5wcKEGBqf7VUMPwy+uSQOB5TQoKP8SuMnAhVEWxtQXMr6mNJ
86eII5iir+9K7B+Z/vrwzZSx7PgSP6oqWgI83JJ7nHDIXaeOaJ/VS4/E+PWx
VknmMFL4cp1erw+zKwC3de3iAgZdikwjRKjzyoBNGMGbC8SiVQcM1LN1ZirU
uvwTxdErVup+Ah9QrvuFrKOnruO3uUbGoiRXy6lmSuW1oOSz+g+rwzcPcjQ5
SVG6M0Z+308o/Y5EEpxEXcyIptazuIF3snNgQLc5OplJv3COD9479ULuVjQi
WsXZ+4G0xoUR9RdhPGZHJqqJBt7lqnQml3M4M/4A/OrVf7gku/QG2qRt9lI6
irg9wUHdyamKqlxKkTwmry1GAdMjEyHVTxFyqHFhGaVRj+q0tlw4NOn59k15
iYMyL6LubP3+5AlrPTBHD4kl0XbWotonStPYJwwYjOXBsXW86aSQK/e/3pjr
FvOYiFYdYkI9HtG9iGaTmfcVesv/kPYl5UlcnvOBERBoyKf4e6WhEAQlLGUQ
Ffrx+7nM+nIlqgEsAysyTSk37B5tAifjVE3EazkYBPkRqp6iK+/+n9fmcnZv
YqA9pVw64ZC65plwEEI3OqboxvKtqrqDIVDurygFn1pkGiqE5F9SAbHlVQ8q
q2kncDD+1uV3OasmZ5UFGVw9SbUFXELR1WB5cyv9ZuGobMs3VoAdefA55ynf
r11Otwjjl1sB22K79LGkNg6na722ZRIf/XBogboCdyhwXOxjnSHlu/J+IH2Y
1U8ZGFhSdNCa1T3+6KtOD6D2UKV45N0r9sD122weaKeSGOUD1qsyNigV3WFk
x0cs3Zydj0pDEW6S8pm8sdd9tbz+V/c2+07BmulZLKY4+xxTy2Fgi5Owwo7L
pQGRfQefVAzSiCkuG9DfxiQIMuHK/I/sVZO5SCLkMdWstjnm3J7G537vq1f4
2syZONOca9SOaD9VC0VO1n6BRrQTxy3cXAYdA3rJgZtqBi2OW71nbadHtkY3
XDZrjeQi6348GeBNNkrtLdnHD+vRE8Aplc2yRE9ITcg2q1mkp/dOVd0xFrcf
jn/02swYqJQt4tYLmNiMgARLvc7rku3lek3HjtkXlz76Z0MA1emXEzWXATKo
rvph9asIS1My3pjR5VvR2dYPMKwawTFjOwP1gigD40eVm7VOKjUOte9VkLzI
ZPu61IOkElRM4Dkm2pr5ike93vAhVubpkKszn6/VxGIK07mi5pm84c+xlya5
wYfLtaCSMu608TVI0O9yDUsnXoNHKBGUTVKjJ7/ABJa0+0/IlqA/jQfdRPee
MZBBfud+w7pKHjYUaFjIUxIxACfaBtVZ6ElDsL0PNAM5sbbA+fpP7TWFKIb9
mS2aWfrVF0HqqVuIjNZrQ2kZOJn7yipDBEHIFQm+Cc8WiXbNCbkkLbUf91+M
WtxVP9RB+PDp8Yqi+oOSczcjw+5R88VkOOtRPE7Uihia2ELiFhAF/CUOm69M
bL03Quwbjbzy6DPH4xVdafXS2LQyzHDVL1n1X4NltDhNu/3WG8PPjLaiCmZc
2uMGO7dTlwPOA2RNIT4S+Ag48LUOjG+OKDcMnOKqrXrWI2GBzRHb7bYDiHda
gcNQpuk1YJ3QS0jVyVm5I8Dml6jtIsaS0KcflxxMMNX7ZoeD9a12sn67l9r3
alDEnPrEi3m4mi0+FwEhHnzQDJKIsVnZfPxW2C5GFIcni/YnGFnnIE3oajtX
QY/vxf7Jr4sUZaHT/+XUFW+pHEluJ0Hle+3sCBQWykWFaQaqu/xnLJgo8aSO
dyp63OlJs55DCFNNQEVoQEslidKV3T2Z1vB4utGKpCIGYijRUDSVU7c7dBhF
mFn6lMkeQUPNvy28O5e1cWNh0q4j44cNQDndhpPyCeiNnzPdHV5Qeet7fT/t
3FV4S7tvMJd8vMa7OU2lWXqw3tQLBGf9Sano6GoFrGML5IEO+Hl8rMiI7HJL
snutvg3a5EgK0/Lqdw7YD1pI76fgoqVm7DZ8DzXOetyBty22NLd+tSlQ2/RF
mSBoPYnhV9C3xUYAhncW0gbby2ok8f2mOPf1DeUsp1dn4w8KUiHnDG6Ls+WI
v9scJjtsoztZ/WGqiFQ7EskJ5hg2rTkP25ckKRa5tLhaqc3F/pjC+iGgqZgp
QKRS9SKkHCXu7iGWclBnGN/B+qS+lljYIHPAwHsfXSPM1ZRoX8t9eFXVtDuv
1fHv8q98ThRXWps14hEHkK1n0mGIaM9VTGfLsmjrWRGtf/XWndUq943CcUye
KSDV/kH9rwknK5JcnLFBWHFRHfIE26Eglxg+86BHJ9Qw9O9aN62vbqPAotob
CbyJq+t5FjOBYz/EfTDDuvR44S+8FjoZ5QpZmXRPkVO92WkEigXoLofmJRb+
gW3Dov980rLKY/3DiGQdNrDskCpUKbiLPt/3ryvJs6rcbINSLvLBxxJBTBYP
9QOJ/olXKrQnoabYv8zI2QM7NpEDzLFcVrWrEAVnyD5xc1ipZjNO88ampBXY
j96DyUNBJOokBSufGIvBWdJYdLaBQlfex4VAj1TFP/HAmKjbtTRcGalrGV+a
bT/sUYTIW59Z0a2orG21D94RVN2JxVG03YmX7CpPNnhfmj49lD5/0hNfOT97
+dKIggEPNezsbOpWRAuzUOUef5WLyIv33LG81tVB3FSVeiXTEj1IAeVQAHcA
TOQnDSPpWe5BFytK0QdNE7taqj+Fuh44jItL22/VITPE3Aj7ccVJu8ool6r9
nIxYEf/Q9CpBFGjfyPilFltPGiISy2+YXa1eclrvpMzGUGVslOkzRgR857WH
QsdBNv14UpTkikbGjT+2hqz+h/b6alaFcECOl/szKx1Zv9ZkZPfsBNlmzLsx
pyFzoMzP0+WI9gTHYBDBBuEPquY+js0G6x7Xxi3tW3bA9OSOVuBAGZ1fba05
ACgPvtFz/LV5ujGwpgGfukASUe2lK6jhN87hX0AlfTSlMyBm+Hpu1x3zckK9
KtaEwFzJ4ePP2OYWU/AiAaJBgFslOLexSaGoowxr4Xx4JvaYxZVZI19nwtwo
InSO5bqbxkkdNDDs+CEG7dvVLcMnFHAMptyqVJX27ZO+QBkrICsWWgPT1v+M
Q3+JMaRYzJ/OKsAstaAuuATNsXKrP42FCamafHuxUfzgMIXB4js9R2QbpTTm
PsiqVIBwZibDQBYJK56SS2gmW+esQOvjuvmCxbxoLhMQXXnXAi5sg7PADVEj
T9QJBe44cryshp8kiI8tJm/Ja4Kl1KMxs3WLQWUy1qe4TtJx+uHJuYcr9vz7
xXVfLUFImAcdKZ0dhwE9Yht8+gflQ2ilHIKGYdR6MKkA0rxjD0kizNGulA9c
q/1Bi1p2Sm8m9RGGFfkIFO/RUuvmCDcFxC6iHGF5LcBp5jLP7kUWvns1ZEhR
Uj4iVivS3tiV3DOJb+cR+oKxeoutIXGQ6GSpm5aVzC94F/WVK2Mg+xVxJ+di
87w2GtKMCxBNE8oVxT0jqMnyU6FQoU08e08CJkoTbKbuJca8QF2MwlgLghvj
7uMz8eiZA20/fdnXBRLqCGtobZlgjjsNjpdND0U64mF+SjnzfB9HU/Cd0sZA
ZiHj692Fi5JUDeGNOg5nFttJVqsJn2PAUQdXR4YfzDYTnqZF+JPydnMZ6dRe
JKFXll31fqvrl79oZtfsOUse4woBw/7AEm/SRGGb85OuwDXSr8ZpPJsUFjvB
Pkol52gg4W53lVdqHU36kYHCS+Vo3Q9L9M2gUzwVmvY9871mMhuXk3KOI1OG
5wKroVC/7MnlnOla9KOcsAlyU1ob6NhPBpEC9C6gzOP3ubY8485Zlz1KbsOL
3M5JBquxX/cJXdkRo+Sv8RsRPA9O4W1MfWlj1GkaXhvj/v6bMnl2vzIHXEF+
OdxCcghKGyVBUP+zKXz8CB0fwostkv9j/QU2uSx9V9vCpl0ETNUjH6B3kWxE
7tYro9IgWBbU33SSa7XHcgwQodbSwMU5TFanyqJINlo+GPfzUm71drRhcWx1
LU+KqT8XFWp+nA6d2dY3SaqS4iSVBpZkDnUPqglvAeBeXonMucLRWqPqMybB
VJClyTfLtxbAnkIf63NFlYaxqDFne57TfTfYBrOTW6qqj3p0KHoyU2pKQ5qK
ipZxo/KirKyqomf9XHu9xFlTzEnV7VLdHBfbaiF9tly+fahXdHGHIyYxanVw
XtAGziOM4gVB0v0Kzcb2xLAgKbrV6BDfy5Sovyp8jWuhEpW7d0lCxQn1mAoY
ZQPEQHHHuRQQjcllGddgloLv4e8PnDy8DZo4/aOKM3BhmA+y0fADstgCq1Kc
NU1QPTeCJso4CQipFz5mHOah3+5UrbTCsera8wFYCHpdSAUmOXo4rwr9Ql+H
FEp0A6WfBeFuVYklFDG9I1LYAklHk+dmNqus3WzJpxRK2NcyL0ZrRQefMwIT
OMSFLuMPiD3o8lrwx9KKBxMOy3cIQv8cfL5gxFoFwlxdCY6xkK7xilMjNx1z
Su+MYKpkl119yU2XQIghx8Rc6HYb7apHO1qsn9P4bpRoyzmSm0myt/d6rsQZ
Y0yWUVOjHzZtoB88XoMAUa6wtTwAWBtNgPdpiEppmVgm/klNDsFHbGoiugkJ
cYRf3sR4z8Rj43cULmHqqVImlRxp64fB8ZlhCYAK0rXhPssKTjH8BxbXTzLi
nl2Py1YCzBe0zESI+QsBsCAfinjllhLeHMyMwUBaliE+FiDli5Pn24WJlVds
B+fR+OANdeadjfOA006EFhx2b6xTcOB8CMnZXiOMwm7v0xxGOEiFd1QBRlDj
bGsKBc/qwidgX5ZKGlAi24NiYf/niCpzZLlpo4ARS1TEtZa+RChidizMNb74
XItDenMg1AGQpvbrPgJ4jjwLz3AhZqUPEhAWecvzISyF4a+7laL8EI1bk+6p
gEpg9tTKMj9GvIpjNFAhqCfEHqHtCpURYHtPZzBI42K0Qg+deqj+3TmtuB6Y
REKCfSsHz0MIDi0eHk0y1yjGre/26q3TshjffB4NSrTl3+14y6DFyzqsPt2y
Fx3N+eP+JW3nSlnGIqqQSHzvh0+Br9U8zT52IIHXOzlaZbAfBxkyu/kg6wBy
3mwe5pxIPkxkLexTXKE1CkBkUk0ctooDTUUYTvJEYdqa8PfVlg/9+nuuYeKb
B1s1JoCjgHIxYJdtkZju/zljpU98PjcAQn6mMqIYPCRfPs+/GFxwgFhN/5yW
CsXjLU1Q+xVsDySF/SytYhPnJ99AxpUh/qYP+sESPDjHc8OVl/RyoAsaK3de
/A6cpUj9msPT7grC2cXJdtP4CEODPkcIcs8X/jW4HLKZvf7cFhGIrH8CKP+D
aJju0Q4uew6CjOrymc0KYuxtFDYcqORt1n1cC3Mf7e7P8oePXQbwBEJ/5FGO
4wmzOD4UsEoQ4g+J1sdmiZJQOIxdLzno5L5l66hGbEfM9Kaafdz5ngeqITgA
D84CwmVotQIcTixRceO3QJGI6M4bqJCgh00ObUc5ffyKlLRoHUXe+NtvO1vT
PzgK5MmPHMsRqKVt5Caht8Q8z6+TcFoqaggsltccZm15Ayqf6MoCU1cjTSX2
8ply29mL60nfiTwNCR9BYJdyn7U4xP9xoIp1bfmRx5GNnrN60U4/y1IqDBXU
E/RrtnJaBYznw3EEBwwsCufOAoze6fZ+u+4ylGhZPAkvAEUVUxF1Ffb1GCSr
rdgV6YnJ0Pt4HJxfPe6iDgayfm7Yk0cReKoKLT5pOfNE9dbMzjt547Ve99iC
6SN4V+LZDFxc5JFR4vvSAadwWkIhFvoqjbRvCdSykLpMC4+dxsaozdudRdPX
303HhCn7+rkW03R7eQ/yINLTRhKpOFWIMR/YGruzbCvA8OM5HVrxSfL5cXkn
9lwQ27nDZAxFjTeCD7eMa9bLd5CEFt2SAAIqNSIL1dyiWpFqRdxwFQQPI6rK
u3RFDAx0K4vy1VqRJYfNjOXamSizDBb+x4tBur1Icym1A2eLE2EBts4XeWHP
c50yRnVvtpMbX0JvLjoamE+s890ZChzaHjTrP9K60XWEZLLzMr2gU1LKW+PJ
ldiX/uMC9CzhGIEqbDCU6klQhg2xenijxLEPWNzyRAzRCSmxyJecSYccYhf4
jIQQdqsK+qaH87wzMhkmcQw3naO+uZsqYqGoawL88Phjy0aiAzCe1erLbEgM
5N5X57eesK9CFQDB6DWws2nwPJAJZcc6RGWlnLcB9c4yWqPYek8g6lemRDaO
LBU8UTIPIYIanGugdnPlycwqLBbS07yvQuc9KCP8uJxAakinTJWqnJ0M02F+
T6o3PyZa4g3pCu6qwIfq7WAXiRK++C0ae2qwJvKdO7WYJ7P9rrr7doW/AGMa
smp0/k/hNerxJnSnbXMChD5RVcE64YYNKInPWJh4lIDOr9DoDhIAbRI6i/+V
pF21NsOzl+uvOF/3CPZxVeUXxmJWPrkspmSiZgOVXwdrJL/Hfn5e4flAzKj+
mq8hTCTNRyOIZNUOFdN47a/PEMkC9BJSxf+YXqlmTmsCobE3ESYQw4n65eCe
CdNrvQ6J9sk3KZea4XjY1CXaIruyJYMnaVzW69cVbF7T0Z2IxSD0ZehuThFS
a5wba+FWVbxHC4HLK+cAZOEl/VbPA2OeiCeGu3dfif2u50h6eT7YNBFx3LBF
dVr8ZmvjBK7B11FobL13jW2nK80um+5AV/A+BeZSJjM2dBCanQ6RK/uvEjoU
4PBuhH9i2anM7gxltwdTwiExWJTKxL4IX2YB+371bhMBUNSLu+Ah5Qzfk4ll
4jjSwAAZPtKFI7moSlFPzHtSpxK+q7SfJD6sxykPX9gUDZwW/d+fyrN1tWeM
PhbCqaC48QKe6qDDGZfhxl4s0NZPPKghGac/K+osqgrFYkFIJ8/Wu5KGnfaS
eXleboUnrresKykaahYl2ZeyyPy8dwtWplekKzDaok4CtHzjmZ0m6Rtt5Zoo
8536ge+6120brJ7eebWn8ZnIIcJkI51r+RPVrKOLpZA+kZbqeIedZep8JlFq
r6z8WmqPIj5yKxSX7m+5BMLZaJooW6ep9GUFkojmeHVQTZEZ8BRrNd8Le3zZ
vKTFg8RJ44AuIjxujvE46uFi3gSyXVxpRyoHwcDHUa4DwVjUe0mmSPetON6h
MrVHw8pc4GauBRf0rY8oqh+mzYpYXGg3tmM3xZKomSitNMD/r1xYDWtArmcl
EARRBCfHeCtq28IQn3I0ez1zclGvvclwtlUNH3hjQGaZld9xFsg0OEMTJdsp
jgAovw8wJUCiZTXnbgrmAtfy796dJ/Pmq1PYzMByQ7YwmuNG+4YWQ9PXleWh
Kpkas3Y7dfuRJ9bSfoORqTKbZJt/ZAsCmaTmF8qRMSvEXl5MjbuxHZaz5D1M
OKT/mlXbyQdyMO9f8eGOADcVXjxvdlL0RLAod7nBPienYkEIyU0qQ1wszoYz
Xen5jfh7kPHgodksntTzbg9U654Ofyi8obcs/DyAF7yJkaY5u/z6aAD3jDlS
9x8WuxdeIQVZUJlMVn6NdzQ3ot644XMjedbDiewLJcsvZloWSVFCgRkQSYiY
aJBXK8Tf2ifnpWgpEkNauCTg0nViXXFoVIDenEeRfDtrB6md2kyYRn++Jjz0
zMzZW9JCumv7+OExN5pnOeXzx3mI0++QU8T/CB4P/MLDsWprt8iX22fys6E0
rGeGwpW3I+1DH1QhqU1nzCJ6YfaaA46QYVK5P0frvJxziXHY4uW3ysVB1CF1
fO5nFNfe0gH+Rp3h2dIHeQ2aWEEoqvDoN/3D8G1gNn1lY8+/XNCTdstYt5kv
FH6sAt9YtEtLwX7P+JbuOA0X1UEarbhnGu7O9daSPoJNliEiF8tFGVwGDI6+
/Q1StsGAIP3AVPNKRKVCVwrDXiVRR0XMvifLWDxG75GfFGbUHvDuf+95oP/f
hQCsa1q8g/edn/6mSbCmMMnqOz8rbSYVhPeRvwSzCSoq0fgHqIIxqXUMhR6o
IrG0m0KyttmYAsKeon3GaIL1cQp6yvt7Pxlq3LbY25Z2wIWOE+ifnRTaSbCf
sATBFrcUR7WCpC+srcSlsguk4cKjw3lHhkMBHMlNGTihIXo9UB/8VCgESlmQ
EASUEBAAfBOlOijNflv0WggNPDz3tAZq4GzuCAf08kpemiU+zGt+7az7+uVi
SrEAMRFy21rL1cmSQSQ5GJM3rj1ZHWb3D9kYG/xVNaV566Bb/0GR7il1Gw3w
+hPTwMOQ/+howOiatIo2TvhUFcNqH16O0dbdFo8Tx+8TqeKjpWboW8IDfZI6
6gQ0zarxyhGa6l2RE8b1dLjwQ0hFUX1UROEsGtr8vEyfLvJfsnqqVFfFwbgA
RDmBl+RBjtocBNlXl3iFXJCs6tku2OBtfqjTguyb47h8pi48yoiROt10dbzA
g5BbnKNCWvnhJdoGY212+9ZdLetLSH45CjtrMMNdVUy5WPmPL+LKJwLoynlR
4soy/vLIcw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGMi+1ymUkmEvtcAHW1IGc8AQEP1RUC4GziqYUPN6W36KEKnv033AkpNWjd9L4ePyDmd46NyPyaV+3Ybsoe8r8TdMZs90Udnne9/Tn0Js1HqpDC02+MC/ANgqIEryjTufBdWSrbCbvRsl7PoWc+U9XNm4W6fEUDeamVgGKQOYkXoMX1RTLiijUapE1LopFxAD/VgdWbF1TzGYlHwdPLNTvg/RNbXq0Ac3DYJRCd0BgLQFHobLtn3+x4WftaJY9v8mzdY8tAQJ35upi9PY5XapnhSRBeP6ginwsgg+m2IWW/t/0ZR7fMaqHv+czjAWPUIgS2GiPla+dCUL1c/6dkZsYKVDbW0bFZ5xHzFvPOy4A8FqunnNegB9cCHKIGDlD6GZLkMxDKUUU7b1Yj5+kS/8xHelLwgQBMyDQnvFg5ddudIS0zDKHcDtpySHLyr+rdFgqa13boiIlZFr+x0sfB52NvBDaBYNWK+uQDdla5Jf7TC7/hGSSOda6G0vWx5NyKvzohbWl8mRp1ED2VRa2Y/P8u1ZjXiWwqdnkt/86p6JNCFqJL5kpOuJFiXD3aNWfs8rgOg2+mUDkk7xG6+Z5HKxOfoec9mzMcAl9AV5sGVIcwcB7/HW7MeTB/M7A6weuAdSGH0pOE98Kb3ogolAAN5e81cF1n4DmN4Cluu4n9TzBZf+Jgg6sDljj0lCzDCIImXmKt1HPrO4rRJkox3DghPwY8hBioSc035R5nUqP+/NVNB3LJs9PQdgiAKBqdkVtW4RlnDTtur7x6s0dSxJGsT2mtF"
`endif