// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
w+B+hh00hONqQgRd7g4XLTdUxStMUErQa3qh73OMWVkLpdKf4Lzdm/cTRo3m
ZAQKLRqFPCxYM8etIpPMl5sYDBkujZmyvF01IshxPNSQ4wLCJhKuvLyMaE0I
goa/juRyohKRebdHXsvZnRZmjtrMkjHpZKnBDTF+1UfDsb1WCzyroBVfVbx7
ZlcjG/+vbkeNbV/QT+IhjGlHqZ/264WqbJj8JpX3aXDFNWVNjwGoHAAU3bae
ImYUWjiAvWXaVquVsyWgaVnn2Rhn239cGGdYeTnPk1pLWWo0e+Hy8X+GJw5n
yo56vwXpwCkXj0bh8+c7OchnhQj1LwdARWbwIDiWbQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h3ycpADLByfW/M5ipTK4OIRf+cbntXssx/laWhYedMxmsR5I5M/3/MCgvgGG
vFLpkpSLW6P0p9eh31apTjFCGGbRhlqKY/ORxDbzGeeOeazumE7LlHKaTN5z
Tysyrs+ZodDmMCh8jIXHvv/Fu8VY0CDqgsZGRLcIcXC62u19SA2x0Ejov9fw
AdZsG+d4KPv0sAiDe29NuXglCXwcaSXPpMBLrdfefYugW8hge2YMXl0u4y3b
Tq7p5GsWKIS+Yu0w/Yjdh5Esu71dw3XEQTfwAtrEQh2/ID2/tBE5kxZuIldE
FCmGDZUuNhVodAA3mm3qGiZwWymejZj/AMkn2hvaPA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R6Ox/o30Y9AfR89/2j9iFQbZU/lRT8SfNaKw27JMn27VMFfrgHkgG9FR3BLo
LxB2YI3jrRbWHAyxpCWxlK4kD34nlwLMT1kntRRAFe1mmTZDRPHRFYd2BMsk
S1OegV55UeiyK7AdYG1FV/GQCDM9fJvk0tgVOU97hDb0B5XkaWpYJIfot6KC
Qysb+UPMC54Wvjh9cSURKNOpfWVkwFWUk1npQZFvAtifad+tv1grv12mJBpe
k64BJQpPJII5pvR5PYp6yoEjgBIpoGoP3opIzJmErMAoXXLK0V0uG+Ms798O
1akAQzNl1sH6VBPkhvLGuot9kjeIh1Q1RA07mWw+zA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cF2o4au+rDze0TxlM8+5GXsnFxJCcPAOtWOXRIB9c8caJI3W66u1B+AR5+uw
gpf7Pr1AMqpOr6G4mhMeNp9ed9LQ1fTVwX3e1NoGfxomRoWo/ZaEnAYg/6z0
lcEc7tajIywE/YEQ1z2Rs2BZQDwEjJ4duD3BYbF/SjD68dYOOhDvWU+NAF9d
y7NaLUPac7yIOURbv38h/AsVohK9J/oc8o0Vngus+UzG5q8QiBRsSM5Cj7jM
hREi6KNupHivDEhCdu4ZYTJ+x+97xUiN2Oqmdr+5v5QEU8wvgBGrVM7dZUfJ
f0AaQoi/MuS2EBgQIWmUpX1CuCjFG661DP4ZHlq4uA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GLI53xIQULz8QmaQ+tXgtaAydCq5QDB+NhuVUhIB7sZmvaJ1qhHZ0F8nm8mq
c5oT8qQfMaVmVgk9XY53zGOoz87+eWrFdek/d3JELow+/6k3/2/aSpR4ubvz
DGSHD9QfFCFtNm9cYHGE/+pdbh21z+hOtqs7OTqSuSr8BkzltpM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pbN1Kpea5DyqgXifB11WsVe/L6/oSWQK4Yvl4gl7WKO9BDBy2AGUzGDIAvSu
bgNi1rhPA3/owkbkijl6bTsNlkqPA/NaPqXtccuuno4GSUsXLckA4MxY3ALw
dx/xClqnNEd2E81efadDxKUqjF1H0Wct/kleIIImFoRV/9jd4CIWgoUKrhMS
DjkdfLFOpC/NHxhRJj4lFKFmJbu2G5+JTqqrswCc1PgcJ9CeinibDWB80qL8
0M5rZdahNCwkBsSokXOEQ2TDWROtj3Kd9vyyzGZ7QRITsg0hZrq/1kMMKqfC
JSZIZ5kWfqh5do1OEFiV/s+vOHlyoNypd9PjFUcAuYyU3IPYNanUvAit6TPy
g7cHy2dqFOyKivdul75HtnFvd2DWutw/iq6V7N6KRuWm2utUluAtxgpm/Ws/
aIdsT9sOsSVv+b6daz+1ronJoD0D1TMDU7/URx3xVKM73QXvTr/roDsGTtic
sMk4hFPOsqtaqbWpAZFZ6N1xcnBUufSz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gR74/GM1BK43z2IlNSH3LnoJ1AUlNYgf1Cxho0E//66NJoF6U76IOodpbxSR
JjswX+Y3MfCX7Xs/eatM6gKGhjYhn1zcKGWgYMN8qGg2RQzRbxw1DBc7MTqp
rrRxE+qlv/Z2a7DlZeNflROjeQUGCoJlntrRKYK6MQCt9xeFbBM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XQJt+NESVmL2ddrj5FwuWKnCPjGrPW+kN/GB/nvVZaC/IEV/hpVD/4MBsoVt
C07V5D+uO6YnoW4Yu2ioNMlWElTgFGYE9x6TgsjlfACzSE3r8aR4mFAA/hrC
ZxvJLo6615HWPGzxpSEhbaxsBEacXb6sUzIUuDhw/hTBjPqAJ3w=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1168)
`pragma protect data_block
u40Z0aUBL0q3tSmDuG7o6ruYWH8MfyPZDA7DlI1kin0FsThJOvxupQtMLfpr
BAtIFxU7Uhp78Z+Ig8QqCZu2mm5g8NpHclnjRN0zoP663xhgPbot0Cj+m/m1
i4lN+/Fz7R8iCr9wqBBHWqzozZg+/EjNxnU4VFKL3xYS3XXh7XponAMPNtCL
ig2mmKM0aKN5RiKnbxOMI58ElYEFXRNV2i7QVTd5ay0hVikBOpPFnMLUNAtZ
7qyJaujsWdLBQndFWI/04m1A5mIm2jSOgSIJLkvKhvcdBMBx4Tp5Pkg7EP/g
4vHL4WR8amalUMkg0TV+TBL4gWQbwvR5+QEASrAX079Lc9BCWCCoCFUtfTYo
ExqFc15lFV9HZQXPjuB5PhEHpMlz4dquROE40cy5DEPh1lTsPX24hjL3JIoa
vDcp2GfzCT0HlcE+x7B+Mubk02yss4jXtOsDdSRFrjbnTcBNiuv1baEoYTlR
6sXIX7Nm4Dt/p91v4KLSSEgHQ++rLm5oHWfPd4PT6LC+c5gRpuo4+sIdJ3gQ
CVPIfVowFq5jnU7hq1ZNYEnL8hKLQDUpkPY+dsUMb4bnISedpSTqaL8ZiBgG
NoFu06lrd+O+D7NBER37ia3OJjFpYr6/3+MX2Hz5DTZ5ufal11H2JWD/oMlY
cR0zAfONIPCGkKRd96G7qx+vREvA3JnjJ5949WYlBiQAAPJCHdqGMHTE1id5
EwLqQiHuWSAldYa0HJhh7HA6uL9FcOHru2RJq2UhhM12nKj6b5cVR1ocao3v
/U5CLX6vjrO3sUsCOKEzVPwBtmeZ/1jwAxo6Y2uYEylXNynBghC3rwhmREn8
sHiBuqDNRVCQIkIk0aqNhYq/1I63iVAC0xFBKJtXtCdAQhIjclesLT+DZp6y
ec4o3jAnZkBMsgTGsohtiho1UFvCwLK4CeUZRFVGO+UI7XktyLLhBMPwcsxr
xSiTVXim2AYX6YppOSoPAzVGPJISUMjDUZldJ/g4lHhhctNupZJMQ2Vb28dR
CQTG6C8sqVSaUtyrgyZmyBtwkVqzqeIy/QeDjiAwSNFiP08ekYvqYSp2p9bp
KhN64bXLWDnPnI+GAvvzyBsQ0LRfQdIhEO7trhnR7p4hh2DueRaeJ+z/bVzM
q6mxsESGSbFEOUJrS0QceFkLgCctZ/Z+R1u/IorXtJG1WacugJHi2X33ELPo
DHcJ+Wp5oOnqi1faoPjYw8jjEHRMI59EDyEh+Ns7gaWUqvg32Pi6h/4JWRCw
v4dM5/qjcVgUbFfmUHDRLdZ0MzfnPdh/tVLzq7Xhu0v7S0kfYcwso0+gCMp/
iwUIF1nPDVKclsmAy6R3r9Fk9djELl8T2pn+cg71HhLsijuAFPb0k5kdd5mJ
HdhaZGC4xBb2JvP0m9t/sQZFjEMXDZbNSA2LfGYP4ZWdo/WntYSk+95ZT+0T
IeQFdhZVQZTTN5YKyo/CwZNIguZ8Ko0R3KUMOerSP6ftlIRNu7IZTnY59Nhu
GZecWwAB0lJc9orCpyRILbMRQwuq3HPQQwwq0MYX2DJpMftFF9XbB/kHpw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wjsI3zW5X5ssxMVizgZj2axQaDxcoMgwcweLAku6z00aOsyPrjqz0Lmk+RbX36yl0vfUebAW/Wz0KP8nV8CYn/WEuw+yZ5ktwwOzpAUG4XX2+a2BWBwUt1k/rtRSEEwbm6Fz7lZsmFAYqBs0uzwJ1lzgK+KGdrVUEFp2rrM0clUAZJPMWUTOlqH559YrANiUeWnsBXQnWNOTgg+nw50SiPVfxgB1NWk43v3jv8HXV7FksFEN7/LwRdvb00HZbSKAmDiXbbUlwklnAYJ1LBF5EBTm4R+tImnwFVIn8OrQyU6lUtxkhX1LoP6gcfBYbjXPunLl3pAYNbl6/hwTs3LXXzkQu/q4Nq+xZWil5NpvQf17duRcTg68HwUncCOENpW5GVsX2WkaVMjMnSnMGhLtDgnsThSYF/JcuENxzei1DlfgDY8pysKqrz7Kc6McMzX83Gw/KRUlanlGNziLBDSpzcmwEuE+hQqTw2hlY5aAKoo+p3GHTqWg7dKpd5y3DqhR2zJtof1S0kOUvYxGWHPG62OwTQRR8B+PVEQfqczgkcAnDpJBoy5b801FKkqsB5s4s3cbtz8QfsL5OwcjRMMO2dOVhC1gcMhXyP3piwDWWWrP8XXLz4ieYjIzrzv1ofZNKtNia9t/sgziHixCxzVOlmAIqjgkGeHKCK444aeUqUj6w10gsQbYa2pRCTAft8jXpMfSPs4+2ySgg+YyMUGkxzzGwAgyJ7uoR0Y6oX0fJzzT2uJ90FgvCEvqlhzy1kMOhPHCxLQVHOlVGpSHnIhWC+X"
`endif