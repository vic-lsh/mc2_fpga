// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cxAnV1m93PlvScocJl7sj+9bRZSAr5AiFNMus4WZ0PLWMHSAWqPrdQL90SPv
kAsuLx/rBZtfyjyS4G6GyjyiA5Ipv6sPFud0qsdeAc3or69TzepcRcu1yjaU
AltVYk88lr1ZQzIAm59IP3tvj9qNzVXQjw0g8GQClDopAQ/N67/y0wKKv7YM
D2UoTog04Fz2Kz9uriJbRSgdqHKcvPT+95QotxplmS182GOy/+i9E6L3jgon
mNOlbyosdeo55jT6xGCpP4XY5FStJAVTN/Guq4HXJ+OUjdcLqjI81YpdI0fY
qKA597+PXW+wO76R78spHHcw+4QpdXyZ9zozWIoFMQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B7haXwkJXFUuJYYakEQcJPaar6JQpgrx6tLBCFE06gE04ZtAEgTNlxr8rWHz
k7TNPvEB9DwCCUk08DilsWICQdHMP9A0//bb4YFISYDJqYy6qLvO6MgzDkx1
MTwekuMBc7qXDeS3QTQMlHx9/lGRZZviHKhXE9u+fLKBlGfgdLqZtfiJ0Re3
mrf662ls+ie3DqVxqevR7/MybAHwErSMklRDcK9UhBaGcc9RETchL/VhWdSR
tJU+Jbc8nEYe7F2n5ZMShx3FvDg/NUPpTNl0unAF42cvNsryzjfx2ui/tiix
Lxp5r/+x1bgcg5CsKQtgNGzyEmw92o1fmnvpvVSolw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XzpL8CHKd8FoxdmvBazy5n9xA4N/G8DUNmB4VxOjhF5l8PAivW7AAX1Aclpm
rgOZwlfYGtodRWpnCq770Fsl6E0E4m40Tzt/N1pCz+ONezrEIoH7U6fSHSt+
EGQUvWjtaajbo8p0SFBh5fXeKTuien+B5qHNE2kUlSKtAXkbj71Bk101Daas
ECZeaQxVQLz4CQvboGxbqcRfXieJ/JCEeRenZ4PqB57AIPAu1U9y99d9CYfA
/GSfe94/XkttfaTY6Kmm59Xefl3w0epouTWLZVgk/l2KkqbnR3V8/J8FS3cp
n/nNPCHFru1B/WeEBZ7Ed6iMddI1pWCNUf8dl7PZgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jbDbIN4dLGg/qg600wvvgs278hc7M4x/Opi/YHYhZe73nccpMm2siGzK/EsR
TJcH8ET5d2WM0JDu+XzYkFMOtNn2YzKDg7VSZmqc7edJXtxtSAEi0gvi3Rf1
S+5vxg0V8PDzULQ+L2XZwC9ODuZvmxJXAVSkvYVruT+8XGhADZ/pcPVIlVxz
ktSZ2S8TFT2/NEvfG/mAXVkNZKYZPh4Ym7xHfIPn1i7uOzTMsoNxe82Uz13S
/yULHIsRZ+i9Mf+ajREfjlqusTesRIhBE/uaWy1raXvNZfURMD0aYA+GdKtj
ceYyR1YzC2bIgovdo7uggGw9JiGEkYJadYRh7bDrXg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k/1hzj8q0HTSvfRlIs2aCVtBgo47wkwWnwOQalIbrjibiQZ5lwQDgRcLupdd
ePF3dJ/cCeBBky0t7DhFGe/g5s+F/+v4Coz+glSHFdPgOgeo+B8roymtZoAm
RDcFqJrwFbWvB5Aubei/h82bxiTrWG93KHzXCydfOlm7ApokHJc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LvoU5v5X6Ov+zNDFUvbVV4kJn9UQP0KKaAm3xYNQ21sQFZFQZACVBBpPLbi6
LVhBkzhjCe00atg9soQdnM4Zo5+Fo3ovoXaNgAyD0c/WhgaXp2/JHaWw1TEv
LHspc+8P5JhdAY76xO/qiHTTzzs4fh4Zj7LQO6hS1ryWLWiA/nibAT/I0aQa
3BFE6ad9Hxzt9gMmGbfA/32Wn+xX0N4me97jXafaeDJqPV9izprkAfWI4Ih6
19oQiBXRVGVMFvVL9QzuG52N61/KBXZlllBTrGXTeA+97jdbGHeKBeuLu71e
SMbJobQuuQ0sF4kXrrhGdtVecU+efs9fpLcnkrFM0yTNiN2Yj56BEyy6rk/+
HINOteXkgYWgCVgGUvUAK7bGAoiqMmXhLQyeY+k3/A+hD6a8y4OVnwDKpDz1
P2hRkBLzXS5jWUGWis2e5GSYzEHdZ1E2JYTg7fUYE1szFK3Tp8xQg008CasC
Ls1dqpl09sn/3wVgex/vfOr0jM9tShYx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mDwFXWtzmAw67NkBcRfwc+rfnqWKjnUh88EPwTcGcHSDWa2iLROs7shnYmjt
uvgqXk9iQXnOxm/RTQyeIPT6YfJd/fIA7Pf+1BB58j42qvSJIJcZhbIQzpgL
VK0TYw66BW+jN/fbQ6q2GITP8HTKRVukZTkWf5CuxG1v3GCs7CM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A4PKzooPQi3G6ccIZm+yNMqRCz0Rbo+UgYVae/G1fZqQzc/PWeRxbPuiY3Q0
wOFndNZ6uidYOfLbLeA7zCH+zYJXRc9glnA2DXuY0rpSmQrA5z8g5j2EVLXS
rDvRB/Vj+AMWW1fteG02NsHrJ7GTouFwfFSZ03Yuwwqs/EtJFic=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3232)
`pragma protect data_block
1GOeA/bgX+LZoGPIRC2KvRbMcsEmFB2VOYaZ7AhlzWuSjXf1qAVWjkKDVmWG
RtG80kOqdFOmbqVt2VCnCePqrndqsbhY5GDAxJgUQ5JaYbR4bDnZRGHbWqde
09pycqyDmVyI8iIjrmRCWbyv3zOkgTGuR9p7/6woDUPwZoBb1+BAK31xafF2
XzcbpV0shmBF0GmjyfwrM5/f3fmWxS2fma0V9Oz2PNy3tS4d9fCyNpeZj75a
1W24dGO2rCCMYKaTjOO9kXr7N4aJJ+X7OzUKryxG4+ann9hgx9frgcSSwYjM
tUU3dW3IYcPXBn0gVFMQ+ONS3vK4XXCbTgyGPQqFI27vNxjVMWW0O/cOJJKW
6mTR1iTJzGX/M2AwRBf0MsrRVINQ6bLJKbCy2WvoxuJ3n6e2bfCnjWw+33Hk
bYuUCW/Vnc+wZp64YUH+0yZtIGAwwm7YAvO6XVS7nZDppDNe3CivQabdUrcX
nCFIwXLEcjycu8l4UZYzi+KCx5XFMBUU94fbwlFPzj96PTMnY+rKkOrmU0Ih
M5BPpk8aQammDIBeXt7eROcnL9zMejcygahSKbedRXsKI1H3AxdJPOEZ7QWC
9ToY6ctbCaEtImnfyKJamn8HuKBEYca3LlK3AjCY90hVA/kc77XmFzghdKag
0o9ReG6JgaijTqyjTjBEUSS7Q3kcg2l/r+mh/rGwTDnohXQgdfhQRR/NbwxG
a7+7dJgcutsI6j4s5AFH9qze/wA3lQx9PeuSb4oNYDTi6R+khB3URYrSsbsO
wBBdTOM/KOeAzWWpaefGLOaYu4QAk3GoFlIdhZfMAuYUlZoUgWbI3u04q5Yj
/46ibiaxpbOf5OIQRizxpOqkO/MqME4Vs57Uystb71+0jq+mQxy6Kq5uq/7C
tWDI++7MzAx2KiBT2Ecx3NfB2sNQnZA+2ukPifGjtWAmAqEJmOfGUHXWsv17
eYgq0mgc205ciMzKSuAv3bggyt/A5gB1F7lbfbLNxySc9bdjSU41sPrSXmnP
OJED9lbHoOg8yOE4GQtyO/lfhLE+v2anV1i2ut15PMqsr6sYZSjaai6ihMyN
rstabpKLyu2noICT1uFQhjFe1YCkhcFr8Hs9kM2aLyB5+AJIz/p7R/DtxfE4
/OmPPQSEtsi+xn6NpST5Qp93ohB0vw5AuRvBmOSc7LfuVWXtudMBi/9kPlFJ
2nVzJn/CqK43IA6XekCsJxJV8v2EvNGmUmiMD471Xc5qJhmrqgD0uRwNKtyQ
Doa0+VzBV25DJhA3D84NLamviVPV3GQDiLsBZrx3jRkNtSgr6LkgzDIcOb9V
Fv2TzGALmWrPUxxF7JcreqfRKX72jQvKwCJ5HWBd1dQqbtGFaTV0qIaBjDcn
hE5mH5PFgawOKE3xDg4dWwR6m0SukFnIULCcK8uVyIjbqzGZIzeVjr05+IHt
dVU7Vf2mZO6WrqSmw42SDbw95qTjM1WHefVU4dLgNPAOIl/ixbaMSSbGh/bR
IEEJG9lhNg5MXf5iAgghB58qp9wLRtImylaWVSOe01EU3DqrxwljIEqSlL1s
5XM8C1323d0AiJZgRNHGpiGTvz2ouzb57JutOIai7Lw2P0ZclN/mZyRZcfBO
EQJHU2l9XyyZcZbA64+cTbyUmdp5J72Mxx5HLiFA4+zT7TuclsKW+vMbrhMH
loOUqX2HXcq6O+pLweCCclwi3XxEONN7KhCR6SnIRV5SSqj5Db0YGXlSvwjd
5ftDF/Ag8gUwTL1cmpHYhLsUkQ6beP2XuVq17IWM3e7k5VIPNhgQgCVitBz5
nuKaQb9qEkroZwqGBPqtEilR/n9xmXWpD+/P7mBx8jhOolkOlzfDPdbqV2Ci
6se2AsAs1vIZufXfTcTDAl4rgzS1CGCCSqnn5C+GoIlaVM9gB6eGCluBTx7F
kF1aqRYosH4q0KRsZF4shd5GruDnX9ZXR2Np0npnpAj+sM69uvLVuvoHBcEG
qNp0oNDi1OvnADao77YEj/zDOHTHlEwl1qxWHyAIBIY+9MUOyzoKHumJKG62
zaqYNeJq9xWCh2H20qrnRV9o5Z6j7gHGnFuuXdAhbHES0rUqsgc1u8fAcIRX
ZjR5uynn8O5RSJXJZhmoWdm23rcoOS37N0KN9C34hwjPahF80Mr33LTMWSKd
OI8iRB3eVXDNKg9C8V5MG1NjX/1msn7ZWk1tCNOhh1d8te730SzXMbnti+Lh
2QGfrMxbcMeEKcAut7Sei1bNS6ov03gafPxjstWZ8UQAJGiQEJm+5AE0ubqo
UJY0q8YyubDTuBSoQy4LML5+QVjKkPucOwSIBNI3srhg7pLPJEpDBoB6axGH
ukqoQqrcWgP/1td5S8f5Yw03aqx3GWC8oHNBJDyK7ovcLXFU1vMir4r6Vjer
N2eQ8bwT6UQoRV8UKsqZ8qlb+GL+h83r3AToq7ZgxtQYJuGhcCSrTXUmpRZd
VivWDhNbkxK4ExlBl87P4A0Up++yszUkDBk5sxGPdm+tYoGYlaGcKIIJ3ycg
QjeP3boqyjh8jnElI6NVDoS+utDOauB6orE62j2/eumcKRqJGmXynwDn/D8O
XAXb2GA5x4H0Vs2Ri1K07VPFZf1lx6pCiY8nOClBNNdFfh5ydmP7VldUpLgl
Y6nfZ71slIQLNG7n/SK3UyR//jh4qeK1hrFdMbwkHzASGrqWAWWWuVp5/Jek
0Z5qveEVfxU7AgHD3eZxzGbN+nwa3/qda13K++8mCJ8oyq0PUvCA9Hkx+lIl
EC1zmg6NidiiUxyum9iw5OKWzWRjZBWt/RgHxj4qBAQXdYFYVnHkcWkCQfdc
sk7zoL9U8ScWmiSbdQi8kPFT8/C8WHUVcHoSCVnjqurQVQlSovoreUH3+3k3
c3h/dBoBe3762s/TicMkdjIlsR2qVob8QSU8+198nOlyXB5CQayJO4Swli3O
t4v2gDUlF319oaoChmc89zr1CRphDjcc8D2JNAeFaQyDlj7PkpnRwOTYsfZ4
75J8zw4xPbaSEVpwZG+/CGkGshrT7pQXchNiLs5bBmtrmfuhBA+ZLd/NQylu
sfG0x3FzkmrM4YQYBaM61/n0JPavK7GDM9oV7dzEqpOH7jpQkLzOQGdoopm6
aVV5LDJKksgWvs+CqZLXlQpcFIlcMlsjJJLYw3Ju60ObGDHv61yQnim+uUJg
0n0oOP97GOZm/6GiYpQQY5DtGmgkledoyx+ZP+ZPlBBBK9FENL95ZsrA9WjK
GcZv9ad2g7nTMtA2wVd/taXAViRimOwQ5Y11XiBkNjG9zQlWkxL04YMf0Bla
G65UgZ6IbcSejQ1Tb5O/++MNGJdAUayNly2GVCdPjnNCiVips5MbCCVmeeDT
kFwJF1Nqsu8yx8Ct98UB91ws9eqsIrK+J2bdVrpgQLakqtkBeBj45CJ6kOja
nQjwyVUYoqtu94+y9GQY9q6Im1H9GS16zqPHGDUguwwlh3akb9P+GhzyAC21
bN+5dORGW3ap7xguvhty1+R6lq50W8HBJl6ForP5Qk8c93GFcUMEKCS0Lfkv
uwmZZD0jlnHhTqDX4kXPLXmu3o5CXkrVskWftZrNS2d1t4RjmRocNh1WaRtn
DDKgxtA9VCgb96zVV7tUWUbPcj4RrS1uQIOX0vf1dg1WqfyVCqATXvyDNa8K
IkGoYDNLzump3ikGw4FoAQKc6JfcKyaVdKcJ5LSN8ZMaRngnGPw/+GyUQhuw
wOUBnvhk5apEMNika6NY0ZxFjhRtIKpohLUHKW4L0gX8OGCGp8ssrjdrfuWY
ASiQsBnOjbUxS/eFV9aZTFv1cUqPJhTmUMwP06Ku5EQyYOt6AA6jrUz3ULxw
KS6QBcGx7+tgP0s/UA/9JUSMqSkywVBE6tftK1g3UrZhmyfDyK9R+So/Pd6m
au4YKDQU3IAh4zHEuNSpEQRq27zK8yGP4htbaOde8KeyYSBhpbYrqJf3PQ9d
jbxoaK8ChKHsUTD7bT76FQwAKzpgMjqHA8GxX8VbASY5MQkf9hbFMmEHUd6p
U6KvYBPg9obP3AxVSRH99OldJbLuK1mqAW8/JKT6D5SwjBFliVo1qBcm4Mrf
4lW3ufteBSQi44ONEZxgj29Zh0i0KQlDcgpXFsETx3VND2phR/5Bi3zOZBPi
ErocacTiho8SOGTewHv/cZ9kUS5v/DCXqUUUz3vCtefrv22NC6JxpByp6fDq
I2bTy11FzNyBPmf/O8H3JrVs2cq3kydAKUU8wLPUONssm/Yr4ECIpWoJ0t6B
dsIrJbRqIzn+be9cXXXxAdnKlqbSe/eFZfuW8zsxXH1taLXYUg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KFoHcElJk+Yqz0hekpgzhYMCpf6Ky4EBoYZq8ZfNCuxYhVHcBH2anMNaQDTJI/2mxzb27+tz/qUZ5xm04B4EuGmdXuVax8W05AMT9nI0Unnd+G1X6cu9QFk9pd0vkD5T9pQMF2vRUjyPRdiIIfNpBldIp+Ytao/q8mq8IQIg3EJY66F0qy/Awj1V4pDS6WrJSXKB6Ceb8DUEd9T28xc2i1YxHtLiXrZrqPsMHhpDJfOFg0AV+Oo+xpXbjRsUtwjAmQEpwta1NR5BDa9JyzwYws00bjGwCYTBs4k8UE//eNeKuJbU/AjJ0vPvkBN+ZJy7EBmLery8rJ6bc71EOISykpoUdpQzuzehhUkpgFEe55/RLOuKJpcVrqRXmw23yXmMGafWktmLBaZTI0y8n+Kb/PvU+eKj9Y17fB4Avl2PsRk210/MbvJu8WaBmDpINbPhBW95P4zyLzi7zh1c1gaQBGCPBb2Z2io4IJlOXDIs6MiIwxgW9y+A8U3p+k61KggMCVyRhi0S/fIVrZAu31bDnWMAz24OsogOiH4lj264aB29Z+OrYiPN61z0CAWirrwJeu06twBRqg9irsDMYJCfREiWMNbeQqAYczbJH61kfbpjbG1tR48S6fYySLdRl7+ClVwQ5xhqVtNg2dM20e/yocCgMijC6V00/MDrc8qhvACD4jqdVC3dFN+mROwoE2CDsx8eXEqAq8TUrKbX3u/XII0QGE0ksHrlVNTSQ4YX4BU35jw0EEvsn3ADly7QcIRW24qpqEPobquVm04bLzDDzA"
`endif