// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o9EyST6A/az8fKveGaEOBg1q9H/7lBew1bFHDFOy7szlclin/mfVQIKbXy9Y
ZWnCSS7lJ5nE+SSmzB8O6wFI5ecMlqknJzmX3mmiHArbKKgyet6iQl5kqmmQ
m3DJzeIxg4tj7v+FboK9zsl6JIoHnxL7wp6hbU+C6AxUygEb3JSzQEURLw3Q
NWsX/3h7GNHnxDMBjdPNTbas/mNeG3laned+h5HoI9jfwTzkSA1QAwnrWFNM
+kKY6sWGPdf8FYf3uajS2b1Zao1aFxIxqSIan+wSNTKl/cbd6jE+SDkFSEqy
BzvqgnIbt07WfENj4yoixkuaCQXCxwj20P2QMkf72A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OU79hMtQTfs6ZAXHn+zQeF1OTGRXIJiFx/tbg+47Vvh22MdyNuWFMYp7BDCY
QT+gBUt4tSNZk80pp8ZI4A1/2FNqXn3Xlg5wCKke//lx9rvFhjfTh17JggBs
kCaTvkzfqxQM6nUFLcFc1c5Ia056ejN8vjXbyu+uyOXFOS9qBXoCu8c2oTGi
L3HexfNavCgrzRSSR7J/N7SxTSQ35J63r8KqHH/xKd20ecvZQbipEno3Ivdc
uoJvJIGTJlPL/DsHF7E5qOG4bCASGEaEADHz0wiXRr0A3KkFbzG9pQ6f+JuF
KNluo4zZbWj1rSdbEdxoB6rxXNrcyW7aq8193B1DJQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tZdjsHziJeDnVVmgIwPwBk9Dv+A/Q3jeluwF+IWVIF2behAO93w15LIjzkWb
pH19M0Mc+kpsT00It/BwwofRwiLFfVYEllNvYXUHexZK8C8QK9FMUz3FAki0
zc2vA2d9UJftbcV47lDZ6web1Zzticemztkg5qCagFEdGSFHI4NizpvHAVPR
GkiEFw5YIib8F350NPPSmjrFEp8adupPSQiQ57cWb+1EZYPE1KcavO6HOePY
Vp9pDYWdaqyBq0ERk2sGy94QXlAu98v/oqTpwZuKyCv+VjSISKYrfNQZd5ak
kxqnD+x/v6cL3Ccw8fmeAbHeHv4u31N1tSTG3LIeXw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FCatTGBE8hq6MQ4QUBpAoVm+6CnYVBRehJZziyf9kXRSl0UDJfCFwuedesS8
30FDpKjQQzTvdFgAEMJEXl5QyxCqKcdPSVlKl6RH3y9w7j4++nbcScbwe/Mw
WTpZ0ZQ7UIjTh4lMa10DrI6hR6bTe1MJa7ti4H7DeCdclt6/x/CrGwq5ZXmH
UW+TYVtsHTWJ61Hv5sX2wCurOR6Pcm3p02krdETn9iXpxJQ0bmub3W3EZFBB
qUbgkPfbNEGSML/HVG7Ov8vlYHHX1pzSSs2WRUw2Wa31+eIpzOvoIAH+CQnc
5cXjY0uXIlVphwBwk0jG926nPzm+5IE/OeN/gD+I6A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PcsiRshNgELcdX6jeMUBT6KEyVaVR0Wn8MeZi/OcEF8wdWsutPVoPM4R8o3f
MQqZB5gjN91ClOZmxoujZpxyNwnF5mYUjEqDYS13vIvRMxqSQ3VJ0iQMQp4M
VUyAKnHS6eEG1Fo1MAeXGL/MAmespwdpZn1u5TXYMscyYq+5MJM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
m0AtFZv2FZG7EEcdxFR72mckVCFqfMXnnPVXNNWJ4Epr+acyOTSi6LqYRP31
28IipggyyxZaCzAuG1OuYxUmOr0hBGQS0QV+u0NQQK1+YGJTpeira+HEoh0M
Lh03A+4FXFqIScmiSaNBxtsogp6skSNOcRp39lVzZV4//skUoTjUJZ3NHKYh
wms6ocXz96t4Z3j39LzLCzxYBcWm3F91R2WV7Gfmz8bAeEXLqXA99GYkSO4Y
OTCNcdsVArruAcpYrTqGK7CEDTah2k78iFxFiTiy5lWM3BpIl0PePrbSU5W1
AKXiIGBs6aJMKCGHbBAprDlfURwAgST6c1DgTsxFRVZssFeauvs07n3VJmmD
R4HX+adznCeL9b/fXC7WfPbs3gcxs2juFZL0IaP6CD0/AgmEgP0X4hME/K31
K8Vy7lkN2UPyC6pgTAyQxBt0V+wV5jRj85ec992tMeTH/i6AgNl/bCRxSB9t
oqv7n0sPeMuD8LCb/7nOAOofLst4RAFK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rFMa9RrdBz7+/PSzhRy173bv3WcTPQ2tKoh0UlUILBoaz54duiDMgTEtWeGD
dvRl8S5c1SDOEJ0tOJjzrUKKUulnLi3CNZpmyO9FeaGVXGBW5fzoDhrwZR6Q
jAFqpHVY9zvpfXYgssYROhXFme7QRUykUSQ3SkdNxlrccs1elO0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
F/ySLtPJz60C35K6HAolJg39ISuR1ZucYtuNb4x8vrrm+U13C+j/87u5f6an
MrrShVS8n3cf2sU1+02+5xsIg5u0QWHQP4uLzXQ3a0/W+74OTdsFktHbftW3
fxaHXigzVObJXUCHgLg+T/WMdykZfy2YU80p9f6BkFemDn0DxFw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
pjyD+5DTMAq1pmz4xdoY4QK7Z9rTRVv9GubTqVdfSsLwi8ZYzS/WmfWkpGkC
me0dwJaa0vJ9mpJJlF1XHCuwbzaKNWZA+ZBrCbVZfdbsuAz5BQ/kWLHmLItW
9mdPWMMIieyvFWj1Lq/YLAV9RkPXe9863KVw1PQaZHJ5EkRPFxSBCcID4Es4
TaMAnEy03FNO9PQql33JT03clec0ZaZHCpEtmcKaTmVmYqnA+IqozkgKVcIt
Rbs5oT5rIRjb9G2cxEWhU7CAGLWAU5oUjnHgEKT7Tzh93ATtiu2Cug08fVop
TrQpOHzCnaizwku8lQPNqN01oXK5a8brfGtIB4IOBLUf0xwjXeUtjs4sue2A
oI0FaoQ7riHNCjZS6pPSKyGBtgkyldAv08K4y8zOg3RPgAUABWzCsUqulLB/
Um4+A+1x8cvEZokZfIjCWRjAlNT6cXtt8NE6V1ArUZCYbtBp1Lnnqgt43lLt
lgsiJ8WhEcqMSC8ozY4RaH4Eq5Fp9kzqwJSU0FGLHqal5OPdDmyFw2u6AseA
m/dpx2JG4ebw8Sd8PwCuyrEywD42oLjxPs3ng5JvXpj5BgcWDMMe+x7cJ/Gp
q2ZJAeayU9HsoKKsfl/OCEQjQbyuCFVRmO6FU6+7MutgagLA0bHxHw4ZW/30
gaBVPT+zq3J2gZzHUqA/dNQk+DKdlgBMaeoxcQ07qL2X3FkXXMI3O+1oYs8R
9MhbrJ5hz7dUmD+CoI8XGP6nMlNy3DH8qQKpgpOpUrDGbMIjkR0sLrrA+KDR
oypnfEDSIAJ6qtoX9gxtBfln8HI+9L3L1TomyIledLHnOBWllV2zTaIbRAQU
0TNKrEKxT6cspI6eRXaSVpUndehs4mPvI5Fdrkf9FtF3osMt16G056IiGcew
h+UzSkB9nCjQAIKyf32F2z8zxY9yljux+EjRXfBcxryjiqbWP2xTK6JSNecQ
CCxpXMRbTR8zD6Lt4ivnS3xyWtyLYFyNXLP2aeSpdQZud7/EYVEXI5IibIl0
Ttjh7MwvZz+Kf3ES2lBxQeOtnd4hQTVca2HGZasmt1XVllECohaP0mKAgZez
vnUe+vkSCvLBlvnrEmSmzRoX30Ct8gBfycPaqf+0AeFWCj5Uql6UNKtFNrN+
G++3I6mtgg+Dv80H/mccmJ3LLrjrnxjkXkbEtaEZWljR7i5VcCQDzFd2roX+
8VjPfLGLuCETH5bes3gZheOxh/fwV+E3VzoE6VkYlrAUDMWDNwrOdBV0fe4H
T7DU6mVbe4k4AcxMjYS7X/o4KttPDjVZOpYZKrHSX18xMc1i2k50qkZTRc50
YsA1ViO53Vtiy0lA7AW9FUW+CxclOo7R+iG2XQ1SPDWNyTqpGEjRMosolAfv
ZOMzOQh7FyM4+4qQI/4tIEAM6Ef478tMhhDbGzY5vGOQ8RTO85DU9dXOCr2y
vv2g6LBmCM7vpdnK03LaVbn5Nj/V/uyELrGOwCoomQE3Tey8ieZ56BdHYeFO
vh6h7A+VEexQSlLLS1KeoBl3pP1nXOzl0rAoRcHHQJtwjHXe/ZBE4OelQbMJ
EclIuKj891WPJgeFC4hM2zghaIYtUGeuMy6si1UqendL8LReDUg9IikLSvIF
EQKFQASjDvvftuIUV0lTZxPbDJ+OshIxmHjOgWDlWZyrg6pLziCpX51LXQdt
QhqFzH6sPnXgw8taOFwt0S/aMv+yc0Sej9qVhRfitkGb9bKD1TZ3hwzaxl8X
PSkRgro3hl0BSpLwlNJrjWtRVmKzlmmFA0tVyXU1x+BI+g8cE7WHlj6+R2/o
N83fo/edG5JFtWn5GgOGFtH9WY7SDERf+YPju/bta6ODT9YbY2r9jgPMUo3J
1rI8RA5c41UTDgD7FgB2Cqrnt++jJ+BAYVdM8jok5gPTlhSfJrZhY1IYGah0
+8Dnbkvc1DHBCMqr0q05ByaStea3Q7Yky458FKAQIoLrnBbzDL7JxsFgXebJ
oGngvadij3gCH+XIOarH9PlYdAuIx0InKoD39un1VY9EaehCmgJu5NOsTG0h
LD6Y+x5HWfscPX7ciFK22PSmJM8AsAxJFCwqHI9jvRCzHOIjNxxzXOBB5pT3
0xwH9YcISmYOaRfiMvS28TusH27gQFJnnlJE0rMlEvHL7KQC7joRLgzZMijy
QpA2RnsaBRl5twng0kaQbP2t9I6KKdnJwSpxqot6fBLjf22Q3odDPktnGG10
IZbRl9Th7V9+donGyabsjhp8OorF2kQmZ1CQhjlxAXVFdeoBR2/nyYPnoE8L
QiBMNAy0psS2viTJdDnjUxxIKZ8XLsHEtb8lgjRKbevhcsFlqKeUwE5m41zM
8RulJGfDOKeYYGbM7o1XhIITfyklfVdV9xvJOWPEXLyTEO6ux07FtNY7ymM8
6EBFpCdQeKN+Qbavy4pEWvALjaTAk2msPo6CPjqt5HX/BYkX/0qQu9O2WLMp
z8xxR9oNQjzwlFQTE4G+0UdvjAmHL++MY9aT5eSYuU4hWdUsyeyx2WKm0eB/
w1gstIrG1yHSGlf+92KspnOe8UFXIYd2C4+jcXD7F10iemdd0zGgigI53q1K
4P2hAhJFyU4Z0tPl2+D+17O5Zx/3rPw4NnLKWDxHaS8ImL6iFVArp2VhLJtG
lao+xjVrGsXgOoF+KQ/AJvHJ7hBDCtCdh0CTopnGHYAq4JXkbPY9ETtBAfWD
ZrL2xhoIg90awFCpsDZxo67t03YBkm/ZqxePPnSmQrmQVFchgnMTtqEMlEPV
Y8b5xG62CO542aYtgRN4CQnZy/DroUo6NeKo1vmZ9TItxsyYrMf40X93G8G+
qC9I5Z2HQvr2/4vIVkO37FuOfDMA+FpSvg1SxH01b8dYFu0sNlnRi/uTjeuK
lX71vxAN7SyWxyxfxoJzGXEpn7YBP0syFE+SdS5SaMtg7u1xyowwEOQAuBgS
9gEGarNaFsj0EPMG27zmJJQf+sX/dvN+DeqwvnCUvIzpnWD35iJf6VinNDS/
HzI4rPB6OAhhLjj1yETqX+OKlE9Rv/6+iC8kEHwzZeOH240u1IzPvv4ByIPO
IwsTN4ojO4qRkYUDbleoBGRYa+6rMW5P2UUpH6Omqgi/T3x7lOfr/5BjkDAD
oD0wgyKehMDQ+wUywWJObnEjZRt26d3+4+WJ+uj5t+shnrmF7F+kQDESIHxz
ioa3SS/bZGosf1YNv1PKKkJXnLrOrcpN5jHoLnABlhX/kChlhe0UuS/FjraS
ILipZ++GyULf4PyI23MxY9En7qXuODjaOPkb9VjkFVk25Ao2HJ4RWlcUh6Jf
ZD2ZnSQfwO2/tMcdAYh0Lle+9pvJeb1U2yC2pRwcHSInoDjVZTyzPO0x5qTw
ODhIaRXN+Q6j8kRB2HcxBdjHNaXOIUbe+k4fgZWbrrZ1gt2E5ftMv3VNvt4C
dYBO+zDu+TxltYfVZUE7b0wZAVOdlZY0vKvEEkToDMScpg4OkkzWp/1skTOn
Sdf+VM7lemphHLjqYmwdQ7fbCwQ+ld20Edj5uaUk7VymYVXgt+3YzUhHYuJZ
rCrvIQ2gXrQgPtJrT+sMa+QApi/4xxfIjJ6IVv35DTZPMzeCBS23dZvb+B6P
ONv43jueDUTYhxC+h0G+Ix2xasXW7wqbmVQm1H+7/LSZRJJMjxdtBrtfBTcZ
1WRvBCseQVmtFZUE8WTHzMuhUcZ5PDRX3WK25HaCyFEeOIfqS8msWQQ+tT+q
niiLrrIg1aToZ86CGqNMcF7YB/ei+hP8JRLetr5dSsV2Bhw2XFUIRtuC+5hI
DiYaS3bI9PlbjXhMVFrUAsqOw3xgGBBB8z+J7bpAd19wQnqa6ArnRwH17Isj
Ub2PpKp/TRYYG7dnKIEeYcksS+la8zDhl53AX3UY3adE6rwBFxKo0kBJfbB5
rR8Rq+OsPyMklBxW120/j/dIJnUtxEgvrNhZdPImAQtYXRqwIrP3K9mFBqZ+
g94b/cVkuWwkCgDaGf9SXlrsUIZUrV8HQUNGTRYdAckhT1Uo/OSqfTf+p8Xw
ieWWfN2ihpPV9W0xIfeLJNtDO8dTg48RBTfL1bkOKyUT0eOQlf1aBZEeI88/
UxkaoJu9DJEhT+L30/xs5CY+8XxWQd9yj3L3MF4HNPEV9HAIoFYftvjh2+vs
vyUtYj5suVrETHUeHVJmyeDq/+71VwATT43ek3E2iuvuUw0jh5Jo3vXU/sey
sBfkD4U9W/Fj15s71nVag/ILyWOvEmhloR3/adE8imZxTCccmbNwY1fxSfzs
R0LJKbR5ORzhDziDPCuFc2EH0vgat3OQEyGvgCozfanXpN2qVbb9dNYBugDs
nOeJQmDvwdOTw9dII5oGUTs4KKPJZq1cvMNQAyRFQNkq7hFnnan3J8U6GeE+
r2YDefxfCFwQRvFdzf8veq6bs3cDTmf8VhZsI9jgXHF8325dN85m+I/yvX76
SIpI3BKFE9y0HmvIm6aQvXlR5+WkGNzX43fth5Ht5vrBXe6EZkpZiJkoXOvf
LhzSSBXlAeVLzIiMVBoPdZ+ZtEuXtl2j6jchusI1TykONm4MYXSy0ViQxE5l
YjWUyehQmUmGiaXojFEB7EgNsUwCoAsIuhLUOESRTrDxlvtkAw/FFyAS7WJe
jF5cRsiu3xWDaKWHYocqyjsMZVADsSov+Q1Xef/Kw2f1O/X2QqsUm5lSCebs
741MjFIE0kuNskOry38o12YJGa/KwiDYotipTJILXsA/LA/Ahb6Zh3HhZrgn
vaZb68/CiBHipXJwpYVIs0h4TF0YFeADOqaHBiCQBA+CtRE3vlxf0vh1EN3d
BD/987AAe7At8yr7H/MsVwUiVAQ5xJSJm5FX/QEqIvQIAe1EEHt4h5sy+nqN
bXAGr2KDLB9sxph/sg1682HXSi1jE958fE9dE2851m4Y2TJk4H5X/X0s6RTg
vBmwrzbmz02FlEm3HRPBTLqW+pEvgZWGBBtH0DlAmkHMBh1w2FnfjREGlwN3
OpIbEgjjhYH4jerVY2K5XvQ+CAhkjZ3+57Tt9ul0fuCt5xIh6u0BVFuVzUtv
cU4NZ88NJw2zGoWM4nOcsuvt7uigxFeKEtMK0h1Luv09Jn05a4BFqWd3mPK4
2mpXzSo8lCJ5c7wA7gMObMwDd4oQg7m1+eaYXzz0eV+C/uOwIcRW3kFUdt+k
f7iZmCbZqKZ+gWdx8R580hyjqjFzce2kX4DsgOFYRu7SIclWsRMGhPtlYqgS
vlJ0CBFVxlMrGhON5Rhjq6+NOMBebvyREbbncIiAiQzJjVV/3ZFSLjK+tcFo
IzwPaHtQZmOaH9AgUP+ABXw3yhdPYAfGeTZO2h92kgxY+BCbLrZr+YajatcV
Z7fjgHyW2oCrcr59HyGsQYm43GgemnF1l3jy0Usp64W26dj/T68IorE0ejJf
znn+IxARs3bIvpNFVclRpytwlJ86fhbk5C/taKyCj+MeAWzuXVXAo62fv+Ub
5Xrsh0Iyn8oJAV8zblYUPVZwT/MxHkrex35sUDcUEiqDL5/4ChxNmhOK1Dq8
qwpIw9lcHtPg8J9qSohRQi4yEXp4oNkk3/eLa5GbSyQjNjvBib9AKimsZNKo
FPm6qUo6nA6S/c2wsOrFSxPbBCl3+Fg3alcq4PgWJo7BGSmjcxtmr1lQnc7l
E7eJOrmviBc6bqHADGwExdwegwCTYPQ1fXxfNo7zSndG/QlQtE276eCeGf4C
7XTk+y20pjlfeFiFLmvEJC9W7zntLRZ7ifwAusKtcyJpfGkKDV9mvzW0hacz
gYXx306HtPaiwG5mteIz3rM58oQ+PmF916irWqlMfNe6jDKzUbbcoEGmzB1G
Z5eOG+ZQJvVHBASJSA12LW36lORHEuZ86WJdUtniiE3oZ6VHqpiKV1ZKz8QV
1K7t5/7wAsZd9CxP40U9bBOqo5teIwI45DE5iIsSmyD7oKD/ELc0ngxmzR4P
aSUyLnQkj9r4k3XX/hvr9YxHTHLaYWjvspQLc/e8uRGwZorbhORRx4LiLmnI
ZC+OWbz8gWv4ThynxK9ntdOSQkpAK60BBUm05A1uBz3aMde/0SYMMH9yS9sh
RiAqE6JK+5m4eTeCIRM/RUex+LBbowZzK99IFS4J2S1Ka/ZBOenETjIhXVRj
DgwQC9NeZeaL+W1rXHvEHxoc1NVpJJeWfU8hdmRjnRvMTaovzhhj/i7BSMxK
GspqC80auEDxd1+dzmPHKWJJOwpRREAaJDjcHjrR7KZu4u+iy9cyf/hIi80b
zXwoDDdQeMJa+6nx5UP4pUZr/EHbTBdZZrnKfqugoXkzpKSj1UFxM0z0JHiw
94W+7X4I1UQExEloGvgKiyBm2FMV+ejqDKeQalfKowUppwHce95jJlRMe4u6
J//tkfD/xSuo2lm5oHy2oNDqI+jIyJVQWTztdlHHZpuQNU5anl6IZf18V+7k
GY8mfR7N+x1ssCZQzhFiUb7twVgFSKHuza6i2/iKDZ9IAEvFLTYs6HfQTIQx
q0UHjgB7uZNMnkTlZ1+Ppe4CTHfZgQKWTbmndUUOXAvw6OL5EXMhKqa3lHfX
HlDOGAemLGJWMOHQoc0i7F7OWoA9WWHcj37rSiVfBBt0EM1RPNV3B3KTxWxk
FxlAGdDGeIjwXAGRzNhzyuu5SnQfZU19WKisMTH9hlQjYkWellI9T8vDq6fe
hugG96Jby6+mLi811UYL4VKA9J67VrFQhUWZBCj3wBbblkGMAkC+8Qyt1Rcz
nB4Esm7h40KQKjmP1jEUbX0SK2pNiNaXngN3Nh2L0aRO5cpVlBmwPnkDrQn2
zLbiRfZA2bwYMRN0sBrtjQt8ASBU6uEdB4M83CfRjT8u3SvUE3nhdxQAjxYS
HG0NQcsbjvWV+4VxXYfgYY9fF1KZ+30O7lz41dQj0Cd3bqgv/m3Q0tV+QDUb
CBXNWtSbWi3rSc6j/cVVz3ywUO/s0B8PqxuPZvNF/6C3N+M5VZLuVCJ6P+g1
Sp2HschedgifLQPJEzwG5VK6M8pfXUKTeLJnhq0ECzsMchQ6gluPwMEmTwoS
ZePMwbr8hgNr+sFOH7CYrk7YjPxqftpsAEUXXV+e9BVzhj9bnFp2C9x+s4Mo
6qukgkQ85VEw6lN36ZzqnXMVFkgPlAeqqtmT8ZOYfTZrMwHc4x20p5EQaruI
p3eanRASvW61sYy70e8BgX81S1AkvskVHDqhNcFBzbEIwkdvpJZkLDem+yeY
r2zXqstTJNbD5fXXP+EzTYAtjd3QTq9Mum4IQA+3L7f0o+09f0qRXaX/Wyst
mG1vnCwtjfyCoj7A97wFQIGgcgx8GUbyEsrOFbsDPrlvkbPUpfGGm6nk4Zf+
BjC9YTNPyLoYH0KTjaM3MJQU0QyM4c8w36n3ExoK/+46DfzTZglACXvVOFsX
cYtZG7WAJ6PS+YShlG5iFoQ1DXe11sHdWv+i/rdXSHTBqidB6345Dn5QOsxY
uegz0K1hgPsk4jkEpdiR3vUXVYEiLEuIerLFpjNVoRD7TrL9KxX5qk+7/iGj
3s0CYjKmWjpFdx0JKVgWOFGGToW9Bo/JC2IusEO+0lnq7riFThyBvTbqRThb
oBkzmYARQLp024xaFcBCYNTYQWJebz+umjAJRvuk88iQtZAgGsHHqMbHz+n8
h9szCBPjSqXot1teF0BVhSS0LHUvV11PkpA8gkcIVQJ4XT5kD3jJbO8Y5Imx
MlmsIUdqjWoPiSnTBQrXSVjfiKGauJ10be9cdmw9Wt6Uv2NhAOYsDMBKNvdr
5f+HJ1nj+D0S6oGjokhWk2RnbMMThSezry/DK1RZcQntV71AZj5jbJBXHKqT
69ZJnOBaKW+UKdAjRJKcuLsFnDg+Jb7QCHVeO1vrz5iLJbWF+TfZsu9OJYJl
oHUu7OQX2lChpDgVyAFpNxte/1XEe4Qv0mgiWxNtjQqCETYRDIu4KforCFkD
sXoY3F16TSGLgzQECqkJ0j80jcLubtd/bqHa6EQdFb9XKal9F2qLt4OdZ1UT
69v/VJTjg6oQsGEIYyE65/an0Nud/QLQB+LRXV8hWTC4MadyBFKUbhBF6ERO
Qqv52IT5n/kqIv4vXsv/eLbcmvK45578QXWanDKN+Csr7VvUizmFKRdkTpu9
c4s0tOXL8rfeBAHE8c3VienHYLQbpFpWaKsnbTXWSDJgUMmfM0Pp3AmWB8vJ
sfiYMmUBs9ObVaSMsRQyMaLQi29ARVyvxx0+ZnzthyHULptZ4jQwbDzvpFcb
C9yEu3DnyZdTSl6fdPSrmaCDj7MC+ITZRHR4y2k7aELVuff+OeBYU81W2WKC
fVc4St93erkfjeVQtM8m4TaBTDgguqkhp0LcytFx4iLBLGl65w/0CO8yPYFk
InL/7VW1hDof1vg+qKONvuIJo8ROO6HqUfG1kHgV58mnJQb785JrXsJIf94s
8ybDWyia6rU+IXcPF8LROqBhL3w2IhKFNiUn54NbmFEjohkxcrJBUM6HnMTD
SgEd7wi/9k0veCPFt3UUzLH92mlk7NpFuxSU20Fdng1N04k0Mgubnra4AXYz
KTHlq/metVMuuCz5DsLcj2S7WQaMg0APc3NOCYWG6gQ+4wz2S880h1hQkLGN
MxUeUbhxeDieqHUYaobvGqD0mXi9jvBSKHvgRxNTujOdJjXjTZxJs8W4HSIS
KnMon+9VETmHFkmYgiCPdUUQwxgHoqdCSJKlPthakacetwJ5/GfPgPEwdEA0
r0W8Ke1g/N/RI67kT0MlW0/7LFFbVh+yIbB/GdlVSwNvp8DmvorYNRZNdDSx
YHp6NiyDMe5BBtUqdOn0ugOOor5xp8VM6WWM50awxvQS6zU3+I1rR4Fr+aJ9
dUxoYtix9r9/LKRYEUSOYra+qx4VVvdrTzjwX1Ffq2YE4DUjF2Z2bvgyVv3w
ZarL+wC2pdHIkJ7UBJVN26NLl9WsJ5JbUrIZIXKswUN5zHvczEHhYS5uYuAI
FmTbsvfqNBVxWIiFnMy7EK0aBnUpx1XoCmC6zaejpRt6A4mUQa48xvXXZlsH
6iErZs9S0auhIhd11f7dxl3aZb20xTzcudn1IXc5k3gtOVv4NjpyUt9PagAu
va8eVYPaYnFzsX7+vCKQjNUONJ37UccnFePvQPB+GRHfDmWqMzIIfc0zQxPu
2Qdr7RLd+k8khwF0ktbfm2+azqcpbPUURg6g8ESFE/XhwiW6f+W9316184Y2
KBjFkjNbokSWNiFWoycygD9ntU5newLZuyIASKcYySLY8yjrfDbLTD1XeOR+
uczXeAbXj309t1Auo4I6+wigLMt4WQiV4Sv39awODpP335jz9zcs2L2ppZAj
6pXbXAwH1rAVNqPOxNnl/eE7u5cPTF/qgp0XMjCxFGMoMUy3VABEe/8RjGAQ
DA4DDtfXdngtQ0rlXgain1dShRwJkuiuhBl+pRIpe8RqoVzja+M3JNyRVIWv
D2wFsCISlIboR2/IRX4ChYOqqiOoH4kvW5TLU1qtERAb24T/Dr5PI2coxF3D
UD8DvFQALBSeOMZYnhFBRXAgvMlCb3AxHhMJBbYvxrfObUXeZqXKAkmFIIxs
WRNVkYDh6wSjW6oUvjzS+TAVxtN9Ao7JvGMykXUdKpuU+xhYMELssdDfJuVb
7oCpJg1S9+JOr7rm1EDBIzTucy0JaVYWcoP/EP0DBFg9MUsOnZpfTIn4Pkw1
q4j2woFmakBEsNNcaAKTMqDwN8lsrs3Kh2ORYgWL1GJ5MfRgfHRTSlfXsBHq
TX+BIyfHLbIKOOBVO1JXYTSFIvIlEaEdjjxiLN2/cjemREgIGpEe7I3fPLU7
7nWkS9OKYYn0wugUxjQVWtGsKlYFWiJWSshOyhbQIySet9gR5rntwlylbOoM
u2faOP9mgoJDM7AmcRmt2Uc8m5u/NWwfnLT3Galw45B8sK7pYlhuPLyBxoP4
/iDxXBTI5NtsDwZBGb52XqYfDk8IYcGV5BKf1snkubanPs0fEmfp2/rDcQkL
AuI4DYRoB/PYas4CTTpiLs95vvRvnEyH5dv3t2hd0RVoGpUNtgGiZyq8rPfu
iUHlV5qq0RWZu3mOjDTquJYDBRm2zQQD+boTj6DvxXZI5wrCa/enLS8edNtS
XlMWfvYfbCiarzrgko1m0AMKSjeHrRIbbFoqJoaijQCsonA1n6YuLIwMX7A8
cBlcyw+4ZAGJkZZg1ezvR6ShRRsd8a85fDonemtwbUUJuhf+Rxfzj/Xtfv5e
ulT5R+q5TNfMxPIyf4XVBfZFow9rBQGMhCyTI52d3opH9xkWmzM0BP/Itly0
gzcgQL7lFwnFKz+DsTk88RZbACexJnRmLkK3tHVAMiHkLEaQ3T5Hg3pE/8HH
d3tiifthdlHN8W7VBE0dVZs/YmGTAYxIagqqzkBQhxcHaU7eN4Hbm2P4iw8J
7gRU0n8w8pwb4ZTlwVobL32pTCGpDiJ/mYSXTyioibkitBpBvCuqHpahm9yF
cLZ8vct1jrkPwRVmhA07aaGKh8WO+rNvKqspKc69eUbR/KrTieXu7vEQpb0Q
KtIQwvM6nmXeV5G1HOL1pOVVcwAyHvA6RVbecEEfbdneForFIUAak3ebpzn3
gzb9tgVpWiwJAvQCTyiOomz7pv9YSXGxzZ6clxLeFgx0u+w99fYrXGsKy5Vc
xjBElZG3zoRFLZQk0lia/C+AHWSePUmhwL1NwQEvc1V6x0TXWjSqKBZ4c4qh
auN6ACLU8DLgdukJAPsfFoiuXVjqFdH3o0cbVKd0SNedeIVV0AU2xdWU6sYr
6Yc/t+4RELVTnC9GEL5Dty5yLrHV8QUCOHSobxOOgTu8/H1gYp62BVaVTBKd
hKQrSR7GyulWgO3H+OcITd+BNtA7OvV7gdfnHxaEXUBumi5NclCSnnwpuHTk
JtvuZsvUPjvzYijcya2MAxGeQahYcjfvbQP+JeH5avPswZGL+9aeUFQxraAH
s0ipmD1ebdQ7Fq7SPgBcIGd75xtpcNfYyQ4aEcoVoFNQujOLAHqL64dVBj81
GbyY1FSI/+XEKQr3jdtR54Q5t/OVnmfPhyK/Yporn6MUpzyj8K+uD3IhFXUb
IF9APvGxyECu+3Os763Yy7w1GHUVFU64PRDqYC6GgarqtCVK4VEjpyepw9MX
pejwubBhrxxS8HHxkkeYcyxLueLlAjKtdw9fjCJWzQmglCk0VDB20+f+2PSD
YGp1eW8ue4BkuJxY9T+sjcsCWNcs8drtYDSRe4iGo50kJ8Jb2ll5OXtnnw0A
pP7cyv4oQaU8kitoA+XYUyX4AAiVog5V2blowCWgMkYf+pJsRrMmX5R7S8Ef
dvZU6X8WupsyRKPvt8PiTwVM548hzpvD3inxQwjz9XAHCRpi

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzc6UPZA7nwQw31cdD/YKXJ+foGDjZc24J38AY+VNMYQV0fyAhlLtBNl6/aLhMddrUhTPcVSW2Sfb7PNlnlpWeOc+XhU8fW0pV6XiDiJ7Petu+3PEwKze5vB5XsCU86l9Xwb9aDlcQAUkbBDbr/kLndSsLfNemwX5A3iRvIEm61pldponq1plmR4Vy0lLWiYPdsVyffplMTM0IaJw7y/J7wsGsEMB2PTt23tRAz0UhSB5GLaKcpEo7CRLc9B+BEAnPQ8cJD0+ctg2RF+3E8f02/C0FWyglNycC1sIuIQle7h6vFB9n6LSlwt+uj0pfZoT1mwwe2YCrRXbNNZunCOV0cUtq9i6D03D4nNRdKiOSNS+CBVYODVbQk/FjVqSE3kRWmG3q7qldSg5Wux8ruT1KYbWfqGDMfU8PSmaFJ6BcYMVMZ8JxEQrILDw1Ae2M26lGzgVmdrBQWdUNe7uhnr2hlZ1j/VlJ7zAFhQmQCF/2SGR+6lhzDrwLO0QbD6NIJudIQ/DFKz7Wsf4KGjQTReqOR+G7AIfnBj6gjpQ62S4EWF1axdUd2BfFWTheMC5L8wcQrvfsS0vmDIMoLQ8yJdZTqic0tlHz3BU8XS/9SMbtKEOJHbrbxHtwDh/IJ8NbSYCJG6jJzWs4UQlvWgAB6BfhPGKAvtQjxkJ9yv6528pq/Vzk+/nGLnmFcZe/l5J3yDzbrHCnaZvHLi69Z8bQYFMbM66IBSTtyjEHVRGe4W4V/eypoHm3mJOYQ4ew462IzRrKbmtj1gro4duhG3fd0dlP/N"
`endif