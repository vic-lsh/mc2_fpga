// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zUw67PoMM9eKbNBeCyCXU7UsjIetP/g/2PZFpFB3O5nuAGlIHBrvdo1yc8EK
LngaCiO16mlB0MTrHYDml4JoD2CROjdeKpO9r+dJhpAcqw0m1q8fVZelynNK
dncNE+iTOBHvfMBLR8uhe75EC30LTMN8VKTiK2OZ8K5VjxGXuPOrMGkeR9kN
vT5Ib16J/AywHufHx2TUBVm4cmH9Yez5UtVWztxMW/o5LGxzbh9UVVTtsCjr
VR6sUvA/y267seumOiLnb2FNKQ2L3fNB1Ho7Kjww50VQvColjVnG5wVqOist
PIGj4d9J6hx+/5LpzbAFlFRbfKkAyE+oNhby3j/KSg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HqSLQgHQoSDBp5C2K7c8Z+rllGGHq2JUcnkQfPb4rMaFFkkq57qZOg9Q/7oe
GxWAOZCp5JToGT7J+Ayx0v4racLqI9LHIQ5V1TOy+27ty2fcEXEhTQhKDh58
3yx38gKt+9C1NazwRBxCvXnNrJDjALc14CKJk808x3gx7A9d83S0CSpwYxP6
stpQlDreg5DWvYT4BACNd4yjlGM67ub+IQvx0PMW2euENxijkfPYfIZ2roe8
A/guO25ZqPSMlo/wc3HXUGln+Z7DV6Jk0/5wIfrMmNwxjcbAY2TPTnGuvbS9
hn2LtUB6ixm4Ns33c+USzglG6tZsgl1mvRtO2VSHKQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sYDw3a4HzeMAwBy+g4DgNqEODn+zIzkN7hAVJBhupwXmXcmzFTVfqg/KZFhZ
oIgNRKjPZ9vN0ER/apTPv4ePTGyTSGxbgqwPINhVJZLQvGOlchF7cKp8ikGc
C04tEoqI1lHkM+N3NZ0n4fQ2nFR84smQDWGC0481fCd3vc/EIum35+skUlMD
i/rNF23u6rmCEasSP8DZ2tjSp+l+z9fFj8Ag7borobF/J/DxuQPZLRvf5TPu
6qO4vjAXzSdwYeBNyY8ShNP+aBtRXDtPPg46kZIGpNXeriIKW1TFcpCIIx23
GOG8qq9fDU7qY47UWZwBSpxkLZygrwhVX/8z17M/fw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E+YsFXqFIJyFBibOfFthlOXnmL1vv83FC+3LMF9UFwoNwbKM+YPAjE5OcCuZ
MZj+McML5EpQsrYbG+mACwbkyNuh7kl921ibFiHN05I0kO9SdpF1aZi5RMBv
1vjcd1CENK9FweD6BsPadl3dTB1dk4kduVZr0qzB9l1/zcWebLlyzzur4lSs
LHUn85QJNg2Fe2vWDPNi7vbfWCgMXyOuJ2rXBjSgrx0k2SOIwdxJVE9wXDEj
GlQk5Ha0gnWsXU6w/iKZHfVfFGfGCsCsb6aDg+rFReaEW1OObXJ2fJRNCWQr
MbIH0ud5IUVL5zsmBVPw7qVfP6j6sVs6az3Kl8ltbA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H8a23uBZNJaCCav/uEAGrCQaUE6n5FNLU3qwPQ3t2SbhSPECnPpntk1T2fPj
8KjQw32/T6BF2ABon8hT79KnWc23DDb5ox5BogPbgi/4fm5uWDdDqCMv8B+e
lZg30KCsEh+dZeBuc6hS+G+lx1KxV/6QkQm5Zi2Es6PEC5e4PH4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kTAZn7h3s5N7XGo+Jr/R0pdbb68CuoyNuSJaIWKbavHNiGRjlgKE+SJPrDdf
Y8hO35Tf8gft2ytNT49kIywsdpZuJyZYuA3mimR+oSR3c2daNz7kNFXUPK3I
cgLSIU3ZKjor7ytvp2EoohbvfFjY+cGIZrypGV3z+quDbQavmv2Bbpas0a1e
/KPGSeyk01Qw0A1U5U7pFKB6H3cdW/Nk+QVmHjsqNRDxFOOETg3IecRnIfI2
Cy40rbvqQDVlZzPhkMNyz0JSiH0BpfXf7ZsW6oeIf3KbfUHHryJrPuR1OBFf
tDHaVvK03lxJU7eNX0cXkQG/REGMXWvK86q9eeYtKarxM5FR77wtOkvYEg0N
fbdoADraULH0vg8fKxy93Bcd3pWhxnbu9tj9MDI7o6qPKYn78WqBwMZaEof6
XTPQNn8hBMDIETSIyFZ/Ggf1SFiVQw1SsdL1B+QelC6gaGt7qhHGeQOz7oTt
Ud9I5wEg2FYVMlRO4fL9M+A6X/BMCSPP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K48A8rbph3L2eA4JAykMgYIV4NGi111nvUzV4X8wNmVOK7vAbp4pMtpQVcjf
r0TZtQjXs1cy924aZg2aRWKaxvqa3iQzGS2A+eRXYR3J6/xPFTofo6TvUzW2
vlsTmZ6/hOhR1hR7NJnl09pvTyi19ZxP+aD9hluYegMR4DRhggY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sTZPgdTUzlUgqBEU66D7kRWcdznJQMzEpxOCEJ9xUaPgm+5+YHPzDaDdWTiw
zlxrfSXFP2DxdqHPmrec540BvXUfICqXeean7sppCEyJ7NkQwVI5poFKvpCc
UniCBKib0EVzPbwxF+IH8iFtjhu0Ev7PwBTqAzSjobZmApTEOuQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 30944)
`pragma protect data_block
6WCulsKTSFCq6uBYsYV48+lwWkESIaUnbXfzzfqHata2ts2z53P54MlVqB7E
O3vX3gjtUp2lprxMtLfBQwFKCiSDoGb2fSJzuixyaBUvQDkUZcDfp7tUBSuf
TrdJLFOUNoE3K77YNELhkwmV6O75i3zeobXKOeLzoDjFClzYf/bJYkEH0wca
AMqxTqYELoAgPGtzZxxHYXC8fTUeAZZ7BG5oRpR8kZ+3QLDhw4yNChGEKX9F
1F21A6lDB3ad8DGv477jQvfr4Uk4UpErk7N/Vcvhu8wMe+C3V4rAqDBEs4fZ
071vS8Qw7ZOgf83ChPXjP6/1XUs/NDw+YXcq71AG0OinGmSb/aYKhKudM8mh
putVOz1p7TQL0pT8Y9icrahGVidp/a2qIdEX3Pr5kGI+ftuXBZYeKzxY2F7O
+67nvE8K6jUrBEqxTOStL3BsTFGP4QGJLTl/bschVlbS9XtAxP2Q7aIaCyse
BUaoC7OYIHOUpiVhLrnSWhmseUR2sWStg+cA6tcBwqf0p3veBbUVWwZwNx5S
rOfrE7gwJd5kk6QxR9cbAQPN3XTbRw8nnAxx0nXhOInRm9jJT6KdMI6H+s3m
tlz3Y3rA8tE1TOkSoDjSBOuoWPy4iTsUzEpI78B9KIkcGs4uVY2ITo6W1WjQ
SpYRYDXzmKmKH4ab3VIrfZpDdYZah+fAucViO31Hue8BdWBhvlbcEsN+khPq
8J4F9kfF8oEt/eNCr9i84aiedeyowqroU8aUMgDV9yujQ5c4w6eIdomTqAJ4
6G8OGXudyU0euAv4dw4aYUVpwSJbMJnHUJHX0kovnsa/Dzt4a/xJ25yielIs
QH1mvIIgYsRpKHSYIIE0jVO3eC+vVWtOcGRuVwHJlYzDx0DcTOZKiNIl9UBR
MhpnZNodbvrngV/o4vragRz4uYnURSdzksGjKfSNHOJRtNi5G+rCigU2QU1s
4ZdJgp+t5epgI3/ZV6sHvCrIw+EG6HG5GeG79ktYe66GHG2AOwiK7HcOVm7H
ZHvKfck9eYTsbepEKZwSqOoML31KwA2Sa9+tsFVeWZ/hP8gmxRJC3e17sCQq
4HBTsNMwzCq9FOSAM0VkuWdlYin4IHnZoiF+K6siBimeVqo3t/iijqfDVsaI
O1OspXhhZLaZPFZW4Li+SkqLNQctY7qFgpkNuyOne4Bbln4y0n+Laya/jg65
GD7MrZ3XzLSEWePv7gwtcnElD/M83agheAxcSWubztr++n2lO8jJwitkiFF9
YAZgYSsUtebZGnXl6CJ6TyVSbWnhy8w9MmHIfi+QactLMXy6vzwRVTcBJgS0
+AAeReYTPuRT6SY3hCKNFLxVIiA5mfHQOeS2KmF6f9wbjhVbZtJm3Zp+rHsf
x1IKLizt2FiTjtK2RA7lH2gMpaeE2yDo9rMQjza3Qi7OmDVrDbUxkAPNfiR7
FbBKj8qyloHvXX6jRWW0Oy7YfbLjw56YM7b3MEjafDwmjCbivbhdXbNzd0ZO
yYe+xMEwleQ1MX03xQHMcxL4i39NW8ph0TPRuoIjlUF0UVPZeaXJpl+D5qlU
V33XSEzB80xha/fPvWdUViaHbU/Km4Oy9swOq+RxEThf8D1Hn2iTjmdE5aQw
552GZQ6fIF2hl9DM0xP/VZHE4EzXoajLegeS9aGsx0bvfOnDpAKOuODlJrij
4CzT8dueKKY3SSO69HhoQcnAaXDs8K7/1dGbObdMTfTz7HSj8qAwZ+uXjDBa
HZypmhjo0LH4xGsKo02WBEZm1S2TmNajbMeXabFYP9ab5krTbx5qZ5MbEgje
lCQ4qphmiyoHDbl0wUVg+3pewXwKQ8kRTzZ+0hHtlYate5YBLfgzrpmT0GvG
UTbVLfRN6C0hoW5JnT/Ox3Jvydzg+diu2XOn33dJdw8QWpcZrRCCAM+EAtrR
lCOvSkW7C4yq52mNEAUDH7BQrmNuVAsOADH4gBDVE2rMogzBAAFor76hx5qD
tkFgkeFLb5nDKODIpnQqAN9w6UEoYTCrJBeLr4F9ozFn6saecW8owloh3IVP
93D1rmO8fijdSEl5YdGhkqU4XdQRa8OGg+RJq6nLFFBdf3O9vK054wRzDlCu
M86O6GJ+SU8CML3CV4sSoITeQYtrYYQV1kMtp/AeKViS4IRpavMrznLKhiNy
+Lf8NGSaobyaiAeJIi48zjSHueAJ9vCvqzp3apEvA4/GnHHk/IqmigWLzRTJ
nn4eexUc9+bd2qs9YRyPb3xVJBW1IryXEqvBCf0p/WcKV8BbPbmwoLl+rXpL
p7dIquOk6V9wbNQ6BTPIov3T/N2w0OW6MbcySX7brzB+8xb8Dzwom7HC/bpW
+PLWVH8rbtaCiNbNXnyuK+Vg8PQTLL8vUcw/cGrH6kxUt5kEUpcBm+w7teAQ
CoYdrYxDU6Tq7rPcX3wnQl6chypEUQ24vBsn3n9HBsA2gPGSb+4949BGdJtc
cqvxWcsBNKBi/clkE+l4KKrkTuFr9Tmmo3yDFTalYR/YNCEPMMW4YBhoD2PH
LcTVXMAg5vtDDXI+WOcZmSphnF5QyRC/UHsiL5KfAoSjxH/ZIjvolYdmv7/Q
+ATX5O3sdn9/u35PVTdxTz9itRItpoUIh1FUFRoSGPOV7YMFYnEJVUI8Cdx4
Jr/yeDsj0TnsDYRmc4l029viBNDNQlQZfMnmDfuc4joy12EaUby5gTKw7rlA
p1MbiTTFdqJFkXUC3R8AR3iMN0+LoPDMhK0DWVgTusdLZGytrma2p2O5pDGI
sVStvYQi1yFXUHKl+fBcXpOiUuP0tWjH1731XI2Ln6Q2di/K3V12vwYM3rvY
QuPKEMB9tGCBlORoFUEhdE7e4r8gJO1UzSS84skp0ECQcoazog9PdHy5fxfX
s1Eg+PpLo4B212xLZ0Ct7rSsnYdWH1ENiYN1L3p4a+RCtl6IuwNRX+nOdQ6g
2AQRIw67RsI7QLH4A9Hr3mr6dnIs1pSOQkKh00R0nBJLKGATWcrD6+snDgwg
Heqe0zSlQG0Q6Vr55nF46GUo7dCUGwU7s1Ig/LYiTCYy7av+2BbCElaEEKyL
7Lx/R2m9SRxwqHDiCPRh26cnYz+O7bEOhxA3BQZ/5wnptJvtDApiqIKL4RMN
JdaYRB7rjoAeduU/B2BEXRlLu7qwhJu+t14gMtz23tjH6gCQaDGFP5SA8a/0
BfDDkF2N2tGLioNNgplE1k9t1pvvjRJ07gzXTxTGUPCDRTAJUfpnAnaq/7zg
BBBxV1m2WyzSXuDd8wD465JCRpcIs09EjBryorI1drLaGXtIXjGDSM++sc7K
T2ar8RPmx7Q9w9E/XxlV69WVFiPWEKK0b6On+71RfBD+5Mh7CrDQcnHDJoQV
w34mNRwLv8PcRE34DoznKvRjJpfnH7t/keoPpcMFYzkubaRFoJagoq82pebh
OSDvxL+f33w/GCXA1Y9tRJi1QOATiQHHUsCYNXF8LewviT0NVditBnd9TIHJ
a9QlcykeptXZppwd8xpSwpXknnGY9y/4ZeScIrwqZMlE09fVABmPVxuDRWYU
p9IABuFXwYlxsQIc2IQzkdUDt6jZ2sWiazrUt+sLXAn5e5YEF9wZ9sVagDj7
nmHs5BPlGBDHICoS+/xb2rbM445+HSLbq0UQP+hgA5ELiN6FwhISy13ZhkOD
auiBCUkHGtpBEcmzyQNIXrZieSde7fJgNd4qFwuPXbl6S0EJmVKu2gQzWfhi
iDZBfIq0yHo1ECJGpqTlmxONQhJjO69Qb4gwxye7+uQoxddsZTrxT2bMq8rz
pxpZQ801HZpU1KmYpbjqk5OIPR/z5Qt7LophiYbeDGENKpdmm+fmUmJuzAvk
OUkbfXWNk5NyK2ca9em+wiHdb+oCqYwgwhhyOMqCG6kbeP+waPDw5I8vlKL7
1RtfmHCP4DXyiusY+J8h2Q66GygEuWFJ61WT5RDZ8CN7RQ+bf/FBr9MgeL1Z
V+P8X6xjoRwIVqmlJjXr7xld4Cdf5ZzLX4S9nXf4d493hSEfzX6MbC+yCLJm
MBcXiLhCsz9PcsccpzLJ1A9BxTHHigp7GfDXhbZkEYKm23Rl2eSEilV/Q2Wm
N2KhMqwdow28S/ChKnU8YPu3ADdz7hgc/osWrF7UIUJ5q1CNEHJ20/s9oGiu
SSeZC+ViBRpwljY3Wog3DQIy/i94i3JNa53FFBGXcG9HZ69CoTTz62s38XxO
y5HmiHBfm3hjnqNTS9Ixjh4ZRlxvhWuifBA0pDAJ5CmwP5Jp/ty8ukJf+YaD
tdDlDrtecVRqjk0wDlvArKCtBMeIoXAofvItLcKwC300Lo6HQ1YLzfSHPs2h
8ogK7E4pvguK6R4z9SVb44oFvzo0ja/wodtfyBy4KcFjd2sVGdIYi1WzO1ST
hSiZVg8D2tQEEXi4Evk62Exo/Bh6Mjj9cYoaaIzmUxElql1wJubJjZjBdGTd
T7NhsN1YU5aXJZiyvpu+uVgqIjXLR8Nxc9h5wIJaRHhFKCOg3sPoUZeSDiUE
BPVVFg4vyAeNVcDu9fsdm42t+OsiOXKeRaCU6eVf29QUP5t4lX6GbB/IA0t2
zj3xVfeIDH/4plYIr/p6F8ektXuj7tGmIvAZG5OvA6DoEsmd6vnHSQnRoXNq
FJ8WC8MwyWlKB/I5DRRgqr14BBDDdHGwdx4kEf0/Z7ND4xXNV5jUnY3LzL+Z
yysNun2aWz8HyoGKSxyIMC2y47AG7iZYbqjy3WWI51NpkgAEenxVWZZ/mSfR
o5bKnBHxZC0yX8P3jcxbKQtRjsKNvR0HsoB6JNI+StZ3gs3F2I0nA2ha9rPt
+jsrT9LwC4DuKQ0u468uMHquwnnbmkvZToWYMxLJ5sjhV1tpcsj7Zx9+/EmR
GwVFFyBexJ6KV7qkmosbkZoNd57p4sMKr+MxlKYUU8mwomS68XewxoA+KkGn
/LW5lbIqFb4nQb4H7Sbq6BNwwsZxvdKvCDXSedmQMI5gc8qxCV8kJlu9bkDY
Uqf1N+sV8igO1g8rLoWww4M9RJaWCdZ5JiplxXCmGIH/N+s8bUQrpy5XyBpQ
/FU7XrnA/tOOGrEyKITZZJEBBDVKWHhseqb6/fYGo8O28pbdh0u2kmgHuTwd
M0Mu4jZZfjElKDqbbZ+0OvKbhmBcdIZl+hgZdNpjyLuEnYyIQ8OAgGZuNZ43
0JG0+BZkb3DpguL71lVPA3v1VPEND6GlRe0ACaSC/CZvOHGYWPW6rpJWzflB
8Ezn4g/GYLUFfoEy+KiDsnHjBEGb8Xjy5x2ifretBoR24mCbywaDybP2ZfWR
BWZxqr/t4qPkRIye5RWvM9LbIBKlAWevOBz66o3FEqtVP7H2jE8aMbALgk4r
Dc8McM17HyYOw87yKTxe1ilhBky7aAb5SIrc/PTqY5X66lrDP+j10YolOH4T
+82VPCac5ggA1/py8ibMK3185JPcPGMVStBSvmBBR10h3d4sB+RsBXd4WGWz
GoTZsiRk4xoz4/aftYG+R/iiLIzAX8i1ECK0lP+YuFsVTFGMsZqjGyhg4uxZ
UnTYw+MuDqcevc6ar7oCvZaBVDiYjcn0eNBbjzk3JCmfclHu9te7lKOazM4i
nCldnmrdaagGq+jEqvhLJhpvfELaaT/xABSywVsJyyq2YpuW4QCSTRdGZ12/
VHlv6W6yNCiSnYioXA/y+pMrTizBoX/zWju9VAx3IaqJ5ZLrmspn6htGruHl
2pP4kBkuc9sE3sZeGS6p9G2UYfsl/UIdlpsae4+4Z8OLkJCHv1xCyIgLmUB6
mmRyfd+d+p40Lw4oEP4UTcNc/7jNRtPCr9l5nmxBlYjPRdK0V83MIeIG1N/i
83UbicD+vr1YoNpVZuHnnzF9cWJNKoMF+m/HOnVvn6fJ8OalFD6Sy0YXcOs0
CBXsOiEWUh+9RLpNqZ5D9/5SUnatLM2jpPdG22aXxqHP/ywz8a1B/i0lhNKH
k2nP9qBlZM0IXZgbLyfCMwQ3Ot55s1CJCvgz6e0E8eebnvWCoEMvNEuEAXVT
H+1DTyjF3QaswsrqlhmyzjHqskl5RolW04Rwbte/cMiIPKQ4v8Qj+mYcAjNv
nrVwpBY7kTlStyZLVmoc4VQW0LWU/08uhJyO61DmdQAv86qxWTqHiNk5zH+6
ZpfLiMOgRCpTf8nYOLIyBGpt895KwNeFBmQzDNytCtpTC8awLxD1bMGBqwvc
S6y7TMzMpi78o4RWVt7TFs8YDONmYlmxpPu/fL2LLlOuIqsFtX/IOPdazAUz
L5inGerdoTLhDUkda/JhGS8edIk3kNu+YrpewSZlDR3A5w1VBXua0FKEbVXI
Gj+pWK3m8aACNc4CB5plr36FWmRfb0QWw8U+sLSm/MzAt2blhKL/F4104Adv
tFcQHDwGROdPeugvi0DHgUEnSVfI7nHBn79SrULNUOlnyiCFcgkc6GU4qV8j
X5L2qRSyFPk3Nt5jM7vApWinPDiolOkTn34f1ra9F/n1oFoJEja/5Lx3KVgE
ayCUM25rorWvaOhSO8NPvEeWWI1wq2ghY+4DitfbQjYX/5iFl+bZOYJT2AqW
OPvyNZoDR+6E1ptShYWFpayMrBcBQ78AwoWG4tL75CAEMn26+CSQiXZj5/wS
qV7e7/+jox+q5PWbzPUrYarZUkFekpj9pLqpnG9aApw6hYfCU3NO8Se9MxI1
FSeV7zbGq3JF3I8m6eUhSq2LCMnDS+lu7m83jdXeTWYzi5TmgbuCyjAOgnlo
UKMmOXQunK/NXG1Mv1HXyonBiJJeBoLjyhOmpWZFSHsxYJRyzJLY33g2L7wa
5sPLjlLLakXJKL6kcg5UpRZX3jdS1MnPF2xOMkiOu2TQKNztEj1tRiWe+eSr
J/faurBQOAiX3+FLYtJ6N4PP6j+aBVgwShbLmCA69rV6ZzjoASFH71YDAB00
G3h3bfKo2rZAhZuHC77T632FBAaZtn3H/zhFvsCPWhJHqJmoyBLgo2bIw2Pr
Wi2nGppcB9o33ZBcDWIn5XTTNdnhagtm9NNKslIbAng2umykybvWMHUfpiGE
9tBJLS8g3qfLnE6JaM/FDBNFB++59UOle/szZofGwnxFK286ilhde/uiceju
6Ov+nVnHjNLULItv6y9Psnf9iA6OcYekUlsJFYamqDcPnG2Xcm7//+08i9F7
dlxLGcGChXzfRFP2xSXaZfa/8QoSK71cFMG1lqoqrUOxXTVrHUy7qCr+aYEz
SMyaHhZNF614i93dJfJaxhpPEuOB8gx1wM/Tur9lc9rZbaXpFMKis/8NbcrO
dyhNuMsd7WN7BGzIj9GShmAFL88elINeHfazku72BQ4KH34wvgiNqYzNKw2M
w53KdndZ3S39vIPyrLNsydLtbm7w5r0+VGz5zpImjQSVD8ekX9vX8thG+Czt
vkl+wsKnzp91+w8to77PEmJkyy3Ud/+axUS9aqyFBbdBWSPaU08rqn2RMETr
EuVYpIY1lUF+bwX63/Lmj7J6wETI6T69XMaZ+UyjHKR5k7aRCJo8Ka4kHBUB
c1toNwsPOaoy2SRb8E5bpgWNQf7giedfKgb8y0Djv5Z/qqB8JHy3aAqFPcBJ
1rIwSGcDoXS88a1WYV2E8ix3bFMsAwq0xwRygahnf/qJ89kuvjktoTb4Iw1A
rIFWZDZs2RtOiRucLxXSDtvKuSA9Nbs2qKzpqpbRk+CocO+JkMjox+3mBzXp
rH2kvwZG3Z+FPaTVESxlWNqE7E0IgmsbZ6R6Q2c+v7F99hCkAhVb6MZYRsQQ
q4GGB0PpNO3vzKiuXExfMGvERyd4TjCaeyCy6+t/VarxJ0LvNnwFFsm2xGBO
MpZas3rDMAQVIPpKFUu/7epNc3br5pObU6HamdO2Tdd/D/Nvtw9xD1U+HlHB
mJvyYW+tabDfGDoXVxekR683I1AN25BC4tA0A8iJJoQ6nXYtX7aaK3HcqpAc
NL1CtQ+mjDfLSjM5c0plDUqAXLUczxmlIwUKEblph/PW47Tdf9jwdZGoVl29
bk1MTAORrNPAtr+IwmlZAj1cw7BN4rXARHliB/WXoT2WhUq+NNZvCcwXD6u+
j0SePJ7zg2P0GE09sPaV1jAscgFqrg2sNGNQBH0c75eFdgtLsHeIIPQUSIgI
liRZof70uc/mUgcRqp4O7odZfBd3993b3kG6Pq1A+fuANMAYK6j87q+1yXxx
QEi0dNU/fIlKbdltGETXxEb5Suu/L+17BaFfcTTCrs4GV7iztXlE6zbDXFhm
vyuiVt8uXT/lKIrfubrpcF01aUF6/RNeDUKBRbReihl8xCEf6XOVLiio38Xa
j3GxcVse6RZjncj0+QYc86OoPCd+Wbq/RZIFbfv2vZCkT9G2AUV9r4u5eAcT
noReWfaa6qMe2T8CQFI/5IYivbmVZCcOUjXVAiOFCjLpsJy8TRq33PNJuG2I
VzZy2yqPHy4seqbLjKAgkSrDAvTXCB8rFVs7imnrX+AnXtCl1+jBcM0lqt28
eoV162/f33iTzZFsSvnMTnWlx/UQvPaqZRIbeLNECZJBRHgsfcO1/OBTqcNR
HY1HXljY4/YTUx2+LxcO6kJdr5KlCICAndj5aEKIVNt5xYaJcPpyAoJtQuSN
TjTD8mTZLHWdj7Ue/64/Sd41knV2F6/XCNxSUAiMBA4RZ3UwAsiXzPBCj06Y
K8U8txu3+B4Vkqhz/Qf0xw+DY4bFUY/AKc50ZuIPrN+s5XOM68xmSenFlbCO
ow8Gnd9FSk2kP/NtulNgFa78g1Ap4Bn9rtgHpY0wkPaHgDwRzjkdWNzIdTjn
CxwlaKO8QO0n30Hw/PEnXMs1qImDaTwglFuD9GFaAcGa9mMRQdL2YFv7lJtq
en2UPEpgGJb+itLoE+EDex8xQFOOdHyQ11Pr29/wlaPqI3wqLOkM3Q4D0aZQ
uBC1PUeQhp6iP7FzSaOYle4IDWY40BOW+OH6mYF+o+HSjnMDfOVe1wHKZJmd
cLKiq6gxQyVc+Jt9LFVP2NChqUpeWKBvgWuQmKBV+THGng9yFipCsbuKZ7Ec
8eonQpKPb1fp540gIr/dJ+fSwsH0uPd4dm9euug64WpJJPkczlPgh2Nm6NLB
x3Sj1btxEnR5ztv6VN1xyoMvMK/9LWAPbj8VKHxXgj+r3yDryL5VpDsJWaGH
d8TacDm8mo6RG6fxP6qtw0jnUWXeLjVmPbcXS5ePs12k47PmsP+Uz4ZTEy4K
wZOgTM9mbP1H7wIW1GaOCDrcGqsyDDUJhfY6S6gSu4stlHS+YL8665nMLPKf
eGlzFgqp4jIlTBt/nc5vK0bUEU7E/0W/oFJ4Ku5YqiFRTsQ8BBLNBa2ElBYb
/WAasdtanOX3SGUvYxl1wHZ+IJq2YiJF5ZILNa94RAXzrDoPQJZ3/LROTfkj
bBTFEtPH8fmo0aZi/GoggNuNf+UjwpeM85ZKas08cVy3WSGnC19dDn2ofLlq
MgyKrZ+lxE9JmCcn2uoCwHecXY8ZgIuz+PJdg7ar+iMNWhonDIITNoxGGIN6
kPxAG9XZJafpKYe+m2kyVbOdM59mp+2JSkAmgw4DnR7kGPnh7E0cHZxs5aEq
tV3FOxfnk2BVm9HUdteD5qekJeuzPj0bUjKgG7KWhdIJ2iiNL4IQcJM3KnHA
szHguACbqCDvfrX4ZXUcRvPQ6QV7oDSnrWWFhDPmulhJX4VofqUF7gr4aHZK
rUrGgSyN93bfVejDfzW+ndeZXvxc8OEiM8HzudGX5NWEShuAbGZEC+kuJ0pA
SqdOJHAPaOA27VIiZSAC0Y1t8OAnq+Zvatk75nDxenuulrxS3eViRTMgKRQZ
IO4q8fUbRST/rugaOFiEkcWJawvaSYkHICd4fSjdLuQVFn4Q4f0CVb4LD6dE
UZrjJwttQvmngKhTF7Hz5XLFS+Bx26c++RLRYhpDiI0swr1BIXg+o+I91m/1
iwF1sh3ug9DneAXtKJWUxBdAoeGt5wsa3H/5CleNEGkslB0XVRzZqoK9Q1bu
Wwdome+atDyEWiSxGovx8hRg3CmWJPSJS5xtMBehjQKmruyX5EPdqqhLOdlb
sb7nwMmQfYdVXjUjONonh5J9FQCYym2JKBVML92Y/eLu5BeS5GsDja+eOhOb
kUb0a2tJ+spbO74uJaDATVwao+DSRClAnZj6VPgJC4Y6SeNjBdtMNjrtQuxO
cfHwSzZnUZARQAynGved4FloI9vVOQhdRuPuvQuFcqhMm/chbZbX2mclbGOm
xinysV1bf7TWScNFdLMbBsqLSoTUWgcTgZY3UG9L2xuKmL5Q9dq0xANXhx4B
E+F1Q/f8FIq+4/sjPya0y/DBHvzLkXg8V7PJjcLp34DdmhU5mGl2nJlQZk3i
BITYKYa5L2FcHZW7s9sKOmzB5nLX3f8qeFKSM9lEqWdZyxauUlccblbPt8pE
zFyIFz+19lmn1E7dGOxpMgAftQUBoyST4bFuzs+Ej62Nodmof2cp+C4Ry4PI
6XwpLvcMVUBtrm+kr3ttj9Sp1xR7LWDsoizPYlSTTj+e4davt7nMvhHUVSYU
dGDEHh57NuQbApRoTTsj3aMF/cpzKLxLrRROcPK9AwlnRhSXLNqk2KEH4P1d
YORjBM5ETFK9FVRAjshZfU6i5hGY/bZFQ3k2F2c1GDE9iwfMiIjjTBxpemGZ
ybXb7rOS3LK3ocQkl3iDfe8VKurzVzwnHf0ewinE48g2AIUGrxUtPZ7AtENo
jncZgeu95K3TVy90avphtQ8waUSSyiUAArp4y+18KBeQmAgoraAdkyAdaHRK
O/FKSlouCi7SkkiG25jFQrX6++vw1CqVM8ZEl+5Mmz2C4pTYIy6+xzSkyd0N
qfR+eKyQswsryv1m1v7mbMAAIteDch9DXtu+C6wjup0LoQEtUJySvTTKyxsZ
DGPk1wrroVU6pp8r8bc/munOX5GEARva1iWeBYW89VfKTJsObCCm8tKOhdKS
GsGGUFczxZBwu86xiZF7M+AisVt1YcBc0zK/XCdQlilXuCSxF1Kv9VSY4AkE
Rti+oUzMdqe2Gf00EabRMlRNki922ucrpNFlezWCeWHVM36D2Zs5L6aNdlBV
DkJ04KfTlhMam+alZUttuIqmO3J1wss5X8lKMzE40+hyZHmesxbLkVlAOvfD
dI7tTbWhbmzwJLWXKlmb5ObiTJ4ktCuRN47VlzBnX++jTEAh2/ZGIeXNPvfk
wZL4zyv6Um24+px8pqSEdhAoU6SdWv98WIXVmv+9bAr8Y2UF/53ls19x3Xon
7kgeJtWj/3x3EjhnIxUDk84j+DvymFSz9/RmzbnoISgHT56nJlFs0pQ1YgFg
PQFZrrCzT4/1QGUQ/9WepUN9+O/FDaYtcu58F+UvODS+GL2Y9F8fiQfmG4SB
hKe/+zipzx6dJWT4hhZrXKLhUGYE7oi4feZC2MpmpoQaNN1r7E5MrUqPdVgn
wqjGMMFmMJtmD5HI6+vqpqI5sFYPWMtQ5kCK/JBURCTkDkOVHW5+8XhSP8bz
/+euy5WfE7YWitX24YYuSWPUVsCvR67683tViGaPWYaCZqEQoINKD0Hj28L7
yFDX+ZthRyhBAFm7Vb2hIJxlEvT3tYuL2GYiUgRR+r9/A9s5oze8LXAg+xNB
gh2qkOPbzMJEG5kFBy6FuNMvLTfiDvYyvZ4Y45LRXbDKtfSOYjwDYxsqkdlS
ADDwssCcoCDfftba2qVqpv1+QWufOiOzb5VGzeBh4EP7J9DkYKF8opoL7IXN
VkJrJ2EqRgK7SvHjsrtU4QD6iBcCYRE5+7r3gk+svaa2erPS6cfGglpavaUV
HanvZxUmI69wcHVgwKAbPqyrlawToEFa+d+wzkkINzapxmA/rOxco/MoyiiT
UENe+vSno1xy7AvrqPqCwhs2MKQTna7hVgHgAew0x+1s92xD9FSxCgZQrwZc
0pxGCOjAexHqR/jsQYb6KGdgfBjKmHqRfwhPIxXsZbd/0Z43nm6fXmyBGmro
rXTleT6lBQs2Fi/Zwb/EaxWmlXTKTk3sHGPts6MMlWCwExX2OjBn3JwIXSTo
RLu+Se8oQLrlOjG6Ct1ukRp94DPf7lMbwJWbYpzdWS5DPK5oGCgJbuzUGyoI
grrM8MdQLLoJU7t76YDYsAC8UVzQvYTvNrFszwda/1DR9sEW/YLrsfYqNfEi
W3X+2AXn4UNqDCZ5ixhC3OjdG3J86KOAsnT+0qF1wcrtokpt9WQsuG4Xoe5v
UCgEQFIYXSnRx7XaIS27h1GtUgDNjb5v4Rxd9PAGYG7SeRmEzWly7t4RGJ/I
mGFbF15ocP1LYq4VNKNe3fl/ld/8XFiR/fMNkLSVZRAdpUJh9JoWlqoqJzOz
i+9VcYkz8jT3XjNs5xK15aArrI+MjisrHcJ6oYL0RB6FMgyVXlpRvTZJumDf
yZHhWHeU0rAerKobhhicsWPvniqVxK3gbAJPJN/4Zc6vNZUwpZDmFR1dZJ4M
EyQJGUrJRAeGD9dEqUN58p5L0z2rXtO68DjwPzXAFVRXPhear/sHENXMTnAr
yVbdiC7zdwB5jtjuzRIq2pDLRu9qSUSRci1B3c8StFVQTH2rPtirnQ2Mm8Fa
MVe69sgZhkB2NUqYuJ/RdDBWW14tLohvDGoecrYnyjmFyLlpiDUHR2sFoGZe
ppLji2OppHoGiYxkUpSulgwFG34dc38abgDMh5VOMTbzfgKNTTQ4sBCYbvYr
nHkFfGL5hiOI1K0Fj2MuQBsrp/v4r70OJN1YVVTekllAagztNJgh08rsCeNh
qZ9DOGcN3ecw/7WKF+Es/MERZjx5tGgZ6BFtiK7XM2suD+WKvr69yVKj0lGj
/Qx12HmQjvqIs+OKWxdtQSVVFa3lJVjUOWQsDNjlShDRE+yzdskiEKZqPQrf
glijKG5yDg4jfT1BX8caLmvdklSGx64oNvWJpUuKlu0a/4TVwSA6UJnh2inc
FGA7ev3BfO3j3PocjO5UjZYXzBcGoXc2nNqE5+krrVnDWtnCcEJjeWKlRUGK
VD0B00HWmSpmxOJIDHsB4SMBVQzGZ+eJDSvhJTAS75aKL4W/o2AR9oJwdUk9
Lw2xZ+FOYPo6EvujJNROuhWx7KR+sKDP1Ps4LThKYKemax5UdfNK8SqyUIKZ
BP9PrKaaF0tsX1YjH2oPywSD0cHgKBDfxsSMFXg6Ut9fwKAFdCl+eTDgep5/
+mLbRhHVKRttL0+1innioEkfFS7fX57/7Z4L05bQaxHLQ27gnvRR1qE4edow
Hdqi16rERyiVvFyiR++JdUD6oF4BtQAXLAM5W00Hbal1/cvoiEq3UBDnQCqM
WPNGg6O4YgStsZit9tdyXFMnlA1UadD6eJE3oAJCO74h9tTk+Zv+mTVgQKL1
TJ8luK/53l86hLW9HNLUbKLNCyBZfl9R4Kqh2sGzSarpqJKrsHv9DS9WPpig
dFMFOHelvzhltpmZ1nzYy0IHx9Q6PzOacu6FGOeZXLKDVlo2vr4W9sbqJ0xs
drn9nv27ce6Dhr5HKy0MHGjEmZFlplddkcfSQaqCTwEPfoTTGk2oLj33BEx+
jw8Lp7D6vP0Pi3DV2o8n4Jgfoq4f6L4WaGoX3l5QujmSykgSv0Klu5t5F9aX
bnhnztfApvjBYYPlJzCN63JJMTsaa4zRNJa08UMb909LcA5H2v8zz9bJr8uz
wldG6/4I15udYqWX5A5rHO9JCL6LOIUOgowBk5bG8/+akJgl5ZMXtp3yDDRf
CYM7O13c3WPXZVGZx2B5rCl3qlFjFVRqCm77+v15ySSggEjyzQ6TMv4lgsVY
6jiYUyd11uQP2XblfGDTJqQtz52STmyz5gcueSd0ObKtOv8De1+YVREwLm5h
ohIk7wFZvTJIE6xqCkMVAbOop4BMqobmbYU8aS5jkKQIJFn6fz3eh3ThJtQn
RTsNVXyytL3UmztMwWJ/XVvq93NVx3Dj35T14KXFzMaO2sLx1//KxRHiac15
ymyHrsL+8ISRf82P2clZs3HkFltRmjjeNJ9fCXKd2RHLq/OGXzUmB2YMgixN
+E0URxpmKfoyhGk3Qi46rNfMh7myDB0wB2Jxe0yBIJyT9e1O45ykfGYKlrWN
Bek834Lao3hSM7rewJubni5abuZ2MRaP82kf3if1Xyqeoo32WW6UJlucQHW0
XNE6a27VYPgeqz+0Xmriq1qDDoBoc7Vgd/MXX7Qx6AnEeWqfaEwn7yEMdBuq
ALseZkk6E4NpInD4jjYC03N/6vSfMZ1B8aI5sFTpVpQ0QOVq0ywtlEfpnxVK
rPuRORAqSIvhynyrSavJhWaQivs/2Aq50fQQxx/NGmZIpUS5QB31Ew74T2yE
Info8Wvrmo1IMDRLIRTlLExCNLIbM1hXIegy5LeVuXnh4oeVycS0+vmbliT4
eWvxZjEhkI/VXh7vf+PIxYb6P4GxPeJjWknN18oTIQPaN0S5m0gfDVfMtQhe
cLSp6xC/KZ4trie8gKU+kL1x9FjuIMWM2sGXxsdWKvMoht/tRTVFejYJCJFp
FlQlRSqWYq3ChDngZ5geN/t9XhJkaGJY3dnqo5JVlwpTYtO7IUgm3fgZcuOj
yiveMiHnQzhhnGK8/pia8RKmfCs9wrq/SbpP1Tpb2MCsmJBHV+DbDttKzazG
GjGmCvRjYWwDpPBsW/nBvATOQFnHttu1RSfO1NkiDS+obBVL1nZx5kLbsr0S
CS+ft0nV6G7w+pn7cPumr/p0e5pLZbf5Rs5i7qdWAAK0rGDOfM6FFm3QT6DR
VAPQC0+60Yld/KXnFsyvuTmjgslF31lYbNvQcF36s2rA+KupkbT3JUs6yv3S
f3qEtt+5W/8xR7cnnvRnL2Bp0poDy+FgKGmrGkWjktJXWRyfrCEdktOub19s
sgT2Uwd8DqNmpTjRDWWImitW002DxmdltqKQh02VMwPctp7DblIADmWiqXVa
nX6oVibmPVwyHqdJfD1PWfdh9kdATLd6pvuCmYZI+7CouPzbStpKd+lZ4SbZ
SMJzv+gWBTb8IhFnZJXv4rgnliG80YtRUS34nvrVhAGcxH6RwoNL53XjoC8W
B1OltbLfk+eUzdVnEhohzEwf3vOQHibSDquZryLDaSqIGr7d0UIJt6pkYeoU
DX40SlXbtrxrqB/PPone2TKX8as5NQUPNdJzywpPzGMKGo1KHDMpcueuGnkn
DCk4BLonTf1qwBbRHrqXdEbrze5MZEqgTAU+gMY7i1y1yAZsDt5bksC7HRLm
UhpOUwER4QYHyI4Vt3Lf7+K8zvAvidNQTv0XArcxAgiqLBHwhUOsPeX8KPFR
hU8huLhh6pj8QGn3HGATqivaGnBzupK9ncQSuIBqRUAYYrt0okNGWiyFiXqM
GbDVZ0Kbu14BtNk4Io5Fqq0na25TeaXrRFoizzGwrH5O4A2sAAO2Xyr15O9H
qoHfYUNQz+OePW0ogMd6PqNNYtcvMiDQeBWUC4MrbuHaXJMw7VnKCfLs86y5
DawY+Syp3t1LfTDfhCRreRtVfCk5yNUXbTnd73gZaPfwK6mcMRFudtz2xtJb
LsFMACWPjxUO+b4SDzXXB0Z/qzk82zUIi00L+1Td/MqMMITn/qhsJ+GQvuSq
m7OpRY8T4lhvjmV6vrDO52S79PamX5YZjj6S974U6hLX3i5+qLbO+Fd7MdLY
oqPKYXjBqjX+4G3Zx5ktMvz35bdyrid00dnqURaXVFPKv7gvD0Ub7e/CaPB8
TOFvgzsG7qTLXfHniuNIj4GVkvqo2roNurJELYvyDXdNq8ltjONKbhMWFGX3
RPdWbYdCC28UvHDulsg1Fcmm1a4no8AGq0ET7YexNAih3iIwOiQ0SCOn3m0H
qEMv4AJJR3KV7mhrGv5JHb6/JIePmqKSDXFTdqvzuWmXddLzVjtpgHoQozUx
BI5AomblQgmBUyW8CVw/wU49uYTlgJbgbYPqqHzVKps+4uKni17JbcGMlywf
fNOZvtFV9C14Uo6GHMdFd58VL4W8PnqDB8tb0uqJhRk8OPfbc2+2K3iXFY1H
iizgQxkyhES3o4IFVRLVtjdtSUztZXAWwm91qB2Ux4mWTEYOnbzape0Enlai
hnIw2T3oNuUcGlnTQm9Fmzr5SiV26/ncQbqShm7PY58G+YCxOVb3J8CTwwvK
2ofkl8fu5R2/gSS0oIO5kE0yV4rl8o3lcHE+O7FXfmQ0+6mzRa5o5zrEajwY
5RbyEUPCA2Gpzi6RPkMqN3CHk4MYIlM5hv4I8kBRnpxfZBfbbUnz3L0BGyu0
BtljvlkeKtJNIDdBXGsgQojReo1VQOPIfnQ6AYvlbthd7xvI9LasyXDzVIOQ
6G6R6Vsda0I5yPe3i5x+58hXjFctV8z3izo4+AgGDB6z2vhGJ1MS67gwK02Q
/vOako1CgjeewAfnhlKoy4pm+oxoC1tPBkwG8SDVBQ2ocIMbf0jYD7o9AEma
oCy10Av3et7md0cvZ2y3Ej+wwaFS8VwONbtMiiiU7p1CaqbcbcbhLQh/YFlP
xbZycm0taSkuOL3zy8ozjXGrPW++PzW73/YhnCPuKSavkn/MNOxG52QbKwRI
svTRNexl8sBJiYRsrmZuIyTjDm2VwbCxZKcffzrN/6sjrLS6MyLpT2+aNuka
ZSRWY3zsWOBvJynVWKCzD1h6ulwyhHorZZqnVKQEfmC796ENUxx2xcLrIWVS
42vQTYczcqRsuxEHCO8vZ/2mwV3nQJOlZF3Uxh4c/gS3zp5a0aKpUqTRLVAL
FtnKC+EllsIbAf+MRQloF0s3Z2jK9+eQMIJfHvwd72zrXZYpOTiUqJ4NWZrl
bwJvCmnGUJ69CdZzcLjh26t4uCe5vGIThBtcfE7FkIEpmFL99B3rbnlzhlST
cj3VVMPsrb/uCT+t1Yiozf5RTjYaVN2NqO8sn2A9SsEUiwfLXRtsG7CzVr31
98NlTE/VI7CRUhTIs5tDq4dVaNEooLBXPkxw4SgBBslXeKKbpw7/zTHRD//h
KySJcE+pSaKEv2gNJ9btF9HpMjTvMlC3EvwwkzZqiePAXgRNS+ZRAmZW95Pv
Xo2X7fCxCiyQaVHvAPpjd3gjM5Hv6uxuMAebf5y7cVo8xKtHdtJU2qsXvuiE
TxA6xNMzfqf1qdBdaCgQvfA3kRrskOAIpj1GEu2mSIAZP5LvNYoGnH5/VfFX
fVEGrLL3cY+0wq/WKAfZLtiDJZpQq0EuUbnlSr+EQcBV3SD+wgDFSpmYJ6Uw
enPIEf+QdLTgt59z3zmyBswk87g46EYB0xzu4Msa5sBflPvPHpG0GmfJ58ST
vS72kjIqbtqpg1aELKef3DNU22WvTa+3F1ur+spjMvMJjgjWemM3uIuddevX
vingi8MWzNUVui6S+uiVQ+RlqR+RTs9hTqeq2XaVXqllUuqCKwB8JnvL+4tH
N5axzuRI9BYirvCnh/vGjTBvhSN94Q/f4OnIU4O9qPS5biUWS54LQ6900f/8
cKgVxprbR78S6ErwpIxjd3oJKvEqZWshmSxfb5cLgIel1fhJIPSSpD6IDnBs
b8eQQ13Ae1IC+1guoIThLvpBc215f0XTCEtfZ7qRsDUS2Nvvi8pp8FyccQ7C
5GYpuDMF8TU1nFsbEt1rle9h0aBFDL1vihpVBngNFyfaNjPSdGbZF0ZXKwYd
/itmtuhGqwT8NGOmTjBit3Y761BDBNDH5Dpo3lIhkzsFIgzySvtjwBS5vfn1
WOdH4eJRKwC51F8poXgX25P0LmrRg91lcA5cahWSX/PE79gDUjrqPtjnrTj0
wqOlWygeFvcoqM5p9+qMytw65Clna5n1wfDrrirFupNYb3HkJYzs8xHkz/QT
fOeOY6NGt3w19W+75lvV3Dhapl3oloodEf6n29UM2isTMJo0G+1Kv2QnfTJn
ugkkv2IzvXR7YrgFHf51qcxTSNpoVV6p99A5pXSiqrBehIrZlxJRoOb+oJYs
+hqBXGYH2rv9pBK5fVsQ68xeSXyP16+OYLhD/SktxK4tlUEeQCgvNIHB/lHV
JiKcH8XAeRLyZ5M8kl1D3MydJKMjkpHB2Ysunqs58fa+/Mo4KV/W1YOTKduf
3/un6e+p9I3qkZEYFjNKkl5sWtC5MTeeB3CQyxEClqgY88sSFMt/fuaqdZ6X
luENZ1BaNrX3IOFPff0uBH7OkoeItxyoPDBb8Fge8aHlbhemQmPfrObeCbK4
m/oQQtj3PxnauGo71CVGuUbDZlOquonlR5a4npUQ1ADEnXeWMDaV9YmLlrPi
j9mzQU0IZ/S6Qqcu3Atk/k0gFP+ISrZDhB7QwXhMD7Vj9SdwcpkB9yzq6NPI
6ZA5rrhAtIth+7iTQzqgohzOoRS60K3p/e5tW0LNP8008iO9NK5CrStuyULC
UAVe1Dv1kI1HrSCzcPaGlgqKj0a+WB3MwKENIt1G9TTOLPewJ+RCZQ07RzKH
5EEBydAzcG9uKb/s8Kagois7MfqKUKhe/LGPhM/Aj1GA0WSlIBHqpW4pMuio
A2R3qAmly51hG2zGtnDUPT1Ru2T+GvfHMsyIzQ+JpqI4CCF1kxRkuLc3B7Wa
nz3O5q/uQS/wjnKDGvcjja0NHDMYtBX31S4HH95PF5BpTnTaocGUQQ+pt3m+
G4bmlmx+fIVt1D5pRf81ko3AUpTOveTll2Wp6qVSSAsAdfwOaBEIu3Dk+UHH
Ysemhwmu0HPehewEoIA4tJkryc3TRFLYikAwH9d4RtSIOlhYk6Y/pnUuwLDe
fFCRwsri/2K2vpVSyzPqp5cci56Jd1wcpHMuZbKQt9nwY00MVfCwtpzecdkO
qEzswzvKsKDT3BC/I7/ZJ70rX6bJadjepvyKjXHjIvEPeQwzHGH2yW7+pxBE
p8PjLx6avXsEdjb0Xtg7bU0+in6pqwLDD1oVwxVz/Yez2ZZ1xV9JSibBS+6/
2paCb4LEhPPO5Na4i4TNIyuNdG5hqNO6oimz9mh8zibaP1lFf1HZ9pg0a0oX
8NqlYt0B1LMRT6HqXpgyRU0NQLVsdn1bGA7yRi3mHfZ46c7VVc9RhSpPKxVh
MrHnZ1v7HDXG3GBtTfmWIl5ZZSWlPOf+lZhE/eigBN8F/HKVT0AUyoR4T4i8
Sitpk3RVgfE1WrqYf1RjgrDN1/PMs4xjYKDEH1LpP6Vsw2yeOW1O7yszalcz
nKmD3i828hTbN0LZVerdRGwFboIm0Kl/852a6+FB2A6oi4Co9pf+vA7ZHtdE
COdbUiofxyd0t++c/Trwubp/MTVoYVwaQMyOtKqsdE5pzDGRIhyJFjIYpoxY
bG2Pdhmy1K/b/hCMXeD57rW8N9NpDUhLnwdWQJUZdgEiEcW5deRY+UN/aBVq
bMDuVU5K9Q3AAMmmXtmFu+OGZPPbGnZKxNOw1RHXT+HmjPEDKTz9oGF9k6pp
t3r+vk5ClCs+U4heKMyKMFd7N/McshxRGRxce0UVTzAwyerFVS7fy3oGR2KG
x5m32Pv/5OWN/Tc6WnBZbGTl4zY03X0/pRb5OUG6tBkfA+wXCJOR+N3UOlXb
jN+1GFdp1xcleB9u5n0GSgnlnNy/2CA82CzyrlqLZVdWxzNkdaowfsnC6NUL
QRV2O+T85RDmqwqXrV/h8rXN5O9SIsOI9uBvNKyy8MwAgFWkuMT6CAivJlA0
JxhDo5v467hK6DVJbDaBOWJBSnexKYF753oiItNzTs+/5HXlUIiyNbjrUMNI
GFK3aPFAzAlLgaP9gimrfnmgpBl64DY2AFQmYcVV5AvaJ21pBDu1swylElL8
ztKK7RIMu4CN3RlrMEt/viKsguTB8aqLrnIFV72/Mwz8y+vIcVRr0oFhRsyz
PMwBXa+wkWxohtRfHwryF9CMpwAeHmzE/Sbv1472gbhdlZROA2T2/IH3D50q
xqgUvrzJuYP0MlgKVbmP1a5i2eFcskqDupBAXBRTZchaP2qfYFjsf5U3XROv
k6o2MPQjMpe3LK8dxQvMmC/31BZOFCH5FcgUYx+G16hKdDdLqOR9+BTyxu4N
84nRe4ZOEqeNYTKiDX/BtlRjKhGklKzooHqRGt57cAMe6wR7rscBhkJGKLCV
PTKvq0mpvDBTTo2AQbTcnOBZ+o8HKmP2Z5319l5p1p9QEmlJcpvZVb+507Jr
3yBeB44VDlmSWltW9ybsK6eGOux7pbVVIm3v+HXm8GYEjLSbLkABiBGy/YKw
+NzwYOMCh5+Fy0vvzWJ1GKK24oX9FC/NlkmN1UVbJ0g3KAEauhzLvX+O8T+6
ygktn6fOFi6VaIUczQalQ073fHkRv9ndnplLqGq+5wfh9k0mYH2IophUnQOh
hdgHp2qthGPWHwK7wbfQGbMcdQ1vyu7z8ULbsPQtVTgw9Tx8RI09v/3nDw9a
4Fh/IMyhIXUlSc3DxhFWo3Nh1U4fFfdKYYMRMQQ+711vpd4ZBhgorbaqRzp0
z84Kht98R0pMi7t4WFDDp4nNBD1biPbUqT1QpUiz0qhdARaxdpWDPHJzHtoi
EP3X9wUfibAYyARJp2x8ZBDpFFkKrTR4NQHvNd2o9NKlqL4g54/kZayAUIKb
LRPKvFQC42uOznEwdIucz2Pg9ov05Pcsa42hEnANap1+jKrcH/HpFz+fKk+b
K1GI77qXFOKIY3aRtWtM0SqQANYvB8lqx0QfrszwxLDmLZQVctyQ8uvljT8J
ZAv9TRJfiYATKbQPdvAeJagPfmCPBHa5GCw08TTuvEHAcPEE9xUYfq777+jL
CH/S/sBeHYH1NLgHokWt/njlqcr+Hq5O3IesTPsp/9IUsF0d6iFRRuik300c
htA0t6HxVRyoRcCBT9wXomi6qpYitvZDJtli8qTMclyBSHM78se9dLaEyts2
JKvatgBZPf6I2ywoPqO9BBey8ieJV8QBECs4Mg1ks5ws0Z7npOQPZV1DBCPo
DaF9EwUIH6zOCd88P1ZyEe3ZImJOm2AelWzxXVvxMtT9/KJyN7415deGbaBJ
gqWh3gXJupEp3J4hggHd2I01dJM7reIT+ptfetlg7uYArDVY8MwOgxmCEacu
0A1DprhYUXHxGheh+D7OMIPSIFfJH9bXRskUsfVvwgVipeCJp4lGh9HrFrup
Fuo13KfGGdZA74LKtiRhofQzeiJ0V8lx3eYiDLNx+DBy0mcGGc8PYgYwhc2t
sSN9JlfNr4tOQrw4/hiHVAOsnD9IejMI9YXWFQ30ABDcku9ClKDqoSib6EKy
JOKWvZDQpLYeqyABoEEAyfdbEPj6/lvg3WrCu9ReBGxjMpr+C4UE6lykeLi2
KWr4nEi0pb8BDYtJygBJCpmTbDbuuJfoXfc+os6CyHLKYtq0bwitXy0U6Wh7
SVYYF0T2Sp7I8EFOy5I4ropf7hfj4HwnjiqzJYJSnrXnGvcehjaLXQ6uZCDF
uORMxExBbyd6WRE1ploYzHH3aL7wPM8guIMRc+S08JBHzpa+oi62NToEVCDe
z49eDOg9Iv/M+9lHygV54yR5ieZpsfLjHYkIkN5UnG7p0CA7CvSdbA+Bu+Mm
Fz0HdEUsUk2PLyapeHKyNQeiyOwZIW1o9DcBTJ0Fue7kuvJVsDhH42YW6WCe
EnXiiqVchogqgH4xEmCRdp4yIOpgRbDoeRXnNyx8iwMlyuKKHoQ7ZKZTyhim
GFAw9niaRKzt2hcv4Uf4dXjZkH9dnomUEwbIVcK6JUO8N48CPu2thyq1QIMt
GIcL2ZM5H1jLscscVQYrg+eWSuLipSrA1+UGe/U29f1f72YmHpxcVIb2zk5W
0wgIVgpjSoIVx+uy9S6ZhtG8SoQCxa3TJrbdiIH6l+L2M2YruxlBac5WB3PF
ZhpdnI0TGEnB1DBuuyPuSE5q7VufRS9nEc7YgOpcR9h5VrBSDwrqyr83XItn
WsQW0OLr4ZOO7FRlrglmNp4GpqhzCxUaDldWWTeNqYOlnJ+1VuRPv+XuJt1x
frdaWSjx90GQYQ0PEm9iu6KWNqH2/3AqDTu4pzYDLgZIO1myxlD4xeqgTB1M
odL4YWbvXYGrxdne7V87s3F+SuIwi3Y9rihgBesgeuS1hnI8qrBztr+/bLiz
ZrgSbynDShf5CjdmP2J79b9RTrWR18K6AA3/odBq0sxPqq8KX9Bcjzz0MLBk
bOLiRnd15uhZ22Ir/KloGmCq7YEQUkmrBlQ+x2687Np74CXkJDyiiPuyYHn1
rUmpjheUSffPFNu0AcW5ErOBq6LA2X/O6ngETIdhev5KOWRPQwJM+N+BG5bc
WAnYD7w17YjTuU2KXgSMFIPR2FfNspDrsl10aojTI6p7CRKTqpxstKNdFa+t
pqpDuPPmSKDqAOyDGqx7mksC1MAdBrtxEAmQ6RHNGuiyTEwXQpIIQcHOzP58
WM6Odg01AFBTq+cqThX+CZexdjSeJWFPXQ8HY0IwpYZENicZzBc3zzxBaxa7
m302JFrH3PoozRsURvJM7Cfw1h8qQf17KKEJF0PHe1D2mrKSm8nSBB2tmKRH
eOSzqSlP5KG22O3V400lVG6lbgk7nEeICsSuGoa7aZSURE/MVWOWCNgIlq1X
TUG9On1tfoA7fHMtM+XSE49JxWktifsRDhwz6064TYZCSh5MIruJB8NBvfx8
zRz7685n0388pax/DFFS36WDqz8eLWVIqNv3FhldgnkW/9cJJ/wDmoWnKP2S
pHNauyWkz7YoTzbq1+SuRgPxJ6cYy8FOaz2U5u9W54I0wg8LIaS9FXBopfMY
0GVUrmUMp4L852dAXNkHv8zLUdGF3qGEPkZ8oiha+2TDTuLqx/+xWN6ysIWZ
npimhDetTrDK9wTf/QLzr70SWfrPzLIU9Z+xWg9RK1CGK/f2LXZGZ+QOwnXI
VPXg6Olo6flepxQDrbGJmLywzxbeAg/PWXd5LONvAsMvO7QIKMIayalw9yiP
AbUtZdxn1oGur4eURkgRlZWilvoqF+JTZkBs+Bxknl1CfCT2QctxzntX2TlD
x07kdHzXkA0Bf5Nfg/rGHN8uzCYwD4tH+cBpmxSh/+BiVMVWbTu2tvGAgTa8
Q7YJfkZA4MPWYzO8flAqwrH2mIVKS8rroy2pqjcWo7n9r8Ppx44nRmTX5bIz
xaxwnhzze4nopMH1KxdnMZsiKitCI1pz9517nZi8XwnVApAdVG+Q96roQlPw
0NAIfkFpb61BQlHHpLrvj3KH/4LB6WO8644cG9KzOiyndwM4Aullwa8Jb+Yc
Q6O6WocwDD2/h+4rasjG6rIgZv97K+zA0Iuzt/T+sbkCL1m4cO8nOUjQVs8K
65MJMaAbcJxpRFJTBNMNLd3x8jBz+GCB2u3Wr5AEfawbEIsQ3AQkshlWats2
SBLgNtvDNeNGZTT5zG91wvN0CW5ZiSmKExOso8gGD1sFGR6S1Ua9HKd8dQ4U
x4PsnRl2Ktirf6uY5PrGUts0msI/mhyRnVx/uZH3wI5VNRZmB+F8bdk7hY84
d5D5Ng0PELjXG61fwyX1CEm8puaJrBEmr1INYbhaV2MMeE9Y5dc0qiVoFhf+
c+aEtxQ47A9ROqKI8tyOd0rTM6M8TewL7G4LGN8XDTQtFHYYBCPHWxUOZkPv
e8199pNc9PlDuSufL3s3Vnq0MiXDTEYFolwG2kTeROu+6EUVbWdzpyoFx9Kw
4e1u4p7b/WmIZKSwhKevXbb2a1Od9Qz2GkCdnDfCcG1aJQO/z3haStrNTEgs
bErIs8/j1wUiW56VyziKEjdwgPRxTT416VN1N1yP6TvF+STiVPy/O1vgtUPl
ITSNKV00JYxGbhZ8RgbjjG8c9MmwWS+inPGIJ0NS93x0gDh29o/43SdJdLpu
4GetuQybQ3n1UEmxiu1PXctIfwaYMMh9wNYIbUQNxBZEL2BdJOgKcBAag4Xu
V3xXYGwbrDM/56Co5vLZYTYX4for9TT/59hdY3AkzTbrLDU4ZP/i+2jJ5OTS
TFYUQrdBO/d7Mt02tYEPh55i1laV+16EXxEB0xPMl/PtTtn8n2yVRfynxjDc
AM/iUHNyp/SethiK2V2jaxH95Eco1lGxG6OFRINuQSxbRXYWMZ8AuGaB/ijL
AEXtaacA9+102oSbYYRySfYeQh8LOmMAVjHVE8xsUQISw2k7zZjae9nvi/FN
HB5hA2h3r3vJ61yL1pYMa1Y0s05gw+Hd4QXwEPYheTBuqoBytWCkLC+8hVKI
RnoPFWUg4CSQvc/n/O5bOicInL3nanK7UgIqaRNmOhWCyD6rKMOvcDelZlfe
XkAvzUKjNw/D4MMVnI4XylIxShtvAcJTKDB5idySHOmjup9AVHeBYidSpvLU
np2bimGzqIMGJX5d+gz8D8pMR7LSFzVLpBR9Ni6LD2dyaPr/4PTc0R4E6FWc
DvWbS1cOtWaBBneo5pkgHhjXakSgceN03gIoi6uERw1RE3B68Q1BznUzlRap
I4+dM6fay1ZU+eIewI8BXMwjaDw8l2hU7KWSX2XTUdcwuhBesWPSfsA1jta0
yXUudA9fOvSUAQGwJL9gsm7qKqZpYM1FVbY8dZrReThkRxEjOlc+Rt3O1cEc
vcb4hjUzC6OhoKIwuD3gLBnWX87MX6tAr+mNnrQGBIR4a6cDaoYJKC1oPw3N
K3VIQDff7lMD9zD/vlbOGK+hNc+77zYbvDu7zkjff7YL2T8nGOvAWq4bdXBy
D5OxEcQT0ZNLcyksgXLD51g8TYOo/q8S5s/f5uUAfRwCLYolPtwAeOM/alEy
BAkTGzeRE3aJVXXigBO/ULs+/+wrNEzgPSMfbhzaMTzW1mGplCd64DGflm7F
VkUfmrlgx1qJtN2IyJt10GgtFg5wT+iEKgX8wu3fqzMSX2ZeBwOUAeGJi6ys
RilUIHmMMkH58oYguVoi0Ot9FKRKMHl/biTIOfjzar4E1TOs7P8ZIeS+ZlHv
+q2nTsQxHnfdRm2XwbWX6dPg6FH+sz4kKs1+cLqhFFiQLi7coNJ2JipWA5Pk
jahD8GKxsH4WConK8SXAjn1nYnRcz+ozWn51fokqxv6BBu/JRLQz7dr8mwd7
bw0j2nisMXcOXI+ulSECO9Kep3Nbj29Mcf2sXVqa+Cuk8tNKk12JrwF4o5z5
HO9xWHge3XC/bk6YxGogyMWcY7L6j5H5C50+m/jyUV5t81/NgbMnvBebPr0h
oYsOcJVR9M6YURZ3q1f02q1dzVy4iQM49MYTNDAmZnqrT6wDaD/drFqO+nyo
qn2TFwo2nvSWpDKZWQASiYNzdLdMy5lGg+TRX/Czrtyzv3yvrCy78XeY1Ch6
c9OtQXx7RA8/dHXWc2vYSVQykaVkj0KMTKabkGh9ywjIUOSIbFVdyf5yinPV
SFiAUY4YpgPZucEG5WiV9oBjWmM5Bal+uSC7HZxWz2gR/Uc0hN06uG2sBKMo
GkBTa8nKAyTayulHeeZKjgca9IxjbxAC5K3gNhZ3C4F/r1HwzZRHonLi9ICc
Okth4DLlKSKwj1L2rWiOBLWyt92by8PCT97p3oIwWcR0YlYbknAB/TXVVKRj
Z6zrxzojUv3dS5p1czh1J95rhBqEYkhsEzjUGWU/0Uv+zJke3Fo9Jded1bpA
7BvUoMd5TyvfIcC2YMVVg+S3YMjYCytcUxJGyKnnNJvI9zsN/Oebfm78f5tX
NxC1No9FDbDX3S3q55932xz+uAK++NrM6g5Pt+dqdT9cQHwRrO8PFc9Plo2y
5RYoh5MxuZyzmmw2p/RwsinPqVX7BURHjnkWRRTM46KxpkBWi6G3Gf9B5IDR
e39UMfCp0VZQbOuc+vLuF5Iv+vOiFvpNppSpEoRbeehzY/cN979F7NQhOM8/
wzImb7tcohvV4v47zYJAOObQtdAFED/WBiM7fO8MuC80tderdorO8d8ZQZuj
KYNsOmKWHwq+oC32/6GjgwQofK7BVUMzQ2YXgs+n8AEy8kTw1E4endyt26Kd
/XEqncce3kLC61cpLAHfzWANAQus5rGIJ2G8nxv1RRFeYFdX8K5232V+UgG+
Ka0E5i5gkSAhwTpespRFOgVPwVsGiDJ+GaDAMyPcfZKWzWOJtpJdm66XJrGP
FctMan8VW6Ev54ltKF8pfQCpIOuPZQqIfgWNlG29p6htSshNe28gHtKwaQdX
cjuZd8IP40fOjLGpLgnmJHbmHm5SvZIntqEvjvDHaspaPoyhu/vIYUGMfIVm
qsF2VDIadO9k0tLwoOyBAgRFicCEU/SqagIQ+g6HPQV1MJwR6uXlPBM442fr
ADvtQfpybZRPwcocQgDO2v5KYtiuUzVJpeOhZ0dAcJNESt+q1ncgEmw+n+zz
cbCmMnfCX6YElWbzj8onLloMfyvsN7G9yza7bFTc+fnOGLj40eMJYqW8R4DZ
9o+RgZsOZ/fpVau6+M5AnsbyWxjBg7KtqeofToIJlbx3ophR6Z3QPGxp0gSU
VdWNqhjjIMHdcB2pSgNzF9I7e7pK6jfqNJkF8yLIcnv+8rcuZfs6yqfoY03w
1UnG43LqAQvEmOlfAGOdXvbhVxvVEMTBtLl0XvuiKk23/7/EhoY48dvdQejp
MnrB5UTftoEnfEnN3Wju+tYGQ7WcH63xj43FGLlSzga7UChl9UGNs7UwCkZm
SAM1SiP3pDC/XNlKkHiMLclR0FFDQORXvnNQRPFHvV7aytDJnRJZL13AWIuy
pJfUgMuPOzSHMZMiCMKaeCT/UpFWjeOKmibEMI2zPPylq/svqns6SC5AMEl2
c9zsMiArzDl44aC37TC1K/FNb6vXDyXSOhOf67DCQ/YivsU8BKz8IqUghgA8
Bj10hRfkUsprt71JfkRMnvGydP3jfZZZUO87PSgVWsbVcAn9lbmI4cf2sqxz
ktqf6ZsuPlN7QCNFo+HEA8R0gZ61a7rcP+Fqvrs8X8TB9d52cdzpACvXhzCV
61j0DDvrPd/FeRtaX+dDf3czPFlNBi2q7M6Me7pVw49PHJW/PHu/nUgZtRq2
kA34oJF006za0epNV1WX4SAevrvKkYVOVZZnhqzx9VRVK5t72pU/MEBTSk+I
FsUymy0g/2h7OjqLErOEs0KwQqdDDr6+A0diuAs1SXXpdhmypPTr3zpvVok0
qEhnkiz27TOwrX3O0GQVu9Qe2fpToBqhrWVrQ77jjZFt1+wt+YsbNKFlmGIV
opP/mem9wRMKYFfyQS4ojZrr3Y+m5u9WIMN+db4WMMzOzigksqaX5mRqmh22
NWKpBcmO+XTpMLCWrQvln/0uUZPdoS5aMuisFEPgFH58Vw/ocY0rmHc9lwFr
uVAmHYjgQ7hZu4J7bHtXHg0ek4DQ2L8euenXTvLgmeFEQkQoOkxv2b1Cpf4e
i2fpJ8GtenJR9GQ8vV6vL5eAbUxXMPlbxTRqWLhGw9hiP+zchygxssMsPDPt
4NWU83sv/0fBrP9wOFmf6bYiQvB+KKGtON6krLZf8/V8XUIhfHynOKkRnoyy
UJtdBFRaSkpS68favBfF+9rIjVKoFxPI5nElOvBHOr4Hr8lVBhBA32WPDf2s
y9AAaUJMPb+kBpi6cMsVeur8I9bUB6WzSIUt9zDexlT7RuKm8Pv1IGA7Np6J
fONoU1XPeLvxwXUEno85eTqEt/BvUvn9vggr59JWgK5FxjP1g4pA+ZEdqVVS
8PDcpIOEFXJ2QFZHORPQ7hitG0jZdB4XSXl8fGG8XdUW6n8R11OhliKxVOpH
dDt5ewmfiqLX6oVHYV4YQABauPrDviIuEvzyYRFF7xHBmAy325nAq6ra9vOs
z1z1KxxAyL3RMGAFWcyNrhMFfzvb489FjH1gmBXM8AZowgDVNvPzJeZ+bjei
xDCxdhtxgyKNwbOclfIcY1EAJrw9Q5HlQPhHX6qHmn6AJtvSyb2Hct5eymkg
3IY/VGGks/vrXV2+3kxHs0s54VrM7g1JHkYwTPhmdUJq/R42kWQJuhEYDzsT
FdweZTWwJSj7Nxb0jhoKbGp4HpPuTlOWFoMf038oyfMlTRBWufjYB0uM1CCa
zdULjT5IUUHFxoByAfmtpNrookfJ3lPs0wNkO060zfthPaxQqjXIEft/Vq3l
4WEo4r3EiUGwm32XAzGdOB1Yf3Wh2qxP/QzRKIOz33JLThtxnulUkjC7Tpr7
J6ODWTorOPNjQ6awyJ+wt12tIhV7vPECLnxE01str2iKV8EQFiLJd8i7GkGl
g6FoNhThdaJ8VLWaEkZEKsijN2rBgIAPp8MiWVhTeV10Hoh66Ua8dSnWnPep
Q9VJ1Tzd1N+3UBiUx29a3XajFdDx130tjZ6Gd/I/Jk9iiOWinULi0Xo656s6
rKCJjMXPF5GEtceQPq/NoIySecSHxdRyA9w7VGC/L0bUFfM4igy/d1NbFY/V
2bNWKDFOldQOCqyl16lZwGQPOQ/U63Lq8invvRKXScJO8RsWCdghr+5EIibj
N+d9nNgHTwtLlXu+miK38XICGi079FxuMPpAtXlAo3vfJ7Uu9sZKsuZucCHa
dj7R3VdTuJ+ujr3vHEvnOkpFFFIsKPL8p16yo2ZQ6X1ATLnoCzZUIwUpHd63
MViY4G6GitZAtlFCU+B43bJ62IhOyKHTIOMPs20ag24Xl6eOtdbZzqFdeK+6
mJ8F+EcAP7+hadnNyS9vno5qOs3NRaXyGLVIX1z+Qxi9MtM77SQS7b5F/LFM
482dlyryVotjVR1BE4AEPFrHj2v3btse4RmntuM6tFOiDyXQPvzqkb+icUur
ETT4xhwhWokFeYaAlYOgb4whRGbcMKJfWB9r8sppbJPyPSEQzF0XuhOOB8AC
5MIq/o8isbSqSQdkxg1qWH8yjDPbPnGvOLcF+9/jcGOvUZAToSZptME07qk5
EVl25eqa5J2V4c/awpPd6hjMsbIGrr4FHWOufzgpyDDuedj/fURoAfzJ0iWi
+2WLZSDz3I19O9kEvXA2aghNFB/XWBoU8pqhIkR53G0RpRyZPQz/vs7wYrID
IzhxKU4XDzsSPucyTLyD1EWzQQcHbn6giMMKgxaV2+vCIKTOcnmuuKzTM1xf
dBu3xGU/fJL3rWYGsn5t5e08NQffA7MzHTatpCm5kbFGtAFUKE3HUqbb93Mv
8IB23lW2iN27KQMheykia0M93CxNy4aiI+RwaelBghh/YBKojs5Sw6cBDitv
2AzPa6nDoSJI30Z/PCrihDCiMIkzc+J+KxHS7DFtRavuWQSlOq75Mc1x42pW
kYXRxEHOLEsnEdPlTP5W3U40dxpvSW/nyIrBMBWr6k8PcjxiQb0pUa6zZi6L
tVJje/+0Cl8XYwBiucWxVdxEy6G+fKvOSKfGdD1k14rxS46Nk00L/XqEcD7N
/u4k7KVbjaE6AU+8W+P+KcAGORG0rUkJ8GzHkgRd0MCWsu6T3Tf66d4qWfnR
zfW7y/ND+WhHmO7MqZUM9Q7s3X9jaZWEe3YHVEdAki/SZicpn8pPuEPU/vS4
5nwTPeT9DIklKbqDBL/X8CPRLo9srlYoOCgnKT4J61OAlNkrurkg7QfoIG+u
+Jeb7J583m3WDnhPUHl8yZzb49IDZTX/WqI5I7TFAwyMpqQU6m7M5n5kJxns
GBJlm04/Kwf3TLWKoDdvTpD5gkfhoQCFKtHYhPx8C3GhH347JDuEkmtCIsI8
XeGJ9tbnFYgOW0YMIO8uMROHVIi5+1mzQFafq4DAd+k1OmqaLT7Y8fkC7nOd
B0R/C7CkiUYaZkV+sOsjOArVX5Avg6e/fTgV6GA6GXK+BUeFNnnfFrCoRPKk
RmhJ5LJIeyP9UDKwCxCqAzvi4rHewHCV2XDTSpLIvJU5W4Ps15bHXG4f5hTC
S+V4ovh4VbFoYsV5GKeBVK7nMZlfcxDeuEzk1xn1IO2RpC5iBHc0WBD2Uo6f
j948NdsGvJVUH5n8gsL+i9qKumA1notK1dplm4gpFy2qC+OkX8ssShSOBwTW
YUxyxjW20cyVG2LOWt7NMTUT4PbQYEbYVOJoSr8j5PW10TKZnzuu3ehvxLNk
ZtYjPa/2ccBZM5KNbPo0j/5DVK2RmbqAOg+MPWsy00F/QjlRsgUConFCJkp/
6QXh2ga9JInm4MRICPACopCn1aFLyc8oYg12Ac0GyDgQmmx3dCtzcSQBu9cT
spZUxZL1VXsznSmaIq/qxUsA4SyyxNQNFVNfZQpFVGEfaFGfLB79HqEY6AZn
6kh8UglMgSCnpIV1rQpakLXW6OdbSEyY9xP2qd9Ga1Kz4ALlGx/enjY+obsl
cIgKze3ltuzOZiEnwdW+dbfSONCP64FXhApELCQew64NCFNyVvEESFhcE4fE
1TlE1lVP4NaK8tUEtlW3fR+C7tOZKMmsAXYSrPf0jrvIYOT2SPBACg3FnhyT
2rchft+f5nrpuJ3yrvMyrFRglWdMZyUqCVsYkVZ+pjYGJR6HpaNmibK7x24h
aTbkjBXAEknTnnomG9alAeETu8FOjoGnkoOYEHA5WQ7p8I/4M9YfyiUiSyKn
rnA5YtM/4s1nSTjcTcA6eQR8t91eusCHK4/2cQrE6tXzcli9vPRB1d8PKb3o
MfwxyKTRs9WTLfEBQO+QCgizn22Va+tb29Pv+f2bMukzS76CXMcWf/tpZ4oc
cS9M4b71OnFwVlWAzvI/GwmqLmRuhqQcR977B8PB/ALoFuykFG1PAN9cN2tw
zQqGSAUGQTwCGepnFhZ6NDpKzLZNxsZqoZcx61woEIXOfvX/7zs8CjyJKLKL
vd9oYEjypaw08zEnveO/eB9yKEPA7M1W9hipCVXfO1JwoDmJlkiFRef4QCHF
sQBNIzFRezhMc+iJ53teU+n2llG2hjOKY9XftgSZ3pfvxxf0d4r8UZ7xoEQl
k/WGw0/R9nb+4qbFnETUOEc615ESB096OYFPbyu84kr3PRvAZ81paVeIGEQU
Q+TMLP2aNlQTyq/rSmjc1ZEph8nGqIPzLUZO1tNKmB8OyIFTA+RsIPOl0ZPm
/Fp5c65/oIUHmqmXIkvXQy+t0Vl62MCMHBYyqgPudjp0VshgaNfgofsqEVzN
ANKkp4xywq744eGQYlJ1NNoYPDhzG2ddal7BTizUDHeani43MtZVeGHiu8tZ
Ar6g0R1FZekBugxjOgX6LGDEtbs7R8Q1fY97+btaDpjN4EkBNuOO+hdaCeZc
YYO0y6CK5eo4tnG8NNcmQK5uDjxrFSg701CyMh/cO1uHu4G5hPD5/aspHmVq
F6XRKAls80DtgLCYCFrKA1nWjbR4QXZ8M0z1t+ItImzNS2IpvUlX9E53a1mA
+6JPegIfgT3aWnI9FfaVnvm9dsP8EsUFhegRC6bT9f/YNH/ugH0BMo+IhVjD
0V4wwWNdLcyM2nvNArFXNibRdsBHia/drNy37cklcMvfXOCFODmBX0FFsx3D
lTFjxVG03XbplCDDIJPb9uhnrXEiluNNUr7smDApWMP4dTgkLmJNaNyfaM5h
R8vFibVivFdrwVXgLZbc77KnNGzIKd5PSnYzj+yYX/O3rDNNLH/90x7G8bHp
KaVGiDmjJvfZKj6HdUPwEmMcS6YW3qU3M3+o6SVmcZVul2GR5wsW/EIH4Elr
W2DtpDEm7A25EbzGWc6DsFz3i+/KNEippe4wExiZe7mSmLJ6g2Kgqj54rLGC
d1uBqhWXUlwHpCfTONig7F4a5kJht/JJUTiXQUCZb9nhv7B/XE1rWV2qOr4O
QoD7lTLqowmKvey8B/mZJHJl026s7fCxW7ika2VpRlPOvhdrcUI+9AMBTp6U
colBrubSRa0r6LLE7Oyl7c+qhvXNOYG4BHZ79gfF7Y+8EPD4Y/9WsDrcqtIX
UEXoWnCzdMLuvQkdbx93kXHlxYw1hWOhr5iWPud/CuYTrvELQn3KwisKagvp
OPiyq4GgiZL/XOrq8LZD9iZW/VjnvqJPHBJK7VsIgHiHD0GxMygtSl4OwHlH
J+mZtpfxVsZWN9U4KIcVOptcZEmQGeWu3Xfh8aPmb6uuOPlAO0xxH8Lg7R9j
yCuj1nMC1HByKCHSXNkJ1rk5Z6Fc04xQn8J5B1D8D8xyizcQwPBwgReZD3Kp
BKaIrvH6Uhl3UblC/7/1z+WeZosYoa9zPQDlkWbnusY6bN7xuHCZ8EN21GGt
7CUnPx4XeLFETXfgAR81Y4fGDP0BoCqssHqkX/BrKj77PcqKSxhC2fPi97NW
o/6rLxBF8ee4T0DkNcEgcT5c7w86/Lvyc9A0M2f9Nu5muEEJLvV7+K8XlX0o
JwxJSK26cJq3u0L8jFY5cYz5GtzLmDpUJQns1wO9zvJt47Vow/x/++gvWJdl
TJf2gDnipHkuT4mGj+aAUrET8NShI6bnaVJ1nrFGMn8+AfFg4iiFTz6l/hN+
TVsPWkJIgXlM1qZBf+jblAheNAfgadNu7uAKfi2U209uJFA7qTeKup5MikOG
bZd5eQS8BVCfoCKxhIOJxIx5OXtXABlTTN/XUEns5NP0S5OX/PSoKefHFhGy
unAQS4bZsvbpmjj/LtKZyIVsf1UexCeXA3JtGpYdDGJUYuRZNWZBCOAibRVW
9cwu3w1/iKop2Yk3acxfY5HZ4QOTrorCfttfq1qzNo0/FxXJKtVSTx0S1Cnr
aaO/v2DkBFC1wcLHLLzL87dAo+SqG+LN0Ar/cfjsybyUowQYLPcUCEbcaqAs
OVUzQK/T/XhW/wyqQVLJQmg2mMWgoJ27W2dCLplIB/9PCQFB/NvUP/l81Avp
pVUjdxhrVK7k6MhEzubkU+rKbdVgAVR/5RTysvXnm3e/bASvR3l7sQ4Y7Pv3
Wx/Kl+jPrAtPmL+WrlihOpK5z6yypFCFFbXeHw6yjRI51sz24cZ2uHXGdqPS
BnxxUtV/OD6W/Yab/LGcs94WHwp+EV4FGWVFDB01y9GAbZLZC7cgysWq6HXQ
sV8/agN47nNqqWJKxIBaSsEWw3DXfsHUq+y45hplhfodx6ADZMuFBUlXyZbN
N2nQq3XXTclKdLkSjLDTkolEkNBMUD47kpcmAlWm+RnFp2nzup4WaIRk67kI
yNBK/lEeFzdIi2I8TwyiWBbHYgqcze5OH2S3mR/2fMfqngi6DqUVkbR9mgLx
RCsRSscnVBpaKtDkmfBYPe4lzUoggnhnrpSf3hScl8CeW8haOQXuFnkxoJLg
UQTXnfCARmtVh3mIubyD63jLDSiBkIYWo1MtdbSt3Xmm4ngGVCghZDQrPmpB
u0V1vddHPETlJcssU2P1ffCqNKQ+P7ee8wCssWj3OeC5ZlB42zLMmv1zmFwI
3TH32WpH5YQGoinSwwVE7vKGLHky0oxfj4rHDuT881CEymrqtZmldu8+hhZj
CiyyDin2d+o8Ph4CXbIzTejCLUQJh3LVPOV2FQZkijjAC4e/bhirjjzbn1Y6
AD1JMLkncNyveKGRfwqjYggFSgEl05i+a7QcUw4WtT0dU9/KPvHr7P1YFRqK
zz9a5n6oniNi4yBgbcmWia9Ln0rjywdJrr+JDYD6a6v/7PK3IsNYkGrjQey7
9i3PEKhEbMl0j7hQ+SwRuOY1Hv29R7EFC1I8KiTeGUVqLyga/FjX0m5Nv/4j
KQfALCpLhbiDNuaAOciVEnQVQzENcu3HmgqkBms4Fxk92wdtCz9OMqClKszf
0FcA34pbywbqFIan2Y69JssVoqGUJPSIOGD/8xAHpAjnu1uK/eUOpZ4xYzgy
jt24ghugRyuVnB2PWPBDfzMCvXl/Pg3JT6AHZT9yaXqp3/xO8O63GZ36vwrr
4kWuys5xFQ0QSpRMIZ2t9Z1leMP6jWupaWdUSfst45a8U1OezVbT9RsRX+zO
Jiuu3TkDaEqmFBZOhcNTGNA/l0NWAJiTwGP0nKTS+vFcnJfjOqcEeOogR5h8
LEYGQ3Ih5LpUFj2h633WiLgVqtTi6eQRKV7PwLOLWhRb7IZc6uXAS8Ppzdy1
1w8dFdPe5ESCqg/EiZkJDSd8ZjM4bUTzfMxuO9cEwIpygmBPOUut1tI1fzkP
r9Z68+4LCO+pcM9Emx/S6ErVN9pJFi0B8kNAPtmd2KOtSSSMQwOnuC6yCw6R
Xv8TKdHLzd3PPnmX4/q+DNtCZAmiLaajpQazNQ2DE+c8CQ9YkIOnNh0vPbZg
icm4moT7m/TCRaizV9B1XSGA9g8BvPKpXzWPZPdFIaDFNG3hiYj7Y7aoDjYt
r6E+7WMTl/6sLVJLGvCPpza2gU8cDvJx0oxi8OEASRapgY4jL3TIq0i3L/hu
lnlWx16j544jCd6nrjWb53AVl+Fw/4HZfcv4d6dcnhZizTXFUEg0ggYDAzqp
TzzjFHCxABoqbG10gcyIkmPPW1zxaxDYEfolsLwNtfXpMlvpjsLk3sAu+XCQ
BsW5vOsxmxtAPrizWBV8b0GRP3BLxCQFiXz4YToJLtWh/yr2Ds/P/hSEZGZ+
IXpjTyP6cyVvT6G5UYNgBr5OOqxqTtZ83D5jX5JoV7/QMTIhEVtR0UJlud2X
Z3DcXPHdsn7V3RezizFVKw/DNifpkiRYp4x5BmUtSrYtksTrKdYVcjQ9kRVo
dmoaivOxP8hzobRAVdNUagHcHIxH1Ar3LIfJO6xtVGp6Am9aLtBsnXRVU6ax
ZzNaHJnFWG44PFZjY3Wzd5N9ScxQjZQJuZd+/7EiP8xVrdfKhbtLj1d+zNy0
YRivnUVebTKYbjClq9+2pye0sZL5xeUOoA528rGRDfIRd2SWhftIcrqJiBTE
IP3eCeA/yHE0MWPETqTrkVIfH53MiRSqjaqLLdwSOtmsgvUbKyaC7iHTvawZ
f9gWKVRXRc7LhyMEhmzXxLEWrqnCEHMfIxoDpWW1HhHDYojJm0iW6+47Hj+t
uPqpvyPi1bY+HKXsTzvw8kBRO+feS/3/LP+RKz9M4R8HBL026tGDLxoto5eL
gBkxwWwtKPLti4rg9ZE1cc8HTcvBtSaRPDhgyu66NkHf6SJV3Pcl3ABncXg8
oCD0hikrUR4xscttli8ctvkvS1QHjNvHlzWsAdJjHFIrlVdIQWH/5N4pvjdF
Ik/rHuKefJE/GAPSJG9itBx2VtVo1AV7m5W2l4Fx9UZaAfyalyedJ/H1XtEf
JtPy/g3vYCJ847nJPbiMWBAxyP85D+vFo1hA5IecMHq/2dd2hPBeRpkpG2H0
ALCYw8R+iXkHqngegQ7Ate+iKh+QHZTiOig/j2IgrDpuSbb9Kt7MBAyr20wD
RHa/Fo2gXSjuMX4of9JRlgUmy/DkM1dsWCz4CcdusbMU2pEOriPibRcHN540
oPaWMluvd55vvDi7QOO3jhJTn+GR9I/b4/B05ttK0YOj3hotA6Ed677yzRrr
NF8cRGag783I4Ia++xPLRPVtPVXuRJqwMGGIxooYRK8IlCi5huhWNdwDSwS5
/y87/8lJkMqdTYIGRQa2QRZZimf8n4vEFfF4d8NGfJo4oU+TTUkND+vIkh/K
PwdMon8WWKm6DcuXzHvvNlnP+dkgHvCr2ou74Z0C5oGaOKz0Uxh+XHQAuErs
VE0+bf2q/NuzUz7i3q0LdU+b8OcWa5nXOXNAqTCAzDOxQs5jF+V843cAE8Rq
cJQpVM5ejD5Yne7iCCL9ocu6hre9sD/w8yZ/dFqjf4Qe+Ger6v/aVM3IOEyU
veA7iu8IfNYmdfjoEkPyyhlVgkqi+L3xKXARPXxFvZjQbfOc+IesdusrX2xm
XO/krKYJZZ/RmGo2CQO+AI5EcAOyeFR06j/Pn6UQBjz2ACyqqw+3AZEb0sjE
hRrf8SYRCUCVUjxkWSLfmg36xFUaXVlxlns0PQ/ANZmogXPcbs02nBFfHRfk
KkJdE8DXSrDsMh4l/DAvkAwF1Q2mJPoOwz8oaf1aIpL0rpfXTMo2EVMD6b8r
4WTQeTTfKwRe10S7NV733zlaspxNWzUGfmIl8S9+CvFDDHiHAU6OkZad1QU6
kBDSOOO9abgOSAXcSTQrwVipE1NabvVc+4K8OqQ7OjEMrMxzgV5o9owHdWsM
comDW0S3S0xa7Yc4lYNKn4RdmoLsHK1RtOdlGMqUfH09eg+jiC24O3X2h7Mq
Rb3SYuWEMA+rdiL6d6Bgf9doQuV85/eqABjorWQDAQo9C6T//r/M9giAC1Pd
HSlhewHD4YmfV0xA33N8XZJyjCA1AZroonzqi6ZoPrZBiqbrdpTod+FZXtjO
ZJ8J9j3HgsDTyeiYV4D5Ej8tHoUaGdb/AHDKAmElqoLyonWkC10ofrFAxXJN
m40dEQ6xGJKDI2o9gfg6mlrJ+GW1dVDFQ/crnybbpdBgdUv2+TgwFtD5I9bW
SL3C+KLZiD3PCB7bkzzxJiJPEwsEu7fFQH06IVS8LMMBHA4i296UnWf5k9r9
NjNzYBfXIoUyGQVad6WZCFV/6H6t4wFkxHPd5XpKUNKZ4t0HxoUjIFPyBMSo
0BM1G/cRtFRtf199ptTuzyJ4Wky9qBS8Trc3J/yFl4EsRi+0E/JMTg4XQLIR
f3Vmj/MSaFqbPrXwWkkUAa8zPMRY2yhH8z4Xio0UU5/PKTeOtOSfXlBiE+cz
Se7LwKRJCrWmJca/r2zYBfKdYTlzdYvR+ZxOTjXaMqvVay2Yd1A60rpn4PnB
xAD0spZTNMmRnqKF3NrTnroYW6ZgrWylY/qeVAzNqhsQVbfylc5lMZS08O5D
8cnk0AGi41QuMQODZotQrcjFtQWgn7szkVbcPCu6iOykym6aSipouHlY4isl
hYi9acMZ4pLoFb1rpktJmrpZqeEf4enwdJmK4P1IjkzeYda3VQJ/vENEvAYb
/jf2gQQ51Z151I1kdJCwzTgcm3VVTUow4+cEFULCz2m0zov61wx2x/l+VApK
jDMyeHguwOnGfBaCfNwg4zHYFidJmAMGa9Hv1aAe8uZwrJbZGy2Pgr0kOg1Y
z95ny1q7TceorjW0jIAeXH/EZbAvnhAaW/ILTeDYA8hKh8t6sdZo5S+Q7su0
rPkwL19SEh88U2Vp1Mmm1xEY/sVvYuCuJSS9FIYggEuBqGolJ1Ujxdi6DAL9
yuB4C3FFICUMv4Orw+LYVoxHcm9a26qF7DXI9czOpxSXDkXwnEsmRto6ZZs5
oHl5ncsvMcDmnE10/jvTg6wA3FYvSmvsWrdhHuqGvIvLfjYqFV1WhwxoQ2Os
6fhFgZ2cuZidbDj0nWvuO0zQ0DFSPB1irg3NIJl723GP+hE1TMQCo22UbPzX
bE5HrxU4hNROWpzIveJ05WBCt03AaX+ujEqaw9rhFqtE7FgolF52sSeUUwUO
NArSsqtvpk07L+LcXQx2IF1jhj2RYhtqCSZvn4L3+GAelNR7Mm3qsiodS+Jm
8WDMwpPDKiIR1Xr4bFM6lhg/IjC01gP6+XXKz5QaW12NNlqsUxZ/JrOJu34H
2QIEZpM1a/VuM5vJB16vBqpmfPJY8AMWm8wgyZgdaS1HjIVojqxgmeLRLKWz
E2vT8hUKwJfYP2OxZ49U+nvhbFftZl2nc6nbsQ8PcIkAV3NmX1skVaZIJNf1
6kWyeqcAyz7iE7NCehORNrpYjNSrYU+sdXBg49M9pjjoPjJ911hw1gKQSCvA
avgrEKjE0zUWSRvGeH4YPuqnGHI5pbg9WzMCOj1FFlptx39WjwljhZU/oVGL
h/M6woyZUiq/WrnJN1cjUlYTuEqFh+g7TWomE68Mfxsq/oB92KMedsoz4yFc
JqPK1Z/9bQ0/UBBb98jPRaqSzeQLHXk8YfxOLpweALCWLUPzPzwN1MolK0Qc
jA+X2ooyBk0TpUllRlQz3vpVkWG0DUWR6mG2dbIFQDilhePisuNKEr3omXV1
rEOi5MjChBy3YPucrwBjHiOYhpj2dEtV7YOmXT9uPvlzqaVXgzXnv/tl44ob
EL7yfBGqejzU5WkNc8TxnLBoDD5FYXt2WLdDTW8mybOfyN/F7D3JhLD10H4+
E/6y2Z8ca1e1RCuc7zhpPnuknbtp7ZB2hYHXG74fVKwoHShLcuFHlPggOICx
t10DAlMWURAeGueYNCiPE04gi/6qiADvs7ggW9+T0sGb1p4wsKG8xjV0q34d
qHqOi3pMYPXn9oSiwHyWKKHp2ndz1OOoFW/lde5owALJVKR2PsEJWUi5ZKcP
xXOsMWCyrK5M9bkW7i/a/biCNKv8XChdb7TqWehNw8JltbR/0TwZ+DSp72dZ
ud1nhnQOJXQXta+39vuBbD1ySv0ttBdUvcbtFX2CzaclVrQGytETL/rk8Jlc
7fLF2SoEMRoA6Jo4wRTzFikIcoDjtm+7TdJ6lpmftOU0e1DNBfoUouZxYdMT
x2Ul5yjXhxP2s+HW5ZZsLdk+dEh7kZAFQPYytMLgrKmCt395+dsjlawDq+kU
IolMLtsz7nhCfQqQzhXh6kjcjezINE+WMIHNeP+vCmhhxx5PlJM8HpCWnqju
rT9C+P3bpGwSWlNxZHetnGDo5ELpOhAISDNTFCvzxVJQS8QJDbtvl3QdT2P8
Q/OFsNfY08O2WTHosFYXHf8LEQ9DbNmL2sw+Um7K0hJj77sVnKw8xYNZN/ca
oEXj5DqgGTBpmqmoa37PBFgMPQJK3STISNCa9LmR+FDFPLizOiLAIz4LRn+n
1IQQidSAK9T4r8HWNGNNS2o1tGVWupsbvATGOSwC1wdLGnv+klk1NQ6h2DLj
Zn6Nj0bnotSmeIV4MNjp+OYZenXg4p5TUmq5IMUHaZUGHosEvPMlVYJI1J/Q
chL2oe0N9/lY1VSaStXzKEwEV+1J1cCRKx4CIgrODoT76fQ5AN6QeyWhJDAJ
ngDhZMAGcViyFm7C8ZjpH57BZ0R0F/lgITKujTmfUIraf3Gfmscz51HHc1In
nTHR+JoC0LdNLCZdkAEybgFkQ3sms5LmL/MIa3IfSId08PrFG4KRLR7ietvf
6rS/pNTlNqn7uaG53+FTSpefYhrcSVhW+CV08D/kSxdxVV8Nimn1/kibjHWG
2vKidXqMvHrVmYwhmPM/kpU5zahRzln2IefQ4pFTrs26Zx/Ghxiw9CgAUwFE
+TffYiNhzbKNgyz7hlCuUO/jx2Bu2oGggQdQyXisigxFnCe+2gvNeGSNZzfR
lQRlVvVgJwQXzrrHN9nCPMOtYj5wazVYCU4fBSgExXfS9cEmB9IV4sAMDr+S
QjoVWH93IiZRhaUnqLwyoOlwJK1jNSFQnQBR/DBE4pjkjQ5T8xO3KUvPXQ65
AtTYzqL6O/ds7aLzXHI2kq5zuD8TfGj0FhYCXH+77Sv22wghjG8Mo2gkhmOg
/8RCYYy8u331wrxMTiZcRWd6dckcrxzdcXLtGJc3PcOH24LgwNAgG+VKXA/9
OY5pFgmrcsBY/HluezeMYOJaemisQQ1mBZWHq7biLY0p0nsB5ljKWRlZ4epC
7rCeX48UySKVPCH5W/TLRW+yqPDhx2MCq4GneJFXkIMY07iVeL35ojexJVjh
tsiF4l6f3JQ+DTiLAKCRhGZ7FD6Xrh9Pem2TynPHG/2zG1zqyrbTpPKVZ1TT
n6lGjPHUtLWKclbj8dC2kKsx2D3Ya/NoIKDPsuS+zMosHc8sG+UE0/BVTtHa
Kw6txoWOpQn/xuP8a+xmJ0487M2cFznH84Cyl43ghONtSmQ7niDVVL4HwfMd
4DBWu99MWNMyueVovgikQnXW6kCuRS6S8x/UqDtn4NdCEYs/bqM+BGL4MuGb
cgfSTNMou1W0WWi071yeIvNeNcfncez3KFrdTMxkwEfs9lwsakiPieba3cJQ
U1TpKXTuVhcQXtrDHocNEM/m9/IOGXrWizYaX3DO7AGzynnFBd1rtz9pMrJg
1LGgUP9Y8GJTOEDyroJIAQ1fDUzsSKWyyd1C0U7PAXDWL6DH/Q1cMnyjbFUK
0kP68S6l4sViQQZpjBi9s+CgxaFKPDLf5Fc7P+ZRasNnVaZr69LoQtCw0YHd
Y50N6eCCKhO7Q2d4CcN9Lcq8K5ss/J4kJVOvyi8Qkj0p2e51WmWd5JGgDZJr
+sUqLlDJYoJCrp4ItdjrGl4taf/iEzpbC/M4e5wR9zJix4j74e32oQ8v8X/k
CMDRqD73X5Be2QD5moiv/bkRSCLFX0YGxHF7DO6CDcOrYO8YeSxsppSfq3Am
HSKQssOOR0evpxt24T1D+X91tY2fPUFTkoOQmYOQ1fuFUDdCNI1ME5Yab/Fe
50uAROa0r3iWLaoZUk57KuYLo71rZsxwhtL7QdDExOzE1vfP0HQxUJV8bh2O
AgctTp4M6M3ppbtb41aqi7GhyBgW9fjNQDhwFy7P7WEcneEJO29WcNgJzKff
agueSDlgJ7DPTeClXKqXvxNg69ARB23rXQbLzc14MQPsWs/qqvDQrGwl8Rx9
3kxTWzkG0c2FVKwQVxRtSI5HrNQpdu7M5xR/anQhLREodHT8UKzxUjEhU4mR
guD6SV/CZk0JbCQaJPUHK6+/k7M6s19ShbQWfjZjSLZlYfHOgsOcFLdwzXHl
W249+zT1aMMQqXfqu4Iu0zSCTNzE9YeZN93HCJ3NaZ0EII/joncimF2BSgta
nt4C4lZc8QQI8qmAWbjXr+oSd3txuLv4SJEcXuETMjoiWbGOJpJOeM4giTz4
INHGaNKZLy+t9x3THucxpuEZ8KgEaPWqp8uy9jq+g1Fg4DXhsQxXhRRAYlsH
RUWoUgtWlmSITDd8LF3feFOv+IcFO6ceZC6lui9M6w2TywnI30ldb2fQRc5F
FZ7dDWjyhJQTXj0QKLmhOcezod3DSSYThl6NJxBzOxDFUfHJPMzEZFKmxm/2
EpewNPFU8lkPGunPgbsEmlpjZQWVDDBA9l0XBq21kOvCroLk66N8UKA8HEsa
okrCRDH0AyVdGTAVYahtlLW/+1Egzm+Z3xzNhqSkNm/L16w6lY6V8b4YvCnB
NBA9TRRqQiNSPZ28KR61ZQW0E/Gv44/79KHK9q7zZeoIfzlkmQvVVSXK8+qJ
XGNVx4daotwpM2eCQrMEcRC744pGkzPRMd14MwABRiGLaPnhYEAY2K2HuLvN
utJ/sPa2jV305LatXPe8rwqu95ZVsYxO6xc5ZrgwoUsBYTyogOn3FXcq6BCO
z60KtaetOETKKECGCrUScBgOOKbBACqPAzqAUsRglDPtkAlNfJwY15Etqi7M
xRILmD+sFBeWX4K2Vi2YIdtAQ8jcqawH8qqAd527gbSAQT/8AWQP7ujrpNBy
sStY+aW9dEb6QshW5Mv6ejbNJ0bzClBxblD1wxjMbCcK0JZlPVZnsVTovD9C
+p0nTMVXjkBwijVLzy1+0HRnhfB0y7Jkak5lBvGDnNoRataHa6IMfmlIsFI0
O/21ZwATNYSlTaDe4F4sra7Cuy48SZtwI2GIH+kb9luaPmRZONsRttq3oTUy
YLF3zPr+cFvd/xoM8GloHL2pnJYUjJw2d1Ri+gQrQ3T9H7MFb9HotI5CFzfC
TOCEXBQWdWJRUBN3YT5btqtBZyo3jgUKQMoBjil/FdsYKAUAl5HqDufSjNSh
pea8KjdS3A4p7r4UDgiuRI04piAQIH04PNRP5Hc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzeMYqgLz9/gEtRr6fo1zid4bP6zzjbdZmnrewLgWhxCSFxseUs4sZIgshs2QvQ5qEFv6m8k+wtngP9XqhG9uWiBvt1PHvQZTr5fsMuErVaNeQL6xT4U9rdI1oJtW+z1Fsb78GKnmRvV3nPPToJklcm/acEYFeqT3gcmzpa/mPgCKe5dB2q1u6vuwXFLFXZbzJM/KQUW0nnjY3U3I/b9sD1FS+v9VpILrkRC7IFrKY3UJa4xz7BB/Jbh0d58x3hsErvVqbobhw0mEF9O0ashYSCn1Om06S3F1pROx7ihtmfm797KSiilCztdRjm4d0MNyAczCiLjx+dEzQlxvMil7kHhs6QbbkuxzAGk7m/8SwYo58ft3lGK1asXQOsUfH2wEqXekp33PdRdzwh/U/yglVgg7/2f+JRS/aDWFP7ejuVB3rv377UdYZgquTCsGLxXYNVXX7CTnXwS51zDQMahVLg39K0kQGnHDVD+DDo2UoMUJ49JZfx88rvMlLckbVy6sEvQC+6vwOq9yErLBCdtRIsCUDx/62YljO5HCc8Rmj99YjqJIREKe5Ihe/HtvQ2ZZFVbq6v3npL0kQH8/grdUtz0AHG9b/Ciz21pQ6TTHKL4JeLkwKcGlpJMoCivouNQFxAsA33L5loM02a9xGz1W/ev8iUqCWqYnafFmEgd+YVkjCBzhBjcD98gm42swgLQBaTbSKMy8PkJ8AdMeQYauQ7vLzBaozUHxDN6Z29QFw/AOoiLFGk7K4Fc6cje2hP37MvputZ8rqr9UkIdc9FF5yhj"
`endif