// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yI1pOSE70Rldgx6VMbB7P2Ear9r2Ah9TDrQ6K3Pbi5XJ7kYuCDg/xVJVPrtC
uxe6LQ5iN49ppMZj/YEVjaBRPWWW1pMR9RqPz5A+F747tEdQO3DWzJGjMsrB
sEB4rbEG7WrW/9TQZmE8gJ237vT7XNxRdLEJrq7ednNlylEC0ackdSoJ4T8Y
U1OtUR8RB/BtAMdOdXlpu/W+NzLVCXRAR5SLOpD/F0yBLM2mC4lPlkay6BFo
190ZPvRYj1AdR7UEgW7a4+bISoeWviHptJ2H8+dMsbq0FWKy6QPMezAK1TXJ
pO/h5rhzyGXT7Rzz8gN/8aoPtZD0XiC+1mTzZsToYQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
om9DmyuCLXG40Ef5G62rWHb7tyv7MwTdaMZ1FAMPrORg+ub6QdMXddeBLlKO
yrEk3i13uqGlc3oOSLr5w2nXb5OpO3qPRJvb+wmKNLfJQlC6UCQCiO5RqdJx
NHkcCToFPlOMIpTVxL+vFB3Zd1S6iF1Ct3evL6qahrbCRH/yiiZ81EQxpVAH
jf0JU7bYstBBJzhYUfST2URKDfo4F30Nz7oLCG5b4mohh58+K1l2W8D9F94c
xi3zPsfbM73TYTvs9judCudtYVzxverioWBc2NidTt1qv3JkuxaoMELkMeIj
IYyWl1Xkw3fRreT0xEkarR4RpTL4bKTR72WQjVipCw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iHkJg1bmDHjZrvqG0eSknUx1FbcHQG3HRomryOZbj8jSdKu33RUcDrCze6ou
GDDJEL7h2IZqVO9d5kxqyOwP1xbQfHXTISB1ilpDMzhXv1DiO/UgC3TnDvjc
eGZAer8402ZWmB+apsn4jR7nm204APZd55etuR9QghDGbMH5asSvckPxnbKv
WlYJ/ZNTmZEDbDuMdbds1ZCoNKlHJOCLz+hropDa3FdOmIa0uO6x5eMlBioQ
iw3MLe4LHXxTcWQBpNcQRmoycGC0oN5+LXNEuLqreqQU9TK0YwZ5I3H8DH1d
Qxz34HSYZU/c0xHaw/p87/SZKd/Cd3Xad0LjmoNWEw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eR0shMe2g1qBB+nMSV0tiRc8MHk4yT3k1tdGFi65aBVxW6BmErHJ2GcsBczE
eLm1m7nQWpQvoT/H+JKW+tIZSfRzF602zzrmBZQC4Nzz9ufpmPcbajrSeGFV
3yVuaW0FKoK6Nyq6L/OKUy5fIoh+hFsK7fRTv4tBG6B5zWY8iI+U+J3cWuit
CVNSVReZOkdn2xpZEpiGxWr2lFCKJRtNNHQT5ZWg7qWCRjQLK1hN9kgkAfcs
7xKA8ILw6dkE50e0v/oRZmjo+JEimwgP/h+XHp6vK2JrcFXq++MTkiTOvPMY
WRiXmWFHuGgw+SsPavfDpn/KwWYbMq/y8gvUoZwbOw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PAAXeJH1udcouybYYNRqBvSI1zZB0V2FkPyE6kYF8oz+eJHH+oAquzQeWBbG
7VP8bB7gTxuAEnNooPkIAkFNXfQ2QzcfkcxSaY7awf+sYdTX1fSefparQ03l
vgAXKUGbI/Ix/TqWB59t6ZwwRvYTrOdTPbKaqlpQcAD7HSxJtU4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WakvKJgk5gWAvL5/7V0dlauEfm+VF8LFlmPPL0IfuHTdrpXo7eekiwJ39FZe
EUtZszRN1Saz8UuVwZ2WbMACgqRaDkbOufWQ0Gq6zN+/Ae0+e6WfJgEwywW7
DLMY7qO6waPUDrLRkf6kA/MV17nhyv5/aK40jRYO01YZR+VUT1hUukFo9Zme
R7wDljDOUQ+ZntjwVK534RY5ZjQ6Ch8qyTbRKHcvaBzTYK2j+D6SQVnLEY1j
3safI26ooFAdYZLprWVr8B1qPYXrsOieE3G9rGbobcW83shTSOJf0jg5e8Mj
yWHP5bZBaaZAjIlQoo/LqIFNvRGq/XfnwwRUG/XcWvC1W9pRcf+T+MvASR+4
S5D2aDPOlJ8y464fpo51NJYR6+TSfV9TBb/k72QpKhc7ELXv+RODXwJdCY0d
k1X/xdfu0V76/bM0hboy1Ciq+19ijvKlhW+4oVYhOydT0z4eOJsjpUPLZF8U
79MfiPzYIE096fmhKLk83fAnUIn2XkjJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gGcJgZq1Em7Ka1atjitX9pxh5aX0/CWWz019Rac3HWTkb5ofEH22JO162V/O
fsp+K+VwPLvf6Gnn+UTzbUXLlX+npY7wLHNR6dD86+wNhS2fUg0YbsrxfnQ3
9IxIC/TuuoKykRkUKathjfUrXWNaTDg+9F1VrXN2AapZfGAXPzQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bw1nQyJah8X6futwb3TjiCaw/0VAxSTRn2vz8WAZ2HqylMh90EEEFUivLKhw
7zGyBhchilEgZUUBmjVFQi8zrFsxuOOZk4JYYdIyj3StbbWDGc8x4I06uJAu
uFBJ2CF6izvdK/k3biMheXGCG26TcL+YGbAirsmS1PfQAGriiOw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10560)
`pragma protect data_block
FbMmp/v1Ah5tpRyqm+cCKRBbuxhDgIyrRO61f6VXICjUbj5E11r7nXWq0C5p
YveuVU3Lq6OFGMM1yKjAH3y5b2eEk/ER6yi96Q3I+g2fBqMxjUa40pea7WHi
lLQLBY9OrSq5bJM5OeoOCTFiEbHLdqVx/swonfJUQ6tWUt3tQ4TwvGPTCF4m
9MGk6HQoEIpGB6vePwSoKfvXMym4aMbxUwZTs6n6+Bd5DyBCdnAmfQ1dRR6G
72cFdrmFA+H637z1o/re2M6n9chTeAyytl3lgfgH2W8nKEHV3hcmyi7xwHB8
+7XoKSQUCGfYZnIyr61rG1RPYaUIdtnBPpCO0hskshGT6WEKVm2owFWKfosG
V658Msmkp78SulFFbM5KCHLdLEjdHv5YEdwF1VjiuTrAQ+l6vuM0vjhmBFGt
HQNqIWksYvSS2nglb6FkPu/1swd3B0iG5TmiA21pfIVINwdASo77BSfRfb/a
Grt4s4bs0vxqYHvnM4y9McnFS4qscjrniyPzNJGPr/BOgUlK+W56Tw4Gx0wW
qJyCCU+wk3LaxVcvlYev6DQGL7dPw9SOzeSjJbd9ZKZ1PHbJ9jPF3i5AJI12
hA9Q3LjscQ37Kj6pZrKH6Zb4uOTbrRHjDWIZdJrZh1euDzhknpdywjoE1INK
kIM0BX6XI/d36qG3TG9InK3DmZUnzW/JV9nGqcgKsXPEFAeH6XziTMOj6Lnu
eYsQaUI1NemM8ZWf0UZWA+gF0SKvEIT25tiLaZmLbXrwMzywZ5nkD6RYt8nC
zbTHd+Q+Qz1Toke/oqJZ+ChnQARHaLOunHVktFbSXi1ygk+/9eKtqL7mFVzx
FaFeA785IUBBSRAarnxpsIh4e/TA03YE4aSZtP0dSVmmiD1XXhI0KheSAcol
8tIed0U4N2GdSh/PJ3UBNMXkBokHY8GXflAU/+IU5Hw8xhH+bA7qE6Cp2uFB
8T5hBecvWVTjGFFh4Mu89PoY+Uj0JSb49SkHcr2UFLN1BRaWSLaVWIxzZgdr
Mim21SfgfErhCgcbrKxeDGlsVyJGaW/isD+plqDm71M8v0DkyInjeiLY0rRp
+fJi9IzKFaXELHlDPIX1qyddkOdyI7UCn6qKUV9DNO4k6TJ58BO5swWm5TV9
WsMW0Hte+EADTT1tVdWr8NOsuSyrY6+yPqWbEJv3SqnvkEv/zNDhdSirFvjX
40JF8I41zFcsWyIn2jMVnfbWLwRl8NnSxYfRivy01SNVJGRWNMhBU119e/Rb
nurf2AbAE2kvmJXIZhVrdRKM799jbU4Zf2zqSFtrDH4q36QVAqeLhYCqpLhi
TVKNyyEVMoV+PGzT/ROv0L1ADWFtp1B5syJgGSa54ZM63RZnj+3juh08wgRk
XTj5Q91GgZXukE3he6k7VElbAp9u6s5fQVqz2eKV+HapWJUK3MbxqhPZT0i5
KmStzdVSLEvHUO248MZJQT945LeSWeEt5xbvFRakGd7zG4uMLQ9JKgReQqnC
QLTu/XDVrv4K9Df0AuyqS0vefsnO/iTS7CcrfVMa+my8Ji3LzKo1sXFwhOhV
ABRYKZv7CYI0ioEQmjWPtXUeHr+w4KedPRHMnBUv8aIGng1wc5RnUZUWWTe5
NLQeQFeCGeMXBXfizC8x8sZeILXyRTt9i3mXwlMiysYJknX9iwZFLQHccwmd
GYyfV3he2esI7xMATW9cbH2V4RrwWfMgHuU+gwpcll3EhTyDtXViNBQbo2nO
A4Jr/MLw9DiBnNq1jRtsbSQUC2TgYde6uOXPN7nWol2UhOPYBaMxPIA+Crhf
esd0887wcT6oHOTXI+vgCHWLf7uryeoMFEQLQPDVcl6N/nI7tutNO0P/IF9+
Cp4jVNPsTZxt8SuY4qI1B3GEER8funDaGrkf24HJnIVHw9ZQYuA5Zz+yFkLi
O5Lxaosi2Nbm73N9V7V9d8BCS1Q/cl3b5fXuxRqKcmipm4G1wxPFXi/VQg/m
H/lj0taumQ0c/aYZwZsa1ub+E/lt/t6ZXI0M2imBp4+FL4GavKs0BZnIRO+v
BhmGHXL46EsNk+/M8zmvCYnD/KhoTqAJfPsZuy6SHqMKa6qBpA9qqKgTbgMQ
EBAsELCxu/ZUQW1H7BmzVRsbwqGeroJNDLZmSHIIykQE0j/tlIAFjSgaYaTo
GPtSGYp/XCABsHtdID2O/yFzy2vutlIF59XW/ZD/euOfAO+qNeAUuq5HhHGX
bYAM5Tb8dhxtXoXOKzqIbqm0tNuTs+Z3Zg7NwtJxo7JaiLYTQe0b5s/C7AZ8
4eLgqMYA8O2NZltnGDhoMyvCuOe6tq5A/DQ/Bn/UEh8jxWjwub3AwcHgiKg5
WbCcAUpn5T3POFLfs1N55dqrdeKPGbrBVfT9f0jYdTfnBf8567jN4n2m65Xl
Vxm+TZ8dzUb3KhPu0dyolTOkooygZb/LnE5tMk2ZSsOzQW00o6zI0C5wVgAO
qQW8gyG6k8Y6dWUC2ufZbiOTWB4AsZaAjFWF+rhxnoyofmx+Bp1/NSJwAuTd
I1VoMGHXC1bO5CUmYG9pf04UgU4jXehUlC2RnOvKs/VnBuRmDsdW7uIO+7jw
n+hEFLmJf+U6kWYOW+G92+plUJQnIhEPWEt1YBG1etrakE2Ol3hwO4DcQIk+
DrlXBW5UFEdQPAd9QtBW8QXc9ir+zS4yHzcVf8e1x3MveWJ3a4uO3CknBslU
faV1zagV94+Sj+X8uK1bbyCdcsS98Nu30jDp6P2gL6t4auwGZWVswjd/PZMw
GKexspaabmgVZ8XL5kmYgPmAtQex1F/9GSZ5LNTPcECIkZcJpxomqcj+gl4T
PMuajVnRWux3x7btJXfhpeIavuEqt081zAQXuYo2CUqylmh63p+HDHKW/RDm
xVM9JEspZRNv6th6nnumZOBo8aMNzGwxJqAjkyBgAS9JaywFGMgZGJQMsLh6
lzg2hEj0cIVhc4PpWp4uqH1AZVK3O81uQxPZYSVRZ5EYC52tFZiKji4NTknl
6BBTYhenPikxhC3BC8jKlWzk7Bl3G8rQMMsZH/V+0sudZnkE+DEArvVMkGyZ
mSJOP6b8Gr9GHppduDy10OaxNJBzH4op+JsCBJTnuH5ywARRJqz2bxB0LS3o
8f8A5k3PchCTQGLkumbE8f+tbWALNk/BXIaowmE4ded43KQweIgLbUmUIYHX
ICZfd2mVZCVHKhuulSm3I0zPrLVNIvew+8HEgGlJyYsFZRqmbhA3kvx6mocm
NBSYUjcJj1KVnMbe/oVW8k6XhHXujNq4+iry+sSmmHZ9+bSAJhqhiEnT3Ubg
7HeKqIAKHnA0df2rO1kzJWvrlOHoDX6s2iYyIFREJh3fqYL8YQaHVhgdFHOx
u0o/BCYkxoWuUHlBnSw4A6mDxrY3l0gjzh4QwdsFomWe+fPq9a+02NX7Xoc0
Cd5uSTiI1zuVEqUKBt8HJpzwCg0+JT8tVII/sYcKw23oaIFHO6rua5X4MppJ
HT4MF0UWvocRUf6atDh1fisud95NR+TAAptMyJ48sN4NjUqkkCE3OA+YtPNx
+kuCSSwJQWKgCIhML9OsIQdqzcViixtlMksu9qpM/OeEypklyjxuHzP2UryA
kxLEdWR0rka3wARUzvlzz0eJVde2TmossFTEcLt5CkbgE8W1a1bO1NJjt4kn
fADIWDquNRBVCBoJ/UKMrSMQnmJaMfM8ul3s8FrevCvFQJhZbazU4sWjnGMP
KE9njDe//dKNs11uZAjBIrejKEbd6n0DMomR5X8yakYfKjl9AxzAaET+hm5z
V1e27Vtdf99oATsWboddA6JKJ2I0iOjssPy2zkORjuV5yCwwGF0wL/bzFMRk
Q0Y9L2i7v1Y9WyGaXbY8jfZ4Gjsr8OiqZSmJ00xt2nE1D7a+SJv65dCGU+B6
Z7R8CUa7lV9eXPUiVmr5fzqkUZx0NCJJoNGYUQapKgB4A/qoemg8PjYib+Vq
yzYi0AzKFEpXpFLtYFPz1c3d+2XaHW1dVoOmPCKp2V1hy2Xx/bTsmIGZKzHQ
booz/wZff/boN6fNdbfcUpLP9obRT8KYYOukUg4402QeqfmKeeqrU7L8+Rv+
LMJMy74duxYTtI4OpOIUNt/2OzuXyEXPPdIhdHnoR+ROn8OKSyqxbKPW3/p9
juA6Icq2/v6YTijZXLYGvDudXN6ULMf0ILWHz9Zy/zuDiO8hlJuEscsrqEHf
O9VDgjz9jHYLRQf5X1UpfbEzy9WieSHNHnePz1g9Hzdi8UpTycGVF2uybT1E
kMDPHhgsLcqphYLmMEeVk+A7xEw3j6g1ymAP+dtoRiBQeD+Fx+MeOwPLtYh9
q9W/q3YoSWq3SkIl1oKpJZYd9P5OxMvX34OMSJCVFh9IRw2oSLDpKezXapKM
3hl7kmo8L/GfF4ocy4OxJQk2OlkKuqYSwD+P+5LRU863b8p5Z9mTIA7MSmS2
EUy7LO5rs4jLYDBAEGKOWzI7aglpzQ/hNsEdJaf2kjPFMScgTCXH2g/ep5Xu
G+fbBan58r3xG/uBj1xeSCEfgP7hhovHHEJ1PPwrmbBuM/7XIPgeBXP4Dwpd
eygyHcvOJmKUvjLIS0++TBqVqDplriq4M2cDhJWXLG7TvWZbCQod8sdbQY/j
RlE2uxFQVGoT5RK3lUjXzczTYwEUKin8HIb2hBwsaRk8eRSuVOXaS1j3kaog
T6elnfYxh+nELd+c8kGI3wBHO7jGTYAx8VceIrzptBTFT5tss5Jn/KpkNku3
160uFJDsdMybQhvvMnxn++3ZdFbZefrVbiCo83PHP//gmWT3rd5XiB/mYUKR
qwVu6Rbxy9f/a52LW3/A0/4O6ZwJtpCie9ZZOCmzmQM17lady2fjhLch4lBn
omSasC4pYbeLtYj8qh8LOh3frQWB1cwsYVyNV2ETLV0wopsqq3Wd6VO8Q0zQ
uIydjbrDDOj0BTXDovL2I8SST1atMvqBstbewWBAt82VDCmuafvBG6NOpwrD
SaTpWwjmhJideKx2efwRI5Yqc5j4B0o7jX9V6zoofsR3zzNSB7kM3bysU1fo
LrJcTUEkBP7V5ncxl4N7gm4+APBHVwsMdkSu4H+PAWC2xZ/dhaTiZkUj8uRh
0KfgtojCRvSBsemadyFFC52zef3Fw4XtvZIe5Nwr1SyNOqGjoAzIx1/G98ng
QSLKeqVzGzISB8cJPNJFiYo9xQaDarK6RNxKy+gRRKTqJE3FqdMVFiXttmnz
LR3O7HGe4jR7xgcREZYTjtKOh5mYl7Ngvi7q9pbfOVTzG31kluAy6E51adnO
SsDG0xtQEo7TuO77nga+JSjJMKFb8DxeAv5E6+mwFGlnkTAUApaRQG1zoU6q
abcEY1IVkRgbX2iMc9dmyiR/ix+r78cmSTv/KhV/JVKLHt28oZwCTaaTtMY6
7iWNxsWM1oFDveL5b22kdSGDpdmO2g2Kc35EWo332Ygim1ILcxrW/Gt0CP9D
rlZllctZQ8iStuZhQSa63z5ePoKjE12OLD15tuvnZIjqVqrb7hr4FkunHrcl
iozhkR9mGVnDCfTbBcQ3F7IQzmSqpgRs+vf4lfBd59qyyNdK1E7tfwrDDg/d
oJ9zDgPjHgrUp+DjI6zVmF/+NdHv645tyTVbt0B+K/fxA9cUT8+OmvQDpQRc
QuLjnmhJmZkKJJ60LSaIFd0eM2Kw/8/m86JdIcQUvYDj904m1fWFsUT0tFw7
mD7Ai+3YiEEJOGcKyjgo7jwkjUtCuygXSikPibbRVGJFA8cqcpHwaf1FQ8jh
Peeikjwi4ebbzuRz3yB+ofW7/CkbGXZ/bzLzESWTi6zR9v7tIbShdpZkiGlx
XdMDWN2wIIzpQ05r+8EKllGO7P9FcCvt7hqP2STil3vDj9suaynePN0c39JM
UdKnmZoozStiTmfydhRl8dWRo6b2hS/JY5m8qtm1KOqrNRxVlz9vGmfmfcGN
h8xPOHSGao4bIXFBEGGFKLtL7tq1Fsx3U7R/Pi/ltUkhHT3yT2feswrniBcV
itrEJu3OXzXCLrT3yzfXeAfpuaECvoJETumQzep4jGL4dfVOPxBDk1NdKpwS
cAu5c5xxvqJQcFxaPGWmrnkqO1NdoJgobD5/mxUnzky3mqpS1jRapsce6dMm
c3nixTCGYJASHmkxgyFjyxCDOl5+D6dPNp7v55xBYnbVies01naUMa9gH//N
BIeP2BIErI8SRQ+dmG5OHtQ8/yKPfMslgA+sFuu6dywDDQnFyFg8KCiQ8Ds3
fngVUtQYptTFMosMW2ux+OfHBXYxrxmoGDcgvQDU2qUwjxrievMTyIpjq8QY
NXS8KaVlsw7BzmK91zRpRCFdT0yhrHnUaMHrFdkSrzen26zoDAh9/jfMDO+m
oVxLE/jHwiGyaJJaVt8SBqdj4ZoU9JqeKg+ke+aApl+2a1WHWqnefx7c6NEf
sJMC9bpuR4fdZDNUuMY9rIfWGJEnQKkD4r6uvcea53E6TYrmvM4Yq2MTChRk
ddcFRBs0HyjO2jDnXG0DVW8B0ASj7Tp0N7SczIAoZCKpDUdz5VUK/sGu6iKP
2S5UKtoWPdaGsXf3MIppoJS+jgPIvx6ersDo81A1xjKtrBZXo0N/zN8fCB8U
mc/ucuuj7q76rxT6NNgp1bgkc56zWmVZ44Tw4iNeQq5xD+3X1f7EyTiZBzrV
qM6Z/RJ9xM9jvPNjl2OghvzeItSKmWou5av7fB+0eg5lxdLGiNxDZIcWx0bc
Gy4v11WPItKOaLYJtligcYNP+VnL8+RDsNuxTvGd7t75bYq5rhpZHNbvxH7Y
HYCXL/zt3bDl7c7m8tvpiNN7RoszGoe4b/huOakJcScGI9W0KUk8WTPeGMbT
dwBblXb7dM2AO9114BFA3klq2fzOPW12Lvtp6sAAtC19qDRVzX7ate1ouYJD
ffOkG01CU3JiKGcaZOssq9+SVHpmtkOEhUmU1UPdrBsYX23u4BxjvL6ho5GQ
2zIAv2brsuonS/x8OX2LIR6CzrVq217yBgJwhMh4YtiZNOOa6T89VT3+5TKV
1ePR8ixmpTjAvWRq+6eCLrZRjqBTW4V2CTrEd8C/dlJQLyI7cHRZrf4BMfx8
2nu2VxhMI0GRCmeIFPYZsWt6MIp+F1jQfmjRzQoGy8M5YY93xLRMBPlYtSeh
GBGrmPUwN3fGA/SX2e4brg6gl+VGKXA52V0LyZffcmsZvNiN23wZWnmxQbKM
r73o0w4dLidkUVQxSMvFlReBzk0wUQBYQ9tr3BmCBS9/IlbelaR7WmQ/eWbr
MAWZiZq3ysNlRUNi+emKFPu0SnnCR5eaZr+5GiR48zJZ7lWev/aIj7Ybqcrc
1bfMFryOz3I8XIHm5YND/AmY3q10jspwR838u+e7Pb7FAYKHiI1JlVE80CWg
pJZZp7sCkBKUhYcvHWxBAQdqhcFyy3bI09HPG1eOhxKDWqprBOooFkl/iaZf
TN29MAFBv5tcPrEYqjw8giHxW5ITGxC99DMEJT2R2kzzsiMJa7tS1yk+P17P
xClmuYLJuF9C3x6gcYfZ9iCDde1pLrgRX9FiI7oDbVKpTXyDokX3ih3Hl+YW
MmYk5JQakXoBFWdBU8GbDNIwTHiz8jKGRSzyfzv2cL/THV9oCvz9FNiT5Qh3
JChSh1iHBk1XZ6QhAiEctOOW48RW6vlZVtiOFCk5ynNi8L+qv3lacWYxKvK8
oLHwEc1jzBUiD/jerjbfEH08rHWbBTSlhBfKQkowE6m4Y2/Ugq5z/mdK0Fzt
EoiezHL6U3JeQiDbf/2bH+Xou2Dw+EUBtZmUzXqc5TowpqcevA5H2EN0h6Bg
zuZeEAj6qzh31hE/rav2BYkY5nccupZy3Vbc6x9fjywUba1iiix80x0s+0+6
zCcbceowIRFCSavMwVb+/f6vJ2KbTBMTkrgsd92YYObbreJTfGR8QKHhaD26
+T1g0zhi3AZRdzOjYCZYxPWqU3O3Uaq7Qv91L1mmlDfWnKgroNREdUWlO1WF
3XebKP6EWef0IYKcRnmIDuUyP2MeKJc6hZyb1bbde68DuSjQKjn7lOiSJ5Gw
kOt9JYHRewwXiW55ObQK/E+LX7S7DTHPU0STAqqGdw5UtTAux3PIQ1C+C6oT
Z59ipiMwrikgOPjH4nEt2051GDWui94ZClpLZbDGULYmqSqQ2dezNZuazaIy
fK5sEglI+j2SjTNcsz2ELQ/Mu//0GCLUps0fe3CxYrrL6+5xqmfpgagYsU9l
MC5PTdd2g6Qph9R31nfy9uhyA1SmAJ30zmLKFGC6JjwuXWqoOwKOcvpjaDai
X954rF8dPlDk7NleODRW68Vtjhqkq5mkFFmq02kjvTYwddSu2Oj6qNvqyHb7
tqGkGGhF4D91xZiXgciQMKQUt2H6RAEg2WQetxsWClco0d4LbtKhwu3MNfLi
lzPny7OXeZ2v5pW/sC4lr2ZMvlE9nS5QDS0eoRV3kY3yVJlb/Z2kRTI18maD
R6kSCnlon67n16MbAxvdXB6kIMSHNHtr5w+D+usci4WwLqJ57Hqrn7djRaAG
xbg6RY7T0kyJVDc2pReV47+o8ww1xbfKsNuVfOAW2eM2CsCxVwKhHT3xvGhE
RlgCRK5X1+XARk0r7fxRsMtt7lGd4SOT/SFI1Yz0JTnIlxFK6xneVbn0x0l5
j5UPhvSN9AqfICMwqdFqFbJ2Q2Ooc7KLOzm52Ul/SGH3LveuKMKIngQcpLnx
ut2g+HpVJjeDqIZuCkTqcusvkGaGcJGHVqOVl7PE8W6zbxCcYki/0AkJ8COB
mBECiBVnHKa5ETCT5XGeOCY/N+H9nzJpLa6TDj54Ga20mBS+TrTTeDcDBEtZ
VR9s17gufI0yCGTkon+Q3I9pVgYZvRnWhCxnTT/goC5fs0zjWWwYvKH0srZD
ZSN3islkBelfahtPnsIa0UTCV9UCVRLGXvDFfJs3LxB6qSi8PT1hfZUv1Jti
tXukNyNFhtYliaY4zcvcnmPYm1o8AIU7BRujU9P/O9Eyn6kCqJtn6UI1rbNJ
iH6maLybrMyGkwcsPcnGBxmSxVSUC2mRSP0PsjMkfG1pmOlkQ7Q5YfwbJwW7
CbY60hmL74Eo8PQ0DOU0ArwX3sLnwXLiYynUGKaTASFT+FypF4X/V88zB+ft
cl4p5Hh9kPl6dvdIHJ15AkQa18E5H4QlsfWp97CvhScBdbbxIaa6NKzToWRS
zeQQMl7beDXp77PvRHLF3nAKpKIzRWZYK/biF7vAVKk9VMNiXqr8krKkTCVu
DB/EHILDIe51+BTssiHMXqMu+gkP/taRbxbyAGR5hAohq0WlGdKmhEZbhMV4
sm0enF1PMsqKn//4gjPDqcdTn60d9jYCcMRlBm0NxH2xCR0IM9NxktPyuiwe
KoNOwsHr/qutUP26W/i6dTtJIJ3Q3CohLtBBvP3WrUtbVXwulpn5cJJT1FjC
KL7qvTBUyW1WZjZyXCIsxlg8xmkChxpd4CixHzYBDDCay4HeCj1WpFxRqfqR
o4EUASBBUM25Qqru8JGmoGtnXZg6yuzgAn2939TjYZybX3gAqFr6RPPBjNOk
jUJW8SACY+wEdejNsm1vhI/uY22Q1dshA9syh0ZZylnD1AiJFLhZ5Ehew+s5
6MamBxLC+jzeXSvJa5z3JhfTCQjbEKbAwFaH6R/exX1hRikRLu0ulxybNVqk
0bnvq8/TTHPrhyZ47HjAOzl3xCYS9cnMZMKQaV7n2JSapZzTL6oAFXi+mwE2
SodoI+4xZA4ereZ9hmFMgPB3t9QnbeESfnzcPQcKLslphfpJhbOOin8gxWaw
VD4DUHi50M9jRSz3NaC6jNhNdOAJpbI0kBhjV7rEMxUqOl15O9oKQt1wXEbD
g07hhM76lXfRIBeM7+6mIbp8nDsaR+/w0vRoD0pcMMV0uVEP/onQ47+B614e
EMfLXpHV/n61l/RdTzxDg1ft/VZ+ajxNHVd/MNGzjcExi3Gxo+vDXa6LK2MO
Rtwifvam1/xpEx1OEN520jvuFDdzlPiDxcjSnewIVBbokS/u7ByyqfSey+LX
c/8J5THOZTe9+oCzeMvworRuTgxjq2Ylc+xcVz9HDqdDTHki2hm+GGlL/vqd
jbhaTUGtxYaHqFcaOx0sQqmuk4OWIdJ2UcYTYFu21yjXlOREeEuLjz9DwRtC
IaB51DXJG3SmWLOnMsnYyD0W98a4AIhdB+rA446Fkbehho/YnXbZaHGVcNtW
z51TTsA0mKUsm78BIlH5k5cq4mJy/dHCOdAMPnhwFQ0dvqghBDktYfM6bsKk
q6SRlcZytixJJbcXITFZuFi1/KcK4CKLL0zGYBX2nQwEigYmXrTD/Qq1B5gM
HZ64l4Eye6f/KhMQKc1aGir+CkUuoImd0S+70mLLlL2QF8kGaas6o8ec/DS0
RTtwrM/93PmLOcvnSkdFU41YJTDgvNQFXQCoJupllkQMCjmXnYe0pRDkH3BY
lltosmwaZRAhsP728wNqsa18Xbdkb1VbR//svj5aOwQ0K3EfsXylpP3/Ie48
sIvSGHzdC+YUsq48VxbVukeE+tBuW8pOWC/bAUqs+7CUESqE40sVmQL2A3UK
b2OGPsi6djPpDyw4StOznnKQPSfySF6aPoI54nA5dlbyk6KqmJrV9SGWoPwd
mh1KPeDBiPt1PrAhGNlbw/TdLHKTyMohjRmA+TqFMp+G/IDsMUgVL9No6WE/
xhwBrVfK40vyTrD6zdm1oRyfgN4Sc9FV2gtQ42BWTP5sDB4K1ysIRu2zNDI1
aVR3eHoZqfFEx1Qg2QZRtxoO9qjacWM+gAC5nJ1gBo+uxbtes5CR+Zal7Vmh
9oF3bgWB+Pe6c2dRMzVbBVmELMH3iYRL6Ehs6nmioIauyoa78U7KKn6dXTEd
6bmHQr6W84FTCF/ZwfqrgH4BiFtXxorApG/lDJzdXpWGmz+vslZ6ng35rCpz
s+L4b5AVLFImPxJ8MAjSAOnvhWq6ia4xKPS7LHtDCtdL0alYh9P1Xf1ZInqp
n8HjsZkHkr/Hor1/YESZeZi3WWDqEnqLzc9ODRx4knys2StxmyDIXMWk5urt
EVHrG7yK6UlBqWwM+mQWO072g4fkj2Q5KZbbR47x7UMOYJ3x/aWZEPe6+mMY
uPzZiX/JldpQOK//xoPAAgXZYU+vTXFcHh8W1/4l2/NSOupyPKGNsWfmIsef
GC9oob7ljMD6wS0G/iHMIstaH0zxWoyCOJBiUFz/5ZbQSCO5mXDBUhhcXGyY
jNmxgj5SJF4JuuDsVY0SECJDv51CNj9QfarSB9a+JH4tqERDRBMTKbFr5zUz
d+CIYDVzI1WwrJgoMy60OP5OfBdPUlgIM7cbvs6qqkiM3mckiMBS5epSGLB/
yjluegwQKnxV88JPsNpCG1HNlnA8RjoykYp/W5g7HmADC6RFiwcXB5KQV+fd
vt+PYj8sGxMiG3k4CCjsON23TERoaxJ2y4APx5kV1KPPjlzFlcGClLyuXjt1
4Rqvdf3q131ZgP5w6Ej5+w+IhBmTUH64PlJqpdzK5U1IeVKdzQHRTQo7L7bS
GMVFI9hSI8yY4Ni7ucGhCh5ZnDuwY0pGLfMBvrFH1cKPSB16ymWs4oeCKNtA
dyNnW0js13hmxGfdWQXAisQbdQQKJ69khC64BswF1XZ87awcRYO8ZHxXKf+1
QbHDFBf0K05lc86RuFS5NaQRXuO3w96ZpeBuVqgXghZDBHdACmWzuwJ9B17A
Y1vq2cXqO4MWVPoAScV5deegjafjvNbSkGNSQHr/kcjElOZ9EUlEjlSv7wmM
BG9nF2p/rdcC0pui4CLvNGrxytj72AWshsmvy4wly7iKgOXNJn6bl8wyWd7y
2t0XvpdlWU7IBXELna3idQhClQ9zAdVsegcqtLx+T9GCKb7wph7W/THqfq9k
DGhn0Iuvy5n8uRnjCk1//SDl9do09z9O5oYWestfKJuv1QPFrtoS2CFaCKQu
IRf5TmLWFT/rWV3ednKgMCtt4JFXezXzxGeYWME41OT5eeiZ7w5BuNBXIR+i
gVdOHe5tRJvsB6tH3EFCHBkyl/jWoGJ2/J0G/hsZh33ooeD7llCYjnkbzS0g
xzCjztNXz5Y9R+NGIKSDAdK+4uA8DHXY68yvdKioi/ZEJKd93FLheP+D/uxL
L0Qug0CWB59RwnFmf063K4AEzGw0fB0PENKArmtPyMSM0miVkM32mJVpSPjX
+RGva1yaVpn8nQqKoWHb+f/Np/bpYvljWXTSZQjzAkIFFcKTBoPv8xGlaP/M
pYdVTiVl0y8EyUFyb8cat7q2Nn4aXeoAcL6/b93xlOCIq3HJDL7hZg9pn7gB
1YuLP5qaL1oDJDbGeR88CdS0ov0KIkR5q4vtwdhDj4SZQsUbM3GW0o0A/eTW
xiwZ1A89z7TRq62itu2q61zvp/3CLIvv87KyhcBhNU31dw61Hl/YEyZb7Nmo
3QTNHt0+vJnnsPWHYiHtAxVFHvSZ+qZ8QiFBsYpZI1fLfNqbTuxH6UrKoXi/
4WWe1P88+eUyzmCql3cyVtVDG4j5uWM+uYCr45C9B30Fg5ONTjS/YTC7wqsd
30wfJw4VTik81q2nvsYQFiBdYccFDQdzgS9w/2ULQMXy3KQrBQ+bq4dMJi/L
cqmON9qaPiKAOSwu4ECSEcnNYpS3ftqsncyKyU2zXcg0bjWBItUHDY0oto8f
hG1xDQweLex+LjJgVgCWdtWNknnbo+NNEy/HQenSyeDZeXbAYSS7Pn5hkZk1
m2zmor1GzKBYCQ1FNfsy3BGPmDytojzIAiY//FyCMpoGA68cdDm0SHYNKRIH
IsuCFDO5g52Kcxfa46GlBTsamEZeG+kAVnanPYhEngODnulkWic8CcBG/MAI
xmI8VHoezmTN+vC72jHoLF3Yx32T6Q14/+IozVTT3CYsKa3fpxNtDWvkTPov
pETwKB3Tq6AWLY+huBAcpYajf+PqS0ZfdVWQ7CcDE7ZR/t+Me0Lk7OOAQCmK
7USS7ewJxgMPXi/gj1xSohooQNygw1UaQVCF5Njo9/40KUEuy6jEB5mHxvRV
WjByzFHnuGgo3rKCKbIYl2jkbzRFEgJpSRLVsr3l+UO+ha+ERDi/XafUVBkW
9GTAgEVYjvBk0AyPHq8AFnHl+bQS9aWwrkmU+mR6rmzqX3eJ2lH1F7svg8Li
6UY/PXXOC4P11x8pYab5Gwtm+VZxVH+Nl88s10H/KqKxHS/PE4stBH9Z7Gzu
mYtmhBVjK9OTOHQbLwMDYAcf+gHbESSQhYzZ8KiTekzOmAR9guqKRBrEvHmG
AYAtjcHkhl+6VKPpdjkjT3eQSdRvqk+61cyyMfPBg4Lj2lwmch7JoxwHPvTk
fru0s50javiBhlK8M/B7SQq2QxUHu6scsxues7c+cnog79pk3y388Nk99nc8
/fCq2OV7KhBilhoUh3p8cdnMbluinkyA/Ms3rYJQexwfb+lWkMTaaLHgAwTz
f0QYC93WxCLtOR+sVSGdB1Pw/RmBfuewSuGxJ8o2k6mvCi++WIUPXPdrO7LI
YweM+4a2YbNVTqMjTCrZcAZk8y2qEoF1wSHq95cSMwrNfRdGlKXErGDSMCIS
pmkYxkeUEfNZML+7PU/H6y5IKSRzY+vH9b2Xnf8L0rAmZG6T1VVyHLJiHt9g
xEhC5grN+xGBFIP146J71hDtcBnbIbp0q5era2OGYz4qseD3YQLR/bP+FVva
fR4m/yDvX966zq4kaZARuwoTVx8OLC5y9uPjIihRfILl+OiX7X6FfGPNeCwX
S2es9rP6RbqcBvCZAsq17BYPUL39LRVSm1q6P7S6uPPn1jQfjDUPxx/sxL+v
9V6pcq2XEGxfWNefYXhZFPFk0amZluCR9NB36hgo6vxJsYpvWf64CV9Jah6Q
AoAInlJcWMBBXfL8Zy9YcrJkABU1G57Sfc5Gt7mwzo0m6FMQ1Y8uVcIKj4DI
fom3biY4ekjK1vLPkFcFQ7XIhGt3BEkeIf24HGdY53L1L2Fq7+4WVrFrlG9w
tE53rw1C/gIrTMH3574gJE0g33feqDYa9jFwqhuZif0UXX+MdNaRhuMvTg3W
UfskNUv1TVYArj09VL7TxnGr/bMp77qAwEckwOMS

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzeSyeEWHgbSJD/3MAo9PaEOi8DpB0eXAWL6ZflqKd1JfXq+JRCdgWCvXiGAXTEIZ66HpsBsfZ30BkesykwgbXHqhDcZfGskY1t2O/b6UlwKCYGL8537Nl3pBjC878Oas+4ODbKUSfXMXoGCRKxEDnkMrCkazFfRskEQWV5iVKaw63gCdAlarcLIALPMtnTVVRJ0mD5NMU+dAR74VKFHaIIWnFj/ElqKHb8Ud94ZqxukhkpVhVR5kdeQoCPY0hCKCB7m9hhLCTn9OGPao/hZf/dCvu/F3xq2cdK41tOFjSNUc/0vex6jL9ScNdBXQ19zcB4fu0pAAzxf+lmcj4C9X/3krpYNe0Z80tJH1NAUTt7anMDlWp0OGE4d20lqJvyzIt2IsDzgjMMH1DlmZWKLdGlBQ+lD++f/C7zOw1dlK6inOk4kBLdjJSBC6rURf5pil4tuNUuUkRkUTesVGxYe0a0u4QLTlqb7p2eqDK1Bq8+V4Zy1PnvSH7Y9WPCbAyo/RLCUIbW2Kddh1Z0R3jebygdaumt3+ZHCi/JTorTiDRzmTlviNNEOY3iBJ1ccdOwyhmGaW6LeF79sEUSrd9ywhxnTN0FaR8HdPmgbIISDsTkahzxcp80g0rhAn8aaDdNdDuMHzpsWe8Ka0dyRCpRPAaiQRlzBqZ0B4cioa+kFQQ5+0jWXy36XVQ9hfMK8qyZtTWcaT6UxdS3Mxwv5WTHhXAMN750o8RNPMTu9IfN8N+iYxLSlJo4hQLXCJ0b7Z1q/dgAhsjwsh2HLyYw/ktUXL1YW"
`endif