// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ExnqgbiEAhfing9vesgUZAdhqW6qS0CfUdE7eEm+yPzpObXbCkV5NPszmulN
nfHxoItifkzCxqxChq9TM7kW2VINnx70hj/qDjSlwO8GqUHb0S1qZ1nxULfy
8dmh37sY3dv1vuQOVPg3Q7cCysvAPPsBc1WpSoWIHiYnO7gnqBIuTOMRE7je
4fvu4E/LWcyvihmHG6gMTZalJAQeD3mclmLVP44kFiH1HW/IrLD0vlceGv4a
kw4TPZUPcF9A1rzp2oyVk7bk1Hd/+KQsQ5vHDn8r9kZl1pVlw4XR+k6pJPlE
gZPziAXg5R3qdWA3OwyavuYhgXHTsDpcJ8iw8XPRTw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m0KLpKtosW4uA9tWRrjXBdCtt0b/dzKzlkKMjQDR2TsCoWH/+zoNuOR9KyR9
VqrkVTe91Pr0cUSPbUY8rSqvQC0yVvWTe4xsZb7+j1GagmCvhY/2jBmW3tNS
Ue8fdozX4o5Nr+iiXTXo6h91JMUwFY0pSuDhmOtxCZKN5qQcMijHDJ1wKRkv
t+1+SZW1+0D+f+lCdmDq47RGRUApGEwRjsnsUJurZbDBTsrZXJ3NCuV4eE4q
HWglQzOyPPofLkx4HUlYDauQTZd4WvHnpeQMrd9TY01OJxw4Dz+uVFJMXFIW
Kprr0D8whJZ3qYl91grhINt4Kt9OtGH2WzTpAHj1ZA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KjOqjEup8w5Nm2DLhUy5CMS2W9l188F5re7DaBUgehdny7oziqiolvnhDmLY
W8yYrzgRtVi0LRlY3FNk4lgeja5g1A0e+vioAbolB5Ng6vHfPdXJ5U5shAcG
KAG1ldXeWj6pUz9yT/xM9eBds0xeODjvDG2MyySiYz/PWdS+hHgWjuLVL9Ez
rvHr3zg8mtbTiGqwTJjqey7WY1MnCNPsNZpuvJ4yEedx9a2DEM90fVcR3und
xvwPByKh1/hbTXk5Ts0+DzmbdfVmzxuwcVO5Lv+/QfgXSfxL5KTMS55XGXT1
3C3vxQ8xGyIXIytn0uiVqYpsdah8Ylf+ml4nUwSDng==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iYuMffgGNqrW8fden1UZVWCLGpsQiJGXdQLERAwuOEKE5TllBvcLuTf3i5na
laQX8R0uAqiCKyRKznw94SuDLWQqIfqMbeCEz3JI+B6CYIZepGHfDud+c/UA
VVtd9OFGcq6TnJBcTCuaGcuGctPNrAMNTEp1wIsxNfApRtTees8Ja5/jtV0f
oJiBpBZcZeZtUiv+ijgKmSg8k1uPQzULKOMCyCr4LExjPyaSgaUYXi+cxw9A
mIBlXzyvu47kkPAQTdhuyxJANz7LalNsNqG0fBsNmLubaPO+ULHM92FzIWV0
qPqplCskUeoIGf8K27gocHOvRjVF8mXz4jBozGfdaA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MYbruZNzh34P5nHryT/gj/De+iHLBg8+UN6mo2K/XKRzhhPKol0QsY3w8h7/
8DYZWBMC8jHCuwOdYGssJGP+ersCD+W9IQnfI5tLkPch2mawOigCRWt7ecWB
AfKC4ZSNfXbtksqQjxkDrh1D2neBo0VHe0H7mcxmg6csyKI2pIo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EUpXRI/sReX84RpiEi9O5i5qydb+ik93KcJUK/Vjt12SJnfGvNvxXviJX5s4
zqCuXfBGk0kj8nEO43Tbu55aHBvXcTDvj2+Fk7dFl6zNeK3pEqy9Mazt5LKs
XxsLoOqxyqAPQVZxcHWS/eWyrHVao0aQGp8+b/viN0rYL59UNjPH1McnRnRg
pjRipxtssvIUozaenmosxwnI4R73cwZ4H8q6FNa4w090PPBySLh5tZueNw9z
AHrWthVFoqAasbmd6NgbpviKIpn5s/Ch6+JAs94rgB21Un+IHqgnwyZcZmeL
6leIrGc80cH2Qwg6B4LFvnTBhg2918r5I1k6Hlw/SLMh4ftkX48YfKJ6HiUW
wFEduRBMa6bv2Nk/3n+EFKmsCX84weDAVwk8tZ0Uzn5p1pqpwawTY2uQmg35
s0uvoJWTlTFmnPS3KXcOtLQTohDPtVB4dbClnR+X5zwOVX8ink1O2BXV6yEv
xmIuaIo1BfxoV/c360adJN5/cfvew2es


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HJsC1eoj2SVSaIgISJZT8odH5KXSiRFIWyr5THbfQlDACq/T4si+ddYgNNnr
sNbJ3dZjfIjr8SvSeVVYEH9ZpiqadOa6hhpxozYBOvt4421XnG6a/0q0+XNL
qYAVkFuv2iPDpcBoXXuWyC5gSvbLccSRrPLz4hIdmEnTqMpkNZc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e4uSiBoXPv5mhha1fhy7GE6NnUvRS/a7CkSilklFpCSJEn0TyEJNcc3G4jil
ltlQuehyO5Zcv8Vb1HWvd1JuNKPQDNppDhgluI1Qn06S5De0jwOEg21aAaz+
cr3KfMowsJ6JILaiLLV6FDBlCXVdQYxG6JBakem2OeMraKK16z0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31152)
`pragma protect data_block
y5uLKkt23sOKqCKBVB+DvVR5uhY2oMxTFTwXVVJG7UvpnONZnmyvcSaWiScx
XK9jxBgnC29GQcRHttu9k0puQDdlz9JNLz+7LPiUhbGakS2NSMBb62Nlr/hY
vXCaaAsBPqxeEFAorBDHvnZiGzELHGEiNnOleyc7dQpn2/YI6H6/9glf9Lse
S986oHzk3uxSMs43otZD+hPpygoVwfxisdwf8GyogdgLmnXqbgQlbdO3EXmo
8JwwK2bw6JzpmkUlC06l9CxHSyQpmG11WZexSfdqbJLm1KgodOwaXLn86cZc
XwLGKro8ntTskOW1Bi81hPhtQ0kCqlJIqbWBaOj2NYr/3Kgf559KAS9Pog0T
tK0thC8wfiRxGtrP9bZ+ccObikrZLGTjUcGQ/3uyPCCZ7qGMyP2jFXzXfVWB
aAVmHrKyFcke0P71yp0gPwBL6zXzNoo93OzTxkCbQV7hjz4E9qlRP8SzHiqE
0i2L0LhZCKGkZFTc6AYQ1LtH9BW+5ZhUYWX5+Lxg+8o4uCKipOp+y09QUKmj
U2vgIYZBPkNVCNG5xZRiDkzBy8opBwfV3HSZZ2hGy+yQWQjS1qLC4Qg6HRK0
R243z3fxlo9tj0Op5gVC6KbRK/hQ+ozIKsuVL/YIbd6UztA9yf0Sbu2fegwm
3mDsNcRcA10txav3dYgl+4YlLHGjLjlB0N83bIoIN1WIVHzKThk29xeh2awf
jbODDehxQ2QXws/pf+w1NGoaMUJ0J+TOobZ0KCjpcF+HQkAFu4U/Ry/PXsen
KHWxDlIstQ0GiVlMmkteBMIRe+DgrGzSMwYeoRtMdZ/aKGYV8iBm5UekQaJa
09CQmPbSUFBxycQO3ET0D8rXOg3MD+j0hR6MJFL7VM5rHQVy3Zrva0YnCXhL
RI7BijTvmYRFy1Xjg3Si+QOtaTERcneKf/6Wk9AzDML+gIyoPp+lzG9zm2IZ
GWL9bo2yrReZ4QIRyC5TYRK0gT3BWLcCnX7kWt+w3yHEPj60g4I5BV9bVeeu
2A0sGZywk3fTlHCKHRexb5aCkOICXMrp9AGA7fv+ZZyBOSEYNemN9mS7fCU/
jeQG8YFwjC0vw+OPwiyMicnbQhAyBVHpLi42nA6kBo5pX9BZmDeDZEmNxVX6
WAHIZL+ZTqGt0ZJiKuGc+mambnUEXE16TZcB31eADbBTZq/VpAZUxzNi/CI/
JYcSBv/lkGyI0yrPxgA3wCDeo/0aUM50P2I7IO64GLzr6zlR4OIQaA9TbyA/
vbIKr1tY0rqsbsm22gi0+CChAlBWSQZF81EzYCpN9LJMU2hSazyAYAY/UAUw
BvcN22BsolGPkuG9C6bjoBtID77xS2pZzA5yuwMQEghJXBlFbXnh/gSWzXZS
70F+zZr7hYwcQ3Rhw7jvmL1ozw81NbBXGwwqVOsQ1JLzDyKtB85i95jV85af
lktJzB9d9C6fVlnLWLXWQ7c5toOdbPy4bV7mqjH0on4Cay5Eci8O7AAObne9
LbcE3dszsJIkzSGvj2TZk7B7ee6Glcv1bSioba8OEPfeJLotK3C1LsV8QwwJ
VAInwgwu/LqwW57WEoUWCIMjLCNP4NrM7gIMA/dZCgoEvYIM0/SyO9+6q2KT
MppnZ5iKirtdCmD1Lh84RQ+++hoSU97wzy8brB787pHqS5/W2sNlTv+iY7u4
2UqCcXAqe+gGuVwVkQUfx9SDDnYIGr1coHy37ddoMRDaW95n1WYNnQZGiyUM
Hb4m+nO3PcF49gePbbn7GtWUPy0LV+/+ihX9Jdw8FJ1i2jkdI6qkunT+PaeQ
bkK4hqHxiqY35CPap74wgXnOvInp9Nj3hit4tiHqMXGKcouUt4Wt57PWRdsD
cD+/rLvjAumFAtag+80b1PJ15LduV8tdzPgx5GsBBekiSMHqKyePvoSVKw3t
jK9yv6Xlt9R+tgQuj9Sf9E7ealosvtff8fD3JUqysbjCkV/i8GsoYYmVOSh9
CVV6wCp2Lyf66W/1HNphF/MvXvYEw0WIBAt8UovfBnP1tnyFmEGmZb3VO5xl
CkCITDsuqDJhMUkBubXvVra5ZZwxczW9D6813QWhM5QL6crSGZMMAjT78ytX
95tFcean/GxwNB3fsVfbh6tVkGYFPBNRe0gBI7LMVWkp8M+OWdySoD681iL3
w8qxC+BaSkLRWfpgmNOxg+IBFtRHl4bzA2Lsiw+rBY+R605mo0MEBaxUvWfH
6uwFLsZ310Pit41on4esZUOMZr8sVhvhH1HqFFzEHVbc64ts9BK/pBxqKOdY
rvR7Sk6xjtJPCs1XwRGpJRSJ/2y7bTqzgevBl7S7g+CCfpjKlobxYJPk9P5w
iVr8RHR8om5y7ulh8xxcJJAneU32OUhqQEes0KRkhNicE7rEgZwW4U5J7TjK
urNwBgX6MGz/F9PTHbWi+/lKQYFlKKN4pspsqYWeYl+jvh1kUDq5ExHXTqOj
icumAdBguJyi+OSSvmu7/ItdozunwSVdsl7sGgY3BeTncduqAeak+sHrNPuS
MnmLkwRpchUUmhyns3bqkWv4hTWZvLfFaFOcqD+Onhts+nXJAAyTZYT8Yzr8
xuXwkOHdZcDNbGYJePrvhgX8AIm2ku0et7fSn3vWPIo8Ul9Z4IfU7PUbbMDc
u+qvVA7PPl3t5BfJNM/fM50/lJgPabZvkI801xVDwpbCzZiN7/v2Y1zqkq+j
csP2YvYdIoU1synm5Y1KwG4VR+Gw7osOzrFF6ZmAh4Ahy3JNiK3mr1F/fiGx
dUnsWeejArBjlyMXsXnqr820HcxvMu77OpJF+9zehzOTCLamnDFr8PqX0NTQ
9NIulOef7DPYplezMODMDAFEWqmOtO4gEhBNONPtdS8w6w/063ZgzLSH3Mfa
/tC5LPUlXDh+Utq4EGCrxjUBuWrg+6nyhhPpDXEf2ZCwpaAJiDorS0WtdiLg
b63rBjO9X5xWYk1+1QbTyROAlXcbDJ5XG8n0C6wL3ETR4oX2OXcAyd4JdPFp
3oTgeRaPW3DiDEwxWFhc/t+5UeljFftaeT05I1tqtmSamZZlwy3ji8zhcUQv
o+mMqTVbRErL7Fc+6tMgTJiPy2olF0g5y/+Wgw036WvMI73neDnDaapxkKT9
7evuPCjKKChQPgoW74zE89ShgMsDr5+6R14QR5xOh5Z3p8Ad6emzlI63iw1I
7uSzZZ2JBD7eqGOpuAlZ/tdTi4JRiSphHVy2Lj7iN7a+eoiu2TGMHLzQuJ8I
2xE4zCm+aqK00jC2eqQ5VlNsiERxgirtbhmc0m9+eT/Fo9g8shfd7/A9g3Wr
spw5SJwDvP548cUz4T0SkHNO/nRVnGhI7k0A0rdyW4RL8RpA1pKvXBkVEcBL
ufU3SR7EDlX/3/04OitYc2pkUptipbD0lxtHEzqC916RTFuxfwL9Fvq6DxTF
RwbyO49zsy/9el9qJOY0A+5VFXjz5R/89I49tG3Kxw+klv02n8V7MHHuM18N
jVwVN7Je6QiI7NiiEGc2y1uZ/fUodaHq1xSE3OmZzGzVMVfWrjVXg09kSaex
h7gY0aX8NcNR6VPS6EQl5GuZlu+AOcL7ClYpESdVA9eoRALVrUtz09d1W0LW
VujNjpnhu7z7E8k2lsFB7UHaI3ZOsAdOC1SYClbSS/omMnxbjU6BULgOG/Ya
P7OFDwvwcSVAwhEwHo1A6n56ao2x8z8bkhuK7ajAf+gQFcC0mycSbJwRar3n
Mt874BShvCCfQ8PupX0Ssuf0e1m4+ee+VUkQQ94nXEVS2vpFxALuWsARV/nx
Riwx6hguB7gclhbQUYJqzPOdRLffTkg3gKWiICbCYLtupB/S5evNo1Yu18vk
+0l3Z/98YtM7gbE6cz8DKOA1kgvdTTOPwNu1Vi+K0TVKl7Ec7+MjNy0Zir6+
m1swMxmX8GkC4tpkzWKkTcEE0X2terYlM0SumPf6R9E17Lw3MIWWONl8Tdtz
JVLM8TeN5BjkkXzj0omv0YxQp/ditJAWPhwNUSXQNxW0oqT2XMkuERGshKzN
FzAZoHEO6AhTFL4e95TfjgItt8ewBUWIn7/fdvB6wQoMiO4JvaUA6MnerkkV
+uGNPCp64maufUsBgStVJcklp7sOoB74+Sp1xqwtDfeBsQynNqe/qywa+eq6
iaEZm5HPLNl+8cLIs7UD/45ZKOUvulAHMPrSmoJUTv9Cpn9iuyh4smtJtrPD
XDjaexY3EfpHxJkezkFObyJRRWDSHMV2A8wguAk7GdX9Ou3DihouizBgruZH
QJ/7M8PwkbC0o9yjhP51jyTu8ARvWWP4PZ02REd76twFktq+I2L6mEnYR2rK
PqnaAVuNGYu+GDje/FXYrpuZIsyTHTGMKuoamVAC5KlRF2/uUxOw6qPjH1RL
zv4gE279m0CEmuK9u+80TDByjaCBfBWnaBtiO+tYgCefJT4qDw98juY26SE7
ykinIx2MdgIt3Kv42N9NPVBMBtyx42t8Xsru8oZaYGJyx0a9wSzz8Obb4Jtt
AE8gUGvFeA+nyt3Chg6yZNWpkbR9OSfwnRq0GPnWgi8bAahRNeYt2paqSJ5l
zjjUWnrVgo4wRx1ukxnJCUDmHjN3AXxpRePL6SEYH9vTMc0gLK94sC9QuOiP
rwCqBKBUl7n4ncIq+OoiBJbDa18pndQOUem6YbVG172WqzBvZRMGHhNJoEf1
Kq1pgd4gIjf1AC71AjQ5H6RDZdpVrLuCoi3W2qpJs5laTEo+HRyHnzdA7gk7
L/+X5VWaZJd2dSDB7gooAxxTWhVhJNkVaPP4Tdjg5MO5MbtM6XV1E+f39a1k
328EekDOJRQMJmAe9CFUgpOR6tdlSS/kUhfci9LJ30DGTurJE3rGHgMX3+j5
uPUoXIPD29YgjvpzltS21e1bJ6kb3iOCOKcY2on/swhiz+kJrOz6HDcjW8w+
3EcjuPVHFcmv+1sk/Gj3kzF2uk/ITSR8lj4WRvdwkXKsoTX1CS7pFjLhVAxx
D7O2qiErj5/07wCEgezI//nEcGomztKGiLDBuZ+KR/0KY70rAFmNYZlXxPvB
mftQMP7EzdEND8ijClmxm1P9OHE3d1a4gCX5gsqhBj01/5o+NFyidewbvuVl
AgcGfk2ynVdRuFWxf8/7hAyYW1Xn8zuWaTJK7ijRlnPDI1D5K9mHlQvmtIWw
I57Gsj8aMWNBzD6i8FWR9SL8gdnc+2BiIQQxgLjVquTZx/GOs8ms/Etup6Gt
IcEVeWk/Yog+tyBu706mYr3U/qoOF5LVhpjchhYhFNF/Mi04i8p9XVQvWnay
G747KTzycENACEaCLi3uOCURYphcU6z+M3N3cZASBc7/GX62LB0mdmrOFozv
dULQ+95xgKL1xV/dNOZJDT3IbW72Jt3jsUZLObe6aDaMuppWkp9/ZnMKIBw6
XeDMJAEr+RbqaqxeqYTNfo5QoUMtjF3eoMvAn6H/O1lTDBz1Zg3ja8Ngb9D2
VONngh7d5czhl3x4p6C2fN4GJsXuMhnQfHrTKqceoaDwgMJY8p8rfZwmfAoL
tVL00/EAyfQ9auSHdB11A/NZIiU7oVikgMTBigUyVHC+WND0X18u3QN7+Kwl
WFezMnmrHud4HpuSe0AKDwvVFLqLOOuQydeJy1cJp4QCS5+siyZfhauadEQi
f+LMix8qboxqasbBw+dtderJZ3PoW4YSOAy2OyJN+KVRR+XVG6V96ZCeT41w
V1E6+UF5VkI1T7RYmcVtaQ1//550IMsgB3EmFovy5J7xVxC/Xq8nClPCbzp3
kPZIrQmpCGacd5LGt+JpWdl4w+kIey/VzYwU8kFP8Cpq0G0C15Pu6GrHkMzH
G5hO2CKtzEisU3Qu0HumK9tI85AyeOvPCy0j2smDQ+OGjKsCrUKUP3aQgzg/
dqLHcXgBnbjLnq1IxYwhFEDWYuySoRmrGM5QJ2xriZi4NpPYa5feERrcHQs5
aEmCfLuzvx4btxO0mzeaxesrXKVkYI8up7hsCYtq/X7lhFji6hxSi3vrT9MA
Us1xIQPupi4fRBI06oZAr+OkNCK03EDxwxZa+tJI4m3leLD47e4Oou6p7yS5
i6Y6YEV5jwL1OOclRDi7rSZkzicK+C+PidCowWx0QSEWTIXoSC8v1CFC41d5
OQqtGq8KCynbEijPCEwDJToawl4RGCuuWO2/URQedl95ch8aQT7UBZZT5wyL
rP16I9DxE3iPJI2+zCU8/lEgtPfMz/rzPfArPJPHHqb+OgBU96VpLTY+LMuV
MbSJbMt8XaLeKD7WRk65N4aXEMKA8jZsJ51PvqvPcLqZcNQMPSZmZetdzA2G
Fjg3r8YMVxSNLUsAYu+lyIwsFTOypxJyBM0mUzR+zc2oxvVg6hpI0IGLrkj9
GVbeWe9n47Qmt3EjI6o9Fr34thyFxDdTem9da3eEenN4cZ2+cZ6Ou+/9BBos
usP3Iot12hzU1cdsBuy8hYqgeg8E7LcwiO2G2RbmQ6AeBtL3eAQB8lkFSATX
UcKqKq1WanOEeiRS9HhZ3zBQkzgAtnqvZAzS2iQXd5JE8NE4fRsSOlSIya7P
xiEvrxRWBV2GUxKOpZF8MDDW8ietwezDHRnZRsqYZXFRfVqqDwUq8sFrVxhY
ayZMVpCizPh80AO8lwwFrj45h7BFUmyGeJx90a/0d5Li6Pw0FH9gWghdWF8k
y6JeetTX3xRKRcEzpw+Ert7PkCRctq0sbq4z6e7ypVXE4J7UwkiOXE0rcPSL
XxlMdt81+FLVs8TdRHz+mpTBhsGsOqX1RGIBtCIJcMb+NM8Pu3JPtAYaYAwT
BG80dpF76VE8k45xq37ZjBM1JsapW+kWYwYjdkmQ5q9G+7qVa2xjjAOT4U+B
uR9/JHpWUsNcrIuhw8ovzjJbkxjxrqCl4XbI6/4ZljRbh6IVxMvGYPUw3ivb
ZksUWTdBple6Ai8nulH/YfzHSiuh98lP8h881wj3s4+iLt5GWG7rwYZmHkQj
+ooxQF2JOO1F7bRaBsPprvKDdrnpQOJuF68UiKjEKuEhZj4GPutTKt2thTJE
FZ5xHxW91sfJCUNLS6elAaJST44HSQmrkRzT+W8xvHWs445E1dnjJIQXXwkI
/BHjOvytlnbOy2e4PTYH/8x1zGwgre6xXvoRgpG5w0bIc4FvjC23KAYk778L
pcdT8U/xxhLme8W0vVchH9eI1tSu3ggaXHfwb+iFez9iVhPPuKwSIvtLtxh6
xmffEjFhYemQBGYRXahzcVkEDX3OBX9ZdXg8tnRsLSucsjva79nGrarxi0RK
MGG/e2tAeM8UEJlJ1EHrk9JmWo0LZOl+CK2jInRCSC04OxZuWbBOLx/O9hv5
GK6y4D5ADa7Ki7gkNwEV5xw+nz6FHnK3Qdo9CsLxLY/Tz/UTdOXbg/41+Zo2
WecwqJRjmB7EM7VYOUKeh6H5sE44DXBXVPN6LX/wCjWy43wrWapzrDOviayM
KKdekji9tfPeKEV2Mi/mG5c2jhovZxKSKO3KO9AZdxfLtbHq/Y3fE2d0ev/s
r9YIDumZIQcqGilS9TrxzN/tA89+rxvTYoRNk9nvxGs/W2lr/0OKjg7kCZn7
wlxQQW+9xJHW6Hs+pC9OxsVj2GHtqdS2cuTLlgWKCbmhDGdWDFVEG2pAeiw0
L0jvlIJ5Ot+gd77KftBftARhfBYtSQbjIxZ+n+JtE/U9UAkSOyjmVyjWwUZl
vMRnvbe8uQayfncDhs28+RVwhSQppFoTZdyzuAl9/CfYJ11HQJkTXYHyRAYX
ugnkspXER3JKPmheZJTvBAHpkmNrhfPWg4B484Xev4FYANC/1Ci0gj6nG8kf
kjhMoouZM2TXl0ddHJ6XpowtsatN6aHQOo5ifg0uL97ZSNNTUhNL+3szCW+C
/yOEPwYuqhA7wJlB6J1Kinp2C319Bq7HJDzhaRkMJHEwClgeYzZVEhM0ksKF
/kM4weFhYvHrrdjY32Io2xqAXdXUjheGRJFGnGmoj/rcfeVBA8iSazYTwS2W
9Mw/fFmkutcj7EiiOrTiXwGGlPJezrTkyLo/Du8ofyQGxisgZ3KV70ZPFEfu
J/VE8WYTlebdF3BS1JrkagxrF9+7hPLK+fevjfe0/Z9Eun8PgNBWsXw+kJ+7
ynncfLBwiHWoV8r32S0kPMAil8jm/Lb0bWldrkoX4Zggx+QlKr2afIeOQbKM
GZqcE0TQMUpM6aBycxqwzmKHAtI3lcsjdwcR/qwv21Ww7qEKKwUuRQIH0okv
ffv8P8BixGlNiyAmI6fp8JO0U86wDludqCR3g4NO4ui/BP8GwgmubnHF4tBd
/OwCubGW0HsC0iFbLNGdGNH1wpdwOOBYT+xUo7yPlxBtFwfddOr/Ap/Ukw8+
6v8BnQj2Vp6oTGBitOSHmt6UkjeC/UTCQZJUnUgH0yAXyDwzDm3z34ao6//w
55+JLPhYQ7rXWLj1a1dt4MyHTIg6lnWBOQn1atyYLO/cLae86T6GxiRWFlR9
MuuU+hYYe1WkVxjiA7Msv2xND7qYdnrNmQwK5HxQEMJlxF0Ifu0oTkirQ+g4
Da7oJjlf8Vpoxsbq6qU64a/ryXyQ+oDq6ZEU/xIgSzUJCDr6fisYT/6PaLLC
d0zU0EbY9OxejZUPe86A7vGbfhag0+slOpotKh2Aet4gENuiXK7QPDGWgojp
yCFOPntxNiM/b1oWK4ZjGz/Ba27yF5ngYrEJ8UasID8QMZu2bNZOxlKe3Y51
5LCeBqFgn/hZKd5cYHrpEy+ZIy8SwX0x16hTVOHUNcslP3rAd3H6tSvJYYSI
d9sb3zQgCgTerPUlKds1rrU/7ES4+3PpFgUIlUA74aHUMkje9cMt11D1y2wm
IgFdR2/mfowPALbCQPOHCOOiwPC8y/KoOgSalZx+wI3MMX+QO/7O3PVfh3yA
5QYXrYikXucjLd7MQrGeqP0/nYkAAQlTFpcTVwUDkFrd+uXHFas3w+FINqJB
EOTsaCQF6YV1ojjgR50iJigJdcAstLe603VWPTXS3tXrMYqa2dmkzz4thGkK
euVxEh9jIo3aqmSNFiDbOjAhtyBHjNK7wQUon3Ykju+Aq3kzWQJLUOt0Ozvr
2oRjJfPqYrzkvOUIBD0CveXPAsPMr8Ss+PLb8Bt/SabsCVmAu4/8+HnUZq2d
zNL3HNHS7+KIJeHTUGkhMK7PTr+BSI1p4rZXTZx7d6lpevvLfRNN0hRbri4i
28rjRU2MZmy1m62ypmljiCOMqUvMmxBqLVjqhteG9e2Uvz0Sd5I9rjAsC/Sz
NmvVr+itzZB7H9tCQoGt9gspYNH2wnFINfpczxzdTMvsC9uCkMCCiZP369uH
YdcHZKpmd5BHLRh3a5Iv+nEifHH4X2VZA+c54bFD5LYGFpJUxMETBL1CDkFr
2s0mUv8wvbtIjiZHOsAODoyDIm3xTWc+x4l/A1dRfK/Y9SU/+qVPYmooXKpQ
Ep5eSsD73dEb9BdD/wQkB4MBaAWoP8b0INUmPCt5+w35QLVb4+W1d8UsY8Wg
jvADVUY8mhG/wn5jhUui7cF7a62vVhvrd05Sh5AC0mUx2l2KilNNqSTqXz28
Xhc+PoO6I0yF7WlLikwm3SNzJnQ7JUtFnoMZo7dJmqdnOOtWxkN7jXYjxxs3
j1D2Fkdgqob1/JXB1UBUdd7aa2z/PUZxpzsHcdVqJfuMawfCcvsdLP9WwXrK
DvxmDClFRp78EWWTuw+hOUOQkzomVC0KT4yOzAu1SFucdlnmI/w6Sl0pHKMw
SzE9WGMgBMWrbYIhuiyvMAKwcx6fhPexT5gUZU6GNOUitEnCvm1Bvt3M4kii
sRfSnnIQVYBYsqClLHAefMjn6qHvuvSl35AqEcC1f+2naOcjFfMbuzYyIOG5
q5BRzJ92G7QV0Coc3COMLnqUJ6cY5+ANQHr0VV94OkcEFos4+CHGK41kR5sD
VhprnZRltxEr4vkcduuYUX0OeNmm9Bw+YiAa1L1/oWmnodz6kUUhDYJ/Y9Oa
x5c4c4C2IJt+gXbKZFotQZDALcRnf6FdNoQxCQ9NvUeiZJ1xr+Q/+0kgoe8a
SsmzsysBFf0u0vVI3wU2UhYdlfxbz06tzrbbJcwIzqBddmjQVFB7UkrkJYJN
Yn5F/UmwFd71Edwkjdt92d9uwwL78kZiqcwiS8ruBa8gGh7K2FVUvGbnys3s
O59djw8O72Dkwp1p4UqLQPKamrKUpeO7wJX0K8rqtrheKeP0OeyDj7BPmfAM
nTMKMiLrEoerD/MTZt80HjwLQikV3HNtpp1fb0piCLG2hNLMlqk1QzQsep6U
Lv0OS8BGjNiZq9CJDny8zB3vvYIXptBsnmStlFAxDbdZurUdMxMJLiUZ+yU7
HJ0rUeKL/swGZmfyajg+pXJxu/HDtZ4uujK3ptgGjlNkQ9IzTfXXRlpTyDon
GXmphz80T/qp8LEU9UIQXcgSwG816N2kKu6yAUwCDOp3x9GRdHAa8jVg+Uu/
XhqDowpe8qJ63B5yQDRSRzuzTR4Lyi223OurGl58emdvlSulSvEbLminGjkO
6xW+OpSQylBAhgmLPOm4enCnSqG+2o9KbbqITou+Bh67NqixGwC1BMvjrHqH
u7BD6AYVZmPmrgT4AduwlmCg2ja4YdKjSlqkovMt4je3OEPBSAxYRcjJBM9d
XIHTBZ65CCSceF85b7lHQlRaeHgkfBmGAA+WJxfFfXro63CRFgjpKi1wMwA4
ypS+2pozkjgjWMSoY+tXvCGav8MlcT7u0aUkRXOWaYsSxvweCK/HoR1zXhHh
MEi8cSLeyeNhGz4NTUTWUQeYB2fYtQWyQxv02y2f69Ta32WeGfIAkQNKD4Co
SbrzWTKFPa/jsWLlrc1104nYpxqVsCg681S2UfPJVzIkF1H0C8gKqa/5Cmoa
FFPENzfNW0B21du/A/qlvhVq06XROLGglyvj1V9Z+vERZsWs5w/e9s2wXRaY
+kalbklw4QDk+gepPP/xuyq0OhkaQR+ZFZcZgDYqGhhP2mqWsSiI55V93kIE
jKzrWTRKknNXytyg0lKMKdH4x6ikTdVQSF7L9pWeuSGtA5qffQcbS/Fe2yTn
wG9qUTik1KfKnbu5pan+wXAtNREKX/bKXcurqucFFDVXtbvi9xcPOqR4SfMJ
64qhM5ZRhqamFfuF88KoMUDMJzJTtRYQqcmeRJCPkhc6jsOBkwGcvZbj3rjN
JCTiNgI9eH1gvolpZZiVvY3flqVBtsTp5CO1vqF0BCI0R0ZmNEG1W5uEEftw
0BgCGxft9nS5/pLZsNuPcg1nBTrk6TXD6LZYDmZMZ63HZOKQ3NAPogtvOPFP
eAeNi1C9dEXqFNQwo68EwuBUyS5uvt+Nc9+TdvuOrKJHPBJKcg6M6PbN2N2u
+tnOLUQfwnojEvJNEl7MYP2EPB6NhumhQNAQii7/AKEiIc0GsfYh0p1KDHIi
GNqP4pEFiEphIY9n1SteynUr4KIw24V05sLGg5UBWRuY7yOXH3Br2XQ1wDjp
SaTDDkOLLdC9gIVoQg95f73R4PxViRUkVV1KXJkGZjFS1WfpSipYJGkzLgri
BB/H3R3w6o/MDtuQYGgT6HCyxrBq89qcxwRMsLyo5kQ5KxdmrDgjoi4I8kjQ
8y/N7IRqDPNZQTOaJdgv1oYKhRnKl47g0n+tfEEDxNbFjUsbhH0pkvTLraa1
I9WRfv4dCf3nkrZSEheflneP29CkJzb50qi/WTqjsm/lL1XsmPObQnCtr7ha
sxeppmYtsos5SepdLmWxbzzjLCOcwwrzVYKVnJ02GjL3vwrMdz/d6gSeYtOm
nKQde1uLYqVuI0Sof5+FxffphkizlUVxvr3wkwju4NyfEBGHhqnjXHhxuc7K
3onfM/utZ3Ov5fhWxTTkOImULVV6TUCYqEMHRJJRutI2HtaJtnzkMR8oLB4x
8qf6BKGHzv8yUFfnCpxzZLPr2MF/rqwktu9LzDEn5z01MYwmARGmlSuz7/ez
CAuns2PuG4DsIeS+h9gRwZJMrrZpCcWJ2GhfMp9hh5gJtZZ/1Q4w7d0g7y1+
KnP33J/IBSIMhhnQb1kE56z2p+XRL1aX/lVPl/nld5fU4FCVTFxqNrMutelw
nlnX6l7966DXXd5DiGsriXLvQ0IdEyu3WZPgAJtH9n+l1YdhBq5x0YIEJP02
mo8nSDZsK7LcBeR1Le936jWPs0d7Fp2kDlZvi59FIpYfPE4T5QuOyGbax9oB
tC93Spr4mqqVh4lM2RSstSoQlnmaaWDbQDUJ0gbTwI6Kbq99iN5xnDKTdTnX
JFD0pDpgRyR/k4pwUIGhEXza3JEt2s3lHQypqV/xtSM8NS2OI8jio/kDcvaF
erAds8gVBUgT6UYjtBTjPPHjJxfTEsKojAe/9TYc3wV1TFJW5rfEOiWlfLQO
1RH7GcaZGBkmNK+/IBghca3Xt66nRTgXODcJvK1DvIlFnCKMV5V7Uce5r7sW
A2/mkyiI9gfs4jIvz8iXxHpbXS99kGbaPPURA4Rjj9NMN4UfDrubJdgpn+0e
tl9wUmFKWR+vYrVCNxtfHwtUjBaLQPmjQB+6wyqYmYy6mqQQEGW1ThaLnd5s
PxxKNZ2+UEKkCXSQBoSORHaxgTn0TCTWT2AUhyN4cTM6R82lqxds5XNGNuAm
KgyEWMTg+gmPXGy/rD1i9yYPTcH/H9/4vwAICXp4o1SfkPTgBzRUnJv7G2of
lyucZiYAfWS5h0ckTlUNBGXrPA/iZp5oz+tfitW7r/sjWWiP6qC2phHz1SHI
klzoKrfz0m3D6216otk6ZqERkVugZ3tb3YKLwEGLaWGVaEoFeTvZshu0qNag
aRhIVnNyRlBcOQsFdKPOiHMXAhvvoxCYX9IwCmQsLV/7xuyLyBjg+RZZqPpf
0a5B7pNa0TC+aDRfjT/liZuGoF0RcDiGa0GjarRnsDOkPXQzZQPBRbtN9V1j
vxtWk2algdeQ9J5d0zGnpj0TDcOoWq5F4FIz0P1Fp7XmD0zu1cecOKF34qg1
ifXSRnKr/mXnPeJzE5sHweaQJHPSS/HkgiqV4Pum0n1NXTZ92N/j0Q2eZxo/
Ke89RzW+0UfMlU4PXCKBZqxe0RrvxQITdeLNKotM9kFscCxxy2hMAHjdoPUB
TlsdJ9m+IouLPpsXP86PW7Vhjx+GfmgkFJtJS4VEqloy64yn6k4i8mFw/sKU
Hp99RTsuHtZ16X9FAeqYRqhYJLdKNl+df8On/vVS+j4Jwf/rmJwbU+Ud9UpA
DO1UpdK1RPzBxMgetsecdPvmZfz6ScXglRr9nyg4dI1ZaZyhpRr/2VyH1yX/
NWJP2SPVlQcGy+PvUlTK/Ak6h5QYY0e6UY0tXBrd3sr9zSqhKyuZDQ5fY75S
PdfVwm2ZH1L6V4csTaqvnijYmU5zLQU5qdH1i67+TmA8I8wTXKsp/XrDYSGC
cMW7xB1tVGgHHOK3fMvg7GQ0jfG6y2LVtX2dwH6Q82sdmFLwNKWBYUAjcwxH
XdZJm4bg+8rO/nyNunYzSYxcPCG8H9DEtwc5vXCqwEe7sCFeZojhWTBVAJRd
5SwB0XwpcavWd2lZU+FcxjXLJf2OApIEuYC2lSblyYspojp0+Ww/Y1JT+Hep
yaFBlw7peQ7Fx/iUdZpWLtfRl6/jUvi9hayWkvpV/+QWWQP3V0fudj6Dk++/
ruzLTpiRBRhFn+3j1qEhcD2bcNJv5EaWFfuiwx6r+EADGeG+fu9lXpx4nHc5
zxjj2ba+i1LGzf2HkfOgHhFHAFTYsPEZdvHQ1tutkjIuA86Z0ssshFBAKFXQ
XW/gOyOf2oNUOhLyngtq/h/k3br8qvLNfpg3bHcss9SbRm/CgbfYa8jnJ1lS
DudWzc0Ff4KOUSxKQfxkqsMIuB5PLtTpb7Tt2ChPw8xLBuGcqzF5mq+CkXzH
nkUsWCB9EpWywLJPBjuQiT0/doX9CWAlo0nC9GFlKxUSEOFhkY8WeQqMJaqX
UkSTWrhUQuRryZMFaOw++ilP5PYhErTkZR3Qxe3noOfLpZyN95i+VcodWM9K
umR9lH9EfvYZDjLAZ3gLyLV6EjQ6zDNrb/ssWe1JP0cmEiGCG0IgfsoVG9xt
ufJKHx6ShZb2BZVqT7qLUcUJnIv2ME8sHKHECtv+87N1vKEctshpKQh35eMM
pbww5a9F0Ewb5YwNIcuMh5RDTB1l1JRVlK2o+OVse1mgR9ZYVPL2X3B9kxlh
FAnA3ueq/IKvudMUtrTD4cwYeLlwj2vLEYijSGP3a+DQ7FojG6sEvrFdL1jC
ZRJqOX3t/Be/g/RSy0pmznTOp+LkohmRo7AV2bOV9VxyACXIruMKf1ua4urm
OIth0Y5r25JAQQ43Qc0gJrpFABrcPkjkxdqgZQRlID07eZJrcEl6iZc+21SV
2sV5z39kvCW2u84xEPLPF+eS2SdzfjKgsQYKik6LdY0eUf2yVP5thi4CSjxk
9Y1nlAkqL6XGtOC6DedYddXWKpe/mL/UTPzprdKHQJ5aXptpVNAIxf9B75cc
+h0kXDXSSAfDy29J3GiNnAgAQ6bxLgXjDa8aK1alPimMuypIVU5ZfSe5kiJ9
61jeEU9UKlfo+jgyeVw1zz0GLV1vU5BXnoMaBJtyw90ZD6FMZxRDEJH3g9sj
HavBXIhKZoqa0U3hsIjpOtLRZ7NTbNli9WKHVOHFc2WLfUSM76bfUrZJ5bMK
ToviFHGOaB0LVudPw4LmtdTkVOc/mgSP3vEvyjENVEN9kLrqlW1KJDsQ80In
GBv8Ot1U8YPk1jGyraSAtDC43OWQ4hgFCziMgnhdZEcK6qiZmEpNslIj7wT7
oZx/e7+QH8DxE4ipZ84V91AdilEWfyXZVW41r12hj41WMUYHPqFgDNvHVI7v
WVyMZV3t11jQRFzPqmA41ni328TerIs70HoV6yZ2r/5u61KxhZOP+9FgL/Cl
SSIaMUo7tN2s0LEBL2ORXL9wVrU1xIt4wOywQoe+4YVBn2vqi4983koVe7FJ
7hiZVKUSs3OBIjCVUhCQOqtwxCoW8Cbbofl/vQLPHyh1STp1iFy6y/+p4jKf
n1rgUbd455kXoEw8I4+e+n8GczfdkrblyWmkPUwWlGaf6jkMxqBKYfV1x1yu
5JFg4Y1nnRcBznGlvn1dGVufB5LSwqe8qy7Q9125sHvmyf/78yGKoFHEjZRp
s8wSQ63lP7CJJvdQ64zl6z0Lrr8ug8jmQu1e0i/LhbDPwBMLb+lX6WFTAqFF
0vqIyKgcdkJR18YahXMMm9AXkRqCAGeBvxmwwWhdKn2ItjPhfdp+iOC6oBDW
YlrwobSvhjZGveeBIPd+oin+CvvNe9cxsfYEAz/ybaUxOTG3hX5Ors9Ims2L
iIsoBF6SLa1RNKgWBhg4fj+mdvZvRyjWqD6AoHCUD21KMIobKU9LGj7wk4ub
vAZ0cYPxJC4wIi2C8IQF94yrMB4uVc6L2I624qZuq3NEjezgnCA4uq2i2zfy
5RTGW/9JEhEB7j66XiUDqge6HqFdmu7v6mGuA/BmEJFYJXs6JJWoUtty7fpO
4sZWAZU4/xdtBP9tqWdfppUJJcK3o7LzadmSaB7nCOfluGen1nXatrBSNv3G
1iM6ECDk1weXJj5UM5jjzP6lCiL5Z7knnAlbJeOzix+JvNhuBNPY3NCRXsA8
dNdWErNJ+n6aayovf+W8RZDYJ4nUQInnvG6bb1N2zsUB2JwVRweleanL2scp
ZVNsOMj1BQ51i4wrSZ7gVV94M+APvMOBdtlxu0/48j9d1rxmsFw4pVSakPLc
OcFrmbuGbBEoRNxz8q2NsmDmAM19OgfQ1uGa3WYVExMPKFYvuaQUaumcp7j9
V/CjhxKXkJzD3tbJ+JafV4uh52r8nlSbNUomwtQMUmhzTyT5uopzPDQla32i
dv8IjJrpN0/FzPjmdmzIhkE1NS90oYuUKNUb9lTJyhXvpoEsysBQo21+cIt4
2myMYLNRdua/GLmPN23oZtic87TM2PNk5+vS/7AILCeRV/LYXMyhQTIUQmhW
iYx5PO3FyqKLlIsjo4/5XQbZCW2ESPKvmiSa/51J0j9YPROv/gfxNYVl3eHP
NSWY0vm5FVFUvFXZUFepwCYyp8p+IC1PIu5zTIOAt4ANW1Ar1SN1zZAaWzx+
xaXp2vai9Y7te163PX3coNWp18WkxZ8NF0Qzb8j5Iy92yTXTW2GeyvW9Un7c
u2o9v2SkAvfaNM1FAgQsuJA2/RBTASvhLenjzvSQFkqN0G/OkB1qzqXI/lgD
4oelg5H19x6Cg4dLLCnp9Q4fY5efoN4aCsB8PF0aEBJCrJR7Mh54N9pH+/HN
6CxFoIARgVlHnxx9nvHCBf2WGMvYtPTrw5t7wtHuQ76sU2J5LwST2pR4jupU
w1Y/rsG3yj9LNtKVVwpkIv8goOUo7vXHWReUWbOJeD20PotKY2KCOVR73SPT
Hf724/6Sk16hnpLlPqtA5LMHizpMFFN/4lf9GN2+GzF2/AgpiN1OvweDq9mf
NB0aENZ4T7C3CmqjhiPU5+9GlvgaL4tyyy29UZQQK/roW3TRV8Jm1qwgG+Sp
sVsmQ6To89iYn+w/W7P3/yP0jxd5UDlviBFNuQDmX28P/kYzREqGkc2gHL6u
S2tGtl0yGfObGIffCWcTxHeQBPYl4d5mY5P0jTR9xrh1W/MmUyshZRruvNud
lCA50dGrmeCGhZzCn4h5EcBQwvOrZ6MTQwYbvUAguVbf9Rb6O6PHI8XCik/E
c/YryWOrJQk3xBQjbE0tir/p4oWkJ3Mu7Vku+E7KBQ2OLbelQR2w8y3HnSLy
6YvSTr9TZqrot+/dO1Jr7vlq4uUkjM5yxyZ7WBm6MAPuRLeOEIVrpRxewrjw
aljD6ZplFgQ52l9MA8DqXJxpYd3z5FWUneMsjJI48Gcf1KWyBbOl9BqwCfLG
DnVbAAW1ZsgjTUj3xKWbQAWjs/RONQSo7ttI0hB4fOpqM6EKvJJsn016tjTY
Wlq2CKVBFpwowXvsdmhkvUWYbc/sv5Oxrme5xqhB6NvlggTRZVKJRxX4/OYp
uondz8VwreFdwRIoifcswZ0Hos8dxNDVY6wXyyKRXR4mopuqGnkEHYxSE1va
XXmYrPjY2ZbRPhKSFRq8Jjmc1J3kGojv0yH3siPKJbm/li/7iY4x9636A5HA
qnZv54vwt5Nc1brbnKNErlA2lxOWjaBDjlVhi5/lwgtQFzJYodVC2SmTpPL9
BgYX4geq13esgVR9PvJt7uCNcGEgYDyJkI/jWu9i8s04sWp+9oyX6Z4yoK4g
H80EMbOfATPCMig96d8u86emKVjjXTdEIoUCzffzEgEee9ZlOOP8jeG0iJIe
BMiRgUOeYYnjZICz28k19IdXdDVdrQ57StqfCN0ywOLJXjOcXQLI81pYAA68
o5DKfHKioMKyxS3S2DYGJWgaA2hz2LFlxncEbXdyKxCvPsIe1T2E08Q0mwRS
bwQqou4a5uVEzmEHtfAw4gMjXrermv+FjZMq7vlSjH3NAgVNuY4qhJqgzESG
I+8tPKXaREwfYA66rE56pf4bwPk+unFNMjGnlyN7uUXa0VyphwRRAg0DpxRZ
/DMOQmDbwFSOm2QRHXGN73ZdLNZA6oUYVXycWhaNP62qNXf49CPND6WRDrvk
M5i5KyXJIHVoPDMZ3eMVg0DcrwDqgYMTB/yqOwFS+cBhg9juWJkHHKye3u9I
Epql6UhuLWdVgV4PSamzKmyXU8DBfgLl/RRbzWFQFODlzINH89m+jYE3Ay1b
SrCjPokwacavvUX4pZYB2usj2qwio6TiRcaoc393sM0oWbcw9e0Jxp2nKHSj
QiBNKxvGjCdrWcGyh2IsNK1oVxNaQLFGtxmtbESVp2dXFQR4CqqyxuGFCP+Z
4DS3vsFUq7Z5m7rHPqbkOg0lv1MZ8r0wSdkN/aAfOABaJtgT81D0tvawNVex
7jDfwbrOQZzDzujTxA2iepFg4FneM038VyxdnvuXIgnPubAeHsJeYKn2cvaq
ak7bTHLCf9dVJJAVhyFOuXkj00anE5akw1bJJfqgPMGC+9kHp32CvWYJydHY
vfan3+iBiY+HburNpkaBCz625ImwheUuU3+ATw9e/g9J7iDMI3DUF/wCapfT
2dW/0SIEE55HMF17KHaYM4AGhwlmaWp23EYj3kxCrPbsaKWqNOamOgHO8Iqe
zksF3FP2Bakxc/3ZeNaFLJrQ33Wu7iHGdrmZmttAxexAJG/NTpLrT0HPq7ED
gA0XruoqgmmcsxJXdodVdGf/K0Jd6rr2aJ5vche+ZBt0fzP5bkH/yz6UPKVK
XXGSgXHzl+iFORd975llCd0aQZ5jW5NaTpK2h0A1iVN486GZbRYBeEiWNCeg
trR57O03Kg38fFE1b8OgNpyoytwIKeXjdCf4gb/EwjkW+Kl1pCb0RLNYjKf7
8TmDg/SLg7YRtm5Ig6CNyCUPh9zQMIpevfq9OWSPsd2JO9wC5UNSv1vyeITM
WpOM86P7I5hjKdPn8OMfr4QCte82i9sT+5gYQU62aTqJOeQ9SSHUu96jrwvw
lMtltXNf+CjzcpJk8Lip4qCIIjgrjK8+k93WSfNp6Wmq4nlxxDx97KP2IKnJ
ECkWtaNLXdlXu4mmXP9kuOfUyokRbWzwGB1MC4WIp6ntmxVgPxObFj1x/lcp
sJ9XeafA2IUSsnyrxe7SsdYwMkIo0Gjvd/j3pixKVUszcXDs4zFCxnx2f4Hz
xb7M4RTTGO+TnO7HlOE/2RNjlAdArn36ApmlhQgEYvpsT7J0HEClnAC5Ke+T
IQ1ItU24XXuWKgil9BKJLIYXYWWGBmlR7jp70wa0sEgoqT2QcgStKnWO87oS
6scIfbiY+aL+xTEwaDRkoYBpnwcHng0fLlb2B7CkqyIFWhNP+yr6BrYJa7ni
997hVtiM4wAbkRdOUh9X85E5q0ioajnuoK+TsMhQF6VY8HQmBaT1R5qMdvwS
mHSjjZuqcFnxA7IHGJMNSTE4Z8iD+4UlKVT82MALTQFjUf67K/z1SiLI43kU
PrKUu6WD94P6iVj2QP4zkWtllBWHpSBX934TYSLhQHx4OB54/nGjt8ujd9J4
0jKsCVdwecgYgda/ZK1eFaccyNDkXyLIi2PqZokHJBK5DCu6SkxBNKnienY4
1tzg8BgAyy21ZZu0Llb5dObZh92+Rx63OdYi9O3CEbFs0cxBrdULkzETTOa9
uX+muPZIJdJgX/4nSDg8TgTMcdfcKcY6FvEbH/oBqPKUvhWni8f86uB/+CCj
ThaBaJR8jfMFcjzgk5uaP7dUPh8YjlgUqaw3CZwvP3NnYcnN3s9Q0wUzd3Ba
9q8RbRfTsPTUNwMVFI3vMbS/LCk4+b5Z0of3h1+vMq7NW8HQMa/bp392Ah+F
/f7ojNj/oDmoWd9aApVJp7BvKcjE2AIolhbnT/uP93cRc91xgMKINPf69c/e
iUX6usrBrV59IEHyrsILqcXELez3Cvmoo+qc0LcmvoE9x60ZJ1WVaklwH/wI
M3y3jFcRafvbI4WGIROoIQmF7DQ3C1IK0SFyYlBKo4Tzb3D3IlHim9uq3Rey
0coxdYiTKfkZP/EmqViKz0orJsshTQQuYoIgSiTuTsSZE/2aLgbI7r0zJexJ
setxZ2TgXpX0+/8XqAvcfFDA+CMAcISYJYT/y0iYJlf0IfDT93Cz0E1kiU7p
rVfAYjAu48XmOUe0NHfcmmjtfJUMA4sgc0GiBZH4Yd3Np8PcVUWexZbtdazV
krl5BrCGUHEalOi4G+P+Diu+mv/vtP5TRauDyglNSMF9i9tILGbFcqgVWMUv
jq4LbG6DqpJCIVSJM3R+DvT9DyFvO3wzxEiV+mjjB6G11mCFXi7el8Bgtm+n
7OP4+WByW34uLc0iOnzRTE4xnYhet5a8x5x/OqTcTzCNYUO5N2VCuAVtmt5W
vX9rfIdGtHQOY+SKv/MZEV9MP6pBFCcwQpJ27JhWYuD45EAuy2PBYXxL2FI3
eqaqBF8TgTS9YQCIlZYs59CW70Rcfhq5yaLnZi2qKYgAHDJNIIvpZDZEALuA
IVT3xVz6VIt4HKZWZLI0sRHQJHcXV7WZcO40TJLs/GeP3mFyQbpkka91W+tr
h7pb2kGEmESRjIA1pluDmRyh74TqMP5dj0+31Fa4zCeU+KSCzCrZcdiNtKH2
VJ4uuCewCSxAzBgovxVOh8ixyX9EB3maK5CtQ4bRRHS68Upc4ozsfBlr3RRz
XNYesP4XDgrc6vfs+gNwXRWU21DG8VPW7is8uSuAXx5Yq4WU2Y6Fq6up9Yeo
ttD5G1Hzg1J2zVZ15DdEj/aeRZzzijuwD6GMWodRPW9mFzcZxwQs45SNWa+Z
7fe7omyTyzxULD0wvvA54JlpdND6W1M8czQPlwiEKHcGf99Q1G6X3eFlFXYg
Jkl6ORt5AlFhf8Lt66K3ZgBFXltaiAkXqlAqkPiAtuUWBOG8mXWWsTbRbmsE
AfkBZKDZJfvGR48osNe1y825n+i9ynUvxCrwfDXBvINvLVtu34SJcb8/AHAn
lpk/Hq+q5i+XCD5vISc2lWpCNvQrisxqIWZOVE103x3lhMtejVfYx3yWi9Pi
bUiahD9hXqZiHhgCNeioPYpMe1kdYDIbWGG03f/Lr/uDLTDk/ELkqBlliZdZ
7rQqCTTE+o4/tDfNJm68+5gp0zTf4hRcdPj+32MqSLteLYbrhhxjxKI6HJc+
o4M2s+ZCUyu8xr3wjSZ5weyDrhKl+xzrpC2hf0aegsWnGjjfptg1TPJVDe7W
3Dslgg/oSMd7hQXiy7DECrQAjfjbCtJRwwG688FJumLuL/dMX6MYtaxcYMfb
Eh7nFhxazfxnC2fCsE7/ETN/4ryCBoMhuk6aL4nWgiDmuskjOh++POntrAIn
DIuzWtOwcirS4JxPykMi6CIi4twxlnDr2B0QqR+IiZfkszsQ9KIprIFJ3e+F
DlEQ9JmpsBFdwweU60IvITphwvPBlqkwPTu+VrWjVgCLBLgosztrk91L2xh0
x7XmRimrSZqtilrvcTTm5POPvAhW9/O7oNCJF5Qt9ploBkTz4M61pd6RzN8h
bfEeHH6qmOFQHMJK2coVyM6Y1GP+JspjinVqBxV74yaio0DfocCKZQyNCbCC
VJHZVCtuquhDUQJBrVlO1XHKtJclG1MXdaV7F7c+D8hE2vekQ6pzTpl+iI9y
GvaKVL0n42nBWmfyG9719aLqjM3g0DcNIF/WZnHZnpG7HRfdst2CGpZ1N6V9
xlfyhWIL4//cFVxhG6PMjpipQ6ESh/LJU+5Ae6BRwFv+wjrF1Q0eJqdvhdhW
iQgi3Pua2sMqFFjheZeB79C8h+YUaEaOX9b4z539ir6S9Zpbc1NYkX1ypy+o
2azRd//nXJXN+p1/UR5OZOvxdIZ3+BwH6jBjlxg2O1uo6PHjvlwrFpDGIxeg
cBJMWqOqoEk0VV7WWXpssIxSt/YNLtsrd8OWotbT55hB9h0sTePLt99a6YpX
BEPMiy0UTj3OkgH+DlEQC8LeGML7PaG2lfRtSYcAp5UsPpUIxJG2Vz6HOC5y
ymu6p+Pnire6K/5AQGpEXgj3chNm5JyuFmqh4Fkaa4HL5FmQX2Sj4AxPmwJO
OoePWdiPlh+CID/UewT0Oww5cCEBiON8XRiE9AKkCW8C09V6uYMrUuqJ1Syn
KovpJJD+XPKMota8r5mDiEddUGwKCqqHxAKKyprfToC1jmbOF8KEWSrnIS3x
6eVFJAY8PZpyWk9Pc6o0hfuEqO9n6iG7owQ7peV4UdMdVCJWu57WQTBr0WbY
y+N4/a02EqKbpMaspmKkf7dFmjqbSCVlnEVojaxLfTwpNLVYSWmbyOmUf01i
w68VAbFr882EDQaannHXsDOS+JsFTALEW+I+sWht/7jnMZs1LQlGtOSnATQf
KOCdkbaAzMVj/97dCvyPBSVWMDULwab7eAtQ/wVlh82kkQ19XuwRUHwUi9xR
+4AAcLkmq+ppmecBaP36qvMYv5UpUpUuhEESfLPxfSUgyRJs6QtGzC4ggChV
3Nv8KKCFdnpPUMe3Qc4hfIewOZ8SnY8wt10iIgqd+NU/OODRJ7AVKx57YiQt
7F6FuOlFNwKNXdJ1zqoyWKQlzsj4/rrwF+VY34QI3mjDUWLSblt0spF6aoHQ
qEiioONSXp3XXKd9qma8sBC+Hi1gyDbcrkhEKW+dkeAwJ1SZmiciiixGl6V2
AlEdzK+dmIuyjPHnSU8bvSK62/5BwMuNEjUdDkDI7FgF5/A3nS/QCBU110EN
/TZZyqqC0UvI25UW2SxMILaHRDSJreHxx7XL98Q+AveKGCZ3xESLNXoWuukD
njeWN4UgTJ1qAW1Hu9oZn0ka19j8whMs26qYsCuusUlUqIwWwF2XQJqAdutH
E0hD+rTGWWmK9sLWG/7IvYULXSuzgEiywHj29YoFOtBr3mG5q1YDh9/DFgxO
uH4DZL2XCgRa3VOfCZ8cNvf9YXhINj4C6sOM8wKtBhNgFpBpUOpSRX4IGm0K
4i31Tqxbg+V8lGQhj16GFnFgzhDlsY01HW8ETptBT4Xlpkks0jUolsqPeIht
pBb5zMMI4vF20bWG6HP3M71MCpLw/6ulj6+CmhSNHiTdX0auraW97zY5WdPF
ZgyuehoD1471LpCrL3H4yG/wjudUzZilHvp9xkSdHSP51KPfTGVJktY/wsrq
se/Abzl+azIeZGabHs3tb7xnGyVqOeOny+A4f4err2jXip7+yRoePe4gpaTT
IF9QLnjiPHNZ6iTzy9UD6M1GV4cFsohvyCnQq6/GSd7Twk5KsOtkT8JodEKe
dSZF/TEBLhX9U9if8sB66EODYV0YBhtY5Du8s1QczHgFBMWsUbHb7hR1rk71
SeBk+UYHpwr2kntvPKKoE70ONO9pimsvjOz37EAfvqphfs47RdnPFtu8eR5p
NK8fXcMLzTEQvvB++i8nXX7PrMdX3/nl663M2PY9Eg9u+swDgxzyvipWqOzr
RlnaQJ2QOCujIyCI6ZmmIGlljptYuoj5b3KcZmVPOsN5Rqz2EBux88S+pDKz
MDNdbV+zjU/gx1kQNM3+2IGT7GfpBhQ6SsreXMPxMB6AL/8cMheH3SnLEX/T
d2sVdH2S8yAPzLLhGCZJClF+a0cp70eCJGI5/+T7Oy2o8Tb4dn8RGZK6bMkw
65gK4TM+PFKP1jE5eDpSa1oYZSWuHiR2XIxnNfQrK/ugzxvPhMBrWt1N+aFc
edNpg9/xyj5+jSX8ob6KYDY+kPlQGGmibRGbuYTGO/KVHKatkcI4ofqCSvKS
NL3svKtg55NkqLpCdhXeInAidkT3/Rj4tx9xM39kKXxpflamLAPn0Wn9W1+D
rDoyALh8qEy4rPL3u9lm6gKntNMLVtye9KmPZfvfz03KGB64zwiq/7gEtv1o
OpzeQCvfmcBVgGIey1EGPnto810FE0SBZW65wg9JvmnGRRh+usoazl6MQJ/Z
9LAJtIj5b6ZxHXhKiAVFwMO3CGxLbxig3cAetXuDFfqTxaBOARbd470pjQkc
JJfXXIFz3n5tFb8EdtQLgORMd5/uVl9ZZmbbN9/hLE503G+EHOpkvPfM3bos
BwROVCGxWfdjDIoQLeZBrJECntTx5rk11pZ0taJtLMNd6lBEn64SxQUTacP/
upH595sGSrqaFt0+dvEOeH06jT2eCIfwN+ztyPIYg+JCQ0SD35B4Mrr/G3rZ
hO9qd9fgdxBctsqC7XkjYY1fpCEhRAxaNPM09KB2am06O65wboPiaNF9Bidk
NhqjynSNZxrRgo+/eeHJ3zxFvFIJhTWccHgP5OxonqikLwztIH5aEy6G1vfY
lnlp7+lGi/S/9wI/GFtpf2PmaBhpvJ0GDsTxUUvv29TMj3PmOhLyZaO4K7N0
VrH87rH91UwoHvJUp9qfWF9cCLm8ouNiwoJ4FVLVsnaW5lKJeyKzh5S9kOUi
hwGcdwiyDyJEKZqxxmB674/0rm2sSSB1gCPtJBj8k3VjIz9DZWCnHIgH9cyQ
hMLLVSPn0B7yXCbmu8ngWBR6CIPVNm2j6DKmWP2TpIejVUXcumXDTpfng3Ob
6Lb6bEkcb83BdXD3fdKoW2M80MNWcwxdxFlixVfHJgeXUpFRve0YtuX4g/k/
TQGk2+gMdqqsyqYHMAbh3qkVR1I57uD8+fffdbMNt8tfMdJcRWmmH90IbCQY
pDkb6JVORAucDzdxyXkib8ncBPiMZJJ4/PxJUy0F2V3hMHrfRkcsU4xE1vXR
ZcbWcgak84Zlenl1PE1vmU335QO0jict5CSf7CsrY/+3EM4lFYe7fG5c6rG2
oy350NQ6eZdqdc4ztK5I3FpsH+62PRkksSCw04aKgFPvBNVdN6R4vI38KORI
7lFX2t1tebij/ceckmKh3fHRhZ3k0ZLq6YyZ4SVm5r7iksE4rx8YuCkzynIV
VVCHHoX02z1yzgbKGS6vJEJxflx7rquCnUha8txhDtesr6cC7EPji3d8XkTu
DCE/V9u6YFj7+H7EDcTQ+9iBpdbhF0iOaZ+T5GeKZXMVBgTlAHCJb8/YAeqT
iy+RNM5n2yfb0eiutjqiyiIyUtPayhvf4PnqT1ZMQIBCjJk9grNezLVGzvPi
u56fw0N50FD3E5ig6RLQ6/yf5SVfKlqKbh+8stzdjKUjsBf6J8PP/1hEjAIM
lcAjHD7CTuAdWD/cY2wyNbbTmI54mqliGPWWt9me+nZaFQv6Zr2/a4iqonrm
i//mFVAjDHy6Zj5HcSHXM92QhKKutBZZqv5YBdj67BVPHlxDVMDAU3bGhcSJ
ZGNf4f3hx0JVN2GTQuSOPuzWahr3nnsvHx3YZpDa4HpnAewW2Alwq6Y+ki3y
6jIza7Q0O+GCGnUEP5o7VDN1ugCiCHoLRdE8IIht9+Fox8i6TnTzsIpQsESE
tp2jyN3JJ67+Umf5mw/p0/7E5EkcnYn+TtEt0NICecDlibQynlSl2grAFt+E
4AnP2s8OS6PxPUf21g/to0IraMGd49oiq2i0alK17HJ5kS5nKMpviSXb7cRM
4dytuQzuQsa7ZDzLxeDCcPX53NqOslMXvEUJDZFiqg1eVWzMmhRDc5nCAD0g
UZFqiS1zO/0aUBRzMaOh0B48V9XhzuR2banzo53x6qsAxwmVp7KtN/9IiTl0
9beVV2t1PBVehGcuzl7IeUJqNkiROFzvEmvlF372KgLlCtFnnDIIIHocrYRS
VFlUaYHrymPSnA6WLhut1SMGYEt1aU4ho/1e+9GpDSVCJA99RUG6zBb/gghl
puFURul/5fMoBxXUxifng0QNWnkPrSWD7TlgftsgX0ZexU6UkiFIaDvRnpQy
vfem56hf71CHyUJ/XQaoj8pGuaoummi92s0Lh2tOzb+zcrY3SfwB7+2eZvN1
eQrMPdeP8TlUoQSzYSIMh4tyks2YuNl+Goj1nGyatLuO3zlz6a2IZxYWa9Fg
tD2UrTOMCoCzbiHE8/1SsLJYbmMSjbWbTaKL1eNt0hcvFB14LLZ2uWQBaxdp
EWR+N/yIKzyDtlZn4uM5fPlTqOp5WEuNKflstCFgi6CBUlYhp2Zfjh4V80nZ
Sio6znk/pE/O3/jxWXI4v+dUE+41wvTSfb2Y0C+TQ4c9FWyPHu0hsveCGuV1
CgSGN34UqRpXoXsqjgp4novSmQdQsvzCpYhrapr6gEIVYfqYri5agetP2yVs
iexyboVpO4vohu+5NmrJ0IGYjPc9DYidEqAURZh/v57Cr3Bdh/740vTKW1hx
k6E5WcO4/ubwu6a5SnezGhb20xkNAN3QbwTIN4ZZ/RaXoGYI0S6qSdIRXzmD
KLVx6h05oEu9hQqC6fJuMTvlLWh+S+qsGWJxzZ+1dQN6orCCNx/b/Hh6+7lp
3FAvdKvvoREKqetac2+1JgMXKjrKDlQ53SxeZ2XMzxWKpSFfCqsJXH2TNAfE
2F1qXHNKBlGZd3biuUQ3/Y3k3vWX5GCIWGONBZb6RuMuHsNLgwvxR9CoqqOT
5fXm1zh3qU/n+x0avVMTucL560yF3ItHy75TY83WE+RFe714px0WjLqxZ2z7
XSZvnUWhLktItDgV9CsbzzRn7y76X7RvSAC/UehgotbkZmmx6qftIBcDWRzM
jdZ4nXQ2ms0EYRRIUxHZO2S9sg4jBccbotJAD0hl/MGm3IGgYYDddLLy7fYr
926A2hS8Ch7GkoCjdI0RNg57ThT4VMlQ6DCXoCmswQ6ikmBrd/o2kI6ELxMC
1pf/iyw+TxhR6PsqfAeKINDw+JXMKIaDpBW2+NLk4sg4D2DQMgFXjU6wrl9Y
hJqgc4bDgHTwKuWTehjogxvup+6ffgM/6qq0JK/o4qrTabOktRVeRBa3m8ye
K3/UPcvYxRIzfQEQkCYujjFMWmPKLxr5SBRT9SW6+GEH9t8qnnSiUKTjlJvz
lCjoG6+VqTH0DtJpM3zZjMWC39OOHYTuX5eCzyiTGiTVKga/rvuqZMmnPA+H
rmow6pX+S9GJBECwi+okN+gs37SB7LYI4hYliVvHU7a8BDVUc9NME2cPeOaI
8bSe4Pl5qYrfZZyiTTC0jxbFcl1CywbhrQ+tHoK1XwKzY6CJsXX6Q1R1gxCx
hPZ1aHU7SpUI81ZkYt7FhS5CnDG1Hb6pnTvTfrI0PurDuLMjtrYutzsQXOqk
ZZyz3FtY7MeHeMvjfQdK3v85qhCbWjhiFpweTMWORARghqnHiRScGLdhR65R
7OK+1P4UK5jJBiI+5onrsZfK/s+mOwv9/Pq1zX6yC9hpGAmfF2ZyeMM2D+Ri
NQZKiIleMrVnK+hT8KEJKVq4xHiTmqNsG/mEV78L1SN0q2B2c5px7aD2Gpc8
pLfq+wqrfUKclJZ350XEe6zVhuEQ6gXVC/0Gm6kyQX6eLGZervLXI4CwgiE6
vJbsDmf2f0CdV7Aw+WvMrWiYHOXlA2Nx0KpMQQJlHC5ST8+q2BzdM/y6jFqf
zgbhkZE3y4hSexS4Ad1HwMvE+hznkA15d8FR62HI7YgdXXe25sB66VbHdwXK
P+oAnr1vNEguDU4bomAAaevyQgQdytnrOwRLoJdJ1LshZphKTd40IPDKJul2
yn2hGNRv40miBBRO1dcELGUVNFRuu8tErykZwXBCEJzsFvIpQ3IeuTDSLQsK
o/av2+zovHTEfQ7Xp1Dnvf3VoMf0u5v8yKNhL9yZKzyOfsPtQG75nB06mnO2
fbjF4EUeXC6l28rvUlWMIYCCPaStFprkIftfk737zzpoCel31G1azyzghXVC
m+jDSk5bUibWNswcwznDrPDLcxksgCYSSG9EVL5cEqI6oLf86iGjsi2alo6B
k8PkNNICAinqiKY1mC7zvy+tSfTHKFHPjLGsqYerplv0DpvSCbXx3ThdEVJs
KajvxxOadfDntL029ZOJIpJEQM/ku4OmjUhG+YPbpiwc6QzMR1yLEn+9f3UG
31xpRakklRbbzYWyQWyciQWJQAeRXplML6fryUdxZ9VbJ4sjTMqhSSEtOD9m
2agvob9kbdPRjpQ2ZTzJDQrUNrYoR5ypZ+fGKUyjBSLUDCViYZMCVQTwmOce
UaWqbRp4a4ZPL45zBj9jBKCCIpCXe9JOJOVFZRpxsdVCeBwD+3A2ZXNd7t8K
PWwWqi0goatB6fDfw+6FRxKi4PGlh4l0NwQGKH/6W2DALC6L4w6bcuS5TAxd
NUUpW2K00tbw9ocppFx7ahCOES+q5NNpns1ol5MxDKK0hCeTC7zdMQXnLBQ3
NIsyHDsMDrzE8CAAYIbxAWOitfg/Q9UrFc67z1Sc4zVfVuP4IWQXiL3dZ1DA
CXfcwgJ1EMWMsTEunysdWawCZ8BxmjXaTjaepwYr1FeAfU2rw/ZiFR210yAR
3XNoTVsHzknooRmiC+a0BBP4IU2KQEvFoU2YskluGodYQAg+zMeKVqR2iujT
ZEoG1BNdbuc4p+QZ9ZUCJVEk2dAdGXcysSx0WcNlvC4pVhf8BPoolTbsQIHn
2uOFtpKwXfrs6JVbnETvNv4542GkYG4YKNieU0T0n70kPtGJ+08jfU64dR+x
By89X9fvT7X0GybyQ0FIb0sTImIxLn5tj4rKz01S3JwuKXmhr6kLK+4ChWRj
ke6sA3t1H1tHqhIX30HIXUO9oGiZ5gml+81mYAXo+G8DrN6/QfOTKyattWrr
4hvL0dOOpJh8/Iz4P9A+PpV64UsKKFkjNQ0VGtHZfLYzZ7rIDpqBHEhdD5/v
nldqhUGrWDfwU7eFPmd0O055Lvz7lJX2TYt9Oqgj/LbiUvufZ8NjKqKCW/uy
QSIGZgxqoxUKPnxQfGNStAh5fWeZ1LRx2qPf6jmmO6FomtLKJyiLHJRHiqLm
MXkd1f8bochF9OFkGe8n5zEVv3/BXrSFE98ndCzjIa8saZJRTb1cTqEpHO98
snvOrGUVFgu7r7HCFbFR3deOD40bmRxGmA51r0NdfI6QrlulOHA1aUbfIFGT
iEmpHRSBWYMwVqdkhwWLQM/eYcm0Izse310eSlWUdC5+/L+4Wp0XNONOjV4k
2o+2VXVbpxLO0dG5uhi+RQUP8QuUHMko8wiOdl6KcJ7d45R9QZbhaBat2kHt
Rbyq6EqeCN9JFZXSX8aOFffyAEkdAShhmHUhF81Eb/aBrn/UwVyIb1tYHM8u
+ZgE/VZAsHyU3du6NAaraq3cLxOARhi6cHGFzfvcy0t0pM76kkRxOr46gK/3
+RDj72l7hWVSGmVlS/epLyRDc/p9Y1ZAPUhSYT62/bOhGysp9j8pow9g9nbw
wanFIokdL+PiTIjpsREay71foTvf1yGhVOVo9Feao1ViW1qaCvcG15YWgVPT
LTlBEVcwnsUrq+6+7OPUhr1pEodf8Fl7vltvPYR57FOrthgDU7wqdwA+LtIe
VlEctY1JtuVpJlRFN3ra84A7dg8h3FZWFVLClYg7YwA+Nl7yLvPLuyi7XZL6
muG/YhBHfLhXeHUaIaNbdh58jGi8MRG1SbddIqo2JAbx00AHhYmtvMgoaxr6
1zP1O6/Q6zirb7nhLnLAJGja/NwZ/d/jaN/XZKKRd+iy0r4D4KqvUQCuZEo0
/McXfYu0Cjl4S19fyZMPhPvIylLmIeysvK2hN4fxM6ulJWMwEXq6/W1Vgzp+
oIIbkgho6LenK2mTjQfECNZ2QtOE89IvqtSL9bbiWJMMYxrgfeMh8k59qQpD
Q8a4+8hxako8oCyid9YdwcY8pAPYdjKjTjDt97PmCq2OHnk+BZ7U8QTLZkJc
agvnvYpUpWFBz2j3+ApGVWOP+Ik0V5NXSRgu2vYp06LmCQ9P4hWt4pXCr/Mq
GEGQdCaV32TdV06eA4YXqANPzF44csQeXnSNZVrxmTqzsjO3tnPYUdMSHtmW
yk8oB8qfviGSoDBC0sAld47C6TfIrx0hH43gHa0b88sY6ipqSQo7RuZRNOIF
E5X6MBH4ZIwQEl7aUfwe8goZmhtpJ4Re0lYPmELKVXS1PbJLJY67F8FrfIhj
jDbfK7y+U1z1wqJiTamDbaL0JLQRCC2XQ5VnqPrW4UiRMylO3zJSQg5DO8DR
1UhIybqhIdkVTSc2sTigIb4dkCmn14XOBkqm0nBrgD5WFQ6v/n2O+LLgZIWu
ZJVTi5f1UvYM/FWbR4x2K5BHmsKnpJ7f/Hw5Uzu2l550w5IxOp+3iMG2NGwO
qj6w8NzthJt4lO5ajZBWDIrSrG6ZoypwFskeEKzf8dj/i4KRLHfr0qkhgu6R
+r0pRxSkcH61ddl9+uLkhXhxhdXZf2nVk2uhFUoObGdOgoksQM7kaIEqzVaf
s6LNk0HYR5/nt0kSwYa/VY/GgJPOrLijBNA/bnxwCMmUbeFKClFxI+PCuFSJ
H+huyRFhdXaCEFTVwJD3PUaoaL2+crONqjP7ScOSvP3i83SjHike4wmm1WTw
nS9kQMpPRN8i8iMKa4uO40IfnlI5PPNP77HrH28QtCXH8Sjhpw58QyNgAefY
onnQlrnXSD7GUC/4frdx9+lvy1d+S+XqU8jpCOSlrSr+6xZqkjwFBzkwajVp
TImjeUttxxh9PnuI2LR1+dz4ap4IvHkR7fzrW68RcZ/hZk3b3l8z5/jItW3q
ZEabvdo8YR5d7AIsdIsa5SvM2SGTERhBoh/0zbsXDRZKXLgvrn5hgyJzS9xQ
WcmMDb/XCCJGD+uRRkg7jbVQmrCCPzR96az5Boy9qRbd+w30kgQ/h29AhU/T
aYtpOocE/qNktktCndBwW3fAuB2ygkIAEMHHwvf34bH9Zgo0azTGB1fiFXDG
dCsNk/LlR5NBC/RyUeMVgTCH9Vogw2HVdEWZy5iV/6234UvaPAg8pd7F5KyT
nmicyaLuC2/YWlUUI3IW3+BzzsxylLyG+YjUJHI92caKZA9BSV3f5mDsnMWu
x+mKDFavTVfov93mRzizXEzPcCf9gIBrPKPOiuLgy5QhGgmfYtyOtVQN2MKv
MMM6R5WsSJup7FPHPY/UfTX8sGVgmTSIsJPaUMHqjfR3ftEFU8+fk9hNkd5r
TX7TB/1EBB2sU1LwmbDv+XC2WwQk3LSHASPPUPtDngANZfrkgYeyN8t6WXT8
OC/PrWUD6t5NzzaB2zcmC4TdQCEar7pgIPlEWxZp4t5b+R3dkPFk8p4zfsio
3oxk1GKjtXCLVkfevJJsQqSboCLpOdcAWzzu4dmUAOnJoCiD4gV5Xd4QL4Ic
dlAQe1bPs07vb7Nhdd/uWZzIr+c9BaYR1ihycHVY7EihcQD2kA21aKskkrau
5CzlmDPiBA37oSxfJUHswWZ0tkWsV78ttxCHbbdlofDQ49pquew/nRpLzA10
Pl05rZc1382rm3UQ2/+QaZQkoj62jdKQIYk5EwQaLjGpBSHygFyK+oquM9OF
wdN3JlcRYnGzNamx9Za0irgMhsYMnz+yTY4LpB03U2Tzdo+FlvNtuGZMW9t5
peARt7O3mVo30wOVTsCPzeMcsR/gEsHPFKkxEy1e2T+wcWZkIUYEJFeVc3lh
B2O/LsmsCCpRXzvZ7+AP77P0MliZHsN1lpiP6ZywrykkgITnExMPQ5DXIYCm
+hjAGv7Qw9b/3EPB/lnXQAbnUi9wLf1tsNWDs6rS64r2zCsY2JyKqKpIvPv0
ARsFj01VOlba2Ip8EThhlprrliLYr9zHpvGdtLAth6beFdqiyLFNcXZojScz
ESM94/NlkppNfZEb1yUoxdw/wSpGiLCpc0SPIATP59RI8FiGOiMN9nvRoHfO
DCdzfiFwD9zdpSWAKn4Egsqi/NTKvfKEiqN4oVdVZ6CaA/aBSzoPozpvErLN
zPvguel3GhArYdSMcTiBHLYIONExWDxUfexULrv/tMOQJCZjCpE8wOooMnxv
y1SAj90EniY5FQCpngFdhE0QtisX2yrcsviejjG/Wx4Tn84Enf5wwjsEdyh3
2nSTEtb3lRPUznsRvJXjDGonHJmPfVqOMVK2moWWP2jq23XsocwUbNlVnpdR
g/BPBBlIR6stKKKokXXddEMI5q4CiGdA3gxVKXJVAkkUk1U4HdkK009w7zlw
9b46x12XcFruBmQ/qs7kcujqlbORXmPYTmfUjYlFLuFzfi0iCKaIbUN2sbiR
+RjxnhIqXjtgWVoQUmUFLdNAT6EcALjZuNZQNyYQ8bUGVtGnG6CX1/B8qfr4
G82tqfsxFPv7/rsXQ74HgfQ7lvDv7B8xkru0LRGUV9UvhSw97PFqEhM4JxWY
8iEVE/Uz5AqGFO3WHLh0RbHdR2ME+/8jww6FJ9tT3KXfMlb8wqx2BkCSUqPk
JjeDLaCZBrfUFtzEOJS08i0xvvNZLybxHoSLojqKAlmiu3cn1lMAGWrKsCA5
bAdiES3SE+6nueFbbVSuI0ppIcvQVw5t1SsJroFudFGtequk4qPJPYt6Cez8
9xHn1ogVPb/KBMiybgzZ+HHRjJBiNFWrln3CQtQsNp7TeKd1JJBRxPPatiK5
L+lqtNTrriQ6ViUJ2zbD0Ywcs71Ea898DX/zo4gQH6cTamUhbklu7YmVabb6
/5Q3I9IEJ/dasY/mTPYDgMWa/95rMSSZxsu1VBm6p7/c7BZLug2QsBRjPngJ
nsP5dchpnG1LiMTMCRyKaYXJ7uadXQ/l5wJh8shIgxIxWYuvM1O8tA5tAIYf
EF9YKoV9hYA+zi7Ypapt3ev22bGBHPuzsHgwhle6n4VEKlTFH0gxNNun92mA
fsvwvk64E0usUGDopXDUmevhrONFuQRV5L2r0EpjCiYvhNaCMoW9JYM0O8SL
BWF0/VI5FYqZkct0MNpwYQMpotOLfejWjzXYX8SSF3d5BUNhdnW7krAvZCA9
Ce6ERV1DZmWM1omFWu33ynOZV7FABt4JoR1PD9rG0ONm1I3CoRWtqzlCS1P4
Ff6ZKobcRgOdBkGJddnIRMrjWcv6Rd4edZLIuDmEnBf/3P4xndeN2WNUX5Fn
UbqqwtYuqULSxpsk1y1OzXaH6KvOjL4W4oRmrGNmGGOLQxC+GPmdJh2f4xjt
C7wwRky9oanqjl8SrjYj8R/rRiMz+yUWqgnEorPFr5xyhD7p/G47LzaZFFAl
rCphnMl4IzvZ7lntP/eFMTFyLzXOQlW4B1IUmGrx48kewCeMLzCUqvTQpRZ+
gKRYVUKvTBBv16Vtf0JDNNGUipdRUby7+un4qYyxJSdoqlOeJqN6KVCyZVJJ
vYpq473sJAivqHEAwE4eo620SS3eLwOu5w57azlqTV15eaYpAxlOUj0WjNHB
ymOp9IEvU1+rV/iLRTzWczdYIJE87hoPz2PkyWUFa+cyDP8MvGlHmiMHaaET
94LLBpLpEOb4ZPZs1Fh0ehsmjkW0VOLWw92uq1orhgJbL69tXKRsu9RdBDA3
1Et47R0WmGyIZK1vZykFITLsNlaWbwObIMfobmacNqPDVwnByc9OwQnj/B6E
W01IhwWi93HenEBADWcqe0p82XltqZZGju9HeB8zIbLEkephndkQmKAU989k
zGiuneMaMsmYyLrrtJubgdFy3m4QKtPEXACDmNw5BItFxQWW7LNOD5/5+/e+
+uDdTs9fjj7lz7XmFxFg2KirY9I4zH3TJKh58ngn/kGmaNB3qpNWwYsVMVYF
mwF3sFDjRt3qtkIOBnZKcfQlgdl2Sd1w3Mj+jSbtOqGAQDSNOVonOG3tPivg
yojHyab5l2Lui2qCsKjNcCflsHsAi1+FWybvqbnBfJEkmddZohdD3T9fIdgJ
bgvmLu2aMw+9bysVIqENVf25aWj0tml9qhEf3sSvI0M61OwA0Y9DDgblyMmM
uURzhGwUqajg0SBYTgXOujF6s9hcPxcZAl7+OL9QC3XNGh6/ES76GrtDcJje
MxlCXQN/KyHglaIdVWZx/6F3dze0PfpGneVPR+M7xu8N2zMCaoJAwpLNSink
40S/FsT+z0YVTx78x2PbiL1fnu3OHKi5deH195HkT/VXq6CzTs38FMMooqze
kpQL/cUyKSqvgHnxwxa0VnxRS8F6t0eJJW6fmS733iaPGdoWIHQdbCySLdFp
wFb1IK9vz9r/mtWqYxW59EoXDBuEJSVJDQO4aQM6slZJLvcp8Ied9UPdeDXE
XsXDmo1g9MX1L+17KkERi7skpDWO/1OZX/NU9BI72HrYEJ6sHyxsUl36ZzB6
0C2Zt6aKH60bvQZedjUjeaEN8HxiA6OPWTrXpbJvqznw0a1JUKoMve5NUKzs
1g6a7H510a3FJ94GcRf8KJjl4OempKyvPoyJroL3tGXmC8ahiOVxpKaUo4rr
H+GvzzxHCurJ5tLY1yFn9q3fN7rC3znxJTjNS/TCVKuyHyIiARjyAXevrlLD
fXAm0ZEzPyzSDKIkYf9xVylkkuiCeXbQtG9lVvHj7h++5kD/B7jXwrON4ppD
z4pHHe/5LGpDNbBBHIdn1SEajpv9aS9nGWMkJMcxvCYDMTOZvA75K5wQQ6QG
HCf9TfTbylE8jpZitcKP9DEEtXS9QYmuWlHxx0KRqmwyAXOtv/ZtWcmc1Vdd
J92Tp8Sb5hvnn5RmGNVQWWzXoKisuZi8TATPI8IaZkoz9Ws738Hs97Q/8iGO
BKymXDxWqV+xVTOQ5wWhmQ3+kGja4RhRb8uBM/xY927fcZioLO0lD5oF2Xnd
ZvjzOOIswQTn/NmTFeaD4DrVOIxviAHBBPUbEgWI1XUZBHOzEw3Nh1LPOH/i
RqtF3jCD6Yh3l1ivFicvIjUEmy6FKT5JnVusawNHOWoG/B6CO4zvWOEasogj
EHl0NgM/+mRPYAlfm9qgTt3J9/K2GmihbcCo486YnpffGZgn8er2HLCvjMyB
oz71PYI543UDReVW3XX0FxMWSSoT1RnZk/hFYH36sOOs1MGtCqRkXib4pfB+
zrzb5SYzRLj4UkVAW+MJ619/uZ2Iexkkh2BEBOivtXbUCGWgVNMDQMzv3XMO
jpXftjAKNMznwfyc+6MAjw+HM9mKUwRTLOpnIVHJ94yuqiCyu+8rz4DKXL30
pWZMMFcz7XgzlDqiUXKMZEivNMkxbXONdVBYLFQdausW7C1ukMCxy8HntExU
8bh+V/2LNscuvtkGZwmjCyKJEVoT92yXSL1of6E9Ktez79mFWUC7HBDSQUGk
HWUvgrgcQqAEpfgPnuZPnWO4EVHNYdJgPCE27FgMayoQytYH/iIgUsbc8Via
+KvAdHFqADYkQ9Wl5sM0xYyKkT0t+hbEO04Ewcg5AJoO88tm80llPKsucilk
rcwu/BVXtL+Qn1/rz6F+gXNyPz8o5UaOR6rls+GwE/ulqnOWSssnKR6ULbDJ
1v7bjaoeZsNr7QCm0C+AM9QjOiZ2FiriNCHlAzaauq88HDSNBTsmI4cUPvMM
7yUsggxS9xhs70qwuBLeaUr2YA7PxMCrzSP0slhAeOOmVIWhDORmbU57aUDd
kog5l41bLv27Sa3MF1dfMslR+BQ3r2VpjJdX0GkwJRPqt4PEWH/ejuxzE6DR
vqi040BxHMiZvmyfDJ875bMtw9Cf9Kmr+0Ow86TsdtUgnpU3MnML4ud8Adr2
KH6k5vTzXJDekkEAxJfS9LkUQ7BfOxBgdfi8mH+EF1gxmjsKRCijXvYF0lDp
JEshUp8O52ZyRw0hG4WTnWNaYkhOPxWovg/9lnl3Yypj0iUordkdTKPnCLd3
hZcQbv7CBdXxJR4qsbLA0yyeyTZ+wVyih34PvHljJqjvjSwOddclvpJGWlmU
1bcEELcqBAijP7ovLV5yY9+1LPf0CUFdNXRsSnEkSVqrYIMQwYZCLtcCFO8a
plrJ9LS87i0V4YfdsHyuQ6BXUB3eMK49EqV9UtNqm0Pm0gcls/aMtNobj2Gy
gtkw/K/N1sVHwV3JgFq2+VnpJIZLoqY+NPpN4r2vP0mkY/2QvduuGVNJTBNO
dxRqlxuPuE0l8NinVvCI+hie88G4pi5XWssO54Ev+NMn1XTHsmNC562FxlRw
Oyvzc4lyoaQQaB/SRuFkJWLCWSZSwh44J9tz8FVkHIaOL/D8m/76Nl9AqXr8
FOLxjW1NpjQtvzYIoUWmd5h9zRfAlkgtDbadIgLWLhoJb5mCZ/lzpFvmX49l
lflqRP9inzOb5TEb7WT0+zTXOS3meqAZmJjcRmyThWyEseOfeho5mM2n+JkS
8wpTZ4b3XqPZiakawohah5iH7QBbwt3hx7XVxGPhVdzNGh7hYP01UOT48DXN
zCHInmG1DSGKsXvW+Xkcj8Chs4gAHCrK/nLd808dDFrAlNr1ifZtGYhYJsKL
xcJKp6lwDrgbJ0plBJocEsikqv9xyA8dPm6ud1cf/IivgyUohKRbesInHXfO
u8BY3VIm+ZsswYy6+UKL1zqL99Ka/O3vBVlVW+zkHlixuTkminZn3A/ISRlo
+BN0WUh+HTq2mnBHRb7H6G3ydy7oOyteheNJBXFhAcz4FND0KaZ5Oi6R/8Y5
5CZJZWN8EwFGDI/b6Don/dvFiZZmYMHftdWeWxTcrQRGxLduSR9rQaymM9Ry
8RgBvjW9kYyjfogFXPE6wMGBYcpHXLOnLOoPPO4hfGSNV5hvAPJk0sBY13Nt
UArn+S5Aw0w3y6zV4qOoL6G3WqsD5WE6bPtUWfFUx7Npn7Bv7AGQzp7ZzJlw
hS8fpoKMuTW+DKOqYlour/n0qlg2NPbu82aeVEBbdW1Z6ncs3KpdYBj6RXui
ZkfpyCicuQLGfYHEhS4ncbui2fSpatBb5jqyl/KPXpnRLT2f8B0I36IAjPO3
DbJqd/ONn8SzJTeuzR7y8CCTz1wH2d5Eh5bS9KfeEd/IC77ejr8EpAuYHVIX
o3RtNONd1H58jfNFGTyjFUJOUFNMiTlfM/mhb298iKU1MA4mZG1Fvx3LcFfP
UbYspTi4QmNP31KWjGqChOD6WMYM/P+OOrONBFBHWfLDSJX9Dr9cIKd32U8o
ybd5VXDZ3yIH+5wX31lWi048wOBRRJbK/IG5VUxNseJGq9Kt+5YvtT0+6PQ3
8I8/KIojRyeqJ6Zw/CywGSRP8E0oL1UaCq5yuy7UpTuZXf5o2oJakPdMl4PJ
pgces4Cyj0fnrHtk0+YXc28hvIWJ0oqHiE4zrSSfOLSVsIEhBZRNv72tagSb
MPxEipudkDJhTVdeN145VvIb5aUr7j23B1HH4DidWuWPl4KGZgL2Svn3xz0Y
go3cFMqwf/jcuRMZdehbDit7cIUFuwJosZEt/FM8r7DSbLEPf+SPTPeRPCDV
miyOm4JtIkmQkdgnx6y1Y4DmW1xrKeHfBk8XP77BMh8fCqFfPK1o5ftY/KVc
x+oaW+9IrG6+M7sgjfk3sRH3AWK2BYLXWkIb7CdRGh5YkTpdHvkRnM0l5Rsq
kVeLGi1ExV30wwVYfDDkOIoHPfmvkhrILqIZjBMnaN6VP5y0iqdX+2QDjKYW
NN4oyxEvSACK5C+0H4aoHmFr1vyTkfrDUg6c761EsxVEj5M53AXcUF/MKg2L
U22GHs4zm99CeO6bHsn8DXZadX3cCvd9U+pPncJd92a3ZPeySr1/sNKZdqvu
JN/QXP2PZ0mqGgJZuK4ho7CX13dRGAorrlrV1ylGWeZ1yCbDrJ+K1KdWkl7w
bNLRSmAvbu7GQalp0U7rId4HJTs7ANWiMc+ubvzCmhxK74BdCaXAEXxXgdRQ
8t7F57CoWXxJBMDjR0oSLj3EjLF3co8Hp5oWrC1QP5vN+VeH0Y4ziIzhwTbh
xx07B56R/f07tGx5iOk9lP17CUxMaF3gGZeSRMHXAUwgcFRbQqrRV6G9B7Zy
2UBgZwh/omGt+QmC1hQEQGCQZru0z3AUc7xhQQv15ClSUBJZ14eICiIjtC50
s7U99H7WsohE8yJ8m+QKZRzBz25AbISZqv1t2aPY11lgFiC9raFxZ1zzH2eG
ZIMO3AFPKDvJC17qYv4z3KG2sS8owAMDwpgWoBaY6+y7C+oZCTs2WoR37q+0
WYNIIvIPpWqUOG39FKmfew3aDBqtTnnk86sh9VIfAM+vNXzYKBMg931DF2c7
+Hi0nxkGTcJje6dzsB908HwcJe26je3a1srcBTm2zL/q+geuwSbnNs3XSzkc
W6o28gJ0t8li8PqLm+0NiqtQSU/kU0jiGkgd13u2PMzXNWp6qkheN99MjPkz
YhSaTc5rNYLUrbU18G8yViuLZi6OBOuLzdiGD3Ed21sR8Cp6GwXJpr+irWrF
nu2pVvtX18PdyZIP8vUeQI3kW/CULMXvnJvYwLTzBA1pzhDY+FdUweeeQ6Rx
a/xSxEyjROpU7+WxxeoRClK4HZZshSiy9Z04FyZTWYFaF4s6YnqT7FsQBRx6
XMnKYvqjHAGOkzys51Vf+B7J+nQuwx6tAvyl3Qs18lLowmCfDTVGv0xlHrE+
vbPLCtL7hgq4avqC20laxH7DBoiEQ2kzg8H+lUETgNFrQ3hERp69fR/9h7jX
6gL61PhYY5Zj8kKCwbumf7Uzn0rITmG3DfowHOEAVPvOoNMCscj6f3w8URmQ
w/X4BFLx6W6U0Apz+OM3qbSjwgof/6S8XGC/iL6IhcVbF5ih1XpXkFYwRkol
3HGouNsAtePiS1M6yWUSwBS6roPbXc6xUazPvmBVDtI5mhhG8btC+s/vC4L1
hS1u6cMpKlk0uN1vOvZl/iqN41x8uayZ+ZZAu73MM9r3qiGhbuj3p2wklfU4
vzmrDmIs1INxVlyP9TrYgo9Csjj9HYrHw8JLZNC+CX4xGvRVDsa2gsw1bVwr
i1aaNRcFeK84y7LkF6VQcSthvFQOa9N69LJcSMSWCysYlbHYAU4KMQFd7+i7
ymXKU2KFtzjTje4XfFSYyUNVd+iAYCOVMznXdfivQla89TVcoN7p2+rvbgiV
tH7aZlCP7OaQslmZiB0ebjOJScIZI7qGA6UfANmi1v0SR5ysjsD663bZ6tQD
cVw2RdiCohahxssel7PUpdJoebmC86K3mwluOsQ2oN1fJtCbI1rCc/Yn3fcD
58YR+mnB1XGcS4He1FgGX5WB1w/sPHJoQuotJCkKrQxu+mMj7eOpMiEjLFHg
ZKHnBw9lluSyr3NgRvYUmIKHpBk0ymInUpWyt6EBQwU1p7vNpSUPAyqDBhzx
lXl6WfQFptiMBKodCekyy4ueQGX8HHIfpOjoSU1e1kFw2mUsShZ4C/8TRRL6
+0B7rNuuTi9lT1nA21lREcbuShL6UKjnDE6WEtWV6m9VBe7obS+lIl/+u7+c
xIvo+rSdEMBhJgfnLPNuZ7+LabEZKBD3ffvhmLKducB9UP6eqk5tLGlCnEkE
IFd60VzQF7O4V2fqPTeQ3RDM3WvyVVr8isFMjg7ysJMwhNYuXPhikqg5WMrO
pyy7NWPFZdr84p8Wtaq893cC6zDgdXZGf9keUd3QQwv9yB04AFIsm/heJZ9J
hgLjxtxNSLki4S/4un5qDRqaxSo0udy3XvS0LKqKLr/0SU1hsXQt/BgRcKAi
I9t5HYYowvRymqxa3sCxinL1JYCI7ilHORRXL2VI1GxqLZd3dY/83EqHIjRV
8xCKp13E6qdz3i3DHEipWTG56N/gqdQzqMysaiqer539GOLBfSuUIAJmXM8w
alVEPgvxuaoDSnckaTQYdp+rbRN6fb0V4ALSemr6q/VqO1zhVjRXPzb7IeNT
tlly5NwFKlYZ5K8PXtITXzfOy43sfUb3zN4K7GONdLxbRvZclijOIv2bB23S
GdfeSJIdL9pQ3LUh/hAZkjGp3+niDk43NmMo4wapJ9LPFKi13nRKQGANHZkm
8IownUYcLzuDofhzeYTrfJqXas4RDL1ZMLAB93lXWlJndkrt/F3Jkzoo2MmG
Td0AWtxpGkFRg87Yuj/zMa4QVdCTdhcKR2C5r8gROAmNQfQR+XFA/scBURrz
yXiJEoZ61V5DKXh0EsIPjZsRBQDT34vBtuB4jQtESNnv/vFhOoXEKcamLNHJ
la9LkLNGmr1Gj5Djsy5EA57jg2gXhJNV6/v9d/9k4rw11T43VAWjp6cxRcID
+944hZl0sw6cPYjCMNxAWbFHLxsaGIIMGNdJFv5ka6N0vVxWTcWd5Jtz4FTC
0xHKKjI/UnQfFDI1R1U5lAdpvv/ed1JluPXe7XhCPBnjr0mWqJP3Z7s5k760
qyPv931dGQhp4K4udUMYWnNr1BqKKvYE7Ay98v1YH03LluWQFR++XMCAkLq8
mbYOO35BhrnIsMVBQ8Tij+EGtaMaMCyyLpu9RKXNNi5petlAUTi9r0E12fKi
l6nlbZZq8swENIHXR3tLBRQzHzElDfwBb87A5pdcyozEGF4RExRpMVrm2XiJ
NL0l1CGEgsL3KL4n+7L0D5OpyU+cl2g2vsfyiWPRXmXqbwIkQoKdynjoIuKi
K3tS5jVsWGKDGEdwOkXojL3VJjc1jaHhuhZpmOV3+Vwof4waikcFSS93mtVM
TFUHRM/UmtXbY77mBzbC0zOpPZcxXBjkdg1hTcft9jJaC/7BT00+bP7lyv45
WYV7nA69zSvxlwpxHFLUg+frAIoj6ilBtjCuMJMp2SEdnVUYaBPdISqc6B87
KGfSKutdK3MjKug0H1KW3fO6RHahCjLLTEEh2uX6YFOezyqV/DxuHoqFWw2b
L3p+SocIJ+54ONLkfpotqMnRBTD9qFnkrg4Dd7Eu1f/vC2TvvMpBmudVfl1B
uSryalANmrbGNQVHj6UjcyB2DU5aqPDbhT8/q32JBNp7kqDhZofLm9BI/n+0
mDA7rDW1wkmowOn6we626SD63Yo8doqTY9YzmIbLetQJ5UxplEDVWSsclhiY
puc/RZc0EFhPYEhFO8CXN9sIj072Jan3pSOYg0bgGf0tkisKY2m13g59nKgc
HInoh3QBOu4QNVOw1IRDBpxRAz3Xlct3i9hjpuoowD0NQXK3GdLoLmIqe/L6
aUwrNga2ABonNxBxRdpwkHPCP6ot1nHjTup8lejsQ5ih21WYSKyBGrtSS04X
+pKvnTIW+4lA2Z6UFj8WbgoniXXATpHHz/SXflKwPe9m8VxPSX6GHdRsUiof
ugDVE93ytHIuWQLaGLKXd/QFcp7594iU7QSnZiXzwwwGZSNhXpAJcU7N0gjs
S48XFUCrdpuci8Txb7OqouVl/yrELXcvRwSHtCVCixi20uhkNHBIGTlYAm1f
3Y9vgyzTkBiqxz9SYIJPZLXMwleHUfIB1VQHYS49fKUa+elOYwA4Gc6Bcrt+
6epTf5rbYGv1v/j28+McEjvG0KLwwrDHmebbI9zJQDbDCzvkM+Mcxeae4/zH
XHkX3EIO+tzb1VugRtEKk0OTW0V2FX+3sTZryiou6cX97PC2efTYPF/FeFdk
UpPV5YohtoVdXBDJkFBNUCvhlQdTZF7/VuHOu7zGQL5B1agx9oHPl14zM2BY
s7FEpoFosbo1f0yjAzmOxcCwAsmObNMyVIVPvZ5GSvzdgmVU9qP6z7N22URf
CrXCk6mVwh8a+TDO8Y6wkVvnh7MLYfLkvfAu3Pzc9ijJ9NeOfnkLO+OT0hw0
vExvODZgwxNvbaZncs0baTk72t7F1HVK3tkm2HCUipenjTyCIVrlzKWyYU4l
DMjdZUCoKkBIIRwNDdVs+Tdb27UV2gXS2pQg2MiHWcVEQ8PCEav8jvUmrM0w
F6jfKe7fkW6KWR2qzXUfoKAfEe7LvtApxnws927BPZGdP6geDLqonO7tfLVR
f6CQ1c5yq46ZqKgFMGOeGturLZmuRkjdV/5yPZIibbzj32CrdN8WXmTDBxhz
/jur5BvAjo+jTu6wVMgo6VniXms/IbIXvCzLq0OpIaveAIoG1d/Sfl5835fh
S4+5dsS8wPpgSss6XN8YvHvSJgkR6905HDkrO9GamEOiBl0xmq2O6BtztgMo
dmK6+fsTj/MnQ0N0hRIBh/YRjO2TKdvjH5MXgzXTazPuX3FcoOpab6OVJ1Sv
L38cd0EbC75BveXBKlUEDRr/Fn8FlbbSkrVsXSYHEIZS7jQz4MWitDh6ogVl
y0r4FWWQundQBUkeM0PK7+5lRaVJZUvEsrz994/KQOxRV3aMP676L3mZQPwt
a2/kO6Y5OKwYkF9sLNlg883jaDfqHoZ6ELkQd/E4H8KI25p9TSdoh+c1JiZa
SWfm+qNdER4lTHIzMzVWD6cLEmWKtC+5nvc5HkaeN18vil+djpvp6gt8sgNX
z6p/jaUCZVykHbWz

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpeg22wq+Eo1UxHW/QaD9thBXx/09VPqcSnUcrzsUp76bQCAR6nW2XG0cy+yssO4JTgFr8QiINHYa02FuW87cTxn3OTIrxs2yaaCT54m8EX5Pxvv5to5XBfnS5nyllqcFo12QJ8gNBvWXZmWCl3skfxVMf5sFNZ+yLNI76srFPbmQ1UCHzQ6dSlKtbrAYCUK2thnt2N7FogCXctVZ+UTO8CPdCEyxw9+uNb4vokS/1HnhK8OzMygnXufMbkXXLU4D8KJoM3kh0/ksDgb10/a6efZRL/sk4bhFwxy2MQ/LjrowCYAkm5I0sjs5YrGbdbTiqP3e05iV5vBB/48+MjRSn52N/Kgyd/7UZSJMssgLIQN+1dvk9jWtQoM7za70eBTL7VI+pY6UecBZYNweC02AdiYT+Y27PirrBMdovlPjXP4Wit5Mc+PSuQzg7LelJwRjjxe1v9/YR5kNMP0iCdW69/Lfo6lyJmufyk4U10NfIoEqDpu0dTiY5Cd41iMMTZJPzHhOyC56PEtG/jTLFRGy1t6Bv1Wxrs7i7vDQODJkFLBuNGr3W/wQlQPhj95v53/11aJJeCNLFLj8qDUWf4C6Gw60CzOcUaCrBosXjyhX4U+s9GaGU6QQz2aZXqQDJWYuMZ+9aBS52lVNDQZpCrJVDZzbDJcbIM74AAgsZhgki6DZND0X6obv/BY7NFS51kMLLkkze6Ktn0yVNWlvfMweHmYXdKc5QEkqTAnlL4kTXL5WY6/TgveaOvppUj3smygGj4WPd1h7OY2YCOpGA4bbXvwf"
`endif