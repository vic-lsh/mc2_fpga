// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JrqItglmhwaezNFHbB0jyxArWb7FaEEAzqWxD13CT4eujakiSBBSLZXNcqdu
RvnSnCugAEAPrGDkKKNV8yC9bQIY7C7SMawOqRql32Ei+t2rdTkxciwEmMKp
OO1xKHVYtLrk15PRrNo3qFbLnTC5onDo8T2nuAc7RvySgGe4Jb8Fvj3R/OuO
OVxWCmICSGxPpkw7p1agC4S3WkRSzq1vodTY73IBz/a1ClSIpAf/cQcNKnbk
LSJoi7RUaa0VdJifGDkHdq1D1MccRJL+e4PmRVWol1hS5P3MJUxHOTJylcje
7FIcAFOvD+d8L+c8PEcOLgAZzO/0EVPInmD6WMlatw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kxQ3xaDoCw040npbrjFC6rSnrC8QeLh39iEKJ0brb4oIDW2bxWrF+xAHZeZb
bltQGvhzCs+uZNpRsOxtdjL3l+c6qYa3j9Bc03IoSfPku3HNmutKz35peVff
AAvnXMSuimnsFu8EjHlfaF72rezQOpRTvSyJiQJaW3VhhE9yLMcglDqyAh2a
QeDhUiar2Pgt6W2Zlt9hsDQiMkJExCghwGSZZBD+V8r5+DvjjoD+FEIpwzhu
NzSQmOjKOKBkLupKMuTOU6j+t6xMGRoMih29R5vysVXfwZ/DZgTcVTTKyfPY
re7hSrKGV0Mav78g1/WxUUsdk+KXDAiYbNlWMfOWhA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LMAYLDRad7xsG3EUwCqrFchzB62EtL4wAe6JmaAW+7jxbfP87bdgE2NcbgRZ
V+TVfcWNjClBX+IBZkrt5xA3qypU3oCR+PInJFGhWkE5SVtNxf9R/c4da4Nu
Bzg7NHOE72Zcpk4mwRlw1mkg4Zv0rPTGPQpBGfaaWsJDpZYMXiY+Dc7wF2FX
fgBUVOHklOj1FUh6GjIfqeIB2ZY6nMXwcZdtHMAha7sl4i3x/5VaMIt8x1wv
7PJdRye3OSgZvwTmRBnNq1Itn09+qhvsTnU2pBOW1xBLI34fK+WM+K0IBtuD
LbqvHJ3pSpR2U7982fiQf48FmaqFDjeybtw9PsK0Zw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
diEfM2U8Ai0L0bx9hLMfMuMWzunw5V0s5zs8M8BGJFMEhAgJvWKJNPmSIKE1
sa7d1cKs9KeNmp5tR4Oirhr5GBBmyAgBgwiVeLAqf/ZTjIxfDvCUeZ/jzXWx
qY+qoPFmus6SAAgX357wew6O3jncg4gH8gx35hPZFuPRMgraiUFKWeV+qrnO
1wqT5wcUhKNkPwf0ofghcXg1PmburgTsjdb0ABRDJvkJP0Ex//athXVSJ0A2
zMOdKDcqQRulXXoO9mExfM7nt8c7NPrPkbm+mTdj468XpuUlnBTwa2peUGgf
B0kOrC9mL/NvgRt//gYtYAiffa964LDduAsobhPcxg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ovFAnZpRhd9bY+YgW8x2Isx7uqTOSOLdUE/NuFLSS/BZN8PF08Qlg+2p1Fof
uPMquWPOpzn6nui/fYN3IfnhqYz7W0uVpTWrW19KD/eP9RcbLM9kUM3TgAKs
3vXkttIKFdHCaoCjbbvTXUSzj6C/ikOwe6GAD1NKU7hK296a/h4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bze74+bg63h5BNPHGdjuU9LcPwU4WVSIfxGChHAsm8/Z8eGm5stnFpaWE7wn
RtgtQk8GbAiVtI8h8Rdcy58NluDF607ucmg0L6NgNBgNerjoe/wcJhkEwSfd
BmaJr250v1w41nJu5LQCpqyIyUH/JiYyKegCSQ4nBqF11lKMW7Nx/7kS1PQE
gQVZ++qIMMZ4l3+KKq922REZ2Cvh4E64G/iY6kwKVLFZpoBvID51YytIun3Q
Hl8DZH91e7lRQkKGzsnXdVWQXxCiIxFh2wshngjp3/WJtfuAwmwdlX5//DmA
jlvyulXQTmEVb++W3DMQJPb4nIgqBsHfZDQ6bo8WdgyM6Q+0JKaDRINkHpYJ
19Xplv/5Ldk+nYVGlsvNMoXdUjsi8c5HWUbm3kFJ0gJUW5ZokaP7mUvq49aH
2q/51q54Qh5S8KmzlKOu7eatfjTNltb8ReG3ouumdGg6QNE1ssRAkVL1EUtp
gbyorel2Jhx621OAiTWypoRaVcP88PdR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BPEN4o3uvEKKygPfciGl/ONne7nbvdLY9ugL5lehn8j9WnFesu7DEwGXKsHf
TPvsZj/ENPUuPIXHEnws5gZCbsj1MsksVCD1zucv+tUFgL9y4XHcvhpXWCzG
qt3kuRj+oyxpv0yKInIjQuF/fPa4CM7b28bCzaRJ6OSNzxBdhEY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I6wc4MJ1rNmMxNstN8EJF58G9Wqax41z4NL6ZkOVAbvUja1ZLfZIwG+FWE63
JPaR7/Wo7TL94lWAmtnqg/JYojeUtpkiS8g79AQ1exZKLoEvJF9SakVlJqwQ
kJJSEthcPDzCZSggvVIRB+rJM4HM3MDNcyaMS2KvYGVCoQhQhp0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4736)
`pragma protect data_block
K3plrVYKVLanTe/cSdinWFGyXVa7rRX26j52TGpXNTcn25BTEvcoOOIWwz2Z
Ig7ErKX218fNM/xkLIByNi4lPHPAfXaG3uranec+AIPnNmgUVo4+pRRZFel9
LLPeB/MPvMZV1kJ42kNpH7CsyyFxBrm0F6+g2XrBIjUhk1kgN5i3Iiyh841F
/OjHda74IFq4WQMA/O3mB4LsJUlUgEvu+GI9Ef0MEAT/uVUj7LHHLON4Kcv8
2bgeM+1+u/QSQhZGROuRHbZgS4chsdEglL0dAZCsiN4brFBKuN8Tz3ZGmbIu
1oPxUBAvjyE6jq9748ERT8Mq2fx+pqUYH/+pVXAZiCNkGPloYYTMkdbDoXcz
qze1awOloch1qytYJ3aOp1S07JZrRrDmmFIRBo1F0Mdvt/M+XcjDUSAYrini
yUlqRNu2EtSsmi9RgjERG2/NAbjUEiIatzOd0AavbGyv13+Bou3ZOoxLI1qi
mp4xV9rxPUTDKeV3Q3AGk5X7+W6gzXu8rJfF4GM607SJigYydTbX/cZFhaVt
NO5SNLhxF6tv3VhFhSTGCEAuvvSk6XyyEcwrtfgF6m2ToP+Mmlzxy/iroxHh
pkbtV0u+88Dy9IXphhWeZHfLjfZ4zkn+b4IvXz/OEVGP4DP7qMpKtT6D2EUJ
fRJaAjpcayJTMtQEnoPtI5zuoi8w62ZYWaVhE6Pzv02jUTXZPDgo+lQKcnxL
vlaAxDfTYNSj3wVUBEdh0tsKsDE4OTwBl/qHDHoAaeW1yUPe3la9LRFPNdZj
thb4BMfIO99hFlF2V2yQ/6JngW9aY5hfq7YqD+SE7m8NTm58njGnioMCi2Cf
MW9c43qcket2Y3o3md+NLPpA8V8/VJIwSbwNkkUvupwm/wkjY0CexuXAYTHy
lrH+xk2QX+ce13lgbqnH2wYih92SSirWksFSTt+G4Mq/GondZyQpu47Tr2Ov
LXgrsPc/tBSg7sEzzCO2Phv7bm8AHd/8anzAwBFO+bxvSz1dlkZokjLgQatD
Fd0fpuH50Exi6UYksXntHX1Cobu6jJAyoa99OJJy2wZMOZ+C6lZNqpnu7aKD
iHikDPBWT5Mj6mjvKpF0mt6RNeTdVxv0czpHDsTyxjyF71ugm4WydV2HBDde
I8LjxIJMD3yzqCWm4GciDrcwQ4xyWAWEOMlJGFOE/nZQ4Oq9atXOj8bUgR3X
tl9P+BsEyFJe9epO3EEmIpuRc1gCNKiAo6A3eGHjQrU6CktpvWt2c6Ah1bmT
Wr8+WLvVNwt/AD+W22DJZe0FgphLfEPXUu4D/9UDCSLaqRECWYC5WBG6xWdb
xBnd9om3nUhNdzy3R39QKWhkDIko9ITWxcVO14vJ2sPWXS8QEHF9MTQfbF1r
8NoGGxPnUoC69RJAGKpxlj+hEOZGY1c7OSmZG+Xw1LHa0OUVrFFzgyTT5sqh
sL/MoqYooNNZrAGExvyuqmgAFf7JTA+jDG0FYnLalnYsQvZwp3+lXkwuWRGA
Lp+E05DSkeY/BWNOZFpAfOIaGwI1CkIkeueTrGaGPTZzgLJl5mwsblDnhHg1
dBErwSuJDG4Ua63xvxxSb/ViMu7+AOM2eR6lakx9V1EqpS3IJQQQXdAmOGMG
kWAvlMn8kWF7BJiaE3TZxwBef5Ed5FR3NS/psW7Ei8Br8jWymhUkU1Qs5Jhf
NhkVoAPBxfvLfZABWq6/6pdD4MMOWayOKcf92xQPRgCNJU+r1IrK1wTSPfgx
xlApkXrTfVbUtX9xlU2EGivxrZXqPg9Vqjk0wuUjaGrpMuMT6W8UMCGDjgxL
T4MtnsqED8TG+jFmQy3cSJC7TvpeRW+pPCaj8oaiJlOzzduleDF27FdbOzXV
1uVOGZ6fSd/3lZlGfds1WS7R6kVZQKUIZGluAmNDUDZNpNA5PwHJ7H68WTUE
7trpowmH5YsSApEDVPxs5drk9NmDzAsJCB/pRH82SNezxBaMkMJcoLJmfdfO
Ef+NhY3/IcoSO22aTAO7egNDyNh7Lys4DzL0kmN/zBtZ6blniSapO9LNjXsR
lJiLpe5aI2ISqNGPTFXS+gbCJKjpwIHCVrG+ZAeu/aVIW6JqRMZ/JK1/qk74
jnvy/8ZpJ5pusnt8hviggSS5qFx98FwA6V1d5EXCFEu3Pk2h2MnIC0rvWJLH
g9wid6Mbja59J0bpDY38C6poYdl0+veS4gv3IZ82cEeh8a3Q6mPSK82m4Lwv
dofuQpuGZ7WyUDJazgMNESmgevNpFEKihQgRWTaG9qVbFuh3RML6SOG+smGC
sIqivDlWlivrX0AhAJRqFjeDEN3ZVfO2diKhlGzJxsctO9C1Q6LUjhW6LBp9
KH4G0+jQcCxwu4f5J6gzG89ETrWrKKUZqn74kO7di9jymCwSBnfR0b95XkGq
YiYSKzuxLXOuuXPVyt2/S+/b9S0P9rzKv3bR6Si6THep7wJazJmico/eR4Lu
tW6rqzo1pyCRXGTLQdT/wsY32Cz5GVHvW2wffl/u86XbdFFi1WiEcuKRZgTA
xEOp0TMPe/Zm+F62rnmEfEBd2iVmUCcyutEwJ5sb/d4AUgfwr73j9Pye8zEx
g7xXZ3Y0/2tnYSsB5mk25R0vUgO63ZRhZ3m+0m9dtkEot5jCfdLUkou+FjXL
hqs5scrz0iTU1GtMePcHQXqFPtW/DG55aPR02wpmbod7r2ZAFtaHXi1IxUx2
MtaSnxG7dG6MGzsrHGWKKfe8Fqs5IMBNz4ERug8143aV5z2sLZ/TzAWWv11F
dPIHx4WQsdyp4ExoCOCEPbI81lvTpX4qQ+9xFgq6EzzGjCO/QQGVpzPAi9NO
LM0iJfhJtAAUuiKui9voD9rT1/WRJ0iYxsZdW8fKAcTFPiC47/DmyIEymZ4m
cgr/rwKkLDj6K4iiNM+jbYs0S0PN1R0ooY549KiNPTc+P9ut+snXh8oRfovM
z/+IELoRLEJjope5zowbJ51GW37Tb9qZy05i+5rSmBeYo23PIJzeEfNwsBfd
tOGZurilABj5FloVgvdSl9bQYKClayR7rKhfm4GAF2rK7ioTjRy7jSpY4p/s
LbalfZ7X1pLMyFSOO84SFB3zTaeJYYmCzU60lyH7GT1zsF8o75XYp3iILhf+
ekKR8gyFuP1iSC4rc9ZWqeqtMXgo2d+kmkfKivUssQE7BNaH7KSh0FwXQghZ
uCKTUllmBPZreNHsTv/k3TbqyFbW46mfKUaJjPlq756xh5DDgshkwXNswexQ
MOaPhA0T+CuKJeXRzMBZZO7DqOnTaorxx36gRsmw3IgmKciHq+5B3o6Md4lh
8q1XpKlxXgEwDd1m/14iRhePeVG2g3q1FsuS7P5daDtTxCU4k564Pu7HKfKZ
TRe2iIi6iIy4gp0bIe58PM4AklBU4mAvy5Rg3NhOOA8UMhbpMJqQ2ZilZ9Sc
0HKl9VHp7YObNcPt4S34vwfTqFY5jeM4xP6KATmUk9IBflxZzipUHiobqGEl
wQALGjxajZMaqmZbsXd3dN+CYbDRGtXkl2NXZTovZrDuIRkxfUnZgAtxWlUR
naVBnIynkMy6nitDxKEwFy2mxK/B7ByMjL8MXwxocZS5ILsBqBvgqoZ0OPn8
mhTs/U2hY+9zouxRYyyB/hNdZkKYFT+WEkf0iAooV0w/+blr91rEDZawVWff
gvbc0qt4YNrtfbFlhxjHA54j4MCu1a081WLL2T3bj0mmF/hcwwXqQ2jFRvMg
3EUcnekzANbKAl7SwJScCQ5pmiJBD4XnmNfw4j/vWkP+eqFGCQxWRYinJ/mi
QKAsZv+8QfZEje+2d1evyfyQiCrk4MkbSbJlbIuV/SezJOJTpirAgsHO97OB
/l7Xe/tZsV0uPhK3JbetNNqD9LGQRdzpmhz2U+//zi9SjYOLXaaV091or9LV
7bZvjK0adErQVucCdnU1H20g45Zr5Pe5UzlibrQgS7BvvUUPn7cO88a5q7gG
kpOxbOPE/fyOo9RlwfN5fr980pABeZ2o2bFVHRSY2vYZZVOzAwtvJki5I3JC
RBJb0vfO/jhSk919Tv0WRsG50HKyAfVvxMhzzlXGe6iGqagq7mrB8qxEq2DE
srYmRBpcaxKUPtx7S5zbGbZjJtkw7o4cmnYyPku3YSvm/O2x+3SNygCoBs80
UqCBwXCWzLAz26iJs8Cn0rQ1wiNW6tb9wD/iWFXYSjXOG+r8TWv/jkVPamsl
jXwRL/tJ5LYOFo7bmGCYG88ck0rUcWItlrKUbhseqzK1uM0c9ZRDkRrDA605
tCjuv8zeU0uGkQmrc6wizE9K3+xyfE+EQElbYskZG4EyNxSf4BdWTV36tkKa
CLkanAL4Uxc8fyhJsKNoZV7INXbb+N25xUkn8lXYaEpjjbOqPNJ88azGYKCl
bqE3o+pzxeW6Wtwkh/rJK8MPeon6Y08OwfjwEiWNa5U6AppBNoGEQwF8LdkF
FEt4Vf5/1DMqA9Mq711t/AazLUmdVLA0MqBf+gsm4SrNrgLbsS/dEO3A0oJA
hMRlVik/ihowE7N6SALf1ga/pNe4TY4fiWx9z1l7Ob8vD9bBg9Mh6ZiwhNTz
f8tX3FYdGeB4N5iRWNYR5X0rTuqgI1ZTOjTp//mw5F5cyu6ptRti2UMOcYiE
yH9swNVjTa2wxbXTStD0LDpICQbr3cWsNwhVx9WC0JYBNwIx+JOx3EYk7Wjs
xoy2LYD/EExcH0zi+8de/fgbhnhGOHvxkOcgWEDm0VmIiIep40wftCd96GmX
IcwacU5KlLHFSrIeDoXVRtbFA4Ha672RdtnYqJudkBCU+JLyY9lBmKd1f/bs
zdQKgiYdutqhRcBYRrsDtwmm7PJ5Nq7h0Hvh7BZGM6liuBxc3ucJflWGWuHz
U3UNEIPD/KvmfW2GoDBiAZzZivRnfz2eDPKO02Zwqn52fL2R9Y2dXEDRQgRc
q5oxEt2voO+cqldjk7/h0yUOHykYoWTtCJJgg4fpAJA0aO6rZoMIZcBUlMdR
4lVQi58PyQqtEy+KNHrdeD0w8U+ETlWalA9UE5bg4VpSMCPYyK8E8KOMAUG/
/VqWnp/liBNv1ieHlQVpdHSaOCFE2s39VVYlJlNx35qkqaMipT/j78qjkEK/
sjQIJWtxlbDJwTfxRMhytnrndEjyWei18GuOg6KUh771qSg81lL3qwZVKD0e
7Z0abnuAFK6zIhWfyR/jOawFm6dHMaWfFWBiaOuean73FJe7lA7V6XR8Hr2x
exhOv0PyG9a9P2McVo2wzjh8LtS3Qd6dWnchBOtY73OnOQBo1acrDOHPOXEn
U1/nzRbrKJKyUtXJxx7qIB8hgXR5f/DkRXrcy31dqJWTEbA4R5MJrzaRZPqE
WWmPRkgOkm0lQIZyypscToqnKzo84f7SJxRB0EjZheIKOCy8RQ8mSHmbY9Ss
67rKLPFF7onhd0xvpl4l9uZ9zxGbWz0bD2bOe8HkzIN+y9JZhH3AHOq4XmM/
09oxD1v+oEE/wsh5eytm3lpN3nNJDCakMEDSHlkKlqH7VGsYJDzw7KAC4yaw
Qmmq7DLy+XfY0OXcYGN7c7hrBVTENMp/RA+qaR31H+J0jFvzypIJ6Lj+DuV8
QM2s7EtrP/1ZQPb+T5pXNtVEhWFjovIr+3OMf4QuisZ3YFKnbNELqRxxafV2
u12WD9Sj/RmbXME9eh+pvIScKmQbjb8pYd3gWsH/A3/GUKJXAcU9FdF468X9
mhCRFxg3bOhA1VU4Wc9/UfxXZb3bT7JWrLZ97ITHIkdczFn46+PwGlIRAcgw
tr2LUz0e/TbK+pBcT5FdfRM6WLUnAN9SDB77a19OFRXXy4ZWENxbr7uU9rxT
I3OXfURwOsNYSkZCoYFbj6bESe9ZFe8rNGGm1Q5F19Rty3eaC0faY3THDXFn
QQAlKrdIz/mrqWEko1LLaAn3Sw7Qkwx43D3NKLbNsXwzu1o4Kxzqe7BO1Oj2
S2GjJOuNb+z9CMaFlkOTOYuhSpchJjQ/IOXX4eh1IzspUso1pxve9MLtSkhH
9x0n6gBkklfKvU2yiZYGoXSXKOkaRYTdlDjJtYAI7YahzGRUJLKH/k+rfQ38
S8yg29bceFySguzukjm/sptKYt2slOzSxl1nJ3i96m6FQY1DEb9z9J6x6i3F
GWDI055r75UcXlVOASxDgTCSzFTJbUCIQy+bSo72a6rmVUzOscD34wPeyl9k
XyDjsfeR7QD8V1sD2C8/C3NJ5keXsBjkxGcHMM+wQNia0F1pr60bNnyaBsZP
dvManJdGMAnXenXs5S764ctySW92tZHDde2ix0Y7DDfGCxFtP54F169Jjwdk
Q0WfQ7t2Byhf6QA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eq66xC237TMcwpZFF6IQJ1LwMH17NefY2TcjGxjlvGiMAWE9OvDzZDkpZ9XOx414Mq/CbcbLc84U3lt6Syc11TwvKTXaIZL+GY3l1rrttse1MaV1o5jd0ZDGE4ni2DGaE3fI9TK675Wjq8+jqCz4OYY0cGEwHCrbFgyOpmBWeMVxW/kFMpEHuuibs6S9E9f+F7hJJAmEaQK/jpfpD0uZJPVUO1X6ODjIyIjNEXDCj+pC1vufWTHQzyrCyA9IP89UhxCJmkYZi0vYo1nwVaP+CavrsDIUBeFYJouJuGpz/7xxc4C1ZpU1sH6iiiGW86A7CoQtwUYf60e75BDzqTRxMRkw8OFkLdMN09YkTcuk+B1a5Azs3h8bVaj4S3aV6jnwGJFtVcPr6WkdVD0oeys+dLBd+sjktQURyft+9YdMapDxP93WHfMs6DIN2Zc5AV7xijeojvE9n6fGlbTuV2OPiTqgX+fOIEa1RC+ERdrFlrKaXT4xXjcf458JIR2o/RXL41cTvb1JZeW2OTgfeLNPwNHtNvjklX6gjVUEZY+dpoQTEo5bAYztc6Mhqs4v0Lm2DzD2AWnP7RQdsbuHV2c8E/9+kxcHZ2IyAmRK1639lfHkaFr+zhS4MqbEL64bn28HiQDOLfNWNC71pJBC1anFW3nMl8eKlN4A+l/Sl8ZKjPhQYv+BAbnU5IPChAsHCEi6t/5STBoEO6IgI6yp10hARenkitMTKXkQ1aQY1xQXQmE4Iv+LfRHU3FXPFk98F8c3THnUaZfYNRo4eOkXmXMzRDn"
`endif