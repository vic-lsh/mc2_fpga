// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
urgAuDAnWcvKVjr85VoQ1lV2kaf1gnSIV5eJ2lxfdHmSqNSxCIptoo+sAHxa
3DZVmzC0O1CDxkFvAetoJtd4rsVR+d/BFWRfnV2gJ1WgTPY4pbySW58emjCp
DIarCeuwoRrMAtUfDZvWt5oo7Y1S6O6PnkDLulGI1egreEV17pNXraICS/VU
PquPWYFRijj19WXlCyLkwe4pkiyaitLft+h0ql/Dl5NNulhtVStp4WyizQPP
o7c+4RVreeeCaT/w1HaYMPkdnQ2Ys7oqYQxFxx0nZ1UoMkIu25Ww63lkH+IP
YmAOPaKxCqtqO6dr5x7sBJ3ivRcmAp3cwu2Tj4SJ+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xaw8I3d9WRJlZXw7WvzeEm1xCRfwuyzoy4qdnyWK7WvVdnev50oZNZe+1zdq
ZzzaGXkcsp4cNIk0K/j/2hZrihwVEAActaaUP4vcU5t/16zs7bbnVA75+H3c
H+c3sYPTkgTvva0W0D08asFiOCp8WERbhLAVIiQpX9JR2mrX3pEzPZ35rasj
dvCnX1LFuVztJyhb0xiUxwT7HAs1T2CrAicqkb7XDZMmaJkfgwpP0RI3Zvqp
pvLXV/Glza3AzXgln49xxGJ+gq1h/A6y6T5YIgC6c8cv5FSo3xDYOdalaxG8
wXwHs3jO5bq+t1ouhRYtww1sFXESlDGRMqB273O/nQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JpU7CnNY8/Mbo4cKOtqEIS5AjXN1zbSu+H/u4zBOr+JfgvmYuMEOauL84SiC
Q6wNSABHYHgJ5DNLXHpf/Xa1jA7wdaU8li4cJlSGz3K/rlxOw4mWBeyKMpzn
nabSyMWK6/FyLjtrDIO56gzt0uvbiHdGo9b8URJCqayLAWm2KFMCGRNPrueo
8l5FItCz3gT0YkO0JrXPQdC56rhFLiJTvWXewRWpWqxE/Wik5UMJQKyMfsGH
7xNUQSKesOsy728tD4o7d7mmz5Co25IPhgxnjHWIiOhQvy9/j1DCcTwZYOu8
eNQrijW4u0Sx6ytqx6U8WK3D+vf0g5MkP/Aud6an7A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lAn+kBZ8j8II4U1mBD13WEtwwGfVS+ynjgj3wPhxOvuAjJKE3PtIzvLD8OgW
TVUqFbyvLTjbXMMODglDnKkWCfrMLewJLN4Ni3qWp5TaBpQbV7VjE9c7WjMM
/UIAGqbIT1OGkQdk4IsTiA2OHhAmgSobWZpXhJgQ6bcpJLdKXUu2chIEIPRI
JMqSZr7n75ws5z/ysgEhxVI5+bGpukYRskfzYhk97ZHntfoNbWdXQUt0Gf2c
oq0E/0lorvoQn76dNtKVF/4fMTK8Fg9vRPtCM2axi4+IyuDsvZlz5+SZxqhB
ShL1jfwNpOOJ3UerHQm85EdAspSbsGtn0PKDjDIdPg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EprWJ4fLQwe/9HGmfxyxRDx877OrvpH59xY9CZhXEQbxsOsvAPiGPMuOrH5N
bF+dlSpthdrTIvQ4pd5B2K/YM25Lw4pbbvxBZQzM3kqMnpquzsev9QCz5AcJ
I0cxARe92h8BRdLA3Q8dXHDJYoZNYRisXMBGRmO460jMCnACFhg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cQ8qIWFHtmqiK1WbU44dafVeGnDloCQ/WKonNJ1+gSfvC7H1/BWiMrjsVzg/
p4q+dGahcxxJPCamLK2UUdnP9efnn0v4FiPLW/mmIA49zQ8QAkAQbQN8pXhw
SRS+jAf5aq7+/qNE56o9uVfFPP+2x5ewdHrEhkHajPZg3DMeuF8DO25bh7YE
TQ02dUcc5AFrPqX8YHSzIZ0ebSFW0uVMK9mEIhh9EJzF7y97hm503FUx2wt2
KIBGav1wnBmj9eVbHVCm/FQzsUhIP/vcSdzej4JNvqoZuEGMxR4AhCs17SQw
yG2WMZuVyZ5nvG8XUMKw8+iznrm3wsX5zoUPXupJZVRLNiAHz8opcblbR5ce
VA1wFP7N8d6QirqB3Dj/98xk6rc8sSUEeijlmeNCc42E1zrHrrmUUu8j8c+j
qLeeq9PZFJlr5qvnO7uqvGi+/EhHq/zkisLOFeAEQA1+k1iaT5vnxyg6B34K
duZF0IW2i1IMzf9X4mdYYJYGyXP/fEU5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mnALoW7+vm+BzjhzMmYIXlJ4auvjmtdkTl23CdXnk+XqL4UpqYjLKicEXGJM
+AH5kn3m1vOPlBSwi38oFiPEVc5tzbAa6++6KJHOrHPNqp4SCVCbzcEJJxSu
6jhcAR0v3+3podF5camszCDsLn/4Dc5MuL+yQnkdbdumJGT73pU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IYzZEZuii/iwN9MsV+b8+0X/V4kwnyqSIOCLYfPV2O7s0nt3fM8vv/dIWu1Y
eaC/XUcuSsX+V2wRHe0NrtYwXGFCSGlgifMxGnmhWcjebtleqh/YTLcbi0m6
Ig2nussU835UoA0AgRaXrv11uLn68meSSYf0fWsf8GmOuYjHirA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4400)
`pragma protect data_block
kZgKa6fTWOkwPErYC6k63FiOpPedb+sc/uySNmXAD8P0++FTpH/JJMdtCwsT
hU+vpMuB8veiyltKTedNPzQ3rMEGvsJB/5lxvBaZPmF7w9c32eC0IS+nSoXg
nPmn9NM6qGUAjOYD43hMf5z6kfYXhUaKEepW32spbJNH0E1eWSiw0LVr1Mph
sP8KqkrnD7ZWdJIVzICkrL4kSkZu+F5wG6mgI+e5ZHUk7rWiO8suKvYhASu+
56v40O3vbQmH4aoUk8MyLmYFWxwRxCFjA2TL5UhwcXuIzj/pEVdjkTRZ0LIA
tP+qs3xKkIZNgzXbcgML4RfZ6OyGIO4BjWtEkGcHTwCb5lX6MlPSkcFcrHdG
dU91MtoaYciMIXd8nCqFnebxaZt7ArFBVKlZr46rqlvILepMYW0TMH6Z62kK
tjTIUFZb45MEerj/l/s/H1nvPDsCtKnT/VQfoc8yghBNAuwRz3yZQfGtI2PO
1VfaD4InxJWJHy1SIWpzsiISzpMWxwADLzgtiuljwD3Dp1FeTu3hSssMoP+f
OPwyGz9LuWUzPWzsbFxdVchAxFCILO5nOB9gwxLNUBoZUx+MZqnV7rD9cUW1
MFtpAJOWnwKXA3yIQlmU7diBklF/fExH1bk9E65H8TNgiG2+ZcxHDx2pLc92
0/sgToLFl/+gRsvXOAFnHpcoLL+bQcRfLeQCOfvM64EDw9lqj8V5z5ONS1HB
EvhgRNddEUeZLO7SEs888a5jnuLwQcNGh3cXatgZVMZj4AIQAO+ft9tcBhbE
HhoMxGkMwTtF/N7GucfQqL+36daUOql2FcprE9ir5dc3N9OKzKMtlK+1hy95
vDMJf9Z7TOaxHPCJQYhbN3MrI7EwfjmqIvQzXR/GnZRbCF+akKBt7F9XHgTa
xredtYJ70QjNU0K7FMH2WSIZy+zXY1eeyu8cHoCW7phsr5uENLe44Ji/ecGw
U/gUfFU+IUp4txsD8R0WEXodqGG8XhfhDv4n8VQiGqswow0+hnJEEfEmVy6A
GSqRlgI/ayomYVNSRywG9tVcAZqYFReZwpAz87oR+DN3pqDp/rVPC5XCv62d
r0UP9gBGa8z5pcEJIJtsyfbpAr7ezrq0JrOn1puLRt5w4k1eE98DmsqO1cC5
6J5llGS1ftB/rdq2NO5C6g6vGwewD4XFjhpMuYK24uFx1FgF49uowr323b1j
/Jfh9O9nhbXylBAe9GHtPrXPLS1FkA3zeYgTG4ZOMkm4chHiphZ1Es5k799D
XUTw8LfUj9MT+PC4aWstRaw6YLcx4pKcVzisKTQHUIjiPZJfmtB8FwtdR09X
QWMl/qd0g30PFI4itTd7oPxekj93LZROrgoZz1O0OilfUKtLv5+yiHnYKYRh
QQQWHQxL2WTfTQU4O98OF8mnHjTQIiBOwCkaoJ5CPx6DplT+6mFqVq158mUz
o60IBZQ+julLq+QrsbbFintRPLIDtePGL7eC1rH6rgMrlvwzwHmTkzFf1uMV
H8QiHClByXB/ttKdalbKsCQwjXQEod7z9OZgN3auSuSVBCmK7TuJ/gGlao8l
LNOlQlX/DSQ7AkZZTEAE7d0tE4Sj/0si+6Mii2DrogSw6NdSaWz/N0GcSbA5
FUxgnISH2/Ogr5NIdPz4bJ3cpQsq/tVL2wIYm+hl7WhV/eyjRfElIjLD31Ch
4tk30R/s0gfZy+uz+W5NAYEWeaE5sBDygA+jzgJ5XU79exOz8KhHXnDkmRsV
DiMXjCEEu34TdITLZnW0PEzV/Z33KG7d+7gH0eReSvFw2ywn4aZwXJuKZGM8
IFxY2sRTRJtBIJraSbbwm/VPF6U6A0EErMuipjFb5UfYNKseIkxPjdxbJtPn
UwkvNlIVFRL7XVzWE8HaYYuscuhtmJXwf6chzLngI6p9f0V/3POwmYpTDN4N
gpKxL1CuSlmDNPz01bPCDUYHZ7wWlYMUxLoZdUOmdGVBC3WtQ7Yo8OHcM861
p+2DMZY4V7AMxo+fl0lKN0BBPWhdfYlcHQ2dhRGdhmvCfo5CLX/esqEb2aJE
A1d64THqLGmKmUaxDynKzUgphBfDiERlh0CW+dKTyWEgRjleSiklFMuF5fBP
t5LnPgYGn/sgQvwpDHiXLaz+yT0vvfO5Ax/RUs9tIe1a63bsb7I6PRTYJwSi
Y7TXD+QccMjZROoftVwQmLTFzcsWI8melIq+tBrOpL0gKZlq5cpq4No7uISg
Q1D7tvNNiH2lcFmPlALhvVDxV4b1kLipC5OtBw4WBxBP0EM4cwmxLDD/rHWz
D0/oh3Yqomg07K4tnw/DE1HzaFbu9qgn0WG/6fL7YL+1x5LqqOfQsGlegKc5
UC9zrw73lHq3fQ4eglHhUzCQEEOGV4yJTn4G/svLF9s2v2hSXczmbvwv9sdq
lq06et+N6O4bq4Gj302dIxKsUhx0DcxRhpirg8IpBq1zxdtkoSYEm3KfLxsO
cdO8S9zAIiKYN7hNSHYih303B2JPoqP2UpT6O6DNRO9riZDq88QQEfN2s83V
KddVsKOaUcXTBKV+s/0iXXNSLVVaZRU0rei0Op6xPjem2jRgPOIrxYV9bOb4
/pxGJxj+x7lgO+7OEQKQulhEqeCx9L5iJ3mO79G/wNo5RbMViEjEekyKKY9j
Vh7xN6BVmf/m0Wl1ZNQ/dT+DNc5YGCtJkA/wKGhnP+6b4o4Xaf6C3bbVtZQv
XOd6DILEKonsESrq35uR/BvZG/nPD+vZi6YExYqviyMJ5J/BtMTUPItLUBa/
IsGF8gUNDb+UZeAtDqrbVPWanEVgEm3bem+7om/0gjoFn30I9xhDlGKBsKqH
SkvNlAqq3/91FVyYxIxvr/tHoKjL2L2vuILJEmWX+mH6bkgpuJol2QH/5pFU
NZrRSjIa1mvK68wy+6HDd1TLBdc0zSXC4wOH1RhNsmJRO33Iesl3cuapot4p
TfNIloNlPoVp6aA60iRqHTgsngNM0QS7+JRGHnhfhePiWKTZom7mSw56II3B
k5/WxCktpDXu7Y2ye/IN1TxOE5xLKi6WCD8LJHVvbkYuRu/fRS8hFJbIkZJT
9r0VTMmB9z4/kmOI3ku2anbDPCOG7HbYQK4mzfu/Bwwn8Nlr7UfHLmqgyyyT
zbbtp4lp9ui3vt6wZmvZLkq+lkwkpQU7CPgomU41UdtiuFL29abmp0AQp4Zs
xd4y09N3FWG6+QcEB03tyog6vdmTnAtxe0zxOkDt90aahzUDt85o2Q2OIhKm
byQT3P8OQ/kucZO4N4jnmxe8giT5x6oLdBborJIVXN6RQoKeHwl9XTYEHbOo
aXxms4RFWgsecr8qSp31MOlC2HamsurGG/8o1EGxrbfO3qOmFcHkuLUW7FB+
XHY1N/Xu6rFtvwGOEckO7PjV7ZDmzXxuP14lIu13Pgz84ImlQiliMNv4A7bX
bd3j/X8ni1kg98MoMmLEMuN0rB60koLCg5gte5QFxb3NL1IvPHSp8HPEZD+O
D4cO4cPTRgxlBQ3XwoS0TXgQpFp4mCW2MIIADeP/9p4ROUUE74hxe8SmMJsY
GIpf/JOMdbsyeywXPOGgze5rMDVXQUA2aPUUbGKvXjkSBdHd8cKm9GjHK9vd
VC0hGk/kEu5sxKQ2YbRic6g5lEqdUig0qQRlponqGkG8T8Wcr1s4zObX2L/S
t2c0wuZkCbQh0+IvSnfCHvLqcfuWGTfnzixJV9xiHYvxsrrNrFMWSSPXT1C1
7dnlblNng7lcG//a/bjgRwnPgvw4TRNdJlR2F1e5K+ot+2O5kiT/Kbyg5cSE
HIiHSjusKKMkgtoYF14FrarM96GPASLaX30xeqVRDG/8I4LuJh+CP1gVqn4y
eq6NJudh0vLmyd27HMJv0ERPqHXRPG3Egv/bdW5T8Dab0GXWJGYdrrtxjErr
2PpAKURzo9vwtkm1+KCXLgE9qYLynh1Em9enhqnaeapzywAN5Ep8dnrbKb3z
5r67x3xGcdF/JLZ1qZApLelcqtm4nLhPJE1Lb6vV/Da2d1sUInMENAiFxf2M
jTzBENfPu8nZ369LwJUiErAm2l2CQswLQLZ635r2NHgeHEfFbrrQjW2Ylyos
IKOOmsoADnZIZ9ZAD6sq5SHvp5VFgaL1nZX8uJ+yIGJkFrFTdTWVaOTwRLK6
KHqHow56lmTGwxsF5aUYnRojTb99w85JuN2Uin2wYaofjUAKqDCdgkKI5JOf
bsPwLsRU7HmFbR8nA3rTyQ5wU9AZieMZz0zWykLn8PkuMqZgxPXx4eFwVCQ0
cNZOgPHpTXFjO2Al5oGHL/aeu01iJ7S3z1jcoE4tOumiaZzxPYowT0h3bkjf
LYQcG0RtIeJ5WhLJbrl8JIyeCKhgHCl8D2PXGL08o7MUkNAZ6NbDtL5cO74m
1IQ+w1Q6F7pDxsIKURdNrZ40xQvHJ853dowbIbaQJaprKIeBxvmTl+HdX+Qq
TCZ0wMEAFbvXu5VzvRWi9YLWIXnSSY1IHRBicgKNLVAQjurq2ffMVrEH8dk3
yIpbNBZdz7mhdXA0clEexOqnKh/R9uxOpIQMQJ4GUGcWU8sSaEms0o9AFtZP
YPYlrxSrjhdaxXSCnDQLOzYPClStCXO0DMM9N32TmFHeKD8+ocoQoPYcS0V8
G0JCNPTneMFO2ZNvUdKGsqlyDH5xDooYA8UKxYX2Z553sA6d6PAarLi1JilG
ld6l9ysLbyqXVQf6ytO4R12GiC3BRTVpMYAmWpg67DCVtQJLyly2k+yXbVPV
z/0uAWDpGxsnOo8hkbHKMkzFcHD+MnLpJKwVufZXzKtaWtiibIlkWlNOyTa+
+V9+LSOxoWBl3C18h3jOKUYQZ0x5/JnNU8dwNKnew/f+XY9OTFJkQ9Cdhy4d
zLVUOzVwqLkIvG0EC8gy0X+LFHXuikX25PhEKr7SvLeu6RUWplqt6yPUCHVo
sF34BsGFnZWM5i/9JIiIXqCL6mPNsrNvupb+ZQ6YnlBlHY15EfmJuYeZ3nVr
x/9RhVaXGhzaA4tMqQqTQQxpyO3XyRnNQ3LgF70IaR+isAcVs9QE2+ys3NFQ
zQryDXKsUccKiceS29FtnfcE5Y6+S4Qi9GLumI7l33nlG8pzvVs36FdaIY/B
q2WfQQV9RaRFDKjqCnikXnS77F/LaC85T0MsFxdH1rmRMfOk9BL963LgIzer
NjTnVm16jISM9V5hOQKkypopGr7fHZgXLK0zdX5AWCWbB+C/kc7t0SKP2tZL
Q5t5TZ/QBDUK4p9C5TAdmMAumhTLJLNFeal9VCPLL9XcTAlCctOulu2aRw60
NYevcl6bU0OpON9ZCaxNs1f8R5/R8E+EZGauRzL8CBoRSU4Kd94klIPtaegj
UjeXR/px0/SXmy4d9Wpf0vLNfnu617P3LxNNd+n2GkBCHUxVIjq/gCEAY1VI
fy2oL87xVQ1NS/QOg0UKCqVX12EgJdIS/m+yoGmRK2M9H6+EEyLoqaWCGCTA
8ag6lRloq7+5tTwuM5LGa1Jl0jyfmpSMeMR8WFetvHtoRBkCLEMHZgNoWQY3
I4BBFWdWaUmcYBybIwlj7mqEM3eIRYbYgLtYGmKafFiHzn577fT/10a3cUq9
BKc5Gzp+ss9oACvbruf8rh83N/+hs7Een+DVZWiOpNqddX3N/FFRlS3TuRqC
FQQtyOL57loMEG7oM1X59WWEOA3GVxD6qzC0G2a9lnl635LznTf+Jf5vcEeh
PS/THpb3PUVgYDA2aKpnCD8Pvc1EbkH0bo8nvYh/01bTmom+YgT3G9nQqLK1
7o9yd+fkyeK6l9QnT4ykG5tsQpaQOWlVw8oqIjoXSJgWCWQggQwTlLUgRMVU
A0l2iVBTHCyKJEV8zfRSwqU0LZWH8FSFDM9nLwdeztOcCps=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpejIEJbdZDaszfa5GUdNjk63Jst936YPwz9LRmnn7A4kqNrZBJ75WzdUsNGMPlFpBDZ5Qwq3/XIStXSxohcG1wW1Lc0zX8NE0dQZE+0AJYjLdVm2ebS1vudYYxB0exrFvztGSU7JUsuxUAbNXcFYjRhl2wx9RYzlNfDTyZ+i6qDGazGXl2zhr97tQz5M/WbBJkAwmdBdTP88T2mMcQdyds2+/jCSAyv+NpJvRuIOiZlwaIEYfISCzLN18Nu4PMDPqQ0OXrD75RYumMg4GokbxlWUXPzhaaUOmEjCnNwrv3NfE8NuNhRaidOB3zGHAlOYl71E/o+KT2PX6qE4/59yRKaCjACdHwgP+SyXFfmlRcmK4PNHzOBA24KQtGilSaCsB9mKJwNVk/At2sEBrQOrOM8b/chB065Wvn5aWsULlbFXuL6Uk0byldc1LnhllLKuOdoLR7gcj5SK9BWGnx5qkcu//1b4/zpLUI2HLAxDr1nYpGHWOcdgsecf1GVt5DMRGxV/Ta1lwXcvjj9oKT4WmZL+lmIjEMyP7Kw6lMgCo+sN1j6Pdp7LWg+QuLRHa/kg8qswpYMlqK/XC2FbfZ4Fu2y3JZMkgxLYiqmyZ7rAP1eXuPY/GHDRdAbjHoQDYLl9c8zMBeIpfoay0pw4QwOmB4a5XSZ2VYBoNxsqvAWS4OLO5z7ohwi1Jm/hZEH5tzd0E/gdKhdN0ui8B76ipIcaULQ5s7QrddywKvkLxKA7cBCxnr839ZcGIZs9GucT0y9rV77UzPu0hm9cUAOC3fG6zgL9"
`endif