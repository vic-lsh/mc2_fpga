// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FhBm4oG/fyT6jVFZwDRXU9zgKV1pYMC/W9DT/Exiyz6FUwzPDETEdYkz/F1R
aUUoLT42vA9BzoBYSxLixaoj0WF3vqwMM3DeUCQWLEHU9DhJaYnlZ2Q8ZdSa
d+Ip4JXv2diVFYzBe8uWSFarB7r1liz/9Ora6hWI+qB52dszxL8Y3IoYekZK
+fyW0PMQuktgvFP5QwxJgFJQJCBT/PtuS1yCr731fIYi2qn57c09kb3ewjY6
fJ0T9rcZOooJs+X9DwOF9nHO/SfrJuJh8ID3QOrtGTk9okf/553QtnXF4lDU
RcYGTPeXQLeDasly/07gYKhJ8XoeYJfhhvI/Mud6KA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hbWWQUZ5kmd78VRiYEbcAlQvMgoORS7Y7azNjU70N4/LKeIcjQmxiHidgZnM
vfTbe3MWAzJL0TYh+iij1AhA+l/07pLAVjfJGUwt/YtGK8Nz3lsuS0gsfXD4
L1Z7nRouPFOJ71yxgzOzkw1asymBI5cEP6cDnsUZN94tEk0cVoZqo6v88ZKD
NpcRuQx3641DZ6PwYhITDbT8Eb5GUKiym4iorGZZsiWxHMOTpsZbDP9gLB3r
LLSIoeAuBDEDqvpLFcXi4pnHdCq67TeUoc9mAReWRuSzDIB+XFa1rIPyK4x4
O90F+rEd/W6RLmh6lHLExeoABMb/r9l+iY6P8U8+Ew==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S7TrB6EZnc62fZYwhXlaZViMzTjocWXpc1C8qK62mmhT2S0l88NbT791JRkf
7vw/8Kst+x9MN/r9+3WAcfesVmu5h9GsdOPOChg2rkckGShYTbOK42qugjmE
wcWKYaEKgTa+kcSfr53MSaxv3wuXozA6sDGY48GrGLektKzvjAPN3H44VsuJ
9wbzXGAuqO85fM+sqhdBQ89+vsaSqjSvKN4YXQmLC0xfgXyBNojLsKmne4a2
GR/sTHUVe5CzNRuskvYvDXWnUkOGQo8HFHGEwBwBPAOofdTkxk7cm9+pSXNG
i/2ju2YryRBkpbXaOCOR384gReciRuh/MUGEJBKIPQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jTkq63obegwd8m0Qb4EePDJEmzwKce2UqI4rxV1HRSKiSTbrUJ3PWY/h0Znd
BdhIOM/Zq65+lrjapZemF+k0+HuPzA0tMtrVLgE886lg/7GbQtwA+ftP/XJ5
+mTPbH8HYuRfLelbFFrWvGquZfdxB3ImK6xm0IXQzGeyQFrqXIvaCe2KAKNJ
XWxevHkWq0Sf09ACa8yXaZUcxRujzqM0a+P308jdqOdyM+CFzMy596iavnaV
VBGEaZzIOJHpXEa5V9holheJrqBj8gXy6gLJoUo2/rFxksBHzWh+ZabLhUZU
5L0l8VwhzG/DwuzBW8316z36ER7OcbVWbq4nUmZyfA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SF2ASh3hSYHo4EreAXL6YgU4UqHzwO3K5J0udeE3j88S67P9fU20FnaMZstE
6DWDfgYGb17KBKghHdGBJ+hDyVk9xQ0QVznls2bSqVHFaulKBg2t2JccYLNS
7MmrgnqF13OfxhApRtgdXhd0WgOuqcLn8d/1DnPQZC2OKUBw64M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RdqW3MACW+ITohU60bEbAtDuz7fMX04/SV7x25EHJ4Lkb0oHQ383yX3I8iG9
KXVNWk9Vl771mBa9IL4Zd7iTJAvrPMQl4KL+m91iS5sGqKLhuxZmbkJ1PZWP
tKW4K2mYXju1bMTVB/K6SNfLGBKB8jdPRndYqBmXHw8ducDj1bEgutyDKH2Z
cOZ1nxvk4FljWLET5bt+7a8SYRp9KBAAsG0C20Z20G2KOixwNHKYqGQXUEJa
5WsBawVnxu/GCM3k59nbYK6Zu+CLRXwSThGZjfPzxCMz2BJplJP3ifUVsAmH
lrWuKLZ/CNmTjFuPZGSH47CLLy2ZnbYXW5sbhS/mkyU5Ylq84nVEx1KUjgc6
EiY06AZchPnRPlBhXch7y4SBdmzE30patwbiEPfONxDiTN4asMjt6dRlgOLg
ObLtQxsxUVeFAzVradGfAnWfz6sfDP+j06GY4vtT3BffK1sCGAbFxlSqhVZe
YBz9FN+oQyGrVL2bZflfjX/tASwy/s6q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UvXg5fHseB03Q3DpMySU24gylqgudLFkLGZu1ttHo6F/D9AFTOq9H9BwWRa6
Uh66DzpcMq9aYytChhibMCi0uFai+krTk1SlZuSJR+7eGkXzjaQ7RwqyJSZi
ncd7ntOkWWLZ4nto/wjzchxrKNurgLJ5UzpISadRpfms24PHS1Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bfEA0tXNDHPlma/ccY7x3naLxCze/jNdp0BbQ7GzXHhKZaxmq3NSH84UaWUp
nbzpjHd1JoLBSJVBCKCMR+uN02yY43/lTvwVRtMuuHl8/tejgVrSvU0DEUXJ
BRL8Qzgjv5UX/UYU0n1QrsSpaHGTUz7FUrDzKLh/Hivnp0KN2ww=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 247152)
`pragma protect data_block
sDjkQWM0FoPf6FWsZR/vT1TETqiyBvXDR3PEam6IWtjavKEgEMUOwzImmbDV
NwCUC/bSY4q3l4Z8+SZ/h5oHWgoxtFowbjkp3HzQcs7D5JpO/XY+iiqXIWgh
dYMhaTN27W6nRnxkjGKmzwY46ScLrUOVUtBybYrgQgy/TLpRd9pig+6dI0km
egjaNGWqT5oqwtl8nfwJTnQWICN1SbS45hoOZzyN2UkQcJS5zdv8sw4YWdeY
0WhTFnCH400C3/Jrq7I/OTT6qgjP2LX6Ga4Dn0dXfOQp1pW+r1P9Y46CPVyc
GK0DPCb7zoqUqjwY8fCacJPuYZmcKKma0RJmcA8T9KdnF/F7S3azd2iXSP5m
oQdAafLmTIAgPYbKBJ4E1eUYu57JSHo35fIaq7GJazd3KvF+UUvQtH9TOvKG
f/nncFrycYaHgoWD1ZuBTiEb93nhwns3S9NiP6gm5P61IDK9hhD1cNt4TMZU
PEoo9y44wF0ztKqhsvgoBADsjS1nSwTyROr/1w1KwvQ0/YKaDtGk7YrJYBSt
m8UfmdaTc0V/ePy+o2n4IPb/obYo/B65BpqaDxb0hcuch6mAQu7ojaIQqCMJ
ayAvH6QZc4V7sbhuPGikE48rawHi576Q3vU6vJFLkFN+pqtQyLi0yMahDuCd
BySwWshfhjn+7u9jEbHK/Bvt14GSiHaUJz/6XJ1DhzBBYDnDad4qL/Cy9KCT
hbrIquVRb2gp0YriVDc9r0EoCaMEjBzilNjUB1OXy9oEAniWxkYCAc5wxg/h
scQuIL6lFllYZMZ4LzBAwvK7C51VRtRM4e8Hm31Fjb+YzzLc+pxH3mp3KTVX
/IAhXjNgxt3GC1rzjGeY+UeWQJcGuhFn7B0/94AZaRo8RrwHzRNiD4V8VJd5
FOZjKAG/92cGplFv+S5TTBSyPT0Z/y64oSiYLYRfkhG4yT5Xiy+HoUJwC64l
B5zjKq0PeIfBbcDsZinnG8tM2Tb4+2wuqkD6l0dfnNjyjaTa70mCE2pUXeaU
9EfbcqkBy8AOtGCSe8l4zbwSt5G4XhKQea3PNEoLhSLjgSEEGtN+2gl2SVPC
OsWnbpVXCW3X7j+WxMpJgpHxj+gpXVwqTDnhG2+K+zW+c2KXZ+Nf6fEwvV8Y
V9vALWI1nGBslJTGgKKwhKrk4Alss1MJshu1N8VSJwlUm+qKQT9jfuOyY1/b
jYS77MwK+rxpD1YDupiBmzhMbJEM87YYkvV5in1ccVYy1OE8N1IJW+4FkrTG
rUOe7dVqUrh9CRQJnahfeV9HTOzSSifd9/iIhtio4kbMyW10Ys/HzgLjTKit
Mn+TwJ0/0YUCKwodIphL2Tb2RqasbcsasAQX+awD1wO+MvWGdjTDUlwt6q9X
72418a4trl/WTN3OE2QLDRn1eHex9efZVTVvoSg/y7AJk/EsRjfMdJH57FWV
7rq8W+ekfIz4wIk6M9uxf6vdFj6iNII0s92TrQqWvxYnZxHxtGbMLT8tg7ae
T9MYXKoQ2ZRkz5p6wgLGg4l/lB3T/bOhmn3UPBtEPtLRd3mG80R9GroVhaWG
ZNpo54J5uG8ZwiqEeUXebRwruv3gBWs5LwEC54tJtCGqW/le+Jc2EYex60dv
eg5BRsQhdVMbr7U1zWBgHbsJaHmXEYvLKHC2bYckIS8+Hs88oJRY7kKN6rTK
gdYxVb8BIWyyZXjH1swyEsZ+xufnW3z8V9FqcK+nP3/j59fM8ht0bENuTVNA
Sgf4Xe4YEvSmcJpwAzPNY7JkrFlMhVG9+79AXyadCIHNg9rbMjaf1Qy/EFfn
nJMqLOd4FUveyZ6D4iqB7dY3gkYC32kPyooreADm9Upd3HykmDMpYXKiQhl9
ymwIgfLjMn+LQ5kXB8fH2s5Tw4Xcpl+Axx1dJuX/ytLCU61UVbw3k02v1+y4
QmSUNQbUy7ZL/j/mqbTylIR5cYDHum/qdiox5/rPlyrX6V5I38r/96wI+7yV
yHmZ5GZmycD/yHEiNJOZvG6h8Ty4md14NJsjLKM45IACtzTOIITtzuZ/0A4O
QGNEVmzcD6ve4840G8S0zl8lDuMSP7AMJGUUsFWecebk/OJi7gicuo1lriSX
4bHFT92pvFbyPdnwhn8XXDlvmUrOEc3ZLh0wklGJu+VxLMMCsz0qx6pR988f
FKgdlwvB2NeNRXRQT8EzUG3wWC77z59VkRblWJ/ZFePqipVasgiHSypwozQU
WKnGMwwrinwIfOhlFA2pFtF+SV7AgSvjzmbRrh5pGIRlsYKTPUcORkXc0Wy/
PqZsIpF97ocz6jnWPmCDJN55ozlLeWRFOB+TI/VqIUK7WR3mEQwGGxFdxNNq
Wass+iFfuLtDLE69lyqsNzBDzTGjEZoHav3Drs0pm/xZWHQkF8u/JtD0dJhY
mQEjM1CIcDnCB3j+5nXoyXxrXWlhHpsy87/YBp54I31/ZMd8dyUGFp3d8tnj
cg6lmsBE7VBqOeZWjHBCKJTOHu+4darcUUMFBHgUCkzdOQFPXh2QYJbKGRAd
3sYakoO8beDj1itbcLgEIip+6H9zwNcKfaqig5L+VdpTs5zFw1r1+93SZEn2
MofH0WUHBA5hR1BfPElrHb+Diyz1688z8A4oqyQL6K92ahEi30gO32n7lk10
KoncTj/rN0YAR/1gkUCy9sxodoJCrTyyg2L0ZffqjydB6Xr+2PFyaEAT9plt
kfZg6GA5XlHE+1UR4DHqbeEw17pvWKIdXtNt3neMNRbqZS2Ai6qw7XxemPf8
BJS9yhqjwo0VqJ2cH7pZoko4Ufaav+XQlnPVgJEziUa7lSyO4LV9BqiQ5Bbz
87JaoI/PFzgh1iiO5LbUPCeDJVr62wBq1hUP4un+S9teNUR96qSDiauc6Ry/
VjA+4rj6B2i//ITSTE+E9ilqG5iguou3JGmP6MJ4nPyCAyhBXlMTYBsNLAy7
/N/xedgOv1HlSloYHAW4g4hrfNvC050WpH0M2GWksrQFi6R50uHT9p/Xrl2J
0nFbCosNv/jyp9O7IsZgZOJXY08h74JkGFIXxWr66sCVNqb2WS3SzLPw78rH
A168hOj84ZKVztCrqNGMfNuzB9BcRz4gbEYot11U0D6zx26TIM514EmVuAEB
FURUve0SEZP/hZnf5Dsf1J2MzBqyQ2wtUPjl6O19dWpKUAwVwXlfS/AhKxJl
a1VwtGiOSK/7dOXlBcIZhgmMDntsdJ9Fk0vchWELwjg4H6cJm1/SeroQlYlZ
N6YdTL+DEkd9wUHOPlqXQWPrXxM2aEtbHBL6wm124b6iFsnuhp8ToGUShwEF
aoiMdtpE9rL8aGnTnstJZTSkRP7eV8q5e4d1+ayXy9z+gKTRtQPvmTsDnOFT
VvmCyEGKS5ElbMTHJYC2/Tv3wVr33Bdx45fdjpYCxhQYFt4G9O9YxkjvdMw7
+Dm0DDnzVCN9abguNdtdCVtRNhHKsMBeHRaq3J4HNWi8WzwL9TTRnDvvLaax
/gTX0DfIPHpEquNdQNGsEf29cU8FY+5X+XVL9+oGH5MlzNUAC/WPf8bdTb+Q
TNvZkwDZwLY/9x0wvTTro1JHM93r4qloM/7F0IrF6EOLUQRmooTX60WpK+Hf
3D/Uy3+NdHG+ue58gve5dt9GU/dimU7GOixhSfdLerUSLoNekCgDSEFDywF8
GCZetSv7NB998VTDbcSsS7GQd/jEXbCSAIdMcPPGSQHKa7NcbccpH04bEe/Y
4iyKZulb0XnRv70q1yA/oHCuKw4QTXASweiIKd0vjAImJLB4H6yWlsMOOZPe
rCtxjf5FSvq68IykKDFQV1DkmFbqUfAss3O/54pt+5zAKIjuomY0cRF4L9CR
/hVxPHb5noH3jHwpOMfOZHrnk07Cmi5GhXLW5aMbWKGF5pSk1dN+qG7zOW0G
dOWW0mWujXq/8Am55Da1A1JwzH/dmiNP/qo6SIcvC0g7b5hnPRD5uFlSzz1w
jN5GDK/Y8ASHYKEH04LdpF0aRqNEnkzDC5d+RiTcF8/CH6zGgXDUGrJmqHuA
WsOBGNn3OL18cXGsnv09gjf0lFCQHl3JEX4jAK9/uIAMj6vll2k0wPAbbth+
1ufkKOCazrR9VW6eqR8kv7SP7kDzFJ+OEiUPY43eC4pCQO+X8rjymyR/Oce5
2DPP2gkuTdhuCyb3gqPYGFC6OKQVl56K7kcBUmCbjB41NJXz3YBs8YCJvtTj
BWVhc+MclVuV4UsbeGwTYUAED8t4MjdEGB5kV4xNkkVU8UT5c9BTPoIYr/pp
8ejg0QvauAnQPuHWC3Em/q+JRm8UwNR68Kj7x3DTn5aj0UMGnxt52BsAc6N5
d7G7orqxsGKB5f+LzLPoUQaa4A/44pqZOzDWRSaaFdFURIbj2YXRz2STyDYX
/jOroiZNDu1PG0Y5mI6VfnX9/nIhglxLzuis0xhVDuV9N4OiHt+h/vVds373
OhETXB9FUsVpMl8Le2vqHLRQBKxFLUOLvFEDyUW2zccHNl0p34CdsgOYCTSb
Dj+GX/V7TKpSnv3tMe5RxSMMLMT8Z8yap7bPRRLWdG5/bjBrjiJ7yMp5+26/
NgvyXc+NJ+zt4i75hWXhe9lDL8+ZFGUCl3J79ulX9dIgUkn6266L6JCJ3Sp3
fps65zf9cLGqnFt46L/luOZ1udRFSKtjcyluvMyKrMdWyYiWdHM5UJLKlOs/
DcKEDMVeq8It8aNO/p21jPzIe6f1NEmvbctz1fZs1LoJDj8JAknR5GDlNdH6
logA6uIu1bALnL+k7khL8P0Dvnx8SdrHKSfta8sbr0khHeRYCLpO4URWUSAF
GNKq/CLkLmVWr+ayRbQMQoCFBhsXny6I1bspVAVR0YkCpdcDA2ug3QzYlHrn
l24EupUKXkmhsMy9h1XL5VYyMVwMfGURaa5hxS/3RkwvIJdwUqvOmCK2+1Px
lAL90UC+2jeR63Rh5kkRhNZNv0tN9UcwvTNee6bDAyyeqk1sUs62HDBiXUBU
ejvMCjjCABLSUPMj8MN38RCaHWQB5wt5VLeepX7jP6e5JaomfyvMK98/JGG7
KK4C+QRgXBZYdGBiEM/Wto9f++vBCCzXUpgqEnZ1QVZrVStIJX038EDuR3K0
JoPZMOLzBf8N82uUBL3Gmh/fs7AlhrOHYCLP2Asm4pV6vaJfAfVQEDZa1u29
D6+DYzAgqHfW91EeBcuZPtdGxpsRr6FAGkogB1Xc6DtjYH+TRY0XNkhGda/R
prSCT9IwgxxoaH4jKqKvJ3FnjzdjQPHOEa9iKadSGj9nMq907vHMNr/wNB0f
SFozrWamDx4+6MEVPx4M896G/Bu2FVf+lLPzh90xtCM9nWSq0kYhNe2o0yoA
Qu6wg2O36aI8M0bDYLhC927uL9wmkWhgGetPz5gSVQdhbi+I+mL1N3GM+X9Z
KPiE4mnJZRxI47LA3PdP0jxc20WsaDNOlQ0VUu4TP1XuJxz3R026qjbrcd9f
7Do141kaP51WqBWdpQjDIqF2lcZvIyzSj3i53To8btl1Hzt53Lp8uKrObncO
b99DkUNiKAa3MK1ZVHuxVhLqThtVInvUjeZL4nfZVHrFi3FSwUJ49n/SvFD3
Fwg2E7yeQnU5q4uW0lB7ok69jW0sAK/vTG40RkmkZuNM0m+WJW1vtfSdTUT+
TdRgZSKseCRW2gi4yHXloNkKTF3apERbuC0ZrQ4gN2v5veSNvfIMU4vZz8dl
C2p5zAXfEmi3Eg+Ejc41J1EN7xvILiWHmIXC8gHn1Y2WHUiK+et9VdUNXEjg
kWBGxMH1sXVvWq9PGCu84Oz5ZC28aJwGTPXRM1LgyI2ZCq10ZMJfRCPkkVOR
JWy3RuDAOQzWbXNR1jsoPb0rKlHecYEF0UtBq/fP4s8jn2uVVkAeZLU2xkoc
Y2rfgJ1FBhXXF0LLF5ICXpgd6qHFdAoYnNlWaAz0Ks0cJ28B7Z3SWWBat2Aa
n0YEMDemMpRk1yRHGtqJACZKMgfpfZS3GN4zqp6b8CTS70bb07OAmuz4vG8m
yZ1lETX0dHxxQkIe6Wnr/U0nSVQP1WDJ/QSIxRFNadkEc7ITSbDDB1PoxQBJ
nkaAUAa+9JJYbfycVzjBg6nUoSG+6YwcGgRrkeUPeS33UlU7qfRcPgh8iid7
3X3uEWygtp3gce67jMhL7ClLg1c62ngm2OiGTbxkh0euxHwAlkh/phVRIG6y
vhcK8/Uji0/byZm+Sa7RNbPRM9XNhbG/YmNdCO5u9X6QAuZ+ZvMIvBEOOR1C
z8FsIMmh9CH0GMjuH7CFoOhu2Rwu/yXkXEmg8S9Stsc8IY3Jtgg0VK7gV3GU
nv6p0Kuhdikz5vZKw+Mjf39qE8DYAZ+FpR2Hh+TdyPh6yAhwB9Z+1ZxT3HKu
+by9dHSBJftZ63xMu4a8ihCyy+hzWV5iFc3SWlZ06hlRcQgWA8Prrq3cp39x
N5C0nUmMV15ntZbVmZAG6KMobZyPvsByUpIEbeD/mLsQxDw2+osMc+e1yBfl
pXp2g3/mp54/6gAltgEKRxnuJEMfMiGY7bgTGqRFGYMikZDc9iPxRaGz81La
qhPQUvljRYbuUdWT7OJzxPcsEKbv6hpMeTt5HBVOBWS0x1ScIAhJBG6K7xVY
BSuF7G9tsuoPZfOjlXqRAgimwrV681axyR6AjBmTP3jeaKzvljqWqfbyazKZ
3iZscc0HkefuJoyd+ekAxmdDcEXddCsyWFxVFhhZ49ODuqtNpMR9X749sk9R
tLNpXXcEiKaeMsOpLhClyD4x/pdwcwJE8nMlBKue62LWKpxO1J8nSEIvsd9i
GKSrFdoXxpUjBIHpdrcBBimA8rdK1Lq1K2bH4WAjrsCka7gylAdLnosxbFrs
ara9/OKNryhcoVpNP5ZmfhPjr5QKu5kjTwGlQZHclKA1uEB7IU8Mt4ZmHniJ
LK4Og+r3+XUg69A39N2q3HiScOLkLO2dhTpgvbmlYEBrftZoB6NIUpYmn9Am
HUhDVae7II7fmjrTfbZ0WG00SthXKDdupRh9jwApbxhKlvNabhJMH5190asN
AveOmU9tfksDaI3EC66Z/e/8MpZ/s4tBDULe+IYmXZq7sikd/AU9zstTiYfl
nzB2h91xEBPdcN+EzpJ2CJM3AFoCaD0YzUAoMAxjJ6nBBIyAF45Cdir6U1l1
dbt/PZIEi42br82e0GAFN6f4GbK2SVc/sGuO7IX/27U0Rm6ACYmfyAVNxXNJ
j1NRPG6jt58yDn+xCccasgpVW9OhiApYGUfEY/+vK4dA1Sxw0qV83R6EeHyw
aQ4/wvRKV6u9X4iwd0Y+KTT1/ejD3gxAEQEQ7vUE5qYD436mM4ln9Xhnc/KU
gCzigJy63MUUfbPh6fMg9wq4h3TTXjuxKWEwHKVbY7fSXzss+qTMOQ47LsHv
ew4X8AhHs/yFhIZ+vXt9c/9Xwe2HDzZDXjhecxoJGlFr1jHJJJp11bNruWBi
Y+/c0PDehdhXn9K5z/fx3QX1jFIF0K1EAuvA/v/l5txbmZIlU+JagbEke9JK
XLdgVDltT34v2W4GGy8KQO6NIN2k4RaPYcrLb3Kp+yiCL2S5UzzVrL1EI6xC
GM1qp00nbv+1QAh0rr0Muag4ZBkH+t3xdRlCpcJokuNoftTcm2dApDVcDzVS
SjG0ZpNQtZpWsEWC3tTpN4i7aucW6+zFvfavhHq1/GWUQtlgRVuPPuFsrnsP
SxlUFb/34ME95CPGSOXObjCdrWmuUiq+NyTW6JYKQ7L29U03ExM9JVaQRLG0
TzqBotnh1EwmaLBFW6llqmsHVTVyiumavl/PG8GJLyM9yrJOzScQ9zhg3DJ7
zw9uf1LBLlJuO4+Xddg9ogKAleSwNbqt2/PRB5CRMdtFd+PX7icP7NI5Xb0F
NItjh3/DiuV0W6QHS2PqNCj4y//vqJX2X2n1LyWmcy43tHICloBH6q8CB/0k
zrFoasYOa0vhZ+9g77Zpvx3XUA6DpBAQQY7pzqi3FaXTc/QBNMbmkz/xc93M
UmGHhId7YqgvjqhyriAZrC7QIdUswTdE3/NUEtGG8EHcBmmj35hrheVzR4ar
TJaIb5gk7Fdovr5Mh8qxNu1bWUErk5PDAn5C9DYZ33+klU4sz0TDLFpuXqzL
5EhYYJE0iS5j6bUsKPc1adUUgvECMAyNx5OoCuWbo3+n5XYwBj6PRd9qyFoT
dAT4Mhzubpf7tSWZWFgVvdxf1Q9kUL43XdYa/MetiUJ66YiMFoy/8cdBgk1T
X9P8+vTcO/c3LbX5cmbaf6WunfH9gAYXAfhxf3FJuOGbIvxc7EAojbeTx4Nx
P4MX8Wet4kXoMq4jFllxfXXDDnpysQQJm+jPh84pDSdwRGFG7QQVxnCr150a
TqaoGhF1EkMM6LCiPKji4YHZrKbMCEu112Xa0DoBg8Jo58cyIp+AWeo03mUo
XYxQaELU9qvpiSRyeU0gTN679Lnu8yzeZmZzI5Zh7wmSUMMG5Qzyzo/A1N7R
L2Lcs7YxCclhYG91cUDyduuXUDHLG4gbKH2qsgHK7bAhgzgRNf8ToilEY1B1
6qpnF94PiSJAsglKcVdF9oJOJoSiNBx0RL8d2/HGOJxhNl6R7T+LBH+H/WlS
IALs6sqDzKptKPxUCvOvX24LO7/P9ztKYLv40QwpyseR5q7y16gSJMNyTSvf
SYpvyS/APDvonT/rIuOF64GDls8IYmfC/V7jj3M8E5gpcEF7E6qTUCzaMAU+
7G1HiZbRmL8GIgL6N9/YUdANJ563nOj/15dXC0lCZlK0uAXThtz4lEKDYbYR
Y29NECH1RgOU0NReqv6MoK9AppnCMovRq1kYgfzToXdwaImwVfWMDjWDEunX
fxDev2S/gKsslUW/Kmf8daoyUPz3Qg0XMWZYyAsXatO1iwPqKLoadiKzGLqE
+CI4SMm2bTdlkF58z4lsg/Xj+FGk34vXq/dqe1AjVObKkd1jX0qW1WR1W+FV
1KLgD2r7c5jouRk7y7oKmmqGkYgN3am/FOBcq5KcPorBtAbyINtzOunNgo/y
UPYYsuP+W15oBz0REKboAsJuekCbuqAwXpY9Z+zDlRYk+iHz4rX6KpHh3R26
YF7OvN1NfffTcMxQbPSXGmqzvPqcvzVgqd9RCrb8a1Cd96SmAu+sRI5OJ/O3
Fe17IFMb1CM94DMyzYYaXRKzLMONPrwTYL1CH4ffWrGnxhD9nqTaAPVCTROK
AZv29/EkJJU77rL3C1U26d8QULWmStqt7ac5CaeWLZdgaEp0SgaOziFbnom5
GGCSa5U6u5vM7BO6wAog9TaCGHRg8egPnWy8Pw+Bvc7FLx6vd5J1PAc5lSgW
JV0xJvmrbCjD9iiIbCDuImcJWcXDrdJ60D0NrGPmbpCuv5vxjGtvrLqr1imX
LaQB0lCUP146gANvUEpDNnGRDSADCjPE9x0bQ7M63abFyPSBc1wed6ibwoIi
eHKlNyPkn2+GglJ/5+x0Pg98+ooBDwwJKd1Rc1Y0SPwrtQMQAC2fGJcI9gjD
Nlkl86iMp75Vt1Aiqym9r4cK46tzrort/j+Vo0K71EHX7OGj9Qfnbaz8wCEs
YvJE8HZD8o3WYYrR+JpBHveKWhngqzYvjka2Iiuxq4joOnJJfDw+dSR9YsiA
GbGAC3jYKDylvJwL4bLDjoW3yy6pS52X4Eq7zmYamSg1a0EQJdiyJfDkqdV+
d3Kb+GqqX8te2tfRP4t3yKCUL/j2BxCtS+OUfboUlbNFGavBgeXo4sQ/xhq/
qMpgtK9Js5LEoN+MeBA296cGkxzTm4PPFSMsQJm7sraGD6QAHgV34dEFCwWK
WgL6Ym++UtIPfBP7pnPUqvNFrW1Mz8zqtSdieicEq1ZRszWk5xQumHha791z
q0ZvzrU/PMsJrhcFVEUxhEoVB+6EtHWIhFO427N7SsMfM010+OqUYXuMjkzX
ySLqlfI0+M+woyVIjvqlSq3zP81BePiCTni9vdkwqFFM2nVwmaUZ80ryizVQ
du1vcx/q8hahH5U0I1vVTUcO4DSlmiFkBPeExsk3sUoantSORxs6wRs9EoeM
ogg1rd3GRuuadMgVVgBlzPk1t3qsf7f2x9Qik09ifDHdEycIZSlvq0t1AFJ5
v2ZPaMbkQstL/w60KTTHqOasMrF9pNrN9OtxylCB1VnIHb1XN7/XRMwMihen
pS2ETIkRWxm8YvDZAc8Tz/u4e29H37w3QHJR292l0flF2iZJk+x2JjvKJeQG
h8eHw2rDjIqMLqdT2LIthDR8ZU9bZ+ihvfEYFnihu/Omqsm32cUO0d/1HG10
Lu+brSkJv1wEyi6PNERh+14iELeVLAeZhXhlnd87X/kvj79AirmE2O2P9J9s
jJqZZOWuzORYa9YZ/oZPHPcuiPPXkCbJGrU6GFkthtLUf7sSYNJvQeaNU4EW
Cx51KOFK8wN3kG5SQP5zdkga5B/KITlygSzBMkOX7OW3uKRnuLBkn5SAcvwo
W6f3WxeKj7H0wq720bMr287QQ60ONvaUkbXD4rQIlnYy9p+quqwqLlfCiupi
kvVVdZm3FPQtf4nQu4iGpr/PoPs0CqUeTdi4pXlFzPkExYLQ+X3RP1x4ogCj
8fUoOY+ZdfQ7AMOYJCc5sodhd6/iNPXHmeNjs258pAwrhxBltCLX66/vYvvo
qBH1Vz6IHPe16UMV8/GGfilNjBj63KrvvgDp7jnunJxo+VFPz6oMUT+rq+fJ
juysR9rZFzbl4TPGeJGZyY5TkDGidP5TcGpSnQlg3CLWVmlWrWQUcIz8Mp3w
2OUrpVPUc8vNDLGkxRu63/uqeVCP+Fy0guk8D93J7/FpJFGB5IElqO6xHIkM
tytfDabQJRgGuF6543FOo3wGz4SuoVUUCBUmpd+CJIcx5VTULW9IWvWcIgf5
0SlstnmkjQu9cs7wKMBqErjJbr1ePW9tixggoukrlTO7Zw8haFzy2l4dWo9B
uKHdPzPU4R+PqrJoFAN9pwTV1irK6AaLbzx80yn25s1ViblnWaq3qUwQFEoO
t4uTGjqX7TwV1X/IdK3DxUvTvZggemN54mL8popFP6fXQG7RyrtKtuh71Iiv
Xs5vnUbFHj5itwYGXrygETiy4DVC1TuDsgIrMmguADGVreNxAZX6UC9qQy8S
jOZk3AzQrX2unITNnPtgoDRy4gS82jRNmMQUQQ8+RVkrbuQNN1kmYJcL0DNy
uVJejEB9WkYLZ5WzYCRkhSLbAbee3UkrqinREdHoldaqV6W6Q3Uv719jY1/t
dM+Ga9+qkrrishy6rgHmO8XINO/7YKPI1CQ0hQbSHXNuvf3KszHcX72ITI83
C+W8x9EjtBPdPnLgZd3uFaLXdtjqNk2ROwMiY4iRYEMfq0i7ncPXVS/H9miu
0jboDnEX/HWCVSc0oQJANHcIDMQfG8Z5Zx1PF4JyIQnktAoNBz1A8JBkXlG4
S9zzn7sGceihlZUSiXDio3LVQ+s9J960UoVEJHz2uel0hH2kHyxjQ0HLl7sk
14HjoRQBMREub0BdQSaruxgziRoIG+ofV2GwCUsXEM759Hc+OXOigNP5L/ak
I/Dh0tQfgp8TfogUFIsPfbgCo2ulIOw180qG2CibRaLoFxJTnrpR8iI6v44O
e0Sep32uEGrFGg9vuCsl4rRLoMoBet6cNHwqwa5LrSdw+vfTLuSHAN4mSQ3D
ENIFltu0Yt1ueM0cU4kIiEN5S3GYb+HPwKUZMHpQRmL1Z7FXPrpNlpnD6ns4
6TpO69kn7t+ZlgIq59OfZvEk5kJjZ+jWHow5NTtyIMgTpiMwwIRNzBN+pEni
gbWkhAo+eUjTTMGsBrzJ7DcR7sgsVtMLoWRQO11TUMQTGv+JXdFPyBK0e5BG
wKyPvqjN/MHaQOK7n/LtfKM3Im3A/S5NkDt/txRs6eYZiMu0yClLFpJSp+/k
X6vqlCG9dTTFhadGmLcS8oPIPBnc8sP+/jYtphWR4APqkjCOrdjcU5jnGD6M
3rw/jXvrdfTDQ679IqV5e7nHe13ZCAGVIMjYS0mNnO76M4acmTV55He7pNTM
8GjhMb9P4TJN9Mey5RPO3Zt3p57skpuywH+kwnNwRFL/v7YToReSY7ub6yE3
8AgzfokpDf1UJ9o8r/diuKaifv0OIApbWEJZkE6w8PAhy/JCiJvvGpIm6kjy
jHNuNTe0FfP8W8FwX0FaBLAmqYJme7vgPKVLyxRTgqM3T/O0GoQu+U0AW1ol
ZVrUcT1cXnvzfOyyOgILeQwbQjzYS6q0A9+HJhBENNTvks5GlQNLEl8Ly8HY
FZKEocTxI9kEhj8gTmNEJeSK/ZgNjowinloCbqIXJTqu2gOe4kcnIOOlROCz
knEKyksoEAvpgph62CX/jPdaHOiIFY5bKQArsYpLo5HayV4Ypfdj58tYjiNn
YULcw8lpu0+DzpmXtIKt61L6whEslLHyFWtoF6tagcfkJ1jW0tWhLZ/u10Uu
PCO5kHipiJl3rr8Xg7vd36fE2jlGftUdzpCQrYi2yQ4BlmMJ5IEy6ARW7iPo
xlNLXGcI9S1Q1ue7W/4hyjDqTz0vvVAmWYPMNrSaig/Lt8RMIMHh+az1Yw3e
ANzkPYVex0ioufjdcJ2YPboYVuj0+lHAldLJ5pvdvEDUCHvVV1aU/59PLV8L
rzMbWR+DMZUTPtm4JFduW4ZWARJmG+9fI1vYwShV21azeXR1CFY2r0CbnaAn
diwO/CAyFT1LKH1G/CSVpici2kV8D0nStn8tei0uCS/radsjRN/9FdMdr2s2
z+khzsVN4icK1Sl1L99OjQ2Z8mgmw0Gf1w8GIkJ+61D3KrotabRXz94LjMvj
N1vWn/wWv1ABcQjQxZKrF9UbxwG+nHEPODe+yreQ/v8E3cgs9pTOU9yqZe94
guQI7YMHEIRFvFehFEWQoE2tQpFPi4iMMvC5zOxPO0HNykVZWzT4sLQK8RqV
V+Qi5QVkmyLO17Y/u2QQryvFBttr8epLdW/LNj7CM6FmP7E1WKq+m67RmYAL
P9djn8cjNg/AdeMzpnQfsZHXV5sRb5+uXyQG9uFnSn+wukOkc/nfeNezL7vP
aWhFatgPuiezCPCfaDT/54MZ5IRFIey86SvijTm8Hz01tUkgsk9h9bC/+33b
dH8xyyr5hseH11p1o8HcAKsh/EdRCk9OLV0JzytWwk1QbupE1bZ7z3X/Px8C
sduikKG0uIqcFSvr4M5an00f6pwlimfHVr08sppJrSUAqEjPto7RMPfm0zk8
z8uYFXJKFN7CoJELuVntd+s5oydbeKU+ABASUiGD82u9pM7bSo/iH/OC8DkF
3vAGtERu/1tBDotWMb3B6jhThFcC+1p9d4p+QCZUwexs28szsInR2UnyQJQV
Wrb9z43TNhxiWzCbTb9ClVvQTbG49eTI8vaG5Gq36Gy72lYg+jXaDL2vQRBF
6szy2hJufq1QizvNP+2As7H0pax1RRNcA8LRtqtsxYnAgYqcQhrPfbelHxYE
xuU0q2+mvzBYeb+vafBb2kCaE59wHi8WW4sWEMUmbm0GoPciTSAYuayxgl9M
QEGzZUULIUgtf2Ev4wu9EObse91gNf9r+96hoJsnWOKATa+MZRNBN4AWKumo
x0kNgisV5zYXMETsDSlJgGhOVhH164xhRMCcMeY1Ud1bggzMfIDvBBB0ATyg
vdtK7QiUMkRlsyI+epNcchyiRSpY7PhceNfpvn3dgeke++EjIzmbl4pgi1EM
QwcYyyyt6UU6AFAV/+NYT8ASjehWiRs3FIovPSMC+LqkC0a9hTA5VKk5twu4
G49gbfGuFZ/Pk+n4w8Kj10h3TBrUq4iQFrSbUQlmjYrWs5uJ4EY5PqmKlvwa
e3UeBhml5CuDQcFA0XYuxTMV4HR/18Ti2trRccV6WN6GzsxpdMO0xZAco1xw
4mE/LpHlEbg4W9LOXvmnHZDNu0v1p+2Hr/aqhC+eFklPy6a2Dzn9S6zmq05R
J2th+POvYzqvpYrtPbTnSR+emK5a1ztb2wKQy9BWwcGtMkNWq9mFSszZ8Yei
OY4Q/B5W/mKmFZpC94mVVBi1jnyqHf5ePE15k44JoLwZTBwxFIakzuj0e8on
1qYb06inQxB79/oNXbaeZd9Ura06K4jdplQX2ezf0K0V0Z1K+Lrh5JcOh1N/
fCYqfEHB0T3iIyrLdjDJqK9pquiUV5nkHsHXICHoWun1aywa6Z3WuDEO0OIC
1hx9rSxlogTRGk5Q4Exle4r+oE0WK2bmQdNQyut//nIzDb58ubyZrtmz0DUC
biLzQ2f2oadXAZKA1d8TBrZOc+TXd8HORVb6h64WBl3CPErK0QZe4hn5Ntsb
gl/ijE2A3aXLkCM6KzhK1OJ0D7+95rXqsQDuj1S90ZfMAhZAoL5lMqRkTZkm
GvsJI19TB8WfBfav6P6LzD3+UV41157S0vFM7jobnXz7iA1RPrsRA2a3i7Gk
c54CeT0hB4aneVvMFRiMcFuN4iRwYc4292AlQvu+X9NrKJq+TyIN36B16/9B
UZ8K8KrhsMGmWQpZF5o4iKhWhW89xEk0ZZ7B5PkUfrB+XAryAOSDMFx9mKRn
vUaxGRS2dDcH1E0gMDOC9JNY1z835Tc6wHWNDOOz4Vow0YcVT6WWHCJbi5mW
Zkdk+0/b1rKSWuRnezgpkgARjKJkVvGfNbfOjlVsQdOD9vCVRBaiQg/SC3y1
bXm1qJTNw7995CJCObh1NgC95pY9xdHAmW5Mh6/KBYeLLRnAPX3EwZh9gZnj
wXAP8BwQszcD/MmI1RQ8FUBDgEipYqiGcYplSh7frOZMtPC+2OJ4mvKvTmkZ
iapoKKz4R45OEjhQCcwmh8lbImNPvQKm3anf5njfsM+FCe3SYNyFCH/1KFeG
7zb5mqFbUa5oEDzSEFNYTCQF+V35Hesg0HYwv22W0069OxC0tcyMzAWf3KIY
19dhb5M1GA7JEGP+hl+PtXULu4dyFU4xqbZ7CVEY1iqQXkZ4yKTLdwZpZnQN
3UOQahdGwB90DqJ3h/EEa96NIbX70dxz4FwYT9lQaO6bBdV+Rlf+eiBt8F++
gUQDc+r3Z9KSxnkS5fHUfT5rcvC8V94kv9j9p0O6ZNctSUcmuZntd7T1z6yg
FZN/CVAd+k7EzlHmqlstvQdDhL6sJk5eWWqMZ7vGbPKW20I3e1eHZ4oLNgR9
onsDmkYi7qGeb8Bstwl4C1JdDSIBCA9ZbRe1InxYAwUOBplpjDxTrmuZoi04
myHAjL53FgaLYZeQQacu+sTCNP63uo6wQIotiWNp2BNT4QSnZvRt9kurxCUL
7a3mjkr36w8uy1RGBQpsLfmaa/1p6qSEUgzIW8JhvacIxSfzk5Lvr36EyX0s
2cghCuNi0eHX3U49vrO5jQqmIdKVwrs/QuS99kLLkb6lP9rBNAl17XVqAnHo
0waRF2zhnFOukqd3CFX8uo80WRbDYCSYqQimZvhboZKkmGQacGEXDApn7uvg
RJr/TvcgUOeP4/u7uN8IHbPdKW8x7cgFVwAr/oXdqkv7Dg0queEFD/zNeB3m
M/F/tUv7DxBQO0Gav2v11H53Uepk6Sp1G1DCFaG4KOY9Jq4ZApKiUa+jdUo8
Ns0lP5yN156owF4vlVmvJas1hhCVe7jgktd/gZkh1LXucEEOfr/h9DvB79iS
vXd09RcVuKwwBbEiTc+RNgB/7Ti+ploN20FL/0Mf8rbrxW09nC3vFXBkPrOK
vk7hKh/ZG26TbsqdO9xf96CUG7A0nDm72gSbFLUJS53VHDeyYOdI90qTANta
/L6isy7KufSzW+UCC/u/1yuuTCDVvqn3MukF+D0epm5wDdR4NVNI1YmIFaHV
v+O67ogF/Sy0eEB5hC/4jbVkGm8iDA+GBbhgvjiTMp7/N6NXkaZGD/aMvz89
lpcU1dFrZ2vojWnhhz9s8Dw1bv4eLhiHA7zL7zNqlJGsks6AorCoDqYVkpgE
9Wu+3nprT6MzInwCHWXp1aV9dPB7FSX40YBl5zZZbJtzba/6R/A58yxOEc4Z
czgj/HtkD4ygEki8td3a/cqvVPMP5vkns54NkY2nVpkwz+u75wSfN6ORCPZd
jKyBVgXUDAe/NReFly1dUh5GgUl4ATNaUMqWAq/dtJm/ia+y8v+Uj76QXGIV
S3b8MLoJsS7hCwgTvDgF4e26sxhTCLJjpn7qmTt5K5/woTem8UpF3njPtApT
O9SgqpjQOskJ6/Fie6V7sxwMDR9cm/JKEoMlkpDkHb6vGQXtWyEUTy6KMbLI
x+eivWUjcmA1wd4jY7NkkE4bCmgU3JQ1s2xp4gzR2Dry8z+nZmbtqiTRm2kz
Q7Ilb21xsEUpRPfbORRqMO7dScWCZAQRwOQsy7FqqyWTnp0iW/WG9RLuHKoY
7dZ2eLS1Qu7XUPgryL8Ufvmk5K83dzsVfrjA+B5nA22LlvhpTz05XryHx01Z
2rMnfwSvYCNzZpGHhaKbNyjJVJxARNH+7+Pmierh0L21/Melz4rJZ+h2ccP8
60fz4XzXsZo/N8b061HWk59cGAtgGytpZIwhtQtMexpBj6Ti5ly2tazjZNrt
9Lj7TEv5AwU1YRNrfrFsotSwJjE/O1xwX+aExV5je2CxAbC+AA93kdBNR3DZ
rBaY/LOri8QyTaQHmflNkZSSnuT3aI/hVoUthQViUM8fb6ykXGjOOstjcXFZ
1IiSPeN4g+KwueOItoTEKoHKqnGqybw6DUBzBKjhchY6T/6Chx1tzpERu8zC
x5iM5pNHrKCZ4AgHvUfPR1hSM6mIOCe0sI9366BPa4qo/AGQJOXM7Fx0SCUX
ysRMA4spgSUR/ga0Ip/j9n2VcyLeVKQ7PrQhZCYEPMKTo3ZK76EkKqwLDHM1
c/CWyrLQJyDKW6PA7KVbdg6GqYLlXtUyORUc1/eLdsI6juoqgSEVNh8fFBpQ
m+suxSu5YxvtP3KhsCq/EQHLqLVdquH8oDntBVNro6WihIrLS5uBi9BFpyKm
yOA2GBOaF65stcMP8Xk3+PwJhoUQ5qEnrxnlRTwNWqoS+cT1MMpbUe6yfHKs
MQmtZCDOJC+IS4sTAqLbaom7Ac2N9daLIuQghe9UTAT+HuVV71dDhc2fZ6Ph
dZqLnGZrIEejoPuEJlWKKggoXME1lqZLGDaKYgO9V2dIDZIn1nTK28mD1chA
18g/xh/RsvIu6DORE4LWpabKokZxZzZC7XjoxXSpWzO32zLYOmZXbviNYMZV
3qt2VpDtufX7TIzrYgj6kzELJAhcONu2aaUeHI0G8493fM6HhV5tkBsjDX/o
D4TpMDDVc+Ngu9QcWJTL+c/P/fF+qLiuB/3PMy0ykN+8ZnI87VwgE1CBC8Nw
LWJ790e+5ZusC7mzDR6j4HCctTeJQcHALkHRkwG4SjgwajPL57/2mZIWcTEc
fEvLhyefRMj/Qw/B+/nr2Q0esGQ40HiDgqXoPBx0dLPJbW1cACuI8wFSHq8o
WOeAoMN9eKGd+a8PKwp1ebcixuUSPNXOI5dCLk/3jvD/vuNsP46PVyPUN8wf
cxFz09YQn2pH6dTxqFXx/tbgcho6QpSbCcPACWSqy0ubDS4pJuvXVecs2UA8
zS1lOsfg54Ys2Zi9jJfOYY9+lnFPTWlS8sOGJ2ooVTokSrzlWSq2qan2sg95
JOgK5EqcgregjgxnHH7Hf1dEPXRwfRbYsRXH5fOI8SEwyjidCCQKkDqOD2nP
dCqvF3cyga2bcap2H1WHMurBJwWbnp5TrJtvH+0fwaK14l2GTCX+llkkF7XE
nWaYf7xga6NBovVREaMcU5UfhdYCuaTyhZw3j8AO2bZcWZ2wyxW1I64KmQ8d
HZTbQGKUOMmrlCzTSZ5PuWy1/A0yR6rKH7Oj70LITN0q3ewOuuCeAqWLaMoJ
mDLOSVJVVwKn0F6fcHOCNgg16ZfHt/KzqNJ3YIowOVWJ6wz+IImy7wtDY86C
bvMj6f9Gt8ZLRI3OBxwRmTzCzkxG7OaLf5gmsVWZbZO6dvDTSFabZlH+dylI
5PNfmLV4ugp68S78vCv30Dtz3Cr51Ez+SvLAoTebirTA1sRvA2Qa28h9FhiE
dlDl66lET84rMOv02KYCmmQdGjLLO0tpmPMpKT/RlT9oIL4kskY/+ZSzOTql
oIbnFIPruigWngfNoSC0hjXH/B4EhCFNJTTq2xDjjMNck76rQsMx3ebg4zHt
SG20QfFfp9eslpDsC7FY31UuuapGcNtxARZoviNu1qVzj3I6QCmKW8LsZ3xL
+AORgv3qnbKf/DpN1R2n0VoW1DRffYL2Mi7EE+irYb0HTTuZJLOEhmw8E9PC
PlcnWIIeN0JAc/LIev7mecE6XnIi9fyJn1Yulu5SaByAFW5vCOCDar6Pc1Dv
Z+8bpUdr6ASb6PWm1WGgeB8TYmmHCFRW0gWGPZuR380iSFRz/ij1gaIb9sUk
OVU7KhAFFkthuuKcr2Xx5KzpbmtpWq0nOVBi1geD7F4SU+ODsl0KollXX1xQ
Co7yGiBuWdzETHkB71cL+s9PH2w5m0U056umZLaBnIeKYbwDeLxb6iLEbLgO
fDk2Z3ibcUp5VYlQslGnPLAUXJmuKi5PVDfyKD/pokV9J/8usIYHhoCpLBhk
cLNl78a9WLk4zbVPPBzBHALmHB7O9iI/6w4JyEwiRXagrZyVui868tXFUfOX
GnjY6nuAynhQWSVEGSLyRHK5IpzJ+jm+t1BV4uK2xHxeakmpKqtF7TRFIEKG
66KchZIm+sBgELVlBd4FFzxR5BhH8gsMTvwT5Vy+Ykxoro/xeB6NzTfSrLb/
aE4I1D80sFigfyldeILUDBLSxLZgQGQFoNImbsq4LEfp6s2+1SveFneDvHPs
TjTzAKEID+KrDOu59O+8EZ2Bb3cx6Bf3oe7WFMuEZFU3zOvmTU6Fl0zN2Vwt
F51Ml+8kgtSkvIKkU1lK33J9BCyFy3svMDDVmbinAmau60xJhSpOSN42gSjS
lpF4RuLABB5iAx+s4qAcofznD8/SXEpn9ytGoHj2hDu0UHvmuBjH76mursxe
dyeWuepokFD12/TbKFYKiqCdRr1E0tifauzuAcEJMsYs1HVRzKRFsJ0Owd0a
xb305BsGXr9gevlBZ5O0OB12t/zCOBRQbImB2XzTFwQrZsh/BJFD3wpWxWE8
0ieyvX/CrwjpQb0jHL2XL56Ok4fwahl//l+nGf0sshHHAA3jeKgX0kas9Jkx
1sq20HS3z+B+lTYiO+4WaykE217WdtR/r8ThwGlZ6Auh93gStmEU8rYhBzCB
jvevGiauvXBnjhabhZgrcKi2NPuVTHPN2o9UTw+os4yulP6b/0Exb2Jf04gV
ovYJ6HSOByFw7SweZ2JDuBhXRFDQpgwVomRD6gFzVsLDhz1dOifWV5YMlEQq
ipbIzu8x5r0NMsuA/WdX7Um48NmUx5fxvj6CJnUTisUv2nCRnRw8zLbeEnih
GiiqUUmZnJba7wFrqzaomgX/a5Kel5xVvySGbQU1y1g3CQfvB4K2anas3GGw
ja1H+yAbdhhwzoF76yu2J/uXntEobi0uvB+fpnDs7MG7zzMCqvOmQ+xd8cad
MZWFr3nYrGiiLdGhjatTiCrIjc35F4KZzIGZnfCVXWzzOoIPNWpRFILeNER4
w+oRi1DrFC6WIQOC61S79ZbpAWyiNijF9Bph/C5EqG6QomsjkdEunYNt+OE1
7nLCl/UzC7gh8ZT/dqWBp266syqWFyJFYguGD+s8cvTWDK4tonQQDxm6q71n
g5S35dkYi/cr11lNeXeSQ/8ddcQKQbuIU4biUv9826sWkkOgr34zjpCRA0oP
YzRCMp6zxePdcJ0gKvvUl4VLw02VrIMyhEvMn+thVTc66wpl1xDSG3N1HfG4
IzZI4YHwuBfrFuTe6LUP/3mj/v5EuUyAPzestLTVgjCgu9r03yGNMGCdv4gI
Zo1lClSuiFT6q9WpZsGZ3CQlw309m6V8YB/EmI6L8XemDK9gPgp5SVhf4sd6
w4CEliPWwJu2caK5aF2pdTNe8gnmwZW1f+WomOoOHGjGjdXBh9na9LWnXhCo
50c5KVeaHhjLXIAQG7wuRGpqGVsM0KEoJ7iJ+9WgT7eAwya87jJ1+tFb2hQZ
ntQpuF7tV8sqgENEacU+4oFx4siQqPD7JBfnYP4uy5xE9I4VDOMQ2caagyBV
AaopTaFKXj8euVCT+aP1fWPs6MAY5WXLi8a2lYfFtFV7MZ6Ea/sEnTy9KS0r
My2Qqb8K54/v+6FC0TBa1FfclXQOjCOi9RFx2YCqJsc0OjlRrvDv0ihyyXcE
hCTUk87yDFCDYJNpLlTLh6JDf7R4mYeDlVPuvvnVV2swtD0ZZ0nOfwstLEg0
4wpQ7GGtsKy1cBpckMB88Ut3Fb436SxGIMkgUrr4pHM60p0Ki3i7Zrn3qxHd
TwAgAH+bAQHFT6ynY2L5scmrAuQbick80frCqb6oOXTbPVWO9TtVJ+cNTMCM
dMzzr9u8X5PDrqokH/oczNT/sidY5eM6XjzWfFPJ0gJMoHN3sI23ntjJmfd9
bTnSPoha8Uov4BRLapdJkaDgY/VSDEfP7N8kVuWpppnfrSk0iRm+XV1eBY3F
bIC7GbtaOzbqCZv4GR6Vdh0jYA2s43Utv1Huna5Wt1SLsTcd2S4z6m9AA7Le
9XjuPr0CiYH8eL/DL/ATD3lQmEJRIlLl6XCaoDvFkMMXC0nEzEy0xFh1eFnw
9pvzR30k8pn+hTAZyFHRRdRE0pIHkSzrKEOy9kUoNOIl5y7ApTu8Y6Vtp+ZG
N0Fh+GPQHnb+U7RusZzqkdg6HSMoOl2H+ydHF+dDEbG1yntWCqTEs/95s85H
4rAk2H0gvN9rr9LTRaIPx4Xr0qBwzgH+h0QZaIvjPfGAmocGyFBFNsU7Z2sV
hcjDQ12hozVO3ZknCZE9h/lLEG6lsZdN4GysTxqNkxZVQyWiRjotxKbAZMNa
7xV8EbD7NquWAsIi4/tukTZ5pBQNgwlwgaMDWV7r3mSNLJITdTMO1tb1Bgpf
XHdnlmhVz6TjrHHI+vJEQQzfc/hyNVYyseOOpRAziXHLzaAyZuY8Bb/K2jmR
yKXAXEKmKGfsFInd7ESQU8sc10aDiRIXqyJ5ZWFXjTwzMKWhEFl1GTrH6loa
+owmIdPi/cStla2uPeUX7XT6sRL+oqqdQP0nKG+HofnT1NadNFywzixXyNtk
uQ93FcNTKKE0kzFQgKUupNVkG3d1YP8FOGld3hxGYXvNxVDRRlLj8u6NfL34
PwvOqMf9UgSi6gSKV+ha314gNw6KU5iys69wMWYvVj2m9Bcj/+YFHbSEhWWp
3lG4RWA7rhGlRlqu2scKiFg5k65/2lXWXquqESDPtY0p5mdZ7FiYlM9Jtlx9
sdSqce6tKnb8G5YCEo1WRbt8VSES1tsFgDWMRT8mRrglzzUDONxAJ4PDOYES
QIj4miw9sSsR6kx5LBwIYXz9Dmf/cBMDkAueGt4Bz87lByuHsw4FzV3mbOP8
mctl5cA7doAtHx64VHxXkiDaESKqd14tBeJkc32Su75NS2RzDEoqhn5UwWUK
ZhkWJbSzKkrcE6rMi7GneO7LXTxdKcsEAJaV3arc4l4GdGWXHWVVmGYUp51R
hcqll8YQLYwL0o3DjxH2IIVWR8uqkw2UomZBw23t7Rq6Ql0C+09A8kRRaIro
fV+/z7duY2qXiDkQ5Yxz1BEKsIOh3pKf1SgvfJN0LmNL2UGUtTbL94ERx71d
VqpvxOOK0OtcdqeoizgAa4/WzqDUgRXBQy1H2SmGLZnqF7S7yL6afA8fNXxh
b+Qk8k9Saq6f2OY4pxwFZDp7eUV9/1/jW1HsQ/lis7AASrGMKMb+nGkBSG6V
L/WDymxJtGvMWpmDrg0Hop44IitN3WtftYTXg0i6ga7H9oq1qdd5Gjpk1Rfu
Fn1JK9h/ppppuDvV+/IFKVdrgdhDc9Tmd2fyBjDbif79coKWOph+BNz9Ricf
NKUdNn/uz6+11R+FAkH349Zpt/Z3xZH7yzbxvmBq1f1Gd0bS6/KTFzlKq7bi
vYcUCMN4LDLIzOOVn4IT/bE2FADreIPUgKzBPu2syBiMcVJBOh/jHEvgLw23
ancLlOhhMBgGrYbNnrHh+PJQ/+Cn7FDIuw5nTXu7pOQ/e/U+09DmpBv0aJIV
mGURvC+to9MZHwU1zPiEGMJawiv1KTop3l0+a2T4qjlCTAh6c+Hk9X41IFSG
QiplspT8fGP+DDf8qA0Z2g01bKMIJhLR/7aUcL0kW8z0J7UOtAyyIP1IBzSy
It169Wy1UyJlRCPhjoe/+pXO4DGNRvyRu7amWxS/sGmQPzp9BLbqhvNp9LqT
H/evHeOWU+1NEKYPC6ud1TCyc2nxe10js/Grzps2CB6EOLPfKkcYg6mdBwAs
L3rQjpmc8wNML9B5cBFwDuIKQRdC4q98HWIytPZ5RMh4jmV14LYnnpHN/plB
+gyzjPCwe7Wu4fE8Bt/939OsOkI2SyutxanalSjPxXd5EbJXjmUcXNzn1jPv
aY1KPvs8gETw9nY3rvjXm7rcN2+SuUD+u9VR09TccaryaZbB/XX9Kg8J0yvr
xPFhfxnx1NJpK3oMv0jsgAg34a+E1/hCjUIplu+LcMDgAwKnS7iTfhZcJk8m
OG2Qwa6TWNKesdhsfWC2N3Cffp+eICHIuG8rmGvf7wFZqXNTGbYd7kfXqLOt
sDt3gSvBBUGEHFqREJ2uwh+0omIvPBZOEaqCbHqdVqd0tA4ADTCu+b+xPV/E
DuNSo2kUCoXeYy/IFOPffraN2fnUHNiSp4E4pbsur4JO/QLS/Zly9wRCaXk/
3jV9isXLKJJtV/7zcUDpnl+6EY2N3DKtTU+Fg/QWvN6eUX0orqPPTIqB8PFa
VUcgHKCYH/Bd7emyMw5YXLvJpXY84KGhBda0X1Ui/ljb+4YYcjbkncC/EH7P
aIl8xcLr4FszCpt41yUpJYEs9ez9wcInMcAkQK8fO2ahAryTSOllJ02QD5XM
4OLLMl3El5BMiwM81JmoPyttaneVag+OhAy9UJ/dMWExQjeHyO3h9NivitIs
SUpzCPC9rGSd6/sNhjpxgz2xuVs/7LgTq+4XNiGGv8pRjVrcCrp4Kwq0EB17
/+97Jn5y28xoaj+ylFXW4KdlenSSafCX4OltXq2SPX7XhlViBoMuIqVjX4Ky
iIO4jCRypahgtDW+DvnwhEzrCd4S2m0f0iL06GLqFOUa9uRsnHV4nvoyA1s5
SZ6GXu1wzx0xVF6I9s5ZtZHqCB2xRyXx6EPzjyq63a1Fb8OANcei4x1yAaIg
s7xoUEZofo3tZVUMEiBbTEvGYw7I3J+6G5aBAnTcQOSPAzXWX5myEzXIS45b
YQ8bVy7BIabqMG9KYxR0V0nDxwnvXbmhfYMM/xwqBzDFVrjJ8Iw/VBEzeDE0
wxg1HD6I5IbXZOjgBDGHaITw3rHpHNjlBy6CoQst7EO4Tv9I2+TjZZdBvYVK
ewlOu1kDRTrFQwzVACVd5Qox6oalG/T1gjL+rFCSn7oQJ5nu7TUforMgm4Xi
EDSfhkbBwaEuUKmWJkAqafWuxC1pJfFKNuYIGd8Oz125wGEQEK5+VeIzlTfL
pK8jzQlFPZzlpsmkdFoYt+gDyYY7tCPJmHIjRaJuiYhewdvJODKJd0Ibewrx
5SxKPckAcOfmr7uXGyoXplS0JVOjc+uOk3l6/T7Y8Hx1OtO2zAR/PKB+uPEG
3jQMHGcaxyip5V7tl99vUeDdqHhf4cnNeXR9LDjdz5Qtzby6TrLp7Lki0tVx
jnu+GdW56W8ihRvBAUOkO5mjF4qCqBpgHIzmBw10EkkYVny3XyQWWE4XXZgA
z1H19BWr5wBGWzMn4YUpFDLW/LGh9fh4goTxMgMzbPHzXhcc8v12H4csuvWr
+D01W9mmr/7YGnHmCql2P53hPurOI/XuKO4dM3Iu3dKqpQOfRKP4lbzqu2Qy
g0ePI6D8aqjr9hEMyMz3sKpE6KLIyhL2qKAoXcD3T637Dhre0cw1UDcP0IiI
kPp0Vme7Htl5yJWp8ODijfCkFPHTRLbZolQcw8Ps80yppOY/MPAPq16QbWok
wTOpiUouhh33m7sZJfAOkZ0hWES0k+nGiL4hzPqt4iHkLH+YfALjHqXyTX5J
hdnch1X7jJegp1tzFJB2zE7QU4xHuP0RO33eFRcD5br0bGrKbNVeEzz4cm6U
t7+G0vNM3VGyWJGzYIeiqYal9ZXe7JZHGaLARvaofSFv6kitTpPme/kWaQsD
tQkK+Jw9j0hwyoIvYp/RhFMIww8xyLoO1cmNOC88gK7Y9c9Fs//LB3LjvVZc
2FiPRImh3swpeZGf+XNJrK2TYhUtRYQBbpGsc0/K7a2zSfDNtJ2EbyhuEhHE
mkjHwJ7V2cTlXagr6VF+OUCgzH9drIdMQxyOmotJUObq3DFEoGVNeYbHxJKE
FCwHWnhEzhtAUVC64hjFt54AxNjMVQPj1Z9ypLwVx14J9aCBNW54GDF5rglf
7vl3WFwSXAyf9NanpuI2BOPkLww1qBPcVdzwcfkyWAiW+77HTS+nTvrFRY1+
KA9YNbbC0e7HmYSkCceq0U7V0Z/iR7f/3IyifQs75q/uaARKK73HdOVqb3Ah
K6ceMUJrmdPkGdzqwzUIbJ7ysACO4pjse2Uy2Nuh8QlFtwF1fZ2BPEwsgGyR
CXZFGAV9djEgiBIkexwP9H7d9wNODvdBKlMkbuGAhIaCCr9ZYGpt3KRfZjym
4a2QzPqkZEn5/ex1bm7xcURk/BMZXTWPKC+mmGllXX62HGpWeaszOi3pTkcD
wo+gC0y49VcNxp4KNe6NQZMwQz4QPsl1nQqcaNzqvqaZ+lbe7pF9SXB8Ma+S
OlfhVxfNFUk7PUIhctNKXS+UFOIJltV2IWHvzrlDeT4xl9PHZ6ojIgy3Nc49
OAlHgmoXg+OvCXwDV4jGxlmBh1q3fnWbVCaoVKa5vVZIhBb1z9HjuPt5VQyv
gYTZiAXXwEBFaDyYzPMYIOFT+bmxtzO3O9ub7mdlAbGrBM6LsXvbD70Nxq4Q
V0M17qQQ7uPzcI2qEaSancJuf8mfwHGcpMk0X6kMbLDsJiAIfGxgrco+LKZq
p4pzrqvQelo+V5yuz9TtvQBZJ3/prqj5Mqt0WWlP+/tuSsNcr6xO6iXy0t3D
zqmwubzFRyBm7sB4ArAQDtE3Df2Gn043k9YfLf4+GV4o4MP7dLdQYWYDzX0q
yEnE2aejCekd6/IVkiYRTQje4OmirIaZqlIQRRHBb1ZgqYH5bf2Kooq9SIRf
tPQtLuqp08e5mhz6dU9sBl86cPUcxHCSqvkPZfqmJb7+co+fZT716ECshL/p
lUekyb674UjcOLw5NvlZF51ULEI1xUYr3JF8pcO40aCn0dPF+rVKfRGphUp/
U/wIINoOu2qkMX2HFucGI/GPuJvRj7NiDJUC71sFgzLVWHatURyUGCYfg6G7
shm3sYVQ/cd9n0cAwBs7+BseVl3DRgoG2Bam3E5wYmPky/E45UMKbBcnSQZV
WiALyVllBjAhJq7PmWdCzEVJbZ8AiowBPngOw1I5dNYUDz1kW5NZZV1aesDV
oCUC4axkjUV0YLRCFJoLrmGiODkjVAaTPLgR9AhrOr252rLGgtFxo7xMF6XN
Nx8w9Fqs+eyz2AYRp/lHIgCj8705ZS5pWBDHYRP9O1OWLAt+7Z0gQIU0Xjyq
NM+kmVaUfos8+si/Hi+VUEuBBSFZZFu8OyJz/iZh8YoxA4dCgYadEn4L4Yo+
tVBLBZjSRLTs0QSzimrzbNmfcVl4NOrBIyEVcAl2VjOYDT9Tl6yaJ+LwOgeu
VRtYXgj15ypfU1qN9srLj1aNVHbIuNwBRzgG1CKFXPOaqfWa2h2ijVicrjac
23rHnE6GmWU1IFaDtYfu6MYl6BzWrpeJhu6SOhG+SuSTvIlYcf1PgGzCiCh1
DYUOtLfvx7zb18AQMsoDY5D28Kr0wZbUnmZsaZwy/vr0jA/NSBJVi/NkwFdz
6KsL1mdOMRbvQCa5PZiVEcbK6+0GiG6HLF4Kg4oOBHwWuay+nWpArUFhiQVi
eWA+Sc+Q2uo/GB2eOQfQtKZapHVBvuJTUBaeksUPT6XjalZe5aPDn1qQd6uH
yxCAVBvCcBN5f0a90sC7qxMOwujdD40GGH9c86fZiMvX/m6YmtxuR1Fqhh7u
ajm2uk3sKE5QybvL03Vx82xsVtHDQ1TP5oXWOTTluuwZ3I+oQzmIjw2C+Dh2
BK5VDBlvhJ0bZgmFoWx0xx9gJylcGboET9oD266k177hrU7uK4Cpl+ck6GZe
Kmcn2cSpxymfgQ2NxavJOB7Q7iTl4QNdvlwPYr90yVPJbv9PPfZxL+hP9LB3
WOMQvOe1oyBppKiQEFri8keeFuCL/8FTHQQ5UrNM/rmNekgFeNW6uyRNy1dL
5xxBSUbSvEYBNy1Q8eX6WZ0+/F0NS2alcy6e1WFTf5k6VxJHXyTg+lWBvTwk
RSCh8wtv1AzhFWBHQk+QVdYWAdSAl7RQTrYp6vxlTZ9elJAtD2wrHDfa0PgA
3At+Db4T5Rcvy6u+6LYuzR1bfzOvaq5L97lxRwS0lNOvyORs4faOiANQm3NE
2lmbhcDfKEVwvDy72KBRK3zw4VjFnLkUXquhrYu7E3CAJQohtjm7oouAegy2
PTxK3uNkdajUZPJ4G13TztWfPi7B+KqfEveDLSKWDtB8GHTxrNbd6CVaR2Sg
oP5H7Fzyw1R/PF5T04cGQ4Q1nw0gjDOITtEeB0tCZ/PuC1XU1DICMJaU/Ug7
CVou90jEB1NK5hS0kTffmAPCn3KpFaIy5gnrMYp3YNvAr/xt7euxAeORX3ij
/UFPsAvozwSmt4Bw7Xg2vedqGIByJS0hVpoSjmHGcchH6bTTmuBaBNU3y2w7
I04ry3PFwbAyjvKCjlJcazoSAnXnvaSn0ESeUNxD09bOCFgoxP+A5FRjXUpn
fZSmz2VdKAdhZnwcmpWoIHQkfXIQnwV6QIFUmOOPG295awmE6VJvL/aqj13O
ZcsK01SuKZrbBCNNzPB6JMBlceAsheaynL7nmcz7kA267gzM+j4XvmxVk2X5
JMtCb12MvnYUEq5U2tYJeji7JVNS0hjezGTZPI5oHD0Fa1NEi95uqrbqLJk8
7YmyUiKgINVKSFGvchS+KAtv2CCEIHq/nO2VHE9qAF2HYikNs91YAPLcIAGG
TavJ1xOLf1cCTx4WSJtYG40LYPYKiHmoAEzid59Uyygeh1+4xSM0inDhX+Nh
VnsXPRSGj9vquPn+GdC5W6WMb+rqfZBeV2KzJ12KNy+gmg4x21UzUtmu+ahS
IjiNG9rztbHRxxBCEYimmmfrZ7xvgUlm6g9GVLrB8P9b+hWn7n+zI09oncpE
8QDRho+dtE5f8n4zzAd5nvrWZ24W/um9RnppLBaqn0M1lMBWS/SUe/BEunGy
EfFuM0xbbkAFRWZqConb3KFmDd3aQmWSHUXiUnSfhNNWSjjdYT+oSbwI968f
XCgCucoDC8YjLYqRq3ID2a6e8nwf2U31TNm5ptvWvdDqvHF4GL8zJUjqxPuA
21ZHTZ+KLxdCj5x//5XrKD9OyVeEEdYzG1OGRhLxslWQyt02a61ZrqYPc7g5
k1h0MqJMPHDJPhWi9OYKP1JvylXe3e8rk+wZac0ZZO7ev7OUj8nUwagEkfRU
521v7tDvR5GZw9JU0rqVboNkJV1UWyGfjj7NV0tSjrGwzoGuIqIekb+5B2Le
E5Z5fBf1IjwSP3ZEUok73ycqpfjaUm1CEKCANoYToep4Yfk/BHyaMH+vWhps
wdqUi0h7fQqMvfbQxmW+zCzVaI2TdY9YO4gqL91SrlIElo4RWqWJdCawftxa
Ct/cfAOV+2p9BRMJzItSZ0MHb+VygTWoaWc3GInZid4pVvd4iq7mCB7fdL4Z
fuF1I2efrrPe2eCDPWNKr4cgWpJItmiCnSt6+olnUa27og9RDIkC7+XKnzTp
6FdvHWE05SYhPNlw4xTFV28ukEvs08eWb1ly9KijhgpGjcqxlNDmx1qVs7ZI
lR7l+i4VDt8IkJrMvaP44oYCvo5sNAcn5cUY3lnU39PAJ0ecGQ1uXc6MuY4f
WCueC+F5GWsmDIjZV8VlWcjfZyKAFK49wE/T7027YAgLt04GLf1dh5T5M0u5
9lAGQPO9IUA44m4U7ER+HEtk9GYRQh03iihp66ocBfj4w5cX4/DuBJg0h44J
xGYPceHgs9hI/jjEU7CRYcoa2KTqupFCDZiWtfIQwKWgNFyH58nr4NbuCZw0
RIbfHeeINtMb9oz4HXODKcDBjLfWD2K72RJKU6ZQwn1T9xBhPXPSG0lRuUaL
J7K7hBJwWoUWEqUOZOn9bS2rstOPUvEgGb/ByHvSPZnJLW+r/wMpEHJwpz+u
do+RyzFL8y8/NX2gq2RGEOBFT81EZmEk6miQ/ZCkbcET1Qb3wWEQ5BtfKnqs
OZeAkLi7hABlmGcJz8bSbCxAHv/8JBV5PUScqbXdKT0Ey5tsMmys9CKtYxJZ
7zl/nWpQ+S2kgGt4FGTrabLgdhU1YtCcB2Oaojd7v3vYkN8Fcb3xr1QNmfRz
HUDf2h8stCspcGSY9vCD0izWYzhtuStcvedah+g0gDygZjc6NeIG17PigI3u
XtFMnOPgHY547ZvPaauFvsZ/8LX7EFK9z9pi6X/23/2GP95NkpLBhDA9ler+
MbYrliHe1P49Hn0CFLpY41PCzAbnu1H0Kl7pk6qUqBglQYZdOnYJ5IAyYebO
lNoLxef+Pw+dgubem9mNDZdXWKnFjaC4vTur7kQIdcrYJXDvvkruarV+qpEJ
KFViQWhZ6A6Z52GZuHMYXzjxhjp/FpGQZ39ZzYJewyAvc6veRXuR5/i1QDRD
O/oJFxkLJ9vgYkkFGCRJLCA1FBua6NWeDtwxQSMBWY8dk39DtJF0qnz8ZY88
GspcO4cC60xFR/HIn8rQiJhi5HP02j8Gb0XE6yDzJxVvoiwnAK6duUrrxt7U
7RNNZk9l2KFLUKZzRw7Ufb9YIVwMZWUhou+jGTdkWkfk8SsheXdIcOr6budq
Z/yyNayrE4ROT+hMmXka8mWuqruFb/dfxYyKkJ71w59u0t/0lTlhYek2W35U
DF2xGXgD2qSoQzqo9gPhRqZsuTNEUQqGEedVA/dnVlOubfL9arxxb1CWLWmt
Cr5hvdezLNrZ+RpfHDfo1IJsSDYWjU+0zGAfnMwtWpofmY6EWIg0eDsLZmKE
Er5bk97LOdiy9MkuNqaPT+MYd+xLnrQ4ahmRl/xNx33EkciKRxr0yHU0PO23
WlIVQ6QEs5Ax+/buJ/Sq71e8phsg9BuBokm16QaK4Z815KZvCYqSJ92a6iGB
2b/MQ37sx+mkJlZTbSGFo8S74KG+uxvnYGCPZPOCAq6lcmgBgNoz/vTwHAZQ
Uf0Uq4VCxKUoi99TkJ2Nb6QvmhGTlr+ebLQWyL3VgdGmgoJIjReXTp8/ebKu
24ohscaOqe8ssucZSp1dY32rpvXXny9q3PQwY3iLpbfAu1vR4drv3dL560NC
GldxqDd6G4viyXyp1Sy6nBxKt+K+DvxLbMVDMgkPI0nJznlnePsE74TUm4w5
q3RIHziA/5IFbS0N0DtGyFP6E18gJVAVm5a1xj2atyvxYLGbEl/qFNV/ylnI
LM0OaZGz/uCkLPh16hsjyADfkNMDU8pZ5PyD+8UCVJYMMqIP/rzSPOHTG8e4
Ez9tzhpw3jzmPfuRZcllPgxqH95m200Uffwfgt5flSNiJ72HAUoHqnFpeNGf
GRm+x5ycbFdDsd6dEBlJN0zV1HAyVZy0LW50LiyQEg1Q0x0R6ORPrtNTAoyy
ptCcd58FCI4Ed4AH9dhiGg9yNN58/1EhI2R1IlcK5xOg/sYdDB3QB+1AHekk
r3i6y5raxDW0FnVn67xkL45TBy8c0pNWP9suyQQlCXKRZXkC6UsvdNh4wLlw
rFKAANkFmhvNtFNthlGKQI0kSH0Uus4IAA/DrZs7u+2NJo2YOpJQUIhre8n3
alJsVCwLvlFm5rbp2kWLzwRPSnkgw8uwNIggalkhJw4IldaqC4QoWzK3KI1r
FOC5+i6paJGHOyadQ3Fc866z5wUYqFrJ+r7zMWIinEfU6HsDUeKjlQfUATtR
cBRcb1VtT2y14odh5dTf8PyxVvgd35XtG69tPfy4vYvm4DN37sqbI5crddn6
cnSx56hP8gkH6WlCnPlbpdbQ4rKvlFt6u+YO5QDIPHNLdXTDGb8823BODoeX
4PuoIZnM7MC5SL0fgHTPH0kd2Lwf0SCAxq7I83LCGee2mjvIjhvC6eq1NBPU
hBIjOf6i0bK7Ej1qjBxcnHKqnVbtMNSOzYfY3zhWD8c5y0uNoO5Vx6/AKE5k
TS+OwCwnxT6DgzHoyS8Z1+X6L6DJuYW9IxjGEJ9NVDWLm83z+xG3RFTBAX1H
1MjaFG9I3AriSS9YtSbazeXzvMLmMMQoKyYYsIyDojOFkyOxm+PaRT6/YfUo
8JFThGZfVdRUFJFBQpVC3B1p/LE6skQCL2ThEkAw77ahAaAnOiX57G0ACuXV
7GhmB3a9Qv/BAGU0iwqtfvtW5aed3cUW2n1fEykE6eoxO4k1zOhjuKyMr7mX
t3CHZWJkWxyBZ6mhVT18iQZINGfzowej79XLonpqVjkspaB7zgO7NpTkTmZI
k1H1cMxdU/zfXZrRgM/RJrQYytznJG7HayWKeiUKlCnXGhpvP1MqsFBlj7iQ
QjgVAgN+PH43C1ioAoC7I7GYCh6SMWhtsNq/c+GRVsj7fbnDNOr4gNx/dnzd
dDEYHqq96lNlbFL0oEUIokPqODN5HY29uAyOr1xii2PijgQBUibYZHuzNv9l
wuzP3EcpOu7v/u6WQ516HrW3bI0PGOM5Mgsm0rlDaVgvvNoKkhRLXWYqD2io
eXBTlxBhC+D3H3X0mmL9EuSm1SC3szSXWPMRwmygqDntvflwtJYBBtwb9XOe
kingC2LMggIqLhJ2MCQRLwqtmFlB2Z1jCYH2ITtxHSETg6qI0xYNFYjmQoap
j7/MRCdylCRFt23jw5uWRBD8gctgAxG/sGEt8sRnYeJBtG+WpiIvpuAioavc
hi6yylgzDkaB2rMPVI2YIe4jHZzpuU6GjN33wHRQNskwvPbQlrOPDmsBT/ul
v+v4JwrvDVckY3+NsV6u5Am5yEFK536Sgc0fk84/M6m3/+2pfiOuCt5+Kemm
ea2U/bJFIcHKVTrCzgg8X8T/va3t7G0AbIrxAGvXf9Yd5tdM6UmqLvvsFtcN
qdQaw4m7Fd6MirNsF5ovDuC/FzM9akp9ek9tu5EJA8H/7s8aGoqFRgLtosgY
CesFni38WsMhTaNTnCdvTlNxZkpVIV1wp29QV+xt1sshof2O5l7L5SeYpYhA
90iZ6fFuD/w4/Xv7jZ+16H7sSd3hBhFPRIJn1Yruqvn6Jk5wTeivYQla2h/Z
0Y9/oD5rIn4netAhvpW8uaUIdlen2RbMcaaR4mB9LXnEVtCvgS47Fd1tNErz
d6+refS6WW2M+w1wpCtwdeWd0XyEDBNQ8///V68nZeLlOoPLE8McdxI2srzQ
Fga9/+VmqvSpHvOPtAHK8JQ195acHCneHEOK/xm1ALUOZBco99sOnYArZqUI
aFX6kfoWXyGv7VbVbAloiZJdErpthBLF3qW5i0ct+gtZrAC2giIurX6zzVNF
epLCTdDdflx0RbYT/VC8rlvF3GotRX5HXwkSq8O734SU0SCQPC0KVNfqnN2n
OrKRalBp/Nsdu/30wl2ZOLPA9VlIm4KATcPRqakpjvWBaR/hrSa270N2xzjh
JWSiwNxOLDJUUuDdVuw9E7T4ClpYUzFYAKAZQ80gftD+IWN9wqBT0sV7SvIO
cv46Q9qPWkKqJyhR7yXYCxXP4gtHK61RHAtKCw7Znuxk0av8Mv7R40d+PJNm
wKAlZJ15QDB9QV+0GRuQ0+AQL1RYk54WT08hH8FZ40Dr5VmpjMkK833E95Ar
HBAfkNf6CT8kgyd0LKYsLupy85L/0pGRhSwjKYcpf5VDiYxtPVG9MxVtoykL
o7z/vgvjl9xDHgscmHKfOOmSYgY13IXIgyKjmpb4gvG8LSVw1hRLaPsmYkPi
gu6xNIX3pizfT5mGoEXPJuK5f0cUE9vf/hkhzahlIHI3vUnjTHDkL3fv2SUU
eGg9bu1bxptedBKt/TRWNaHNAHwnXDWxbVp7FRGjaR9z+sVD2gTwxkdIArym
JsuxC8xTLK52EUu4K72ygySYzRPQhpdX1pybGkBEGnThzzHIpJ6SRn1c2Qx5
KeoSabm6EjU0e51PcxiPeeeVlTuE3KJjPEVTTXgMLjQP2fud66ikdLGJc6qV
epFDN+kZXMMf92XUH1mUc0GjOx4zTgmtk0ItU3wvHm1TjCkM+BKhTKWnaUG1
AV5pR8oGoEG+Ns12POJgh1MUaolaLVzMDlGYv3C43LaP9ah2iakZaOdhRT3l
KkjO9h419KE6nrO+i+GE3SLOmPXunN87X8nYr681jjOC6ZLNvMiCCXzXyD5L
50Ai1VDGtmxMCnb7DtB8J3VG4QJbJ5BlotVIFTdCar6orcw3a6CJ7l8noh+x
NRAHMgxEYU7qjbxXQWywJTQciqlpVgAo+icRifKU0Xq2jKVMdqZhhyxcNQIR
IuOAm37cRxEWRjbWHKtfkBquV90Mqh5/6F0o32wMPt4S77nTsIOLOfAuCq2R
eYjgKZfqnmyuJmcg5BOFWYJPcz+d5/SQFB0j+r7NEX3Xam7IIrW+T0NfFQx4
UiEaAtSRGdOZbqOEXnzH8yrwMsGv+CWzVDjB0V70y3pAIwqY4tAnUHrOCr5N
GBkwahrLCT6OWexhp0hWX6weYeHiVzVLwhIYuQkomb1HtY8ZK9uLAtRWGWQD
W27IUjkVyDWB2a3APCkfdEg9m4Hmrpya8kOnbsoY4wdss+kk5Vca7fspSkU4
ajHwEWZmHRhs4Sa5dXTVNVyNvTCh7ulEIxZ4UQKDEUOmIvgzJbUTHTIWCGUr
zQse3dOCSivINgCb4zIEP0nZwUT/3DuZ4bKXAgockzsoNvXnABVu7Lqzt0hB
uMiHQgdAoklH8wRVj0wJtEpA9utSUSz3+hXediMopxpHj8ac6Qhns2wA5Hci
msYBVILHI+pt+vnX7h17wX6aXWMTiOzC94T7nVv3ZGGeuOnm2xq48vFnZBgd
hKvzMeqEr50LVdj7XRuyjOk3RdF1bzzICf4cGtRTn4gOTOk6Kfrtx5hRTloI
tEQyL3rCJzMpc+8wNq290QqTKkS/LeokwSKfYVY9tD3S4dpZ3Nmanbmcpt+m
azxTSxCKgz5g/YFJUoYcEXNHx4RyIwjVCaqBKddseJcZhEwH4j300ghgqLXC
NWTr5upIzDf0OVPP3b6Ung8bdKywTK81GfqmAJ433MLDj69mlCzar1qGlzl3
sc8p957vGaXjs21xFTkh7nhOL6+y4NvORKslsxaYTMy2MbqLhKd8j69pU8Wc
cirVHoLFgSV8WEiz+a8CUzgds/4aHla784+pY8oOAZGhsP5fVI4DeaoWZgob
haALO5aZ6jHDnP63UAQRQTSwCK2Wsxnn76EXQpy8D4r4V9WGVooZRn1U9Mly
aKZpV0S7LEIXsqqGnbfgipoips41cJakyrCCuYgiWP7vohj6HQvjbOdJLkqO
oEJtqj6u0FYbQxjTwHmHELkuZfVihdDSYX/DzydVx1JbYwUGWVeyA632rg2T
2nrtIXHy3pN1fbSGW/glkKTBKkqsR9x26SfqXbQ2L1PF4WBb7UCnJt7/q/xd
ppepCWVpc+tDrPlr9lQNLgl3VxUltyg/UoRNptwfiwMqKxP2oGeznqfOOoc1
TpF1r2jCHY7TgM3vhACqH2frkKOhed/baWQEARGDal/CQPA+Gvuyx54S2Dj/
p+c4+2gwiZDTB+TQtAWEEVlYiSWIZHYpY9qSL/OQk1nmtRWLnEyfWM92iwJt
Vv7Y16vh1VCDLcxeIGMMrAnE7+DAeHryzIE43O0hntBk3QTaxbPC/f/gN2hS
GU7A3g8fFYj4lq+HvQTAmxyy4tVifmXl5npi9YoVDrtgGt6vT2q5jn2vLOqO
JtyCLuyV3hGKufUAWCq1MkGZpScbWI1jXT2ZzMyt2Kt5I4C6GWg3cELGAf92
pdWmMbPes8zeWs6Fkxw/kWnnxkEYnVLEpuNorGOYLc7+8XDdqNoLZ6C/yS0y
8JGFS4MRjXoBKP/Gu/buSbdCMoZLVstWRS9n3vh6UNeczICdojTPAYep5bF2
T8O/CTabJ4TvJ8nrGfw9i4RgRLrhtedlAx5Jnh6UodnSe0RN6Cnu2MKXQ7R/
FJVTjMTkkmSwzDtPTBXDU7y+6i6ukCKzkKgHQVzk+uWfeFOrkbdqDEwV+07d
zSGaFEnEKUCsjPAddM1vcyZcyPgs/d9H00tftXC7qTEGlLQPG4srAQPegDCs
BUjeZxtbm79kzKfRCKGpNfe7VcuDzEGEUlEJOUnMdzo1ikrLYSgNKMkvpGqD
gMaB4lYcf4fTfL6PJyQMPtDM1/9A9CaZJil5nqNVB/oUrtWIATywZN5trd2q
7Ups21EUiM8b+cfSiGiGgSeLXOhnJg7UBbc5AtD6xRqsEgIaFlRDx92TAhe+
EjRvRIxT84teYHz1IkIhCb+r6H35PXsYcOjD9go+uW+ZKxKQ2NBFsCzcjdlU
vcEbbM3rODA8SpvqCUsCqt2vQOAWul5T8p+SvMSHlakVmXkkmvzRkvEVVaI6
OUom1tRAk4nNaS8kO51NitxDWDKXhUEQUpd28bgo8pa5+eXKPVBY9ihcs/VO
/xQGJDOGnxNN1d8fnNAynmgCYW/WL0xjd1RcJBNrtupDNXD+0LUAk+0905NP
EYMDCsCCJM6NMNtYhhvLTDTqHXfrqwnWF2RB2ZtA6ThS8GSd8dC7mla2B60v
V7sdvN1i6vyVFSDPiJ7QUh5jRMUawMKlVi/ZqdZqP2eDsPmVty1++rlO3SlI
FJUozfNUHH7Bl9nv37fFby1cipyv7qSJYdB6QlcfxN2bNwXOx61Sjbg9c1Hs
yMFnsN8tkeIf0CqU/4Ho9qmOA+/AF2SrG4r0yEBUQ1TnflJ6LZWRyhudk4Lo
H0MNfujfJNnq2kwBDAi0Mj4p+qDThWpna14/UM8nGQB8hCzx4ttoNwkAeIFd
jTNn1gWg659r+sy+D1x7NeZc8N6GdpmWDVZxhzwv1gIB7OZjrjq3M6tbTIhD
VbFpOfJl5eOciNSxdkLfAkn+aOPAbRE8snxb8MYhKzjbJe29Do35y2x8EHuE
HJI7OtB3VCnoQg8OD1BMKRx0SbJhxcvuECjtkW2aV9are7nOpD28DLVHc27B
VERcy1vjjwpALJ8ab4aCq6TFDAKksR7vX4ykcVvRpAM0PiPxPNnSvL9/hnh5
4Dp5oVj0YyoOP+SaFlw/XJtE1xKQMICSS0ssx1JDHBFzHpCZcSzuCH7D/x6x
IQie3aBEINOAb/jT8kAAkeC37jSpDkrqruXZzYApgvhaQxdMG8qYdKK7iqh6
94Hdjsozz/2gmryd7MZZqILCCNbpRF6LQ0jsz9IKAAacfIPSVwwXzkoK2mJx
1DhWaWAlaqpOzwK1R2fmFvvrocmrBqcfzWl6uXsi2JE/fc/WB8B5Hybl1qSJ
eDuvz0ALeSsGPVzGCfum45BN+sfuvZutNPM79439T6gUPzR0Bj1MPuzvXdm/
BDM5QB1AmQY1/R53pGNo1EpILRNnKddMbK8+ISKcawSPOPT9Pqg4uZ8o0Ioo
FO9F7WE+JrEyx4RY/NrcaLewl+rb3YB/WuzN+dWA52yeAeJX426HQaNT0c+M
cXtLuOfL1JU9hGDuZyI0EdbzvVklFinWUE1WL/WsWGeZW01Fc49KPNs4LB3L
OuvbU/91teXZDQinILfvATqPm+cs5XmEnhqmMwyTCYWTZOvcCTf6ZfPyHXIU
b1rAJYDplTiqvfPpcfyH61w5SWJAg4Jm4SHpdX+CLMs+4TFo+6Y0T2SSX01Z
BsNV7TbKuyUimO831dPgCAqgJ2X5aMKAu84pvHLkvr4hNAX0jzlBnRoINPf0
ArWqTPbmmUbDoN2rfWRTC8HNiyLY4LVLhbHAPOiS8uQilIIK9pOR8MI6ivlJ
8lf4Q60dkLQvksO6N0DK3sa1MghuR7G/SzaXOoUcQgi6Nf3kaOFQraOtOtfa
bQovMUmYTx6E/8Wne8bE6hXYc392aHV8If67+eQ6PGJi2uamBAhvRDfSBNqn
GSXRdTK6zGXtyfAq8Q0xPts+l09mnzblzkRJVFk3yEXG3GkmGkCLJA1HKIqR
qdlqYbLeBrD5qOCfu4VZsTWS88Dc29nIbGOiA6bmwgRROiRn0diWLUr9gIY3
KhZOK9r/K3ZBm8Ag/crX8Vn+tsEyvsH1dmccxPqxQ77GW9paMCtzUwGZnQkm
9BiQ79lmMfdzMlJxQX4iz7CvkhFkTSBcogb4H5kEjPz/zlFylURkGsRQUvQH
BPOhQ50yRlJV/oEVQt8JMB4lyMpQn2OYsKSt8Y0nvZNSPDJZUFJMbwS/YAoV
GsUgPnDSctPjug8xlV+q3g6DriiDkbde31aaS3igV2mJw3nqTofl9L+XcMCX
oqwA+l9btzNUR0qDZHIHDyuzJPT1kUynUB7uEx6LgftZVFq0jKhT3Dt0iX5c
CP8vTEQZMmzeuvvVOHd8f4jw1xor9n+yqpTBJp9jwJqqHOB33kvNnR0AMjCp
VWAaGASAnDfGjkK5Lskx8ffwmb5TF3KEm7Jm1tTWfVjAPXe9OkeLG/A+NNgF
d+9TzJJS54qxyaNzpPrkE0x6zx40qsRW6uHSGvtncJxA+GHYJJTLGTr3Yvdb
QK+NYrWiWZW9dXasu6OYwZzOM9vzZ+2s/1Yi3cGL8RfmGgr442sAQpJKdDk8
bq+loefLr0XYqxprD1a4O41dIW8CaV5zxSzm/0f5IZGWGBwcsEx9dQO7vTmI
JWbGR451Fc5QB9mK6qCdlOtYntJUKxCY8IGYj3gTfAVyne/A9JGNvQMhsGV9
haujHNq710OpdfCk4B4Qf2qnyfiHRCc96i/7vP3617lLEKL/OrKFevwix5Gg
Tk0S/H7FQrCvkXjZRsvDtxBss7K8SaYsKpBOQ9t16aymW/c7uHq0jqnd8Sae
/SKN8zWuYcA3rsnorTdjlNCtb1OLPXjpXF0e+jmQYIaHdyDBEbWdY29fEaLT
/qvZrHPaMs2G7yU+Q7stRSIXEYUalkKD5i4wHg1yAr0dq7QcQH9GJNgbb26A
2mxX3fyPiPTeRX6TP8VKUqK3cytTdXmRd4smKPmTzMNoF2Ihm4aeEqhUp4ab
Q1PrpZD2C5hf/jdRoUInd5eAl6iyQO8MiULQSewlAB0A0Uhbu0dkNxalxd5S
oSS9VyKlAUPA4jsgoCgGEoKE9S2l9V/7MHuhxSdt7mk2I/Gt13DvTJxnhOb0
W/2xESgK5d9sIO1k65+McQNbgFo4W5IRhtqRXNjeTHgybAmteUCAJvBODRE+
SSTUDd8h1+5drcyt7Q5NhioFyKbplJCGgiJVftMYmpo2Gur7aR5UirPoXfU6
bs7++HWPeNC25aAMOntVrqOEYCHOfTVQaABUmgOsEn+cfasTxH7bbvNGGARO
T8JvNAJwXKQpjy2vHeyDjVMQmjqOTZ3puBXyoBMV3BrTw902AFMKxp65PzDE
rGMdlRoArEqHNMbO+WT6mCCFipg7hd/dKfNORWNgEea7c7imyn3ZkjqIi8lT
NdQxJ8V4ofETOgfYMoDZX9FvdaMQBKIzRMT/FGTtLsM27bWuorM2x1ia8Ohh
Ke9A7T0l9n7CEXEiTtcfUoTbVjR2+9t7cVDhwOrtAOqzVoAjdRVB2Nk0oKp4
Bd2QAaKNcRvNlpXr4o3CQZ6mljppUJE9qljGjV9Oc5HteL6w89w0cBbc8NRC
2qaEr65DQirw7Bl6qmuh5k1a7K7plkMxZdNz9anSX4vHgxmm67Vdazg1G4Ko
UY4QwOSwSYy8UTmN4oCkQbEj2QthOoDFGvLVqFq7MJBn76vDWLib/ioXIEz+
qVztvp9y5dBRCCwsZI5qHk0uGQfAKPRVFdKlctY97GzyAQL+o2n0CgBdXovk
ZhEh4xpkN0m5xK6uN+ztse2Ah0FUCiA+/1TDnBhoadg4CkL82uMp6XeRUMb1
2zjVg55TxKxRrjO5jNQJNPLFlIB9Ouf1i6RtQvSMzAkTw+gm2gXejFwLOozq
0dwI8oBcxHcbW5VP8ViJ8MdW3ZnuTY8zXxxEshjAMB1Ni3VDCmR6ZGwMBITi
lAAoCPtDHYctZHrwjH2y+4WifW3RVRGPAHh8i5R7/oGHioW4VT6Bfm6eBLhM
/bM8sdjAb4Aa+XGfa7ZdxgOlPqfPI7AeJrAdXWeCglAwT1K6wlJJzm+wVQZ6
g74GW8MuVT4x/svLqf272iNAT/RkCxGVNzEMcCZxPTieNjohxAc1OeAPy2gq
rfGx791LGjlzXliapwmbeI/aXoSBRbPDXBkmjil4LtlQucXBiqz1QX6UvZPL
+bi4kYayZv+kR+mBZQeBtHGDVwjjfUYYdy5ksXokUEl2B5gcvV5JYqPDq7Da
+Q0M+dffJjoldrzuF6rkf96QFacBeg+OIUb7gietO11V0C9mJMzSTOuIcplD
yOIxFxY3yceyX2jXUFAr72eYKxANydw6e/9s+QG/eZeS/HClcZy6CPtscTuT
5f0DTV0jdm/eYIGo4Cm2QRCem6rKN95t8HITNfmXeN2p6XyCl8ylfLXyexgN
42k7Qnmnba0XA3dMkjfsVI4LxrLOH9dy8JD5nqzwnNbRlHzGPnyNLIzlzHqi
k31F6xsAE7LvTnm2uoM0Y8PRbSAJndxM/GTJ1ohqArKh+5I1FIEVX3zEjatC
RMotzTQKtae6L2vRGkYujP3gtW0juEJUcinGsb2Se49ZZ8XNkTsvOra0WrZI
wUK2d33oWLySdWu2LIt7G1LRCCIf8V1QrL9dGpGowLXh/Cqmk/mOndGgtfcV
eH4FSbHmCLEKCirdfz9Mlz462HrHOcKjz4LqCYuBl8U654xK4W4mFh0g8XeO
mqyovAoso6H3ckGstVHdoprRu04zRqll6XFgRXDrVzKLQSH+M/+h/Fs3BEEf
anr5wNtrI3KH2nQMpJl8/uqg064XWQA8d0EqCQdT+0GrmrOKkNoGt4uQtU81
rz6sBPPq4cfuqziEKrnObmBdJse6MC4tbneOHrF+IfIYPMIX1eFwEa1yRsGL
qEAC6etULF9fNtUH/+qEQGHr5a/Hh3uBS2skwhQMAtfIgkZaeK3J5Mc+tpxs
BDV9M7EAXnrpleLpC54AZDnyo5NHWOE6zr640DonSI0BpkDjoVPrwcXLzhHx
Cm3M3Ltbvy/UDKoYH0fx+DRbr4yz4oMxIdyib/c0IFQOZpELW9jtQyCkbnhf
B2Ct1Hq1SZ5kLkWb/Eh3Sdws+897Ta2boLqd2PKrz51/qXfVTfzKeK7C9s/H
GY2pY0a6VZYjrWXbxArlkQjrMeDGRWdPB2HUhabHwhWJDqsypUho2h49cPIj
UPN/kwFxT6R61e1ysXIn7vK+6HLhS2AQ4LYyOCflqR3Z1REN6sqVJIKx+rGA
K++fCtVt1rSTa344khlQV446dQQpYXalRXGApqALvzAvy+8HZ7duGqbkyI/d
fDkk5TKjQlZwB722pgKKyg/Wvj6tGVaWdR9G9OpjiDWQj3miXNuiUhZQSfnP
IVHChqshYpbDp3kIjiRwrMwJpV0fcQfEz0qMgsS8uIti+rmvQ13XJGT0IHEU
Ha4JmhvGehp+NJj0jt2xB8ejTzAgauCS4fqldZbmdXid1obhDHCoXNtkhiGx
OVa4Sc9H7+xC7uM99oR8xELxR9ihB/LIZzWzZm+xpD0e3YHKpRSCz7hT2zfu
/v2JfI6JsxR0qDDfqytQ2R7MH9GgVHmo6mVSjv1/spOu3yYPmGTSVv3a9Ivw
p/aVcsa3kRaMrrUkS/PLZzAVg+hHLC9NLp6e/NI72+55Ie/xADkDXz1d2efX
e98KuMkBzJZft43eh1jrezKsPefoGWXjgS19EXUZwwGah3nD3qPGYxpOhr6G
3TFizV3JRAvo6YSuNKDTPIhtjrn9YAX5wmxZxhLbnAEilzj77fnFXT16ZsOK
uWVFRozElOTAyiTypvMpO76NzDbJ1NsZahbKNc0eqbr2FGOCfTkwazT7U2mE
6zOuHTsNKCSMZwKEyFERIHBJeoGOAJsLqSb9WzA/bd1gZYBDKYJrMxSUSHR2
a4hr/vCaTlw2eGDVru8qBWe/NYJnbg8tfHf6690fQOf5S5xZO+v5HOq8jXV4
EPPmUSXv0RbUH/PSehNlW7NcPRhq+fEzId45f/7NbXyNwLvuO16q9Kwldsb0
Tt3mpjeZndUSFlncZ/g20yZQQqZRSDGGsEpkufQS9YbFJhb3CQP5GjF8DqaR
k1R1JF1prOz1b8lD1JIXTDabYXRJ8dDl9/DpLismj7IDTjYeoHbGsairRHqD
HR5ezFOte+gGj/KItdcxYZ8yR50vb7ehxV6M53eRKk1Ts/cwykrqofWHJ8bC
ic1OlVRbBJLprvnJETjC1r5xODPh+Iv11K3ZDXNK3BYLdm7J4HNG0P6VroOT
aa7l4ulS7fV+iioXG7vI9CzSKFTixUZe61QLEkS1ExhkeGx2jpQeIugnXG7h
Ivoe0qHj7nhXtpaT75Fm1Wl6C1VkV2b3fuhgbL66ccY5R2LsQ8SVPDKkKy4y
cnAAEx7dgJ+7irVsANHZKiDeBNdjR7Vy7uUT1CBHXsLNVXzhT5zBEzVzpr4g
IuBtUbQGUNJ6vwzey2I8H9Gff2D9nxT8LwlOtU7R6/C2NlVSbzFvQ1JhUIHc
zlyPgwEsUrf/WH1J14oE3qrN2nIzM6s6E+KSqbgkaYgTlS9QbJE3hSyTkkTx
qXi7oZPh9VOzjhs0USJjVKEY9JO++3rUisavXc2MP0rNaI/rIxFh8G939BpZ
yCEgOu0eiJ0y/f20gaaFxgILP9C4VCa63W8kyRFjBchBCSZYEu6E4GskPxeC
YYC8gWFDg1MgG4cQ0d0y/0giaxYg40Q7+94VFvto09JkhwWdzo5Ll7PDXb+T
aC4MG7sWfvfaiA/244c+9lgTgsgClLmlSn8LrJ4lirWIXyijJvcNYpwnaRSI
kcU5rq92z6YdijXdXpbgNLDDowpGpYTIPzNNibgKqa6Sj25GNxDsreVM9jy4
hyWFXtkv8xuBFNVR2E1mM8W/cGjFrz5BleUv8HTf0PAllMvWCYoqafHN1+Ch
TNBgRuS0YQidyP4j67xHw1LiaB4xgumwJoL6RSC0XDJAUzsIMs6qQ2Px+czx
OCqpej08ierAegbCWzrYOuf/C4fhM8iVDd+MQKJg7ugaJqxFOCG3T4RC5fm6
lgWgkDPWECYQ4NxYDXybdc3yaIE0BTD1A8L8rTNktE9pQ4rGKz3NYFtZpVdJ
uXLU3CN914WzLiJArw5cmlOdFbSteUx1N/YopBjfoajUfICJWPcwQqP8SB9A
u8qQwd7/uXe64z9oJmcvsypq7bc8zmARYtzL53FNI7td650k3rdiRM2wbcSa
W51mmZ/Jpfpv8TSUDk2fKawpD7+0hJKYQDR0F294Q2h56Rw72gkROnRCqdgx
usZi877SnJTjdy5pKPS5Hmgi2wPMZF2cKVcpTywNhvXsqRl+bpx9OH5UFCNO
ZuyZZS4IUUgBKQk0SX3bJDpc6u/iQeaT/JpNSIIDyYRivzsOEUle3w/RG/L7
KOa7S1xZS2R+TzlCmkUs+njpOYAKllPqiZ9YMiRL83sqri4lce+MRn4+S2g0
oATUAiBMRWa/freu6t/YlNdLyotkW+HCnvj4j/QA+jUVZN3ZMjgIu4chFuOE
yxeW9a/KdpH5KyBfgUQUcgAzbjUzx2/8niREfm9EthlvJjZYdk6xMhtja1Ir
XuN/7cZk5ByiZgXwIUiF44VrxgQm+wvRlh0Sa/PjARwUIJ4Rj7+cWpSR5w5K
iK/oiifvUUAoTYnWnJGWWJZcpaVTt8vxOQ9gUOiB8GXmz1orcOWisWRB/dQv
mU6a9/Aw/azETqKOI0YeokbdhYF9Obv94JwDeMICqDmCaeuqWsyXvXuPBfo6
ILR8r90BIRae8wRo+mj8d9bvdIwtkrPhtjQgZdlL2qIE0TMZ/gLczwgON/Cf
dVFjv/2IHlHsZpkOqbFbSxiBwjF8rVWmkby+04gOieAjEfNz6GEdDJ3IVPY7
M+VYwBD2pBfdmYf+CTiPzQ425FJlsImnIJZ5jJzIc6dGXTBUp2eI/sb6tK7U
IAC/9d6Z8A4WmtPUc2ZehNPiPZ5c/NkTG+8/vJn/SboQJP6YjKYqJCDq3Tx9
x+wNZyKIB3TEkp3T/12huJKIInLdpk+xBodOxwvWACZA4VuKso+z5plhpsT3
TLrFzVeBykT5foX72XU7Rfq1q8V4YJFqZyk913A1clvLjYxxX4Mzyolau15+
NHTYuPhlHLibxGFUs4tZdWQAQF0iRV2vyyDt8nwYEbabjB7UAPYTb55lkMF+
qyqT+sfnNa3hspqb6sTen+G+vl3fyAZPeP0doBUdwpWtkf4Ba+29iSwsvtQ+
h+hH63WDvx7X+zZHX+lSWQLVTUMblv2rgR1+rtFttKmSscMix21hgLQXWYea
uUjKMJvtFejQ38PBNyh34l3bwEm31+uulxkVaE4V9WCu61cbRufPffgmL/4Q
09755PDOXq3TM42co03O/2XIk91XK7qTg4S4vMA7TXGLkbGk8ZFT+/dedgac
N4sx7czJI5MJMlBD6lN5zI09tVkFhxzyYD4K6HbYL2CmKjiB2kAvQUjxSM0m
15cYm0hIbTH02+yrUvIjR5NBRKPQSL0/TernMl7NH8mh/AOgHpUkKEFiz0rz
p6qilEIXfKdOy4qbmDsqDj0SJm+/615xw3wFe8babDMdscomt7fFS05mtmAx
X43tlLMvzIsrreOeMDc7mGLc2Uqzw3tyu+nIxZ6joizwvfvMA8H+raqzWAWL
OVR1/AOGk6K1oYK7JjoBEB0aRO0EOVgtgnrlXjomighfWSqHNh7O1qNztZu0
ddj85jtfuPngc9yv33xFT/qC93vaxmDV7Ty+d6MQVciljqtNLjLbRZXZZdUz
RptpzUz4Z+X1qohC7YA9biMIwr3NeZ4iIHQPeaPL7b/MwZ+r4V7DAP+FCh1m
CDjEYLrwMMm6BuQwT7amwDI6pPhHcTh7WrlVYovD1wVLapZ+bE1T89Q7YZCC
mOHkNusOCOECzciwuobh4TNh78kDtr50NB2sAwg3SSalPZS6xojg/fb/Xj5x
gkh6fNDXWm91LfHLJTatXGZSIkvwQy6yrMkX4rQB2zah4OoBtZpNCRatVU5y
cbFwp7MJyOjTNrHOOMBbhqECgbamQzDOmzGvOkcLT3Dd1HMCCV+L7/aMFsdn
FScf6F6VMnk84uM53/YbcFQbmhunp3D+Ckf6qKN/1z6okujkrra8u+tqtzA7
S+LskA9ROjStpWhmbnuEUpkIXD78GjFBPGCDoszXC0eTcCfxv0RJ6RzRzcDC
4gTnrE/4q1vGo8um3yTSVeBUh1GyM8qoIAsBnyfw/lzYIVS/+3XOmTz29yhB
o7piftza19ss6DtSoJiIvahEQBOZ+peN4kVNID1X+hVatEGU9xAvYh2XOybY
S+qFIFDB6w1NhYFigJvFjD5+PJPPKGuTo7ifxE2eZ1GvFstp9c6HRguj+mum
klkamSZKDqKl4oN9lE9rgu+QNjABcx2DnqFpESHtLV9O1u8x0jlTUL/FPxWx
96eYHLUMbjZO7bdhDulI2nacXeVq9ceZAVCVNBbuVeTnHHR1r7942DmWv4+w
Dph8j4MgZFSxMzGiu24ZxiAh5EP5SLB/gTi4/lS2sBdRR/0L7yAVFLPT3AhD
Y2piE9HYvumo8NF4dMwQD94JabH/Be3L3p5ko+Eytt7Zf8+rP9pdhpsvsBsg
XHi3h5d9UY2Un+2rYqOGEMjyr1G+Daf/GRgZVXOkvj1RfRJRFfqtotbCfJjK
Jxw+vnlmCG5fWFPeTgIjLp7GFtwoWlcI7nr/WEdmxIfwWWoPQCF64irKPo+8
51XntKdzuKusAHVcwZ52Ejl1+XaMyR9jtwXYvM3SkMAQyy2e1MeyPcaFy9xe
631c+JmG/5g8PaPryafcBASrPBF85nCdIv5DssH1OUD5H20HlvAHPdP2o2CO
BhR+7m0Y5nxvTi/xLa9CQUZMDrcEGKJlYUPQcNkSWhrJb5IceYpw0bfEiNx3
z3ftko7NFm3ZNa37tiYXIVVKrZKdm1p7QpXc4MW/FFrYVYSh1T4dAiVxFQE+
JrlIR0X2gPIs5CUak7yLkjHHt1mMSCWx6pM3avhC8M/w6vgn5PLFUqgvz+Sq
Js85/6Lt5IDFRxWIYKF2BBjPsWNw6bV9oJ8qihRDX1JvmHIZ8+l0H+LlXzR2
J14KWHXmlinmGvwMWXte5MzpH3sgD0R5DLPT5QPLo89j1oSccxwBMFjVMQYW
QSPC5QCD0/4Ce1YoAMWqWcisGpb7tedxTjwlHpXUwCKuHHY4fkvare7oyv3F
o06nCE0maYTKdZC0hOkGwmR3Kv9YTDw1eXztl8WZ+JFJWCrPUASo5ljtIYUN
VOf9Ogvi1Px/SCM8pMAC3o20h0bQ+iOr/4BGS3YRnNfPcAhBD53fB/horVRf
cmOb9E1ChPR9Imi7fsEza/23ZBPdaKFPEZdST63rqoUpS2Edrqj9FM0lSyqa
TEyHKAnZdsUryol/LZteB8HI8B9ZIwn6VxrS6i7wgoEGWx8sqHfGesvRvUDw
z71SX149tvlopfolxwLY2y+oe7Gluji+BLfxPmCAYF+3J/aAJWGr6/1HYpMJ
AMgvLdyJHnMxS5uc7GC/vJslNK/blek/XJHFPeMZQhggb+qKe4F5G8H0seIY
4yRnhGb3N7BLPL0DJbDsPqa7QWssVoNVS4G9J9WxR4EZD4H9z8frjyogaDkr
eNk4bXLA5lfWteocbUEaW+vPj5oDjnpl+iSAjR2k0DRC8RGCKkgmjgaKNG2O
3YIYSwQ+/BXXwzKLkzoSeK1cpnalDBwcTwlwq9GeKLjtedBzkr8JR/nBHTo/
mKgIUGsPneImlvdbarK0Ic1/LBDZtGFMKZ1Ls+xj08t2N5e7b9KvChDr7KZe
uVJWQBLWJwi+BzqKrxoGM4ATs9NAV5yoDhqEwyJmMM8tTnoYEmKR5ssjHLYa
hSIeHDkVp58hkwsnZKms59NzP34BBKw4np51NCDjLNIWUXds0hhJADj5yelO
J0O5HnyfkKKam1SyhC6h2cF/HRoFnfhb6fzy84Yi7JKFtJYm0gpnIMnfSK5B
0y66yo4wEiqGh5A9sRDdM9TmYEZyFoLI4k3Cw1Gngg4aEhKtj4mFeIXhJf4G
RLkat5hJK+20Lc0SnfK6ypNBOam1DWS0pQBmw3zPSi3OYFHQgtQmoMrKQxbe
xZq9XmNNKgRWe84Vkn1WhOtfJQSwZcxGyQkixQ3NU2mFsHc5QQu0VBqhcfuk
PJoJ+ZidA9KMwmToCDzVzwbgXbYv9r3vBylyJIuzTTYwFZVKJHL9RjmBWdql
XyUwsP+2NcgYclxyegMEFh5TnWMU+laI0pQeGREYc5dSbAVk3R4RLyOxwZwX
euHyUJCvtjX/pbCtK+8xdOTiwjWJWB0VfiVhoe1u199mFlztDUqD4YPGzETe
3xg1le33E9OmuKL4i1kb0OwgRA2Vbxs74whG9AR0HT7jefkfVsjslHtr6Y8N
BDDw6/smBe1SYZMQ2eAhk9rFMNsUWUJDkBU2/b4XKbAa3c8GHLsAUyTFKK8w
vzb53ytL8NEz4mpX45nmJ2V0vvZzXwqP6lfN2qD5SAAZYdHNn3vSMMkHOW2M
JFZqE4BZ8obihVwdZ+VfLC/v8GLs9rKEm5ly5TXSpDXWSi3KUnFBdvjbxcWp
0/QWtdGdQIK82TAix7rG+IbLHR12wjvtZXfk905CLHOgNrsKSKzLuXbgzFLe
7ajkfMsPXbIDjBb28I3I/yDwmW3oken76L3H+h7I0g8lAQFUzOBHAeoRf9qr
nq2ZC1d+X3DRZ3vWdno55ovpp2imcAONjeVc25csB24xVXRF2QNfrmG/wDnp
E2enHOL4zYkwyLGfGxKDTLmVT/JsXNH5fT+NmMdOb0Mim9rBDITq/SDoFYa4
Iw9vXjbbhszxEp7tDbA7XOBWirus7lWA2AiBHn1Hvtt9X/1qvWm8eoKexCed
DJByLVw+bjkbgtZBg7wEjS7ABJbvZg9Mm3vhGe9aLU+NMnzXGk+kOzk2Ojii
sFx0GQOTJYyzwlIdU97jWyDolLTjHAHmgafaNlilFQvbXFYGdyEnJ8tixdk7
wwpItKEC8vDJKG+F2RcJV6mZBa5O0IWz8hzEnTnALNlcVnlQsEeHYnYkyeO3
Pi2cQht3zhkRHjmOg4Ke6x/7WYI5TmVP4VYRh+ibFdLFCBK+a/3U4peomGkq
JlJlx6mgMEis13iXGiRe64LUN4KzfBn+Wmft2iboJL9HTUHP2iV1Zij+QzWU
B3nZUxe1rXkaWT4at4njOcLNz7sFB8NR2YYgOzXruqGEpCITy/XbEPlFe5cQ
M9XLaHAlGOw4XDGxQfN9zE4wwsDETJJ56Jlr1l11ZCYyWtBvZ9OEJTR98MQJ
M6zMW74beyazjZgfeh4mR3GHy/ZD2M/SuMyUD7VqJmkwIGklfvN16cXxOKQU
9F0WRAPmsD73J7JkK15d7G7cdpHXJy+FDfdNXwJk8QW608W1VaCcG7WZGkx9
1A+Ms9b29FvC+mNrfFoQuV7pYF3TfMNV2Vmqu+n3KUKH4KFWYn2EEo5Waggw
TFMuYhIiS8zBrbP6+kFSfPpF3kMN7Zvxjx3+jKMb4guSEd/GCnBgdo2rkJCW
cAI9WDF3CaymdViqViI3SxfaBvD+wbuFgZlIVPg5MsLbnE8dnWV1pt7WQmyC
nHjyp/XOm8t0VuWtokAyZ27ad2ezslj7MN2h0TvwLw9rusJGBilfQEBnGNfg
ucRx3y0L/pAN4OqGw5hnuJy6dxEkyXOU8DzmK2fGcLHHKor/Jd1BJGFSu7mn
LdUlYKgQOrIVsoM74KkqJi+JHlokoffkcDHDbLWVOG93PT5ZaTrowySovXld
ereXgVNWsGE55HUfjEE2Q1tu5GrxBpBLH4gfkZnr57isUh60Qr2ikH/r3Bfr
9XDnyu8cHPOM1huAZExWr0r8gNFi7+L2XiX0hGCSLMlxr6AzBhFdjiRg1Pht
VfdQQhrhUTwuoZjZmsbMEW+Gx6MdkU7cezZ5JDNt/SQFkLBg1M0UoksYR8NT
MK7wOzydS8r63BytLDYYxz4rvammABMMDvj9b5iwEdL5JhCl41Uol8OtqG2w
eaO5pSHCSMeQYxK+coZGJssbE0DDlhllRiri8IZCVopYkqXPZOMPP438d3Qc
WOtq5usbDKsOq6lraXpj2Rxz3V9W7ZjDyOms31xBvaG44TyhJe88HnrbTiEB
PW5irhZP+o9GfVWPoS+nmutk9i3HxVu/S63ke9K0YrAbFtTE1Aj+XUVFOD/L
t0QZyVQeaziGhwYgtVVhen1KlBPq4uUPxJ7U0xVx+e5sYHhE8MTaJyvsiNao
d+qbGXxgHZxL7LN0j+xcgf1H7JUglLeeJgHFXWz6UjanDzY6YrcJ4t/xEFUk
enJKeqe213BxnmsGJ7XGWl8l97HHwzEwdt9jxoM5fBRgblY9bYX+VMoR5AEZ
7+CVNPmpzwKaYpym90quIbq68NLiJ3wOzJgQmqujXqDm2j4OuPMw3uTW93so
+SJFJACHLvJ2ptWNqg5zLVgj9kBBBof1+LatdKXvKr/XjLne212eKr1chfnq
HPKxW7jF3P7Qmbc8G9Le8XSLK6n9noro4uShmfsOskinqkCjlLMTTwKk/cgA
NlqDaImJ4RejM48YKkZnzczz3YpoT98ZzV2FEmFfAzeGFEadsfrvI5mWnm6e
Y0wPFr5/XIiKQ3NL660HpPg0yAYG/+VcabG9IJaWaV02CM6E0hQ6OhrtWuD3
4hSEL5jXJtT+vJKakiAAETA7riIphaZzFYCcg6stVjkZuctpqoHtI2Gy1dl9
guphwVKrULz16VGdUJLMOopNAWjaEI+0vpPFBi/x37Ws79ZRFijyhlfZ35MH
CqZjftLVOvkrvV77U8AhHrfut46+6Pdk2zGyKl/Zn3omCJnf+7PMRSycxQ0B
lc/z2Cznq2iOv/le6KXNmb4RL0Z9ThacU46CyKhLHrrVUPL7QsSxNAQQ4yQb
o6rakq8y90/cOA5eyX+cSR07PKFKx7co0BVbyICZh/VZZUclDbraeHgjv577
5us0Xsx3VZAXe3UojWRk4CdOAHAMWcNB/bpd9XrPwxY7C/m8BIj4TcRVEtAS
882g2lExvDZCxWnuK/dMG5Av5/D00L3LDF2EN8LKu/AQfBICJgo8B24TQTlr
/KNSBuGS7+X+FC6VtW5ac8Gv/B+IVtF4qlySi+ZfhQeYMC43udiVxrVCiLv5
lKaX9qUNzZRY489qLMuS1pn1JUwRTgtLZl63MkoKPd0YJKMDMmrKclZ/8k/X
IugxfGvSDlY4lPXLGFxLGAkR7A84u2+o55aL4rcNjcPPNcKYe/TFOj7lVL2v
AZg69t9SwuctfFDzo4dJRMebzUKIIXZmL2dmvbtx2Z+1I/hqDYoBcL0cj/c0
VQjS8g5jLkNYhNOH2kRgmNcNn6GV9ZLmNRcQhYsg4deaFpOYi5IZJQRw/q8l
mbrfBpsn8cN5OfuS0bes6ErSPXFs4Ts7T82h3HdrMmoDmLG+LRMnHt8CEqbn
Nb8/JBnODhs3lFCq/bEcqhpjfqqew0dgGOXHnV5A4hTtJFRFL8w2hEOzmijC
zQSn6Vrd4tZVaIRrbfxY63lunTtXFrwDyK7vTWHjNeif7Fsp9evnZvwDHbp6
/ipprbF9qjna5QKl/YJYJBu2aI+tK9A78x/rtBrCig9ohHaWOparneeIiFdV
T/f6hSOY0VrXmY+CbAn1UPVE4WInKknR+LregA6SsJG5ijVbMlWDHEVO32a0
tPCpivmrjnvyaiHssZ1cKa+Rl+o8R49fJu9MzUnoXQ5H8WuA5+AiP+sxaaOR
Oa9pip+inIdf53mcNDjGUXIhUt/lWDOcbTMqDBzjJj3YZk6K8zC4fpzUjzue
VLQ5werSL+aRnwb84ehDpjafy0x54kXkNLM5NdR9Y5H9MNq6fOHJC9g6ytOZ
FVOX+qZ+eGMpbUJMWBNTj8qRXyyiop5s9fgOVhvP/7wnscZ8lji4hY6uOU5D
MPmql0PAWSLejus6G8euGDg6Ao0tjGbJGL1PuPWCpt86W5hnSdwT+ExV9n4z
QkgiCcpDpCvXFaA06ElI1+FvCC2U1yuEL52I4thXGq/Eg2s6FeTRfJCp8RSO
9X9/7N9gYbfESdBnPAZj9r0RZlx2JrWYlb7dguVeb0h7yNgRbY1GAPFl4fz/
Iu/Mo2QLlRcdzypQM+sEwpcDt0d9bE7S62cKhCxqEXr99Tmu1ktGGknN/ABG
Z8R6/S0DrwBpl0kGor1AJhKS2/uucQ7Xw+d852uoZMztnid/BMNcvaBH0lQd
mdz6p4D02eoBxQoSrg3hxOcHgZjxdGAu36twaIT9xvQX7+2AjRuKlrufMFU3
Pt+6ZNGtzrcmULxQbJQqrmuYc+C4ajxdDu9JTGmK8yg8C44uOcKUaebmvDsQ
LqQuEHz2RMrR963nwpdMjwpEDH9FQYrsszYCU11Lvop/mYr3NpSE4x3vkNOA
OSnSqigzWUidyD1iz87LW1tQZK7v43fG8l7opXZR9I0On2lBdBBAhhl1IV1n
SAqTXcs6uBU4z2xW+JzWcE84IvW7aRupRWqtL9srlZm7VeIideL1GADHiK+l
m+hH9aWeAXWwCElCnsbYvKE9J0yKE263Q2xDfpt3BeH76RcsScOcnZLul9r7
OCPVJZya3YsLsfRtJYUTo8nHS/hvjYEyy9DuOhAPuZzpbr7lJC3d6pxy5ndt
T6f5GqDZoXdfrKgIiwQPerDilTO6RoP000KFsYWSe2hejaWzqAconchZaXTw
QGePK4ZWVKRAPXCDegTI0wpgcuWoS53a9biJAgX8VTXCx3KVzTFoAARUPD/L
ZzQh0cmRWcMDUZEP20K+QAlGVCPjrzfIPyYa/eePXT0GfpCLCSvDtollPd+h
U8BnvnbZ3gCNdOPMrnqcjb11G7tt1oZHYSyrF/gq15X71/Jpu8b/KTvXlqGG
IBmjNd7t4tdOQoxqYo7BkCQU5yneojCB0nkQmV/ikkjHKQMucM53Czrw+b4X
65L3JjXvv4xBGa1PAnn8Egj8dim5y16Y3E3pnWY+AamI5ESjdetg2FbwLEi9
xgZOd7CS/aXea25PSlI5pMK+iQy2HkNdd1G9OeJ5aIKEOJBGNgZBiV17dG+f
MzlI1j/dx01vLyn7uZKPc2iQAXwJZaHutz7gFOuWqS4xmratFgux7Lgrp9kf
8ohtR6ZgJK2QLqOp1W+cW9VQJ1uQ6uKF5Nec1omNx0KQJbPpS3AppUwRy0JB
uOmXgaIxr/jMvQFWNtX0eXyovNhOHOhXhJGF6l12Mz2n8whO2dAwhJd1JZhF
3SvRwuQt9+cKwQiv93G/EefvVf0TSe7NYOudVbkt9EJg6PH97yljEPj7cg9K
18J/dZgacQLoGBMahv9SGF0vuJBkQUQ/07jxw9zMEeZK+YzCWpgGrVyYz9PF
r4+0Sf4ImO4FBkjSjSPoZJngHJOufm1kHUCfrQDIF7e1evddTPRwt5NGeUyz
6kSYv7XtxCy6ag1fJJY+egcsbpKDg0ISYm9Z8heDKkB3LgN+jNgyHW7pp0+i
7t2VR0ukHVnnWH5359NzuEu+1TcvzLB5nA8xBVaOQvwB3vkxaIND0BWUeoaw
hA9J2PEsVAGrowh2jld3xHhFoGs3MJnEWWdnbUp7oPW8JoqKAtp1xNeJh5hP
Y8xGAb715cOfCNTkjVWFf/lUiCk5gGZZRFdtHOCfWK5o+99zYLyCQ5eNVGvy
Fkw7ObaeBQNC07HtrKp5VnCg+R9XVak3twChHbTT36G0HFMBegr2PLkJIN3V
qLEN4QblcOd9eRmyUn8MQ/WLwpNQ7bepuURLuOPG97SXMacw8lF9rmdXz7fl
QOEimNyfPRvys4C5JmpA1WbZmtmmezVTGsrTjWOlrvEvHiuD7NR5Di5VcdMi
FMrIuftAKquRQYKfQdOMh/3hvON71nO0xI0SS0cwcEKuJft7mpBhs9a1C/75
v8lnTeXfSyIFtViEx9xyRYHPu4SthrL3Tj/z4T7u9XXb4tyVTGp053maqzCV
HY2eddc/5JTn6fBwvHM8WQjuygXteDIQigfE89q3XdUycvo+Dg7mhBS98JuO
ceNypiWKgCujeFdw+qV1nn8Oruz5WiLyNb+pacyhDCFmsT6hYBUYNVyw+Z0+
GXa/NYpMDT5eQRmgKotu1lFtqDuuvwQN4cDFl8xiLQYJw+UmJKSZfB+Mc0av
vLe91dl2R6YtYuUqxo996uMNU1sCJy17aFDNiDdQ1NNGPQHPIIpqNGaEuXdl
c3649uaDjUBRsv4V/5+HRPAWcBQu/Y492LEh9g3ce1xkoFXSC69OjlGtN0Hv
3F2nd9GYlFZqsSYHLT5QYeF6VpT6c51EjRixvyuiJWidoV41rzX5TpDiJJC4
6q9cpcPrto3u2bReqRe9/8QmhXY7L09G3h3Efl+TVUGtGXNdszduB750lQLb
1cV05IQ6ij8nTZEKuwekmT1174BPqUK3LL0+epK811+mQQmWKLitVJ5DYLcA
t+mYSXOTKZQIiOyotvTqJ0VgJ/OkwJ+984ZgMPH3F7Z41NaZiGuahbp57ife
rLdi7oUqip/wVF9awoHZMqXI/A8ulekpHJA89A2Gm69YFar9rCmpcUyHY8MF
cm7fBw0pa3v6zsv3CNCSKJsoakjTYiyKRSDLsGTnYgqdwiZclS5LrjGt9PEQ
6LTnGcPGR0vhXy0egl8PYuqFtIg/O//VeqwKgDcXuUm0ZmgCLjqXYsbvqfNl
rmYZcIvJDMXvRwLUvY6wFcVPD6gnr4nal01GXcI59ieYmXahkQxbVRwsE2JN
Vd+B56oqeRq4BgkOzBR9jqYmGgoyBpTWRSKGKXcqby6zjDDnIM63d6gWUs0x
yMfuIxQIVDOUBT04FISdyuMVHBQa2dJaemOCDRpOxom4d9XupStRHwdfSzlz
l0R08STWoykNni6z+286IGeVir/mNurOYfijs//Ist5o83A+fnAkOuK8FUXt
FCBE428a9HYcqI9a2m/pTCl9a9BWa2t1cq/3fjzF2oxYpUZ/PaTp/zHESNbq
nRiQ6y3Y1iIRqPWfwsGfQF0Aml6QJsEVGtJrSbeCtCP/9Q5oX8dGLkMQ7VQu
BWrNxo773WiDIccxnqgBpMULZd30bYUEWO4AOCj5W8czJBhi8/e2V0+Y0CDx
HFQWdiYtW0oPjxkJU0prskA9HyEwMBMEuNOfBaq1j32cNwdS4wMqZGSiKgLm
DjUa0/uexONL+O57OEzWQp7aiBYRe1TCMBADnvmKB1DkVEThRXEOaEc91pK+
TZCZkkzAMpBGtByeDkmS78UGE+Gz6+piuSPO0KlbHbquGdEvO88YLli6Qvf7
xMScbdM/NNuK2xCnV96FINZkVgkcBDgJQ1ndqmRTeew+KF/1EcuSiJs3eiyj
FEfUaXsDcIQX8N7thCcqznvvqSpcq8AXt/GFNWl4YNsRG+y7r1tyJtoWo4YW
R5PcuGjelccW138h7mB3sTV0zo4DZypC8Crudp+/11q4MQTCvupUK7KjG481
3b0dd484UMhXCoB72WnmQyAygcNs7NUNO+ZZJpOITTBlev3Z7hSfE+cNFf0K
rT0qFkk/NiNA4n0ZKyvgoTFmGsOGiAswWET4OaKX6iX9kyOkTmonlfskwiAM
fV3HBbyGmm1kRTfxuKUE5Gj9uy1hjcLvVs4VdCH7ZciL92/6ctUw0gVDMS/o
sFCFU4ZAOeOc6YXkVUxx/WnFjc0dqvmppsrw2Tr29nsGOm9ihkpOUpUBJifu
B5mUTf/8W8uUBELxMy+ItrCE+hWtBQ0FtovTqsJ90JrFwLO27UKgYwDkwohj
f1ZWXQcwCDYHDHkWf/5CmFwEJBq9gG76ohAvpPQklWM2yCUhJoBLpwlpdqto
G3a6d4k8LBKWuB+m0Z3io7ICVe3bV1Yl/+1KltvUq7W++tCn3LXbkB+aSx9B
BEWfAFxwjVxvhpQfe3E64Kg6Vy+Efoi4zh27sD5SLL8HAUTFUqf/tGrI11Ou
uQBaA85hzk4Z8uyAGbvLQxiGtx+gwksPzK/CHYgx5vS4lOV1bKY07dC3aAz1
alvXAxmmbV6Qmnlu+xx+rIkuVHuaNuNzmVc80QwrOS9b825tf+mHfCQP7na4
QDSQCYejunyr0k1gp3EQK6ExGEB//PpdvhgE4Qab348nQGME2FQNashp3nUe
DZTZccAHU0LHc4sGbdrzNHaSwkIDDJbkEoo/sMG2wQPGayVRJVIQw/w4VZLJ
0ZrIV3tiISXhtTH0uNo/IZPqsS3B0A9bOg9yr8B3FLQbYOg9x9eW7SEdFmfB
uU+A6kSmXlyTmntdwe3iGzJt5+vpIHMBHHzOvbF2D6sUe2IjjMgM4Orv5PlH
OqyP6YJ43A3jKQoMIP3Ld1TobaMKVoAj9dJaUb/lXc7Ov9ElSFZs6f5uHz/W
6FE6pBYyYHOlNgz+NqlfsY0gQoxEEFSvdi9n0FOHWt7wZcQvXvVkbshmCFEU
sEHWGGHJEfoKyp2ey68DSbifY8q+mrGNtMu+kWV91t0DGza7d55j/ZVZVuuX
EpQ39FdZLSMOO2omLDJjhQjNd01G1azuihcGEkMY9ofP9/JGN3qH3OqPB0Ry
Rfr4S6LYkG459gPM5JwDBSWgRNgz1gNW5+1Ol3QU/LMCQy3KZePnic0GtJFM
1D5WdofkEaj3mqczRLiuKaYOhNo9QY1kjVCqBOk4ic30RRjffGvY4+BhBTcG
KMBgkPBvszU+UjYhvCYnJQe/zXwaJPGrjWyE9hdcAC4O8HJtXJeq737EXqdv
H6kbixnL/vP+jai3BoL0dWY8hO1TXnEaS5DWIC50KN9/qt8O0F2ARX2qL91m
0MWV79oyqZSTsSQQ+xRzYIsPzuIMthhmSYOB3OZ6tl3rWgxN7jc+a9ew6xv/
RMOKoYYVlyUoGvLVxPrXZcYW2d5mRS1Sl/G9OF6cMSsVI89ZUpFqSFC+4W32
oZGOA7x9HJtCtFdTiW9V8evVlfM53TMPiCRH8OC8avb8AtKoL+RdL4SXsQP5
wp6AB9N4U5ffDLGGXYrMfdPXqTGoKivKx3QonL0fP8UMWvQTN0xP9CE6A8O9
3JE7EtF14b6Piy0fGe3rL765rf0jePJfmqR2UpMXMhT9Oca+JtnrP9dz2qwn
Ye5x77vVcPYyRzN/kagS+NLjOfQBI6Nj9fLlbnr1vzM6FI5GjjwRObg0aW++
8zDabH+V0WL7cKOKvEYHzdqIPULWZEXZ+joCeLlRBl3thF1DTX4gkbkOaRMP
F0dS3qoXzw75SZQm5D1yJ+vSluiywSJ+SQAf7uiMAh1lBcItqZJHo3B/uK4f
JrEni3C8ikwRS+QHNR1wPnQMFhitBmrVsWJAwmLqU6aqUOhE7ArLVaZBMaqH
otCiTfw2EF6IexYdTraI2RZ4gV2vKyKWzDwvQvBzKtsfoPyCtJGYAnUBbp5Q
WOkkTNopBSsj48A4aEAuUpHpUux678USzlJ4gCbknXX/kB2aBBBHSBXEGTZF
jzzBRF27u5UcljRKo4Rhs14qe14hF+j+QmyQk+uy/sGIzB6GTqqG+ten8abE
vPvlqOy6IYaSmjIy0bu6XAj8lGzyEID716p7pPcQ6rA3ryo3bsUp6viKJLEY
3xmx0cND1LIIT34rDIvZ+E+9IqAYlych9zlhpqjFVTZwGZBX5F1oHPbPOaUx
wLW6PrL0qHYPeLiyuMjobt+zAWkoI+jVEkTOHwVt/MXkuA0Xj4x53uzpdKcb
VOwwlniOyiq0EwJEdCKRuV2Tf4+748z+AmNCK3cNa/ebQvb6TaIia71NJG6f
FxPMUbKcQMB6RsdOyk9Eix8M5V9RaKWg/UGgup/86H7JxkI8lSRVYNIsGAVP
6zl+qbB5HqipNulq+lD5wuL/B11OqkldvI+Cs4yL/9Kx7hjKpo4AGZYVyOmI
Yax5C5Oc6tXUN22sJg9z4ZL2vsj0rP/hLYffj85os4KRQ6j932BJh/OGPrKE
DZR9yJ9PS1EKxbBD2PcUWuc7UGsIf8tfsB8F3ouX9ApEOIm0ZoXpexlQlQnR
znum2u6/ICvHpVpIMerZusUfvjxShQHSGePsnKWnkBXxOmGknWFhQt5ShFbr
kRzx5V963Y2ALhpN32pW3hvaSqDiNzuuH/EXm8D3O380FtHV6tS4bpnOpWuk
NsDqZFaiVH97kEYs7MBrCafImy8iexp5mXDMM78VD45och/bx4s+fQqD7HEV
amrMSEMfIBu123bTAbB6ZzWkMPvEQFQzb9jhaPZrbKuKFqSKSmJ/bg4ALkaO
Lw/27gPxR/6LssqJ9ogFVYPLPnUhId86EtAipGhn0OUJ+a7kMBDyUhHte7eJ
piHSVnE17tEoJsu6ox6bvRs6J4+LW0OhJrvDY+3IiWGV3kR0+mHtNqq1Tmd9
naectA2WVN078dyyUXxIevbRmIXnmksill68oTm8osnj+17BEWqkt0th6d2t
ud7IuCKn7/NwvdsKpPFCSctkr6Ud22b2F4loUmO2ELX5DVDRmTPK31nGiIk+
Pf4wjcsFOV8VJ+9Eps19whCnLXNTq9Kiwn50YpGmFaQYjxN9ek4Z8cUNqkrX
pMMG+HuYEhhDETn5trK5teWHOnOCt77oNEmVdR7VktTlqvN9lUC2PyFjocVE
YSSM0F8gLkyvEkvFI0e6a5IsEQb+kzrYVV7IWMt49oR1wNWXJBF+52H665Z1
7N11CfnsfBS0FvBMw3UcukdaUrTQHolcUGeY5Rg655Hzv18oQFwHhlbvRW8e
qXDfFRcW3XYpuPyWRMpi2Hx55lysevi/ccf/0NOZLefAqRbA7KnCBH9QijXc
O8WqJ6pKSwEtF8FWX6odXB/0iOLH+2J/Xn5aCYhtisi0Xz+IoGnvkBcBGrw3
7I9FCDCxSzoES+DS4AiOLGgmxUNXMVOcNTHH0jOyvWa/A/lBkG3v1l7fE1xu
nE9T6A9ErzFVlcn5kue4uv82/OdpdrO17toGHJ2yK2pJxHjouXWFKDKfehu5
l0RuCNLJxYpv3Xwr/Dy8p6CWS+p+U0rk3zKuzzf/r0fISZj+DjHPs2xAV5/n
H/ZRrBF30WVANVR71Lz268g+wz+dW8EiFBpZujfXInnyYwlNZnRWBWtJaHA5
Qzpbo4DusdlYreYEM90DdL0lpOggfiy/yC881yGJkz20QsqezemYHZzBxFxD
7o3CshTEj5IU+A6/MK/Bcyr0m8tId0kC5/3DnduEN3wHmHMExgjUJqD12Pbr
ShUp+Bk2OdmgffklE1t8TBi7C72Uw8xTaSW94QKu5hCwW317UtomocWNFPrX
Us3Ev8WmoJ7TAn6HRAwk/GmDvq/XosiKSRLAKMqZMBZ2QDa7nc2K8dujYnEI
mh/viBLMFgp/NP6ra14UE24bSGlq+DTuSa09qRs2xRAFsFWqHTeQtVAdZ3RI
jywQmTQr/wi5klU4KFzXZUB1Qe8FuFG6Xtw1mmUbf7Y5cpsUdjb4EKNGUSUl
HbkUPzenNkQfhcAM6SFEmvDRSGl8AF+5TAklbKLZ5VcsP0IvWIK46MCxM1fs
cgGpNjhDoJXOfDaAkqI123qPB6jpnULPQMJgY0szqlYqGdHtaSYzWwXXXKh7
pMUuYVb0lrHAPFwvcybzADednQz6ap/dBQikxA/aVxoTTVE7A5cQpcJLrVdI
xgXssEeK+ZtT2QOGazMCYOuMQ62WIDLcKFl5H+DTJGegL5O+8+G3HFTcz3X6
XB49XeZGi01JN31ECIOW/JFMn2PFQBgIS1ofF6TBzEr/Gze6nevCmFdXUUIN
z2syCXfhjqEa0dhGIkbT6BVmLpSdnO/owgYXs0iPpkfIuGr2j+k7I+x9f/vA
FyXopGrRgaV7cDleSR/rZqLUveDZBiZ3Y3T9169TWnicnxJRZant6HijrIo/
cULzu+XMCxMZBnh17wzit21Ziwx+vAUHHxrjSk+RnZm/z+RCxaYwCVdgxtMB
KPyPo30BxiHCz4Dd6RpOy+ab/ik4L0vP++4wppYfLegIX47kuMPzdLEyLAN9
uCpjT44yvZ64MVjhHe0zACKzOpBXLXnyu6kzm0Y44RbZ59FfwWbEhumeJdyd
6C7vOwz7C+moGVInmrbJXsxuJX4sh1KIUyul4mCQ6qn6VErglAnM/66bPw+x
5Le7BBFb+8Mcvv1YjSXmNXkyIKz0IZKwPT8yWjcuxQbb80rH6TEZBrk8Ggkb
xSGrdjX+KKV0/0LIk3ch8shEN5vpnhrUvcFI2Ko4M/sZFwq7ypTd5DyuBIJ0
2aibMUvKijS2YkL8nSoq2ouGm/nB8Xv1nT37ReZD0DlR3ZJs8uH+CLzfYK1a
hTDAm4lZIXRtvc7cy5j76XH2x8+O5d8KXmdZ1ZzPveryiYiWeJIneEmLN41j
NO3G6MM6ObEBkSyAbY8REM2xHPDSQiMs3E90o1UlGd5bhxbaIcj95Edebh+Z
gANPRFDRsu3rfOfzASILNhUxeYPi5CxRrbhWS3OXi0BGVc8FTluLQ+AOblMH
3wWhjvA/nHASPY1AsqoU7AMqN8H10HWFtZjY1iFPum6jeXheZ8UfC2bnbQk9
HcnUOxIMmhWA9V3Gtl5Cja8UPt2sLHOcoVyIDcP97ZjHYkqOksPVhqQpAA0q
bflySSf92g3afDbJY0W2VmRRVtwaJenBPORJoCIUaaYWUabLIwN7t4ejkBE/
OTge6hw999gsbe4+6Bh1NQ9e9fbFLNQ6hzQbp2t8ImJoqhl7otLfSbjK7nSX
eyjAf6csXn9XIBDsqafLX54gi1HwifxSH8BeOsuVIzAexDnOOV4Rg642/HFs
lARZ+rRVV5Z2fqCcQ7ZA1aa1UqRaKLF1GbQ0dFcgv5BXgNHLaJV5nrnd3Lhd
6vqMyqcGe5CF9i/ko9e+4oahxadd/RTZJ7kG9nNB0hn2zqs1f/aTzXpm8bqF
zpAqwVqhVhoMzewPF+BBVw1w8G+yeHkrBcFT8fz6DrVN9XKBetNlCFVYo9gZ
0ERL4DzDf8pDZM6GjTE4cfhNYjT3YBAcdZpE9yO2mPWHNibOKRBJ/Wg7EH6+
b8yAm2Ah2zQKlAKRIAaHGRn9vTEPX1+GzQHobOm3TgdKV2X6R0MY8tNKrRr4
yOYcSHR4zMyfV2GealzNgmfRj3qpoPUX6cNmNu5AmGYLvQEI6qvSlzQKxOBT
qsqHn3rsEzBWfssOp6GWGZFpgu7GK7tQMErGsRMFMiJuy9Qu2gmPT0DhePU9
T+Jn9rV0PAJD1k9ymiTZnqT+TsI2DvUscJBcWRxtFLVqZHu6zHNLvowh6fdA
F9FbWXesEk2Sv3Ms0JWJn+V+PeAQRZkChtOu3AXzqM0kheTsVYj4/+rP/yZU
3lDGHwGauRu378pt/oCHRmI+na4ZmmA+vukTTOl0tdjGHmw/Yi/lCzkXFkio
Q9K4UUvyjovJgqBFG+NP7pwbJjKQ5Ag+rYUMHTkCSbxvhYX6vGH1iM3eEc39
xSm8rwnfwHfLFgIT2dMKz6NRmD3C3GzMrNtrv/S6Jkbv6sFr3azCdpOt4SMU
oxWA7ucOe5B2nC636ffTFsYJI2CHa1uaAe41pd76XY9e5OW+3X3bcg7ejmX7
CVfurgCWSnbDQ2cSHbTlDDqTCNViRdBPp7/Z93V7ziaf45nVq3fIJUl76kK4
BOeLkBMGMIGgPDWvGs9gCYH4BtccngLfEpnhTPvx4ZL+fzCxkBG6CfnJIGUS
w5ziU6yeKJS4EmeXAhwBHdA9VGt4jpLeu3dFfwTVMshZ9er+AqC33esC7eXd
ho8v/A81TT3tijrwTESrlrVOrl6JvpbsUPNnC3uc7u7ME7iHDRFIjLrgD+9S
QqjLV/NiI4oWe747dWcN06g73G/xsVlOuORimj+WDrkkSI0vxMovn1M50UW+
UJfk19qVRHcggM1bdgkVsP6SSJnlohUzQ60r6gH6+2ZZCtyO1oWBiyS/6aeb
cirUzsjLvFL9D/h5drT/lfV/Q/EGA0IajJo7Roc8lNeXfFWEDHfYuDSklGnx
nkD55lCCsC1ROr/JAsonSBU/+Kv2ugXR8+zA1rmnZkqutDWaB75/cfsAbHYX
ttdnYA2H6dC5R7HBIqlQhWV3z/1CVU4otVez9pIHKIrU7i++Ym1SmhNita+L
mWkzvoZKxfISzmiFv2KtFNNiajRdPTVs/NIToHJcb6ptksQlmixVrqDmI+ez
YfwBJtPZpviso/Qf5M15aNFMYm1sGELeA1h2c5qfbsod/6aOatrW21s14ed2
WbGjO7R4Eqn8dHQ4etW+m1gYitgxVZgFm/0l3KOS9yCi0gwD8Er6HkjBSoLq
Jco1GabWx6kK7GXiK/YPUz7sSAjNKy9ZGHco6xUPNyX7XE1CEtQpbgM4D3g8
SieBHDkKS3SaahBIQK9VnWY0CywiZY/L+JG44M2ajIgo2v2rUJy6oGqLdkd4
zmEDU6TN9x6JO88kF5AMK+pE8OxbpcdB9uhYB0bDAoxipgviNDF6f30nRucW
DZGfwxGsLG1k0YqXLmUwwAMhXKR/wAQ2r7c9GF0iLABjTO+7r3B5sD151RVF
zshlRzg4K1NMsQ6Dgbtk3NOj1lyx45UC6BBQlE0gL0oWHvTcvEqM2pka2uzd
mI4QESlrSc92RwcuVwrk/1q9vM7wVPkBAi+SvHG/E6hzWJzQ4Vtep8zPIE0B
Vh0+SgATRC+6C2raGDFg5X14klpfwQ4jUyLNPQSHcUifczEXZfdjFD1hQ4as
hmP0M6oI/uxTLBoBwhRBTwHoApxLauQAovQJG9NMXCM+kiap6YgTDiIWwFws
G8+l1cCs8lz216iMhawccRlDaOn9rZAPdVnIVdF1YR/pECUnNTF6p4jrULwd
Hk/xW9cfeidnGlI6hRE4BbCJx7xUEXJe7CoHJ82QQu/l3PzCZxpavSn1vIEf
ZgX6gz0F1c2EEmArd5jTx+/fa9NjNa7tdTZNvwzOVubwyPPzBtEOkt/Ta1V3
9T/eWC/o8N292VlLatlVgDSkVzJ1PToyDakctouAnX0Gvb/AFsJRPxkTkBO/
1RgzkTF0qYduQFqzipRFO3hU0uswLpSQuxddmJEFQW3dDPqxnId9fPrZ9z4W
i2IXi45T9NXY6s/NM7Dp5kTzTlHBKtKtZFJTOSK6aZ6m+q04HH+Kkghl6O3d
zymJ+OJO6334Z+2l/uJEPFBmCG5TTx61f3pBWKV2GKLoD+S1QjyDTCWqfau7
M0HtUrMvBxB3K650BN9HXLUidDGIabM2a4DgI4GHtGouoSWUulvHngjiENv+
3fG0GWHHLjJ46oykw6+Whm/otbHgdyFhf/PkB1p2424/jX8J1UgDcRzvB1Bs
LWV7NBV07vQZa1hSUL5zsjfK+MyYilCRuiv75yKu7lEsKssK7wc/44iI6bM8
bG84LtN8BXRUDnoU0qfQm8JNTQzc562o0Ss990fJVppo8mczcOTKYLA1HVIb
n3Jwl/6koeA9wpBMhEQXBTDcV/FAdzs0GeRjqjZ7eC2Dg9l1d7EnWyIsfvhM
hfW4Y74E2UdllEsavb4PAZf35DNWIzGHeTDmuneNQPbZf10sUFJ+RXenLqoF
5HS1YyLQX2GDx6fuGQ4AG4QepN8aAF6tjzJb/X6oQfUIdGJXdMZKmZWUc1Q+
6jQHVPMlM/kNpZYuaZoC6OFn0gM2awTSbceZDLF4EgaozieI2pufm4taILKB
/KGiWuoUxb5W8h6EZ60DadsoFkqtyhOGoAerOSz+tFWM2PBD83F8iiyhGj/o
SOQ2yK3CR4l/mUZYDwwezbd3MDmcwgXBvB5Jf7f2BAvlHnbF+Mw8ZUXGw7EP
hWoVCshS4M8xeWE+Lm7A/8lSuR2681oXGsgQ+Xucmhw6UqyvrXRQsqfij5xT
7fmg2fhDGZlj9yNtfRxsXHGdySx6/jO+6Ey5SM3N5F118vaffomSnMafDrSw
5yfJi/PlOFkVvpkaK9d/73EWqFHQWnknH4C79iUzmREZ2B112zbYq6tzlu1A
US+857sZ/uNXli68j6Bo+guIgyRsIyE+Y6fME01fpqcxvmaXR3FriIp+Rd4H
LJhuA91Rto7/IBr6kMTX2gPtoc4KNZ9wi5EJH+3Yz8EvS9GDKQ9Vbt6po5s4
oebl/WZE5rDh+0rdgC9R6+pjeX4VuP6vfZu8mUHvp2pOKHH7DUCbBD/WIfRJ
xfpCqTIIYvtRTgB6PNmJJZnkHuuq/8axO18fFQSAcEwKiW9ZR7/GDQ61fYCU
CxlNzLWpFrPG9M0fFUb7dWjqYsiZyjoLcSbunBl5bk3QOXQR19VtL75oh3bX
RaXgbTAV4TSbpmSfl5qk0Hv61wZvI5CGMPyrebX9/p4AzqLmMJrW7UVrSXUr
4aFZtYYfohtVdaBQU7kdOdaHWxWuf7nuI2g9ssxKpP4BjLeyg9ldszQDhsbJ
+fYgu8kzahNVM1rlthIKEAPjHrqrhraRGfmTp17KaQYExKO4mb/4RqJWF/6p
vu2CPxdQfHORfu2wbNVeTcvXgkRs3ugrNaY9VfvjtEYCVUzrGErMwIphtr34
IPlCH7WeecOLLHmTDYHxGEau5wQy3Uc3dMnWvo0//xIXWZB2gSt3Fdo5lxZA
WoX5+rmoVxM9kP2W/5xD0rQs5JixWWvZDhlZGuxkaahtqcyBB6FYEf429YBW
28tsGQKeA3SdPygR05d8UgzARDO93bhXV5eCoP43312PY7NF+UN9wpaFwJdv
D6v6j2+ttDTs7IyLan4x+orqbGied9/NUfz5XizysyCAFYj/BRDSjPWdSjJl
MCd/CSnAj/ZwosQXcWcUARXVHlgS8ocEjNLmkyDNsJufvI+FIVXM3+HkIm/U
xojtPS1b//h3IPe/woalHtY7toe3FT0h7+fGyCxbhmi+V0QGi+9TniQ8A3Vj
zXjPEODimL56XBV915eF4Iq40ee/kF10xOPUv7lRu82RV190zE3DnrSBYcsy
4xJ5FPJL+b5fT+NCkm8Aw7/yRjR5TReuTBV3w2tYvFBxKMhBxFFN+1Gs9M4r
t7ZD4Xze/8n/HncO7DkFQmAGkoGmUcYYgpca1A3qSmwRTlI1WKj7xzSHsji6
MAqaQ277lZJRuB0dsnUxUioN+YlImnqjqXFHz95OKsWInL1lzh65hSTL2wMO
CZSoMSZrfl9zrME1tuiePoPz4RZulfqjmYUdxgKKn9HT+TsOepHifP14BqoX
9DnPT1JhDIkATuC1jznRMXpNEwjkkRag6fUZoUn6e57vWfb2Id2C5ixUZWmE
/uKL+Zz15dboQyvU8dzASKyR1x6SERC/MctSYy1cTh9bemJeSzUs0z/84N3M
k3vrSo6LCJChiK32Av0Af0gm+fH2AlYt9aPz+i8aVRPlcslxwZD1tmqvkHNo
v4OvEuY4496DXXkw+fqN+gj4suiTQb8vBMdQW4oAGGkEY7M7cs8/qoX89KWX
2ZW7VIvNMvSV9p68kXWqHX51Bq03Hkfp+kw8LS28x5ZTh9sB3Zu3at8eqxmd
D5beB1P4dMueOc8zQnF08IbHVLg6DYgyQz6JTL7G+pG0QYdDAzuzopHLvXpm
uz3keYlr5LPiLn9XoYEkQkdH7ehoHXGaKZYhoIBVRX6c1Pe+KKYR7IfezMOO
nH8TT9r6gNWpZPAtVNXSmdGcmxaEHFdjegiAHZKjbA3hE1pdKjn1xafl2mZz
La0fmcyKs7+h5V6U5YwsF954Winb9SiVhxhhYMT7QlLWVFVcsKrbkHPhAjtJ
tFjWGf6GbDwon0uxdO9H/hmbUeYEXAhKba3zK38CyrzqvGJ8u2R3scZdPlpa
AQe9V4w1cGdWhQL9LG/+NoXf/fgdTorY+Qhq1TNFdu08m1UICChmRkdJuzsU
d4MDXUzBPPzkCuDBcAppUsGHfx9AgbwgCEwFf/FlMVgoQ3slo8HxP1uBPBSK
j5hr0TVDwfiSmbP91sIslbnMD7H0BnA8OGefsEGIRn3qQG3QNJGl6rFbvufD
822qXjTEZ4csrlrB2tgPPD2zp5zVaLHVXk7iIbmWmP+1FV0hLBdlrYfzLkBF
GWnxYlYHfYsJwWBsv61EFTIbKsWfALravjTctJDl5AP3n9dZ9Z2fvDsr7mWh
BDVNQiimFni9o/oNDvIK4rgTyBBcUhpZFpyOpo3DU6RPMuPRfCGrnuc+4rjo
nQkQArDZpRlEaG2utaZvv4lGY3aZG+nn5V5qN+eSst2IGib9olKIOvNZf0Mr
DKz1jutFbpiqcxvcYPbKDZ0OlASQIwdPeHTVKHEUYVtCJCkhnY31c3nQA3CA
bGJxgpjhQ5q8swAoh4+9Kcy8wU9HaVcgD0+iDZ8j/Hkjg20ECFRger9HY0pe
Sqme9NpX0V/9uWVST2KXoX5RutGSSiIrG/v7JU5W/z19mQc6rj93vO11xQvw
w7gGp4qDELhFwyyJGOxVpHOtz6TikmrSkgCcu9FfzdPGbP430EgyRDizjMNX
qWx5IkUw58kPpi/0KKe6+/BB8Yd4W+jlFn32agM7fE9k7UnLQW9K8cKX0vAB
NSPaYr5+ADy5y6V9CQf7QiQKClR9bAkpvUPKd7dDx6XT9nAr/MFoBiQP0Xgi
zliuq24pZDaxZnA7rj0naBfLYLuzzgmvxgq+c8PkO7ErByLEq+xf8mZnWnGk
+rO6OZfzNRnd9wgoVC+ZCM7eK05aATq/esQx6u3gqudxQStih5ZwdIxPs4Td
H/DZaDgm+ksoQDFvAIqoBIO8pn7iUIFvaoYOR57tb8y9Yt2podeMJ96cQRrp
bgT6RYNPdtRHZVAU4yRiQEhh5k19n0a+MjsP69i++2InuXINVAOslrDB0AqQ
iCSiES4Tz7N34xtA1aG6Rf9/8Zrth9JwvdHalXXipoc0YnQQqL+cXZ/tfAbF
2zxtZlJEre0Y4ULRFk78bbFw/J8gsHlTx1hRG0Nti0GNKm4wW8bgiSWITbct
7Ssgida1ZJ9jn6lj1kECdICrpg7JMh98fmEy9uF3NgxeU3sEDS+Wq/9zA+u9
hO4DCj7GFyLUOdDcwT4Y5e8OaWQADpUw8BMrRu/DOKS8H5zSE24y2B8ODuFr
gxqZ4SYmh3C1jioMgSrom6iPRNOonJS+KGclI7YNh4+wYEcCwUTWECSf1By0
G9UEO3a0dYsRVR8gNUtiMuIi7m1A86Oe06RXkU9/yTKVUiJ2w0NPUp8WbAMs
Qr5tMmpD1btpZyyjdn4FoUHrrI3t3Kcy62FDZK6JR91wC51MuzM6EknJ4JSA
4eclVHj5xCPgMPmEEZoOnRF5BsKtf0p1MurqqpTL/tJy1OwW/j5Vhvz+1Eas
++ILxIr3kqwHWfAxerRT7GYO56lniEp4buoVWEhRjrV9hA5MdiibfvNDakZT
j7n4DvrudSweLMf7N4WVZ0sH/XU17M0SXrCWLJctoi3KAZ1V16MrYEevcfQU
W/xxYmerx5Kx88iOPQJjTd/ZCzNKOq60hpUhF0R8gVQckCzc2UlzsTBqjZ5Q
bhHy+JayGuVMKGZIXMWtJEwxjOxLuorkrsndGfXF5Omit3K7Rr1GF7BLJPQc
BV7vFf+LQDCuXTdb3emfvHoJmsgVmj1O+tBryM53Bhtjpat0nY/USFYPgZam
V94dC3vylCJ2SAPrYN0yADwGJhpStuyi3hLvmWVmxOTuO7M8BMQfsj+Yky6e
taFvmHptbBoLsAyEWsGbkvNkl1GbDcco7vQw2bmcbl3hN6V58DlI3RtXnWjg
h3lxQGOBeiJvdFjeSmSx0gjdo0VFSj/iJwgTGmWgsCpB6nfg33WkzrqHR4ax
Y98q63p5BvsZdUGXVgq4Ow6KZ7WsuwOluYtlpLzpDDsjOXasdLMAKA/VYXp4
+XZfKS/Bp7NvAr6jNDIk53jT6/wJNucfJ/gg0HKRjO0WhXQySrceFYV6pKGS
3xcvrZNea2f+tjnAcY7ehylpe9UyY75WrlJCZvjRONTL6HuLwL9ouj7xSJGr
npqkXjOEazPLyBLrjyZmfwnTVknE/kFNTtXm9H0pUKj9GI78nvuJ7F9LJOdY
dnaVnwbYdNNtx9DO8plyLct7m3G4IXDQs1FSz8FR8FkuFE45uMUAULdCUyMh
2WwVANeu6ZghVBOytWe4lF4DZpY7cHYRexhdnQbrPUgxnNutrXBmlD3NWZlh
UFfxkCzJFLQM/1l+t9o9Ee9CWJnlxGfNk525pVRdhXIVD9E7PWaoHq2Vg6JK
LRqM2ifE5OY81J48MIIVstANv9EVKy5NEMuUfcInEzmpxilSegEazQr16xKW
4R2HwUAKylR/3bJxh7O8rR3lq/FfgqPCCN9XwWYanNle1JxKiAqG+jlkR1ug
sNazolTR3m0znhJXuP+EFrPN3S/qx8H1BinBvrrWYBITBmVS52PIMSQy5rHo
bcLEEr0vDRLM69gEDQ7eBTEVvagsGbCSK5IvCBIcy/sStrdwahnz7xdD3jod
EJhcc3oZliBHHuTpejyxodBAxSqZ2asRJdZKLG5g/5/Gfl54Z85fi4aq8xcB
t+BacwjobOAegu7296fx6Z6KCioKAa8NGm+GylRXfzf7K5cs0kxSnyBBPDFP
n+JXb8GQENhoVxfiYT2BbuG+2V1rCZpUxwxxwvZjsrRAA4BXzbSeCNO7MiH6
6V+PrmadzC4wjKI78CrMKvrommJmoHH5XJulWKtMfw5Y1fmK0xNv7yF7qPCY
AGdtQuvGfgik3JY2zK74EL6HWZVL7dqiQwJAimGquhAlW+XOn92+9jUZvCsC
juZYARfuy0KOLTYc5sTCf6TD3pftLHmios2thVq9XltZjF6U85i+CbzSN9G0
C/91vuK+3NWgy/+/aazhdZACJOawJTr0T9phN1myIwl8xvRpPgvvV3VIKEl+
m4d3yv92gFvETukI67jCyFSqfqMcPT0vjermAlsahlwN3ww34Ec5Jj6+xa5k
Qu47oouKGVJHKl7gkh9MwNAeH6MIOlZhKpuyJISDJeOdNeSotzzzxOl+8JoK
DeRTk+FeivkWaZADUgZLMMlf/3ay4hvNVES/BNYBuSq39IowpdrFdsfN9OqA
ydvZWDX0GxCV0A2RSA27o1OlC+NB7BeLn7PXqcbezVQ6f/UTn13p3Bi72ZQP
VXTwGJJbkL5xpGs4d3W+9yFG5v7Ii2pTLgHr6h85Qu8y8r1BKORrQ2SgxdwM
QrowYP9tTLH1/3uQ+NsgS102XpZSdUcHB/wmosEOoQ4ORf1Kl4HI61fHhj04
zqmSZQv5ce3XXdoJdU78mCXCp3Fae+EqE7/DfpWBWZlZzCrTvDyQ68LouJa2
Rm6iCrvyPnoEMRr2sJoKYIJdcC2Idm78tUrE4Uyd135ppR7jaOfhlbdlOn+W
MYBMmXypSXW9JSrV0vnANuzOXvw2fZcmMiGTWdPaT+1kg4Z/Q8A4LOo1NFGr
kD4UsItDS63zzKqRj2dMUjeJ3UOdZ+cyHurIoYl7eYaQ9fkqdPNb4ozujO/0
+/RudpMJuH1ElE2v0wDxKtt9FC4eBhfzmvH7QSVnCbvt650BoaeKqffvGFPs
vL0IdgCxqwP2qzpG64c+LwLDDRaMVF6H4KyNEFMRE4Poz5WK+DhBYJ2mc+Hb
6TNrr113ycbjNWyCljFdIH5q4lyk6Df4suHy92Zba1hojWrX8VI1KUTBO+Lp
UVLwjtJsqZsnteDUle/CdvtlfFaemBklLlbPh4MU9OImns+v2fiHbpG0HDy/
QEfZDEvjK63pw7I4MqnsO+VckKd6TueD6JHu8Y3ovpIwi28aYu6xMYTv4BS6
P/F49rMIACxketxJYkuMOFkAoNDZgzOzyQt3+MsQnQ8QDWTPwPlMRj8/HG+O
A/R55I9bKCu7Ruf8iq2fiIhtpSXZozQzhauwOviNZascrP9Tu/yNVF0t0LoJ
la4jVv/5+VEjPg/+BYOn9FYf+2nc9uTdavv2uuMASh6KnHQiJfSWK5SLd9NA
tzSxsybqaWgQ0oTpPJY1WU+KXuje8lSLi5uQ5F00jUHVXGAih145Ok6Mmkvs
kKTmCU7dfsO3Zt2C2bmm9JBzcviWioZcNBpWsNpaaZ3ZnS6m1zb7NCM9Y1AG
2QbnqXHRM/njrc+s52TtwmDjoQdzLhATs8VYD08mKxPeCBNOYkNNvx+1xQYJ
8GTpOowYDaR3iPe7fLyJ1dybY5m5vPXRAmyxwoe0XenuixcNGHAY8lryYHEQ
eCKTXQXtCgWlL0oIMCEWcbhsgMjN7SvyrAvIhLuwk2kv0BLIDC+lSrm0PtkC
fetv133Y7cQhypqQ2+uBexamE7DS9Rh3EuEiFGtfeQPUTlaPA9i928UHA6S3
Y0fx0mjH/5smCUmHEqsi4cWxROjEa0BZESkF3DLI1yLDReMMT+DdzMG+zSqy
YC2oTEEeltK09shHJgIEWtkmGGA3TCXnq1yof0zGiI2seyMQ5VQ3mNV86Lvg
6s0VLDFV3JX8RYpCz4KPnNhRHxX8xUj7pM28HSQDEjRx+Ia0obRFkk/+wXuM
NEkfcKP9iPAMY37dCmk8h5gpBdbsqtsjRTDtdkMmsGaRVIzwGuMpIVDweEDl
TiCHUOKT9yBtT/qt2JgVHsDKG/nKOKr26P/JyaWxLnDP2lz7dGSssnEZ45Fe
r880onmsr52h84bvNy3DVn18sPbp1GeSs97v23OhWeIfNGsRd4yUFi+mA1yy
pyzPIZana7P+SYh3gHWh+oW73NHXm3sCBJyFvgYUgezVqPYR3OkeavQD+ojN
3dxQhMpgg/Nz8odhW27VX/LQg1eaMbcio4ZxRNmROR17Q1IeXayYw8MgYKdZ
iSjq5IDUiZQGLZiKg69VRAr36RUMuvkEdeKmmKGVvkU5r0STVIfrIShTXvo4
/sGv+64s7LPOzF1SrsRcO++sd0CzdF8A4hVwdlXpZksFP+c/7t37jRwPgGZK
jAJHhgCk4IfGldRNCclpUAfnlB0Yw0syxRdWh1zU7tcYzj17M9/mF66d7NYV
DmVSU0U29L+SsVWFZiYoWQX4m1xgHzymrFLJxgjanhXouqecv3jZtNYQfJSf
E30kbeyia/k2vHw0sXWSMKVF2fi3Qp3T/En+SzuVdW7fB0PvYgSVhXntfrzO
LXHHJMZFX49Sgi0Bc5T+eQ4xjp3ZY86SYcWGokfpWCWZBkqGYX3fAPp94UIm
p7Gi7tJxtf4ylDWcJBIFrxV5ewmd+RHZTRpsFqJeFbn8eqyGNjRx6O/lpQoA
nv4NINatWxST6I6Bp1OYL8JDnK3LpQ6nR8fY3kk/B6edwFmuCH5QxIB8Ne5o
nzrbmlsgeSazrUN7CRmYgjAVkNQEXIvMmtHqr0VFGKB+BnKMQ85o6tnC+KEV
Rrn2X/tejgxQeU6nXYE8WdGFJd1JdfIDs9VA90VrDIPKaJlPPLxCEMMupp29
5ENz5PFp59Nfx1tlK242UJY5n3NtLlDddAPt49T5sjU+wf1VVQvICCq592Lp
VN42hs4L3hr/vEKM+HkGQesFujViRCnOxBO9P4YP1Ny+DasE9d4oxnIg9nXL
5OYMQy+LHiil8jk7mtELwYDA0iV1f7a/5SxsMm48o1r8yKaWwg7K3K/QcobK
hqGKkLnUzsnvgFVgXmaqTkxXG32ZUrCnm08lBL5tMTGiOPBHMXVHw/pbmcWA
UTpiPfwJ+PQGeafcFr0LDXU4wxxbyfw+cCORtiyUHS3VeEd9Y5rFu9ZTdrVK
mpcTAOaLleolROd04AoE5TRz9yA8HR84IPd5tbeE0qS7D9zzTs5tE9M0IRut
RTk+fUVOEUZW/b1Ki8KbJ/liJI6fBz0R/xSaLsUT9jdWlMjOpEe3I31ZjYPO
0scUt3+pRrUPCVAxeFFl6OknYjj0lwiQSg0HODwUXXSboocF+H1emIzyrDTv
+lHdt4uqDHIHhI5fBbt/VP8wOX8uIPHs43jiF5ceXGr7KZWkaRTf4v8MN2YG
L+Vq1lKaTvkvLXPKh0jX2BCqtrWmh5U2oadpzHcjmw/ekGpJxu/5UnrlQOuA
cYJ9S/jA5F/BPAZKfbt+Px9eJroyMb7c/wDOyjW7vDIyKEFlR4mEhb4rY4xO
OOhI64AM8Y5TPAGp8ZBez433BlxoGMNoke3jaNHKz7CwtpZYcLBcI5Hz2NTX
3anD2tK+ufDVOEIfDWlR9376GXE4Xym9TlWRYBcywAv1YSU2K4RkSdLlD/KO
BQzVrAzJeTi9mvfO6ONqJNy5zHeHfNDHoYTLFbw1s2RrtnEPswiZT93HiwRD
NdbLtOUUNrlkE0JqBVvbbOucxFG1Xr41t3I2OFW+YcV9le2uO7d8CBwOKtjn
8/zaPHAcgIBLWpVNpoltJ/E6lkx4gDixVXr34yw/xW0yNQE8rUD/GaHPrOjo
tyj/pqCmxmVfQ9A22fGy390R8vfOwG1NzC/x4pS60+R5Y0HAyLPAnNO5Jht+
Vw6I6VNI5ta1Pd8IRuUgdRSdoagS8peFx3dyO4/KSenSIepVaU9LCNoT/zxM
nPvhkdB+K5zerU6pZsf8MDYwaFTwNA+nHZTS0Zo0okG254BBO/3u5kirtQ4O
je9NquuecegEGhND3bY64iyjDCdhBPKYzbv0KbxJsiSI6NWTDnl84TYMnHk4
GDO5KzO7PxAJS9WphvgV0l0goHEivFEF30B3WpWSXI32edml+mflLz0ijxrW
mIZJyZ5zLWESkoK1RiciXWpugaCHUclKB4u0q+L65+WDzSuZ6yTO4G+dRc/4
kosKDc/9zL92/emPM4ZhfNxvBXpadjiYCLlzBQ2SCCy4bvVAVeNRMk5i92TO
KohnTm7DxXdJu39A2DjLzoljCfxFHOxmnFc2VA+R8VA7OmSoCofph/6FfjaI
YaR2nzVsslTS2/D3XQ+SYHbc/bLOl1Oz1f5m2OaVqtrVoi5RzpgiDiUgJbS3
2UAIV+oFOiZzA6oV+FB83Jj33N01rfaySpDL5t24dcxS2tsuMd7d6gteigSF
4uyXzN3oFCyquy5uwDgtEC2Xcqe/e3D3P0Wa/tTBXYHZMEeJr4KSMQXDUdHs
Hdx07qLALWtN+usdPU96HeiDQtmEYhxNMs88mrw7ZLEjW1QBy41A9bWFPXsX
vPeY8Zl3v2V50uPr0vTbAXVIA7Z9A1pE5I6Ofo6ji3z2dzl1N9yXu7ZJNxVL
mXGPCvpxUl882/o+JJ8KQevlEkugwX+b4ayJybAflpEENoMigIT5mdv8Gbpk
adw8wH6N7s5y987cGKQkhFk2uxXhfvlJA1YTdNjPqp9GD/voSh+SAPc6aHZA
wRy4DNrYVhLLuF7aCmHQXLh01DSOFyNFtVjrhNZqyterUUjTSMdvfq1j7S+y
qt8h1UFA/RN1TdwYzy3wpZVVHSSjFRUOwGIxAQwF+iOtUEu8nE3SgWwCrS1Y
ecKwep2pkMTvCWeOkQeTiVvxLMRmCVA5Ic0yyOoRbFco+x0e3+AIyJLDuvx8
555GJ830udjblcmgHuva4L5qOL4ylY09XF0Nd9f9+4dKGdF1Zm3rAE4I5+Z5
N5fB8FSQ8flAvsZNLTNlp9Nd25C8nEwnk3C/QROCynj09QFc62o4BV25Bz0L
QF0xP9QlRBryRixhId/Qa+gILNsrSjZevaGzaagt953BfWH5XM/1FBe5iez0
p219FqLJRE+s12aenZWLLdEEXPEgebRT3mbdIWzBfMpqO1IlAUJZWrKJonqN
1uBS4VOBEJ6E+WNIv6e3TiMBq2SIgHIRHCuW7qz+5L83sgYgGDK1I46Ea1Bp
QeubUa5cmiMSGBs1JkXrs4JvIH4Gea5p+k8NqX6VgE+NT2MX/x7nZpHpy9AQ
++AjoDFvQaJVzbwtm5/t14OyvqCB6S/NPQ9do3bO9ubCTebUBIMS49xlLWYR
pJqnapxVX4GSS8xKl4TeNiDFoINReqStYXYcKrFNONy9J/uvbQhFCJE4z1eG
LXuCL8jCzm5ynl2B0LMD9EOn9fUDaiFTiVdBSt01zamOYOcvovRQBXFSNvW3
8a9frlhKvZrx2YneEvW/GG4ToJy+xfu4nkPZSLux2AYNpXPMGVbp6lmBbUcm
eAcWJBeABtjWzzeCMK1WuSDB5K0f5l6YvIRANAr9XrnuhnFXtUq5DUss/46s
ZDqoe2BljE3ts2XhQrJsC4SKKYFnfo1zMBOwA0lXu4Tc5G+EfSssFLo0JduO
8vWUGCnpBMCQV/9Eg+ryegpn3yfWKHPnD3PHr1bBXydJhU45cJDYjIvYeRl1
JN/4gA6jVqXwvBElcr4s6f4+RB4SM8aEVxXZUyVLjrz49xbkTKzof9RXgi2l
ALFuJw+M5cf+6HKpZZSEJ/Ot9ZUgrpaUyK+tqXXHG5dfx5ckArTUkmd0ej/M
yEoI+n/PE0gsPg6Ng4DnMqIWhO8C09cgtvln8eRmcAJ/pTOb/rimQb3TX1/z
0WRf2fuEtTKLUxnzMPBDSvPx3BIF4GeybJ3oag0u6gY/eX0vhHZtkEN2Naww
x3aadIH1p7nN1adQJMljxlLHO5E+VGg+MH9gzuazmarPjEpRpz1RSerhSCAt
YGo4STZHFiqSwyQhdaR6hop4IRO1e5GzQzaziclmRFFx6fKUeipieDF3DbSD
g63/ZAnXKjYduNH1VIjD385B3cl5Q6N0aNZC6iPqDNMlPenQxqgaC/PoMviT
r3faju/dznV39CJug5BNd5wSUh+ThhKOj7PWN9Ecf34vsQW9IlQhYrEylmDq
ESQqDe6bYco2P/Wgi/C4loWBPmfDtOPRMpoaHiP1yJ5zbUDZNWSmba37DuDA
cLc4flAlcZPnJcPTnMTHfWBLSiAkfn4NLKbDxLZsl1XfZfOYPn6/Hi7IodAx
0dqLx946y+HwzH3r2fs9mM1S+lx2k54cbq0xTdz/mT6zLdw1CACRRZRdA17t
40LyeWO35gIXT8nyqjDFGc4e4kHz2Ni6f8KMTatMkdF1uFfJxAU5LSxAOSaC
bhaVujxwAsYyy9E8Zzg+XOZ0YjZiArH97duZpm+D/gU70qozburEe6BxxtKa
fV+7mQcRtwynbjztC1jv8pTOfNWA+HXQGt2LYwMuhgc1k39aTIG38FWnoMo5
ThVjdpi6uarTX+mfNYJ4MvIecWRiB9rneCOza3HLwF/fFGyU4SRZdUYPo+/T
5brVXFBmkNbPCuv6/HU78xM7nDBWU1KjMo27FZ7uzUUnf0Sj9EU2P4fEromw
ENoEbfKMU7jWI3mxX9Ttc5yMMe55amLGGkL53xUTMg0TtINbp/u2fuYigfR/
ZpEIpR/Fi/QbrF217A3Tt0yuq3E/Ub5K++4ALtl8AAmv1XvuI6IaFGlAFP7i
ttY+q5otpqh1admxmlSVzLn/2/mvmw9ZmiYgVTwEO+lxQZB/IvhF0kGk8TuJ
qiLfKithCN+c32yZsOfCL+rp9kMYDIOmxm1s8XHrwiE8Xnr+SnvmgjXtBw1Y
79TvEiLlSxXI9K7fSVTN0OLzKXn9jZNAVBSnvOfHbt2g+XhjIDUvByXYRRy5
2qwfksVaMTehQskEYHijx4RDEIfrfOJuMtA3eBYQ3fIV2mPzdEtCcwA+JdnX
61nq/f1mMIvArNR3IsC4Zx7RhMdhkiF5gm6DdmYUNxIATlthQUw5Qld3NiIo
//CS2irk5nRj6m+UvoA3YE4vUVl4x+IjOnWg3ucliokssBKh27a290u7Jfm7
NMB7JTSi0uenIcqnnQ2XH3VizWH0e+vZW146kHQfGjDMI2iegKD3vrCwO10I
dt47mA6Iog2ot/DujZbPM0VngPZBK2IbA+E6DNOHoAkXM5cmtriJZ3XW/A6b
/CXI39RFHEn89UVr5C0BWUR/Pae3smu5DLvO6QvlU2wQpByCoTB9xD2Cqe5W
yJfXq4rJ7LdahpTGCClm6cNfBThUV5G+3PrLzXGWNrh4sELYQrNfAizN7B7+
h7t/7SVUpZtN3D2UTMKXYfeG9u6zWPA//AW3Xw+L3oQp1WCUUf2R+RCvwG4R
YikiyWEoxbM0T1q+ayDhOaQFNDAD+zrzyAwCmP8TgOPCLYMGFrPANsY/tMfW
ph+J9ahb03Z103bV8iz3xt1RLVYNlTkyNhbEXlcA+OWB3IiH70Tq89fPN2Tj
obTgg9AVoz6QoAYms5ZWoXCpbylQh7z2jLzp3Jilgy0ohrkT1N2FwPBHHhHc
Udh6wldlUebZcEO1Jyq8yNfnepWXww9cYVVfyWYHOhtPrZ4HtX8tK8yFed2W
1z/+fZ/7V5SJEffqE6CfSjIw3DwQjwycsPEGaK/tXG/YFPcrhONCEZFJQSqi
mcyYJjmBIt0ubZQcz6DTBPtbKFv3TV8cuLnIRFZ2OYZlpK8KUwLmJdLdN5GN
LN+9ErNnqgoEFBxPJ0VzyB+xSlcdsw5vbFkgoI6RB0cKFZGOUyUq+ni+RTos
3eygiJ8hqR1z/ThC3Y9VyVEHSoGMU9xPlhe3ZQBOwuNFDiA98CnZ2mRvwhQS
rVptZ68CF9DtceXaxoBqPWZJo3FMlhdBc8HQZ7w/GGY5q5RnwYSuU8qmYS/+
A71zfBg/WhqP27cOuv7piie6Brql7d7ufC41Bf+LMtqXelfMw8/pv67LQPnz
p6Ap+yi24Waf7fHdAsOFkQmheZk0k+0FFSJTPzWf/FT1M1t3HFtg4UdFXodt
BIkY21uKLRRrJFat+OBqfEP6D18lZBBtcjZM4haPtQ2ZAIcwuo5U+uxVce73
PBdCd+V06OB5qC+3qPbuE/1S4SZPLqYXoOpc9hH6eW/rtpR9PJz10SnXQZA3
B78BoMiMtOF64Kj1mFZOd9ufqw69TRCpMobfy3Ny10AE5vUWaWIW3jDYACtu
8WC8jPEV1GipyyAxBTTX/WqQN4pJR0MEZ/7t9e3BSiPagiXdiJuoVJBRIGX2
SrWNik2aG6R9lzbz7mSAtaDPCzdzzUzNCjsxHm8Upp8+V99BlE97xHNbzz9j
nKJp3lbOXUEkKYDJsdzQzeNAgI7wECAuKI22ZU4VOyue5B9vSOuFJhFlqK9M
1oY8K+n7ch3xh3APRrPsvCj7WIyXJsSu8We8f7q0mQoCSvFTDbiNzaSgbluA
VmGxhfsVr/TRPFMCVf0peM+nT67Zxf6ifU4vjAE8WRJdfamBfBXlc1FUm78s
4nexxDYjOCI7jSPIXe9TkQUki1TA0YCd35Tpd4P1z7Ga0loKbkhp8gkGu4Oo
0lyyBLTHtYQF/RGQYFqPBu0MSsQ8wRKepigK0Q9tuEQW5++3DeSYleLhGdTO
cthIx5KkLz07GiOqKDXjiTh0iCb+fukmos64y4cMU8ByF/qtFw5j/ayhPn4Q
AOKgz7dSEZOCZgf1XyuBkNFP8sBgT3DUjfNip+ghHOXrSdGXIOrVrblioIhu
YooaHm8gzSJACqGeWzYVL11a4tCtNFNLYPGdKS52iLDKbVlYuy7CYVSiAd9+
rY9b0XkEkSMcwqbZC0tfLLDup7/R3uZvAvD06U30hKps7PwuLVsfpYgwGP1d
0lR7e+eu62VlGAfMLd6ftjOoiKX4S0rHTY30HFzYMoHN8M0Ka/roeokzMHOp
1Zg/kIGcJhzDCaoUxxoneLSPclVyxIvKhg6zHdwTXnpAq2ggLlLGE51kcr4R
DLbiOK2wBnV7TPijHP1dcXo3HdV9bPtazmPfyTW/7O9Tjl7y810SrYMU/PZ1
dKVSXMTcaVKNx5Br33Xv++3qPLiy/4921KAUdu1zgE4E0LRhfhmiUONXcEU0
91emTxKzHdls88zAWdjPBiLXyyHoNetwuQmJJlchQ/iHbdoGMMDxNNB73PX6
T2yhNpn6jutXU+3LwTf/KlcfX/ZjNInDcc0uMRKvfmTfHdMDn0wjrRikOErV
397o2dVozAcIf03Z5UeqFzsix87elvLqmiMHaO/cAD9DsKGgZXUoLMutgRMB
yF19ABmEeqZpN351hAp87VO0jWXi4u4ERTFlBonMs+qJ+r2i8Ozqf/Os9Inv
CVUvm9I9TQ5QXlQtzzdijqnRWLYhoO5qZZsP10AMQ8h3YExbAoZ5T1vQiO1a
LSCBeAKPd/VVedSFO9NEWi1NjYArQAdbDgUpEJ5LwyYTY6g8ORP3OszoKdKq
UJ1EeCv9KJK0EYNBY6evSd8pDB3ZpFctE7lI5rV/F5EPzr9QqPTI01Lmu9hX
nZUUxz6rAfCXrLiQLRRss1LpPX73plMheHi2C+mwLhEhwAQXj5G5MDc75x1/
rMMYZs9nVx2dRktRRmJYTjYUivGBx4P1oUX7K3qV6GgVFf4Kg/TrJbW0Y9r7
P2GsFkvjBnOSxieCE3GkcQYAfP0hWQvu1JsXVAWpewWzfbNKUtoMrswzSkGK
F4IyhrQFZq4Fx/5QhAZ1SjNtf4zikihUVBAZJRE/ZKR7eTukI49GmXF6kFHF
y2jcya0Ut+M3b2V1K096gw1+h6FoecX4q3O2/Sf9cY1v29XY2TG60MypNeVK
b/hNzDjuss9sRDdU2eg8BKHl7bg9WPoDvxiCsHeVSwZEVODlrX3XYEy5Ms4W
cTMMB+ah7k++il075d0DZwX33HhBegIyxC2gD8ytmK0o7gz+crVpeQStXAXP
3vY7dRTYbulMYIj8rncXn2rqEWJEueo6H48ENYCwnhG+1jSLK+WKZgLQjkSN
rVRHPCykSkowUDLGXVoCoI5VexUbvXJcIh+H6sjk5c9m7T3xH39DnMZI60R4
A4HuM/q/ueSTzr8qkWKJ6eQD/Dg4QxLZOzSer1U8Zr6Rzza8s4TXsVKjZeWH
uFrKpKu/mh7b5BVJmevuOj+dhBeXRkg/OV3fLGDwJ1Wj1+jBxhLrsbt7Fd6c
RNyHjS3CfDUQxDMufUAjutAy6fEK+nQRuNriE1DCJHRipCn/gPqA4TpmiMEl
jaL3gagaOqyn5ft/hjVXworNgjhR3L/KApK6a8uyMhCO8F9Z6S7YIQZtsLJ8
h+bpf0YgigANSdY4QcF2hlNYHyvcAhyOqHb4Y6R3HcfDAx8drPafyU/uL+e2
kpixR+HvcELlRbfzi8LavbJTolFYKk2XSpjh9Ypn6ji8d7AIXjjhvCWYpgeQ
brNCjo6bQgGrYLgjgZM/GP8pA/CSaxwSvXKzVhxF1PE9XGsa0MASh4EDpAZm
Kq2sA9OrDm0NFYwMEFJvO8RfcGfwKGDpZcpqhWn4b0+GsbfQh01vmMdimfvW
GSRacgkzUniy4MIdmcbDpQJcY7dv9ORM+kgiTkbl3rRL/2v6MceVg0Tw0WKg
eW4gLj4YC6gFhKjQ5zz3LNyYx62pkaUgHJQFvkPAPf9khVhrrfQhr9QKRWXJ
y3KAYgMi/bwFaL7MHa7IUL8IHfj0CdzuSUXaLfYxmZbs7hAHPOJ3JMUrUhO2
GktoUhmF04B1BWNoA6hm54LdLr1tyzyp3NNmvPwFbxxFV0SaSxCR/iZ97HBB
jU/gnLz4KgznGm3GQM2U3vz/N4CS2MNuK5SXWjshMEWUDoFbBJwHdSPx68BJ
cIQzXY0+7iJb7vwMA0JdcrHKxwsj2sFm3tKx2hS0O2+QwWRQppOwGzqFP7JG
wNDQx9yMGsL5DuKhHsdaiqI6diNCIQozdKqjXIEWGd8xbmRB5umnr4XuuOVB
s2rQ20qvRJHGX/6vqsX1tUs1XI+tH5H6rpknsPk0kkQTeI/NCnbBPsbazd1z
LAMBNMgMM5USWRHZPBZ/eV+L4RHJmrGlSajPycujs7mXOOpgfgs4sdKC2I5j
ZZEgdde2kzO4BY5xwrYRIJw3ptSdkBbJM6qxihDlpFf/d8rOdylsVbry+9uB
AXEy15JGTyRgd2U8vMyor8nYnx3FYlXkT3wYzzT8ddI6s2kBkWVkBs9Fq/aW
lxagt2FSM/XZ9szwfD25zA6QJSTWKOeHSAFfwIQoK/4IWpha9GbPoZI/ND5B
+VjKlpKWkKXM6Y0vuvt6d0JMY0nDbiOzgKGXPRjSZ+Pj4dz3q1mK5Zns7ZnS
i8Ps3gS0arn1H2+rAJORu4o4lppFe4Jpqeqp65BSndSd80f4iMPYGEYITdTz
Y+jCbQ870VQ8w2yKeDKFP6Mva3sZk412Gw4xJOj1lDYgkDHTsky/vZfnwBlt
MaKswFFVjQCyVaRsCWRy8P3ak8nVUs3QpyR+N2mjrU0wkxFUI6gR9EOmK9Jn
B4Bt8UEiylsY5HFuMLANFmXOHb46d3uEJD5/xtsUZ08LHHy3pIvoXoN+feuI
rVbQPNv2mRlnx8c8yazfGDqfiaJDpHUK/H1esLZkXEm64PvWODEoyTaMUETW
nagdEp/WJgbL221Gjkb4Wi95gOSiEQJ8GZCqCY2C0tKF1RwEn5rNVpGY/X7q
iuItaJW5dDdp6Ub7wiDqnWjFi5++q76o2qwSZabKftS3avoLRd+PG9rOSiLE
jWT0ZBy20x2Pyit7RH0sn4pvz17bcRTw/BFKJgQdxl1fzjy2S6clFsvsf93G
qRce4CZS7i1xwsNKDHkMnbfhssoy/cdMlSTlULJuicAMEcXVIQac9LNQwqKo
ZrxXFwALSrIQO+zMgUZBjWBffCQgpIszqNTY12mFxv9KVDHwiEXSTY3WiHll
MhJ3K9dPSyNr6pp859pDAfKzktgoHzInKMFG2K50tk/bai3TG4RjWrWreYXc
IrUnyxdH4S7xu25ovg3q0OIl8+G83m7Bw1/swLHtyHRjEJjDDF/mokkGm3DY
9QyDPDPnZYdTC7dcBiMDn4K9Ixp2eOUh3TTnpOpkj+kpfDnoO41t1SBnTkbE
QEhXz0T1tRwcq5vSx+4hxmaDXHYkzrC7zgpIYb7FoYxTn40Q0wTf6gQ5r0I6
Bx3MSBiq11YYpBEJDJ/3MqLNMd5goSknTE5/ELFiSLqr4Oyi6X5q2CmnikBq
vtqnLIiqPl0cZrdQv68dNhstgFHlq0uj6zAZo/761e+z0wzy4EdUSx0zsVGj
5IFC+uO6vUd53eJ5PpIeOJpEe7b/oknztfje9VrKB8YeJDVEUAPJ3IDT8cC5
aJx5Pl4y2nV7VvgtopDLUA49QFlmeD7AmqQNjjgG5C/yY+z1lgX46Wjcu8CU
0rA3irz5YusTjQVg9t/iQTss15t4g1k8Jy2Y6lysiq9VPPhYAzXhP2T1WGGy
YGzqfV8rT1x0pm5osY5LzLmufeIXczKcTqVirTp01cn8W5A10Z47o0ZeCxcA
Lu2jMILnuAlNmuZKSgkFMvNhDqJkcssZxyMFrsUk55ZreokKSc1y69Mmnodo
BkhMSDN9lmq0hmt6wtSiM83RuEzgRYyUbdeOEu2XQVuquuBXV8CI3dHU/5Tv
EhmHmztUzM9oSyDwP1CJQkKhJHpYXDogTB0kldngz8IHuJ1ePKazz1Caw/hv
5HPQWg/hqh8mqhoss43rrO0e9AFaC3btQN8EKtYlvTySbRZG554KYdvJ/ia/
kNLyGwB7mjwF6BIs93NzIa2mTQ335Aao2ynDDY1W/xSeY66ncEwvYM9t4aad
mL1rqlKseazz4JMUDA7AC25ipznELmVPBwpuNnnApieNcs+1xbBa5L5Zajox
3jpKqlOb+uujcFpg8M0g0Hhf9kAmnqVCoE7w8W/TqX7YbhNx05Ojp7IDyii0
DO2TE2q4zdE0hSEwEwqIeRrr8M3y3dIpy1JQqzhwAvUpWchJE1iUSgwZtFk1
GbSGCVO23q4PcLHmrrHF4pXl7Xyirmt/2UoYJW4N6oMrOxaMP/d/9JmcJRsq
J4r9U7zVb8lO7gjttORX2+UxqyaE9QF47ycFKCgqMRNJMRWJ7u5jTOqMEf4o
NiTYL4V1E18azOwnGE7nyu/JbpfX3tJ3SrpTsNavX1AwdB1N6xc1IbYH5nKj
LbhYZSyJKN9alHbnmSmg/E+TEujIY5bcsT/rwkJTe6xcC5MlAZhF4DoV0pcl
SEFnZfojx0VzT9vQQhBTcREHcOa/H9FL9Q6PNu1WcS6qnmYy3muNDxy60Kt/
fWagsyOlP8TLx8kTTFfZT0yT7X51lmmsVvfBktUY41Pl7hpWG1GplVd+vTcI
mpXs319ZhqZKO481XEh6JDn0XuVp+zxMu0qUn1gm2pfq3SHHcOY9oBaXMyCR
b7hb9pAK27V4fGSKfZtgSLbEJusOE4n2rD7fW0hC2VBXGR1TBP5AubZe2w6C
C7yXHF7Y0SDWdTiiGTtPZHROW4roZ6Coxi1wDRiKRNYSkV+kKjvEEdn9ssez
to8bSfUOiNnC9WQwm2C3MQcq0D3oawV22hYixW+rKE6rNVWr/42wLjX3NiQI
WtMjGS8SSHVaenxjWo677QvPJuBrpOUyHSvCL2Jka/fKmmyd4OMFxE1iZIbW
tLcrVdJ04rDCS3WZJIbmQRFWYhfNg9467oVN/f/bux/tSSh1t3tV/E3VPBVu
Bx7MR9FhmcPPheecX2EVeQvAhngLxhKvhhn+PoOjSEt/dqNRL4a7h51XduJu
ErVjBi4SJVz8ohThDoLk8s1KTOHhVpDLaq3vquvykAuyPl4shU3ulUbsskJH
Fryw0TPecFJmkedzgk2WM5bfV0Bgf9zAgyhToyFR49HoYDTi4biAXtXZpc21
Ty0SqrLPEX2NH/tWp112cpKbS23o/vqlzu6HIR2YI/8+A70rCH55QwXBmF7p
Gb1DNKq7qUa31lD0a49bjsa9ZhAfBwUNb1oV1O7B8uEsvW8xlkJDxwZnX9yl
Y4Yyk5OX5lvRXkTqY/YNiuHEcboDBTwfvqTX+BSx6ARcYxANayLk810rnOVM
BpKdbMLcKAorg4cYlNSkn79jpQX98Hy2j6QZhKMemyBwIlwR739v2AninYiF
1l7zeN5lvO9Brc0ck27buqhj4xffML9s2ye3+Ddx910ePDRtLv2jNwFNiJYR
bvKhG6/W5hTnhNIpqILJ85/8a1lUlKJwplfS9VrgKlUhoB8pNQJFFQivjrDZ
x+r8by6wHbVTr4Y+pdDW26tYj56kSnjI4R15BACXThkk61XxkRBPSoVTG/Vc
8ljwzBuFdqLg1MdDd1iZPKC9LflGdFPDq8QV28Vq6aiDXvR9kFKDfJB0ywdc
z4OYzLiwixsCxBKoCg+9SxK9hPLr7pzFx6bwL/k1zen12M808bD7D1SIrptZ
o1IXDb28yjVP+E4XCMH7+w4CoegtzqAXFUBtrh5O8siAGlmFsD+hQalexXqa
bArJkWKCS8iVP6wfd0GI6Wj660ZO/4Lm9G+Z6W8Z291PusCzK75Rv1iFio2c
U9DVo4AAhetQCpO0Ri/xCVfW6P+YyXy17KF9TaMuFyMw98paLYwfX4y+S1QR
97WdB4mUiIx4226w1lbkTgdvRUI/LUIHlZQa39rC8PebBmVIJxJGcRB3jLEO
YPPm2t/1N1mOtajgLz0m9YKWRcAJm6OjRvMbbmY+IY2gA4robqhOYy8Wnevv
jXMsRf6vFPkK9DyWDSsK0H9TC3IIukDC7gtmp1ARNNKAl0s6czUrbYttaEu3
Hd/hMndVJS/lqLg5xcXvKKOQ/r4ZdvYnxKw0APJN8QXOwaGp5yU+7VTOYgVC
cmhYWfkkNlH6UwkFgYr43lX8WW9gqHW/PCEDBy/TTlBe5yu+Bs/dgtOqzVF7
lIZ/tiCymVd53wycYJgLJiAhmH92RJhzNgDX6dLu+GcGiLpdDwzhNiSMeTZc
9fwROj/eCGirq6ZA8rCtVSLXiNkBf9oMmkWaJSXVN/8gvqe8ARcgjmeEYUc3
9qdKoDXQvxRJ6RWHeWSepDRkcgH1RIY8B4FQb1XDGfzvMR3UT1n38Rpqu9Cd
LaRkZ2m6N/IMmDY13dbDnlLCMq3h1aB7HLt9PFTJgxirrY53pYEqPS08AMZR
1tnNgxCGV2xEjT/ZQvUESTN1jhYUIg8CPArtVbFg/O9nCjSjE7iRT6Ps5YXJ
a1wXi6HQgCdvmSZ0NF1/r9XJ3zww+wriAvX+8X8B7v+EwaH1BAgcoR9yy+ED
Oy0RpqR5Q8o/B/o8J7kCj7aqkt+EQUJVRDpiY/EkGAOun0ONE6bzAQOIYsIR
vr0OAWVPsbFo9CaazaLgFgLDzB3V+40SW0DOD3+/cYYzWQhOehzn+2plx6cM
HuF5HorGs8HpvGNhbkqwi3ZanD01G/24jhlvnHXPOtBcT90S4LzpqVCSJiCo
gGnRY5V76DCL9bGxc1fg/UulxKK6kn5gkvffl9opBifMtGvSIzGSi5CNGVYv
0dWY932BoHc4DXZnfgfUMXwTNaOFYhr79mz9nPX2XAiDKxty+T6kSGaeMhkj
VeL/50AWLHMgqgOfEop/KM/WMnQlobx6z/roBAWwOXqblF+ExmUV0R6mze5S
3hAxLgNE0NwxHrVwIns4o6CC8U6uG9qNcRiaY41uittS3fQV3MU0zfAduKX/
pdeP4EDOPodHPkMoR83xYMrWYjGbHNCQop2OKInjWrcH+caAb7pprpnk3mxv
j9Rx7byqrQcIVzSfc+4jFZx0b1ycZ61T/nuY3qp/FOaDFLhzX+r0Z4Vffl01
9Q1v7pWfWhtN4vPKdLoKUGj094SOWSApXMOwgiFwxEwdR+DSu2IeET/H91lt
/oLeopvH1mNS0CH1uFaz3tLjFJLmqUNWWRYsiMcJFsh12/OzCgfizIGkTTiE
z92v09XSATcuQ3V2Oq0pgFx8XQHSnyek1oTqfci08CBQwBY+MLziqMQl9VZA
af5gGX7P+2wEpqzlrjYW5AlsNqWPaUynOjiOfUlOgEMFbF0Krd1dKsvLIO1X
Ja+3X/cRQ6H0gX2dlfkDE99t+b2D0dxPe4Kc8YhOEpzyUQc6wUs7U7RmXwpC
pHwP8teIUgs6j8uwLsPiNvlNtOn4zKghXxFbO8EhYI9lLHE8ACREeOTSLfdh
ea05/zAGZkp1mVfN+NvozRpSfTX1WBC3sT0I1h2u3Wo01q2f25kpKa892Dku
5MrsT0ID7UbdHYnbGz350k3pdwTHs+rpsqpaCQhv36yhSVSOcFIJ+TgDPfMA
JJT6DhOYshTXFDLg7/S3IicJrRCfDHaHtYnSSd9BT/tJUqVj1Kml4Da8joSK
FBCVuttC0YiB8+LBZShyIYC6mYvcJdpsVk2v3LKxRplqjFGGpQKOW9GfCPuj
PJ6js8bSlgLn4/FnYaKeEvXWbZTh5vqEnVEDvZSRtzw6sfl9gGWQonZU1Utl
Ic2mhX+rC7yYFxnshCxUiVjMSfCaQv2edLUZZ8k6O6Y/4fo/6+ZH7g6MCzib
tnP6FPkbFvGKZzB2dAdANeJFwzy4FKdNXkPwukiwg0q/G4+CUO+hPM6oHcXF
MlUSPWQorVPGqrdlHY8Mgplpk7cVNHQIWIpffpWbgmfa0D0EHF3e5qZOJrKs
g3ylVwuVlzRYkBE2RQ3xszXysEZVhd4atx1Dvy31vOXH4aCCsWJa+briG2BU
EOGEE1HkNhldN7wmby3D294fyHCV38ZfALLvtt3yOu8V7EKHpOxt2d5BJA9K
Vd7u2yF6+L1Qz4b5Po1ur30ZgiBC+S4X0zrgumtIxY/1101Iesdu9BkOgr+A
jNkMwh8wWAkcVsKBPpdJb545uT7rIvhlkWOVhkEWBhUrW3JCrthK37ERfjo/
oEyLF0X2DyJPU8g3nd5IGRP6myMiVeE0WAlJLx/iOtMLPSD/a2PhFjYIoOW8
aeVfy+HZ57c+ckqeTbFKWqojXTxD25L1ewuAIrCcrOrt5KwJAV0P0bOM3tDk
/UG4k+351fdnli1HHebjCJIReRsF68eEaRrV/Xj/QUuWeX4hZv7+0s7kwQc5
idWi/ZI2eq32nvLV5aIGQ7YJag0B3ZArKr9nQYvJoVH6PRxfk7UmI7r3CGSM
ReLWKUtmSdn1WJvmFRMQke6EwYeIGdT6PdhVrnGzwKhT1e+GFcZje1eiXbOB
d7zq84owBlEAM6IenkIJSHCrmACIv7+MQ3x/1SG3ZTmFx8mlJnbLzKcXixYc
7jLyyECKLTRM+4Ns+Cdlk7JYytdVe8k5yIq3TOcLFw1rNSSxZQlTxWKq8lZk
hG+sEMB2o0ZpJd8rQHnlx2nRZM3jjZfTyRAq3NjjfXkNDRxrq232PQgJOcp3
vylmSeILOWxqyHXLigpeUzo6/e+/IAfUmxd8XlHJVenjHd3THaSpCOPVj0nm
j/Yapqf1gaDGqeOsxOaf9jhGH7ZqLpgr5IfPrP3nQ1mPwS9oPETRyNwIj1Gj
obuqf4LphPrViFfkrIrDtCh/LHenSmhIutN5Bvz/3w0zFESKij18Avvndkc2
K2QHStEQyJVepeFlT7AyQ3u7I+/qi5HPkTrQGkgzRTSwfnnRwDYS5uXG2t5x
9YsaR0QI/YL0i7YTLLrmiiwViwpQ+x2q4znxaqu1/rceExLNao6y3iAYnn4G
/JBskLCP279Ct+p9574DT16+194LumG9eY51DGMUVswCJclvtghijFxUG/fp
s3WkNeITeUB5JSUi8mLKsuTj8NYmV3nuaJXq502sez7mPkFnBsCNWFhPA0DM
/Nc1HEfjdR7s3oU0PY8+VGz//ErGx79Zc1QVK3JoGa5TozGkdSRuep+a8F4N
oGA/0uwX0dUmKrBM63NmpNn42+tvfQlewWJQ6EEgJYm6sUKsEmVkmZxxFTc2
Tp+ZReiUBpvE0J2/bkhgtEeFppMXvWsETgbHevXTkv5NZdVQIL2dRNDgstUV
vN21XL5gkLR+YgtbXls53ey7kqkjTZqh7KdY+JfthlSWbVQfc10RFMa1kIQ1
GtpKLqNxOlqnG6cBdv9HRn6unrnNHAs0cLqhGuZrXu/1pAT+tv+patOvcVR7
pB2d7iG3Zj0tSQTjtFNAFZGpFcGSOUW+oAw9Wu3SlBuWZTbEwysGaDQDgwW/
ex8lb8H51L38856nYHEs3Id01qPpqLJ3kT27nulySNS3JzFHIMpZmxOgcPZF
zBh2o801iqgIMBVuhX8uxJt83tjrxaCeFdvI/s8vFpNE65DS3vXnJ1Hl11U7
1bqPgZrFR6aXIiDm6xFqtrUqU27yiB3hoGPjggCER3yxadwwu4dnUhLim4pD
8mn+tTxyTib5sPgGcmwFcja/Y2UK1v0dd1l9oPLLluTOaHsnOwa1HRcggbmQ
i9PxXL3HAZOB0wDHhEWkeaMnqNEMnkCQmwmYboC61bfHalYAiGR3tTwrZ00o
eTjnYMPijWIg1GxJ+PQCBuq4rWvYQwjZcdVoPV7Bbuoe6miTOLuCFT+7EY/t
k5dDpgOrUGzTd8liqRk7eudPLP1wNboyhpNdRWJokEqXdNNZPvpqQ+yWS0Jq
jviBXIhHQQuHNYmq65YaXQPMfdCjH7wE8tD0x5IUDqSwhqWxjKkphZW7PJ0j
oSuXLj2TKBMnNHD9XpDQIIFw7/3NQ6VTR0HEyL8vwOAmX1EAYPqZDrwvp5M0
1lS2pklzerHzdieIuLYeyxFw9ZjJnW07rKHGz7Ska/N8ELD5+hMbywyIaUPk
w/kz251wod03FfpeFc0J+ukzVbsufKR2akiGhwPS9CM6vIB66BarkaQb23TG
7MNalhtLrbhk5yOhUiubCQHEjLUwXaUf0xIMvjNymM68bg87SJZ563Rc++q4
d7pTJvcmeQoBhrWCF9LX5UxWAk3EIAYsVdHXqgalRMNJzFyF0UPryWigErQG
8ApkVcgV509fnhaKmRHSlYKluj1x7zlXR8ECyy/UwR+4pow5hqWJcU26yYXK
iDV76uq8+DiM+hZKtqhKyEZakbcRxwKHJT/9HAUJfDv+FnREBgw5WBzduT8L
G+phTeZKswuHwpRXwQshSi1e+FSq5/iY6MSqx7rXJO08M0STOKJhtkLo+MaH
Zi3+W2gTOaxSPKpM0fJ89axy7C0eubH5n6mWKei/r2+/77X80GO6IWld+9TS
p1HNYrgf4bgpBDx9/gTQJsVTcvI2BnyhORFY9C/Pj9IIytdv33y5EyQo/uvk
EfE/Qj1IHSPpSCutKdbhG0GDgoXYd6Br6ne2uw6dTN8eJawPLLjw4g/YMeOT
tiCDBWECCW75gVd06py9LC95GVXut3F8uNRpkjv8MAHkNwsJhQpsIeA9URMA
byc5rIOybEdQ6ZavnA86pKUvwjfpvV0HwakBJnH9SmTbo7ZmcOHKJ3+8TojN
zJ3Dfg69RhWINfuk3vAyZUW0BCeNgnJWWrKIu39w9YY2nxfiKnLL/KBcE7tV
fk9AIKUgbv+/f/7C4TePlZ5axzKisFmlKqc1v68ki5hOh/T8ynmF1/6Rkqn+
Q60vY4GN2xxnoRWE/VJ+QzqYjGUtWbq048gLaU9DVwWQvUlvf5NWMEJns6V9
7FE1zJK3YOPtcK2GZFCxJeKXxOsxbr8BKzJozYnUz0dF6v2yrtkWbF+hgOX/
RRJJP/a5ua7wM+O27jWGO9nIZb39PABuzhIgO9lS5qx7aeZMGpjUYT09MjG5
eS/Wy+Bg2jbb92Zl7bTKHyBNwl4J1h6O5pDk9mOM58ZoKUljBIxfZyBIRvJf
zcmj1gVjN+VzaRBr7OVrVAP/E9wDG6EAy36Mf3IdAmeuUXnW17qkZgqRLQ4K
NxquoFiJpMjAD0aAuZGfZjE7662pKIOvLlif8DgmsnA5CAzNTuaHVMx2JK9t
i5/ttlHW/MMMWyNwnIWMq8wphE59anqlYpGRXRU2/mgcFNr2Grt5gyi4L+iK
9Y52ICOYk50ILpwsWBpHGwpS8uqcv/EO54iart+a5hGhvQKyQKOfFaP8Y3qi
Jkmf0xyEFVqUdq9IWV+TK5wo55XvrbbvDT33CRXTa0czZUgrz+DbOW65u22p
n3Ht3BDYR5iyEfYXeGc6BtHmAudwIfSfcZWRaCLdA/rOmLObZQeyz439LYgJ
3qJAhKsj8LvkgzKwnzh9CwCi0KX8wHnxnZ8rxKcdJKTFK3drYkYFdu1+Io9p
/gKTuGvUqUfdg/tBJ8Fj3VS84L250fH6I/Q2Ht5fQ9Px8/+2G9uSRaN8ryzC
FezH6pl5RpQkFp46FsA0nniqizI7qrOEaZNixIRWPgPEvDq7bQVDyj1wdX4c
M7fRHqsBRDYZ8qC6IdIxm+Ol2jNudZo+uUnL92m3CrgD5q/R7V0NtKq4SrQC
tZBAqDOKedr/ff9hfxE7tPQ6HB4j8FuEhWgnBKTvaXzNmo86HN/VYqZUEtQD
7cRO/tXzJo2CJ9LdOq/J13jxUsiAUw838IUi7EC2XIJwpXTK/cF2LIruklgN
jOWXtdjvq7XNUAQ1XaxLj86M3MreZwXlIhGNKYCK31j+FvRPJ4sTJSA04uDy
kz7Nz6viQpXMkBmXyNyaxoKY6q2rJkdZ8qfLIPkCa88hy3UADYnmRlh91cHd
K1fSbQL13eHQMdP/NyBw+23i0aQ+DC7AqrAar/AtVzZWMNCL7b51z9Bfgnsr
FmTD4pPLdRFx8F46gjEiUkk/Y90jP8bipyLIfzmVWEqQCwCPGMrb1fgTBVE0
XWiQPm4DmCt4uGQibw+evVQ5LRCRAxbrKJ3/lognmCOsgFAivu55LLo6dPuV
1u156yYlbtwBnAvH03swvE0hwL6Et6x6gS5Ye3vmgZtNQ/C+t+4w4vWhEIsD
w5i7h+8nl8A2yTVPob7moVUcYP/oGkNJ1deo5Hr4jtZ0mkkcCL2/D50UP7Ys
+MiIKaWm1bmZXNWn+J+/JSJAm2f4KQQf+Wba4YyBG5s/VhkWVJdhBlFbD6vM
wVhCqqhDsMLDAYzcAXxztNskFma4HibtnYsbJpoW7ntz7MfnT0s1X95IVPsF
cyiqvcvXZvIcoXfZc9n84DxxaXgc2Q9pc1q8zdUddkwf6H3k+X1KA1tyV41w
3hS2YsbJOHLsahwsjli2ZSMO/D4VYl17kh5BBlZtdorDmAR4VtavJgk6J/iZ
2flJfFzDRIFvEq9xkid6Q/Z1Yo0+/1VrUlbNaaKmZlDptOtNmMmJ5CuCYvaY
/efnHwbouM8mXIKbXCav7t0TrJRcyOGKjvfE6e+DobN73BfehsV+GRv6QMjt
7hnOxy77p7W8lM6nXtME0BVP/BNcryJ1mO2etVSNOkb1myspv/F9r3bNRFqD
foOr0Gv4k2JqkcFWOzGfzkZYXmtE4l5RQbVo5VWJsbRqlDHQOnzYGQEgABBA
CL+IXRJJg61+wqgJYnYNbYmE+n/dz2wmLBwV4a2i3CVglrkhqodyXqyB4Bby
N6670lB/BjxCH+TEbh0jKttFfXCbiKlwSxhxlHKCx81YbmqN2RiNekx+yuFx
+Koj4hVqdQX/hTrMta+ddH+XbG3rQayIZMXL8T3FiiB2ZZPvqY+9D6wbzqBg
NWOkonBee4fTPEX8BdxwoDtAPkBpdTvTSTVAJZWSBmWjqYqwxSFoMcnmLd1Z
Yiq8l95Xrd9GLHMcHsWlJIGUKid6jpjWK9fm6/Z8DMZfWGIWqycjLvbQnn4u
BeW0AKDVWIw7EbUIPYt8tg7BrFgzC2tZ7FdDpCo1DfAYW5CDnr6CG9/M2HFo
JMIUREAGvI4+e6lKiymGAn4NJrcd+N4nT35rWQZZPAUGDRHaSkYV579Q1wxM
cMAhTFFSOioaVnXbNtuLakZ3Wu+BTkA5rywda8lOPTQIgkEhxs1Wnf8/dc47
FvJYN4JB63VQu8hhipmgglKUsg+NVHPmQU7E0cBzo/Jdh745a05SSIDf1yoz
cyPvxzHG1YtO7Vz0cAI/qpMaWATEZxOecnH5gmepAmBcVruTJUHqhj/Ne3K+
SuCppmfxWmuRKB3YiAe/wQb3G8FOXsjl+bIl/DJ47jrGpILY7elFU9Z718N7
2iyWTKsA/FYsjDQnPpXBZHu3lnNSdmIHh1YFAYLAmHDNgszgQbr3Z9wPD5Bo
ND1IbHAJUyfGr9zM2HC+10sPyKw8iHJVVOqaYU196XP6fM3ySqAHofn5oAZB
yA2jBl28xmD/Ibz6kmgDx2Z4006y6rmRdOeDYjUZcU8asFWYrnT1h/F8EIip
dZvK/ucBpzdK1Cg9tuJiPhnLPRXiZ8B+EAmwrO/Z9HjijRcPNgJNYyISD0Rm
tcy7TF7Vc5gxCs26yFiiqAczK9MXK+U6UbYveTRh2ZtAVpbec/Z1d69Jdn2h
yOnvDurm5R08Z/BITK+K5o699vBNoGFkWcuCJQsTrRsF/TxHVtKt1ruRhsw/
LRqG0SFQp5cIz9IIzIM2s/LHbtfL5WwG4PfPnhiIaY6jnpVz7Av7fIDnQ5bE
ZFrvxMtdGjs9DUrhDowAVdCfKTcngp+rEv/lzpn3uoKezzMkN07HKNBjGCWX
Zz779v6tj/OyVIqoiijCBqCYnpvG3hmM55SeY9vqSYJ1kYmAm7ks8TT3gyH3
WzTeenUw3c7qFo6lVTd7sVR/J3SewUe8la+M7+yWzRrTM1RYRg1wW5gZW3Yz
/eC6MIQ9aFPHhwAujKq/Jt6v/fV4DFRiZkV1p0eahwnO8GENlSKwSQLbku26
txpp8nMU/RyxPW7lnvPh7Ka6mLSDL0iWER5TKraJf77eqAnQJqfzhQpuuPj8
2Gt/8ONPPOzgs4X/zPf4pT+vFs3mkuU7M39GD/BK8TzPaF6Zax0KQzs1PIMv
al6x6YDcfcHKSC49hhLhNQj2OUxmcSpKoGRkK0GJtzDEyQy1eu3cV3cAF21S
VJZg/t1iW1NW2PEXr1HJ6IrDA+x6UEXbgxz0AEZxSvr2M63Rll5jS3scTZON
+kWi/FBktfW4sGUmewgIM7ufAMn6AcOGY3j8NNJBSDNExZ7eFASU46EM0+X+
OCr5epX5I86i9yjw0/c/yk+r/TjWB3JMkYteSMzgOn25rJqkUOCExjyetFVY
H27+HcFU29N8qBejhpQNe9R8rTkgid4scRYLTCWEAVso0K4t8wMuOgwyV1RI
Zt9B2OClOIw5/BCqxFUGrk90ZfoNoYWyrg/xb5h5fhLrn2Lr8U4KJo678atw
6SLIsu0g5CVksKs0htkZ40od6++kyS1tg5sJtsmUdlD6uDWkkVlzx2HTpk54
Rvt8XCzsu8YwpcvKLFPvk2zqnkTCFXVR9tl00ahsbCkXIYqywxZc8LDmWHhO
Xu7auz1XZPLvfsixc3Kl8xcMea82hDpLPhRYPQu6gkxlwnyuigkF+X6kUKch
UQHam1M+OAKA5f8SxPlOLgWkEDqLV+L/K7ZSoscVq/dOin/Oz8RIL+ZIuoPw
hSa3GOet7+MxFluOPUumeGYFOeNu/xhjJsD5vZpoV5yRet/wxGqCxYFDjGci
i3QINTtIvPxcpqh2sZYvGJcBKTVnLNVsAlvtlNU/18C+TmUVqqP+QlJuxWAF
oaRfzxvnA4y2jIlFCa1sIkQtZYnVzbY/KtNMhI8t7UeQNH2uZNe3NMbTS+Zn
jW2z0quBtws6FiA7cTOKYcGB0WJFCur8qvVAkfgQ91XKUYwFY8+KBoiqB9rq
bHLtHfEvAoOEWm2Z4HosoEdoFxnNOc+AF68XwyQoJFAJ10wGr3/pdyVH6ZSO
tKsagU0ZhjSrse7QoDYrCuKjqAfM5ekdR/CD0jSibauDhXQt3cuHQCk+cm9S
PQ8tRT688ow8A5FV+JNlNCgsDkhoXFSzC9+77+k2dkEK7P6WvoG2+YSeP19y
7kx1cQRiPMwbtb9EEl3jEPKOztn8KZNGDtdWacYeI6ZCfXwpKvc/stamKg7B
z4Ytbfafy/PpwXn6DKxeOkKPGngxsWh5bS6VwAgLCKVjvZQb0tTiEUgYIVt8
H98fIdRoE1tkAXr/ZhNKE+ykeSRzYJ+GgFsod5FOhCVKOkLXT2abhb7pJgeD
FNQTshcZ64ZByvkLs4JxLe6fQ3dspvtKdN45SJZ4WtS9k7MHYxim2ohs4E79
v4sIVItNfbv7R5h0+HAaQDuUwu9hSF2G9WXzghhZYvYdexOMhfc4VG5T02i1
JYa84O8RREBwvujk3I7g9/Ye/9J0YFA6TW/SYas9jBtdl8KPykwDeBRtzM4V
qgQSdna7hOeXJ+wPLsfuCr62x3CowpeyRMmLdjC3q7AZ9Ybny/oRGgSnyWoY
wPEwIO2kGUV35X/Xn8FG4ZbBy5RSIwBiRnXkMkhW16i4zha7agA43AnD1HQt
TKJ3Q8f9N78mA51o6ac5SRkvyNBiC6zd7rD+DeIq2O3uPXlY3XVHwW8zRR7Y
cpFt4e8593PPnag1yB4twr0TJaxu4dkYigkK8nhInrn/nPoEDKLlJx84wMcc
tbGJNualiVVEX3Tv2t2dWNRuYDUhamYw4AGTp2DfVpAtj1ka/AHPXOE4NUL/
5X5yHeKU+vZtYX2yMwsXO3Wgmhv7DXN5WMH/MJYe0XuWdpVSXQ32RlpNz3QL
DTiwo4jSjOXGkvrZvc3CiUIPCOitcTmr0ZVQsrqTFUh8r/71GiW79QFJelhT
epiDRu48tttyYgDKSJACKU8QyYgZojmyFRUohu1J/KGjGt/sIe+DrA57tQW2
nOfD3u+WCbN4LXxfqDzMmOEwBkz+DgNhu7YMZFOM95UHmMOB9jXQ3qL3TIIL
/iw3xb3yTiyvUOGm7HJ7PMX63ZlZWNyI4uLCGFG6q/3bNgoZfmyX9+gV6O8t
6zaWAFd7RmK7y1SktGm7seVELc+oSVDLHl0t7tXEig3aGVL4ctM0YkchlGq3
87n3j5giOQ/KlmjSzSM+u8jHDio/sI1vv5ogoj5T7rvJOVPXHhpDkEYxHUqL
yB3n43cweuts3Ka24zU8s41OiVvy8XbdOCUl7aP+3KnE2K/7aFf6F6Icddbs
62nvnbbiPMIXJkws1l3XekehLgSAe5I8DLFeS2p+x0OyDCsY/RloimBbyyke
dFfezUAN1MC9Sa2uweWO/gjwNFAftRRcXP19rqxIw5SaNQ2aO6dD9IUsG3Ut
zw+iJvpbYzJaMSsNAeYe01d7Vctb7YbAwLfCUGOBR7zb6SzZeAittXZ2ohHE
RCMXazBQMVSwO2xfjiULRisl3QWDM8VsRereC9Gs+10+swpB4bqpkAaCfqgx
qDqrI8OpNTmp08XOutvDPKnaGn2O1Uhe2LQVbyhwOls5TjOVbUgKSwHtI1FW
HS8wqJYUKHtqmAixqM2Sld9gNHVTih3sd5gv55ulSBJzoRq+IIQ9Vl5cBdM3
TEvQSYAw/zKx1CVV7dy4UnRBkbPpZugb6dGrexlIhZbXJeHGQMZ0qheg/Bt9
GUIHoONeUq9CZDp2FseMMCjP9BakPnhfo0kbEKCNCkBZ2GFpuJhTQHiqGDwG
edeQMiuN6A0tzjpBnX/xYHJ/c8T6sM4t2Q/AbafTOhMtEeX2O8D22igSr+Dj
73FXUGzMoEIAPsjWvTuPKUV5uMIqCbDSYp99CiX7HsQ3/uFt58AuTEQY7fYW
HF+6BjkT00SB9QF/npwHb7BCpNnsfX4dEURZu+kyBIEI9HgWL+cf7unlyB5g
SB5Km8wY9C4E0UxeKZHqB9eoNvUdrHvVWBswfNcU36Tn3v2kxRiqUsreQhOc
NXo+oBdfZ7SKZ3fC7x5uczUhmwe+GoKXByn4iyKNPTKZGVosdMx7izLyJg1t
eL0dJsaB2pgEXA30J0lJ4KYQjlrU/1FdiB/sjZ4ySdwDvnWaecd2N/01svgt
uPOGdRrsOjocjlDU15rnFKrWJT8dBAcZM4q4stcCOUN5jXfnvL+0biQnTP0F
SXoOWdhT9zt6+B3R2tGzZpwLVwledETV+iO82nPcg2eoTvU6yWgEk2SsJ2a9
pxlvokkkvkS0toMbgu2BLuZxrHq56oXw67UyyFQeNlU1MEbdlHLnAatRfjI9
wIRN3CuOHydrKea92g0yWSPKhbw9Znk4ibL9dP70ojkc2PlcvbmdHlse8lGW
TBRLPWWpbPLBoVA1RJ5FmqZ9Kix+BfaPvJfcQEA6rof69mOHf/h3jBwGf/hE
l0MqpUlPHEbfyPuTOEalXs40pPd3JPyX1g/DvWmm7tnsISyrq4Sls1D+WCRa
v6vJcjkOnbgG5+u2l69vYYfsie4yYHYH9rrxljSdvMvub1TDWVHJI86Olfcd
6XD2oXJukViJsIdL7u2AfZKJ8qVIj8e7ngfxYN28nfEP47YYHuFYIAJ+c6+q
J9ulQGWjJ2/SO2w+9Bi0eLXQXDJfjkHuZ9GEFHpE647ID3xQ6Kl3wGputZGy
on4fx6p//38T/alZlX0uyd1KM7C3bb5vh6cKzK1CiHG4Opl4c9FHzhWT3TgB
FiHR4YalapsnP1D9BUxz0biJokIPRNCMGMVplkuCXRG+JLhN4etsT16CdaGb
CJqVPZZX3mFJid+KIlwGxIZbEwdKqjwzh8pYXkjz9MJwZCTjkEPvZsMotDGS
Ao5nsnukSdes/bS0C6q6TOepKJFdMZDm81/wsGOp/a3gh4y7z79dLEuxStUK
c2eHgDMKuiAUrtQMfktaYRJath3ErQ5n+sxmkDkac7zvjdAiypEZGe8Xxiua
DjD/z2+oObq87qscpHTyBZKoNiAVpCRx5mpvDZ1aW8ccZcjKN8FBbv7VrToy
Zka6LTtfdA7gAtDWVJD9d53l61UHweWPtF0T8ja1E8p5VHZibRfKNCAGxQ6/
sWubgM9xMvUxy9n4inxDdTJgZ53UyEcuIvsWLvU8Vf5e/HZaXWCUQ9wM3USV
jgSFEia5rat2vKWstHLqmeIQ6CPnK5E+GwZ4yqQJ6+AFIUXLFSm2a0nts4c3
0MijDDWlXPMOYczWGd4r2x05CqZ9mZaFpzZdaNhnOOoUdHQ0r5TfZ6vSFqUM
2irJktdvI4MNzy/z55qDjVg0vfpOgwvPpWo8htx14YPxb+8yfFiRXLuE9kgA
sw3VQ5mOiQ3TCzrNw8fvzSkmYmHc0Tw+7uDBTDNdMgBvIwpE5Wxk3ddFb8Vd
4+cZMMHYYLB7NGTFP4FXsMIc/Adbsqa7Zi5KMqGM7sbekrfCUbynOc3JvnBq
hNdZs0KuOoxCEvsxxlWX0JKql3L8exNbrbXwU6IxSByNbLNz4ovqYjqa2DZs
VXasddsAw2tYztdy2XqX5Qh0uyiCAD4tqYi6KlgYW6TWZR+jL+eZBPwOecO8
QtckfMf9Q5HUrHvG2v1Z0Njeq9kZ4+nlQIjVgfwe9a4s2Rw9k9o6P5szR9XC
gvJyy+5DkAmdLSoWCDzgHzJsQOVSgLHhmHOnHJrpzmz5C5xhTXkGFTqvDMTy
bh/CghwVS105lyxtQsLEWnRgFerYfrwAXuyDyjQnVjDfhgBkyklwT7mAYoMr
BBGn5g0bzMpvCKLBg5bIwPpyecIJNOS9hB/ryetErE74ZC32k/9Z0nCHSM/a
dWvr4EjUhkDff5mpXA1bTqCNmWpgdqt/JuNoHjilwxuj7fUOdXWbnUzkPSVp
f6h3lf5bbMPCTtax0kxwlGQP0WBHgso+qxNbTI8iXHQmWrLV1QDEYhXaOKYi
tYcTZiX13/2pFud43UgVnfMfMLGfKNZQ5YHTW85KKYfw3xIQNAZS0EMRukKd
YtXT/2KWQOTTO2V8I43NkhIveBApugO0evmyLWIzFl9mCZk6cvnOGdpky+y3
t9KCaQbVSXEHVnzUej7uzOrOujcnkfOPeGWfkr4RpE2eaYvAmCQxB/Yh/Z4m
DWliJde/KWi+ECBqkGHxm+GGD98z/Jcv6yeuhS52JtqCxXq5vaZH3wlVs8/G
TwJxrZ0pmR1yc2wB1IncoBjNgkqC293rEcj9eUDq8U7cvTuNpWHQJeHkWy/y
576vwzEdqVdYMAEwSi9fpmuRSgDdfFK/dUEQEPx5a6EAH/ud9h8vyl2c28sB
Ky4cWpzXejYUtsd3cOEMvLFQuoQSPbVzYkgyB/T23UwipdJ+LMpB/Fl8g6JX
bP/HH15bs6RdTEerfntSE02TyiNCXNnxAaoXOKifEQb+18qO+m0M3NKsdWAx
naooiqXUd8B1oIU+uaQ1b47dR9gK7x0k/l9UePPDXTNeh8Dk1261A+BHpFtS
fL5OngbBTNYRPuNMtw/tKa2e3pc61PxkgTszOqLynUXDPrRBQ2eURbTYf+mu
tEdp4R1BUu8GO3yScACOGFDaW2Qf4Fhw+etMoYPKeExGpszwGhN+ps/ZbJO9
kqE2ym0Lu75JnFJnPNLMfmNg2HB7cz15pfMHkempmDYKgt5zRl0+zSnSZPcE
7iNHagD2ByXsEnxmG6WakwTkcWOXvHOhU/9lMKvEuM+vhrg3lWyHo4aEdnYW
PE4bscvDtI8EpTlibCqo0VDClFe01khfzJ7NPVqfnaw+0PvR+GvciwxhchU5
jMcPBmME3w6pWFbCzkQaqbWlyzdtMeTtig6HUHZCTrvOZ6u9v7FQnwENrnPk
NT2+tWWEEhlHgDw9sHwk2+DyDqrprO04CDcI1Ym230Z05DiYLMErIRBsMO5U
T4NbiesqwD3CqTZaxLY+yfMM+HV378M9Tl8PNuP5A9NVzYSkN1PsnRHagBdR
kcEe2e6UXzFDT0vV2qWtJnUjI0giruPZeTnkzLobiJuQkK5ppRVyg7niVOXQ
J70zCqIzLR37U/QGthsDQxjPyQ0bfM12SEwwQ9S/O2iP+PbC32p/dqnSER+X
vFFVSnzl4Q2MgIdItJw8DMuR5kE5SQsZ/tbHUgoL/HVFJdDTZFGReLEYRN+U
1frEoxSGGg0crHKDD3VJIaInHww7yn1lFMsv1vptjHNDc5KeqRlgUBr7xGV6
/SPVy+KjFVKdnZUisf64PRhMu08uVQLzb+noSn0CtKlaFpH7blKBJ11fOtBh
8Yn7j7/3sEeQV3xta76BIX4Cm6lGMCOAPDn02iG5vunvk0L6AVZk9p6j1rP8
uAtGzjM3XyB3XtIFPvnGBd/dg+5kHtQao6JjBtwFnw8LspRLNne5aC6r5wKQ
4NJmYYiAYy5xidp22XQcf4vshWhWgHb4XUqvLNpXYgXX0P3UDJnVu4M1pQKk
tdjl059RpvIOoFNE/SIz269K2MYpwAcoupMKA/doBtsZ9rU8WW7+Of8UKoo2
ovENHe9o9VnRlQ5PGzZL+R0oykc2oDJ2wBf2RoAzQAwVQX16DSo4tVeERTz/
qvt6loNWtfLHcQdSXrInAVur4nYZwFEm7GEgczM5BwnO890nGEwfZ2IFb6Wc
Da4GBCga57Vxxo1mFnFoN45zeTJEQGVTILPUvW/dmZsqJpa8QKmhLQgxjlm4
2wuXkf37m16OmlFso/cc38ronmG4e7/9RdfzDH99X53Nq56uFS6QdcGaaBMR
V/H5ZRUO6Yv5OfEFNovviaT/vskR/h94RpOqBGWtvT0FLybKh0fS6QjqeVlY
kKZ8Bqpu8CHqLt8xosxJ/qSYAhgdk3N9akEPtdcW6jQ9aHlV5g9OTZpZSvFA
kiTP0GPpcsAdeY4a+FCQe16idV8cVwiGodPaL8j/bqfd+PVqjDXkiKgYuzjr
QVyyouSTFxNEmsVIhHGrxTQ8uHbFJcwDmjCL+LbbExB+xf2oVujNV4cPKkK4
H1OdyGIeWoJ4ukJGY8YwdIduWOrv0DhT6gMocW9wqTJbyKlYWrcJcNifpJWU
PSbGlTHZkRn7/nIEegR5Qsi60LJ1EMXBq6A+BNKJlGKGrZQYEbg0mPmNhe4d
DgOG3qRsXiKCPZr8PgyHbNssbuo2bmbHjRfkAn41iP7u3cO9li7oYmybGv+2
ovBhtP2lgQAe4boj6s3S+CGiXXPTW6j/AOIs982L2LA5a7UC5FJdHYPMrmrU
Z1AxCmfVn8qU7i2PwS1JbRuCGGUhx3xPn3BDys+Bro0pa2goUtqw4cdJ3ZcC
O1PJvY5a5YzlQZJXWHg+Y4Rn1eSG1ChmMRhoGfsKF60QZLN3TGO09pcAu/ga
53acmYxv/fCCFLTiG95AN+3xXjPjkpFwMVGoYdGn0+GeVJxwo4QDGxCks0nP
EwkKfuwB6vBTPBpLePyzWlff8O9hoiuJdL8hiy0vDo8+vCMPZ7uQSIKAb3M7
ukX1mt+CihKc+SieZzCjG9H8RtWRLmWsPtLbj7WFuPNs4db4SxPr2PtlIpA7
SGdY2XgzGc6g0ZdKKpM6JY8dEklvjLXA70FcR++29/FWNs2qRFUEz8rw1+PI
C6hPkEvJBhZIhIoS+DhItYzku4pWOOxsnRAO4kxAEvlxi9rC3D5RJ21DSVAG
+hgT6YLExYRFgiAByfavhH/rHzQ61kQGGUt4KQte2jyJaRSuJSrJz+mBI4WS
pQ4HGQooU6ocvTzL+MtB6DFzEXOBVugSUpJDW3BK6HeZ+Lbtp4LuNY3B4+iC
2C9UaqdAc+mNN5uvNJO3OpXhYUsxQu+zsoTNePOqVaYcAe7k5NkfdFBe4IYT
/Vll8PsIRC909JJnBBucgt2vGh4/1kSWAmVzlTHeBf8vU5FqfEPC7bcxHPl1
YgTlzGmhbQggKimT7BSThf/9kXLLqxv6UeoGHjQkQ7gvSMIdmB176dEWyglk
OdRq1Fzolfx/0gL61Yyk9YrjJBxzlWzt7gVRABxpuR81V+5woBLROVXvwyUd
irVpCfgRL4RTc7ne1WBFohnVq2BKryyun+f3TfgPf68Y68OeEtm30BV/uH+I
yCxN+R1kTl6+36IS0ZyaeV/8MwpEmG4QHJg4Uc6OYW8iBHDQramj5mGWFG7A
KmmAranHOrfllagZ6wZYZJ4SkbpUunnQ02dpTDGfnBxISFRdSk1tCU7pyFWW
B2tKo+xTh2A4RUCBUzkvpJWDOPCI4WePWKhfn6wrIcYKTkH/Xb621tFL4jSM
/SmLKex8QIdlwjVm0bnMNOMexvTZAJWqoDzFWOaA3602tu4wGrpCPQoJ10i7
reghfTT4dxCcAuPKdrf6tHlsVTQRCUOUdqiMZz++GkgQoL29Vk1SUz+XzVOI
+llBNHxSyhkPSa8To1Da+xkwGVwOaDpdjHAHa0WsTruE+Z1IX4A9Rl9+6FRs
lEyIN6Dty/y3Xti8nb4e1CsRyiLbAd2+0Ff40z6E1NkoleQ9hSSqgyZmDOd3
K/74uRvHz89dKFuJJ3q2ZArLKMIV6lLoYdpx5LwqDhMXSdKL4tJOWUyBYO6w
pJd4vIn32vOCfK5D2cC7I08R9HBdZWutVxDvM1mvKNLAPwaIeF+KCRxgtP5v
+lzDKPEP19ZaLkBf6QF2TWNsrRYJArhCQisH7sRQtIoKr2nyGjGWS/sk4MME
P1VoCCJ0BY4Q4PEEl1+CcsKFJo0F0ad6yMSUppEmi4OMVUje/MXMQ1FKczKV
a+Hfi6p0Q8KXGU9zCspwYOSnkxBlek7YHnpHzICOGDiexHP7zBRWIvqoAYKM
Rx7n1vUKVg3GZx+AJajRKs7XRYtShWMsHv3UoDZ2Qi+cYB2d9iBBx/KMv9DE
IhBuFL03EiPpBQpOobU2raRJzQlffzqAM2KJnZdO4rzpf8HP6k6RcqPfG2Iy
7132XHUSaPUTgth3EUztFwFpaiqckR5mMwe0MC6AofRKiK5rANrCuSoOKNtl
FeEPF/w1WekjUIAV6Lx6aznGoyM3ctmcXA7aO8k976oOMmuFhpfWVDe6r6CX
QR3WZK7RJanJSWnhRUQ0kUT2Edo5CUt9pNF1GvzzN2wI8nMhzAt2koHRsdWl
UwoSAxjuHWs7hJOJq5xwtF472riNvgYYyfHlHLNqmAw53QXXVC6pN5a7gagp
AfsxU8W3JelRW52dn/fna/Ph6lUGfcHR23LqQUSxJVM0s8QnvN4iYr2rv9PF
3LqFF7ycTqjoYMHGlcW49Dn0sFwMmzwFfWfJH3CJVgLvAi5DnFJGkTTIVhXh
GtmsXLIT0RclP9kc6s3DKoqRq+Y5K90kXLLtEGWgubdsOlzHqGdE8k5/iZqc
PmeTbgBVKKRvyoBa93tKAc6yCXVWrh+/xtoVSucdPMg2xJNvd5BMWyO6JyYg
6Qn2TfzqUMBf8uUk3h7nUTccfPBGyvklnPQP+aqJdOlTGJ4AxRrv0vKIyfGn
4H+xrI3yuRDpAAIo3ZF+77taStzwY5OL2TyHlC3YfoL9kt5G3vjGx2VgfXV2
U8HySCeNygAhWxzoadndUbi0vubYAqC29ni25hSjgoMNUdsROx7wkHOJDasu
IvQou76ABwpDbM4T2Ve+6P0KGqGeqOl0bY5pa6nfosODJNeZN76nv39QUV0s
8AdAZBnS07PJKkvkgkbtFfh/f7E0/wWOM4umJkjRyFlNVKHZbiUEN0kUu2tu
7dOSRcs4k4vt6z7h1l2r9bf9Q3jSDFPfm0YxRMYfqZKfGWrRpdGRSwe7qqXS
mEpQKxNpb9iI3tn4gaGQyZm67x4nvn3ooTqEmaG6DBwpgHs+P+cACSOjLgD0
YZ2ffLD3ymXgsKTTbQvv3SpujsSifWlOKDG8pteYIAkvbwHCuliT/XxoKrF3
zWYLx9es89PCoA+tS3XzifrpG5922wzRXYpjUI7Fo3aLSWg8yo1/64Fc5oAw
p1C9weICXQ9SUMPD9J4cx7OPxWR77A9wT8/WplVnvUFoMOSeGXm/OLgJIazR
wyZWXPCNHV7pKs29xHnirILEwfEVVfXdj3piUJDHjLiSRrvXkzGhTbFPjqOb
1sC+JPZCmW2EoaW0slbspJ0bICluk0aXj6YRp4dTQuoTc6hdRjrPbdGzOJyO
bnNrG4ohgjhAbGjANFTisSbDTBZycLARgkG3mbeXtS8rGSLdHH8UQzWgC2WK
a01DCVxt5Fz5DwFxrQLg2iM6lZmQsmyqEFzsWiV7PrgrOx9408lcV8ddRSLo
DMhkTIVzdQZJjP319tOSxBpT8dGKBNJj36+E6iKCCw/NZKGJ6GrXCuF/qvgQ
ltdRfPv/ADe9KyPKNIpkrKbxzLdflQkoajVhsyjwc338R+WIiDL6lBHZwNxj
YeGjkoyaCVsKLzDEaQGTB70iVpcAtE/Tt+qiTVgkFEJ/9uo+CtWZp14N8Ywv
h+6ZGV8k8VsVsJbZKyN7OlTJt1/LUDdM7srgm+ut6X6tMyWpKQelk7TYfqMl
wV6P3bv+yeeJIpuvRJL2inOpsH45j7PUNDWWSfZJPf9lQ6AENmA4JRxVyPPY
ukVfHFsPkBHg6RceMIDQgxsZVFzb9MThunljqRWEny4vJiQL8VuwLgsVbzm9
mJ9OVUfZbx7BCAw5/NOCs3OQn1QCP49re8BOaUOcASNvqhpD1Z6fnZHy4gtH
WVSS+utgW6Q45gxNn0q752fbkp/VZnShv81J+0OK8+sG3s4Tg1whjQQKYH3O
Lh6tZR+CjztyIqMaxVCczT009NK77+W/PBeLRPAbvkyPVgEKz3h4M8+W0Pak
SgK8XjtiVQnbHTsU3DK0Hbi3onqKtEFQxTklrrRvDNMq5R00QmWalWTGJ380
WihhCP39AUXKFXZ5w33DHP+oD21iU90f/z2ae2ylfGe3ARlwEhAyWxJoRy0+
DQ4jNJU01PVzciJSGWkpbooLAQQch3ixaV7pN+zuTAZenRPIHZrZdyRNwOO0
aU5/xNXVukl727AaJK+JCLmAZKBoXcGTEtnTkJ60MQ6yLjYPM9yx2sLEyMFr
NsLQgKYHRcdYqQ+jTjadknE/GdvFBjgkE2qQAu59v/BfaToYO3frLvvqrZNW
ZpAQrJ4gluZWkUdgiZGt9dAi23j+V3IRL8QhlHXPyIagLEAtMF/xplp3mRVx
mfoEVgejwjSNQoASetrY8dsBtMLqUUOrPetEqRNYiqqUD2jOUnRRQ6zVqp8T
jJQistXzaPJAbOLZsxz1r3E+nrtMbx92ZMeAvQnTXAPuhjbj7AcOjh87gu0o
RuS8YKAbxhf+v+pFiIGk26WFaK1AfN1iYrNO4IzTDp+XP1xmwNZ51EJK2mvQ
/90X+9YNl6ICQkDbJ9KjgtuOsWaAv34ZyM8j8GwL+TLyKKB4xciVwyFD93GG
KwjHdSD1uh8X1MzTS244uSzBrwyJD4QxgVMripDFRiF/3Kmk11o/DGK3LFQk
Tesq9DsApQkbtQF+45CyZc/QIEaBtgG2DDGj3UL+dSEdNCPt62GOTakld9r4
yEYB/WGKjb3+vW/EVvdtQI8nQ0SABPUlw1SzqnPsFLowNgDPuNZbIkqI2wU5
rHgklHlc3/csKN1fFz39nHGYK0pLegOml+fqmmwzRYysCTq0y7PswHNJgYH8
dMV4DMiXNSBC942KEtHHS0pHkqIfZQyLm9tZJHm3rVvJzn+MiW5N8X73vUek
4H02RlLbmt2kaukO3i71YPEzzeTtT/QMUjchYN061wIqjWo7S9gFeq0DZUNV
qbxOhFDi3PYQQSmBcD2rngp+dHnzXHWiEkMdblHmI9Sf7d6bCH8gQH/a5MDJ
usFFdOWUru9DNvkQC+nFUky0aNgjhqpZdJQLtxN4nSObqdmt6KdHS3vvLi4K
Xkqa3Go3r4MVdbdcjWVhsvRcwPPZov2HPKjaX3BR7qFHMMDP9616/OAKHfjM
Kkb4/qOD6HlG67AuFH6LyRsZLenn0z6cFWr/xIqJ//PD+q+j521zE3sQD8MG
tXDRMH5eJ4rtm/bZGVerzyHpxz77E0XeetF2vR6DXjk6XQEkH5pCJyiKgowv
3vL5iRYDYaUeAYbCaO7yqxKV5gmVqPXPk6pb2Ap+4KfapigcdKJyiWUM9N+D
NpMdcBpDjO1gWX8bmdkMk5fKULwBF0mVoFeJEJCEVvZ2gr7iaTI3uOYiNXAw
ZHCagVVUBxse+hxGmF8pGu3nbl6Wkegt+TjvcZBw0iinLsoSrc88qODGTjwh
LlEvqpVYT9TJVwyYbmhV/fXTrBdCwzHHtZDbycqkcayHQ9mXnZNOJ+LawHMZ
OwKikQqN96bThd5s8bh6CKpg+a3SWVk5VN9QHWA48hUhrHp31JIC58yVaaCf
owQ/yScRNGx3qaFADpTbEXDeHWBi75uLrpB3Bqj0Y3eQy024MdwmtOja31FZ
w6Qor7DwNNLs/wBpMmsXQ/2wo77ySF5EPF0NiHkjnLzty5oA1+8xfCOdWbY/
E7UUAunosFbVfiDfbzgpPofkbHgnVJyqyqwNXgvlyiH0UL4YqeRhPU5/kLl6
BXvh3WCICAFaB9PHTKsLAewjYcAeFFqWyGgRhVfiuPiXNQtBxecsAZRgQAQA
XO8qcKkcFy2R0ydZFYJ5dQ4Vic5zRMhE3/esH16tioM7Z1CV38x2FgML1SE8
F4o+dNSxehFDt8Hb2cf1XpJQxq8gK6wptSgy15VtZ+RV5A87NtdMqT9IhPct
h2XA5gWOhNf5xQKy+7IiMgTniIqozwY7u0WS57aj3fOHIY/kh5D033DazXRI
KZk46m7KWI/k+bVoZb+El7bD/pnLcLYSpAlU5woyb4ch7g4YCEOVQLRZSaMj
sHvSC10d3MUk6E6afjP0iHY9B7UnK2U4qSOGFYpYpgcP6ampGTrHFPYw8c4b
4u0rt2v6eyWm0uXg2BmsGyiBPzh2wzyb/ba8CBgOLLD8Meom5F0EHDFCQWgX
DD+CRIAtaAag/GzDuF9+lotytrU7CG4qYJi4rlIfqIh3PFSO0VNjOb7ggNV9
ttJSKhkRVDRuZjFgI6yVVaAxh/Lv1AYhnGKigWAcjak8pQ8c8wNoftMElWWa
Ng65sheTt8fM97Zlrkfo5y9UmDoe6fJUgXQmkKTmOGiB1kr6Er/NJeKxkgxz
ST7HpeScGlfmZpKTEZT8lc4vW+2k8icJBaiUfh/8l3hUA0wEME2QlA2q/XWh
zciwkSJkCy4VjDssgnqun2XQlc5Lk5iW/991eBv+iLnS47QwiuEdLQTK0ZJF
uRozr05KZikwwIqdhH/yEQYfL8Qs5REGYyUCHYmSoZbA/kU1Ajutjhl0pHCZ
MafymTqZkaT9trZWCmL3UKSacrC5SPHOyl/ZX0asGTARumLSTgiuJFdeBQ1m
SYhwA/TlQ9/seTe8ol2sHIlfJcCfZBBPmpHKbtpRplR38HeK0FVYU/LY7DVJ
hpuKh/rtHcArB9r4VD3/J0SUPXjTN1Hjob2uMW33qh42cTZ+FV7XuiexW3Vc
g7mhKyKo6f5J3hCyGijHR9jw8+PoK/tJXzy+ilLwhc9XKRRV8/H/lIMlYM0L
2n/wlLyDno3epmGzz8ZgPo4Ysykv38QgChSnLA6Z07zI2ZMDjduYJnCuHDw2
Y3XobgMk9HgVyN/R9zHyXRcM1iKkgMVO8TA3TPid/RKfUGll3s2jWHT+oJA1
/L9ziVOdSIe56FbpLbEIjkn30hpdfNewMdc4XP3axESAFIjyrpmutdXoRkBu
rLQeeNW9Sg4PvZ+zf/CcTcqVlZzkwPEq3vjAJW+reVZj3d4PY2Pw71mDvttA
hf2wPAZEi6lCSzxOWt9Zk3gg94BTuVcLvF1ahdVzns3zqM7rVtfM0p6Po1IT
+BKd6JgCSPnt4XzFV6HcuIXxCJIZNND9Pm8RH0vjMrXHzSBmNaElBSQYkkE3
x8JDB+vb35zxhZRDgzS1Ky0dVTFP+E6TM5K9D+LyM/e2LjA7FggP5MjZUvlp
FGyVwhQjGy4hVbUvD6Ox0Us8Qv9EeE/sNVM+4JojbpySr37DYcztFyqL1We+
u9g0E6bCBZFcHQqdmm43Rfdr27aJOpunksb9r2XRrd+2eeXw+shQSLB18D8v
KkEmfyZ4s4ariCinmfvvZEF76xM145GIS9fnrBI7aSPrM8BfBU3q6lKVQa1e
EjxA2NcTI08+D5MDwPEVHH/UTs8ryQsA64LW0hh2Xwsx2PRQCcfwEGUcL1rC
PW6p4pLFxfRmTcxKcanjDm0sUxPYs2n+XeXRMgThYKnXE5kd6W6hIjCcIgPD
+xZqGfCR2xJIh/1EEFnhHcrg0zdcTTQ14Q9e1OHvNnZJVPaZbhUyRcCEKI8E
TP4JwhUZwZbUDLjk19REjRywUpwJEPeZVULeHkiWcg4FidZbZ6ZXb7ifPtA4
K9748qmQXh8vK/iPoWbp2N5Ya5JGr+8UrfWwztMp4PR7TqgQdfFMVtE/B4Rs
2dYSLjTR8q933DjPGeYdV6NFMLjpzuoevNKhGOjJe7qdhjaZ5qnL+MdVmOsP
Ygwdj4Ywp5uzinREILeYeU25ijE1t9BoQd5ZCY+wpRDujPuDIgqAy6WhtMqb
EpjXcZEQ85Cz372hxLXrG8Y9sG264tbvXxeQr4+912QljuNYgWXD1Qu1r36t
4mkzapvrTFyRkV8xYCZ4lMcqGe8tOaT4qzMR3TqyNknLfsAvsGbcrcwkDjJn
vAoTJAFae4Wadr3AGy1k1544+A2oOnL+XuISN5j3/jxs6pk4k5G1g+zj2JrL
dqZQHt/TsFmJxMRrY7COyvEzLUbRyC0Aj7XB0/k34niKPELL8+4mef2cqMKE
jBDWsxWpfO7wxc5SZxU7DB5qbDQn8jl34ts/Jmv3GfMF8WtKS0uubb4kgfyo
8Bu1eDYBMBeMn2cbx5KA9cQ0I6ytNuv4Z7Eg1KSji9IcdaENe7sI4CBtz265
BadG5GlkF7D2s1KwjmXVrwPGwwBDOraeELwbkG2/S9ms5i/512KrPIZkJmf5
Am1LaZPAoCuwd9FboreEBQvOp1o8mnmhM5rchd4L+umE8TABG0xCMDURvncV
pX6sjFt+gjlO7pWcKYfO0dpbVIP061c26JfVbX2QiRcbkFC67Cz2JNd+QWz0
hva3+/JABMz8u5JI10AmeGfuR3p+RTYWp3ZZGtJ6xsYx8NFOz/NnyKOzgKPk
qqHsd314X2EwXRvc8J/QeEKTXXlJsdFfQ6wG05elVd6+o0PvSB+/Vg8F4jV0
NxYYJ9zJM4NgLJA73zOZTSaepGLEGEPBQQAfeeSZv+kp83xHBNbdtJO25140
BwtTFXEtpNx6J2iOZD5KKp95wdLUAnaUAQCck2/TJCRIQj4i0gPTt41XQxOM
vt0QZyQWQxaA0gginn7E/QRSsQQY6jwwMxKCdQcPoMhobPiuiGagWSCr/oNu
awZaBuGNIIcyIPjlpJdvHD/mPcf3RF1gOOfS9tX+7Eo47lhNhVLZUscP1aL/
wmZBbIQhmC9lGtex7zjEC5L+joK/JrVKVekWl/TDNfPqIxoYaJh+dsWiXh0r
m6fTm6cUUt9V0rY8EkhzzZaMcUf7/QbfS2BS7W15M6+JCRITml7EmKJPnM6C
d5HU5W11ZDK4Nzznd1HbMZFR4rF8cfPvzbBhuCYTvqMX3OfMB24E8IX70BeU
bMDfPiDVxC+mvZaJXD82VK9QA9LHALLfKyXnas0d8hY0EY+CeW1Lf24SC2M+
GSsbfIe2gn8m9Bo1v7Cn/EwujMi5ZKZiic5efwS3lH2p6t81039ysPNfcm/G
idrfwY35fQH7jb13/BmSh5261h43ObBYIefQKFV4thbtTW67LG3VZoz1oi8r
xcS9O+yIML865G2Eg0O1PfKPFue/HYWqdNHxhs3FCSqKdo4cOCsMX/XciqiH
7CmR0pgXGAbMPDwX5rdpH2yTjyvTQyzaEoZw0d6aOF/KxVwmlMSHZu0gnhp6
aAWZjebV5lBxkEH/EdYL6+yZf8bxgnVhIo9w3Gq1ZaLVqK9G/lSNjnQO3pjh
ibHF8FlSZM2Yl6ogayOxtPluqO6YXSjomGBeRhhv0UKH0/RSRb2ZLyAJvHKh
bHijlRl5tjtH+ME/GYXgcX6zdY6QVQZowm2yZy2XgsljKFTseO7jpb4iad9b
GFxCvomVXfyhiOCpltihY/cenqVBzROhuetJTleVFlb9WFrmee/hQP1CIGXx
2al1AUne5fmtW6dTkIrCf5oSWVhtTsrjiE23WFinUIN5TPOcORgTnJN8o0RH
JRQRH5BDsC2u17ln6+X/nmrkFUkm6pbFFWnyZ4g+Ha4rtpuZ7hTrPdN7/8l9
TZQsHmvIXI/CdATLkh5ADqQro+IraAof0Qw/bNSs3RYhPdmJZN2lL7Qu5Qr8
Ze8v+HCs+4f5XLcc0untETtLrx7eOOZT/uhBUSOOommhPCe2OoZNzK7EmtsB
YXJRT5cRBd0zUGn/UgK35VPF1wzrWtlYL53Wm6CVB/79lCpjilxjhq8uJSvk
JLwFTqNLy6e2K85c68gaKH22CohiR0SwL3fmZKQ+7sy29v1kYC9iY9NT4j2n
o80BtIHS7WpnokThQ6UpBzKSa3p44dHc3sGHumgS/NfbFVKPg0GXe4yJBzWn
pczjaxAZv07PJ6lbGDJsYOtbwp6B1oFO0CYEYd9myEfWX/dFT8sUDjRxQZVY
n2+15H8pK3WghheSrmYkWcEnSe5QTPPf1GgpR+1AK91cSTcoAOTChdwSGwSN
HHd4CR0ooD3y9wYO/gX0Sey0TVlpRT1eBGAbZsYnv+wc3km1+E4p7Bjfm/ll
x76KUeeM4bHG+AGsEFmOIOsGFtvbWrBxZn9RMMMNwktIyJZ3HK4gWBStlt46
RkIa7EOVavlQBma1Ann8MCXfhDAM8xdMw5+D5XUTXNPIN0zBN5sJcrGPtx1L
KeG9lLZ1G2rpor9Bc84hD3gutHYG3XzPrjBM2cgqohNY/wxMiCxvQM9fZshG
K8mb1kVt5SBi4SZ+ACW1P9J9RwKhoMZ9jhYcl5G42ubkSxexZXzm9OA7fc88
NqPnaGr0WNimsiF9M1yD4yfc4kz0o43XQFUsGG6Zhiqa3Ln5+tHycwrVi90F
RCed+xxbH7pomHJsQHdYARDcJNZjV1JojNnBduthLzQo8D/8x/yo+8AFkZy7
py95irsQTLRS6KD6W4v4yEMF7g9Twy+XE0NugQU4Mp7XzGhWqN/2NvFoQ9H1
lcuAdS5aPqE2wHW/5HWEfN6CW9yC9z7OymTRSWPVET+F66i6ETCWtFq6YR5X
+M4Wqinz3cc/BXrzIGu9C8y99FCsMwbJce79NaH5sThahYIf4jtgJcV6WRJO
U35y+hhhdZ+Klydzgf8Uy+6+/vlh3ckEN4H7ZZQHUll+ni9BUUk7JJSIDR/n
cC3V7Zj/zwkQYaXRrJOS7vRS593QH06f9E7UaKlxkeCl0Wdmxc+OZdKY3uD1
twkGuBPAq1VjKv4GIRcvhsN9/k4/jqJSYSW6lsQr4y6ns4Vv7SzhNKZrFsjW
DmC1os1nrLIRqoivYuqZCIoKbVC6VpVhL+BwQjunXvC0rmC2KUKuxQTmDPV5
yS08AutcN5JzGEs4LBp9xLz3iRA6GxJYRVm6dGwgvs9YniSqAM4Y2kTDE8YU
eDOiqwjWF0iTocZvj7nTt7Md09Ew18JskzaCPSr0f0XGwXMIItNWHzEQ9GPZ
Ji7uXxxKp8cMrLktU+t5TGa39A/zS0PHNBDUaF5k2teCb2SBM+o1Q1+YhdaE
pebIo1I4+o74tpwScXoN3Qn0mUjR3q/+YobShoX4jXEGpGmCFdNkNmIjZDta
e+JtVf0VcLcgMZN5BLknJoVC2W7CQ/WiJFQdYzj0tll6CuZeypN34kquz27/
3EQz6Pr+JHvPkxndCykSAmNdktiP/wacKoJG1BshSuKvtRmY8FeLJtMf9DTN
p8b+LVW5vfZ4+KPGCx7AFca6+GTE0hDohWyxk1TyR/LhdtXe6LmA/g2oTK7E
1zG4G+ChZdn4MWS1aezx5aTT1vB8H+g6ay/zj5s43NYBQI5WeAfv9o8rBgr5
bJaSEzeMk05etXPsjljwVM0T5fhW3oDf7zZ4MgnE/GOdgS0f09RGB49zmgGG
1C5WC+cAeILsRLjCKMMn23d3wAj87lLRNDOzeVJiPej8s8MZ21c0EEfnqKfd
kPrslKNHk+GNq7yICReV6AZaoTDTxLAbuDsZ0faAHASMsD5vEn92hNxNEvT4
U3IpL4FFjxjqNBB9+yBFj9AV+TrIP1tlsOVsLvI8yHjLh3fY5tdBGZNvmzF/
51TiWr2ygogcDCH26CVn2BytDbDZOzpFmiLx+fWnyAmn9SrIqMo4ZA8bEA0E
coJvRh2+Dz+SKWyMUpbUYzHtAsoZTusL7YKI9t1p0nwmrhKnKAVEmmtWd+wu
744NpNqCJPcKtFgwWouMiFUD14lEOkeYuHvAiXt+7edJx0onrWdTrmYmIb5Y
BVbVOjDmY8lHuDg0s52x9KdXFvz9PRVcm02T7OvngSjgytdB42VR2jLm3E9p
zNa/N7Gpa+x2bvMFDTxZQhTQ/M/XMH3kSWs79cVp/51T4fWQ80dAFUNRVaQh
tmYufeCO3zCtkkRJm+KopKpvph7IwhrYKjpV6UYKZ5XsHIKbk9d9qw7qHEj7
S2lXfvhcw3Lr2WrFXo6JpAc+rayjDB3oT9BAFgMXFAd2SVMuBsfMI6Za0IOP
mjslKXV+R1C2Lt7OzQTT/6UWcrXuh8CjXmiCxWFCi6eOynSP+iVEXe8aeCuf
O+8/TOeOIMdoMz77n3LsGPuWT6Ga57jId86jR+KW2y0n779vdnvCYCNRCctq
ITcaAZwjuoSrRNOdML40L37OsDynRL5gb7uw+SDVwvHfKBchiIDGm+tgCcRM
HRUgAgmHigdA/yogWIMuhR3NbNCaEQfaa17hm6NZN6HiFhJ0NBQCWbWIOeIU
nIQ/60OXL1ZJ+G62//RzglQdfsq+bI8m1DfTye9Kgwv128xUKxrC22Y+FPGR
htrED7UPcPmy+cly2BuLeMfG+3qhGcYa8eOUiW4mih0wn/Bom3d3zl9DxX4e
Zyq4Mm+qMWAl2xzuj7DfQ7K0iNeUiQXLR1RbQf3bPK5PWO0F2VmDOHWS1SM5
Fe4FW/rN1HRcUiJEuGq/+8WaeQBscFirE+VSLZcGAHWLoSwI2/ZUtcRV/t/4
kp6UrdNOdWIXXDBbNQRWAWRT4u8OKrhFrOW1+nDlgz617qYPhREHoAxfrYSq
TG39olmqttM9A+Gg+VWr0rPkS8UbeuUisozoY+GEfhCYizraGSrqqslfoWVU
fdIz0IJz1m3SpU5Pa2+UmqE3ZCg7nlX+xg9WihIxK7c5/0HquV+UW9lgDiDb
7AR2bJRU7zkK6bxLSTZe0Mh3gcdArls6gQRzHnGr9rCjpUR5XncDZXLKLLSP
fzyUqwlR+9u7veqWS/t2moo0cqTfblb7I8WyPqKeQsn2jr3S4B0sWK8HtJas
lKX5qbn6MXojPz1Q7X54NcCY2hCGP6gzptq7wNCh4X33FkSGA+A+zLfaz4Jd
I87JOkpAS4l+KEJPKUACr2KfTZGBZWbE3esStYF9SBlHJ45leGneSAmGoSWp
hRpG+fPSSALQ61WA6FFRx0nDrFYuVmE7zHypbt0YmumQPthioPx3dvcXufjA
GpZl4DfDFaT3MgrnYcoDRslS+04r3diWFpRyXFClM4p69R8f17tpUPQcnBQB
x2NwkSBY8+NGYjb04nzSI3cY6e0kcHl8i/QpZGpUauM75Pm43stoTFswRNJw
gKBdHw0C6N+ffSq3mVK+GdDHNvoqv6fqmgj1MdxgLwzQhzqNH1JODbP9Ibsr
+Hy7ahMW0eD8gWUweS4e1gSBNGJT1RgLEA3S0tQM2u14+oxdjL4QLZrZtGCZ
7bPWE7CSlhcO5XmR4wKq2OgXoHF4ij2z84ky6+20vPpri9qTSDjfXXzWFbNJ
xc0WgUWI9sGLkPVEv+XAttWdMb7uZKCraUXuTVK3GKtdy7DiYC1RISit7EeA
Cjei/p3vCq3KTfjHmGpItE87ZJZ7qDkMRRNbdt4Y4xfnOyORleR7xaYka9BL
q2bDG+vuQKKTTbgREldDIP5eP8G4brbxaCdVKCnpSdnZOpopn5RXkJ6IzdUp
5seFNDWyi7KskKNkkM9hNu+f/XuhB6XXpPLZ7P4rRJMRdUaZGTYFzDYhxrOx
WwGp5uyeWNSER/yi/LGJVNP8qMDc7uTkNW9qyz+EHo8YzCRlofir6aDMT2VD
RgWtqnaQy849f62DcgTrZ4ar4CjF6+SOtbaMnki5UuFCJqA4f69y7rsblrf1
NeXFI9Q7JgfGCHTTG32LPMQ13+L0zNjpFPDWk7kEJ35kyogG7+xqIReCt3bC
1Q+x6rWbPT8j3IVM1eQzZnb7iceQK1VX9Ixv3GxLh9D/8zH2xbSH8KkOBvIR
j+mJG6HmkwGEuRS/6xC5yCj6n2h2+gY80rhGyJCNIsVaxjp74j3x0PUuYtGc
vJeY4trw9Omc0BCHANaNCDH6WsbTYvGIL6p1KMoVgsb1IEHNwSiRK2RBAvPs
cCxeixXzbZ6ZyWRK1pCOTbf7gYz+1eyM0DdvdLzjW7sGnoewGkrXwE3Xe+9g
WFqKEX58JoB81Ust+MqcyoYy0ExZGP3Sff6UyxIHBSSL/9/ICxX0eU04gGsn
97TWh7C3MVOVE8RflvcyOUAGgFnBobb33kQdqnyLa8kYgDUEVCApnoVuAj23
tfD5O0hKUvcf1WqWS8K+wrbpGGASTza2cGt4rrectDYJMEWFkG48GVqMeMcW
DO+yCL+BGap1n9wr/dfTsknWw9fkfGmbytPqcj8of5evQSv2sGKvGdCK1Te9
T3w0kPZc/hzmQ72NUqYdPbWOl7qSiOUj/aAoswhM0JcR9L3shZGcBll7tckv
tMNzp6YeBbtf0b2fx9WGy5vepmW558nTjf6TmNdX4zIs98lqWV1Uxc1RukxK
UXaGqX4KehC6xuwHwNwtcizML9HiKlRGUoNvyhK1lJqZ7HhmqksNkNo6FRwV
cz3fndWgqX2jhJDp50AOLjYo0vOuUQ3aOdZ+eATMRAUq/kPL/WWt7V+k3K9f
tfV/uxlAO846RW2RKRznMrUIxogbp97Xe+zNO1SDzLWaW6CocINO/6zVeEIy
af2tdcJnOJGE4ILHV5pUlvNykYUijps3sbOyxPGzwMUdU//khd53vLDBaG/b
XfgQl2DriYzN2cwp6LnjApI9XVEGP5bIPm9/17VHttIgtaFhsM+f0/2U5as/
hwEhSn3g6BgESpvUyvKqrdGzWulum92YfPQ8jsMtJ5PvX+MBdTDkYCb2XWxE
kJQM2VMz935LEdfeFqCp9hbj61FA3c9L9+kUJiaaA6+eJQ9NqDckxAJS8M7s
LL0doRPlo2qWd6Rg9yOEqgqQA+RbflrV2AszEsyjzSaOk8EBRUn1AHPLLJrW
yEVYb1fCOkAK5SNoiaIOdDXcXg4QFXoKmByoPkMSB79M7jCOpsRfu25Vnnt7
9l6UfkD/BSvZTnUJGV89TeIW3I11yWR8499dRKeJETyMZGFvyjNezNgo60xz
07crkg1bSiY4zf2G6AK9qu7bSFtf/DHjrpn1evmUsKE8HRuvqsTNDgX7LUzd
+Jgth5tI0ARtQW2IK4aIWY27EI+lKpcayy9ezT972MtQN71UyyKD/i/hv9Jt
5C9UmS5tnn7sty9eqADesIcvrgmgKEjfkrBTr01CWzxK4LBQyhn7cqld45lZ
3LgBVqPj+S/4x7k83BW+yRADgJoQq4sQMZMQEb5GXGs9BnmDaDcWC762LYrA
/CEk0sInk3VOI8fx3htGpGOgYhNgVWF0YTCt1LchJP4TKROvy5MSoqAeBrz4
C2N5MaxfS/iDtNGtVUvt1JqIFZl+W63uZBsCmbh11dmMJnE6ZWOJzDgn13wB
yeypH1uwYZI9zgXIuUcNOmyT74/s0mvSq2pw1YEAnQ0qDEijFe0fj8liWrsr
Fg8BO/MuviuAlXQNVC5Ods73NZDeLM0l3Dk5uw74B6uFecSEI9OkNfKUslaB
Te+xWgSJ9ynIZZCDAAYNpWuP2Xk6KxgGPde1QyWLQk3lb9W3HjCEkJ+Q0DRC
21LIBkfNjC+04IyJi3SN/F4KF2TiaTQMardqTTZZvbv+iJdWL8c7yeIEVIPu
DrdET/LCsNAgG2jkF/FzCjrNv/X4gJuYXx+fXi2Hwuom0sSW9CqHhmu+CK2U
V0vKgk0ga2MOgvrKJ7SnOsJwRjA8JClo44KIaPHKQ+KwW+2BcH48B6a4Fb5W
LCdU5f9YvNtnVniRIKEZsNgpPybIJLVkMRrntjVqb0n8/58iVq9gpTujj7Y9
Oa/ys+KCUqkNFiRjHQeOTxj2JRxub4l67yE1QgJ4aAJCdrFLTiM+F//dxisc
EsFSSTEEPm/5iDgiIka2t+TsC70r78qQj7BYnO8D/qJqmo9+lr13zYDHa+PS
tQ28Scrc/2lwJb3cwCMMqDzi395rF3vh7LnA3UtQy5K5COAPIwgHoyYrGo5T
tfrbqruPQCUCYhLGS/GXbskeUPx3afoO4RfiCCS3NiVqHX36vcfn3edU5JNQ
9GAAnZ8FkKUrh5MkZ1U2jiaG/Qz9pVaflqt92Wa5oAlwsDACIE17mxbqGhXx
dbEskPg3mSdsqPzm1vUfvbsdhngvWD6v1MK7xfLqxV8Q3wtCLvC0yR5vh5rR
bN94F4MQhPIYptPIhIh6oV/ueYAnTDdaW8NMqqqBD6BmiT4wORyoxCONtuui
UbePAeNdY/P5QynvsJ5mi9M1eYhQDvgJZsPLzW78ORx0DCLEPM5HvlOsTkco
mpO4ZsiDgHY3Ytl/IrYjc5xIJOfCmm7eiwGzQyIQ6Or+DfvglCnNg23yRtzz
B+XErzpgHp3v7A3NtAJw84vJ+fyKop5uaU/M2bqOfSwSETpttgACsmnKx/kN
QNqU6H7T4zJ+PCgleOJ5FvkdYcCbR0HuTlMmDFs7OvgudWpilc8IxBKUDpFP
kAO+Ab/f0m4vtmx9/px0JnkITfl+Fl8yjdOfONh7r7YmbM6dUMdeMYikLQCD
jvvEtHeVrJk0Zbjc/c48mR/a/W/9wDQSWHwjpJjhRx2hzq+b7RCBuu3k1G37
LkM4eZY/7HJFTjHS4zZjsuYi//akiCFyKpDGEjeYJZl661sp7Me6phrow4sj
5Y+Od5n8Xzuwo5W8UXpusneK47NvXeXTL+LgKPA9pKn/kMLBjrX5Jehy5OdT
LJttXimzcqUpatwFwDZaL/Ip454HRrsSEw/1RE/jXu4PjdMS3gmiBKWM1DA1
MYtfCCXS5wRsYQTwAeA1Pt75pkjRzB0p9TeaYzPXaSd7elzRbNeng/ev4I3A
XcggugdSz+5CF5Drqh4uBbt7e0ywq+NQscOL/X1Awr/3+x5QzO64jR8ryPwc
TGwQ+pRoAnYqTAOsseTngdgNq2/tgDe+2P9H3aYDWl1rB79AbW0SBLNNkxrR
5e89qoQVi7vi61FoI4Vw0uNY042o8d14a3C6N4t/XOM+LaGDby2KzsQqM1bd
XGyh+ZzHpvwv461iIXk4a3ySzxnXfvrGp3EexKCwjqQeiHBmh2AfQuYk2U4B
Ubua+n3Zbl7DaSmiM9x/AdO+HeuciayAHwZfz29F6z2bBIwur5aGeSYnDxGQ
LZPmKE0L1iIdZc70iAXAg9HR2Uncn5SB7QRJraG39uIQiKSraXyXNbuMH3uF
TlIbn4oxB91bFlKKnFTA3vPcGZ+UPY6DFAeW1jluK019yHwO+C81Y024aAt6
hxcRBGnRDvTmfH6+CSuoBLxrQKjGu1rJyQ8Cx53psxvEFXQHWGoPT4ARWh03
0pF9OoF4H0PmMgrbAKjwqARChl+wPEWq75tYaKXgdCwggDf277WwRXf87XCw
pfIpOubBw3Lwn+qFPrhUgTCDgDLcOz/F6wWo+i2h87dFzZeQPalgyY8hkoqc
HS7IBLljQEBHMdhO06Ykn3AquuKwQ0dhiYSpsf0YagrLS+zzl/J/XqnS7zxu
6VzkwPl1AZ0zceIJ+lMrMBsqovdeY7jwMl20CsBPh8rozdFcZGxQcv7reGtr
TIss/q7+6WJkidZZLuCeNuF7tIkEqFVpDWGT8H6N7L9JxYeW7t0rIyIlTbcm
/3bmm1//XtqBC+E6GsskhVjfJ9yi8gjkaIlOr/+As+YfKTn6jlfOb4QMY7ao
3Kcj6uYGlvZZPzVgCc1m0nO+r9F8vT/zeVPm7EQxjYvPiznVaDyCgdqCb9XJ
Z/AYHFSzaYCAvVc8U0n9xCw1xugWqQzks4ieW4oMN/J5uvYiYxX63uGgfuDw
/M4SZOW+6Zmj/Dji6NhTP4Tb03WEcDsR5c5ZPiLX8JMCWThHgOAwPRwAYQu9
OKuGDSegcCTYDE8ufTBbD1PwyjpyPlftSmKe++A9PEwxbgrTmflijhRvY0X2
A33LatrODszV87bao91wyytpHUHWPRKS9wsWkwF8z5XV+DYFwJumZdAjYzle
+1JjNY4eD5LtMV+LavzB9aEfJ7+WR75lE7yy0G96A+Ix9eHRUpv1ZECEX8mM
aX+LFTaTCVIlZ4P59NpfrxoIhlvwGTY1YJN+S/F5irVRs4EwPY0USSI28F9n
tAGDcZcJA8Je4H+Vhv4U9nvMyqaWWODXlBqLCPf+PyS8ZTWz+D+4MIhySB6r
sDm5cK711KsifqO1TOOqE1NTtb5RcWUsleAwd9nGohPWsP5MBtuXFVXA6/Ka
yrygsNM2O8N7InX/RNM4RDaJiPQFGGuJ5ribVuMWrWL+v9ioqr4AYVGQ6Zd2
l9WpWV3azbZHeyyOsR17kcdbztC8oDPtvJFMWBtgBkLd3CewbE9tjsbHosku
F53KRr56TDALki7xj3cQ7SNv1zlcDj088ythCFGB4xvRaO9mzN3OjxvAaASF
EOINhOO8pEQZzoiXOZKYMl+TYo3VgMf3RQ+ldiCu/xHEGL7D9Yk5rPkqUTqN
bui1Oa7kaxo6gFKlZ13e7uPvo+HfYuo4XiutPdSy1b9aNR0dzfuaImou68oG
qkAiAFOALAGjz87Q8j5YCzQ+IcWm0qRvS9obOuj/Ep3zUHkbtbub/rrz8mRI
E+TxdBy262QT6WgD3fY2L/uu8uXyPeuj4sADdyVfgyff2lammZvloqi4QqoQ
/yyNoHRF+U4bl1qAcBryh1VxQlpqE025oB2CxnMBW4HVP2Yn4KQNPIraRgvt
TLA69BxMP+1Vr1jdy5JKqH5iqZmesJGkmOga1m8WJHU8GHY+HsuXU2xHA2XV
wRUIEUNa4G5Ln1SaK+3HVWaL0hHX2Tj57cEkcizt0CmMm4sHd2HmsWPOsa2U
ngkOq6mbXeJeRBtZz32eublYAOs84msiAvRBxNnnqd46EwnIQZkfIR68RuF6
Cktos8PNCIrb2sijaOUJsN8aTwZn1KJ/+qpB9L7i4DDMDYKPiYIRlPEIG+Vy
i4qaMXWWMiPWjDgxF3pedyyGUsRFkYsFH54dK0+N2hgWGRUB4jZ47QPnCUEF
5NWmOvccJiniSAqfMY9RNwokdT8v1WSHkN88lwedgvs30JQNn0IIp3HAbwYY
Vbnx0W1LCljSDYWEWnlzKKojTq0sIOyzu5Q8Tj+oMpQELKuFqs12TVVeEsy3
HR4U1I4OYsSch/jwY1S30Qp0dqRJLk501MwSHmE6G6zFFBYcCyieXtVEFcoX
EPQLohJiSB5ELvIj9VCaH4WyOWzpTM4A+Hbme12efWCtK1Ehd+cju8/QFVAb
R90e/5G9j901rLFJ4laWMcQkStHPBhhwKGnNxnrIJK2R1wdniyuML/A0NK1S
l0XRviGQj8MhvJOoIfM1s5mqJ3jtXX8BTt1p1FwYIswTC+dJrABaXr3QnVwR
rmU/tDGUjTql9krovhVkv71DIdJHv+zqOZegJyjDctX//QMD0C4kUWfo0ydo
MuImA7ibfgfAP74yBJhSiva0AuE/M0uELA3Z7BRBRgYaE3+IyMNmEuoiP7IJ
iaTTFCQWV6t8myZH2FIfeVd7k5POiHtOB4cRHJCVFPppw/oNhNAXvK1CQu68
sgrldJtxdp0DwpckQYHKg6rSjH1FufN8HY+hoct2DmljxbqFSjWveaoF6bY7
2pRjzjGwzkbas25EoNEe93EF1PKwxVL50IHeEFtTpxqqlI/MvIJncb+TDEld
CDf9ATsbn2BlYc39hxPSQT8ZB5JLUFTrUBWvKPVVHTKhftUK77NZ7YOSVxcS
GWZoXpCS4yl2Mv9nYdcQiouW+2tJPheeh3kNHbfcNST7/DGqeDGalc55TRrr
BPfO66uPeHGWgz1/i0ZSGIe8l6S+cOq1GZgXhksoGJxAQGGDkW+T5QzX9vg5
l9HeZw5f6TD3S1fTflJgh78UYwtYe/b1ElJrDuQxpxY1oPkufz8p5dOEVPkZ
V6AarAJ2BMFpk3NcavjRrxCttpPEB92i7w2sWvBnUDaREEscCKgzRUvjZwig
QHMa6g3D0QvDTaPZKotJzrofgK+LE682Maq8Zfl7Bvv7HxthtoIeYabM0QWh
ZZltA22mhwsaWFuQmHT7h54EYfvLblZu9W1gKm7GHKcP55RrmORa9G1nR8OM
Nf93x39qj/bmSqRlk8PCSQtCtWTdDZakKPkv7uo+aj4zUkJygu1C8e3rijGI
OAyLK6I0fY62uF0tveVQHkrSyOYyO3tawFeLJs6DmqFwjagaJDNYUSSuHi2Y
W5v13LpFxn+uv4kGOe5SdKx+ysxleQl8EvhJ2acV1Wrg4EUjCGpFUlKXJPkh
KjUuJ1KsFtA1tVOJ0n8f2kkDfs3Zf81A+BesA+Tdp/DUB4IPZThbKGUmQv6B
ORC7AQBYUkphpSEmzbrELPDtgzNK2oCLn/fpTUNvKIUi8V0UtTnVro9Sx1Mf
U5jrBXpD8es8TyxusSh1m7c7sHgvjVEcOuvSLiAlLQnoiGP2XLOQpOxk6U8D
ydU67HOzA+JWOjiQFWwhCMnRYXFPKMpewWZAEJl8lRH9MKGxEQv2OtuATD/8
Xkx36483EQat/2qZDfJObrOPRNtkwzBgS5RhCad7xFPAyGgcHSZVHJKIi26A
K1i/WN4YXmwfr7wFSNaK8gxjjlEjLS3aT9VT/nCPv5UEyn5hfsrPZ6nWqcdg
BQwAQHdD9kNpT22WIz5plGe9RW8V2FVmkLCtwKPqXB1cURz17YMPVO/pw8kw
WdfKMpaUlh8bqnM1PCkKremLc3DTRhFJHWGYIm6dSREAdPPrO5DqspDqrYaE
M3YChP9vxSyzENK+jK182JQjHMLAGT1DTU/0krD0IA+e1EdiklBba1cKRj9t
ftIpdBzVNoM+e3BO39y4RLemK1OBWrGwvcNk+fThbvPfnak9nU4D1wLpGXTM
DaSqzVgAuR1rCSclcv1YojPER8ExmCzMYqPcQmW+Fp/ZQqbaT4QxRZx865h7
m0OLzz9MA6HriqpMEAya65eR8ES18oOu3ioACvws/Z1nINsCIDDqx811Javi
pe4kyk0FOJnjW2sGawBNXdI7PeiadSz/sij5lYpdaWMq5xnmdRAB8p4rjNy1
9RGVxVgUHUbF4025UVNDZx1dg0DJ9qWQ923NHUnn8DjVc4sUnZg8+WOhBmEh
nDaMdxdqMtOTufBAJV3aVNsRZ6QDv9pKtE2DuWvcAwiQNeJ1iqUm1Lf+epDx
u7OAWJAgz5YRBr7j//hF5YmrWStyWD07EXoZMP/VdfofhWNi3yl8qx2BFVp7
7qWaFqLEy3nwmuOLFlPWx429UaBGbPB1c9cKXHFBxzoXruSLTQqDETbpgRys
TKW2potxHTVXa4Lvlbr3nKX/hGqDVlSAuMWlpTgpZCHO+PAS2gYowm1L55Xi
qGw0ZYU9jIg2Uk9Kl+IS3mB+fv0eJQk+V8IH124GEsF2b3Pm+yXKyzX8yJ8C
9st/G+MDpyztBtzvMmJNg1U2h+ENli+6Ea41UQ2aea3fix6/Gc3cWdBwJuIa
udtuX7OhCNieD9o6GRy6CiNtFsq01b5udpZGJh0Z9UpXZUu7/muuQnc7P3G9
qW/1A2Nph2wOT1lP6k+4bVtKTCK/t0qhrkhiY5NJSScSXVJ1U9jyVrrPga6R
/BUm13OE1PbyYCuMu4Ni1YZ0dntJ+OmNYX2smKJSpwx/oxWjN3a0uo9UG2OX
CoQJq2Bh4pyp/4MoSj4FFCvuzdW2IYPA1wfrfNu6YywogO+KZSZUFdOMhWjc
wMHeTZcj5mF+KdM96Il4fZhRLtiAedg0t6acXuutsb5epw6eQfcR/p/6ZsxY
0ZpKOwbp4LF+vgj7x+Bt3lzxKX09CuwZmfO4OrF6y7L5SkXN/t7PFOLlaFOq
X2AQSmfww2uQgMXiTpmScPP5ID1QobBASzzM0zMH/UHvuW4+fNUbq7fcTXXm
/bSEG8bILEhzMhYqv52B9+eV3UOOpezMvDpopMq1Bfx7zy0Zm64g211bLkgE
q+oVcZTMFgskgaGn9vKMTLSD2BODryRTzCATYEOT/supgmMD14SIbkQoolBw
OkDVURiHT7RWCJbT8BaybnZtxnNAi8xR0E/eReoOrQsMIvJ4yEq+AM5hbfjU
x/lvRRzmfNLJ6odrI5CUmypbLZMRE/o0Wlo52HM5y4BuYsbbH++2H2g5tGq8
MeNNm03hhHM+FrylzePMfsOMEMZXydsJEoTEsJ99gyoH3sJVxNT4HJ4ES1q1
2Fy/rwlY0FO4aNqaXljqxmY/lrM8CZ7dTqvaqGL87IxPY8WA6T5M95vzpAr3
cp2Z01F4JJ019kOZvYv8h0O26ku3mTzkUu1nxO185qXEX7+tDNWzcYvMBBgD
QvYUu34Tsakr/GbiTgGztawiENW3uV+wD0Q6tWJYw8Am8gHGEDNDnx6eSWTH
+aRTSeKAdxSJk9t8wSbJPnTXTsIhZ8l7HNTCu7czChomVToCv6bIaU9Ul5Fp
EtrTmRoEEYztm16IJhxtUQgM/CTtYiEwMLH/YN5oiZEi16YdjoFy1bOEpqz2
eea76vM4CfhAeWjkYtEdgxycXq38bpi1HvQDlLq+KBE7rue4yEo/QHvroUsg
QhC4uIyF9+F0TngbAn/FfsTzlQcSwbKOzd7bEmf5wSMVSchldM/M3Li7kAjn
gfTgx6YPtKJuWGV/G/Y2EvUiHDcbfNxSLMSRfjARVhdeWFFwbttLko0fQf8y
YzRZQ8eTr6z926Un8vdpywo3LZ5M9NRrBU9psmG9L6g7kFHrZefi1siuCVJi
Z1ptsWNOwRctklS57eTJfBIIPdMPhvyx0UjDg1tvHvbpNdoA+T9Ly1+cNUsZ
JeNb+0gV+kamWMXHEkW5/vG3dfVscjLOevv7g4GMdlpiA2SVjV9GluwsOOdS
nXkKjoWywKSB6if0IgbG5r+ioxG9V3Ge48zxTuk/ys3+79pWOcf/GdTv2Nod
M90HEOBuRyAJGL7dM0bx3hZUMFnz16LHkTQXjlOwnammLvCugwcwj73BltxV
+B4WH2wrsaahhKm0DKC+qRmSSocTLeVX+OQkaR/NrrfGMtyOWamj4bMLFiNZ
vT7jop1PXLigxqXlTErZ3DGTnrw/1obd49wI8M0FRTYp3WmElWsYuQtLpjP2
nhD/ouHXkSN1sTjYXVw1N05pv9CF9zcj8kfGPMsT2WELVo4YodrGUnhpC2aP
DmjE7Yx2tdbFiBgxyIXqGRbpGQyz3aQWngkvitJZjponLnIhnwPgiavg769+
0JmldL9E4EArBViyBoWnBZtawGd86yNA5Na4kuqv3x77aOK3RZNn5qD+wLVI
QTQoKOmuR4lk6b99FZopVMIBodIL9J8EWin8quHFwLOHeboSiYKbL0O+OyPv
aP0LSWYS0trShqBG6kECS5UD9qQ4hPvIAsf1AyBcqCXXxDBX7pYgpT4Dylaf
mUNzYL+MpKCt7chARb6nBj33af391bBfiBnjcwzhuVrX2/ZDkoo6DvWnTLDL
eSN10TeOJ+IBLtsJ3/3T0InkfJIM1eCqjI/uYCllIoQP37r045TCUgJ/kClB
PWQIsgTLSaRZYvus4iseT8X4iJawkRb1qdotSxFlFHCPRSAgqFvuZHraM8lR
12aw2syctsOZw5al6YrFW5pRe8gj+RroijLV6nSGow5TFcO6R3MSXWXM09IG
06nBKLKdRo3wY1MWh+G2y5bI5IVZbQ2HkwCsSA6UKjKXCunaF4uMwrzrzkIH
l4kx8WSmCLDzSPg/HFAKKvyi8d9i+J5PZdIvHYoK8w4nVIm9XR836kr7bSVC
4Va3L/x8fgnkkzl7mrJ2M06QfyXQIpJ+qVSzDl+ljpTag2VHw4sJxPgsgJZ5
YK4L9Qhd1wOgz7McbrZFaSJg/6q9pwM63cwv2eNjeXsuVHrzGgHHEuSjTtBr
Yfg/ZCENUZkdojqpkn/yPp2q184SJhnJaZai2DRbFV4gREFtMk8PCrN9afPo
tlStSpk9xquxfg7Rh1VDHtFbxhhdJpDJOfx4Pey96BPcY6TTRGjkCHi9Moek
MD0y3rcv8pHjOeWYcM2zqlnFxLgL/ov/NchSyl2+u+jWmbnco52loWsOkubB
HdRFS30li8v4E233p8eWXyjVDlYccnWn7oZ13J2cV/XACNq8SieUZtCvV5td
JWdAqXVP4bV0d//lffRE9kV+1ymT0QPGeOH049rrTpzwmiBhOtQcb/WOKvzh
bIWJRK6bwm0YFlVTPidxU+/IgYOBL9v1uK+8IGi5FxGJito3tk9QP5I7Biiq
QYtEIiX96f6QxMlxuc+U5zKzPswWPAX0B9jLKABYDIr9qZADPcS304weY70s
JFe8MlPu/gsvWvcgdKu3Gsl9SPrUfewhL5aQx/5QQhBpeVcrgV8Db6W6Fmhv
9EWRLke23DQ2VGjYKuNWtijjbUt7tUCfK57lWZ8jsEZT2C0z9wrofuEzZVEX
hZwcAxk2/s1fbx9Df3O7jnsJtkleMq2Bx/+OV10jc+nhlMw55qc6er3LDa/2
CMmPQKTqm5FTSUNKSUgxwtGQqYwQdySsJp3EO8BcBkQ9eh5XhltG0rzJHzL0
Pv0PFc3+/ruN3jb55W+hcNvAeNKTN6rm5cvXu8qujG/0iNR9Q+ZSORKaQ/hT
unw1Zvzm+fRUqiN9309f7k16a+HkaSzdHryjvym5je3gb6UpKgyjCyoNl0vU
d4F+dJqbeJbqz3GXrxBMqTCaFcjoTuBmDjZUisqc4BH5/2OzIpe+25F/2rNo
C2nvJnlgHhfwkE0qYO9W/wCzLcNnaHr+faaWVIG4Pv4NmfNBrypu8Q4wNjMj
6WWCtwhGG5WcZR7sOhuCN9Hcu85Eun13X+xFfgaR1GTuS+uSCiI9faHCIW7p
0BvH68EhAn9Fe7oi5EpUwoKlPGS9FS13pp27rR6PdORH6EZFc67mcaBNni6Z
KYyGpzuYcWUTR0S+PXCw/49RNv/bbR2fnZkR2a+SaqA2LI6alFkFU22CaTQ4
SFAkhpeQu+s1UJVRCMhrIxvtkIbYSedA9rEYea9fVumJxMgkZWMoZum5W1eb
b4tfJi+pyeN/GaFIHMlx7KDeiimUKajfJnlyMMTry7weQJLXUwY5Y/gbFAfn
+BhZNU6YBSNZ1dzhzpTUpljFoYo5/8HgpReWzrcgDVC0beXmzu4zkF6nHxRZ
fhcqFF37HbEu1rwUNxiEFJS82VaGH4KsiZ/tBSLvOzx4Hkz5v3VznwH2QVNd
L2bfV3J6BsIC9JxcesF7AXYGZrnueuVw4fbjjGJsP/7xMdXMlXGemoQPj081
BH0D2nEOmi0MRH7mUqm06vTdo6mS/ycS5ZHLVgg/f3Tt6O8HSEydoIeJTZGW
0PjlR/2s0dckkHoq/XC2jlK6/uYaFzXIrf9pbArtZ4dDEXFTih4qFbK7LunL
wA8Op8tI/J/A7I0gCDWOOrwcfh1O/iKojje3JNXgoJgnlMVnFJLV+mXvFpHL
o4a+bWnfSfZgNRhb0HmdQ2diIH7ARXPEqFesWcHdVX0ECv0jivF+0ujYrwI2
dTRtLfQ9g5ShLsF2YO8mxxRtAoA9EaDrbqjmZ3ZEGiulVV3yq1Auk6HxCwG7
EEcgWpVZ9V+PIp3Ce8Xdau/JcmaFXMZpZnalrKHvWQ6OFjKFicKaQUGuQyCq
XUuLSBL7Odb7YZOkXVMLIWxob7jzBoywlZFW6Q2OEgb4biWKioVy2uD9xxTv
0TsrzSlU5H8EZ+xA5VPR0EwVlZT8mQnyOo10psu421sCy62S8jYu/0yEtWY0
NwGr3UJge34T9i/QjPoqI1PRG5Y8p7PEJqjKU2/XnHgGNyrNPJVtuDtqFgQU
Knsjym/AdZq84yi+x7wztlTRvJ1cCYpoudb4l1LhLxy11lhpKMkVpppLJee3
IqEYy8jikZJqQhYNJ6PzOgEjR8yRUCfO5OJg7L+SOPim8OC0m1foUOVS3Cn0
jxnHg+8K6dhlSPQT4BPtCWaOa/nHRNwaAZbEgE1Js/nRbwAAxwSJUDEkq6p9
bWD2/VXXF2fnacijI0OcBXv6e49z+htBg5LZgZdtBhuwMndaLbPJE3rVEdHS
hBEMFHghC0PghMHweVGvzxUo4IqfattwsvE5H0YU86RDMMwkAFZN22vdUHRD
DvrYL7zmrxPSRg9YCR6gqBgcgNJiyJUS2+UiV4hO9sTOA+e8z2kLY/6Q2p4c
clyJa3cDXlud/zPBzmz8+bdEVPNQQtiUlM3PeKHy3812pJUuUQlhvo3/+O1r
xK8PLLNsXucZXV1mLBmpJqdiHdtKmUiXdPp5qH0tBkWnFH4k9S2E9FEbTOsB
gQJclhGETRTNtK0JEwRld10fn2xfcxLMnFzrKvq/c2ckkDRfv2DQALCSR+DQ
uQG5P6V1AkyMtkhfb5kfhRC4nAD73BaHulMbk5f/A0JBAUdutCjtlQ9I/8yD
d9RgxJn4nNQYCt8eyYPkXtuQi4RyXwlwyPYoxShP74/nPMdchW2pvdlPsyHN
tTAoelnHrik9MoEj91IXaHacEb4se6axTqD1EfsjPj+3+oF0ZDe7obcCc0fm
W/fFEemFvEUlSWLG3pqaIGdAoI+IfK60bKSBXSKp5xGb+ph8gmhh13fqWaRs
KM8WxU9BnyD0ob9XPNyc/wp7FSnjhii6PSBSXSFN/qAcsa+kUR9HEq9KnzAH
mdzt8byPSu5kasmmo8Kw3aotNg9qJ+RTme7Gu+TPVEL8chdLCyFtoy4GV9NA
8xXm0fHQiWnKcoolKZ5UMBSJQ73aKRKueRPiONNXV/vlVNGCQO2doCsfDcCt
vhfYPALbQDaePJpgJO6EWjlLuV/pEhD5EV4l4sx5oyPNfCI0aktAJNSVG/XD
CBjHNvrVJxUESPiJjq4NcUbOiFRiMTZToNAu2bAjJtXxfnhNxJREX0byEUel
yi+lpti54TMH4D//QZwDdpt7HNdGXIwSQ60St5SPIf5hM6DXCE3M0JY4uVTO
CtwgfX1skd3lbjT8i/aUv8m5gL9LGJnkoakWg1g0U4QfRsoJEbK5bOeywPPj
/2bEXrOnZlMcgDstKzStIhN9vCiQW2V3iSqrX0bJg/QnVWWlizI8cjHriTe3
uNAkijiwTmx7h9E5W9WEl2IkKkRqXe3Pf2VguXX5nuQyD15zaRHdHdE3ujfp
SYBnE+9P5DnyuSZLbNLyb2p0ldwTC6WVtonkMRAkudc0zRLjxQZQQMUBBzgo
5UMkcVLhqEsWNbKS0D6vMxzOpabn/6ZdrRgrUX/3jnWIbKtUs4kONKq2xo4Y
48MIVu7vlX+341U5fPsmaQ17cuT4ZdDXUWoJfhVmiHlgtMLaDDDYeFBipChA
/bwXp/aBbxGBG7LO5nzEozRGDLUvvlIT9/d/Sn2zNplEGGqNSzffjOmziVAd
PjAjDKNWrtls8BHAnGoCSMDqv6GC5tv56VBk+QwOv63hCxsyNqGkGNzM75d6
MGE+OZI+HpYGQHNbm1W8NCvkPGLIA8R2lgiJB4ZRjQwwQEFIWG5Ysk7n/CX1
/1JQZX11QnFDfU+g5rSSvUssIDKlZNvxgKVtGrJPW9gFoAwzRwxZjHwaP8Wx
yon0BBbJflIRGck/ztZg+SxO4uSF95gnmvORE+t+OISD6HLACgsqh+etuHOd
y8fUwTAOGinpnV6FnxymDKyetw6XYFTTMMGWO/zd+Kp3im+qLiHwnfcw0vDl
xUEYfbk5yM9x2vcI04xpYK6iSWhaiO7KGO41gebJ+Ry7a7sMd1Be73XSlCFF
eDiBzFfISau9aURPbpnMaue8koGv1cxoeDYZaTsGw/Sy/puInE+GZCBkP3wP
btHEaiHCz+oKA+0mLS8DnwOMs1BhlVADcAFrF0HTDmNnoDWrHzT98WB9pUJn
14oJlNWTHtPRlCJuZC7v6LTdD1xgU4f0l/2Wxa2xNJpz6N1/YDU71jNmP4QB
B+jWtxXTPT79/YGqSWKwqVoCfAyyoD7Ep8x94KUoAVLWOAiaYXAvIat/WOy6
TYORgFEt2PMMi6n7uAgf7v3BB9WOcxiWdSYwAUEZfT3kz1fPxLSjjjZUlVBE
OVAxFjpgeYHRASXKkefzUgv637k8lOSVCigo/JjyvmADtR3yh7tL+eO53hj9
nlzS1lttiTutHe/rPPTPmETi7kShQ8R49lHdgKfPF/1jmn4vZgjwXAv0tZBR
i4S64H9aXbInp7/pJTO8kFlhLNGNh9Fra/waoAWI1iiXdu5cgx74G2Gf5aGd
e5OJjg1owNt99o+eST7uUpyQrMrClZgJ0L+6TiapSf/HgIHn55hM//5E4yKR
OohBZmHODRsVocrKsUL2Ja2tCeuIJcCH3woekJx2hSKArlsquxn9pSvZuomM
ZXJlOa3v4d8EpixaWMAVdDdWkpUmb+vWY6P2jinw7GUut5SocMntWelOwW5Q
IdyjnSTfOQsviw3/9gc6zhA6Ncst1674tCuGW1FdfC1CYEJm6x6hIWUFzS+a
0k/16zH4WhC0Mp9XMctb4zAOPgHeWiJetD/2Kzd9jExRb9rrIIYoMP7gxGYA
D+r4YLt6nHLY87wbw2ay1uKU7syr1ps275HVSBTsYQs9MioNO4NqQH31bm3y
nObccnS//HqWzqVUvYTfb20smyI+GjapdaKandqc3M5NU10v31M+r4JGdw8j
+6xewFuU8VdjxgK9znDO+4GFnVJOSvuIk32RfwFDofcr1keCTI433Ogu5Xfj
8fsw0i+MpmHkCcfrNR0MuP4qdgx8Aevhe7EjK9AC1nIi7HhPNqms6t2jToc6
7LDey26f14YVNL9A/+Rp6C5fH57GygGaJKGFK4HK0uOI0NRKqYA1fBvw//vB
OdNeDuaeHLUSrHPsjC1bWxIuAzh++aybpz8ofMF/9eJJJF5mT94k4INfnkTa
9sINKk2zPc2sG1suUuU2kT7TgPCQ7YgsYqscvhWsGV+l7W7qWSR+6gnlY4ra
Pzhnql5ADNkHJfk0yhWPV5jpBBocuOT7kzTcs7BuP2DhVLFqs7xE3rtFpJ1P
Vc31T2xpYx7i3O9996t7Wzmo0r3M8RXcp+nVYBpoRw6muwseo0BCau3RTc+N
SGFEdPE70N1zUnVrmUFNqnmOzso9hlItTyBqK+Z2XDSQT7ZiUT2JZfDZx6ea
McaBGTgh477ciKhFSbYhgYB3ADads9iZ1CMaxMMWtf2QDNxpjIK8Rpn0V1Gj
zudk+/26ZcstVeDOQaOOwlp2LBpstKYiZCTnOBxLU2HhFep2FSwpwgaoiGxJ
sBOriO0V2dz66YPiNtnUEAhXgfMOlqIGlgDXGRsVtXImIVJvgAsVBiQqq5oL
qiaz3fZkTp85zPXB+WDrRu7FUEiproUX6vcQNiWkpv5kmXmu/G/x33I6eYm7
Q99RgoHCG5O8m+d3ia8FTqKYsXgOYeKsIrtTMPNKT6xQm5IE+oSsn2Tb8Pdm
UjxBu+VlWwQwevQjHpDy3cP4DJj1b0/+BLHeksUzZG/EehI1ChxY4vCC01ay
aHuD2SSTPgavlBfWszdPK347jHJpWFG1eE2VGv4nKrUJ4sfPZKgJMffecGAP
NxAorj246JKK9vCDouu8PEnBHu8mNpoJNAJPH6rG6TCM8ThCVKvO9b4ErsAa
CW4eCuwss9UVONGV9AkgVhDtkGHPdE9iiXK3sFMYRW5g64z3fVk8KWxD6WTW
vHT76iSdnd49X5QFfr/+EioDe7TWHLqswshA3yuGcskk9/uZwIRTOiGozENj
RLT3zGVDAbV57H3LyNhO26blmh7jE8EmJ1ioZJuFOu/g0PYI/fhpuSgidCRR
N0LjMhc3X+4T2zG+0libfTm8Ca4ipiJnKreyNQLnbO7I29VxzgYKC4KlrFTb
bRdFMJAAdxdrI08sGJyL/YnbwsmQvpbm4Z7qYLhXGWq8frpbgIEPYB6SXZ6x
uc8SX4iD0CAs/qgL3dI9C6E8TQLO/UAs/bpWFANqkffCy4qawwGaACj3mjWR
x3qQ5DRfHMbcotG+x0hhp05d29t6CJJUM3HCViakjlPSxYAWqquZKnrHwVk4
DO7vfhp6Uc8+9jnCAVWTfUAMhAEl4dGpFasXj6gdilc5NQDfsIbPyNFaWaU0
VfsPV7UOKyi+gKjQo6E+iS1TcfyV+y0MXQ250lQYFyEsaKdtk+wraO31Ea+6
Gc8Z7JzDM+l1kkUXddnWRWU7jDi0giwkxOVJiGz+1XmymwwfeRcUCkFld/EC
KG/TSRbGGP4mjlK4NogvsnQglhL3jxgimWjsOt+rh6aDTYvbvgD5dDJiPhyF
V1lUtK3RTy/bRcpjGJuEEPcd5uuyVZqGrT4XahUR4TSeRMqLg3mnKkycGgjG
IFTbVfGSzqNStyq5f779vkVoR6EaIYbTQN6NUJMOKecmuL1N8gwd+J+BnocJ
h6tTnbKDLw7NVEccmDoHVxj2j9Oak7XeiOV13vVWZBZgWGniuCTGkIFjgVoD
KXEqNcVuOdYvobkcIwN4Z6++K6x2mpWJIKY6eurk5mlh5D2rblL+qfl10rb8
pfc1Vxp0/gYXS7pHLXztyj94oD3+k3BoyNCAwTMJPUB3Nb8lcd6ZYTHQ+kra
YhYWv5fBBn87IhQGW2xj0K//xB41fD2TM48qE9kjlIHa1K3OcgkKAhL9xlhE
T+yBz9UAVTMafLy+k2mjjBBUCLjmvTtxtS9MxEJZlbdKmJzkFWtVJi9tme4N
Hspr7ms5g8PCC+/mZlByU4zICbiHilUGw8yPR8xVdXKJQwBOjJNRzxNMYhnS
71uWYyAAuiJDBv0OacXm/cgE0aF8qG2OleQD5LGzNCSkeEJeNXVilYqJFtzp
vbQ4Q4VxggCtf/j0DaJPwv1DYMMvczFmSz+6DqNqnjVh20hCTwnU07ZAF4zX
9R966pHwxrxbPgAtt+OWAFbHx+qKtst9KQeZ2bzBfB8oo6PINx9EqeFwqSRK
X7XVgzuKI38sqBrmmaoMNFv9EnRWgPmRhR3CL+PR2guwlZjObGlsF8ApRsxy
ZAXmXnxK6FV0poLehSq+8Hjje/vg/7d8BpJeQZAWDxg731HfWQpb0yLeVL6T
H+APR+gVH2OsTj57fk+1hI06zMDNG5EUoBCV0bqjUcMWijS2oCiUgqqeXxvG
S3O4eYdeBghDXVd1S/l6/LvUAtS9200N/eQSRQ9E1eEGQeIcUMyQUqu9tSGd
ui4z/P8MtANroyQw692a5Vo4wH9LGVJnummzvzvw1IeFOxEI5/9HvEN3uevj
JiEGJRriKzgcet+sy2Fe58uuql3tNW2hs/egdZxbcU0j2SStfrMGTAcNsk1D
WXuyPjJrl5DctGpquBrzEXSiQ172eFzaXl9Bl3GXv2B+HiK4oVZoFVf7mlwh
gOnD45s0e++8bmSPf+0+o3+f5fjm6KtG8v8c1SLsOANnH4CjhU0ZTw41Abaf
gnUw7mzkX8vXBJvWlVu2vxz95QJP+Bn1Pj3zhbMfgL7w3Jycx2oR3q4vcWDr
mBXYvB+jwFi9O2eHbnzVF2ggd1CEV2b8utIm86I0TSDErd73eg1t1BIPtisb
9HQ5cKpAh49iz+l+OrLgKCYC5+NC/yl2VjwQZbDVK7UXU103rxiIAsavxT/k
ugLJm/G1NGMioMb6nnv3Udu2TR0dbbdwrTbRmUzPrX8l5CL3KTwsD6w9aRxL
/M7NipfNtvmwV4oNSU1aevtwtF6cVPiCHRPac21ViCKyQ6Rfu+of7uzFGw15
+eywfo0CMXCSzDUE7w7EAJB4gLA3SzQn6vzU2ehgOumUl0vAej8vhBrS6rFq
1TXc06PNHGrvxcVKsO86rYoMq3a6QYrJJ1omUSk0Y2xCeGZpFwQVGiG6MpGc
uu0Sz7AbUgJ+TFNfeVaF2gDF2EI1rPpmYfHy7Fh9jcTERHQf+RKkuXSfogJK
KIoiWKyLnbKo3GXdJ2McElooK1oiuFbUrXH/P1NLKIWWSbIyl59dJjIPGvL0
hBOJxlC0wqAE+xEU+X4gQ9riB2xOB6koFHNW2xY10HNQK5Xp4+DUot/8zkT6
XeLq9gm98skiRXIMfqmZROgz+cB8PCpPeOuI/KmFv8WTxX94MZ272MM5w/i/
NBsZhjnhyOmO7LYH76KRQpfQFgxY12TFO7PpkUsUk3PwTxa9g1L/7cEGWJuz
zZugosAbObVUiU+jq7BAjKSXlUdMscqiflYdrEWtn0fBo1crWbPokUFpMb5J
QnypMgMRcP6bmfqkUK472Tl9q4ba40Dk/VZHhjavAE57+4fJfB6KPA3/r9Xa
Pn29niSS+MKVIwElMVjgb8sXFLEx3Zs70bVtpazxMZ+EjPz5wBySA3skglqk
oSMO4h15ZYQsRqpIygD3Cmu5v7hzUC5n4cbczBdjOsyHudZGOWexVsHMIjop
k4t9MAkInI8J6X3Aji9xj/EkVfik82U+cKb7Jxw7f7unh6wgJ4Ht89M6zjK8
Vx8jxP4hTsTprMzjtjhqVQUByZ7AjvU6g0CtOo2AEUuC0FHby8qDrwBr35oH
59L/+4nqdxy01eytzKtJXSWra44Q6z76d9HV5h9g7C/Pfii1vLqiNMpUxEL7
f59sdcUcKRqmUHnw+/dGo0W7sTaVc8v+bSmG+ukRGE1fZaHyDE5ZI3yIbD1F
+SA3eLDJhEdPQ/3nTVlqEH0BNT1fbT8zVyC5ufEl9ytghz0i35qdlbmSoyT7
NelFvfDIy9gaV36qplaaetN1raCZkVDFFbJpXhyjSdtzJ9KSThh4Uz0I6Lnc
deDW79vtWpW+qW13NKBb08X/ueYqNBoiO+azzXr5qnsq8QBsdS1fAv7rOfHe
czJuHXVQ+dnQdQievAAJzul/+YkLZ0dG7ZXoM4o+bXt3d7n74hzQoKJAKvOL
KZib4wexo6sG4aHaCxnYu5yYoDNiFAEI0qW+LmZCvGECky9/BLoB3NLc4Wz8
R+tTcNQjZXtj6lboPVL3IbOc146ue99WfJsFnn94zIvGPo4OWlEs7NAfaTye
9dr1OIYWOLKnCOc0vImdsXaUwFBjTQ8BzZCvzW/D9K0wBo+46eoH/eibvXr2
qiFGHCSMnNyYgpaxvL/fkn6ljO1nhlC/HEwq6vHNg2UskpDrDqC9DShS3CQ+
DUtymAq3Ag9gTQjhg0SstPLM8YP09lz3dXJ2qXYyKnmqq0tmd6eFSjfI9hBh
3LPWYknfCxVCzKoODBSxpmHk94dkkcQ+cOZyTjgO9Bemf2FLwDGLDadP6zhK
KpE2if6uD13T7lCeZV2yBVrMT1wVHbJtoDxM9wwxpekZ/IXoCkYFC0ER7xJ/
gMeCDmGTmNynC5o84h98HVseT5/cKM6MPt1RN+Do6Po+jrHYwEhFAAf5OPat
KvQmf/2+J2uXnUlUlbKet4gNZVeztu16TvXN6LXR4ln02H9fZR1R7rFqoaKv
YMTuwsrCtNmhAQNL7eaai2jwxqx7VOcZCFim+pTZsVAEZ4uyJKeYAPQl8SUm
CTfdXZinwmnxr/eAKR5HMCcidheefjMRV0jj034JldRlR1+8Vs0FLkDz4QC6
eo2mwRpyUBXUrTVkKliR/G+FymYiRw396ROMJNm7bB5cme/jlSYVukhA/xIp
BJhf6Wdc4pirIeUoKSLHq1f4SUfszFnymHAo2aRe0K6z/jHY0t0jYz50jJKd
MxvFSPEq2xuBJgzYdVpcKYvGhKwivyU8dccgYb1bdez+WLHH7rlLgdIVd15Y
8GKep4Sh6YpjB9cEqSAYsj1TzhdMwjRBH3djYC6Kehelo7qzM6GW3q6U6AmV
II+hzLumw4vVgobkzrOeTlPlmMjT6cSv6bzE5Rcqll2fU5VjkUEx9UdAEQmX
xMXOYjYsw4Zz5ervhaH7zM4k6pZvV2dKLATmCj8tUl1Fv6+QQf96ICM0rbIa
YNqEL/wswAffi8MwFL6AdbyNPhxQVGnO4IrgPAOssSjYDVMFftfStAzwsKhO
BvnwQIsxOTrYSTFXCznABaarSS+ZU5fIdXpG8dS5D97DMLPCd03ANZy44tyQ
3xKSTepAinfz1LXrB8TAhuB3BzoHEWM+fbs2vT+FbNGc4J/qr0hSsbFYx9BD
1z8NNv8jlH/dNlHZu/lWfW5BZ+i0CBqAgIwF2Zu9XPKxUe8u29uH5KIG+xzE
EQ9sDhJON70UF7rdmUUgopb35215aFy2LgOCuiM4VT3MQtR/lVEhXZHHExnp
CIHoMjq8/2jtCu+FYu8Cdjescdi3ewrJhXtNGfUPzkhpbmpPorcSuZ8DQB2Z
1iAhnZ2BVZwPLhl/0ipd9HXbCRhDtaia2Tt8bK6T9gObkbqUDGB0tfDH7wbn
c/zCEZ5DeQP9c1bEQt2+H3+8z/qQ7bhTwYVtUMmfDJanx26ryn9sB63fqu6N
NE7TMW4Dq16Ml1Oj6Q6pkHiUrLfQcPm8seOOPle54MVlQJwDIcwR2RGqP+rI
xIvN374oBwAd4dd+EfQoQ+Fl60i1tABKoHpqHwA6UEurxdAnOll7d0hS+bJL
XYBsEgV/awhpaO4OURPlYeu9D6O4lsx/tsl8Vjp9I3Kx5HcXFgB6jBFS8+7c
t0S7WubgV9To3Ipc1ycaOxF4TV+T0iLcpMkpXQHmrPLyZO/6AFow1xt8ryfz
eCHDxEpq6exgtw0qHXG12csLan9NTV4N5gO9Y2o6VTIaAkWJTjlzMXQ9CSZv
sBLri9NiVJ+3LlHxV6S+X1LEISo1oV08RX4O21YCtKJZOOMKbpaYQXHjczbn
eda86i48Jf05quC1nzp5u7YZ4JgvBJTJHgzD/d2BTAMt1zhgzbNOoJL2tOpp
yC5ysdzYonri8OOIfAF7lbcYBwiIYViDOUbbOh/cTYNZXVImbqyc+lKvBeIB
LBbm+T4jK7vUaZk1AO06sxz+VHRtsQtnlX2UM2XznNjSS0hH3ZtyYDWYz91r
s3D1Xoa/UI0ypoFoxkV+XppJuPXsKW1Xr0U0YV57wK1npUdgogQJdwZi7o+9
AwwOz0SotZ5VBSQIZqq6mAuIieD6un62xuK2PF86FvJ/k5VRyndWq65cqRLE
a9O+64gtLWTKin8JUzuzDs5M4OWPvWwEkfe18EmvR3L5ei00DBlGxJBD3l4P
n9VdArbd8W7HZoNmsYWyCXM5LzwcYW5ejPXzIqgZWrHVCpiXVC3s/wGSkkHD
3vxPqVvzKNZEMIO5UO0YNE5QUkHsHq3qFjLV1rPgws/wTZcOTvMiPCXL5yOd
Hti9W2t6Pn3QIjw4fQKqmfKCuRNb0+APdZndOXM5N/NtsVk8xHBNrRAY3DCc
HdWk+zcL2H+/OessLa+fo1s3C37sbd58dZQl3T7uuIiAAzKeZ8WO0EnbeeBD
TzQrRNrWOAmJAzVqdf22mDRNIZUGSZdr4fB0W7BRxQ8oV+tFHtciYURD/wVf
B/86HNTN6DXeG7PnuZGcTR72FvbHB7+1aMEItymOnaf+iRP/CYOMQmTGNzcW
LHUbaAOIhNbVbUdltzq2C84F+ycrcRqopjGSYI9IWNIJIj1CzijreTQQ/cRX
cBzlV8WHW+dyGiYQF9/ZmAT7mAm6nHqqgkIdvAiyh67EbHRysgMVkJVupbKT
LYIF37UabQRDGp85O920cdwSlRfbSVC1rSVA/EymJ8eYaFKY0aDpvHTdRvzD
/EAjD14gSq5cFmL3f/1NL+Raofh1vFm2kejU2FOVH7FNUuez4bQijskOlBWU
9K41S3SyU1SOtN6ImA+Z3uf/A9k3pBeg8PeKAw2QJzKfxTihBY7IXCOxWkJw
pecd+YQKKJlYMs+OFypLQPSyMq95Ywuavz6YNI5ZdKzp9KHyKPmV2O/zBfnG
/x315V67BjGs5f6zODfbnxNbMUHjyStQKjnHMBsY9nAUDO+8qLyLZ0Zs4xiZ
tTpWLsXU2i0WI+y7NYaGDcWgdA5anoDsvdE9bRVgLwKBj4fCrT38/410ZXFF
dQPYLcpdpwLl2KSLstC7d/bklXzi8pgfRgi7fXk5IBqbj5tDX1H+lIFLWOMZ
P8f2FOu23+oxOzozQsLzC9DQdp09L9LjYInHDqVgAxQQUlIbmbNAstxsDHPV
NHPqc4bUCcR6oGCjdDlz9NSmeiTy0c/S4LRLicKbm/qSieNk4lxVxfIOqvnl
SVymdGtpVi6a2X8K82HBqVEzKbYbsgJnrE8wtXVZl+wX37RblRlZbRaxZfK2
tEkjVLvi5SdjbrR60GbdzqYaRg0SDqHBzFhT65mAXJL0RdbabvLsME9MXJsL
mkPuHgUDEABkuj/8pywpyiWlkFYYFXVWsSMSoXB2UMWkD6Cu7kPwABRefuNe
56xHlPJHg5SiLr3m470FHouU+zIxrWQ0QJj7tQUarAw4oNl0TgDysdpaT3Ds
NewPnm8bnVrzhUqJgEn4PAfReqJHMJ9gWAp59bLeByysvUnUUjm3zBdrY+Kp
Cs8FVgkWvtCzAcWU1WoWVdBMwFMewpTz5Z9YmnpTfQWQ63gl6LSr6tAPlBhN
hlhTS/i+Jp+oS6quCxaOABd2Dsk7Li94iZxsK7RXm5nnnG/Hrg70gsBbDp7Z
WtuYUEBLDDhjGHI+4/6V4PKCE+ML3BErFlFldP8c7L+R6XJAfuCdhhJ8szMb
lJY4SWCzSUVJ5Wxae99BHQSIuhUQRP53wKYOBLTazuxD0ItXx7R1czQae8FT
AsmHJqlhB2pGsgHGuH6YWgyrr/dd045EElGcwWwR14yYLJlhBWf/a9ZCkJ5D
Y3LuV1b6CVEHacZbz+xcFet5EPH+kaWkigQw6RyqrlqfMczwgNgI/HunQEAe
abX+NryalGM67/OBjiWpiQJfo73pIsOZlXgSOgn7n5xkm77mREqG9DoAdKtk
hOdsZq1GPi2+kf8vd7F7I+UjmGw4CodpgiSypODowMTXnKJMBXzSL0U/ZHMW
QDJRP8YzvzJCBTrESJoATnJagpSsMiFb/X3FHWZfvUcQk02jkt1wXxf2AtEE
iz1s6CQVlr3aHpRCaa3nPaJtLw4n9LJp8yJuNgdrLLuifsLB8guW0PnHXtHD
DA/0TzfCLvDAF7nkL2gzBM8XZYE653pDdBH3jzpYi7W8e3kPKXa+QTkqhIDY
1GQij8aOpQc3ukpv/RNGc+HKQa+6uP7Yace5gUFSeaRBKS/cX6Yk7rAejef8
NYL2oF5d/inE4Kt0V7kEqaReBTslpcFRNwStThpGlHf4kG0cS6ZEKq3jplIp
vd2FyjE7veBFCyuwSLwBWOHxDXSRL1ihjIgPly43WuNhTW39MOyoPT3GN7Yf
p4Ic+eCDjtSwnGgrAW0XrvddwHqDe+rCedkLRSALLa8DDrAG8R2IMOxJsqex
QjRwXLa6GHiZ/hSroBJhXOzPb0XD3M+pqVy7hCVjwwlPaBlXz1awiLL9KqTu
WiL5vMZZY9EBUTBJ7GynqT0j7mLoe8xoIkp0Fp+zxIA63jpigxdX36Ko1oaI
vtg2mO5fGcxmMA9OIxCEsuiOwS1DJVGnWtZOE3NqANpjMc6rvf+/aVn279cO
tNiMQqixb0kFcJtgHVgBgQUix64smmMEyNv1zCtTK8vTky3G3HEaGadwOW4N
RIxB6RBWKTJ4OImpidE6OesnkWgF9YO/RFxnoNc9mczXo5oVlM8S4hqvOa/1
lu6Qs7TkKt7aQPgkbvTFa5CvFkjMXO/tspq8DyfcYhttPR1b5rlZ8q70E6fs
I0SQ8tR800aZzXEaGcbUVz4gsYawiCJU8B6ErjT/l2yyaRhOySmB7QrKQOAB
V5/fw8lfRDtw4u99DensiDdZ2g9N0I2ELIvWKcHDQfcbEd8y2UWaINLZW9H7
7r33pPZv1JEhpAy9+vveodnJ1kzrPiFmdTwZZynsyFEuPf9XJzT8/a2poRDH
jauxglnItWHA//46aeRjL4stM1BXWY5hrCrxXoDBr25k5I+io4z+2lbGOFyg
/Vex0DfmRxSDfAi/tMQ3kKOHyp2HP8GmRsxpea2hQQxpFkHiaUsh3pj0ELZ4
/dj1nKjPikHMQP9sNGwIlkTx9jgCYCYNtava4feMBL27zD1q95tcmZpscfm9
5eSqTqFp4GxjUYVo3TAiUJSOukV65nfMe59wfkxgfBMFj/M+y94XUby/eNBf
uIP1Eaj/hOQyAnsVWanuXDi/skYoECKxWuWggUWkoOcvFbHolpc7KsO7oH6F
prNCc2QSqpWMIbhUwlmYJeT1v+GpHYNNOhhmDzDHB5Np6IRg0Cyh5d2TvHtK
ZSxewkChOxz3o7868hzygL76neol1ARAejY0n7EtdyYTh70riqpE5kGYBsgy
1vd07/+8Z7/UBG89pFvtKCViKKI4yfqRnVDYui2KyAZnT80xR9dbFY+YaxAn
bkV+zHyxYAP17DJCR7+qqsN2DXsbYTwbs3XOLNXB8L5hUj4SoMK3PcafrVad
vGwHL4OwrE9jQKGvJXsPFXikocoPPktWVx2/P+Y7xYKKbYg48az5u3jklTUZ
sr2YQRLLHLGhOYthzlSqFS1bDLHJlEZ2CsF01ptMxd3LK4ejLn7aeosVxGLY
ysPHR4NheoI/rUQYYSErTwErO3Tt+3zM/NaelofmbJ1NrnCQY4CKcb9uH14L
DJ7SBR/7TXu9MtlxzflriaPDJulP76jXMMWsMGnFZoUlGD+QBLA3bT1SImRY
XhyIkss3dTqdn+E1Eg2hrfpclykyGt8aaT1mGVT403eTi8qSV9qwtpz6euEX
5M2ycBBdPZnv/4zmPXTEcC2cRo0r/KaIYGxNt5o3R/sFCwIzvdSK5Lhu1lkn
HpdXQA0xHC3s6+oM2OWiVDPRWJReCJGYLL/fjD4qzyLfbpbyEVOeZIUqER46
A+gw+UrvE3E7MeLnmtVecpfP4rX+miwZz1FbsNM95uJBRaLy7DziF/SmLKFc
EjcUiRJRO8ut07E5xGAVIf2cvtdbcMy788/d2bgYOPoBKBj5NjfY7jpL8KAK
/Q9Ut73oTPmPSEPoS7MoFlwnwMz2CxZB3syVuKv/4o8hdfldsMiiL0keX2bo
oZcbGZZZAKvmHN4UsfF55RjdI++PScT/mqtN1MU2CKh+P3/SKR9Lq1R34yTX
WxJ3dDiHHtLGw3v7Tzf+rp8vcp3072e2vAu2oTVlTnRot9vu3Hde5Anp34TN
ju1dpnbE81FeuZsAmbSk71UB/tvzeYWiMWUEP+BwaqHDFl8TLaq3sdteBqNL
KcuHuh6NDziZtAbkea0eS6htyCvL58Lrnq6J9VQPnD/HOPBFSfnlkbGqVmH0
v8LIaajpBweYfD4zUwkr1p5e7rgDomOG4Y81SOGkSfwgzWOwKsHOVVh3ydTh
hwFipJO03mWB6yE1ISqLK6i3QcpY//Ajtokbc0V8UtG7RaXVevOkNc4kESbW
eWWss7FONN7Gghf4wLUc/gzZ9Okar4RbRvxnfISqVyqU9RRwvtzsCX2siIvq
7W7gxI8BpDRHZQMpVylLcgSBaXMnNMXunjqMAzE98pSpnms8LHqfbXrQvl2i
STO97yJiHrC4AqGELO7dCceQkWcJA5lSvPU4bkg/+ec2qen626znB3kA1Sp6
B8+dSr9n6X5la3JAg5VenGDsQkA/Uib20GQ5uYDFbFJgtJFXa6nefcSUilCt
qrjEdg5MaUOp+nLXXbVXSEpcnyzEF5PiClMTXxG3voiYpYx+n6LhKsg8O60l
tszS6sxcFufqXtGUGamXO3MDkPf4KBEpltglGXDuudHK7E85RSbuwU6nlB8A
pkhEg7seovIEH1nbb0yJLq93+MYAOJiBGLfZng1ErbK+hFnVdTANWCY+eSA1
LQTQdkL8aiEuphrZ0nQ7fcM6MTzxEHaT9LNWUMx2qnBNTQI+u/KH6nQ/nt/F
oTa+HmOikp7scgEh3ijuYmVfrt0/m/6RBN9ujb8TqsSM38jqA2o4P/Wl4O8l
7EF5hwePXVjTACGdhhYCkZKdyhF8SmY3dgwdD4JHTjRJwWwuCW92bE99gTge
dSuGIaD3vTKjLnE8+B8hRuZnrcuqLmvpbUHxxp52w4jTwQJiUDb28suVADTL
WmZwANbB5JJ2pfi+eZVW88v2IqjkiTRs+M2bJj3dRR0ZXEZManRA/V1FY3LS
qebkYM4Znf8HnrerQwIWfq5PwGhIoCjZpqfxDge71sbQufy9AdZaY4g6mdZ4
U5hiltTtAYz6cTPqViyCtsrJ2vT+M+fCcCqBD/ck4nVbdy3ovBLTcRADLygd
Sawec1hX/dFqthbfcLKYTgGVhDcbsK1VVEsYdyeI4KkD1H7Zy38Da1Y0PtMv
nR+IUYGO1Wq59whsfb47VgGUEOcnWQdoLvV8wSYedK/CtuzygDlegc1wGiKh
ahIcHJaZdRgM0ZXXagSvd4AQdQ5ySJqxYcg4nSFTquQw3kqmSbgCQls6HZZX
h1Y5FrYy+CMSLUbKUlkmQChc9GyfaU23YZ/Af2ovQcHtNl+iFgJegm2ssVzb
DNUi+PZKy75BaEy3zb0ZiLZH+AJbEC13zjaEj9cNWoXnPQXLbzTMYi2bAg+O
OCjhgDOYmNAfeYNYv+5yHwPhb2V8I2q/mvHy3VYmv67APF1L/9k821Hd4vZc
9shHLnqdNNwHV52g+BGNpdVG/zK4/KOluuve9RMGyoxudDkD2xbpCALzQ+8z
P4XfPRYSxkYARWhlWGyF89qJffSuH46PChy+jFfIuejL3aHghmLLS5Pto1f6
SQkWilsrx1OYlE7Z3RM9ZayZPSi56LuT+lZddqjis18n7+myN9S/jgSLEK0+
gzTI2JFuZhc7aAr5IAuNmPrL+WR76u/nWkMRlS9bd/js+zt5Y5svQ/1y78Y4
39heh7T1/Wxm3KHI3q5NLEtB8wMMU9LiNo5UMmaRqtNUb9A+7jP+Ev4UqvJt
80QWsVAjQduTaZVD7EtY/7a9qioaY2/THY04RAnk1q4uURgqB/cvSQFKVL4W
ugbk7WGyshiBa41V1gMSy/hhtDEEz4HJ+2B5Qqc31/+iCuJlXeu1E8gHWCZV
469JboL8QGpB4IpLeMc0x4/3QAKLJ57xtbwZ2msXZ9CT0Jva7hrPSN8oYDj4
M/Oj6wS4xfpXEdAaTUa8710b/MxGkOyqv+zuU2y7U0IRhG+deteR3oezrOhm
Co8OT79VtdeDDUWr6LlNAXr53JGepXwqqvt8hlwEXJ9EqFGy44irwjwm+Nf5
Lp2jPHnF+fbZBeWejS4UHSh2qISZ1hNMxCs9aRu3fANmjlIGzMFeydZkMhr7
sSj5oNEULP0IiFxCm8FCPqz9/Xsm9JHcSsE/iyhB0hiOfj+V1D3FfRIqSzLi
D8B7yCIsq9O5gPuCso/njbtWK24QGWHokTOtCQDEi++CoQbniSR0SlNnBazM
KSgVghVpliTs3Qxi83gwBK4cH/NlKMKyvyj8XoGV++yfTyzNVcidSgho00Ku
tJRuTtkb97JHwTHGzeTOUFqFjFYUJN4MnFrFFx+1HcBjL7t8KkneyTBW3fsW
AxGL+bUEu1ZByGsRGwz28uk/qeL0pOTDfMXf2YiAqcwLM5T4g3kGUA11gJWV
8njO1GE5AF8gUevpYrqiKCGfdxk+ksPFKZanoxxYJBsm5FAvGoQBzJ9GrgXX
78B1NGY+2lSs0BJtzhRYVXfVyOAQ994WIQEF3R1O5CB4FNGLNxKVNtFsAbhe
C3YyNpNzFXFWsYpRjC1E7nad8+RNnQT6HKvxGp9Gq51JuzSMaIZhj+9E3nRZ
x5JCgaKBM/7zq2nWtIr0Ez0cg/XOCm4mtRucHGzKtdA2EQbbyyagHWa7nSsp
BFnd1LiA6gFSsVE6mG6AF8NkdiIy6d4+s1ZupzA1zR8XOW56jeY3LtgQ6q+W
J0vqlHhoO7seccduUJ00UEC/qxhjDKfMl3N9iizfGmJ24CtEjkJj29PxsZKW
Pyc3MEjcoQxxP1LD9KLwzusCyYx7iIbSGH0zU61kUBNvh5K5TPmTjio3p6mu
6gHtCx4V927gtmwBiACYMWVBl1FeE7/ojv348UKeNxLiuDRWKDxztig/Q132
0fv1ZwIYhhoQ4dEooQsUtDZ9kb05Hv9hZLu5PMM9W7R45UtseT9znsqGj1Cn
kNZz1/bANdZAexep7pZ4oPCcnHGU8HFglRqHgivcbNDpOFmx6ockkX6e9zGW
JtiJoyPC3wJ5E6mRzUN8LOPnHqBqOFDbh7C5S0tMvNJGfaht9PQv9MTCSX4s
wv2fggdXQNihrtECBB6mlzSCeVjVJKs40CrP/qxhLp5Llt9bpfKjYkRQ7i3w
lx1Be4hohDi9fWrMo+8zRUrhOMMQOKS/MeFpMIhEm7MpEgxx1JdfRaSodqVF
klJGMK87QmsnGAyVjXqvR43C81+pYpGOwVqThFHXTcmyA2vhOpFCbcjkTvx8
/pDQ8XgScZWBHp6g8nQac046EqAwbovhwnb4nNPLrq+1vIc1ZW+lGXLYkV89
lZX19GvSeVwbJ2tHsIqiFpoVBhN0vnQUB+Y1BgLDXrl65ptImh7OkH+d1MqY
wVCgLbEldl6RGZDuturTfDFCNjgHFnlVk46G1n6KTl7Jn4XAwGVTdcHbbMok
bQG1tD6NRn9ZaRxMDjcmCz2RXI8Cb95kOVJIihEEn5wgO1SlQhyrA1QZeoFB
PJozuY5/tpxJCDVtp3rxrjF+pb+CBp4vsgr6/5YThvRdTXwpW3wtuy35cOil
jddbWIviw20/r0yJrnk67Sm8bgw8DCv0eFGeBMANxh0p84rOteg7Xav2mkTU
tVm7tEv4MNcRqa0rDAQGGQfZ44qFQRx9p1P/9/CVOPGuHoYrNXe/tOaRBIKm
LfJq3tNkgf3bNRaEdlbGRLEYzk5s/DRXmXfdc1JGONZt8z3VgQH7HJGIfDYR
v1oXXGLYgZgm3XEMZa1n3LJy45cpoJAZpcM/CIimMiebWPmROh+fbza5TH//
2yTw239yjaOtyTMhuX8/DnwgI2h9YqUBteeEBE98AEH/MqAFSlC1jethsGHt
0KTmYzAcMe9xdpzOrwRAvtNZZB7spDD89N4p3PamCAsvcI3ZpDZoZ8SwnjFz
wtqqG1ejwJtrev7UPj5drHelMuDTfYaVXfvhZvwHyx7MggRPbK7nn6ADAgSl
PJtmpQZIMfB/fqLSWxezbEh0Qm9s7Yy7er6nmZS4+OuYJ3018dO+pQD1R3gY
LM2tWmaqlAdYTZ8M0EQVK+PJNuP9YGwVDxk/0+ksw43/7k6LugMhEFEA9NcC
NqX5gpv7hHNlMSv5S5jnYvM2uXbOPTvu7MmaK9TaAwXmm6DVcZ01EEnE/SlI
7xmO9iZ9kTUqqpbjO6MmkxApaM43ylZgechZySyZrXpkefPh6pI1PamIhCdT
VwWhybe9xTsgl2KGzRslNQbzGyzzjkiLcTYHiYSdsaso0bPqmYnVSAwGoOiU
plf0/EomXQmdQWKaKYz7dmGz3nX2VtHA0LQpoUDv4Ih0uzqztYY4zHQehjbV
zZm2hIJWE0UzP80D9eCMr37VrO9JvpjFv+5G1qG1BPizzjaI52gPdhclx026
XdBWVsLRHNw+ZFaN0bzJZrF/yXyhwUeJ88RpOQwzzC/2KXOGDnjy/CMlPj5T
PyiSR7+6sauiNHSBATM19BsSgtZqSs0O/5K7DUbstbdOBIWfVnSn5n1Zdz2f
1VkZcnf/klUB9bHvzpTqN+KbRRn8hITBLuip04YLGQp6o4/f9agv1WgxW5zA
FIdMXUIQxVyB1a6slSRIHz6e6VeATJku+fJlBHd2XYJsi7StctpOEKPOVCtP
+1gi+NIfOfIKAv+09UqZbDFp+FnMRJW93AcPAhAEyNMLlWQ2cp/iWRyW+W3Q
VtvI4Q7O8gCI+FhAOnSFG/wDcvIVKd8iUblEdhE9s2p6wEPbWdw1BVH5uE93
aFSdX/ZADRb3+ihkVs8h+fXezv4I+k1R3HRUtZtjHrzjLEPxycdz+wuv1EAz
4krVmztyaX0jvwa0JDx8Y2R/6HrI39cWITWJGnRvJvMg8j8yb/rjnYMtIqB1
5f2iqFn/dprJqFyeUoA8z+7LrLUV1hDNK+6FI/XBMO4+VIwpbIaRUcGdjisR
VSkAGM0jKCVpfoYh7Tlv9JjFE8mHOP4DOIGGn9wzufLRyoNtgjn48ZDi3+Wz
8Ww0OEjzgtlxWF2qs/q8lIV6uDyBOfWjXJRVzbLeV9kD/n+rIofb3ei0KnMM
7ybzu/8tpcGjtXnHYRCz965m1CFsAmG3se8ZgyTyboWYXxerCsz5fRVlKD73
2QiZEzXhP5coS7iOGx7XFA73xSg+IC/4FNRNTsAiKNnwoRKZtiJYrIIvLCzj
dUpB0rpbtVxNcXPffY+F1dv2OVkStjQwiZf4ZKSJ7Z5FYdcQGYMBhL9Cq7CV
vb+CND2BonaoOBo7dIYnG/QkIlxSJeowd9CQD94/dKeowiyy7SfKG2q5Y68i
T764oxCd8tRrdXMZMIoJviSShR/+ghknzLfDnNBMQy5B35CXl667BL57wdqV
ZfBTJs+o9QQCxyLNJF1fbxXxa8/xS/M9BCEvDCNKYHSKPTXFt5sbTGIKAq8S
pdo+s4yOGgHqO1FKN4mliwkpb890XP6byo8KkAnzF9/48GvZMpLgish0soVA
hGFrk8tjVK33dkrzv3fkYMzR/y4wlmj6lAoMPQa0kM0ync34gI+jVISV35bP
g2uHN3pFCi1osaH0Vs7TbTXqoiybuCpKf/63P3ZKGLR9wtENmDfUF+9ze6Gc
4dYeNWOu6DgLzBX+tgc5IYIR3v158hlcTnnZrZ/zXlO+2bIgWlmez1yLWIvv
Ou12e7IOZTyem5/gxu//sMvbiSrdKyNUaHVZ4RMf/iE7jX+3zkbqecfdAoeq
3FFEqsIkVHSHUfzHYO6/R5n6u1a9kAS+kz3B0x28Yh/mA3ISlHw253sfmMIO
xXz9H+MD3Lum7C7BKKQVGvq1o0GXWzG3Fo7Ub2Z2l2DXWZzRF+yC1sXs3tSw
USJL9cd51ndn6w22kH5DyL5r2i6JoVauQ3Q4O1Q1TmhkZCXbPGyKALl0cpsF
A32h+nZp4R/JIr8zKDPF3/Xi1ySKxmcoe3vJ/fdrr+FpZGCOGbR0YY1+GzGk
U2ju64Kx2L0Ruv9kjL1Fkd5XpVHbzuD/J4CCzPufWVnv8sHFsT5AxegV2pGr
lcStg7BTqy37IG5KiPialViVeVP+2gZ8JJAPC1jE/gilAjkL8M7wZwdzZPHm
LDhd0ypY9nfCcEjRi/uPn60S5sTQ9XbstI4AoVdlpKgEPt91zukdopNWqxlU
toME7+8IJR3hU7snkBX8Aac2grm47H9RCL4NPm1zVec8N49Zy+QkV16xWCqF
7HdHG1stBrV34KF5657Le2CwhmPpMy/1HmdPO36GTNnV5y2FrofSVWHUBWqn
6iEJxuUPvo/XyRQR2LupH+koAcMkFBFInG7crS/QByFTKpUVuyYAL+cm7yQx
yKLYCzCyKJYRsuo1l7pmd731n/+J0tlxOfWctmVJ99LGrQZJCWWp6FY+dJqE
xIcAgqUZajbxKbNLLmLtDggHrpiT9MAMiTrJiNEnr646kaYWp669IFK1LHm+
cgmef4pQMcDiCvQ3mp3JJSAVLMPfdNS0TGb7d0azbiC2JktxUNh6Xh0G7PjF
WYPejgcpt1RMf9dR3KUSElP6t9aX7PSb+InQ2nvj2D3CCUDTAp+/+sVMVGcH
6NWPoFIlkgdG31RFxUcbFripD9hRI+ru62azyBpOheQshgglI6M87qQQbI8o
N1aRFeAnYOFI3V0Jth3dfnOpae+ba5r1s212Z2MiQVYCRSKVOf+faedGfMh7
nzjQDLvShdz/saI9uTcdWCP73yDHTFXFuHFjjSXpRcqxBEGzKGkOuvqonBnV
Bh8bkLuPcacNCJ3YAGF/1byew0S/qZ532LNn5tvf4tms7TIQ8KS+HX99bbUk
FWUocDMQEEglrgbYAuIx/tNuVsqh/wivjvkNGNVtCdBSHcuMdciZ/nLK5Wt8
uH/lqiYbCVFzv8NpinG+18/NuuvziAteLZsd+uo6ctMM2Vlirl+21PnHFVKt
S8iVxwhuVitwKdKKX8Ma21XCeILr8/ymbyJ4wPY0UMAu63w6aup3rkxPyAbf
7sMXmrmzomdHItImtuu9uNgYjpq0aZZQZclzIxLuEZOXkdjBdfMSHjNTFVIr
YT2kIcEZ4DuFmrPNWUizZoLELL1VjjTxuHMBzzE1nDtT0Q62gq32x1gUXW3T
oQZu97hPpwz6zk8p4fIW85xI6qjOQPAONFF+nKbmHDQT3xRqyNnhrjCWwTlB
CNJIjQcjnSqZAQDqnxIM4Ux984PpRy+y2sBUMc8H9qvX5JLEnIqopw7wSM+d
Fk8cUhu1G4TRDkZVf4pwtDWp2ys8L7YwKLv4S2FPnqTJYxOthZCvBWYwF54I
7Z/pCfUfIfH2gc9NPH8Po/TnEZvR0O/6tfSdt2jKBr+apneejVlUAkr+oa09
qbfrk+MKNMa6AG08KVBZQIDKFeiFfwwvTHejT+p8lucaj6x1p+1PYqFNyq9v
UVwum1zJVAi4q0+Eb/B4v5PZg8QMfQbGSLCe/P5nXMYgXFSkaYNVRP8Kn/JC
3Z9IUFif28fB7QMJUXrNpRjw76is9VzvBrnC+JDo0HBHF3XhnkMe756RnkRs
6P98/mzP9zp6+D9/CoWoDJJOc5XpjjY2eu6yNi0FCWC2sR+7ibDL9LAz5Jz9
Db/K/OGWYARcehx4xFwMDNsJNo/YvxG/kMck4kYQh0B0DdZMKSTq/j6FV20A
p/YbYX4VcKIYlNHuUPLhyn60Ur/nfAWCWxl6NdHihAo9kJgR5bCSFAa+9Nct
N+4zAzJ3c83DE04p4jnYCreSHppqSsHENqK5lil+GeV9/R/o8PiOcZ6/IiAX
S9yCN+1Gee2B/P1859mHs+toZSHqZ7MpAdbzujxyFNfsR4O3F6P/vfFMoY5D
19pcURsB5l6ZdI/kxXW1vkXBIJQNU0qY35ROGuM2L9DUOTIg11/Ijq3heKBz
wdWqpvyZDKqjRs8OQYy7CzuFQgE94e/fHL8JP2DlZnbTowtTdQ73ovPTawKr
b1JC+rJTh++05A2LcK6/rVn8c04F6vhLyxI//40NALXS0yT79Xb+0cCxl1M9
hNEEK9jZ1I0XSrZbWDg5cXZ4Z10X/A0b+Mn0295PszZahn2hMZZAUnVHdx7s
WE/tFAV2AR7TXO9D5aA4rRszZZWahgiHCPd1IqTRMxxIqHU2KfYw0Dcz2qgD
fXuzsdNXRaOnC01iFj6pyJNhD9dot1ZTiYOZelcFMS+R7A+Vbn7OrheNZMoj
70c/xOY3EmSSWKyO8D2DqHuZo47AHT9gS5+UIm5Vb3x1mlVj7cS2O9OBB82f
/Qb2tUW1JYNw9fSGam4L5DTx+saqCALgGJnUISMxubxC0Jwwsqqo/j5eQ11u
ZtaZOigFPMrbpsxjqYivZpwwfUAW8Tx0a+bOUFrh8G2a7Ff+Nic0fW/PHKkt
zszwY8QId3YWSNEQqSj4VVqWUFzrbswXMKa2U8xVUD9O2ijIoBqOvx5Ct0e7
aMMHGr/34b++7gyfYMjrh7Jnd/ikof3SYIdbgV9w/d6B/sJtzrue2bUjhIn5
TP/7mDrYQLyPDbDt9SdtD5Fh7jqloNB/P4fljM6Upk0SySuvPhH99csQKgBI
vPvn9mDFn7vDDp9Vi0EdApw3C7TdgCi1iGOpokizQXL6M4lbXXrtvLmcV0wV
DuiNhUT4z0p48xboj3foWrpH7ARkfctWsLcVj62mCBJ2jbBBSGOi/wVoONDX
2qZ1gcFQVeQLuDyb5oqcZPRVANewpGD24rtVbfpmUWGdt1+RKX9xsF3EqUoa
JjGy8qsXc+i8jYbfZ+cqlO/idJLqTxm1j+uqs/+dTkRiMNUEngU1WIp0qC9H
u16rnOkkhdtM+W9S6j72G4/RTDoKfUgfoZrLIeeOktw+0s556l7/rr7i9ejp
4z2SsSCbXPf8a3DHEqUqt7hXl2SrW/8pnP3+i1z05ZiAh73mr9CME0KIxUda
W06/zqQHLpaQF9NX7i3gnVivA8B4scJI8yPag3Yz2R/05Om6kT3xpS+7ZsFE
HjNvhg5eODM2MIWG4iv0yVLI8ctpymhA5zROrKuXi1clic0nsoTApGr0Zsq5
Ey18U/6ui6v+WpY+DQ1bp+eZW4B2rBVFJIVud+oD3vpl4DYwleLLLTgV4Zsp
9KyGiIkFUUnB/Xw+pNqrl2TUudAzKV5QBMnrqwYDM64qn0Re0dyZHUUFN94C
zlY/Omf2e4zGoiT6PeyJdshqe/zn6xbexm4rPtyvA4kYfC4HZWKjXnX7R4bg
4oQ9q010onjbQP0IlNiW0/yCpowKw7wtuud7MB/tuQiCf09fX03XcLJfa5nb
78gjRv7sGG8Cs9ijytky4fiHa/Ywc+2rme6sL740qTY4AxuqCpLjwuQw+m1r
D0/Ocj6d/LwMhHyzFz8WdRAgQ4BWFW1qV87bO8WAee28JeS9MwT9xTHi0PSw
w1vwcukhUDagU1TMZnzU3frEYn2J4YZWzlk04ofSQkepPeQm+uwhiDms6scT
ecUDi13+KjV8eOa8f6QWsK1hHnvP4o1Pk2ElstfTZLX5w6d/tHv8PW9BwK1D
4GyUFonA5P29rNHX41G9ggAN3yLvaBAI5bF5CszpopZ2CkYsgPYWiB0rARX6
ZChe3hu0311ZL95RnywBoSNW2d+EHobkgRy36GfTF6jz7SuogvK4GAf+eMGC
XGPtdIPL0yOqexuTTk8N99kXkJ1xHiqbefoHgEGKh4BDnCM8Iu+qo9dUMH72
OOh2doKZAgtp9kf2MBqGFncfhIRlHhm1fGRJnZzKvG4+mnSa3oDVFbMWJbXf
plPyAQH21h7E0kZZLBpPwVSzpx5ROlZPWWpLivQlicI2es3nWshUb0nvwkiV
/hQeyF3++VbM4qkC1wETPx2JJOU1A3WqDZ5eVKYfwayHjuZ0biWS9t1C8j8P
HjImztz96mAKdpI8EdbO/Zz/OfPVMt7Fa4uV+BKH72bK0KK1nbMr0KQyLx2L
ZcjqD3Le2Gz3tzKsOGleGM7moQ8ypSmQeRKEDHZA2ouhJxEx2Ijd8ElJWRlT
TM6MwnBqYBxZRiXYOz0bufJTXgWyxyt9O377/7ujw4cvyI+O5421TCQ5qh/3
Qqws9P42cB3K8RpEtc5JOQZdh4iYweMfEpNzULMaIFUnPz1O+onehb7lvQIz
OV8aQlthIbCYmctzQZk9++cKVKjo49uANhcvMW6lTDp0A3KFRWwrQkGfn5Ws
Qb82OtQOaeUAdfbYEj1ypkdYha0Px4flZcjWQY6x+DcnhrKwLxLoeFWnSKPX
5WDJrGGSKg+V/OLTPUoRqRohVcoBpLbIBqaF1UDxFjZ9XzhHrOsg3h/Zl1z0
5bueVZV+ByW+aWyh3Jol29bqJoeSuo02QH1t8ebYNJgpNF/rDtfqazm00WfC
QuTsPrU7Oswk5x0PRgfOu8gxn7a0/SRIe3ByuUx0a4ChkWY3odOcz5NtNg8D
FmdB2DiHFUcB8RnXGNBzmZqT8Q44BrSjC3pyLgtGJtw4Kvvd4h0+qBHLzJWE
aIRQjYNsab341v5AMFUH7Ze6Q+NTgWqcnMm1Z4r09k0w9bQAJ4oOPj3R+ZmO
1vD9ZXjzcGFTUr4Y2hLAMZlRZ4NVgHmuzVNxiZakmJMikvwxleJj/12dd2GD
QnyKM3WJFsDquyP9mvw3PE73njoo3KkH/16uLJ4Yfvc+x1FJrt1bbna16BpG
K5homt3IopJ5/IrBBxpvqI9mrtogS+lL7iIkH+dWuCP+/kwke0wb5ClUD2sh
UXnsH3ti4GuvBA8d72jXxpVQ6tMltjsghfGHbOzjoR9FtK3REACdG/qcQMlz
xLEJ04HBHLg01uDawoXPU6DUzWPZOWCnoDKU1dRJOsGcDcSEz3IRpKlY8Sme
mDqnxD9nhVSbaIMnNxfLVWHaMVfvXmHjtRg3oCbm2A7OpAX8WRsW3lj2ZVZQ
laSicwiIz+Uk4gjh5Zj2gVMg9Hk5T7g5MEaHCuFGiMQolRPQRrVNlXsrTIn7
Tv8kwvJ+wxdhMnAnNTBJY2yrcNrsHWwgD4Wwr58z0kzrVgCbwJpC3JdT8Uqo
P5ORz8OqZ+e3zqS6j1jlepN4KLb6SmJZD42YwySTCMsBFvKyxw0mr5/VcpC2
GnpcXQYdb7cSCX7z0VRuiIRkq59bSaCP9ccDPGU51eSLM6jBh7ZM6AabPvvb
jdB86eViY9d3UDg74hEB7AIA+hzTp2J2clYifyH3FagELuVzO6Ra+k6R3bUd
+X7tXukvNtdLPNL/DUVpOVvYqGZ8cq63L4RF2ZKI7Vdo+Xkw1sblbS5pfC1u
FlHXFeFy9KjHVMUm2pGyK52BkS5Fr4o6WoMdZhq0MvNjpGr0i2nKX6zbq6mN
d1p7DSEgExuwwyzNFJYEPULPs+b3H2rQsksjY3zP1o8P6WYkcRVdDN5hMnR5
MWXKa/wFugYvt6WLNE0+hpvdrpZLdzCjUqVJfEDcl3X6YIScwGShqiodS+EE
PJtkH9GQsYAXNa1GF3/aSeJ1I+QeuYw+F3Mg+ceq+APDntQSZonBD00rmcLx
qADcuMOwkWyQTbabUrcHn4fIUE6/r9gG/aGZDzURGIkXMG6yg+rZeUWgEOeR
TbcnkrJZVZ7e/knaVDKlv+R+e4rPp5JARhdgKPQTr3eLtOxJ+OwRq8LUvHFG
meN0oCjpMN9/ZbeU0E8DPZAgL0RfXOBH/H3tMa8IJjd2veoyKp9EcGRxdfdZ
jU5jipHLgR1JSsMQJkWYhUxCIcEs2VkI95thlZ0hLON1qgBt2xuDsBoKGPh3
KFgPwCs6rjusNCV44TZc2Z1e8xed5l9Nqq8Ig/WefI3WSGwHDEibNywMopPF
vfJueOSEVP9pXAFWrWVHDkORKuITHzWLTjhntsddAGDx0u2dw42HS0YwlSLT
ZnIoXq3vULmoclrUN+9Iy7+P/qAgCSaaDIKtU5KoH8a8J9d6+0NWitrsU3UC
u9dUjUAnYhwR2LcUu+V740LX0+5deRyrVK3B2Ga+8Rt3ugOZ5ckwsUPKkULZ
+tcjkeHqoAosximKvAoNZ6glkslr3w8zA4anl+gQ0zLd/UmQ42If1z5cI9py
U71zcKtZ+S4wESYMO/+Q8wP+HwsTLwT8xJbesvhSLtPoCjUo59IK+99gimwW
UX/T5ReSXDDkcHwT1506xOZ/Pmb1PmyX/JUq5d38AQTcSg03wIlqOjsyZaCu
8F79wvrKVXK8rn3KgrvDzIj+bvxENgrbFqf8xKrYTZEbi7bMFWW9qsWaWP3P
BZEiYLNgE3XDNk1kvK9vBy8OkcGu18cBXTUdgLUEu3Pg+zWz5l+LWD4+mP/n
GSZ/cPp/ICOSh+BE+OZsKmfpXW8xkvnKypkzvj7z6G8B0CqEdZni9Us992YM
EnMkLg4NX7QrXiK2MI5DS8XlB6MOj3gLzPu+PX/tDWQIgkcLhIlzW9iy5xMW
7RJtPO7iSzFoDlXdqbC39ulV7/Wz+hsJtn75L80Rj1a9vgqfFHZP/RL5CMJL
SQ+gSWAY7c3afoHYEvVPKVwucbeK5FPrHdXhyCtHmGDKyKu4u6HrpARc3ZRn
dskfyJcjIav4FedWqA8dFWu5YChFi0sGMJ2VeJwks+KEeRES9dChR/FMGaDe
k6Qw4fFryQjQbqrl7GwsSVP7C9/54YUp5NaJgT9XOMJmLb0aUh6Ndo7zBbJg
IwpJsWJPMLFiBIsT1Iq4PSrqCMkpPu5236UQy5dm9FzaKnCU62vasce4cf69
NuMJtr40bLYSqwwEFApfm78QS4PIuxwMRKZp7yIKZ4jeLbC20NDS7ZYWkuzv
yQKwPab7iQW6QSi/PbASHa2+bFnP26xCBbr1lnF2k20A/lZyZUoELlUQxbk+
RLHA8QS/Opph+U7E8hRKR6KNjIpF8EKc75/xouiXeYcSgNERctG9nSZGwzfE
QMlbrtSXL5KjT+E56lrTx1SFJVs2/WOQjDRMxc2ifcvNmv+oRqovUft4cO/I
4dLh3tmI0ZIerbxrRvVdoN5SZdDX25uC16/0BvXxsAZJ974hmcOrDww1DbmT
PYYmM++kZ9QACZSu+DxzKB8GGt+jBXscU8fPwruKAivuI89hOVidwAg3ZCpL
4Ke8V89e9Cm97jbl6tulJXfXuVs0KcwgQYc/tQ7ErNLwa021CYnbhBs9KiS7
ck5J7S4sGCkYLQVLQGuXtj2jVv4fehI0n+5NQFopzW/MdJ5OAOFw8uj9Ecfc
hxupIXhJqtJm8hKhwjD9oStrKTihmpdNy561r92NSZi1984WQ3r4BWAKQNfc
A0hBz5m2CwT1NnRgovyTCFSuZzkOqTfCLdIS+nyoy5ObXbOXW/PTAx7I3QUU
QdjS3w+hXOC12C28BbQZsgzzjSo92WOboPXgMKJpF+Nd+GFLw8TK2v7ZX+7v
yx0sAEcHna83HtH1T3RZzknmYglgEKvBBqJKTzPIytdHWj3wLOC0YdsHuwpM
TYCUpw0p7aivScpkCYJOdJMf1zyq+eFNG0Pr43P79VSxZddHCm1j0iDFDbmn
ZxSwtytF2Yc3TL2bPiaWczRJ1xTU9PyIoZua+uUM4+ovBj+mCRl9+dTV0uv7
7iIAwuhk+zr/S8H8D9ULBPr//ifLV2EGPWF/WmlYwHj2VOhfqV3LjLTqZiH+
CQCjUfT+mz/spgattBCxhXTklw3SwJO8W3TS3OF7CMLzjRDQTq4qT69c3H4O
aOA0UBSqYDaCcvEw0JKHMBU/jGuKctTfejRCEH6pD6nvQqWvouC7ahoDsAHR
PUiq4SGW8KB+dIbmXJ76jOdAigL7gcH7WXlXFQpsD1YaOTZnCdzGlaZpz4Bo
6RQVTt6pR4XP4ZiDP9rn0xIUMQNBLohxM33I5cMYhVPPd39QnIs6w7YbX2Rf
RV7PsSZx1lJu4Kn5piyF9CYkACkHTHZKJbZ4aWWckbmJCljBIuE+ZIxQM8OE
+a+0ZlJ+QkoTh33/CQZp1YBUJUmFqGCoExSRyRPNpOV4zemN0x2dT1f0db0+
AwwHAux2qTq11eunkbE3UyP5aRetsCDOHL9o9PmbwCcW6YxTAUEK0CfMt+M6
wA5RjlkY9MPPrPL1MfFSEbSwjNQ1XRv5eIWrSU9NvZNWwbo2Tbrenmk2quU/
qu44uonaXUmPp9oVdFXIUOW/10VE/VFN1arSBU4Cxd4xdpxsqzJBZ3PEPiPm
li5afPEwIW0jWJdKKJ+91VHXW9GtVZB5ySxUGUJD+a/55hZwI2QvWk0tXyEI
vNweYFkSKjA+10QytU4f0i3vLro1IxFTUE3TDKqke0Vs9k97nCsj+LZm//4o
gBQOqfuhEOizqRoIzH7mkGJ5/1dypk8ZcCxBqEXOV1bMAWGHrICSj5qgAg6O
2zT+/ozJiWExae7Kf7J6iau9dWYqj0Bsag/L1ZgjYxW69jr81UZLNBuvE/8y
eHtP13cFY5qKP4/C+Xns1r4l1tuNxvycTX4fDAGcbVwtWR94OpBj/X5+UuIh
IDC/EcDa0TUOdjXhBggU0oQ1D0TgCkuv2S44Ju87MXRd2nSkRRxkXVqY+t/4
4I/ZKnthqs235JUdLuD6oSUvBcB0ywI3MDrRQEJZQavuf8kGvuXWnhemTMHf
7eHL5n5p7WgqC2TEXEyF4s0JOb1i1AxIjWYeo64xsNhw97OMs6XIfWk29wSS
SwDsqJEHis8FaNvhzDRezdDtXsEsPgI1ARE7Q8LGZvAAMAwhFUYlF6w4ba4D
pP1o2oTMeEWJhXePg+FEEZavtmor5TR2jSWXtKsCGC57xy7MGufyUKlccjA7
mo/sxCDJn0kRR/wH7pSBMm+TrHg36d1lCROyMuffN869uZtKGHdKYJPalsAE
oUc9bwM0gBouHdx6cf6+RU8zefQ2HGZ9B93SZHWqXSePou/T8XSMQeJAVBZ0
03isKlZsCqBmOszJOgnd/CIKWLO+PT45/QwxIGZVnp70AzWPED5BYQR/46Vb
td7v+kYZkqfSwI2MuXI9YBZogZLWKzOlTGgYOB8MIqiuVvjy9F5atviDvlye
rTbAjMDBp400QUp/zrnpDwIVm0SKshlELOoPWYOjGUKuGUYMT45rAO+8KTRd
Egow/IEDETrYROeaTLrDWTeu37yDhTx3JOSAJkhLk1wq4ewOArMihWoulxHN
ievoyPVTlhylJY4UmdilzCncpkdYhccrIEKfuWE9djsHCrI8aunKSfCR+X5H
o4TnjAbXP0XJSyXXzuUkfcazfdkgV3FbbiJKJtJyFMi0VrExnJSQFM9Qxo9j
Trn8AjFYDBaTffu4aekj7swBM3M9Y688JTYmrrU3W7I8U12VWzhrtp/YHIna
13Cxep5NR1aY5ScsrSFv+yQvtpscqSPTB7EnMoNlIGSpCBJPnIHSIZm5UfhN
Ad6bY+nakWtkNlMAd1jDjqIvzpfHbIkxT7o0s9/sQhc5VzbYJE/Xv4krPUfl
wrigob7d5hpJF8Y+Rb9MQlGbQ2BKcXxsHYC0HFHvlo5HcZlTDS7b3z1XtM9Q
3f3ctCZkHqDzubsTCrQpRapo3YvJjPMXcBqzvB0Py28N5cbJtXjsa5WBv+eA
RHBZWHlzU8rlqTYI468IfQjHvMEyBfwf/LUugWdv7vSsr9gPO1qHPA+lTLtG
J2uzqnupSBshr5D5x4gyKfzPq1J8JEaxqUNm1XpN8wugpZwRI5x95/sMpMSh
wB+oAcFNdyzYEarZURcT5UgLMCAULBXfvZohmIX4CjnUlKzK4GlcRFFOAD9J
mi5x6zNg7SJAcS70/fQHXZJC95Vh6QUtW1SvMbejYn7OF6qASsnRkTx7nyMM
Xyh7vgaMzOH0mCfWnS/0M5+iWbV2VRPyAx/O44BrpgL0vGqOGyZ4ye9SRouD
MRw4AUvc6M2/22QMde/FU+15etA961uoS8X3T4DEWOQ77sDIGQJZ6SgfAHCM
YiE4vn0L1XV+C1k8nZKMW1oefOzTtFyGX3j1tJjLxHbSeO1Ot88DrYYQI14T
Y3ziWtn1+M+J9V/FCT0K39Y93E5lSGk+ftcjYUpCqdRKg2b8z2z7dNTi4Vb/
XC+lfkQ5epUQtGT6kaYdQQdqWjeDzmyuPCEsgxRZTALZWcT9veo6fsSjdnN6
NCL5pJL2Kh1jVXzdZzopy90kFZGoIi29fHrlaY/Fb7hP8fOcdDDWLC+uSDQD
jFEXMkmgltbWfQn/UiOYTUDYmzH1MvGN6pOarYZK6ot93qPZ3ZDZjkYOmyFi
vLtJSgp0TatUyIGCFaQFioSS+D/NwOwvmR1bU7Ou6nMcEeTWiUMAuxZl9kF4
3HNfkcVKa1XviaoonOQqp31eCCY8oubdt661yde5PDPJjxljCjThYV+FYLy0
p/c+rForUTVl8nHUE0yZOkWXmxe7QyNfoXEso5Fp4RiIrBljdC0jWFclkFw/
5QAWsP++gr9VKF0wokKKkeZWqmLx/GW2CtdvP/n/jOpm9HSeGM+x4g/wjG/G
P7blMR3kPSWNOm3zb0Em3LP0r565+kjkkRBUGWKhUluXU9Pn3jdb5ObAIa3i
KeaghpwlShFITl3tsbOoDA8rwjQj/V09VN7w0pLStq9Jxd/nFAtEVTNgCHhd
A4WEfTpOuDK0Ea3XRWtlrgaYHUwPkNT0auE7TPm0jK9KMp4mAH+nhVhHmu2i
LgJoBhWkZd15ZoqNUMrUqVGmaRVXCf4TtnI+YfDYkiefwXIocujBzRq+ueBN
YpJp/mxD3LqiRMYJPNJz4BOFdOaA5Y6NBxhs4fGaqGfz+9PN9/WT9VxwMLG8
qcqP51zDSewwbOLJhbCneNmvWhDPbRwRGuORH9XJVXtwn4v1WaUUDfaBJgSo
EiOyvvjgWDcMY+T52AglVcut+Z0IFyD4K84lzb0+2cSDrqSYUON1Wq+MwmOL
AOlHoABsGkXUYynbLCVCRziXzYrnyUe+kEjYfLyuhO9Vp0LBGD5PphreznUs
QGKU8A1gbPgcTMJAf37XEJNkysZOWPRT5FiYHrdihEl2Ivq1on/xsoZp8RGc
3cYEdWyN0msx6iBR2760B2/3dfR6rvH7WKi3cx9dKmXsI22di5zFzJqRTQhe
12/ckoOiWiiWQRzcRbBNJ880ZK43DnyIgacin94jjUcxkufYTCj8t05z6X2o
vO3ZjgovhSP6gwL1iHSR68BNJc6TI/XQOcERI4I2nLcQBdqt4S28dB2Chlzd
hNbok+w/0ebp7BtiAIRJaj+DQSKDxASGAZOK4oC4Gz24iZav0ej7TR6Gwo85
LniT32rCCj2U4MYWPtu5dk7ovlI5Js9r/hESxJml9GNCsuz2KJ/GI1KX1Krw
Hn9uui9O05w+u7XckLwjqOp3CGCUXxmwAZWTOhIbYADvYln4B2sQuj1x5Gjh
hqp1FLO0TZTX3UWxqcycyiF/Wncywt6PrnxV4owa7n6I0dFn6lmMBy4QzEcn
CJWdtLV2l2XPfYhX0nl5814/HgGAOt+yC6FnaJnMSQFu0CLs6w1dleOmhnAK
sNfXbmqtYaI0Ebffc1QB70OG5+DjOF1RZVYqwBe9LXBociobqu35W4ku5gqa
dceG1DV8dDm90NowRxDcZqioSTkBlagfKzQSqSRAP8JHbXdu0Ta7ReZXe7TR
up4gBmX/t1iQh2PmhfwMgmrQTAh3gRstsZESus77st7MtVemphCBQ57tfgCm
ihKZfO27tX5D35uzpXLtXC7RcUbmR17gpGrAAWwJCKQFhIDXnEmGq3mcT+ny
uUiCfkpjaRPWhm0V9mtLhQQTTH7TgekIhWP0148Ga07o2lhhEOUeg+rxaIDi
+vNbhTkeI02PAmfCmgsYhsHKHO9lbJ5JKjs/8Xsola/PBmmiHkXlDBtBbkrf
cfZFGZ/wYMTznVdCKVujnHl7VwTuHTljEn9QzaAn6QPYtEKZvjEwIr4gVRxs
O2ZT6dYEUFIY9L/9hrToc4x4FEXyCZyE4/JTqbTBjQIEgd3bapX4G9Dxrmiw
tar1rkq5fCHozAzQeJz0gl3lbU9Y+PRsDcx/RcFLn6vWClyQDiaI+ctH4+Bt
bR4KRtTeV9B0lk0eq7QRpCnfy9jknEMOCVxUlvMFzcBDs8hbcrwhE7KUmTwY
fg001G3pIwuZLwsemdbHTT74rhZC5rKo5Aa6tbNlLnfDbFVGQtfTTLdXTTXR
X3BkQe/UZojAQ+2xvH+Kd21cEjxnkPCSpq7qfQD6vCbcw1k+unxip9tsa3xN
uZqO+61+m/wPU6GqFaaSkcc8IAR+D0bLcWwxVE0fM0+Ce43erYJ5KD4V0JF3
9B+2wPg1dF5h23L/SJfHqHkRa0T1Ln0wzTWbujKyoHhPimHqKq5cuQoZCYU8
VWchxFMY49rKp4kWCzvWIURPsWdm8He4WS4VlBb1BzFBEBC6XXjl7T9AdfV4
0KzPJhZvneEYIIQZC/JyySDYecAUPbu1K6xDWfSd1bMc4daVi+01xLhhM8rG
vMeDfWFMHxRnPe6oiz/+4uHel/1jkOuwJ52966DbL5BKYhRLAS1hQw2jgpgb
qJ9nIaHpZQcXrPCzdsqxTrqkGRdZwrINBQSI7fnP7HONGbaJOO8Hb9+oRvSr
2Ial+ZCRHJCdRePqHAY3ryml8it+FArihVMCniUzAl4zSePKi+8b6aoMu3Oz
T+zGvwefeKo1lsUEdlGgMpypw4Pq23SPxhu46yYxhlB46UvKc1FfjP09vZrW
pikssp1Nu1UBFoXZhzObKyos8fJ9bavgJSx+Mlxr0ooKh4me11bmJy/Eo9bu
1DOkgticdSGWYRAGE4AwhiTI+bdTsLQoWzhUbUB29AdkhetzEbse+4gImKeQ
gCDj38cJjCwn5ZZRDma9hPehsgL8ZOA1sJp9a+RFPTF2fK6/CHoXFNqMOyTb
QQdudFzApUsJdIuIgm0lDhfjLQJ3ZoteCkpl9NTEsQEa3sVucnipv4DMUmcK
XrC3xYIXNytGQ8HWFPtriN+Cp6wHfaWcefeALYYlTiy12rd1874Kiw4W8WSI
ai+/ANzT6xACBx2dt1jR5wQv/VsV8uzZvhUIAYRlMUShpXn8yU01XYiMLrfm
7kZPM6491kXSDHd5rWYVV0Ood1fXcpmITiNhC+M/LPVuhr2GmrL788hhilTJ
qVqlZGsX97w4ZPAUleN1ubO3V9gs1FBI3X3He6ydVsiBFBGqQ7eKJ/XHhgbj
4+DPkj/KsNfAh4WjpFCFjaJuiSCBdKrMlU+gpPzNQjMylrR++9FD9gC+w6/V
ZDcrMK5WIn2J1dQeGZQ+uwLuyMdrOrwt7oGv9A4BKPTrPAhyd6Jw+qf7E85c
3XepoDNyMhlnvcuyNJ02BbGirCZMDrs2nNATW5OQk1fBoukyOLW8PaOLsmWn
y6JYBE7iE06bJbCAfJd0uTkru48m5Mu6X3Q8teBDmBeEburJdbKijfYdBz9n
6O1fzFI4PhaI7Zloc/jYolPx1FMWvT8x7UkqvGbh5Q6jVrJckDD26BUCtq+e
C7SRwzxyMHl49QzmgJnFNmMEzlkWHHgzxdzBZjPkmG5PEhfbVCHGCWpicfAM
WDqCQKHiVxZxar3TYOl6+oEz29PrB1C5l+X/EiMZyempRQewwR4aKSIs78Mk
vlOH4hmtecX6IiYjUc3WHFCJQSkeBpT41f5KjlOcV1D2H+EkM+WU2I4d8Qjv
pf/zcUj461ikIp+bzrkejDNm7pTLfs/sb8/gRVNhvjzfaMpXebz8csBK0irA
MgLTyz4XbLdesiHpUZrtfaA6Z95CiHTzy5FmR1cyOBfinrcznXHQcRMKUUY0
hhdbcKll+oo9XTVPLyZwGo+oIlonYx8i4gY8ItsuISAtSLNgkdnGWXUme8Sc
BidD7KdPHA6sCfN5e7vUzA+3SjPTqKKfFjEqT6Jcu0HxTZiGmGWh/HXYAoGE
ex1x/V8J2FnodyWqGnEJklmDTznC1+cMrfKur9TFsQktsvm3Tx9OdEtt5I6H
a9EHM1U0N1QgDt0ZVP2f5nbBDEx5SE3McSIZ2xZJ1ufll3WKFB7ji2mpyXUU
GrHSOH2J465Q59Sd6YEPJv7y3m4wgysEYqqlzrQ4VK4+/d3/Q6/ZmodWHyHh
WxuH3ipWZzfmSrttPAkCBoBuzT6h+qC7kN+Bhs0WBML5c86mArv7WrqcD7W8
+jRPRK8QdqZxVpXaUVB3k2dKqa1vJtUppNVJIUZxhn1Tnq1SqrjXpktChGqp
NgWOkaJUkr+nFhfwG1JUW9g+r2vk7FpI5RVuXk1smBRNeupqqa9tUP2QzDMJ
M0d/nI06BuxSzTDnQ5BSav85MWyJiRai+dzT2jIFG120A81IWsGUYW/adX2Q
iwkVRtM4/KJZat2j9n0fViXfP8mAGPgm2tNtWJAFE9xZjD2G+sT7vmKhjpvt
H2gI1B/ZLHTM+bC/fEGQ883a58flUtxaO2LUsxbcDBkde50uAyKcgsl1Wguq
8e5MjrTfjubGPG28Pq6duOItTryZQAEoCtldFPHWq1XBLUXVjfqeru04umD3
FM3q+ZiUR6hT6QUHHWsjJtioCiIB5jqbK/yx49DztObvkU5VbgXKhsVKtRYB
KlizuXPKnmDvXyvfHvNxYCp24/Bbfz3eZxIPauhC/ZqSbasheSW4Xh66B4t5
Dy7XtwK2hHB9g3V+7o0YOOU3dwhq/HWeZlKXJqtsHubOxXm14ZjMatnI52ec
P5uZvGZVJrhPozP8GHYSLeeKl2M78x6EdFx0FfCXtIYjz/VkFCbSCAGK1Vpu
qlFsJPtkvwt99yY2LtdWd52+umZ7pK/Zh7WVMDmfY7OQTAP1znUkESvvZyF7
I+XEWQ7D1aOkigJddI2c7cpX+ynZTcvsb6b0E7ohITRr6tK921LhUoqX0oLa
iUN0i86ygmQY42xfWaMpM8pUiraUiA6OK/Wu+cBOwCeq2VGu07La8XGy1BV5
j/eoqZwyJclc5wofHs5IyOqMULRWuuApk2I2I0qQEs5mMb6zWmg9bQk/yRFU
IwQFg5Hf9EYnx7EXJgnEF12VZitABi7TM3mNtiYCA1xtSw+Yv364CKNhNFbE
Ss22BCWXs5f5v/QN97LTsh/IGZ8vEVrgHEnunEJJSdTT8kmkYmTACRtn0haS
2pBrO2PUcDI7IQMDu+cxRVNW5Vjww/Zi+SU9FuWBj0+yQZfKIlsxDDVyOIsg
j7iNxCYeiYfcCSQOcFwu3fzsCXJgOBjkACqIxw/5pWNEyCJ1fJM2BHeIrodx
GhIw6VfbOH7iUpBX52CgJC+lLMFkIG02OyRdmPexvfUjsMvgaVjNwsv3mni9
0MqoQfCw0yNV34xyFTiXlXsd3e/Ixz0KZcyRfzgk9u1IO/Q7xUdIta6pzv37
xQevEPp24dK/hiYaS+m/DOT8bQ141Tw6Zgfm9Bomh9jkRBPhMEj4kLe7XNYZ
E9agk2JHSQT704naTDyiBHRx17b4lVEsiNZJxr/zvD+0nV9JA6IDZiLTwQ4t
bUX941sBBph1yknP/H5oqTVJMOjmONQeRbYonVWMpofVh1c/nIW40oD8ki3J
alZXCeBycqaMxKjH3cgzHJ7kFpZ/nYNMOZElI3Puz3sxfFqWkuwGifqn8c/b
ucDLBQjILnEOlQiPLUWRHJ4Po9jp9G1GryJao9jq/7iJyuCfDShz3QX0d9oU
2UQXUQBz6GHiLprSGpO3+1uEsdklnHOc4B9LLiW9fA4bh3l4qTYRbuunkCs+
F4hVMLkyJIuPzycqHjeGghmd5X8Af9+R0zERnuem1ej9ACh2FOWALv0YsK43
vxUbBiudk51V6muWhNIkh5f/AFwxWSZcRZZAFml+R0w349wvIRRGUOfIO30b
SPBlSCXdXuWlccEOljLDJOIEHOk/X5QaWQYP2iFsCUUNWZ7oPyC8nDWB7nNF
5YqfNQqzIf62VaKd4NF7iiEKnhGIHcAb3Dx6VNL3qSwT09YpTrG8csblxjL8
Q8hBz/fktFdQoHZhuIH9fuBFsxueO6jJguYOFckqBy0cohwzOTRwIuPkHhfI
qM85h0F59/L+kuZXhUoG1THItnroGsfGC7evRb0sqUDvhR5Vh8auO/yVJmxa
DuABkDtrzVzSnls5avb5Amb/rvaxrNrYmsLbK7eowYpnZQwxInjs4L8FbyAH
yk082qV++7GEX1n4EFACAregYi5FM38hw9HgKqtPmUSf7OFnH65DOeYSvQXt
UIJu7qkjUni17b2tSNdDzkouJnUSASTNYucvqvJrzYpnI1S+FIyKnb1mZaTg
QNSd5ix40qBHzTae5LyDD6F4MYTQRm0v3C4fo9x1YVRlWdyR7cdgFDgNq7TS
YLw5OZ0fIS2E8vEV7szxx7FhIJJiyWkI+IZnXMIOdzBewIcDskPIg0SmcBPv
krehtBKeMRXqnCVnQQ4iwQ1xwk1XAPd00B2fb5cQ8//1Eh+ZuqIzYSRYPcIc
ukT8IMxB0OazbeYU+flKdu5MPRWebIj75jZkM0aSweie3lI5cR/Gr5rrXQqZ
cxt7NN/ieryWyORkJcVqy+D2KJ5frhR6ug19ICRQyWRIWZry62EOQx7aTClJ
keFhxAOwU1o74AwhmBqPGo1K3pCULvAt0yyb+JNCLBPYfJFtQSUgcXqtBTS8
G1E/JnJJaI2/IRqfNzth2gD7wy0Itb/GSDj9QpmxKOotLg1IKeDx3A4+cFo7
UxaUEw/ItJTjM9NaeiITVRuYyFtsXEmLZedCuywsG7wWiXCnIfYNm61/3QJa
FTNYgeA6lyhyIgY184iDzpEGjMQnc5aeYFDCUCTIrHkqi3Gt0eIJV/IUCHd8
QMyPahoKVVk0R8wFqElpO1/MBLXfEMoFnxwqGI/hFvXDDMuWt4PU7v1ZzAZJ
14DyI6EpbV3t6KbhgWyTA39BSu7Q4Hc7f2wriJnK/07M7VmZOZUb10pJl18N
OK7TjaNCPJjSHT04O4ic8DFHv7OEyvMzSf+Cmre24lYsEI8JiPOBi6mesr9U
4vzrTkUEySyxjGichx8PZWXwa80WLQARYEoEzJRbjpn/Ahpq2gFBd6TUVLCy
Y1eLMcQPdRgaup7AUoOLUMKfP14Pf1MvKBwdYIvH6ZbhHQrNR7902/R/J70h
GUKlmRuWswYBCp+TxOEvrphyR5842OYxQNxsgzcLJrKE+OMEUyY+FKwbR8l6
kv0R6Lbt88L3z/xDZJWB+6DULf5AXkXXT4pod/042cezOfDFPtJz992jdI8M
dU/hPyDasEVVnxzkS5vVXWHA5LHB2FW/bvqYRR1/KYtVMOdEtIk/2hUMub7D
lhUmI384jHZHmWaC3VXjbI5gMRvMM4k9TBR6PUpxGWUms2FuG12IFY5M25VW
YXQKBZZW2GmxKlhE8tpr5tU5HlfRILnFFbID0HqYxihOFjQrMO7vpEdi0ojB
9or8ueeNDy6t3BxsQc9jrIAKkmBlW6qVKTsfGWGChR0+5ayKAiy5orIHgr+C
8zoHw3vAqA9yHcF9D0mZ4cMX37qausaQMoqseSlIIYIRmnSgRHEty/+KBIRC
UUidQmBjNxHbX0iKN9Xj8EISBIAMkhq5i/Si72N4DlnOlPAgVY5EdYfL8O9K
4K3ZLcKtcqyOJ6C7WqJ5xMJAqqZlUBdGqSDclJ+OWI8hmZc6esiVAqGC/psW
HDMkPOS1nJNbBVlncdB9vd7cFRUBzEBXtgsMft5KR8nxbZLPp4XUhT0vEWlk
51I0X6VfCjQ58rXzj9bJDW0bq3P6nhpSpJgMmWo2fAANW/MlFdr/di+sMVa4
NtAFrCul23jOkToRBGdouxHwHywpUgNdmt8QoPSWGXHApoftCCErP0YXKI4J
5WwGG3Ukg2Ju5zgt2NXfIpIFWNKASCUmdN/qC5+E3ZioC7aO9u0Dxgh0UshA
G5/3NX8yfMvvFl9LzJ50NeDyi6YRg4oPntLSP0q7Sjw/9HJMmN4ORFr4cv7G
ILoUiP+edPZ6tiEB+MtAbdtfgg0CYRNMAUT5n/dZk8P7UQHOEMIW7QVOg0W9
eypU2Um1xt8f8N6upzlG9bTLvxW2gWh0KKmSbXHVwH4URw4nE/mg75rmp0yE
dvhLLddsJ8xc8/T5V4yjkarbRNDkJMCS2OAttqwmZPXJ0PqrwN52f91vwp14
wzgyp61ManpSwnq4JIeHFsRf61ErndaZqiNlhzDQNR2UcFLd6pUjFnuQEWZp
xRCLW8jpnfZsXmDCpCaxI+qEUNVm59bAYapLjBbtvf2Ifvfe8ifKvBcOxH8h
G2umtsfCkbUYTpp1FwX6VkeNsQbNlgJ9VeAH+qkpmCbE42ajqAKz5oBhWiKG
CXs7G++aaqBionPC10evjVFeb1hDt152vx7tjGZJdonyN9JDrPSn79mTKaWd
bUZHVYvqihRZ7V2AYDY/H/nspuFD6Fk83xoC9AIEA93quyLZHA8IwADDQ1M+
5IUBzMXe8qaSplQGW2rpR0iEFt1lL/XXYHoPNHUrxcGHZREhPLXWtmeettox
OrALy7Da/ODdQxO+zGamwDnmZCKHjDWKNK5LnTMl7ujNI9yQd5uSUdBgHyKR
9LPG2ThoKw8ffFUyyAsakLYlbMtbbzl+TtF5HtZb8sD43j/pOkfsib2Qn7ab
8a+SMZJfALOxLW0DFnYTp8Q1oZUZFrYgoGzMTTUXov+DeHh8B1XVNwzFolss
BkEhARZOA65N4XWGAHEZg+/cjjohoWpZo9DkxmKj9j193vfFKKKsm7+4w8vc
ScPJ4NWa2yPAzWuzrc13Ugapb0w3yLQlVpTMwRi9+GK80R4/SUC8AVQhu8Y7
BgcVfah1o3J5h0/MKkiy82Zy4J7G8k58+1s6rh+LqGU2HJUcEiALSSS+amzN
n1aGlqDSqCKG7khV/w0V9MlIn0JRjGPNUZb5rlXZbbPrpSK+7QwtyLr5dzMB
eSxvCAMkSYc4kdzw+BDp9qBu0UniCBucQqage6bG7VXEbZLM0GfbWYKIBIeG
deYjQ2O6kHACx1ri0f4ajh1Y+2qe9RWsdSn3DjUIRPxkMm5M4/72iAJjIOe5
dznvs36M0qT7vGicawHIsUnNnxHMkAND+VrRuCZq7hjuYPjoLugOBST2RLry
m64C6slB1lQ6ITKWz2BVhBjE4OBfxae3zTNyXrZaXsSgu1Y4x6JCD+P3KZAJ
cOIQ5TuOn7apoqZ2X3KL7CoW9cHVZhKhq0eCbOvdrdTV0J0SIfp5Fd+DOCh8
1eCMOgAV/EfMDWhlxsUw7Y1jHHgbLlw7Sm5zmj8Dy4O0Fg5F/9PrE5TtnY79
T10TCRauqWbetyNr4ISor9BjM5+M1zyOxDrGm5GRIoAVm1wTuOvGRQaI0Dpx
i7rnm0W1AxYP16cvDAj6LvK8g2elUVTNud/0MC5WvPnwpYyQtGBuaUmTp5Ep
m4iJXf0r+VNFGa72iFjsCyhCKwGMBsKIgNs4HsqL/Wnbkxl9wXQzVaR7/YMA
fxUHCYPVSGr5aSNQZClfsok3ZTOkmlkizO+LmGDl+qn+1H2qP+gGOwnfNkbN
JI/OH//HOCitiJnXeJ/yGiyKkOQXhswR98Yz36NyamWdpsBS9zgqbSqD4KJ4
VcQdzR7h0jAcNFNh0U5cvRmNsxDE93MMS0Q/BR8OLojYjULb+hLJEOgMjuej
6edjkKTYtGudMpIZ9gbYm2KEsLY1qtE392DGJD56n8VfL2gQ9v0CHw7XuodQ
Sn3dN/w5udx0ebqvy04hatBPAiJD3U+qSlUl3zG8KHvGCh5MxXQm7ykxO5Ii
zq7Vzib02Nv8q/s28QXd6h/+G6SKgTF+FZczAWRC8o4JRRwJv3ErmsglC6b+
H3Il9UmKJzQhA7Y1UH4chP8rEA56I8bSmJHhUlrcCRi5dqjC6DhI/emWIJBW
LG+Pa26GfNuyTDxiBJWvSeCrs8IhMDupkIg2kn0XB2IYEAHPWuWso4rS+jBu
qILMTYc08trZfZBCow/Wo3SaISUb1A2pQXbily62PR/oF6FD58IKEHDz/YWf
G6oJegi4ZoOcPERf+jCzV4Rh8GKT13FIZBiP2is+u9lqqM1FKqRU87zDB+1n
XZan/Oi3blJV3eVBcP8dnji9v60cdFigMc4/Cw63tAyVCRVHFuxEehxn+8xs
O/sQRO9LaJU65ruq8BvRj3DgvFQ853sROocbwNEtvYTk3NOCjQx27nVER+mE
K3XVEIPI2l9wihAVrAKeoVzQH/mXOJllvdWdwEBUlx7KGG8eUhBSGnOUutz3
qpmAUXG8deHSoNTzN8aUAf3jDdgrgOXU/I/9HSvoqJsd82KoszDdC4rWylHi
cJ+09ZgLgGjiT5c/xuV+EC5qF0DuZmKwvkpvRh/ma95bUTnXtK27Cpwm+4ax
y3N729xIsK6/O05RwTDm65QrfbRoaBXl4+jCT3ILScqIf/FFpTr5KPTzuJuH
8o4pHqU1xsDV1jofdSZT3bfCft0L5Svzi0m+O1QAQnrYT8klWHuHQdX/6zBS
VeXUWTK+PK+CXeA2a4n5tJ5r6/7wRutug36jx0Xd+oP/l+jw1eACkhcFNOwG
+3XSWtBlzThnysDtrRGUpWYT2IRLDYvmZ1GN3vWwg8fg/nN0YodC2rsVijCt
+HbWQ34JKGHUJ1tUdMGZEgLlRY0lb6JsI2mC/RvuCch7zC/g90cNOrxGtpRI
Zh+soF1Kqpjw2OGwqDFGDlnCzN1eaTCmydpNaKcy/hpXeY4nb9qXrw+pLOSc
/QXnt1SAE1+TEuXBiaDSagLqCl8pKhY85Vy5H/XJc6N40vRSd5f5dAxus91p
UWo60RuqOkkzSm3uFhNIuLpMBCIX1aEWywmqP0blYEyodWxj0gqyrbikZ4p9
pzzXUeqseUVil0LFSzF+d9RMrm+kipgFlD0DRPHMTj06vRAem56iizGXjfK9
KIoOlpzO4QiEUUti2Kt6JUUm2SUxhxV/eWSmmTMunVtz/uRSnIyuvr8M1rMU
i21GWpXb5TJEULwFyo5f7cm80g60eIc/KYRn5/0ffxpJfYKOKamowx2rv4/A
LIgSEUWLpwz79x8BeUUs80j25O13sY6IcNz3r9mjsD+Ci2dNpkFDlN85q46R
ShF8wrijFXWUnSSNoQD2lGVX3J5aWWUQx06aOyBSOT0Eqq1gl6zLhx9W7P9E
ex2DlWTxNcu6oxCKJErHVFg3k0BMTfJw6ClEQJs0CAI03h6l7RuFWJ0A3PPd
Vf1YL7mHVC3LX4ReFwjsmaPGG4RphqZkekXNsZhgFmTlq1G3RCL+JuWir8w5
YPRzCHlEJO7ltLXW/5GQB8SQqnlYoqKX6dLjyIxZfv3vBpaif2tlbLRKuMVj
RNQYZQxIzSqkiy47RFsSOrzvV2GArW2FpIRajcIFtmoQDLhls/02CrPV0iQI
TDGObvm+fDlmcJQIx8+00u05baW8ANB+6cdAmPjoGJ2xV3Db24qeNQ4Qr/IY
/gDehGkP1CyKcrpynJQ9m05LPhzgjvFfLOaxr1NXWcTdNGHDQbChusZLF/27
LWT9C73NdHhpMX845xR1ZcNk75K/yq++XNmJyy6h02muQOWvuDOM0vCy9zS9
+RquV6N6dk7hqItlePJY2TwKhELNGPeMGFvYIPWPcqUFrmYOZ85Ki2SSr4u3
6huBnOZqbqzNOHxihwFffqXzH7YrAS3pPXPeL9Sd8aqmMXA29WdQTFwHPZ4s
w95HoEI/lQ2oMRs4i92TN7meg15bqXrH1jYA0vPQVHRkuoam4DIfLY8KA2Rg
8oMbaKxJW/DHcJ1ZGZZoPsa2npCqqpKLpXOiV7eflAYMK4ED5fzzuXqXObfR
gb1+VgBTSnj3KeixbvI+TAnUSpf0jTJIhwMSnpVRV/9oqjKuy2Y/KEb3IvwA
tWP3YY2Qh7rX2ijS7NnUWvZ+BhosLUGLqu6I0y+A/K8djStxnzP+s9DSeuLT
UOi3MLCtFE343GvB7rFDElR1GGeY8BzJp3qOOseUP2BuVlAWgeZDhWE4//t2
p+NUNVC+ug3jml+2JsRNxUWR7vtdK5V/RDyeu8ge1dq1LaqDLkFzLBUc6o3q
IcGZSPOn19OjKzRjQN21criKtthPwqs9SuABltoQuKqyCovCYv0daAw2HVa/
o/Fh+26+fej7siktBxegFDlXFU5034n5RFiQnsmDWAIGMVmI+g4sSzAdAAoY
U4Ie3qcNza22tBmZOBpsE4Fq+JxNYJPAukWiOO/Dm8fiG43kHRJjiM+4gBbK
3TRPz4RDd2n5Mk1jedt2tIy26qkIO1TL+k3TCplNvxxD7HQgsKaqECneSgK4
+vwH8I7AvBls4A8zUc1NwZJj4X/Gu3q53PN7R8FhuHMnWvNA2aVKbQd/PZZC
ls0cENixQzps+LzdTZ6N4lC1eKLLtjxN70zK4ZDSsHot9OYuQMM5HEcbNCTx
hoRj8AsELYltakBXLJVjygdIsYntgC826LGEHL4EGobYtajoBRYrU8C4MZvA
Xcfc5XyVrTSCOYuuNajAm49yvU+7T0WkK33RfrQEwWt6hW9THUKrvtXQZPnM
NJJ18Bv2SVIgT99qMgCNm+MigqPOCITFP9NNNBzWZpQIImrihfYKW8jyxl+2
I5OBjSmMrX2ICK+OKaEsKW+T8lxpBmiaPwL3qtoGhwfz3sO2E58smhoJvYJD
NUIcEDju/5xSoarACt4iviskzBApG0GrG79cvKIDY0lCeH+4aTotedpfmRJp
rPxb04KvHL1O8f2sCLvhlbBVXxZjVHhIf0w3gfFe6CGl3RFwbmyt5CIGTsy+
HQEHI9DDjkYL1BJ40wOKCn2oGjDoiureJ8Q5B9VLtXoOlL6Ui2ibrZDXP5NA
JQlFcTYr6VwERFBfpegG5YxJz9VUdlTliolJcQTjKcFysdbUzmC43orSm8+s
pdU+ENvPtzARCD25VVihNg4AKlAh33+yI6RCQHHsZtd00CLI6ojXANas3nSE
O2C046LtsTHWjHxrHHr21OhS+1Ozta/AB09FWdSHzEyq3m1jQt1E+XriLPtD
HaSiWTJ5dKZinyeyOczrjkl8WX4xTF5udy6li/J4vrSDtn74vHI4mqKKmRiJ
mLzHYGt5OJP4Nw5vLBZ6abN2NcBs0Kw/84mSL24sxspI1+brEMkTwVNsCtmk
9nSbfL7VpUVz4B1SYAGmgnr2jfoLchIxKDL2piNr5fkzMEkcBGJO1njrHl6p
ZGd2qd3IO6CQZnIzKrWrdYQL+qghhABwu8ndDlFvo1fwXsqQtvXEGZMSk5Y9
xvHIr/dQY3hBWXaFtwcHu6SGbpfQb1qu2txbiQhukIDmwVCi3CWSIVS8gO8N
NVoWLkFH00jrmAdXIk3AjiIC4aY2pf+rP86e3Xyfzt2th4l2gCj6Yhusgtfg
/QI1TYEaigCPINNZq5SNte0Cy0NBfWXys9qdllbdPWevXZ6D22GoagqYAEPf
1qBU2IU63pUkNrqgdrbdskuodx3+ZIrFeh0xbp5lDrquUm3AhyVvgKQTWvIp
gqFb9Mr6FMausEYDHpUvnoM2L7R3Lmo67MT0+sfM1p5yDwUTftYkDvpquRUS
sRfUllVDndWufn5GJAlZZzdkIfUwggESfXK0T5kH/SjAh+K0TiJXKjvBA0A3
+rI+Nt0zkiqJBv3iBwkKtgq22tLxlgBlWgTmChz3Ssw8mC+Hh/72CxP6vbAL
eH0XEjIUfVFVVGplvhv8NuZl/d6BkAi/beY0m54/OtCjFPamVR73B5O6ZzgM
DbQFrbPV9JRmYwT6oDOhKxbQUrTYvy8lXp3Vk03n5LPaaiEU1rpWVtsyc6p5
OvSqZRxTIypqutUGYdSi0QafAoX0N8wabrSAUj/PHip4uR4jJVCzyvTqvi25
R069ozgE8WiyRIAYE71Wkahi0wHLxRrNCal40LMD2RL6yw29voIDBqOX2cbD
+uyGyEkZkcvCgaVL/Duj9lnQIdD5EztMhoVCCe6CFzP5USjB3TuKu1yW3tPB
aHmhuJRQCHYNT0BzvW2++uAOVaZZrQ/rsxN7abi8ndap2vDx1gMyln1qpKVr
r1xslLV/sTxTAIoM8dgF31yidckksgscoSXeYjOWJVvMIxifYqM7tjVamjy7
SyzWyTOSiFg+ORyFQhkWo9smoJ6qWzqwNi2zjoVl2BY8bvHBZJSwcsvNzgSO
9kceWIpqNhQBI+kqaV+PyICvoRjakraMqlcqCCNgmoJFRUFf9cSr39tGBpu+
kWBVgK01qTksgjP71+7AFepViewz5tHBh53P3YIWpP4S0q0RaR7bhwfT3QPd
RSSSHh4mu1NDhFI/qZUGwDtCR9DsW184D4WNdU8yB3G74ZY5O23MqRfOsgqo
O5Gx8u/7xczLMERy5+9hU2CrKJ27PAMfCIiLmClaFcniDBQlxY9ZgNeAZWNf
0AlDud0ReKC8njTtaURLmXYkY7eTaGGB9+r8w/s0SqPurHoQCBzto8NpSJ64
SpZy/OJW/kJlApur+P6LGM6S9kmwfL2sP2FYLX9h5WWAjR673zBHsXMxLtey
Ktc8ZHLQToAWTgWhGBMu8F4fS0rhUyhMpac4pPCKgY57toIbQEe8TODgJNq+
cOCjvjlxWgildqKVtvWYaLUGrzmTw2Q4fw78NJsugk+obkpMAIu6NA1jWN6v
jmVfHmYi0U/kNbz1M3Fr6YJFx2oG8cMXF519ZXKaocb4VQBaP9IoLRZXvXJe
P+zybZvvl31iB0quNkJ9faU9+wM7Rq87/l8fWjH2wXd/gihyylq7+3Gj6xNw
OuOcCXZSI6rUUqvymYY+U3VbMIzOTvMU9lEwekUOoEA7qOoH/Eso/jk+unoU
r9JVjR19MCqs9Y4C1F5aM9S0CjNt8XW+hR2XTD3tQJ8E1HrtQKtRvu+1Og1G
2pJ8qVSNdgRGTMPoLOjJPFtnfQl/lgqS9Nu8Q3oTQEHLBSFwV5AJRI1brMvH
JsvuWwSimuQ42O+gQVmRtSZ7qCIbxnTxGbKKgXmIReE82HK8Y4oyix5VoTcE
yoicAImcUHn3H3oeETp7AGl3Q0vRtBlfG1DJWHlu5P5P0eP4zGca+qJlk0sR
6h5F/O4QwkakFpoPqd+2JY44bkM/r4gUYoiwAqVgDEdGzzXb9pEs77TwVf9+
d0ezR6TiACGpnjKkfRkosVdLNjjvVhrrcixDN99rVOcKdyN6RUlC+IY1Qr/7
YlfhgWHc0CZfge/4yHOm0dN6mWoEZyythJtVFY+58kT/0TR+44k/pSaB9/pj
Wpaz9vpB5cnupRh6LuO2ZFtp50WtH0fuVgCE7lKxUjCJaLZ1FiuB3ou6m8zH
e0Pj6966khSJM2bRsRICQa7/d6ai+c7JbJNj14KPMwhgD14GN7EOYw7Aso6s
fMcHeVIDUfcsg/hv51UlgeQ9CAd9LcHf5qcO4/wyhoNAuyNZ6YMB9348ZKMO
NA9/n55OGKY+0g7gU3z2gEiM7LIB1ixNWRcSnKOmDtqRnIW9miQWKJhzqHaz
qmhj7iFPv/ittFuX6s0vbThl1h5vrogS/ZQp5s6bcgcR3NPyYSgQOhFHDstI
V+yxAdyiq1yRLcVSUJvZd6wHGDAcCUTylX1QSVUDCafgK1atbUDw5t9dPnM1
XFQQXWf2vCa+fMarXlFpw3TulFB1usBTzFx3uStwWY8nLmlyvlcYh2WaLpKm
Q7oIqL8TXfn1drewCZGXWAjWfdAR2N9TsO5IWidHTXHjeegTZL0LAxptQ3DH
hydHwLsoDjuVaNh9VlSW/w1UAcZ0foJpQMqwRl9jVCFe9NE4zlFC9/3srtXI
wzMFBGpwHRK/OMX1xqufePsKBxlFJvx4lp2lv+68u7A9sKdIxAn3+94izu3y
9urL+D0twSCFiHlW/qLvVqmpU3iEeXHrKqjJK+atcDoON5scpWKYIobm6uvm
uh2JoH4WN97mCtif87sCOu1k7sVYLSixTxgxc21ZM8AJy/qQHASireYDfHPN
cEDj2Fmyd/KWwYjWeOKwDLsCTW9ws1245PX2bqroukBd8N/LseqK3XCbW4hO
DePFW9NxbLl21uZbeENnl8LlMlhnG3psfAHottKLprTRv0U1FthsFvYSBEVQ
NF5aYG7wmVNj3Vz+vxWoS4CGhv6eAgRedTew3FUYoGzcF6TfJfaoLthrp8c5
fbRGD/uJjBcWZKqroVKeTZ/G6eXF+FiWWpJxD0lpYt150WLCLOnXqgCKW1XO
HcFAAfV5eTDOApuJ7yKLMWRimkblfMTqkK5c/+pVpPUptFXMv7etJHSnhdOW
ejoLoEqgL3N5/HTEQ2d0x8gfOLdXyk4R/6xScH/2xrfZX+hCMA/HWc8M1MYf
2qF9KaWRPrQRGpE4rgmHWB21EuRmU/wJFYagxZOxXMh/HTV3TvInr0Aw3YbG
kQV5r0YqcN31bXEyLXPWxByg5e2grCMrz+GAUAk/mI906IXF/enfLeVS+nCf
56LLMc54LXfy89ci5jcA4/Orc2bTAl3lCqJb3m6r/UgnnEubBF7DUVDariWv
LT5NrBG9jouG15/NDT3HpwGMPFMyHN1IN/294RFGxSSYWb9PCibqJPzejT/6
oSxdpT0WMPiZKXHGcYfSXWCj7xsZ6Q6fvNQmYH/vM9AYZUtMms0ZFytRgFSn
eBEDr5wd3LinxNB4Q6s3hyeFmhk/d/j+kgw6VVuW9N1o86K2H5SWUvwMDSRN
z1Bn4ugyX+o87T+7ih1if3i6GWVMLvCLTDtGfjbfZ4nGZ/xPZkTqdqasvows
v5N5jhHPLjHa1UaUZ00l7d/yDcXIhtQAxRJJg9pffqSuoHcQ+/yAyuFuPWY/
MRAnZTci4VHtawt1ra9pRkKLej0Enzusr+EBAiV+0Pgr31/5e6texKVA69Qb
+AGxItfmXjp5wM9P4mdSEguAa8kRLMb1qT9islNIxxSBP8bCZRaaVZDLcu/v
Kq4BIQ7oi+vJzwYSKl0WxVTawc7oXJ52g9fAwln4IbgJfEQ0Un6uwOrjKCmy
Xlj+FVtyaIZ5r6d9ig8PcAJ5pA8R7sRk17cmSvuGnQzM6UdeYc8Ac6N3/QRy
UDBZpRCrudbE6LWGByzFnj2vQEjQxlxpX7wd5msnny0oomfMGAq64sPGboxT
LX/7K1PXZYcshMPUIYRLc+3LyW7Sm2UA6yWr9gwAuaYr/22nt+6i1UFQKtqo
9bFgKXV2IE7HHN/QNQhDIJni+9xhNsR+KbhjwS/Y23/XyCqEpEtaazKd9Mzn
gFS2Ol9tDZMqN6oa64iKPxFyCVG9u4P+9WcDmg3wqqBkQP4j459GAkHZ1tK0
CCTc2IkZ0xnFKpTQhbApXZb/ajoCMfufLRXwzv/XUKIu0zLp1Zs6t9ZgPvel
CFuOfqK1V64uTjbMXdba/pLgC3qeVm/hq3r9vqCljSzfyfFz8FUdNWLVWD5+
ahMTFNO9q6c06hKLeWvIm2Ui7i8YSaLQuzgIWCEVem9UuxG2dm5cJean1J1W
l+nQWLCzjF8ySg69S7SH0pGBeK3cIAR5T4nvhyhKt+3FU/4HkaNNXHqN0lw0
UA/LhuR0g6V/MSITCBlD0ONGHBRQxqDLqnSXnSTEpiSuBh+9iQSEwpxJmjsx
fWKfgsAaAuNXc1wzg5GPbepIlYD1jjMgNoB4Ai1gkGRqpxVksHEn/7/bx1FC
e4r9R6041ep/2tKJppGkSz1mBYEOKoBzNJTaM/Aj5KEtXwvofk7R3wXwdHYM
bV+ArJtiNB5wYkDCrs3IgAYUCr+aqsjj/W7h/IFHh/nHdtZSnkrlBInp1iP8
c4Hspdqcr8dTeW0dxSKYodT6nlqxeY2xvecw1Lx0SJNwUlBk/qehg2jkYZM0
7iBSKxbgz9b1yan+L0Q2BjJUr26UF0Fpu1bC72Adin2ekElX564iYtdHp1Bb
J7EL7qvUhx2xqrqyAJn4GHb1MPE73PMgBw7NqM6V5EpZoVOV6h9P/NegaeWw
yd4AP08mYZpAt9ya6yNebyKm9GmN4+ZM9JIPb/wtt8RsWM6cfRpHKIuG83wK
SZ9Gc16VQX7vt/SqCDDQig4HiBnuQ7XcN8YZHgADhhqWP4kfBbFwsvSMIQyR
qJI+Xy9OyxS1ZyVBvaYZT0IPGIEKqzGfM/yZ9sWWqLLExudRNCXBw4Irv6Hi
sWTtuK9mEHxrFfO6OMqJhtQi4xl/kZeffQs/5mA6L63foa7uOrKdaZIBvmNk
uNQcHEPqKYBU+e6mUx7ZOvw8XfMXhE83mns7RPpdv9/V+OiB39CKsdbA4ECV
i6YwO5njZwWWB4m1W9chs4BvtsLlSSRLNiOFuRr/f8vT7A4O/rH4STFpVrpT
eNXNLGQNiCX/F8JgF8zCBi/0Rj0ULiOSuRO0Idev22ocWehhc8UWVkfmBwVZ
5C0lvCA7cY2rHuoertmOGdzce3ARviwhAEEacIB9cqtJ/1uiyjudOhnn3iYt
IRSMXGP9r4BYfBYQajNvWZP+aUJB2dFKyfQQRN3mmFyVyKQYKrrU+RhuvBH9
lXvNBK49CkwmR09gL7sB1GMM12IKoe/Gfxrx6p7Q2B2HGQS+WBkY9BLPe/y0
rc/RTKeKEz1n2ppborMZhw4yBK8R6Xv9ATiPADO+o3FZ80Q7LT286T1NCD3V
pPSS0qadz1FzyyhWWsExt3uCgL+CnP9dzz1ik+pVYObhrhglEsgG0dnxdlZm
Jgjlw9op/VtpFXW3Eat3IfNhc2bKq43PojoH0Ag0uvX2XKowj5rCXyuJy5x6
GFVZaLZRnb+Mckn+4uiGOBv92El6qW8FXk+JThFKdxJP8h8Zx8YuCiv8OFNH
LwuKD9hww+dxe+9uuzzIlOCI4e2i3ydbFORU8I28wZPYB+GfJn6/mBi0UQV5
ENNr4wjbAPSOYdiXnO1ckpclUR+sHYz/aEu0C2w2Nn/sodUwSUPiP1s2n0Rn
f+JGVb4aPPvkhTp3FZcRBapKxPaOAsiopReGHRbv673Hwo3oBtezUOAHYe59
GR4kLhslBKQbrABOGaAw558rSfTgxarjHZM/WNZgGOY6V84yhHZbtN9UYdaB
9cpVwgg9KD1sLwFVvmJd/ziTNLtq331e7gd9I3itwtCBLYIYy642Z6T4jZvz
ELPUlQ32713U9wv5PmTFzmzfw64Wb2gb79XmrEbfhu+CgJH/bpgzBVKC+T0y
QVIcS55+xKcWgxBjLDEajAwTX3RBjy2aSy9NZUCXpUcMsqCWPyklKj+2zI5Y
0yZEIoU6aDsNS5xmw5c84T215aXldPYfchIj7Z3do72wg6+QHMhF0ch3IZGe
6LOOA2wnGefVt9KWnzJhmIPwpd56gAqLtFPrjqGvM2pwMKd1tkRKrYZO8aO/
phXvBptC2WXdyMjLpuzdNfi7xey01uVkoIAFuLOrGA0bMSAX0GpV7QXqfXMI
CU1luaJrIkIimwpCZ+h5BozIyOnKFGnoP3AZ2lQ0GQj4sD3wuojk7QPwIPDu
n9RIh7Wti7Pvj4ABOZr7yz+6gXSw1Rcp2tJD1Qja1IFWSFl5uAJlMbTnPMhG
AFyrUgSxTQA9lU4tP/XeJicl5gV9uDg84m66Hnm79DGEFkqFaeSG0CndWzvT
aJ4N3Q8otNqRmp5ys1DucG7J1nUNM8QMjMzjMjhi1uWJw9i8FCX866fExVib
jufOQsQhRtl/rGZRd2I8sQuqHdbXEPdK7Bakgvoko/hSaqEcuOv7DM8NNnp0
WeQinAtwKz50LotUy/H1/7+8AtPc2l//kw1JvTDHuJ8l7pPMUEz5GE1CDmY5
bZXwCvbgRZqvMoPfqa8XnSCqVjTuLrpzFdVglC/QLyQjWjsAtDSd301Il0uj
ryaNP6T+N90pMTI6H2sQuj6ZcWtVnYL2Z+OjacZrM33QfSzpgeUxrtDj6J3q
x0/AQp2z3hgkkzNS3MY2dBCvk2kwQkuY6j9R+0yaekk97FcRRnIauGOZMjbO
I3M75i+DhRhpAYzd5/sOkYnzvQF1+PfKQrx9WweM6M5aWas7223BnENMGuus
UG9NEGGlXD5st0XdJcFAB1U7yLxiU3qNuDyr7UZvQUc/Z0H2+GveiXy6bzxR
ge49SQuZiHqdx+J0k/oBuW/MY3Ko26TrxCtucagXOdYtGqvDANvhmXStPKzd
4x5ClslSaf5HVvoCTIDjCAHG8hs4cbhQhxaekbHpygsLQwo5a06wF4fEu40k
jw4okT5hr8gagBe/foqDT4DZ8v0MbAxawunrXdEYcj/CkhmDAXk97eSmJB/d
sNiK97D9Eig/IrabyFGkXvMXucpEWGf4gVsfZuQyGdr+z5awf3ifW9TV/Yuv
r8D2srv37aFgspIDdyTt4I6DQXQ3HeyIAro8pxLpm2GGRerA3ePYiAofRl2H
QP6nC/+U+W/3kGlbAJtfsDFdHrsrweW9BwyWEsb2jhqeP3VeQa7BgMlhc6pg
ej6He0wVSbgsrWHkFGeFgKwff4osF52XwQqO66wKvfsgKOmUWk2GTgNdkgKe
yspQaUJ3KgpNjn3MJcCHoJT7nAmUIMa/bmhtclcllBXWRYlJld2XEWQAdpX1
m+em3VNYKj2Xv0T1lQdLHZngBZQ4OZ2mxkE1/pHyWxO5Le3dcfz6sP/B0DKA
//lzoX3zXwVoTTEEb2IAMpjhR3RcWYvNuvaZPZgxiOraaSKy6fh5UdkjTQqP
v9ogdeMvBadxdEWK4tBpcrmWCLrXCxy2aVR2vfV/m97mgAisHa7/V3+MlJmy
88Y7ifXsHJCRvXjGXjBf6AyX6lpmFSS6qL/ygF9jOt5R6uD6QKeUB34iLQjC
cx1PYnY2O56miuZs3S1tb5YML1d9aaRKj2yN4eewow/lbUO08dzeKYp7KZUN
i0DFClHDK2dywbzCav/LhtEszzRGtwSW6r1sIzeA2Kw98zaiVEFMNqaIFAUE
b7aXBkdAgsdgS82TtKDvZ22nlNwDhf9+A8YSYwOqs9E3qcR/S3x+ulKuqojw
RljeCF4jbKFrKxIxa4poQlkz8+/H2SklW2g3Swbvyn9foNLeiQzM6OYuTkIq
utzQIowVwFGrs7qfXEownH7po6laZy4WcWThypbWTDJk0JVqCldF4d7BO5wb
LBIKWhHUGG8dPdrZxpHZrfYN+SycGlmxE1+/Ab03LECiCKaxMw9N2VPYjLQv
Y1KKtaPmXgSCCV1RPpCgAsfI19r1dq6QV63XJcyUY53CNu+QKkq7FSpOhFWg
wvJK5HhG82XRW94f/Jn9AfmY2NJnC/Ws0K114wTFr+dttoaFurwgBZKg8sGo
boXxIazjDi81jTYEQAMX4MLhV5Mv6kELXx9u2Yx7FJfmCSibd65Lb98Nl6Zb
lSH9rx743fElamhl0bjw8h1UBIJ1IO5H2toFr70QX7KAWBmEnThzp8gmJabh
ajuzOgFtSzVuufTjBBB9cYWB2DKzxXxiisocLflwetdWQs2A2eLQaZNrwCgP
0H1cOnSSvZMnY2EoX1c6qgqNAyPpYmx2t785zDMe9gsBe+PNYHpXCB60CtTF
klTvgNkhqou5Zqij+s0DJItDs+aBbNX+MLoYk0ptyNwpoT9tXTfeYE3/1rhv
xdNQ5YC7+eelPxQcJOmNniCrY8wlw/zrVv6kWaKd5BN43oKJGPSlIJim26+g
trM4Il+hZFqNwVN94TBDZz6dqOfhJC2smSQG6I6L8UfqowDAHZhFvU7itErT
Su3NgfHtusnZ4kc7vIIPXv563WZ03Ilt44pKHa6WuR+WkmRi/ITNiCkiO/5c
wHkkAHh4zPhewNEn3xNkKL6+CPmY9vkbs0zFzYO/Gyw/2qCpnle5dL+Ri4N5
xtx1kZGaPOmKCZrzPvJyScEKyu9Za0iKqVDAgyYmzLiikpRivBXDoYNDB5WL
aqxfvpYwM4VlH/MqOH4+2SrE/53ay/0e1U282aXcIJv6+joo5SXJfDOaVEjr
XW8TDau5bbNNLE25tGp1+2cqEnikHjCxGKVkFEi7v5QULL3QAOaX1REh8qHb
w70SWyn1KRILF6ghpGroAuG2qhBK8CxYusUOkEEOSA34c1v2/lU4W3uxfY68
Ta/bvFQ6UBCiYVd4u39F9f92e2+dN++qIORD6NMeMxGq16Aa8b4Q26VvqYxw
KU4mfN+HyEN5GZ8facA2f0f+6rvc40wFg0Y1mUqHuH4t7UkESNZf3qtQazyT
d7mh0ryc5C0xPk7WVHNOPKpElhPWYMT+XP03nHKnm3cNGitdrkhugPZ/E4jL
kFZntWxZYmTOGyhUyK6OXOnuuosPAxjWxHiimP8qYla/CnqZaIh3V+8zaRjP
YcJXkUDG7jiM7s4knRjte68ccRIs+VvySQcl0MUMmYXWuR30QZVlozOzzEwT
kEFj+EikOGhP0StIWW6EDfjvh8ZujDrAHQKInjveVuweWu4/tCyuZrqmpNog
67qdkDmQDWSYdiX55dxviex3eXoeg/RUPHYiqC/QnjF18lgYS+U1TEVHDI9A
MPJua9W6XrVYxkEtJtOswQGPR1uq5VmyH34M5Q6BUhP9nOLpkQK86+1rXIYQ
GT5G5c6KyRUJjsSUW2JwvsDK10F2EmwSLkgPv33B6bFvZ07k/P2526eDYKIr
6KwL4py9j3bsOuQb+7rl5US7IGQYYPrnQS4mTNVLd2rN0DJ5tQSaQlOcH6ea
waco/nnJ6L9YIOfceijqD3qVrjaXVbmO+m17vSwjl+5fJ26WgLYiNv4YPwEY
6YKhzoz0v++pTFJWn9RHNAVEwIxZJTueSSDYMestyMa/LSU3/yO4VyYUiI/+
g2+QuVnmpmeMJ32Lb+j2fUklM4OwqFrTnrKeBwqxpU/cM4koZxN3hFra6lv5
WAm7bgMgIA4ru74qlGCaq6uO6Bil47Ld3l9pVvCDoIF3VgKxFhnQC8cILiDK
tq1f6u93e4NgG1e8RMMdd6oQ5tPqAg3poSzSt3olB1mjLUL4l5QqzAyy8Lvm
wOr8y1+pXwfQdN0rrFpMDxAEjhcsrSKLSSEkqhcIidbSo2cjdVyDHlulw44b
WFr6JXy59JXkWYxUV38lGZvowGkJl9kWNCKQNY5hSx+6Nm6jxnoN/ckq2xNY
MvMPB6TrA4gmjyBtXdXN2PniZxOkoc1xgqQvwgff1pY+cd/Phnw73f7ZtTAG
UFnIqYNVGbYzha4PigjQ9pAxkJLTux752a1UW382Q8vCGBpXLWe2iVEbagOD
vJxhD5ENcL44M07rrVzx5f++YOgaU8CPCQH8SrTaDF7eg8BjqyVQxa5mOBs9
PzvVdFLp+T6PJsEdlRu920ssxsmjv9ZWx5GavYCGFPRO4ltjg61jeHe1wIO7
KxOQwUkcvjYcqrfMuVfb6bujApi09M0IEHEdk+gVc7xMgycoj0Mqaxi4Wiaq
9DvvbkarbdQPAxKVrqwb3tL3xxTl6O1LL9FGRKjy/ld/Q/VxCGsFre9Fewos
9CoVsiUhLiWfbL3r3zFb6BPHAFgOREUr3oCgN8H0MFM0kLciUKPH4mJjpQD/
B26KbnGUTkVoAC00cInYaotoZN45LWOzaGXVWTZPSp+vLE5CwS+9xyWyDnRp
bJMiJZg58+PB4ukFwxX4ik4ZxErHPdSS6RjfUZdUMm8Zrwo0aueiPa2CJ8cG
3REtymPbYY1Qsib5TzWiCOyoc1dEyl+7gsL0tvtvL518QYJMPWWXy+v/oi3+
T7GqY65V63y52vwoxFE1gs1sfajz27RDKIpvY5Aul+wBH2q29HLZpCK5RSHn
CLrycMLnNBPWA5hERc4LJFSlop63D5i/oI75M5SZAsBIl8fJV7lsxteaxqfc
1S2qnuu59GAd4NjKZD6CJNLWxOrE7nAZ9OBRhpLXlyONIW8A/k6W8J65FIAm
W7EF+phyKIWHbKLS5kowJoJa6uwyIvVhakfHCj2xRn48Cds33reye6ZOYLwm
tgdpaDEmw0LxPYh4ZWa7vtzEvH4IsSpSoBVapLxqMYiGtnnkmsZRMco/J45q
HwqoDr0L7JaWxMTgTrSxXwMHsuhkwDX2TTY15WrQV5MMyYdNefOiEjdJSEmX
mBjLdTPKm0pirkjJ+B8YZDR+gA0bcJk2guWz6+l3CDfk5ndr7sSVtTjiFt4v
VUZz2fqGXKsfq/AHTlEoYgMXJQbcVe4Ad8HRSJZfrMoqCHx3EMAaA++62f6m
4MXBDqIzqOz47NqzBOBvB3+WC8uJ9TvRD8Ug/9Ga1uWocmnq9gBQc5hEAPEb
AnVCjilZ5x/qY0VlLgfCs5NJmD3fszW+oGJhHSD9+bsvyWN6JUe00wTvI2ui
5Drs+ZRfqHqVfmmtEjsZ1ib5htMVA/BsXb24GBJa0dZvWLVoOjBTMNkxHtYv
KFlhyAgS8nITOhQS3L8IEg6uQErKtP0mWxHWAA+B6OSsF1SIC58PMzAQqOZv
jcCBOr2lEEdjGGjQrKUS4noqDZilsxM0+bD9AbTMiKt4vjnvIb9luH5vBT1c
qG9ZPelRryWJU0IGuCJrkj0m3Pq93mq7CIMvh7XtnmUGvU12yK3pmKxx/KHG
P2JMmNN1tocurLNwTZC6ibPONXl+Vv6HJKOsbE2fxaknV/BzG4aE6AFzDoGG
YSkPvNv00XyKgW1aEImxt5nhMRrAlSYjF5mcWffllvsE31vLc0Ohjcbno3cS
o6M+Ej7K3qbHJuuH/PE+WoT7SWT1OLnRsUnqTEbgQmFP0MHpw63mdDjQnnrv
3RkTOCOdaOWTtyrQoTTa3ZfPskC2XV24Q0LMTUVq9IP2bS2AcNWAXuMXdSoc
PAHXeFfwzDIAuNPQGAHk2NjNjnQJA+LXCmYsC+TlQsMRRG2AagH+9nSYSht+
B1I3FJwUqRLYiv3xtXDnnSCtwHi5se9GJw/OxCzu/psZSEQDkendT44+WF4S
85AA2eOAYZcfNU1KG0KR4gtIjW0eWY5K+XqWb7psw9jR/FnGB3+s0586CYD1
1QtIKnSJf4i7UX2D4smffbvhEJREoLw/IQSu3Q40TnBvg8JWGPYUk/SjAB7f
ng0Plz/A65mHdW99NgE8iPrkmGI/yOuCXEhiuOozPI/zRbczaUkUnldjMElN
IAvYLvAZZyvCrAq6tQpQmXocdrrZ6t8lkHIXz7dNRXZob724zP5hycuURgH6
h4/DgYSbRmymtkapaHk7yqcdXSusJZx0OU9v0ROmY87rFjzRdYchYNmG9DUP
6zkGS/hODMcCOW2F1FetWPPoZHhHs/VNgD6TQjzK3licVFWSCnYPTspPgNXu
EojYO07IJu0U5DYQYg+c7uLnfQmVJG/UVbvgG+LCYoN/gB6Jq4YR+ESJ6ARf
EVMf76EVNuGMkoTZEwGkIk9aJUHF22bKByEwpUMoe+dGI6fCiGJeaVof2COl
UqDqXPOkwZB9eLy+YY1uhuu5osi6vewhhIfPKiNcpMhwzhnGYenYlCXXsp7Y
FAqy4QP2pg7gFy3vALa8AsrPYdPoPAMS0BQsKuyNGdYEmFqIYDRie0+mvf4Q
oqYPuCoM/kEeE8l/HiIX9NcApLDw/ttqPFCvH0jeN9WMuv3glQ/IbgDx0KD1
kIzqFRq/mZeiGNTmLDMm52SLQOWknQ85tEP4XxvG7lsIJddEpr7Wj8stiDb2
fUNr8gzBdTHDzMqEsLTpzdpUY8eIyuEbFw7JCbrMdyQcHxfnODrMJwixbRDx
MI63JRBGbVyJR0qWs794zAKAN+ccHyCXYBRjtzA/UfWgcL3E7+e/YM63VTnM
pQe2+CdqInLhQBidcU0GWTbwII+TrbphQFhlDHm45wa+Q5cvdmOytGAqVAov
cmmKjVh5cb7vfqEP4AUPI+BwE8h/XarYW6Wx8bYo2Z09NeAq8ZO9jVIHc73X
+hh2nghPCborV/uLM80n6Bmu6KFkcxXjtinHGkwAoDJGS1tFko17aTfOwiTm
v8Sf+orlHheVF4D0hVBHzjbOP6Ei3G/lrSSsxawHX7KnSEo0bFoEfP7TvAGF
aqDZwS/r+TAys4O95aYOr0Z6e96G3LiQRjn/Re1J1onknmZSyaJY4D2jZrB0
5T7+Cf4KVWXt7NgdMIL02Vu+0ghBE2+3ItujFauxSpsf30bYgsU++vE0IhPz
/Rsx4HvGMi+k+aDpDF2OWlbJCEUDHUB8RfpYCWpUQaGD1n4YF5yeH2vZACMR
dmtGlrgZcUZ88ANGY6gId3bjnrgLQ47UQ7SiuuKTnxXsrhU9pVjTTDzDSd0p
dpj+hV41RP2sAxxs8BGt8/NU9uoXGSqP/CezcdlJFL2BGaRbUBsEbr7PZqVx
J8KDcKP/+f7x9iB3mSRrQf0uBNbeyC8amxChIbNfgmLxx7eKw3EZQVXGyVKr
Ck+RrWiAbALOct+XgVrXgH90ycR0rQy7L0EFqJ72dRFrl2SPebqTyVfyzdSO
/fy3TEw+prEbjpQ+OspiQxWQF9PSYxWvO7phtF3kL5WvidC7u+zE8CCzRZ53
ckp4b1LAbJSIUfZ2jNpJe7mQEko5tBGBPj4QITCC0gaGPGYt1iYpz4WZkth1
gRBkRwNah1Ij5h+Lm/Y5Y9ldHTEtgpK8YyiFQNyoLMS7XUuvlhrjv8MQ2DHG
TZ5TeYYvBakIAIU3LHfKlnmJX5MNqelERXNQkkrPYObHdhfUcHrkrRR+JqKy
W44wY+aqVH55370nnckCBBL4WxoHo1UjKJyZkEBtB7NJCJjmMcDG5P0iI7xO
hkXg0U312tzH2ZeBLPFqIY3mtRGCyiBV6OsFfMBIIRh/nP16t4vEQY6jfrrW
lurQHCV1ciGByW2zEpus8HolxZQpacc6MpKFOlw0eSAhhpjdq6gNzBVrp3z+
roMTYiq3oj4jeFTkLidkO8KdiAd6tB3CSd4lTmTnxX3/bO3kn8ksAsfa3TUP
0RsmrcjMVGEkYMIDncNgoWriEjBeE6LWs4jnJdpy8fyrsQkoRHK0fDi9xCae
qr8XDOAIP0YOOoBZEj4HOO8DtYVNSVL3dfMLHL7rGgrjO/UO3F55aLBbxO0f
Xg+PFyYYcUGeBnQSCFBPWTF+phHPtlM+dTpChLKh/6lNNRexUjUHGafbEgd/
283Z21eDeOXAYue31LxUsqq7NFA94S9M71IfANPnfYVS+X8/qg4ieOjRQLsb
Kxo9Ed1Bw5zEaNQeSWYGOH1AavaZR2z++Mb//bTL7S4aM894J5v7UW3PkhhT
eTphiKZQwd0oUhKLmN+1s+mHqjnKtVrmskRn9Pqo9DTT/hDovNVcvC0dno6L
NsB7mjACFWS9lfZjZUNdSv9hcEV0HfzKQhI0gNG3hJuRQKKCxffG1Hb9uG42
FOQeT4/uQlI/ZzyoPqrayMd+AjH9btSavnGm9OqIEeL5N1g+GZPlG50GtS1b
XIK5ChQxYndsowmJaC3QZW6bpucArvvenraLaanXUWfCDsZqI387MvKNQHjn
FOXgMNLC+orbHWB+nfiKy2YvC4LqLQE09f8vBHSR5Yt70qweYiHCAFhgewmJ
yWFnzCmlR3XypN45Oj4G+yxdJQ4cUc4xt4qy6Dm7lJCGb7sOHIJEMiAEzZ6G
LzW9g7jwP5WLkvlOd0RM0uj3JKN6wl+NpkEMj1Ge1p/ZuIfzkv8czLf6jMDw
TQrhoFhePHjau12RTtKzPjGIJhtFrJogXFziowGbYUPDbj7hkCcZ0VHmA9JE
j2awC4YAdpeR6JT/vU1tK5X0vwFrwbQbaR0MOT0tu3mjajWHJWxov5FEmEH2
r6+eAmEX16K6HJHq0ZDFhoVPwfLiyExHC7jwHmTsFLFout7wI8nI3HseHzeR
p+I7SOpiRC05kUOjDgBcROk62s7Z3RApDi8bHUOs2LSaz8EiobgaQDtYF7d8
ToyPxg8sn0kWQMOOnwQa9FgUC8Nd2MhQPzOWkUizcSLhXwCV2XE11NcHD9vn
FKfZZOu9bwgUEM/hBkE7VNaA2jWpBbrAmj9dV5etFzvSOjpquRYf8AKaG4EL
kKhqMalDlWOeu7nZz0+MwwsuSmdNrMpEgHQNm4DYVXrxbAmCf3VmEec4okca
0zcDZ8IDk3fAL2Z/f6bBOCs+sGVyfKxAH1/woJNZ50ckcB+MixM5x7BxKEEP
UFfI6qgamBNqav9h3I88f/m+ak6ozr4o90IyNTNLNz4jRVnmgif9DpASlXBO
oo2UWn2qE9cU2nL4Tpih9nyl1ac9UXg0WTbkoO1ohPgbNF+a3lXdlngzZV2H
iFAMVXooXqNhYVLSYH7o7FKibt0j70Glf2gxF655+FLArDkLtZCncgpwEPLr
soY+5KvDcd5cJIj+YgEVwYwT4xTZSkv4gd407OLsr1isOrfVCD403Sc+Td3x
D8ikw22p/DWoaslYReine5k57K/xUmcWNIWBOuK6OvKkNlp9psqNWKFCBtDT
Rj4CeA0njGSS7lzEsuADE0yRlsxb7ffNM+424v0wfq5i9M7biIsX35hWL/0u
K2lqxmu177+Jg2uRNh7vNFbdL9PYGqbzW4o7GFIikhzkUgL6IaBS79rkDdK6
QBr4z9+CAMWi67RLtMGl11kDRM7rk1vAFNRc4NRxmo9lTQD8LuowN9DRdsWE
umgCUdtR0WUJb7LfKgrKv33sarYI33OMUYvfs2JKZa7TX74AbGUH7j9vZFiF
wgLRVM411FEjw9lqv9n6YLG/MA0zuCDgkqBzmT07XlXBZEsQlRC7YkBYDjCA
F6mcD4jqJ8jn2oV2sYxIoN5nxKuiZSrGY3v5D+YPJiBAQX3+GOYSboODkPlP
4Wjg5NgJQyRcwhwbwY1cNkZFa2OGrPJP7LpFJ2T1QTOKWYAN/yevqMaQIPZ+
ljDHVtTlbY+4ClhM8/2B1p5lTM5fFnK79NUPlTPsS6xfpbvCiKM0cVU5D+0R
/Xw2ntVgMcjaYLi5iYh303HvuumToNdaZINquCSREJjBWN4bUcNe9NpNmfgt
Ah3QI3vMFG+a1xUpDX1YE+DlEM4e/b1NM2Xh1gnwS4RwWjkLSNzfYAC+PH45
rU/BWmXeeNC5lLeV5wiHNCk27NHosvRhoDm0pAaqLSBNn2YMZVgCjTS7A+Q2
zZYV8MBf0lOujxp26gEIMea8+MyQMBnk8Cm57W79GE4oGEoc3ni9F86V+SdD
OKJq17RHv1vZmMay7BLXi0aA+kc6uC4hNhDKyMcP9WfXbq5UVKCtJzfITHOX
MWxyc7b/Fnd/tf+GRSIKDa01oUa7nvVlIkNwpurrQr1NbJDTlAhvyeFt37md
aOceSb6FCLL22HHP4SHp4nbU6vmNHdmRC9BVLQEjeTaKDHjvnWCgHnXEbqPI
zhLir3Pw4B513j1XGA/OnyHvZfWkX797kq3ahaNifO5uhmmZZOB40c9BRRio
Po9Y1ZzG6NLVbJ9eoyJKIwqYpZN0lbv4GjQL3Fu1fD1/NB2F5huzu2FbYke5
OWmQxd6huyEuCTEqGoVOcnd1cqYBfDk3wicIPLlDXZU+Jh+pfM5Lr8VLVlJ+
MqOcppWiLpFfHZ2NTyxo1PIae3b5VYSiOc1Sz64LrwC0HFNyY2Nvgi6MHi/0
TJQ/ozCJ2AcF5ZO/VHZTP0dR+37IbqsTf3s5/Skhs55bZPeY7MJwkoAxQuZ6
v3ZeJpE+d/IMUKk9e2JMHEp87Dcm7TYt4m1lLp+KtbftF2YrXiSnaKhvqitO
5bU5afrdfMxDxmsWcTC+0v8hl38GwByiemJlHQxWU1Vcuk7pvFaQUOIeFMJd
joC8Sax0xWrh/IAxRw6rDkbZNUARyuHSQxG++I86xv9QhchaxCzp3kP3s2qD
iLDx+juLVP4y3GtN3d0eds2dKPP1Yq9I4BC0M1ztvByHUWL/jC70RGBDqoOE
NJEhiCalQzTGfub9xuG06r7/IYuFllKtsMoCbItzOoVSzofSPfQYItxlG7XE
EHrWUOQ4r+MEsGogGK229sG7AETup9p/ZPgPE2uhaER2TrwKaZtZdR7lXyAN
QCFN6hxBalx1ftUd9D/ygl5YYzmZMjBSFz0uZZfndDlY5MgKJap/x2uQTda9
pRrexMQNup0zrNi3TegA/tnvloCDj0hFhov0aC7ycd5kkU+hB7lmjhjGjbHU
lAtINGnOD5yKG7CY+O42bmFXqxE2uTlIyZMnnBVkqoP9k3W5SqWjgSBt1tBc
SJGveu7rVftVzkn0klhHZ8YXhePO1u4gwfxxucerqZjkYb/zgJGCL5Lwxbb8
FcJ/M22ZOLjGlKcTMdpBN8n/JgX92hnwwUn/X6m0XK8Not0s9kj9e8aTERLn
waNkvQwefRtFjhKsI5nRFOj8iSoe8oB27wOxx8dCJ8pOP3OibryoOvOfPcDU
0jTbyJyijB4o3KwlSHQED1RIeE0b5WenMvbQMjHniGLyAV6MOqJP0umCfpbh
l9bI05C7ivVZYDMthpmhwWBw9i4daWvgpohlnXD6ijmYR0n0BwOkc6WBw3cS
J1AoWIAyklyXcgLpNh4tHF3cDmBMD2OeCWBOLB8195LPUIxyaK8VEkyK9xrF
KiafKhRu9jlNrfH8ABy+PY7muDF8Eh5JOMZyXxOxxv5lfn5cUyUbXy4Y2QoC
M7CUb9BX2BygxL47p7Z58H+oLjnE5f7+HlQbjzZ3vCeWhdBYlwPveR7qN8ky
r1uaucUfZVoRtAZlkd3fIB71zsbqR0SOYqnnPRXqA029v27eN3GGEnuCuJvA
c+QbdwN3wllXp8T8wUD8wWSyUbzvQIP3CCaLfwpoQHh5fWnAwBeR1oCbQlij
7Y3Pfh7FP5+jPakxIJweFd85WFc8v11ScNJKdTTptULM7tKNx4uQaDC0Porf
d1sfnKTfN4MR6haAgBhRzk0QAS7nrya/KOCblscEY2Tv9oTwT8GOGfwsS0ic
7Z+0Yr1bfxzy06O+o4LIBDkibfYthE0HaJOw1ETEpTAs2XbgXGA+RVm1OY7T
CGgJ0/4Qo57wikWhBE7v+1uSfm00Ru84WD2iURsJnxL7wQQnhu79IOPSkMwE
hfS0ymzT6oTRQzfgFuthOXxjZ8n1FshSK0D4f+1ql/X2epnluRKzBH/HCwfN
InatX/Kf/KMeQ949nCkAO1as2NTmxTQ6XZWbInEoIBWbcpuEwvrrDEDMLMol
v6NAjSWgnies4HwTDhXdPTRrcnKOfNiHFQ6UnVAmMyvc32WT8j3NT1fPNXyL
Rm7aObA2q++YGurwV1MbhpXDKoQ9K/qlq70cRRLznoKAzKGfQiI0DDtiCC7Q
SJH5/03jxhFXUbjwJYbF/SSnG6Ja83fXay/7eGZTkFbKYOMiJnaXTY/Z/0Ol
96YI4CrsXIer7ArRknJjJWGsHJZCjRVHssb4LwCzpzIW8ZS6wlSmgxDl//ad
jVLCxJg0SBp1A7nBBQPG9tAhMevcQsPDSHwEqeMbZ+MIGA0gKdDOQG92MGgS
+ileKSEQtvzX3w9VhaTW4XsP+d0Wuq4m/lh00xwigUlr+wdVSHnbwJMZ2/ip
K8jX5peVW1w6TW1PjzHjNmPCJx6BbbaGabwfsMdzl8EnV2E6xUItGrHdE6du
B35MBUPdYuiW6d9N+ZUVqr9S40sebwODweUnJW5EnKuNNx68qhtKQVQ4P6eX
UzNF0s+FrJvi7iIZmaoxRf4MLW/uasQrGa9NGWcFzRRSnYZDRARr3iq52fEm
WuCpP322DdD5VY33fct6mYiyfU0QcRQTacjnSC9CN4ZusOIXtpqnptRT6isj
gSxuQ9X7hUATaKG4KttdvnY3vZtv90kot1FhsWTKibA0uIvJUxnHe9zFTyZk
xybkntb3TgTWB23JR/ecTQPh4bocBuoa6au8RTxAgagIf0r23IYj5uGTDbIx
CYhfCj9hlPU39vVKbvYl2zHPXeeZKlC0tnOF7taw2g7wQHORJy6iIqPKtWJd
gBZZ2o5kPyztYUKm837epltX8rO7bOjsv4VUPSzrpjAiat2vZ7AsS7LrAfcN
vW9wwQGn+IpPhRxXtsWjs9nIYXP0ZwcBJUSLzO8ZPnvxbXDc8S/SR13ruCko
5hHHfL80L3GOik/hzkFjA/0Ypugpm6Ll2Q3bEB7Vlrdb9d1OvdW+bwsOwyI1
dVt0e3QNkpQzoExdwUO7wAgcHFmJKGxGhGhfb5NPiA5uDRtgfrQsJcZjsZH0
KzpOeqpUlafRmzCIdxfmBPkkWw6h8M21zSJILDyB9hB2pSV2n3GfJRR0DZwn
Sdq+vq7FzjHB4fCRgnqNR9WPTneoPuk2fpEAXJVix30dgYt3wrfa9B9ysJiN
RTIZbaXrcUP8T0HIKFZYIqskfHrBIwrOdes2OxpCUA4adu4K2BkOF8YrivB6
98zXZDsl6UD3xOWidsF858RuMEH8MQ8zwJzbsc9jaPIfKIDdjyHVPmC95fek
h9CGb+Is7ajMJ0CoruUNCXnTMRcTJH0M8zGuoTyt5Gp85eCu/cOUZKxEPPMx
8kcZJbFx0zQec4sSErquqNQZgFyLgAuV53DVrvpKKoYoZ9vB1hLG7PfwngFi
X7Dnt3q1ad6LkZL9UxCMbSOaXvu76cV01KzXmp6fqpgeGB3mtuEIV2JGnCs/
r1DCK2MJpx0rM0d2DvGwlH79IVHnl+EBBizc0JN7iCajDE58BbDwWC2a6jBp
ObbqZmKxN+wuYxjOHJgDBwzCsg2NQxj5G5ewzKN5JXozwjnt+BGUCGs/O2Fp
R4lnbQVyu1rusZCij9qEjXawMH/blEF552CTlqa8j239XWtr4cI3BMKegRkR
jLHfQVvoJrRCjNCWTEjRmhKLJUiUem1u63xqwkmWrd5FYYmEGMthPDfJgJJ5
jdDYjzeAszZMhfqCPEr9IN9e2hwCNif7DFQ3N69yDIaGL1MKUkBKl/Sgibdn
uxi/7VX7eRqOYbF3eF3CNrlrtQyzHy9slAyAZ7IROO9EwEkZoaNyyndEY6vO
4QVMlFAb3zm94GQjRWj3QYzAQiKCWpVdg4gr+x61rG/g1VFhK0jn0Tq1XNIm
N3cJ936Kyi/1aIyLabP8O9a7PSenMF9HCyYDnFqsl9i/7voqfvpevOeIVGci
MHUj+pVxY5h41APBf+a804yUNQ7HiQXsLxwbuRPfZxezm/AP7B9PpvjK69lV
2mg2pcuNzV7t2cCJePhd7jfbF8TkMXqCrRa4U7bh9ZX7YVVa4nzC2/rmQW4q
al8jjSLxbiQrM8Ht0KroPz7zHhBq+QUh0IgWzSHwt8UBw6vZiA86PpFIgUDW
ZzoP90mXzJK70MIIbc+u6tmYEEKU7ONJLmaSmCqXy8DodLVVrKdWCH9Lfi6q
NAxGvwhyWDCajOqdakdOxLOC1tE5oxDrEHB4/8nBLRVKX6wW1Em2Gx4yKj9v
PPBWt7Dh48FKVM7Q2h72cVuSeyC/WfY+ZLK0l8GLaoN9VtHwffVATN2lWYYq
+nWrzZIvAxtbb8e9xdmPjRbxSrvBVI/pV+P5asd3LqD5UXb5kcw9O7PP+ylZ
8Jh+8Yq7ikGjScuz9MG3d/0eSPOC3wEqvEIfwHDXfNiJxg4rYjW30zY6d4fw
uGIyznzJvTPR+jXanUorn71zD6zGwCr7fsC8pWHY5EREIbBRt7EbHsKFnhgO
ybI9joNrEqW43pBiALbZuH7/7WyDgFQx+b0Ae5XTeoM3JFd/l5ZeFwf4Y2pL
YaWNXdqIRxW9NUa3hC8DhMHicg6gzn77k+19GQmRynwZBFZE7sW2a8Q+eglH
BX9fd8Ga6kngEvN43EvKFiJSxNa+FFmcs3+vtQEn5fGAOBy0ohVIeabvuTDa
qmaA8yZzuKd7XTN1kON66o3NCvNFMkeu94eKQ4YSymVd5mRujCXUyw5RNU9H
S0zaOWe3sVffyst50zgI6aJlpxI7U8lOw1Yhz/ewKHhmQCCKibvysZUmeJnA
lris7df/RKyG4QJ7Ir3vRob9QTOeTPbb+1Ih8zGJ5gD1kMdgMlDKWwfQFgT4
tKBXdgmehtrS7hztY5KzhwvcrZvPFAmXnHCR4hVgU7RBUJq/QykkysKYIyha
N3N4CajxEdSZqcpIlj2BAqNDgplYRK49xxLry7ghMIeoWC5vlmqZM4mSGcFm
Q8qLKApAeBKGMt7XB5jXrlHJiPuSLlZTieGi6LJEAkLVQw07tS5E2zj7CYA6
CylUSgLlafKOYGiDa6WoZtAaon9oOReUAPcE+6U4HgjLvZskN2oZjA/i9oLP
HINhoy4dMYWXK7wR2ML9boEiblW6j7Qps/PZJOvyvoZ6f41zlKCQz24UNjbQ
o0wJ+oXlv4dcqf95ljAr+ssilF4gBUjO7AmLOfb8N8xxXHVX0n5cNtd5mhWb
xuWYK+7dQkzwYuFbILF85pkpFIdMiTHV772H7FynwIqD6ESqIh+hyEDELlYC
q/+YgfBa+vfScIzNcHPupcX/unC/91ckQYtad9GS0JRluiOKpllCGQMu3kBh
7xOPMKtL1GQsijZGH/XoPn02P4ksotw7WZIfMSU9jGbsbYjH1xhZa8t6huag
/kjTGV2tEM6P4mhMSVaKGKd8n5+GgJN66hLS/z200B5psyoxJKev/h9cncxB
76nFYH58MRYpzUJeHk68wwr30QfTvMbzszVsn0UVsMe7dF6IgRhfZW3Zt3CV
JkB0x2ekUM3mcicmjVua3+Kv+dezuSv5L4+te9VB46UgrqdrIqAwcH6kwsh+
n32O17ED8oL5WtYui1rJvt1ywoNqxBZUku2RFaqOHZWEL6PUaGxB3Ug7ZDb3
Hat3ftA1kPfU9FrGPdS9axIQ3FmLZIZEcFRFstgsFLMwy+gN0T0cSNrVWNbX
TLJtBFDp/Ri96WqFByni8gSD9tojln5SolmeOTg3leKHqlwoDkU73caWJDQM
B0oO2D0OCALFbV1SdaLffgL4/UmBOodUs/dpe1RCFpWNTKzi7PIZx6Acao5L
Da+aYcPH7HzCNpZD7cW6XnWwFgRnuO/ajFGaOHyXNjkix1hHlSZwckLESfn+
QOaR9iIT9EhoxxLyGp6eTiVqOus/NqoAcR0SrascuMnQ1Y8Icr+pM2CUuAdP
i1seRMazNWYTBTNH4n9i/IraYP3WlvIR8IwABZ0GYpagXLcWlVrDBFfjQes0
t8r1JswgedKaqoz0Bi/p8YVsCGPTsl1Y8Ja0pQcbRUvGPEvA/69k6deTX3SK
EFRqprZKyifa5u4IWn8r5KmvsTm5uwbud6cEn19rYteYXaZLeJPOIesUKrAF
WLGIfs0f8yfT+tw0ZjIVO1EZQaDOLxqpqetVe3HBp6jeJqJXS4yZHmSszMBO
rL9tBMy61+K7vAadTDbLooGX/d9eGq1vaXk8cjc+S5MN/NiHRHd7OXmRpxXU
OOrfn6tNFV2zzxIWkLo832K0ZSvYEyx5A5sDfR2h9kO6A/liWhAVhxxt8hGk
zS44OLiQ1K5Cr5tXE31Dlr+w3/e94AHZXf/IkcDoMCd1x7vwFovqg3LBEu6n
x7sfpG8Z9EoG0mGmQImACu40noyrDKd46PwoYyr/7T3VhNAMGqFOUietjw0q
v/wIZMVU3AMoKHrGMf/UH0bzpW6hcKeGiD9/IpexddgUj6iJrxXmvxrSDLZq
JqI7m4aZV6YIS8MWd33OMHml2LZirrYEq8IgSHa8C8ICKJnCvadZ/NCgEp+N
o6zqmxRUtJ1LVHeTn9q7z3BfnvIs8x61ELLYvNXbeWt7gj+JeBbYDmGTAas6
3DDACtCnwhjnZ5E43zbpUpRV7Hv+2l+WHH4IxjrRTF8s1/MGgbc8vuJzeYSv
GSPfuKTl2uMhuoD641BACccdiEdH5L4UECWlw0gjddQg0A5NmZJ4yGhE/hpt
qGCyyyvL2XIOGBz4MI4ZEtpquAtxPm+T7IA19E6aJhy4l3DBqPaZ+FEdnTVX
JEFeHokmnJIiId3oRV5eTxrQQlZlp5m2bzhEajs2qGyIlZFMGQyhP3kfaTKJ
TPwA3E4XTa53QPFe+MDVaT6yIaipduqVw25uwsUCrraPaCrA9z+4qGrsKkc4
lIlY7VXeoy9k3wBXcMeXchGZmMJIvLH2mClxaGVWFToy0IeVrgMSL9T5lvjx
w4YeLW+g5WQ2nlAcS4T+j5CZ07R2AO7Bg6y/Dbv77fzROr25LKpNFpL+LJm2
hquzxozKoY0KOnpmVuShbBovFfVEiFCvOR5fPbkpf2+ZhXyTBaHENjJiTjri
CZ3U9wj86trSUWCY+mMBvW+HLclOrC+D+4SajSUPqkVsJzE/RQTumdEP9KK/
fpnQmJCEXwhvAVGJRHXm+RqIeD6OGvPfLlNexHUj16fD4qulHRX7IOsHlaVx
lsTtb3a2BqTR0VISZEk9l3gfmXnjKuReYNXHIo5rcwv4R/OoOrN0u32AaWE9
7ITzJ/CSJnRZDqDcpen33V3JesCloGUyER+1qOcem+RQbdgrAFKhVZAoseQ4
UWHEahVibtfX1N2L65hQa/fWRjYNQohXjTleUzqmPPu7YZ5pj2WhWun2BeSO
WqDSt0z5bS634B1K6Ge2Chlpv6YQEHr1fpW1fqF34rTWnnVnatB6n681pmET
hk97pMRnAtG1sRmefEPv65dfUaQfOwTm0D+w36Rt0JTyCXblRozKP9kMgFeX
Qxkt9xM5WtqeE5RuTmUY8isVjtC+6S3tjUqCi25Wh7cgTuj1gFfwwTTJ6+fG
cziFLHFaByB2v+QC7wYuaseHK5mj96LwRrjV4hYG5hLh9e8EryiIMhvv7hfP
ANRp+q6es0UY+CfCuZl454O02fnJ8ZEECwIrkzM+XD9tJYc87/IoTfuksmfm
OEc/cNdWoBXk02JdZWbgQViF0jzxI4pbO3OPXCC4fgEYSVZgyW7Of7Fuf849
atqmd8ynZlf158ez9B82LCo/CJeCAH5BgGvwkDK35JunzUk2j5AdPcG4JvC+
KZSvAgOD9MRp4OlbmHqfB81LjWjdaH6waRqah/S7QBwwAwQY+3Cy3XzerOES
9LtBFuQMBqSkGIEUgBaZ2b1DFG7r2oHfjMfqBIGH8GTwpnyNl142mi1nmU5k
4S75YcTC+NGfFRBk78YS0Ci84mllRdWLTQziNuXzZp5z1DuqLvvY4yOl381l
PZhclDgScyftFg5ebqvMen2VeobU/tQiwDucOxMd/H36SsaU0pc9m1t6l8d5
1194uW0oC6cJk92pBFbx2Aj3yEpyIzTma7wQ96KyFcek4wqxv4yUSygdJcrj
ePkFNWOdnksI1ImW2/VSQcmDhUO5ln4CvWFIHwdsLXQYAnnBpd+/Gg4OQ3Tq
bYplXI6eoNjro9A5q+4CUjeR4yGqmqtlsVIWe0vuqnMOSBjvjHIX7Rm6/XIe
X53hPUCGwzLwkQr/dM/IeCBN12NXGuZ069tDWIj1RJuBGN26xHyuLYGELXDX
tCZSbNTn69dpPPC5dwmyl4SLxfl8XGpJuG/da1WNIVT/uFif7bkrnEANOzFt
Z11yVzQ7dZ2e4jr9mwuZTYnEkwJpww514ztQszZSv9lt0AU2unUsymUbsBvX
z6Yi3qbFhyUkV497xLYo3Q2STu7ZRG7UwWAmm2Rqeo5gWY0JzxKeKuiP6agb
p5EhF4fL4TwtYx0+q1o6G9HYs+V2tY7phX4lsFeDTLS9zSXUEjTif4BWp/0Q
ADvvh/D55JVl+MAz7lCnuzv88L6vbKLuXPTZAT757Gh0CtT8WBwmrzDSGArA
SSRXu0yXDUIpjgw+W5mc2FGO794BVz4DDZA3kwxeV8f1QuNjIGXdBKQJOEah
1qs7o8x17qnaLUb7xMP9LJN8oy5poH9x+bEPd7ytW2uJoaqb36p1+af5+q//
CGw8DFkcZntIadLwYoi4VOFrROXQFIXUk6fbn+fALX67Su37+MRki1Ns83RD
+UUMzkrCifu15PIVKML5kcDVj1DC7sWr5tn4t9EHV7ta2bW+OIw730zBYjwv
WFZZtCPikjf1i3QVQAJ6jelrrSOLiBJzZgNKpV4efMFVed+QsgbDAJShEMLV
THCmbHAbKjVBUIIX1WNJF2vNJ8kWyy4xogImN60PQCoplnWs6jNCYl/aGi19
9hx5zKTvlKqEXaN4iqVMljYQQbsg+2SnNJ9hw/A5byUWFbERbJIHsBy756gw
4/KtLMPxlRCgugpbO0LQA0Nuxp/WAYf//B+uy8ttCCUnB0n86OxH8qLthrI+
RZtW0x85aQFNWQrNp0I0T733fDun1VhNHADjUtITCK+ax0/A/D52q73Ian7P
7r1kRwxHT7VBCEFX+Fw3bA0u3nvuqc3TImssWeGgoeVBMvvntZd1WJnMGQIC
F61PNtmMW3lt04PaMC5ETipuI5K3lrTjeb3S/eughCHYKaMEpyC1eC+rF74t
EE2KrNLVp1RZqmD/vq6d/kA5Ev+roYRXKkT7MMUXIKqJdX/YkJVTUSRl/CQT
52oUuyKCMTNsAvKqEq4GNVWJ2B/CUg4Wzn9U3H/7N3xgXktsCGHOiUyyjfkq
sKveJQV1EFiZCDbpvXtLUDFxiL/WYp/HrP/FhOQADL05HLza3DVS3AJZyWiu
AsYPqlbLd+/iSTTWbn1LoIVaOf2+3IG+AAozf41kvMlop7BI0OPJlF8iukXn
Aghx/qSCKv/VPLcKq41wOldlqAJAvgtKH+PZ2K5hmyr10OdzPvficvtrbi6x
7w5YznaxIv300RFC7H9O9MWWGfIcLNlFk2dWg7s/M48ZE+dvDea9Yy5UNiL/
TYfx5TI6x1RwXadDvplhxUDI5OOJKwUCS5qfW78aywmO9JUZH9seW7BP3Sv+
IaUF5KI3lODQUIloFniAbVUPhqyUsxq22bpNVnuxWe2vQfM114OSgDXLeyEq
HMZq2N2Pl8wBy0AolBSeODCcLyPuU4GFC0qOEhLAjf5XB9yWO3QMZaTwCsnh
visuipewFHkYGP5nuDFgV1FGL5jDzMhjZmGdDRXK5zbCvCD4WRZ4qC0AqNrh
VIqKXAZs6zT9k53TE4RAWLulRoBdux/jMu9TMjtlSqXlj291YrOYt/pUbd43
7ZkhOpkOu1bPjI0nQBI2hr1JbjpOglb1BYXYUMyeHE+lWcR+GzIowK3eI1D7
LULB+bV4urGwT17m8vA7UpnaQ4jHesR9xkubn1X4wgfbhbu2oUJcvlIZrzkf
JmDgf3ujAQhg2OblR+g3uk5QYffnnilE/dGWY5iF9IqC1XUMV9Eu+C0SDTzm
raw4VSD9Vp4ZxFZFWJjPSxkBVAuI32tblpHSLNqb+ZVXnJN2NyvF7nL+yLmU
WCD4N0kJqylqLCgIqVatTgGRWYXJYUpnlcndw06zH6auMaa8mFFfvAGTlNjH
l9+5DqUEwZJSMCPqeyaPwEt/UJiNdxxmFaJbHEigN+iNgmeSjrfNsQa6OACS
XuhYpKRSWhpMo1mpEZOhwJDfJcInHMf/LC69fH3bX5masrEjFVl/M9wYyvZa
VsE6MtJSnzoF8HsLYjEpfNZFExy1a2wWneRdayRPTRWEhPLq3sbxKqF2doPy
rZxadis00pCPPan6ghJwRax4Bha6oCXbSGKTC1aLYfDQKCggcC0XKz3JIZbE
ZPIbaEtMTPRybhoahUPgrM/wJ6f95H1uMPnhj8bQRUJNQ4rcrdsHbBGiPSdC
qZqggCL0xiag6HSn9hDqY1/9PbUt8nhfaV/V4BNNLn+eHqe/6tPFVWDy5zsw
lKdZrMjxxz0e7Rr9SsXko6PhoaHrrxFlTw2+9cZ/ATgyvP9JqpF+BMCpcLUg
XNMuvaXgS/fPDODS1XhKObwKPnn+rIUXvMjlLeNRvzCVb6iMW2aMM3SfR8mt
MDKvd6aC5Gkt7F4hlpBbwzDZ/bhnyPgPV6IybL6hw++d5mPit/M678roKRW3
m2lFevmP/6FMWPeQQyA0rGDOprQFsjzvzAy83U1HBg95T7P49gY0yUqytruY
LXFeYfKfSXCHhU4Mq9cj9US3vSRVGyalJE95SlD9u3e69O09RfnhP/82lMIp
x7wUtG+ERpa7hEIWcxwqLV7+lGfjWIY2Lcuj38PBFU45hmh5P4BVagW923LP
IQpLhQEnmur0ymf9JNS8WUacHr/09qBhNZi6e/WNr/8BE61jlLghvEhMM41m
4kjKjXBANS8I476vCsddAKiRLiXgN5Yj2W10mMIW8FvOeHZg82uur5nt8F5H
ZCuAfCKppuNQaGKGs4oYJd6dVFipgTKe7r1iOs7jMDorh4yf5xgNutKL/2kz
Cq3hNS6qgqgTrv9PzvQ8MCITFxRlJodP8W24rtZtDwMq6Euqo6HqFPvbfXro
VxiTX8bK8QfPjBE3m2CtqM1EDYldTrOFz6mQ539CY5bpuqOkhNzp0JTuphRe
lDQsuyk0+NHall0izipUkckgMXy0c6GoSUUg1WUDkAIcb2kgKhSzxQ5LOWsR
nm4lSr419HSIqNi4rnWQF5LSo5wZn88kYd15IV85iNEqN1/xFN+cqH71KJ80
7LNfWktKQHSXDK+h9Rp0fPdtfDUyy/DsnCqyc0ks0rx3KEGxKGvevtp2kwlV
jHRM1xc7rvHtucE8z6XUf59icz/pYUB2swI1njyqdoRYm3LbrqvlTtXDD0wk
NU8dxosOyGShWVLKhDoVygs3jrU1PWOMMO9OjqfKHfE4sPBMlUkNWHgNPgpi
AbkUFIgQsn8xOjDdI77WKjkbibO8DY9IskT/fepdpkzEK3GwoCB3oyMDRMyS
Ec6FL3u5h/3RQpoWfcAGF1hbf1O6i42/FyC87hL3qGBGACjFmvfGr/qS1qVe
DTARr8cnvxjGZlKJ5HAegEc452S+BeiD+H9SKoo37Ylb8CxBFjB3EcI6KAqg
ulhF6YQC+w4+zK++D0IIy5I/ZWYriBioukpkumMs8hz7rtsloWE5XqjW6sao
W9P/zVsx3IWLId4hqN0fAYumBzhtqXLx4/EEmY+N3F4E0cmtQ0eaZpoSIHi7
K71y5Yfjdc5swTjTb+6Q4UUd0Mq5mMORsAI7sH6OgyvGvBG4qiw0T0w8iGAt
6Xix/Xp51M+EFsDhhwaP+xJL4g0mPDh/ct6vq5EnipQ3pxLwTBGQI69oxHKS
Nu9710mnKlzzB0lGfEF39Ru3zZkXAfrDBOb+4ErVp+h/O+mmTGWk+CGk6YUz
SbdW9OotVbZwqOn6tEMpkP9UtxTmIW4WJXcTHrgiL+gwXE81nZ9RTdv65Ye3
/xDthjLMrBAuSqbdEMMdV3FqJP0bk/W4uMn//T9eG3Ig5jhkuAx3lvNZ3Oc3
dz9Xp6+HFsjGKfHY1/VdJ/noJ2o9U4wZvatyu5W44bH2pI4oBPitFc2CRzuk
i6pJtpBjoufXlc7omY4plRIwwa3mqtY0twEnkzIJiwdlgzLlyAYT1xirKVYy
qnF+3Q0tDFFm8vCGcnOEw9f/glnVXrTWIVWvb/Ida3xnwYDBpj6xDt2NF753
Z7E12ZPjlnw751Kis65WfeVys2GJJfE+FevZYcHdOV9pjtF5ltacfEtCWMga
cHsFY5YkxtpwHpOqXzquUQyLP8Ae3LaEmbbaMyKYWQbGNGvAZZOx/v+MzZ8C
piEwx28Z7K9/xVFLQoHkqsuPAazwBJkQ5KofMWzxSI83GwI30gh9ycrmA6SU
KQdEVbgJIAqbbfpH7lREFIA+ZiU5wNo7fZvd/N3OG4A61TCcnqDXT0NIMbzd
qI5Ak9JZbb93dLqVG2MYS/d5t/Vtw5ZjR+2hF9f9VsjOzi0Gbq7KQq6gV4Dr
SSfIU7G+omWf/BXzVEAfsSZGtqEGnL5GAYkP7D17TJet5Q+5kS5vrjhuGhUA
sy7F9X3YbQXIfw6egYfMkaqXk1wxZ/UUOpnBDBy5qGuPbcgymig8eAXmJrWb
P7oG9FkOnL86cQWRYyzJKmSQZ1lVU6GlClZYsmMxOHIwCufvTzHKXGVygwre
sU/oOcRp471E4pjK1P6xlO+F1WvVGSA4dLcVJHzNg4V1mAIm0NehJ88R7qq7
6NXibJ5s/cvA3bwJT/iadggPGuNhwdHg+RTVWbYe2DP3gHCx4i5sKL/VA7FI
Q2IU+5VGcAcY0Q7MHl9KuPKjK4U0jgmifscV/9MhWhVeUae3hugWm2IoXsXU
zo4xzUQpr/njr/ab72AFhV/ahdRxVAU5uF0nPQtPUcYPOatJ5h83wEGsxeKo
mL9Ipf8j3THPI8WONXF49qiops0mGGQ7b7r2L7plq7YYVmHj6Udg5Qr8VDYC
OqWIsoJAg5khi5eM0dyo5OqQjl6ne7WKmWqhTCpYi04Cw3qQf5fgTi+FGMho
jdDfOGWkc4KHKWp6fBpXbclf8S/IaZASPqmN8Q4eEyKLZ1ZPx7okbFd6rHT2
fLuJl14QDo3T/4Xx0iJ9eiiFEx05DxTgcKW+y3PvfZD0o1iQKrsYOMzdSyJX
qq1KMzNv5JuRb0D86s3Emw7pYzwTZD9WOa5eLDGovHJKfB+ikfbAmFL42enp
aXkzZcVcTkWV2p7dh+84IxMqymQJmUz7G9wym5FLZAhW5UhHC2Z721LnXGVW
qPGBAq39rrrf9/Lsj52KR899F4m5air17Pes0iJhguDV2QfwRp3Xe4faSjNn
FKzfR1CSld7OS/zF/yx3Al2CFD2YrUxibabktXjL5ap6V37d5Pl1JqKjg+Fq
4KRZc8ZA5T8r1abYKO+w/rsU6GQf/acXgD56WfcFKn8iTsQAfiRME3bsDbVG
hzBQ5yBPHy+P4BzZ9rj8Eptu9lobmtfYpiWycPC1XtaFipWeUdmDJ95EnNKv
Zo+rEqx+1IGVl8LMqtpk1m+3KPThS6ibi25BG2Cv65YDxWVz4bkqJasCChji
nPkHoLbyGHiTMO3L68tsAB8m+LLDTQdE8zFIrmUWBWWywXiJpK/J97nMPurW
mTlBn20jHlp/nTbNi3EZWaqbPqSu/MTp7UDyrNmy/yGeW2hHL3v85r+5Z31Z
aT5jMPp+jAgJbBYhRAwDowG1MlADzDp6ml8J0J9KNzHcMzAAcGa4pWH3Hb1F
XmsqwQE7TQjSfT6kqePKGboDwyhT8biNDCxCkYtDUzrkK1kR5b8HypaP94mf
EBEu7QiMMjgJSSD7nKHbcEk9bj/0+9mqu8i3i30fRKKPHVGaej35sRD+oqx0
32mOTQ+ay9qvOiaJ0wtKRDPQWfaod+RbuNxd6iB4WHtqGUeVb4ZWBAd8i0g0
zRlJYAUciTM9WTs5hv2Y+qioU/daABpeBAIFpcS8ZJr4FimEKQSfzjg7fZsr
YDJ4g5edmf2bHiIt6LS53ytQDUpGisT6oS9gtfyRVPcZHABSR1Ihxbc20ymz
Dy91/9U8lcp8Kdb6rZhY56nbOr3/RXkDkAeM4Bj2k2coVYWaCyr1IBo9ffQH
UCPe5cTd8bk1+M9CaRSirayPD58opXEm4NtB9BqY6y/YUX2p2f8Ic+oQztXX
L8U3f7nHIwHUn37R0S5KkqmqwNu+WLKcuKbTF/yb9sqmgY8MUdPMJ29vlUB/
jS0leYQU9sOgaECRnMQ7xr8ZHbpX8LvaswvB7QnvKX1GzSCZWV5NhFCYead8
XIsPdK7YfBIFqlZ3E/WBvWyGcAQvJa2k0g2n5VDTMamST63MvPmdkcCfANo4
cYoK0jItUP92CrSCO82uVUCBzNwS1b/i/NA14ii9pFtUiD16vRWL2p57dtqo
dbNAUca1elpHppM1AogsMn482oll0XFDpPLTxDliT9Pb2QxziHPZOwwaE98o
tMcWKbgZE3m6U8stbsQlHVzagNBZd/PEHB3A3lc3sQkaFJJn6suh4/08Ihco
kkuya29Yyc9qDNQkshv9Abap1Zi4YhKh4h2Q4dCGdm2WS9s+B43Uw6SuPW0k
4QtmtDbg3VaqBRbvhmtsoA9N+M4jFrKRczwYPXp0wgKLjNhGSg54lHXRe0EA
mG0K+JJcDvvOVutfceoxwBFKiOIfLdbkYRFdElRzQsy/vYR3T3wJqoKF1KNa
nUZjPgVRPnkKIkuyjOlztv7f9q8YbPT53uwkvwxsfAtSosVjmIpDtweWoUEG
0KlE+q2gJUoEDpPyms/TCM1D3eZJdBpoaLuFYGIM92fod5ck5sVQZ57W2yxZ
KVH9rKl81wB5boXi3JZszU0qGNbhXwLid1yhSAOV5E4cyVEQISJWO0dOFqNo
uy/MxS2TtRzQXkpz6dBOF4MK/b9Rof1qpXzq3F0PaQZxU+sJxjOucjfWkCao
yd4xb+JIReV0dzemVpOFBC4v5YrugOnfCmtegdzuGbWWxvCdWSTr+jZhZa88
ebPIUgW5TENOSDUqwVhDycFdu3g+SehSZzmO+8MIw2yib6CI1Y247gpvlhNE
PwnAz2289jgeGZVeKsM5co7D9AG9cmQXq8Xi3cOxEDKprqCjWPlh28RDl/yT
maqENcP13nlRUj0qszJbshC3OOxiW8Y/Kg8E1ej0qaedGndO0MB0MbYgzFhl
V5mclB1Rk2qtnw3We+0fiiJCBWdJC8/mGJgX7jYv/UswVvuouKyMpPLnoQXn
Yk9H5cgYrhZo3OZwgJAEFQ68pCZUPemZ7sqOk8M3NY9DM/twjsK+QsKDZgNQ
jX2YLBKu+AfygPE03It0C9DUDTeAPOp/embpjMU8hnO0u8kU0u8gw6hq7QFy
eqS0Jqfs26lzr7bYv/otRQwiLtH8gynFx4eGb52W19cY1NuZwhZaxFwCyc3d
1a4WaRZ1J24XfsyPSPlhEPJbvM8LrBBSoahxfOLXxGsxenY609nFLKdVSNb5
GUPtqcum0bdFLr+OcxdfewLNYQe/7uXPTPOKl9Em9Q/MM9rVcUT1JAJDS0Hb
KHZC/uaNrWxLg2qkpG52pBEUyHMbAgSwoFsd1tBuG9C1YMXmhOihuaaCUO42
285WjLm3Vva7Wu9IptanQaQtOx4yp1q02KAzVPmKigRh5+3YyhZBqek0TlCB
rKj+Q6cnDPcbJ2HFSdHGiciRX2wiUYcxK5mapLgzJYMb0oFij+cEk+44Zhrg
d3m3E+TfmdUDJor9hrfudMQ9n0GiXA+9Y5lJN21CloVt7IyHiBTbzGV29QEI
YFjEoiemjGgcQnVJysvB7qJfNgwkME4QXxCpkIeHM4XWHEN4OJ0CEaELk8XV
2Vt8+sUG3/r8Q3y151hgokf4hwnRmxjcO9F0wLGcTEZ96qVjenD6qKdenqHf
m96qpPnXdAwsNFNCkJd5udgLK0HuiUZ7SLwh1Ubboc9zMl/2pHjv1Uci+mxH
RYEOS7seUkki/kEkdfQhNBzAl9V0yaEiD8lVNgjGlOrbHV8xHPlfApgrXvC1
KkAUZT17FRdZ4N1joUM75HFbqDAsIXEAsl0Zx5pRUMdtxdF607HkmbmNVMuJ
FCMOqsvMA4R+G2Z5yMsy2X1oogHWWa2SVNrrcEspVwsooiFIz17JrVwNbdHg
U2jeFE7JZCiOuGMpMFzJG72lkCO+E6Z9h3bQmCymObFL1MG2XbLN34AJl/qf
8jUL314iznuU+BelU0ywnX9TPBM5zSRuO22VDk7WS5CfIl1CYsIFw/3AAFU6
b/Yf50IZpRk7SDS0MuEBY0V7oVm7+EReT6TASIrbpOV7CnWFkzyk8+YtpPbW
r8Op+K+Kkyquu8rUr4S8CZEPdmesP7T/0IXkUK1qzcL8B2Wh1nlgRvrfZLS0
F71YnY9CH5XLsxstqMHXsD09PImunIIdK//NzELcwrotC+HumQmt45iqXuvA
SnQrbpNFclQFnDxuEKJSbLKcgm+I8t84yagJhUEDfuoJzwaWETvjtdl6k1n8
SzU77VbM5x6TttblhnwooUCa00I24SHfO/e4koxgDGEgYrEiswYdETblvFYb
SVhP5E5qJnImHqfQMuZGPFSRVrLxvBxLeiWp4Uj7rfciyf4rkJhdiCc7fIkE
eaO0CtWKsNbNvDs/qZ2lT7/+42XLShVzBZYfjJpffV2t0JDuF1O/VjczFyut
QHjvqb0BY4SfiY/NWjg4JMmPZ5AMnvehIVaqktCzHXMO5ve6zAW5klom0wN8
QPph4tnztrFKuv35+YRDgxSSQGD32dpe+y1ksrTnHon9LidZmDWk2hKkC/wF
pzqLMHxFZOfJT9eWjerjSKiUxCbCqZZ5vK4mUdMHye37lcfYMzYebTDeaLm3
CHLkxIvKdSxGn/nBTB4ZcttzpuPmSyHD2ZCSykZ7QHfct3aY2BXRSLeMVhMg
ks4CyG2Z255j0sm3PRDvMDB/OkJPhErKZcmAcyJ64133iYXf5euYpsavHQua
hF2tOrqsXxHUU+ti3OR6P1v3uieFiFX4BIJsrihE0AZNIu8G2BIK7ii3JAOe
IGiJmCmqToyOeoZiBjT9ZDfv71rlB3E2YCbZju84xcmiK2ZrWIDQOZ/P3TWY
aY43tl+aRofcfqjjKk+X4L1VpOKwkGkOcmqW93BF+BIw5Y4pSo9tM5opiJc8
U89M2j4PCmiH9x9Tv4Rc/oF2bTVfMIdO7r88bDJiBYGJgswSiDXZFyY2V5s0
vpcxiRQG9/C2qCLv7Da6hWtiH9swVQMAz2fiw+z8Rd7FHwOZdhlBwXw2MgAT
AYVnS3Fxe1fKqqrqKxCzb/SR/R7XwPxd5JjuFJ+Wz0MaT6S+mJ6Cb+QyBlaV
rbnXXAGFBzQ8IKicU8L3g+k4zh9vW28xP64s7S899dM5r63J8SCxjd6/Svau
dCxRkFLQtujW4URK4lABZmrozNbtSUjjfjxsAQXiwGvo+XBRtCMk7r4CRz+v
CFTnV9A5H+wnjG3zxQP2DV2XL2GXVrkY72RRQoyaQwggbfLYSDys/eJN5kwj
E06xlimQib3KP0nQ0S+7dQDKqR+kYofraMHa61F8EWiqQh9/ryQW1i3H585w
Q4sDvN398TpPa+/5b/BKYvFOjPw0Bw2Y7UZvze359qiLL0iIda/0gSdxrxOp
9emmTep4+krd6D3TSFNjrZMKXpot5jkfCiUTqRmBghyyXRAL6RrLyfGNJZZm
NfY3gh/PJ/JUgXnWz9o9jSW0s9OudbaO3W8jD4ahNf1sVWsRNbEerD80er2l
tzvK6EHQ5AMbM2EBGoZqgRpHuJvU9bEeCsxC0GNBXi9KDnx1gjBIHygadOtV
M7eDUA+1mzDP+GeA+fcKLHbWhYUmw9F010RhxU4u1Htsoqb/fgaEMPHvNM3d
ehJmhRU7Iy5rzR5sPI1JOwPLOPvwXZXIBRMX7xKLs9IVKoT35QoHzUuPiDs7
D2LdSNAXkGzZ+Eestde2h3GOE7/DTsxJXRtRbNUqySA1C5W5TLBXsO4OxcTZ
B0dhDCHrfPwxY4bq9CTh7nWhlATxv7YBOaxo8sdOAVBgEPBVYqgROwWu/eIc
xSdMxmLClnoP/VJwI+AC6/ItiKaOoLGbn0vvWlcccCzXKeVyeBKk0Bi3XcnB
y677DLj94jqAZnz+YyBHBNWviJv0KlAPiCf6CN3SWBoyYcSwCyG0wlg2saHT
PIu+JU+0NHbI3QujK/4n+8DaX6wwXi969GcmV0jJYJZUq32UdLNto9YbH7+W
FBVQH7ODjxXP0RkRD+aXaOnNuiccZOS63PwtI+0xg9ZF5GlUhStHI5O8PeRr
v/of5nTMuGGc+0lASoOyJfv4+KATU1ipUgxlD+A5wXh+V0TXUciRnrs9Q2cs
5DYlQjOYZR44hwZrVF4mDpGiKoKMy9SbfQ2BsZpV7Y8NEu7/Pdv90DMIKYCv
SrqZ6As1wR0wiIJPk35dUhQKt3YCOCnWQCZBGD+WTKVRKr/T32eaKPKvhAlR
qgGpgf5i4hjOZs9wFhuuXJL/dMseFBb5mJyO68L5CJdxpua1skl3XL/uL2gp
z/XB/PnDEZ4HxSfta3nBJty6BFPHwvp4M5vE9MLR8iMoWXrWJiQX7pgn+EMK
gc+ZXclV1eE5NqSVxE1kah5Z1ifXfn1etQ2U9nr6JgvqmtroddaTeuMUXoEl
wbpguM9YKOKVFh0eq7tMyEgv24r9vjSkQvsEY+dfklOixDQCTwQdxDdw+k7R
ohcME1Ajx5yPVXKit52MZ0ZDWVeKq/HuRUOiV2UN1BBpSMScbI7BjiUfL+YE
iDEE1f4N19BRZYFF3NpQI4mftq90RHoZT4fBUYNjBURa4YdcfKzK71cV4vVc
kwd5VDWT8KKwKjNAniUm2sxaJcB2Y5GHJcH+mgsv/9wnHjMskUHb4IB9pQaN
IHkZh+V5YjtQgQWzG9hKDaiToaFXtjvwMT4VlsDsXQo169gObKv61wKo83Mq
lgMMUUAIsmS+JaogcgvlaUsCyHJ1xeUhMvTT3QdQwW8zsNr4Z2T5h+YWSuw0
ptPMv8PN6rZn6dwga4wTpGUTt9bzHienh74XqOu4Dd8yByf9P43RQgUG4YG/
61og7g3Sv1M0fsRVK/fqtNQdL4vQWKTg2AmggFoHmo7g5Rb0UdteHeij8/VN
VN3Aa4b79FxGHLxs32CLrMfT/E3MZEjDrCa0bSjbpE1XTO0g+h2ziRb5QJoN
hu5NJxLPrqhP/xYLXzm6pzz9ziCM3nqlpn7QK4RlFYVZQc/CHyYInbtmnwX0
gJti5U5jo3ytyinj5WIgEoTM8jFHBP5xGqIJ2eD2x/lGt1Ui1UNEpVL0GTZx
sMUTa/O+xQ8NLZfBS2Lba8Wp+3DgaDWNZSOfLKC/5Z6DrW4ukzTn3/tQyzDR
dYh/b3VGq/XH39KrcxjFHhG1TmHeXSsuKdN6WPUP9BKpd0tTv9W2d7oNW4tx
elI0drrQh0UB95bNmbDWC3r71eVksF9K28fS0abHOqGfSx9AmrzVVHobbygv
do8sO9wpV6oqpNwdMOOZRs7W9KQYn3msHp1dZ080OBKcsRHWf4Ce8Ej+peDP
P5PDAAFMbnsauuFDOS0NECXN8zSZE0pECFUwDubh3DEiC2UDm/2PpJBU967F
ZDv5WGlZUUZPPP469cHO46c/F99AxYVzaOo56IDRuwGMcN0F+5M+F0R8B69p
M2U4zz2GXgl0NXEWGvUK56/5vyBcjJ122cLQrPDbKi8YvlWaiqclom1XmUvt
VN7QIewib/i9G0YpieJhN7OUDGz3lfjEWuJ+rSLl/4CE5Op65Lrdr4PpwBZg
/kfcR4ADhdpzEeAmbbg8/acba+P0KGslSmEqv4Jvzanv7Q91bbkoQL3zOXUH
WCDM6mvkcbfDk0PaaseA0RwvPkrfFDUvJKUOmqV6yb+sycW3pKMv0sgMIK60
pYc61aWhacM9v4YZHhkallxW2J7xZxopSXWCxYLlLDl2MQ/1Tf/cMxHyp6pI
RFBziqsQAYn8iGN+/WDf20MlqbuZJzYfAz4vrSJ6JywQsQ9z2MLplrlRdCFk
T/kdfE6ROzo5xGtsHmyynz91/8C+6jHD33EhDS8IqFSZ+ganGDyZbZYBEfvJ
lC8LDkAFu6GLb9DQx1bwWamXn9IFtoEFuVUS0sPM7VsHkurTHxqUfVQzWI9Z
LjV0gc+YZ23Cns9EWTMMR4ZNTH+/mJ37TtyWEyTT6a6leCJaXqNa458NIaLX
fwASGhOpIf1wHKTtsatf5R3C/yy6NcAKThOX5QqhXRPJSdDPSH2KIViDprPi
9jH1lMoZMQa5Iak3deY2jzpK0xPNtRLzromRjLFm5/Ts9MDoRFWnLs3IB8Y4
0Y1KzMjiF6lJL9qk/eGyYoDSZ+T+Pzqqd/qqORRaWpoIKINaIxHFNaiA1E+7
gEzEakJm9IIN09lkhtxFAWRROMmeuI9wL8Boko02EdFZJaEecANZ0eQjTqLR
5MtrcipHyB1Ke1LZg6vGuyua7nX3rOjbMq6HI0N9ceAei0qugx2whVnvpLUH
zI6NXJehjHJ6kTt3EbfG+7iYU43CigO3drTN2oN+Ru8TCAYeXM3lsgkE4KVe
0Wn+10rqkuroudSJuv1j90/82N647pLXLyP3CG4VFe2nh+/sfLLWK3CL5T8O
6eSpEt7MSqGEjaDVJcgLyO2deQy1mwEK4YI62pRqEOdLHdi0YCfPftTGsH2l
naaNt9UlNuvBAp+vVO2o1hSDxHG3rbEl3bgVoIRkHvOHv6W5c2Q0mHvoc3oY
nQ9qHIA6PybRcpGm8GXSPgRcMdr1lM0KM1Cc8pc80X1rbGf13YfwYxytkrYL
sfvw8sFNF7+G0plwytpoiuCvuD/yfQuD20c6fXkQSDK8+0PbAKpUz00nGvff
6ChsZP7k9umdui4HdD/Iwmqk5c+bZt+agJMlKT25LSD1/7Vs8ABsIXtljXyx
xmaVPQuuGfhZAzHecz5yYoHgFh/EGHZL0qRIzmFecnOYBt8lhJiDa+bFdpp+
d4sp+U6CWVNGyUt8OCZpR/S8gE8Z44jDpxdRsjoJVFZ9UXNWWClqU231Uw8C
hAAFT4RErucGNzPCkE1Wbgcd1lJ4cht/mlA04KCizzNW/JHKzbg1+983v0e7
Be5faWBP1BlsH+LvMPMhFnXEaX27YWBpnKCtpt6gcSW6+6VcP1tLoOaHKFPz
6ZtaF0VMxePlqbnxks9gaoEpLYEw9oNzm+u/8Ua2fvqllqOnRWYbKKTsLbb6
4aAq0+TQ4UQJz+koKVDY++RRV39vxQHmZVRZCcL+bn6zC0P7E3BdEPR1WsiI
04Pn58P037XL6YlqJBq7uBtjYyUKYDWeSdpDerZ5/mFo/wyY4hM8pc3SX4WZ
DlKHXU8pe7gTa7uQTVOY9iAnj8LP4dc8f6mKGKxJW80gyvt965zNo9eI0bb6
+eMSyUDmNAngLdS1MTRG2XgkEfXPHY2yxWyhWK2ng8+HeD5sCq8/vOSWCC46
47c5lHOWLCh0DOBsUBuijoOj0xvy533kqUH/6IuFWHsQJ8pQcGn5UqiK+HYJ
EjWVr2V1DmI64vCi6C1ZGq3CW4dGjAN8NJGuVIDNhYkCOqs9JPQ6QR0o4LPn
Kt3j85iCNj8XGT5sYMPFYNYwlS3zsETnjJEsA8wQOdwM6XYcdY2mhRPPe1+B
tFcUEShNfGa9dqm3rfWj5/bw+vXXypvR88jxvsnKrZzGgbq+5GJYwpHeREId
j2tMvcfVNKlhOunbrmhlR4FGc3bbVBPa3t/WMqA6PkVuXOEp56QoqcYKb6nL
VICxHBQRKW/2+PNw3F6PCOtXode/wvMoDyhmW/IG6ex5C/A2i3fFgYcT65RF
rLP4I1F3fMSL4VIARQsR8cKEuGe63+ZZIlxUN4+8YlWrSueHiWQNH2m51QPS
5uVL+rd8AG/cfyN+bX6KAV0/pF//Vvlvn8hAoQvBR4oJc0BO2AgWua5K3pUf
SjxEKpJgfBJHjPQjmxYRBRB06jkKgmUGVX7LeGoPgAbruak3fzcuHoJfi1vv
g3pbuFL3wMSWiUza/waDDryUYtcAXjFNuWBx62mFNrzkqEUX78yVDQ6Rlv52
ctHyNaXen2IS1ef6GQ9P2Ri0nV04diXitK1xk9ZLNUX+B6agl07LiyYbnFz8
PX8xZkvGptwWjlo8qVp3pUVR9HuLnzAvB6dACEoOWmzxu8OPhmlTiKZZ/+6e
Ul0wHyNO1ySQMElODNtUs5NIdcC7sSd+Znxx36ivGadEIq3/6eBQIcv/TMcm
sQa0JTMbEXpcYPDKLA/DPzXjXh+1HG4qFliG9M2l8X7FfG/YIvN4SqDF/R1A
MXDrjrSqTIvyE+YYi0jUlzWkL8p6vCJgGluFq6yZs99j7jOwF0z0b1vXi6OV
EjQP6YPM4TwRUGZvhzMVYzYj8IpdrDi06fu+flPfX5PQtPag8Cmqnd6c/EeO
ZhbeXnPncCy+IRYZiSvO0Zw6jVO6MPV3AdZzUE/BaHjlv0Ru/V1tIUaSwVzF
bGYPyrc+6TDEoq+zttJwqf3yncn7YfDh3rl7COuUQrneXfxH1LXpRq7W5jm6
0PGDLMLjrU7HJnGpYYgbgbz2SwuQVDmmgRZBNwFmrzqbdF6MZz7ek55ntgmz
fT4UKXAR0wdeiFs5wTi5NJy6aiGpYznCfLRDwpToso4W6dBexrD8t93GpHvT
aa5kEnSP97m3rzSR8ThxZVvCFORzMF6X5b4NVRVQa9toknIQADmEmuCIRCf+
j7aPknHXT70nQuMH1L83AMzNM6cBifaIFGluhQKp/NZDqMxfhivZPHKWEiyS
nSTn8iTJXG1z7x6ZXnlAzyjRG1PnX7ctCY4aluwtA8BOuo17nvYpHvnlVv0z
jhD1aA60wV674XPr5LzQXa7jbdCHMnrwwr3YZgNSBFA7K5J3BhydYcOaucYF
7ksxEa/agXpZyzGGV6mjx81DniKSu0oOl8PGqrHg50b48vqjJEtMeIoLaKPQ
+VOgIyJs9+JbV9ZFNuNNcl4lu1kBMd0FmPNlYST32IxrgaB0V06PXq1htuVl
uBEIz66Bj5LOKGJ5XHuMWs75Jk9Ilmw4drFVcIak9hBpC0aLGq+NmlVyHunN
zfIeo7ZaWXZ/ZQauo5JLttLh3qTWx7l18QkMZ/yXDhLZ/25vpXXDA+x7Is2S
CG418qXNLj9T2nlirAq92y+fGLlzSE0qNL4IvJNsWAzy8CmQQFx2yF/S/VeP
fcPwbzq2Pb9/hlRhBA5wNqhRSEmg5yqdBjVpSOuQVFwYWZTSlo6OZGqN7BCm
6vvSr7yu4TJtYvIYYxjGr8mya+W1Xd9kILp/uIXxEjudoD4Bkyzf3I287ZwE
qjof2sK1pi1hC7HPBDc2RAEZGM/936TwfSlY+mU/Dd1BhRYI9rUEJyEgJ96K
O3oz105guej0URcusnEKepFDQmUNtqFpDZaTKuaRzXNTBw+/QjtSEqetMC4c
WVEJdQDc+lNtIjisHebmqE/PXxlDC8C47kajzgfDGiDJBb7YOrVTPGFqSx/I
KTf62Mk6UTzuNzw3ZX4R4kUSaslZ+z9ZtV7hHSD59HQn6pv0lm+y0gcyy+cR
yDoNejjDJBAN5Sph4mIm0ZS3Q7zbR8NDF9GZcidv40tLKScC4QymKbg+NwC2
2uKr0C3lB9jFf8lZkD/ruxvkrPHuGvrMWWjWClqPO+XS6sQFuDmMr7eZmS42
pBa18U/POTGw02LFQ+DhoBMAKB8m01ai/8Zk9THrooO1KLDr0LwK8TubYKrK
axD+H+2/0Bc9qfMT6EIiW1AbxVTWPo2+Vp8acwETSOBCxqo3in4u5UyRZw1Q
7V2QRXTTWkW/dJYEZDd3h5ea5E1N3a3EEIOHoFuN/AMyq6M/7BecyPqgTjaE
xOixKOVH+kwqRgVVPoRUnf0dSRVoIxJJ4ZXFzvmzCZEqZDTcILT+/KMSGBQK
x61DACetleIIIh/IClLiaCWytzp7xuEV+8Ys2U783VRsQQ5hkxgz8l8fJamg
1zDMIg8f5xNIo7J2Zj+Q/OvKlC0ol9OirkZ86VU/JAE4a3cbERSDpfeWO8Kw
T/HAmi+b38WOuuc7WPIaJxfNP5w/bnYmhOwhc02HV+c378KWeghJlfXMve6p
Z2lf66U4OGvGvIWwQpBC3l34l44nP4xc5OONp3ezgJZRvCHK50IKx74QEzIp
w2Dyc34SafU1M0jOq4Kkd7UbTdOz2rJLHyJ0w//v49FeGAnxlqgeOZXWYS5t
7BnICZVeYUUhMDbLdU3WDvabT9is13Ah2EdPApKAS4mf4h2qJ/wcYcDmqMXc
vUMuNZ2EKmf0zIQ+mRyxdK4sM229PZ10VXCIDW9RPa/yAesa13EENp9s7M+p
0u65SBUtiRlwMUGKgvhuEm+xPmdi9pkvpPqQT8S5jytQ5cZRfgmyM/2Jt8lh
gQ0gSA/7wgOPWFfaEwnsr85jvA+EiAgZww63nCZ6gdGu3rjJ8JkmDB5hBcno
uAUJpW1hNtpgi3SrMemcg3ixnhcVQh3wX4UwC2fmTfHpxh9zjBKwc3dZ9HBb
hRHuvlxKac49/nZN4K1jv7dBFFznJrbfErmfgwL6Idi46+pmmYQKeoSBcmxe
DxxtBIkFuceCz5Y2WwRSwz6x97IdcGfR17zxHjovOqqY7WGjMXogf6PKaCAY
yxK2qgZg2asYlRopHt0jXYaQwrWp/ZnErDw4bLSoeC1DPwwZVuGdFMLdi4ig
wTSwyhbRzI3kKVRlh2dI6x0e0Z5emKGbV0faT9nM1mygIre6EnJOaKIT1BWe
ToByAf04a5YbxuU/zosRYbBULkugeFWjE2+NDZ08LY1UL4Ayp6VRXyI+n9qF
vEgJ/DgFtNIQCzQSvjH5Zw8B6lRGqPaXCReTaCPcaG2Ox0AgMq2KDkkreb7z
Tp97V3fSzSElHTUAUGcE1CEOZYhf2NmTC0/LCaP9FVlMqEtuMG7HkKWWwh3C
49UvJVJV2jr/VIQLu25hnJqHpUPKY/otjfalF8ZB95mfcTvXR0geJLJkOlHx
ghvrsQLTUsXkK10NlJdiqYs4UqCm9iVNIvOZOuaF4B6u0fUw6UZJ13QOQs9c
6hqlW9yI9RQXLlcoNBmZYkSH5eShVb+0w4oPmsfyuJI7CcwVeannKb8e72kc
+tv46c7G/hI0mp9HLY/kPMBjGjcLcZ4ZSqVCPfrAF6OZVhxv+x+9+xKn//wu
JZ81CUNH7RfZxZOkz5hHQ5IbHxjMEMnZn9SQ/HCeT2BhlT6wU10XODtEoI2Y
KCaw2PJheh0lnFYMwg9eXsaFwzi+okG1D+VsfxANFgdqmvChM7bjdK6iL+S4
qwREab2Q0rfVyRxtXaWdLIoTY3M3SNXESb9pu4jLAXyDJzzEl9a2gbKhl2+o
NLA3xzADu4nA762VwcPjh4+GPfvifO6W8EmuC0AEENqaHq/vPyD2TIo464Qz
R+bf3ZYaBm2AB9T2jHOppG6xE2N6MdIzdC/YRPJUDU5ULzZCC/YPifLyErk+
gm5leNcaExwEodTom/5T/0tF3Lciu4Z9oDBWumJ8T9ZfDyP8EavrfyTDOa6M
u5B3qNNtfMgYEWE71IGOuasSbMUfiI/ZtGvIpEGBlXlyTjgFVKr6PoO4SfpJ
Nyarpd05eUNnElSGEZPBoObzjn3607oX6x9alRrwZ26wYOwCRQjL2uV6jbGP
6P2wBjtZ4LA6O/PPXippZMb6c7FJ5UZzMo1W6/oLD6KJF2mkfFC4C1BILtyh
slraFoF2dgaVRT4QpGVR06GAv+OcSl7EWZFN/K4U8KZ84SgTx8ZqaHrjxW5g
G0932zALmxVVF9XFfSYIg5blu9vQUsl62y8vsptkEdAbG9Gep1vJXDNqB+At
3jQJJudD+Oima/1+340D5qY+FK6BZmgC+7b3Qs2KHNDc+E3WcYV4z55xOhMw
U/fytd76hBWnGbjEeECaZ/rjRvTVrbX4qpurxaSSPIIzMkOTATQcGHlEnlnf
R4/ZdnHMPQQ6J5TYsVOovuLZap/p3bPpEShJoWj4+joALy6cpRSErYH7Awxi
X7vvw+0NA/fr4u6vAlm4ei4uQOb5INYV+6YzWfP4ATP6SVJpqJdxV5YSLPfV
D9qGwZHikI7k4OFwzMatP/QmcQ0gQkZYI9gEEOppJC7W+J0tVXeJy8Bn5Bao
V5NCIDBJJQfvV8sp93EktPtbgIQB443X6hq+tXNJCxl9QKuwaM+EdJvjh/S1
HtRPrvlzyLoCVoLa1w0rwB482gIjkJ5eSGA2QF0YrCxV+udli6T8LMiDvDVi
RLfLTXMrhyIae7qKyew0KT8SXnoJaMzeVYfaO2BxAhRBV8H07bGIVvO/UEAr
RmApA4vLbuD6JmhSO4cyCJHPSL3Vn6x45oEuxPhryPi8U+FkWU7AW56nTA0l
K/mrUTgJIBzhUPLChWlQGRwmP5mJNPgSj9MR5qGqWM/rw8n1NlrVFT6LR+qB
b9cz/BEP2D5XgyIUW9xHFpgcMRBZGAThhprys4pnzwjI6YY6MZYwLsQ1S2xY
BSFmugbvXKyotxlSSfmfQ3bs7BuF8iNmAaNMlltUKcMsUySZUzcZuLE2UYzW
8BG1LLKJxivMJC9jlL0Ki2LGd/P7eAs+HaUlu/rKSG5rw0nTlwmWctawWw/H
KBa+XIQKcXmJQb8t18fSpHydwNm2pDLyrEAzAsNtHYz9Gbog944nzkJk7nay
QD+AzaDbY0+hmTxoujNj34pxWkQ+7KBlh7BDVlkjO1RCgZXI1KZimPxDmX0G
ZV9oPQ6Uz1CNqMrCJxa+qrtwmQygWePuqEv/b5pl3z6XbqWE1V4Jy4rIx32F
m9+4SoP8+KfA1XJM/Df93ZnHURgQpDYfW8r+KsFEj3kcK+dnKnq3NZ7hLs/v
VUnTDSTkdR9PeqeIKbt48YZTc4UDFxa9qLW4r00ERCP6xL8hi0vSfmTKcpPz
r1INa/O+aT6s9kTHk6/0NsI0U0LK1Y3pvOjARnwew51IO1W/e0Ylnax0Sl8T
yToSdg5WugghqltlWa7/sLaZI3dxAKgxb560kePBrVJ2VJzuqGqa4uTrw8il
Hla1ld+q/SjQ+bmlrwkZIBbt4zNEuEQfw6oxNH8AKiylap26w0tq7ocekNGk
XpduYBIv0osb0JxhBM5dmR4ekcRXkcm4vg1ahr5insjLiyy/aPDrOrNUXmnq
7JaZF4FXiVGSrKy4X42glTyJKTR1v7V7Yk3BZIaGmA3vDtnOUzZgT1nAS8hJ
v7Gu31UeZ1x5npMkPxtqBc8xHhqjuNxitQk7j1r4+pD3BAAHshjdqi5BcoWS
Lfz5Tf2yMYXuXFJ9TDkUhvtl8muam/rj/3CZfbeaeqJL9lbn28DKg+MfELU8
A44VTuJfLdkOVH9mvWnJLaWJkzeMPg0b0oaQ0kGhFH8DiInL6dTTLw8D3NV/
JowmsHDPK82u72/rxjPSaiXHIBm0EIyUEo9FA3W11BCtM+B5ber1LebTRvn5
CbOYBr6NvTTLf2a6dhpKHKEgel4ZUvko2XByx6OJZ1sSjaHX3MyHdB+kf22X
tUjMCiBA+TXLxLOPAs5r2DPJ097vJSre8ueqPiHnGtrS9KRzaM2Zoc4+4oFj
1YpkewuE6uA+KryXr03rB4Vm3xn0aBKQ6mpThvTknEbIkNn7it4iqLFBFz8j
gJlaL97DvTIHMcFlaXbCjw49guN+dQP5FFc6lxXVW2tIOcUtjKnRlvO8fbIR
+oEQlZsKQYk5UsHc0/gT5tO6r2JyKXq8LGHF9ntMPPY9SE2ZaOzs/Ajw/SDG
Ni9oGpVQuY2JQzx6pXlMgDGKnzcf0uBT8Z3MeCKmk+iunG3GPjfNKYs5Yehs
+TsCcAMquV1Tg4/hFkwPy7ALK2aYQbgNISD2DK1d8yPhOIQQd/y0MpshgsN8
WVmAmGQGmCKqsl9OZyruvCLVkZs44ocJAK6LD4Ek89I32B5GsKfRxVQfnCti
IDvpu06KjFb2SUm9scGXuov0PRYF9ZXxQ4W/+HfVN0f+1vrsgMFPz1yw9b7S
SUkM5VvArbsJQ/Pff6XyXBs009MizCU5c9PEXhoOM5B4vGXTSRqsLj3k3Cym
wjpQ3i+C9AuxW3MgVBZvOEZcD8F22JZTGgPUrWc614V3kqNLq3wAlS2jXASa
YmhscAuAh/etbShK/ninNpeRk2hLRxzTnav+j7EbzDUm8Wd0hMvkrBFjdmOV
pKjjaMC112groP8fsuQhLNYzP4akWDjGzk4B5h4nRH0ApLsonad7lo97w0+P
egVwYZ2MTMe4kDretyiV1HQfdYM8yRDpdxcgtZtgrfwnNGrpO67XCVO3KK6M
xlATwQD1f7oRm/g8/ltGUravD0FSKDjZVbDGodO5ZarSz0HAQEjiek/cQgwa
uIh8Ma31/VMNI/BT9GcLWfi2cdHSUv+oWVAxic9WUOcmB0VqCLHFOtmrGcRU
WVHTdHm0r5M/d6UQaVLT3KOi6cqQi0gqRKA/n012k9jT/Fbf9MRsiHzOFIkd
H1rMRUMy8H3qM15XJZvKYNtF2BTU401no1UCftsldbMd4p7KratIkEDi7UEC
7s2y13DGQQAFeqr4AFNBno737C91aXxpY5PPpL+xcl8gntoBi6vDmz4bCRVb
jSUfAywVP78T2kNmQmp/MZi96VuhMq/XUvMH/Cwa6UECTggoyVT9y/WTS3T6
HA4Bxi06sdF13ko8h6t7bT75mEevQ9TLkMWI1Aquom6p78PX653y+4bvPl0p
lp2T8B3X2sq2LjtpoFQqRjEoblirKxXT/LUaMhIys4DK1UuzLrU3XrSQzT/2
L17z+IxfTVfCNTet0FQ11WNZLJ9xmlsc9gzBeaJzvY48oeXqwK8plavFm0rB
ALtU3o6wC3pafdmJIS4CSg3jlqJ0telsg/gdo2zKj4TMTHuLl/Rc9I7b/nmU
mpCnu2lzXxw0MJ0Cq1gDBHB1ZPrUPR+kL6tTu9z5zE75l1ucJwYpVdelO3GQ
3XGpWgpKU0viL82m4OAfDYqdrskbVn3Qj0T46Ib+MyEJoQYG4iY4AgRV1hS0
5Kt3qgbhBvgDlkhD2XwQuqMXF+YcLtv/LfyE0u3NeUjmOFARayKiljpY7ySK
/Ldeb2uSALPx5jc1N/wMNkDFBkFKMq1Iqpo33V713RHjI5Xvmao/+r5vcwJ7
bhcA6n/8WWerIA/V+LK0hVyeMesv3hg4Zb2a0si3HRXStFiZ8e65RwrX5PEG
RB7/+/Kf0M+9eM0BiTtfSfy21jhB+1gmBtzoq9sUBGJonFQadssM6023S85P
c9dweBtCOkdaxkddyvjNcBasu/cNy+dMIJb5tdqWUXgMrp7oA28aIK+/PqFv
16yLz69ME+3Q2svsBuOKv/PgJpnJ8OCm8inqZzpkJ6qHWm6ewfkyadNIGNAM
palSNz5om6S+WGozsadNhc90c3p0V3XPuduDXS6W0X491JtHJ1IKqFxY79xA
/NF451rN+saZxf3u5V28xeTylPcf7VPKhk4yBEEHL3pgCJzC6xvRR/dWRN+q
QzbeyT5On6a0U3FDVhNomjFuyT0prBUGDX281cZhiP+e52FnTrQ7QhSHnbys
lUmAmAOISOw3fsIBQxeNKS+SqPOYDhxf6O3pjJicMSwzGka243QUH+1paBTV
bQ4Z9qc6swHsqsABfSGh90M+jSe5LwoI0aI1D4zFctXHju+RVMO21nqkF5WH
6IePBpTjAry+GrlCkUoamYnGi6Im1q+A3/ui1vjIvP9TNV2AuQWNAYSMdMwB
z3LJ7vJjN0QURKQhT2pIQ0dv0aVL68mQfbOvpaREEWNhIcrty+sypQU2+vun
iUMta68FYGudx2T71k1ty3i3p5XeUIpy5cz4w589X+S7R8jI7qg05KvTzjYG
nh4p6oHudUwNKvPSAwN8+XGq757KfL7NxkqPF3hWb4Bi9EU/8ZHdI4Veok/N
C3xQWtxEKdS3SqhyvdhW6a/zq9DRZoQvMN8R6nm23azprh7gfWSRDCZ5/FvK
IMw3lpaN0f89gqPdpubK94t6JVNADoNg90Qcl0Bqfc+q9X0fuesHwLCa38YE
P6602qvr67yPRORV/OmU5QbqLdNkrBN8Sobc7dE0dScmY6gHJD0Ju96sJK/M
RoRUkfqIVZrgoE/EVQSU3IM9+sCxOIbpvtWBvGCvkUmCEVqceTGdsR32erNT
ujokEMCTQ+AU0EryXPrf1shCSg8YdnrxQ3McbHPAC+iZG+vG6mk9EEPHC0Ap
/LiGIO5bkzmBil8Xl638r+GGiD70O7wQN4CE6vqz8qwQisre+9c2oQWAvaXU
hBLx64gXOBSzLXIBgNw3FfDBvLxr//nq9yInzzY/G2ZNLbECiB4v2Mz/giie
ZXznqmXn5oeKCDxBk05MxEd7eelcApRZFLbhF7fETwOg81RFTFDouJ4M42et
Fpw14KcTqn5CSiVc9zx+u3QTeR5z34UG5RL3H7hX0Wzt/Zmoa1un5bXw5Z0K
DdaIaQtcfrM9H0xo6esuGiCWP1cZHja71GlbunyRMjqlhgf02MVA1ivuq8ne
w1NM93iFgt1yJ8W2DpXtnvuNUnWPtVEPNhxXoMg3x4kkk9p0txmqzUBTPLa2
HvHlqQigTpTk/T+pDtMH+zUHQUAjUr/Nl4yJA+0QObp+4DhRBJzDg9IIHwop
/+SMeWYLn54+8gSurdIKEYnsa6O2QYDHzkcKHN5XrZ+e7IyNNYSE6bBNG8K6
zh84Wdv7nG+zTB8Au1MuUVbHabvAZOQ23jHtrdoNhzIJYM5/+wrwcyErXrzu
OH3AaX1HkDgWKL6fsFENbQWA6cM+2aV9Eb+FyuJJa5wOVPf63F8Rze4fUSM1
qnCzXikR3L5TZFR3nLdyKyT1vC/1oIA2lw0kVjmxOqj57QDaJoQYN60ZuiPg
U5nOLIo+O6LvtK1vxr9XIgFC4+RZT0sUJgaVz/ktEXnDMrg+d1tTyjb5xOII
3x0cUs+NX4jXC3ZK48qc2Q2GOwXf06JcrwssJNZohnsJnS8wBXNGqVUGj1DC
WXAGNBXwgzjgqCQBy4twzgq9MR2PoHJD7htRJ5HZQq86Rrz9WnFiy30m9lLr
Vxp9efOlqo7jn+AxGidU/v+HZcbPkrDxxCsgmg7qpm/d7SWeDC1CjN5T7bYG
KRuaJ/NmZPvkQIH8i9nbz8AGU4qq82ZNtjx5mPQEPpuAA9BuFWG4YaZuKPUf
x76O9YVmJPq4HqlVMse5oMACfL8g/aDZ13M8u1iS6HvzJacYH4V5med8zJbR
4nRWH1qCWd1rdl9FuMiaiSk8og21QNuaSb+f5GueiN/5c4U/Qe2BSjEbANpO
KxXx1svUu11mrmU9tikdXfkCjdcoVu+1aLBQbgbtI9qEmPKmQLRwBlSLKogM
RGWImWTj9hVndKlY2fR5YLLLKjlTNbEQ3PFEtN51hMUpqtnVJwFiveUq6yho
mAgRr9bM+lmjhXXMW2isL8hrk1xWYU5KgPANI0n6NyBuuPfCa719hxOqhULE
4+PskaZkdZ6Nnz7gaCMo0l8vCVjfBYZose13UnBT6MGO+dgShQCYwlBHkl1U
RzDFqxlIbwq8FoI27aNI5gZBgUIjgIk5dDRYBajAZnh8KaAz3Zy/4MRSYH9f
O1Jr3ea+X5/bYcjsEtZ2S9GrVVV8W8Uicy1fg1s4Vd+Kq5pSTWG4AaohbbAo
BtRyb2ynY7SFtpixVdOg2Hl9mer+QMSDm9xG4+zCSZJqbwEMW+4DjrUykKiT
PaMCaYTmwymGrkPJnjTRWueDj+iR/ztbebctjTVKSk9it8074Ahe0nEaAIhh
JTvplpLYf5pnY3MCovlkAV5Dp6lEq+9nyg1OiBUukPbpROzVUVcBszb9HpNh
LMH6aULjNWUqm7tlTIBUVr2aLuFLsnzjo2lk20o2LB0an6KWUpRf9rlPUgwJ
UhvJS5Ax0CcsBEowqccuzTS/cS+SE5OmfiTv6KmQjN9TsSW8of3sM/J/SUBl
vzR5n18bxQB6FMU6CoMooMevdoyxURVxRBp14n92ntuNrimpVkNPhFrP/bgz
ERnwbqu2rulrsdOOe33OfvGJydullgsdSJW6sVP53aGJaaMIeJkfMQoAVZGi
8sNPxgRGcreEPx1SJTlTrMz4a4KN3ZH6tBxHgQnN7/yQqYvTBaZb1QXWa0v0
vTyuVQ+5AdsWNZrYjzKmOkHLSvIQw6taeu1gLMnbXXvHfA0xH/RwuccY3RIM
MQ6Vh6MmiXSIh8JSI6BAIDF2NhpDZR66jjWdoPyEp3QgI8lnxeyzxMkaC0J/
JqJYWL+wg2Y6amuKkDjCodyLfu/EE3sdJbFGHJQ5UCvbngF6H1gZKj00jYMc
88g9jfJjjy7OP1c7EV1IMJzl8awUKEbgJkaTZXmKuNRJA0NgRcpiBZxjs/H1
Vl5ODJGCEEcPFFXX/1WcxZb4EzooqPnl9X11kvd7ZrPw29+pSIXdUdKg8780
gI2XVQ0KTjMy0euvqN9JhMZeRVGdn1p8JE24Rz/tEIcZrn3u5v18PbtD20cr
ffACCBwoMVvM/DGfnptmulG7xZ4kGonPSwBdf+SozSRHj4h1TDTBk9bUrYSr
gVO0D8eClvta/yncW9Dkvs05ZKcUFgFI7YnLXZhBGW+l3DqejRFtolAYtG3q
sU5VijsYkkMEv4TBz2WY10xuwlde1nAdHlOfohvBITdjNdzSWus3n0RoQYTv
lw7YMIhs73+Sqco5CcQ6Y72cTlmHnrCQf9jIsU/U4FnXl5yHrSPff2CwKAQQ
Jf9UkSJ8kDaullViMHn5Oj1rstop29Xt73aXAmNuLEaBG6l+Zrx1wkXkt+l0
yY41yRLti8a/o6LUZv06bYThJS5pV63PzaSlXAJAtbQ1Ut2/Kz0L7KKUO640
A2f1nHt6bTJbYJumtcgqZQpuiN2/TWHk9GYFnQCglAWE6TeKeKMkmskTOQyR
x+suo9z5LtRUPmwRVeNJgLTCnp1ke9B4jLgplccvQgIfAJX+ux07wK1lIKva
uOFTqojHJnF8RpxrapSGEKpXQMFvYZ4j1n0rahnVbLMen7R97YEJd7HlaptO
zawns7u4PGmpPBVt1aVpkQ+6uQ/2zw9SBvxGgmKpxYNJEtFimM0C4zABe9Eg
KzmbFKQmGjIFbpMgR9drPz3J641mt/q7eVr5ZGT5pVJr+5EZZaQGXEw24/l7
B/Kd58duTyH9mtya1grQMCBDSzb+FpgnzrQd5DHRJgvMKFotkkaK8lR6N+nm
7oJTEge+pM+4bhPLjTzBFRD7KcXQrBPmjlTup2xzsxb+WGD3sx6vRUaNWZXm
6n8hKNk6LVWX79jv0FILmeJ+Le0ARJVso4vmd9iaYBzTkKUtjakIJmpFB7FK
Nji2z4yPjvcpiZQ96gvw19NU5S7JnF9x5pISbbVfZ/OZ1VgvbhA1bDOp4QhA
yaoMaHgXWGeLYVmrA7SHo0YGS3crhrQv1MxUYdCcjsFApYbL5V7O8B2zyGFl
M+rPhRDg8mc90FZU8D/koTwgc8tIm6WWaaUy/gM9XZyTaz2dHbonaupl6cGT
AXYZCZtuCsYA4yU4xAZVpNx+nw9MmzgCHmkGeH/XldsNmZYXDi+Ay/k+LmTa
x+KsDC2YQHtz/RcaGb8Vu7eXphI+m0ACUAaoMNDOjdCcOf8C4bbbmy6ugaTM
T+bLoK41bhN6/C400kV7e0bbUnhYZ8/3LnNm/FJmbW4o9xoVMwRaxAZM2fJ/
2vUv23oNYE7xpBXX8AZ2oHUmc4OJVOpx85Owd3KED9NyRXX3c0kgf2M2g1Kw
PIbKbsofZiyZrTvECsWx29OgbSkwQyLGCZSMSG8v9OAL1dLLAeijcz8oiMVj
JaZnqf3sKQsC5CdcfilCgFqF1vM6rdbKEYPEgHSOyXvmRkZ6XSKLV0bZ2EM6
uls8iO2oJo3+LIWEEo9xTXiw4BwrZV0+AwLzymv1qL6SGyGnITIq9QLm4ilM
QIdD/5d5OBUTIlg5lGhCAhP4vBX6EN6Od2qA+P8AwPsV5Aj7QvZ2SZjmGjww
otGb5QNUjC8hjbpnA24tc9MzDJgfE5uCFKU+r8HxqXujWlGe0EjqRg91nrrI
zP3cJGIvxrPgD+3OyZV0vAvhyj6nC4ssiAsplhjrABKLoduTLmTIRfR4dRBE
6EXIvf1ar44/a5r5kS8amWGHqVQFrIZ7xcxaxMmc3zTeR6fgZwdTRtgQBGpm
Vavk2LB4eWhhI0N7PyD1bSUdQJACQu1QQArbwbDlw9xu5RJKz5kqW12SbK/7
t5yXwiLPCye96mp+g49jaBOQIrYIetlQeCRSkPhFfreaJYc5hffJFPrVEBLd
KpfS1onRfAyTaugCqkhJxxkVqdfO22w1vaTBYr+iDq2C6FifayixJsrjekcA
oWvvkROxEyKrqs2K68/rWGlErn5IZMAz5gycHUmDPxW2p4cvww/mSCxZn/xZ
fC8Ux00fvbLbxnrYYS2GJdHi4FLQ9B1pq2P4azNzS9ZhEsmJQS7FqRceOaZ8
29JAc2Vn6icqWsI5ni1eLxT5ktAtpPDm3LK/sEW5YbvALKLLzyL0fYYEUYEX
tzi06YTaJ5FcvSFUZKxn949372Kn4xYi2T16HOGqaL4y9fdzMHb5R94MiOdg
YM0wkkHQ7JILXXQq0ak1jHwSHYz1hSVKZAqohU0UNi9iIsdN/1s2peV/iEYS
21nZP2a2K5WZNxmFhOUesys2u9XlzQ6Kfjlj/o0TE0rDnT1/hTi1hX6eh8bx
mcSTTXZW4/ha7qd3OJ/+Nmd6cF0NwzB6f0Dhrk3zjEwxMQKYoWDBDHJSKbV+
dxXjfsubZOu5dhBMyigNn220XZe+LHOJFcgCxFH5MzNTdkCup1Q8ZQgoJ5fG
Sroory7/V6N5puXlUt/U1QEv0RYGp0sOv/pc/FAKn+3V7BcYCqphVg2v1WZ5
Qg3T4kGdJjQ60G8/Or5hbGRai9eeTUytwFuQsbOa4WkgJgLWYWZpdAxkvhej
fzHlMPKRXY84+mOu+TlpXOvg8GPTYGpnk0lt93UB2/YdW6S30MP7cZ3AHUSN
h5DjszoJoRYkyWT27bKmjvFONyr3zXB+O+XHr7IgTzI3m/ZwFnGKbBHNDuCO
hk6G5vQeHGwQdM5g+ZvLLR4R8cRtjUak/IYItF2GqI1uvSEk/kwTtKBU9fxn
quQTZizCmjjVOG1zvLQeCt7CBsFe58AC1+F4X6kYoKz9p9PqmGuzLky2nPS+
WA8+Yybw/vaUT/awZ1DUeYUs0sTLHgvlhWbpA5LDwXCJ21dsqQl+7Rwfmdo5
SAYqaqVRfLRrrKI1gmF6EIvpNqR5zBkPy2GPcyZ9OeLVknDrm+e04ajnsLbZ
A/Pj14X/2w2Kvd/ig1EBi6LKhApYHaZ2IkEZWMByOMwhzxNWL/y9QJHURPSX
OBouDTEkzrw6kjYUdwvYXrSA5L8PHuE3wcZilzvuwwC6pFf2uk3pv1gyNv20
hzKrLDegy6v6KcrDfCzUWPYWPuqF0VnksF+dJZ+kOmed0wiigcZzZgFaDs3q
E6wDrmMV2IlOV57Gn/fwzVxrM7k98OUBZg691dh5mmEWk6KGf8FYqPwk/PYM
I6VjucyhvZ8RA+ZlRbgHnTaPhqiOQ1YKzX5P4nUXKFjOdwDfdOHWX8cmc8jp
wWKpktXQ1pwMvRg85670U5d0kMDKNR7/dcwYeGoPjxQuXSvodz4vdzqedGda
oi0FVkJnYTvNyJhqByGNfSk92ci9jdpEK01TbgR6eTsniNhLZaege6Oq/Ev0
YE9kBfxUezlckSp8w76OooAtspF0eFyUddxL8K9nkFTFDQlTE/lye3BJEC0o
DRuBmlHBhPBrWPBoWZM5G8EN7XhrWVzaFahDv1P6zNf18V5dHKtHu0cPoZZP
ukhGXh6cBJPK34iWDyi66hnw92tz8jJNDykRQxNCOdbmHuAg/6FeaCDpP+xw
MR3WnpNYqxdKqQ+zYheQgOP5q79T2gJgP0MiU/19KKZtAS4ZO+eC/XrnzA/9
yyjgCTKioSFx9BjvQhk4FG3LF8XyVfjvXVRAKURuXTvSkG80U+OhUh20p1Pt
XiTwSZIt13hEgEvRXKl3pCBvqyAMGXchS36lFslDwW2i4NL9gpF0Z7Fl8utK
caiPQ16AC/Bw5/nRbXRwZ1EozvH2b8fkAIlfF0HWEVabOHur91XXRf0PqB7p
qKLmhvS5gcBCgAocuOa8a4peT1cGtCgWv8MuPoabnvG5f1RYBT8cVj0MCbXH
BO1V3BY/7x2nzlnBoobjdoiBI3Qa65tJfCcRQfiwcLNUy6E0hMNy6wmrgH26
AoNI1Vd+mwaod/m/FqQbMewsMUAF68LIIjP7Kq7x9PDp7Aup7gewkfFlv7Ft
oJ251/IOuSFn7t8qXcLbmLkLsf+iZLO4y6TLUrxI6NXAQ1EMW/YKZL04hcKy
XlEcl7VSFVGEJwtPeedJPqdPfiOPnUrt6D5GYw6B3OkBTCXM08lKlTpVsgdE
eYBfdhgywvG9tbDwGISZhtt6KyM8OWfB5WlFbSn14CyolHxWHj4bLTeVg52t
IK2z6pHYfsFMHeb+noVcHp1genZC2/fNKOtXRZetTTR1B5SSetldNgNsz3I+
QPTQwrWXl+9HKDBo1UEd7O2g1+OkXMk1HqHOLf50xUr1zQPy+6RQzL0S7N7v
48YRnDwlDoxqeScw7qbqttyxSrVlGJlHKr1vaKMMWY/SqrwOr7RsTVe1ELbA
8Go0qTIgW7d+PgyWkS71Rkqrcdt6WM1hyyOCUmSrYnX6WjVNHY+O2pwi94h1
rqHItMjVcvUgYe6FZ9nB9yBCIR8OBKuUmYY0QSU4EM/npNGHgOhIUP8JqSfo
24jFAxYedT3B3LC9KYjmKcs5BgiRO0z178uZY0EOIK5P9prWCV2YEXYh04dk
Yt+V3WMendUQmaQQKzR+/OcvA6UWzqnC0oRgZHqdoOto1OAI/OCM9bv08fbc
HHhDnCGfLLpxCrUYmlBUCIFBmUInxSfxLYhfBpkJyqRZ3lbK2tfCd6VA6FBu
e6Fc5LswJrl++u7A39em+D5BXY3zAiulv/IyFkoFzYdRs+84sg17xrxyfdS6
+QYKCHAswpFZcQh3PxDCg/TAT8OujpmJLqk36iJdRG3SolxUtPp+Gmx15bwR
K0u0M+C3aXkxU60ceMC+C2kW6PqbLcmF3rntq74AVDOC4S6BjaZF0PGqFZvm
BfDrND9KMNi3/zqIr7PW7sS1CXUJZ2ljyZFlTMSTUODiI5XyA2/+x/bSSMuJ
28O3DmxQLiQt8kBWxYJNQIwHXk1oUWq5XjCgPZ1aEtlGrfaSHhLg2h7vgnUG
UCJVOO48iGKzYsxxS0mMKGXs7SDzp9wLUDcO4iREstNsBmoKUh/P3XmC9B30
jm8+aOh4m+YZv+BYAAj/+WjNW+JbeZvQT/0rDNfynMoBFmz1yaND4M3149Y5
GKy/ZltP7AG0YhZ3pb9Y8EwCuAhfR6QMKb6vp/4OUBrpmy1zGemhq395NzQ2
W66PWkYdCvmqIdS8dAaVRjXaGgAYCAu2X0rjrZhjdQ4uyyYoJuBugL2uOfSV
e/aJbyRAKPEeaCnVyWvhEyriEzrSizWoUlVnWqRo2xLEkbR+cwX6WvemEyKK
ARzOtK99bqvchXMw+kizmuz5+Hfhbz/yuDs+VHrfq7NPpciRD+1cRZJoN/ad
byp+nvDF1iobVgHmakjrRnmf1uyUQ+LnKpOgLnyrNhGABqrmTOh0binaRfcs
Rdz3+P3QZ7xd1kQIqQFzEw3UVq5h/VMTlKm+97cZ2EoezzpWRlFRpBMiS0pA
Tly8JaCedStS34iuou8MB6dI+2vO7Z7HjhVz0oynH5+NPY+CZG0NNqkVImE+
J7yxPkqqG6148GAHDPoD9kDJzeOAdQPJIUrtO1RgZ71jEIHyApPpvhKKobhV
ocSlOdvoH1IcfNR8fQ7czjQDwqVnqnNtOtoYM2DBw344m7Hbmi6tcsz6MYX9
rTDH/Q+fsZ6vmdqlzUeM6Xetbegxifqj//itQcwEKhuyiKhuqYiKtzKza0LU
vJSgEQ0vjhkoekCLarjY6SlTos/00DlDKgllDBEnxAHX3gMOmkPox5WVjCnI
o9cPflj/iZ8/F+tY4PN0C3d/UX32KpkvPuvoGT0LoEZQm0EgAmov/qOvrxvH
MSDr/KQwru+MMlnMsrgulOTYo8V4zgJ5q3Pz7sx00lyuVw9mMFuPwt3FoHhf
9M9g7jyeBR2h+Debiy5fa5iiHCLgbq1W5b1gNQU5jeRt1FCZnQhl3Z2ZTLVa
v4Zc1N/TvbmQFQG1VDigkKpRDE43RHA1ALCbRRQn1pfX+olrRU4/DUlAcwwy
O2/Kw9JC3cYW1hyVq0S9M1VsE2rEzpHX4AlihGCsnYHXPJDcuGkfKKDUa7tu
d8aMQiinBM0ZO6B6mWoVVApeyZrtflnl38NaRs2LWCgRAY4JtPfIIUYwHbxv
CiTZmUktq94sTlfSaLmiSvBCxCvIMoqXldMc84+yicIDUDPdQOv7DZu0AndP
dIGdKNJamO7CFRunmOqdwUGF0yx9YmC/vc++C8jGjLNadPflnwjAiqwZ3MPW
shNn84LEYlZhXQxKPINa6Ky0/ScU4deutw5o10GhX6Moq0aD18rkVxFOjJaG
ETsbEnpoBDpb6jTVjJKPwo4uBizah7eCQg3bbPqXLn1dB3BxMIOyVh4l488z
yJXshK/xHb8EZLnjeHbT2YhoM8a/EnUgPEEvVqNRy7yx5HV4j5sGuSVq4LSg
Kwt4GwBon0xwPHxOD4Tf7anj/63wFCVxkFPFcWONuxM6hpZnlRUZn+flQ5iY
QqFiJRtz42YqjwJFcxPjT8oe4h538h2WEVuZREsml0l3MaelO6zTqOQCatty
sAMXroZLU7TLdJQYzLvZKZCIORDFSSeT4m7S5g8NHf8QxxuD4uzeqbgluCt3
Jatq7LO1WcK+EFwu5I1V9dqsXcr4oisxZttgPGO4rNBHay3pIpL73zmc1kwe
1ZcVd7YtTlM05ebRqb1I4oBCaBpyDSM+6j/XJ50B9KUoWugazRdtL5fMyRY1
hqpRFdSRG4mJKd0/Dr/Ri2FRoC0rjA9lvD4+vipV/wmt/WlAwlkIN021op+1
N4SPbKJr7mPSEwD6v6cLf9jh0kzI9G9VGruevVx5N/Kl4RdXAHTqYY6v/gnW
gfPFgU+NrEijDHlYXDoOuFal1gVIlZRdlGEHvCdzM+1A3mQ7QKOJ8lHL0PNb
sA1U94ZqajGtfXlXypee+S4kNTG2e6/8+yb5eiG9Le5AILp2JpAoOkDjZNH/
VLU5QQKN3ESW2IzmbBMXL+r0tP+T9vHOQIMuefnbfXziJelDYcdacaADEYfw
BmfTPuPuZZOIOfMN37rQOlSjRCWhCngiLrNbk4pocYnXIm92PHCc+RwHbOP7
Lzg9e6JAxrPlnYGQ62EmjIBpTDf8fX8pCG9pGKjqCKDuxGKGssFEkHXLyel+
QyFXM3bTDOq1ZYKnqjbnZsS7Z0BZ03kVUfyoU1srquO+WZZljswX+InAZ4ma
QQpZ/Lnmux9RgxdJ94A87RCQFQAoiEkXpk6ziWUjxdsfkPZ2tMXNiREEbc5B
2FMANCKFthKUlPQKs9XZnH4XVjMNCoexK22fXE1w6twsUW/Nfo3GIQr5iD8m
71p9QHRsezLFfSX52indqRo9vYB234LJM8bN5ZYoZrWS1StQ/g7Dlq2uVc81
ko7zoR9usKtM6Rm09b/mjo4iBgDP6qGMkAXM9dRkWpB6cUgj7PYoLTkDA1T3
ahxKwwxi965UaBzf9CMekbJGDVn3rwI0rUQu47Yh0GpzMGdK67j5Txp5aHwX
LYM+QFE4PtgfhJRP8VPWfIrXhsFOBpMvUZVH6rODpxewrF+X4N+MlqbGNZar
/1MaJY0j9L4LHjGAg9PbEd2C1Aj4z2VxGAIv3x9U4aFH3n3N9osQ061Du5O1
P4VQkaLzlzfBdBUffxBiRpli6vE+KEd70hnsZcCswMnqvD9An/zvBSpyq5WU
4F1gqnHIvKrk5L6AiL9czbu3JDj0KpSw4KxB9Pw49SY8GW3xvyN2ykr3OsNQ
IjklzM58k4t5XBJoyRyI4XBgykwdF9UC3yAZMsZnAL+wiMUnaaIypDKRjc1Y
WljClDWd0c1sB30O+BtS01GdzxYjS25RqFcN3boVswXVNfBYLhO+AuLO0Ztx
ybSUCFc/ob/jPt7e24RGRk6kvL0JefF/acqgaEmUPNaKG8nojgpaESC+RUHD
ueNnHHziSrZc713pJAmQEM5rommYTH/LiBiKM++j5/Ih9iOcEL+YVwej6m+a
v4Ff1vQP4xvb0ulH/BF4cPzO6qRoR77bfJmcVwg6W799UhJZbpIoKEajWVNb
z/mTw4HHsY/OTe58DhiXLEcKLlbwfw4CBhtZMCl2rIOqMu/t0wnNQz8BkyGo
EbwUZ9F5+FiHk70kuIn4X84TairmETR/L7awj54Ypqxj4yZ9z+t/u+mQkD7J
NYCwXDvJCH/gfxgmd6Etw1G/E7gqnqbHI/3kSWjTpSWluQNGFYAtBBcRwc7H
moNl7iXiJ3yBWOulFhXTqkbPPOId0bGg/4a5v6FAYLnKPlYaHGtSZp3chayx
mIprqJMpmW8foQAt8Wxjh06193tdGAUGfHr6YtW8B+icBUyg+MHklnPBsmOU
AKcI2uQf3BgeoKMlCxRAnVBDNKiEINuXoeUI8XC+/yYBJp1hpbjkhBEurcZY
Rlhroh3FNcLvETCfQbCoVUyANhXbfO2vbXE5cPgGYOUWijt4ZMTRFtWyEfcB
DXeyMtKogTTopDHDzLh28Y/8FUrSYzAMsuZ/ns7ukVgwoFKwJHVDCCzPR/NI
DIYZyZdEtdHhOBzL9mzn7lB3IcHauuZZ+lRN/ebUgnmK0gmgGhMFSdK+stOc
RNxxtXohfia6QEsM//MmC7xeSYbyiSWIWXkbO41pe2qFvipyIVKO1keelIBY
VtxXdIbBafjt1xfNAO3pcuWthVnC3l+FvuIsKkGVpB0YYgGRkwfaI3QQ72pM
BgQd24b5od0ABqcj+kkDe6ndNqibsoCMf+Sd0BDTt8P/+CmCrprszC8+UFk5
hf87b0gYYNc+wwQS0d6XB/VlHD5B2AKroou/WySTYRK4zoKLeCh5ZdMT4Y4I
Ue51RskED9vdK6n/evjzA24rrARzlrn5Ort2tkWv78fd1rjdyoP85JhMR0vY
nIjlomb+2r0wSjlj6BWeya1O1A6RFV+7gJZu474m3qw/pmslQ7RoRK5ABdEd
5g4fpptvYp4fD3QoMdgXwpU0c7RzuryGZguJG+0TOctKLllsohWxkP81FYt/
qE7ftkacSnxdlagz6ssFbDTptpcQ+WRw+cUyk9RvhSO335cqx6LrXEf5k/Qr
RIy1YuJolNw7w5uKzAzGF0VSNIA7MCPX7NI/oFNCXRfbzepJLEG6y+7uaD9M
UtQcrnwttmj+wPuVd5kJygjo4++8sIwbW3TlB5dRXq+bstmFRQpPsvfvhEX2
ArzrNf1Dgz1vHimskEhoHPRa0e38yvjP8VQJVHAXS5/+FXxvPSlRg3HwhOGm
3MditrqipjDoeJemzTzxFTeLnZsft4RJS3oCSRjSIq9zXenXA+uGmnDmvxB4
35SdmrBL9wAmv9S30cMXALr/KRmzWFKDgERIQcRvdY4RFQ7yKZfNzkIQ0Ew/
1rJ1Q0/VxO5ldRCuwJH/eVMmGWo46UaksLQ2qq5erIu67NWeFChiABHWZxWf
6ESYzO6lk8OTlLph/ErYcKVBRr+Nj2eH5VdUiEiaS80X99UfB8y4w9pMVWBM
C6XKsj41BB37qym5fYCxm7ij9mieQ7NoG7+Ow5HZwFmwdzu0w81W+nF1YxsM
RGwyjcD01VXx2K0ZFZx/ohHLt3MvB1B/HBri8WbEdypIn160ZfxYoOURUcCf
5AFngAXHW+g5vjQ4kCyCTlW9/ZT+5XoDRfdPoxgBa5XYID5i6kVvcATr8bxN
jog8097eioGoDvUn1PIEjZ3hK/dUTakuv45RG5PLMz1nM2anQpnURtum2n7s
i4evg8A+vsK9wE8sDpQaHJGZKwrMxxiEbC4Ay0fx5a4/tcATMgliTm7rGMMe
9tGBq8nzrsePTbTqAYixgzUPj8MBoeVGgyatzZn/Jo3Mfn3826mgr5BmfXg0
oobImCHGLJ/109aRaUZWgMOEdUur/m08M7drfsA4t/bztc7rQrnvgkncYGtQ
YwQavtN1cv5d/PPxgE4tkCCzEu3R02uQvMq3BDVLt8AguNF9al4KsOn+oIAN
/8vbbbk1fZrfNeJbTBiQlw/ABK+7Dk2WPcHLTnMDcm5pHego+CXKahfC+E7P
P6CTdOOYtHDGtqH0wCdr2B1LouzoX6GZd5jnmdZzpcunlY6y5y7a2ZQnmD7c
o45Dk5PlzR90KIOaiTAxM/dSIhAU+nLXwWKHT1W5kQeyZ4jixvOQYI+6+XJ2
DtnnSOhJU7SB/e5o7u17t93ZvqC+TENwqseLGlYNdN04bfipJ5AC0hko3Bdn
po8hCKt+kfnB5LohKx0kT13qW/+P7xjLB5WWdsWprpNR2+lX/WDOnBerAPot
qJWM1czaoV4vRNJTqpxWe2OUAE0MUUuyWaBN+mcgLMXb7kmu7JRfg0QJaBbk
vyt8QsC/HOKTrMx/abGdL/V9eK0vr+/hTXdMq5LKeSiK1LLpQQQM8F4OOVev
d0q+V6pzFyAKF0g+XKMEVYAtaaQ9gccRJ5drSM30Y4P30DSIprb6Y5EobLIH
wZNpMbljCH8McWZmaKwolnNBfiYHBX0jvsdwMfuc+yEppXfCCgs2WpMRWCrz
ykkKzttu9lMKaKHluVJPzr2fPX02YsXCrVkd50wT9CSYkIXNTL3w1FNGey5d
z7G9pRrbHDR8j3W1cwuVlrkyVlNLHLU/V0AA153Az2zjPsda4b6L6HFVNpfD
KrFrDSc0eamlUWsiw+VSpNLgFHTdhucNKerYrFF3CAd/N8MA0OpC7mn6jSO8
/O4+I1XFUQedpvNJUAtDbOe5TiIanWb2flIpukQK/Xu5w9QJCiLlwf8vnDHg
VrZGtj/6/VRXD0nmThP0ElqYXATpH3scVnAEaPTaUnyOWbBXcL8FLf5M/y5p
97PqXcmJ8iItL+EZ1+Ax6qe5wFwKFCEVIT6ziIskm4g2dZB0w9f1GrZ0PNG4
p+m49++ifl6c/EySzMfMCWiFk0g5/Ie8fmA8etrPbdI1xx/qXs80TOCOYBJC
TCqLmAVaxk9yLM7LXS5WXqjHXKdH8LS2HYU9MissOvokNOyGWW/mSUap5lEc
ZJTZf8nCxHFxoKsiT0tL7jTyNUf+76dsAX23+jObuHhuKNGS0SNpKMjWKRB1
SwcJL5qRcWvQMuyXsXb8ABPbaHfDzP2h7K1nHPq4jF0JiXqerS3IxYyJ5k9u
MhdGjAyytQ7bxsG+ccMZ/VntebCvdwrpUkC3m32u1sFR2vvPhtYkKKsmp9P8
Y48UK8t7DBoswHCiGT+9bX2BrahRv7jGxx+DO/NG9mVgL51j8Obe8wgtcq9i
tjxaLucFrfqo24p3cphpI3oaZDcqdgPWiEf11RpJbXJgKRFO5Sd1FlgJKP6d
CDFNLu2S8W5UL+4mCP4JEkJcd/7uBYmQM+CmoWyvPWRm7l9w3pfleThMJsae
EB0w8IQMYK8YR1NCBrfN/nhaSQRAzuBAn87Ru0JPBPGSysMRKoLrRtjksd8e
xHtLdHX3AVS71OPG0s8sYMqhpHX3uM5lbRZE0+24IHXn7z9CQDLNyj5NYwRq
UX35wqS9sOuAuNjn+vDnwlAjoQLqZS4ogAyJ6TWd+FhJssI5ztVTNQPD+Lij
rZiMwSrmiCYwWWjEQc/mcrhwZ2zlS2Tdzgy8bd74Mv3gx2lz/9s7m6F6BxrI
LOViBf3EQb1SsYP7SN+K8w+g6YuQRshfqvBCC6pUFLbcF9oBba85IqRkEE2v
XH+Voz+zFmb5hP0zTNcPWGUZQU46br/GhrarO7aps/KDQBF7pqPwZ9a80pwH
sfugKdhszM/MtQTNStX006BTR3a3+YYf/P6GpHiGhQuxVU0+FBt4jOey5BqG
+3QVoIGpsYL8nR7rSpU6UhveXEIIJCN9AjsxXGru7CwovUblp/s8apYa8aA4
94JJElDmY1f6pDghtKRWlAy2T/bzbygTGI2761+7qOcmKOvfF44evlykdCVJ
a9z7xYRNDJHUdThEnG6KVWAD9Q6VkuucJ1u6+nWw0dKvun63z64IbxHjTmyZ
HnTEk4ZGZCPbBYEnoB5me7Xnw1XOXNy2SOqZ5DlhRgsVZin1DIZ9KuZLtIWq
NXH6rV6m8mRVY/qK4C6nzBFa158JSTb6T4RPZdaveoNvPRvBE4q0W5YRybU4
CNYOlauwu5IbyGwN5KHt6QG6xs7dIutyD/1SQMGRB1z1ckegXHnL6Z+pwRvV
Wl0nkNOXr1PDtBOX8ZTDJwxFSfep+3CWiYFhNpzwJibRSVJrR5J6X6DMk0hk
k8hhlVm1JWh3WXGUh94C9swSZ+/QLMedRLS7tSVNDQsv8BaCI79L6VEoesPJ
6+UXoHC3P4qZX1ktK5eho0Rsu6eOpG8YEJidq1/QAB6MQzL0yfosGZY9Qlms
x2gRSQNPSWEbbygce6fPc2xD4CZXrbo6yjlzQCdsv/HKr4T+8Dx9wiC+5a5x
N+oLRTvp+rpHDdTy7MHrdDGFBqGWsmRGy7tWxFxTa6XlqW8B+9v+aqGmeNu7
IJ7YiSZn72bXSgmLPZvlBfGk2/28W+8kjQrd9VvfFNuK2SSM1hcK9950Vc7o
oDFJpuNJEMBNC5ljog6yM+RYmnPoMzQp6cEv8Bkhdc0n3cbxUxjT14UahoNP
Qj/E5EPCLjO0jcpZ7g9W+ncj1Uag/yZRw6u5sGJFtRs9Utd8ErAxgQOsFR4/
rm3b+COBK9H/+mqQKpy5WOgHX1Gs7XWn16qF1aWm2XG5FNG4BECy14DBw+Vr
xefz+EdQgfcgrotoUqENer209zX96iNwKubcpMkFeGx9xfrrL9LxmY/CghIP
qkaQznx0DnGe16e3nEfhLnNdRfFyy97RMKVImEFJSxB65rb4SvUdMsXjAEp3
WVcA7XUITFg+DHqEctcCuJclOi3qLPfQwLRAvTHI7ZEz5zHgjghhHX8DVtXk
irASn02A27DuzyCa6gK7xkLHdjtpbQXwn5+b8mCuLHsQx3+zE7CxnNNdNKYw
pwd2pu9TNNAR1/wkB/zlWThT6iVQUQZsAiNTi+ikr4OYSHssi3c1ewqhBkp2
DaJk2SjKR1izlSDy8rSf8OR1NwWGg2T/3KLjRCNdlpU22YgyCwilarz6zemY
e05a2n9pbyYIZqmupIX/prxwq9PueRsnUXuZ/Y0k5ILOVHdNRnLZxC8K1eYQ
dzbw5t2UWNKv9cm69pA1YPSO9tiWH7KyzHHynxkv3sEKfML8Tm6TXIpYOozy
HowVOgcxdeeWrhUjQlMKsDMe4ODGT8/Ksgtj9bYjJ40BF9DiMKz0VMLdF+/s
sdLk9M4yRz2fP2gR4zgYpNZyVXlLNsPbncyfAoROEn/oBT3KiHUBVxDmeKJE
iwfGbz+WV2Lq0e0wrQBSVC+4lZhp1ES5mmI8gV6qSFxJIdIeCoqy1z/Djqzx
4rDsGMIiEK60MJMSlD6ctWva9xeOt2B9kTtCoHT2M3EZkSkM5/Yb0vVyB7zL
Ry2xgJhQe8PFqBCN0V4iIMtDjWbc9/yHhrowTVqb29tg1bBw91lXKZpy0dxv
czUp3J5Zkt8MzdxCe1m91yQcmZMpMsV8mcaz8mQw8WufFPpRd9W/a6j9e+Kv
9CON7Q6JhQiUB1M1w8zKdDPFKNYiO85FMjStQgXaW1TsSZ7Y+KtMvZ7IpDDJ
03PBKHdiNZpStAqKBHuCLZ/Rjup+uSxZccMtUIClsWcJHJzTX6gHGclLqyJC
HatEowXHWw3TvEE525LiY66Y67Lc/Po7jLIqkO6I4DiRyKVOXpk7LICSNon6
saaMqo5Aw9PHWdFTrNwIPLh9FMTb2MIPTHhO9t3eZQQhAUiuW+A6JGOzwrhE
g/f5eauCdjed9VdqIYX79Hpk+onRnk/0AGbiNvJlnxfv12FuonpBQye0J5tR
gboo5AtVlY7hJnPrX0q0JqzSb0VSOWaOJqt2qxc9MET+Gm73Cgoj+Hd7DLHT
BvvocVEMTT6ubrSsEjPUeUMw54+qIqZYABc5SxKOkMXUtURAqhZZ0ARaEmYb
YuG9YjiMn8TSJzAufZD3a24g1UqseyqvZykrjezQc+vZAm0EUJvLGbXXg4+z
4KiKs/2KdRIqzQi1t/jOfYQu72+dCtqYr2Yk/ZdEDQ+8Pn7USFschehizC7N
cukJCXTF9L3cKetclHut02/3/HKEriEX2dbi33odh5hkyd36Ehor7sUt/S2a
XVtZTP+ad7fnSs9DJlvIxkyIMmr+LfbOMlRpMDasqvXUpr5v3w67gL/L6ukG
RSb+enr+Ey3991DCuYdNOYxB3hVCK0Plq+Ygel86FFtmyhH4EDVwVle6lsUB
yEqq3nM9Xsi9ANRllvtbPGtjf2mH1IGaY8yk1PKtPMJ0AtAlUt9okGIRupdX
FJVsAwpd9ziiYZ1gy6/1fkLy+r+zIAgE7fwisMST9XAvA5nwP0nWCZaD52Kv
YCuKt8ueP9kTdFRRJIzceHfKKijQdXix7DD+45VDSNtHytE1nB+xkKVSkvkJ
pOE3jLgwkG4YLuHCwc+duIWHwgVLvvS8eyb8ZAmCYt8OJJFa2nw/VKmRmjvV
HiEGlU59NIP0FXqNMwcKibZxwFBFlXOUSkwKK7eZkAYxzwy3VjScI0VLmWKQ
qIAMMktyxW6UfLZdSiiwS+ZNYvgDPCFObXKdanH9rxRyEDPv5mckUbA2mQ98
9edgnOCKKEbIxsvABseetj2gzjL9oMWo8Ta4VWRqWXbHMgA/TWec7AFwR6uA
uK96FoIJbvxdiFPTL68oQBKTAbdihDD2laapaWthQdJSYotQ7yfKbjmLu7R+
OOvGd/GwFW0HqBXr0GXnMoZz+blo8fJlDCvLL9J18f6DogasNg6jWVgUZGPB
sJeyFnk/cNTsm2D0G+zAozsv9u35aRnyBRS4J0dJ9+qblrXxy2qri0vYimrk
69+kHn0EpcblBEKKQQxEdlfzBJeU1z2H5+L6Vj0A01LiFkKUnqGYvezWUidY
cMOIVaRHqLsXFCh+SVB9L9I9MGgYF2YwPiqOgvD5iz/Jq7T/T4BmybwrcH3B
wv086GY0kxH7V/RYt9ETlfHmZcKbe4HQ7IVYbVwgv4QiNrfiwx4P2Eurvv+m
TdAiduADYtc86G+1yd8PAfTWDXguJ6f2FWWkHXTaBw068nQKxm+lMsYsOWK9
JNRB4elQBAftd+A3oyE/GSaJmMhzW15Zy0BdFsghjQ+K7fKqmitHe3+ATkub
P2bHXvqt4HgB4caODO72Hh7/v64w2pxWcpyfzsPd5MasNXceW1HFvr1pm2K6
y7pyxOMfCGeHUA+tQY/45qdAvriJhMywKRDKmyLPs0kV+wz9c4mE9VU+ZqKL
zLRVub2B5s0WqO10Tg2JN3agZEEAp3SEbt7DlTy7YJsA/kr7+dsJ9NhRRQti
k0WtPVumusFnjguLIkWPdixRBRHuVV8rGkAHAdsdGj9uvFi5VNNSmxIsU/7i
1TF6lf54e+qUreGjRmiOiFr09O1zyQMFVH8/rJZ6GJ8eyhx4Gb4DckB3LFwn
QmvOTK/L+kMJqgrlpcJTOtCKmvgX7wB3sNoT4TRSw+eeg1a7woRN0slgL0LR
Hhm7Xvr4EFIHFOg4dGF88sqV0V+xyXk3052SQeDOci2IC/DaagorDDyDZ4eK
/22BuqIoidzwrYwIFtoNcNgJJjvZ1KNj71V0bw7MJXEYtePvFySy1cle8uc6
+kFlWQtBFeSezmKZufIQKasF+zNQlg5tYKKDaZMY+B/scNA1Qy0gR9eNP6NE
PQLoacjtQa7NnC6adCzOHa3Lw/03v2tSm65zkOTyjWedSvEP2540X1D7KXHo
gefZD5HWgqQu2tJ1GQTJLM5URGKCtgF4pap7ZpBirobFZO9kcbhu9QR6YnEz
ORfG/rI7aM77ZI+gcpcyxu7wnzgpPh59rI69APLrWC2ZOgkrw4BPwQUU6Xml
ST7uckqboUmRm0MfBP0BfTPWhFsqwBxm2jemY/uarzy6QykBr2ecf2kAONgf
IrQPtfrbQcQwhTvxkHRMxJcCJ5J2ELfXgMNAx0D8LgKKgIjn2ObcJKD1+BEE
uY/Ke9mzOYmpTDrMczLwtM+QClulrIAyRzZ3mv7qnZOemrN/T6pMnYPMvbLo
s1YbwYROfnQ86CUROKbAYDiU0BaThisecn+IG3OLyWjEq9Yxez0NUCBIsni0
NrRvvppnA4R9Hi1L6ip3JIVGkTwVRanS2AHAiEoBsgyUBouzHCdXWEA2Hp/K
3bvMYddZY3oe6QBk5C9zoQJZLoX1au5M0LPYw/x1Se5MpTri0M+/NojI9idq
dHcDCLbQNideljmOQ9LAiQqfKeAtyWu4Id35h9P5cAtnJtd1SlrYTpoLB6Co
BP8v2fMg9w9igBwngKsJ23VLE5awHf8+Wzu/8sbmKksBR1o05yH2YSMmNtAv
clFCdHfsWF7scWEi+7Z3yAo5vYHhMhMDpQP+af6NWXfvstHCOlIpcdIlhHsm
Oip72KuvNDojc/5Q/sHdeCG57B3HKlZJD0YY+kjS46oDehx3H8fylQfYtFEi
dOr3Jw+vIz7yOnppVJxPC+2elhrR4/Lp1vKna91mfk0BydmX8XpTo6DrQogh
J9nEJ2DeWMcM04C/AHarmovlJ9PUe51M166n8EBBDAUwS0brcgR+HsLRHbWq
yi1k9Vo1bFhBXATSWKqsS5ML4ykrr7HKLE/kugNGQx6AXBqiAOqPPEpE8nz2
FJs2UXYRxYC01G5ka6Wi4k1JkfzZpTdRc+YJBOQ9ZzRZcXSxHwK5yxllaPyt
/gacChthCQwtxlEl1rDeQE7B0ZnUVTsZ+/XazmmdhNrrFCDMn8pWKahXLK8C
L+1XuGK9xWr+71f0vO7DTjWrwWTkRRZwB/AlJPtsYirYf6x8TjY4l4lpjlHt
kj/N9c2KCRtwrrMcUlmdtn5xMfr9WSDanU/dwj1kxA+gEFKph6i52namJX7z
Qoy7WZy/7HhQe1k/NYYwug6XdG4vePTEAm/5cSyFWc9vlt888E9K8HiPQldV
SjmwxoD9wkIT5v3LT/HsSheaVyrE18UhtA0u+xqJOMP9jvShJGxMoLljQMhC
Kx3F8zbTuG/ukzSuWNjxz6cumYo0rrd3H8Xb8Gks/VENP3fAcBlSTyjPAmy7
2+2+LQoZdn1TvtNuxGt+n1c+uPfutz77ZLIMhlh+RTIi36DRRudnz2lq2BMz
fVYe2zE4NPMbgXrUjKJv6TPjn50DmB8npKJ27fzZGCUsJoacDpGhmFPnxKl7
2HjjL3fgsJQ5cln7zVbmGe3N5+VKrWaB4dhaLfq1hMy2p43fNySB7XiC4OWV
up9w5DizutXfMan9yUpYE2DSwsWdrsikDvO0+piGPLqemV9w25elA7cqHTC/
NHPJ8/VCi5QzMQ4X9dXykinVdElCQdndXQSuN64Itz+CzCX5dZyVYRr8oNJ7
s1WTkpuCJwV9vJLcro09lgc8yNXzl+xZhZ+Kvy5SbBRGvvOynElmTu1Dq2QV
2zdnhR4pk8+j2pDvZOXD9y3wc0RqloWQVrw24lkbf29+MLBw2vnnY1Eygz56
Z7iO/3yu23gycfTY8gQp/puzLHmmOtrGB0hPRFqHaKwr4890U/T8I6hSKc+h
DyDsvdj2fT0sjjOfNjX+j/7Zd1NmytO1/qrlcDHWOAR2BqwbQsl+yQGwfCON
uSVQKS7wh+n6kxSQJQgC+AvciIMEKkW2IgzVY/3bsLB4wvkEf6WLKgUc8oWw
bbYS569VvkZ4c5aODE4cNM+mivP645FgTcvFDRlckoo39zWMfKLMvATuL4lg
ap2fxc9eNo/+cNbZ6OEJd+RJy0C7+SqL1rME71XUc2fPu8qb/6XjzG8Vcy1T
b3vBboXrzo+jHzVv2AunbfqkJF0tLgvIe/QAkqg7aJqEkhGayf6vCLLblTMw
0asjXci59c3Oower5ZfsXxp88U0S3+GH0GD25K8uy3VC9CLRf6Qo2v4e9qv/
3aCh2Hp9UIiAtze9XmKhR9a9SagowxxfmjXktnJ3srdyBPGtyHc+GgtK6kj5
ZxSp38jnxm8kHMlN0Sby47Ul4EBqC8fY3dnWn8uYBbgdin90j4NYD847hHfi
LGqmv9waKJaGQjNA+oXpWw1PObAowDe3xFW19wr3hvlHHoof0hOJsQQ6iMPu
uTUtcsvfcjXAr1CRY2v0R8P1nUKx5Qic2cfF2CYLhrwsGIXKSPSg16hsgD2V
q6YJ71Rx66tGohS+LVIJZ6UXWzYQyP40WjbmQkaG9/rZMXI5o5poTfJEafum
OSTmjEffYOWW2nRqt1z9KcsloGCtVjTdGB4KoD45p2AHJ77WyJXBj6FQ1AqZ
DSQ6kTJUsohWRsRYKhOmm+HllFAcaQFtQoLVs78IV44n6ZEm+YP30YNpNDOk
s8VlmrZeKyoXAmQF6dbYC2YuMwa+qZ+y95RWoXPP/4xhPeLs+VVbJaLzNO7o
mjF9VZETzrzXrdCS3aYVFSyUz2fDF2Uql0HU/MKVS4jWhZl46y3Yqv2azkmi
siMr885GJZ3K8tozX1zPQH/iCIMAcBW0Lum5Igz6kCjWcXrkXtXBi0gJSsqd
kQ7xZm8UXDu0sudlzchnQ1Y0YcAvzTURU+6kZAuv6JbVxzo2XaqJgw/jifa+
tz9IB4exAtiIrR/aB0TSOj3yGYmOuOJToX+zzl/VxasKMZuzhKuXP8zeQQcW
4XE/Rc59Rf1gNlhqs8ksY77utVSwAOni8tglrMfDO3wOnw1KERzmBznqo5r8
UepcWJnj8FYYbi8AS/Fz7nA/I/qEz7ByXhV67nVP59SYdUdW2f+JkUuriRya
7oue9QvPKivr2DP/5QUsrCzvr7nXjP0k/eTAnSNNh+knY7KAWppTeBWgKXQc
zTP5t0BHjdU22JM7W1isFdZnQ1RWBcNs+gmulnqXz1E+0/FCSWPXyBnjn5An
yYjWJhaTw1f59fyWWHYDn5c2rW4vusjEpZdEyiOThoNUQxWJVw/StFgGm/qX
aOYUzgNiza82dEURfrx3FKcXCLLfo6h6YWpx3MIQnJ3PJ4EiPM+8kVfKIYfu
ECyoPgqXEg9ugp6LXcRP/aOXRCAqN4NgWeOQTPt6lmxnPOmzOKEoNZ+pjzVz
/BFv4dxMIZrPJravJdREDx1X1lxUgS/uIhjljRAxrAAf+CxUe+Z4ZBbM/+MO
EV8uTcdRw3iu3jkf+XA94rRoTdQes197Z6VcR2sla53V3JlQ9SpnZ/0o129k
2GynynlaP2ToytacwnxpQsDQgNM3lIT0bGw0xilXxSyBnezjHsdzNX6uXjLA
tDvl4eqLK22kJyCGBbMZUH5cGXxtogXvV//F0JxYtStH0HjUFOntqgXwyHWG
hCyggEzA9vzj50AQDb2g0kRFxhlmchvbeSJ2hd76Ot7CoGjymjksZwSDFgO0
Z31BP5dx+jyK8YLSQLFuOVPc9E+E7oAbNNvWtPbk0T6AewWhzPI+JGxdCwz2
ZBM2YLi8v6YX4ppAQUxuLV3lc5dSrTQroFB3S+rO6nrphJHHuvCFdR/Jmyye
vlHd+9hjSTr5U0iCeJRETofGKlVm3MAEg15i5I1WR2mBcahG01FXQGmLv2Zr
umV2aA8CP5iTk+zFaeio302LbhID7y3/uqhTXEbNhYEYgb/c/GXjCWJsgY9u
hAy4mXLwwSpLqVcYPz4o5N8+l4uaNq00N3FaWh7EHW5pXecGsC+Lo7zWTVdg
LBYid5NWDS1dTE9DBnWir2DzAX242XwTDFOXn2t11ncnj4IYck99u/PRd4Ms
ybs6/PZSV3BJUZK3vntZb1xkOdlsJg+csNGOvC+CUim2rrYF8laeX+2JVHwm
tFGqdWBGgYBotrD/KcVhH2PckyUbQVhonroo27XUv/TxHTL652pWRC+qOYbD
r7mpzzkcD7NlSmripj1hlz2k8MgdNE1FFj/VadNBPmmdA409z++07Vudq15b
7YhF/3675hZDfAyexxbhVICHAAYsIzQchzTXRjOShcXJF6aaQIX+4DNr7xZP
kCpFr1NIlTqzrc1ZhcgaUEOURPeTZ4xgH9ID2TzEvq/yNsejJhTiNpKxLJfp
ZuVn4wKFfiJmDSniL5P7nJqOASTqrd28H4qT6H5vO4ejiC8H7ABeQreVabOg
tITZTR9j5zH7ObL9q81wpgXS3hNAC9X2O3aga3FWfllRoKiOWwHCOJAiX91o
hy4Wdt446la4p3wYAUHRUqgKHdrK1K/UVcUw28jZkmverSnkVY/gTj/CHx48
RW32b0LyWfHb73WYqrcU/XjEI4cfySYTzJSIUIU3VixTP6bOAPCG4+4nKEke
mqPZM6rc6UDryLCItJm07ISRcEfyuRBwm4czjF26QyRqcz7bcG9vpUM+wIai
2dGlVgJy+4bzf/RpWDtkr52apumaD7OsuMaEu9um8oyehiT7zouJ65L/mhVE
pRYv02tf3o3lBmm4oXzotDAhQ6Wj+PQ03iLbFFcLIOcyajo+Hivx0jwDd9a8
ELKM4WDEs6uKZNeSnibQPClCKB0+U6dfEKJaH/lhYTUvXx0r/ndQ46Ag2pOl
EynK7OcTjilP3PUwGXigXsAWjYVVJ7qvS2ON71jPYMs/PbgmZgiFyM0T+Lkf
G4ja9MlezJzqAVHXYawqV5jcCVknZ1XPeVEr1BINt3JNMl4Cep6b+gSBBes3
9EPJwLNQuNjweHmy/n3k4ghrnND6Pt/elUlI0WCutI/nSadD9ItyMp0SJyRa
0XFbMEZjFigsG+mbDmG4gVQSlFTG8Dm9FccVTeQ2FkjAZFmm5Jsi25+7aIVw
L4ZGfLmBrsf75swMRdRpQ6kzy4aMBrxIcIrqqd+8QPhFs/2zm6q02wjmLdRi
d4v4cZQpCOPZhxa/jHmhbLkKfFTHgR8NDjY2YX14C4iKVCEYvCRFPbAlHtdL
xYmeFcUKwgJzEDEv3nVHA72uMrOIJfm4DIM2JvbIRG+iWXIF9T9cKm5GByZ+
3uH799KVd6W275rdizwZToabicicVAJq7q+IWmvyTvyhjz8Vx1uFcaZQRLjF
H/hNDkKmwK+9MDJww2nHIUhgpg72T4PlFtDuyFGTQWVXAGvLf1zx0DXCwnI4
VddYTY/eKUQtV6y113c2HU/y1fDRyap21rNouRJFiv3TXWpIyCBe0U2YLByl
vzqNI7LjYckbRcp9bBX/xriwAHmTPKi9+s3j4W/c6bM8PnO/51j3VkqVIrYC
Ftca9m3fjCmwrc9nz6rzCDDhmq8mQmGXo6wTeJ65IgrZcZDCxr3q9xR4WoDT
0feRTo0PzHbjOEv4EqYNHXTHm4JAmQxJF7idIaXhZ0y5Y33o39Q7H1k19tO8
mzu0Nehta4VMTyw3prKZ80RpJgaCM50eg4LmeB6KjCfvK+hBDZ8DbO5EaIZC
P7HSBeMTMDGV4/WB3QnJxjf3yOKI5FW+I1WxIAouWuaSBY2/24PzcoWuE0FF
rcK9SUG2agx37KLyWgJ4NTwHI/Q5oGcBPnhljVwK/BcMQTmK9jWXn442ijXR
WdShAPcB276MDEjYDhxYqgMpqkItLm5viYcWsRCa/j3A9wyHjslpkmFXUF1O
EOKXGOXhSqaocySQJPO3JYGlbQ/MDgQFlMIIj19noWjR8p/LwXlJQzSOSoz7
bOn0EyenTbXLSIi8lGgZes+ss4Wj7LJqfAyUNK5344MnVaTwfY9jFHwNpc4r
fokg4WoOiKekgcWuRmKZWJnZtuiJvd2H17NVzFAItXXXNkdb2wRDiX76BVlA
0BgjXD0G9v80t0M7Zuw+T8rvvH1DqUDEpYPuA3YGfj0qn9SuSZbZ4cxG5+Cm
l8P8Jf9555WhAt7ntUjHtVuJMYJPaigRA/tcb1gobhO+ELZ4JcgprjbtsDah
/uTXApWX7+Sq09trH1xWu1xJyaKO6C+fq95nQYeazCOPDWK8HSuDoOejHuVY
cC2cRnTz9nD37LAuqxx8AVbEz3RP2ODaAsvAHc1xB/Giihiq0JrJRRlkKGwn
6M2dwlvI0e8jK7AQ3sst/BCe9nZxoML8btyXJLYS8r62fZ3O2B88BGPKyg/1
9JiuL+WwpGpNzS+gN80t4w4zPxeDSy38Lfw74moO4VmnStV5VSFWnuHqnKlJ
LfnX6d6kF3cfX/AVZdoGNHi8bDDXQJMRrEWtDWUkOlRhbCR/LC3L4Ff03JlC
99ue0a/gUqBAFDhTdHAsKEM3lezUThCskR9DyxfOGgAuTCyYYwTyq1jl+npR
kgoH4v3G6e7kDezeBr9A2Ywqm9orMbdcviHyOat2hCuZu4jRwuTE10EgcDv1
o/hgd7Ea5R5e+Vf6oPVWPYnsImn2xJEJM0hdV7mEcxJZFk1sbYOrhRGE7Xz0
tC46dTa3jBQ/2NNcXtmhftgg9MHMd9aXHDBThQWwOerqACYAI48X3uHVeOx1
FY84wLCdudoDvv86ZQOMlqc6gvDPAesN2AaqnWSXRDQdGb6sFxZggiyV3i6z
k4rri2BnailoFYqzmXM9xO6IuXAY+TpRNyjZQm5XIfE8Ipxb8GjCePPlb5Qc
0X23G5+j2oDZBlUXmDYX9CrCweiGkvcXUIT3yHaMB0kXPyWuu2HlJ2SGW8Ho
tkjtkmFuf2xXCMNRk2RyJZK+j9W0dMukMJW0XbAVq89g7t0dh5tJ53vbawY+
c1sW47bD0eqHg7IL4N9QzKe61iOntI19e1DqHCopb0p0QRd+y26E4NGMZJMc
wUJYdwSGTqx2pTF2g9+AecXRXNMWHeEkFWEi6htTkeZDGn7rgV4r1NgFqK9G
H1JS/2kf4Vp/ZvS3GYzyBQCf+r+LGfneHedzf2HBgez+icZ7B3B3S1/UMCn8
0d0bHKixJX7U6v8GJK2rYQXk/r3+111u3NG9Y9kGv7QIQA3eThAEr9V0MUzh
eg6L9X+XxRdqhZhzfr48jJEDZA9XDVKB4R1gSRGoFdQPk0JBy1d4k0pk+wcQ
qgJbpyULLeMVuLRu6PvWSEEgDfJYM81AuYM4qQND+5OC3kQONETvwcKWbxF+
S6cY6ocA//SZB5n/3ibeOmoAWf/sFhTNqY3AEtgQn8IVxjnl2WjVFu6dHYMa
TDkXl8D6C7mJUW3nWDKumyJNDvazAu9i+Mzbps98VXbVypvBTuZYYJBQ/nJC
TbjFJZsNFRM3ZYi09Ecxyl1DXZuozmUaKY9kosYEe+qJHmMesEsirXZIlZIe
UlSkCsdt4K+4+TGpIGS4DNwsEdLTWHScH1r/wYhRU6C59EFxLEn/tUlBJwO0
Sqm+gZTwpjUW46LITwUhNlWcUy6ziXzuAjPdHcvAWbCTPjq42RTV1YJLnNUr
pnLKMVp31BbP1CbJi24CZfsxM27eXTHl+m0Sfzqp3T5Zwhmse0ZJyP/xigEP
q4vhS0nUV92x7hy/tUx4vr2aTFWwN/tLH79NxLjb0EEGgBDOlnVsQuZo1eIE
fev5FRDZwS6VbTT36SuEZpmn+tw1XrFCSd4PI1f2683xu2u2QDYgRYe0ZadC
1iLlg+YMFayamUa3Sr7rBsJe3ZDTOdUIHXQI9d+mCilOlCLzHSx/X32Yiy/k
DXHMD//h+2gD/pIBG3Yk0yCexHpQBeSFlMpp+uV/qSn/ImOHYmgZBdUBf598
DA9VLhgWBp5vHFtrqzrFcfxoeKAikRxINybkG3p7pxZaN5NYJzDmuLo/o3aF
ItHuEdCon0aBCkYQC39DBg4vRe5AtDUYuWD4FrHWdLe+MEVs197dHEtp6d4X
sT/m1pPJRq+ezqHyQyoqcMKUpQKgs4qKayVfr/EHxHXYrcUZRkWAhxI/xQqg
PEJJHWXniAT9qdho37bFd0r1UDJHf5kT5F7hDEKcxMtSd9RFFHo6tAiRCBzS
0qsVN39tahFY64gSXno/tSInJuL0WmKEWoQAbSqQo9lcsyrBAWmvsjYlXqFy
1IjdjLwDdqblm+hivgo5cVGk8Ax3RZ1qxrHqCUPB0tlZZgJT4C28z9SZOjw6
CJ+mnsNYxKzOlvNzLNe1nV30B1DQQQjNBljGiUsOBppLkDDpGULP7QC/LMK3
zk4pg/0rDU+WMaUsdXxUSdiMcxKwUa2MMSkRTt7RTgO+xfzmif+0SH1MCGMV
4YHJDcMFxoZARcdqho1cQNNciKydb4ro6Q5INzffO6ga6po/hKo1KkI/dxG/
wuhQu5vMNQKxH1zr9knkxhvL1hn7/UCY6bkYgegeHrkGoeCkpgsR49/Niiu3
eQKjrSdHmeXXWru4yz9pVYYDj3SBNVKiN0xJszvMqU/2fVGY1i3ij+vEfa9p
WDhWeI77Bcco7m+sIzozdMakDBISZEejcWsUU54zZUSBJ6KFXQo5D0sxzoPH
o9WPEIcPifP2V6xbWBpzHVqYO5UpJ0tnhWRKT2x6MAozpA+f9WaVIdRZ46vD
Zw3OfjgLaYc3Z1K5t/MgaivfNhgNrfktmn+leOLCCwM55OJ7s7Tp195NkzKI
vL1ctYmx1ZBjNT+JfuXblQETNDw1QoAOAHgfXa3CuRyXUsghYqHCXUIyVxMO
/v/OFj5xxRT/VUufP4goHMPiTenCVzsbFUKUZkOWOAYESbDvOiJMCQ2Tw2hf
o2rKrugcDKdtlYm69AaJFBQ0Io7zrw8irK/Y66jPliPv7t8unRKdYNtoL+EL
oLMYg3VyiJX18GqyxhQEBKvGfsbqJbO6qbc1KhPAzKzhrlkhMISsPlkUJXsD
NxfKzgzXWANyWNrHndUKITiYZly1XZ2CuqXn/CZI1RmZbPo7W/s41uHhrGXY
Vr/QG/qYE4xHAV8E2LTkH6L8deaBavkjJ1auPzqsBM4sriEbubnxMPIA/xxM
4J1yM0+TTwSJt/lXvdotK0Rz4d5TzRzzk9mICCnLBH4eAjRCoKJmL0t+YrPx
OPOyE+MZLw8S+Z+gXmPPvX1nnoj8TiLyHV8gVFrDNBQhyJNSqMbk8dtzy779
l+LtnqE6nNECw1mme6OV8VbvKB4FcQ1YBjZs8yqRoQYIFlAtALw10iUiVAxE
Sou9bMztg0cyUzEXbkNnaM/XuNlHPwfvZP594GKZ9+NOy7YgBeNCcsi28ykr
8kkQtTPw9v1s+Biw+b3B6zwz5C0gARsurkhdstdUR3DB2bu43n3v3V/zjmKa
3TXFB6JAtfVKh8CODDgY+Z5RhovEoX9JK1cGMbVjx+re7QponAx/oRdOjNDI
n4bSyRlZb5YJG6cVJRI2ZnKl2P1puLpT5+ZTbBjSTuch/jKUgqnKH9A5hDsG
3J2vPWwxVEAzcXUjc1pdjZCUYDVDvFL+C/ptPuDxpdDk7tBdCVY2TbITPv6p
oyWhMEYPMS5MaEL+6TXNLlgXlPO8wcZvOTrqa+NTb5+VuMTEhuGPlFLAw+2N
Fq4miGWBoMianfsAG/VWMNZGs7SfxVlk6wg5JHgtXwLUMmBZJHTz0GdBfH8q
e+oFbfeet5A7DtAqLgMk//HTVbJsQ668CDAXP/uDZN/tkcCAndBY5hrsWZ6L
+OysJIMo8Zvm082E2e7sCm1d53OIDlScXW7he6Bp+yIMxB+Aru8lji/ODXm2
oGkGQXNbK3VS2m54zYMf3ZNySvtxdES3iooMqIaSnyy8NXH/QyFhZgD9vTfr
NWTW0qV4HQJnD/zr+ntEJ4D6i4VXZMCU0akP1e+IFBgsYSkKKJEyw+I767G1
HPg9pvJIIAzVAA2g2ISoSRi08B6UT2gMV62UUoUyR2vvv5xnnDRFXywj8IL6
agIuDfwdZX8lcWI5FA+aS/OS3K/g2OIxIOaTyxaJp+wwf2PHvtT9cbH+bNbl
KU+Q+vBcdVs5xxt5kQIepia8JDUXk82J4nA1/qKgmdFhfFLpks5aoWDCbshq
2amUMDqppLhP9g355adojReX3xb3vKqX8AMZZfnnRQjCvVDPeBzu0cuSXlF5
tcN4HKRQa5s/7DgSUvtNf/GDSPqYG0UH73ay63Mf3T8CmMtqr/Cqmpk38A4G
0R4+wZccsSNZdzuLQyfqanL49GOWcjyiHtGkbq+OTwedj+wlqxYg7fQ5rMRb
7J2Ywy4qTE8OP7zXatJSB0jDvio7HCbsuQxStCXgUUVLPkqjaBwadAQvO+S4
MihOKamJkZCqDB38fxgz1mAHqNHKA2Mfi5CjUcmE34tAjtoTwXA6BGUET7f5
63dmpGP7A4Mljp610oJpJVTXD3KmO0s/tYkQW1XVLP43W4tPdYr5NuW9ITah
WAM0FVHwOTLCLE4f8BjmcJ5qqip/PXaKRW3mWMDFZXodj9L6dUb4iw8rR2gW
Mv6oOMocRwMe108wViw/qzBFX5Nm5fBVRhKioSHwqw9lM4vMRTlzJczZWT+l
/68ecYEw8NbwxhO72ojGqOzEfGB3gjMDgFcNE0Ea/5jGgzD/vAU5ngSgX7wo
EmVtwUY3QIwqBzbcidVjnxY7gD1NpkPE1dJ70tjMz2yk9w2MJM9fKXT40xL7
aX5US94aNkGZ/iFMqy737d933O3idrroQuPJlXUs/nP4dqav/JWsNSmnVJRe
Hrc4z6nApE6a5U/dBSoKJmVuojEsOiPVnKiNA3QPn50cgKV5XGU/cDCs0xzY
D5v5AX3/7iixIl6Ixq5ADmUtjX34Er3Pu/m1jfVtMPARI4qkeUHooXxgHALc
WtmQBy46K5qkIusLKXuze63pLh1Nwb/oIxhTjvpEhSkR+DClWVBkgRjbXzXM
kLpJmNJ1YhwvGI2gvcmnYpQJbPYMbBL7/FvendicyRDOZzrYH0p8XfkPdwye
WIjh7qFt4caDnQyWh5mliE53YMIlqLowSztfod76r88Zu4fv5SY/B/jiGGJK
th1fuc1zqjwF6A9uIhafmHxZ5jqLLijkFmdVTKihi1ez5J9XGQ5myAcym0Jp
PVtPLW86XfNJLSLBr6L//RxLqjZb7CU3htKoUTu/zsxtMqVLB3455Q8WaIGu
pqB50IRUlJdHbzzojUqBPczvU6iAitQR17zNOSRif8KS6egyOb0gRUIHeBVQ
6OgY22qHSgaVyrQ0aIClg1V+2l/Hth82FQhi2DYAv4K0aa8310RmXXsbzQP5
oOudTJ1n4pduQqb7YoTlwRSobkL1/GRKq44y3T39LvFhpcZ4dvIYc9Dk8wi+
dPgAYrpEb8KG3kRIwrE1Qlw7dSDBn6pkmEoDJiRsqZZSFIVvkR8pF17KNUgJ
0l+rnj7JV68OTcCFI5WO1E8sqxaKx7oTYljZRSw7eLLWw9ihhLdiQIaQi2Kt
clhQOorie79XlJBdw4r5M2csShElJFtaC07Ek4u+KHB4e/B7FnrikcrKb++K
ncsgeo1godSkZiCsgurdUjvMlRGgkNZ5lbamNBxcUwXWUa2uZ3SvmB+BBNFx
7WJkXmkcFcMcTxdXTCgwlsZ4/FL0y51v8M0nw4TrUuJj3S2M66WG1NEFF1JS
WjydiEmZlZviZJRfL0RuVeMzV17Jsf05daYGqbiT49vu/ecFR3vhjl54RyZd
LwnngOO8ViAVJI/8Q15mls5jZ6O0+YZL314+hTcsEn/cBlGJV/peDbHIOifz
of44rBRCXGpD7adI5ysZiM1y1YYTrUDibxfb6aZ2g51k/2bHaqHGi1S9MVH9
YOGzwIdXm/EfYG1xeI/J4wskUkrPY3BWkPj9/vsn5lRQ2Rf49MyAyLSKGouu
Kpgki9D38/WB0oiSMVlHS477dcORrH5p3W7B0X5K5EJwpU3c+a1X5EzKdjOi
07Dct0hZuffx1sfaln3G3Whju92DZwsox+2dLAHHA6lhhQ1oP683CtBfzKPu
RLd2Orz7Mzti4R1OsmCsTvH245EpCQJBIChY+yDI9GNtQs8+6tH2GdUyKPzC
DBdNNoGUrtismo/WPXNPOKsa8GzxjtG762QTAp7zQmKbwYT3tgVLyzQNgk3u
vmsV+RbjrqxQIi+/hFp06fbvOkuOANEX/yb5HeAyp8XdkPuAtPGlr1F/L47B
/dZRXhBbn/J8680ONxj1V2gA6ukZtJRG+c0DvNhFEEwp9+rnZjrbifhIyr5V
j3QY7q8tcF9/NS0kYbln46anUm65UX9DN0GkX30rHrMvTVigyFGpXDNqISWr
6jQNxeCNAZ+bI2Qo7HU3XdrPCgTdPtDQ8sEcr/Bus6Ngr3TdSACdo17xo5qn
Dfnc8LOwYJtnpRFUbsVP+gtVQHlpFVqyogMIuWN9xXRZysxA1hz5k7d6e2/J
wd2MLlPl4usb78AkbarzVABQLtmWObzAtEJg9X15B+EdQsxxxxPu9Cr50F+N
sTPgbolQ74Acm9eLKdcWTYJh5U7Fogg1hLsAf2XmW91JHhG/DhnAnGzFtTd6
OD0jwATLGgG0j48dHwBm8R1gnxFOsIS3USIWHnpJOn8dNDeMff4onmWpnOsS
BkU9+mOVJq0T+gmt0TODyz3lqthqc7j/TSLZVbjmZf0UEePoRSWn5YeiFdMU
98AdHpwr3pebNjBFQNPb9j2xF2qNq1eagzq0xBpCrhmJ6PTYKh5upNXZgBWJ
puPUjw5f+zE6W63msHpTEBen7mUcjHh0SQos/jHJa2HvrRVavyJ/zKnwL7zC
VgXLa8Nwi2uhPohDNiB9kyMnkr14vVExw3GyhpRGTNO6PxDZfdltODtryf9z
dPB+uKrQbhQ1bnZXnaJRV/fZ/S88n94bQdtYm0go4V2yzWhL0N03WPGD8cAY
ZrRxSMCHJvUPBxO6nPq7cqeTZUI9vrqo/CFnuQXqnvyG8X+lNkQ1SPszYPmN
HiXAy9vZBufDY0G+QCRE7wXdskbQwh1L0ccDS9loNT39QFNhHZhkvm9A36Sf
mm6bGP7cmaUbvQYtkHt0LAUeIlPLKA80lsL08PtbRJQjlrRYdsvgOqyERqBa
8kouWDUvFOCITycYxQnB9EhYWsfCVH2yvGL/y3o7IB6F9+2mw7R1mRhBEOFH
9n/iPga7M3rjcp/eP2BXZnJdUQMnWkLgXz52wdtWxxOH9iD3uIQ32aX8QaVB
6WOC/sx290jLltvbdJgA2C4HGYwmeh8eSMAJLtWe5uuF8sbq2tly7KtKCcfl
kSVj0oT0sVzSm+nsQ/PUf6c3owC1m9nlTjuEYSTI2Xp1Nd9DuV9n7V7bIuJt
81HjJVsPkQJV//2P8lIWMV2PNbfFt4Skagjl0DwbptX5GdAH0yOgFyudomLQ
vMRxI8Ar7vLqs5ae1LEEIH4k/Ky+DjH66LTedt8VDISuDUC0gfY2YuoaGK49
mdcdo2X/6dawGvWkzPHwlv7+woePDuGqz+aaSmCpvoyeF67gdJ2XvFYgR18k
yI7/VUpUdcnL4k6WY7vDI0UlvHtSSSknsx+30vngXJW7KdSfWvkDDpfEX7oR
h2mdaJBo74SKi5sAPQncJEDyTImXKnXUEwu5y+nv4smLNRcDzVMC62P/S1Vr
TJTZUcCIhTNWXbI8L3BnR3SdANvmeugAm5pzhqAjOHFWxjIEqq+xByHB/BxS
yH3SD1C0DQIM6gdgoUkaTMrm9vI3L+4aF7JrdE6IAcQp5KHI9NoayOLHuEYJ
kiYdysK1iD1wts8cvBVmtgLI/yqMI/FXoshq7JoCIuZn9zkB/mKCfoNMQKcW
h39mqHD/1/7848OaFVCXJew8pfOYlsV09xt/sRAtkCOLU/qlXwsmY4vZQB8M
X9QPC7HDOXxReh0hwpb09UcXcDRmGrmPCKdmx8Ce15zTJJzTei+8era/Wmc3
tRPpMJbQw3pio6QMUOXtIoaPgJtJeWYctOnrKtp+PRZKx3NMYt/DtZ6K/FgT
YjT/sXl5T1aQq4m5YBLvu4cw75tme0A42PqUYNdUcnGh1AvltiNmgFmJq+Bn
jPAjCBE9RuHJgjlwXo/Ida8hjQljzErKQaV0QRQSox32VGPqLemlG51yeILo
xaJiWHpcYW0G0yOP8io/DSKger0TgCMglIy+V5t+y9rjOUrx+KSOCgacF4ru
Ou8yYsSYHB/gEt0bKtmSbeZzYzpGugU44Vo/B6AP8NtMIFd2NxjFi6Thm1jd
1+H9e2No2lutuR/VcjT72hEj3jpqGyaNTZwgCc/cff5EIxsYWqUh/1cKu4tQ
LXxdfwvelrG7w4Ltf9+dfit5fT0xtUMOb5OzVILOJ9ZK3Sze8eOctljz3hOY
6BRTxmfGYlGHRlow1K4Dxy4/BEEjzXXm/0csxjZGjdxhgmVTCyNAdXbYLEqF
biz/GByhaETXKJRlgKtWmYzEZYN23NKJP60OXexNLiJbF+Eo3/mo/XISY/KV
rNqLIo40Bs0eie60oYk8LcqVtwpG+SZSDfzLB4I0/mzFtOKBjisqPBv3k8x8
8YBZgmptziiBGqnuV+fttQjbaExu92oyVb2qzwMFADP1KeLo9/rYV33GVLNw
d2edHz/yWrBMo88RoGdbKYymKn4vAej/ONz/2nXg8Jsw3c36ewMphmkTxV27
yC0lk7/6LQ8+ezQ/jGGMJ5IGc8WET+H4jlPBAjoGiXkAhKUvX+Qtsgv5aYkr
zToYNMGj8/vt/2SNasC5F5tAQ+iMTJ/Ju7AEkbQHr+rgc0upMHbcCf+HerbN
dIMUNFKKooCaoxNSeSPsi86ZfACzV6cI4l67rnBOuxFFY3p6Yjesb8etlHTy
E7ALkGIalaZaWgAnzxMzzZN0tXyNKNOg/swXBk6+53Dwn4MSBlOQgzJLbxZk
jDdBBGiRKz39kwTtvHOsYwrexwCVF6CR9qV0Yna/cZdqTQj3wlpumpF/X1FH
EGBw0nGcsLfeYvv0aQVYaFxWwgO4cYijpQ/P3mwgUjn4HV/lKf5a0xaoFNpi
GdZyd5GkNIIYg55ej5q1nP3lUsxMNuy3nBL53Sf96g4cVcihgvqwIl2ovO5v
7oprg66lZAAs9oKqQmEdy9ZABb9bDrfbtHoeEivC2vzOB2oyktQds5sV02T4
Y1Der9RPvCGs3AbKaaBxxMJChErwU00LBGJsAkf4jhh6m1gYtIgI09E6uX9y
L1qOSGOev71/gIC3X2SnXdcRG3CsBH+8tKMYdNIlkPX1VjgIykhN/AI9Os4x
qtkS9JHGv0Dnc6eUbznz1xDz/Tv+lS/xtj/H30P1/IKJz7a9Xy5RssLnUh07
sRIGUKGDN7uvdqZkk6HqG5K/vZZwDMCJDhBZQTKFWLCGn1SKXtHd6OJEQrbh
lbYxqQpDOQbXbMCpncTeUkqI/7YoQcBchg9MQ2kYUEWaPmvSTK7xf2qB2yT+
UcGfSuQcXMOvbD0BEPnnajiizeDXjmaVGAkSzR+0RuTE+cMuf1uI5/g5GJhk
+4eQ1vCuTLsyXL0dxhES71jbVBLALbr08WXE2JuYXzZMgs+PqyO/7Tf5m9Lt
jWqBkWMRMjMVxM5vQcaaeRY0gVort8fuVlMdJIe8d27v4blH9snMjNaVWKno
sVhhMTGZo1ESYbeXLG4kQVUCfjrxoK8cE3kHlBPNiGou0WcVyWx3D6yU2205
M1o4L8oZyRIOlYQRaFIJ+Kx6pUTb/0G1O3FDwKipZ9zWoY5jp3rrPHTwFP8b
h1AMk5SAZSjy9TIJZ1257UJu8cbyKeeI5hRm+g1LsXULo7ZM5jYLtVCUZBP3
MHr+kHonmR7tOX8B49IEWbfoH6xmpx1gAnQJB7EW8RXsaR81CCFTQBtaFP3K
PRyCGOtF8VXchJHxsMpTogJhSmrC1QkLVGBu4/dqBamf+g0yswHeKvfOwVaa
OKOmH1xICxaiaPG/RvT2lxl1zgO/8gjFiQjpnzv4yGhxoME6rFIZawzG6ddw
tacPSjgMEoKfDi6RVoRhXABFPwQIXg5WhAQ0ydSnX9JX0AaQScRnUXZV1NeG
DUQhH5gM2Gm/xEIgDqza1NQeWrdMoO2fXw7/m5mOSV1rQ/j9VKaluIxQVGin
th51eXYyinI1w8WOW/VxmxBqfFB8s9hxFcYYxxntqFN8J1NP5kA9ncLCguCq
HdorUw0t9pSLIG1DkQRHTPz4Q7hFH66cn7IgCOqVh/DhnUtcwMXbIvJU9QSk
Vvxdol5bBSbPvMILEdNQ4wVm5+eoxlco4o+AGPY87o+UBBWe4H8XJEW6MKIx
V6ZVU+EuBSNV5RUu60glXaYS07dSs0piNuVj0BZn+NkSPi2au3pmF2vPludm
P8o4fvuUkqx4anPXbVYGFoCDhsxagohgNS1lNO6CJQW+J5kjQ3CgH536dKuB
SBsWQkBj3hDUHdJaQAcM3QoXLRk0HdhvtVIngDoeYKDliGXZvWtNmJa+7bgm
RB3cOP5KL/PjUK+J24wL6y4uqk9FLvuAKyg0guOUYxNULeIUKN4TbImGiD18
ta1Nl2eNoieeaSR9O8qlXUWjhwFgLYmn1WQo+MD6PMfQQAoOFiUQc7FMwtJ7
OxVxYIl8nihLApZnnFCU0AcNvSti3EG5zjjvDBHZos7gYdgX6r0bTJATcIIf
KQIrKG1dYgB86O91YebUor3nHUsgYsyz50z26xO/54EoqldIZWCZphoQkV+R
SbxtroVLxdSUGe2PrjhpufOUU1mLePlVQZlgiiYsh5feL82Fmu9EDnV8H9pP
l8FwBKfMNCn6SflGm/MtLd9YKb17iJv8PWfmPoPdf0YEEUqpmih1uruIRH8v
t9SXEToyDl1CImFr0iFbIc4NEpNd0QdgxFyMFRa/fosuZXoTu3++BdNMShkq
LbCfZIa0ZkGkqnxNB3TyEigpR7FRd74UpXfDNDcDH+ZC010edO1NPSsFw/1n
cZ8q/MQXuxKLeZz2Ama1ZpEhfasFPzuhGHbiF5E9G5eMylEjGCNbP9ILq4c/
/lVSzLQgc5ov7qMxidFH5+o8OakIBzuQZTjx2D3UisoPlZgAWtkpZmC8dIet
C+eJQPyb7maquKN/Z6H/5Pr3XyM2FutcLfZ1EhmjFpXAkF8YtmvadUYRBT6i
vP9OIB3LejLd6IVpAIDxDG47kLpa4XB0H7Z8SfcRWNkUjE2bQSIZSu43kHQ4
Py0Gm/UUpFE/eRj4U7WlDcLkDqYmOKjVWEzUod7SK1PAWz4ofGquyg9MBH4E
7x53SKsVyk0s+mz8ykCvsAA3P6UoyaWTS9xoeeuRqzu/tvEC1urIXAPBaxx9
jHIWjgUx2gcyIhozJBE1hImVgiht6gzZmPZ9Va0TLicKXJRip1UrwonaVObn
3L7XdPIhq56irRxxYDwhaeVz+H/JwwCxIB4efisyMnQVE3kPBt8a7WKW7j5i
un+MNqZsxotSR6bdAwPahlyazmRqgv8N40Xq3ElXsQPGAntlmPisvV8BZb8z
svlf4neDacWFW5LobUEaQpNXLpK291ZdDy3tkdiWQAAj2WatpL3+aOwa1JuT
sNjDUvg0VVzcJLijYEuEM8Y22d6qFJeKx9qNF3ez70fNrPYweEgHGg9WMVen
7qFjSD+pLI45BUay0ge/AZiMtWojAkRHQNHekBGBEUbcULy76f5f3lBlozqW
ZPXkYcHRcZAGSwu3IDmgPsjDFxhiOTMKjAshBCTvePdhaMZ00WK+n94IB8dH
knE3irHPmbDWhxJ8jr9rSpG+gX/ddk8UdL+76L3Gh6EkI8wJx1HRvytDVg3v
rSJEK++w9xrwZhCMLsTh7KT9/One2JJUZM+AaC+JXxTvJoTQn/j32XhuCkP8
S8eFh3Lo8sOZLD/ZckLU/WrgjB7MbxuK1PAER7aBA1ayivxbFfAH65pCzc3p
QThNJ3QO0l/2TtnDcGWYRFNjTFeO8KfN3LtOEGaBRQdRRGVtNK+23+0HLzBy
5lSv/aQ0Lwx5a0Bsg94c1SRZ7o2es27f6s67j8QHL+Jax7yzHgZqW3WHSmuX
TJ/IRdBJ/rDYtvnOC77bdjur4ZHVwYzoT4keZwo0Eg/PhDqNrQlYlkCmSoiy
gicYEf+G9Z+EzlCm7Uo23kHfqsaoLKiuTGLPw1BXuIqRx1efcxlj/qpm4Lic
lV6h5lKUMJxZGRWN09zfYjhp1BqHxD3lp0fyT3H35vPnBfYuARRc9XsFsBvw
kS6qgn6o+bN+QeNjrQDz4skJtQfSBD5CfbksBNs/SlJ6QfKAVufUwv5gRA/x
j6qP+SU7+ZMhg5VYXx3fUnl+OAMJiDdDYqGDSq+Gh2Goop1KGvTLSuniEP7O
3B8Dwpsbkex0FhSIh3KinyV8j+w68AGCciPVnpTSr2o5DxFeOcxaPfiPsziI
Pn6oT2Bcyp61Rt5sSD2QASWH9WmBh5JxXCkGOf/A9xOQrRYKikRDu2S5VUSY
RcMkC+vqjZtR5BFic9ZJdHv5TiBg8mYAFf46uzHhDLJhlye/fEdSaqAOpJqf
gneMIygtiLJl5WPGp58LtNDTz8CcO05S8LV4VkDQvBtKYlxuM6GbbMr+5TKB
ePHf8DTGARPxmZT/fegLBtm8VBiQmHX+BhQiAn0NyCI2xNPYj2caFOhk/tmp
PVaQypWHk8PsHbC3SprGxE5tw8leLMtQTMat229MylOaPTC5oAuOqkbxXGbk
+XJbPpA3jUuKG9yI9yZ3pRbgNkAUS2lkG3tlSRBOA6rqv0PJZhN77rZS371+
qJ88ceUSqkVZmypZuAILtP/fr74KKaR6zBA3AlrocAmQ3F8NkJITS4Gc5Jkq
Fd4xod08JkIIh6n3pvv4SbzjSs4kCEpRTtSu2hd3GMB47NIGVazyGFydDdM8
QwVlibHPhQ6gTmnvU5E98og5eEQmXwKqUWnXppIvl0zUl4NnelBhuvw2QHsY
6P17sDIBpCz0jOZdAgrcHws9rtIfyLY4D7DAQD43HF2lchVyCUB/zD/cqAP4
0Ooq6olYvuVG5pzURVc7RmmvmRb+RMA4qZNZFHvUJt5L7XbytLoj//Zyezpx
RV1SzJQT8EWDXip10Cper80toBLHiLyKDz4QG1DDf7NRNcm50xnCbXgm6yi6
vmHU0igLdbZoFdiVWZlXq8+g40EwUz3ozaDOG1RYoVBN2w77gYiGcwkb1tcp
GEtkDRBkSTamzCqjEG8VjHzZYP34cgyCtu9nDyc/YDGmH+NchEzVRsAQvwB7
5XoaMVsJEZvbDsYuhQBbXo3R8HsjEeLfAGUeRFVGCGu7WPX1Ue1qi73x4DQh
gJipZ2mckPvVva17VNeTbs/4X+QLVyIWkT0VxETu0l6GBILQj6P1I5OEk2jM
JAJjZu22NJ+JtlNJRyNJhpEys676twalrsLAiYJdusVL1UOooUWjXWnqswFK
TU+FfOLH1s1KbtGC9WSE4XqRfaUZYmSj5jjrLt9K1OLf4LoZL27+KsYEIR8K
WUWOagPzr9tKNZkVdTgLLwj56TWyKPTLUroPrex7Fq4kWg/6k6S0joZBg79a
O1BaZmXuez5cBAino6dck0GuXNDu6/aEbNHf/ztNPhglNTnIchNDeR716FKE
LuWAM2OzxYN2m7/DGCI+at5qHk7gyeJbMMzWIXVzkqtvg3Wqlg0WP3BH9xF1
qezDyNxapt0GQLss0fWbSyc1BM8JaF0W33yHrQhnZuFoMQ22vKEvR3IJfUDM
etNEz/1l0B39gZrn20/vPQ8ZpqYYWRMFXoXsrLADbb5uyAbe3zRTUXnCRsX/
821gn2sceT18kijkzZJuUUHCCU8nitPItWZkIHCvD2w/d28uKsnbSPk+8cD2
mFKJkZH3dCD1V8p7wkPjeZY5WDhGPOlDZYhSoJfZ6SEgk7YPu2fxjBZKOxHR
EjzgB/1xRiDO+xdw1N0NSo9g3pk7omQG6TxwPVvLOdCXABXY6IdNafCyGjnz
BGKhz6uCsVCO0vuIxrSjtJl1MRLyIH4fMuFl+qkkxs5iKKgzaSPiktMfj0sY
w3GN2xspL9OJ/MMM4N0r9Cs1gn35zVYbFWfYaMPth8/fxvZKfbmmZ2/P61YX
rOnIUOtvYIXDuta9RVhtbZMBQVFsjk+/emFQEGnc33yqBhHhxQ7yK4LXbiuk
mVCzCiBjplh5noUO2l5UKuN8fwg7cLr3rzCSV8uZW9k+2e2PqEnXeoiXpPv7
rRTCWrVShDzB5BaE5PWS8yCRS6WgB+HUX+NM983Yq4cDi4ymXlWhV2m0g9lS
gpaz5cnYwirXrYg8wDYp9bDQl6bJs9q3/fOH+79BduabuqkQAzen7EQaJ42v
cCyR/CKOXGEK97TjKziL9u/v0xrD2oTA0piYNj22mQUUlkhRKfhhnpqJbFhY
Uf2vG9nhI6YOmRYXW+fXud5Xro8t8xmpuHiy+1JvQtsNQZGZEd3VBSiIU3Ys
mv854SAfhhq0qRkal0/nX2hIWzJCkOWf7/Bg5K1U2H3dh21JnrOwQ5uSpy2O
YuPbFMUgxvBQlxGRiFiv+J3eqZy4Z176uQmyCMSMHS49SysdK7ejYaM4YhV7
CyQUUytsxODxLGOaciwV63iB3+5B4Q/jpUlb/9w5nTu0hmPFNw/uJtBfXeFv
lbpOQWbnNJKAsTAalIsNNq6fb6sLmNvS8Wg8uszpjwvv1G/Y8uWuiAdElcSO
Efj2zDlyLFFVkHdxmo/innRbFTXd4OlVteedd3OjAJDR/nwa6yVnkwkQ/ga7
dF+iSyDwdOr4+OOwyK5tWMqA/44dpulP0XJV8+jOry+7mKpwgYEeNM4hr1kX
+cYBAUcFQBfzYOZoFN/PgV2OhZI/o/LuBIM3AmLW9kXX9wvoUF3EFSA1nI2x
S/rKaFIQYcHpNKMat87L9AXbBzOqrzCPUm452oJarnQsCbK8TY0riTECeWCc
dvIZyjYxVJfKmDy0FU+s2DILS5lUCXmMAvYNwHaBn5/csMvdCvdATOCUiH/C
DKDGYXvY9HHLBZtZngXOp9/XYgZgd5sSC94BAGLkPBiIm9YoQEVWqOlFP3Gd
JEeRZP44fA5JD1c2Ivf8EkOR+F9yCLRvuvU/QuaegPYtCvUd0sCgmxhJrG9G
TMDV0Xu/cbXKZak5GWsEzuqHKqCBW21OL2HCZItdQ2l5j91WhTdA02gRLmq/
btCzKThxyl3zq9x5n6v60CbmfydVLyNPnHGPQ1/0Ek3mT05Ydzvy27WoSyhk
scir1NnM1s2tCVO3Xi3Bdt2/v80TjMU2JsbiJUSIbCINqs8Cse5EcFt9CrcX
8Dwo/vCxZYnL0IpKT5NFvrFk3ZuD555kLsFrAHdVPOj3J6fF4gEGSO2kWVWO
lgaHkZ5tGA1QOICmnxSsoTLnsxi9hLxYdsHC5q21k4GW3KZTRCGWF6AHKnOw
I/DcJpoltvSCtbwNvBob29yiT0WLmOWDBrP21I7AsP2DiNIdkqcUJi7IkmLk
NnElAAw3xlFjzO0yt/PswoT7b5j1BKdbijhS5JlDVojDlMNQLGUMA7hMygNH
Jjdxdho0PwJzSfCVz4cFXz+zTe3NgJI2tDDeZuf1n4KK22WMUtxjtIcqLUQo
Fk6Sb2zCxoH8d+nN96Vjc6u6TGQJXXNCaaHqWEGKun35Gf0EDyrcK+SBsyNU
7i6QRfNn4LZ7sVp0FNugpv99pkKm80Tek90Dch53q5I3qGoc0F3jxJPimHiW
2knYFmB64DYkQ1vMtYdDaejQB/2jYesuEKYWyUIumOoHy3IYpMwAwFxNoR9I
PdjxZmiQfd1zgWvR1UrjzFcyyZ7vkZr8NwY5L6KAoiYF/tL4BnU3c4IMxcAN
jLOlYd+PzxuZ8lMeCIK+qkGw/n18bx8M7yQrBOOot2MICgvGrprjDr+zuLHV
KLwWg2XVyZi6EzavtV/TqVw1UciQvs7a2CLLMQ09TEHOVjBfm60MnSTwiJNi
URs4WWgf+4Ocui9xiNH4dPpnbpazE2Ed4gEQm6msZPvM6o3GyqDpzv4Qbp3q
0CdXN5TyTHSRqr5sHPRM3kddE0hDsUq+ZPeqcYZ+ocpnFKUOsTQjC1JA1EXp
51myYKvhu9GmnG2NFyYBfL6Or5/p3SMzqKhOjoNBI3UrG+qTw8B8FlCvRuO0
/v+gZjveDpr4OviedghtxJbldny0NGntNY57x00cQ7as3/MwHzDXAKfLd2f6
N7clCEUma4M804JRqbKld6ISpHblNM+wWWaId9SHisBS0fV1S9mDpnoEnVZk
NOdDtKHMqlnK/dJ4yvKvTi115G4ARgZGD+hi5MpTFFDywghtw/49jrzTKHAs
t6oe/HoD9VNLFi/+SnZqsxAD+SRbxEkpR6ZSUJafMtHljKr+Z01XMuZfvrxu
YDh0UZMMHkc6y5IyIO9p67n4TaEplnzGDTOtQSs2k8fHdocs9e6yNlDn313Q
kGGohVJIWUDfWYZbwC4nJ6M82/YojlIOFPifzKG3A+mO2nOVMSeJUzlD3//c
CRvMKvkouddRozEOJSbl4RO/xaSZE2Q93kXUyQSjVW266dEjGwoAw1OjILuw
FaUllrE+FH7lWRTzaKUbQu5vlIQMBevqv6KUfPaLrCjDhNr6WQ0YkNGWYmlv
W7oQQT1fHa3vnfpZTaJ+/DB+UqZ+MFPART9CPMki0UJ0ImGVJ6FQ9Pk+7hsM
bpF9gRrkduoJRaiBFcc+HLeidhG62Cz4WMuezrLl/Cp6I0Ly9nVj8kzZla2v
o0DksFgVzq4xyx4IRUZ8CTJ8pEfu/GVA0IJoeP8CX11ZuSFTaubfkNUbMNu0
ssoSGbdo6MKT+RflUPS8YEjbSjpQyHI0b+5xCo0E2Nobdf5ex9ihXOOk4BXP
oEvm+h+kJOUd48xWLc2na99siuMj0X2+CTDeP1oCa8EH8pdyMtccRKSV/aso
aHg1CyR6eCun8Mt/o8foNlP1OpPh5o1/Knfcwuf/B64ls/Vdq9qdG7UU7vpf
s9NxLgHRowbOkUuhlhGsdxi8st4lft62yNbNdtYQ0kW5cu9uB403pNiUQf83
Cmg41PIsGsFGOq0jYzG1SULuT0vMP6pyLO1UQRFj7j4BiE4RxEpjALZDolxS
RtCd8QUy37i61Eipj54S3ZZOZBWrwwqzbI5KonTiY+7b/Hq7lOfMndils7+o
9to9XibqTd83D3xkjOsVTrNtluDG8EomgC+aQN9BaTKiaAKVpwOxRkv3L2DT
KgZgQKCCVANVF8RsOGFUXMLZuByM/uRXOeHGkVzr4a9qr9DuZ0X3WCthtObt
lgZlUw7bVfcSjeIJyZ6JKQHzkuJQGxDV+JUx2ek75Dv0fEPZOmAr89OMSvpL
4IBuLPaVygO7aumXqY/f/NkwpRlLSy7ikJAMh0o5BdcEjcDMh6LhoH+DwhAZ
gNFfcYuRK8lUOaYB21sT4o0Yc+cBePXa5twk+YgRBYKFWqCtMJiY37C3qJoh
Oih2YaJXB4z8LIkHi8G2E0KGekr2RjknqelRQQXJzXmuO+RR9JAR0fElWWlx
cii41jCySJOVzLAN1whNjQOcRxyOYSPLfOr3w5B8QwkwOu9OaA/bEK9R9aEQ
QYm9zWLy10Iv5f3dD/Mv9RIhDC6kJZQa5YKVGQIh9CtbwKQuv0Jaw6tqwMJc
wSoYftGoUOEPry4nVQsTnmOatY7EKLl05XTuMYAjU5PkJR9aRjsNMl+AWiTQ
lftTtkaSDg+xCgdmhhV1V3U9U4OjBoAOUi848/tbwMuyP3wP0X6TzL1A6Ez+
DSXDySYFzzJmp0ZQ8BVAGN2lFhVXUNgrfxyznX3iq1gS/6wvF2kxgL9ZylTj
DQpMbixwH1TltEdv5P/Uz3obgj+N3d5vJGIz9DjFcTkcOngMMVjXV5eEZR/q
tq0wSbZm6KXhLCFoxHTPp3M6mEknS6l8oLUqCRTuH7+Q6Xnm0vCf8rsMAFGU
koxNbfXksSlDBxuaMBLtK+8jN+w/HFxcde2WGcKehxb9Mr5ZKzOAwJwvrMBc
SGv5KLPKS8EGqhA33UX06Hii//hYwst2EHbld8lWVG4Bqlq4CDyh+ojR3Qwb
TK/w9bMkgmsCKgVprqpgXSdKrU/GgmBKRmdUSET4fQKiwvoKItRUHi+Zyr6C
2UGwBXVdSYa3GoIryzGti5eSVwPp3TspyHqKsStbptabqZYwmtuo1VZ+oI1T
+NVg++u1uIlWpWRaRe/XBC4GZ2wkPlMFsdO7bN8/uLd1X4uYhrXpc6reXsoB
lm3X+hRD1q0bjtYTs6a4uaG8KYwVQ8XWcdNVzDmgaNRH3NkIVzsJXnYGzw8j
AXlWpgYddGDEg9FvMS1KMz6A82F4kDjG173eaNtUcKAeXaA3PaeHaP7iMXVh
Dwo2v6a5IhhFA25F0EqDZN8FXv6Wzg5KLslgQl9u7qj7XjJEzXF/7K2Mbg4V
S2fiMZstJ1a5/g6ayqQ89J8HNnG0VR8D+Quf9Ii/vvYTEhq7vsO3yqzfrFDe
IuSFmeA+c/a1kmqKV0hRbyFwdIH7zuCgxLEWiv2ABjWRRVqnOeqHx9jWaUFg
liJYS0PbNgl87T7C9gWolp0XRUKyetrNjy42cUmK+acTleq9B/SQr3BN5DFR
DtKmJa/sEdUrTg0xBJlNDi50TKo26WHlJBa6prJwtnLKmD3l0/MypNE1G5Hg
T432geWU9dR6YOGC080CzvqrDLTgX59hvuaTFb+Q3NE23ro8XOZdJbUvTpcP
7Xx4Nnl7H1SyttapjsAq5dJjgeAPxMqZUNtukeqrWe+moNJF4JoPpINWAjwV
5RBJYt0L2NTAswkXbkm0A5eLrh7aPSdShGhH43aUt7eEiWrT9ZEsEU482bXh
7rCAPa2iWdSLeFZy36RojhV5a4snTpsSmLfGtROnMYHV54Gi5lqT8K7G+Aly
1juAY1zTlPkIBQJtgJlDbewa4uKtIvGhdd5+cfhXDMPyJwBbMEJatuNCoQjt
kUpq46BSRlEbdIF5/Lnea6/4FgPVsK9BthwzKHiPFJ1ii23u2wCw+oxlY+of
GpI2g5WxINW2OsVd6pp8HExAfB/zxjwcvIw7N4pcKrfVblin8vbViWuniISF
2dAOzmtDt2ZEfS2LX1zWDcA9QdTWy4ny6p/Rhsfnay/MjPT+WTd36sde7I5k
BXbXFh18ONQiopFdnynUUUx2+9FbqwogPAMXG6gPzfx0crLBMfXuEXLV8wVm
eQFyzqoBezXZ524IJpD8dyxPNSKfN6od19oTlnbV2/yS5WiYKM9SpUL2B9Gq
Uu0nh6TgYetju3zHy1+KEJmJ3XtBnsEm/JRPyIg+0mdWMO9P+4TfB1S6hNh/
Mq+0/XhbBrIFfspBzm8of0WHZuP/iXy0xarAoiPbTYpGtJEbSqoyRBaJWWdT
ER94hrTsZuD3FQSztVdAEZxxU5B4doEclo1pgvHXTbp77OqgDWIYowTW57vp
gkxl6hBdz5mJGYLra5K5LBaS64CkMtesWwHqsf2cPCeHrlOJF/BWPDpZ4nEC
Cm+ksaR3i70udgH+XDtAQErek/HVut25EPiKwoAuROj2UgZ9WRUMC+6Jalr0
UGYkEfXf2iYS3PqODhXQWf1QRMsZxLn6ghpT2gCfkr0SHSaCbbtKAy5tGJbx
41G93fBIqpTr/3JtmLDaVSfyw1hAdC/dovPe5+ecNCLZ31pirM/nuOC9wfPJ
Ir0gFlaz6XEN+NhCvjCtkuuKIiEtnDeRH4cMlyByqCCIpDy6+AN/jXiV6r4u
Db0xPhA6RPEdqIILxXcTMsmL7VJlwZHGcMovgo3sPOJq5/aIMp1c+/ud7jfk
aex1Vaadz9UQIwlySeKD43LyrR68ExBqgg1l6s0kFp0vlgIKld2ZE3s0HvZA
/Li0Bfdo1OHODWcuRHu4rE3+l/UTrOIzouK4Z5hxCsqaqJnewiBwrBwCPc4R
J2Sh88LwjDqju+LqlDYO4C+/0TWEbGr+Ub/uxdU5HUWcDA0xPqW9uMlncDb3
dh+nMmHOQT5LJm7S6aLSLZ2qiVFv3n+K+A/DHJRLb6o/klrArfwiqV7kKR5X
uSiqsdQ4Dqsg4QoRcfdHneqx2G8jI42Le37YBpfMPZSJ4V6R6wWpk+4NgFKr
PmepUKPlU4fc1FI2tCu/PBLEYzm+1idHAGY0iQ4+HQ9N0fqzBTsSZS67twSD
XQPuHjGb3ZsRjbTXNQy+EM6E13KtC4crrsGSkH2muEZZiJXeCX3x1NWkANWD
8Yus9ve2HsBrC5hsUIPXniDv/aoxnNDKkh55GiPfzcNxM37kN0hpIGXFJ68s
pJT6hyK2EDVp+wZwJQAC5BbGPY/6RQRqx5OXtgtgDhyGfWMh6ud+ntMciWGd
hUPkOZT+jgLDIgEZdEPgC591O1QaeJQpLCZzF3sG0dnvskJ3w8UIqSs0kvM4
mIqjk+Zl4bmd8YyzTm354h/azFDxYzq/uvQO1NntBWJkhSiwFS4I+xoe59IC
jYUS7ifybVPXmc849GeA2piBC11WHU1PvLMoynOpzvia0zNw8618LCJ6xzAn
vL9OirGqGAY/jrawDyMDGpFxK26jw1k0Dyb4XBLhzWyi0o7vaMMASRdXXD5Y
aWqYxt2ArxaXSVFAFXzYS8ILMM7AFxbv+V5u0iTmeM2wwHMlyPLoRqshkxHH
BZ+24RgtI6fvYfEGTj2TfiRQy1Mi/aP+W19L+EGjMCUWh8a5SX70XUK0fLMu
X+xJuQqsS4pVislHM0HQqHxKStrR94scWWrEaw1Lg/Fwsq1o6PfZWRup35v0
ucT1Yksn8xAEBRa+77kK96T5Th1Z7e03N4bW5rCLWC+bvHnGKaPJJmFDrvEB
/fAh/Xv650tkhgtveJ4s4ClR3TCwiKaa5f+bXkxpR+GuSTBJVpKYGElg7nCv
qqMDLuTnU356wEnkYDMfTYi72jybSNI+5IjC40il2/qpYJLoZ1jjBMd648ua
9fpfzJWc3+XzJCghG54z1gK1kpA6TMcG50U9YUzKT3w+W8r97eUSYLEBoGzY
6n/4dPtGHEi4o3j3eQ+h/qWAAGL+URxUdjusXDkWsXf9QA5YTSd5NM4v6dRE
rwTgW8bmGZUNc2TC/5aNBnW3Ies0rg+dX7wU4plkzyVEpcckZpmT2WScAhl3
ZwIqUPDN8Ip6TpxQeIhL0ffcRS2DpJU6pARRCbdzOZDFl9lDCMA+RLK4BE+k
BTjbrkzBL/F3/P4Hv6HBri567fJx3fCqpEM96jN3dvp5Lw2/MKntGOQf0QJG
HoUediJYZ4ZdWJb+clHvW6+V0m/UkREwPlkuQLcmMJdLxuGIUuHym/XzSrqj
9SRW3QPDjNQgeRAv1VaeqQjNDwPl6YdLc3u0QIANO3TK/ageVSPrNNOkFJR4
zm0EOS6bRga/PshuE/0oWlW5UCiSe2f8hzz+aCaWS3qApjcHAjfpWp/mx/nl
BDJTOaiFLQjhQmMHY5cYvvhp5ZgQ7m2Pl4NdJplWWL+EIVyAhFcgst3Lijn6
Cvd13s0tK/QjWLXgWwdCJRN34yfheOwSJYjbMj4LHLcZzOnCJuwLnOGuqo3C
CbeqckYYDqDkwbQKsd3lbq3Ojvo2Vr130BAavgF1geLyzqm7FSISdnEgBXXz
xiqY6vVoC7HqEDEKhH9x4w6OKGizJoHWsWd3jWcC2aOH0sCYKPcaz7OCEh03
bX2+NzBl3HBYCOncjmdJmHGBAmD6eh0gx+XXfH/IcVsYvLxW1aAI/rgbF7Vy
wAbbCGeRAl0b/s1OpthxilGr5SkdFdVbP4FUt6+asK5IVKd+JjKv8c4cyDkT
+Qp2je7Xpa6krJ3msOGLOkJek9c2cEFibhyEA6NdYM9v7si/GxP2MyUbxuTu
0R1fiNQr68VUMJaPDYaBu7WZo8zMhxk5sGyEvABGfl+N/9MxjFjVbYsALUWQ
eK+8sJ+G5szaUMqM1FuVs+Se5TODnK0dKJS+XGgX30RaAXwVzCfxg4baciiA
Yu5L0AYTTNYcXvJ1piy7YKYuxjkVQ0Dl9kxPtKc0hZc0m/A9DivBUtddXN2k
6NIhEN3y/hV8vFYLpM2iXoE+SOoldM3bVSzUAb3ntZskvn7Bwtm1QTIWyiTf
O5pR6ke3ePNBm2g4yDGChpvrWFA3fTXisiUbV5bmpnvK/wWe5OqjmMbCfdjs
AoRen95bmbEMaC8UXm4Q9CkcYPROVKeHRoP4sRLNqxqAuTcIErQxBOOyFk+B
PS0RIOBLiFZqX4zrGbvkmUN9ylW4CRKt0QX9YI20iKlZvenPV55Im21Fo+Ew
om1qJ/4EBOS67zCEKacdTAlmEMMKIpH7FtkQMMdBq7LrUDBWoyyZwBagM8hR
qhbFn8UJjbyer47xPAQ7CymKUYl7IfSOF2koDumq6CNyH4T792lvwf9NZgDB
qoJaAv9Fc//lSdEJ/eI+eCcKLYF6+A/HW/9EOdBgvRnhYauOcOFTJQatJh0U
ySdO1NLiX+59NsMJGaXHB/CmcAACs1OVzVTeQKZ1jR07fIzZrRhgGC/lx48k
2uuvb5IhV+ZK9xiYPB5DmBmd7Nwgyo0+DFM2X9D2RZaYxHrC2caGgqBie96y
/ifrqlK9Qq2bXQm7pQIyg4o3r61twkR9oM3dpqAmRcQHeE+YQc4Rmm582iFk
t9Bf239C9kAdlDpxMX1/SI42EICe2NqCXgnRxLshrRwNmEsCQmpAVbgtRCym
7Nveef3Imhi/vkXqQqOXvhOB3YRO4gYRiCaZkAadm1vCixnlWFoxfEuabKAz
FAzXuaXuwN4WWsO2PKn61MjjMlQjyBjmICkvihrN90MPdUoGgdR1GJyFaDdx
nVVcg3uiPq6rdrZbV7cYYh+7vjB5PitPhja+VdG6/UYoVPxxWNvpgC0oemog
7ilSOD7pFm8JTKS3kspZPf1ZaPx0kdE323FEA8ejSUzyTBPYx0X+aMGZ9akb
HE5iqSWBIxM3gJbt9xZRarqXF+YZt9/dg7k5BrUD3idc4fN9cQKt68r5+OuR
pKbcceBIhx/kocI8wZxEznh/QoyOCBfmlZr0LFYf8y7SnJGQ/Ll29al20w41
b4qCM1DB1rgjaq7wKIniNbkKDoJYR0wwGW1WfLEKUfHSOqHBZaHtiYynovqe
Hpxpx9RVsKVzUAtfe/jZgiVUvSQp7i3u1PvPE1BKlavXC0LX8dwesWS5Gt9R
G5YLLKXibcbzDRs+MFJstr+C9EGv5J8GJnnqA1uYUhVgpuUP7dGuR6H46qFz
uzbfe2n68EeVktUCOqNNvsc/0AshEW/MgEEiL2mTfcX7OorZoOTDhFRoWJdM
XtVOaUwpMeSGViyvondz541vGAiJeR9MhffW2jS5BqbevMsjHJji1zfh1WGo
XMfhhucJllYuJUiyGOZyURTMeAaDK7IzmUHMJVXc1qCUavF9H8iQL4d/67uH
1D6rpOJvZAmOr9HfJWX03zfU1B9le3cAhklJgFzni16elPtX6KDySn6vsJPn
niAg9W9mvWeeu/LTuek0osh9dBAEh+JH3XoS6RBXgyP6jCksLMgBq7nge0dy
QwG0MBYG7bjasP2tPDeKUd5Gjg6SVw2Z6WwqS431TA1Ap17ukyOqPQbu+N27
wvFlY36wDHG1puyZ1kPIdpTkB50mQg5TgVykFmteKI/2iMkjrvR4oliCdPhI
Jqhd4pBCre3P+BNagSG6CPJ7d0VvLWw/J65Px/qtX76NyRJJ945b2M2pV8EW
1s1MnU05FG733gXk5q59Sq+WZ59sR5pZ/vpAuWMf4dP2tVxgGNwF3Fm6NXwr
6s307zpAnLcZ5GY325Uqg5P48/dr3F3EZNeSrkynlDNKsj5hY0hRDEM8oivp
G0IXDGdsiIv033XQzEjHqlM7koG/6AzwAuCPfQRkBWbczjspwXFjU+QXqZ+0
BTlUX8+ZjVp8wrzZ9PbT2AWFFOBNP1V+dLSrqQOR8s1+ZW7vbugLZBdWEHVa
HGdYEeREqVLRWgijXjfQ3f25PKIC9y/09kzk6+yFaz27p6HlFRCiF0EZ5Hza
6bJ8Li7lzz01nkVv5sMaUjNMMloaentoTdNWwktTdXR9SkQvjjyMsfGPai2O
9XoyYedigP4SWK0Q5jvp1G6LndOF+ybkJoz2EKF4Gfd0vYL7tMTaO4yePVbs
YBRlWRHkPzYujeE3NjwHAuPn/Uj4F4j9Pa6bG3nzD2ChcDUCRvnuepCaKkVS
TWXH9cgXTO+W+2I4j2W82439JcSexwNws6rDCbIf0QiJ4V28DutQLZI1j2r5
AP+p1rmhkqZyvfm3NWvOYPHn1v5QjaD+ZhB6bU8aT1LJG2VExnrF7+WCKJrR
eQxFIN7w6qfb9sMACBDKdR+P0bCXrQIVziNgEAYSdckpe9+CAGrPbXQHnb64
Govo1gz8UAZxEAVcjS7tm8+MXpUZQUr3V7cqQgLo4pXjHeFRZNdhbZInLHaW
tolaqtnwKdpRo+oQDixHI4UAQUFfCN8pf8sbebNT+TjZnkxM9KU7rzdIrbmk
xECxeq3ylC60P7e3fTUhR1J1+NJlXmRrtk5KnmWtqjiein7xfJok5GKgH51g
ugPwlKfaP2WzyQSu2qNZNmGBsnC4qWzJvZhtB4ftsjaz0wVKtHg931W1UXoh
tWrF5XnBBzMi4XxDqT/0JHDs9VWEtZPQhLPaUYmnjceqGfkqvyqBIX2F5jSi
PbzHwrE1H1FnSvxXfE3ZJf13FxvbI+k/GaKJm7T9DBblxLwtk2DTQu/HQScR
hjYQh9BJsqQ4+r7ooIyFgdnSO1JTy9p/nHZ2HP7h36kTLadUuRGwQ9wdXTSi
ASTmMl8qxoxreO6rjkztXGkshZK4T7jeqblFQPrW3U7k67goSKZRedWQLBBc
qYd8uhX7kZBbypxhZY8tAmk1laadfcWNrNcb69GSUiimsLU9IqUsCl4qSxdl
Sddn1jwhistbkdIt89nkkis8z2+iCnHcHaHYCtqHPHUhf8qtgLbKRITvvO6N
lgWW8u5xiybT+QVOEoJ+4QGXxRa5w67ElVVnSr/B57MgEvxs4bEs7AHzSAHB
4tZantKLQcIurww3Ct+fymBbptOE8A8SNnLWshKMOQLoW8od+KAC2I3mOAYN
CiOmoRd43PNTKv5giqxfeFWGcwfYqP8kAggb4KenRXH12H1679lD4RAC6T2H
PygxRNvTuXpA3qbn65Yxd1eqUFtdZ35/sZ6z5ljqGjY96pNIbSdC7QNQqwZD
dVI+el1BbX9K7TZANxR5NQVWxb3jlCDQE+Q6rbd2oi2rmBnI8URJscE0bBvZ
ITKm77CfNwaZxHtKsFWOo/8ej8Tj5zDPaN6g+TD54ZJ07u3Si2hf0j5SA5NQ
jIzkm4XR0WXixzqYoWk0VqtQwBpIMbed4RqQfsItipILtoMBBqQwdnzqDCIs
MUK1o5tR1a4wahZz/luMO+EtA0ym6HYAESNgUROq190aLrC8kQtvha66EFCK
Mdv/qwEtvLpUTplTwkG+J0OwtC7HZpgjn0n6wLj7xqTm2Sgb/p7aBZVZfM1c
ZkSkGa0Rx+IFY6M1RI5RElpmqdy/rVvFRDNOiOYRWsxsrlnIKSrE51UXSPh3
f9Sc8c0RsEt9AzSQI82+EW2iUwkRGkUQwZto8XjaVKeqVHTJD76vyfAtP05I
KTkRxKfSLzqAoQgubG4tc67JM3u7mVncJ+1X0TKIKEdzofpD6Wd35emvN23M
dxwFJW6AZn+xEDbUfOdUPnnvB24xeYmMjN0402ZiqUEMlMd9+O47gr9ChAsT
km3Onf0FN1oADwyeMnXW/TzPzuvTenTkNQXIFFrLB7J0lnSnUzHNi3OB1uYP
VgwRuSEafRDyOQFGo+N9t+XwIVHRs5VDJf/jgeu4lUHqswiuiRtDC59h6FLO
YzxHrKPi+YO1MLY5Wf4X3huFPv3SiA8iMP+9JsIz6ds3z5HfoyQlsUyW4JYR
rr8rppREqc4gsR5B+THCIkWyp1Rm10e8MDv1N4AsVNCLpdf/t4ri+6HM7P0o
c7tqidefGIOjHhKoFPnxc3qqyUOIWlMgja2NxgZ8GpFhQwiGrFnuAZkBw6m9
Awdep2P2rLoACCsE7Ex4+bvhIgQtf9wQ/GEGF9MVpSA/WC7+olNht6B1pqTv
yqHkKkNBK1exFp21JHt/v2ri8dDZXX7Sq0m2utij+cSWl0cGJw/cI5+mFvR2
0n8ckxdJejlgpmeIJ2/lkbReksS5emG5L63+EDjcK75vTwetRwLNvlDizfu+
GVQWELuyCgbqZsIM8ygJCLGmCT6pUAI1DtoAtyH5tPHu7asIZr4wd7WxNuhx
l4XdsagvsR4yRUbTNY4aUC7c29kIH1UXxW+CFicDMFExDRkmub1k/Y7MaZGM
GbvpPttmE8fj2KFW+5majmsh59paIa5S4auns9o8ODlD0Dzi0opp+hSftPJK
olvky0sLMUbV8O8I0wUQ5rYjssJr/kSAHGArgABCD5evfML6MlToeGzM5Wnz
YFx8B2nAcw9MArZx2fUCJCKkfiFi7Pdz8uYKSJdl6P14HNSDO6ew+coQG1wy
ET4tKCamVuehtFk4XiOdkczg4Pz4WnoKZMsoHAKwk2iN8LqZhZzJSz6QwRud
Icrn5RpFvv7uHNe2JuWlKVKtH7pfc4eESMb8qOmkaI7Y7klVU7oxoNTMHvDf
tq4zuwcHCWKRlgCWqwwALGMcOpdmfAPLwmtV0duL0lAsNttc4HJYfQ8+ZqAV
NL8xXkd477Bj1sTplMJMozcdvkWH31OYyjqlNZPIW7Ka/BpKjOmIHlDlivc5
oP6eEdD2GqaUo/bKdLbda/VQglK/f0WvxBdDhBTPBC6hJyjqKveBlsu1VYrg
9rLBHr6OSGMvt5ZfnOoC8moGx9wgcYlmV3kPCdp93TmAxfadu9dOPwTCywMd
2VCjC+l8PAJQYLktY8ov++M3gQTAPKBT5MSVfedbVlkKvzxiCXdKnDwbbEBx
ShvnLpbEQhBo226aOhEsSYH33864B4VT60L8UDwRpYQu0ufW3qW25C62E/fW
+qP/LW7/Bm9bTEqF+RxRl+cFkkInGiO1zKJTP2MKvP5fQ8Wu5PrLO9+jqlE+
QUsf2CkUEqibPWvSKuE67Byx3EmvMVA6fbM7PvtCSRKjF8VnAk4l9JZ/OJrd
ZuV5taGtmg/RglgXxYkqKrpvzbgB2fZd1EojlymyI84oVG4PPyRmqqmUairQ
Jgou1ly/1+zr4kvkKgW0AJurCzo3LzkrwGCcP7o6ibYG3DV35ty2UVUKwj0I
5ru+FsFZEMRyIbu78OyHeCOxhBORNUO8mgirDptTfq1Xc+N2+0YA5k3feQpA
3nTnT3FLezfe++Oh0dJIMKftWtZLsEiHESQ9ptwdWfElF3sKcRZEuqmFlGP+
U9F5e/kJcnDnrbTvqyei9Osa+TF8EXXOUN/SI5kz6FgZ2ejPfjnnh97DPQ11
InGJOGpUx7nYCrQRv1ZeYaqcTQVfTXT5SYGILQisoPmdXP84TuIhSmf1eiyO
U10QeNl97NzTxSBWM8A9cuIM4WssNR6ab56ZKyNXaEWT6dwaRZqKyc1nWVtM
1vo21xgvcyGxp8UGgNBibqlN5MB2ujkGl1EczZ28xuDIjohBg2KlLdp3BWa7
EmE7nurhgr74OEPKuNFN67zR2ug5kGwNwKUURpBWOGSfU1L5VyHS3bo6RD0U
8yr9K97u2XWQME2vi5efpNRuGTHJRrOPHDPF//MWMlIiqVGzDbgsQVzrkA2u
gxM9usBxxyQdNN+So2xcMOxUklyAwIJe+fAbXTijLc9C/QfVUVZZpn75F5zb
EgZkEU+r4Y4xgwsazsQ47Tt7wNaZZEuObgqKqjtjieQXu8r7IHOdwYQBRT3s
ZGFP+xFayh26vClH9jeWL5ekVA1jfgi+f3GF0K7jbiveWgB9RrC4FDrq+0AW
Lr6GkKDCl2dTJW+8IyosPJAvRpTKAwha8I/3K+HoNesSiTCPHPeizsA3SsGX
ka/l1ABWDFR9xSj4AG8SbxybIoM8G5n+X2oowueXH9pGIWAthFFDiaI8hFhH
PneYolr2gH99he16Mrk2tDHK6bRUjfPMIOLA+jQLAEjHHh3rZuBvVQzUvolA
1tksPEx69E1lwQT3RSckwa1fRpBfBUJ9X5vRz+3Lap68H0tgB+/+wBC2x/zB
EyAMNTKVHGMTK7xbxUz5U5eIGGd9iag5qR5mMPzDzFIi2hgAFrmNQw3ItuTI
fg0oL728HT2yJzThmRXnAoJrgn/ED0hiJ1MGdtweAm7JoMjXcWI9Iz8TIq0H
cPQ+VUROHJrCKvN8+ic4qHE/96nUiZOyFBp5f+wgPs7RLb8Qp9MfBCl3tAC9
+pfUxzHCiuQQ/vXWkQJUYnpYPvWgrrXRrTrR9XLMQk+SbIF2HwSUO1gVs38h
9D1P1ZTAUI7BfD+0DUOhwZdSh/NBn47bquRCwX0x+GVdnluBIXNeEJEsLCZn
uzAqiSu0QGL+lGsk8GchNHh5ja93TrvBzXVZKp7UREK6bc9e4r1YkwH04yfu
FCZyxOgzGx16el4c45EaAEsVbdjlW22sLc8R+dLt8CrojFuuhBHPdv1w/S9T
EDzlXhFGK9jodFgJYnW5IpVRpGWh+XJLkt6a4okyVnyA9dPWL7dPc8B5zXv7
9/NoR3M839+aMe5XnajKaThKtRrUT6LymlZ3N1Gn9feIpUxU2jb5U0qfPhjL
OVBfMzeFR93ubScz1n6DzzoNOJ2RwNirxQJoglocpSwpPDfX7olPctoBA3xA
Se8kCyec8bjVQ49hejWZGQFrOLE7aKIieYHoysbMAlnOPOSjY/cvE53KabWg
aNdcDcLEc5Iw9qL3RSKY4pGrfqEK/CciMZyegSUmdOdhvGFBrqXakPzZLN4y
qNVs3HkolTH1EOSfZVijrFGAFVJ4DhqC6IKrZ7rXQhq4i1takZDNWCVkcfZW
g6I1Vd5auO3nfiR5OfI1b1ToBWfU9JcjVEMozev+STjnpJGhxOzzgLzCKhNC
Ihs6cyzaI9Ko7GFbq5bL4C81xIH+Xjzso/D2q1dKaEXOJhSuhjz7R3FRoTC1
RMXa9fsXXweQ4t9L2/LZWNRhU7JsAT0T2tpP8e42bRl+ryPwxmygjXgaCilm
8ymsdpR8axHBHWqdCddrb812b+6vGF7pOazpLaR2lJmINIX72mKfoa/zQ24X
RQOjjO4p7wFupYo2oi/xR/zxUSiPIhJqnSG5YV8wYXahlvpNgWEzQe2USg/M
d7dYLJxXCqRB0J6MJgI9uWSrXPbISl66J9zgBmDCR42afN4JprK6NUsL6mKU
HUtMqMaFxTwalyxVMxVjzbfPaEeW8nnGNLI2rsIugw68DWi10+n6ksZfKEz6
to+Km5JW2QRsD+BUMUs9XpOYbIM9NEvWgsHi8xP1B7jLhEbnPoBfTVGi4MqE
TMzP1QL+AmufLqjFoL5xqHKzCC9YARcRsFDU+JdYcAFvc0B/rViog4ePwYie
AS0WeRyznHsyiH18bZhciDY4Oe7hqFnZDREHhDGvjXQl7hXYbqPltdaO6Byq
QMsfqkizu+cXTkhsLw3H5Q5ny2oY+8fxK2/KWYEzi5HllLwXOxl7RHpNoJ2s
Q/XAlhBseWbdXZtyFEMtBDg0ai64y2Aby5eEmMPKGATJK5I8XWaZsxvhAsyJ
Qm7KVZ2aRx9+8wqDbSUQuyhRZfX9fAwbytkvborjNM/aHx3jiGtChon4sWq+
aGxazn1RBxdP3yK348wQclQFP6M1kcsd5KYQptp1EmBaRoxdnXcsW2QCsNX/
GUKw+tcr7yrVxHbB/0PZw4p7KfPY5lZxjWfdGFi9F7BCCYhkm30LbOvHvrWQ
ZcdpsbYKQ5YngjG4Sm89NLpUC7HXPV8lu3giEIa+OQ80nQ/SZy0G76tBzeh4
zlDJ9sLJRrShENoT6/3yBMA0JKowudjAuC8iYuDSU5yFm4hf1eYjwHAsLzRq
876UuZhBGFhJx/nMQQDhD3cUheYuidggH586ZHf3xWOqzuBTDbN7GkQFpVLz
WTpDnomFwlMeWKiz8uFHUkZq7RUnv815JE75k5x6Bjf4gRLC+xAzKSqkVQp9
Y02gfLfrwqrrSvucuQexWLPm5fisVvBfR6acg0lIzJ75yC5SQYr3idoiCDqR
6q+PQkz+NVP3nZIKkev7c48aA5eBxa2jEovYpnRlLTbbJdUgc10gkJdTvKqB
vTaXbWf2JYkY+7TUVg0jy8AgWLOz8gHHfDIAiPjkBYoHP/9tAPVQ1LrToX5f
c/zfcnYkOOFamNGEtyhjFBG+Um+caxIftJ1CXI32wIpa/fpa119+PE7ouvWz
egkLzwDyQBHk3VXG/XY7yyeFh3tmYEbSK7tFYDH0dx5AO83Pml7g9svjEE0n
Q0Z7KBcjnyUv2HILJMxEY28c/BxMtxEZuYRjSZxlTp8aSqjcEK32W+48jHVW
v0e0k59KC3U+1OoRiMfLprthk1TkDIIDEr/2E3XToTJelzbQBGYvQgsM7CqL
+JKanYuXIMDH16piPXlu0nYR3k09bWVMGjEnUJh9i/m2vuptAfUhjIaREbnN
PMReDWr5QnwSnwSDZH5j3PSZ7TfHglKK6bDdfEA2q85RX6uxG993lHT7+PJD
JFiVJVcNa4dsIJ3zu6idQ8emyIktB6QTypcgAoJSFryTdELLPaug+6ogKt3r
De9dbVnmdtHzaT1fVQ8eDdzEAq5UdPAnrgSHcHlMeULSC8KXJeYaygL6U664
R2Ca58yJPD9kaKNqdnbHxR2jYoA3mmdu6EMR3S/PgmrCZ1c6ezhmZVWzI6+L
QLMa01YJ1satqVQkKeKYYxp+k4OfbHqAmjDewFX5JkB8GHXiVl1DzmfZcmcv
eyYlzqD3m+pUF7v/JF3ose8zcW0IhPAHLKDt11Ab0IQ6cR9BAhUW6rAN9Aj6
ggzv9slSqXY8VQjBwoRpmsiDGOyf/3S3sMlrOJmp2uwa1CCZWGQgsXaieH0j
w/d/6/lKBRiTKfvMkmiXYdeVNeqNS3Hdmt8Z+6rokhe5+myzD0WbYN3ENG/m
KaHlcd42U6z07yVb9Zeor+pWD8GHfAHbwNoEZc2jMBArIiDZ/2t9jvw9oOwh
30t/tLvKiT9HNnjZBU2Cq5JtEtXOMbc8rKuHfUvF6wfysGP8qzqoJnXZPlWg
plvfKjp1nS0Uu7jJB3pcXXWn6JJ4wIj2J1DfXIL+MViqSrvrAyItR26xjrCl
XIvY3jawZL2epmyxjovYE6RDk8/yrXBqSN3Aq4amAiokJ3B4RnJVI0syfAn0
I5eoObhe1ygw1DpRSxY4ZjSCiuD9knzuPuw1DM710yt0mwXAUcIhzrsUmQOU
EzN1Yf26DcNuEAc9dHHaiEEpZxx2OaXMTw3gb+dfd7YdLT0Ik8cH0VwD9WyI
rdgLM6gl0q8X2VZK0XGUavRarRiy6SawbP0/48xjBFUdkejVYcC1wIDfj6ry
6oiUA397UgKUDgUp4b1LAIjtpf1lSFzo1arTQZYpCOzkbsN0U7q5aIC3vOJP
9AFSbUV/i+Aqrry4HOc+70sNg1AA9vkwafFsBpJ2ART52tqlojnxRS684DG8
6+1Et6WRYzPMy9DU/duMaL4QoXzZCLHutPCaf+mZuuezWYauNofqH2PEvpr5
AMW++xq7NAFtS84DwT0Ot/r1Fr/0S1PB7d3AmCoCOpQFmeALst/NCtL7FI8c
w7rBdsTw4gjbLgRHEUZTi+ky3KlPpMmZ7dXDxjzd/QB8VRwa1FVubpm80qOs
83KRBpaJjCPTDRUCGKJ9kbl139HI/0w24DYakmnVrIGF5CglYxSKJwvRnysa
/dsuHeAWdSwghbuopxu+Li65SX7Ncmb+VB7KNaKo3VUiYTe73Cd5JfVkihHj
CUXpS2Pa9If2aDf7BB18vAxJL0OdvAqnKL96HZSudofNiv81FBG4dT2/Kyud
DsD/OgPVm9P8+s6CsO5pdWWJrKvlGm7jAvNU17whhlCwfZJI4GDTZG68DFZU
fIPtLb5oLBk07NfSmpSBlk6Dnn1cQZ/HrNETUADm565ST7AglSgeBzIlKESy
+axgpMzcAEudwnseJQ1UqtyLhyINP3ZsF1zzBajv+Xk9oGKhkFZL3/HHXfzH
pj40lTZKgCtAO2xBmy/qmlDCz2A8UleGhxA6UJ9P9Pvprltma47SATsURALE
dZ58MLCB+sF9ZaAHmfN/rYzVTKevXDaYwoArOKAaf50mBqP4od5FST9S+W9A
otWc9tzzgfvcSsSM2mO3JOcrK1YKkrhHSgt3sOyQz4HSO+y3PHF+0SU12Byo
Lp+smPdF2Tw9ct5ggBaA3xMvl9i3aXsmcBBo9L9av8ObsrnDvgmmGAea+0B1
uucTSmtrykxRGtcqhGyfQx4VcD8DARPRFxkzopCZi7XtWCeY1ROt7uaYHCDv
gIiSp4/jw1gDnQod+8RaLCojw4wjpg7HgjKzscvUtMH0wWNxmmojZQjlbNWp
5+l/GSiUJ2vIEQWFrR8fZVwlo6WaMPBLAvaKXBhI+VvWZ2miWQtYJzx2tPgl
EysUBshu3uZvB2DuyZ8e5IOfuTplOSaVqN6oMgBeXzhPTZrELvGr0ya8cD78
VuxWGG6ur8yjzKwpHZk2iXUdUgc2ax3OvLiSJ9+NBAC3n3rq8zowgJgfa5kN
s8WAo9ECnO15xnhmYh7qgPNRCoCEmAmUv4L7S8MxkXVsV1ZzvRQ8FbuWA/tu
fvs3zOVOmxfq06ORtWwGVOyMqnnux86hR6EL2Nvkw/LOnQYff5qKRoatrdWX
VAhB1RHrhuNPIilFYy4QEujTzCQfi/j/MNxwW7AMUK6gQFn16wsPKUDN2TbH
v+jqy1JB19HwQcRSiMoruqx7w+e173BahvjhdtppX53CldO9zmaSFGLRwfa1
eNwrzvOt1AlVThFeW0SfXyKHoTqU4uM5DCb6C5vPHC0mHRUPw5G9JpVN8Npb
I3pEb+J5+gBVC3DG8a+l2pO92vCQcBLDQYYTs8UTzmMtacZ0Hq+aiON4nOzC
1KabpJftsDrRelBcESYxg0xNowkfIAkqFE5Wxw+gJ+NpN5kvdAfFcLcbXDL2
Fo2AH2f8jvWR1Oyb+SpzFfVT3UDWOB93l1Bbwndy1/95hFZwrkAzSW/HJRMa
/DV3qHkRc9tA8YAmBYB9WABhzqnoCeGRrYtHkRUj1YPPhnyA2x3jW6p+L57g
3Q2/7y/I0RXSYKhusXGOGJqVuqBhJPBLto2uJGO59JS6UO5NDoFIeQ6zUmyJ
oCDPg0lFL2hcCIqk36SMZvNTMhZVfj9N66pss7CmR5MlGMZgpEz3IGajZ48l
ovGqFqM20aF5eCLgKcdtq69hEvzTyMgcPMHDoiCuStniJY2Z/qpMSKuBzLA5
+SgapkY+IN1cI1LgvqX0JNBHa58yr6OJ8BSzhZ2brkRjufdFX+eJJUX0z0Ze
txniG2NTcXyRbtU0R8e6EZQpgA7PBvdi+kDH/3Lhb6lFpwGLju36iMVVN/90
Vd9FR0QYHtpiskruBiHfz/bM/gxnKl3eR+t2I7NCiQrnfZWl+gekf4EKyG16
gi3jIplDVB2J2GXqpq71Ae37dK+XxGehrl1Db4os3iyq9wZTLKC01bcJgslA
AluWwYVI7wMuk2yguO2vjmL22VbulJ6TSIViGgUwfn95eT+VO8WQ1joiqhuU
09JWJrEIp4Uly3oC1xF/awKa3RFWiqcTJXpCWhda7tkQVSBgKHCEZ9ZZcXtE
TNZoT2EoDUrl83Y4qXHWoe8ejDCi7smyqCSc5NS6jyecoXOZrNNlBq3glXo4
rYrBs1Q57M/r8wfFjUJ6wuEIFr7Wdy3g0LF6kH6O1MPQ0NYThCECTxMh1Kl8
EBuNamHAS6TWeBvPwV7qfXL1D/8ICZLK26wPalt6sRnsnrqTZyKSUIjLag1d
Lni0OEsiCxjqYDnTXCs7kUbjiDJ9Qqd2qyPTBbTaQc6btfOqqbxehbqS2wkg
PRFepPbe/prNVvD31eflfZFnS839245tAZWdflR/7e47WxMjoB38Id9MO6th
HEl5C3wzgH6kUDme7QrejLi9AfCOU4bD4eYJfYNGnzCAnor8iXIgA7p44uDz
pZi2brSrXI0LJ4rvOAXH5rCoH9r1fpShjsuhooCqLx9R/dt4pPnKloVWUKRL
GQIpfP4PpNpAru5CLtPa4CNZ3PD4dhaUqXX6a6oOw9da12ey3cwv4pA8953+
QkiGDsPmfwZotkTEVxhFM0QrmYj8AAXM51/16/cs2Q8hHqW/9dPCsLmZXWQv
f9ATeXWpYQOeOjCvGCGKjd3vGTuEdRfXMtGh2Mbv7Lf8Jj2IXQo13wvfPgEQ
Zz9r4LqBvwlQl1VKYOmbqEdEF+XuJ6F0tzcHfnsPKgUWMOmyj0tRWdwHta3c
lNNa3O7zrvAxaArfcBGEHmD2y0O0qCW6Ao6l9FeN/onyclAMpIyOiCEhXXI2
oeeCcneEBafcYWGn0tHe4RydhtGQLL5RZrwPNtbCU1zh63UxX4iiqYzru9Og
kcm0A4kNbTxtJM2Eg8I1enFATVIRY2Y/+AagMYvlucS5o7r0c0jVep3a4jh0
2SOSqXmujKxdHGJpNFgZVbh5a68iQtZ9y0tvQtEtPS0nyS3EyFUW8XR89WKk
q970K8YFyAj2NCG7up2k/R7MBe06TDGAE2xYo4oo42wM1jdVl6puH0j0wJkZ
Xy7DLYsAjLJ9RuIGXdobATy8k2OmZzYbBG80RSstJTLhuMns5b6DOq2w4qF7
f2GzBB6RFohnvQfbqn4gWj6lt4YRlYdMjhAv1S72Ay6obXlEHKjsszSWSian
+jpU08bhd0ULp0AZLm9EGqQh1tW+nuJUIJ4Zfz0XT2uF5uH+uTDS1se4HbGD
eu49+m6Woacwaavbh6BdUfGvZgXiDVyicMjRnOvuRKAXh85igD0u629/F8SG
ZPytazlgmEMyq8BvvQgC3Xc62Qw6Uac3LD1A1/nCvUTTdgAJsVR/ksz4oHkZ
HCJcwsJqYHEshV1jOoJgDiUc/Xr7POyyXbHQ3Gm0x2qi+n5Wp9UrlwrII01h
68xeJ5NCU9UimO+oLLVH2qmNKftbic4peJs5aPWZ5nyyBQT8ZyQnpJm98mAT
GDNCyBziSOR/SUKOzer1chKZagHzRmFS3yFtGBzLDrrWzJmoyZ1zQ29CJsaR
6Rm75owofWROjLvtVkSrFWhEZ4YAlPXyll/6JN8LsHe+sSQJZbe9GRUfZv/E
2qgDV6lIywkNypaZkDJzkFMI4EVykzitUNKkVgQWDcPeasRvB0aAtNzSfCM2
omDA+4HVq+BLjB8on4tyqXDa7dyyj1m3Fy8/I3R8S591episItUZ6+Gwil8s
FlDGCKC+QwtAV+JDuYXuX0sTa5eJXkPn/tRsJeNPRDe5f8T7qG1TdB5I5TNa
DFWE5Ffw2cA63h7HkJCUA8fgvJvxVRYEwDgY+FcuKwiE+1b21WQHvOVIG6PM
tY92MG+v9xq3NHiuqIuhMi11vD43nop+6XPVAhAWuocKEOkMVS/mRAl8EF8K
xt2kwGyR98rU2Gixe3ovaadlDZ4m9XoWRKG0jQv7eU1xaioL87xGgnDIM11B
Tg5B7wh6sGpkDoua+Bv+aeYFEn1qpeduzigb7wvAncUdwKLtIaiqumRFaqP3
GHGtbII74OXQyLC6suOODQAjJXOdUO7xrUoNo3v2Sj265Bczu/MewOnAQO7o
/X95xdGiEeSUbcsQeKFzafhbN5nw+NmC/XH6oWmVt90bNX3g2qrvGccXIssh
PJFRt9AKIsaZGH8SsqPGVc6iMANLrvsW1zieASRBKLNDlf5HPsZyeQNKVz8F
Dx8gLVHihzImC22tF9YHLXKBtMMT6DN8JgpgejUV+lAqWpgnVNV2Nl0oOC0R
a0uUq2un99eKjoZgJv7g2C4L5b0+31cIGsFIgNjfE8NT+TDuq/iEYB9a3++P
uYOervF6B1EVRK9Gt6Jf50YhRCdH3y3TzRVRydYqFbZWzSYMSewP4uGyXZlv
Vm2LPMuRatT4WtYBgtI/mWPMzUQe9/o/Uc5J4YkPVysHohBuAJ/0WP3ZOlUk
rWnOR1hmcxMTXvWtLs7p34KWVtMQryP8SXT3eo8y18QIRg3TubogVC5hucN0
YR6ZYLK2R3yR8A/LWSsOyUQ/xtKzjUX6hotqvDVMZNQYbfESJNAmgnSHLdZe
TkPiz4ondtkMzAHrCHK0ewOkTFE7VUngLkt88AtmAjAMXYSWZhlDLjTeE1DF
EJ1ZhI8Oevddb3V/bTwelLZWBYOITQv6gRt2nTl10dzzbmYPbuch9qpoIvQe
VlVQb8Ochf7+ovRSHClFgnjJSjhjjeSYGGNoWSoDNapkJpXFwlrS986A3/HQ
BpC9p2hXsVxm9CCQKI+fRWw7RcpivsDr1IgoTrAxxP+6pI1g+7IIgrbrPpqV
gdTAEFylQ9OxuTIXY6CtUY6ay3iqGBPtQsX+8JB96m6SrsUrJM3rf5rsRUpo
oZi0GnAwymBjfkE3jcJdVRLr77aKOfW6VdPuaXxvrXpD3Cj+T7dzcTU6q4e6
Ev9vkcE/p6F5OHV2ieP/wTHfd6zhI4ASCiSoyK5xdZZ2Qz1GHYORgaiLnEhe
s2wPt/pIy3vNlbF+rhbFm3qenHiLn12YGMfXVuPuVWzNNXZ2sWVOQ5NcPz+5
gq0ZyAb6wMej9uOAbguzyXKDIYolgBAe6o4XlOSTnNLXybyqDosc+ebiU2je
a1W8zSzLXiCe6Rob1WSz5CZlrtllqQe5MmF+Qpk4F+LWM4fILwgV9YlVA9RW
EgN7x3KXdCnl2f8mXEOwAmOa0Zgi+LkoGRdqcm7P1xeiz0TLFH/G4Jvfk14u
5goKaa5d3lixTSt7JtOce4aOTaFibM54AsHJ3YQIMmmyoIkEbUQ3XvStz+J5
8JAUhIfUh87YabnP+20FkTb9BBR53HLcmlbJskn4Dbtp/A/hZFCNuQ/IF8z9
WVo2Iz1rGa+WEGE4qCwkE7q8FXHAECfN8cg8zSCk8GV/1qNS+xmTX3OBPqp4
x95wq7vIVyMQUoM3XpmxQy170+2ZK240/2VCCngp0uLn2y0dlft+LucuFbx4
aoHMiROtyz9gaawztdsZj+ZZ1VTmqUwopRF27tkfB5HWaRYbvMckFSqfVjZv
C54hHC4iHhNi3KgG567gu59WgpUUeP3YKjqaTFQqvVu+kkcQF/atyLj5hKFh
8Z2rwHpCS6x54Bx8ddTV9ONGtItImvbaOuEKqaMuhAZ/JgXU10uZkV1HpF8/
xLac43Y15fDziGDqSaxrvp8GE8/1C/Q/gigXRZ1P6mfublqtosZucy3Uf4oP
LGc0T2Y3mmoE7v1GaAI/vQgeVP3HImCiK82Fp2QAqlCXFv6Y26reniQQXVJ9
d1I48hGRYXI9aqsAl4/pTdBw23ZekdxuUm3UeD3NvAjxsZLx3Tt0upsMLivv
B6oXee0LfjTcB0rFgQH8sfU9TZnb7il/uNakvdsOmKYP5daPmqyhhKyH5+Xl
902MHUNMrFo49bI1e7C5EawUpVd9ZixMdJMpVfk1+qg/9ug+IGhexXTJoM2f
M5dHINqraEJUr081gg+9V2Cn7J+6ZtfXxQN3ff/HvIGnZnEPu/uBcPHWeL1C
4UbP5T16FmRCs5PEWP4ZM8oDPvopsCKTD6Yv9QlnmXZRoxLZuOm6yACF8wvJ
s2HLg1lnp8mx2F3s6E0cCAAO/iW5Z7I42pSH+6aSdZ9EHUn5xEz3vUphAIKu
ajxQT0wenO+UE6ZrE7nakEWUBPsLBMIoTa/DOEu6uBNIrBqDJ6FRqqCxDPeD
P300385EkKG8yxnYfskrmTo4G99OdYG4IFa/cxnfBgX54npLFEA/8+RwKrft
9sQGd7ZScl0kzJVC2pNMGNXBsLSLNrBR1gtC1SIXo6UXGu0WaO5XtPYmHqZX
R9L0x+bRr/KKj6vDNyoxszIFxOoCt3+lcYOwrSQCH4iKG2y5xowk8+PR2KSK
H59ygTW3hHpxZEfaHt/ednr3+VNEeA/6qvJkcFgd6mciqS3e9ta2tUOFVMh9
avI5N2VXhD9N5zjuMwIgnnOAGX02ZyBVDYz97cbiWnAZoHiHzY5Q3dhErKam
TcMMFRTKHKlQtVZ4YoGlAxCzKlYHLj4oFZOziwJmrg+4J0D9wFSi5OIYWwBL
cofZr7i2gLQDz+/+o66ZApGr1VEYiChV0S8T9kDHMChGHuTfiOKsWjpttd53
qN0eKAZ/o39Is8nYDRdxqlJOOu/WVl2pMwOHtqPVwM9B4lcdp1vxULOIoZQe
95cSSb9gEF2OvTlHn3JRKu6lm+hVg3cLSLMoIxI+hEn1QmrXHyHS4gppsI3p
mqKOOEW5ZIOCGeUPMHO6QrEbAPQ92ji9omtBQ/VEIwB3hYw5ioADDsiV8+0F
nqMu9vbVvPArVmUl1pr9qAHRV5joQrJ+WlsaDdiAO8JZ1hdu76htU+LEEa02
hHhRYpczwVBRq3hUzy89825u5fiz94t9eNBS8r3RIjwtsEFf/zKWiGPICdMT
2h0WTw5d8I0I1XlOQjw2mL4wnJjHQml9jsYhywmxcIsUYEyY0XZy5ebTQQVs
lxVPXehUqq4cXawV2pukg8cHwcvxT5etp/IWq5OCS8RhsPdIYkn5ohZTXoSQ
teHkEiYn3xN+N+k8zIGBaABsOlgJTnDhCEDTtomg2VITd5Q3U5BD0Wy9A4Ju
KaIoB0CtIe3LEBIwiQBCvu0NGtN1WhIdcrCsi/4ks7QTD/VDutyuZXBxCl3C
tabxC2X//SVTb/csuNJi7D83d6vtfLlnKrDu4ar4eXzrC+tsLy+s5m2c1gD4
QTZhDcPR4m6pp597tvjt3idosuIDEQyh/gyY9NWAQePLOZPx2WqC2d8WpX5I
zmK81lJVeAv/sQNCcis3yzugYd42erZ20apTcvVDje3ASmsvP68GfS/MDinL
HUJZo7GcGbHTxs0UqT3LQlYk2ceLSFesjUHIy6A6fus1WO5eeMyvUhll3N5B
Cdzmf+eESCB2cqzNAhCvyXG3oL2YNlGgkraD3Udmt0M4s+ZjKzOGS/rlPBu5
Vd0iDsJ516AtiqBrkAP/JOD4ruhhuAUibjNplNOAYkjvFcJB8mITNN/dpiH5
PbadBQ0SFabqaOl6nkPkBcws4Zisns8FV/0bCKF9QDQ5P3lOIDJQp49NAsTv
eTX6OoRReroWSJM03i+4g3J4OBKjsyDgHwgZnbK7zG6UoM1sxHIyp5Yg7rZy
OkMr/GbqNWxGpdfGAnlb8WUrvAG+B2OXPAe1IhdWw8GZnwEYA5ZOm/nQwRZO
IG0iUuALiJfIwqS2apoYzXhuzU0cpgXjmyjHrRUQwhss5ueMfMVf6quispw8
l8NXe4R6p+7gKVR9K+KTTSppiosqzF9BMvYSb/6CCgW6RLUDheIXCGmlWGQd
iVFZBMzOcXAs1Wow0rm/Z1UTg8pHA/9UzYGPJH6S0KRIgycKRb798oPVvd3N
+aRU+aoGL/5UQDUt2PR+SMTfbdm2s8CGGUxUlSjO9y/gGPg2kgUKE296O8zy
TR2+VdTfRHnthY2YdbKp1G/5rxBdIbfSozn5XGcEZ6EjCLVvoyHRmKAwBLys
0OuoXGA9IxpQym9B8heqNHJXDf5RtcFvqi4Cpco6Q8T6osybiAVevmzkL5G8
NXTuFjV7clfsIWTuyZxK68/Bwk4tj+r3+rCmFMasssFk+O9C7fT65SqHgQnC
5uwIE+mxZIFHijLUKXxZUSWQL9SpOwPW1hO/M23N5HOVOSwCqPKfrAUXS9Jl
MKwVgFQk5e6NXiml2FG709zZHkzWcVVm8b9F2Oh8qELQ8rcR8781GX5WVcT4
OTgsbNdGdJ4v+R8tl/FMVj+gAJr2SozAVCdA1ulgjeQark9ul4NsTTSXhi0z
A90pbE6PmSYZZ3gXeyklPqGpRY3Oq1HHX+mNCE/CH5Ueqg8OuUHA1Zomplkf
gf7qWQzk8gqQ3hcvnpdD6F8/7c9w7gRRwj+8KnAj2YDxjEtG3V07unVLaev5
JWd0GRDCxJBBV96zHfn2SQYDvn5WET0N5+2VIhoSQRDKe2R7SAD+6fidRY/q
2E7ARdENOwDCd3qQ58+J7n1HhYiY2IWlI9myIrlS4lMsJYRhKUXRgYIDakCs
ljDUriXaNGz5ABl/lLtHDbOnraZw8bsgAJdP6/bMuYz4tjwqqiFQO28x0zo9
bwLqwULtLjpeUuWjtwsgEIRML8xLF+c9m5+t7FCk3dAfpzZavgnyW6pUL62P
cM8y54XO1TtxY6YDrcuwQPJx9c0S6MNYDGp9Z+JiESlAjI6U6IoE5U5JVBEV
muypfbJlHJfdtfRiv275gzwE1K6PKhak7rO5qSPpqtIh37w9+iqYmMyCBZwR
/pGG3cjJa64SwwpaIXejGazzf2IkrOqLP+l78NBOQhhll+9fHMLRgk9vbZ+4
+X4LbkElr1Tr0CzugMtuFUIE44ZZ5c4jgt0CzdlFWxz1hXejy6n8jOhtEafp
2Y//V0j//UBz/Dx9mfWUTYhHLaeAFezHdI3GDcj6sRJUjabyGDZi4eQhcG9f
O9lyuczVl2SfnID7947QrEZra3U631q9i6IrsXxbjiHI2rywDNkl8xz1F2cz
G3Wj6TB7p3M36hUS0y7bt6F1i45dWl12ZTAQBcmKW5QVc/e1KUwj9Uw2q9HT
LTWglqYjflJ6x6yjKp0plL3uqQ4/pUceZgLLLpfVPztn3Ncd3IoJb3xGnbYn
pSfFvXNyttQq42mAeQOlpANlsk6lKa7KDgpNFikm7Hts5C3xUmI3DlbA79aa
ZVMnTCE0yxqF4xo1CaTPyKhdDg64Yugzv5SHAT7ZeriebjxgRJttfVtp34XX
WAlN691R7TOIEisrwBywbm5OKs3kzdFSZPyz3Xa0RGwsHLM1I1HA2ERFwalD
gMP4qdHTsqel7sqtj6s5dgmbk4gHihHXZlgvpmAAMohvHIL1JqwFPaP/vO6b
3DCXjkN2pNiO+AWrVD7meA1PE3Wvvoz5jZcwmtEklQMWXbPurLJKf8CmK6aJ
42d11yrwQebBzT7l31//8pGCgzSIPPnmdcfsG59+i6gDkuK+VFW2utYYYb42
YIHPve/q9/FOtM0tFayeB0jcAKIitjpqnghVMOmJTlqSw5Nhgac54pR/Gp6x
S29HYxWmHRD1tTU2d0ZV2Aguh1zQcYPmy88xi9OGOqKPmxJYh3AnGTwrXAnq
0ViNKt4P8tqjCCN0bHfNCdsaHkob4VrCzQ/b9IMYsrjAEwOW/U1s/OdTPHHm
LASHMLUu/KDK3MGGHskbPFUwKH/IgFwauOMwnAppTGkrqlmEtKmDhCQUmizW
WS1ZAGcn0O/PKeCSEY800q+JTSdOwgkfyi/u4xh73JHVQj91zCRMngjHAIVC
NYSNGc+u0FE85lAIE/IZ6ybFIIZ3TaSjHJ7SmdzBZROW3+eRgy3fGM5ouGzP
xIXb5h9k+4/PvsUYO+Mil2pHApKoNAcr8jscrXWOT1R9BDgcclxeTo0odvDM
xWp59hg8Od1cr8ylC5FzjZ0DJ/AC1VQVR9wzaymzjWjI6Ehm8bVRIUiowEK7
djr/rYR3jeDU3niAMAGDiD1L/iBc2m04RfQs8pAUh2CYR1C5QdnM6MYQIhl2
2OqEoQQqWlxkoyIfjekj0vmPYkNy0KxpEexSwudTJoeSHLxGPRJAmHbE/C/C
Q6bfnmmfOdgLuhP94XQfxSl+OXlDjfI9bzgyY9i4aPyGRbZBTqk5YmkU5ZW1
4nIlGaMEo8LQum5BobohIG+G56fnvKJa9asenuc9gqFbhPp+Zyn4mETzyP/y
wzq+hp8ErHLb8NwLdJBvGyZdXU2i5oTQTvXNND4T887xsjyrNafe3ks/kbs6
Pli6jgMxtIjpvrJSRpMbo6NKIdVy7yXF1sZmHzCdM1/K7Pko8p8fYe1c1vkG
SEfiv3oT1J67O4avbdDvrpkPzEDZPXfbBvRm+sqK26gySEYzFLR6g2Wlpcnd
L1ssApUoDiNnhFJ9iUqYjv1bb2JU/4GFk3qtNnFV0lM2G8cdhaDP6o944hYk
naKEc3Jn2+4PPlm4B4PHehTmKQv6VhisbJgFOp6s8B+MjDVNxl36pcw6bb+/
vaYDM9CYiNy6Clg4+iWBtpjJXAnMZwCVvYFCQnDf6qgyxHbE5/wYosu3YMrO
wCDyMscFvYa+LHc5l811cp1Qm1aUjpSvxMkIoLbS3w5Kr2fGiMbd9CBpAZMH
q5jyp6gdnwpJhBrTbbYGkNNdS2CZDuA1XGHUu4kloaxORFm0GazCy0Xvn9ya
sQG2zy28/urEKsz2s8S9XY9W588YCQqlKfCwDKMFnEcREC3HRcBDudbkF+LC
dirTqYqb2YUlkxULtuXPrVi+AkodqynwgseBBI+SSyxs1NWtEPfrsui19DNP
uEozY8Gm4EYTNZLvQLH6ujpra/WjxsUlBv/Lhx6JQP89jhLXF7UKs68BGLH1
9RoDrN7U3gOSWc5ys/h6blT7Qwj+ch9Ixhv1OtKSggqsYZZOpfhwyWpNm2Ix
Poas6sBZ5wRPf2x6e0PSJ5CfAthcLoE4fHNTR9+VsC0+o7CfS4Rimm2j4juI
ZcNGDWSezwyLQLclZRUdqwd9QpCgBljwg/QZIimFmPN52wdi+JbRY9T8m8X/
3oWiIE7QPBPlbWanabTsnR9Ui3jNC6ImlP4ODEUbx29091OaZanX5I/GlPNT
aV/bck2RfkUfFzvSd82LHQb6Ek/2vVDp3zksChfzzRUHdXmKqq2YY8uWqk45
S281r/M4AIYuzNdRWMiuqnhf8e0KkVt/H/xX/uaHeY3jkp8u3BmOOojiQ9Hq
S5n9Tx+5S/vtZskh3XT8EqoyxPGtr7Z9ZM5k2CwNyVMGOloOC+I6K+5bCBoQ
sdsoZQz4KfS7hMAGcxVzNv3Hc6WoHzglf9in0gjr8i1DJpJ27Ud5j7n9Srn6
d6NrgAG1hlvg11yrVgcKLuC/Cmr7HRQvN715CZzgxT+lf0imP9Buy6iDnJwO
VhFZEyRk6XnsvdRT1xAa/nab3492oOQAfh7z5/Wv6pO29/aGjvcv5uFYeaoN
OPI43A7dUncZEYtVOkA2OBqAyw27jR4CJev2O3GPzFy/DZ8i+L5isYT40rCa
UON5DvXxx4LAtWjU93uCnBjQYeBgDByEZ4fgviffulNuXNioAtmDYVRfF+c2
4rVdTXVGMV7ciJA86rQkuSYq01OoPt/asooNvgzpHhsOMz1IENx54d7RT6ac
wRnXyy+FNhZAuRmSuc0SSuthgZrBNPHvs0siTrS7tNl1XXJl8r5LOc+jC9dL
l6L86hRQ+WIePkPPOPGryGXgHc4EVcrQcepClaTzhfa7Etp7F81IcTJDjAbZ
Jo3srJwJZI4HA99kjsmJSKSjSAirMNYmPdHzOQ+AXPt2tDayyFb4Tri8V7wT
QrJuovc9LIyPwYIgVNc+rQ9937snUuQNUHmgQqnlEVHfmxLsO/NbisRu5C5p
O1df25YEgY8E6xc3tBIRJuyV9qjM8cHWLnFLUel09t22cxXNW4Ry1J/axVln
EdOZ/C06SODsAZAU/Nry2d5Y0TTe7fKgTWZMViOzMdJhMQF55oLwUCuMxKQV
Uk2iBXFk2F38Aul9KkwIYbClHpBltXA88kla7R6nLmTDBB159yA/pGzcxTlm
qesS2MDP9I1JeEc42NtybTHiBxS7VhEbX8T4Eh4mnhATXD0DXwSIjoeki/4O
USl8x7F8ztJmEIgGifD7S8LHTArw9uy5uVt8EMHKxtsBPdpOkjJuBFMcbzG+
4BHoYtXQUjKwejw6hILidvtITL1S8V+eNa9Qzs7PUfuMsP1oyjaDtbNEOg47
zfssqPFC9O38e7FwbDi34vqoSMB+0y8qU8qnxpLecxn0SRBorFKVJbrx8Izd
8Qf6PLGD6/Fm83DJpqDGs62NfK4G/fYY+uBmXruh0LZM8PDrxiZdGXtqYJHW
HisPunN7+QfVQWmeZz5MSL4gPFC5lR1CpfQaehH73jEFUdZG5IXhht1mliac
5GW/JA31FcWJM0ZxQmH0/paz4dVnuF6lLY9Gmj2gOZQ9B3uLazvQJcNxrGQy
0s24Eeu4Wxx52Vu9aheKogXcaxC+fvbxHF3NW3CJAgKFFKDNAS26ELxO3oIQ
Pl0f/Zj6CuN4Y7S0uwD4Kq5ptbIikP8G9tA+f4irhsPiQLjFtQ/zurmknnDY
xygd6e6ChXtKjVrVpSkzp+nMvHab08mLuME85M+cizGKVjF4J9aDcScXykRy
o7y247OtCydah7YI/oyo2QsSHcHHcuR8GIxGqxVp6QP9GLP62Fup6h/rSlfH
EAZrLMCQ9yhs62Y7FvT+Ye9xKpfYOIwDsKIErxX2HWK+wzkZRp0xZarY+167
5uQwrMcw9ZHP2GACprYOAcZ4sFiWAsc7KrkVw3GfKHiz6Q+MgXHZZPkcLsT1
fbyXj9g7lDo393XopW+MT6382jO8DrBD4nWIbW4qa9q/o4DeAei71afyiPjK
IvGimbs9fJeljc3QPbmQP0SLeC0+C9ExpVYt9gFoSZjnpa4bfRROCwC7O6lB
48EvL60Ps4ga3XC+W4ByBOTUBQb4ZO4cuPUstDhbhIF1YDREfoVASrAGeqrz
Gxh1NHGfDtV3h2oZ/HR3bFKdcZlZM8kAeFRkCTI54BviarJmbIfZksM3EWkW
TwSlfMrvGByxUmDlgali3XbNRy7qoTlwNXhcc/eWJEBOeDha0KmoXHAH1rqN
EQgqtSo1mjZ3y3FHHi14TO7K6zUanNKQ1J9H1yVsqG5x042WW65H6Z17utFx
bkByHJvowc2bOVYzo2ahRE8BeU01mL2vjWOqPV+R/iu8VWFNT/ekaFSkY6nX
QAlYkYw0oiD0M8feH8GADrGBiGMkpQ2qRMhV8WyGBneB+nDGJ48PLLnoZZGi
WL3khuaxo059x205wn6KSv7K/DJjyroUo/LHeaW4zrS3XF3ql07OMtUC3UTk
d+UIZukV3Y14F7G8XvuvWCpYBWeGrLYJYiG0p5/aYvO5ZOZ9EYFP+8GHxxBj
l4yZib8Mnsv8VWkLt4M5aKm6RLmzL3l0AvjTBEowZbdzMRw7qWS3n78WRwgg
WRc+LYM/T1rxoOW8+/gD+QjxmFj/MKmnlrtHa6g+5bGvwdLQBlW0sYnSPfFz
pzZBXuuzo5F54hlh/MEIKrvmAQbcr9y0X9oy5Zd6bw8Z9Qi4nZvoUNN7zgFJ
FsMwa0TTw2GLVmsyIvAPnDpn61WmfYgsBYBzBM1HR6ntqSeGpBYSvBQIAxe9
G8L5pcq/FbQ8PdLEj0A1NUgfft/T2qqGLm/mbCbAYNA/LOk/flqYU62e6iL/
/Phu2prx3CX8x5aRBmiZeCmgTn4LsrQj4o1l4ugDnuTe0VMkC+zv9DBmB9m2
ZwXMGREZXIOmzMr3EIV77C18QeNhi7ZvnJj2632jdE1EL0+sXcNPV30DwDXN
y0fWzAuVkNAuwOUnHwSL8+H1WwwcfyH056w1z0cKV9cTn20SIOw628UiYsg5
NqfQHQDu52o0Qbip12XfwKXVGPT6ZQIyXvopMSYGM5MGR/cFWICfDjWziyRl
t+pKg9wQWgaTkAFLKWt3OOK8J8oCjQtMYEHa5rA7I23xpm9ALcilT9qM8xp0
sti/fR5eo+elBykmIESgzX4/EW0npkz4aG4qDiwHdhcVH0AhzkRc5nrGAYSj
2m6jv1gra1VB3lexjbeWzejfD1HKKPTHptN8NKmCbu4XplPaHUyOxoCXwvVN
vMQeV5Ubdy6+cjjEmaY5jF8WVPW0D4LK5qkb/coYabTtR/qmVI8Xd+uBJ8lw
NFAvqljFXFkjkapdjd/iNvIl7KrvRNSDzbAfashgPqWU4Mnua1GxRnrsTA+w
GwdO0JUqUVXolCuBYBGLMHmLsld6jbwR9bwQYlI0y/xnoUonxMHaXUaQAiLX
hM3uhLkBeRwlrI8nSxPq7VgeAH/mAXkocz+EdpEiM2kx1QuDkrWVI+k4YXP9
mUfKZUnCTgOZ8jMXhC9mr3gCTq3W+wCe9p1xZpBn6UuoQdn7/Q4kerJJwxm9
VVNtI/mz5vifzKQUIjrCFKyWq+AJQY7w/ue+JuYPRR0mZQ9Lqz2tW1lKeo5z
t+PV53XzxiW8W5JfE2K5vG4DbSmdE1qmO10n7w6WjheFtUhwPHaU9rD3g4eR
D6HGkG/GhYYQBHsCpe0UfmkYy8QLyK7t2x9+VJDsn/xEEFM2Pdv5r1NhEYhr
rYJXcM39Ql0hAFA1pIYy+rB9A9wTPAmtmFzrO54c2KFBaZxEHb5j2O+Fqoif
W1ZHpPTD6B8kncJDSkUWzNzI5RpQr5YrcCGkQvqdPlW/foMEIjvlqBgx7y9F
0Wlx93JnMu6kG7+1E9Cb5YJluV3Tl2knzvOJZRJ/mHqD9Y+ngxOYFIpKPYnD
ogI+Ct8+kDpxTUtt7owOsy2S7g2qAUE8pAEcGtQGvFPOxDvNEcArWx+ZevO+
48v87wSDl1PS1UoPmfKgijh2dWTB/GeYCSr6eovOKAoQYo1vjVYzsuJr6LU0
FSDfqlsnq2umAnrcMRTbvr8nSYEBiqqQggqV3NlWq0kf03mo5CrfRkm4aEUH
A6cG5OxyqcV4uAUzXQ6lqBh9WUCfP6yG2+Ncwx2LdpZRMeGV4m49so4z/Ijy
8hEL6pC5nhpnjSLv9CFBMGKue8Tfo25aOhMgssYWrA+sqgywTuekZs4fec5f
k3w9CTYYs5oPsLMgwm+TjYTY5KewIrcMzPOv+w3SIp8PEEo7KN0eoU1lJF+r
V6SE1vKBtrrWDCVVx4/F+6msPPMF4FVTLwFiV9ssifuDOOKcISZHIxZ8g1qY
+CU98QaXs7DGlmOS+1+UQWmYk1bdNHzs23HhgqqVXNN4aH01cVmdYIxcCApP
jDYFgUZUyxl/tzpisUFGf2biDA4vArPTbkrhPVeCtOrusNS7fEGAPqyxcFNB
XZSVsziwY9DXVSkRyl06/nFdsEbLcGoKf3m8jt7aDSMbdtU1CEnUrAymsnJG
kYJsBgUW8k2ZMpOgF1dOl0lW4Tt7xgDPdwliNtbg4CxGz+6f0Pd83/1RmIED
u6Z3Rx01rEe4Nf28hVySnfT4mU++GQ+ca+Rj8RXJuJdj3lWXsAUHVMO0Otuk
jproTzxYB3gjBgqS1g5v/KNMCD9QDEAy41Or6wUbjlXsivN4nF0IPj0s3M0p
m5hp4GmDo0RslT+UcFOTsvZE9Kqgj1RU/KkDg2YMwjynN+g+WNiroYxjZ4mt
KMJQ3b5nVzSVhNy3iUwddn2wPyaJU9wF07SEbTM+tMHIzxt7/mH37Dqsn6oI
ds8/p7FxRxKtiCk6YCspyNR0dMCs//0YcJo7QvaTG/TK3eIGySrRjAGhVjc5
WHFfF4O54RnVxpOR0DpZxklk5aGEGsxEPCunNe/FruZK/5j/y3f7Kr0gv/v2
XbZb3NzBQaLJ2irdtHvwoNchHEAfKvwkcxglUcPkA6jZUzo91dkbmhkX9cAp
SLKoD9BmieLjXy1gQxRa4dYVFfEfKOpFnXs3aOSPLrxVRW51CQ5w4IViqkTV
hi707n9a7Ajv6SoKiAh3jv1KqBuPiUTyaYq0pQNy6Vlf2z3N33aSQgO2WpUL
lb/uhIUT5Di2OZV9Xwom1uHTZhF/ykitJGlXoTpQ9cJX3kFqFuOjDSROscMn
qhXGn0gErl/foV5gSEnSrSbPgV5+O+j9w425/LZpSZeduJktAedWwXDGlC5T
+o94vr3fBOk9E78SICCEQNRW3Cywm6+JJ/bmsnthKutFlBP6qGVTuq2mRyN8
lsD6zFlNo94ZjtwYUSVLfKV2+J53Y13kDG6S2PLgajvPavsnx/KBcdev9UBx
+0BzaKa77TMKe7WeWpaRj8UvTBdOJn+75IeN3se13v1dqG6tSdRzDmzBP5fH
4tY+FWrPQBNrvY7WM6Til5XNN7011w/8iiPXFqfTY34kfJwwV31g4OhtpAgt
U4vAsSohxcyCcqYcbBSec6+3vgJdYf64P9vWQ2njUrvU1b2BgNQEJwcMG8Rm
bzoNSy/fUa2FszYAjfKWdUeKeNrifsw9vukLXoNYbyfY6RayggYYtwkNy0J6
fr1z8322b4yvqh+ns9IYHnI6bGx6xGQZdkM4/XbffmALi7iiK0YTM4hJyW8w
aWdJ7B9ZtF9tlR3JW/R4PhficBnvY8kY0zHldm38eZX+bK/7/dLJLSww5Eu7
+/PlhLJAdMSqE8oX7Md58zRKsYxdb0rBnSEig+2EemBGWTUt9XtagU1OLp8I
4m250i+l3GUM3cP6PfsxRIymmRfD/Oyee7eTwFmCX9kbBYwR9/qX0QDT8VCB
x9saDoLCaHBUE97iGGhyCKD5Aw4g9BpkrnpggXp0uCx/nfc5yVPw5ObN5csY
TDpcHh3aESyfpOSI/4/yJoGlL/ripzvTf1/1qlXTxMQNXoILQifhO68d+P9O
CElSGsBe9LDl11h/+0d6n788O9jhgWx48O9vtT347+uALfqwRyhKlzD3Wpj5
Q/2p0pclHAau5QyjkjboL5S2V3lqQMFfg7j1rl0sAbjDqJl7+q2PASMH+FP8
n8TLQ3pjXnbq2s4BVqU2XxRdmGDP4J+0PSys1ipDmhwFCa5Yc96XQiNYXImM
iOFA9+YDm2Pkuindlwg1j2+n7v9fIGPEcPPKaBjDuZ0z4OMK92YWAiMmsep3
KveTX7WUp2cNSEupMVkgQ25dU691ZfP28Im5SD0Bu7VBNyK7p/IUkaduJskW
eaeM5JAyOb72w9s5RDGumSFZyQr+qg4qUoWaiIiOr3C5d3ZYN8hsKVLi+MlE
IuBaxM/fTKZfhRXFxWPnsWKc/0wkre2M7NJ+PyyLd2UHH4My6G4WuXTZTd+4
t731PQLMR2y6Na4kte+y3eeNGBptfiHGHi7K887RwXhoR+XChisP/2I2dRfF
weLH0PGKQGhgCWEH4X/CF57XLBcAeHlgV5rRhZKcZJR9D7vn9PnGuNVyDqup
eGtbIooHwq0AqzF6CVM3ugnlwh3xz7iZz+bu42+7TwON1KPkZ+TInoPFMMic
OVP3cUEYjxRTv+ACn7jY8XI+fR0wZ7MTcgJHCQUyyLn6dibWnjcwRUbsFPgY
qGsrkpg8Vwbp8oTMVkG0jRg2bhpMGG/Q22O7k8zt/EXHtlIsdY3GHdssss0w
GLQ7kC5eGJymC8azwqzJnhNcJdCK+liefwbm5kRvo8IDqmLNmnOc/QwG4wDa
3Q/V2+wiJRC1qxkUqpoLd24ZMyzA3L/uut/EVEp/i/xMESgU1d2nZROWmc1K
tIeF/6NoYt4GaBz6oO2+DtwsU/eYzDocqDaumk+H2411KMi37GakP18WkxP0
8p1dkndRRAen53rVqN0W6JnuWT6dcUT42ZCaqIvPqYnEMRA42Y+9vVP2u8JU
KDTnSF10+wA1RVEckz7+cvJ1vbZL8yjEMs3lhBLi3RBPwQJkyXD4sd63Pguk
pr+puzKUtGpFLVMZ0PfMqUTvThoy5OOC/s96reMqmYmvj96JGYitAEvm06Nb
d/NPXokjluwyZVvTTSE38jlU+K7bsMwJ5vZgOkn18weO3a8d5kCSkTODIrwi
v2knJGjX8j8knuuX06czTRACC/EFsWP/tVPOcrGYRONGxHy6Mpm1jeIvxNo/
DHoKPVIM75+0AnIU4xK0qJfFDtCqd0LNVivn8EfmuGxlQM7qhnjSD5QvcKpr
bt81yGFnNmEWsImRydKzikQ/oHfvd+xStT1qoI/GX+9p+yhtuuMvcftnATK9
caCjzkHreCNqUHvnanQiT2nUXFx7SIeVhnwAnY0MH1YhzX8s1w2DoqVZNpm+
N/Qyudx0NsHSDGigjncmmaXeTHMJYH6m1DJxOCIj1z2kbJjZe6b/wT3S+Nw8
ARcwE/QOu+vSCZeqVyQGtv6bgy1HpYcRFwCsG6jY01cOxfPVVOL/XiDZyZiU
S6kwB+VmP+d9Kl/xBrrx+IU0dSalZdpwt8ms+QFXZEa35fmrEknY9mUB6cOT
V3n/uUmcl8ZrDJ1lZrK6zGfyNSCYxjQfCr26beLkT+nihXRO0dAh6+0foFGo
VYr2hbCmrco23iurAND9DttmNz84ULOqXIpiC59VLzDuKCtHHZSHYrh5D4GC
Zf5iSFF4aipV2yajBoXH6lIWO56Phn1qmQNrntIEVgvHs+AvgOxrcrrzE+7F
5kgpZlPcZbqb9sbdxgtZTDXvLrTsWMJ/J/bUxFwSOKGsppWSXmeYvcTlkl5h
eWt9trs9xFkVlN/Jyp9Zxm9I4d0/ixnIjyWhp1rZj3uB9QISHHFxWIaB7jOJ
JQuH0s94ART/Shmaq94dVi3R82a6GFD90iMHqDyd5hCtrSq4y0ZUd5NYhsC+
EobqVVQmSgVC0f+ZbZ2BU960b7eIKzsTWjtTWcg8imTT4G8rIFFth6UNLu7Y
A5RrHkzOGdUxnMeEC1CvReAAiQzElKBFXQHJyPw4FcCgdbBozgaXPt9oQF8p
7KjwXDfwATkUBz7G6p9kOhsHlLGLKwWnDSiHFOtKo+3D/DepMKhqVvKY4Gzl
gTgfeQeVPsWz4sFh1kXeqQMi/X6FR1Ipz5KB41v6+qEFd69OfApllx/TEALD
q4sZ9VSn/wFmm/4l7MXHXQB25Wy2krCKS3BBbP0WoTKkW24Rckn5ahURLL/Y
fcKD85hkfgmxT8lOeqw4Fg2M8xQm+rzVQ30peJfbsisA/B9z7hi4gzycPEgl
eODZ/4BeksMLFi9Z/hKN5oAByvL0Flw0KIWKwt5WnbkPWVQ0BegOviyrilUk
gvLdT8taVN9zZw0jb6ewjzrwEqzVwvzsny0MjB38u6FCXbRw4xkh0i9L4krj
ekTK76H7pghYWk/KFRJzBnZZQ9P4prBvY5FE3GmC9QypAw0LLXByMvLcs1p6
MoQetSOMJFbkoozgv6xpae5LZwUiRs1dpakr2v9IT+DXNGDUUepkyhLEAR7A
NVY4/0ff1NySb71M7V4xFm21HpuF3onbGTSuihLaNPkhBk1h/xU8Ek6xf2tE
N3FqDPSQjsA4PWQQb9suQQhWSDF6fFX8vbDLb5Ise8OxImnK2OV7/IU2vVvx
KMDIVqmlSF0hGbTkFt89NCLT8644n0YhU6O9zrIw0OG+gy2AcxTSgqkeoddt
pJ4afgvyrt0JShR5FJ35RbcAwc/09JpMdolHfXyOhnj6MfkdWr76lJMB9707
zu6AnWcPLD+NHQcJP7JSd8OV8fwlonmxbQ+b0RlsWW7TEc6JMSfrX03Pxd5L
mvibhBHYuJ5Ezfp32pyT757TNEKGagVBAhqTewVW0V2HU8sDPXi7/x5XgGvG
nUU5MDwVogibYrcakaHtM2wOWRVLt9PclEzI6y4JSqnx0YRI0s+vvbSZDgnL
sXmbLDvimNX2FbEDJOE7Vja/4TYFcrxIBK2m1c2rtBNOf83+sqeKD2qiIXTF
TNCILb/pOlfVIZE2vkCb/KJ6UI1Ao6nHKWnuTFFOv5d4g/UyU/QxsT6U6dnb
hCln+fj9FlwZlNksabYt8zgzesctCcUpS3Kx8u7YAIzqZVMKbYkGEFtsFqF/
gARdpAQ9xYdwn7vUnuKyCX9yNbGtnaGBEq6TOePLLlMwVs9XdFjujXc6C8mV
S+X1yZSd4LmcCb48iKW1tHz864mKDFgaBmMU2+Bsxv9pK04suY5xfK7t230u
fNpM7MZviT0sOyxWONPvItGMH5uY8tOB8OJ51fuSV71qYy9KteyMizYXxVWG
TUi16893T5HxHEm+2fbpPZx097FqFkT/PIyZpL533RaC5liXJIXTj+hKgbJs
sIRYHYhyXU71QgAHsnoo6m0xI/oXal/AKRuZLe7mvwMmLsuJ7eWg7SzKIraj
CINgPL0NeK1wxf3FKwCKFjt5h+k40n7NFC4by/uZk9MT2mtdSIeXzsormjZN
GRIEYNokdsosh2FDNIM0lIf6GjSdLG5BJ1doGNlE+d7JfQjdzwsGFCd+lXsG
8uAw+eF9flqNIz41M6osu8r4/F3vTxCgNyL33OfZYXh45pF5Vq4ETvFPw8VY
1kYmolclbPqb7sPhwOtadT6dncWbQWp+ATYETvoVCZqTIhBaNGWRqlZGoHOr
ULmVBmOdVpK1saX/nn2oonatqdFmcA9Ij12eEWK4Y/wcwJAbA+H32gcZ6m9r
RDJGI1r6mxHz69wOommagNeOl8oNYsw+XzO05L61Ee86I6G1Jxq1H2cjFEJI
UmPnSEESl77xPCnl645zHwFsl8Ozkc4gtg7eMVfsYTrYCk8nft2wAmI89OMs
N8V9snV7CX0M5wxKG6btfkEaMnZtDYb5E7SBRktXI/5Ms2CMxTB7sMqSK0T7
cUOSS4PLEAKNH4TJu/6xSnnQbmJQ8b+ASc0+Ad4ZVSq1s2CF7E8J+Lai+yYa
C8oPtK5F9Mnqj4ODlIOnaB/Hz1CPBoD3wSw5kRumeoUNS7xUpWRw7xE0KvmO
1Cvtjv4LFwwXqAqt32SLlRn5qU0Lnbqg7egoopqFLkYorJLSMxjwXowPOqmm
YAlXVdE+Tj9qQsNwAtrdWzz2sHsuiuc2KMCxCzz73o/uW3b0CThs0qP3GI50
lSrlJ/7YfPIkyuElFKFy+bKsAMEMDwxq3RJg6uGB1eNsJ5MzLL8cJdNX8Fgy
0z5ENj8JBIyGu1MUeeazsuPvXnh+oeS6375URX7AOpXB/DKPJ0bduMW5IBph
F2VpKco6dyLlboUByblDlWVnIeg9NQpiMNOGQIzeOpzmGqCVHwiqXIpu7TMy
SmZFwqK0GWiobU6LkdTy3okHUY0tY229WUWh+SP/K6AHsmYAQLUCcgKXBx0/
VFPMv6cW+Czal1CwhG3jMHeYZ7+e+wt++3ujgtv0qq28v1IJNZvKDWnDSU2t
3VA+d+S04a1/NKtyYTPH2MTEfNwP6/7lAe8orChuI9feTTNazxZr/7iaXt82
9OOy3lR18sKgsxC8QpxdkVpaDeWcN3cvFgRfTKkSPsIjb9HjWUh88dlKeZDa
UN1y5loy/zgxCLI4GCcLvU/Vueo7hoGOeUeelvex5D1XdH0F8j/+iOo+6xiA
KO9pIOwJnGmBjCUqxckJB7PvLYxYYv1ZJge9DpychdkhVoFZNx4S4lGrqb/X
71zSbLGEbaJoNW4TGIclrKvwSyIX6I6QbQJOQHVWrqr2n0nVHCUDa4Q0+tU3
olcbEkh+j8ZSgHzNr1MIsVbprVxYP0aPOsUNbX8ekXIhL6MVg9JeHVGX0LuT
9jETDotDkxjg/OLsdURMF0xjH4QliCONhxXs0eR0bxYEzs19MhMSVrwrzf4F
/td61LC1RJMgbyiMHl6vvwzaWItWrYihMeRqSS2b3HOTamG3u0nHm+am3O/A
5pVgaXPH8ijYBeAe+UTfT+2leTZAk3B8WCapNAV/h5jJm9VFSglaDhDQu/ew
mIkwOh3duui8SjLhnMdOJrArCaVOgGmTxYjMf9HXK/eBVphkmf3HrYy36LpT
r2Gtgc2BL0uqdqVUx2xBN8BpsAsayRHYAQFKEtWFNOXajLQOvoRxvfL2BZXK
7nXclF0s88zkotX9c/gyPdoPbeOeosQpaOCZPcmT880bo0AkNxmTj/jHd3ht
/KXVcJGh59G3liI44O7OKcV0Ojsm1navyg7A4sywbC0rkrhQVV1+EGNDjiFe
S9W2DzSj/MB2IOrHmRVhzBxTZGHK66MDu3TrrYsCBJ4ErMzt8/IvlDk5eNiZ
SGanrAPqxYDN9FpST8p9rWVpgnJpMwqLLKHHOuzaw2Z8qjlL8+2RmUwdjnfj
bGoszcKV/5sJL3nBIz5+WCkr2SfP/5Old1k3OQagTWOBA5g1XnA926RVaSsH
xnQXPpw3tvlg3oiEJIbhfr69vbC8xtmXKhldALNl0T4h+nDBk6IKRPvVdAy8
rL43/Ucy92ER6Ic8c+II7G3XrBr8mtG77wT8Qksygt4hxjEGTccF0edthNK7
ZwJ4LEWFTyHEGj6aQoyesqu/W1QC2UN7B1QtY5VxlRQxdzt2EXd0Hacb/TUE
Of79o8TuOrLcy7hhfcyoW02tTWNC28Ab757JefzqGlyF6MT7DE6yedCAW51Z
wyROIjvOORnr5aAJ3Jt0i70Fw2CWVPFCbdUlMlhcqP/DYm6adSszDenB8I7o
P6flVeGuJ0zoqDNJ/mctPv7Ebed/6e+/Nw75xzOoj0WXeSkV4fii3jnGGm/3
JqlUzLi2Q0hrAe9HyqJ5yCQo1/156p51EuVyJdLs44ffS6uDRj9Z8akY5VKX
4B5qrRuJtGouAY56YWZlO5XXdHx8/L286b+JzJFrHq2+WvAebWlJkZQ+sg8U
n8PCwbZcR6aXpReRw4JINsFjP7h+zDeMDFkILRIv5qXQXPHsuqA1jlOzFuOY
u50qCdg0IZnb7Fu1+QATcHQNUoNhU+p3hSmHf0S6xnOjVoCqm4cvq0X4Lrep
iHkSMZq4cHc3+K1t+nGtOjfGxyossX6yb8G635VErmbpcdLY2QNdWU33zv/E
ZkJrYgf+CHHJFaIrpb3d84M0iDBf9tAWj5UB0g76FP67OVK4vTv5PfWq2RLS
vthowGpW+xEfR4Ke2aT6rNDnB/X1/TGbcLWltuMadoQzNv58hAVKfl9dbJsc
2yB8kSPRjvyectc4QugzTVRQgdcH3G1X/Dv+WiT5hU1ufoe1E7KBzLBY5F2N
wtCSy4YnqfUHEDCJR2C2CPMAgctygRDvumBkFGqOWffL1nELCTgKugTcJ7IW
I5bOylqPvHgS9Q7VqY4toq/Yj/DFsswA0/ZuGrAtWCIrKu7HRtQcSTZvyJTs
psgCfjmERXrY+27xhCTP7xpgEwiMCGZ8YkPZcTreSvnxQRG3RsO5KOUaDFoq
4J4JgfQiSTgcl7LfN/roC9XQqVcktC3xtN/nJTnAVOUVLEOpWhQd/DIVfeYd
onuIKG6pe5Mh64rc/kqOV1REJGKThabtrS8J8ma7xkbZ/k5JogOQazrjA9Hq
G6H74cBL+gYwrJa/j008PTs8eCFNjVUSV4UO2i7GsG4chdSU1RHTOrxTG6YT
JR6Toedw6OieEzl+Zm6dlj+zqkAW91sOxXeOk6Z063Wttdl5lrdKe2Hq/b9X
BJsag0Qi5jjexI9Gq/MHt/g386WiRXWrT4vbhgUV2NP6OOU+vxZDjpuBEbQH
iWQlU2FCD/XcyGoqeBhL9LbgR6u9eLdBWy2ChJft+6hKDmsg6vaICjXXXCHv
FTus4hElI42TmgZYngJ9XTPA8MW+7+yMIjqzwFhUo3ZL+ftNvNGEl1QF0yjv
qsq4OFcEoKOQnQXJwPLKLpi8m/XaWs6z1dn2rErhFVciVHtRU4RVd6Nslyvm
tkIbdVz/w8jU/iUDY+KpUJF6uBNIVlLzlrmkEI5OBr9AL0GH1kJrjHF+GzOT
oiK1+rAuDjCa7UvnoI18zluGv6EckMFptLqaMfrk2mIYl1sKoDAUKzuxDSe7
uBDEEEO3WQyfH92c1mK6YaZzx3bdnf4iqaa4TrUVFoGTgXTY0hQ6Yrs/hQwn
XKYYTNj9+ojiigySYJ9++LuMdpHnXeSnKD6nwv6BikcG6gPyyKMy9E8/LbVV
uFA+bdoGnsmvtxAkMJQF1hj8Hz09gU+iFRY7DZ+4p9z3/VWVLErJwYdq8y/J
MwpTIK85qIN8f41o5nEnbkY4f0a0zykDMhTo42eMjNK3XfmnmjgvHT260iVT
5Kbtr8bLrj+IvrFkKfO2kottLNYk7T+YIqJ324eW+1UxD9AGooUZzMnyQYg4
qr/TJmMw8jFVJIe0ah2QwYDitzYq3lbLNnHvjkmVodhiqkNbG6rDadBbsT9L
cNSksv+k7sMR5WWFNNk+FgZld4KvT4lREOtPCQcqkCXUNaFI+qMOP6W5yPBt
fFo5jg76NM4lSOPbrEycbt9rdfS3jj7FURY8YZy01CQChnI7OKXMUBBjJQIC
Bj+8aK5U5V2KwKfXDXZrCl1FCUyLQOID+ztyJeeewvPuTRq9lVEenZ2IhveT
WfIIhfH/P2ltvWPxK4afAWnbKkCQCcHcrAbwLDX0TtMqGuJOAjsxOkczdW2B
vZ5rQT15SGRi0Q7+QyoJaqcSguHhc6HEUlb0p40BsyOkSsCuFksAQo8WHFzJ
a3uqOSOUK5DF5zud6gspaLjfPrtPg7KhL0EqBuz1aCpKcRG1h8Squ5JQYtF8
Ycy8ee7RSChK3Ew4jTKDpz5Y1sp7eML0hrgbbDlzUI0A6Ioo+NZO7ueHedP6
epREfZHfNCqmnpubqc4nKBC8SrixO63XYQd3TzYK5vYFYTXCpm3Fh00nXcSf
bAxBkc0WS8b1950lTZgYwKruRxJrc2s3ZEtuTkpJ6CvnGTWCHrAa4EZ4kSvu
dfEaQurA67Ww9Rl38b1RJLmg5Oro4bNAG0qMWEh6bv8Zmz+gcavbeU3E4Nrw
OTDKCSq9RADRacoTjxkHwGgaJQQ005qgVvOTQJPXtxeVw7D8YdjbdqsX/wQY
ik2gPnmwyBun+hXKgOy2SHdL249M02WO2K8aEXs5t1m0CYRhkExjVn3Cbo3+
Seqwyhto+71/XVR3Yv0D79DxzftIcm85ZQ2ImUYTf6oz6YRRto3ZEjKn34DU
iCELnPsFl2cemj0WsCYfcF0YU4106f1AXFF6hoo2OMspzXj632AWYflyjRoF
IOMYLTKexhC6nvIfStm5iG0E93K1ztbPbT5xnNo8EUW8T+kpevrZ2TnMMfct
tia9gLg2KfL8clc/ZvOHJz2u1cIleie7Ix0bDTExT2f5sIneWQ9I2W1CcY9Z
Sc6Tni0RiTlpKXbYN213Ul5BsFeP0GeO8jAxaajyDpgXjSWMmiBSvgGGpoE7
MI9Z4h3VqsJMPSIcwtrpcL/29lCiuc/dCEtcpy0KrmqS27wVHOUmpBUywtJF
V2Jlbe1Yx6MZx9+z5AN0qd4Y2/Hu4Bat7dNh69Cqtwy+RQLVR4KmA+Yh9Htu
xQXVCJc7AakoPqv3DXiSOFlPdvTQ7kp58ejC3ZQdfSKBbbMjfEY3B8KdmH1Y
vBAaz5KBbqEH0y60nyMlEsjlhV9SLQQ+JnMr79y84wlv4BTrzHu7NgfW53bP
uq1NLgZMg+vkjKndQPrj7FIZ7INaW4zDWof6cE0GlJz+xaI21SZBPozs2D2C
TsrL7EYEz9chJ+pHNNEh+9YSD/jVBv+KiKBwD9pfuYb3ZdauXNbGE4tlHKF5
bWI79h2VVWy80h9KQXEahcffvOvFoQsJg1+vqvtB/vVVplVphZTpZaiUuCs1
u923y604wCmYhGbYBjKczBYVTM33fdXP35RC/qbw2OqOtAd0aHwpL8b07CAG
vXozCZxgAviVUGA1eSe5N28G1IAUe47JT4TZBcoiy5xit3vz+3GDKTctVb5C
oj3T+LRLog0oa17ns3vNt5RaLEb8IieLG+UdoaLIb4ErpTaRL+3W3WGNRXf7
8m2uhDNuTHl5bynHWCD8G+20QlWCFEcn2QU+H1ktcZ83LE1/fMccIQEc13hU
S6riEUACPH5Wz5XD8iaLPSa0PbO/86ID4s9Q1d+1MNEo3FBYiyv8Dg62IoHH
lREFVgsxaz86IMemNFZc8K1IDIpygRzjq3nILHYuH8Ae5K6y5Hex94x7ylPh
lq7hdzHKK+8lk9AmU4Y7m9w8yL9m/n5RogHWlWCmyAENB1F1B/WLI3nFumgk
k57Ikm087k3mliqM+a+3CvUwwFRAqZ+EgBiAYIX22EXvS1KlGU9ubT0C67sA
icDst8xZsVJ2uyYfLIKo8qixT59rrcSDace5L2P2zT0Yqw4oDbZLn8ifCvSN
2BjcjPhqIQTRb+q42rL+jesQgjS35ohYzs7N4Pdj94k8+ZCv2zErGUJmAhFb
h4AOjdzTE7AQYO4kBxyf4mcHEnlMH0gU3CGLNu/+TW9luFzLH2wBgTThOTtP
+hhNthDRqCRZcwofFgtI98VdhsVeEqOKHLUwFPLafyPYsgSVIVYRwD4jdV3u
VjSieiLN88jjT7/TdCQmg8ELSTyCDxcOOowutIYAV8DwUe06q9Y8Cy101Exn
A7YkSyOJ/omj8fX8gWz8CvgVnIsb35pXQ1E+xmoU6Yg1sRXDbpWPi1cMFwYD
UJ1p0dV1GBDkY+pvml+DE/EXKmaaqWN16NoFg1g1EfkJe22njgmhJQ6Vn+8k
9APadIJJAgaRX3r3UaDgvfdQQMQDp3cjSnGoOo1MYypS+GNtG1+jD2nUhfv3
hZ0JYX3NL7uYJuDbItu4FiZJKwVFyh8aGP4i7o69Y+PJUI7ekYPGESRYtRK8
zZUGLH23/+lSMw4BmeBBa9HSJ+TvkKMnjj+dnWmrpuiw3Yx7LIlW9QP5BgOc
lb6mERoF8uuY/vVYJJZBa/cS61P6lExaSJwGI+K0hxTaI3kU7MC8WGm53ayC
MN31mn01DJQneiCB1z+tom+7dOWy0TTNaQ88LOOnutZJ9Sh+pT4a7QPzK/Ra
rfCUtC0mDmgntt+C+dCA97iueoWCgfecQ6avPYXTa7iTleIszkJhiCMnNNtS
yp67W1Kt/uK2UOi178cMyKq8vDMd/hRzZgJpvGUiZH0ZKtdNlCfwJiWaHXJ3
ut9C7Mm901FG+wPtG7O4Va+23H4J/nXXhxAa3pPTTfI82gDGxQJ8gKNCqzYJ
zGoEoYIU6FNW1Dg+y4MJXuixHrC6dK6KIrUmg1m0fwkE7bcov2MVrpb9RsxM
ZUTm9U3nZiVTlzh531b6amj2z/2/tJoxoaNPmS0zVb0t8Lf9zYRgrF00h+iU
9mFLzwdatqyO/2+lTnD6xq4lcotJ3Haj8PP7hVOfMTPQkAvO1Z0rDWJbHa8H
F9Y+nxKl0ZAWSQeq2qDnS9lqvBI8vmM9VdUNz5pTnW8+dQbih584sOxYpO0B
xlvl6yh2gHinmR57nu71tKxB1nRPanI+8hv1rJK7YanX+UG7vQ/caRQI/Hb2
1XkZzse2Jk25n002rfxXH+rGLTT9f4kxwXLaDEe4gx5l0u4bmSzB5Pu5wz0q
glcBx3se5It3dJ1G1dr3TGfU/LxKA7jK0GRrwyyp0pz4OfL9ihAvB+xiaaaQ
Bgi3zZWREK1lvXHQ1wXPGLNnzPJZ+DSie/jf6CevbEndFkY58N4Cx1sUmZCT
DXznF9MNi7ZKr2K6GwyRddrNi/dpFptBHPet5OOBEvnaq1GPMrFA0851xT5l
Ry8jqViRD+cxH1/iD4CzY04pYq6kzYHr5F1EwbSZBYBhdgZslqmlJXlwT1Ad
nrviDcZDRgkFDEdUo8neaTXAG/ya5bDxkX7Wv2J1+WMbTelOyK4jz2iG+5VX
OAFhUuZ+pSElvcqPRiIRQtOvLaU9XgARUbOdORHQBcUIHJpLI4u5aUsDz3qc
y1kpV5xJ9meOAAXXvhAUxNcGAvKWSY58NvHnAAHjdRL94LTsQD6rx4zH5HoP
eF6uln0LoDcbq8w36D79YXaW+BpzDYHpSuLsb0xgxD3Mo/47TUOeYRhs3pun
rxZXOdzUfWVADvJyZ1KncP3djI1qRvf0zcSAzwVLLNvPDicf0GonmmcWFnxw
92/2vUR+ChVboE6SxFMtYb1ON8sOFgTogI/yevqw20AMhF7P1+/Jm0YorVAk
lnzfs780PWKy8E4sBWvCQ2PoccSIOwm564qqShyGw8cyN8aAOsHQSqAH0M+2
VLVp+KZWbblsI4wFmJUYZ1xaOyrwn1BkXXpFsDrZRIPleBwgof4yjrHAghUD
G2paNnpMti0oVv8xAHAOkiqfxQiHIm14edOTT8+x16B1xXO1+veCubLwXEhc
5iSw1IOvojvOJv8Pq2HCRiYXAx6t6TJnuvk3pwgfLPmPBtEjVfrjO7jAnOZw
2Rq4C0Y2GS894OYRXCpbTDeC7NHoNnO6bySPQa2OKhV70bViVUDFohd748h4
H/BOAyJ06nigl9nIFJvBEE+SIR5PNTLQTZlBct8LLhfLApbYbqYPd5QMpg57
pLqnH6kMY6mrO12hqHG78ZC+54LeRXZXwxcItrDfKJDyhgNev9DVarbjFpRZ
wosDvoCYsvlp6td8oVxLGmEi2PpfeCef0rl/N8udWLmNIZm1lyoBj31PghWD
UJzEWixZh48/lGYcAOaf9VO1VDXwvTJ/FzR9UrYobHl/2c/rgsCk+tIufX+y
QHPoZbzjakIdCp3HlETjPyv4YEB7GA4eO15uWlskV5F2rtLIu3YkM0ErcNc6
oOkcfIk4lfHDbs8jqWnloOpIGBVKi5iObdetovlafzS+JUiqOvYKsuqkqpSl
tIaY6lg/is5xnmiwk3A5pvqfo9B7zQeJgA2u/NCGiriwn4dwbZubFIBnVREC
MGU/CNQMibkCIEz6llD8ILOlx4rWaXkvu1kng9ZTzdUHgbZ5YkBy+FTIk5dA
jbOGgKrGPMxE8cg8mC+ZkxV6KGWh+KwFIOBWKa87SkiHCbuwTOcqwGjunulU
RJcMQs1A6BZEA+t6GZmEf9Jaz8rlgOcpnHUpmXBXspib0SulyFC0Jx56pM2L
lCvXMbCGCmXzWyNPCe90zFyHQBuq28FBwvprMC+PfDvqvgU0R4FRl2GY4HpF
s9tNUKCRgcdm/6nn2+SVuYzz9Om/NCcpTtcoh8FZIz76gFfW5j7vjM+43/BU
x5Ap0uIzAOngHrk/Jss6RinMiNv2mq1jxzMAADAxieLM/XQv6xO+gChnH/13
MD0DU2xDGmyV3ve5KBCQdeccOfdwAwycE/7UU+q9AB9pnWM4QLtSHiY3a2IC
MvPf0bgvJqo6oebUAbSzvY1YAuVQM9BxlxObSiQnc1E8Qlk2HOLDZMkTCYGt
gUwl8nHKnD4uJOK/urFCtz9QQKcJjRT8V+pq+ypHvHV+ukrZg9+y1gXz9Lm+
zPcNshNsfCbTWMeciWklMXwWFTfp80n7cUZ4Zp/c45t7Zl/fMky5JFMvx3dO
N3gIOV6bq4jALh385y6dZb8y8PzAsxgqflCILy16yxGQjqH3mdozNpaxg2my
+YuG7beqORhIjgPXjyePOsSm7gCvFOgpnARAFHUlmPzNwCgzeIF6i1pTlle8
92LnEIFQTqYJ98B08plO7u5622AQD7v8p9bcBTJcTWnDZ5Hc0d9ds0NKjT2L
PrzCVd0Ie1b+pMtRcAxeULlfRbB4p/u9v2oZc2JErm6O+Nb1og/P0KpyVCxW
R6XnXbTtpgUqwNtupp8gGMB1lx2IVult4sGgbt1Wdrh2J/fpr9buHc2L63Dm
57yzlWaezwaIiTGVI1IJaKN36L21mp9YueW8VohBFQkap/gUP9fNOZXftl3Q
S49w4LDY1LkFoYjU5OzGwMsZR/V65xKD/XgqLbwLnr7q+jW5zXn64kyIKgPc
Sg2gwNNcyPKNRj2jL4QfGOc2GknRMvgoDc2kIjDPNBG1vMPFbVz7s/JpU08m
+/cDdma4qn80OTpEExFN0QcBigufBIWN/7Ea/Gva1eWzi0Zx7xcvhitw+441
kYrr4j8HyEdC7djxXISHyZnfRMQA+eD84lcOOehWKuVEwMCpPk1G3CXiGxmh
/a3JCp5j7D2UreDi/l4cvbe8dUJ16Fex35Cteaj6zA3fbfqfoW0dNRUQoNkG
RoR6rAPC4km9a2MkT86kj2HaAozuagStqMUDzdaXxK1O8/omgCI2uiVjeVdk
zevCIJVl4ptymZnLUoGeR4/UlqxMVybhHP95h7QYvm3UN3XPrp8xNlTWvGK9
0s0itqfjsdU9a/1qdkz+nWuVA97koliLWs4aQAnQ3miPDiahp3eGnzmz5Ozq
pSR33GV43D0laEvmWMB23GXiOn0yMVv+69uCS/uN53H4mLpp8HwHNyYKyYVg
NxZnUZC9YfoigUG0Oz4m5LHjcXTwneE81+5zqtgd+okfie6R1eHsFXGrcL2e
29HdUa78VIyAadoAoegzG916nsxW+cIXlD65Yb5EkzSu19DBp6ESI/CjOMDe
8s9QhKPS2nLbvPtAcq/hsDDNASBsEymJZ4j7POztYdT/AzFr3uaa6T+5Nk6x
7SemVTOL4sDots/cWI89UDxXSgjyIEFnDzUZqYZ1xWacsQdGZZt7dh91lqeW
ODCiK76v3R7nMKdwqrDLZx+VVRgZIw5ekVFG5Xgru7FM8VFw0ndC73wDf5al
8561UgDC9nALD74CJ94KBwRN++sXd/0VeFBQHwmMMLpUyH2WJu784HvvOa5a
iHVWKHjOgfYR0c4McIqAaEKuKM8P6vjzW6gqy8LmfZiAC9dKh5VUUj/pHzCr
dVmjoZ8dOBz1nQqr+KWq4Vxtsb3pM4SQmZSnW8MELbHKj6Nw4TKKuKXk8O4R
ltfI37FrF27P92HO574RebhwdkLdeuGO4xe526j0CcVRlTNNswY66JV9A2P4
MbON19lfzVF5E/N8/qj8FG/f5/FdDAqs+rBJ5sDH0V/QtNT/AP2evSYhx8Er
ilygqTjpXr+PHPWYYhDn84nwxLOb3xTcceVaF+OhTNqHsX2XGFzgvl8dz+nq
6V/Z8JF09+Di4tkK14sd29dDqbWxFozekSIut1AjhV+0y21nqj0TVTLVYtsI
YPWWFZm+/ONeeXbJ0Dn1NdfwHj7Q6wjej+o9pf/RtPZQq/AH17kA56Lj33pl
vK/17opQAvtpWEMEkPTAyZudPSxO9nd21LEKz91yjmiRtjLiUuSdkeAmoxi/
eJgT0sVlo0u0slwHzCBWMpgFFbyB+LKEUn1ehK1H4EfAPM0feTMLHC4GbzL8
bPNVh+BRh3QuTYHHyOf2MiPABY2sl+Ul/H0GN7xj9u7m4Kerc6x1UHbEPdfQ
H6LZ9PeIlxn91jfBNUKsJq2rB5uNBJYY61dguXUa32NNbsneZ66vDiPEmBSD
AwNlsrr8tQ4DH+FIKKK1Cj1vEhadzMH9F4vThrfzEahB6/tqFHMTDqZCFtRb
gvU3gtnG2bOYe7inFo4wNTJgRnLmM4EAO+W0KG6TpNeS1TNVijMGvACOjTxf
cHr7N7d0dagrwAVgZt4kY9sAJnF0PBY+XbnPKpVerN9R1sb1J9dKa2amUMjZ
XEsOodi37U2JKP7fERuRz8qR8Qm9oGMXxjubRKZTYx7JrPn0+oMcDMt+vQi2
fQMtcxFgh/vIZPsdfcedHryYsR2bM1j6SHSpB9p+rD1llF8IeebVx/TWaP1D
8SGICfMBh6R9EXTu+ec5EipYrbIAtGTznG7hjsX23xKcmcDzNcF7R7RH544C
rVp/m6JZYiOYI9y7uQC/F/LQIjEjX6psBuiOhFvCnvDMQ80bsYccg40E93m4
Qnb7K55R9raT1Gnig/E7RM0fDuYhRBEzCFtR2qGlMUlMWwWPOs08q7oY8BDN
98L+Xhwp8+bD75kfA8CkuP2O9gGJ+egB94VwBoy6qB85G+CHravLCjwTRzBv
IUqSrpP5jwXrakepry1NUJvYpDpP85ZeKzWi8IAsNO3q0SHpj2ZdeFwikZNB
/p7OUY7MRcF0uQdz+Iw9pugBskS52vjYwL+34cQUhHQQVoL9n4NdjHBEPjL1
uCdZa0qZxZblTm1Kh8rR2GoCRKrlqpnQ01n/csyMLeNhLXLPQwIdkzmdb2er
Uok5xZpi3+/mdfKG6ruZf+H5PRsOA4OsDNDsfo43XSviwNrJC8Va9swQq2OR
un1y7pVp5o28f0+PfaiJ/oiitWRiHyMFNaqEYfovV5BrfZVbsTe42tV0zNYU
tlNEelRv/g7J0XTJwsOcXkbTGew1kz5zFFq4QmSFMTQkURHZUBGudGRnd3hJ
9pIMHrHo3t65k8hI7EKSy0YeDFMFTOPqh7EnzhgnY5FcE4mhGDVVyJ29LqqC
BC1kM+lIpmX1zq8CpAxcP5Gj1xV6MVrNLtLoJorEhxnDCSTaUpmzSmp+ZmN9
Uv9UvaYbCYhZoJxc1HQV7kLE30N8UK0Wi+C3KdjDcXzqtB6CvJK2d+Q4PxS+
aOpR9zaOTUe0xUHBYJdVqV1gEz2YDn1/6yc0W0BRfE/uCZx5756xoQXSeASU
J/SNwViwxQMUtImgFu2qScFRXloqZM5Y7xIjtAdGWsGac4Z7gOzYxuO4IXc3
uPwc5Gjgc9iO8Mi+3eixK7HSpBx2nb2yzbSdU+L7tcI9w0ccm3Wjf3tQC8Zh
DtjRHxF3IiFxmPQegu7zjJAh9mnnHxXjiMgnnqyFWREEBOB9z2sv4aF6wF+6
EwMrmxYLQ/i6rzlzWiexOHjPA2JhHuWowK/goUB0SgWVwB1l7JO1woPEmWvV
rHFDsGnrRm2CxddpFWb/nB0ihqNAnQGNPomffYihjw+KjhzglKg9d40z3s3D
K93O72ptVGkZDSRWc2wrZd3CoWD/0tffCq6ymm1iDIv4RDv/BOEedhtq6joG
NjNFKH8jl8BPc0+HPu94pxfpguZnMiFWt74KSU0gvVALGFW3YTw5quqG0ro4
vVJymPc4OWiJ0gV9vZkYAj2eF+e5zDKTR6Sjdp5+Yk+ySWVoFcFtGXI9+X35
jp+yOB2SsI5CfmTRuLbSub4wAViHl3xEVY34wZnyW1IkenglPv1+1H7nmsQ4
OHYc7KgSJB1WZIO5xWdiWA3B4fC6ObHVmqP7WDL/X8LJB0KFm6rRVN/ot5i6
5bi/hxfwfYeZnBdK9PSz0L/AZaXY8ZsVXeQJ48ilnled/odk76e/aTtvL/Es
MgR9U+JxjUeKzoUCC37NHBGsVtziimQHKfTjUzrFUe2ipveVNTkWy6yuRN8b
7y0/12WPYaCHYlMvOtewsM1ptxKIcQhUc2VpaY/Ie3CEYzRBuOszQEOIvoWa
dPSnOWFejmfdCZULoeUFd68X8GSMuuZimyDsA0TcBQ7vvKQE+xqzSQ05O2Hz
0a1YI/j1OFlgywHQc2Gi3/YCwPLuDiqE6wWsa6LKNqzj4HymjR872ouILdYr
iHvS57udRTHPHMLRgNndBa88hfdNQZwWTmxD6+YVamfMSeZcXsJSLAp95ipL
+eSoS/riaVc89h6c+7Rr4ALNyQ9VqeyA5D7sPnH//htnUOcIvDwXm516+kVd
+ohaVrMKydnetriRUKPQt1TjKzj8/GAJnmsXMysoG30PDqzWBFXD9rDKqEEl
hgDVFJdoaemzGrAG/Vx2lYf+8c8tKw37xE9Rmz69S4xepnBbrHxfOoPkiWa3
VLa/xCCFCBD6l0CZcM1JVy1U/nG5seiOrbeDZTwL63N7dnkW3MdqAer2IWTl
d4jUFb6gV9mcNSOMnpy7yEDHwR9cyzxNUI0kfp4DpzgbEH/d2QHzC2VzqB+Q
OFHQrvrSsgN+po5RRhZgM7/pvB5c4nIHUDFHGxZZEdEZdkJAANLYzl3BCzyP
kB3MuYNB5wmDcm2+wdxYK1Z2POsDffYKFdQHpN4g3S9TA7JytqS4pZloQbIj
DWQDI8S4hmN/PqLr6nKRmrH6o60zD84JpmkXGQLt2zxoMExVDUFovQOP/ctw
dTWDtYBW7nS440HwQ/BMAfHmEdrHG5D6wVGorsO4ZnqJSQOWS8hEReFBnARe
DjYep1r9a/zrtZB1QMyRNssDeiKz+iUIS5Ve4CdIxU4aeG90jbkXI2f2MiC4
wh3/BwAFsmiPny8oMaSKWpWLCZUMwK4G04PIJwM7dnyo59J3v/5KX3jFL29D
dFERt9bnvj/Ga3JzPt2FBCu6LhQ9pDc7U9AaYPFt9/X92c/RsJFMuNETgmqR
iaxppNCHf0G5qlSRA5PTBr83HzQE/8uJChPJZZw7+ibbzok1ZGRBkPf7NtkE
4AhMFX/I4Aa75AjVAFaniXvpq02oq8jmHD8DXx0xS+YNLV2CChJ/3aoE39SW
rXnP8w9R53WyvoVlKIAs+QGjEXeZKm58Mcjczb6Ijekyc36X3MSlgUJNGEPc
O3zA/m3Da77MNxKaql7ZFaaU5STICo+cjwnrznUm94xRzCEv7hNLQsm07h0Z
W/JJXXfxBs4kDvq/2jMH7OrXB9DN/a9QqqCiPSq0S6Mn2IizCDcYQDKPatKO
cdAJGxVKg6ZpNVh7foFCGC0mvXnO7rQJ2ithem9qEeoHzR9595XLeJ2Xsf7F
Fch8IKQ8z99ZtE4EHbVt42J2JxangeW7HjE+WvYBQA0gLtg+nEhKjGCX6Ps/
ZCwxWhk4MwtyusTMzE7Cj3FZAkcCSQ20+xiFCM2eQdPOYiccQNferWqkPhvK
yk2V3B9dwgL/MEVHVUtrVUH9bd+RGqE8HWufhyah+aX5XuIAjo7t8HiHjP7n
CMi7FwVttP4awF7sKVBJ9j1VtjLTKXACYypf9+0JU/jOOgmPKL/IC7LUGGGF
OR39+11JwsPRi6x9o0lT53K/oNif/pbi/ojDCs+3jpciIBPQGzj+ec/lGYEX
O73pt8J6yAT8s1ADgXFxocfapk4/L0pHXHqa07XntDXwkcUQLWlT4w0Ux2tg
NBrhScQ7yIwvzDNAvua/rXUJAuZYk11AxHBV3uSzUFi1McfcTonK39Yg4wMi
pCGukX4oajEKBOgFCviQTywn5inytM7oyd/L8y0Lp1ow/sdyb8voj7BxYChh
iEDk0VnSq2Ku4Hj+o54Q51DRLoKaft6x86e9A0xoYzmlDleJXTWdGh9QDgVK
n1MF1I1Pc7g3/zjn1P6YxD6/Ixu8zkAHE2d9eCP5kuJfuEtv1/WG4aofcheb
sGdSyeX721eMS8gCL+YSly24Ph/VvbfyI3L0ahaZrCmy8Vv5yAIRqSk0Zz45
sEHtnMcisd+8225lP+zDIVXH8x8INauCr7GGNkLn3+Dw34jDhDV+JQZgOVKY
oE/gs6hj99PNA0l5d8euBD6ZHBcvwamc71b6QWGIfWP/CkKM3EObfwPUAJFy
lZo5FXeUzOSRqKH26P/WWs81MKTPNSNhtTuZYF7h5yXyFBSFdB/oIWJJaUMT
+ltXnwJbQYoFgJu29i7gK+Z5rf6yeF7vZO7SU/PTV56Y8fUkUkWdD8uUE7vH
XM0hRa9CqhC3AMgm0WC+M5X2WozKty7TW4UVEEYL5MYxEyXi3Jb5L8qydV4e
BwKf/H4saIxfzwefKYdqnh7yUhu+LYuTqaASh5Ra3elYnH/w2SuvjsRYG54F
6kK6IPK2vv5HxEtVT77/wCx3sWYiSqMJKXkf2HRsQZdm2GWI4LYnwZXCbCNi
A/h8IlZOTgLSBAkSCuv/34MetrwiX1KpFHIp/fOg6V1MadTyezTp7mA+tl7I
ENZJ4k9bhg3vAaXT4aw+nUa0G++BfVfQUKryP/mr8XYzuwreZHuCsNiaf/Kb
iczxhL2559Pe+XLi6lfpRR1tN2k+V3HolWU/N+i6uqp/jTrvo1OAkSgDZUw6
RHYiymK1GZhi1bFOhEGrFwW1YittuJHkfNvozXxXkvyHu/muu9GrkiLQXYj1
DS/2cJIo+dC+6NJJstS/f+4qnDP+IRSMtEoZzd00g9HjfT+G9N0khxxiEBuE
Ahr7akW4bAlGzMkN5jnviqXUgYXXd61/RR8e4Gf62i1OKWqZqFv1NkICUFiA
AsOvolxXW7RhgBrlCbRJ/v+4nvDdvmh8vcz5UsEGzbrYaRZWR6eZf0SAhybj
MTTgSZ2hWYIDTaW3SCDJ13aZgGJxwA4x/yo621NM0skIpOxr2aR8zAQw9tTR
IEAGJ2SK0IZwxf1WjIEXVl9n6KQkQnpnj5fovTYAsPdT8/xlkLZJARgslVQw
GvcPTncCgRyjcMqguuu+CCetf4K0oK8uYHnCIfxKTyQTlVrJ4THbb0jGLwGD
V1jwVSKmgJdjWNtgAI8lLjNuC0+q/jN9NbBmq765r6Tv0EL9/lryfPLnMjHJ
YB2A0TqmptU06OpkHdDLoSOnrP8LbwQTfZezeIfepDhyN/dzNvdHwcVZkhL7
8N3wM8HAzmP9boMuk3ndjEq5JwrF1iXvGZw7OMmwQOTrDDmRAYm+HGcmtVba
fAZh6einfqIhxvnjplrgBvdzfZRNZS5grBxzPF580fZwFT2V9yPl1F6Xz9m3
Gdo0VONREJjL+luoBCN/qoGFSLRFAO5ZGckdWN0nwjQdvvSiijJR9TdyN9kF
1mqQuWRsrvX8w/8WrIi7/icFGmrcdTRdvaRlALHQRJYlsSCZROTWH9zeyBSN
3H+n2nzB+wXDhH5bpBqzasmWj9i+5A5m+OpVeOq8QgritoBQSd9DLeyPjvjx
p04UUHXFfFeeQvorV6HecJiMvTpGucIWESKNvJ+euY9JNuD+ngYeBDjG0nbj
P3apGudP0Pfdz5YJHpkSVqTY5S0uxP+ciC9hV89C7cSTkFxQHDYC2Mbo2UWO
yV9ka4QgOtFlFtfTKyJPbvRkIaPab/LUpCHfGY7kIQcmtc+e/zDz1xZe/Pcs
IOoYjJymmY7CX4q7+Od43eMy7tPG5yTl94bLeaRkWkZCoso8awehF7GkuoMJ
2d4qHJ6bUeQMO0SXhRSjymXfLIDZDKXNWemT3XnCPDx0QYzyWCYsnASSzSky
VUphLg6Eepg0KDFk8M4lse6W9l3UYlPyUdu4CNbIjnxwkkzcC7Gn4fAGjJBi
zMd937psYXOGXaEI59CU5rQ05KhqEv0iWzBM0PwzRfkxwkCn1Tb6DtECribM
+pQxaJ2AOGfVHRE1x3649gm37sOx0smnIJ7qjBqr9fnN1iaweqN2wKCKS36D
TpjqsCAsYazOe9u5OEDyWcGeBEp0ZkXQ9xL5tBu53d4VxSq4mKy6KcuRd/ue
Rtohya9O1wNAJ3OCaGrtdvszkzs33J22sHbeM3k63vfkh6/jm+vhsvMYzOTi
WOcZAn/mi7nKytX2zDF+7W6DrDR/5VBtU0zd2PTvbQDCYatwNgP0RaVzVt6Q
r7Yd/ZJIv0Di3JZ4x0ZNHjDa8GXyjb+rq0l0YGm5bBU12LRWUYw2weR42Z2d
lBMRR1LT6qsQbHsIpuWG7iRbqHPauRAECLD0YHwjwkbGLtLf0RqJoNyFsdHT
8Kuti9M5BdEGYfV/tkFmHeUvfynHheRHwfxx7zkuxukY8GHLQ0is0FRCnRv/
cicwedjO1nE09ucjJhz0bWyf8SNMWXFc3Ac9JbCP14X1kZM4RVqJsRpvvLPl
4QEEn3y+djHuVyGzrDDD3G74apkPtt774LchKIF4tS49QGQ8EfKvudV3QWgX
q/cEB0dd4xemhzYjmLjaBH6DE4ZEMeoRGUXd6YIBVRRn+AtGRCKD9GVO8oTY
os/nfMVrBWGED6wyt2GqAXIT7uoQgEy5o0G63ewSlNlY4u9vgAUbNEJ3/NST
j6fq1lqHRtSnnQftPmVhvzkqfZZoWGjagXuvqvla+Dm9JyReBjEP0ulvSqn1
gKqKUz56bA6PwdBGyNGhV5J7SAIaFA5RDvMw9wYbwA53ffPIxHHdGCyqH+bE
E9vRsWijsbc7YaFQXy1jw4J624P2YwJIklC7+huuPba8eSoZzznjLdE5XYJz
J7y67eI3pmXwVc5hqzQjB/U/HZYwseHcVQD8o2O+OfOpY8LUMqBeVosfb283
XuZKUekAYd9gh8WbFdERPeAnH1SFDs5kGCcUwYB93ZQa/hx3ll96pH0yNvdH
gK7q4O2IEFGL34zFBPNxauIVL5C+qDiLufbMS/pOUBItua/flEGH/SlLVZHw
X9Nhwlgo8Wgx92icTY4LU4MBrIIRRAhbyhHtJU+TBaLDmnk1UMpFbzMDVl0D
x/i5mslJFpn8AOaVsyyclRMqKmCJizI0342JNQ9yvINR80JTG2H4TKIqKyze
g1ZMS9N/9Wah30+0EAKBgV4CbpgxLvvDAJiLZIRPmPwfcfqyz6i/JKkVq4KV
4VgFwniq0E5uefnEySqmWP3gYNjtusWpvX1ZFrmUIFktONKR44c99fCJD0lC
kx2n2UCz3DUCM+peaNC36pfdzS9wjC9yicSoeSmoDzvrp6EGk9XNdfZXl0RV
bxFr9B7y6T3OTry4RzV9iULg5Sh6LcimOYXDYLQFaJnYQUhqg6FWBIt8tqtg
NAp5kfapTv2aX0D6HNWDKmh4RCQ2Ppfmr4nlWwT2pKwZWAzhHq4JS+jWypP5
1GB9SF/pIUb+GiwYok39SGyhOfK/gJuEMF159OS9arHthHUvlmggCuTZ1fJJ
M+WH7ZYyArhfCzYLiv4d9WEfiBvZPcbjn3Ar0GIp4kKuDNPb22I2DnvYGIub
BSaeO+wvgVG0EyKZJUxAs5ZUhsSchlZrTWca43qdFU+WL14PqJzWU3UIWU8S
8oNjHzNthHHJhfHiz4qgGRy0sYcyV2OQc2dhf97pTd6TzVQSNSHJPuupvJgO
Eg3dspfyuQ2c3K/YrJHFH54k6UvD46ZNsr1flDSOssVbjDiYUdMhtlk/bgjz
q4qI8B2SRiWO2sYU+xhsV1el0zh2sWg8J2hh933U/oRMzOvJdTxOJJuw/WaV
pl3ZnEOtTzjE5xaGYa5W3H6yvMcF+6aGGdvWVtBibibwkxDdhbnh6vqEiN28
4YCWkI4QkmTte+aAuS7T8xhRNEa6faBmTwW1PuEl8T3TaJOzjoElh9Tx8Blt
pPXE6OBMBQ0r7Xy2boPn8uk5OwlybsRpA4j6J2SAlwEOnSEeGs2rY/VyE2Qy
0bSo1PpVdH9fHexGFHYII2RC8XVfpw8jwY9KQy7eS+GgvVRWsfWuRa93iVfn
dwwnZga/H3kT0Su1DdYyYjsiMJynVXdhOTHEPdtzEbzGnAkewEwmG8NcI6R5
bCgJ4V3iBqWaJboGXAnanB3GfdEkrBzqvbDIvKUpStZ/NbDSddrBbQASXDoM
drAYJwMmQKgw36ShBDAt4gj4hsfKA/BEd/ldZRcgo/q+wgEpFtGug1x/t4tC
Hw+gZI7QH4ji3lRIUK2hbPMwEuKFGxbJidknmO2t9pElnNpsxKmyrK+gPa/2
WuxW1L48WAZvHa/idm8aI9ttKtkoV6O3rZI6xHAPtoSkcOMaDN7ic+XItM7G
1sksMzHEAe+oOcmMkW89cyVx9Fl/PoPZj7cfEmXUHPqu5YNXbCUgnKJDM+9I
FUwDDVQL/xsUjYMWDopAYVnPSFC8LX30GsfqB2ulNiARXqBWJdRw9aJZh+2d
epgVkeq3IQvH1He82m8ND4qAeFLIykrJeUE225k+kpA9JdaIeOFySj4ytZtV
wGY3BuchTXnS6kFpwIx9f8Z3BgZGxLGtKOVZyHTAL0zaIjzdNOfHR+ZBDMee
C9AhLyuukRohhJ4W1t1ZzRclbDZEs9Sq2363Jd8g1Rw+yI3Dfx86muvTdEua
0qi/zK2A6aiImrVRRrCDMxAv9mSIxwFa6wgbvlhvTDprHPglnPGi0vJxTK+Z
29ep6EzEp352bptEsaKyZWgMLUvFLJQO/nQNCOPPACXcbDcg9ugpbOBgeXR2
vKpuWCpq5JBWhNQRLsJX6qH2zFnlJkwKl6ijCnSVaRSaLhfB4d1ZuXBlybCv
QgpAuD6ImtrpAJfgiSBb1NmVSN1Jk+vz+LJFe+KzdmGzY/kzuxUzyLeUekdf
y5GEJSlwk1uxo5Kau/fe4ZSKSjBodjNQu3lf5SG+n6btd1cUh4VYhP//1OGt
eILmx/56zxW8kCBnerRcHE5gireUXzScv0jv8WTNpRoFUpc/r4+bYBH2bu/g
zComaPDH2xg5RVzOvOXoPkxFtJdfJ2F1PVY7BZa67BBlXLHOmOKH2vKJFPWE
a/u3sGaQi9qBP4RpZkqqnlIRRXaZJSo1ZtbZBR4JrCY4Pwz5jvkWnl+BQeno
EVaWssqFY/Jh50br8gkqKM6YnMsV1p0B7vhMhwnHoY+FrUBhub7G69xH5QO6
cyn4u5TgqEPRliFho/CYGBQj3/A1foBGhjQ9ft0ZV6waxU1xFxwW5tvdyhhq
TQIKcGvtrVMUdb/KxSgU20IR73iEWk2nsn0jZR9AU6kHBdf0gedNwA/1LHsK
BZ4/VpoSK+cjXgC9sDOYU5jz7W786xbUqnasDaWnAg+pETqB31LPKsODxUyw
BxP8NSrOiZ9/1vXHL7HBUQckS5obqr9FTnVRLXssow6q8vFrGJl9AyQEuUki
Ffb7Crv+scuT67wm/WyPKJBqVuvqQGItX2wS23zRIrtI+Mk9ly+Gv75PJ+3c
uTAVtNvD024Fg5bZwtvjqy+uMUOnzwh4G63GIYG9HISANxOmGw5o4FfOm620
uf7Tn6aR80JtEGX9g54oop904kCoErShfWaNzUyuMeFbczZQWZjtFhJLW0LE
7uy+yXJVdU9TNa5DqOMxndM6AsEAlSGQmsx4QC0G7QFNUKXCwVbXo3I6ZrFJ
Sbi9Gk56FL701rcbTBOfG8xe34c2ALq5dsk3dGOPrKJFSLXNhTlBz2VHSuJd
0wNvyX/6OcW5MxtIrWbZX7PAECr8SNUB88LY8+EELB+WJLKB+b2jKKHA17+X
tyTzB0+UFnwTZQ0cROQzR6NnSZ5uZlGL4G/T4HzWvQ3CPrE660rHRlSYR1DG
hiPf3e/Gf8z4F37uoG/SARVi5qYvXNoNotFzAsmyPg4SFAsBo2fy45HHrbjY
/aELQFIRb1digwWn5cp7g/anUx4wg1ksYXgt3hBin9lQHxCeOLOPHtKlyfru
9hirIpmmGcDqHXFtQmXR9mqHuIhWdzy/SDmcRo6Ly54Lbdmn3hvTySXYxG8A
n5spE5imGsbTqODSfECYrXgUd/JBbemlBM/fypAy4L0SLnazr6DEeCBCNqly
98YJFQnVyfzmp/rUfDRPk4kUwOak1CgdZjgkSt/CJTKKBqSt+yITNI4sGTAX
4p8+5ZNfO1A3LBr8lp0tc/ZRMtOvKuhlTLk7v7zkFJU9KTPa3Xhs00tGz0np
8iRa7XJIJxw87pAR/1kPOAIGyNOWATH3yHyeoBZ9NKFQ/hzWYNb1OHurqas6
e7rIKsDSaKwSelmKE5rKCtm4dZG4dEIMkFjVzeKIvjWm3EWcipZ6knYYbzO+
7sWTwUQ16Yz90Ze/YtTFIpAD9OKyUPMcYKdiTHAc0qV7AXzxZhyWDajnxGTq
bOfwV5UPe0MXyZJh1TuIE5kIm7auSy6JsQfCVIgnjnD3rxSFOdPGfSBVJO1o
DE40NmqJBdWXf/JNAvUhTrz9bgjWgLdbJZXgrIH+Jq16qn6N/nAGVhPB3Mx+
K1jmrKgOvKwexH3VSb1/AlVks5D67v4iuJtmaWNBSB2Q4n+JhsP7f4LM3r2w
3W99ct762DQsIET/+yYYsXhOk812QO8T+ABx1iczTg6rxyEJ1s401vj/Yute
NODfJ2Y3CjJWLea09CLOg4b8oU9Xx6zES6S3eCjldNm62/aTK+QtIGD4RosT
lmRbyRu5RYKF4P/Ldf76jTDzNysdgtSgRznAnGk/vpg0wm0KC0tObCiF0l5c
vimRxr1WVPMu6JqzmQE0NwNSP/gCExHH2pZk5KqJgCfyDqDbmgYeuf5gnfIY
gpaqUqWJ7kOgHdVvBcEPU1WNIz9RUag3k/DnGgJ2KVGJBW98XnMXMw1LYOIP
iYTeyezLcJMHOsyGYspbuABsSq9q98jUbxzLbQaXCbBdvLYWs2kXKSqIXIwM
+5do98a1z+761wz1ct8wOvayYdHjxiSpQGv/I6YUKqKd7PmvKKfnTHeeYBgp
XS80KzpT37o2AdT9KxgVnkxMyp+2psTSpKGUAgJtmR7lij03eQDZWxI7+sMu
u33uehc/qVjJ0EmbtBt16OBgpiYtcwn0QAS5MNkXpH8veOk7mPmRGFnoNR9l
E8hZbDNVsDkb2z7k2s8Oqk13YaKnvMse36wTjRNCmfqkepHqtwg86bY3EL/U
+FRa/DUu3p5WlAJXhrUfyiPbWLPv/0bxjcT4tRXGlq8zkQSbAFIQSFwwphQf
4BNnwo2q0OVd1E+N2IiW+iy0oXcgz/0xnGUe6qKG3C3tgwAa+gUMER1ffI8h
Wb7UoKdTm53ya9nRZntIEVdsorI2utEqDRXwokwkd8TwgbwI0NOaRTr58H5e
r5z+wFpQExGGE6YBs3LAJnXqaC19WnvK5np8ggtlAwK6jMPjGd+KBkUBObMs
TMzXWgVqUm30mdB6t62CLsZKaHmdMMbKs3GipwXwaIKHYpZxQl3P5o9pGOJ6
pLUWfGtrcXzwjMfKUnbm8TBPZWZwar4XkDQEr6k0gC24r98jFVxVj4gagxal
vXjs+5o/LBXHWE0aJmi4VeLQajnZwSo59HJWOSEQBIy6LhApOP12xal7OUnG
tfe2/ICPwhoQtAExn8AGLeiwyNwKVEhMIOp0oHlLwgB9hxAWb2INwVvtStiC
BdyHXnOnOWreY1dlihSutEm5iCpx3CjaMMz1K6sm7PQmF0sqFgWqtGk7XCBb
m17b4QHckUJkOzudVg+1Znqt5ieA77rN2mMxnQWrhTPT+s/ZmLW/pzSXXMPq
fE7P/T8UDy0hm6/cEoa+RSK9ryGvucusdGCbni5zYoZ+f7DexcPTDA9JuxY9
ZsgQo0dDaDc2qJfUXiIweExTLu49lo+Mp0EhYFu7qkhhzebAKhYm031jrVY3
0h8iRdWVZ+fTI3xkg8j0T0IPqL7bRF43RB9aaIjyYc/HGcmptETGCpReqNEO
nFujqpnSJUdr+/mFVf7gudZdJq7yM70VtQPKbdRzQhg41ZFjAiTK3FPbcVCD
rtDgIrzkfVhGsxftStA6+5UFntio5xshJACHiMHkxyBexhJ6vPN1bl0d+601
FHN8VEZxjo8mgnJNRsyfzN0+jcfkWSPjJoThAdjv275RhzhObnHPznEUCEds
s/6iE9wbSKicyhJ8FBfyaBvHaDXa9qDQdOgw1rBK1uqRSF/+0Gtb6gKDJ1LZ
TDMYCTij7qAI/EGz3m9QMU/8Gy/HoN4mQ1ktWtrppZiEgbiy33dPPxqtutWe
hys6rWX0AoHSFmNPCS1xIj1BaegBiZapAOlwsGNhD1TrTzen8tfMOOObZwWa
MaAOz1O22yeBXoihYaDi9uv+0KLorx3/nVAfcEto7XCPMme1iYFm5pqEiwgK
p8HpHJMUYF4TSiRpl0jxjLFgqDbqRTavgkhUAc/qZHy7pkT2Q0DzrQJJQS2G
b6ZHrV2u2WxB/XfRp1WVNVr/awp0t37dQEy1MODTMQG/wJ91ptRJQpejfCBz
0EaeXk6zXTKHtDkyrIGpqep+8iqPKiBJxxSvJNN2lbOsP2qP+21kZEQt0W4D
YFtajfH/fH3i6ZmwkhiqQnOBoWxIhnWHn9PvDtW9MOGL6AV3QFka366w6HmD
cZXiktup4phE3BuM22Bz4H1vEo0Vk/17uCk0J7omfp4iicyMIMkEAP+6ai4/
MNPQmjnszHUD1+ebWoyY3/E0MVhRWWZKksYnnRv58lzb0mkjyLiWrv8LQgng
WaK9mqlV3w1HZod60/2a0QLT5diyFEdhibeDQ1LrABEiIFoYPRlQ7nfNqoa8
XX5tGvN/2aHjERfYdaS21YmNyCp47FZahLC2wNZ3hReF4ACrR3zS4TFhiVFI
4RBYLwLfPxLoiRVUNCAQfRQf/6sZB0ajr6d9mQiaVCiPXZLiqMKWkV1fNBdr
ZtRIc7a0IBidFGQDBjWAvf101c2UNaNiLsXY47j1AxlBlHOrTuHJbAO4yAxN
frolIB94l3e0B87mkN+sg87ajtpyEeXfCWUXENDEwduIa/iqL+pn4dm4vrdr
AlD5YeE5PWqj5V+wfP8ujcZhIbQvaHkcWcY6laESYSfSr+gI1ai81nCrwQkW
Nm5LtE7PjjFm5MS9CR8ZjgV6mALyNQfHup7knvOWsz+BX2R5W9cHHX/XGK7l
JhKQV2gsgQ/zbiY6UzX2H6LUimGdNpZIZWffxpMGQPJXz9RUGzU4IDPeb0ON
J5nRDvQzoDVUIE4O6+OcrDyTKI9uP8gCpv4/7BDvi2NY6o8DfVBBIqwK/I2r
KTQh/oRrJ4I6WOjLJzEHp3s/5sbM/46nUnhDynR0cLqqtSJo4AVutnej4MSb
1e0wDAr18K2D1Nh09HBfdzlhvKVNKdFD5V55F4ctaCyHvocwoOYN/IlLZeF6
sq9iuhrUtR6yJxYqIrLvaptL5Wl4uZyQiiaEacXlXyNGUz6HJYxpLFfNzyJ2
rHHBjvqzvrhjYkSVGAjSiAaE1kqz7Aigx7UJCDmmDzYqK8ZCGHxoQ5n6+u3h
w8Djg/F3lEJEdoguTvWspBvI144JHXzhAa+RSzDekY79JDVrLjZiAChPfcSz
aPJhoNJ7JdI6a6gbhxO3uUzrO+1x9u4AKhf4R957MeHkO6kCXdjHBS8OmbdI
sXoIozlVArzd3rz9zTsfvF377S3AbcSW7k4NVmRfZt3/3Vhd9GUL07vdUuKm
MukZ+Q8l6Mrp0nKzRqmR6HVQE0JpuFeaBtyVsFRH+GKl+txqbOtxIaRX/Wa4
OBC8bDhcEtFvIG5WI8kXdlnZOwDiN30fQ7aBYwe2YZyQIu9eTySNLHmJIFrb
c2wwitXefMio72mH+ECc8eFD+MdTv/TxdH6Qms3rLwFPLOZ9GZivXzCMACEm
E46AJdx8sOjJuUk35+bTBTurLysqdyXaGsEKEVU7C0w4336KevS1HEWv38FR
EA6O9rc1muZyQK5JYpK8tqxTSpQx+EHuMf+lcovMsATjkIeSQv5Xi+aREh33
5jhy7B5UqbAPKtBC2I4M/a1gC53BCHi7pgwi5ifFzNl57i/1gjdOzTyHMJSA
w97ckSQsriqrQaLakFAP6OUCxcHKE4o0DfVfzZhm0GyOAMKLYOv/oJR05SIG
BzCfa1gpW52a0kSBBxnkJMNtg7yd9Z5Z+Sq7Tmv9MS3WTSadar3LJUyMZdQZ
HMFP3u7A33BjmoyKrXKIGn+cqeKqDLJE/p+4C2qdWIt58nS4fsx+N0u4zUZk
x19zS/dcM80mX+tdIIhnAaiCpH3ITHy6j4brqMyj6p8YxGYjbyIUBIeaqnV7
NAeNZHi96NyclyntdqE6VqB6TNy++ggNVKLvr3dwmWYVsPNHfgYHm7J7edyo
tAYUSUzPwk4aKFwVOCHUEmbzpbKuZpIWtVjyFwM0jiUSYZdiLDmeGRb6BaMP
2ARAPsED3Xk7fU36iGP4RR4i1if6itrdAnDTuPdBDKFmGNv+wZ8ulFlWp3Vg
MmKWZHAip3aw3Zhl+Z++p0M70eTchxvh0v9O8aAvzdixVEAI6aWel9hFIo0d
CxmUacLLNdx2kMPg5h991g7M1AuXXlZsahvyn9wKzpkaKKYPOQd8IWuko1Y9
LrOkQjQwvpsAYJqJLN1CoO0TzfIjIEsHkFj0SxLPMDV0KX2C9c4Ganp+QmZB
IROyxTS/umxfQWc8Qo0Hsujpyybewkzo/2Q4hy+OsFLpiwtejws2ZsQVelPf
JbyWOd2QIlYWq3HcCT/MpnOv53u5rBWBisuxLKx6OUmUmaK7UVhliudHsgA4
0fFx2Wkmq4R2pk0s0t9Uze8osm16edbQrJnOf34vx3jqVbPAMoORTxS0Hmsm
I7YCinuRzSM6fQnp4X3lLvT7pcspVVQmEGYcDy35CNslxS7ph6SeDKZrcXuQ
CLYZDHq5X7KEuuaj2OVDSWIbRCXlAo4W8lIIIx+zaGQJPrVPIEqTU49+m+hg
Yue6V+1wAfyvf8xlfqgSMCoBEkurV5AI5UEHHSDrKEeEXLO8K6iik7S441Dm
Lw7f5cTTYEDbQUjZnhSrwJwSQup3lvMj9uTrNTrjF6mEzdwUmcb4T328LHTm
Pton2SmaRFvryqXpYq091GNFyL1cZyHFY8AvEw3KbwDVGQ/jYCcOhfbJ/+ns
3ARAxFWL+G3DFUzogQT7Sjd5XpeVqmTD3DApWYJvjnMk0ZXwm8wzMGnqpDLo
3o9BflFK2pFxisChK95nKa1we4k+8jk/Kc+5QFU0fXqw70dUh8BMP9WR11rS
PGBMBdcPp5ELFkhVG0QQkXKsIYh3d3q7RhvU2SnImTe2FdOD0+MDaO8r2C0j
2wVIDbpcRY+mmbxtAQ6XcsaVonpV2tqKUuYgjxwJRvlwW+E9JLvAdB381qlF
pONYRWGnXzNIXR+jf4lWRGcvmYp52c2ACGx9h282Wn9cwlTs9GgdENzXh8ZN
ionr/ZPN/XtHN5ufWKJ8CwRxEhjTTj4muT5pHnUchmF+dGsaj7A2rygyS00L
juZJbgQ3rtt1L1K5iG+U53aCEJIYTyfJUnOhAA189hiRAwt2FW0Oj09dolsg
FEXXOnSPDubfjc/w+U9AID0U6M2DbTAywaQQ2n9tmN3qhIQEWqG0VF7tOigq
w0GMImHoKN1Hw0fzTc4v7VUoKMfr3Wqa6NM/WdOp7aaJNZk1uZOR5Hgh3mX+
jdUKX0Aj0RmWRcl0pZJ+gJuqvZO9zqKSMiu8dyH6/uUXykn4Vvr/DW2ZYaPB
17/wGtf31qDOEmrhgoUvD+VCF1iV8slaB/edykJbESUCA5EQsNnu6Z3EtDkO
72M92MSZOjqF19Cjf1irfbfn18JLiuPlhmgQOuDgWWi5w+UAh9HFR6inq1L2
QTQ1zHqKOMHsAyJbfVjvCzIqNPdQiERlahzOURMZqPflra+2acKkBfnAz+AN
IEKsWV+bCFS+kBkFNv5oRnC2svQniqpeKhSyhDKfJA7qEa6HJX0NJ5/cZUOn
LahQ+t1bLRLkuoxaUjfV9zGWDoodKSG0ix4sSvjQlzM72QgT7LQmfQqBB1QB
E+jbYkUEjl0uv4Rni8mgrkNCY4s4ya+bQwWa79nHuAeTG6w8jFVtUkZtJM99
DWvYTigQGBzjwR8LbMlerKkaqoGN+RovLz8mU5ZmLbhOdF33jtylZaLU6jlp
HlI2WOuLC5kbYCAdiZ5sgCI4+02J4pDTXqtKn5cRIfffjUhRnrxr+BfILsda
vlyRpJ3C9Rwx5ggJrHKRhBzQ3MjYqZHaHoRGJNpvuzqQrf/f0JY4C62eItS5
IDtq4W96QUEYTjsodGafTgRy0IwbpM+jw6Qn5IApy2ppFy5eegXAbhEZmYRI
MkVhTJLAYgPgDNqeSfakqIfBrDI+YwdU/F/fKiF/Cw36kzrGzOGfv4S2p0By
8mm9mttQVKkqanOrmq/tvrLL3pTIPna6JytQvU5zmanCtRfiH4uOkIyEoSm5
HurxVsuLQsXZwSQ1h+18GjgVHpjNDn1cdRIh+Hr9H642TPl4KQC2CLurecCv
hqeeVxbT/LaqaJfAbgZFO8LV+Cvt3dZjJMyamnrWk6rL7XHw0nh8lP1hGPEr
1+zr/CtG7/+7vCZZYbzpXApiMPMIL9pyEl7VkG88WgD8/1nwuGLAyBm8YRNe
eo73UIZyMc0qJ0+08QqdxUr3sMxMY+tl6b/h6PyWAOWPM9UeLGmhI1T8xV0m
eovCwr9KO0ZrusZKaMD6O/BuiZfPkDhpZSxyLf1j5Je6mYYagFdt/wzqxpPk
y67sGecFdG2uMb2gEinL5xZjSVA85Djh9eTuDmuEGLz4HeeH5tnyMbQo94X8
ScnP2XlqogDq56fg97DHeLdrfWuU63vPoAkXEa0+pUeYwVT+kinT6YSBKpnQ
d5x1idLIP8a7QhSACEySPjj/W0TL6UtE2y5zNfSoHpad8HDKGYLcJaWth6+o
rp6Ue8bfTkyo7gB2gZZXH2RgLY36ZZTf346tkcs5MM8lGMpByoqcUGPGTfd8
UkHlAb3ouJXE5vbK5hY4Kpkyx3HoRPJ4WJsKdCuYDWpj9bTQf9zFQCfyJvBs
NZGsfDyVPztY9R3u81TmvIXlgkg/HPONClFznk9mVuFfeaSMsu6htLdbITNb
G3N/bJvH5mqXqtrqnibXRpABN262Q/RoV1MojR0JS1oHsgG3sJYhn1ZyxIOH
if2V/GaGf9UlIU8kZcg/l5B71qoIhHnK/7h6LkWCToRWQbR+UjVOTuM0wiz3
yOtIf5tFe5KBZeA50xzY6Ze+huFLoE1/L/hagET8HA3z30j8t3r/q4bKNHFR
kZNgg/I4OnIu8ATtOsvrjNjCiEiZv0UD97bSpW+zLv+dyWem5F0JWCv+EZ9w
G/paEqO2JHBHIGfjMLfrsDB9Lu2smynGGQrgFA9BBXZtjJoFidqC17hzIJxN
a3oORR0Q2LtTwNIhnLV8Lhdqt+eJzOX7X/LcnvBtItsYvyVxCVS+9iQ/J7CW
k+ogyQs5wIgyliJZtBNxOReL5SJof7Q6EEhePBKGlbw0S36CsQHQMAHNga41
PJ9/9eKcVrxFsC22Mz5nwv9ca8dEc+MLFrcE/ucveNoBZU5df4Ji9gNbUIOX
Vn8ef/P89Yhw8/UJUlFJpP9m0Y6rKqjqkSYfDSBAfQ3MuIzdGVJ8l2IPvGey
3ZrrHLHiPIBxnXCWDeKvCiYgquXEF1yarHROs9CteafSjST0APYjN7a+/iYo
KYnSfOVtSQve2Nvf5s52Zu+uQBkvI5qNcPEDNSky0KX5XWZ4I2pFZ6QcwrR0
+Y9U18yxb4zOfNSmjKgcjk8xFjakhzK+QFBFUsw5tIPvNHueOeQvCJpi0ma/
PgTSdnO8S0e3Wo6afh+J2co8M6xlEDmEF3ADgcV8WI8+/EbII/CNXIk2aQJv
GyC9Edo4ogyJjZxoy1bPkNRQVClPLv891rCc0OCV2plM+ENdVPWc4C+N4+dw
yj2Ym4tG1OSNKyLxp+ND0DrBf8zEX/FKokcyzlIwbNO/4g3aCN0+k7ibx4pg
fIVoUBFWTzdVun8i6y0BWDMvl2SCNUp9tqgXk3kHsTJ8HPKr/SIKgKKv0XHY
YWXNVskNwttYxphT2eDiW6MRALmyTrl8TINzPPX67+zpz9BjNT0rsenPqamz
YXO3j7F45sPSs3bkuQOFu1GqySs+nNYkP+ktrL6rFmSwEQDLEZtUr6r9IkR7
Xcy27EMC/BTGPw1jzH3PrCujTn3Kmb7U5due0K/+gIm01q39cjyhSSVeohdt
UDqibxCbwW+AV4aWTuLXt9y4of8q/oIT0VaO+cXO2yOL6RcknKuRi0fAHKkv
hWfmqG4o4+2pel4Ou/HCTdIllnOuQPHTcUINwXrM/0ufl6lEEWynZ8OxyWaN
gC0r5xmLB4I+6WsNF6TR57uK1rc39PIvcwmDCuSJQ+4SnFDeV2F8g+MA2Bj0
3HoBl1qyVZvRXEelJmr4SbPNZ7IvpmfdrhPpHd4hNgH3mhtKElLZJBYf/BSy
6ObwTV+oaazJcG6SgltmBebwqsmnG+RZxFQ2D0LdAYallDZ1Nq/VOHfOlurr
EcUATd69SBoCTk64Jh7VBtYj5L2rZoBeKD4beznYek5VIJLE7c+v5usHjQLy
r+0fOdLBECmcZabYiQ4u2ySP2PplXl0nYUIEBcq8tuo4ELnE+YV7SDWkRGje
mksp1DUhXCH0r334qv+oUeVhoZ41Xxsk73ggX72fDZPAJ6/Guv9x+qKIvXC+
fh4GnjwxCpNjXUXUPyQWkrx3WSaW2eh+80NE343OE1JtflZYRSv5WAJSX8p7
qEKNPB9B5yB5XgpYXtY2AUhNcceTIoHqhDP96/4J9RNcZryqaRUQyMsZbjYX
qeUYQMkhRR7q80Ynj6USbi7YlU4sMTF9Jt2Xx+g0F5p7YyIjAw2oPLySTQRj
O3s3AE5QT/HjcBi8+gwpmRHPnDZ4ZPbuKLAR333enQ2IzIGI8tR0WtdFs2Vk
hb+abOcRKz3tcnB/vFzZEOPBMDcoIGXldgbGlMTnd88WVj1O6ynvYaYKqrSo
dfKhQbR6tqhgiln3Kf5aEMtXPWJXtQQDVaUxGqGT+P8NjZUD1rndmdqjqYbB
Q7Npcq4sXXhZRbsUV7UnrQb7QomZGbop6b3m1UOa13fjdeWuaVrIxeuuKjiS
Zpm7wey+20cM5J28SxEsOhompvEwMg5eMwgMqbjrAuHcP9LihjwKimKULSZ/
j0sbnTs7caKzu7I683XxDYYkLVbh2zJd5UihD5ofwDvcxgmi1JOApY2kea/o
j/CSY71Yg9X1twKLJ+8SIbNW8JsI9AO53fRJJbChTdjNuVjjfFAKQ5ch4D0t
ShDEpX21bdAZOxC9o/yygsZ6vMzpyobEsXBr/K+j1AFBiNcWEFkRhXlLQ1te
eOirZ5UrkRvgDqPMSDyfjasMX/bsPJgvBYF90+ReURq3+EQFJCugArv7qWTN
zoJbMcHZGxKe6R76yDkPNmsbTHqtyhrP/kPg+n6M0qpOj8Z3ZggZiNP6fyXr
I2w/vGbu1uBnmFI66Rd65UCzEjl+enfUzcUvxmiylRjsff0/x11QOFCCoWfQ
XFyD/G5goR/6LScDpQx0HWTuEuE/koiE7q6UdUmNLytO07vpWkVygwKLUH0L
P2yk4bW5TEyXIXOnlhBk6exSaeQNef+1VS/qBM6z2HRPXG1ONw3D/6zAXakQ
I8D6EMAa98Ml1Js0JQdPKfVuDPTEfSigpNbBBWREfc6CuaqKbf/BnPe5MEdU
dSazwXRdXhjLajmJPIwNfbMBMjMI1m89uWt0mjamiH0dodag6389ggVf/pN3
OlBbQQpZ0ew1e5ar3RVG8dGLKqpQYKOBlGtgKbp642IE0FAZ8XSlmkdIib4v
UPD8W8obhUMvoXvsQsk/w6+x+kEqz8klbeqMWZ9PZSaT5mfToi7uulioBdoy
DGgbQt4mQy8JcaaR19wFZHEJWQxHHwL1vkSa1N1iXHqq0iFAq2UF4LBK7HfX
UltPo1ap8ZrxTyqubG3lP5FtZk/18W4G65S6LS93P6TSGoMSiWBVxB0XB2Mm
/KY4z4xx8koPA68S8+84+EGDhupgSuoJ3jkgDDt5YyGqjGr/lIIwE7ExtH7L
zL9GlkAN6iVqvo48nPrcQAGTO6BWCK2r02tKdg2hZkcSbJKF86W4fvGiuUgU
5zJeqvC8YM2VS8q6vX6KBw7fybsqV2NnlGW+EWhvdUcIdRdx4onyd8gp1TL2
tO3WhIoma+1Ep6wVXrT5pAQEHx/N8V716twsupsosLJn6piJVsVxbHd104fe
fiu38qbcvU1nde5TvQMTWCvKVbsylBCXqguwEsJ+6RAA9monXfbkit6djPvx
eHHVY7FJvH4sQ1iYYIR2itJt3HuTEnFGuhJe2PwusfloHSABq1M3q/Cl/nUP
fKG95EW9/pny1fr68v/E5gngLqUcIXXwDbZ99/kZj6cwrYEXHZGE3b34v8gq
Re3DsmM9u+16UFA0TEu41/esU8zk5cpUJY4E6hBgDTgFAV+Ea4MWUBGjwqG0
ENSdX9N/Ni79DvC3fFsHm9COGy6KeS8kwZMovil+stZs11spCvEBCEY2M7hh
K4SrI5i5jFDwKA4JGGOkZjx3Wav+bkz/wG1lxJzBfBhJCFxXA8GW1Xk9n00D
D2XumxqJYg7Q+JoPjJ4JA8GW7NyGdsfR4Q8gMjFDA2GEVPoAGJ67yIhICORN
T3DlhK/BSyjTRsYUVtZphHvfq5LZTCoPQSmW/M+yTi6ETjHqMCUMXm7tx1SL
NLKtOfOtsMrK6n4tuYaO1C+kptmoBsBMBtdIEkHhJY7+OHUBGyevGMs7QytA
cIOpbMCUa6f/X6R22LrY8VA4GsrmiDt0PPuvBQEgc3qEEjI52577jxO7ATt5
BLaBA1yINmqVQyUl80Z8uNL+lMuIzUhA3kgFgfNACrQlpPHs4JstWWdhUt32
5XRExjknFBpscxkwERw+ruJyCTTd/WT8GJiFCp7U0TMQbQ83eHLgMvBIs+fd
KPe7EQ2+P8veG3TUNxNs0hK+hafQBBo3WRap2FJCFZN7vFjoQiMYaB7kO0fu
tv5h9OE4+AlRsjMspY5VNAHDDNTPuA49DaxnDEOWHmmuuX++ya4QHHWicTvt
yFtrbXziafZfQ8Ftd/vv4NgJktCIBdzxIS0TaGhRL8nDQSyBHP3zqtiUAkaR
FPm1Hu4kMKWA/h3ycziw6nR9vzyCdIkvFw8iy4br1NRVTUx619vRn0S7uvUO
kg9+HIUTnUczwWRKAUQiBK+1BqenOGu2QshL60UFwHVAdkf98LkM4BAuGcvz
gzLNrWJx8QLohwYQS6jonzhrpDCjIPzJWZ/ti4aS1aIwm6tmUwyfnGLERUI7
CjeD/fUa7OQ4j/Qdvue7v2r0tNgUMtPdm19Hz2W2sxwsmDZCvaUk/tcAj70Q
PdlW6foS4kkrKcYXgffATU+cZ5RpdpEhcenKVljtsko7NeLSe64BzWQY7yfg
cA4z2TpwhD63tg50Zr/3SJpxI5XywwQncZy+TqD4DdviAMZl2OGxL/x3TACn
yeZW3GWqseTi6SzjzDmTJoAwG72M2ztmD1zwa10MLoefTN3CUNRgTuI72y/q
cWDHg5YobC3pYKEz6y7fTJuxb1FVz2XwT1v/O0TcEHTM+v1kXMbPLKM/8WK4
kre/ChoX9WvX2pwUZ7pJR+SmyZUXWiPdo1LCAhRS6YckcvfhWgWGGkWUvC27
W1nrGSKClUy5Ld1GQMMzyYbb1vD0CsM8lql8aYDWhIufytoulCIQXZm4jPX0
TrrustmhwF7th9g3uI+P/zKpVIiXvkBXFITiwWPdWIMDAOMnyW9y5fon/dJD
s4hwBbYJQmE2KW2m3kMbzwPVvTbeoC8Zpr2AcGqVvWW7Pxc5ASEUWs76+Mj/
aMb4cGs5x6Yy+c60+jx5i1kG7qVqWjuFGAOtwYbG1O41woE32DAQXuoJgfmr
s5K1xuufpqU6AHqNU3tAck5mzcvE1zRGUCucRv+/9aHsaIiO+i/Dy7Py6k/J
OBxWYdKKUgxdiMvmc+jVhtMSC/8J1cj5wyuTXhXXH+9jdDmvVrkc7iypVnMj
hTURBm82BGuPnP9U2b2kb2lZ96NNwzHa7osQEPjzg3YM4OAk2b65+eXtADHD
gCbP9L6VXrTICZ9sezxFV+DmmA2FoyyrmVr3hyR6iqf/UzC3aq4qF3r2TGBh
aKPC6lcIQlRB2FzNgtCm6eSJkx1rtJ9LkJqbIrZfIFHuYVZ8PmvR0IMXzIyN
EjmiWG6t/w92T8dzBXengI5XEsG02K5qp8PPMAnItewzgfemThksrcR3bhmw
GZtr2SUFXQIoMUwgYnVAA+Zejwoag3ixh5eh9ooaASnGksIUANbExp5wkSdR
y5VXbwqSK7fPWt0agwa6t6zYAwJrz+4On5s046rtCd1fn5IDAwuQQCldRYkn
QBVvlR03Jv68FrC2/FOt3iTlzwOYBJVmk3sfHlmNrd1IFbRZW3DaARsoq0El
QEVmFDCDQJ+N/29OTe/HK+VYm/jlcBYeiH+FZh7w/KQ4bLjaVdDsys9D9Y5o
9pEyHuOBuy0Z2facAIIlFWw1TV9LdsKSjAudoqDPAZc8ImDuMmPYKbsBVSh/
svUHygo4wwkRtp/lx7M+FCM0hf2IwcJvWIPJg1oO5QjCRH5SYicycvgz47XL
mm2Yx5QiSzoy1V8DI5kZuMWxnMX8C0vhvbkrFqCIx5T/7XEOQcIUt6xq305G
FkU7e4V8G4Y4tgAhIAwQz1HjVHKoMVSBTF/65WTlutmeclEkCb26VM/yqxTr
r1QSlQRFeHc6ttmBeA+IGXUZ3PwjkS1qkgu1gXT4tHOeeAhurgcl8duCpcnA
iIvAwSaVy5INcKp00NjpLe1IXoOI0t8RzlLOcYlP3iSlaKDEBclCaBhocvT1
6SAocfWyEzP840GnIy6ipXWBiBrivslYvYMbNfHdeBXf90ra4H3XPpI/vgsw
B/fMLTBadmPws+bEhL6EuvMw6YEbWRkCRZORbYnEiP/EGyzK5DynX8tkye/s
pdwWK+yDhsl0/HxqENNtbkSXrjETX6p6sZ140CkGFQ6hWKoQIqnDebHplNys
+/YMOmasdkDngnduQqt4UKRM83iqlnJqI5LqsefCIiHE4aamhTEazrQM8s6m
U3fI7DC2ULJCHHDVEjRQt4QLvHQp6sXI+Vreya9IYkmVeFMfwIzOI2gwinB/
NrUREUAEpTljJ/da7r6zYVIc/ocktEbSucVb7K4i/qeWdGg4a7cKmdVw+s38
+RYIXLXegFIAOZ0XVkZVBm2F1YYUZlGpE9gTcUq4LIGosmZCMr09KaYxnlKj
N+mTc8uOyX3O5OPJQQfuxthN5v9QA/CG1Cy/pouxxWQky6t2U7pQmq8m3SPW
JGdY3RK0fTUVTEHF6kI588fx5DlTjBdSMCqs0GKV3LE94T9YS5/zGtjxiZaO
z0ydKSxKEGbjLE7Vj0WIATqSEWUmKyVblHDSdlZf4CAPZoXpA6h9xyWFnCVz
nnBrsyjf3quOK5zYntYMh+nh2DfpxXMZJIBYDtuVZvRdG2iZlq5jx2U9E/G5
+qIK/nSb4emcXMuW4NmN0oWhethdEWvjYfvgNXHdaVLZTIsKAuP7mzSkcirv
o6wPp+h2bE1enB8BxgruAd/QcK4GT+F1SZNOsI38++dQfIWpkTPkTuxZCxVZ
Gt6CNKxyMOV3v76fjUZ7jfiHNd30wTu4qdD8F+CRii/YFONNITYV2wJ7qT9Q
o/vVkXNhrJZAUrVeLmYmsLDfp2q3NQ/ZWIDOqV5Kf7/IvyN89JJAsM3SEd+g
DLyJQJTd0dbgPKaYCMtaI52RCnxjitoCWNABZ3uxXz9GnDieOC7+k/9d636u
7GnxRepEsHPl1L8+QOZ8tUi1xqye0nV3+Omgvqk+CwbR2ZsXpSrUJN+eNzMN
3Komz8IK/mw7EukiTcCtg2DHiwKlAQiDkKqIELxFd/RPmp+AtrRZ00B+c8ko
MZ21MvrnW07HfYBOgfsXL4hUJlTLBazS7rBvspWUKNGP1phH9JpgbFMXV+7p
r0IWXvA33nNIr4vu/COSzDaZF8ehhavCg2owpxyLNC22u9BILRHqXLaOLRzt
KvG8ncjQqsygIGWviePB/h6l1KTKIhET0NMP63Na6R4/QxW878tK6Q39miX5
NsnVcJeGLRh2oOEbfqtS5WNqlHiOHLdBC/mQYz8/0mxc9GGvR885/YT/shGp
rChwjBH6mde/YGjh3AUHlCdIEQcW+AamkjcGqQsT75Hau+fVayUYDZxMebbM
dBK2byLn29zMb2P0fuMQGjcdkPf1+k+BGQZ8devpnwB/OzU5iz9G1Oagolsw
Z58HnOPFsi1AodGLKf3S7mftWLSi86xX1VvNI/JLrLDvHz+AOLZTx4A04BXY
Q8F0AobCSw9cWzhkd48Sex7OKcb1OOy9UikDTm3/5pSCF++CQVdFs5imcfto
4p6Ho8JoM8tSX9Gv7QdkL1Y1R9R+Yd/g8haoUNkTaWP5zjlVOBMR3FjtdTkz
58lxsDDRUcHZICFL+NyCwZxN3QtMfAnjjQFAv2+rdJ1OOLQ3ajfLq2SN4Cuw
0WUfQCi+hJgxxLZQPQN2e0pKGskx0qLMfB4057UYcfqv6P5Fvycdbkd6BAvM
QB3kE0n0oRmTlVg8C/4DNxXbL+D38RP7lGrDeyzRAEIYgM5szrdvhHexhrOo
5cvRyYy59vOKr0TfB/vTjMta7IkT0CK1ZtU0mquIVDLLINsYvGdURhrQR0iu
aCKgGpsgS4MmR+F1D6hcy+SCA3/cCDfOuOqQ3ok312c907z4cW3CaP343/X2
edGZ7FMNj5/KCLsSBBtHpVFtsg0Hlm79NQc848cwPvtkCk03tQXIlRac0j9Y
2f2u9+FALdrbbrMYsnXk+xFsMOxBQ0rJ1CWN4BPCt/oGAhLEEn4KicHER0bi
pyovNGytWg6esK9CbR33rqGCHLJ5eOQbj98Izcg6j+0knoe9Vgn297/zmWZH
AQurTiYQhbZetS5y4p7RaYLs98eWYN6my7I7dmfmDvelPc3VVUd669YE11xb
XqJuMEo4p0Aica+1bLTa99u3K0khsn+mVFXcVOcz9TXljfiOV567MPSHYnAv
0+otBaoEtB85XEwNYeSypUdG05+cB5fryQ/5BjLSNluqNszoAdRMFU6biQlr
kYIIMeuVp8ZZVbVtZ4T7+tqvEJv0UeksBMCU+qPY+Jp+y20WKfl0hmKapaOu
ndaC446gWRbKIfjLoiAfaLEUxAKGezNV6/HPiw1nfxN0DiDdJaI/OIy7mUkK
YpQLgY8RUmMSTm57wxLct6Dq7lXo75QN5kMeJKyZhQbKKlXV+KY8NZBSCvOp
hlvFSxRt4ysxL474rtIz1TtisxZJ10kdxPo6cn2Uka/9KzyWrZm4GhVloDB0
vXrLGotCYtUrej8Q6DHOtT4WieUppyBn8x1HRZyGsOuF5VDPXjmkt6FxwcqL
0aB/ne7F6nKZ63mEUfTWahXhbvqE5E16iM4ob0Jj5VJ9i7+ETxaCseXLDM1c
GP2QIedbYdpIRsWeLAHIO5fXiYulm1McZVYA5PRwoxne5nhHHs+l23M5P4hb
w49SBZ/ZN92BsHqzmFRUqnL8B2YGUpJYO1VBPAqH3h3WBHIa8KoOme6EKZH8
5/jgBdtQRgW1j8Df4fF+OFVd9bbhQsl0qOVFc4Tq2RRn+pi5yqU7JXn8G+ib
Rq5luD9ltf8Hrk2C9/8LTeB13w4F8Cavmchrh4nJ/4hll0yay1sJvOI/n4xS
OWUnnOPca8wLDn7VBGXHnYf+35meMKjSNKnidtPGYJnjJC5yNimoKqLGB9lM
kXuZdr88PQ1DQ+DsracO52v3TL2D/Dvvjr3lsM5/cpLWt4rKwBEL/f8dD3eg
Lr3t3hmmnbCdnVscngNKZ0jacXG9LIOyBfJMXxRc0Go4hj4QDE4gDwUTcdZd
c/JURhgTzr5w+bgfQ4LG/9siyvxBtAWvePzeDuqSmtGVMZRUCQn6+5lEKaBd
qvO3jfwYfbliBK6jTaCbCAqNF4Fmv1dOgtbfocgcrBHLfg9otUCx5qNWlC7c
C54CMF89UkjZI5FpuqsQP2snE4RkMV5+Svf63bEryVulkbXEDrZ6gPF13155
CFTDvSX4PD6qATKbGnTZUcQhRU0kxigHTg3fcNqZzxmU2ueJMJIsCdomeapT
dSqdCQoRAYb79yQvGzc4OhOecxs6aHJ9uN08ZCfI0zCfg5sMtwJA+MtG1cGj
TdXeVy+UXmNT5nn0Wofk32itsHldYIkIv7WnpEDtj4BViqibd8wrHyvPZwON
kaSNWmhrQJwAJCogQX8gl/QKTNGuyQgbgHbS/jIMHOExF0iVsmSkRpDRv9Fb
NFXpaR9ZbWDKMvNlG4sKKoDdHkN2mmsxNqw22GqBX72zMHxttfn3PYXDVxkz
mxAVtPdJJggCq8YcMHMBTAEEU1Fyo5PW8PJe0S7zkKRy8xCuKYD06KqGvCJ/
ShyaEAAMLtp83EZzsPYHgt2yxOfvxETRLsR3VtDebKXgKaV8iY8bvrAh6sXh
AqObZVlPed2XtIuNEQtO9FMhVZSOX23jlGS9KBjg0Sl8LYuhMXjB7qV9y/Ht
o6JjVMVaQqsJyb4//uNmnmk0jmaek7gREhiYNNCdTFph5pgUJm/bqSskvRNe
IxUam43hCN4eRypQZPBIG0ps/xXtsC+jQnVNtFzadNU6W0rwvwCeOAVGwiv3
MojcTdKyVjfiiXl0q8G4rax4lDrytgXOqkw/jFkiGwIOpkz9F5pnONn6AA9w
hQNAqdyFozj8m21hV0ekKdmU/oW7AwK0VRouW13cnt7XMBIpij2oO+Hfwr7E
YHa4bXIIEqXhSN25yX0IvRoTAIwEOGr+YC5C/eGrZvm3TZyCOH6Mb54TI/bw
79smNUZjDiRhptBYQUMZfYvtLNPiIgiJNWa1+JFsjRroZxKe/RwBh9TPfmkH
d90xdxxjZDB/sIAplQnblLh/mK9/BfqeP2+Y+reqTxOWBk4nkcmqNWWedqYF
7ifdVfR3ZfgLD+fyv/UL66Ur7v6HNjhD0VBYpjTAjHxKMJyolzydDKTWwe2T
EQoc8bnVUJ9NCR758jLxhz1GB3X2V+Ye3MOJPQuLYCAx45/Sd0NAkSGMyVNA
CP0gjZxo3ki9DMhR6H/QIfEbs24wjvEGrSoEuIuRm+vD7E3nQeTdo89zCX44
gw4MNy8LKIdmAkOr8tfWgc4mNU5+cTAjgaVBHepRIAooW+Ekw702WnXRBC+v
OnkPikEtG1S/L7FFKBotqAc9Fg0PqDq4m71uYPk/qGOx8umeRFyEh2xbiaEX
h9rNCATYCBlvL/6U0/4jsW5rsKM1ef/lCUlCmLYMg/B6OgS0B/5ZtLv5F7ud
QANHSIKizweKZx1ER4ufKCNlavoKB8nwwcdDkWht/a6PQII9xKp2IAKtkt8d
vleNyCBni3kjSY+FseKwvviQlD84TDmy3vCyxNJoleXDDCSMSR65qiHLS4V7
NZYeLUJvtOX/NGdKzCOOO0Ks1anDgB4fKJJq42VK8SNXSERdYLok/Lsa9U5N
FoPM69XayDg0aouU+B+iPw115yYvuKM/HjkXWHZlczguRYoCY3aznR5kRWEf
DMtNpBFvuWFVoTBHMAxtH1CA0wDK6hXXc1DSK+zsod4IsF+r97Rtif20ZTJx
taUceQD03S1h9zVv7J5Rwau+pCJtKTezy4/vT6xI3eZFPSc6a7TihgcuUNbF
TPSKLDM0rywFR12hb2jkVD2xDti4NAQx9sKMZSaCuYPDIYKngF4ebVKF/R/2
5rjW73tLuLmFHB/VfWP1XLiTnEWwpJiq1mpUhvLqBxUtmom1C1HRFklZGQEG
CdI7Psk25//eb3IAKm64DuV1HoEZkOXaCRrWLCNQD2pYxqAmlW+CSRopSmxk
YKEIiNdvub8qiZ482ZN0Q+fttWyoUX5wVpzfd4oaOfg4YJdT7stZEva5GTuG
VGGt4auG6dvuUTQd1YLppMTXKyIJnbxG/Abtc4k9fANAzDL4CwGSRUmagNaR
M2876hzFpzKCFM0+knjpTNB864Jks4ULwrJ6ockrAK2NW+1vwmjyAxTcZBkJ
Esh3uiayl1xT96zrZJVY/+pfHQbb0Xt66EOmT59FRO1uF3/mRAlFwxP+jQxn
K6vZrxK68kaU0tLVnx90IZvrwoMue/YA0rligZqJWQIeKwZEbYmFaCchffFp
0iZRmAGPmVYS66oVg95jXYJhvVdPytmva3knXWNWQ9o4FP13rG363FWeJcEi
/jQ4TxuUAfYNIQ+MJ54mQFrzP/ooFJq/vdzsrMkW/P9f9iLofzcvbRyHZegS
sJpDgmnKhKojwsg9klc91n1jpinYkrFB0XfPE0qQVM+avxP/9CQg69h1G0Wu
VTUXxdwtRA1bX+9Nl6GuqzCgiUZgI6X/HDMIHW96kYIlt8oMJHgtU/jIRWtX
h4mHk4IWz6uj8HmUHwfW6BBVDu6sWCmZ+Cc6VINo+mDyYZbVczpi7jv6l5EY
9ZoiRTpETnsTdTQMtwjWHTGyLnW8lOYwYvrDxomgIljbheInxqcZz7zQ1enN
VZ8X3t2isEzgHCbVWCQTT1o31ltOgSthYOfJ27PGtY07UtYvkLY/+DhERj5E
SC0GrH54utkIyyx0vHg7FVF/1zdjXFfTco19XUYQC+MFLMhHi1OATfQQ9N1K
Z9xf80jrpGzP6UeqpJPn0zrYZwMtwniaxDTF/0LNqRye4G06H6si2ZXdDJpT
Qdq5Ru2yQFtuUg1StwJPjCx2FcRWr1UuSBGwSN3IQcPW+ZfIrrAI2dctN3bb
N1dgsvgAMtXXzbUUPu15Mf/2Ta9nTpH9Ae7Iqi1isLo9MTR7i/D4Hmjjhne8
3zaELhUNhmVyCyyNEI/ECLYsdf+peWojzuHGG1r99LDcAgqMmEuqYwowVki0
48aOtsjPJBPCDHr3cuMrjNLD3F8Ae/zjls6IBA0EuaPX4VJ94KU52jZeo71X
YY4YPDE4QudfzNJ1UTA0D6bb7FpyQF/afNY9UGxibCCnJBJ+/8M7mcJFWMUF
hN5w8g5g8YkwXaBm1ilrE5RUWkTChMQyt0bGLvPeX5VM+JDPJPeSmh/oXsk2
i3mVJASUKZcahhvgKTyYUQE0q2w1SliARaUjv8chdeEaK64mQV7gRqGZ3fBM
jIsdnj1jDO7iYZSHDlZb90kZwEikrwmacpR7kxnuHxU4stCbG3HrLGHQ9Ymc
IcwF8QtDOV7iHJDdPygcyewBnEp5iWxkQxYSQ/1ukbciDjSQ49WiPDlxw5UF
sdF+NrO9CVY3jl/eYD/61Yv2hYFeiw8A0GThvlPcLtsPPeIMwh4h9y+4RjMz
RpSUdONWms3owzsE22qNz6a8Nz+poBXwFj400vWDoVFfT3agYlrH0OS/aRgU
gcqulpT346nKRAh46FGXbAZmoUpGFGaX0qoHMTtqtPDVTHO4KHqNKvwZXAH6
5CA6I7knGzAD+6VXxuSB7BecV5BxC7+oIzixLwv4aH1/l+xyyCRaZzMDp2L/
jDtfj5YcM7GQGGlsIzPEnEh0d2pppCmnwk3ZQrc4k6DJxxzL4Gvu36om6P8U
RX1igGQfU0aY3zOVuc4PKtJ4ZKwE+ooYa8xJJBouTYLJQgq1KdLxGaBfCJ/R
fspp/JMA437solRvR/tVu86L2VqIFmBlTpAtz3GdL9Qh+Wmw7E1Cp87KZWYc
39pJ49yfAZkUzxRw+P2LPvu24r5k/Wrg9RE7BpPAELxp/7GeHaBVtZHh5pQo
RD6YbOurW7PI+lgt7aqvW5kJrE9U2EcU6FVlucg6p4m6a18mGqJFA1IG5DaW
lFhWjpYkQCv0EMvKwZ6ztV7NxSRCIW58+RTF9cMlXhvOlbhiGNRYs/CQxu5+
AHaoKs9a/Tj8MmJcg7h1sK/VXEaQ5Z0qGO7JdFs4PDtF9xlFFkx9wKnAk+14
kFcu2BNRXV28IgSig7wUULaWRlSz/iypCI5AVNLFzGbnh7lmzij8+JV6a1UX
FnDo9KkW6ElvBFbBTjyUuGZWgHQhB+oNkbLgmj+Bexz2Fi6EQ9HqsWkNSSPp
ZJO3cD1kTflR4WcoU6gimnHX+L1RkXkzsrRlbuC56we/RYVUIsx/HHPF6e+L
I6t8ZbaABjOZ1dIN8wnoXqMNg04RcXCcZuPV5IpHwTKeXoKfxrJiWkH58BTv
LeuV+94p3eh8aolJWVGYs2+81I/mAQ0P/pG7MaekM0E+uzEdKNw0cDx+uAah
OFI2QnVFYe6AnpmpBXUyoScFiNpc+2O3GvujtbL5EwBHRbW7d4FBp5/Qws2m
zinWjkYrClySJ/QKdmmomBFZvsB/fbf+QSnjvoBwEzkC+r+00gN4xRXDgSwl
sJJqfWncZPveZvFp/aAPGZkE6Bu8u5oLPGAvT8XbTE4Uhgaw6QkngTAWapbz
3nGrwKvAulPndHv8Z3xML1DcD/M2ghGCsmZMI3CT0FMmob18/G+yQqaD3GIw
/Z9IOcE9EDx6cperSC4DiDcNBXASFD5/CYgICHwn5XjgFJUnZD45m8C7n66s
l8jijq1EfxgBzUv08/7rb9IwFxp1DYGpcg/u/o/7GjvPFkSEJgThpmfGmrSk
aN9lq2M4sZbJTM0yhq0LuHzOXfMczxquvKYCD2HK6WLQ5p5VH+Tw74kN7IUk
IXLELxHnyExss2RoTvBhewejnx5S2ex+jS0eKrcARphG9/Rw2zMeDpn0nbfK
62SuVY532sElb5Zvq5YdG53Z94A4D9gLAJHv6Hmc+ozhxurQUraUrT/wMnsP
Q0iQVnlXfotpAk5oxBlkS7bQKE7kyC9OaTxdVpusUC4u8k/6MFu8GTlrDLoz
sjb4ZJhrn+M28ZohrH8VmEXdNKcvQbHhCxFQ9DCyDjg8yHjSLxi7IWotYF3I
3pWSYtHEiQl5f5v7hhtcequbozzYIT6hKWNc1ex1TNvz8TfxeDHyzUPVRDL1
gKLrlgyG9fmPNhsv08i4ly47ur3fAIEBeMNAqhDQvbbausSzjNxubYUws6+D
fSTQFm8/gZRFni0LKeiydIt4P3MWHaXnN4zWmTcUMWLyiPxKZZjzD2AB1i2+
AxpD6b6zYsKFrhlbRYhxZxierxEmTte8sO7L0p2DrK3B6KmCZF8j/xm2ioPm
Pzc69s6NybgZtcpvYEQ3oBv3ZLkWjOSgsqYODUi9K6RKbWTKILnQQgKe/NLc
SzyE+G4fB5ZStWE1ZxpQM2ZvHFkW7z/b5h55cNMEm2yzf7YZdpoF7zchr4o5
IxQL1l5PSRtJsO6I96bqcfgj8hnQPcqcaUFB0gv46Att2ZKG3qmhR9Spzrha
gTMsOxjTyzXYXS7yaH9JjEpHVRvCJwjPZ2aTg87dRRQ16hF0cTFiff1BhxOv
kbh1qeU1SXOaLqJ2AkVfOv33OUcs3WFg0j/mnxsCEpaYw72ww9dv6e6UJXuo
jAV3sSo2Hr44ur1EOPhyZpZW9MiXgiK1D+btEgriMSDMEkfRlRwWW5zErrJj
Xyr5kZJStfygi5N3hDKuvY1Y0PSuiMiz79V//Waui9VzEBqJ7EuuSZ3lhq9M
74k0GSnCuO+fAE4DNyiMRSwrDr1SVUfeJK4GBHEvbQ0uCNdv4A7HbvlUt7Oj
AixEyHPymlrClmhfMFW9YIDYxFMrEf1b9lVBsv9ff6UK4wEsLsMAAfX/QITL
xzYGIOLdxjWC0gu++FbghXdqvU3vf+Cd6yj6/tLjZf0WChtF/iO2OlUNI3yy
lnI0qwv9sV7vBsEIUzBhFEtlAaFUoaWu7lNwBZPlhMkd97nSAIzzxnBnUmu5
GAQNy+XbM6SA1L0RpSW5EoYS26aEjowIMjGi/sogKlV9xvT4fRZqYCW6aq10
hQmzWDD0qetM8Fb5OCe7KcEBwwXc/K2qHaht8THb0yIxdQOaZO4VoL/4IEpm
95ibJ+SopF6uc5JuzG/SaeV4CUKIlR8g7kocl4AXP2CEoCH8zdgo5GNbG0km
K4+LsEHtWVtu0tD5bklLQgCFct5z7OAxZ9ACARCIAlrmP+KroRCrxictXxWB
JGfcADz1fOP6ktcuJLwvHOpfmxrv7l+KKBAnblTXP6diV9AnTSD8+eyXLoVJ
XOpZX+CebQZx1p9XTeL87Lw4yyqpQi1Mox/+48Rq1YzI5FbD6f5yA323V9Of
Xyi9V+5Syqjzmzzjk41gDHpEzmdyU+Ou2EpBGNyFhhPeFL+wwA+Rh/u7WRAp
LpAHhAwVDunBsasgjZ0NzMALwrKOQaGXSzqZkm95vAlfdaoPnPX+OKD8qm78
8v/67DmFXPzeONX9TNwJoYKRMMsPYAHasSjTX1L6ScUL9naxgNAF5lDISZuq
6a4tUpOcfjv0ykOfPn0vsC8r5hfM3wLsdnajEynnyVUbbuWhJO62PX1MSHuK
dPXXqnhyTQW4vE8SI9Xl5D0+eTNgCQ4sVDSyVBSGuI0dF8R/Q9a/QhYPPjK5
nNBDJ/I2YDjkhPZfEu387jn4XsGTQQETrmkiMEtoU/9Mwq8V82zahEE+rM8X
Cl6hs6QAZVk0vQnJ2P96l5AVS+U47x6PioGCH2Xx5ijfMtRR2AysblLGepio
q6ge0kmzTXNmbxovS/hlRwfOMj9GffaqJIWTTqlPcn2iT+vjT5567D4fUoft
dVWNjxUHNQpx6W0HAnk9yykXlEpGZpr4zlKOEJKG0tEl9vcyc70o51L7c7Co
eNMTAvImrKddxSXdTVLqbgppOLfQ8Pod8rRwRucRUCGbvufjXaXnAUdlhn3U
D0/ofU1UFzzMtIpJlE8tVLMsz+zsLEBUahukF5Cf9Rm0Ww8kd1/xHloHG9Jq
E4MjEifIWp84izEPWh+wNXYk/wS7LvXFGtjQ0m9xeaDpFfsZHB23y0fNMgaI
9NBcXWAYQ5LVAa/7Akos9eRK1eMrMNRA6sxjvcYJXyITdWwv5P8Eb8OdcjuV
Z+KhwQ3Hq4YPZOGbk+Kr7MilU+DFFRbnFpaG/oNGBPb4h8EYnlbnCMb64NnR
xUJ95tpX9F/wSLpfSNuE31nptJX6RzlNuq5Fzqqaw8Etd775HKIO0NW7LIfV
S9CrrsrzWSrApxaBCjYsLsHznMh8D+i2bbO1Sm3hOk1ue6bl7x0e6u1VORSz
UVf5Vilwh7l87nsckRXBlzmSOMfdJ4KytTUgf/uykaLuJ/o+7zquXwh1odPy
o1y6Cvv2Bevx7hQi3UqygTepc3HATGaVWc96Ev3V+1ShjBA0cvrStKJeFxUU
U3ICNYIqc+m2K22cWzZbkyk+eo3U/XiyN83rGQPImEE+sQNFqlfmPu5y+rJP
PeX/ClNSqpM/jOJjfB6BJgr1y85/HkruBf0XCjA61Zmo/GeDHKVfPOTq/q/J
fpGqHCg8aG87vhc2huOzxsoTGg0aa4POwn9Fkeocx5alNGxVXrnotyKT4U5k
vLTl38PfMVnOUIJwrP46reruFnLSKO1o6Oq4THo8UP/SamCNFnLK3ALIWYuc
lAlfu9xPL25U8zp8kJ1TTL7IYlKepg7H9v4M96XdA4fBZWDZ2g/cb0nyKRuL
YuVwegeGgLfaZ25J7d+9u1XE15ULoOZtJ0YNjrTYaB+sb5+a+cqs4e83Yob9
zX+KNE7WpmOuz4Yj8q7GU7aHMBqo+oekii6GqGtzC+OzUhYAQI4egftfFZUE
f1vV2hUCQe4no6enPfmDPuD4eaKnOn75Rm5CM1Be6+yNFJFH1Qal7GgmyOj/
zuRBqiCreuoXdMoeGvoo4nj5i5BQCSAIXoFRxPDzSW0Si4uWeYvjgC1vKA3y
AiozLUYAITTnYmmZUg/40Rszk6YJjK0QHsc4tVRVuMSFdo7rz+3m2MOmltxa
xng9G/uEnLTUD5yYfm3dyN3Kg7KsHaZB9tVkPDw3pY0FTSmaIDrAtYE8tG4E
JuUs7Sm5/ou05vHg

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeieC+bakXCxZCdUz8JsAjcVX4ajoIut0IYCHsHxbgdPY0SoOD0UnA2HoOYgLoDF+OlIvCu5fg32HKINM6pR0QQI0CoTJH43GY9K4wFEhNIhrO2tZW58k2E7e0fSzD11B0jxJkVWM4oTnnOzq0W8R1oA5aKRcznlkwq9SFRYYVnFZoylIjywHnhRndE2b4xlUzERky6tUg12CXWAQdw83ptfiH1zykv3CyWxNLgW82XBjH/Jkrj7EYIlx+wAdt9DE2VByqDzNzgB/IcS0ZccX21rbGyjk19+g/+ESHShgSxHaSqrpB9gaiBeVk0CgKU65sHfGAgYjfdmeZ6Iz6Z4xbHhzlkq032e+zmmkEwqjixTeFAxAg4wOQ489OkqaX4mlBID+wUhT08FdTSm6lRpQM4orYUhG2DFLVuOTCWXaf/4GTY44z96DZkM29J78uCTSqps047HwJr2CKqCVCl2zrKqLWLCiA2k8/jaRtzDjVhaQY27ag1rYdVF/OHKbp8TSh8O67lhHk/tZSGKc6L4fEl9m6a414zil/8mBmYWvRv2wg9NpVpLEriXv9hOlp3q24RTGdf0JZuUgO4EY/EtLJSV6hql6CTvwmIZeQbIjHkIF/3mjS3wY+D5834CbJLHWs5bT4fTPI5HTcUBXD03jWhnStTTPPkxxhozmJbLR9YS3I6eYOqZHBAeOl5uVdEZOWbPcvzzME3yiUqrwmzJquTKPutbPmaRYHymPsdAlsJiyWScghlPOE5Onf1+nV3A8b165gM+xYpjJ3czSYEuhRMJ"
`endif