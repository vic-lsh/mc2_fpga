// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iM/mpnyyFi7aAWYcFLnSm9jD4sIjoGApek/PrnnyQ82+Dp4RMwsqhS8vxvI7
xg3rh/GjnlDK+4dYrK1zLi45Q+by67ViroSKhL7kmX6U2MUqVn3brCK3/JKR
mD4EaaI4TE0JJNZF69pZY6k+Kay0c+FULvtWZLdPfsUCM05zjieM+qQlC7e3
kVAlxp5XqfGmUD74pJT77JRSKG737aoo2Li+hLXowLXOCrO3HXton3GO8I9a
HrslCyxJPbbXbgOcxS6Rqn/XBxqwp0llwDdjMO6H6TTGg6oYlMKNSyL7Gx10
Pd7ovKxzJYVWv/fRYTxrN1vgV3IyLcmvnr/BE34a6A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dibrT5zxdq7OPGBnHxGg0wvJj0FD6S/49all5v2uR/jmJzkvCawXXQssX2HC
5z520w25LMNUePuM6FJ8XAidfHsvyzCM8WS9n96zFrFY0cNR0K5aKI50kuVU
hQapTkOjCo8+ueGBu29myCTv0rCn9wswHNScAvZO4FtgJo02QlcoVFBcPZTB
y8fgiuHcEgemZpbCSwJZBgqGs/HKSeB9Q73xH5BfTFHIT23CwW5UmupcJ6CW
KliKJ9nyP3Nsmn9Gx46eiuv6TMRaaoNoG9kZkpNM3EYxtKhrOFDmxmXEvSM4
yEi5gQvNi69Y1sL9A/U/6r2CPuWS56/3HJ0HxDHtog==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tDyScgQrV3xnE9WNJrLRYfXUXc/cnDMHJoJ7pzj1hGLB5sJfWRGLlJyVU/bk
zC0fTb/yuklOGEXOAQTRhvQXpWz6rXLClLYWFxmfprN8IF7Ceyngkmk+OZlG
ETei8Qbyp5f71mhG7frBamoDfkWUKHGrgm9wVeohm+9yeJfhMNFnvwv94K7c
4skH+zNHWld3MaIw09xp8193z/REUAO5B9fNkIyXr7ieiP+PLhtlyBO/MCMV
Ibpj74TDrCl9Px3qBuNJVVdnol9huM3lEDMFMo+WBEPUgUwwTXxAdYVOE/gX
zdmU7vzVvofWELL8xn6tyharjmkWp0nePYw3aN3BZA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QsQ0lTc1q8sy+qcAEOza+yQnr7+Hn/MWUI8UkE7B8j4QyUZB0dyRj667rrAc
7MYxg3GwIPQC+5Y+WKtOHrvT/BhnCxZyKVrTuy2dZVDil5H7zH2v3yRP5Gg5
SZQ1oH09xDwGN0F6SY9fyCfne8AU8F8XtroDYT2Cm17az2gUHyQ5Pw6x/0ys
sN308eVYvQu5wcP6RXRb8E+W/oruoDIKG/bFwuIAF+d1aQS1yEPYHmbeDoX/
9ibGW52am5XbMv4GBVSIRn7YMjIlzEI0DE0Pd8IAwPS1VbsbCgljlUHfOZD/
l/Bg4BzEBVRR7Hzdki+kMbpQGah4luIpWD8hzAmy4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TIlffLn0dyRXpUd7kUL9qu9IBwUgfvL85yFtO8t2hvfGmz3O3GEvZf59ejMq
9iusy1VWTFW8Tqe5Sl5hqpGBmf2huajz+pLrByXfcY48MdZR4rgGf8s8nXUR
N4SXbz0APjekoq6X6f+pHev0n5zFl+cPESlOAw8iZVYIufKwbiE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Dul9jmVEqPtTB3jMze4D8SrTZLHBzl0422svMH+L9kULUgrllgMGLqjhoBwI
O2vVnHfH7UCabJupRSzDi4RpnPhY+y49tOac/ODvNHAfUECHWoZbPM4lE7MG
igGokJ2f6fYCJA8Pqo2A8hMwjiDLWbpL2FxWeTuXiY9c+WvJsqx6nsurgQbu
d5ru6ZEt6Z4YC6S988Yq+F/Ykhv1LPOCbK0sKBorz9aHXkLZjXObS8y7WJyb
FVCXRsGsKYXwKQoANuhzTsvHQ5MtAMwUr9sb139TdiHtxJ2hDzs0wUIS3KCr
Ws5kBgXiJjxar0Dvq4yaV+Dl8/fcuM0U/4vrizulXlWaRajs6cn09bf/Sjd7
aqvijF6tR/npI33kD8ZNM4JjK/rtMh8dPtwUjnuXvAymgopmEvggppyywIfn
2nIuEMXwSrEFqIT7PGJlxZKEZ+0zqc3adzX1NFWYWba/wmgKSAOswNR6GAkl
u96YsTqouaKziaFFiPyrKry1ErpYsn7j


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XmeyWSF4yfu8WMNcVDq6TaQww4+iUAUeIG+qbjUtUKk35Swo2udqPAqHVqyF
Xs3SInluwC9kXkvgCr+kToByjd5/onfdUUwJnoqySW8m3fiW8iuH0TaE1QIG
w0XQdbHGavVfUDqeHVae0SmrxoTAJ9U1CM3Z5lac1+1ryqga6XI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J4soRPWg0BreFj44hKUSLeUUjLzjTGBPxdeyMh3UtRRRZ0Rn2XSF/jYPIE6x
KfgErL/aKTcJIkEndda4e0I7eFzspSbpQSzZvJ/46Ng5t382xAPNygmgRqVv
Xj/Tz6rNIaLgOIj8SaX8CGWdIuD7gPwfd9xe6/gfXklrgHnS2bI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1424)
`pragma protect data_block
aiMlnN/NYlhQZBr81cOReHSlPyi9obUWuiKHMJRtREqakuzwAHRLkrayZqDt
3RNFFae6+BQGIs5w4/JKRDH2N3evgsg2XkGggchgNWi0iFojN66V1Sk8L4dt
EzPJBfB49CiJ1/nvMa4jgBJx23e/TGWgAEZuS7KksR1FeBmss4PSHODvORQX
PnhcpJAg9H7N8Xjcl6uTSSlcKEFYhlCeEUCO4HkZ0eBFsuAXZRObkczrpkWf
fTd2B94rXRtxlBpKII+5SMaa5Qw9Lhy1nNKKciUxGj0zhSQghaha+h7Z3vaC
HkIBep8s6enlWXfj2Xrn40aSvrOTZ6u+trrNHYOGO9i+RMZHSeHRvUgxu7mX
mP2sJefM0j3r+ynnohWj/ZRNHO7mQY2Og7QqgEP0W7sHXbr5motaWEXxybEQ
FmDzKgXuphjQACVYOOyidnJEKp3693fltaKe7AD4R2zDyGxK2G1070Ot3VR3
cpSZ/d0QGmMJgcIYdmi0Nj6tYUkTV/C0J97z87YcUKNJIaZ2cRh7Fd2L5hxF
vcDt1OtcDoiOaAJicrsrwL+jTQtONquW+4nYMBni/LwSZpjWjrFtpoFRWrK1
vyBgOHdkoM0syWpO790mR2egl4PkgiqMVkQnBrpWtdqk7LnJp4A8RzBtUfDy
GQ1Y+t6mGn7HIZcSvdo0Kvt+lPDnmpbmSzvl+4ND9L7lgnhwa2yVYSUT3uOI
T/tgLaHn5GqI+Z68FHv1AdtO/l6k2mUI23coV51mr3dYO84itv1OxNH6ZzPm
GYgwXPxjUz3cu0ALJY930cr6encXSwC6nAQSb+ysgomSmZsiQ+EnA9p3ccKp
5lSQeTsU2RK9a7BZcZ6k3NscfxmfodrOobY8BERMn6UrZGtaS5Roh5Nnx4Vt
s/zDircpYsynAtfTlgS/YuxkoJ/uCLwMHz09+7g7jgGcInXA9qyPVdMhgaqJ
cfj1WOyoQ+Qd5OePDrPqcsiUL6JDi/et1mwbfYR5Y76PMuZcWeE9WFxcUgZ1
01ZgTY7WEkZSsGXSFotPqIU3CplI79NIvU0cRto0OEzWFx75KRi/k/DuUKne
p/2ff8chZY8jEwfGx2AnaMoSvUyFc4cs23J2RRUmING4jBhMBoUK6bDSgyoA
7IDgXxoyQ/MMDQIzIYA3FlU4B6HLhjtWk/BYzBfNSdbVTuxw9uBVUF6eXNK9
QKwHC5z44jM2GMrB4TmV6sIyvf4rI7ELuOCiwxdM85wZ5hUf511RRVETfrXE
Q6BFSY7kJYFmjWC1K7IkY3AdNsMeca6daLpJ74GSQfkjYgyrkJc/VSW+0TWP
0bYZLAVMd5WjwFYWJ8zG214scTOVNIGKKk5xDC/ry+NuvewBBPgUIOZXilpG
m7w4QbyZ6h4iiV7ljWG+RKFmm6hENq8S2wDMxUkdzW/BMS5cWMfaW7WVAvI6
/8BXewXOLhKoBo244C+zFhpqI7HBILzB39nyo7P/T+xN0C495Wml4kjEBkuT
HRndkZUXuqR2ejOSTyxDLQYTZD1VlwIdYCV6YeIuBRuxGMwKN6dfI2e1Mntx
hpu8aCKUDy0j7OU6HXBUbU6l182Ru7LwKRgk6hCuvAfk2hnDHlqOBx8cPDo/
zmZBdPRF98K7xgRh36ANo9BEYnglGI5151v4n6llIdwZ5BuNC8mpb+Q9iAwA
YOdWPrRYwg7ZNmuf7AFxA0moaw3m8AKTcpcpGtNSBlAk1T4jOwApGefEX70S
X5NmBoJXNLwqEpZRF0IEK5uZVldVN7YbmtrwCNYyRSehCZJ8P7g9GzPn8OcJ
XrS5vbdHTrFloGQQHpDXKxZUfsCvKCiypBOON1xaR4r8LMndlwPH73LYHo2Q
/oIJOQYRJ3ceYGsdLxs9czUl7lBpIYtJ8IinfTk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQowC7VynDAXpHhHULTYSJjMvw58pxYe3WVxmJHwv7MbkJ6PJoFvzZS1U/Ap1whJOIiOdzhmGV+foE8ze8vqsgmvNbal9sUvgwg0uOfOFk8jfWKiQTXlsofNReVbW8PqYV5D+zs+Uv60wpe++SP1Ew+SCbxpe69ovWYZUMXiyX+2Pu51sLLeOtgKtw9CQnMNUKVBymvkfOFaDnFwMNfcQwROc0m1CZUu+gzh9Tx98NCVC8lQpqixESrLpitQzzBDPLBxti+9xxOq84GAW29kq6YsfB4aF2O8F4hgxyAS2ZDT+LERlrF64MnEnhBvrYGCffPPx+ChWZNnMauALs0+Gv/5sI+iJg6nbLRMpTGCZTCDO9ef4OTiyu3DUb1ZQ54lCG79j8SAyjc3svywIWiLzM4s8dSR7Sy+pwR29PI2Krgy2NKEQ++sv82cgSljqdWf9XvRaXLi63TVdBQXodxgDqa05AMbD4l3L/CNv6J4eWMx/hjt8cdKzVQJFI5pZbvjdECCOcyBjFlaE0zXake0/P5uM0rqJR63c+T6KEYJiJcWzO/KLQtyxlY96tbSHLvbBmeYkgDv9kAArWNnotDR3wdCr/zdlD0E03m9yWM5G/FBPjUi+6FqcwD5TGLmpDK3ncpWRKJJXweTeGxcBe7K9bSIaYfImfs/I0UfqlcPxh00ZoURlOQX2t7zNTPbl9utGQoG5Icdz7oz+cgxV5HSQoxtR3wuQm5ekO7b2mbnoBCLPkH1o2s13tVmed+lG0aSOu9dbYMgH91KKm6F/AKyi24jO"
`endif