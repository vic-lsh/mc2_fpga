// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R9k7pErL1XJFY9sJeDTEtvKfyCR5QnIfgD58qJdKoG9MwJwQGNlIn3GITXgb
3DO0YQ51X9nwk0pAPRuwhMLdAyY/Ix0p1DcK4lN2zrQFidLHLL25AgTNbv3w
FkDMN/nNDyLHTc2JEB1CgZg612VT76/OEZBwc5+pPLWCCACXkicGLiTjb5oh
peFqG5IJi7hRd3EN6z48WWjKZNsTWmJf8Qcv4GJkoAMiVlyEzFE2sDCBi6+l
mgwVNOZfTzGVNEbGoiG0vI1Pk+5qy5F7Chk2ptNHOk3Ct4DrscKv/1aMaQ8f
el7FjAW2Y/4vSmZQ9iJoW4cDCZLdDgyIe5E+9gvS4Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QoJd1VgqC5QBkFwC9rEaB0HuBriyedf1HMY6GRogC0t/IbKRTnrxYDG9zJR+
iU/M5epj0vSJYa+Fh1GEbWk90rpqFxxa2w6NzDKzgXgU9u4rUH4VAa5zGgeY
f7MADPKKn6hZ5BeSpb6BzlRL3aGfty8pCVDXB7L0JiCICHO8cSkozcfq7TNA
2h5cO8Wy2tpPF1GrIZoFqrybBDgmjFAauLwhCwd27mBxR1yV0Z/zwB32cb4Y
q7JEXOuci+fVnDoClwTGbzf1h4TYUeq0UC4gmmzL5MjFA/DD+MP/E/yXamxm
kDZqvhMrJQRxtaTrnN25Qmj8qy3weUaiLP+2QpREdg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lw4xo0JYwPenC7fYUudiEZRotSKSveCmnABOUVLyjQby76HEveW00IY+06DO
pSY4PBtyNEU01w199ODsih7dFO4b3hDaQjm32fnszMpqlAp+Zt+Im8zyEBNU
+1aJLFU9EsyQtAbKpIM74JmSkU8d8jkQ0WQ/UVhGSL4iK/1zm3nMhlT8M4co
NKPP0rkxGw+G7rPWNNkdITDhK9GeFuSh4OerPkBxrpM1mSjJJohuybL6NT9/
WPvpBIy9j64wQsuQITiEM9zfELD4sAYzJQNN/f3FqLDNp9a5LK/vZdYx8hge
tInhTKw4Pd0TtzVCGdEg25WbsXbnu4ZWtmqhPF5P7A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Kz9DU2MDlQm/Ql4K88CwAsx76XiTOFyz42qdUgUpPQAsJrySUnJLxklLHWq8
HJo4TWnPh7pOtKppQbl4ru0H9Q1J5gYfzlrEvQixGG3tgBj8BpTtrMMwEo0g
BbTApAA/B86clzNRhG3ea4s2R5tpvl4t5JNvxWaj4KeRXk+C1Y0yW6G9/4qC
IItWVEDn0qyT+73pI78e26oa+P21jXNvy8hZNHj0EVIw4ooU2zfjoJWhnupT
FcT0L2iZW2hSbBsWE7qb0tXam21+mtheCaibQpP0vDPIrDltL6I0b6cR+yEi
d8vy8jH61kQxITMqqu2ybuTBROd5ALDb/U54qnJlrw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GtyYx8+VA5BkeZ/vUXfliMCrq0+Z5SThHoaFb5ZIrJh3j6xhQ8z80OXPfzni
+8EJupVxg7A1jNipliXDw9wlz6aHsk4iCr+AHdtygBA98RLtIvi7x6nJab3A
NcRRVNuEQx9rNf8nS1Zj9RVlqimgvKSs7Mv/PvRYWUKJpwJNJpM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ObcctJVvBUMqyVTHKhvK5uZvrT7OOBeRkjp1Jgnj22Sxmq0e9Os+w6VemF/v
kV6Nq6fMjlKwZgzm0H1CNjZnbD4S2Lcz9nqazFR+hHJx3EW211zKtIIp4bF1
fsgxKfte9ZNtsIyCWavcQFtedHMpX+l37udKkiLrQQwxeNAxwbBGAldtZd5y
6PqN8iWMo6Pq0iS4HLEQq/VpnYWOBxBEiEbKIeQEO5URwjipse0GAynxNlGT
K94PDbeRNTEvfRZ6ZULkSyLohAZc4utDKiEP1xeTJC9SGz5j0ddPUurtl1vx
HuEJ3pQzBZG50g9QrUibOUW2Tm/QFEkEj2d9K8uSrDe/AF3Fkothv6vqdDC/
hhdbRxC8Ci6QK9r/pp6PwPTPbPOe+EtXeMgmZDOeRaQJ8i6bAQp4gj1HmmYU
IfINVE6cuzP9lFi1nMDweuG7KA3gOX59NUP3ZGkGoz00FccnhGGztk5IU+t9
Nii/SyYU9bNrYNZ9BaTBBURs/GZwFzAr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
spdBfyFjuyVVKw87J5GkEyj88tjIP3iPryEhCHhY/W4Cxe8ibBl0CXNyECTt
6qR9MBG/zTzLorw8vpjYcK8oMMQQUWVGgrzP1elY3YQFgm60TcgeLNhG6GWD
tDsP5ZPQZ58g+R2y20nViURy0Z59fKV6bhzZUFAX7OMJoEE6bUU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AF/NbQs9Gr5KY1Ic7Un0SPsq1Rlf1QlhWP1BNnzxFr4P6krp0JQBpzYxwLWt
xOsrqPxnFYD6cB7yUGb4d94tOtqVakWnNECCRJ/rb4m+vA+T48T5tr4BJ7/P
lGX6O7w8/DP4TnDZKubGXSjTDpMOfMFtpdpK0YzCnDVyU90IUMA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18704)
`pragma protect data_block
7XJXXMf6N11eYdy97FLXMj/LTeq4PiFQ1d4sVxcZfxmjw8dSXIb5wk3+amd8
sbXRr7gWcKKNdq7eADcgGXhwGKXJEZMUykC6aWBLXOz7B5BephcRbcQpxF+N
toSZe1MgTlPIAz3JSuqjvU00sah6Y9hxBYX+it6rL5J/OZIUSV3np2IyZRC/
Ow7pDphKJy5QjoYY2OVF2SawPj3dkKKQEZthiXl/eA4Lr/Dmh2QSilvc2JP4
3J93U3OB6z72HvdyeHQ/he6R6GaqHzo3RL9OG2vDK2smD2R1xlMKagR6ZZcq
MeMr19RISpktwO99BIy12+zLaBgumeEu3X/P/XynULNpF3BV3osWEFT+bfvI
s4rUCh/7ckGkEvrk7G5fVijBaxzubGNhSdurfQmhe1J+eDFocuLxbnKP9wpK
mL2mAxM3R+Ewjf2fhIuHYMKpepsylx3T3J2qimrA28OFM7Zpz1Q3eXvj0xbM
nzGZpYb2c+OdWCkcIJRcHUCqAbrK/y6rNPIXsDt5wCeWQUr3Dmm2hwfblb9d
jHK7kl2Wu3tqScFJXo1+B0NNO+MR1ghvdi5iX0BKjMjoKwJ51OYilBbeSmxt
w6JnppqpN0P+kw8r4QkiK38Armen4km3L2lVutlCt9/H6vckxJvBbjirSjpQ
KfNDDvKSrXbv98CADxrq+3v1n/qlvImlU7HDGq00SzKqjGd8AASrNxvdL7Cq
KWr2AiH6NNrpGQh/HbJBlnV88yiUoRn0pHbdrRaVPdRmEMkhZi6mZS0GC71A
Nr06gEeRK0Ix2v168s3xJyOSrpyzMLGdJCmjY+hUDvSs7A+lrTLypyFuLB+4
UnGZyKajrm6AbFzfVf2zi9j/oJrrcD88RDp1vaHKjbFMJC+SHCIHnfRtRGTZ
aeRcaFrIccu/ROR1udYvPbIY9VR8EUj6k75xQMQ5xiiN2etM+fkrtqYpIB88
IxuG66wm/VPQGXTsVSNInM7Jz3OFsu8m2sL3E7VoDpx3QI68EKr06DXrEmCL
AHvztBdH0ONU95b0N8VPYjEFcZvppYmg5uVBucSVv36dL7ClG9wBXOnBOZIp
heTVTPHYbskqnGP4meYEMRl6x2UEfrGwRkDLc58K7ruYKJdxAXqU2qPU2p3a
JKQMQwPx5F9xb8GCqv4PKn58cDvtrypwH478S1pqHxCTMDAjac6n5SkR5UXo
R9cAI+AkRco+fbdmoRwZgVZO4gM7EpLRDSDA7uwn9zF6DDj1ZzYJYNH4ExX6
BKOeYbg2JhAyLhZy+/GE82Ti9uuDab/3hXf95LmfZDsvNuNHPaBpib7jCF8C
NeAy8114RJENZU4BpAQeyF3pqk6YkVmdznrRNyKQPoxVRWiIG6RM8Zhg207V
CSpjaK+jXqLixT/ixoIo0ZcMJr9v9w5QEMpPPcFYdaJMswcRyZAo/ebaaIqc
HjVxgLb0Yn+AlEqWWVqYdI7nqS38bDPzUYfWgzb44AMW8+LsndGuNyA2i7xZ
twOmimzzb5StalcA1aJhlY3PRPOyjFlt6LnR/qXKC3QU91VWMmvt77QNgKA6
2WHZSItq7U3tSez8MkjCWhjmvcV6MFFr7JTA1Kb3JItYyX56kTdCJ2JHh1Ca
XRpMWxpe/oZzLh/XEvHkYGt2y7H2S21XNqYuk4gTBakNSNrK/eYjwFOipo3Q
nt/JJxyb/FmAl6AfTUlZK2Ds6LsNcMpqQNUI/+QilhZQxdojGq3+BCF67fAv
R4Fo0m+7Nt8p7c/+VAu+WTm5Bwwa0UVTkMWyGc+oAv7Q+fq7JvCzB+Hc75Vg
ekauUoIaReN1Lv1xkzLKDWKFDJad9+43s/VROQE2OmSgIe7wLRKukd8kBjNl
36QUcgJLUT/0W+utaBK6AHbpLnkFMSwBtHFREfCbhEtp4BxsL72Q7t8OTL6q
yPrYIzSGzGidimNrbVbuuzaHHB+NRtMSSYsu4Ojd5bUz0R+bxQRm4NypSFUw
z9hDQuzIRlRbRp2y6FL5h/VZdWw/PXm+ilXkpomhNy4YR5Kke/ogjz2TwHLh
wBA08v08VyZWDgRReXNjF+qfHBCWfkrYTwXBeFHHLepUJJM45iunxKMmEjVg
abRbTxYmWiSIOuFlq3XNoCllpc/sWJuFegV2l9yB25CNqd/cgwmcXIF7mlnY
tF4a7LAyL+Dqoa6ccy9+d57KbMWV5PSSMEx8J0J8f0rmA2jEQB1QXDnqK6RL
Rbz7uf38kyHQuouBaTsWqew/cvw8M5n8FVCw3uXPxm+8BeOafedpnGv9TrCH
oJGnkzNAqp41KmuAjO5mnGA9onSOoM8oH19IYNZvwUwerPIbd+XcXkA39vwe
FzRO3APx18H1DRHmHaAb9a5AqOMFlf8B49jNRAFVJS5QVVpSWRJOsyGQoCd7
AjI0g3/w/hTvBqvECfbtNOH5pJBNO1I9e0QQrkdzsyRcLkb3u4IGBl8QlIjM
ycXKrcHTHsqneyt0Yn2q9bMtu7oTwtLYRSYXepqxG5I1lin3V2NvJjMAeoA7
cCWMP7A4vH6gVkH+H205Gp5DL8c6O/p1y8pvjy1EIab3eWzsLnHwkU2S8x+5
yVvFwBceWkLUDHthm2FvWUAZ0mmq5lazF/SXFBwxfKZFVyApuUahSX/COr09
c7ZbMw+HL3jAuQggHk0gPIU63XUIKzjac/qYReSTg+CJn6NP63kEefPGgk7l
HT5cXucPVRJfKA4TG01/eftFW74uQjbsSL8eD/6PYlEuvtk4/FikIX3hxSNQ
gQ4m2qDrHfajK2auUfKbJl2Ah4aQZlVeFj7w9XFWgUOUvJHSLXE0av7Bqqgm
STsqrC6WSgJJnYJR25Cv/0pK/molAgLJaCdDeY+Bs9wp3WkKKQ6fQqNHQDY1
yREwnJcV6KNxwK+TFcbUaylrWCX2ghJe1C/hNn/5x0sjXYkRqH8wN766j9X3
VwycWd6XUPpQRlj4Odn9S0YaeFaywe+8RX3+vF/Vhd7kvC0RooVG1hPEDf9q
WvsJ4knRupKtM5+r5Gi/PJCNnzRX9jHWb4zgq8idJoJMHRBaP7muNHuQnP/L
nSUY62VUV/7UQtG3Io3v4E0QScOYYRfSWLqkUFEfmyBkIgkXeGYnR4xpv2c0
iQjCO7+B1/alo0XJisH3wbZGv8T0LnZ1O6e/kA4/MC3FXfGWsIP55jEJoF1q
N3T7GC02eM/N12o2p9XRbDKoYZ+h68w+yqChWbXKbe0emP6IcK7R8FROK9ln
p70CAFTsJJZOkdNqVMCQuf21IuPL2mwsDw1Y4BMRmC2ov0dMePLkIte1MM2e
Y+jJ/HpqMjDSBmMT95EJFr3jYWiKCCM+wKmVyYXNoWgjAfJCAEfQ5K6B0vMS
m6X+QJ5lW7ixUFzPX0I/vt7wSIZ1aPO80LieLr3K6PvD0lEiFwHCJEBaYtNg
tcul7DjR12IkIFzTHkfOdGUUvVIt5w8gq2VVvtKHA/uasNYlg3u+QMsBW8an
246KVq8XGnqRJSKwLJ0ugjoyRblHZj1Q5nIhT011BN8UCklWeiuMmDv732rF
A4mczJE/PXnDp6NiMCWsN0Oq+ozZZ8Ze66zlQMAkk/8cY4O4rVJNVSCPTRCW
tDdkiXK1ouZheDuBGkQwx9ZXxGgOx8YQatt38O+2vLSrN+JQSgIcjO2w6L7v
ParbJaErCH2C8Jq1Y63QfBsT/Bq7Vo/gnc5yr604iuZ4YpkbC1Kg8EakInbM
6B4xq7A5pvODXBokOc3HYjAVs6j8Iln82T/7PWHitBQMXKJdq0AUxCTic8uX
bkplj3+xI84vcnuT8t0VJ0eutXaEWnNcTe6ZTENA/HZXANLH3B43mJdEMxNo
xvb8p2x7ch+x4bbqzfyrJTP9+DtpabZDuE83w0PDVcVxa2moI3sMxdXrWcUz
hEx0maKhnSU9FrKGdKLtaxseeWSNLHjfg7QzdgFsfTPE2+lTeS8/E3CBJsk4
sY52MH5SDIRvzIuMA5cxN4TbqjG5nS74JjzHflCekTKfVngkycwEMBoyPif8
fmZpz6agchYwmA6hOGGSg2jCALpNQOMCYdJu+HtRpVRu/RYNE675ojViFJZ9
OA5CmQMEpnGahBxsDWpCsEsCffFQbwITK2J7nhgoriSnS+iTaypa95YhMafq
aszgLYNWPMpOLFRkqhZRT6QPC4xqTX5mthFbwgQ2MX5fZ9+k0za/8ZcgTafC
i7CfhqIKBqKWwjh0Me8W8BXjF6rZra/jeU1ngwYIUgWGAyfdC8rraNP+38yq
55lzibmfplHJoG9IIH7Exazvp6uSfh0V4twhwp0M75hsAPV1/kO780g9ySUP
+urVSdY34ccUjTrQRPl7ViKWi3kQm7UeX+HRWElaF892aM+wspgzaDW2VPWY
EBuz1oNdr35mKGTuIIBMSTBV4MNl8ww2vgsnq+zDeM38aHAUkkJ5xPvf0hqq
VcnMaM5vkB67OaKv5PFke6J2uVkTIYVB20xjcH5L0E76UCXam5aYhzPK4zK7
dESfXNiBUmlePHbcJqLlLlst5dxYZGQSe72pRjDfUsBPSzK7pkesafi5mfub
jGyUeExFwSZ58sqY6058OQEj/B5tumlBS2C20wBb78YVBiUL99cLXaTAX5Tx
YKX8/8tzGB36+mlWkERcDjY164hcV3dsd16TtVwVldBb3vAsYDbsJ+gqbH6u
XRHnT1JK9IlS3d66PwhqEdFAUvSnnD1AVCRwawh2wLCebOkZ2qf+P9S0NLUK
f0kuuBO0ILHwtbdKjqoi0jEgegWBRT7eYLGXb60okSz5SCn2P7wgzoCJ1pFO
8IS4BHhOCW/5EWetp+O1duocUAxPNwd//O3bLZrqc9xMXXdaYNjikxl3oNxv
umfFFNaAXqLaH8HdBOgyv94n2EpTdP1KpwY+AQ8etI55589jTMwjsIJL+7OL
l93gSijlMrNfUkOg8cTaDEOsVdNa46VhVTQ7NKeIULCOYUEehjrcgGEdrHzE
zwxlUNVhV2Gv5Nz7NzUB+1tOJG78jzKvwDwztnx3T0wBf+bQn0Hwzqc91I4V
TaHi404vOsdzfyPJh3YyZJ1EDpigQE7NbqZ+DbV8AVtzsQV6cPjzFqK/PpPu
03vwiOr/+NjRM5yZF+kCTRWSD3v3TxL8uyb6tGksciK3n8NbmkPz9bHJTNWA
CnmaddBMYUXL1HaSag3o0Hq1dwl0hxQCoAmuZNWIzByqQnINMgx8kYY0URoJ
g3XP3T7zjypCnXlH+T1qa/6MgPDhD1iLpk26Q0+HNbpbQWkuPcHCYxakPgNZ
krnrzCePZqnw1q8nBQsII7flHkSJ4BMrm6saApU+t/FLEqeb6NnDHyoiJh51
ddhWr18IcEGhW0ZqLFfgZkEPbIstfdoZ6DCVlDAtx6I5XMnX23hRbDerTpLV
OkZqFwK4jx8UQVwRVEIKGR1IL5sgd19OB/la8gfL634ARUVjaUxgNQSctbWC
/BwD4J7qQHQY4BBGh7ojBwdwrvwkyJYgwCYXVuBgiLVHxfxjFouM7GABLYdG
rPYLudrLfoPMbeO/7IhpvGErvmCit0PTUEblDsy0jOfCVLleW6HXQ72idNMZ
2XbQf76cdWe9JEzzE7w3Ve0L/UwPz2TWNka01z2ZdUzMvxPcmTiu/+YT3NQK
LZ0k6SGp8VptKq5anGo1oe3DeohwZU/wIZRRXw/xHdF0lf8LIR+PpCehTrK4
l+pRRux1fz2agHWUAQuRdYP89nSo9wsKtyopCdnSVuHalibAIbJCdyu4QNfY
mAaCyoOQnT4PlP3HgEavZTrAV5Wek4pQW8uEg6c3fp9ABXgXj5BPJEPAudtG
H51Xd15yGphwCPnZNd7Yqghp9FuF+ADgX+qWECSMTskazHqymGkmoLW5w23g
qQ/AL9VKBgIzeyPmW5qQy1fTHNn6jLux+BKkt9dHr+pcSgQL940manVd+gS9
ncYWFjl1Fq0e7u68zyHnU38l5pFeNhyhYU0u1cYX0/U2La8VKH1g3Frdvs5z
dtHnQS2UDlVRCF3n474ZPZEDtyxl0KOa9Q16E/6oE8/7e9/msOgsopykZyBf
c51PXEYorYpbXJjYzW6kwE96VH9dktSZPx+9IoDvBPRfGry3UsQ/hcm9Ss2f
5Z9w3GurRcTUtkuaLQJaDghNQDerX87te/lERN4ysYxs6ZhPJB0mRW99PJfE
zlrYwbjmiySgonQIiz8vamM+Nnrm6BbPvlRdiyu43Pk1jNsqe2DzTZ+2jJCC
yy+T/E4cBDUINjnB/NUEcOcA99QPKEosKiqQtBhj4epFcBDMGKY6gWSfHhaW
GsCiqVVVKl/B2ZqWaKK9iZCSCOaGtegASjmRK7bNhfPm/OjuvwC7XmDEi1W0
Hxa+dnLB7hRXDFm96+e8Kf+KgVqMvhusjawn54g+mG6aL/dpa6yo72DNRVMD
BdVNMVaaWCnOMXTH3v1J8wOGX6LWlsSvpSxXr4lysnBWwsjhVSpQXpBpyPta
l+sQiIlOLBGqbKxrK72bMWD2PWTl2n4xWT5m8vdFBpnyhEZwB3jVBzwJY05I
TTjkuraS0jHj2Bi0AMDWiCskj/wvj9CEQ4dxlQr4SJ3fX+QjJZsHgMAGOdxt
OxauIamK8x+ZO9W/dGArObq+FB8KQGNvEXORvCgQ4Aq7/dVdfxoX8Nln2v0s
kNT6BoEUKqHL5U9SGK2DC4vvXleqj0e/qsX2boDKqzxaJvzYQxmaOe/fDSLf
H5rGeNMlsdK0c3BYxcvkGpB5Vm7xa2eSHxpLqTFoLShgyPv6F0gCGMb51eSo
Oe2AIsB7T1QmgKOQaMYr5muiodn2v2oD9JjRRBkfjk1ogWM1xNRjBWWexw3k
ylgAFxiHEu1DCVPPJuTE4dHnlmpAFKyQZ1vLnujsZjQDUgWaR42nTd5nmWzg
wPdP9FeosaW1H0n+983DW9h1Nrx45b0wiK5JaD+HcIlu6IUHLnETvUi4caJW
ycf0XeeQMesjeb7qTTTPhiTZDDh/n/DMxGnYl7mqh8StKJabLjT+POvgXrg8
q3oyH+mKgpsH0BcK7nDEdbuOYYhZgcSPW6pkR6pZrbEX0Lm/31XrymRT5fOc
Jpf7Jy5R2b0N0jHWJYSD8n0FriMc1Ncg8x0eJV8QTd7T3sXrDzHEAVdOfke9
aJ6SE0GXQGW9wdty13Vd/oyY0JLK0DAPFgeos1LtG2m1UBhfSxVScxSnrVj8
LLNK8zhGBYDATn2M3DSpR3rDqQb0YCpvDSxTfsOIK4VbFOWaLIXcvuaS2c2S
LDpbXJyBj1ZEu71dY0O3HqBRHuyfUUSn51yvw8mtM6JCuzHvwLf/7p3u8i4H
VNLMI8bXyfIvFUIftH6CLWd+G7w3v1ugNp+jx0cVWrNyobomuFBPBomtGMvA
qg5x2WBNmks6BeJVqwRA/wEPI8iUHJHXrT+rI5UWXCniRi7nnU32L8F72w0g
8fyUGozkUTjd6ihwNWYNl2HIAxvvSio54fYb6jcs7aHX/iQQCBlfz88mxrHd
dlglNlyhnbCq5NFlUSFr9PCKTA+TJFVBgVTFEY82xUqhXfbReNT3j+oOHjC0
ScOYvxJuvIDBbiJbFIn7mZE9Di76ncQ6INL/cK/r4nt5CzPwQ4JLapCIj513
OVRqoIJmdqcgEJ5uKPQxtkpE0zieh5/iMzZsV7INWNQhyqqbICLgt4ygdshE
3OfRXusUTKbRfIpfr+hknX1MxtE9LvxRndLBsdZubE6pjYu7NGuVEH171LRu
xYw0UG6MsLtWdRMq+P3AYOjatVadcVStgwGfXaf+h/HZLF1WFUGydDcrIJ+9
9bFHr+777oP8pas3RKBWQ55AxeyTmNAaMLEf2fXT/qLuv41LEZ/BG3IYfacN
oTepxAgbtdiYd3Oqn2OsLehtciR9HXj561hciW6Ktk13LXSfveIuwk/b9iMC
uAUCqkiNytR+YOnCq1dPCspO3v6jV/8Uso8lZA80xeUlJGW3RAeal4is9YNh
BGL7uW+ZGJg/JMqqaS/Hy3HtQa5R2BC4rDVL0xRoiICVYmo8vNrAmU0VvMwn
+dxOMWiMOPw9SCjyM2ZOObXsPR6Nk7JVc5qgpnT8UHq8p6WwU7kl5Q4MYskm
zFva0OYnsWVHdi8wLrYojNqf5hyP+O+40gbhX+Emz6EYyB3FkTiT57n0xdXt
Dx7pBTlNN4ZD2BVHBf9FEv1TinvstH7FmwkBdPpuWp6gBt/RrLyTN8zCO0S+
A3mVAXlDzai55rrx6ueOeuxhYasRP/TZSFzoh0fiCIQ6nfD287bIXp51Jrxc
kKuPNii8ozew16E1jU+tNqF8vmlOh/w4X+NPbet0+cbLMu6rlZZyc3n5dJ9Z
1IquW7W4rOLAqxdMI5Qw5fOKnd65xNe7dSl/ppo8XCMb5LM71cYY39TAozYy
Qo6ngWnD/ZUyszCJszoGAWFcz4q6y+Bvj4278CEq9l9QaikLorVl8EnaVBjS
52k506QYV/eXppwIllcXcU2pQ35Z5z9vgHHeT+aEztQNwP0GzsQrk7RvJqFa
NKo31cVrJtukqHd8XQ0oD3l2+64TDqw7rjoVKebY4/MSDO/xUpWzTAF8A5LU
d4E52FgIQI0Qb+dixO/Qgn5dTxwlUGZIFDDCKXi7nncg4PV4sMsUGJRcLDiX
gtNLLOPHLGOVB0KSJKOanWnivg2jEZajni5+zy04KCY+BjZYFWP9xpeHyc9a
0yY+6p2UgoOxSopMHgoo5anXsxr3O5F/aZwG4V3oqFfBT0mhvnKXsTL7MCSR
LvOPr5Mq0NbzsykdJqgfczVlEci4VjI3svJg7F3ZfWK1L1wVxQe+yOsD21D6
msxOS57NupQU+L3lhRT4SkQrH2L9alsh7QsNdu/3sdHyg0M0/6WOtj7XpzRR
ye8djF9EK7p8V4DwmpuS9oWgM/216n5+OTYeA0w751VfKDc+aLe60rIjZz9X
tUxGxzdCppw10wNqZoThsATn2pNdhso4qvp+Miu+sVnezno2McLA038V8f4R
8CUz1Ew/8ah7wSDaNSrvFxaT/lOTsQXeP4ai4pp0boSYDEu1tmjA8VJOyRj3
mIKMN1BLK6pAi8YK9HMmxEW7RHWqV63ppu2WdBn/OuQ+OGqtqacxb+3VceMc
u+hAWM//vOnZU1yvIXYnMnUi4CJ9ztrZyCWpe5mXuZwZ7723cJIYGe804yOz
VgrbdXMmdzFZcvj3RtuOu4dqvYtX4Wls5BqrgJGzhyFfzqC4tMOhhqh0lfVW
tTjtJLMxhjBh9RkGjlxM58KC8x/W9neQZBXN/vQ9i2+zUs91iXfKM65UbPAj
rLMIgdHEbyCEi15qLeTgMcFI66EMcekaBWImHvkI53U2eTxzYyiuY/Us8VqR
QCNRqTNCK6C0hcsULeEdTHUDpfpq2twm1KY3B5sJCDACHEPbLW+J6C2ITE0R
rkAMInS00lURT50iXd3bElybQ9JP4Yqxms1Gym3bYUWz6Dz+8+z8tbM89g2k
VjR73hTy2ukCesqQ9HqC/WUtZ/K+7L147zhRrxS1s/wEvcGxvnC3SM1KyMIE
IPuUyOwckst0YFyZlrYxAYuGNg1P8CgDfVCmvBIG8e8CGRUqZettFpcCRN/V
CHzk349TfT31kIbT/qBVOt6IAnBnl+l6I2G0K9EnH6kOfZiS12X5EEwqiitN
2lXYNPLSqeOOJlDHaLQhHAnEszuXqAW2I66NNT0nxn+e43X1B3Hd+a9CQrTN
4/3PnCBjc2DnWuRUhFzpL2kVErAU1JcJDma5lZIRZ14GswmPDj+DOCThMnC2
sgyV2e+djBapdXrz0Nq6QY3hFBK1wA9MpbVkKEpIL1Bv915WalqDcx6UCe4u
GSkBpaBFhMePS3t9S5rKXhp03+5N+lxhJsQtSwE/lrDM3ozbWLpZT0bnfbQd
RJJUPd2vr+kkDHSWma7y9Nw5Jy0LsY2ui5H5So/J8Wv3eYzqI1Tzzwkh/gP2
NUAFdP1RxYilWxTSCyejuPxiRBgwzuqVvb67hYbky8p1q5yTWUlOO+zMmJla
GVAhw7ZIRbHiXFuNTKdeP+oGnRmbdtzkU91n7+rpPhwANu1aaSnZYWvMWOPD
7bzwZmt7UljS1523KYW+4KjhmND6S23oYaybc7gpgg33sHtsWLLk+jh25GOZ
qGrK+CWJ2Wmc2Lm0GtXA+aakxbwx+B/OIJb9osedUiTQRV2g+zeGWcUnDjo8
wWsWBfbm6p3d70fVytPQzapP5DxMzV9bJBQRwhhJ0E9qh6XTHMEkEF/mlGLI
9RDzIfW32Z5SP1Y7Jg3CHqEteRhkfc7ZwnBSJuRQayF6lMLHPDjVN8DjIyep
hq6kmXa+jXe6SeWmr8BAWM9LluXSnKh3EB6mS9vdFZQVsZJABYSv266geHwg
QSUYIeSlyo9tOVmyuUJwOst52nBbzXNjulagqJfTELvs9hlVLN0zXGMSxLs3
7X5joMAo4mH5w3ULuF6MDV02hd6nZ37nUDJRr/QzhZy3tC6NXE3nfdjCad41
dtI1AKFeIu5qzKkPPuojHOyS5kRujnh6QNvOAlFm/a7bjibeinJ0ruxzYbpr
A5xtmWC0yxvWyl4jbB5+M0qzbp2w5oH6Ub/vp/IVLQnEczsAt2DpmaoOYHSo
EQ3QcAJuk73jNfU4X9nD9K3LwVih90x1l9PDTKvVbhWBLv4D5TNxJmYYPEUo
EthLPrZ5QzAzmyj9W2h3ey+QkbQXB68rdReC28b3z/hBVdvpA4hHs1e1FBvl
WR/HacqWgB9pG2WnBq7k06utudgXvJ3UzsLVegmM53MRDoSssDquo7zESefM
3+feCA81pHq/NDuMwAQVN9ppVRgMAWbtcFPlXViMX1G8Ve3zIAKnaUROsmZm
homS4vGEsV+ZAU3+7BhZrT24e+GNfKk9176+scGg9dORme+YGHibk4Fcj+MQ
V7JFN1wq6Z44Jdm582D811gbz0LDZF3U/15A2J9+u3EfWG4XOPxwNMQ39Zbg
W/f2BklptUpKH1lSoqfsYNw9oC1RSnYnh8IK1nWpvG8Bw9zW9eLrWyRRRzlX
Uj4orV8GMBtRNVjLqFgA2g2O872fyBYjgr8/R171s6DG4uzFQ2yOxFo9N+qL
a4w7DZEqSVNcaNec/YKp7lP8fyzDH84Jnv3K+KCBI5EyvVkBbihPjhcCX7hL
MRasCq1FXPqirAYs0I9u8Q60PJuedFt7avskmLBnlgE53o8CGhCOt4WMzyPJ
RJfoeDg7li+tXNB1xvNbkVj45qHMVIst5YhHok8HJPL6JlVPWV/6uNXs/csf
zAuvz56xu1zD59lxH+y06S1hApcl2Go1/IMf8emDZ+W3WrbWWdWkgVPMt9C9
vsMeztarM8bVbryZzWvqXQX0i3Wps+sX6uwtIQJDunJZBRbJ0JafvoLGElFj
b+8ZCHHzm4Fg/1r+asufeMUI+zXA4rnDrjLutjA9LaAsGVsO/dmCRvqMhyOW
2PFim7hPKxXzf6LeuQw6IcBppPIlnShTJ3XifApfs6LIl3QGj+mRtUYrxQuZ
NO5N+rW7WRLk0OlfCX0/WnvsBPN+IAU8ZBb31k4vxQnIV6DqdtgR49stZDMq
6SCtaS2WVy3ZqvmG/N5EhnuN+EVpQIF7mEKhYgv5wtj5SkOJZFxhTCGItgIx
ENqGrrHKsMNhxWdOGygKJsWCZzgMA1h1mbBFVD7wweQAxDRxUSBZsF4rJlu8
ohHZ2hWSZwLrQOULx+cXL0XW0agiYfkCcA8Vff7eAJ7uBT8nq5S2WQi6xnV+
fb0bcZ3uWD4WwdkIesgFwdlfACc/smGa88M5YSZqR/iDzKS34pGT1IvtkktK
gV0yVt7WQDuitTsa5EWqtoMLYf3+gLexeT78e6rehkoxLa7hWNe+5x6gSUq+
kZ6TtlSfy/RFQ6yaCpYXwPImI41bHwV4tLGnGuGwjfX38IJN10fAm0bPEisy
CIhX37jHj9VHT8LgD6cDlzX+17/uEA2knm1n32JAwu8Z58Nka76WhXs3Xw1Q
P4RvUuENNaXMeFX6qJk6jvMeKO+c3HTSS2HgSmn89nzZQaFN5tMnCo2yynVq
V6DcMKBnn8v/1Wf7SKrJdStxxFNedkokxjq2/89uhfKbLOcvBzu7CtXW0G4f
uk5qL/qNtBVLaWK7g+x9mQxaBFvEGhe16WGsmljFuYx0sFcU0EzA7t5idjbJ
7FJOE+tmheVsLxct3XV5u57s1JZuE9e2ZMACILagT4CJxELD05ky9H6BM/lV
TSdO21bBoOzuPIIra7A8o+i+49bnfbyLerjNpUPJI+qP3hWblxwwAm1fvJUA
gI9PAMCMw17RUxHrFQiRjGArLNJm97TJ42RlhNkZKWPIpdiHiI+qTyoa+AHk
K9OYS7nCjqf+QLX6tWTgIP+Hzi+nZxPSZ7txIFSI2Ov40h+YVmWpNwtr4lCA
+sQHcnNLv2+GvbfEsdsYQBVYP8bkf8hxV2rFhQwpIf0UVCdDT9JxX10mGIfq
dMTXHfnjDi/aaLhN7a6ojslZt0y8+g4EgtcuzzB5kgKwtJUBphVxxj1xFGVd
U/bGeZF9vRgUl8fL4d1op6S7hmTI2S5mwQz/kOIPQzO7tU8iw40IcjiYRAMo
FpuusXBWFy9/Ty2heXe2clIqgsZ3QUbC9qu0bP3cwvYsEfcgowRUFj5E40cN
hbTKVNV7jF8jB520X7gGJVIz0BYOLt+kthII0xlrESG+SnFfcAcrEg1diBGW
F6YAnh5D1GQRdlWHYzMYZuSttUHbv/oymvITaXiEtatDuBAml5zU4MwAGKea
CxnA3RLhcG0K/BIgIMU7KWEoxghxaBGEsCeVoXBi8jBzbucCMkxro+f/ddYk
7ozLZ/BLdpusI7IL2vNB10yrL5QkMvEaTrUCQP0+KNa1knqIXDnRlFgvuhOU
9Y1PpOIIsRRQ/35gBkm4H0RJOwOA1rQU0b7lMFNYU4f27QTWy62gMwNbfmS9
74dP6R6bdMNHKyS+/lrvsz2M4bM74FkVsGe5GqZBonxMDzSkpP6Xc0jwamhj
BlQZ5DYhUKio1XYGjnRP82DzsZf605+GEizRUmry1Vac7Sik+lq1IiUwUmNr
4lS/nTXF/m+acPP+GmDB86war4Wuie5EdgpqJshOyKOQM25OJvw1k2boGvs/
ePmZrUE7kPaLrybI5PHSZUN54PTQz6e4O9+ZjyAojc82NRGF2JyOot11Dt1c
klUZMFw5wQ/Vvv2rHPPSl/aDAE232bUb5LeJFcqyRc4P1thqwN41C5tHHWbj
LbyxHpej39bfiiYsDN6d7Cz28j//dWrvO0w/I+y1wiidmfcp5x1lmnw6h3cR
FmkTD7wDI2VAvvknPV8cwZZrGDI9OpH5zUyuEBWPMZ4F4UCS0IKVHBNWD7B7
ufO/v84trjTibR1jQRT3e/q9Am5FCHeBhN+ZqmJShUw0si1lCnyd/llHJR1f
VZpWFkwC5/OVXHdZrILrUBBIn84Q1nPdayAJ8X/ZvhYauhH5+107+/xDHrPK
rfVz2VojvUIRCTpHoEnWaHaU5ZKX+e7YA6+gtsglOfOE+xb09QXj2GExHiYa
Xl44pI6yuTd2Y+Y2whOCDcSNjqgaQ+7Ep6CUHRJDPVHnf5GxP5QeZvVGgHQO
A9zZ4qLJjaSGd3SiDQXIQCR1ja791/DGke5+1PyD4enQSjPya7uxH1YD0ELH
VLWZnN51gOpxDy/vUYWOlvrNuorhy7pb+IqEP3OtPejjL5riNYfmMeZgn4Lq
ALJ+dugIQ/xa5EMEtJwrBW/Wrf5Wz2X1ZWU7vmO96PUvZJxNlne/9YInMRSt
wI7YDHeMb6YlgRonxQM4lavdBe+ryF04K/HkldD3rmgsgCggziy6nfOfMyNV
La2s/HdBDIRIJMXbefYbX8ISPbGRnRjnqKd/XPYBwn2DSFqhq24KoFqzaFlD
3FCh6vOVCHeU43DLbwBocAAAvE88v/iTEFyC1hSpDOzMGQ9Q7VV2A8P5Kdya
MUVyYiOE2wPIU37K/65I7xCtyQs1wUvnqvRv0T03l+U0+5fPtKfHnboC5oqc
fven7V2r8s8Sqk0aNo0tdKtvZJysuGvBYibiK05RpxVCASxIslbrXLrO0xAT
aEcwL0Ztb6GNI7RvZQNNvd145gWIyu/VYzROlyywp1+rOK2f5hXepanuroBr
Mffq5EENrPurt8r3U2agD/PyH3Lm1+8TkevhgIwvOk5QlSY8xALeaVMNdCEr
O6p4abJgRTFhD9LQtzHByck5d14Y/B5hcU00BuX3sf4SQonHhpbTMJqQAuMa
dfzS7/k4RenKRuVgSQgCqCC/yykyx/0o5ZK871kvQYmA5lrX+H967JlRKc2D
YYlqP7scH313qR8KnT2OAHxl99uqqGlIscFDLtkuloucxIC5cbhY3BvebErh
uzIKmWvYKASTO1BDOZsV3jjTRtaPkwztEyYb3OSV3H7mWjYaeeP1NmNdSRug
ipWOL7N9vCkr/bnxFLsb8AJwo+TYpoQU6aYndciQPJTJHTJLLaTIYTVQqVfs
utfYHUGCKPBOpf5SPYqpbXHljt+FFyUGk4pInas790tIx7nG17AWbxDU+HWo
2cpq9GTrAJ679uvJQa8YAE8yG4ejUAV+TWi1bq3mLNXceqvfMEgipHI1d5Lr
QdvEZvaa1JMWsMRhEusXSrtzFpfivX3bqO8Z+m1x2+d0kX9j59WYxsFnhspg
bRq8RfCX/DgP5goirDAnOF4zU1AUikDuYRGEx7AtQ3kLD3RsG93L73Uv4MEk
JuAaUJBPwJKRwZX1SifbM+JvOCO47d/xDYZnA8J/2qKTOTTIsBbJOhSv1O3q
Jfo3zN57Z+5DYVe46tFo6UeaDGKtTOPfu2SbcrhiDe/AYsXhW4nWvFQENYlL
0i5lcME4lx2X9dTl/ZGuHUAWVlIrYXZD3iZ6g9vBLzPlbbAryr9DmmTUqVSb
JSSYe+X9sZeET9TVdRaDkBX2Dvzsvp85oGRllMizBXI8OWQ4ydZZyaLwpsCj
zaY3b8b4SkCrk8I/+vAlMtS5ZEbGSm7u80UqVHUQvHK48+VD48gdH7F+2oSl
A/FC4VSY/g5qtuV9S3m63k9pLTMfK/Bx1IXfJ3hLUjXqH5gzckEyfiHl9Qji
YxEJ6Gf1dRfJzVTdinSnASRskkZGTY0NT29xOOcxlf1sqhJwGyA2IHYLUSCD
+q2Z3yV50cDxqr/8UvW7ULOgU+zGlts+WRQAXBZ7OWg1BuqvkzhT4m45fNPp
+fnpA/YUoneClvqb8Iz4atQIbo93Y2faE1Ai030yjQkr1ahHKM35yrUGjNcB
no+PgGw37j5NxmN2SSxQHLl+bJduOFkWM/sMVGBI53O6a5oNCkUvYAJGzHpJ
WyYSHYLlzuASJB0JvygJyA2vk23sTNQ7GLUMl9dNOkLh32R2IkdHCRFvY7S0
Wl8b+vuypdlZnIovbJrq1es1IUacbLDhSFS/eo5/q0bi22YnFcqBJ8fr8jhz
8a4ax9joQlf4bfP25D2/wcVt0bW5yB8YcrWS+Jr4ftV3nrYSncNMaFExnBD/
oK/3+PLdi9JyidtHh9d7vhrQtbetKXVBnI0xQjedDtN5irl+XRo05nkpJljr
yuUldonu4671fcIwYX2RvL7X60uOOQ9BIHuqUc1/OkjjbYNXKojgd9dDEFTa
mC2SxRCc95mi2oKJSH5p42rZ+gSghjUDBGjOogjS/zF6jW6lIuMR8EkZq3eN
kRZbsl3dER8Tp8o7p6p7WLsceiUYFvwu2pEYvS2qV8IYi35mbHELoZvGHFMZ
D5ytLkK6h0HWDsHT6wSOxKBrnzk6OBoVVfP97IasnJr2gbHpukrtPdQbqRj+
arVEJBP9poykkwrEHiBOt+YrZalvkOBB7cWR1GZuWT0VoZd/4cVnLdnH63IS
875ESEQjS2K+zXiBUIjeDCNqbHeJw/ytJIwJATzZHetOzJSjL/2K1+afLOjW
vJc/jdRCxv4GYjAgyAJ6vkK/dQI0YLXxUPXeUQvoQ5i79b7exmmlxs4+SnWp
eiwnFwoRYeVwbBBjR3HfQtqJH+2yfhk2GQHrTuMMmgh/xYcSFtL3cLg4ueQ+
tWxSIu4z5lzCChY0kiTYd/eFurvaTv/+73s55/PxD7jc8H4zbZzj4Ov47dm2
PgrqgC0MzfYSQrM3SfkOrrm+3QNb9DkFT79DJB7pTL9nHoALsOKvWcUF5jMI
/3Pinbsdqf64AbRKYDreIun6oSEsjJWwyY/ySxWcRVey0McqUNX6C6t/12pE
1Ld1F3S9Jpisd9llWQxO4XTeSw+sllDj9/dnhuCzgLfzJ9Vv5A/bsLcFrTDf
nxnr8gQsS/UaHCj71T5o+LXda4ezLwiQGdChtg7NuQ/atNK7SLDps3Ebzr1u
ONSPCtwEW9i+6tHvaaWT4hkr3k9fEM/SAtkmRdolCUmi6ufTrKi5ebkgT+d4
MYehKcGD6PNmeCJcXv3qToUQWFQJRlsnP4zNJHpggNZ38M2ugZ9PAXSg8D/6
Qg/o/8BpcaROf5HUKY6gmg2ARgZI09XBh44JFVNDnx8luJv1N/519pdaJPk9
7WSjClaclw0eGsYwFoPJA0NHv5J2+eqTp9zMTlAGICJXHruFkUF4eS7g7mO4
yusl/cXFp/zfZ8XPpVARhuInXrRqGQH5/TqlsdH+QzfRK1eI9NmBn73z5Pit
x3ZFdof5/CtDCtFK7PBTNS13bU3QJbIFLZvqcWB2drKRpFoAopAWx/0yLESW
WnHSx8M/3pgKdCMTvrQaGcPmQ5DzaynSSFuobHX4ZJJv1Gv+PTl4wggBL5Bp
/lNvnbAzUwFRhWhOi/pvj8ALd9QSYQuLUgTmtZWOztqkC97UQe411j7kyGbD
YlvRG53UwqQvIP9fRLVqwUw2nutT+Pbgl8Ax7dMApH+fr72/+4oN+WlWfT7+
faZEX+T4CN+gjJhDHvhOhBWPudUx3m80HvoLXhDXKoxXdEAiodYXT8ENDcpW
+k/A2WzoDozHCiK7gOkzDJ5rYcCMiV9hpyXO+HkIOk2+S+ZuxnTG7nOhPiSN
guyjMaFOUG42dgCNr7sHLg8EM9EffzunmIa4bnGWzHBKWIZdSFMbEj0in82t
byPXr/fB7STF2QmKP0d5VF95Uu8XZLGwD05QuPHf5Z4srhdtxTQad/MZ+yRP
fl7bqVxCbwN1ucC8KPjPNjDfk27l4ITqfbfuUHSD9SOHMEUlxVa/0XKdRg0c
q+HQL2ZqTcDptmM1ZFahqYqCvfngC4mJwfQCmF49dndtborvWdGjz2aeKBh7
LlEXOAonvXd6dg7SUewHLDk8q/2BVL9SMTYq0+jwV0Xoor5ltli7d26TjvBM
kfep6D0yQbER1MvgXXrCL3E6rqLsoCZWeMC70qR410iK0ojpJiDUi7F03F+5
0lUbgpvUi8GGCGoTaMXgPb4Qa2U9CmIJw12g38LphTfTr06z5B+N/pL/eMu9
cwQ4hfUujKT11dkwseuy+DVX4iPPB2+KwFgRqlmDPXbjpSmOkyX0x+gtJohr
8wVOCu6TqI35lKbx6lEKV/CgHipW2ejBDXSDY+oywBJ3aKE5Mc4OnXrdMgHB
ALHwsIIKZbvE8Xd1pnKsjFwCjcpSiDYhincx94yRzTHfBfk8H9rZ88IO2IeM
VSqc0WulkZCNqVqarJrtnI4awLcXFoLyyEPJ6qj/sRLt/da5tW5D2j9bsPdE
xZj1kH9S//lDdpggA2PnGt+IYHzX4ED4fdm/x597ziU9y1FCZIRLhyDu+62h
3ulo5RnsdPtbA1KVSh7oWJ3veoMpkVBkM4PPV4nuojxqrvHtUllFTfH1gByk
kMt4uH8LsAEx4K7hP/OPMa0Ifu6IrsnSkMcHLWpaeMgem2CMzJ3M03jEOtpZ
2XavflwY1Qo4TQEKbqCjJbFxFgK7tEGwou89phu2E2gZM/VP3NMnHeeR8O0Y
EJNfy1D0epf5VrRHKtWFqZQ87Uc1UJUahb7UTd+z4oF9dyoKhKKxdz5vlgH6
RkFVplywaLISx6VKXgAyb62Fc5ZfNVA3MGeAXHnTQz7eMOdS2TmZTIHXdNcO
M1kkRUHl1jiF2SB9WdpBQx/MTedwi4kmc2fZ5W/td1jL038NPu7XPjuwNu0o
hpvlnTkbO4/UWF33KbPBoVPqdjZHUG+s36asfzCgL8oZhJn9dVyjtQ4vdPNF
MLDIdkDvn1TxFFD1R/iV+R8T8Ay7gDDSYnu4AojMnu5XGIPPbpn13+QumI6W
l4rlC7fXcm0KhSzlOG007Wltp7oEGTXOR7eaF/5MfiaGAFHTGIrPipYvs8J3
qqQlDcue6HnM3wRYbtTs6pts9/V2vhZUeidncb6Okl6CrWNbdxKzXy/k6q9H
kroPTs6wbHJprnZ1S4IxQRx5j6NsODJzVSHU6bifqFBvhLk2OgxYTmx6Bz16
y1E6HmT2HAuGnix2ck5Q+ZHVw+8BRpc81nh/S7AGrt244JqjXt4JaHIYxOg9
0coUEbc9g7fEB/CqRA0A/diYxsv0+oTY73H+dJOxpwmv72oNMGTrL52GpR7T
EXkl3BNXyzbs1kPBsg2jRftmYbMGdH+u7lTE118oj1a6DiQmQqY60ETwzkGP
bbVRaPCejM3k166iSH3SZsBwPH25+QIUIx7Lq9FmoVpdf4JWPSNX0necwexN
GrRlRFNEV5V3bOitGEnmR4U6x+hTT6inKANsifyP7D1TR6P4V689hbL5WVg6
gQxC61I8v2H9gGqRjE92VOjRErIdALbtZ/4WqFnHjMtRtKRsO1z8ovWRHdD0
XS0e14XAhKyaTyjjHR3DK6DurehHoSzhATse4R+vX7ysjuqkYsPW1CPlE0zq
SidloQL4GRRWSaOzySGsel7nDw8smmcp68b/LN6UuTySCg0KV9M9rl62VCa2
7TOyUK79ho0YA6jztmUvboDwnc2hdFEeEfyBuU/CU2ZwlWYIpBZUC0Ys/HZo
+Zz3p4hJ0DZXzfKgb1y7Bjmb/IfzDHLNneEm5v3KsDv4eufJddLej8ALAzl5
ZYtvhtKoUFLwO06OF2rYghgd2HQ62cXLoT45MOyCop+pGfNc6+tfAKmViR3G
qLZIn90XwwfrUSMohv59LP+bIE6zI/rFXRg2b5/LEd3yfkKQMlE3clQrnMyn
JjQJ4p+RTO1snqu+AqLTpzLnMcSqeg/gsVWmMNgwN8XIfvEE7XU3DuJ4gHGb
sDg+H3BfYqvfnqK2X+3zO4KdcBikd9iV7IMs7XlCkvWrllQlCiFTcR6oIf0O
bVOObsV1f70x9SvwCegQoYsvNtoDyjfWFBKsYjl/8/Cnznnlt+bSvexA5HFG
la+lab2E/H8fkByDj5fLXiIjl206PS8nMHwxxTVtTe9ixGbAtvG0AUdcMUwh
1oT//ghqCHPcM4vWXDEDq/CfjKgap9BJVUUThWH91wkSLFrBBzTUxisoXUQb
YU92dQZWQkzrhO2csWc+SNe1lDPUmulVbRyzrzJwH7gb7uMfYM26eMOYnJAx
DQMKtGZEVcdgSljthsnoC5H9NCElZoMWOsIvUGHg1jK+DGOoJ43YpsHOXzJ+
8u1KKn7qoCeoxL/pRFMqyxmfOxf1p4bdBFQX+K19PoQKag5kWXYClTocpCiD
inJKXFxn65fRxmEudEqVhZkQ8lmADzrJY6VlJu1SydODOvms3IDVl12iSVq6
b+VXoES6m+knu+AtXysW5Mzht2QL2xAG/mFUwfq+RkPey+o8vuS8c4Xzqn4O
7+oo3t5Dsf3DDDvFufqBIlOeFoANqMv2bhsgVZOHnFMsqGNoGkcKrXPEQDFu
XKZBpU4ko9slm/c3NnSE2GDsAt4FvsOpqgAX2JKP13vdmUeh29ZwaS7iKUA5
MLYyK76H6xkcNFUAMeNYDFCB4aUIRpJPQiszzWp3nlknLZhYqjwzKnSf5m9K
IRAAIMRMwuLPgqpo2hWn3vET7eS+p4AImwzK5kkkkgDLeq+9zcfeyu/cGzCc
ITzoKC2CX0cDNbUUqG7kkIwzLyq2ahJ0JVIe9pSrYDSRv5pKDePFOQMz7lBG
4HUhbGE+2Wd921WNJWa4tmc3WMUsAIZGCqjWJLMThQ2roasqP47MYkGXrqI+
FUluistmHWm+3dAwXvUTAYF4jnoGGW8Yd1gjZ5Qev1pfjNlJXRj6irr9T5m2
28BkNT+9E5IV4jbOVKatNhOxbO5XZV0GWa4w6pdm0CUQGYobyhV3EJd1LmqZ
pqSBXWcGc+JqwU3hqcrG9alfgMU1+22bhZ/gDEc4Tsi26cNIIz87+0rsLiRv
9//8XR+1dSxKKVoyqBEDmHJT2vzP6d7yZEnyEWqpR6tz/ZlLZK/I3rXji0hw
sLQLeYAA9Zzxg6LaJgkBO2SA3Bc/8T6DBItc1zFgseXyd/CqEGzz8d7lxz7w
rW+dFQEcTJFtZLKsoSZgquW6i4/X9eTkno3IukPoHevsusNukVn2mAC/ovK9
WBbYt56ruy9wI0JmYqjm8toxCHiLibyaQSptXg8hlYuDqtmC7YPSIEhjEa5/
rmQ5EyZKGwX/sZ1XITjeIHpC2vQf160KgfDjdWs6fajGCzJc0ZiV3I2bWu6Y
hWCpT2Nx97BHytMDNDLU3E8Ddr5N/I79VhrdUGIOiUPbR9wut0eE3CyQYyB5
jtxDt42YiDfLoin0L5LbPz1x3NqXqJfb+w8K8Swd+CL5PV3KkqWlgx+ND4EB
z85ctPwzfjC/qokk5f08cRv8f3lFVc1vskgBq916fRfBbcajqXZ1Goiq0flO
AnfQlroE5qYdJfUrkVbF1cKLIWoZ9Mlw5ZR2nNU76h4Z1Fs9e17aIS1XuEWr
DX4Jo7xYYg0FJtyJp3nrrocAUy+226SG/7twWk7GfTIqIp6JEkNNBGj0Q6Xq
wHee4rvStOHG/kVB41twDS298HiwQPHulE1QktN9ckItftkpe/vA8pqkB2BJ
K1HiOQ2Py8y+RQdaB9DUAc6EujSz2paGENQuocjH77E+d8GhosmwfdI7e7FK
2o+KV5uaQdB4Fy7zTX/5JtA1WxoUqPzRucEi9FntO+MhFzga9p7KNfgR6x6z
tfPa/YUeOqp3OLvDEQUBCNSZN2Ybi9QQY4V3ihZk7D/FL3T8DELg1nnabSXO
k+0UVY1UJH4g/810aBS3VP3QkMFGFmVG5TaTUraPYSgrnc+16ivNz8ptCthG
4V1EHv7yVTVTxPJmioU4mmRnK4CHZZTDnS4TSsTXQWfEM/Q9s6XEulvIZ9mY
gfwYLteIvPiJyTRy3dTF8IkkcQBW58FHXOqG29lw1RLQTK/Zchm5Ec+WeszB
SQa3pu4kvh8f1Omc8wv0+DIYm0Wp663k8TpEjY/f1DeJUYzRL3pxTC/+kPCs
KZ+5cSi00EMjOC97tyHW+deL3GMmXrQ1Lm/cREDcbPuXFWagstChPT/BYKbw
ZQ4/tnSSSBiYk/I2sdT/yGvLGRFUfcxOL+yjQdTz6jLCTTQDGMo0cY40Pfc1
4iX/bwzccbTM7eWv5kh1uO2WNcOHLyCZ5pJxlTwVdsbtlML7wUuQQX+LT9bX
oVe6pgrNZwbMOfOtGfydZJ4lLJQ/jdfsCjzSBtbufjy0h+yY3lyawwJl8mKN
ptmOGpA0Wwp845Z74MCAK6HLJ5iEyAzuiDM0B1cIW76VhhtVE97UPv3jtu1j
x6NxVFKfp+mgL3U4fk2ZyBGn2F3cdtBmVEPvKut+8anjekYYe0t9RjL58qWu
w7ZPHXp4RY1MqmY8spSO0A8NjqFbCZlDerpiB6ORZKckqrWK2YEfB9ctZZJC
7+4yzSGzSgod3TSpz76NDatLZPwtkNxXKPKzp65xsLsqw1U4UsptJChtxiXy
qM2bckKXCIAXToW2WKTd1MERPwf0HiIm5k0vm6F7t/ZyPeH2uv8rYB/F+4Lp
CLFwFypD/522cnGRhVze9i+Gk3J//vN/dUFvGAWDUggVZuWH6Q6H2czcKG/b
2eOjnwl8oKJ0ywXQwZ4JMrS8ndVzPK6sBBQwbHY+n3bAtJv+z0o+j+F1uBHr
lYdBKw2VZ9Q0R1mC6Enf68v3f31axHcMumuqo2RwaWvXh07sSCkkQiOYMWt6
ljnlXEqpzBgXHLB0dwruwO9Snf6wRI4Yn2Z6cXDF6KDb/1cxRCKc8xxeJcae
T8Y2JjCj8d9ULTJBnrRf2lKm0TwUozgjKOc+NKp4R0+SgytCix/j0Uxu099U
ntoGJMqC0BId6bOSXV75icsgo1LTrrSLPn0MZTOoa/khb47TB9eCGKWn3dcc
acbDvrV/GUVVplhT79Xl4uCvvxh0sg7Y7KlT0s49zlyBBPHRYZwFds1zvm6l
VZnwcRzI7VRqgYxvN3QHVJIbN0hnWepE4sA3EzA4zrIfs1ChKpylfEq+2c0j
udARwUx+trud/pJdyhRjRTI0X9ZpZ7wzoWMml6GpgkpNZ/qIaUm+8hcUPbSp
G7FpWCj74NUcti/flsjsI8vdDxe1AT92rVf3Ed5U0/2Gti98tgVavi3UMtlK
Eb5OKBEmDDxvA55JOBv4csy+t9935RueEdSaDPFQD5RPvlB/WF0ED4w9AcS0
kGduEoaqHXzWVwIDgfb+3DzVa7mRjydQth705mC7vNtCYOrJu9xqb0RKQie4
0v6lEQ50YVJP6H/IfcF468epKR49+x3gc/LAAQVe7eB7z/JjrKIoloMArSgZ
3J3AunJc8nx/6ML91m+X1XDQLjz1irt6xs7Aqi5hLjrBdutMzbZ2dLkvGlsR
pG6batlJHkiS+kleB+tpQ3wQgCttAUj7TfxqFbLt9cKgtheHSWcOZ/ricHu5
9Fk9fmdUpjgwGjHb6CD3U1Pj5Iy67qCyGx8eK1PcusWMalp/kt/nwLlWeqwE
niXGXguQ25rfU5+uhhG/L3GXHofotTrWGGEqDWMlq+JERO1Nq7IZsdJXPooH
wFyaFfegF1ns0Ho2JFIfyMlgt5JQiO4BC4tSA+CBjR/1H8N8P4LR9K4TuafK
rBInSpzYAGwcXmdlgKr6JB1Ci71yoSruzp2KUgH0cOM5+yi3u5iKa+kX7Tgi
XGRxMywNZHYto3X54F48nQgMR5SUE7OGX369bhI3zCcDgfrnQ72vjHvoGbM9
/Onnj229FApuWXucQyf/WLPlYKQV20FCAvG/vhrFFUeRtNQAMKSpuTTK447u
8ClDFoMs1c2UTSRda1404WEUeK0ZVilDFnYssenwP/xoYr7SegkSzecaV83m
8KUc60h8+espivvlTsgUqNMY3ms+FytpwTRfuNYrylhm7w9GUTQLVluZHKV6
yM9m4j3rBtxZOuc3VgGq68e6l3/4f63Gf9riLBltayYY1QyPCoRpjTJRz2ww
BjbpzW2hOgIYyOutYvATOufDn/D/OZXbC+CSbNXhgAaitk/XquD+hK4T74Qf
aZ4JNk5/kiwYNG1xvwuBqXeA0bJzbZliLcnKMz3OFL0rgB+YsaSSpXB69kxB
HG7MF/BpvSSlAEiqVg1Iz65GBE5KeF8JJ6UnAz+RJ38+sO2Vq1dtDvKV+qA9
wK46N3cv54KV5weg2t66HNAVlg+xD8Xl9P9q4nFqehUHSUelXdlp/njFyJ60
VKJRskyVkHzH7as63RcHkUD3rlv7lTB9VOFLqFtsYLMqRcvoZNQ9Z52brWMI
mOLLXz8uTf5LyhQX8wxTQitJYSNr/JKZ1DvxACI+AjCGj/KdG2frtrA277C5
7n+Mvyyiz7WI9kNb5xE3hHqWhrm7TUnebmQqRCon+RvabSSbugWGywsYU1fr
JrQhHx7O3bezVZv5bMiLGRJRVY+uyC06SlSdma59y9g/JCQt+Y0ePsxzQftC
5bd6AC1ypk2X2DAWeSkE5vH/jcE/Zc7fa/K3Y08v77nqwGSF2UEklgKVSaMp
g0X/Qb8jeVWpsB+c0XS8dqV+4caWQ8JL7MIQB+cYC4C/uq61K8TlQ7dDazmc
mPKuSme+YlcaeNcmi6JJXcQC2vY8vyNH+OJ2xEZprVLvTBODVb2/dzl4jqp6
wZWVkViUduO8lq0YDrHUrGpYSc4Vjt+jhFRCKNTe/ufP7c6BEWpy8Arc+NMt
n5RAN2d3d9I6vSsYYlW5ZkQaRzsq2rrk382g66aZH1yCqQ2OXYApcltmzKAm
VL94DHfQdmx8RP5IxK3HIqP/HBlPlTrIunZZiU/ho0n5S8PTvuG/averlyT3
ig3483tUn9Gb7eJ1oBMvGrNz3uiyKXnsc+b2iuH+eUJeKdl2kDQwKDtIIT90
CbqghC3R/l5HylT8hUI1QA8AQtLh7VHs9BdE6HBbi+glqGoBhI6oIggJccPi
5arWWmux0WTX6XoXA+cywQ1cbJlv2ZfqVqubabW79ulsK5eK9cScUeFNcxEz
hlmDABT++JgNh64hamcJIWenpdfA7r+rowaeMHMqihOsXhMufynx7PqdNT05
JQiQ79t+BUlApWwkiLvIN4mp/CT2Bh6HhpQBPJ4hgE3Lcm0dyG/SAYfgHRAk
wDXRWJarMUMgTggiuBrgqTpAzaPmFjFg0u/tIv2qj/BIgWyyxZNe5faGZrKQ
SNU1MWP98E8POoljUoJ1NTe3IzS3sben4815AaiWuGLfWwCz5UeHWRsx4USA
ZDdDShqrpSpm+F8PhJh8LGvCcn+DmCnoYfl6BwQMRh89PYg3A+xof38UkURl
3BC4mXWWpgqJ3VMXC4SpK2MjMY/xhEfcPP9KUokQkD2NDEkkSSg8ke0Q0l06
5SWZzFMuu7z5B+7SJ2PsOyMlFOYQEkpYNYPLD9zMXieL0m5DcduVjcf4hCJp
2LOVL4xb77LXoFQnaJEKWsSpukUaMyMr7wUKo6Sxy1zDobuvP4VBMeVI1b2S
DnDJjGXcnJ4d7XuAdmaP6C2GjVqkQCFRmQg+cgienKThrVSJbw1h+t60cSil
0DxsSWsGSWQorZQnu3OPXuhlNvRYkqJNDk8H7hw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qQwqtD3sZGdDG98lzdvbuzeC/YWcfoTeJPoywuxopIvBCWW7FoZ43etQWYYES0StyMNjjmwis7kAyUqQRd4OnvLrMwhu3WPtHvUTHlNBriTXJhhjBd5XL6+JS3qKGRw9FFUWdVbvDzRCzGQQfYl6BtYkf8qeKzFP0KjTgUavmB2oVYJ4Pd96aof1P5ctV19LFZZhI04S0IU/q4LHya5+dPquzZRRLgZ3LmAgdG2a9wjaJUw4HZLhD2ZUMomAKSjO4/+tUkaYKmdiElgdHeATNGfc3ZPfrlrbJolmzqfxggDjhvhI4GTG4yk+kxGWJ+WmvN7YKNzNg2tijls6jCD2h8tfk5JjNhR9P6/iNA0M9SsU72vDulKjZ8bY4Iysc+K+9/swXQ9gQIV0JlaRGnDDKiNXg8ZD61fVo6Le9TBY6E5CINn26Y2atZ99xanLHOe2+eNyd1y0A73RE8wF/OZatL0qqegLuOoIqJ1746zgxXvtAUJ9bTiBNmRew2oCTcNBP6P95YY+cl0BMPTYmPR3DN/873BbrZshVB7AfKLxY5xvdQNf777OqDzrBunhs+WyXP2u27y2jMb9T8dqY80VYq6eMzqFGzJBrDz927rZYhzBwbtb0Jy0NZ18kp2fJHosx0PAngAN9CmxMUEkx0q9PlTd6FSfjq64TapKnnthSDQZ2YHmv6CudkxTa5+XBfC2Vpv3gqFpnkLkAZQ/tSS4rve+BKeiitojBD7rd57ez9ecMtKOKCyRDUd1DdwL61pEgnA2QMuG+LQeP44drwUAwrB"
`endif