// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J2kyG4H/mJ41Q8h3ZOA4UzXr/ZmDV66XzsdWqqU32empNVO2AtNWrJ6UBim7
fjYbrMWb9HYdwXg2xQYc3VhmcOHDwp7X1CN2Wt9Vb5O++7Rk9gG+6JSyw5zx
p6O/it+7lnNVFRkp/3bOvO/zB6ItuzaOMe5RmZDgSIccksDJSHqeuJJ+qVgq
/FZsNslQhQRjT5LFNkLCfFfUMFsAJl8uZEY2kaFX3TVI18Y5ZeqEtj7yKg+g
UcG4Kr7XGp7xvQPhqz8cWwU3wS7SHW0hyeJbS/i+tm8EON7wNNV3gCdv3m5p
g/0MbT8hnip4rnptkQmZl/8qn8ZDlHazda5NYR6Oew==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MXtw/rm5Fh5J0yye5SfQEqI/0rtaauYHecv8UGHcXIoP5zZH3TjKdqfTTuq0
jRnQm6RPjWPP8RE68Fw5EhSijZ3mvtt+hMdlj5TaI8OZw5eqfFDJCUS3/dJE
DuV4QWWZ7sNc07UCK1gpkxuvffYjiF4SGUK1lf8oFh+HnkwPjupc4mBADQRx
CjJn5FFuH3I8sVeLBDp2PisaD0wQUCJjqgDS6GFAziyOhp8YjAq2ixs2DLAv
oY0xGG7debioOB8umpLpzeFZGrMI2QuUbIFJ+iDnG8ggffULoBiStZ/GK2Va
ihJnkgZIW5lmhrFrXzn/lMMrCjI5jAOmBw4FKYFqbA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pRwLizpDAHNsYU3qkenLVEYNOyR8B2Ndtsvmqmm/HIPzFVZrVinR0g8FZsLH
q+qZYyc+mA2PcfYG2w4ij4AmBn81yzoPutnvXFzCFkHgbEdVX4HJp+Wdr2LI
2tEccSIXUNYcz1e7FOp3EdQaUZD3bsGSgkJMnZJDKd9SnfIXcErGe56V6Mg8
NMu2MX5wmWZVTmQGXH9jA9F8GWt7+P94HWtkHZrLMzPLcuGLZqFTAalA7aFU
VBPkwOWBcWwcXHHPEeTbazF4p8SyYeU+R57xKwdWNOGNR/1MRIkKkhvBp1CA
K6KSMR/4rQsQZOuDMLygHUpDffUCoFujMy9lXmMo7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZDFxMHNE86WpSAx2tM7rCQIZf3sd7fD5/UuVwW0uDHwVJzfFd9DHtcIFd+KY
s6iYjnZBmbbuBnlWhCkmPtjx24hYyyQsk7nORgp+6RqiKD6FmMEw+CqYc/rb
gFicZFjGIJJOHwOGfEJ1ekD1dMoBlspqU3JzdQ9sIOWePov29qaRGAsKPuFM
YgHluxSnvRKVYyShPs6C6ujzHeZz92SZ9OAdW0TK+RNDMeO0IYk8tft0RlkU
kMLL0rYsD3957Ob83J0so50upr+cb67qtoPkOuGORKt2ZBHNrItIHa3qFg6v
zu+05mxGNp2QRx0YwTJQ48qjSLV3wXHMKX/kz2+WXw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
diA17l7MXw2vxyzyioNA5EIpDv/NEzL4HJOsdOUUb3hggd3KVrzJ4ylWGAxD
eTEgQ40rJqWFeOHbtxCj5b3Fi9YkTqZYJPT8kZ5AUPjA0gGnEoR1lUzMHhkP
5ndyUObjfaPG7GM2VX46W2hGKq7FPWu4Lacf5IECh4/5w+c0rMk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
S1g0WHPtbGK1GIJTuZ5gzkWS65TpBQ67+q24dHt4pqbnEv92K+hzQA7Hs6jR
hRShSfxkf2JIojvCoDahuq6tQlcTiXdHSbjRqHZXAIxjJ2vHA25VxunbOScb
QVQnqFGCaLxAnMtfb+HQQ5yankUAn7QTqQyDGc6Bu8r4dHuRSRZ1b7OK1tdT
zl5hE5Pl9h5xsf8XX+BHhInU+FwF+rACCdaP+4yWlNIqH6gxrA0Slkkd1+x4
8T4SJ7ve38GrlA2X43go7Kvi9nBy4Yeqf14dju/+WWsEHAdjNis2mCk9ktaN
29kmkodeggdnEQFphaEOHAJEgpIjyDPhtLPh8RTNx9uN96tWUkPq0URW2uDC
odQjBwM9XHIDc/5Cg8vN9fNgEAqYhUfMAMUTt0h1jL/NidBGKDNEh5QA169H
pseqdXx6Fh2OCByqpVOx6jKC0JCUjhv8B0CA81VoBMFGf0eQfrxhHd8eqg8y
KWkilw3VMAGYwJ8QfbRHepHAMvQVbgVQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
at+XEWasi0Ht4WJrECUIVXWkzdH8DUa6W5pNjapq4UBYzu3G7XvBlchlho5i
dAWKwSh8Vqv0fRhPX+9C0AFvRlGXytN9e5C2+CI3XhOtp4NprsslXucpwZL2
62PNnulghBzsm704Z7lynpcI5bKEw2imAJAXA7X/+pknMDTOHaY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aXKUyU7D6AuZmazgIqpTw65l6xkxFQHGlnrpQ1oW4d//QhFRDFh6PhgUmb8Y
Q7EI7PMKpoatWQO1ZT24VnEITzoAJz5ti5xREsBxBGj/nJFK/PnUh1VYOB6+
CxBuOyteeEKcYMLmpcnm/sNsGBdkFW+EiobdSrI469BTyj0ve9o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4688)
`pragma protect data_block
6M1mEthtL6j0SAqWTeAZK5ZoCECdonbhJ6YczzNRxUia4VfgIKZAEnekipll
SE2RIgKIYUl4+i+6aU28op3m2lebIoaBzXanT2fZGATDx9LOBuyuQU6x3Ihl
zBtgQ9FqwcPsXaK90nkgAFfcg0XllZJWKjF+fGD+f0pvz+KMiPlXl2W0b/79
tX2V8da1/cT8u6m/K2UC5eyKH8sea70TjR2JmDRTWdrxtgrbBBgvyw4gdgAA
RWd7O71oCl534i2eLrOmuhs18+Myp3nv5misULvtoSzcT6MC+M43rq1H/KIh
PzOU9zRplvMcm1N5MiDKmOE45uB6kGjcg3WEAg14qBS0iW9zkaBD6/ZtpZRt
61jCQKjW7W6ak7WYukOn//IQGaaHTuIZO8DEju0SoKP2eSoWzGtW1Hno61K3
X+UOJTljzWsmFFvSDeoAi9kpYMH+khk0mcMZDpHolwKsGX+euS1bSBrw8CBL
HqbjaP7mzpA0im+Y6jTdgmC2aXvcQN4WGXJnh7ps/9ukogNHI/g+WFmkBhQd
JVbmac/5usYu2luraQE80BNkh+MHwu5VQl9/kIWEUu3W2xbWYfuYBZywANcG
IjfZ6vX4JkwhRSsp9IDGPMQbnkTXQZC+MEh3j626xGtoN6IA3EkR+YAC57Db
haqcsIC00nNQcyWCqpQIYbX75XsANPplsnTBq/H+ZwkEyjN9ioWCv2x3XoWL
HwYTab7AikSZzTwl+Y5sfJT438j2btS4cXa2OyTLz01vQe94mtTnJyjZkHnd
KaK1T14yA+tLbVGYxd4HT1XR1rminEF6oPzQFqY5xvWSuA8nfw228yLhXEMG
HqXFxQBQzET/yqQZ9dWt9wLdHblcQDZngRuR6E86e+ybuwUnNOvhIUWNljW/
YZigVk0Oh/gLqppLHzf6RiI2S2YJ/jq60/ZRTLV0UkHPAsKB3lMnC8mY14pn
X0angQeniOcpeNDANXwXP8iIwCUnEfGB76VXpqt2ZFRkht6VFH9CfuWXSBw3
1cVWrFBpY10AuJkxj1x22CYMe9GV/zrN7ue1WQiLe6yLdWKNNGU850Bd+lon
2MxiwA8paty28jPiFgeOb9xiCA1ttEbdhg3KEL361KTGfbUSlXxgPCjf25BP
ESo2oN9Z0s6lAuCIV3QMKdO1IwotvbDHyUho5AQqiFWrlb4qh8CsybCTBXsJ
afHHf6otHJj8w/b5GeuYEDDD1CtvQKbpnyDy9/ZArAhoz9TzSJDkYorh7Yql
ze862cTtgzbCCDpaNkncoONVSTdMmNN8/8kxe3iH56f6Go4FMRkwsdR7hBCw
tJbMqC0gGHjPWmTmeU7PyVbeq+t7Cnxz7sjOi087hzWjfZBBcp284pIpOaDM
BhIIfsy77kLJYA2xTgRHDUhYKUC6VwVTWbdqxo1O3iEAQVWJGrz391kzpBJA
n8yB7BR4GHLm8EJK9sJMT7VtK/2Hc+pBM6uJlESvemzfcu2kgb29qH+RxanC
Mq1QQgVtLdtQJCmeHzhUEFe6NtVI1PxA45nUgWY1/47mS4iDsPUjtGkEyyUa
m4fHoAR+qqdoKXOzYUdmRFaUEuqtZNUIxES6YzCKam5QQClJDXNMUmj2VMXQ
msP/HV0cHv/5molTpPI7V/TsURPRnlmmeAr3j9FZ1X2wHT1joDmbkodXFT1C
LX+6XzGElhss7yY9CpuB3k7EsSj2c74c8XQk0X1u/37ToZPMXM1365SVEF1C
97lfQsNKdWJLG5WDJZH7UEWTMbx/YCAlye8svudx24Hse5Lq4dQ0jK62KSAV
MzkwAiHPI1gAUdPygCZpbDDBGnlQoJifyicKTc0wcbNAwCZz1i7z+NJXcmrH
VIhoyhLBl7qVd4xTb8K55a7pH+p7HXgnPY2ovze/kfzvL6VjQzvFE8YQ7yxN
FwLJupSO9+IVYzDUQZ221zUcJb5ZSt5NzJJRLLxwcrmBFb+1JWkxS4a+Eo4T
HhgP4fRX+RD0pkjn3CGXLVNazZWoq2l33UPSJTttXV1IWaFcGeUewuNgJc87
iCIBj5ULc4ALD2vQRvW7WqM1zRASOWU+XfWvGcpTm+2j8LUSqofvlNzrh7qU
cShR3dQdYJg/UaWTNQhoyhzrRQNl0DUCSzOQ2JNZFjShhL3gLaD0bl0I73Gk
O3Oh5jHWkmDOs9qudkrUI6IDscUkq3QBuJDXwG+zi2g2EzcOrlOVvC9VYk9N
nQ69eKqHj1z/IEfldHwZyXzEyaJjKCE5Nvml/VTq7O3bpmBOPplD/8MPPuD0
6V89qD97/Mmy7DVl9QbOAGQNFHJwsRzGySd5cHP+XCq37nSA+JjJvZFozMDf
wvlAwFU/u8r0OZ456Hu2Qlgv2Ml0imT32t3MM1h3lGwkdSf/1F558G+jSbh9
h54C8wj8QGb39PpL7tw/H9/+3Js8IeG3AJaXFoG8vFC24uJvbHZ4eJmLt7Fr
ovdJrwEm+C4YdhLaYCiD5mpIzpP2/vnVoKcj0kCd7gSOnBXbA7RgCC94+IdN
W+j7XvOEMv5nhwagUXXJDFkGXwn0WzV3oYO9PV9ipKZEpUTUbkPypBYqVr6Y
LKZF1o++7X1FWNPit03dbMT+Uq7mq5cY+4ijGksMsTGWiaY14IaiUezJTbgw
umEChNFFBYCEsf1+qVjl6uRPgq7S+YvnPeKU4ZaFGTOcfbLX58n0pyBv5awW
wwhMNTNwl9fdo8X0reX1AQbuskzNBrKrGm0nZfBEbcAPespMuGxqyA7lGt2d
4b05WXkzMhtwshJhELptm2Gr/p4Myj8cfyUT94T8kcDVMn83NKiZC7xamb4e
ZPepLaOerY5i3mwYa9sVcb2HvgH1c6Ad0zj7gvI6yGPR6J6wJ1NwOB8QTqbS
R8ZY0ZyMzthWx4oIqWtdxORBLc0qLjLENemWQoPMslIQ41lzQ1jUoc5ZRQk8
sdLmWJOWKZPto3eV/3VnkgXYeN1BBh4G75M7/kV89hJNrOcX0bO72WGNhFRT
FKNLvRbFBOjv5hzuwjYPY8ih8kjOgT3SYgVZtNnA71vYW4MTQhYVsnEb80Bb
NzbIw9uxQ8eZ446XKl8e+YnXJ0YlzYv0Uzixl9s/txDxrlbbBpgyBkM7xxfm
y9Tyo7/i/PMI3oLRDwx5iaz6+aW0rLlZM+k2G0dCbzZWDG5xWfYuXMH54L6v
HjXOqgiviuFSub4Y0bViYfahKGGHTw+M8/MzWrJ5vQEWldfRnU4/qIxiktVz
+Q4kJwIWyzWKXO5LVa0S4eaTlL+jsB+9Zn3LudSTbIuBmbeeG7y4szjeG99q
fK/JDNRi5mSO0ypXae34KM5FGTtE5x8XVMgtDeW4wbAMYK9c/CW6HJdYu++3
NhTPH5dIXyiQi5EFpZkHDdjLsXS2JsFV7A61IYqSlT0gVV6qB3PjcMnPVdIB
Ykwr/mzE6/xNcy8ZM/0gBomiUq5NQGi+4/synFv4elN4IPPT6k5+CGDy2XL+
jfFFwa0bzCTeG2wDg83JkUsw7B4klCjAOKnXlScxW6nrYrosoMU99W8dKmCq
srwN81Rj5zbs0gvra1PRzpTdrGecLTqFjloE99MOWRTgJgyJ7Fq7QOQ3pHIC
uqGp9UFnkqKUM99P2lYwrsgI5EihTbWcH1vY9ab/PP7pUOR5BA8lC6mxQBVe
ogtQEqjDuMnCBIVsWkHknxEDwgudjQ+eoVrbbijC6hZ6H+egbNXLjDeE/MA3
CqaRlSX3zv/0wKhfPs5gFDAhmMsatOeuFqZoWKX0SWv/cC6xgvxfKuvwdBs6
TujPrRsnPHGG66QKXEq0efHjUycDWnSUxEygbMBXyS/+Ps6XmfvHHARLwL6J
QWS9JAt8Z3tr+eBVDeGIE+NXg0qFiwgAl/oFNfxqHUN/8pF+zaRA51LGxgtr
WNvt10ks236bb+jTd3SLl29PfO/64znJsU4lhZozZocC3G+o8DV6UTcxxDRh
q3+uihpOS0ZhbPTHuSvxG4pn+GgstuTl9lxOugZAfQrpJ/rV16w0B2BOk7wv
v8JEXbfUeTkYrH7ynSamCcCATxevqVePT1C/RR/L64/i2V6CYaYtKuV4/UnO
JWS2MTwiL47WmocjhU/KYXpGZpR9H6q1tqzy6TKrjoGo/ur96n/ls7j5CnbD
gGoTF6xXMre6SHCGJfajV3oJouebCjhYHy6bxyRJqvTICkjswu1gygvZsmFJ
1wY4q1GCVjkjtCMP6PT0fQ4Ng3l4ms44I1WXbmPxzIl8MgMdqNYdBERik3+E
abBwPgwf85kL3xwtWFq8wqH0H9VSfR2wIwLGf8Ipxe94FqKE5R4ptpRJ2lsP
veo8RUZU1YHhYK8cSHOaEJNRfkT2tPlhsZ2r02upK2I6vkbTg6+qJadtnesg
kLbHYRDSTwi1/uCPLrCXGq6Gyzq29NZILRxjCSvgYUQ1cDUsIBkOge8XLQeo
ozIJ4f9Ev5jtCE5CTDA2XVGIGUE6XsPbbfF2MvPTuBW2oKCCFbx0HjNTjTmz
qvgbU9nBZtSp3FUJwuzI1GCtlCt2NKrV4WjzuGu39QrHJjDR/Q6YFH4VENcU
MRwnboxztwKaide2xC06U5EKP9eIDM8CFwF4A7AJmlsbNnONUGLme4t0i3ji
L+oap15AvyTyB2cDSf5+atG3/UbAN/+AtVRLfDeymdqGFhDC5D7u++inb1e5
qe9h0Zf4AkQZQU5G7zTHQU9qCRJKeqAF22re5UoWjogtmJd8VZUjbShDjNmF
TB8EUHLJA4ES9/cNK7nt1QMbr983cDxMQdYebV5tZ2wRmhQwaRLCKpY23rwZ
xAG6sUd5SS4khj3OI82p7PaJrwVOOWu9TyIcD/lhh/f7D6EEUF1X/u1guerK
KfwLkKETEhI88cXIyVymwZQ2FgGi9BuCKapd7bRWdnm57M6peK6xCeGrtSb0
XRScJuRCRWAIlyatNY4kf7VOYirbxJqp8rJ4W/XeRDqnP1senD4g9CLT+cgP
HRydz3SvyB8zXQzGuJplgS0m1Q3VYynVY+ZZAGI6u8Jm1eeFBSp6n3Bvozee
G7hoxzwgguv6862iT8Ddp/I5hGl1UyqBP90lxD6hAZVs/az7gfgi5U4It9XE
1LWunTCpXRctQdmyIyuVPbaT0JX/r432eGL5lTWP5g7wShO6owd6oFylxquR
R7TvZoh61epw/5opEB+e8EtlDfsHM+wUw6I6EAatzd0vmtr1oFYqQybfoP/u
3g3xJOaXQAIDsjbxoTwKdd/358zayj+pSGmesiRPAZBv8XBvk1QVzsv2Nk4K
GDDFDZcYVsFUh5d28Awtzx/nvMVlMWLQWgwAQzEy6eJFw5R/S9XcOLgicXWt
+UWGMeMuP9+fv7GUU6RVh2mca490ODM5h4cetFupZ1JdtqEMx0GRHfJkFNAg
7gtGiOkFZ0CT81+vRebIfgfrQ4EUyOaK3AKUK+iMgK6gvDTNWABVCh4EtXy8
b1iT+wgAvWR6xvlz3HBReITGbbUdLb/47x2U7R+yTcWP0U95Hzk25ZQ1b2OD
SKUNB/DLUeEyTKSZuqUxx2WgMHwZaYX5IIkuRqP1jZirDle8i3b8eWwUORgs
Loxb5H5ipDupFSZXm57nVnFM9wg+MEYhFdze2KrFtNU90ZHH+6tYlXXos34m
ss6msV0ZYqcxZZhnDNPoLt9vdT/DZQtjZotlbyZOHKhbobjuneCgSxjE8Lkh
Vb+WOCWdDYkiQCvY0WQdO6Lr0TodEkEDKuYKKuZYCQfPj2Src0dkTxmG4jBy
z+w5HpTgdG/wYEWqilpGZPCgyxl+RWFtT4Aecd0eW0dk62Ewc/onsMuoqd4R
5FRXWb7XUAIKm6bImKbdnHRLxL4sg9kHyxbXc/RtQDR5F+McikqMITRGjAwI
yjzucSqAsxV/34xJRIrimcqAfyRXyycjiL/+HH7G4RwvDkfpUP5+vXUoYfuw
t4BcqpztR4F4bjWMX8s86k+3ZQwiFqqE4PyRwJ3aoqeZaC/9/tYKFTGaP3nQ
XrVubKo1X45FOAGlbU2xE1R1m0Gn6Pd55L1n0dNyKfQ8ZvyDdjMuIO2JNJRc
YlYFfo7kO8uKUQgAzuq3yZ7WkixiM0B18Pb2fI5Zvl3hHpPZcQAlfxkp/oBD
A3WEdR+0jcGHhjRn7KFNHalLs3atto+i4dI+rJEdcaS5B0nQysGP2eVRx61h
Zj6Ox5S2yd8Xr0xZxJmOUHMgB8C7WeqVRHWS/g3KVeXbWex2Y13f6nkTMjQx
JuDBpBzH2Sk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1L07IUn/bv8PU2d2gAa43zT6gVNBdK76+fxtlXiGvVW//Pu1s9AjzotHbuws6ViuTGJ2GBH4IafUoVP9uVYHtJse6xrbWx6yqbN/+zAxG7mgwriI5C8OXhQbdy5FfTUr91easMWM2o9QlmUFzEqMiaeso2UV9hUsSBhcJAjb5OEQ+pmLjBQH81EHiqpQ6lrzSGyUh88YjUtKKnzdToXAevl1ADedxlNkdImL8vcpmMuJj25jWy+UxL6muAgz+/+S/m0Hx0Cck3fCBBCNnxERsqxVrqdLWguqpemKc6whwr5czNZ7Ignw5rkwwbFE1iGxZAtjF/r5e8QXu4uvcJB1GS1uJsG3ExQWYQxb24ljgw2yITds6xyTxCUCTsaMRbNZY/Du7X1CbRhw3GWvTdYqRLWK+DO0i3Lz1jznd2SWVPhMcBZm7/V3Ch6/AOWwsAtlvyXarFHAJ4Ia6TmEWlo/657wPfMFCB0/PR+EMRllba/0Q3z+5WmaG/KnPelkCRblfgzR+Z3/of+VADQDxDDGwpHTwcpnU4CI50yxE4Lsx6A525LOIsF5hRRBBc1Ud+3Ue+RDwDvk6OjQz/RCVfsptO+cgBxKpyrHtleTHt1AN6P3mm3j9ZXMVn5yutHByt6GaHwGXEofQH+ay1T6rscBRr0fIljUi2G1d2bJmpIQppcQ78CqH+yo2mGf66pZXOzOt+cXnPd9JGPe/tX1HWLA/4GDyEMg6F09VMzXla9qgJxyjJGLRGkL735ACmcQZYKQYyOMMEofz8xuHf+jZUxrB2f"
`endif