// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rIdzbyENdP9YldvpRZvlx53wEbFO7t5cG74UQB3ums4NPS9qFbgUH3dCayEt
UmJApgr635CREy1/RM8uga5dKDQlWBlApMAqNU6hkkV59x4Y0wEZrEDnab+r
rHqS+ZRPhjF1sWgL7fE3fP/1qQkTYcHD/yhE48Ckhm8mb6GPAsxQP4wZRnjj
qmqW8mYCgZTcFUzuZllY3F4AWEQ8yL9oFvR2mG9mTDCIrrQLzy5Y7Z+TVU6e
HsVeLR5P4xdx+b6KC/6GIB1QU+/ukRdibigkfCLOL3AAdRkovqr5uXJ4tkNB
ha8xlXQeP1QrOS9Zm8rDRoG7gzjaxDH+BakZZCtqGg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AqHdXOCaLCnOiCYFYByMlffDRHU/kkh9p8d0wbCjXLb4eJhSg2tWI8uXLZ0z
o9F3ncgbycR5IP5LgFL9fIggbYx720xIJIrbM9XkR8nDGnq8hnqgIRdiLoh7
T7Rxtl+0kKUWNOjzlgY3FpOXKlY6UfdsLIDnuJq9qQb2TFCqtMT+uCfwwNmF
2sYacaLZY1jibaroUPLMRL9N+mvQWHdfaEHLX+6wlaiFuTSlcLebKhMm17cR
n+FY9BXbK0oOjFNEtKBT01qS1669W7/bdBOmkmFP0okm5zU78FV6gxfZ82pM
3J8mYv0rUBcFF6R784E/6cxWhkDM5FUcEB7jnY4+mg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V2bhFtxEdLtKaIoDKAUeB7mmo2qdrSM7IbbZb/jrbHJ18kOPlGlQKjyRkMtk
58TVWDobMNK3doMZzlnolNGG0020PBUcxkfL8BFTREfG/rrCND/AnB30QPY8
Spz8VMSZsBvOVSUZjbvSqRo4/b+E/mDnvQEpNd05eWO8UfK08ejqrk97pryt
oDHpv4icCArj8Q57LcLYnkWgziW3eDeBZ80ezS/VwsTR+osHTn5s1PNeeVNs
zy+X5Gnv2JG3vlnMDfLD+zEeZ1CHivVI/sg949AwUKsYbbcJ6Fis5JSLlxbN
t2n0uyqwOrgYdhg653AAXsKuDY/shfwKn1cMnb7miA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i+K0x7ZXL+ejf1O6J6EjLgkKLnXM1RqKww+3DxvUYi6qaZL5/Xw2xJ4Giwik
wno/vSyQ+wv3qt4ERUqXgc2+pieq61uIGL8w+h4TqE9/yL3AQZJYrCyJYYWp
Zwn3D5kcWC8vIMXIXWf/rP6SCyy6YI/+salJcZ7YX8v7WwkQb3ZnzYpNH1VU
tZs47E24oO2KZG8/DWml1rfwJjctIJzGxEIqW+axlDQFUahVY1rWT0WbTPu3
wrXy7nj+43Dd2Nzee8lXd4+Rq9f6T6UsSOd17YaMnUMSca7APqJAic3+tqNJ
byPhOBUci9RpCRQm6Zw+g5oNcV+B2ixrME/DNepwkw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YdWNHoj1HdvK8bPOcOOEARx6uhCJdAMz5Dhy7p8N/k4M0VlvIi27w4G0i2Py
+HNoSbV5VR75g4kdSOa6yM8aN/HYeDQCDaUGIYNjXlHEa6NmI+oUznXG6CRK
oXsSyizPoxyGbvh6F9VT69j7dyUysJHj/X2LWpwwQQOwvf4LDf8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
x7pV8/BcNOfrwhMALBSROvIoJmn7oslnEOliHQCnw4qMYejCUer/EXORco7f
eeIW+Y2v7Qx1HoXdT0tjbrVrI/oOENbV011mN/Iq0VTXDSUyGNaFMeTwDwn1
zN+py/9TXgV4s2Llm8iWPwQg5ulnUGbs0f8nx6FXlgF2tgEGpTA2Y2kqqojg
N8Vmh1TFP7ehq9p7scGDk2Msd5Oim0mkPIQ9YJl8cSFYE39zOCrqbNZLDBKx
g7nRJdOikBsSR2ZcXG1EQ9/FilJFraWwhzlA56zW6F+rURG5m1tOAdUFZMbw
ne42tDfjT7yPeQBaiPaFy10ahLcr78X6MKMbl3FY7TSj0Vm0p98/cHKFG21E
iXbvwkQ4+/b2DYwoctFPy/Lq3uiz9hUsFA0SAk21TVWW4tYzZfJIRxc7BZL6
GJvsd4DSB4CkojKJHA4T3652oZPnGLQKU6Cps97sl52qQmiMIc0sSvL0abbU
c+0X/F9K7q3vHOLiDcflM2CKLIAM6tGD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KsPokpN4ofJacrsAdKFx0FyIM9E77JBwDyheOPP9tMahOkXH/wkS7D7JelzQ
BG4cbV7MmVFKgqWW4zQGob8FOJwuv0M9gKwgQgI1Y8yS3UDbCE3cN1D8iLvd
vx8PJq09QnPddS7rw4iUQEGSYp6k4ocf3/r84HC5dc3ZOaqRs9o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cakISDic5SvK0rXzeffYsS5mYyTZhuYNybmZiV0+vgCzyND8uEwW0pQv0Hz/
4tlbf1NSiTDe+aKxxjnSTMNEsVVCg5/vyZp2qYuPFPkXd2xmfRzSwpdu4Tpm
8GyAhe3AO2/lVMJr0gq66RIQZVLd90iKpJ2oZw0kU/9W/T7aZF0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1456)
`pragma protect data_block
E8Ecsp7ltPLwYdvAbqoOqZz192JPEjZ0MMgMsKZvK2mtTc1lMJtt1rqqJIeC
TbIdlQ2lUFB4+bJjqyTTpmPy17hWZEUVwxE5lLOByfXzoT24CgyoWx4/Ph7h
GCyrWOXeSzOZeKUHZvw79dEWKvDBTCWlxCbCX0g5Aiv+PnMz3Y10OgB2tg8O
v8MgmrQbuIB2kt9jzdTiLZxs5cMORfxPKek95x6bwlK2c6iL1sjY4YQ45W5U
wfpqhQqkzgvgiZo3KqctoVto4QYciorUfUOyuGW17/jpl1cNKaYNpp9Mm7A+
Sc3dM3tIj+6oX9u/rsdOl9jglhEOLJwl55IX1hDR6l2FiH/RR0aaRkKd4IAD
ouwDv6gdpz/JOndb0gAAj7PyCpEUa2EISxjEkVauu7iV0x0Yr/Rz0fyZEDmd
P2lK1i/csxEr8JSZ+A9UEeSZE11sggSDBG4tEsaD2tt1CMC8VdSIWXHDrajO
42Ve7FpASr3iDkZNI83W6WXFEj+ilJHVMrgEiWM1zmEhCnw3tfFAydBhYz1h
1OUfl9pnlXPuxur1gM9wmAwc4X1vsLnSx26JFnNNvttKMzblAAzf6g0ACyJt
K20yB42IWGMET9kKjjFxqlpENkHHX7OM1/1ALCRqFODSQfFMgyi39KArJwGZ
KJLM4dZ/j1YvpftVH3bGovGPSXwuW3j2smR3NwxdHidFu+adp/F+xOnnPwUz
lxDE4uEzT/vVCsm1Ouzs1IRe97VYicoaxCRZ36nMaBaHihPM3Fk4REXMipJL
Nmfl7kQztnE7GGGubh6/nryi4O41tKiTgpY8oEZiMKIRyBVx7epJU1HSgcio
EwBcygrCdt2nmX6pmIeFoEYqTapl3+wDtIJjXgmL6YESSlLXrPRpf2gQ/6c8
Zv/wFc9nD5V2bXFTRe5KMYE6sFTJ2SpymDVD5vz6waOH/bwAx0zPKSVriOG1
6WgIMDfIb7P3Avs7ry/GMOpw3csTR2pdD5S9ZEsRatzs8jv9R5qAs+9/PxJT
xf1bs/J5JiAA8cPfYei2eVNJBIz4qRvXrnbYp+AcNX/94RMspOqvrqyRBJ0K
2uzLcNr8qWHitKj0Tf8NtUYayHsB8Ep+oiU+oy2GVEPAI8s5aT3sy0hpUFsz
mnyrmgJNL71rQzjgenQXbHMqWQ6xFBzUZYRt/urdOTJ0k1+APJ3dDGOHwoHQ
CL0tXdwzc5qQY7xKXDC0lv6Sd0ec+edtT76Eg4vf/0uhrADKS7jEr4ArIMTY
ISqV+KyIwSO6JC9tUdSXomwHzl1fxeZYPs38HlOe9A7zxYk8+p0ekcWkm9DT
NVB819ZthPeTM32jAq9K2OBXbkQYPRu9RHJj7u8kYaL+fJSnzdo9/c3oTiDC
tSgVmR4Tj2EFXumkt3/b+yqNkqpvB8lf4SyRuN+Pg2Ic7O0yZlg6J7qFEO7C
DzB54QSe51qbTgAa81fWgsCGmlq/zTDeT570DXEPUu7mAIopdQd6An7cjwRI
EmUaHboGCBvMuL3T5Ft8H68697DgbCcQHYc/zFhQ+DTR+FBZ/thgIU5CDHM9
jZoELe01Oz3LM+4/ODUIAEQFGQ9mUIidWXU/kYRYeoGsLE+xpxUKLwq3JGDm
aBQPrYdzLjxnyksh+DlABRBGdZNmgbxjyzx6kcAhVGluV9i0N7GGFjnfwefy
lqyYFS7pRoAAG3sJHt7xe9VaGPeBGyBKBXcxSTdnPHhYK/3i6u4bx+aSkIsP
oyzg7/VYq580JhtBPEuBdPwie8HhcAfDzhnvIBZbfovU40UYOv9oS8ofIESO
Fvm1/i95pAs/hXmzs0pQIjfo1QRNvVlBZzmm1toNChxXjiKLjHA8gv4LY4/L
cXFSh6i0oo5x8NeVvdXayA53YhZaBTQGZVyeIljttEAJA65cB4MpbogCVbCl
kIWqBFMbmjZNzRKbnavNfA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdeCn11wUt1B2lBCFe6kv6tizo21JRo5ljtnf3BgZXdNeQWAszMTm+nxvsD9bE+Od01A4Z7Dm/9N7iBhbUGxdTtLLYNZTONWDkwviiifow+uNQA9qarPO+phlQbA3/i1YrsHxw9b8MTC6YKZZHJ9x7ZiSMekpolrT1sKoVwYHG22zErsuJl5gfqlCPwZ0Rnp1iOvOzRV1FOqjjsTCI6Tny2PRfOO3GqAyxnpOlgYLNFhmPSZP+NDa6gfNSsiYHuEDzm7Okg+TfaqvCBFxXcN2Qn1IMrR+INzQdU4ZxdQpNW/8e5gVzGKjNzznMaRgxl4asQ3GvLdwCA6M6j5/JvFSQP6XMn4dVKSnA6CqL39pDexB9n1QxbBTDx2inGCTSGinitrGcKJdigAxYPa6yNNytbte1YnhxcsGYKH1VEx0OobW7924y9jpaDepIBcY8hYrRPl5aHKlResaf3f5YCpWG1henuSGi1Zo9pzhlyD6gdCERt89FBwJCRJHIWY0EPelkZJ5GcV6c8+amb0oC92JbJA7BIUUH8nTLQ7NsypxOnxm7AWiLGcLzBkBdR7KCewyjZztBuM8FlK4fV7Xc8Ko+BNp3XQdb7MWT4rqorHwSZZHISrcTvsidAxInuBfEEgeXRdQ/26kbNUmFEa+waocvHFcXiZqaQA6waSO9FWZ2YTAqlmPCZ9HHnvgJIQpMab/6ZHCNJwkGiFWCce0d57kxOeelHyYV8V8Qh47IGD6jvGBg2TPwX3rWK29Ecn475S++ioJ1LzUq5Jx/0oxnpzDOE"
`endif