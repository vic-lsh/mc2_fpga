// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QI5u6iAYS2mS7nl1Y3blHZQblby239kU+h6oDHOV/geqOb1Yna1UP9hrdS1K
ca063abvGsF+q2/8ArAysafSiswbTc+ta86Fj+Xr6XUCpcQCvlSDlF4zmus5
7NEXoN8J0PdjS6fsSHPZFesPU66OgWPMPHeFWzCxxtLYZefXgWdP92Ngk30Y
2Pb13DJPcNllSBCdekjebiC/7+27OhLKslhWzZXh+YL/T2zAKLNHDgeUIDyI
zdk4kc8ZdVJznNCFLF0smD0J0NGOaXNLx6i1B2fLLsJOcjScyamXOEtijsDa
wyH3KytBGonr1zlvtezkXyClER12vp90SX1+lnV9vw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HypAA5tZsePLown2a8CmFPb4UjDBSMdqqpPLYlb6sH6S7JZKeeFmBDRAUbEO
MqKYLwC3D2X0MFXXtsRfbu1xMqyWUV4KOgxeFNc30XhP4qMGVUU/jLQtzpQA
fiaqgcB3ON1BgQkx/ND2qpUYNhwXmkRdb9qy1AkgPzQxa12WLU8Bd+XB1nS1
Yjt541eA9s1G5wcxNAbGgANp88APVAghOIOuPI9aw7C7cT4xZhzNEsOk3+G5
fFlAXj55wj+ihtYlLeYxS791F5VUp7TyKw+Kn/9eASVrqoVKfyndsTR22LVU
BXx2m/irtarRqcbRXsDyfBSBymjcW1tqEsCzMTzSZA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p9C6UD5+WwjEtstlWlBOll5tnwjW/Ob/jaj2AH/UEgOiMkAljwQW/1WRYS+P
Qwml6DO+VQJyiVr4uUJGV7diFJg53mbPBGtHsWeaaTWAS+NPZ9A/8zFVUKlm
5LyAllsXxQSiWEDLvOLy4ZuIecScIh890E1Zfu0DEv3HB+TXLgKhEZEdVE1Y
ndppDeTtCyKmYIXeFWyjB81wko6ctdUKXipPjiPz1SktEj5U4OLag4ZUaveu
tKVaMPTL57tab8wiwcXM9O8Wj4m8ag+99fgxyHTnPe44nS7/JgH4UaQaGvef
P8uvKdFZvjAEsN6hTxqAuiinbp/ToUZAIPYpDu0grA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gIplbh+fw+d9saD6o7U51T8xwLQMVy5e5+WD8cnUBJ2HTj4Ni+KZ6U/a7xK7
3DhikH3CWMHz/xJYqyW5OCnwcwrvY/xfqF8pFlZdsYGeoEK1M//8vAwdah5+
3nSmLedSLIBA115F972oWW9SJ8vfOT0uA9/mkG5k5jajaFa6jLXre45v0Z/T
e8ttSAn4oDYfmZrZRpRxdHSeRnpFK+1+sdB/WPK76fMsGwU4YIur2zjkj8bS
X09V4HTvAOHJi3sDAGDBbpQ43V0zjoItm7Yv6c1LMGyBj321oyONeBVWntC2
pmuZWZ/beEZuyiDE7T8KOA1cG5Z2Vc+mUVO2jXLFEQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZBdoGiGgYHIE22W/UBkdcPDYu63K9MU7R4yp5NkIr2w1Fsm6Sfnwfv0e9p2E
Jbf0Wn8wqS+9+rah4b+Ewh670pDA6Bu6uhp9XQRk52skLlGMByEVxtzRbWoR
mDa1P0R08uKOpc98YHlMhKsNwnpHurmqF73VSdci92qOe04r1cQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
fDTbkrzPbhZkblUIaH+aHxIgvEwe4/88yD4NuhjhiQjPC5f7xLA+znLeM7c+
UxxRXhd22xViYLvDmV7rv5FBYe8AKTxkNKKEftOX2JKIUgZVOBtT9RyCui1q
jbUs69yyc99FDfvPwcFEXmrLfqtIiORre9knHFdh5bnsuYmy89pK4xe6ogre
Dc4zz3yWLTUYNr20IKQFogjTcNuqHR08+fimil2qWaKJVP1/d+63Iyf+a0q5
1tqg/f40DywV8zTia1bMWnTy+A+bRMaU8GKixPKcm/AnicwZruPsX6KJELhW
Qirdj1vrtWSowhmds5Iy5GMnkgXqWhCo7PYy7p/In3tEYdW0lw6+IE4YzIWY
Jeuc+y/XEPSkldw1pAe68V8KpfmwWz5qo3uHTQuux9MzlN0K7Uxyee0LrW9m
1gzBXq+R/tA1DABAzNWWYbLqsWwy6RK2+itSx//IE9NBl6U0JVUYy/tefsSV
PB3zu1gLxt60PEulAjKoLsz7cSwWIiCP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gqM15BOKHK648TLIqY5BF+Pn5LhilkYQbfqWVIpRbxllGrXhJvMFlVOA/M4g
Tfnx09IYlAcwPJQIHcNgUpERrqXoxvc22PtasXelQx9XsUqlKOn3for2iilB
x3dl4lB41nl6QRIlL16oadCoFN0So66LS7JduRY5xvZCmYjbyGM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JbKDnZBK4L+oqUr9EuqeQBjqTi8OcibkU7bSYcl0m5FnO00IH5SHxvGaXUph
rk3MOQnl8LlWxB2JujULluPre0EetnnjM8GpJ4jg4v2YmSTyUMlRD7JxQd0C
u5i+Gg48FyOlec83sxamNSPjTCbnjcP94CGIgiocjpjD2q1EbeY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 29696)
`pragma protect data_block
swgo1PTvxjQHBIFJcQ+wK/4f7VnRu76rHOEbs/f0gEDy6yox9esmRm7Tsv+W
XcvI9igADMJJp+no8aycVcIgjfVs5VJz1sWE0pKHlOtEamm3trx+eMZzE6Qk
LW6zr2ZzCI3930Zi6ktw/qBmB1qBaCgOzvGJf9xUorOeMUQx1KimmWhLVRMR
Ku900JqZERTZZXpqatglrEj+f1VgYuIG9l9DwdJ42o7/UxvAManq4Bfk39rL
hiXMDBi/1w9x/ea2jHnW5dhKW5kZMfs0zKY8JXBaw3h2bsUf54mmFai7bk2s
taz6bBJdw75yc4ZtyFZHE7i7GZVW26l7Jl/eEayngwUUW5tz/87QtKrtgrWr
QqtjuTObJqpaeUX4UQcUAZiJwRXhAQdRfRkqZsuLKUx7uY0mrZAUmkclGSDr
n796u8toFYmUEQt/ocmpWVqcdEpgtgnqEGsiiB3+pwdbQrFQlKp7rFl3fTIf
6W+pb8msj8jz8Uab/MhEFvliCrCxHtb71KabcBMjFrvRu67pW6+7zSRPFiVw
2AaI99uUP0kn4dZJSjDUE1cJ2Lx/MOOp8n4amSDSX7XjZibUBRhZJoMtOGKg
OxN90odXGm/gISy/RSMliTzgd4yGyJMCfQ4cS1Ja8v9N14vYI+M/yC0b978Q
VtX05gt/xy8bbain9fT1cOGCiwlJMtRhgXLn4gFJcIBjgdcZliZWNPiHauhk
PQs/iCS46oS01iolVOawpVYN7fNk4VXQFD1HYLjvLyv7lH2ycvvobvU4qFzy
zY2qh1sOl0ovUVZwv28Uehot5Poyh2iatDYYboLB+r+8vR2Vd12O1ERI1lKw
xcqzHfqsvf+SYspWk3JwSlrkw1KwDyJxPxFU5S1JSOdBRjl5zX7g/tVauMWv
ysp3dNXR1wlOFK1aqVEdlKSrnLzfFrZ1ZmdKF8VfOyXMi9umQjvtqzjscWp2
KqwsQVVl9x8yk3IgYX1tHgHPOZzg5BPF5+yX/OEPvgF696pT6Mq8i4EJ6yY0
14u4avD8SnD8YKLWPCNcdhY5TS8dIa6ICkeIP8AE5/mL+dbMJYxgZXpWGf5+
esbtG32xMrQl29GmSxCPOMm1Fqa7Vg/GjpgTn1qX22z4+FbDBjIx5zfBkXmH
GkaZ8BG1MQnkQsBtz4mGsTb7sUl5I0Iaet30Z9Ea+QKWKmURyzOphYTlKV3a
jCygEtPUOwbvHkImnV1HrwA2/VTwlsMVDsdnYGWU6o/fmA5pWgxbBgq13QEh
pHTnFqVD1qj5wSGxynh4X0/w2AvE5qOi5LXPNCm2ZNgk4imKoagLC0JB1aPr
M/1J3dv8BVWzWJ1ZlI6jFDPNofAjArkhdxmnXnzCOJXv5Abb5ZH8EnsYUmQ1
+q2GyoF5EayKUNCkAJ1vKoSom4n0e9vZlb5EUEVQW8n4ZS6uWMZB/CKCSGaB
pgsH2TrMIMg7FGP0IZ6pxQkisjA66msZBIokPJcJl4F/oIZh09Lq6K05hWQi
lLzHNfAgSa0b2oTKvyKj13ItFELoJPMBnlZZ+9iY6XFwkMggQpKJEagXfBQ3
RDhWKNQmQERV71LXevSUJevwXB8dLwB2EoVWLeQ5eTvaR0c0QLm7c1PyVYEn
kBZDF++RtqwlP27ej7LljMi/TNiaIg0HXw1Af4shl4UBSfZbtvmSwrIhy5Qy
QMqOLlNwWNbqd93wMl1BFw9ynMZNhBErvd/CTSjnzlKRc0I1wXpTIx1QiqjD
+TYpA8BKaE11qOqloN01E98kOthxqB7Oxm/3Xd8v8N3X1tSguF4D1BObhI4+
PBOaf7sDnPjOuwqLug0XSjqcfspZfxfZ1wxvJSjFnZdc09++aV+ri2H6OlpC
fWFYmRIfId05OjzcDWCqJjbChmKYK68V3aQR6QsRIsJroA1JyBAeh+fUvcaC
HAGYSCoPohlaCcdth+YC5aPLYhx4C7gZ065YAqg7e4u+gCnAVuQXuf/t0guS
azDrv0IabAaEZmHM4G1uNOjm5GaScm7+CEsnC2aI/BWTFqei8eOqMVMKuyWC
LnHni9C6Nddg1i4ae1ycECwzxlHoqI0YO5ylBwqUboU72+2vs3BBRYwP+wtx
8nvHqaysHbxWu/+JelmzDlPco2D8N+ZEKRNE2JgXh6GHSLLJV6TjY14uNE+X
c4CtSh0UX1YkTI/FMmzb4+hxXBfYJ+CBAloKN56lmxPMItSaSzxZNGWmDyDU
1bRAfX4nHyjmVYBeOR7U2SunpMrHakB8me0fuVY1PhzkVAlS2xVkBfD28piY
HgdUxwlR6ts/36UWrzbOi0dg7rzf4zmGYApIVqgFkHExewliUORX9XLDewuK
OVnMBBaZWJK3CMAbJB9g8hs73rkInyaAO0YHxV+sNXB54cxWsSiuXyH6q2H8
/oSBfxm/bWDt0Mo4KrVRjTHoTV+22jnIbI4+nfGBNvSew6UGp+kkf9Lw22PT
+fjpk35EISaMjWhVyQZmQgdAAt2fDr+7PYevpVz2DCE9iyu6Dl4THtrBiR6O
Bn1PUSrWXFPoAW7MpS49SfZdyfIp7xU/k5sxn5OKgdFtfSvQlOGBlXtrO16D
cRnsRnG7qyjmvaWlcr4xEaXMOkWp/U7GpejYRuuqMVkOu7ouyCikOHNUitod
JW2dfcgn2PVrYYOvcDiWhmgmwrM4eFOTNKV4ct4IIStnst3umHKht4L/VWoH
cpSVpL7JnALxmMmap7koHxiEbRRl1jFYa63kqywKQ4m77RN5wH/Lbvhp/rzG
ycoJhlpUJhXmNxqQtsOFgSF3uckMehWdNHVxc7ObcRJVqH1gJJ7ZzRHYcqII
aDKv9YdzwtuHzWuNS0SWXEPsAV316sra0U8fmlKvAOcHoSrURF+4f9WKxDvA
A8pJoJCM/zLnQ+fVjVge+NM/0H6tBKFTbobhMgpcQH0MOHgQiA8dL7ELCzI/
gB52oSg3BcLeePtATf+ksX2xXH533ySVSBgEBp8xdagjLKrSmCR/9HQG1nNa
fJKrdXsvHx2Z6OG/QLOXKsgxBgL5oiP42tjyuYuGojAh1CFIkpW7BSs59V43
deOjf4/W1wyElKivKDjqFsf5qignz5Ge+ch/OF5CekMbA+8o70B6509IsyXw
MVF1Y1gUmhS5m2vpPZ6C0a5Dk5gZsJF0deHYVyt+krxPsHixmW0YzzDirU/Y
xVPvcqSFGM3qbnKnnJGGmP3Hwyo27UAzRGD2YIWatiZ3p23fAYPLRNbwdD/v
9A31b8PiWQjyuMhOV1v/OX7f+l5fouQ907vPaXDwjOS/hCKO112szc2TXkSI
0In0KQNcj8iGybZDtonDE3FN5g2GaGBzzLycUyJsp6Yms/If3u/9ISAIblOL
A127NBXLPSTxIhGIH3BWJvEEZZVMyIjaPLe3Qm9M0kMl23eqLGJyFEneK9se
fWerI8cUcmXFLkEDAfIeYtYZSwmVXugXAxyq2MAaM8Q2y9q4WzJHUGCh9cj1
GOrtVu59VjXfOUZMh/dKOOx0AnXunlfE3w6FiQS3PVHzoyj/yhwcHHajxHaY
RFT41FKx8Ythi7Ih8jj7bK65trZlPH65QGEG5VR80FjDNxZZ5Us18aDUqIvJ
dHu5CfhJMF4dfGHD9MbnSm3Z2+1SdBHZLVXJ0UblqnzQs1CgX1pbbp1JbD2w
UfLfZ3b0cJWk/whXGF8OLXAvi9klEkTX+bXOl63zkQeYFFwukJc4SN1vpd89
jb+P2rGA/6dQBaYdradjVQGL7h4tMzX/1tZ1CDVvhDx9W8yvMmhLBt0Mczhx
/cAlb/LfEUOD3j0d+nZLpP8GisnGR6ElNHMvAwWB12Q+eqJQiTvZvhRaBXxf
ehaTLuZvLwUvJyFjzdjI3DvgRiLhYnOC2IwyZ1fTK/3Wz0ms7oNqqGtJ460r
FYrD5UnoSdSZ47pipo5etS0KoGUY+Um/IMjdcU+kDmHsjHFbD1nxnxBznLbI
oCIaBNv3eISnTGRxWW95kEa7oXWvjJN1TH1D9QJDv8jHmR5vNM/FZ95xhQne
4liJFhtn+CR8bbCVXGEkLlpf6FdYvJCXc2f7AERCrZbYX72gIqTgZ3XT8T/6
GHTBGTfERnSvsqHKS+hcsXlGyQmLCWy8uPCw1c8jDXYWicjAHL8Otv5Ut0hi
Aee+NSTUF8bSlYvzQBT+SoW5SXS6hbo1gdnp4NUzG1HRbqIhzAX5RRVskIY5
ILPgjOztQeusGHe2rn10THJKVZPlkVz2Pd7TElN3rbCf1X1Vx58iRvAUYmVl
OoD1n1sPpS9dMEtNlqGZzD8xnOPLC0NqmbiUsAcCT2/JZKQZ4xCI5gZZtwc/
vvSi1G8Zlp+ofYqNqQCkinMf7eYmKZDETwD4ejcKNvlfrROMbmWTCElugh6L
rr1XX0MGG7R+na0bVBGfiR0SvDZwRPFMGz3A9fl0C97FogrftBTH+slo02vG
NlMMZpyTp5IoyviU9EAjCqPRTCE/g2MogPoffDruu1etQKIJtDb5gk2JbjXj
5eyMbKqu0d50wuPKeQ4oDdX1tDCRaRpd0p+Wq59oM62SH+QfPpZU110MXTLU
JL3hq/2bL+eTGJO61Y0zj1IoQGGr93l62PrSP/mABkjTu4c8o0MS/P6zYbEd
SgvbF/rGodTD129wt9FvqtVfdYDSASPTuSdP4W4smd6rt6n8ANEOqtUHTUrQ
5BfKRUYlp/+SPe/aKEF9vzuII0VWm4n/TelaMYgH5ee/5cs0UWPUyHcjOmZR
kyfCLkjtxZ4+UwkstqnoCS9vPIqDDgmA6UFN8/XqKCuqqiyCGBCPI/PkZXEp
vLzWFyQ42smA3BYj5akSzw/0m/r1LFvg4IZXtso1EdWZaeuBgcFFgLLk7DOB
Azpo9c5UqnUpDFE5TiH6jr9yYdLm87mWnq+9mGIQHDLmws366A3nUfHLWz3g
khzzvvelVjbhiA/mvPcvrRWv5/CywlED9gbM+qyCzUZP8tFITFHqyuieE8vR
DCQSHtklbcGmyyVT5wYth48fZEH7CQimKgLb78EoAfl/p3LBRw9YHtSlPwbR
3xQy4cyUzTByIlJPdkv/nZoXus8aMWwTTJL856ndIQzFgdh0jj443p3Xd7VP
CmANNC2kD6inVksCcDjzZ48tKirJAcJShulgsUFVGsUTvCZWAymvOQGLlEGR
8PR24O5C3FBQLqld60mT2ahikLTDd3LpY16qF5jtiQnQzIjWibloe4Xex934
UfhY+bRouzLhmRfj1QAkE3bGXInEMEUCsDm9dKyTXBUUgMITQMWGCw9I4T0C
Jpk7P3jA/ptsahClobf0ucvXnuz7g9ILlhIvlRjyz17lXSTHqiz/osb2hYkw
OH0ruBN2JgZ5trvrDG+ktyxSRWlxC7Iobne6tLJrTMwswjCJNK9UFOVv8rO1
zDGsrtM02EdjZpEndDPMOOz0cQ2XGacbTM6ssT3vSyn7k+jUom2HcD7K/3zX
zFX5/YHt2R+AohNw8TXU5CQTer6A+L7O9ZWGOAdOIerpwcqxGxs0exNUJt3O
z1Kweiq8tRDf0s+spz3olvWprZY5tuRxUce2ow4wcXwuyxQ160ExJn9Z+phf
JsiD/fp1rUa8+ihnObdCqhsdtkMzLRbivmKv4a3qZ+OD4miJ/Lpi3mNsuwM6
YW09p6DgVHMizaqG9w3sfU7yZc7Q5Am8adjoFmVJ8zi1ofRe1CxvLrjXG7xP
emPW9cHMZ40dmRRDn3sxU4VY1vmiBf2AYj3s4tCRXOwlplVvyYHGRuStHisV
I6PG3E6BdYxXmrpyhGyS+T6IM6LdTo70dv+9E6EuUGmc+DrfjreeXnUzWBS9
rL2Ynj2I5l1g4X9BMJzE/7t9/uDTSMQQf0wWOv96E4jWM7wl3aBaB9VdMbQ/
Xdst18t5NcbSlWhzUgalqQXCwpHs/Ipzp8oBi4MRlt1mRdA+mqQW2hI5K4ZT
0eeZuXiCIwrGECJVoTqGhdm5Feb2MiaeCEzTICPIQ5fr2ar5g5G6V2Tc05Hu
EoBCKkMVrZjWzEVL4pO4XB3KxWZdI8LdCBju3vm8dq899mvL9OgDBdMlGDqD
4WuQhA/SajxGpsii3hfjOEKXEg3m6uuw2y9zjpML0NSqIVpIHf0q/kpEqIXE
TFwZ4hadu8RRI1SdkjaGhS8zBUW+cfK7wPQe3zM5vaXhV8FDfH4cA7OWCoRW
KjpyzBS38VzaONeY41DP+Y3a36HBfTnGodlf7JEK3EMYwFzF5v8u6+zUI2Hc
jEC+HxVfxsb+O1jKG0qL1D/nIIz1eLXjp5AfMGlnQRu9ChGeXrlb4RNs13RB
LphLGB+IXanM0sp8TrEQzOmdZQ6FKmp6wbJ3El7SpCBKpAXOj0O4oM0HBAzW
35RPHU6FsiLvSo9yw+6VfMYWrBmmHw5LVwc7TbWO7I8hLiT/San/jRMN2qej
98z4g8apGEvuWgh40M527toFE6jeobA1+hN+omhj8bQh6P0nM2B5PN2WIWhG
LhPwSbkczhhiNz2Sy0jPR3JD5bOAGe/2yMoq23pT755ZYDKnMuiu7VUq03ba
iZHXxrgkzLcPMskLGSLp7lBA04dtotaceVLHDcASSaoQEV7udi6vSV/45QWJ
wN66+q3JhNTd7pIqXuyxHcvSH/uHVumoD/joV3WtNMmkRrj8vbcZvY3hXO9o
ty0WVRgKDokETp9q1/xNUEPrHqHvb+CxkN28+EUP/NSLoszaYUK/afovhigd
E4rqnBEvhNYV/psV80ftj8kzlvwufQcaXPJ82lYisdfOP55MHEsZ1a6D/QGI
p2N28TC2Uf335VbJZt/6dN1AKn9MzKJglObaLdUkTIMCk8KKpJ3+bmHv+fFM
AgHf85WkLlFekouoiSzgS/p+B5//z3aWwD5ZeKvsMoY0UrXgflwJrhRYeQRI
Lrj6+Fxf4D4MPHf0yn0IO5tx5gVwIS+UmltZYEJenatuS27QR24kTi8CI5EI
YOKI2WM/5wwYoq5hMVHxzMnohaM9Fes+Eawx6R5oS9+dt7+KMTyF2EOYSiA+
TcRvzt7836cEq0WmtrIhMWvXwexumDqgI9rTLKJjNKiBs75AxEQvNaJ06G2L
xvnb2zn4DYPfFayIX2/oiSqgJ4PxpnKCdLccVs2MBkv7huFGukArXZ2+rxjO
1zyIbCXPqez2gKosZFtPu2Xr0px5axVRGjib5NM1x502nXV1zzhmFHjXUxyy
/XpQ1mlQF2aDObFPehEiEfMDWAFqsTpCJOBas15WPpJpHLEpkJ9iShTQR58w
h6Gl9V/LwTCGrWusJnxYcnsYeauqQeXVm+jauU97uqVq/OFpxl1K4gD27LuF
LL5STrJsTDO57xYCG+1IBq2AkIqQ/bnjhJECR8KQYy5KHYpx1FM8Y/20jZIf
wTrAK1bIVNmibtSZEVZsFyrmH2A1Z3UniF/fcNHBdvWN5g5ihUnBqdC0bcJY
F24mRRFroy8ZNNVJfIfFUKfil9QL6KSv1ZQ31b2XrF8LhiuL0riZNkI8ELrG
5q43kfkozo26xEnKRbXXpZctHq+7VR9bXD3FSUcRFHns6vN/y28JAfwzXRwe
VfUpqDfpHWzNBrGdSthUSweh8Y6qKso88UssDy94hMeHqkLJLHCCEvTZS/UB
/7AWpqrJ06DDj8p0y5UJAd1Eey9jDNrXG8/kfiHj27WoLliTLHNm3gjFEHt4
RuI5SgLW3f7ZcNDobAjF0JNHRiiQ1+r5lMTIg9kS9Zj9NyqPsHgN97Cy8Mqk
fAdASie7mzlvsXQKZW9EcXPtFvc0GzM6hm3IP0NsI7VhDw4q3vzb55wHr9Wj
Fiawn/R5zzON+qmAiN2RuAzZdmpiCz/czxN9jmFZtDVnunj2uKbrq+Ef9WYh
/tm2LYIY39ilM2o7aFrfFNQTZpbiwfZ/3hgBe5b6AV/7ww/lxpEgpClMQNlF
auFHp9lTC2VQRnzo8REhkztyCol5iUQ+wHHil31SzmKgGGL3Puw1GhPAEU/g
hP9iGjL+1S1dSAWpvifNxtXG3vvapaCm0I0CTHo2vzYDrpBxGso9OskfiS/Y
kfilFWuoXZ8jKUWbZhk/Xz+BYA8Tbk6EVZVm2z/uKhLZERnZeQo0P8k+bQ6M
+YjhSmWy6HGq7F48UAusuty30xvllUYmDv/soSROA67nJOZ3hYRKLq2DT0Sn
2tmXwnFK1+8fAmJkrBTSmBz++nEXQAhhFB2lc3Gdxp2ItifOILWtLwWDpd4j
CGwPHKgVWooBkF9pSdTOtLnkdPzekNANcq1FUrf15p+GI4Y3iv+6A8zMVE7w
mqvkjzY6pUVuarlpuZq/TvXdnDm0lByK3VhhAoSu5rDvPUZ1vqyk/cHPGsKC
uP7pcXY5mXu3roJsjK6wXXp0mJHlyY8r9PVgxaIWFo1kGJDOZDy2bKnS3hXB
IEqQUqFec5yLmidlMxiO2DmQeDm3HPNYbyfUtKnWdzQr5pYFWRikuNxdMalE
uUJU/l/KcXWHNDOKZgnBFmQPTWpO0/LSo2oMsuNefEtKYShDHckiulUENUG7
9qXyi+7OvVCtocsZ2tYYYzRGk4a7g1LFWvvZ0KrkkpTtmGMpdw1MHVu9dP0N
BZbdprmWny3nQhO2bjlTHReHjiOfNvpWiHJmK3GXvkNUhcsRRuauniep+QtL
HYpUZnBgxQohTlv5asn7yaBox18LOC4UF316nOtPYVjzyXi1XlduczxuBjR2
YDl/pR6MXlV5niCwqxCPAac8ytel7wPkbgMdcT44bP1J36sgOrU5nXUDvyQ4
iY8uvfq7yaINAZxa03ZYF551fZ9F9TXMSOD8je/Vi06roOO4Zl2X5s8USIlK
AmKLDHYf7yaoz1I8cSCRi7C+qKhJZhBqvoHfKx0B9exRs8TX06+XzsJZKMh0
ymFeOzt6jFJsZ0eif6C7hI6NAA1NZwm7piTzbV4HdTwN9sYNyuDNffMewDoO
lkI+yN+f+peBhfDbhnXxc9GVd4OWEFZ/gsuXhbP1iJMJX4KvL5M3eLMejXLc
afR8hfuDG9zLVWFa+9ki0psFnjx8ltoz3Q9yIOtXneMgchn6wNVEfwS6l1FT
1nsx+6tvCiSa+udlggTKmvyamt+4M8RcgrXbJJ/s64Ua4kDR/sr2qTAC22oI
+CF3OjQ/saN0PaVlzWNO+vDqXT6sW/HyyE0YDg9eHTRoyT9xATgTw92ySlSM
LzrN6jdDuYjT89BB8XY7kBDYjrYUESXn8DP49AZM6dK3MV3+S3/hQsqXM4//
vlRubY7BVZHmGE+m2SY/22t6MnxvTWqTaVRU1JsNaCmcaVvMeDcI1ssmHwpD
nnEMQQrD2gc8D54GiEYDPvN960fqzxJuDnJ6nZSkcC4sdNxo0pXA1jGmOcct
ruMlAdmJ0UckaqmKpoXHFFH9wmJO0Qc75Pk/JhM4kVF4+YkWvFLcLNuAmoG/
7kg4jMVIthTO555jMxJ64GMLRUJO6eEOA2+6aiCp/R9sT5O0YsczPDy9ax1f
iFa7JghOdlFaKB0seTGXBgejNAQgbIfAilLzO4fmiUzXBzfnfLzFvZ0fPbgm
MoqiPQ8uoxtFFLhWFYOkU4UXdELhYjSCaRFv1j0idLLqb6c7cfRsRLh7grL5
yzVD/Wp1P+fGYU33kP0LZWJxdfMXM+pgdu6DhZ5jDnKP3DiG7LndLpKemgtH
Jlw7He7ADMF520p6OnhDPk2d1ToPogGNrR8B3ZjiSd+48v29ZQxKMTJASa6P
boBqDGWJn/d9/HnHq/2OZrJz2+SUGMN/pbTWMjEhkN+jhR5b04+T87TMFJea
c8PW5Sa+Y3pNohYOviQTQVVIxMyUJi1Y0XOrSkg8cCnxJjlJoa/wXpaCjdh9
DbLbCDDJwBOyc1XlN8Wo6KYjZ180LQgup944OQ8bddjLbaqBUN83PA1KikO8
6RH9YQDWQzcrqmu7rUkMO4jSppYioJ7/+TDknQMTKIDPGzrY40eMNBL2OlWz
MS+gVtqQixYaKwK1yDPoUr0uxpk8HL/dIs+gFRYFLaZIxqWSsQdLH6UEeZx4
3HN0/XcSRfTRRLlXh77/PtpNEFhLhZX7Fj0w4ydviw9gQbxBJiLomCCLS8+6
9hTG0ZeVQkU/b/m3GvXZCzScbbnR3YRtW1429Pp7Wdx2JQpAiCBu83GJ4Yn0
EaofgLfW2bvwOLeNZliEolJSPNesfqjfynoGVIvH0Ag6/NcHK8wxR9H2CbSf
22Oryttkieo8y1pErTAFZW0MY0MPpWMsjv3+WXDUFGuV7duF0+ejqiNZtRUp
KUBZVCxeKBxFbeFi52kCkunUGcpjXGZbAQu/Jsgxd54xBHHQo6+tMu4Wwqvu
L6doDm+sVOpaPZul+cD9nP5Rc6zRmQp2X6qu8eGWoWiPUknFKZHkUcwavb6H
LYswR70JmGmbzMqvwHayt524vnsLvdiDrLSCBzsWJGM3smAvEYYU9I13aHXO
K24VLQiFjIUYHKnSiZKFWhLrJuhnrZS8ZXahUfbN/7DiItaoJzsDzb250S0s
tguaMGC1hTkAqT4gnNdod0ovT1+h5OyefVh/zhC+dsFEvijUlCBqAPqivNYE
I54gyDtthycZ4Ob9GGJbXCWoPc6G3Q0cTp2d0QU1jJCKPpPClIMlXcpqHN3M
M2PmLF5rVgPpl8xUIBXlnsxemY1aOBypPx8IVQqCtOJ7CFeD4sA9lSFEMfok
f4Rd4fsg2JxtRMB1mocsWFmEsY1z9ToTSK5gBuiAV3CeGpORt/rBpAvxTiRv
uvCW8A0z8YOeQdcfzp6XUn953fllCqez7FlW0GPP0CKbfghYRWkTL1Ba7Pci
2jrA0crTcCO04ac7qw4agoo2xl21eW0t8WsE9EZIIQDgD5glNfIsrlBM5bIS
ad0Y0uVnrigJ/PXouYizothbh+2fAn6M9VZseDsJBXD6b8+MGeFNpYMM1+iZ
pDZyKA3lssMgU6q6La84zvQtgkzHXEGjZZ7GRcxBtqjvb83DR8B3uynvlEYV
g2WgQqxXqTiFBcJKIeTBN5P1lmoxR4CUXNVtWDFDg5OPN7uqHaeedWLYDI3C
T+3iapQf60CM9gBVAwjvYP0kzOl9tJnDEZWERtclDpVszoCc7q7m3Llefmux
sMEUV8H+XunRtiQYFMTDumFQKxYZESqqRdXFL57MXCn0pRBZlfr+X6zndc5v
Ix2qQlY8kC4T2vQAKtierkZ+GNE5c9hxldFeABPQk3loleysOGtpyXeXzldR
1BxX/i7QnSSxPnWQb11uF2I/EeAXADC4q4M+QtE6hzdD+57zhtew0x7vfzu+
aBL3PD1V0YaeyuxWYC4ZFbB50k+hkRYocYrgI5k/g0lnVt4n+wxIyV7Vk+3L
/GUPN7ZmpH2AEIT0+CLrXyR3mbDMeAH5OT+v+YOthYru4tpZxibUBSD4kTmS
29jc6EYuwdLMPd6gkqLUnegsyPAsTwf4kEYVusyu08wjj3tNP/trdv74vJUZ
gYNLyg54uxqzv1uIAb1QFlthdrXJ0dbw3ddD3Y6jQpUIEoKgRinrJpVr6c7f
WOj8OeeLUjyMmZNphoVqMvt6za9Vt1RXB7kzMQS7djt46ciXMKbqwiur3Pui
R5BZtHSYxDlxw3+Q+iNUp1C97o1HCj/YfkDK9AYsOTRw6/KMZLr1Us7cSTYy
iTct/G2kGyfWMorPhPOHcLYEGv0RBw8K4ZaQFsGe9oa+b19x67blvr5/jqkO
iNrqrECxcHY5Z+3bYXGSFDz1ZO288Xd1rDQbG4yAuvfereEs7YbUn87jsT6K
hgAFBpL+Ky8UDj4ThwZh820BjIKETl0zyxQWqc2me5DHl8KrDt3N6pQcRpZ9
zQw+lgO5yRnUZL7HCA4YtfErtvdmFP8CcSsP7MrUAIFTilYAkU6guBCtZtD2
PuljNFLElQfi5RSc52TNYpKUEDg5AZok7Lut9FuTSc0EfvsMz1K2dB9uz76A
LwfEg9FhPrlfehY+hzj/4KGkpZIzQPBJgLV9blbvL8X9Y/6GWG1/YZqAnNg9
uY9+IoD2aM49EoRiW9rLnP1AicFQZo62kSoAqzjGHf3UEw035Ot1rrKNEA0x
qx0fh5FAP+r5vQgOYTETiPkd/2tFPIFVXB+BTjrwYRcnflMp2xN7c9IAwchl
Pvj5MT//+3Y5AutgfpXcUQ/181UZ06FKxTCjKlMWPM0KwcSn5TqgfO44gsQ4
vu1yTPVB9mgxjxx8p3sHzY6ahyNe51xk0uZnvfoXBnbv+Hu4l1GMsO1X22R0
bojvwL6ZfILc91juajdXXUq+Qld6mo2ycOAFIcOBLPerEjFyg4x8jZoBWDuZ
Yp/ZQ9accRwy4C7B5FXySwKQWeONf03fAhb73ppw77MnYbAMXYduT/bOxjwU
iYv4mNWO/AryXkNX6PsSXCg9DM137N56I1Y9vaRZe5vq+mSce+948wbnCCLJ
ejYuY9MdYbgWdq95hHHHFpj/J7asfgmMESgXHB4Hmvj7cw6pqgpUcQNvTQNn
ieb5X9SU7ydvTDi0cUWJrMsP4E8Y9jRIDYImlKzbAToOvzdjtAgEOMKFCbgl
fyoXbs7jtDURpqnacGvPYFtTo6JUpm3Qi0thB0J1m6ouhiW94BCg7gn6YZ2g
TvRWChPb6Abnsr3vJePbfwS1doIu3tZZwYfwZJYRHu65gBS7St2Wzt5i+U97
P8x8pyz/dp/HHiXaQYy3059xFzZVBGfw30tyKtIfh62xgHpV6b1St0rPwUku
YRwca0QwJj6nTiQeLRK4s/dmxNbUtLrk39WseSiaLBaanAUH8b2UPSgYXgHG
mr5kukHBNdDbLGnZezOsr3Id23j7iJ4SlXLbRcewLjhoN9epnZ6HLmP8KhoY
TX0d0cakBvlmZdJmHoFLe1d2wLbO42bB0oo7KCQ6TWK3u86u8Q9HyDuvjleY
8umVFymMqaE0VhQUbThK9n7J6iiceT0ORzqiMEUEJRvd5vrkKpGcs4q9+PBJ
nuExo5WYTUZfmFaH0KQQTvRUNKtOcMrXhVE9AQCWjsk/l1Jfy1Q1O4bVr7ps
gSF+GhiuyOrcjM071lfyg2j3gHab28jQ8wDlbJYu5VgpnqLkf+QgwckmlOBI
RPd5YnfWxSPHP8oL1+LcOp5zmrOc0XY3LowZxpXxwelmF0SHgc1xIFa9iSNu
IBAoBqpYFFZBsbgvzA7CaHwtE6lkUE9jXo7g5ApCYBbWqkJgTwZqrk+1ZEaq
SxqtjL+EFsaJggMxxCEk9XUfS/mkN6M+0CqL0KkowU1XkyyqwQStIl1KBqxl
YAapbh8lyQHB02aiuFnX7gxGKghSW18M8nxk6QnltDin5J7/2czJ2kyqqtI8
PvvuXXy0P2zCUtxKP7FaVVX6YxUVOj1NJ1bhhjfKR8PFS8wUlONtlawoLpuM
R9K7sGh/8JfwYw4xKa4kiKJ2jF4EkNraFjZ3P/D2lJVW+8hxJ1IRAqCvC0Mq
ZOCFwHLbx5QyMHlU22Ff3mlPSVQxSlIS2472Ntetux8ZhBntuMPGr1b0w7yt
wgp66FGlIK5tqBTjrTZvm10hmAISPjawClsqX8cgic8DqWZWkZ9zWtBrlMga
j6AMnZBfNi/oJ2X6eTu+1ilFLf1SW5ANTdMRLKStE1T9fEYQpWl1AeZgH93U
pPg4eRKnRfeKDOQ3RHqTr0ujlguot1oj3RWzJqc7EkkK+U16sf7/ZlJlF539
ZTukXKkhukXkRr5673f82Xl5wy9Ja7aLkKdzAh+Q6z25z1Y2D+UvWLYKRfSR
ipt/rHJjeRwvx8UTigRu9S978y93+BVZh76zk2T2LADkChsOEvmspG82ZiZw
Ik/rHIhqKtmvxr/n6FnlV8eqChJA/8tXyBFs2b+Tn1nVoZ6WoeFjctdwKGum
K0FV33jsagUBSne4O95PkHCaR8CE1wrRr6F4inbKUErvyL6mc+sLy3bRYlvW
5I9ecfXaCbdlKjidkltcWvvNdpaCEavNMwt8Sh7mQCCbjRjWisF9UGY6gXVp
dZDZqyKIeQ1bmmHShCuxqXCFhh8IHexhs3NGSNKeV7Ody1TQZ0RqeVyJbnkA
2PYSy4zlZX/uwh7V24JQazydInKRycWHdqemRA20iGx+m4sln5HZprk9SpNq
olwHWKrbjqr3PVEftuWaLQqcQ+3ljUNu1jNZ/41xUJPLWHIYmhBa438CkJlZ
G2G2G5kfZdWaPqvN7I9HJ87oC9MrvNB5bcQh7CCNHrDk36kW8FlKFhOGfn6V
MG4GBwIJKz3QKMmd62HjBXNHWhhHWMDGb9qJDRgPVio6jrMtF1r8RDBe2tiG
FT6fTsUB+AqU5/MFB585w/zIn1rS6FTKw7Sn0W2gLwSrwOzAhCG7egU4Kxpr
wGZk6x/C+g2yfa6s8ve1ZAszG/PuEyoD/FHmsTvPTuDpH1WW12T2J/bvYE1S
UrkjOGH9YEPm9NDm7oqkGFlhmrLAKTbxpsSH5XG+vKyxGNTNAPA5Maq7uFFC
znQV/PBDIV8PwMJI+Y21tvxDjufIdk/QV+D5qyA61iWz7uCSAHPBfVcB0OKi
sbn4aVeAnoFUpDIZRWpxnClsRPkdE3pyCF6coLzD0KTfz7sS2CwayRLb6eZ3
knhoTEDNFGp3j7we1YwVqonuf+762JS3bWQpWMDTGaqhDW46mwxyZJIf+l84
hNDaQTU7VrIQs2rI8TtcEJ4w+iS+19jvo8BRF2GC7voZ4sOJo23vHXtsGnmW
hZecvTzOd+GEeQoNfOul0GM4jbiFW/84b5usO1ICX+edfWMy31XDU8e8YOvX
bYt0fO6RLkQYKgIcp94y2rKUDkYdWyIHbTjxqpq3GEIRIuPd4bdUw9Q8zSgz
DO+vDmr0Qpgn+1fFPLdE6TnfnhiLtnb5CKtkOnnP06k5XGQmhCc7hA5wLNmk
nvA2B9PDHx9kp8Xr9RX0B4lV67ZhQsrTj5MVSij2TfZsNc9gBd2vjYN6d4h1
A82MYBjs6R7SvL47i5F2FK9/Q5OZe4OD5z10XHvnwvkjJVdhMmNbNJCaSds1
QTcOeImHI377JIidyL92ETLNI+5j3MdTJVoK5KQ56e6npuN8tJ8ggoS8tUhu
oBME+lZgM5g/FsdZWvSUKlPEDANLAj2eC0CHkT4L/m2puq+pr5Gb6/o6mE4L
DnTyor1JA2xrb+XkMYKl2FNjT6HOJHv0q8Wbou4f9+TSZIv4rqc8AlcYIbKQ
vKc7dyTsfCqWV+5+/7Et1ZzQLToLYqRbigs+2fx+FcVtpoCwGux+IkvlFk86
ICaPRdGcQZouieCfVvtPjk+IqiapiTHk67TiUVMhuvm9+sWGd+arjtSgpqg5
SxYbg9FH/XdZP7cgtD2xgeHacQWv8ADbCIP4b75gMxWdBD2wCvcb7M+ykJix
S3qySSBqLL/DZgt/hy84beAo2dhDHFtNCgvwJ1yrFUbOl8Y3hu7VKbs9QUXZ
yL/2Kzgzm3/ooDYP27bXSEvWHcmBUrqjLqCKBMscqpWKjz7Mv81/FwK9KovW
ccadjhOzzQivIImtscowmAqg6fKz+F3iWlXZICCtR6yiOVgJJd4ZhfpvWuQl
XnJJcAoQKtMDIGfQnD7INaajRS2gxq2ihHNC0Vr3i/vhnMDoYkjqk8TdQCxz
J/2Y4ybD2dbqeEWxDJnqqGSBZYROBIFvmfoB3UKaFDotHlG+zAgVSE7hIl1f
3uYjF9W+aH55+s0uhVkKsSebtjAyEyQ8kXN6sku6dOQTMnZTKqDGp0krByPj
zRLYq+FpfZngnoE0pdy65baaHw0rl1v3uDT3TjvT+7FobIQ7yROIVARQeNIx
WLSQbMewzruyFSU5vEpON0FmbnENp214DGiZ+s53hWPJYF5bMg60+QlsPB30
FggSpkQjdkW57gLIyRqQ3xO8V4nvUd6T0zbN2eGu6AlthW9HliNQPrrO7gIP
akYf8Gck6vbJKk84x0ubilUKwXS19Zb/oGVDs67rKskEOhzFl3QPURUmTNk4
kieXp9Uz/SUxj2hb98C90PIFosCVLGAbyctq93/N1RKdgpWPoJwqcduVpfCg
ZTq156EpVgBpsYGCIvUMLIUk2nd+xX1+u1ZpF13KwgiGtRrIWAY5ZBEh5609
XiR0WN5f+OOvlSA/Cfegk4apP63n7034g4wDwTqnuPCPqt54WzUR0BvZ1WSA
/4uTMjHlYV/imxqmIusUWLY+j+EcxILeBixWt5Xe5aKF1UnYMkwkC1ClTz1x
jCCm/V7c/ztSGWK0XSnx0UCF8nkkr//fiCTz/zz2O6djsvr5M8+EF5d7jXzr
F0C3TKKHfP43mA4jwAWPm3I6AxHw2yoJXApxAQLu9Eo9LU5Qu92ibS9n/7J3
YHjnyEknl6/D0A3sU1PG3ysRQi8lV6c/Wr1TTacfT/gwtQ7gdg/ateATzdar
gAdT5rTcZD9B0kE5fH+DjGVfUFQiRJd4z5UFxcXSGOkIgtYOOHceAJj8/BaM
JkpROt/rOUMF0F8QavPV94UEZb6HN+3cEuSwfq6fw7YEHuKmRaWLaoUq75V1
EHTHfEtf64/XGhtCDuBK2Z2+Id8LFAT9EZ61Ky+fBA++VbIa/Pczj6+pCj1x
2n9MIxGmQjJ+YCcVBL8wayWlAlq/li77SF9MzUmJ3SHbSxE6ouEVknvmWuQQ
UIHx8VnIzKyiAPtQwNQVkFTy026kSTa9vgblbUwsmM+s1gDPuk1Lrag/30dQ
cj95a99QCs73TLArvMYOLWa39MrUbFh8K2w7GV8Et/kZm7Jmw3Kv6N83VxqP
03xkCnTA/nETroxMlpqGqVg0znouujO4lRmn7UH3que03ZsEXAKrb9f//Zqy
EvCQheB7qBTZwjIemomtvy57S68JkktAOHwsr4T6/V3DjmA7EvIzcAfxlm02
VWhFv3480CtjDKndxKshB4JVtZ2uRh+XlxIOquE5glpMAnptXONpUclx6EqD
geM5ytIEJqnz1JKG25wXoItnXIid7JfenOKK4ncaNONtx3SFLkTYZRWLBgpr
1r5UkXUX1cZGkZJDM6Mo9gQNkxtk1NQmSoP7ahaQPpeEpfslalKDI1qI6RY0
NIIJ3fDK8869zlYDfR5lTjx62vBD8h2k43LYNq8lCJZYGqMjwhU19E14ewNp
yhYOfGYndydSjVc+/CWNeome4OvSpw706ibxgm6E2wujQapM1D+67YFLyuO/
Wvui39JdJwPCXNKg5ZrwJcU5exJlagB5HALEAXcdhUsInXups6ynnA3L4DAV
uHkpK2U1IHlgSigtgrjc2ttEDxALX93eVdS/MFYCd6lkPCvgSqEuqdlqgTPq
/64SUdm8Li6D5g9WfvCPQhkHnGkCkT1Nv+WNDq6aq55pjNU2F7Rnj5FQ3bLm
gGeeWf2cm9g+AGHPuNHUhxk2E96uNWhniHZP3cSA9a1gIuOxnm9cNntfOAC2
wd92F8h3zAhrADRPLRpWiiei1s/z30fyRD7fmYigmYzWJNJ9BshgeyL8hUmK
wtlmkOX9ve4amUItu0nP+Ld2xF1IbNyP6uxup+SKTGfOvzWveAD1d8P8lIYy
6B7vHekKiBPI3GipbqkRFKdsRlT5sLz993BXW0UAaBW9xkd22fpWugAXlc8+
jALe1yGnZ+fxP/w/szeh9C4Pvf34RTXZlIhE1xXx8SXmeJI7j+MSRUgU19Jg
QMfy5AWvPNi3Qo+lsyuqedefQSRKOhHzHyY2DPfWc3JJMWQCXjUU6Hhzp8Ja
DTm2eGRhcfsMvs6/wxUW2jVDZxfrUXv89zESe4P3qNJCxYyEH9ngrK0Yg+dm
zrtjWiEIngiCHe4/6Gy6GRzfLWdtYpT1K03G6gLRFSkKOZeTElFzPZ7Lkryr
01Iw6sYzBq/pt7khH8tnESEGhkgdcBB3uUxUo+D64YndaaUOKBtm4IIF5zk3
Q/j/zyOwLCpz9EijuZ1w6aoSj9Zhkcci9LrKdtN/XrK4TiSDrvba3xk0Yl7q
1I24T3o7oK9ZIAfecx9hEn/w9RD7BJTZE8DyX8LZBu9RArGa1S9mBfmr3I8P
BPEQmw7tP4q7WbH+/aBsIX0Wm0BHxfzEEFBBnvU/MCsb21J93ZKZ67wlmri9
ixk7WbFOQECLkghdULJ2qG5PG1FJUGGcKHqHZ1cciwKZzVmfikXgAEGMTc6M
sOcspMmkNq/CNHfSHzd/7Bu2teMeeOeXfL9u6buWkdsuC+sZwP6bH7i87Kb6
dJjlQtm0VAZQLMzDvuvt0sxxgzYHoccC584UaQtZoaRY+akN1LipYxo5WpBu
UF2kkyWmOmOY3kA4Kiw2odcZFpI1Z9aMH6D9BO4ElL/hTz6ZT06McPo+XVbE
CUb+yr18D0Eex1qN2dmSDI+HWcbBRNtxuMmfTFMHVLHIfeXhhdEC495u77AG
Owkox3VOFvhK8CAvycDlWJqrwZTC2DBlOw8SY/Fm9pJ/3XJfGiS7L0Yw2zgb
yVd57bDZkyFMJQLIrR1m4O1AfOuH33AeYAhqC9RNtOo1GZJQU2uHExfXXzKg
W9lQu+Tm6pHf586SonpSv49/ZIcO+1P8tYgq+85ZirXxBIQE/tC0gzBq5PIT
j5z5JpYrFLlslmg+twCsrBwebuDY1YUKV2vDh7m77z8wI8YtkhX9FQzixA9M
j7OTIdDE/CyybsxqrcGlWOwBv86pN91VmMYO6LxtVjLuaM5afyhZckcVoDUK
MzZBII32J7FoXkuiBmqnZhI7BTk6QqoXo+ahVqsZ8qyYrdRYK9w2qj97tX+s
qmW71aZszGPAt7ScdVFGTqpLHuLmHEsISnOZWzQt00WKr8obI9xHC3yKApSE
8ZZEQf9nQSUdFkov93QcMmh8EziQH4L7xe0EVjDbl/vgFuk9HQU8+B+iHCrB
97oqhptblrlvSSyhFrEiqH/upVDgnpuc3gYHF8UNCAAa+N/4EgBrbDmUcOp6
NLS/k/Mb0WPcvjQUgkSgw8iTVAYzoh4YF5/kdYES/OEKbO0AD5VtuVYXt8xj
Vzn2AbJJ1mxS+bYTjD6eg5mRaJq5fENS9671HaRcsK7VPenY0U2yLJoEDGib
88LA33qeVtlecEr9RRPvU8RmUqeXv9l6fWMxQmIgZ2/z3ePIWAJRhgblGEPK
5VXwXBH5PG/crA/8g8pOU1DwfZ7wl0fXVWfrHvfafiEm2RP8fXF+Whcvv3Tc
mXxqLpI2AVMD+GLrsYriTEOTyXsBtWW9mksYMpHNpaM9Xre6/kLIXCz9O57C
J9yGfV0zhSlpff8lX2ZwhrG/Rraqtxkfxd7leA/WJMqFj988FL9ymeEZpLfF
uM8WEDEsGQrJMljRzrolYNy4Dh42hN0muPtUC/6gHPbD99evlq7rWXvc0MLT
FdpXNbSFVyPMKhtitORqtCrRI+A20FcvDfF4RrgB49Kn3CpsKuBtL9Sh2QUF
hj2N0d58f5VW5PxT3wCIuXM9Q7S/pFDUJ9OzLhG3pTDgmkGxAs31sX7b+Ka3
zU/zJV8ychhtYNjXbUekbaeCF+4oDoi6Xoxroqk/f1EY2Z2FxrNbmTLh5bVg
uAJKVg3psztWTSLcCKdxu+XDsQ7zCNdBh56pLJs8UR2MZd/1RvNynnWnPC11
ffHGQIixr4AIIRKgUA5WY5QyQI7wWRzlhXk5xeAfSApDLaQxiucRcVOwpjRw
oAa1NT/65Kxs/quqzHaa5BVKDBo85//ykEpzFs9DasemmPs1bXhZxVZEATmO
nzUtUuFAzL0ZvaII6rbmmsv0zIf2ShbmyfsSftZidw592jW+47CluKCmhgvm
mCwVMvEgRTJasF7zcfVQtN8YjopELscQpeat5DrypGTf8FS50IKBGBxE+JiR
Q8VTX6lbNEbe8TecQGRQihcWYezCzM5wuRp+Flt7YO61qvwU53g8BeskuNMY
eQu2iCL8iFu/9CqtgDrv8DbxyMwerCz8S6oXsvZiPDUjTFsncX++HK/wxNsX
cI3unBELy67cZ8H4ygYYjAzYNuOMezPTRtBGI9gOzcZHSLft105mvMYH7bBE
MEYqCgwY8iuy/RzGdRavl3iKm2gv0d1eQv1/dUqhHyJlGqNIVZdRhCiix5XD
dDKWpPgySGcbV8vXkYnUcPnXReC1wgmALEIL6ImxB6dcjgUtMXCBTIouepn6
hfz8ckxWRvS1EHTMHCy2B8uF9RTsha3xNSzCdtoB6BzcE8OkKJGpwh36IsaR
NQEBACzs+dVXFPROnX7DmNSDJX1nGcRD/izGqJ0p+OEmkFKOVcoZhXbCx25S
Ns5SWr/oihEMaBf+xHUD3ke1UbQq8V2iEk1u/GKvSmgTa/rA4cIDD4ZG2Xoe
LGTupmfkwKSummOYdYpsfjtPgeyYvXOLyYKbHdtTqxOlOwYhI6RNfYjw/DbW
mPkpegcNb9nEiHIXr6Z5J/bSR9oNgx+zxGPMEk0gV9r5rPXudxlpxsp+NmFh
JgPAUQsqbjRw55wMdJnRHM4vEKuiAyfJhlUCP9oX1QgOq+q8Jtji8rls0TOe
khFCA7RHrZn0g858UwwX8ZDFAn9/b0bpdLGXWiamuRlH3xvMmoir0Fdcxa7U
HzI4La9rQI8LyXsHWVQUdjk8tLYa7RZBukTnZXt/pLUy5U1qGTWWLWacAUim
OzTyIxwuqXomgpSwTxofeK5bVs98xxZYCPvXtU99FuvtUT5ANA/8ovN4oBTx
ngTmOdl5iP+D0etUvXpxn8VbOT7nDy7QXBC7xlRriSmHDwizjfD27+ZBMa7g
bCG2VN95ovt0hJ7Xt+LESR10/7U0tGJPAtGh9WRahAh+HMtoab2w1uBA5b7G
TakGzBZzB+Sa6gN6z/UNKmZ7+TrfPF40X3vyMgcXr3isuhU7DwtrhZGkAxU+
6E3lpgnhAyUs+vkYy/DwAiHkuFhsOemhv8HbYHE5rJsK+3eqOLRU8bhVSwR7
TrVdxc+VD8TD/7Xy3W4AlA+RPX8oN6BIdNvfDPhNpxmMDZXQdZOvT+wK7GBo
IJCdtCNJ4aRFVmMTurvZ6Q4w9emtByi/3trpXnr53l+zrTJyTe4OmQBSoBVh
cDmNsObJ93aQELy7ypfLFUySVJrC8L6LLRxfOk48f1YPD8XxD3xrs65mYmT/
mMmc3RcT+AeNkT7BDbFka444PzNGdYzje3xm9CQVoHVMGvjHJec7MLbMMh2f
eECcIC+WCPZdiHepF/67/bJQDO9x04x1KTUA1o52PdOSBldJm++d7aFzVcHB
mEqJRRPHoIeLnlhYu0eRjDava5crvs28NTDl64y9K2UcZy61TVG2sI197FTQ
wTTQr/TDENlcWVGjQU65lSOwO5eNyBWV/D4Y4udBOq5NvvBrzIYmnQyPWHIH
1HD4fkJiVUBYt+JLVJp5J1qMEOiWD10gXJw73gT0kPo751L3ahiXfZd7GNH7
K1nqn918UxEgelWMA1RRAYPxBcfmZTuLRSACf8cJx7nvF0q1AXiusx58yPfp
2DoyrsW1nl9sf0A4eq7B2xXrM5rvmNBTwwBf0pQfCo2GuwXJwbPxeV8f13fc
mGqmICHvV1G4C7qCF5xmOHqrFUd6kOm8Tx6Mwe9ZUtEg/m/fYBaiMvb3wbu5
wlaL2ZzwMIIlVUbpOLrahmQ7Fy3RpwbH3DYxHc9eWp52ezHunB3u6YYMITNa
JPvF+FMIU37GtDR4yxyca4fFIbt9U9bfzAYsjrhCy4N3Mz0gH5kYPHwkJxWW
9zDrwo2TVGMVjvNvTwospkfGFDdnPWb3YKmLRsuC6//F+5WhOqVA8yqH8ZtK
st4WPf/YsOzSMAIhmJYH7LIrkCI1e55IstkLFol9qbibuE4PfVNNair112wZ
XQ9bzfd9bmkLSXrdqcOe+CW8+OnIApxA78ppGO72mbkZw95GXQB/dXDwfPwM
mJuH9ET/ePQvMWIWu2l+289VVb5/+fp/Tmsb97JXjAKrTt3G+ezZJEoWncEz
qOE98OE7l/Ia2zmCtKzveA1aP0vhIzXEB+pgfCD2e+t0jQQvKH9FuTnYOoSp
Cx+SI4F/lm+ouneDmFqwPDgWzEJc+TynUk+c/nGbEd1zaT/HFTuTH9jb6vzJ
YGH8bvWEWcqZNMf7Sxou4Mnq/0JpSY8NGi3saYs5+EVdGfXocDpXwib50HFZ
xNgv7502VrIRB0iw4Z5w9ZPS6MXqkZCrqNGLtytoIQpUOsAD8K91RukiHXrh
oCZZQz6GWV7ROP8KkFKBUaTbFGjU9ZsONcZfzFmSA7+0Y0MLLL7SKgCWEsT+
SrSkFKAV7iPrpGhsgqQue6AckIg/L/tf8B2BlhV6a7LZ3rZY3dGF+0qckrOc
+iXxrwT31YNwfBWi/CCYAXH4sJk17PoUrJIAo6Mp7aQJpg3Aciv2mqG3CbLQ
BODwK4X506xjXUFdKyZdmUefmdluasBOQVtR7Uu4fgPi9M02m1DhfIcXKkLP
K6vKOaCO8qPAujhBpqDPkdJ221OpoDnfkSxFZdvRJ6Hx24pH5XwfGkgxHL1p
dFUsMgENj9N0t6eKy4gtVNI7CQT1O/qVjnUzqvYkk12cvms5IHkdInXYaRPt
25n4808HFbvt5s2O+RaTtqcDRBjGc0bXLB7kX83To3ghMqst7E+jq3cpxmUx
5WoGChYFu6YXqXospNU6qlc2tOj4/Osig5C5ZW1hgoEMtPt8e6cqearYUE9r
baAkj2egMKzBjFG8X8/voPr3T+Ieon1J0PzzfVSqK7OolYmvYhGH3UVVfiYR
UZvRoOqh7vAhg618XbHjEhMWnvYyuVeDa7l6Wb0vMDQzP6EpPLkqiUD4ybex
onr3MTu/pFoib52J+qlFA8N6YQMTISnBw+tdwQdmabWvE2E1UUUgdfvIg8vS
QLdPo6kC56xcBnpdBqrXhD6J/Q/SlpPfDWyE21KsIXfMmEbne+8HtWLWljRg
cvSYSK2QlOr9diquf5RrYVFoViRpY1swcgzHkwcxto3e1wqcvKue8jj3VJYN
WXti6UtZdXU0TfjtpEXqRwhrjzYIsmazaY6OLVTk45efKY0jSlZQR+qo3QLM
5FOl8F1m/rAiFKcx29Gtjk549opFvcK2//4yyH+9bAE3K3spoGjRvhjGOXij
mGcydgvFUst9UAFkYlmNw9m02ZUUj04Ko3hbj911Y6UVXcm+Y+04OC5VO0DJ
TngGPrx1Tg8No+z5NTnZp88xwnOlelTW5Cz+jfOiICzdIK9ErlhT5Yh2PMSe
4R714+oP0I/j3c/cQ2JOo8vVuQEZdnKbqkXWW7qBOpn5DzCWlOZCXl7v1cx0
ztLenwo1k0CZ0uZHsXvWisMRxJZ4x5oyHBPTPfztt5sX3a0XERvf64RxEcRt
Bbrlk3rPRX4Cntrz4PS9p5CxFK6kLDxmaDOJsqxMU4ZwcrKRftN7k+rsWx2i
nI+7jrxX5OWVdJmMXqEFIfMy2SlnBdWxWWtrGkM+qe4hmMTDux2LAfqcmujE
YpG4/HBJe6MRA40qIJVqU6kIcqHRo9pdevH0HX+rdYYzMeG9FmTSBu5JqERx
W+vb6FjGMYtdlyArfz21uQel2yP3bRcfh/aqVxxAWJbNAjQdNbi8pUV2w47Z
eeW1x9IXXIuyDxDhlCWphtWX4X8o3nTwYI7z7oKZjwOICeoijp4+jLWXuzZR
InjoP6pPNFCgUvA1bmulQTYVAubYPpcwq/uDOlcbd57gAFHSwZlBR5SnXr7N
jCKKIzvwmTc9Hh22B/hYQjSaZsSwATfFIVwD07p6sXRU7bX+n3XMfHfB15Aj
a2g0XNHFfaTALEm1+g8z/S9tEHwsA4CMzgo/sRtGY1bBWu5RAF0atBwRj1xC
cucPL5gkPOwr/JakfdeIDuPRANL/dZ9oqJR/EjxRqyc0gjHPqbOvwr5oxqdz
Fxv9x82I0theV2v67HAjiaQdJVs4DAFTHSdda1eOrrIvGJaefiovP3zzK0ok
LI8l9EbZuAe+7Z4rX1I0zXW64VBii90SdqCqMBdO0GvxT9FEYCLDiVpdw/fz
oIYge//39rqVFoRD7743vTVY/bWPf0HHwVHZIHTvkmWLBgEyaPI/K3+/C3Dt
mVTFVbxoi+nhSGoTtHj5FRIHisntUnmSG0zfTC3ZJpNj+fxdowhGh5sW/Hk8
oQixGeIF2JaalALbaEYfJqc/iBOtEbq9YAPjqrAaq1KWGsre4KxDUP/fXwXx
iLLxuONuLp4jjgnTLalaC4EHeQTqizvHyMadXH29qjWxvySj7hLpjSlsvLL3
GI3+jNmLC3i9tM2yNAjFohBrjVMYH+nQqdYqntDz4rnD8upfdHfXVuYiALu9
fBkpSHLKPBTLC/s2R1Pa+U9RcizWS8ZArM2Jr/aZ17F5QsgCGz8oDyiA4XFS
mXV3aDo09yXAScGNDmtoPD4LAkJDgfVFONDI5AsTj/qJU304OR35GkEfDb9G
c8V5wokuhDDA1fB57s17FL76HlRFwGKsxxD74cwlRZELURgr5YP2mnzbV3Md
n04cghGbxBmE55U2Ck/V1f68clGjQp+F05r88J01RVGpWL2efv4GRpJJz/Is
0XAjdyb1ozQNNfSWqFNv8zn0nvaKtpTvnjwC20X4wg/gC1jWdNE6aIYTc+ZL
58WJk78oHSYGD8TaWEbSmsA03OhlbE6SqYILlV6OxqCLEoD0bhlbSac8qzU0
GV9qldOPQvMHTr6HNlqHVpzD2wTopptn23E+piWxxXgmQwGfT42cj9aoV44C
+xTMjG7zYqFEoOza3jpqYHhvJ/MrtmgdqGApyN3ywuvVjYsN4+NudPi+U7uN
kjS2vmI4aWz5Iz/K+sdaSe896JC7OuyUKnOeQ69/JTvNKFTLaOmboi4gA25E
vUv7xJ2NIa3aalGT07dJbgY2GToLyYdVsX4Cw51IqHBlQP5RCEjjSFPiJwh+
wEAN+Iz9gqXzGg6Guf0LRF9VsqXwjp6JYQlOEm0Q7Znf97oy5xkZzzAD9zV6
H/KpGNRv+ybnOAFBBKMwLfp73IKV77g4zWPmnyFHFGFXlGMEJ3zbaoxAcA1W
WcSMjfeYNYQSurpmjaK1tZeYk5tmIBjaaWIy05bTK07aTnnIogTZwp+GrxXi
IdTUtv3616CzXP6aYXtLaeBPiv3k3bDrfwNNZ7avz0PMMej8NttOibUU+QZZ
/cmvd4eEbDMZamELpVU2OzHGSIxW5xVlpgzKtKAjU9K3GimXEDq23QP/2fi4
w+sx/lQyT3JIAzV5r0aFcbTxzL2TvdioaVPz0nnua1kAwbikavb72CCujK5O
3gogs0qvHvOgat3wskwA4g3rbuQ3Z+3vDSxtTDes1wOGrLcILreHZR28NOMD
UweEG09i+XsXfAJFU67u7vVn3YcPP44FtNv8RKJobdoXFpvWFmhAr/ZDTinf
VXFf5hnIajdyS8dz24ecg2hSVUR4Bd1+ayZyiVvdhRA63SP6JW862HfhPW+f
dDGF76kZB14ypKITVb9nLyHa+w2zmu1Y1gPpgNod6/Az0bXml1T+1es7gE01
ksnfdf3sKnBahWEmL033Qz81ZQBWPL8utXP+OLZPmGZWPmfzAtoOAH8ga3HK
ND1K2l4iDEfVQcdGxBAlhO0HbjhB8Nn3x3F5cwzHa9CZjedLatFrE8BMfWI1
grXqREAzpX+8TpyEdcxL5mBYzAehnfm7iT8zROd/0AYWEPWfDB8xwv/vDI7Q
oO6TaZFm4NJ4cHn4PNtIztLKgjiSYRp+QOQ66KygJUwcHxUoaJwWRLQ4t/xo
Necjvtw01aR+xPS9fZJoaddj6Sisp9Rk1zcvS+7LGu7zdU/0nlSTQeSo6deB
c9D8AXV69t5Z42j0j5pM4yxjOYMohsKasTYFLKOTdPabUDvZHsT6fUl+eLKk
M0MZ8vITmMlwEvzPqKDbc/LKvZre55tYbGsORssqg7jsOiL2z3rQGClTkbaK
D1GBB+VQkwTNTFDXq0cUmGEYoA8fQb2xxdTm8imqR8s/UbQZ01K+s5rfwDNL
NBxt6TQiiEyzduhOR8Nj6TLzmeMFp5iI8rgef5eHFYCNyoliY9YqqdGdl+tO
Sw6SPiCGbu+E6+ITWq5LEbI9x0vmshcTQYQTFRiPL1DT/BqkS7nRYac3/u9G
GHM5dCtHbnHL/jrB+mnNV52n6jova9RwLWzCEVVdNnjJx5rzwZWy+PEzlWOG
3SUcE0BO4wpJrDyX1XtXdqF34t8spoQORzFyKB2oGUvv+01Q1Z3Zj6ULWP1X
0MSOjHSvVySiV/452gMaY3oUGCRybKC0MZaFTa8GuIC4k2R1OGOwV3BJDaMx
7BxpQ0BWwcUiCPPZ6JIgm0KOOGyraJuUzxPBFB7ujMIUTqvp2lm58jThd8xL
3VnkrCCL8pUjgJKDWDGPrZC5ka04c3iI8ZtKZwH4v7ol2GL3Fpyx/5yZIVyc
7604W6BeKomhHuzCkBsVlv/nV+2S3NWmuFIo+xtREAQfnVcFXHPlWSxbPcpp
Dpb0dwPF7KY96x5c69+lzYF6W24K2i/vY/22q8iRqjziEwJSt3dxmriXSR0w
1MZhUo5iIZ+Xdkiqnf3xCOYBfraxXFzZFuqNsQegnPiJT3Qh0GOLXjuScQIm
+wJJTatdWPgfDwQReaOpZR4nA7LPTxt+58bGcPLdTt09O4L7JAUxj+UyIRtX
Bch4OkAd0+pKPhR1kJEO8n5ZAtEtBgXODFkdxTyb2+xOV0Ipy4quLxEZ4/xb
6nhsFVBKNci/wwAJw6oxXohy2oXxuAg1Pi7DfaqM3W2WvuTyj8Ogs1SDLXOz
yFw5O21AKwziL6sBs7yz6Op80u19sCHcTq+3odrx+4PIon4c3HU6t5WgyHYR
sPtpgyso8rMRC7sa1vhYDG5PaUvLBGCX/Tf+0CbuBeo86dTPgjAPhM10v7ir
AfkaXst45Y2d0tOD3L1s7G5UnK9KOL1z4gpZ0QgeOev9qEfVJ0/OhtpNZdup
yK7MdslT9T7uvvkesOjS6EKP+Xwf7KfGpnefNgEI/JXk4SCmASncywDo7xVC
BkALiJfnQb91KCOLvQcvUiuRjLZUsWaAvxz0Vw9oJJkWWLiIc497q4LpoIQh
cyxrzAhv0brnr4jlqQzk/2l5xoamSO9OTooDk8voFzipQM+X8gP7VPRWEwiC
stXGWx0A4Ki6AANNrbDr7yYATvel7AoEQvxFaTgxtein3/2u6rKGGJoj6oPY
JMA39PjmK4xvGFckmx+xW74OghUEx6yAZwkTFBn3AVLxG69Rqoy51QsfzejU
SBr7VYjpLLwTQV96s9OclrUWzBbK0+zixOlAinScZnNzf6EhcpNfgm66newu
IYSYavPYjo6RBSAu8m9CwuVW2FYoI5ALJAlNNzQXueBEzq48BVpEcM8J7gRD
AQweaVNfkE8rSG13rB4XffVHy9q+aueBMTlc5vDglIG+grQwe1tyIEHEkk1Q
QapMRk/htNUuSHt94U0k+eGif3HAAl8Md71mgl5aKG1z7u+ZpPkGp3mTDAMP
gU861aBdrvySuAql75Vo8y0R8vW0NaziH8NEQxMuV43b6mCO20Pe0nsi1fRD
JJWxpOOakVvng6OCykqL4hx+ig0JXUbW/n4zQ4Uz5yZ4lIL7Eh16xGoHL65u
prv4b5lgvCagBnR4yR8L9+25APHbIk6pGCkgbb9wJ/Nhrd7w15XTPOr588Ip
hpG9ZTMG/+eFvXA5CEm6txykle+BqF7PiVUwOBQpO5xz4WVo0xf4eQDt0YWH
hhBwW2zMHleEfk4oXKIH9RY51N+o3+YHrxEzGxOg3S2fsHe9YB5Fb5JD+jd3
grFn8CPN0af1KyS+wEnWSBuKrp3gTd1/++cEToYrfFMIqcgQdoecB5h1oBML
ip205n0JeXkkAxo4PS/9Ql9DTyUPDLfKOpbk5iCXLy/nmdfvZM2kRWGCaOJO
OtB98on+y5w2ZtrLjqslnT8/RpDI+CL7z5SHqPql0qiS252D7yda907SIBD0
X+CobfxKUhnbaXj8yNj+9T7OHwU8KIpxeeQEezU4dnLWpMR3IiSIneNSnMOO
dJbtlqLzEYPsxQwp6CH9sa81RICN+K6wcoHfxE3/7NTxLrmn5MxlctZX9Gpj
Ey1KMUuvCDU1oVN5q5ntqx/+j986Ow17tR6VSUrYhgpNav8NxC1zfvoqlbIu
j/AV7QUdKyDILIifG6lOLisUumsl3+MaoNqosWeiunDyd1BAwa3tg+aso9wg
bXayoVOS9ShScUYHV2VHhze6wl+THe5UNdG1/iT6qfGRxbqjQj/DlWwoR5xF
eR/9Y8sOWLm56wExul9UY+U4Y6rnRzXfnNTNztbONhMsIo0Fywy+yAylipEc
1xuAoP7M7OgmyEYQy8GpDUamjf8Ms72wPbIj9xwbg6yBydU6HPNLjD/hcoGK
BvzzDu6/sFxOdMVvXpfanAtHE8lKVr2gW2mRHDZIQZW55OSYNpzLnj4vHFM+
nRCfuGpZ6K3GmePMaxHWwk8dOm3GIaOPwqRs7EHyz5MdPZrPwS4c/a5CwGJ3
WnA5pwNwKHp9uMM1nhxgCbIuU4ZhToxI2WPmX5QXaTU03TUyGuq/pIyoCGmU
CDN9Q/FoAF7N32tDYLRqHxiEL4Ce8mdpEjhgG+EmyxGuL2+KZhbA/hGCZ7WI
8HDDa6sUT8pmfk6PMJ2W2voRkfK742C2x+5MSYCdUG1hzmsO6execXJsVgiq
9mUCtsDudftLjFt/hM/1M5Dla35mNHC4RbiYDWQ/KUioj6arke+hi91HfPTn
nma39epEYEsdz0SFCiZ21SJ2O9Ci9geKwlh275jggGcLP2UiE/qSQhppApdV
Yo5g21fLH+SwP+j1RjD+CJuD/dgXMgQk/J4qQ1232X5Rcsiy+ocue7Ocvgf9
Rl6k9eoXp1WfpabCLIll3cnO0Odwgmah5Um9NROeojWbo2+MX5xCHXqZOtN8
LG5YnJv8cfiJBmvnE795RWIA8YJ/cLapekrx1J0gIWpPue5IgWyR9LiiMS+P
9do6St5cBmmICppAl+/sEflDs0ICxf/map1WzaDZ3DYAjoX+oeSPdWj0smwf
9B01AJAOr6cZMDaB4V/Fjww/4Hh+rx35rSKjwdRGS7R4G/Y7fsnm/rOPtIgf
mbNGx8amEEL62Y+OBbnAJw5WID3uAZXeHvDOlnbqzjCt1r0cVZ6d4yzuiRlX
jfFC9oajM3NxfqGYjli+xaWhkKaTcqFeOX//ndcQc4+MAe+chkcRczWo7Zb+
e5uwAbuvsxBtFMt6GDPWZANyCagRzD3hK75m/vffXb6/rGtbkEiNFf4eAu5g
2UvA/hz5fcjUsqPZTQCo+DNKTkDdw0nKGUU1V5GeAxhs/YGIWpHlOfAsH6/5
13H0NjUtt62e+UM0X+/K2F5k32+xpZlaOu3Un7gRkuua+I+vDObqJxafMDoY
BZNfD5phm3h3k7VKZotPa9FyDAzSYC29nlRoWkkPo2/XjlH1H6QZAc8xYrjU
PyPdWC3eDAlqpOZt57we+RCd8dUUkWxJ4NvlTH1i5kDkLb3wk8iPc2tHB+Ng
bN5aarIyPiL/mxBnVc2tA9CXzhsr9uqK/11vNMkClynoWcar7mPeIIgkKdPG
nzoqVOrw0Z2Mv3+fqKVkUiB9tWzbjB0mH1lEWY2g8dRT0ehtBZ8fMzdEctIB
S46Ybiw9vWvmAdpHEARvuhJmy3yFNzgEjSFD8Pgo2VTOE84nres4rZ5+1+nz
peSNPfhiYp956y7bMaIr9Y3RAvVl9pFYViLPQFpXVbYw82iFAfydTX+I3jEV
gOG8geQxZveWP4nqr2eJckuQxS1NYRnGeeKsc2AiSLfqWUnc0SgK+oXiLzf8
vLDHCIYM+9Y5fPo3/si1WssALXXbbEjguNS1V2ktZc07N5uzmYBaHMaw2I+K
HjQUDQVmpXF64d0nQby7PUQzBeg4jNs+8XKTgthL6nk63Rct6vt8osV5Q9GS
MdSuMxSZeYDAL+EV6YPK26JLajgU1mrTKoxvyiWFS3H+HujfWYf72mvS+1Kr
G6H+PWYmF+H5NoFkDtA6kb31xGDhCbQmwmovOGbR7c0u9hYOxADBzP4mWkAq
UnXo/+MGIvwZshIscJazQMtzd8l/JtXCr7MIOvni8YsPG/Y62lFIq248kSJa
nM7Y3tFm1a2rjLgZ7RPw4M0+3V6Z/szb+3Y+emD4fyaXlTZVdX1D7UzbgpMh
JPfPV+AM5a5ipPpqRb++KpsrBlCdfLib4UU+xJXvzSWZQ8lYnTTK1194ebZR
j2zds1u1tphWizuFa9uZzS/hEwg6ymnd6fXDp+6JYLzUwSbEloF5hkoQoSqU
b5MoOfWja6svIm8ZFeqri5TxSpVaaPqRSp9N0f1w8/RuqAFf+zOA6pOPllLN
FVVmj21Z8XpvIaUho2v1TJPB3Rz0cFpGK/EaIqzgRfKtFQbYWRq86ObFvDF9
EvyvAHN4GhH95iHc7wvV+fwCnT/ZBN9XJ0CbsI20nNYUN2laffjP16WrKuUt
MCwWRWdLYvTcbJDeLbpPKVaiasklZAWcpcy3lCsCVZL9u+KMH6Ke6Ggji2dM
pnSpj2vi4lbWFV5vRJvVn+L1UFpOyMV6pJElPbUoDR9d/Czis0SnPNJ2Zs9n
ssotMsERVBnJtXv8Bx0DmtIrzLIpm4wIF1JrxE/YExQe9s4t3VoZ3J5NqAak
Igu+IEOEqtUjzfHplDVDqjUo4rs7A+I7EpJoUzJEvDhRioD9uOeLgAoY/KHP
sSQifI5wGQu6a6diToYFCfe7jUphYtEDmo9HCIFJ3LpU8aAriTU4hZOvAXkS
DLHzU7yf/CyCSirzbWRO9F4Wr/cn6nW+cgEF+AcmrakF440BjpZcP+JXls5a
LIXmDigiresDhlHh+gKlROcfu8SREOqRnlBZHp8lQ1P/Bfxgwfh1buh5CjXZ
tW/gfssQx1apTk58pQ4H93qn8Ib65Y4qHtfNdIV0l9rGrzrfG+Ifz1rzAJL4
9OhOMgZE+tzh6J0maMiOjPWuHsFgG/TTQEg2GSvi05bfdXSncRdR9i43yAZB
jyUOkHDaxQDHNKwJTV4YHNP6MLmpx2cvqNjLxxhZA1o+AX6WHI2m0DlvBgAw
qxRzwYbMM2jQPjfO0JNJBr/Sntugan9Dcae6wPGDQIQq1YmBybMSFAhYDgRJ
kSYtN19FZ6b1nvMxU3wfUmaokFC+37M2WA7ScXHM9EL7zuuv1RwwYb9Gv+ye
j+Fc1YJ5y73mOGFcQrsAT6siT69PGuiKTECKjJnqcuDwD+yjhupQQC2fLqxI
dXjl5Yppm75n9FlkJRsRut+HoRWJzRezUIYQqojPDe1sW5pJo1i57B6Qr6HH
87Fx0WpKTXbmagPyF864yTWwk0WyHm6I4wTraCW/f+yaknzZvnKxb8Ex7UlT
AN6xwFZXb3RyeSlkt2UDIE1MZbmVknsMxXCS3yEKffy2RFmvUZEWDYV2K0DW
UH6ZlB8VvJbyRKmiyRV+wNi7qY0o4ysMgPlIXfaVG2byn2cApScUIWRiQP2c
gsM25B6VQ3pfsxxqYsGXkZ2PUQDfJj3F+PSpqEZViRZAmQdEbc65+Z4lpwwW
NeKRxxHpUwrZju5Ue5puyjX4J8HBm1132WVI0iD10+2fu4QBQAfahleHe5Dy
JCb9tRm/TfR/2IxdLpTcFYS6pMYk3dH1paXQHiACTGPHSHMbyiUPmSnbW3Dr
R2UAduXJDz6xpFN79KZ33vPxXUf1i/W8qFlt2KZzXTlpiprfpUumyZIRnYuN
iSIqPLHP4sOIGFFs0VwruylNh2xXeMgdwLaqF0EsFvA5H4roTRzi4McQ3oMd
zmUBVcCP9qMwNKP+MsL+/xAyspha4EvfG40Cpgf+SGZaV9Hjor4/hH8+DO77
uY9JcvE0a0NdEVBfpjJw3CkWTmR87fJzZ0jvq/RJTY5DoRtKjaYuME63xxLu
4VuB1+KBEx+lE5ArgDGqVzNcTMDoeb4gOn7Lfoh4E6FGqvt85tDgyA/9SGyn
RAkilz2K9ZWihr5lFzFJW/6Mh/g+gxVTPVU7hQ/1Gu0vDBmgdEXU33eHpoNA
es5aOh2mfQnN/7nd9qiPRjMWU/jtn2V9VVJ+A+XxuW13sPh4GjEjPpUXyZ5j
OfkdVws4fv5G5/c1sv5H5yhPScyUcQ2AjSZkNoqy5FoL2z0TE2PSmf6EG+aB
IuYP41TElrsSG4hWfp4RrZ1jVGCYomrlD0XIGkoZxyJ/DgxOYz/V78qTCAXY
jr0+y19lPivoJU4VH3I9PpH7kWWi6CSvXoych6LrrNq9YpDLPKXnEFSIyYoQ
A51otbN4TsMqa5S2uSeQL72kh4Foie6zlDXtuIzMPm9BgYzdfnHE4EsJKjAr
Ax6EwJq+n9caKEq26ZhhTi7BlFYkSE4dnPmTRF1HMdmDOxV5jkM5Nu0er5DI
khQXVjOnj6gJBClRs9o4oE7wyDG8XUq9+BcCvT5csnH5g6JlQuyGeWuYVqdd
A/ebBq815VG9NzcH0VDeLvxquV9ObsmZAFQXAT2kcEaZeC9cIuvlOJWUBD7H
ME1Vy6dLBVhcvUIwgi6vtzVqW5QnicIX/umHbUl9e+FfYaFwPigUI2ivzmWN
ggLWqBUq0C0Aan81Zk1N8jEdSrYLMgwGDg57ZNnLFvBdFACJxHlp6CX6MCf1
rxAI0SvKauVEA/n2J+njwvUhmNR+vPDpk2NIT6QrU4rqAB6251GTLcNIQ1qn
P1x9bu66M0gBfbmcznIQBdkT0gJ6xziUqUZg46SvM0XjIPpWTOad4fDoWdyL
gE6K6E4jympDBd9DnsSNNj7mGG+z6+p61ASyrq3NT9d5P9RGnmr+uTGqL9Hf
cQ8Y7/SO873hZnftKGde43WjtZfyaL79tFXf89Q4YXXsG1XGpTBnxTg/zVq0
bKn6qRAVS0tA+fLufz+/EpULfLu6F1TUOzSPJ6MsAF/es3tlYMTMLCu/+Z8x
2ZNbuvBpCs65dXBqix/QSdCTfgDdqqzci5WfkCOs6Dsfozhs0q15RxAsAsBr
dk4p5aLN9xUSoVlx0s99kpR7Tbf0jYJEOqZi+7LrJCZrc0JlnlGgjuBJhJqG
9ITV/8EzFfAZeZNoFG4pFzwaQyI5cfhGXSMpIPFAg0h+ERGjj9UIECD8kgF2
NnDLKIn5LeGWtqvEDXR29Q4q60YcifgJCSO27X68NWXpDl2miS8+/SWzfi1M
zpsdIY3m/OS5I2dKkb2uVkRFoWH8KHnfaVzpW2RNk6RLgSk7ub0NygLY4d4D
jaiHGvC7wNy06ath9th/an7vkNZVcV4DnbQ9Qn5k4rq713yhKJHEEkTvISjr
GjEoxmMGlQx1OqO9Mk1g1nqn3x2dXrsJDR1yXEv48LB5CA/inpDu9tfA4u7V
hZ3J0GkODvTx3gytxyKP6GJgAgXN3pDyTg7h6L1gvBoXrsCwb8UH+6hJSoKR
grJbhx9PG1K9rjFWkjmDUm7/Rblo7Y2UvQaJqtaLUma54o2YyrJZ1fTEA2t2
XOoe3fdgWJIqKDAEVxX34ILcNdqG4vXVlfZ+M2Uh7g+4/o1RaMlVoO856jEa
B2ZVXSW+tgayqAkPEhh/kT49O99j1mboD5inUBhkAp9I0rdFWlh/GngpCZdi
tQOsiyPafQvtNcpK1H2jeKiUyz0weGqk83p75YtFXclOk0oSaY9yMrp6l4cn
rqpyPy2r5oAO10yzDHuUNvuvKOWzw/gMAgtIw5NTOlzVSwPSM/lE5PrlPrwn
9BOGg0lWTGIYN8upJrpG0V/H+Ui74vTEJ6F0WeZBkmxIsSNHQKFRupD+C5Sm
CtE3Utw6/3C41WTAzeIsvznanUBc349qdgUL7GAkS8uREmDIqf5iU5T9CCFV
7b0alE6lnRyt8fXfSZLqPrN6nTwU735EUBpFp8VQgly0Ft9TF6Pa3DZ95K1/
H51pQMWeDOuT2WcyJTxW9hxpzEUNYirTf3Xt8912udZ+y+H/4GtuScEsD0mj
wJWuwYS/MrlDWko/YY0yzx7s96j6B6iWX8d33evbSPf4rJgbwsmNUVGD/A/Q
ME56qAOPT6pReQFeHPKEXB7TSLg+yLdmw+LRV59XKr20oBCPM1mskuhdF0Oq
BGwJeZCpbRu+udvK8wgwo1bQTg/RkLInCDOKNocmMC+7e2PMq/xYJ9EvjkS2
zhYJV5gguBDf7icC4oZyrCMYHiZHqzl47jLdyxOpYR2wHioI7s6xxKpqRUmU
/AeNcNzZeVvTs23JY6TyEh2T6ylBy2710592LOCz4/E4SmF2koODbRlmeT94
ZaxtMKZFlysGOvtLNnGraNRXK/3Pf4tXjcvOS3INVEdTJZNoNmLg7l0o1k++
lRxbnzrdfFlBduvssGc2cdj51x5xAK8cOYlQQ1rBUnsJfUUo/+6plN2LPx1K
fY9fkklduU8666hCc2Y72/989Cs8cjfWwRebTYSmSeUsi2gp9EDJgITR8h5K
IFVxIU/yj0EJYhmqNPvR36mlQ+MU+w3qVeSJHPzI2f0nTAvrw1UbZRtHawLN
8H2nkquqdySTX3MIH8m5KmxjDi9WY8JNOUS893+4ZzJYYdcX+u46zJMuJZiQ
o8ruyo97rYwVBclKmDno61Raa6e3YUn4qPf/IjzNaP0nkgWzwybhH58lOEOW
yl/2Hv7AavbSsBkhi9/LNqavwFtl8wQ1mIobSANkwTy812/vYRkgKVAwdx/P
kCOOq9WrFX9sCJTYb1nJIlq+7WxLgSrcxHJ1yPaXLEYPK/M1tiFtFdGGI47B
rvkK6vGjSFvkE4HZV6njmdwYeSzENqFHkFabmpVr1zNIeiqOpMr/YCym2qzD
ojzJzRdn70bFNt8zJzB8fEYf3kE5JsG2Nfp/PAqwEl5U5/snt1UZJwQeu67k
gUrrPrUc1h2bCyII2wHuNS2v7Z2/aeCt2AlWoaN7VvsqHxVBnsHdWmKl0Yn7
4IC/Ynq3rLfBZmoZYoSp6uj3PvD4PKlUNbEr9rqgmWqbCPyaPr3SVKM26Xm6
GVcRiFTi/Ea2JaxPQZkhVcQ8+edLZRVgJu5LBpdzFozjWz1zgHZX7D4IHxl+
XQDXjJtpdeRYb+Kq1oSaRAvwdO2k3Tz23RSKhaXOQTmSqwcA6kXK4ReR4FQs
ya6SXssYAAKem7lP3meOMTf8QOyxNMSOlDzhDytteOfnMBO7fLwWxPImBp68
wsbjQ2h0kCFiwt1MfP8Ly31OjNMxTu6tj/LWufaCCyMTz0cIxSfsXVYVqPDh
BhjTcaUu2m+zwPfqGCiXJBhimQk1j4HORJwlBZEPCb97c8J2zEk+WIBzVwTk
6ABt2U8YJRi9Vz2wM67tuafp0EJBQeiUGhMrw9pP3WZwW8OBMYFS6um5vvei
p33Eg2CLrSr/vKfn5u0Rio+hCIuhgBFemSQBIOAHxA1GWqXaW3DuDjLVv5eY
A1lJ1K1IFAgw+opYW2QR/uij2QOnZ6V7WzMqQBx+I2Hz/O3y+hQPXICwtvUb
632vLo4rMX8KVWWpRixmhvDfrGnpEDOkLhVt4BYSAupiYY7gq4Gm2IAHOSDR
RE06jwwPnLlekGleqwBkqdBdDTEnVwoMKp7DA8l9Uak4IhATmbtoUcEX0yAc
Bh6HcEvW03gj4BoiX2Vquuzkz2Ykpc/9KUd1dBkMeSarIITjHaSe00YMKCOi
/9wfj1bJz4+HbxAuZllrkdtSTAk7MX3MeEHlMay/sabKkDmCJVj4mAHJt2if
oePugTVHc/WFIxrf0GxwD3NZw9dHo9+6XaqlYzu3TcSMpM9U1QyAm3kl236c
amZnpKY24Hz8IoeR7Q/AM+zKtMDdGrGRQYaJBbJuMe2DUOe2yD4Bng5gCorX
NRWrJOmYTACXlNoqHHv3OHrGfTGDhmPonZQMCxQCREx34mO3u6Ui5oOXDMX6
x6F+B3EEOtW5Xz8eJbEnfJBEkBeDo+ujFqbURZ33cAfPP7Xy2W6ObjkrjTsr
leqmQGS6M1fG7om+KdHXwLTj+PbU6WCwkGVSZCYequB7oNEuV4vyoiiNRJ1p
Zpe/FjXtpbt1bZxOjGv+H/oZHDCiGRtu7DzdCCnKf6AEcLL+i/gh+mZMwXm6
6oXhD8PPkrDshCKyxZ3bv+/QBOGsIqBFY5CEi81JpPSTwQ6EKTtlphErq7tg
vDRW2/n52toBNBldLEQxFHftfIJe68qiGm/bLtAbD3OsRI8/hciVoBcd9jDl
Y5wUqZSgzhD2p3dIK1AIG3GyfHVCAfuid/z6gqGmmjY8DF72mrkE4mKd22re
FrbJk4YVtcsmMP48Krp+Wt4DYvOna0BKGtesEMJayrkwJiRxoovGWFLtOgEu
fyA9AajY3IQqgb5mOmabT8RhHCHwdrBI0uxaodUIuMvvnXQgP/K2QtC2kNlS
dhiyX62WwDyvNAZoiyY4cwS80F82E7Wdwxc0aKah3XmsfklXnuC6nBFl3c7J
3kj06On079lz8sbsxwVvBVdCtn5i2mZGq0c1wCOG1V3InVDMUHWi4e7sMFBg
EQAB+boNqA3fPrNQ+8ejLEEX//F/Ahsi73LqsHcLkATfffzTTKnhrjN+mMS4
wOH/kvPzRPqWvAGvFx1rwgRN0v6C66qpSiecNkP5SSEcKFFiKlvsjGo8NI+v
/o9y7mHyRYw1sAE8L1apv4AhTN6ivl+DBKB4dNIFQ8Kz2RvBGSrpJsO07CKq
e/M96kU7Ly2uG5WTZoVkPDr8Ts+poCb9SgaekvdKwl31IYe34dYqK43uezlh
yikGcTVbIaC2Jhvb/27SZneteltn2j9LIVLtABy8MFvnWkHB/DxLLPXoonUA
ZJNuSP++qLeg7BREJl/I781rlGXTfQvzS6xMNOBKejpVMfsAONY3zqG7gvTE
Mc2ab/X3n9KSsnzDCZzkLnw+vrx+tjdXJ/5+X09DUfCTMCI4HI03ORA59GFo
VP3feOwleSqDmiTzJsXZn770kNsjAGEVLV/6R9nkLn+ScZFdFZnQm4I4I3Ow
bF+BcChM/3qxHie4cU0C+G/5ANyF9sWgmxYbHPs0jZVJbrj7y4bdF4+fCVnl
roSqvGlSo/ZeUPbn+uHz7xabgmlY0T4BJKAPVzqRd917Q4nZnbaMNZpbqygV
Wb6OMr+AGXq39+RRDXbDNhzRQUkCoHVcuQg5UuHdjcG3a9ihxthI9+Fk3egf
l0XDxX9K/JjlISXxqUblBQ6yn8dgw3QN/vkge9Pg9indakCPlZJNmmGvYYdB
pIXONwFU00W6w9uhxKsEl1bhgQEvO7zxmsHeQXz5PBBm4sEJppvQTFLpauzB
CmUP3p15WWSLxdohfIJgACK5wC3+xMxKKrmcWRjiRuBn8QMJUY4sFldZM0ZN
FNcCIzpEwiavzUFtfdBWCse/GU2dToANyzMwAhH+AQYrgUy3mQi3XJrdRuXw
PU/9kyeU9cjCJWi/7NUoK8m6rVvjGNXjlRdsaf8cAUJhAsU/+hSdzgx641Xf
Myrjcy0CKvfCC3S9o5D0vBW/Y1EKtljDGtkV8rMmXIUV4qcxLix8rmAcgmPn
XPB9/9rWmoOX3qovbi+kRVhB7aTpyRcz2Ks/U9V77FVusR0n/qVFaylwUjUN
wtCT664FRgLiLgrXdpaMY0HtL7xcINLLor/7XXOY20qrBHRhkBzJ8+5KU6BD
/cXrufVRD8iExeEUNGdNdVXiFHBEO2Oqv6bNorYWPZiuQrPOEg7jtdG2Z1yt
XriwjEq2vXTf04fb0agTTaycIG6DKKF8uH08o/sefRfV+44C6OHh8z0lOp7y
9tJWwII3hOZCM22NjK7Zp7+a1yXGUHp4NIvoDeikp/oqmNTaKAba5JauokMX
PpV/o91MvyhdO9MVrfA6GTklBPtIYA+PNWR+ic1rBH9t9y75XWGnCyd4x6NL
nHU3snd2V9R+0pXebgxf3tt9SQW1ok7MYSHP3IKAqiQueXhaqNBSNQ/ekbaB
r9jVIWpOsy9zILYVX94HbY9IsVUHB5Wsw8VTZRWn8VgoBSSSGlUnUY8lydi+
G7AyCuorn9hOqKsHGlOT3ZOSgZw3pY6UesghsxSTf/5m12XBkXDBr2FvS1Fn
zR9dzmSmT74fgI0ocQxHYPrlKgLAEF5aAM2zJVLrCOezV63674+XDPEh6Pli
F6uq6qSBnPzf3KxRFr/USD9mwii1qyYbuVCgksVJEqSgTzV8NSsUs11QguCD
YUjlWJxusTs/8DYQm3C9G94fKIpuMKro9IOSyva6kVXgFwEnHdR3lzdjSlPJ
48diNC13qSCQyoMjXUcfmIgu57BC14jrKsG+1yZgQOzLHt+s5GPV+DKkAMbm
kgP2CoSudWmBNMbH0f+TxqB3HsQNnCQXjKuO4bpiHpqulDAah/Pac9g/kzJ8
1E6ZJvF+EcHdgKPk//W3RD6r6HeHaJzswIdCb0ICCOPqEQ15gZUGgodrD+KD
7DIHaFpSAqjoSR8OwDfx0lJZOsb3BeCmLlIs2bhWFQ9yH/ONW3uLcfP1Qi3I
JtfcRBJsyzKI1PFiHm9bFcPjdx2TBND91e7PioomF0Elxgusa7qE7Yh2NHpx
5+AQprcM0CyetAKEaiOxU763LDk9We4Gr5P48FDePtj1zmzzjhb53KT55V2U
8YYGwU2gQrq6jm7pBCnqbOaiD/fOAjr3SKtPl4OGj01crP07Hie7mYzoAI6F
s93URPuWeTQS4uMeWL94jrSuRPLG37lw8j+0K+8lxQYtqHsigXRjt9kqvwbn
Im854eFolc9tMqGdEVbW2qaRdzow7BKZaXIau4RgcciYkYBJq3qAq3uv6TrM
eq+sA9sWDeOEex1WTAA4Jvu/CdVmxRYyOx2FYBnd/W7Ij2fXyOMsiHljo+zO
j+MEvNqd2PstB4zzKf0Nhpa6lq3lfxbdqmGDM+e+GkmthkbEAEEAT/3ccwjw
5+pp0oxk/RqFDM457deIFXpiyVajdhPqVmIEkkqc76z76uJ7+lMyiWMiNxU7
NnCrIwb/u7AnOlhIqLSaFnxazmhhDU15kOti0AdEzOkqB7Kj16SSizEzQsPW
IDRRxCsRkWao7FvRtw+X0sYayATDyJnzy5ss7Nj1uNpjeYpYufLSJ41ovTyx
pc8UcwlMAaK3UvkFHps++k3XWkyodxhVwnYHOadWRudnXMJtMkU57bYX0tRT
MO3XUHTgh5p2YOMdVSn2/9m3FqZp0auHCb6vqIB7VaK8dapuaQNkWR7KpLCU
xq3j3Yt5GZ+PQHXQNBSQmgZa4BCZ+dVu3971qquJO5cEWQ578BjI+lK6iRvP
cejTY4D3m0qF6xo0k7aiOr5oOQJKvnG5orfZf4JRmFfXTG5gJ6ieBoHAuOUk
r0WiRLGDhx+ac98mMpPHmWJHap17yL5mefqtxkOn6kv82kj4NhwS9438agHO
m0CsY6MCwwhIDhbxPdii32Is8WRk1OYK923Kw7EU2OBcwPl1kT2WLmc939v/
Gh5CZUtgeRpOc8Y0CvmmhqHglbnDgE8BLQnh7M3cNpWZwXUtc5M6KW1eYo/R
dVtfDz2dc++9i+xPnGxHOTqyzQtVdAJk36172AqdGhzCwnNWFzpmlp/DFXJT
uNw/2Y9EIkU7HHJZPj+akSso1jssbukw67RpIyjEdd0hL74Uej5CPY3flI3Y
msnc6L4Osfd3007vf4RsyheMt3ALmD/dEVcuYgWevkH/FiCD2Ws8l/s=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGMQdak4aeN3mzASjKx4/WOhxWmNT3iJsGCEZZZBuLO3ARvRjT8itb/HIArOGCorCYrqQj8khltYn0IgwlAkRt0OC6qRgK0Zv7p0kuhX0MNZdXjrm9t6w+7y+9vRlKnJVMWVWRq++HfVMVbpWtQseaPgVraf5Jd6yqIH2q0SgVjSGhWFbvBaqYsibjFSbi4CJUXAOPrXQ0qDyyro6JpSJaZ3eaIzQM5jHeZ3pqylg8QR4SYDgn+UaR60lO3v+4ULSzZfjxqdXPkDkWXNDAGCv809Dr9ccvGkSQrupPcI7KVv/HqWEhSBLV27v3uBv140qIU67YO7NT22UmSOS+jN5a3QSWXw4rdzxBXDf9gW98FbWkyh7Sz+QvUbqlbXQxsTlBY+YBlqdzWKE8CNDXJGRYOxc6vWhNW132FeO0EmweWzoNkPzYJBxPUbmtIii4qxZGURwWY1Ulu70fjS/jgZR6+1Y23oQpa0Cq+inoQVXiz9nLX4oylyqgP9dPgz9xzrYy6ou/X0TYj1ZmNgnnFuzUqGQlhFSuMyOKi7jpcNNIUbhRsrvoV4IAatdSTDKQq6J06YbBkkKkIRLj1w7OA75gho5PIFuZFxUjQHaGhcNNXpHGDOp3vwW6td87z0IFYwERZDZbafIeqmKGG0PojX8oWq9DLH+SKObzmo25Jbhn1H/D5qBI97/55ywVdijPwGf7zy4piq9yS1BfPNFuAL0oafJ5rcD4zfR5frp4H1W2ms67YDhvGYa5XV6uaSkL4wwm2xyEJaDapiNsKsmNgXkP+d"
`endif