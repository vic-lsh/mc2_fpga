// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vmMbj1AnUdqEwyLUkSCdtGawm4zo5c8L6iemVDNslDg75NU/nk525dkRAa8w
fCXtGuDMxe+JdrYn5ncKtvdlePhZVbHXUTdqDeuKK4NtKFyVPaJLvpi5+pZ8
9vCTVa7jV79xomnpmQsFKmPgnQH07pUt70yfoWY9zyNykM0faN6VldIr2ZS4
TdfB4Qg1E8pOj2DWEFGc+nD4b/mD2OuT+Ip+XL2rTfrrWRg+La+PRfeJDuzO
SsbeVToC4cC9Az1WVdNHH0Re6ke9HVqIXxUSptSrI9ynbgtHf6SdQt7qlGBU
wxSN2Lr2F3IdRTtilIS+ZLKDLNoeyZz78lBdeoMU1Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AdLxs+yBVcYCXmYZhOeuy9ovfuz8fncflYefKrLcs8XfGT4rQ1WxInBq34jI
7OjUzzITXqhx8hiIl95TuvCs8VkYfVWGQANlvGNAQyTCvFsvmO/KMTxdD3Y9
kUts5gd7f0CA59Jr3Ly/x3veRhf0itjT/Ea2GOCrv1Ivj4trLTHXAh2rdqC5
vmLP/yvE1JPo6kw5fv01WDUwWCsrrbzWnoh7cLUlMQwTd7sWW/BJv0UPG1p1
p9l7pTPIHPKeTW1gRzzy2QNCmm/ZbmuVSoTCu0cF/3KoXH151j3CzIdNI4+s
YpYrXqOY2knLUYi6LvnkfAHJziGdoEG7JBGhLR41Zg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OkWFWnD1E8/w6pG83sYxnao1MZmw2TjJxXpPB90+BoLHZgg5JGEuJNJDcdkC
FGZ/M/vsqzSyhtc/iPIVTG3ABiDMSg8e8K4AtZ0nLz7u0daNjuVQ9PJtGDQK
lrUygO8DVq4k8520rxqOd+pS3cLa0hT5gA+da5s8idNCTpn5br+ZDxexZcsy
jn9TT1nFaBhprFfP0UFW4zNWf+JapESwqFNfjZR50xhEhex53ESdt3795i32
9/t0id0xj5j6g7ysgHeBfKfBkuIcv7dlsOC20/mIqfhYjMdGpqV2H1CpPsdz
dd6jFnf1+lx2eivzpOx0GPXzH3hHnti+YrEohRFSHw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZSB8++sYfstnpdxJQI42m1VaEPmHo9jYpGWwi57r/jpr0suYvvfdpalPHRZN
eyE9/9SbAESvn/Qu3k2bogqEWOMB1914/WdoULdh0z8Aq9QyhhLFerYGUCDs
qFc5pklSYEzIgV6pR5JQb+3h5sVdCvm4EFBem78spt0y+X4wlwxd5R/Z4n7T
Q0VTRD/Y2YuEtTzmlfz7yrb4oBU0Xu1nHIgtxrNvu0doFbq3TEnFEOgJnSUA
vXZgwWCSMLiW/kPiiCmdG2KYDpseK4bIu13YxxnEo7mSLJ3WQCfW3Wn/9kqf
4kgFgpHOCc15O0bEjWcQypeIzG6OmNj2jIzzMavs1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hHRbW1uLtk3IfnE2bTtGSgAz/73DTcWhaNL9Enk0yGSRHPvYZir2Pvyz4fN+
rTVQU+Pl5Nalx3B+VjkT0t4FtRbfBUd/ELgwBzZCrJoGIY2htJ3ZHBtgd7HU
Flh+fbnEtT9RBHWXhr5l2QDQUcWuSPXln3NGqqE9ozGC5A3Q4lo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AbqhNJALW3BEmZfd02dQ+Ik4r0WHUVbb/wdmFk0lFs22z/PFGOayhdp2o/0i
iPhLZib/JWdar6vmkDYFzgXviuarfy2x/MAmPfouMF3+nEavON8JcSmyDtSp
bAdUF/BhdF7Np1R8ZTm+hJego0cOWgbkDYmsQqiZCJEK9gHJBPm8W9W+IN67
AZP92/FSfaaB7tDJ6ZDd1XTcYM8z+By+qvo2tHygMPP8SXqcSTplPuU9pE3s
mHiJ9Le4Wz9MfJS/yRpqmQjd41aAvFtYMuIhdNeeHH4RLYNcjHOJkjbtbIb3
GflCHxmJ3H9MZr5FTMU5Y68gYwfdXWevhhXW9lRn33f7W4NIuL2NAl2KVqpj
efjNJcInQon+LEWzZ+GvyB61KNKoeqysjSuptFnJrp8b8k/J3SmxbL6iG6yo
Blsa/U23CbkE7gpCQAZHMAGAVc0zsdmlCrNFI+ZwbTEVMVh4uZOw/ERE+aqm
iEC/NS6garYQWibwQEPQgCZQjRoLXbud


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hb87ZE6aWQmIt4eAfTu37RNnyHW6ucCkJUbd99yoqgJUMUOe4gzCW+D9mSD5
KhsUuxZgqWac4rNijGWOXNKO6J05MoxWRjHifSIlrOA9OprB3uI3y23Kn8nI
GwLpARID+OzklH19duw82N+2UR9DP2QCxqTMNPf52727FIeZusU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ByEFpUPHTVZef6t0Fkcz5XKOXkvhVXJ6I1pIZJg8KESlLDWW6XjiICK3941p
cB2f6bGmNSnET/CJ19ylhMzFKJyOk6mKOQywxF5oEtQ/g0KMFy/O1O4lrlud
ab/hQ7IzKYQvZY50Y+zUuyYTtN2ACKn/yrT6H8Njk+LRoi08OcA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
gH2fwJu964sXDsVBgNCp8xtx0dEQT4bGyGK/8oLu3VlMgYWhygdCuFyrAIdA
P/IEaUlwINe2YClimeSVwYJ3cFMZJF1VhjjVJzvQkjalmILv3u5KlFeH+KRW
be9EynkUSP62na69lpN/HWq2Lo36BISWsHZEhzyWJ/Rjpr7QOqmUgqJSi8og
yWzaV2j4OCtR4/6Pwlhrw2pVdsbbj7Zr2yzMwIdRjIhtY9P53xqMEfYN7fh/
eELIT/FGRPpLO2CnpxNY45tR8XPN7TqbyDPFTRSFvGKmo9Mey8ZzUnVtFAZq
X/GVQZ2k3SwExs6KIZVo29lNzvrqwOQEGJI9u6m8M+tVcLyQLiVesJvXvueR
gvco1gteNSlphsF102d7GQWcEjKyjKArefxYDvIlz2Jv+wzXuHwUBJ8KfpBp
BbAixJ67U1/j+K7Vy9SgFoj1EZEKCfFbF/seHa0ITW3tpC6i4I1ClNZ6nHRG
RLNXI6p7u2+/gPPpUJWISDDXWwqLMc19ySrlLlOaHrVhUbVHWeorbzUylrQO
fg961ADItYIAHbEp2S2WeBnmoWQneSw1NOXnHu2RaI54XLJrFeEiVQR8vokU
u281KEV47uCWIqpwoaOzw5OkdPz0tayddGI9sOmB1HqbDIpEKOD8m1UmRfug
jRxgY1RTSs8JCq+oolmuCNhtJsYVOvI07sddm4ko59AjazhHceKErnBg+fhC
8pyD66wNzCEJKyLEyVL/U9UdCgn0mIHHzVr/2hdpijXfC5oWzIhmXssxaXin
wO/FqkzLsuqRa1jjQp2avlfE68eR4nibyVIWezTGvzRz4iYp0VMOpMLr/Mvg
0+Td4ht40Fy+pch2fHrZA+DMjxbNlw2UsCOKSN/qD0EGzDnnypEFWozIOxQO
Q7q57k/n0AP/eynGxyajtLcNwK4mDaHW46lsGjQOALMYID2XUyPCxHuwduRu
zBl4/yqums/XqydHV+Pog3S4nQvdvl/D4JZ6VOifaGXd/LezH4yKAPtlKo4A
pc3ykUktrhJgSqyf4HViaDYGdKVpcEwAIf+Yt9Hvha1UN49nfZCGamjOxGQm
LDcZ8qU8SA8YgEqzjvo9Tz2vaNIEevMOvDmdB/MD01C5WG3C+BIqRaiN4d90
fLnKS1gYeKEt/VkWB3YJxaIvm290kQcEHfgmk0ROE6hR7WHKCuYCXHz/gXPN
74y3Wnc7OFC/yK3jPgIiEib1SOzTId0iUvIFow3vlZPPyZlskZ33K67jrVHM
8ObWSwuU7DpBvFqxBReH3TWSblHL4zLV2Fq/zW2Bnx4nzj/YrJZgYcK9oSNl
N7p8kZU87LudmQve9ANHnmMYQw7lwsEGN66j5vu4wr+1vxpDUC5dSJvRvtxQ
8t+y0jc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqcTIYTaY8qvMoCFZZWBRl4ZWhSiha+4ChWiB05sXP2BwExj1uWQDQNC8VHlvmrewoG7yqM0lYJqMx/6OVaHcO+TX84nuQLsQNpP5mADVQBI9mG+Yo1NO+qW6pPHIwcHdZ4cx3YuKCZESwXdemH03cFapnSbsoP56Zd0HF9h7YRGz/+uhCGEXOTMnrlK+3yWYl5Kg3EHaJE1p2JbHeTS3B0eCN8UdDsKUHWDRoeITVUXnByinNQNkVzBTB+fOrV5RIwAE2Ye6XG56vrbl8D9o/eT/nowCiY999PEK4komouM8NAc6QgxzWKaNtO3wpi2EbZ4QnJuBktgLCG0JuhkS1/LG6cSeeDJBigd12pBCJu7p66+MupyKHMheVSmTxntYmiN6O4kIM0eS+a8lQZaUkyMrB7218QVPa0sIKe4hnlt91yQBzWsIyfvZQ9a+A2CTlH5EIBgwVLeAdLl9r3iHej90ay4QwNDdxPkeKeFa8cYJ6njmmZugv2P3OBaYwleAqmVf2pPR0gn8RPuHbDVc3LENvu6Nla88RLgROJkLIk+SJbL4VF7pZrtyt/FG/GAiRmjD0S32rp/hkGRSGjsnYx4gYx5eOQ5DSbe25oiBJgYbg34eTlagJtyHmpag/1quK7xwOo9qkOu1ASGk6BGlNZJ7QQb65QtEsMhH7stUT8mTy1tOMy8C4A7lu5zNJ+r3BJxWN4s7tJx2h0OT0J99n+JanLJj+6KORf/4mWSA/9qNhmdDbHKOGdloK5M16KNgt2Dp+yPdyw6M+9GsL5kNhrJ"
`endif