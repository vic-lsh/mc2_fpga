// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oSltpa7eL8LZ6E7P8lhsmwOrHFvBk1yF8ivWpjPpogOGdPV8Tfpc+kHGPVdd
l93/6xdL5PwCyaItEKY6XB/IiY4ww6sPpuG0q+atJUj8X4oMbbKG9AmYzZB3
i89US0FtHqVZsc5KodQdb9YxAtGDmBnHZBQ+77QCxw8pM8sMU8TM20NDIX9L
muDj/ny2G8SUfeYVKHoviJkena+sFvof+CK6q/rDlu6C759hANUuCp0cpoYR
2O3Yq3b2fKmxDB0uWCQNk8pl3GrgJOGRqxEIYrFPFlbHmasy+YWqs5Tnlzqs
e6g26tY+K7AqTEY6ml56RUAxoCa3fjHrGbbiB9X6Og==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BDSsMUTXCyfUtohVHPd29Duxk6qWO5VHTC9gKxBVZsP69p4kKiQmfG/ShBMT
O/vSBc1KDNXBdXTSotiGHM8/GCMkf7yS9nAwDyBRZmiuV5G4NDKD8bEBLg1d
3ajfBWPJP2YRu50+mPp8riwI8NLsWl+rqN179Bn2v1Re0rfqyehRYfUH9DUI
nt7XjVgCrVQfOJZRCYnpb6UPj8XSOnB43K4ecWWlAYQnSMOhbf39XjTLg1Bt
0aKQMPbD83EGmr/tnzdgUzb3HiHqoY7DzNaO7gDwC8zJk8GDY515bNayHpkt
uPKfZ1Coy8XmiHOYrdxjMYk/azlGFd2Cl3YnJKS75w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sMnXqjuiDMjGfmr23LSTFx74+qMFKoyR9e/kKER4hVDDFVhXIgIKsyVfhgpN
vkIV/g0K4rATgjapn3lU5ZPQZardZAcUfNDihSPstsAjcsZRFpyNC5GgGT4c
2oTc3MdI6d4dLF26XLanSCu4ku2g6iOcPUajXvCXrSWDPVijvDEOJk1bLdQH
cpKjaVQI22RpobAJhXuuVPu6wv8TKjNYczjeXQZG2jDsARzPNaGo84ts4A3u
ksYQ/j82qHQ0/xnd6953hSUZuqmY+KMrnEIXd4RUfC66skycCXG/WkJO6S38
gXX6Rzhm6+JhkOe2nXdpoSZGvQbikl+u4vofCVb0hg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qStxvxze6LC6DDuEBlusTEl6dXbZatD1qaQC1g8NGuzl+/dMt+1NoxW0rOFO
sWavGHNco9gACMFC4WyULLd7wZdeKJeV6kE8n25Q293hq3ZwXrWA5qPb13lw
FmPDIL4rWFJjJlVwb1C8gUysQB+oua7NnaPXZ+NPinK0QG0LXM65YuLn9lvM
c49B7fakwt9O00AixqQ75cNyGn5f0m+xyWFYjJQfdvaqoWi//QvV4Ua9mvc+
sjy0sucKYIP4+K3x/gnn2tr7clfFdtHatRyAcra6/aFt4k0pdV5ZzgEGHYjO
gWUTOJz2hKQUmWL64M71Li6yP7vgUwo6ZMhlnzLnTQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XgU4TMY+T7tG6Hy8oNWid8Xy5ams4OC6Sibtemq3KXcAM2e8iQL9IWYmTkUB
30tR5KiFZEE+zxSLFDuGpfkPcnFqSRcy4L7v7hK8DVkVJsdjBvTNsaOFzT3c
8YuYqWUyKO/+g77kJCWvowkvTSz1ZzOkUwyN3Cv4uJbg/+Uzqns=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Mkqq24lMNUXVQOjvdkfzzEb7Va7q6HW+62ku/UjDBmSn/EEQr0ND41jjd3t1
8d6qyLQCxKXKMn+LuuazJ5kZ4LMlteHk/TESFwUxClj0/HwqGWmni6/AgmTU
m6qu+7lb7658LhxPvx9k0RH9oN/JTlq1hyqBqrOHuNmSvXdQa9m8Q9Xh2rQX
ptGO5jUpNwwVv/ZFcyc1GE7d73cBIiXmWDM6k0Erng/1J28tC8qFF/lHkX6e
cto4K4dcBXlESs+afjz5h9JCkL48qpVnfwBkrIZ8+RGLsNoh+9b2WEdXL+xP
f+5SblqoO42FM98sorqBWw7+cbv3GkrxVRliP+LGuPck6Cv72ye8NprLFfaL
PmXEUrx3ecUkpEqLBOId0fMVqvMJl9nsNPpD/Av0aSB61cK83KN2DnlKxnKS
jgZ4W1iXvdvc1fBzgV/EnnSUoN/pgb5j8X4CdQWqBesPbJ16fLA0f9N0wW0v
OGS6rUBa/u1sNFTLX8ocNlvhE8LdoCb5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
l35YkTezqKndV0zs8UlDFRcX+OHkOatd8qk2LB3VdQhU3qzTeTqXGd8TRAhG
WQMrxdV4uJaW/WsCTlxfYUsvHSrKai6mSQwM6jkUnhiaNQ69vJOq4Bdxl/0j
8HkzoAL6uIo1g57Y0BLmOmJuP8c+jqDuhTBFZg+6VLkKbf9PiC4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lsKPtiIFih68QfsntjkPPx42VHfkCTIla8Zucq0phEnOWydN6WoXJYi+UlJR
rjThOUdFCdI66cQOxQoWQG7wZ/NK7g1N5ZBnVAunp85Cr5+3uiETra2tYZtl
7UQqdRcz0emRXUgIg3wiIoPJUa7+LTkLBz/QwnWDR4Ey+onkQ7o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
mkOXY56UPvdmxGO560oBqPSE80yIqYJRkcC+KzWtwgHRmjmiVAK7gUUQJ9yZ
FyXoohScOZ1MFAl6gCTNxM2JMykCeaycwykXNYP4btmzyR1+0NuxTvuD8X5R
i+9pG9QFa6YSZXOeUxzSmFZmJihMZCZFJ3ruYmF5OTaZTKDOtRSO0720SYxF
GQtXX+tmiUJyC5/aym8+CHpbAPGHeX4Mxcd5XCwz68RpThj3QsEqJfX+vU18
7ZwCbSlFATqIiIFh3B56IGLOnx3q676qLD7xMcnEv1CuQX6D4/nofFcUCXCv
LsyACLTZLoDGQTRVnUYJ03EcojMJhmOqqllmd+vnd1/uByuGLp+0OB3IX4Sh
+vIxuwqr/+XaIq9Ig08cD3k5UElzDf0Mc2Uj6X4EPky9lD3QBu5F8AMXG8w+
H0BeAPDeDoC1WyKJ1BTS9Yo+Cl7VMMk+p2xYx3OViqvD7ubxv5s77b/QLEO/
kU+hTlrI16J3avDwt7FhuHompY0gLMq5qeSRwolkrXpNY3R/61gfwEqZm+7D
aBWMf2yjq5RnSpbZhv+kWytVJRhdZVJf6jtTOpQEeuhipPvZlmd+u6tHQVmU
060FjPRKFzcStjLFhQTqMp21aUoMtZ+IShefu9ye0/3EE9xSLY3E6N+06Gxx
J4X4Ry341JyxyNn8C97w3IAzxMUIRWLNzmjDuy6+G75iBARKP6AW/kdRtV3X
cWIXQIsBg0AKtkPvxG8OvCMjeAzZO7oIvY7rkBiXT6XFMV6nupGvMtE9vjPn
hfdZRqgpkbMU7riT1jlE/x2ETcUKcaLtrCwH1wVuqEjmDEX+5JWzEBIALLOo
AC+E1mKW+sC8bC0V/drCPIfJT9bfYMAB6sR4Aqn+ryLsplg0IsVN/0gy6VpC
NMl3juOarXUTws+5mNE1GXSMqAM5Pomz1sL/A9b6SurSTe1tEjJnMnw+jy9c
eBLRAzk7URtxmvYeuK5yqKnDk9WYI78nmGTRIzgrjHDnjQ+D9RyWPhkDo+Eu
hVypNIKzfideCGyJXzeD6j0glSg0UtqV4tSSQXse1wD9cFDEdat0pKwjOv8s
aEFgf3Hhu72GarUQUaRGLg0GbVmhRun0rFwgImHaFoEihE2ksEflsnwGKEXw
bXU0ONvwD+6XXqq8GER2CkvXrEjXwIKrdc3BqxdnQH1qqln8pa+DMmKuwwee
jYtwCRuYmek0cWQObB/WroXZyd7O88p2hVX6htygvzoXJ9yoYIZmFSTcun6P
GcIbH/dxAePM/BZey3dQcSePbVgIQigaC+Dv41iCF3keez/c9hCNq4H1r7p6
bx+8G7Wi8OPU7ddztRhg1ICz87uBSnI0z9/LnQ3HNjrHEAg/OFjJDieiW//0
KRYLIrpvsa17cBZkvO/jlJxO5aD3CUlpIZiAmg3mWZEeGolLKppjNK0GIw73
GMRNOtPhO/hCnq8BWti2rbZZteLCxOK5/RpCxrAgy7jWfWoRmi/nuJlRgq47
tRs6Q8u0USVy8D6mSgMmpr27vcQSCX4me90QU75HoauhOsOfoVnS9u4CdkdW
i8iMGBmGZFwdjLJje6YGe0TwOb7wmCXDSXtz1/h32q+5d2veqSye2650wH6v
vW1v7JWM7Q7qlcOtGCYit45rq7HYQmnHP6l3lIFYvR1nuOhMmIWEaVe3XtNn
+Zn5esGP6qPYjD0YBJXbHTxd5tP2Pmye2PEBjMH/V8QHtb5tofDtXza4SRfY
N7npMaVGmMPWmbrsdVf/Ry2BLaV7xKw3aiD2k7FBiJDZWnLRXhdH771e8nPj
hjhECLtAIyCMkfWyRuLY0QuyN8JM+SjsFCv6ONNO7vkRWGh4UaAxVJMCEjfk
1+HsI/S3ogAnOVChOrd1MWyryN6qfdehjaa3WMXG8U9xTqak1zcOSPcCZ8eX
xcim1ggqOLBIL3oYSikYxBTjBMstY1/M6Y+0toCnEBCP4T9tBjSU6MDv0tpL
uH/M0oe2f+e8i/UT5JaR2t9tHfdkDdhcPJij85vcT1C5NCYMrdr9QDyRhUkQ
0R1RRb9F7IUhsXQ8oUnkpiuX/CWB7iqMtBTB1ZxEoCrNb9njmvPXu6u/BRwO
uD9ISRRM2KX/RSJTCls8PEhfMOTpkfieYe1sJykxAK90TNRXkyPrTXx4wf8e
txj2hMmKfrHFMqw8tVzDiH9FWWPy0T3D3JyX4JUkSo2fBKaksfbsvTUQH62+
RUd8cjTcWd9fjweB8HezcvgBNs4LJV3gfjBnvDinIBtO/gVTpWE2FLTQuosE
bXUohXuwajRodXtdy5Zak7PsF1oEBmXANeMYVXqRX34qScZYiDRCIQJUv7Y6
6pnfkx3uIbszEy1sTTAplzlcINkDGnXfRXFf8Uc0EdRrBB89clJEuoT+Ypj1
TmvdFjF5poz5aLOClwhVzy/WSFCo15HkZF61Yj9iFZjFk39l+Sm3y+EL9zgW
IDR2/N5klrMs05QCqzFdt/m8tayLr0viJzVbvB2D2FUnrJXh+lEHJaF0Z4B/
oPLtB8EOmQ6X7BAVLUfo723kR2xRePht2yeX58VKZVtwByWmoYiY0ckJs0Xu
oX7CNQdJ5L9LeAmp4PkrCZZj3YcRDlg2tLT1O2miRbGsyHglwIJHuLIKvZ3R
QmTGY3hxp2Lv6iOaWVU+gKwOY2iflBfH3dnX/++xhLaTjtDrdrpU7D77fWUT
QYy2jmYBBSCO9jm9+ptVweYQHGyctNLlpJ367OAnqB5aeF3a9dL/kUcBi2bE
bFsR5zgyYl83HVjfPPQqykcIM1cZMDBlRMpxvxx9RjYLCY9GWl3pzbWhOCWu
yDD4kLSYVRqyX2EdMJeVB6755WdIbjEqVjBinZhBIkl35qIiHebZOh3I8pE7
WTu9J9YdHo283PC++FXZms1DGMnJKIBjqp3VHHOrDynPYD8EYaFaZrLe4Sq+
nlA1+6X5Mw68teFS5fDm2542O5nvBi1ez73m15Xwa+K9yw1E1jJeX4vBes3E
yFXQqPHc4DgcCVcJ+B9aJt6IfJhyOqJa/AINbbHqSj+gXSXKQn/XyDLGC6yk
JOFTqEPyZjM2jQI1ZcOxZZ4Y2ts6j7Dr5O7wCcZpeKkbJBLwbx0GVkHW8Cr2
pTtR0loNU2endoGjgOE7H20W97puokGpUSBJg8YFf8j0WcEp0qvdWUJB7hqV
WVW6nfcj5HQUSzNqsfomfYy06aGs0sETBp2cO6ZE05mXUYUmhxdfVbVB0Y9r
CT4OzJyNpkFfik4VC+k7tSrWVjnV6CV/W0VY586c/AzrI/RCgR6ppzogTMMi
LCIN2N1IR/g+kX2GbLhbnp218AL80I9NccoGwUmbjpPIwZLI6S0demqg1mib
nobtJkB92gYbKLF05KiTcUK+AGiTRzoxL4rnVK0tGsRfA4yhneriXx7pxkPw
ckt7tGWCoCVTGFPVJr8Q1a0pCuhk0cqJZc8Bc2FWehxcqbBE3na0gBDbiGsC
h4BXLKQ5FEzUF6oyRoAu+Ksh3b5iBcnSMpvlZtF7yVd7MUsuCZz7L7q0/2av
3mMT+nnKdW8xOUYVey/K6UZEzmMDaaXttTF656bTOPz5u3B6A/24BFBQmkfP
+RiZooaiPhWJgDPrMBNIJRjTkKLVl5ZYs0v/H4t/QuLbvwuE/y6Nd/X6tUzu
wrQj8XBkHqGg5zC1raBsefzk9II/DurOVDnuopjq5F+hKAa45KiCG+L9G00J
extsHspCQ9zXWAadoMxpzDKfcUMndtxNdEI/xX/OwlfZsrwflVz6t4fqw+NA
SlPDu5hquAq+vUT1ApYjPmH7KvVhDp8CW7HAxtNWr+yFW2X7LAgLJRChK2SW
52c4G/uw/NwfGvtU4N+HDMnmN+ZL4jl0syWOUxr/VRs9nF8pb5yswxF+BRFV
Bl5/tVfy4kzlOAAdWNqFV3xZtg+T0UE0dNBwdWZbKtv4ZLuMjzklNAaNZYyv
dNbFOc1BPyuhyv/+L6cd6u8L3lxaXOoecxuhiaB0LtwMgDiHoBACqaqabVyL
qhL6fJPoh+8dSgClZbjT8uvHDhs97EBbjyE/zIK5/oCTJ0sZ/8fv7GHPEXZX
S90UqXW8lswlfD0jaBk3G9qQB0EOendE1vjlTJGElikPGLZmLW/gOu6Czq/U
zVSS4SbRH7v2KDmPCeIVpkdOZdUtu3JnDJbXq45nEQwF4VfpraMYEfoquUNE
gcV48+FrSqqZQCph7+sHRCQqwK5Net+Vd0n+joU81yfVR3gecykrdw/WyIeH
JOuAEqaLDTLCH6DhtMbtocfQocrQ1IaS/OjS1r0C+LfDYCfTQ4PVIURTaW1i
jJOJrVlWYb74RyWjsJUxGXjiYKhb+Pu/6JWnsgpmNCQu/369rmz5I4LxWdkz
mzMliF51XWrMLinlzNPxd2lDYyIoYsFemBKq+Ib9rINrDWEEqBujf3WVtj+O
Y6tY4eBOdj7UfJ4WSfvDmd13u9pxIHioj+hI3PfRFk0eIjtcRknqrJSpkhZ5
nZwy5dc6JN8tN193wGO0oiOg7wUsGFlGPMYPQffma4Lv1odV126j2vIydpH0
vNeaJlEyUul6oKSbV1BONeSN36GXoHfdry3aCS6GCARWK+EfJEpLmIQXy8he
LLoFLWctP3kBgLEWDNDFGZua12qQk1NnZ3vXs1/twtYsw7ZlFcR35JqFbStr
tqMEW3yv0VZsSToM/Z7P7+CTHGTdYtpzOK/q0Ue8TRLbr0/8OAbOhx3sevIH
djugvbzYrhfukP+++XvrvohpRNF5Ue583XR0tqNo5Yx5TZya0xVL7I/bwgaq
ZRT85XlDfUSri6gnfX9bUoFryTzFqmZs4Z4oRj6jHUWyludqRS8PE8HK1SE7
5uR6sd5APGYrzl0HWCCpcyHCU/5fIEpa+KYBoR7g36r42UI0lpYxI74Dsy6m
VKSBrztL06FY+/z6VKiIAd96PVQXlISGsfr3DqIwsLlTP0gg2ju+pVRhM2m4
0FDa5vDkKnnKoPybEOEYdwLb7V1scGGPScUcGwxwh1IqaRZ7lNP7LFvnTPHm
C9G4cmmfy77DGJAtl0BMUbxHmnipdtUNN/v94RLJ8I6uakrBo62HHKflTNrN
xtkL6mjcA/KAqDL6soZVPLVd1IJu1z9GRSk0jxLel8idP84gmEZib9Wv/nu2
uId/Xpz4DPaBIRoL9tyztmD1+CbxCUQ5X805wdYT/bDQ4pSRC1sl0K4bbm2K
e96oidYN46R9CP305Kr4Yid+1daw5W3BM0rHD8gX3BolOxIfC9z+uo6KPAyx
7oxhQtklmOo+9BkXkszDQGpFwRMCaOBAJnBNYR7MWy8LErcWlwamhnQrcEta
gY43wQPgS5QnrCJpcaHiIVySTkgdVG/4Fhn1NeU9rkcKQ3NkGDt04de6MG+D
OplpgduvXQYxk4DylRKJQ7aMYSIKwdLCtGZaWPIS4hZEVXxZKPUpwjZME0u1
dd+2MqOJDe1ccpqGHv25QMrkZycePEB0FNw4CCUXLmEZtXMzbqzBy9jSOJ5V
RkzjSMQ9bTfnBrZHfuCStv6r47cQMMB4ec0AhlH2s5wqgAR39Afcw6Zt9tpt
1+8OtUfUD7/e+yK2c58svxncjrk2/k5N45/u4JHkQCez/E57OGl7hOqsuTib
xUyHk7oeGExe5wYYQRHalDFG87v/9Su75K+4Q4hmvUCtj3zl2qY7LjAxQeMt
YaSYa/0xxIo1Iz7MY6E9B5reS2GiSndbGX5SPKOYOnLUHQTjCP/+t5d1zvQj
CqryxesfDEXFUbJa46JYPdHJeJpGJmgXuuXczdJTzbrsnhVE4Va96anEDtCJ
hnyntDG0Wv4Yusdhj9IQyYC93mQC1/70gpQVJQl0Fb8zB/nOhoiLqOfhRMvH
kDet65JPBXka8KXK7W/KUayfOsxf2vep4e5MeYjhde1QbRSZjFLGgHPdK1ey
JrJAzdv/IVhnW/jbGqm/CrJ4pO6a1kD8gGuQIIro99PsYEi7/sp8yUXSPNXR
AiRWsOzEJmrGagU3bOE31JqfbHMFK6zOWScQVKwXlHHfZVFtynmrimfbcj1C
diyhm4sqfrVySLXxHCXqBQ9ywbB4Pk45SsKQTeeycm2aavi/rMmCG6K19smg
tbJuSVbtJigrVuFML2TipcsbonZW2jUV1ytU0HsX40sS3pS2iRzltUNe7ZAh
vUmmLg3UYYttdcnbeHwuqMi2+7w9gSUTyX6FX/azi0yHQ6S3qJOiUqeOtJxO
PZHkAj/mKM8FBzsML3xS0PmqTGRqqcGtqEuZHEa9mJ54KqY7fATl+JUK7a1i
M1xXe/7l4QeylpmTNDBNXtS5zrCN/t1DHtR0trxDGcVgMUfvtDbiCOF6J6Hv
BPqcJdDYxzQoOeIb84rriZ4rlhV64DpTEsYlgPrqHcMiIYyOSS/aaeK37xez
ZLDceFzsss2adD0sYCey8FnxuGrZiol5BH2yMGQiyx7GVLYLR8MV3mgues/F
wFF6ZT/VWC5lqgIxNcvFLPx3l+KpHTPZhxrPrpMimfiBQG9rDKDS9hCQvh+j
jHKxsugg+NyPW3QeGKWJ7wEvpI26te2BUhqFvHkQPTCRWiS1PLejwWr7+++l
Py3JM71bm0oGQ19tNNqMlZmd84b1J/0BF/iE/7imhASwOGGQBHmUbttIUOy5
Ed+uKZAaLMczzH/7Q3nSo4LjIskVKzj9RGnTTzmnIImNyn2KN7dWcTADXxWi
+Vm2+4jQCmfKsJ3U57j1DYkDzIfcv7j9YOO4zwN/bSdg15vtitnPXYH0bfHx
TnhcHAqLXpzISTh/FJgNN9UwqRqCAHbbwmRH/zQzY3+1uI5jAvnDw+TeAjfu
CKTekM+rUa+/XBUgxZJkW/6GZ71wEGKBPgj4/YbLnXFeynrD54COhvihNW5f
9HmkyzAZOfGWuIzoA9tr80PaDGKPSslphs6Pi/MfEfX8OxGBiyBV8A6+v/Q9
+tJFnkOTP8QJ29Oy40D6rJeRfurYdJ8TkT2YJIcDutyBPzjRFXpa6d952NdJ
if8DXualPah8hiewVEURhDqv3YegkCpZN7aR9i65DO7P/OzjYfK88Viqw4HK
aQ0T/z7KUTzJ9PfLqqDBOwgVBshJ0RAHDmRnR1aQyge5f/HhgNtZSsc0qOyw
+vhzdjchzNXMlWMoNnSjjNfYoqbCfyxcRqpZDjSJaTGC8BD927LOH758OSna
/E6OlmX1qZRyX4n8ljWYkRr54h5X+iLsl+1uYTq7lg6EkG7/zbAp3bFvKgJo
h5KpEZhsPUaFA5zQMpIxWHWVYKZvI6WdJoOBCWR64gYEXhPRBLRhLmvm1Ovc
8pODehYS03/HjE6+o7wbP5ExqpUSBmnvyKve7kAV7W05NbxbHgIJHXxRm/zQ
qEkabvIt3qnE2EmU7Rb8z7buuEpyAtfLYgrEaEGAGhRgj4Sjvc+9d7E2PeIY
D3Aa3ukxnJxAFDrWQTTVvXe3srDNhkb5FbCszThj7AaluSJi1sIADehtS+J0
RDQV+WqJmNm7mp9Qxm6a2LCFvTPcoHUiWfP/ces2zFb3pUN1oMR3RjhvCwSK
+eiJmHixNi9+9t/6IUECKxud3f2L6OWGlkc98PUnfeJiW0PuAjBSPgIB1kb7
yScOuspYMqiA0qrKVqoNeH6eQfVylGQD05AAYsuVXlHXVzbNC9Yj3gHjIWUw
49Yj4Qvuzqbtk7DY4TpIICzF8UBWsrl+lWHwr4ZJy2tZHBN4MkGaWEoTRzTD
EbZOiNRCrn2i26yTTKqRWEVVcky/JMzRzS4PW6QNZsVj349xYrxsVYVhk35A
u8MpKqVN16g54UUHkpxsesr123YZUEgOXFOPgiNNaeq1OpB0qvGkWg2YdRL8
XuRRtHYspS067qtrel3dO9f59gU83ZzjgkOCPefIcvuoG3cJLR1/QK0ecxeu
2hGZba3p+6lrrj5SHpXBDYF+X2AipQgFbcK+WEWOEabehp91NCXBeyqwEtm2
V6ACDbYCNaSTk7O1vZPO/RaiM9ejwHZsL3eyv1Sv+uZESGqJ6MWX6t/OZP/7
x+Nu8dkeBjDm/nmluf/pysRDJi5dHiqNocg4fKUlEpWF0sOxI2GGzkHLPna/
JU/4RzWi54vq3vYXGZoh3lMdF9/YWZhPeRJZQh3SxpMEV8hN63yWsBBAz0z6
ZV1cyLwQVQIaSsMe/4cHTxTBSy1dRTz+IB3QRDhXPVgmct8pAUzcAxBSwqCS
mdHH4O/VgiAu4dVa3wA7w2QN9GJiRXADVBjPH7EESlzn5CS0mL4EajMp+rzB
yDCKtjNrQJCTz7w2A470CB680sm9I1tjplAfEJEaZ38qA+1p6rAZ0hXlr19q
QYPdfsv76exSWCuW7X8FzQhdb5mXEzUl8PfPl4eAOe2lIt7GnEJl85A3rqx0
pQaH407mLzVJwTs9s/ViuF149YOC/A9z4LKIs6XymkVfBVOkz2xvVCxU0Veu
tAz9+UsJ9OCT/V/l1EqZA66s/doMHNwoIVIfoixpI6xxveEKgkYELSolXiD0
D60uTq0z/La8Pcb4cJlc4szcU6ul0CmbqVu0Dt6iptoQLK1zO3Ik4cPLBid/
sSLiFlLzTVh5kyMUIP51pLLRgao1jdVFBnnVkGVcgu+WjLL7BX9eAhmK8t6g
cqfI9q4sw3VC6gnCb45uyN4qKLBirpvUkVxCVvnY3xxMf8IhEcCXpufC7PEN
djauKT7rkOMYf2yU86lRa3/+ExQ2WN/NlpZBJu1u6ESpDDoQLffw2F+ELc3/
41so5tjpCibC7JP1zR18QxWbi5sgRCSDuTo+R7T/M12epGrvIhJFlF06GVT0
QQqKkSMr5mYiImviQ5nSDjsC37WW3EmfgSmI1xHgPub7eRO3VQcGZrDf0f0j
DvtJJITtSL4AmUcgZlH1ANWmxdEJD+t1HzHYMj1SFQGXYRPXqUmitZcvSBl9
E/aC0uMixi0l6ziZr6YhJZNcQiTWFo9nVgyuP4c/ggCmSyQbxaMM8clTa00K
cNqMDSzo7NGKBOWc9hE6PNqSeEKdAyz8dtq6gotxPLRw1+OIHqiJTXvsc6S3
pvOd4Qf1eN2nFYzmNsX4YkGqqNTnBcqz63gLyoZPJ5dCBjc0ai1EqmVwRL6S
gnHY6i0o5qrdmlhMh3zYtoL4nh9UolL1vMiXPYZvf1MzfZMQRa5C16YHabDl
Vilrgn265IpImtqYi1vRzwLzgkpuD92okF0GTFtKaND3bxLe0G+LYgC2OJ76
p7L5a7exmZLWxqxaOpZ7eUMiDGQEC3V1EwFsmgUfN7Q4nzdW8rh69J8FFLlO
qxPTVD52Tt3wuTedUD5EFox2qygoS04rb9O6lNZMaiasvDLPq43/eZxz92ZQ
A8esxfwkpssQ3Mdd2ygBNwHLq+/6UljaMpe/onpnCeitMJgEz2jZaIGJ8OBw
/CzK8NKrG+X3jrwDvaYJwQXEzRQM0WFWO2bzY8Lq/VUS1xtfs04y0WWMv18f
2WpKIW1HfX+b4zK7sgLNY1haVZxDW4uol12Tk35ZWnIAVd8L8kul1FxEmVS9
xHN1MOD2hqsbLKna9nY5WcP6HGUxfOD9FE4Z8V6l32zaTQxurxXd1+CCV0/x
Zw0I9Fci7wBmMqSpCuNvW/3A6VmlrooeLQoEg9Yi3ATYio/soSJRKABnH3wb
njeVGo29s4suVXSOYHohjhuGHCnvAZXP/qigrv7rT3Gu0ZIkKTo2hVyLnW0Z
D8nR0z9sJconoGFrKc8d2VhtcUHJMvn1d+tBmP0eESAsbTxvOW6P7MiD/vIR
uO9JVxQD8gx708vUmsJ/dWZgaopN235SUXuyBYADj4JVAoC/aHb4n10/iWCW
onz6HyD6Vc5I1pQoaqjlQqFx+oJhGzmSz8fQFFWKNDgUgL14AQa3rxWW4y/5
7JMW+IBIkNLPdPCQxYKsWkspHgU6CJK6z4D4PBy6JVjwJSFKAqofKjCjnquH
kUzkPi5cwERiwkpbxUFYmb2bB1r4z6KCd6xy4LNpjxY77QCb1TF/qreoqq2J
T8jQY7peeqht4Fc8DLFLUGhj02RGXJl5RyKsQ2lNMze8UxYqSLTyEP2R5XHn
oQ4Zwhk9Uwz4z11hAGA6iFLDTVdTZ/+VKN6C2Qfu3qJC+hiY1sOSQDp+gNP4
0x3jJ44ryKXzZsPhBw1gR/mEGsWnHzG8+cmg4u/jWBYQERWii/ccDsccyL8Y
Ib1Esn+/fOSWdruZXJjbPQ6qhc2YYLQ1rk4c11bamraISpQ0/dghD+cRuVsN
pkkJMP7mImaKHcw7apxCL+t0ZAoV71vT5dwgduNF2Jx5EHXhQwinvlbDRxE8
EFVbsZ+HmI3Kk3xKMnoImSBc44X7DdX4ZgLZ6XnygXx3GNbNCSNtj2zirFRM
rGsJPjGAs8gr7JDNQYt2Xw+lK0ZxORplY73gbWvgPB3eUEY0E6ZcnjvKLqx7
MO+zl0tdTm59AAK2sW10S7JLE5ItyxFWwb0pIclmlhOj6yAKWkMxJur4Zmwa
xVpwIQbL02aeti4X4oLHMAysA9yKGqZkDnRL1L6KEVUZY73KmP5MKdCzeJdM
L7JYjVN5OSLiXBehGcsl3Tg/nK/iDO9dj59JAoQhnPuLk2fTFDK2m3r6ISmg
P3/2HmRNDNxqCElLSty663JEZiPdilN0jBwY/rSU3We3uh3Q/Hlj8PLCg7P5
ZW7a5cVW5dh3fWe4qQ67Ltkm6i3H1IU1p7zDt91bVmGHlySh5qU/5lmKTYI4
ug0y5eA/ELDcY4E6QKuckWtDu4e/rU9Tie2D5hmWOQBrFRqA68x6S75WePe0
dCvpcmdQjSnnM8EN3qEHQUz6EglzqTQE24+6f7pO0T2VrULANxWyxSW4/0+I
5JkVEcaT5RRydlvvRUUSQZ5F7qi26ydYpg8ZC3sqp96a+XoNKaU29MzBRMH5
RVXSTCJ/tllmVEKhiLto2Z9l3o3OYdpZq/EMudoAFQm1Km6dCTfF3VPprqlb
8zGNERV3TY4NjwaFZk5ZvVR+j3gSumwfrzkIDTgPMd19FSrV7d87OaaYUEqq
5DAig7OW9yX6Kqa0GtyFhqhhkO7uuimap67+zNtm7cdRmB52Z7fBCPBLf0Ih
kStmZQVpzOjryXIq6EX7UpZmB0MqAEednoUuXJK4owJxhC6p5j2y9QQYWqgB
9nJggdCpBokD8Bt0cgu7QqS/uyhrRIXvwZeErE6i6vlSxNXvZRCnZvtCO0Zo
MVqps8Bks/2w6OBumqEpn6uv3AoG1STfWSjdFO2v77hOWQ+MP4zgEK2B5KbZ
YgHDd1R8W8Rw4B07LZCOGpdIyFacZ4dY4hW6Mu6Zc0IpoGH0

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfZv4DmBX0LKtUA4k2fl6mOPvGc+Cb5V1Uq9JK9frKI9Qug4bgmeKyHTNFbLZwC1l+C6TxY0BZ4UMhHmwmdBLbAaXnQ8boxzNI5f75OKZzezAXli7MKvH/F8NcZT+O7iv18CHAWGlvZgEcGyd0fOAhHCadkud0BcoOPtsuQVffIJYjzXWkj/l2aN7gwkbvdl7vATTOJltXRVhjpDor9cG6lFv03m/5kh2PcM/jX5/NUuRR4uy50Ei7oZlX//s5aNJOJIpc3QIqZDIPvuNgaekc7qsSBiBjqOdKYmeFk8MxcmCCT6CgxFukMJRW8/esEB6tA8uRSvnef/bxMT5PP4rmi8JOpCSIYO55V9HI4i8nsZ83Okijbs4dgWtqMgg3EHc4lQgFLKbSW8d6B6sn916N3qrA7pr6Ht24TflcoReIghuYucFu4FPA6FT4V8WLkcDGfxFOF5DL9MsN44KXfRRklGFDNUpv68RftoTqVyhZHMlMxtWiH9GTunJe2brAve+yi8k/yGrSQoakKUt/SERObR/bCMLWedghoxBRzf59g7qpffOYamdq1dAToSP64l6D0rdcATDZUMEYesfZw7DlFgl0yfLYf+Z/41i4g2hT69jQ7KeaPTRuEBO0T5+XnNzo2doQBNw6JKsdY2IToeZ1LcZh/4M+Ao+fpXN213oYJ08ExOpbePahi7ofXbULp9s7vgQVgsJNTSOkefF6fBXmoIZYJgxhkZ1W6m7vQRHUZdkbYY/sOliylTQfkAT6fKN/L33PIEYalz7DmwzhYnpWP"
`endif