// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UXW7ISdliM57L7s0F0QzldABFyYFnCSEFKRKkPl9Kgm5740EKxEivRPNGU+T
l7JHJq2NUhSbYAjpv8UklHOv+OiA9lhEKWM+UnppnN3jXe0hr8GyPfwAlJJG
lKmfaDYTK0nbQ4YijrEaF3NNfJ5cAQCcTn694t99akwjaTxL6byN44j2hU4e
qwFoage/soOpJpl00W5BUEfMc7+zocebXtZntSjC5En/Sn8iU4a6U9fIvE0Z
8BY0Jq6oEYcOcaWwFCGVyUkzMC/h2nOmGQI3wleVlkcZcgJCuBFQRdO6y1np
jPaV7pJPSlA+y6/aNeJudyiqJF62xHyzvks4TCKMyg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AWhSUyEWFZ9YR8zcsLzdzh0SCRLFUoFO3nvT8OSJadBUr1+BILUoM4y0KtUW
+Crsow/BArCR4PG3+5/MumZ2wzqFidscE7f6wfr29sOBl4IGcSGe5Muwqko/
X8BP+dOnjjhTA59lla1sE++S1WFemkdixu9PpSwkfThvh1rl9iUcNRWh7HGC
2OiVsTUukqNj6E9VY/nSUAuXLWOFSoQfdUgOxvbjucHY4Fpmq1FXjjTZN7uB
tLut2kxDw0+bgBhox1iFGrch+ZjaVEBpoZW2bZWaEROF0YBXS/6D6tnZwzK+
/MqUSuJr8lO+Ise9qtMTibFMCLRpovIwKE3tOcYC6A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t0R/Wg3LrVvlgzoePLY9zIegzzxDP8hVdHY89HRDkOTfEDCIP49gRTWivjM8
xb9TSbXGbiKzCrp+dOE5KqJ1/dab7rHJH6XBqrJ0HFB9dgs1gdhPNLosmn34
usW/AEHtUQwsdzNYpVfs3dgjkio0izYK6A35DoGi3kj5SFuICH0OE8SennMe
K4pxuv7aSavfcv805HDRQsqAnIu09IcgNAyRnxbN2zMzoQsSK8ppP1Ofz0SD
9Ti4qvldC4nDOqXX0/ZZuWTni8igtVe5QQXT3ndRp/7EOWUZ09pn8nO4dlK7
UJN/bISWETIa+ZVzj6BUv8n+J9uErx1bcrsCsJXg/Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FsAzyRKw1/Zr6NIMkb+Jt1tnnNRLm4tbBk3ddZeymB0vNZMEyTD+pGKdrLYf
OMq07VVng2ynK5katvrDTwUBq1hpS0OTpiUKjHSZRrGPHGC5Vwz/w6tut+0i
+UANUtfaAf6yRNrnzwBTj5eBz9AHU4+YZVTYh+ja+VEI3Qw7gVWk8lxnwoJs
WVt/AGo3WQDklHoQNbhe/w5C/WW2zzMnYjMHAdpziBvm2bZN+lvsMvG3UKzJ
0V/QObOsVi9HQbg9VoHmn//EA+KNOrIujrbpYaJ1IHGNpt6N9IwycORgGa94
u0oy6/WfdjteF2Vjd4pzfkNj6Pu/rQdQVyWhNdixjA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fBv+H6a+uQPoi/D0G5y/E8phi/I3o4L4jLkGAUiv85KZm4jnZZT63qgY+HQ9
kQVJV/Fed+meiyALtPucYJViGgySG5mcby0QlwwEOjeDe9LlnQA5NWn9E4nR
pYnWkKTAtsRQNLWbM+imGz6Q8pQyCO4l5LlZx8qK8xCCKCep5Sc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rVydJFz2dJ9qvPJluqLRBQs71Y5NGCXDznN7qXEkoYFBmn4vuWQhx6rHWR+W
LJF91q5vkZC6tBtksT2b1wEbHVt77D1QYYqlSYBf7h4pNoH+gPlY5X8OyTLw
aJ2q6ZyaT0A26OpjIVdzhJ94J88R9p5oCBvj6gN8VvC5/4LofJ2cYpaINk+L
ceq34HMvaKzH9CeP9THmBxDFe8iwN/W8+mR8obQVE7aMuyiybN/dGpCe+iYU
wwrbzKuYzpzTHiLwmoM3cnvrQPGMl8bjukvGGOP/mYNGtXp2Q5e6ijitXNxf
j0ICdNpRz/6a0ZPbpP/wCtnImsmtqn6U0gc1AV4mAbAHqGT13G8RswY5q2dX
7ICosdsWDu5qW9d3ZwQuhP3DVBn98eY5JxK1+YOSvcmAZUzkDsWr7Zxtzs1F
lmrcLudjLYYfj/B4yIhFkwxZBPPEE/b+iy8MoA5DfvSxYkJZ5yC3BlR0n45b
7bprUzA3ohM4n5abr2kHCYXZm08nIpr2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iXDWI9OZ/CQbh+cXf6sXka3hwXUa6MvsszoLRPNn9QnHO8ApQD2WSXAJX5id
cp2woF/R00Aw0AmteEqDMfk6ommNSD6j9jvNBFRMZVNOcy6mo3PkLq9DAUIP
UePH2v1LQ17+ZdadZd/PyXo4yDvVIaezAbfINfoBC/VonncoNsM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z+P2aHQXsbNLdHmKCETCjTTNeYvYkJ/ch5LoWDC9PQiMK50bnWYnCWVqsR8G
3DbuTXHvA23MyyBcmvaCb4lJQq0n8jqjndw7CsOziGsNhAYlfe3ZNsquw18d
5OZcIJSyox6dcH4Oh4m6XKW8FQWoQkRYKnZgmJZ3NxM2ubJ0psI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31632)
`pragma protect data_block
FZcqwdlRM2h9D/dnDL0QT8Y6jyVVk4EExzQoGz2EMCm8B4YI/23+XVXYryrZ
Fj2X6tx6olbqS4d93SZsOhzb7JCl4Gbyr21sMZCW5jmKqst1+Jv2AXS+Pt+m
2ez5VqEIZAjCuAanfhELVfAvw499Jr9n8I/aVCltPWG3kFdBRZAewab+r6OQ
PJd7QVpq6yYmv5aOeM9Hm+5o0+4LBRxwDmavfgWyuov8LCn7AGWqL4xMWzzf
HcwwGvDmVMmEJGYTJaRJ7TwU1Za6WMUBCtgltRCf0VX5DBzq6pYqMX8RRy6U
4YCnUE/h8HwvH5VFKeXd2fiGDrtTQseELaL/uIq3Q41cSy6gHNQrvEXpRwMN
N7g41Oi/hbOaPKkLd9I32Kms/GHGpt1u888AvYOKLRkMNAY8o0nyAprLQdUv
fEGowVqBOYm6DQx9wZ0PIY/I3W0eczz/qY8ygA1gMncdcVaXfy8Syb8gqWQD
ticfDXFCcgt783h3wcYeVG32IdvUcT3zdDrnfdAWvLPbOjxNM6QWDrpcULDF
A7J0gz+PONBIdMbVO6O74Iewf2r0r1qSAuFVn6EpKGXzuGWFfLx2jG2gLC5J
9Md7ohzt45jpZCVuPZxaeYp0x5UBs8SZFs+7gtzGNwnr0xrRefwCpagPKljq
ULyjxxyZiKaKCbiT3PqhS9DDO0hawCANUP2gVK/m6/xLuSH9yEN83hM4gXHV
mnut4pAGyFGEeZG4vVnIAxaWC/e4FUwN1ciH7d7HUxBIohhxt8RhrW0E+BSa
6/U1HfHEX+0uNSVEynZB1aG8IqptrkkkL65zAFRjloYvwRbLXEWDXbXjlwHk
wjE7krTvFtZ5DkZAjTEp28C66ZYY/fceNcNbiMy/r1PCu70cZNQzg5B0wfBe
F7TbendfZ40Gx594KkGPf186PDtJN4TDZuElgMx1f856gHGEfv/BjxpXTXk5
qmmnIFIWM82b2myJ1kZIvKlANqRRLblkRjzTlyQgB+4NovmSHmQYVV/jq4ey
jKwACDbRNdpDU7BaWK3UAECYib5mXHgGtweHMuDlJURBUs359+GpJhHbcyhJ
DHUnwJruR0LI28SOEJe2RrBwsU1jAPVZAl3VqCEfZ3D/JKYYGvxAWqgRJeoM
T7t4N6CqcohTLT9NHf5G96kd7uQPKq211sWTR6ub+A0ReCgUyvdEC60KGvIb
+NhC6snmPrP6/lfd4LJ0yrthfEJKoru0OSHyg46zIORoBSo5O3y9FcYwqVNN
o0rW401XTwoS2IMXrcZaM8EFgz5uQa87uwVTWEkKmdOI/63a3VkbQVYWylgc
ueDCPfkXcvLSR2gNEG5/FRe/4U4F7qmz1YX7XgSzIfKFVe1Nh8FvbXzZAtxW
qh7wBceMC90vY+yT5mSrGlNhr58d48I2rY4LWZTbOS9HvQqg6KWv9RNlOUQT
jruv+Inqxeur/Uk/JN+m/wgfTq9BYu2DymX1/PCl03eakyYY6YES5h/jq5fS
zSIuQJNqDoC7nxe+kU9UXrJXDf4u6qi+J645FmAsygmnhfAsSqvVUE0RsVnK
fb1dPMURuYS2pCTF0SgQMHsvCoU7UlOSDPzNoqADw4FQbwClwbNu5Ex3tBI2
6kEXO41Mt9hSe8onBlkXq7AIoz6/0cLGn/RqjcoNwJgvncqJk69qBxyiqpRq
/leY384gUbRdNbJQGErAgbbZ8D67orHvTtEJk3Yl4r3IVaKk+uTFRSrhbAr9
PBNhRjtSjkuQKwxOLCtL6Qmuk4LaHDrgFnUGs5iYGUX9sL6NOTPxoTMwSKDU
bHdVIfsN2Z/igHYZ+woBhpsckytnXN18XJnxX1nUtCAWUC0iajD4ghNRPmHM
g1n+j7NeVjO/Rd3UQkuzFf7UsmrFy1bSzNS1Sxw8+dJBHBADVEmzxclErae6
77XpaD3/uT9AOEuOnr7V37A/rQT7xGMAHHQc5CX4LEqSiuJ3MnKgu8ymcxrh
ySZdb8B5z4Nx4lCFu+Y5XsTekwBNJzuOrR3zMmu1v6Y4aYN5ZFxctTESh+EW
Yl4rS6RYvkkzDoVyK+074yT6rekDGkWrV6MsCXvuYHqa4drUvpC5RlotTJNL
S8HjzrhwkPo6zUvkyMpjnBdwjdITIcFRs6h7oV0Ayl2IOFwasSfISDN/AISc
tu9q/sZWexJmdSd8hwvRQ8vkd7zedy4XNHu6NN2ckum/o8T6psM3nk5ogh6W
LxHmTpQKd64v9ZTzf2w2k8ybe9+soowGz07AYsW766itYKGkkNKLw/m9bfiL
OO6nWOR35Y2YllfbBlgfwEQx4fYXY22/C2IRkL7VJC96DL4aJekX7550+xVN
DBAlN8Yx3PskvTs2TmmcvL0osaO0TYK6XQmi94lJ6U6oAyjtb90RjZLvYAsY
kBou8Qla9jTyPMOcqealUYYJl+XHrBtl7Pq4yZpOupPqE8CEq9T0QqeJZ0GH
Ph/498glztI8WbP55QBD5Tatpo7vAikln7Hp0FqUYdSqvNahpbh1rYZPj5WD
SV04Ub/34CRRA0/5oKh6agNZ8deri4Fnb7Fbpf5ZiW4H90sVTaDMdGDVG67u
xBxSt8j9u/Cs0KtKPXV1+hpbNN72AkjF+bn7GFlbOzX2OgddlMWXEo1ZfZMI
AvbBBJt74mhhVn+W6BcHAVei18aOafDeY0sO8xHbznOu0x7K2/B/5YaMYoUd
gFBrXAa5zUGV/Yp9kP7SeKodVy7YGEl0Hoxvr//4qeAHMlp1SvIpKKA5qI0o
IYb7Lkixwaoo7qRMWSwU4n2U04AFWIPULGBr7gKiTj1nM0QDRj55HIAlsYRD
cv7WZ3qnznL/fts2hGPgfcDDgUb/GiAurAcosgIEk3NarF4ad1ODM0mneLb6
CkXducnSsGFGMA9aK/wmtif6TNYJfCWxUmERP89VsmgrbDsdVlDda6wUj+Sn
Z/tBAn+9mEFQXRjSJcRsHyJjLCR8EOgzzxBU/mSxGdbdEhOimaUOq+poHbfK
nrEb5gZNcyAmM8LvsFKmHtcvmL4zBWES0zbpeH+br4gwRczPKm+OybJ74qNL
xXdsJThFThAxGaaIfwhvi/ohkziLCGwKc8lIeQR8GnkOhexpfdUI2GpwnlB4
CFFI9dYXqP3wZNPKzxGpv9VaLzrpMZ1N2Qk1XtGPQSXdag7N8/uigS+9NEFv
F2jaN4akA9CJsbCnMkAAWNEJwfDZ6Rf84NZC/UVhUpo8++SLye03j6kxhrh3
HG0SbfxHTKTaPKDBeG6x6SA/ZjXNWeZyMN5TxYlRcTvWGgnLgE7WmvmY+Pbx
mbtNCRunVF7+CY8ySgKEl9te+7I33k8X5F5nHl+UQpu0ckzomvUkxHpNGJeN
RmwqvKlw5VIIwaBNa02ULx7IzfTh5riYNrBkY13YgpINbyEibXtabUrGDOsM
tO4nRbYMIyE1f3e2tOVlh0HPkbd3+fRVYWRKeS9FrYiEtH0dDInWaTup+ayP
ANeW/fyItYgpZL+dafq8EcasCHMt2vE+J/aUqdDy8QQwdGymKt9dvsYW2Iel
hWUwCtwVrxLINbqeGTpXG6ktrjyaao+gs1I8/w+6/1fuyMFyVw5yr4VwBUIq
ctg9RxYuSvI5ObOgQPbTr9YVJY210PgrhqTaC+Y/pgyYT+mlkXVR7/LYib9L
C962I+Yygxuaj65K9RyKHiWgK3dyuAuDMx37b4z2XwgrG1qoeAcnv1MqqNUN
CEi51Am1Vr4edN+ckFiQiW21wd3+piKyjgCnzBnz5THFdHQYqobLH54jB9lq
Rx9NFj4ASYX2tUGMauL8QPIlQb2Iav2j8N1Mffw7XXEuq5fgaefBizwGloMY
M9MGH8Hgr7UktVS2Dbc41qMnTTrpm4vWaqZR9bIp0+jbLxaLUPBL9GumlimC
2lMejS+ELO+A7jAEx1gJSgaSKcIHSDMuCrR2CZCG7qz3Ek5NnaDqggqEWLfR
2p8UZw1JIhq9tc3iy8xe91VfNYBCTLbt3eTW1zIGXmqLw5tJKZ7pSWmZ9Xmt
0TPs6bk7b4fwcs0qOE/Hna6DVxJH4jyQikjFxME+u3TmscgycN4OP2CddLRT
Cuh+LaQJ0rbloiuivkZAfs/UBl+IfIWUkWF0nQeO3dbysuXRbcDlf6TneZjg
5LNDmF5L6GeZP2zwQFxVGcoq23Yu2QRt+nKu/GtPSnYThPJQQ/DxAMa8Ol+V
zpV/jSL/4BF2j6WW5HcUq5ZKkUZkUXn4zhXAfd0vn5VIIvFQY8L2EfSdnhvs
ZyAzIKVUp0u6sAahGZ+5fPERLnMwVpfgduSmAasPVlph6si/BrQDRTkH6Wp2
0/Z+7D4KpaxlKcaose+pgxiHeeBuYVd7hHYoYjUg4w7zOABrpzkRF8wUd0AB
FCZXNbnbHY03aC/Qxw8eeAkVA6rEymeSXlz1UJMPwUrVMz7s+ei1pP8tkPTE
bQIaAM6N0NTaDv30Q25WFLqFM4GGiHSVPB3uVWQeLF05AAaXWibVybd8MB+r
ArPDRg9O40uyYYMgy5Y6oNsY9d//Q8XF43bqqHDG4mNbyZQuwoiOxo7bXRSf
pa0ArS3yElbLfq6/kDFY64wSQy7k7udGLjGKTUpTIbcgHBdBq39TjR7xm2jS
yxOyXzjBTnIuuYdCJ+h9PSGcw5El59RrG8vOo3NITkrFY60Ke4koH5rqIA8p
x55ruz+26wrg4y7HwfycEwBcTq4nZnEX8ozLPTV3xtSgs0PszKYo1EVoMS4q
rV1OkSF+cgQ2W8I17j6hFDK1UM9Z90GAf730cjeVhxVLqwidPOZKLIt7s5+y
w1E/9AgL2/33LMHWMXL9xKAJZNFBzBE24fc2g45ovyKyOLsYuPgMGw07+s56
7rIckRMKyuGPwHBi9nnEaRgA9t1kD/1kh9mcyIJ6HF/nMcAM6IaFk12VP+D9
bGUP8G1bMGot49xhDOw3SfOHkNHDu6Uhvb2XiEt1h+TZ7AWMgA/uR9wK5tiL
zLbkNIhfwlhwQ044nhFIXgkePTIo1Jrnd5LTDbQJss6pp5NNzOu2VD+LdLlj
v+5W8z4b28KFVGsE3xk2LVh61tzO3HA2XtHCIEpdrYa3eoDEhiHFsEfUvX7O
Ep1fotEf0sovnjyMyOgIzSOGukTHuUMbpGoWtjHfm1tN4qirf5qhg0n0kZC1
+uzcfsd9sp2i0bJHOQrLpoFGIaSxpG0tiTicYttsjr772J4NiOFOoinOYxnc
EffUIj5vxWFg8p+6nvXGZ/rFVHiIUzyno0Wd23a7rcgU3YUeLvhBR9/6wTHy
+Fv2jOmlLlPjVn03YK9JzS5LkSQd+JEGjiu7V0VrAc1bT67hKOuxA0y+s0aR
CtUW0fD3dNRHxPl1oMFMJMzyhRoiB4pdR95xuVayRzqgrBhsB5x/7hxMSSge
IfME6ePvjpUifn07BCUDxXTpPALVYcDbooAzdNB27/iqaydKwvdRH+3j4arS
VkxtODh1xy5YQCjTa1FvPFRyvSxlBj2nyqC7CMYLo/WXkdvIyO+bCqSaO9FC
fgmi0qW4epNlgib9sd3U7uROlPbk+8CORj9U+81OCSG0BQenByfTN8CKCVhT
6APo1+eSYwiotWN+E95uH5y4Vsd+FsQ2PXrN2gGv3PnjAFPoP0d1Q4NLvu0R
iYLeL+8unQWJ+QaNXNYKpTAXApcLgCylH3Ne0DVnRda5fi9xUNW/WmmPli1a
fFYEcRlV5TUVm/oxBh5jo4JxXCL78DM1D5DJDKpLf27xvUiCjdTgPmWhW6dB
JU0RCZYruw3OCJKaXQEgXz+bgRIfb+d72kw3CoXpiBDMuRaC87TeVZR8guPA
eyfwRE0UBm+8J8SubnjSWMUN7VVU6qqtSXM2dNh1HFHES2yuM9FQqhFHIAZx
yhEnti6PEmNAtpL2Y/EmVbHUNaTpPwS5ICn0cpP9os2tx0pdwR8Tt6OWH5i1
YYHYv0cESpIoOfGDPpJccGuFQM/UnO5dljlAwe+kpQOiWoKn/zrHzKtP45QW
4NYI0lqbLLkIlTcbLDPtDNqXbYXOUqxpD8Ce551dcx/vuHVlGHlCiBTv0hRi
2uck6vp6V+ktPJ8Uv/WYiAC8TQpmlk0D7mKjDXPgdTECs+wZStPIc+tG5/G3
BgQ3Y8sS0ep73P/C9ia8VtOK3AjuQTCA3PTV3gHO+pHDbnrdaKn9DtXixU7v
xfNpsSrc+/wRnZEZIvrpfHljqOPHeGvbc46+Pqp3kI3uvvV40u5CS2jZ+wJE
JBzlBI2FXxn/WDvj3PViS9swYlrdJruO29425NI2BefRszn54W0QrR4kKj4S
m9BhaPgfH0Q/rv91+8/VHy6R0YkWebBajtzAuG5C/lWVlrXVPk5DX6FQNwls
wcxonZRuq7AbvFC1Kh+2AkS4G2FzM/DsSqVUQaCo9dz+x9o/Ij0/7pYtb6f/
bzo4hUJIfSoEZHHzLrbkH/V9SsFjDzqgplOg9c04AzNiwZElIfTyUBeJ6fkg
2tprRnMa6IBYD6bzZWXmWbVW16AwESa7yAELR0Qzp3VOigeUdCFaIih4jld+
5MO4igLX7HaLzXa2hA3ZojgRbF2+sZagULEwmabKQPav02AQbjCDYegDYNly
wotb+XvV6kaVRaL/yQhpe62dlDgBDd8QshZkCV7kzbq3IIe/eOr5KT5k3DN0
et+QGJjVSIq9jTqWKZp3X3I3jEFav21oakXh+sxc/SioMVF80a3Y+5dWS4AE
NXBZdLr3luN4KlHJokx6ssfLfV5c7X5d1U9egy1LsRLDFSEbchmdRII2HzCQ
qQcQl55WYQvOwylT2TxZUENphsI/qq9OxkkrOUnFa6kq/8vhiTa1MvI24qAQ
NgWmN08IGe/UszA6F48gVHGM8ZNlMbW+8tYxy5EbSweAjZa7+wQfDEV9mSKg
BI0Qkwz5t62+bPdIEppevHPwGEbMA5jyVJ1tpe7DGz2BBoq7nRQVQ+Oqt/RX
h+6AqdSlVHNzgvhECe4H8UZIRLoat1tIyXHeeCUsfxppqLC+N8qFUtPgqWUl
VhWXR48Vkx30jS+VNwKbZTGaNbKXvs49/V8PKDcINSQl2i7wh+1+xMK3p8zA
oSs2d1z+QJ7L4wwFVqw/bpZ5usKjvcpSKlg8fulzWMErKXvMsCJ5onlWRG+X
2Quf+l0jgE9MZtSjBdm92ucF/pXBTJCDCmcgWZms/AcdrvWnLfWRJnYT0ZMo
13b0Hqs9E/krqMdRtQrfDiffpPTk0GoRQrQBSKYJKytziQpqP6AxcoSH/A8g
E/0klNdBuBBefZu9sZy03ijzPBnyweRBrg3sQbqDSyj7f735ax2f9ZG1hdCH
HafRnBsEFEvrWECc1NcqDQYA+8oYk7iCKWjKVk40udu6MAJ7eIajhl66FVcY
eAYoZRbJXB1gJktP6M5mEQTccBpEoQW4uNRMlMlkjGaoqZRrTeQ23lh79Ey5
UC90gVlOxpbvE4iUBRJebXsdi/LI2NgnJABcDntMu07U434HnyGFhKIbVW6P
4cy3sNhqwKxnW4CU+aMdZstPyB7Ub/8K1Aujg9ZhGzm9ERPSZLvigm3QnUS3
OP2I/sUCa3vHw76/NpvpL942bi2wm/nkVlW8Mjq3dHMgnF55bxvRO84+IYAj
dIXGkfo8X3bHsts2+H3iICHjAo5UDOjjalsLIFoQ9+8B/GdM4Olg4O+mzXT+
KHJzF3obvxZOnPDTPFO/JEdI7IBjn4JngVcSw9mNtWqVjqiZKRFABkoWvmfT
JvqsP5saDev3mT+AXHT7W18FPkYRgz6qnPl2xoL3l08Fd52/5N95/HVq2DF1
3Z6kyajJefo8JKBWFvm3DxcNImCZU2j2uUY3EJpDS+x1Y3G86vjHVa6NHAaI
82VR4gY9rqAmJ7Zm87D5VKVF6eRr02dTeYNNl8dl60sJ30ct2mgv7E754jAD
zc8fbOnlg89bB6H3B0srdZ82kbdknEpWVfn7dZM3oA1mv2T45hrT8DSjZGV8
SG3xgOPvwVZ6tp8+8w0jzRPybisiZrdGefIB21IVf+RVSIvuuCPAfYSrf5nd
uXvlmpXyKo3G1OAuZieeAehMSNnKYnwyNmIi6d8/a66P2UlxenhFp3+xxmk/
vMetcaikYhaCd87ZVqfe2LtDETcv+zzKbAd905SfjwBXacQtC0Fbx/A9TfDE
w24NyOicKnYab5ESvmOvxUpQbuItk9SRi1VxGyEdExMbyXMOsgaeyBy3mMMe
n7O7j7Iiq84zTr4fl1bP6F+au4nNFVWehsODyhpTwfLRjrv+SUg+Faer3XVG
QyzvlDmHIX1Ahafty721+dmc95VjFB+WlJk2KXLghYusJn16hsvYiG1tyDQ2
CGXH85ZiUKi55MyjBIuYZKYLP7TCaNF/zi6TcKhbssDTtg1w/xVLZ6lpqX1H
Ih817WNNV8i9UWLyqlqQq7MxKZohqOjQFYSiEAUuvyICArUCtrjj3upMNyup
0xzt9c3VP9Vd3QQSaZ5L6gPySvjcOz3iLD8ja8rxz5q+aLj0c2wSJug6LMJl
o75VG0SrpYynqsqTSY4RdPVniDnVWCft5BZMO9CxU9BBGXU0YyOEHrAqYdsQ
hvL6wl0TIn7occXcP0P84vsU/KrL0puZ6X8l1JHpxuyK/b1p5ydDr9zQmlBE
EYkQGPvQGGBLmNk7w+9Yh6Z2IyOuj25rCvdGn2A3iX6WzRyGR9vaUd+Nufdi
KjJ2Y1g40Zvti4llouN87dTAdir2L9Kv1Jb2clmJHn8po3S3T9hINrYNnkyO
NsTkP546p7TMCGiF9he9XQB5uxamLz+SaRnnMbUCl84J9LNQyH2nI5re2nuF
LA4hSgsZhiRS2GBHy4pnZ5TwA2CHyi+ocPlKd4DlRaBdVB0zERNMHR0pbNLp
ocvYm3is0KtHisILvnXNVGoyyr5dvyIND5vFMTrMEsstbjOZYrfDC+DMXvu8
8jqOpdpmyw2kyWTXpbKwowqRTuQwrZYSiA5lm4ScKfjnDLauH6J9QIJA4LcK
bzTQo5UQx5E0uAB3HMdyk3PoGTX8oxvQK1er/f1ausPpy1WD0n14kZLn4hbG
TsP7muonHgiuVYxbZvMJxJF896IYdfHrY0p4IsyTh4Yzebm8GWiexxFxepiR
awGwsAQ5sIS2p2+a86W6jJfceSoHizKte6HkVC+2Rmn3dd0tlffRZpHS3Ahz
w7eedn5Yup1O2dUrX+4v+FuNjHGxLpXrfYKhv6qnNwfJPvCBtTTuQU9dAAC0
eMBz9aWXCFYZY/VTj6Ie1ab16/Xsg3edv+2wuf80owb7aoFPWSdRMQXvjF9q
VMG04L1Ovp80fr+1fzkjiI7DNsy34sx50R5p3Afq7Jh972Ovs4PDCEZwBHHl
OAplzWtvzt6XZwZ2Ime+9QqWVqGTaTolFYsvnHl7IBdE1ArRUs/6XN/lpvSV
b4ST3LBL2Qa6B8JvIxQRbnnqqRoqjORu08NRgVap+gcEIaoEe8cHj3hM+eoi
pQpdVTMwfHW/wJiX7h4clk0hap28ZqmIbAQGSs2Plu9DhV8PEnhU0ZIhZcMv
2IHtaSMF/5BTM3H3+TV74sD3m9FveZVvB638kPNU83BtLwcNF8wRcpmxKGry
ZgTdIEVhJ+T8O1uqhKNP34Ndf9Oq1OiwbFFiCdP1qYa8C+PUx6KONpagxl6y
Ze4AFzVk87NvmWMEJRRkCC4mD9ldsxObjmvmOCnR4wfMYNRbhPWsxmbzoBW4
pQ1OD9ONCCXhwAMKwD4mDSGFXzcm2IA11L2WITsbF0iUPBp7boT52C7LD/n8
LDLxofgh7/nElSVr5wDmpKXIumgsQTw4tB+sllfIeuuMAF5dUmJdehwrbHIC
d0mmenqSan2B0E9WT52F9WacuXGpnYfBJ6niKuBpVKsqvw8XN/+vw1fRlIc7
Z2Ihq+LzqzJExgH7aS8ar9OKO8kKfvlGukOA2C3BUE+LTB9/zlmdgyX7/jth
zT77hfbNblwXDJChLdmlP/lS98jYqpFVqge0VAEOV5BpA24a6fFpvCpwYXnf
/VseEOxnryABZvjV8dG1QhdGUynxgiBEIzYgh7YO+fBIzI70NMonUxqA0Gzm
nzMgw+Lp+e8BkatO1MGSn44BWNTrV/mc28NBSSEi2vDt56phShXrzKFIWmvl
RvRw41PXuef7pxZf0Ec0aKNpF97IZ55Kt3O8AqhTVAAxRu954SJ8VLYNG96r
OOMg6U9kakXYJnN/8tkgo64NcutsYvM/IsTuvLz21B5FMzUIdwqC2MZEeQrb
eVdfjhAG2WFCUs0XYZCWqUpRTKYX53r9hb5FC1uVUhKUvn4OnRHbjp43Dl7y
KjbaJaOXAgDIuYsAX0/uxvIDVp3pdv+pI/aTnaB2zeI4Jev5cRkVI8dYoclP
6b7ZmBMGCuc7+T8NP3GrqtNmNb/7tYTOKhfSWyC9LrkFzwVLUSoRRNI4Dd1S
ab8AqHrmk5R78VfQ5Oj1xsZLDgYuFB4uxZ4+liD1IvkuRPdTQ5G994WVAkfE
hqiGGD6hNWLo4R63lr/vnsQwMXJiWriyQE/L5UgGeYzHqZF9BME2VUKiFH5I
LzdTcCQkuZj26TnO3+he7wYY2qwc2g0GmKKhyG2/Ucu7u0WCl9jb+G+z5MCH
uht2kK+bn5lVuxBBG2MHnhv5ZYzFDgaZBi4ne2w6ltlij4/fSDLlILaaGhI3
trxsaArYwWwVvs+2xdTry+GalQLgnEW79AX+/AlLPwJ2tYeuLFZAEpMBeQhI
qHKIj4EpiZ9FwX4qrMYkr75kUEM1uaDmq3CqnQGZsWbL6RsZwj89/vL2f2Yw
ljliqzuwXZmfLZmxz/96wbqQWK3uwN1gmHwYsS5xwa1S9xZb9YLZadpk3LQz
dENv9/FPBE7b+W9cyn4/YXAuuNm+h+lUYNLJK5UOITYN5BbEt12cgm6KYJtD
6MpR9za8h6pAwXQ+HBmfzPXAkedCArP5TmLFojbkOuCWbqhVNqcCrRcAj93U
c4WoUMAeFHHNTbeYswPX5W8aM506ZVVG4gbrKceZChGk4YTfe1CtepWOimfl
y6YBIe1aDPJ/cNbBdrVMP9GW/hAMCmDabcVxiQVHjFkdebBb1GAV7fRJDrTI
B5K00qv4LXX2EEeAdO2jccnqLI/HbGhz4raJsQPQKCbCg/GNksfizRUZlazQ
VMi/KEqFt6IKHf0N/ez64VMlRzLsk2bP9+Pdbmo5RShtPD6Lyo81QCUpLnRf
wBfALKgGXjYtX8cFawI2EhllTK6QkrIwFJh9BpT+TqH7BoPRM7tUUeh3XRB7
8qfDrwRcnrMIM/ap7Tj1AlcUUvV8l7fCVd1c13wCpa8GYKTWmBYb9G1cTkG9
2KzlJ/EWjB12zcyw9zVXlTivvHkVIZp8FHzMgT1s43xKf8Iu0NXVyetB4rjl
s5g9F9dttumxrF6RGkOmjOiPeXmWHbHz2Q/CAqJCZdOOBiyIbeN/oPK5ZWiw
WpydHgdrJuLPiJLin/5YP1qjOawHxoKOHy/h9b6UHu+ns/0LWvWGXcsjaPWW
7IHyvMxy3Sug+YRxBuGMNCRwBNIRWfDTfaJhyQsBh92xE5D3fpwIMG3/EDpg
FK785Q/kAUyn+qnsPjOM9XtSytVtNKjF5Gvlw9XMjqbfKIwGLymnCXlBoAto
IEVfcgDJEevJVaHAfy0P+VaBmYVYsB6zWHOQcRI5+6K07GQNmBylbygMSTCG
f2waUj7jd8ipCgkrVYXHjxzyMH6LxTXVWQkCk6Tmz0uGSknD0tLmGnzk9+dY
OjfsaDOypgncbzDtGK5Ismvm99Ice3iEKiDe40BVTCNZRXtMT5cySw+Sl4c1
KEh8YdwfsyP0hsy4Zb92+u0OCziIMDGgTMRfRVEquKKhcxiKTaXksdASG/5L
0BFbd/GR7fJ8wa9gpCAJsrHcRk2ZS8NhWU7Kd+JrCtWgtNjpFJWVcGKxHFuC
2a1oe+WYYgri2qBQmVnk5dBeuAeEZq7/XDY1g52BhRvkVmltf6/Jo9oPcPjo
kOKNSfGQjWyO5S0+XWlEr0LR2lGx550JVy/g6TjVFlq7QN9BiL5FbZqDUzkZ
LMI/Kosp8iOG9HP0ld/dOgb1ad0vqt1hMhZOAleq1foaA6zFvYtTZsHUQAYh
zKM7sP8ku9Lm7jBrb57tMlYw2bhpE8V816SgdKZPr3yYjA/Jy2/Xw+16EPwX
G4bLcgr+I2v5ddwnciD7Ur7r9qnSOxF4SmgHOJGTNMjjfeDjl6jzMMcyy7Fo
OxFDSX8jI4BfjrlVxJdjDeV2NjsiG343babOrg825RITEb0H+nnWHEstIvDX
MX1QVCOREV8RaiYVvjSmsDcYYr61rxOCwOsC6U8bvynR8YQveLjyd0KEuQxQ
ZA18JVKfO5WQq/VXAX4ASVfOpTU1EeCD44wrsl/Nb2zExk2JgdV4okHTUPRp
+32WeQcIU0cKnU2IReisywvix1Rd3Cvn+Ge/NY0hKRG62DibF/rYU5x0E6vl
5iBvHJcZgvuSpbfWat2etXGBKu2DLqQ0jB72Gv4WxetN18zxyBR8bxurDjTq
O5rSvVwZwf8SJp8ylK8opZNCAw0nv5ZS5aLLf+2A6DftQr8zNq0NQ13C1Cc0
W1B3nikyLDE/wA93Zee6TXupWcbXiEsuGsJdtw1IFB62+hb8Dhn35O8qraM+
vZQziPr3KwtQUyFMFzZFLf6ndlnz2TnHhRI9gagjykS9oX2GG+P1o+6LhS2S
XyijbsL59s+S2aZf0EagOYKTEemEK4VUbv4itoZCJX5hXBSskeqkGL8wYUPq
gSVLwC1ZL3jJlCzrbOrxTRynM7TBevoKr+teNnqQufxxispxSx22liNL8dXO
EP1Xg1cHoFBRus2eYyoaJUeNgkilek3wT2n1AqISfDAXh2iqIBan1l4WdAJj
1uM8TRJ10jxhMh6bPcViZgDJdQ/1Bztyb0WYNrmBQV2qaLLikIT9kU7NOknq
fXVLIgBhyaFL+f85ClWPklpxzu3l8E25L5iJiXb3zyAyG96pcL9EK27QElbp
P1ZtkaMtd8dj5Sje9KgnEBLEa1ytWRsI+9AUPP5KLu9w7YEA0wxWVTTfnYbi
PiHNicaiFO83RAsmYdHQIYPZnbnFT73DN7Pf1Jgf3yVE220UYNJYF1BYdNCF
m6qBzCzcP95Lz8otQwu5DlFqb9BnwbOtXesDX3aP4JRjlZ/MxHCltr51/HU8
4SIApC9cmQ2I/HP9dOWA8OHi1FzDgfEyZTobyUfQk1PMwiu28sJVAarWlJBa
7go8dpkkVbvCQyoZuQMEQlSO5ZIW+56P0Qbd+1FSf0COlspjhFGo7GS9xyxG
V2TVMpXI38fCQAk9BwfPSUfRiAZrltd2/MEBLXIis5azGhXR1bUbl8P0Kgjq
OyVBOBO0UcMIvbxz4FeauFd0gFbpzSmgZIE0hQFmb0HxcrRCsd96UBa486uN
/mvGT1Q28H3okhpc3aEAEWPS/36NFNKORurnxNTwq9bbxCOi7+jXGZFP1UmE
fD64KsvImuxqctTqHx9d+2E+Q2sO/Q7WQL4YcpcmY2w7/smg9gpiZWGVwAvE
EvVFOth75s+to5mtnuWv8XNscLYk70oAMsvgWjKGw69Ot8bu8fd6WYCud4Z7
zKGJshE+gxfEjNQL1BoJRpkOzWTBero0Qg4mGC/fdtrZzigrUvbwCtzQISfE
Ph+6xdZKVrlXc24tM8CwfZn1oqO7UqrDQTknzAY8grx//4dyzHVH36rmnv+g
zQx6t+w1OLark8z/rc/EgJhXTKz7YELLPUOmJXlBh7D/1QfsOVQ37fhxd1I2
4sL20SH6S6wylRBMEJmjtpo+gJzOVyNKRN/JnQTfGA6ijHKxEJAWpolDtKYV
JYM/HqwWkZsl2GMtyljAzbg5UXaAvcNLX8G+xVLd76q7itg53WKRZsazth0l
sCWxSXMH/sUF2PL148SnBrQXLk6iQHqqc75C26uNEkrH61j+Zbxzq92Tck8g
L+Lmz1sENiKODWbIkFECTptPktoESATZqXTbjk64F7fMZQroF5DihE2jF47r
8FLjcgjrAFqZ6Iq1T0aZs8MCYXJylcCGOSHMXJiGVq5dVTPTURblgWdtfRmr
4MscYtzky47Ve7VuH/ftjxDcYW1Lckh2usR2LR1BYfVeFkhjwh1lxY1hPo4U
JbFDwRWOmaArwXFpKuHSVJL4nKhgnii3f3qzB3bgVdD00aa0MWkBduPMZY4v
Oy0uYCd+KkLw4WE8mTpvY8nYxWy5467MGauZDREzCKjHfLapNyxE7b607S0J
shyOhDomsgs2fqzgErt/mJjeAssKefgi7CE5v/2OW8g1+Xxh2xoP9eXkPng/
7ZLeML6u1md12TUe5EEDGZEnmH6cLdvbetnfPV5/gv87Er0ynTAUW2ZhXWW3
NZDAzLHjVNjiihSWBlThlLOipPoHEi+Q9vZbhEXupc53xymlquq311KqrQXX
CyPokdYotK1KDEJRQ9kyctuii1tXPexpxwxcc9uZl14j/k4OSfKK+yBCk0eE
0Yz8F+58AYDfJ8ix6OFCDLcCvvP6ND+ycSKHg3SUNCgdF5h+WzcX7WX35qYf
n8xWbDZGHJqLfSLEN2Om1/SRaDXHeHnSDU07gyJP55Ds4u8J/4X32XtIUKSI
j8QaSZjMaXHD1CDpUIH3ILEqK5dJgWWExuFuEOH7v/6teFqrEo4IzjehDMja
OAK5OkSlSgxDX/dz1WRLzcwxaNJLKOfE9Xrrl+3X4NE1yXdJZjrWrMIGG5Oz
opsM6RiSlykAhj0b+xU4Mf5TGHYReSzpnlpsXm6iL1BFmtQzYsnL+EBLAvNs
POr45Scxn4utxXXGMaDM5Sk3XRvk/2Hlvj/5PRYpwj1Bl1fXZUBggnUR7rh7
8fUAGoCclm/+aSREhJQIJ7K9z5FWGQYD176sixNxWveefBNR5cG/F6dwqZGU
3Jn93RBQuJ8kFByXkfJgzWevqnmLk999qie1YswWmA5YWyBI4r9nry2VDWEW
wxRKI3+/6vuUmRBHkXypRZxOckrgaLK7XSwu2BwSMdziwsukiP04XSm+ghG+
ka5vvZxWnz6NgAddZ6pIwEIt3h40pyNOLT4MR1i+7MQwh6s4s79E8i3Z7GGv
9diV6HnyExZfdQltvqFMwcVpSYmtTRQ95kkv3iuVKwW28Q3WF+a6dZk6ws8j
53bmu0rsorzbJsv+aiFORMto7760lRcc4kPFLmWOoG9tp+QXFrwd2EAsgWtF
lPq2rQG5goyoRqCtsODbFtvjThjxcCHkA+6NSAFxK+s67on+amLeCP2gAqne
knNJb+tUrzPKyAgQH01itZAPI3dF471Bqdw5L/Su5Y/AgI7rLz1iK1HgV0Ab
5yb7DzK+gXo8gyPL02XiAScpBUMPBb7KelvD/9gRJP2b4EEiSXQCKBM4CbRq
ZT5feI6Vt70nmTQ4kqv/BiTgEF7L9m0XC2pHktRN6i3M3cAga/gXK/qPk+O9
4wtgC0Qo+aqLOg2Rd6A5eTMcTXmfPS3mOqtLWktxBkjP+eSNJbNaDP0/xEsA
IGWetpwcxZIApsG3uwuiFAF6T3zzp6e70zR9hYyg6FJY3AIk2DeQW0h1DK3X
Yep+tx4h7Hv3mxG8AvODwNjVDJqF3NDmGdtGLp7CsZBduIBL/RjPCnNyvtZS
+zF/4Az57JJRRrD7wuPz1X7apDeQRIWUNK6Bwy5HK7xXNvkVL3gOtF5wRLLV
Oe3qUquFDEMaWzmWq07Hz836jPErVUEsI9UfkQK92sCR/W9fMb8zsZGENZ5+
Vk7+jMpa83hMxy3b1Y511An33ZTwQuYcLN1FQ4V849VXCansjSFBD9xLW+TM
Ht7ePLIFY35d35S9y3cZOh9T910vgLWbgIksIqtfuQfMKJstiTqgvW3uFGFq
gvYqVksmCCUnYKeUWNUxqiaD48hXvforoDRQlw2p4PPpp4xF3/s3y7JrF482
GeFmT1SSk9/VHF/CamJoUeaa0FSuUxw6BjEEnMjg4zlP7cIhH9zd3aVsY3bO
R8aSZZfQxX8/8AcWDJ3D6mwzv5vrm/oUyZz8oD0ZIW38yHYcgeBzKbf3PJAG
UvYC2TWGmG2o9IuFnM4AJ+XiIYF1S9A+gpFrR/HDmWCFDhWMW/xlYqvoD4OE
tQH5z3Ds2IDmt6WEgPbGQr3Rlbg3HoM/Sdqg9ihcAExfEW5hVNqbYUMAM37y
t2XE3h65QQvECyexue05rsdHXzyRP6T7HA5gHltYcqBb4WXeIe62JpEcp0+r
kbGu3WaVlpWU7lpK6oJ3p5vko1+utJapbHhTRk5+CUZ4zjgIsf10CJbZzuPd
XvGttyfoTaXQg3iE7G6RIiDwC6aArpQYrXPFjW53sM+kBw4CLuUfCkVZ+0dr
tm32e3dOT9O1yLTH0X1Huafm2XlWYd5LkItrcyvkiaMgVKaEaFVKV1nuspEJ
SUmaNL8ml00YiKmstvrKUH99CPqt5Zc18sm1NcAdDPGeXKi5UbQODRHHxPgk
n6ssyoMhxpKxQaN5bjOptpwgkBVzEN9+iK/LJFYZpM+Mxla4bOhSgu0EZmGm
Ilm6LiI3RFejfXqQzPSL/mZHNa6b/qEy8lMCZfLGu3aKObutWvK3nn6dYz3h
dy336HZ+8Tcjrj2de7FHUaXBiM+a2umga8AVc2zMg3SWXbO1tlZaed/bUve1
F/ohH47xHth/RafetyF8Gy+t5vYv57gY2CB030F+ppxHMVvFL16+UkDrR774
qxZ5K/gSM/9tIEgYoM76jJhB+pQ3LRVFjlkOSbVMGRX31l7yO6Z5HvkEhLOt
Go/5MQ4yB+osSiA0qPvqrtlj4lF902NfMQarl/y4zFjIyLXDW32u8vTELnOa
GDt2vr29x4C8ZTpL8l6CM8H4Hie8BDqLfBt3p/Nmm0h8FlX5fXziD5hz0iaN
DwvaFyGqJdBTqVern3mzsS1XbuiorcFZ2/GlUk9BGLE6cauFYO4Uu6ak8PHw
BS8+VkWDy32LUbBrnRulSgV52fh3y0CTePNQGOWm3MBZ6Lj+HTh+LcgZPlnH
zoBgPAxCjV3nWjuVLYR2VGoeg/WZMatXaHFQDJchhEHPX4U/2hz++3QWY2RX
whw+rkMGumDgpAUcFHLaLLIbIuY490d17NffS/zapmJtDPsQ7YgW0uZJjM1S
qkfKOyKPPdt7NBpYsvMWqkfSF+uNDoFw8/6PnnXADkQCmuARMMk9DLbhtRJh
Q4ga6Ojhms4uf4deJE9dV7ljX9MZoz75aIkQNuBPmFMlsJiTagbe/MqtP80e
Jsk/fkd6v7SuHXnbcqyX/5Y+GSyxyPRs+8Bxc7gIrVYcT8MBZwrPP38txs5w
Brl73tAUphDuhmTJJgqHNep1GWD2uM/J1YJ2cwJrYX9mQEsRX9N65dP8wEkP
YD1ddsLb9Zz7UmYf/LcIFohOWD+wfa/E06D2AmwsqJKK65dDUgkwFRI/vr60
qM4peS9Hh/9vPsQg9EtDKVehvkscLDYRfCpuCjQNj/E4PPjOMAW7JkuedHBc
JfDlHt62F8fjGPUQzOheu6hmeO1Jocbk0L/WmbUtrVG5LHYygFQIUe9Wu+sj
6tahoOsCE8bsv+xL827rfqy0rcrL9qiqEDyAnq3gWPxje7OENpzlEG1yB2le
4fF2MBeeOVCXB9Nuh4fjDwKu9JILj8zRMkofZH3eJYGsGfajlHvJHXeE7AFy
kQB1U1mXFoAJ7MEJjXXhLKNERD9pHaleWoy/m2IaXERHO10ofz4S0/qCLbnp
UBTtKMEHfo0NMy9v4PALmdvrqYyr+wxQdSIdMgnR4W2/0/Hx8Zkbz4wmtmz4
Bh/d5Ivluwz34ioVMm8KAptbLZPdERrzyH7dCC5c9kvsZHC/22fnaEnLmK6U
dOzPlwR2VfYFdnWhSGPUV79/79BOqDcPxAhVEpn1zO/AfyJAL23rEYaJvUyI
11UUVEeNFA43btcmXOK4GmVcluSqOc/mL6lp5S30na41Q4xE9ELk3oAFOoiR
gjQXkKqnIAKXx0Y7YrEdZwOaMuUGE87aVqi88DSlCC6xC0opnLNwvFGyVBlk
DXC6WmGmfEpGSJWDOnFh2OSyopTXyAXHgNYw09GpWyHl6flgIH/BRDFtFThs
txvoqmbuBLM2yPf4FTzd8gE2VUfZAvY13YwhkbbS1AN49DdoNw6bzWoEzgWS
9DXfk+PvL+j9YR+S7t1S9AInsX4NQVN3YGbq/175TQ7tKxBwLUn/ZVLZVjiR
jWni/UYLhdBEV8/lrvY5LNqg/46lQGLoLI2W03A570EvQQ6cRSqt5wMkRNzq
QVAUjgIsAwA6V3/HwdCuB60R9xWRKIcQMtWnVUfeVM2IcSasONR2TKHWoB93
MSEs+T90NUhiu3ApFTJdyd76BIb7UtewYkV8c9O4dNAZirDbYkiWaHF4kqC8
E8195wWYAOz4TrGmhSGQHMwVQZAzFaiecnZsiYu+qUhbhtMt6D2Jz4IJxVf6
RWhBbPETAJ9qYpZj98nbn4U0nQHHmJtTT2tzy+PldpM291zQl1HCH3giq9LI
t1+9XWyH0LA3b/5a4eyY0NDgDRulN64wQ0XtCWGdE3fydW7TXWEG3FFZpR1E
ABBCoEM5s32ItH7Q6QltL8wwznp/fftIeg18O38MmjeVz+LoDOVjzSWPxOcK
kMhe7I7waE2PUeEtkWsC3YgNyYoyn1GiH5LPF477e2uB5/ONbrLcztc11o1j
QjXxScIYeGHQJHvj3sECdy2yY0yd6h0nzfB2JaJybgpRRm0Oo8qkpFqVwA31
DjzvUdCvAbGDaiKbUHc//rmJaYjLQItKjS8m6W1XBsEPkB+4pZ+oYrsOo5WK
T0usNkWSXKtS+fgi2KALr8aXNvpOQKSh9223D5LO0ieFrpDYDMHc6Npej+bi
i4+o2ykDqmAg49rV3Ht4XABsGuV4kE1E0fUnBZI+FpLeuRQgpx1MdEtPXiKk
W+OLwfBfdZMbu+r630YBCH9BxMvKJIpgqPnGh5RC3SH/QjSHwPyrtLVSMTsE
W5FcfOIX44IRFGfQPd7rc0YuEAdpInkynU86FOqcrJqN1zaZ0Iod1+jGKBo6
OUyqiBLPnDqZ2NH9Ar1qlYx81MMHNm8b22uS9us/bUvgxKn8bsRC/VtLxeoh
8CLAg0NAg/70oF5TgIyipEhRVbRZZ6g9hdmOiW0xnOIdj1aNRllLLJ9eGMZI
/rfjF0dZysgGvoTH9xpVJSfz1eskYWico2gGFvkUtKID/TTRqgcwJEST863m
EgnkjqdDeNkQGMvKDc22SBvmd92vBgX8UHkVKHxKuAmqoukZfypfBpkmEOxG
51bqLVyVQqCIozzA4htyhvl0qdvtAULajtabq3MGQzxmKbroHuwO0fO4YsXL
kSgrpqNDR/wlazwP4sJ/Clz0UYug9aoMDHGScYu13XAhHE15yBUi4GJPDvdQ
Gj6gF/fsBjIJPQLZOZ+Ajc0Tag97ONLGlGOoyo/+Wqs3/mZlWDRmbk6s2ItE
z273jtT6msouR3wOWv56YjWUkXXxLYrFW15uxNVDhmCSyKs7VoQREtP9u7Uz
cIyZ04xJ/Cp4G1TKqF8kTZOhmejFtRGDU+C1j2zc8K34SxgLt9K2trFDLz82
Yoj3XD3YQDTm+oCnymMTk7tyoafqWgzqvoGBdtiqJF54xxkX7Y/o+q5s7UID
9/r8IB3DHDHBwF6KXDQDXwBVBOTmMVapXYNZfQO/kDdq3pRgYLItvsyeFJMD
fZjdP2u9Rxe83xGyvyEEk5sZcEpscF+IodNn3BTVP2jqQOEHDnL/JXuhTWvC
dgLcxLUdJfLJ/ygSz08vCsudvf2GWI2z8fbsjaWP+rh/vCxmZEC5QjAcKoga
BQ3LypdojHtAm9WctmWvfj/jAg5uFmSHI8PiVuL74QRYU95pYQqYon3KiS1s
oi/IRLaGljoyMa8y/Rz+OeD9pPygsLYfz5dK0UPMEq63BnDJjqgv6e2Ap5p2
ofK2t2mVcP6qRXNs3I84RfTxdjWUH2iKeGyKZhZA2y+gP3pCqOvLqls/cPzZ
3TcWX5jUgnMHhpwJpUFuuNHcph7FlRyqKZCSCQVDMI0rctTeT/qQuS2JRR0o
dDr3tRy/yS8vKhOA+h46q4ya969WGzbp5qarfKaVUnWjkVL9RI/wCGGzy1yr
B+8MwHHNrFD4rcu/38tpTYKCy1u3RWNm32LNI/NoGr/w5CblyRqimbSDHRzy
AXm6f97BZqR1coP1QWANG8UpKaF0Kf0WRnKR9JiNzVpPu2BUP113Qk+RuFuO
6NJXZ30dXbxTYrhBwoKZ0syn+yNCGm5qxKjRKjtv34tDn9ExtT5bgI5bKRCR
SYX+jGlEWKo6IrK43sPYp+Hj+Hg8UCwXp6unIGA5V8OokN4uBVOpf4Nq0OyM
JzJF37O6h2VFNBQo11yQIUNZ1GOV3LNg/fZvNor8Gs+lX+SsxZtZo2AtdcvI
KO0eNEHue4t9pYvdbx9osp3i/rX8vINofF6BLb/H0Ufdc7fIEXGnhSZbayn8
/CqwnzcoHHWEzodzhRO2FjU7ptpQi9fmVBmrVW4jNo9lAVNX3aGUEEVkB7Ol
UOx/gIPSsHgUItZ8ltq5CFY6gzmKSorDwIu0smNzLaWRSYd9R6Hf7NfHSKC0
MOfIjLpSpZN1u/uloCE0+/avgNbG/qVJAnc0vqU6yYvT1oGPo8G/MFidOnbi
LMxYODimtnX1xTsBc3MmKTC+6DzF9zhlegSSpbFKicDQX/yeAfl9mwe4YFkX
Qi8gJT+rpuDK7MTa4jbSCr9+K00JaMu8tRe1CwepC+hv6YQXLVp5Oqk1GTDc
JrDD1J+CgACYqakg5gU6EFVNaaaPlv/c979c3LJ/8I8TXlg4qaKHOIkLxSRv
ku9fTmFa9o2pJ0GIdldXgsujmhxLDoFEtrpFpUAQx3nMuW2hFtg1adEKZesM
QJmW02Ff4q/HuSR9CyVjMB3BwwJSVX1j+mvgvDJCsuISTpXOUt9vLC/nXgfi
FdHDePBpMpOlJMGgRWHPzJopD9cX20yBmVDoBG0izs90snnw4pUjYL+Cy6L4
1UoP8o3MDoA9tfaIF3HY/NfCHz9PP7LZ9QEZ/1BOylskeBcA8f3EDJ8jPaI0
ZudURMhnAL4m4AlOf7CPTL8XI1CsGcC2tmqjTVqSqhBNvPC9oKAn+Waretoz
nceu9KtyUrB7vALgfoheqLTmWRb7NaG4L0acBjAdzDMzyGM0oeC+MfY8qFrE
aRf/3XiEe3J4IuYOrjYwy+2tDbMbrR8EhmgZr3iYK2UKK81Qidh5xr3ozjvU
1E2naOJpfYfmMn/7oeAfz5+xVvOR0Uiv67zhA/CyrIl98oHG1kT/PQFmovVT
BO2Kd1QG07RkbPVHVg9wwGBrfCiN8m2hKXtyB2v7w0moylmeV7hEMEor66Mj
yAjnuOxubxWG8WbzJi0IGrq6RbzTlLA41hkTYChG1t6v3vi39ll42iyhQY+4
OxwmVNtTJE6n5wJd4S1CC09n0EMbgELeY5kBt1XErvgxrj288eNVY3O7cTF5
dEIZXBr9KT8C9b2xYUpPrUdkpxubXboVrYKwIIttqeWg/CEnQrbTbV6lmOhc
kZwmGarYagF6vQpKUQrW23l7hhpEmHrnz59YDuhAsg3k20eJtr2t9yZkSSLL
7WAB4DIvcEbwiH0a6MXd7HPkI4CjfwKxzO0j+tvz3Lt8Bwwjg2kvE58QR6uf
Bp0OW42gYW+aa7n5teYCRx5GjkbdpTyPYPyUkm08VVMmFY1iTBR1XVR3+Rx6
Q+LnVVTwPWuVprj7J0h7EIfkVY8iTiCETWJsOAiVFJpBrZ9YN0D9WBLOUfTf
vkFWfKrJLx+0MHI8/XtSxhUZuebrO2OyG2/GHZKiHF4XscR1oPX8l6KWK0vf
j96DXFEhl3Ru7gQoG2/UFQAnS/378lLyy2NE1eHfqbi2BmxFn9NWYwG1Vf+I
dWDhp6yvcHWxgwSbEEJtJeqwBgmiZq+C+5Vwupm+OBZHyt0IygcLT5CgpqZo
4RNaTDnybEWZKEM8RcR3G/UcUlqoRHHteWESBL41A7hA91w/ZIRfP+Idxz0W
u6OFj+Kk2EavHX7UC3INR90derOh+jWNi3mp4CRnKzpqkUhsgK/ZXU7phmyr
sBysgOICtQKzpvSmr8O2W62oJG/oD63Uh2U6p+rbf20i6I6nWO/Iy7vFcfwx
5c4iUaCzmjks75mO+RF6n1IPTomi6hw9HnnLTjf2yP3fGNDvJX+nbSrQ7vDq
955+DodsdieQ1YynsmqFKdDPD/Z6GwI66UiEK6xp+UHG3DpTGd0F77T2WMaR
Ts3kixDbc5teC5gI3jgUl7pBCwoHyyE9AMaQwzB4U6tPogosHhXCj5x3U/Sh
iFy5fQJwiSzthrBsFO1H3Z+OwB6OwFT4uuu6cpo7bqdy1KGgDD2KC/0/dqIx
IFfDQj/ro3kT1tp2CYOaOxFB2aFhjKOw6gBV/vbk40KMXUWAbOz1SIUrEvRa
lnwjaCzZ4OmzRvQnT2CCpURbdZXgQ+afoFGYXvQBnXgv7u3zVj9f02M7fQ3u
RMqEyrO6sHKEuyJKSd7nt3KR+DiIPJAANZQL6EhhOUkoj+oWxrkOhqN4x7vf
02NPtSidiwbn3Eyr02TuIlkUBsGeXGAWVr0/kyI4UcbjVrjrrJ5CIgXexZlY
TBRCxFEvDhD6NQ9LCZg+pzglt29uEtkD6BopwYCMABSX9i04FG18zPDLuQyQ
UufzIP+EXLPkf5jBiI6pR3hykXaaFGYEe/Ydic07tjbMPe0gh+abhNxbKy8U
DSliUYSWKicpazqxastMgL9dTKvOer15olaskaGnyjlkOj2jkxBv45UgYtPC
HktNXhcGJic4vAWjG9MiBOmRwdpYEdavJRyApNoZITDsl0Yade672aXfe3AJ
XQMPLtzwb3hjaA9cg+NBfqq/oKIo+q4F9SuBJ28LT9pDjGHBPo6YC6W1UIM0
Dho9QS5AkeXCriurw0NoL6IG/UUE/XLUD1/qRG3wtIy13NcmZDQ/tqFYLNyI
6zIMdI5tcmydf/1ggjiMzfq4zAZ52gB2YfCZxPnWUvwWr40AE80pDyBS4vVM
/TKCN/P6mtFW4Hl3GtP/6fRARwSeEzhjIociNc4XtZFcFNzdbKGs3qbITH21
m8pf4POKABeBXm2qKzpAF90hzkRhB4WMbX3W2DKz6OkJydOcfWByEXucjMG6
9GVH1io78kCuxSEEwFFRJkSKTUs2kXycH/+Y2wslNGb3bcjTgYNEjc4VmsM/
EefpaBV/TNPi0qCl5i2gkj1BP1CJJYf1UkkLy2kNubRHaRSFDZx57RZ4+ZOA
xg+cpMpole5qOGplmoS/YvPXPMxK8Be2ed4+FoCbk4Yc55KQ8Sm4HG6eYeAq
bhYM6mITfsH2V6tDsL4yvSgIwC38kmSjYt4DqodNVGmV+VAeA2vJCsQFeoMv
C6b2W2a4eEPAaQCfODyRu+a740V2Sc3/NCvcc3CZazzuT96weKKzdfiXlBf1
Jx9NodygYHkRSp6O8VK/CA5jd4qpIFq0atPQMXyxs8mCXnMv6uv4i2+Lindm
SPjjKX1LuJjVANkGf1pjsRKbyZ648jUBoHQ7/T4rgu2yJU6Ni95UT7nBWext
WPmzHSGvfUlSp6DDo8f/xYd/4/P4IZ9dQop+uts6puXHY5Jc/jNIpF6j32JN
FfFd90HuQHOMV0zikAjzSYpO39/74a36LjxBHiIwh0gH53KVW+672HWpd/da
pWxsC8fvXPq7SKg3P10i1wB+cEUYVxelcdVJT50kNdNsO6vVLRQmxvY1wvJV
XyY6toAt8MnXCqzRIyT4WAIqvnViWW69bcVLe4DdhOnrR9y18bOmEGpDTdKn
lCqwbcmYWuLFGm1jVJ95b6CDBSMh3sJBa2cSUhSWsWWjRcuy9/NsoQ7WiSmP
ncjZ2A7IZcATx2OjZym2dhY48gu4bcd0TIJCuUbhj7c/RteEtqvIF4cNpQr3
rWM3IHAbZnd83hfyw/7r8wQk7+2V35Ee9ShFgEEpXngQXUR/W48HXSpIjLEU
rf4o/RGemvvU3USWIdxpaSJxf5kYmDL148/4sLeRCdfZSmrQ93LCXcJ2K8ar
CXzNgeJqiz8Du/CB0Kmsn2zePx6xHZy+alN1MqDEX3wKQn0dR/C4xlt/Uw3I
gc+9rdBZkqN/HEu4965fiw0znvhw6jOOMMuiv0mMcwoRjIoNTzupV9RyAi5K
4fYJKcqck0Ch5he3hz8B94qo+MgA/8i+NyoZpksdByhsvEqnYBRhmW4/iGp5
jGflzlXvj0ymqwbVijmM6R/hBbYVv34WGRCeX2KEQADqOnemGxTcXahPCjau
iYVkOsv8VdmcTcIWLDZO5iYTd9SGRSgmV7+b7xOTQvwwVOATty1xldqJupHH
WTPKYPMd54rWQihp9lJoTGH+BneyKjAmjgA8NqsXEaT7eQ5Dpgb0N9UKnrqp
fJmNXeOjdDlMOFB+0a1BMPYARdm4bc56BUrBOITSvyqey1AnCxWpXEFhqeUA
Run60SlCtmwKl/WvBdfU1sVpE5SVLsFRpLxKNZATcmYwbhxqKfglgSK5z6gt
gkvQgcjDq55PaSBYhQ60FsIXKXWMCn8oXqSieGtvmUUlNzT36LQq1Xdr8liQ
TFUyhCsn1KfUsqHQc1oIsYz7uP84YDrdJlorb3kaIdSttDx6PtR4raXY20eg
wFPNiyvFeWDQ7igkuxf/iygbB0wKGLjYYOBwMHZRhn1+wiXMuetQ1s3D/2as
fWXNwrKywiQIKAMLYzOX5Alv4moMn0+vdaHH/FhusowCs8QVrhIKIfcN891a
ilwXiWMYJC4aFGfHTghpRaSud/p81yZ+LkjI8WmZmzy9pJVkDQW1fDPijLtP
oodc9C/+QJ1VRVgi5jPSqww0Oj7tXr1tAYZ990i03avlYAdAIG5byNjNSdnE
u9XIhjuOp5CdmYaMy0RaVmMPHc+u0+kYOwqXaLdJBjeFig78hqRfTKKx5wN5
4RUw63ujAEMIoOcp1KAkHGJZp0b+0DNDkru8jc+MJNSxqBS92Gh8rlGuCdqu
+JbzWHFJ+32ptNmLuoKA3dgTdUQendtB86uwzRDVb56iKF222vDEv7YS9Mfg
4szdZqT5JSpVVqmIMILIfLsZX8DB9BevQjoGZXsJ5ltbhrrv66v/1pW2snEt
PkUIsryt1+KufaQOwVY48a57pmXlWKKzhqTvG91jJMuI346AmndL+itc5jLA
pc7ivNOxRxCiX42TFKDVmoU7AQ8OgouogcaDC4QCp7sHGghUqhc1wFyA6l7A
HcuzwRKa7V1OUxOp0To0FdEPSAtKsz4ThnnLJfH4JNecdYADms/ZR0T+uc6c
JSqdme8mZb/7/cS87uAnxGTLif7VjGVwy4iXfDt6aKs5yvSJKxjfrzXNBl0z
4VciWiBcPmf9zOIRxU+zUT43TdrXamqy+x+objbAK3B/F+4bxPbm7WKWjH9s
YkMz07zHZEm9J2P4tqEyEfg16PIbs2bqdMlm6MS7gQB8VaD93B6Wurw+xypt
G7/ifGM1mu6bNQEhpb12wprs51aAQdQP9cUHpjpCYle6c2mamHU73t0pE9mO
36RX+VDl8zdnoICThaW214cDgwFr12gW9zAZjWqJKBuPxP+B3MFfx0KRaw8h
IyH56S+dWNOwUwQn4L6egfSj5vH49nT4vGluh1m5Dbs1enKYH5ELHNe2ryRY
Y+/fKBbbpYFNKuDz6ptWyot9lRzrTdi4zE5+3sFY5v/s/i3QfArHHTeMcoiN
WyHNBY5Hm59QJciUcZQp80wsgroWh7WNiArfqxaEZ9qCKBvcel5oQ9jihloJ
uLACOtih0cWoY4z0Cqrz0wyoj26y8jlbE9gY6nEjFmc5k8gHxn1nFMYZTQrn
iunPFSbupUxAGWUcp7jk5BEgSTeJXzTdirBdJUcE4Yi/Y/WNwMoZfYEWA0kH
ab3zwOoxALReEn4Kk57pcygkhVn8GpHVkUSh3cqCofubQfRPTs2L/qt/oa3T
D8vZdIFGK/OLJmqGMA4G5cPSlmZZ5TTYv+YL2Qng2PFZuMY2GpC9QvjCdbv0
2TnQqzMHVLKkJ17FKwu4MTs3BwZxlhJQyaprNtwOnQUnOUirm8TK5RcJxCKz
XKsy56DDLWp5LuhgueREuGzOkjqEfoIG71GNhxChjpQuUb1oVWyDOsCmzFim
o2qmAUAZ40pogXSvxGjHKYjWgjn2UCaLg71QbFbSEoE5l+jMIJSX3jEd3zE/
TmEkZmf13+8GL5x7U4mMqyfN1OcbOnGy9Ack1/MsoVGoBXm5/8K8WvR60Og/
ACY+5und/NY6CvGcrqQdsfNt60I4TJu3bxNlDJkcJZ+f3pKjwTtbL9vf91g/
XWX0vkKMXswy4rFF/FOYWIbVKnYeX+zQ64Uz/UuGu38d0MNB96sfMKV6kbcF
KMDDO8kYQD09O150/kUxb7dknYL0eTAl7gnxi7MoFqQ06cHKT5XlCZiTZyno
TTDpecusis82G4IhUDNqoDQoz6Py3hzRx/E4kHfUvr7UaFL0CVtlI4PVeu5i
tQ1+vaLijxw1k6/XSdAWLu9mdomS2pEYaTVmM6yHYGGEjdXcWYywnvYiRFe1
zD5mQb/WfTgXq3vBsyKgbzkaZRK1pw+mz1WI4fKka4D/gJE6Sp+GNp0ZfqJC
/rY79EJ2uov30CehZW8flKQfyMK2olyVEBafO0w+jpdSXyV4T2en7tPXhYoI
xQARSuiAKfOOFIDJbmrWLlveYe0GuKd12tI1a9UE5PvpDNk0GD3P7VpMjFvQ
1yTgIQR9pV0sjo1UUALjBv1mXdtgi6MvLKjwD+vL7WSc01JAJRy1zer2lUtV
1KkZLotWUvcMsFCDm3St67nPcAqyMZs3MlKtsTs5YnFnR8aR4LYA+nwsxOEZ
yjqcWnZNpadjhGmPxIcPcO3MwD0xakuarKIZ9JjwngtR7ctY5NGS8Y2QF5r5
EvQkliVOcec2TL7krYOC1FTX6pIEmg1oEuesmHIdG1piOgr/FGW9dDQZAm5C
zNhZWeeQNE4Eco+jbm0aS7FD5jRF/bYQ0KjqW60fmsyd3vnzYKPHhptsR1+s
o3FbvqwYBxCdIqd162wTa0n8KC/BA66bKxntl124LSFjLpXYAgHE+cNUgrYD
QrN0PpxVVs7eTq9Q6h/euXb5Wzy+yd2ry3w+H0F6Ueljfxvo+EaK7SPdAZQq
xxdVco+ioV6C35Yjkt+XEo2qiDZkU7YR+/iEuYwdiSjNJwJOXH/QelFLNwDu
YHBLCvdtNWSx2jHkd9PpVrNqhHGYUY0aQuhLsTS0Wy5u57hSolKs42sGguQX
t7ZbeIZfwr8WSCFOBhhSmR87j7mCRZS/l+QqQLDi6DKwxR0XlxrwyRPysoJg
52bp6DodFGoS9nv2VUiXkrE1DA6egBKJzw+xQvh4LbcR6fChcHEYpj0tCq0a
L05lN37gsx7LEWOpb8QImJnmfajHKc0wYOmOpYFgCYluFx2yAfoop5X6DUAt
g9IlMKqmUl8Ww/EKA97wwThrEdbvczEKYwlyK0ibAckRNQxShJzbxMxOCbWw
tYyuVM1z4fkeVKOFwbRD9Gbm8ARvofyqTg9c/PImGlddJv1Z6Gn7ruwQZHng
vdogN4tw/1s2D6cB++RSsBfKcYsFWNH5sqM0hJIVSbV9oGluVo+8QNi9DUhM
h1WBQNs938mfz/GT2LJ9iupBZclq6bwvNySzYG3Kf29+vUpxmlQ11oIkVLFt
ZZ6rhdSFN+uSLKwGn06lX79aYKpub1XMGv/Qv6IhgHC06AmIQtouTPCptqZT
+OLPuQ9lX5WhZxHTCxtLTFyo0UsvHS2BxjeYpgMoWE7zi34O5xl3M3HVsqnS
zoTzCVg0dIh3PHqXV3FqbNOgqbo0BLo24aeHs/QRsZgimzrVfs8khJHHVsDc
Z8j6tlwnG6tBUKRQmiosisSdB69mjN2GrjYvG9VLU0HsVURVB/lhRuAwEUmK
L8JDMkdQ4w3zLAfe0CXNXrF+s3SryDy5v4b/bW7oGfPk0dRKyOYOB5x6QXpM
yVrJXEfVQ1wb7abEkX74M9dH6AO9ql5x3SkD7anyAECPReKWwhy2vwlMjuVE
gubpc+rIutHYnKo5EyqRSRMt8Ys435YrKk/UXk0zkG+LHIvhpjndW/Nng27C
DvfChOENRp/E76Q3/p8t3KRZTTOzMOmGOUkRbDNA3fhgmdZ3qhsbcni2XAix
xqi9yfo+m/6CpKYwxpN8OBWeLDDcVZRtNgGVyAuZc/SvG1fMo9tZiF2nA8Vh
WEVig+RJGAJEm1V32bbGpBbgV6KqerRc+jxha/zOpZOuMEgIXfzKAei4ifoT
hCfTMIroCC7hSwph17DV7NZsvT2l6wPhd1cLKvNUoe0zO5JGjq4cKRHlrKm5
7BtjJF/R1QUAn5rCfXfxlEN9sGLZt9bM3vY2/3zuqQtF1p66nSqyvWdh4bwx
3JTie4N32Zp4zpHer+SunPJUJiyTGXEr+X+yVNp4vocNy7UhzuLHdGucUQsc
cIHKxfUJtou9Esx4HxdgvYO9CzFyd7syxMRjkl+QPsX63VFqCAoJmUysajJ/
bFih+gR68Td8ynHUdAxQ2iDvhUKNYr+ysUnlQ0mat9n6xMmR4og3JFiZ9g/S
ZH2beLgJtQZEDMOHruWAyFd4W9NHTmvdHutemVHciTSyEX3o+b0rC53meVB/
tR07iQw0v4PHTshbPfhB0AW7u7W/2QOanc1UvIT+AyXgkHr0Wyjnu4si/ksz
lFNHKwgd8VPtcISoyDhzgvD87N4EmAyTSJx+lFp6RLRYnCi0Xq6hTGiY4zzW
NXEofQshlDlB+6Ns3KFaNe05oIaLsmq+Tej5JJSXZy+pGohXSgn+RxZxNBTB
ZdsxO+RgU9Bwk755/mPkeZWEb7KTDFi6JzV3fpx5C1jmNxtc0psQ1i39XDir
ST3PxrRtNbZENpPIlChruXjUj88CeL28ocosnV7ie4K3WycX3lDQCkys9x7u
BmCyY69x5WcULeo+mZfwmr6VL2WnhiqdxlJM6N12GPg4zv/7WyNrGMxKYkXg
9WnlQfDWEjLLokl/Kz9Wlh6SLhAd/gTgf4iI3083Ibl/xzKmhV92jXdW+vVY
2V2ayRqpEJ5Ge10OzdGR6Zls/4vdWNpFar7yv1x+MmU267No13ZTL771Ncwe
+345GA4P377oi5pAH6YsqlivmylnHqddxt8ev6ti/I63ItcDNbfgotoJdphN
VXbpT0zVGUFQr+9lAnuG98Mu4wKR76oiJyP0ub4jW0ccmpE7mC+VJaPdXjg2
wLDRcm9rfa+qJoddn+8w+lY1gI8Ndi4QqgLOfJ1Bjo/55X8NhBSkUZcaDwIo
XY1Ch+95esLAIILI7CymQAdaJEP+jBYgZJDao6zcJh69au100I+TgMgXvG3k
qAXIjVPQJIQ8feXRx+2bmlWlE/oPihy+Y+qz1FS+x2zOrOJK+FlJfYTT7+J8
xSPdIuprfGTCrMN0qzq+SAxqSbES1UcoCDf1IQ6HFw0bCRt4Idp7+BIPZW7y
lXFMgZFtvLcC1EJd0BMbsSEMSiDjJTA1M08a6/AVwMAr2xD9tt3xXqbhqmC6
JfRGz5aIxMEA3gP8Z9RR82Yal33PMyLZk+pzfPzPWD6VvosfT/sv8X3cMWSw
prXjlzcsprRCQNRuA7I3U9/VgUoNvC7+Dykm5prERTNNxvgtMQiVwHACr/No
hTRTFFwKraa5W6zMlZ3x7HB4j+qNTNvIfxre6lFFqHOivFzu84EI049vjH+w
8AomxlROqA/eaYJrrSxS3IOL0P132/PlsNmkW0FaxPj9uGDG0RO6Kzx3rKhf
gK3agSX0d9gtuan5tsPhGiN3I7BXhQPyVLr+tNZ/rYc7WbAZbMFZO6MmDwzo
oXAVMqjXJMuRTbxe5JnDnCGlQ0DrSOGJUoLCSLn2GPCjd3HLlWLiJ7KwL7qu
jXrmevqROaaRbJ1+HhkoMABv/5jroZNnabgk6mK4wKWWZMWKdJB1saFX2HDL
wr1/jBRZs03QbR6DgrzOw+RfZ4TKFfXtU+b9agAP2n6xkCmn44UPRbg/6MfP
7pxFiR4Pb2YObcYAv8dqyaw1bTXvV0I2ircp6+9mCzA+nOB57VUJh99PGzL/
PHK+JAdJTFezXMV5U4e17CI8oS5KHMeGnbG1doy2Ysb+dcbx8I1Nx05hPe9Q
Oiz817ECiUx1bAFymlrB3lG+Mo4bl1D0SsxrSsDvZvgvCRBi95yzsNKOxclm
e10XzEjuNkHdzp1XzCdP8NTy37JhGqLqZ97AkRA0vvpLhdrjD9Jy++8zUnwo
QGL9x08SWVlEKbXcAXEHs9LkEIU86ZxVTMRFmuyFP/FC+hf+X7F0v5Flq+Il
oNTs1STAg7o5P94FVkGkafkwoQmc5Bu+t1jG1pGrWUa1XJT9npPc41bhjESx
ssx+yFrG+6FrGTUvcKiHHeIbU3G3yRJ74WlkDGfzGBWGMUU7mgvftuQtI7jA
x7xKIcfyInmnQ46we8aiQrvVXU3z3nGC8f7K90W0HYpi3jZxkpr4cZLuED4j
e8BlGkkT4aQdwZqTootYy/sYcb0yaScSQye8N8AVJA8jXJggNXzE2wZpR5yj
BF9XxaOyaurgHOIRmvfE6KQf6DKQuXeJ14dNlLfOU6CLv3ooBRqr6fR3KClp
uIkO4dai/kHZIEflDbBJcCQ0TlsDOXgm9sJeiQA78kpQ1WKoLHBC3nfyFHYG
b9BNn6Uwp/z/idCqI0oAFGTzzhDo4SKcFUrOvoVqnLtBsEyqnXRa2OVYTkgW
Xuxbs5ES8uXBjamnIwVbKH/zFK2M7rHmg+7EhcxkJy7WvDdU3cAPMYz7L9QP
peDzR4zkcc9OE63wfF38pFnOM+XNHy1d7sMPMDszS/38TqP8mac25QVHdmtz
3sJ20J5Mhu0IiC0FaLfPT5fevvZsvbZOA6f0Lvob8LrqOn/r5CCE+sHq9IK1
rGkY/j8giGYccfpNtirgm8DhcuHezTZnDL8V8pENveP5IWNGt4wDGOblplRP
z+h3XNqh8CNNxXQnnuWhdosoWqZAFNrWCI+uc7EEDxAwtouUylSn537LRAvt
ES8FV0jfN0bLQU/BQOX5nA7yWXAsEqUXdmgTEtBCgwwG6iJ67EffMsiE4giE
Z3ZcUVFE6dMUkS+OkqnW/ogbNjlKlMeKkm7Dw6o63IO8kpR0xevgdgVCVw3l
GXTq6Cal2Yb3DzuGCuulYFEAxTIP7fvPS7KN5iVjoI8KS1I/QONhJLfPReI7
kVEzS9URcdw0DReEJTKLBKRcapBOQjwWKdwbXMpT3BsQW0iNGGkTYhlbc1tp
gkFfSJ6BPOutpQbHKPGIk7U1T+hTlH20FOIfePNYR6Zv/EPWhtKHc0F5Yz3W
E5/uvc32DlLI5nFJXm/0S7VusHbT6LUbYRYY7d+oSnv6Ncc+/ULx61f5K3/6
+pG+SZTQbATSV+bF1NL8hBUdu/XcG7/YzSCzXi4L5+ab7Nh3BEPBHjv91hqu
dcmLUR2eogndln2Dx4MtIob0nROZERh9doaolpz3ogx1iP7ASzF3vGCyUSJc
KoTQ3pQyg2QSIp0pKBvhBGlcgx7JakFYPVGAMm8VS4Ief4ThwiWjUUep6Uzc
mQ/VAivNLlHhpnyzoPxgD17RAWpohD9tlDdmag0xnZ2cDSHJ1ji+oxc9/t3t
L/hyK8IVrzw/MFfpxkXIqV3KVgPaOWVNX8n8N5fbSe01wmn/oeDE8T+fTCPJ
BAnEdjHRIEi14xjklHGcuS5F90wxhyYa+Hh32xXFtiXQERh5oHDsYbV5RG/E
8O2M7hvMV1sUBadnlHnwHSIR7NydkG/TKixHHe6Tx/K3a/JxUTpX21qNaFFt
uGwfMy8QAUqFNesRMhM0xwSE0/K2eQKonXKHS9MLHdlnMy8NIsh+QgUV7Spb
WruI3oH3J/m4q4aefbazUcATg20I/QEE4q0MMeYRL55EkBA65sKPIa/FuyIH
Ak12zdfZTCKOdyPg4YaH+S2zg8DN9rVRDebdJa8BKp+/qXyD9sIRlSthz5OW
wgLxSk2f2sT2z9cn3v/stUI93GDnOCKmQ4IDLtD3pXPJisstDIBGnPD41+bv
vkvN/qIGIIxqaTerr2r34lANkiHWGCn6dlFzk1oi01s97g9WE14DUprqwCdC
5Z/UqT63NKSyfcogFiuueCgZJgxXREt/DLKGsvf24CwgCbjM1HhKvkCy2FrW
0enKLLbrd1ORDMCNwVq64HgCB8IgQ6/eIN5TgO6gxSE5GE5zF9GOOpVBbm2h
dxcbpfh7P7gF87RKaL02L+EujtSyNkCvX01GKPlWdlgRmIrYZD0pD5TeCpPH
5VUrj0/a3ayMMfNLcEpR+tQOBfp4bHKQTDna0LWOc+WAbFRI68qmwPq41iQz
BfVDdAJqsX6UMHT6b1Wf4QITJ6TGM/yR08bMqtBI93uYkriu40l5v2zjn9qr
bnc5WZrp7sc/hBKT3bD5cR34EcOQ2nx+rgRp1WoJYTlkJU0NCSPvUPE7PBST
S5asyR8aNsaLMtPJEVwuD9T61xKmzhReEKgm8yrcQjS2q7MiKMTMlmVUYxjk
OMKYBKf+XM0UKiI42Iai4t1gtnOtNfOq4qK1FnNQGqVv1KUKfS+DMXMAZ18c
72VLoK82E7iuF84LjWB08C8UfCPcuxgJuJ2IuamGQ3m0iBjv7+1bpFnmVB4N
o1SnXcPlO8kqOVdCrNSXShOc1jAVI0AZg9KO4QcEpUGB6ZFKkbvfwwh2TNL1
3ORC2LkLhiDANbYChYWmTcqoQxo4ulPYzpu0/loTG3JO4xvU1wM2l9YtkZcu
LRRxF9Ck0xEWQ6qraIveXZNywnzvmVcG1AYO3c2jzSGO+5McjwHtqri3A/2V
32ZCzOGrOLfJDzts9u231JWtFzeH0PADRZslfGZHLu3FeJMLSghQan+OV2s8
tpuoCQTmbzmfgqvC4rC/61YDnE5BjZwHK7dJmbss0LzB2K7SlxC8A/GFq0x3
rWkAPZw7yK/mC4pZxkyK002ANkEotFntTcN3rdsvG2t5yOqko3SuctSDJCf8
nR6GcRbfDZQKca4Ly4ANeHnYnQyko4/Fhe7YdaTjQ0v68P2CABW91RsFJ68j
2fcG82fnpSecnTr/Ev8lpQ31veJbpIy1vGnsjNA9OpW8edv/SC/0aZsh1Ykl
YuFZ4ForbVsGWmTqlgmX0JJDzErQkcVNGOYZiuDQrUYMnpWSKNBV5UaTCzLC
TGM0o1I7NMSD9b6WRb96sQTSdNI/P0w7FX0o0zhJdd3WfwoRC4C8IRXbNr7l
+R5du2TIpXlERzjkDqUCNneBzOVnOUa1WCn4OYBj+2ROn937fyIR1pott0OH
dY31T5fvpZVIRFTEAjRsmuAce65K/w1sz2XCyJ/OLg5fzrUoSmqzy7dwvdBY
HDupkUARI94UiO5Yqx09k35Ez5nJLq2ImsEZRm0ltRWfQhANdXeXjNAmlMbu
WLbyT1J1GwSc5Fh87fgEtqbzz/OpCsJGDqmL7d9KPr4rXNQyV5nS9JRVCKl1
IFiP9DTOxtIVEVcV7MCMlX3gBTVmt6rzk++F4KILT6O3Wqetd5kpXDo0KNtw
i6aK5P5rhGHMoZ/HGJjptDuFDWDbN7KtxwomJ28VDgluwNsrblLYsiarVQ+Y
FO5VdGGOXVwzjUZiB4gTGccliqi5TPblVb/Be17Uuzjn6eaCvn+8xcn0cLLl
jmCfoSDExzBVfxmn1QUps0j6DCAgL8XQNrIRKMw/YY9TZ2dm7twQV07d1DTw
2xTQ9o1QUwzKj9epqUQx51tn2QHtSHp5zMJV2mnwen+UnA9fGgYP+C8qDVqR
G5+ULUe7DuucrXelXEixfyUzvUvdCxbqDC2lpjgqJY+lxQ2vuEJK2KbWjfxB
u7dVUpPsh1hh1Jj+hsYWbVW8UnlwLhHiKP5n9RuKPP6LmsVcoHIMSB7mg66a
yhCMs1Z9sDRPpufqj/PohzY1y65ZpSRyQnHmE7QfZpOK2tnI1lmz4OqGvj7L
DBt7gBaVNKLzFoWK9/xrHor0BdlSpV57shP+c7PH8hlZy+kyQ1bSQhBSBYW3
3TrBcFIoJgXKh6lJnKVJ1p9Cwqd4IsRMxhQ6L+ekvxjvrAAYrKv1wl7cM5ZK
0G6Jlmo8+hllDMJkAOYb7EjUITwXVGZoubpsqmeusjiBrCrmTIMQPGWjD1SC
lIscQzVebKiqvJE1P+anYgoZYEVvDNP66mig7I8vAeTOea4wJbWFxqjHvOst
t1J+nDWqNbTcCk247ilEPMkKaYrv6+fCMHDIPV6bCARDOrwSHjhDMQi69CTO
GpIQY1w3k7jCxOBLLrr5YUtPKZwhzAy9gauE5M7gK0cPD/zW+ONvqW35n/Oa
vuRHJBScp0p+KHpgdGVYq1o0vF7xA5FWLgjxa9TSPVlL9WvgK8hry7RvavJN
ZKxf49MAMhMB7rUFCkiBgDqrBeyz1XKQJux+Q0IucErVkwjUZlYPryhPUJYs
frZ5F7InRi1cYjmi0vNwS8tt1tGAa063NZUOJKs4fS0l7mcOEXLPJQJTINFg
4FQA5n/NXzUmXa5m+L+vCkYfI4KwMFFljNbSSoMSJY1IBvqmo2Ho2xCjxbMW
OscEaiZTnj6rhBu6VTPZoVpAt0//uRS1YjtYSWK4xdhELvIl/rTY3/bmNqt0
FzuXdw42F/rWyBY7OzTpF+heAQ0Ga5Ov1EUgW98EA6lhKOYn6q/+0KVEwJYH
kiFF/G49ku4hZdqmZ7bqX1qqOGZV7jGbWarhCjzcCcy1LzGYod5YVoy+QCCP
GJjxKXXwuLujpQBfkqogeMwNcAgs8I+uRKQAeqkf0U/Bm79UCY+93Xq9CjTW
hxLuMOwtYyLKQj8yHSuPFB4Vqdy9KsXYnMcRy+gRWgwN1nke0yaYHilyB7O7
IegPtFJz7wHcOo7iujBHkg3KTHh88808nm+inOGY+qa8JL9IPkMyLyrpEtGB
vHHKCIJx8zbwhJ0wOhLGfaHeeXwfQJuTV4SpSamujPJpyJTZDPFUuWcka5vl
+x8ocrr28vXUPqIxswZGGMWeQJILvOYPeNqlXJXwmznh8gQ1kodd5/W8m+45
yRm4tYD8JIc9nNftIgaBr3ueuSF4XDKrsi+ZV5kN/ubnQCiGlYoWFiXSBpiA
C0Y6O+7CFPoJR4ui/kNPvYYUMOJ8hCzOqkTCkz+L39ADzEQrkyMouwKYKSL6
4SWMB2/5JQLe5WlSGMldmVVzxYeWp0vZMmmN6jPgUW118BIlbCk/uaLLydho
6Iuax2FBN7cH+qalEN59W86UttR73Owe/xIzz1oZ7eEd5WGqgbCA+7bgCGP7
yFZBts/3arLhlzJNvdPj2uJtbXrBSL3KLh05VlN0QuA/2jAm64MrSdZ5a0XP
0jATCsQhSk9acygEX497Ry53s/byTYS8qXqlph0rm8IgTfh8pXl4BaT2A9iM
A66TAxQwPKAJhByqcjm5SJ3g4VzzBtmso5xlNoYX/cDMgJn96rtWJnX+jkHm
yo3Wcymx6FEHnMS1SFBSpSOi21zhWq922pBd/Kq2v8YLhFfoWA562xU4chyC
qyaW9/1uJBWknxrYmNerSr6jf/AfNNeErSF4vmJclFWy51y4dYkqPFR07dl/
5nP7h6aZNLag/KwzqE22b8QG8kho3r8WK68IUh7oQuHYQnFQDxAsUhI/P7/4
N1SYg52KO2lgQly29gpNOV4ZpUxKTU6zMjgNABWf+75GzUTvXSIYdBbuFrek
2XgHdozILL5Ct04+3iYnjZbtkgunp1wdBmMtykLTMlZAjNSItBr9V0TP8w0P
9zNHBJ8RiQzvnFtPQLWfwXxsWHGKVix3b8wnqBEQ27Q051H3lKk7IhfZsLRO
1XIpSpPmVQLxuJfAw0+SHWWCoDN4w+qyOxDjRe6E/GiGuPpHNM1667g1F5TI
ESMcLLWjC2xU9Ia93foqbaWCpr7QO/meUVFqZpRDERzeZnKLQpqQnSXxvskU
dlXQ7Zp7ROu1MkuZoYQJlLgjyqptNMxjYUI1mPZHIg0ibdtCVtIRhFnOcwGn
0gLOkkBKw64r9LUNqFP7hrl+ENxp3Mp+H3gBMFA2116Av+7DrFPK3a5TSTsh
2IgpbN1uS4GuQQA4uNa6NkhJ6rNkMupkVIeuZM2jaT+O6I0xxRXnM+OGuLoV
TfuROROJ4N0iySvDOALtbxCYtVM1V1woFsKJF9vkUoXssq64Eqk6BBvYe8G8
UlR9pr0PfNl4XG/IWnoWOBqmz+cX4pAP8smoK1uVD4EAaf4mdNDejRKvKfNU
H+uRYw2AL+rjvZw4GSKok+Ptz5g8CZwAfuBemeoyMGQLbnJqBTs0CErwUYGJ
a6NDbxY3CrmUsquvRfhD6y1Cko0G15QqJia4aYuwZ7lXBzpWlVSxHezwNvNb
3hD79k6HVWesMppWM0+jIbhnRCA3Q+bpp75oe4D3elQSg7+UA3b/0ZZW9Byh
0uS/vwb2qIv7Y/BdTrTk4Ur1MyDDfxFRBF4rE0czTRXJRuQayj/fOL+7PTj9
ifAt/tbdd4bi0y2i+6+DaKx8TyxCeVZtSoSGbTyCQvpi2UlxkDRxExLzUDlc
BF7WzfaVyAoOEjNABlWO5JLsa6gN5B9J4b5BwYo/I0IZZENsJJkROvWjcZfs
pYUFbW2BSJu9gEfK+zwYbI75xHDmXjualMz5DROcWn4fmR/Qzn60FK4bOGwb
vjMk5jmj1fNtSgzuhBABST50XkTCpBWtVVEmkukNQhEMrHyMwbTg3vB4aTtK
qbM4drQOkLZU9ppuwwwjT2f06YT06V0s7zsh6T4+cNetvojuxEH/pSji7++l
qqOiFXolrwP/uPhlg+9vMhqvC4qx51+/m53O0oMXKCSDo5phsfY0813kwlTg
DGCgeiAbleXFoW6vC1TRdsaL342NDp2rZFX8KR0XrNWPSTW+l4UjqKIcdoOa
faCoDiNagGlRuS0fuIRbgSHIsY8/mvydlCc3KIkPgKHAgD9gP8/2x/IV5+dk
omP1Sd6L8P9tp2BMQ1oIcEJH0aTWx47LlQdHPbe7vTFPsaMJOZIwhiuLd7gW
K56DXuUAHJ9bG/Hgl7NOtkBIDtWuMhMrNLEHsnG+4EZWqDS8xykHI7enSjKW
szQZbkz+kuGN++KlKxVE6GwWRXnIyXwS6u8AzRyXQ3nY7Z45rDz3A7dqR2Cc
NUsOq2O/pYOz24CiffqeKkXhfke2NxgkYBVHzXcmbOBSaBtjQhmfz8EdVaRx
wxPqRcOQcUYLXeJgZ9bCT9y9iej8EWTJHBkvZBfeM+ETOmWfXP2Ftm2ROpPK
JPFEpyNaPOGKjXOedp7pncHJJrkhvqO5rnH8oFss5AQv03CuPCfByXaHlqiF
23iB/ngVNnq28mYpTu+B7aIaZGO/Z98k4FzFdefi9y4tiXk33M++mgLsP8Kt
MGOwWKWU05yFlT3LMcLihkmROAHoA/TZqWi0mP+W3b31l+sRgJ+ku4+z5qdw
h16tqBTGj+W4XVkz8jdo6fUcPwsXh2W+08if+FOzMRkPkYhYDu2ULrMY49oy
ZvZjG7mSmn6Q5DZTCbTqF9NyVGXS8LEu14xFT04zDXBnYLoJO2o+ZZSNSEod
O6+hQYqEBihgIa415w17XwDCxs8Mynm+axpZrDvnG13v1DOKRl156rJTcbK/
0sLjt3/Retf0OZEChwVmPG+9rinsz9AIuuROXOcy8Zojt5k9MXxoYg7LUQAP
VD+lFIH9IR9hPlmfOUfz99cRbivfbkYQfyHJAxizTJeQYT1kBla1QQfyiGwU
iUhx/UGDNk0ImZGjhIDlyEVUof+FNmA2LHSslHh26s4Y17uJ4cfPXAEMpZjk
kjDsPryqu7q8DPO43ZdZkQiwDm1Sl8sXdjmnr4XUVEhY/9GDJcYdyVi9mCfk
EGLKtiiqSWyGS4Rle12NXOwg0yjR5zgCK2qnQ2wnMFWl7VFHkrZil0sNvz+B
Gt6vozt6cDMJt1tL6D7q4hzyjpXE9nZg66sfSDS2vOP2OQbuDZayTvrae2a9
UuBXPe32N7qQjJAefMwtTo84F+7P/yBdZpr6Ry96mTIEPvuMdo93l5QDts1X
p6VQhmsQ8cHssXqtsDmODTcMPy/u4O499QLqROnJ15WOmSqdPmSFHYB4mJu/
9622WJ1r3KD4tNpuZYeydeqdZBHYVqtyUk1QpweRVXqYZXpyRK5nGiaS848q
7Y1SZiH52jKe9uZcHMkrqbMuJMlSlgu9+IFUv6gTDex8Y0t3+V0ykje6bUkV
8Bws+Fi107/x4FZON+0oMosWLJrfk6ewBLR1cE2meXLAEVjq4RJblrBBp3XP
jeGx3OPcxWYrUPOy+bHVtoeQ9mXdx3tmk8l9x7NYc9evjYGLtg+lhanvw+EO
VoNKNFx5Pp+DkQfgm1Q0/cZDqD0oHBOZjUQGR3Av0N7zu6g08ULIEgh7sC8P
/C6D/YjB1s7xFPfqewyQkjG+gqDm0nbcVMVZx9NKicwnXDVDAO5GgcL50cbk
4r4foKLkMzfylnw/qzHqFu4hiUj4gBzRFgoQtUpGja0b8lCdpmt5I9YXJQb/
05ctP196Mp2jCyyQUnaIB8e5drlP+4rsabMXQsk38RU5fhU6bzb6Vc1GQ9Kv
DyM6Rd6d92MoClwlgfcj1yubdkF4XMiQ1BNVmC42HTaC3cpp0bXsRFvrceNz
fD0zZLdh9SrFzBkgbc/3raE6GK3izKa3s2HXJmOEtO0MZu9FeACMDt90gUSJ
32hk+yvovBNLszO0EObU7m0BvN7Kc3BBRJarH+7KrNaHHJ3oWzaFUejRN6JH
ZBKCzjkHS0Wtdk7LmzCySerWTLbQLMtENKKPUz96F1Arfv0NmQ8QgwfBEaQd
pj1yaHnrm05doVIDAUrkvzc59DG/1te/5GX982rZNOlFv+CZhn71fCjZWxwS
YjcoJ9CysXEa148pD4wJGokkpJT2l5olx94tdBJM4jVRmCtW0uzqPskQi/Ok
XJhquWA0P/tPaJ2dJAulW1LEiClgvHQjgjDgZ4Ad4GFI55EmE8ecdgZMhEMo
Yd9aWiQiVcQYobf8IIcTexi2z+1A5oudHTrALrthyaMZie03B5IWBiY/ND8B
HRgGKzfMLLM6fDaA83mkK2yrUuFLUtcdv0ZeyNevTKKzhsJTrsMzl+OkQn4N
Cyw7HyUuGBZB44OzXcOxPT2u4E6Mvhncry/Sy7seTowmlRXM59drHIOCtBWo
fgmZORWkRgGp+yv3owHFJDV241LJYUFuAqpR8NHAIoELTenJOPA02pqjaght
RIW6mjFXv2jC4xHoYJvhE/nxbI78FPcWl9zAfM5H8pivNYSQFTg3LaAyAv6b
fUK23eTuHLCb9qPiQMZ8P2L4RflJI9PbdMiAqezlNLro983D6k5UHMwrh5wX
gCvb/EkWyBQaRkDe7Sd9D4JLCMIuB8SPIk9GIC/llJ28OcGNdAq1pltq2E4O
Wk74Drb7214fo72/hZeNUWNkHhlTGrAlmbZd+Vee0lHLTQzDOK0ZugCrARYn
dXi41PcDmMWY4/S57x5mZYpxT7bFnBpcGTC/5Ns0jEJgXaFG/1Qi0jVNhSvN
4l42H2RsCcbJiiTQfuEBfWg1TSgGT7Ltm1b6t2QKrCHNq5oqb7mRE18X4jHd
2hazeZqS4ACYmUxuZ0/ixy1kH4fgeqABxf3iQRWpnLplxVOATp96/Bby1zFM
DBVIriy25ufYvZJDCVrXrVn+NQlB/bS0wVg5T/wqGzgeKD7Pys/CCPh20LiJ
VKCsaWAjpVE/xm05W1s8U2ieUt4YayFWn3uZ/olGx8nSFeT/YuFU2suQFZeb
rC6j1zU/9GVPj2Cbj0Ef2ldx+spLLgqzY0y6AYkEpcAn6Uw1Vi5zFRVOuPTY
F09uP63H8ocqxs3Uso6h1ilLhZbMTR/VDinsIjf/ja8ARgt47gVfw2UrIHyo
OgQgFLD3AqoqFX4GoYUMdGSN59Mc1jTnERcs5rP81/ALyLFaytRz/zXlQ9QM
LnWy0gC6w3UimH8QL3htuusbSgf2fyefBY5m153Sevk9ZI1KJ8eITViPzXN5
Mu7ZlWqnr0GS2Gl/j1mMh7K5hNc5tAAh9jcngRnV6mB/V6NzfChUR7YqP/UW
fSh5fMosuplZ88DaNsw+PTqh5e3/dbCeCUHvvL2jX2LPtLky+zLELkf/UjYV
wltN3/w6qtpE6XLzNsHuSrM8+/jVHz4jhG9RNJ5oT1kY+kTLvSl7axuySYF4
MKyTRyu6OyyBbUQUBVu+sDZlp3a/kGBaxn3TmB43ipzu347KFE8taaZiOxp7
ZndHMT7lp504iymd01NPKDz6kxXO/dWHauX9xKaPElIaV5SsAFgvfqw1gXD9
NfhJFGzcSJNjogsWH6nrMAzehfmCna3I9+KF/d26qeVhI7sjub36KipuSlUb
yWs4n+QL1O3iEKC25oKf+eMmg44I45fTXcZPkVPxLglJXj8fBPNu0vHdYnjt
gONoMoWiI5EyNVu/JzDmXV1cReIo5re9ec7eLLfsFFKlzeUwmR1X4CyphAXI
jyg+UljKZMLQARjiVFpj8un0KYbpuXSWjo5Kwh1fZESb77BIDIofVSv58z8W
ShAVCRpZcBgfZt7A2cg/Z1QwdRV7MzRnhAzEPuBB4wBC+nf2xe4dQLacBeVu
Wv7NofZEU9UHkRWb5I9u6Y4JWo4cEWoj0h6A1Q37Giqd7UKkmy7G3Q7+7K2O
mKViPTjIoJMFXDNKSswgAFyo/aMtEpqNee9t4vqDiR8lA6I1TOztV57yrtdE
u2PhQgsVcStHXPJAmVrEy/b5V2RbPGUrxN54KUe41SvyiC54B57a7pjfhVoO
WnZyTcd36jQJPFH8D2NObLOwW5NHzQEpxzGFjOwZG0bv3CkImIhTHsvx2oKJ
Q4ztwCI0wFEFyzqmBf5drNQXcibKnV3PTrA8C+WbeEjKr77xBQTm3tR2eU/z
tidha3i71ZuvRKmZIh56gRCZ0tlZXRt08XUAPpdS2EGwXDjXzeMyU3MpsZ1j
1PDy0Pfv5Vplw19w32JnfZapC9JfD4qPrv0K/oQfwNflPzj/I0BBAEiCl18b
Y23VAs4nNRMrkrYCyjjQdaKjleyEpR/kQIoFXe1m4DMxZSU9qAp9vTxa1H+T
5I+4zUC7MCFot5PiCyHEZfYourACbSOOsXJwfgGH5RjJAwZjPhciGTvqilQ0
z7nSlHgBsz8h9sO78QanslOvt85XDkQ4H7STFbuUnYNE2XP+NbONoozsMItu
QIYIj2Da7OQHv8i0S7cDQpzSX2t+e1Prd2hNXVGk9wJMBKSr0V/p/QewfFO7
EeEKMKI1eH3eC7P5LHzPaP9vAU7VJhRM+mK0xrXN6mA5sP9lLuMpzRryZbzZ
ILPsdsCDiJFfOC37LUphIPpp40JKMWDA/inNnggoxPM9pADlquXo2ehpH4HE
JPMQwugG412GjXh3XWbRmZMQwLRjI/uB7iUPmZ7jX4QTI9jPB8hn+GaYvGhA
5B20aX7Vo2m99uqF2OZgfs5guu+AG9MUTW0YfEyG06XokGeSx0p6hQdmWXYU
Q2qs3ffFbVqbl4f0ztsXFBs6hFtc0hEXDCf/1nXKCVOaoVqYFYlGoWqNFSWZ
uWCq/WOqZLr5CxPypKsvuM8wF5rXhiBXd3NzmO7PXzgppfNx5CV+4yqoHz/F
UcXrQf83AJiTvBF92hsEXZzMaThkTLqMxmldTTu9NiaNV4qpl+nC//MEfKBv
wLRBjApD8tPpUmmSlLZSuwkJjfOa/SGDJ5u/gKe3+QPkxmpAfoiVQ0gMYIJm
GcCnh318KHxWe/AUsKEcNvwfZPy+RwCzI97HgpGo9JrtJI/cPr4DraewF/0Y
zMALPw/+ftsMAC8SUqyuFUDolnAfyaOkfUTUBmOm5WONfnNcGTK9W/5RYAOL
MUXbBezPzK73F5i0deX4rcbEbR5bhiLBalCD9ylY+XTvRiNCjVZjvvuXX48p
JV1fe+ruX1zqSvzoeDFQ5navd4WGfG2wXPkA+7dPA+SAlJkIfVJJeTEb16Vy
evc1x+0wcHR5RqlhR3qNdE5fDiovqrgNvn6WjcoPZ6HZUb9l2Zz4gtVG

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJsmnt2iWtIlKHLiLrY5+X8/vfFTH0+zh5mC7Y2nOQVHnoPhPhSB6IPgQ1RdDzcEGnoShiegg9GRogmzAFHOiNpm9kOlLLzOqEoVncuNfQzjzxNLD0Z9X/eXDsB0EefTtJM3vM8yNpSpg2FgUdXvzdKZxiUtrqDxAbov6sdROE8Ywi/DiRc7ZTYYT7LtZZgZmk8Uh6M384oebHFBrUlbuUdISIho7sLYqIVI1f805qHKoFan381ELCHtO5tkeg+f2GOv7/wsjoZfZMvpYRA2G0Bt7fLQ8huxPES2r+LyWeN7hWMjWxlu5KGjgut8Kw+ziPJQObRhtd+xYhl6Cetf7k0NF2WfDlW5e80asfjHefAQXvJWIzsZaeQ2d768waP+/U2iEB9tQ6ITFn65Y7Md/Q4UT64e8cusE0kZY6HyCDLz1RQJqNy8hI3y1NPbFgdqLaTZzKWqxfHCYq30F7LUlOv5nxgG8Lq1MBIP6pag158svXoh8kFaJ8vIM5z1b3/7uF66yJPURr4r/LFDDd6ynFfD5pR9KMK37+Kts7LeNUCkXnvexD9O+egRe+gnh4iCNkioaSR3Q9nBjDAdrExyXkntsNn0OujcU9sD5NhQFKlP+aE/zZx4S2TfeK7Z/xdVDydX+kPGe0sTErDHI7PQ779EcFm3eefHySU4tT4u+i83eSaSlWL7lD+VGWiu+5DAVLhh6q34jdIez9fIVuTDWX5ZfqjsmrfSpxHAbyJtZZrfWcgHXc+Yt8Qn5TEMiufIuJH+1JClNsqCAeYMmLjaiIy"
`endif