// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yktMmX6mHI/5cZ3Ry6OPjvd9nWmJIa7xsQm2R2YlY71y0RKuCdUu9GlFoFXh
sj2reSLDTQx9S5IT4pxH+dk6gm4KODqvLk+UzLmFUdcmD2EgzmvYbV5q5GTU
lKRDbxDHwQxS9wMMPTwXdiri5yD8zgKdmGn8LWXyWtWA3evTscvZSXqrbiA9
BP1Jh3iMC7ADTHRfd8E0muVu9w5tU9d0XQaZsXHq673BrOZ1uny2joQAAc96
iHQ5YE6DKTl66CUW4+dXz+HW5ep67R/uJlU3TAmc8okvzx6DH8VmwRNcw+te
+IV8pQHw6CceRvyU81EWUPJFBgJJrGQ8Eeh1vKdrTA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Sa8j5GmN5VowejBZk1lUrbiOWka/8XLxUZoFtBzJJEGKsw4v7BxOnz5IbqB3
CD1w79nCobiOoKeIz3QaRta7VA+i+i2/mcqCyWV4YX3eRVMf6XzZWQVMheWm
1AV2Fc56a51kUL1K12IfCQ0tGvKxZhJGXROOApLGlu165k3Mm0rJ15KnokEt
eh+Ct7lK7HYta6j79QyzO51LEhD47VA8+fUNEvQiFA85vdEYNoiBDtQreuG1
vLlacU9pt0klzp61LIkhtbn78hjCD8qM6emK/Kjq4qolIo0ThmDPLRm4sh6D
WZeGSfdJBszx+Gebub8j6IAMM1qJGE92asHzZMuUpg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HtkJ4+7zwcKj6nWwAEegGsJiMcSqDS+qcDRTaHGT33uxdoI+bBpsHfKWVoCs
nLgYAnpFZOp9Onx3onxrjG9y8WdmgrI5zqxDw/PdL3UMMhOiOf/rsDj3VRkK
E5meg0QAMl1eZaM4SvWYZG6PZ1Q266TXBuwfKwUTZw3m58WyXSGgtTkObGxU
8Y9o0kzN96gotbcxguKXlxumyaIMLmEYSC6tTVV1Q80cSKUNsrOC/kt6YyIi
KUVgXUa7WVr0iviGNCkXXAn3QiAyLkWMyly3FMqQP5jHReYopdPFH7R6+ZT4
ooAEdfGuvp9DY3xZoxqoCCgayIsia1MqGDphjKxU7g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PVeQy2CVeN2oqvju0gzsBH638EFl12/w9gblHNgzSpNo6/5UYdqSI81zgpxy
CbfhlUFKAeoaLNrTDZvsz9Xkc3SGFMY797LYIQuyO+dzH7171cK3HnbfQSpT
rmRBecKhTL9BYcyPFmRRDE2PBqMamHpq8Y9I9kUxf8ynjPWxydISJE6h9kHA
5SWd7drn0KxqqS+mC6bW4dNARc8nHCoEq+RBmrdUhrC7tRu6a+X1iLGgLxeA
cWvqOIWooR8m6HL9AdbMcU19WsmYOdbzzyTxRhYU1qmI44idLF2my4kpf/w0
V98lzVEAkokYAQL/mrsqe2+hJlIElOc03pmpS9NQAw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JqZQGR8sGLWQ97hewn4UDpMcMCE0H3paDi4CuiULj0riGmW0rAqJt7KI1u2U
9iKC2WFz61RCRdnu7epfOtbNo0bxGnvcInzAYv7trua/vy/+6zSAsV/yG4Cv
g5KdxXtmUzjKmJp/tcJmpahA3S04w0xac6rl2O9BFQZzQHoWCxg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
V/bkJHDaVT9AMVjeJoXWONAyvaoVVjvXoURuUrnrk8ugoG9Temv3XMIWuSRo
jk6OYv7Xiv659jmI+lrndLzbtxRJvpzRHp0+7Nh9WFVqgfWzZnFMww9r3ekx
nqs+WONgB4aQhSsSS8O1+ifUo5wSWQNR24CoKZR5flEXs7m5SX6l2U1JYVWy
K3OuO+74joCNe6vR5rdg4IAfCmQ/MP2ljHEpD3er84yHhxxkAGnZhbxf8/Ya
4C4ilYUnZLwKE4utzUu1jgepmDUTbq686kBfRe6cYr1ibYIg3RyTB3oL2SfP
cG/2aEx+/nsdQBcgN1ET8Bwzae5pdMryglpw7w88ynwtE5jQldUBWHS/VjXF
zXpqEkbGnKlLh6xyHyFIclYbG2DLaKVrW3tbCMFnCqbHNDxt3C0TugYAWGnc
NtztiKNaeFQNNb2QKiuWlFMWEE0N8xHx4NgMRSixPPb+bDWnPmzS8Uz9oqIp
CohbMj9GpPr4NmKFnasMJ1/tF0Ihao6n


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YnUDmx/NbZQDD+QBYYf/EA7IgQBspIs/n0iYNiJ7l0I6n8IXZs8YPgCUnbwJ
/WQPkyjHMK1ZwEObxU5oZUfAmhGF/BvPeY2MkD+HGqYsY27J7O3gR6WOKcCW
K54IrnZ1rRRXKje9RdJ2iteUMjyKlFC7CeZCbAEGPsuw/Vbul7o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B4j/gAzDSntircLSOhUK5DRjYQ84emUFHlqh7NcFMiTgV42fRQ/3UFJpq9m+
7QrwzoIRqwXI7oJeHg0xdT1n39cFqfS+RudU9hA8EsMLtVKSz1S8PSs23Rf3
CEsOk9wZJt+Jjxd/LGlrmLEc/kV46ecQK1kNdMO9ayoKPgpB/3I=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1232)
`pragma protect data_block
4Cj1nS3y6LvHa+0cXMETrrgyZm4r+nidGCOi3uxz4WfGqr+9zH/RHRobecAt
Yz0rn3lt6CNAuYmR2wN9Bgp2ZCrgORLQHTRP7nnYl45c+F+iPLRVX76zxloy
p6AAnPpEPU7lrqFIWPoED4oIA48kV0Ggy2OzF/boNXkfyhYK8tYnuLNsXj/t
dKPCgEJXxKrMJY8W4VGDTUCjWdRKyFc9jD/mmT0dgdYgJjSfcZ5bc9U4k8rc
ZO6T4vq+jjEcr9O81jn+lPDIQTVO2Vhmg/WFF1FrdPm8szBV0CyYB3mVk4e5
+NTu3qADeS1ZgtMzY/Muq2vtili7dvS1t79Z02DMSf3/19k6ATtx1gHi89/Y
ts61uhHTg2gh3a9dwejwvTy6ISzeevEHVhrj/bMoob0Ywkzl5O7VotdEbkbF
JMWIlWgJKAeztlBL71ewCy94dyOrltoErg6imGyBRZcFzc1X1+xaikUvLXb/
2zKz5KDdfGKyRNYAw/THarUrgGXYppBV/nuddx9WFrPEjCYVvPQCFxlRnfIO
TwwE4yzDSWlVokl1+ytb4zCyaeHe98fAv71E25oXsZOgchqm4O3CuV5jmgiL
CxfqI8USDo7i4w4J+nzXVgRohW+YOZZRzwu+0/QCiN7kWsWDyPciwhIVo5ky
d52+0SSdkswXtrBniy4gfhjiFRmdFBA6QjAygwmnJUDYNK5If/Js3foeU/bu
GFLqNx+d7CLVe5U4QNfInBmvM11QRwc1O2nIDw6BPGejmRzoPE3ZamZxIe+P
FmSJZ2xyYJHS3UIBrNTtTPJSxNjrQcrFVFswd6vl3MJXj1H8nc2p+dOHebI5
HIIRVNHyYtHXJBsSgEObDJvGNIzqGoIgTnjIjRQFlrMlpJiUAO5EcsKg0dp9
LyxJoTZU/NQvVZKlTqINFdr4tofUhferbxagyj1rSM4d9akrnsCQrl5yfUH1
1KaV9eYJTW9QmMhyoXBZKSZAvXi0AqB9nsJCNZ6Iqzs0JzjsQRTbi2OXKXmB
yJZ25y1S5U8Zj56y6XPrdDbsLYGrbjKHJobB3izfELU1bGUAzumHCMjahkyp
LfbtfJXluiFe+8D6U8bQKpNoFHZb4JlRIFXJ44reRQbcW0rBUEeJsxnN+dXy
yFH38Jd1HXSCDUMvGb52yZTbT+I5pZSX8IQJpB4ZH2jslCVxW+0bzQ64VqCF
qHUp0ct62rEznsWt2/D2Qd0P/utz+jsNVNGemF2EgDBULkW+myxKqPLdFPoE
NH01Q52i2UTx+idHGYMdpcDFj9bowbDkxbinVd2k2gCrNOdeIK0+uW5jfYLQ
741dC5M7vbvgMCawZzmWUAWv7OMwpdtOyVBJcDhkcAegGe06Fj+V9yQdF4Tc
bSm+Xg7LcLhwaucFPJrBC0k1ULYb42oA/edgzBN/0hpMB4jBWZ15mhcww551
Iwx0OoDT4dIi7pZBQSuhQ4GQ6IVdwFDs+w96Lhalf86IEP+qyV1CNNEiavXF
BrO0l07nKmr8SthRSEzRs1vjipI3z85DjdUC+QB//T4VOb9QH97AOS/52AkV
clPzXc9sq02vRnslZicmjoz3lVAo79BjyuOlQshhAyvczm6ioFN7olXJsodt
lnmgtphkCtSd7tDAkbsBF0c=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdgCKF3vJMbpWWIptHs324+att55M7wSdSbpCsbojyzOPEhKh3f9iOjZzQsP07yrCQWiyWqwnpTbSPiekVGdx2yS6zrahKKfgpbBZbUJpfZB6MKrj/ZmoTPpcVcnIleMw8cmWFeBpJBKxJiMAY8D6u/00flmwtNWstH1O+QrM2p0BBGhgEBI8ei3m9KgTZki+MUWMiLl2to5LLtebunL28fBEHJwMU4UGAFSIASY7pPOHl1evGz9qOVqNxrwqf37/AAYF1fkE37ruXDv5e9IV2S+Iut0C5XIZuMpwc7SAO7md1ZUMijxjwWMZaGYZiXQ4V4vm5n+lKsBda1RKmEPyc1HqlVChj/jt4kyXr9CFNJA2RXvhfrwFv655CaThkWdq1VAoOIy/XHpyWtlAKt8aERoQNyEgDJArGUu9zRaO5IXV1X7jerTSMmtUvjr1LjIjbuSNCTJy4yNCQynwXKQG0I4YPP9GV4DbhWNYeqgE1smLKcKPycwQzkSXJzw9MoiJzG40i4tNJRQPCiY7N8quqK5k/q2+n5P3w4zcL3G8NLPqF/oWbBrSoToF63uFAHnGSM1MxuYjVZ84IrgYZjQMKp68dFB0wwtm/HPSLOHGNU88R53OHVOuecvXhsGGfGXF1D/GIgLurV4lHStC/M3iImT1OD1uwfQeC6b4iHkmkTodbhWsIMohOukhKqvbXKpITL3tXOi8NpI3bDRNUSt+b1W+xRcSTGIfFx0unZSEng+P2qzIXefn+hfXenvXdX6kkFRAcb4RiDv0ZYifBujNGP"
`endif