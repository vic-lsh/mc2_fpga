// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i6rSSl84Oodnp8Mk6SpQxZD5M6HLCfi5A5l6jKsleaC/KrVSo+T8bk8iie7b
bois6M6F1dHKAQ2pKWC24kolUgX1c09t44BVemGMtvJqVqE5TzyjIqanNEJZ
S7qqfHma8ezCj1JCv4prFXWnVcicV6cjbuZKpMk1afJG3W6gJvlsHK6/9xLt
z9BAZzwWlR0Z9WXStppEducQK+fA0BlyzoONTSwNVVhiKq5IzfSgfymj4cOs
zr+23QHgk2pSs1KG6BF3EqGaxv+bn9Ew5owXA/7WtaHXNnE0xW+kbMiFejZR
1nEIO5zbi7GxSOZXq+qZPElJmBmQJdf2YFjyQJmWDg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n9bJ37sfxv+qhgbycQ6heKcZRfrPLWwO4zMTtdj3OupCl8quvm5EsZKm/ZDk
yEzg/qyH702+Lurr+H3je/Ulq+pceYh8f0PPgLLryREyWborKGulv6rsaQCy
G4aIu+UZJc8hXE/Yf22gvz5356VMHlhVWPRkoM0NNaNDHdEffk/jVyktuo1m
KpG0TGYM5CHH4iOQXSotVl6GaXpkK18ZlczJLAf4UO59HVSspQJe7mRtXiLA
R0mpMA2Xz4XUReyVoWjnurF5YHsMmyTLYZwpak0awy+tPics30Hz/eLIIeft
KwGFZ+PtSnRxLXhGiBzufBQhLQXNOm2Uy+uQ7WTgoA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cEb7DRq2eysrpBPh84yattNJEhcxVAu1ylyQnu49VkvyGmGB37FG7kt3xsl4
RtGpBY7M+JSuXEEhdwuruL8GZF81/zjumZ7MGvRpQvPDCrUFhIs6YC/g3+13
UkpSSIMGrILamcRk2GjF6PMJ4kub0eUgevLndcrIZXXvJJXjJ2eExyo0FLRr
d4Uaeda33lHptZp8oyLr1Yt8T8a3fYqldVrynEJZfmCOO8ehKJiVP/8t3XCd
8GXyuDAnoWCHFZtdY4FsYnxIRrvGbqotSBg5fnfi/ktll/kq/LddWyghWsP5
5WdRns7wTEllXAGN0Ly/JL9RFgAAkBsrWjBLttULmQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oMtP0h1XkNhBM8VYh6muAeqqPVE8HmY6bq63ek107wcjrkTiCRL56iYUJIbB
Jqq5oNQW7IS257mTkZzcrfhAJtMTFhM475GXRlkPpVTPvS9lz0MFYid7I+z2
fDYKbGVbYqGTkfhpp8JughTpoL8oRvsflxkGn3nPrbU0CWYIDMrL+ezrFiD+
tPYMBjdj2YHkjA6iXP0C6dgiPd2bSpY7VZRnLjMXuLADL3ZOl8WMuz/gMoQ1
6GqKtIIZWa3TX6HuHMCfr3o9mq8Tc6Q+4qdLo7D+cMa+WCbDKefV7EaD4kto
Y7mmN0l2p2XrmQh9ElUejj+l/5ekWGihLl/0pb5tdQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TCp5dVF54BaLVHqpSnaJVily9sZM3rBIkdQjxCxA1Kxc4FO/LU3Qw6l0cT5j
bXwNDq6nKVtFNnC0cuUr/6m/OGpIj7Xlqnj1oyDWUwLbTa9vAC/NjKBGk4wy
jEhvF5hdfsxE1baGxdq+B1hxtyNBF0nomvBQ9LUWa6xCn59wmE8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
K5m4fN14vVBCTknDCmBH2I2kX4ihKg5Vvgt4sXS50qsoHKj7UGsp1plb8oXI
zpl9ZTjV4OkvwmR/Sz+3i6Mf3BPelw7v3eOg6/I8LXbazCsUQNsMRoCMtlow
7dyp8o7n9zYp9CyMoSIIFdohRk1BPigusNYBTnnaGnWZVPijAiCRc/QF0xra
HxY0jGOGRzFknx/9Z9W6AzFUpO5UNBbSb/f8ejv096/3TEiy8Fx3kNxJSPSb
51t2FZ0XAnbXZAk8RQq84fp+VS/HpbU1k9zornBHPVd5jxb8YRh74hiXCP+5
+6UNNo7BU/vLjKY4Z1TFneKh5XET50LCTs5SxIQME4e17lkLCVgqf6ApbCaM
lKPM8hInSCUTpEyPmpws7MwCqyFPoy95e1ZTQftiyr4xiUkeEhn+U3n7WYuL
+wnqgqxh9bKWLH8tdnQVt0w4a0KL6VM5arGyosRm2r5tBL424/LEFKEIAdma
4fbfH0t+A63ZdrIGAZepZueM5LsfyEgf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Al+r11YQwnM7209RrSqFxmMLjuY0/n4OrkyHFJ2ixxKTrAR7I60PUUNwpW2/
Xo9BFuqOxwFm3bAbeUQtO0bE8tsReNDVyGXpdQd6DnO6T2tFJr/B3OedAY+L
bM+1ol66y+97e1td7nIsiSywCiV3ymWdjcO83UqOIF+9uoSUUDY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bbKq24qbO62NmxuVmSletx14m7/4rKMTWci6JoXXOpYZmpeBlEwu3tVWiQd4
hq94QrX8IOQtPQLYES8DLbb24z1pfV0qYY45+hzEmixRMTdzmtLoAVLQndm1
kwREsmCG9hgmyFt5QH5W0yNDnPElLMqNz2twulKi3d0xVeXv59M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13184)
`pragma protect data_block
qZjegdtjtP6vo3YVEeHoEzOVWt5a7dyq5mUyx74/jX1Z6rzvF+S/S/s+MO+9
xzrpw2bbn2l/3oxw7Cbw/cg4SjTtBgJb4BWztCYet8Ore/8OgWqOFoW3IEIV
VrzesyunM1fOGDv1Bg12iNdWq1v0x4NHprbPnBqeYLSTXtRL4g5n5UoKt+xR
JJb+AVne4yPx7uVeYwW9BgqZQd/4f5WlNabkKGXvmVNKu5KTotTvHz7YvLWY
ZrNxglSIbMcI1Gcau9Y0ZzYJJ1LnkjQOxIg0nP76Aek0YfLVkSUFYrMhgzed
FwZXxTMSlw/X2jXYa3dIUbp6NaoHZLoGutS+xTdgago7BiKW2EVz0YpGmO96
C/ewRxwkybyWxM9e2ramdDPgnHMvsg4vUGzwEV1sGJDB7x0Zn7wp1cIKec0C
VwJkm+yuc4eLlk9ePDxteiPbVpVaMBEaeW8CtRlBCefsY69n1C7Ol0bGOlrj
FYfc4BOKY9tX5GdUWvbuhhHtHHw44qO20vXU9hBB/IDKmCdofb7VLLKsWfGr
Yi/SKoOZe1mTV9i0dxJveER6dxj6WCvhDvaIZAoMR1Ypt5V2meYZGh2naM3x
/sZhl6AXP/FCxaQqeJaRxh6d2EbrEoQxau7PCvyhqrt+/UXO2xCiow/oKOls
TvXujCM1tQKjd+EECmLR0U+YaxA7rpHau5MkXqaNHfcFxgHWp0iZQ9WRSZtd
qJgeG23WYCRjGYQ6+DBWvRph7r0j8uwbvC3G1hK5v5CC47UYKZIyjIbN0edC
k9KWC0Rt5YDN7dkMEOij5WPYIFsYm5YRkDqIVFUem7sAHo4qPmbxGx+eKdzH
LuBwpQfkfQ9uFSdmBGvcJkxCljMV5CjsmfAbkWACuIU33nHX0VGfyB/9kqhL
09BtxdQd2btDVjshmVryJNCljNxGWOErlk27vIhS1ElYZrjoxEw5L4L+DQa3
ZdVPTVW/RumU+v7euKrGryC4U5Gqo0MWJ17n/VViVSab+4KIU/xc3bhT2KUS
ygCIYsZCg7+e3ywB0uXrlldmYY4b/3IVZrH1UljvARsPMFiy7gSWmJ/RTY90
ThHxUpNe5pha2YLG8Z6zVPBURTHuLx5utuM7RNEntcv4j7yh5YPMt9xWjGlU
iIm+jf/6XNLqF+ToE7R0U0K60BToHeedqECctujaFu+Chx651VEraPvkJs41
HFWeTYZQzRwYwH3LOoVMg286OzNjQdP5I2Rp3ul6tTN5bY0WzWV3gcVB789G
YGCGl9byFeys4SpJd+IFTp91ZgJrN0KbwAVlDRJ+QSZN9tqaiEtYAtW3cw1M
cjn95/c/7SoziTGZZCN8AmiPH2i5Flndm+duQSRjJKxG9Wn3DZvnzhckqItf
Gwm+JKr8oEmbpvvP21f3+q1fW7PYOCNjDUhWqPp2yPzQbNCnOEKXaCHNLKVz
JsXdYZb4fCFxy5fHvuNXYwMfwVvXJzXSeq+Rn6yvwAayU2mpDgEcrFQ3EUJU
e+J+njt7pa6GTUvRRYVKV/uZUl3Z6dmAasO5idiLB6vOrvQR6StOYRXLJtIM
Wm/iOyttQ+Ljio8C7guOFlVcd9SwOvtJP/Tg5nl+JRQkRMKzGR3wrQ9GJRoM
IWSflc8Ry+PEp/mwnAeZuL+HimCTUp97qrtZbimdSm8NtcvR1lN12ynG5/9L
LFb3FZ+90IGdly0unXXRv83YzM+4oFrBA1d9kQl8RFOaRXguG8ThdUH1lifd
958Cg15xLytixSNtQPmk7LWYgtHMTGl/cKlBw309SGxCCuANlVCTjXW5S+RU
/5IkKFFZrSMcGfJXrtQpm2XodJ/WS0YwiJ+h+uxRZ+LI+rZEJYXcNZcD/GDu
WZBQ3Hl+3fUZLq2O3bJqxmkWHWGEI9v4xxp2r0TVnZC0ki4xASpnpyYFobqo
2v0F5JM/1reRhnz2U6/qsA+/zKoX7kwLU5Co3Y5lU5VkWay1sjBRn1KtJAJU
oj+qVz/7dlm6l1aGhBUz/2dkuE7SCIsqkpIwQiobNhl3X7elndWIIae++pWQ
10fzTl8AjCjH/HKbdPaeR53h4qH4N+qjavX6oKzLHJ08D5dKDzBgSpxglY7T
GEcADItI+KkBTwp46yYlaqagwlcbhSGKTVTSAZB7SbwR0y5GAFomzNywdUyd
bmlCweNiFeMPGOBcig3FybFhBqd4a6Arv+oSclEFC50F5T4EqNShnStnsV61
z/n/5jkAHgDQn+AWgt0QF08bAq4n1Lzv9Ts/Tv1A7HjwJF+QFUMxxHbTqY9Q
h6bvSyyHnsFFlKdUDJdd2ivaS+HIgzlYZYMb2AisOBJ+EEkswEjQFNlxOvXJ
XU3/I3uqtBE4jLO3FZsu/4jR5pQqYD9mtMqm2J3Zll3Pl9Ux/BXq8FBU4NNw
RWATCzKFzzA8e5FbNUpyJqEehEjGsgoIRr9MR2nmC5fyIMUFXKb/nopsSTlC
vlEzbv8hMkAHgqpFd2ODGGTdv1Y7PcqcFlxn8akeCTRZoNDTEKjMnrueMATa
GaFmdIGgxfiyz65bzINh27c/7/TnPg6fv1aYpnz0MudEpi5rTFRI2d32kSb3
9ECodbqmq1TCxjgxCDIBRP29yxZ13Ib4ez8TuBdxNeYSVbFFKKXIqrHjhJT5
kajJgaUOoF1ctI+zP/U6msjIch1zfDLzIU0PVezT8jJSemrvITzalJVH92Y8
o7Yo/XEPLeMKXocDjGEEL2lLvYvyEYlWtfl9kW5+6CRzSqIo3W2Sil6FibUp
uHwYfVYIzZiu8xSJNni1/jiDGXdj6RxxZORKNrkoROpLXI3nPaKGbVzeETbT
YLrRXiEyUkimiy9IgixyHTlDyOXxuNzZEq0sxMCpm8CP8TEBTpQt4w+ax45/
T6LLml7VHa1RpR5HXwKgIL2EI4Vz2LjkzeHx/V1zS3iMFZjmpu8bZpinbEyI
OrE1+XNpV9KULvei0TwwtLjRmPn0e/X7Po0LDtRqIbmDoDRkv0gHvvXtB5of
GP0Ndg+vmrwc1Mf+Bc3ydyBHu0We7imt1+SwDaudwlOLFVNF3DSG0ql9UgwB
vStGsZ4JWF3HQSt10S+KfjSlCm4OdBMuniv5uS6FaXTlorfQXQ6X9Qvq2/MF
x4B5fm7YyyOooKVzZHM/ahWxa2ciEP5EVfOdruBZw3ukrNuQQFICtumBmww4
bY9paOujzxc+/57/O37SkGS6F0tmFzoTHduem6HNYhaoXgKfamdnxDXv33fi
lMaSx/TMAZagqYPplNVKWlwikZxyUEDJY+m3z23+7AbWDgOruuBwYnoHyKm6
2/wFXsCObbhqLFyXe+IaaNXBrOyfB42HhIpaQCOf6hUMm9icJpiKQO3rseP3
IEqWdgY+fcVPK5hphdXsbraTXxpbXOLH9mT006mphurKhr86SdQukofe2mK4
8q4DLYT+PFhpSy6iRYtFSbentUMOkub87D1b03hlpxA1GcdYa2XeJnOKrgSi
7zC1dY8k5EPTtEG/CazpoNd+RHPBjzKK2Xzoxg0Sk3p83AQH16odUo8PgQeN
qK0xWMJQRs9EEyr1o6kYEoprVwZsfUzioJkxTX7H8lHYEn9SuuVZWRgnbnpm
msnbpPxkBF9pd0QGyu7D1ZlUfQCpIpJhmS+7G4xIIWrel92tAMBqc3AFLBgs
kngQ4/S9BuV3c8+a35oeP7PFbUCZ0tTjCw9cxLKoqiSHGknG8UmQ4LJ6YM2H
XrNGzDai4x4hiTVCauXq/bqz58ROV9ZrG14hVI9kT0Od7Ynec/THNghl9U+X
ZTDiGE+XOqYVPrcSukhW42JA0OY5gs+sYWEyn8NMxBsQgecNwYDXAGyLBH3B
L/H/GM/QGGUqSBkjig4kQS3sVJ7OkLmrOjD6kCyqzkBl0tFYo6eFzQhLuV31
JAJY9EM7IckYQ0MTyxbz5VUq502I3W5Od3zj99F0zeBh1indI3wZnBVlbpPK
iliAhQBII7uJgovmshgE3WHhoFwm2ZrJdl1ubrJcoyBKQ8vQRxns1k8nukot
a6RbDZtAXz/ejSoy12XKG7ya73KSSeW9ZfkgjfhonmqBVH084PG0toP3OKG6
WQcjaXQTkKL+YfwZB1hJuvKNAE4iZ40tj9oJ105mSUXJCO45bWiKoEKTmqLa
ealGVpZAoSUX2w5aFEliDVVDsDRKBPCpkHAIUZqIcMsnxWlDfKDBOvh5oPiS
gQNdm7f7E/iZQmZDYdsagCgQLUYBV3t2q/KJJuxbQkJurLY6Tlw1xZa0TuSs
rF5rkDIuZdWryMMCHStfTF4R2WGen9AlvzhvAahcyto54NRvjd6YwWEigNu+
VITS/MIJDA5YeJDoGXQ8oNEOen1sDj5jHQlLBaSMqhdiEyXDbs46WGPN1pzu
Pc1+/i96yKVCuTn4TFRURVQQEeQQ6HDgLWt/GBGJ1mua4xJaQpqoMzrV86Bo
ssBkDGaJtQF1CvKsuh4BnVqo+hK8pRmwxCWyFZ/F34v3HKcr27PiZDWYaedx
Ej4uMScwRFAfJ6mwM0bQ0uw8pP6IDAP1Q2/5SEgVs9IZGOwzDIlOrlV2jIFI
u/Ri2dc/fYIO/8EfdLtXAUT86JJR0XA2ixJm8tx8g+UF3BnE0qQJ2iG5OwDo
BLkoYDq/IjMbD6QLtOuKfNZpm7Av1UCmJNokeWVKJfgDQ/LbxEk9Tc2/GYXt
Gwgyy4bb3xgz51+oUYy7MuaUk3AEgwIZgmeDNUON4mfK8WXO9H8TQIJvT9qz
FbSJFsN6SyCM3TE2ISPliAx06XVZHBZpuAPUf6hIyc5fDFxju8uGloRHmBR8
CMLc+dMYHyBbmTxoHaMb5gD0E2/m55IADrbb43q0E4FdAePqyp6LzpZB4CW7
fzPKeAwdlp5mJARPpDVyZQLtdcHwsuRYoXQc/sjOyk1QhBz8ZBpSV9PYRZLJ
SnOaWvCOf2X8xiiZK8K8wEr20wMQbTTObFyNsbPKfloKb5/3UbNOpM0Hm+M9
UTwtRTPAyE8nnRaCTglWLlLKOgAta29+W+SclpoaALuvuqCO53ogTnt4aBFD
acyWS1gQdGvFkZ0BpAcUecNrzyxFqV/TfSdbuD1W9EZlOPMDvuLqNVbU9g2E
/ylTyl88DVNsLvDZn67hRpk/7IE3Ah5U2gRpzmgISESA0LOE565uyxGs/D2y
JyQnF6i3AIL+iEnH2vApzcdBCpeuOWpfoXarJZ4W+gQodkBoF+G8JnR/0s1d
I5N0sQiytzzl4lF/ESZ7x4Jr11EAWQ+ZOB9e18PLsatFuwpll0nAcFLgcWjV
cqF7GDBUbb/6xj3bYeak/pQBbPBLI8YvRpB2ZNx3ssJZMALkB8WwdVf4XDWg
wSlzN18tMs1cGLjr4XUU+dCUfBNoy9Yps9IheVQom9GZqZ4KaTaO4r0EqjfF
Owr1GeiapLpS0nhWgWP8CNj34OwRa0Yv1v0eEfdMphkHRKjk3xRTcr9mda0Y
+RoYUCaFGdWnK66zoJbpHwmYoOb4EnjSS3/lTVeDl6PKinsFi3wkppzWOR1H
QvDuKra1x91GbOKw+sDcka9/MiAcLwRZKUyL3QkSq/qbWtH7y/aR/Zn2noLd
3Q9aJPtm3YWo79EwyByYOTQWhLGFCwYHkO2NOAOk0dF/b/AdtO0f2QZMYBtY
oirGSo0GQUs3PbbGSeOpRPk7BQy8OViTtBzKbo1JFd+v/+P0BPchc1XD7pWv
UlFvboxkCXtIiu5kCivE6r1lYrPcPpZPtxEBuH7Q3JDIdHj8yQcu2tNy2+H3
oVGDtxL2LVYSuh6+uIfJqyZGjUQTgRs9C+dQ/mxrzSCXLvdoe4odiMWprFMD
Essta14ACgYGDirD1ypfattlUTTgDM2E7vwb88ABU6F3wFInvXUMWp2riRU6
Ln5IhAS97L5nHe9P5Qv7wNJoijdrfx9DR8QeqBEdxmrPnebLvUzUn5Yv7h+8
ZX3q0Vj1Qh2ft4+hQxcob5ZS+I93zFNoQNmxb7rQbGPUeIWYl6SyPRy7elzG
TJYwmEhxt7ZVnSuf8ArCgUb2a0M4bexB+gPwVSqTDSg5EaVcnBUNwGLLr5ue
lqYoilWsTs+bdVVXY26Yob3if50Li7AbbFn6JVEKj4vSXbkEQ2oTG77e8958
2a5mWhcBvtNgzKaktF4s2rcMxzN35TxwGtXQbdbzh0edShnVcGDLkX3kunoV
A5eC/QnSU2QKnT5WH0w1vt2badcNYpNYXRN6tGSfr6LV3RqyHYGHCnwhcUVw
06uaSfeYWzJE6OXbBdpYnxNuznEOrgdY6XM1b5rBHF/Fv5Np7O/0910wsw8G
DkhCdiWY0rGMqx8BuNAJ4lPrQ0q2NMxfEuEUkb9QPhfPAdPrROsRLZKqQslb
G2P5/tAooCvYN2DdMKJfGYQPwEL3pnPkhhFz+Jas+7vxZn1a4qLlPuRTD/vL
rifBs11tLfMi0ROtONorUoukdhVDb8ohezHA/JRPj2lA+jdSrwqOntmimsvd
w6dWgX0lvrtTASo5Lp2pnbkkFjE5th/99KanD/DKQr2iIpNYb933eY7qWqie
XUh6Pjxl1QZ8SVxVMoUXQMt+vvWfekITKqn2NWqiT2WxcPIpPjcTC+WwwK1y
jF1A5IeGqzio2vSSLekk0tn87JTXh+TjyYSdbEyEVgeQOYgDu/ULi2sYa6UZ
IHmUyMYYcjlJqqQPLIkD+SNul4SYz+2+o+ryu/X0aJnwdk5trSCfunrbN1+E
SYBrknKk2A/2uqY1ArAFdNRtqWaaBQFL/+ISQMLXjPAPd+/BOeRPbO36M0a7
NJtVySr0UuydLV15aG7Fatjlnd5JyyUHW7NbTyYt7xdfabSF/vZDoiP+Wva+
+guR+IGkL0GrdY+/SwMTJeuA7J+GdX7wnrsKxZnzIWKbSllFfnJ5GScSsOzt
FS1gxktCbX+N22sVxQBryJAaePGEMBVI90NljSUfG0pc38Usi3c08mMtY9QF
zC1gn1I6gD4a+WB9f5pai80eWqV38HCqin2T2IFfKN5+fBlaRROcg1YPzaSU
8wp9H0oRq0MmcYivFnTsrUafA+YXLF40+9klGLP5clp4wudetu7I5pM36nSe
8ZNFKILJuvrGhiwsJmkp1+rHwADx9wsSCge5hsfgjE0zzEkjbIAq4UcMFq8N
B++8jhZ+lMmePpmMvPOQCTaEnL5b6IEyXsaUqZNL6Ts+UjpkAqMu/UQ004pZ
VCoZmTlYxSjjLLopq1r4ekleAgyeWIaTGSQf4wlGAqsZ7TEuhTJ12P5Dvat0
pm44xZ8Fzqb9XQ4V1QHyQ5LNlfyxRMJFZz/hpYrzWnoTxAjstUj8RxNGDFu0
w5xv/B0/H60MumllT/WMqHNFiRtqmjKwEwAp212OIj2O40x1gqa5y8UxhL2x
I2D8cpDxpDC3FWQK/BUAftHgjsMh+CCDlweTzAYi/qLUMNB+Hw3uR+ubU1Pw
EnG1CF3QikoFiEIpV7FUjSnKjXobGvQi1BoHfj1XUYhq27guvRcopiQ0sodP
DMJTh8M71JpHhokv1kQZoVFBxS7+VHfA52DgGcXnjvSZV/RelrKfiRzfZJME
cGCyQioFcuLKJ8pr+ldnqtcKuNDnwFwB/9tQkKdQ6MkjA78VvFVo6dclu99y
/oLqyIcofWh2MbY/eAxaPj+L3zB0AdLiIGVb2QyIzpl+cSFi6XcHFgH89ndF
1H/d+bJq+SAaWhNrflKaqbVHZap7gOvyUzeW5lOJFRZmq19izGreGkltRvui
/t4J7RdKh/vAYo5e/hLQotDXLroWyOSHCJ8KbD00YhwpDVJQAjS6rig5Wapz
wTTECqnyNjpRX9bO8aYhK/G8VEulRl7UPEbwH5quXnqCD4hgbjAnN2Wjl/Jl
e/4ItXp3ep0EyRtO42kA4S3JOrHnKu41WbryCKm0IjUB0vjyS3Vx8Ksve79K
nFVrIopid2i5dtAL174/q/1XqE2shUljA/QvmL4JAecWiQciI86VFADEQBGl
PnOsG30L2EGdZiH4cMyvhxWztc7pBpW9w8mQydWP1h3aUii+0hp6uRWj6FlH
h6Yc12TqAqTyLmFHA50JhGDSubGcQ7x+ztIYqoQ2AhNiWEEyHEHmwVXEEBoS
RGSICc/dSks+QFStYh6jt7Cn3tko6y8mczdlSH7QUtG9iP+9vH34nq/dx3af
4+ti10zDbzt9x/DoBQmHD3qJbLKMlSwEq9maCNu57Yr4/u0tuT0l0gf535t3
dB0GGnBAELOTZ8EWtCFOr83L1y9dZcRGOwAS8X1qX+al1OUnPR+LnqEQOEVc
hHEDMacnlh3nM6aLq9scuYnFPD7sohTrMlc+EwbCVSvMh7q80mR4ASUJ3aN6
b/biw13/edG6cVEVqzEdAytWRtgQADHIjj7SvqR3axNWcaJ1y2aZTj19kFSp
sogHKZmNmarpbyWuNQmq0rtqDGkvTi5eDeLj5cgfDj1Wnl+JP7jNCiWrva4V
IpiIawQL7u4P5nph5FazZKSCh12Zt952ijDMmIDlJ/6Hze081TnYotCi4GLE
Ht6s83jkfY27Ag+jf9XtYyQ/GL4z8ftlxeRVdwGVFmiV2ne5s0UvS6tE1h0x
rflWhNs1bFF++pq4hAefbnqfZmK6y50Brz/fi+4HRCBuyLsQWySHW4mebxeD
MDVIAeT/xUU4jpqXQxUr1AoLvNajF03X7IIBe5MnFXR1mKROVomn4reQL99Y
hnrABvWx6lzInF61Jn1LSlsoyoAGy4ccUahPaLajFPwWJpvmipD1Zj9B5FIP
E4+y3jLlT37b453nU5jEgP1vV6BjYVT9at1dSxZC7FGBiSGU6lMPUDPnx4Ci
QS+UgBNPib8X+4M+dx01MMYqMw0INMZQt7WVszYh7WJB0wTJ4rwqv2ILwbq3
AsED7mfXUN0CUhsEWvhrk/kH0/dno039t6c3tma9CmDIAbA5GInf0xE2bg+Z
Es0ZhkFETBwOCHq4SbPPErJUHXLUhn2J0a1G8w3Ng8j6xUj6j9ZECclsWaX+
E8RYxt21Bqfa7GkN1p2EesMb6zV2OtkMgKlJUFlR0gNjUfv+wvUFThg47Va/
nngc3DhldIbyacDVSgcVIGn+er7Yh8TeoA2c5Ev8Qh0i1OmDSvFyCG1veUEj
9FmmG9xNwJ5yMLJAvo46A1D5BIICIc3PSe8dpi/AMxsvuo+SISXKA4ezz2Pj
icL0fgl3DSRu2ybIIjfKTfCKbZsWfDVJgwB1eOUfJlGvb/YiTkQfApdYeXz5
EJo+C5fiHlBTJkMk9dov/Uo+IWgDSm3vOpo5+dG81uTni0WSnEaszL+Lygvi
qJQ4oOzWvSuwX6Ef5YALVziXaC4fb0YxD+7+n2yXTO1Q7vV7F5XnMypcUZ8X
fEhbXlv4AxAjix6VUj8/EldWm13ehIsEYGMAUdoImZJDzzogxjs9UbUNu5m/
Ud0MAOEio/QV8jkVDOb6xbqjNvnbmkFwjq6hbtNM2773zvtwmMW2P0km+dOg
LjCCXIQT6+o6VsVKpYV2GCGncxU1JqUM93gWrvbJ0CSvDSDc3pBlQ63uEobT
swaLOWzs5QOUaR5OvK1Ijz9jx0XO6JZYN/kGkPSWx4XwOGaMHPbdsWlVtxrv
PIqY2vnchI+ipQl99MipMaVwfuRmORr4v8ojNZQh0GUdg8YssYXbr9pSse65
BiA4ohn7yyknwLMXCdzEe4jE6D6/xrusyz4UQf1k3fL/Od/mNbscCRzPcjxv
hEoNGZebdnAeEyeAW7gFokU6cctRYOvAeeA+ghLfH8KS6ByIIuUz0iYd43AT
Z4/UuUstpswXLmTYkec5snb89sYLQsblw3ka98+KzvsSZ+iFBA+TGFLBNdn3
D2XrOZT6/6sbXQ1ruOX6Q+StFBSKy6NwCnNK2Wp6dSJnMtPFgsJp8TO871zg
1oJOS3xn7jdF57dlKRsa5zyEXp99akcPrz6bKcBR2jj/ZmEivTQdBRxlYmyb
kMv8K+RvIzb/EplsQ/E7wzIaOHA6DAo+s+qaNfkY6jIzNsG/bYarFmKNOh7e
7n050pZb/X71O1TAUd5GoiUIgYFgJFpMSOU3Ap7RyTnUAlXvJfte7HQfGL2L
/eLDQAMTKzPoBKjcx7wdni1rkqSHtcU1togfjVtt5DpMVlF3E/NMqengCM1d
ehjrL9N6v0BGQ2auBv+OI+fEywe5xs1AqAv9oJB21gyVSHhayKclg6zoJpB5
z9qZl1TTX6H0oVuYtHmPK5T7DPbuxJS8y3QZ2GHVxYa1R1uTSQfxNWzjVd/t
ymOuiFVFYmL0BQ2ASLuCY1FMDqlLJn6754l7ujyqj2Z2nRBbAhG5vyUkL6ic
7otKs+0uvaTGwugvr2OHQNOqsDocPRRQAbz5ApNH+FzJvt5uf55KgPBTlXnA
xpJZRGy3DgKX/OZnnjKq6CcCl3HDwIqPNNsmoVaouXES0IVdEH2p/FomXhWE
ERBf0cSdNKvoDcQa9F/z7eb6NJ/jqaof5Yl04IzBS9Wd+evwqFY9wRaFZqGQ
euIrnii7Ignk83qvda/qyxlem+5hkk4Wx8ZCAb5aAoYW5MyGkw36kVNT3n8D
6gHVjJMBTh9MKUNvyVjI9S2F6q6GDhWL86jell5NwBIUOqJuH/T8TZz9NuFd
Gzf64rsY00vNzmuAmV4gbFZ3VLYhCj8UPE7PlsxcnTpJ5MY9sc+bfRYHvMoc
+W1Gg2c4eZr0eXsElf9gv4e/oSD1kCbgmpUjrffkPUC0OusjDi26wooIk6eC
L2/1MEOQzZk5g0SX2riVmvQbbIuph1cDcZMbgw+fwrunfn5hzrr77mlPUABv
sQwKkj5b8PRuxxl9HQEuzOxVft9NgdRK1QUDTWU8oxGEccyZ0bMlFYeydrfO
9Mlck1elTDZhm4cQqo91dAwLmb+4s8EfspjJ5f8Q//b7lIOiPjfJNByH4bng
uDHPWFnFI+lra846YMHYEILid4XOEHe7oa3qJ88MmzDkggeHKVxF66ic25hQ
XcMBmqsVG+1GrBEWaTmxWA2pzgfvOx1c7naZG4jNZ/iz6CPxSGW5TIr/CimH
LrUjJEuNMOjjNltESdmKtzRw8DmzGRqt2OsVdBwlwPIFxEHA+0X4rSyiDgAb
DTBiC0GNGifh7aU5jZfglLmTHPjtibWpYHZvZn8wuFbc/fbYwRAczZ8YhFx0
JSf7vLdoONQbaccz+jwEV5vGXnKTwGO3qx5CU0ItAZIAxg7zuAzVsu/TTJec
mfFuL+buHPO9TToNTHlTio3pYEDAGdgpv/Ek/2Oc2kmr/7eBXvVw2NiUcPUS
W32OU9RtNBb6YXqI0PgkUZiihB8BXhriuNklkfVWvPK1ASxEQ3KAsxO0QQmp
uYk6j+Ie2JfEF544+ljGSgHq6J6s4nzM4veula5aCMjL0lcx9UNL9PWfznFo
b1iuDo9KA/r0sP6huPa8tKLI9thFAEQOK30M+D5XR827yj4lxsyrGJNszgFN
bkSrEIVwnoYSuYCDGOpUCxew6eQ/sUoBqLtG6yDxaF+V5URsXmcD9zMnsxYb
VYbwFMweB41s6DOE9/3ajtMV9wAmP6cZKYW5DHJLjc1piFMGdVVkcRboqlNQ
gR/eD2L5uLEEGBI0DBuniAVJqAuMzckz28RSkxYVpsFb3j8vXcOANNKPHABo
M3ElTVJYkfOtmpJGqagQbI97mgpQH4EWkHSWTELzbNC6YnWOwtQHjheepR7u
hbQ94Fv9TCjZo7UnoUF8dP0vFIChKCoEoCInY14ca7Vvrtn9jeaS6cp/3iVi
a/sWC8haUE+BaDH1KwbbKf0Ni2E2cr+xgy3YeU13p0Bd9Lj8nnZLyWro8YDi
zVkHXBlyHQgZer8v4clWs41gWyO36B0Q/KXSs9vG8qn5J85QHPOTuRB2N7sX
4Z9ExWaG4hD8bWK0GovI3DLquFRna3SsVCLLTTAwj9giSLAR4SQRL2CaGOE1
fohI8z2E9P+YyZH0QBxVkUZdq6PnhHt2eznZzhmM+6bYahhbOiBMy5ydc/BT
8T99xRcTfbjK86YrOjIgomyS3nVVO1zcs/HE0aRGvT1YmmchDolj980G5qrn
58W/mhB2wq6ybI3nvKvAeNYbrJHNUHWm6PqIWQP5+dwf5rFXH6unQFIjXIqt
r6pdHAzBTU/UFK02OaEj/ZKLmfH5w49RomhiLyw2rWmf3jicZH5BNCeb2Y15
KLpPu5Xts3up3zphJMK22feVT1ILil4H76b4H2bDBuZxezm7FV+X3KwTxZ0K
TEZArHE5dfwYaBnT/BuoKyIXfsOZxlqXiKYd3hHCXFwdh8OelgDI2cBa/8rc
DZo7aFsUeYJZhT1mrNle+i5J+lax1s1NWQ62/XcEmLjIl2eGbZK7tstqRe6r
7Shev4EssjQl98O/0dVZAuMYCcU9WLcZTLNeOdzGrMduM6LIXCHxEK0hHs9p
0pqa4Mg7CjPdQrbn2AoNhOfpu11+4N/ofisSkQ8d/anJ2j92I+/o1SLOlutL
Dji2pO2ggluGgusi4yg7Rc3NbbSFVLYh7i/MJxZYSJF9jAdX/isleGuQdFD6
e0d31qKmx2E3A9JVaBkUcgI7LQ8ANeb2lojQV7zP6xc7QUGaG41VYkRYjYeR
BqC8Mke8B5a6L2wFO/e+83AcOtss5q7tv9cB6q+WxkakozziPVe0dtsekmKb
O/xHSJSiYpQppDTdVbbOWHIacIY5oNwBkLGIhPsrbdea1rRFMMii4hnEP3mQ
phv3Mz+73IXR6yrbIxnw6nGbZ4azUZCZoFZ+qWdi/GkjiCV0+vq9+xQrgbYq
Uzo8Kb0KRqwB/+m1QmQ+vq/1EcDJXj5vV+OITXJqP/stPp2QpGUGsqUe71jB
XzkSMz/Yc2nolCLeFRFItFojpjFlEN8w7446c16Qiq4XOMmhyEY6Ns74tJg8
q1bvLlHLRncaJXssgpgavmpw2cU5weur7VK/JmSlpEVO2Sk55hfQlordLBJk
xBgsx0qUoaGjTmQzTzrhJyG2YTrJimcKjNJyrUo2rHfPwCPnHZ//NAZ6M965
IutEd+qOFJEWMk1ca6TvmABtVia1IWrPNFUHXc32wXxYtiQ0v0oJFL/ItxxM
Ss6FHoE2FHXb12Py1DZN38mCP9v3nXEc0/1SJWTGOaXzI3n/CJdo+nogXnvG
21PJyv+KLbwURBM0ZJDY43OyDDTf00ltAj8E1VNw0JC7mmmsGC3CZoCw/RBB
GXC5TUS7DRT6yl9LxQdwAqI22jYanFehOXgg5X/ZJgc/qlOTz6D48Llchhi2
5fW69YMKG7gKa6aU0UGxuwY5DA0GDbtg+vwzrjG5Zqj2dJausRUiJsnoEsuI
Jkkf0tJSb0qE7ma0t1/Q20J6Mh+at+BmjL53sLfbZMOcBYtm59rIv82n1m+A
MRsRCtmEJosHS6D856WhSreqGwJeq7WyDQ+rvh9HZsTmmaJrKkNhy4uTCvMe
SJ4i2aYvKPqlBZV0OW/vJjs53xWYKculsh1xAE2NFREXN2k1CIf4Q8k+MG7X
TtDzD3/2Cj6d7MjIbJQTPgwVgVTwgT8S77dVs+mM9xNPVsp07nRES1j+WurO
nHRLt7QqLhx/hKsM/Yp5fLZf1j62j+f6bpZlcTpOX+5QOfYVF5hkh43gT4YF
wgVUW+COAVvVn/5LQp5/lWOwKNyIai8Zo1aY5kW6pgSr6GjzbBvodFG9qNHM
U2OyCGQRkglO+DAG8SX75gf+SjL7Riu4Qh7scPT3MoSJxA2oXU4Io1IQ8QSE
s2w7HxGtD2RjGWLtbKYhX7N3b9YdE6q7ypTtxc7w126XyK/V3OGK6oKTB0da
nSVngBaOumFv2xHtRIy2WRg4XZrYsT6OGi/uEA+g4reoD0hjnVrKCpqg3SPc
Yrr6zJfIZDPN6UsIjDE51wsm5lkHKfLNhTGLXcOBujvQWgDcOl+YvwBLRw0m
ymD7+swTzYLHMXSPJvUljln/f0c8eVPfwLYpJYL8u/j304IBjJZvPvSXkj1t
/7/ZZ8dRJjgP3hdlENrHsjhZ7NS8dB5bGYQ6yQ58xlt6vWR+qV0vt/eV2fKE
cIXDWTd38E6Ayzpdwr7czF/FiUVfkhYQDtJ4rsm0USAvQBpz4hyMsaJMArvI
tla5cBe44x2PNivm/McU3CYTLtey+QPcRAk42dMED0xZrlKXEoyFKIcP81WF
s8c0f2BTtsClQhKIVS1DUj0fHAXkkPPBVNkmn8rSCSFbIYPU4ZYtBWrlcg1Y
9PM3W47NwZDDgByClnhWQLqOCGJ2XVx7bSRg9U4Bf1+ghybb9iZA63Q8WPW5
1CJt1IcvSq4ALLwth1WPrw2VEoeg6LXaKvA7Lo4B21r83bUsHOmBNvEZBezP
taSd0fkdo2bcG9t9DdumcvOyrIAonqNc0NHDxUGUc1GeXZWyj9UifF6ixDNi
TxPN0gr0UwOxb89m7x8Jp3MH+tH02YSFR1Px0/Pu6ll/yIJuB+xIOvmSDR+1
ppENFJwxyof9lqJPEHXLbAi04KP9qdPmSZHDy6iwSKWTn5eLat+VQSHDCYYJ
sqqnR4eLFerYQ0+qj9yjMrR2VRF6orw+09gO12DsH3/IhUR62e1ETqZDMFMo
63cdTm+/ZW5JIlRQ+Om0IlLtxdRGBAjiFyrafyduTca4UUOqZ7ai2R8LLxPs
uKKLCWakkcnP7VMrwZ3IO95mBMH+Z4ueEaaJ+FXeZ8zcewzswaStNkWnG1hC
0DOXxL/vNNo/BsvcOwSnOVFkLbsZX1DKE0HQheTpcYdEgWnoV+fGL/uIQNAW
C5eOVgNZ2TBU40tUSy7rwBBql+HSVfLaDOOCEQqvSJ/SqL3d7J67P4yE5hl0
NTvKHeb00Kg9B3Ef+36DyPMj4c1EVuAvHHjZOMzniGZkZmFxYdJi709KzJZA
vXayPVZR7LBwvVpE6ejvNE3a+RejcBZAkmXq4uLfBrVizjErD3Pnu7XlE2f9
qSW0HqidRFjjaVQYJijq60uXKPAszuAyVj2KJwcvZlqH+IxJUyTEUa/S6F3F
VTkp/i3PjXLhjwkpt8YtSVI9/EtecT74YNHHaiapRAG4JIMQAY6u/Hx1atCQ
doOo7Z6iEfCd9615bLEWtP4glT7GI7A5C5W1sxx24P6O02a8THbiRYuUYUWr
+WYdYOHz+wrHqewH7yI+vpkfzbkS0uIj+sDlVvcHQjR45+XLWRLy10aqimpC
WlV9Yf8VgD53Wbs9KaqEKbM4jMvtstfV+s3xGjp330v47HVIxIiz1E36uBPG
c+qsdICrOcHGVQMQfDJyCSVxWjKhFBQ4t5ULuP+l3tjG4VSfRfQQyykm3ILN
2zTeSG6XuxcfKPCkKIHpVWlEjj8gb38FfIoosuci31t2Tjz1lZp0sCMuB4a/
essmmnICFukMkWB73tGWQDKm9vVIt+CFmUQxMnBKchsxWpFjyBdPMO9K9/zM
/gictdpMvKrHn8U69/JwBTpyGFPHY4qvdTVLo6sxqtEhzc7uxCtWu8Ni65Vr
b+K5A3dqsTzXNMGDhk8gH6/iDc1CVdOREKxCHwjqXOLhbcubJvoHUPtYc+5P
ESDi8YtPRyT6z6tf3wxw9wsZ/2T4SXNkrXuH26qrJIVgMyRxHEKbhpjw3HEt
8cnBr88nVz/T2eZ9awsCcRGq/aDiLBAYkbPzvKnrDw2Ut1PfBPR1N9Y12Q21
flP+EE5745+F1ReGeVtxizFwSrzG3BKt1TNczPVg9Zrg2iBz6j7SjGem40yj
ekRpLHTxpnIwsF63ecwp16ZIdEF+jz3k4gK6o2hG6eE2/HPBpCFprwPFIRv2
uasem1JHexPIezjgItW0eUW0Z36UtQL+3COtA/2ZxBS3Wy2o3M3PKxYZ6bre
KAxRrOOUI9N03E1ckmMz26EvdVWCzh8riqpWuLkoFDq6Pi6bOsL8UeW5x++O
l0nSmoX5/Mn8IOB5N9m6b8qeXN/KxWXsWzB9Q0fyi9jF1fNReCYrDNBaUidO
i/xog0Rn9zsBhqbOucRaVyc+Ynzae+9tXir0jy4He1dpqLloH2eBnX+u5Np+
nEwdTG7vEslIwjVkPJb7G38F3/oiCQg7fSPxYjuZUH7EDix3biXwJ1zLDeZp
du32rf/s5Xp/pRox++OmEP8uXbG9molHGnTZi8o7/efIn4SH21gvKanT8Tsp
ihARLQg3iEon8nNAIu8WT3kHzd42Dy5/4cOB4w/SE4Ja2ZmYYiD3CtxnFOCO
1bTjsvGRngrxJpR1MjiSe9FILE6xn6KYwznv9PbKzzDOTekvrLhIOCUiJKHW
LbClsEmbK4KRSONzXdTLU5Azn+Q+NGjOQuUq1Gg3p+RBhB5YrnygnonQz7eR
vuMxvMwAuym3AKji1THZ56+zYGK82AURVAgmzl0q8jtuX78G8+K69reUmDBO
rxM9hejRs3Fdm+o8bJgYaum4narIy7e0cjihUhomtRaCwCUODaBcTxUBacE3
NrIVBWuW2gJbR+AFuZq9NXiq38By88qIL6lgl0Ol2bZA848AKB6KShrSswY3
IAWMAZdKFEMnv3zmGRnMiZzN+TpVwVvj96yQVoOOb/Utkjulc6hRdCeZYqff
on0Z0WtZJwTq0jg91AUNF+SlhIdp6KX95rr0NFDL5RMR4BGhfC2mS4bXLAJR
z9Wk3fNx1rXTX1FzhIvyq6i6bYPBeJgLQEtYR9gOa6chihfJ83xhyNoneoGN
VRrN9KQP0axgyf07lDA4Rfeyy6oHWWcO3oY+zh76PKW4A8Ue1CKXDJW0NjXr
YxJB6Rrqo4eqwxTmBpZZpBAEDjd5AiDrPaJj6tg0+z5+KcQlxA3d2WRd71u6
BXwPxiQtDql//I6Bs2ku2/jaIOVBXEu1+cECk9TjDVVqg+1u7UcZ18D23Dqn
hew68gcd/91EHFzDe8XsdJG6N/iz/A5ZvpwIeFBi03JdG24c+8Oex8opQIN4
t76WjUo985bH50KQcm5S4XNTGQz8hjqZPDZM+GApamhizHmct0F7vxszKTsM
Vig6lFyQxGjcJ7wC7uKyN1J+jMS/6kYj9miZD0IgFt2mr3BPWLVJjjNXgILn
J1D6zN/SADJJmu0kwpHnE6DiSqNobfMdOEUSE0taiGKzFWqAXQJi8U6ykDn6
4OnRaKmE4nt+7QyF9pAOzcol/9s7fzJE+EDQFTlOOUB/53VV5timbs4XTnEo
agUZh+06ARcQLh45hZo36eoJxk948mVrao9FTtXXHWxDePxiP2XnejWCI1Tc
QxxsiPS01SiniGx50G0p9+L+uKW/jzM36bQJuRC9Deky6jNrEI54UkU7SAo+
apimerA/Ca7f9QFcsY+4A/KBFXy51EjllTh5sELtppUDPIkfrIy83vB2kunq
HSzpK+YgdUp9Zfde+FX3+C2eh7cgs7aVWBGsSk4Vy+ogIGC/Mr35zgEdQGXl
Fi6b+8CgLJh0+vpItqmoLdNkIpMioXHYsC6Y3TeGcuJ7l0jv5YxdH11MwKG+
BtJOUFWOgWUnRZWZWtE3VPsgliXv9u0qpUkGGgJRYeuKQrpSwB40MToNnksY
drgb8cjEriFLvlsSiDOwR+MiktQSyMAzOmv4DwJVVGI9u8cMY7TE2khPKX4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMMWaUsu0UYfOVzqzFDfastA+ZwC7m6jHVAH0D2s3yLv3MenAcvxU3Ja4E+R2P29YPsI1vIujVDWC7PcIQyOBBGUO/qpLxt99RQlIK9ojCLvCxxXwk423nRJ4pIL+u0yKIagWg7NmKqiVQuuhrtE/RyVvsjHYNiEW23Cx/CTeuv+fdfqCMWssm306T2blNAwdEYZa7LhMoBGOkZoaeTFdVeAw5t86sOOkw8yVrMvHxXL74WCBunBEO/syxxvZzNcmeasLBAk8nPcuiwGROh2mVDbFeyb7A6C/BpgVPqLdkDs/raLY53dfqlJlGDkjF4NrieAPpRFEUSd+iLaH6X/Ynr2j53jM/SmXsAp9BQskDUKT3nnHlAwtxWfZWv4D2Vly1pyuAXLHmty5rpO0Fz6Lg2n5aj7XfvcWgERVIake+5H+FFiko/0L4VfBJhChkar37LQ6iBE8inhBusQFkz8uzp0hr5MB2w2RFuTMKpxoTDU23gilzruA1Q4RIpcH2zyrux0TUuP4pGHaleftleZGiUWeyLsrsSsNPY3Q3z1w+PAA4kWby5pq6Y9FApMbtBfKXtMswhrJpCPHnnho6sV4viKiJDouXAfTnuH9ihZ91tXgApfAB38g9gJPnImN1wlZ/tfzhKZHYkXF84BeGyxKiEGXhkVG/aa6ODHOaGqNMEVAh5jgrp69q67wxqTtQCZqmCvGOoQnbmq+J8si6W/i4cRVA09ReKe8MCzd2l3ZJ1D9qD6CTV9cJADdkoTkvtA1AHesMxHlTKluXHJE6Phc2BB"
`endif