// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CaIZXngKntRQtAky3R3ihRz60yYxJ866leEZV4NQj9gL+77Dk6lMrDrfJ97R
xXVJ+AlFUURNFQRUkZI4tPSVvqcdwu/rqdcQQJXql1rxZCAjg8hKQNAH4ihc
b4ORc5zT6/F70vk0wxm9kwf4hGbiZz1KsaUKNHJ4afP8nJoF6glQcYXTing2
Ha/XwWKnA0lruJkmvJcLKFCO2y3bq9zwZffqxeW1A9TcYmacGKcpM20B7Mzh
+MsMNqxgudrH0rCBiQhcK0q6hvbFQcpIzg7o/bu7DKSlr8pjoO56RoVMz7oj
DlAeSwOw663CTkId5Kbgf5sStx6NzICQ810gAA+XhQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aKa/18KmrCNOrvyOyrGCEaDfHQiln6Zmv54mMGeN9YrS/hyQ2rt+2xUm1RyK
Au+OO3fO8/0a8IlKRvRxGhzxZWAsIrDRd0g56/rnemedcWxNayyLPO8pHfGq
wCpiO1/hpmSQJ7W6ZfperoI6P6294hWMCXCOxkBUJUVSRrlIg4MMvnVfzhFb
bznDmscsTA263CUijHy/bhPYSXfCu05SZ6HwUoHyq+KYeUaVQX4gJ4HtiqTn
nuxiJdKgxs24Na1X9M9Ak6OrZvr8NgnHSGBfElTixrAwhznRCUdDxH/UTE9L
JCMFxG71Yc1ESY6dIU69+z890eXzGYh18oUmMbHmZw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aUeeNSsSqpMWYFPiF5KXe5cGqVSjThb3kAk5ECuOB8C9QLogJ0zmPgHOrIY0
wjqhinbDTOS8HqH3Jrm3EGJRDSFU3b8OT6rM5wzb9FxH3XdOv1PT5AMsIi7t
LigyI5+//YTdGu5JWFsFs7IrTdFq8LDopao+u97ns3OB+f5YocuJQYXj76ro
+QJncwOhQcTHXLc76TrL6U6UnAtPSBeU5KEah3P2EgJV+hU96S9XIgNSYn4I
mnzsPdBzXU7xDTpp4ua+PFXlcCuGx6smVKuBlbMH4pB2PdC+TFoXvbyu9NT3
M4EMCMDEewhlsihEB33L8hivcmwFQu/zURA/K1Rung==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K8g5fA3VlPqpJs/RJp5IdUH2ZhD79TNXcTd+ijBfypIDRsJddOw9uAFbW2/V
GPkr2GOZcPGYluaGKVQw3FOs3NkvdG9EvvYbbE+L6LUO8QU69461PwZrKTVz
tEUwwjUnb8p0OJQ5wMAUn+UfF5tZq0s91cu9WqTWvKrgOM0RHHujOCDHJU4y
7TiT3JqZfVu6PcwVJcNNof39gFWO1ysv7BUG9+/xHdH00oVgd89ah3P2Mriw
6bo6FwYrXwTpZ4Sxp3L1L+JnTMSlSKf7H+YiPjZiVGbqC6mdRblE5187g6YK
Isws/7DWfp1bO7j9gXsO/mqy76nKknFDRTaw9QQiqg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EmGP/wVEXxcbufEUO1l4iBtLHzBmGdk0I7PdqkypVzjDHQWdIiL3EoC0GCwc
v6W2Gq+oH68euseRIL9U+a7MPq5KGpR/UD4uUaCAURnpsC/vYv4pDm5AHpZZ
iUmac+g9PEhBN56Fr3oGG5Ys9+4uHuQHoWgh7vMGRRIDxU1/xVw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wotTtx8IgS5vXCvs4tdbBMlRcbkZfIomxqZLgVm/CLCoRbgwA0HXVtsOJNlm
zxlHQC3pTdLSpE/DYlyP/9i6SzJYOggOadIZnWunRi4EqBwmjVqW5AJf8X99
yvlPXvHl7e6oVkj/EzQk6tCKPbMJfuuUQwt4opdMLXZfGAioNSUXYpjiw+8M
osfa6xBdDr8gCqjUeNFB1FgNSCTRYkBpVfTnnm0acPeZW0OgOr2HSIxdxZBl
UQqfe6pz9LxQ8gftxq8yA8uKuUhOncckiMRlWKchWeqjsRSfSJG3sfzrrCaJ
CPW7phaI203v4j2C25+ZcrnJVZsJ0X59zThITEpwOx0sAhHBTaDVh65UrO1V
GGi9JBOIS4+b+UHscw2I+hThSuAP3kwYPl4ZNwzdutgzE10chhUV/zaG1lzt
4XLb8sN5M6XKo2plnPsFVNfp0vuHDJ/tpxkx0w1steIeLCLmmlSoi+96LOZ+
JOizlEvJkqlgh/9KqwuiRFj/oU7tajf7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MpvZctIT2xFTsBRLK/tKsP1pO294eR63kPiOdvDoKQXhrcHVYPP3dmQHctwj
r81U+0urCHtcOQ05bVUaTvZbErHNFXWehFSEWvoxP15YhtWqynsfBmWH9Mr8
/R8NARKdo+Nql132tsIpKgsGXfRE5LjO6vmPROyJd8xP8pU30Js=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nZ6KjHj3ongCPEwHx7D2GcBp1V4NZ2HB/8BPhvkkiV1WIy2xUM1iAgrhR5uL
YjqasSFFVm86SQsMauzJZxh2Qn5cIY/AnAkOqGyoy1X99Gp4WxDwZneVdIvv
y2NqedVjIYk4FwjsGthjJfFYSMD7ddfqrY90j290o5nl03R3yJg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
r2RJqRYYjB0UDtI2BznLqxr5pY8o7pnAhc2/pUBvYJ1sUGXezt0HPAk3mMNJ
WmQRX1mZS2udZs7apc/GHA8Kwii0D7rxhwcR0SFr309g8sW8tMMtLlCviD+5
ZX+e/E7iUcVVuq2IpyE3K/7K1KwhWAN51jzD2822HW+TFLUUQ0e+iUJ1jn/F
8uIC5kNZON0nq/vxhRO5BQK1xm+4rJJ/DkVjbvDbDEaWGKFXYMvFc3cXTyuz
+MvP5wOdlcdbQ4GF3u7NUNJ9H0VDntlDhbqKAkGcrXua96IQ2rNKD+XlM5Ji
EvtIkUNfHZCPMUGgBlgJgeFflQLZR3NhxcKmESKnGP+WifTIWggx8SF9WQmC
OBuUmWnqaNkmAzoO9DSTYIRLbpsnX9l2AVjIR79pG/mFfGv057ejP+wcJjx3
inmZ2d7bjMnTxjFBepwEHJUMNsBvtRXRme4rc849NBLEBfcwlbwaq88+LLcM
WiVKCLEYYkC3W70iz3uFbylGbTqk5o0h5undfoN6m18gEAJ24kKWjGuSqij8
lgSOmphhcoIximJ85mwfKwanbA2MCIlwmEqFno0QnCYfgkfRA+Ua8KPwVnnz
CiTB4FbVxUeJYVCPxfuok/e1bLKByTgBRBIs3ZCcyLZF73Ndy/xP1d0vZRH+
zSGVXFjLouVMD/2LBy3rLWS+aLViwg+awgtUpgDGggyhpXQV9Xsq2wKWRuXJ
D+r21lWBTgM3ugPtxv0S3ch8ctxxA7opINpdg0On4d4sURtj76+mBtdJiG11
TLnyD6E5aoRmsOoySYsk77yIRTkFL2kLhSILCIhe/3O/dSCrxNo3JW0bZw7Z
PkdnxCSAyIxr+9mwZ33E52wE59KdKkIEVpVdBMbqzLHszqlqK4FzqViNMO3i
1D7mag9a0WA4PgwqcLX1KVwOxHU5oK9EFstdR6SKi1c5hJOk63AXTlLW094e
mwLLajiuZNrdGetEtSdMzPkfDleOcUSf7KripkdjECr0nXRvcAfUVXu0Cs+s
77D40anNh+FODNn/Y9pcGve1U2S1iIfA3vVDywo3RzJrmJsvXp8cNXq+gOv1
3qdU8DiG9VfzgiR2MJFTPh44hpDYUR7Z0sNNuaRfHEDvta7BIVFD04S9i9d3
SfL9+ut2LzFEkc0AtXpsqpJOUPbeZ72PyXArQzJMZuryU0cdwGu7uno6qtVl
c/mWFKZfQ/3Cn2WmaSmuX1+UdJOWOS0yXiLb/1uAuAiuH3dkR54CdncAcTqG
03v1Hkr9ShMKzXgEyfPE8AHiL5zPsdAeELHiAj3cSRZZJxQKCX5JbRxPWflz
jr7kTimel0wfedqOLAifI2UrQn9LNfxTZKWe+3DQ84qkpGpTgefkwpJ3R9tl
T0weR+w=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqe4yARYOB5OEnmzjImTv5C4+fN/2wg1HVciR2l9jhOO+OrAWwhCgrWnwrq63V3MaONFxVZfVswCnxaqA4ydqyatUSP/s2MoC/Q6Rss80v9XV1UHdl67Ps1w3POps9duG3fyNjxEqMRkDGDu/oNvP2okXpovUBt9a5jOD7tN4GzeBVFN90Z8b3n0WGqPySPbiH7Di93cnd3EztJDmYWVEUrqBkWxcj9j4rrlBmOB4hG7YfpUbf3BgORkz/uR6e0L2RL6kWkCr5kxY0KiGBBiDI1OlgEgy1/ocldjyDfL7w1qgqusG0ZjDNe+qMPRwCIwMALzs49zAl45mcV2JaOlApaL6iXAGVGgmAgN/i0gHjdynF4zBdTuZe5KoV5ToPpGyBZwPzMT3GLQMuT8u5xDmas/wE7uzHC1wWfIuoo+PI6C0kC09EDyEtadAsjqD/w+jSv8fupGLjO1jO6mYRq8JeSttATl66fKOxR3/kNnuvDPc1qxx59QhXJUxMueLLV63Gk9WPAb5EYLDoVk09m7UNtkGxgtVi9w9SrGesiiobVt76TJdRjO16rKNuv5S2xBrUoLyQm9E05JTQGlRD8fUl3VVtgYQo/xWPZ0x94xe75DW1rIkbMbbSMEGpzHIHLOyfQs9GBsZr0K78ezzsq6eEOvz3Z6DU7XCNMRDoSPHY7Eri1KKgnKctHPfnyJ8HC7/vga4OcQVZ1Clggu+Ln4jExCVyacgH9OjvA8+yaWCbjePluFluhkOyW6ScLmCMi+nrshqyp8tQvR0Ir1jyfy8CGU"
`endif