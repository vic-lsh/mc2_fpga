// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tw2HEnRKBW+w4cAkpuVzMzIkQgIEJeQ8aakra/9w0j+Ut/92Y8wrhv7mN342
sQK1NxRJeerKFsObs4w+V8r3mqcI0Y1PfcN05Th+6Rd+xjBvtd/HM7TOwRMD
AHrgBN6lEr02UB4gUbCnv5XLUCWHf7fxqTFd+F0PmqoD9MfxDQd4hAU5MG0J
M8QPYRsZ5B7u7/RwWVwzUKwDV1wuGW6uDYtacD63NkilW3jzpxn7cplE2fh9
8WYowAlkNdiPx9kxD9wASfU0m5kAuzsk4FM3ug8j8djUOiEgHT9Q1Mi5+d8s
p1K5Ski5xgyqCSk+RujqHFDHHyv6wd8QWHI+hy9J5A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dWf26OKzGARNiEBuLBhksVOCfBnfzLkjPL15R8KP5ZitvSwzDNol3w2TtH5X
tWXRHGWZte0YPUX8Z6QH8aLVU/9P4srRqPaTPtlNXKP9asrb1Ipr69ioM9ji
LTyLWGvzaJ/cToLdgKoxjzCT8KfT4mPJ9VPFokqo5TlKAG22j5IdKo/hz03A
KX/t1xaE8tA9LwK4WBE0MvAZ283aJnZ+TVHU2UYNwKdNnMNixUc2scwmIaHp
WriYuT0uTNswZgeAtKcsW3pXQVUvnKI3HUHzvgLgLsQorR0NPeVNrZ9jkbZu
VuZZyWJfulAJd1wYJzuy8isEBT/7ZgtQ9i3z0k/uwA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sKgxJplWILJ6RgxUuEW/KQf76L8SudfIjkjWIMoBHFYeDE1JX+LRE7hF2Mld
8QUJlYIfZSxN9xNZVm48UD+IyQ/21B26AnvOZyNKRrSuxJkrmK7Hp7xePfxi
wb7IsJEanEZm0TdtvmBKFQrDxmOppSZAyirJsEJsbbaBAOvSjvKCDpvgPqeK
O1BkcokGV8YLNMLbGiq8QAXPDAEvR9iPnAAfs2ksJPt+PE8ULJkZDzfTxBaC
uRaRnCbReKxCOC6wO5D5zhUTXHMlXvQvRCw32rOSyL0UuuB8oNUJeIYsIIJo
1MowMcaOXAVnjyUbCLD2DC039rZYeFXi7dnFpbgVxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IZybrEzjbp+O1msUgL35OtNs1KrlApKAF8SAZLrj3EDxec0WsDvxSptm+9lf
bM3v9HV83CRsW8vonBszSDggvo7+QJEicaAXpAInTgBOQLpv4x2nSIzKKXDV
JiVh2PEUCEYmbv5pzhNXSfflxr8Je9mPFDAQFjdfaTF1ZFryK/ccFt0ZWK8l
B/xRPTh1ytJ4aSAeNIcFt2NZ34Sv2qMreQ3LPqS+gfas3uI25ZBhxIk+fJmT
qxKlrgRXrvE3/+f1nv4M1oQ4zhL4AO1jdzYl2bbP7cz2SbUjyGpdMi5XYYAa
FbbIB7vnkhgan2j6ktsUrfHD0cfF+JCXEG2BDmrsjw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nTih16bl+O+CHULXDaRV9w/vRSSc6HHKEH3gzCoZ9SgEz/oW664f+W4bWya9
Lz2iFkHskx26RD/2CwTo+S22pwYDFyAdY66wLxL3ORn30gViUNDGvQCz7gKS
W7ocAk4HMGz8trVeiieelBYljSP/7YP+VMyfYogN5HpJaaWA6AE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XvFTaDuecuXqGGi9RV2kE2rrCOacyO7DfhOUDlZdKLyAZTFn05waiqa7S8Hu
nQSrMP+I0Ixjms8+iJUv45sWQ8pjVnhJMBAYnUwgmE8h4zs6UiPnGKK0CQlQ
BVIUsbfaauCyl/ffRCe9g7L3R+8bKXTwRI87MRruLcNueSM+esLCMpiWDMve
yCyHNJ5toFAD4Ztsrff4J5MoXgFquMHFEzZRU/pUGRS1Dk2E16z1zilmnN3M
KxkPf4XvFly7vQZihSWqekqZ0lG4yQ5PBhIDOD7WnMbmGCz8tGPnDFmAyiyX
06s4fmmz6Qie1SvcnpBwx+Ybzjvjc88XolyS8leb7zn/+kcrWZtd+ZYFqpm4
Bo8HVuav1rHaEWlMWDh1ODapIlIxBvHOQz8Pc2RtOOnkt5/9GvWazRrLhub9
Tyh6Kl17oirXoAkAttFr+r4hV0D7xQGBr8fH+ZQXbWviVmEGE9Z12wFoyzKT
X/1ZWO2Bvp3Ku/4KVkW6ovZAL3EFoOVy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q/fBaWh/SuJud1l0odHEdMZHpADkfJG+9jFU7fhDFVeaAWkUm07G25EPO/nD
1v37gZMmG5eRv9i9OKOP6NGJM/LYnPE8Ldv/pzEkX0XB8abH8PeuHyzT8yuG
hki7EBFuzMaEh07AcArUUNDxwKkPBuCCFy1KIizZzrBdlvJtWCY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AAWtRFKOjL6inlMmeFUxOjjYX+i0ms+WhcGhVR1k1N99dIXCgg829gIPJ60N
Axds6F4kBVfHSlgby149tbi6XnDh+l9cWrjTEKhEWn4i6Fv0+zTTaEB9z4kF
zPnf6w0TYUvqRlUrqXlHpYJDiWiPxYZafnp0LjSvHdvylhv6oR4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 34352)
`pragma protect data_block
lpiybYGulHrC39JFjepM02mEZk5offm8IUBoW9CBPJSra1xGk7c+1o0N1Skk
J928tt5ZnrFvCgy1UVYnTBB943rg8jhHBKruVqrqqw/SnQIPPpywzcu7lwVp
VrE3Er89uSKy5F2f8cWa+VvDBoNh52rn6VWtwj4D9qS52qtDt7s9nYYIFeM1
Y2LwV05QHnqrIyy6CqiJIkostyODt0WOKvvB8z0pBKeevLLOspzRIdPUkWDv
YOm9F2dXVlHRf6i8MGTL0EUjeINkTa1n5zJ1VD1dvE4MjoGa7Vdw3CiI+oly
s10TJ3xO5wwx/BjdE08NALHTYwmiktdDIPnyyf2mA7Xs2JbfgyxsMkPmjaru
Wgj+iiWBFQZ6ldnF8dO8QODId/nKbMDhJ2KGiilY6RYNOblg5bM6AAk3b+eE
eCZJJYfewidngticaMsxbunL11Vs24GGGxcykKJVphtncw5I80HmPY21U79b
L752BKEXHVZHhgBGBjyWT4rVENmlgWm4XKDpUCfqC4lAVkYxEYI2L6/Sh5cG
4ycn2F/me/B1M1I3x5VOvpoBOoH/kb2Q2GXouiKktlIXa6CO557jexU7Kvik
O1IMR6o08pJEb7+9s4dfap6NCdW4K4zMoVJ1GgXxLXrHcxIHRDAX6SQ8ASgq
o7Eh5hrSFgytBSJCXrCiOKc+RimaCi6HztQInHV1OnwN3NIJ9iaufg+3ZN8q
slENPiDVqWs6JTrPg4S/KimXJh9ZTMZu6nLwc42P4vr5y+QJXafxLQKh1Mlq
5gXo66x6B+4DA03N9RrBMSp+d6RRG1ONowYOXutgBMhVkC7S5ssT0IGmOSlM
WPgNbDcttgf9pnxbYV3nHffRjCMnef9/C3FeI/enhdzgCuBVMfqf0bZ4C4iX
YNGhFH6CaF37NmngS11w3+BTVpFQA7ES/UnfdQ1VhdHn/gPZeZycHYFik1q6
jNxwb4sL3S71Dh/CzkYtgyUXkxJ/NTqJ6cUUitbhQzwlWGtjnuePjR2ZHSUo
QlFT5MRWG/8u9pAb5DT/yzJVf3cslaC//kup8G6QvOBBUKGoeyIbZOpHaZmw
yJ/iRVzmPoje5+bQfPT+vsEDfaZZk8yvYQlSVVd/VFfTe3ufDIkMwrB7N0OB
/OM+x7K0WAbrJjgNLrrUlcHrKYnRlVum7G9xOAbaJSL3Abc/w5Bv4/opflvW
SGY9bsNd/IrmAEMb46+fvrfUYcXoRKGTifot2qLXbJmXcRB4QM3p+h5mt2TB
6FJUFeV3jNmEZAERqJWKVKT+LM6QgugX9v6Bmci+T8ernXOLVKX9e/jmEWCJ
TqXtx4n2bQ5bceL/6ARj340esT0EDsGq5zODegBYmzJ0hFqdOj7gsThjAEUr
4/ltEikghsp8zLGwQbOMyrXSdlu5F7u+IzAF2NLssKBTvG4nFK59LbzrUu6y
JfgqalR8tnq6hg7v7oOAyc8WV67y9M7430d1vaknRjqL8NMTK0daoZstmci1
AS/QSdf9jHRM8a5ZYqNoZM9BwJQmdo5RMDzRzkSl3Gtz54p8lRdlnocyzNrq
d7/qRb3pAKYCK2xxEUhcldmySAjtbT7/CitoMhTJs/Nsepa2muLFBBcwaq+U
qphdvV+GiL0c24C/bANo/5aWanzGn/+J4+Z6C5mxKcVVv7AYXwbAA3yJSCoK
A6srQk/tI9VhlSxR98gGHWCDk5dScg6prQMeNMEq3LldUbFixKeTNQ8iHgAV
vVtokonidkilU7bzBUqEQ3CTYFwpAB6XD+Tj23j1aQXHjcD0ZtqmKc2kSr6s
IHldhmpMvx7nvYWvQBpRaK8s11rCPeTzgfPUDVPPZtaQTOfwbREIL4d+EhyX
sk9HUkOiOh1d1ZIFjmod4+8n8edlCVaNxSJblwJGeXUCGUMGPUe+sfNBKhUP
adY6TbK9SVhMiq5Z+GLnXwi+cKxUvAGH9+9fZqcV5Sld6umJ+PM31U7QA+/L
mmIUHtVItWyTPdblQeH4X+9l8mJI2PkBhaJ0K680yhjq34MnZwR125HQ3SUV
o7przYfj9OS8z+9UgxEjUUAT4xdCDZjR3sRHtCdL/QM0oC0GKOXHlr06Xex8
T1tOaSfzF835q/eOfpXZ3wyUwjJj1/QDh6EQdxshr08j679Quak5JpL5x1Mi
O3Fvdgf76q+AC1r1WUZO+y9BSb7onHmAnKWLl1PnUlKgEbKKZtuCEO4Aiz8f
/beWD2E2XRKbaUviOijGeWUJH3xPpJ7LzOqheT19yWnqcCn6L2A6WRLNz6Fl
r9cTMncdvZJWyxNsPk45ECoNCrfL1x0ASyUtKTWdS5OVpU7SRe3pGJXskP4b
HJa27M5ysRMQ44o1X35OckIMZSn3LSUVPDnAaMJMtM3OTaXEQrKQRyHlDR2W
zfnVrtgQ8P0Y+rWcdtErnEE4xOX81VDhqmvXbcCWo5E/AyYe5KB9/bt4E19z
2msPZ6duzpPjKI2gF9VVQRtHGU7CkIT+mByFJxgTKwYsh6tq9+VzmkpejwGy
OCTcJWfOUxYZfe80ekKO+3NqGSCvLp87p9Jk1VCbwmDDCCq2pmVAxr0A+sdZ
eE+czHG4ciVGR9m6iVdshpdHu2f2sVGow9Qs5NXgLAmSd7VV49t4lO/HHqp4
ksCFxfYrRFa5DjTs2FzFJYEF+JI5CYrIeRLU+KaHqboTYe/Q8TGaMtpJnOn6
FHIY2ms0kQ/J63S/6QY9b9/4IuJFxnV9PWkIDoK09i6fE0J33WFdOmItUQYa
mmsH/4MPkIl2AiVvq7vXTsXx2MFRqE86gUS2s/GTtaPp0U8o5Dr9gJulbZqX
6KAHJ3mXayfB2izeyiK47oCs5dfjUqpaM9A1KmHnriOUJvI8kb5eYeBMUucl
Rq/aJu5y5dXasllDHNex9a9kxHepEAshmsZ9Lkw5F8wG05ObIGTm+rbgq3cj
OrN4vLo8/kTqRWcJvsR09rK0O3Z30KZ64Umy3M7PmOQ1edmFwXbyzVJwEqxp
ovv+r//8eBLncRUAJ8je9P7DuZYqyDvcipbcIfUwXsYugf+E/LZK0FEVNAk3
XgxwtWjdj2r5w+UcLoTJeRrpPhzD9PTvUqBzpsCl9Q2T+RwEG94gka25YDTt
nSDWUjC6qrr7X/2zh+TkRXIVuz3/KD6qIuIiX4Xu46aLsbws6QyFFIEUDHFc
ZzZW6DAAOnr5ZIb6LHzzrGRrXldG3kCKGFk8+0t1ajJIfDDAZgTkoPi8k2cG
v0BmVZUPvR5ay3Ce8h3OcNJVXRmyKaDcwFBlT3BVIkawb5dPdBzD2ThDNc6y
iaLSCC7OysZ6CWRP6pXc1bv7Ngk5zsZ82VQx1g+1h7UVqexayN8Xe2DnfaPw
5syURpFa6sYAQ807hrVF1USSwryvh9t9vzGS/EjbZ5Euvl0L5lwzgMSY2SVp
jhbbHFJq+B69ZR5MUfmZxpwf3YHchjRdYdRvrWGSxAU6cd/3fbgIGR8WXw/Z
E1Xqv8mH9hPqhjFxdwBMtytvV67GdLHzyURiJcuUTK5CFWyqljlcMkaimlrN
8Cr8JDo+nY10vxix/VfMNUCx0eAi7oRM9+ha2Ftw71H4vDTDxpuJ575wHX6b
cYqUNa9FL3f3b0BxbcF/Lg9F79DvkpAHEsckvXux0tdjYjTCc0xTXqdeai3x
pMxtCSk7cDOR8iG0DibxxZGE4EznS8nL2R4t/WCk1o/BzGBu1/izrrV5LyOc
a4/YTOenzBW/o2eXasvBmo1i9PNp1VnXOZV84n7x3syDSfE1BVEPqOxiRIMt
z6RNhRqYH0R6K33hhNXkI/XH7rZEegkr8Ja3cap9k52dIk1nsMbXFWYHSzTq
O7VhgJ0/IiUWSNjr71YD5jf11wYtWfr55W7C25ZDrSk2M0W5QKbMDyB+hXhM
Xw2vltMeLz7X153RWDuUhOZJL2SC+C5RxzST/0MCNy7jGFUvImyIholdldqe
aLVKTBH78PJpacS6sEQ6aiAyfcm+kbYFqUqwCAaAE/wBx8aE32YCtO4kl5ON
BrefiavIvMW503B+f6mkNuzev0kwW42O2skWCXVCiJhfJuUSyOYcSnmq29ZJ
SR97KOx+MKn4OxWpMGr4+NF45PZmg2nF1pi1EJa/Yt6Mle/MoK980fuBt6i+
h8k4dMZ98dYUA6ku93MVGLAsYiqf42RLhlfCdiLopSBw2LMzFW+kJe8gkk4T
Mw5PeTuMe8UirGTLr1d9E8BGWbH++q3iiak3lCJNe32M4Z85BTiCDKXWQJrH
CSO0MoB/Ah7WEpu34J9GiANuP8tSZ1CH28Ag0eaMUdR4quHQV6fmxPFQ0dQ5
bbJzRf0oVitJ9p+/WllaP+XdVotkEgN879qTL8PRP6J5XcCSDaFJJlS4575f
PS9cbgtTwxOWX6hVRVCYiKzPN0hJnL8Rz97qxJXy804oz6v81JFj/oFOozOQ
ceIkqmB4hpmI+jXhtM0yCrKyPXMllMpj5kAJ6XY1fqr2BEl9KmtaDuJfpxOw
BjViBuWHBxJjqeT2CAJk2WZ3t0Ce/BqPHMyo+LdogZP6xpbwt7Qv7sqDXZV0
TJyP9eU2zOkjRIhtpR7y4RYspdSdWhvunJBdYmTt9eAYHPD1E5vKjL2Kk4R/
QFGHNvVeZGbQP4wqQr5M98AIL45DQVwC3ORT27WS2JNXDowi3u6nhyWyqx6P
ebb2SzAhRhSHsK1mzwxsEpVzWlnwWyNHWup66EDw+VNzOjczuTgyiBFk9Cgp
EI7adc1+nxCiLpqke51/fN0C1CbFRcHxvOKpSKDzF3NWtSfnYrIjVoNvDQWh
bfehX5s0mkKdw/Cddnoh4tvcqQXsXRXuqVZFwV3+cRilz3s+/PTlX5b5d7rv
AKhnx00t9aIjxPKwIE0+stiBG13GDq30YMQgzXHkVdKwUoq+rcdrSKegYl6d
rSF4TQFdCa3XJYbo4Vp+TO/Ye1VfKIrKeqHQj3Dd9EM5bBLV9ngFvUJHq4vQ
Eoor1ay9qcCprqeJFxN/yZvSdXZvOYRJSrDUdDGVL+ywEflAOsj+k+kE1yq1
GZmQ+6Gd4IjyLhtHhCfZbFTcOOrE/0ljc9ZLqdOGXmgCqg6/dKRqLITuRtA1
/EuJlzWS2eq+JGK1+0nrIA1vh+e66PMXwyZXEzsQJsjQqj1g/jTN7PWOyyHO
6dQ/+mzDzZA1pqfyDh/KZT80x0XzAQMpsxgrlCfIlh3Ze+CY7qxZ/q6KprVY
U715YnTFECUY9JPu5hgm18co2v5E3ljjPKQBXfzRyr2HhgYHPPN/p+qE+W2D
XLpQ7mYCZ+qRmOTL8XpcaJBrFf6M6xnCO4Rz0l3i6xuZ4esqVxUgbzjP9Bxf
y/XsTxncYe62x+C1T5lIsxr1JpOR8zdGG0pq2o6gLB3i4+boiEEoVEbfOfP+
kcWMiSn1Msp/Qd+Uzr737P3m7j1nnXnnntbFetRDs1bE8R3hCGGMs2ciYVMk
+OJlkHLzzaMfTx8NASz2VHZTcDM2CBHKvTN10wdexc/n4elTlWy+hlBj+tYw
uPhrriLCH82aUiHceOLApMtAV/5AyfZOdRqhPZ7mFesG5ZU9VTBKJwClMlzj
NOaf95PGbBzRPRfOcTNMyzO2obs3uSi3YCa8yyWTXYPoOmgazM1f8kquSEhR
eMUv6oXDV0PWTf2w6jbcqOH6LIJdt1PXlXWl3CYW2ph4eIzSpBK82Xldbdai
ZPYEwcwV1JSklvgZ3OkdBGu6TfUUfeseiv87SoPn5QZPKrSPjp2TWctxY4yM
Xv9011DYZvPmg6AG7mtwD2iiHLZxt1rtKJVbZTKn2jj+rsrdCQ7J6Fku4eLW
U3Biu6Q2fSkWboIsfNEfxJTUTwGlCgGSIgqRQBZimhhHVcas6d84A0zKbOwL
/txhm/Fgnz2uPgadIxBpf339mPi14AD8oVH/V9BZIofJjXVa16mzuLpT99p6
cYRWNFJ2dD51yOyPZiM/r82KN1H92K1V3U9/NmDGzEz1qvMMWKz9G6P81SQK
qFL66ryPK/pjiZEHF6Oqg2YrOGNF1BRQJsgbMLmzOhlBRaEpW14lcQiONadv
aXLS1u/6F3BWgb/z0KkHJq2DNAA5RwXzWSrxXpWOSIzCZsX0H8rwaqMyRFZ1
DI7wNJBRzFF+zWK+MpvILk65/25HXx9eb1XtKzzGP3YTaWh44JqQbnyWI5H9
VZ2DnKcfykCX2v7cNXPPKFjTRcrJShwesE+SXR44LdMLJ6+D4c5Tb+XSp8B/
akM1vKG7XuSATeYqIqarKb8LRTtvEdAOwfamFzUsNkCliAQSuTdDt0N0R5Hv
jgU9eHynfgybCQi7Aiy/SIuwcS4ByYOdgeTz07GrpXTKI9b01n7y1jPzU8El
qZRELE2FGm94rm7+FfUJjtvj6niPK1A+lNqAMU6Xa+ejD1Y2SCiNvGbUYCV9
sN+Pgb/voisoW7+TOtiBfP56hxV1NjkwOyKs5SHLTTp5Wrfs8qgwWuGBvNjR
mXwJGoj5z2exMLNmyBnn+2c+bzr04VLnQpf39XFXcHBpEij2BPXj/8ug1fd9
Nk5DCBBiOtG8BImKfLodiMTRaCYDs3PZVTNOynCzkdczzqN4ApCjvR8gFFLA
Akl4T1Axyd7KZ4iBK0noEvb1x10O4toedJOGR7jsGd9qUVf2Yo2LeU5YHuWy
RB0zumnR8DrOngn15sl1bD6VVkzk8b/9LPU+KRxqRf5Y43+PQxy0sOUHUlcC
3EWJHcvWoQObB2FwctRZIXo0KT/8OJNRMLwEOfqidqYtqv4ZW9ZuMQvCk7o2
sJlm7GtZCUuOG1+E17BsjsN+BS96dHtaIXSmefT5Fsx/s9ln3Tge9Qdq6EE4
uxb+Zdrno/7Yyd+Xz+Vpnhg4+hGYLn57jewo0CeeK9SmGvhCxY78F3uv1rNz
23JQBssLkcLZTCBTboTFXPghxHdXYBAnAI+5I4Fi021Ix+Jc8QPCou1ohBtT
DH7I6oJYUm4IhXeUmC2sgJHrFGGWLr40Ty2DoaAjj7RZ0afJyQc1zX+vgrm8
MtizMGsAs3MZzZBIBNlhXGyVqw8VxFwT6wFoHGLRAqk5IJ7ODXYoUY0/Ccyv
Yj2clgUkhWCk9qwJdSy6ikcHW3jZ6XApA1ZakJm1bDJ6CPSZz7fkg94us6l0
BZgnAEvTq4IoHWQlT66pbbrWDm5RURhGl3IwZoFeD0trXUGsC/3cI4d3uCv8
649wVNR6Yz6Nqwf9+VJ8rSuc66RZRRvvlRu+WioAqC9Ow9tHy0tSVY4Hw1N/
g4yk5GiPwcJ1nfPna6LONEN0KBgVy/72tr6mlLUI8Fl/8UUPqeMPK5UUCPT+
tkTXWXxYj2IOZb6LiIgkVycahDAP4Ekf+D5mL8MTHVCzNoJv3+M0w1by9vZn
KJ7fzlas/sj6zAfN+zxjVomQGkXRZg3N/+U5ysqmBQFNw7+6GWmndmj5f+k8
tPOJdAN9B3coOtz7uULx9gqJz5H25PMA0TxfJvXJ8iveQHwTkFr/iNcQCx7Q
RV9saylu4i47PV4ibKXJNlf8PaqXB2O6u9AcoBFBTf8pjNYJ0U9uZyn2hlXq
XhaaQp9wzlegg5yMnbOacEc73Lrf0/dxJL5/EOHrV2Fx4ngVPYzHY0wjjmWw
LNLGHA2PcNomRXsvhwJfRPPLaR1/RtZPzJkFmxCIXF6CN71vIXdIkxEY5T3N
00j4F22MZXC8Q11/k8e5WnlDiJnlKZin8ZxVbCTgPPVSQN6l1SCT2NMZ/Ibc
V6AnKeNAx5H+9gBmqQw1hDE0deih9afvPwag4Y/svAqnAGnu6i0Jdg7E4+Ng
pLdMicmM0s4BGgQecmCIsr3jGBprawgk6m+PFKYWPj9iNnNikqOKlTWBQ8LK
DM+2GUbDuBpCFvXXc5q4FcMD5GElONKR2GJJas24yo+zKwI1W2Ny+Ak0MEkl
h7N2WFxC1iWjzsrARodvJn6/iq3sJKwYFNH6RV4Bp+9+EsTuZZs85vltBve+
p9E12bA4zQSh0lA3n5GsSf6Zy8F8mrWB8neEmVxU/5rDBOiOpM8BI52hobul
SIshxsHISS33AjdMfGb6SrsA0HdhyzmI0B7kNaD2HSlQiOIulg63u1psj2Ya
geN7rx96zVtlepWqcHt+XP8EDe7RxX3k8pa8gFsgrnMfUkDtpnJ0bJkZysHa
hbb9BpTqzYLZ2/msgeLUJvibBKUyKPvJpgbqyoU7UBniPzBPOOKN7uCSRkPc
U96Vo89Sp8xKgEYBYrap121s0k5O3WQfc8dhfNbLPP+LAFqUV9wsVMbXiG48
bkbM9NctPFeKdqXk6uGTy+0BLSUlWVHIJyTCqdYQUno6ITpg/JGr5KQc9q13
a7Fq0GFy0BrXdptPmwriqPITya98KmHTZ0JlnHVQzmsE2y0DwmuRWedoPqDa
183NoPogfsK+zT7UjwL8FA0ox/7nyFq23aPgIewobFjlINKVQ4fb2XxTBEZo
X71V69vaPrETrpjNHzeQZ0hExdrNC+vdW4P2aqfcY0s0zk9wY5xdB9kKK+6+
LW8n9FgXGwik3gB8ciwDvAyDawAmNF0AxxTXeYd0FuK3GjGbqc6yHnLoojEd
MNcbt1+cBPiGY3Daikft9H/GsD9HapLssSw7JMiDqRS+uJGa5avrOFk8W0q8
PHI5tZ2L0MvrUExV9sFsepef213OSv8apS7XRTIqeoMPRQbAuNdLFaJOmb4O
XS64KwozKV3VH6861bNiift99zJ+W6B6bCq4YN+f9mbzA0rf/SezxfpanwQ1
2LHxKZWl2L73E09ILQjXY8+GtIh6pqtoky8vP0Zo8jUD/rCvNjvEROmsiJSY
h9K2NUQGMzWY1laNlgLCAM0zZfrsjHtnWfkjBsw4086YXSjhJ6RDPyMydKj1
JJrynD0sJaN7srKoAO2p3TflRky7RiwM4/kX9B+pxF0rZ0zCqIsM/3HPsq2b
gaZvT1ox9x40W0iApGjczk4rw/vttjyt1+9yWAIcwLXiPPVybyxJc+bTUaph
jowuSEzYpq8jwO6xvk3cX9H/124NAt6kGNi42wLkyBm+zoI6jn7Gh+xRzR9V
pbhuYd/EzqfDPW1jM2Eg+4q63fiOCQ+q2BXuIue0OaPOL0CjBpUzoyRADHE8
r4jSZuQ/OfZXBTd20BZQvZC0pj7FHQeN6Qn0QAAnaqYqeQmn6K2QckpNq08u
oyitJ165ug70WCnGqobJm1t/J7ExMKUMnw0zKeGk5gXTHVLQHt19vdGeH7cD
yshIjXuEzTMLbvJuM1UL7xmjcJUtBjppNDDbpT3EV9co4+cSE1yLKvW8X82s
+RBsvEDzfBIugkHcrPEF5zIR7gatIlLN0nc8TgplDFqkraY3eXOI+iaUKFg1
eauEJkgDPLzsb2FQeTgXGbZjTYiwy8SYWRKyhC6gSRAV+xMtoUZotD6kxYZB
8yuDsS78ogov6NiYvh90XjPYb//GE0doOKcQs08zP4yUKKozA0mIoNFOpix7
QAgHb4cGHAjKWYxtaDU8/pSBXRRBz2JnKriaubcynKnLrIBhP71vCF83qktK
ldvOrpWIt3paCFvW8s9vtWragevc4qjkx0DZ++eZhSXg/+P09/VczoWIhM62
lrII7XXNVI+nk2kre2OTURHuAii9S7IyAN6dvB2+mC+ZoXGoKTbyfACVpPtV
myczsFL2cu4OYpMgAWqDP2mMDx+SpA4vWRoB5JlH+JAwiDplDvGWNChwDjvj
mjJh/x5ixvZIVZeTJgNr/hUpI2JqMSWlZtjiEZ+FC5x4tnYddqnVcOdIgG9A
n0x5PncL1sN0mDcK0IXx3yXm4BG6DTosxmK2OLDebzixHY0a3hS8y3t2L3EK
AdTP5Vpa/4mEPHeW6fuBThkS0W8r/SOzl+9yKs6cNudfHIZbt1IRRukC3b1N
4nKKg5hHlRV2VKCCPsHg6/4EzLxRusSueuW3Ex9M/7kk7IuVlqe1GFpY9VV4
og57w4vujwzRG+rvh6r+n0EV4XBSbCCVvxYuLHDtGo1ZBlWUlE3CSDAR4tCP
EBGSzy8wjlXiwrKpU99cQAa4t1qdpLBGHc/NWV3nDuL4ph6g35saSGATTsw+
5paruMLOirl9JN8Io2fzdEOjX9w9LVOAn9SXTKBJ2FTPQgOFS3GCSBTVkH/P
sGoEhVSkaQ8RgTKlcQsFAOpaVubwwNMzCak1CiMgdXD7sXwm4dpVDzphujD6
8h1yjuAJAGRG1nb+h53TZmBBsrDdcUMZjUEJh3inqIsz1pzs3WP5DSBW4ct8
zu3WIt343oK6BevKsmJiLa+neMyxQRGq4NSuRkugN6DNEPpNFut3nXktFBs2
fGqTEcXMYhh/yjkLYyNJoDsNwk27emkJRergR0MyCdMqxSYJ5+e1j2zDqOJa
RkZMI7SfcAVcu/M0vlahHkK9raaHYePO3jzYUivgp2wA9PIFxqXioFDA7Mvi
v8Y7sg0xk400ok5KP+3QuETzDiz4c6ObLBQeNmToCDc4XQnMxBvgaDfK6YzY
a6LribAuKAQ8YQe//6LJM5xSlvyptmyYA5QuPdcADikRB5NzI6KpImxF5M+a
l3z+c+Fsd+jFFGPvsZx0ztBQHsQxPz+N/t0HESsltsqk98lNIvD5A8THX+bL
dy2vBAt1/mHKk86TC51+rtCnTnVdKUBzTynBgikSftSYDsRRIsaffbws2OMV
p5ZD1oXAHpOTxcEOVxKCHMBKg6i9FeprKMbq+xGmvrN3RfqdP6GKDFSMflbT
2C3x8MZVoPSnaDvm4PHg2HgXqNIObnEPat0uU6kqeHer8VCJBGecB+csiq3C
TQy62iBNEGOpNbsjMtM8+Oo+NfkWtZklDtVv1HZtLWrKgIchPrlqY4HJXrr9
m4vXnoWBnWpyDB8C6EywH6tHHSw3xO5o9Ki6TiCo9zoQ7WHVFamAPL3U1cwb
GKiB1xMXBYKVr38uFTsTSe1n7fKKWLpv7dAEgou3oYpwE1uxUnUR3YGG7qVN
/rMgpByAguuPxtfm8D8S5veLheUuOyP63L6QIv0WiPSxkP0r80OQb5CprBfY
2KHVPokD0t8kNX8W7eYJsm2B7Hg9i7Jn1BmQD/r64XMW8OV0HVyzOQzgKJY2
ZpnMQPxUA/ve+ODXeBwIQ5k1Ym6QlD/K42vlSlKG79YWLr/lor3w6wJFYBGg
j6GbBwCkMsBdD+7GzSGVyF2R0l7oPlZ0vjU3VDiEWiYGCNQ7UkblTgkBcPRN
/X1TTkvg2V3npc/rIBEuSY8TjAIm2v/plR45dnkLlAIoIdwkqcMyhypIim2n
ZKYAdsoKs+KPh06UIIO4h+7vL/RDdU6iQbtRP73hICDVGzPLGI/1Gx1sEqHF
UPV3U88wkYlEv0GpAJnVK7oW2CYXebKMcGLX2aENYT5NzHdk0puoHRMPsOf/
6q0j0UEUeGKjkTNmVk6HVQ6IL/a9vVPMmzx3HXOjVhDVDfR15uo9QgC/lJvz
XR4HRsDtw+AW47Niu+56zjcvTLuJD2Mb1kPVwvvjOyrpMAjYY0Dnl54Cp86Q
+Bohkb16xcePUnG7NT6xnV8uiwYjyxtEmdXU5XrzzDfOP46GIHiWdWsTyYRB
m7/W2plUj/uwwTHFLSJ8hcXYgAQCo+YSPQL1ZKIFEZyRD4fq15FrHq2smPTt
BwEcG4z6472WmPAjFfWW3bspY3BGndndQBpqMbc/9H59H/Z/egWN4EewFnml
NYU7K/Yit//P1HdU2tQGwuFHMKqfxq4oUuGIFOdz60Hc3TOZZALzN2Bbnach
alZvEH1M/CfYgITwamFzLlXFwrGLRCxo61wHe0Q0gvXCcexyG46Wut2UDL9U
v8M7QNRJmP9U201D01XZqNLmRN7B0CA7e73AMHy2eWbspVsApo6PHGYK2yYD
3KRMPaEEYWSBw97z8XS0GGUKMgv6I3V5rTkxbCzzQEHuKjBsQaKQ4L4mmztc
HWwmz9ZL9qq1C+F7nkW0qkwa+tV3yVyof1krYr2d5Dr7jpALw7C4GQTd1NOd
xJYaAOG/kQ+Sha6EOu1XQQdZNYrrOfnFvAR+mkBxwES8MR8hBg4kjv6e8/ti
3+FfcgGndIQ+ryCf5H2cP5SWatzNcQ//I9jV0Sl8y3oSA+D6ctE+1xsbz4Q+
yPIaEjwJjPIdx89pPVc6Vmjagt1X/TDtevqBz2xpFGZrTRV9T0wqSfFawzdo
aCxa+cEubFHGQclyaLsIPaG8mmf+40tQXJenJxFnw81unaU1IoRxL9bJEpi6
TQbeNjcclk3J9WjTf4vZYKcasIwofuf1HtyMUZ6MoUtYaR3KOLFXMEhxrnv8
DoH+bOwcBs4UUwoMNO4jqq7z4HmC5hb8tifqoGSOtB5koiGNn5O9pkaIVTQH
qpYVKLjz53hnIa+tSgqjaT2FpCUbzlgR7oG/oSB3dL51AdUXQ8/WXHW6/xdk
/Qb/hJC37Y4RmNGmNnPB+ZpWLXpYQkJ/8pb7sG9/l7lXfJGfnbjFYT9O4bAS
T8uh53Yi/TXwuDwEoRafYsUsQ4+lb2jB5uCYzr6BnK1esKPX8yDQ5xKcST0E
CAyO5iBGvKzyL3qyUVgjidix6uP5kzYwvisJBjQTHZgXxI/AKFjGVRkUn+pA
oIPxIqopCCCpBVfHzfKN6vMEUlVG0DD92H/LQozUZhwHY6P3Q4pdttgr1jq7
+gglaVx6snX6QU116MotWr1juLVV8vEK/GYMjeCvoRRIRgMeCZn8x4iDhaj4
Gf/K9EgCcaMxKaz9Tgwf/SOnQwS5xXs8pK+cUl/DH/G7ObNStb3SwvOtqbd1
Lrqcuh6LGMz6X+1aCqkhZrwLDDvqO9Kjm1YnkSqbWfTa4Yfui4ApSVa5cQ4i
ccjZLoWf5dn4eS2kDoFdyQlsNSJReGlVRno6Yd5BWhbVPeeaXKWoIpjw4iA9
oGDZA2RaugSzASBL6Ga3YOMnjNTzkmd/1OO/9mjLRIHMjvs+TB+H49ak8bA+
M7BD0BdrXKNnoAdkqmWfBCDIy4IFHOrmkKFCXUwsWJ+AwDiX6dxOd/JrWF8m
oQVBkwUMlTr5qICWSZPGasxTDixfRnEGa7vgHtl5oNY33JWRXykuoAPBoXox
Sh0LQaRvKcsElqgrCeLuJRtwU+v28E3mZ8mXnRTfvJyndJ+rY4oZqfAhQJ8q
k62fQjTJcLJ6QVGPicwNI8BGjmh8zody/Riek6EqlZOkHnpOfW6v2CHj7zDc
6HSlrho4BsVCwN90LKicCtKIOKGBCqb093vmADoup/rnAo0itNcFUIpH9vc4
lPEQOJ3u0YUVg5ulBOHZyk3UXgPdhzo/WdjYStcNRU04QATK8P12CC2OB4M1
6kxdj4gbeAv+j0q3tFRG0QGgEHo2osWQ5rccaa/HM3FxlACJOucNW3p4VeFv
MAwOB1wEa+RkzexR5d88XJ3wH6Er0MsLWHByhbME+FMMwhCIm++3yegk5A7h
KTizScAdLrQAOOxbJaO2lHz0P2tRZKx7WUMEN8EOOso+Xo6n7ltPap5OUod5
6+503iPLxuJ3bwhfucdIXDOG2lxUyXg6XZTu0vatf8DdkCeRT4XsmLDCbeCq
t01Ka5oke+gm0dpjnUNdCzt9YLfpAsJIqhxuWrBZqMPR4zw5W4qv/2NgBm3n
PsM1IjWL12UycgV5AAhD2j8V7JXOPWnZM4YxGaB1h5VTFlFhm2mTe7g9PeIJ
GC1QqAcapRCBd7S8Q0opl27dl77XaFhRF4U2r5PJN4I+Z8yx4yP07FoBhfjW
b3ac8eJN6dVD6ucjSFeQcpKQTqz5c/erX/KbPMf2xkC/lpNaztdrIuo+ZoAX
8ba7wfzYY+MtOOw7YIpwDt7sRPpQKnvH4fu99+u7fb5vkWvJo2hbfJy9IKfX
5wML27hQxhe+qEASIxdMSSWYIOiQ20/Z//UhyLg+8d7qUN+Gw8nqBJVktqQ6
fObYjkVHkEZYl0W9ar/+OgQlIYAmB0YLozOhfeCO7FCWV6TuUN1K3Y3W1mx1
7a9pHgCNumDP5cNMUDTEHCNoL4rZyT5ju0RPc/RliU3o+bpegC2E0cRBZWRj
bnG9zMFCYwaGO68uCpvqe6wUFjYQrlOzIQ+fxat7zryTLSwdahiKDFHDxLrr
K+eJ1de7QZWh6zoi9GHKULjWswlzzzTeQbgFNFhffNV6/FRmaw2r0o0v8tFR
lvMBzz92KriPQYeP5B3kr1tAgu9K/MDWt2YJ1qNl8EV1OFA5wmxvmg96fSEP
jhiX5NL52YRGKMQMwFsE4Bj25CNDTqfih9yygttsVpYf7rsFbm5waE5NMx5G
pbPGbCIWtiWbrZeOKAJlVSzt7s5SYBZOu/sodKoVKfXmPlYZ9nwTBNhKW5Bm
r/1h5byfNOccztwm/8lDKxYYd9sLdN8N67MOb8D1RPe1veKLElwl2ClP+ugw
i1AbNodiAsGMIaHEiste3jl4/8iS0HjLJuIZw5BHr3La7jSpfSeIMnKoWSA/
8JO9p82iWJdPfiVxRex0y3V4Q8tCiRu1zmKN+REHOocqT4WNEYF/G3kSD5W8
UOnJNxcslnCb7e/0BQ4XfeEO+5UmHvCYMLk87zJOPJbU889iBqHBF/OFB4Tv
3mY/tOVF0SArO8bga2dzVzhFNhCEno7d8y4o/9bGgRplDKSxOUEAlswFIwXx
QncFEA38DyFZE0bmpUUyL3vHPAR305GXnjt2f9oGSnB6IZZE9Sku6R0TNWIA
w5lokp6zviOObX44coSkf9q8qltx96mZ9UU8+jJO2E/8v6lZ8mcFulPtQAIO
HlDS+tZltsIp2/FIYjWOMwHatgKHPzJzrRVChX0Wloq7y76UBQCdmoxa7Pbb
6jalCChNFWyP3aXqzh7b2uewfM58axTHWm+1M8BhIcsSDoXsO0epruFMpH94
/U3JFI2ztEx7SST8+Bw/CAJrz6rztTrl6/Uc6/3n9UYVKQY+73NnoBo/JqYy
adXq6Hh2Xx7F2MLfsLa7zXmYvbzsVOEGYescap+zdFLozoLEtAC9NYO7XH9x
bpTNnVXwVNMxtQMks2Qx3vCVt1m5fB7igazw1BJNu9+Utc4n5IWo2ZFuUj1o
lhjNbo+g8GkC94gUsHdo0W3fl3gp2WlDh+q6iDAH/fiWVGT+yRPHcbMSsgXM
L0ew8NYGs55KBmyiQCj3IFS7r0wzN2bu0xzuksWEH37HP6a9KlvcVwfBX/pZ
0S9hq1kRci+bacjFJAvvT+Ir24UZPwZVgtih1EQIAaUaYMKAd7amVte2NZfb
zvCMpMAFLB5u2exkESMZKBNGqL4eemWD/t/qq86Z+K/MkZBfPMPM9/4CuTtK
JOm4GtXsHAZuv64yt+9h8qtLVpBwSFTv7h9HN3GzoBT31MDnkxgMhy0kyAur
B8FJVSheraeIWLGXEUrbgMjjXMg52gsL+Oq5YJAPTOyfA+EJYruWGZz5ldA3
vvPeSh12GMKFAYSze09P+VCtVxAiTE432wqF/WoIZkh6UfJ4hjt8o4ivHkT3
W7noGJgJU8qaF5SEacfOQptFrHTTzAvluBlz7mk8H95UUBiebulOe825uXJm
2tSVixZOH7WWtHeToHSBL3LJ8hDzj4iJZ7lW34ds43ztBgnFoXrVpDimuDfx
hP5mTM0BjBQa6oszk+edKkjHulJkppu5ARJg/6JlkAneEwMdDt7Xb166Mgwt
utuuOHbJ0n6L1Cq3DFNseJoPLg7lOgSBR9cbJQZ//z+vfsvIEzHwRfi1XlHU
G/ZIgClPDkFcSAFyiObBAQtAXDpC2k7rs/kqnWC44ga1hvG5d2ibAjXLVkUy
HweERGSriRdiBPKIL6COWrRc+o6IB5ctHlhtOnsqSrxuGRApmzZsjfh/xzar
t30OfBLfHgbatwJiq0YisxKjEJVOp2sFRfQ51AU0caYhOX/qme/+1SU1iku3
L3Sp9zgNp6SBoqXzHeDEi7TB5qysP2//CZ+BFf9JKupmbzq63bkTLAI6LOYT
P5U+FTdLZR/kU6rto5xabwR9eNzCSa26TS6WFEK4LZjx3LOOh/idoXX6JcJU
iPvOXNh11HTwO535lkVNA2R0cGEo8fseP3/Ka5z8RtvgL5zDP4JiSvdnLt9q
Gtxpw65bqePZS6TuJ4qSl0z8atszF66mpVMLm/woaE81H3yqv6siYV8is5Tj
n/OVIeOFL3yTZws3cm0hK8hcm2X7eyps0onBKd+JqUiwrPQrLE5Ny6/Zlv91
Gq0bzd1SiNIAhm7dK0bu7saY4fc1utUXJZLR8VY7FTsqROhcIcIlGAHQv5MH
bjfnfG9EXpn+J0IIUs67CV/KreJ+kmUMnkM+WBgfnUMcbZhwmRNR0EJ08Fqu
lipslBtLj1emwnfaflZRECGpTs+TbXXrqPyISOvzRNmD1YB7VRvqOYwuw+3p
NokyKkS2V1ajQ1Spm740kIJWSynov0HV79sHq2dWbUUO5xrNNeFINnTw5pz2
XiCPCSOE86FCBydVn8v6XCMDgqva2Xl5O40KByGefbjvMK48fHXsel/L043/
IHXoEbq83ze7bliM1aXIeFIFxc4qNGConIy2jJPgOhiYP7HzYrc8ucDfTt/3
SDth0IQ2+GpLEZ6CDpCwIYvws5Mp52jAMv4AEVszUkwiGbYaRd5txRngWJTC
RkyXfxJP9I5RsJMXtJTIHoUy18VHT9vo5DOAk3tDHTs3Ik8cC5v9V33hFmt1
RxGb3w0lChyrrpj/Nh+VQQXaPpp7kTOkmzODJU9SZ1GIXm/AcYID0mJQ9NS2
P1JIKhFQWo3hE6iBVLxNApwx3T7c1lxm5wf63iuPBmwg3ZxmOMhLFYucg9aV
3MurmWmPm8Tsx5U3dxWBmCFNTO5Lss2zsTmw3pdKVBFJz/3bWhMikC9bdA9n
b2WI6ptc8XDOji/Pes8F3aN5jKF0RW9SZCdRUmFa1RMGwpHaZzQbRxdiHZBI
c8u7aaBd7UnHZ6AAWaMb9bUAUma5S2909FxxYccuLUanlKKcrQdJ4wHaqQyE
SE7sGVWrDLr59Op/4AV4eBN/ZsWsWHouC2HuaLeyVoy/8RQ4qGm4FdDZR9h3
dwmgvh/S7SJmJea49oAUFxESwPrZZzUYx23nG9mnxDL5JQKqf6Yf4PfUGSZn
qockDr341ENx7Prnn14XPDRLJGtp+hA8pj7LYGrupF8poTh4RtVXY8ibX4/Z
Au/imixkvvP3CPbpEubYhnrqwoasV+GjCA35dvoUmzGhDp2avidONW+/XszP
hulftA2x4Lfex/4nhz4Vv4YybmFrjujTyeHYqhOGi1sHyMxLl0t9SD9gG/eJ
Bylz3WV7f2Es4nWd20hITu+MvUXkR1ygsMbR+FrOSC7U/OaVdKIjTFClg+vU
5QHVGZgNr2rJUi78mPkqC7fKzclLN2zyo4yYZQ5Qm+1udYFoQBICAlWcJGMi
+dWXHcWhG01O5FekVLAW9ha1CQ65asHYmqIazrlqaxGsh9Zlwgt2zakv4RSf
JGXCGkMhV4D3LZ+0pIYntk7IlUqG3tWXivFANTX7a8NbCTQoshy7RSJAgrIQ
eM9nW0+XgbeGuoWwzZpuH+JpS/zcGkR0Ekj4MyFMlJiv3ZGWG/YPDoG3bxYf
LBjVtPzCXz83Bn9P80p5kJDWECNHNqiJ4ff/utm392nYD+hvMaoimkAw5XAY
DmV+tPnNpY397loAwFZcNXFO2yT2ErtDiB2nDKQSFMvZU9N/k0OA6YcdFXpj
hBmbegpmWQHq+65r/7QVo6EQHZQ/rda3hNiWwK2NBS/o+ZYlSqQwQAPV9ZTT
tzT1q9keWS2efanckscRofCKZaOnH3Lx5qsWW6FLy/RI4X7u3aex2uqYLQxW
MKG2kpln+wtUZKulE3EjZX1Q65FEBNAWYb56NO7A53ef07smJy1LqYU7hM5G
ydz/Iw+fER+XauIWg+KWiq3WBDwDtGOzYraeiRCfj1ClkwzE5aHdrY4fnyPU
tIIuzTyhmy5gauqskEyL7SmaLLRckyEQ0LHW8jqwD4ObFENtqkE23N08v0YS
PxjjZ/PtsmAVf+UdoYbd70TH+XpEvWuZomHc7Kj5YX0zS0bmG40owDDhNRMX
A0tpQG83tKevsgwRrlijAfXIBdcYxdG9+mreuUYjE28gOXKtRc4KRCv5SDdY
fIthXZ+s0KAvkAk9Cwi5D9vQXUxiX1fZtoYxmDfW7FIH9eW97uNIB7jVxURo
b0v40V5Bmsb7Cq4FWFg+6nsar/N3JIpRc5XGn/01dTy3qKc3hc7Syn+4I1ZS
lSFs++oc/m3Y3rHSzIPV56VX+MzNWE2p29gWiDGG+BjXx7huoIYNrZai3Z8q
8/rToOeCDVhg2rrw7TBlgz9MaU8uqH/m8bq8EnhchBSzZd0YRU5uiXVJ3155
WDFi+fnf6nB49ONeEP5+RKBHjDmpJrmEGNHLtZHyDAausNlckZ59kaM63CCF
2O5ug5UEKHaA55ZRByHQA6AhRp0KUNNV/ULmZhwVnlJri80wSfMYmpvTbcTz
Ue7jatlZl2abB2g/u5PYuydxLrB9AOR27mXVRERlbo+g0kTNUGfalW2le0G0
FVC5Kbvw3WZHo8Y54OVu94LLHrDztSqfDODFUZP+QCNSpX+nin1ixtm5H4wk
GlL5MIZcyNPhXA5pmxTEV+/1smSEQaTEoicD5qDyQB/7NsnkOd6GntA26Fg9
TuYPN1avEYyKE1/m57lAdeKzKgAFnym9Eqj5OzEn3foIzBWYvHPtS9fnY4DC
do+dJdaHi+pA8YhjKKZokLo4R9v4Vjp39FqmTqQ/N4SBcyMqJAupKchZ8tju
keWP30CEBWuUU8i0mpL8JCnGEApIDsYlOAi0VHxfVptAIyZejSGSTTEoalBX
DRzJPZ9jSDOSYAQ/nJZjg2KTnhx61r1+twmxWrjozj2GFmoJONdQqbjU7zWQ
8QpGkKRQQ8iD4kkrme5UKSCL3sc719N1kndG4o/1MS2ON5JH2d/TADSFdVYL
Ra45GNUoFK9ukP5xB3sJDs1zO4MoKgPBIElzRT9DJYX/5MMngImSOzo1kfKk
ONjsTbKS0X87F/+qEn2nMQJKI7MYTjhMzUqKeRYBOnbDxz8z2n/XUJmyOdQQ
mLgOx4UDsT1wzw3ZtFtlnKvmv5Rc8WdzWoa+Oxgp4kL2NPPnp4VJJqnYpLL/
/h9xqeO3LFYE1MpuIhCXDV3UzAvM8htq7e+bT6q1Dp4GvoeNU/G9KXTs3f5y
lBgyfmGltQikNloCl70EAJvMVHjHPlFNuxaojq8RSc4rG5gTkv2YdSi7kxjL
6/spU1bQ4MwMXyh89OJldMo8hnPhxjBwG5G+45tIxxImLR8YeiANi0EN3t6e
LdlC1rtbhzm2PvURgBEqcken+OrXf8Ztf/2LfHzMUeMqNPASSePhqupeFkEK
eYRNr6+GMTKxPutq9URM9U9kH96wwMHHQ35hMNSbBIylhEw/przjdgCkJOqd
UM55dQ04/AlSJhkDSPEFLTkKBXYekokSzyEDfqpS1C6OnGEFvDGtqdeh6t5I
u1nlb5pOzgejQXCAOOCoCtwON/fnigqBvho5xXXsqp3Q22+aJpk7UXOeF+g8
gVSPKAV69YicDo9MyYX1at92UIS7otUf9EJittqVnM3gz8FYzcpyv/QpzTjd
12LvcEuNPCoVpuNbsJ14ehimId97MaChLFHM3uTeALK/kpy2YkoVepK8Btvx
2zpS+ZcjLURwcCotfd4Eob9j+a/Ac4DTKQp2LwGCqrEDYQwmeGmoiEPZO6Ki
OF9ohoXRNKwTtXnEu3UHxXp5uB0F6ze4e8RHyZppHvPw22oR4zhyQ88U9tgY
F1PcZYpi0VsRvTd7OajL+P4Rs9VAUDSRjEX4gggFzSQygW46f0uTdIcRTjje
Hj8daqAGtKyyJJy5JTYfv78j6Uxfu0vztYyLDtL1xIaLYP4HYyya4/omLE97
DurCxH/bsrLEfttvfO/D3DOzcvDymY6LjmVcA4hEF7lBEqIgslIy/feEIfu2
3sLsLRQTF0uFeljIma/uZlAmR6YiE3WrGLP5KkHaGJ90UEBKOU3/AXlIZTVx
WUhgayp3+rmQTCSXzhHpGl6IOy3ZtUgiFKR2JB4ZCTKhXohmOlE/YVWgBllB
kgpiEiCJw5uuN4men5/wP9qW8JtkFT0XW3DZsHDEus0P7GJppeug8H/+8vkm
Ka3+knwx0/gc+wAeQBP+hQZtA+AwwJmgg/4eKDHN87Kb61y6EN1KJOyuKFTH
AJDTW2mdKs9n9xtz5F+Iv7jvdI1tCw47V7P3CDmdFolkPFOGMv61j/fH44wA
/Jn41ZXVKxk0yonJ4R4hbBqA/SUSkxuKyN6cv7vnObYNEcyxFRyYJAiF97xJ
eguJsSZiIrj/XSU5EksIi56dsnbd+MfQ3rVFBpctpV2I4+Aero7BtyvNqBFR
xedScgrK2SDoc54ukaBSsSdNT/a/d6DJu6/Bn36yic5LXOatxcSI10c4y/6k
ARTvD1dJvOCVTGLL8GlqSQFxQ8+UCodUhK0HlsHr3gq+8sbHBTmLefcasJOu
ceeOFtBaktaNVoKLK+2e//fhhhOke0SbR7I2J0GHd48DDAMb0Vw2YPK+SvrT
azabga8H3rFLAz5bpvpZ/FD+sCa8f+JhEdzpovLhwc9ckX80yf1OAxM3ydM3
Nr4qJzf74abEw/n0Z5sUB/+IdyhfDp2m990d2ckAW2r68JJDvWI6ALgjAllO
PNm8ZBDhbC4lWuj/BJ1+AouW195DcN5CcUwfWyJN0l6hxztg/4i4OVPZs/Ln
hDvq8/jcFT8+sRZEiZoPAAiFwen/BU1XMMcJjTMWmrq79DpZ7BX3Hh5jVcor
PRIBaBBECw+33hKgUSRpS42jdmVEq7oKA9W8PqpYGK3MIr+AyG03EYZ5EVyZ
O910iN6RNEpnxSkMv5MjGOLQj7Gn9fWOvHZAl955EZkxQvTUETJkBuSNREOp
swkyBuQqOoO2TRWik9YPS4M3x/1mv+e4NhT7XuGHNVIEE3+XXuT5hvmMViUf
J0wStW2Ts5sGUQmvIsanCoPdqlPSBZj7wenhlpO6Sz49iyedM55rTDzo5dkR
2fYfKx/7PwtOFw90rAfCz+G2BdMG1DhTMvzNScFSX3/lj0y5ff2148Dtst87
bIkJ5+5G4j+v4FrrtkrdZb7dtG42HK740KdVdssSirpt9Jt6/sWuCWwYj/iy
M4ZSmoKtOpz0KIgyV25mpauc/kzN20HxpTZL35I6NyT9VpUHqLJyDe57GPPG
JYiDxW/BTawmpiIp6KSFe9306puS+e28ISR/+ep914mLPykiRP4/FsAJUwye
akqO8iVHlUxc1yy0JWPnmy3ptiH36CKhoKBiJ5HHdboJTZPoNwBRZNpLHo9H
y+KqHvzNW0DgimRu91JO72EZPFZu7rBXbn7aq6I39FBNJsM3UZHe7hVBPf//
7EmUXfl0YUtdNOGIlXWkIEuYbnwQkSEMfXFzSQDX25pMJQ4dc4dBfVbmEj1+
RZ9h4yxNWcr4+nIssv4BWfESlk4Mw7byCoaqZDDqrjIddE2vNEOyxM8q/JHw
VtX8AEkge60Lo5KpH/hPc0wrec7IUhLBFpX4WPVLNSGlGfjwVt+TG+GQJW7t
b4SUZBFfw3iV3mKr7+YYfXEY2sD38Wx1Nhux/jZxTaUiV7WW/Rk5lkTRRvLm
dtxOiw8hWnFO7zz5x3yKpUX6l3xx8lMT1H/HNlzbjwUfQVUhBWZv636WwdY2
b7TcI5wWGyVip2k7nWRhV+9p2ghkI04U8EDCGLLPthuT5Eko54mYTBwGyKV5
bvCpsbH8gYDM+NrfV1etvN06o+cORJDTJNkfYeBa/CVtT8v8IjkOte/wHY05
9uenDoJeKRHBiuyxPGXv2pQvxqXM96TXfFpmoJ5ALof1cNKwUyJb1SycWX8J
O2I7lC/P7PNFoPmZYOYeajIQoUH9R9YaURYFNSWNUS2WTs/OKzeu+pE06rdX
t96IbZx98X/gdrouzdsVimDYzzKQjbfoZqOhJdTLwPjHA44Ywnmt+puUaPic
VR2LLck+G/NshdyBJeF5fZ5/l7qsc6vo8fx5QnnHKKAbtfGxe8MEQgH9D6YF
LqVb4kQrn/JzBx1/hGypOcdOvQKm4JfvVkH1dNvZH5D1fvENo4jxsWG21ea4
Y7D9beikTQ5VUCHdjHcQGY4NlIq2OK0ziwnY83JGSemXOL7V+R4Zxvvx95NI
kJSHYsHweWVrIEYtk5zsep9bhBKtt5bNBeZHJsEi5m4jPXH+QPDOK5pgNrm3
k3nMiD1kPIHe3bi1uEog/T9mevEe2YNF34WrCwMYvoQpbtN+hV7f5T280bGz
mnZ9HLieqy8jVX1tdSBsBU9n52fCrTHD/FKpyOEg9aIxSuFIOtP/JlDGI4N2
Y5NebLbcWoY8UiXbiWtQ+pKPHe0VwryzxDHkjMrXSdQyOlmfeNOHmu4TFf0b
rvc8d0ofyKcBeqIt7vAT0T4dLHRgFc+1HSwjeIuZhmPCaNmZM3i5/X1NVt/Z
YdidhOUyR3KVecTkJjZ9ARelAx43CjYGV5D/G8DDwMCN8MoZuUGveysIhTaJ
Y+4ZbDbABAv8gVUtDkuLGN5uiTPP2MEKa5kYg3Z8o56cUP+cnUDvHOeWwXad
OeZ867BsSmzRpT8RcfeIceDxv4onuuNIhE+J+wFyPgseFC+iHiAkI3ZSpfRu
lHXyGDtWezZtCuusmiP0Tldyecoehv43uHkOOf1QVPTA5iufA95bQ4tfwDl5
5Qk8LKE6ofu0qRknxC85YIAr5OGiNw3qFYxJSpdtgJnnWP/xVVKlrglcrR7b
R6mP39K7Qg1CMaVksImThV0W3xk2X7vK4PXoZxxFDPYHYG8+8/luJ6BPK73A
1sIJ8eC1IMpM/OZWoCDacyPH/YCdavhcwlHmEuh6MjnR6QAbchq7LHbOC57l
6yRX5M6ZK1S/gZBqDn+MYJSGTWvNQV3iouME8SHzcG+qav1ZB7cg9PFdxQJn
rW7f1HaD6t81dpx9emZZhm5HNMDi3J55K0LQbaNOivrYvgIeZsqAzDi7PU31
47QSylVfI2N3hneiuKYs336jbLvIFDmz7bUERGxAcxSM3KHxeL5Xr7jz2y/N
s51kiE3NH1x6aEjjrdaUfY7mdyO3FIVS42U4dhn/7985rSvGTkX3iXgZoDu3
R4o+9/R3InUyvwsoWgFtFApzh/w1dOl+IMVMbLteIptPiFtelGs1JpxKCgl9
JM/uP3pMLpjhLk57LC9ixzjGZirMh4EGR1JTetdi0SlzkHdII04P8NQBHPG7
iJVABMUwVp/8BqU3EYnubUYmGV2B5vfefZfL9wvPLJx/GYzXf+XbPtIJblEj
cHPamBXTbDdxk/AXQdPGkmWEqC0HUCHFKtjb0QfzjHSDhJVpMFYOeltUal7D
YP10REkVRVr1bFLWky+Y8bDA3cGAVd9yaFhf9mazBBHwN8J4pRzIFAE1leXC
ybb1g9Wz+5n8fyQPhoqeQBhvGZoc/HMb1KH7gyOao8ZjZZM6CTniypvU8fRz
Yyx3q8EbMq7gfP2Da89SBas/8zNwVbtSRqoDRc+O7fP5UQvlbZj8UKnWcCL2
GhRpFJjX6Gtt57R6sKzjbFToiq0n5OP1uKdO7NwRTKUMIT7a0t7+eS/jSrP5
ragtcRtJ83RJA8iBGHBT06BybZnvaF43XE834HbIYzETUzsGlEji2U2tfGAr
vrbtevEiZs+p+18a3LSKKkmIHRDMeqS4qtyUrkin/lsEj5dh5dphEDUJaU2G
phjmMss6y3Q/1wQa0b+/AtBEIL0TP8bhPWiYcwZpBuRThfwE8djpgpctSzEq
X22GKvTLh56ujoXOvsKPLJHhkPCk2yRLrEtQ1AJD+H3yqmx9S8gXcuSZtQUQ
xAMBAdskPdsqBo5bOhKA5b7ss83cnje3Ef5gGZymnfmpJwHscpXbP0AYVrug
rp/4n5qik+kH5T0vwtkYTlXUoCaZkp1/gPxTg/1uLWcbeMuEv9RvtNk4OXpU
X3hzGWpPYfXoS+EyWRFXJYUALjhQnsT181pMI6kfrhoXBCIS5XqQ3EHUtuQO
3KCPjC5D3RhSdQcxSlWMfucmUpaaxKa4ubxEAN5nIVllQjRKGZ5TekshMemt
e58OUrmjDOrzfMqu2DPwuj0bNeDiXwbebIwemj/50XQvwKtcuTYeTv2e0GJA
gxRtBz+0/gYhVdDuHrYES+z0JZHWULFCYDSOZNu84wHR3F6eKbiEERdwpZ3u
Hm2zsxTuJPS+s5Jn3MgbTDakY6WEyXC/raZY8SpyQe+aSqdX7PknhFhryRun
wJZLM4KTaZlJQl/GsotfH2JhlxsSiU3wkK/AfRJCCr+y6rDyqHiNIbNtdKBn
4UFplDg8r8KasGgvcy9os0loKxpub+avFrgie6AapSERRwy9vjspHzLDLknL
Y4jYharOuytsYuRcJnCpUP+tGiT8B8oMGqx1jyWIIoy0YvON1rhj1rYCAyKW
X17N0AvaI46DL5V3n7tOn8zxyjRyEXRC1PdzxjXmoGiHfrqA+rE+kbefikEL
+vVQu5+uq9IPqQiwp9E5pS8q+y/r0XCWlmt5t5F3ujwhGJnkMmaJQ7u9i6HI
sXsMp6aqdWZlZfLK1//Qh//MQ4+UFCorE/bo5uj+OhNkdpIKeYlBpehgF6Ny
kVhwHBIrAURG4nUD7q0qxmsq49yuzkfGJNN1K94TgVpBFb1uRMET7uNirBb9
/mS3B36bvxTRzXR4oxFzVBfcqTPqe1r9fPcE2VsC5WJv8i3+4hb1QN2cBus8
U1CZ8hv33/AShUT1mmnPqjCh80OHDPB+ofvrJrN8BGbWer4WsmrTV4E4HazI
V3XkUuD+wXwpZcfTq8FG/jLz2H7TtjamSzoIzXkFPp6b4YHx31stGcUER0Hc
3ROSMZxtDOH9iJkNTs7hibUoa8jPd+a+NWIfxEpOUBdnVcPMgkhoPuZcc8At
W54uoh9FKIuYvRFacUpamGHbvQIXsn8952iiQgzlx6QkwVsXo33QHAjrzVjW
O0FOs/SX+AhYvwujKkhSBW92jBkD0+yIP9WPgVnOVacVpsGa2Jf4UVVUcBlH
d1kXRe2WEomsVK26ETEqW/MqH6EnJI+BRVIn6R03EfjcTii0YC3QoSTS2UMK
a/9vjIeH/OLRobieHkhhJkgzZ9XVeUzVwzIBCCfpOZ36tt6xaS+997GaNsda
nGZ6RiJg384hUQXsVaWH0lYn8kLLCaHeGz9t5motqDiE80Jc6oe3bye/OyjU
xAhy6pIB47iSnRwblh/c6S0XDR7Lqh0Vl0Wv8QIiVJk29v57a3kjRSqpm93F
7lK8j7Qisp1MdpdZu9OhXsxb8eQhrQhKuS6f8q5yknh2OzWdP+wW6ilbZ0E4
MKpJPoIhsIUpADsTketDlwT+HfEa3lC61XVnc8zstE+eK8zXCjXJeZVRIvaB
TNnKusxG6Iiodfr5kg5lhJjnuNyqyeHVDjyVSYQSybjrG105JMKoJczMR1hy
EnbJ1N8pkbVdwxliy0H78ayVKEThwUsw0VsLmbvwNbGFnTLE8ewWKN4ssfwa
HkXTpUeWx5Rp16jI0ivhBzX9B/Wf+MImbhy+SnKKD9Wz03rpFdaph9mcbrR0
ocJzvsHo313uCKyQVzenzXBaeaDXICVgiabIW70EM5AANiHnUdvCrq79v7C0
cg8DalcmJTOBeftjK+JsbzbgIcVRDQs9hwSz8Y38mgcTFMQImlZwoyCyI1hD
BS7DxV5NhaGZChsO8+WYMFZ8ERkzGRYZ68UDVBlTH+rsOUDl4ghbuF/bSXBK
/KtkKeGIVsAqJsdehUm0uB/KXkvsRSGPzipUrsAj5WeyBIYb1nsgAJLmTHnz
/DHwL67AD1x6B+Lg6M7/ySZ6yYrLLCXQX/fYp1e4YdUxijDzDyMgmP6TlwL8
/5HXus7MZZPScxX13KKuwVQyTOwSxKD215HrzOONRy898iJMvihCPEN7/9b5
1FCldOQGAigGkfenVykIXlhp9TavspwNLV4grVmfunIDFdrCuQWEQRm6m/Wl
tZ7MML6yzxFpf2bBobb9zpIdnQtEZuYpO8WyVUFIniMdWuV0B3vayI12dt9n
o+4PVHGd+OVz1bJjhFKswvfpZrzaL92kwbbkekGM+wR7Qv4S3RRdKRh53TrT
KpYra/m7/Y2R66+n5+ms7ENQ+N64Q59nNdbuNpL2goZMwgT4mlncQU8tOOp2
VxbvC63jFanGf3ddSxuxXQBNW7f9TGK/ev0Pk4S4UCCeXP/sd8m02g7JCktL
mvk0dez+dgLLkmMmaiuqHIvwt5A2jy2r85ZVGaVwE7x8wKa+PQ5YiMqcldo/
7VLMWk3KYSmabC5D/it8b5+8UgGsNJnNcKva9yp49Z+UlQ+W0IUFzo1nGz9L
PYN47ASTrW72Dp84QATAPoEbhaHJAek3s3+HtcuRhTYdfNhUFhCT+G4VRuLB
Cq7aalEvTcYW2cCOPTIQ9ogH/qzxgOM+sC4I9yYdWBDdktVzXtu2D8kV86d6
07vbDrbkVuZERL8HCUEzSmGjGKTo48g8OkMYC34XthyWz/isJF4UL9EVJyyV
VahuOT1vYw2tfmBOSnplN26aVFM/fKSR/QNN4e3J7QC5ZTz/zVO5gXhYuXmx
ounjrWN9whUNhO88oIb9yjL6M2lUMN0qybKmM+X5CZ/xEjvIKeDxODXTdSP5
SnuBN8NTedSQlCioqtyNtrN/cbV4rRojLgxheVP0r4BE73ABhMN+M+YbWr4t
m/3GrUu7H/4JHpVv/IJ4MLAGRjVr1D7KRFSwprpUJaqkWh4KR4Ui1ra7v4Mk
vRirspvoWqCE3NZYG2IG+ydEZ60/LrCRGLqFV0vKrHvsz/2iYhdhv9UWkTgw
5EC1ZYGt2FIMwu1ClfgoukYUpjrLIUhXGlqkL0rurmL3RhGqP+hpj+sve6nQ
+aChCedoL10LNiWskMrHX1V7AbHt+EUIl69FODo9GgIWXKPo1u0ecTjHyQrb
x1QEfN7y2xfVX670HKOEZa8ft2cjy16PTBZi1/Rwc/mwqi7UFZhfM6NCsTIO
3mQVrsn+lVfZBAn5mAtjPQ4OKYM3Zwj9LKQ9beSKYE8bN/VKWLksJKOhWxOR
9k9wn0piowi6dFGVYl1etL+h1WEs7h0d+6TnL+u/miP2uLlcm7ythASXWwYH
lM1Dm1hckGBOz6ea8DCZt+WdlI1nN/9525JLPCvWosumf/YBJESE20baJy/6
/hg0rTcDiKgyfsZIXNRI97BafkBDZLpV7eD68vd48ca9V6gjCS54i1IvpvjZ
dGLaoGnu3Oz39Xo7t7dxo35/P9oiEq3S18cS6BzEV+GofmhJeXildZF48oaA
Kl6GYF1bnIL4LtOgtZLkcgVO4jMzuIpihVzJqehC12QrOlHL+jPPXX60b7vp
7E1AS5bAB/vCV4g/Bq1HAsl5ZXfYIk3882TCsLN7S8JL/v1oPZXa8qOyDgPD
Vmm7ovkPSsUpoAFr30vpcjx5dXd8JCOsuc8LmeYf8dLNJmyTPnBiT9XLBcV6
TCnRz72na+/5bBeABVF10wUmqWlPM0Gt9Eg3lwp1ERl6h8pCyPotUfoUfInj
4xe2UpoRk+PlNBYtNsIxO15Msw3tdce3ionkDNlfy9TWLnsxXRwsqc6u0uL9
rxq1Hc7reGSObutalrpZgymYFyKJC5I5c2D7fwqPOJ6GI4QH6DJtQGucYXp7
wJUhtb3GM+3Cz+B4pfbH70DaTVbxe1Ni+xzdNR9+86uvWqs99+gQz5QF7Vhe
s15T6Ql20meC5CssCO51pXOVVvETNiIMAUSO4w5uvgj6D/YmKe92JmbWFvRV
Xy9Ppz8RPLMyQuILAM9wwFXbCv7wKP/HbZapXbiSBkU4Eztahm4x63lqtBkt
xEjWkHA8oeypZpli97spDTfpyV6YW3/P6Da5zGEswqJL+MYNfLm4ekL1gkXy
xGA4nLzimQHLu//OKla9f+GYh0Qm60o4K1siADqKfJLP+l90kF4wokjSqQq8
DtnLHqtaz+m51lBRJ7O7X0VjW46/p2waEEv+QAjWMJxpMLBDQUDrvJrE7Ua1
bwwmGunS+cCAVqnkc7BHudY5eN6fAlY/yVZxtlv06bL9QFv4ERCMH18oom+o
1V3Euh4J7fAeoiYPTQD5KTvPaTIJopieyl6fr6q8aR1JVk4jz/JbMNwdE+kB
rpS+ApgRcjIvr8jNPlKonpeZURhn1v6Aj+4lUDpzD316f6ctpkHm2hEX2rW8
O/mMloVNaep97sBuhlERTk7kYC7lbsfNCIAI1s2p1zQrqn4XxcqXfpCtqcet
JER7A2AgI75+mmpjT4Vm3vIJ7SdzJ+f1tkhTQtgGvcbPRT+tU7V7YImADEMc
szVLGwmQbEK8MweaVl2v8QlO8CZVi0KbCDT7KACeLmPb6bmNgCAhLUi/dFON
6fNHDSMuF65mEugsteTy9Ke6QFtjAoD4AYjxtj5CSPVFnv121lHja8Ti5pLt
k8n4Sz3Q24JVL4twqI4A/9V2JyC8N38Suhr2UUWQ25r+ytDLZTpGqBbOu4QJ
vl1BJnfxPkoMBdV2cugoOj+UK47m5Poae6bNn2Z3tfbtvRFUyNEwjwQust0W
sqGLRXr10gKQUDyo8uiv+il9+2DT5qJ5nqJGHq0qweOsHY9i4xwNxfsVtYEO
znebisjj9pJfMF0Qz8pthf8LHG5pg5dK3k9PC6nsi0dLIGbx4nsctJFF/I+b
WaTN8+50pUNUT3Pe8fq63BkScX71sN+MvsdeHknpsqKA75y7TlzU7fseE3NJ
iNvp2wChg01LMycim6uoRb4b6TI3YBpvSxjP04h5hKCyuxT8q3K92NIgYgkb
hqdfMQIlE7jInwto4MrqbN5u20EpotdUBOAxEkvCkovvZThnSdwo1mABCg4Z
1/dKq+ZfqGt2pq/qPSnzmiEj9wVFLcu8OlFISOCIqxf61g8ELM5KHFwSIWf8
y8XOmXJjLBjI+RTuuPeAmp2xt/3jS7rHfkyeHXHyaBekm3ta+mMjM6qrhhIf
EhRulU1Kjv6ZECA4ZIdQt2xdMKmEcr2PzjV7+I5INsN6LItmNvHUA5p7PvUY
1OERIXBPD3HjcLlpX6sUPte7ThszOqiWizsZvciQwFL5EHAj3WKLTfeP5DNj
nQn4VTmMC1wm9UdZiYUeml7+YZ2LXOuX//4i3T0G7XJ7VjRwI8CzSTh6j176
2SuLd7IFZRUaBGG25wWOM+yAt3R46XZscKSjudhO+kgWZFzTRtgHa9Yvvt0T
3nsmLV7qFhvMa3ywJpKKz2yXO9fYASlZme0Yu6vGAkP0W2jzpyUSD3YVcc5G
aNHLqBBFLaLW0E68R1OjLWH47GWB/zhJ3DxcYR8wArwVWGDwROMPdbyNya9N
64/TP1ApbDTUjYQ08VHbpIPfJp1bszWTagejyXf3bNW+fAYd46D5sIw4b9hT
UdD8PiEUZB+4a3BNwPI54KviW9KY7PYMrHMgSRL5uIozlvqT4/I69CkWTjgJ
7mnrSnubXTSzB1ih0zQPO33BBHnhZnpuhsoz1rANhtNbFX3LEN1vRb52z8Cs
BJFiBwMront38jH2w8kz0aX8Pa67+uIqZNfPnrT3rDXErS/PcqndPiklH2cv
w+F9e1N22XOgZcZZw3FlYUIf7mmAdnj+taHjdtfcT3hhcVejz29PN1/bxzH0
kjtDeGy968JJ5FcC4g14f5mPzQj0nea7WHUdLQgwNtUqY4tys2FMLMVQz0wk
q6sgTeOU3PkfvaIPT5SgvukfCABlte9JbwV0kAY2s4p6F2mYy/Uw5AEcgeZC
A6TL57gD32HSwp9LCFRUkTjACRJKCbVP748yBghwmYD8WvLn62nRjbQRqh+d
AAHTzJUtSdmxHIWB74CjsJ1EAnSzzB3qU5nfnv10A5EsViPpXEJyanQBD4Cj
Y5/32Zn4wIo1fbnNjAxEkiksWluxQMZ7WGicxEOE7LygLTvY+NM5FFYxHBQr
RmK6ZCszJnFBJyMjL3rGT8qTFfJCzlOmBixqRFIkCfO//KLLKF4qeSpTvepH
uVriRCtNGFpN2REyQ2pl+BSTGLOBnb0YmVS6omFsfQYXDAIvd2a7Q+pPlGSh
V5Jv7QEavy1OxvFbPOTPyRhDqLx2Hz/GrrCiGubBXInINB/v3a9Ccz95KFcF
AmrICI7Z+EosqnLfRqQ3XP3YmLglrtKDu/F6R8PmxVQBFYwlXoOq6MCSkva8
E9pq/wlB8VbQ6VS5AUzY8RJZcoZQypOpRl1R4ovf+Ozva8jxCFND+DIEN2be
TKhaVDa1RRhDIi8W+AF+LBKzl4kRCbSz/95Frbb+iktGuEWcq8caLYCO+kY6
qLHHPEyYQqhdl3F3My3iPdzxI/hvi58yf0L73ReFQ1S9ih/L3xBdtyM2MJoY
aCQYfgF4mNVvvUhB6wPm9D4IZJ19h+JZJ8xlVDM/HNQvIEmR7I1/E7oGhasa
j3Qf7Apg5LXvVqKDoP2eBgTIG+WB0RNwzIIvl3Yehc4NDSQKRa5YAuN+/hB+
6aA8Kt5YjeMuBUAPmVPIAyU6CvZ9WLzp9FYwwzu/mbWKLDJOkoWuAmssCiQq
7uIqYjdTwKOgvWRQ/guz8Bx4SM/Jl7lSBnYOeUgGhfaF3zpZGzNO9makLX/V
jYWzz8zb/1HsGqpm5fE/gfhI421UbdDbOSH+X89CVdzo82zjjYLqNHLkR15R
0Rapr0bGrNfZxnlpiOEMwq5ORP5GGCgFeQ8XhNczPDmrk/PLZ6C+FfYzKLVE
uzRKskwG0XZsg9XXsrxH31EIvdY22rSHPFmIWdPykGO+7K+3NW+t4jL3mvG5
xSAKv9SgW3RR5BwmkqkeTlJ2tFhZPiaPDel9vi01Vs21Gml3l9LAD2qN2xPA
P4p5h0lqYRT1MBtFf38scZkpwCYqwSfbzhYbxYF/1vkTOUmTagOvjcSAJ2RJ
3pbUTqnRZ23rBXdub5D4f1+44zcToznwAFZGDpx9YCB09244io3oqz2qXXa0
tWZhgBi9rh+tiAoyDWT5DLvvMadxmAXGclI1ypVo/Dk2R6QPudG7A94IBACO
gdytrEnQPehPeUz84pWS8X8Fg+P95n5c70lskRWfFePq7cLGn/3FB9CM0TIZ
MYyJsCaM+v5Y493JSm3nqHr168Avw4vJLtmTmJHCwwota23rDZPaYxAj/BYW
7kMXeTV0AVdEq1sYG/CcKpCr1vcKe2SU3Gm4sk3Rn/0LxbdS0ues2j3IOQWt
aY6YQVa1hcrbRhk7xP4ohNKiAU0hE0CTcpuzi+Jgno8XHyM/gwPKy5e1YZyD
u7tItEbEA7RA3AwogYQEpvJeWiNwfnEXy88GeMa4hGMklrlmxlME0ss6ZwSP
IzziSgBiaA/5dNVkB093KDg/BtonoArzGyqGdkVE0Lxq5qlr5pYH/YRSJ0Zq
xIS0NZp0S436kNtdU1PdNrm5NHTarwcKT0zZDqx7eTX5KgLpDSIBAixKboqK
KN4Se5yI7QrXHbFKuelwtkar+oLBvbfIZUki3zUxoidS/rZwGH9tEB/9PMDd
HdAPODZqRciPOAopHXkgJtcMZizWsemOiUa+WntaYbqULWVqz0scsNrVJk2q
Um6DJ8qzekIVdHvaAwns7dUkAC8j8orTCVsQrEqIMIS1bEiz4qkLwcS+sOGj
4ZTCwMIEcHliKs/gXe8aRQS7yhtCHvQmDSZykh0wrOH62HWpBjjqSPbi33wt
qeb/2X5GGE7NVQTege9ucNNAeBaYtS0KBXxi5O0qRqZ2UNw64nWw7oSIhr0l
dLkV8WpSAe6jqk3cPKYKbNbWFadfVR6XS7DYNjpUhHN1K35KtMOWLGEQ3Lwk
pJpxYFO/MJJ0Go9oarLDVG9/h1ufGcx98Q2irW5Dqh/CBZPxP1s5/pHComrq
Q/vVG0CynQF/qBNeEFghq6w6H4GDCfCE/jF4s578bnKEby0K3TCfsp2rxmaX
d8WDySBuCZfQLwOyRSE9FlWf2+G9DjVkRj0orMp9zK9BFEsVMnXJ3+LAhW3k
bAPC1Ratuf3rK0EEibZPtpWaYVyZ3bG2YklDA8WFr4sAWSEYeuBJ9mzK+JJk
2HToGRZuQOGCb8N2toUjaSXhUEBb7RwiYLnRpofsdDemnmsFpz2GpoNNZZtZ
WPGhRuGLA+0oVWnD4o7v/0GSrfX8lNW66XOBjOUYT+3GDkTx77vzaCvA0D+E
Ykx+etYjFWS3MsPD6E6DRBS4sC5iqRGIhxLvUkK6/IQES+iKUoc/fwSAVUJb
5mK2w72p10YHlVRQUgS9QbtsfLjM56linMvQZ8cyVOpU0m69nMrMWx8ue89i
cM2kjZDQXMHTlpMFPe6AxpmBVGwFFd+l3Jc9AUbuig/DazbR/OnFOqv+nxo8
SiJlKwDN4Z+12HI8IB4MnivJ+D8m5bl1TIjkosD4+acuDeq+niRj41rze1L8
WtCtRlGOhhWGESQtvTOfCT9Y1nJWnPwD6IJQQaKI1lFy8lIDaBSdjBr7Q0Je
fbXKDjDdoARRi4Zs9sJdkyS7xQW7QqCA3k+o5imKwDGMYpxXqesR/Feo0MHO
PkYLQLbu+LcSoE72iiZmyszh5HC5/OjuouI9y4xzQBdkifuda+zCNPN5mXzx
JK/wYOnvioXS4kKiMzHWDZSG4mZzNXYS0An977DkskslwDowaQO+kqgfs0QP
UzAvHf5DfQ8C0lyQ+w2LuiMSMJxiyH6xv1lHylHsMyDT+4DutX6KjQUaugw5
YBxnzbVJaso2xSkGMarpuagbX8FBc5DX+70yp4kjfZhHIPg4W64xLPzp1drv
BkanCHNzNrcy9dJLp8Ayw3EBkSFdQggHhM0iE5Fx1Yr5Tk0h4bLIcsYwuj2j
2sbFheD/Fab/wVMT0Qwa+zJahz3QIn9+LIZOf/tHohnlB4bbSLwGlyUcN4hc
097TEPtYuOOKrZyKeSySROAJFMig0lCOLXCFJvCYFPwU6XTKchaBiENUAUoG
rJZiArJ0mATYOFzP5DhMzfd8ZKdqpA4lMcxyXA63wZuI+Pak3EFwPuU+wnkL
sUCrkbQaqlE3W7qwlXEnYur7+FzXnlkcTB9WVRxuEcMClQWfBLSAkJ3QQOYQ
gBhYJtM7pKthUB4HmEfh1OLbyp+pmXEt0CyLEaiIykFH+4/VjSaKW8jJ7Jz+
B+zm2Eg2vIEBEihSSfSuOyN3pLBxJeQaXSra5uYVHOjB6sxRMTmaxRxcCFn5
ADdkcQNcXyyU+172LJgDPZZSN+cnxw6UwlOs4WtkwTwKnQCSgsh9VpL9syFQ
FNhAeJMbku3XxKkmidbv7jF/gFPHLDoPwOqZUNb6f2etdeK8JtzERaQHeKoe
LzQODY0+kIjsEkPozU3p24r2D9db/YXq3ENJOJ+3Hlty0KHbksU+nOek1DO6
0esqVrv7pU/Y+sNO5LuPOf85djh185j+i8uuYYVn9EhN2H+Pr3cMPYZCF5X1
G7+iidr1I6vsbuV6bX0iAokzOYSFDUEO7QonpmqDMXC6Vd8dGxsxnqqXjpLb
l3nBAxqNMRfE2JMVA5XjyOwL9wKGWlIy+c5K41hBnTuSo3BU92lK1LZsd3Fg
GwvUYxJw76KW0j2RJr9WG7EByHtqqNXqlkkbOyoNnaB2Mnp5zIWYQWrI86uo
kiiXvx2vkXsuTzI0BYlrEkbX5HkyzMUwJetwWbp0NfrCnSPQ2YllP3ghJRwV
kHA6rrnrw+JUXzntd8http1JFigpElA1v3Y9PUgCR5J/ycYf6QJIB5bM9uVR
zpA7gtLrS1VpyA/aNTpOlbIng9GSokE25N7i7zo2CuC/ki5oA33I7gzX+hdg
apKaRBMF8mX6vu+/mh30oBDZad0PXEz3ZAfQivnL4LSZcDEpOAoFEYZ0QjAj
CgUWM6vQlfETp3RPxfXC5lpa1TuxDFnUbHT/huf4U8SC9xklkOQah+O3lCGe
DSTyF37sPoFE5HoJCsFOZBS3Rz3NThoKgDgH2PJ0026Ugnlr7Byje4vD6ZYM
unZbpiNCPrxiC8u0B7t/xSdBTKcPLuwg2TC5V3sWFRmHnoDGI2DgMOdalMAQ
SHcAYgbS8L2MmICarH5NXfOXyiFM+rK1uXbpbn9GrqyAaQHq/Fd549QipyOj
IwkSPgQMrUdJ1Lv61arAnXh3TVVf2dhmOUhR5MK/JVm95OP8biI2C8s6SV6t
azx/SKe7plLaQPxxUQVqkkuOWeruNxKQnyYaADVg7j654siZlOgUcGNKNuy3
GvUwzSsEEl9q0ljRxhHJ1YUCGmoLgHl+llBikI4fE/m4RW5M7gJE6IpZTN8H
x6YcMggfHaEIrn9J8BnC5Wbx0LyQBtainRPMBmelczZx1uDADdAuhpCA2dAH
D8xu2eVEOBAprVeWmbwH85rF9GszmEv0s2DB7N5NOeGShmYFJjbOE/muzoRF
9K0DoPrMdk5DeEriHFDtjt6Sr4ga0FREx+dQ9Nuyllftshg0Jtgy9UDksMoZ
vs/oOvD2CADAiOZlaah/GrqqeFMefc+9xcj3FQrbWbe5+G1yPXfAclF7MV/2
u8k90Yfd5KZ3rL6rnIodqwG8wK3/h+62wXevVVgAdLwkddDGP0ECYRirbcB1
x02TkkdtRB5BJPgfgD95bm2e7xfAGjZdE/5HP7klXQudC6W9mPaexpsa0Oua
mW+NexYuBhFF6dosRBgVWiF/7qbOkovtpg0GwhBIn5BlqVuBORzCrRTTwaXU
L4CFQOC7We184uFHFhZQKatNsT7dQan5LhWjI198JpwQTgAPsH2UdZ+nJYs/
7UwCazCHixpR6ZfUghDFr8O/pkKVyor2MMgv2iRAAAACWNwl6xwAalbnGWgt
sk6IIMNStSn5k0Wgz8npRjs8vCxoKNA9kGtgcVCiAQ22lvGphmi5QCFSHHTf
Jlyfd5+BJndORu+hd5JYO+c7zhBUnjNl3V9bVdhKaw3aLSFAeLkxxZtDqpor
xLnRgGU72hKzMRjTkgOQ9e01ql/y6/7bZZgoKiH4Tw8omXv4WmgV8dF1rSYv
NsDhb883I65duLIZvraWSzbkhvpzAFO9tN/HXguvqKgziKviTp8bjUZ7QvLC
xvZrMIpNUGbPqMEm26ab1XQnr8PnBkSiLoMUeP+9ztlERlmoJnODJH7VmwP1
mchNkNnZISHNphzCotkE9nqJHy60g1MrSZG1BgqjUiShVrragBnwrtl9btN4
Ayam2oyUos3HncHg+kDn2xyeAamyqcZEb+5a5cL3lEMj2JbpQJftRvDSEBdo
YfNdoD826x03022eBaKX6OzXO1TEUmTQkEDixdlWzW3Htpbpkkrh/fkv5+Pb
wHfKvWiZiLi+XQ/e+nMXP7FkAazibtaturfy8mvcHpbGEY3qdBrvTXt8ejvv
kV3dT9qaSnNYLliQ/E+yt0v3maYqjaQ7y1SizbcgzldKsIs0V1V2UMctgfOr
VnTVVJfmauQyAcv8EnhWH+UjPHh6IJYh+/0ZJyfPxoFa7rUIesp+gpDVo3Fy
B4hP3CHv7gydAKAfTZnewXtvLgKKAb9XEYkva6uHo4ApqJ1/HbaY2UkLz0uH
eHKz6OQxEYM71/H1VdTLNs4+bNBKjzmqx/BasXymw0J9/Qg8368ywXSGzaIu
V/HFky+pkd62j+bM6rq3uoe7s3eaAaCejxVL6x7cj+VDgjaSW34x9NWaKrBz
BKUdrioWlGYelcUNdnJp682vaTXiEgxEmas7YwCz8rA45eP9FMI+qDgmDrwp
/AMbtWXPoxBzqH7F2ykkmM/ruqRNq+hBRNAtC0fT28BRt3O2se1KuXGwXqE9
qj3rsOEgvKgpWQTJ5DVFcZpckRlz+OftSmfwRr2JJIdQ7n5uhdMtVrgQq1q9
yR3xENXiIKwg5TZCJiCT0j57aNyOkIbDBGyGqJf0Ipuxw0J7WbQIF3spq5OB
Y0Tm3LsUZLJ1DvhAaX6t8SJgnWyMHboHQBsZ48raXRMbXSYlETiNG94Q8zhe
7mHgTxlRla/NvvmC1EDBbLzi4K7ly+f1HBjGe2zBW+VlIhzX7SkTksqYJpg+
og9rqEZ1hDYrep7aLPESBk1KxrdIpvIbgyDD3h0GPuRZ3eWOqWlXvEBkAaf/
5RjPx99sHZA5lZuNvAhzXiNgeekjsapIMDBVoB2+YS/GJwfvZk/jJzPSHkeV
8IQZOAGM17PBTN6ZR0iDv4nzI6H+nVyUGfSr8T6zht0jMe83FrmldIPMHjov
jVdA8QI7PYRcJY3ywNp5LGWnD36aoBHrs6cUNzJ4sssQC+M0AaDi709oidvR
Tk4Js+ze4kMjBMCZgIiNR+SLoosvEPXdexuLBImitUhtGmt5YrNkMVIEGbFH
eMlal01Pp8NSEBex6M5pQI2EkuSntgFUCqD29XlW/AykLQTLvtG+temayYYm
ENs7oP4+/a0T3QclTw88C2jBh8kSeW61De/pJHrJ9FGhoTB9TV/Ci87YcaxS
HXBbaaUeeJLng41327iv4NumGEJ648dkqxM7DX6XQKtEaQ8Br6gLk+AZGR+m
GaBetEO/bd4J1EzQmVmpu8wq2gQOdV6aPt08eCdZAQcX7K9Ijxpj/P1+cPav
+FGJiloxnHJx4LIjq987JH2mO5Et9xKZ51UiqeWWoPXBpGOWbBKvxIQauvEl
HRRcX4ua/pZit6i84lDI2e/jRJ2P59vq301jzkOULNEWdVrp8p8C7/eZ77nZ
qAMJhZmTKLQ7YHXUs48OoQzXUbXbUkqF5Tjhpq2/mRqFk7iMcZcIIu7MQcsZ
8GIj+dtYBX4iaYRGb5e1HNef9k/H1TTWDZ1wB4G3QHHuh3oYb8CLRI127b4o
yHGg+9ZhhjhuG8aF0FsJst4bq1QcN9qS8AtdfYpR5NyVNYEyjLDVgZIhNR+J
WhQ2nwR9eKAJEKQS03CVvK0FfYE3F/S0dKw4zZfQ1Bb8WV1AumTypGKFsJXu
sJ9gHVo754cMK1XZAQkh8MB5tXUAr2Oayh1x9j8n2zA5P/ty8aErszDtnUJq
K+nRqzr0tY8wpmUBIRScmXLyLSlNrkv5SHWeMw2Fk+Roi+oyEaZDr7Y+Ri3U
AmvMN8bJ/MPj9iW3zjXQvhx7Rataq17aIiX1PgBdaGuJ0pdwLnZ9DR/b7G+G
B04RBsGkVh5LfFMHpWYFQcNd5jW98arA47/Tc2qHpGPHKGKzcJeutyXbXjri
djYgvvpd9/A5vl9g/Dzbc1xUqveX4pv1S6Bfzb2Wi1XzltH9HAcybOgiAHYF
+SEsXwQ/47EXXDwi0Fu0edBuq3OEFXGowXRcRy6m/I6wnPO/5c5WLAwqjyek
b7Bp9LAd1LdT0jm0HQZr1sDDC+G36LO5uDILK6KrcX/ftvVogQtWBu8uHR25
9ILvcY2qN35XPRyye0OQ4fLJ6/EH76/Le4fCKgRso6SVkapc7r6u9U+c8Ob7
5NuvSiYPZW+zOOIoUqaZvhp5pun3i2W7KvMJU5sz5iIqSlyQdaWqDyYngOhW
YQxunm8ZAjx4wE2zmE1nOXKxbHv9garRgxnAgAbtuFnFxpGd/jsz163znYE9
cRmw4PUQjGpZtD/L0637OB8KxAY1C6A+dnwzCLzhds1s7PhiFs7bqiFGXVWZ
XsoFQypEqkSBo/yu998IQ0Juyt+Evuqm1Ybd/MpV8KK+BRrVQZk2hq04Ieke
QyU1Xcl/GH+iUUflMQC0w2reo4ghNKlj2/TycqYeUflP//Bvp1zXM6GVLh75
30kqntW7c6bXP30/tc31S1nCWomMVZuqntrik1FwzZMQ6mHXlQwKduiKFnPz
HN8zBpmv4HBT28Zm7HFGdKa9P87boPON1xqlJnO2CGNWdxNHAQgvQBj2/HgY
w5OSJmNpDdGv2WprTpWckWlIRMC6rK2hrbvrbw/S8uXxr/YqfkI8hnuJkW3/
l8jKkhrLbi/K0lWa/OK6MQGKn6TcEhXQLkvFN0eyTfMuhZ1Zke5zYo8iT3P5
JGkdtQTcud9wHhNWXRkpPkOo9yG3bAAKQiHTpENPoufl9TVuJ5kmuYl+Sx3o
XYASMludsfpQiIUsGYT9rXBlyvpP+TVhyloA2vwUkJWc3BcW3leMA+spxgUw
mtzKD0DJZHL4NPgYib6k45vTh96eYrb9jjWjWXXcbt5Uaz/peRV3HwCjUblP
w8MngjfHHfpKMTkUmKR+pHhuSu1XLM7TKhbK0/uqEQXQai7cykhpX/jYz92l
0XGanIuB0LivspGA/NcgWwAXL16Abx6FGPDCdgRGQP062aI/+/HGgWft1YSN
maau7BTbtVYupEUNtMEnV/iSVNYFONGq2J0qnxH+qTsgwUc6E5kPHupiqDLu
DLduqhbWzoUaObDVK1UiQZehQoH+/hytT+Q829aBLJcwclKVMeJhLaa/KITM
slOcgQHeiyblJx3HlRUpSHdbGT2psBm5+rcAT+XWvs7eLzGJ9V9L5ZPhG+zD
yKKSpViZoeygq+ULbFhr4U6YGpKSbCN1dOhVaPO223TM34eSxnvt8/ewb1HI
D1RHzVEoG1LsuSpFYRy0Bfc9ksKLVGrDQIVXcFlclbE45qjyZEvIsBJG6SUO
ksslxbr34smSYSpmpOzNn+gbjhf1Nn4ZxDK/wZ0mW3xrk8rHsjITERlOUZcJ
BRACuqQwh9lb4hajSobbnpQn4duY81Pl0i8PcNRSb4oG0FyyQfm9d55AX8NQ
/n1v+FeOn4yCQz8YMNo2uagIWP4xCPMOWv1h1xrJB87sRmWuDkPual1FUWev
xuGCx3m2/ZiItS3gAFjxWRfmxdYIHGRetXX10d6jT1Wa5s9U13Yk/Zwc0Wo2
PWQyhlYe4Xwu6NwkhPEzyFxiqzxdzE+5Lv8qgcKVU9id3R3Ee0Eumuk8Zm/x
O3h5A4EpACdnQVUUCpGn6Oy5WJUQ3wNPPGnMBlmclHbaEhNDo9lNCEoWnWrt
6Gr2FtrWsyjXgoSOH/ljbeJAZcp8AjRCwIci0HK+Ufhy9S3HkZ6xXGPd+LBY
89Cag3sjQGSRnePMqO+ekmdKKnP8fQAT2RJGsD9qUw+svUIGibJ6uSV1xOLb
+he9uCUOfoToubrzA/57SZfsFKmox1J43QdG9GwhTh6TqYx3dJunnmjw0RmT
ezEwRhOwGLku3uLVTtWEJjBJ+6D1dkDKnquUb4AdaXcxm551czBDggsEcGrz
1nj0dYCRmIncMJm6PeOGL92Czz/l7uCgaAsaLe7ngqc8vesFtW7aDWhYKYJ/
x+AQC7If2e6ev2FoSKhqCl0LAnCLM17SrPtOJWIL1Xc7oThmF2qzhdo+Ftxr
GSIXzOfsvVfLMMNn/epAYhO43pNGiSE1We+zdycYcf+7biRo1TiHWT73L5YF
oAUUHwFSITFu1EOhk4Dpjnyk0tBoDxyGcA2CW1rLy4TlGNflCj8MKnuLz6nZ
xAHcfzWCEPFwLDCVgkwB/ivhKQ96Ey9gsHoRr3DUHALAL/+07m1TWfZNOh94
EtgnmQfFavmgZ3cttfA/SmFB8wPFeC5WsmFOOxnOD3rCUgVY4FLVesLl6yLn
iaFdqGlaOR3IIopmoseXo41zOHuXfN8LbG/vi95+VXTct27yJpcJjTusYtBu
AgsbauKURgmmbgsRv0duxeLe7alRgx3FvGFKwcwq8TzBBSwRkAMe3oIvcor4
VAlFTrfWW0Ca74wf9VoPIcywWU9dXJfgge5TwCnrwSdEyym868fSq3ql6oEo
GubVEtPqffzsRy0oHUKB1jQtn+KqiO3gjVPqCe2CjWE2Bb2a/bhO0sinyw76
c/d7otcRQGZfGoFcCKszPzx85vMY77tTiofliWMQ9PGYaJ6ZIlk98DdsaKUJ
8B5iNzar9El6KWh+Wt0FzjWPKLyNzoISPyVJIa+OLn1m0pxq6J4UgRxaVD99
LgxEajZFq+mjro01oQly7fpcRdLGFNEOGJxmiZy/CJBGlR6TuZWxCA4qSDsk
EIzvifYNjc4uqQ/n00hcUD9wsm2s6wfXEB343Fb2wciGbc5hZ3BgscWd2cpB
QQG8Kxd5JVJvDHAGUky7R+59UjXmCBAb7VEJuxDK0Yg1lcN+vINpeYoStWWA
nbHlPYLMkWzOClRh48YoknPOeQBS/m69S259yGd3w9ddnygPov8SrXZbUTdM
3WPkyPfAkVKs0M8Jy/p8TTWoh1/sGTD+C6j+qvxBLyaRg/2jo7Y+1ncXHJsJ
98TZBIj+y0GhGMEddfeUay6DvsP74omEfTzCXrMBl2C7sjujs4fpN764iXk9
a0H6KbEEkQGxwREyuleEHnrd0Yy+5KCd1UK3HMqexStIxgMtBVSus+mgVcRB
MP8A8kt9aSD7++OdUHQLYy2hZKhrvjGfbflj6KmZl0JNwOGUJMeHLB8xCy+w
kq5f63hQQ/TKid+CgAvwN92FnL4MMHNZJVzL9p5JQdlHR3KdaAWN/vdJb0R4
lbPKLIwOaRifqeDkVCqtcYpJ/UB8kgZN3CBDeqAZcw25ttBYuZbhqNktbc93
3i2ztdBg8IlVgI5TRXEM0siO/henQ/lzRqyYc2ruIvWlbaEolxYrH6K4/i8H
5sLIuDuwEytUKEJBW3CREN/1VFGmQK0as8KMhm3kb/vIWoQMP3Qeozvrq+cn
y66pLFzCO4Wy9PIo/YNff8NwHdk/VqLx9KE1AjMqU0Jdqs4W3baXN2WiqnrI
ExWkEfEeu5ALhPiIacexMA+dJxVkrzMklHx+vMtqZTRbtEQorsmf3PWARc7m
R86N8zwaXKzTe/IiWnEohqItGmfpPxCWpz+B/9LkbC4lqO+Sa3RQSqXYqOHq
SmhRPHBTEzcX1Rse9+kXQNYUwDGEVnzV60ckZUd13VjZcLP/+w3S6nDOV0HP
ph/L7MwK6mVKSLvXPBDrSZNbAD6yqEZXxvaBinKy2pWDnUWzj4sHgHRCXa9S
uyr/4P8d0DPAQHL8MtLDQHZQwNPWe2y4tktSt5mtHKZQI1gCn631cDSfdoQy
MY3RDJdnw2zivd9v+/aqHkqPf+pqfdVzh/0Fb3U8QLyhyGQlacn6zDQxZp2Z
f6J1Os5Zlf4m8LuZ0sBOmLzozI090diC1uQhfXz6f6RsliCzvtpep8V7wsa/
KewgS0Yq+sxqEGxx7ST++jrKrPiZgvNGnBZPED4Edt1NiheY9UOJA4Sbdo4V
2fhMawT9F+uTjZxXXTePlItb0qqh0rjQ4cmP4kufWo4LCa2astWRqdWCh072
7MdYojaScaFq2x1oD7rqUpMf0O/787FVQKKWlbp1vsreLk40bf/yVEmLeB0z
mPVkFUgN637T973Kqoj1XC1LO+fgdqN2/YV08Mcn7AT6Nktqhe3CrsfJjIqY
v6g9mjE2NxKs0CGSWJ+E6eUsICE8Y+qPcbf32Gp0Ik3rmUwpz7PukoISuhD5
gRy0SGNHq6c/VN+S+n0h9oBVcbPoi0ZMy6YeRqGTyK8sWq8A+1AAevhSbsfO
Tj6scgVFdFcWE3ir6cp1yZId9zKHFtZwG9/sw/srPmfiN59syznCwvMdVN74
6PSIjPJS2kEz1vFIz0mc9yzA/8pzT4NO2hzfcJP2hYm7/0+nD2i+nurMiAO+
UrxiHeJ1zS8Kk6Zb/vYGgkM7FJJnRxtn17NAeoXX9UDR3uBvFVTNs7ecqzd1
vW7XfzsDXhouWPHjPeO9bC0KPHxVmBQnXMoDQn6K634eYpiLBTQRGXjc8ZlX
jBj0n8UNCu8OuPXJMMdbLi+rnsuxfnpN7sMrHoonaVh6zoJOjHF7v+YhUkVj
yqh1voS9sMzCgV33XWmfTxFvk1Z9Wf60i1PcItDnoBFtCnWL5qyK0IKmd0iX
aA1g7rXi4DH+O9ieJvEDhzGx2hp9/8FfaehokM595K6ohAAjkRIANLBHCqSU
frb8qa3IsH2f8QHSWz4AkSFKidtlHbX1bmca6/5De2jtQUjxj6FDuFi7wBcV
uUkQS3M34xQz+pnDQ5pPVITOQi5qkNSOtJ8bzMSmg85MfEUk1kS171Gt/5vq
1R05/JO8traMEKPWJuAJ4eR2buFU63CPUzQ7qvY5QgwCJyPzLan36vwpgvig
Yf+FpOBH5eWV2gbA5OBDMuj7onTn5l4lu3Bk8CkmJUkRPuaRP+xXehRQ3E5O
B6QpdMii+B7u45Xl5z5VII7hWkco7ZZ+YTI8O7efIUZhWMNF8OgIM63XvdJ1
oPbLtyNw95fcUE90dg4TyQHSDbyfIyW1VBh9aP5AnoWvfHelE7M3lQYdcok6
XxPpWx7VtJ6tg+T1ff1wnxTamITBKCNzAstTPcpnZaYqqprtE8XP4fKbGHgQ
LWXybPBpDU93uEwW2URjBTxdyQWc1LMTeofbKTQysHFTiEtZCqnpEIaFpJv5
3AtpICwaE5YpBnaxQlDz2mi/jSGVNNs7ZUdTKTZsOT+sjrIoYFQpTvJmnXPO
xzNTBrPuuiAEtOu312lDAD39VVe3UsY3q0aXCdt0h6BkV4IrJ45ZaR5r3HZv
i0x9q+cnV161qzYreWvc/Qxd7eWwQgdCiXwZ60lVRb4L+lzeaxQlFRpEB1gk
fl1wXQf5xp+B+PGu/mreVKItBIPEV0u1aKVEJNxH0SXYGKxTrCSmXYoXaN7v
xflgdLnyaebmadkLRVvCevZmoQC0/D5U3yHDAUJc7KasPbnZs4Cl8M4zHhXK
0KQVbSGgJaJTjL0761yqugz+zYRlQCDZwRPhUUYpRDZh9IhrNF4CyCMrBS/v
uR+qLyfIvpqI9fogKdYgk8OS1UqePMaai7pAqV5Ya3TQd+ZqjUiPBKAXgJXt
qWaDdQnSRR1sqW4P+5s8kX+TGCrUD/bvvvfgDCJhu1yfF1hHZ7wJEWkweKvK
BXR9DVmfY7qhuZ3tczNMXR+JRBPRW3mJTeKsmdb4guwTRtbAP1toeVSgxrR6
VAaCI3bXsJZD2lv3VBDcX8F4LrM/5kbAqTFX9AGHln3IvXc8/zpp541mcPiw
9fH4l4w7pp3NNOpwhx3PVUxdxxSyAyH20tBI0MwsLE0M0OVugMFl2bNmqcyF
3qm6Rz6voxawj+BY9uo5lzB31Zeb/oq90qOLdCsjoSnl6fgDhoFwDfA4SAbw
/p+elO7N7T5kFHgM+v2KCWQ2hOJc3uUYHEHQILR5sybUABDafF3PmWvQWmte
vLMQDABZfNW69hFqKzuK0lJYI9fQ4brWhQ6xgsdMLKvcE1jD9+V9Xre9sX0X
JplJI/icpv5XFE4m0FeWtvV+JfMBKsd6618iZtWVXasyiPklm6ut7gSyBW7M
HopN4tRWpDfi1D4dd7FdNuUF/ogjAbaFLMKxl8CEdYbrjeIumfET8vlQzpjA
aHaobG9qAUW8tSeHA0wCGaLF8wQif8tmf7j7KpJDu357JLMN9iezGPfJt5z2
MNu0iq/eY7yPUCLwVIwdt9Yjfzk2m/gMLnP2zjNBHztkQg3UsJZaSaInHSFk
BUIMMMuvyIDDzSkPCqKFP2sg09UY0RU0mUu9vpHovX3H9k/pxHoVE8/fQTYI
OvtBghtb0jXsw8lUEOZchJBSVefAYI7xiY7g7JmcYzgAvc60xoVprCuW3zaE
5JlJVJKrh+vSc+0hpQXkjG6ZXMrHqubId7Kyz6B7g/UQ96TsaEFSN3RJJdYz
+n2nxGdDpWWsSaoMHC181Y2lCD5PZcHer0I0fTUHKgzD8VadGLkr0jxSwW8s
amAxXd2Y+p6Bb9kJgcAmd7qW29yvm/15bxB8krl0kfk/VyT+2/zRFDXgiYjV
cd87vmK8sqrF5pHC597vRsbg93EXnyY80mK3D4A+eH2oAtSS9Z2VJlyjtLKf
wPCtUxwI/R750/le0Ykv2kp7qFtSO0xDbFJ/FjXzACwuI6oIS6MrGVNT0Jmj
Y/TiUZCF15/tVkhxYXrEX7AHE/PWQBZ4fjXpEHIz2ekVZ/Y541t8Ck5M6iKe
qFPUiJYVM0DU1G0DNdWOF15Oq/fE7O7uNyWYpwFlPk3PGP7Z+TAeVM8fLE14
oWrx6YRlgLMydsbCvZwbROVMxdk/lK7QfiW3emk/Bdip89Xu1S2lKozopk8x
UfiDsDf6UmJKUR/i48aiponThRe3ZCc+1JbQLnA2hIgTXnylEN1U/nw5Wt39
Vhm3z/Zns1RVZ7uPzv6jich9tk3IjfcJLIZcgFVFE8s0/S90y2siaJq2AJpU
QP7CKrH0ae2RqRWN0fla57nNWMy42jcMPKRCwZIvX5RXT4TpLSprZRTd02pA
6k9l35yEisRCncjsu0C5sg6DJ/dTWReA2U6E6MYIZdnh+jCNnReEasMxlQPA
f4EMM9df3lY2pYAiShJZG8r5h3iOpa7ZRVEK8EyR65HcP1fok5Ly1Mmsl3T1
kr0bcE9yp17L1O3J+CsY46TjRZrrkyiyd3tD/1HwSD4IkpHcrAyeWytZjpCr
o6U6PpNV6cIWyLFcKhvG6ROJZPxWdibNocUoCFxEj0t7beWpf9MX9d5stoDE
b/CfcbSUHeU0KYfYpM4SMHGYQEtJ+ugj1Y6h/xwHSduHnEW21y4q9VlQ4kb0
PcMHHgjRyi9xlD9VYbNI5a/F7TRKj02ccla1fCCFyUgCU6AL0+/SWLUjvH7C
1a/oFEx1t096WWHpaaBOfl94CQBtc2uYqIExiLdrW9lMPHwnlo/Eowez+C1a
5axXqxti3lYDbuvcAv23pmNo9nJ7QKpn76B+/QxF9emCiUuZXdjsEKe0i18r
EQ+re5Ax8qEsBmLMHUmf3wlnkKt1cBbYmrmmBlMO9WnBGGv0pjYRuMUECMGV
+rxhWGrioLPA5erbOHk/uAa7pr6h/asFMSC7KP5On6tULPtP11PN+7OgnyyI
lpOrC3YOQ+UutjVWr4oPFjuIrNPzynYNzoZ0nFXy5W0JYYXr3up+T7r8N+AP
ngcG3r84ixkmqxaJnYei3BIkaIOwC5H7wt4H039ZwLPi98HAHJhgPXrlNgXv
uu7j57ENs8hYdSungcK0k7KN+Ci43jSW2E694qQKVeUWNFt4qNAJIflVsNJ6
1ozLbtdsEPZY34wAT/fVUphbW9cfs64ZtUTwG9c0JkAi72HgKhZicns72RJZ
coMnRADitrjdw2ngBhPTD7RF7Mit4f4NUMxHgSpfPFmA21k8iqXLV4bZCLVc
+ulO4+4yHuFYVyN9Uc7LtVRk4mTQSru3DZvicYa4VadmTSAQE/rSJo5DZODv
ew7KdfUigjynyIQenLiqrPblgWXHq0gXFLheE2eDol/8YLr68lYYwfEvZdSd
n0CBKYO6jA6dWlWTN+73IVCRAqKNP5bpBO+9JzqTDHbPly7jxKMX5cBl1fDB
dTAICnCY8zifESyNEPYxlOPl/RRyzY1kzOdTpd0Z4jhgxqMj4UzpyeWAtpA2
AQq7gKDyJt6dsBVKTTnxlXASLU0uBmQRTlShO9zmMnoGIBvfApJ3XjCwM+JR
1h71yQsS2Etjr7T0HA+Vfh4gaXPtsY02Kj+/UmlLC/J8LXb3ALXrnkDA0Sgy
BoNlLeOt+6fn40pjEfxPc9vMaruALrblKlfexpGlSMjTWVCHmG4eEv228IK6
cenHfyqaLio6u7qD2lXu1rIjmsZHajFZzYFEDjfFvRZ6io/yhkFuizMFDLGw
cZhmyM8QU8DM1dk4A1yDqhiS+OQeetLRduMVAMeU6TKvopoJKn69zjoFBkxq
vKAgy2gF2i1bh7Qz7Iq7nyxC9suxfcVDaH0Ix6vL5wWxaoNhrJGnRa+uWIAq
y/87IfTXrWoIfufh+Hcrm7qacyZMQuOnbHr29JUGXPWcTcVksEAX3pNwDUPV
fkGKLIoTQVa8HliN7mBT5/8=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1L1WQ/B5p77enC9Y6j4cYfDk3uBioT5K5zl2N0zjlBjqz+XrrUxi/HC11Wih7GLv+2PyxGG+rKibw3tEsgaGBsaI/UkqzTymqkXsk8JxFNBtw732EB/kHzFh2SzFYSELR855vg+Eu04I8O9Z+R+dDiBzqwCIZSBRS5NA/IA6x1HPQXGXtQqAuCp3cwO9MB6Jjsg4anV6ThzttKvf9vKjF5xCwniZ0hoqW+0VDDiNi0kIeuK8u4lmsIxxftBweXYLrtpMAL9ZMz/VDWEUIIwO84OFe6rq/8lVM2rcTBjm9AC/3ryAHdOeVg2hs3en8uBRQF8HnhX5evWllZ2P+3Imt0HfXqWG5uD0hLZZhJ4mqLwxH1WORkBD4bcT4MskwG5NyCw82FOfPJpit9WNd7Xxl9Fs2oiKnTO/dxudFN26Kn16+6EynZodNW2bfoGyZ5clQZJdF7Sbhp4tIXesehPHuKm4DT8KTXFkDYNJXedm+Oc+FwTIm6j/N/VJ9eUvBRioxKSrzN7+Ey/kM3FGZFwRNjJi8a0B6H62+EKdtrRM0HHiBeDRvXkFGt3+cpcq/wiIdtFr2SBirRM8HICAnfbsepo+yDgi24fOs/LvNC7zilhfSNZrsWTe+r/CchwGDhEIdMB4IvdcZJ70yFFuQQmv+SVCNrwbKeRkel30N6tpPk4OuxWv9HusPf1AGJuIEPlA+0ohd5BUAFiTjzRUn59NCL+DgprSKt1BaBzH6hzdP93NpTMht3hmuJZNDtgCtQKCxLQnsJ3eoFojgvOR2cXtukf"
`endif