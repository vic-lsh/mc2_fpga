// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CzAI8XObLd/OfWI866Lcq8UPyIHuMNi6yQoojwseGOI2JyYrae9+usRIXsZ/
rIXj2s9zHIhF4RPCkUxVUnMr3d+Tcb363UZcOKCYsgckVPJEfSIu8ACRr7ry
sHDVLB1dZhuOlmmLHecPW6vRTFnXR4nQoWk8q+1X+4yP+tbb6yvCLiiE4nd/
cTQYldK+QaNuVmM2a9BQGm/HYiKi7WYsyOc6vPyekHMZzF2GjigjtaNcurxz
nAUv7mLiHUHowOf/S0RTFtyv5u8uFZMaDAZiXe1HN20jpQvQuDD71xVVZYx/
l1FqphZCLboymkBBwczA2v42COqEdnzYhdPyAwRytw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C385OGT/T2A9hdZWoab/5XjT1c0Ujql0mZ8VqVSXuGSfWXw6oDg0wbJXQ2Wk
/g7LuCzIEgF+k3j7JMIISls2Vkh0oyWr9abOCrs8dVPQ0Lo1g9GmPBf01UDs
cTOU25VEAB90f0MJBkyn0oGUMJStHM4glWwBEsv3k+E+RuWIYHUj0XjS9/JO
OfTEt4P0Wl67KALTF7ogtzVddyISKU49Zxdd71P6Efa5RpHjSPBw16mMM7on
yjjnhBz+P+GpS6u1G5hmKi6zrAWB9ld4p6rVeUI5YBLdD/OfRPfRGRbEZeCm
kd6fEeL6eKNIQr1cG2CZDJQN7qSBbbUDvy8wxqFAqQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OPzblk8XHB5L0RGNpo2VkpzrKDgS0MdyEKfkUebGs9OfbxXykZ3RHlW7R0bE
Yx8HpZvONx5N00c0qYmvnVR15BM5Y/MQKFL/Aj51bpTar+cv6e0go44ShHi/
Venfg8isguKb4yuf6sHel2AiZ1jHkjsT5M6LbXzkPXzXCgbYL4YOKesI6RBd
HRWhvNeEq1cZZMbgGMSKs4W1wASRia+rBDXpNiPKGZRLV8PB9Em07t/LaKao
seS3BnNKkNgQ8Z+HENKhR979+aqglv6uQ+0AOoAyJeaTXv75pBtxWFSSZxCL
D5cBeGBk2PFMbzzAJ86nfokXwTqKIxXqASJrfwU5Og==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PATw0FzDu62gd+eG6LTQqknmthUVZ3gpZ+PqiLXSyq1qvbm/XiWFy4/VmsAQ
ixStYwVPUrUs8Q4J4fguGIXal8KBXA4aL7w6QexRVzJAviLngbkPc2RT5fPy
yzuUu+Oym6FwyFRxryMZM5yXDf+5ogFbYipFBhVzshR4q0SheMsO00kqrGyn
aaKSgzVMazEoTOgJWb0qS2cCcaGOIGfWslStoQ+CZ/LqCfxbDsgHtfnSwJgD
fwzFPU+yZrP0exSBJCmAGtwn6Hvx1bQDYxFohXuAi2ZuvpSCS3ZylwTdxuOw
8fiBu234IzehbYLr6o5Kcrbpeql99oktwlhwqA7J2w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W9xhXH4BZDYVr8jLzyX3qJg83gGzftjMhYTlEj0retEushuYcBx02uTnuoyZ
EctcqcFcH0Gsd8ByhVk4qPa6GkgWr3u4xNJQ/l5kQzdkz7mlq/2aUENpgPB3
7ITYohB+j7DHp1sRf//xdnH0yEYJZDvLqJzsd7k2f2qDj6aboJQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sVkxRx1XOVORjvYtFcMF2bDor886UxQ5wyjUGwZqfhJ6VQKMMNEnBdFYuNkD
ismMfHqkOkWMX2yEy+UoQ/QEsuLT91cGvd+eLS5tBaHYkiM9/+NG7NIekug+
yk+3/qdocZ3+O9iUYXEWOu+ozLf0htdUkUFyFjDgSPAy2aRLzMCYuKE2lhKH
Qrp5m89ZuYil8ub5gZYarHmTpraGtuuGrx1lRBL/+a0KOgtuemhgk7EMNq6I
5pACdoqRPFpeV0W/X8UDwTWa4MCo2oN9ufGAtwbIyxDvM6mCrk5c2169Nxtm
NVO52Z+oZC15E5YWy2uyV/h3iWQ2cLaCjcGQcf60eQwi7BiG2d20//7ht8zW
+atJLRuLWNEDZg9nCaoCN1q5XRS9JRjFmucU/x7FkZMR6v62xFJod3VODtIh
QdEmSwsuJaGXfj6Gw/ZDnHwTmNHSeoSC93pkhbcYjwTSMH6IXVs2puo+q/Lq
SAgujKMkzuUypbpjYJ/Nri6BopdUDroZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qDudO8HVBmdZXl6Cyz9soX7AgIxpwfrQL3+056tpHU3i/+bAXyEqZyeRLGN1
PJ/dPWGwq4XF7YaSUFZQ13dFxtkGL64u0SpUGsnt0czBHf7gldfTBdV2z5L8
bmW3dMcPUSDwziqWN3vLRmY/SKpBwAxxDIddMuiDq4vpF6d15+8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UIMtXdUxWs7S2D6S08YWW8pmH1ApN/13tFft4UWbu2ejDeZ7ZvjSu0pt5p+f
dIya/IPUKFSLpzs+xEdnTux5B8QF3+I4hK2/rRxg362AAF8Dm1rPdFX1Ex8W
O8l6Wyxq/Jaf/GgYkqYYTtcvo0eBxjgIzq7tiQ7xgWS7zD5yea4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 71360)
`pragma protect data_block
0bTIbCXuNJTthQmFg5sQFkBP8lAZ1Ta84RKHiGEaxN1/NIn/VrLWkYkr2M3B
sFH499KtcSwX8N70higCAmLZPKzWdofYpZGsajB5/PZXnk1eEC9MH/nCFjZt
E8nfdHj3uiZYe+QjYikFhyc9Rw/PzHD7uFn9F/w5fRO/9QRMW2du0u/oUKL5
68uaB3AW23udFzTPeTuT9Xk3L7L7VF7m8TFQ6RHxTwO+9wuXtDueeZAZrs4B
+SjhQLBC1QCbH1nSaMW3A5mI6f4eb77QAVZllZmr/9w2U1FZPwfuRy1aaC48
RkqnQDZFNy470xxt8/4/oodxsJ10kNFt8ZF5uqCXwLvBrBkShuWLtIjVG4KK
DxWTXGm9MmCbj7kr61arPRXOq4oYhIA4V1iAq5LxcjaioiPEPCA2Qo/ygTHu
JoRYzk94gcTLEkmOxO9/Gjhf/G0ZOAwavd3jzHdNzgCwCXAzCMrtIxWBcdrn
xZdc0+0VFb7rKzMxfjF5q0fEjg90Gonxwljuw3ZH1lKhToiAnd/U5iAKB0mb
J5isOTYgNs52+OfcjoH0ruR8d19LHY889VbLBgqblMqQ9ERI8RJ0huhYMOuY
fdC7+C6ekiFJEfEPQ7VceMZbppmHbKuwtot7O2yYZ8rLOcQ7U0XvT6w/XMQb
d4vYQAYuZaavjPlvxbRja1bxOJFI2vsiCxwZbXHlXQxcifzUHLUcIkunk6Sh
VUKacitvL3/ObhSskKcPYXTkbUGL305FV+tkTYIE5dcKHEr1ZCRfhSL+XEv2
seUFPPwzQ23betEwnYsr4D5jEUwzJFvza2aQ3apiTT6x2flyOj95kx8MtXgJ
L60Gc/bkSi+RrU//HdPkMS0XY1y7BO12iTEAfWrv+2AW86zG/YQoJLpcWEYP
WgIFSAbGufp+qCHWYePp+BbhGMJMWoAPzSOqNub+mpF4c+IxoRChLNK6hg73
OOgAYM76OEr1CR5sKjNStApqYu0nqU9xLuldY2kIVpwmhIZ9TKqlO1YDpYDY
J4SFUmyveCJknCO7ZoolVznMybGhyuOzhROeBKpXAbBTHAmM7eMC0bzU7ai5
tE5yuhD1/XGYpsRJYGUzX6PmZOWgfwbo+o+snIjEjGJDa5T/TAwgym0enZGH
mNZaRGlAx5TvncSDsA5Tt2d4SOFWOxiAehYCGab9TlmTBq5mEQ3uGlx7R/s8
j++65xtsy3ihV0/lruzPhEyV1bgW4nVUvYeXhyxopgJvaTHF7Fg7OpTjlAsV
yNw4cferOLgQHmejgZ72sB5CePd6u0bp4bPNlIb+Je+kxcvQ+mYIEsBAUCnV
/6GneErEJyPSovpSh883xQWaOAyMLfD59tRRNiMDygdGSbt4/59UpspPZTcY
/8jKyJf9FrKUN/a27Fec2kJeyFisiU8gXus9VbXNgxv9qkeXDBZk4UzxAbNU
OR5dJFEtsHw0gGGaBxCinnXq8o5gkRLAUfkEUKCH6APcd9XpkRVedyLJPOEN
3QQPNqJmIsq+IGkBJL4bNLPbFWvaLXgvy5Qj+Lfl7HLvPElRxR5s5+55S7fg
8kyK7CYsa0fUVJYBHFjQcluvjs6jokT9cLG3zIulSDz+Zg4Nx3pa3yoL3kGM
987lgjL/p2t/6JvKfipyki61cCGqgpNyIOUOCZWgds9PtxyKocUIKXl7Gaar
BZFCJ+wcKPim8cEFvWDMGwQ3JTAap0FIhVB6LrxndH+hzLfrM65nuLJ637AQ
D0O+INtzVqdFDqkGX06OpunxTCu74Rb3PPdUmTWA1gnBAZefrcIh/+5E0Xfn
Yy9rFzXlWXvk1qgkYwm6oohLKWrVbl/1RA2fZvRTFa+q1iTqC+Ozxe454Drx
T8kWLpH+Wd5ueFDYHXsygSwrLnU7x6q7wdcUGJq1AQpoX8KFdrV/yW8Zn97w
0rj0FJtFqQ8DhUScGV1KlTbLe3CCwCtSHwTsq4VVz0cSjytrq5X9gRQLhnv4
BVrpAqkoKwX/gXMA1b1H2kaoNl1120XRC5OkSlSGfopq/75rRCeUl/EjM0WM
jhF3CjyXCRE6cCBzI4IGTaCw1XQQyFWmhOCPo94Kqt0kBKRvv8LxwL+NX2lC
+IoUGo8EjQW959ELhDyDsi0wK7KoQ3QDR+Ps5yoNavpooZj0gYhaYKEhkThC
5C9YvmlBPppxoC1mRccJipJ2ZRXPBcOGDu1TTdHgxUvUWJVi7PU0djSRgZfg
5IW2ZPu1uHwJUW76By8DHtTDfHoX7gRFGOY7PT3BagM9LDVtgwG7eq366nE0
ztJ7rmNsE1PTo9hwGSmMXsN5cz9vcGmHjFwPkrTKL3NC5ON6bWY/3LlxU6Pf
46zVQJJyMAw+97kbYr5a91+HMSypUITIIwSdfFPVOBZ/aB1VIXOFAo+NmADp
C/Q8k5Fxwm6L9yQItNGo52Wzrvq1bOItGIPXClfN1uSVPyLgK1av2fTqqoYr
I4xmA43ssRympZQ+e5CYSEaW8tl8cLc8C3FuZQWqEpubOwtPHnvhoS/Dekvn
azOEdR3tkm9K0ckSTxmmgi8d2OWmuH98SDePxTDmKRyLOJra9WfQk5ybj1lk
Rw0t87/sSUumUcc/FicQwWi0siZVyWm8qOVerwQWC6r9Y3sHnb8czxsvTtTW
kY+1ys4wi9qA6nARQeqmzGr98ci3/xPePoFx6iTvCycU1D/qHFwGsi/DqqBD
CIk1htamOS0jvzjBUNQvW0bnGYm30X4FqpKbbwEWDeAzVpJZwXOVboJ48CCD
e5qZF50y1QMyM3Wqw7jkTQla0TGCtyfhqJWz2tbBIZafTo6ZIq0MEgrd7ZMI
1pOwKSYqXduA5jcjIpxk/a59/vku6uoLN/W6fzoDIahCyJj/drd17j65WHfp
jx9rBcAq4I2hwcalE2QtkKvgJdcs88w2980PP3QkCGxN1ClJgWv3AG0Pz3zR
Oy6hgqJXzFk6ixJfuqGjCYDBI3dgKdFFRGeQsYDVcO82gFdpDUy50JFc9xSz
EE1oBEeJFU0P5rnwtJW1IF450r6F6JkCH/fdCPYMKwv4VxzGuGv3Ji0vU5wQ
G858gKeD4YClRqaDGtN2tg7vpU8IyQD4rnITHTAuWolrJ3DXqfPjn65seOBA
uUeSdxkUOsCZ3W5l1x/97H1v+oK9QTlctzoY9EarXBIC+YIwO0prMGugqAyr
uVzY/EIqi4osHe5BVbChaP71OHK0mjspWwItfNr/ExS7Xm+jEGRK4QJjNBtR
MU3TwCeiNaSrW1FU1uJTyxq1dfmUduFAi16HmRK0GJl579rN5PIISZaFnl5B
CWHjR+DX6yA+y1weq5BlmsFAbZp7zHpZn1PTC1nUz1T2ANsMm0UWEDTooLRq
atJsrT1gKeoX3LUKy97O17FKlucxRRWm8NXGd6a3Vhm0hVY/iPh3ZaQoQjdY
ItjmNW5yJ4omgyUU4YKUfB2CLBzxbuRZ2S4wnukSuXnEt7K9IuzeWoFyy6xR
KxUVlXd/X3AwoUSRiL5uFqKIx9qs94/A3gRGhiwvWj1w9sqsASC0RL0dvVJt
Twp50U4aML9XVW235N0DMezGdqoW5c1861bHJRPYpxIMXCUYDMDDmfIXsWtZ
mFokw6NBoeG8vaxf369U0xTCARml/my5/pzOrjvg71kLfTbqQWFPyctEhwNc
GWGHiJucWTqtHWiCuWn2gt6g6ZjjWV6861ATlWyAr5eN1roQ/zw7Ky794uke
TKTZZ2I47bvmboIrqJwDSnFGxXCOFu7YlF9s06ysGVDCFY7JrKJH3NXDjcJO
Y+P/Tbh1IZmwjcEeWCvF6Sle01DTWlOpZ4HIoiNIjio7AnKJKmTFTbLPzLEI
tdGH0I3iyYXWg+fcQNdjcby20pzXAXc0aAtBJDf+gIowXndQVeyptFoTVPmA
LEoBjz0NdKGnk1E2MBVVIRn3naYY7fxfrbQ7bApXVEyqorbjowi4TMjrZ4SE
+Iby695ACN5M8lw7QWZlm2LdffqQyc0txwM/tdpkFTb8q1VCTLlomtdw8b5d
j/T+3wBmP+GHfqN4pr0SDtRJduH5yy1JF28z+1mFUFnThaNxwNKE1JF3LINJ
YDOFQiF9rb3I98307pE7glZyTKoymONQsvR3k+D0XsZBc1G+ekq8PPsDVKx/
hGPKy4E29hsByC7idamajWIBeczwyys7wpkb1T7gLGBRglK+d7x7qnsxVQRE
rvc9vhJmH/V3pmkvaCJ74NUNz+0+WHVtSHG43BqcCWS2gY4qm1Q+QbYT4G+6
8jeRPGNL8d7frP9reDpId4eybY2lzghq/ilZUITn5DkjCxDh27aOzn/pRJ5r
TSWdM0HjJFUmQ9cV2QsIGY9O0A1DvMtk40oXCLhgmFqwc9cJhNb/CDkMh1oz
2CMRlyqr16RKWjqyO+ah1OoF4OzFsx5A/va+GgGAK7cNhwccVQvYluv92gVY
4TCA8N8woD8o2OIapBeQSZBdUnipdyeGOTpBOFp6CJbCOzELQieNFbmqZGaA
A2TykRr8SVnB6WdJY0XiY+bfDQF29IEpmo7iwXwGiwGtU1Ba8ZIc9iPT4s2I
4snE6U08smdmWUO/l/0lmQ4Wk0B6I89x28EOY5U4K4EyJkbH8PmE3lhlRwBd
ZpxllNoyk6+oxFheN/SciAEFbX7/whG98Z9gN24LqPHQSy7CBCWq5F+H3HTF
YkTsR2hMTr5rBMoE+Kb7QOutd938nJKe3GMxZgXzIXTvYGzu3zUcgUmVGiUI
BU3+bTvov7r7SAn2StEDcvjbiGoUDAjR29onaE2J0P47Ic8gfUdZWb0uK2jP
vrtv8fS7zd+rICCqyiyE3xRwuzuW+OKdwKcBaLYgZ9pBwPl5aW2a2FXM5SEB
wf4vIH6pvdBIt6nQ/zEEawtQ7VfVA+BpH/+tZxwYWiEZnyfzbFAsdsFizskc
cEg4ma83+OiT1r/8hOnLMYpBkeT8jOOORZiAcfeeZ7QtUYuoqnbKtPh7VRE+
a37nSQKNVODqEFhQzxA0k3fBRUijpb/xywp0zeHTABpNTG6olRpmNWHI2BCA
8ZsV/CyypOIpo62i0IPU0xbS1fnqh/QUNAEq/iLKxIE7I0Kw0aEHwnbovC20
aHjuUgTDWXkwe8xJuah7GsTcrAhXdMSumxieZSWlASbkKLKMOO1O4oCHaoHo
IyyhdlCwLRK6gLCJ4FKFPNV+QhUp4cbvv/Eq8lsVo6YHE1qnIZnjTMEDJD+D
nhTu+ILKIzcGvX9UmJdjEOrBVY4cGBWp6gVFMR+F4Io71mjKU98VmAeILEPK
iVRjre2P57L4OZvodR9g9XQlGwyn2diK0M2+qv54OUblKHfoe8iCpcaEsHR8
SoifGhDuP/oqznJCqhyBoIZdg/WG+CdI79EZiVcr/4kNjH+5TRNzTtbYZkxl
vL4scDVn+Uo/WTquB6EAiMeR+NQNJB5UUWj1MLOfuKBA1+rTkN/kGx//B/mJ
/eSvlp4DsAjYGcTQut/fpLH0zZxkXlS2cf2G2ynAp0R8UvymrRTlzKfCIAcF
6lvIk5ueLqmD6wXTm+yEK8Vg3iuDRuTDcqiQNMjvZA+yzzOgzMJ3BxdN2NNm
8nWYG9Htl3k/ort4rP4MYfAeazpFZyrcwb+2rwu2EjF5tx4BwchZpwrPwQyI
haZv3wMBr+SNzkYhqu2jCcay7yRqAfWQlGcEhiJc++Ha+VOAer9gulteGpjY
Agevw65gyFnxv4gdxqYBJW7ZPF5+Oc+QEzaM93I1awNdQqbNzD/EClYeBoNs
RQ91SsdTrxONGf9a6IDJME1RYdYSGMTlSWLwNO4qz8s/fQ7IjonSFv8321Ac
x56e2fhfDrzZDhSpYRFluzgrNS3nqvgr/Nxrh7wrGPWtrLksyIq7emcRbtNJ
kyeZ+003D0ZSg3CJdtnJZKwzjlNWrFitHUWl3eerySgCRst+1YpMFOGxPyVm
zPtYFoFB0AP4DJlqaoO7WssvHnkHG3WnQvPxlzFF+aAtULaHdyccnt96G/uF
/bN9wtRDmULs5M7z6TehqmcH+WRejumBx0z+lmiYqKYrmkbrJT4xuKViL5vI
mxAu1XWrExrlIfH5sSlALCG8rgrMDbh+WSq1otqGP0CxkcYIXZnIYRJk3Q9n
6UruID7u6K3DGTt8p8MzTNwW3vySohuQuWeoThkpZTon0AUxmAExTdmYUHSq
WejrcCaHE0/9YxcPkHiD1wvowJL58d/vXG4VT0OqfBHs7j9ABqAtde243AVN
SUhq4wyibjpvSyn904+4vRX7r15xKGbVj7xLimDIP4lEzIrEmJmSbwBVHgn3
63sHYciPdwDASqophnDRT/Q9vKQXGK6+Ogz7jAWkXD4JH2L4pc3+VJJI7vWS
HiGFQqpjaDHLD0ZG3FL13eaWOq4gDCDD9K8uJ8bPUNj9PpvBZOkSJmJZ4LS4
GMbSBAsvoNdIrTGIXE+4pnGs9uFssOf9wR9FL8G9N17VtF3/Le3pIrUta552
elsNK3NAm6iQf91YYprrBPu3tZJmM52AwXWcwUOg0Jh4Sh9cle/gBli82UKn
Mh0VOHnGVVlIduDuMgx7ECxnEGfFwWOcWBVmhY1GHDtcA+4e/r4ktsCkp/ua
r+UGaZU5QA2e+a/KtOrQTZchGV4BOQocIiWqGNRMhuS75mSpmNoRJm6mFTST
NM71YgbBqVCF/J+PxZwyOsXsbLX3Vc26jyJGthu7m4YY3c3RKAw/2XT4fShQ
z2yQF9E+a0LAr5outmR17tsYs0d27zGuGEP2+0HmJFVmtuOExCAU2tYshk0b
AkfyE6koSe/qSL3DT+3AuN4B0iuDL4HETruqD6Kngo2rgJhernas0U2v8MeO
DguhJl5BtX4nRetia56No+ymnGDRtSCqnqhrMhdn3xXCjVgx8gUX8XPKpTqX
PD71jkERibOPVLif60X+jlOro4hyOPYWQIS0iOvHIjvozFOJWSypDSQ76C0d
kxVrJfVa52ukaZOWnGUvp+2Z/TXZLj1+fHFQ3SNDLzGdI/wMgNcSrEU6LVvu
G1T2L3fJD5hc+XpPhCGFiUIO3p3o6y09wGguX9541+UaLbhtjhixrqYSMGKw
MYZnkAHuZMncpyHNmVdM6P/VOEIrORu1GIEuSuBRKBLa1CsuMD5G3kRtKKqM
x2Q66drzWuGp6KMvG+NkJ7oKTOzsB+TN8RvV6aIq8NfSpVTU2k0H0bhoHE+y
jk3htXZXVf02Ph+ekn7KcGZg/EcKXqh896hYarZHg8v7B+u3mScYTj2Sa0Wt
9jw9CoLQhwH8KaxESyOrHyHeVfU6iw71ePoiyAn80v7+A+a/7cgOMb7cuMtl
2Q6tDXQ/49Znq/AvtaSPaJ0I1MeO654VOkt48ri5L9RkKRNg+9e+67BsE8ui
gHGX2HeC7jTpzS2yMfJCmXO8nh3ir4aYeERBQx/UK0S1oXlw5sai1nw7LBie
9xFnO0mYjJCHGciQJNxb+TUr82ZbzowqUZAV7NFwMX/09WkYhkksRh2W6XxL
BOvYUbXEHLFHAnhIj9b2S0k+PRyHgt0162agSU4Bc91cR4G5Z+XTwZtxbACf
MGaiP7zxQ9puh8e/bMUOD1pvSgviIS+Yu0n0E7DXhYzu9IVr3/tpgnvWXurW
iieEGgZbzrx3FG7STHd1i2vvYJMytfq4OE2aR3hm5Wx9s4m4lCC/J8x8FUTX
tOm0/olx41Ka3vIcXt7DDdTSz31ACnLzXf+OjIqBj2SYlP00b6Ev/Oq8HePb
YRf2BETpaH1wOJ8Qffw20gsxCfdhevJ6ceppa0PRuDxSTjPuPGz6v388EjEh
uvIZsjyPuhj2EJWmdNOYSlz7sqO/6d8Q0hWw1RLej24fmjZMxL/ARFfQp6nK
bNHQle7ukLA4P97Ka5JgyMa9NEUCybVN+PxS6O37jdkPW5k6M0oDfL+V4Yt+
fGEM4BoxG5NRrNAQJfBYPXat9/jeWdB5U+hvM8FEHF+UV/16u/ayRXfs+scV
soYmBEMl/1EAHwvOBaNjCdLXzXVrPyuWIpT0sIN2klUgu1FapJjmUC0cr2JF
455nxe3OsIgQHTTqnPdW4mujr43JHJkbpYzWxHy9YYEsdl8zYQA+hXLbEp3i
5z6rH2hqGsr+N1IcJQu99MV05KhJVlUqVPNVyf64BHfLbrAp6Z4WrY0mAAcB
olVETqiiAOmCgqtm3KCgsypHlznAAh3ghsJcq7YylKw5vCz28BoNqHm0Y7jH
7TgohABa75SJDv5luYcr0otqQS5oPWUZQYnS30SHLXU78PUFq8ypuZN1QdBt
fUPj23NwxxVYbnyDgM72VzPW8lncK1MltxBwZvfZLWd+knv05VtE5z6KEVOe
rS+pTQaLhBOdSaRYvXCO3AVdUH/YwyxAQTmJ10BJp0vuHJ6QkuSH7Sz3xRRJ
d5HAIMg2VAa2gpBZrLK6tiTZg+KYwSdR6aOK8kpuK7uS7OjXB9yZbwecTSe+
anrPv4cvMB+beZzS/RtyfrdlBaGilTR2Qtgj9TusulPhvaqO4eO8zA9/nBce
P/cn7gJkgP+ViftjdC6/Fai0V74ELteMsg2+wWTz1RnDfmXALvda6zAVQiO/
SWtJQdGIULdVEY/QKt0BbCMwHurOKfmj/sORWT3wgsHF+/MjNrI90Ru15O43
JkFi1vkfjcII3f3ilINpDzrU7wfD0D3UpUgij9I7nrhniAHGw8qOZi2JhomP
+BrXej50Y0JBkjCWtpEEv+mBErXFCHJOV+F4VBQ8MLi5w1w/Z0X0xQ9bkuEY
C6NdzPfO6BQYlrCPNK309vTLA8MTuk7hHQjXmtPjPqe7lwVnhRVfpbX6RpOE
qZjbEFcrfUM+rBIkWDlDlmNEqT2SqEmho2teg6Lp30rJ+MM7ZEsWkxgvA89Z
P2J3UhvQVki05Inq2O+adtwumbTWDezGAkoXgRSK0DlPvl8W9X/7idl4jSeU
XU7+ZavpSvndqBeN4VZsUsIpuyiESZRE3Ob4//XQ37SMaDEIwfG+Lyf/EBNy
ggO09dc9EmLeozeATydq5WFygiYiF1/z+sXxxNmF2iBAfrxXtcX94IIxYusl
1wfNTehO22y3wMTwczz9h9feGNo8qGdffI66me9HDp1BYe01zegOlnA6rVva
LtXkRxOMPtHazwO/JgszcM14wy1PdE37jPpFrcvHsZF/cKF+CnB1rjmVi/b8
okLdWgR5cCJ1NgfrtPQuK2UXsB7EL0tSE/FMvcbiLPsoJbUC45YwayKWilze
AlnQS15PvFjyT5tzm8Jm582qbEyc3PCGmgEUhMZ+fPx+kLNe53dUPKObIpHU
wnZicXdYsFAI1t55mnwMD8JnnsEMj5Pexr2LNac62WNHurRAxRgug+5Hk2CE
PJq7Ffzh6VLxs8WH5aj2Rqt0CvvaX974KY2qa0CqiJQ87yHtk6j3Qj4Anfxx
CboCxIlKTfRMFzpuatIfqGCouh2/6vNIrR6TpIVVZiN2HIxjbDNUaTJZxif1
d8rQ03cRdVrfuH9TTiKMX9Vdqb4xxYePi+HkTQgVw8+Y9UgmrtlxXZD1lpo2
7Co4kL1FYB2jAiNYvvIZs1gHGBDhV0DogNMPtDwySCY70p90q2/8fF235URB
j8ZLgOWLl/bSOsAYDA8Xfp2t6Qfjmuy7qGyz6CTH8+wjOwKHNRew5rmWW3aX
U6iyiHd8n71H9HkXEY9VrcVAV5ODVEO4Vzv4lFvDi3oxGb8MOZjS61x+cNWy
TySiIN6gPPQMFlbREoOsCc3nxw3VembL0mczf56IGJh0mEps6Qw6l3ovGY9G
Tx5U6bBMj205Gwmw/HQ+FDj+e8NJCTUpNf56df2ZcgFJMSn2NI6KZdn/f8tl
8GT6VRpln0hxppHBRR1TZio7TR9swTsg6Oc/i0PVKAJ5k1RmzqanosGce19q
950Uc5e2KdVaRt6FKRtgenqcXV/5SV3J4/pRCzCdtTWBuerTmk+/KYmNL9BV
npUP7jmphcrB8azehhJhMLkCDMlSeaVoT6dpofv70NkAQTtKApxVsVyk5s6S
tMsK5vSaDKga6SuIovboqaQe6EmZ3a97jYX1v/PwMKf2rezct22W1+43HS4f
VFyQtDV8FAGA4Q+Z1wov30s8yd8iUudMEZ228qt0xwC2U3rny3wpaPy/y07i
X2GkYIkMEFt978ISz1JciFv21ZqWlMyTgdEKR9KMaKmQIRjkhR5XHVg4i0vZ
JaGnIVxiyEOFZRjCQ5yPkE3SpgdKZmbgJ+ZBVesP9af1pcQZskYlQ8/X213r
yVnAyQYTqHNPviP2trX8vpdiLBIjfTidYMCUWFv7zYdRuNYSRg3sMme2SpBx
Xlw3cu7dzSZIhRF1ggb4RZViL+QPMtOPbEi0kZn5ZmVANVxHIWnosUA8pT2G
RZoNyL9M/ysYMeCw6abeKARq4SpDrtjFsXCoRjYyu3EBe3ZyGFaoqMkqHQxb
bbV97Xf+kTLvviMIomq62dyN/XQwmCxQxZFjpoiO0tO2qwQ/OzTHZosvCvt6
molu7OKu/KxK40GWyZErxqsxHwJmbhbgxWy0NGfOyGCDZlq3V5Vy0HQ5w0kr
+Q9Ug2JeUQHBTJ0TWITERugvymWPC6/8bXY5fJYWDoMHqJWJ/ggrNv5qe5Z/
JwC2l6h/H/fYJoYFYne0HqALZaQ1XYRYJBlfBzORG/HXOUKfNrxA0rGXw7ki
ag+ROeVNVHJ8rZtUbFn9CTBrDts2Q6us07wvy4uxuGjHBCEpI6feFbIrMoyd
n6kD5DqWgC6iRRhgcZ6QoRnoME/hL7rMjJEw6HScQJJDuGflbktSaAn16Bja
pHpPlk0N7lO95e0bc8XRxbuD14Dk2JaFDEiScKprPlyHu77Sp9Go/jtNle3w
IY+ke131/ehmaYbSIqhEcOgv9z/Fxf2zqXXC62RAjzB3qydwwRVKuYpS24na
p97mFqqy2UIq2GwsQ3ve/FsyRrBlxAf4vjxTEMu2sEaAaPH1HHkEzgWH+IHu
daQli8FKsKdHqwK2k1Ppe/wx4a6Tm8K/011xAsIe/0JT5+kQh9S9g1olkm5z
HDO7nMY2z1FELY5ZA8wvzcCqM7IVBbvBZKcIehVAwHu+1e3wcMa0corchL9v
NBL7n576Fewii6bJ9CVtJnL2MS22qfD2fY3CF5fuABsvUj8ESyaeY8mYNq2B
0woZJYtPN2AmzfOJ212yA/ZcBnHuOy0ZvxVxivCMIdM7slBb+8qMLRftIVBf
okSMe9ryf38JeQqIk5J/JOF3r/C4HzXAncIoOFGjPdcBte1f3K7gvvNR+Nj5
vIahOySGXO+mvhp20QxcXWYhIdY2LtDoE5pRxDn6PU47XzQfJq2j5BQ8arzg
dNFzlzuA7Xta7NQ6rC+uqKPPIuOq+d5k2TQEeBjZf3zIaRUrxEuXDi+puFRl
TDTmYdmNy7Sbe9uGuYRY7yOU0cAi1iATVu8i0Xw671XXId+7igMw0HibVtn1
E+wTTMC1xQheZSZhD8Lx/WoJynK7zOV/xGRYIpyZbdnFiRqXP1fJG7caWr4n
LASe1GkUJ0cIRhQpZANkkQF3bzpu5nk1ifByS7unNzoLiRHaMyOg0jaPEoMJ
QbkDzSn8MmK52Q9CCoc45Ic1CgwZbAakJsYovez7+1oh9sxUaBAaquVQ2J63
iaGOO4T88vzdJCXZLLAdB88tfDxXzh7/kaV+caManM6tFiYbLL+XtDlm+BkB
1bqsqWzEPu1dgmGjLpkDuzrJQrj89VQfP4X3MjJh4BmGl8OexI/olVGBy7PC
DsPphTw8SP47/K0ZdACIyCr6BzfmEBrh24zqUhTvR1tuHP1R9qZ8zd7iwOuT
X6H+Uzx0pVU8U3ypGQBXK09butoOpDJ4LHpU6ZT1PQ1s4v5/EmJChLJ5dIRJ
NzNEs2ZXStzW/Y9hX1rDKqWd9mhVTDoyv3BGLapMCp/9o+M/I8Ggk74/BHdf
hqYjhgMGKQWRfkWZ2TioUYy4DV2D2veYPOGgfIk4EHMSg+dJbw9rs1tKXTqX
z/BInVkKm+WSSaFY6UP/bifHzEC48bs38Pzjb9A0jWhPNh3ZacCOwoRM+7xf
1G0TGUWLz/NjBa86UDVEcUc0sLzof5ZvYSmHwY2aCeGFb46KSuINzjiQUQzn
WnXNcQ2H9GaB3W4q1JBTuo89YojlSVSYYkqufCdMMYtG6zgBYZuwqitqJ79o
4T9dFQA/axEH/mFVF6Fjb/qXkV17c7L1etEkMbjag7ZOkCGNsW6X0AnbM6oP
RL9NYySP8ahB/iv6gPpjhk4juE4UzPJYPRfoCbb+Ee4t7wjlmLFeABI4m27S
EFE2+5ZFkCnlgXLfQK7CfjZVUAxeAAOMjwtiLqqIUYvrgRsKpgbUGijZhtUU
DNXurutN0qGd9jPA6+J+s7795M7NGTnkrjm1N0Y6p2ItB2+oPm3X7RP+lQ4X
mln8GlvQl2TPthhkQfBK8MrCz2WgbrEVe1yRBfd3qpCXCzepzWi1LLQ4BWMc
42LoJ6NoF6okBt53k+5PxpnS/gCsJsWV4Dai69ztr787r2FIKrWzvcW2+ZLU
1Spkda+dPSNm+awSxPzzjL0nwtqD2Mb2IRX7/ZZp13C6YyOZ54enXCdImYwz
ky2YG2D+BO5Er0Wnm4uLCvTz80PiTSp0iJ5uAgGgqv5sPXQT2Y3Y6r6uDmNr
+9XbIZHvcBq3eXOfpHRDMxtB1Q8r0ZqATh3WjuMKS3SjjOd+wXoMGkBcDfUB
ueHeuR0dAbt5Hza1QM8c3mQg/KW9KNk+0hCCYFCpZ8yAcMR8qulB9jEVrU1C
wtnc5Ghaw0IFiFyGNDo3S3HQUQ4F77mrmkwhf26e6jlDf49vZwJr5B0ZVBWs
u0MUM5Q+sGH4YhXe80CGzzQl5OP0Ee4HkHFfG5Z69qpHgZ4pPUlIxh1KJP7k
baKR0LqxI8mbArvcNmsV5I9PReH+Fj0lyrBfxYRwY32tZBm1QvuTV204QgA0
/PrCa+ICo3FjZ7ePsiSbVteAzdILLbKoLDLZlI0776qETQrVUE5cPOCT23Fq
e9xMEAYJGrtE3z6jOXcbLpp+00OTCRCqOdGUT5osi8kDuXr93tI/GlwVkAbX
EgYt+3MDG6WuNrFv/rJfxJSwI+9hj9yVuf2zNiNrt+JPHtkAyvWg94NVBBfq
8NJX+NeSB/SdvQBXVhEbKQEMRYIIhrixoegHhXXXzWm0ZltHu/8CXgOCVhw5
h1T6ebcWvq6YLPFXneUAUYRmPR72JdwK1boZNfgW8khSHWEgFXfFRheHh6+8
dzMwelsKETLORooE5YMno7fLXCJv1ZJHJ59GWVcutZjPwS8f0sXTPqcsk/O1
DgbqS7iHsOZ2MQY6p17m7/oU7CjxN5pyVKbDoxb+RFjHyEXSplvJJTTAuhVg
a+8sMOzuOnP6F5o0n0VvJc96vF30NMSuL/TiHTSjflMx49TxyZkTzruwPtlq
CYNI1k7dHzG9ep2WwAHK7vu9/w+wOmNKVr9j1khhVYu+H/qNG6yx9OB6in7u
Vil4R5gbrJ757TbsGTzhKtw9o2OnuqASHVRVOgC/WqmWBrGcLo5LzpwWi/rj
vJimtMqOTs0w+bH/5ZDNpisWO/jcmhURK6UH94ovI/UlJYh+yj5l4u+3RU9V
eZ7oAGzOqsGAJRFg89t5jBtm6hvOmbhnSO44cKL/cS3lzGgx8O4VETfLqDw9
Ct5OZNzr7zwyLyUA+aa9LcWU8iZVG8G0gcAxJsfzU3mbPqxxZ5Coy7k1RhEH
h6sn+7bQg0QBfVQuUEQzqu2zrkE/q9RG19PXUtnEOif88rOVkHOowbXhGIoq
sCjzWAhDvo4MbWztIsFZlRoQj/es6FCKLhVgmdzyHVXuLohdwnw9KJw4d+1B
ADJ77N1WZlSCE6JdBebyNRWXGHZPTs3ZwNOyoFSZULlrGVxE9G23tZFpU3kn
ADGKxtNWS5EaYhKvQGs38wKz9OGD2ok8gkPdz0WtnjqEe7J91XXyNDpgR0lw
JuVKdCGq/Jsf5ShGtNZgiPfVX/eM3fGOgQ4PwiCdZ+XZ7J/AnCk/lxCIyale
RmdDEDFaAmibw9zXCJN7+3BFQX5GzZJsp4NA1SGdOyQLvamZ9UEt4geD5Bss
s+EQL+HW2QPCMJPbhDiWJyiDGgUaNBqA5E7x0XaPHO60Iwxf429nHrtEyKPn
ahS0tGd8B9Nr36SaJ8F7DnqPt6i1/TpCHJl4idCBylWVJTXaI0rLwCkwWHjb
3+b+GEdBII6GQLJX7jrf7tbzfqVvUsfEUvhk02DnAsjRwmL1C22NVXOzk0H1
g1JdoA0wWUueW5av5J9y+YlXkK9SJy0E73YKzffXMMvMENushL+/WwDxCy9L
LT75AIfqPY8jPgguBKzHrAy2zXN/4OgMDoMOU4U7oUP8z8hG/LDl9DSPM2VD
OzQCAKBZgQJI/ouo27o71yvgoOKRHLK2TXx3DKA1mCYgqtXqKIBJK3dWF4wF
cotCz+tDMSTP/sc/neceBxf/tlAfft7ohH1zMmB650YxFRWfMZJ7Sxaa9uUH
3yT3fxJagxtIrSqzspqeeUJPVNtFOagq3McaOEWhSkjdNJ/jKAB2vfmC3Au/
RGSbPALuHanXoI7eII8RDcYgst6kHxOFlAf3Sk4jfDq0Nzq/89DeYgGd7RZt
EDQ/qoNxf+0XF2oQtjhc0E48gQVrOwUFfjfKxW467LQLTjQ5gIbPNzEE0der
GAsqsU1R0kn8MVKH7Fckj3s/jVtY8/+qssTuU0EavImx/e4VF135Qa76X1aw
tAAgoLQALc1Zxg7I6QJJcQtsuK/172TYcfvcI9EiyiooSDXWB+oGDQ4bY6GA
lZwrmWtGomfza73yHyRKAILt6IG322f2MPQ3WZ9Nu+z/ePhbfFiFcFgmqnAP
tNO6VS2lI4fklzdDOUuWZl2IEptWkdyvMT/xS+l6Jl5jV08sfltfn0PIQHem
5Q4k4/PPee3geTZcihIMGuV+QwdR8eipeoT8qyOOM9zNBFdaCoJeCjHb36KN
41JHZ1xjYN3gL1pGf4PqLQmENILG1tZFR+PC6P2x0rHqeROd6wXMKzwL42J7
igZoZP4QnhVDeqziupeb/f9C+E34p/60IwOkCdr05caoVUboN5RQwMvQdl3S
t4+c6cLT+3MzyxfnykowPGFOSi0jU1UJ1sKj4ZcVBjuMFb57XPl2Z6/TGgWf
h4AZafXVfB4Y1htElEQvJ/vdX3XdBOrDN/R0kT49v6W1voeOJUMLQcR8sbLt
KC17l8uoRm6GuMu50DYu/pp2cc+3RlcsO6fsAlPdH9zR94badjCCRQj1MjQu
ymEGraDPGWs9YotAn1MrArVZRISUXR5Uqtb1+M04o+XeBkDdWhb0zY75Nvj2
uzPOi7cjQ+Yk2tY2aJ3/nC201pdilPKrtFidBZ16TMviYCnCgMpkUZOvQfXW
RRwHYX82x6cym+HnpvAFt4AWIjSyY5B6RGFRTUWhBKB7klSeWFvj34/hm0GN
FRI4nJrmsTOUZOKkCVbKFzIC3gw3rBSbU7UH/Kc0+ASlj1MMa/AQJAwRkPtG
/9JIG/tpYKVeh1NvNqX3z5sf2OCn07XGS822OoZGwTKX9mRJnZx26ry+wNIu
OwfXEzH9UXpIYhf++tijkYBAsyLhNQcrbUfpgCDcikUHCudqKAS27GsPZeAj
3uPTQIXZaTRp3hs1vJ7+eXowqOz2fE3hMmT7xH4qLf+WqA249esHxFbd3D5B
DnjXMOuzdB7OzeQ9YsSD/s340iqUnWuOY12OMEcSUoYHIz9aqWSwkNO0QfMe
R5HrG3wW1cmhJwfvWOwigIo2D8w3PN9/4BsK10Iu+QWWi9VbU4DWQh2che53
wDkQLbl0QMiz/TbmFrZKQPCg+DJu3omw5GMr7k55PU2NcupV9w/YCug2QqZz
F8ZpHIwS5pow0hJl2UJsPI14iIS7D5g7+Fcc5OTtInu7GFpXWLvIasqEivwK
ZA24cGG7Hk8NVJX64XCZ2ix1DGW+aZ5nX1Hkg9zxjL9Fe7Ajyi55uy5LkSDI
fEXsLshN9QvCBRlWOsGVFVLDPs2z1sUqE0PYgmYRlAwAEkhBR8c9RCluKe7+
SKbjaQ9TX6Ew1yJvc45HuaW5jl0Es8HbnOWxtgX7paZLkR3Of8eTrMo9wwzs
zkOXBkiqy/7xmqrU2E+t4rsm17vaDZk9UpFas51kG5ahs0Vdq9Ar7ev1J2Ig
xy7f16B0otObcfKlFTJ7ptsF11AldIuOPO1XJ5eu+C5aApwQr+aQHc2DJ8bd
oO7bRdL5h/xDEBzEtfjOyQa0M3dRrf1yUC1qfbw9A+jocQakZVDYraWULJoC
cx8+s6oLZfcMosEHOcnnrvZOgFmVrSYOfwRbNJUL6+6961qjX8c9c5vMIyj+
BxQLh+D2EgSR1aCULmzTSfzTkCsCrS2f7XzNMcgsNx3KMDbcTunibFEKJL/K
UB72FwD+G4GQx/kMBeqVZW1CYTqGcoPDV0UfcfAAaXNPxOMJcYyihIDSQ8fJ
f2w0fkwLdad9sQiQEscNdmBDG9fkZH6u7S4qbxijV+s4ZeWTz8qenFgC3RXb
cyZIdaQdGWZ49NKwmUJyjVX9I/ZJJFLf5FGBt6DT/VA5NuqDl0LOXQVs7bu8
f/zm4s8Y3KwZqogk2GqMkccCovhLRKvzSdhxuEKmKXi9pm8KgBlNiCvUhgTc
XQXStng4Cjfdyf4qJMnBvaMWn+jAmy3As3Ro8XTSV4z6xqICXvAJHUgSLwbS
8oUHIQJzW0HsHqTj4jXsVfshCKcLe96E3XwknxuldzWtgOqRnGh/brsmK5lT
Ts6oBJSGdCH8V/DmCJhl7vT+jF79sUZvobdZY8JdxhT+v3UZSHtFLA2zG8Wn
9qax5WswmtnX/CxnPv33C9KzyRYDcNBP0zowdzx3XCbyrz6YevPt3L9XElil
a1A4uCGmEZBz/lEYTdLz4p13qfvksdB9SY9lgDfbireWyST5hD0IdW0Wp2F8
vU4Xl1lyTdqZOY3WcOV9JDtMSJWY4r9eNTU7v71anukfxc92OhxL3Ndgv1YK
cUsz9hv1w2/kSTV6nyLRQKW/TwEXTgj1/CbjVFaWAhxZ/lL7TdsIJyPZeVSy
h9DH9JogpC3BMZBf3NjpiA7oKpJQ5abzz2H0UsLSBIWCjCEhbX0bq2KV7dCQ
XDyPdNzKLy+R54BcUMa5ogdbrDJ/pYcYEt/2WBzmqJzAnUBxTL4I0ozrG2AA
za1T6iqMulMDC1t1YCrHy577E5O0UOxPOytHp/PC5pCI0q5ygivSENhDRq5D
2a2LgGsB9fB2JicH5mzBv9aoICd1abvBHzo11to6LdXNHtenNUSzuS4laOyI
GGDSmyQQFw/+NofGb0QocMmPvYha4NQi8RAhaCpGeadMJ/qWX4Iqz9nMQZ3l
UAMDPtq6oP+a1pWnrzVffKoneHqJWbFioWWl61bW3bj4limWYtM+QJsVACog
DVIP5H30JHdbLtaw6r1Iag1ywGyrzcUoxYjeCBbc0rr6PLQkKisyYs0Bjd01
ybUaf/TO4Kadi/mkU6k22vN38VlelBFErkwrJRf0Yl8HKIwiv/eykyT7k8Ym
hCmeB7n1eCcZO+GASd/4oSarFd5+T8mzrJELnhrBqGYGXrq4lY1EMhXtynId
yNLhvWaU6xF619afVGul0KmpIstmoz4t0K6ijfAiqiOD5xSzzANy16av5nbg
eKPG8QYUOPXwALNvgmimIMRvUuIKQphtBbzjnb/R8EUz4ZapbVa23b1sGrA4
3CwfKn5DCz6OxBKpYV2UwTh8VpgRo/XhCv/NjZycTEQ9deIMcJunVGkjU0Ii
JBccZ87+xmY9gEmYAIsL5SKJpCK80+m4kynJSXT4qoMtbudAf96R9MA0YI3E
7eaRWs/FkVGYglybLWygxeLhywssR1rrzNSsMK9xTJ6Floz45dUAKvpq6HOm
uN8JChElc4kXfD4jt+q2XlcLoR1S+zoeQxH0WK/zs//Cnk8Am/xv2osP+Q3C
oaD5BJLGJBJwZcA3dU2a0fAxJpJy1aC+7mUBH+P6EDNGejajx00NALJKFmPB
M7/Dlo8woYcpXVKPRUxbs1BQBQjJDSuYtwLNBEpNPDRUcbF89BNhJrTbj4da
ijX4Gc/jaN00Wc9m/IlbOLa9z5Cf1QKiOYKZ//0rNSmRP++jmZ+i+eO9/qsJ
vTCgJKivo3NfXitg5uW2XwSV6nuksy22LIQvMqKgNXljE2Vmulfm//lFwXcw
gvkuk1krfGhisP5/kP2qIOlqVp5BomkmjyWPM50ZYqIdoMeCg13XZi18gzIT
oA2r/xhTEwu/pEWtsQ7zADYMC0TxG+GBS5Q4wV8NjLEB122z2TX8n/jp8Mxs
rnTuFxNO5PaOhZcD+qWwtQ97rpkg+Hv8MSzmomkqDqz8JqafCyMZffvyJIhc
FE1/RJ392/lfq4B65Wjhk+l9PHFIDLCvKpw8D0ZQT8kMcqbEn98wBeFmwyQT
UlhDcLDTM/q9slEXcwEx3aqQZnN2KdSBYeV5IKUOTR+YF75a/2NwThL3E3XP
aE2kJ8fnDeYy2AQqps6ty4ZbRMTTqwH6Pr9vVFILnn1xSLm9cCaAykm52SlH
PoWeI7og8mWAOI4hMY9YHoobfUJkLxhz8KLdIijC/ZrRJB4XMX0yHYdDtRVX
fw8ZoEBCyaN4hXxthLeX/AZruh0G8GYh6J6R7p9MQcEW0eE2HAv0OHNH+Y1K
2I0pBHmjBTRq8MZPCvLviBkAIdBumXkY9tVbHCtVoHHDcqjHv2ulwq7cMzDw
p++37WnGCrG4okXalqNEp1pJzMtJICZjslN1suwwT2rppBwpYR3iskOLxON7
dPoCZSi/NyRfHpccl3hfcM2j/OncnvIb/R0WUGU7l2E7AwZoKM94A1zjWdMj
LO0RzmXVim6OP8LxcgZrCQ4pqNNm3Lm7vFgJdtr+k2/2t0KkF0fNq299RyaY
SHJOK3Q4oKLQTHt5KFZOiB7sC+vc8wbkXaJIGfKWtMd762r+RfQPq4w8OB/8
OvyDuWFPfgBttfX7g1wj/GpADlJiwPSYnbvcFEiw+601sEgUAl8je2PIpqYf
N8zCI0KKJq9HSM4IrYgFtaLiuqusZ0l6pjDvgRCe320Ml6cuarGIMgdGJzaU
eiToUbnPlFAbYmFvUCZ4kKw0jg8cwOYsSpNdNzIfmcaYmnnr3R+xoYjrHOok
jddOVgNSlUxzh6/c8AGZwy3TN9YSDPCWBU3x2nXoDY89Iy2p02P80vK6iRA9
3EqUmFuT/v/wOELWwnvy4q+J5jZ0fKXB8gsEYOrXa1PH/P+Olf4Fy8w9VmcK
gtYMK/EAt9Qc4keBSn8/FiBrDXT34jVjjntjGowwfZGJkWSnoV7CBZv5DLKo
6zMrLM448eLXB7OlbB8rmHWpIvTLsgyr5PntAxQld60rxsO0Rk9Qvg+dlw/M
ZgLSfri2OTBsiwUo0ksZfHlNdmi8NcDz2urQdvtzCug7SLjBHkRk+haLj61s
71XqMm61MNYF7ichmbwX2yDb3V49Ln8lmfzHU/KgkmwfA6f2/xW7lsdSJUs5
r3ebA3jne6cwxJPEFclQGD3QoUD/3lI8qJvBCipS2VJ/MuTEJWAaiYvcov9n
JJssKqc/E8xG8v7JbiBF9FXDCK5h3xCc1NF8M4V35mlJKY52I1l1kpLWoB6L
6QkWxoViy31kXvV7oDl8qbZOtaJwdcimVKnEfpeIDbmPJzWURCdqWcWehc0Q
vvoCjyJBtfJyhdeGxH8ISUueY8UuFyxUqmVvNYHLUqigDg5Z1qMbKMqmNPC+
uBBcl0qAgI/VZCUiq4M/XmPd1INk62McWHSt0Z680v5jIJKmpVKkMx3Blr4G
+feTGCrzYMh1iApDGaMK8xa/7A16V4uQZxCkurjOj/JiJ4TiuFg29z0i/fGA
2A1hmjRsFRlRSG1FICEup21PqsrAjCoKhoLjDv96Gqhxft/YcE3Ib32In6V7
bI/3OFk3uLI+ZQMLA197yJ4c6gTNJ8OkomJQRU5QA3I7Pia6crfpJryXg6fs
Rmn44FVSAW+t2ERF8FWa+3uGv3xRfESNpEFwS710NKT8belRXmjNKiAPWrLK
zjJlCwKFlb86ryFbqJBnlmjlQegSYTdN9YiH0zroXGZxFnXC68H1jqdwxjYi
XccyN58sG2Bts56FGYorYG5H/VcKohXXpMg0GhjvA+H1+gNxNfw//5fkwR21
cfNAi5eGBiP+HyFqb6IgRr6+Na+3FD//n8mps8flY8NMzSkMVCfUrHp0gVle
OD5LBFNKgvwsbZNEP72qDUQuHVSbOSObqfo7/QUSJvTojNvQ4FVPjmFcqVMp
ZOFEHYCrze+fT4PBEPtmFO073126tsUl61f4hndFTUsJkPyYvG99wh7A6gF8
Fw758KXs00MRl0MLEvvmDVIXXhxlmQxZXWvYmllklmbCY5PYkeVXtMaekzPj
RHcObdGmhtpEVAGhx9DSJfeL6j+RzaPqj18qUuwtMtkOc/tOoabHJB/1CJ2l
hCVHBCSKsInicTFEwPDVzUnrRo61Mtktxzl7uPnt1gpMhgbVEaj5+FpZ3gJm
Ycgmu1FRsXkdzWkTIyxNxWgY/4E5fXwlW9Y4jD/Kni2pouADWGI8ghERrjKK
qXqk2jJZf4mGzGYevwUtfW2ofanRj0yglfb2B6Uv3IcMMaLc/jS3Px2AKgIA
4iavLRbtovoFnxq9XQuIKkAQEvDY68QeCUty9j/AqLrSjB4WDJ9yvSdf8AOx
ts1wFqupDFE9JHEASC4LQvdNRZ7geJbewBdExKIf8wTPVEhFiWVVCqUs8I1y
0/Rn7wqmHBkGfiu3cFH34wGfhekoS+/WRN3eOa6BKb54IRZRAKQU1/s0lXhL
y9nVeDZyXeDYd+pf/sGodjyBli8q2hSHPMiJ4z6ySMqc9zAO8sDRsu7Bo39d
l6F09TnSASrLL4X+xE52YmhZoWXnDtYsJeVzXwREC3J3qv400becByWa3Eto
M9C8UViK/q4755TfxCeYQuGClP1Bp6VkzdgDwze2QS9QMlvTl2Ra8v3wZQq1
Yeqt/hVDYA/vVzEuomCg/24em8kOuVkwyNCXNVJJAxk/cMUGkzht38jCpIWB
cUfzELgQuInxywyQxuJbipRsd5fQeX+NfZdZIDEZlwe4VI5ydj9dYexQvFGl
iD/wZJAUO+SkEgyLJinBKWrVQluH27G++yUGQgvht2x9J7iVZaNZ3XCslGyE
vuAG18fWK8q6sWmSv6Xos3mTs+vkRChQU5Jkw2uifxWLTuC4StxGMXTyH4em
TQ8GGQNrbbssuwfhLO/3Bp7B+paQyVlKXDtAaQEqjW/l3paI2pUrlgUqs5PF
TfSa40YnaBVxT1HT3iOdL2MRFaEHTz7nwYlSTeqRXy+NQ64JrjbyyNFOWLBM
46roki56AwQf8rIJ935hyw4rDXxtnB1CehhvcePY9voQFuBs55juABWiSLRo
oDE9yzbWf3gBZi+vzHjY2Hc1WfFc8BvT9ZeZgXE5jCBDX7P2LG1KQ3GAGLM3
QpPdLhaCgbA9qCguLOKfEt+f0dPz4UqnFWn32CnY/RgtPTtC7y7JVDDEelWV
ai/kwgIA0Wb/4GhQLX6xKL6R7Gf32NzVpAYLZqCBkp7mVz+K+kRTDg32oqIb
/nrrMfdpurSpmvhqoqZKmTUDq8sjHw9+tVCpXna+8yMnZIcG/AisGVb047vt
aKSPeS79DpFs4yzISu5bh/z3E9Eho4D8ZeBYcssV4Aw36xKNpeKv92Jz5Bh7
tQ3qffdelrCBJMzLxmWHjg50SI9rCNTvXUuAQIhfjyQt/T7a8Qp8L72x0qZV
xUGjVCFJuwu3Jxg/fw2X2vUuxw2PVe7gjxxRsCVqeqv6l9r5cODUlGxxbV4x
s1ol9A2n8NnU+obXRphGUvw+dbOCUGMOC0RFHa5WumPEILAM6b552XPqnG5l
ouVPasie69BG62xFHAfJaihS0Iu7r2XmnHc05ET5PjZ+SqmQ9cPkIfsw8GMW
HDbKgDdrPeE5zuvKhxUgz8g04SYyWqzk/skiISqpxgAuv3SoiCuwBslJt7YK
BIuHh8YsjlkperQ2LH5HuP/wUARsTd4ueRjduzZViaqeO1f+Dk5Fqw4UwREQ
mi1yownPeuFGdFh+tWc9i2Ntl0/MYbO6GYBPqt5jrFm0vnVvNGVIVI1hwNwq
RbqgM9hcaNSADETQmbmis4CUfAS2vM1rngpzx+cNqwt2A/Lh274XuBMfdj/b
ZotMWjquDDMeyLC1lp9RiNkqlp6W8JIVyDSvMoAMpNMsc7oe71MFqRzt8BVn
NOp1+oYO+CdNoSDCoUI0ttn59A9E5zQRv0JTuFjkBLUPywpGrZX+uu4+BTaW
qSnSLakikxL0KwibFz0c1rCgvpnYO//BZuR8yrAe87sn1M9aqQOpYlxLlUWi
KOOrZccIzpuXHxw3nyTt6Break/AypjcT2Oo1ZyJumNUxy8OsMOJDL1nxde2
A/KV5lD76ow/LrXqtXy/OKV9LvglCCttcI/naRg79CxYKYMN4d9E/RdKtHOa
/nZ2YSxcoI8sK/F9tpXFKjK6bBfkpjDbooo+YFzmKQzFiBpbyYniNNxpQSxZ
XR94XXkZFP4C+wulkecF5htWsC5ltoHn3JzqgQxvBPUmbeDOoIy5HMK6ZTC8
JXnigKLgztT9YM7JREcXr0uzg0gRofKVtMcZjpFzut7mL8FTLOVmjD0IfHtg
kyOFDsizqDxioTGcXIPkLPz3umUv6Hvtukkw5BLPK8+l9Bwg+1lX7X2zGADW
eiAnhGsPSb5Gd4pqJqMtJkUZO/MqGTs7XZVnKIWfAB52+IUkf8fzBQfNGoyL
EbFmFRsv7VbFiQ3wVsbvKN5jw3Nob6TfSd+1BbueeVI17hcl63/tBj87cGlf
X825GokwOi8/DxPOvgzvgsGmNmQZH3jUr7e3wpIH1mtncN/gpNxOgi5hJXwP
efAOOi3A5yMipxHoC+cZSkORphjsP611nYCy4K/EtCJwl0OmZdv5p4KdgSws
WhvNpBrw2R1CdrLJLVUsf9N0evJYt8zt2G3gvx/2nZCcnagUPmMp/cztbkrR
dkmkGrLTR12vEHLQ29s8i+kRMXpDHtcgoXIwhtgjm4aK7dwgzQQTVSG7taoO
Rb5/NQI2DxRnBx6ew/eNGn2TF4t2dbBdkzFIAkPwDU5ImJiw1FcmSSFCB62y
dy5yIxf0733CqS9nWHt26PFZXXZDb9U9ield5zjYlr5P6BHS2g1sC1EC8hvB
9nBilev4NstELOvho2WAmcIXFvmgBGNB3XLKYEcW2y5GQjRtZurwHTPG4CuY
6fxe9UfcKHjxYe3buEWW+qIDk22bf3fQdB6SZvQkucLpwUufqGm2krGeZwWE
GWzBwc3MTYI4eQ8zic5iCM86hHmYdXK2hnK8Lr8hrwl8odrgLeoinVjcjIAR
BYPb2soEDA1iOCJZ9pYuko2RhvtGnGL+DK9RVHWU0426r4EThS6TaIUSZRFn
tPvO3jAxiGOPqk6yW2ntFuu24rUtXYEgn1ZMaJgOWfUSQCGbZtHccf9YNEx8
HdNqwAKUjiJBEo2927HyQWODJcsrGWRZX4sQcAWc2aOKs9NtnhJ7sfQXraAj
oLz1Z+TEQ3L0985FUR+YQ2BebwI4t5eMEWYvZr2UVPH1ouMxNjAMNzatKMlY
/4JrpiCl6VPns+WVB0fBcYlkOXjHGRwYshBlPeQEvSGl+azJWT7sLQ6wxTeW
qAJPoQBorRYOyZI5dngMzmbMmp81hGtJsVpr8B3S3vdYyrO2X7pJJgzcypy4
EmThXenn/7sieIAZZl96TdvHcnSU8b+4/CRKoRGykAq2Z+PEoXA++wpSenKp
QJwA/33FZIOgXsbqA/FtETLie5MZwTpj4IOE1xeDttaSSZ5AYPPkR6LsOaAl
kq+Rm74w3pS1xXOqXl6LBQeViRyojPjiJiBEwG/DjuMZxKQ/KPVZnbmVKJ0V
jd0MLmqxlau2A77hVjoEFiPWLoWgc3yJMEPUFeF8147VK/lmqBoV0BG2O4dT
rP3s7p8JbuGw/H9efl9FPYFvviUw53bJCOgWObKJUm0CCxi8+tPD0OMZxTGo
XZmp1xMyLlgnbLXzqPZSAU/DawoGleSlF292Q7XpMdEPYcbB6MPg1/K4cMMk
XP9yMdsz1rMJgWme2YFow61Z361vCmNgNTHeq7XS8TV+HQ7tj7+llZ/SlmUA
mPtg4KEXtFkKxNI5FDhGlsALoMUcZz0dD7Is1PisnGcCwUuuwVNH1CKJFBCk
fs6/eGii+JeOja0HvedyYVwyrx0Svt7nx9Ld/JqgTWWf0PlF7kelANY3nIts
fF2RvifxvMpD/4GdHfQgB86rfazdyMVJZgvJUTsDrdQeTqfX7BO9Gku3XM4p
cMXu7eYm85orF2iYZZh5Rq9GiqXemuHaGF3qbdrJqS0XDVfMrqya0oGorlgO
wiN/1gJF4Gh2Y8zKPU1bqnDPB9Huh3axNho3xFQCTXh1AtpoxN/6tGZ7pXfr
BzO6QYLCRaVOCGkjVQbe88aYwcB6RpFo8DPcwsJOzFk21vOaRpM5c4REYQgq
MWpRuPSYw4XukwqscWQGmd1z1YWKWm2cWSEfIOsfPNkVsXThKBSnDanQTYrI
U/uiUupT9xsLAna0pBzysilsJAMnWQ4seJF/fkZ4vpiNZ89LquqR+CV3KRt9
esGjNcCLp8EN0Qug0LdK9dYUZ/z8hukRDOWfnlIWhSIU/QhflHDC5xWtba8c
uPoU2ZdHVUwzLPGNTfwmZU3lg6jpPvpIA8pnOhAs6vIBY7OAsGMkBpnFYCMZ
ToWoO7A9CLGuodgBVlhBY5aRhT924JJavqVECOKEsKlwDEO+0nnwMNQqWyIC
tHlE2m7o9yNfsniduyxOvgnqEfLQy4/ghP1KgZqdgYCoQ7lSpY3HS098078Q
fCVU9jEdBhs9yWAYqNgQfUcLb13gq2RBXC4chz8xyVN1HrYq/7ZjqBKrS1sO
ntb324lusDyZcgs41qpCQ7hZ+IW+jT2O32ZbJGwSEUN6g9Hb13ttBYCmmBDa
6aNfMPq83KJvPcyf2oa+LvXk1u2+25lnO4AX4P8GM+CLQ+BYYuGDY78NpAth
p04Ikodaq2N5TT1rKafakeKA2y+P+Dz3BGlK22y0qvRgVIe1vS1qzqOr/sfj
K89B42ML6UEXnGEM+fqb/3DTqk4VwMKV9Iwciy2OhrbiyXCKtLvJjI2k1vtW
X/2zxMI1A9A/IEEL5Y9CAA/HmMcDMV2GQ7BTknGzvJbaj8bzgD/JtA+tyxyn
eZgabH+ygzfIjUUdeO+1O4tnIcxSXeDBq5MXNWOxWX9b3z6VAo+5KvZcQ+DL
ok4fmtI7EqSZqRnslfmV68fXbqhk+Ia7wRPQypGKpfYAIPXyuiiKx1rDgL48
YfMfahRefDUkdrQzRn3weu12Xx2zRMI3tZRcqqO837i+Lr8hZKm0xASrjY3X
AeovLWeMjK1JDy2ofXUGnowMBkC73T9vnUzPzOdB6xfQIKgIXcTvfpy5dzgp
SBfTIKp1O5rlBzJtmHcOaMxBv2lhY2UsABfM0Z0L+/7inn5tZ08iOZQ2vRCK
hKgVCeA/Rs+a4RXGlrYw7bJCD20YBuv3Etkt5TukKkJ00ih1+EUTQIO0lcvd
bbsqemzWOPJhvmeIPK8k3w+l4jucJFQjqbBsGdoyUnCHezWKwsX/QySuZZvV
CcY7IqMfJ2rKkYUb5uyBGOvjjrgyf36GFXxEkj+Uws+1RPr0vDE8zIL/z48R
Bq/S61LIGIjq4nzmpUq50NauPHlLpc1//yLMUt5IG4kjWe/Keo1avfXA2+yW
jgd7+040PBdugtFVzBV7Qx5y/iQTIy77psk+Vjn2bJN2Ryjpb/vt5gRktk/Z
f9SM0cgQlLy1HGhzyaac0xV/jmXZcRAsngaB5VX8h63TLKv5nPQRmw1ccoCc
7PGX9WDmDBW4hw/GOfr32Pqo6q8vpnaHwp/A1zcoOPNIanaHPdsnDx9NbfZx
2W34gjILkOocDUVSRxLSgDxTJRx2uUypx5Rwz3rTJVI/0tsdca6t9a9pWi/t
J7Bk/NQaOeHqmmMg54in4BxdnDZNiNcch1CdHbRnPK7xyF6vTqiKpzhlV0ZH
RTHpKKVSjPM6rFdJpld7bupBu4r1LMFmNLUcUgwC5YQLEB0E1hw1oIdJi8RZ
xVjVRbI458Pdshfa4kCkeSVKKRbP3itUe2veq7yMZ5oJNWAHGj3gYH49xnZi
dWTncCLa7LzdYEQNSfkCOc/muUCnFNdbWIoY80NKKbLiVIBif5MmHWzvox3S
7/5vJ4n0a7M6/nm9tNUHDt8L6hJ3YhcqB4E1eS3ypq+AignaqxGISK+bc7Ho
EdQzgRE/raBQ36rymnuCL0JA5l5T8fMOpAPxTkvWvybktDlMM37yeyDssgCA
l0rI2UGNIoID0qojbI+Y42cxUt3xE8zZ89LkUDbd+uduwqH9UXGsF5Y9xqbj
ncIDYoGbKRLAVGQpGXahigbnM+Bz7tc2s5+r2GA2Srwg66xWre9uvZj1MB4V
x+83tKQLwOiVLqqAcIQlzviZc/1GGr95G9urgVGw0K9d7lrgaDMphYItUD/n
HAu1/n4m9Hbfc5IxCPP3JoYJQz1wZcKCxb96PW+CEfWzYGMJPy2DaPftS8X5
Nwk9WZMFWF+zOaeEssL8K7b3NBTLF0NFSduX0pc4w+kZott8NdvC2NoPQAlj
ltzsekNiT4LFo2F515b5f8xfDMz97nk4gAERqrLIuh7fquHrjPcEyGB7b5Oj
vBAU8H/l1NWkc+DB9ejOyOMYwLf/KJGDX0NvMAO3lw7gkafBDInIsAyNOHPQ
aPmyEBF7oPNG+eJpCIJzUiQG3D17tcOCJagjmULgFvw96SztXBhsn45m+gZd
8MYUFF5V4B2ObNPMdvTTHWwFKhkve+5wGNupGR/Y74U7+BFTNBWxoBIIcno0
Zn55takvxliYAoEb19Wi4VXWNuKKWEHBzgonLz9QGzDG7HApgn6DZ8FI/G9X
q69fqx4LMn/JJ9xvMQhrzfV/bnIvdMFgmMC/03YNbwS2soCaliMnTF3mKCjU
O5V3rJWqfB4OnSsQzOi3d1Kokzr7pR1abUNDpB8WzWKKmfbtVmQJgRZQa+Hw
SJGXlUvnTpCkjhl06Dm/04TcyqlyLnp0sZDvldah15m3j0dZNju9bwbNmqUr
Mkgn5jnzZh60BshXk3IGy9tN+nL/7582D/kHFKGqvcsjzUl/JmC6DGZCF7Oe
AwkIhctUAXKjC8YJnoVeUPFI8FCWs6edl3gsZWKd5/o8ujKtrH6Vqp5imhmb
PnjYFk4Wx/gneA9pApNlU18I/8r4MhLwAMyrKvPzsk1T3IDD72D/DlF8Efh0
wCiT2elbbQFq0okcn1guhXgG26z9EoH45eFa9SX8Nsp2f7kDbUIZfxFH4nml
/sJ+98+MOpRj7WtYxAr6BtOpG9n1ej/YTt8o8SClVyVi9FRMlChgc0HXpOOV
7CHg+EvH0pl5lyLJou5OKy7n9cogWu278vMTsGleBfAIa6qlHhqSZEi/YYoe
oKBu/993czCW8IuxrTCIhzEbU5CWS9O6NoQ1UKa3CQw+Og+cyjgEaUzma2ZF
3bOs3Oe+SVWg2digJxaKWMikk1OIRhbnDySCXVWh2IN0+SPROPS5zcIqxsOM
SLweV+MBOUXItDhz/Scni3dvOm4T5HWC2ea1awZE8YkzWDmnze/i91B3Ucow
oKNgOtIHo3usqJ52lcTx7ns+xcKYeq+W/D49aSRm+Pl/dHEeVuIaE0yPgwMg
/mM8Bc0KiQZ7AmMI4sI/9JBzuAHKf8GC3ZT1U/HobAoT8OQRwd+uGKo7OcBB
2oYYIVlCUlbSWaH5+h0seF2qpE2PB+BMeKQ5Bw4Kk6jNWvsDDeRH+OFmtPrZ
mUzYogXiDlF5O0i/K9OUaqP177pSyETUBCxQXB10EXrwsIqAXYSHjRME+phD
hvf4R8zEAM44SBpLtg/pQrg/hEdYhoBuKkfVdrwjEOe6BgnBWI2VSvMy65nW
Z1flFRwEdWhRJKzJpTFBFLmd9izivaEiFoOVs+mxJS8p77JZegHNxqjWp6AN
lVi6soUB0p5WSW2BDS4qDJ8cZwhx27QBodDmsYcyDIYAUqPUqgOATJqff61N
9sO9cn7ZL/YyJBa/slH+v6OLI3ToAKBrquYz9ysOh+/32lCTNU3Fb2E8tosZ
wQ+VgjNA8ydxzs1XG0/aHU8b8htFMi+s4/5iWhxnj/YhJjZsuLQ15G5wWH/s
AymDNzo6v/lP1Kigar8/AbG+mWAaTk/Cu2hrL8kBK49vqMGx5EsjvgkCjBEh
sco9OSEs9frA8c0qkhrvu5ecyGB3wop7sr/0LfTYmY6TCgSsdvP3fgC6Gwf+
bY1XuDnF3vsBcjnC/JmKhHoinwaJVVFyAmM4ZjwUBWRk+9r3KmP1RLdQxX4i
k3esYJJ0tErHMk9toHt7y7VnWxFtQ9Iufu+jOiCLKVKUrtM6QaiXcqgQtc3v
vKYUd4JUaFQNsb0GqKT05amBOMcHOUQNy6HtiXb08tYlmHlchxa6+a4zxl90
hCHKiHAivyznuLoTOxTmYSrbfFet8qYSUqwvl1E/lqhajt5XIHB5jLnMHNta
1md8oDGdOzmFXXQUiIdto+yvpkemKYRHpQFR2CPeujRLZcZfDdN4Uk70Q3Gl
1HFK07chS1+WGoRwZxiz2AnFltcqzAp5q7TGYZFAaQfj8QuQx06I2mQFnsy1
BYSQI36y+U7TntvbWkuJcYNi43qjYRwf1eXAxEmlTL6bOMjgE/9xfUscKfcJ
loRprDylJC5YnMQ5+qL0hETj2ulkg0CCLodMUcM/JdDuq/fG/hRMDJwMDqr4
8XozD57rBwlXq9BgHyXOkyhc10cpJGvbAizFBscrK4D6uQghrjD8CKnvYKdV
6DtlUokWFhRlm2wr0MGpsRxnkBlrHdfPoEuqzGinU7xbIJGLp7QFVSU2TYBF
GYwfhHwTe1HrEZc9WB7D8sNe0LiLTUdnjxC6AhrzHngaYiS/EXklkfDvENYk
wioYA6H6I2k1vmWZ3u646Zdd29jzxQFvS6Qpjis7/fLet8udysaUSys+rfZb
wqkhZsejljThA8dHHTuqZ65UFrl146nOZeE3DMhhnOn86LCWq6WirL+SZZW/
KdRLdS1Bb95NZ8jnZhgtVd62nYsgFlR0ZYvWruQK94BZMD34LwFqNaTspiyw
DQh/vkoeMNqVCi0U1kAhQzzTiikdqB+ef5Pgn5NYZ/JYrLS+oB36y0M31shJ
X4/vAgx6fKaczZAUoXr9eqReznwToECYAg3Sc7TSXiitMrT32JUHb1qKTsut
z+MEL0INjfU3w0jM0/lhfzvAV6HS9NwXLoEHbZgtxUrEPFf6pCn60UuIIIXP
gDtRJYoweGnD0ROUl+YbUL2kO7uwJf/HRBzMurBp81Nd8M2x3XmF1kzkQumc
9IRnQCIG5KeeMh9CrGhjsjCUsC6SBGskOTKQuqRk/ykpQrLmzqT/oTMQXwAc
mxSUI7V41TsA5gaPWyH5xTH7FCkb7xb5Hl2OhDbSSQ1jYm+kbDqJKQROlDOC
WVPIyvpfjkZPIAZ+4r/s/5n1BrMrY/E6V4kmVgzTbYDwAQ73QcQAwCuWJhHg
Cu2l/dHUOIxoCcSNoL0IgGf7BMFylgLSpTSfLNFjJ3+hkMvjHF4NOuO9Si7a
ZNtUA94e6FKKF5OAoCrfjK+Diil+HmC6u4w09q5y2bqcHiKE0HBFLH8Oshfo
qe5sh0tSoqkXwlWg8y5UFzYfVvZFyZoMH53EK2Vak4O6jlTl/4PwB8DMqrja
aXFb0gq5/gQlWkNOgQnjnv0aqrqmkONkWQDwlWl5ippgMihwKL4uj597WJ80
v/N7IoEgaeyKqMkj3hq92bG3zT28w2Sl/LxBdDLxjtL9jjrk/BA0u4/TrONq
roLivrjGXju/HmT204C0LZmCs5btLZZXqTAArNeUDE+eJITSxCGuBy0yGkU+
nHeTBVPuN/WsPOsFJeZSV7Wcs2h+7qd0aI8F+i5X8lET2Dvn4OwueJVZYoNh
O++LWBL0CUszNI4aWU74beNNmVl/KfaPEiQZHT3SPM4C/84bdM563u5fZXPk
2RncYx2R+CUNtxJ37a8AYZD6KXumC5aImoUkuQUflXfHfRLOeu3krhpJTEIW
WicZ0JMfHW0BN1vi63JYw48CjjBUc+mjK2A8KKrV4iHi8OEcMJX2G0A9f+UO
5nTJUwxWQmyUrc1O7QCY1nsZM32HZRtje7XdJDPG+kJ1DbcFpM+efjG+cXMw
ciJTEpg91RNetDwt7puDut0jJ7hxXl3ls31+tZjCvEkZli+GiXuihsDEutxM
z9F0rK8kITRGe5PfUQ1P1vJ9pIxt8525FFSrOw6ttjh+452MV09QMIsTqeqf
SIweuPQDC4hEcGcw1VQj9+BTzJla2IV480ytTS6lvP1ByfIwNMth0NiYmm8k
u2n81Vii19IrnDQmuE/dNIQkdTRkjgqc07hGHLkbn//AjMAuLOclsH6GwnQ5
vNr1H2KQ7HVZHwsmIT1zGSPDxScu040PbI1lCBve6cz608Rg3qeTHrbYMB62
QehXlEROF/sPbqhqgLz7o8Qz8SdzJTacGx50MNJ2lfMfmYZ15eFEomBQAa3w
8/N6emKQwzTNd/7FAAzXFcHAxMQkBZyWa1VOPgFY78keElFzm4FW2jAX9pLr
npbl6TcBmil1cEBNHzQa3J5TV4fqzrZnv5vV6iRRP6m4uEwVPp2JNQNo5sIc
qk/nvPmYhoviG0uakNVpEU/oeTWP6Adb/mu3FaEAxdlUkU9XoL9GQ3xW/Jk+
KHltmvIn85BFxougezBp2ZrRYsxAilRXhNy7Wl6Fvk/M8DMf//ynhlhclYkw
hzjZRRKCKI6V5dShqZiprhc+i7QsIXFXi8/gCvOKNI4iR+J7p8JUYImLQDXu
7RDnggHmtVv8u9PN6n9OzJCJrt+UvJuNMjlJ0DZvLyID2s5LA8TRIM6Z35u+
jmZrCAO9NKOfHusUWf/esz5VhhPA2k4ELrEU5oy37iiyVs2VUPur5760ysED
5lqFKQpje0o7fhXA+yUHKYOLXM1VHo000gJLc4AbCZ8m6wekgJ9AeiMXxPbv
ISIe/hO9NMy/dohthbAsA7L4mAONmR5BcHMJ3DnLYvxyR0pnBEPuAzj+lvCW
u4xQ47axzx24llipxpelPSVpFdQnDykCLQpsrz/PaOFO7azqJy5jgO/4igDU
8PKdi0+ABJyB4ybi9Ue6jmkois/5oBZEeQ5W2AxA2KhZ2/m9pjrYdJ7XQxA8
OtyjHmfOi55YQ1k5EJJ+JToVYEMI/YoNzjv3LuCfJmdjkLiRmd3N12jU17jM
oEr1k5BVOmOeA1qS3LtEET+0KJm1qNEPk2IP7YArENl2fhPzdE6Y5rnjW/1o
k1G4l1XYue2/65H38uvexkALcgTtdbeqlcKI4vqFOGRq0yxyY8p/fCvzK1v3
R5KuZgBt48SgW9kUxKPFQHhdue7bMzTCWbnpuXv8gbv3sWdj0ch2RiRgXVTj
1LEV96x2F0i91O/hFA3JvJiCrb+VDYt47ruqxDrfDBn27y4QyoDXsE74wLsp
m17/IRf0CzTD/oIoQ743Lh0sIsGlfyPKFxIP+pS4eMX5drCznfvTwMZNfj9w
EaYU86B9upZIA9CsqSo/7lFRguqB28vffOSx3hnFxtRtKltM/OooITJb95e1
qtk76i9NupmEyB96zSwLfjwqnzy1UKBmrTd0gMSFjKcXa4SEpqo5grEA7KH5
DmA94Xvroppplp5YFwgSBco6VcHCBagIdqypo6nUB8bCm9BAI75+P5fppCQb
S52vGDEbK35xo6PkCWxc/y/dMjOeF+NVgV8PVPkGYF0VzkLXMp/L6Yg9MoLh
YBxMHpUsOVkYkxhlO2B7FSsueNqS2vFHajniGlsrCe0HflUGSoo8XF24pZGI
Y9BT5SyaqB7mlqYICmkqI22UzT4PmR1tRIZy0MephErL/AAeskADNt7j/J9x
mS50euOvkc42WC315TkYVvOhL+RSKuroFKlgCj+IopEFvHJZ/o0aLhEz0Vmx
eJKEmQfMPaZjYiM1HS0x8xUCgaegVSE8njaYR4gPD71oPThldf4QeDasxCUm
WzGQvs+b7fklPQMezEaF2UBdu1w8B5ukm2A+SstscVbMwTXd06G4Xasp2j10
+9u4jqzNcdVjTwhwuAsJrgpLZAKQhBC4zRpTZTLxLYw3QLLQDv1nzM2n9kTm
zE+4UjyPGHK0YWk01mzyEmUaqERT4DTjUirpBaMtzXro5oiYEOqyzIdDiLnN
VXcksQwwCXilwUMQcdStPwsnpPfwBkgzSJro3c1bOKhO5cCsWzFby4hbChgC
6+Meq5lfHXOt6Fn36OkDJm90YyWMkyjJ+RMz3FjLi9ZLiZSqkqorKRPhuCZ5
abDaYpaEf3/KrlkVLohrn7mFH/hT9IDG6xIsikvDn0Yn1ewDyVXlTj94SD3X
+3b5ZRGWsfDtQ4azmXKgAl132B2za4Tpv1o7Q6YxCWPTSEW9HPf9WmmUKN6x
BVZZJLcCwRMAJ5mGKHWQsw7/OnQpurnoHvLaeR1aQfaopFGcMPC78uaqivXY
LFfh5ulklSOZKzVONtD3BvTEsxAfHlJ+jDTPtgx77vj+v4UtjwSHjHl0AnX6
+VllgHOHj9hcVOR05jW0RyYsQy/Vq9ZzKC5HBAgvIa+AkSqNx+V57aJwGnNa
MQmlI2lySu77Tf3pm/cj4+/vmicI8SIZbkycNjOU5/uopuXO0bKzTsAqlCId
KfvdlL7lalk620JuVDR3QglU+L6SYBZdn4CXy1B3O5a0sOTt6t5DxORzmdIM
ZQXTiVA31T5GCDBlHPx1sVi4v29lFjfjuynaF9UBXdzt5XH9/Etf0xq0YZuN
51bxngZGFpk3TgVI+bkJjcSU3dOTNOrbpEMtkW+umH+IQo18y7hTzeCqcWhm
4KRMWIF/woPxVBVyCIyYARGYDWsdURqH1OOc72r5TtFluFICL0VNY6v0yI9V
w//OBZzArvWEHR5RCXntiRg4EMVQXM1A5f5zVEl8KoUmhhqaqwXr+vzNdTbe
ag8IjNvQivUrQAXDU6bDdJHKUx12TQI0DIv4Ba0oGkHZwqvru6ONGTWQEnqv
H9JfnyGsLyD0+t9QtLz/JiHZAcmkVGEoZBAgw5QyG8a7eRZPj40fRnz9boEb
wSDhTyixeaR8KcZ3WLwYPPLugsLPYH53wDvXT3ls3vaLJ8MqAhkZb05EfAgs
Uf/DvUuN8DQEEIzLh9f6gihN19WFiMBmOr0yqFuIYPJSdVGyVfVk8WgDHmTu
NHWLXLTVf/mMSPF2w6sdfB6hB0lJpD6XTcr78pk1aGAh+ZwzaRdX8K7yAp/D
5mzzc7To3OjmO8J3BKOetflqBYR2qBjapAjLFFg47oE28CDWGacNW5+237CU
rRj6Ouf0RVVRCE9d2z2T9rxaJAddfEjR6j4/QnF+JsyXev7ueTA2/PyXw6m+
fWrCSRzP/59/ICIlDR/KnbQRYAHC4Ezls8+Vj5JPiB3c5LsQ8KJxRd5VoQDq
thIHp1/9dnK8tl19t3rhFdcoBKxEAEKo9/ndMVgybnCQU58aUbb+3AGmKZjE
6JI+K0FrSy7tJ16BYYhjg1tTYIlC4gvVuKbEIG31ErWtksn/ONGXKxDemGfM
s1IFgf9LoarcdWm088RpXTk1CRjJ/cwFRj0eXa883S8rgkcpl05BJvQykUI/
2J6V1TFvxua52XjGn0quBwHAFPnJe5kRWpTOvkl4MyJJAA37a4RiELhDe8W4
GqfKFAciyic/Uef1entHFFyz2NLyUIO7gZVoD+wIr6bwYH8KkWLSghlytsGG
Ip1BWYfVwEDIGxnaZJjU1iKnej0IEJ9Dc9SFpGT/fEtb3Zjda69/UDLWaDpX
CKpLYMh5lSp75FuLBrOZ/YcL7ujrwzYn97eSqRdNpARyy2dzrDpIaRh2CLmQ
osBwHMHjE+HpRYEewxDGLAorgzF7b/tgMjNYNxBIkhyqeABBuvGXV4YW+vb0
XC0GDNsxzp6Oy+rBKdFWILM+byg91GSFX29/HeSRt+hsgLeV8pQFNF7cLC0I
7SaCwz6q0bTTdXCEz0r0xwmJ/4jNKM2IISB9D1bE/LLAjglVKmFi0hzSrc7f
kSuJvGv+P0Pr4VmEFWlltd/sxO70jYoQgvfesIIVctOMm3MWr5/TSUtbB9CX
g5czXEP9aBtLDGO9rgM+2EIl2p7CHb+CGG0OyhqVFyj4CZI82dtEIbe44bMQ
Lc1d3MB0BqhIcO1yRdBenFGpCRXxGTdU+ijDUCmB8eISdt3tVlvmCdAldcZA
f4eHjZSRnHt5WIi82y6d3Jun8bwyoyu/4B/uUNZMujcbvsiWyb56e89MbP3/
sceWRGh8a+PRoWCUi2MHEGCft9pnrBJ6/X7sxelOyENKYXjrdWktQ19pAJDR
SoJwvMFf1eHY/CkGImN5g4Qd52g3m50bXuNV0EFzrPDzDvqOOQGUIDGD7/Ib
710XWRxVlAajzvAA2PWxEmUP2kUAt7c66P1I97oTQ+DF1n8S9gOgILUZipZv
I0dYBrcwrR/ZoFlyOXJU+XUlRvYzKoRjsx/6dOzDjR1HR59d+MZBV0lWdopy
afr/Rro6uDBsvcjHw4+DkRUh7cE4BRjp3hmIvnUv6aVHlOfj8esAkpK5K8gQ
75F5VpjPUIec4MnW7vg9eg45WV4bE3MXlC6Pk5eUn/oibs54u1qHgqzOUHZM
p8NEyxUBuAkEB1EHPbQSH47n82MSRNfUzCNym1Rf9+NEUNtzt88WOByU+h+T
9IlmuLwukeSV5M71KXV7ZE//XZSkzDgtXjsCaSoX+XE9JgpbexexlucLP0cS
uoRNOoBF8ft2XWIRj0GzJ4gt54bEvBXdUAk8fnGbynOru0AVN02D4bKypyYG
mI3G3LeTWrgWxJFjEaW7Wq/VUBBZklY0U/2horbfJXLC71utHKsugWQmqdAZ
ygLS6NKl179UyZPjchPME73g6dMZDmNubfhg1fMe2IqljUq6sQBQnIL8843n
HfoYZxqRdk7DHCQfKqPRCfYMZ3nMXG85EUWx+kcXLHDjQO88Mt+RxpldLeM3
bnrGZiuSU1KyqiXnx+9xCBzIzUzqrrl/iwJq031a7H3R13KCOQUT+IkrByjK
8UuchpPpweok7kdsigxAHPag9wAUKVM5jae8DjenDDi9xMt6RgqnO5R0E5lp
UHvzd621iwSBEJci9OrR3soY9fRVDKB4baEuAxLc3widaS2ykZQD6uZn1jjv
4BxjkUdkEYfYJRIJ3tUXoiS4E/U18nUKYrQVLlex1Gaxua5vF/NEa2/yc3Tq
rdaqJRILf23OtCcXGnOPTXDFL5PurjldNgfYt8u/w4cUkKh19pMLQm8x48o6
XGTcQCsYGqyk3ad6JZQ6abFzf37L6cGLPmxaIewIb/yON9ysgTK/Kn1VwZIA
IzCJgKBXp4DSfnlMjc9Yy7T0ez7s6w0htUrlXWgHH/AheOjEUpKc8fWRYroZ
TjDnMswj4owSGreWZXrpL5qM/nb8u7CzPT6KnKOhAJ6utmiW+LRrb0Yrz5z4
tn8j/LSC96UdvBFoz2GGd9aqBAAk3KGIrWloJ21fpwO+GGgGVYv8XYyu/laA
X51z8bThC3Y9h6VPCud0Vooxpx8PZtgd2+i+EyADJRnQNTFQhkWgfi9ubTk4
hxXM1xB59AyFhvppSvkdFZP9a+tKsWFimRiGIAG/O+MbkIx9mRU37Omaq5lf
s4QptyCC6KvUwQVH57D8GAeTXp6AWe7qafcx6aN3989PLlaoULK20KGyNS3T
BoBDPReEc4tmPuTHMJ+7uYRjat6Ejz6A8ir49FWF1lvdCLB/mW2ydW0svMd5
H1+H3KVFzyLwQLlTiIwTubEDfVC11t/1IQ8tUob4yLlSvvPUvjUW3Ls4OPQV
J4naJC1gRrumx8O7sedA3hnx40QhR6O3Qchpc463p/yVtG62jBjjxn7XLZDz
3eBR5NYT2kHs4hu8hRXtFJxAKYTid7TMhjm7Q4TAtqR3jdtGAAzxDgGX50G/
+JiUvKr0kl4Ug8v7oRl6/srE0aEMmGhwXhLeGYh3gXBeStSgd5SqhvGjYhUp
1AWrnzqJ94I5+ISNdEgCovtWMzkBlJWaYR9Cp/FuAUNbFKvetSA+UF3vvZiX
z+LAAIe6IJ2UHEnJPXVGVcVf8X7qzTm+D5or8QV4g65KHO9MeqW0s6E3eOl0
D/4kB8mkBnJSaYgkR9dEuC6vAsyiQ6YNyB+3fOGDM5Tad3SbJ/N/l8l3SxkW
jnnMF1V7SrKmqyOkeJMymeSUYlKa2Ntc6dbG/WThpwmkzYKIyvcjAfaI3ttK
EfVMUthiCozGIwi7khqZN1gA2iZhbioi6yjF+47gLzef/jAFITna0hCh0BZ7
s4fJNhEC8FbfGR3iDqNDD4lUNtLu/oKg6KK2RB9qmmMNwnMqVrmnB0w3JUyV
oi/l119x+lkisGxySgEBOZ3VUIR06dl7IawQLmdvm9gBvPUDUO+CvLun9K7O
D6fHrCdIKEsbL1ua/fHHWqiyUw4ek4urPFB/Lcky1eX2+E6v05hgrp0UiSfB
DShAIHv7OsbOD0gwDpnrCmoCrJB+EIRQidNb+kl+7Up9KM6yLtTZJFVFobdA
jjcGRP1pITCZjOofm1P5FzOWt/erBNfC4MA4Y7et2IxsjK6qWTvuuZ+HmqyJ
A+l3ICwpg/8c9wfcmp5aZUMpsl4AO+/ust6k14aDNANzEhN+L0hApu8FKFZK
rNayjQT/iFsIbcWa/+npozJmesA/ha2vRLJlbgcNhZ/MTO2R9BlpPRaVX/HV
LQVkNtKE78HY5rWrGEuKMDjRwct51+eOcJq497EOaZvPsvYB5eENfVBPE2Gt
2Cm0gYITEZPnHyrLqM0i5NYYJ+wBPdl6l4Sb7ZUPFywco47TVv9sA7HbTqkF
vFcxCsFbSAzaEacKVPmFDQCdTFmwVfICYPcuoTCbDA4okZ2Wc8vksXli+09p
qgQl2Nil0slJHV7ONeAcArv2s+Y/hFKVJVvraba2Y7d9XFE17qLQeoKoPRqT
kp5aMkBVzixYCDHUlARXsUtSA6/ORqk+LA3jp2sUQVnP2raYcBWiGdNuoWHn
NpocGuUTqLPn7T4IKzdWJfPhhU5IDbrciQ/u6FTGXZ9cQ2/AkmDlDX5GxI9O
MbrsnNz2amm38pFjhnuGB6Y0nS4crfNvn9CDYH1+U/28T+g7MS8gQL+ltZFC
QORTgX0Q8RAoMOJj3bQuhyA+tXqaXtW938aCTxsqszQ+jbN5ML9v7HuKYwV4
a0fPhSxtn+UWas+0TCa3uY5qgN+yz9hljnBUOKj8YIcWBDMc5FqLRFQde6NM
L+oY9aQCpxl7WEmxtDnGRc2tvl23/gAjd23hUBiMw31EN9k2Z1p2K4ory7m6
p3Xsvjlnlt/NRwfVmhltkZdPGklUos7mGEqskcge2wgCmJqTHKPzcYYizFys
AZwHeMIOafkdvoZsVMdHeH9QJ0FTc+PBobbfqaRjz0v/YxSEYm9uRXeS0dGe
xYrGhs1m0Kn28gqArLUIqXImYUW7SFKRnoNQs0GYumpmV21zDHA//tvryf2W
2m6Ztt4BYBZDQXoo8ejzX8hpoYBbMsqP0rP12bORGx7LkpMDAl0L7AXMn93i
4FUiGX6CqvhZLF04QTEbzKYadg4tGvWkh5+elmaGn8n3tFc8YqCyRAQ4h1Zy
VJw3kOBpFP26M5bMsKwq2fUt6gmGennoJRThrddv5uYjFUCi9r0O4O37QOMu
zpyoNgVI7uLUqtmOTFbNIozE0sU7zZm86aXcszTEr5o2NqWpYw7AEzo5A6aE
1CnrziArUtqDzHT4aZrbaXb/585RPUr6BdQJUYyV8rRZ9YU3q15vIBMUZLff
SCeD/+IW62u9JFAuH1akMJsYpaXZNZ1wvRlbOLgtyiJRtrC5NNtxbG/InfZ2
0Aks0FxwTA/kEUShLSvTnH8vm0OJs2H+jN9PnF1eeiWk888PvbYo7AfAH/QN
8F4rlYqLOZDWRmL0/0nQi3NfEsecN3bIo9vq0UNcpHD1yWL4CTX6zVwtQSOz
siYq6vKEveIADFqoMqVixpTu2I34sZ1WDC6ZHPHt2A4JUPT2e4PMDSBRqGVb
Bu6d/IUM5R6AxeoSzq/OLoioxSXPhdYg4zGRfunLV210337SOu8EzJqOVV2S
GavfY59XxhY7/29r//UBYgiZ5bJQCdAbZK5VIFJH6R1ys7lJ+YpKKoYSKLs/
EiUiGjrOm0E0ZQoaotyHOllUt/3YbnFsSlOzoHRRTD5asjf182vlDBZLqpi4
o7w27+db0ABjK37lMFQXxgh3h6YVOPfIwzBHOMUyzwuwA4OC6akKDXZ7Hai1
DNvaN5z7a4ONBbKoJ/d5aB+tk8ZMUJO2J69jTIe9aUaGSOdFoP8ZAOVYZUMu
+eAh0BP68mgwftXUckNxbKlyuDatB+Ob3kU/1caPvt5mX0H5XtOfcys6mKzH
2MHGubn8AXllWgQspEQig0wz3Mj7ZI19UwiCRSJ75IYdHEjZJDyUt6Gghk9A
QqvOgG1Nkor3NqPhUTuds6idie9L5wjWa17edYW1pv0YBO/wuOPDG6akKzjJ
2SpVvPlwcHLhL301zr9Tm2UNJVj7N1MSk1PGenxOGK75yQdEl5RkNkBdtM8A
uKC+MOOQv2W6QcH8+uLQmrImZdFkf4tv0RP2bymcgcpnQakChHeJx0DV5FlM
3dVKZ/JoVsHQyXbQ6UBI2Zrp/jY13otOX5KpBuTom7Iy+fnylj0TuX8c3IPc
fT8iW8gOHnVrEGl+wH6AG6mHo/3pjpWY4lI1xFvqjk4/V67J942hiFGmNH6B
xkiTuSCGvENE9icm8mB042VpIVEcI1LCdO687aZxEtJT0wtcz9D9/BH1qoLy
7MzyhuI+KZGkYRirjB5QpTB9g+s3dIEbO0dTI3tX2GSCsvhzj1TzTP/P9CDp
M12Te4efGB1kebtMNuj+kvQRPS0507FECHBXEevjB6lWWWrIQILv70U0pgqq
6DyS6xfBNZZj68rm/eYy2/pI+kFMYQQsrg6nkFdi/bnGrmLm8i/shpQmClG0
gD0CQvgyoZPfv33CW2QYUB6Rp1m28/ByqaMxrDcnMY0aw6g0wXhs+O1tVJM/
X9SmElJgwAuEYXDOTtP1rR+Vun6X0mTCFT44wdUrehWkv7L9qNGKFTeuaoAZ
0cMlsZNSfWI8DodHmnlpPKgR6EVgND7W9RTo2jQSRTYCx8h+uWuYDGysNlfJ
m8nciADBEGDLMvjLxonCQqUQSJJfZmA0Mpoc9cvZuPbykNKcP68d+9sbZUan
NkXF9sAs/pl2yfJHDrcI9jjizDWtPBhh2PsGCUop3YSwNJVJwliyCU4wu8gG
TJlnn3aQqZ6a/VKnAOeCrKqsD4yGTO8zwtbI4Urwd9aqIGo1k0+rS9Ml6AwB
FxOu/Rrm9+KoX2G1M8tKXXLfqgUlYjbivg2uh16xgR3smYQ9re5+vRaYWym/
JdLIx5cwSJ0qynvpthjrxyBznFsbLFAQD+7zqT/UfA/SwUx1vlUU8zZMOf2c
qmIiC8rDZ+rTdbEEh9FvqgF8vvv93hZhHRGlfQMfdm8xAbgwnm3zbwKFd/vb
UgxC0RF6A4jwKoaCyS/wXLbFfsAHgAGut+LAp4pcM+mwWppNbbN1qAJdmQqj
qRSMHNwHOMt7buwzIhG6awzmPTg7WUPLTdlCoVpZse9NTPpWo82DrI37Lqf3
Zt2HyoO+6d76d/hEDLR+T4X/aSqaEaOVDXet6g5otGMnwPxKOPVAuHoHdAcG
UoqdM7vvPCLTRUq0Frv6wlj4VIPeQ88Msj68BrWQKtZtnr3NNZrNGhnNarbh
4sDzQmwkNPkG51sHwZYomQQPHD2AO8IPWRAlfw4SaVT6w3dgmwWlf3cUml0z
5pOKGoMugOU/+Z1nrK041NYUh+42bCkvDse4QLmGtp7bMd98AIvnHMkt+n+k
z0xUufH7bRvEJR6zHnraTfYjJaelOj0bJPNUgybHeaUPNJxXVLGz1gwfeY3A
yUHN8eCFgaSfScX74asxN3IgKo7Ij1Aroo6AYXqbchC+hRfHOwKgNvq0t/y4
0jfZCUHdjysxa9Elv+/k3Klf12YkzVXVoLY7lRS66f5tyhb/oiY0o0FFSlFa
HulznSqoipvFurx5L1/gpNSQ3GnxrAvWgiJFgIFEotwDdu4OM9nYL9Idi5/6
ga3gxnML3ba497tQh+XoZ28EmymVjpiI2DJ5BqGM8aVZBueBnRCkIpGEnHjd
ZrGGIATiDNW4LUk7oo7lOwHeDsAgMXVXUd+c/JAPMngCCTRudbU89vga30Me
2SZRNq6hG7/H1BfqXPBzL+5cmkgZxUpbIs3IctnlCHJLYsHB+3QpPuoJEGKJ
8l0d9R+w5O2aOD1A4tGUG6mZxx5GGRqO/Tru5PqUVEDV4sjzxsw1iyup5M9j
msVDE26N1dyWuJyS+jkdjk8UF8kh3ddq0EddyNPB30lWtGIh8ZXxaN4dYSD9
DLTT+vfh/zzPJrk8t9YZl/zW9SUWquR0UwMKTCwxyGGJ38Cp9zK+Gd1lq1VD
EExiIAG+TMLi6Kq8Ywp8IT/UKFFpiYEQeNlWGV9mBzVtI30BBMqo+/qLDL2L
ZI031XpGMazEcEi/Jd++LPMlvMtjfcfo7seD99xKSwtE1MkpEefyIlQZZYxg
Qpm+YafNwWf9PIzZFWwgqJZgSVygPhLKS0SfyQ4/4gDHJdBM0ZgxUdeNUYQ1
IFlx6tr02Kglv/bdWJrraglU5aIIUMGlVzhcVFmkunQB7dUcg3wYF0PZ6Hvj
MP9oIMHe057oR4G1EbAmp1TwE4Lq1JfFBk3O0rCVG0muk/OhfwpGC9Ay9skN
FXfM4GbQnWVN7PoKEy0OSXV2VdARIF1rPfy1f59nw57pmQyJjchxEQ4mokC8
8fbHZiOPk003/56MaR5vp8zC97/k3jkVtnkUCz1pR3uw1TRFpkZ51cek0P1t
dtCnF7HWSGbcMXjfUfPo7tfEgFgZ3RNcv0QY0tUUDzu3XOjHUuJg91w6nVTE
z0IFeO/arCzx0pupADRZhWJZuWxWIkCrR4o52DYtfv98DNoGap9kTcQoK8+q
nhafoJDgJP7fIH9rXOGuWyOjzp1dp6FcXDFGAMARftVlty3tbYoKWz3gw6iv
Gi2hn/fGLueCnL75JpbUJGei/VA6Ts6tdaU2EY6bNFkRMP7xDK/uOJBl2gpp
WOLKHS1Q5U/JLequRAu8H3gVoN/hUG3NJpXNXdTcir4sbqpzG4rGu1f0cZfF
XqgyYIoDxNRxgrNwGItve5IqJB8+YK/O0Sb/i1pv5rGyrqw8bCWi1Emeghzu
098HreT3zr/oCmCUajuhm+/aKPHBVAgiaoI6ZOdQ4NlLT0bo49Snj8Rw3hpl
7yfjBYcFi/S66IBNMpNN2glZmic2cLmWF+vGtMgm0kOGWcEBeeWl3s7j6b4E
cjFB9XEE96D3XLMDa9vJ//DUqa8BuHvrGf2fjtudhnfcJKUG3r5Aqe7kUY3F
nJsOgVqNcD/c4swFyqDd5WvO8skTzxzgAiCAWSoRx/MTtSMWdU0avZr3tYCo
SYkAOHMrjU/PdZXl9ZbpX0CG2Bayyr42AP1Pj/McudVpRmnyLbS4viGV4nTd
ECw9rP0drA7kXgJDNlpgMfexY0cOL94ppV1JiwFNc615Z3yrx8v2IyUqk7ET
RNjNKpTGAezLcWl0A0C3EgCl8/s3YZEtz/LFs1nb7U+NbUzECxseFSAGDG3X
AwrHdBvPJdJ4TrpW1CFb53iP9J//oen0nTZxFIfYAtYvz6Tp2DBaqzZFaRkW
n7Zqu9a3FUbWunCYqdEd0BMfX7YF53Mj/wd/zcJ3JSJSbhvm2fgswY9qA3T9
9M0ZOEanJc1GYWPsm1/Gds0LPBKbZdtG+t/rAB57zfrHeaKRnhdiUVZtko2S
gkLgKQ/IfeHFwXcPAkgRCzDcShKXmE4HFQM6RJ3cPc6CzPpi/wJWWQV1IoSy
2SV0A/iecVbx+xchM9dQ64oNBKiNupkGiClzmJkEW9ElLJT765g0o8SR/nBJ
Iwl/Tk1GdMg/CrMpN7/tcABo5ItiBUAXzkjj47bclSXysTede7HpSzr2idwD
isTSxgePrfWG+i6FyLztSRlShH/tzR2z2TIIos8u2sRZyeNcOKXbL9PkebDj
eSRwsz6HIfWMNm/mXNciMtZe1L6xhkg+7hWw+4U4pUMjU1as5QPaf8VL1EV/
7zSF1u8hrNzQowp8bGTrgbAMr2cimFg4RvZVjm07TB7aoxa+EJGO06LhTVHw
sb8CC6yYcH7cEk2DTJG76T1RhXdfMAOw5rlCSeRLwiKfszEfPezCpBeIYdR5
qc4L3S7rrrjEiQ9nJCqkX/1HoYx5MClp7g2/qNyP79iud3h2Uxx7RFC7AWQJ
D8MW9iN8dqA0wliIKfVEh4HKNuiKjyDoNWPK600zhBL0BZPrZ8XrvfL8eXBl
T9Nv996gNh89XwSzIVERE/xRlkNePwdAjscRgfa8Vt7EfFUUU5tJtl9lwRDA
3e14xvgKPgBkFrBEU3dCZRX9owH8l0aNml82EgB9TDeIhp4bM+f3Ai/b1ZCF
vZYF9c6GSNhA4Fvte27eA+4N10VlXoDVlNidUIdrde2TvlvBxdm4J8Kq0BpT
qEo/UiQ91uzj/sDF3hvYmked3D58LqCapy3qhIf3suDzcOUWVF4a/fVhGh5F
h9VNFWiVHqh4Zhs6GDMxI0Vudw59y+p1Zv58ZcMdkqXUBCf5fTYvHxBHfY5n
bMVJKhrFU9oeFoOMl//iQnObM4hm3bVVgySDn5PljK5gd33puXNoowPYQFdS
5P2tG9NJyGgxY79J8zeoSxc8Cff5rftS0RYNui4guUH2YR8oNcJYCRKKPBf+
xF82sXe1ibvuhu0lA44xG4wgw2XL/nOhba5535/ENEHvjBH5JW4PRtkOYu2g
utCVPmsYgNF5KavfdjQeOILaZU2VZSyn+zFy122MWSqi3UPG+fX0ZgZtNV9h
0V0+rL2n01G4Kai7xOS3Xv5Kocf2vr2japYMOrQWKzQxk/fJj/GAFNkaCuvh
H1Fcxb3J5fgPNcVVKa9vjw5McstMXU/rvR686oPWofyj6k2S+MYb/8Un/ln4
bRWoAqfLlujDjRgBt1udMvF+fIAdnMa6EyoDDGGJlumX9HAGciKJLDLvF7Mh
KGJ5uzFH3tIDT36XVfppGMA8zPE7Ev9rqwQBVUY/yIix9TU4D+U7ZakXPQn1
KtKBHpJYdfNrW+MTZc7pS6u4Ye40/uOosVKIZX8IDNv95etbiEksbphEgOQI
S2u6BznrjGAvu2pZKGC1o+T46pShAFQHoEnf/QRR/sqrz6RtWeMwhF5ZxVsl
bwsx1/1FOMCPBg3w/Jq7n08ASok8Kb8x3W9Mw4zd4ygnlYbwHo5GMOaAOCzZ
uCLq9Gp1wMiPmw0a7TBtV66frxlfM2iN9xZ5vcJXHMgpqFdbQ8QznzGiO0ju
DmT1RZvP1m7TmMJgBb3BAiTfd7t6gmyrdR1co3AQd2QicE17z4vS5PrNWolI
kuq7D28ogQQPVdIpBmXGWTP8PCFllz3ZYSoyKwQj7n2Lh3tPicHlvGtClLeI
nDmq9FabvIwitxVzT9urTSyCYxm0xYU65NGHLq5vVuowQpcAUIljoTdwgsV+
JiBKt0A+rcaQQFOvT16gwy8hcwDEpsvcIzR/sEwfWZ8WEnqT3k1WQeP25ker
MRPtSVcSw/srewGcoFt928XegXiVJzfG/pREhdPNM3OGzGO5R6FWfjL3LXx0
AOT6zjGaiGHiqAtxN61dIh5zqJK01N7sw8vvaBXYJxK20Sam8EnswD5RuQID
mYrUeYsdci5wb8a9CyIJ+Dia/no4oUyg0cVIya4SbRi5LbGRRG0hF64+lhK8
pET0+I1HQqlxOUet8ILARTrJTqBgUe7IogJWMnd9pjK4jHGEXFsdP+Fqdo7+
WvMoMPd4zZMopKeh8p8ddBS17HS033iMKjIhqOZCQ3Tj5JAHTYdFmqzHY2ct
KM0Zq+t5bvJcPI1354kldK3/9E92HCFqzanU3ubbB2TpIvIFv5v0qi6QJ1yk
ESSnuHaKuCETd04dKujCM+ZCz4MupM1QdDF5pp0f2V/+j84ve4OOAxjssD1P
1Btwb1CEGI3xLMKzwSlUThfgpzJ0aflIRWIxnGbB9vOgU7jHfEbsQJfJ79V1
k9TpcjSwZgch99JvLTbp2nMqNq8vfelArEUtKS+JF/1Xz0I/m1O6/L/zprJh
kpOlKKT9MbW1p79Nz1xVmo36LPsry8eNmWnJY9QPMm9P37nf4UNC2txNqP7h
DI+tjQGpp7Mxx9bPtvuRMtHsOwVCUpw6aiKgMkkm0WkFtarLFIF4MFdpiTfG
fzLmi6ovnMgD0dSONVrhUrCitbOwHmIZwOEa5aw2GT+So9e479iBc7Ntm3Ns
6roij6Hwr3t5qGHCm040f1USQ/iM5b6fKr6LA2S4bn7VkG1lJ+GUWW5fHgso
VPTTTcW6Ca9q76e4ZBuykHy3upfhqc58+vkCgzmzFaYGP/cbwUlWCPMJabxo
2bal2M85NORh/MiTQde2OxxIpe3y139u76tGEnjxNbBRAVCxPOsZfbjdqmtr
hqzYVS8sJkZcFOmhuMkLUA3xu8j0ZILE/m1rxLiIaWZpYzfkVzZwzZZsjIrL
9pehETVetOxVdW/Hf1V7lakUath6RS9hkiqtnPEyJZni7XT8OP5zUpLQgjHZ
RkGJX0+l6I7jhrdE7ke9izE4gWuc5l/LlU3Gl0lTQ3aEDhO2DfFSKsZZHiP/
yRXsebnxdRDPWICZGbkTdp9IluaHyc1MaAya4BBnGE3E+i3RodpdBwba6Okf
CiPno5eMx5dQNZU7HU0ql9RMarF/TSnepArY/DeoCaN7/b7tN7wx8sdTwD6R
Pem2XZP2rPzY163AaBkqpweP29Lb5EN0+fkh6+pwJCCi/DMyT0Zg+zUqc02l
a6Z/A4BK+3owuYHxOxft6OGW/oekqZRu/2wBlV0Z9OmW5xp92xhm+Vx7SIol
RwvMcXf0aTywFt7VwGcwMDun1xX0ehV/robsNMhvni5HZZbor3ecvq4V5Xfj
TsnornSJ77XrdIBNsOBd/51rWL2GZ0FSGiOar5a89oLz4+CVXSdXXoBTgV/r
ruJcHTywNPX+HbRGoGFBl7sY5I246NE6BBTF2RPxa5Ob+Sim71yg/r+7tQYD
g0z0wtdbHCpcwRbCxxWrSEA5+JVvCJwhKqxxZOLBbWs1T0lKDBZLCse/9d3Y
eljvO80p/EJOD3bh7v2HnxRTpYKQm2nN+CGhJW2907DMjg+DAo1RnI2YJfY3
UfpKTqlKR1RlNn1Hj2gw6nqnngDQet6SsVDQB03idOEuSyQ4RByuD05x0u2c
iJRuurkg5SYKu3rUocRiccf/BAnQnOit3ISE5P1TCGhdggxPcMaTZoXhR2XP
opWJZF0tLJz2O3lTbKp42JCGqV+/WWXbVPtC9NfBGpQku7DVSaw0TPhKhKaG
qLzEeuBh0v+IK3oaJUf4exX4SCt6zezLn7jIjkqMkdoU68bE8gbcCc4gkbZR
RMQlf279AmXEtH8bqfElV1hKO4R9Fyz6pFa+Aa7HxSWGPGtmJ12BA+M+/b42
C3lrK4XfV8BLYHWv3wvI2cBLHTvOUapgIMRKJI76/zwRbRO4T5Pj0tKQcfDb
Var5cicT+0mVkck2gtFTpy5LbEbp5vIl9GQlRtaCyjae3S1h8nBPauPVzD2w
hSl/Kzj3JfVJ9eeBOjmLB4aOSZy/Lf8vqKhNEIPRirGwW0ek7j58C9njOhYg
0T5/ZWbeT2+Acq/eXIydnaPj/lfsUUtAvgkF3VMuJCjzexNqVq2mxXqNwIBh
5/SWpSt4VI9H0F3k574g3cGGKR4P+x2WvgxIOUR4DVRRTENkNLfRLuvGUdZ3
gG9F9rdJZyffErPdq6kLcdbe48tZ8aMDhlT27LbGXKOS+55+VA+efISd5rKP
/pz6FfPb09fbbitVoQn5l5KZJsEWkXxi0jq3fUgwg1WqNvpeCY2BPWguXphS
/GXyvWdV0IcWH8ITCyKX0sKS0u9u3BEPwqddsN/pJYwOCATtix1UUe+3nVgV
CvptyA/69lk/2HWf9Fh2vn6MsYFiJiu446jYUGrWqZABm7k4dWoi1EkQnCY8
yUB131iEG7/wr6KrNecyrveHVZgebqA/4KMKwWHmKkn85tK5U6sSwhqrILaE
bJGBrxAIbEDKpTc1FhAqQW5EucE6iVjc2kE/FDNoneYBh7iY/8esSKU3zCsx
dIAuCz8AcjmoK3Ev09R/iXfDM2FUt4X4sLyeS8t+xzfg2TfbZLHboG8f3VG7
ro5zL9cyfr0rzK5JIusW1Fb3hXrJbmrKxpdk6d27xlDD4N5hiNCioMNofh65
ctM/5x4XrbyDik1TPJ6PmSrqL29T5Kj8FEemRXkeGBCx23jRMlMtSgTj5BdU
Ykv08FLZf5YDXOD2C3XX5/eiNI77Po//qiaf6U7u8O7qcvDLFTlpS6RhoRv4
BdM7at580S8Lmukc5d9PrYNrSSif5YAjBjbQxLVHniuikVvvxglOKsba3LaR
4fgDN2u2olIHAJsmuDPW2rXchXTTQzrDANVz5m5Z8FZAExQ09QqM82wWGLHl
kvhYhqFCiWTr+CiFz4825jZ1tYZ06bFz4uN0OZVmCI/UidsHXqjANkpQYf34
sh8fYd5Na40H3cPeiz3Kk9v0FfjsRzp3qodukUh1OI1sgknF3j9hkrITwTy7
pSfXYUL8pw2wg3E20otAFHHP+OdabGvX01NYU3mgD5OuYKdv2hk9nJhGTmIj
NG2QtKMe/OctWxAUjYDLkiEvp9UWtezsc0GKN4Vtd2PoNqZ9c9dlbDxZ8U/z
IVlYCPIVMXJitAOgCw4dOCyXfIVktJ4WMqfNjiwWfwTX/lZ76axqTA6Jj16p
O7mxKsL4jcUrVxQ14ZLcYnaQloZwaLiL6YdYWO36Hy0d/Yz4wazhI/U8lHlZ
0ccW5qSPcuWWBefa8MdvymAlmXJpmCaMTshxqMD2ybYeaMI1joBykWMZX9NG
EaerxPBVMl8z+77QmLklNku+QcCY1e/MRUHJAbot/NuIgbRzgKphKKz2tbz1
vd07KGtA41NHl/X5oGUelIS4v/jZds11xqSJkQFH1XX36t/MjaDVeXANVwv+
wlO0Gqcu0eKmcV/+ctX/GPANv7XLsy2x7p+i7yu57mkMiSKVH35tQNCW+Mv/
g4mKEZL1sWMNsfl0QTOu2f4JAI3LmzsGLzhNHlvx/Rp60/P8AVBseE3lwM7+
1P5PilEmCwB9CLU0wVhvnf4blgmm3Tlf/aacssVGFZDLFYeOo+zxkn8yJmJa
MF8I353JN6MV0ntjpAJIupKgkolrFxfd/5H2zwQBIBxI4zymhPJ/mnploMus
kAxeC5mGdbuGed58wmawRbdm/EgnDMnFwg/oNoz+uyPuFirWW0OFLC5fnX65
XcUu7F469OXyUaGbk9yOOedEizHv70A95Q3qjsGGiBJMNmUVs76KbkOqdU6P
UFIXlF//C7Kr/6C7JGnS/frNWrl9WuN6o2eftQmoVFJaKWOJAcAvepfAJjz7
VNH8d+/wDrZDgIsLvaPaDGDEkclswZ6ZfCLefk63Vaujz8cXkKE9iJ7vYiC0
KCuWne5CwOUVzUI4OdQdTJMdaSxSxtvY7kppwJBJQ32WWc50EPFWDMUjCd1j
/a6eMcaEkJRucvpLo9JfKNW6TubN/wg1WQIfZYVlQfYynch4Lk81CUKMJFaz
ZBGE3K54pNQaRyAO8F147HoP0snLLzbTfhSqZJySqWZy/CqbJwxFyGQt+Y1e
C9paSKtUT2lOm43cfNmKCg9RIvu3L4g2Q+UX4dRlmR7L03azPgx3E0tXvrtX
NwQ/7BrA5QlIJy4btGE47pf0M1ypHtOsBHfuSqUSf3EwNJHB8v+DJArlJ5xi
qqhq+vAh8ylGJMk8wV9J4l5Hv+gyxO3pRDt0ich8JLhKGLuqElK089tJIQqX
yGF32CpaTnauCGI9WRSWj8ZAdjwciOwtXZhuLi57qQRy6J/aSY0f4ykKOp6p
UwC2e6hBByDBB74M93tv2HHpO5qBLV6vjfGOF3I3DBPwEqhDvJoL6Hw9b/cz
CIHHRHixVfLa+PohYJNyPcQEwr1D5DvKM4HRYacouZw5ndweAZES7x439mXc
q7LdIX17lEbeQMUHeckq2WabWeedOd/X57Gx64R8M3OnSpItDd5isy2qo43d
hnALaOyt2kL9cbuj/4EKIqTUJuOMvS433qpvedQnOjQstFSrlfpB/c50or24
n6TP0HI7fYzR4gbX8auq3c1w7ptSuyHiCLP3hBY4SxN2bssUW+AVZYzoAUBS
cM0gzEpoLbFG1SmSqh93yQKBukhobRbr2pFG8VB3GfTNWfb7GnD+WMLprA1p
qjIigoc4OXkmmHm+JhZqPTeV1yHOsmi1gdvpCC6fgPvkmSCVRdeAAQqgJu2L
oyTnb9MDCGTYbLj1E9fhYFeMohl3mKbJc8QBPtZQRgpL6A/rKk3sZPc9kTdP
T49zgp8pRj7Umtq0Ku66QyUSyEzlHtou/njM2reBBR9b8fUxeEh/Q3IYvK/A
0qIJ320QBwt8ev1Nfg94M35qfZ5shKqRmZDv1jq2khbSFXMZ5RpCovteaiCY
nhzrfRGMYEk5sGgmKO9lt7rtTPFNk5epoVWCI1NzJYPRmrH10g7QeoToQ7R0
yxwVxMtuBcd0adTJD9txbiNt2I8iNa+KY2H3kAAca4nyYH7Gk2RDeFIdpT+q
K0+kgaOGMeuzt8NszJfuNjYE7+jHxJxaJoaIQ51euoKX/o1+8+aJRRHy4Mps
bDgJyz/xKi1APcsHFv7YwZSJD9nt7gYL9ajTmgkkGxEYLgwa/+Das6RlE+F/
Xk6Ok3U83gnwwQgmevcJwm+modMKcwdGdI5euBWohAPT228NjLdCs8BIullN
PNaWJUocQw39oyoxHckkAzp+gmB+C8pNOwZ2WtPd9jSEffZN/HqFNCF4KjkY
bG527mDY/LfUpIajlqI7+INUKBdNQq//NT/shEAZZNBiFaNJEVzDweOoLd2i
IOeDEQsKRJRyJMkYtj9hPIFX69CSrJ1gwDiFFTsJCyCMCwN5GGFVR/xfdxx7
QBdwoNwVzVFN7Z1rE+vhKIsP3gss3OuAzHv8eQ/aw6sZt/LadEzJY15FXff/
MUqdV51Rz+U0f+xapa0A6wh4mHwXpZdpy38zKHc6yWgrKHWJ3nOjc4pyewGa
kWhWGHYFQpFWFEaorLiOqwZIphKlUliiEyPbJvUzJc9FaLW3Y2ggXNUZHKu7
HDz3JiyG80AZYZxnLSOEH7DzDDK9F3J2pcG/DcxmHKCBMyBdinVCVdFYEf++
iI3aLx3+AwTkcXyUAc1FYtn3+Ql+aWRZmefoxsjEQA6f4fY8k0NgRn6ISsUW
5XTnPv82scFQcY5hEhVoXqNZN2LaWlFr3V5fcQnhrbUvvxxRCGE/HvYQbpgf
xiZz8mV72U4jKcbeKQJ2Ug3T9V8jQfRXzLxVZdX/VpViAJoMc+gS265m9qTO
yoOcaGdGqnuPdlYhQGAYS7nV+SQ37YQdG1ttnn0Bubps/q32XB9F0wcSjx2q
eL59ifMXbvfoErxEc8w1usJOYrx42T/peFM7o+5TcKhkuli4vFhbEczgs8/B
Y2o49l6aKGK0irILUnErjKn30y532Lp7PXeNcLDy4p9gT0IxszMPEWyPlui7
eaVgn00xzJvo/I+14Xlm4j0wh8XHWro96rTGmc65IyBVVDGD/MqAp4t04vVm
jFnkK+1lYXuxqgHpePtV64XhSNeuDpKVUdV2VTJzsyFZqNSd3Kzs6EYrHTD2
MqGrzf9t/rnCDqLXmYOV2udxIURvVcumCLdu7tEcaqGBe29qYlvWsqmoPnNK
sOZxKJUEHOg42y+9vb5fpJLzy4B4MkHtGY76oAape8lYZgxfcobHjeszN2CV
/908+ljv552umu0v/5pJ30RXRsk7VY93/VvVCa69hvIwNW5/wx+wZhHxXpQh
MyU3S9Sxs/Pk5iqTu5spdyOXRPaYH+NhoGX5cOKHNZndGEi2IS5o+iko1Mue
fC7VWs0DP2G7JXwGJjyMYjgHLcSzOLJLu4NQSb/3n7LRiIox24zhPsZRxDsu
Hn9tM/HzFfk5x2jmVruc2Br3KZt+u1metRCvKdCZ1Zitp9jUyLMcDsk1kRYo
T+VEO2mYjaoMKiE6m/GH5CMoGJeaInh8RZAqI9rNRRlRsFjWrjN6+kRYTbuN
va+vXN6CZAkrtdkzqS9S4RqcmDk53C/T3Uzkt+lzHjCGRFKaWWGUpSmp41fT
UoiK8rcPk4K92Y5ezSHOzv2+SvNIzDSUJJ90UiegAMnNo2yOpmzKNmrmURqU
GKuCoC101Q7WxkzyjNH8kk+YQb/wUiijsHpOcv9eTw6kPt35Q7VsBzCoq/g2
BhH0wzAOFYBaINbbYhRCeqgRlfZsqtQjz10FA9i0Tq27B1RozfP6JktvVzK5
GFKUHTu2CSbme4nQzAzHDfdBPnvst21yokPyclfEOJ3OsBzudXwFWwj8Ac5o
pVx1GIVKiOcKus+jV9MxVkXaCga6yHM0zDI+Vz+k6mze+2hFHWI7HFPTfJR1
jCh3Hio7Xw+WZkzfLku9baxS9io8S2Y9WaIbeLeqlDpRfmIrx0tvUCTv9KAb
T6I629Kx5/kfwxVuCMeNuKx932vSDIQBNmKOHby6i1FkfbNoMkPq3Dtexeho
D8pXercvicIpWPCaVgKLfmfbYxOawcmO7Zj+Tl6i+WgNobAunSzNdWs3p/Tl
QHYWL27mDQFQoHIf34/kNoUBUc8eHwXIYceBssk7EgFHQeU3ieTfKWtO3FXO
6l3DaqWLgiuMisvHKp3/a5eIffNYmqK+mQNKDV8hHuYinCWTR0k36Kgrf148
0nL8cmDUjkbZ6n032wbl9txvGiLdWzimt06pT0sHlphCRt9LVb9ZEuI8ecDF
JAmfyNK3QwoOxj4IkG8JKxxz3N4/QOSajcQuZcasloXYJ2xR7ETmcXFmAWUW
MYv8a3ydlu2GUcjfDyCDrJwaXmtllWLHudpl+FQzzFNlAy5N/x1fisnGINBS
q+MhFbwdpB08rUjFX4t6Mh0Lvf2BszBh33swaDCapZdAfByWOjBvNKhXNnfZ
syDHbJ5gcE3xtGI0GL9xuxdCJjsq8l8RzR5Opz5/bOJDuX/RlfDiT7fGv7EO
tVyzWOzmco6K/d2p7C+hpaRG2oZOqCTbBEMfpLHkyRshSDiBcozEdtrr2NlL
Im7Clox7sVlR1mk/H3KulukRbUpqHNEY+PTtfDEZU2YKhysi5J4RnWfARAyt
cstfIve4dqqpDEC1HJyFZhgo3vQ8gbLiUeAi+4k+nDLU4yqI5CSgvK7In0P1
CFBPQiXScxFhv3zvT7zQGXnuhRhTU6wiQP7kcUDRynGmOmqZN97YJShbhj3m
jg1Savg0xmoEQEcHGAc86hDQS6ZJ8ds31nE7XQQmE3z10s/Df27/+OQ9355y
NIQIbKa706KperRW8NWu+7zKvcxL9wsKaZogtLyIHCZb5buE0g3SQfrT+A0P
rTlghtwdO8h+bbRJmbva50325fdJecYuWtvO3F9oJJRl7lgq2wb70P06hoBq
/RlG4RXK+Zm4pXPegcrBCiKrZMwb8RChraK9ERUrj+wCfnTHDOgxfNaR4Clu
NeMLWarEecYBL2sew5/FvikjKEJ4Qe1h7wWWAXTDo2O1sUViNuQZwA0HcNO5
EF4Kg4BM5VOeuDF2HIBikRkGqSGolZFj3qPi3Mkq7lsOGylFb/5QUM5IuoYU
eCTuVqxTs89mbmHTvKlRH0CJcMRxE2CHLMHeAIGqrkdWLcrblXMK4dOk4KHP
OlguDar/Cdf1+YsAujzyyiqPKwVRGZuIja9pCSV7ubHtkGdwj5ilAPQdi+IV
ihZpDoldkLQM+B2mxk8L0frIsM1D/FUJsZf5biJfdWvrVJNLM1L8Lde4Ttyy
WBQPjh3ZdC8Tg/ZUJw6g7dqGcDIaaezXYkHmc/2CuLaCRYId+y8RrYWxGHCt
x3VX2xTSJ3yr5m9hTAljZ40QBgLAgtp35/CbHknlpyGbN19aBM1xR/XE4uZd
2hLQee/ApiZLJw06ZXUwpMWOLM6FPILWwG5B9Cj/ngbrxLNK9UVHse0CVw7d
vM4W/CUy68E9FzWex3yhsG2w8hqwxs7IQsYbvyzGYyZ9DPzJ8CPvkRyjYWvv
vSfrZfLlRS0yv3IQ/d4qOqPhxJc18Rf7TVjJ+oJwS1STZDpxBufmhVMYeRym
oK/ptmODQXvC20jGg7zwCNvfZuqgkQ+RT8krgPbzbnGWZrqjx6VzkMxVeqQO
uP+dcQVVTOfxPc7rtKfnxdMN4hXDV/IUR+LXvDIUJ08tEITdpY2F+id22dGC
c6ucMHnF9qEgkaMKXi86elzv6PIBQJsj4Yx6up9xnF2bIUMnHl3l4U6FpOFZ
XqLz0vz5Zpx25KWq2yy9FhzQVKa2yUtG6LW/rjZGSedhrScH897n2gIsXQ1R
qUljzw4s6DIaGriByZsCMFHdtI01EtRLUpYy25ROJaVAH/N9TldLnUdiQSas
pgquyJt1Oh6GknqWfO+Np58igObNcHcyclTwcRj+1cQ9GGVcSkDiqQRIgPbg
vzkSz2iFH/bvw5XQ6n8FCnoKYx+EokAzk6AWltWZZEKqnhDV9nQ/PnDeXAsH
LOo2vdQWJGQELmxGT9BzIqhxSqd3U8INzdFRId5mPBvvHXkbGdoNIX13oO4R
7Aa2Q+4QnED5ZQpMHp7zGhSy5rCHV17utznTYmli3kiw0jrN4qH15k5UhgCX
7kCgKXR39rDjES6ODE38AJdYx8ZZUXgbbaOZOUsd7F/swVCvzujLhzuKm043
zf6vaSWnUoAQDNQ6kvACSz0QBqpgHnmTDuyKCxEog8gNga2GMMNRuO/tDI9S
3mH1JQO5DsfxQqYm+lQUZfESOIlyFStzFSNdJIkiHJ817IpN3IfULR3+4uN1
gRqCxN5wxQQmqAX4Wg1Ze3dmOj9QhAFwVYuXizHHtlkE8aQKthNbVUc35X6y
yJui+PXfB6s390hiPKbMLaaRzSzxohCZ8zrGbfOzxUcX8y8IF9ANwIh9Xnes
U0rMXrgKWmPy2ixMrgjBYkeRUrnK0PFGEhRK9vGPUynLqnSChwF5jPKwhWUz
Oy6Zb53vxmmoPcKQHRnvAnbupO7N7jJS7rPXjkuo0HMa7BQMwwk2jlXJLGSn
0fnGPew8QvHfcRkbzjUI16EvqDwkSNVi8ro/nwK7FtIkfwNGP+5hz+A5XMwo
PE7G9oM3MCgR9cDIVLRn2ZRk3Lrgwawvwh/js9qRxUaBEGgoDs1T+7C9PNSO
hNt7SlvGOwyxJJAqhGki0nmjvErAUsjocLKIGAvLZG4WlbDbYavTuIZbqg1W
M3ADf5GvM+SAeaM2QHkZpqgGF8l5ICrgQvdpdeVddWXfvSeBU/RaWv4pGeTK
55kgsEoHrsY3Vv7ALIMFjTu5brldeNJGEQl5VH2DCSJz0K5ieIYpd5Pc2aiU
CmDdDDHdqxE5pRAmwsGdOzBcbxWAGsTMRIFqCIhfQmvwrwJqrR2pEBxNm5g7
qwbkSjX2FVEQiiYyHn67AfXFF9StTvwWD+7lSPlJCdWYh8h1Pm3wiakHEI9J
74RM18YEHhp/ZSXf0j0NxVvCzEK983XYLK/LXN7OvdFX9+rIzebR9TDwMtSz
3vejw2WvU+0L3XbNYJyWdlmeZV0IDvC9WQKErimkyMRCLhiOJAEKWPMx2J1E
PzwR6aH953XfGPm/y/okvdZcTt6vxRsT3xuRiREjDcJb3jAlSxnd8hlxBOn2
OGT3I/ZdRPdL9LlikRfKR/zV7kItsGVE4lQxMLwT9mAeaumdo+5BQfBeRWCA
EKNcg9bcyALog0yWjvJgeWM+J+B2kQ9J1BKqmjMVNyEmO3o+OSxxzBthJTeX
NoURGC5TZQ5bsmSz34u7bS9zp7H1sOm6VXcslC2NFPfi/x0i0FOuAeMPeeIq
63rGedH5+UIdgSOCkkaHwxjCX906sj9u2nxgdI1p3l9YVYOAvpEGVPSxD7kY
7dnfmyyLLS6dCbqfjF87muGdl8SF+6lIidM2Mfcwa2KgqvSlKIm3jm9hCsdJ
2PHIl8SPiOcdMlLgCqLm8Tnyfh5JnxRRpIWgSs5O/CA+A8OtXgaEkDUC1y4I
Sre7MWWc5q6lPVxn1UeEZj/Uo50IuaZsc56/8pfrylwQnYr1gGGbeNqEOu1X
ZucUsj4kuc1JnNxuCM5fTlNp7D1MxmW1qE+FSvHFDvBnL22OEjJZWx21EiyQ
weQ7f4UarCIt2ucxKrkY5wwAtHA0oJDZlUt8pOyRic37khyBqnVY+ykgSuk6
HSM1Ea/5ip9MzqM/NXAhQZyne9FfoIa4ZNm/TregI/ASSA0G+jct8/Rx9rnj
aWnRx9bwpPTNZxspwtMLNtFvbN1Drn2ca28fbhJqNzl2X7jh9uURrW7ajpyw
aoanA3JG03QsPW772PDCD3ikcK6Nf9WU2MkPU7YykroY0iqe2btEwMwIDW8f
UWYfMQYEyWxkV1/L+PYBXj+OQ7/fMq3EDs5gnUXbFwJJOuA30oe0LHZlE+qT
zs/khL84yYCHekgABdxTiDyxfiQWAdK+y7m4WErGHTslUrKWWOCDcqHTo/YT
PR7eiuWkZuKvQPtPLjGG88pKJpAzCqkRirgqZ70u4Yr9qeV8VKdmvvzZvsHI
3+cufHGn3gOlCISsGkDXyGDFHVwpiFcrAMcLeSBqXI9y3zjX/1a5JrIXLjhg
C0gCfHMJZL8/R7+ej1mcn7kI4WTUOmtVRCTVK4Frs/SBHsSLyDnzsfcAb/94
xfu+DAhOEtNS5s3lImDj0us8YL7FvbgRMc1qLHqkxys2y5YOrHgqI86hDjd4
OAChowG1VNnl5+8eSO0dOWC2T+ipSeJZvAPcvrJUUvthEu9HlyGzkBORle2+
Ww4HsCW+xd7OypK1eVehQ2PhtgwQPIOZdcgM5r5c9nr8nN+c6qotfpnxXYCa
pjMyJPhSMcm8oD47rwUCRiBLGPzimjjxHDDsAGfrY4Ji0RO0ECJk0HcTJANR
YDdHcGPia1t0Vkttr6/LGSx2CM5DVjuumFvLmO7Ql6jfR0pNkbuFMxQMtO/M
O2l5Uq8F3u+pCp0Q2yxHJVh2QGQH4d28fTVxga2DP7uHC+77mEgwqH4Fsq57
dbQ4SutM8Espw0k7jZHV0bo2UzpToxR1YmHmj2KnCHGkgz8UVjIPqVm1Q4pp
d0b4oVYFJyrU/TXiX3wSvt/zI0UNwA1LkZAj+peYhl4ow+x3fnz5zMRyF/63
18fhZL1Mh1Pn7ZNj0tnKTOBUTgmpf4A864yrjp2JVXq33b/3/eE/DfNNwTjk
Ew3eJwXY1KZgfP+EGVhUdFeIz8N4UMl6zxO5/6BO02GvXXi1KBKXAgTTUbrx
rXgZq2g2RBMK2cR343o8JoLcqWHOq/dxlJ0Y9bYfYWotsMqW47ysDLg6cRsF
+HXs2kF+wOOTl/nRoQWKMMK+BzG4gL9FlUFmE9H48p58AUSD3FfKcEYun/Zn
agvI9z5fE3aM8tSACxtYPL0S8FBNMxVdlTkLYwx7CuHghdrxaVuBebSBlziT
f+R6f0c4tx8rB3rc0f9TpqiByjhXcb0gMc80l65WLsrn9Zo3u/MDOYBU6Iyc
GEgQjA2aDQsPa8S1+XGKaM+F4MHc2GtLJ9scpiBBZTHQIAiWB6Pm03JRNm6L
hP8IkYTd3Qg0lS7Sh68DMrK1BVbPB4A+sgPttF0XD+kemlUb56xeLwKX+ca1
ABIC0PCO/W7aq1fWRENtMjzrreWueM8Z7rY9YODuJjdbRl5pdVGIVE+WIbsx
kIMeLwD4DFIDSSheGgHl9Rnm/MdoGajIgMddVQScrlbdJXl3K5jCYIYp6yew
E/QlhlJtv5t/8h5m09mXR1vKENI2HPZI1qUNZy5VWD4iGz7wf055f/gr2SfH
lONuQvKXxp2gGw+xW3HLvyPnKQCvePPOta5uqRiRjXE93vwWPNro3jzjW4VC
Y2ow+ylDz/VkVM3BwGMiKcphUqRQDg4TGcEfZ3saKhzC4V7kE3nUiTqCl7JC
UnI3slZiUIku824Pgy2xqzZeWZkl7elnn8Qb1CO2DEtU5GlfbQN6KImuq7yY
BfBue0AgY6YTz3J8D7B808MLq4D2knhwsy23H3dj4DlDbSgWZtJZO9GQmUJG
orUIWTyJj539x36zNZ2HrCwY2ILoj6L3duZlNP7qYKM2R0IKynTsL+z8t/Yf
ojPe/BmMARSF2WV5cYFfJeyU3mAjcqe+lK/f/XHOAXBJzQ4TeuyFUiSrNAra
BMZ7e/zLBFw8yKOqmj58M9mQifvP7HasveoClmNkv8edW6t9v0f7tjr7dzqi
TOAOyMnbn8EiFERnPbo8MncjkIeNpmVwfYINPbedGW1zHcUfkBHD020A0eDj
+gTsX3eO874+J8mKcMR5lMhtR+uaM/Y1HrYTtfKq8p9L2Gu0C+yyVPxAe2yE
G8T+BlcHGZf5czvhQacUYvprz2nOVaXiw+Pzpb8+/wwKobFcK/w3u2ve2CE9
ZvEbstrFEfcLcv834qCmNnLq9k1A2Cj83KLhrsDQGELS7YNlRP2+E1ZYJvFe
TI3fPea4wYuCmwhSblsoUrmPZ/E/hY4LFAeBeHMyMMppdSmTGu+RbEiH6drO
WoxHparvypQGlC+pANs3v5oT9AkzIPXTTjWfwYY5IldRBSREbkybo01Y14Aq
woLtEmCR3BGbkFn93j0/7QR55xnADDqmEo7Jv44wZ4G8UGRiCTo3eEohrOy0
fXM5RfH9WEDUs1dE4uKMv8t3Pf8OSj4gtlkfqCF/hBZstOjA0nbFwbB/dIGD
NE5oXr+BXCrftEonYXpjd+/81iqhPITXljdyn6pocTJjv3sOg9zxkfhhD9+H
/BiuYFEoh/6hBTksTp95UuIVmLIeH1LyYYq0yVWhgjzSGDHw3sHeIPin5NZE
5X9nlCw38KHVRvXyOIG7X6PVknMAGNmYlxHW35jVNQXsLVXcnrSr3Oejmegr
BeCT4Z4+zhkNH2hkI8kastMwEG7V2TwBgP2RZ/Fto2cLUiifF0N9ZOVcCUAJ
mbsqgSnhWPiJQibmK6qhKghbnGh12weiMlHF5oS353cFq2UYl6B83LwLJZ4Y
ePleAABIkJBrOaHlmQzfGewcN8ExmW3Ger0TJIqPEpwgHxhPWoojrmsAWw77
dUEexkacCWPvnraonTi9pc7P7Tua4gZ23DzVV4YbS11TKiosa+AvT/TuDlcT
mEzTGS5IbmPv2edMm/2eSyo80E6juoSDIhEeAItp+WZiPaiHuqvuOgSnwPEq
u9dxRiE8o7fcc5likkw+mM803KFVBmU3VfyD11prwNLww2DJ6d1XoyA0KPE1
hcKNL/bQD1YF2XxXiE0HuM0SejcbvhgGwT19hqyJcb87VFgzjx0MBLEp7KNc
kAGVACVHfOaL/lM/ro2UDUX8IP4hG3oLXoGcTdFo5NBcBJGdpGZI9dXFZicy
+owPGYUZjhqWX7SG1IkdAXz84x7YAZtOaz5+4gK6+NIlrgolrgM52Jn3J763
sOZ4MVkvqTw4qnGmHK88dkFoO4cyLkOqJlu2IH756qho+NUrehXwABGVCrsy
AirYJYSMjCwT1yOgT3BQ20I/Nyz84L2lMN/UFMAhSzeYKdYP3lR+I2h9+8kN
EGVCfQNSgXSkFeaDTgDt10hloldsKjrbElFOWqZ5s1xsfg6GVdPaQIK+Uouj
hrygSCmWlZAuLwf/gkY1aCFTELzAwmUlRBa8V6JrRDrh3ziWdrUM9uSrJsLX
qAE7cRiBL1wTVzzzOnd5mxG8k/h9WP1cNlucKERjJrBobYYZl7+KoI70EW7D
EiKQYNEgxkU/1kZA25D+BVzm42geIPV2pzvClGNc46GXRBxA0J+7UOX+eTkt
3uD2VsyFw+8zYTy72S1egz/A3mDnfaUMRqFZtdP9LWrPDgmnoLN4eL6ZI3K5
vDuKssF9Kh8DBKQec2SAgY7EFPMzqNX2ywUfFS8TGU0ag6Klfl/QeI/hKuv7
iEuSYoiaWRuFWtW568Dcg2kfAxy2p6dvn09arxEFqHRo49+yfSZc6SC04pSG
X/xqunf6JMatF9hTMYwz+ifHasI9Oa5tJb2vwdTDuuQMfM/yJbN59ampShXw
9JZd77vk0Twy+vOXa09PUDcVPRCWItOoH/TDnXnWE4pAylfPwOhkgMdeUPWK
hR8osYHeiPly6U1DmdlzdQVSFJABMs3mXup5WTWTQigY0SIN6iWqU2E6Bia5
PMjyNoxzc4VzCN4rRdSCynXj4tzrTcyrIXAhcSMozaf5HuSa5l+d+W03dkUa
X7/34eMH+G5SUhWQ87DGVKqIiTagX9uIjv9ZaGy1LzlYdXVjtqvGnWw7iGP8
LIMM+VoyjyQLjqBITDVDDEHQhmORh3r49tfyS9i50nl95WqvZy7z9gQDLPos
mpiqnIeJUhITK7Gs5Y/6NLALH77JynwuULxYqwm4xKzzBsXgqnR/L6+p9YL6
jIaHN4v4TkSOiPJdiqLmtkXmBoatdBLqthlaVPq451IyKEtkrUUfsGMjABby
Q3/hJKWeqk4ISpwks40Rc37/SuBlb8EE0TGhqz9Rx4r6ulMArxaJjExmh97G
VFcgicvES20g5BrcS0fCBCCqGnc3JPasHOISCtugtD4bt5+3v6andGPWC3y9
Lah9PPUX778HlLDX+zCr1ovr/jal7tvqry7V6UADDhsEYDYuR6s2Sy/o8VFa
yEndbwzapMUC4+hWki2SfXR29WXXnXqPIs+PVxxGIGNqSY06TDXqnY4nZY37
2Oj+R5YwMHj1b75/vMQGWdS3mh3UgQp/dUuEJinsoKFujfsTG8iRzluxxf5K
hkCnBF4a268PrHd/xPpQSgvLq9LqBIygOsVaigXFqvWJtKvKXvFmarXARhLc
hNcuLi8W4mISYEfBEbyWC7z++Pd9ji+4jBiVE3qmS4tXXhthosWefIjg224I
vN86Lgt1w5T0Uv8GlLM3narzjgec09JWq7wdg5ELf/SiH0rwEtcRzMK6jkeR
Yw+E6fq8pI+4PFUYituwC3d/lsrVV/8Psj48PRoq10fD/vi1Gcrka2Lz0hzh
UzHnH0hxu81w+LukeJsQw8Q/PQyfvLAcMUSP1piqUf//UZBj1YgFSUOlpr3/
/ExwtTFwHkhqHtGf68iCYDiHn3WSykFmEGJy8Bn23C95eTicaD4wna+5pZw9
B6HDK4CgHAnni3VpGHH52Lf8RXa6eFGaHWAjpBPt3rMFNz+Dr3dxjz7EBd6c
aBRHRZzj4fnMuMDj3EgP1KApHxep4D3o3pDaZXBaIiJTd5/c1Spy+lMHRRyc
ICCz7H9ZlFxiHYS9y6xb3/iEMtpUV2cIo2Q2FWYP3Gv2tDoCj+B0bjONh9mJ
+bZcFVWrewom3zMir5EDaD3QlIH3IoGhWAV+kNldYDenzI72PjZHgosqd+uO
5uVso0UMKJaeRwiEClqcmtArANOHSfeN8jck9lCAXoeZA/2DsabT/AB0+ZHk
zk1ddC7l1NxOlM/HtryhNvFwcYacEXqxmPhV8ZramN1hWdBAviU9FAw78ueK
HzfrLU2bpeFhUMcU+041OixMdD5Hq5Bp3piR3O+JfgkuM7Rig50suj2KaVLT
TZ2/Ct9ebiBcUqnmx0xPP99NPOHD36AUAgyO4lOAAhIVtdz62NbNbHfTDfK7
eUb7NMckTzR7P81N3jjQNYhe14P291i1GG0ev9Y7GM6S8ZT7UbzZ8AW7SAT2
vcH+jRP0sm1HnlMddTwBSlfw/T5BVxGGefVtInBT3V8m5E5biu61vsVjsP96
yJyda6sGHh8UpjA1/m99+kgAwBxOZeRqA+RbqqGL/YBNgDDJaMBqiKpmNWXu
R5+0unPjlxYgKw61ZkoGfdfqwon1znFDvOjTxfiY/7Bu+CrjfC9NdMlpxZNP
mbnPHC746w8mreolWWHP3p89J/Pfge9WMReGp5yvfTqHnYeec3nyBVzKtKnm
d/TSfR/vPD4DvijXCm1ioZ6zHw42fUvrmd/33S6cFi1RtmsHzRVufX2YES8O
l2rFol0aJA3zfjLw7i2oQ8N9GzRVKr0vY6KrtP0kxAqpYqnPr2lhzXinK4z7
yKtIkZN+wogjaUtF+abS/xeGU9kn5+9dubQQ/V7GFbck7HmxoadH8S99kvHB
dNRgcmrJVdIjZGmF6B7kk4IHSkZJQ4tAG3Xo2fGwzuGb4z5G5cqcjgFI10TY
bw1x4w99SG0cFXrTrq7vuiNrfmVNQD5/yR7oLNKnSm0iPs9yRqN+9ejb+CWn
CYZM5CpLSBz8swr7aAV8R/xe4vPYQ5ANsvIjL+vCpYyj8BGhLrx0pla9UpRy
zQ7G+ngaTT+itTKfY6/PP37nvvZT+hvAPEk/Z5E2A4mNbmOvFzAjAihswkSk
GS53TfvcwXQVvaGMMx0McPEMVA+6lBKr+JzePZItQ2ZGkQJvQo7rurC7E+W0
dXZVl02VHOfxr/+FB4MrnNzwcVfkbweAM+HkR7bczSDauR/8xY5vFJmWz+gO
UE/t7/cIbZzWEODL31M5d6p88/2app8XqMPdK922gpNyq++/Hnw44X/OO0ke
JpiM5lYJ6hqjEpnxUmKfQZm1N7RDPUQbSNCPxuHoYGKN+11IS4wMHrwTe/My
66d3WLMtCiKIl/UksppEra55SlLurtZtVGvPjm/N6+BCWm+BAWHV2wrd0JFq
izarLhsIA2CPpir3L6s8kASTxtuZIkB8s14lrWsicsJ5buvH15NKuXy8uUrm
vpHuf7SL144YF1i70/FFsbJLnCFmg5P95YoGsNftWPgWulNI55m7jsQru0Vy
t6vZLV4llTRWlebi8rmJR5Dng5iz4XHv2JdEo8Wm6RseWcKV5Y0B13nC9MmY
UFz79yWAoWC72wCPPTCwzO8CnXYnbS6HDRqwaysPWxNrEWIk/r37BPksSYqx
jPtAz7f6L8lNwGeIJiC+F29g0kaJMXQtqQDKWWmdBA5z2wVydSS6OcLlB+mC
XEGrkaKs9VkY0O07u3B94wscm0nFnWnuqLToiPdBJi3R022OmN32VSYLG5D7
5suazRr3L+awcBlcMiFKkUqpEOdv+Jzqu7nQdLEE2aGWtNpgV3Ne9bVcldjG
v8CJLki2W23a8iC6pcPKkTNjrLNQq4+EBxRbA34neDPihI9Z2OKlEB3gNPGD
T9xn48nsTKJ1w12teBK4SVn5EWwLK4erUZ3OhAnCxDoZuL3AaZHQHRmhzYbF
FVbqxB/MpGZN7BrC65swXEsn92WguEp3pt1sZhdHb5uwK6cP9gA0rH4chTui
alFG8BqLVXJfA/J0h/cyBo0nOh9TMntJgiYL2lro6BJ8E3wEj61OfblTBUfw
M5i2c4247jtlmuRxja13CXJigQCY+oQLddq9i3CjPyyQeXsy5+k7KXGeI+QY
raZF+iHS/f2JaSALAHQC/CPN1MuOlyq5/Kd4eAKrLkt9XKlG03lfr8Cig+dr
vn4tMGNCpa5vRbEk9Ooe/2xKoHiZoT8XtxGlZBEVesIWwOyHnVHJebpTfE4T
yGva8fty8UUsgL8mCww1X/tIdNAMqqwf5vRaMjAl+N0cNxiCpM7gHPJhNPfv
sVe1t7cpAKYzy4/3mPMepQ00BuTH1650KUM+LqqzyJdd2pDsIFrdp73AEXgj
MOtusDgWOsJnO2Hxln5d31DeHT9x4X4bt/6Q3hXs9mnf2X+gmonM+cfjCsLH
SetT/Qr9wyAV2co5SmMJx4BC3fXiatdjorRzpExXIZm70E8HgpDe5Abw3JQO
jm9IczQB+8X7oKSDLz1yOQqlSPCA7FlyKF5c1Q1FBWtXQMaH6Trs/I+34/HX
WproTwMn+lF8kIdw+sQufiurhONwFiayHBGH9I3RNh21xgndPjuakU2m1kdl
OqyUTbOAu8Pha9imzSMY03E0X+/6YFVRhwKWqzKnBrgPmjpLj9v7TEfowt2V
S8p1T3lgUNpNoEHeP3bewndj5N6LpM2myZcxoDbsf3TL0XeRKIhjyUUXlUFQ
hbE/PcF88T6VCjk8C6GyjZYDRGK1Z8asU9QIcvbT59TsnB+pmCo0cn5IhdsW
YB2fGHbhl/R6RMzeEm+BTHCXnc1Aph311wWcD+BQDOtngwXgnbn6Jtwiz8uO
H6T+xnmM9Ve7sQPmii7YVS/oTkfDhTCeY6j7vfnkDxC2ZO6hMB3+qbBJ14hs
ELDcdxglJHH5bJL7cwuGbjmmqccCIuuXLkW1Nrcx1cp022YuaPjXB/8Fa10O
XPpcYKspTbW3IfOXdwlyKV1MfyF8UH9Nh3tbh+gbgDO6fA6jBhVl76TTNomV
95TJbOBnQcjnrYeuRyuqIZEfU8eWUVllWFf6GZ49gZ6wPQb/6mgSl5gGKaC9
MUtdyaVvERsDajR/LfhXURveXuUcqRKVRPZ30fHHg6imJDp1mGsA+vLzkRjR
ezjmyZ1irXMoT83ze5E3dhabkB3fpi1VRhmNs2CbnOAoa5uHjHJapH2XSF2W
lNR5AKGh567oFopRT+InI9uoC6tkIVIdi4g+vxvC+cG363+AQ4YnKmZxGVxU
jhwmzSTZwu5K7D06oJVIL6/RoGzXgZRHd2Q8Z8d2ywYNclUYpG1qrd+JIGAs
SiWZF4w0OyN2tOOU80Y8q6prptWVcmxoYCNXm2gYuE0QvWMd9XgqClShK4H+
29Wal+UPDyy2XuLo4n7/pBZfh0Ea92gKlbBuEhNl0SUFw3fRBmGD1JG5wb6C
wHPhcIj1gzsnDw+BQCPcOv/Uy8FBYo29+ek7swhGd5wRa8e9FO258Pmi6xNP
BNKQ1xVBDLqg9oQvGG6/hc8Ect+S18JOpDIkBJ4Yble3nUqom8WrJl/L0ok5
DcpNSJQL9NksNjX9d21uVyi2ktSnD+d5DXNaYBDUSuWHPItkvMlEn7YAnbDP
VKlF5oa2kAwI1srKfoIhoEmW/bjrfBxIpiUNgva5/6TkHXuLnLY1xuVA2TW+
KGCoqzdITOC2qy1IzvG/IpUqF8KBO8mDIt/jWoHs0a5ZAhpH9uhMjGmJjCOG
J/LPy+uNQDSCANhh7sk7IxzKo0ax8KeiWXetVn4N9wwxKd/tl1O5FQHaY9nM
UqDkQQhRQbZODD54O7aMztz16clfLbgZIxmAlec5VSXXsuTh4cwgiszrhwFq
rAn4RcjqQ4ATxPl4HKyVGwrrsVCuRYSd/0zWoa5rN0tXuPzTNfGNYNIq80xh
Vpgtxatol468lXxWo6laWQi0UPD+B/NJDdJ5MYO+yFeNgc5qkU5OuPjTtJye
bWTj2fyBRVoTfhLYdHzx0jS8BfP6vWrW0g/GAObEWdqfDA3DnVN2CpqLweLC
nI/iUnSbvti9oSnc20BmQvfkW07jhWCdo2TGXZkNB2wCaK62n73aWlDtF6fz
OPBteiEhXPL+UfBLqYJbycK0HqH5YkVxkseh5NZgcS6ORZl8RiWbhuOwMI/4
1E2Kazl38Bebe1dT2qUznVqJYutEAe7m6of4r32jdxZQ5hcFhnyXMn6yALbS
3oyrqf7AoA0rqCovvFPww7ATzOcfa44a73fuAfBwnwBI2oSkKj+aTtm2ljmY
dslJjm6RrgpSKpEXReFLkV7FiL3RXqVFZ1jxFisuMLlBwG0muEortgvozWBs
1OSsmT+rUTBjkkusE48WJeqW2RS8v7rtoI1ZjpYuRf3DLJiOWHV8hAAckxzR
9AmAQh2h4/eejh+/1eI403KVYM1QtOJb8kkZU2a3dzgD2QB9sVfcbaYKmTDv
PpyQPadWAjYaQxFvkYN8mHj9pdN0yxoUOsBaqlVpfhagVOYX6Rca3qrGkh/n
49mM4MmerjOxiyH64psBJpvowCMs3g1hiqXl4dLN37V93I+hOCmnNLoKj9lG
JltwsUcwHozZSivlWCeSu8KHpM+IYnGeA/xeVzSJQxC7tXvewdVSuCdkH0e8
TYdr+GkDp2O32VcvP9xFDTXzcwP6nFJOkBChfU7QQn25DIIZg/ybaYUfxAGy
BmA/XyhCmiScNNOu6wNTA1YtC9yyNYoftziBah9BVYbxOf2a2FVEUVqOpaZI
wJ22Am7juanGxtsLEGh6k5xmDeke+BglLxsWo2N9EFAxp21mmy/0Y+D/bxam
jbJmy953tjX299W+e1sHulq2teOJgiifvY3QK7QweIh101PLa4GMCFx6yLm4
kOf5gkNdAHfB7eboqVvWRufweRwo1MEOaLMhHzeEmrZZfDYEv9mlZWlCrrtd
EyJ6NaaenaKd9R1pIlWmqH0fBY0ctjlozKan2vcfSZpB9FCY/rZRBKQuTzRf
om+AZo6HG0f3BOU+AHVfw17oMHEhbWM1EfOMOrqLUwcSSYP77unJ4NVix9mU
wXS9/fAleeQOS3n+8kMutCyRg643L2U+RpftQV5LtCZqw7/n9N2HNH88MCyY
v4EMi1WGlZgL/tVTAJgGMcygEkqzODKH6QjY2P8k/fj4in3LoVAVnXnKSeVL
bTEi4qyDE0aW3z5N3FzFCUx8iEfTqd71rrl4QvKtXTdVYSj0gNMZNuztQGw3
xvFsXmKBs3ZPK5qSGk80pOmDpdIktrBuSOVont2ZrLYfq1k8ZZ1DFTB2SG8Y
Jh8tPHCbqRmxRhgRE8Z5zfLYCcZffwZHHGk7P9XGPdQSxAUw2ZYk+ucS7oZD
IsbsMlex2M+78Q7TJjJk8ewVwVkI7wKqOalqrVOP+BCRSzcanmaapuuxQu/i
i98FKuC3WTZvQUzL/w1XbSaO24fJkNXNUyYmogL9pnh4Gd+FEa+1ZhUzBkEW
/aYPPhIirvEGtXoX8avQ3UMEmCNSK7ID32Z9Lh8Q9L6RCFFzfjpE/Kk8p2LN
54n57FjaQwP6CcMGHMmCdEzmbRxGv9VEYXANq7+hfJUpVcg6GUE9zjQPTb8L
z8Kbit4KajT/WsbeqoUj+Rr/UYBGWlJlt+dDHsOtmfiVJC3jI2E+IgVDz+EO
gSjtZr/LoMkSPTvjMLQwnvIxHMt84dvU0CrBTWzcRiReMoBeLo4SlDPBFd+r
ZirpzRdGOxsT828CXz7xUCJI3cIUw4/X/G3KJO2Fubf+0D9D7vWbX2QiPUyE
ddhmfM+XUs46M6nYAuG7NVI3YGTNDY+KBZTiInenz1NIOM7yeeoByQXYUlRt
j+FI5nrfwMmdDJqi2v4MopLOZ7EnyhiPVPK8IHw3eqbdWqDsFTmNw7YUiguB
LWBbXQd4JR95MxZ8b4iro4bij6u07mMMHpLyCmSyRQxUBDRwgUdSXIA0p/T+
vB32YCGYTQehyF1klfwNO/RGgvvYnMAw8pmswajxsZbOTi3eOnfhSVTMUZqd
yJsS6O7bIPSTi1hDoiT1lyzL6vGjyrwkNprwUIvDClkGCaoW9tWFBs6iL7cE
3RZIG+6kKtpzz2ayuiASePeHMDdAhIEukRoiZ8dynBvyKXYo9wXIVRP1KX0p
OklB/k4naAwJDLC+bN1TC3BVR9N+4EkhRx9mgKuab8o/ceQuM8QqgABlTD10
7ooJhKpEQvW/TRo2cvfNEQRfI78SyRdNGunfCaz+Su/LuMR0CtKbM1ItZSTX
JJXjZjMSRT0UCJwjH1YtI+ExVBcdQxjE7eS7M7lgZ2nrWAyRIhLaRPXTOEkK
axZcGAuEgP1vEoLj4U7dgEL8JvmDNp8aewX6alI6LXd7y8rAOtTScQSr4RVg
6H243KEFl/tRMaNSQcJuFn6HEQ+IH1PjvtLZyk8I6pb2OyQlUMWo59v5+hCP
U0IbEmvapqxYERmO6KRRcqOf7xDT2KYFbdx5Hi6okJ748uw28nvX5WoTzJuW
sR5PYJblMAZmZ/gJL9UxIoulnRGvJURD6WJhj1+jwr4gn3924SJbeNJwzsEy
7snG2IlaFLNpOPIyoyaFlQlOjUZ+iHWUPYuVdYGWhjuVFXYXDmQZbiL1LhXB
IiN4s+eWvXqh1Tv+lRedu89y5nK3FH83bLk1Me/zce/fGa2kwA3LNxMjW41G
xtt/Rykj8Kh1iTDQqfbXBXokddetBxKHWevT4X9AKR8HYCZiPsPNNWFdmXJi
1CAJjN0jKQ85qGEW7dzCyBcQkNwNIZUbw9ZL5EGPKRI2HqfT0G0z/q6ezVmp
Hxi1GLVeVpipAknyFNudx9Asomxqx1E/3EDQgL8w9O8DHp+1B1KXa1RU+QBk
5wj6SsMLbs+xA/4PQEDAdkG8pHpeFQCGWNY5dbkminLcu6NXUSrMXnKko2cR
hfQeoyCgyqTkLV6SBkTbsOTygpQpcje+gAY3JopeYt6+TjFTSuxMjgvOFSsg
JxRBUkLK7aWkCLDiWs6WqDPzFopbA8TkVyr6dt+5270qG/+Y9Lq5JEWMY//T
FPFZVsXpUpkxKJFptErPuVVx3hEF1El8uNNbBlEck528y5q6vLwouAuvaXuh
XHwSFsTdCRoqdTxoR9x2DUaS/ZLmQdY7q26fhDHBUo/wcMfFcl+9qtbqoXtI
vG+nqS0mKlgjdKXApHe2/XXH/6Jr8ae042TII1gnMDeHu3juz3ueSskMAF1C
5xI4cbrTan5C1wMdimtXJKURLIpq0WiZs3mcIEcxTS9+08J51bdOhIUq3rsS
XllmNbolShWeKRyuXBFinI/nzjNlLU8IjxigICNzq0YyT7DwIdC/FiHRpMNM
UEcu4OrsQNgqssRwiDY0XGomEFEMBTiKNdCxLCnW+GGqZ8bLkQMU18Jqmpga
edfJ+xi1slltc+YAzsWypDYkrs4UEEAb1azXJBQGTuaPNNapidpOk/ufZT8t
3WqqkWbpb892kW4js8nAHudTGOjwK3gkq1KSPZ3fl/ldXHaHGenNXQ2cI7hT
phZS7vgrFbB6tIVcbUG7Sej2bPz26zWXopvU+f0MeT5kuEjcUn1oFzmBviWK
qNCdsgDtbT9cqVDj2dzFDWfWfv5hGUYGVKfqvx9Qikgm8ov+4G8/ZM2/e74g
8ytzwH0orG7+Lp+nr6nGysAOWaqgzGqeRl1cjcyzYdgtXl4Abb3Bz3IyAM7b
gSLb4S1p4+taqP6ev+6vLF7AzpAv8y1LhRR+SyDnPgJ/Zfq8xaH4ne6QY8Ku
YfooypfLgO9O8SCqUNlp/47ITk2sLf50YF6FPbfeOGNCGeF83m1x5hPe0V9R
dMktb9qBClHlNwYylq9vEhX1O3GlbNZrxSo3VjpE2QKXIoX2p9LNecRWxtlM
7vZxJW3FH27l4wrwH/o9TpiVVDG9yh7zdOvf7+zx5oy0ekm5ScYoEdp6GR+P
Gdp7x+UmpG6Al0FR4oloxv/cJ6yZIo7VAyXHI0eUJa/BChIUeJnc3Fv+zMar
UsIAB+Y+hYXajAh4/3w9qeNzHsiCGJcgUU9RPWfj0JPrFH76FKXRFGB9R0Ho
vAiB1kAqa0aK1x+2WkF4j+ffpBkMRVuui+Cc8Qcv1IrAbQLULvZDlmFc0qPv
PW+weBCVZZdbb7YDVWRCBe6ifoW+G9888ahQ9uSp3g2bWdZdwBHF4u8k/4Ek
FHOL+ofjq6T8FrpduZk1N1v1FuQHqQtAlBCEsa5juO1jfQVUKgbutg6ojENj
j3xCKompPE/P8DIk7OUwv1Y3itjCuGLH8IgruBPHp2I5uMcQgduVQ1+cX5wn
Eqs4F3hMw/x11WtEpJGIWc5zSvXZmWN0T/5C9Ex1Loh0iIfmZ128+RLcNIC0
LZCIsAeB9+BVXSv68SpOkqOy9rkoJq7RtZtOAzTESFvUbDsC7+b9UtcL9SM0
5CjbT+DxqqDjvmJReVJaEDN2z3znR4S96Bl72cAmCaPhmOZmYLvk0fyoXTwo
Zvb6QjHS1gMrEWhNqBnJyA6e21oGfTV6Ho8/lYgf/JOd1bAib418Hk9UAkws
qYDb9SbMsGOXKAXQ1XCcACnTagbrW+jvUZoYIhdQT/XfDllUs/91w29TNR6y
ZUdXKWwfZIHygkId0GFU4IfUOnXB+jfPsUZ1RT8s8pkSyCYBenuB3Z9m6yAK
oNBYJWoXTvagbj+g664TK9vqmtxLAXCwJFO6JHXttTt3OzWHdRYtRAGGCKda
mYsyb5QF9y7gZFZnj/gcwCbgGUa5N2sEcy3d5IpqpJtgO/dZqhNK9GfP+hjU
jCt5VDmDPDjdyomAK5zXITONJHrK3oK+WHF/yh29qmf7YxKYaMwyQR5ZbbUf
aNq04OpwUbgRTiHCZ95J8/IJ6VG8Wppw7M+NeiymZ9qQum4QeauUZ1+MGReG
f1v8I1Kf3pfaU09CYg9fEE/K/F1ucI8o1g0BORSGMhUdPwIxHkkHP/iMrrQw
37GXlvsYZjiRY7s+RQm09ASowPmjMvfERiDer4Xm2iHIeMYKM+3l4knlnSO0
TrqYw5uX7kpZjQUnNV30CyrNsmxar4kavmZ9JohL7celNZR0w5R5TQyUWCaK
Pn2ABZ3T4kAbIew0Ct01kheQKgn9prNeSvZ7e/XUrI/J8JhRXXLHMdw9cSWo
p4vfnoWMCBsWOO6ANJm0NRpD66boPSlE+NYm+yn7wsv4mRFJ72mupkETHKka
fJgJbmpuIrSX/Pw1zHxgr0tiOYP9DIxmOqSNPrSvHisS1cS1v6KQDi8NHuOv
Fqmd3eCNfaJfyzD0fYAccf3rT7L0shw3hxcpK2pizc0GIYmC8rqdUo49o5O7
kQATUYIyXAoUPwJgZqmRF81C83pTJTe5VB7A350g3p0hF20XGkBuN+1YmrC+
lSIARK1n+OIJdWRyggqjQOqSDfVWkJl74XAXLG8oldbzVZ6jO6QQDRQostS4
3plG+vfsGUeNMSnymcBmFmeBtcTheIpABtyPrguoM4OUzSoxPdIMCdz3IGuu
u3UDDBl796JxuNeBB5OEWSygRix0EYVVU0830ltggL1duqT0sVp6d0T7JYBw
wbRmGDEvlu37yD7CHy7q/g5DEAxKw5reP/kgrfI2/JZTCUWCHNeFlV+E72Bh
PmTvsUL5UpUkaO7RQo+QGMMH9bHP63bAVl9LWLVlzfkDxaK0zuwuPTQg2gpI
Bbv+ZEnuFjzrYPbkTy1GRe5OY83diB79sXFkyQURClTC5JT1eSBwD27f6BRq
YpWnKRZTJzG1DSX+aVSmWnqhPrvNZAeIuzW52v93gMOamNyjlxxKytkSNge/
3kAEnl/Jsu3SECgTU8eZv91/4kmifRxnnXZySmTi7A3FG4wvWTmgC0l1ZXqu
Z2DUddwfM7rM/Gcm9GLDFFar7qB9Ca6KRwzoyIxeWuSmXnIdB4KQayV/r8Mf
lF4KmzCc83hM5LS//NtLSuwisUY1llWPg0fld5TFE5J9uy4cyZfv0OW9Ot+M
2rVo3Ya1Gshr0tIvTlkSuSlNHhhRQDEbjqdqsElmjVbwY/fCj05PXAfllIB9
t9AT6FYLtdA7iicLXtvbJBoUihfAvSL0Z1nUK4skED00ggrCDgh2S7ZaxbWn
NVbXOYecDpSlQtxUulthG9/IfYbxJ+6e4QBGFpBCvuqKguSjfY/cCszPa3c9
xQ3hpS4+iCbVYtCDJjVb+gpj8gOzfkyGUbvsRJlT4ImXqn1SavAT8uJxNTok
VQaJGjiew7g4w0bGWMp2GWfvzKS8Gi9io6a/PooxCSR0HaIL8rZwjirJuOIp
5wcUbCkqkPLXllQmMdZYfWATnH5oD2ZIewZkBs6cgYT9ZAm72GAaZKgsf3Yw
sZ4Jk3ZVtti+zbiCvG4tOg7R6E2nMx7Yg77W/HlfMoMEtMmHCmI6LbXhVPZ/
lURFx9ORrWotBJuOaBQ/NevKrnuDS7Ila+wmEV4zuEEtRPK5wX+8QYKDi8BQ
IB0bx8NpZGy3y2mdRPJHrzdgfSu9SGKx5uHTa0TjFOlRpZzpcaCoxqAf3D4Q
JHvcwMT41WfFdgv9FJ1psB4RYChwVW1Zb/8n1puJGjM4kRDqwUUatgxnvJXk
e8T94zj+VS1OdV8h9EzVANeJOPg7IsRsb1uenLK9MypkgKG0OyjdF63WLR4r
mhAj1fWIjhpyHJaUHOfMUizBafnXkB3J4h/8nx7H78Ndjqelw/WCuLgJICKm
TYCgmROZr+UqJLqtf3oNtGC+n51CqYQG3LlmgFi2M0ZXjyzo1IoJ96huFW5B
KLj+2dEqYVxGCJSIG44I1NAZInelv/z4NnZDRnWYtMD2isPF+zZWGGncMp77
cVxnkot2jGEPN175WdvOJvWBxFlQlMtOWAYRLCqxEyVqK4m3CJ/2VD7O6GCk
y3YL2gwIuBgh7qs/1WgftMqkIV3O8Xck5zEyYX32j2lai60ctRjb3QFD1q8N
byUcQfh8ERKP1JY0FeU/s9adpfTDrXXv0TkEE6ZDwi7orIjx/PXzikNC0Pi3
g1UcNLO5Gr6Wj4ZKtYHtUdAwygggx4vzbEQFtxI2rZQUVMX6b5ku5odrYHWl
ZENueO7/x1/7xGJLHFaMYsPKCDltOYAXXXTKIJ5LH5x8lA54NGmfkzQGWp8M
+INyOLDCmFusB2Mawiwjd5QjEtLJRejSZFPbFkfIlxiVNTs3bSZ4zuraPuaG
W7wJa2bbUnaQT2vBxyqRkrdzUChvTNSIMQwQb7A2tclvTBUyalLVJ3tcaesN
mo+bIUs/mH7NFGW4zPbHHcMTxieDKpRn445PrgpAvRhtk4fCSsEbDZQG9qdW
WDoCPExN5MWXLmqcfMMXnt8E9f43Ozg9Gp44x2sTXMwxAPEa44jlPVWo7ny5
A5rZTYBYxyG/PsktZoQmecmWs0nByRc3CIYdp4URoDFANqO/KSlaCtp3W3Rt
QJEHhRxcM92yAhHCZr+4wV3p31dtXHRarRAHNFtEbk4RuUDuWmey2AMN4eXn
Bh4dQ0BhU27yMINc+uy0/abZF+fiudoKjMWsFOjHNSivfNvjeT9HUrGiIFKb
r8WOKAiWXZrda1exDxhEcOh76NWOWBJ22X77CoSWuNk6QUMHl4bduJwLdcgS
ZnoofO/yaOcgi75nbYCUw1C6T5ni6y/6eEg2t7I0SCC8SOjOedY4D5j+85Dm
+5EXallpbRnRAA80MDZZEvgrwp/B0MKKxEGJK0F4TsNhfASAfIMyW7d1j8gU
TCJZ9WE++u6RzhNeiCQv/jkQ57NckIqCXPwUzTFgSPY25dkYalOqkrhBQ57w
wLOZWkzc2lSg6SflWLKi382m7A8xw4wYGiC2m51y+9IVXoWSOptxWeULE+9q
S16h5KOMhUELBmlbjqMVTI2xLtjyGS387GKsq9soAsW9GUkvB6r8HpQfR98X
ndn+VTLxkp/yzGASr+ARzE6lBA3fdLGcIDuIoD4koljQDd6rjPACDb2ts9Sv
EOZ2nl36VrOp8hptMGxAaezdc0zYM31HrlOm8LVxBIUNk4uF+tRZHQgS8gWk
d1XLWxWL9ZmgAU6f37FIGRbwQWCVQiCgZFSLsgKfx119pa3bq40ueHnBl6hH
lAMLUHQJH03KN+Atqn+gnuf7LtFyvW51Y3xGgK56YGhO6FlMfpiBpqPDO1e2
UUkoZPXP/kU7nlKXoFaHEX2Ez3QxZr6dQMZwkayxYFtt45T3KylG89CcbHuD
Iu4knY5D+/ESWxEb+sV6aFeXdrkUOGYjq3Z36fqj5o8a0O+xn8+wlHFtChkP
T/piHdhHfe6R2MunhEY4Mcl+2IE2iY5gi4F6H5ZQnO0v2jAVrBQ9/Ke7cp7c
DXky33kSfH5CWqfLNSMSit1GrUIb2cASUs/5egpZ4zQFn1+Mi8PGYqoCVHeH
RDifV64hodImz0jXrmC5Udv3OokyP4pT9+wUKYwaXgqX/xNwjUPSK7F3zqxr
7FJMrJG4kON4aUNahP4YM1nw6fhfz9GEIc+d01PiBLtGIYllu7w8jLEo4+e4
03SWor5Q+Z8T1kYGUgI17uFIxVwccEKzWjTQMH7NbNgEzbDGrJxZVyWBHq6r
8KHvdXOYiA1MgLHvNBWgW8+wBaKwHmVTMy1nITe06g4DIhRvZoFt3KfBuddz
Kdk+TroQ/fvqc9L9lYaoZapwUw31+9G6Q61/CvwaoQIGDtH3fzRodOwyv3ty
fB9fquHxGHWAaVuS6kUPK2n6jPK72OfcRV0FGdb9qdC4VGeTCkLg6oTVU9er
+/Hpo6JxnxsVgDOy0MLqKbUse5Kv/5C7l4MRZrKS2MXD/fRdr5bYr8C0WhHr
fMZijU+VCVwuK3Zf9cmvlAecq20kG06swVggbjcN2yDT1N5aXkdIj/9wcV4o
FdRPyRC+FME8hGkMJiPqAatttOQC1fBTVV0vgHTTTGm0yp7lpJjTXIcvsxNE
AXNL6HrNUocYEVqOMJ2cS0UKIaBho0SOTLy0LnByhOlWRfyJepmt6aRfVQqY
Ey3N1GSGMZQZkwlsQ4X+eWiEP2+HiyOmsoA8SK02HX8s5tcaW/t+9WkNz39N
tj+PYKULmN84FD6V6JuTEjklOEnDXQLTamf47tgKn8CKfqiqIhtZFh3ewBjb
JarpjB2IoccSPOwapOZxy5gbxXa9mAItYlM3muToECGJDLAcRTZb4mnbgLfJ
RDyLY3AX7a5pu6i7T+NMK0MthB6iLDFXxAFe2BBvMDDsn/14gPkkq6dOnmU0
llL88K91Q+pd+8bTetyH1rRKbCTsKkbUQcwZyMNIhfn0Jyc+omqQ6oXY96xy
kT7cq/UaDfPO7Jq1LX0dOuX51p2golOGLncK0OUEAtQ9e6zqtMjovow1Klju
63a2O+KXr1tbXKR8uRX63tq3OgqnapqKtw41jez0lU2tgOl+dXaLtUuBCk9G
2OC7ouvr95NzE8ZSfW/FPoRf8RTQi0KY6wwQKM+rofNWxs+ZCBGDnvYxdUGR
NmpGveQMA2qdbI4hjcjYTZXv4RmEOn/HQiog6nheVXTKwF/M20EB5p/K+YS6
RMEEsebJNRt4tOTC0ozNH33RRePluy/7gSMfLzab+PFAPKMNbonXnA/hEPIc
hK6ey1kXeuhx/n6vMnHOuZqV0cF/21jVc7saJBdHnvA0l9DHixqMSketb/lF
LDc2nII2UBToD9mp4YY7/WWC372y+cyXYo16x1Dv4qXfTiX0B2/A1o7ljd6n
BTZjcljB0LBKhwiKHJkuOEgL62nqoAS6cVeidXkVgJ5YvYijnoHdhwylrjpZ
XY27IE5dF76W5un413DLlpFr4UsgmoVmbOQusg14lLGELIRXEis2pSo981gk
zXjts+LhzFk7lrNLXpkOyeu74ffCxNtcFT+aBOmREeQw/Fb4NtBX6FuC05zg
VVFQMOdYJnrv4Tw0FFE8x1S7jbl2QZxIgJzm9MSrc348p1CIVfS2OizY6TWk
Nw/rAtjfZ9R2+9q1DSHCXrkXVysR1/j1/OYm/OX7Edv2cUU6x7Lqc97oeBRg
p0rSZW3/HpftoCZ6Ym29eSgKCHkHNl/v/FyBKR1kGVxpMAyJ52B8cf0XoVQr
WnPgzpX8v50S7P+JkrL2eVH7o1l4XBg3nn62qo/lJ3mx5FnUM4X00W+6KpJW
YFYrjPDrOs0rXpb0G+F3lK0DxEmPQ2AlrAB6aMUyB9fDR/jbAf9KGMvdYaSj
U46FQrsMlV48Qkmr81e+sNEMlp3lKokwxipYiq/qOlAEMKOGguaWAJfZFxMA
ln8n/CgfR3412gBNTnoLVDSNt/GpQUlU56fvIs0BEfrFmjjrVkqzB2YS4A2Q
EFIw9kaFECKS72gnS3cJkMe0QduM+SjQYahtJmTohIPDyUffDWubJXGw8CBJ
8SOdK5R5b570VOyadCrcu9YD7Tgi2mZvX/OI7okzQudj5anWysQQRTZGqijf
JuCQEge4rbIpck1QhdMSSKv0ok2I5oDGQE/ylPtQbM+njbKZqlMiUwllL1Kg
0ZSL9CnyuAz0dr9MY/48cUTz3TVCTOS3wTbIExJNJDAAvvjxLtfTvHE9737G
NmO0oJIrYWKREeh7g0jLtKXq7eE/1FB7VwCG3ZXyjJV6+2ndp0G57iknit4I
y+FB5cqHjDBwyxX2Y7luqtGyO9Gfa7rVYh6VKVAaBoXvsMUyzGoKMypW7F/C
qLCK37BTvi246cSalPkTVm9BXTY1ZlAdtGpZIotzCiCAeCQ0SQ7d0qH1Fqhf
jOX+vxVnkINADn7v51qJ0EPHMnLj647CL6Kps0VRpXIZYK9vzYQbv4hC5nWD
USokeBh+dR0wyDaztZtwmFNM9NHlzh1L4nuxojc/f6CweXWpd7GdDjLJksPP
LJ8LUEHrZISQYNkXrPdXbBH49G3GrZEmu9kkdXNs0Gw4mkN32DXBpfCv/9Qx
npv4DP7x8XzGElgAX897fc8tbuv+PueSP0ekyb7nZaeZ/tEDbZfZzFy3cSWk
4awLrHns7pTeYsszWUt/ViGZ/8G+5wyMqPxw7McCxrSm/9+JgKapWhthyZEw
mp2/GhaNpVIIXUCQjO7VQu6XT1v94M2KzvaifqR+Xw/+Wo0z1N3tYbQwbxh9
XF0PN8c8lr4PmdKAxYZUnoqsykBtLb2EdUptc4Rf2+BSYSHGXSZKOSsS4mGi
KRFMF37myxLsS/7yOOJyEa78PELmQ++q/aHa66ItxlZWAlSZFNQTBvrUCL5+
hwqGu44SUlP3DNkwZdlfcckrdBq+0yX/eIOSoyExpHtNA7HUjpJeM5TTlM1l
u3M9arTSkhI8PSvqGTY9EO0whKDxdhOK2be21mgOT9LgONNrVOGCE5XmYOhG
pSrilJumFXEdiW8aritlAA/xExEb1jwEdeOz0XpQ0aydL+CwMQthMCpZ1SQ4
iDnsdLAwoicaNS6QCeZhwFNlHjJV8hLy6OqYaeot7jQiW0Kh2Au5Zp1vbQ8j
BqinSZLcNY+a68JGRdPipB3+qRgEUdfx2jgVFbzqK1e/TantKBqDPNPdl40+
0LJAcFSm3n0MC5VJHrAWwn6hIp+wvCOT0CJzujnxFcTdMUBIpCnIDzqOxzLB
IAyrVy87PGFhnqLLFxbiw8MZpZ+l3j9I9mcOQ0z91auC81PyOw6sU2OuTuuT
kJNzzKA8obJ4/AQYGFEdADV9ZSO+3cBUAO3XAiQcoML8FtAKCG+8o6ocll43
pKSBSp45Ps1CRtYQvPGFWmzoaUX8q8kBgORfJjjHtV5d7I3CGqNEqwI1qZuc
5NsJA7rxfkohUWyJTNALTuYVs6ZgZ4MxQQ1NfrHVKCv3VuSxCjXTo0bbORrk
mlJCm5YU4on3MQ/qSbagVgzDXi9PwK7qFYb8dX7JRyfhePgUeLduNl/2XWb3
PaMo+83f/Ksr+2ILoZbDpGb6YdBwfdCFaeLYTD1T14OBKhPZUrDyrR7zh0Gb
hFrxpnKdYIsWV5RArO+57dMmqrGKb8itRtgWHSi98n9lGFJe1dDlCQVqDxgV
5bv6ZczgveDomAItEv4fwWf6jEchQAYRTB6NLTyLZYREXUjjIQXnABazXc2+
Ho066XkHEhlYYQwSDJNqWJZBzVdnu7pOFSH3GYaHmUnWT3IzybEJOWzPKXhu
6DlHaiYnNZtvQmF/O0AGqDGnMVU1Yeav2/ITP8FTW6PwoBytyhCTK62VvEGt
+vrsygvCpD2KUAWsWfo4doD/R7YYpGiGDNrZ486WZ7iYEDV+5NinlvNZ46s+
FW0q8wLqDsB1d6gBky4HvkC3VQta5NHf4rm0KrB6l7DR6BDeLiz6hRkEC4dR
EGSRDkfr58U29Ou8QAhbQp659f6m3vfrarOZgs2iJ+hBoQuS3QMeK/f3jpHH
a9Q5enxQysqqUA3yXe23jNXWKoXFZn98RmtVkOrjMrIHWFz+JUhQjvcBftxF
sXLTTgQOgZGuPubBtIf9Wz1ehUScXd/333TuQ13uTEh8VtuUi5bdRH3BjY4H
ATL5+hg7q6zQcbD0J8fsi3JUekOwWHwt8M4+JdyIvL8FHLWgneiNMGD7kAUz
3ink2aLUD3D7HpIu5Wsg8J/lIOKTgUqs8cyHQZJ3Xt2ZpbVFn8XTySPCNBWx
LYjSQMLcy54G4AC6IMvln1p0eSnuJOk6OD26dl2YXxBCERwyU+9fTuVwuyj+
03+yWFwyLLGVgEQXEmKC8+yAvD8x7kCfYoTR6FIxhEe6JUz5pqxfg1SoYi2s
rifrOsQ5lvKSSiOEi4R9DFxPrWvWtebmlkEo+CBTjxi8SdG3A3tDCf8lWXJY
fMT/CoGR8bqOEr+m1gWzJX1LhL4dpn5Hf7Kd25xR6TTouli1h2kUlW6o4zin
HuEw28ZctKJqtxfT2/zH5JR5/885JNTSDNCQg7BY9qJ22AsDr7X25pZ0fRrb
ZXq5NqTzJSKaH7iZAkgz8cgC2p+HGL7eoydvddOk0OQKjz1AUsHnsG7RbI/3
O+j09K348u7+6kfhBfeAzYYnlNM+g6B0AuuGHq1YuvqUQ/79pnN7aXzqrQXr
EtVETt9Yx1AYmcW7ZIhK6FIVpuOZWwlZrYEbvMtm8GuIwWw8Wqu7G8Gz0WD/
qLpCUZg5j7TUKhPI3ZklPL7eVaOqwDJrPk8TuuuwS9/BHsc0+u0GWDS98mkt
+xp+DGCfNr3c3mbaB9ucOO7kqrRZnJ25DXL4nspQEg+I39g/JiS8o6c5Pb+q
iU9M/To1MSIjWQjg6ptONfZ2ZzolPG2MHtgDYx9ZVPV0ICJKLWBaKhT/nYHV
+RyExwNAt0IS+xCWTBwWcyLLAkOGmHVvH/kanP5ZeTLuGnphuh8I9ig2gkSt
iQ8OowApeo0kvcKyK27YifIghrTvGr4Tu67d5uWsfSTmokjSCCRI9JEsKRLq
zYp/kwgFEya+J6NyYBrCx6eNwutp/cUz/6AM0cU36MkXt6fMdKrfk8vO3Vfm
xjnD7nIg46/dlKToL/QMHYfJ2YHEl3nHpy0etvSd4GBVK/1AdM7PeOX2t7ol
CkqV8OIJTEnMSqU1vNjLchE5fH0RYdTXFSAKQMjld9dEJn0G5UbUCZ+mYYjB
1R9lSgAnBftg7CVRzNjkVoy+xgT1b48JeQXFe3TWrfkx2hF57Oz3ZsXV1x76
tJojqnEs6gldAjhmJBC2/aBeVyVtLnapF6mRyiyExysVaY/25sZhxLfNsTM8
I1j9wRxVPvumwqquD2JOzM75e1OUTwp2eaY3s/Q9HMsa3EDQ6ioUgXzNsFAw
n2/CYrTyH3GIxfoM+5FT6hyDnwjrGaYbeDmBhy/S57saE1UAYUbmg+auEdBA
nDuW+ECTWnQWzxDaO7SC3jsqnIcW0lKdRkdBaPHjmUu8AesaFEtVNAa/M/IA
VK4XK/gpIohZNAeHGIeQNtXrXLDDK6QzPoQkz4MeVIZttGExoVXLot2WkNVr
jVCDrUCLGVdPyWNnvPxSDCdGs5NumGo86ruoJKqtymuTSEdKXxEJ4Cc/BcW9
XQexoJMnLdO88Jgmag0RRoGyIrB7iei7PglhTvxOtDKW0/uhR4RX9rQxzPhW
JIo7Zqx1JVXeiI2I/tQFxsvGZwXPhgTKJT9w8fLcGArRYZlQ7fNAMsrxcDaC
Iratv0h3GROHXLTtzhi2as0K1b01zBbiQikw5BXt2i1vOX/0u5t78iPQxXJl
Cd46uV9H8ByWV1GwWUgbZfYuBVWbgueX4vTSfdpx4++/hUAPu+uWQDImb2Jz
HSQMXJo+a0koZtvCleLZxOQTsgcNXqBvDUV1Z42XabFg1vfF0tEzBo1Bmjpj
dyQi9ZK0Z+tAZbHaeamK7YA6J62w54AE/QaHl5EWp1rhLIj22FsdfYTxsLjx
CC2+Tovd+vjCNItne17iVy5s/P7M4h2zBuIBq5Qoonodpq7CV/l8c5XbUa4G
xlUKmycttHN1GnCK5LsfV8Qxj1jmiAx2XuK6BtgPnHTTKx4E0rmQZQwCwkW/
+/DvCE2N6lINh18IbxOVI+mg4EAUVKc0l5tYyhmERJFrb6LI+HHiM/TmiRua
hOuqnllN7qDt27BtEGSMqjnOwO26UQQr7rVxH0iBezZt13Ef5kEC2rYanLfl
oKeew1c7maHBQ/0Z62xn3GeFL48fTnl6Y2MDw6l406+fSFCyYq7X81W+i6WJ
vUjOqPEhRTuuswiCVzxldaf5ZDqkCUHgPKmFpBqSvtbvhcKwVlPD2r/b/GDV
2sTha4ynNOqGSqZGHqvZ0YsD/7ZaN6Lns0t+V7Hy9CGPfd33iyXCj8Ti2u1A
G/cww9H7OtZBpNlRK1/PR7I7aj/v4+8JGAlHFzEEk0bfiZTcfGUVk/Ynd/C5
1+w9WuCKPyzAn2TivX47/Jru4id8OO12XdiZsk6VsP517sjwNPAJRC8jLBDg
0HzpeRZwPw5dNfBRyeZisERHbyBMtCZYVgbWzOyfsHaLyKCTQtdeozollJjg
kQ/m6oPYIrYF/NFgc8L8r0biX7K1yCtMlQ4GF19sH8JJrR4veoaQN3YNYvGx
JWKC9cmKewKwPav9GYFdDfmvydBwAeajy365cw59MLUGg6Dv1OgXWOvRrT2d
asRWoXN+sbn2e/eicu4spuGTQhC1/LngVwdlzeqstK7/4yW4tRrV929QdO01
s9r7NnWSDwN1orPy5/YeZtVPXojmpCt6EVyrmmMUFU8rHtX0YIViCvE9jkBb
Twf+86KId63c5MJddSA9+cjoRx3yATHgLH72he0OMZlXsYv9GGgTblK7qy0o
qTEVRdYmw9MMj72TBebZspR3yW+Pg6IkifTu75Ut4Auv0GC7Y9/bpVAOp2Md
JxUli0ll89X9/whL8rffbtQjGg+5IRrx2NLyVIF5wR/lMvP+es6iyFresUMh
0ngnX97XiVJ4LOIu6UAtGASAF9hkgyO7ZTdG/rmaWEBsXQuZFNoIAOypPyMe
gGuoU+eWTFbW9+9y2zjkJJvnyCiZLIT4qOjcZVLoWYwNC/eVRPKAabU1/vRs
SeeSjepxeReAd3dxP6Fu5MsU1gWxyzKTpvnNmIMuJDrKHRSM97j9viyODsv+
QQUTQQH9OxN8wuKU5HpduSSKLhNA2EeZfqbIy2i8NzjqnGdxBRlX5xuWaE5B
lFRZfscqsEGIK77pK3PWaZJ2nlN1YQbCzK9m8oFocgDlOJsJO347PlqOXBwN
mK7AywWBj50YBT5aV0tETO2CqWeyPb95cjOObuTQnDZyEd9KxeODWlZiP05b
QBy1YZyMis1lkXZQPUV7OhukfL9Z3tN6ZW7iuktMO6iau0U5dxeFrF7Wi0co
U3ul0YrH7/gyDQawLwMF7cMF5LavQHTwM4HVf7HNT3O+rgbjqvYJ90buTwL0
nEaLRxVv+o/Z5VS2dqYvro0Z3UgjUjDsxiZOJQQwjbGRloT35/uESxOokEDq
/382Dg92NZVzFP2tg8/mHaI+O1Nc+F0eBoJF5Y5wqZIXGF/CQgupTAL4Hmhe
h8sLSKF3neMx1SfnzEbs6KcSzGWSOqOBSmpfpczCDn0uw+mzlqcGTIycCE09
hi9ScDriTaJpB01bYERUtwoWF4NWlVRIUiBR72dO3Zk2SNBm4aLM0H+FDX8c
aeiwFMbg25FFYZSEEA+B+yLWZB2gC/+UNvEJhnYc49Ftwuec3ZcM8WxxY3ZC
1MNZcylXPpvXsIAlWsH2ZGmiF6AnO86qfxD+rjMzObmMyg9nE0K79bXuwaba
qU82VrjeBHqpJodWpr+1eo7N3AQBUL8yKNbQ7yp+Vpsboxab+NOEhph1ltVO
JPSBpLkVPIICm4XzcxQ5MLbNrUssP9onrR5PgLeI8QVsNaxyiqNl8nCbhj9E
jMoODJ+k1my/2PwZ7J9A6UIFIBlrU8QpDJ1wjrn2UHPzssrsSzPadVz0zDTq
NegaQwXjGNXwzR1gj8IKz2DtLZj7ol5jUn2x+QCgTyCsEszVt0CkwcYEMgZ/
xRLCDFDGRES5Gzbf+lvoTLkI+qHDtdmtoEjhzbw/m4qU/bp9qxILrpARrbI7
v8ca1KVWq/OBboFE9hEhsnopzRNVFyJobu66AaoB1/L9Usj2T95TRFaFYAhJ
o/NvP21gCr1Z4zH5jY8A5t5s/V0SfT9+m/+auhAK/cJpXUhDK493rzyGXcY8
/+Z2DtOUqXvDvHZsBEZpAK7quwJHN1u3PdKIPW4zsvl7mOGzBUjOUKcGNoZE
hXowmBMa23ViKqcoinma7xmCSlMJDFUB+OVE67xevKe0LgFeE4avZC60/tQg
yXjtE4VdfXq/cmxnyOR9GGkqfCRopiu0FTzGyYLOPOKaume2nz+PKxnh+b8O
ZvyNwCEkC3ZsE7du3usp5SJasP0nAiLrJoftxvVJcFPftoIc6lMxU5YRhTNx
HM6fuxfVokvPzqSWk+VhudUv1LKgJcGO+dxJUmzl7H7kEMTHjclowyEjKFXj
nXGNo53MoHYvgRXAxmZJfwB4xbDuQ5+XzXI0nBKPXy8mT3TsBEmjN5ckfmwS
hngu7Ps1jr9BLWNg9A5Sw06ftqwdL7blU0rMIWqO58GzkzW1XGE9HgkLMz98
T10apJrFsYaPzpesw/Ee+2lVdvcCYwly2IVeMBS138D44CjHa3s6EEd4mSy9
8so0Tx5ehBUjc+yfo8OLrp4x+DG0a5mp5UkFUfWXkX/wzGjsjXhwNGspXuEb
G5ZagWXE7KJD3cGptUrziIlI2OY0cf0OcHias6I1R763aZOCPFNp1b9TzFJM
Nt+6ZSfnWhRkVu2wHxGIKdDYQklRkHJbn2zVhAzExmoxXFVOEpHoKYBVYCdX
HBHwCsTsB6i88rAVIK0ahOgVRAUYMfyNJ9kUQFK+7JNZqc+TwRxx5mfnEhZ+
Z8AzSJA4qEsHprlo5ZiWsHRR3pwYlyFsH0MMkxq974xIZPDABtwXzyZIYdXz
sukmlk4CLVZameE7uECWprOtLLPz4UxVTlAeoZR+rvX+mipNIh++0dRD8S3+
v7X4gFFxUGsfkozIiaJyHvgbVgpGrGjc184VgmQa/BkpKIypOOYgp+iXv2FL
cQrFZZUAz2au29V8scnVFligCF8VpyZKQ9ZsVMmd6cjetp5LSO5W6nXdZ9jw
dvPoAo27IwY2FSe2ePKa4IbFiznDab8Fy/z/MxHs9iJzFC0/ZbqNhJuapaG0
ekc/bNpB9R0rEl1QdktFZsK6V2M6IVe+pTrwJ44Bvs1kPVZqBuDNFOSGiTVX
5txX1C+6J17rAS45JTjYfR/KGAoHMSkr2s5Lo1EIv8CJWR/XEijts+rW+Ax7
GXYl/PMe4SHbmsqM4H+3h7fvArPQVGEd7y/hvc4HVf/iutN4lzkuWPTkppHk
/MWZjUEeIFljahqFnOhTic3innmTgxpmGSyu+ZxV8iFREtGiqb1GgvyJ4j9l
AobtunKchbSMli2+Rt2H5ZdF+yFLOsbcsWylCD6BcSWqovUPwhsMC8BmwjNE
YsP3HyxTSp7WtAyNbKCftw7w0CPhVeteui5uv6bEhYVI7W4gZmPE57rhGCdD
N2GJdh036MaflD8SCGq56hoOLRwJJCfuwpX1UVLsJiZUVNLwEJcDzIN4cFMq
UZeCEsNJFHyKmXW9OtT2J9zBuqXydAreVP/rbQZ/0Sr1j2EKHMyOljxorf5T
WTwePOqaHjqhz7U1F5hGX0DoI7A8PsWMmhIImwSLMYJ+f+3/bEUT7MCQzKbV
GgG0t3zpm3HQECnmr3FDW7YrTcP3WfZfu7g/n1GNuxZc8Y9iRYcKtVAvxRha
u6PXo0x8+cNALXoCI7Bfue7xhx57aYmXZXGc6nDwarN5xDZhHa0dTsPEJgmx
93qfa7nk5sjpWdi/ktMqcZzPuXcTZ+zaCkkxfEbjzxSGSIZFKlZ/dnmuV/Eb
eA24Uw7ekW4H2a/HKIRWMvEPbN074n8KbQary9Se7fQ8r1iSZWX+1XKj1sgw
y0XsPlxWpbLsZ6JIsjz25hB8vpMcPyIcYBqfBJX1XmA4vSkZ0UrLSlSo9wNF
C/9+NRwUOHmk7plWJd3sm251NjgFX2WZ0WxbvNDPKQ6CPre5gEtRQVZ+2NlE
kmstbYFZQ1f3W7Xm7i/Da6hnQnuUSiQ/QaNWPtTT9U2XDid9W7qX84nBaGQN
IG6KDTDufyhggOl1zPUolHNkO03+Pim491KdsAdqnON8klUFs8AaEHVwhJXt
7DUsT7WKy7Hrf1UiWrNYekpbm7JkB5ShG5aQ78QgWJA1LSvrTW+l3OlvLFc2
lgTn7B2ESXLkRo+Bk7efJZeD8yVv5bO9FSzWYuQE4l24oDFQkyfvFA6RvYqm
P71kGevYGx/IrxGCSbxtwgvD3PPYu1Xbft0w5PukiK7meoRx1tV1roOHPsC5
RShIdpCbkx0j0g0vTZETQy8l+bbQQRmAp6ezKw/8fdB+/3S5QdikqniLh7SC
6eT0P5YmK5MVsb1/j2jSymL0OOuZNv5OdkOR7USOtfsg6/AVY6axIRHftScv
y1Y+MJf0gJD1nV+v0U8Eg3fBKiqXn5BZZmwZZy0mu+C6H8+IRg2dCU3RbZ3m
SJdh79ikiPhUb93KfkwKKnrI15RsvKKftthj+UquxEJ26TKlLp7U2PT5iFKY
IKvKYS++qspMlW0dAkvVR070fCP/anidk98AK4AEo5O5onj9LQfk39/FQxui
0EFNqC0A7TlOqP43MubNjEwEBZpYNI/+s6a2ghkLo02uAi14KLPQKUWFPNgr
BKP/QdrK/V2+ZhdQ7Px42KIbe0Wt0Ea+IoSCWq7t1O8zP/KX9J2amBx5GS9c
uftCO//F8ByAkVC1EX1F7WDH2qAeKsJHZA4uCES6T+y/jGQ/CvjZdQQn2rCz
iI8mMzDDaI+9OXc20NV47pNigASiQWUnziXy7NiDv9pLxgGW79OzXfQQcOe0
+IdQt1RJN8ZAFfn0hB13qAvp1Ys4zHjtt+sRIgu33iYcN5KD6b/AqCMixUC7
IpMU4og5pDpUXyZ5j4Ml7maVQzQqmri3K7/soey6EM3Nq6/xWsmjc6/jWGYb
kGxsBp3ywHvJz0LGGduol70EeJRCbMxt6HdsT12iBIOjIAsocP3UCAl+Nas/
R2+HszDWDC+ZnnmndpXDGPYDRvyWvf5YlPelXu8Yb1SJsrL0nJFJlrk8QenY
flcyKuw/LVXl02ZTwaJwPdWkkxD2brhjLl52q54MwXdZc8PTbrNoBJMhIytS
6kkxRGXuxQssDAWoG4nHrSlSuLzd3e98XOYaTjBq7y1bOiAJhOwPgHfQBYoi
W9/kjhgziesYY9iAbRiX17XXXMUTE25ZTKw3JtCXiP4exa07RSpLolVo9K3M
m5HWBRn59zErazPDMcfSY+XFCwopywVmTdw2UOkpYmTeetXdTAIf6yHHDQHB
wTLE+4dwP7lA8CSE2ATa846RAWzdZiAuzSA1Ke60vQwU0TAl1PGpjLjPZvVa
AgN9KWmkOXrzpnXN89sNKlB6xSsiTcDSXZ9u9jiYN73jnUXm5SGwnHPIW7Rc
BeE8wviti7TkEMSsZUoX38pfqNMT0+zLi51I9gGT6c6scoRai0rGLGbPDkap
///+UZWTRSaS8glNx3EgFeiTPFmDPCXhMVDs6EbkirRYfXiT6aHI0k0Q2Ps6
H3/poj0M9MHARDXnrZ6e/mxP9/6OuclLFajxDjeOtJIIivFPkq4xS4dUWBMj
Ycc2UjXq4TnP5hcTWdaVh41jdseVAl4GXeASxKNpEZbL3ZAYovtiJqa1m7R5
mzMsT2N8t+DNIqYcDL45oM3R2WstV0ziR9sisNmArUJMvOz19OZWuUPMQM8Q
J4mfGV2BzeyO857qOMp7nmUU16jXq5eQ0N97p29dqcttyE7mP7iS3vexsDQE
i98+qmiJkys/1gg4qbdvJNCQj2OWjsNbZoK1VadIuvbjLRzUmgPENKbFetbd
nnSm40hlCHJHrTwa54AcYwBwkfmnWZ7IscRNB2K1HEXs26dO12uONVEeNEiW
ThCMeD5cooH6nd+ROVaqTYAC3/399LtvVcT4xxdGeFlrHyvnll9R1pD9KUYC
bxITVjEbzD+hYxOmaw42fsms0MJdqk5URcMo21wljUY/dHITL568v+Wy4ItA
w7paRZDbXy1dD98eIh/hcJFhJEMRZYgBZXevfvnykeD/lHTNhU0qcV9stwzN
PZI5jFUCyJHTKN98+jsO6eV4J6bxcuejcJPpVcBFAul2II1NlESwLiAT6i+F
zRBJx4TFq4kH6DvIq3AJrZe1bThZLYM1uLXHnXnhuREW+Bqh/3HD8ZFYvPRH
P9ZZfIKggzC20NNUw/kLRC6bFjbK+3re5YGk5ovRIcVGF5ODSqlFGtDuPgSy
hkWjD4wSApem7R3U8dRfKQ4uvxzZjmpYl/KmTa4XB7gzqthAZ3ym18znO2IN
wDC3zBdmauKKOK77CwzFKdQzHKnzXFf2WACwYbFjeESY/LSHe9o+/aZHC5gT
96VI1/ntMYDGvjSC9AjFymfzNJU52LKGWdYwpjoXFUfujD8hamoN/qwUZN75
aJjdizHX0pw7hhJBb7SoZ1+Cxm82E2PBzcdHV2vi/aXPAmaKwthBMRDIoR5v
I+/yacTLMfmyx9S4tOwY6eVe1k3MWqA2ypJl68G/Q75tBzLSygud9GJX4aBc
gIzcRD0phFmwsCvBXKJduuxw4bBJcbwpVBAnbqyAINW4I/N1PKbyu/sU17ua
+ziaTvqhDNMzpAgGT4FqcaNfCs94kjUPlGWJg91YaFspe+OCdlVQwCN4AsnF
an5LhjU3Po9gNc5mqLTDIWSOZ12Mx45UzB1x7WyUllhpm9TVUrEYGCs560XQ
mT5eAo7xDxzb/+bX99bKGOZZfsbZ5wXGjV4ik83G+vE1Zyz4svgp1V/2+oob
/aPYOjNvpzijT8hsPMRAFfm8UZTk8sppqLj8kBrswZdOYt93SZ7Ab6PiThCF
JRAlgJPBRybKcTVy50iqVhYmMfuANfjc44KCfjLmR2pxj+O+mDa8Gf2ieg0p
nmIygmDfAla601UljBtgWpZPjfpnaGQXJSF43I+NJuPjnJvgU7i0gCikGWlo
+JF4bbx+4rrsc1n4LQBD259bdsBkT0/n9HXK04TSF/D9pnfhPnF4yhWVTC5K
xV6pex9S+3Hm2O/NT/U+r+A/S7Fskdv3BTE7uufXzZLjefta69st7eLf5UWJ
nbR/RvGkdNBHGo1ZrfBwLwDwUbDsSunrhBwo0NyWuC4gm9jbf2HPi8bDqovt
mX8hmXUnJ+LbuKYqzbomztGP4ZePdp/XVehrTRjOdKQqCGJrJOndTDL7F5XG
DjCEV7qSToOLsEAZfYrim8n/GrgsA0vn3K+3riwIDBfh7cDIYfiil4/7wijY
9dDhcZPDBtu1fQUPuHomFol0rywp+2flqG5K3JNHKVucHossenLdf/NaTuol
HQMmW6ztSjef8UNyAnMgdaI2AGKYxTzloMN2DfAOkrS43D0+y0klQ+m7S8nF
J0m7gVWvI6eB9RvfbDYpGuhB5yfqLaS3lFvY+IxsddNSVlwSz9lg/pBzfQiT
oDQjOZRiCsNE9DjUn0YPrHKTJsQURq00zZYf+e6V+O3es45mJG3CKdDvcnsa
Hoj/0ZNYesYu2yP/s4tm/W/StbZnoBsJaIBYaFvujH5fwFmnB+yF0WE4Kwje
YJyLROd7ZkJOF/1kblsNmo20w2fmXvsHcUukq2qIpt5GmXP9XQQSRok0yt5a
5gZlrZzZ4OADJK5w1sOE0YTMVdRyB1Va4Qope0XlhGyWItEDHZoyFH7NAerj
g4o8irzgPrWtVAjGcv39PkbnyZZmbKzIxr+ZEivlSdryyzKCtrKZdGopNbsm
L9D/Dw8CJ8Vqj1ULfMBCKRQEcRtoXMmNTub+32D7TNhXMkciEY6hmWGJQfy5
sH6gu78+lGQP/Uz349TzNGH+wDMYkl4AxCSF1rewKeky+4/r938r1V9VZGrd
Tm7fK5/4oKsvlv8XEWH1ptENiZySuEbnTUsyUOr12DLxU6xwhGMOo+3vrpnC
aoGwInuafbsOxUCahjCMkeuaNoU/Fw4A5FAUrCtnLfVmjUODCzRZ9bdiQRlp
UcOk11zBEbCCrYCYK8jGGhoZoJs/WLFDNqho+WMpNqbx+x/1m7ENV4+dwy7A
r19wvvGl2nJVnNjoSPht3AMN7Jw5BXfvBOFadyYLUc+6NSpWN+yYhuEbZa0r
7+jvrcB25R1h6sJZ+wBpsFCqmG/pPNClEr8EMh70GFq04TViA9xwlMwuroyk
A65TsR2qMOTdaZ/jSgw/+JU6XVkr8cSFUx8OnZyVwMGkkf+dhCbNXzTGDghh
NnEb5OwJgOoCpDw4RSsVjMp1NNGa8Au5GW4/ctglMEbwRxCDVC2bNrQw3xdc
V4Ll9oxOYjc7L8hAMESd0taH0ezd+A6cAa1sMYbmYEApWT2rQm8NUOHBHvbn
U0y0qww6TanWzEN93ozy65IqMHrRlIFTjOE5KXqpqswpck9a/wQBOpnDgKWX
NRlRfXuoHbq/65kaM21IH+1M2mpd2g71y5u2xn2epKGD6EJ4tP8Kzo4yVQP1
nlam+YCsZvks2XjfzvvGLmmyiUm40DiaHZqYdTAqAZIFuq+jpQd8medEw5fi
T6JAf6RZqgmY+5L3cBqebbXbgG2drHCd6aJ2cjl44GQHff5nZilSMGFiL1aH
bR57KHZOyWnQAqxLQb++MbX638BrIsgsrpyrqyMnaHAHQmJOrvy4ENxdqJFl
OsEqY8zF51Rn77su/Xihpm0ZE/UW7A+MMjk/WLp+X8JsE6ng6K+OYCqRssRj
8gYJDtGFvDXgGpX3TSaChlWMVluqvIC/0XgVbcmn5C/kWwlAAxf/qQCCyWx9
bx/XJIZAIOnp7DbEwYhS+rfE5ZR2KTYkFqQAV7Aukom8J4Ac1aNl567zmtiR
FHLLxMI9o/Gkc6+fZoHB+RzqaVY1Ljosly3n06+8DkEYW93g/2qUvXhn/nV0
JWaGS/RIEsCk2AnplYt/r+/lOKPw77Hv7CSZ8VlBohLbWQv2zUy8QyobQvrp
M/6Jbmb7kjpmUNDHfNzMMVl6SLYMp+Eqe1lX02mRRP77TUIzcyipNPAZGh4E
lyrpoyO8212k44hBe56xAt4JMCIEaBrEN+KKkfzBunyH5nYJlakSF95junZF
uYowVl+1WYNX2u1itdYpKb4WDoI6XnJuGJToTHcxiUQ/jGeKD6P1xcDWuHbH
5K0Sw61dm7Tq2KRnvS8ngCaquVMvV+k1/uMIZkRT7T7CWKzEvZxc1BqNf8HN
cQskMckPT7e2GkIr6JzLKgrz9c0ogA7Hm3Ef/l8szsZZXeT5Pj3hV9LqT5r6
WlhYY7Fb8/0AlpyyqKcgOV/5wmy+NzBc1BWJiHAcVj2p+EU1wju4V4U4xist
DRlXWAO6QsxDYauT/Fyq4zd5YeQxGWoHtiybgBcmYugW2BWGli5thFQsffD2
jnoDmHIszSWjehHrtwXWeR2UFMVN4zdT7gA6tiH89mwuZ6ry/iEJE0eyCwIE
MgS+L895OwLf5BrI0ZR3fQaQIqkYcV5omfhzqi0xCrD527SIdEaL8HKTVVaw
Z5lZBRhNn9QBXsjMnijUFiub3WJVLaoYh7gfqkHEKwghB2pT9KynNnZH74EL
PI0pF7MDKmvGsYBfey4g8qfY8mXD709Vi24yZWiAI9HkVXXDvttmtVFLsYsb
Vze48kbua8qNlguhi7Oy4HOcGrOtV6PpJnCR2ve1yy5xAaooGQ65w4Ep6O87
nsC19LTQwrpzHX4kjkg7kGN8yfXHMhRkEPAyfD/KHWkx+q4BHU6iQ8jsCv6G
5uT56uaA/pV3dmfWydppZcmyfJ8ILCykfiAdVoPwGQYxeK6ybPaB1e2Q12rG
lY7gH//tMrsmwuaH+qA1H4LrDCqAcVLLfFTDhZ5N+14vOilUUf35BzfPwJ/u
mHE4zb3kaQgJuPpSmvhBkWvB2ftNJvCzP6AsXqIhO0qR81lhEviVDp9Gy8NQ
lEMZbjdLqSbH3hsaqZ+SILJr+V3zmdoVz60GccGOVVRFgWiFxBNZzdzCuj9q
qlMgWNeTiXD53/ksFtxlCobRe+hdMtI9dr2d5YsPO/a1Yf5g/J91VQIsAKMV
5ABXJi+C0kb2atwfjY2WHv/r+wHM6ZWrOzIKwaN2bWkCaqPsc7nHjv/kkMFh
cO8gWUydp4Sq/Mj3Jv13BoDWVhzEec0aHPMWUYQZQIrof/5eOdlk1WAXOBSG
726XeZ4bYUK0KEEAEO3v0AAqwWycoPDLqpuJgIM+iYZI76fWwVXm1iusNUWH
41aKhUrylmZojPZkvKXCe+es61BoffNXSNI/mQvJnr7dpxjMH/lGsgU/zvFO
eq1kBkOJNrbmayQjXO7tYOfeCP7zfB40BHaVu3dwTG85iT0FND3OAoAYgNoZ
xzTr5e+OHzqOWbJrD1X1a6RZi4mAFoTyGguX2zNBp7srXIzC+bEPs+6Ar7Q1
JTiqPlrbnjo/lrFF6l1Nj19tq6pzjJRz3oATgn8U0lcG4eAKLEHLYGl3VhmE
eg9Fw0tJdAxhLodmhQr51JMdJYtZWjDiIWp36GPapcQVtbjYQVpiiOcz4vH5
qLSm8moXCbT6SuCnJFuXLYLlwm+onFrmxCp7zxrw6KhKxC1Ca+ILpkXkpxgW
VN3yayJVoSmj7ZDQpw3S+h7Fmx3+insr7SDToMvoq+WfOYnUzoH9nToq3C1E
kjochcwhzM4a+p4OH42g36qlB3uQ2tFhJhFw/HRnX6IX0ehJbvN4Gk5JGdtr
sg5+mv4quVRGjpanHyPZhclcaVWk3P9crLdnyDwIsLA2MUWfq0NyUry5XCYB
AHWYgCEM1yrK3nLh6zhMS/NUxPWPiD506hSYjpEFzE4Ir9kaPVyyowB3E/uB
veg5biUbPogzkx+rkLCdhaJErUmp3GfrymsUezA/W8hZftCgPyI1SBqbFj0v
JVu1hpbRoLFZtO0O7n7UgB5gm8zZ2cQCsPfXM4ob3tib/buQ/eSuVHKY6I3t
OUKRgchV/oxRo7UTIWdQ3D/OpE2SGAnDZEWDl7pAvz4Dp7QigOVJ+306LEi+
XHbo1arwSZNR1ODL1GuGFla7lN7hTcl9KLRDV2wSbWgVwlDjZt7cUBtNXjQ+
5DRgV4PlBfFUHtEj6qJYQNecnJTG9zz0t1pCE8tWiWP3fohJicxc4ORh4W6M
pj8J9Ta6JoP6nv97G+KyWObmaFEvF74sG0UKJPfJpNsUpH19XZxYyCuDpcLM
jtWVd602DMb5ZmhjX/GwwcjiYl7gG6Fy9VauCTFUlfMOZN5+AjsnpfaPBIp/
KvHEiTEO7Hj3YesdckO5FJizkKrhazmViS2y0qKN5LSPWzdk2vLzoIEpib2C
9/HJu/gqCOQ9Dr9kfQ0FUxsW9RxIlR9WPWv2KxK55AZcIgPK4ocKUeA7iwqg
u1DoKxAUNaMCwj7LSFUzQuOBp+5dC8luWyVnAHARfmGjrxWkO4PEaiw1Y9pC
UUolj/SkiXqNZjFwNtSNo2cYAvf+CfdR4OdnLKxM6wrG8b6knu33h/5wzmW2
W4oDsjOtx373PeIKZmwNRHOdA5MKBGtAa3xe+vTPH4Aw2ldwJ7EbdN0ILtOy
TY1yQzxP00il3z7dhHOLfPsxY2FjWaQk9pbvHQXapfzjnJzpB9KO+q11DTOt
Uk0FFUQC5j/rp67VrF3+6fSa65ItGFLFjC3I7Y0A6egXzTQzPz0kxzYHwZ/3
+Q3sSxwsfWg8TYD7zPcRLBwUXs3D/WQB4pKKVYbXvnkQ0YnzUijemx7zZ+PW
qs8M7bf9GVWxaul74BmBQdy9n+0rnRPNRSyVDxNhP7xKZ3Thep+d46hveu/B
BcnyAotdgzWos0gIyTjAYrBunWZHgEBGj2eJLSi9jF0GvidQg7dmglS6v0nE
LYpMTbhiSFjU9K8EFRFaTh6Yy/PNA/pi54RttdLW7Ks0fpX8PKnrBjA7hQvE
D/Fwtux1ZmmHsyeF7zeTA7eFWLGV0uZcpUanmqpd6IuAcft5SVglGsH8cfr9
OC+xjlU0wasyVVQN/nVjJGOqeHl6i7C/yE0ZtmoGszOXqyq81UIvV0A3p2L0
w99hZ/sR2qvA1QnMoAKwJ0mocn4j99Veh/gfl1eLYS63Xy03LxiIRllr2ntH
4HxaFLuVJXSCpHIB/vm7zginCWOkW3cW7vayUsYKhHqL8l0KaysAaNBo5ik3
AJdnwjDcQTjIWpd6s3+6RRN5hTFNgXZS9mzyZMcsLTT8JPQz2y93bripQE1s
gkvlPafsYyL42k6XzXzL/xZJxgdiqIf6V+uGTVU+Mk4LSnD0DO4t6qV0XvI3
e51uygFtUYL4CkL7utXynP1hY50dTJbR4eyl+dreKRF1CcuOyGhbQVbGitt+
qGn3wyIqz2RbDDfu6veLD6X428I4aQy7hIQB9WYqUwpr7yWJ4tpx/obVrLAA
Q2rAPr0xN6twxBqGk0F2/oTQ50iv2iL7Og8DmK/gS88F1m2XoLPQvQba8VKX
W8OKU0uNp1Uia8EP19ZKx7vkvjtjlQdBHqTaT7kTD3hBHX74vfOykY4ApScO
gX4HXtPbdAKq5BaMl4x8Nwl/fD3EpSavC8jKoN9ugUfczjSMEXycHW5+9tet
1+hjLkSqcofPEvz/tpzlBZ/jb2UwOecgoBMGuOGG+8HW9eWQI8nm0fKCvnKx
AagteinF2of24/4R+mWA80M5EqLzM2rEedViAcXHYgWnEGgJMnooMiGABs5B
M3CQXpv9CQXCQjmbPBfaxTo3icGtiT9wOyXf4t/F/4krPG7KNFCQgKr/pp5v
g4zlFt5qaw9/AjRwJPf/3cbZbEzlR1o6ya0WGVKBJSSiS+S7lyGha2lUAQJz
+sTqYVNKz9ki251Sfo/vQw/1wYH5ix4qHv1ed25KJ4HrO2XEMT/3PirHXZuo
6vJw2QTqAgom+WYOU3SvTFA4/AI2NhbVdGZoLEYbV0UNC6ASYHAdK02/HuKI
pIHN0icCNoUqorlR1tOlDkAu53eZixsJ5Fypr9ihFCuER7HTFl9EbagNasAH
9Z8SGeHNuKCeHYGyUHaJIVpMTx1/HTZiyxa3GB+Vi/PimZG2huCY4F4MXB3T
5WwU4Et3vS8O5i0fYJ53PyoLCORbYC+7APxYrDLSmobtM4ZjFXFBZz8R3N2V
OAPNbaog9vEQ3i1OIIYaXnZ7cjQSQ1VD9i7p2cmIsD1h+th1zwN1xS/looZf
tbBJF+zeInefEaLEl9QjbqnMGkUwSFqKKpClQRLgVWbATtxg5vSsW0NhQ2pP
8JFNoZzgtaFocEu3vnQLs66kNgHoUimxnxa3JF6fdV5H784HFa41AEGUuOhq
EdVASDY+dGT7EcZTtQAvkRXvXIUBR4cE6EFZ/mVT9BbuRSTXVTiOHWuGJ1WJ
ISkvTKVdgqwm2wLgnVtrjEc9Ntukcd1Apb39voQFu9WvP4j/RYWA4Z8vMPM5
NpqnC1VbDsiZSR1bcfcd4ybY0RBnExFEXTQD6BVniejKWIHScTR1KG4jonc1
JV/Ffqhf1W6Ctg66NxIv5tzicdXKUwu4QahyERYoSj1XH5piAb1JlaEyJUtP
91lZba3xgwvvINOUEGY62P8Hz2oAATMkJAjEtN+s18j4A+5aufllG5ydrqpZ
ArH733b+U2IK9YkV+2XgOB1XSU4p3ab3KOl/pzVfJoMF9kDCXmlhXep9AiPw
pfvHNwen9TZgj5I/vmBFPyBRad/4jh0IruBiMu5fLP+zrIT7wAbIiL+6MSo1
NDrUllggyoogjcekQ66DnRKh02lKRTryLm1HCw8wpar3X07zqACxN5Qz6u6f
6MLaX+zvB/RfRrOFZTKn6GNJCpAqnoixFIl3DFAbNNpiFn5RWlMjKcD1uI2H
70zrO6b5b0Utr988n/47C+PpjaWtbVMm3XhxpkWGrJAavxteglFoqJ7vkYDc
wI0tKTrc8KIdiY789slrIol0JfjrnghM+vcNxeFLoL91W/jY353OhYs6xLxk
pThQXdppprkuMBwLba4E2l7h2kA5YE5mcLYJwP3ZBFRUGzZRDOtzHzjtluVn
IzMALb/cvj7e/hV/UFOQdN0j50hLBkLQPn516iLK1HNXQ4VGo2LY8V1N0S+S
3UBx5SX2dZQHg/m3Uuosc1iAmOgpGv2K/gIFhBzhFYTz+HOSy7/D+hp0j+zu
ef4anOXwKV5/hlrPuX5X/y3EFgSNYE6hWo1+ihvhWf2CyQZq0gU8SlozPBBI
3zZtamWLNTXMRNb5cTc3JOPfrFT6aKIB9HQ4a+cx5snYKVYCUf9i9cI/IXz3
uPO3BmrV/J5/fKn+Y32l5MO5oHAZ2OTOSIfTwwjIGPKU4kciZiU4uFVOZ4Qq
Aim/jAmLyvRCw3eoSYrjp4eE6XBFhHHzdLv9x8gd4GZOWJhSdULbkGP7wsj0
4B1MiS/16KMeaYlPK4419dBU8DoLvxpohVC+39y2fsQtC7SqFrWul2YoAuiw
U/RZ6SV2jJo0qkV0BvjtHEDPC3E1W+juEHBo6NcU4Ov0VFps09Zl4zY6Z+VW
uwel749uTgEpF8g7Kix/1bPkmsxHih7kx6Efm1TMhTseXwOEOGDeOSw7xMgS
8y9GxrA51GIBpp1rCkwlAIyNNyZOcJu3cK3DWaaajOWh+66rDCaOUH6j1uh2
+QUmwcrYlEHoejdwwqifrzcTIe5JoRMuuvH+IfbFpzTuHEOcPQoO+j9GANPT
/Kgf95s40vTCLSO1huCes0065QczCkQG15oZKv/Mfkgt44p58WpxlMn7RIj0
CZBi8W6DTT0wdpcULPfyqIarAEKJHCm9lF2KMu/A62wiP5J8dPbk/KGPqmal
UaA38J3QtnCJt/oI7oFkfS05R+/UO7LCapCFofef9NMKf2LB4a2baQbs+KBE
Fd3yh9yoggvz/yrf6fgGUSM8W3/fl2mw2pVCTU6vzgsjIbNnIIR7Wj0U2CpX
81Y2Aa1CB608k5M8ooexgUvsny3niKn9BBdIaim24+Z1ahspwToKRe1P/fxW
pqVP1Y6sRqAjT31FkhEsp6NmkF/JaQHsLBk7bAgIbBVK2KcP5Z7ZDvHPxAWC
Z9qjVLHJduZnPfPcGYLeUnwBWrO5MK1zReSmwq41eH0PTbHT5GVSFCTX6Fhv
ZD68lG/7mM/crYSgq1bIZx3s7eBvY/MVcQc7ae/uRir+gQOXQW5u6WsqLlyu
IF7aIoXYf7yGuBb4wZY3f3jhP8j5Vu0ODafP2qEpJPTD3D7adqFxG9NHZ6Ek
AkkiDaQkadcgCp4RAsdwQWfBlTY10RMbA472hJqaTlJg6Y3tLiC6Anpi9cyY
QxN87IByl4UTerxsaxHcTGlxMGq7r2D+Z/Kd/BXEfsuzymCDJAXr/9/GyzmD
GYDry0IevsgDXRnYAyE37gbkX9Ie8+2J2XlNwyvizfgGZRWiRbUHNCSBwpA5
OjIqT1rsY/Sclt3Ufexhn4rkdt80Hh6dO2wg3Dk2eZ6y+YLjIPm+mSquDOqJ
TrbgTdo+lT0j+/usNLm5oNFVxy8ZcFqW1ll106BC5kdBkkJEWU2SWUJrN1Rp
up3QXA2BaWGZ0wn7SHkZ9Dq/rxYUlwXXD4Y4VMEAYx7R+9n9+L8WNt/LtDeT
Ai+9UEPYJBdy0/UsNbTmdM3q9GV1yLgvnnfnMUYS1uMZxc7sdiYkNfg9d0ee
fdOqasCpnLINu/9r+zsLzUo/xyRG2uba7LEdxZQI/LYXNrycz6UkZC3dCV1w
y8FWmr4U2HpxNT93moSHvhZGJPzC13HpWjmDG8fGjMD8hJbeMKWKxVClEVHz
reWWlqzPcr4Zzyz/Tzqq8SG8T2YnHYzeJkxi+twA5lsLMk1TgxFtFEsC0Xn0
Jh14XBE5jjVd2bHUuOkAhUTOOyAjuAxHWqQzDUnJzSlQ6Ja4WaOcizqFdnvz
VSQrSkxR98rQ3wPgrsU2V6StbJKaS0SZfTOdJbbER/gPtxapAcxhtTxFVVS1
+gLgMaCQyT6AyC/suv0gf4qY8eNFdu7w4l4WYjr2/8AT9o6FenAbIkmP4b97
nhCz0lBvFgeBWuGbxRXOaWRZdU/fAXFq+ao27X0SEQ/WRFJPA4ckyLP8jZZk
iIHHPUZ4g6EqUyZwfZVpFOw7Z8HD7FkkJSUgFmQH9yM8FeAvQjn8TFMBctl5
pJ+jIzbHe89BXJH00zIeLApZzhj16d619dFj/tTl1q5BQvHVXtBQloDkSWA9
pP+2uXIO4urWz5ExvXPz7da678F8QJY+GY3ZaeM5CxYr+zK+f+vo4+kIRN06
0ZCx1i8q16irBStoIXz2TsZjQmj28FOsEyMED7NwqL+JB6JjF00BQtxlrlSD
bNanLb0i9aH3DT7ZkegUDE3S3jK4jzCUPo09/uT68GiDNnnJl89E77Bze6Vz
KuJWz22RzZWg03PoRfHOb6JOdOlF9iAXcltzOc2e0eSmr3YBBg8hBFrl2SuM
ktMkrFrcMwslwtjuE4w5GSaougjZsp811m6ZNBhNjpxLrTYQ048lVt2MXffB
l+00joMudblhuQ7WtjlbSsgDg0fnLUdpmSigwsQ4Nd+Xt+9jfeSA7Np3wBT2
0yvykIXCFSuqHH/z/IxTXkasd+bWobzWWn7ANmMHHCQkJ2KC6+L4bfbT9icS
sW90YsBAMDsHYDoEyrFokwP3Lfrivf51CZkX7025xNIAcryDL7XuManeb4ap
+ddxMg7TG14Tpwn1efgOaEPlQxK8zJd+K0T1gexy8vz2zOHpAXp45lsSoop8
tUh1SmlbzQFHXcjIBde0UirPsTsJ+H1rqbFY5cOeBul6Wi4K/XUuuR/2wFeH
mOoDPFyXaR+28TqYzWJVzepxH+oxVGcKtEnqJaTzqwgciTpmzXDB4jHdB0tS
B5hnPp5uxv2HNPu9Z9rfIKGKzU1PiB1PMcJ+9+QYZPGRXmU1p+FH7m3pXSGJ
jdRvZ/bxIBPx69Bv4uFLGvzXZV+b+eaUDCxOZULA8XFmvSk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Z1kxvUZ6A6pwKaxOdYs07NFMnLFQMgt2NVR5MKR5RKdJ8c9hslnSwQz63pqgbJulNL2IsMQbF1Uj0IhqVuqvHik8GKPJT0wra1hxuKAB80yrxPtVbyBlDdvuZxuBjXIgzc5B2XcslaeodZFtBeyMeUYfEN78Sx7u3lzsX2A4IXzLnEWV5U6gYlyO2tGw+1I67OKRfL/w6Pxg+cNr2D1Y/t3pkMof+6e8VFnEeyhkMUQxp1V2Ba4dT5rERxQm3m/NM15XWs7KeYm3iUjr/wJ77M52p9iF3SQ+JEtiwuqdxH87uz+/p8C75KQGZkYJ4U3Ml+tFkpy6mGA2VbV+SCspyPZshoPoOHsrCsBp8ibS5WJxGsffo5IIAElbRHfx/SiPZhHr31Hxr0CUaZjlirxV2UaNC8juAKJnTOeaAf5rD4QlGSHrzxWiGfdfsh2XjacIAiiGQS0g/SVBRQGwugvM8LwLB+EnmOj4myOv6QqnnnkwApqzIVjk4XF1yfHfpH7dk/JhGcPpHO8d2ac7sRxEd2p3mS/AjjLViHG+9DQavRoMOa1+rr/D7sAOQUtsOyPQ5uP/wgMS473M7vHzFwQpDplc/7QfDwaYpGna2ncC73mPWyQkczyfilKRHyh2lScJhb/jbFFTU8LkHBd+hcp8ZQzg5ZIaIwouXThS4YtKdzAYdoQ7/3mDhB5gGACn2vGCGlmY9R2l/qcmAVMJhNR/MmYG2H007rm6+V0FFUUEu2NIooPc7g5ZMaqO2DhZHAeakYZnvsuzBrUVSMix8BpmqGjrjOGOe6udvQY/CDo3Ll3pYwGfME/U1zWTvszK1h0rAEaAVaaMhzKlILdpWFc7i23OF2lWLa42ZtsmD2HAkfmrjKABv2QcpZOFQVrV/T6Pf4pncqNQuF5zIdFyDAkV6tkISE0aTUfrkx2XCqnGHjjnWhgxyqpI2VB+ED8oMPJEVPXa4Qk/m+0JqK6oj7+uU5QePUGkbe9XeuhR2i5E8ZjtZZAYhjF06dcpvMoBBzZ3"
`endif