// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bV3Dh9jhgTgGK3ladTRE5bklvY/X9nnkseJJspvQnp7dqTtVKiE/BUH5N5Er
tYz0XQr8I7oOuW/N1U2yMK871naWtAINXBaV7CJS2hrUIEoymuf/3IaKr1iD
Z3tTvuOKVzNGl2yTRPvkge8GxTXivsxN4G3TMLlz+W+pJfB3NHXIJ1pQszXB
nKqVgzvGTqjo8w4V3bVqba3ZSWlPoP1FV5EpiewoQ9a4Ycgs4RW3nD7qezHK
C5ZenUgFsPYgrv2vGmLY/S026Gwpeno2hvF2waH/8LTkOKg9zOKEhN7Xa7ij
uIGxIa6nt0qr56XIDV2thvTnS+ugNfkx9HVSsATFlA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gbjW/YzE6jbfStZrv+zTfcuWH9XwmSBVKUYSz6IdNb49VDFYDWjXqI4cOMtk
NR+Ivu8kGdpQglVkEfUNV8gTGLZwpP1tpV4aBAFfaOQFMMStagEy9zUIZFwc
FTJ/icJAJX9790fAW5wl2CCTt8X3B1CEwZwBgnHqB54Q87z7pd5Cwjp8ASuN
eUu6hPVkXEBAPmQ3CxmpxC9bWKMSSLAv013xRkdlBIk7/Zv/90dzkBgop8gP
xGsWvDEvSNJNufbZKBdUCoEBpXH6uIDLZvidINBH1AkLRhTASEbKcTIS093A
Ifd2LVaP2x6iSq74S55nxxKQh7IK+G3za7IVdpOMyw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KLZFkTbasxrmJ7p2thbj9AmzWgidUMlkGXuWjycYg2CYr8C1qOrNYma7cGP1
ui9bRdzhQD8iR1Vi6zUiwkTduoeYEKoiSbVKAd6tYDWWg5S2DzZw6GH3Y20w
knSZssz+86u7/o4/aA5KmpcYaqO3HRSm4M+bIapEWouFGbTBMp4v21opiuPE
OCMHD/nfvDR4Tv5AKOSpD5kZlj1prNsksdadLOrfYJP2li/EZDtErExOU7jl
B9+2XAMNLrYely90Ej8OBFBQrRsen6u59ILTcWj2zBnvJIOy4y1sBQAG3/LL
O62e0wnP3sAF1IDCWTWXwGy5b5i0QWYfKnzYiQq/OQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WrihfJTGnYmVWTSFo7G3peRcL4PRELpbSSyMhDevacG9DGjsjaUSyjlwdFit
FMB7UPIdf5etFGPynmZbvur3geKA65jXisiIyPS66Nw594Na4ZELi5m46nCZ
c3NsJGqR/x6NOVZwOO/Q2k0JtTPC4J7IGo5GgU90iXuoezJSjirzcj/79NDe
dl1vJ3ogPmYu2ElsDYwbRkwocVf27zheYxT1Wf3gi9pJ0+890jjOgHFc2Z2Y
DVTTT/wo3vuDZDGC/jTB8Oc8j7rQxmrs0RehHa5FJXMYtgHNa/3wyrzCSWX4
FnQyc6PUnB6+f+ipYyaoW/UM2waatnWvJjjTkWBk1Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EZ54y7gi3O629rRV7T3AAyRqcSkHQA3jVdjJiM96SheepWMKBINiRv6ROL6A
37CDnCwsIIvni4URZeejQVZOyyjkPrZW98WbBMAhlcm95lJBaJh5y9xWJN9Y
qlXHhb1ZIXdSzg6penKBht8AsulAMuhTnGwMmSnJT2vbA2pHbXY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ar5l3f2k7jYRAoNjF3FhhMDG1z5xsmqgdp/dShETwOWeW+HkHvPFlZhXNsmu
2q/AK0r7OjsdCU3bEiEcmncPXwN2pp+U9C6wJr9Wa+nMYYbE/HTBUeWdyo7Q
99jWAdyfstY9Wn+uxXQd+j2zp0QuqaPvE5ewS6ZbuJl8Chs1MsG5YXUE+AvE
CzpufTY5qSfi8QR8PS2wa2Sg/EdPBtLNd8Ud6eT9ERxG5YCTvNrh7qqjVnGI
tKyNwUA+oYH9SaC2qWPUggMq7QuSiggQrgO/3niuw5V0k1TOYCCmcca87MJI
XK39TVHdM6zrw2rxr7hFQPAznwjS+kzNK93WCx9Ap/hfVtk85WNUnnC21MKK
sXJs8aslHOw9JDoyI3n7GNpF0V3VlFIIKH4SSgnkM6aQt6KeG0603d5dHS0e
dlaLhviMagHf+zv8s5qWiPDqfvCGMWDpeQ/X5kbP1HIRbjfJLCwOMRxPA49X
6ccLU1oUjpyf1FUXeJx4Od3NGE93xLC1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eHM19gBcIUrhpG55okygIyDM6O4KU3YLDom7WzGI/Wb/QiASKzJIO6CDECsU
gyoNA5jfgsvDYnVXzkHk+OwB6S/wsHANNnBdp2NCkFUl0xj9+m9YNPRDq8ur
XulPj9JFP81Y7aB8LDmhoeG6aA5Wy+AfUvPYYbYVAQzlJ6anXLI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rv2Hw4IKdfI9qDtylotokB4jxn7ePuqzEooomMRXNgWIlDVLCdYAws9xZ6pH
JeIgtlbX17pf6RtifkYqTI8ZfNCk64p5VpCZQwGGaGhPsgXQJ6cmNXwKnAiM
T6iJoaZszhIZOapOjZxNurW4kmuq1RbIpQBtr9etV53Zo1mvLoU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14832)
`pragma protect data_block
ux+ZXiSxQrUzRlts2vFls7Q4uUUOk9mO79UuSRz4FyH3l82OQaXdg/GqTJ/P
L5o2mzDXcRJcCIiZWr42aGbR+Agk23/KBPzQzaMBazX/azOnkDpHUsup4/Ru
36mf5348v+EhXz295l2m36VXNie3Y4zTt8LjI9B6gp98HvBxZhvJbiDS0RuK
Blz+YtppU74ReI/R5LzvcVt6CpXFdTw+DFJJTjb3h2YPPeq/geWeyRacbmUH
7tMugefojjbNrXg3x14g84KTtoNlh70AdYaNXaj4TOub1/Tf0E84b1feZfbl
+sln6nelXph/KU52o+caaWCY1BJRTu1GqSaWPjg0xKWi7Z2DCivH7RcuxyhK
MkgtaEiFkVCBKQ2bo3+ZXZqWntxdUsX9d1gCm/PRhfqghnx+T2yFjr8OYe8L
FlKNwAWsM3iXrrY4nYkxDEZJsLFovOUM6q0mzW30zlMi/6g0bL0VmAg35LVt
C4CECRNoiKoknIzvV5QPw6MT/FwFkY30C3Qk98PKRd+nXLZ10V9UIqnZGuIP
ZLmHZV6IfHt3liBt4CcP+1EtQs0yH2fgMeW5/5GNdfgh7RVyDidqhDiiXwtg
Lpr8UaVgWvs5gX+ekUx1n87LnfSu8EDLb/xZWh0g5UVEH6W07obxmSMKULNF
PNY8BHSRu/qUOAGn7LdT/3MNUxPWn0WhQwmQoKGtWWiRDNJMg1+L2kXI+mRW
IEuu4A2PSC/ksaAWb4i3GflkABk6/YCI3IwC2TOkM7dLfumInpbVIk8J2rwo
ZEz+isawe0fIGpMI/uW3Mv3XoxwcPahiPWi72puxsBFNJBFinym5//k0bbCR
QmJwjM0I0ufDoKiXIK1YocneX0GffYCelXQ+b6egFcGHhP8BtluGRU8YmsFZ
XOGP0tJlr9/tEaI6ssI5mZRYeNN5Jf61Wp3nAenFolKc2veQ/W5GDaqSlMvi
MbysssIOiGIObvyQSUX56tz301c0nv//u5esYwJftYIcTaGkYxmiBYPCdLSD
DNN5JP81HwVSgBonmpB07tdhHroEMp+q06LomGS6Sugw9+BlykTh1MYY1iVK
zNaWeuWTxpGrlENNtYgMcFAca7NyH15coreX83z3Yap7r2mSC3lJJ4ELrunf
dBVnzOV2MZNEzcVAd0QB11mQ7A0aeeyRAPJ9s6DQ3azVt2GFoRlAaW9KHiO5
kw86criPCr4oVi4E7oqjCXt7YpBkPfJIdI5FEMBfYHzCxT0vzo1exKhC3kvk
QZTWbGT7c8wNVFGrhTuSrgC7Fl2FQFVrtM3JJ6htVfdGxR7o8fIVlYnwzr6D
fwIoSqgR3xPGRvSKiZCv66sf+ou2ZDI6zxT2WnnClIXAxg1BEHfOX6Xdue54
kznufjqnPaBYQTtdSzAPhiM5w82fEgYajiyzKlrme+rNdxFBQQMFwXg8GOBC
jmDdLRarXHY1ktosGg5p0UZBcvxnb4DddvthAfkzDJEbwg1I+ACU9gy87y8X
IHfi3m2zNNZtYz7Cca+p7KKDtfjetnsNHFKSZ3epIOYJL64r5ShJH1rgqFHU
njCJ0yW8X9vYCq5QUcBZrh8Xv0NXBND5MJk2+GoB+0aMvq9eeFIzYewBbGJ3
Q4CcTV1j4MTqxEClsnpBJJ3SNvahstr8cZP1I179l1M5VbjPyob8lU5FHfn/
I+DQoSvAG47VGqmfahI58uvPjj5WuH5faPmYKTA/dnLWhx+HLYxiTS4juFuj
fOeA5n2TsLjw6YxA1bDZ8RGVMoPIWNxIdTuFOVqufqmDvF3AbZKA38g29MsW
CJ8iG2u7VOvNF2hqDCyUISdIZRWXn5mu8pfb+61Qh/2Tg6tmFeB5RTUeHSpQ
c1PFMVxjKrMcWFt5ZNdw0d7vZalF8ZSLPiHvfXO7V5xM4XYHtLx/LVi9IMsl
pBTtBR8HzOAdDasCnT0PzV36tdr9wqKUB7UstCioLk/tlCLIuysVZPh+Nf0d
SJNIelgBZDByE7wLKgiEDQFiPTeXnnKYZAcmclRE7jV0MbfOTnTuPx9fPHvH
p1u6bWIoosiMCKbGUnZew64G4MbHA4iNPLIw8N4JF7JTOOAErwO/2L9EQaKa
Ro8DSSdVFPzwSv+v/bp1XutPwyP+rj/7VBRg4OvyO00/QV7geJDq436c8sGB
96OX0+JaZ64E5dB4Epui6UZ3gGTpHP9/d7h4y3isbOLAu7LoCt+iq59l4mQX
WUHwJIMEtX6lc+/vLmB4GfbB/LQYZWoiIj4Xj8knJEj3KmqeBvR0rBseyFCu
6LRfRPpfteNCiC3muYLjxHl9F6nMIrr5xHI8a+kh5VD7oVhcvOOh4PDMHDOS
xxCcdPj2Q57BmN0qRzeVHT0uRgTz8hK8VB3Fnkvr5c8+ZG2OHK3bSmQ/rjbt
Hfk0o8DzH4W2R9T0A4U6KJKlnBEBf4J/QaRbk2efqcvTrYhh+iDGrlVZMNiR
LFaW5A7eCusdGVdsasXXG1sNwOxgshCrhvPiJzkPXRte5mXHbK1/YbjFTTw7
tEFZprFC8CB9hQOCDQ9+czM6VmG4npjhsU6kBaPNef8p/7o89/hT0lzdLnRS
AzC1lwBPwRfvwS/H1fz8+IrBlRNYIrxUC0NAEhT7u0O9jS48XB6Vv79x6SvS
M9Y+o/YRv+TaO1Sb7cP6QmAxpyA/hSzGFpP8xN7/VV72LCn/C6tbAxHBfUue
UkIoOh/AbfDpQixS0jmXjtadJyeYiviICFIdgu6VJVDBcsc3EL/qXOGL4SXc
+PXeFPPArrjWeL5Khmn/8h2YDD4xt1ReUFkGAWzKqaDtYVeyFE4KnZ+630Pw
JsgAY49TxqnjhH9R5uQA8sfQ2yHIsGCIiixlRJY1m5Os4dWtVeKxnsyS4OBu
B9Z4DCcm04GMlS2wdUrwg3krv96nYJ0ds5Wb5rbncYP0o6dm+18cRCFV4qii
b2vm4LoDP4XUsuaM4aQ97UYzqSylsncRYYYc8vL1/WMF1r56sCq+Sl7mTUzV
SOzfOxmBcWH6xvMJmSYcUdsUXBZo9UyBmbrmLwhZeMbSo7y9+HN0j46XL0TN
P6A5ibWhv1KqbgmtTL0GKDCfEM4KUgd660JRRqS5K3fCbT7eA11qAvLCw5db
R3b+pBoWB8iQojvHIUNLV4yMK0DlEKIkUSgYoRFd/ngiDUeG6hcHLla5VSMS
WswSgd2JPQiWUABNHOS3lKJOGD1KO/+8HmpwKoWZUD09ICzLh1yCb3gjPe5t
kz4jN4nm7UcKexotQvtjnvRw9EF7YaiNRKjwARqvY106R7leqa69KuRyCwNQ
9vq7Q1Dg587sfnI7vLS8D+ZlQ2JYxsF9hBRLpBd00qaO8AD1LNxCjE5cqdNU
wiixx4PFZ/O4/LfpsXErWjOvetxxQarOqBc2ZyULjSyuHjqrZZfPDMLtaedu
qpbGiu1/pAu5hIEptoXB19dF5WtUJfUf07e+mMVv5OqXjXxphz6KDqvRPkxj
aBvc3xLZRsA9hUBThBbujPfolQzWcasXbClio7YJFKvZ+6os6/BZTeY0JTqk
e7knDbq7giL4RY3mmVlX+oo/0DJ62q+6KGiuo31X2WuJVJjQSy6tQKPjlBKm
LEKOaf1bJsrKkfoZdOzXyKrrmO0BES42jpanIVVbGHH7ksynW1poVKDkS8/V
MxSHozmUZQ4BmvSPKf5XrP7130W/Ul6rR3fL56PfhnwXGsdyT4rgDFRlEUkL
3ED9kzdKmm5KE9p+2TuUQa+TbeO6Nf1pgwbA8iIFwssd74hkokof5KZm1d1D
1WQ67VrcR6LB7qufiFvIapUeuMO/V4asnPXbdcr5RIWAHfr45lHLPTFz7g5y
o17xPJqE0n5Iryp16f3kbnKEezTTqos4N5i/2Z/1sptMQNzK7321kS5nH4O9
Aiqy0CgABYejAEvWoef12zqrCP+XQp3mCKl1GqKeEFPtapeaOEniEfQ8GwsY
2e3oZRLZibJ9kvI4Hyf6bRlsRWWV/4mgUzlzMzjky1CZCrC1tXkngOS+vIjg
6Wy9AY4xfDeoWljJ0xCdZJoFoPB8KGDtjxBFNdRt8EOzTiR8TiHo0dhfcwJl
MfTybZbw6E23lp3jE3Wy7A0cdAOuW1aZzA5bqgDZkA1QaNK24EeqoWC2JR0B
3rCi0wELb9f5kbmfQK+7NwtrTb9wOj/sKHxg/10rhUaza0zPNe/2NztUiDv1
/bmhRR5ct/WKISW75R8GVaAHk10SV7UnDvEum0hULTYGWTVCLm6Zx7+74MFu
ceddL0OLLyoZGmDqVPKi1wLGXAkWNdx4L4QNtItxJb8eHwxbO+FTEyH6z5KM
CIUQsSimfty+N0B96gP7hvndavhjTiVDPT9YzpbyeavuQw/cDe7/28Ks5sTj
e0e4qvtBodC4EhvMK6f1gVsxJA9PZxZq6ERZ7PpcioTUMFxoFFGTbiAfWqQB
hhjfULW2nlxPUAtYlRs+n7UhhyGsc1SfTfGJ6l+HiboJojeGCBYWx72r2+0S
hVu92c8TGXor9I1RSMXJZ/+d2j4jONrCjylpoAPxBxkCpS5KsmL38JobJwBe
H396TCLmWSKaTd6Ylbum9Fv4GMA94jKn+nqx8ubYGXmyT1p6FA2pzX3oRLVU
EVmHPKKDEtCET7uEN4MW1RrLDTxqXTpKwOUPI3ChphmnrXLxg0OTV09TTUhQ
stFi6VHthFaG/b4DTDeA0JzgYYM5v2OKigSzCmbugbt+RNLx6BFPVJ93RLbQ
1wv/I8rJThtH/WKr6sLpmA8U+cTx3WK0fTzMwOEx0jn/Z6Yk0pKwRE69nCRA
89qUpKJMuD+LaSwv4UVIWABWBCb/ZHF2Shq2Y2IWLhWto9WlBff9aDcjeDxN
t08ZnRO9KKTJ3H9V7BcxUG39JD+l2xSnVxkPwdFhp4grS3WfnHmG9QAOueSf
0dVkGRuAZV0wS0R5W89O28NMW1h7iEcgZRp0OhqAjgsN4rVL1/ZwpvukSb+C
9gj2djS78p7WRB0zAXfL6i/kSQEry/57BHZMR9mvGGouSzH6V/QjHn4W/Zah
49uu8RGDQ/breW/AnRHzFZFr1m0/n+cVcTNmYpy0f0lUY5fnIhVCGuL3PfoB
j4jyU15JTZEmAyKeXdZR5wuvQZJXWq4bsdw+8y4Gruc1pb6D68AMBGQieGA3
JPI3ykK4iCCaWo8yTgPsSF8rGigAIUqFpv87zBw3k4EL9dl7vIeI5JeXW7cl
XuNEc5X4gumjZ5vq8/G7yeMl6ULLoYnBDspK0zr+IjhBV5KEuBR0+Zw2QKni
r1voLTesfkd4HKWSSDoVV3Mf8rRDMQQFkIc0PcX1AjQjnAHehtEPI2g/TGu5
MFsZZSP8otuJ+oBCaZd/3vj0eqhm0JXEugpaTlRFlgPwy7rBUjfI4p8eL0jF
R7tfQYPmGj+xNCdIlAa8CWnLqWo1bX1Ohml/xdliNCE3PdgahbPh84twD3Cs
GzmIX6hOwaqGX9rO4ZJHFKzXic0UTq0ML4RCRDm6DKGnDflkFXNbQx0nsPzK
IAEjnmOQ2HMJTxC4Cu/4UqNQXihD0c7SYM27CXiHjwT2pk7m6HCdZYRRDw6n
m5QvI3ONyh6OVgCfEUAjUQC1BGH6P90WOq1dlLFA5x88QCqyvlhK6qBIJWzw
e8Dg67ubJjEeBdsXi5LaGwWyfroOds/GYM/9DkqiGYZ9lhELVAuC9j7EM7Xr
PGSe030DOWkeqDcHPEvqe1yLr0+18zXlSEmZTpZKFZ2HgIkI2r325vhgBeqC
HlL953J6roTrEOaEAt0ezjBmuA2j2e4GRv5aX1gU+13V0Eym7Xhny1MSatiy
zUTLKTx3SxfoniPeyWPpXNHaj+A1JuqtmrW1G0ZwSuRq9nmaYW3pFnkclAC+
nRTYtWKq8PDVoWnHTS73JXOY8hIpKggL1qa3XCrp7VBxGmhyhvOgOnHY7AaG
WPtW5d8Dmrw5ADo760xLID563FGgVoTMF0Ukp0qoUkLPUEF8mDraypa3d8bC
/m2PRPGyiWZqBDxLO+RtlzoAz2AEacE2nNGndpW5M7PXzTrHy9Cdzhnt7kMB
5bq00GizEvMrHgba1jlJJVhdI8BHN1NEbj6waXxredXtqkT5PmzkCwUFXreu
RdJ8xESt52ufLtyYwVSeQlibTt+MiVZ9wWsDmaCTjgpZsL5DgfgX3fvNqZme
0srB4bqL319dA8nbTzbmgBYWQG4FjBmh3RhZY0xZDr/5jaHXt5p2gwXx/bZb
C4gTVymcqKozjrP+rkUfLAfeOS1S4rg8Ie38fGTwOcT8AeHcP84SX/dmZbwc
gzY3aKJARmUWJZLaaQfkQ3MeEo9dDTzi2WD4NBfz2Xh+bAaEhr132EOyt0U7
6SWpFWMBMf8jCxrk6YMMgzgjEI/OiPpHoXDJzVUJIYG/5umGFcEkjh7fXCMB
whtd1Qs+pFgkmBG2AAOLlO6OYzluOZ4yHuM3AnCqN4VUDarj01JqbJOo4CSp
G0Y8REOfo+ifVZYo2iwxJ1yUpodUYoOgzHkGAmKqL4ZIJVIMNF+vNf2cE4tn
ESk6U6t11QL483lnnWMl0mBQOUGgq06Adzjtg+M8aZKGMkh6EWSyoHWSIATT
miz0EMiDh0AanzA3xnSphxM7lD+2qeprJE8eNxkh9epIrLOAH0xe+96KvY8m
TlXKTg3in48eupyfbY42eQcYr13KDKJsf58U/mz6ZorzTco8b+4gDDiVEUNt
f6c83i3Xlo0n6qOU6bUHSEJyLozUAaJf9ck37F7e1hnQdSZVhjZ6QcMNiep+
Ky/Fa3254HMMakieLSesix0eFTucQYBVgUhG90GutYqFr28smOgwoUbjUCAv
oe5i8rQgQ5cmvehUgIM5Htn61ojF7QDTHjo9OISFWrrcZhgV7xG8D28neduE
KSVSZbDhilG6NeH4lSYRWI3d95LdqZBLOAHxjyyEDrmw5v5o9/TP+y9zyhkI
s73XnO1lRRpkdn4q+B+09OxbPK1Xmmrl/awoIg7bZ5NujMJkGGlAkbluH65G
e6JUqyEshUPwSFlveTV3JY8BMGAoAR/+ga6nM9RCGuuSVfbicVq2AfJTUeaP
/tfZMQaJFKnGItTkxpIrOLlErM8muh6Davlej8VOka9xY5f5N7cJj2m+/sK4
Q9FqUFYk7UiXbDd717Z3HTTemH1y62OrTOoA6TwpXjaOcLmVVvZZEqcZShmw
dYoksz35X+ux+dEK5O09HyhOvP8e9LS2gHNeg0ABSEo498Z6hl3euzkKD6Uw
bPxL3lIw/o2K7LFYHFxYbgpWoykuPa/f60k4v680DbkuE05x6AKJt3ua19F8
lx0JnExZ6txKYUnq4jtpJ0HBob2iyLjsvf9D9uJHE43K62Y5xMZhLMvnX+qv
CrBzcr6eHrS7EflBHwD1QEdYSsBNvkj4SOnwLPj1n72dc6GA4w0EwcnlogFz
xbLK6yvN1CcjcroqYXss8jxzvg42C343jgONP04shEUhjZLvijjz5Wf+NNDs
ohYtpW5HxJyFF6V4ql3dkNTll1Fsi5T2wI2GGYsfgQe/qlgb0jXc+JTd9+MR
f9QfyE/FbZdifDNMEpUDF5aAZNWw0T3c/mYPPJH5B7sssA9qVXIkO/atyNEa
3kmzjX6iVmEWPxDzD+nyQ09rwnjUjbzwDwUBCHJni5JYnjgxPDvYZz9sjtCR
O5A7sa/O9ejva/32tzew4TO+uZ6JTYxOLHV1wEFM9Ov8i6p691zl7h9TXyAf
5gEuLLBtEC2CR8EJzQ4x7CI3RL1gaWStfIrC0b87oJU27yyhMSP0stNGEPuT
M+0lk36he2FAz9ta7tcyA5MbYcHipRF+gDsvTaf1BSV4bvnZQUCz0pRbtx8m
RdNNRvKX+HXIByz0AAiFm6j6QP06x7nnQIaXwNJlq6jyO3C7Z2jO7P7zTXOZ
RKcCfQg0u6WJGfFZyDWn6OEf4Aq4hF/P1tfwz1+dHSm/Y0VmW7Qyz/siSSbt
nMrVWXDJac9eLo/eR6LEHBkSCjgzngvb2zHU3yToXheMlCJUdPvRMTEa5e8C
+GlC+tw+hezA0+0W4rVCtQGeRO44Qwn6OkK5TDiE4Cs3tKm6JMhtNfrhwJY8
kFJFrn7wEUcd57T+c680mMWnXIUj87IBseH9tGzXDfoGVKawe+8rUTRictEX
gQnhXE4hNrxSPZqI9N6adZ4WeOggSQCWU4RFbsVEWkBEHG2P400WymHMQDzu
DT4rix6pcuyBluPi2z5AXzu62hMn71dDNjxzXDJjP+vFfHlH0bZwG0OYWJ5T
lK55BwZPKwJMcPFDthVDXUpUUDjZNXTcdMVUyezN3fztY7Oo+Qe6gsKKPq1O
rJNk2Zm/hc2oeUlKRqLdGkWYdI57zjiYXCe+XopU+F4+cfDDjBFxmHCcHzKf
OCDQrj/Xnz19K3j06H48a1uP8MlEkVtDXUnh2R3mIiOAqmSp8Sou2Kgqcf7y
qCIVEtcHqPdvL73RKw2AvgGzOpt0irgxx8b8LSbeKC4wBf/J17n6QSmAHqUe
Zlw90p6pGBsy2OqHLn02vYSKxyPhOmnIuuKf+9E7jftB7JU2OAzDFd9iSzBG
MBgHIvTocLhNu04mjrR90KtR/cFCYg1/Ie6EpH9/IPkiGKsD4rxs+WuK35FV
QfHICs0F3A1rMOECpi4L2ozSAXHFFS2m6UFg0Og7ud6oIazGnnYrY6b+XgUo
PMpNNlhnUgu8tvz5bCkI6Ma/w7KMNplldu2KL6l1F+P+mnQ6//velZ22W3Xw
9Ujbj5PRSm1iHzho+VOBI5m5QBIY6lMN7eAlVD4bEq0L6Bor+oBiGlJOuuLi
+AeNgTNjJzOfPSVkhoYSlvYvhjsSYt5usj65v6u7A8sBJYpHk7OatwFooIL+
N3ar5PRD76mNaoR9iPXO5cb/FEumFwjR6M9jlxXJoNn6dkcC8ODobgYfM0J8
ZRO8heBVPy/7vB+vcgr2H6hX2ckZ0zcM+R5tM8Eh44ikI1dL68mqluxFo7kA
8sCXoJzzcSTqBHtJFJIu3vLaq+BqMAkdLrMoEb+GVUZiugGEVeWMJZD5ToDv
PvfD7UA4b5eYI1jpqYQ039Yv/R3PZZjS05ZpIEAwTJjvKNDODKqVihmzOvnk
UlbatGQNfSU+i/N/U7v9fZQnMQkuxvd78WSco4ydGLgL9/l+DMIOvF/uq1Yk
q8MoYMMPmrRfNVfSTpNiX0r/DEsd1pbPzj6T+bYX463MvVLdedDkRSky5Yf4
H85KU58cZiK6q/NVJnKj4/HYQn4UXMfSWUomBHC1FvYoo0TbXEO7uZHI9dvH
belOGlNxMNtqm2HKTIRdJvH3J2oq+py1N3jgugcRzH7TAVsjZRnViotufR1w
FBQzkCYM90WPRal16WiXnD1qBcaYGMcwTSWOx1Ox0vEtKoQw9IHUZQMZk0rd
amhEYqvWsC1dZ6GOTsV+kA1rvT4Xxw36DPC/csRpPNLJRU9WLK3VTBIY0L//
hS9SQDaq8kzBPr2fGWp55JGQsLwc/n77cXoZ6byRI7+4RRUcEvV7hFdUqP4H
MVerjNrejs0rLfA2UHgoXsFPWifDCDrvsAHoZ6wx9mgZpfES9N2zVq3nlQDW
dS8m1SG6vQgNCzUCkyzTgsMytVvSvDwFN52PHSqdL8YZ20qxfX3zWiU+jk0G
vsN7m2n0AFiZbaGw3Hf5V+lP72Sn9zdxZKm3PDuLZIktg4c8ti2Uj4rqp2+k
vAWwhsV0oLHL1Gwom10mGksz25hssFMMPCqkxUMURYw7q3b5u5alHXsXKn9j
LLGIceClN/rCLYEZmPyp+dMU+YsVuv4YKtJqT0JPcnnyahKttBq6sKzkLQi7
aUr3FC0nMn7drkWiWYTGYlmvtWgmUgsGyYT1UvnYgcXomMbxQEp5QytbEQ4x
UpUVcy7/qzUX2a3fYJMNZwB+lm6mJ5uFJN6H6sHY+1BLAoPf3ZjJ9nULRdk8
dX89TRz3BnLqGHvf9p8bTZgd/NMp1VAwPEo5erp/NHcZFUagoQIVCIWHVNV2
WWvloh46aK9AfN2/dR70A6fbDIKETQGnkIb3oZ+c5CWX/vTMhMgo6PJ2bw+1
cxGMk+kMA5LjdSoQfBVmx0Hs3yLMmMWMr4DKnN+LLSOmuEadnYX1tH8+6D4e
VBewWf7oSzTVUs6VTbvvl+ZSxNVvhqau9Lza+6fnXf5JRhwKYGZDHbNI3hm/
XnqF7WSP2YPsU56ryMERHjYCCmY+QdP89c3LbbH7cNHDpLrRJ3uw7QS+g6J+
NVewj9oYI9W0XyYSME+s2658Rk7meIrE8vLG9IExSVKbjWy8gCkR3caQdhCq
vO/lwV5YbeJK6u9eoQpT6jA505odxEYlF0zUB2q/9AS8ZA+Q8AgooeOo0JOL
cDchNA1QbmdJKwVdbD+pu+GujWaZXmnI5/hgidHzJV8IqeBCiALLU2k0uEWk
GL2za1tHLDdcmeBBnMaKc/uPJ54hZyheZ+JLgXKi/m1uvyseRbf8vcYrOa2L
toah3PRy6kEajYlkxePPqA+aoNRDnjhUhXu13u7ZY18kNMYNFTguFGVJmR/W
I/IMXinPwpOCpR69JvhIFmtx1mmnvzjPl4Edim7GkDCWyswsocEpH5YssOti
9ZVNXz55A6pPpF/wtt5HkZgBv+H9ehlHZGsXVzFoOjtFUIU24zlc88yJHXgR
EgVRhhYUgZu3idSiEAr3Y9FKYBn07MhVDV+WJ8kIffGqu4GkHeQGFjnjysSK
c+ctNo77JyBOIVgWpO9v+e7NET38nBs9lmbcY9XS9AoUZqTYLqiYRBY5wTGJ
dRn/Qjr3icaG0p74vXukwvyQ535KaslLP1xBHPIgn1pLQTYmbrqvzTJ33nsj
9OyYhOfYpcPIGYctzXIMtudU/a01fJwzTIL1p/RbHt8hxHi5O0aB92fwjY5s
K6cN8K9R9i0ybt1rVKEsnmLYgSBUDlGZ8YtumeJpQAgWINwqkAd3tHNuVwJ4
V+h3yLk0TVigONt7oaYOOxdighucV59DRHWLkiNGbTbQdR1txK6BMIkSHMk3
ccEUQdNIBTtm9A/WpkX3CKl73eXL4Ew2+fa5zwaNh1ShLw+8kjU9xg964UF8
6/9Wrzi4plDhign1KQNqYa6F+AB7EScqqaY6qkq/zDIoOVAgUtX2/hNUcljl
iwsTRMi2rIMb97xdVbfEPqxShUIloY1jGDjC9Zwftd3aDN40fXJXh/NwP0uU
b8Cn1jFO82GKRaMJBWvE8khCr/oLufdVBZLlMOTI8zYk4JNtSaypGZ6p5do3
IsGOpXzlLF/lOZa0rERzG4/tmpAJkXNe5UEaK7aBALF9utiPmUoAlcZR5I1k
Y+OBHCodcDaCRH85rh0NgTf1ze3v4XVzp5KUPqU8MfXPnOIY+07ES3qePGci
XJVeKI7/qUJhpMeqdXPIsMUIj+pLdUapLOX4OK2i1sX4i3cEeZZvghTVbL4X
OB1C626Wn5BleuUx40YvQ9lAdeSe+z1tbDq9rhORKwOvkDGqD7Uvpsz7LZ5W
AGypB5RGG2/kn6bhAfoEl1ndr5XnWV5B1ZJLI55CIcG6Dj+oSraHCM/YuQSm
E2p3cTWaGlvbKv18p04wjL42BbrIFgTEg/zbs8PWcUDGtzmh1xB7NHuyTzEZ
0rHGzzsuBPzr8+8x1JlT2rJP66DI9Pz46mHS5AhyDqIRcViZMjlKDVacEWVO
PcSGCsByIlbDtzJ/l2kU8hvoTP2TxrPsIA2bfpYDCxYCvDnibb9x0B9vsdTu
Fe4PizJwz+ocPP00hkPCFsvKY0f+8NktDEGSsEi+tjj5ZHaAW3P8rJb2fozx
CqObSqkjlSP9spgrucclCGWnGx6a9NKEjS39OGHM6kdJrTUPKy61N5u/AtHb
TWrqz03pF/Pwp8PSv3GDFHJGB16jhBn+57IFhvB6ZK/xVYHB1rziBlvmW1i8
B8g0o9be7OJ8k+5xq5mFwp3V0G5jp2kvbw3Tnso8g9ihGcIYfpAGlnncbGrM
t7cjJrUZEdETLEnCJOj3NwKzTkt41LK/EuDNWL2abVigrMoy65vKAFtSRk1R
+K3pFksTU4pUxiWm3tMnCX6NAG9EzmpV9CQCUddPBFvtJCAVdXmx/E+k0k0I
O6OUGexOy38kNI3uCjQgZipyd8I+pSLxY/JZCvjE7To3q4Rq9qoQC9NiBoom
hBhCqUAf+C7WSi4ya1fQ0Y6TXbmq95rwR9kLbLb/DTatZfHZjlkUXH8DkBk4
emgsZMmv+tSiGBoXvvaprxCGco0ba7XDZf8tO8VhduRGsvGp717qSIXKc+Rp
ZnAInvWNvbZSCo7Dz67ggxRRKalFAXgBfiR5VOPuRayqWz0evZXztT0uLObG
pSkpV5M/BdMBx3kUR8XQ9UnGQaum8onqJTksvH+r3YzwHRotNEjnhvH5p01f
z280CKO/QXXrp6OuOmNTDOi3E6PCoQ8qSoHkdAqfaLqxG1NCb8nTb+JHM3uk
3UllOrl8huGzvRIplL/pjRrDBnjy9r/0u8U8uK+v3bZbWSGnhNI/fhZvRqH/
7LwDpTtADh4OBSCpeQTK/NjC6Rio8U3AIdf2G9eBnZ2BXFItDAQtT36irqiR
JKj4Px/8FnwGItwvBt+oPmZQxRlSHrKevN5nD9R7oZ1M0FfIQ24Xzbn+pk2Z
DjW1qiyq7ZnVJTDZbcBErXiPbfWb0RC4amI/eQpd/91rsgmliIwB3hVRQ2Zd
kSh/TVk2G77miNzeNzd+/m1Jtl5BtFlW/JwXPMBDk/p/upYvNnDEVqwhB9Aa
QQChbCgJIW/xIwvMbS57FHvHSMv9kK0rohLeXlYUB/hTexK3fkLYacbTJeOC
PYqALNHsm37qm2z+7r0TjdaNX6U9DKSuPFs4v8lr1yYgQNO5nIab8gzM+kJp
ajsQikCcyieHhXdvNv7pt9opGN0DO3pTNjcgSrycchbbUg7rZw31116IUdry
ZmpXytnZvpgIrE8+4zNKj/iZJvN3Aragp+oiXeSyRPuc2I1KXN4g80MgdjIE
rFyN+CxQi6aNMwm5LUvaQbtf1h2lJdDyXwJaZUFNGBkz7+lrpiucUhY3A0+Z
pP1cZglxmD3XBSp0c3uuKGeN2OPolKrKC2hpkcTXwatelaXVeQK7FFgLYzqG
tswFdiyTsCz2qA7y6bmJH8cfddMnKytRYINqb/6jtlE9Rj+E1TqBs9ITgcld
HHRel+f5q+mkScG5r0Mxiu7cbojzl5yyswYDqM8C2GvlnDXwYBo/u7JU5CMc
VJ0eOGSR+L4jerEDgWWUeYSM6HMagOtJhEKa/S2vgWSWL5RX0pHCYTSSnbYR
OxSZy67l6jZrSg6XcugvylzVMDYh6BQcstMENwaR14mInrb9oeO0rHJ23VsP
+WLqcwhemwSb6+PR0u8lpWOPFyA8g8Pqz0mpB3v0llXKz0xwBbdeuNFMQQYd
vf0Dik5rr7ggVtdVxjv+k+f17mDdNvdNuoro2ufFl9wCxUucFpM/EtzRswfF
aRMA5ZmkOOECWuQIAwquj1f+1zOogBzLO3EudeoTNFxE8b76zYn5Stfp0c2p
XXWrG+lVZm/hcyTq4+QntCny5yKhta6icQc3oGH81fHKMSGRVImkB/4+MnMj
J1B0uePWVbUjIq4/Xgqqz8LbAcBtC+TvQW9dQEdyfUepw7p5sk9Mj8ismo1q
Yxgn3VJFhSZP7fYZe5v0d3rlIOt05C3/LhLcnRxuNA6yUQFl79ZbMYgOJYxw
CxVC3BZCFdTMPYkGVW/vdz+BsS4AdQwwBwHCVLr8dSSv2Rumr0O9EwxLTNEc
gmvd9Sx4m1Q3eQUiaOPoAX63aeH5gK856RZS3Vv6QCaAQESOgE33vz5z9bfY
+ygvkTE3CtATXb7tEOGfT6N0n4bGiGrWcjdgvcsJ0Dy2tf3LPHtDX0MyM17o
Vli46u4n2GXCQnOgi2HQ96XF3qzlQ3BoATfN5K9Xh6ycz134sQeSQL0OKIA6
ZRAk9scsvAUT5gmrJbeABPS+ZrKzA8hbgu5bbBDhkeQfaZtEL2nd5sbLDfPu
KgWhkKnnu5GeWsLZrRhrs9wINmJSKJUlbceZr4nGoND5+Jwc0I2S1u57mb/m
TghdDRPtUjOE1vicArfYbLrt1WnFhzrBNgOWQniadHX8s5PS9ssIzUn00YBf
I7EYvEkA/H7dIHplsc2zbdxciNCmdAL7Hz5wIyDzsIzqeSklDDt7XN3KH+Nb
iBUBmogn7Mc/JaPb8OLt16ps3vaImEg151Dp6G2hHivjNvQ5r6FD8Ks/9J3V
ZtgZ2Ck5fqCwhU7u+36uerlVi7TCpleA+3IfjB7Iflr8jipBC6OYWhBGKtaN
k1QM115w/b3f71F8FZaLlKwMtqtPYw97j3KYJS4EpTGbajbfQsRs+SLrC7lH
R/7gGYSNnZbsC3GWpSJSv67NLQ2ieYg9vImKOi1yqjqnK8Sx8NNclfA9tdny
dJEfJXdI6zJvVK/Yd09IaDxNBt+ezD0U+D1fmKLmC9l8DYyUP26Th5Tf68Ly
uMTnJJwmmjVEarft1TGroWHerjndw2xVbWfoIUXDfuY6wn6ctZougSV6jz8f
IFNs0n78+0NiQ4BQF7XkibvONuvZCqUcO0h2fIzY2q6BuQxwhnRzAw+Xf1JB
BnyLOTwXaVQPfQPC/5EGIuWUJ2JeMVaLgDO5yTn2RbnRM2bv95m/aZMSe25U
9YuNDRegRzJ5yVtdUxmvtAyqWtAMm1fZ60jnv8zpWajwiwAehkpt3AUMAr44
20F0ExXx8TnW6BVGGnrnO1WQ/GHxL7uHtTraDVaywrORCXbWr8/VO5xsmcgT
uTrz/uUK/6e9/Bkqv0ELBLIWqHtiUEcittOmzA9ECzJDUkgjMWofqNfmdXwX
DvRE3ElR1/4rdvp+fOeRdh/ACnm+7YURNjLglO8Xh0/b1wQb7dda3D9RkIRT
r63m3HbSzRd/I5l8cg/FUULJhKQUqZ95FkVOFnszOji7B2IjrXQQsvG79UYA
5dLjrLrRH5OPZIAC6hLMXggZLLHrcHP4F/XlwcY07HjP5lntFc83SAmPHq8x
6kIb+nXYBhWkjwIiOBNUeulpA0FDxJbc20PhxWxKgf3/CeRBMx+4ngjXyZyY
eKd0Jbj3SHwSYZ2nr03FvzdHeOeBTMdJdodUJGX3Ym8D8Istw2SKdNznVbH0
rK6muYSMgWVy4D+uyRh/m3G3MNcjnYIF+Ejrfj7B6Hxgfdgz1mOlp3gW9UvB
F6rUMgbCmC8jA60FWb2GPr+Yw9cclsy8IzJZ1R9Krgg5KuQ5J094c2u8u55k
o1aeZqlYjfS1S649OMoSDTMD9ys6fzVDe+7KKeCqPoHNpmFlk06RlF05HeXj
HWegJUF8ZPzo2glGEUZC4iyn91voKslgpeZlDV/ZOqeGEOIhLY2Iq2GJyMa5
rW5rYaRjAZweI9tgHrqQe7+NFarSKWaD/5aCGDdEcOdltBxr8WRQrSp5twfH
IEdiyB04iVrTflZxwSXX+LSBcDUGlwoyuaHYxkdhDA+YwPqyBs7URXMWY8Cf
XcY+kh6olImukECzv5ocSZyeUrK/VT2Q4erVKLLfQtZy3O0CeGKdpp20iM0i
SI6MoQHwedRA3mRL+1s86vecsR30QdCH4JB5usLe410Nh4TYVWZYz3XZRtHM
ZWXvTqd00qZ1LZ+B5M0S0P7s3amg1vpbdMnraDBh0FkFWifZO6ne2SANtQRC
fHEOntS9xufo0OGMSHPJGX5AFKyPyRaQJsB7TUCMvmdHhvhwZvUD+iUHps5R
zT+7mKUX4VU8c3csM/pqfRYtUacztG5OvehMyCGI1skOICkdNxWrmCv3Skxy
Un8URVN1MqDQhGxCV0pBQeVvvtfX2xoG+2amCy0z60Mm8b2mB2dYNvHLnGoN
6Y10LL5J0vha/ZtcxmyZONfzbHhY6I+SV+FOwGPIDmYLgX4sJwxCDYWK1psp
R7pbGdtOccDIIhJrPs/MnEA5zXK/v/L1IReNvK8FqiYYwP35hdpF/OwW482X
K1r8r+6xTThBXx7XcKCLEzVceFBpxc/AXT4fRj0ApBlDClnkyiugp77Qypc+
+HkXx6uuWlzaCRE1p21/0IV3CTnzijZhnQJqftrVT1RwHToM1oaYDVxFgGn2
BTfKdATYRWdD7hnWCSBJ9OmRqu+KFX5CBP/ut6Zisck397yUTCD4hB1IqDTH
x5Lx1O5XFJZlAr81nDsgKjq5WUL1rJuXoLs5i6bJ4oWk1ZXExP5fQJkhzy+W
1cas5/HZ46OWMOln45ZN+G57eUWxaE0vWrWOhJ8uGBzGd2r9mRmCLtLV7wGd
pbWzq35v6MvX3KqUfcKWyWJHT/yZjwgDMYFdsClIbeaubFGAsESh8Ba3k3vN
bWKmkPAsjpDmV8jd6qKrh0/4Jq+wbbhSrgNssGs2PnkXrY0mVtQtnLPL2Xpn
RScwLKL1wqthXJU6aP61pECNhiIbXjnLeahknqhM6zbty8JCzVD6FSaPZaN2
mSqDtyQpDeb667AXIWqw+rklE62MC2BIeFrv955LSBFN0wBrXX3ej4dJtHg5
wm8TcF0g3yvbnVjvAzH+Tq3HNItE5Ltivlq+uSUOiZ4ycCT5TZ384ZRKyXvU
r1eIF9g7KMzXLWdMtU0DuNSUVM/RPrIbLTfzNYgovLA9PwnKcdpN/rzZqgRj
1DOW5xx8eZD0u118FU72avPZbenXgiBUxTJTEwIom1+nux5roqDAeFkqYz6N
baQepxvAPp6NTvK4d3G0+K545q4yjgsymdEdKL5WdygHTiKAlithbX/2PGh4
CaBmllrS4UTe3E6+nlYKXqL2YBEFYSuCWxvlUkzTZmcuoJ/zTTvlw8l3uLBo
Dy+H6lf3YDOEQb42YCuisHp6mS3iWEVFESfEyTN5Al/WLjjLo/glEILe37tS
YeX5ZQZjzX/Rg8huLv9n+29ITI34RLmiTEXjs/K6UMVUPHD5dCwnQeHYTnZI
4m6mjO8nSh51dGzpldWpsrD8tmVF8kBoG0mCoI6ylbvEsHNfT5uD0ORP6ctd
fwqopyfimEwGlOeQZwu9UuQUQh6TF+2UBmFNwZgbFfr9tR4wQddaswqdwgQz
LAyEyhuh2A1i/AvIzSQvyYbqYmjAYaIZDV1kfRaFOAci8/PuwQStrk6eP6bu
mh37gCHPD6gTo9YSSwH0Zzz8vqUyW3jhOVesKifbUYemBSBFCqSvwzpCcWLq
VJMVWckpopUFiWy5/pylAIeM6rMFOlxPUbE10OliwDJAxmmDYaKtVGl3bnyT
uX5wdYPnDyEi0lmyydO/unWrNny9Ov6cZn9qkl0JVTFifg/lksMp/3LVGQJO
wRJK73i7u6f8xhKOUpl81zybsFcwp0RQ0q0oKd5NNlKFx85+QMx4CqhEMCwa
E6h5Os/9fWhpWx08z3TEsFc4pHiB/gFS4pXd+skyzJwMmq0+qdgfX36NB2VD
4m+GaFye8jOarz7hBzsPBOYYT5eUhI7+c7zWNToFTtXoOfnHnZScQBCEHMD5
h6vl9DQM2yEEOrLF9JaHhRTDy9YaMqDeKFkCtq+DpRTHw+HaLituK02SCWr5
eKo2EVs2Am5imkUIRzKpZXNdVmzQrGBy3DqJzCFfl5g+1MecLf7SIzRUII9S
wvAyay5eq+qZXoLRsLOaKTwbRiLI2vmP5+aoEya8xb0mQ7ahOeWrqDc75GMB
viyv1iJyEAa1GygWYJmASQs4d5xi6gx16zA5XEQ4BFzmTEl7A/vB96JEmYGi
jPK3lAtUeUkNfLLxrakRx++FhMbrfRpz4CCJjq/gsS8t+PDIkojjDHqaV42P
3t6albAj6Te8GBz1V/2unn5DP4sF6sUoK9dMl6rSg9gA30H8+Bmnd5ypf8lK
ex3SBldH0DV9tuKaI094Uqd//dS5Er1QRNRdyR22Qps73LMHhDl9ZbvIr1XX
kmlKk47tWEpgjVX/H4mOLoDp9QnpIWB6QRgg1abS4WJ8fevhwTSMBjWPKKpF
n2XtmY2SQmpn1lBf5Z7a3M0stAYH48j11CVh1FahUYiMXjOZFUnpIx6pS9hR
YoUKKQdAodnn9nKS8Da8utnJd20ETGm45ES/73cyHYjblAMVfhF5NT1erw0/
t4FKgQvwM6GBZbprSAyieBfZjqgmYxjvaxjW1b/H7uHEPptoS5ycpJ9h8YAq
bFLUJ9Y4l/sw9RzYVlXGNuWoqJbLDfEnFbAwWgVRSOg76yUq7DRa4HIicPdJ
z+ryUbUwQVpSWttzcbyvLjgegS4dKzd5sErLfbs1jhqMPZcKZp7Dxk7Xg+9e
kIn0+Gw245V5GwIJNK+6LI2Oi5qnczwEOVzVsb6f+lJPeVbTFxMnTZcHeDLl
RYpEaAo1eIm7OOR9v7we7AjrJfB6sGhPEdFB+fN2oJq8aQAmiBrg+nv5x5mU
prAW9uQ+QFERp4l4Sbg7FDFBcKVNC/JvZ+jGtATNeIQjUzZkpUUdtBxO6y38
FThTgAJIyIL00g5UIdcD9NdDg5+jxsZ11Gw2ptLuI97/zSVz2zAhVWYks/IK
YW4VQRBZQegOZcDFSRTsYjg5pklzcZYEoKoRLio36pwh4qWCyhIeoAj5Ce55
NBoiCkroG7gYn8N0Y46RaZckPE2SKLHs7A3epFX5g6i/xjhhIbKz7wGAHkQq
H3ud0LXIG0iZG8U3xZSUpAhc91SKLssS0AcvVRPThCL03lD4svsMCScngIXh
aLQS/xgmrhxMF7VDGRCwPqrqamT+W9ZHWHeqj19D6KpuvW/1b5Zb8isr4s2T
UmifbOgkc+qW8U5jQpoOOJxXSyafXWyeefR4rRcn7gANwmLAD0uNUSFzp5TV
8YqxHL8p2xueR8tERqL7S9F1plI+Tl3ndDK9tTaBD5Cp6t2ydliJnJCEYL08
HEm/vTvjE7s7e4/JQSo5kZAwF1cXjjq7Qgt27XTFnuTgQKHVxJ/4cqPn20DM
BvigBjif0DIqdF6L6GSwU3U21+KwoGeM4fEeTp87NgoPrQoHhvjouXaH41Af
V1dqpZdanXsFsKjs8W+xcVF8F3+IB7/hCUXcGoUzqIv3YXNWVNy9MNVfDD6K
j3KwFTBP7q9y2twnGMrYRi33xG78MjiUxqrGfVsU034DaVos8R4k80HjVFd3
KyCsHwfpIhL8qEMgp3GygmkSScqI7Hdvrhq5jzyzXqbgCAVZzqdYsaGuXUU5
XhlM5/t/K+NtwS66KRtc0t1cBIKu84TuO9a7grLR6tQu+GHxhbalmQWf9e4N
Ab3QnjeXAxOxO6Rl7T0T08VJHFOKxWX0BfpFg36Q4YOkfRSM5LRABDq1HMT8
ecz9ii0JbgFRzIJVSSH+k1ehQf6Ztemq1Fs935csilkfAPwbugEhBBwLTb7H
wJ+ktOKczqaKyhEAPBqkyvOGN124Fpm+H1F4zQBU9JgcKYjP5LOg4BiZJuQp
sh6UDuHxdAxskW4TLKP/n5izoFfLVumsOyvhqDgD7p574VabKes3BADLMuhS
vSynDAoWmRQsqBbjbwt9GV1E0o7os3pGclFjoORP+c0mACe+bxVkDBfrE+0k
QZduVkm/8vWGJKyk3IsaYDeRNx/pu2euQPjI6U03+4lZoruQo8qlhsKmnQap
uxuEzmCeUICIwfg7gKMh5b2cFQEMBa8S+iiU6ZNE9XDJ6LompnitYF/NU02y
4e+M4Th58CO4YZW/3LjYeZmGzdfv7ysysBU0D4kTOXMIoXSWbBLKeZRaGgxi
3fqf6zaNFjk8uuJtiUDc1/Q6iKrkKloC/Eur

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzcTIqXLIzG4G3IcAEyrcEQMrQW+QzNrsyY1QLpkU5fZfNCxzyv4Fx6mGXBlVLO5qH2e2oHFeEL/b75xiAZtvhm/Dxs6Fy/SxnPt9IC3RMWlvUuRNxcNnmjbR+ZMo47WxLtVqonl8cHX3q0Om19OW8HeMgAlXCVSXe8NO6dtgV/RV0B6Gr7ieVOziFYAeFS02wST/4Dj+wmeVKQGbLpJX8UcVJQlMiV6BMdesDucjJwete438hOSJzEzRtNVlrI2rdSH8nXgn1dxMVRR5ztYW8IXB3UH+3DgDRvakqcQnJdkw3x+ePz1TKkEAvgCR8Zdaby4kn5XnoUuILG0QHCE6bQT9xzsZguiwtj2ieFsNWlqhyb5rVEiKjnVIGbfwPmlIfswhU1BFon5DQ9Aby0fv+aSililQuvXHvoKQeKfBWgP80pQuCV/rIbLIsgMIUJzyBuRpzP2lRT7mpq+F/5fFOMiv3qqwbKUaAH3MK0pUsKKIgSJGkTmfBwP7ULj3UwSnZw9VTDTU3ESXkZFpx0qp39AoSCebjrBG21Jw8NcluCjNeXbPl6BVM2lu8tJ67enkzC89Hu/OhB3qJwiIWotyr+euCwtA4W8Cm1v1JjuqJEv5kB0WAhbNR1CpK/y4UeoMLM7zMsNNaT8YdgKxP4MD6ed/Kwk4UKLjPXJcjSH+5PuwTvMXCHUmw3epRHcT6W2S4NFRH1x62C5rI4c0LA+FDMukq27ot44J8TP1H5Ju6gBvJOVZ4mzThF32Zs577iGOwxQKAyNFl2MpvbjV6TgHVD5"
`endif