// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ifRxZzAobNJxxMWPZobGaKtJNDtjY+iYBrs54kymrTSXJ/vme0NvIPsVaBCm
zI1MCoJiG9pbHxbgQ2HlSOEC/MnJBCLkiDrZ54gVrc756gcsN3IFxb/lI9gs
kdho5azZhO3H9X4dI/eDaNY6ChO4n0Txrq6iwQpVOor8MkIJytAg/FtbJH+J
6DbShC2hiZvPAA7jjOqH9/9ihxIfw1oNZOg3T6pe5BueQ1dJ4WAdbuXPNDEg
br45tuonkNimu3WrMRMx3E+ksDU0awyLTpQyx/nicjON6DrTeKGK2XQxqGp5
eThn+HxLoYHAL9zB2QsfqUvAeWnyaEhzdckmPgsN5A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
irrJlSaOmOET40XZ3AeBbQbL17QovW6a50cumJ7Z+FqBXDda5Tz4G43e1lVV
UaaejfFu2QDarFKIkn8oxHVXtK4bggudWmIvf3duyUWHa0CtJy63IWnphwGd
DVjndoR5FA8dgY4znY48UTokbqPNReepxynquaKs4nSHXhEz3dPEqW2g9VNT
mcrae4E/94zfjVFv+/eMd6WjHzj2eP5iUsvSCYo+p65RMsQIHlvj5Qz+ENo2
3d2gYx59wHP4cN2QA2IO48JHAf1hbl4DXRsS/NT2nsfEhVJ+2+UuyV/01fW2
sBmUXa3BS384VS5ZU/ZFH5EYOvXCmxsema5m2U4Acg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PHvVAPA9GXFGi29acF/ZNMHV76q2c4Hxs3YG6BWigu6ZMobaFQNbXvPnwwuX
2tLDSB7tD9z/IXvdxd1G3DTteYYH+TgYCvMx5ocVkYsfarI2Me2AoK0qNSrV
3TPz9FMV/Q+jnUsNCfR+Jv2FnVGajH+QToaIqynSmRrfpuFxll2WNm9HYCOs
jgyVRjP0LMvH2pLa/zJjbdvKEo2/uecWMbEXWEPEbu1d0gVzqQ5N7NuGwYsa
9ydDEImFtnkePgn9UAZQvuCqUTyfw/kBk5mSkOmhXiVn8CoStaCjYYXZS8hS
dkWQdr5d/EPZSJnBiACOQ/FswQDqJEaPDwNlPABZlg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gbBQ90ZeQnPUQFVb+Uv50t7ouPZosXAp85AsuDxuBCYt3uZpznUBNoNPnaAk
pjQ5Nu9R8TBnZiS+gVSKgfqT33+OL00xT2mF9UADeNadAD2zf/b2AGgyq5eY
VBN0zkIn8PssZhEqS8GCIi1N2VQnESAwuZLnP9acZa4Q0BjZwEU+UkTFRC9O
hWP9XlBl9g89XJ2m+5lh6/6t3SUZZawAwA36ValVkHlT4JB4eiH+ALtighyI
ngjgBp9aZ20uCyoX5f+sL8rHI9lCfeTURnQhCAjUUidi83DIvIf/ZyieuU8N
dTGV8gvH+TNne+D/s2lmDMxVpgLq7e3XYx6kKmfXEw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S3gOIOICB+JxFAB4ZRyx/xoyK5KMRlRzPYSVRRPNB4aBYBlKGcPQn/SzU63Q
QYBV+wgpTDbeGAIJCOkPO1ksW2j5iY5bIrf69wiV3iyhqwHuogzduHivIGMp
GLZLIYHvtD13Rlht73/Hn8Bn48u+TVtfAwDQ+FlVFurzyR/a2nU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aKiU77YS0TjYdw8BX+LexTs7/CuPsTLiBKtrdP/b9y7Abz/P/WUSGjogQdtE
7YWZ/SCnp+rGWST7gw0sE9dMoT62K593M5kysSwMWn4rjWZymTaKTkn78rEM
CSatHPQqU7QUVgANkeFx+ssCKkyQ5icdMEG8qhFWGbfvApF1+Q/6JknJlfpk
liHarkvxSqkvUl2HEYw50p5fdHn7+MNnW+E5BSY9RA1hk7qD2T8Y8VpPlhXC
L9ncSKUyCaYbph0uZLztgDoFBOMM/8E8DHrivej0pGz/054Oh0zsEZ/+nFFu
ea1C6+FuzyUh8jydFRnAuM8xqEKJnKLGs7511KIkP3aBxDBwRNfe8RkmiF8W
OLuYUDZa6/dAxysDkZEUAmQqRZrC/UrZxpPCBbj1EyPA1ZUSy0dqBOrcNkzD
tD/geX9lxbvUJ4IKqcp4i2MFs/+WZOZKXGSj+T1uyEcr6QMmbc53EgaoyRYo
RzAgH1TzhBXoHC7HK3w7Io2mUv740zjE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IKoRo340BJ5C8bK00IWL7/RU1Wf45WJVSt3oVYS0Dh4E3PU831HRZZ6Zomyc
M+MnSf4mfIn2tqwdEk8ZY20Pu0rDAqfnnvyeJptIDjR4PwRSvu2UBLB6LKRf
oK5h8J31QOC5FWHaafQKCIjVptrczZIMGgMOaVUXGuBvxRIQo/8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FE4qMIj8RU9L1Ne3YZnuVK5ijg25+ns9NWxh6l9oPq+Rk5HV5BytaKUG6FsA
20m+zRau+1dmGcyMTHF30ILtK97OruVwms/OREJDW9xjMJz7LzW3ZG8YYYZk
k0TAqMWpWYsxp5Fe/+LSXiX1gB2qhQyCbLisvhyqxl3CDZyOZCg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4640)
`pragma protect data_block
9A4G8QEU9NMsQ9fqK3XgM2TI5d86Slm0JurRO3Pd0CANufwsOV1u08+M8mGh
1XUc/jj4VaCcalGeHy6Xv33Fk5cN3jaOtlAW6PDI17VVyaOXsppvxBT0thqT
oHMu25P19JCG/zMrI71XiXjlXLzW9xVDpn52BwvYZhkuebkZUOwqAlnB93pA
/uImtiEp3b3Hz9W31BjLSEGzKYXw3xBspTggAWtfS9XqyzydwvIti7A7Gx5G
+1/r4J2V2VsFrRwb43Gta9pXseg1ypLm0A5uSed0k1YAbs9gItdSUxJ31/c9
qT/N3bhZVoF5U+ByipYhwW7oIgrf1y5wMc2ohCTQwephI0+bUnMvsgL1GcSW
/TuCxfo5CWJI1KpYCn2GIt5N5yW1Dg5mAtKYh4kZllkuZKmCe14qeYAjxbx9
o2AS1l5KfZ+npfsA5xmTebea+xkAN4oshU0bozbDApWt6ufJPE5uQvOPA9K3
b0Nnnxffq6L5Q4+dM1/9o7UWLp45aEZTmpmoVcjFF5wlRhGmUlacoe/DX7Yu
CAnAgr88SKOHVV1VlWs7NuAxkNSebHgxyvHkM+OM9280r/8T4ptweK/SkQ8a
qUJHITM4CUJWpqldfURB8CUP5JBGCU1By/LfV3BjJqFScZWT6XuSl/3xo9sd
pIvbfUnHyP+XGArtQhg3eCwDpAJCue7S+1v60JKsxAQED6vXK6sYfuVzUjlU
sDUCYEToH+lUK5h9Nf/oVrXnrmbmDb+/1lNB/p8dXxpkbapNRUVpkkdbr+Pg
B3R8c39KN3QYb/CZ46DGtnu2vm3P7/t0TB7InYrV/1m4z/5+RfvRxXpgPIVT
Ambe3iN8WawI977RnN5NMM6Kwqph6sLn0m84FNSRNp8EwUOiiTQ+tMSwztdm
OGiYgbEjV1h5zI59ULgtJZuIrLzaThaxF7/qWAd/RU1LqVuV5TkGSy4od79H
RswMDD7ESOCqLiDArJ2Evf/HrRna8AfdoN9TrjIPWVzbKrVtIggnB9n9xtMz
73JNi+9o+wRPCZ1wiVw6AgD3MVlqX45aHFPggzvu+UMyD+gW02f7au4NMGIf
5+KSl9wJsl9BUNs5KHJHoFzy31ZazOrsFD1gOuyX547ypcWc+8wcEeOWaRMg
zBKT0f9aMs+CnGUhkAy/c6u/Nr8F5wmr7s4GSf3obwPLVGL3UtTj9Y/389Om
ssZYqe37nKKQ+AuHuylPqYy864R76KlLAib4L1pb81TdkvQrlQIdVmy6qoww
vWKX7vTaz8RHEuRwmPyHn6yak4yQTazYjzTLXGr8KtIRWIeUKIHkWdNkh5wh
MwX0gHNoxvOCMkNVWUFx2iWj5/Kr8RpSBHTQf+2W69/BP1CG/jWxX9Cznj01
jFDpgyBsmpqAhRpRKZhmIBC1LEY9FwF29b4EsJWvSgGpTdhZDCZL2ciXIF6K
mS+Xx7fY1Ng4dFa+vHgN1XasJD8sd4Hfr2PivpWWEki27wazQWaNfT4jHLTO
tl+jnWcj6zmsqWN8tmo24r/ijbBVok2DflY7fYLUDze3f82DQmloVzIaYdsX
0S+UrtKWom/Xra6ZVvQq6phNGh3XYVumdvxCjxK0xDnV0ASWTupWY3pwpSz0
mo9Wqqv1PND4uPCxL4z5cyDQ9VkIi8Mx3xNnN6WkXeeqDhO+k4K4Z+Jej0Kd
wTs0oLbUigK0N5oQP2+koC2CliZLeCpY7rdGGoLVdacN1W3OhUzXzsPZNOKu
FEU2vVCdmzj/2vkLjCK6aiFN0A2TTKjKsx/UaJvy2PSlJmwYh4lVO4/wdzcn
OODZKT9v+pp9zx0+9hs6hJO2UQP05YI2o5pASIYJhhHDhvhzbWXK5hz/N1yy
GPjYyPx2mjcVP+gdZvH8FhIO+tdsK8xZCrG/ne2H9HVF7vdGjxOqi8PFimzJ
iR2XiPfyPHe21D8796TbmIWS50kWA9gyG2mFiZpMZbR1doeIS69ALl4S1T6w
Rfl2LmHqVEJjCgvDm+yFMmzwUEYoD3/NqvHEZk6X3wvobdB4we5oRVfW0fQo
JT+5niy/IsKobYCYKzcdlXhPwVb2R/CbO73fxK6XiEVBZ4InnEDL8sXFbCay
FdWcX2j4dVgTBzdjtc9xaz4oqQIaGu8K/lS8oUKjAawCXY3qg3koi+X8uGUM
P4xnvm0uw282F5kIRZrQYtfKLuAcKl1jfpjxOveDA2ncsXuf5F47tpFp8Jdp
j40TvUX0MGIHeDLUX+UIoEKKwAP0LuDOLmKDLDGmnqhMn4BST5edaFsbfpjp
KnPL7EKrSCTw5ImY1ElcPrrmPaCpjj/a5mdRe+J8TL+nrpw/6UqkxgdBKGef
BeOpWgWiUmDDXEKjy+tebU37CoJ6XIJB+3zQpCyWh2m3fS5Dj8K8C5SMd+9e
toqUcvHqOhS8/k6QZu2+1sJ0A5yEJ6n87K5GN0GHn0XOcycm6fodXEbmXntK
xfukypqQP2IyuotAJ9FTvznQnvwR7vlSCBRwCMdPjCJvwhRA2AezAn9UzHYc
ebRBO0tNms24HJlihdR/0OHZg5h5Q1OdXce9X5SMU0UkJfcOA0R3yTllwosB
FvciyPbG0X8g/o2BgEOz/fXn9B1zTXF3DKUKsGeLxC8vvBsJ8QX0KSv/YX6w
U26oVMOv49nV3IiUL20fHeMAp2BBaQKoUPJbBD5cjMKGqLjsBzOiEwyAHYul
eLMCcKEyJBQhVZ42CgO9KLTa1TGFe8F4MnIgm895E0J11HCWklpCWp4VjRx0
XVfBDrK5E5Bwt6DfsqOu6DaMFOXDj1tyygxRS21ZsPktxhpsKODLjV3uBdPT
7HfpyERiCQwnsOk6Z9A19siomqojkTP8gzJ3YVLe3O7Oom/QPoCWsS0EOgs0
ER7dPTvyYaEFdbsLy5OkwqY+MrRP+kkEwm0LI2RYi9OxyANxDpqNAGWbuiTf
Ud4kIQPvKZAZNGBIu6w3BxOXqF15ILW5V6Lp7ILa4CmezsXzp2+tUJr8lWO1
iV3vda0ewTJBA+xLzBUsdf+SYON2EgL9GSn6RvCTZCRzgD8Y9fBuE4f5DZzx
SiunJjlgD0e+Q9kgmhDpQLny4o29e5JoAOw9ebtE0CmYAPMwMZOsA6eOsDid
rzXGZDpwlkKmJJKjxi/9aeZ69UBzjqCudm4GWMr7XYNTEncVXoPlrYQiZ5v/
MjZCf0hrNlOuyyOca/KgJdJsEdQgEEfGPDVZioQ9IzxRL46VClANtMN8aADk
EzpWsxuqMqv5Oc/N8f7Kb8FVjMNmm5MpAAyxvAhzQ0nUinX9HRiZD1qBs4ie
+ua0iPECnU+S0GAvCOid/2537E7DokQERpBej/SgJmQZCOWizSMcH0wW0Ao1
x8lXQlmh2YSUi/fnNh2Hw092z5W2GNqTzWMWRZ2D1xm/ggzENN9fiiOB6eUj
GonyHNZsZ7MB7qArYbuS259c5Uny8egjd751BIwaE2F93iHg3VLSGbKEli1W
v71OExvEt7Ra6R5a7VJkwJVoyx/uc6gk+dfy/bVsFMuefVDlnXPjIso40A3E
6t2oxaESGaz7y+sA/qqUxRmcCxMpd2GPpodKBFgdae86ve6Ay58qFzJ4BLRS
iAOtbl1phNCe1zIAmsnyLv3lTqG5x93nJa1MR8tx7/P/mTC5NjD6cSRI3mBY
9eMBEAfP/ymkFirsak75KR6cbSBL4LonkyaKq85nS8TDYSOitulBpkdxpyN0
LS6Zu4Kg7Up83lj6gWy16rqh0SXKRuOl/63UlMiE9rfkTgdtWv0y4ffhDhRu
fOFrAkiBNZBjC1lyDmF0MPGR7gMwbEQjO2nxrlU0kBQ2rWHIRS1ZBueSmU/o
SyVFsgD1RPxpnmtUIjGrB6sPCvN5UuKHveNnELErsvr9pkph3Fqxu7TCI809
JEXZMxhSbvLjfLaD42fPlKkZS51XwWEaZrJrhDDwORgqDr6/JhszDwTIyy4a
VHT+JeGh62dBwh0/p2LNMDMapP3ksqD/FB6R/B4M2Mo7bHegP2brh5WIS1G7
arcQ1HE5iu6PnDTlKNkm67jXQ9FSQaxw2Md7vVBBNHmguci2s64hrtW4QTU6
Z+BCRV5bSrR4SbgD2tc2Lr7C65Ziovp3HHHLir40YE2AZHjrEcCyQsu/otRm
cEYzCR9t0YIS3K1Ta8uFOTGLtUbhDZM9/EtAnPuSVzVNVGLvJ3gkJC09BSqj
pvho898jF76WAee2I4ogc9gdPasbzQ8mH961mD9VmyQm+Fdd7C6vm/5EY84h
pHJJnS9nBcTxDmBsjbBftycwdF37mYdHXCkNzK45jfGxOXwiw7/sDMch3hxZ
KTgWmQKOJGeA28x2kGsAjp8qvnYcuF3ekx/xm69Gx7lnX/d0JZTenXGOKh/f
anfwPV7VgDVS4EnUhlgA3mOY3nIfqMNN6UuGu6D+vwMVzlnc6d3rc3fZesgR
Y64l2KeH4KOrzYFjZuuRyVrVZTCsGYF098FiI1iEEpa5P3M5bciGbDR+SkxN
wrDz3R+81hNhbdN5rJa+Ryxa53kD0GlEyLgFY5i5w1Xbd7SKs2ha5xxSssXk
jO/xC/oiOTdq/bCRlFfwy5hPI0Xoo8f0XKHsJac9t2B2kq5wF9S06khrA90G
WIPzKOR6QOGfIpCFjAQTY1v/Iz7ERiv/z00UCJB6ibIImqTrMqY/9kip7BGk
o7lFSHy0Kw7MktATgd0RhkLqD2/fy+vFNsYa0R6kryJk/q6kQ4AKLtyHHw/P
WjOi+JG5ouptiagatkXDmm4JtJ5JCYfgh7LFrBlqT6Wz8Sn6GTZWKYkDEhJN
+MTdVOntgDf6MiEuJLbwK2cZFdYLXQufC2dJewsuXnTbOEqAINO6VLYH1Ymp
7jqgxu+13EYreqn+14xgZovR9wGU/6LS3Ykdw47SO29wBQirGkyf9/9m0eGs
/CaUZxt40NUr46WmgMix0z7EdVe+9hwtHG+dWVuUCmlzpUeu0rjL+w2FaVjL
wsBIUveg5f9BNf72acBDik1uiH7qDuqkZs8mfEZvOg0JPQFD07RVMx26uBRn
02kcoKuJZMJ0gNOggu5H2QkgA0esa85GCVAuI8fcTnC0ZL72n2LjHfmqWKrM
aUNkgdmc99ahKxCn3oQ5wno+uqrow4MdbRnTHNfDXQ8kUdBtZJ9ECDxAcaXE
mIQRlDDSuvjC7y8UtXlcj8yztBcg1d4kW0YSg7vUV9TxK6uLXy9DVdXpR1yu
8QXzBT08Eu8RqJ9MMPCKJ07VDAnnffT2haHHd5/7+c5tV2zCt17zffOFcIWN
ELnjuvJXQtQLOFF+VfUy0lhDLZjCEWzVK/WDAPWSir6V9bSzbrAfQMFg0VVz
ZKwvJElD8tRppd7HEiShvSstlHPwWItEErS8dUCpbba3sPpucURwEYillm+B
Y8zYr4fM9w2VnbuacGCMJzeCltOyQS50O6+zvhouoo44ewTMT0bZbyQ+ELHA
M4YhNxD61VPXmMWe763CKMndbPBoZs+sWYDyInb2d1gZc0lf4HLB3jQoGR+S
qGh3ULgYfG5OO0L75wsnWSnfM8iuPLd4oUtsv0vZKukjn55mfNAt37AUkGUk
GSIgBbT9MawDbN0G/eFKJXndEK6GsuC2KPT7/A6Z9nMTuDlePPnyIU2xwQjN
cr22TAhVTihD6SlqFw3KvNgIvM9bchqLTSTBUycb4rT8wgBz5SB0PIVXGwDw
/dPUdPFccR0EE+XcOBJlXkEFU5YUpZax1Teysy8TvQewAb6SOBAd5V1moeXH
7Sm50STRK3tLz95gbj6BKhW2DFNGBQHGjAUYAXnOvjK/meNr/HNUwr04oB+r
r473a6IjihXVXC5sYsJ7/kmAo+TL9Qeb5VaoMfOE45KmcmUQJaFIgU9rqEr8
ghJyuvaGWz+vYXpBwr2S+mjGebNnKDiXoi76nwq5TIBr0N9IVBYBHDYiIumf
fZ7qp+g0nIdo6WpIF5fT4t/ibGFKLnZkWJ0kJIXT3xkCcawjBxr/QEyCF4b3
gMOSbAlEc5FNd5PIzESKjviqgPTTg9uFA0ufK1S0VfIc61NbW+cBWxTgroM1
enju2GyTxT5z536qMMmIYWWthqr/nLrMUIjzydA9INKvzUDVnS1XhhkH1Xrn
N+T3/9EEySmiIWD1NvdJQRI7e0R5DGcemeGTjSS349jx94aCcp3Bgrd65tSe
3ySX/xY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJPh8s9pVC9AHA/lm+sdmTKNfI1G2iizWGnsOPe8RIxUm7Ildd4tU2TPUnkD3OneL0OOh7pggbGEbOOVnM4wMawwGJuHrFCU4V/3u6MoyVQPfsvYGSFkRDbaKdno5RM3FWScRMgwK/c57rzuND17SwoEq03/coYOmjAxFBBynbWKDuGdpM94qe7QIa2unDDfwiUsWzHz0x1izBXk224YZrFwR/YS+fHIytfZD4Iv/FTJ4Ac9QkSIKlTcEQIoiqybnDsMpXc8PzDCdH3dzMLAGPYg9T7aPsfNh8UY/5HOvZmzEs7UptW8TfwSfsH9aOzRw7nIciWPUr1wkRwWB6fM6PYKnTMqa5KE8ddFmzzRlJ3PpJOWQLawUSzTsaY5vJkOHQIgO0uXsPETKjGOepNUDvYIr0iEkUNzME+UD84dGat44+JXfE16VIXPMVhuDhCAJ1keN4Vz29noRXCgx7Te7zSASukQEh7C0CbXWVuNVQGRKi8wbpCTjfkpTGXHCpnusCkD3np5gMYgnfN+dKMsyg3Klgnrw2F2YVTSffzinF2Hk064OyAhfx0xPl6BDhfnPtF59K1DYTo8AJPwPbU1d020439qJIM5THLPfQB9HRsO8TQ0dK64KZnCuxe1oIOrVqzLQsLHONX+Jv6RDXumSFQo0KNaDsMXA4JhhKiHWn8gaPVBVrtnEF30BGF5sXyX60B591Naj2RGzd+T0N2onsPZ/Wth2ft1FsHSSYcBoIuHEMrTmQwDnrX+PHb5arBREgnfYQWXF195YRI/jSUn2M/"
`endif