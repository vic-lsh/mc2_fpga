// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cJsZuUe9H5HYMx+SnB6gU4vOT2yO0ld/yEcWaE/+dm9uova7QW1keqhcdEYL
nWDvJjOvKBqeZhIfg4hNADaiSiMXkyBlYDc3eiNfzt/+2Z38NWFM2GFwz/Je
s6n8sOswjWR2dTdXEFuVF6khlm2/J4MiCQskV/Sj7QgpHZa3fSYjGG4EOMDT
tmRlhKV7YXexLGh8M56YvDLTDJttbgublIGGME4a8CJHEagtXxfWkEKTi0tV
KSDIqo8aYXlrUBU++E6yh8dipg0kTCrZK/b+N8biB/MTH9NiJocvRkstCjs6
YWN77oGCKzgX/gxsXKpc72rUQmERSQD4LGgnpqTXWQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I6O2AF/VQXhKIxmyUkM8MFCBlN0dH2FzzrqhMhRQJ948nm36Dzt6+Tixajw6
7oDQ+IP8rdTHQ6h67pinjN6oFitiLbLDN0/u1xYElIVKiYkfYrEBdI160iyb
I0sPeGjXqZf+Vi4EAGy1qHDDR8BjFOe67HIkLqyv1MpoZXX9rbQNFkdnJvSb
G/MPgI9IFMG7kdCN1tlHmyBOvzPfGeHoNmdCzssspjErp+1/p2uUQKrktfVC
ZMr1GcxbrGVv384YZ+fVexuQARj+fBpFQqd23ISfj0yalesNdyGgNfvkY6PK
5xX74JAQ85iKEWDTFwWz10H7ujFMCp0AQXCRI3IpiA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eBPrTIn3rVbs7ZPE2FPGcdmWsSomb5QGpMCg/VH6ut6cUc5BIkhZj9YMSUZa
CAdCkQ2O5HWOEvrEPB0V/E++W5TW6XtiBQ4wK/5aMn00xs6/OwpKndGuVTYB
q5G2qDIrK+3MrDcEtRhXyNSDVzcBYLTWDyfXhThdaVrcwJ5aclbADpcEXi8a
IOzmoZ1k3CeqdERUZh2ufjQFLDVgCQjkMHOp7cTe2pw5f+QuPGaCkGqsczGe
LksMMH6ZOmhHU49cOOTaNHz75N4ks/eH+5AIvYkwmGoSla3AK9vYgADJxsGD
f+Dc96ACWBKyDEtYlxoQ9MYc1hDspPccF+76++ZUYQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oUOz50mWqLPs4NyM5vepd3hbTiKoWBN4EHgMiSKASHrNdotJYYVBL60cBn6g
/eLmiqMJ+JLLaIhi+jrXgSDpRYkWAlbfUYAMVDafWEmeuuPDuCwzrjElGnLL
/8venKGgQeRU8K5xobOEL3TwqMWMiwgvYH749dLFNH2HG4/3mRJFCd/Xb1EH
4QgSZLQKIVGUGYrapMnxwQrHFN1Lr8tzQRGCf7+kljyhy5Nw27QfFtkWPewb
jHzdM9ldmfNydmUFTtwECjkROB0B1J1aTgnZgmjcL9RD0aYqRWwaxvEnivCC
rQxYJ1BwqIMNsp7dCtuiLcLQQM1Pcs9x46U+hgkwGA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FB3aMvN9PyhXFTAS8ZhUMNON6Zphb+nrT+Xob0+S9oPs3TsMlBwLf3Wo0Q0r
zP64lzbXLt473MgLQl/EBtoMgrAPdXQoJ4wrjET32Yd7sD9U6uoDk/DaQTTW
E7bObFqeZ0gjDX/wguVIF7YVt89HsNha24v0xLet8+FEmjuZghQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ju6UUfESHy95DIYaB6FXHVbC5am3v+iS1eu1qDbz9tjYaOGGjHBJXiKOY+BP
uutJyPd5NlXIwyZt/W77xnKpA8C34/Hr5hHHb2y7b0OzEqdch1k3uYOVab0R
bHOs39J+joe6z51wL3UhtdDfRBILT+/LGf2UNbbcsf6z/qUPsSkDuEF7URY0
xtkgCXIsnMR2rqG0EOxqiJ2AlmpG4LohPbNmuTOhLfCou/wTgLr6nJJI6UyB
y7JyisBCDZxsE/Xnyl03JOEIWhGuoVsRQnLTxJ2FHJmrE71uabv7QbvX09DN
/uXZqhxQhyiwp1yTriGk8w8JQjxFgBJreJGXCsP4qZgrZGgwI3m1y/4zPMyr
JOU9tQpDzrPqY7lLI/pDWK4qXhsIwgyiz2C0axgSrhZNnlxnIgUloGnGfUI8
nXpqQ4UH50Y9/n9/Q9Oio8Rwex8n9/okOpts2cm60Rpjr5/Pcab0wJQIJutz
6bgeNU3t8nw8AQNNTjS7LxRXZOxzDEk4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oSSFs8MD3wYoeoz04qYLceZrgj/+dbPRnrKNBz67dgnWtI30TeLIc4GIKMqG
a2kS3HA6yDu1iw5UGJTCax6dF7CuXQQ6IoHpPuxql4Mv9KW8KzLDby5sf2/d
FhU/dXAAGcthYciloTq74l3hK2brO3aTh04dc6er0sy3/BZtC7U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Iv3iA5QWwUmvwUntU2IKO8s8vsg18ZoGzckZq1rsecW9XVY1ibSs/374Kcla
qMOpFhG+OyvOODsPuwbsTcMIpAt9VDC0iuAUfziH4r54oqHGuQv10TOFAt5N
5+31E4uGzSVLQaFlsSYB6Z/I0Pd2t7posVHbjFZQ4Q0zvqQw2Ss=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 5568)
`pragma protect data_block
WKIvgSVejGHXdEDM7UPctIkY31F1HGz6Em72AgPlm0YXok1Fafc14WR/vgEB
CQjBka2XKlVjQgY+f34gJ9hte3o2pRak/IxG3dawR11H2x4zL002fVi8JAVE
4YFDP14T7S53kgxITMvSHPqQXtI4rJRdYwhzxCCerpieYyJ0VDhbkv0gl+Rg
pW9+VJFBeSNVPOF8YzVm89BYyjdSX0YZ9C4Yvu3W/m+Lo2djKa3zEkACDBak
6ktxCeifTmuxiTFlPVUGbnUmLGHNtQHllcoHBxxEb+vJn0iC8w3Pd+EXmxew
IB3Tt3LL8RLArNYv6Rzqfahx1r0SBxX7JVKY38hMIdtQIRU/JLVcNf4Nz83W
4IZ2ifEYN0vS/y3/rM0HLE3/dJjlflQ7yY5zNz/D1W+JhPhoZ3ylk3s/kZSV
HjWkJ5PK5yCzb3J799MqxWIAGDWNHt9o4ahiXkcK2v6BpD2BfJUfetGgDG03
1tFqkXN1BIm1LQudPi98GtvN6sgqw0aRsbYIzM7if42qjRUSXG+4EVAbl6ex
tAI/THLmBliMGVjRjvEKRm+AJYA5tBLVf9S9IUY+adKS3DLO26dZZy5q8Aai
IRE+jKHMJSAJlc1Z6SCSDHweor/ge4CtebK4Iho4GVJ7N2IMq0xcqXZyKO1w
8FHCwNFew4K0gfkS4YOpa9I5W+dWLh64M6KC/DtcCigMTKJwVgTFUHduo+oI
3BKroD4OQGYNuWp3rXP7RwH8sMHagu6ggTj2HAsltKaSy47T78/zreyfJ9Jx
2s8wO8Um96ESXT2rs0GZOI4urDNW6zCKFrurI7UBbqsx738uRDLZwi2DZ0Gf
NE+qRcHula8AwhhZQ2/rOKwnmUuzX5oTVWqcHPYU/U5ZEXKjw8Wrk7AeTYou
fFXiUFkPKVBZVLWH45hc3WyUorrauKqSITZzZkURIKnFrfXjVWi8SyT4EnZ5
q8LXaM4CL7Y/q6wNuDs74wIi2/nDESTFqaEvs/0fs1SHZDKutS3+NiJHpZ2f
b32CrcMO7E68pCc/01PM8A0c+5+z9tYJhCz2S8IJEV//Ix1XdiGKaVU97y+p
/4XQz2b5DfD7i4hkGEJ5qi5RS7gwihm8mlEb3MQ8fHbSJgJPHPAadpEzKmrF
ckwS6tOfM/ohFfE8vfbfKlzUTYkID2qofVjLN1HxW7/DSJQEhP3ubkOvz3w3
GJ6/QJYMTqic1JaeG50F9eFzqWxYkYtTecgOklb5zvoheia7WEF+gblpBOPT
TD9p+54X/PZxFvqNTbSamTKPgqVe8+MK7S9NWlqFrxR0HjZuy+uIjo1tKUt3
h4fdy4MdBKe8XxoUyOq4eqSGX9lCJeobqAqqoy1wHBZCDXuJtiXZlDxQOvJC
RB5MJSEUB0s/yfhVrtViGlSEYACjqb1Y6hu68k55LaOkzt9m/YLJyaH9nkvr
KAI8yRyLpkrrOm4p+fqpJrHUxJ/rTriIViwMMc0ChMNqvHJM2qSEcXgKxsJr
6fP1/rFPI/bi63Xflj0lN+WBDYCuT6iNW2p3IUB3wBSDCSmPTRYVhipjCaSz
wEo9x+419BsfkQ5ZLbE6uvwcsFz9fOlz7QFY62YFkpQ+SVpu8SPuzaX8FObc
e0zItTre4NDsn+UgJYOkCJkdwm2yiSVgfB+Z+qGcurDnKLSANg7V3lhqxOUH
gQdMvGbgXM9JqAjDR6uT+vqwvoe4cC2gEBzvfky2iUKp8S5iugER02z6RJU+
aFyiqiADI7XH01Q0CCjonKSYg8Z/ZUM3Wz/vq8PnLQXrVecVl3ybyNeFfKxN
5tAM4o/CyEw3QNUZv5SzCnQ10lYRmahjDgk+5sNYn5N60tUFp1LeQVVMmMZh
isNGz9rs4KZ3IDZdnhBmsRinzGTIQDaSv+tNEagycTqDqTgFRUVi5pK7nsPx
jPMB3dgz4oCBQl3DTFg61yPJLyDZoxqUSpv8wHrSRwP8e/Ry3CbM88FRqk5G
X3YBzlVJQcVGJpjCSv+bZatoow7+rJOZBIQ0B8AtWwCGJ9CEVQqAoxGygFUa
WR3vz8GxYYMhWuQY0csN05Sj/aw7qjjRZbEiJw6P8X1AvUKJk6lkOOxS6dLz
RIrW2IlFFZIrT1DIv8Cdv+b2HWvRd/GWVLW8ncKAG+pEcs93zzk5uxH1MVfJ
w4A1+KWltalR4x3o0C7ca0kDkKchDwdltxBw6OQNhFSumjYMfhIA1EA6At5h
ZCEZWOtYZkvnVVLmBQ8dBB11EkqYRlS3SLfkkymzRVqvWEfXnrm1M4AnrA2x
D43DIuYle0ewBJfnPJx5Q8em/NnRu/ngnCmscnUoMdaSOz4shh6PI9u7vOOk
56mE2YeDCg6/z0qZ1hH44QVtArZy2nVkGBVCIuFHRb2Mp7duF9CH6gQ02DmA
N8jyqROjxu58VKvHG+mhL4eIHEtOf3UIPcpDUG1Ym6bG0sSIXWiJxX/cH+78
E4i57EHY+oK3ijJG8TvE1OnC3criX76inznCCGJBrDugapwwCFPiOn+WivwW
xMYdRNBj9ep4wVJXhJPNGwY8iQR5x9JBIZKyKLvNXOXO/MwKNnpPAi6xJvSh
ImKdxU3l7qUpRMSXEtdPsqJ0MQQH4/7MUpnen58/9kU74M1HoMKiHp82ZEUe
U1p7t1xkzAvVPhgwktH+i6UM9hceaH5OeZvmnJ0evtO3i1kVT9YS4K6yq1h2
y91TaT2bbKXIrRnTCu8FvIxCFgIFvAoTMeyioFc9MdunsgCXbq85QKfBGJFp
4p+KuzwylxCcmY8bum1/alpLvK+mPu+KN4wtxPN/8n4zigf85wSGYlSAWNwA
7CXB2g8ffK46Bpa/aFPSGf3Op5n9sX948NLDgPbxkczQ89PDXSFwf3Tp4NsV
KI1Uz9RlSvc2EKijq0BQAtkXhz3xea7q4lP88x/L858WxSCpgZWXGNFH0xTJ
XPMuFetB2yvV57MV/+xNoqtqFjyWnFFyJrOxyGM+wvnj5f/8qYp7LpxRbnzQ
GsViDlcI8LfDvT2uL2GFqhb5WYKcqMDCqjSSvrmit8Ubf+iY6g1ralhEiMxx
Ned/74r+rpDZswFh+oX5au8OXs3VrxfIvbNdVHUFz+tLEVo1FcupVUY1lvOV
twuF8rWhah84lYyaNfpjtkpFLi7I4NopCz7L6yyhKmlQPkxD1ro1dXj19PgU
kuKhSM+kBGoJHEsO65pDcVQ55Zwthxn4i6GPC2AQLbRC1FMZGM5+Upsvns/5
Y9eGVrBj8Amd7z8ZmZKfDJrOrETPcycUMDxw/hzTqm7Tab/0yioX9NPvq9OW
3pQ19BLGuyUZDAxVNTOyZgkjmWsBD6hUndrsoNo7rtqc34WT/cMjjlY0KFqH
H7vM0G7XHB+qvog5MS0v/wYaeVkGj4qMI20qmFOPPMUo1N8X1dt6Ab4OIREw
fTEikhGSnj0PgMagE6UcQ0yidjHH5DTbbuJYo8XGdIQ6ZJjaXxOSu9sFSKko
1FrJWatVU3hY33/Nh/pTbqRvdqO7dIDMiXZ+Bon7Nl+OqSvX20YEGOzUu2c3
AD1KdE4NtA/atciEOPrUNtk3EXXw1Pi147z/nJOkrA4ZkDowhdGAvkaAPRbP
W7NmcJyKn1+dddoNQ6ne70rN+Ii7fAungw7p761GkaTA1fXx1IBXr1BknRbt
y6xZMmTeFxMY0WPotIyXVQFZHvhaRlEXyZ5j/DTn802DFad8KnVdNh9G79aQ
zVikuLW/jVUG3eNpaNQxdc83XBaMRM+c+Zfq4r1q0X9xLrVZ4nZId35vlmKr
CcUqTTb/ugCQdirFR0c1eYQUnnKARYVYH9hOV9n/sh9SGcDRCGX5rpX6HhoN
L4fFhaa/uZanFneWR8H9vAQsxomwgz2L9QvqK6Gkpw8NkyBbHsisAPsTAaYt
2GzDRphYThZBe+zfLDaPjacCbo3DgfQ0ud5SsHMfZ7qRIz+f6XjUhOqQtSUF
Jn0UtZJSOPqWnf3fE7FDvfeWXgz3leZPXkbwiNtySgw1fgjrrnX90Q7VlY3B
Q+4lEw9sOk1yyiug4XqUn9vkx2p9FfrkAoVjxZFQSMs4jZQMO7rSY5RsjU0h
zhMs9BfAMTbbIqK/RilxZg75PfDXwjXK10ht7F3RGKdeoOvrtXWIqIPMhKKI
UPqvuSrR9iwefMxfPw4WXPT8Rh9mCsDmksv3kIHvQ7D3wyvJtQjHfONpou42
t0Ifu1Sj3B2tyJ/5IxCSWWwGy2kcIC4bmegw1aGEafL7fmZQHN9iVosdSQgc
GluOZlk/axE8aX2HT6AYX6zkejE/H4VrN9mAUUOwrpzpPlr9p5BylPbok/iT
tQnuu8apVxBFPAxVLMmnBwzNS3HRDIXNgq5WIIznDEM/58hSm4QAR22rKmZi
YAr9WpgXQPRobnOuC5POOjLGeh/al+w1jmwUrPGs0Z58l7b3Dpqmj26ttSN7
wthsttARxBYHub/Q5OShms6UFHISGexhAlVpGx9ucrN8ip9mWCc3vHfmhaPA
qAnSrJZf+eSpP21bmml/3S1h/6gQBbfbwAlp7sXuuxhfO7iu/DB0wlEIBsj7
wGxdfp3zNOh3xZburi8h0xRm1v4mE8X6BQgppfw49blT9XJ27CWRjyvFO0q6
BW7HWfzHVsE0fR7yj2BArEBUzJmUuTT4h5LCMvRsI216/dx3OwQbpaD4/9YM
cxlhnwttGfBh3Qpkgy/DJ05k15v1u6OziBt6UChfNEhTiiJ0tIskZgr4sCEw
smE8hlF4lEhfafuetFARkxFoel64XYTT6N5RQGo0Ejx1Gf5jFH4z4G9dCg/A
05IUz09lATmZhQEnkFXbCSSn3slRQMEzioQ9Izc6jumvDrRb7C+Fywx1nrLz
DxnLZKcBi+vjR04eXZ23i+90Z5jCVCvXwCcAaXAD4aNrtOAU2aTXW4Bq+9LQ
RQOctY4rCW0lGtPUWLlOX1dPT1YlsttDbOdli8k+fsB/oOe+fJa9bq8KR6Rn
Mf3eUjNJMBN4oKsIbJYhJ+g8N0osV7+URgwdTOxHxadzGMbACzIFZsuGMhIC
92kS7rIP4BMqvfOJWgtJTzkfy+83CYLkG3NGTTxvsbFuJ7QtuBbtY32moNwO
gc+PQXwTZzLSfCmEktTxJYmVaxE2g8h9lc1u75631H51RESafbxBXUqwyZhh
dOPR1hV8iaGvzpxwRe8wz9Ra7atDYgA9pr5U1n8W4FjQhYKav/4vsvfvspDt
gRn/WFcg1BhT/a3Y0ubwHnwPomnhG4nlplvLdtAiINmFGQwAJxBfUgzy//+B
bPH3tO5WpApvOsqHBfBXFUBj3RD/yS177K4HhMBOFBEGvKNzx4SnUquSxj5k
A0DemimlR8g6de3FxtXNqwAXrPT5m6z3TTUNGRmYRWw+AxELncZ0tZDlGylP
IlEFT6KCGjGxKbIzAOLGJ4Z14C+lr4URH9A3AIOR4xVfPiMsfpbF8UoA4Sgt
/3FRG5Yv4mwiQomkwQdkDbdE+sRkSlF4cXJtSmPkkH8wFiJWg/tfjn2Wvziv
XulYy6EkH7GlmmS019+M+X/B/kyjGhrl57dplW7odb08VCvDJV+OD0yKHchP
pYVnAT71GHSKO8+HiaMKy6aEUmqRmPNLWQ3K64//nbJhWyO616Ui7H8Ok5tx
MCbsQVH82kcW/BkahzN2LXRsXpWQ7XTbwxoIY+2s2BlsivQ5zZpRn9Vc5PQm
aTi6YCGY6R8tIYG4FBlnndRk7oldMfxopak/3ZDm9XlGVc1pj6pPfThWGoN1
U3/aed4hryKDqxWEwMqz1fYKV5+XmaB1tjFcbhstrW5cT668HsWj+6nU9LOt
WzSLmsc8cez8YAgku+RB+WnHVyLFsZVpExL0/6tv7ArPUPA5iJon2tOKmGhr
gdKY53pAkIBYVh4PYW4bHzcPE4J9PrnB3ILIPu9+8WWbqaz7pNuTD3B0KHTP
94s+xAOA0K3QL1y4F19pW5/g3wqtAQ4La2eW0Iz0Vnf/3rRmSFVLJ6X41Xee
qubPy7DDcqNEYMizs33xnywsr1760IvIh9QJWM1ImnmL3O6AIhrS+U+X2GhP
Wz+0Bs8pWwxyJRrVQf8cy2ER3QNflu9uGOBq1axOYcgRrAS+omYWRbGY2uQX
oXhIZ6aAjDtw5tmMAn6tZ4nII9KU5KvSYZMSpUPkXWT4oQTYN7e2BKVIudXZ
fYZh4QemglHxOjd1zFPc5qPoj3QbA5RSe6/GOsKDd8hiJ+GPTX97LwxxoW4n
zB79ImSgRWa/O9KbTVpvnOV9ZaoaiMc8bashe90kTo3AzG++Gtsu/xTitS/g
o2/RVGVgJXzueI6St9PTdCC3qWjd011z+trDBUPM4rcTBLHB/rZg7f1DL/Z0
mBN0sOc98H2DjlsQ+R2Z09STyoo9Bao9xStcTp4eLOkBkiFPZknsFeMy88zA
/0ehAf1baPw97g1BRpfhltlstNen2YwGqDtmCvySdLGVc3wQoB5l1yDdx9KU
dHVs2Vu5qsMOkdNpQdi/nHSNYSci8VU2ND3WFBx22fgTqbrPmy5pqgTczNRC
mkHk9PEv8RN6GTvWfp0LVadIfkxX4UDsns0ex5kXuRKdK2axFVzfsLXTY6oY
buJGbOmn7hgThyBexh9RlcPiQ0lwpWEBkGvDo85OjECvkiuWqdv7odyO1jf5
KA++e1PPFwoKGLOq+pm+EpbPN/EqGJSOdc5HcVa6k1U1dbdOH3neARlcjnwS
A2p+AzCM3IFqGwxC5OG3nBZ9Ts9CB7CtTcdJfvh83w2CH6HEmk3JjmnYGZ72
LHngx52Ao9r/K26OR5nwoWdw+0zzuLa0yikJIsVe7PNo1eEwZphoZAxQrY1b
L6u1H80ATZaVCIpeAMUXtExw7iWtYxf+R8QozcoyJJXwK7WHuYz6YCV8zMvG
0F7DWqSB4cYK6kk6WIO89nPUPAuu8J276glbLKtnqJoDAixY7/CONtpx+doz
WgSy2F/PS20mjGPsvGg37zJE7G0qv574BCrBQyDdibq1f/3Gdq5NjA45pfpq
BZTl6tqaO+Je3KdoY7nPppZyR/JfaBA54DJUWf8I9PkfwouRMV0t7/gzHwxO
yN5eQC6XmiULDhjhWv10yCZaBk8NHhXho3NZ/lR9D3rU4olLpKsjvyB0nOCl
FZVNh49t+P7jDqpb0V69ei76xuR8pazs/yC3QqCeHldzyJG0TCPo2MDIrLW5
bHBWF9K+KwaHo0mFcWqKlcOn9uirrK+5yGJ926ZLnsPye2IoLAF08LPXZ9vt
oQLbIpMRr2vcics/7mC1ANq0OSPA3mjTZmNtBLUzzyu9yQEQX4xtFkdDFOKa
edCJaLSpDT/+HomnC8IHtTYhith9O300EQ6+Zs/bzJ9+7a9HrnDJN8JAbFln
INk2kjnTPgtJH/Y0ouIBcCFwZUyTv7nK/l7cWUAcqSIY

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9Eyz9ramvBBER0O7KDTqhvOEuelI3y8/h/PQmbJL7znHpR/PVOP7Jg9NBRMxdH8fP0fWyec3TXpkddHg2Ys1CTv8Rurrwmm7oMzcUJjxNvVTcSzKoXnfFAMJo2dnzyDYeZOJy9MVFGn0N058y70109O7lW0zf62BRnOkaSGoWCNpSrKDgn0RqG6elxHl8Yg4777M1F+z2JNM+pYueP7pPG9W7q7dXo2IhzyCPqVBl6iEoEttdAg74nVmQF6JfRzXchaKulgDQkw/CG95XbVb5mXUHoeOKGT2z9u05tT6W2MZCrHS17rHYXYy8nw/UYXZAk8cZi8BNBlTt/9mOeSbZfKrKmt3RwU0hKtPVIE9uH/ztnLSyrk37oSzdjWjA19fjBjf/sR/sCanuZ57qGqVB67CIGaGkH3qZj05s6dWTSySeESWFHMOKyxR/8KgVAcKFhcyopmypeOXiPGuxVpJiFHnlRsKHJR0Lv4KIG9YX06ELK66U6IM41WdlbYlB7Jk/4ZylOdLDrG5V4ewZRtfbDVkNfr6A1ZWTAQPA/WXHmBFXkC6RYgXA9na1NqFzwHuZwoTzvkAKizcsX0Lzn0TX/lzFREAGX8djLMa+X+guQN+vquVgYzoz2iIdn1HHCsRJIeb6k+8k9PNopfYi5jnLRGWJ8iFjylR2CdI5Uo+04tNVo0fHnnz0uliV4Dw7UIEKD6PTrYxTFmp36kEVSXLaZMt0JEMC9F4WUMLhO8Ms3zbU5T1jZHc8fB6B2cA5CVaxDzq2IDD+69E+gKpOHU8YiBt"
`endif