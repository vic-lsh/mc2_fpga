// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vbLGpGkmY+6G5Rao5wZxb/iK+tROKLUCh+ujVLfe+5DY6M8n9pK/P29CrXFu
lCK8VfkHeLWcKo+leIqMOSbXg1qaFS5TTnFI0GJ5LPie4BTd7jK8VzjJFq4T
ckk+NcVI018zrqpl5bQl01Qm1hJPpiBXr8e6K0lRKAhGZ6ePCCJm9jNPY9hs
NVQleN9NlNwR4p/oIyGU5csWIXVxdGhUKhSp5TkdNL9zepUf2xmN+7dQN5a/
0vVsG6TrNhEqPkmV0iNohx8qHULXADpjxbO9h4oJHAUNU+XOiC4WNypnN5fV
q+eg/yJgMmsjFKtpDyh81GdNKOoOtN9ZEPa0DOd7BA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TxdO2IKCgVrAWu79BQOrqwalXD1HW+v3RQNtTxML2abCb0Z6LCpefDGSRCGR
g+Odmkqz/7DleJtJ+jn4tqZ4GmdeQIqQxWlIrEAaOJZBoTiwCtnEBd4LdGzl
GCNad4XI3wdN5IoUWWObIVbEu082dEQJkMy0+7uM8/ecQ28W5qu1I+It99jx
xfe3fM6yJH9LOsApmKXmhbXfaqe39VXS2+UF/Pcaysxu0mZp2/n2kpdyIfLK
c0VFaOYEnmrcA/bAGYdbCxSpSqBgA7U8rSZZcQR2vpFHHGKOGw6JHD/jYZ4A
fq8lRKfdcWZRJdKAheTtPNoPUGXpF2XOS/ljpEkoqA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c1U+TBuTBf6jQwt0WbXl9TUqeNmBWo8gk6+wXEug1cIKm2Kl1yYqCa5g7UoB
ERR1IVM1pvMdp1vOConal36fzQpkZe2qIVApGcW0dwVonfJDAjOTjaGfISl0
d+3fGjRh4WLuhSTVJnIF1xu2bfamKAXXcWGeUtwIEW0AhuszLPhXEMXosEB6
zu/HlgI6ZTm0yWz7bT+U+iqGxuQ6IDKFKWeIzlX4qH801REisSnhsxcEDjHh
uu+E7wjdJHCoWBHLmL2IlZWPOhURanMoiye2k7s5yDHrShySfiNDF/cX80yz
IU87X+ci9ls9qMKzS8iaUBZgS5gspgTVrpgmu9rZAw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DJjKqdjbWowiYhAlx8Hn5tc23oJWiTmhoKjOefoAjM5aVjx2VXkLlCjqo7CH
exUJHSeRSvQwj4bbqFA1QxFd3FxrPrJBJc5EUzyeL2pAweu1rDg9ooLp327C
yuL+pP//WqoVqnsM/BvtfINbD1jiI68g0l1C5ck5spm0PUWijWaot2CXYZOQ
Ja/iQQm4nq5z/JLA60lMiXp1lV/MJ4/CjMC2HPFJ5OVelEcyqoOCexDsR6aP
Ml7oR+ZjEYQ5emOWbiWGvqGrcfvqqgdFfiA6d36bjwmPJCNrEh3/DLHnLYXE
K22m50Rr6/kjAm1lOlDMkevn2YvuqxNRWDuYBOpPcg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ooCxTPp4wyPgRbQQR1HtDYfl0DN8njlf00ihWcFyf8fX9ri2TKRrUDz87G6V
nmSRwOKHPXsslkq+vMBI0ohOZkdyC+LTYdSEVS7CK5kj6B8INYX7MwOyXJgC
IZDfQL+iqKVAdcJAgRr8wR/XQgkSK7GZteSCpUTkxuAUzPOlBxc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B89dBrr+vAqy+4DoilhqSgMhxDNCoO7t5yKwB4kPFA5qlv20ogb/HRVqDmcp
hnhScLAlfqIlEknFOdFXbpTA9qLOM01+c8IhJoHtEvwbgDKMiMYBPNYxphJo
ZqHaxSWOSr1Efol00aUbYQcovlXxH/OAPiV5YTrBBaJWkw6tCSJqrrHC6deX
ygV03OEzbLCgTJd5YN+u7DC33Ft9wLSCjcoLjP6d4gKQBheBbD7ZWkFBxJEn
QtorU2uz8ajDXD+eMut9EG3Bc2zxtldWnuENHoL7q1N+gVZFuFpJOeOiSZVr
VDFvDMMDxjXgmYIG1ObnkOLSF9Nh9XL26SH8Xh1NsnoH0J5eoURFuugSf07k
FWvJDiIjyMjjbco+1/3SNAQh6C+6BKfJxPJhfMjQkjI8tgWzM25mfIAtx6vG
nxvcdRX+GVwvSz4uQ2Nn0d20xOBK03J+SyZc3JP1JQ2H4gTe2FO4jAf+8iaO
ctLnKE12Q4cpEOkJbOjL/NqcFEwtWnmw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gmV7SxO7uW5AEYaWUA00S3Vzf87YWDMQRINWX/Gah7sM9zVE/3cursKOHjwj
YgesNGd/0Yb2nymZDm/AJMqFdcA73lFDnvxzhFshkEZyc49I4aTBNszNkgGR
kg9Dk2Pe1pOjoiMMx+cl6CTm6f4iN/uc6H8x8QI5zl3zjSudhnc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Um0sdkpHNKawPPvicXfjih9er2lRvxoS8wlkX6zTP93BnrGfiZAxLBi4HVQu
ter/3firOxOnz1+dzkYFW9bpIvFojJ7zW0drr40f63iXyQnwV2xWMedLB8BH
fHahVhm70uKOokySGVQ7HeGyIVdtCbdLM/VstYHTPfSx/FIxtDY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10000)
`pragma protect data_block
kPcd45iks8Dz05HJWwZKUD+zd0kGxh+8141ubh+a9ohFeLZPZWzLWgheUtdp
7GTZh6e+L9WcEAIJFiCbwIdCDjx9gzSPwpSCvGDL1tygoLzoQHNJNaDXsfqt
3ltvIEkmYxF5yoPfjO7YKz4iL5uda58CLzGnGoKayoC/P6UBJzjCDs1uFZeu
RuZTVDWSTe/MR8F5Vpg9EHycNsWdY3fodEm6A9QZLEGm9xBwNwgtrfemOSo3
hR/ZRmb9j0JVrQjOH3Jo8DJBISKjEkrG4UQaB7cGF2IurWbouh9dMkWftzgH
jTyqL0YkQ4Ky/icaY1RLKnOVB5iGvEoczhkkWvxQGMxaF8OaTVasuze5WsCw
ouA54JH7Uoalu9o7yBomPIQNCmUBFdSBV6QrwrUyeHJ3qlDvDPJzbyg5WZD9
O2NK5QtCO4YG7PP3a3ZFLlbBKc0UNSoY3MWiTqA+3r5gKKEgD97/C5m5F3qq
AQ5LF6dfbdfu1TtclAN1JA5sYRdX8SxGDBcGsEQLiYzL/Di2swqS7YrQSgy0
dKxCY29D4V8U5OZW4mG6V06ac/AILH7Jq1srO+aqyyoNwGqnc+r3bgrMOJph
TutoBE67KVdarYi9jQTksfr/ppfL87qFsDpSrJnhom79/OdWsb4sOKoaQSjD
a9gKx8s49BCMUOC83srwNCK+1Cf1N8lf2m6ynf21k5/FTjRyELhxX9wSa5iN
eMiztlHENDB/ePdgwcxsshdyoaA9fWJZAw1YQukV/fv9UkYD0B2frrDT0maC
ZI/39Nca4I6v5YGjSYi1f2JTHz5yo5tdoO6c5B7KJNTQdVWb1MbHOe6lSP3e
FwkubJxTeVgUFuAc1+vHA2CeP0uaL/nXbBECTy3Ls0HFfJfb4Z0kWS57KRwl
8nMXM38vz8jGxHb9kM5GWSa4BP8YuQCf9xf3p+WhEnJXwNFO1/VJHzLlws6w
vjBqsWwIIZ2mAr5ZdKRC7Uw0bJB9IV2PNty7/7X4WLInAG7oWGnGrnnM6Gbu
L4pYLS4YebDNQFUcx/fnmgf/C0T0TxXRJebYhhaJ8/06cIMxlVqU2Vq+3eLM
ncDdZi4bUH/0vSNI8jnqfDcq2Kkjqd9+r8beG8rdnu5+Lsh5+JDfdfke6FJs
u5rAS52Q8y+4S7R/wqsNLYoJyBZJYIxkZsmNP14+0glJyVe0QtnT57V1X5cB
keGMWkaqZLwFKvOoHurq17u1TU2Fa2DQ/hY7f/t4xWirq5o6WD2++lCzNwaY
0IX6d2tR4RyOHPdefzuGjF8uirWfwJoqmxtSvauWASXuCLRvqRIfNCMglWzO
kIrTwEyYhl7NDmobiJDCdL6ByVcsAEoYyAtWrq2E5Hr//9IiitizLViMJxcH
YN+1/a5OKkuDidX0fa/4Q4KkSzjGtzNKUzgnhNXOB2apsYx9PdNh+FVdqekY
oRjN6MZr//0RvCxwhuPDdBuUyNWCaoxUFePFlbEmY0oyJiQzzSYFIJDLkAVE
2nMph8I5q4w+ADNw3HnyS+ryeZ1l6LP90hs8aUHeZx9z2zyaf/YJ3y4tKgR2
q0Z0kT4vbow3fUVSe1ryFi+kosBOcunXsNHRA+WaVBC0Ty0iAvh9ULx37sDz
k6ImPbN5gfzBlmb2f3gubeuCnXTzSOFjC34aZ+p9wdHSpYkBz8H0uOpaz8lc
9JDp5z2kOU8s1QTNqL3DOYXCEuVnxkt3R1o6O++3dZ0hQEuRK8FtY4EJ7YK+
iLeZStP2ZWo6KvJOxQGl3HE8/oHEgjtigZKNm0+RxnqFf519nYFbVEcJuAZR
kWLGmt2+hwmeWizGvPR17JJ0r+PoHv+27wsVMko3SoxSEOXt4IIwrNUvoFdA
dR4wumrgM70bsXVMAx7lxNvl5Agpu9iW66ZwdHwhEIlOGde76HsGgZnvSZBc
YUYXQx9UHxxTcX4yMH1aZV37F8yXeif+fjhMujq28NUD8v7ARt5QoHE37mxq
bdkUR8Xwj9ffUZ+7vs/dTsOa6mRK/sLDUS+/qe17pFTcI/ukL5xtDckvKs8+
5pQFYo6/Cc/gSSXJoTVtwMqMJBaLqHJoLamdlCXZzF3iLr/bk8Rx6nLtDaqw
W5Tfiy8urTD9A+8f4+FYf2+RWhWcihDloNy1bSSruTbp7nQhtrokdadrswIb
YxMHIKc6aN6IRBfW1hInDndXlBgyKno82tdUGssZpo1T21tnVbF8vu/LSIoT
jA6n4pA3ITjgYX7h0lvn/H7WUOyrLg+KKD6IhYzlqBJcjcgbA8N0dfKlmaaz
nZCFMIOs1BHh8hp5i/Q91+orqb68IfQiSOqcfBU27sWKyCfnwRD5tQb9hkf6
8gSGLHUmfJURervq2TMfw4Y1KtRlpo/RG6OzAbHmCUwvyWAm12NkzCw6k7Ty
xQ545+OB5yJkQY8dTcFrl0HjsNuK/CcAMmEni4KJWrSzbi6rHqwkBnZtl68D
b019bIhypA0ty53I0xH6eDk4tsR42udaQSngNyLiv2V06/Y93SGDKl8qUslU
Ob//LbkthcCBiXcG0caC8i3TKfyWHdPslj0FAnONn+nfBxYQ5YsDKFtdtSXn
OEgEYnKvVs6c1fYA4kvI+L52qkk7+f8MANonQkZ9iX0URGQBdZpJ/q6wuWWT
UohRUnR6nTLQYCh+MFLOt6dz1KkHRZh2Ey4Z/Mhnme7ekMk4WHTn9B5BmFh/
rL/S2CkDVtFnMVcuY29OgzXVnBGcr4skFMyWeMTt6BlB380Od13P5p2TCv/6
jrVbKV/xwT/wauZNsIIT2H0/x7PUm94IU09iWaEYidR4+i5sL0jKbQVtzjWv
H+PpdYn/xqDPoq54yIwb1PF35+WkzQTgxEKiARd1GHCb3zCIogRzUNNxPfDg
t4PAzpE8R5+kqKSSaXL9k/g+etXuNYPMaSfHiHLmBs2NSyWlNUgJF0OShvxm
g3XDVUDTx1L7UHq7fE3sRgYfzNAlLW6F++6zS1FD0o5Jy4hQ8bvHVl+2Cunp
nVxzM27Gdt33xBzV1rmyP3fqA2jWwiCwEeXIrjElJlEnqfG76kriSNCUaDg1
/infWUzVs1D620IqNFc2GMOVfWIVrb8Q8sPMCiZAY6Z8uNMCfxT7bgQe+ChT
zJS/Of8hS/dnPi2QhlC+P/HPhggyFnv+ETgoBDTiW7KiFD9sml7OuQE25tSL
V78iGzJ+9LhyG3mvqRhVmJWxOP5D3u4QelX2gJZFT/10erDWejHRtfZ92PDM
I2EKHup95V51h4IwVzT74HF5ke/IFjUYbpaL+tyH2GwKm/DQAjYq9ve8cGjZ
kmhroI9UVdkOA2b4SnAjIZyAcOmSRhu9WzWDmcvOqcxGW3ilPx8UgPr9ro+N
6vrgye773uOigb5YclhZrCXnOvHAuxxrYoNYj9OjUh3gys+7yGQobzEnOgvy
t5e9RIcbyDFSKizE2HdO/vpZ/jK/7Qcm+9NQrbdehkbYdKEXJqMQFxtGIiML
nArICuVjAUQm+V0aU31aJgJ57GUSOtggHdm2J/5UDj6928kDfUDalFGaAXig
KZG+OhnOeNqtNkTioBARS02GojMR2UgWDZyKavUkYLcgUGJysB9xuCP4LvkC
3//YMdWoDH3t9WeJTvcrG/sBP8S6pxqmDq6rJhiF4a/1j8eVYqCfJzGOnM/p
4N6CWIw9EQmfjzmF7YOsju+M9yex4jS1WXiodT48ZcgBM87bwciuF494ot7i
Z7+DUAeGQazV69xbpMlvmRm05aLt9X1EK2Kn1BnizT1BEnG+HVRQ4kwr5W2A
3AxTheziUf6n8rk84abG3uSK4I8/JdqCsHiOzrZZLcOlwkb2u9zfhT9CFsfJ
kEFU+/4MKQZXrqSghCiOWMKiSnMc9ntYoFlXax9OF8sjpgU9CrwoPykrfMRs
gNJod3MBcfh6+LfD6l4MqNVCewvIezE6dXd/0Wyw4MXXaokio3ycenwZefpg
pvFr1gdQiu5GjaVarOimaqoIR/S81xikZ7v/B2+xQr7tU9plPGOFTxsOJUHc
x5J4g31dqcGCTA+BNf5XB0j2LrCfLCwFPZhnjWlPXktFo5xwKHZq3tz5bVjc
GIYKlifPylbwWQ+ev7qtD2T2+Xch3uvWXxTCXB93uszpeSyTPXJ9Z+6Qe/zH
KJWhb8t8ZyflRaTwAfkkjfUvRrSGLsSxGcdA/7+DOuhJU9zh9bRR1j2rzqGj
eKrxFMwSw6q8o3XertMJs2XpBqhkd+jFuj7rQxzfi/+4uMQEWToN8NOSqs+c
ysUzdrh+bo3IIh1mLnSUDiTmMtzjlx995U3lHmPeaBcFJq7zwaHAPWYTmqeE
9D7cotBCDqDISaakB/29EOMxA/KHou4iaewSRQ1MNRmjNCJWe+sv1Xl5Efru
n9jm+CzBMWlFMUO9Jv5jkeFzPMtg2/QM0BjsnTdAOVoc/c8bRCnJfDfX5sOd
A3on0HlQGg/uaZaNviNmfNgCbVThumOkMBYAPQODNb2PUQcZp41iBfRZM2+C
g3Kcl1P/0wXuNa8QFrJ+bci+JFrKCnuRITYA2lj4QvAMM3s0QYbUpFnqDvwe
PoAn1w8sswocuS+2CyHXJo1zlfOYbpfZgf/QFLtwzQ/RIlSrn6r9Yz0BVm8K
5pUEskWagBm5n8R8ruKr3K5qPvkvP77z7kWWgF7gbunWpxpCIz1n+/PH/6bt
8RWquBhFFy70DlX3/tk16v/7VXqxmbm9lU6k7LmTtWNXtUkDpFiz7V1vC2bY
1BPtrRXqfMTYC2qOekxj9d2OwlXtiNttgSE7vMikMOJzPvDdDY0LPL9bpZ1A
BS5SgfMQSVdicfNlIF3e4BqwZ8TpmwTHeDTaCjlwWPjtKrBmXUq/Ca3qByM2
qXilxI2zhq1leHRzfMlZk4OluqVJKqs0F87XigIcd6ZJ2mc7lLGNruMbtDA6
8Yl8VR8u23fDuHzYT9okyOY16pvBKR2u+Ln8QdMP4PfZQ0ctmnp8osIUZ7Ii
RCNw+9fpGPjSUiGVUR2z/Bx+qIquF/qMgl2cA9mKs/Y9migZRpUl17UqY2EA
39Qeg57Lxu74zCCxEsVXzL8A6Ky01ShNg14RAPYBbb47WSeAkWf2wC3pZGC4
gbQMmrAm4yWQzgsoE2NruKUeT29bPEt2qBf9Wr3SNKuw0zyvBR7MEr+WYEfR
vuXR/D5xbhYEF34WVgNIcF6iPWx+ayewNwoKMgGeYbWq9AnfdFFfVYzIGWCV
VfVYlfOzgA5be3wd2EzzZAP6uGBIzF5xn2fEhjeg06j3gYzZ5Vv3zQwIsboI
5ZLc6GHmfRM9Ny/EtyvMgOro7l+ls0PUOKYUR3rDk7j6TvJEElB7/Vla947g
9LiFURcBuENbP4dCfGPydfJqEiG92xF+AJ+zKIqTzfH0I4Z4SjXE3rfUZ/vW
tyTfwx+X0m9mB/TqhcjMdjIbwopZZGT9aCBtk2rcUuEz6e4ULwGxSzVzn6l+
UMiDHQLrbcYh7e1MiVWORTv9YQa08ei0gkv3Ze7XdhLtkL+KWKOEhCw1bhO0
SE3pbD053oeWwEMO1SpOpR4JuKQnfSViRp9Q2OWjDVa9Vb13Txl/bA8ZM7wh
YwuvrQmFph6YqCXy4Pf7B8aSnFcq+2J2jIa4fo4vExhVxLe3Q5W7FvPdCphK
LDWIDrukdSQPoFpxAdN5XnIZ6jXMwkVbn8LrNKpwrJUgphxqd4x4W0VwH4F0
1g6YZeqUDIeaKpn+jVxeSV2xavIKKN5KYJeMcakpEOTPcWKwRylUXfcqK5JJ
NNphaqMEFaRXcmqxl1xNPmrcs3+RCyH7Lr9pvivATRuj0pbuw0egcpauJeqs
AZLugW/qLwLPKdhyarUx3julCfv56esCw+PfNanwzA91CYzuIpR7BmRRsh7X
QcusJSdV4O5p1u63563OTqK/nqX1my+CCRimZFTTmBFKe1pHVWnumW9FwF+F
DDt5LnVlVhg36X9fUU8+weIAJLsteHQsOsuX+CNJkTrh/V6/7yTJCRDrCE+s
gyUZG7HHM/oXxlz3IqtqfVJrVr04mwxqmJ7uIY+xGpJqckKV/oRM/D6/TNco
VaWsQPe+EUGEWF0kQPRbTD4tGQD8SzntVe+WO2ZAECwUXkOYeEZM84CQCAnr
8326ukKmEXlRnLUAf1ePbcgbrJUudRMVH9rE/OSnONMZZ3Q0YpA56pXEGqfB
o6LPwT+E1HhS4yfBeu5oUEbQjwzoUWW3rJXDeIXHKeoStQWbZeg1SPXy8uLo
UTzJwmYQwCdCzk5iGqDR5gn1E5B+f795z/5bKAh9OwUZd/a3gNt9v70qryVo
a2AjnlT/jvS4EN1p/164gxweaXenboOfeT/HGeF0lr205hCcPbyKFFOtBe0v
Wguv9Tye8+ZkmQU5t6P0zAMQkkPT+OO0L2r3UO+v7avAIsPuWc+CQ5ZJb6uc
4MrWm9qJJIGRVDo9ieEOyzc7/XMgO16Kz0SoEvjLTylva+nVqw3c/mdWi7Wk
0EQUWEwy8dDlTZhLjjwq0nmASusB3T2C0WQytgEsM5wC5teAOUeoWsVyVLr7
zMhQx2pOfSG615j+HWDj6eimVHcecnp9E2rq7xofhiQrlOFfqS6fl1OqTxpU
jNfsy3ehlohenpateh6Au3c91eLLfq5j/nj8WR/Z9zw2bERl8e1PC4dDd0/5
5+wgFNJJYPw5KJAL8FHRg6z+enDC98why8vukONu1i0cx4BZd1HO+csvylCT
ETHbMf+t+P09vYgfaWEDoVFkHRIbL5+mN63ztAZbox69lwnaTdTBrG8AVpmh
bvfrPZIe5G/kTZk0IK5GWUUHJpo+YP0tgGggqXeFTc+DgESmFpfZ2OKCA0tO
yeBqMBaBg6Lt/WR0ZCEGEnqH2LyGr9LEdc/4XF8d5hj7y15xMjOIrOIYwefk
YZ+abVymQvcZn4OgdAO+GP+aI229SRoarMeaL+5mgty0rAdM+v67Wm5zmSGC
+2jiGA/t/h55p694gcGitukeU9iNVPxN3GqNzhjxv5INkczOU179kj0YLP6C
yxmI13/EV7V6kLeFLpmK3YbAqrXmxy4I+x1USlXSAcQjNeplcAtcDNbxK+Ex
LEZvHKUNKxk4ev09hSRgwGE56SNT2+DmaMWIOixzCoe+b42CfWFtVx1aCGjz
mzoN3m2uAZVnDsOWHMxrM2rmL3l5zIruUOq2FDnquVfcYyCLwRbT4UeRSYtO
ljj5cAo1HfavIauTQYxx5HgYsLk93eHzColVFqfuGkp6ecBa/W5/tEt7/w3S
loUs+SsIJm9hmUA9BTxfP+BdAzm5Zd1yHTFwRS2Ci++HhG4WR/Ap9Ul9iMFJ
TfuWCCJCDlTpzyfrHerrsLu6At70Wsy+ANepqA2VBF1aWqrJQ/lfMz/hY+3e
WUDIgKNYdz0DEVi/wjbUp/ZVLFYc96lpdoYqYkgBSpOAjKBuwRv5GEeH87al
5QDi9zl6jowT27nasPC2cAsn6lhoNa3flrE2ebwBEOx2oBr4t91ecW/aJOkY
xnj9XpnTL0CWF6tig6Wb/uUia3XaSbVVqy2xHqQCIOQ4oEEl+uFUMISpW2zK
FX8V+PlK66mh16enSvk5MwVdTFbEGYbYptr4YK5aPuE6HKLinnDXVsUsBYvp
JGMDSSoLcLvRbVkWGVKYalplUuOCRph1i7rpyT/m5ja97DCRZrwVlaLjhI3Y
EZdujOBgP08yx8vDnPzHPYGSP7u+WAmmYIfL5daxK76qZsrTYt3umWbJW1BC
apZ5Lv8VyYCeLoyURt2k8ZkXRfAXt/au9dz8mPHYlxSechgxQW3FBIynAA1J
ILkhKxW/f7CkZmtXaaYS9qkYhtXNPtdoN1ps78pqV74MfRLp9qx2ccw6Gg1d
S6hPRIlVBNxNuVPtnxzxO2lC79g0RtejaZFmQOeVAXfU6HOTjonZLpTFzlAe
J6WdG4VEoQANZHq2tBi0kFGspLQ5uMCFG9Z7rrz+Ner6qJpxNueJjVEpunsQ
1yOIA+1iQXOZ0QHykjmRU8p9KCHeeDTyXHYYvwJ+RdTpHVwwE158QIqb/Qo8
GTt8G/Xuh5zY3QNKerSIdiFJE4JQcUC0w3t4sFDXiAiY2rY5SLfKcgxbkVph
3eDMl5PQOhbO+g9AqSeqEQVw0jWN8mSB9WxczRU+mRbeOs7OKP1m1vEeH133
j4uCWiJN8/X5yv3Yw6p79d4YzXLzPUV6P9uDHCrWSNagyRelJqjxvKRUC94O
zshmS+owa4d5SylChWxb0Juj/kYDomwI0CYJv8RX6UHJCjWg9X9e5ZAFO9mj
C4Z1z+fAM47sFSb2LXBzy6T8S828NE/IPM4wJtsqAILlC7IGc0s33CXpnIOu
hO/w2/JgVJhSgGP0wUoq+9Tcx8+Kz5BspUS4WNq/hhvuXcwv1EIQajYtgP3v
Tx8sT4eNYciR79UYBGyXqtKkw3jFMGSBWTIfxdDAtFLRf43jovWSp9nAw5UV
Ys+o9n8+bgM0720/+W0DiT31QuCc96ckIHL8ABwHW15dqJMqs0E3IeW7JQM/
11bYiGY2eQ1NGRU3x7Y21m2pJ9myhcxUcPItLO1YkG/g1zm/gDUZB5vnr8Pj
MkpB91rJCkOphPAPkm6Uz8foVRkBem4iY6wO+QWkkD4QgPpRSb6LJ5A4VkYG
fmpg0nAwnmSPorH1nsKLMZ5sf6eNSU5IS56r39fJZKf0RFtL95gHv+k2lA0k
4zAkMgdxgTJDDiY7BjszjdeeP0EaY4XIFM3yGnfoj36doYYHjrzU56C4iX0A
hQRN25538RpehTsv8xO/TGUanak0UXhAPIFfNybdLIYNV7qkUHhoJgkabpIZ
6s/z4NvmY37ITIShe+ZklIpIqtY48kyRfh0Hq3YuwFZSlUfuTvHl1nEt70Zy
RwUphUgf9twHqFm27wHV6Zfs0hwgtLEnqIO1nyaSWtoM6tfRWGDZLwwIFStG
kZIVFi0TgPvmKVvvfg9GRdYkAnLtv3hIsRDPGxJjCBhYDtYfVriS+ptFmMds
RJO6m7UHyz80FJx+4acB4Z4eEASk9fxZWdPxkwx/m809afOfFab/de7Nv1DE
fEJhUCLTTs+IgT/ms/DxpOsDPEer2wwYuE10jhgzJabK8G3tL8+v9Emfo3I4
rOter5m+gWgVYQLthCa7WI05gq+wssIM/ezn6e9nN97iBq+vdXJvDgOA68+A
7zE68O5ZWKLyPtmdoyrALVNGsPFVMjniEJC0Z63hY1mOKAOL5cdLQYaDLRc4
nZPjsoYFgcw4JT2u0EKzPAxsnRNyA+U30mfS/Dp90dqwdJl6KwgbB2zRpNlO
UB6vxmUyZrGbSsGQ31IZ+IpP9kjExMkHzZd0XnUtKa6IkRE6GlZlmMPpzozt
xr4esAo3il7JF9SzRuuZdoY+eg5xYGDHoJjnDL7A7bDECDP9mq2LJwmEnozP
x3WNh3BTIyjTEYh4lDdF+SRx55UagmmNCT+HddD7Sz7K5QS+fZQSBirKQ9fM
EmAJBmZqntOuW0/vZmdUGe+5wNc72WzBTKrg5AoLOl6MbeKlCzkfi4rhQgO4
oSxyuB4mn569u5ScNlKoRd6YDRnlfimvnhAhY5MpubihAPJojkNPTMfKsJO+
K80D4yMyF2kg3jK0F+qk4l2hPz9mA6WOTZaKbEZjdqmX11OYdd3gDkqrtHX4
a2jJyzb1noM3S1YYEGZPMXMWN9Rqqr4INE5hS9NGrJBv7cVy5eQnSSePrgnz
BOVPkO7ctkpA+9v4W494TnfrXOO3wFsxYCeFhvaRz37ZCVm/wC7IgW/hamex
/m37lSa2T26YJ7M3yVVkKTpA/9oOXCjmNMoJs7HgtS1nQkd2jmw086FK6/m4
EJKlKeO2yoingjUBkvqAUAkY1PQFY0eKUJgTzxrR4LAYgJSJNg5Jvfb4/3cH
bd81ewbvxEXnl14BbVoI8DnPhwqzlvxAAqhkFSlDRqSUKHG62eRNMKembKsj
xS6MNab2jOgUVr0t0kgdzhuno8CNjQ3p8Sxo3XywCeoR427+qrn7q2x/jtGR
jnkyVtoCE76Yc0djZKsGkD8ZpCqdFFHiUExafF2aZkfQDBsCqaAcLztkvYxc
rwJI/RhgL2eLGzXPxvV/3Q7Fatk3wuaNxIInHcKSsa2zIorLQzuYumzTNcVr
agUrLM2zxEiqtt2o3s85VcBld2c4FDFtV4WqAwBdDa/d8W1Uri6ryqyReh5e
RvbFN5NAK1GL6YG45vLJnaMCdbTc1GpOR+hjP3mO4COuc5UVRrrV8vgNyhg8
s8iABJL6Av2zYqAYitFUqsUc4DP3b3sVMgQmbxKC7yjcd/w7ln4R2yju6LjR
b/WxQqV4IQ6PkfJOrRXY/TvUJB9LWdwiXMAGxKN0e1xnTru3OgHUt/AmSHfb
EB2iw364r/Vbs2vNeXV+twv2ROrmhIidZiZ2eb4jIQ7jGw0EpmpE57i/Y9it
4vY1I5tztFYsu/AGCP12hCMLEnLBJC/A2I3jUzyvrRfVi2GrPmeSYsXWgak+
I3jj7Zpb0cRJ4zpsj9cU6MoB78VchJa11hRA4XUN7Y9Fj6GF7o6pQtuXtn1i
L4H1p77FN9ku3DeSQ8bFc0m+J4tLUxmX+8Db3nLUxzzsSLcOkCDyW8EC1EPk
PWAZw4kOMTELSlwvqJ7Y9d1LYg87k+Nkuun1+rDwfMpKYVriDkOBizSP7I8z
lArD6XNqlnuHurEtMQK1PJHbv6/IsiKltYNsc8fa+D+O0ODW4TbNklvRzDMy
HflZ9MFLmyRW/DE1rv0JnlRsD1CRJTPZzJR65rZR4HU29ro7FgmI0qwkLqTg
aWsJuMpseghRa67XylRGUFweLpB9zAEFLi4ydQnnaqrM+kn1/JW1oYTzx27g
0lxWS5T0Pz0d6JF/pBBzNqDqPeyg6L0D/j0ZQe/CWRgjA1alioxpayi0T5Wk
vmsZ81v0NP7cG/h2aLFqKpQk3R6eZ/YfzGVpbZiJZ5RX4aJKlaomytB3icVl
sBCja/jfMPbAPikaTp8eDMUXrBbRJknpOTF0nlptez5CDDq+GHnCGEcGCNKR
KKc3v4bFJv6VIpTIxbS7JlVbJ47Cey8O3MlRmzDDR5xcYqJGnlFsTlFTUrgI
XWRwXcESSLUnADK99h/UVqoZQhD2s7qbKOux+JlRxvp/1hTrUZXANLrrlq2R
odWoMIbLEf/uJlA3vIV2U2SmmGZ6ujU5lD5BAq8q7HMY3t7zhfkPsjaeyAvt
nQcf0KMgacHi4YwKEBmVnyTkLMS40o4V4PiIXhu6XjjQGEKK+axkoXM5NH5L
u+Wua/nhRIxQnn5a4SkTij/ftvOdDYpim30a8sVt5U3G50zh9D6VYS+l8+p+
ZufP376MSx16LGOpFJH+lmbMdzX5vGhAqerhEKIwpys0QM1jb6FWtXO7UkEf
korM+ysnYsasIgVQRg69Em3AV91qpxeRITIiG7qmJal93PYq+f943+1ojKOh
UuieXK940j1RjpNDojh5dYPuyHPx+WLK8DXkvVe0DHvXwPZkJeySVbGVhdr0
5+FvihH9ChXRHvTjlKytcrzizDBhQVR/f4ZhaTr6P8rYJd6HXVXNCcnftS5C
BuzFrEyWCkNaKbVEDC/nyB0LmDZnO8pIhNsJUSJCn8F+7MwTwdJq3iMzcTF0
8+taSuvW4uJ2SPKQltmj45hEaAhCPwWM/1KFSEKWFK+uGTg0kfyWrDJij/Zd
sCoPE7amhfI3Zlmr80cqNmXl3qHCwMtGVWG16axt7GoLHwdBciqIbjdkoQEv
M2YTCVHWatEPUTpHmG0IYGQmw0nrexL7SP+5MAxLNC3VI3m99RVDmINyBWFe
eaJZC3XWxBnnb9zyaEGBasaGq7yTFHW6OB/6VQQxU6CjxL3nTpL3adzn3gCr
i2IuHfj5f04BHA0ULrILgQFCs/27xFT5DaX4Gxh7EqHtRTtCmkNCVQrNIdZl
tWdzdv/QEr+b/WkmDA9Y3HbRybjyS9k+FR08nGcel8E5h6mAAu6fy8XfIUQE
E2c0/1LkJK8RIbf/NvX/lIXzUnmWdLi11Cz8FhMbatyvlvhER+4kxRuLvC8D
mqrYqXgQGsESokOLB8l/I7uj9gOE2p1NfNauNfo9BoEJPadeXv1MCGcgYg2C
QwUCgObXz5+VXLzoohdEfcQho3UvEyoDtjwZYn/3BMxnMXTII8+Bk8bCjvYG
VUPplEI8H7WpuriPQEp6ngA2PWjurB/TlugzZ8cEh0IeGC/z1gKeIL6LFBAJ
0NvZ8i+vLMRTtS1GOhOya9fs8tDiPVZZoAJeThyQ6fmpTJIzxZP3J28SRqk0
+cCtL+Jse0IjrjhdgijwV0mfVC3FKvpqgoURUUOLSSZ5tdn33YyIppLNXDop
YdmIVqVGTItRrzvlNuJGnKYOcllCOQlJrc8684SkkD7dtjjuOvaD5e4aAVMU
MS5LZaQqUuvrYLRfvRezp/Cyyr46NdG2qWpLluojHvvC+b1ajeTTfjtF9l87
yvtATvvamaQ2VfKbdg0UDcOw+/NowLeeZhYyZYXiV9KR24wPrWXiY530jCcg
b3Xi9Q7Jq25acsxI+UnLMCqHgtrhRFzjGdWx+jJkg/hyJhsdB+2aVPbAsGVi
QhX/CYYWsX7nDW17k25Deq21EtEL690Q/Uo9ivgc+vz49f4/JayA9TzkLV3o
GITeOLMs4C6DqILASSfk1kGRdKm1ST7+zfYHp2XaBr/bKZf7uSr2Kd7V2Uv2
QE96Igx2R8bGXX+1vOdAs5g+k1Xh8a3/W1wjjhEZvWhZ0ECmtcbmJmz2goUd
7ZXZwMCdD6bX5PVuLBZajAo+D2ScgIgy9a4Ddqq9Lubd04sNNFP0/tb5dXxA
+i4+lA3M48NEYM2OEvkjO5Z7Vv8jzNEBdF2RBLSfiPeUuhFaPWddA7nWQnQk
g50haDfxuBwcWoiG6THHLYHy7JXV+l/EuvesOLZTr09BvVBdtee6fsj+wSfR
t8aGtjIJDHuT+0BvlFvu2i00rSQRyRmZeqFubFoFTD8T4UdYJphDz53E7YRQ
1+lxr8tv+HnFA8jUHzUGOtcVG0ZXp62BLMUohrF2ABcIQAkB6MLyJx72mmX+
q88pEU72iSTYWZtuaIAAN5eAVKPkvMeKgRif4VNdh1mQtITcPtXQWSteO7q8
Rmi1EuxuPx2fOMpVtLdD/Cii2zF/oX/dsE0icHyO+VGYnUT/RcXArgk09AKv
8Dyc2isl2pusrUddZfK22isV5AYj/3d7YvfVomwoI3/mSQBBkw/qAii46bWJ
x3sa1pReb1C5c/yn5e1tFTxvOQsaFiztjy/bjIeUsAESCWoZIdCUDLBOpFIg
bmd+qeOylDgRzQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfTBNcL1nUW1I97ar8CbFy04oCXWEHGSyAjQxFo+Xif2INzeDWKH2vYoa57eDFCL21USkUTmi1UIMnpi+l2ESMgk+Ze3MHbvuB6Egi+Q44oFzfYDmGjNggx5cWC9B9YEztNMtFglRei+eJrafSvc9Zd1J4ry+TuBfw6fHzdpuuOVGSb79PGQqVpl+36zytBqKinDvav1buNXumnlBbYWqo49NiR6BfrzpAb77ESgdewsBxlLgxBGGf64r7icGrwZyqkDJ8XErgygNjdA0NdOdIZPb42X4CG57n65P6SYVprzVWXbmbu9aWrKS2ZTmpJLt0FHYj6EgNkoKkL1VSBM6YwTxxp6IjD0YiDMvvNa5V6N7mRUOpTIdSNo3POX38iiyi5F/dhF7C5aVIzLs+5IVm98UFjAuZK9H49oxLi5XG1ZaxplX7S1KkSfC72kVg6eqHgThv0QNbrCTpMzQbd0xOD1MVH0KwgdG+C8hsA+s4mgJfWtAIg9JYas9rU+dRCHGH+LSagyUZWdpzuVjsZVMgA67qOa86RHiv1j/kgGJoTJbIMskL+UbS0bTvHBAHbNyZKFXJhI4/TjvCV4h4lj3TGbEArPUEDI4Fm4aHNQNvmdt+qVGfXWZPKXoTX5ahkq4GcQ1t0e7wCJhTYqPO5UHN94TfKGj36Zyr6QXMZFv+LIrCZR2Eca+NEUF8Iyn6ICD0wLHZWTZ9ZuVv7hfIKbTQuCM6tc/2UIwcB/Cqwu3WIac9HENeLwuicp+ZHxbEZGdrOVcrX9kCNZ60e7e9Ghzmh"
`endif