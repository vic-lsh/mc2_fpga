// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aJF7Tydj5B9b95ZlSd+Leg3low+H7D/eLx5Yyv9919SD6OXoPUfjUvm2CuGt
TDtPtSWj6288g/uOTSVCcSoEQj8wINDQgSmZ32vZzYr3at0R4L5dYzJTBYgE
q2puWcesv+D42Oa/g9E0/2QJ7J018duaaFxAwFjpSKEWg3V8MNPSkGreI0zl
LUIi2e8ucPpWxxI/7Ububofs7s3Zmn2tWQncVULzg2JPADKGt/jt4fzb+oJK
M7guFq5dtuktNv+rX4uJywIGGBkxpkQs1DfYELSrFtffATHZVC5IxLGPSkAk
chzFTJdsg76AYfyygjeQHAocN1Ttps5/mmLIThr5vg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f9Xuedmi4DJnCg3LFLlD5SdZvJza98ST9WEmm1PqpHpSgd+rzPTq4ZHlRDsq
fkJR048b7b5m6D9drDqoR9fzwQnI0GLMtdkTsV73ZDCbASWf3aUJs0sS679P
DeDxCBMPVVYCgIMeuO4AB3c5Y5rqKgJIAw3bOIR1ZWuo08H5AXifjQKc4dc+
jarMHfpNIuuUMtsPlCD0ZAgo9mrjZiIfkVS4FA0xjorkGF667OYtSvGYVlu7
JWZ4Oai6Oam66BIcyZ9o60kg7Pq+0vfGATRTf5sTlw6ZpgF4FE/b15nd36E8
Ue8qVLla08UJ3XG1DAFERXetKaddvm+PZyVoE+YoBw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MIT0KYIfhuUIp+AwHK68ay5J9kxp0lL3mevgzRScDCd4kRlzX+CogLZxPJRR
Xt+yUqZW0mLCn9eDC/5nN8doTTsds6tfTnEbBPP+RFHt/HFLnPsD4zQSm+ci
YurNhoQQnvbm7qDlulrMSduweJ3b7FhsmGwomXp9T7d8CQ0dzu0nPE21UqZn
RWQub4pKnDMBRQPLjygYu20aSA2dSV47JOZaDsoQCvnXFVDHd4Wwqn2pkJtv
daXjadkitm2JXmNOLHv46Kyv0g+mkrpCJ4BNyUoyQA0I03YbF2T33nLA5kDC
nT0na3UYkmIABe0NYSmweEB8Da+eI36D13JkEbyLXg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MwSeJbXGE7jObNPo7qHNBKcklRHC0C3nYqcqEwCkeedEJOegrT37vs0wuAX/
0P8IheOH6DoqbkWnwXxdWi1tyNuAchwZiyB1uOVVck5fhtHDdhrp6xwqaozf
6L0g5LiLsHhanR7esYLybFRUjFTXAfc5snAwSf+R+sdcY/lP7vyLYcyKHgMd
VrTQFJfGrIAUtYsaL8f0YjOd73L3LCxkeQEVibFmeq9RKjtonZQWFSbysRRu
mqbStf6+1BZMV08nWcWYX8AZWEW5h36j68iSboZqr6momLswPKT53rssifCx
/h1kKXnVEv89uwVWI1CG+KaLU43wEdut5VwE0SjE1w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HUU30pVJB8lyKxQeLbfLkbbhitZEs9YXc5LvYYXJme/YcI/tTxES+xCptEmC
DMdbrlx4ZkQLmYakZ6fCc0aSQ/rlFDM68bmV20yO7RL/yi0HN8dib+Yl0WO/
upXxusFrBVo40okHyEn2J6a7cCv7nVshunpxkcRu9Cl9bkMKiuI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JmMALdhGgzCSnyZfup7jvdf2ZsHEGkGSsbeEypTQf0PJuFFB8DIeE5ODViMX
pbCzxxeZWzxSXWttsGUDaL3o+iSs746Qct/XIzolhI+CecTpIW1J/Iw4eZ2V
nGDR2K21NbtYXTrc2YEouSyAUVzaYfDU5ItjkwldesSYvHOyLgQnHzdQb7xC
zQ9GmNacaMiSDU4YSzvWb58GtwlS07OXVkUHFTFCf/JaHWfhrU6gdtzKVXC6
YjleDtECJchQSl3NvCuLk19XClfYGaOksWgajvXuv3nAvL1qU99Xbn9zeMiR
0oGpZpO7OqAXYG9tz8PFbGzZ6lv0pezjWns1CHmSkl36SVhVbMe7gNgZ1nO8
KN+zJm9OIGJoaZTzmUzxWQDTg2G4PvbOCaok8V/q3qy/UtI7SBQqSw+EvNtK
BX92d1vjoECRbpay+QIGM9UYpan0UTSXKagvuLd9k7pkUe6M3cqtFbUC1DbQ
CoRGzXy4PUcrAw0AWixn7mqvJQrP50je


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VTmF1TKnW/g5uY6yQ655xiuqzQrtDwk9jDwp5kc39TdL8EKIGfbJ63SKxnUC
W+qh9FXBYuHX6LRQ2arO4N0PHYlXXAzGaIw5w58dhr9BpTu8Vx5CQscnle8j
TvBQz03rfxZ/FZkOZM1PJ5BtQMxk4FNWhTEaWTPUvLUqzK10ZWY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HBK/kq4CAzsO+j3kmBkiuJ2iuaEGeSo/JNz7/OWhd001qHmbH+uGYVQBdzrh
C5RRNPMoLVXgsF8bgRB3bIf75Qp5KX3WbmPMNnWWkiKQBnW3gUhdNwdqtELf
A6tKuBw1TqvRkCOKZmq2Yiso4QuPipzluVkyojm0QvOneUCi6dw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1080496)
`pragma protect data_block
GWV8ce7m0esad/5JDL9R3p/tQPN70KqBZgTlH6xAUOBD6GnxDFbRtoDkqIXZ
DqnmJtXzDWSBegULlcB5/k2jhM+UojaT0bagUdplNSQmEeX0AFTNXMU8lhnO
DkjZBRjYzz+TKguOXkydGU2pUcZn8pK47uWBF2lkJaKQ5GuHBNQKezBGa/gY
xeqyto+TdDZEudXCuxQVY3UjtwS+2d/vAbsHjmxuWmCFzHysBr8J5w6kl4md
hW8gNgyvNKk6wtYjc1T3XZG30OEaYz0CNjWMkanD+4Ow12ruLpYtbespZl11
dr2Gw17NNRK/w2gjnqeW+XiL0VhheMffIVidEWf18TsADxdgj65xXglyQN/2
bDJrgZqXDKxlRUQ8TU+VDXiVaYw5MdsHpAhBdChKywOBE5rvGXHNOV7cnfVw
8ZHnkndfyM1pSjrOE9CAukD+/56aMQeJUle8+G0Yivl2GdrW4EyVHF6b85bP
06F3yV9SyO9VRL84v/5SBF6YhmTKAPH3gBWevnJ05GcuKq+B+PYaTr1LBAAV
VAOPRdsD9f2P4ZJYnUjVGtVkgAksDAGrWH81OVGj5Iyh9CzYGfcSle+sQfDb
+O3rv9r67dOVOFuGlVBjQ0hM1q5KFdBVJ1ZwmDONEnbS1ZBebe75wZ+Ha9cB
d4JMaKiUDdy9Pm+M29AJGqC2VaCs3i08WiOdDSOHSOt0sjCWwiGae2sRkPvg
tsvAwxgtjkuPxMQzuinEuhyrrRP4VJKwoMiySltZDGVWm+RCiyyqi/AUfQR0
vTe/arkuM52aji1neleU7fCKsH2sFzmqiYt2fPmbOLPgpTNQ10mlpOIQcRKT
6ioBurSUFP0o8DG7tj8U9+spJ225AbiRS1krxkP5A2+29NTyNaQDGqPaCClD
JeIheZRd+EpRzEZeccBkjzsPbu6ZFqszfdjW6XPvynQzlNLQHk/GIztCXLdW
p9bBb31mcRuCG5VF7PMiIrbEyOSeBbpFNu20/g0p+jnzPe++SnsUmW8qPMy2
ZBL8b3//zUm8XbX/sXaHfoWkrmfOugPjBIT3p3/d9J/FB38pEsGioOzwJC9d
WQTDJiBO1yFa5oFUw3VhP708Qr8o541aHpYxbNCLBnMo15fJnbXSJ9P5e5Fv
fqR6CNYhhgXgUmis/rlsex4wKDgDE+vw3Z+jP4LwRnqur9jfimjyJLe4i1Fq
t7/cAB2iot1MNt9Caqeev45MmUKuXkDszGopo8ixXPf+1Kamw06FixlAq7Tt
JX+IJm8Q9V8rF5G4y0Ygc3Hwd/+nRN/F3T32wRNCp4hgOTKXOMXSPq04u0D5
dQ1NMQYGqmsW6ynyp75GfJPeCEaSSqLzXb1zaLchpkeILoD1vEQuDUG+7Odq
hDa8oz1bIxAjtVlRe+Yqn5DLs8vsWlntgC6lQWF5pFkKv3sdJOuL+JWd/yp6
ul91BFIWMR+NEbQWsGngmdkYVipwqITk56nJOCxh9DRsf/TRG0IeinlvhTNM
hehzYcNKQj2fMIgrWBJcyfnbIPRbNdzsb6BymFuFieMeUFDxOKN9RjGFv39M
mj5uS/ccfIF39AbGV2kLuypNKq4wnY1YB0jsHB1y0LCLJMZ15c/XIZZJ+2rb
r+qYKy+lYfLN/pNfTVIN/sVdokri4PPGW+c4Sf/4Ycnu+CeWkLAmJGL4/goB
jTHwiPKBESkT7/lJuUTsT7F3qz3L9yURhIlmWt7pEUxR2R8xalaCIyLS34B7
aRwoMz0JiTy9ruXKSJXTLCsMxwK5NWrMOe0ugJuj98XcaSa7zyGXlUYph52C
IfCZYHGd6U7EN5mfg6EYJdRAQ4kyYZwYVfOLAKWQXpGybFNwt/g3y3JlPkVx
RZ6SbnY0H+7ETTcPnASopLTOuamBz1O2/Ib/uuCYHBuyUnqUAgq9Jf7V2HQE
YGFKQ4S2mwAKP8wafk900/s30mQXa7lzOkriV465Pi/rkR8v2IjhBYJjKRmZ
1FpTHQgw6xdelLllMZRXUZ3PNPnJzTVV8DTkfMF6U8aayQtf9xbZaIlgpv03
43Wpt29Giuu4Ukyxm7V3yJEPw3PJVitMPlVPgsX8og/ii0VpvrX+w4Tr7hGy
q7yN5q9dS39jqoJlzoZo2zLg5hsKbE5ZuiN/NjljJVWF4HWZ5OO0cpYUb85M
IDkHhq30PndHFGON3B0alJzB0/c/9mFELgcHG+ZCRoyNtaMGD0pCwmGL1W0U
KCqOBnpuN01P2MWcTReWhaxTJjnOW84OMwjURtWTrEJViDX1VVPIMHceRLKi
BD8ihdxfDsm7QCnrTRtya3uq2viZ1fXwLTg/d5WCLAZmxg7pU5+oE3ANkHq+
l4oEEA0qsJoqryzubU/+9m9Ts+LFm5iJiczrvLg7bfBlslUUAEUcXBJ/MmMe
Gdr5x0OqIJ9wW/s4+jq5nQVlkud6PGLp04bVPl3P2R6jSAWIQGZn4lqqgh3E
lcp6lMmdP1CsrMkNGN2DoJ/6Ye8LN3xohAPRqTOM9Vdgp9SH02DaY3UIt4WD
vpq9MGltKAkbuZdzWHf1CFtpiqX4TIaKLnuH7lQgssJUed92tLxBEe84jetI
aE1IP0oevNIOfbrpSiafnvXJw0z32rnY52Al0FYz9dYy/9RrST3yJ/8ynlI5
O4GncxanJxsvF3nV1VtSUS4tKW+Old1iKt4wsaaBuiVl8dP2V8V+GUqar3B+
Oz2RQipcKBMR2cjuKBp9kmdZKiiNCCGsr7Uv7w2e1bR8UNnDN0b5wVfM1m9S
c1CJ7xZfZNMZjByEqAv0BKfwzCtfprfxhr2F2G+uB1wRn0c+tLMksfAwZgNy
qBa9GYN5xtt+iXVMJeB15rY8ubFQThNKmElUVsQKWpptNrWMcUOTF1zTek2m
2Vt0JsSt/cRGuTNSq+Kfv0W4RiRaqRfU2vsoaYE0EPt7pJZ84xUky4o1h1ts
wF0rj23DnhbMYksQKM3PneE+o9K3r9qJXyYwDEsWG9XvWsmSbd3hetLAJoth
sJO4UF5fUS+s7BsGxqyexJyqRKrdx8BWv01meLm2W8GPs6brgjCrdKKnAXgt
Mny6jL6spsTcdlmz4gewr3j0E3B0iicUzIFdXrCj/s+GTQ7pLlABNAfqE7yP
NkxeLh71uh7bqm0vLdNhz91kJOF21yZsC+c1D0vGDChjaMmKf6zFvUiKqL9v
2n4fDPsdtv52BqHJq3jIwr/a5if+ia23tN0KWPRASkm2T1JyeHceNraP5V/P
Z/xZWb/JopAr1BjXbqQWwr+AFth+Y3poybXfd75lorvYLTc9LDI0EHhbwwgj
k6G1PKVNkPn2Y9oELUJ/NdwtJNIvlT4xhxp8dht5F34f2kcenEi0oCKq7C7b
Ud6dbxj1mAxXQyRnM0CY4//vRCUUqNBIR8gPDv7kJdwW7+nnsMyXBrxIoAzZ
kzBFTyUbyfPNxevW82UQMEtCKGJ3ttrywL/ew38zEn33FKdlVGowFlj+g3N/
YOzUxcn4ddBoVJ3PPCaSeB9kZ9TMdspyYkHZi07PXi5nyxHkwWIIuHek9a1F
ZBhmZgz6PwnVLX4pBRkFgx9I2aXuiSRgNLE5Vwai3+DJRldo+hgqtxi4wD7Q
yx/KNVwAMm/4HExE2Cw/JnQkmH7Lip97fRkdCF3tWeAMwMpJiW2KRUylJbCn
K4g/O6RPLKadtm0sh/28zPd5k7t0yjpX1I6Qc6G77+FK4oao7cZ0HiLMFJeN
R6pjCADzLnywRrPG7CMTLBWtZ6JpK5TbDiCzvn+M303EG1rl7yC/iaZteZj5
o10p0rBsS8/kmublxWy2bVLGdf7DOm/3R8wI2nOmTxGpPjx70yIFSqA+DrZS
X5/k1mbTwfwe/UhMziSoT7hZyXK4l5+StDYTQ1Kt71V/s9aVfBivhIsMm6mD
SN8cKRbxmCYMWBDNKhdgdLOk+fSTYzSQOiLNNBvJyUItUn9r3KsEiOdQvIdt
s/Ewq0yvk1FJLiWnpjCuKReAJSoe8mk2i4WDiXOEwA0hm3R3mlp9XozrX2AP
pkUTT+tmc6U6L6Dw+rF6aeIf+TdGDfxd+COJKCg8Uz0EvxvK2vErLZ68/6pD
X38YsoCk00erOGQ38ceE1K7vV7awZzahOHxZFHTCVVZ4mV50EuaY3x+hvzl3
3pPQ7ufLWpaoaJs8DlhVQo0n+K6vpP4/19AoDiYOobqQ6GtXQ5ngwyn2xE2F
MyGCZsGeT35cbVEOzcfELEE0EXIyXmdmmAgWBSqMUARTaihfJ1YkJJ0vG1Ml
UCsjupAExFbM14CLA/Z2NuB/c9E8Zrs9F7lLV/bzcqnkTbxeKBVxiu/coHir
RMLXqV3ugzN9UiiPpRu7U2oT6G6u0/hmOOjobk+39N0un4ygo0UfPI84gI8t
ull+hjPoVT09uyJueUz9i7KQJa1lsyGLgeetY5sTNlYRG0N3KxO8+uEL4WzY
FHbl6AJCC0rxRDPhjbLPaUW0twqis7QlyrFpko+mB++63Wiyo1PsFYcBLTYi
X2Va3SctxJTDF0ZU5BMkQVfebcDJF0t7F702YS0v+GA3lCikE3EszBO7pXU8
wukAverlYUQ2RFP63PrD4+DjNB9oxr60UqpqC4Tx98CRDIm8M+TER0nEtGFh
IV+6diE0bMhmcIZuMQEny2d2JITm0S2Ojyf5eBp+Fa7vni29VoBsC90D76XJ
F5y2LEJjFAOxmb3EUclbWGagEkIzSm/fYKWMFqt80LG031qaGSvwYLqY4A08
3c8ZT5etOBjEn4i2sDPGhX6P9QlXs2FbXIRyVcElJp/Qe0QAi7lLAzUzGQgF
Q1gr1AcyxwmddhwIRq0R4elUg9Q0viTEVf3WjiojcThgP4p3zsW6KVh/f+Sr
0oGvj910yF6oNNA4nf8jl20MYBYPOSJ6tdTO7Yt9rgPEN6VFvzR5fYzKQOkb
EqpJ11bFlL6OEvrd3/oYGN6grlw6jXNE8sdorrgw6wDd0XMu5llemAFQkGze
yYqXiZ1IltqRr5tuQKqg7x3bjazSbzFAX9d/vSoXbTzkn/6vJkvMqOa9SCEN
stpFQ6Uy82CpXC+xbyCsmsi9oI5qaGnq4rvCVjCAVecNUjL/jOUMg+QQ9wQP
fpmaPNqNrb5tm/n1owxLIEA6R4NJh9199nFFWpObLZJQjpf9ncSTQmJ8A0GG
iHhlXBtU3s58AN9aVdFK9fySJNtdHmaUgtc7U3WT/CVxNLEjYKfxUVeDE84f
sbN2Ki9sDgTuMHZWHJaZgTfTShfdQJA+jH/cewwH/Ry+naL4riSXM2kEvIeI
kZhMvFEf8Xu+Luc1qhSqhe+HkDKQl4FZmI3zCPhukQzQDJTUHBmGf4oIgw4/
HA51oBzKy6Gu7aEYEGVLHdQ2mvllF/z+GVe8KHjHvqim33jKWW1+Qwf3/fhl
GiWuRpY+CfaH30wYiYRUThWcz9arEDOtDFVMaBeEbiRS+kyNoGx5tQJQk0/S
E5HgWLU3810LruM2mwkpPS38N2IcX65FQ6fANnpCy2SIuF7FsDxJHaLVIPPD
FLygdGsaHd4kNf4TLqf+bLkbq36RIqvBd3JPHQENJXtFzArMQWmrI5cL0nv8
U3ToTIg8BboTRudJWufYXTr6mcuCmsnd2CyOqFde38Fliqz7wIivy6iKjjFY
Jy6YGdnKU9i4yj+o4cpleI8wFFWvEufJX8gpPzJbrm4dXCWVo3zuSD0f5w6U
AMxQrmLcbKpHKgvjZTH5dtHlbyGR3WbXe/EkU4AOYE3o2C6eHj/x20PEre0e
iwI/jBJIxbC9zjHOUNNSy1Kj/KdBCyKFGnxPKwcONOXFt58F3ZSd2H6qb0tw
udIxwkaaNXoR05qnf5x2sAqNIxEA265+V5SDOUx9/w0FG2G46ly9cWs+lbIr
wovJ5qtu2qvjEyND/+LtgWnm+DzeOkuhuAitLsyDZVoQq1KH46mzoxwlZCGi
iPTKZZaN3wec7nroF6Zm+qQ4bEn33PpxT1Y7R/37RCJLknMcWBr+/wkbK4/n
0O22jpMgdzgDyR9npUEnWPhFLeo+gdsuC3lBZBCyMKHyQIRkF9PzgN6CrM5t
m2I4gGPZBBNy6wrfbeenrmHMiy1yvhiLt8Vv7WTI1xGMFhjtwESp9pveTuF8
CoGblTQBiCLt5tT0c+KgbwxUb160HqORuCT8MjUCdyaHIu1u2s3tAELB7Kw4
HqSrikO7ImTLVALoUoEWKYQ+M5J7tBMpPoLqrlccpE0Pot5+tnvvd4n4tsQ3
eaAohRlcQPNqATXTRPBw3H4TkNGYc9ME5zTwVfpF68F6E0AJ4jI7NjDhtWyn
UgTcBIkyLTBLGwnzFZnRiI+0Ae0dHRpX52axIVlR1zal6U+l3DuA3TeRwFFw
kWRlDASjJStX7To6ccznOYrAz1nz+1DUcsuY/MqkpIvNHxCA15u/z+f1ebQt
jQF4Hys3lG/199pFMJxrlhf8tE5DMoMivKKMpUoop3XF4MeOZrrYqE8b9UVm
tjZAN8J7WjQNSu88DGU3VoGPdDtj2728xvLiku4/TNR3YPPHOaIWOjwYVFY0
dIN/xheKZIQRZ848Mow973HSgC8mrenK8UxZgzSLgNhxSPnqt7z9m0wIYqm5
OFarJ2ssqtTj6uLtLrQ6xOQVVECJByRvWg3bN4jFE6++YSmcvpmxuosZm87h
e4eGxVu7DAx1y3oVArE2BLCa7d699owuNWSL4TIJTrMa0vAKCuCGuMhL9PZl
Ogq1G/WIou7ppbfMhVHn/dHlzCWjC5NszEiExuXIOfvvllTHAM7Yzuh8b2Nf
wHLZi+3iMtuI8iOjVvpHi2q22MVggwSdveAOKweoGwYZaQLeJ1M7Iy03CkHZ
KFubykg7BTn3lJn2BHuUnD3UtsqwuznIf0LcXtEiRRRERKLP3yaF7vzUego4
sqSHz8TiFPvjNlew7yqohJfVAsRQI/aH4pwlO+vYC4gk7gfyB9gcZHoipMTl
U2gf8ySztC/V5vvs7OEZ9tY4Sa1x8OW88QUMj/Gsd508pmIs0ZrsG/BbLFzW
dys7wUSa9oQ250HHEVYmAPcEGPLMwiFbGICnzUnNp62q/IJENuW6QdWNqrxr
Q5FXCga41hZeNGGwET1SGrrCg35hlnlTg/UdymUz2+201Eusy+AuuMrzrU7x
8mfEtA86AjDrrk44Sij7lZpmTbgd0SgcVIn6n9GdotBO8IUeCc/7nKUWeo4h
IeEhR//ToFYnjJTGluLq+cc4pVB0lvBaamarpSI1HasUirQOe8610uaLm6BK
LfxQ8YdaNybeFeS/k5ryBaR1PK3wIa/95lLpsHOTNVAs08RmO85RURHN6EE8
c6RgE0pJVqXLmF5SaeH+OO9iTbZ3jsgmUj/uOv0OxoUaIjOwSHnMh4dNV7/o
8MT993fU/HJKLnFWROR4wzjrK5aBJHPiF0A2pftuKg1b4IA+VzksavjmGKiw
FTXa8TM6XkW5/yo0fBkw2UaTayJZPwdLA1ZoZageo9qp80LkSg0wwyUSCFMp
/iPnszDCCg6vmsC0VWYAvuzuPPKvyOB8CE55ztGsPmzvOWt4DpgG+v37WtBs
jnkcqezvYqFBBe4bUHRYzcOonk8LJP7kt9EcEft9Holdxtob9kwHC269noK6
bGXTmKGVcwx+k3AlKtKG9pPhFLjRc/S3Y7Xjfbeb52yadmpPTlljSU+6iico
cVvCr4VLg40z/Aa2lvY0y56nyj68FGNpvKG27I9I2IDEm1wHmi1KfO5VT8BY
ydO78jmZkwyDEF3jhrCqjzvfJt+1m2JXdN13rQyhz+aM9SXKSeitTtTJuIJI
d1WEwQ0jkAMgxXefY7Is5/RqDMfTuMY++8c/koA4ftazbXZMmiULQSCFrGwE
McsODGfStZ6x/BiiGJwSjLixJ1+IJIU0Tmv8GP8vKi3fr75Uuq2D7mq0k4Nq
+9eXZ/i5vzcNdB8NgVla8Pkzkms0orqHstn/Lpj2UxWFavRy3eOcWz6m1hnM
xZ75yT0j/TF4d9SUVDaZQtSGOGlB58pV+g4g7C785VXoKYNCncrnGdeYXeVJ
raqFUI2+DyMBIR7EMpbRQ6LcsJg3n6vfKw8bKlFNuf0NUAouR67iTU4jmuAG
00jRhRzXk1k8EEdY+jJ4a2HCqUJE4OuPYND84EmWGP0aIgNNdWlM3PJqNSrs
qa0VA/z97W2zWYjRUVmc4jkS36qfbJG7lCNJnj7uqRoHO4BLNdzJ/JGk1ndF
xMRHW8Ym3xzm5HKTTOozr7HWhs/ag/IzbfzSiHI9eO8HbMrzrsHHSbfbj9WG
VGHHERESuPn+zUnIdNTJrLSNJ7Hsf+VLnkVgKF/QCz/APYl77TP33+8XLuTu
46/qwO9Aq0M9/ee8QNr8swZzRgDulX65H8TSYGw7oKVy1rLUUqmo2IJwagnr
5lxHwlDm/lFJDwy0uu0eZpdGW2edCtfuH2D+ofJlnRUK3N3xqTeMIxM3RiPv
2V8blqbu/yKExSBVw0m7oTYPwG8BQnN7N9RvMjlzFg3DZFrTBNtM4s4LDSSo
r7P13X7Bd2Lh+6iTmpSpfAVDTwR7Aceg9RNlgtSRhRfpjnDj46EuS07CZBiT
3Cp1zgBtj24CkceChENCBaORHHeAR9CClCvaMlrmIX1nwT1LdLOkXcL9/Mlj
FDG8RPZ/Inpvi+2GNKAsukiSN71f4yO8CA7E3skb5jxAFdsjD3VFZ8poFVql
cmN8aKxU/UswP8bXjp0RnRo9VFLI0whcROAyjGwt08fsT6iGrsI9MmDjJf6g
YeGbCYfvcb71DTmhn9tuGeOmJtvPp15mjWC9biFRvOVnOrHDieTFTzCReP+v
5H+jFlGLNYuAob6kCiAONmo/4BwSCloyDno6U4ARjaZKUHxkaHzkXWzD55EK
CrvfM4OVUnntqlWa3Et/9q40Rwf0CeiDHWgFXOI4xNHFJabef1gCUrE0bt13
VUCQrlK9j8LsCq0ZiAo+ytPvt08eOFr3wMpL/hbCL3XHk/qqsBsCnOuDKyFQ
RidvXu81ktcXvcNjPRlNbth4GQSZw9v/SjQMFxMnZEuXvuCmVaaTerMkpCLI
StyWp4bQqbubpc/xKIeOz46QJoQM6imT5T1zvxQzkDjkU2ThBfHSwgR6VBvI
FJ3afzz78OMeCNy/hzA2itzlFmlJSZd/Nz6AQSXm5Qj0qgU/HX7fEmkVZAFA
1hV/58ZZYfhmrspqAtztFfY8DimVtcpquVzg7aindAY5s32PVHzfYlSWedRE
i7WN3H+Vk1rC3GjLkxyd9EaahXs4JjWkXd34eb2UuB4G/ZXUv/rvxZM8FdFJ
mNIEuEyz+DNrAP5Gr07ENukjigNu2atDf8WrSeSt1n1D3UKzL36UBZYqjwxd
eIUKoS/vFTxP1hkpN0nQWe5GSXMgO4SKGfmENDxjC3AfqsXM8Q5PIo24jUvl
5JKq+9LmhTzAGJcsdUESx682JyN9Xs2MZJbSCsPHY+5zjETsedpToY1ZZmFI
19b4D0SSLfRWBo+AQQyOWEz+pvgCskgma3QFMLA47EiJcbr73tkPrMuUmM8H
LRivrTPLMGEqNFJ/SD48i3ify7SK4fgX3Vq0q26gVeOonrI9tEIcxPgjt5o0
skDuDyMZnw3dN2LjugRsDoYPqlKiZQS1skbMnntFvyPMSpJB4UymAqFTuEDE
ecdI2RBFggYFU9jf7y5NrrTOHKNI9WNxyAKg4uHv+nErxi74xfotEzLmLaZ6
EAVFz7KmzCmAoiQ0Rm8sLR7nqCw4z1qXDX2t5ECeo1j0zJroMeogUjvhHL6w
kefg1Z25F57XMOzf98qh2vAeqHwSa5TYSKZHrlizw7Eyz/sNfEAr2ooMbU33
7O+EFnjKLBvh77rTQMqPEsWWE/QU3LJ+IZMOM17s+wfv7ilmMsX0IENecuIo
hJDJM9T1h9EaD8fDebcRrgdXA+nILODqTknQn2yex2RfvWedzVk1N5IEW5cZ
frPjwUn7Moa0E88W7IUshLBqLy1C9KtGTxpSi5uuTP8Gv2plpBr8l6A/Wv+z
/oFL7X6apQ+nFMLRb1EWnEzURGYLNgv/9sLxWZiT74jf+DlozSqiO7P0e8uq
+LlvcuDUqm5oUMqzial6wo0zg20lVs829BKj+emw+aeDH6/xjqjauDD6+9VE
VoQApGgsf+w5Kgs60STRbnDnRlPYaf8oXJHz5lwqqi47SA+1zLxPG3YBWNnQ
x5WNG6H8wHwiEUB73nYcRqW/+uSVLFXAJ0kMoUq6Jp12ffu5UEzKiVLT+Irk
mDJvKySF68tt/UZkEI4q5MxNbC8HYleqqhXSjsrVhd8IdWUrDd0sMttUOHqA
PlgInYgoJz6+jGzFlEmrBzF4KhYlLUPXZ5nQFBODs7y9MdnBpOn4Ev0SnHF8
dw22WC4o+Qmhsu97Nof6Fju32639U9IE8WZkEFnJKJeG78xKwbwurG6dGsXZ
3IUYRDbnGIDi6fcSt91jfTmIAGWI4o5UaP/z2KPOzSpJ3sK5pFNChSLYShf5
WQTxXlXTis2CZtDd0DvsfE+TAFdORvSB6Eo1SIZK+7J1IUa0ipvpDksznMZZ
5BhHuGnNHf574Ia5/5915Koeg/Md5TjC4RO6PdpesH7K3fM/pBNs5pd48jbm
J5g35ET01N7F9wrROooqU5Dmcl5QN3l0hbvCZl6RM7wQDLxSY4TgsiWkg5lt
L5k2TS4U8ImpZ3dRlCYA0a4HmgFQbjurfM0/YNDQqd0L6BsuaJiU6AKbziGY
gHi29Qap5pKNZ7FymIJ7jWYK13XHPJjSBv884Nk/Ryd52Bdi716rjeLA0SJ3
q2z/7nAb7QcWlJgEeQifYSLJOn4wfR2oJyGjSoBCLjPmUE1z1m6Vt4EH+yL7
GjwNLNaSZfLqwnnPURy3XKLDlelC4J7OhCqfZRamqec8yFOyuDSIuI1DkgxR
QGBh683jN8LTzgjF6eQ/KGDP6/8b20w0r0fkGMpWkdm779yqQfjdwdU/730Q
fTBDQXUGc69eGqTwNFWm+EXWNQwllYUyga7H22h9Ie2bkVxLrk9/mAXdEuUe
0CB0h/gS+1d4tBq7YwHQXN8T6koGtDK1sSo9AJO244vuM2CVz4ipGbXeRlHg
biY9uVFGw4WYMlCKnuNC2tzsBhHawwRnmxIbBdGe3KdMx37DccFTjwx5Omez
ku3pzxUCFoFHQkKii/qz+psu3LLb/ornuowzw96dz4TkUYgpDUDs2PEsZLnc
7a8vwgRt3tJhhwXgAjbMahqX3UWDO38vArawAdknKj8m73ePVIJDgrbG3tz6
L9tKKPxGgBV46qGsoAgp9z8dquvmp8OepS/GQE9J/Zg9b8wqIas9wIaQoQMX
1N3NTOmh/R4cqNBVP5Ek165J1R7iaUPmnTVdMxhHdev7KjFesVMKNNUYgeZ8
8VoKpAxFlL8buWpmhplaNrD8SX7RfSs7PdLzikZ6VHCod2xLu9bV1pW0xBog
NwO0PROklMLjLe6/i3LvAQZ4KpTZhWW1JqB6DPxPxrrtpGvgh7zV1vn/ob+H
UPY7vUU966N+zhs5GhrHZpImY3X1t9lqDN8/AHwR7BeIupXSIiyyCgrS0mmX
PqLZuzKB5d/AcPeeMvhMi99DBWgPxGn/ycBBxe+QecQi8cKG0iEwaxYeI++v
A6DocLYZxNEnwD4oo5ABIIYB1e/Q/O/6fX2aVAMyb1ao39p1CFdP35FXXsbL
1albM7jSYpEKBkd2xoMIqcKNIB4umot1Y+1BFho21TvgbegNftP1JZ6xu4AO
yPISL/SedERz7Zs30A0jAHWWVBTyoHaTVz6pR1QYqcZxxtiG/ffSnYqIw69c
bem7QwFyOBokkB+tDxggVT7mKwImIgYkqiC63t/8J4xc94L7FUFZl44PHYGS
U3flSxs0u1vKRf9PCSnlbXUTqv2N4NG2AUE5RZdBwx3ytZTvmlNpK2cc9Vog
QqTc7KTCO0fS1i85usaKSA59xiBbkjQGlsuOk/z8/BjmZVSfHiLQhmO4yv7U
hN2ouMFz1B/alUpROx8vRg7H7/d0dz/mbkEYz56ZW9NkHGsLe99EXlFmWOkz
kd5tpw20XQqh2wtpiGgvi02JKDlRjSdVyefamlYMwYef8ee9rT8DeWd6k5KF
QTRnk2WGGLZMWncrJtKT4OnWwn6SMG5KXlx45YrMIJ9iyp3QAwh1XeiM92IC
2QtWrZDdfglmz9y0pbm8z4nU2mt33CkIVWazcqbLcBq1XxxMrHq18xsv2YYp
2fdRX+ECQp5VrD9IA9sPGYxfEucmfoVjWyV5pZqXAcVSaTuT4ZMAgx5pqidj
9EGm/7zsHUicKrqWOiwkAbiX0LjEpYSbPevIS9CbVjqZGWX8fveis+XL+ZpD
WShmomyN+OhHqzmic0e20Ynk20z+jyvuNmxFejkSjvSrO/Kvjcm7va4LrLAv
PzSSKHC+7NFT4/8lxHk3EyPKEB7ccyjlcAiUCiKvdqx50uiT1I4IhSIg57Cf
+XH9BxRW7o69Ql1M14z8BNrUMbGuV5UslSvwMyxqIVycktRCoXrxOFg/fIhJ
L3EKaTk26+QqZMetaerQzxM5nvy4b/T7h3Zp8672OP/Evs4yTt0RRpuPSwvN
ZueabWH8ogvKS1goopUXMTBxGTi9wea+3ZL9e+iO0LPqfG1meXhju9PFxu9v
uBAGEneG+fdL9TF3WUhlCmHLiehsSLevJwFyvaLqwbwNmam+moC7aLDjtfnv
3jhW9gl9maPRmxp6C9zuwOo+PrgoraLNOxkVmEYpC63gYXBQYxP8GHV8buF+
vCWwZupoD5npGMTD1TXEmvL3FSdsLbImGoZIasLrn3YvZDbDrygMy40j2iIw
fGXwErEsxwIvh7T2VjdiBGk88iQ/cyM3sqIzxeulcvhipcZdDZkLPKeiuFPq
p8YPe6AN/l4draeqIl9yAdJuv8xBCIAsudR5k+7uGQYEc6UW5s9V9SbF9lMW
PrRzZZhPgAT9xxd+WaM6UFNylykIYJBElNInHRS2+RfQHbgir5Eh6pxuPx23
ErifzfdrCYji9VQv/SuNSEhKTV8YeZFCYiSr5pRi6euZf/w9wW+h45/2/ibe
GRyxX4kGQBiadWiDkmnGyiPlaDW5W6CydXWp5ctQZO1Q0wOXflLNKORbis3d
9bC7cneou+0sInG2CgA4RCbvx7MSfzOXLC2gG9WcJR77lP4Vs/GIxCoxygvo
irbZvlYL0WGnB+3C8O0TqzTl/pL1wdFc7clMoatF2+eROouvcHO0IL0KchHf
MtsP2eQDV/9OPxdIcxOm4tzg+aZk3szli2guppzxf0uAAjkGqPWrLZLjFn1J
xxX27+RrqyPLCgBQpUHqGWxvNDgeT9o/RbGm74iD2+WYU22UPh7P2h39vt2u
YFap7WJsk58xSuDwVC8/Roqvy1Q0wx7au2HI7R8kWKh+QRkTWd/s0RfUHYTu
QGjC7NIVUPkTmeyIMPvF05rLlsiJyaMT9/h4Zs0Hw9XBrxo3qz6nTQc3lC67
MhO77OkKyY1vuTN1T/T9szljo1W33B4KGtRL3z6tFmBo1DafK/a0nvxyNo4x
BTHXi4ud5wGS37Nb7hmIxtx81+noml0V3L4CYntQ04w74zfcpL2+3oKlZrmU
GUdqFGXQn6/14b0kY7uoMkZvTyszh8ruyn12URYSOn98ECCkTeIqCqbaA61H
r6hRyk4aC7Cq7JnDbXSMub2lNmsWBS/hrmM4oQue0e1Za9aFiCMZ/WjRkWpV
B0iq5SSvRo8lRcNUoosfPBbUFQILjSHf6uZpID77/uEpGYv6seAf24ZBehB2
9xRCHiN7f1DBRg7DJJcEbVjdJ/pU0os96+t81cNCynPE1cdWheRU7JswaynU
qeEOQw3AgUQ2pmXeJcychaSsq0946dBhlJo/el1HA6Xey3GzzDMgv72AV7gT
wIAKqPXdIk5CNo+5dCavflpynVpgQRgE77q7Ga+fj8APRtwhJDRPAY2vaZ75
BCI8Gn9XZRlAWir2vS3GDOWCtx9Atp1+HsxXHnN2v3nVJSwODToP7bUvaSxM
iE6tAk1HWvlj7ZYAIRh6xhCX8ZwBWK8XATBdf4OFVJNBPzjytDZInvaVCtLm
EeizdEF6QjCt6Q0Re3qBtmUujojQ8FSERLZJWBLGjuatW7zZ0khqga+E4F2n
5Mq7e7XGd9tOvfklZOIDnidf4sO6LX91TPW9f2VU+L/8X95cD3Ke9k0hx2Vs
WQC7en3XcDNnne5mPVhY9YLdzC63Eax2DAdOHnSfNJj6UfLRo521/4vPK0yK
iVeE3t2wXiOtwJUptarOYcaSHZpHAc6m0/su6Umn9eSDxTsczJ0Su4XgDikT
Lh/3XSPdXc3WKJpToQyKE1J2IrZGQiXNchOCc9/zuttBmcxTqj/wbehhDIZg
h8vC4ck14SGf1fQTjHD3ajcNpefmqz1fKClYjpHLTc6mNAy5Ada1E186pOeC
k5XC/1RF1ociorvB6YW2dmi2UGrjGputak2NSm5Z65hO8bZyTy7W03e6uzeP
IbjqQKe3CVOz99rsiMNwUVy6fhrb4cuUY5rLrasQiTG3vwbF+0sOmyfr6niA
XZuUzR0khsPH/g51ZGsk4mKLsYcrrPrm4jkqAcmgPfSOM680y4hhFQZGMQwo
rFbAm5n7b9Y8AGiHewiAKCdPUmB2DNd4NoXQ6h6GrlMcQvkGCAdMn/UkWAzr
HHUstPq66gfH7fjSv549UpslKuZxOa1GbDV2JIG5iFYSkrNpYRrRhZXNvW8b
qV5tuK9sU1j9FSuOKxjqpZBkWg39KD3WBWTnrW1OofmYBPNIXMHHboSy3Ps6
t9ikzRcSV0mB3w2SgnRfRY9erV34tOWonYe3qOFBKX1mb0Kta9E+3ctml+5y
WVdaz7RXZmx7rCz+OUzHioUJcGbTCMND/ksI3QdanZ+nSyddcX9DPCxZNKVU
PoT2eOZYH1MFFTMz5hjOf/03SNUXb4CrFd8NajJ5hnvGZCdxAYyOPOL+akyi
37IRPEVMI2sxDQDuJ9OPFXpMpQd76zBXGhPH0KpP2dPcuWZM+mdbDFN96RqB
UnLGxuSIYFCpC9zFWNSvY+NljE/Ece5DL9AxuWtn/L8XZcD89Gfu0p3tvEEQ
8qdLOao3zyj/+NjHgLd1LcQ1WdDFrZaFsQi/BKhRXnI5BcpKh0S+gqlE7wr7
aZwOXl2tuU+eW1kgsLTptcJ+prSR6O96BYvcY7o7IPAgkfdK3XP7I2AXsYFg
7XQhiqwLGmDbX9u1VTuiRD2jWNzBhMUDCqNtSLNIDhxkTFAICIvj8Bzx8lLt
/7QTI3WLD9uT/7gwHLYNHbt4j+kYshqacaxxIeb3S1WES2QWRpdlhpLfW94e
Ui3HXw6mlBZUc5Cn+ThAdZs+hUDR23j66wGX/F3Ay7tbIrcgspIqfLINcaIH
MM4uaTVaogM1XcYhi1dfKPD4b0C1DqeFalvAZI7eMOkpbapIdSBMFBokmaUK
e3Zigr/kI0yMDG5B+badq9+lyuWypkqdN4oYEl4EXWqI3k2ziah5isW0Y36R
s5kpEGdIw++nlCss01OAsg43hQA95bJycGt8uEsb62hVBbexUNusvSwzE09H
iU/aGEB2pGGNsytTI1R0E3HT9ubd+KVaXs+rbvz/DLaI5c9jWEFotUAnTVtD
0Z3CDr0bxk+4KhH8ir8GI8RltSkchgiI88OySVKjdBRA4t6G1CRA5pb6hJFv
lzFSOO2t7/vpfoGSlEZlWaqOvve0iw4Sad4BZCyB7b0RIIFxM6v7nR0EYjbQ
G7IIwsrhJReIg6UG9C01wecx4C/tcqh2QE3JzZXe9Antv52UX8wEhvrVs1Dq
wkuSA9th2+hcdE6ezPzGYI1cQLUB53z3YFo5fVzXTW48vyedFoxO4vVKj+dD
q7fX9PlwyB/Cx+NnLFM4bENCYarwv95lEs7IBzJHe0ZGGNekw55EsotwQMAl
B6RwoT0j5z5kP45udHvhQM7w4MIk02yP3ATE2kBE2uSTjKXIqzMxfnRLe+bN
GEfyGtY8JwiJvwTe8qqBs2lOQwHLdPQDtFPciHX8uBxGO5xfSjj+V13bAWTH
zcRdcNlZNW4IbrAP66NltxFiy0pRbWjpzU2E6e2tc0DEjuuRhLQunXw/8QhX
LLN91bJgzxLThQMSRcPiGlOA3jDDCUy3qpIhmVzTceZrYiJlWKxLqqc2aCYr
t5teEExloaZCcJIHgwA5N9OE50BM8ewFOJv5Hk32fJv0uP1ZES80OvVos2D6
+oXIvWnNM7iJ3wNDiKAyfFH3MpnXJ2XUdd60FWaHDlb36JJGrIKIHNojxijS
M/m447swDDO56t/3T4HPBP8n4HLzXiS7Wya6PRisQEVakpDpgAQNpZJY7jyU
iGk7Ehvg+LpytaTkgKBu7y4juDx6OcCGnbi9G2B/lygt6dqBfSUoRP0w7DmH
OXW2MUd6z6QkGuW0nVXr8VGkFYg+g3A3eLX8PzxMixXsiCrV0usei723GU3C
ej7by4rJHzx4nLIjbLJchhmDBgwlX4zk7DvAQWuf2bWWyOi3YZTNnxkFgI5i
m5xsGCNQ/xb/6YG3rvLTiBazH4t/hc5020tl5uQ6wgbtm1e7pdaMKT6fEVBM
R7eGUbpZw+ugtXe76HGOvYrywGayflL5JmLBHLN/U6y/Vi2jPCYiNXKUeguc
L4o8y8ira8FO25WFg4r4OZ5XagKzrBdE0JNfufPTWCnjPbXMZnbYEhigGnT4
CGqaxAXo0GduVetdWrJQgqwJXpMiLjjk2zIsjYH4RWmGa7P7RhE4kb9iO/5Q
NJ5nrC+UJRKU+UET/gUhKpJa1c/x6Fw23Si6DkuANChTi40mU8csl/fYyS86
YyyDDiNIaa8f88NkqIuOd7vOmWj+f/adpC1argiABMaqAklK6QeIhb5VsLxU
P9j4Ib0ctgVlCU/2QkQLep0xaGdPFUGvkCZYfocH5Q75lD/2qLGFj9610mt1
iEs0hAmA4q91JdUx1bWVrqnvt1eYZULfaViqtcDn2zSAEK8PNW+/m5hLyu/O
rnBiL84ls7IXlE54FDwiGxNbZ6hTeK6nO1pLcF2NJXPOeS53cShM/qTEUZTT
3tRWvu3rJ1WiKZA60IkhFWybep85JBiFis3EiQJLTSxJuKmfwTyLNscfv8uv
FB2sfyRGR/CPXKsswM2KnBZo5NOBJwGKOlIi60AAsICOJNQKs7neqWvasWlA
TvzFX8FceBki0sK/6OcvLIgDbknO4bSC3zPh2E4Une2XgRjD3sLkCGtV7DuV
O3wz6d2VcJ/s9Z0WG8+TX2D+6jizKordFyfeG/PbaoIuKWD9TU4Mq4P4+E/K
PXPUgFTTIMrxTVvWsbypZ1T4Icfqnh+e9g3q6DrGsXdLJf7xHsI9bG11lQzg
/ZUaU0gncWUe5az5TOhrs0hTFgd6aTuZA8pW4VCoq5Pa1NyMQMKg7UWtLmmQ
TUS5rjynVaSKLn0tahLsOK2S21lasdayGUriJIH4uIXTAV+cJemo2wX+4oAP
FTbWcAFGjnK+fPqmOrzbSUW9KNWtoSJNPYJi8T5ljhbDJakBw5ofP+UVSd1E
bZaBjabmNXgr/OZWMM2oXLuiCUHetpRjjLbqY3ITGY0ktFsfZ14IFlLMLg6f
pDrw1YTE3oPovKnCSHDqL1H8RZe9jCEpYv0M/LGkf8ZmedN3sh8NX9C6MPFk
pgAFflzEd3+qfcb+aKeKK8qqz3LXuRKMaqHC8Z8RSn1KZdr3ElnTjSM1v8h8
3R5LVS/eAXqNBy9xbBMLfkzBNMpZ2EkVw8qWBSt0qVrx6hjOeojb5Dt3CY30
T9pkkuUAfvjzL7g2ES6WXpklQ2qxPKeDsMLfuxzQ/UPxRmD8cUnxqS3Lx578
t7xP9HoZvEaIGbH+CI0371uFmXkUKD0hz/UqBPEeazzK+2QNbqxXae2nlNGX
HQjCu86T3le5soB+6Qax8JEi7/GMkA5RHRgs80RFWE15/sTkKjNS0zbv/yTB
GQdDp04gm0bU+IiAJeJwPJ2bTA8NzrHlQiD79dFbHXSfk2JeM4vIg9A5U5+y
tyUG2qLMkszHS9uE5sb8BP7FmbokiM/Nm/uX8HV9jNMUjW8+ZF9FymqzzVqw
BBK375hlu6EdkSuJUrG02DcEslTZIcKr6UbWKrU1WMNyfGx0zikOge8nmoo6
DOXmsiAOtfWQSv8Rm/bahArdyzdVfJTI4zP9FJxrWZTJOpW0tIwWXXyPTRb/
d4x+uw5yizys3GS8ZImJYEisNHEx7FvrERnWgIkK74hY5pFwt+atpe/Cdl64
38qkYGJdT+7bfKwuLaXmAuTIuASdJ3/aRum1Ex9KnLb9/9jT0p/MGct+mFhT
lDuHh+1b0WiWIgm2WMAcVd5RcQIOxHUnZDRMk7jyHZax0VV5+HWWjhDFsrgC
ym36xUhHfwvCXEwvrxLknvKeENuCrfkQpYQkIgUCQHu/fH6JeMQ9/U8jy3Qt
hHys58zP6MuQaCxba3c5Z0OFJBcGQI5d9JndgO8OQKe9bke4E8oKfqRLvyrH
/YPkkSyIvEH08Jijqr20aJeZbDk7SlD7d9/Ks6ejI25xnUD6J2cUPliSYT8X
mLQofeVzih8u3K2szBKtO22AGQnw2kq4BrjW/XDD6bskYeplcjiKO5pnb7Ne
fKy/9KymtJ2RCJGluT5Els66uVC4t4XjwFyDlsT03tD846iMm6owWOCzz0jb
pAHDhlkhKKY16F8SDUQLDqoAoWdRTlbPD/Jyb5W7T77wj3leZmhTnsVXAc6x
iksiOL71ZV+9eqst3+qEp7BCVajCtalioGkjf906ldv0FZhLyT0Wb40THaP/
SYDsZQCqj/vCWGOgOKmWffuSJ5u1PL9GI/w29a1Pb1G1FCgkDQ7+zDWaJ56x
fGTJbUQ0kjCJKbRaUsuVPUNxXl27pUfxBtLvrMnbpP0lkuwdxR3fsenQI35D
UBYMJV/WnyTaBechg5SSCikNslBlKEiNuwAkiQBLkVgvNbEWye050iN9QXqL
FWMV7xbxZ8N9zcakU7hmqKmrvXSU1emnFBPBtnb1RHTpHskxpBfBE+0CBIYV
KttreLD2vh7gVa7d+12veVGVHsIpXzIx50vBZQEP4K7+7GN0RumapXnU9CZH
yHgZBD66fsWekhvxyjIQ4GHAXMSBoKPh0RXeBfMucLgITuoLMh0maeSxIJnv
ikU/6jn+dl6gUqjtRf2Ku2KisYKCaDHWolKPgXWrpyxY7n121Dh6jLugI8/v
wm4vGROeWb4eQLd6MEQM3ouPI09SkQqnNxNui/+UWg4plZv/wn+aNU+V1k46
ttH3Z3W3KTk6dcdvWzLD1c5qbukHK9LGsS5+LET8ELBQShscjswmzrSBlbNs
MzXmdvysf49hnwxo5+KTpdLjX3Cufgcj3tSb3xlvx/cfdXndnKuU/rAHDMuI
MWuCPxIx5To0yB/5njVacJ8XIzWB9CGLFuGhqpQDIYMYASmBmEjHove2oQ83
ykutwJziOaHrM2Ypcgu0Lq5uITSr1LSM037ngAWAfuiV1LTTgFcUuIauZhtk
mI8YjIao6BtRqb+udIPwya1F1KihJjG1tVrbD6j7K0ggygakIGyg5uqXWV7F
0Uojz/hz7wiTF/Ktk1g3UnFW+cFsOYLlFx/kH6etMZh9wlSwy4Zv5xEfzane
5UEUr73Ajca+MKYsmDZJEbqQqYpHJ/4yWyOxYld/r2OqJX4WgJ5uuokf22lB
zYd/Br+4gSxaZhreGHqljQk18wL7s7oiW+m1aQav3zEkmI0t25uvSpqUutWZ
XkYapwX/G5+vpwK114wfGTcQp3jS82lWrlZDlYO7Gozu5kkzq6gKnJLWES3A
1ywYnbnq76u7iA9X8W6E5SJC4Pe+x83N7+8qdDukONq1Bo0Yquuv3Sqlhuax
lIqIJ8L+m5W8tLGT5M/wbe4OIyPoEXXnXZyYfWf9YfGynKyGo7LDGr1a1gm6
vocr2tj9SMYrhFKfIWhw3gEyEk9QaxvffmdSzQcnWslYDwQrYqqTjykJsqbN
ygX7N9TN3VwK9g+fZsjr9+SBTzpAXN9L9+h5ykUhuTFKzDgDejv5pzUTuo3t
y5H8WTcMf8bb4tSnGhcw/qBra+YKS8ZsqHoeFAapO/hfKB/lIvgow1ULB2Ud
XXj03vufcQHFxC3HKhwcrGBoJsvuVDPy5XVy4L06JlJ7QZNbepUvpUIt8Cw2
AXBGaZiNaCoDIaOtRfdjlhZtaDpdVW09pKtPVDETpnvJO6t7B/Ibgv9pyGRE
cSymIBauw9zREQAnXJbzxtJP+KH6wYFac1FI3fiioJPZrmk9ZowaeP4UbcSm
SKJgJM9b7hB6sWeVDMZxT5vB+FfavGS+0Yb4qO+LGkaOB8qLta2s/ilpF89S
bs2yG+QxkgOgB2kXeHQJv5RXq5ceGBK2tGNnomdUWJuSXyRWpm76mFPpp0mm
oA7CdSPxp6lJFHfsa6elN3h5bs2c+TWLlrZgCKJ7p8iwt9ME+Ry8LonAafE1
du7fmri2S+nTtR3kXBzlQYtYEXN3LShpEu17jvpVqG+CVvnaUTOmdDMjxCKc
tPEDrNwbQIHodmk9gBRAB63fiBit86j+182AfdRo5GKO1N7Q9hwEU+d0GE0N
bRfVXRWqRTlL658LDyKwdCg/4zCCAPP6phbx+yzQ90rp5QFaWY+iNQVHRbQG
DNbolpK7DlZg3HF68or9jSpO0uOEYlpKP/cdw18a5abnS6vMgeeXSoeFnQhY
cTtIl60ohdVoXBxYE9e/hnbWBJXz8b6YKCd8FGAZsSJvLAOd63YTuvOBHvVy
Qh09UdQhJyS6CFBY17kR1ivGsw7cwdVX/btnBHhVH12fzcBSnVehfx+7NTbA
tB9/vw3vvZe7sCyI89PDqeDWWqW03IpWeZobhaJZeSjEhLoMQsQDrqNYBDhM
x/N90ecqKLsMq3ef4e3xlEeVKzUrnCvzhy/xn+Hzfog3XCXe8hCO8rKgwe43
mgZ0Xc4VBwpe5d98E1Er0Lm/kw2gEu0+KIHnfGmLk2E88ba5qXXDR5IhYloK
xcYcgwGYGLkYWVy0JGVjQyehnTKVVy71Y14bsHKO0jH8qlQOlXtkXA31FG0Z
YwUB/AOQXs3Ixy6rbSGJcu3fFk0djSy6LNMc+Iwt/hAzzmSXFAmHDzT7m86v
CT2knxkjeIuBUOFc8u+ry3gZz7EzBGh5hL54cwfDFeq1EWNVijbzStyppXYo
pe+GXAJTCdawAtMQGsI26VlLqSuwkpsJsb0QY9JAIsbhVTJUvcRckN9qpgDf
kwsMm1LbbRo1lPG+3mQ1F51yUBbEuDVAVX5M/ISc3OpSqyHhAIaUIxwyi1sn
+tLUMfzaPmn3/YadXn2EYRm59a9qKZ/94h06l7yz1pnvvrMQidIkjmVgvE+2
my7ix+pOvqNZjz8MGvSvyW+0b5UrC7/Adlo+NfhUrfx9NIqE85LHEIU1/lHn
4xCYSkmmmnt9TbBnsmZX2GapgAaTzcV3tMyT8XmBzsKrOIPCb/4l014GhdM/
73kwGyA2jkuqFHLAw9Zyj4aRXVAbGjSQoEUwzQcd4DUwqKxEgsJsG7W2cUrs
EB6Se1taNl2YWVu9v1Jre1j0HoQ+siF226V+hCuFi0T/zee5yeALeoVGQZyw
BDIzAi251kWagcOu7EZfYml03lbbqcOP2GjnsJg6MwWYaH4+1OsmBpeFrWmD
cqAOneWWAII57ltPK9hDSktkbqSb6XdPcSFORi/Jvd87bdXolLGWU64WGyfS
JRNBBnNu/30rE69jr1XurpbyY8rbxoORT4yjxfPMSBLsEHQdb63l93z9NY4y
Foi+cp17N2xUbtesSnMo5a5aQpXqSc/m+KQOqQpbQfy+ipB4kcAkAG4l3t2S
zeE/1Wls/43aWH7Wt3M47ho5d3kUUOjpBrTuPPtZQcYuvNh4V4LfzLxbBTrs
REuNUOnQyeBq2rTaUAQLY+D9bzMOZldd66Vp7AGc4i9CYBmXhG3u95JHKsdc
oMPokgR3/93c8MNlGlPVatce7i+hQ8E68hutmaAdzD/DPsj4l61N0eV6dPfK
4xBiFN4LgB4XbJ1cVi24eZYXPTQ0LkmwvpLGLOZhbKry9DycaX+rShPSOcrn
ESna5rscLmxYn96hw6bzM8CV1zfLs807U1+zuohOlOpzWnHHRXF8qiAFji0t
6QYcX+cpW1hwZocXDGcEexgB5c9EUur1cPE79H/88e1t67pgBPsFKgJ57xtw
Kg5s2ZYEFIvXc01fzjoG60a+0BiURFWAZCWdbUOOgPPwmmXg4MWQBRfM+x+C
JkKci94/PZB/CZ4x3Z4J4pqNgkZKmSDeokc9wq9NHQ1Q/R+Z5ZPBuA3OlOnC
UZgNRogIuy9zuTAoNosDrEBDXIF54YYIh2GD+wTur7awHL38ogZADUS+AGqV
ylEJv465SHFF3wqdBIGmCYb6jlweyEiZSdEgQRHWwQ51YjH4alr0tsdIh7pZ
o6hiooCk9OG5MJKlrTs05U2Smcx4f4cd+PauLeRgVzoBtiwojKuWBCwj56mH
mS5Xc9fC9m5fgYLg1viZrPZQffoZldJD//SXmGwXu9LvxChtrhvWbYhHnPpg
GYytcw0ldCduqqiKGLXPCWfw21xjBWoKRGor8tA7KxGKZX08rtdYgIyZo11Q
30TiFUhYagA7LKCfZVcCB0E3zXUZcu6/4js5LV/M989OE+jJRxn+viDAEjWQ
kz9gd1F9ni8Ay+UhCSa4M54xid3QhJsFieC7cPS0CsAWm8mGWmUI8lKSUiQi
EIdnRAnb9qpdTrsA5TS0FYry3nZ8iSc+rDfc6KzBNIUNmuU/Keu1FSrPNqO2
hFp0+lwP0v/MmKWSIDPWUgnF/PO8yQdbJ47EP2hPsWmFj2itDhPd/3kepWvn
juvFSVkjg2Xfw9nkwmOsn+dXmiuqzUEtJjOMFQKcN/34erp3Z9jhoaNQKWl0
GngGivgYXZ9XrfBzPTFfHkVn7BXORNB5K/raH8+xavODQb93XyTDXhMCH5sq
oubBfl9YP8eQV3ncVO72qDgzPz+EiaWEEVUmCv9/Saw7JScisCnA7JJlxBlT
9HHKRNv5WT70avgrIhTL7VaeMCV/2OcoLPagFfVlkhGAv9EU+lp1FgTxf77u
KoluaNBhNQyrcva+4FhuLxVQuaMAOlLSwbPq5g+6ZHzvm2IlkAKeN7Fje1/r
85yJw4Hjo5Ag8WoFgZVuixThwb4CU4Wk/PuLXWk21HntTGjlHwxL+1eY51W2
wv7pes8aZqeRIakRn/s9aCUM+Cr/K1nJGymXe7hQgbkTsyDE9z0N2KVWCwyD
ofPRqGWosFfoHxepEMm8qS4x95L9J7piWIHxF9SF+OJp4NbcJ33vqwQ16OyG
msq80pOB8xvKyM76Qk/c0s7GOdejaUibyR28Rk0wZXz77RPs6alUXT8ETczt
YZ6EdOXljRYYIYywH3ouZ264mWULBoQ5NXZktRf++TcNugcJcWUxSnkDF1U2
W2T0otjtYCmBxJY1W66z0eAKrc3nS0kCuAGOXp6BomJ7lFOikJ9Y0bFUlayR
CaHw/VXJZcfPxktU4MaVz8CkOFWU+lSbu9keWP84ZxQRjlq8KgIlX5+MHyvc
4s3k7OrIJtN9dq834ltiBbZOyFYqIFMgkw/bamxfqJ14VnWjOy7XujvXmgqN
QHp6gjQCh3TB7L1jTFfcCQOyLXs5VV1Mpesw77U7L/9301U98RWkx15DJXid
3D7MbaH3SLxaI8p9ePFmwT3h0aLUbd8Ip8TJ5TGfn4ohZmL6m8xwikotunVG
TY07EQwzZgwB3E20vhJ9H6uTADqdAKrb017ZuOqDJftJvJ5X/wClff/m1WYh
fv4U8x4JKfDWnkCAFSWx1igGKyZKJ5TzxGjrpQra+yRA91suSaR//hbVuMO5
oleB3psHx3wSvfamsx3n1ssd/6Rwxe3qjnMoPt2q8bFLZJ00pHSmYu3VCIaM
MrWsiAcFrFSlv9RsbZdEx6aq+P3g/5FkFQ0ZJGXi4S6Is4/kVpEg0pXdSptq
QfAukkozILNG8Zio9yLoOv2tmPdS/4ej8DZMvhfvb9DcNbqISh+MLZ04hT/y
i6KJp7lG3+/h3DsSanj627g+tvJWGEuMW9ZiivSbXjSOSo9iXy9jKXPNJmvS
M9dZC5YS/XuzYXbI7DDjE86wNxUhN7NWEW/T4oE2JiNbhaIgt3LUgsbfDqga
XsCl10HqvB6n8Nvj1UfvnllDCw+cdlWAp6FxiX5jDDnHknVQ1QpysCCPo0Rd
mpgUFZ+L+u2kTKrhWl9KgmKx8cBj1vZwawwuP426i1KYY0EYcAm2rpRFsBQ1
Mqs+JtLd2al1VIa+6Gn6Zfx8lOWuhyTbAbgoTFYlTh7H1x+k2YGhROeknp73
RKoec1IVAtI+RQubksNQ2BbUvdWEx3rBT8haoOt7fQ+8GU8KCAgaUO1ppZDy
Q40OqC86sRk1uOhPmvEjUUCDleoXh/k2ib2GNyLPowlQkt7BvsiBP81lkUoa
NMeQfjz88QpggwnLSJHGnVcTtCSzfP8MJYmeSsgEjO/cg03PYk1I85B4CwBN
+1KJgGWJ6TYnxOXPz2g9hRwv3utFGPLBUW4Aq+fh0xkeD9XqL87o3bG11hKF
zyKpT4Dx46ObFOvMTsOUQDIdV4f8YWF/6Mewe55tTFXy71cRGDZZOQeLMLhc
3j9C3swfMeViYb3Fu/BgVt9lnbcykcJHjTEwFm1dUPuN3V0J9FlIhmJwYmBG
8lV3SeJQyntBz5RBg2BQsm5P4lyMdc6kc97xpwn+F6kqOvflUOXOjP/+syzJ
zbsI6iZoJ+wks/Bj1HZLL/Za4Zxw2wYtC5elAb04IuZ030MfDTfNlcxJqjtR
Qh6oG+KFcPSeD+TTdw4Nw/gUbdngmdV2WzGHUG8HezInRQXIry9TfyAgXY4Y
pmrxZo+0bwVJ3vDt7e1Iryl1wMhPUggL/ZppDa+XwpAic68wLS4SHV0WwiUM
4JtAC46BQlV70VLcZLEZ84a178F4v1s3AVM6lkhQcnrnGcpR+QCkddLtfuHH
y4Lw40MyJnYH25MI4h5jVVvYrPV5ELlP0/BEX2/jyo+GSKRl52otuXzhsBl2
niiGaU+9vsICon35WADXIJyuupKU9zs0I7iX5NxcpB0TZqVwJoa6VTeeUxTx
trDuLOI0OZr5RC74avK1DRcD6k93iORyL7EKM4f/TipXp9T171zKJAKXfkOb
4JLdpJ4+5hbShxjIY0DSy2FdmEHgU9r0jlbwQ2cjZJiMzpOZeYq7cpc4xpqo
dmPw2hMJyyOdbz+8amGn5mIuuy424Rw09q60bK/AeE0tx2dF36wrKDZiNmC7
Q2A51QcMoIQx8bwvLTsd696XvyEknZBIB0MKeZQnzR57rJOxoLjbOEeRh7DN
dR91D8lFvCBVpmmbUa+rPeiiV6iQrZqNFs3HoLnj4a3OdA1gjOk5arpxE/dk
mRCcPjUXdagz34xmOkUg4OZccihxR50OLHKhtXN9R0w3vIuX8m+3yyo+5TCO
ukV++igtUJCAMnn9FdudbpeXYL//ggWJ3HBO+ZjjPzt58H/mjZ5b37TjcLrs
f5AmurqSKX4vAYOpS4QejHjCzzWIDa6r0jcXgKCylfq9tvNUcCGBaJd5wZNs
jSkQScgciZYPVBZnMRSqGCT5IHmftgN/eWRi/LTUxkDWU++JYd6y/wV54c8f
o2wveseQ9WNOxLfDquSgB4rom3B1yhgzgAQTXzQM/Io/2N7uSewJ0Pofb0uh
EvNG/4K/ciuvFMMAzA2WjBpgAKTAN3F8r2ViSUQqZDnJwmEFg/d+IZQIZr9d
KGG0ALOY3zVYA+lgxDfheAU4OSFWbC3B830MaIlVHGvdT9RQOs+reklCIIfo
nicma+Mlx0ON/fowwr9DyqgEIocp640Se8nEdjD/k3mdmcYIYVgUiHGwDIcU
ytA/RgSnbPkr9j2LtEdbW1zHIY8tiWAOp4Uimc4ajuNtnyv3Ah2DjGDkO/vN
klIBSGUquqIvjWrVCru4P6gSKIybloLrHu8DeOl8pNRjDEMyBhP1hpIxMNYJ
WoVL8z0gQ9gW9HuOB5fhOTFeL1wAqzB+Fy63FwhG7oGBtDKHq2R9ELN8rkhG
yFiOTfzXnW9EPvlJQwnEsivtoa03yHf9FiJVOoRHLhjZnKxfr2DqiMsk/Ojn
IZsdmnlYOtPi99ieM/tBy7Y8AJOfizfl787kdUyQ+FJzKUh0h5Dga06Et34p
4ooGNXmEAa9li27Sg5UCVElmURbUqAgkAP35R00Ttcy8Ek0wXMvwWIbtGOS3
nf0mCuP/3oUeKu7OfK6DLBl29iNi7FVYaKq73ly9/wgXZ5a8UJnnF2LWiBcZ
1HuQfAFibA8eNWwfYoiAOhzvRkUKoiWj31Pj+FtUh+snlCZ/9zEQNAY+k3JC
yZHe0uzWtLh2nJOBILJ5qBZ1fdApssQfQO2LSoGfFuFa7MO5WPbYVMnLtfnh
XawDXSbgu7p9m96dZ5a74v+GiRNgr8QYLTanu9ezfJNYv25JW5+zb8KkkTZz
qRz/PV8YynqJzk/H1JLL00GsxxDeZWlcON+m0bhBtmu3TFcfzdr+HmYJC7Of
kuJxjKs2HeQWM1aH2Vuml0rgcD11gl0vCxRMUSDje87gWHxdfHMAeHadHJFD
XIpkBuGerE5JLv+wx07gQKBt9X6Dn6RBKEGKbUDxvNykn19th1loTn4sgtwY
IwNlc+00BSzsVhm2HTSw+6azwP69DqQR9kJ3rAtluJwHNFBPiSEJ1QlKlY6R
IiPvEH5ck8RupuRilZlzqmZEn7nhnRkkDSQ75d2eoWEDFvB5tVMf3G0Mj9GX
ZVR1FvwSbTQNCMDFNauyzCo2eLK10SuJCeHEYAp3kcObjHqfXJWdKfoeyFaC
z4BxTJEIM2T4/JQrmnfx4n4Rujnexg0TOJkfKscB2Wxp9wHjqKhUJCCpWeMC
VHT8vrZQbLNlM7rCphRdfhNnWQq7x3P8GsE7txk0DeU7OstQG/y1u076Wr44
gPFBwXA0FLVKu0b4qDAmUatzJlFoeuH+2PTb3zmnReWEvLGgPihebBFMd/i6
/VyeLSijl5s9jIA0d6eivHYXvM2YsurPZqMJiGl9aGor8zouakC/ftnF5AYm
POYLYN/7LN2EsHxssqL7vk4Uw2di57aVR84md/oeMEngkq2gcO1W0gt0xoSm
HlzRsT1sIfeIzWEKInF0qBLsDUZS8Qr1a5orotLMAAJbaAfJDfsXrfiWSGwo
8tt7Bxn1Bstj+tfcqOC28fodo9ymK4+d2L+3Un2UAiCe0Noc3Fx9LZPtgt/9
rtRYdj7J8XxsvWK5+uHwdYcxbDW/Rsj2/9rEMLsld3aQRoc9wHfRWRZwELxD
xUAY+Amq49ndeDe+hk+Ri6VWASNHc8hudOfSh4F3PXdlw3fKdyUFAd1YtwjC
S9OW9fEc3rTqXKoQDPURjJDahj6d2IRV87j3Pbm8facaDrm3eNQuY9riPpZW
MiRVS1Dm56cG3D8GME4ow5izsbj+DR9ocO1V/LrzQB498Lq33fgomEao+U/q
BT5pg8EGTNGTfcx9OmrwPFaSJCYSHdwSv1FXWGOr7kxoLTOwhwo7i+1G2InA
jY53rGzjdtJOGRj/jdcDbEHuaJD+xdsUimsksoP16OvUQw/Ga5vq0zMIgTHq
Fh5fGbeS6reUMebrBq8wQIsj9oBCypuPNRpHPBnVxTcgIuFaPJB4rW/SuoAr
IRYOsgCRfw+c4JS4gYYbIexcwqd+Lw42Isb0+KVD7QokT7IeoaFYWU4erRV1
tahZeJML8WQHSkUnl0cSNnmmtO3RLFIEgyet0/jsUUGs5UNPLtniOAlCTks0
CNyfI+/beS7QM/27iQLgX8PcQTd0rovWjg59XdM95xNCHUFdFipPTZHuu/eR
P5kUId9n86IY8PYVC2rD29fls8iEAoHYQ2xtSXY7gpAapGKNX7ADIANISY/g
EARYx4e+tz5roYv2CCsE0LH0Iy12WikCbTLmDi7kQ6QD2xu9bGP2CfubDqEk
t/f+POVtQygBgbJSLDjvMOUDkjJ/GaBe4X6SDRK3phoG/erWoCC1+72pz9h7
71djHNoG72bRCdJZp8WADMGhUl76SrGTZwj6ggCufsIG0jChYY7mr1NEiVg4
hniwhw3ebs0CZlVCJSpDWXqjh6Z8Y2aMgIfqCYbURctQMkbHLLUMNTKOVsLa
vKKuRCj7Udroe/Tsn2Zud64saz/2IpqRamop22MV9z7Cp0PM500td2E30Mav
G6OEKI+bzxFW7pLoWP5gbOXl0Pv2J3t7yt5QkUPjk2dM2E1RIvFa4g7immeJ
Kf07ltLGFQEdgIcN2efdYva2lUwwNUEuw7oUxxPFpYGhQ+fotyNKDGTop/5t
CvOiTPqgMLd6QHq6D6h+pJ2KPWiQplDCm4yaOFw6tQ/U+PeGmhTpHFSuQRsa
BELM5P3oHtQrR6KrNhdQQX9ylx3DneusgZub/x9nI+PHUNScYb3JdewE5xz6
SZOJakDDKoVL18vUHNxvAeXD2BjMMWiLc1bICtmrVbU/9scqF+nal6whQexA
u+vhbTYGcOcI3pbQj1ZsfhUQemTxvSfTZFf8s0rva4PBHIyUaRTBjII1yPJa
LNq3mn+7wuDAuFaC/lASgKD/C1uDYZcqDhnqBh+9pw+fcdBvS2HrefcI7rC7
/eiBtezqwoGY7DEofJ37XCTwmegvwANMTlKK3ASDfOx2X++zXFZ91SWMaOR/
653JjEO+gWWGsF2arpA5QGiZEUVJHqk/PZDPb8bpa8IMjQijl0+GgsctV5BC
HZ9cvjnJV+qAStk3eyKbyKNSo1U65oDMIqH+WyfQ+F+Ne1f8HqHcBdBdEFwC
0oxz3ftpCHOn/RCyaupNv4aHlaItu9o+fx/ahRFntax7iviuk7SgIpb+86FM
u0u/7rdRtaEeLMhah0fR9ZCtHbltiI2UMUEUtzm7zCxifMv1d7m1zL+WrMWf
lPcuAJ+H8g2S8qIA/uQVmRKHJO2ptt15255o92j5r0MKu5WG8vlEK0B31OY8
SgBcbuDtPkTSGCBC1mw36m4peISIKSa5y3USeViVY48kUngpI4/W/efDB/Yz
GbQ7o43K+B1hVtkRCM0RoF9M/LjbHrE4p4bDdUT1B/8+9un8r/8VQcOIMKau
EniRYRdew8ZrIe5v+7mNYJ0PTLSGLAy2pxccG569AM03CQS4MLqX53tLx50A
m+WM3J6fPc1JKCaM2gvlkql6d76qAXTksyz5c585o+qhtG8I3DYbvsQKI8Hr
VjihgvObN+D59glIf9X0C5ibG8gcGa3ZTDtg8N1cA53t2msdatHVoxCZYfqF
4x+BBAcbO+kSPotVpygCIGYY8hDYzSwo/smnoZgXK0tddW7dPV169gHi4GPe
D8YVb15Xb09xQbunxe4J1IbT53XugXksMPqS5YUOI+51XL5GC/vE59FfSsC9
XDEuuA+0xEk0hWgJYDbuRaGBQc7C0VmH4fzYOHiqeokD5TxbEsm1qh9KFy0j
+aE1hFDf2f8S8EnTgxsquL7i/HGXxpJC6kwbNiBhR27n748iYpClqNZ/+6pa
W/hDIJ4MrRPJMtpne3p0ARhFRGc2JJflawFlE0uU5yVDJ5QKlWMJO9szRqkG
6zIcQkpkHBT1NuRtJnMCKEZzVOfBdm/8YHEiTRm4jtcm+6nPF3pqoOAJ4cls
6tc7sbrGqLqA2kZb/4ugNAS9A8BFr+wfPMWyByLYfn4WCWuF6sIqd0NDDr52
wTOaieBeitCGHVB2UGDgn2rrxIhNJe3f98EQpBVJQ8g7PIC3eBNFxy75wB5o
llny3fN6KNNYUQAgHLPAL6aSWMkdA6MRjec4j0PMJeEPvSXmORFOcZz+M1E7
1nbo1/3ccafaLXDkw5Boka1EYrMFI7p0Q1EocGGO6qbKXkjlhT24zAXnG/aD
UQ2Yu19RxlrV/hSTbzKi5B98F0NCWVy5EU9ixyjuCF8xIhJboyOrqT+KzWEG
oCE7/aHZcyHlPjV1PPLQBxTK4rwbKihT1kr1qKXXj29dtJF4wWj4jCFCSBXm
CWUHo9HzQcARiOhmDKrQNxMDPDneahG7in5WnTVasZwHpL5bU060brJELNbo
eO0x4ZdTJ2exR24OYx/6yKi/uu72TQlIOpgJUHARBrrvFKgZbpm8GueqbCDf
LidcpZcsIuNvETTRl/CV+icWJ3tmzmr4CtpHtuMA1ONG61ctq98eTJjc8LwO
i7+98lqEkiy6ALWlNLzA9OjXwgGgzdZCDhtKow84nqGRpBtCWeQ6NqBiRfF4
szeCyluyKo/Ks2+hpImVkaUBviJHbl+vy7k1W8unvNTWHJJpF4a69usIX2FI
MeGzmlC4JlujaRq48v0ajRB8KNrh55DO82+ZcSz5l4ofesQFRWaD3CO3zIg5
5+R2HVYpNixE0mIFtDTiK8/UK6mpWf2y1u/RElR3w+TydIjystdfA5Rgfht8
tfiK50Gv4ZeUfxvBRMA6xWtxx2p4reuB8sX5QAgPPgBEzEndMc77YtG6PuYm
yOGSMmC5Oqgb70KsXvpmX+iXobzRT3WR+5jkIY2DOvt+zd1ebIYlVJkSheAT
MXjnW9dX+QLlyHdVuRAOHOg6LX8RWrllJlG8zsr21kAlhsHl7nFt5zQPmh6m
WTM+7Kd8fjVxwu5M+Nxp8TWpOFlr2PU+TqzZ8PgagHq/0355/faDPnDhT3Xh
z3j75gxe3pvG7wn5ZjSH3hRqK4GBN1i7c0vAPeFURbFMgwHP3fIlqN7azW2/
sh7hsfZDR1xRkEXC4DAV0l5E6GkggyjEHnLWxKjoSf7LZDSKwmk6952xcrss
GlK2S9Q/B7ZcEHVwkMpmcK+fTLI3KQK5M+jbFcOEa6iYzYmv4GEF8PLUoJQH
1BcDLG6zZ5/45ShNqBYfrjxJmPF9NE7qheqevy5QDE/67UZtIhHKYwJ+02Wr
cfOwsbXiKCof+Dvz+0lSQ7AduKBTTwc4mg0YhDscIEwuPjwbIUiUZNLfz1bu
0J5ZymyOGcNWdzqvtfmr+HwmlUiirfxUabaBxGphzOoFKDLZ52weKOLSnRNp
GLZ1ldk0yWEl5wrD5yVbRxcRQ9rvdRdWIq65rtkYT6bcqiQmCUke4wlkbPuR
Uzjcokn+/fdwfnzuASmWhYj+nnoLNasNwvVPfBer+0+FASbr7k+fQdf0fm6e
UmT7nBKxawENiZvOsCt0iZ2mX3G/WfLuWZOg9HfwtH1w+i998n/9qEhNMrN5
UlGlxuvlfHLQT94ulEgehoW75IyH+iLuHpCGhYMa2sBH0uLp34AIWknkxPF2
sBaRSpPsuBljp/q4X4Ri1bi5hyxGA6p5fqE/pEEliM5BzMHYzGcwMg5yCg5e
4WyQ1LEmvQkbCRO90GW0Toqhm6hYA3+3TF785dzfm0jYxuWtdbZDccbjTAr3
iMVGXS9tNn5sekCI3UhvCAdWuzgHK4BTleG+s4Oq/X7KKV46D0IWgnGqDsxs
wakRyxVK/cOtTAjnHhW0ZG/TQuZEpPCVyVO4edSa5A8UO1QWpB6QNUU6/Vsp
nXvvl9XHAdEtWJAlZWcrK6lHd5GBF2caNYWVkZZYUW06H+o2bwwwRSRK0c64
E18REZMTq/0hLwwJ15l+6a5eefnu+pn8QROPqaGihR0WMHH7gba1AzOG36d8
ggrVeLpeXerJf69F/+CU4AsQ6pY0MivAFNgOF/6hqx4qs4clX7oPHtWcbiRo
ZFA4ZOITuKPXE3NLm93nJyIaK2jLMqROJcmsbXrOi14elk4BpV9xhM5HL1/W
kfetlPpRCpOMupFaAUbPAgkWVjUoEfd0Ow6GelTOdwdg7VZHVwVJUVS7O1bh
yAsL4cfFJoYs3jrS2eZqQxwgag8SeGkpny/rhsllHe28CRkS0plOzZLPcOe0
ysO0Bd62wBHB7BSk83qwTcpAnxB/YBD6Ius9ToLSk7FaO0S0/FsRh1U363dj
E4RaDjstHGDHi/UM0VZhxxqP/q7Xg8lFIN/0yxTkSI1VJRpFML36NwFDr9Fa
V2MIwOQRZjegaC7XfpjqrOKImDeFSttWMTlntX6XTa8Pz9cF4qNs2bn6egqW
kdf38rQYt0BpcoT1laCyvaYB0B0Tkc2pGScwTauGnP1EAzN8HlRtr9JspS1k
6TDIvxf4Sy4uSAcFaZKjTy8oSRp02+DL9J1t93q2/S+Sy5fPt6oS+W8il5Nx
xoW98+AX0n8QsGzoC3lHMMftgtJF9p2mt6oTcjb5xqFbA+/hnNyLxOuXeqng
xzs3QiqvbFD00a+vZLmituCrVJZACqm+YcG7RB7FM/M0aXhHjMqlF/ltkLfx
R22dEOgsPMPb1DQf9OV7owdkCb7hgZTyaJEmgwoI8pul3JfUMFGAyMP/J4WZ
ufz1d2Bf1xSKn88xYwzoIJaDZoR4o8PuU6s61VODREsGHfvBvr79MrJfE1+o
yhHCi1AQXvgSN5Usv50VrTfNIk0DsZNN6hEuhGCB8rJbQwykcd1/MZiDNCsm
B0Fih3/jXICPxge4pdQi+2cpVQAPYhUyBDngfmYS389th40zrkEzVwVcvSEh
wC6sGWSmX7TeNv5w9HWOaZ93kioJsXXfwO2OkxKXywtWF4tXMzvXPpEw1vk8
9kdTLN1pb6aG50cJV4Iu6O4VR4vgVns5QMfO9aezgajIG3rP8xr0RgNO+YwN
8uy61WTH0BvT3tRE+uvYEGZFVlrE6cKie+8N9yW4sZxhxOIT8XDBobLHOtvy
uJZH4OODI0JuXSWFHTLvnhBzViXfBosduOd8MqurP3b8IqEGxJFqsjhzMkrz
pKbnpw+FETMW5nHVUhuqJwUhngb1+utBxIUhQLC5EThbM/zzajxeNCbTbIUw
5OXmjSiAy1hVnoDgCsUpihCKMnA9iVPghi9zla+QoNQtNrLIXgePcB19YkTY
B2bKkXPKycpwGhO2R8jFD5yISA9Ut5SY8WDrM6m3cmFW9LuWiggZzc3GdK/J
ch/md9n9NTUPb6gB3kVer9tIdWdcqmQIDsoVIMQ+aqF7U5EKga3vfdaBU/Vk
EGxmW0HK6wLDyPMpPITe20q2YeqRsltgsvOcPbEboEG6jm8hLiTLwGTLg/Vg
oxCCdnfxx3vtmLlhpzZNawoIU3r9skbaF9aqYfEWlzbBbIv++hZY98lC4BAc
SLlbuGQZOGu8aTAa7aaIJfA2K0TPYyDajEC9Bb8j7tZzvnjeGlZFpteUzskv
J2e4bKqw3o3T7rhoqgp2u7+G5G4U2qDkRwOsijSvfVKc07WfNx2rZHJx7a8s
g26cPT3koq4ABpyS2MxtPpOXY+qcb0fHMGgsC5cfdEU4MbOIf5HMhSDr0jfG
CMWNMLQNk/ylnWVM9JiYkDrWIHNz8qwDx0Dcf8mhivZRhIxze44ZyzzRZ0TK
RGT/v78O/UyuHjdoibHw4W4StaxLY32igtasO4utr+XE1eqInIk/fl0As/CJ
+BWmdp3ul13ceTJslVxeD1sHCuT4ZflaUejos5XPPxGvhs4ocMrIOgQs5j5H
1OwcLrrUUIRgMsd+8vIME5f6gXdCWz450xEAfHoOeLGWkXv1qbQpoXezDPPM
yKXslx1r/1FvcNTXqn9NMpcqwlwsUWAO2fdA5/LdxfT2aIJZ/wWWj/dDAdqs
ye2pUMtdOZBqc8fR/hUe2SEyv80FUGiCAXl/1udtIqlYPGGCTGsKg52/trxc
2LY59uuwwSJhqoD561r6P1UyUTOYsOeDPBejsPnc9bZeATAhyzCvcQKeFK1+
LjNCznnRHfJGGIPIXbeXEWgcohNgivdBqFW4RKzoxNBOrxosabqjrDcnM5qq
V8EBBmo6sVvYMvITFX5C589/T7DBRDpKVJg1GXFwcf6YAoWMN1oYqGTupolG
Z2EgpqCX0rFAXS3YE+iSMSleDU/P+HH0xT3cjwBwaMW/HkqVBRu7H3ZPYGWs
iEUe5Vw7K68xr3/R/zEx7gIAFGdspyaGurmUtGNInwhYtqFWTVi/Et5oykvN
yoqWHcuFhu5hlUfQ4ia1m9zltqIA/U3g1Q3wz+Qed/IlDbWEWARsIJvubrQj
+hwT0KbOiYi4qigrEanygad59LLpiVRMsAji+jh5m6F3pdmMVfTi8B4Ah/qo
rvH8ASRalR0Ee3R0g6W4prAro+e1dyYi5jBOd3Yi8yOPZpnLJbl/fFwK68eO
6NJFEtmb/8zVI6erCqTF5GbvW1Q0TpuMSQJ6fPQsM+XNs578weIfKqfk4dow
UbabjPai9HlE44FOuWdFb3PkIVCL8m39mvrXepPm/laZTn/q2l3JHaI5FzzX
vYkqqL+Jo3G30mLq86e4PL3kPXJwzj4BhoJrq9P6BnElHSIlKoy7dleGi8Lu
1joxC6d0JA1QzyovmVxDPZfolf5UqYP35oRTQV8s3EnQ582OP3sHx/A4c5QY
tQL/nHwd5VIom2FZ+WEdJqD1go3QORAEqaVQTBM7EoXORbD4KkebguxwQO3n
Aw4LOGCcuf5QOcBrmsPBMejdYF8yb0BPR86bG4QcKX5Z62g3luD1DgcBcT2a
TiWVC7/Em2bvIVCbfu8+A2CXUJFFUbrRTkQ2PQtIHK/TTgNhiFi7qx5SNsjU
/nmgnq2UcnuJEM11VSZ6NWV8dv/TR1YegrUDALD0P1kUOtlnJJN2IGP5Sb0A
JkXoaQCE0cUOTnkUlFkCk1rJ+n8LVOsZZQktBeAyxiKxFjrdUZr3aG44YDjy
37C0t6wr0FdvxAXZ33Pu8mnm3hfFhlKplCfyFePlZCiRiE6O5skBOWDD08XA
YGQ+JccAW/jUiaxHYL2sJ0Z2gXgw758lyP9e3O3fe+61jbWqSBZm0Oa+XZWK
/2Z1PyGgYyBG3ketrY7Wb1WAMsD7V+EIV4D12BX9PNX1jkkJbWc1gcXtmHg6
mdcLeYSR/yHWgzCBusxXC1cQ5F65mZwAXRBNIwy60iD1tTG2kLf+FQ2szwU1
FuQkKMPZGWOGDajrGWMMpWBgjTOV3lc+AFt6+adExywoqBitKjGnHeFRTdS+
6SwwlGRiQ2m/DpjNsZMfXip9A859c7qBeSeKWklunt19YsnGK7M/uCfNQCEs
JPw4QJ7Xe8l2tn1l6i8UJquYSpQGLdgNXhnGE8DhGzHrnxWdiu6Ua7ioEIUI
MzeOmBxf+7t+9Q/0K+re2ZTvA0D/NgwN+W8AGWQxUF3dfCbM2md9F6hCpG3A
b0Va3AfJeLVuQHO41wk1DxdRHz0jXzo4it36NT1rIRZbFpcn2WnK8p42120C
dbI3/Bl/yK8ITxHvxZQS0NTJv7YUUkEutCjTT/1JR214FJAV0yUMizn6SdKZ
DQ2hzNP/NdRJAiXGM+ysoKzWl3CU8TaGDa0RHxTg8ggoWp/FrdRR4wMGJjQ2
qD2X/vW9EAn2XRIMNHDNZt7xcVavUTdqTD6tQOLoAoi1SEenJWx9tKUuqTB1
8o4dNfs35/Ih19FB8qNUpQE9mWvlm0E2mMWZtdcNaweaLhKnRr/e/7td8AhR
BKlPFYdTpz5RtqfoqxS45SGtiOhJBbecYXTJxeLSKRqIWO2clNaIORL2r2Jx
Kxl2qj+z4UXWQoiTS8geqIDd48bEWzw07W/eoIv6aTlpLUpjDDIp3jgjWsYJ
d4JuQQK57jjFPuaV+8qINjBn7gK5SFBN82sep4PHqx1C8srZHMy9STXwPld1
J5pSCy+4ucf0ocRls2x2Ut7l7bJzqmRnj2SHvXBttB2nM+CRKHJdUMby6miL
fQteh+RY6ZRqJed21BV+eAB4UyW000vqr5JXoasYVb8ajVzHba5+Oqm79P6V
yxl9r6QaCD1Zwfk7P6ArhlvQ+P4TBD3+uXWRsdRGHCqSr98Suq3La7/j/ufL
6UJWckhagvcTBbktS76G1LDPrTNZG9ZjzVyusUmGdnCbeN8sCowVHpwobypN
tZBEWatIBwk3rD/nY9bYmeHvfzXtEy0+DbXUSCcNcxBKKxSgnQkDFyhIY2LS
oTWK+QS9ezEPh/cVSgPId6sTTZ7lbKCshdWgLQyGIHAT1lpq8/KpWP2AvLTS
RiYXu7BgJcXYjaiUwCQv29iHabyOCTM6UqL6ieP9ufNO0v4UctaS3caf5qUa
u0nESKAiHDmqHzqQ9wqePqGscv5/8z0hRT1dknOwgBOtLCEKTFQGNStV5G1M
Sgjs36iNinZetDhyjw5WoqmCfltzdDxMy2ix7lxZ8ZGoU11fqTo92oTn5siB
pdn6+BLAv6P/xF7zkE/cSDDpOSH9/7sgEKHo4h8MywZbnF3q0+A5y+/3/OMo
w7EUAxkFWnMLbMgundx4CSFVE1JT4BpVStRjbtJrpXjR6UQLSRoUsmRPZ6c3
i9vsUpQqSFwnKF3yo7JTT3l/o2/U+b+McfZYOZiKVRBooGsyCGbivOO6tKL1
w37a1kaM5Dxc4RRFKq91geNUGt8mdIMmHf+ItVcGKpgsOsXSU5we1PfzbL/C
2I+JVcQlaGoXoRzgZZvXMzb5Z7tnOjXLxzMIz+lmBcSUlYL0iiNT0ilAgqxd
13gFNPJHZ7RG+2c1TwIgpoWwUoA+AqLYg0k7mHN00+xmE9tY5EIv0TL/YXUP
4LxSG0Q6TpB6+LPMv8CZLUhOtA0NZaBAIOGK3eSV45Zfem9RMysmD7fMYt8w
haX29c6gKJC3TsPr/h2Br6BjvUNiqaAHZAu8mQ29wPY8pHoAep5XJUe1/D3B
ye8HraKpDSmGrNuHikppJctKFBqzVqMWPsQ0kqqDJgmCts8PqvudfhSq97yu
KDtBK3vCQkOsbUGnJHX9LV7xslepHwxZwNsuAL62JVphLglaIBKv72aOh5++
SodQb0+I9SxktYSDvU0oRYoLCLwSQN9SnIPCmnA4eXdCv0ud3DQI4oIbM0XD
se8/4nxnK0oHPJeG7LAEEULCAMn/jy6Vv40lK2WrzGvbTFYUY42a/iYqVqep
6n9G7hqRtgKb1iheW7FrN5rEGoaeudJczyXnc5jrhqiLs44AMJ7QQSO0nLuT
nJeK0azmMA2OdXdlD4enVHtF2+YykoNDD14DT1Duy7l1143DZqmx2YX19iyZ
dh04bGT13e/e8tU5d0EQmo2a0BqHTAD6EA5szGojIEgW65eIn1PVBYRSokQQ
Ut8TV3Vfw7FcXUB3vVn5WCxJwtJzVzwOZv2lez2hGf3dnEN0vrzy31/svZKn
3wMnz4JhiSIIsXGkkWGtbQdaZRauot48Q6cLHHUXCi2cRmG054MpZOlUJQph
WJAjPsUINAz6JzfJ8fQRKTGxbY7BCumz3kmNz6+5DMcFIge5j7Fp5E1xyYqN
Ausw5Q/l+gVBibZN/feLSDSRGnDvgO+CAMe/VwCU48jCNFzkamezLItWt2NJ
a5cTzDkeDdGRIXZk4zH9QzOc4iZxvRK44YISY1/ZygRY0euvQMfn1kNIfEfl
BcAudEpdJaobBX2FwU/qj9pAgEd6xsK9F4TJhUiScKCT/VWo5S2ar47Xu4gF
2mXM/DURMduBf9pSmtBAhzffNUWXpaiURVCOKL8J7uUgmHgDCQ6BW1usRoRb
C5pCXgL+vxSny+HkA8h2Nnw60EFUwDetZuYxPh+H7Zz/+7z/mVyokt401r8w
ONi1gy0pHGt0X5T3PlFRIN26HCaXn1bqQltKuSfnN0LE26z7eVx+DQvnBWzh
wxrT25a1cF3oTPmLZn77IFEtjDtTeyZ3UDS6o6onaqBe4derxFry2MtOmPqB
gvqxzaEo47oiBU0JnqT+ByglaHMXVYzZH/CzRlLCF5o2O6H4gCpDop6Gq+JN
zHBu9h6Zoyda+U3y+aU06cHuHjLHHaZa1qOFw/UhR5BHX0BHsshC1dJvBMS+
1KYcJUYs73w8bJmF0ycF0MSzBo7uw/Wk1QToU4wy7m61zgSIK9oSk85uxSlg
Jx3HcpiXtCjLWuuyOrAloopX6tDIN0TWqiWV/DmSFV2DQgoYF/zohs8pVCBa
T6nns5WcXhAPSfANwWLxVzRzGthGud7bOO9roVK6xTvYLEaFU60UMH2Rcqe7
o+exAWLibSYDmrYdve69sNoQFN28/2jHP9Unwvzjs5tap2RWw7x+s0OrxIel
KPDH5E0mWe698zd5y/lKHq3IOiawbC35Lyw5KFHTG+dnDXHYKoZ47IQTqdWk
6Gj/ek5tV2yTiGIOj8IEhI3cEnDAewbfKszhbishdgDXx5rKDTRln5HYpLrN
ao5paGKLxyTQJRiD+oYSE2cqbNBzaMEISEQKPmiF4vLE0QWoBBMMiapTZ9/E
km6bQsk2hfncn6YyPpNPxjtSflF8+0IIsUnu0qxFTVu/JirjroDpJXaDx38A
D74q0hzXtfMlvzl3fI9KyxeaTXlkaG8xpHntMbtgIupqVkjv4a1l2lRY9+un
HZayIQ4bP1pwpPGJQ3JsmTkNkux3zmy+oLChc93SlOF6HAQqbB5+kfjgPK9O
ZabVVYof/KlOQkO9hGW9CBRMeBvbnuQZiHtgaBB79cSuTHW82YSl+yjxsj56
THBYsM+T1bk0AsKMtwPQ5YeUYrJS+PWASz+mnsfZRyRYQ12SyensYRzLdWPX
Y9pT0w/BXSVQ1jhD0Qr00mow7DisLIjiZkyE4dvi06tyiSKkLZkx/Q0hGpFc
7JJtzvfcl1vq4oAKt/UhuQv0N5bqbeKPUKqxV2N51wEJ5pzK9rV7UlZJFabs
Ih7uw2750d2JJnZVQjdbankMsrU50ypNZAGZkRzikAE4XLegSNa1xjp2GhvQ
3P0p5nDYbQ95VQ2RD6ic+TrZNCWJPaP7SEN180fpDYlihNozUsL1EKPBEjOr
jfCuqsY5MvOi4xYnwkCKiCBuEkOsHcWNHbqIORd6FkQ8I6LeVOHMN8Joq/R0
Blmv6JnmX/MF6UzGlZaHGGjV0b5F5nS3KikOKjhAhG+iZ31QpU9UFlYfP85n
tIZB4/mIT9SmoBM4lmlR6CMWFrHi510ha5F/kAPcqpu3XyC3Wg72iO19Kzqb
HakXg5kEBu7NpzEQ4fAa5HPhMK/NfRl2h4cqAXBcdUKz2MYu3vpqxwBd0iLn
d/A29d+3FKS93QS4khgu7GmCSJg2La81hNjn3MuHs+ffZNTah9yQlb5Rio3j
Ext+WlTIZ0bwJmzEOf76w5WaKh2Dl04Q6RLbNCwo6JWIh824Zz7t7tBNzULH
h5VId6eAzVKkn3CifwlQGgfn7H7d7r1lW0J42D2L/ta6Aj9ZZh9vKfjgxZTd
sHXNX63jHa4E0Z6eid5ajfSxiDeOyfDP0Qgz/a1C1Ok6V2GUcOrYKJj4jN9/
W9yX/KpIDzBeNB1zxk/nghtgpur8buHDpssnuc0AmnKORG+q5REd6lIgkSSX
C+SAmohYS318cBbl1s/nMs805dsNFdIUhAa3tOxY1CxOXBzht7RJ94KrpVlO
zJneaE6IMjJrRxnySOn9kcGtllCagtiP0O5U22tNUoUqeDHbsg1DBH+1LMMH
F5i8dlKwTxVNeg2oqMZCDNHJXLFTU1v7tXyQVKpTnOnz3fe+JZmsNR1Y2QoH
TOo1e5dHyeOLTwshKRnm7SEmgt3sPxhXV2rufBfPy+oPNbgQGsWDrQRIgxAf
T6OxUdSiLwdQ6f3fXQMx0xMbap1/sBltPu3F9vAwZn0kZ4dsi+aMneCqi4OD
qs/To1l/PMN3ajZUOn6Q7gTkO1ZZGSdZfFmRkbJ497xwn7nRpzlIafVNP6K7
P3N1g5gGZ7o5nZ2fW/KCHNsCJ2AwNXm08XLiWYzfwytU1+Q7llO8Mi9Raxqq
/ANaBjTFlZ41KHzTyp+Ef7BJJhb+tQake93d1gwnMiA6W7rGDP4Y4iqxU4j3
UA+CIzwtOtsVF6a2m1h1Kdh2AMCoMIkfEXE9xxThK+xCrmyydarxTB41ors3
2ydi1ljI5efelW4tL1V5BCy6P2uBHCbZraZ64aG02mrGVsqYfpyUfz1qKGs6
MQlza9v1ex67zLihUw4wWZ4y/8NCH22pSjhdbmb8bjzTzB79owZ9v3ifB9Xd
rG+UKU/77JDCjd25nwmv4EqPTSoWJg7u2EmWysMyeThBrGFCU3n+INxpcBuX
BsQ5PS6jVAs0t5HC4xtWh4cAqV3ZHknYG3nWOgmryPeJIkUmc0O/sRZZOW8n
iKnPY3mUXkggDTfbdrIbcXp2MGVxeXYJ65BaOM9lz9IMR89ADIPx5WWNDLsE
fc565TpcmHtonbDsWDhtLG0zwtnulOqiqdR1Fok6j6LDt2KZzthE2ERC6twE
8WGaV2awcl7al4M2xQEKdPnAF+qjXC6n7NXnIhdnYOxofMlcWEWUVFQ25QKM
bI2wAqqIDzhMFgJYGW4kGGnayS69b0KzlTqHqdnCDs9/FqpMMGIHyrUNucOQ
s7rbGm+jna+/pCW2KXMvZqAwHl6MT7DH9gtSILXG2mA5ah5QJHMrux1aXpsw
phs67RgnP6u1iLI0+K/r7t1YwErzYgrTv/aD2x6NutF8OxSSvsjQ1pKCHvrv
+tPGfRut92zTMitzZAaIKhY5vEXZEVcPokmIHXct2WGaA7r1LtsbFPWDcHcT
nLGbP2TnmM0OxO1MD50400BNEal0UW/NFgOyKLkfF2Ldupa3beP0lYWwQtgU
oZCmVKd4SCrrdBvJHZr8BW35rta9np3zM7odD3Rxyb5SLFlp9nkzmWe69aOW
zAAhyAm6tlbNgQbW6ahlzLQoLw6/L329OTlHhn1rBL3nRFDJwbUMYj7ug9Xi
Ol/Sh66u9g3YRpT+8rkbd4dIh7jAfEUi+mlPDNW1aBHtijI0xb7EC+BvhaWC
Fqg2XLZVqLZCxR7iQIEnLesbaf943wi1q3JRWaJFMAssKRGgKwp9zUfOEzr0
AjW5vTrq5+lifodPU0Q79QbODLgul2VLTP4bxo/zSDqbRfpqsF3m9DG/7LVA
7ECldrKOThc1G1Kqe+N6Vjmf7YNpmQSkiIUAXEbaCJH7LqUKxCKPUvfZSZUJ
Sh50jk7UgX83GPaVHBvScGVyGh8nNwJaUmP4ZSrDOWvNya6Cusxa/cFqmivP
r955TKN4Qa6rzuC2q94jqHeteVBY/NXaIhBU8S9rsRo5db1bpm46ipx3cmX+
Rr0Wmwga+qF1WBA5Qmw4gZuz+Bdr/bY/L0KJrgN29ox0AWUrnpxP7Jh8x5Uf
+G/+wdz8nBP9tjftJkhBRL0wQoIUqPU/gnsUq2yfSeN3gxjfWbOUjypMS/JZ
irpwhpxBNRHklZI2+GCdHZl1cDs6zHHq3Nt+P6J2BAl6MJ7cUmFop/7HShKD
35uxIEwr69PUl5wMYRV8ih52xi2ySA5XW2mufC5p+AcPaMEC1cQ9PDDdCaQa
Hrojysu/2gck0l5eGQil8zi7ZpjuKWnw+bP4wqCXqzzusjnpmA9uv61MLZDY
EMAEoNcvoemkdsEybSBirA+MokE1vmvz9QivI/bs1JsxTyphttt9LHs+0JZm
DVPynRSPXFmIcEZ6FFzHArZi8Qp6wrhlx6iTNhNeHP+FWB9VKWiUWPgQqNzK
p+/ERc4Abw4X+vjT/Cleo4dS5Yi/rubJAe5VIIu1a1o5DhzxKvxjxSgjXZxQ
iaFoqRCQJVVR7EgjkQT8AsD6vtAGK5VexTqbArTJkZd1ZWK7IJNeQTrGEzQA
KYC/IAezmaqXtLP06WH4JmT2R5y2sC80H0Bk0WSvcErbyoiyMeK1FH+52x41
hAGRVRGoHB+QkoQl1ypbeX12wxBd7/ZhGkmTRcIncpk/vTIu6xyJQ4qnbQsE
+eueMvqi4wJ6dfMaODk5Oy9NvMODN0tg6Mp+grpk/8A6uny48zdvn8Crdzux
FaR6iSM55Z2pHE7bFTBI6hjXppTV7xd9hGvYIJR2y1F4wKhJ6XlVPD/v2Bcv
iMhf+gOBCZ9gCbz7Qn8ejZES8IYiszA//Ak9xjYpTZfk54YqYMCz6kYHRDyS
i1FIJQTm3bsnoHvcalllN8l7/i6hZ/dWrBYrs2eYIzcKvBRH7GdCvC+g1FNr
78QTqYKUIYvla5iLS5Fk+xbE2vzm8LuzuAbHSSibpKkqr84Z6DVpboWp/skF
FQajvgbhPD5z1WQOXca2FCNGq7kXVuSsj3OCKJ+XYiASsiJBUCLPl6PoBaAh
5oHI0rgEwgamU49xiS61+lSo+NRilUX/deI0r38/FIHBmV5BbLdYyW4yEmdt
o3NPiXVen+nqQTzVRrBjYMCjp0+GH7+p5GPshXO+ppHzuvT1ihYsRLxxPt/B
iVB8mVs7Z06G3tkJfL8OJrJfcEGR6chfue+9/an1wfuc0th7PbbA/UlPCRvi
DPrC56Kv4538GqzaAx9BvwkDErz9/VDJRV2220dkStzh+p0IiUpas3KpAoaA
Dtj4yv40YhJQKTp3caNN9182+fi0on1XgqM7zo1VkDkO0Uf2/RZzM+D0/O/O
fhyasBZtCKklLsLnofGOoQ/h1nfdAuPqf472srHpkgxmmpRA0CoGQf+eQMqL
EbNg5XJaii+Vzt0tRV0rKAaYiRqeJI2ZeltwlfWay0apK13HgoidfnxkI9Y2
Cgjh7AkyHPTV8EQsZrk1Hug3dsQZu/rVSRCauL9mXTtEsIHI32/dJcrhmofF
zBqvFjeBERmcJlaHOw0cC0DjCZRpf4XVsapHrmvQv1P0S6dMVP3s8oAnvaVW
kTqdqUWayk6pJta3CAEBgT1TZgsJdnWbPKP+H9k8f4XrEciwBuvSbfxVLCyT
XyeczJeiLFkwZNTTGRbLMyHginVNztJ+1KS0mItjuJMP6rES3cI383oC5Mln
4oixdHKxGh3MO4nAD2kgh+UfIkKMww72flPtxZ23pfEE9qtUNVjk9qSTc5Q7
oqKynTxcvDyW+Hy3grhH152bJZIOwyMvJIRBKDNLAtWioZqHyo7dEn+gdXQr
2n3LPoxqWBpTDt8BpLzlKJXEeGpHe33XfevOVAZ42ueQ8iMpJ9m8WiYmkEfX
q/jZAhvYDkB6zuxoNECJ3EriSFBHTzcdwCK9U9J++WiESgRDfL39iQoxx0Hv
EkO8i9+I6bam0wtA/LrkzvK4ytrp59tZsO8RMBGKfbhbAAjCc0uN3u67Pa7e
0Vyw2ReYudZXd3KBQtLBbX3Qm7zxSFZ6izoxZYFXH6TA9V9wd03SSr95FT/L
N6EvZ6xymavylnGj/Ypyx4kArwgahJQdpZH+0NSsVafgNYP6eoU/yJa9S6cl
S3V1PqpgzUu4hvp99nP6BJ1YM1KQI8wu0mSy2ZiFpJbh3F0wNeG0TLcm3QNP
K+vtcRoIXgsyxvM0nAtHeLRBYyzRw2ljByljzFjfQteKb3AnB+wTnGLhvm5L
QQ/R+6zdRMpa9qKHr2cPgDmefHZznm36zmzwGlH8IgJsw6kbnBBub/wIxd9l
m7F5NycB6cjykU3l8OohU+mcI7qE0tzBZ0+Aetqhq+YyOYmd5jATZVU4qSD/
mtgX8uh4wslJi29IUkABTV5LuvZX36MrhowPW47hJqtfkgfIl5oWHfoMxLK5
ld0pKsF15mJ/GmDOIUHA6qo4djwVSBBk0p7fXCrGszhgvvUGWnOW5/BWr2vE
38AoZFalTSLMbCpbsF/w90SChnX0SBgHOj8/51JvgZCJGYwMavIyVzRMZyOF
X0WiYi6PbrKUjBf94A4sK80gdU5IwkHe5Ol+vtXRE/Wlyd38pLJ8/N6kKIKE
yLJdJMybxwQeB6j44G7TKGzyApeaHq7qqrm8eMOMRZJRLgLCLE+wRTKj0cuv
CEztZOemG+w3d7H06NtcLhSJzgAsP5N3S1CdqprXD6Qqi66NkT573ZxzDX00
/dGFJv8tH0kobYri/PMnaSwMbr9Gc0jUpbynWfWwiJxj1CQUKqlOyoix59TU
ABXspsJAtc2glAsmRmypCp85v3voTZ9RCr2PLADWFMkhmK2ONafVaaBz+7uT
QVC5Lk5Xiw2g8yIt2EK+gW+uytZx7W3LnvbZtSxgXCYrN7SeEUi9BbVCVzsX
fy+L5GouKShjRwPGMjh8Wu+2HmkhtpEVIFDiD2nWuXYGBVwknX35CXXSKqDg
i5ykE6SxZpWOavk1b6ADrxsuBVaiL7Gsnyd9JuGVCsHkmu478ZSlzE+buUrI
hw9BJ4SpTi5TI+nYcxh67S4iSfXNnRm4aIzyrlXlFzFO79bbnVuVF299kMTk
6jK91sIYli9TdDVAJ5WPLm9zqOULYvQ6L8Yd+Cf2TBqVKd0hookMeJRbljVq
r2WYNzO17abSHLm9YknrBlhv1dGWH6jGFbc7TCarah4jxMCo3vuLZW+N2nOJ
msBWeGcmg9bDT09wu1lvPACaraNQqJHg1CMKG4HNJS3tvLwjbMzjvemcR2n9
VK1nBjnABsCi1AzIvttyTAUiJtNLeAimscA1GXZmc25JfAG3+wdtZ7Zm5bs6
Hn/1kQ4r42JgZGrbiRowjhAByzAoXICr3rIPApTlpqJ4654HGXFHfNVoCX2W
6avedENFAQ678QiAcxGdJn2YJM9EeWKbR/3TIwlQFOADwJoPT7QbOJpqJy4h
xhXigngu5QD/RABp0ZFp8SImxhQh4kGKI2xyVkSndhlWuirMp0To8lDCojng
VsSRHGImbwDJIs+GUhbqiTHNmZYTi2mTMWmWcJYDm7FDJXwZbxZuclNoN482
Nc5zleSP+9RxSJSLw9PFQw0MGWcbzPGm0/eyJaaN78ZWco2S5IO4H48C8K41
1/dOO4LU9+xKKiIO4dk6DndqfUW1yTNwzdJslEs8QCfdWqA7kuyheCLiY+El
d5n4RCJS+oPlZGoMEH5Jvwyk/mIoCDBnIXE8iAySa9zgceq50N/4x7+lWTlX
xvdVAwSiHDRvbY+S4OjGVQ3xlCutDfWGf82JQV6j/SGvRpoiYOwrIZyYmIkr
4OfXq7eqOshFMpZoaKutB/PpmamYho5i1MJ2ShT9eQmgx3UtEYeNK5b4Tips
0rGiyye41lPkmytAD88TplRkEXEEib0HdlgGgwngCj3wZ1S1HpMd3Dftw4Us
32/GmNnYq6yGAPTUD/kprv3xBBhUSf6WdcFrcAaGA8IDbzwpowN34rLJgNxx
0PDB+c0h+RTQjR/edJ8jFyLnmaeT+pC5sDLZnFF8IeqlxelRhHzLzwlIHqNG
Gng1amWxhSaDOjrSQVTpRhnUpJgAoUTXPH1OEcY25q45N1uM9ZX3cM7Rce5T
Iq+Ju+/Vie7JleJzprFBsi4PewDo1iIEjm1X1Jcps0YHcMY5MP5NZkhV+YMY
GvF1lBiFQMZL5gXFT70PXancWpk9GKm6FCWLDvDwNLktELvyaXQIIyEh3W7K
WiVhSGnRHPrGM7f40F1vb4Smp5+0b+0s9JKI05+Mc2NCKCO/Z/Yl/ZOy9wMN
flWOgU3/mghLwh2oVXBj4LPaMLEqiBF3a4gzRQtA4l0cv/B6gtneVe/4dSOo
ygMYcKRUBSay1AOufxJAsHrNQR9HL/HkdIP0xCA2F9jxY8G0kd7Yaf06DQD2
5DgD9moRe8gZHFcCIl+w4jLNdZEkbMQ/JNvoHNYPuo4Bt3c95mLfYaqnHmsL
29yy19YthZkRFduiXG1OdaEtXEEsxV/9HR46ItRG1/qBGyv9lFrELRp9rYXR
USE17dGisVUQq3xNVZckaXJuxPLJk2uX5OfM1Q+bULoc5GiInmSTj6v9S7QU
xPt4rNcNRJAAoYqJl9tRX0E7azA72ED4b/kuj3X/9AYu62uydmTfyrNiKN2D
Qy0aSoMP0lE6RdptiXwH1Ft7OgZ7Weij9JkTwM7fgtqkqkwek2xdjsob1zjV
flPwZxq4x/NpDGF+9sVAMvBXzmlGFyQPWdo4kVybqQHFxi83r4HfV1V1pzoN
YKBHFFmmp4qMhUBqn16HBauE8jIJ2qViPuMc3rpp28aeGFyupMh80k+yU/DE
whQ80RPdK0w2nTtzTB/a6XIGD8iXYGkDKe96Tsr3SVO6IbjqhfT1wIzlQXxT
UPANs6/iMtfsXx9nFYx77TZswKbZD9OLXPW+oqB0SwPGl3pr4h6CdV9zAZTv
S27ibwrsaBTWYJ/GA3Y5ZQ73JnKPnexB/Gkp1dpwTJrQ/McVQBdixnWpzqVx
cFN43EkBW2SP4b/Al9OqWgWfDNizMnRxMN//+HEPC6jmsWFWFLSdnAG1r4Rn
YSkAd7EkelumaBSd+PsLF3jafPa2yXe0RjjzrHZTgtMqOVkGeOikTh0M6Dho
bsz2aa/HQhJjIBAZ/btdU0Dj0oECbwi1fIf/yaWzSCZp7wL8kPog+iZ6UdXl
ARl8MKsc4eWbps+thH8U26Dv1d6oMJUNHfkbTyc0jfzS/KbeZcQHj7QHXU8E
zn1KRlApll9EJXq5qkAo+3T+axZBx9/9t75Q18EVb1orrO8Df1kF+/8MaYtM
/QrJ3uPiVHgiGaGtBvncwRS8/P0Hti/mxCpJdvwif9KPppBvCb2dKE6i5rMW
SuniCsvChwn/v3nWtfdoYQhHnfepEUOeYCsoSlvqD4puFHO7hB/UzFgXjj4f
8+IVE/YHcL9KgBidiQztgnYca/JzcrqE4kyd0JMfI40CbLSvCIKHyq2PtJ76
Nu/XsQl76AYNE/6ypp1qRwBwkFsocJdxuRZxrh/NLtAnn12HdR7bQXs8LUTL
lPxprN1ixDuaLhkNqQRfm8WpvYDRXmuZWjxFHs8q64JJu0hRfPy9ucpUp1fR
UEkpyRijyNEWBZBJq3DbUDMwYy+9J0xWp2dYEUgHp+TQWzdTow4phA4stkIa
ymky6NqsC4EZ7NJy3e++/aVhU3Ekt9JTsi4xsjr1n9E/+KJw90vZaDbbJo5T
qTzG6RkVjbopGFH2f94Au87aZ34DN8IA9UqBICiyLhrH/uJ7dNhDiZzUwj6j
9P03samAj3uMpSQBpge2559rNPoX3NdvaUbZb3F/dZrmlzmPvP/k/LGymi0q
hShPDqOqX/mGwUXxiC0TS2I/KiyO9U7KDbejRCfZyAB+3zpHHmFk1ypPIGLd
P1yIswQyC23Nd8k+JTAUNG26tAYHqFeqjlPNWRUJqihuOBQ1pF4OuGe0YO4d
oIzrXHpdIfVhF2eBax54u+6t3OqUB6Y5ofVT6wl8sD74qyoF8Y9tY3Gitk7U
NC45OhBcdPhcN4uFi7u+vmm825JQG22coYGQ8qwjzgTc3IT+Dyy2+pFWueeX
yfeB+4mXDHc1frOWS7QQv85Eb5keaPxqQ5nkIzpiESCib1B8kNsARyrTSpnf
/6QGRBW+g5wgOZdK5Ch06ZNMZ7ihdi+rCZh4/SWJHP0h4iaJgfshDt0EXxDk
h/Wq2acCNi6RkICsZj+7/6SaSnWDNyfa14bQDFNykNKBYkyLKmyE4yjx4r/j
s6y6CtCFM/+V00bvLD1STXyX0ph6rMYCOx9vvnWpZskrrVw32uOgwTSHHqoS
9CI1Vqt7ewCyS6t1nwtevJ16rYEO2puXUTiCASjlCk9a/NXmzZBqATzMgC4w
gw1tygnCVB2z+tgFs66osoc7ru0iIRxduvaKUJKuIB2nAnmWUTXhT2b16CVf
9YZX2lTzUNlyC5UDEa3hxQ42IcSBg8Yc0MXmFZ+KWEvL/6Zn/UkTmL0u2VAw
tamMj3kOdLPY/UwCbDGAyxyYDbn6MAIO5aY9+Yk1ZpmjH4a9Ytw2VLAwbKTS
ZvX0byJzOKhmeSsqiiP/Qfn7vTRNfdsK/KkbH+rTQKLS2x8PN7KjdgtLUfNs
HCVTRKV96NwplLTI1bjoJXauxvwBGQ4dz7mpVKn/wxI1f02Xsr8PdQfOxVpu
hla9hs+UOXMbjXvaHz5d227vMPTM4ZCzctWSJa27y3WmKmxfBk95OODpmRvK
qFFgo9ZCwXaay1Y2xe3rDHIOV5e6KVa/WIJ/4F9t3Ft59hWayfJdkmXfpHHi
IotFZBMJ+ko4oT56aWGAIki/LezAwZ2SVvfel/PA8NlAYfv2JLadaXw8IzIh
EmOD5SFsM6LliMWCQsWFgxJMDobP0joIsIYjSU+ECrDkcHAF7DMVqG/X+art
Jcsg4aEJAoqsLjjCWjbni6dmYsabUQOfxNNRCz/GT0VV59xh7FY/2n4x9XKE
SciF05lk9ccpfjWshlHbVq6gkesvlI2CUmSkGwy605m5yR0MCjQGZ/nGx+QH
PiijzKQXbcVr6tlMgWNeJt0y/D0lN+nBWavL5kVqjKh/wDkrlQwX3D02tz/w
KMynAAqzLgvjSIU2KWtw7n7Ti6aU61ONxs/fOe9OTl4Q2sTiC+OLHTC1whKl
wtUbqnDYsK5jUTYaq71swKP6zdNmAzeqIlU2t2yekzskaAp3jpYfGfdFH/qu
2iFTAI0q8ieBTW5uhYLH57MjfXxD9BLL/oGihVj/YRDU/gcdJCSmlLk2YHOg
8h+94OCh7wwrmfHc9ktkpsQAAlhg7RieQmhDNRLsDBxUzs9+ksVue9Qc8C19
6uggn+LeM9TD2BOjmhpH/6/LVph8cb4yY6qsZJLwH/E8HJ0HKCP1/D/4mYHA
zakt2Q+b2S4NTKM72/5sLVXJiIZ8xmF7ME9rYJJ+tDt0b5h/FJ6IyRZ7UCpv
PIPKpCJTF29t78We/8SVmzoJtU2BPz8UlkRVHsXBv36wMg5DoFsTz7Q2koy+
D5KxbBUhg12uqIbe3uPV9ESjGmGQqZULA2RWH4K66Zedv2D33nE+miXnsias
SzHZwi/yK+isfYFNKwC8SQvKNZwlUnadjStUZ+VoZfsaNXYAiY+fPGm306jk
nuL0t+dGeS0+CwobWAtNvKaMP8UxZCVpHDFylGKREVfQ/NDiLXrsAHhuYh8l
f0oaDL5CPzRirl1pDGzUE0YDQnBkGQyV5Tl67H4nYz8AuNct89GFugPiqs0o
JW+e9TEV84KWpsLHzXHk18NmT4HQ3Dg+/H3Xry2xHjWuCJdAjjdId0Dg0nys
tq9X/zKx9qt5SyPgGeBuqpcdMu9F/r2J7OccywoYqSG3Ny4B/JxwjsSLq2jX
jP1cNmGZem2aonY0AMImYgNw8FskEXIlm7yMwo0qsuKAKDZMxZ3cRqiUZT4c
n3n6mUT4kDAsjUmDpq24GuEFdXObAHHLTdG9nmZB2TS7CBf0ApCHS657LFo4
LU6Dm30wzSIrajsHQiMR4KKcz8B9qV78NGwtFpa4atbfZjh9Dr6zXI6qC53C
hKIphuiBGnPqCd9RatQdqtuuPh8lCmLiowlUc8GsmqQQbogJ5+ieUno7AR0j
gmFZW0Qcj7gXIszHdo+Y8u03zQoquYW045ki9dXcMGqoHggH0qcfcr72fBtS
N3pwyEVP3f3Tb0qCYeUUJfmyokCZh0N+JNk16G9JDS851sdOvb4Pd4G1hpqx
1MUlpOE7pwVM7LOyEuhGlkYrtlJ7yUzIfm2EhNTepbMDkxi3+oFVr9MYAbsY
EA3UG3ECp2Zgvo7U1htXeVFNQ87wpt0bBA6QoqaWt/oCcpgGdQVU1o/5HeL2
BOfqkCUXefOO+HJWzlIXKB76Z9E6h9nLdQf3elzWWzWKZUHUGUjwokH0QTTN
W2pscW9pZjziiQIRgUHjem4Ep9ON/XJZbDC0CGDAGigJyr6w95BuzHeiDpVy
26xXEfKf0odtgh7VBpP1vLHH50siPy1cGRMbWkiKBstuCdiBMTEmSqOd7Hf/
7x08FvHNJMofebJenkyoUar6t8PoNKbyHhTuhIM1YA15AkMSwx7nPDmgM61Y
UWfpzw33YcgyIO1tsTukJfKWf1+FDZxLETm1NdV+ou9yq0BdIXn2I0Pf60Qf
DW45ro9JDJ8YaNSonNYEXUq2f/yrQqb7z7BE6xpvkLoeEbUcWIcWsFA1/wZH
M9JDmNNkUiDyaOWZpTcltGQbWdpCwJ3Dcp+5lB1ZzZZvOBkCVJiKyhaoN369
4cBK2VYV0VTxwkkhIx26JyWbw8u0B+hPUJatX8dn0lIY6bEoU0JGUIgss8lh
czhAjv8zqL/a/XLl4Gqdg5MgDnfHLFMod5/M1glPWdqpyl1sUbPawqodmf7F
ZLX96uNCuomvhIeT4X4cSzQ+nih2eqw35ArOmgK//y9g9T7HRu/6uJdWEM0t
CXytn7oxk/uH9ft0bVIRevqrKKkXLKCp8fcm1KPf+zKquJmlGacZQYPSCJ7X
i+tHGvnbRs7aBSsKNIhty3JPoERny7RLscFknlV4CU+XfMoEnsXPPKX6hUo7
Zm149GmBzREY9L2OIzdVNJu30M3002kV/pho6V8b1eC6j+Ic172ROcJYez1l
Pw1G4ovArfo+e9hu1Bz/EO0W549RrcE8IqiQZ9jQYQLEFISXeSnt1Gp2OTHP
JPCNTnEWeYUf5fkUD1yR2ITiow3CfxHn4i/qRbkPcP2JskV4APVpH+P4hiRw
gYcOaG7Fb4pZeAJJvKYuL5O+kr0FdafweIGFo/k/dNB0a7cG9b5iKCwlXQFx
+wbQOUAPzXI542ZIF/CwCDFvg/4wGavooqlWUQe7M44Ijb+BaQ8BLvEGtQIf
Mw1dHJSvwqhxouFyT/+/aFwaQlkbur1HCT5fVtdiyQx39SO7+aqVIhKW8IJM
yli0e99vshahzNiaVg4sk5srOQwR2XmdGhv4MR91ViEykDu3ye2k3ZIV0eCH
NKrlETarIScYQRnN/a/YC4PvSVjFUyibVh/8vuAERk/4iZSIbn7I6FyRDs7g
R/0XUKpV7hd++nDMWWDHfSeriUa7B/TEJ15ojY5llJk+hxfZjH3D12stc9Zk
k1H9kvp4vhS+gKxYx8hCwhghJX1viXRd4E3DhKyaqP7r8+ZYjgv5ly1uSCL8
dl/z4qrH/mh6FJL/4n9luGnLW5Og7gogScv8y3qUMZkKk5DPy+CnedilE+wH
OUEJ1W5FHSGdMpOL47fMwylDqp2xysBapMsWFx5gzNL+gyXF6f/lFP5qPbng
Tprv9zoIOgfIkoijIWZmNK0GDOvYOFJ+3060fgFUFfWrlV/H5L/fBfzFGNv0
gliHgrHb85gLwQ54pIFOx6sVkqb6/pswftJFa0cXct4l3l0ZRN44N3fcs0bl
rg6i1El6HkM6uoXQ7mQz5cz9RbLDd3u2mh5Ridc9tdWynARw0bvTJT5idkT2
tD2wjeSI5efX9waPSiRZY96fumhaIiSqd6L3fIM5a5unJM3occtUaXV1MDEi
Y38pE/XKl6Y0CuOtSEb/8aDQZhN+ubqOx/SMp3V2qyUw29hlVEXbCpf7QEni
B8if44BycgUTAzJj5C79mlkv9QRm8FoSb8O1tY05EqkNAqeJL9wUXfLsmEa0
KxaYEt5ZSOEw8/on1nxI4fZISCyTVC32LmOz/5vuUNFz5BBD1x4UOUPBVsTo
MscmTHqpQkGqw5iRWg5rF+ukxqS4IGfDonZ349hZPQvsA58TjYxXD+EfPb2x
HSz4h32DkoNCZnxdtctDuGoPNvr3YjKaG0bVzjEQtufB3tTNcsrbTKXicB3J
BuweE1bHkdUz1STIgLUXOizrSF1JsDZhH3BGnBj/f/aX8VFw0hts57jYSLdr
j+Chlrsk+YsV5xa/8MYJptB1ebhHvhvlh9h4ctBWvGH6p1dz03ptHhJxpvXq
A+YTTavZs4yYObCD5ZkphxyaNr/RwnDC79qTDM1ddrkUr4FAMjDKHqIRCs6A
xwljANgsohp4OcDSyLwsbxo0HQLD/yqqaZaGNKpN4/oed4x9cxCDAADl8w9S
dRGDIDk9vY3YqELZhjUox1ZBQSiM8wuZjizISgYBFxDnC7G3SccGcii1AguY
EcIhlVT90uE05Pk5tZOiGoE9kYWIS1xY9+CbtQ9wfnmE9kcAxdUXgvVKmi5e
6JSD4iNtJoP1p/5vGaaSoWBXhNhYpcgJCJdqVH4W0VRCkCmMGLR3zEJZahvr
i7MPE+ngUvhzeEy72hn/z/R932eLzBRD87sQXPmFzwrld/LQD7cGvznzci6e
54jBOsI3LDYqTxmXxxyLofleMrU4emuKA669sVyp0ZXNg9YzYQQh40Q7LgzO
NVGnbBpWt4+yu38eKLVxkuDfdOhgjM4jatAEKYyh+sh6nZ2Ac2nLHGbfJ79O
jSE3t3GV16NfhNQtDNeZog1LVcG6E2k/2DGn8GEfjkNG4QiKuFADqGGwkoWq
igyfSFvt70Hfe6nKvsG9ZoD8RFe6zO9CnUHk2qF0ZuVtiVQrpg9yBgoJAAyE
TYR4yFBcj8eFuAOMLBNWzdH+zVZsdkbPw/zeYv7jMH8R42j5l1/8AcMnH5HG
QRjwm6LM/tTIZDMAf/fDFuhDgFoW4x2v7oXMUy7u4X0RMr+vLGipjxZYZinM
odtazGa/J+yEmIl9EX/XyVwofpFPoFZgaG8dQcd/PIDW168ZwtC8WLsn5KDg
LQKH2BVzfAsCh6srQiyPJnulECJP70s9p+rApo+iIAvFUua3+XEb4+8nSA2Z
ENNOO1dNQ+HqRpIAmLvnc3/Kmp5u7PZJK9r4T/KKVTXF9WTHxH9lgvhnxaYp
7MAfrhb52GXgfQYDUNgD7c4Cahb13caGgtk1Efasc2sJNdEuwnZZmOSAAAS3
7yYjj8PjsVG2RIJJzcQgZiF/rPmq478L88jGEGyqXGO1AhQx6//Dc46MXId9
Zb1E7b4TGyD7Q3ymyDEl+SfX5ocgaYB+sGsD3mPIA53mVKnnwo1Ftu22WaPg
czyi6UtcVdb6OT74zJ80cbEu9FhN7+xlmfFKH+bh7Lm54UVFuHjYAYGqY6S0
XpngExR3zrq7kdL7DwUwITWTwOomF+VmVfwFqBRop/61+W+ijZK3f9xZ+pTF
2JMLciWHcQTvoRHiXncOEtsN42Ls6T3qJzE5rsa02umIenOqeRI2TavFlMjr
LQJC28xUNf4cSU+I+51eDUdI70dh1kuFoY46AjkKkFT8i4G5c+BYp/3nWQST
dHYOTQZIlHtmR6DGfOoSM/kZ7K6jCLxVV00L+GONXFu60UVGwP93wiJ6moB4
GIdJPd7cBk3MLOv/8JdX172UBFXc/uHoMwKyiFfIO6UpQDSKpeUvZBDVRDku
y/L3k4DX5S0Kh+jbjtHQVZRQZrLMm/Tatx7p/y6tAN1LkJTfXIl/cHjXCwky
8xbU+95rTJKvc8EbY79rihJJ67WLHpnlazZqCLjewuab4PIyx0MRgtrDHvX3
tZyFrv/Qz5mrf1anWSTF7Wxnz6C8SBkPy6knkCSYnxSTumt1YD7CSQ5Y4MBH
exn7B6Gcogmkis9fYWwKSO0gjR35rPVQdfqpQyjxXgHUgRyYNj1JsewTkzMB
VvjihmRIA5E98aiKRAb4XLGuQaOeSfLO1FiDIEjrbogi4UpMv7kPlrYDba6T
hEzE9CUm86k7vuIptxKZ35U9O4S3GELCa0So/3d+1KgzYn+Vn0Ng/TXRLuRT
+qZ5CjrNVyBhGFxTrxFELlSLZ/BuyKB+aTDhcmePr8pe+sBpZ7V/gqRZUWt9
Z1WHKVOZUT16/H5U/gIlyaA50gOC+04qM3+cZ/ZPdLHaE3uZ8poD8ew30Uae
TtiBfQdMzFk35xV1ePu55PgMPerettoJBVPrLNY/6ANjGwVpjXsphcSHfTEf
9SdjJ+yaZZvhttSl6XTP7COvNoKzDF9SkP2p/83UbIDLQj6H2KYLNONBh+xX
xzRxunOpNtqpMe3JC5AI/xYN6JQ1upzaHOPBMvKSJ73hy+6chW7ZwjiLUlLx
zQfRjbgB6lNPk6158YX9TdTCvIz8KvFnkZQq4Mjttqg+EubHfmqDIH9dn1Kw
EN8qLAl4RmP28xgyGsz1lQnilGrv3zEALp5J76EVkAfPmetTxthxrvEuKdK6
0qEX6nsisCYf9cTgtGWzVKV4WLdGqEz7BfTSd83rsMvZj9NqrwnhcobXqGDm
LIa7IDGAkxZ3WQAIPUyG36YnR8k7GB1F0cEsfAdzabyF/MYYDnyG/9P7qOxK
XUArDc3j9oPYy8JYl54tsglEDdJdHqoJf8x4gykqelgvINN3eM2xdN9/P9nR
DPS64KMjU99Pjp4H32Aip30JJr3c6yl3qG5d0gjpYDCZg2M7aEULTq6n1+f2
YCYuD+nq7ocKudl6QBfMgAnzT2MH6E1Dag9BiSIoMv/c+WY0GRyV6Np3wxkD
Di9fbafznHZYG4t2GmqOXKPwcwUHm/EPTB66CHQdqUvyvLbDQXpKlPyd57xY
SPT7hNWrEAQY1EYH6pjPsVBB17gLqGamwmAxUWHdlIgIs1zbz571FEGN6md1
J1dThFvxQrZ9V4TvVuaUmOk4akJa8zKdn1aDab0gYuvWv5awkFiLgNNKCG8E
Xz6i6bPS7rbtSr6NG8TxdgA6O+jgSXGcx9COzs8lbDKzeT46m020RMdXiG9e
bzrOfHbHeAbWIMG/ht0fnup33C0QbOEOtM3st3FCo24AFtC1ZUfpGaQZns2g
zKYTnFnZsHHh/Src773cGrIILLM9PXb0CZ9ihwFJ/zWSJkg2NEkU2wZtP/OS
H3lKMVW7xdIOcPkY8Lm7Neew3Ox7oWxO4+vj2uTjfH98ValYMFI5mrmsycPt
Jp1Gb94oFqgt7dhXRFOXa3SyGDmAgcWEuXA9zbWcjappU3psQf/R/8RVTWKV
dHWMhWju4nf8P3J5kMmZlGlTRxnYJM/jKc9BQMqaecRUTX159Leih1C1k1Zs
vwWMN8vqA9kmp39Y2ghK/HB7+aLOuydaPebAKZSFL+/m0en+41xAVohs6qoj
MMl/5jRzoEu3DLlCIA+B2TPFCnwFHZNqWwLo3J9UuCWQ6WTUBrBnPmDhgXfN
jY+oCl2w55a6mduHBEBANd1bKS/K5Iq5oaCt2y6AcbYNbqG6739rb0yBH1T8
a2PSTUOI3uSVs9A8sUiFPLVF2ufxoJ3sfPfSLQYbqDUm5u2hWeJhwqm60cx3
K0JDTqKQuXCIYZRu7DBhgxoBniIAyLJcac96jSI+QvW8X7oKI2DNXaOHuUuM
LP25FTKAlpQoDu4oF0rEhOO7pSrWTOk6suAxQAx8rrc4ByMPfCr9edaNzoVC
4MSviOInTXkscHMZXScTd6zrf4ApjBIO/FEDoDQE3tnzIqbgXCaXU1baMzW6
P29UHam1EsWqw3jCk2cS5KuUPo4kHdfbBAzymdNpdFx/PUlviKzeVmRBvIYg
+QiZF6lgTRApb94qLStR4h6CTBmQQ6l2L9UkAzQbXgrr4Fm6GcYxDB6bWzE+
kwIj0qiU8C+bFDUN1n4WFCrTvW9e+/3hbLwhdGpBg+6QMjrAQDmDAOT5Zf3c
6ZuGQ6daUUmE1G8cUWTbj1ReURqRLVIrHKwNQFwC/8N+PmOZIuvjMPaRiYwU
XeHGjeWuXbjs5iVEOsfnY0j8d85vFShtuXHfNRVcGt/zD9xZs7bNwDj3UtWi
cQcNuy65iK1p9s3cb7yGk910xovJ1Z3ngNc8aDBThDlllXlw/GfFlBrug58d
6UmbXm/mYWwOY+33JHov+U2/BdUCB7VIStmUPxmv1otZ8Py3Y+qUiU3OARzn
oYyX/NSpCPJ61FtHjAnsL3oh00GKzAqa01exM1iWXQAmUtC4nnZ/r2MPM2SW
xi1RoaOtO5UlGSCg2ldNn9KtyUvgm7ZoxgjTHsq8FDlmOPG5fOB9zN/oKMR+
+rSUgy1yr3Mmp15AJTAAqStKYgzJHmQTnXBFBmYARttdCRTFOMlszewsdRPn
J2QNq9isDIsbu8jhXRXTzDz1/WqARLdG6Gqb81o3+jCsEY+b3KF5/R1PU5Y8
SBQVJrbekaBHFq33Wj8bTcrCWfVk5/FR/h8sqU3KqYGsUp+90M/nJW6NWpPJ
0WeLfRLceOYoRW0fb40sJEGiHQPcy2rhG2bbzq5v/skxe8gguRMgK9MOIFTz
PU5hMG7aDh/RGX1DT7QLuoAo8TjvERHwF5bPQ62gawyx2vpPKDob6Yp7wf/t
fBhdqq/dhRXL2YN7/sWojVs4fciJONhRaR5Nu+RIliKiY1Ivi67VtgkyIRfr
SDVG6f+ypk33pkHufGjNXnP/yaIaoAMVsbvzBRzrl0mmXogT13lbvKugupg2
M8tpwqZJFyDY2YGGXFj+v3HUyWTZSgWI+YKA8e8hwadpu+YesoaBxRMz72Kt
fmaKStENzbi5VegN6UzInWi+E4n8NNxijGFj2JpI1Iu54H76zOTwAmJKS4Ng
gvZezAETwO0SNLM0y2NiWeSr8GeDquPlz0BTz5iuff3qY5RPJAjrV5lE+4g+
ZwooQ/JsOzFdigb92+i0Ed+1uPrau5gbg6/5XXRi0Sr/9+GEoQYC37a69lV9
OWBN+sKcHsCXvj7KVnjPbTWc7xNx4gl+T45vURG5ZHSFDD0lHMZqoyQ6USay
5FaxJ6ku6CELgOjyH9c7FASmQGOB56mIeSGMlJDeZQahGSY5Hm/xTBnjxQhh
x7BnBzueoH0Rg8UVBzQa1es386a9HPg6qCNSHoKA18U27QhaHzZYWA4xXAQI
3nMlq1bNcqTnAAh1QgJNb5dAmt7duI+9Z95Gdj+hlOrzmrnUMGftSd0JO+9W
EFCJKyvSObuftAUxJ7VNcQE0ycZkCqY7KY8iUQ8CQ7Ys3kakW6PtTynWnS7E
nx16k2BVZdTvmCVD8LH5DsmBJ0BsXe/CUX3laLsOFwn1+QSnD27qIK3ZEYfX
dNPd9je+0BXqBM1ue0toF71k+GQNovI0BOxcOQKfcwqlsTsqn1UeH8oYvICV
cuYrdfOzzgReeZWxw3emMMIXqCJnzf2nrKVKXOztpcmh+y2S+xywKO+XurdT
Q6PmBfG7tcp2HOVAtA1SSxrVHEtGfZLez0X92kWl+sAIQ0h/4ANq4/sV805C
wOQGF5aYoIE8vtxavh5rYN6PZX0OUoOmZP8g7Hhkuyl8POOy3oWZFaBxABbS
0Gi5Ca0VMvJYPXP6bsb4cBYIrtVRK0pGvscQu8qd72OQXyLehzILbWlEUSKc
Cr7w2h9pmxCuzcs4prbD5RuBDfkP0xjcgEixVjJ1ctTa0dopSY5lGHOGF7qB
GNFIzhgsjuOrI26EYnbP2eJekBM6IwVfaUJbWJVdeBRRReclnelq9FxpKGfB
irNWcp8IXx3S4t3m7UjySvDNcnvqq9hErj8/23qV3De8Ss5DAr0bmED5da9j
MF5tHbHKvOrc9C0FuR4rMA5xI705bsmTTqCr+N4iG+QHRTxNkRNJXMl9MQZZ
ITSKNrkv32elXEncmhygxV1lJnx/IEmg4m0pFmk+yXC6+nm+sAPwtX7/pgI+
i9hFrzJ6mr0qg6+OhkZNisY/+eAk1ryfVfyQ0tXdHkmrocu4OkpRWE1HWm4K
IH6uttmeECEyCOrh8Ggdm27fHENIZ4GU2Iqp+FA6Ngj/rbTQkZmoeouGo0oR
F3Xnt0ulAj/jp4u+/RuKuYssf0LhxlGimfGygsvTp3cdC5WmJaZj4zQaCjiR
X37c57ps9eu9tMGtqZk0ZaPAAtRavdgTSc0ms47e2b56t8HgMOLZQMGQrzMA
TS/v9E2AlR0k2d+qBf64v3T9AjjLUIhffx2OGjtDQVkYjJdG7ThbgHE8GOkj
vv5Q8bzVHNopYnTW98Oy8SpG3uPqD4atwv8hu2O5Gs/UGN9uQBIYhUzvoGDM
IULtQtCFzdzX1lEElbIkrd6wef8ht/lGdSpLH6Y5cSVkc0vSrMWBp9W11Rme
1FelFH15UoDi9R/LoRkO0yslKDvGmxQNgOWisvy1JMlKSQmVdBWc4/YwTMy9
Ssz/XjNVVk7NfJpKcIvv0WVB7VZnBHWKJQiF70ZG+RrM3SJ8VZP9wCm1oVy+
RWh5n0OVm9BAZb07YdPsPGC+TSG5SF578EUZGkolpw4BgVUQX3210BbzNrGg
LNJjalKq9ponxC3ZgXoFC/3ZZ+U2mhBDvx1FYeXW3rLXlU95QZ0Rurc1wnNi
UVbJOLrAEiYq0JJp4dX6EZWnGA/EpphUnM7u5Z4tmhJR+ihS1ys+LS6nt+Pw
tDFTJ6J6lq1RnexmRADjyJqLpJl57mDzw3SIpPikYI/zQIGFQlOpI4tSCMni
+kNaA7vjV/hwm4dvAj/HkXe++2O43eug2Ism3g8buRvza4NZWVFrZd0FIxGC
vYbITh95/JFp8MMF0hcWNuO+DFFZXY8ddPkewtM231nxDnKeIYe1gf1jPg7C
8IqniR7IiDKWZQPLs+7XcM6Ao0smTMjFAcM8dBnnNTrO8LOEiie3rAfIDz4g
BpbrHwMkgLTvjjO5XAUAlXy2a/Zl35QL2/boA//rClzZHcm4lf/UGHTpiUBP
vDE7MqYxGKpYQ3gW3dj4k5/vLxKMq9FL2y7+pfy7HQmD9AFwdUCdtB+euhKS
TWfzGE8VzkXrAjVDpWGuoIsHP88EW2LjfR+ZsOyH8rILYvqj2Z5x6g6A49lY
x3xzswqHXKNA02p4b2oSgWvpKEhnbrktEMxXRLt1ATNl339TsmDtddxlK11E
d4eCwgdkZbU+DQMWZv+c4Ic8Nvk58baihhxKoopE5CGVp/x6+mjx3ibqnEkB
VmocoxV/p7RnS0aDIEeAQK6mf3qEk+NcIGPvVHHHoTZEwr96qlqoo3HH802y
nOzwpf9yNP1Uj0bcM861A2h5FjwN836syfkJ0su5J2NJs6rk98FR7A2YI6Dd
PFCIl6BIv+xRJwiWzYTrhqTv3RYqODcwQUpM6lqc77PFoFV3zaosE+4HPlz0
UZv9S0c8+hBZU8x/Jk1OEj9URj9vaf/wW4BO6khoK2vBrq+yC9VyMxA+dP3x
y6ZYbw/Hx8Zgu9/j7cO9eAFGSsDY8c7S/ktat+8scHD+eg++PPBwyZNUcf7l
DBIBza/UxEZzYAF873OXOqIWqJP9uF1wcNJymqJpweXvAWosQXYpK4umAc7a
YqSN5Fr0normgj7YwO6lQVLbsNOkL9I5VaFTtGQoqE3ILF9B8RS9AigUcdp2
7hMpQJU/Ud5sAhgYR26tAiDq/POipcFxwVEXXAB0PklJ+3abyRJ2X/lBh2RY
m20PE/cXg0lXS4L3mlgGG/9OQ3pHli9OI2j4NpHwiXorchk172cmke7B/g5O
ekpK7nnTXUzPZiMVzrechvjszntJwbBX572omD/IFPdzLHxJYm7gdtYYA6dF
nxzO74++Tdj5pHI7mYd8O8/h1HBLtPB/pFKh1J/oHihPhzlcHogXp/oRqmmg
CSfjOoDnhiUvrwUBfW/LgzjdIucwzC+gkzr2ZxS4voCmi8CPBOvjg/57uNqA
nCVqUMY98Um91DoLRsu4FnK1+ELKEqjgl2lKgMMzi8eXFzFFSoPvcOCi2IRI
ul5Av+HDTcRU4gMyS+sJaHoFauBoEKzARcCA23uEsqUzfrS3w0oVFs0SyNmc
UFHlBV+u3CZX+4b73LB4bcCEO8opHQYax0pTp5CpQP1O/xEzsq2OKAabXZuN
K0zq+fQSgqVzs+CqmJQPWF/SO4GYa7k+wfqDv5iz4dKJCUIj6yUDvpc+WmDt
8PDzctFc3gMSgxxKXuy/oWI0/kvCCr1C0u7ZBAWRNWpCuf09wt41NkvLBEbO
/EGuwcj8ReMm04fkOKDdC0SWVeMeBDIRn7ttZLrOprU8sKnc6W9017DNkNEd
U6dpj9FrMcMTZ6lsb6tj3wDnS2vCAK42uimUuHAwKG+WCCG983OJu1EHl3Wa
KMWR0c4YYnabY/YGN9W57Q3W3ls1L2EYko18K5++KqAyN/fUmcHRYgFnAqWi
JiwsKCVZQvZwlpEcwjR9T2SzXv/GWzpSf7Ejxki3ClmDJRJgcEQtCjU1kRVa
rl8PIhnJ0ybUruJD1n5f3C2o5itVvpJNM2bFnvg788L5bROhvKE7P/zFRweP
ypMMwtUbLButSCtS7VDMiYr4EOy8nEZBVFG9vlkKmpv0sxnGWsla8XVYJJH4
hkFJgI50QHzPj1vbuIha2sma5vsoFJsjMyHRIz0XKr+yQPiXGtRyL1PyZYgd
BG6RUz0n4vucTK3lOJbgYEeFeRvS6pfRnASOghVyXEldSf+wDC7py/cSw1Qu
Upoq+Ka2BU9tF2HL23qClrz1YZskNGMpoQQuiyMydYG9NvAYWHbhdC4MgW3o
0KbmE9DaJZ46PjJCE+W4eQifgDjXUTwO3dwYsoEgRpMXJ7OLEP8qG2rYOmUc
2n55Y1A7Ik1XYidrr0gK6RYb55O52mfs0OJoCyq9H/r6ITp5omdK+HmEx5JD
LilqlexPHGKjXspLTIzcS3W5ONxVDTCbt40IgC+v9LK8MmTXdkvzMjptHLd3
dJcsbZGbY7ERBB70FWK4Yb1jdxwvDPTeGeyCk46QCQfAb/JznVmKZj0wIHoE
19BHcTZWYHXEGud9xSv78xzIdYvnqc6mesziOcnsRABp3YZVggl2JGbn9yHV
ZIZnQoc0ce/nrMg8NKMCOEqG8vtGyIlihfFiUurn6XuREnJWnx82j51vuYI+
6+izcVyXOl2bvYjkGJjnFq5HxMrWK9Rq0kYW0fpA44nFgOf1uvtY+8WusTJt
YhnWxiW/O5jYa+apt5h7xQ+0mIalqTYJtZ4E5IOSbt4G810QlCT6g/NuhfXH
qiJbX2dWK2mIIl+HJ8G/oY8kd+iqgvvn4R77vpiHJaaDs9A3nBG3ZMFLigg0
A5blDkhfczPSw7GOJ1Fm7UYPl1Ke/wRHQXr3W9eNj2Qa/6V2VRb9AUt63lg2
Lzwl5A4vFEsLjzxx58E1ch1aV8VZScryosT6oSn5paADbFQQVLzR4y4aNfpj
jvMOtx7E4irvYvWR2CI+QmNppgURF7lCzau/uLWL7KL9QQMb+mCvR03J5BOx
ftfVbJkgfve+y+aHc0q41M2rCsAcrnwXSx7w0MCuzjISel3IaQUKLjPGgvfV
CcTFmrGRsb/+2ND404gDQLQoaOKAppH/7l+PSSa1KXto8w98BTYMy1aNTzII
XYcoQzdYg882IVLTqjFC8xbVlP8NK3JexGJ0f9G9m2RMGbMBhIrDqHJEcvnh
UL4+9iL4/oZ4A+WQ3Ndmq+i5cdTeXpdiQ2AMtjyaksvuzEtJfPwZG9bfkHBV
Pe6iIgpGL/mlGgCnIKXJla1Xfe49vLsVmug6H5W2G3H/IIcrBIo9jSdQzsTN
DrpXWnJGu7KM4JYDRgwW8ZbOYqMpeIz/GatJnP5oC05NGZwtZsPuHeBf5aG9
BTx5ZCvGira9ekeu8Zg3dZ21jTwOGP3lXgTPvBcyzWrZ2jusitV55/++3fIV
ebZf+Xu0S+B6TfgwfOI4EuI3v4fN6eXxkvDoFSW4inAOpMmCWARL4MJtWuXS
DuFklDFe3EGeBCFV+G+6mcYjNEu/b+Qh3WVPqAVpPQT3xbT5jNJjxN35WDeD
DP77loAFjULhddePEjAAMF4K1SETJw83hVvklN9SMw2GrxIrMyCJUknLyo7e
8TsYy29F9TRMVWYJQM/pDb25QT26ZTec1S/Z93I4E4y0YXjJW/yqRnLLe678
ZK+oj6sXXq282Vh9El2bFSVmwIAFXaOPoGZbkLwc8AohvPiteQ2dPQeqwM8G
uFxzbQf0XC4F3z6deML8V7ZweCDsnDdZPB8o22Yd3isM9xKLlagJt/0QMGM4
l8WGcOTO00d98fMrCSiCIZUy5upr5DdQ1H/NMgT/DNLZKR3QxVTGUUiUclNP
LB6tqOBxR9JSqQqvY5H43R2rfnOm0H+kKVEux7kCjehuGCRUcyONK5xbVGHA
A0Q1QbACwtnKBKLyD51OU9rNhCgYsBKhIER3xbmvdLiDYFrJqJsKBvQA4PrY
RN9FLTGY07YbbKrG1O36NbS8HlUWeSY9m67Bh9NU8QYCybmyTtn1A7xiN1SO
qaNy9lbLEmFaYuj7tN5+XpHN2q5kcUpjWmjzuLw2ueAyIF7BW4dLv9bJVh6z
Fj25iY96nXi7NjfLVaIXmBsxHTOCQFvV8vc5QDwp6yXP+tAqlyL1+CnGB29/
zIlZtbYqc0FZM7JsXdjlNeJ4TRXVgBMbi69nV/SIpr5bgNJWAJT6Hr00nQhe
f6JGeandlMDQdQEGaQTBPDe9khssfHi5JB8FVcRkxNMgUo05o8NoWQVK6NPG
Xt0KJ/WV0tyMsplw4cjBe3FLPYdd0vDOBddOlfMG2XzkR/2LV7y5XGbY/0rM
SErYafAO84+3lzn7g/F8VSck/RPOSlEfwOnDcHIB4JGZmYx8NaSPs4pg890Y
bJ/c0AqLIFxj/rgeFLBB5pvf1yVh8b05a86Ys2bFETUrjQchUq5a41BXQ5kP
X+QSZM6qA8ceq//YxMb1irlV1AEJgLuV+pKy3uwYR1eJxLm6zhrZOjuRfkgv
GRlcNMyBZkRHJRrZEwjNPIWagu+StNzmZSywXdplIWTX0NkUDVH90Mk6VySI
dduYl7s6UNhvM2G4gO5/bksCI0KyIZwhkmQHKy+UY9e+Jt4elfvRLhWRp4Kj
pGqxHs1nx4K2mZpeabZD0J046dWsnnBQ8uVE6ob5J0DMwh/lurTZdwkybAPg
x3XgLbrq22GtKxBc3xr1iqhciY5vNMSEcgFDCxunUe7EDs4BShCbJ0RSdi3u
LntOlIvIkRcV14bRULMBqgRyUsiB782y1dQDYBBJVP5UqUc0ByHOuyFuthp2
X8vDEH/EBtK04PMjwaNqH1mgARCdp9Mhox4EKvcKscKBpUuoLsK2BjLWyH82
gPdYHNBCeyGQBAUi72xtedohf600Tph105v+8s8PSJPtdFznmsGvif2y8YS/
H4Disl1BykMid+44mU3bjHO3C1QZjebkLiEtHA7W2wWzqMr+WAeXyK8Ea5Oj
Md44iKnfEXAELpkPt378oS6VK2MT5K4RRk/II6VGOp7bPbr5LAB218ak2OH2
NuQ2HzG0Qx6DIS5ZDSZPRxHoz41GXAEoBNvvPbOj1ly64ZpZbdmYVEYy6wwT
PptcTKaU3tQmKW5mMJ9XPJv9u444gN6Qx+94c1L/TSWUYTlIf40YWb8DCblK
ATyX16H9IzOtBroqMH6RG0vxZV83TNd/WBKhIAVIWKfhecP2BgRmN1ZdmDbp
LpCv4GQpm7kz4kiwKsaPRuc40iHjlyGHUpHDKUEJ1vgyxmfSesYiMQWc2nPV
mIIP2SuSqw3otq57w28QmtZhimREBP0HWAsr5AZ9KSHjw2mhGuCp6K4/6r3o
Wrj5PZMM62QXrkFebmMS2G58QLNOQZA3zuBQzSqGwEsF3JE19P//voqKW6Rt
HOB4C4pMVnOvirl8UOJclYm4JYuC8FAj4G0vIWMxYmI+EiA6BKT75pDL3Ef9
OjJzNm4myMtMNbPu5Sv9OZw2/RTf6REJYPNrsaSlC2ADCV8xNmsp2OOTDed4
3yVkVIBpEafortk4KDid4ae5rZ/YBypFEj/S95fG8xjNQaYyU4SaryQ1fc5g
gCwlwX+bk3+sTUTEwHYQtkJ8bjl27iF/HvNKULYUC6ZSYUkwsopMGSBhAKk0
wCLfJDXxj5nmeUiLM64wm+6cJ5oAT4uXw63oNF5/o5NRZSR1JElt8mOjkomS
NG3M/WhO7UPZTuog3Q+VmsdWEhMGnZYOW06g1eAFWCtiA2MlSzEff/Q47jLu
yZkHw8iKgG6pK3UJ9X7CCf4J10sOiKYlMAxV3IwPRp96azDSR3pk6kOObk/L
iiwE3nxrBdHP/JdAKtLVzLIqq3tv212/PBpTYZwA8d++6nTQbNKAfizxEBAY
5jpv7aDKLjlrJiTXans1Bv3kj5nMBq+zjn+vRY53cdE1/tl2RnmHnEbwl/kt
FH62ny8rys70Gp8RhAcMsu4Tzxz9ctwQ/8BLQwEx+XDK8ajEXi7VvHsSV954
b8Zfj2R1DcllQhXyZDr9Ip7CEuzsYNE/mZMuyf/mDL9ahRvnsAXRhgGzeJvI
oB/xX0i8Wl73b1eToBg3afsAKtxvJ2kPIsGH0cqVttoGlcLveAUPQwDZ2E4k
E9JRi4kbcp40u4sgfxQbomhsbvu3tpRTISc3ZE+ricoPNK1ta7LQKGIkwfHc
PiS8KCbmWk6HD1UYdah/ZgfbEa/zbXAHylHYIU7fHVmLvVQL5U3EWNtFScD6
R/AUUo/QGsTaHIq7f6WSyB4cmqGUM5+X4xJw7UQygDzNoMvfkPBxHwDzfNul
01XH+rYw6xHCqI4oLBJdm488Q8sObXtAXMogHTxN91UqvJUBb/wnpJy9Zf1i
TyPFQWFkzoSnJilKNGi+LRg/4qiBqXNCbQkTpVgZZZrdY8yL0gaNoxn/w4tM
13Vr2V1vrFdSXQjS3dVrtqZCaeckbPkWXpEriB4mFnrWF00wNd4MRd5D/RTU
zO10r5ZTv3EbJ11r7r9HUQXVabGmve9kwMZkskTYtxBZPyTdXiMjVeWIlDeK
fNh6GLxoBsDXq99smuigUtr17LQ7p6e8wt0s7C2yHxm1iq5h8VRHxo5CaBMG
hDdU2Yn2ybtO2H2RhNG7wQRsZGsE1q/CprlXNSyVcFo0kgWhi9COCrD5tYBw
ofZKNviYFWGR2W0L3nr79c/7oxyhdZfElyxv5BMosXPy/6aGy75BejfULEaB
oyQjySh88clyyTQok/WeMCx1tsozPKLrCy8XmrYCaoBtqfe5ax7kTdSu3hCR
1ToGEIFKti7nO4hM7vPJX64f9+iI6sGy+/MtFmoCRhVXO76WBZ583/lBWBud
+ZNsVJHWCgDpojvM8BKsfmx94SafkVT0WrYcsppLgmbBPHCwQZFDuRLoxllN
0k4xkmpN635NhcW1DQAeHkAXWfN22d03JJOqxvkLsMsbCPL5mGF5EOF7EU4Q
ArXJv+3TONuaz7eHcyrgrRkgqlN0xakUxdCQBgmZ1YIdLxau6m0EbO09mxxp
Cql1XAwnQuWTGFaMCFDgexXCTo0uiWR+4OfN7fgy75KWLVyiT4cnzXkBhYlg
tX78QctKd2bEPiCw/4gZ6r2/LPhMDNSrm3eHi8PkUh9j9rhisknDR4OIXcTQ
v2JjdvDnr15jElDTyfh/tfWC+N4CQM2+/fSs0IkpxbS2X23NTyGN7QwIqvpF
8y2SGQ/R18Gp3I6AvpAcnglegOJlTcZZXr1urgLysvt5oYEco/Xia2Fmjxum
v8/VSo8UC6/GXltiYGEsJ1qYrEwHBkGLDEJ0VIgvIG1apsKY955n2AR97BCl
m31gOqHEzumztaodawOpTAztW2HLa8w8GEuCPBPbHU5tqREEQYGI/7eRKgpF
jaEGH0HEUaQxSTGfpx96KJnsrmDfi+picasBH631KeGtFPd9muEhOPqyYT55
Gp8LQ/wrn7ITh5Srk4hvVuzA5txYnnMXN+xKLzqmaknwfk5Wr7a0jeufKvBM
iEMXx63euX0RAzi7uDLzNWMzpPr70ApG8Bv3aAmyVzWWkvAQlVKHodWbxxXP
oR4/rM7wJ4KQ+k0K7tkpkAp91YQb1mgQe3nFbrRGRisuv+BYwyTPTKZK3qSu
hwVSwSBZC0/014qxXVakFMrm47BtCWz/2LJPX2lIxNjWU/CdBoARSQ2HG/wP
0Z8K6zb58+uIe7iqao213ShRCjW/ffmazX9OCofpaWPi7fqr55XRWvUzOz24
xFri/4tRbw6/ZO+PqTC+11SIkl+1AkUK4XTHhS17isO+HrAqsNlAO1x6fFwk
Ava5Om1z27Tl1ltC4GpORvsZJL6/1pJi/G3xFvGSbocWcB+Pni8cBI937j4g
tJ+QRqYdjxuQyCgxi61sxEkPr+WIjLaTRJbcjR7Qucr7/TITy+OYSuoF0oAV
lDp5MwsXCaa66XYCaxKZOhoPdIswg2MEV4aEHjAv6qqILKRJtvOfioqxKOx+
C4AMDCmmq/W05m0cfj7wDquWmT5XUphK+Lsepvyi6U+X/rPc2L2AYOSi/QEz
VdzBxjuUQoG8br7Mmp53u/1HBLMIJypujcojKBNXbf620rbla21djqQOKNZt
YV1q3Gsyn1oMdqgCLELBfbg8SQUMoaMVPnN18Wbfgq2/xGGKGytJtShCrsjG
csiGicXGsKjl/KLT5wQGg8Yg9Dl43ho+9RqlBPY+ogN9xullMkNiqlMVomTE
JZZ/TDs6pwTZaIJSW3Q3j+bgwn4mydUzKV2uKQvTCnlR7byao5183MoSc4/+
q4031C+YJrF2rbQ+edE7MCBOksGqb2TWheOCO1XUrUcr7v8GLg+FpQyd+obV
qfMZqjnuSwEt6HO5BAuquG1MogXRpEqgcpu1SIWZDS0QOsfKJpvdWBNkRh6O
BosavBN+GR/NL5bbBkbx+sRhql5s0uJD5cbcvt8UWNAzomXA0fDJ+V919d+6
/9PduYIEr+sBZaEg0KjwBXizJOL1qWoARqMB0E3KJNc18ppZ/vd4yQ5fwIH9
STfUAwgJQQN5tp05Gt8Ug/EId/MjPm5/mV8b4Ar6DiTSWtP/SxFes7xJOXo8
Jc1+BQGun1Xc72yDsbnl3QJoQn0i6GO7gBDHyIXO7A22d7Orf7aHYp5M9qal
D39Z6j9ATq6G4L9mREaRdP1d38Y4XbZYKin73XPBh4FeCCmmdgUr7rt1Rxop
U37RWDw4V/qkvjDQJoLDdx73boBbwQSi53cEfKXRZ/QCRzGIIA2AOcEash8z
oxR6NznfXCbi+G1neEHX2aFf4aKyn0atefm9AL9Sqk4UJHV4DFkE//8uQEr3
Hx0SP0T951GSmb1hj4zBwyjoorv8lNI17uxdQBhQe204FreUPs3to2wgpMXY
wJpRQrBxmtVuMBGs9hDE3DOoYdxXuxb47XCR8aPk5N+tT/oDUGBUl5kTZO8a
w4e3gHysFMXh4CkQGSTjBfRSH3r9NiAyT79xJF3al3HrfyT9c3Tzy1epOzRi
PZ1DDdkR4/n7mIHkt/EOumdP9YNlSXVIITSUymU8MrR9gqqhdT4sljoJlp65
/DqomIRtKFsqpEQi8ey8DVOY5aFUcKW7D+n2PL9OJ6mIYicuKNmS3QjK611M
O60r+loUFwhlyULrZ7BpG234kaSiTJ2N794n/c64kus6J2p5jLJV3Vi/iDlh
lROtNUsKU48SwBRbSTfkdWLbBWd7msX24dx0lUsnwfTadSqtf1trLFkoLuyK
P+Db1vgkCBvRrqY3IVoflbhT6gIjZMoFTQZyC7OERc3BZNjKq5LkQFRfsP1+
FIY65QNPFz2UsVnepYYAyesZw957X4Gz3GR5U+ELVNd30XEhQwZ7b3HbOxbu
23J13IyE0p//NheYA+w6dAOGZD8+ICb+zYagQeVT3h0U+91AdxJtaDbDWgu6
KgSGou8g7iXC02HgnguL81jAeN5SrwX8f6vt7SQXeJCjqhBGdc1oHFC1VUip
xIezSKQGIQwwM5AlkXtEGg5qtgtzx9EzReSupPHDcUAT1NiIymA4afDU5h8Q
rn5IS8Cbjczbse8qKicLZHgqXdAlYPXyfw9bx37P1+/YfrUb6AH3cxWNClyh
7HbxDtXMO1c2z8ImzaUuG1DQCqFZMXYRJcWNiHU19WeU7M+EIgpKmFt6OJaP
NaRWkFbBtZ9VTUKJ0NwKNZpoXBp5O4BvOeSh3cCM5H+XD9/VO0TD2bC17kdN
rBfmaUn2Py4hU46ezG9ZlgxDRiZbF66poft5UYdmoI1qPd3YqWSq3Bg7uOD1
aJLyWZG1+ajcYXDFuoyzrOMi242rg8pD3FkNPWCAMNsFCIpU5sYEJvguM+gJ
x4G4MuX2TgtoSvaVPvpkewFkixM4ScGgjC0siZgQfby3WqbriBjjqoNIejpr
aM8DwvoviAciFECq4owE0fhRxmR1Vuz3KGSmG0MXNu15nNUQ/c8kUZwyFITD
Sv5gDV7ZE8cErKlsfMEd9hznHms6htf8r2ciQPt8qZhkKdOJsT295+EdJWuK
XLa0YWG4HjkDFBe4TaDpRKwXI9CBnzUeA8H3qXX/NzVMGl+grO0+zDo8DXgo
uG2AwU0s9erNN1LpV/vP1NuGEeIx1EO3Hty13H5SXc60TI+0OwKPTD1Hph9t
CBWDjzABPuIbZNLDxEVyiLtxTuQTWufnQXtVVmiMdDnEN5fUVxrzselkWVtd
NB709VZwboXIrqA1YH4/8KRzCjPae2KWz2axX1vCHj7Qh25/rbJ43TEMj5mi
3T3IlshALx86qxGqkE5oSiWjBH8L5F92mYXhsPvoemXbIhFAuLhKW52YpJag
UyvR9iKmSQ4A0gmRlacR/p7+4jIBVtpX2RBtPbhQP55lYsUBDC0eu1wGYqcR
LUNKROYMASUstR/NDH9tUT2R1prg2koUIHnrjQQ9VJfZ/5fqu9QTfExk+j8X
WA08h+VXqqqWzXjBa3bfQDO62/pHrEmDanesz0g5Q+K4vFa9Bs7NM1Ow/ohY
QUR4qrY8IEBm1XEdZahcGn8ydk9uMtl9sKpipIAAUg58MMA4KsFlqguDosx7
Oio+fnWJB2kOM7Wz23ATJSzlUvl+X3ueBfIgRbB5lAAFpewsK8GINdGllEgs
XSaE19QLsbEY7CJiRMOLVDZXO1gmv8+njuCf4gz1o815Rldh4+vuZEKwGbHH
Ztu0V3fepwoM7zUhspotZp6tmbnzjLylrlfL+m1OHqLhpJ5sTXGnNxYk1n/o
LqrueLFvqlj3x0E8z2FJdJiqZO92QKyCDvNwryXStAGW10Q4Xte2/eDQhFdY
Pb+ip3sQn66YuFD8HKuztCge4cpTEMeiIuL2lXvyJyt9bm5tlLEe0TS+VRKN
1EbPh9AyTL7YrxwXfvTcz7AuYdwBdrULsvf1IcSPkDeJBGkfeuceDX6xbC66
kHeduQn4A/2i2Vy98yC3fpK5lrzoNcWw8GccpO75nI/d4vqrId6+dOnrzG0Q
2/yjnRfo6qlQji1GYzOt2cWdn68GWMNqm31U0Rb9+xEOauvNDHyCsnkE46KG
5Usie4Iv1ij2tRG8+YGwcWK2GrHip86zgReCPJrLeo80LHXV8frMedG3cPQ3
jwscGHL9rrf+99NPfDuVkti0rtQ8Ki5kgxsyZVQpc48SNz+TvUEgdbs6wID6
ND+5HoGTc4UNKYV+8f/6ttAQy42pyEjILNoqVjzaYfUamd5o9KvnC4aALEhz
yQpmYW4N/lIMXo8AzV454K5UhCTdOgxk26+jGc1G2mocrTCa302CQl6gjlwS
C7Kxv3m+rQt1MWZneaf/nYdx0yB3KFGmC33yOjl7mN91bUNTb0J9jbI62OA8
TL+HK/jq3Rzqftc/w11Zp946zvGfM6S8wDWLMWaQ03Ne69dgUVvTfe/NElDq
+NnHXo0QuGb6Y4kIrF2dQNDrxrZ3kF4NcnaNQzI71QgVpKa63gnmRHSuEFul
jwstAswuIu3qaDpc9497H31LCi80C0Lt4yecpOSl6bTMcm19PdRAm6VJ+MaI
Kk1em6pzl9R4qAEcB770unejtciWGQnr6CA9idAUwTqfRB23vKGMuNUuUj21
M8LF4xNe7/1koJjzTLCpxy23xzTzt6R4S2vYon/xBAViY17oLGac49ZPVaZv
StJB6j+o5+BBn51T5Mze4qVHPUnXA7A76i3LWOiFg6+EzMH6uUuDNst+4NSh
p5BOOW6QZDM4QsifBHrfQT9KcxWqSQDmTxbmEbrG7ga4dR3dmi9HMURWDT82
f7A4aLtHU38wVJdNPtM6zplO9PwvxL6Ze0CFYPCsG5goGrFa2SINs15ytfdX
3NoLEhT23EAoqAvLV5Jbd9xiZJVsA01Cz5VXcrSXuerkN5n/SubJTPGSFqid
8u6JBvZLKzTs2jRDwJ2xazepssPX1vVsVcxuLWs1OtA0K/YtHubkOuGpnsNq
iXYoRqP91R1SyMvvhxT6OMi6pcToNeZ0vKxsJgEsN4+9dqiI0TAy4tp4p7xa
fklmkeqFcLutqQhQLFLFfGUF/a/BUwqNddJd5mhbYtGOhGN66XSPIwwTeoRp
tBzm1f6vHsxcLGTDusSPvSaUeH/ytx1fqcurhpPdQHzEcqnpHZjL92y0ERs2
/gS2gsanbZebJUrB1QIhZ/jYqG1lbe2dC0PGeRvY7QMYi752owXKez20zDxo
suWSuaWhW/WrwMvShLYvR4IgCzZJbedubz6zZlm4hvXSrsjamDuOGd6GHX/D
vG7rQ+SAyDmsEvyVvLH2TOzNEcuPFa/m7RamM+PJqbSAfoxfK3XP77+vMDIW
cseOiAOi1kfybyAshyg/4CEdYFXUtPWW8zPg/Ygn6Nju80lGziGLmc21ZHa9
/M7Y7YrGdKoQN+zhfm7/TjjIra6HSc+ch4CcfON4gYsiFFXCLNpKuI0P8jbX
ubvi64piZQJUTQhj6I/9lsK8KibVb2VzNSUwHYTbLcdcFfiAIekb9WYYhNnB
H7g/SwNGh9b1h+x8CjLDzluAilalBcCz0RrK6loeKlvq2vMHCGX+R28ZrxLB
4fpDnfT6g3M46+gHKuV+OjOqcx2cQ2De25733wB6Pc7bRnAkZFncFVrJhCfa
MXNu4A5FRyw+OXAMbLSvnAYiunLArt7rE9yor2clavOUI/matNU0sFCGu3CA
scHPjXA2cNJ45XASfsBa0uHwsSac6Rtt1TO2NC+3HptpKNr54wxWljarLqWS
whceR86dr8hAJs4S3Wbyz95CZ/1EHdmS38cRoAK2iDWtY2veRcPL56f/Ej6J
zKe8ROfeO3+0ijJYg7dN9yF+L5tf+a/2PIyhs63rs5xD93ZwwRzhef9D7c7W
J/f+b2Z9xrkPnxKqy2yxjmZ5COgukiKwk0VK7A1SfhJ0h4xr1L84Nu7BWgv/
LT0V4AZKrDHh8j+Tiq6YFHdz0JKRq6KyJCIyhgZvxpkR6yri0YI1sBSRNRqk
Qyd3rBcl7GBn/mLTnQQcBMTruFPxIn/61FKohkCEjpVnxz042zMX0VkHjEmB
Urj9rVHYCCgNcTiqabt8rnbsjL1anUNY1h+sQYTsM55OPx2FDnQAu/AHIYf8
nJOCsloGKqv0jXCLcQjn3DaJysIHJmvZ02N7/6H9Gs121A8xbQiH44PBKwjM
iPzJaKeg1+ph6RpM9QzEbxIRt+Ym89urJ837KXaz6TWAtZLYHrsESSL0lv4/
/+DaBjA/mJCv1KGScET/Cy0Y80bYSjDhF5IvZBHR7+bUQe9D6LZsTtFYRmmA
JgVzBOyBwzHSM3JyfWI/9pa/1ru7FLesTkUs105OlvRlmm5jvmI1JeDbNvhX
pU/OVVm/hdii81/+u2k6Z/D1ZZoiCqyqLPs0XjSDU8RSWpe7Wq74FcE9poL3
JyWp5jAdFKOJ1JaeKBBa15l8RSNWzKEppBF/9mqdaCBpnwWaejpYw/ARXwB5
p2xFobPL2vkectjqx3clh+ehDmk7M4D4+Ps656U3snOeG0+6+fqlWDAZI6HL
mbiug256Ez8zTnNhOLnA7GiNwh1szc7h5x5JMJAatAXw+yRx5GV466N6JeLl
/iUspLnA9s4kOlQOZqPgD3tGuHnUsYM9uaBflFNgFykXhblW088QYt5fMYe8
IkggfV+z0GJ3RLVr8lDbY2eXwtmhBVgWt/pQxq21RYcrQuNaVjhU6NWd0bBt
pTGQSwk7yecOxGNEI5lfEA7+1nt6p20G5fGBFejlH9GyafSn+Cz51sc9gnzu
FbuB+gtPbh8SXQTgt9u29XvxQ6Yljx/9CiujVPC4U2677/xTpLNMwtR+5Qjv
2DHQrbYS9Rz1PTre2Puek7vooTbHAPCI5EJIkwLp3FESl2l1dErtRhxV8JiE
AApxyA2xiVVEg4KCvBlZ2ujaQaFIVuVdXQfkRkBQVxlwQ9p5ZcCeKTMrqQpZ
zIigfp0bfLtdp6qORt3Ul65K+mnv5o55R88xP4/kOUlKtVeV9qomj02BjR0a
FdXBOTE6/JrkHlI10Yiqei2ujxaekV/KZMrQVygMrtLQqVCzhjmDVeDuqQ8u
S0/ZxubwBuc/zXx2QuQUtgmjMnbFQoV3iEazwN3O+myJyzDcjSCAbSy2OVIg
E/571cskAI2QnE3NPewIvfFI5SWSHCLYEWX0k+iREGOMfEhpeSPKm3VQI1b/
Os1X/8xUO4do0uGf+H/egUAXeRbC/1+N8B4Q40ptJ0Zmmwel/EM89NqAeBRj
Z/zBS0RXIk9pjI+RrbYLL+tFi2bAJ0tQ64wWt8hGru0J8xog3uioJQA76gqI
x5JVDBExfYzh++711mqrOXdtHGkddskOmtx/fmuZ3QHRi/qugppTOgaWLqoI
LjZBy6m1OegpqnZ1yPZLkt/jCF4zZBCiQnfL0hN5lFiflQQRxxi+GuUK7C1M
VnIy+5IkYRgPdXV9JcxqRZyMc77cHymRYmjdErPgg99jWJtPPv08M+wMEVE4
SBsJ2KWc4HuUUviTIjxPGrITmsLezw54hBZXydiKHDrIgsFX4pfxoQpoEmTn
DYngTX+xaL2qLrDUD/MXihs3PM0xSxufxfRwESNQ4mu5bbYgQ68K0PYkQahK
+lAMpiMCBiUiGCZ7dlu3n5T9eiK1DXkS0uwd+z11JSyXpkq9HQ3Ydit/mVYr
kL/+iaROL6q/bdSfl7V58psiaW+wXFBdUTp4M4Q4N3aq9qXxCqCzKnUncNL9
Ji9a/rnpeVDPOE7blIsg8vSx6f890z5oto3l/B0wpvCTxiqkb0FbZkbhCfti
Ad8a1ukYHxRdiGcb9FnSx1C2AVV4LurVyPprItPJ2oVXJz9w0wWxl78HRTzM
nmo82G8ecxMApAAT8iuOJ/qtd3sp0oXgT/0Dv9iqqkt1VfkmQdD7Cn68TzJt
WBLkqF6I9YoQ8CFxIen19KVZCbuXYfg4l0xn5bkUwhwOtt3XeyaVpWxMXdxZ
LcqkjEBuo/Ne2rghjKEy2p0ldcs4LKPTqSIfnUT5UBYmtKpfpIJHrBNSoL4/
uExsFK0Ifj78QlXlKq7oJ4ad+4pBMos2eEtxE7KQM274gV2oDcMYb6ZYS/wC
C/GpJbu7dri9IGryraK7FfFwIgDTwel/XjiDQtxU2DiTQZbiZLJ2vfRWBgkR
SKf9+rtDmmUcFwMxcZWFEzY/6r0kjj63K6UwTTgEoI035zlYu58/uh+c6Pky
poIy7BfkK6bBp9qnakC4Zs1hCX6ItdIFgrOQufCVDpoZ24oJHywijX5UCK6S
c1zL8dQX7E0vVmpHkf08IYTgSQ/SUypEOIul5/npCiFcn9hW8grdjLJP2YFA
6nvfMtuCEqyPLa4QE4NMRQem8S7FDxmp4CbyPxOZq86DSzulVShNjCR7biPI
EutzAI38UazpJcBvVdEzGmqmCJ34phQ6VrI5kPQvH8QCV57sn2FXCcgk8B7M
tRXcSGd5cuqzABcELikK2EXfcFk2I2Jj9QvxjBjq4swbjUXJUuGTu7VRLaPw
X+hmwUqzHJ6W0PeFebsHNAQ46nRvoZkjm8txuNp4iyTDTxhjfcJGIuWSz0m4
GRp29WsK/XlVah5+l9IUrcIeq5g/F8l0OPLLE9sgfi9VhBux/4bIRI2ZHAeX
wHtJcbkub8e7jyOlt84dt4dpZAdu5ni0wy99BGDumO+eplw2r7N4qtCoKmXS
B/rTTdWxWjeu9MFlogIt5GzCQ5xtOJMxad7ZdiPKX7eEzOfKuWCyTR3BZtri
NSObKWFTwAZQvQgQ110azUxVj7zk5iB9fVNXudmuyZFLVw2vGAMJiKWt9m7Q
Eg/9hje/V0hv+ShLrZf/kOgAwAJTeDQu67XwNz0m8NNJBz8xlWe4iZABhFsP
AwkS42mGcCaM1T7W5BIKVM/qaFpGVAg39G/KIjbKU26iQJ0wZ/s2nuToPS4q
GZzdTHURwg7yp67+SF/sILWVzLZjuw3gRb/I/3+QFDaUheIyfIT6xOHtb5Xw
LrMmENB/vxzGYsiKVE8Ff1C6kHfwNk3t4IMQSsezfa7GQSgCy7wDxkxIQd8K
zdA2H+NhUdWBBjAAk0Or56Qvwj8Y32TSii8993nneSOBLcn9WPl0hylyASG0
blH+FY8tc0QnupsqEulxfvg26Qpqq/P1SujdvH9eFmQvbBBFYMAwd0l8TrpH
VL31aFlwd4H8t45+4EQYeQwaw/jb7CVJf094OFPXROv3qUTE2dnxCCeZl24u
2K2JFFaeangNhJz1hQv5J0Sa4x9niS53avd0Dd9Lg7uVUZ88C67rAXQfjge7
TCTfeWie1aDhW66qcPJDkrnXaE4VNnjU7XPcGWICx0/YyzCS4KDSll+5nnJo
yxL0D4FxsC3TGwKxZ8qgkN5kQk8fObP9QepoM4q6i9ab+kj3P8pCt/kHEc8R
VRRm0pcVM/2LGat93TfMiUj341HSOkicvf8e9OQuPYhc8pTA1lAHj4gkEHK3
SttxvAZz6iDbnrQVtCsGbSyihWCtuIU1oqmzCmKfZvIVJ5Z7fwgCydRS53Hg
sjeJ0FEMd81qam/og/PEBqXz+h6bBVaax58tSbV2Q3UKxcUHwzxIcepYNwsn
3DxT5obLxMmYXzUtFFwM9ccIp/hTmYKpj5anQjMyMj/B8bMZl0ws2eMzjGu6
l3WB+Cyo0++NLIcuXwzwI/B+guFImEFwqEVcWpARctrAyc1rTQP6ggoJCVxP
lhyfZqqJcZMujaQAQ2Giov7THoPaKS7ESupOxnJzryCG0l+r2I0rJQN5+n4L
Tg20+AMjKI9WRYmzIC6vCHmNE8T/7gMyoCpZoPXWIISPffk5HzZn2cq18xp2
WoTZQFOllmJBHCSWD0qrRMr73Zh1vUC6Zu1WFNU6lxg/AVSVB1rWtHGSS7n7
7kPQ3HDECh9n+TELWiQqgIyHSba3i6UEfpr+1u+I/P3cpT+p+tsCVCsSXcDw
KU556soqgkDafNQ3fui7f31sffHTEtExQGoUxuBosgEANmgg0vvGWUt4T1KL
39u0TFJ3+ozrJC5RLhqdKLNCnXIGhznIBXV8ngAwmxD921I7mfH7rFKTabWW
OTmAKQlt44PtEgPn+uc76JJ2pInhUf7oqnQKKRE3ED0+aZWotwd5+oVFtvHC
57cMBIHammEPO+NLt2uwmTVNm0m7rQU4QeHH0c5TrdNSkocmgs+1KY7Ur8k8
cK+gPtEAxpHpuxtPGzJv5W+jwJdPkzlHheXkSPPp7xAX0BwdjDDIXXVHU7sU
m19VWvzSv9VkTtt0OzbZI9oqZ1XiuZa8av6jsr9UMXIUIhMLAKmPcHz8xzzh
ZZSM6VczAugSDaGp50FVl3P+WVsFT/SFfq5G4Z2R+dk+bY9cIn7u15bfiwH/
oG62gcJoSDe+zLPinVCp7Osqqb02jYkmJ/x4YpI4lbOqJ36gelhPRcK+Z8PM
1sjku4v+kSdIaWreHPBG4bkd2nGkO5VS+QR0Z+ukbw4d959JMd8VwVhmVabk
xCFrO2N323mwRZAiQk2PjbvOqeOzA48Rx0/0zw4GycqbDTqcNHN7GF90oFbC
W23NFJ+EZNtW7DzR5BeyHMwRQi8o94kO23VgYLkqFTOLJGHdPkZFO9GDKYRx
5CJSfExl0pg7xZgbH1UHmQPEvETp8TVAhpyJXQxVXdsUu1+BpCMAQ3KUwvz6
iC1lWVV0PO79tcP4Mjyp+KoItueYGjDKOmwTs3PX7vZ5XAyKH3/3jZ6bF8uI
kyiMumv7uImuSBj2zjZ9GS3UnvdaNHnOMjcoGjIivHN/G7c39HpD7emLDPF+
d97g3dXuiFxzJaPiTI80isGkb3frPtoDop9VGc4F+DQmdx1MEmB2c22/+yBk
nxnz4wExDd8Sjv+zYT78nd7YqnLavga5RtKYI3/fCJ9/DSbN/Het847a3KSQ
LVn9tLrnUhB+EjpziWh8lnuhHJJevfNsr1SA7zHCz+PISQAAq9VDh+Idb/dU
0IzECqNMjC9SG9gwp1FYNUmUCg2KGoT9OAvaeZO95gK/TeYgnDynt8kKZVAA
YdmHb8z0w0ekcPrOPn2DMuWrnblufOxWdbI9ZfSodujkQyl+860bh25bNKJW
XsxINypoDo1wJ0sSC/N7pwCElKtoW17d72pgRbYFXjxLcm12RtL2OOx3LPyv
d3WN1jffoa1yiaWXaFXZFRh+8/SbdeC96Ip9MGKtFz0uQCn4hz0MKA0Fj/s6
cMMdEiQJqpk+r6itdI4/R5RZ1103MajF92s7gbVHtnvOHfIGGhg0M0RyBvlf
K+Rs3y0kW1+sMh60+c5vHtDYT/kj72/xUwGj5MmBuF86mc0hpkZxi1/ue8Bo
TcqLZGnRogN45CtG7SG2ne1toF8aBJrVMlvDGige3ZqUlgmQk/hYc2lBEg9W
bbI4rPQXlZCMHZ8bv2BjxAHN4MQghCnssUDthyvBnK12T7iYIYZ2bnvPyKz8
0hpj3adtwAGmaYVcw7w/2Ux63hmXEV50+a/50G0gd7G7YEJ0J7JTHQmCS2cY
8mBnIrKjhN+26MXIF2o4Mnwhjcuj1RNej8Ps3uo0ZJrDAeOMQKyAuV2K3c7i
t6ojawkr8seSFyNgXV1E2olYWf6vksMgS270uiLiOS3ZTIoLUPBe37QSbuSq
XwM2mGaXILELeKRufWNVsNSLKxJkWF63be2uBsaSV2xE4STptU3LQQoCdqCx
6zPfu2l4sby7iitOUYfVScpFMRT+7mYzYFeRJx08CdUFn/cIPciNIu9Sd8X5
QLznsrc0sozxoSR41LsICXWTgm/Na+ZShO/G8uHeBoYygf8qhUM5+J/6uP9P
cmjzZ9OM94CnpwS6CT+Wykj2qRDwzzW+KuMf33RJ2SP/SWgPptGWyEHfca0W
FhuRBpoRlJN6KL6gCIojEj07WZgz1DfsoZl29645wm9NzlUG+YJK7Uhfufmn
8GiuZ7zqpf58wk4jjbstlnl6SVpfxtY5hhc/DRrpMXi4fHbo/NvgW4oTEuP8
upYZDPxquKCJXEzV2Rq6r66WhxGOEpH40eiBltY+x3G2mP04Ndj0n7I2ESRb
wkatSbi+60agZk26fqb7x8Dt5ff+y0VizeOrlnhyZrzLEsR/0VlBdPpam6uW
iEDODCVjfEvxY6EoFIxk+P66MD1urlrhLQWIoc5WRTEirqW3o7DE00MwocF6
NtZDZhkymilan2ohSU/h/523ObMULEyf4mxfxt9REU7UAovr9BmF3fd/kP9Z
g8ipHssT0rPjDsCjvzTfNaAGu3728MdfvwJHirl7o1B6vryu8ol9y+fnr3Yz
+92DU8PY5CSND1tWfFIwnlJLfuVvdsDYWzNNXjia34J1i6xPTGS5kNGSB8NJ
e8C5GhYqrgWqs+O1XdAtmpVaXZcm+zEGsmKDrvT+vpZ0oUbiV/pI6Ct84Wqg
QXHI90TdN2TeXhecJn8p7fPvMljtX7tDuAyaUDHHImuihLtorenE58CN/bEX
Rs2QYtXQ/n5w9+ZbCRso///QBbumk7ITRBuM7FRv/76zO32k8V8zHizSTY1v
obOSqgYZlZHsTqTe6aKBfGnLnQjGsU3b1b/qlo/MNFVfWbrLM6oL7xRcdCPU
Q/MRf2ozx5PZNRQrl8nqtSYZEX7TPCmU9a+iR7BTKtvrGwG+dVwfczxhTFV5
TtpnNI5ZbRfUgdvC+QuB93/3KGr2P/3IHQi/s+TpShOQW4UGy+oWWO7qXEq0
bTqhWthSWEC4zFwNeOgPg4y//czPk/SLCvuHi/vWkqWc5/mPI0OJiJGIMTnJ
wcMSyZC5M9oF+sUu2khZp7NbejmVGaNA8mGstVgfxJrZLbfKenqWNd0895+u
iinxPvBWvl6EB25gmeUUxYaHDenZPjovFfVgO3EtMzYAsfuCIcp+IiLiv4Tl
qTnaEWzc3OWovxy1ddqGRTTSXsM5oTbKJoNXryhgWcQmcnqj2JnpEdhk/Rqf
vJb4c/+W5KGoB7r1EMF0ZdIPSH5dp++bbukUefwzo3/NQ5VmxOUJHO5w+dAG
voINLxn5fkJKahmXRCKZseb+YbuGd0Q5mOLOugE/AWNcjqPtvOxQ1a6OSEBT
+XyG1BPSye6OyZ2U/EaHevqmmHGUA6UHVa4Q1W3FbTFjnf4XTwKba+wHoiSr
chFYp4DJkf5iKz8PvCMQQisq7OL+KPsQcemFjO5ef0gZfCND/fUiBcpXgTt0
1O8RfC4ULs8axiZQga6153z4/6Q0Z1/oVezKVGvEQAQh9lC7idw7SEC9D922
QV7FLWn9QAuW6wqBUKikBz0Lk3WC+bfpVfQPpn6OOGs6BKVNKGWdz0G4q56I
9yXgmyOK2LOhZVoJHgjEGDTdAoTxv2373hxEW/WIfnWLhhjlz08eYCVN/8HG
BwHgrz/WDh1N0dgGyzknPkowlbAlvyOTXvBLKn+vb6qi6jxzPtunsGlSGO+t
FpqRJWs6/gxnmM8x5qSKoInOmENumQdgDklfK/oTZYDRiW0Frr/PRic5X0BB
nvkT8IRCqW6dBU71feO76KVGLgBBik35pKeXArxyLtQue0d/Co2l9gowqLsZ
pfjat1jP6Y/82YvAIcjLYmr9LrZugpUAq3Q7RQHdL3Njvbi1gX7XIW6uZvEF
0EcKTBG5tOEMgOSE1VC8h3XcSw8rWQiUAWUpoDzkQ7kLQl0/nOxfVJsBYzOW
HIuDcolg6JbIkNBrrlGYCN+yksSVxN3vULUlQF5Rb2IiTuomjlQkGm6k1MDo
Xzcgku0Fee8l06ATgCTtIy6TUTfNcTwVL/fYo4U5owty+W/Ivfm0w1w74oj2
5779zGwk80YE3XOgODAF2k5OcBVBXAxi/ZVW/8j9HpH3k/pY/rLm5hRkoVJj
98h6LfAh7kSElAVPLYlVUnbyJ1eyMgDCZ/WWo8jKpQZPTAZ/c4VfmpvGlCXj
h/GdkxPhyYGZYWOm5bGFuNN2mOkqSwyh6aEqx+YGGF8yzz9pBTS8r4CrtQ6J
7vLVWtH04TZKIsBJa3WYmKhsJw1KlZuq2WqNX90r/B+z1w1+9NA7lQw7LMvU
g44RvDUtWou6Q2cXFQTOiy7c90QCaMttBBSreTE1XXT3V07CkxXdWWc4kgg/
VTX4f9uGPyvocDxzpev1PKzo01U3jKBsQiLptR9utwrTvTF7EnKr9UwL+AYL
ShJr7WjM4c72ob4KbAoPwIWpIcGTklp5nS7HifFdS/CWG2QsIDXfCcOxQD3a
9MGWcxcKCabYNXrWqp0tEWR5eqRRy2/Nff9l18COBj9OY2xJsZ4392tIGNSO
GAjsSMvNv4yh+BhFlzfD2L0KBxlqxpKoP0UeUffsyE/kUosl34HaN2K4KfOS
8d/Qk7CrSE0WT2jsLbHgMmFFaLtlnMApnclZYDJMEOUwk5FkkjnZozPvrsj9
7A4BNd3a0Z9ljN/wMnabqiTgFfSRonxo6QGXCKWnq4A/qYH6aPdabye88E7U
ewAexfnJDBrkwGJYYXUELZA7pMREQ8VXFUImb1sGSOjQGWcdaxbe4NdMDTom
zwUKrKxXwrQO2RuokAsPTXg1zhyitQ0qUE0lfK1cgocLEEUP0jS5y1tL0vG5
tQx5tr3dwGkIZ7F8dHONug1mpdZNneFUvrrZeYuZEtQtJSgUGWzRfFCUShOR
4RXn7by5zX3/ThnzAQulTA91YNod4VknUGcYEq+LhBbe1sFU3MC4dZtnDbp0
uL7EDnV9vraOV4dg2dsFvzbOszb3tAS+pmpaLsSj16d1bEaVSYEH9gN7eoBX
IlSYiBRp4WLp5kzynxuYHAUhIaZXrT26fE6sGzKyjbxUmfpjpNUoL9k+H98j
Who5mZnVothE5cSycBZXOGoF2aWaXLAY2345QHb5eZa6/yEPVa2B4zWDM8Lc
LfciUHnHGFKkDJP/f6dbJigxPXT/QjhMNqp1I79kCOaxj6K4FhAyX/YvVsV0
cPW3CHitGHoIMdlGCrxJt5x2/tnMhBKoffGCaNzT4udI9M8GbaRQZ71EQbgC
SkdXzHlrGJ0eDIpmIrrL1T9DmBfmtPd06GZPP2086RkD4QjUT7OxPrfd78TN
5Kz9USJBH0n/rKf6L63mDjZF3wEdMXwPs/JHP8/1mrWpsLJD5FkX/gSnavkt
7vcChwajR1dIoLFP2YUyFQR4Lmh/2ORbISwNg230km86HQqE/p+oYA/9iH1+
ETRx8+tyvvM2qWynym8ym6mf618HrcbYijDQ1P8rbTGm5P8zSVMrlAa6/pFk
H6dPVqRrbQQUK9yHAq99TqY1OWPjJrMpR75CYg1s6rn4diATllqWEcyU+8DO
tljqKqQkEMJzCK6b2AUhu3ClmcOXBtxjFta42+bBn6iU7cOYUPzdXVxdCdNd
DnaXBWylBpPiSop87+NcHtzoJ0iv4+lNiAFjDFKT4O3OOqpdHZmeHNbOhw1f
QK1pZEm3cM6rQ75Lr5yl6e54vwqf2K4diEvagpvWUrh3Vh3tTJPrx1qYHkP1
+a6IlmHLF83mABbL2g5oq8rAPD4eF+RnJZQ+sQwQR6Xaegklmm4aCkLT1Rgj
aE44slPI8BCsldZ89STwuVicmMBj6ghzjmqGj5rtP+0qaAf4aTHLtZ0EiXB+
CLn6vLw6YJYydLkK6xeu8tTMCgbF/WSD3tSQ8NmSV9G5sX0XjGYbim4dJLo+
tKVjF925Bqpt32W5AJCa7nxDhXO53sD+U8DDDBpLCJzkRh4y22tgbcz63Vxx
MDfrnbRhHLQSegCXVJtzzKEoDVha7XmMDfOfQQfgUUUplWcciq18GKwXCC0N
bakD2m9YmCUZ4/9/c8Cphc9uS54L/Qe9FaNhmvvoFZCLe6KQR2yIhMhxu207
IMRoLaGCVOyQ7oWcvl78WxLd4PW7COOJmgQRpLq3XcA3KPDZoPyJNEuNtdSN
epoJWLB+9LbiNi5BTbVc4WHjsL3B1slmDPr+2jl+hKp5jj1ffJ4OtRGs/v5j
oh544wTELJA0IFwIcIgdOBV45VtvIjMQW3C0mGha8PjVqF63RqK/AE1UwESv
p44plubEHiRbrzBQGrzXtKSZUyCPl63AOOVZSfhrYDC3Zx+yii1fR1ftP4qx
XsRIOM8IWFugcfOeGwGgT0DDyOOEj1HMtKmwghRqaoN0VCQlPax55MZNOCyQ
9BQR360h/cfhzBFyiyAwRHKlDl2JpRMzO/Ap+kPmAYkY3sWe3fJsO6z7im/u
+dhh7iHAxvKTVkb+a0CG4oDxilTJ2BgnFAjj2q0k7y//EuEbvZAzIU0tff0U
enQBUVAg47AJOORXzNDnD0rSaQmdP7u4rEnoZhw0ldoOsbNvgb8aaatOh15s
pL5VhrZNtd4oTw1Lbnr0wtzM/nHwbMuovKuRTUmMZaPtHBv5iUOpxYokfIwo
OWHy8sPh5zJAr19TaG4nyyHhXymuyd2AKL2+xLDsdR+8AY4YjemEa2Sm/fAl
j8E56O1WLVxUlpb/jPXwX90H0tUXlSGeoNL6Q3rxjbinJEtb3AY+y2u1Ggkl
sj7oBcHidVZ7TZmlhdIzuLOGerV/Rc7Mbtmal4VYDubz+uEuYyy1F1OMONCV
aFGxcg+Kt9NNV9IiSZUTAIK3o8799JTV+YV2wlWhXaVifUlGGh/5gHF4rA6X
gs1isZtp0VLzOgZxjb2Gi1bzCFBh+U2wZQOdYoDU5njIjcvz5BxVJkX34N93
zKWOfrpnj/KDrESqSUfarub9TOn4xqncxiKdc/3g/J8snAfq4UNfSx8g7ro/
w3kZ8u71HLhHpoPL61+mASQ5qLAME+xTFwcyf81t8vydkt+Jvs80OSi2+lIQ
cZxn4eS5LFN6eqCdC+29Q8Eq15DklqMdcNaGkhpc6vJYFZnKEY7W9blGsJCF
2MIy+y57r2UZyJYJsn0nODpGGic5oSmwVRXlfEH8gU4t9baXDzNmSsLoObno
xZhv5brBp42CB5XXct2YR85ZI8F9w8VWZ3aTLzmQELEt8agyXz1wTooj0xHu
hDrRUfBe/VexiGTjYjnaFdggfthHxJefDGIlBQh0TiEfxzBcs0i+IpmMwSm/
TOTdKbwGn5FrucGSUbxPEBQrbathbpKIQTGAOjx9kZpAeuQESSfTltlvrC3o
Z0uretrKzLo3NFvFsxR2uPHfur6As4fz8kt5YW7Id5PNZ4q07xCXfiazZUgH
DDzcHx22tmUUQCAguOyKPoNi193SrTS40i2tu6amKLyo4yDYfrdlNWUdutaA
LDy0LMn8706K0Er3vLxKJ+SOqsCI/m7aQ1X6bKobyH+VuE8JUcmhkxBGNOzZ
btz6/JMxEm0huiYrO9iKSyRjU2cWXXOLPDRW+uE+mzfK68GstHHWuR8rzRin
2RPcsaeMqCZA83Eaq7Rvl1WTE4t9Vzyxu2Uv5Tp/kaPiFJaFTKwqyjGRWqfp
tQHK7ycqJ7ZV+q8nXwD7EehDVe13s+dA/g29eBweC+gwnivWzhq10M3s4/7h
mYxnYD8TV8dLn/f8gddQ1XLjsBxBLCl47BHf9DFJ4fNEfOkAPvth6P8bKXSB
n++a4fp5kqDyAgOid0sMe2C25Zeff76XXlXQx3RxiUyWwE0PnGso7lsZ9N9S
TuMMHNRpQmhr/WvPaW3lHk5iC+Cu4ynm/H0jaIH7XfbZLm/pNBfzlMYluAup
9jE+opzve8n6ZNl8+s+njqdDE2x6K+FSCpF5QLeiYEU7jjiFtOSQ3D3vvWkl
oM9toeF7UJJVkibCY8/MUSdYxjWAWFMlUgc9yKF4L1TemYCkS1ch9kFl7J9S
T3V353wQ5bgh8mGtq8px5Rn/pyYU6EQsOdYle6O3S0lL4mXyUMxI4x+kZ/VN
4vMweCJzbFE5mZn1SDHkGSq0YElFQOxW0BEphuYaJCoqZXezXBv2l4IzaMmV
WB9Fu4JFwmXN9jwSiNhwMBm7Mc1O/+pJLOnddMxV1pfTEBgTSH0Xxdws+nPI
tdl/2crMNrxAlcwm+n0gcs1RAHP0RvcMgZ6AEXQ+U4vljc+90KUWy+I3vnGH
3I0RRZd998zhKWHZD10ZQ7gWzgIEztltmh61egn+mrs4YhZpmVSU6NEVX8r3
r0obdKkUWH1XuYTb6Akal4/k9onIRBgKIQD6IZhcrTeMV+pmPYBYrlpn38MA
fMYJ1OVcRMwGEyBuRVNHEGB4WXwMa/ndsRpAL3c8M04DunJ9E71JJT8BwXdD
4aLRyTaOvUu0wMcN+nx6uteXM6GZw8sfF2Tei1ucuyVeBFzU43pOYN4p8KFg
dLSasUT3pOfUSDgfKBWYcUDWcD3iuN6gpk76sR5Z08m5zj20pwCnf0HpTxya
uDwIAKhPZbzePHJ9ej2wL5nKzkpDPX00EGTcIH98D/NWo2OklnyT54ojthVG
R0UlPmuPDKvqGn5eSH5zm6B0s5ziCabIEW5hN80ZIJCLtF5+yQR0L5k19e+e
Llk06NFV5k2D02jpRoKb/IQhAyOfFw16ecWxEPB1DN4qTRuFo3DgLXuM/xvX
bBdLUvzKDeMMaiVHgTMZ1ZklCtuBeuJdCs2+VYkh4sGm+YJMcn4Inv4r8QIl
N/74G41vbtyHYkby/iYlGgu3NcL2NYTMk3ceyOhjw/E7Rofj3p4F1pkMxz5X
GX0YJXWJGp0rDOUKiy5uMLw7U7lka01qSDTF99Dh6z2nprA6x2BdQ8axwhZc
AOe4HLL3BUoQKQ+R7yg2wUXmas6Nv1vno9GsUN1SoWoJhhcC+Kdc9TLXAuOQ
o1KyS/8aBQ1Lji6zoa9KNoTyXz2wgWjlBc7gL8RxmUGQTIzQKAT6LysIflUe
n8euKFAjcBUb86s+a1l7B3KKotjPNxk/EI45HyV3s45o5+S0Ze2IK9OVGQ8I
1Kl3fMXfpqi3lTf7s/hqMR7DdRF6z0Iz3uyPJBU8pTK9UlbY9bxmCSGt6GV2
Oc8MvJx+lMtOKHjIzgn4ER30Ea3j5+gF1hfVeLspRi1fb4muk9TQaODSieiQ
STtnnI76WjACSJGV5JMStLUOw5DDFMBtr8YMBF4FKGM8Ez94TklxYAizhMTf
hNwZbRe3XUOlpo9Ai/rpK+7Dkqbq8iN3KPDKmnZvaiHn+wgJT+lk01dNvaGo
QOFQQmIXRpdbXDWF17VWPBn+nZztlwNsv8fHKbZUM9fQJl5lV+qcNi9+b8AN
N/EMXuV8/fTEXjjTLY++M6VPQ7Wfwh+Zi45NR1S3hw2zw05vHgS63YqU5qpS
1bfhp+RH1K8lEphKw6OH6yNtvvUUhMTtGkyMTXt1/b9ZyWj2ZSDijCG97Tox
WirwE6CCfXrSj5cFpFlcnalkPoT/TsiyFOYISF0psIbbbqiSlz47GrLh1X4X
XGF+E4vYsP+5Opq65qUVJRvXTLrhvSvQ5z5u0WcnPrqhGDzZ8fton69w/S5/
lYqp2oN2F+kXAo0EZwPABftJspcvHXFGHlRjE+3sDv2OZlIggz19TzR4xV9u
0dB9zUJFCedCPklDIgxcPhPO9cmpo6UjlKNgxN5WoFtvcQOBOLrV47O6ZlHL
tbZ6SSibERCabCg06l2hWq92K3J5K3Yl+A6QY4/nPnthZ+3FbYfTwSp44NUf
uX4rxxvsvQ55HM/uJ7ihPzJBoRoWwqQe1zK5/R4pOirXhGs1znZHCc1WGAe0
r0WHrw6D/CtKB25k9fbOVdFPsmEvp9qs7JqK0O4GYHz1QL2dq+sfT1XEfWWg
vTqVwLBrxUCCVPy6er12a6ZJaPzg8nP23l1WCfjFV6OWmHx41SEkoZPdL8Va
lCdp2vG0/XOLf8uwQnvWTsnwQcHjQo1wqBHzh1I2XO/2l1HYDou4K/TIuVr/
2+k0bnE0Q2sNGAVIEEh974TIe0Du815Wc6N0eL8BWIEN3i0v3aM0/qBQ0Oa7
GXqTMAKa5WNqhYrXa6YW+mSggOuXNRqX5b9rOyZ64/w2u8csKp9EU//XZlim
TD81rhNEZ/0UaE1xmK7W1rSYR5nf7NiBeKgMAC0ZNfkWnJsPg3V+1lU8fsEl
YDgtrixGW89QVT88rP13YU/n4U/DX1PpkwZ3IcPlbFYGARD3/IOeZ68a7lqe
0A6qvE/Po30hmOiNX+Lm+6k8oGz9mzJ4qAqq3TQn8MOpjV7qzb6ZkNtPCn0O
2mkUSgkUQM6fYYXOkp+nc1xTws99NKJBq5cKqX1486WlHu/h8veL88PFm+UX
M8JoYECZxPt8FfpLImEmaEhkF/gOC0i7gLDlPmej9phA8kfq7KCMs0RW27rp
ziimxroSd/ZR5GEpluFQ5ONRvTbBF/dz2d8/GP1SBT9/hvfhp189ShyTQINV
dpDufbNwPKmFKd8RwtogebxrsA8OXUKFEa5nm2ifkTJx590LurCW+HSotccx
rNk55oFPbOC3YW6c1TgJwmMAjJLgxgix8wG5AJy8LkryIOugXtYawHV6zE6x
GMF8cIckdLJD3smgCZeKhMBqf0ARGaxp/Iwkn8unZmd5aCCzPmrqKxtkMsGa
knWMuT2oCn+HTqPgPFwISct/XrTQall8iMY9NgAoXTbSGIFKQQli3REFzk0K
16YHm4ZR1UR1kFLph38Qm0/MxxPIWJsNZlDsIVNcJJK9uUlF7FuP1cSl8RcB
o3BQnAd0n7hzTik4SfTehxCDhwc8Vzx5UTbABV/BNo2Ev71t4zmoIXVBCzRT
GYkcKRZ+0U3HPfDx5nb0D5FepyaJs/xPjGK3SLkg8Yc4yhVE/rIq45M5OauS
2FSvM+Rzk7BXryWhZgXY0x+0ey9BCN9IG4YXOxDWqB9APHzElzPphgGCtLnN
WtBbYqZ41PPYRjubY8a1ZSh9ceIm63c/KOaPzQRK/ZmXwREf4maBF6MrWyrJ
XcnnUtrlJNcb2HYa3gluqy+UWe466Wl79hInWiCd0ktvC5ECsgMbRzgjNr87
M27IX3RGbAbboHJzsST47DX56FKtu2wLi5SPy476f1X3GL8k9bpdpGtiQ608
F6jiNk3MP6kwPgsxUzyh0lMnrfdfJUOeqauV8FBA+rHCIY61IsN9T0jCLjRc
85fmrzN89Xaf5fstKl9T/o3iWr97QL0Sis9rJRLPK/32iRDTy+CBxT2zUwqF
H6jCRPE7WS8NrKSXimr6hmX49juOoV/e2zo6h5lhi9SxaJkWGgO60pZpbMRg
CYrAmWi03jjO3yTVrGi6XyipdT1VEZbQ+vSirQkbnLv79Y2ih8BI/rSQyLij
ZdXjPJTKETWyPDXR3ITNKXpmrEkl27WtUv18IRojjmqozIR4/denLFJoSh0K
eDbwZTVrcY1kbPR+9yZQ+Ebcw05qHYkWPyDlYSUbsPf9pyBYByWxukxzG78S
7smL1IHjBbWQkIpGHjyrHUiN3YlP+724GpfJPJ0+BWWwjho2XILawKSoT4gW
hMRPblPZ0bIFztpTDrBsytSFbY5yL5xyiuu4wdRM/LeMHs/Mg7+GgSCkBBOM
Cf0i99mcW4PK0Y3sGEq4T6CgRMBKnjXnIDHq5Khj7l/C3D0nrnLaX1ceYyQO
JfGU50iop2y3UxC04lI24bXwAD4LJi9F4/9jhVVrG4Z7Qznv4L777KrvdwyC
ImAl0q3zzQYDvHxH34diPy9q3uvHa1sxVrTHWpzNz3I4zHA0u6zElAnN28O3
spf/Tf0GxSgknYPVwamzR7APM5EoEta1UMgxMBraqspUDlLcL4U8o1eajs0e
+IAsBWHJP73wRwzN0c99ij+yFEotR2LuYiwKEzA5ik0ZbaLWik+4pg11Gw1b
AiBlEmMlkbkBFyWSnxgMbismhZStBhrd7g+rKDcfMOhbuSCbJCUqeuj+LJ+l
QKsclQKOv+GMRrh/SyhNIVnQNPzOjCJZ6lyV2oRYlvTJE+FLN5iPTDpzICmB
NkVPi8XUGYhJCvvZZl/b2rKwxe3l5469iDdIAIr0RQD94rJwYlczBRoZcQSY
2LLb7xjAtw/RcMyaMdavt9/8Qe/EnC+D2foQjHSLaGtLdBKQZGhPm+I1tbCe
Nx/efHrNIiZtzaAUTNxmuEihxH7sR5k1womQM4n/3fD7s0Il8VegKWH5GEfu
x1JC5oN+sjueK4tf6GN1nXONkeybRYkHdrUS5G/EyKib6/hLIEUAVUnx1SA4
ApSgYdLnyJTDprJsfusoO3uHFOQNqhEYhs914Fty6/dRqukLKGfvlAKFXOEP
jG57vcqD95+3xoaVflYfZ3J8yV8fkO6/o6t/xgAiUBnp0MXqwGCPp2Jw/y0i
uB7bnNDZWxVx7HNbkAiJH3rlRX/yhgUZnXdijE/s1YyutdwtIdhFnYCtSIje
l9PCy/E2Rz5cne/J+u425kJXXNGQVMjPpalLSfgS70Zdjf7oqe7MLv2ZK5rA
Wvivc0AfBS/wrM9EGK8+cNe2Qw/Y/+0Ltqw8GYgvNxXJqPZGSx2vk2lZFB/2
TKOPJzcafzCK0qf4HhK24GBRbyI9taLborl11hlDLOpXA3jPoSWpzGHd0tZ9
NSZlfsj7RMMOrZZ2WCLZpR29jMMBmy5XTFyh2ChVS618nH8AjAp/TgbIjtDs
WNyXkiF9kQQkjQsDC0n4MQJWxtE451q2kb6Y1auRpUajlRq9KTcFzp0j/FpM
jCGuQMNRtGDMMa/ZKr3qpKT2M4qIK/LvRfFOIMjqFFuVwXy1+1+XiwJBMRpB
J94zg5Vp6Ujj48sW7eiK4PKKPfx4adkzH9IHMZiPEM0jpo+aEKiSh+oikju2
yQwlrlCgxOXMYlCgrfLyTZxnGA8SbgqxPZznOG180/MYEDQjYSSu7L5Vmh31
VozauG12Y6V5gKqnIYmFgbFpYIjZ0TATztv+c3W++Tf4i+MrDQaw7mrEdPsE
PNLJG3cSM7dtsupDZNOaI7QELddSqMVfLR50LOTxqkoUs+LFvR17ezVDNOuY
s8OA2T0DEVN4eriJb2F7kCR8ChBiKZF6Y3OaP7QOJmuZD8xrzbL5wv3yteFe
C87P/mKKVLoDVeg0YYObF6cLLv95YZDCTnvuO+OYsD2uyjWdeLjyxLNVzQR/
edbobg3m/nULGjbWPCyIy4p1DrXxKdXA8BZ1PD3R2RSBBKzd8+JefskIHn7j
unEtGCtS8jk7y03nwgX5qHhaGzWRzEjmD44mLeETS11liqjonMQWlZKNcYFl
TDSKVg+g9pcngNDt8kSm8ORFaeUTWFUybr4OCcE2S9I7WtkbAT9Xhfuj8E1c
tzHzjDt3uTsJ560XI210cwRSP9cS9NGiRACkLtA4biPm9YjoVJzq7oKhnbjS
WtrJHMOygB+eG1dIEezDovbyBpp1RjpUKjmt87qHXdCsVtA9ER5UBDE0eY5p
tNmBuGFgTJ/pnkoYJumEOJVh4OV/4BoClhaoe4klNn6kIcjH5wo6cZCpdSfd
fz0j9t5LWnQqh5aRE+pkgeu5zVR6erqfb50oTr7uWOPXgxY9bK7WGrg81myT
+fiBtIKnqi/2YKjBmgBiN0tVUaEpMO4Nzs8Wckf78f/klgVn9FCR7uU7yMTI
SPTr1eWbuJn93eMjhxirB1c/4cx4AZEy56M/X4qcy7hFCqRPZHJtpqv4eHvC
wml9ZW2N5KUzwPeLrvdbPqMFSItLT1ankOFzqygexA80a0hDdo6XaPg9w0t6
eebV8PHhQO1ot6kortV5Yl+P9amYzjb+tCN4yaXwJSnzj4kgMbuedVe+uAsu
5bE/lIdS/UqKjmWvFXgs5KRGOCY75JsWnN0sQt5MtYg1eLTOdtQhwG9rmhqK
WKecPUpk0Y1gpUthkb9TLFmAuII9lW1fIjxI9Z59iReK/IX4Mbza49K31mdb
Bw315RjUqk788/TOimxi9Uw8voIf3VP/eZImlXDYXbM2CMIIjEZ1iZEJbND5
CmKop2YM/P4upV2jyGfxrQQF7RBQb4iSJKWwZRiLdFdrXpGmQAfiWaTk8Na2
UsZIjrmjRK5RVRMWdmcbFfKR1U/qpXXLZ5hfJ80R7zprAy9uxK6ps6Jor3Ld
COIn0JCb/LqG6dRSMxiKC+gIBq42M8xO3IrQ76gp5lJePJQQ+FFSQgCSgAEG
t/+iUWnPlVyVIozcI+BluBOhpMC4xS4FrYGqJOM0MWVBpBvLOkqtSXKC16Q5
nOBqSY+eu7xrjGM7+n0O1Au1baMFH6F+yxIRlrXyHicrj6Ax6nAsWd+USiXg
2LVwD6tSJXGxkaXlZybxBh/oxfNaf4vx0SjYcK59RvTnScspJ+6tRI3SDRen
8p6mJEcznrhp+sGTB/1fdsISXtJygMIUHKmLE1MP3UZWET3tdbp5X3A7lDgh
juLT5MZP6czQI5IfMgqo5gYW9BDq/uSvOlA9/6WQSCfmdeM11iR8YV0sokGx
uALfS7vbacwc16nhLHtATilRQXjehC30kqjmtrxXzSVKeHAPIp4aqmeq8d2s
1zpjBZA7dU1RDQwmFQU3Pyj05ecF3DmR1hsAqp5Vul1DSMIPP3EkXWf8pObl
m30J48OacEVfz+VIkwfr/IWFxfzJVVRONSsQFOheXYeCOF2nqLVeHEHJqdQP
ygutkyUJJSMdV47CJM7cYSJSWdntfwYPuNNHKKByFoxVdnPR3cvsYMlrMvk5
Lg4bGRJTVDViuitMXiRoPoM85ce/16tYloRHCSEnansNDlhJcM0aYlyXrNMK
aq7n0ZtZgJ1XfK+AAKlZ6xHrXpwL/L+33IcA1KzJ0JfwhJsNIYACUX5rvjiB
1iixA7+QhI8fymxUx4bL+ixE/sNCH58Ep/a+Sd2OUF6DJ33+lsAdVh0AnUiR
beXzNCvPORbyi2bwbQe/GiL/UbW8ja0Dh8S2ZyQEWFl2jPcMAnrrHrFRmsrS
k0rypfmczjhpOg/cJNPKw8BKsZ34mEtaoSbIEmXHx0NVz3rGX4Z6NtGWcmo4
2IWZ7wlFmKEmb86XjdySXRuU3CG7KgtjjsuL4xMCFYv1stv0XaKidtGez7eG
4I48BZNpN8GVzR0cw1vj6dIdZX566AHGmUf0YhZTSXEML6uhi3zfLnqKIfce
P+mtqP/ZQRiass3oLebBR1uE8+LwDLQFJqa3JfbFBkT8tp1n0/T2YuFMQS1h
pOMxyvhdB+ZjSmQajKAIaeeFEYdXLntvR8ZXht4jWMgd/cFhkKklJlmjAlbB
owK32YLQ0WkwOSfi/KYnR8LRB4J3/4rPO0phUfWmPGMt0oWt18LgIgRSbeHV
aY2Gt885N966quQTWeFvP+mGMZtrBf4tRdtrikrs3uhEDkLQLINqG/em7DdP
9IHVY29/SSRUMrBT6ZQ4MYItepfXR+7/paqdrtv3WM0suyeDeB9qMFMHUNmT
LDO+brtmbrKTIAWe7NyyDeUzBICL7NPC6nUbl4MDKuS+9IgW2rBTq8CEGvbX
sqzS1nI8XwdYrSBTwLZ3xrEn96rwPIJWXm3jnkhgVEtEnJnSI+dsK1P1Pxzq
MRZKU1n6X92RD3vbdbj1oGOAGOaPBNlhev5wgb5ln+Kde+4b2oTHGw7epzkW
cVLI2Uj5lHZupzx5+T6Jqp1y+WdhDFxrl7RwnKY0c21KCAQMDE6NL3CUINwO
Sc0Sk8W5REYUHhakJJ9xLwsMTcNOl0PwqdMqcq0RSWDINGYoJXbVgLXrND7e
dIsQF2HeqKIgHy/9aVvuxpnu6qRT8j+xYfmEVrMlorrLaUhceA+sdDC4jZyn
B5f703u8K7iRPBvFUxZ4T6xNCjn26gGB2Kv43UjrrN2FG4JUwELJvet9+qVL
jSjN4zTclTmzGcKPDLULoGeZP61XexztuR45LIOCx0dqOKtKDVm5O6Fxb8uC
xhwVjW6bcUjoMale36DVB7imm9eUlbUD7iR8A3Ym/kp0dXt9SNfFX0W6Sdv6
KgerXX1RY6OILBF1WX9lq9JgG9rNIqbRnn5o+6ClKjkezzZkBMjZQUApAor4
HyFzoUoBldapEZetmnIqMEWjNE3nxgBpT6URhicBIjSflPtli/SH6NAlucqK
w3wH4uhE06ol0P929e6BiVVN4Hz+djd4vAFxYZkg1fn6zikxOKYFMFDDmtHM
tPwB7xp0V7J0+QtKGfHvHRHDOMcHDIi/8RazFWmRb0/Ae88sdy80cqmP4wD+
KNexB49Tq/zmluO1BTatcEGxFiXjERwKce8AZPjGeUJOakJ0vTOA+arVy1cq
9YlWDeozZ+UN8SJrPy04mAibDFJDSO23/N8N9VA3UZ9jnkF8avHhuLSTLQYi
pqhvi1in3Jmqc6bmi1A6ahzxyGL3UqAtqpvcLOQ0VcUqyWXmpSx7wAxzMS8K
oTskOMVHiNLHv/OxGiysB3AK6k4xw8qAeH0lLLZPtnFNqYKIUcDDL3M4XKcL
awv12q1svD9Q7MDkffbQnu4df3ycNU1XDdUtzkjOqV6fMtjyegiRQAORSqVn
nvJwumIAn6dlnHpo5R/jhiOJXlI9wFNFBcj530q24a6WSoKOWsMoZh3mdRRB
b0GQZGaj7o1mi+b+ubwekYEr1m7hwgXPrJwRiV/mvAAI1fONzgI5BQi4sn4o
VAutrCScpCLIYetax4WIRzRg4O6t21TE5BNa4zGhQHXGKIFlZidI7XoixBa0
gaQL2ECzRckDZNDCzWrpEfBmcwXXeRQ00PMJlEf0TlLHWlPEBWrCDeaSy1wW
MF1vAb+/iycZea+e1JPBisKxtP1b4kktsWk0u+6WKQjlkcz5UrooMrYoIFZD
49TNO6KKbkJ9DKhkEWYOX9yfJCwwei5DYE2EoPGnsnTAhLJs+ilVWxtTaxCA
NHmXn0H7wj6R0KQu4J9QEd1Lrk1HmqkAIe3hiXbz1r7E9Hr/379i+6fvnXVp
D0A6rsZ3upWgAPkN9SULu2ZQ1M82AEeVFgn3PGbIo0jhc5//jLORRxzec085
G0DMVG5Dw/ChNbFAaA477doEzFT0tF601KdkdJRp8+0CLRnIHXxlzAtANiX9
ngxS+krTP/eEQcrKbhIgiTtwi7Wmkr7EYVICuuOQM+iCqJTgner8RnnJOryj
/ibYHywumDmfy5vQQMDnyV3ce7Mg9PZN4Va5F+eDUp7LJPRtIxIAq5WRJNAZ
RsDYEDqWmijbQFHAXcDIKV0KRMR19w1M2oGJWsQugpglDr5xa/W5MmRUNGXZ
Zf3hLiOO7cGgEJdckUFQHbOOoiqQKoZnOs/lN3UyCheFq6UUeC/jHZ9defqC
Roegh40qge2SOcANBFLiKuyOEou3bOxVcZRnTA5kJlhL2ToLWMOjTbUC43ps
9ShfV3yxTnYxpqckNWj33o5DaG22kkuAzQJOiYcezQaSjYMMfmkN0Dcd+G3O
2mXRS7CdajCDh7fO0HyRxNVv3FSO4FDxZNoEA3s/RY4lgAiwiUaI7/zXOcRg
RMw9nv6SjHFWUsID1DySPhsiwbMOU0E0ldH3OhtInCusv4TCHCBhSv3F3nuS
UjsczBYNCcwdcx4+GNpG7t8MCE20NtleI6Ea7pYNYFJx4HPRRzkwQ2SxYRWo
QMjWAXycJ59I7wB2xTDRSPRF0HgZhNmUD2ffQ+sTF0hYghzAC385rMc5l+Gu
I5youobyA+VNmkBLGsD+And1UAwI9uSKHGmHqL579ryNL1g5iuWdjGUpb1Dz
Cg1gPdgaMkm5AhxK6W2CHTGQ7mXsHbO/driKOvhUGDttKO2vK2rVMu/M6LX4
MJLpxDBQhI6XHPTFOcx2RBzFkWscJMvtMXToFlhMbo5NROxtlw+tOvjXOnRZ
Ln9MgnUNEkyIwgTOYU8/eu5jg1lOWzcQ4mzIgaRD93ZVq4XV7PZMR0EMLFpC
kW0evWDfrWd3fx+PO6nRQ+MvEuLnI9y03YfnBd/XwNg2vp/Xwd5KTS/5YVPc
M2iwP17nFv+KHaBUAjArQ3/f864M+Dj0IUXpuUKKyZ4bxbBCV6vj2ZAwxRQT
ziYPRQIR/4eo/8HElfyyAcCYWhiuYby744Atrf0rrDy+JBgLT30rbDCY7W0X
VkT1GZEDmUzbdh/wR0Wsud4oiqCkCWom8AtGu3NKU7BA0vKVdmQ26uIKEMwl
B6tg774fIvGx1UvJxqNCvwACw+jBlPzvg9WX9T6tgAmOERsLPMZ80jPnL0Or
QNzYJp7IoG+Uld1RKKpoRUteUfhPaY7GI9Kzc0nwUGLs+TVj3ONX1vHZjTNU
8CMFjcQS8N1Xp194pzm0/hBNBDNw8Gfz5EAScLaf9PEj50F8aB5STwMmaZp1
G8H2xWjJdZWJd8/JtcjIT4iVQHiGgIRpGM92L5cdeNk0an3wbau8zAkvIk4Y
q+L2eLBoRe/Q60RhEnRdr4BHZ9u1bf7Oi9RxtYVrGIaVqAHD0R4kh/rq0Zkk
3Qy4czbZvrRb7IPR3WDFhy6KzeuvPK69HRcJI3/BDOZljju+wuD5RjvJrG3x
80gUXhBopTlzeQ1bzUwGjp4R7WsSZhdw2FEj2YhYolY0MN5fvdyx6+7iOgkS
PAZOYCMnLsrDC1uzf8jb0vdrLKsoq9ZyHkT4UU6MZIe2tT4zGtGg5GBRYVAZ
04m0Qa4LmJbqkAHanoj89y16LrbqrzupJbDZopVcSbaJ87oNuT0yxdpL+eCs
G8vpXsno3xAf6WPgKuRZ5nY4FPHjMw/XPADSOOtnni62P5FkdTJ7reFLMM0A
nuYMahcLkCTBoWDeF3ayqMGwC+jElOspWP4xQZ1i6n0bMBc5s+9s+RtLOt0v
WyoikQg/G/U5Ub+StPvpq1EL09kxQ7wwnRMUy3AFNoA+G5Igbcg13xlnFiaM
swkcEcJrJaCNCcPldba4n5XjV4nnxAJQVar1p76B9zS05JZKj+vB9jhjypxO
AHVXT9w7UWWaTLn/5NNV6cpRgXCfe8dz5TwZea5YlfbnSVeq8ykJb8b7Il+h
mdeg4EiRvzU5ktHr3jtoPkLRwP+wMbBRtIQOLfxcHWy2f0rJuhUurTJZ0bHb
Jwk5fW/C9plVa9DlE6zG1mFEx7SPvbSG6Anj83BL1UBXX0hmHNCCh7wT5xqy
XEdy8nrLQ1UT1xHTQRJ/eikFpRfrANTUGd+V5bDXbY+NZkEcrkPxEyNuinNj
a4y089gheS7jC0b6P7C/y18qdYbcGiu8bphShUqtOenqN65GZVnuqcsmJ6bg
+/wnC3GZqoB0aq+mty2Qd+14rsd3vL25Cbo2uPNAxUbCDUm5HNIsUszM7t9x
7glygkByprW3d0CCEkWPQ+TjeRx2nXqcZnL9OUwCoiNgJJ9uN57Lxu6Sz2Pb
wopyLedCYY1xoGHaySYopyfOyR2HtAH/zNYe5SxEIfGmQz2pErtDHyZ7i0RK
S7HEef01RD/K/fm/aOQzMqwLWUN+2LNuhgwW3wH9cS9O/n4KBBn4CJHcMmhA
O/ctwJL+q/MQPDCLiF44ZCo8MBWw3rFT+MM+dVVomnjFrXjJwxjTCrWitHlw
vm1AEjChfB2j3JIpcDdMkT9QO8nzfnsl5XL7io2RjAsjqBKBW7he73BSntAa
R0V6My6NF9YoaEbpKPNXL1mB/krL9ZkcyJiNuDnns2uFBI4Mls8aUW0qX1oK
QTe+F3KZw3EeSdptTMlD0fvsdo4dTuEP/EWegl/Xrbf5LFyFDiZIV9vMzEZ9
1CVNnMrhWMKbPBaUQMXtfDkGXstlNRBt8nNJdVpuey+r9/Ctt/qH7RVV2lnl
jgnX8edLDQAytxd6bY5uY0so7w9V5VruKkIOiwE0/FX6IQaVlruRvKgKOBDK
q7bVKiVZGKr5K3qppm06ARCCImSOVGcMaVLfwp7t48gmXDeg80ISn2E/dxls
Y0jutDxFTmvOsOUnZ5jN8FxI0VPzlxzPtrs3QQx7WybrbApME1fWvRo0Agzr
GGkMCt4E+0CRAQPMZXCGIClek8FA28vlrK5a+rulXawEZFXParO0oWan/mvx
BSAFFPG0F/GuYUfVdsdz0b0uf7WCekj73Ut08/XMcwkJG5LKKdR4kPCZEuIB
995qAtBq04OmVfX5Qk/08Xk/Eb6VMDAeBiVvxblHiqXwfXNO46aESrRBLc8G
R3XyTFSm+Y2bythU3wlGr0Drorux1XERzDnyVGVpuxs4X9sSeqAndHKaJDB5
kg/sgBANuiy86cJWMpDhXOGm7d/V8Xn/Yorlsy3snPo1DJt+HuJikb7TRojC
zFYowPSJMjShIZ+5DPAHW8bYtQ1NX+CbsyLNHjie1OEg6K0ogVGm7hlZOhU7
6DlO8bUPvp3wdG3slqpvfXMQOs4DMsdSsLQOVM3SvwZmNPvnv2ltSLfE29bH
OreqfY/TSl/SAoQvR7a4PHRouZhXaPniSolIAas9kn2qkhoMTltk/awDnHpx
DrG0nfxHa3N50r4ftlhdi0Efbh4NgrmpQWaZ7p77MRbAjQDiRKNptDT4S5NQ
HKZ2itr20wZ+NQY45y+Tq/ZbaeKJ86glDAFAbg0G675OMr6do3+TyoTyrKR9
scMaknXv1XiwfVCEWqax+GQiZGWvkdZ58LiBeoethMCz7L3uM5MAg5+LAgV0
2fb33/2W+jFBtGpV18/onyvj3PnJs119eHzMNjxyLg8hHFx6GkNd1AfewZgl
55waid3gzeso61MDOGR5A/kiUFZnFJmksalIdC4V8YgwVFsFXJIDU96cDTyQ
Y2QR4S2j+M59UnYR8ZE064GESXozRnd2xUH0evQSP6NwB4F5zMqCay4/EWlH
D9ROeOVuP0Qx3a30v5+9SqU4M7m+VM1+/6IpQfmxC2vqCLUhD92EewFBGdBG
z9lPy+6SOIqApWvcwwv1Nvf3CK5O2GUW/+N68MY3efp47Wr0OG/fQLsd6wh/
FOf7N0UmCg3s1ocsLMadkfde3fCtGSR88NtNXYmRYIh8H7JpAoImQSnqAFX+
wpkaYUnAYVBQHFv4mD34HPgYg0q2+yeidjSLgQ+OAzhHbEoxxHgE4HUDE2wc
jQnGAZc/lk9g46rytrqq6HIKQkRSbrhOooi4FN0jQQleSicsqVNxuSqIfVvq
bqvJpdieAgIMM5/pEfUjyr8neBto4Ar2CaMOWkfylwuPKMizcDW/4O6VzQms
hQ/AJ3do+Q4zU+9owHEoaVjBV57PbOzKgVcYfG7NkltICnigdiOI9qo0erd3
aiHFGZQ1RDQ2Ra30dZdIv7sF+p0O7b/hZHD6mI5Zz+d6lQqC9j0ztTDBl52b
6dtgcDnogzo+rEe70eYXDiXx3Oc25zvJ+DD96kuKFS0flQVKhkvJbJpv9k3M
Z+GA58MP0X1Xw+hl2NG1r7d987jlN6li7SBQ1h3y/FwtCGnW3QQrlmLtESLJ
76uX3EeRI0tEmqc2CMiQifBA45rWGGTdgzoF/Qf3BEv4FXIkAwsbTiKI2gxP
JFrG6elCLKJCrJPXLSmgt3kSG3oDbA+8104kpqsK+buuMACCp91G1h+Do8cn
n3/NvOqDD0grXHBNkVeep0NWjlY1P4zWJYBfbGe1HvmaoThJrFlxa7LlxWJ7
/412t/ygkqYINM6bLrfsRju+U0NEpZLFVnMXVUa/SUmZkUb4jHMqSrMHIoZi
rEAbb5HaFC0qO/xciPHswXex8gcdkP77X4gcoqXHMjsvgllgi2rz6RBJkwFm
Jx2WyJSLpFxSE6X4dPZjIumjcyRsUCTX2gIaukgpp00lzHnHLKCQzp+7sf/k
u832dCmFehj7VoSik04ZuHBEXSlthFYyHM3xloF6bCTYfGo4KhDX2Bbh7JsC
+XGBu14R2jcOMC65+v6pK/izqL7ieUXb77UuzywSJXpTdyZeV2y0cdG3SHqc
cUERXJF8McypPHuqyGEkB5ChBusT5er0PLTtkkxosTwCziNqLCUATJwIogx0
3cZonvd1M/RQmJLm3+dBfR+XtzHC6NXl1eylxQQAAzcAyReRsZb2tqI4NAnh
vALAM5sVU/6vJRwoaex4GPsk+2HiCmDvWKU5ivLM9ioOWUefLZTvnIdcsJDY
iD2u/GBc7xAlu2ugl1Wyd+zOHD14AlSCK8TImE0Yhrdu6n+afZxNh4Na5DWE
GG2KzfyZD/tuKIk27Jah3ukvtVBIax5y71AcumRY+VhVOjXijqhsJKgaCzhy
qsuGxVEdWT4dmk+ZgMUKBJveKrLsXPuTFs8NS0CaBXKF8hm0L94mO2XlqC1a
EQKYaQrQ3RYGsI+HxqHuk1ZXSzNF6oYnkBzn06n3UOT7ohiaG2pvkL342rju
YzUiY/P/LdOFHiCQ4m9UtvCf+9VOTVV40FG58dT2PQqi1ffki/bF2pZHSu6/
K27dSkqynE1FxG6gESUJN1Fe0xxj96otwQbYHGdRi+w3QKSyNUgkQyuk8qop
/GfDAB7n4JWoGJQ9E4aUuNRz7iwt1Pci5QtGq5gXF6rHF6WcishXk4PdVmpf
GMU1UCGm+1Ui6EOrCyI/bfSz9opLtHbWsNAg0n7m0hi5ypqGD6/ya11r8zYh
vldb/BqBxn32UrUvGfHPYWCL+G5rcBiRT8pNxWiODKevHfqYqKW2ri8cyBfV
NDXQDQezcCApUQM7/xS8wecuuNm28B9mZPYd1qzuABag8T/H9AIs/nCyaA4t
ifsyAm4o3X0dimTskM1lC5tlavhSQh6TKixol8Z3ZjFo/YSf7D70/bbdJMkw
eV3HZsn60MFJzGdAFJ9bM8RTzM8rTAhqYml2HHEktrP+jLip3NJWdFSLPftr
RTDgAhpL3+gMBiAUoh+ntd0D0T6UMMMCV1i71uMlfUhqocRfU6SSB2+5VYq7
3SIusc9wCGYuT5SU7rU08WDMZC0AQp8hM2MS33rP1L3YdBIWSIDX4AXt3LZ+
X8oJxFBZKJLhxHRAJOO/7x8Esrjm4wuungRdU5vOktX/gv7SBlWkeC2BKEiG
gtU+87cTUvPDhNXUga10oitl7Qn8s++vU4gr8v1RNQ1QoTRqGQ6JHFm3+3px
/7kFbbPHV0bqEOpYNfxw8KNjQUjw3vXAKZH+OurJuUao0JJtvjjU1iKTVy3J
ZQNlpulhdifBdMU1SdcxRwvJtXmmmhphK7W3KDJ/V815iNtyMopz+S0q5a0W
dSizaTQBZKVzvUvfhJK9EIqAWcUolpb/giS9UQaohO1m5xBcIbV4JGkKqVjN
zaQjFr7C0MuNCSuU0m6cwiGN4xmBWrdguJdLeAwuFV+X9HNwpgJrcfwc7/Z9
ajXK75zZ3RzDeRiJbmdUw5DgW+3BayUXem8Z3nehmUoNZRYaiSvCGlQBZIE2
l7G9K31sTiLkqx3SZtFdp6lgFU7hv3vIxUjRmuauvU1MUfkmsr3EIyOmdtOx
zI1rbVA11uUwtz19M5aeoZoyeUkXQHscDaHAowIpLXNVFKwHLQqJE8ZUibEA
zqaJDalTjppRRDsFGafURm2DbZrgBfzcbDz2UocCaGiLf0MlSUxX/dVB357i
CFYGUNM6MIvXerB3n1HFNc2o5/3TjdE++tetdcUkNwtqkS9FA0QvdAq4Euz1
N4L1GK7gRRk1RIN4JpmLlUtrlTVJaFi0OHut1qxf7KG5sJtELtf70ZWMpH6i
UEGi8cHAcjBkDF76LV3V4z/OAtvApYw3Tc+Ig9x2L9DC/pA5C2HNpeQHrFld
fmYFbbUwk6gO9tJib3pPoFvAY8wgFjjBAFbP2Ip47NOuu1YHBA3wh99dCXz5
/E3pCSX1MzyWH8m6Qol5y65tq3Iib/ZDf42czoOUWP4HeiDQ0n1vUM5L6pwq
Wi4VRFXeYtkVCFBL9pipOoCw7b1WjHSQGXxf+RelDLa3C52P3ts30+x6f/Fc
zo1vS7uKD1mNTRb+MA2KdcG9k6AxfmKqTvHLsmnt0LnZ6V8w4jPQLI0SZ4Wo
wbCwy0cxMuIrHtPg68AhY/2zesZvmi+dTt1KXnyp4+atMU8bZdO/CAW9RYDy
bMR8bpEd4X/jH6f4FUVAHWY0NdjvR+RDZWQK+ekC7PGMX+wceU7NO1cwRwfY
Oee5qKXjtXtMz6+ipUQDEEGP+0cip6Ps26b9mWJaOvNn6d21Lg4qVChxqqRs
6EoiqmDo2Z3H0wdvQgndAOcp5PJgjW1P7Vm0txsGyPhdv3YTSUd3IoXmWD7f
WRsTVqVny5lSFYxyUL0oTK8p2CTzrhDW1kzT9UDD3j0sfWSi9Of2sMdMJ7V+
1wOZiZEtkdzejZU+T86RE84EkgrDWXbsrKr4bThl6wDflDV9FT7ez+A8VQ4b
9Amf5MWUW7JNbhxbtsTes375VEu1mNQxWt62whDVnHscqElH5TKOkJSf5ILz
oazQTllTT9KqmkPdV0SZPnjA6nH6MUgFk0Qs1PT5ObwzEVtUfLNXOcfhUBjv
Edj/dOJpJkuDgugoJ3ia8DjDtMnrLQLLfd4tNARotM/XMaCJoQVM+JIQYgcr
xDSmRac067dD7Qk47j7rb00oUmKAa4N8m0brJ8nqcPsqfVsdvgdnG4OqMSnT
9T26ZycTe90bC0pVcC6jTAgVYRRXVJxkM3n2Z83Ad/MgCDD8cb6MDlhTNGr7
Bqp9BQuZxAh/bhJ1jks1jRu9U5kRSf7tcnhWaHMqfIv6om1YZcAIXwHUvtBi
X5Ys4m+VA/TO6MVoCADN1EZpm2JyTS2RkbOvPi6hFz/jI/U6deYHDOaFnXiX
Xu3J4oeEIM7tVhuf7k0n5CrOKSm25xD8a45GQIgvGiljOQ92LK++/OTzgRiO
dUcBJL3xQBLLrvxzXhppw5JXhZs4y5HxYPX7MXuJyMAqHjqGYbdKQZhLzTl9
bgYedO84DBa4hg6RTp/NZpaoZjUWk7HwyPIf9yUrvGavTxDWhrhAFag7vTei
iYiLCVzXBfE1QCqkyrNSYJm6OoAOsH3Gpcz2Krsx39ATHGkd1tDkyPAAjsiR
3YKs8OiYfGUAJ62FemS1gPtrvXcaP3CeSJW38OHsfCAMY2E9baLkyG/oC6Rs
g0gdatxQdHqn2ul1L31yzDqNHU4RiUj/y1c5mEIVbtUYW++cfwsWRG+MCOA8
+UY2tTtHoS27Q5ffUu6E0kp9SLf7ncFWNvqJbtMBTAIlFh0nJuTNl4JvHEzf
PyGrMGlw/pGf3fay7D0MmJHHGsxAntbMjlars18wJFezO4p6e067LihSYQuO
G8tiDSppirK1mO82gH0RTocjucvT3iXAHHWK7ntYweK7/dHXh0Psgokl2G58
TTpxnpTGfObueykKN6zvy5gZKfFozc1l3UKJmRQm4fjk61l1YPTk1IN3RhtJ
IdSIu/bTtLTn/NvkIliU26Pg42pR98ycB0utymZcko6XYaAMsQBBSeUbIHM4
mFxRvVt7GHDD5BYteNzg4POeWcTpX1vxHrbvfVcnS9khUxvy1rHhAL7Cc9Xo
/mynnzoV+2n8yZqtT1f5I6ricPcRFKS9V6leZWiHQkmCeL3AYHpWgRVjHgF5
zy9BKuIIdizjZyPb3+pdjKfXKLJ29SWZz3Utd6krVsRaR8eW2F2zfVmZ4eWo
j/ufjcZsv+u9wvMJH1qKO0PQubI5pg7oCn8noZ9/YJmhpMRQ1mBnbJTy3O2Z
AzpjIVDCe5U0SVoeS6M5ByJclHicdX/EAHfDva7+drOxVZFoBmUblUlhYADc
OnTz6abKE6gH7Qp2VOJikM5YmAhrBveEgLpid1KwsUxXZhMK36/HWygwm6xA
bVgkvYL+vRjZq2wvx4YIuUGBicu5uJCJvVj2IABOf4jtVjt5MTe8qC6MkYgi
pQlnyHXFZPLgUQO8vOCHUgN2F3MrbwRA2RPbxv71wSYjcAxZGgbp0y5UjEQ8
alv6uGHRZewd28bzBsIP5rTc44w3WJq7PmyEv8FXyGZWRICXp8fAgCXfL/KB
A178haT9otqC7u9gZyKKMXr5aXSzldfSZe1pzjezuCip0RRdgpt9QQae13Ru
zK/9RBoc2g6MxvU6Ax/oPg3U5lJDO6lzA3X+XU+8CxTQHP+hCJ/o0hrcbJz5
xx3pJENqMz0rV98BnW1DjjbSS2ZjpngCrfwUgkJ5HxyWK12w9Dqw/n+gnpRX
p3+eYcTgzcGwDbQYingRg5KOGHaigKyisc39iJvGjfWFmWnkjU2dO1FXDp+r
VR1onnIKMvu2ZSqJvfPRR4E/ZL+fdk+QPj00ukpary5W3v4XoAKmGGqkm4N8
C0W7BgQ/HlgVBMuujLFs4reGIZ43VgRGNOAYE5Usn8QO+rq7l7Y//fKsXmw5
kUpGD6OGCDiiOmU26RU1+GArfEofonw4RleKNoTEPS+T7R2qkxWJVR6ubQoy
73jP4iXYeIBdks11qhR0AmYF2s/mZL0dA31dSP1vNA0K9dTyXYqeVRU+mIUb
k/R77A/PEVIXU4s5iJsSUx7q02b4dTpH+Vfl5IhZAqfjWCBpHYsPc1lz79fo
PBgVBcYDK2MjEIpUrytPqX+8fDEmoHrciIR29cXW3DLN/4q9/Vn5k3IAEB8F
pcHMNOmMKvwa7dh68jKI53BRaEKzfeSyU4zoJu3ifdN22HRPemdLEURJ31Dr
AJdNHJPu3U9uhc1x0OyL3ao4xAxdHSr8jsfJzJUfXwn6Hh12bRS/neF1FFip
xkhaRf1bRd+qRuPEMH0sF+XZbM9pQTsRMQDQDYt0/l6VSStQFkzAe/KTYQ8f
VXKTlxzx6vF5FxlP+RzznbQUfqJFgCIyPucaXFyjYXZ1gpMGFMtGOPylk9hv
m0MinwodstaiEHwd95mMcuqx4dcCzuKQlc04kXgpq+gqykTeqM1hE9z5JwSR
Pr7ynfboDvvxv9fW+XsRi/NK86aa+VUa2qlTBFGJrJV3mKlMMHZ6I2gIUqWC
v5dyAaHpz/RmLTNtdMWEdvFlNfA6VpQw23b4NCxmugW4GcYrjdcVoDaBAr+S
7kA+ezolpI/wpqEUnZXZ30VCBwdt0mYPxfqYNWipUuIjAs7gy+W75+2OOYUh
+I/xR0ytzne5+0wiOLa0jtM5dNx0MlTui0mr653g5Y6NjN2vFcEQLRvS8vc4
y7g8LEIpmB7AKMicd6Q/aSLYSzOKuU8VmWRlf1iSRZKZFM3CQJAMyVVXfidn
g//lahpaXKFrlQ+Gwzh419ek8CfPQq5rIo/NOjCHhauiW2cpxzzF1ckrpQ4B
vYRYvV8hid6/eRQLY3CO3I5kEVn3daTd16N/Qa0n6mtt1t0qUbTseLTFhJCD
YZwCw+MqVW+GMoqJK/tSg9ewBM3RPS0lJtzN4b6YV6DBKxldCjQhqDRMQ304
Zw1UYCwe3xqeEcKWHCBgKA4KwU2UA0RHZ06W7GuyR4tCHTNqHBohn5Tl42Hu
DXp0VN6I2tGg1VggZb+qb1ejYfGda9xg71cp5N5fUxfihpcV+75ycRT72kWz
GzvV9NU+mwVVDUmsWoaSrXbfj6hvHY1YrS5g2jt5aAbDGUx08q5lEm7EJAmZ
4c/7lEkHxLKjj8SfGNgmo3zorVNMXOCmasHJfL/ephWBe9KHryFnDp8jTc0W
nKRMqqcIXWPp1rmTMVJ4frE3zPDvLGVgGv6q7HhrH/0+3O8pKDt+vpUrn9S4
0aFsScvT4tM/kDuwyImbRu/nIcAL36w7vF1/Jm+dK3C2KWRrwNwUr/cDNSFg
ehPIVXui6WyVH7qMl5wJ/6QsqyE5lcxbeir7GjjsgbZkL4Lq/w9bpnMiuCFS
plzxRt+qi/bhCQfRoC36rh6nReaFC2Byawau4Fo8OqTtFTfL5YmDWQQUaPa5
ZRhrwZPvR4lcPF9k2vP27PMbp4zm3gU0mUc/Vdy3t+u1+sbA6+SXC/NN7F8U
sVhXBz4RluS2E2JdySPKeI+aDiEesJzNvg9IbRENeTBSEaR4cfkMTDbe4XiC
98bONJaVxrKW2edalXiSdBU82HIFNs029tzY23xIhkmrTDdjxDN1jHd7R2IK
fizA9LmNRlGPx/+Qjsu3MXOZM7lyA5rc7Z2gFhmsxVPPBT/vaD1N4gbfLdQs
sYDgB1cTTRV7AQ3ZkeEmrf453S3y2JrjYkMFfpqCRlFSL5fC9iGqXGFLHZ02
gCwlFu2YyEQmYzbNjCOIw29pucvGRzbllyMy8BubMeP6f10P23jedj8pqKXi
ed0xhFi8yPstOOUqgEaDAgTTgqn3xTMmunMKZWiQzwT2oyJv8ZpwxJEO8nXB
V4Cy1YtHP8jRvnpZKuZupFXb6Pt7mp4yzFn+DrtUT3+dQNqdmnGtEUGNYDyt
tFAh9ZFhdYrttKmvhzAadxcTUZ0YNCWmuv5UQ1btNEKEVrJnUpmD0fU3u8ol
mgEzi2gxGAc/NmPtFBkwtDfie2a7hqWBgZNQHn5jzpiujNiIJL9+Or55VZ+1
jwPnNMzakfpmVdoXqHa2cSosRj57VO+2gu9ricb1ssWw17b3t7Cuy0oOSOx4
vMyGNF0eibFW5xyxo9aEiC4E8DNZic/dZ/A4nKoQrQ2Vu5uJeSL1WH3yo/1N
Wkr+bmUDt0rTwOY8T/2oXKijPGuAcqON63gfKKY++UEQbSlOvG1VMC6zo/pJ
Pq5Gc25M/KFeJzli28egSGhMQ7C3ur4Db+noowLEM1Ak0tIEwvdNX3H25pUc
cxcYoCUuf+4g+BaMAHnkb2Y+b7e2t8pRU8mjpAmfIbJ6LVtR+DWSh6PvcV5U
NqVlXK9y6d5HGDTvB8A0VJEH5I5iX0fbzk8N+lYihLKmrEA/5mGjPSsISJrK
Dm5Je12SZKcbO3aREQ+GKyA4xpEQ5JiJmaneBY8R8I8UFububgOT922Ph1tO
Qaos1tANkZWxEAhHOWdgmPofy5iWVWaJa4C5dNx3J9+OoS+P97kkUHuLwfDJ
+9YYZn4zOaG22xq3Oin0CcgAkDLSJeao3tPXHHN2OwT38sWD2aSp7Sou5G0E
mf0a+NKpzolABtzzYso0Sg4gc2ko/kMYnNPJJK87RbEi3u1OXJ9YInLugYM9
7Jcs4vZKnWpvm2NVEbGXdK2JRPvLxuxETtIg3MeaIpjUYqv/GZ56TAuBDTjT
ETXu1tfmzbyN6cyfdoXfAK5E7OKWl+7Nty8B4CsYthKsvYipCmcVCRwJP9OB
M3OVrpypXp7v1qscfIpb+Ic4M/Ev9pX3VpYO+ktAHlMfABFvwwKH5odU2NPV
YYQfqlmAX6AUD31TIm/5XWjYZYjYKudfph2QcoXS5zo53R+hh8rHl+L/4lFb
w8TAgUA1d5K0oxQQJj52M/8w//30C4VE5zhs4nQPiHvEU37eIrGt07bK8Qrd
zWjtcyWk0xLQwoiBNdcwLWVKftGYOHuHx09iaGKnk/bh47SsTeXcqy8Jf/tb
sEWZrMneTIa0JeioQKQNEpZx7IYU7vuzpCTX6iRSVskILSiDBRH7+9SI45cG
JFk0gIC0YJOGW+A83Rz9T/MxH4kMeKS7PGKCiQWIjESY0XyVIiiBlXRcFl2O
3Mq3obtr9UTLIpuLe7dl0+Lq9YwZevYWmucSJJKd+uM6XM2mwphJahXb+jHw
3cCze/KBCGFp2rTnQ0uW3DYr6Lb+zVvGu8J6L53JXfBZP5bOy7hQXXqsNCSu
H2CgX5mSqh/V4O30oHTzdVDrq29Lldo5n/bVqMgSheXfr73abfggu8+kCdIM
O4RyKhCCQSNTT1IFhYE0B6hyMsC8eSbmki5Wy2clyNs3tEOWWH0iIpgYLArx
49qJXCccANizBRv9J/mH6Spci7AxJ4iaQrpFHMCUnnOLrbiuTiH8PD40BrFw
Wjemf5uVzton5xNqEgZIO3TwfOipnZu6pFIDDgULQQWNBgVM61l0gjVKC9Ji
FpYinzbRzd6jDK/hDe6dJsPszB1OzN5hrqdc2zweL0tA+4uqolumZREbxK1u
LT6qyOyCyIGgA/qLJFhJGdz/E0WzQJ2N2E4YLHAzms9eU+NAqu3zdvO9HDOi
TRBdHtQrZl+BgZtYNN3JRulMIjQnnhayXrx+Rz8xrbmwjY5i3yPj2+qypgWh
5NrwhRegUZEslgxLJJ4qR7OljK8e3MPi4O/nBigbkzPkFhws4zk9SGE/2Gvs
b5LDveSOgB4rnGRCxpuuj52DQ/ufPQ0bozJuAg3ooKBz8XpmepnKNnFJ16cY
X+m1L0PC0YBQL8gNZ9PpLGdqEmYpcEb90sObAHI4VXeEB6oSwQl2kXTX3/F/
t/ptBuMl+PFJkcaP9hJ1HxJHTzCNiAyZNIeFYnjfSklQnGyLvWkQE9l//SeO
pTwzpPdL5S/F0Yju6MMLROj80MPmLNRmZ70+xV78eOgSiWkSHTxL2TyrKQ1I
R4NdlCovlhNY33dFuQfrAuE5MFwfzrrtPI0kNKxNlSbOCyy4QFU7u6sCFNxA
ZULZCAUfGr8tKRmqzPe5CerRhIkvKb97mEZJ/GlZ2mvQd7/hXZjl0/p8YPWY
Xh6KB0YMHTt2Ix/Nu6CmPE+sqS+/g8irEYq/jpdopDn68qajLeLxHBXAhhwN
1Y60fG2ckoExHiiUZjLQVqGnybk1n4baD6SeGbln3/kJScZlIncY4LVa20w2
rLFfnMnr+NSR4doBjqepjmhmlYpnDui35xaiGm1GMP7o8j78V45Vn8Dk540g
iIgJiELcShZMGJ7d5Sq9n4GmIn4lEL/kuxB862nE1c3mKNJO9qu6D8w2y1a0
hdw6reY11VQ3uadAesk2+AwTrEphGQ4f6JTkfC2Re3uh7reodAd/eLtYI9UA
yFnO7jVLZJxVwtlvbH4Weq7bek6OaGLphSvvdeIHeJCyV+L5U9kJApACY+k/
hbKl3UphTUype6hrfHvivNV+9YoKuBtgvXNfNH6oYV1XqVzsTRSI79oqyvyD
jYbXuCSitPdRSIGO9FUSn2M6io7AVQOCtZhtgQveDvbPF9vS0Jc0q57Z87XQ
uB3ASRLpMQhHUZj8YjCk46b4GnyriZkuKqGBo9QamcC72fRNGJ1yMSwX0uXB
MB8mXBy/Ijz+EM3oMiQRMGX3tgCPAn7oSynd83KmdBKzG8gvG36cupe1IGVB
Bw0n+8ypho25/PK7hf7HQjr6SibFlT9bfXKb23mafZV4/dgB4EvteqBtfxVl
NacgZNelld1Qj0X11YnLFWNKszSCYwQZjpFPX/Zy5t3hO12GXF4HtfDpSJNs
hiH/36TJtbSZG4bu2yfbAq5GF1JvwTqLmtELsEIztwUVCYh/52UgBNMFtKFt
1Br81ZWolU19zvzmz5+oudMB9S+KnvXr/vPmkcjtajIlBeeuRW+UyP98aAFe
0eL5PaAvZSlCGUbaFQhsARuZJaQl/T50CoAAWn7ra3uiSUF0bTnUpGSvp/ZP
pLuseOYeZzhaJf6fXbHo+IuYxqLwbI4ichKDCvtY9LqMOE26IjbfQw7L8VZt
Q9RcDDbGSCwz63JwHHT2ND0sOdoFw+PwV2MzBFgFKBhSwqvBl7zyfIpAnNtl
U0FTiyVCw/h1kKA+fWJazfyl+IgbLPVWhrF+EQ/2GtmWYEr02rZIxtn+YSQT
I4WAZNbTVHjqvOXOBZFm7N4YRZaB2HduC9d6/Di4O+7eGahZG+pFw52TyQ/8
mISXjdQ08LwCXCn3VKCCJEvIhh0LK/bEUmw4fuNgxQevzVFbZ2TWTwa2JFWS
glEjkMpr28xuiiUSA5KYrc6tHfWMVQ/F7EsNBReDnDcw2lYW7OlogZ7EeubW
IwKsyY39lEGrMmIJCDhvc9QaridA/ZqJjoTkY1SOWcbGgx74ck1n3kYAaZpB
GHNvMnE6NO+qWx9qbzgHXwXdH3v5gMh2NSDkpvr/9kbNepTUNTgL4IcjuJRx
KSZckjqfWDhTAX5ddieumK8lDVJiTHQmGKxavZ2u3oIZyTiA4e0tARIOh1+2
m3u/1NfWJArD+tJOOVe2iTmblgt4r/rBjZx8pZQXYbtZVPbawtuIr3M/QETL
hWlDeZfdBQrahWYgoWYY0zOQEUEw3tdw8Da8VxJtDcNaT+XJSt4ij9X04y4W
B3Rii7nf6OWjlKDmJFe746dHIBQESeN9OYJeEeTkblsP1HE12+2tG8/BqLOU
FxVqaDps0j38C4M++bq1AX/e9nXt8melRo6KHfple/otIY1iRWlL9ywr3EBg
2x4dN74LwPWcp7Q8dXzkGXt1WHzVNpkLep8PPEnXY1xtq1yd+XxkONybYMa+
G5rGeTDbK3nOBIRqHRPsDIROl1/jqjuqA0bdoSU++oow3AJjpF48Xol32bRe
I94pNiFRlnnysuGAfF4p0gOFrQMQ2gWc1PLE86yplrFLj1mV73rIibe1k0EA
YSzvkp0tauQjVgSSDIxlY9MfLeUES/7v+umHK2q2HC35+8nTe56sKr5nv290
yHp9Ep9loK4NwLpY82S0X4+9qqtOZxHNcAB/dYMv/Txt0wHmQN4SUgoz+MEa
AOiJLtsQrINjJufpavqq4eNcycFdBx+xcFZSurvwci6s6Mafj8LYlzi1bkbQ
SBxG0YAoyAA8Lcn1HC4G0rQXKtwhtI5KqRPivkKXgg0XwPoJaIHiaiyWgEgB
sEdyr6K/rU5hp7zaF1lN0fmPBrtQq+0mvqHrH++ZMEfQbxhgD9W8xf9c987V
T3U9eThfwz++v/7OM/Me+TA5ytvmZY5Ok385i4Hd7FzIZg63FDxK+USNSehx
k8N+D/z+Q/MgjlpsM9vPwZhZDauifGNitsv9Z0tZRPQrjc36Rcw9FzjKP+gU
0YiHZg2N/0cn4a4ZENxBMSP81cS10CeBIF8iyOndgOLb5ZCI3umIVOMIGGu7
KZyWpmdTU2z2+z1Ut9njJDzi4L+ELCpPyrr+vUnxxSjPrkco5mamSgOOV9Py
NEWH9ScCWsbvjoitYt/uISeLL3XxKeWvvqeyXm0gdhBit1yRL2QK5wt32x5k
wMukOm7dKWGUMpVOQjnc0ltsJT5qE/8/o8aZdSDZzS8RP+k4OyOG6jb7JP/K
qDrgZFNMc8fFbaIXfJExPSVLBVdYbBRtgryBzZgvNPH76lurDkoaaC4KEjOh
kxSMyiTEiocnmNB1TLIPp0EjZJ6nv/rbIY9AcXioepYdiu5XAkfqbTtF9mzS
2FNF+PIPeKhEGrSZ9Vvx2YR7VtWw+MbNLijIb2pxRh6MMaqVLZ8DG54n0XiW
b2aZvvd6imyI/dig4DfToRAIXzOigJEZMstVqoOlsQkaDF8gugaVpUZEAlZk
x+WvIgHL239VDQ6aPL0IBgOG7iWy5Cub2UyDad2UDCFD7gZxAcR0dWfOja8R
WgjB3QCh+/YQLobVlGjUnJAeVh6qhreDLEEDpWKLPzMFokR41tTLp8I6prQz
j6pUirl+5cDO/k1c5pwk94CPBYWboDeOBcCkSRpttHopVZrbe1drSzYEvSBd
4BlYTSlQtSnfMxjfFyShQSpdyiqvz8Jpz+REAFUBCxvP9JMHnyBJq2tDYMxM
T4QsouL3ZsriJXo0bZorbzIEibqL3vDtcHCl9mCt2wZjpqEwgo3Y/YEhCEJ4
JdoEIS7vd1Bve/6ob9dDWn+N+vkw95xgIJvgl5mVzbMRPhiBIsIgqfsGZmjF
GkeqlgBejK84De3Hf7DmAdkfee4942ENOxOzsImT8wM0EMb64/705qMCLI8I
o6wQif+B44SSqCAp6KkOCDbk9iwkEZPheNMvfMehyE61z+7h7xjLx5lYyxg/
IxbU+bI4EkERmjL11vTAdJvmxtphaHV2IPQ1p7OYLf52va8wKwj8IMoLvyyL
TW1QThyrfPlwP/+gTO4WyrZqCGtDEjmdEF8bDE/59zGn8r/WpqFwEC2kIAad
909j91R/xc3AHlMXBBC0zAqM4+3b18epgVMRKLqr1xV0itw3r0YBkJV5BqQ6
8dP+wKp4CnySahASloyys0G6WwaJwxaNVsnouiOap03qE6eZZi/L3zNkrF5Y
gyxOjAUTXOLr+vfKjzWfBKuaCcz/y1NCGBMaYRosv38QZQAcdxVFf1A+D+es
4GFcH508Nb/egt/hm3Bvb4vkXCkgtSV5c9rQQVth0IURE2HxCgxomSbixpf4
36GL0srC3Vb+MKbeK4r87DjkBGo8UO/P5bZO+xRwmfZErVdXs23qIlemw9Rj
OFwiVzmrnXP4l/NfK9b4eJGK409Vl0FlFXQS4Fmwgr76/QCdObOQX3tCjunp
tzdBdd+l0WhT++0d9Cqhj0lHhIAoXYpFPEIlNVY2SABJN+NOSrKVIqfUDEC3
LT7WT/gwH+pDYHrY0SXw4tI9gtSoPlvMWtkSVMZsAYT1j6609eoAWinOJCZ3
7ZLsT1FmjHYjs2a/DMHbEpJURMXA492FFZfKzJMuh8ro+7cfOM44KpIfjyfR
NcW6El/wvHyw3v74mflSz4zmiUJBPPWkRzzQf3z3VAYI9C2o3f0lMBTanpx+
VnmY5HCkfKJIXVx4snyFXl/c+pN4eB2htXiOUrm1Rh9u9c/P4BD0Oe0IV0o1
5AfylrKqWsFZDdcKbMgVwibFN5YdWakgz5E4c0Qwtn0j7PDhMHY3eLncPI/q
Qis6TfmeMq/ytZXBhu3D4fDRxA+1vQijgpQ5i/AazAEeaiaZs3lDUSWHbQcB
24Y4JXM7s24AaCQPSnu2yMiao4qKE2vBlnGo0FPyRC5Y4sB2W8PYodoJJ8LC
tbvLR7anc9rM9J0NeN4nQm0PBj3H5zt/yDaM/ZX2hakpPPCIwS7wMbhbS4T6
ae5COAYt1pdLYWEyZhG8c/W6HC0JSFfhudzTlMbaz+Qdr1QZ3xuwoO4K/uGV
TPpGb17dkxf1mKFEmGmHd60twbHQV+d5kim7kWyP4syMtyEvL+xvb/XygCBu
IZYB6H9GmL6PNNrBUekuwdVK83Sj7dNl0ELwXYGA3c14MfReHExpudOKrYZk
UagLQWEg+anPc2ENiOD0p1LVzAOHNQs0BEhBPmyKmW1a9mW5rmf49eQhzZ8l
jssP0iBPqA6I8E74L3i6Daklo+UaYWOog0xOo0WaCHsfdU6Y64tPEE/nM9aG
88ytYgWE/McVHibktbk6gaEpeJ94Shfzd/r8Pk7P7LwYwWz4sRi0sicpgdUR
r3Y+9h0sq6b8FKxpEuTBFnxCEp5lK51rufO7H76ZfOAJ+vnNHC5hjzknzVb5
ZULPh2Bta0xQrBm4sTswpMFfjTC/kQjRSEh4E0MLtoFX6d4z1yA2bRTN+5Be
R0UcUBzrtr9r3d8N/pVHbXqK0nnY9+VpLFPHmQRvpvEbvueja3C9KPfFKdQi
ucLnH1ghQd9yZSpZ6DwYVclrDQWWuQKqdbpK+JYPOsC9oY5fChjuer6/Lubf
Br/Mzvdsa16j+394looOtEKEAyDIVXEqKeX6skptJksRpKpDLiIb6XK62jcf
EyUyom+j/d4Va8Lflm1WEwfpsVBEVDTcQ0tsU1g2qZs34Tt27oggGjSAB2jT
TGKRVPtj6vAT4uA3hSZo6oTsSsagpV9+lo58rdu3tnKbIgYR7RpmOPbswH2e
6Uzb4/kVZpB3LAC1krbDWAhCRjJ6ckUmK1KN58Iw1MAw3AzSxA6kh9iJgEEQ
9pPJ2H7U8sJfd6eqelgj3fNHFLqHEwYpLD9NstEjtSYz0s9SLtBQyJ8ZUaY9
ShnTM8TcXDjjoMKQGnGfKGG3hDKDHkoGO2Z87tIp93nLAUH5Y0zf+k+VUTRY
UBQM4sl9SK4iuxjNuzHhBoWELEvxM8ro33yIHT0L3u147IPyj9q+w1uVW4YV
k/Ax/jnSW84Jq3cKDGhrUZs0D+RfTW7ah/7IcM8B1ItDLOo557FYuFobyvyA
UrEikXwz6EdpaCEXNbc6bFn8sksDeyJUUD4BRUL5nB+hZi+MLc17HuEByaV+
VS/z9wl5h2ns8ArJ04QUgIbR6A6y/pn9LB8dZUJQ4IDLX9MZ2rkBdbV0CQ30
+9c/KRqI5vZgtvImiJN0ZtxLJ9TOj2TSI0ymQ++8yS3XN72GC2ZFp3jX5Y6D
9hZkAESqLIktzLvFE5vwa93o76XIL0IinpgYIlgivl0fDRxtnbFEMq3hs7cR
Gs1+ysWlOXLy/ahdWLzxuhgmOxH4VhFT4JM+XlkRQq+Fue1zdzllSNm0LcqH
pNepBaP/AwfBgDO+fNZkY6IMYSivEmg0GRCvgtpdhJuPTQALNRYLDBcD7iug
0hdCNBovcXv3uSA3DqHdwaogXFr1RNphPdm+2gaLBTqFve+iq0HYUaQTEvWC
TWbKTlAOu3n3EdsnZtNavyRjExP8mxQHJKV1LzYWyB3GFpO+RGrxGAIK6/Zw
QOXBNSzEIviDMb6HL6B5+1Lda/qMlgdzp1M6IHo63QPzkwW03EF3Gc2Om7Fa
L6BwKY7esYzxpK4qPKPpzR5v/jj+Q2jlVIfC9J44KDQT0+QJg5pQ0ccD+A5x
H/YFQ1Dd5BsyeyVXFnz3JR+yLMKt7h+IeOXS4/yuEWc3iVGpNK4HJCWTJC85
Du/4IAiLWCYzn8XJoR5EfuZ4sBlXp0PPTZQhUY/KxRIKYGES8B9YSDguO+SL
v8rTMg53VWHgLKbl+qbcvNsQO8N/ZIoMHtDXDIZyy1Dvwx8hRYgGwM6IQ5p1
wFabaqnX+X/VHK3UZvxgLIZ4qXSbvofI8hoaDwyEVEIBZsIhGYb3TO+eiDJJ
vndmxmmjvwYRO0bWCXjFnE2F3CERQKFArT4b3WdJLTdk8bPPu+3iY/l6ZNE1
DnEVgkdq9YHFVPXqr+xvdIVzj4tC0UvRIkJD0atHT+XHmUUTpME2LJgMw+j1
lk/D83uviuPaPSdQ3XbywlzCQI68BHcBsfqModAqBo7O5F74BpTeBnqjsTtA
hR/6b4cRRdXV3K2lTXr2VnIbPxlfCHf0imIo3KScakoOYBD0eEw3/fCbiyW2
JWEm+jXRhAXm6n4HJ44L8J4gBKrW3KLZPudLDJyxVnDZFhby4DFHPtg1mZ5+
6bxTB3gRKG/NpvTaPTxPn4MvxDKY7zrffHinqoob8DI/JBMYAhzAJhPIl3pK
hZT4ZnhcPFcsUSasBZBoLQOPF4os4qyfg4F6QLlwM3+fF5fSacu44XDqzvou
ZWCVBZgdJ/0uPgzplA5hyXU1Pn+PDzkurZ7U11wt+b3CQhgHaCoi0ggTbNF8
AjYIELa5aFX/Vy6ieFrRRQmbJdK9VTouXDba9YJ3saZWZQ8miDaiwUYIifNE
YGjHReupWO10P7XMCT+KsAX5GoRf7rCp0eg7IAK9OV4JKr+xgj41HVTbLtRI
b7NTDqTPe4kmjrZkznuZiP4I+WErwrwqJNwx22v8QXaHBUEYMaRbCpLDUJW0
dvBKNlRfUcJg89zDnNsFHTjqHkw6qcr0L03ExQixsdZy2ZxtOccvdhpQUrb7
Pt/I24emVUlcHm6TuAKkhDj+lrrnzci8F1ChuMJ4DY0xPXsK5KxNr7wF4GJ4
pwv6alA54A/JFdPZpz5bgfHJ1tWBZkAkSOlxLTUkc/b89vDSUXLMnQKJqZmr
8bz2H/vO+LWRRusK0iX5NwjTyz6VB19wL/i5vMupEiCVBdx3SHbuHs3ixcbX
vuP/HszOIkSvWbMD+1FmkUPefNsidUxQTgaUkH6gicGKe3MveSNHZF3aA7+E
WPpUThllk6DDPEYuEy/HmhPOru4m0cnlO821T0VYjclknU4TWl8dl476/is1
vcsCjMmu1bBXMNi2wtM2CDov6uB2jVF6RZstKUTVC/64fqIdWZE+xUhRQQg2
RgFx975JHnhgORdj+toGrh89A3+3Tnr/NTuTqDfm/leWWcblAqL5Wka5dSMb
22UVZUmFvNsYQqtlTQiRe1LGASqvI7wxcVbm4hhPZuXCfeYG3A2uSuzmVie6
xAANDRw9lsaKlqIg++sXgez0X4/5vHBwjiZw688IThm0iMWqV77F81orqP0P
CsQEIGDbGTWMj/052ol+ksbHhYEgUmX/gd2TgmZJxe5ejzJgrlptsimjXNW4
PKdar7otlo3AFoLqAXHgn3g7LBfo2rwBEYJ13m9OVDFER4egkm+MpRyYwu8U
Okpmk91bfigDuYowgQ9UTikbbsKd4juefGL6mBg0zxNnUWVLxVUcVmP93a9U
zHwY5dqlCd+hUk5sz3OEsID62M2+ftyV6cWa8XfNPwwnOTuToXIvpzSSpEF8
cu3XtfOfEAZmoNcYTQ7YYILzWaVNNgRRjXUKTckr81t2WAiN03aHunOFHP3I
ErRa6rvAh1bvpFhF75VJniZlYkhv31HSeJvYcNqxwK2eAI59WVcEgIUIjlA5
OSocdSaQD66KoB4l2Nou250sQDcAIM5+Hwb8zA0J4A1EjZlxUkgLrCtAVuAU
6CQJM5RpjdxELLv6qrqUUmPVaOsNsuF8kAQ5Fed53qGgnE3PxZJusFg2S5AO
cMBt7oP3W3a4bxTsMmhuxdz3QYHljPWiMh2D8R3P6DYCgUpI1y2B+gcY4wCg
8/9QTL89sJejhoHFsS0PpayBQFq1kDheLTyvdF+uMqWA2d7nVEkSv6y1Q8fn
A6KeFa8s8CD6mpqT7M2SUmEFaYHU/ZiIkIbyNr6gXvTloyDOPPzOOKgvricP
Y3fCNNV1QYrB0ywkBfTMSKf5xsMFmivr+z2JkV1RVHnxgeAiSAa3cVcz98lI
RzOBofe1TxLus+MdgfeBqUIKEpe0kLDrPYJUY4JnNk7qPrmzzI3ERezn6YGD
Q4mYS/OdbbLR4kzTMVUo4l9cG1TD7PSRcwTsM04/ZZOrah8LzlrX/8h4mTz9
Tugp0/HCxo08iu/OY3jUz9BcEj1afpbNrMmv40LUIAwTSZA+MzP3PZL+Ezvm
acnp1utL0aZaiejdeWANUdxRW7nv8JZSDrx7Mh/70FGPex0sVxKO01W8Xwfg
X9lzenzYLKc5k4L0VR0BbI0YkmIf9hgBlSkWLBzu5xJ4+5AVHaIiEHKwWEYn
kEUVoRR95puvgMvxynjIuIz3so4ZmJDOyx+PeZi+ZcLCB3TYO/U+bwYC3SHo
BVBqODK8Ufq9GJ0cNyIJ5Gm4+RM/pXxzl6YjLPOjEMqPk1z4e2QSm96+mO5i
pmmT41NggvpcqH1z621TzH2tWAjJw1zTLXfoLJzEK9En5J1an4TLpAEIypZ8
L1ieFRGJRKcm2h58K5IoP+hQWavxO9xeMWSMtyEwYGWnnO74+7HA33FJyJXn
D3/AAtDEr0tbDDCkWXR/TIuznAK8cif/AYtH/ten1hmeZYjY23E4UoAzPRvr
OBHh+jmHa8hlR8IwflXpSB12nnJSzysIWKfiF7oGEtQSGmQZPOFFrCqyIYSD
Mr0IJB+Vpc+wgcuKIBtQi7aeeeQUECplklZNEx32BHSFc5yJX2buedek7QQL
GvGui/nA4aZi6/Wul+dVJLmKNqwsswUDU9eMnVfnkEJZgSEvjCGa0/za47Wz
BrFD10WypzMqDLJ9yUaMbzxkATXBwKZRxL17Ju2RUIor2Mc/2xCnwECuBuzY
mIPdpKsmWZhIaU82tYQms9s9YYDgqB4gxxZTOIGZ2AM9a/MTtmvBIZ3WfLQI
+JK+ruGbQKEQAUsNHyA/Bu+L36V1uxoFEgqtHiL/o2XhtYpYRIzr+5xQ7dze
vzvKju0cei2BosFN20MPD6EPb5N6O5pb4qcaOl92Evqk3H5E8yI7dgm9gQJD
NJjyxTGgDc3Y2TtMrnKcOxxB50cniNuCrtdXIN6o2aF3pX7V2qALiw7Fjn//
s3UDKAdNbarFHW4FCMUbywQ6T1inarZ55oyfVXqhGwOTPhgq5fJPqxyIl3BF
3dWnhi2v6F16utiBuXhaNaLZHNCBttycO5wWS+1jsFtlNdldjhk0J8WT6y38
r5HhzdG22pwqdHZ8W18PG6jpZrjLGrF/i+onwDQ16Q6CFJ/VzUNO34nJ8XCi
6zgGpmPMAk1hML10K+VhMgtnOBW4bW07kH7nREVmScrUopFWne+lkbMTZ5A3
CciyvICsL2VhXRwSpXknbRTqUTg/qZRriiF3T6pKMbQWx1POvmeFpRkgK0QV
KZ+vNm1hjcymMkA/NfzmEqFazx1oRWmvl358FnHRi0InLxaDiMaG7K774c9T
nUbRKd1YnF0H0hFCOWF4eeZvDFJv2NJX1PEOPPIvk7lh0zqSmtmQXEwJGkGD
IP960eaSgY4+0HpPMQsyqJf1r7PYoZ1pasSwtaARmA5ncM5RT7LYFPbVcy+9
oT27OBO2fIUEiJEY0B/KRKsfdV+i+C3yCwNc0ltC6jO4gN5umjn/HSKBYkhz
NgjtHm0wtlAC6LmmUia+XkXfPV1Q+nC/3SjhmjMsCX2TNqxuo93j62UP1f6s
Ieibot/xyDVLrUovg8eq9Z/O7kENstlY8zs/z1L8fCwvaFbLrQbtQI5Te/K0
9vQtvhGM/IGJC2KELFa0Bw7QgiEYg2t/BlOiTIX2It5XITrWsfFsXNJ05frv
ClDHtNPSrkGzjKoefEn1Pv523cwl4T/d/alGUTjPlMjKWE0yPcTycnh81tEZ
61a3FfYZaFZJ+SM0pNbARGuwqAHTa3IpqsH52C0kuyAVDdqlpK0C/b2cmfuc
ezvC7SpiQFO0JYPohlq4jj+lZmqBJtor/axmgqTA7Y2NN+6ieR/9yi3m10Vo
5edDZKsE/A+iHCT2swqJG6V9jiUJ2RFn535cDgxOZHR4ZUBNdUc48cnGeC6T
dXsvbBDc7Kr4ev1xzdpdGhT0v4/YnsVztpdX1jP20jPx7JqhbXjOSfzeq3kq
GPBxr/hNTLsBpl+fzmW9tjcxfVpFx9yO5ZGiqP7+KPMXGLbyW0TXDwWbbEtX
nFb6JlxlnVs3jJTR44dfvrXWa5spM93DDZle9BV9lXjkNe8r+VbOMoFVBhQQ
hJhj8mMOsacEu9Y6jFjdBDLmBJmyvDseTMmXDEjHoTnD/dfKjeTe/L4mKAG4
H3XjP1+Ila0111MO2eK6QUPQLnoYdg7hH7WuZzZpvc9RaiWUB01RD50V+IE7
QIqU6L4LtpZuvXSKG2VOmJNKC3iALPd6+ne3yj3V/Yx5Nh/7/zQhLOx4kmeP
OAnurICTgGnbEBpzgpG8F5gu7AjG63pjGJWHYCJGOxz1xrtYBH39ebcqIQOc
cHX50oHGG7FI5wKjw9E4/ieFEJQxJt64DMRCU+D+HaimMwHZslIsy/3G92/y
EJ1Ib67opo05ll/R/15IecumQbCtV0LU9aOC1MJSUoQDaGv+GxUV9PynoI0d
nFoeYHvGzBhOOXU/zHo1eNdh6u8Wt1mRIXqS/JE+kyrU9W3bIGdlX+ZkMeM8
9YXLXP7G5On1+5CO3L4jGjMZlnCMqEB6rZvaYpazPHUBWYGzD0P4/fTcqOX7
DEFxcAwRnT9OZCdaLXPuTO8NdwMjWQxekyHamZEd1zUjUJWhgj4kb25i77Ar
Hkmtw/lNXfpkeQm+r90jGXpFThnvQTXZBy/NFa+/hMgR4K25dk4BULDhpJmd
WVpoMKrS1mzyHDwP+p108EMvE3gc+aXPL8oK9tPlTUivgwB5xnbcdmEPIZH5
FniUXHnVJOHmpnYJmph/idrWwp4bKU6ZCl8IiFf0+XiF7HkrIfsvuCRQ8wH0
DO3tVZNed5VihaGa4nGrTArHflGes+B0/yz6YseR8odpr59yYV91jmdxGJZS
Jwl8g2PlAb76KskCAvwHoK0CWGmmUNYA/vMFUuLzfYpbV7UHT1zud2sVZIg6
t7gjgugZD6LX4zH9IpsAk5Eko00143A7XZryEnNE9Zs33IAPVoHGGSlvWs80
Nu7GqnqYMF944iO2bwTDAfw3G6AuNo6pauZd3e93frhlT2Z3QNUttC3JU0xW
mziMOMNobB2RxpTDaTbutLh2Kre0jlIbpsPwb+D8O+xwVm30BM1qxvoCNOwn
FvNOl6b+QdSirOFTfv7CGkkDgfItT6/cAdb3YgtWVbORBt8fLAoU5cUR4BJs
n4MAazgEqT3xPtJvfaFE7j0VukYxRzPMDpQqWR0j9kcihAFQhEmIPY7kH4Ae
vTkG/1qd4+g//7M/6g+gB6RiiPY8LAh/T/c9sFiKbKPwT0buDMTaPMUtEGwo
dQeltWrJNADensPqK9dfLGWHT3fnn/jgzTqsw6JHXEXFV93wZhyTO6hndnTF
GelCucH5mJHIgG4Zn29AH0F/Eecs2dYYg42BWCHfacT5QINIGofAC0yfKucz
5HVxKKxd8JN1XbuTdJTwYdznTgaY4Y1npiJRt9EDlvzuetM64bIYsBtfFUa+
x1uRAoiEGBgr/i4J3R0etGfHiZnsCU6CYKsI3x3GErSGU7OXQGL7W/E6vDet
Pn4P/MVo4M7R0SRAhF35CiCT+9oFGzmuL7Qmt0VDkHpMEvse8wkb7qQDJu8x
7jOfo4A5MxaBXRJnGv8qRqOPh092Fi5eXTF08zsKYGNwizUVtQvbnDWIcvNh
fnWGzFbH/zs7/UKCjV4P0yw7DNbr9pOX3MnPPwRPdrbdyY7qBTAD17ptYQOx
MxyqeyqnFRuMPVOyUWsJpSzTNFSdRptl/rHtrdd5IBOuOrOw6Cr5gooRhMNZ
abgwgDiakd0JrvbpW2yUNgZ5W4EezMWjY6mXUamQw/SLPFujfCT0df3MHOWs
TWYZbUcGTfqY+7Q5y8pzT+n1S/+DWON71BQbQH1f99ELHdvSGaL3aqFcwQJZ
rAhjoVWj8Qis79V0/j0JrWMzdF8viJr6LKtqVh+BFEbbJhmG6jsg37clrXWV
EuI1X7ElkIt/fB9UcmRLO0O2SQfvBBbEPIYz18j5Yo4Zchmzxarl5W8VjjY8
hP2R5BIVitlnxy+a94LtvRO3j5f3721SH4MlWUtU9EbELKxx7FRg09qN1x3L
74d2Abzf84lcrs4/7YjLISboErns1X8Qvj+eZrzsfoCBq0mRvj+QBvjy1huq
fVGLhK28p5Js5OI14peAnorGCpyl09Rl9TormEbz+vwrk9Qws4DVARKCjOky
gFKh1BOZNsyc6NLqVHdKwyWOIvCYXam8KtncSM6XADNwX0NM5FtxYlk6exVT
wC9ZkErprxHhXQVTmy+eMnU+hQ+1xdwqLCfC3bDaPwjuVb2ehUZBq6D5haup
o+HFia9gxBRGILWwmfKKSR27FzMiW3cBgqYyZiolMl9Jl+k1G6+iafjnE/Ee
xOO4d8LtSRjH9pKNIlOAsUey8tQh7znsSPS4L94yX1Uuc+8jLVjdzmZ/uZal
RiDUEUUP6kkJMQIhesXuj7GVAtW59PJZ6pQ5RiaicKRGiffbRLZAoE3lxFsX
YokaD12om80CKlnqy5W2mWwiD77Ae7SL+NHSmLYBNZFlSDe6xj4QuyKvuvvo
fPagLnk6Db39xJcGByU0QRtDvuux48EC79t/wQlAA/Eeh1GJEf/j0stuQWh6
0M3aQ3t8I+DtkyA96FEKwlNe/W2LQv54FBhODHt6fAhRf+ni5yjhiwQrKchn
9rhw7antQyq6yt4U0eEpw/rx3aoBY3NWwtiyD2O/skMFFBqEr7y+K4wfST0X
AQ7FI5pVbq4j7wnXOOpwh1poVfoDztra/1PbxyOSDKS336TGmXe1nNW/yADB
C7tBymOX6XIO6KaFGHHUV8ZLymlpEqn8j4COwRVrWbcl0EFH5a/6OY1yfoky
qonhVBcyLjhXruKy0oWF6rwhYG1z8KsvPER9e5K9l9NBST/bTpKEYUIY5SKv
kTj796+5QQzmCYf5HNmQVToq0yY47ajjP1YYCK45IFVfaZfOoXzNvdt1ylTK
v+8giKWAduwVX3FxcKP3uvvabhY3u3YSu8BfjrHRZEzFhst5HnX1a9aYbNPM
sImvDAe79dZZNhRTijG1eo0CZS8m3mR6AzIxwTRfR1IqnCy+nnItSf1CpigP
bXbE1PYNHMwtHqiL8+NSwlMKGBFbCwxVdrUJGi18Svng63EBUsG4MK+/oGrt
GtoR9aYVeucec1aVY9BEpBfLNQpmmcJz8x/HRtS+5c7pHYti8l8bPnbc2p7S
X5e36wGPnUynxiKv3iEXO/lMarsRadgIfu17WaE6sRa03MlwAfexnTfrv/t4
jd6PoB5XYIv1dXq0+Ct5Cfpu3274uFlyqsBckhmem3jVr7YNSNPXJL2ebCzk
IZVJNyt4GfJemWpVF5KWCihVTmJCjQaVEUOSpVNWY4WvCOfeDeKVzFlOCdfn
8L/Y7tplhVFCH66nsXRywonOQQtsTyZt4BpllnPBF3urQju1o+7rxuXaiS7W
rTD77SOa8OMf5iyX/Kn6Odxq94kSUidT1Dcg1PrpBrq3fLf9g2k5vR8AhBTF
IBfEHpXGa/lSJnWfAcXuLAwNnfaXZGRxP4zdnP5LvgPDGQwkd5neye0X29vo
5chfGQVcLirUvB109qb8hhrGg38RrHexoJzI0XA/Ln3ZXCUWhQ9jHZDlf+UG
XzQ8Pp5cPBaYZU8JvBN48FOBU3/RZ54XNJCUUIM3ZBftknT8J1IbV+1piSwo
ftxi0+uJz0uQ7PpzFIfuQObbHABBXKMKGaFvt+N0lntK3gB0VAL1p/GV2QcW
75OcxWb+2LeHCWSWdASK3Ro2HdnU8FUKYA9nnFG7D8r3TezJax56ioDOCKnH
L/UDDzBkApkO20v6JBRViIGmfLNwdTYIR6Js/KQyg9bE56QcT3uAERAKjqRN
JnaNrQZYTOIR5ZoyolPr8VeaBRvq42up1a3RyOeRN4d0IUT755/i4qukwpj0
RcXijv97C/S6L0hzCSWJ+EhVPTogdSZmKMvQByW4ShV1UmR1vUf9pY1tjDuH
dsWYyDnb8uEjgyVmDCPe8uvX2Ovulp3QXKx2/KvL9ax7XjEtiYHOW7aM/Tmh
aXeC7A1LS2n6t6BSwDSrVWNEKMeL673IgJlPUFaPF/CskJPVr/DdhbKZADYV
cvd3NRtT3mx/qWCUSG+JsmNqRkyx+a15w4RWpqm7hko0ef9gNSCr64pKWQq1
7EMbs8A3280wbiPrkh76U6wmkwhhK3yHea3zvAFBeoQ04f/vVZcnnKXEGqHf
AUQaduYaxTaqJSJoTgweY68qA2oS2nKZ/G7OE1LiZHstmp2dvry+ZjP8OVWt
nOzOzMIeGnBV1pPLFQJE/on41NosEiRXV+ogShM0bynlavt1Vluqu7ranU9T
BdwbnXPvUse9x3JsypuTf67EnpCr15amBMWv342W0ygrhtxY16WJKeNHitOw
3qPMx7sgIB9VCY6s8uMr8U83V6UWrsSJfsaH2NeKtYTbyX77S7dQtknqmDsr
KgamhAf044De1sANze1namPNO7OemRc9orcF8hzMZAXFctabAwaTW7av1rOp
8+Tw0amXwCsMcaeyOhAJ6LUgyVu97I1NGANJ0eXP7nA33LTzFevEZbXDCg7O
oHDnTFsM98KDFCcYJDFAddK6xf8hr7zFGkm75OIo6IU87vmW1jjSlPtETAMk
6nfSq9OCSL4NKq+Ddft+DItbF+LXPQ5b8xNyTSMknx/5+Ze4VR9mPwEJuwQD
v5reuTWpKV5cINEcBXVWKjR9vL6e+Sztkc0vu766oMbT/9NVd0M+PuUtADyc
Ob4dnQoWIYjCzkUzNkobztyDdPv6ef5nFFxlCYjrjp/B7Atu8iTIIhUisrqL
UlzFCBXj+cyGQYqHlH6q9G7RgcYH3HLi7IeWhBsOggy1WndvOM9no3VqYRdh
5IowUpcTyIZ2m/sWmXDF+LwJW2Yz4LtgjFr/wxSNG6fUmaalDmQxqYjNBd++
mYRh8PP4dhwwoqPcPQuUGLgU7Cxe+raQAzQ9JRePxaLIdy4TWelxZC8hwZTt
HebYzPCieoD7ofB808BPjsCNK6+uiRmqhcm3wvYuuECQSHKtfwJgIWYAGGP+
bGTlXI8uZPHYFQRQDCBEsw8bn7/IZ15wjOEd1eftc533UNftMBwHQhj/fKAx
F+I/ecRfLenfM1S84B5tWxkHRisDez0eBqNpyYfMJk67QSVl7swmuD/wkbMb
hynzGV9uyADouOO4XIH8Ix0pY/QSJir7yEcZT07coizjl8gRBF8PrTD20io7
8ZiIGWil8thtGNhiCGciA+2Z3I/RMS0RhxD1W6kYl5I3VBtwxf56sd7ms/9U
r+3A9+7NMTFobRvW3QZdiJTx8rhELYVbKHNwwUroybyVhFWa/VD/HSZNCTXW
zW+vCwIqn7fPV6gjlAH4uuIKpDZ1mOSOueeLe6qijBB47BTjmqHCERgrY4tw
4Q/znI/B7TlOUnXyJkINVwgJ8zW9fKPfvLwYHk+YQhRNX3Bul7Uq0KPB8qsz
d22vZ7eOvbIvizbaa1f0aqC16jtDwPDBPqusyoTAUuM0wUE016qL6c0ZyLqW
NKgpr4UHjbMpzFWLL8aO0F0eGbzvESykjhLgIEF7Idr7QPC0Y84ug9HXX0t6
f3Rd6+PE95OUDoXWCnBLoeLbUZr2CAYUmnkMqgqRg45Krt4L3W5DjjykFqs4
0q6MIGV8G33roiSIQk4zHzu4MEn7l8CgL9GmD02eoUvHqbbwpiMUrBJM16n0
09TfF2R0N9LmAuRixZqL7eXTzSzIzMMW+NZ8Q1d9NWP7IAJOeSMszeytMLy8
+63QH85NgpiLPl0MPzxoeCI1eXiTjWjm1lJs95LfhikUs3FoXl0pWhOq34sj
ICmO3Hm0AJWT1TnECdIUgV+U7CGQ0FKp3w5VNDoQvKx+A0L7dQ9qm673Ufo5
JPn/GS8KaIZL59DskcPNZjmh8ALg/mrGyr0RdeJ0okpjcHR0OEMco0CC0BWi
GnP2IwnRLiZz+UU3nFESp6GMVXfEI0yXRa47b1Rkvh48pMjuji0nCQg7twB/
tL7jF58L8w2MFmI3aAHIFtZejxy1wO4lAPPP2kMzKLT5OgClVqXETmkIvPLX
y2K8ZdmcNmh7/jWaEzHE82A+PsU8V+2StZqRtadFaK4SUMNvqSfgT4yrwRSh
XRL7SjC4/+F37yiKQOHrJxRVfyMnfmwIB2sOJud/Bn33K57tnXGkYeE5CC2L
6HHMaacgN7Qk/UX+zZvZfaYAfUEvTRqEfodY5w4CTwYKumjYi9tMbPW5hxgE
wDoyTV9mh9eU/fNJ2uaoCJJo9qMWLIi1o6kLV1/EoSfrNSlXndZ221MgOhOz
XtONuJq2ilg5dcyoLbGsXEtE26xTUmr2UXC2RSaAK6AjUcATvWgFDzeV3IDL
J7dB2X9Q8qkgAUO1nHFKopfn9Mh53P4hQ7k82Cn9pRbWJD9Iv54k/Tc2q06W
LHAZS4tqGs6MuFgV0c1pTk7NUeirA8ohQ5qe4s2DZA0SxA1NyG3x/eepQETu
qwTMew8cmdUBIxYx7axbqPbSmZpoDx5KJWAne0RmKSCGYp0H876O3iMQKpDG
7kNFeqw9LriJcKRaa9CYpCSIcdYAbr80YQ76CkHs3VbPz+iTufA2HVvy2u9w
MfVa71gIo8TbO5KWbmynSf2SdLbL3oU1Tumo+p+qoA2Dig840SmKNjdSTAD0
cx7pg1YP/ZM/dcqq/7KR3Wa5PXXCqR1D/kwIb+IOtJAnLCibBIroMLOXHxMr
6O3qRivED/q3Am+3q35oLMAC9lrSKUPZrr8P93TyIbYwbH8OLqUnWl+c3s8k
Yi9zE1Bim9Acn8wEpY0WMb53QpDFYRh2p5K0FTuLYsZJnPaIQ5nCnLCcp0ug
PuQaw8ijiTeroviwSRc/T8TnwTQDvDR9HVDzyqrOr0JeUZ/L2E3j9/NzwzwV
L3GF4Ri3phKoJatQzm42Uwgkg7JK/8hdjj5aUnlbyEKQodl2ty/3J6FEPCpM
MjxXolD4zSB2CAilqnp4gl3JxJnYZEJWNSSL+VE0NTDopcAWVG6fHeHFqgd+
Uk+wZmuaBceRT3miLEwdxSyhzbNfXPX9v7AKmfUAZvZTmOzXRRZbhk+CCcL1
+179MyzS2lJrHmJlNt1qlLH2LYcCEBMCpeZsEUsC59ujIvS7r6vJLcyge7JQ
sDoIKNXltCf1c0pBMU8JPAALvn5WTdLQ/0/uYW7Rn4jx0Mm3P4czJJvHcdLM
RF8mxMy1wPXJb37tpHqXnvKKa6fpo32DwOMKULw1Z03426QAVc3xznk/qylr
HBQic4tb6jTePFwLSvVqoTaXGsRtDyPC+/80aHaZ5ywvfXclXWSS8vFSRkOs
d+ef3OHXV927OnnVJfyupnj6e13DnEY5jXDQWikMT3dKiGC2FlfumxqPZim9
tWoO8LnxMAfXiTsP3ypkESTzGW5m62W3SW+G3kSfF2WPBW38UxqY4XWmz3eJ
Ve3jmxZY5tn7k3AclLk9jdelNTqvVC2LpkJ/Y1MRFchAo/wh7YspYROV4GUm
SVsMLX6FIym5gKHHbL3+KVJxSziJi/NyyAi1MnLa1xJR/o9e5cXwffhJCA+z
OUkODInnw+fahbDGcvLhfh9DLooZUizfrL/1G4+xP42lms3MVmJ010P7DX8F
Wy/O/o76EhcCkFpdJOlUfkqmOWyOtbqs6UMSAF5uV3UBqad+y3K/20e7hpai
5oWinW6IQ6pscSG1TYHYaqR2G201Jb1EE9B5Gdj6LzyLxBDQkLAn5ZFYtgux
TuqfANqqT4phWgdLQFuCxgFPy6GJcyj/lS/iDBLXRhZbJdeNPNQNl+okQbhD
T1MzOZipXakK3JRq0QS0FfxVcMBta9ZXy6fY4inCVZIyq/u6vu8petCLWyhE
uWXBTbpeoOhkESLC1+MAIbY5jE44zEz7X2gjO1X4jgbhCmBkAGla7Ebt7BQ8
81+IQU4oQ+1hQB0rEtoc7jMtpwLkaJsi5DM5IgnppSf4kVl1S6NjJ8a1uNrq
3GNo5uOsIYntmQ2kAoRLH84Q53/HW45sbHKi8AXwqItXvtxGcFKfWRG58eVo
GP/e2DHu3ZMIyq06oR+yeBIvjwwMsSu7Z6n5x8JrSM5AxkqMPlO7JBPhEdje
hZ/KwOFjecNtebuJYeSEhb6AYV5o4pvF3+lCDB2XbSAK4Oy7JX6R4Ke6n9zZ
B1e+nu03acUV1KZ5GUCo1dKsei/iFn/HbGm80ELmLeMOMsSLqGcXhvDsFL8c
pINMuTfEfGnZ0i3P1adk8j8+qURwOZcip6inw1JDMsvcrhOp6uHF2s2Lv46z
9QF9/4XiDNUOkt/3850r4WADpRBH51Cs+KHxk7eF9N90OuW03mPLSz2S0uUX
OeToifvNnnOAsIxiEjCCZ9Eq0jS8mxTnl53GAlRmdMCG5a7VVXCuCfm5Tu/v
B2fT2HtYk553rRgChufQ2Q1A1diWpSUoyYjxq3HmGy3/cHowg/Qy431/I/+/
D/vBoLKMsGwRJbmr83iSlDp5BHlLQElJYnczIdgXLEsVU9byg/ybHX9IDTzp
6Ajfdnx3Dj4Ii6H/OFErV/ZhnmptuvaKSAt6Ykhu0PFgB+iS2O6h0EkB1jcx
qW8vnH3htKCZZWtiYkdxS/nkYVgCGj8c/EI/hiDr0FWthZmuxXP34IwA7M50
YrAKZh7RUJM19o5HYB2uXPhwzPCfZ8Le67Bsmf11jUFIxwWwCTyBn2/YyDFm
j99Q5MHRrx5dVAwt/VUrFM+qtfeWJWTZBLCwSDNzPPlJYVHV7O7rrKBgcebI
JZUCAlY394Uug9tBmIoXf+WDsdcN2wqGveSNS03Th2YzZshiS/aV5ha2oARo
AUVl78vcztMgKeeUggqYDewNZ5DlYVnr7MSjAGKJZ0Lp+6oAI1tOxZDdLjTm
FAOQIsJ02nVo9TwfSofARl663f0WOB2aBuvDrLCMqkqxtlZJjXt0HNyFXJyd
wqaOBw5VN8KYpiTK2psdxp/vRiFKhXN9cOVI8exaFggCZHBDyfmrzr4S+qL8
R0FHv7Rv1QgAWib412RQ02iWIvlYdDKqgpKIZU/KHyzio9iDOabavvr/QjVU
TzZ94XVqDO3GtiUxl9jkKikCk/Hmx+yrpAdzj6jxjg8jJKOmGhS1BvgIeUei
3BYxczxge1SQZRKfueqVLa2vCoYnkA+GcDHTRUb6E7f85p40gZwMEUcI/v9X
RMIqITMQX7KjUntzJY5wvjTccJQAhWq0NN1x5a9ssH349oGZB8gebIXwA/nG
x5RXhIZM1E0gf4AT1fGiZ3bp+I7pmRV1Is5d4FLpgG2Ke0yE7pKYuKs0H54V
/3qxnEkkFY3sVe0DOjDULC8Fz/XmqFkhA8LY8Cyq1xMojML9Qner9L86425V
FUhoxIOO690iwlcRTIibYCMSWE/VXrUHBoibH9IDIFaRXZve6Dqm6WT6Tj8n
6wOfg9g8xWhL/08QxxHl5obUPfSJOXCDc85qoqHOPQ7FYElIk4OWZ9ylGdZW
YQz7OFAY1dHRbijkfAc2RFcz3cOqJRI4QkuWp2OOnaCtf5+koRf32HEh5HAl
19SzTrnN0emztuDxb5fiQC5jmdc6SbRZEvp0KhhX/jc3E81dV5ABE82V3/Rs
lSjlnVmUKJPR7U/mLKPQi2UoohwqtdlTgW5flU+i71sZaH6AlMGDG568nya1
i4sjPwxvenalCUUx4rlib74XyOCl4j2rRbDt2ah81mXijON/P6wGsBj6oKvF
JAIx2jHLenhlcdP6P0MfCpKWHHby9/99xVw6nPlotbngGGvOzN/cIifeeF6M
oX9aare648mWDxLBaN9DSSNdxM9v/JsWooqjGMRkc6JH/H4zXn8+NnVEuzXU
tij3mcXmO+HR38NiJzf9aqe2wYxDJqd7fVUAk6T05Lq2Kk9k1Anxgv03L2sl
glovBx5sEKoDH7kVheBkVTeLA9BzggPQtJ7YXGXEpiob++BAqpNVccMecGzJ
nKzRSTyw9iOMlbpkrA8zPjwyEhu3gcpRiiyhyUScRWb2nicPfskxQvk1w8zE
72T1b21RSkDXRawqAAgigNxNgIzmcpbSwEK7MY70fAN2sgfKJETbprYqwTzz
cF2K8VGq25GbQTqnPX009MidJfi0O1mq/0+BCLWMYtrXKc5MDW+dED9C3Zqm
LkHSGPK3HFE5Knb1wTPQQ13K7mgAbVir/p5zQ9rGdI95vS4A1KOipeopkurQ
afMTsk+RSZFmWv6UMwwPQCivgNAUPupVlk3HOC8R14MS92k6Yto4FfKsz85o
CJnlOQuiImUcDaQv7HV2GGTkpFVbXtDC2KOO3K+Wpy4Qz1/VmvllyzZzT33m
hEXsRMdAygAfUyZKJDXi8FnPK8a592ZEDMWwLIlSySekui/UKjaCwDp9FoEf
8xBe+niE7+HAtTxJj5lAmw+I+Hr1e5/5uXoA4Qe7tt6Kw48lk+lqJr5+pWLg
bP+uzB9Ch+G7PV7uy7uQmSwD1SZKvmQFon/SDeIG28sVCflKDL4NgIKrHMDL
nUtT5mjNk/I/aLD5uP1dUHv97Rd3Q04i8LWdDM+yQcgNQORdT3eJq+UUwjOz
Iryy0EiRDk938v6Jthn+9pSLY3VGHF95kqjWhBXqYiVUVPKQYHNZqRyU5og7
1U4cZeopIcT4c643H1zTL2mSZneE3n6x8wFeYcrs+Dg7Ifvx3UnUXGEgZpL7
sU5v3Sw9aeVDnOJEbs50y7WlFEf9pGNjoT1Js31H9OQlBp2W983Gn6RgBxXr
OTpclt2czfzLDy609ZV3i9BIUthR0MOmnv8wCD0viQULLUCNQ5z7ZSGawTWj
Jx9BwlVqOX2Z5oJiSf9vNN7GCa+5kQ07oUYjnJEKcBlxBW29kbUyzEX5Hoxf
eWwclWbmwoT6G/dvpiSGgobeDshi/xVoYkYZotUpIw0gdXA29L83gjh0qhH0
dSaKgOaiCDUQ1zNgpmvEEJfdPrKwjWkT2SQR4Ue/PjBAj07OCUU8+O7az22W
tyGAZcWiiggO3X+DiTKexi95ghtiKK3+hl5JbuMzOF3fJfFyzIx6crqB4ime
0Ytkssb174/H+npKpR167rvnY3kmH8+n4LSjlqPGvTSbDeFdrTWaSohTN0j9
4W6hGzHSNcHTid66kpT6SEw99aQTZglnAY3AcZAoZ2iyJvOOmt9Wvdaos9DF
4m3H5+PnxUU6Ig1MxLsqmO3md2382hZSWDekkvPKlxNQEv+a2+Fljyh9r0Jt
oQC9z76LL0CdSwMZ9VK2k1z/Hig4BayzMIFwOiRatY6kN23KV9dfwCFDfBAC
Nb2uCgrL6xikn1ecKWue/5jqNtJZwVP1Mbt6kip0uHZ+ff1QK64bl3NnEiVZ
GnaN2qormu6UkddN906ZYZOI+HvhObDrKmE3HpEqmyjipHu54ASrFyZCVeOt
K0Adi2EDvgfrwHH7r9j6gpjvbjRbTs3ZQwF/+BbRT+LtszoDrGRrvsKlCDnO
iP6aag6M6z2kORNb27CyCS8rkmkBScva5Fb8bDlfE97HamNIVR1PhhyIsQXK
tv3lj1ys6cfMimGFvCHsr35SCB/deN9uFhCtd+QmUTH9o+Z2tCVAbC102Ypp
mN6nDvOyAMnixOOuZaNuo10LXXZMa6Dw+Jba8jvl9owLdgca/V3zFsUg+KDU
OzcDtUC1Sb5lh6zSWi87JyFMyw2mM2yHTGEb3RqRP9mWDwqztThYXr99qhYQ
ArfkOm62qYpPf96eEyxwWFrJujNX6htQpJIVI0TomkV4KFl+8oKOD4XfhqwN
o64v7N/fL0rNdnDiC9JxllG5cMPf9NlQP0SmkcEhISRtS7AaaBQnlw5QbB+n
KOxqFPlbcljIwXCbHTmHyAd1gw+On9u78gdf4LKIi7h4O7x9ljwm0OpXRQo0
EqEN0SyYlQz3/pX8md1Qtl0cLDX3gZyb9wjgEafx2BQSnAgAt9DL8e5N/Fkk
sZ1HPqdNSWdNBqo9p7/46zzgHopcK7paTyi5VE8w0VQJx+bZFSIIQAmR2Vg8
bOdQBRUWtpd0LabGCSSKv+iu2xq+t13POlvovL7bag9rD6ya6seJeeTQhkQM
n11uglD7OKGeu4pd18R+K9vh92wLi5itOQS1yEzNgyad86MAL+F9D4yTwU7H
q6XpZKvtMU5wD93U+YySUQZ8U7DtCOExjOkKG8yHuRHfD1kW85L8qy0xPQzZ
hw1oEKe+xlkOTGChiIIwGj8aS3KJsRdZg449Vkt52dXauMF74Gw17yJ9MIdb
lQ12SHFYNF9TqC/2fKCyWOEkKF2ZH/3JRkf8Eqy9mMqdbjcCKR1NyL3UOUJd
SEjLIpUpxUeX1dXTDq+tV06mQVenmdtM04qJHyET+lLnL58NgXiBTplgahU9
wpYHAsGBYR40nYCHxwNa6gEf07MlXH9TCcOZL4Al8sGX+586mZ44j1nz7ni3
tDvEHRRXl6RRoiGk1HmsmGpeX5N/gDJyaLjULLgYw6cQoaT+wg1N/vlzsNyQ
cLj8iSPwseBD274xge+xiOJ6/aCPmAxJ4hRI2kHtnXrk3XIahVuzqTN70eF0
OgLnhpusGaTZcE83omLsJAUYxGFa/acMGwpLbQiSinlG2rBFSPeFixahYyhA
FXQDQMTF37jTyxEOfk3/YmpPkayyj5PzNS0RTpU/RiC9ZwyR6tAQa6QeGKOX
m2WDhxP9NBFcK9TPe572xiTLABOrq1WbEbzEsrcwa2yJuokXoTtQxnwS2/Of
6Xrh08ab4twJ3up70GEpgSnOPZNvNlXpQwjulfix8wjNb8UniUgLNRtoUibT
rMpolnSg/Fk+P2Zz6tzrdaXXICyzxdNAc4jNxoOOiyNm0/whZZOtkuuShiQv
NKETh5THKbyGgVhaYOIS/NYfMvg/1uXZAmjaKsrHwflP6Wv1HOaTbHsBPy9+
KpjCAzxwAy8QpRdAyhArjE204PYoVmauJTcFOgitlGtcArvJm+DGxBdamw6u
Z1Rq4/3NkZWNii7qxrO+axTotnteE0etvgd/cSU+P7Y44hft8YEHfJDXF5b/
tT6Me3nqH9ucj1g8owexiZmNtuBiK7Vh8zJXBGKq6ORfim9BBUolAnUqUOXc
hzcq/zqSTlkkggqmr14NDssUR1Di3n4mu3aabVBXoQ6q/AOyHbBl3ufXvkZ/
3bmbqjBw3m04oL8Gso9StKFaCyyhxQr3skrDumxeafni+6bmtEipOJrjQFPN
QpsXKMWw/akLcbQbcOHA8eRkHMRQ38DW2AJcu6JUv/S14U2EnNhYZOoXLeeB
VaE263LBfF754pUJReyQj+NPbLeURz+zWYbpVI4Nllsdvxzt+JS6DzvLRUQ0
TmeEzA5xqcmRURZyE1yZSeQaogKMOcSuCfJQHPwMzA+dXZW5JiTycVF9rD+O
SpVNaoZmYJvvFL5be/P/dlVFFWYKYlmywbzyxcHTc1P5UeGayZ7ZLcOio9Oe
YoDHuXzubvq4ibRtv6jo164Pj6M5fPJ7gOBGNRvFRb4o/c0WjyV0wy/cT/rI
af6Sc7Nf1ufAu+KIsbv7LxCsN4SmeXHEFoJTrsJdFjSauPN05emvF3yUxYkk
kSJI/XxbR6rl/80A30oKBaUlnLFBMNJZEE+fFJrMIBiO0zWxcd0iDLAVfy3k
hUCZPOcdOhzytZKp0s5kuIb68AP5yuPkBdpirQM93uEp9AbxY4u6Y0naUzuD
JI1sLfNXLDGvlsza7ElsTcVqW/TtyNAZ53hMFzDiYB7Bqt2056Ce6FlIyW34
hFnUms9oozDAkg7OM/lS5c6HgDB4wxQnyy1b2SL8JCp1tBybS2ehcPofRRqo
X/rFpvqwwATHZVheaSnXz75EDlt2L9vyZy2URJGiwD4lJXaaUf4sOP7UGl+z
bDqBM5uACb/E5TW/71DROb/R+J25Shq/keOmEfotlUgdAyOta7NA8FnaMS63
q+3vUzsZA+k/s6xBPxquR2OYdsddlW+XmzISN8iJA0h1UvTCm4RX/02MORwn
nGMIPQpvs94IM6ud0ER8FELj42ghqfLCjt5nujjjz9lMcffzo0V5Xb8ynGi0
NNzmkJl736TsrZr5yzs1NeM8P2zZ6jWkOvagQx/zUzGBr9zrIluiaSVeL26N
w+yMVJMp5dJdpgaObt9MOnEdxM6GJuT8IiH6A9fQWalgBe3ayG4PM99AdCjN
mgPfW52kAIO6xX79UOs+kW35wszAXcEdOY1w20ZrWAg2EaAxaQH4oK0TR8X6
cZYo5DHeQU9ODRcEVyc2uv/EcZLg8QSwxUVGL14xrD8jp6F0Nj/SUeZ+fk4j
xMjV2NyHTJrWKN5pwkoeigIxxbkVw/JLONj7bS4inF3LKH71Wt75bYNkgQjd
/TD37IsiKXevBRoprwcbzQeeCk9vZPnl9qJ/oSC2YuxzqjYPjQ/aT6Wsfxi/
Bz7RtqqYtrt4V+KmG9Pt4OKt17vI+WNfVZfAml8jDGSU4x8WTRdm2RB2HGfD
NWh2ncoLpoOOKo5AdDsTXB0/rcReS/qvr6XEs1GVG59y6dL6bUREy/fOZ9QH
wKIshXgNbPVrtpSTiYBBUf+85PCdi4gMYV+wgtgqJOsl6CROJMz98iosaxdd
aPEgEovmabKYRxMvKANh/da4sHOxee2DV1O/vcOp9q3TgT0tGekC3EfLVrEo
I+SIAeh/Tz7d3UGpHs/TuUT+ulomNfZbx7X5krsVCPC0k3MnEnRA/TBEY7US
GTYK6JxjIMXIEo85Pa0i4kwsP/lqAwbjZWSVlIAPsXqGZfzndyVeRj+GXc38
3Xuk+5Mg4lK5j/F22URAU9yORZettsxvL02TvvF941/IsG/IacMHocIFbEGK
7SwJ5/R0gvAh6fdLYMSoZjqDHx9zygPGhldlU07sTapz8UaVmG63mj8hJyx5
v7AO9XIiEAEBgAMLtfgTaMo2lovrQik8Ikk3DS3uFFw71A8UCN8ac9fhFwH8
W0lCiiH/ABWs/aE7INnZ20Dy+Xxl+7QwU2jCvQSG2mMBqg682aDDoe18lEiE
47UBHtAz08NDI+R7AkBILhhAsrM9JWC8bEC/CWC/YRcEZ7CEUawOj+EMeCkR
FGwxtPdolg3x7EI2MBXVOWD2UTzJScdyzvtPIY7tjkKD02aAOpVRi/eMPgL/
TPeKNBiKFdAdD1PuCCGesI9OMUxwVSVHxEVlCfJzhHwd/KFqCRjAHMabivat
ODONo0vs9UAOJo20+/LD+h4BTG5FdmwwSDlE/SgjWynKJQkxke5HXC/PHYeQ
hjLdGxtQKMqoV4I7FL7cVErC8C9U0IIQoj57fibGLcThkfJ4js8RSBKYjQU1
s6rkf3AElJa00p13N33MuOCOlFcckS132S5bdZSBO8pSCvFdh4/vhOVUI0iv
hhg2QbREc1NjWK0IjNtB8tuSlQ1B6rYAVbL4oYi1RIUO//FCBHZerutN+f4N
86dDV6KZ10lkFwlx1Q/DQ6xUnBSErypuaioBREQTfXcVhl4xY+mEswPXvmYj
sQzhanyPwCG1j7XSQxo4olvR2AUr0iG7K+16rOVc2B1YSPe9FAzJke9T7DT4
+i5Dm5oL9iJSGtyrpBtzgmgwobctdegfuQvSiSHMX7S2So4FbpczNIt0h42B
WU159h6SpOv1Vcw0znk6geYmQg9TT5JzZCYkdj5Y+piCFqKL6bwrK4/1TwjQ
fcHksv9kpqLk9s6r/qRB0VGMXN/O6AFU+PQZhGbk2+dzIEmve2MsBo4ZbxaG
yJIoC6vvPDLNDo2Zr1GVvasHVKMyUYdYt8Kg+Sq7mCgip3jHomWVKdk3hCV5
mxWre7rPxVMa9bcRhAgg2fwrZljxn8tQJD+9O3TfT2md2XXbcEj+tAAdTwFl
XE6kcBya0DRA0D+BLHbJUuJUCmtCGBXJ3kiLq3PfMFWYraQSnsQiScBYFzO7
MwCmi4m5ZLvylkDapZRd9/1zc6ZCUA9ypRqMtkrsWpGEKJsnm3YPt3hBTi11
F7ujdPOMcyXoIpP7k6ZZjKiugghyDEgavEUfZhPhpZ5Bcwo8okjYnby6ehZb
n6w7MIgGddA+n8Mw1Wq/TWIrYUgset5Hr5aqsvsLhXoYiJER1IGA+FnYktfC
+D8/NDIX0Nz+8CsuV0XPzKi3S+6VZ9U3+QbWPMjGvXHtLbX8gqUHTnJYfQkS
l9TTH3ESy47hNNDgVDr49Ywwx587S1rNai90rcV44Rm+CWF9idtjBgcfFFmt
DnyD+dUpir/e1O2MHoNBVWmd86yA+10jEZt9uwoubhwOoem2rdolpexJ758L
8miZr8FVsBcXo3aVc3axHAmjf+qdKg9oc2iXnOFfj+RAgDvnhHPe+C6GnCLv
zlITb2dUDcGIXNLkB1PugEajsvyNr3Gk9lZnTBV+g0sw58JgDymc+MVF3YKn
sqfWPmJ5ELUGt3Ei87fdN/KUk/7VmMdNgTCbXygjBJsCZVMdNbU9U1m3v8BH
wM1oUp9oIML21+3YDH6+hIPJ5XGUdvSJn923c2VG4KSXsMdItxbxIj9jdY/K
9PQzqw+kejY+qrdFJIUWNdwKrf05uOvMJV6UlpT3FgzUygZdT2jw+vgmwccx
WPnOQGhAloFsHNOPUbih9FkMclknHFSICs9L4di7r6l+MGwqR98Zd81sYyEi
fBjjfxL+KlcByQpM0PMvKUEEh1fYYFLG4COUlEeXDUesrsHHfU81vJOmBaT4
sPOlX+7ioriFRPJMcHsHlSke7hGENyA7vv/0/dpKe2jfvE7jjlqOLB3HT47D
bRvQippQhLKVXcu0HWKwMr8ytZ8yIBay7ozwlF2c3GMUCpDpAHZFwNxRGk4h
wl6ETe6FRHGJJ5LAeXYa//nnXnIfjAg8NVjcT8jkgLs4VJU9j55jmvQWWi9D
tVLXP3Ji3qK7dbdJW3azrEijxNHGwLqoxnxO7syGyYS/MkRDPXcweN51nR83
O9fW5SDkvC7wUPBVQKMZJZHKwfoufbCiH5qHtPjgQnqg4DHAeY+33+5HdX2g
1jRdRT30ApGjrCXNmhy1wNvxmbQwaVjz+sLk92amen4tjUbM2Lbb4m0LtjYj
p+En6kYck4+sJXQBFcipTAfhBrpjvOOC73fGZ4QWXJKjaoUB0LcBkanT4wiL
SpiicdoOx9asEGZe5KM56Es25IaFFiX47obgK5CGMLiHxuIi/eHL0hrIbiXt
OTeW517gtQuwWC5v6qlHjTKrK9HDJ9httjEWquk1AmGoLJ0y1TItPHjqEhrs
AWHyy8gIyy4B2oi9iWvYqHGWnVm/aI68BNA3cIFPnHOdLkQVWQADSKMlktku
U2mJL2ynmbVeDGKnUn4vYR5aDd6yoOmqGg+bJfNQoG0Z0OnBqqZ8BaeSzxNH
IcCy5o4Zwmnd5dz+SKU/b/C9vFFb34bvNFxcPkN9mGSzdhTr4ew7clOEbDuB
lCWMxe/28M4MSZEzj6pllEe6M++NbDLSyJWRWfYWowD+v6CpS7z9xNEoUlRd
dGM4LZ7Rcuzfs6/f7tCAOmA89qG4EwA+4Furk0aG7qcL8duhcJbOJ+zKSK4g
ZgVJQAw1C2sDc7+KXFdC6/AkhG2bED8hmgLStEg/xjwVvQYDF3MGGL6niM4o
DEGvT2DSDwJRDYf9Ju65xat5R6Yh9NqRXGwR8gLkNLsH+khRv9OKHzSdo2hL
mGagAM3LWmarTmzUljdR6r1OHWQMHV98+E+r8IsAog5reHLNIsE15yiwsRzj
GPrp5b2kDyvJN970/UqoPtRUHntwsHKpa6F5h7ke5qbwWJ4fH/W58ym5EOQl
UglwDCQ8SEKhG9uiLBUoqEXOH7e5KiENNsmObHef9MAIEVo7tglTjTQkL1fI
QBNBSVw9ILpKWra37BWw3O/F8oVS8T3A2AMtr9gGUJnJGfPFIeGHfCGd4yN9
mJpPYzXbHD8TLWHXhEIoaT6plwqdsivbEJe8fdalpEvt9yp4mOeZKQm3/p51
2E+eLXWlPCQtR3Y7SZ14ebeNl83BM7hjC5r+r+iIdGvcuZBY4ab42IUf//8T
Dt0JkywTkFunqyFp7lXAMgysXoDDUCKU8e4FVcLeHNTfwYvyVv6alZa1/glp
DP9eOWq2jPGQG5lOgeERsJrzzcNHChLuSbPTnc99bk8b32t7nigGzkwCoFfD
b2DHbj01Hp7TbmOrKSznWxaBLdXvhmwO41UyyXKri2B5Fy7Ilf+stIhmxcod
xQtLqaf5s2LePF3fwYG/NFHfZJ7kDD6JPYitdQ65xdOP3CmeWzKMLNoF53pB
91suiLOzv3uDq9JLcv5aRaVtmqz8jt6y6VV2E3g3+Y71ydFhzjwZyiWOKF0m
3yR4KRnZYKuCSv0eHk0REwHbG5j2U9Rro6cCNZCz2UQ9hzIFmivnf5Z6byY0
NXvLM06l00dSy/ItqQfQDBqslh7OIy2wKSahOemxWMoTWqldCKqtIXzt+z0l
asalzUQyU7ueQqEhl+yUeW2cbCuD2THBgZ7dOpRrhs5A340zwtRDeBMKSGiK
QOkDdMvDND0wdh5cKmgbgRJvI7xbbssUvZRrOfCXk/myKFaHhKde05GIKUR9
nD7ITUOhfoxGrUJcH0EZ2wMpSQlIKHZoB9/COKcd4AnNu3wv/fhQ/Aze1aXL
VfGgljMuZlFcdA6/fkpxyahSWkIt10GQ5tpky5ywUV+KOFIhhnXJ400mmSbI
eTQkTChzGS1bxh5sdXCH+Z+QbXiHp9hlVaehRFd93DvbK/GzAuOFWD6neZR2
WP/lBDbM4nxAY5hvL2KyP3129l4cEtsdw6EAaJc79Gh32158YNK0H2JCeJ6l
wSI/PiPHE9A9BQD+5zRYJkdkJGKiWCtUDghoJ+Rsc61OKrbGM0qymCYdEFEZ
PEIN7rLO2oEJoH9tUoC4dnw6feCOrTzVrn9SeAq/CDye4kVyK+GJ/U0nzQJJ
oA+0zJbx4KEzgnR5ti7n5wYcOwE3JAsU3EvilnrXOLXBFcoEqOXF4uYJJ8zG
xZ0QrETrQJhB+OxEIHx/E5yKg97oRfpnsiEvIQf70tISus4sRgYvCrChauRb
puzmyyBxy36NliJhSkGfc/FfXJYwc3mTNT6i0DSu4KQYko9IRSzSq83j1PIP
lfl+VZGfjfT/Kq6znTZCkJIfduv8Jg+ge7w6uLi+0xNy3MgntUKq/UB/UHUa
4hdWjrSahS+kWeGfQPc+rmUKXNYiDtm2CSwiRxVRMMuL5XftSOKJperGwDaF
DPRIFrTvUywAQJ+XPitLjt+23NIrr1vJyucAM7uRWb4X0JsdHZtJorf8pIOg
6hywqH1qkPlpr7lNKt236ZdFkA8A1Bi0/aMsvWjielndDLCdv3A2mu86rEgE
+ReSTKttCKYeJ5ocL49UdHv6aM4M3Bs/Wi0lHY+yKuk8tXyJEa2b75Svbxec
jMfPQM1fodUJlk3ezSEKg14VWGAlnSxyczUhljfChAQAh11iJUXiOzJaBDuO
Xyd+BOsnE3extyO22y32Eb80ydQpVOhl2BvHa+cW5XiFGdQ5/FpSGMgN3Ca5
yN3OhEVdEQTvORjTfvIDMWEbkixSJl/G3CtwFjERXe1B7vNKnRB9DhrPnogr
EpUAMVktLDq5QIwIBa29Ok1XF5lTK+qF58z6yxjSWLBVUVkybLNlg+rkRZFb
6LdHwvLpyH9HuWVP3o+tY4sTsiiK4lzqyObEL9gtHJNZjVJL0eO7HGjQM0dI
/q4GWKgoFk8DOoPzTJmVw7zoGyXfH9xkdhkzEQ6BT+OlXW0aRMDk4/971JDQ
bxX+L5DpHvAMnysPPFGQVssnthCKt32vzK2NtnVScDFtXaKK3EndTtQjx8Ry
HjgIBxPxd0c9fmyyqL3GskJ6j9MOfZdEgg8oHnlm5ZudHQZ0/u6amuYMN1UZ
FPsNUbhca5IjspbfUGuMqw84U35eGRtAh37t0t+nOmxhrKarwAR73qw6tv/2
2xFmGGmWoqxztKabRu7hUTxzI0gQJ5uIRZHlwg9lnYUHyrbgY/APvk9sIxHk
zQMfxuQqVTk156wJEaK8RJfGsg7OjdwMaX2nBURqVULdc23oDc87LNrBtw/q
qqtqZK4/qsmoFSewdtpLGoXehABV9LCea5GY7eYTtmKxz3bhjlbohXiO4cdw
VPXa5CnbIPpp4M7mHHQHcFlKwxYpEBREWhqd56Ob16en2VAtypKxDZi9T8u5
9oRNAFejjphxSIycJ2H+SfKpxC9FLp7p9faeXHRXusxd2GambH7jvJ5se4BA
gp7CgxzxtYNGVFh/430J9fKv68scodwUkvB3poHfj7UtjGoi6kcxJRKCmLSO
cJgzOMUjeRn8b6fuVZ+We9VF6Eb/4M0BpT3pbLGvvx8uxXCE94Wz26ZY+ase
FBF8iApUHJBP8SYZcudtKan7DNvCWgyJHiktTOWpAd76nF/lPNuMm2Fl/qNs
KxrQxZOC+LwEcsSRMpaOhVfFF5Ooyf0cHJwx2ycrmYZ+UUvnPjzKtuRnVzyv
/40zHTw/xz1blf/yJwHibEgiybiNOabcPXpchg/TwGlckdFedBkeDs76z+C5
sWUlb4WzszaFH4e1FnuIa3kkLNpsveb63A4f0qLh4ypFB6RTWU1R5MftdaVb
5aQgp7Hovp3/dKP7ge0f7kaFX19maCR15LNG4GKzm4R/biF1lee+CFBSLgeZ
vrcS//2IEruDR9/R5VKKc8BB8F0ivGL334hCrcbPu/qkbvRMNwAZfHJWh5V7
YD65VH/yL8eVcXPNvmBmwwrq1p6IMeVqY8Ksmw4hkvegJP4fb0q3jUfxTqDx
1Qt0Knu3Juw7oW4QHeAPkNUQLO4wrK0ZoiOUsAZFMacoQkr+/mjXx4izoWBY
usxQuSQUVEIRhEAv+PQMD8B+YtOzrjPvE1Bzs55PddljR/tEIv2AWCoiX9/8
y4Wo1+T/oDtZK/ysQXC6M2ox1cuoYUWjjjYF/g7ccnbqXAev3JZMW/jfMqrW
qkgnAeRPpJwOZtopq6ayl0nuNSj4pZA2DIibWhEy5zsv6cUe8fPIgpNYtJn6
yfn2lnF78Gv227Ri+4p113jTkw1Ufs7kbmiXrzLdIrTLhVkLp4NQ92wKuEe4
ObXCMdQPGEgQuPq8SfC8c/9FgqzEmiplm0sx/w4w/AFQhBS+P/EcDcrPVsT2
aTLkSUZB3bmArJEsU/qycze6iV6Qa3PoOEgjyDDTVGJwU8zcNeqUvMbkHHnG
1gUWVQn2cQqIWbJK57Sv3j2vt8dEuoS9o3a3gEEJ5vIef68J7C7+RaBoryRS
jbw6FNGEaziXQt2UYngeW/Voeq0pJ6SJRRr6mhWyQvA/1w1TiPmtqQj2T+Hu
224nFmyKOxTQu4i2EdwiAy/L1ofGHRgPDLuE8N3g+UwbyFqppOYlseo+d4I9
kYgnOiweXkkIDfivOfq2wvXlpn+p4McpDPvsleLmf2vOMGsYKz42+eVTMZi9
ZA+YcPx6fL2DHl60Jq4/ALyNirBQIRMNfRYkProhAV76fybV3wwmWct7LM0X
Xa1ZFhHSSVYBuqR4pwagQicoTP1sigOcrnWTcaksS+Xrz4vCdnKxN3rcnH8F
l8KXpviIFpprI7ZLJ9hfG9MJgEMD4n7xJwdZOixb5Nu19KgvRbGP+BvF2+3n
t6TS60e5BLao3RSmdWZoXpOIKWs8+gxIvLJgLfP02bpcH2sHbU34X6YmDKi/
na8XGfV93WemJvesUVs7FWsUtTPQ+O9ehBNxPP3Af6cvpYLD2qeS4k8ncAxa
o4P/S3yHpCgYfdRrvjH97ocCvRsWwbKaiVVaEpgJc2oEdNLkw0mP5UgoD6A+
kIqNcs/kdv0zSs1zKa2oYejGRP0u9LzLNY3WpHf+TBbPwKIn3FD9Gambcj/2
4L1uEGUKn6fRlXbKaugkwvDTFvYyrJpGQtlDNn9o1m2KDQpI2pkiR57Vhmyr
50YW3CV3ucL4HKlH8RDSwhbT0azDPGcF5arIsyWlUO9yd1NOoTf5XYZi5/2h
N3T8gnvo1bNesiIRloXfsDDZ3RftqRvVwzuIwtN+8UOSZT5oz5zyw7hwDLn4
zxS344Z4melkGyeJU3hMPQ/4SA0V7SFmtToepwP+FzuY+aW/Zr6+UN2Dmx1L
pHy2cQznrm7uXXMrPG4i/0hDnRViJjHrYEW/KlILnctsZPIT8v+Q9s0kJHQw
F9HyfUqLOhNNgNVkGISTW11xED48yUcf+WjPPXB/UJYmIQRSxqj23k+uiCf8
QhtI29ydWLEUsKn8HnzwjIH073W5oHm1GbqIWAJ6WNUgVuPBHFheKjMNUmJG
yFADgh2AW3yBl8K8Zv3ga0OaOBbD0QRvWHeon/Gdf+gwBE+RpXpNINfwLKJ7
FNRzakYG6xh3jxcWq03omNd/fDcRaEZJPCiwhNUGb67QGZUdyHzH6nfmBtse
dNozEfrsX3hDZ8BrHe5wI6cKHYuXzUb60ZfHYFi76JQ51vCtM5BvjzXflwiS
jGVnYxJG/5Ahyx/CrlmRYvxmx3jsCheovvOMD1sS9qDO+B5zGsvYjyROIkG/
v3PiT/lSEa0/4GxK3Spyq9bgNMRuLaa5ROKN4XvtYsb566s2CqSX4gKbzGJS
OuhBux9sVHe4aZU9Qv9d55u8DF5/FC06dt/Q68x7Kkm7wh7kgzXSngY9uqyK
bnLDyzF8rt/yYuyTJO1ApNQk2VdRxVmTfDYmGqmpRW8gmMBs4xo6SeDqbV1t
ZICZUhsWNHNEN7WB99Qg8CuA1Ef+FBEWaoUnlTItCWoUYts2oMhIeQjou4Sq
kxeYS76S6spz/+2ott7oYxyyytP9Q2mSRg3s12bbNXsLMqd9FPVVQDjpfcg1
yvELIp3ftYLuPb3sHS/fldUBxj4cX/DK7BIolifTF/OylmXZZTRrMe/yrGis
azmxHUgVBx1qvgcc37NhZDc38s4ipdw4YBGVjxUL36D4oBm3QEg0CHO19SNH
gjzvXt6lYWGnFhpscHenjZGy7RWGbeAQTBgEvWAl29JU3J4j3GAY8jBT2dtX
n39IE3gLAfFTco7OSU6deyzHMqbyLyE9ZYbTwKeTRxiVFkQKCDqdMDAzyQXi
fjV3dqJT7NTVX8gXwP3thcEOs+7Eps0qHMaSyH8TI8OpF8uCJNmDMU5RM/4g
T1DVHt+5jNSapm/6PxE5i45jmRnedsYzbYP6IR5GnDXE6EBQiFc5yKjF8X7s
Z/S8ptlvfgnY7tvjcN1l2CoUFt0febSY/6XRBdluoAiPfm9sl2U5liIsK7ju
Haqffa6jSfUWzlU4I48jjofOR8NC34Of4Tu3pTPmssqir60qjtPA228BNJxe
9bzmFBVf+b7Kobs9i+6mwNCzuhkW0ftBHet9/KxitsPffehVmnGIyfq6Db31
H6fYczytaBHw79p+0xxNdkBOCUZOylodLiGp9h+ohI2GoYjgCo1PSvuEF7BL
BubbtjpNqI8rPnbzyN6BvXZAq/ldmB4Ea59envrsbOToHcMHKMCsc0ea5W8h
FOlKoTz0/R0KbJ86G3Ffv3628r7YvdoAy3joKwZecb2KjBsM67pOmD+QuYtI
euZLXHujyVnU+JeD8ehISFQJaR1voa2MtNvzsi59rv/TRQUA9/QnW9SfW9kS
MwRZ1s1o9jxccCbeqhoohTHcbNaAR/tFQyDkRsmnOzWHWkNqH5OWiJ24td2O
/gWA4cVccFOn8w/MKf2tt9JGwlJD7dQ1NUsE6cTYQyUOoTts8Q77FItfjoC5
ZbSTGnPssDu1hF1cxRVBdoMBWaxXPee60uF7DzxdHBDfaTIFbI4/Pf5JE6dJ
WmO/Haf1hZzZkkYnMfEuLa9NZciAoJZc/vaYjEqorcdwduvd3x+WCJsve38f
oRTh+aBmg3WN+VxpjSVKaSe2v5/NJpzDhEkGeYB4tTYENojzvLgCRvLu0ouR
IDcDLXeDFzRTVBzqMYSDmosscpx8m+W1j/aF2GXQZbMBLika+EY4i5P2pooK
fWLkRFa8jbzxb9EthZi/rSWxthZGnCGOAvoKeDl8OD6PZdn5HVsik5APDJnY
Mz1mP8eXcLOC5szBlkZ3ft4APwDYhhzinne+j9saqrL3BBw47Li2M5u545DS
StYzopO51mIz0opA0DYq9AxE8Jo5L4van03UrESMPJflM9AAjM81IDW49u8y
b2limqGyAXfywZ8PfXmbAY55NsGzdlNJ1PWhw6CjZyOwFt7bX8zXUBoYI3yx
b+nZafYJcdLdAbYNXOugi0EvXItgHpROXstYCvanXwdVhxgcQnbWMfoQnUXN
s0zon0MEAuiwrNZvyYodMZqcT7wIpasqQXrQ0L3rqgiS2eOAWKcqGqsa4S4n
3KYJuGp8P20oTDf5fL+Pg65RWYBDwV/ZBicjzPO5rK8481EY6RrSFoZbXAcr
WrMQX2H+kGzgFS0skqDl9+uoESbTZO5iFRcH7QRj3KZnrTjBJSgyRayG9k6Z
PXQlLjk3flTfz08MxdcQWxHXCH+FROXisQJeCNBTkr6uNLSuCewEzcdi2fIx
ZcG3kU9qNT0MeIDfMLAORBTuZbz0oHfItoVxX7/eIUVsEhqTVYovgTTepBI4
uj1zXM9et2jwkRxJ5DOMsUim1Zctfg4Ugn1OFuFqGP7ALj2fVVl+7ytZuUZY
WSyK2fy/DBheNfDCxR3W1PA76NPtz5MXYZ8HDm2zEAkM6O29Jeh4k8THP4Cd
jeN8GYaXn3IOfDN6vg22VQT6YKzjES4F+MKhANEm0ZLI+dDQMKBYYXuIp9l2
pFfRy0AfZl0doI7aq7svD2KGvlE95vgxHGutcaahLXzTdAy0J5Z453Ys/Lv7
Nef724FzYcFuY0Anw3776RPEXoPrx6fDOvvrmO0Lp+yAJ0ayzuPXCrFSTNZ2
P8WrWMWHwFRgWgnFOxoB+21yw+BNWFq577L/GwLFfX8XI6vZzS/JOTQEKbVb
lt/PSbQTbXCa8kL3uxEy33RWtnYerJvhFD3ubhETsg/OYS20DW+kS07e+509
U3+lmy/lNaqtcF/4ezj3l2GNINRiFc2IGObf9gbRZ5jzrfWngt9bi6iCTujH
TAGtd4ZDL3ZowXa4Wh/97zvmlIvCZ3TOgJ4n70UaF4cFdiDN6mbJyuRTbZse
pK9xr7Mbk0Vrl7crpHhNoP1CwtdQvzL08M84C9nVfnnj8F+es4A0N81OM3kV
Mp7BSdTMjaDAJs8zRPl9m4YwU34J4QVSqo5oK8HsuhEpi+0OGDS24CRhnbIV
hotT4i5LKW8HAL67NXlmTxw0y42ytMk2LTDIamZewnfwf7yVd78WhsDt7XBi
MSseruGnp9LNYCIyaxa+vArvOk3LwTeWhVibDha1mvlchoYxqyIPXWPO4LdK
iaRtaNCQxmGiI2XLU35+VDpVJARqTAy82YtJQdnWDb5Xgj4jRWRBlJ8fiWF6
/dFtZ4jvTAwqkW9qhfBVlR9e54wgzgGToPEwsUAmEVKsIMiw1OCTzKmfe3Ni
91/k35UO5cR8QWnWpmwkah29Zx7fNxy9UC2uZ3OuKjpONZFtZwJ8Ls1RB1bX
2h/N6HpBLOWIawsXZLBlRrwvlcd4+Ca5EXHJ6Zr75vtB9s6It0xoOXXS1m5X
yORVtkb59HdvL92DqfAmxYK33Vwmx+Iia8i69/xye4Lj/O0TIjNzRy0GTfDo
7LbeIGa+Tw2RyF9JmM2z0WFIP6X03BgU63E3qehJFS1WIriqXBpbOjqGqY+V
rpNKCWneCaZZ70lhxct4eJxKVGvICUC8icxRP++XtD65ZLztvJvXP1D7vcCA
Ca0s/pjlUizgeTLQ31pQrfs8jqx5RfOsbAUg2vevjycjIWXIX41MNXZeaSqr
0pxoP4HcELT+2LtZOMv/Q+6/2bsINPHVlLNhOMZ0aD0bztPLv/Xlfm55vPLw
oMIr44tv9Jo4J9/XtO9E5U1fWK1XQvwd9IC1xXfk+x1QaTNbvIuraPqvTJlF
qjS1YV3eGMAtFshtDF9f1+E56jWL/XbKVpCi3LVOMRpH86ldHLwU4+l7MmWr
oZlIldik7hTF6z8M3/jKJuIyBqUIE+Us/OCSnbAL93hAzvaGkyjTlZvF/dbF
keQhGeNjFXjkGWNLTpx1nd5zO2JLmYbAfwePE88ond3s8oryd4p2EGlhPwLm
pZ6zfqFu9aqp9eSvSee3+UuOmK3KKzUx8BGaylIbcL/tQY7s/zGet1KhddZD
tW/9ZBYC33Ym/hUqG/vAE4uCA7PrbuGdTkFOnb/4EQ5oDsWvjsFquTb2MxJJ
2v3FcRh0MKXr1D7uOcfXcPqlw2dIjz452MurYK9DRJ1V4j/wwS2ExXKihb1n
coMxUPA7gvZBQpExwDoM6iClV64YVkCYb3JpgWyZ7mHXpXXQ/1b9gG+Z051M
7jdLUiqv8C1ywoSZRZGJ6hXttcVTVIG7NJp084mrQlF2Bxe8AEQ27DB+PRzs
bcpMLHzfJLG7rtwY3bFgf1ePWiL0UmTJW17eYoLPq2ToN1dG8kHJk73JCmjQ
PZp0LMEGlWwUj+wdnthR4wxw/1/gQwMNsGtGoiUnK8MZL71JFE3v8oz9F41t
SN089PX772OvcyoFYJeCku3qkxdjOR2MBSz9487mt4vW6W90oLlxcL1mR00G
Z+0eH8YeasddKJU/p2F1Jev9AcQCDGliF6mq3gP+XgSn9xA/s/h26hLydltK
6FYUb2VweiLpUef4Y3m2M476EBQapl8wdJpLTRGu822nQOquBrXbdYt3crLg
YTZMueGsqHO1FvXN5Q8IZEiEGhajaUw8O0VXg/1KkudP9GBpeAOYj5YqEV14
WMzTADuH3jLlpvEKmYG1P43Q0ywSiffLZx5BV2VB5iFwgoMYCFVpxoXMmU+e
ib6cxYGgpHwmPwrqoOU+DBZpSBxlGEE65I20VlhZ3EONYnKsK1JNnzTSoFYx
AZ/YI9SuxR5dhFqXx8Y01W3ibZLU40lU5gSUpGyaVazIEwKXQJswzMW0vOvD
ocviBB7U1WYkf+70oSVd/+4iTPzshUbgbXibcl0+NqqtczWOS+AjvkJMIDUy
uxj9fewxDXvAXMe47bnRmoX1kUZJigH22cVnL88qG+GB/nLNe1Z+Pj8bLDNm
dK6vz9TAm899PW9jSyX1S63NrYBahDYnnByavhqVV2IdixVRHfPKzorB/Yll
jQRorzyBPGS6Cj2QpVbkLnMVAs2zTo73vYBzuFK6YakaAcO1aVI5TUi7mUl3
HrC6iXQApxzQ3KzAfGfr5Ar96x3ouTjT41UO2eARpBQNxCAam0ftsASnjqZp
kPif4tB/X+UBhToXdtWFHS1xd8fME/M5YUiN5lKv7xvBw8BLtXKfBX66Up4Y
awSSq8sOfiaP9+f/19R42uJEvHPu++DLc5wbTnwnuTNGZ13JCOhe4TzYd9HI
HlDvBIAkFFDFESfnYi1bk4quYYH1xMFv+ZFIQLueNLsVxxXs8jSxYGYZG7h6
7hyebP1OdsZn8vnnHq+b4FgQX54QQ14wLmVuoeEZgIuVDQHYxjScULBlq4zv
sTkA9NWg3nJV7wxS04/Pty9HrT7GXbHSkdAy6l1D+suAMpSd0AXsJE67gjSZ
rMPfsFZK+fLcf0Go1PrZ+Cwc5xDhZxPEfzW7QeIWoY2qcf+zt5VO9JuU0bBI
uzTSdklIcOPEquYDX544jBALS3Zj6qPtQcrLTo9pGIi94Q7X4SG3zfPsZhkt
T2gA85TlKs1Mmk9s4bGkUg8jtZu8kbWAJMVGK3Ux/YT9PLkJd4CTn+smNuUS
Ysce8ext6/L0pEVq/fEnceRD24TRYpPhxu+8/LKGf+tV7e4UwmbLTqtfMjzE
qmZncZZkDR1tUfiKli0Xd0UhRO2j2OOt6YATtAs9vJjjWrEBckKmJtiYJxot
5OqD86BWUH6+TGvmvdE0sWTaynYU7i88LY35HABps9fCLm3jk+xKBE5rtjtW
s/HWCEi+qx0pKa9crRyFyf64qW+gIB+VdAdJpimGFlN7pw+Ild4Ury12kUgA
0wCfcnvilmSCkNZ2kWlZVu662azOpGo3UZ8cUyl0ozzysELunbBjumR2ZLN1
G38Qqdd/WeaXAiYgdr0kYsHJdGYxKvtvFveBO7g8mUVe3ZHS/i5FyNbg/wKJ
166uMd3yNIp1rLUvlIq0LFsfDcTA9tqM0ombBEnMeolaQY1O6eAnQPd9YqVY
380Z1cZnPZJ3h4KMH6s9v/s4g93Rak2/uKkAa2HoQfBZXzdaofEoIEx18XU+
sYNI2AHFz2YeRMVpjGklxQNNdRbEae3ASpGTsRz9y0ZhvuaTbWR0DjawjziS
i3Q6+QSxcE9Z4mUCkDAleNypV9jICWBViUnT7PjS1cEGs6UxIHHXqRtAH/j9
MdxKY82cBU529ZlqlVVzENkva6644WQbgSgdKlJ5OPrsmYOmI0N3gvkJJkAx
UElPQxI9MpjCG5LaDWxzDESxrydV4Rjgg5tSDXhpEZOaX8HZiyPDRufmYJV3
uz5yMfYBf+kxZJ4AoIdhDUvvqyJLbSmlpLXmvVsLahYnppwUQTta5w9ymI2y
AEIqoq5vc3lJhDNieSBzNfZ+50kJqE7VuEhALsDpO034auwKTEkgH1xp1L17
9ajJg1fn0EmeR4tmptoaHnooXexB8/LDzrDgHzvKb7kCWOG7vmKM7dhd3A7l
jxk+94SUN+M2eqRLCQm9FWpPG15d+YXd7L6fz97Q6fcS1jXGKY2htufh9rnP
Whj0kwBPXbqPgEpGlAlXVnTqazJ8eJ5vIefcEcQpvqjhiBakZBn37aXM7Xso
CA2SO8UKxfKJORKCkr+QZDGOxhZYEwFVTJNa+g1HnsUBlPQHTZpBr8cfG2P9
FbBTuYnDMjxxfIBsf9d9ai9d7jLWaFsSn4SwLQ+UZB0WXK7vvfXYi3Dqsz3q
Q6CcldhsJuKOmg6SQ18THQQVzZ6Etm2gC/yzTdgZAbo/wssSmGa+qAcA6E/2
eVlUywDUu5VZ8ktFKaLMjjia+qIsq/zyG5LSgEClZ7M3ZtWMIN1RXKxs5FUE
QI9l4p53TlErczMxKMzjmA2fliSY3Vn9V8yuLiKOgIUlYWoItkZgNYlIqWMk
dbzGxim+40JbFGJRMfxG1ipFuP1YRKRNpoDX4HEo1OPEjV5bIhTZgmQOuxj/
lkJN7bH2TRmdyP4IJb5T4GZZsgKPf+nSnkJkcXMG2Vo4+vCPu0JRE0XH44fB
unrPwrnM0ao2iNsRx+SVEA0TSh1gbze3yMOIwhi5MsUU9r5kQhdFNZAsXtW5
MmGt4Dbj+meI/N3nBNI4/DLE2sZDa99wbsOO+s2JI2cRLJRe6Q3wGoJ085DY
CXvV9pm/QJ0p3SGRMkMkkPIuzu+EC7qpTw6LtDyzsGoCk03JDxrwS3ILBuWw
uKvr53+RkZP3qhxUlhR97B9cdc3+1FPX5df1VlrbX44l3nTb6AHHBEaVD57g
zAm6OH+lwz76tboNgZWInpnsdPcEA0toLuNSjpTWyd2nfCgq8yo1brBa32Ml
yRQZFoJ9vPknGNfqAmLoDtRN8Nd9d6M6Z7A1Wuaj9lE+U5p5xXh+mKtPbJDS
07gw/G5ow3Z8BkUtkcp79gMYYT11tRU/7L8yJRuAumaVejEkZEOJZoTUa9z4
tKKDUu4uuLjZU39so8KZwMVaOoJht9D0X65WjEYlkGzITHLtUjU3BK2Iuctq
ndqRuO/5bP3VXRbGIg3e6YDqdYcw2arizwSTmvYMx3u0b/RVl3/0d8RnkR04
dxDI4ss6HazmDeNwRpJnRxYIN7SgZTmujEHBlNlusCxCHOpeJEs9r6I1X7Ht
4BDlcpyYLkXWsCN9b4/zrHU5/OxNnrgSpGL5BnAYoGtvCheEabfMRgeNf0/Z
z+Cxs6WLHRYbFPvhTqKEewX30DJ6QJPYozZqVMF/FQO6j7TaoXDBvnWD9eMD
c93fQ3Msf5rbr51QvXJZ1YJ+isAS3pJjVi6uhnaytp7FHl/z8eo94+tNk53X
LYNGEngk4YcXVhxvgSyxqARdXaEOhBXkHU4cOIS/2K7OWtqRUG2/mzAC+Y+W
WKxS8JMbPEyNSP3jO9Q+GsOdemauUlaFXPM004ywo/FStRuR7CXXRRFpFImg
eEn1zAHIPDJTI6fU+M8wzEE9GHsi+1/JIEkO8bAXkWwKpOMfIIlT9Ew16Imn
DWZOhS0V67gMOrC7JKKSlgMenwpTDVepgZqjuTAsDw0pqhq/k+YWMp50TF0Q
QRxMVwguONe+MUyQRMHl1CEtkOhWkI4PpO/ix/ZB3FCZ1isgr6Jo0+pBcdbb
+XjDlkc9VZRMR7IlWBXi4UDOo/mNrdVO+p2V4kMkvmN2HL8hhKQzRIbWIle1
AAd7+9cCfOLtViAptP+cqlPfRoZvx5GFHHDgT3dzPS7p93mFYIPXBPYYhjrF
rSbSHEqwjf60PqeVM9wLG/s2H1MU1uCTBq5Tj5pvqRv0cibikj6x92jnxpww
iyYvS4sXJaDP+7D1iKae+DHhTupcPa//LOrwuHYB2ulpMGUSrZ74JPj+GQg2
JfGUvRUg4uzgpROQDFsOMhonOLpR+ExhTYJkWVy6xPjR1DrOkcvXo9Q2/ICY
zI3iLPbrWTzDx2W/yQ3WNEhwcfJwY1YQ/GNDHP9IyVwHNb17xLFgMA7AO3B9
dd/0Nz6X46gaCY1a0AG7jwsXkn51mydYTEYgAZxsAaanczGmdKwJ241+HK3m
E17Nt5mPcoOzY+H2wt8RtzlewFOkoVusP2Eoro9L9Z/ES1CR6Rg5Ux0tNBZt
IojCvAAElLU7GG1B5LIzdS2K77aJZERvA8bF9udq6Y8WPssW8HdkMq7pxarP
BEWEXpm7gitDdgTRhp+fKQMLVkD1WOlhZg/BdbWbzAAYBxZ17E4IP4KQuivk
/l+A5yO/L4BzfrYZAWbJMDcqGpFEHELxZw5p4ORz+IjhEbfuRzGYZX2dPOM8
NBeLUxVKQu7A/RmNpla59nR55w89eo9pltUMqmI86AWz+wBro9JNfw4t0dJt
OmBlnoV4bCCuKkBD6IB3cCnWO1Ip7lcAuLKM/xKqfDj9Zwwxbsy/v3mkt5JC
diux8iVR848amUEYeAZYz3mPufyOBtKklMpvvf5MaxchOJS+AKvDiOYi7Kye
CEgSIfBW+RR9aChT9lxVkbo1tmoHYZltUCiWg5/fcRoGMoe+uqLHj9PdOKrW
HLplLY8VH6qOrViUmf+3XG8P5/ykOPlLhKXtOSZIE6AVIkCWwz8fThQq61pQ
mlrJ0oZ+in3mMbVQBhFIJU05sM4YnyEasG2cOxHf662GVhRcUUcbM+gIFgcr
oX0VYB/3M/GKNNU/YTuZhLtVubhV0KElx9sdb3eqzX8KBy/F3AChHT4q69PY
YEbBKZCDKFDysNPkuYVxHOQ4gXEwgKiXr4CJ8sxbm2hsd+zhXXu0pVsLDxIC
SkjlBxHHOIvIIpiBnX+N16rKyV0wusOkrT+Oh0n6PG9r+PrB5mOAcGp0TyJ2
/deEJ3lQ4lLUa+kKGApEW3DTdtaoj8RdWnCtQLBn7F8PIsD76BBN0YDqf5Ac
1q4SblBUi/cQPoUDp78PnBVHYSUh5hsMTJeYdHelWb71a2gwtIRQ+eZ2rqZm
gjTV58sVGXySnyprRHPivtA+REociqlR/SmclfhQE3gya/4lPNrL68h4+sCH
9ORgLo2Au8I28Zi4ZN/rB0scsti52XUwatIqkKnCzBfOrfLzgCe/ygEDxtgS
16RzLnEmEA6CTZ3jfU2Yl63RKljzPuDZYFCJN+ONu2QiokIY8yVvpyvlUvSS
G5nXjLNIWmSDmwQ6VkNB/BY9yO9H2Gns0LJ0LvdMOfVohXZHMoFPoleD/ck+
ZWzkKrJ2UMykb3liJFDcEPTGSduf5O2+Pl8CBTd4Qo2LfT2mOo78NaIyLJYu
RW8blAGsYOUIv8LgLSnPr+5TYE25Uuln2g+YLJZ2w48Ysur1kyYu2D8U2m/B
irwKFxG8ljl+Hzpu2st2r8hmqGl/7DgJil68TtBysGlgRyAZUgnnFq5JOfFU
1O/4EJjdihK3msdkWavLbiLoBmqHx3eTa7KWDmdv4Qt79FNjRTp+D+TvgC6x
zzVSXRURDKl4XW/vHv3EN35MiwBt5UFn+ehoOsKE4+cQ2uFa5CK5MjysUEOz
zQUzEQVZsoWJDb9J2T8BM7WkF10IfCbpXTnzPd0pZgJRJGfv1PCUemTCs1uQ
92i3hzyPrth8jpOr/JA/TUwml3XeLXau+X+TWJHYPRJzpaKNaPWdRRIgfmuH
z7bceW2hp+GcK6kn0kdN6xjxMqPC67lsXd+iMqvyfVwK5P4elvLBOHiuki7e
/ktO7aJzlUAmB/R8zJhLH+Uy4ULjoabgGSZlID1q4TbHAoq6VilBuxXMR8ea
/hCyxq3zQEJC68Kt8m5RVX/y/ugBZh5HgfouZXS387L6xskC+/cjteJct6sK
RnX0uH7Ex32wPMiJNPbxVcqsyJzp0s6AN6Q88VGCEGTfL0rWp/hfh6x6veQ3
qsuyLAm53e+Bwyisfh6hP6xvOrHKFpZSkuerwl6/w5duhoiq8VS/Sc8jP8jz
y7WpYtdJ0Xjtqkf4mubfD8KMdWHL3sIMw1+cu5cnMc/HeKY3PnuOsdOdXIPn
kwa50QMf+f0SnwnW9HrBHXCTC21es4WTae3dLBp0Tu5+o3DouXJhSfQ0LbAL
+YFUgGkz6HClzKvm3ZkWPKupckyUZIX9ap2gf/Dda2qzLpybjeBs8VYIWDCb
XxpQa/4mf5SNuWhzJzFSIW9HB42UZDiaQFiHNu6HishSSu3XQdd+VlfTqGW9
w2jcO16sqx3qQK4YKAvgAgYX5/ZtBw254H3Iw2+DOkZkyKMu6Kk5ikU/SeLx
zGynhJqogdKFA/PJ34u9WPI3kXt4qmrSU3PSRlxRvXGCs9fUlM2N3PAZNp5y
8JIQnHi7LmeJHPwi0EoXfpOwyYmpZaSE2csFH2VCgLFqENrT0kLJVhLT3l2s
fDxhtiFMX/3at+irS2WFSzuPrfDbPbTv7M4BdfKB/+uZSKACMTmuecQq4cp4
sBpedVsqr657c7p7WXeZ6wcqu6mXqX3m/DRSoG/C2UwcoIqe+ZBLlO4D3bAt
YM3XmUSCvjVboUvk5AUChHzjXDU4ZDQUKUgVIH+Ki86aAT0lFSoVGZjgBlz+
A1K44oO7eAOPrwgNMtofGDZ1vjVhfy01JsYYprI3aOjRl7wZm/aXem7JH9vB
zpg2G4mMEoZABhtS8q0RPq+hwqZHyT4ZZ0r51ULWevqaCy2qD/6qq/X0zHqq
sIDkk9j62fQTHZZvjOrKedtLPRe4z08srzO46p1XCkLuNSnq3plYQ/XxrTiW
U5mTPHjvNdfJg1YgEV8+B8qp/Mun7ZJX96Dglbh4sTS/uf9z6hI3Udumhryw
8X6Jt/CD+aTosHH/K4M+VLLeweFfG13R8SFvA00Y5zqlTXP4aZ/SOpX2pTj9
oOaENx0r9Xs+SLunG41AhxN6/hs/FmjZdtMZpJFiZcOFax37y47/ggnINU2c
xPg1jEdizTRHTbuRX3AbNAh/sacfmA5cN9njeg035uL9gR7eDtdm6tYzN8zR
ht7+RxmPmOwRyx/Frh1dQKSm2Zkyx79696q7HmAL8oN5pUeqfeAq7cVDmyoy
rQFowh1SRf1hO+QJ1G9SOl8vOCWe23jT2n4XNnVcYyLBDSebxpJbutwlDQEz
DWtUtTKYcuQyMAJZk5ToAiEK7V1rCO4aTPSFSqw1dXyK98eWkMRa2/y6hQ+w
ddRjXa4WiucgJ8c7g819MZH0eZQ77ZLZ2kAtGUcV2LxBKEHlhPS47pGiNqQ/
nPsHqdJJt1jGxhJcisjcJmC28HUjR9my9tXenT3njzLhROIeSgqDPLIclc0X
6vmyzMRggUk+CUx2S/U9yol/+iuqJD1uFofh87OavOIlBy+NhFYsiYXwAHQo
I0JzAWERji59tlGM2OvSzcgPLTsxyh6oNo+O9t3wGwXiHS2vZqWiWQH58rtD
d20IXcGnqan/5JgApQIzFWlduGz9KTHELiRBJTiBnN7Ug/yA8CKGzNoXaRY+
dGfDIiZqJ7ZcyYBfytOVLybM07UAkeCfoQnANQpPPnSd+2Y2KSHMOQxx3VaB
HGVb1lx0cgGfgkNKrpy80mJ/WkLAtiNCbG5DN8dl3hUS+n1h/yKS6LOLeuq1
0MmW+Fdl5OvJNbhhknCmqEvsQ7kr/UIaESkEjV0sdhALlXkOKW3SPmPjbpi3
VD8RKqfLOzepRcfIYh1UYH6XdKwneBFZ85vMGkjmR72w5jP6qbTY/5IB2c+h
/4dJBGcXzCbi8txPc+Ah6HgV5svPlyMf2UMxLc53BcQNE3xjTsfcqzhPECNv
EBC19nDTYUCWC9uXeSyeaesfkP5itmveCj9XuPjY/XjSKaIIuKJ/7Mjr/IUw
CPMHtJ9tFQAqn5Uh5WNujQgSEKIEXn9qox0WFI2SxUZ39ysFK59p34zVYIfZ
+rdX8TtmVwwpu8RDEGbymUwXp2/v5a5SALZ0xqh9c3yWGckrmFUA/2v2inss
tkH/aLORIE6U1p/VpEQP+Ocx6M7FcLR342hbb097BoFgkCcNokDRrCODGzUL
ZIYMo7RJwKR5KjqkY84Ok7BQLaFCJWR+uAJwVIeWMUHmgfoWmK4JtUXgNkH1
1Mas5ZPWO7G612rubxaO9jw/SqV4NADELyDvd4akbXo24mui1AeLpQh+xWED
HumovckD/MwE2q9zKK3JbYZWqnjCH5L5rhfIv23JV7N5DFkrsl/cuGyDtl46
HETFnXXgmpY51C4GjZnzv2RJmF7L3a9E27tM2bOtx7/N9kpuUmTxNw64h1sk
/Czyu9SKl69juEnWSw6c69M37Rc1Sj3TlMIcG9XA2YGAc6ai5D4QmiwOmXX8
2/IXJKvX7TLQwmghLWktssjGVFUihodfcY6cnK5SW6VEIodWxQxlJGRKfcB8
1xYl+MlRTQwk+YW8r0ub2Pryy67FnbUc3HXb/t5Ys/Rvr+L3oXw7zZUvtEB+
Lf4JK77w1BJ95SmB+FtuGGmB8MsrIfemg+0BeBWKAroajdMvMXxoL1gxZTUI
0nsYlbFMg2w7zjurIcde9kUYqCIjtrJdBn/7T4zNi6hMJp5VpPGqI64+bWrM
xwiA46gAer6s4JN+iEfwLF/T55KMAzahNrLIS3nSQMS9otEdxM3uY2vnMoKB
N2M+GfFO22RqO3wl4wXnAQPAxM0CtmHNbh/MNy+qugaKa/IG+7N2bZ2nRd5/
jsO+I2oGXGs4WoIe5UmLKYMmKhjuxGyniC7s3mDYBzpfV9umAkGF7PTG6u0m
0VRXJEzrG8ocIMr//AqTfBoOBdMHhgixI2Z0yA+/Ogb6l49m+HN0CUmDSSYd
6GPkX9LXIjP8kKl/MS7JisxjeTmsZjBmc93IkkZ9ivD4Nyj+pkhGTIYzKVu/
p7U1bixdQ5HBstxB2zOzlXoG1d4ayRXunAUEUsSbH2NZDqfveFoTrCxWn6c9
wUmCCtNr6b43OnwoIK5CfWnpcqeth22aR7YiuTScIyjYILbS8vX7VKjQVmbH
Z3H1V8thLyHhtC6PA6wAGaHQPtqhFrW3DWQxyqd7FR48UFJM536QGv6CIcJu
wBhHk6B9hQTisYZU0fUWq+wxYbevoarQ7o8ZNbPM9tDUIcp1OAHSBBNcWVed
zs6lGj8j2sOusSgDTegxCbg/m46A+rElp0TBvtasBTP03kw3FNitPMlkiOIT
b8uuNnnD/Q3n55lv159Ac7PT0ralvnCah5WKZzLBKABlYCm08yhVC/wxxMwD
/Zvs4wMClzWNI4ez9B6q4sSy8z38BwBGd9RiKWLhqK9vnAWIajiHPLfynbb9
cbyma7sLUYejgWpiJESrtdyiXrsmxK25UzxTaLhYxTO1FwTdsZk9Zf/nEt+/
8EHHy7C8k+KLyeGafrHhmQDtPtRIwd1t8JzLDkrO8u7B/bWa3kG2Fh0z3pjN
yUIXv3B/CZJH/36qtZEJoVZQnTMb7M5nz3xU5IzZndrjP87v5GRBckeQKnLB
SVFJhiPHKpNM+N+a2Xn49xMRH3A+ltYVJ6wR3/Kg+xg/UB021nhd0dki/wpe
ApPtsa7eli69lmCCYiWxcnHiMt20oLj9Zc7FOUL/b/Cw3LMZjjnfWTZaxPfy
1DfzelWUX+bqnJWhvbBGKdjMqdHlm4Qc9mxJqOIyM5Y2MoSNjVsFMIfYy4EH
129tyFmJ3y5xob7cj5yK/jrckpPrecJAhRlGUvJEHmMsZouQpOMazDQOB3cg
R9eaDMfGTlgaakubABFloq5yuONTvsFmv1+Yq4uz0g7QjQrdgce79o0m71Db
Cr+20yNDBsqk5lQsO5mBpAwlzYSpJQFbxSecmA2R/tLtJ+0KrEn9tIz/zksM
6/vUcjrMzdXO+wXXohXRI87OQWFBOYQtgdSW4yPYiiRNtGDs1yL557VVtDE2
aaU5jDB+RHEhbCj2i10cBwrD71AaXyfgiOEzHNNyPHQaxpQtxKtTg7vrtO4D
ep1AP83KFVsUtViLq2Zm+Bxd08368BtTUDLRJUVMzMtejMhoPrAWDIZiV5UN
7Mz4gWfL1sGeI9CtKrdaG6byYPsqL700W11LeRH5TyAJUPB83eSMXY3RZOL+
eSJCOA7MHZqIVxSd4Q8SNLDfuGQtmIbLix53l9QaFn77omvrugTBlTSjqOeJ
uzyVC4B5Dkqzpc7Bq35RY352pKDfxAbOYeiO/4vMq4N3lp/bq8ejI7PHIuP5
kcBNg0xF3iu4M/mpVyT2dvPY7ik4HfStocu+BRsE5G/MGfnUdNzcp/jPrDlv
+aFskqiZuOpm1epnx4hbwm/LQZKn9ehLD8mtgYCKJyHOq/Ehue0ZkmdbmE2M
BpXvAz3zMMxNj7ofbH/5ahzOgUUbv+IamQGUo3ZKY7EcYWQ6u3sNKGaRHC2Y
s3DO3RoXgtk3asEKqATPnyD3zRCpmTUyGQMOkrN0dDQeQkf81lGNZ4/G48OF
RkBUKWACZuiUXVABFqXKSH6sFGRbykyOz8AISs5t5vZv/dYv9de/dGNZ3WF9
j01MdFP88eLsE5AcCfWf5j+SGDpTXzCnaKR+eYicbRluFKQf3VTnM6kiUap6
uJSWPNjNhy5KABUbGNS7MOETI1fiDc0lMpkwnLHDCDgIQrLPK9HQ7oqIH8+0
zLEmbTuqONy+Wb0zFrEMavGl+hZ7+oLpve8z+3yqGdQSUdWwUeXSMuGzeMvK
i5AESzPBOtvSJIXvt3Zg99QWd1FICLoQBRIz46o7k5Fn48Yk9E1njw5l55dQ
drr/nTffu2IdfvyGxaulCkpqhgrWEwTsunQ/r+JKDZqjiqAq4S8oDrMIge+5
3Oa46X3kLqahHjhCKbnLphoEcpYRCqU2+9g+1IgN0KOI1C7OQKwOSQoodL+h
1Tg1ziWoLA+PliRZjPlo3/4nnxTjdueMBd8fvG9Z7RCGJ+ykKDJnx4Tbkzr1
0fVQKLs97mLIiEaQP1JNibkwvH6T4PsfJKTlGKbVuFHHWdmjkatPogOh19zc
JC+dskZA28S+QT0++Jg10eS4P3tK8DMnV9DsIPl5egEIBqzpmKp/POKJuljD
hObM2pBc/fy6T7sbG+1jcRaZWZbgDxkdlHlSXdS7f2wQ804tdPYNpMWXG7mW
Gzh2lLEUTdjIqydGLXcN/TmwhzA33VQ098iCoAIcbFUNaIOcUvYPvLfUz2Kt
47Rv1lLQIBzfMjztdPJfpt6LcZtSw90XLpGPaMf4+aXdYqNgFB1YWo96kO3Z
7Tf4fVt7t/Sm56FQMmoBIjrvu15S9Ia9Fr3APT1e4Hhf9bJ4obnaIi2Jog+h
EN1MwlFO+h+FyjGXd81klcsVpo6jUsJ5qg6KXmxMbxFJoz77sVNVhb6w0CrF
swdHscKNawMICPq9sbZJU+4gPr83UcfoLpfZNiIOg5/Inh+J1X94Skn7MNko
F5dbMyaNavoY7fOmWk0a8WVDE1WrntsEMLqFIu+PkPP/5B2i2WBqJ1OGJ+Zd
AVrcxGFX9mzX3+PPHC8X8h0bB7sT9bC0+zIgjlpxCMfATZ6Adodr8G9snkcC
w2wmG2SKzoAXjaj1Ki7LTkpL97GGXXdnXxfB+Y95VaTS6nvfV5S6yO869RyA
WxWVlGDR/tt/k8D0mtXg4Ats2zvUluG+m1KS2mftKSMw2aromXZg77muUCqC
TrCfRVv2ryz1qM89TQ6Jrm1PlMjZi0JJ6yILSZTz/QauNBaLPAbvlqO+MK6W
fGfAw/SEm5emkt1rqRCHd9XH3CBc4OqmbFTo8p7pRohoyMB8lRar8rlCbNtq
8Lat4DBbO4+BPq/U1mvRzJDhYKnLqTbhvncTMphLBpKxcukVze1ihlXCmLEy
1PTxd0XbDo30VlZC2cLKY4LVrawG0JWO8eHsJu7raUjyBCQjRLoEuS3RVqqz
y5pIAAbUt+B0ex7SRKQJ+fJ5iFKJ8CLWSQ/qdps86kaeXt5p+kstGGM0bDQ8
AitgYXOALrbX+E5ZsndhmVVSNDI8XozEzo+uwQuzPoQGtfiCqBIOYOQG6ofX
xuInXODv3ZmCDZ3ewE0ZEAYRWLA5R/mC8uWASRzHjcuKn01gwZsOHy6yC+ea
Duplbti1nnnODLWEDpilXFk+H6KbRIxN/X8JPEfhgTX4M8HWZqEsoCC9VN7h
shTQIFOKYmS9t3eVESn1Mc4Euu7y8e/FAXvee4EMqfzAnsYzdCj+hm0CJkI7
gIOL0COtX5BqrgydLdwVw9suk+Pigg5O20Eh5Mw92JFZs6v+ZHxTqizApmrc
eXscSxtg8bqJzLkl6ufEf8VYjvN75sRxtTYeBEvrd+Nrz2bINRgY6CR+toyo
oBGn0dfahpsoXsS1aHEaxxaHK3dsdISZGH/uRWkNLnwdV3gXuRKbZ3Lxcn2Y
huYgexmr4EJZV1RwkaUS9zJa5liyPGZaeL/o3qlj0QMNxjpbpCzI9Bx/8Y9c
zM+f9HxN3DJXQEGECAd6yQHBtoPcVjqYGB/Esk9zFyxXSvgOKgr+eg0QqO15
x0AZBQb3h0gfP9a0YgFPkrGhyr3huCF5t2bydbHa25wiPTFsW+3onRzYZhMQ
NwVusZ0ddWYmVtX3umL44IxF/I0gBIIVeXkeeWO0RS2HgsPiUCdoi6YF8x/6
ggm+ftVyQHjLYbOLvlNjhwpT/aY2NDsfTf0nW+YAunWj/X/+cYkfwEaLbJHw
xOCv9rel/CU8tBKBWioBq92ydSZs8LlXoIK9L0gdRDkc+mIeHElY1R/GiGfo
AsaGwXk+in0J0AY9r4w+A6T6tX69dIMsgeG0XnYSuE30XdayRT3PX6nwdApr
7hS2jt5hhvSUT8gEhS8Aq0e6049Apg9EbXgWoFeGK3YgK9CmIWtKZjRHPd32
3cVWwdOxprKpn/Q3z4R4xq+SD6SzvV6XOVVjLu1CKAqZJrLU233ipAh0J1++
lVm+e4+93hDx+YmCNwDp88cbJp2pQDO3ndDe5FzPbqzQ9nLFIZYnsVRooQhL
r9LwcZ+4mHU4RbxtyzGHAsn8CMlymBvkIvwPqnYAEKynU030IWmOJoHCpMS6
CN+pzHMv1MygEcC+iaKapB6m7LLUKOcv1GJ6J5pLXbXw6Q/PFyav2vT5Eh4E
8pXMhIBhwUm+s591/ZN416OWpTMrRjLiGMMlsREJncKEeA2owaYaM4RCOIar
67tG8pW9F5aUMjd6moozbuI+FUMiW1nzHtjJQ92he6hKUd2acJmkhRsNO6m2
iuuh5CPP85x4ZP/umYHc4E8BPALpgxgI+Ly6vcsv9dmLI6mTu5e5147jdC9u
9Wz0iPr2niigDnmVLuxqMmTcmYsnj069XQSz4PoiFOl3OwjX8X4wqA1O3mkb
J1Nbo2yxpv79K1nXy+Se14o3TsY776PRih5/PV6F4LV5L6PmT2oXx4X4RQfS
80mTMecRO2o6cHyuaahsHu8jrkbHxdnIh/KyfrFzu4PanBpjwF+LrJDVBlpV
7bx6u+ulFjZt0yrysD6pCQ40U/GSrFvHRWh243VUMZBvUwt+3ulexuHZSr5d
qv+qc00TVH2tLDEGTPqR30k7dvr5FvBbMvzpHD+rNOvTFOTn9PFcRpRUcD25
3UUQnwbBXOioqPowNNwau9cOlUaxxxjjT+0CpLB68dQqzC4HsgJ4LZwUoAIY
7KoA8j3LUiZZmehPfzpEj85Hr30LcCyck121Q6wcQJa3mEsgmVO/8An2qlDY
vWFaowlSyAy3Shlyhzv8ki3Na9GWZPAjsJS7VBBllWTkQ6eDTGiYzxzJbMUz
q0mGan4q1vK09I3FZxa9+ICatFCajpzP0uaV57y7U2dwZou7GjDNw7DHe8W4
A1euQONs9qh8vbpVvWi5Nbgi61XJHg88YcH51lOR9LFFPVx9HUxR/mCHcg9g
vpxBDO/wd8a/C+JYceaI1PJNOz+u6pruBARw2n2LY30Uh3IvoaVfLUBxhOHn
d0RuRqnF/kW3miKyDF5f/t1HzOd+dqXe/QTPuIxheOtp8jcozonNDAp90Us8
8GLEkwn0I3wZYxSXrRHpLYnEHLBNbTeNYwYpqneLcCLLURyzxpbM/Lt7DXvP
li5W4LUcyVsf3xbjSMx+Mmy8HWwqDS0kul9qkhYgGbijnSbleZ7AkVPO1qC3
8yrANO2OsLdQRyO281Bdq36NHlCAjovA+GFp4MXw8azX/V3FlcwVq5y1whX3
k9c+IOBJhyTeMZFGPZqPNFwds08JwArcCDPwmmDZwr7U3SSX8We4QXdxVLJf
VO9YMqmOPiUtDDofata5e+PjNRP96D5CeG/8Cofc39WitmRQk8zQCV3ysu3b
K63pfq9gM5c7NcNKU3IBr9ORQ06z6mPUt4DCEJhF+EJMjq4Rf7tKzcS8nHAq
WoT2cU0YV8lKZE4PkBmsBAsN2Mk0mBTFbpvvzSCHD3gikJNJkXqBZT8IeeTj
1Dy0xGRrlUmqgoS/nV+GSUJdl0JXgO/xvXuh/vaRKpHetT6F+trnD70jG3b2
fxWHarYT9QE6zp87jMkX8FzYhsrY5DfTQUt1sD1DA1kDbBTYZiXHipUUf1uW
RraGQeTax7bDJ99vM8+Qu0z/JgKWm/16NZ3OdWcfNU0lJejrA+vZy4e+iyPt
fM8cn1rTKr79TYUizc5aB31GMHn0z0ewm9sty+rVOfhM1Ssq8wZpTgwWwaQj
mtG4uRV7gX6/CXy84goWE8qYkwCF+E3ZwpLaQQejmQHmHZLKUmusr9CLQBvM
8ag4+EAi62MTICB2kgzP4VH8LdK2AF/arYG2epoYtknWAbZoMCln4QiD+/If
OUBa4ZWk/Pq8bhc3xiyTZuosAdq83AUXMtO/naFIljQYWO2bOZrwUkr7ojmQ
DC7BTNZV9pOoryXfwp8jlK8ivFI+nh+7PqJDXWwwMXIYtYFSNCFMfZ361E0g
0F1rsKKBulM/LeCpMwCjUysZRvALKV3ragUc97RthxT9Ltn/2j6eZ0rGayXs
GivfuMQjxWqn2+MjfJmJ8YfnajjrTfY7LULxVjQ0gE0p9+Im2VEISsb0gdmq
87pCpnz9ea5Dxbtxg4bkQyjet8EiH2/ort53InAxobwB8sPM4wFjw9BkSrdG
lS7gasIKhb4Clf+LGonVha5MzQDYDvKwO2jYhFRtJSJpnFoJ1dxDw2epQxyU
f2zWQwayiA/1Ry7miIA99SRS8FYU51yHCpNAg8R2CgwmVHXrFBH2P4C6yh8/
TdDjCB6ihW9CV46yUFSCXuMpQttyzTHJV21r9MiTDYSzm2SPE59IAhkvgwQm
fHtl834fftyBBHVthgXYfSHYnGzmp4zPzrHNzOVv6LxOyYtSIHCMRgo+Uc6r
806eka5QXaMpyBzM1xNWzAf8uJIwvXG+7gjfRikOTyqe1SVwpczCZF94MqCe
XFjpL8a1FWBLb6mi8U3TbvXovq3n5pmxt9eJ2+kxcMCqsiNl2nPQMvgYX2x2
AOaMRARNzQDOn35M+9y1m8x7uh8YhIB8+Z81FDpIGPH0M62bNjjkWIWJ1cUD
2oCkKzGXDPaYvWAqd4RO+bPnrYbDpi1y5wtGgLaIAILebW9cp5vpu/KwQZdL
q78Ee2iikPhDQ1/V4x1DHvKD2WNjj6SnJkXWbQpk4wWanmmEaAv44HkzC4D+
8qpFUoH8OBEvLMazglKPNWEn1zFTwJWGr5RmDsMz/1znzhGwHCABWN2ji1r+
yqgP00PIWLLBUjIiEiaXeorsCfB9gvLTDZq9rQFnpJVm0HafP/myRj+xQo/V
1icEgO8qyA3Uk2oD2ODqamN8afMO/lUTfGYnZ/T/YD9jj0BAN7W9ES/ykNPn
CYC+alXvjqs1HI5WUAaZ8ki2ATQGwgDtp+2kmWzgpYyZtPPbqnloztTlO+q4
gVWbGf8+XGCDEWTY2zB/vjznWOR+s6pHEt+vDCus5GDe4gB7/ibnKKn/+BIT
KxtxVZgYir1luQQHI0JgUGkMFmQUhBlfFncnHgC/VjU+KxU9q7SUbnTEE6As
N+xiDI3i29vj/gEnA7r/WQFHvh6AXK1r/YxVfyHaARSLgR1wQnLJMnkWSy8j
htPwDDzqq93iekoZiKjrTa7Wj3csHArJpnvP6XWIAUwuDrZMBITFst9MGGA1
RiuRcwOa+IfJQPkisyvPefoUNBUpFdzqjXc9Sc7zQGLbpnhmVZKs5Gqbcxlo
boUkgcgoLLYTBVrpEY94Fx00e/gYeOODajbHOsMKlSxfsVcT/UwIuMw1LdHi
edW9SRsFu128PHylcGBPjtZq2mkElLEyJfeIkGq1ZE9NWbUH6dnx0nT1feCY
mKPzR1n9TMW2T5rgXP+niuNpGQfKdMp9vqSf60UOAWxDb1c7DA5Gs1WAgKh/
goemywAhJzpEP95efZmUSjOlb8gEsPMpSygv46aUjMy7mIUJuxpvdbLUynEb
SyBAmPH6QTpc9vHyFQkwrRFcgtJd07YGy+r7NFLk2/r0qVVzxrLgpF0Zbt5D
j6SlricOx7S38qDqZTFxmLzoOdhzGJrfc9xdvVRnqWsQwbct1/Mmy7nCz3Pi
TLWpUckKWv0CeLab0wzw/li7103HGUnBFgPEfDhHrAdJDW6lLv1MWpv+R5nn
ssTdtDhsopR7lFEG4qut1Qz/dMz9sRO8+47ZvkRxqKTq5dL3KMwzu7/Sdy97
C3qhTleqJ4eoIdZ3XmMcKKf/ClD58pJp9duFz8VCLdWwtOZc7/eAc48HN/mU
QaEOXJ9jsKyQn3E9k1PX/NJdPE89unlT9tMyUXvylfnaIzo4Hoze33VqYDkY
HsnH3v4Bn3ZX791v4F4QsLiyilGqkYBR4piye0r3IJ46MQFAsj8EwhSihL+n
VBMGCJ4ZA0rS7tBW4FLnxGuXIhgnBlyQnhT6TwUDZxCfykPzRJtsSUbEzmEl
QP6HLby/4Dl0XPazbIGS/HujDaRTZg04o/O4O7AQsmF6t97OCHBCm9plbmvl
lIDfZsBDgKBCWXGS+poGKaZOVg0/+vqu4H+iTQrMq5J+JQoE8jH0E7VWLYLr
TG9cc6kzPE7UrgLUCrvJbkcLeT/v1JcGRo+NM/X5u8nNGj+xQoHw4gZQs+w9
C4uFDVMvWuMZcdlfNDC1NBxehZAGcFQntj9SNucMEW+VE8m1QJiDh310te98
Q82RZpbMI3R9dZVnzlSbu+KgM69LkfJJM0zKqqlsCBBgMPEUiFEv+ItJxmVY
qYIDa5AQqRzrgxf9EjjZLWHp08dfT43n5duXA0G9HSDbU5drLoy4pWt9ng4w
X49WSMuDik62Zl9Fb9blL6KxUSeFsKJp9KeyxbPIW0yi19PaByk3K/sSWQ3E
lc2QgzC0zY8og29H0wPc2QYljwXBLUNcbYWeDpqvDcrCH0OWz6YW1JB9G4Kz
1WrE93OkkEuoWBZPLbGeIAJGWHvFZUt+AaWsWz1yISY8JbiJJ5zrvOkpdzWC
JmBGcJJjGFSZnpU/hz/tXECpa/VmZNAeJEuX9fMiX8rgl8uZWvaI/0LVgCNe
DsvUlyih1j9TI+VUjUFrDuoFV5DizeSSgrbEvTiecUpA+dlzT7mWX07uCxg+
9V/n5F2i2XU4ghFjkC4JnsYchCcJptTtfAL7+wPj8BS0GdT+n7YO41W63kwS
o0HW7iEKM//s5Gwvx+8Hor9iKSMc8MprNbi8buJKIBCaow9sAS546zvgBuKx
Bmj1kS2VM56coeDseKpyyiQ2kYeshxTRw/hKOFYdVHf2HXH82sYwlBQamOxI
PRM7XeI+K5AIFtcHS4Q4qs/DcsygB9xJ7pdiu584uhW4XiMMPjU6jiJDQCQB
Sl2+XPlGYDidyPPR01tfT+1DBbsiUnl7vYy/woJG3E67B/LzBnPkZ7oCsIsp
uVln/+RGLo2zsWiHQpBrBmtd+GWjz/CeRDipueuTWpWobw1u5g+6X1buMS7I
68pa83sIO9PQhqlFj45WnUOp5GO3jGODufFmRIHHxZOqgrZqupz8C+D2/Khl
cWNYZvoImterKciMl2u87XtTTPgixd9zOsqb3ZH5jlLQY9qyZ6lU9vmgZHFJ
qd0ilH5g6/XhCt7uw2rM4Oa7y1bNCQicYesinE+UHEY4pquEej2/TIiN0W5y
aVKDex7dVI5GgAopIcYwf9AU3TYM9dcOGZJLI71lID/U42qJoptqg2YzYmnU
1TYNEwS409lLjIqU9XeHffD7K2+rT2zjHlCVRHglyXpu1kPLYRSYZEjdvYOm
ulNsiDqvPRDEM+fZ6W3A+q3k2G/lMPSlX8z3fZfu9ZGIgsQBBvJNLBuNlsLO
xG77MtCTglI0glRobaIEqe3catcIyQxWnAriWKBD+w40Bgjvk/FQHEojZZ/K
IdGZau8TQDs1f1fwEZ8tCvP+X9wcXThfdywvyyXWbtsCNwKQdCJIIlYgu63V
S/8y5Pb4CLQL0l5LYOH+vBMXl8luGdzvEcWGSVRPdH7RYoyu2+IJs5ATyBJz
WpwDxCFlyKZBYL8M2UOAZmRlDVM6fQ4JzdRYbs1xphajFenSSHYlqfjqsNzw
m9R3jvKP5Ts1m9BQCcsYpQOJ2AN+y59jgTWeVod1leItvPMFbr8pclh9OcLA
1dm/hnHLzhE4imzOxb+uE9plisIfNKuNihWwDaAX+hr8Q7f2o5AFLIooM5pg
Ha4kdNtnzeWZ0X4gRD94EHRsl5ghdlM/uZwS7jG60ksVhyHbcYidTdmvfpHM
3sX+TF1nn6A4pjPGdzmoBwqPMgWpCppeqItf4+FwPG3R9lsYXqQS8+36onCz
kZ0M2EG6Jwx8941HAknwuJiZ0MyYztocNDjPTPaDL3AwQBTi78x88GnZYWAC
b1JWLKDAZrlpt5kDcMjNipbRH8vaqgL2UEgOlLN2/vFjlowwq0oPESWbGc/K
IPhgA9sXgB4J/t/PhwudoZ2DrFduFoLleuYOqYvs+tG+xlVQRapIUverNKNU
Yw1YzOyiVtN0n78NGC8gPiX32Cye4CKcRHH48um3FV6gVHlEsoGN7VOmcHvY
UyVHPC4xTksTIYusYqVZMWWhvcEN1/Aj4FFtHR5cj0VYpgs8ZUOxyXETffxf
CkNaaXOycFqnaoNSnDxx3l7GxQ0NbWBDCPVkXWkBlQSsePHGH6+XXYZwkdc4
XYdafJOs3Oc+R0UmqaE6ukkRnvOWfmRLPNa5Re0W3n2J0ZkC+/O9ziS+MXCT
DWXwHuzPfXpY8rkc6EY8m4a4531d4rPQtuA0YZrs1LUmBDiRM4z4sSOwQWrj
OPs2+jw05PIy2l7VujYf4Egx7IynP4YW74hTfDazjc8T9d53AASBWB5QCvtT
11vTZ/nrmw2dn7QIdMhFgciif1/TZm2sN+osNaD+ZrAmQWLKh6Z5hKns239h
sqhjuYgqeraLCA5hH9oSnUbzQpgAmUai6MB5rsdAF/XE0U0IHDoqS1DLjXYb
melLS7rPLlJd2Nh66+S8RQTJD4n+K8xkax9aS2vdd49XhgPxBefNxwhUfX+C
I2PGA/TVBKHWf8brtTDebpZb9/71ze2I+UGxNsE/frq+QyVGog2M0f4dBHH+
cB56tKZX6Ta2dQ5K8nRgWdgJ3RhuR7MTxNBDka/SshbMpJ4RQ3TOeFwdTNdc
7wNXW3HcfNpeucdZBaFxoeJTkOcz5xTAQ13T+L7F82wgXSIy777FtEDNRgu/
Rhsh9gwUMwwnQp3WPrTUtHAcsNtHZ167bSZimClR9w5hmjDJU8kfI/JiyHJM
2n55krnZzq8STghoinDRZl9r6p63BJFALrwQd5b82BuJ1nT3/pFBseYr+VY8
7xBg7QNUCAV3Ebwh+r8Cay/PrkJwPidJCYrBVosX0x1GKw3VrQnqQnBHUORZ
VHJOusAxmyoK27dRpLBpF869KRqKW7A8XfYcvsD44/f6aYjexdPv/z+iGpKq
ZNsw28CX8wLmczg27oSXf974OUG01MYLlGBigWMwl3M1H438gJnR02p5Lm9p
JauRrh4aM1CDm8gekG4u+zLdBpsGAPx2QQwkpHYZJENgwbqNPPBM2xj8F5IL
5ULAzB7Zt0RvbGUH/SpfBDWmwupZLs4Oc+nJlvbv9qSVKuwe96uNmA84NU9T
tWBGRxui5HEzeJydFt/y4JGoMqslvvFu0tqDmPXUK/GYflW88WPHz/dt7vAd
q8qdXAmZtofguq5uvEwQdXbJtlW98Uly/Y7ojDIq3vHpbA7gbtvl5zUeJiNm
Bt7C0PlJ2YqnOBJKZtl286mkITP45EBz/NH772Y6wnXIPfpmMH8GhHWSrCaK
w6CyvGYVllVTeKfv+anONYf0LwuX3T3BHdddwdDRE5Oca0w4VSPAodZghdWo
CzJQEDzM7/Cyzeq0v3lCVCg58UoSmUgb68XFSmXUrHiuszP3I6tuZge03RbZ
V3eXezxm54lfYejqi0efvNMm0MOi75sYAuZWpMqjvWCv1KA2zv7Z19Ausw06
++NR1CHwrt4EXZsG79hjxLLEu2DTpw8Ek4P4/JhubNz13gPyly88dmsGtkbg
S1hLmasLiSfJH0LSX/1DhiQymXS4FIwdF18JwzbHSuAz/H5+ZfeMqmfW4PwY
pLE7E7++5X5vpgGMKzUkH6NSRwUb6UruC398K2ZkEzW2Snp4Nh6Y4Q6wSy55
OM1eYYPCOHyeR+Tq2CC5Aq99QxpeEldx5ih5R3WlALjFr/BEqL2TvrpXn4Tx
MRn7FSofvZnoZkgqs4BzHI6AHwwKBfZ+eCLGYVpx6A4gdqW6mtwzw2LtahKm
V6qUEPe7vyCk8+Dery2OSIkWgIqgfy5GBmupAdNwJ8wv3PmY2OnQhvpimvvv
Cn0bGq+f0Zt6XtZUEE4LuptGuGOvGP8P0chGkA5AvJDAjsJpVK8/t9bLp6uW
4svXJ6AHl99qBCHaIq3+5mwt4nsJEsnGT+FNid81HV/fy3OSGCRt+KYdFEyG
oCOyIJ+8oZm4cJ0f/Eq84+xA4cTMqHZM5pJIi8AQCOme1ELFJY8uw2eHWmvI
OicyF4t96CmIrOyzyyXWpBEPF7CTfSptbJTJYgBE+1RwM6+pN6uNgkl0MHnb
O0e92xwDOf9gXFjI+LqGZz5w/jTBKzA34lQI5OOWNiz04jwni82074Fnc6JX
JSm0At+Noeua6mRopgDhlIm+aQrKDjG9z4FQ7yFsVwEGmqYQzV8fA4r7nI00
l05vO/XUBCHvil+AilTsDJJ0ZmEAkyo5vly5Hms4gr8SfoTLjMkIVxymw1M4
sRzTnyBRnnfQIRFFPziFdu5PCF1sEZ0luOS/4in83c8Uln6rJet9PlwBlYlN
j/ZnuJYFrilGDySt/49xOVkodaiYkCiRSbxBgdiCibwWKb2/cno89DLKugFc
WyZC1HNNmB+IgwgjLdeYw8FnPR5JWk8kwNi7jjf6VQgPX1Qohmvei+ooX2+n
nIb/RJNSC1wVQsr2cpgdik8jQkDFXSPHQ2hg//5Hp4dnTyUlMCNMJXtMaP8T
cZibC2CEMSCv7fiZDAMmzUoGOESpYQBqAA96Y0He/KqCCy1tsGijYDgkYzUL
OPvWH3HxpGb4ql/hYiP+4KKx5hA+3SCGLx2Yyujk6fQ/Px1aSqKW5B2UlckI
N8DaOr8imcAm/zc0M4kmEUP2NYegit4RBfdQakarhg0QlXhPrzZcNx2rUbqO
RKlr4qaSOOUCOLryVbBEasUDzDh3YdmWJO6R3RQ+C2ohg4fWUjhurDX7XO4o
fFYvuYewpHIKIcNL8i04bV3dcCsoXcSnkWjDZE44P5DGUEQqrkt7P84VCQVE
/RkLbbdVWvDn1OYZGJYCXeCxcTHoyso47pumCMIHuKsheec63tVfqAJB4m4P
WfgOpNw+jfBSzg1/MIXL7ASdgaS4K0xCRGv3Lr5HA/F2rXaUuKzrDi9JKR+5
ya6BOchvZLxG0cFk52Cmpb572bIMe+rSz5j32Q2iXYnw3IBVc0kCjAynRhVk
ROPcxT0lLI8cTdM5cc2fv9M55Uwqr3PlXyXZcWX3A1GcUFq7wcpeVx4wsWFg
t9gIO7PGs8jICDre4yVjs3sfZqjRpc7J39bMD5qSUFESZKr+22JTcnCyFaTA
xB9+RAEFYV8R13Sa1lZiwEmcCEDSnkDg7OD+fSMp0TEM+wgY7FW8Af5T8CGK
Sdv5EXVOrPNJSdT9WUJrfXeULrvmh+2K7FzDt7SJtgXcOGLLq40jPIiwVl8Y
JEN8ISVUwxLGhCcy4tNvWBHPozX+Fb5x8blTRIE4bOdvPfW47p95KmQMEpZ8
M9wHTgNTdDKWJTGTiq0EGxfP0hnXR8BxeTal3K3rAM6Zn9xG6yoviWRwTXc3
P1ZQ1lKu/x8rUtbbVFgsk7Sv2JfaOtV6vuNsfgEy7stgvGJt8NgjXvDvglv+
i1KTMbOhVmEM52++27duqPlm3TgenQs0XqLEX0+Yqm9XEzssy0p5R0DUTuYn
zuP+Rdh4Y2YuXk9u3rzG4OzCBhnCityczyBS0aZrRxwqsxwhE7yKFYYOQsq1
eJBASljECfV+uAxOAlxL4z8q/Wg61NDQso3ljICadt0/w+Zt+ZQuvODJDqaF
nRoPo5iDLnZB3r2/nHF83W1/ADGXvoFPPX3Z3D4Jju/s4Fw15pkyhiAZTIGc
C345o2lHM7BO7DT97cT6Krfp9aaTnZcscaSB/ABsSMhXHsr3gRCZ/DeEpZor
b1jq7sOAhHu5pqJcRZ7MqktrnxoYQcvmfMoIEZ+0ENVZEAd5aItbN6OuiwxZ
vMtURRktIIeN9fJKVvUBaWEocfCAl5weznrCdjlR3ZhLHzIswnzQSaPhnBAt
9sk6txbaaDGMEYY1cSfS36GczEa1eK8UcYv9PNRjVZXdctxLe2X9IF5F1yoy
OIJRs98naoF8LEEgR5iSmXmdOfIHjiUPEehXTHMFVgbzJbq7DHZBYEuQn5BI
mIWfFhAvJ19O6jMxZXO943uLmOVAHR0KxNurH/Ec3f82Qb1iNX7YSx5CKlzW
0G96E1diqequdFWbNkcvr7d5L2QSpVwg3PumpHhUy7K7tvy1pIXHVR4nDCrS
Fc0XDCzsJ32aYBT9aJwvt06TlzVRpCuGohz5vSA0gywAZZAD7JichedyEnVX
xUhhYA5LzQf77ptNV+0LEZVJi5gPIAWEPI9KcBPqORjW1Fsr8kFdTckWByuE
IrHzr1drcVolS5f4J7jSf5BUXxqKsIZOzIzEpx/YaV8dnkpGM/3YTcex+9a0
8w6qCVIxfbMQtLDc3WC56HrzmuhwLc3x5YnNqSfimKqlIJQqR+keHDfgdZuo
239R9f2NvKejIqJ+mXhJpXlxky8foFIbu85EX3/myQqhijtJNC6mpIYCRtzH
WIdpZxfxYZ6D2mTI9Ti6+dt3Gw7A6lniZ3oVUG/3nSSyoN7Csyckqm9xYpC+
xO9hdnmDwVpzdpWpUoyfwZv5JUwGe6tStAGB+BvM3oD28jzhUjCpVzXEz6v3
Uxs+6JwLaVv7zcSb1qkJS0VZi0bsdsrPtxXGt0Q6mb97HGJVW2url3+UDjPG
RGe5tCiBdXPdKsmVEZHfVuyltgCxXvvrMz9Ft9SsCJb5BXsTB2cpRkUbVmQx
4DIo+XmpCvae/1Gq66wQAVv0FI+M/wrGDq++C2iGAce6XyUtuGVpffuKipO8
6KTWC4gxxLDo/aofDDpJRfgjfR7h4nwXKvZx1MQ7+GhQWuMG5QbOQJVlL60G
BXBZmcT8Zz6IGEkmYk4g/c3a4Z5m2uhsfbtZQLb3yBl2bQEldLpOfrmG6fnv
/35Q9tpK0N/t7K1oL6oYcupg4rNlQp/lnrwU6BhWcnDisZM90MpMFUztrf+Z
XXa4raCscfunB/uVsipD3PbTcgSX8FLllJ06sD1Zd5KkfmNzakchCvkgZGDg
cO/zQAXwvpRVIZLic2RvmlLg+bpR332UPS/pxJXGN/KhsTrczqwwy7aEgbc8
jdM0wzFoEbbF7A6DbE7ePHop9IRVNtOsw3ZckzDHAuLMAoq4VapA/o+NfLC2
2Kf1R5ZBUCG7lMUphRFOtt9ErMI0pMsTP1nW8eMO7SIyNCMw3kbep+wVSlsa
rR/lStKhgYXA2poeS0s6YYl9pouBItRd3QmCkh7OUps65KD2Cd92AviFjqzV
iorw5m13DHpsVZSa7yhgjiTrHjUypSx/piz8Ft7c9UXX4ru0Oj4Lu6/SCbc4
dmCPtj5dtjAeZNtDSPzA8/YY/1meKEydE7R8+A33BPlb4PvLdU5FUXeDPeTh
g1a8Nqt4Wnu0E6tB3PYtALOXNdMW8SfOYC0jDrfZcti0l/cCpRlFGGzRP4jQ
OQqu/hl6SFGniA9iVTRROxV6cdOAGvl5ioJEy0BicYR7Gk+SfiKKZcwYqZDC
swR/bGb1dae+xa+RksAlx/3922pc5L/vCDqKgN67Y5rKWKtuP316t8PyOCvY
oxAyZF7mTPrtyaFbBPGgu22hCZWIuG/Uo+2sD0Ae9KiOSN12fk8YoTf17vqM
pufXO96FTGIFalZh+zpw4kdduqvOtep2KwmbormZdZwj6o2HAqZiTSO1cJwF
DE9T5+/WjAlIJlrGh8tI59bfA7ysMMkayxWfXDGjZ4Mbh9aClb7B75+Ozk0R
ezetaf15rqnlFcOjvLY0j5ffn5Kob5iE5fEaOYnlnmvU/sQdxN9MqYZO7l93
n5Aces9jp1E4JfW8lXv8Q7RD57IPBoxbUZNthDAsB4/eYJHpbB6gBy9kEG/C
38/owmJU5YY7eT+fLzeNBou5Xp3uAd7zIg3W0Y2RZSBifchaiV3s/nxEbpxo
8JTvmvOHMdPSb9ODRKK5/fAq6v+vz3EjRdNWlR26oDwdVMfX7esFnz6/RYt4
keC39gZsLjklrICRchwiTpIjrT1xSSKXApoCq04wkJlWnNlDiwRQg1djRfZH
xhvxkPyUSP52HMr2/QLBcPx3Ff8jXjOF6I001CqQUKSZlk4aIDTbgL3MMU9c
ofp3yDQkyp6Hs46CZh+G3ri14zTS3ayCu5mDtb19+tabiBwo27O9WRipt7RA
v0iLfDxRS4XUKIGWNfCEuxYdFxSl42q37eAKVfjBTtOUHacCFG7es0Nr8T/c
OhpHoHORR6/u47tELHtmsof/3vTBgU6sH3hrtQmraS7pSYM+9RFAYiGSCNqI
U9oJFuQ4faPENgx6gi++e0Kq3ZUlpkutIEFBckQsLCxUuQEiheH9kyBFjI8z
l0Nq9gBdIbMwy+VrRWlnchUyEoGaBObsxz+xgHS7jnjq9BjLmSal0s37bT+i
3QkEj+O/bdBv13mRdf+7maals3LP8F+wEjfmDSYNuHpORlY+pm9XkDuAQuqd
rKjg5KHIAoj6tkeSBMNkDmekjETOVAxqt0Sw0OFd6tT+PyyUw5HN1OxgWxEp
Rz056E0LQNdA1aK55MnrT8xWfbdEadCJTunMJFfhx/v0onz3qX8bNuXQsmVS
QvFYYdoPr38Thhipu44dZeQ9hcm29TnqayhioCWgUzoFbKNXWITpXmc+lur8
0YcMQXL7/oi+aueN84AbH4aDHPmQAaAGYKCZEpSiLikn5I++H0Krunfuf9PL
NYfUfbtzkA+mU1qZ58jkTWS1Easdsr6JblnhfizbcqRjQC9b4G/4Ai6oC71P
bkOaDqcpHEyYu8Oq74vm8RPN+aFfirM2OoaEMiXqenuYrWXexcdWPisjACcy
SshI5fpTnkbQVGafvPVYXd5XK3/HnQMfJVxWaJ7I2DVqjhstEyl2TsjmBXwV
Sk/SaFHKq9Wx1/r5Pra5XeyA3mh1sNBSa64OI3lSMJpjj25Zo+kwxyAM90Tg
LmhZ64uLw6m2CiYFYo8JI+YzE833GvJdodeb2MAw0VlD92MnpuZRs7C80P34
hMrxP/nfRgQrCvkasZrJxiqg+S6L5QVgtb6YjT6KV6kW6gTDgSJFsLn6dDjl
Swz9lRWno4xQZ7PKbA08T1qjxUSI7bGCOmdcb32osdCUZlzEsa7WbB2R4XW7
Hdr1BmkiQOmp4yk9z9L6KYwWQyzN0T4xd/RfYf6CJjMdm72GjDoXUNxCzawI
uJPl0kjahU7Go6FbE1eDCt3ovVt7BaNBnRJ1a1YvkomR7Q9tw/4BRlimX20q
fNRpACbtHhLOakbUZW2hCDjTKFQgKdeAOsXDMWBMWZ8IR4gLAGDQbWIkmnP2
SnPj9h3He5Xya+QnX+l3TnZ+20KRi6CQy0dBqg28puYbuotdeIMnpeencf7/
9E2eDHAtQkLkzObzL1l4QbvFZUEDaGTUFk+iBZ36LCDdEgOUMJ4lReaghBjj
JfkFtFazAUlB/Qs08iFjHNhJPbz+XcXUbz4qC7JxGGE63M+8QkZvPQ271ODB
9LtrqTcPcQmAzM3ZATnvVwe1i5usFmHyZlolBH4L5LQ3CKVidEY+T2CcDaNt
LgOzHBBexSmSGvNRqiikdTyEsPB957x95ExZUGequLGzesE28fRqy5FiOy+Q
kdxQMnbYlykfefuyc3ZzFznN8d6KA+o0VezVjVvohLaMPZsBrsecMjVhCvnK
DZzd12qEklJAtxVh14SWDKK4/wazoBa/eB+CqYJpBUwnI1p75ODPoHw7zdJp
TyRhgNIdLKk9MnUF3HEhFq9hFNNAPrW567ZQa4JFFxBz+eXfjqlhVXExvcPr
lLefCYS/78a1G1owX9SWUV+8uq3ksKsCB0TVzphIPwnZ5mtjFSiZeMIuuhFJ
uirzPQnNazlh+uNIaT5+LzfhiwN7QwBhgrkKkAc3w0+dQM67qDSLdzG2El7O
iv8YqzZOxHe2H5AjThQJ70xB//JH3VMq6NYzstm5COALY5TewoiBQbE3W5z0
LaB7/9rXMG0zWPy4iOS7pyUWDPsuJS/Xbk38NsIk8BPPRRSQ3xBUtfDCX5sv
udTEKBX67MynLNnq9u3L6OX6Z28fmpF61xeV8mgg+fYn/bVBAuqvb8Noiy4T
B5ArooKRYsy26R0AhGr94aEtvN0UNyfZ+FXC2NH0YnMl+SdVhDex2NSEFvTP
viYU2P/p0Ibpqr86a+NFgUMbyJhSQ7pLDnG8DvD4GiDZ2OjUnLRGFB1kbM2z
P/lKEbaK3kx+jYKyg4WPQeMrmG8iZ5JiSQ/JXmQnWKOmZchaN6+deTsHKuQl
gKkE+j1YRpcmC2GYWGrW/nQmNXCvC0ELswC6kGTPb33GIrtVhXakX8mEF8Er
gyka4HdnumXxbrGHIPI4kzk5+KWaEevw4+bSxcqBtRvBhf1/i1UdtXkm824N
WVQRx/r6hZJSQbToKrl85UquG0IfhUPycwIL2kcGRaEIRO43U8oDCqKALWlA
z0r+W9/AG5rv6zDO2gaTPidYQ8LnwbuT1bR3G0BT4YUxubZX9YUDitHuqG+s
+JXXdXHpAlavn3p3/VaGss4hwges5lJ3sPnB3K7J0rsxw2LGOmbMbNhAwCUc
ehqb7B/NaWGYT6bmBhMLzg0r3u69zCSNipxAQ4CRknkzuIky3FaX9w3zJpxv
WiAp+wT9O0IRb4LSs9kgmrWWzNrXObZpAWVYJrMqKh6rKlcqXJyC1EcjkeSu
ZPecAumu8AB39cKQIvdHnbJbBF0KNOtMu2h4xuzyP30JbBMCcFfVZt0uwGc+
HwJsP/H1uYXchunpJD8DR1awZ6DNuGm/mkFLwPWMijaeP4W6CSVRbbR2YWSI
XU5JKw+uGkrpp7JCdLjonXqlIZeGPuLS9OwoY339GDBH+kPjrsnqhDsXg/bA
QyVTI+/Z1FrwdXXRkuJC02sDTm0hK04Z9GYILBSim//ZkokYQXNkXaz+lzsr
Qyos2Z0mrbKJx/q4qT5XpPc6mi+t22xP2vg+jcyKyt1sMqb6Bq6KVg7h4tk4
gN1cjWrJWMPu07rp+W62biXuQKNwwfSoulhABnNa/9Oj24FgV8qiD84dqTH2
hrh7E/NQqFWTYeBiQw08kAvsxWxUWEjTPeKoP5/4Z/oNsaQOVFU8nolY3l9i
sLp8dDAwHkhTAlxMfTouk5odlQY+nNSuXMtviT2MGGlF4e205z+e6RFt8Agz
9sNguq4s0vYg3Gcp4unQ84qe2BCXwpJrIPrzpOyFBAfwFHZFAjkNkC5F4WC8
s35/T/gmn68cfQlH9V24vx8ixT74R6FjHCafcB2vZw5bT4OopCKdIgx2Tk86
ZXV8r1yWnN0RZt1gZuYZlfv/n/dpWzO5+vNZ8Ytyf3DTCfUkdfEqaXkZ0Bv4
s3oUgriNg01kFUoXNIA8ECA6WF6iKG+vS9KhPtK2q8WlmkONyo2xM1LeyH/s
auQfG/8S+KQS4b2VuyIfItsuzUsH7M1FupGK5eb6pYj3WQbkwpEk6W8KqjTc
pCln3FtvKAN7h2cokOdu8UpNIxZljwhnr3tdXLjVN6ieZRxSv6gCii5Jhxdp
Uzkz1uQ2lCYZPIntLCJ6cvPPDGw+PcuiJDbACgms2Nbl2wjUC7X3BNDNCZ5F
Kko5WlbyeEZyD0vSTtEh6YjOYgWfg3Qw4m0O2eubrbWzI8MFvZDTwOONaat7
kV0hCLYpRToO62j7TulnJQdPOkmUKdm5+ZLGGvfSx5e9jUsAzVB8lS/90bYr
oexB2g+CKvI6H1NcgtgCIkZOhZPtSzDwuTc82VroPET3J3UDIP9/RpRdRrWj
P299YEhkIoDh2/H49rsSlTARH1bqsKAVEgQBk5ndP2PD8yBKTaKVZWsQVH2r
Uq0z838KWdDdKnj1noDAB+dq+OIfkdXtDmPmo/K3YFgcLm19gIY7BZiIl2dk
j7ipehpEd348C2Os0qxmoBJcXVKske0U1/pGobFUCVTwYB+RlC6Sb6EpUiIa
IXGXN3TQWbXNOGj5N8Xi5ALmNla6PYDcGLIW0utwX34Efdv17juCT3NPjGMW
Ncmf5db3yIdj8P5Mc1as/QT5IA/lmGCM/tnNtCA3JntZ2Z1h8ouu52vFX6G3
uHZKk1DRkP15j3A668Ij8mdmGA+ddd3pQzEtMrx6X2NvRxZShRa9ptQInrwm
q/I8ab0YWGyFkXNAhP2CbO0Wf+mpnp1ibBoAhCIrhEC3WolhUbphVSGO1NDh
KyjoDZDkxj6BlO8EKBV+aV+dxOi3373k1K37GWyt6cO7mQxHcP/lAPfHAmJr
ZGZ/v0TIzh3i6fuIt9mSnXqKxBBExowvsW1Qfg2PkKNNXjeD7xUp8JSGyG9s
DQQRceV0mRgwjipGWZVRzMb6UAk4YQigTfBGwYRZ90djeyT0SdAnvOCvTKnx
S3cqg7WvGOFrPHa9VDyR3Ecpi9RsqV4aVUJjhTCmpXzVPMubdcb3Kpn+14dn
JETXayNfwF7tk761sNcgNMOVSjpRoeplHV5CoZFOgw2UbUlbrHDtW8DCPkZr
AT+gokDVAKlA7nYEbOvCb71N/EmgPwkpNJ5qTpt+XJ+y9NfDcD3FGc2CvHva
Mmv8zILg/vDhwJSIFRIQP4zX2YYZ38b2/hE9X0nMyU94ye/310tUfCvQlRCS
LOHI/FUy3jn0so2aRVWIQrzdnrROfQCvFSS612a4qPqTWuObBesS6AcVDLlB
s+x5vpALD4VH8ofacD2ZhFPZCisPTHnwJEzrYTa8E9J7ouck4ExT11rgLN5G
O8SJJBoW5aG+YdcKKLM/5Unp08mdX+Q0TaGYv7lyT6zqQeTEsygmQbLza5r+
hC94EEdXNdXd+a5I3V1/7AmqGYf4sCv5ehFHQJ/1NHJoZoCLRse3C9Da9LrR
wBa+mBOOeZpXCF9PCNRc195BgYIr2N3AlUm3qRGgCQBOBvzjHBYpllQX0WDW
o5SwMnSu+hO6byUDeZHN83rcrFRYfRmAopnu3mVO/qe+0BU/GgbrKNAzPooO
DI8W6Uz2tmSEefQ9LbfgIELDyAbC5tBEGELdPEFvBHUIgOdjdnSpu3o1/HyN
/L8ONd6/rk/TyDgeJe0djb/q6lXSeUjEiSro8Bf0v7WDaiMEKEXDSvI/RpZf
VP3RxpGBL3UwrODZPEFLFUm8LNN7CxMTE/NyvLGg9fMlcL/OCSX1R90H0L+K
uBWeDY2ENvHeceKBxBhvcCFUcAdv2GV7mrgmySH7vWfOD28deJWf4UEOiSlY
fmdoTIP9kgpkuGW6SYTvTkUq4b7074vwtPl5AAiSYYraVTe3/wNp3BOg/dlN
c8P4hLg3iobmOkAwReMfSi3Loq5iDyIYMgiLIEnmYlTxwiAzKEmvFrENpgnL
TXw8hz/R3mLznXE558EgYXahwipDVjO5Brvi/hioJx1V+1fARsQTtMFYlaO1
vzf9rpHEbn1t4TWYIoq0hgvbq27aazQGm8ZgUuRCMpPE+O19+Su3ug02u9XG
hY2eKajoVXU/14o5d95hofStI3ausOBSbb3Dc9w4CY5Im4z41B8KDuwpEgvk
97FiWrm2qoxexH4buy66KWwp4I8kdqdO1nUNayvGjHFszneUEv3BUrHuCVwD
09rSDwUAO4vVUd3005vhlEPO1Uq3gxfKGy+HqTAszbojGwvWeilWKncn0/XB
6xogJ7wAOGhFFxAnKzkQt6Vu7UWXW3RkRSVoFlNdQKD3WccrxEaUAasU6hoJ
77CWAgucrXnvBvqqKzvFX7ZF2DLxX08bDkzlhl4mt6b9MQiAGLfLodILwYcU
vxCdepPGEaYaBKsTCBMgKgKLCHXIVPlnDCja4G3+Rc4zNvoR0r1BNAQqYfgm
FVXvEj/TAv5DyTM20+BnJlBfAP62ELUsECqveygzmzeTW8tPbfX0R14yxb9T
YIrx5i/l2yVHLSTBHCKLGq/3kNRUP5fqgPCZe24rYKqZC9dQ9h2/len1gB9L
MkOMt28aoUKaoaOPads34blZPDs7ivXjMipNMrUxUsFyCLwWyogReHWM1kjd
27BFPSVuvyGTilaI3x5CD/4O0a9uRJ0vPQB5/uRWXDyN1YVEhE8HX9v6qCKJ
j8zs15x1Ehw5fS8FWaSuRUam0Vj7G1pl1+sN3Rng5JhEOng3rjEFkPsda4zH
ddbSYy9t2QmCArLZrXx4Wl8kAK7uVfYqKOZdrKfMzwPSiKdACVU4voKC7ycu
T9P6cKLuIdeWLICUUvP0LpU1D6BrwOmhLkxk/v0uWQ2Nq79MJiCx/OXxZqri
4ROgwNOBkXHtymWJ9cEhAUfquGLPVgXT0Ccdv6PAfXv76iXM1isnBgIckKii
wj4fGxvYT8lgxcQ6r4eRB2PbwyyCQJQHCBLLYBD6XOdSXZTDj65kNxVXSrwK
JiGEyMUKMzciU5G4sESmKYT0UELCdg0mHbWJWHSekCYxfac0Wx5K3V24buQ9
Q2/q7z0dvPVKWrwDs6Zoz9eQ6NlvVVoEiyycXeIjN2HSYQn4Acfpt315oDwo
7CArxDZMnhcyjlcBWyGe1kEKc4rZ4of9yZvKKS+dV5Bc9fLIee0URvYlriHT
kd6KRaFD0PP6WEkkrGh22LFANy7DHqbpYLQxZWSeOE2lx+sgb2qGKVXqL6El
wjhITq9/yUJexrHxx5llHzfHr12j90F8mFBqn/SYEcx4sytwAKMo3IBgDcMN
PshbYp5Cfc8bvlVoYtFmv5mr9lEZNtKAbNBtVC62AzLJzxQ6SLgdnJNqVIfB
0lF8Xv/3bIfxjrsmgDqYUKlCHxcKNgbbSfu+ZqxGW9bGvuFUZuKRUfbcra76
+SyRq4cMygRcUy7AA7klB+cq2VrRzShxwKx4l7qer3wRj9OBHp2Dds/YTrhJ
nPBi3Wn0dU8cMAXPG//oyLscXkAPEedAxQ44zlY4ZvOgQFJ030m4yr2mVYhM
CDD7yObc66aMaSfV/MiRzlZQuFzDPCvC5BejAXd/Y2GMmRgEgttYFoNuI3Gd
cwSbuwGaVxDFeBEaNg1d0mY5ws35/5tYoo/xc1/ZrvIhg14mJmdlo/sy4KE3
zRgEStsVDu5NY+dN7tsPpMjp/IL4ajw4146MfbhMWdqpTnHekHiW99uOpoY4
eDy+vFu8EWK5qSsR+1vJC99+otS2C2ePiimsfWhYd+5mF8/+j4Uu1/VS5S6i
XZz5x66MLT2zij1NZ2JWfx96K42t2oPSP72WdHgzfv5TRKcE+EsKIpC1mfI3
uYv4s+IwUOB6iDRlTSgeFmD9bztIML/8slDWQx0LN4a96R87CnttkDFeSwD6
qrQHJubBhUxe49oz9mxb+jL4H6nDquXC5fJBTRpfRS0tx3gaP172bYeme2pv
F8BbPQdraLqZe3EjiFe5XiZM1hQONejMLrRZQjlyDD/NOXtcLqk2EyuWcdj/
h7vMv/xg52HSXaJnLsdplxXwrO9YM4Y/deKOyMliWKYAeN4WRXdlSjh8M7Tz
Y6RfPr9ipagy84heSWZ235Bl5K+bJKMtF+wqIFIMT3UBGYu34KivfK9VU2Vp
vuV5Jas1Pmww2iCkYXxpzUWAJ8hjXQ2wDpGg6EaHN7qCRdA3gSLT6XmCfL/o
YB7J/SV6C7K+tZ2hY+3mPC9HTyWbFdcl32T1tfYJJNKAAwOU/zqX67JqfK70
Y8gtVA9okYydrb+DWQpz8qODR8QDVsYYXSOo5dZR4hxm1Donujv4STfW/six
kVpQLOvbXxfSro+yod0nBQslTz9zYUGb0Xm/DEAaneFaAvVVFNOF4KXuFu3b
BDHjiajchksPRBVjHYmU6mQfkiFacrANC2H+LNXsL0MPbW//CaGt2TTdpi+h
4wJZynWGh+oHmr4c0T3E1B2J1erXrcdwwvwN9TkteSJfXNJ4ptnBtjX/4dYV
BBFIb0Z3Lvi6ZJIrEBeSPKVwcvBmboesBqk4guXBT89rqhPYYhprqsJOf2dj
M2M9hNO+kpDeQK0C/QnhCoJHQJSfspRYL+a+A/WOpV94Fn7VywZA6hzeYZvL
Rr87Xouzf/PrWhMidgTxINdqOoidJL0TOkrWtbs6pnh97DhFUa9uJHFiGiqs
cv/YkZ3ggvJ6K91dwm+HfKH5RyntCQUw5blgkwwZqbf6g5A4mHgv4G5kq5AU
UTfzEnYwHoCmWU1V0DNT+WP43FBMeC7bhvEWFL8N85PHU2tGzQYm535rG19B
HVZo6XN2D3IIjLHtIf5pvYRsJUpnwq1CXkDPZlOKZabxzfseIQi+s+fYjN5C
lyCehjotiJsC08ia3fJaMN8nht4LLu2CvkQf76pfJo15pnFJeOtEtlyf+zHP
RGrV1HmjKGkHYjWlOq8RpgAgYWKOOAL6xCAWEHuI5fl2XK7+gixARYTL4JAC
a6Abk4JCW0XRP/N0nw7WVRiba6klKuCKeDPO2rsONPywt+aA6rxc0Y4A1wAq
ZXoaMkp527yer3RZArv7RRDx1Fvoie0Dw895ZA+imKCUMZfzjq4Ike/noByL
xTc3WDCaKT/CFEvoAcooYxIUoc9y8FnVeheAzxnFs1iu4KJspgkOUdFznSaI
9321BzKYuowF4xkR+1eNGgrMtK4ZB/HBiDpyzFk1JPEFMyEZezv7juP/z36q
03K+B7SllGFkmdII/QqRfaVoiEa8Tc3D4QuWygBlUQ4LLf2+h2htShSRf+IY
6tUl1yJ/kwoEfiThMn8vC3CBXzwLfHgIE8GT91wIBmAjjclxp/I8MaFK67w5
inWWTzdXSTDJlBS0hiMuSVwa3oYJnb2tSf2Gaa5SuEpkvrPv+LCZ1JwrwuAm
Qifb1tCkUm4LB/aMjBexD1sKz1TAisrVsrvkDUnOK+Nng2+hdDiFGVRrGWf6
AqNOF8I7rpOn6Cx9wOPdPUk89191bTryDsQLlbwB9IFdoxcwhYtCCARi7f/k
YycRn+OzTzVpjnx9WzWSiqyzVivBffy4W1XpclYGFX2Kxrk32tbg/cvJHKRk
wp3chZ9fm6CcinjYyo5KBUWXZe3JzckIoW94ArZNDb58DVSWgApMXMdEroIt
Z9a+Hqp/6WGp4Dr74DOt7Y0bvyyw+0mwDYUNsshUiQiVv0qsmd7CNxTD9AuJ
/UGrAUrDdqJJwv3KM8EmLy532/TYMbrUk8oylovOxelcBXHHPfIjJBVvETe1
RQPYCUFLp0vyq8SdnyI1ebi7kZfk7u9m1U2Z7mScazUduuVPpAKHhcM23z4F
7qX1rxEmnp1iJhOSRgm5/IjKRdnc1S6848lugxO0ZfIt0Mh+LAooyvrUfyXS
F5gD9Yf/GMXIo6EfGdN80aMDyl9dk1DpB2GRVN/2FVDM2cOMwmL3Ok8z+TLX
SHYzPngP4pfq35uV/H+dRvf27/3UZkGUiGJzHnb58nccA4o7ZHviC7HpL9It
xkYbhmeOfOAaJK1EduzQafU0NG4w5xpsl7DtabiDI+meow/HfbXOVuyG/QEx
ylCxHTVyzaTupfMLxM5r2IshHx6+ijY1/wF8AnJybYgqQTronKZIdCVbsEc3
88ptUxTPgtkKLvhDT2MR2/yLTpwHySRBZHI81GaVIlDtflDuXb8Yf/B9LChr
Kbu7+TyMA9xsPb9xJSqsCHIfq63EFkz6nTYFkpLlke/Q1xf+pM9ybrhmbGJq
l3DaQD9+JcTOzJfkMYBVYSjP/orSSM/J0/9sbx56TNJbNBnKY5+ynYKCC3l9
UKnytD4ONadqpcnSe2v8kyX+SoXxlDQw8tkwOXO9HYzHfK3fc5+eOhKjawvm
+MPmrl5sm4hOGzVwNDtbh83iwzgp14wbntmHr6kWiv3iEGN3sxFBY1KIJY/P
lgByP7StGcO1yVuek45c+pbb1+8L4MM7MWCQeAYnc8uIOnWEZhuvF2m3krxW
x93S4WFfIp9vdCOVi214WvIDuoM3p6Wh4V27anqrc6wQHjvcPEgP5K9GojN/
WYsS+5LNic3peSB0Fq/s0nhRsgHTmTLN7A6FdnMjiadoIJ5/r48sxfJWO36R
OEbuQxbK8mShE/BRPsEVfPFTiOe2aFJxodJSYeBemOxsV+qIL7RdoOuO8ENh
VxoU8p4I5u7naWlnQEHR3ryrSACLUwxTavLQBRPpaZplSSumtI/z6v9UWR3P
au9jzh6MbZrkBo14XUe3rH5K40XB+MNHpLF9qU5EYvDuwh4tRrEDGRH3K19L
5WA++NMUdL90VMMyf/WXCNrs34yJqhYGAO2NDK+53BWLUdPyT9UwdBcFix6B
6jcClMxRrE0PDz8WclocFXYuuGmN6hOO8vKzWXLDhLKJ6Gf0vE1T5BH50Uhn
1OpQFnLBtZxTakdTC0QxBiXmKVvDKT7BIuMuvb8PlD5Rnb/Ze/J+vD222Lge
jxml7QNLs4aVYk0S9sTUgYkpnIeB4qySnaUB2sFKZLz/k0jqe6YFxel7hBVO
oUMxWr+bwxpfbr5PSCM/Js8sOm1fb2EDEcIDJAaD2tezDeA8U4YuWtsyntRz
ZGIPOb9jP8syCJdqmZM0egXqqyjGUUPcr3Sj9HhCBOe8swxkDPTv2D2KPTMS
i1+u+0YHoHUfFaKhWg9hdleKJG+RInzAxFfMs023iRIqVpSUyQ3oWBYOhqA+
A9iaBNfFNJkLAGl57mQpHN70+IOcb99u5ysGekTZXNji3WrMnfjSNVCGCvc8
hg839kmPtQ6UAPcLT89o/R8qtnOYhIafrziswh7E8QSu2SAVpy6h8YTo4a6i
AtGhL/BOYXYORcOtr1wPr1d11k0xQf87J9wQnSjKwTipknz6xevdJ5HJ6juA
ulbfDM3q8V29a8oJOxTd0UXTGtELgWMnAE+l4bABfPlSMD1ZfRxYRT1steYw
Q1INwXT5Q4q8S7x40noeTZOSTaQe5TXIBX7h7zRKZSQOhjlNu/vA8pkSfYml
hWR+ZBxYmxkjvByvw0gju2NA004TAbVsWJkpVHN2Mp/b3NfFYRVSnmowV5h5
8Ck+Jlsasds6GJbcz5IgI1zZnkf0hHx0VUizbzrRZtXG7BeeV1RCxr4Lmh6j
r/VBaptCSwe1n0wFRxvf9CPPSh8b8WjiVBCVK7OH1euLYDUc7D8VGnBPlgSe
btWORSBr4hz8wUZ5fegEcfyZRQxLGr+T1JaJNTdOLYXd6iizzkYxjdLNZHxv
Zv4639OoximZIM7vnTuVuPLyX5LfWxKfznR5Z9rLmYLxChtZHW52sbW11Aih
j+O3a1BAxl6lYumBYUzI7SEWH1y7YCPBO9HvfgZJTvIo+YnLtQdhRPxypoZx
eEK3kCwXieS8v4qehDD2wyReXwv4ojKg6o4GM2R4RiH/a6x+B+cM583QpVOx
Gn2A+Ly1i1R2JE66XdXGevtTTmy5HFsjCK1x+hi4ucTt+Odd6IbXZprEgFmL
4VIyqgRMEFSFB8OB2+kEBhZ9Ou/HgQsOfLWP6UhDuD915k+WgHa1Qnz9EbNC
B+PMbxhdMADbyvyQYcdaHNnYdZmgKEyfceM+UB6LE5z5lxxH26MaN07+UErG
4GP1h2rf62KkvZfDaV2PS1hGR0Zg0AtDSGb2DoHodTfTR8/JvyrPHWIjv8mh
kLQvrTQRZ8dlXUw3rzAu0Hr0ecA5bbNst3m4VYWOp/FGdZ2/uEtWDWO1+Ujd
RNTf9fzE+3hxb8vk+pfI9ET3ogMBgOI0RxNvLQhhSYAdtnqGpmzx5LDJ59IY
xXJcs7+8TBWKriBIPcZDAPnzi+c8uMUuQQvEb4s5luFA5ne6A2qkUJ1hEimJ
3aWFMMYX8+DblXI0HjwfBz2+vvVjKnJaQBGM8dH94SJEgWNZp5LTbBMiO3Ee
0Fm5i7EOcXb10jXwUdT2x3fZ0B/VTNDz+pwHyA32ZK50aqNr3YT/PRgxyIjr
0vOYRxt/+Svkk3sUf2Ftqnd5KqhRZ1Vr9z23k0rCx5DljtGkVSVfd01/Ujzy
JQ2aqPf3b6G4HLiO9ZczveHsG/hWHGg0DKMXzk+pP5QfCnZrIgbD6khOiywK
hzDiD75zHdHDuXqriuASN6VCnoadVZd9gu3/eWDMOu/82TNfq7DRIQMK0/Hy
7BkNso3FkuYabY0ResuHt5/zyi61Y9E9jrI93g4yygx4H/W46bP4+uFXsTdb
f4u/6rvRZT0PH9nhsLcNVMCWlWPtjvVFV34rQsSELbmU1kQhjV3miCRtFZZr
n+Ir0cEvN2kCD/rc+AjofZgaaQ77U9DY0U3zzeaMfBPk5CfjGziCfCpJrpce
FHvihyhsihY0u3a2xDFlhXix9t3tbL9VyVlSyjHKzIeWkcl8cEYkCIrojCGI
SE8Yu6K657XnN/PEIY/zWY5rgQWfF05Tkl/lYApUBmF1YCX1L/2x4uTyhAT3
IoUSAH77bgV9/rOKh0iGv3MwNzp9d/G+hvgFVhRFDLEi/5bKx9jI7kMOKFSe
11Gn9iZeDGK3a0SOd3gnKH3EL7RqyK5dRaOt8KDmw5fDG3CY17r+/Cd+i5JR
g93G6wS3rVjywcLWtHQnnmSIP9xHX35M1webkLRS9ANzUXgFBx3yriNnKytn
VSLsanBaUIXHmr1F3rpKiHj1pFmmeqvMjD36VtHdN1VF15aDx+Aa5o+zt/hg
gGsPYMdG9KvM3UX/jdLhEKBplkhgvN9xjl5f9vs54maE+xt+VedRkUlNTydE
0O19aA7i9s+yASrvPZVx3GXBfFzWdrqLL3fsiORqNtGs6FxhUmAuBwNBT3o6
n1EUknaznaemvjmllIt2YLvU0gTYi+sDf0fPY4KdnPYfG0uOJfgzAGGWTHOw
SsltNyJZ3+i3inglBQDhjrtmUhVAYdN9wACvOLqC0Nb7ETXx3HYfdI1NZ7bK
syQHJQEYfhT+q7b+3RrF2sq0wBpqLB/9QappJcVLoee+eznGAxyo1YQ/lJl6
3P+ummT6jCLZcBACi7tbx2PlhGIFwUdYrycCRxa5cbO20Ci97IyOc5D9jbPH
S4sPdP95U5mq4YLqF+LRKi6kuWVOJ5/oYHdkCXqnJ+gr8b9QNhS4V5Mka2k+
biaY7C88j8D26AFDKxHbYC5+VYIA2Bn/zEIvbzlXN4l5mh5MNqn8Bl46iQP2
jryi2B9j2dHFGgar/+Ij4Tqnoyfcqjs/mB0I2u5JAF9RSp2h6UJAkMkXiAn3
x0efCZ/EoJjW/XcKzXsPS6UKc0LoJJ8UsXlqmPw4bpb9XeFIQyjgBVRHhMzc
USAeJS/MSDKUb9+oWAtXRWhCMGBo9ozC1eLDxtLG6vvAu8W1qCiQQiR6RYwV
GGkE9ZOFZvIgZAMiI7zgJLK20C9YGP2ZF2+1uDUNxNfmw5IxnFy7aHbrmMiF
TTT317HboyBm2KJ0xCT72ihOCOtOoOfh/vEsZlovn3c5VUsbI/eJsTW6q1GI
aLy04xsTS+vzxXZNdDLhf1lWB+3RuRJWKhxR9YxGfLVWOdEC0qkqusjSFhzw
sEr6osFvaSIpdtCahAdoqfETcWhLJu0lpTM8dn5wuHzSvtiOnVGjrFCtNAct
oveW3p2+GPZef+/cpu/dd2YAxwKAopptQ83mTwvQhnU/rHRQtFWs6+hN55VU
KuRb4thk22oV3hfRPmrRU3tSjot87asxyb2gdFgnrKQQO3sHA9ms1km8b8vt
gfPMKa/kj9Fxf6HZwf8ZawyIHZgEJN3W9NE9IX/cwZpJ3rhmmrBfavcYUNea
fUpPsc4mtnLSVYn7HzDL3Mpr86Fw57+c8UZ+Pa3Z8Rj8/aAYrxF9YcBVPJOA
rzzmTJ0/hQJrlwbdsyzmFvFFrnPVSgytdXUa4yzCAWaFEPAMEJBQ1sJTfJuu
JT6B2IcdrHfo1LZr+Flman/u0KhmdfR0y4fqO6XnaDT9ZeyDViDqWCygGGTC
lqFXHuizAjVtaf8ToAPVSbhEI2ZJ/V8LOIyLS9kKmzxEvypDf8CvKA66Ze1d
rMCO1eELHqTZakVcvmO4GiF10Gn8xKEzisT9hBAeRgU2Ps1GDwi3PokYpsp4
6yFDWOzOkDWIASoc7IBRvpyuWcR4zv3U+/YNjHO6YBVPmA1WqKJx9FRr8w7j
rEthF41F8uCDS/aNZBSa2NnvWG7fPTzszsugQRDthsA2f8DZa/KxUndrng9l
MexsxjZ5xcYD5NL5tav0CgjNNVo4SPPUry5N0KEZwS95FnrBIVL78A5Ks5kh
ptELWhGi5901AoEuwSc4Xg2Tf+ViBElvKYJSoe00Rmntrs7wYN9rhmGCT7Gk
MHs1VBJA3+Aj9+obspbtZFTRIiD03+DmzWCfTOGSypeGoCkCmM19wlJavmCg
LeWXr5rcGvhv/74AADq9GQsF20xcgAuRjuN2p6QY4F+vIjNvbkP4cYWVhONg
svLB1B1mbQ39phU2H/UEysR8chi7P5gytQhuZS3L13RE6OfN0Laf0NI9+Ur4
4lQ7DKZoYIGdZPj+QPZRx1Wal7I/QMcVQTJ9BDl3S7UidnXpsoHjrAQLcG0G
Nzr1XB/HHJTlKEGnNfl+QOSmQ17gApfkN+2K4O1dlaJ08YhrIqEy0LpZu62j
0jifXEzYwsvMgxzlCZpYfTO9qUKRHD3cQdSCVnFlvFiFz8ZXzBCInBQzRsxp
MZa1gCt1vWvlZbj+yJ5m1yLeOuUFx6C2WW4W/dT1/SITtSzFUOkKdF0+dwW1
E7yDPDY6QRa2V7tx6r5QWYp50cV2JWuk3SFAsBZRsg5/UKkMgfzHmxXTtz1l
fK5Y51blBd+aYhAE7KuXIrn3FwBQq4qQBBGISevapJNdrBU3X9IZY85l108h
AQEpFqVp3ZZCaq0gDSLJL+VwSzWamjCIycPwyj8ZSVBqY5rxlFl0fwmgrmvZ
hjIvbUbBZOKv20YXzf/3nlshTHgMzBGXOZdyKiU828AyQ3AYcUEy8JJ9xMAA
DHmQDdznZr+8AJqN2TRxzj17Ic74W2WV2yqSHg+C0t6Y74LYNPZcx4OKPUYZ
pDGEga0Vzw0BnpixkziDtxkbvAwiXNQverNt77TQewrtChxSzDhgEbfYmOVI
AQhh5NSY2963YyTa4tQSg2nVPrHObOGHaEdIcPQ7Mps84t09pPOLi54MgqdJ
s2AnSx8y8gESq4q07pqxm7pP2wekjOmdGsOD1NcEv6kWCdv0Al+Xp5w38/j8
K1+V6cPmKXy9EcoV722pn3tTP5zKXo2kk14dHmEu5UL2jqdRU4GmL0LG5GwV
T2i1hHkGSKmrNxFn5AVUu3xKssgEHEv6RrJ3RAezVNtudTJ14+Oh54lAbwlz
tbGlOiZhfjPrLPuvGSkc+zEQUHIgSHVe7fQFr/K2seaMuXmTD9qGmVuGdpYU
X2fiMs5reICC6GbJ8YG4Eydv4lbPZRSyyDzV7UWnhiEUJauV3jY5b7yD1I1D
bZeCOJyA+31mGy9JVmcsaUyQbzqk5enq+cabGB3fAq7AhDeP3eqqr62w5Xju
S7+f37srlZSX+uEMmMZVPBQQEpZLddiamxq6xgfWLWV9okWNknpVA4PH3v+h
gs+vHd0cYVEqQ+hLINq5PiQNvWVG3fB8MX+C65f9w+ey7dH9FP4QaKzIMk9L
o3wKP0Vk3NzoPcXpoxOPlqpcFvxpo3xYb/hKeTJTqKISzjSmPMs1YIavfQen
JHNY9SkALMfhoAQNHzTTxqNoyr0gNPRF+egFOzRNvkWsg3mhA8LUZ97dvw5t
TwzQFKaIbKYCEwZFxQWCoJ+ql3I2/1kJsIe0trlNv5LUsvoqEHGoiUL7vKQ0
cHkKtRJlITF+sqRJQjXgWEfxvwFO6zYqhO33LXABLn2jNIkNz/BbCw1VAcpZ
5lxJeo4vA85t+WBicncdkdfMTTU4JRdMmgIWzZBl2hcJVfDKD/JYkQVD+3yW
x0Y4ab4we6fs+/X8Dku7AWiMXW1pId5V0yvoLCfacElRu/tCBNhRm9LABxAs
JWwSiqqJBhpPUEzirldny2Fs4nH5lsbsjtr0Gn/Pf1Nfw4VwXkQBnvbC7f1l
a9fN651dqag4KTl+2iNRq9oScpyoJuMW5FOom6w4yt3IwZfwwzfAyr2c9Xu/
HfoirE5OCkSX/wFA9iXYHm+mpOLz74EeXjwV2a6BVOpZg3EEFb1Iuf23qxS7
Boz7s87BtBigQvKNp75kZoQ+JiO97Utfkelijl10xl0h9ozpPPBq8WtQZPQg
AlLTnzLLGrUvcHLD8xZs/g/82eEsBoRHPXQPnqSomJMxWcqD4PyozbOd+jh0
1oaEX8WXgnRJertrxOp+weW2+gzyLQLuACiCu83i77YSYVatAKv8hkqA19xX
145Al+B2tKw/EDg8R6bEXeTwk4KetB3y8fFT/DrE04CEGFWkpdzBkpvcnunl
UPPmSk+xO6151LruxpKrMDah8kK4Yb1KR6hYtANFx2g2ByDJdDPpi27d69dr
BYm0kKYej2wOroGm10Z2jFE6awGlxTweqrfr5Cc1izClzZzvGbR4EhlQK1df
ZdZYmA6LaCeaIqKFFRmJ5Kucbs/yyDhMY8jd/5vQnf5gn17JuLZHG0+gTEch
Zl6SH9R3c2LNmpivgEnLQwNMn7TxNBLVXmQXUgUFdh5/x80OlbJlKiE6yNZG
V8YKsE3+XpqX18jb7MjY/G8funnfwK5xdsH2pdJMRG097o13hQdTXykFOj2m
TL8itCX+0hZx4zB9lNKMbqM9ne78nDXDtz997BgGKgYWwzMCWWbqjC4BhRuk
Cc5uIIkNCvJzzUS1HdgHTNmLesL/F0l4ElckyppoBhPCmVUycPpxQPDIVthh
NPmYSpjO+NHN06FGxK7YbR6Vt+MTOyEukJddmbxKO5xOp/gh43nrUdGvAmyW
Fn6VKYoI99XHWvcSJ4K3puRo4Rm5T4ff6+rrdNkgIpvmQaQZ9IEZqUCFNy96
bFatxYZWVN8NtmeL4366CG96UFne6Ibhv4/Zhyo0S93sRaYatHmb0VneXcxS
pfGrnbop+3kBLq6XHgvku1hHngWcp35NRiZpuzdgh9CflqfzUU7EObZhQ9fG
Zjz03Mpj9vVvvbsS5Q/rUyiIODQjK2gpP6R6EAJYsp7+v1V0WZ3GaxKKOCcn
oi5Q+EzG7tHYrrKJ4u1bqFDJaYTKmumSkLp2t9CD97vrFqwF5iBdX3QgDk0r
jl52Wbo2PvOviJVVZ0L1Mk+xOyc4+PvmlsdYqu4PqnPslrcxyL4FERhDoFSQ
UDoz7vZYZvAgX2ANQIV1n8EAZ7E2HmrYbAZokHrrxohu2ygrnmoh2uNPnnNf
0Jrxc9diMAPRZXdp2mcz5rcO1v97hAiKsO7ouMfnUTMFG57dbdnPjRtP53MO
poPF7TyrV1pzhz/dmNMIzxSipZZD46qY9BkOb4et/LV4k9ZJwWbMymoq/QwB
w7+AzOakOfsrqSUIYQKQthxprOW/A+qST1Dn70mrtl1VA3JTulY4CDXxd/co
Hrg8BQP1qDKq+1c5XyY/rnPtgizey7/IyvyiXQe+ejWV/eL/2lXkPQxCLtgA
aQMw+Bnv3q2BcHCo59FCumLHtzDU+0ZAcBKN5P8IxZcS8yowFDG0hVrtXBx4
yt258ECsdR/CvAiF3/KOnbWpu6LOsf/UP/cYMr/xO1fI0AvycrnYlE8LYApc
2vHggl1K7/23jNtezpQJQSoJlyq66uZs3Dptlvf2qZZBuZP11uG9yd5OZY9m
5GDs/To46j01Tr6YiJlo2MR7/0g+sQlf1P6iNUqNvYCidn2WsUcD6HkKo6me
wRyXyyF1/2wbNLqaK72WQdMpzV5kqb1+rOyomijGF6wMs9cJEXrKsk9PkvHG
MXQobZXSdGVw5jYGD2ENiMhoFSXfbDN4Vu530H4FPkGSgwFwHV4DFRe90g9a
NemAFaQ0AWgXfP/9P86xJqFgoPrGHK6n3icJxo8cuk2SAZtXa0aa9l6GT+TL
XqGCMNm71MPmDOtEn4+XkQcpUmPPI12T7JPcLx0RRCBTNuf8g4zl0WERZXqM
9AHHZJVl73Vzq+p+I7dL47AGaOb2cJkbH3Hw1iLq1+g+cRbd1ah7miwfFUW6
DXvIbtidQW/1zwgct6JCQgxcBnYjk85g7TWnVqM5LrJryAH6bFX22zRrU9HU
gq2YIq21NbPYJCobIqEfwEBOo0RtQtVZRzGuBeR8Jiznl4qRNs1oxtNDYS7m
BUFbYli8ga1Hgm5Mpr2b7lU+P6Zthjux+TkS49J9k0luGNyjgCl5KUXqYdsM
kOEA5tjTi32+p8YOh4zJ0PQIrwCFzBi1LJpb8RTR9M8aELs+1p0mhuJgZEVM
fpwGi6kiJ76jZNNO7dnjTgwpZxXaQB8jWr1JaPhMpiXqgVI4lkSLRwCl1eBv
EFMyQX1fgBo+0zpJiUcCcxvxMsbL0FllVfKke0/Q/xbPLGGM0uFY1FQY81Lf
7QpfO+URK2jcMMmb4yI9ONJxUSnvDEogcPIz7cM2kDaSjOvYvfJd3Q0N1X0Z
7dE2XstfL3zaDe+KCxMPy86cB840y9VrtzycJs0n5wEuSY7DqFl7qmMupWPC
oKuhq4SrXeL30Eb6ZTcPGdw2gtz1/pX7+7IXe4iW1/Cq4Hdnn0M/hW4CR/JX
slwUnqJISLqvAyKGiXK/gFNofTLfLmpv3/EyKc4SIb6eMxWS8pjyhg6ZUAXB
t3V15YAywvn/Mp8egBYM92ylyBCf/l3dWqMnYrc8BSDyGHxbZgj4T3cDvkqq
le7kWiVUpLUjqKF7NsBL4BB2CGYh4wDSWT38UVsB2mis1Ik7ScHNqebFQaCy
SlW0veuk7XZBqFhgF3tZQj54QM4cBvMqZo3+8SC0XKZ+9NokqT7lS3iMlDjR
ijyprLmxeEdY9j+B5QpT4ylLuAa6QKjsTAsxKVdjhIi635BrA449M0DuTFee
i3Nfo6FhkQ/aiB7mpFiA7QNUC1VTQrkztfuIn7Sz9GqiNR6JrGRpQ+WcqGAC
L5LOTrj1MT9CiwUtpU3W14U+kkoOk7333QqGcYSajcedLJ6FvxI5qIRtAkS+
Xaqgsg8e3x9H5pcg+Ax8PDXgdS1N8Pa3xmOOfKEScwWUznU3VOzLkEEEHrql
Hh4AqHzHjg/vbjTSOiYmi/EU41tZXhend0eSk40Tljc9c171PdVZvuXjN4dt
JAf7g6H+4jkCUujQH/PWYXQGDP7G1R8UyG0e8dJ2Q3DLfZykbGyJJwZv+ylz
OurWLN8S8U2YsnLKhyL0Nac9H+ClBUrhCzjBVi/+sm+xwY3Z04Rsh/l4qkKb
c6t1HdgIvWpZ73/ecCvL5m3r3CtrXUibN/N4yLp1YLRuvN7h80XBv0JXYQy3
bMkYIKrwxqqkp568ZyJRV6pPEelRrZJoo/l37pNpol4fFulIW/iz42vJgwhU
x9qcRjhlOCCWv8yN63nMwzzyzS/drsqm6Ye0EZxWJ6cwvGRkcJLy6SaVmXGB
/mo42VrSXIAu4rVBUXsGZDWTfAgG9zoX7ZeUkLz63DuHm//4lH5KkV4gebFY
Wa9UvJZsJ+7cBmjzhhFmq7fPiG7aoC8h5PErI4ty6k3NpOXtKsFfWiGJ9XDy
RLdbZoxSvkQc2WD1iM8UBDmAWtUICtOrZcLLX2/XS+oAlxd1dQ2l765nMBfZ
t/tIgWud66KHJp6cAp+sXHpTE72f2eiYbpzWnJnrVpxwPp9p0UcTBU/rRcim
mddQmbAt1ubOahlVBJ10geH4na2DS33oJSC8ZxqvjmuF94kcfFuW8EMCGYVc
YXe6amMI8tu0LKJe7+5fYN2iFF7lPv/0mmgnn/AaG+9PW6XhY4prACGS1tIW
G0gVb8cB7/TEnHMS0MWol2n+7GZ0Tc+pBTOXJh9pnFrxsNUBB0/961M7e6FA
IqWF6nHcLj2cFrIM5ouKrxB4sR+192J4MM8zlOsa1J+We8gSRhL5TSpyKXbn
qbE6+C4RGhwAHnF9WEya0pgCcDjiL+STck9vX7vSKYwTLj3D6e5oijNWp3xg
40bc7hEC/kYaIa20gSvxs+6C3aw/khpCwLbJTnBkBns0MN+5vqLjlI3a5pN2
U6bzet5sxJFPIqjFud1MYHqEWzeiFP8ovGRBcFdaz9XDmI/13sx2VqnsZup2
tnu90UaWlqu1NU2TAiHQ96m9f4nONrUx3PiE2A7cfq9HIJqg52g8x7zJYUaW
o/EpNty1SuLQdoNoHRuNRF3A8hyqposaN2zAXgYstjXYujqL1hqJxdCZHWMx
tmQuLk+EtFhMmCpjvh3pwLlyIwdaosMdTgfXdhJSzerrWRZLKe5bBbaZQjGm
+YbbuFnWHWg4Ekj2f0JTR3CQL+IoGHFPa1kiTcl5tHzuRzL77NYcEWR9sE2m
897LHJuXWpC+7ainGGKSg5mhIsxQGSstSosiS4XnQtnLjtmTSJae6Ul+tb0x
q/LRLiRTiPRPO8IOgXXnfRN68GC7h5+U1019sSqYplsjwjEYSDsbCf8y2yf0
TWojuhHTgl+dFGnUlKud6VFNYAzTHg5JrTn4HtNxEOiiqDVY/CutlAp067Dp
CnI+SjbhFCtR81WJxLXg3wvwF1HJZi6H0QEqs7+bXCJ6IyvFTOsYVPvcomwR
rIcvZt0xgMD/7yabQXQqwtFxtQHJzmc6/wjbejJwD3bT3zj5YGqA6mLxqcac
UgCNFGxTnxD58O3VEAUZgim3PKjcNzsU1Y0AUryp5DUIqZesyWS6ixmQ1599
ciA0lmoDgAULS+U36x3SobLgH0LYB6dpf79Uu23gv1Ac4K+IiOQL5NrEQB9w
wSD1+e33NXw8OvTQipj3pen8c/YLEy58g5YDHk4/70iaWs7alSinmsjqcJrd
xQci+XBB46CbQwXcRtFrvxcxkNLSesenIzVkd7xRLtO9A0IWb1FI/Oq3s+1b
j7OW1R9RsRO372IaZjnFUGiITRm53QWpya15QbdEla46wkMXxUBCYrIC0U9J
yeNmFWZkMZ/rJNxtYzQ1ySXloL8gSY/4wtuwIwNau90PxSpp4h79jCb2VGLO
DvzzD4n6SLvIrRDU0xPWx/o5L+dnqMzoJ3uKUG9xl6ymE39lb06TP5QSRZGP
vnyPAYQTJxHqV2V2QdpxmdrB1XvCJvXQK8V7xnvWmM4ReNwCYRrJUJWNfwHj
Mke8Hh1HOfWOcn6z6WA2uyhAhrAZl1Xiy9Z7a0VxJ3O0GnQAHIfFjQQPv7fe
RAURNmgBWbbc2aknC7JnNB2Q82D6H2KNAyzQ2p9c1CeR5zG54lUg3otAQor7
iHu1+HfXdp+j++BMXJAKosfuoW/pJ5bihYIsGyJmvoyNETMdUmbECf8JVT2x
HjUVzMP67bfapTFfa69HWUR//nLhSFq3ELrxE3BjYpGmHCMR7Qrkxv64dX5Z
p5LqkkjkVW9AukYKqRzhPJPEc+yUehPyDTygTST4OE2+mb8f/5BcJTc2yG4C
heG6ONzAlvPGSuR0hYdJsjOmocRX8Mcd64XOm6Mi4/cjnt8yBAfcXnPloZ+K
n4q2ME5FYSL6s1IoRqANRoiua6afQDos0xI9qNv+fGu9cwspfWIxoyj04ZUz
klxfzH8QM2Ujv+s5MUC7CM+G/Bzn49ygCsE6l4ATW+25q5Iv9PEdz+wIVHNv
N7edfj/P709K9IIHrMRXIwxhCQQCboSjEMhQ2l2HfZ6pgf5cXEO5yxc8WJ5g
PXc8WEITVeyqSYfOVAvei/yDs9VelWhlT1SspJckO6O/Ir7Y0yJDfY6ofe8e
ExgKWfqvvE23gqruJz3Br7unEDO9jyCkGEVsqoAewlxelusEQWqCno0V5aAw
x8IZnuDUYTjUDzYFaNO2lI5CpLJ6LEX04c6x89iPvR6CFIzj4484qq1BexWb
TfcgPCjimCcLDSWUMtMlJwSLRUjD67KdvjuVHqEScu2Yr97Cy4e+o02NbtW0
Axj0/QPtnoIW7b+OKmBMODa8mbHjdQK0q7N20g4MvUch4e1YCPoUfXYa7UZd
WKt12SEPCVGS7prkpQ8Ie4Trn+6oJMJd8RQ7Zqme6UQNq9SsRFPtj5LSpNrm
YZ+3BIup/M6eDgdzBstDXs2YAH5+wNQCCDWhRLrM2Se8iv9uxU9jNn2HQ21q
51OCj985ZB+qCtrnXcynRR3QPvwU9ul3O5V2IGBVpstM+NPgxY7i4e6GeGtS
lu+nugb3KDKkJRrTZpnXSfnBMXqlycaY3l7ZpKmzis1TKeceIjaez00yiAb5
KTwuaRFzOvTvUVxySXbFdJw/cf8uuaDSK0utB56zdrOpAu0lwph5Z+G/R67B
bdOpyhZTZCqwoXMbR0gwegpktXJosyY5XEE8ErgrBbDsCh2SZmDYB2XcOKxu
5P9JV3A6XT059FHWcBKIlf1xW8SEMhI1cOJs4UX/o+RbVCbAcUbeahZ8hsVr
X3l6uvFqT260s3Yld/HSckYDxgXrNwm09LOV9mCRDyjDZi+8/6SRLJCjW0IH
y+NFrUi2yclv+Jkzb1Kqmx5ObZUUW/D1jpO69avxVYY9P7XubBJoKMJJWgze
GT6xL4n/8em+zs/nVp0PJRU5NuzviUk8auLcPLLv+rmnk5eyzCTi855V7WTm
uyhMnN9DweAXA76tv7PLJHvWBJZdWIgdN54qI8951Xywahm9iUbNulU3jmDB
Tgi52W2aCE90RzdrtQVNmMctxVlswpkZFHmkvXCXDDJ9Ez4c887Gm7wuQ0CI
4DeRs3Vqh+Z8rBjiFkE/Zau4fb8eLIXAPBreu+4LGPNIVffK2bo2oNfzxpzQ
Tk5UJCYbECNOjk56B0f7evVR8Gyq7TIMuCzLxf0BV01WOLYHfMUxjF3i8uyq
gXuPpT6snuAotat4A//knJwfhd2VgCUax4VxO8G46YX+DRu95EPjgs96DPqa
Spl25u7FZm3lJFIvWjWhCBLUYmWjwbFQmySSAQW7b4zpfM0J917uo6eEMxTG
d2IDlIuZlSBl7DAXXSYYhaUBWCdssed6OGGEUggd/xpvJ0/zGDrzwr4iNOGZ
+9TNFkxTybA7RtWaPZBcWiOKtdxx9x6dNEji52nZAOa9uV9NeUHEVrrtJrpC
DQ2GKI8XTR8c0ClChz+19O5QxZsjZ+uDnJvrHtR7aLdNifWYYQbnmx06cUFZ
HzsFQ3RScrX3JPaVTOk0YEVoZCDaZl4HOwcQm2a40znXCPqRYCOKpNGHW08j
DrWwE+1QE8PXENZZKzudnml0r02WliRgssikH3SEfaPDhHtH1ITSbB9LII93
uZOH9p6luoP0lYQlRaiwJMtawxZFMjHlELqhMw7wJwzjaAjk969w+vw5RXsU
QoV7lWc5J3i1+NuYxmmTRmVN+mnzaGKTLvHoDsrKcad+dSBUV+OSfa05/Iqv
q42HAsOBNmCjb7sV4jNJ6W32F/ou6YGJMU8TtF6tLCNdZErLpz19xQaomEJn
IaYD4vHPMLeOlgjMLhzvNmBPyc9X3YRqYqHYzQLqBAXw/Ky9DkZenlrpkleS
SeFwPpVMAJ999ZAm/z0O3x106NAb7JyNbA9HkwAHqU3GHlkNzGFypdCJgYZC
85e8VavagJhgkSEDb2DSDPj0krDLVC3+Vi//xbtoHiDf+o8Vi9HQBCnZSoQS
s9Tll8CdO701BxjO0w03cdDq253n5s0EmK/9th4JXHFJ+o7pu+71tEy15TA4
4XHJ3nruibX45ZRLoPhDQyrkLX0LSc/o9T48u+0vda5Lueo8ssXnkaggCQGT
MjXxoCCOvb2WY27/yIpmrBibo53RG1QhuZKLRyomWOgsLRT2sLX41nOLkLJB
VjAKHw1n1MsIm7EVWEW2RXDE6+x3WOLwxqYLYUuboxeBkEJKbSW0158yRaaS
8MY8Qs7D8j9UKVfx8ZTfgjk8XPXaDO8AYPmBwCroXb/6uX9YrS16B/E58k+3
exfMx8/RRtl3rEa/HBYTdkgGzsDjdW3hhtZCO1JMqwiV++VGZ+Kiak2l5U41
Mx+p+wxovdh4vg1eRy4ktB0z2Suy13Uqc1mc86k+gK3+9xy+bqzNcrN2ljQI
Jc3p2b80jpjFnd+/9ETEiawayf70V3wB3l2ZE2u6EaqRiKIT5gaAOxVd1WDi
UpghgeXg1lVQoAqlJd3NfHw3W0D173W68dHUIzCgd1QL2WkHBr+mIZILzbkV
FkS47wcxyVUrtcg2cJSC+PSQsSX7wn8eMEB/mWa5D3RLED2ttrpOlvYQROdb
VJqs+aOG3EtQIOCX90Is37d9dlQXl1hlFkpsG6D7xmmmcbBW9gfM33ifBaTB
vNjWqb5T+GhOeE1SsA1ybpbpyCdWsvX0zUN/LE7FD0m5jWpblIGJn6c+UmYz
9lv0NBV8Bunc3NfOmCSQceEa975W0tQUEMDCrh+ELYMYZNEgowMH6M0y1jVl
jqrSYklk4D3BPx/Oy4Nf9UhFsifqJ4D4BpFA2ZxuBw9PDVGK2tKbz1cC0ON8
icASHnFlHH0ekt3ziQdGJArqis/y/Y0KrY/Bgis5s0TwmTlWj4at2TZGjSWk
moVHLF2DVa/s/cTGV65/qnisUssJwasrg7AhBDvdtKbDNO4/rtaYMcplkxzD
1F7LFJsQ6zU9ZRdax7GsdrEMuuhFI4STkxp2mQF342HBPkjV8iqz3yB7kLoA
die7DkPouIUr5G/eNw8l3txFxJIx94r18WngTE8sNspqkEUsDdTQ7ZW8hO65
tlyY1MQAXBCAf8dXTBEgB4EBXCO6b/p51wQBl0nAFtyrnv6fL4V3EDHRmv4s
bb2dzZbVxMUWsVrdxN5aPR5XTOlOxgCt/KxTVOjJK9wzedLtIUaJv918lF6W
+YftudeNtZLuzAXoRRmDooL0ToRJw8UHAU4lZUPAtDsPWmAG/afa3trl0RYq
SGT5iSOvktgKwrpO188HO4DbPo+Oe2Hx2/L4p3rpbrokZlk69tnbukWfNCbl
9iLyFy3tCN6DnD/FbvLvUvki1kCksF5YwHoirji1Y5Hv9OfJ5fIAJVb0Bdm5
1gzxmHGbrsfS3MACFe7VedegbZLHg980NBiR99z3FtZu9xrjDK3tVJXcIGhM
V7Tmq8TgYcEKoatbp14m0oaGhgdllp1rKft/m3YyOy+rBjuqLKVFCJ8nIYJt
z/77bv5O/Y/GQMpZSF1ntMpBnofdGwxsdwR4CD//dovJPA/9fICbDp8wu2RN
me72DWMe3Vp9V+AkZ2G9+YEe+danPoru/XMwp9rzdj68dbuSG5biJuncg3k3
n8u4kDE4TwK2AlM/HgYHQJLvz3YRmWs25LCwMfrKOYQBaWzVCRf7Dv2XtW2n
HgmiyK37hLpKcTFkQXBmc4/W74BwGOIDKcBxhwlWSGv1r42gf+kGIba10oAL
i9/76b/37aDYmCyqFrVrs8HZINT7wb8cpbAvv41jlUzcV6JgRykvNENzcdIB
ll/S1VwKwMeR4qEDhDmnsI+nz2C/oL4eqlnFWkpWVzM5k9pDBFn/X+askcud
FFWkv/nnqxy8hYjCkY+KzC9V6S+CklK1+vpn8gki6WkGRtkIVQQmhtplu+4w
lwmXehnIZPwb6IJ1TZhPflageiHr0wfqR0EGfEiY7PsTRCzbKVxoxWvKlfv+
nFbP8uuzuPkHLsOYeB8g6DV6dMNnn8PIqCSQQRSNxjnTDlzuNVE0qfgdea0U
8KGpYqrIN9voirGL5iipPAPYv8IGZlpaJsHclOxcIf/O+v3xO+xDWLZ0VjuZ
U/UyjTdtJhvB07KE3fLknxGFlsQS3XSwi9R1AH0DJ+kmoavc2Zl4/YwrPbXD
5cTInaqS/3yQ+trF6FguE7ggtszSempED0QX83jWk7gGKa9Nfp2FH4oflKci
hdNghjgA2XpeCrhCr9hUJpRLWbO+m+RXa5tgaEM6MeeKl8TlKQvdlGO5jl/w
iGa0cuMEkYI1O4iYSQmrzHFf9X1I5WceK4S/NJL6nJ0UgX3e7xDSHmkkDUw/
Ce/KzY0yzl44Y5DnlOVckEdpvZeNEALMUK3pG0d5h/BwTuzaueYeCosY0dyW
qhzQ35p3oXEvEuPdr8xfU8wnZW8W96o6QX69njxGWzcnqVOUbJRNw0SUG00k
eynpsOpNNmfWlLFouRkTU/WBmi52i0wXYkMOp84fyYf7w5vFnHJAYdKZemyn
J1QlSdaHT7N9XMx5FwpPh0pGdoqHDHxv0jHOI9l8O0vXnf/xMms6QEe6+9kB
amt8oGu5qYHRAgLTlTPjrU+lc3SLi0I1Bt8oA8FimasQy9ZdnBn4bvBtBQum
Ui4/JTz9xofpVU6zJ/7lNxyTe/4NjKfSKLi2KOLBPibBVMyv+Mc5U4URtMgi
Vluyl3IFM17Nu0W/oo0Xif/mnewIuVYRd7/Q4piHt1TB4rI7zDXQdVkU/JD4
5IYDSyktwaI3pMybPzymcmywbmuDSIKLhzPNb7cbZ2WFzuVz8U/s8ztSYYB/
of0VgTpmPcl+V/lwIXEdxnqsjcRYVbaaXsa9505glKZ/Zq6kyE9+JWREpwVF
8hnIFW8YhnUNxGRxvmBJtCq5VXC3DD68XVZ9UFNJq4FwdPZVO8XPwvvMPDh+
qQ9I0IyXWLr4Fl15cEsHBKDl4N8K9lsP/ru+8mCYaDLoyzTlI5N/ecMz9rx8
75U6S7netDrCk9C3hY6q0ncaXlUEquDUlamJRTcT13m8RaEtk52BKEC9eiOm
lbcpa1D5sJsAbiKU2ivBNUoo9VihRzDRsDtsE2SSfnUOXwvgzP7m0ra5vgqr
wkIXzrIVwJZvzNJE4lI/bCSKQB6vbOys6OBG8SC2fxVIfMhxDgCnlLJz/iu9
iLvpryMIRR92HQVARQYBvBPl6haepSBwDsDCfkt1KNN9Vdho6N6q+1H+TkWg
YLLVwaulUzAg5ImjAbKfVpzps8+ijKn/VsNT4tMxAzlFczPNzbzxc+3awG0S
2uwKV6N1C4FI4z95G/lFxZz2vLRZiTKh1o9bZ0UoPz++XmR0SUxtI0IvW0+l
Yy4bShy0sEoi3opEkeUR5U7O5S7LgASMuwKDCebOF6lke2JZLZPND/hBictT
KabrYhM8d/q50AbFM0x7l8G1K+AQ5MZ1DXqPJAwy3EWO2fu6wdrDA9LRg4h6
P36Vlb+az2qnTp+Zl8yXpf4ObzcAsJpCmFC9lCQTy/F9LsMNZhocZXaHfp2e
hwgDOJLi0HF7N2p4mUkfNgjMRjd/RKJYAr0DkY5RHGZIdLmBX6o9WIRqC9JH
zFlrKUyiid6pCfGWLmSOZw5ibAhXkwOdH6kK1U07hBnv0iUygUXOKJ8hgyEJ
AWgAnoaWQjSXWJ0grfVR1q8MsmTjx6diGrdjBWBmDdSF0DuExhl8wJWAPLwi
WgorMoxVQU3U/pRHGzkQ6A0JfR0/46HDlXLCAYIZ39aCPA8fQ/WGUQEU3wls
ZBkixaS0dlDLWAvewIRxK+jqT5QWv7FjyB6I+z6QtY1OFPaskgdpxfEhxBDk
ur1hpkwEjNDlMTOr05Y9PUvy0wLORdVfB+YFZVKIBAmPlUu6nxPmju5eTtGc
nm/Yxt6AtYEZr72+m+Nvbc0hYi1VbBcJU5A6mep2W/LnmZuXOd1Hnbgsp90X
/qstd68HQyyYnxrS97lZucxx4mShpRz6mkITI3weHkrlSUvHoDJerU+5s7IN
00Sw/ENXqhsG5c8ly8LgnlXAs1L+EOA8iIY3jxaSRDt+uZoek5Cb3XALqnBm
5xJsFJIIut+OzmwR1v/Kkg8yvUMVCGItK7RmzVIIZjjYkFLTIqQ6Uhl2eTqK
bmQaJCPbHD4hBWsjQTGEdoUSKSzN7d8d1vdDgamHNxYc+LRS16AKU6WEPiPU
tPD1fImrwMb7Sd/5A1gLwSWtGoydKoin/u8kE5ksedeYi8cyR7g3YjejocpE
+sw116YwQtQ71PokPr9q8yn6wSBnFhE3BCL/+QMdLKCEdws7jlws05zUdJ3u
G3srvnntn/ArHrtH+fav0nR9aU2rznmvZUMGz6Cg+QlLgT4XNiofbyOuNEkG
1XDlUsyAtd3rD45C3nyfI1WkzrGXJ/bPoMQusT1WMKpCmSZehYM5o09H3nK/
nVOJs3z4LD6FA6L21zm5u1HCmEpTJNDVZGTOGcf3I+XEMV9fNGjQtcakyhfq
Y7aU0yhb9vVDL3dn8YffDVrHXUoVlUW59jJ+blB18hnl5jAQkbHVJ5EnjxOX
bFTGTPrXpzIH52nrNCxgZEUaHxmwwINRtFOy51kAX4RB3pM2oWFHMcPumErA
YqM2J/GzU4JLMjAh3EHH78WiX3+eMgdibN4WYDCVJPFmYh8IefcFumsePIwt
6sKmCVfuBwlPyLWqPmDtXo9VthBdkj22G8uaoVOUB9FjeLhd7qZHN0/0lgez
k6MQFOtHyKNsi5ONDBjPDrACXwPHrDL/pkdqLtz3o4ESbEYpJsjxRZzGrEgH
v1YB/MqZ7CPJA2phRKg6ny1W02LhyshOisWrKxzcjCqjQ8iTEy2MkZuYkNjz
QjKGok2/i2Vbh4Dij36cHGUIs3a7qgKZr9PKD7pWck1+fsjVW9reSKXPvdWI
YIjg75IzTXFjWNq4d7rMb5mXuuKcqxadNlKZvZGIQtqfvX4h+8mXs2Fxlex4
8/1vZxq8No4QPled8gC52aY1qlvUbx4UpalACFEqiuINQ/a1dyyGOuXcqiz9
R1EZlsIlw5waKWFASZIoVW+UuPSauWGC+pAD8xx/sDETj01Wb9RT1xcOWCqX
GR6D2b2NMfxU5kyNKIkAxtcukQQS4hGL4H41auvGXhCqTYOZhpkQDT+3I5DT
IEJK+POVSKShvEHfG3WslVAltobYUkOPlsfkBaApJJ7nGCnCT65oWPvsSFiw
+Sq/SWGcWu0wHAuSGSkakP/l2h9N6VWbNmspkBQ4bWNd0ymWIxrz/RlINdJT
7hEj7udsjgyxp/jH/0WJrZdhfwpwBsVmpd5Wjy+VelSFcxVFMkNbtEN1Io+n
dGAC3dhuPyiWN2TzQEzUzgpf6QnXcFZ0bpEPPI0jqagglOnokEkVVwmUyQ6K
r+IXt69/CkxpZkTcpp+myqdierKRzURMiEj+ukZJ2O0WRJt9l7TU2sxVHEPK
3dURjKgn/sM5JJghe8kp4NfnVJ9iz/1YvZy7+MpV+hokVn0bd+zfFKqvefKN
TK/Vyqdz5U7qYlX6jARrJyvlT4WO5CBoROGFCEdsmITVuOlqb7HfoNgCQ+0x
pDjj/giwTkfsT2723dLuwZM1sonCBuK+sQyu3c5WJANbax7/j8fM3W7Gzyvy
+0d8b0Sd5ED+YqfBNjLvJQkzuWCJoSiBUWaguQAvDlhvio3bmtpP8/0kRxBQ
JhcliFLzh8wyBKvFKCCRQsoXSTTCDOwa38mlI1fMl8F1exvAAkhYZGqlnAow
TcuIEN/GywT7Ex62kM+er9IjQjlex9iauAPC0YfYvvGYotTtAqh7iqfa+IuM
jiIb6SJ/NQwUShGjsDRWIgTWEiNswbXhnEEq1bfA8Rwv+ar+XoDmdtlkQnhS
kF3fqnxohjzcFbvcAgsK2ih/s3cBK+dSykj4lyUht577nHxrt+QuKucyySoe
k6Bl/Yxf6AtJxVOe6tQClhIG3VGsRiG3JU7WKE6WNjEJzbpxBRivvj3b74AW
YsDUoQNjWpxYnpwAlp5IcqHtTUAkMPZhf8SZyuRuGBV3iOmDS8BwqbdAHf+S
vqUh5IwNyVBaM7KaPwe+nq/vFtNR7mNUZwvDs9uXjAMdIWRittybYgiV0u4i
/n2rCzh/wunxK2jr6WY/SEsUaO8u10RtRqHz8wUst+KfUzD1xP6AfRRGIhOA
QyimG3kZ903J4m9xwvufblnF9MlL90B6RM7+Uy1FMIB29MwW+cU1/+oq8W8i
2JUSta+rIPBKaoouviLFEt1ouWcgS4wTatCORo/Thgwp4kVpTSiZXVroepdF
vFNDKVnAKBlKUWpCCUeo2D2O3rck0CNLzyMxt95FaVWksnX0ARroIfEo3Bly
/qHJa8qlzzRFRx9TfG7F8ew64Thck1Qm8pWHqEAdY8AOrQt1051RIhDZcDhN
08aX8Pn3xA72kl46PSRswJBuINXRClbTq2BpOMLNp5CLYeJy8KHT6szmkjyk
6tI0X7G2xOsMasEdV/RZhkQQ6xeHHdQixyHaMU6YVSzix/fxgaNJfepV7Hl9
ORtqrLOoY8/Stg4hc3BWobyzEvLiu/DGMTpPgFrwqi+hxOWWjxCjpLogfEkm
vPtAC3CCiIo8oGXHD1rQYin9E8ZU0wDUv8h5+AIISaLNlLFqbuNZRnOzWH16
AepU33aGeKegwLFgjAEuefXKVSSs2a0l/NxLRMFcFXCTwwUODDyCtub0j2r1
NjwxcFiTyjTptVcYG2A3PA9KMlA5Ru8iksgJXU3ACmBOifRPleOCHYYvrHg0
U9oZSUvM69JxMzrfMALYHyzjfswnOqGhuCXtSSmULVqsQhfxDSEJSjtqGKA5
wRVcIJB68W1jl0tNFt22Qi3Vy+0RrYrNDMmA3NY7ePFfW950VVnR2493mkTq
Nh2n4PDFOT5fzWhG+WIHUyFMnoFJSZLOTYwWXBwEuD1ngtNsRgTTU86s8lo2
EoyuCj2YOTo81bjS0TwnWmpEnay6dEBJr+TUxzrxHHIGgsIpY1mbe/v/yhhr
02sW8sbXI5nds8NV8IP0+q4SnSyKPSDEohdHDBYm0NXRTBIckz0FOLC33DT0
7ohJ1lPk+NcjYYO7FxI6DHT4kEvY3JU8ltSupvkwBmuCAac+sXS6LmY2Mx1P
enOZ5JMKMKJ1DtwUyWhHLYktQ+ta1zG86BXYqjS0XRLUTdZ38QePybQUl4AL
7kqEKMetbDGBxg8/EDB+zLSRGxWpX20N6zoM5Pqkg3ANx88WtdiI4Q3oTt9i
Zyq7ZKRUqAfTj2A182Cyxj8cTgEPfwLfpiJQJ7RMKUGmju/0NcinBpKkD6wJ
TraJ+DAajel3J4hcqkuQCJCKBwZagM6f9ZDm/e04tcKoPdFt2whQT06m1S/F
zAK4Nt1acnnz+QK7T7VEuGNKqPyZTeqe1//fuWgSTvOKMISww4PSsSJi6G6U
iVAwU2ssXWt+n35w6zCuxYnNrxdlLFq51QYiG8CwypO2L7Lfcs1PEdZPK22B
fUA+OcpoAXK04YoiPjjbRvumOIJBKodM9plWkHsX6t/fzrmaxW0Rh4Q6c1PD
1Im23DzphMmttWWvgnI5vGyZgMwJTzi8LBKVWxwu5lRyrY0FTB4Frhh/6+en
Vdi+CwOQfjmMAZHFFWEOAc2Qbo8TB8nfJoLdhK2NLombHUJge4Kmm9tu1r9S
DtGLUh0XEE1ScLb2WDsVuquTsLjl4HlYJvOvxDJlmEl76oX0N6RfwHiaEa8Z
zf27SUtLYcz14fVmazx2e9YpsNSP8cXcGKZ/rz0OhaxIu/RMPUwNA7DrqCd5
S6GrviCIb5F37Llt+Wwp+AJA6WCaDjItob83nUtWLKOZod64jyQYkOBKZ5le
Hrz6NEjck+raeCBG3Xb+bFgZiu0N5acKIvuBXilqhzWDiHwHKoux7hUFpIt9
7vsTbP5rZCdRDD1W3p61ORu6LzYAeewU+dIAfzcnJoRQpkKQpc9zrEy92QUg
m+6nrXnUC+U7jEzWWQvYjZDKyyLhXKJZZzkNFdcW48BBeq8Yl6lWqgdJYqXC
fpFhMYL/+nLuyvxigLeP6O/cGpOhoCIcNrRB6dUEJqj05JBtt21V48oKgsaB
kk5o4GiixS7FWYfv8ePrtYq80myNhlf1vpPKwOkyzKeIEm0Uzu1H64ct0U/g
KRLjLrc49Zb+bDbt6/5AcxfIB3NT7EqJY4a8A6lMr6CaPhNhDg+fEr/Oqwfu
HW/iR0QodQ1HXpWkkUJV/mLJ8H6ju3gsasPbkCzsGDay/DnD54+72wFW32fA
wMYu9YzLi1w5N/fyMcVjZ4CIlZBOUyfYgPfEFDofnv8xk3goQQFGlotisdOd
nZRKSEtIM4Kb3Uh4ORjtRZ4yQMKaVsM/qX7IFUjl/gm3OoXhp5PTNus14LQl
WJF7i7PqWeXovzi3wfgH8xDo6Dn2Rogh/UOihbV75vmMQ5MWGpWBHVRAFWLw
mSZ0VcZlCNYMYthDUeBj/3O9j/cBAd2tGODjlhWY2RjMB9fAsj26NS47xcOk
gE6d6oCD3KCd0cdIIfapg+a3Q6wtw0GaoQnvMbJpoQAXerp9G1uOO/pKg6FT
9iMM4GoSOgBXV59AdDVZIGTGR7fZbIhDozQX0Kpx0DU2vHyXWGtyhDTHzwRt
bk/9/ODHIFB4m6ZMnzkb/VnugoAHJdnBPn8jIJGQHTiYuZniOE6pJfpvnPGr
ayKkBOXPyyn20I9majwBUNI3MI/jea4240bgb0Oy0yqpOP7hkyBnb6HNhHH/
fMW0/MfCPI/XHvzwCmzcRo/bQU76MSsD8wdCtx0ZxBzeCMYc5tWaA68OzyRO
pywIMNULGZMD2qAvigsQeJI4ThoYKeOYtyChMZ4T9NC/uSzyYHlabxISrnW9
AS5t4vCkNyWEe8Hr1J3EUttd2FAesdQr4SMT5CchG1vembK0cYoICci1nL/5
cXCZiUVolchvXYDtshI/pzjQOaYgLzOF5FC39VxZVUU0LerW667AIxbFgQQh
qWxLJay/oTLQoiUSXM/XUDFroHu3WB5E1t1OL2fXCK4kpnyi98TAENG+xmty
ApOiWueQOBKOpU4vLEoxJGmNc42GF0+K1kVuZ9APyoo4LBynYHucFY7yGZ2F
EpAo1tF9WqCW1ISKWRMO1XPtaS2gZkKK4nvxBbdIdXGCbtubnRPoPy+jCC6d
6UT/bAZtT82xUw7AiJBpl/fBq0Gode9AjA4DDPfukHWqu9XM24f9WZcAz0G/
yhS2G0/hY7e/0R6A3rhx+dqz6ryPwgdaIfaPgi49aLyz5uz6qL2mnQNa1Ewt
z1XhTLtgkqi+BrRg5EvB0ZQvoRt4DjXBKkl/2uIGmP2yKA/rOwAn7pZvP29y
fWUrK0G9BOm/IcDKQKxphX/bJWSn2uyWqAXU3Hi8p7Aid1iLbDzz0P+Z/4Wx
Fo8eFXb/vErDgY3sCFpIChc2KJ6nrCA/3THPTdeqWS+OLLwwwhWBffuVA5y5
s55Xb7sO4LX59Ov/gqeW9MuX+t7gmuaDXzjN1eCotuLTu5C0BEe0aJlbTt6B
t5VwiQqFobqT8gdWtykYa2aWlep00aMwtOpyW/XgTdQfJF+jBlBcf4JXC/IN
zSmfkJPePIj1ix05/Y8VA7qfoWCdxa0PmLgpO07M1MFK5BibwVFqEQArbJ3z
vu0/p3HiRi8TGSF5XmSzl8uIsaaiPMglZGVgyHzeTHnouu0np91sgICfdPGm
EqK6udzvGrtWuBR7aC5f3+/qhvHVJgZsgjeBv6zAedw64qCkFszTDGvxOMmn
Q4mHV5THYfhR/EXZfXLeMaftEAOEVvkXzzod5UxKGJ2fKif1YzOQyEgaGkH0
pLDN3expLmUWZOB+XnpUM44MBs/dw+uW5mrY0ndRGLRP9kkOugsh+By+IEse
YPSIpL4TVm/S0cfQmxwT5NGGFBPHqZScNzkYIy1SaG5BikhBH0u+Y3jLJQDM
ihwgE9S9d7SOd0WDvdD1Lj0MOAxy/pKQCqJhj7XxKn/1QqF2ZEaVUamladDS
Bmi09KvUB2sVENkrlHR9eBexssq89jVQNdcZBX6Uept62ZT5Qg70L2lefn0g
jLfOFvHCgxAOGW8cTwr98k4PixpYTV2BIchGg0U257DhRo6rwUdyc00qOr/B
n2NOY7XmFgxUlpasU5hyl//ZnIaFmwNQijOc91hgMTbmJzlbzE01sxN6AAkP
mv9JLFWuL1J4Xab66Hq9KzAEdPRimt2BzjiU6d8KBrT+sfKhFnMQhpLtHHb8
7yh8wxAw/lkE80SC0d2q3B5HONAHM34i2zQ23Fc06NDOaULB56IrZcAyOyuO
CNsXJu68PXzH5Ad16k+jdu2HnlfFjXovQ6Dh7ZzcgYlIsblkRJQbE7a0HxQC
BZt5zIaorSGnct3RUMFo5TDjdbCLpfuNU9ZsuYX/JIEeue6OiuJtuQpGz4E1
zsRAjkauX7y0gZA/8N3Ha6rOyjYMoJLWDEFii7cULQ36SxUVbDI6w5UIPBtx
889LrFXpatgYRArN0rtCVaFqCxPRXpWCYiyfGEKz0p3p1mE/8hVCJ2y6tp7c
Hp7geIFpF+KTTV5tjkN1QP22g+kaFuSrs3BRGibDJHZVqN2m5VAkFRdGTCC3
5y9YplIAJw0M5mKNhor/3Bz35vSzzltD7O2KdS9c0fNtYDVkpK3+FqPPOBju
zY00N0vFHREyosmk7R35X0tGNhPqwzPuB0iNBBmJ46XDjNiFnENiEEFEJAnk
9Uqt9kk1CQz2D/KQsArKItwncJ6u1MdwwoT16VwUJUtFrMBdIYPcp38Cf7E2
6TA39ffBlpN9qAFFj5ksgtwjBk48fEkc0MycODLlean3YYDHw/XxGTYAOgvj
31ORDop0scdu0sxWV+z9+H9vTO288JFZem0zfeevOh6Sa7BBM93WBlCc7a7Q
uhq7P5YsdSOmrRgezDDxE7h1vjw/aUKIamlTN5825iFZajofNGMV/DPnPZqk
Bda5lJ8YeQmXi6CohSCv83fRdwuQpbR1O8+8NoehvRhkS0x8TVjeJ/27KvOe
rkA5wNpVN/J9TmJNbMjqcJj/vtNhXF8l/7ozMU/ctOU/HWjh/vKbwTfGNFY/
ePWW41vMaswv9gwu2lomtecjlrroyMMwbj/SgemJ5UYhwFa063rdT5z0kWay
008oIZUg0qYdPD6cun7QHlVYNVUKwyDSbvViTe2I0ctNTeCGEvJjNvdxpqaF
o9EfWvLsteZSb8B9boDcIvAcazukjBBD0iF6yaHQkD/LjpgieIn2NemDtl13
1UcDXDY9j2Odq/RuUsemgQQvXQ9u58f2CdTrtoAHF5NxjOZFTkZLFCi0IoOO
PEalLODbLrj1avL7Lb4Bs1lhwrFUqG8jTxTtoraH6W5b4UcNFqCbfVx1sVjO
k/hUikRHsDqdl2OSIGkWWiTJbgXCGPHOWfpuBb/XG/k1V46zmjxORgzpHwhn
M0YKfroG8K/fg6T4jtomVX9S3qmhUKq0TT/7DRR7y/Xl+5auW5K48MtaJoQL
TaGQ5GJMLVZKKo7rCWmEsppgjt1dQ01AH70SN8vOCFlvFPDpYNfSX01OmqGH
flIhWM5+ItA8ljlKDL95SpfNpcc+NRi4sXmZNWCbvjg/9D2o6y9lmZkfgnXL
kfZT3GPE3c8XW8d3YLRGcFwQ4hveuL7PDAogFyJ2cSx1d4TIPhTumECPWapI
qLU2gd1ksdm9f3Ltu3nuvvmvkM+VcTphz81QPGw9I22V5GcoaY3JD5iQq3vO
xT3ObKHRbuSlX7T4KPDy1UDwzgPWNqaiv2spUJtLkFJ9x9qLIYUX7PkBhI8w
eQmKdLnrQ6smVBmD/YDnnqoVzL3mT8j2eYiAeqb25ViTHXScvoh8KZDM7Ngt
1STZpmh5K8gpD+FSV61oI1bs5AW8D2jnghxGG4M2u6br36z5vHvCwHipi5s2
D210tDSZlpnb6ed6H3urExsMaPsD+DGv/myEjJCoIeA3y1Ulj4xhkMjUBT2L
VHK0pK7hq1AYHzG8CWRsUUlPZzTFIRFOwIuulwzuIaTze9VIwcxtP+7kayID
1h+9ArBMvhK9EDpW61MnFuJ7oPXEBoFbGX4ha8vpOC8rhFzwWAbC/U/9+9X3
nm5unBArJhqtDRqcqH1ZPOO8hNPAa2x6licyumh6WC0UvGKTkqqyiqsdMvcr
qVaWZD/eSUsX4oWB2klWzYzw1iedd8aJVrNmhOxmCB4br9ooTv1qkEZOsJOu
AAXL5SAj45l3++DR156WYui0r6APd9VQLiol244ZuuykrwXbi7BRc2G+UaTv
lOA1NEqVggt2DFu6KMwjgDpOr5Ngbq/WFntLHKsPeRTAXAAJietDhLUeAiJA
Zg3s8NtV1n2N3OaysRIO/8oI8k9s8gNIxQ0aQQGRJBImMr2bTvjwMlwyUr4d
hHsqV50bKjmgAz+c2Q5HFnW/mkFh3K+eEWGq4ybHP0fZFQqHNpA764lnaq30
upuElACmtAs9dLX6rgp6pJscZWki9eslyBzoKV7clJZiVfQh51df2AnTuSwc
RcICNOeXOj2vCPVvFciB4dgruHXWV+M/ut53gysl3hCtpaz6S+fjkDJv8nZv
bz9MJQnrZNNI3edBG6OfTL5AzuCTzgzrppIzkeu5ANtVUDWSY05SHu7YBBtD
Gb3MGr+FPVDMM75+AKwgS6mP02hxKQr/lt8WP6mqujv3w+atMzgRkEjrsPuF
q0ttsnmnbuJM1iBno+FM+URv1pjEkT/LBqbYAnAXHtjmR2wopgo7mNTwMLaJ
ww+pSh6KE9ocCQClgaLA+8s9UxcIUYDTtarXZE0W4KzcmVIVSrMpRg+X6La4
o752Q07kIFqQmFlBVgGiJmhok36AD95WaNCF9ScLKsByY+96JGjwoAonJUwi
Z6Na6C3m0BCC1XYh0ABwt5c39uDFAlm2gI43CicGFgGzxReLt893MgqHwHYa
65CGxlsBlVLcq7nIun0Y3Aab93KUYSJYEml8ISRHL/IvEfFYdCvZv0HQbtQs
nVks0xEqko2AjGu/93GK6aujpoZMxpsOnfLavXt/V2MFR3fNUzsjwpsEPRwG
UrBa4tPuxbSq1ICyOesE38LvD5fy1pXGNIBGWE7J84DARHq04WObaHYcp8cm
7EbeoTo8aC7Cxm3Q5bEJ20EHA/fhmKG9DOurKWPkbfVHLlRgm4S6mmsdAMiD
x8s78stUAXDAJ/tBI2U42BN4Vb9LwVsZfz/+sCjwkJ1OWYr9eZzsFyw62zTm
fjQgg1EzGdrg8FnNyuzBAvoc338kB4QR92o7UsAhT8gNgT1uqZ+eYc5Udr7O
0fs2/TBFpAL+lI0cWARWeQZIhOnUGXUCrjYQpfj9mTjHXFwK/2z/NzmgdRF7
FlW+q+ICGcl4fbuCXM8jOgwHiaPx8lQ2TCv3bxUp0xSoBHIyhKkSiOOr21yk
PSAWrmzKTGHFKGR9Bxtqf4oSjDNKvzQN0bUWkozxcgvCb/J2FoUrUcl22PC+
kirDjYv3dZAaGd6UClc3m0pz0bSsqZC0p5RI5m9V4UHLSPMkLURDRZBlcu9/
NByKcp0Q9G7UbY2qnAZ9D/u0HdJJVb/BCbJAUnsexYj9jLTnjnIwKFM1gV3o
0fp8zzd7JwHahbkt7Iv7FArrOXl6/G9lCZWfW+rnWGBy3ov7E7SMGOMS1G5x
CVOphhmcsaNPcKPmWIVUEg0HsbcofZS0oIytRrqQ4nGFccW1Qfb3Yw/nFI8S
b8Jzmo3iPlbb8CxDlH186Y8YRVeZGbSYch0Fdxg0fnzh+LzW2X1mvODcPqrl
aovYMWx+FvOioX6IASZS0ELZxt5sKGntoN/aIaWSn+fXg6xETq1BBdHISBat
Spmixi9Ofnd395zuDi88HAaasHW8GPBhWHMCR9NAsSMVMjlyUVQQtDYfV1M+
mAaHXwbzI69nzxg0dHjh8Oqkjeazxk+OcklIYJG0zFtFlqbuNBFnjMcnjfYi
koCr4B/y3zqt0YHbUFA+s0Pu5nJFwdRC+qbLd7Zo3hsue16XgDPU7jVt2ujV
hplAkbc6Sa1IkVS8ya1Sji1c6thpzfjkH5HuC5KUlpcaN4nMNhmwK+K4JSqI
GSNVXKg2sEB/x81iW5M5dhAUUo1zz18pHiEMa5Pda9qCdHevH4Fcvd0SYdQV
DBkf5dyDpD9KMelNfQqlveiJnyVbhtvNtrnd/MAe5s5+1bix0Ef6eaHYuSXJ
pEGqWCsS9yyVcodq5DqkZ6eRAoZRSAc5Eizi7JKfbp2LmtmsQEG+pB/1dzQ8
FyeagS8gwuXP/zHGFCyBggsbohHEWt4cowkBFMCJa2ZJyRjRAJb5YUnrH4uZ
I9c0bq+vaa1G0Jqw9hDvi65MDx7dksctn8SyMUmfkgblKp1pqwcIofcP5Vm2
kwFd3vAQf6wg97zq6qZhOeYMrxz/F8pRpKlTTFYg/SLFO0R44RkR85wmMQTK
BMhyNl25nPnIiQZN/bSZfuJk9dk25Dt3zAqWcsQXT5lOT6O1BTp6tkE6L3hP
rmwsRVNia8mCc8MeeWb42LNbLbhAtTDt/zLlOswD+hJFTBmMtAV+1WUOFJMk
esV7SvAXgKTSRRzmhmbOrmerWpeUTsSM+XBwCZDWynEkc0Mq4QoFDo5yYqJV
9h23Ta5ueavxPajJZV3f7TfEczmg4fSxP3Tf2aYUvaflPijA7CGGoA03S9j5
vXaZVUKwM1kKhOKVwszmARqtsgNT4vptKrNNvwEbsKLheG+fKTEViZgfquwh
6TWNHHeZ88AfTCEDup2IyFoRQ5j6RNKP19I4Aq+/jz/LDiLbGigpNOqF3ZaC
fL8sVBwudE06gocjFzw87OwCHpzGoRFozy4h+dGrfzHouxEUMx+3BejuaPJ/
TkdapK5BWWs4ghnsYOYsNmBLP3wpLS3Hv5G1He6vy7Or50Y8MEkcAKQF6WYL
X7qUu93yrzrITkG5l5JnwS09SVWA5rZP2d1TQQFLiN77DuQadSbpq4kXZNpu
4nKbvNPk2R79YCRpgSthDTR/LztSRNkZ6l96EOGMK9fFJDTrZcSy8QjMa66y
Jn7AbQ8IGENYBaf5Pi163rtIAcgnGYE1WnAFuLt0kALdM4l3Ab9KaFlxIaeG
TIg9x5iWmargJq5fkNes61JGxSLadIoQAbwdkkgOI4/FreQ6iAlp+MzEeAKW
V1U5P87d/0ejIm+6du8ck8/N3wPG0GluyP8RK/AJjcr/+WotAyV4BkPLien7
SajXRWHZu4DoQZz4QQl5xoaR0vVnD+wqo0on/05Wm1quo2c7e4WAKB9wXykm
1EMtpz/ocI1vd7ngOb6sslvQfK+YRwWt+qFvvGqmn5McNmhg22rMtrIIGHQt
jbzqYwQiDSuywf8XLMjl+NIAFE1n0cUvhyDNoSPjR2lHl6YdAJX3azBgWCLf
54PoHImc6YwlWI5qFD/HRvD1ErEkyYFdJQAcySA2o4SOmldliXrCDxox3/qv
pYsnS+RzF6aoTHqpK/t+AXphVb2rUjFk0TLFWe0ZpAh3aguxI6z4GQX4KXdN
cys4JEmHeG2De7YYRtaUC2ERkftIq/gCc1BZ9h+eR0JTM9CgHhXEQTbr99DZ
izPvVx9tsc1E5lTyRSgrWVkctRw+z+i0FqivVCrPjtu0H2/lVQaM6Bz6YL1z
LJkDbUlNXPo6IfQESVk3RQJ+3qo7UajnP8av9yeF0lqt4MhRVCTfWonR0gco
uNq8kN2iGhoLXWUQ5F+Nasldp7PCElphGcgSnRhCIx28rLZ6OL87oQqnSR9v
Qg2uIgUqbG/CzSIe4COyntCn1zXTMWZ4v2rHbuuvvXUfL/zUQla33da3NNe/
3fIy0Y6MZwGQo9c46wQLFBb65mTOFofywSCSgvkf6vxflxAm3Goj3Ym4XQwB
MMexYVwWR76lsaOjuOWKHf1GO8rDJKj0UGqhDmwIzhwJKb6sYx6p2LStCHjV
l9fVugewouwDg3Plsy317Jn3Y5HhbmqsJlkYkyCl9ZGt1JkH+WIm90HeCcp/
ZreI52fj3R4oH9hSDAWO2HvPp2n18YJLh/Kdpx8EyvO+dzMLgka6SFXathwQ
IaNoOjdDEPNeEaHPvb8iJgcSJ7LPHz9KeLgqezoombewlYdey6NP9nBBguj7
3A3A8BYZIZ/ea9HUxKg0nZqCoieFPFeYNMSkXMGN6T8k4BYGl4y3P1nXz0CN
IVJrDUT3JSKjgm/qC/CrfEpnnTku919s4uI5Sakumcr4OPsfytAeGI3Qv6jW
BxKH+FIo5SRt8mVmSHt+bTimIqlLw7D1XCO627ay+95PMjkBTRN6mu22Nn1d
UnN6f1s6VWCUc8w1Z+ARVi4u3UkthxJmMT8j/RSoky0On34Q7dGShirHzEAE
3UOHptEJJVbuefreiDrEgY36fMLrvsD1ZaZ4JTRfwbyw4YJaWwkgxD7/IgWo
6vPteZ+wVOkOZElvAJBtoFeCYIgzlh2SJOThn+YbfWu+zXeaV5nQgh1+KUuZ
J9qdLzwY514TQFwCvbk6wV95OqjK1OgYElTqUpV9Y6WLwFCXbWHAslvxE877
YuKB96xmJGs6IG6h+VKtWXoIUHb/V1KPRn0gkac2dW8XDgkOlWrd1cvZyfuK
28EAwbo+2o2VOLQQOQ/qw10JC6VDROE3RDzgmtQkIgay2l6q8TPMAsRQ2gmg
2KvjE/jsfkTqzs8jTTAmXt5e39GL+Fw++RJ2PhmBZ+eAAes14MB0KGgNWqV5
FeHBEB4SOYIralPqbzVOorAZKINFBjk3KnoB/QaXcgVzcy2uUhHGcbQzIC5X
W8omCO8dP/+F9ab4wyvkDTRqdvY23XowpT3xOxKECEV7toFxfmnKEf8+dliq
O5ugTSzsLxQ5dBzCIetfwDjqBjAvIAgyKKdx+Vf5jZp93M1L++kVxQQwHUqQ
skU7tSrWHh+Yi80HabEBYVk0YP7VKut3eY/vhzaq2H2MOiAFV2D2m3BkK7vR
Unsjf9nhR9Yl/jtsGQHTk5gJVub23nO125G5zUP1NYGngtbKIgzkO38Utacv
Dg0JQIvnzOpjaZuqA0OPtDzx+KJ35lh2M/ILz7CJxWCJfbyAUhPSpl5cCOEF
SpsrfNZGSGs1V+9Mtg6/n9ZkCbhl5CgV/WGOuuGrHDKjCxZgfRigYlC67Fs7
GHGDXEVs0ig1wuiCkWX7UH3ZHV0uqw5/TZB8JaUOufOYhjbYiuCGvqJb6oLJ
MrdZkWMW1PdACnc+N2YeOK1w8PrH0AZklUzOnW/O/UD0bcnMV2X5BgX4lvIj
OclkWPfY8llw+ITYBzGWrBJpwH2//hWwrRVgKqNue79TivI1cWE1dVaffm6S
FebCmydUM1Eyfz0spC1jcuSgBOfTa9ukhvG59TfMbiP2hCu/avCdDrG3t99m
gRjMQtlZc0P9CuGn8BsmGeqNqMnx9p4nuG9j1O/AuZd+6aqn6bYDPCHar2W2
Hm6od5BNHMIXpg7qRWbtmVgB9AHAh8oNVT+J4IvjLIX3bnIqegw270rpDhvS
uqDmeyviwgmOlEnljRNYNbdPJmLQnEsMFGcYQVFdX7pZtAzyMRYU4AyAFEMM
wJNhofebxSKotlVbbnSgFlSfsHOnRF+OBU1khifvmtP9tQa5QLbjTXbgvmw1
7uaObWCYGUSDmhoRfajeGkM5OV7134TkUCvCH7P3kvDRxg72a/05/cTaO4e2
gop2L4KLJn26HCTSuEIZkj5SgUaFbD4DRKYEDlHAGFs9sPkQsUiqU1iNa+Xz
OzqOiac2JfLAWz8etdmHQODTl59GA7GQ0/lxKFA6ILdECHhSpThOTxbx6iX1
3avyuf7Gbd/pUhWL5UMXAjJKJT4/uZAA0lh4uV+s/mki9YHLGncecc2JYL0h
FR6dKBbYEGwG5ijN0jQ/hK+W/LdtgTsJqJkuZfKhGtOGRubCbJIPTa5gqYgU
wJP8VnBIXVkgid2RRe+EwUlMjEgWQ0MP3Fls/1o4xoJP/nWDqBpO4EQVOC7S
qaT5qpMG2pXIDLWHaTbC0I07h3ONupZl3K7FfjwPzPaftkpreja+/LFO3wAc
V9DSjlRMZf6kOeAtSv5lbqdniRzD7cBvWuAG1yfrWeIvuvxtcdKqZvlazXPO
Kx8cAdXSZWsclXVwRjpFu4vrJngQYx+RJsk/zPJcO3mK6aRZ7GzzbHwfTnZ4
IvDfoJ6HC3pbgz0g1o40DLV3C+un83HtmbKGAqjJcAiFGTEhNnCHyZS/pw+Q
o55O04s0DtQyFnvDyoLdhidHRfhPhB2WbrsV17Pnc4S1mFX7SMGDMxdIU3s6
a9p1HgelgfWp2PvBljUi25sv3MP0CbgEuvpdzJ9vWlneim3K0bxy9jeIwo7G
ZRFRk+GoeucyMBb90RLc5dS3DeJB1iaflgPaoTC9Wd5JgYLBVwmLeJb2jm3f
YW7KYT6wy5Xix+pZ2YB0zRunN2w41yAlumGy9Oy/98A/MbmgLbGpxD4FCu+4
YHcBbBnIJRLisZecIqrpogvuilnXgT5rMmMc1E3/ojlTaRkw32LpgAT4nF00
BGcaUA3Aj5bOgzS2lT6R9fYHzHMRknKGVDf7eIQj5tcudfCnJS9zQlmnNh9y
kQMt6sD49QMazUM6GHVE2yH/3Q5/FTPMhKQVURta0Yemh1e7EeiAoU0/Roa1
Xl9PfxSAaryoNOVSfKhaX+NMNeaI1UF6dt0BS9cclvMNef0WJwOO0OBZ3N/P
VIyBjr1Je/0LkmSaZguFWDPcYbsWrTVjqCSpcDuofJaofKZnbHgFKoqSeGXM
ewFT/nrzKBtwhF5OHqIa+42V6D+0OUoTHpjBnubkifbCZfx874SUSNS6ZlxV
fy/cVI84D/SaWhkAI409Ey7nRmXdc7mAq/2KofyEm0Vo56seZhhtY76EDi4m
qQfdIkzaCQYX9/LnuGPnH7sUHgTT1EFOZacFHsaPx09GkKJNpMGZow6uJbhR
TU4BKiY/Ko30f8RV2gmUsX4v7E+R7YngqmOHA+UZ9RuoHAVSsIMb5T8QQvuL
YynrB1r9G/lzwaZoZzCxIJFsiC1HUnjex7MtkO1G3h/lOuOQr47pEwBCWm5k
YGZ5Qh+K6/37TLnOjzkkGRmng/KfznD0OnmWkiDTpJjRems+NLk14n/yVIMD
2mBz16LsNf2J/VXQfNr3YZ+llPq8CogqMg0r5de7JbYxsIAFRng5cLCytMck
0Ig1TNsEojFKH7QQD+ixidaq9t1abFL0JuBeO1NscmbWshP03Dim7Hn71PJl
p1RcE+uXlV3Zt2T20cRoC5L4cpFO5BEBy5EjIQOiz9GahtKSPoGL/7VvdyNu
GUibCV1BLHeF11pnpnhtBnfYbGImOFaLQ4fZywan73G8dGqHBIrIyIej1Xwy
EWXxlu2fm9O3xaLGYZ+WzFJoAMaP/bdckR+CmE/bBnRLeHkuZbCqEFJnQJoh
wC+8bG+NIfDa0WeqqZGmUNhQcG/+3QIayTxqtQb2NlmwR7+mfartmk97OTgf
7F3vw+SiykZS29/Uf3SYTlEhXy3F33uEocWuTVmcs+uz8s4yp6qzeD6TQLTS
uatNCHgI/rVR5U0UAzU+lyXuHBLGcTFJQxacZygppgOfcEysvKovFKBV2xXC
qXNz2EKSIdE2jDqzG3pXIV1h7lHiDx2P/5Z1J56hbmYW4O8RSKlraH65+yK0
I4HiKnVkZHoUi6cybbfQfeypIPOP6+dXsJrXYGuGIsQLbXuZ2J0EKYhKbi1X
8TPc0Nc/OKV6Zz7425tUzclf+ShH4wDt9K/qh8m2cWyMC9WpDU4Y05Nvl9yX
9luOpbANlg52Rh+0qxGWiGSZZ8tHwDnFue8gGmB6YmphQj74tEEHnwtH+r0a
pfJWj2dzRrwuU7TNfTrDEV80jGQeoYhGrakzopmqsLXf+hSmAypTLoGMNiQf
dFERkp4QJ4yNorhNPTmvlLWEGVXR0FU06TAMR3uJ5adeMiY2nTV0uAc3saxC
P/pQ5WfYDSPZeELY1AT7pynXzKiGKsm27SrRhk/m4XMJ9GD31/R5LoLC6sjf
iIEuCHHy6KPRe18HJtpfjvswroyiTo1rOroKPlaKoydMAdy+UbQAtaH+ASOj
recnTfJDtqWTOjbzRJSRK1SqUFm2C1ONqpPYwDi+cVSQaC0WV7dJ0Qb4AB+w
+dGBvWIsz13nrQT4uFP0wdfsbdAgYfgTNnQQnT3zxApT5RNWxAType6zvSxe
BPL3VwAYmMEn3+by3SYXC+PCkwXXMnFapkZktg4BoZEwlkX4y5TWEPE9iah2
ABgFXQY7htOofgKzPcy8k0GpPpr3aZF5TYCvsjooK37r/CG1UWnoYVuZuNTp
qvRImrqeCSXrvSrWEqAdx7YCQqPRR77pbnJhbXjeWBgfCocZLpXiiSCO8Mqh
Vlf87Qg+FD1/sRx5sR+hidDjnogLfpdMWkNnhXd1WQ9XlrzAzPMqlETqgCWw
56HsGyy4tV0p0GTl1IAFiEFc0pmr4tGMXDVFEkOFQbBKWr8w0br00lDSbiDR
IU/b4UG7Zrr0wb6h8sMirprLehLWbb7NZz8PVWPlFajdQZKpvXxM0nl/W8y3
b0MhMEJVCbP7BfJfyAl0prFOrVnMhCf9fWTL/AckinVneJS67jikTjd+rfjs
sx8RsSWbv9Z7xMKmojS+REab72uibZJKiHT1LsEx6st/Qq5BcuYMnXTdwukK
cNLIn7K/r/LUDHGuatwH3iDZhLhRmusljdoUDb4dsz3jWzRouExcC3pPGP7s
E/1s3rpfthiYZbkQ+fhq7zmf/z+5b0vrz6YuJkUdFZPBlciK9Atxn68tACNv
TKcbPFci3qZRSbSYtmTE8PY5bPe9m1Sxuq+s2aoleqaabnidVz4nsErB+rAE
0NMnN8mV+/FwS09/4SROsyH4U5ftsLztNpXyCCcfN/UjA3DHIuq2V1uNLvqx
qXpN1Al3rvHxE+ndVl6ireGY4wQrrQGakQzGMluXTrF9N7pFBeTYEV6WzIgf
uragzXLz9KE+kcPIQfLa6aeZ1DIUehXh6Y13jXIf15mPQNAmf76UZC9HEdgz
2tMLD9DBNeYgip3q6ocdGDH0SkzuQMe8hkHxDzCgXvQf6VHFYjMa/bV9NkhD
e3K8LsmUuDl+9TskcBXzjjBMiNqx7Z89YXx1BpSDywPxR38axv4FCoFgdQvg
WTVvzVwrqsdtAlmyEDoJ4QuN7n+tYtkpKOq282MkbNtyb8hduJeaZ0hHxjNA
VIT9/UkY4WBPpQt9P3bgBUaOqJ7ghe6MctteO/jdo1VKoMQevgdI1BR7275j
xvKeGiakF5uWhM/WIBXa0q+0wW/XCGlE0zLi5iqwoYUDGb52b5QANFmxGU5M
Ur4Tf+T5/xElmS0y5qUF0TNqkjx8lAuHIuXTjJAG9hLT17vhJGW86BfyEo7n
4Gj++bq7n0dcWRNPpFohN6PUDtq/3sXW4+0emxHVkQ6u01fN2yrWCz1qqTdc
jOd+Plv2KtpaMslxhzcre6SpXMWsZ4NOvj5RoVtqXWpRl06vAErswa7mhf/u
14L5QHGPGMJqHnCdO1w+3siNtqKfKCcgRbTZ30cB50Nu8bSTPDOamYVyBDvS
oz56tdUMFb8IzsvBy8JAz28PPYnaiskB16xehtiiWCt+3uWqhCvtxupdqWbC
aLTHeUfPOe+I0aaqZrwkUFxXtz0mrPIuLEDQZNqxVr/Q0tHGXRSCkINiSz2C
uLZDmhCkYW300eZUuD/sOxOC9TqzQHcl9DULgCmnY60F9eEDorK6JNzQnvoe
lxYvgUuRnJ6gjCyNBr5GgwZ0vi05U0yGMi7LGppKvdzQGCPdbZy9M7O9wnQ1
Rlh2k/urXyOJcBnLBFgpCiWi2o3QC/FtG/4r24VyfMa4sU951hL4f0JAW0wq
xu9Kd+IxSBvl6ManyHLGuaq0MdiIMYfYjQ+Typor8AX1trBJZoxjXj2ogqvG
xPKK3oikZUWRaX9IUJwTlKEcHzLQKpEtnsJ5gcWnhJ1/GdcQwnqnUaUWYvWv
RPhiSOn8ajIdEiz6pN16euUX5Pw3pX3h3hDMFOSLbjYHs6ufm1SSDY+6M11R
tgfE1zXaOKnCFVm67xqXwithwv19sNoL3/SgXyFPivT3aRZEd2z0wWI64Rf+
Dj5rcPj6tNBsDI3ZRtg6dNkfWu1g7XW6QZw9oe9jNR7QxC5Sl1FH/HR5I88L
+hiROCOxPH3uKBjZBRjCm8Q1JSAor8aWAoL3xnds5CJLKAbY4e9kTZ486R1Z
08jlfCwfZMBgK8P/MRUX/zl4WeXg0Q/JTrDwi80UME894cBFepE01CumCbxe
hfYQbDWfRxpsDlIil1f3YRNQWJjQrU+lY6M1PdOwS2386/ijgZFd77ybRktL
si+X2WoDtCceT4mAI1j57axu2hvWIYiK2SDMswOcTO9HRzCm1PsF+WNMQ93d
Wfiu/jM++omwrg9ugdt+cEmDqOsitfMfZaX5BdwqHaV3QWOiUNUcwfyxRIxI
k7Z4Rdrd4f+H2vdPw41KqfIjbNzSXZtoXtD+VUT1F/2lMtrWSdmfoPi+KEzX
hU5up8mnK7gwuHXFSgepL+plXVPCDv6Bz1fYD11E4JWgY7wfWPopIgfY/DXS
QVxTQUxu3QPzrcEGNAojthvFfCOuBxi/r/z4IutCeMlboprkxTqfcm6htE4S
3vOD4++AEpOOo7Ae1IpfdSYUmzQwtfkWJZHGBhZY7zJ0hrX182QoKYl9ZhNa
KpbtNr993puV1HfaUWyGcL0gexE+wr1WWMBVRlmwvdky7LuMnS3eWGj9bqhy
277ixvhRXub8eIHnqPX2tbkOTYH6OfmglrOs25qmuVuU+zK++tDv079LYF/a
CRx+KFnfuuK7VE8E60kL+mJkpW+fyL7RHOKWSEjREfaaz9DhLIOUq/D1PYqX
ZUzBaBVP/i1+TF4NzaDkUmpBEYLw4apFUYjPWDonWtoj9/cNujJ3MZ10K2W1
NRMBBPX2pPvjokDYn5pJTASQkG0lEyJmeN/ChBzNPFkbe9Wz3T8UDmBqVHT8
/z89sqZpMjy7gVlmRHgbJYlb2psaoMwkUGwll/ZTr0nwShxgh+iRO0msf6pQ
xu4kg5WDLFbiEWLxFI1HUHrtQHAYPZmo0aQXGtK9tMNlaQA45P+AL4PvhA3r
WyqNZTW5O0FM1NlGQ267sfgiJj32HjZ33f3K0S53QGY0PMapEGISj0Zkb1/a
O2/+EBSjjnWLnYiALXrAQNUyAiejz1+EYvJpGCTusB43as7bfsjsVMIZVkvM
n1T6TCrkU5LPtRTPwpkZpiHEkFCj8YjPZDr4gTJE0+qAkJU5YNk908trAo5i
6IlXpFVJwPLnAIiqMWfu1/OKzatwkkGA8ae+oELrIUWtD0v9XerHuIOQE3XZ
fcwMr+yBnsKzxhA3AIRFZhwBTslMYEkwUorezFP/k2sW5Z+UvCZAE3pMtyrp
sXoi3OR6Z6KZdQ96axYPvjvqdV6GdrqEdNlNGPapAhQVGFDRpbCcSC4VBkWq
7gjFTILZFj+GNI754R61eT/rZRVnfe/QRG89/iDmf5a/dy3uUuJ83XucllyR
nqr44v/zQ8/FBWnfQWzW8y/CYH9FFfE15AF/ii0KZT/Tz1PaqiOdScoazRv9
UzSVUXmJLNpQkWy0fCgts+WKrPh3ljUsKNY/XC3Cgi/gllq00qbcFC8kQuy6
z/wcGsRsNN+FYkrvc89wwxW4UgnlykE/si415Ka+7bwvloMOP+DRZMLYaYIv
LTmFU7Cw0FHYoGsPBxGuVeUsx1lJjj+3TabYRLrZi7CcK17G2QEik46CHETL
tPeUEXF4jPBYMNT0zQA9BhBSjBkMcdC/eogFlbQod0NMNAJpsDRyzCSa/p0G
slKmluxHo+TTaEi+ih/DCggKyCJRc+xMMJhXMtjzUIttHRrVCAGCJ1bv5DIs
YZCR744irB4xbC/rTkNSLdmxpB0Ri1RmVgmNDoXFKw7e8mg5YiHUDZsqTWPc
h9ltR9M/3TAigC69I5s5lbKIMW8Vf1Y2IDurGMxdhyhZHry3A2dogWn4nrKx
oVHZFa6IYeHJ+IgVYsef0hC8454kjL5mbVUoHYXpjaIvhd1sOoD5FscVT0VH
x+umDF2hOML7aahyPXzKFvBh1MDlva16+4gn+fSDJujhWFt5zW/Peb+R6LbT
uwCcOxMH2xl8MHui/jD0zSASJv6dVvh3hB8bbKOynyYICP6ewdi5a+gF3LaY
Yd5de6VdeGLbTw1/tJPSN/nEwX2ImTSjjW3N9R+r2nm+nhmZeHKT7cmw9IRt
5lM18Dx3FQMGswgLtmbFPMDvTn4CR24S8g13cMIEFMWT8WNybau2qlKduOfs
f2xzgzvr/J63BB7asoI/YCWgxtvqHOfk/E4BY9uG3gQF6IrFbNaoZS00ing2
qS92XMLWhzSbEgGFxiONJfXfugoCXyT0/WyiypSBhajr2naRDTVhTLpKLj9x
lMh94rbLU1eU1/LrqIsKNOxim0Rh5thlldbvFnerHaMgqso9ZnMszldqpBrY
mJMGttDCDPPyDrVWUifuP+K4mAoB+AkqSBFzVCNvvJjFuTtDP8AM09N5krHP
IOKddFxKkkpRXJ04W5QYHlZX9eQ3fIdKi74yw6L4Yrz269N0kJKmv9TJHiJ1
RNBAwL9GdEHEGv6sEjQJ334lcx2qr05tDODkG1w16PGb3P8++aCAA7V1SFg5
SE2vD5v1hawHO2yd0yPMccIthudm0JkrHvtR9qGx7lyEqaFzcn+x0OdP76rA
C3xAV0OciC8d68d5gz3oUSdy++gLQr0NRigVqG+mrp0n7/nLaVy/MAN5mpg7
GAEaS66wIk5z/RWdf69WMNMEXoU5guSqLMKemRaoBDClSBqk01OkYrJnj7q0
Uqgsy4jZrKGCWD42kY+ut5i5i1FiX29PkimPj1Oy5/cqUquQ5Sfnn5p2kc0G
Bo8By7PgZKLZg/W1fYeLUVtht6kBvPccyfs70pu1VNx08pG7E+aVmytQnST2
R1S7EsMg3NPT9OHc8M8HihtkFfzXSnjfdJFm4Yc3nfJk+HeKIuD65unFD8h2
P+2Yj3p0UhUba66ILdgMV6uwoMwjQM237ItvD81Oqq9x180sFcQ+pLmbEaGx
I3ZcofMP1hjCGsoejTI4JUU6EnsX7Rqtb6GhXXhnqqWHCq+fLVQ3wvqH5Dpj
8e5annBI8C/rOTWHTk7SB8KdjPantbQBGKhZ+64l6uzbVYlX1va7jGrdqImp
GvJFnfWrdsPFYU+XKCdtcp7ndjSsWLnjSmbqGhBN9E5W6T/bU/mAA+rWbjyD
K+HOuHOlMyQZ+OxkyFPI699wMnmKxaLU/VSSOT2ZRCirNBDNsqZqbP1RqkAW
CFhPWbsb8q7nV63mbJ1kpsg+NxWDq1qIsPuk4s9BusJyAXL31TrATOFYIp+w
6Pvof6L9WoRahyY4EKDPUkn6COWvORH1msitCD82Q9WUokbZ8UTXz1UrsmDW
2EGRqPGiinryScuunfhQ1Blup8Gn837dSIErmiUpXpPCrG/0t0ev7HGD/Azu
+s+37+dqfi2bsAmQ2GHQNdTJNJig4WSA6QFMraRLCKyccNZ3kU5HHfUg7THt
wjXfFqbvgKl2kp2K/X9EejhaxtAHVVDagX6fyfC8ySaR7WgNU3pzXqT3n+2x
CZW6odnS53VNBRRYNwv+ArSg1z/t60yxLalvt7CilHPTk+DWqjcwoQGkv+1W
UMRNIu/ZX6gUfJExruW6xym7r01U6jyrCZgysOE08qQUu+JIfgCeaVfoxtER
x8C/nHzQnNQyk3NGaQyeJACpjaD5LomnAYlutw18Xf9FEJdtOZeoRu21YQtK
EyPGz000VpvnYYk3c6DEr5K7MqfC4HlBzG9ciqkyFr/fbQ9XUCuZdwl3pYAo
Y6lY3++smUNRVY3ylHvdH53OF1yZKS7GQKCw+vWvRQ/wOMLjraWLbKeKrDZz
9wm76kqQaOgEWMaNZx/5+/mnXkRk3IBqwdEttUQ/20ePC8irUDKUHHS9YKrz
X1Cgap4O8zy6Ggfr8l8pBdNEQxspFiCBIdFH33ek2tjis8AnCsJmnxQhVgOZ
9qOs8ApuhuHK50eTLmiK4aiTasJGWtShU3C8QieI+h2S2G7HabjCDXMe3qno
tq/0a+ZmW566C2kuwntEH+6GiJ/D23UIfPmswgUc4bDSF0NavmtL1CzZHdZv
tCemrJerucWPF9cSGqAKDOYVdADbfHZHp8aGelCorhRfq16jHmxjCUJ6qnTX
vn13zHZQYChcRbl1ezhporRJc7YYuCKmcIKrfD9nIzSGURYS3yj4UOBAWq8U
BJE6L8wzpi2vO3smXGbFnDxTkqj5PmhU/tiG73MTQVfz6suiXBZTKlBr3FPr
M8qisOZqAG21OtOf4oCRs6Nf/rHrHRJIpcbenGO4JO/YLy87OJAu3mmbeo7o
VP1bbf4+1l5lMgCw61YDu0X29RcSQltkfXwWmhkZGwuf8gqNA7gW2wjocW+V
YzUpSJ0A+Xz4b/VUNpGG6YYzD04Pgfy3z4C6eOYt0pchrmEpFjMj0UW4tkEj
B7h1A7MzXwAqsFRMgJP68KW9uH9a6+1/M4tcgrv00L+3V5dVIDpPtqTjgNOK
KJ9qsHnNTqYkuOq57VNlzzGn19DSz8V+GlUVkxIqJOuLRYvSxW9a+eGJb9wL
5pRv+2+k8bKyLvUFAYCPmGBLxmzKnDhQ1nxEM+xao3cSQWoN+Z1p9DhAVqAR
v5fMSf/vq/yv5Rl80awgocXq20iQBMLs8rITGKTDcxYEc1iH1t4Ozhdxol9Z
w/4LLJN/7qbRzbZSX/ywQX/AgrrgaVfXvnM8cY60/YXXIZdoK1mU0yPEdeyN
sbADJe4TTN13FtkNkbc7jK6Hd/YsHwR+ACJvpUnlNp9DE04TZTdCo5/7OVlc
unsizJsZN/xLD99H5IblhdPqPr/+v8g/F4aQ1luzQmwVgwrSdiRZ92FLQu5I
IrBwqsU27Rtz+2P2mHR/8cO/v+HblnucLkc9AFo5boXO6cDJMv+6zczSDJTf
7nCVVHXpfntYq707gC9mTKE4I6npwhYnterjiLU63XnlJ8Y0ChhaF4c1yyVi
e1N9MrRX3LL6jtvNwceyA5G0O/R0ePe5osJXcqTX+0f0ShNuJ3zhVepufK6X
nFyYTYJ78aFAur2DoW2drvQKQigXgphghEF47vu6zQXPGtRk0cmA9vOcX+h4
OpH0l5oO7oFyTUuZI1DQUPjpEPDeeUFjT5nTGwIacDyGlpxmG/tQrNhGvmjI
4jfJ/pSPJ77PRouvRgCOml/TFEatrLXTICuCoZl4IGIpayDqRcgKTsQ1Y7J5
4amg4llD9Axj7n121W54pD2/nwAwQy2YoXM+u+UeATSYJgbMyKfZrK5WHU16
toDg2jM2A6TJvxDJ3x5gF62h+mQ1T2bw4JpOH991Fc/Oh24MsAJPy8PhauZr
F1+fAlDpx+WZR80Xzr1ve/Hed84TbwBObYpcFySYDyCKymrOo42ekFFkWKy0
M4qa48tRchEVX7fhvfQo4zZtpk6SDQiA7qyTToOAQJnyjW5XZoDpMri/o4K0
nfZI8NWF7gZ6IiEa+rIimL69/yZwT+bCMeEyP+MDYtUQJLo8F9qqya2yIezA
3VCuoq+QCkvb7OV7GyxiDriW3P7QbTP1SkO2+PphMifZs7nx162YNyxpmVv7
H2sm9gLcb+DuvsVEXs66J43rF+iMf5Iwd/Fm4mO/w5oEkIGh0LdwDO7D3OY4
I7/UMrDDZRhNXVPnB5Z0dwIh1fGXomv2OYDEPueRXQyZJk6kM38jI3OhMgNr
xTTdY16MeIIqZb8vx+I4iJxCL9hLs1VUhhCw82hNuS4ywS9Y8SjwzS9r4RUW
qmbQNbXgufLaEK32Bh4acd9Zpxki7CIbDfZWjpF790YLu/j/bCLSWSXL/sWS
p0mvnA5sTiIBd4MYYzH5NceGw+MXAXhvQiBAGBnQQiXQ5kowPqhs21XwTyul
3lOuQyLuaqnqZUJjUg7TlEMBLWemDFJY8TQVKI97Psl3o+bXCr+OEoViwVvR
ss7gfQZjy7cGw96tB4gbIPixvDBUn0E/XZq3DeF3OfQccOPo2wGjN16PTcje
F81Vu/ghE0cYWhoRCpmDxpckhGLHGIVOLrZrWKIpmXeXhsoqbykdGnwKsYW6
ZtsukbwmojTUCIeBvsaSPmSO0T+pWevG/bW1MVj2R+7uOk4Om8iJKTG+0oSc
O9UEJ1MS8Bl6XZbz9ovBhYdgWn1iBy8QGWkiAlxWrIRuDEbVVaBMI1HtPGvv
pYr84Qu58d2EEMqpfxXBemysq1rD/Ko7uGy5j5j98wO18kapCjs9syLPnsC/
syz8hPBpdYyAIqOUhwduAFFXcoIIVR3x2eNm0RsbmERdwzfMz/oFL9yKO358
NqDj50LGPNRVjADmCkQ8hN0hqFdu02ChVG4rdMrZXNVwUuPSeob3nVZ485Zz
8Dd3b5LVQ3vAUSqupgJn9WxpGuB/olyPEk8PgJak2WTXeywBomU2PLTfyyqu
C4Ysd8juEtqmzYCltSOLUTHWCPwsZUllqKjSr6ZiSr6ADcoLmPHY3Bc+JrCz
GKBYiTJQldFCKY6vCliWEUmKVYWikO0yvVN7tUfuxgmpmuQXvmwxmMegOt81
v2wLlJln0A8raj/XXPgtnSruvQeNZyIIKhLsOTU15qOYXCyPs8GQA2U0shC1
amHBpCPISWr10PShLx8+2f8fKpqIrK9Qq4nl4tEtOCUKAS4cSsLzSNK6f84j
jvNpXeJ0Aw0qxZvU50K4BVox7yGLtUrHSbhpkpR6ZvQnuxTrLzq5x6elFA3K
hdYRkNcnm7L73vK3w2/Pp/Hn2uMXxIHuzw/EBMXVPcE1ELrle4POrNHb0+cp
uhQ7krVxoxX+fb+dZmQagWB/09SSjPiAj9/Ou/eKtwTHxEG4rPzDVbi0ARmk
fTvNBLDXnT7UmAdl+BPPaQVID8GcUZduDMiSDie34HIFTFp5snVdCwIyXpAv
jyxjzjQ+NqdKyQdM+U4SW+9lRL2SjaQl9L3MYGneFGglZmn0SK1XEckQmEIF
NoQWRsZR7EfDou5PaM0TeZP+5WFTG86TIljh4sn8KKLIYgCQDn5BG7cvzgNJ
lgpilmgw2mFU+r1k0OeP3OISYdodgFX9/w4lvrB1LYkrmtDn8J0mMRtHvKkl
ODj1XvTLoWstkuoJaHOEM90q8k/dTJsrATiSKP2sxZXr8y9/RdH3yfRFcSo+
Hyj9/rUwHdBE7R6YSIE4mgZwC9lEpPrw9eNHbfSl70w2FIu/KWXyjxn8+mS/
/GC+y8fSMAniOYCnJJ7O4v0O7ANm3xxcXo4+NAEKnAUgxCjQ2x7vp8YGzP2K
fZQ5VujPwDH+7KGIvdC8+VJE0FVoaCJcDmFTMTYLVvywmR4E0HBz1kXprAf2
HdFM204iert3n4wtOm+OSGwr+Y2w2HMRjHQ4mzCGuCN2xSu1+ufuSFhiW1X6
nQGWrB/+O7EAyK1FQq0fl91lHun3E3HXA7a0bYA9qLUw3Kw9AcP0Aj3oXWo3
At/+jQUhV+7N7Lqt24VsV93bJVQa8HFj+4fPTvzR5SR5EbwppuJ+jbbuaB8W
npbkhyYwLfCmniWCV8TWR0X58vnYr4vIdAjSSD/YJl5dJ1vZSJ0oRgrDEaWc
LDFF/ny1F3fi5XJCm7KbnPsG/qUAim6McOYR6Z/5c3wTzEL5PxYzactocAw2
dHhjEGGs1dhYvfeDo//hZWZyVDHxr0oLuLMNasjIMqPZuzTTMErNDDeR11Rp
w0OqnvPmhzUSrNKNS1krmBVhr99WMKsly0nDlnbsaDuCm8t6W6QyLsxvMAur
dpp2FzNM1VxGfxvbLYXkwjiafc0RsuLIyr9Ys+51rg6fhSrQXdFcz9wxGs89
2azZHO25n0SMB4eu4yVbp++xLhlddTto+hLULOUH8YuIPUZBoIojWGuNjv4m
tW4uUsmTqsGuABzuQeAruRTHzuVjCWZ9vv3LsaP78y5khmPp9b71oxJTkGkj
VUJSnatKzahdl6qMLiQRfWx5m5W0eNE8drgP7FYseTbp/vIpWLKW66lijh7G
XSyYbUca1Ix6OhGvtU8uAVUC72kv0Ch+l7lngENkARzcVfMPg62D7vx2Kh33
OvlT5DoVyb4DPVt04sI+77AYYxxS4C5DItB+TqFgYe4nFlzWbRBfX1fZr84j
iNKuW/y9J6TyIcKh8XgScWZ1wmcPeh+3eMEj01NdEjYY4Amp9qNxzfarzp+J
Id3bnxYWiVI6C5WkmjEFzIRb0bseOJKc80UlUwa23vclVwvlxV32SL2hyej/
bLJ9P2/npBY2wbiGZkOiugwRyHwtxduOWSZNEilhw9SMHti6WRm431TeK3XR
AOhigfg2brirtDwW4DsCcXmmUA7ibjiBzam3Mr+9grPs8DypzHtAtUSi6LqB
zej7S3lf6X5h8Q0FixPWN8H94UogE0xBDKCn8HOZI07C0TFe2K1/9zYvh29r
/ohwsaYNKfvHqxUNGKo6malmqJ+538O0WY+/++Ym64LWNTHJv3EjHYbyxsx+
ulIE1Ylj3EfSPQ+/w3ZANKgBcjdwvyYkTMkSndE7WTIwYznpFHpe6tkSjPWl
w4HN4KoUmARcsuJf2LaxQLy0a7UjRSgyczUGeg5n0RlV2igRcDggMAqkIAip
Rv4cck+VG2VIfz1S2HhrTcWkw4pbY3DwZ1Lr2n1W3b4rx6GbmnPVlsTt4X6Q
heWTogkjv3lRTXxBGV6dzIzu2qLv0GaiefkTrJZ2h7dfKeI80v8yYjlBThxc
NyccmKHgwUrINdpyia5Eced3R1kQC5SpXxDWERipaU2/D4kdYJcSzNJ1/OfG
10ih5lgkGv7IeU6TLZHylXTbLxJ59NfKemnqCNPwIgVt4S97FW/3KH9bBzQw
tyrkgk+r7Z1ob8VdvVLm0H6/VB6cpXHjOuvTbzG76jqfhVohWBPg7VIM3yVR
R22OPjfyvp8KduSuBd63VlCiaZPhMTInnJO0q4kATfbz1GLW8JucQMTq8KKx
VHNI8rJ3BIR8W5RroJnkFYMvnvZKmJS8XYpjd7dljgp0uVz582y7LvGh85lm
C1yFOm4o6KbVgbEQ6ctA6Ou4acaZZAHKtusM8N0kwQ36LAaSz2HDPxDETcKC
fQtfGiURCQYBSXpavHQwf40+jaJ1VFypbr6391WXqKVd239aou7lFcXrcdHt
KVT2tXjJjy9E/cWCCzAKga/G1xm1L4jOp1tYfOis+PTFZgDLz5Fr87IpBQiW
Uy7gaa8oGPd7bRdsbJOFv1jqTcVtnKr/wvHeLg71XqfvCz29VWd2D2gQZZyt
R4oheT8DwwZk6xS9xo2IzJwCFo3twB5QUJUUTHjvOI07FOzfiSp+4/S50tmm
NnUDS1Jz3hgi7JnTzokKHlPUJaCFHOQ4UeAsoDvuIzF9mE6wbdfwa/IAoESW
fqxaWm1JUycnqRMT6A2Avjux0sDEZqVTHQOFcR2kpeehcZoWW/s4pTkluGcV
nTnbEAlDbeUYmVAbbEamyCMEl49gRlvUu2JEVm3ecpHMFM5oNNhMeg8yx3VY
iI5KfWq5TKeXA4iMuIffWl/zIAqyIvWqZQCK+xEcKK35gxgkcr4XuqY9BGUc
5Ws4AUneNaDNlgfNjS+wobr246DVpGoGx6RXTRNByaiWhQB/PwYXPbKDqMsr
plRt+XZgAZ1Fyp5Gt8kaYaIUyHsN7pCypHUiNQGi5KLOOWCB7nhuenX9rabY
fc+7laDeMrQFweZWAiqatst3qOPpGcOra+V97Rf2Fr4ZIcin2Z8/AgcNcguB
6lLoeBdD9W0iLYDAxaqq/EPCm1bL+QBFRGmNMVz3xIFp5dCtutv1u/M4qwMO
515nXIiMBX/IyAIDEZit8showLFNqSZehDeZ4syJHHm5v+P2bmM6H8blmuJh
ajiX6rJp7Sm1tX0NIEM/j+aipn7g3cihfoiULfDQQSybU/NRl1WJiJ8783OA
67Az9gjPTOaPU6vXW+KkTgaigPylsLNd5Acjnu1EmPYdFxEyixBQ6EUXXijv
nTQeQIODtLP/eVDIrOAeiQBllY0dWfUPSp76jwCAHKsatwcPSBSNqN/7zZ3P
XmJX1vv5UTsAxF5/1YculH6qJFe9Qf8T9z6yxvx1tqjfwm/W8OVcXyIlNTGJ
dAp6F4onZDsaTdiTAzOjvXmcNKNz3wImpyMtUdEY2Xh61hDOkEC11F7OEEXI
V889RVtcCCUniCKD4gPVO1g4mMWyy3vhjzyU7RMR/V53G0Pud0OAmMYfNDzu
c7mEgsQhEU2UjAfAEC19jFVpLQ9NTpTbUgMciRrWU3qD+YQFt9gftH4vIMJf
sbsu9JCgFxZzJf0qkOHkkCsWJ4ytJ3dW7i0zfOXsM1zg8flscztxS7S7pR8w
2BFa0gHJhRt51w/7d13PycYfvdne42k8aOfex288BTvziXGvqulRIDUfB8X5
bxBp11nYMAClrq49lsrzr7PF18zkxH06XyeN6Qs/CRhvGg75+U9PljZz0aMg
/WAXbS4Dz2FTNIHV/FLWo7OVZ0VJhKJyabeH2CXoBL+aNkxZr+liT3paiIf2
eeQaTW1/FXGW4Pr3hBkuVWRGx6cdCSHn+sFBMZm5b8RGOS1o+csMOzvSc/dW
+3IriW03Gg0w95PU1cazHJoe6xETUIeDPhJznAP8nLViZXzAE7z5yxyo0JOX
JwqB7nEHcVCQL/j0MIuLgy82YT6qnC5plskVW5sxhpSDVmP5RUk0hr7nzynB
F/bnERen494XwxR3nh6MS6/r43fu/ZA/DyZJLM8l4pGKLminyUjubNTPGdu9
juQDxWNVazYWPk2BIpHzz5TXPrl45qvhLhX3qRJYYXX0ovLcUjkQnEUH+2a3
PCi0rhsCF3V0kVPPUOLnNMJI9d4BjtHZ1qnACGbC6oEsWLWHzO8ho65LJA1h
dRd/d/FaSxutRS1m9KwbkqbPwZ0wIhNGrdrjrpF+f32HqwKuBMK++0neXxas
o15RgUm23gzj2bLQQUsM2K4UWynqRaa4TCSx2vUtW4lo7z54qmdp0tdfATLk
QEjuwDcL5PMmDJkNfMfQHZQvIDnkCR15dKEmjJLONk9fiuzCL5n7NcwC9gof
w7cjq1ZqK2xWdrXhCtDHXSvnagKwQO/xUx1LOF0axai71yRLuhhJZhaBW3p5
K8sJyPNuD6Xrygcwf3/2T7UIqPO8coF5VrdIxx2RNgFJm3mzQ/75L96be124
L+AI9aHoTsvGYvD9yXoJJ9pw09A6mVar/eynhi1p/GV3nDnd7UYtVfGCW4tv
5+b68CX3cmzpUvoDZ0+S2/vKRIYrvLJgRu3c6rRc9hTMWY4XUozAMwyrkMvJ
MIwLYc3VsO+FseCuC10QIPAaDeYBACdIyxs8on1HmXC6hMgLr3buoYN1Tif5
t9B06nr2xncCEeRuXSusM/ULjPJ8rN+8kQUENNmZ3DA+GC4sPnRNLsKNr8Cx
/7DxFenwRG73aVneK/y6f3RewEnDo5lxeYEhoCyQISsB7EJ35Qmpou9bKlZc
DRmweIRgCDJ9odgrNdt0YVgReOKS64sPpwxhW4PKwDRgcKIRS0Qbn/j3quOT
9vg5WNDYE6Ew+W3AeGit6M7ykHpKXuC+IWxiidZ/0PFlAxbt6ek2ncD0AoaJ
D2FFjVBcF0mDao5NohTDqKuluSSMJr3SVJGSKhtLnP21CMa3LzhAodxQLgY/
KoFtN1CU4F3aSA1Tb4iyn2TXJSExkDSxhWDJiD2Z/xShJZ5sBfdiYYf0fLGw
UZeESWK6HlmST4uZ78ZNYcB5Wugck6dBO3PeKl9zZCYRl9ncuZWOaXLnb1CZ
R6y/uwqvVyKgVn4gh2iskjyEkrgHW+VEwzN4fvqZgsRfJQA6JmdgF5gxQECv
XyMeCgyBTxmNv7oPCIWXYSHsAAB8tqhviwGa98XfLXaswbq1DfkL7DWCezoV
PKxyIpiMkwfugHv85vKT/Bj+tz5Auq0HQvp6K3XCVwX7nkqVZMYNQHk24Yqj
geeLmDBZm4lR2Ab2wXVIP2hscKrgMQZJmL0PAc+XmGVvkWYxzUzYU1lotYQM
OqZfJiWo6V6DDGOqHfddB/PnrQsatleq0dCEUIdUd3G9CVYyH240EN8/TDC3
8AMspQ6vhHe9a614ujLRPJKK+UF4dsdGwHno12bZT+pGREICTLs55GBkihp0
YXS83O0PAIBfif3smsQU0w5LNMqN7liqo4imhm4aErvv2psHTtVQy4+fNrDv
IseyPlZFu6a8yrciwMaRUmfbE6jhRYZeICOrPm6fjE0aGM+O/iBpnEKIH1Ac
ZpO62foCvERg8l8K53RRGak5ev1izo6VuqDYhHp5WuFil0GhpnRHI3spnxZA
YWwN2PoGGVykQSD0jZ4vHLjETtsnAmzqGRXUis44aamXh+MZWmUUyZPf33QU
RUKwwU/Ny1fuGx8v/47pOnlermhIYqqHE8kRQt8DRwcRrvbzzKV6pTv69hZ8
R6dVa2lNOe2SMkguqEmDtzuSs7pMURdDSAjuf8/+7DxqfBwGsXKcH7ofmHAx
Sou1Jx9YEdbHYpArNlvab9221funheo4ABKny4YlpElhO44K8DHU7Blen2Zw
2gsbbJNGhe2jAjlSsJqFcF5CSTMEnISKfyBt6BdEt45NhVtVsTlZLRzMOh/Y
dtsKVqw+N9TkGkTm1chZDu/oYORSu44kpbIJQf+o/XxO5pxKOyrmRJUiGYaK
Q9TzVOzEJimT6ryzs1ihMXwQDuEBk/qCZdAcozxbM8uBdDAhA6kQWu0TH2B0
dtKFtsRxpbasUsdZm6IRB/lJfAqKuymUhiS7Mh6wulddgIvUH5BSd0T/AoKG
ECWCr/Meo2sMux8sEXjlOAow5wWXEnNvPsbDZ+CPIWRsovoP5L4dJqH/DOva
0NKWPEeyYkn8XdcvcRQqdrSJEa88TZYSkpVLdRSc3QJ47KiY789gqMiodhbT
Ow6xA8N1q7GaC3Icp218/3j+SPRAAoiaodghOW8ry3tPGWEciE5KD2zRRCMR
gKurch5bD4bonsy2BQGRkdQIZOKTCjTtS/79U2YrVxZSv8g3xqR/WJmgPK39
yvrn7LlHqKHFI7TdKtCuUdNA//03Kdhe9X+NVsnkCUKIqJ/rIlFSAsZ75PlD
dSYybvAjBS787t4m3EGx/SpUy8RjyQ3jGrJ5kRvxgvmtGCdw18OgEw7P//wJ
7CSTUFkKpeS5/vChOMXn27zfp48ikSAAZOxrUgskr2SPYJOCYELAqzo9eph5
syrbC+tl/he63rSqJdMQdORE4PWIMneAYYjzHwOjZWuiY2XNYg/2BtMulT4S
ZrGOkV0UARN+Gndcs71nbPkSZyFh506xrfpHyrm1/XUjEwLmYAZ8U2GytBg7
gRCp84kbOGj8PDAXAncGNbzsaDrwdy7R67Q0hUSA1HARMSmgp+2jwRyCIO9z
aWOFS1VwgQn0YaKhV5fQ2xemxXJeJVvsomnrSznvOMYNgpRtRVdPZCpbndI5
10YeJOUbqqUG8beDVLoQl4WwXYUt88O9AxPfexabQU/EwG8q1NdJtPB7g1ZL
VNXMYqc/nhzL8If30AyKn82y5qWrvne/ZitkXQxcyePg798xG+m9KQBOOzA8
WONbbLMZeuZPikBsUMCBGyqdNrJ7NkulOMtIqZDegt7OsuqIVnKTsNiPb0Q2
P5OJTX0Eky8SeHnJfAg4fGThvrIpv6b4+BPXf93O5rb0/V4sO58WChwXLmK4
zRM4CvcqPbBrTaAh0iG3G61Cm/gUT6GRy3TbImrpRt2rrwpXjcANuqEfO35K
sJ7DVkrn/AjVoTFXeO/6747EhY688Yv/AmZ5HAl5T4QkbQ5vPwijW53/HNtb
KQmDvJeWGBU8SJ1FMM2S/5Jr4ZhE2TSaJcxFMPl/Ptv9+nKPyTvEN3InlxzV
MJzYSmAKL9xON4tBj/ChzQz6QbtYb6aPlQY9Y0H3vTvqXDAQguQIel5Za103
mm8HhlgCV0pCYmDgmYXuQj6acJEl1etL3htJNZjctTtlgch7MVaCzXw/gdWl
usqRIAI5u7qvstBzOHKYMKO+pPUw+cCKP7zyGjtTzmRs3L/kn1xp9h+vAiPS
dlE9aHv8T9AlK7rk2lnDvO6zQ3+VSMJPbKzrJHWIviCZSPvKqRRJ6VS8Th3v
fMMhqCwaNQ/rHHafRiAvQE8JetXCPSvcApEJYZaemLYU4EF6LzU/R4febfA7
3/cHZqVa+RoXGO0xF0k6gJU6nv/szEdwhKWyTB600g3Yd6P2oLX7WAuB5mhj
81ylcXsY7gs6QzY6eWgucwEIq5wP+m60kAVJ8JqSQR7zJ1ZTvtXe8pLPFuEK
8XCq8wTJexJdw7/uje0+8a4rKtQst/BTSiO7S38OCQ8q6R/ecaFDb9mKEG7r
TSh/xwANFXtfQgldLkJhAC9v10cJqxs15Z73hxyyvBVM5gcACI8fDl8hgEzb
OXzxIsia/7L7eAijRimCou/uZoJgqlYX8EdJcBbfLzlfXOHN0YU2CQ/EppyY
zf9V/3Syhi+cdY0tyHpnw3PBTZVCBSYnW+JpN3iMt8Ix3+OeQkVodkc2PXo8
/hnGbuAlObhDEvLEMd+IY2g8cTwYCIcJcw+0lE4sio8F+IpFIybhutzfe+Nn
Ofgb+i+0ZCgzAn2BvPBds5aAvJ2wpne3ECyR3GD+8gVFeMkNkCfiWeJ/qB6T
YjZqd7M/gLgy6emOx0iLAYkIDzWkOn9M2NdvLSWwqyPwM+kck2OtTIrGwjQF
ByQ1Z9xGChororkUKMPFABD6t2UAfknsl4c3ZRMmrneA2bIYb1cb28w7TbIy
R6yzJUuzMyFUbVRJyAXB6wKTs7+TbcCCdUUNAvbs83T5BTIxDzw0WK1cgvHs
8MgpjDgi8R0DLHCubF0irFY8MfDzWCgNtvE6+RDMdxQioKPG8QWyPje4A++v
vrcWug99WevV6D2Pw3HuJgM4NFJ+hPsiueh7ZUrdl9032/P6Z+dcYeT4p+7l
6WVmg5KDXmxJpBkn2fKpbtJ7a8cVaadfIs7qRyfoRINxEfUs9G+HnGJ4KlrK
AHPHppNy0n2s+gaZznNjItkXz573rnbW7aI5wVpVRBiEuJz8TEpacTrLDIRh
h6+KJIgPZdsAGtitu8zwZlmrdcKkhyK3iinvG5CtIxjCJO3Z0l/xr9SXaU5o
ECQ8Ejq4e8+HT66FeACQsF365Qva2dAUxunAV8WLEGnaJbZqjX2H1eaeyR79
8hte+3tLp3SXtJ7i4/V12OdZbiA946D7SMSqyHrJNz9uZM+B3q3qaJw8sc1L
dPwadzHco4gzPtl8pckKAATFKm83YBi+OGOyhrugY3SDeGNgGWCYwk+Hw5cv
bOOypZJ/gZnZQ2fcfbkQpfSzfgc5zQ5jCnNUoZ9kDqnGkKp27SCDv7CxmpiU
9aZt6ukbZUONJUC1p5wnImGFsIpQBrpqJ/BjqSgwG7EAYMPDvd1zywmt4jWd
ZVI8/SxdQOVXS2hVWKtqMhjlWel6zbay9dNIYMW9RWim60HM9Tb8bfdPmmfZ
HKelRlFfLKwSc2rTaYxkIz5Khal2UDzCpGPbi49MZ6MHOU7eRxtfa2NhUE5J
pYdhHjP+JI+5ZaUvPQASEfRXCN6DPh04l4pZfnWNE6zs0XuZ/Mt9oFxtjISp
YtuoNA5ZWzJNkOIg4m6FQs7WfXCsBrEmEn9cN45m0LPzZaU0FClPNyB1f4tY
qcY7A3CSoNe0+2wTUKF4QPxk9unYp3qn51KT4ehGUJUsZjtwPVTJ5KUwC13M
HmL8+1tUdPj6A2nROgIVA2K8rN6ScZ4BQQ7D0Xqtt1cG2OrHxWC6NI3/22Ld
+BnuO9cweBsKnNQkInrWcPor5oYThWD2w4/QSH9HXwmvs55D7uheUHuI9HWl
cpMqc2fZKoA4M6P3Yt+oRK5no44kBf2jS2G1IwrVYGYH3KmjDLEM7/z7FiMT
uJvOxHp1eopqim9CgEPpniGMT8gDPSc3Vac+oP4cR40yt9e5C2lAOKR6aEjn
JQ3+LUJwj6PMrSF11hmR5NJKnT2AIwtpU9CTDUOeyXIXHp6g3wjiPuSLOjVt
DajjlAid/VreSS5TEx7i12/q5ueTssA3w+RZ0X1v+PpAX9410cJ5L9rlyv7h
0TArzUm3+mHO75Mofr4YO6mRXBJncNV1xNO5qQXK8PeSvGqyEl12/l6XOwCU
mPLJ2YCKhllboRVQvI/23HVSHw2yn2/PmMyRpO4ldma2sXn5oYLMAKmvfi3O
4+E74goGGHXICRb/Jb329I5N3XwObGJyttNh3PtZ2nqOR/QF8d3MmNhbTUM+
3QzNfzckbB+3kTy+HZpnF914ihMlapJBOMRK8l2SIKxjx0Q7OwY+jF3HD/9D
jYwRgLz/gtPBlOmbS1/VEpDQdP5hSWgrakcldaNie+pnaShQs6zu6mAnyXGU
KRqAgKq6BBc5I1r+Ak3dtyG/BrNyHs79vva1z/6Dm8XeL75sbIuHMfHk+Ets
EEUM2kXU8SmbapQSKKUlLKPxQjR18qdqmxC4G0wOiyD6pWs/2dJD/6PV0Xn8
d2Vl3AdihxgcXwd0Ej3x+xglgLukuLHBbJOAX8PWXl9wF7Un2jNU93FfbVIS
d/FtlcUZeYGyMU4Dgsz06sAM52wXeHyyStLxyMGUau5vHklRo1cHYo0Drq65
ZKgXoR/rTatkw8kUulZBz5KDiVWLhL80J9goZranc3UHktNlCvFmqScfe3Gs
sJ8saFQPGP7LvVOq7p7EJ8AVZut3iKZ6g9NyjjixvvQRklm5AgwqtjEtD1mI
6Me11xhIWxfjcZ+c0h3qI0sRVce76DTHVQAQa9NYKRqKw62rAzsnkr//Vs0o
hR8W9Hqw1Mt3t+HzOSbBKF0sTkEeDEKzs8OowOvSEE7LGsYXtXRcmguygPuy
zZCRXIszcsVjKp2B37xQYNv5yzcnZvHa4lLR1uNRxnZFjNVzmE7pqPUMutCI
Gp7dD8z3Tzu/plUYbLQwqqVpjhLdu3LX5YQ08UVYrUrpBwNxKoaf4+sDQNDN
zvpqHD3puOu7ZkEWWdS/zkYgvJkxPNi/vvbAKAb5bDi4nlaSV21IF2iDxxTe
hkpMBR64X0gDVI+Pp/anqs1GLcRNBQxgIf9vXfQNYtQC6um7NuzymGyFJVic
FfIgg51V6NAV0Yd/9OQaxVXhUVpU3KqIwgNnwJe19LNkIxO0uZk+3sQN3yyJ
eKKpp+UfdlVL96dNphZtldwKvjtFNtojfkGbsqlZZtKT0OVhxdaFkvTVfM+O
dhL6QJ+wmU2gcx1iRJ6pd1Ie5BiNzmDZ1rD3d9EN4uuXbg3vbE6e2st4WqM9
6MORUM6ViqtfGL5HbcQd4+SqT2NPga2C3AARGP4PBhYCLUdWgzBBSc8huZl0
+wrT5fMd+igRuSQo0nsEGcyVmkqFS4+A7rZ7lwNLXSrRUNN+lwVabpiksjmS
0GL32j3Oa+JcJMJaY7GAk2I7Ve8VFW5/bVvtrYNxwMl5sWIPLqTWHsF8vOkw
izN6RyaNGwC4A+X7LPuVi1IW4DMP2Vq5/nBOC8qwfnBzR/rVTUbuLgi9w/+f
6LV7/6pb+Pe2iZ0XsEgXWNtqHINarjyrM2O5YvEUtgotp0Y4Gr5ZPc1FnGVA
1tvnLwZWQvUs9+9GreCARq8BZ8vwgvMRtkVT6olM3t9gskox/jbrXlBH7wT6
eLoj90F71mbN24x6LbFvYeJXqFqFxgcbJx/xWEWCqfUtad0Gc2gOSLeCg6SR
b4QO47dmMBKFZOpq41LKvW8c/BSg/n58dHAA+XMYer7ngGFQ9u8udpy59tEi
BNbUjRL4YQ96/ZJWN04LwCzOX0AlEOOMWz8ukIgd0qR5PQlHc9mY6FWhF1sl
KdLLmpxbXN7huWg3+p1wRPkeKtl+G3XRlz21aZSWvkLrplwbPzmnA15odx/3
4n8xdj+Fl8jM7vbnBx9mCG58x5MKVdtzX8DOBICITmw6qdTW+vhvMkgFp2+f
kPfDuWvqeg97Qm3sE3aUdo/NWDOvDz4/0WpUjFRi70MJoV98AcwHBzm2TlkT
BpeRTCSurptm5Zaj6wxSPjAfz4ztOhAWJiSzhgKHunrbkf2mXNddtf9AWU3E
smEd/ps8XQ4FpJGQXazXknsKI3KKP2eCTeVc/o1bUjDuiL8Yrfpf30NUC7wt
gTjDpkiK2NJnXwpp9XTYfvSfDaNkNI1lj3Oy5LdX4WT2tT5eg8pvRVjFqn9z
a1GmYW7KiNPv36S4T4yUngXFOW9EZDqH/WstdvskHI2ZgCCOgegWrxOecFJ/
kbD5fDBbqJmTo/JRqEZmL45pFCOQcBNWKKC/7YMjhyyL2NRb7IBJh7rSoXLr
zSpNajgcRLTQD7M32+L9JYrEIWPTEAECbagqwbTj34orVJ5B20PNJUCJyjYd
kUscMeDnROLlfFfhyMGFLRmSNQ3ZcbVrS5TVMN0xDh12WOlXGDdTVHtcR4e1
gvOj/gbpnJwU/ybeEilxmoKpcTYAEIp4WxzmcZcOm0wpIQKQueAs+VaP8EbA
Z07gisRc1KKNMR+EvZGaNh1Vp/At/xLc3fIWAUyGFnKZBv8qdfpnWVskZMTv
Fgqzg0sN7LgYQyJZewzBwhbe/JrjLU/U3KYS0TOv16v+1Dyjy9vPrv6W2W5F
J1s0lehKKl0/DopAOPuwvc74dPnRNVeqYJ7UjvS0aEfxSJnv+ByXRurWUCi6
4nt4GQHJvCNQIB+8y5Q0AUXoduzkr+nCsnvKDr+SOX54HR+sx371RGnM03aP
iDW5+ZC07Ejywy6emewhLlNuBJ0IQa1JuLGITwHS0iOqq5mnFvYvOi7j4+ug
lMznU53T5OuC2qgiYs3PKteEG2XVNBrB/iT4uqQL33nLgclEKHwfurWScCNr
UiKQM41vOg8Sv7ykmN0kN7oKj50MykKr+Idgdy3OMqCSeQn9U0HzhG0GfNyZ
jW69Wi+4M9njeRuqmPQ8CdudUaFZuYMTBD7jGBrzyS8920xOAhKYNtm35H59
vhNv/WxrpEKVHdU691lwW6AkbPkGtf+qShJS/IBCqMEjgba4sWs/eWZh3I9R
yVCIlVYbsd3qRsG4ten+fExZA8BJ2GORV/RLAAzko1f+LSYqHZeeYgaeg0IG
qn+A9ZDe03Kxu6ops52kKGuhTqH/N2ItzQqFUMlXjrK86LKl/Sb36JNBxcak
nc33aHvn6PAkYHQIYagtEAnDZb0VnbuRef+92AgqbT/bLTeSPV+zOOIPVjfm
873ADY11TIJfcuyDxLxXdgEhMnzh23t27LsUa829g+j1yN2wQO41khhRvpZN
aX7tMT1rwPnOYeYK9AAXBzXvEqCuSb11oA/J3Z1W/uieYbxZ/xkWnXRQHAGB
MD5um6J28poRltIKgRtSCWzmHRoLqe8RHpBwzVxszkY3JMskvkLPNdytdFS/
SjEE/5bzkiV475dm1u6t1sT5O+/QZtXpeqF378o4+Zf2pfZtTfP198PKCUbI
O/sTdJtaUY2REu2frOSKxBEMUQxy+DKHwpipfdW+VR88T6kQ+7CsxS6txWyF
JD5zyDv9GBumFgPJPuhMHhtYKRclYXnf+JoiPdZLQvB/TFgh/AeKPFo3dIic
teYQf2aTvH+DM0B8/+jHVP0/j8rZWfyVX0U5gPh7EHZYjJ0NkGQ+lSK+YkzF
lUmFAePkSuNFxmv527Xzgbr3k8q5oywW2LKA1J1IebhF+JQNiJKXcJeG/LMI
2ty8/wKvYpVmQbLKHvTmI3nFSror94+MVjR7R3DPrcWW2uE3kn38HDk3/aUj
LRUe2BqQrKDbE7GHaZrWwAbzKSu+tyPjGUnrg9ojF0rWVq4ar8U6CDjJI1AE
wQFbeC9/ar5mgGrs3aPqicbKYyeqzVHp15bptyLin+0NSC6MPdr/J7wokxqS
4FHIap7WdqxgfsVPPeT0XpU5OoMflW3CMkbkMFcG8rWR1y8GzRu2SAodVzg8
1s2gNBzQmK8fwx+5Vl65RutdIITBgNzR4MxrFqaB5kyPClgrdP2JLsRyvXUD
B6FbUHWKz3wa5Yf6gFnhWFk5ysIknL/vTQmPxeBT3ftoUaBIva/qOwPVk3qj
a99IApmoW3oMeUG30OQmBrY54g4yrf+k9W2brXf9bRZswM9JZ70J2d7xNMs0
MLT2XC1CiehV/rX7XEeggvkmdd9QiZum1CZ4CFGO6xasnKjAK1sDSJV6mP3b
A25SZdqV2d/ypn/C6onbC7g923XhFyhClanDxEyAb4Aw3RAHBM2prkiQWv/Z
PcHaBg8TIt3W4JPgXW1V3fbSJ39Q4rbUFm9lsT7f8nLYRaFrkjYaN3vdOdoT
1+5PMQ58W4Utqrjt5ERhbGHBiqcY4c7EgN3GKP6GzDitVcI2Cs2lrYnd/Lg3
c4Lr6n9cX262GeGYodZQXQ3PbIfsLuyH3ac5zbvz8CKaYvptpHNGuvXwMry5
V1IbdCA8WgsuLO7m2Xhlgu0IQGSuqM5txsQEjuibYoy+QMb4gK0LxVkNmPtZ
dPHfTk+S+cS6+LtNh3whaDVTOX6PGPSP7QGjE6g3BU0+AbsgzAGizZiovIPr
cadQYlqIhUAYUB9Z6mNoQajcLXxsZy8DIXdV22Wg5n+xQq9fqviQRBBfcJTx
zp1iuQ4sgBdPeKAvTGWA5TIk7jHuB1MaGWjX4yPrACJKzg3q0DN16x4iWVdO
cWgkvVvA/f0cISDF/CZ+vnvFuiP9cHCxGlDMn4E3z5f6kWoNuHhy5WoWS9W2
yN82vU2xyNGYzduEI7SRbv5aMM2zqB/Q/FkIntOwpB9VAGeJbttNTH8GSDJj
pTsYd084JBaX9ESsaAGTW8zbPi7B+gihpiDbXrFHiUzoB2CXYRiiX6PnsgM/
SaXjguM7tL+6wupkwRQ5vklPwQ2BOYJJNJcJaZZFfAZmrW3/5YgXWJDOfTIg
o/JZzypeFa5dqRufMkVhQhywdx6YiY5rOINsD483IhgkEaDomQuFMKVlFILE
WrlJHVeEtfpyB/5r6Wk7cZfEz2oj/Huiy1jA0AiCIn5/y+CTMu3fuK3ZIF5c
CalQTrplIWmscxDDe2zrOLraS1USOZtI3w8krfh1g0QyU8e8YMoIJGCq0PB6
Ap3CQ2cZ4waGT3JmgrWkvUhuvZ27ubO0efFQzEHLEWi6WE5wV7/Okxrm8g8H
N5D9KbGEWkSyxnYamaFv2R9K/Qbz4Sa8vW4rbTg4Orr1monY51cW4G1+UFnl
UGCsVJz4WEsdB0VNUDxspC3NUHYlGXiPS83fXXQzu/wkqcYUHBdW8PbnlLFu
lwTpSqh9lSzcCI671wI+JsL83I82WQ+yyHGsGEd/Cw8stovXV4UyASaMEYy5
lSiSQ1JJ+zXs2oAedsdGRAW741ZZey91x1DJJiRzgu2XK7Z7I4EzwqxwQWWh
5dy0NAV+55eQECQoCoLThn96v7LmP7mm0YIoE2pIDeaaiQdr0QZvnD7aq818
WCWvThL6Qhy7tL4tx0+nGJiEq2P55ggEBzchLdRi/W1sZKY2pQAt6fg9Af4R
Xno1pNY76chhK2AyfNZRxCs4AzK0u8B5mnXD+88sOWFQRwUMYXskxgUnAW/v
SvN/OS3165bgRVvBH25O4DZWhjZlKyFWlUDI9Pzhn3n+PwwHaiZXHW8LGLbz
kgY80EygiFQOn7ZiQjLGbLW+PFW/dSxDTLymi2Gx8yHtcy9j7m16GJEHMv5C
wysTDYO2LnEBoJ8ZuN2T7xxqY1CjgehMmAotciw+FRFGarsKxDJ9XZ+zU+5X
bkP/YAFrycH6HvfkjXPC9XhLhh8wm7shBliojOk9TJaFlG0EEgQSJGmiLQy4
FsecHoDC2S3AvIB/QzeIhKl+IFEDmFBTK54hW8xevSPQ3rmGno0Zq/aCUeNw
U5B5hyD969vBle8Sj2Pk7ASmHTdp5rhpKZqOre5+7zntSZJT3fnBy2VDBHGb
a5bAP88NmnpP/EQ1M4GbTtNc3KosDZvQHzyITqzV0enSlMIU/6fRa5kPAKfA
NXaEuV9liVkgDiThfVDBSC4/kvRIxsknp5/9eT+YUQhCXrIwthPDE6PU5VQZ
fI3ZZynfMPNuneQlEIRpqVe3Lqd8pfU0hbIPK8zAMA4pwfTYRRbCKE0noLOH
jEpTxIuSC3wf9E6Qx6m+jWdUt3TiEIeYsu1I43X0QusbzZi80ABCgryMC5Zl
gKIL3SgJzTjpv5rZmZEeDchW0M2KwFQ/Fc87oE0lD7WWtn2TrwRezHsiy4o7
iGdSzz2WpuVyHTIM0cquB3vYc9e8fCdvsGHff1VBfBGZ71SZVHcm9fJN7quq
jUjqgYnoy03xEsT38V44GLK9bEmAiP87u0PjR9FbBAO1wcHsx4LxvDGcL3Eg
jMGIHAgjT+zj4uyjs+FNt2B4eLOQ6ah/WNHyHTjMh16c77jTPolObTpkPmRV
lowvfgjGq6TZmupi65WNF2bEyhVc4p5ZnkI899dNE+wtVd0pxLUArXmpJbWY
qwYAd3ZUn7oGkA+BToTNn4hIfV9Qtg3c86ffB7Sm3LZk1CLaPkL4jTKNbs8G
KiI4F1R/b5bSPdnp8Bkiruo/261VdDs8zwb3Q0VBHe4tVzd5ItVa2sI0RMOl
oYBXbdaeLW2ah4r9IcsAY4OKwmcwJuvyolEAgenkhg/FCR70JdvAIwC3HF9+
wbdvLmWbDCliEbEwNKTJS2p0oljD1zuTqgzJLM31KhZfSkvVSo2yguQuipnk
uOAIf9sZORjrpTRXTM75+/zO5gqha4MVVsQu/Ewpld9twYoWptSLsr6JFFYs
PVrYq5zS4ZOHvH1XRwKBRM4NA6ZlkDWAn52l/98es4E2YHLOVBSuAfNz4HO6
UNIhaToJzkM+DofhEDgAggTYNyb1Mw3RyOqIdyxMQidzcJp0fw7TEXRXBxes
ax/L8UfgYwk6SQSuhrX7wXRBDnZSjYL4S2vxNip/g7gQlpH+i3QtgpzwVYTD
kP2dziC68R+YRTnbLGEzpgUqZOxefj/LobcfW+Twp+9syox4u9l8aZZ6iFao
drC/Hl4trKQEvPLHqzEe8Dhw9FUm3WtN9JZixMXdxGmggl9VrfmPmlYuqQ1k
AeARUii/q+T3KuwJ8wItAPxwmSgAjuccCO8W2THX4SB595X6v436WQhliv1v
GLMx3blJrfTx9IDMTaHkGeAgNpHHiWmFdLeGVxr2Faa7IYWTBxkQjA4qgR+0
E0odLho1kIM66ZYFoDZHNj3ef1i2yDdVHQhdHYAH4NCMrXFe1Mf7eZFW8WZd
eQO/Fbt+jfIKfJe4LJec56nm+paAV+wrqOTtgJASx2A5qBGy6daYP1WquWmi
oUPQVcZLOv6SN/hYIbrRT8Cj1eXDGg5ucPFNFNnKg4GQ2PhE2ZPAbDXw0Nrk
ChD2cQfSAUiU5nCpvnPh957Z0cKBZcMf1Aj+kLOsyth3G9P6clFEdudoP5jt
vkqrzpnKqpf7v32HzR/7pODu9FX8/PEviTfPB2/9iOZP2kEdeiW+x3lev0Fu
jegQj9hweIdFY+Z8JZAtgOholNmHS8sX1g99cHvZVf9pDNKrm19Y1nolDJEK
oG5xCZxqaqPs0LWGq5O8gDr8RDf0t4JudGPiQ6/2pnZJzAZOgg3f3wCwsjTP
71/sGnbeBlD8duBqCJRp6IdabAhkuVZBLYonFkr60RBXhYjZjeAD4KDTxLLE
8CoIa6mL2YCl3zslUkImwx/g0NhTzPpphDE0K4vKr04XVYYhFp3+/hxaapFi
HjpbdcQkxpwXup6zrjv6L1Rzf0IoC8hdcWUqf7y+hH9sv3ZdbS8oQIQXRm7a
KEtPUMUVM18lEmKAts0HP32IPtelD8lzbQ2ptuHqYMZoZOiqXQxTFG02NXkC
a48s1YPczpyprG21imtg47uJRGxLqn365qVskyhzeqyYCZAJaRgt87kEQ+K7
9H2yzT2oGg4Ax/w5ER1eqPBjEDiHgZh76+bYLq2bbUWIp4sdc1zQUEfqtI7r
W1WvFTnsVLOvEy0LpkZwNDcqGxHzuUwUMw1uwtsevIvvIJy9JJptsXrDiVbe
CyQWznsvgbalYytd6VjCP3tshZdouTBX8ZCSXLH3X9dMx53a9MveV/xcw6rG
ynSc6OcWvtNBt6zBacbIe5bKIPcb4TDlRsHXiQdfMecITFRHDSKPjKGIx+vd
HO/AvW76sVMJswYoL0FdL1KhRpi/FbEeDChcIFSoG6OcV/tuyS9W/emNuLsy
8R9C3V/NpQMjtHQLVNKlq4LZUP/6B+WuoVhcznBrhUz7oe9ZPnPh9ED1rEiq
nvqkIueoSL5Clcjjovk7F4HB6ZmK7Sk9mQCAtFOrD8n44Sat8G0rNvH6z9PI
Qn6O/Ip9aneYPHk0fsLcwVSugbVeOAE4TIXIEZPd0wTNEnd6ueFlbykZ00Ey
+iYfTyi73X4VLrOV3/9+2lneWrHefVit99doYcrvJDiqpi0f1BTGtUIIoosv
3mY0JeDp8e+j7/DQ4nq4hy/XzTa/+6qpMVwtdT7fjAW3voLBVf9NuJrbxhVO
2aYTwlkYy3tDZledfKUeV+vhd0Yn2aTVsLqR9lurtVdxBhfjxlXs+jGTgd1B
ITkC2RZOdH+gCP9aFg380LyTlH7YEMF4hHow7ZA0+Tlkgm8ZppgSJNYlw68S
kqu/DwHppFdodvSngIUfj6mtpT8DN3lqkBxYRcL/lwDO+qtpYnH3wGKL6elX
GpZn5lhImn+s1omMu4TH2YRdBmJFuN3V3wDkVQrR8L27lRSk3M+RVPa1LrIF
6Xo/00NgLwG8ChQcUCIvqNJMjuoQOtaKc9IIeYTGVzELbNpDs0lYFVuWZUg5
E7HxWUeEncqZ71/7olopmJ/oxdUmflQQH3tsF059TgAEINp9rF08YIfPcPwO
T4WerXTsEsy1Z/NWMbsqQHvRoy8NK9GNZObCATzvkL/QbadDppaE7PRUFZvG
4eludlJdo5xZggjMw0sAuuKVVk1hOe42ZrPb+wfOyaqmf0QkH9dRiVjYzTng
iiR3JPqjvfP24Ga/UI/8MMHRG5paMjv1UxzRVkj+h246eqtgMH+4UeFZ4jhX
Ps6bfHRlaAvDRubq5oayWtBNKn6xsyUV/YbUf5we18enHTxyVuPMGQcWBDQP
RpD/OQ4rQ83glXkwwhUYJzVlPYHNWhEXUhQgvS9l0eE8xHkDABSp4i2pyL9r
NwhhjZl0o5PFE3OdA3qioqBRYL1ymzV0tHYjuNZAJz/DTxIbidA2blSp+qW1
iL+PqeYrPskSy1OsSTNxwsEy0/7Ps0FS95qGL6UCrMrMC+g9FhHS56igjoKp
kLlwoWSD2oSLGc6rg+8+Ppq2rVcbxap9oRiaqQKg6Sco64H/hYkZS/m14ELQ
3UyMDv1/QfBgwVquULrLePVoYh93ePyUvO+9jQrMdIRy6lQq2FjJe02y8szR
1Z0L9R9Xt0RGbH9A8Yt28fJvFy3kCgx/Cq72exVGilG/QhGWdDpmmqBkH7er
M3mlVXkPk0NQD6KXtUEMFApM0QO9EDK46rHs2nqS88rt28ULc1R/U79/cZwK
3b5BO8Gq+QfyMj3V1KBFrMQAJ69ePPXbPrSu6ja7JjdRTfmBhw+WQuuFNOVE
0I4nMl/mUuOp4PETABMGGCHLMUgIcRZhyd1jzshNLQy1QmlTgCBMxZIKo17W
KIxBMhYSa0TwQH5OtGmTnluu3JEua3uj5MF9YyMV3zLOQSrJNHIjk70FXbyz
9BWkv17nBH5YyE3cvfsEB5U6QAAJr5DjpNBpSnHWNSKU3Ds2SCJvQrSWRMiO
jcF6tDz9kjDHUC743M2GsQKlXX6YQx2ThMBbYUcgyTipyaTFpbzPYy+8JddO
YPlSS6TpFfZ7OAdGFWzNzEffGqayLxZRuOLu/tdiaAbU2nLESgd5tXE/FtaJ
8zxB1fkdCRSDSWBBJWciTAbGSmH/hmW4Bg7hM3C96ufpvu0PdyV9OvkoHKdA
FZNBlQfKQeOSfsA81KOHmgSDTckTltSQPHSgzAINWBmTgMCwNJXqcwAEaq+Y
hZeFsyLwFQ1zOFPYrqPqmADcd5vOPyU7PuOlECh/jX3GvaVdKDyuLFND1yVe
8taW/zbdEhTrn7sfFWqdpEgnKBF9lq7JeXwNCYc8mTqQVtTjPoIL9RlFnVF1
7KcS4LCWfyIPiBqS9q+Pa53rY2MPwzpm/YWHugkzxALfKgfhrRXXSUOqGl+w
69eEWU2XhN0Wxx9W4APXviYtm3Ooya28QAKiE1zgsF+hr17njzzRd9ecoLJD
fyzQtgliI2k1rt5YWFZ7Y1rTqYnGAEW4lt60K3kUkveJ7qKdNAZCC98d/gy2
W0T6nQNBtf5FGNuTZbDEYZvLvtOcl0Q+jLc2ksy0m+Cl6cJ2rGLXw1mWPgGE
C3apI0g5bNaNAdlzApsyNN6/HDCyqqVzk/N+Cq7TlMqAFig6iomo3gxLvWpA
yC5ohz+dTnaCiMxRdutLlMy8eu/zQ9fsAJgCKeLENGgsdPDPizwck2KLqika
budzU8HJmWK23UOLhUzqd46fiGOww9KaC8QTPBp986PwVR3TsRZUVaHr4kQw
8Z8Aw3AExDNUWa+5L9bTFfaRd95Ve7NDd4VO5gKQyvxm/O7XjDfrTgS3vp9i
HJrGJEsGfRlwDz29ZRB+xLM6nYVGAQGoXjj+lprlDBPeb5tP5MFm4Obwi12A
PRvN2pT7+6PMxipWF1Va+/EnVVVSl4wK5vOoHjMMJNgUALFT8dVaNilr8aWk
MYySyuvc68ejR7eV6zYNHz6MCMgqH6UmwGtAuo+8fO/O1Ve4tk4HlpwqkhWd
Bal/TToSCxAHVhICv2qApIMQ9xK9Bol6uhj4gi8NtoF6xbk8579ryyO9/GPR
f0T50+lUD5t0t9t93ywuTfSWQ2f9Hp9mRPf6Pstyg2jbRV43cZRKRm5Xfjk3
7CxJHehy78T+/lAGpKMkAVWbMKXNcWnVW15UXTivR8+A6G/FfnRCxkItY9Op
r5RmB3hkZxAFDR4v4jwLEz2budsAvGxH7ubkxUSZCPUKzEUP2sZvb0EQ4Gb4
0y4UZOwDRG1rv70bTEoWNURxxYaIoUIEpsLG1W5tW1ndpNDdAwbScyzZTinj
joYazV+HI46d+wfXkX8fDvvpzlhghpMcOjHKJ0DMm/dechY/1UgzAJdK1Cu8
3Z3M+vrnERwKG3L7UOTUXrrJF/2UMG0i5e0Yk7q6OEC7d0JXrjmqFhMtQG86
ENt0cyNjfQPjxyK1ZlpBpd1tlLhDOYF/CkkQd7m/N47ZEKCyAkHjbaKBe30j
BgcQ8925cCEmA5GPmcU/JhCeBpt4M95qYvBL5aegn43VWSB8aX2Yz8z/UCmO
Z76GINhzUHsH12EL9sQHNRG4eNaJHtFj7Gmm9o28a1Yo39dMgjBSk1v6qoNP
fPqgec1dGj89wrwlvnLe9dY2C/gX4C5zIZEl8d55R8fkxL9w9H5EyFji9T4Z
aojR7n2jcGC/AVoANjzF6fPeRw5jhzP8bPU+xCt3oxghwrLsptNQ85m125YL
5RQDZSMAN6IkuYkfkaCUcvEuxP+BiMTgoMKi/fBSoDOsdjPhozhJc0lS+e0q
NAShZLILfC69xsvR1045ldwvz0JdkGVQbsJnyMg2GwCqaeSnpfFneqDWt/x8
E6xN1qLeZYxteiOVXteWFt2NQRRnYFSq1M4zhbr4q1CJMNkhaBXfCmvwxl13
OTomr+J69g+W1JMlhjOAoBKQhtUoVYLFCPRwiG2JlqOm5DCJAGI6Aboikj6H
V1UA3enQOft0z3sZojp+X+nAKhx5s8OWSGHc3ZROPws3wmNgL/XIGJ9wlZvF
fJUUrLWIFcYAiS8hJo+TGjY5z9OSW3M2azaUTukZV4FG1ykW1KjDnZf0ctHk
ymzt9hB2TGL1Ufjy3i1HzilkMCUzEkX04U73SY4ArB4+CZObGqdCw+K7GrIk
AXJqVXF2wufgS6xQy9UXRi9eZ81WnE7TSlE/e+dtZztMYtjKfjKtyuGLTEM7
cmaLa55ZX9OeUpd7SXVZKNKGadiYHXJnwEoUH5n7bzKN+uJT1PGiRYJdNtgu
LQt21i+vCHFlnhX1cZ1KIaNxKO3Ip9LsI+ocVWOY2mI6Ac++SPJlrI2nnFil
4BHYEJxxMpMiilVqP+02ubR+ati68uljjmtK6Urg54Mq2Ze25Gn16EzkRdDb
MQzJI+ma5n3gsB2ySgBSvRfBJqCcO7b6sdFsk5zyPuW2JkCJ/fja7A8zlqMC
e07JlMkLBJP7UtZ6VPaIcAHzEa166dExt/IeHU7xT9CZn++wo+6HxyIV9cxh
grkBjO72/Bu69C0h8lERYjewz2kKnFYbtdq5OiXF0l/86BrBRJZGSYyC3Ql3
SB4Su60ow5NFqrFMnbigKNbNwSqLu6WbgfA5WSnHTuKvnHOYPunzLYuazhMa
GIp0VIV+LBSefdfjXHYJjzl3/lU+uUn+YUVpQC5kT/LvFvGupgi5G7f6XnKN
SgXOB8Cry10k8EOcsqhXUMbaHZVGBSE+y95x78I66sbLVTpiLAajqHHw14p9
XmQu+2KRSvOF6liDerL6AG+BuF+6+1jIxksJZLd+awVDzX9qDRac5gPPlGT9
dOTA7tVF7wYge+15xlK+7g9Fb0QLKd3iRPP4wVd0HobIUUs4+laJxss5qCZV
2GTL1ly+YIRAZCoJbOEpLb8bJjagJ5ZHJ8jrmZQAKlENTlAfxUzNISfwDFYY
KXoKXNtPnUjxsqWYr5rpAjJMkA2EFnzZM5o+zEwE9XGRREOQlRzdPGkuJoDl
jjBE+KDM1/Ed0+Takqg/NovbfNWzQcTHfNaTz8q4oiobnN4GX77TOZNLzGSV
YNVYg12AYYQ6VURQIJFtu7cxQPKOmogMf3BVNeG88Fqab9rqaGgOUu2rchWz
YLQoQb/OltyZ8BREDLlQPseLgii4yUwH70vdyEdUpWK8SNUueFID2ayYngoU
h1fvECp+Do3Kse7isPjXqfiCNAZe1xQIql1R3t8glvb7ESpy96NOvre8SRtG
rC0d8d/HQHDdfBwjjl19D/ox6MhsdTYK6B82FOqcXnoh8CC6t8o/aGc9p9ml
z1ufn0m7U0ZG8VN5nh2PNcv5wNwBCiAtPXXDEuqFDSzO9oGyA/h5toCHTDhL
HGytmwWItIXPiYE8AcfinFvMcmyWaHitHPUMwqUPgZCYFNi4pJ/wlzYQ2E1G
d0ul7GPbS/UG7GcYOF0dYq8KW57C50P4ERT8l2n6heTDhreXYWIpATCnnRmL
SSNxArH8FKSEkHn3ASBCghClVfeaen/FK2nOO0oB/sMZ76f4ZOHNIrCP2ETe
a9zXZtfIkcngpeXHyT5Q3KiDD/2s2lIvCItGflQje1eNvOryKm6t6t8e/HXy
9tnOPgeiae5lBSz04/LRtUg0//SGIrMEWrjXJkvd32tLObc0Qbg2xIbezD+7
RfJENCzkCiWonRYaODiIsV+yg7LIsgY0WQ9j21GSKUXlr5OvHaTaxrIbDBDO
NCxt+uJSJVHK+Ns4rUGPdw1pxLN3R+tfObOyD3nFpkoUfuKg929eK4huuMiC
jlwNb8MSoq1fIjonkst4agJj0Bx7xCpxOCKJHPytvaePsTDMbulRxMubb4zq
a50Qw49KqCG0VNjmXE7dkCZghg1OoxzRyArS2v5oc+opE7CdKUGNcTDqWTSq
Kgs9d7r2Xf8YLQlkc6nQwoLuFE5zwSbSZ/nMfkoFRfx2E6/e/gcarNHBOrDL
JhRC52wi45/ou+9hnvm9+KtrZhu60aQ/XlYDRNpJvbToFCpOpHpjqsNLAeSz
2Z29Xduddrti7f37EUPS94fsCh9wOkXtESeZwhw/iS5OD6/u/Qd35K+R7/Tn
ULgVY2jQg4s9V4mGsh8F6ugogpJr8ZSwPI+b8uwOu+3EZuS6Fo0PmRb+MDYM
um0QMZ853DGtT40kDfEX1S0s+nX2HVac2/q4eNh5igAnKeVRSEZzn6TphJvk
h5mTsUsGRj41+RpGtp14whTP5JpN9wRgRG+eR+DR0PR8iqSs02xfz/oFtW7Y
0hykbtUbTHJPMXgKrl+A7jExKmbK9D95s6l/cedugQvbzNONK3eHe5IRIQLp
0cEm+CtZKZWJbPoihcNpwFPTVEupGadIYiIKIxlLeqJsAAYmJF0/uxJBSWPs
qTEpoYjmhTwX2VNS2op10ZSyEUN0oC2vgzvirMIoRAZPlXbW6VDIDNtfPmoz
pD4JyyHd9QCwpEEaPMmWjdpvGpbbl7na54J54cMKfyr7qPapKT1saz6kvwpO
Stency7UzWCFLr/U1EZkQAGJVKPPvBt9AmciQw/BFlm7ONPI7FFjHhuGqLg+
k3PZYiSeLKHc0gTS2FGkw1fP80+jKFr6M7bTxflZXA7hKj9V1FFitMhR/q3u
anaxuBbmhxO0einvRbe4sFwDBuFSuB4w0cfiSvWib1ESHLw9o3L2g8VPDJKK
V+pFOEv0JiWi+Lyj2sN3U+qFSThhfwYQtFvvwJWf73YoO/o1WEdwjqqHEB/U
ajehdioH47wRlV9h2+E2jXgwiMvcr0/Q6u44LmmVdFxEHvkYs4u9x/kjICS7
fTp/r8T0HTAocLlslnTqhwHsY3R1RZkbSDc1ertPrMs4Us3wTK3FrBzoS7G2
ecnB70AabOutdL6v7wJKBaXN0g71AywraEW2HOpFvcLSOvgoQJdEtMhY5dta
ht1e/HiW3DoTx3/l/sMasb7hIeOIOds8TRfPQ8bT2gsNXGhKuLAWHRvYeAhD
9jWSyFI0FFfGCQSyfCNmBRBU87KA4dLkgNtPa36w1gsmnOqJzFZBJMa+u3v0
1vNKDLxnH98Rtnx8Qf3H55uUBfNfk5T6IA0IsMe1ECabVuoR0QKxoLtbfD5o
OITDOohIkLD2PabuRkaxXYHHnrQYI+Acxjs6rDM5Z8C3aaQ7gOHVUGhfoizu
etMOHGuNFJOzWm8xaCbw49dBr+/M3Za1YLvnXoLuRFiQaDwdP9e0K2OaBWVR
ZPBDXk/Ot8jE6jQTJroDl/z3Nh8f3t7RAZZ1/TNpw/TY8BQb8jB4MUz31kgN
HtQAEeLulb4en6BC5D+VJnZGpYdsC5MTGahJIqxdkbBzZtxRgT3+QbigoxYz
IQcv9ClsXpgJBQGm1bHXF0jXJv5x/CX6oAIlAZtmYj9yArryDRKb2/OYWLCv
e7eRDKf0BwuOjn7Bydjiaav2saXomwjEDtAIjIsO0kW1KlLzWVYzD7EFfBub
jeGmBwLYWyI/eK9R3YkpbxMgof2bqmX6APVoQIFTk6lXR/uR/MlvuMvIph2a
OSHx35fQC+PQmtEWaJ7rl0b3SoARtsc8iecY2Ph9eBznKFfcSGptYyG4RsSN
mPUa1NGvakk9RQ+buF4K4kqO8WOBP54wep26UTv0dSoU2dtgckrVqhtNbqpu
L5DTqIK7t7UPUrltvh4xLDnoSn393jr3PhJqKjet8gmdLj4sggdy175UPfoX
7kH/5MjRYem8iQfILIT7l8s/7N94jWSR31c6j2pAMtQfYhb9S6Y3Ne3SrDgT
IUdBvZy6JOtrwGghKfAny3JwBQarqY5oSYv/5awcs/iGMZ+DBHzfNChmMD1y
E6LUTFBCimZLvGryEOaet/71mPbJF+Br9yV3N8WtVXu+/aSDuGPXmcHbh+S1
E836+lzt4AdNp+z43dVP/uQ3D/4/gHIEcnzNjmjHLwabJCHCaxF0KCS9oTpD
D9Ruz7BD53YmrrT4zWWaurVpvkDXs2DD7N4zSbW8c7v/9/Yv4MC8fGUPt4ao
3vlFy43LVTF33X6bOMm6Ql/noKuN00n89FBBycdQOqYuN827brT2jaRBunLX
JWNMoVD6YmEDvJu+CwfsAOGdGL/IDxj0VMdkgEnZCPsBxG/JD/fTGZDnDN82
lpqArEqdZdm6QAgxnaSt6dne86ONnunyX0kDB/+dvXbp4SJMdYcVWzMGzwzJ
NT+eUlF6sOL8n53GSU/YGRcuT27yjuCdv7ok8fC5b5QGVZGSsuJlJPaWyeUU
0+TnbRGNloRHW/VOYd9ypt9mLv9GLk4owm6SM9jjDp5cOZELz2xk99fYsQ2w
CEcznx1IQcP7J0eEpelnqV6xdAqwSYJ+FLvsQeRJ4qjL86LoPSitEnFcSL6r
ofR6o8R1HinRRhqkkwMKi4ZYbRTyVtP/IgA8bCLO4erGid8HBlE7ug26MHim
S7L/6ISKgXJU2KgjDNz6r6qNF70idw5yJl/ZudSqRBYdQ+Dut4Um551sPwAN
bHuPeIxn2Z4yNKhhI/fd4cXWa/SoBvmmkArB6s+B/dJ4bNo4DdjIcGQxlEFG
ZatCWMEqf75lagukEXrgn4AJj7hiHEjNXy1z9NVnzdiks+k31qVw5s+IF9Pr
RJSQhDCuaLvso7fcEyOFf7YnGdIeynwxEFbpeC1VFIzgemlDAD4i/UOgdVDg
8WG/tq+jzEcoZ2wB996tXbMKi+ajH7hvs5SwS/lBuMsxWBw/GcvVX7p2NrMO
m/Ffn3BcvBuvuLJcnQGuu4SQ70bcPVBwtKZ7TJNLz48YdOzrSjWWO0TshOKR
i065zHtgXruqOgjDyLuQ38v1uCoh/fKLPE9McWDFbQTKdQm3HZzjHwq+vl6X
XZqS0BRPlM8yLYikxU8hA8TE+Oyf+GtpzlLoBpQP7vdz0Kc33+D3nH6SJZVF
+r0M2FL3g1pPNeOTMvNv0xO68RMXkUaT/R+C6aNjjwAj5oLADoURNcMrBGoX
d1t/SRKPDB6x1K9GCOjEoaV7uGB5hSVzxmJCR9vYPuDOTAtU8CPIC9xp0gG4
L4eBByC9mfQqSYaDRJQwBQOTrgGdG1L01358xdNcku+Qq1OfF81nOOjO4JtU
U02QeBzZUwkeEFulyeEaS2/2l5RbPWjHxMCLEN/OqHttfaAmOVlFAw/M4gJW
lDEckmIJjBn95ZAQKk54vgBA4E3KYvi7FrdQjPHPh7gAQSDy50g/Xf5AZuRe
424vdfDWcWTYBDSiNEq6nNhuVOecYxgPVv96PqXRUbvGG2pFJ/PkiX/22HeC
702VR1dhxAepmgTFfRqShK8JbYmC4IRN+RzgSk7Vpbt2ITYRC3tMX5Gw7vlG
QlXyKpLU9BvIMms80W0sXFsuJJIfkEtiNvZJgLhebAcPKpOKLNa4KH3oMgUD
rK/pPT6CK2cbxV0flomjMP1DD+l0IntJydEgJW9oEzZFP4wH/ZYH2cE89SWj
KFA2H488sGGljRT3nKp6TEb7rarGox/pphW00NSkaPcPqsXN6BPUzunmLgd6
PC6DZocFYmqNGHkydDXcYvhOqs5VsWdCQu2YCjJsr29KHDsWxV8ubFsRgwy0
HHKgcsX6NB5CHl1I54JeJRbw11eYGLk7MftIFamV1VAJX/jI37OP/4kgp4qy
LVgMiKov81cVk2dK2MA3eOx6Z/dFugQpT5vjG9FSaSa+ogP1Ckvnfu9GVuct
KSmEJS7LO/6+6FD0JOCjSzwdoe9JoBJcg5n77Oe/11iJ3OR7AQwK8UDsckSk
5hLti8rI1z+Rh8vK8G9hJ55H0nRbn1hT/S/B21iOCYs5UK9pL13ENWcfysX2
JKPLBYLlpV7zNTFJIDQ3K4k4P1Ba1I6HhqMgfJjRS3VAJjbYZFvsOg1LKqJk
2aiP8aLTwJr+FNKHdAR2QVRC5OITMfzeWlOcV9Fta7HZMDGjXmcqPdoHoiey
dFOqohtl6q2lv573esyeC8gBky2a8EHP+P0G/7WYizsYC/nmAhVgj7MMJjw2
gsuVZL6yZm88pyvzmmi6/AZ8ql74JSQoC83XprI1UmlKfOj0uDQbAzWhToIn
FUeGn5t1BOIX3OW6Jo9D1ZvgEuhqiYLJFCdEnCXoVvyVuGLj/pQbt2kpeYWQ
8mqOCC4SbI4jXqHjJ7ODpriQQrHm0VwGWBP1maw4BCqcn92nzgYmBPx2YQsQ
CjVp+7sZ6fAnlqd5TMQXRiPa/5KdHnfDxmQ6c85fxi+izJ/wLkvQiS+jxPL5
KS3lB3E9AcM+c1iXCmrNjd/hhBcEALpd1X4V9aS44+vh1UQ9a6KEX1VwDDq4
34sBGJd/VY61WyNYU/rljnnTrUUgW612WrRkSRwVJ8na+jDG+HXbLq8Mi86S
f+eUnt2EJQ7N8USwyX/EvhwrQIKipfkDsjZ2KAPLGi+tbfAJ+E6wbLakC+Ho
tqqot1H9cTO1tfv+l3hhoS+HF+lAnrNn0L7s3wjEsT0uPAqhnGNihghroINf
aOzPmZ5r6Q2RZRY/TwvZXb5UYKtIQO5I2j4ULhLl9Guq1qK/ufTaceGOQ09G
XVaiW2NheVQamQ+0BeZKiqwCnA2i344sd6zC6I//fiJaN2E8kE7s37CI4I+S
b6qp74baJRmE6rVNeviCokzRbxFwNp+pAHzfRJDxZXANhhYYOF3Zi6errZ4j
AMCQPnoCyYYmJLa4xtYomgSw1NNiildiLrNmEo2vQSmJcI9lNQooQKbnv8PW
FIfQMg9twQHggrKfs1Be0b5aaljug424LdLvBPazmp+VLKXxGZXKliv17kcn
dlzn7Ar50nH7f1CvPk7M+rk2//pbhExUOLN7NUTNiNW7jYFFcpjrkBj4rcVj
vrEZ0+LC9bjY/aw6TT1ZquKWIfqEp3AXnZ9jXvjBbKansArSXIOpEM0zegLF
N4GxbsQJVBebxy0GZQqUze/XxWVlHWAj5zYiuIQxHRYr48POUeGBpr1Vqf0p
YOPy0qWMMjnQ8oBU7+oUxm4Yzph2IXlIYlMla9FGCT9sUJg4CJKsDTYdH3HL
eOvdAeqS8Dn51jcJ+3HNvDb356dv63vpTokb2AKZY9auSeOPG2GrHkiSz4eV
3pJ2j9LAOkZiuZ5ZqnfHXfxm7o2qrRJk567bDqnhbktwTdzZvwDpYhGv84xM
ByBPTCDGltI+AlPOW1Ah2GjBYzn6Ik9OVZfKBuLEuZwkrqa2pHZmMLEkGXVT
Zhri+PQNcUr3T9fe22BTWkeON7AV6SPhn0M9mxtAYXbCB/z/mwh16B6AqNDA
sSMMOfLC+WBJ6BhpFtmXnRvXvWaIAo79DMMijW8NcjBxuDUDfgLo27mgjtAW
/N+693zB3tcBMWsoVL8Gl5KNlelvRpGp412063L7ddWPi9181N72sTqcnRNB
ZJmOsVLkDhxUX7Zsm8u2n0dn7+ekMNchltTAnhNKw8bsZ8aZx/gMGM9kml3T
j9UptKWMEsfKduJBYNCgyPZYIGW7+jMCaoXuKbvPrJ93dXHnbRo3Slzk+T3E
O+SmkdsvP/CfQb4hxnhZc9LPcF+F09FSBUKmnykxJkdmy2/JzP2sqJp2CQkO
45lhFPbogYwkvTZsAR4S6O4Yb/lVASRxABOSXT1SJJBqqhFo5iNoyiaSUGsl
/6kqMLTHOOZyXKZzNKGlX9RHCVMYV6lpoSETZs/Boy3+miuXLRPvFpscwhSx
yjlBRufn0g2rB5kTQZNGAqcwGJNX0ZYh2qNE+qeT0Lf1eZZr/e7zPpcWTiuD
gQtpNdqyLU+tr9+S7ldD8OYrm571osxOqUScLMVrxKW1Q2295WD5mvVuQDcE
0ESt6k37hdO/VBD+h5rHUNy1iOGiI4joNxmDRCf0OezSTAocGxrVfUAUAZau
SsTmym7t3Vuzcky33vL1qwDLxZM3SdRPSyxWwWrN3qRoU8zpbOCmSwDGg/2u
IXZZjkicMr6pCBDidfayKvGY2NKD0eyExxz7HBLKmatv7cGMoK5YzkvHNIi4
p/XxjqH7s4l2wtgk+Srw/4q/rBCJoi/fG1iNfeVpU5lCZq7u+A/DVtDlU66Q
8eomeocla+YACPUlaGBZHQNGR99oqTP3U13YewCzLtcnpfkizcX8v/oz7T4W
XHGvh2opa1bUMAucPv0yiMEwibEBe6nx6OkdfyEn2oEOla5uusmdOcbyKkpI
UkBGCoqvRGLw890FOUFw92Q6+9MpFeO2hD1jSlHoJ4fi//W9zhlGlL9tySBd
uauCX7Shx8flDhmanmA4QFq3ZMEtRlLh6Wk6seYJwewAcmQMpKhTx/ftshpq
gWMzVF/mxnTQYfaCzXIXdbszKP9p8+Hf5l1oPUBJt/knHswnk127xSzJwIwW
GfY9ksZE/BQRj6us4gYg+jqS34fd/iHirm5iUZOPAD3W90zm2AP/HZ85iljD
+irYrg3b7W3H1XRy696NRToyC1q8MA1HQsIbGEiXgwZdfmieWXEAUeheDyoR
UIgpjA3YyNpp4zkm7Ui09T5l99nWRK0EjEdK315np759CMigl5ch76qsFAXN
Iu7ocxDZkKJxwhobN/kGQTZlJZ8ZEBrpxR4t9p3YuNpygBg/Rybm/QnKgwCm
rCnpCXmdrNjBVwi631UszoCyVb3cqRPa6i2aXbS91mc50Br8wW4KHFawAcLR
0Ei6bo6aVhQk3q4/F7pgF5Hnzerp18dXlDp9A88vxMg9yZcG22U1wT43PNP0
IVW1Wbhn2wFLe8yYeY+vqzS07mq0xNvIn43RR5OeU54xS8xPgLVPYV8waAq8
ziYg7tSvWJdhAklINH5qXNSFrk8ntBq7cfPGxJZDWQ10V2EkJ++psxuIuqIt
oKGw+XIo4o8FUh8A0T5JdH8f0rYxlwN9UAqB6K1dNlBJWwzkwOnMD0JWd35m
qUWK67OGwrC9J88M9QWiigEweMjttt8I1sieVtad1SMzUhK0/1c8Z2L8OLRc
lL7j1+qf5q2Twh9dskpZt2f/UHfMidtiZH21VkLNFY/x7Y7tYDv5K9+OP7li
Fa3L394az39hpzj23I6VH4TcTHMu5XBJUuicd2+cm+IWD7bBfKdOLhXjEC4M
GBCgIv3P4mgKh8QETfbhUFBldsS/L7VqiZPG5UwEvpH5+QX957wYGJY3udsy
YFXvt3TvfrPIMlR80DIAHliFyPA1YNcxSoNmRXSGgkW4r2cOtjaxNiU7oqHU
f7TW1yIc8DPCnMJMPL+XWpd1TboGJXMLlA7iiqzW1eOo7BsokKS2eP8lncM6
8NKq5TWXKHHOBfQIJKWLki2u5axR+zVthOeYmzslyg5G8JthsIcrF/YoeHj8
jx0NYAlCuZJiPRUmcmKAGlBXKRz13+xMpiFRtVx+mPkn5tFNEk5PryT6foMp
0pct93WWk2dKnthfKqcODsXWkrekqxgaFuNkl2zNetdm4XK8JxZXA9uc8LtE
6oCP7/zSQZhxoSZQMmFFt/LlXVpSo7cXkWco0/r+FQtXsH5xZbG4dB2s/2Xc
pbp2Cbxb9VU+Q+y+0a5lOKqSBRxTPzf6sWJn2/tZtD0Xk2d0vrjGli3hiXa7
xaAg16Z2DEvQiEPljmpvdYPn2J8Cs72Fhdl2TLWkIQXa8UVr5mVIrcTy6wRF
Yhm6Jc8PCwH8LdEv0Gj1xOs/i9r8in8bidMCptiaQzU8UMzLBuxpsXoyKVA9
Rp5dtOw1c49eeHqv8UzpCTECmao9b1b5Ifk7RJn3mTWpdlgIRYkStlQHUm9+
ViM+HDylWtD724ySobmAmFqLFYBcP8UMxj9giE8WvdWXIMSkztVAox/zZbUk
hLwVgTpDg89OUPJ1PpqKgf2/8/tayHQFSqEeknoEY4PdXhgW/R2tmKpS3LLR
xu9NwqdNRcmna/Tkqif+RUCJfebqGw8hFJ3scemc5GZ54wxXQZj2276mYUt9
OB4V5hYpqCY5TkWAiRqDNpVaBJLEQR21V/AZLq4v9Y0SXcqcqKXptMh8l286
oxlR5VRPVVDQFyyu4GyiMJ6gio7RC7pLjDIctwfmftm544orkk2TSwkgfTHP
zwu6QtGLXDzeuvPSK/vVW8owvrw63q/6DC7Cw9245NmOLMDznmX8m3D6ruyG
a7h9y0rAapcITylkXErVlO00slS9mM2XHRCg26Hrr7zjVmQf3xaJhg1S3UGZ
t6eZrdqk/S72BG4CJK//NN/G8PkJAOwn34v8x5DZnyJfFNz2DQXIsNM5V9Tv
qIx/dgCTJ0qEdZz8MHkZTo7PFXK2osDV9+hkSCO7KFShfJ4umKOZhW68pE+/
KXYc+Je0okHmANowy+00l+KsgDLbHCD4E4M0GrR1J9y2eHkybr6aDA4LC/Al
VZyZhQphqN1KIqN05zE+UfhsS5STJhUOf7u6OmV17FymsjCF6oVK2YN40iq4
Zwsc/iZXIPXXbdB9hrnxWFPx9XePRGGto+dixiGusIfxYjbKbqi0aXnTr4JX
Un5FERLdAKjG1nYw1wVYoYay9UEdpIVVn8kl8UO3F96vS0QHzMZRZ32RDALz
xg8NyCEYE11CEi3KHtVgp9FB/Geu2Yf8zVT9dtqiPbcHwkrftWGxhms6d7UN
RV8uPzA2WRti38hOofVeFhMDWWyYQ7KW/2LkFVr/BkPMZiXaSvATJgn5Pkq8
/hjEm1SkEmcntC0okFkDWM+0/xhAZUgD1ZzqO6fbczG8XT8Z25u+DdSsI/5T
hPNN2Bfb+XyuVYwHL+OpkLb3CrvbhVi4ZtcUK4KRO3RB7SXLVQi/O+I7cO8V
lLyXvykoNaRxFtCctHjXovuE6CEoIMMLszXetvsGFTP62GsxSMuCpthgC6aS
muRIxgV6oLha1s888db1hgPNnNSIOeNznaUYt5EjbR4BzVjHYaR35r/fESO+
mADvBZT46GhBJar5IYjsVQFqM2ESyzdVA7jcwgZWDyeZoYSnei6Ntr9Ofiwt
YPncULB3tn93aeeeQiaZ3pylXHcaIQ6paCbfkZEqIuSJ7E7nLP1ugCjeu/pZ
4KsAioc4lXCY0AGzP0UsPCQDp7FhIGiEqmLl0wmq+41cewaxGDz58gT1kEmW
QhbyP3nG3ueWVRWHjzcVQwP80rzRowTOkGHwXE0R7QAEtweysq0TWY3n8X/f
HiUm3d9WAuEQSqtVMHL32HejSqt9rDf8QK2JZ8nEySUeHqYu68d2/GfhI/wt
zosXJY7VJudI5HtDtJsFVVq3ACGRIPt1HNnk+VxvdygCKhWZM0AABAD+gE0L
GDaFiVQDk72L6buDvopjwdEf40PVCwK1HP3yvP+mTbOvHWcr8zBFXtYNBohV
DSSxGn50/Hr0/tsc6WAchaW5sicXwg3W2v8U89a96OZBQZNmhS+7merbkKTq
Cxr5zFPEOo13UOF7A10PLnSiqExILdbX4SxOH3m9BEFORWWX0mFj0cje/fy/
4TflSIzTsS3YArAHkFUCaDhx+daa6gKa5V4DrelcSPT2/uzxmiK47x+WkVxY
Ux/HpD5Ty+ZBBbVFy/T0FHjvd8AKfUwAZJ7jxgYBiP447JuYpfkHJFJWX6HK
OrRhpQomUD8R91YRPYbniIuB2Qfc0MW2S5iwWo5OC9qzImhV+eoVZPOq8bK9
hivNFm0KaluDWG9EJ8D7aWlc16KZ0ZYJx1LA0QLXQrrZmBnJ4tuMWDESNmuW
FA2O3g3IrpjQjrnpvNYiPTUSN1Ml0wq3zy79r0Almjowllbcx+vYjN8ecpSz
/EFqMBhHhWogsKJE/OdZvYojKnKoJpY6LpOj6I2ZwLZqENHpj3nfTYcKCgGf
v6A7t4ERyRXwvI6Fra0W5NouwmSuIIJLhBXqUGZGIs2T5E409x39MrJfYyi+
wFewpKmx9zlYSRx0GWoM0HlvrjiVJTHQFuCGvglnvYq4BkkXJcBQh5ZKh0Zn
VfvQo3W+bxzDjvPSAYfe9JcqyOi95SoujsiHlQfRtMM0alEdmNuydaoZoYsr
mLn/uDbA5Ct3Ej4yYkRdj1oBMCugOBjNujXqh68jd2LS53oEvL3ymMd1McvJ
wfpulB9juQ6JkIDYw/bzSXv/nJn+CzpVOy/BRrD9CfPiDcvD18wZuPCdlY3j
cgJE6UPWnOvCIB+jlYTNjO80brMeTU/HG4al2zBv07uUb6D44IKTsxfqt1iz
jdDFRmSlD5vTYXgbzWs/btL35OXH4U/bLZ/57kTWmVSW9iMwcr7lA6UJ/EP1
UQtSd97gzTFi3AATUBFn7KM93WdqsAgvW2A095DLorQJtJmgxNm2n1LmihlT
+fPxj66m3scnfUtDTm7Zip7OoUGbO84nyzecEURen4x/IkjPySF+BcnZC8ff
K5DDpYaGoIiKjbAK71ew9R6UOVGSaJ4daJclf6IMille7F5WwKtXK2r9n0S6
XuNkbkUlBZlUF0w/iKrawpFfZGUW1brrtSfFvNoLf9meEgEbwPFqsiIKFfFw
ITm+7f846KxbJwqeyK+k1CaiUqYS663rote3hzTh7lNG9PqasiLkB67MFxX9
XYkFLybjmClC5DtweASKpog5G3cNWkGrJtAeSu8HSDDFFF1dlXa3ihPBksJY
G1XNBu5KtM8XL3wCoDv3gI2pWycdP/CpGj2ldfI3jZRXvxItW0Sd/MpbdkxB
5sKt3p7BUvkq3geeWDRPvXY92nACbDwNCtURqAXwv+L51hDxPBqVGsuoQcbj
/3/4+zlFPLF5K4F8H8iVXenZVZOIGiJRVBcdCMQH97HjzQw+5MUuMGmPzhqA
yxLGtCenEI1hWjNIxFHDwZA0B99YFsIevUwnBDuRlLzbCCcoBYhumFp+mCVB
P/lRTL9NwX0ifUbNRiiPDHp9zwtWTofuJ3m2CcXcX1gsTJKUtTL4I6bR8DuX
JHqN0B31sSp1uepXJ3SC2KjfmpItK4ja0W71q4B8dJvjBrfb7N6hc8B4aLZ8
w4K5sUVaJKiqjI1iWx3yxQ1nUtmsPvUWU2Xuvq81OJFaGsekzgdT/fPXSF1B
dPkN4Y6bstcevOC2DGwSlCYHTNQ3Os1b0vuuZIOnK14zCdyPyTjeNNdKErnE
9ybieg/PzSvKSgB87ZvVwHGlzynf2tPBgDyvgypfcOYMtr/LKqbWCS3E0Fpg
GDPRVg5M5E1z/Q+WIWJZaVxCGqV13F0vFrfpeOQA8xZdxE/WmZj2EW3p+HGc
G4dSB/WTIEyLASqioHD472QFRIrBWLW5xLJzUI367GxKoqqtG4OpzzZrZRpe
apdAi1w22VDG5Jc5zrEv70IcyHISxx7rUF4itYV8Ko+Xo7KEJRLfgXTYlIX3
PvDrHFx0gVidTWSisDwYhY+qbAtSu5TfTVMhJRHHZeC98ezyiPJzvzOgA0nj
E+1SHACYGQH/3uGT7soWSmn5N6sRWMrTa8h62e/xT9UDlGjG8HELvDvkpAaT
Mh6cgfnmm720GBrEXfQ1mwmX6yRbfG/RRKWpdtho2fWEyEwvGEHE7n3czv4/
aL9d9+ESMRKFH6ep7TRk+pje9SyDaDcInS9piHumN6p8kXWoUYUMzZErrBpz
M2MeiOLwmpLY+YA8HFWW/1qskTIMdApPvHsPB4eB/BwFgYPUIHPkNvu7Ioqf
k/+GZiHN6KfbNc/7UA2cfJjlyM5xkivvbe8tiXuBxaq4909+y97KjEVgNo/G
1p0Evq0nEXmwN09xOnlLeg+UQnAhkj7ZV0FWdIzFRYcRW2rHkeCP+tbYfvGj
xYVgGMdzU2wCyi3o9EBYO6eIgQ0P1MPj2Hp6tDkLtsqYLBxPROT7C5kYIpNU
Pn2L2sHP9O4metAS6+OLa8aNe+Bp24dFSSA96KxrLPeq5cZzzdSKaHNhlKGD
4hzoB+3WFWk9aiiiBmkEoH1tCIjaZFDsI34UaWNc1oaNW/qRhWhIFPd0bQI/
rBeChQQIefTS3nJKjF02w8GtmZ3fAtSpvWj/h+UbvE66Z3m/xc28O2QMtstW
CBakQjQRXLCV+Q90GZYftraan9D3Wgz5mu3qv+HakRSdP4GywlvtNK1j54af
WiIwNYl0L8OVYwEX8bo5oaNsGEYgHsu6CLTENfFsd3WSaJDCwCZve9ww7DnN
6efXruJtIg39Ho5nnNNLc0K3xdaPwPnJ1AFUfAdBU9ab90DDwM3hzqYpk323
C43SGs4TA/Px0tsy+WxQCn0q6RuwLC1KtZXExExjOG0NkeU990xysVbS0GIe
2QoDKzksMxy13YOElzRBa+q6TzkHETqsOUp5oO9y3yWRW68LETwWjTFYftoi
qTHqjiJX+1L7DM20R6Jz3+LWes6pV/70w4zZFmhl9vdqEeRTbYxom96qX0cZ
wMe+oqN3Qk8D4T49S8dtmLSPZDlrehIYah9XYAWVtjuh1J798+DBacavFq0m
wZtleWzC4fXMZddPOg60/taAixhaESufJ0j3eSy3X0efrEacXYxEsvuU5PUX
EK4i7cGQS9GXmct9bDiEdcZF87p31AiEzIKLu8g9bL9qn2zq9avK9vveJAlM
VFg5RFmFXckNauPAXOHZoEJlrK5zpvRDVwu6m3QQfbmdUq/dfC+pEYvKIt6L
9MXeVuq2CxZilZ+2HSRPxuvF12kGHotnEfOlu1O3KE163h6FPqB92juItWD+
63Uvq6QWXrA8FJyNRnauWZIAV+KllX43O70p4NWSa9zqgdv0RGbhNHocwrSc
kG/PXiOIBj4MHq5H0OOhKQkTdF7S8CtILX93707xF2/oLLpb4CjNq+cy6zBx
L7CF2b63R3LYOBFRdbLYTXixPgp6pIO7Pflj+VssSsOoQk7l3CsEtD1x8bom
lzZJDqw7aIl4MGMWsYU9Mit0Qkgfh58CL841fFAQdiXgH4FcckKrrTFUvfB0
Llg3NdAmnhcU4xHeKacGFXEGd4yH/cvh+WxdpAWHjOgzIEopcb2+EoFhxePP
4c0UDpKjZ8xi+B1yg3bMHJJA3t2bbFfkfHgmTCi1+gP3JxbwVMrMZ1+h9YwR
2arJZSPg7mDAbakU/9eBmig3WHmp3A6w2jZhX11COIjoyOPOXaOtpafKHbc3
nkSixo262hb8fzhkfX24jTTaQqXoEGwyM/b7o92nbuXAKDhBSiMt6r40VeLX
NVGu8W1gQS72OqedbFVkDBOBkTsM6BmOuYJooXJo7ovwl+0R7r+mmQ6H0aQe
nwCjJvJHB9F+7dOXujRIpt8RSQb82+5tFeK+wrwU7bYuMCjCjLxcq7EtTd3I
Ap+5SJ4shZBzSgIlHw0CWRogueRjUfCWJK1qlFzdhiOKJy2anG2DG+qrWowk
lIkjhhbyHtiYiIuFEtFXj5mQGgsAAmsYTePrsvv32GrjDmV5FNRzRdKKZuoS
Hjqo84c45MsdyKME8Zb4FghfAKbPibsv/ZDi8lk1cok9LoV15FkuWPrWrSUh
zvuOGdaI7ZADMkQJmNVRtJAcjStV8vm9TR24ZygBBe33RjkFIdv96D6EFD1f
gDMyDJcHzuH8BSkTm24h3ubjpTBqqixeXqTKJ6SoDjdlEVZJ9h5n6zSeh6RC
PERr5kjQgVItTY5uXWxmXK8S0lROw+Ya78FeQWeUIhTgIobtdAQ3hiyT9P6z
Bhlw78eRf3BqX7uut/xgFDFaszhwq7hyL9Qptob7QGAJf5QpEp2yIIbvFiN1
rgZTe8OMFB+imXv6MiDor+CvSKIMJAqf6gux0WumAc/tYCTgf8l5MGb5dec4
nPz7zEgmF+/13zVJnLTbdWSPfz5FNBv4MpiX1R4iieXgCVZHUULU2NR3t5mw
K1TkhZtZrtTOyibGRU0h4fmA8ZtPCua2rIkNtWxIqRyU1be5cbMyfyP+zw+v
3ovLObkUcXCciJ1FMFaN2DLX2bdRJKcFDKgpjiauXFlaHF+H40GDq4WBLOVc
94xlWIgWKCwIH+htWv9OWmMmRnqf9wg5Yr4bdzVFTiKSZ3A93+CvWVQijdCC
tmU9a+66k3Aq4eOfxgJsRA5ubD9bOWGZTQ3QZwezfVU33Ofno0grupwdvi6N
F6aX4awmNo5s3cIgJjKXMv+TRWZjLiWmcBAK1j65JaHp1UyG3w4ZwYN2XqpT
5rLNaT6+4KVyvdFWQfmzVlJGEXyx2gngv+dUHYtMcejNQyjNNFuqoG7fCB1T
ci7rIA5Lbu2VKRiczPZTCqrkEpwds/PUbvKRCpXO0MpJ4APvEqoJz9yJtt6x
lTO7Fdm0GpB+7LJ0trk7xlCFTGvh5PWnySoVCvL92KsshMjsHOpHtKjA6DKn
HbMidShpd8RFpmefzToKvYrU4WgLW+i+PTv/FFHsZa/43c+MNO14VPiQvQ60
ABKItJ1u5dJO5AqMKqt9s+da33F327WZiTlsFNcDiMP/b8UPPDeuoFrqSSEY
V3hkpi5a+QT7eAZqR62u3xYDW75cR0bi2UoARHMjy8nibnM8h5wZYlDYHTX8
i9ATkbQAKEp/I/fpCApmZt+MlWm2Z+9mw9hUUSUEQJNwGAmjBxJLK+3y1cf+
oqSJX4jQrq4jhdqef91RU9571OeW/09RjGwHgVpn+9oHpsUcoUhPXkAQwMxt
4sjNIB3bk/T967S9sipr7fcEwGCWbuVCBQ4BjCs/ApaQ+wnm38VeV3S4JkSk
duG+6x96mXgoSeRHiIoLkawihPXwMIuTBrbIYyfuJkPoK7sJLjY+CClctsSz
TtO/QYCTu7bLjvqSSKvo6leMSsgKi7lD28Z7rMQvyqI0RXACExXVGsYSC58W
J90GUuNa7yndPgv4LvBTtsIyXVH/dgh8FnAppWyPjg3klzwV9TmRcRGAPkf4
GbRo36g1C65TBXwKfptMDSq68kxrb5IqSqyv0aaYFcyhFd7xu5bunabBGm6r
9YvvEZ1uz8mIqIL8FjTwmYQ0a+WGDBHJB2aeVgFh+RJToQVEUthAQ2Sd53V1
Ll2hQLpfw3PRR4RPZ0b6RrTQqdPOJO9EzORdbROGJ+EcqWGkW/o1JbOq9M7X
lQlm79WI3TB9/oqDoEVOkx2m/FpR1j/J8yzb3fGIXlaCWWYAJcBTpzAsMeyo
rPDmTMW9g9PDLIVzQ59FaA3rf4lriLDdAfjys/4BVukD3jDXjQcpeL6aD8e4
i1/PKxklbXFQd9XiJXVMVQaIFvApNgVIYb+CXZz645VJWNjXegC8xyUb4KXO
V7sQje5y3NmnFJkO4hnqhmzCNpqrdFgyVWer7Ou0iTMF+RMRTR0H4XoPuwP/
nhT0RuS/jD1u+cj1Dr7RnZntXZejshVHFChqZdqVZKpYHbjCpUDaBmecPNIp
Q4D1Ne0cXebHn4JJYF+8oEQuhC+wqVRO91P2GOyUWbdu+0+uyvC3KYfedQZA
usXVlJ5DO08ctpcE67tNBMfKHK0xyj+XNv3tyu37hgWSpQIxJ1jV6F2hUDEw
UE5llOH23qvFvO89+GmTlxAfqWd6YUFHmwuUZN/7rE1/xf5fWJRAOAwvKzkt
wkSxCzn1y2Pni4fJbnAdYd2JM0Z8ilzeOlTU+xplL5zvThfID4GXO1m6JqRV
hMyn8vCQ3A4fiKvFWcLJM4zWDvbPRm2+aBJe+k+vgUM/mFCG4zQB4TqcdxOG
xLQ1iDCF8qUWzqnz8cquL6CXLInqL8bZSgXZV3Mhx/1dajOnjOzeGnQyiGye
5khuVTS1vJktaLhuWlsko+XCBA5Q/YEm1YpVXaeR0q2MXipE+bJZin8QY+Zl
ylmFQc+TMTn+iHC/RGgaytXNvwQeY7OYA493ScthODue0TRzKsEF8SNqd3OS
TwR2YhRBQoTkOkvUuNmm0yakSFDxyt9UPBwm/UZ1MaeSJHFjx8MR03BcOd2r
rAKMfx4y0OBBySHbDcyAhuUL6PkB6EVXg3RJ8ldVPSBcwUITKOposOMuztfz
YjomDd2SJ87EJCEZjtMdJdeQwal4IC5C594MuUp7vBcS9nOYhd6azTViYZJz
coSbvLdtYkAWT1tANqRN1jxS8jK/xZKP0crPh0QBRuR8TMzE/3/w2ur3fK2V
T8N33QEBP9Mkx0qoHdjxIW7APDEAJeghjoJXyaKLkmpp11s+S5n9WskHIohC
sCtIEH+nSCmdIojYpg01MlYxNpPD1K3DTdrT9G32BcYC0LIJjXVzNRhwW0i+
sgk3byydFO1cNasuE/qTbsceaQL9wb7Dd9Cl0yrHlWp5YhHbjfORCO0z3QIa
ZIv/qGi85i0oyYUFUr10tfIJ5D29flJZinJHiuK/+K7uMGAKFB7+WDCst6JT
A0RdQ2M9RfG51UVajkVJfKwNG/iAsNZyjE1BUBpZt28uO6tzpMpCfRf2z9Ix
aDa39R4qUDz5SqZK2eED6cjM/vjYmwEWK+69Vr/9dW8YRXAZIIVFfLERC+85
JctJJCB+nj19JzzV4IyNnAKjhiAsw6M1nVNE4A3R5Df2C3R9nhArS6U0Cg4h
/8GZtZ3wBjxb4N6cx6SgHuXTY6q+MHLIcFv+EkKa1v9u2QmcSjpWQ2Q4G6nw
ixwlUizmOJTcqYXILgMuH1hPg8RiD0w5zwLNmKh0jvcaFYlmwYGQIeiyG/Zi
6VALDSLsWRaFvQBnWSFwsu1ReDMpZhUdnQnou6XY9EdyB+bQFgwC/sYLhBQC
ROpgaBCE/7IWLF9UJllFTXVU93SpsFQycOFcuRddr1slrviGjvUUBlg9keXO
VtXtNuNXPcJroTt1S+92hRuHV5GqyX2qZP1rlXuy/W3lDo1Q9t5Is4cxIYYu
FckXz8mPCagLfk/5c0QZdsTAmgFLEzn9IbQBlsC9ttRL8wTYykFvKs0aHLVu
1ndLevhL6TN9D8/BamWc4F14y9hf8aN4ODj/86c5II2JdHajBLTb0zB5niM1
IuQ9UUmaUL61QzgSJJ4r/sQG/BlgEVy3Ap+TDcSKPVivLlcMT4WZkvD4U48k
vfh/ynM7Tc2Rd5VWD6vrT6ln0V62bWY120/92KZOSHpnKg0igKFbDgbxdNXR
A7t1efhMkbV3QhQuNZk4YbOyUSm3WnsFHwo7IAfYVvJ24f0bi/f69QS/rkmk
lZgWLzY1p2hNA8Y5fae07Ooq66aB1JOwKoLFdhqE9PRKfpyr3YlrYFoZ7cmo
PH7g7WvVF5sTXHQpw1dNE5M4Ng7QwTwYNm6ccCkvLziwoaMhCJnC2lk8TbTV
B+nQ1CtZxdOH/8jxXA088Onyg9LcQHhMJTRHL3vi0yFK/om2FGq0LEX2SIf9
R7I8hfN3XWkKEJEVn9Nmz4ZWMgAldKo00Bkzs1RYVhQpD+s8MnB5g/QO1eAp
CuwTllaR+bUXTgzB1Y7Y8Ktzi+wGLYFkoSpAnDk4X0fxRl1nwriIfXK208sW
jEjRLuLpuxBQ2j2pao9BJzQ0/hoBBXFqgp0o42m/FH/Hy8B3MtQvuf3X+WE5
iCsOKQ40zSO0VfH6Xw5y4+wCGJVVBp9pjutXjmyx9AEKZleSIfGoXqNwoAeb
8UZKyln89VGnJBFOwTtaf1aCUqpIjreERkUlb+fTmCEbbn/9k1EJpy/vrYXp
/FWhDW7rRsoQBz16l0NRW1hGA32axA62ZUIrn98ygoSDjBIsPYXn4tZG5drS
GSv0nI7IaT+AZO08oRgzHNN3mGnwkph4xOdXfGS7kJDQFvVZJwl+7brOB+nY
Wv03WHBDcvBBKhX+Frqef/zLqEuH1F3RKhxpFsuUN+2EKqVdqhV0Yuo4WDg/
S+3IYCdRaWksbl5/lcbPOkahBrG1bBUjn2knxAMXp4tUe8/FMkTcJSZ8tddQ
+xa17lVMUyIq3t8D5SireDjQPdbkcTecUuzb1wGOOso8sFeU0oP4pu2dHX88
GLYImwa7k1YTUTGn9DfIHhnLPqEdBYwaxvzWMiOk7yAygqFvjrh0uzKLpwj1
gdcqzh1I2+4ZuElvanfrISpij1f0Bx0jz35FFLLMEKq+Q6WMPKfJ6xzXPnRo
tdvO9/TUQ6XgCe4AExPwk7psM6xtQ0P6exPk1e3yfO3g+yU/J9aYK9TXsw5B
jEn8NWxB8dR3M41FsAQJz7bNvZ9HjDHH1EXPtgA2KzR3Z5ZO/tZmZ78Gbeih
kPRLTlzeC+pQvza9xNipUSDVF1TPUnPbT/UiDZ5UnXCc+JVaexHWvjE0H+2U
dg/mAYZuJ5/fyxH3H7Yd0AWWVMvbFLu/52bA7t9KRJRZ4YxAoIA32Vjd4jzF
OKmcTvTqIR1vrXcTNa0bUJCAOn6dcKz+Wy5EBeOFlCH19IzhNahabITGH+Zf
Pt0cU8J2mt+sgvwTLWaPgA31pTZEdYAi8u8yf41lYALWcxaaLWt4iqYiah9g
vU69ArW9wWz+/I6USObg+4wIjbsfdAHbjShQIA2kQBVTrf6TEaNn29L+mGDS
x04UVKjsk2xmUnxxI1Z1/z+jG6w8rRrnQMK26jukTX49QXNE19Ni8GxbHdpr
CyFziQoNmTGy8mwyITsJkGa6zZxNaycytZF/SlghcNYcG174rxw5Q9Rz/yGz
eMu+aO5/jBsywbqbXO2oFPxn3T2plH6YbxuD4cUBhg+WAjz72bEcCEsVBUcn
5XdvrQzN7yg0pHVHSsUnX7594ZDbkyxBQgqp/dVq7Zc8gh0mTBuJkvVFWyQa
JnSGRJSMEEah+o8UEyadstFnSys63oQ6O1VPxx5lSF99XlzxpMiB8KCn7GeE
XBJ+cVIttWeiVNFLrL7uh1G8YyMR5W6tP50CKIAC7EBEOMud6cc3uSQyw7+R
VPMKLPf3Ld8ECSe6wRc5OdIR/KabgzIrVwKtOurJ8F2i+TNq16n43Pu2zrG2
FqtCnow0ideCrTxwF3TIndI/XOyPyN6SEZnDYnwQ9nxYdZLWg9epNAQ52TA6
6vbbzB9agn8pv14Voq0uI0hl7OKgfh9qOCijJsWMDiXUjW2o+HCrwTW3t+5A
YHCGnDANtuALRoC1li3oYeKrVcQ1Mzs3gwqfFODoLuUo78LqRxQ1LNfUac9n
2u7R0isD/VWrvkm9xRTpuCkHfJaEL10SQgTZ0YJCVUfPMApBnjpZfAtpvLlH
jZznCQ1YrXE/HoKuxLgQzIgbGP+01InXarebP1DzH1k6O2FD/7lNeJkqUI4m
48F0o+L3WUWRUM1biu6W6bmji4F7U2cAijMzrhCGPkKS2DVU4Bnhf3R7ct2K
94ua6kxxXeoOb3VUlSvYd26Esjg10sAnby4H/FvGJNa8TjfWnAGekipgtfuw
aQzv8bW2vAX98pqUDW4fCopaulSGKH4pBDJlaESbgi+DsQI66OtXhQUyWSFg
MyOMlnAZRENhvzTl0qq51uATAGsWtojgk+BiU2v6VXlPBR/DkV/CmeWeKweg
UWUW3Ty3rBDmtR7QBLost3E4cBZvieYWmTNkXJJMBUnFOAsB+43Y7b/H4lS5
UE720p6RH2EK/lKl19RoMJhm5aZbKRmMMTTRhf2Wrb4WiaTqMkH+1MzDdlIn
Fgy9DWj13hn8xlWXiXt7HjApVmpRWne1iJmLjqxOP2Yi6xluowyV47PIzaho
fRk5aq8Spbmhl+mmG10wAfYkMP+LzIg+aR4QcWDoJAlZUkF7naKmNg19lfbk
wDLffSZNI5+aIOPxgEFbSBpWNpwdkXz6ujWIUuKTh4FgtqR4tBA3HLi7zC5m
D7wmLlViWjUCFiXOn1ljEQ5ikJQELR8WegzYdh5+FtNofmI66gyF8yE95FQ2
1ouCUwmyw/jkofu7WhIwao5eDj+jK97Go65jb5hjPxPJqAWIm5eLXkuUDEsx
iXMPDycp8+VwrEUL4/7WxgvjQ3UZdWKTK9e4y55baQKWKa6IzsFEW/UFAlDJ
xBmSSiYTe/sRME5DwoYXH+S9zysmP+I2GQ6/SEZUWOdQBENFgFDYaMW90BgW
LemGSc3q552YlpKGMk3JdXJlH1q9O6HkVEMjlfTSr+HDmQDtnEobc+1KrzW0
eSERO8nkyxg6SGuUMMx76zYumflqjQeJEP2w83BWfRMMJ6L/DY0t4eXX/NxR
qlbq2ZcvEdbj6sNqWKIdHzTH96H08XuBD3QyrBrP8VNwMOJyY6+BAbYAi5fD
Dsd7Xx3jEQRs1dp186pqW9sm5BGKiNkQ8cc4zRtxIzp+ZGdUS1Rw6pPhWGru
WNuePIKA7icSE0V5ZifVS0vRmPCmfitX3UWqNYdMS/nkfp1l+LrlE1GZr8X2
UuyI0NGFb4TUUlaBZW5JBrYVtWrmAl0IgeJj0O2hLWGpxMRMBOH99CZg6a+a
OAL5exrwBCTDGIIsCOkseYCgW+bXFoLnN35kikNbswGEDR08ti/DHe4QLF1/
/sRtVcUY8FxgfisxqRRFjAKrxtxW51ns0CeZqvIBJGQbiaVV1yZTiZYaBjRj
opIV6GFd6eqI5VpsmqYLLEAn9OC0Y8t337i4saM5rxq+yhdOoh5buQJ8AsYx
Szmb8rmvgsAqK6YTuwBLIDKpZ18drucHQf7nwAnBwKR/y5YCvjMBZIB+lXXP
Y2jpUWj4UrRSoTdlkEFflNp/cCKF4PLNDwWC/dqv2k9TCwnX3I/Fka+m6xlV
e9TN5471fXkTmv8mt3ZcPYlBqfqTGNLJK7yrhuRnNrWz6JiEvYF+f3+H+6IX
XFJobRdV1L3bwV3Zefj6nj7Is9hvusE4zyM0SEM0PVnku9Q20PMv2cfuNyc1
sb2XQD3npreBgtztLKg11Mxjp8Z3rFEqSh+q+xFIZg+uRmF+S8i9O3iQmYcp
C4FzcVh2p6XGlXFClZ7vdqtQlqBB1o5GC39vLucJQFQ/JRkmbLaFDPT3KFbd
wGqZhs5F6zu5zSaSno9wF/jUkyKIVOm+bckIv4YXBXOhrQnh0wbIk0cBZJco
kHUIc/ts7nsNtXyrh6/fW3zkJyA7F+Z0YgNp6ZtMLVJSnYxjz2iLIeIFizeQ
W3HKCFgwaTudGwOrOtGkNul1D+heMrZbs1e4ggPvK6UCAiNvhK0SvQPdRJox
6oyVc0XasOThW5RqT50M1dhAraajxmmchfZ0UTfNbtxyzGhDbNgzLB8riW3D
KDZaKvyY83T4bbdji/sN9Gevnj9mQT83VTiG00oVYy4w4JgbDIqjMRacR62F
Oe49KXe5wxzlc4AoLxZang9bJp5aC1lj2rw5hLz7/VXzn+ApYE/kGp1W12kX
U1GLOQ6LJ03DXSNbQTy6Mymm52f1l2axIaRIQxF/BCGvmkTrw5f3rcM6kbRq
6BTT1iRgAdtQB4e4L4SLdX2Iw8jjZ/lfO+IaKVH+ULwrXKSFQHs6SWYtZOEN
bZrci/1lJnYuY3I0h9yaloU8UuCQS7zM4oWKlbQO6nR/4c6+uJ7gFmJKOrdR
ATs3F/pxQdcyAWfeibLHvGR9i7icA0iYnbLB4NZ0s6OlRfc9NDDLuaUDFk5L
1TF/E0ybJVg4P87aBVFe8y7SzGC+81yViroyfQ/3pDi6MYUkby/Bgo3Bxdvj
VZQRLX2PQpb9V3jq/NpjiHllFJaK1lmqPjBXFpc2pfuhsRC+pHSS3gvrqLac
efqMj3KeLtoFvWlsHjaA2peBya+k30GEJ+5p7UFTCQEE0irui5PfHvyyh+Mj
xSYluN2CeDXYJDlZnD7pl8M6PZ1qbXK/3lJw28XX4R762DP5Nizug1eaTVej
VLzpLrFIm0GZBrgRHLhwDXypA76r8GHhWpfhvCNh0mBtU7T7kCxE+gzKtVRB
EPxy7TiBdNdFpe+qYI0Wyse6P6SfThGAKW41DAIRQ4jX4nCBW6d0bzu6GGgl
BErT9UUPxk8xqri5VhmBGvl7ndT9xr4ax0e6iuD/czKJrk11DO0nlaYYjAKN
zJmIXQhN6e1RuedMUFtuwIVJTjJ1TcNdHuK39EuhzYvopdL5vkAM50szz6Wx
MLSeRJJU4YtXS7zY2KGL5w27XRecLA2TsNxOUg4p7L6MpqgidmZNxBNGNi/j
285wzWR7nPGOUXMDvd9vui9P/GQTWeLgqewaLTzup7O/lEUEYiCA6f2sUqju
CepC2yOZY+NPh87FGAajXKgU8FanjSOWlknBbm2Xwc96crfPwfggOh/T6naD
7lipg9HXv64xqJf0M3ZeN+mOpYZ1SFE/NpNuUxhvA/ZUh0hDiQFL1u10Kn06
kr7Kc6tYA2INGgUBbj88/xlMr9x0uJyhf4nkto55tc6VUyzlSnWZ8aaqjiXG
N4eaffpJ6A4o8xs6vYjH4KPxj2YVD5rGuCHhGGm/U07zTHsZfE+WU7C4V33g
8N71x7+JNSJwbz3VF1T6p/dViE7+283PQym74JcoyjAlTpStB0kVX+Fd2RMw
VAkp5RJ6ejTnRm3nxD00V5/nYOeSqnz36lDG8f4tIxz4ZWqrAuCPBgA3vdoQ
0OdK9SftESPc0mhN/XEuHGnZrbtb4px01Z/3fmZMzQ8A3eQUcqHhs8OGW7J7
SvP+/Tikq6VHgpvQq1+b8hN8yESgIHaenrdrc1hyajAAwe5s9ubpP/jhSJOA
MrjE2fk0rOtCNKYcHHLZ01WpsupLJ7by7LIC0ZBd5sXyqbzsEYRZ8y/tC1SY
PEjZsH+I54aLFuUWdsXYxwsJ18A6Lqf4KlVZZ6CkaVQFaWhUvJKRslRLh+2v
VTfCvwsQEcjEmva8U3jXrcmjWxDNakvlZipKIoG7PVUeG4ACvzOsMaxCzPkS
lrQnJcbWZc+YqyqyB++luTvA1ETW2Bh1D9DZau17nMLJNenrhV+d10sy3uoL
lGpvS3nHul9MXP7eE+RfEr2L3YjDliIBN4xxtRMNm+1e1pHxXOjT895RcVsX
RTQkGjv5HfZm37qLUSHBrRTWzEAB9hw8JpN+HkNXq5iG2oeGQEu383wDdLJC
0OcgOk5LIWJ48s6pcsQg1b2SMfA7HkExz4VY0T7bKEbeJCJUYOaFT+wMMj9N
ezckeAhUmP7oZGqhIqeNaqUxn3hULzD5rjMOpC8mAQCrXuHOu/2q8ZWdl5tL
M7WNkXxs9cVz5hMz85vXr2iZq27J5lH1VBxNk6Lolqp4Q7oIvQ6FsQxUA7Bn
wRygB9jTj/yBe84lmZkDTR0T6PHxbNPBnRCRNsfMEC1QDHKH6ET4Lz5Q32aq
U9kG9UsL/GB9dy7nw1qdQFn/iVUCjsUXZIRNj596NuOCLlo2tMlGgZQroEdl
/T0EeHaxwo60/MBzcTlOcmvNBWJqCF3nI9h7CuhACTT6lh1xVUzzl9UcM0JF
4YAbd/QaDbXBDi22Xt3v/yZ6PdxZbxmVApYWxxXrXvCfJ7E3hRiA+wEtby7A
4rhE3csPsrsUxkA59a2BTV2SF0qO4IwvlIx8jezTl2logo2wN5DThx5BrP8+
AiNx1m9MWrBcdKo/uriqRAiVKypqTd2KRgHQ6+lfZhkK6KMR3WcDAWdSH7Rn
JzaRra3/nf7z/c3e/Bme+J1JDwGLRWFJOgGVwECjWd5LOIrUb1CUboxOdqQ7
rrBaqQ12UELRaygBkV6DU/A5Op6/u4JYXSol8mwibaN1z4zU1I3IJxd9x3hK
UV2JEgXnuAM6bbH/cjqqz/eQecpXsu4wuxIgSbIopttttsVzAQjNXYJ8biap
WJhHhec7TvEVHBjkM1mo0/aaaKQy4adtpJcLba24LtmDnI15r2oGIn3XAbRd
7pfogb/PMKoisjz9e1gTF60PJmX5lFXMeNtmJsUd3N/do5wOs+ddjOSjfmiv
VfUyEqaTlSw/W3cAH/QCUlSbJ/wWF3vAgPiNp/u5yrNlVgYfppYcI7csvW4a
Ev7M9Wz5SiY3heC9tyD0YeTzdszvTaW84emoiwnhQaBeC1c3KFHjasrynuiK
GiwepxBW8C6vDq/gYqtufCQ5YzhbDKaRuf7jsFjeCigzxmwsgpiiDOobKdka
fXMXWxvVzVdIaEAjvK65DbA5X6HaIHKiI7Fefsx3WNkj86Cq7piHwaJPt+DH
FJXi0e4CKhw+L2/ozI1Y8WmOvt2yyVKpoby/dTAV0WeC35WRqVgbwTXz+l78
c9ibwtnm7gIYUfcDfypQT6UncoxaWl4osAfVWufkfXYzGYM+DOjYCYHH3NGh
7STZ8OqTugZiGF5o0OGmhFPyNE6MB5ZmHZ3t90Xtoq5P9v+v5vVGuq3Oa3r1
9RlT97VsyxOt4s90OiKsTtDnQ3wLelyAdLUcHrqCVt4elQo/r5M84kdDe8qD
90f8PaSqN2qLWEsvzVHevWo7lEq7NpevL2MaeNt695Y4zhfAns26RvurvA/1
CqDnSwbPLZw0R4gJXfPuQImKSE2ymrDsA/PPOrr8LRDmAVx8LkE/Cu3pJvAT
9iSsPSV/kxoxLoduVYa4xE5zEmW7TcnEjbpnf6HsMx/3kF9iQImeT4knavwJ
F7eAU3Tf3Zuvz+S7wTtbp2SerqqErk5XVZZCoihnG0r3eYRLXKgxPEAFnDD9
uMxL8SS2LLTk6564CBtBWUTmghWjvPPNEBUIKhqVgmYZ7Cr9d/QdeH9wMBCC
h9RdyIgIXZozIN2RK3W9R/cWQ0XehCYf12jl3cpJ7LPCNu08byqi8fMbfBjO
9dojISXhtiwybKnj4BxeB1fom0Vdz7PXEZac5SoepVZRn31PhGIu1VN4ZVN0
Jv0Ivd0OSml6WN55Bi2G9Z49ILyTwxeVHnEPb+iNTtxlTYHZrXem40L4zzxL
9psNvEB/xb9HU6kpkypMlzp0yb41sreHAK3x0frjr+M0SlK/f9LT9HqoxxRE
80aowz5oIyDYZhQ31g1IWergl21gguN1pQIweGBZFeVPX2vHiZnPz31xyXXV
hQljKP4XltZFEubew22h7dR6HDREpabJXgwFPVNyhIbC5GTfP6rhszoLW4lK
7pm0wtWoFFt69oc2ioR7Oo8Pdii0gf72XrCPkH484CMba9o1v/SHez+0rv7g
zCD6yr4+KqoWAfNSTHLZ0XQ3pD6SHq+r5bW7n5doLdt51pNu65zUHCarEIRe
o0HkkMcRHHsY4Tadotg9Hsfvpqv0WpdtEOtI8IRQVHzSQoK8JWcDn9qVSaTj
HdXrAgD/Va4rEPp0qhEWRx4rDnxMenkV6f0sCr8iPKifiqa/TEIr2e7fSseM
U5aAbq1HlZSzN71Z7fRLZYp4mTV+dsiY/wLK6G0X+Ny26sAwZComLO/0OyVo
lAwm3EIksJ/iGnEnAn5WLmsKdyf99N2C4/c8IQipcl3dVz0koc4Q/wSS5tt0
ZOAXxsxz5QQHWI+StEJW+NEUPpCuwfPnDEo8lhMtzXTN5Hj4vR2YW0xDc0/2
Bh95l0Ah9elyB6t6lrmL9LqWwRpJd7fE1rELuWMKXZ9xu+XY2AruuSk3Itc1
fB1fOMFMpeCoyj8yvSVi1Y8CEaT1cCpGbCT1/ZlfKwr44L5kSgEQqiYix/EB
o+Piomg2tHcnQViniOe8iqpmYIiCwBRmYBjp8ojO9iu69XmyOUXnqFUiyU/B
Q/G9FUpfXjYpsw9qSOk8E4u9d+A63B2jflcapv8BSF6CADaoN2cAiPDLLNF8
bPrzfFhEumWiqzm+eDAoCiKAPZcqb8bzGrt+DSDHwNiJen18DA9J2DSFk0FP
kElTu1q68w++tnvusO1cyjxlp7cXlfR2n6OYiBrE12P2IYY5xpjuvDTtMuiX
RujinvwTLvF1UteoaTaBGWgcQX2hI61wYvgxlJM/D9b1INxU1lrtKeom+KTp
sEA11XvkaGYt7lWlkgp/LfFUqy2wA99FGbr7duBELUCCfyj4swC8SxEXWqc5
+P6l6ivzF2GyTTAxa0J7WPEJBJMplJWakxK0nP9cDzQbTlIlWxL01Dwv2TtK
uojKyoTqXXTmwD8HE+QTVvVlnFIitTFkezzf8NLCAV0Iu5d2GwrbtGMcrrAi
zuIFRpQ/UD3Ndt6KiEw7sodL/QdG4DUNwbCRpeywboXvNpHWGXTRLRzXRFvU
cn5uACAYs1e3kQiugba9qWkN83Sgid8CZB2dgD5tcMg8QleAM1sUyB+PD/cC
yCjdfGGQVvdEjkvKvhq+2Kqc117DpTsoiYPl+uG9juk34r72PWg3zMD32O9X
lDDiGNcbdikQhJaNnV6ckSCQp1Ax8wz0rcCEnt/LOxHSeLRGj/a0Gtq4GRwT
Oi//S2WcDc5YjMqOOWOl4yAeKb8YVpTNRWEi/E5/oiDKN81ckxu4WXF6TcjZ
3CFM1ho8fIbu9YW0/9TpsSTFzc1A+nZaRvVVoSyK2G0qX/NmfIcwMMxvWlX7
E9ry/pWQTT62VlvdJbfPLqNFN498uNkpiaHl8lUrE3Gnsj5gFU2v0nBwIDWe
DR0RomN9PvGWMILD+0aWccQEC0+fC3pim+vbpKa50ER3GYeRHp++5IPnRG3Z
NK+l79BlVdsBf0PCPOtwENOvR0N4UGC4G3g+wbY3DkwX+On3/WbMOy6gVfRM
oHjgFn6EkQw7EqnK2SQinN/aafaQ+stxmAWa0PLD/TvbOTOGC4wecqACKdFF
ELmYRgikXGlkUXDliUmtXr93UrOUoCdVQ4FRepsncEdQICIdlXbKtnBcALoB
zMlnWIXwlAGNBt/RTOo1TjtjYQVMBQRrhyHO3gQkV2Nt1feZeuD1oPrB5G5E
JqbhEjRkCiGcs4/cEXxpRza5ZZL7hsbhAu6FI82dehAPuOjvPmsmxf8A3B8y
a9RH3LFpi4MicGJ5bg1P914dcHGvw8fg7DSvvcxE3/fAmrNmDf7XWuvr9Nih
OU9qGif28skbwkasSzB4tKw76kiiA1DC+rKFa82bT3XlB3ieoClnmn7QJZKo
XoOWExVVBM9gYMsa4lkaDbwzVGiMKvOx0INzFtAGIUY7Q7o4jSBeeX0UhJ3O
Ls8kt/4v4J3IraGU/I7Cm/YaMZdx5E23+iZld0FQWY1qaFlfk++VKnXSGO3F
VO/ovNktrQZUTm6CHO6V1Ihw9qGHziNu7yPS4+6DKQoMMIxEZzvS8YfUqJtB
+57bNoR8ZaGkjIXyVrXYvQP9Q7ti5Z/eq961maL6n4evtZpbyCqy/D/Xt1fb
uhScsD8iDopqdHMvHAJ+gFLKCFGljcXrtKOM10DF68w+TKZfoQfMsZwNDVJU
MCOeMv6a+J7S0qkikY11iNtbSe0mkgGmGE7hHEC5VP3AIt83fM+cK0WcQea2
O9is6n96H3djc0fZJ1Evug2IEWYZhI4nY6QbHrqf9WK7MMMhJb0SSCBg0AbI
nQa/XmL8R0Nt6tK5Mu+qwImSA+OMLmLttB7Fa5Ec+8IitLnzMBlBbYmDgO1M
tly9qNQk6OXxtNdVHq6xLW2KfHu/ikf2VixIte/ZrxafzaWX4f9zWypyb0Mg
VM51aRNYvuNCS4QybabqbW0fF/EpqzibDFig0YmQOr0VoBeS89sn4rO2imt2
XCj1C3fR+xuXSC9Te/zhzDWCm54TV1/zmvYjV5o9gFKNmI8V0LJ/ZFDLHMgK
evdd3Nz58lhFY5f0Jn7s7pX7/xAjLbKSOkLsNMk4GNtkfHHSKkH/HfL15Xk8
whAecfDnc1+au/OAYXV/DKQ8WtDOwH35dAJMlvH3wMv//zWXHg6UjJIL7/Fa
QaD/zB5WrllnaeGjki1Ag5BFwZ6V6WVeXI4C7UvKDS+NkaTZta+/iCKebQdA
U4lcfEptdu+pWlGUpsMBb8y3S4P40d1COn9fKv53Oi/o9UvhVQ86rhBZB+ng
nRi4hLDiFomLTQpLLDsXQniAWXrSrvbpVHL7tRYAB0C44zjPlL+Svie/gxWa
jYSuELHkfw4H/5wdzaaHeZbIHNJTaV3PoW8qEHn0+Fbav38AO3tQ6Z4d6Jl1
h2zAKsmCJ/JULmuqdWhyIPapS1Qh2Z85wuTx9FbVDCWkijpYrby6zqn0Fwt5
89X9F2g3V9lHxSLMr9T7SM8wVOR9kfDMMakyf4s+rDZ3QnPd7xoYWqUc+mbX
OkPTgRltFXnY/Elq4OTmPG65QO5pSnKQUUrBfkpflXWqMPGAq4a9WJ4/Hl1l
2o/7Sm/JwEpJ4oYeg6uhPCDVhVIqgyX9TUr8G3+WLB5BdaJ9DZIZ4W8oz4wt
1F3pwGaGEhOjVWq85XeHZoZO0V6lD26MGq1vps/eHZBYY/sNk0losmZo3EVf
UXRTpP2FjqSxxtt72kn+LpW63uNvP4fbw66CJcqz6iuWhyot1d8OStZzS672
RpUuqjzJWPKPQVJCszGuhoRF3Uqkwjd3C7RTtC1E5B8k9hrBWz86DFwCOgM6
DPTc3Bhu1xwjYsv6wseQKjEbYW+wYp/ikaXHNGOnabMHiIuSX8I9GrJr4NdZ
/NQzZvDNM0znC3YjifLfgK9BaHhTvFCB+Fy9w2t300/A17m4zbcr804DwOaJ
8vp0tIZwRMEce0V/xZWaOzfeie6a3vMmzFCvtf8XBSYWH3ztjma5aez0Qvo4
xJ/Q+vbt+ZPiAGvfdRbn5u2r1PUQWLwSoLAcxW/y5Ogpc+lTYjvprwHmc2b4
WPNnhqKOYnqePr6eF6Q0mhSJGffojuD3k4xwUQ4TqvuWzJzGpT+5IhDRBYmQ
ZjwIpXNMnv2h3yg8WveiVWshB5EYOOrZycEfTDnbHHi5rkePvglJvQ9wPdm4
Gq/VxsIo79rMnQoCg5pr/9Q8YVkwT0jtu3Ko1pDLS7JHqnSvc+/RhigYCoKJ
nt8LbKbaGz+VnY9AMDXMeaVP+OZLrNotUzrPDqykFXIbvOwntGrWALUQw2s1
LaNfan1/2BniaJem6gqc8CAGybWusqkrA706huhYX7GhMUA+Ilw1iqt0xRwD
pChK2JxiWy6hfI2DrzQPan8RCNo+8i0M2LYw8BQLw2hJSJJhWv5ulkGNUCla
5qnMORS8P6Ue1m8M01iVxSgb5s6W0ehjbzYwHELK7xqcJt7V/fyPZpRYC8e+
QnT2B8hVV/04d+QElrdVFNdwaoNaDRT7InyhJNRa4+Jh5DFvWhcl9+GfNjHi
wwRgT/GID4dYHrGk/JxV1zYLY3wH8NYcy7FWfNClhJeD7aJs0tjme9edAmj4
vrSknvXft9xmZ38wu8lrX9EHuLsncdPmtxpZYm0dzR7tsBXEBVukqNDl1oi7
3S6G4zP6V3Kz81ViqkyZKuZejFEJHnTOiEwBHLBHVAbJsYJIk8S+QkL+iQ/a
Dsz0tcONVX9IP/yedy8rCDxb36a4vorHfR24M5EvGUf3Vk3YbwJlICZqcYEy
t1hccV8oxC0dixF4CXJyhs3paqYIYYrkO7mJFzGDeWYeWjCOodoFBQFaVqyx
cWvTjijctlZMO3DyN65iVm62Tu/R0J4Dnqw0i4S0KrmBGgN8KQnHfGSlBevd
R4tT2MjK56Ri8Zd4uHTmQqWZUgCrQuKU6NriAvBM99DySCeDUyLIRCwuJNL9
NcMa3mG+jTmkKGqk157uXpfs3NtR5+UZ/dBmqout23KBc/qvDVjwsCwrQGRm
gIj1vrNs17vWqVlNykFmx7ZbSt+tcC9iANZ7Yu/eS/sBlqw8ZxwoIOC+nWq4
VX9PRHVxUlzyV4sjrdx4FnfuxI8VkUiYo+pP7KORjQFUPmE0fqT+fSUzBKaf
XhaLoVsBtmdDN3QvY6LkT1axUQR9WVQ2Uz/zuj83Xv7UjNKPDOWmN2W6FQEt
vBmOgluCSPHT2WBElAqpbiyhHeeW/8Rw3jG17nCoSEHI2nmt65nSlxSOYABn
Sw4ckgZshuoFUasnlNEx6AiNatKDOL0xC+gzD+StIqRidXnZAVmWb6gSYPRb
jE6UQ0zW7+CuHKmHWlZsxWJ3DxxAwkBA5GT+gsRA45arZDVNqnaHmo5lkL6m
lhgb7LJuYlO7ZfM1bsuhHJujy9JTus1m31tyAQvkKss8r2Dp8Op7icNDX4hS
j51axRG+SykUg4He1caPv5k+HRl8N2ekWgXGa+EXc8lZAmmtGDIeQ6W8KhdQ
0zuGy1tpo/tpsiMbxPNOu0DTUoasG9xh79NEY81Kv3UxCSZTR1QQeFcLn4tA
TIt6pfzC903FIIp5s1Ek34IufJx+vTXdUyFusCU58WBvPRSY4KSgZO1UFMuN
V/Fctgb9R5hLOYRTR1R1O1hqupS/f5a9YThcTysPAzoi8mMuwy7CLaHvaZAi
37p84VUV7jdZ0qHnYdq/lwyQT+etRKr3As8T6rE6i0X05nM6D5FGK4enDvE/
eUSW+yKobKxCn5quJxqaN+UeLHKFzdXdP7ZgUxJHyCGc0vJczxq5MEKWDs1V
SqiNpz1nZW4hgRciqyfcMTOa7uddAwOXV5ZqVHAkTEpbp3JSzENcqLgz6xti
7gF0pY6mpz11qlUFUtQG0hvgDIz8Zz7ghP+844h+MaYIM3cFLSMAlkfxsKah
/IEhvU4aZgUMsjU3uWWcOU1Jio+wfM+IZxocZutmcgbirR9sEj+9cN6zwiY3
i5KepOR3YwqYVFf3Yn6PK1o5rC9YTnmpPX9BEQvw5C0cyXGWqX10AiZQkGao
RKsg730A7zj7NUozua0bYp5pImdcMEW21Fg4Rg+d6SN1sXFHJzf7vGB1PEkV
mIcLBbL8Ok4cezHDmtje0PMqvq4f6IModoCs/JuwgGRkNpPQ0KlGsZ1bNvYZ
G4Ir7N445hboQikS5dGvw2jDnkYb+OoIKav5ISmuKcTIE0sEJryXLBPz0sQP
2/opZPqC8ljYqqOZVsim//bkBHwEztsp2ElZVkOKuFHNypyIv4by+ZkS4Htk
Q/h52w7M0wUAGJ51I2BGVzEZ3F7c7lFbtqFXSeZ3gaJxntTnOUpDXh4mE4sW
4V7ZwDriPrcf0nr4ppSv4C7bd5efuschMbo2/rzcFqbMMwXshec4ubKsRfnS
kz8/b1hsF1EjLH+yTqvOyGXmUlzInfs9Hthvri62TtbITmnENLYDONA/UtCI
A7V086O3M3wXD/Jug87XwS7UCbbjFkMoOR4pmgrCKtYa5AaD0MbEcGC3ZwOY
XntxiXD684YlDPRtNNYJT96CrwVW33g72GbHojV/RXqF8L1VYU6DCmfjFOai
BSMUUVYXhtqObWLbxkgaIE+XZnzl9WrCTmsmhdeFA4TgNogC2RBClv8gqjCp
rc8K4N72ydvA/TT3vXi4dqdTrThtcBH09K/9cOW7FzfYdVpJ/YH0ol4/xWTS
bVIBoHaS8wpEVmRupvBUONiLHJboEWHMzz0rpVIh9K3XDhxrMuufosbEDqEl
sSy2E5vKJPHtGt59k1Bt1JE2hp04WTkVW61oaeNIe9cS9vgQpyGE95VgkNBy
mmaPlG9d/kZ1zWorNaebOxzzLy+EX+tUR61Qni71rAltVWCK+JBKcKVz5Y/l
3Zyi5hAw103BuNphoWJZPrNE47N4AWcy0r1HicV3G2HrLAKyxflsdQ+DBnie
hk72iV8GeK5ZmyGH8xK7pztaH+zSsHTVC7+pvurL9BUxH3U8EIATMlsiMAI9
rLBoVA7T9eFVt8V9FMNilMJs2DgRwvJWHdHMxeKYuz37KKZX2GKxCsPV0ANT
QFWm6PDlv0arzEypnUwCjs50sLmwLK5Frxs3RzAPBsul4HlC0rZtZ9KCG5zT
wxH1bq0LzeYKrm7k4e0RZL6Rjl4uylrFcxyubZO95Dy74ohi92xhac6J7t5J
hnMyOR7502FU9StkrsuK88OFhWnO0Coii/s/DiMFbfYUwNBo+zE2vJpmx+A3
P/y9W05RP95tbKvg5FYGBx6jASsp3H/DSTRYeQTZf9GxnPtdhE1bRsdhhjCD
r4ir0jsiJXicgaj4vftPVnbNRJEDU60+9N70HbG7QCna1MH59oVDEI06kIi1
Mo5AURc3wRf3S3ESer8lqTL18MpOZ95qssF0gjykyhxUD1vcvTKuUlp7PgTN
vc4vvTCdn3SGzz44MFNtLTUvVrHEY0tOQQp+0V9VzFasbJK1JlGSFCnVsFjc
elNT6IA7j9Rme/QG09F286DKHB6AJxR5i29aAJQlweTPVomKtGyIzBg9tlsf
mgei7MlwmxBefS5lBJdlqmzml2ql+wABcPSo387jaYqvuZ6IHj/KRO5p/RkD
mIamehxAGVV2lYn0yREWJ85tVkaCB5ufDbPAUcTsU0t7ZpSCftq7pFSZ79Hd
T7aulNtWi4Fj7khKavJpSoB6FgPju9oiBC9ywjsS9ZuLFPvLFoBv3ca8/XtP
Om4DSfuhRHqD6vop9GSRLuWwSZQVE12TMJV0zD5kGNLmPGclalEPee/MCrzU
OKZpeYuVu6qMESszT70D441xawWqu27+djGldzLJtF4T1Mcwoa1+vZ51qwE3
uTPeD4uYVyt91nxv01sui/RyGhHIY5GbjRefXkSs0ggT1udqZBFRxYFnHFUo
hqgJoyhcA1N3KfoUBHQ4Qo7dE+e4R7qWcguv+9RHzJPgyyIcp3vGn4HsPo4J
xntXeNVm86bos7JlZiZOLeGppuWf6DhrxfQ5q3akGsurP0JPAbOvX5b7jLAz
bx9O7YgTNVMKDzSLHOo1nPT5Ml6hXyDKe8KTWW+9ib/rb1j2IBtmd9quD1we
MxqnZvpcMPkRF5Uf5dpU9AXmKPTm4btfUfG8s5bgDM/fkQMJfZRJ3RdCd4+n
VINmxXb1O5nrSX7ynuSTW+E8gu6zQKyaCmnQ9Xp+GoN4uujZPb79meZNsMQm
oVeCsxTAOC2TBH7PQj0NPq77csJ3bAwrt41kSo5KerfDv/BYNs4iLaqeTaRz
yEMGKFh45rXyJG3kFe258EA7RJv9qeNQnIG/S7qdoFNUrTJ8djBPSrrYl4GG
S+vy6ZDRipM3/hSdH0Cx/G+S74tiGehRG10FizG4IL3hCEJQ30WIxQFRngDl
iLDiYfSEVSZVLjWDk0Gov8ZptVnsMlJ6jYmVebStFQwcxgmc/Ffp1iKOl0WF
AaT7NZxnxlvZfx0TjUsFbpdxKyWoDLkw6V1kXsN0+z6yXkKGY5F7mgT4f+mS
dVxrKB95r5Vhg17x87Dp3JXUzi/xm4STwKiyjvtqvOLfPJ696dLSI1ReVuGn
D6qnbFXGF0V0GzMhq+EdaBzRLKuH21RSB++F3CkMwnoFgA0mTLP5OBhW4/ao
fuZgMOSAGkvjStJiYHaLYXt+xT77+PTBV1HJnLlztSlQYDvHa/2gRi11FS3C
HdlIdMZurgPEmXj91hu8RGYR3MZ5oIFLsMKZY5F0YrYeqr83hUKevu9bqOSp
WHRKKRa+db6BiWAfjpwkiWep89ujjxQTCFQNbWp0He0QKu1kyRoMPmvDMW+o
FinBhNOT5d2zsB4DHmnf/o472zPajbXTf1lm17Io3+AQQRBmxfYTVGwBqMNW
eUe1F2aRS+9eM5d+jKQ9arCk5CIpMFtVS6vZwY1CxwQQO6hkSqx5PIY+kipa
qOdusrDAacHg4ERE8FSxslpY2SD8yzOz0lr/MvpifAhJmx5BJ1YMrhdBWtKj
2j/nKcnu9hBMSLwl4rfIFa6NYTgSPGtd/rqp3LBCBqW+GM5B12lXUKNqNTPL
zNg+Sd5EngMfuXM3QfGv/2gEJ5exSEWduw4yRlSwLY5Yf0P7S6/fXwKrX2be
sKPCcuDvA10DGZhr7zeGMexs1jrE6QiXJxohn3JbWy2zIwj75WVqOS1kvurz
CekmYyFGBzbLZyf8xeXLVCvGsld8DMFKeQDhk6fIhpP/F57+yliFmzQwMy1g
Ui+I+4KrcfkEPRJ/kiesCzz5NnNp6X9rJjjpaOypl+wlifkPNpmnDbAba7J+
MaW1Dw2YLLej4/r6pLDvrAO6bDZHpYnNV3fYFHnDZLr/o2SWxpO6ca4dluJl
PjcG3hWOoQ8oCwAQdCpGLW64ECAGS20ytaB41tLulOPANcaRQQQZ8u8SUW+I
fw5/ss5psA30QZeopFUuC1QSETbcLhve6l5WiOZdrWizVUQ8rtrdtmyGOrke
jhRAlYYaDUAgrkmh/ONAtC6SVJYYmSOR0NFesM4d6ajMcVv4JWQWHS7txfkM
b6GvlE+Yk1yo+SQUGdOyNQBi1gAKgjXh5NdfdsM0VgDmtJnkyDapI93RxBOo
xQ4ifgtCUoYh0iCC288N2bSN4ljLEzayuMEHf/Cn4QTKBEHwrHMDvQZEnHzH
72434n4Fsm2NHXYEyjwRnqg/SBZxu2BIkYQGFCF64IkMic5pl/lx71irHXuJ
h9k5HxQgl94WlnCHqq9VXZjolnRbaj4FvvM0anTbkqt3ReMRJm1HQOBH/KeD
jSf/4JjeqUo54Ll5P1VvzE7xOOuxXYkBeyuTe2yPE9sAu7XZBQZOH/lw8Lbx
8uskqpefhMvOB5dsTgErXy1Nf9s+AWdTj466fL71IT04S5w9qDl4/ks5bKkD
zJ91yofON2WAa8WhbjsAgGFVSq/aCbmdU1fK9TU8yONHlSB0m3qVi1iL3ImO
uQTDHK1vlfpUetKGG8a1d9cLZh3cJOLA7CtjSUGiGhHViK/3fAnB1Wu6hw8p
hE9vuSZxkNrZH+mD5dRolaShoW3JflQzhzOv23eVa3Cq/mdZAHCi/++Qt+VA
yDbXrnA7BHCeOu7Wg/cTWaUuncGJ9x9fNuKZ6Gcf05AOnMJ7bHxQyiqdnlti
EWvnPMzsi5AC6tCH8c/1eTMTAyHlGCahPAWp7p3IEtej2WxHebZae7zCiPhZ
mbPasEVLDAZ42jo4x4jAcsfYOy95tagGswa1dzspzyqLI5BYN9Mpl8Ly9XxY
AAvJKlzCuqwbF+kU3nJ/2+CCRqq+P3Fs8wkAHmCpJqfHsjF0YEOwVowMEKLp
m7wIsAojSlR5cC7eP1HNGPUeql+OJMoM7zZGjE8p6iyPqsORWrKq+vM3LUtL
wcRBSlzvHd+qQHpgZPUI/uE0ysdZY8/DJygxohgNiLPCNc7/8YPb1+ozDonT
vrzx3qp9e8H6duhhBCJVIuPiXFQFraYmK1h6WAMExGdxoi1RbznwE0HF8I0u
2IajDU+rA6b/AE1d8YhX8AOoQ9WI6NFwkODOp1m4+L5aKTTrkqtR9pK2ZeAR
WNI6MEDQF99pce0pQDEm31roJDufmj4j+SGfKoMIy5UsQQ/yryRuKTRCnkJ6
DSylYS8M4yJDLB6lasXGOJhucFUBPnIOk4Jf/5Y8sM4jd6wvJ1BxVLPr/eR2
s1fZiHrR5sWMNSJXbiFpq6WipUPaEcAgXW9hQkD2q3jUu8Omtst8gAZm+3dM
CLU5sm0CfGLM4MNoCgJw/718JaA3nF0dzUA/EG47E8VX7srXISNInyt+tzCB
/29UKKTYpCsDCIuAov8QJZM5KQsEoxkr/Q4pO7bRKDtaqrT6r6oTFu9Rjwo/
9IQXSKyBoZwCsH0vnSEH7c9tVP/sayfvW8BylNdtE08dM/TXUBS7QX8iA5s5
8ubFHFe26kWFM0/+CoBLDHWZuxUGClwaa0jJXmSD83QdC5tiHkJl2cmhxByF
bs9xAVC7kaHUiXTQ02Q/cZI/OmVU8KP4ikJvt0x+oOUJCBtHJLYTzHa104M/
oX5Y+dR+HH7wfhh2PPm3KBSehB+yIN2MVsjH3x2pb4E4vk+xpeRnjV+bhFEv
6jRrJX2rBEq0P0cDkyj5wZcTNRhOMAcwPDI2fPvutD5WOUC8VuM1W8O1JNDr
DnPqrLLdIU5UdAQp70SL5biX9JJ6rCDoVlxv541opJFaH5aOhLXtHLfpZKqz
l3WX4oZkTMbp2mLdhjvcLrFz7+LZ2nUB3ssiuG9FrNwt720C/LqKAlZV3nkj
lRRO31Qb54iPjE56/O8sj48YPgITZ2q/ZkiVKcqJC82jIotHg0hW6GKcxTKs
8OOgZQDhHsm8NEtaPz9NaLjJIE0ASfSBwRQK41CQGygUadvB0iAh2ig8v4Ou
nJ33zeNz6/Ce0HuD6nLocpP47vUP2YrSUiC/XAqzMmKR6g8nt/ZE4gr5/6Db
xy1OPvosgi9B395sXcOCJpluAEamjIyNzFH5OlGq1uPUXZpmS4bkWz/P77RA
FVsMpTxEialIamhWPCmnCNseIwPtf5u9kICmOPQxXSi9a+qsayz+nk86vKEB
JVf2QxAawApNjJuHKcZ+4tJnyK6FFJ5xPH6zgW66qO93Zp2l3g1milNCHci4
jk5Xk1MNSAQcnBvnDL0Jc4s+JvWwE9uyhJ3JVxpU98fj7nJRySe0jTl9J5lC
xyOWjRUQQU3zAJMz/8UW7jUB3PN0h7l/lMiI/8/xkdeUvDiIOp9OIHRA/P2T
o6nzJDmZJL6wEN5s0ZDpouW7pG0eOWobf9Hy3jcd5NYq1Bzux5OAi2/HCxKT
Qg1eCGuGyefNe2J/L92slvrAhmr88JUnk87TSjWRaaTMbdbf9SC+3StxQYWY
aYFGIyEkAh/OkTcqMnvGbMPyqjuB2BxnhwPzUPenDzEL7f0ltdusKte+0o+h
41mfD/SYmNpQSTJqV2Icb/2neVBOFLjLhDYg/NenFcmPXXnp1QlyMD9V8saW
UdFHuF8LM1B4lJkEmzGlnpp4lu8dIzrCci8gBrJ8cTnXZhFfCL2B9Y7Mg9AS
0+MLZ9uDezFQgyWNNlAOgCzyHaS6wkJVa7Sty9KhxqkXP8dhPkn2MlVyXFzF
SaXijJtXmixdvBxZEhZO4K829As3EEp1yc/mde8TDtpFPQOe1EdBdWhwrBdu
VxyGtry9MEPJaS+vyxQpjLioOCv/Ic5mp9cDJAPmCfj057bsanZ1s09MmXqs
jdhY5CYbHaRbC4nNnY1aVFHKWtmo+t04X11SPpxiOMMQv7su9loyYg8F/Zf5
bmXwsz4ewQnPYrVAdSYVK7Kx68BpcUIdJP5JXQDOkacuC7Bs4XgcjMF0FCmy
CT+oXpq3k/AZNnkofzdMVm4lUiBJCwHcXJeBIF5AmaORVaHuF7OaV0pybyWU
hgmEUomAw6do2HzMmHDnEhCdOoJbNX1d5rU4xHnmDt2B8YsnIx5oi3VcU48z
NP9xHlz/2YXOM4NvNaZfkaOnrjOJLb50Kd8exQCsn4RQCjYVVnnb/KvvYYZm
RSYUW+xvSNJTEmDqjSjM++g/iuC6JEB/bcPro9nbQBOFIzn5BtDyqSMq9jJE
Mjq9WnBkwgBHQ7wOChZKhySX7J2PGl8y0eOlahEF6RZ0sOdHEirAi7vc04su
aLj4fb6fbJ1hObNQXmEXtM67YxymLI5kG1JF8zioEIc/+5w6qQGn5mWxr5eV
EYrJekzr8NfeSyKxWd0eKwfLbhwA84EL341HeeIptHIf6sixNHeueSC6jD8J
Vf4Sqji+WXBkVlyVaCBzNgUf/cOtJvkPXM7ujRh/7DhmznibEmWb9GA/pg2s
SC2X5OkjJgHQ5GYnX/7xjijblvYU4SohkseCfU8PKFQPEIm81ySpTld9GGOB
hgV9KuDsB2S4eooR62LoW/ZVbFTl2EFV/HRXLnl9bevRpoV8be+kTH+9Y4h/
3uBNmvkX56a6K+V78mFdZAk3WaKIRdGjVMcqV+kFedTPoHrIScW2JtEY9ZBP
VL5iD3GSbI6kCtIh/LQEQ3a7FK+VlhdqD7gzFbBRhEXxpw4bYTccWN+zZ7kF
uvuzbopi7ElI+wC7gFvj85HgMOFIQU9e+e2UxgKFKly1WYlfHZUz7s+VrfEg
SynCE2nMRTVAdv4RrtnS5Uvh1vkv/uxn1MHetv0Nw+8ZW/qalEJaLgymOwGs
HPzFfYHxfwjoKKtaLSSzP0BdbE7Nu0l6aO06tKSLbJox7rWUIgwPHHdamORt
byG1Bpxs9mVjSxgwkyiu9wSl4DGqntO+0oIN8IF+WG6oQZW7+H5y/WFCX0Du
Juy9yPSvWNWC3h62LHsuwUucfAD0ndEVv+xyxGV6eVxgds8xVWplB43FcOxd
BhBgsRyVEnkt7dp/uGtYnEUTHcruHF0xz4ybB0tLu6K8AcxytapqsT8xHRlS
qjvLtX3K1t8uMco0xpdIQVnmj15cz7zxZn+oW7WagnpXBFBkq8+Q73ZZIR8V
6OQsYwIeJri2SjZd6s4n2RfegcVk/Pt9rGndkVNPOc4HkVmh5Fbte5CTgN77
7bolEf3BjNRtzJ0UZqKeesQl3cgc+eiFJJuj9kQLAnIW+BtAUVKqvpSoKugU
TYRgi1uGD6jtQNYXGaX0zG1kx4LUsZWm21Lr/d0nrN8ddA++OIfVvchqE8R9
WZsQL4u/eVFE4NZsTHVV/Xi5+Z9HUTcQrqbORiWy1XNry4WL7ep4mja6bJ1N
CB4DLxi35MF9v/L8yu3c39JJoHSkypzyjbQqZ2ffRl1i3AzuGM53bRCc204N
fvpmcHCvHs42H+A6BobWYKu4eM3qGLGPtl7n46SyPHtoYB5P4dUusESk+RKI
02wbKnaXwMD69wBh0Eot050ye7Lo9QTHjZoObm7nxBLgqXfLrw21PMQamskv
D+xVsWsRMYhAViasWiT1+GeCE7jRcM6YmZTM3Nxos+cTViiMlqGp3FynUBHj
kph+EIvRAY959q/uraPCitLCLTIHcdv+szu+Na5FkDo7MlDs8v7tQ9Dwd2ND
2JvrHPs5PCAJDwRlrbT2EeGSTGXyWKehluuaqv+fs7e86k4ZdySmtF8nJpjk
P0kGo0OfF3HOgySEJwEr3SlOq8cOWaEE7W3aqgXUcxhqjk1fSV/he7qZAe/d
dv91l5lVm5FDvJUbl1jd49ngBTMVOEbJCajc+9CzkZDsff8VjdXMhrqu4Vwq
tFdEN8eYvI85X22c11w7d86TuQmHrFjLexo4BdPzH118BfoXAtzXRI3XOPJS
lostQgBBrGK+Z+N+rQ+O8KLrzCV8AjcmOpePG/68J/5HrX3AdgCKRzoDeAqO
SW99rNm0+cck9O9W/1BDzC3anjdptx4TSojCfZfdLRO3uIQhRJdHXY+7Bu93
cPO5JilkfrdRycs6b2SsRlT62TGUNJOZzC3/D5hwVIiIUhcTBncoNytC/GIK
7VPxXcTBi2GORtDdK55gibfM7li7FVDAhXBhEqjpx9bzdotM104Ntl6gCX3E
NLVsEtprnx35pd1O0jpr9I1sNgarv6qy7+M1QjdqAkYC/RB2dd1I9U58Olqo
7qQiMBMOdA0212HJKLtykjdraKy65kAbyKE4bpUE1AWVoxg0ayTu0vPGyQOV
HY+1LvEsTZ8pJ9+PU9phaHNWmStDan91mX91dPULti5t3Z2K5jGc0Ks9vSme
TVwzpbuFJsCGpjZq3kRu9mjlvMkJNA8zt6yFCNc9nVIdPcc2WZXHs/53jiAP
xrdW5aOoS/oOyZix+0m4PezpQ8lEXZ+Khe0y4CLUTzo8y3qsqnxdrqlNtClD
7fLy1gMIvp2R5B8Rw9nXQX6D1NqPv1nprCqo+xsUBaCivRadJFjwuW8PQE0X
UPQQgc5p+UogwA0LI/YYSAGiCR6lSSG0k3kmO0Z6OoPGcMgZQg4Ni7YZwQXo
CyPaK0CKbLrgY7JT1GqAqDwe99DM1SzWFzoX4zi+8stzXxauVnXaP2Cmm0Ye
UcrEjwXFH+ltwT4BVr8Xl8pz2sqyrvBCRcoVlsUSxvQKlZptfmAS8F/VEo5t
V1vMxEy344Iu/XV3mAayKJBhejFu3z2llXIh/7etxlQqJCa24ONj1TXLgAtC
rGBNT2++tKybdr5K2du0R70SyQOhZAkCPwczejr3TzcIDGtrPQWjGkUNeP7A
VQFV7K049zjr1UzHEf58RSRa37+fL7wxX17e3gOD2e1YDZcTv3JfH6Ypdl7S
JzuoWlwmnMIjgqgnSZanze0uqySZIVHvWOEH+N7oZNIL1echV8ZJvNXFVKtV
//ldqpDxYIoi6vGXawCoHG1nrT3yxVSusMs+SgqVmo4mJ6BpuoVuPzazKLkB
lgbWS0tQsn4EMwpXZRBSfP+B3X8Ny5UKcHm0HgUV5HHUZzeA2cj8TmqfEedV
VBV7z0CVyf7y/71dSAUM/e6Da0C2uImVVBV7Y6i2CT3F3rSdo+6VX8zFjMsT
1IqR8FKBcrjuGpM3xLQn9oM7z402kPKquvieNP5iZDgQHo8/PYbezkTCLus7
rQVmKx+/eSBNWOs1/nIn+h5rcmnLR1iiJJw+SYw3ww2NIf60YIMsbp9q9eU/
ZO1/emZRPUjzJtNxoJxLIyYY7Cd8jG7OqYFxZ7dXPA4FIGb2BwUDATQdGHeu
ThWKQHqFd72kpEOq6rNeQa+I+R2goB5guQCQGSPruJhjeqUlMSC8q4DAmtab
E9Oo0MCcAhqQd0O1Orj+ZH/iUXEysfuQ903rdtTVkeCN27fnoKWSpsdQXnbr
bwvLQkemXiXOl8STBQopImayjVfgVw9J/bIHO1+VRE+daKLgO9wSZCfXJJ+d
8Y38WVBtVu/6RrARen7uwq1F595T0BiQMDxz1HgiOP7ONTaJ9pRPZKDECHbo
3iRRRDJ6iezRoB86TzTdm+qYkFxahgN0qJ2bx0yrM79eyZ66MIdREGbRDaR8
c6RwsHxp8FjWSNtGPwPLuV5njWhBIYWbILm1TVTbLycJ8CGCeoPrqB0UVQMg
ktGs6Mf1YcVCJPYwvWKVEBISkfWn596TNSEDOFx1bCJdqW6Q32CQwEj8hIow
hIg6kKCafAUEqUR6419UL+CYgf0+JIHw38zBApHkOqEqIs/stYclBfVrMGkr
qOWWjcxRMFnrWmz/v6TjhZWV3dkH5E72zYWMWLCEY1ia0lSmUgnrPZQYKe6b
IU16OYtexHQhkGX8jxVt2ivBYJIUw2ayQcSgnCvId+LMHZKrvnwqawirZd9I
gBD84BeDJaKO+T4gygmkS9mkyzjW1FLOQKUeE2YwnBhxw7w76k5FO+4ilw7r
D1mJrKOw4xlIN4zhtlOXhlAJeedCCYWCe8EZlKly98qdkAtVBkUcEGeh7Zmn
RKH0l+dTBGoeeZnuRl9DnMETyGlB9fTVqPOSWj+X5lNYmaL4rotjQbjfF/wT
IVaIziXh7pjihtBwwRDhWo3tnHnKgpDUpXGPhzbvBjxvqt5o29NN9yZmytDl
BRzEfVreVP++vKmuAuaqAWfLfF2pQr8yMDXMAtHiFBENNLcWrS3wRRPC+Niw
3pHiKSJkys94ROfUognjWPC6XRH/Uvpkhec+kktj8Mlk8D/HYkpVx5VhmYiu
bpBx0K7J3Xb7hoE7yrlUPqcd1CCnEyU7eggIvhfnUIISxCCOdjDr6hxJ6jHK
wz34HZzG0EJ+rNAmuZkQFx+xxlqR6QzQYX3zssAK8g5zTsFfUTP+od14Wx5K
uyEZW+st5FGi4kxWqzX8v8rxppc3U+YuI6LrPPjhBvZZYcPDJCaiqN6w4aLP
hMIcRJSbOmTlcvAqKWBmDVZFlb7NrnSMUJ7xklvcA844Xqz1p5LBZPEFVr+W
2qJm1djw8BCPHTQ/jGMWsv4qL3Hz7QN8aCXS5EUAgG2CUaJshStnz5y2umqJ
yOOIawcIP+czv9AeaiEXsmeWPF7SVBKjy6G26RWx8tZ6uF+Qw/RmXSPpauaV
vz8GCtgEmzcSR2RH7rXMJlvy0f7Yw7Gva4ZsYX6BTZ1MyG8ZSrrghgLyYfI9
q1mVvOqsIvVKb3okQ2PYSO4yzD7RRW8EgQkITt8C37Bup1M96AqZCNZVjCq+
dMxFCGlQbW4orVDR+A13ZefiLB/9zM38m1fodumpHAOlF1zlKu7CE3nfELq1
gIqSGvdkatXHB/9gNoL+WggjEwFLjgX6gxHrQ0uM+e07AzniKL0ZwOKfFDGi
w+R0PXdN6uc9WZnQ22i2UpVW9lBeyUUUCvpmAJ50QZjoX1yZrP1uAra/7yzd
Ow6LP6ZUbPuxUrB6rQ+vOvcy6u0vUP85TS5SVkMwqUgyb1qVORoegIBpR/HU
PthnLBzv5WysxKfODjWrAoswnyWKoayzkp8AhaYzKo2t5dsJyCDkvgvV4fuz
TnNmD4e/pimLOeJ9zxXTaYrzUgh09Gyc1P8lo+PCoHL4zRSQjDr1SaP51drA
RmZZpwdh34t0BhAyeS9HP0Toun8ak/02E0w+/mI56e93cS6klBe8+2L6E4dZ
25tjES8+AAQ+6dhcD0+7RyVpqhTiymUsNXSRMf5DdkLYqwFQbPn7QJvGkTFp
SRHmnX/6EAflCNxGwESJYDU1sRn3e67GJ9UPuPpFC7AD75Nszla+/hqMy0ew
UuNS87TooKNQpZGtbI/78L/evOwwFpwLITwXkjrKQyF8A6yHug+/FI9XtB2B
66ynxk3tQf4+l6/5DNRzv7EandvKQdhzeCane4QbVXpzKD+/9NPP1uFShoso
pb5a7vMym5uObBkPF0afDo73Ad/7/WASyLXNNQUpU4kLrDEkV4x1TjZqyooz
u0cv6eSvjhknk2IY1+xoeRvqSNJF4UA6B1dV1gmO6inJ2CterUM2YgmDKkye
LMHK4xbgX4/MfAzlA30RWl66+OCV+TaVTM8gQoHTxmpq6BnkfbhRunGaoawv
HvvB3j8jCt4+syCadY/MWZsfgFX9tyx6YPs0ixtMqisWLkBS/Swor08clPQT
qH6om/JGDwXfN8K7Bcs5xDaQ67arhLCWyIq9Bhqm3/jVIQbkN2pBCZ1zNoBj
TAskONWB5GGJbLd9a45jfMq77nZZxA9Cjd5XVaofpML/U+tB8WUZ0tRxi6bq
rBxrFSJBLeiKwLSAk7apceiAf7SqIC2UHiPP7CL/TFWmxzv/lu85z9k8rh+E
Gqkyb8Td5VV005sNE2pVz/MY65oobSr2T7SEad6pFb6rITR+GiSD3ppHMNNi
4NBrHu36M/6Gnp6fn18+rq99zHbn6C6z/674QiZ/OrCI/iV6Jpyc+0P+M0DS
2iH77uy6erOJG+rmOwAFket9kdeHFaZo+oIsFG2jqtvGqaNq+ppfNaxuM3QR
CH7Ps+zupc31rT2NDl0bVUUYQpb+HanTNSq27OlFhsFdMZ0RqSoWlhlrtcyk
fPY3VPeOp2qQ78+rJa5Uv9SzQnGx5qEU8yIyuszxVrFikkU7aq+IF5BOc8vA
zp661dsYlEQ8H85PPG5THaWCxMoDR//96Y9GaeQsJooqobvW/UU5Su6V1IT5
OSFSIAMCUmuRLLuSOCHoR517GiuJSFfCuJeeg2L/Hn7dWvZcPXEe/L1Ted7b
ZdurJ70otlZjnhgWkQlULkPDtUUC1WweTwMvFO1kS28nk91kbg+TSo/1sZRD
dDE2gKZvv142n0HyXg2GVaPqoqdSM+rm8fYJ9E91O24w/RUIdYbBrkK3pfPz
DTld/J2tnE5CxdEZA4qlM5fCjac9flbITg8NwTJcc3otzfLIGGmpV/sYI0xc
nrcIVYGpq76JZCuNVpMAzli7XllhYGG9PB7ifHCx8tEIY3tcdT6mlhsUTG/K
4/roH5vcmliKuyMXmeHd7jU+0Zp8/Z5/TvtqCQ+iINd5BQEhVU1aNj2Imf+M
6rMQMKX14pWW8rthV3R/EBUzXVVL3fIYl0Xy4/QtnNjRYyy051Rb9rhLmEp+
bgg97ZPoQxBOF07sl+GdMi2fbEqP4mfFGqvJtdQqnr3Jw1XAk+0aiWPB/8ps
lkHL/sLuLO9lOYTEHzPyJAezuK9W2nnN4bjHTH7nF8t9OGcY356jlJZE1Nx9
WFIbCZezl5c97NTCoBYRYECtEfIHOBQ98z82yKPImPPI7XEr3lQfDioBrxPP
DLuJyc6HlPzau0nXt8KOm9z5wUGPBOsYzi+hcBb0cnyb+u8LUY08ISUp40od
ntisy9EwfECAOteMkcFjLkHaPnkl0j0ENMe07zxYpnYlXmdcOPCatkCFJWr7
3eLBf0Wi0Nhg3rVkOYXoE0flcIuA8BfMhG5nI0v5wMVHt9oCynq0sJ9KXR/2
Bb9JpPe8ET+ncAzANWjUENvFygNfW5pxGrwHTS1ksmCLaTjJeeyHCVgTZPr5
tP97QiiJEnj9S/AObU3aUx+CI8VDW+WQ9AIWUdaRT4wOX9h6Ypk7Xb3cAOBX
wP2ev0PMh+Tm000FARoXqkg3ZLIWzXWvoYaewHOd9XLAnSg4n2Ge/SsCrvcn
0hN3ShoynHjBWEj3sajvxCbYuTfjXcQCYDuWiip5WTHTtki9tXDiyh4+0MjD
kFA34YBqGuKZUACox7PL8NWWHWz/WGZ8dGil48CjWLiYm4UZO3dBAsj/9O+V
0+vwIkogXYO/Hxrr/QTTtO4drnqItqWV+scyHb24q4ACvrMJjC9sIl3670eO
BC8GKlU/CWj/pCQl/a5JqtWVLGFqFpOIY3ViZZB/RO2Rrqk+JU/0+e5Hi6jo
qIkq+jRxXE4g98BXnw6dHArHejPF2t7ckLA9Y2G/Ol/jphnfGig8cIKVQMZ2
HTbyvZXwYoBajW7f7f2HbjF8wXbt4hpfOLTOgJ+ocE7W8URxNxcqQ3WfoweJ
jEFdqXlRZ81xcet/il9+b9Vgsbf025VcGuhbqu45JcQp6JsEwuEcbzJx4Fdv
us7rGbG2X4JZOPcEYsMOs1FBoAo6+DpaYqEH5ybv1DuE9NuXc6oU7zlLNnGl
pQaQX9VZTo1O+wMdzJKg0dNdcQA9G9L+KvptDjmKSI7VNYQYv43M4Jl5yyKs
RY8FbOutvtrcaAtx8X6qelm+oEnR99WGtrxox8A0p2UT2HHEpca7ILw/CUYz
ZA7MhiqLjA9Le7B2ZInCeDMTrp+H+K+Emz3+1CdUgmwVhC+YqTxHqiHlvl7U
jdyWlTvNkkCGZRB85CsPHy4H2bnm9kMi3+5bfWT3ykmmIV3rxKXtmTXvkbHA
nThWkHfk09vSXOVqj3ZTmyLDg73x8oSOJPNawFfgf59NsDOGrf240iwS9fcZ
of13el+qVQ7kuPF+2mnmlHy/tuO8g1z8GenvTrw57OttQQWlQflaBg5I7bT+
BjQe8mnTl0JOZkz8vHgjvwMw6TBFVwiRdI/E/aY0SORkWgsIrJRAfX0q1kZ0
82nh8KXbIZXa+Q8OSbP1dlx4teeR8gs5T/giiZEIIAGn8dDD2I4kW3cPBka8
DtboqjIbqBCD5AJCWYfn2Ysy/1aYlwoJpWWLQTrQ8jz938b85gyPySXN6MEl
sDI+UuYgREckZ0G8OTf9w00fHu6HxnGB7ZABJCX9fPxO6qWTVb8+6zvk9lNq
JpaK0tzKwy7qUfGnf8acEom9ipPSjEK6GjUAKpv6E77sohK6Ty2euFLESPhC
5NsTapsKAEIcNRQ/yDHM9HQBJ37tfJhWitGjOKjatf008+aGSfu+03Pjc1AL
PCs/fllTNT9fP8jrLj9InmstEPDboa3Mgd7JWR5Ls3xxLVTQQAYqpvYn5R2P
ph8WxQjwlA9QU6/59cxpa5lS1XHh+T2hU79JVIqmx+qdxT6atINjIiLp6TpP
LhEnvkYcApu4o3AsvHpNaNIG2xObBs5PhBPSD3prekb2d2JzphF0JUgWKOrp
IUqknJNd033y1NzlQdC69oxDyhQKS40XJfUFz1cBusZVMVr1m1C3DP6Bc2yK
rsjTkzGNkPmhgXgFB6BJdiQEhSI95q9NTDdwLXjpuQhZHiyEY2jhOFSp+jIv
wsEgqZbF2SruI21M+AlLdwhJmGGpr6CKJgwnAXcyZCOjImrkMnR+Hi+DcSBX
5yeaxoUSHmfF1MVjc63KcELINKhkLktqllE0NiOUaRCaQLgRJI70AI/0gE+y
camP2D9gj5fyORcM3HDBNuEaU7mrrI24FOhGxtAtHPP8bcF4dduminWU8MG7
JdXcV7JO1RqBwCioVKjsuwKaKndYeUe/+8NSJrAV7vPVVwtVC3gcU9nKUREn
ImV34yXxEDXZT02A4EuPZlJQnZXPKQ9D46DHfjobzxlu1r+VQGjRWnN7LPNi
WG4mgBfRrQ6Ox5uZ9WGmUcuD30XVk6x4GgR9kzmo1t7T3qvBSQUbDFaH7vJm
vFdPQ3I9P34wO++ORlrEY5cBiyMi+R3J9zfaU8AM8es69qywYNbNGQxaDeng
+EYq7T3QoTHYC4WwbrVbMcil06KHlVhYDKoavuCgzSKGwEmQGN5p4qFH44Ab
9DBoObKysFFAkIGGKkdkBa1Nmed70UUOb1t/nKIYbFOeWTgr80bjpr5jo/rg
Oxe/H9gohYa3E21lOlptk8BddRxfvZSddtJ/WhuB5tux8xl7kLTR75KNcptV
o9v8HmZ90Kt5U/s1cEWWNKKGuJ0YP3OpQ/rL2hzyR9Nduz+MMQ8W2X9qS7xg
l2jCSXa2WTU1vkfMT33s2oJJBJ88H0hfYSjBAUfji1vRTeJeFdAzzuoYiiTN
Afr16N8G1QMDoOqv6WBitkYXaT+1QnaNWfSOyxKuViElki/5/tM5iAqW1tuE
FW7TniOSbshHHVv4UHLAP+pgqaVmg9eJHbIbWtmNHMJsSPjgKzFXhwR/dbvP
4f799trojnXdHHqsa0xb8vEYqyhnXbiocbEVoAgbVaBXmdSrWjzzYanCCEfr
wLggLG4fgQSPG8OScPnpVoaowJzBORATxxhZt3q+bdgDJbCu5yhXNhtoz33L
92JRs/3YwlOWQ4CU1+fVGk8VMqmsrr7YNuxczS4UpmuQxNP7YSnDrptVjbV/
AhAyPyO72rU6TGobZl5Z5t+kj+A0R4nG4Pk2E0x7WHODQGpZq9d538LL2uyz
ggr8WopUBP9XFsVDiW6DhiL/J7oSDooguj5BbFARdAJtP94JaQ28PHmtTrdn
0FsbbKBmA/dmnfBR/tHVj3GhCkkLipB2EI0PUdmNSlEvQIYIvgxIT/fjkWxc
KuQ7EVjFgdbhbydpaXCJ8kODB6IMr2ehZIRwjM+SuVV1ofU//QBlWcA1mc+w
F2WAKo3ZNENyWA9T9IZbsTmndo1+yJ8W8xxJnSVUjwmXf+UNE+rV2cEytC+6
Lms0v+twkdFHNsKa7fROEZmEMHcNxtqBYr4TqM13+rCIyZeMYDW7n10eRV4W
DWEr6gn1tJG7/W082vUeclzu8Ady30kzjg5xvlrXW6HWerE+Bi9a3FnjFA7C
EoJmxo3NbiWcd/QhpsKg8B/kX5ykZyREE0KxhtHg8F9TGjwRcw4RQvDmghCO
F1J5qWdWnq3pS4bFRUzviLC2OYYTHUYT3rWtdRD6NCAZtzrTT+zAS2fa+qZD
WPlkQgM9jDJsMftm12rKEjQ6q/Un+Epe6wjfRFHZhJsxo3NbF1wuxXF7zzTv
cqN07xvKW667c8w4dQzWRiS3x8qDViCc/DypGVp+ly+4MzEQfUnicPGvuruV
9iubkZc9STv/GQrMhpcaVuDaJPK2N0WJ9GrsTvJQdNN3D4hOJmB2un0AGuql
zsRRgqLek/R+fRZPv4tX81cFLIg4Xq4urSOxlgpJNEAbKUTcSXcQiZ+6yKHp
TRuevaZkabA2jG+iHjCbeFBScR5DtRtHHKJwUr1+zQ+Unvt9x5/TKY7lcIoE
9tHR8wsiuBAy/LU++1klDaS5s5Vws/FaBgBaMzBtHIzlUT5Qm0IOizcfS0LF
R4VTdmgU0bDvT6VKohQlScgdadACvix+qSDkjmfYLFhOFtRnmMMIp7yO6wZM
XnoUGNZeKUWZMBQJercg5Etgx51KfPZYMMxhwqBX6hAjexLN0rlYiGoy81A4
gz5uoIwr5rEQjvzQTwwl/fUlgo8REpq7fF8zNnstNry5Y354yhq5t6YuXii+
F+yIa4k62fsdbAvdZxPohpDx7f/mG2u9Q2sydd2TFWOndRc/mU0yMv3PgTiB
y6/QOwKmfAzhruNcuMRWdyHwtYG8IN05aS8MbSs+XZFCHgLtA1aQFdcrncYj
Lb5ipr0fAEzQGSvfFoWX+KAJ1Dq87vhBB/7+TcRjEgvpGAbhiuyfPPsTcmbZ
lmfbz53WdY9+tsqfCfU1LdKNBJKKKQknKRqWLrVBCppJFUuXsxGkUvUWKpca
CJ17uIGJVe12USkxie6k3bPoDs87b79JOpJVf1Td6zKB1NFwp0qjpccvne5t
7U/gxw7uLSo3kNcvXo3h47s4MvNQNbnVijVNYIjj0JjNqsg//DVxeF0DX2wW
8mTiHmJjXxIs9UHT23MNvC0DCimN4yQMCc76Bbq4k7naS27ZxWswyus80K8W
E4Wpup9DLyJ2D2zHKaNbRznZ75FVHIht0tQ5yTUum+giFs+JBIq5RQH1uPIQ
F1/k8UDoz+6pYQNBEIlIymbrKR6OolZdNLmiUrvi8UXYJeKjmFbWbjSq5wBy
jv1ciNObffH30Qh1kVUhcIyWwx6hAgXKsoR5OAOmR6v30CEnEOEZGUubfhKP
C5/LTLNz5YWnGF1GoDMU2IgwWs8gGHyxe+7WN0B2P/bGzZGR5RSaX23v0xBI
Zdllicwp/lEqO2VO7SB5DuBugoAYjxHCI5fOTGWiYyFK+Jhg+yCii4FO348Z
XlJ0r2DSBxv8zGhcgHeKXwdnrGUekcEtaKJl7xQa76HgJs56534WUI0uc9gQ
SI5LTvwwztBNMYnfE0RoDHawP8fjYP0RXjSJEZGHmxtjoTIr4KXYDcnhVnmc
fIaSodokhi5Law/3TiGGSu3JjlkvETvHJI3lElFGTcLUI/9tJpNNtBkoQnHk
NAkr8fnrVjnLTmTvIbAl1p+tU86EO+QUAJ4v67JNcTFbWgmhy2NnyR9BgFQs
XoJW18gDxmyrrgvY7iRyuUAelhJtE7FA58FOzzADcpio8VCfx1+ZOPXqYPHP
5Ak1FGWLep4CqD3z6MSNTeYAkVMcA1ZwsIaktuOSET/ar9OTpk9r8MO2eCed
YX9D0OnIHlLcOjB42WNS8fRsJrSyAQm7Z5iIvi+ehZBl3z0r4lRcT6d3t9gT
itxvI6VRebH0+CoV5jA3XEm+C/lAlxCyANHLXeXgCediYkmZjWijCWAi1IG5
MaPTS46C4TtznIjDFaSOrAsPDjwqmlrFi1weTs4/ejIZP+uWRrhqPj+dTiGT
RJlJ9+vZYwHrW6ZbnVQ7ZrUnNryz49E0KisL9CLREAN9fA/0MzFlLiCSKG/2
mGracdJN5RRezMIzhtuUyJKwe9V+kNi9aphaayo3AlgmYch4+Oy2jQ/zCVKe
JYgSc/hOV3C5MnwfjncGoRuqqVyo7/8fRv8tSeGM/t8yKqy7Cetmx0aud+ug
nlBUX08yqSUfWLUluXfu9o4ApsVP/oLmcpc8aD63YsCs3vXXv/a3h42yXH8T
GQbfG7Xu15wJ2dEhDwUPs0OVPeB+lMvvEgLdq+2QoH5ViR4WDr+Ea49pgkeu
6OJA7a44JaDSnz0TlG+Qgk9K7C/2BxjcqPG4461UAFopxbG9JGs3lzKLbhyt
S+PII8FRkGVJTPvwkgKZQPzBhgQSDOJN+0GqaQ18zwWLoqoUITUAW6/kzbcP
7h5Duotfz5X54IljALxVM1v5t9SGQ+o0CDX2H6rzaqsgOBcyfs2meBKTAUtH
0G/kt3HV3eQ2WlVBziTjqmaBS/oFUvihdvhn2Meh9Q5yruQoGSip2dCEQtlN
2+d+khbpCTenWr1wQbfA7FL3xdV6jeGmCWvq37fYfRQf976OhYXxYtrox4I9
lb8TqH//TdgK87BKmwIgI2jmqrNJraoE6Ye4sxb7whLUzSR/YxJKtDtwG49Z
mljpKM27+mBkbK7uYLzJWgRbeeW+JKbEkSQ2omC2ZCz7Aee+NQVVljpO+EX0
oF4CJ9W87QDjHejAxyvkradaFyFoSjsMv6uGXdGBkTDFXi0P8M2Q72Ul3IfT
dAmtZyKEtc5BkZPL1TDUuUW+jKpxjt7oI2Xl5pVhN/FUsS4NE+fVuSvdw74J
JzXwsmQfiEiK9rKTDvhJ21RbImR8hAwi+NyVglx2vSIXKeKaBniCLIeibr7U
cPr/RotW8lfdUDnX11rDrGFlP+l0OA8ueVD1mboc80Cl3Njz8xq4KkRUsIRd
fQeI/U42BTEqD1HqK/GHS7XXwRuxq/8jeYrpQ228235GNuhvVK8VlM/6Tfrg
+0Svx1widntCv3fbX8j/O9EyGi5SeoCGJl3pO71en23Kzfk7WZf7JV1mCjcD
iOP5SWUF7tVY+0uJZRd01TFEbHVnI+11r9xwW/rlweXAJRXyPMOgTYmsWIRZ
st1vTxsPLrKuqNIYPn83536YAnP98wm+FswGUXN/ARNGXGXFa7yxhoWRhJqr
qJZK/t0DKzrBCauz2SCzCr4hilGsomuemirxBG6mJqqT34A3dTZnaJsOq6w/
letW/wUT4DdfIG/QNVMHOfnWDkbPX2A8Ur/MqL+LgIRg0BdHMfqHHSVSmizR
gYZt3CVtDHpHWMh7b5mazEp8DBOb8mEezf8QOOECbsHZME33ZJ6Og4DEC1iV
mFNjoXs5usGturoo/E3JbHLfhL/3ZNL2L0TJDh/lgfHA1zu1II3OBB0Os9e4
eowMae3gZBA5t1oT6HzdGejyb+MorokAVZIWU693XgPDFkYupkkFTMazHX3S
D0/EoqEO28F3xiK16NbLVk1SMWF4dc3ZhKW5IFt4qBRgaCARY0M+ptohWu9p
i6hR2ZiiQkkzjd8JmxPzPNxs7/4y3X8H+2IZqDP1s/4HjSFsFm/eD85u0sNX
xqg4mjZZKjb0Z970JwnNUFLptDTORAGm6FQ2tmiWDpdByAuHwVYh2mu7Qicc
UgQo5AE5Euxs/keqSH61K7dBlUfIkIJr1t4pMwM43OgxeQlETZszhxLhKV7j
Gd22zlFOhKgvSAt+oJxwi62hvpXeFpoFNia6LwDY62TaUJxZ2nLXg1oKOyE8
c6fpouqRs3AhSqoVkO1icQ19DF+g0qoht+qh+SvlNNBq3MxBykWDXax7zuWX
2jhuZSke4chA6T/dKwVF97rR6DV+kCtuaU5mCnQCwaIc9ilPKAgXhJMTcHRS
PBFr+6I6l3yW4LAo69g89666yaSmZ83vHGyPqAJcobV/7lwOcUOoDQFChj5m
jUa4r0PP+yYZNVPq1TVocDrihnVjDUGTny/YlTtyvJ48lOz1e6I2eZWi394g
F1BopTE++FEJWvK4B1JgBEGqQBw16CGQT281Ah9gaTNJYJs1ylYJXsVNWz3n
6MEwIuWGrQ+2LUzAu88eML6nf9nlcsy5vt0HiawZIeOPyn1e6xE/jojmdodd
sSGp90v2a0rnMK2UGgDwuM0jBMgFHrhtr5xxRn8m1A/6s5eqRAePI6lTOJVx
D+8nanUN1Qm40N+V2pKhK0qQIU5f0qbBbknVz6oPgzerlI1QpMlUiJQN4IlB
XJROcj9IbcWvXEjxuPrnQ9DkkQ6CLM7prSFd6qlyXxd0byz0Pol4WhhSV+kW
qfyGZNKPKFpvq/Pkx1a8zM2xtDYyeEuPMQWEnaPdAfHloFA4qY1hcy2JIyeE
/8y4GnJ7W3OG2owkBzNAeQGYLfQf1+rqn8tDpmOHikLU7oyfO3bPDU8lh54g
Als/hK+qvCpp7uOKsmZlHMbNxHW0WIMk2mn7tB/GKe1H2zm/pJM91M/Eoryc
7mp4E5+VVnIFxDAhiYFA1lYlxGOp0aXH9dV8FxPpsDkuZIlHj6FpgjbZRlUl
bZPhH6JmUsnd9Ap+9oJFwu1nGj+CyPQREDaP6Z4VnIjepLknA/NqmEM/AeYU
lhrSCWwF07+UvJ95D0qoU7lsvE/G98cBySW7NyjkDRUQ5WBBeE+B9E0Xd10i
ecixS5zoMBhSsNItCWbhYwdmhsE5dUZrVGqOhpC6OFGYZEgJBCtYVYwfBl2O
lfuUqrt6/t0edPqET08Y1ewndXa3VHR6oAYImbY/3qz4X+4Ubh63ZTR+4Wvp
sx+vPFgksajJ3wME/7WtSKgX9QBNVMeax23CM2a8aVWfsoMj+GZiDkfZMSC/
eemNnM0lUxPZCkrb96YJborZeIFmETX/1UMKHGFmS0FFH9cTLyxTF0/qtkEc
NWgMEmddonq66X5b+FjFz5RtBamHNq68ZWhKN7lX0WPav50fca+LbEyHCZFw
Ffkrd+tWsOh02g0LikXyDaPBXNoIBwbuPZ3DK3JkX5SpmZ+K5Aw8pk7ukLn9
FWxFpBaXcP+nPwSZa8rbcObw1Z9hhN0kXrPr1DuJi93loWfruQn0tZ3rLZV2
2WMRE6O1eHeQo1rAbQbG3xWGjwmw6PZGhw+5NBtXiFT6l5jUTWRaacASaoeg
SQj4kSNM+8X2D6rb48nLe1N3NF+nKNaHgPQeTSDP64bMvmMFf2HJNz1tuMWh
yidHaRjfTAiU3xjolO1MfOTJjlq9JB9Nrp9Q7+LyXPeG78/mBLrJkLWB2WkC
svk7xwwVs13tTgG2qYoPJmqFtZxsANy5Fl71mIe2oLJ7WgE/TEAqSdCP1bBy
ZYYICDcIawsAnOfimFEInKX2VVn6XhMzni135cuSL00Zcd+jjlYU/xdP3HD1
fcnv5gB9AJPxiB3k2dZXHfoaPaUSXgrlPXEesf5nbFz44+p2tVZrnbAtzWKo
+Rwvq4igwRboutw1zdrbFvWoQh9WfmppN+CxJwHlJDcbOBx44KVgUg3Ma/Yl
SewsjNp1+vnXbHPFx7XNAU5URc3v0yswKj9OVca3paae2wqdLhwPOk2b06pp
3s03QBqJ/b2ho1GCY89PwqC3X7oSV7Esu2V4S+u5t2lUQkjQld/h08E20oci
EWDJTtDB9E5KFEiMXCaiwjoD/I13HlyASTHRFZb4xPDsKLpC7pMFVSJITYfu
VGV91gFKi8bklEN09zhIDpwuwEs/0zR1jvpZFaXqdQC1hW/+4PfpftvCjVxs
ApLkPc/uSR7nE+kskLdgfpJYjLRKTvh0JavxAoRkENP1Q8alVBtdjNZMTN1Q
kKdq1s/6qizoAMAxF9/61oM1kAeBluOual0LoJm3ZMKBkxXO8D/xKnNJwcF3
lzJxM8YKMiugYFNRWsqFYFbyZ8guXXa7+jpTXFtMojHAYxEraQ/Trs5S7Yt/
z6jMnSna6OATxGHqWHhSIfQZsZnYUj21Bk0aMUeaDCEnRld93eDPunOQ4BdW
EKf6ch9t1X25HDAefg2qB3z2kuQtSAwNH0xyqvpVWhYIRfp0LNBZ/s2CuvEa
qXLF2uAU6Oa6qQC2Ozn3kZKEYr7ZwiGkm8Cf2JtUmTBwj/tbnQnC6lkEb1SR
Ht287raU5FKNnMk8qPkNGRkHt1cXnOyd972fAvnKyaGDH5JxTffQhdRd0cIx
rMeUq/Wgzn3yPv26GKHQTB+nKdzC1xd/7BiScW40tbQzEK6MIA1jXr3FKYa0
q/P7myRm++HXEONsqQQ46MR56tFdaeVrpvlxI3GGq8gG8YYq8WXxENrYLZej
V1UaBEfBNwUcRFR7B1jAjSlTGZs8AvtKDLnHaPgkaFSk2kiermcPDemmDFQb
u/bRHhMIpzfhU5BWdTx/nsNFPIn5F4uJo02/2TM/+2B8gMETjVt4tOlLp2wm
1c4C9bLmUyGswR5jYNJPTQmkjj2Y/ugR+vVKJAJPGdVZA7riJX90NXvmN6eF
FsYtA6OUkXIzPnFhPNdCK4LOpe19itd2N4WwlFMABgVUYcp9gwXcKpv5+mw4
58XjqDGwBZPowlEiWRnJosK06sCRrl/51mINP4OMoPhOWL5JhW8tnxetwIrs
pg2eIvN6z9f6iMZwyMCkIGbWR/haiOrvPG4aXmdqxqpfkQuJZqTJK1FMelkg
EyI4+RORsTJWTDZZrDZiCBFcVHiIDNTzVo3VKZIPf1Ex9A9mvNsjzQPlCe82
lKIraiJdgw48cVu7Yxh5bWb8d+wR3UAa78P+7zHBM/7O4tchwmBXtBt++kV0
SYqE13Fo94MwL3uDrvMj3WvNWYSPjruo+eC1X4hA98alAk20aue7Jo9D3kcO
jvFlGcC2LDS1EGCQNY43stClL/wPbUhRQOWRoafAw6u6mYjQcBi/Gh+7/V7C
f6F08dVO268188Dur1L1/kF34JUIWb0YrGm01UZFfdUzTxZhMZ1Rq7KjN+/n
DqXMJoFaIz7mAhnOWNd77M6uUz0PQbx3w75FdnnDwnVxV2Jh0+beu1H1EpD5
e1svFUMyMP8kAJoxQmCOt5wopDeZCzt7w+NLGoY7QuHuVVkPlXcw7xJcvBIl
6fSQE7nqRZ0+7+4LC/SPopXO3ZMAj47XCnmHrbVY+RuWXstPBqM6RC0eAILn
wf9tybw6or6wk/1H350USr9CBrnDQ6gJw65IbcVOkhMEVYeVa/YLPrN5z2S9
4ncot3tVDdGyvj2XeXMvmcBnyNYuGu/N9jgPybbhtjU/cl8etD+HzPrMjvpj
Epx83gzEn+Vt93x9sAE5ylwqXVagl+L6VRCuF9bCKqfkCb0Bcvl1oAM+G/gI
m4oJv874XjBEIE1EWksL8iBrN1iVrarfUUaT8acY5bog/Ai+deWuYkfx6JVg
uQXATTpsAoU3btumaVOGkH5OI4+OItkc3uWIdVMWhNP7sOZoCJsBE1bHeQsG
EN1HJjeW6Oeo6Axp8/pR5JeQVKGytQIEIMpRCWfFwFrQFV7mi+I+8YJ7SAWw
jd91a/ktfT5iXse2oKTJm1Cur4j+eIuOjrnWPE1odInJ4B3ROAb85cJ8PmPb
rewV7yqvNGqtMl5obwI53kNXq/BoHPWpAPa0EYd4WPENPEJezdf/hIn20k8T
46TNkEJDmZ/m0KcKQ8D6sanLuzcM0FMM2Bh61RpWoU5PJAZpAvwIMK2F+X2F
UtJ8r3ingl7eJ4qkALIgWhLuLmqWuQycqTmijXj3I52CpXI6WqVGiViRB6K9
zjUfuez4sjrlaNgseF8FHbrrelSOY02qLE7c1+tW9/IJ6sOttAgWLD6ktYvu
bR8rNPa5jGxOqGCRLR5uxgZg+Am26CX5mtGuYoKC1t4RHXSCenjpKX5T2/iw
TVC+JDTp2Z7nKJJAZPxwkxC3lrqHw8ZR5xp2H01qluLO5VM793ZfykkmUcwT
BpUk48V7DyDRiFy/NMoXbi4Au/kdAMB78zihK6GEVViDwOGMe2k2i9nAMJ+q
tfGeOvWFR8sbEgGhjt4vQBGZRZRdLdI+T+iS+9wBdSCUb+1TVRbqAynJH0Oo
WhTzDBZSZZGSmUxlj1HWYeGfch+/Dx/VF2e8Imc9amy80cv6hx/t0OImMNKc
rhdPf99/BgcUsFfO4m/cf0kFAF7pP9479csUTCVu28r73zxiybjRedXgaPtE
hij+7CH3PLIOavDZheUlq1aZXLS8S3tkduELyrczKMlR2xGsu51z9YwFE0sr
bbyuHd871zIr09B3wv5l576LhcOAtkicu9HhkS0oVLpWsb0TzPczhQ/4vaxv
UBw43b7onpL+gCnbW05I2y9v/Ol7LUJHfxt74yugk3mBX6DA5j7646XvSKAY
lQQh2Kh1+7pMew+hdvzVfXMDwPX3ilnqAZHQwE/Ws/wKoQ6j603C7P5Xv1Kt
87kXphuUafHIiUD0M4TfENfH5x1U4zoBr731SA3I2M3CGl8Gm4X5KvhOvdl+
XdAo2VLiGGDdi6pBDUlVJB27IjIXvwj4ptDzitFEXIceqk1dw2zFiUgO0ykJ
Qc4ZnYDQol/ZKRoKN070zyR8mLiVYi9rY1+XBKL713VdE6AI+bv042izJJo+
mkbGvHqMIxHQyDVAP17nQ6rqB127kf8l69CVbJJ8UOcw3h/C/fcKgYyWX5+g
tfXRX2fIeIUrlUy+ltIPDt8WMn5Upwuk5IUDlMnOGDPWoyntPH2jCi54JibZ
jBEELim7JZU2qzk4+vG6x6YYoFlpXKvoXarE8QejDrVr09ulGQVygIkxJBV+
J3jYRbmerhSs+u007uUOJidZA6awi6Jol9Z6WlaQ5UqxaH1sy4VzgGlUXIuE
C3mdbukCcVoxyrVbQC2WY8pyQUgEA2UyWhj/C7rMA5IUPdUOS4DibQbVGLB9
L80K7Rj7AB/5UFT0KsLJGUXFrzOViiItw7MYiFCvkoN2ufk0vPulLMj0zmxg
+VE3ja2Xx0i8yoRRbqu/WhuLhAmxyY+sdeDrrqJ3cElQfQucTVkf9LD6jwMW
S+OkL2Xllqjuj2VPEMPprQxDKf7XDPwG+YTWm6wuVYPUWXkSY7hg3UVM9Q0r
RLQGTLd2rGN36xsXgxEk+u4hB32WtjOJgev9EaFO2/fwHFriIiPyFIJBQOKA
vEJkojdZoXZR6RXytnkADJZU0lsbAJx6IczjMrsiHnNlsqjk2eKJvacyFuXR
NE+Ye8I89ZYfOVv6rAW3mpw45ibNtgj3ItZuZpeioFDX6FStY+FuuEAgGBDH
zxFIko4TP7/G/pbhuPsp2MrWiKwOznKid+X7tUuVYVNZWcoVsveqRzfpW2pd
dfmpWSeZGXydz15qzx5yXpx4Anl1obZ8cjVDLhHCyNu2SemLi0K14mcOVifa
2J18CleuT+81WQ438NQeKsz6EF4imMl9B8lPma0yeiNhcCeFkf8mc4BcjCyo
clvdTC3HZqICVzQdAvFS3xf8bncZzshRNK6ck+ya/DetteAfj4B7oT6kPLwq
3g32rFRslS7ud3fl9plal9pY7gr11suLfGbawtfwPIB53qP5NByShIkAGVKD
tgmY0jUzySjii8VboJQooxDHySM5MDFiu9+edQ7TzuB6clOfCuzYaJ/sLPaW
3zsvy9oTu9+OaEwLEveKvqWgbqZ3IUjNBEcLyZ8GllNFpssh+2PLUBAPznA8
Y0CsYshzYvlCWcuea3yiBZlAB/E80tSrPO/MQaoO7M4mMgTZrX/RzJogsONc
Rp4drYY4Grt5yRlgPIL1JVBbBQFxGPAwZoYWBU+h0Z2I+NsWzQDSlVtfJYWz
iDZk+6RWQ4yqdgrxo8Z1YPfNBrRtH7WMGajiP+PYQWIyU6Fon6sUshchbVuA
oVZSWDOqFHOyN1/CHONuCvPrccirWKaidj5/rxqpfUAXliS2AEHqIvY+7i5s
couo+nmL4+LugiCB/2GsJVwBWTY8+bB7vnEH9/UU11PmQ4IvEasJ4AfRKLZw
8e2CD3bvdoUM09rhjYl6SNyC3Gm6JdE4A9Isz3shOXyiWFW3DQ3NA9c3zSuA
v6kUelWb5x+mg19AoI7CvC8OdbME3QfhZh64+Tl2ajIYGudDBbPuBWua0U1U
cPC0My3shNLymdoG0ldMF1B8ZfL2ckqmDXOAbOhJUBz1dA3a1ijd9YSkDXfE
v1ZEGyz2Jjn6ZXfG3zQM8XK2z+5+ooQxqHLMUdM/JD/47/gEbkLd+OKw4z/n
n10Mbb2dl55oDpE8AzWffIavK8Jds5GRexzlfjFivl37fu724soen7QW4Xm+
fLxzgu3DwHcnh9PxwjEzBDmRFSOZuNQXFd+gcJ0MMWuuuFQjWMSd61grZrPL
5nVXCwNBUD7iiQnNko5pv/CxApFZfiVyFY4qdHXPNz+5hwJacTfvIij1tFoZ
wyLssD7jlhDJpoSaW45lGm7pWKb5OkdMtJN5QJRP6VOWgQMmRg2LraCN59+t
G7UgNSmABz9auK3hFQRmQG2G/GxWnhBoWoupIriqPWWOGxLW5eMiugiOUYJ0
FNmUNeHDlf2xmoiXUb9gXDlDMu9kVC/oHN0eypTaMUGG8O6ekX5rwvECRcOy
ctvUMRPSQAcoAXRV4z/RgqbEe5YtJnMbMckGmtvB3I8zeWRDXncP26p4msyL
M1EBnD5iw4NWl3M2GyMV9z2Zn4FZVm4jzURKABkRVKhd0vdeb/T2P6OUoq8W
r0AaKvJpt/Pbpk7Q/vszuH9vwkDCjyGStdKNURGOcz0ghxG+A98YrpTf9lES
IkljDxGuquCVUaWaBfaPgUh0ivfAjTZdnbhUK9PEunCIzMl9rfPLMXAICdEk
a+8PJ7olkc+x7CivyALU4SLQZjwAZuERHVs90IAEHp2s1Wshs/XpPxHNcZ2Y
jqHPBK4KZatJgqmIkg2v5yYUs/ooc8rXkUeg3bbdVEDF2kHwQfBnYNL0yFeF
NF5FqqkBf7alIPdZ6bbYbwaaxnq0/uZUQ6O2Xyo9lPEOa6k3wKrTQPo6qysp
4O/xFax0X9ggycV/ZWvI0gv1dIv7UTEqsWX98LwJzW20PSyJwJsh5X4Uqodx
cLtL24s5gdPAFcOMspMbqcy77ymEPGplVzjdqcxzWmxN1xzoiORo3cLDoHmW
Z1lcPyb6Tu3wBiWMwwDkIFfA7al+aFBwV/GyOFsVqvEaeS/xx9nw3pfkywzZ
yqIByrZzkSiaK+CfDE8Jg6ALEomPmQrQ0AYe5G8nZN5cR+72mcjgFyNAUmbW
pFvu6rDlZ9sx2rmK6zETb6Nyx126UPZ+k82fkrcq96l76yM/2ZWf4OhbHaHY
OqKIhyQi6B+T2jiXaj4Kz1nt79cZIGMOsBo7w4F0Iza1+PWIj3iwIiFXEAqb
tq5u/9cNhN+6nCPN3fq+OXKEfy7fBdSf00W42ouQQs4R8l4XebYcNd0rCHFH
u1rAde6rYnI8YSNIPXur16ZKAlUSyJHx2teGKGL7xu2w5K9YemV5drJcixsV
3XwjUs772+YSVz2WlZB3GyIpSN4G4GPmGqh/TipzUVQpOwkUSkll16Vg28hq
kjskmRhGFbef7ttnq4IQDauJ7Irdc6U7g3B5JTMUxX5xFuvvHkgbPmA2H9yE
efq2Dk920Hdm3g9uOxpsYLSn7X3BW+mhvUDKuq4e6QMZjguPZV0d0pfQVSIU
VcUcPj3CWT2ot2ZNop/44FTy/aAmUmUGLQ3SfkZiR52VimhWIQA3I/v+U9/d
+/qyEojb7XvU2fjx96z1jfrSRMNi7pr2BATDkkI0oyQYBv1rraO8PSwO9ZNd
sWfJ+GVpU4PPwcDAtYtlBykXvV7J0SmN6E0d10IJr9vExciXWc/0B4qwb4Vt
EUkbKxcCwQKgUoSgKHQOiHcXwEDEkpRHjGax8hSea/8q6tDhOwlS7XbdsdSV
xA9GTT729Ib8BElCOnaY4vUCO8yKV5vNFc98crscfYw7WrxjEcsNnrl+AVaK
Zmylf7WI2IvaVWkSMryO7EZAnttglBminnsy0yeh8eX+nv/b/C1UQXAgJ07x
u3YZxBZN8Tzm+Ip4wjolRo3aKdFOLRRR3tsdQWdblbHBSyYM+SPgZ2A9ueTL
wdk4x1dtHYZyNbmeAWY7f1Fq5NIvlq74nm4TYG1IqEaPYVZk0qs0Z7qCLY69
ky9tDLT91vB1gQaDcG2UiLYECPyUSIJURc09DcOphwS7Zpq7marC2rx0WKX9
2igNMMBTl7jIQh8/p+ARHwITSDyXbS/DpGB8Qtn/5581s77cLrcv8KvasVW7
IpmIeIcBZ8bzFdanIZsZAHJUUDxwDmhRFEJ07MMatrt1CjZWrkqACbDEs34k
RRxeCo7EwF+0qKwyCQLiUqgVwgG9IdmGT16kUDpOpvCgdHaMt2X9g60btUVH
05m0+GMnQefjx3RglzsAQvUL3V5d4W9kxn2wqcXzYBsSUCzEHm4SEbV/fITu
xGMlOPm5FzRdOtSfqxcUgjPN2ss7IaNI6iedNBQeij+QbaUA4hzJpEWx8eI8
86OfnHVGra92Gi5A5s/Y5+r8qIWyejthXZkKdwNWx6DayQDiKoEyFhUIkY7B
3T1pgYXFTL9ohydL+yfQLhuGqeXpXMGpfFG5G7AmQsOwPrJfamTgPhaPV8Ff
hNy0VsfNwVsHEQrmA9gNDfg+hnhRXNU/NRVo2YTGLYrRJTKVvS/vS3Pe9Yjl
CaZb+e5Dh1921eIq4+KaIMy+1FRixK5eXbs+23EPPb29EPoXOHoL1zMSDGnj
rBJgNVhgu4lPPZtyCcR0vXKN+piLKHvdrwC9vUvzXoAlP8przAzvgeesfrZ2
Pdwze3GR5Q0zSOwFl4txVBKw96rNyJAZFA4tvjBRsMYGLyxBXwTea/qhQ3wb
5GEmoUDxbeK9JB59KySz9QS+BvitCpYUNSomKwyQik+B94Hzp30MuqR62G4G
TH57/KjzdstytDqZs2FF79mqW0M7Lrj3Xxu5ZoZVk6v7WgSSZfCD59OOSVwx
B5hTqTGF2EVFuWomOAtmlheClNFZYt8/4wddcmUpGMOCOXvyphAfeY/yWObS
hVNTAuXaSyZ+9SGRi8Tz9mxMyVLZxoGS6o2ffl4tzyUZlPlSys/RbyPZMl0N
g/p5v0rHVivpvqkJJzS5T+YKh8tK9gTw+ESb7AuDEkg4CerKG0CbJxcxD0eN
dRRlLQXCH0LCCuclntbGakh7CF/YxNPIFrN12um9kwtfkyM8rG3CpTDf84ek
m6oBrOzKLYYmIDdoX2br01yInGOZbLl8IkEBkbE0vJFzxUttAvG4GnkXsU9p
jjzcXGOCG/JplzeY/qoRyrrcX+pteToD0Df9xmgEugsAjQnKOoCj9bwcgGcG
jQ5kdalhqzjtY871Nled9AmJqHILURyqwnKGZuvpn9nB+ryVjSc9iksnx8Qb
loj3vxB5WhO9XZGPkQkbAw0zuMS5N5rQOcOKvuyXRzQWzvenuK232MRMhdWV
zNMyYwmMhtwmglkne6W+EnCNpn0fYY5Nlz4BqPJk4lya5ylTyy2IeRh+BOSq
7sKQg3B7tgdqwYqwCickCnVVn9Dc4pbdDsp9t8B+J2fdHM+wkHE/q4r/tPX/
nBadsXfbISkaxNpoCO5D2A1BXe5IrNTrdBboKL7CdWBrt1gNzgM+EqlwVvFK
3ixHClfwfT+ReRZbIZOBCepcAkS6wH/6WOztIofl9ybF4ByClJKTZz9FqjV5
Y6AdNzgHDF/+nyTbSSqFBLbAgF/xgtNw+CHYLisIG948fi2yCwWXh9jpu3MI
WXm1yHOPm+cVP1UtnrALVl3GXUzzSakLYOOmmIQQHO0F4dgcVFuNeespoqTX
lGwOVX0c2HtgkzU1kAY0dv3yq+CaOYEOhp1vZ8hnqkU16ckTLA1CgAbzUG9S
yRbbhih7s3j2UbWluhW43mjEPY6AFsIBwGuybQoUT+eMO3ynN/gxERPdRGWU
k/oWB8tIUpFSmchjh/YPc/rUgGGcggVDDYo/ejQhIugc7LsjMWaSsiKH7Dct
tQ05REqEa8iyBEMOpqi6qpUj3ce4s6dei5UKUtKxEXIJc1Gs6uJcKDY19sek
Duza33MBwV+9kT4pteNaS/dQp8HjPEdceLdAaTcXgRF4XSAdaQsJNaJUlkRg
Cbyzb36s4lRLiLQlhe2JS/M3iGLfYcPF0m5UaovV+UaSO5nRpgUmYk3SCasN
YxfchzJkucrrgiake4/Yo+FAGHZi2OqNVRKg8tL2WODYqin4Rl8GqJBzL0U6
U1J5N4vuRxt4cBc/WWNDKNkpKostmx+T6JEvXOQnvyy78T5qm6W82NKtpRsR
C1goBNozQNyOJWkopC+XDiq7p1YrvqTz5sVpThA02SSee42n4UbGH3RGq0zM
jbS80dSlpxy3Le5pQz4kgm6UmPqX0a3gyHAvx5spDAtOjpUwaJ8xuDZzAyzs
UInQB56t9JxyEyI7Emr/6mcuc2K4DLP083XugFsQHqe6vh7Cf3PplkTGXMe+
WOwqC7bFZG8+td833t64JVInWNEpG34wy9aZLVutSK/wEvfH0XxdqFOnyBRU
W9edSEKMjGNipgT7W5Lt+JnOViYBbbSE7uBsMtEec97QJlrE3i7xVDmOLx+M
Xz+QThTp4NmhE/Cuu6jhfVGDn1ww8NHoVhojOXZL7kscKadbmIshn/pMTyPF
BkEobkAQCBeP5KyZNVQ6dta6IJ3gHKCa7wzOoN525m8p1HmHrS/g+j3eDVhU
1dUN+KqRn7NBPe9CkCmH+zdWuMUvgKfXQ9cm8AtNoP4DjEpK7Bguq1L6AGka
ewg7Bc2+HGHXW2+PKmenA4PRYZySNnCdAjkHfgIFXtOhhyI7979paDnLuDOG
F4GH0DED9GPlwISMIWZo3+C9b7wWCaQAoTQ5fFKs8ywJPwlHzzzxx44z8gkE
EJOEMUutoF8I8F3VWQtGA2e5N2TFlYNZVROamFlfZMsgH+6SzpUxs+FFMEjF
a3r4348ogK2KS8JX7drhWFVZ/Dl+rIJ4edgUiBYdxcGntbGsys6LlxQQza4s
abh1SANIbJQC8f58WyBO0xQzjgqBRc9lNPAHUMFwsPs2k7H3jH1hVMpsGGb7
YHB8oH4QSUDyUivrENvoG+YH4BiVWRUkn2qnx3f62phEqGXZYTfKAUW+FZA0
YrxGbU3y3gkGdgb68BvPyM7a5vp07tG2wZKCF/YP17IV7cifBOKh/tD9zUHc
0tWAN59IHyrpmB/qa9rZQi+p9tIdHBxoyQgJ7DDrFOYkelCzx5FLLRqpY5jO
PqRzIufDR1ddj3pWqgnG6cUhmsnGcR2WHJg/AJVXP9LqCMF994cbRzgV4KXj
KHtfAQNSJz+RU8Y3ZJfpIjzFaTZ6QN0P4h4bYGJVu7jVu7Yf5Z9OeBTqQaiB
n+2BGU146itV0q9RVjSa0RJUrBpBR/DyCUf92vtUqpPHYi8+hrKtyBEThnoO
VI7FCAVQ+ZOtOs/wVWKEBqwmE7LYe8oaXRursh8O5HCqrXjglyIMZl9A/RLh
56DR89MP2rw0bmoSwrjZNagSXmLDY+gCkEN0Ds9sWtiUfZ14e/CDvNC5VR23
I7ZCyKZLserfCYOVD1wIiWAbi1t0tFIn2C1z8MNO0a9F1F/iEnO+zyRq+6pm
HoyZC7iQgmnDZGksM4+7W8ug0oOzSwTlEDDsyIo9AGRq9fYU5j59xzJmKjvw
1D1Pl7xj9b/tCD/YmRtNf5iHjI6JismGv0pWN2EfDuvry+htEbo+qSov/cH6
Xh9XHYW5CT2wM0kMCopAeMMzYLK23REkyZ9Fwn8+bUrXv8K7uQo+JH8KEbnf
kXb74MVwvsz8qMEq98MBCjXl9hP0ABWC8DGqgM8hRD6xHkT7cyM7GUfZxMuq
udilPm+3+ebwbhIfHNMIcLS957oKWq+oDUlv06Fh2mednXO7jK+pCL4BDSNJ
deJBVp80MXd0sKhA7rRJ0f6fjueALQEWagwu/rlVOUDJEke9EO94naUs2nRE
cF2cgMJr/5hIx372EmOf0zpcL2h6qbh9E+11ZLE/bkPMOIrT6ecxrJnvDbT9
PJ3We8P4XaBZVZjKtvD6x46Ib/AGXLvQYMLPvJcPp4x3QJCAkK6gQj1aqQ5+
EWa5KgB2U45Dd4VSmfS1jdaOFgrSy7AtD/HI4UMHnfEIxx7EniGJsA1N0yzr
ZXaX9/k/bAjPaZiSAZUDDhmYSbEeMIkBe+lml94wI2dzbZe5dWA3Z1brUJ6/
zYgnGyw6cGzO6l/Eo0XtpLQ+qp8xM8+BSF3hOToGHS5/fsCajsPiY+COzaHV
d72hEWs0pgDwFvqPvaH/SO8Eo432n0WaNNelsEZ/3B4ZgSewibDKRFpEFPQ0
S1YIy/RKOlsnB+iFYItQLR3mYKJgmMHL56mnxh1fKpzbjuiUxScprUTrLouJ
+dU/rcEmaNbu4qeHhNlADU4U14zcJsN2Ts+mog6NV6eV2XwvT0QYizH0j7sR
e5V4lYQAJGsNJ2fxMkQ7AHpWFaNw0cz5yFtux0ULHmIZ2PJTN9PGyvMseLw2
t3oQqaekqGLyKMaejhHnqaVDjA3kMn5bKm8MUfSTI50/dgFnz35fxJGXLGtL
VQQyiDOwQF+8FsdW1RsOCDfcRlxTOrGsuru+NeyMRjBN5X1y2Wu7Eedsq17m
RvUc9uBSdZMmblsE71PIvflQ/DFXiV+Fn3cZwmoIIT0MO3/emDFUFLwjawXB
PNrIXg4yoD9bGkWKnmi1Rh4IWH15UWf0BTlPJ9LiYBmbdY6tN3Jx2Eh6ESeT
Q4s8do24arGTMHv9CLjXpL+R3kmSzNcYv3amv72O6E4L7rhv7HHJ9073z25y
cHtNqP4uD8rstrBQoULcDsowap21mpXAl4dXtNbvNLvgd0jHNgqAyLC6N/Gi
/TmBHEZM7I0m2EA+BifmQahWc3SdYwD9ZWhM/vX8/GX0qOHhMqfDK4NtGWq8
bLptVzhrFiiDORUplOYWnJmuB/Sgbyq66IQskBcU0U9gY0IRogUYjpAGkYnH
VADLeGe4U5mIR+akTeL3XrtXxeqYKA8PSAdC8IKf7j2qZZrJQFNTaTV9+mbm
sO/nKAPzd413BQ+mI+HsGKu6Ihup7XH238dGNB7Z8NSPyP4DnPmg5/7oiWzV
qWWOyntJ8Fwz2iYLvv7IIr8XrlCiKUh7C9Kzvc6miAaVkCXyCpAjmN/kPvpB
v/VxjCC6/O4Gqk0ziJLmi7nIDjAwZPFpQjrL5CgwRVtT+dHC2QeBZ+tcpv+S
csoKS4WGO9uvTH794D3w78Xr53zPu0YJuKcbKe6FhGdAFBhiRo1rCWnlSUsA
efRxHO/zjMTVhHP9pBp+kgG1uZpUyWy4z3SB/jY555GHwBtxRfCVLMl/9GtL
mPfvY2aFYZfp53Xnf214H+ZwJ6qZ55hsUYBxKI1F3+x19Qa3WYHDE5UerSwf
n1yMXG9DHfSd8qXolnxXuZBsjr0o2LIdmn26Ij4kbzBsva8cgGL1p1ASYzHq
AOjLQlAdzpJ2d2W9+iagei/BJ0xJWXQ6FzDgUIbnxSIq2JFO1YrRg2PEvIyC
Weyv54oGONW/+Ej5cDmUZc//jwUxjc/QGmFgaNrLrSdejtFPVI6ZdaujVmt9
0HCWgH4XZ1pNAWCpU7c30KKTs5RAdo+wY+Ro5DouX1ZlS573pX3f9hMfNnnA
6koYSwZ2Nd8TRyjzWknWrmy4J+jqgzIR2L5bVKbSq7rzXEv6ePOgnxguLu4D
G/BKCTw1mDDeMDtew6TAtk/2eXurhkFksBVloi+9UPIKeJyRWA0TDOIypW3h
VbQ9wlko7UUeN8u1go8kVxEY49kFF65wGOi0R+nCS9Z4b9z7+pb3x6CL3tlq
kOB11w0ulsU0Jvpye9OWycwJB0uriYWkMXnWKODpANww74y8EPzyCEE44hm6
wLf/z97d5HyFylyXJORtA1INuRa5iWwP2iSfzs24eXtj0kd26XxTP7VkVVT/
RyP6a2iu1J39h9o1juIIkYvLrUF1/WPOjhqFS0I8xvrViGonmEz+lMb5FvaU
dOfjseYXPKSqXeoFLI5hHd5AbyhugQ2QNnd3RAUkB4RKPF7tStnTHICe5dGv
bhCclvAC9d0bynjz3p44TOekdb6ofFHcZ6PLnGQV9bSm6a2ovBIEYjQx2VG6
Kt9tuAjHGBLG7IhN2AjAui/sTnd20Mq2fFpOj2jL9fhxZNw0FraU0CWVBOvC
8MJrtEscWVzci37XzCtI9HyiyWjQup23wHlq2oPsN8yN8x4VlmZjyjaKG73B
PA8equY3iewsgQAflyqGtjtolFxQIYhWRx9pCX78750M91u0AZA/+1D3MnSq
lHgbwG5DoSrD4PGLNuPTRa2YqevTHXtSwJPN85QMLaSx9jI3mAl4eu8uu/sj
qPKeempU3Q0R2NfRfz70D1YlUUjYNehBz+vn3q2qoZZ6w5xO7ZmTBRIvh+o0
2ZYhhQzogvdPC6zyce76hnkn9jyRKf/kffZvtcbW01ocM6Rzn6ZG6d3alMJK
DlsmGI57Beiqii2dewMhFnrYTvKF5hF2hUzCgiFBvK5kB02tBaREAbz77Q8E
e6S43IOZLCTJMAOXVtJ9KsjNfVOFRmQ0JSv+V6HlxoImy4TbeIoGOCg8PnSy
ofQfa8UAbgsO0J3pZg8sWTZpDXL7AXOGEQafGCih7dfnBtIEzrLerMg18No+
+MN8cf84iafVjpKUG9kJX6zRcKZe2w5kGO9lKTPdg9xuquA8YE7LvhibWkUU
+ugsvXjjSUCMhEGu/ILAnN2wBsyR1gEemuvJjALukiZN6FlAkHQqSGrzqXnc
EU/xeO2LYwsnQQ0Lz3TNLNxlt/8aFzQFoi6G3LMYE20WympHH/O7KxjHysl9
lENdL6D4x0DEbZa/5U+LzkfOiFZ/Ozt3XpbTpfPfz2wIe6lQSNT26o3fL/yP
bpn7u8WZevYkn7JmwPnTiciHEIb8AH9QVgG8kkPV/taHwA/ulpqjbzjryTzz
UNjIaP+vk7KXPJPHXnc/0QUlbUgepywIVLVeaRD8qTPho9ZPUj7JhHypYpPz
B+iORQufAc+R9vKyJY9MYrmsOFrhqENF4qF5tmXeJHHgYXZtP7Iua0r9dy/c
3dxUdFKd5hzT3G+9vHSDW2/r7LSMGtPamMyCFkbe0KfqasUdd00blioBzuBt
22ggZ/obk44WIwdI8IXwbZiR2TTLgmpIH/UxZ4tl5VB/HTW79i+wvRY9zn8a
sbSTbxsRJ5m21KUQM++OwuKhXDf/wrsqs4qQU1SX0syTdkTBAbjKr1NBZ3C9
/Bfb08XNXfZ2I/ljjpffLtXpa7r6u9p2t4vJycZbz93o4jniIeMhnD4YkYg9
FQO/wpAQKSFYWub9WsyTQBHysVY1HLDlPmmSBEpiPJzTYZW0mYPOiBtFfpKG
BLyFVVOFpJXGym9+70UdaNZ+QhMRLiJCMu7Au7HaSpmQQavhMfj+nyQh4J6g
mPlH+BIEU3c2eYCvxq7unf+n5V18RjB4V72qonAbeYxEEqCRrJCiHLoiwp1T
9V5tES8bzZVktJ0hQcis7Y9CRDpZqs35+PMXTjtIYsCpKB0tXgUF8lqCZwY9
vM6hLEz7MLEw7PV4SA4RFNEBW6dO3hyf1xY/Ai1oEAarVnUOcm1sMgveeH0f
8GMqYSIUtxp5p1SLrnitBW2pvUw2mECqHcXJKIxjo/PaIe6fr2dXsKbTs5DS
MeKXovtIV+vijVUbbDoyFUc5A0aM9pOqkZd/33ihnzIHOZqyC6sKOIxn4O4L
nAAhsytaBA4f+N/jwu/cIAJFLAF6srVuElFlBmFTE1Ze1aTWG2zzc7OM5212
qWfETk97NsYLwJGKuZWRq52yRX3+5EF6MGmEdSuJdqeJncspCSbL+iW4feG8
v9KuiAc5kfBmK+BAkk1Q8ucU1Z/zG9zCO+oSGM40diqLhv04hAhV9jmnuBuY
sLln2azKwdIcryYfzcOLbkFNMmwZuPU91wOIJSQHlgGVvV9g1vV8KOszjA16
jDLtFnVPBaJ2Z/2l3Hb5IdIDUCzDNjUktOWoGJPHPP7QPFKwzNLAHpE1xnHL
BbNFjzNJHjwE71R8zhhQQvw0rey88fdvZ84Dvyh0a04w4lg8Prksk41MoGTc
4NK+3V+pfeQoMm56b+BmCvuMJGDIfihEZ/KS9x2McmPTUq7M0U95sL/hmpNY
qctBPymvUGFYCaBy1MQT5kCCiBSBcm077sSSmkgz1aoWrWaZ97xHRDrIWyie
M/JVSMQrELhShAdBKXcX7GgRIgayKOlk1EqIGCO2MpCrG1uTdlBjqN9Zn0Jt
5f8+oVdyM/6PT2u4bmB/ETbU724Dy3FnBmzWW3KwxVMf68w5/qIngEv+1pZm
nlbrYoDxcB1l0XGEwYd8t1J3ZihF9UtmveKMajxIipDo6tvhPWFXjK0bcotb
zhsMgJo5h0ZNjigOiQXaDd0YnrNmkdM3l5tCKzzilVJfeCbonWYBDt0lw7zk
zcK3v8do7beChS7dkpqJSyoznuytbfiAMjZVZkn1sNi49/tYf+S1VtmydBz3
dKiJ+GgTVpbZNpq57846Mf6eR3njjyf22iD8A1d60FtxfM8s2K6v99GuSj2D
LraohUg+6ApHF2rv4eRFe67DgEWl7DEjvYfmKW3IwszI6HXN234/uI/VZ8t3
7lwuaQ+kgvCRkdu66I2cqA5B/TszJkvGOZ8mJswnDbsRaKvLbkPttwc+kGzl
TBow0h8mdx1M0tYHEMTH5dZXNuu2QeQfo3i9Cz4YrEhHhPt7Ul73VgXGEZh2
r02ov/joPMUtnKCSEZJOsqNtnyO1BGQmOIDahhFLRD14d5e58365XqepCq4v
4FQxaPy++XUNGRjc0cuMBm4taGIJ858Sqn6uCLj5V2FbUeGms326+vU57Ft+
d9m8uXTaHr9m0tZSZGO98yBbGtPNqiuq4eRpytvT4WWc6DhEQW92Hekqx0o4
iaGobFAzQ+HHrb2PzuQTiB9cxFfPHX3lREdFIxrLxrzhA56d8qA1rOcp+x5q
eLEpfqVH0zs1a29WlTz9qCB3xgZik1zzSjSigeQHAjsSFC1syJ7le7AuChHA
PT5vtwz3xXgeBR3EiLY5qC8NugVoMejmPbOwmxrEJhcDmsKeFu3h0A+09O41
n9+NJy9wHJQ+JKAzypl+9duEzbE1nd9q2TNIzEZOnjqzERRzjmWs9VPMPQz8
8VcVApYSHD+YV/MzEIYgKllDEddEaPTPoYthbqMyHHUGCqFV6YJ5FPTnlc9B
FUjTQkjCUO8azUWUYoEl8zNiSJQ0d0vGWu31VI/qUZbG1Ds92pwlQzmZ2HXW
ZQvPj1wdQW9ghQLMBr2S+dQM+/Nmoh3b50WiSSfgP/MroNE53NJkMF+v1nj5
X61mPog+WqziWSxMZWqTAQFtjqJ9A4JVJzhNU8bmgv0VUljsYXFreynlg+Hm
WZbrB8ERurZxk4ZnDUi0T7ApAXuplMVim9IUOQClz0DjktSGU1weuF+uaoer
b6m7XAD1nr2uigVKcOKYnn/mIr+wIQLJthuK295A6LX56GRu7voUyO6Op4j+
OycIT2duvU2huyzGLVtti9+ew5yyKvdVAUNcXu5VA8adzLCH4NW3Cfyeo+lb
ALXTTxOKqrHnV54UJ09L2E71dqwtIb1fPcjSyN3UmpDM3v8llHAdNxuR7Yt7
n53xf8B69WGLUERKOkdVZyDOt7/98mvSIrxdASeHlOAYoWGoTANTJ2n7YQ29
4aGr2Qt9rCjw/e/pjhq2/46VfahwcRMidEDtBe8jbl8AfWxNrgghxx57ELq8
Bybrps3hzDnM0vtaUNFQgcnE3TKrdhn8N7GBEeeqQjOmTsA7Lf9Ho/IXkcAk
Vg7DhAi1/Kd7lm4UbKHp0CJmP1p/7JQdm+9FBoWiDtNThu+lTrHiguINLRJQ
OT4Xib9b6gMahHQaWwktkNhdyn4ZYhU79NXoT3nCS5fE9YndBRvE/ihnxk1N
MHdYgx0jsbAIxLZDGCaZwhP6RS+bcZPMh568kOFsG28wSW66nvFKkcMdjQUO
ZXqHCOaG5hmRTyeVnVi+yxyw/xCAkoSfhqNJwiNwocbD3fYo5Rxne7Yd98mQ
WyNGmoWDyJ/Bt398xL9k/3XAosqcd1BW2sCPB0e7DYIv06YO9SCNp3pEaf4f
84cfRrI/+lfKjTQ0EgfaWCUm2nR6axnYMtjbdGPZbg0bSqwcCEDz94GHHneN
q2dfL7gFN7EeDNfkERbUEboZJoHi0Co0Z4ztkHtCA6iVMa3wORm3QlIaadJ7
1LgXK1gCFqA2EI52eUaTY1Oq+ftD/cFJcPCjxjd9nHKI7IoVmtwmppAXfXnq
La97+vINvv8UE6HInF9Y/ROOoYcJCkfic1I/ndVSihu5JR8SmUIeg5hkIlIE
rrHM9DwseodwyMZuFVI167YyL7tT5OqEXQbhES75txnfAo++4i3D9K7mV2Ho
2WRsglDW+lv2IOIyumCszberEDr/B3IgRqBiu5JqjkOqL2PVQ/Audbe4D/hT
NNrybpaljAczP/e0oOtUnOMDiaCGwDZWgdUqpHWXmb7lj+aQeryLpupjsIhl
GJ1sPYzG7+tjJNiWr5rf+g615CZSNOQObBCeqjJdOEkn5+oYXtXCPdpI6O/C
lcVx1fksIw0VeMEESPT0a9MKuNdiP4XiyMJjliuqHlblQ/WqY8hDf96tbX7k
v/nQJGa9+eX6ySk9TvwN5sLGksJKKcRXs1N5rY1tGLRzdISTHB1vHZo3unEQ
ruV8fMPjiCrlwclX4TMzWbI6zx+KhzXgU1tCafYBYnh/yV0FvAtZldTRidf5
wqlwNgfRO1zsWfHq07EWsP4edTmA/GGBf04NIzsjO2GXusLZdNwTwnM2UQDX
Q295zuFniakETW58j/cJVkdW1hArA/YU8XMBB3hKF9xK7KqE+uCkW+0K1mRK
OL41iVF35elqCabF10f16hh/puqFRvsMdkGayVl2xoaS9RcA8VyTAZnSyjxA
POY21vhsSTxiNvDhfYlJVnG+uzdUIV/og8/8FgdCbqnrME5HZU09SkHzcxzZ
v2BrDwlyp3BS807R0Qyj7Dg+bsUc/+15B7BA4dhoWG3oAbVkP5SxQ60WZhnA
mF1AiJkbHrm2OhdZreFfu2mMoRcpgQcd1QPZaSuRm31CeokAPvKlK0SXz2Fl
kEN/DEofNePJparoLst/GzbEWdfrxrd77wy59qRM6nimE4e2R2eS30sLzS31
y+r6OdwfjDbN4nll2HIiKdQ6kh1G0ovt74O+jw56fHuIBYe8J5X/9oRWnyhu
r/rpU5JvjxuAx8zl5K0LSfLjXFohUk+IHA7N+P5OE/CG6q4tCjSq5BezyjA/
FxId9EFa8psDPsD7n4hvBSyIVwtOq0TXckN+Ry5Jiv/GCMx337xfOY1WYvIK
xq1ZGkxMYAiQnnnDRiq6w2uSgyUGkYHWRN35eLqD9AbmNDDPLN5YAYFpwV8q
2FGcsdr566o620FK/Hx81Qb6msQqLsdt+kmRBMIDaso89pAehOWktikdG5DG
IjHNYmQkrzwwqyqno+3oKws1RRuypcX0qzHLSkgwE5OOcCJYfPm2nYdV8GW8
d3iUeKy7hZmyILOcH/2tp0VKIfjL/iXwSM/4w9zHJ2RDRXrOBpLyTlPQ/ase
tZ4OtRMbtCZtT5lusfLYSjpGelA4OWchSYrIwjXVaDsTM7PPVyepf8wMPjQj
wBEFQ+ysUcR4psh45oO3CauF719MfjBmtrd3/KC9IB7kassf25MROgBALUbU
Dep6iR+NeFTUNGfm8V4EFuZ08NCgNhuuyT13KCyIRx795TIEEmG8sje2WZyL
Y8MhPYwATzP8vB8F8VkIptgiEKiv08PIuuGbJg7hhnAt0bG1bn4/c4aYSE/6
SV1oB5iucZlhOzCEU4OCRdn/zOfu8A0wuX1DQecAt/SXznS3W2HQQnLXlE0Y
k9a6MVo3Np7Ke7zdmjyUIq05VYVfQy/7hH6SjdMvo1KRyrBUwOzzyioNpYt1
WkiidGi9XbdeAdVXk7Ib2Snbrlfipog/nFv+6kJXKRcyDkdYkPFRY6ODGnTt
Jmiu203uDsnEbVM0ot063dhg/SnpbYucblfpaOgs7M+1Vpbq2sbONQCdMgYl
UNbh1ql9yHX4To9WjslypecF5hJv92dqkJFbJCfUilbtPtpYunWRMnVDEY7S
pmTjDIU/nVymhhtW2mQXqg+71KuzFlXRmbq5FSdzld01XmNLMDd6eq5wAolv
MHOGAauNzZhr18u3bbe9sO7932EZZUTepcc7G322qzN1NxYsnK0qEwSwvng3
3XoachxwnlIJeBWIu/NhTs+YduAiqxpIJeiKUz4EpqeRAnvnPhxyFKRbC9tH
KRsG6gBgDZ/I+tAMJ+9X43g3xONgasn8CJ2+ojlp8NvOZHru4gINtmO0N9RG
T6LCVqajVHnKh6dJ10jLtkudb7H+n0O0ctcVB+8+1cHfiDoF46R1uoDIoc0n
2m2ac+w+UM5gnzxFeqgeAsaQcxu24MbAixPiExkg8rdQvM1aoi4Hp5BpX9zU
mNbzTdZ0PIyI8x6K+k4enSmwcdAtrbemLT8H82KyOR5Rd/1bbLGIl+AEEBbo
gRoE4O2MaZOAbhD8fdimkNFZls9e1lLLAZiPeiXQs2nbUP9603QAoKQxwEqd
egNlINGjv5METuPJeCqIZ4EPmnYF7XISybz31KiWRWQZPx4Lp2zEKxcMnr0H
fwKMSI07+2AwVKtCX0ofPEv6tgRIyE+D2DJ7ciLhy3TMboi81kVlLb6RKbR3
kUjCVH/iBrlgA/7DWCeQk8cosXAv9dE0jUWm3p4Q2ZmCs8w2/zKUzWThAKIH
Ka1sjftdkyD4A4m29YYgtwlCe5OJY3wJbxHnR2NK90rD8wqImWTxVkkTFRY7
JGIzCPPlloI1wihy0r/Pii9kfI/T9BLg8r1Ox7agJ3M6xaCupv5eolU506p2
iTo6KWUZjxggq3RpCpX1MBkKT6oTNO9QUht1EIeedMwnKFk6s3uImXfWnfkV
WsNV+NxWcFMF6IDP2u4yMXQwLe+0rVtu9ZXcIMeeSPru4NZuRE+eqDpnUBNO
ZIe41rekwAwvya/OKZE08WuVpFhQoqWybJVhEkf2zSSkEn91H/AUfGk3RM0n
+Ez4mn+8+/n1kAsJFxojOF45QpU8LGsz6YMs0Jkko879ON6f23INLQBWhRMi
F3yueYAiLxynDLPbEXBNcZBzyc80vj7jnodNAWVNzKHeMoxE8aCS7bSGbhzt
mwANSeRKFA2jeSGw6TfGEtzSXoYwPH5Q1sgjKN3U+s5F1VKqv2tSfqldmDql
UcRbiFG2RxTvKAMzdStmx1jaelQsicYZQhfHF3VMc2ROCpMxuPKMMmo47JYN
RzdnC9I+NQGOdFydS6IRBkbHpqZ7xNsFQpx4nXWUhq98TgliZJGmENwuc8QL
xx041RN26BLzv+mtvDkeOfxOzfa2kWr7zc61mJ+XQ5pPS3I7ardN0Tt9KAra
/XVCou6YLV1JpOriI5U3mDKDZ0A84acimYseafRlAjyR7WMrpn5qwZ6rfTIV
Mzm08jTgGBXbVLj9ZCkIjDKCex4SjKyuhvBV4QXF0E7RiiE1b2/MwQZQJCaJ
lODWHBoDxZIEdagfxeWC9pSb6P7JnQSpIU+nrgiktdpx6LFlRq7a4yCGmjkL
SM5JWNm9KdSsquQGiDCaDVq/giYWzOQPwR7Rf4r3h/D+8HkpaV2QxizPo5tP
/OrX4yupGEdkQyt+M+BYRAkAnRvx4++4q+EjdhdSm+fnbg0shA+Llsat0xbL
OPKcz12JWIEgBD774VBfLcPU8mPyBrJiaRuA6lV+tTmKrgT7KZTk6ENCebOX
D8FQxfm+NlNROuQ3V3inplbpe6J9gMN5mdRS6pjc05ggaV9mkfsLQlWgrc/R
0KRTWsYY2OpdMfBs782R88j8Qj84X7HSVvVHrRw01WjJMYCO5MRNHHGKVSPA
TV70YBkekzfJJV19Tz3nHAFxImqhCmt22cCtaSkfZCHP81bgcTUI8UDpYsCe
KALAFd+lmn35k8PXMNS4vnNQxNBfF11FNSLCYB+5Z6pZ8js5TL9KcSi/m8rR
o7C3haHhsp/NjrP9bpoeMpSJ1O6ix+i9j4HPbYbk4C0P5UdgCEGbLBR19ogX
1f+qxR8iGgtlUloBaR1ZWVDcvNo26xuhxpldFVboixPR9v6En61Ex1yiZ+nX
0tP188mPnfz0B7CXADAsNJ7BK2l0fj10Hq017VWl5z6dAmYp1wJYhP5CpYFO
cfmZtPQFAn0eNOszq3ZIUZApBqRNxshN2nb4bSUgY/Bhn49mBxPa1r6meXac
utJM4l7iy0ggqHu2SkOaH3B/CLqBsCwRhgdmci3AhRV9c3xVd3BKs4PjA640
lTmtP5MWoqh+kbFHO1egW7aAAocm+3RP749NDWpcqJRSE9tDF3AhhGy57+nm
RWWwR4dT/i5dfZ0Dh+6sokbde+nfVSN18maFdcdVJ5u/c0kPnm2LjZx1e/tG
dm14+jXg1abBJuOHgamigNCF3Ev/IXGNolwIRr7wL7GP7BL4O9L89tgKGbU+
wGRDl0K2J0E3JHqJBctHYE4goDPm31mukraAOC1EKX8uTEqKdE6hAeI+nofM
pel/Q+ElzpAuVduUUo6b8pWU1mPFwGc5uHr4OIbCH3wqvsAsZEMZ0rYc6oVW
VijM94ObBz5Fz+DTd1EOw+6eZjRksqcpKdHzprDccHI7hrXw5C0QVE5TWwUt
vw1ejs2jrB2x23Ae3SiEt5wdxJDW/cDxU+kKCNdp5KU9mtPDDjO+gKJzFn4h
JmD/lJRVc1X+DvLEmO2+lia9oXeoFjz5S1rXR37ItayKO09SZpOA6vRuwKQK
RU2TcO08Sd+1XFPJD6VWgzjpUVl7u7clVh3UtPb80F8zSzD90IQztG2sBugq
alxOhVygUns4NQdZvwE4y2NPlWSyfqVQgApY/K1zzSa1Ff0GwkYOWmq35oKH
uXXkgoZ+5IHT3bH2TQWyFOUE7BHg2o6EC8nyCOKhPDV5BBZTmAzqQBLO0gut
Y/kieMjNh5SwZCTTxt2GVH9NVsmGwm4ZE++vaVHCXjRUx5mwaqpKFoINk5KK
4IKLO0H3kHS/il3P+kwiU7dxMy4PX8e16rkRmyzUVPMNttmbD/b8ZYCDgIgW
7CJd9dT+oQ9nNlGj5oBYvSSOyh5XYLapbz3tHb63NED9HzoH1KkkFKimw56w
jHHQ+rDy48rfqpQ/ux8QrUgpo9IEhhw3B7weYb2Sq4l0WpFcvlBkPO9U9bH6
U4qltt7Wcv7SkFygVZjpodOCwFbdHjCicdLhauyKQKJ0pMcPFtA1T/ekBKFV
cBRDis4R6jv+sOKtdCr3LtpWEsBc0VYREQO2ogOI2FlJZViEX2BrODae2cVi
3oj2T+W1Rydzixgh52rSxxC0OiOeYQYdjJUxIqfIA2HnZooDZnPfiNbwoSFA
zQpCzoSzE6aQ+uC6R1xRbVWcU8dd7xVSWNkrdajC6yJffKI2UgMAU7wwWGso
RwJ79yejoqrRmdr5X7XNQ0I3/PSJjgvBN+9mGILCS815dxnqdPJWA+QL0xnt
p5FoxnZ5iDll07tNzuOQfKT1U8qEdRDufPWE8T/aECPYckuEcTtJApt0Y1cH
h9GfWXtBVfhP7LexxxrlSY7YsPuktGxUxaHIrqglkCq9s2Bl8qG2XETEBq9C
NgqTxvDXCFdE4ErbOSxqodCG7GoLrq7j4QgjlTsSxvET2iWzYDIF+mDc5VaY
H1CCNkfrbgX6j6i9if6Y/QdJj3ZIekeGKIlDlUkp8keTrykA6qPgjbUfM0r3
aoT246ljZvtECSx7jj+OtLi1YyT5ByyRzQe7ZkQcKJ2FRvi0Q4+oDP7Vom+S
/69+PzTZaPIAQdOHcc9jzjPNDZhCnRzDU/PbHDfZvdRk8yiZTvEQXi2vmGS8
fuEn3cjFNKWvRXM+XDmke0jE7PX44WL8d7KeR/i5doG4h8bgxew649e/j9Fa
0VBG7HV2swBiYnS4mlHvHuKIcRTaPJhayUYdghXQsOntrQ2ErkmPEZ42nbeV
6hyxydQ23Oli3qIN4bdVMSHcM56DWVdArtgzKCMpGz652Bi7+BDlud7seYt5
PQGgzIKoTr5A7lTDmi0j/h7F2TLbZRkPnaECrYo+SR/RTFyaugQ/0drZ/psj
NiTIk/o79fFKRocF9BpZULZK1iRuBEmZGsiZcCesZ1/3NSqXw+ob+GwHN1Ph
/p67u/V0P1dr0FCiwVutFT1aS3drvuLib8zn/jFmQewgKid2mZ34+ZtUfds0
ezNV8nZ1JNe9TIVcEpKXpN2ReHVbg4hVYsJuh07Z2pb3Bf58GlxH1kzc6ZZ9
wp3vY+OsWEEopN/u1c9Iiry+A+U4IUAL8205nXx1wwj4zluNXNpJYyt2CBAm
yllHIcXrAhKbGXVUAaryIFA3qDQtGkG7FCxbkJbIjFNtx3ayXBlhWYkHJgHr
QyegYon1EUOFrcB04SYzxSKZcqTHyZJrkESL6vJopCMg6DdHBl+Hs025z9yQ
6szZCwUiZ98lfvAUI/Ry6wj+pvmlwd8iY7ETIkTEIwQ7e483aLLL2eUlgNKo
r88vdZoKM8TcIv8tgqne8Zhmwp29QWT2KV0zt9izFo/DEUgilaRQwTdmq7P3
pcx88EVxSyMB+2o0FLrLCCxjZu3TbhDfTMQ/mgV/btg+jy+ntKjHKp8Ao6AF
mwYV4rQ1Q60c4Zv1NEso3uTS+i4DYTCWnshD+6BNgef+F7puSy8h04uEaJI5
He2JXIX1BZjklRLphyK1Cme+tJiu0ZqNM+SLYuvNzdTFkmmIGValdxpcJ6RQ
yrndYQYGJnAuIqcaarFKVwGgfhWP/xAdmxtjTZzQCfjIgY+9cdqyR/fZPXZ5
vNdzFYK2cEz89bQxR8TSF7D3ZfDUiBP8c3+5ZRpSCgFZxYccI6QpDU6W5PBb
Q0nZv7zRzrZIE0p40hHy4skNX0cyG/+qgIKJoUyZyqiDvF+F6nfanreG9idv
1MnKyIA0TvBEO81nVWo131VsjnPjDEWMuspvUEFdcOlFbbF0rYOO3V/6kESn
9Acg4ELEtsvHQnMcsnRpqmYSZ5lMQBTthBEyOPp4CrO8z1zME+rH/Nef+qyR
Ui0C9jo/riuRzV4lXjZdBdgchRCiTuju3NYLSyJ5Ug100SwxKGOdhBL1KlE9
+Z1ZXW/Z+r3QjGaL3hbu0wu0i+q7QelnxzF0IzDA9YA3ivAVArh2r8Ef8kgK
HWYWQ4GIdaTbLcosUXh1IBZhMjYiJFaE9+40D2tZzgHMrZMp3yfwPyAv6V6c
STXYl6XmDcMYA+RS1x3G/kJK8FNi+ibBzsruy8H/U5R7o9AZfgWZ9yR7OmlW
oXKW8nYXsntt+TSNH3OjNYdwZoOSbN2oBnGaa7V+e+5h1u0yFTmFqm4etVsY
10swRiTRVzNHxjb6i0KLU55l8/uTCL6YylqfIno++KmMzDfLZ+j9r5GS6yEb
Zqdo3xu0/UFLz8Qis6XCZssix46JPWSOCqegN4iKgxnk2unjfC2zcGjU/sWP
7R4L0dtLKtDC9aIakp3hW3ITdgRVufg7Zy4RsZqMMYn/5mBVraOovgWJATPI
nirfqVvB3C7OitDWQzhCoHMGiW6R5cIaFWNhnWBGU0066pbjZQUAx85kSqAN
tz0FvzAZoVpVva4KHMbLS1PWMxRPVD04dAB0/oPGXkK1Tij4O3xLNNg20udK
LAleCgN7Sz4yNH/Tj+o31m97OCvSTvYAb6Spech5AGl++0MA50O6xyxRxgHP
yjDjz1uK1rIAqHq5dCVqSxzLUlN62ICD+6/smemDHB1XFse/B0OHeV7pkyJM
4JamEokH5ZSrHJIr7x29QhiXpoUFLNh+OmeKxxdvg0pdgdkzMKvmip8tD2nD
57VUzY4NdwaxakExWENoEj3Rd/FEcKvu1FrIa1QDnuuRUENytDAiAGPS08i9
A/MXcZo2rd2lBS7xeRmPDtKWAI07hD/Osb8yO6YzB0Wzcvv9pUi9JSck7TQa
d8D6k6/3xPdb0KpB7QTms0KMPVxHFXRKdo1H1Vp9e9GnbSCGz+uJQM1emKwY
ch0pE5xnVUqRv2vIN0G5UgUwDlR5IRdPksDZAerePfAKR/JdN6eowFeHRiIU
DD4saren91HnzMS/VA+NxKTKVNvw2bLnDXUH2ehx3ksiRuKB4JASAOqQReJj
R1w4iXFV1k5ENK6Q55R5SVtxzWO1b/ivdsxdn8hQJbmCC1GUWVAW0KjSz3EE
QbNBcgx03Gm95vP6Vj0juCUJbYRKcRohoi/Qx70kYf5uEKVuIM9j+aRmM9VV
pQCAoe8d0hzZeFZ3YiRTKEVPy3uddkJ2Rjn0XmKerEot/8DFQncsSgnxfjGu
dZ/ctXnKScL+w0BtI5FVJptizkNcxzKjYxSP9wMY0lD72qrWl5DdLZE4M0wS
qU7gfyAohmLRXPkygj8ETjhbv0PL+AYe6RFTuMtdYAVvARpQq11l/Xw9WnMy
sIM20LWP+Mthc+/W/3ogFt5Fioz/cxOSE7G/ZrrSDOSKypsOdVV77yUM6MaA
UwIZcB3igKFQB6SMYsbs73qh6+ZIclBz2ZZKCQBco3JRLbcfpBSUMe394Fd4
In4gVzKV1eb7IPfrUJAFf10F2eWbsjOmIDCbfbCKdgoKBZxofQuo8qGFR6ll
hUCuZu+n9FPpFtlfZWYkcrJOYEesiC7e7zfStK3onSne+qXdXNTqft08lJOA
hbPPgvAlVwBkMZjoNrYfo5/VYLLcCmTNMclbuADG8h1azm6/uQeoTI0oS0fL
bJTfxsAS7NEPgQ22rWT62ACZvVAbgNYCWIoQX92FEzLKCZYFwj+6f333wYXk
TcbpMAuz1TJOphLi9LoKSqH1Kt/7kPveiBhphjjgHhUDvL2d4OlDyQqJWE/C
ns7Jrk5e/KbYSgKYDattFSnV3R/33tMK7ydrA7PLnt11iWG1xkkSTmVGg00X
li7+4bFsDUI+W0E3uDmi8sduNpmPD486r7XX5ml8evy/gpsfxkMMt5Baf9ez
fUCfPhYBjc0Ti83/7JdsCVD5dBxFU6Lhj083bMhIejFZwlD+TxgIyaKMlQt8
Fc+LRsNMWrwVbaaVhnel8W/DW0C2FbGOEzoGd9IbrERvYUbOdfi7A7h01b5c
w0HhhnHpzAQaYxm6+rkI5jMjl7Wti6rpxwlUjJk+IL15oGCAcMNiFky4x84M
opU1BEDsrVlSpKm8MWvJlO+KXArigf0ktx3KnVSP9wg3W+aTdsIw2KFZtMQ0
khdkPOn/xyIvXQTjBS7J4mEk+BmevQl88xlbeGBeNjkRt1nr39I5ZMj18OEM
8N4oLoLQD5sP74tY/ZyIqP74D39TicRs6hC9P7f61+dcX8/QZBJBsubb4C6+
ljzjvFpAb482J5JmTV9wa19OmFwkp7QIrQIe8AZLkW3Q9mdst32Bsl7c7hpd
So2R45Ou/B80jCmsOl36uclWaNCQkybngddVufQN1cp2NnnbnJdSsk8qiIgv
n6+yp2LVfb6iJqQ8txrUa8FqtzcZ29RSfcGsrvuoS8NluB4TK5hUHlxevcdt
+bKGv9RgnGJ8JmveWgfR+VPR9sz1XF/eo8amH5RnOT+pG5kS6vBuHaDidMd4
cCyuuj4X5lXT3VnrmVPUXIB0piV59E20O58S1BtRBXYeVga3Ge/qolKYPuPC
rf+usP2htjWqBFNgA3z239p4zghjhOzK8fcgD2wXlTHo7Vc0fayO6OMxGYBR
VsaUgiHZzMbU/1w1grYrcXtjXvHE/lREW1x5TzzrxVMTF0RNJ4L/vxBkbiBU
k9Th8XqwjOL/Z7Lm39aeaF8p0tJUY6MO3e0ynkLmRNKfN+Tig9DZ9IZlsw1S
M7rks3KFPPCYkjjM/0ZxdhJtNowUYqfXHI0MAk4xCy/3E0GveciGRak+Rul2
5wP4hhFctD2UJzUlaOIcYJUPJpDoGMQtvltmV1t7XBXjOWSRHGimEBNWzoyC
Fg9lJqzP8k+lUe+7fxKR3d4Fr+eFV1LOpLkY1BTchIL1b1T3LkZzAvzABy4m
3EnOg3np3j7tXHqAXODMXQ57JzVUcuMeBCXeBOl2exf3732PLwn2ED/mhuDv
jyJI99yaaq/dZIuwq+yExe1xcwfdrZmEbVYtkyk+A3Ob+8xldp91w6Top7AP
3X36uqN95H2uZSh/nxWzw9nuM2MCyhKgWLGhvJaSlVLcnjw1KXibnOPlgy4Z
7udfynFlDbcNqflaxHZ6IyjGCJ31wKvvts+Mi9zk707iSbAbBY5KYu61WTRy
2P5ABsANuow3am0THx3aIXRlESfaZkp2YBdxnelIjgc7Bn0Qmak61nVNdzuC
SYXUXYz3q1tDQTgMqRy3sQQl0w9D07g+HzGJkHIdcvOLy7X8Ke52dWoTtyCn
2tRaWCVCby8UMKiAnA7zi2uVuasFCAz3Nc6SkkBQZmeGsDWRLYSbzKdEizkI
m094S8o+XHBjiNJMkP0cutiaosWNZkzQJvr0gAJ+pJGBDac+fpIsQYcWn9mE
GEThJm1zpM9V7B2BDEmmNSwh8JK3LmcYl4KM812aAO6q9Vv9SgnELJfRDRJR
c5aVy4Mn+3kE24MEMWg7ZDOHxu89w4XMTAoDrjL3mHKFNotrbvCBIMUB8ADD
B8MOqTNVWWtVYvoZEoMkePgcbn3NpoXbd12nyXacBFQNLoz1JFIcopfyOdVJ
fTqBQSzyYVNJQoSZxc2vbepBofGAUNzkz0UrkkkbuKuDFMNvib+NcfCn8iud
/8fO2EpGOLqgNKM4YMAObIXv5ADzmk2kO5cQ4h+FHCMkdyuml/rL7rng5/hf
gBBvETi+XegJzxzMr0XYfAFasx+zbwWPfqbp0o4EUoNpR3+O5HH6AEl8Cbue
p8Zg3TIheWdYw9S321JHZfqPjyctcRjxPYW3cysIWzvfAsS/jMywRQ2lKFip
u+f1TMGoGjnXlYHbENsRz0rRx3cP7egAR4nH7RaGMQ0qSOBaUW5bQHQXj4+K
Z7YCTZM1C2Xk6rDLUXVQOgoZFeYAezI1/c2E598W015jQLHFwSAIYdRDuxSj
w4ylk/P/C03M4MsHkzmwsjW1VWjmB1lxyr5kT0lwTluwMcww7Qox67ncvTjh
iqyyOSqdQol109PnFI5yiLqT/L5bKqJ/Y0hZGG1XcEqr/INLWW9wdY3yGTjo
QYYriOQ2gjz3LADRD5G7GEsy8KJqIF3RR3oEPVilCBqHUz9k0caiKS+45WZB
G+2UlkBx5FF0/2F77+eouOaSjng9Z0VOG7aMNTXKKPBQYnCj6OVFxtQOuuIP
XPnvA2an2MlquvO+Q6MQf58nasAPzXDgidXYggITDOgyCtiVe8dt/U/xiPiF
TQXSrw0yoAcQTAe/JITHXWoCyb8Qky1vze/TYos8iTIMTkOytZ3S9NTcc4zb
hQgD+Kq2xEfSYE1S5V22e6dMvO7JYimQASdxGA38wnR5675mxR5OlBfxtdFi
qe+L3ZSnZYaLNc6e6ue85Jq7LbpXsuu8sxNLs0aXUSxKdu4Rk9uu61pmvAeZ
zi4cAdFR/ig0n9uGRGDOvoV6MIK6WyfaksLt2G+2VX3mX3JJC7IbxMNpQ7d9
OSSu7XXzapZ1yaqpxPlxgJyMQz93Lth4i6rmYjptpUElLFfOGklURzPwax8j
ec1N6brz9hrxdsHU8AapL4dChND2QdtURrYuN8I44XoPFTeCNzseoI4cVLw3
aXtNoQYkxjzLIiBx69mDiFxwPi5n5YQWxpYkWK9aOs5KAtoe6Amsk9C409Dt
ucy1rfHntWUKiAmWVXViumrX1+J5fiEocCHK0Q1oePpRWLAvnIdD1Wmnl3ZU
TeBmLjxMLsjncom4xFlHyogX1u8hZFmkxcMyXy834V6+9dFnxJI38oOLDXIT
FUVtNu8RPU9v6TZh+pfGGUpABgfknUkRSuqvmftOEAA5MH/0w2y74RQwjECd
26a82ypii921mPRXt5zg/JB1jAxCTqxpCBBCRpJAoUVZ9JJFZqp25Fl0l6uR
FZtXhObysuD7sDl0pAelIdCbVTqiNAZnWTsV4/8VoTKEX63gc/bRcDFdHJ4T
MlvLsaEUbOREmhMo4Tj4LpXj/QEU8Y6cl5OAoTn17On7p9YduIrAIAuzQ2eT
8dPWJc5QddSLof40BqYF5BX205ey/SmSYyweBLM3Int5l9D+wNHOgVzHcVce
jFqc9+uX7XjXP++zS6jupsuBwadYkUIhdLHtvNr9JbDWB0jbRXTjIz526thO
YCbhnij+yi/MVsJFloGvwO2z6C+58nKb0BJMfsPrqmj5kfV0k0YS2kPEL1+8
FmhSfXrFTNqq4I0yPaD4s8tOgfpJeHIZuCMH0V8CIREkZdvjB4nMiSyapeKZ
d27pGOSEMAWbq7axSC6fsTY7auu+rvDqmk7EqDr4BpTn8dtIPQQtnkSwSMRl
Omh3Aw2o4xhRCS2uKuT5mqxUubiZ150b36+Qzy1afkR9uOzWzTABuG2wdIo7
wYYyL0qBmWHEwt11FKPfyHWnA6D7BQbuHZ92VsJE/gByIuUwxpS1ijyfZ4TT
uLU72/L8yK3pQij03GHZjIeZA4ZrRLCSUNkEz09mw2rPWhQeaF/HnWNp2IUC
87cq7vvBNA8wQOnWSdDbiRDhVUYpPlqY+jPmf+MBlU6eBTuKPxAQ1+h9+EB/
0+AFOWi4miZB7xmS7tO5oL60JpyfV5R0iD4Sy7MjnWFU7hOgLkfi4POSooGO
SiA3a0PLqbWi0DHNNLOLKaz5zcIjYO3/KFSGAKm02e/qvkBBCvueBPw5g4cW
7GS4TzZd8RxYjN7uKCE8OOezbHDF1DW6Gv6hYH1qjxqVsSZ17Xaxfrz9FraS
7S5qtfurx7xVDTNfOickBpTpDk/Oxsy6zuqp8n8ijhruI5Xu+XXHEjLG4qHd
hSQ71yIRlxCIn8SMkiujXzoRJ8GIPv6Lz0mkNFGvmslUVBnn+vWa3NI/Ir45
nhxmApKvJreVJNLRcaeyzAoqm8aikOO0OQ5sYAYNsAUx97vkSmEeo+bRMKMj
oN83svkoH2iuosHzjEZ6r48tQqGoxcAyi6+zysCBXegfnns4E53clSwBSzDw
LaEPBPvqkeFPWrLZQoa396soOi2ZA0hSFLxuqFIZ2s/d2GfW5bOGJNwjl6TZ
/RkCLiU13AyTCvOKJWc2z+J2LkSnlJKe8WrPkq6D6lZxTEcK8vqV8DH51TZA
/pF7y8EZBoZBoutxVwQHee/JXK8A4XAKlbasyWq0luloHxJ+6tCVHLYgZxqO
vE9ic/cgDjZ5lKD7NSSOb3O15zA/uORNxrxvEE0oqo4JObId2Wbid0xR2WZd
23qGcu83wFEPfw2ir06dTlQJ9psTIsHxs+b9ptLC5cT4cQOJrjZ/P3AZ8kho
KKR4e+rRCZuog7SZO0G7CzMlpjK8tag9Mql9BbXn/y9lLVFZhTDGmGw2xNQ4
Z1FfZJOXAdDU232AiBU2AkOuNZxOuwwDwCutccZ1+Hcp4MNvaj/XMjZ/NcWq
6w7k9fd7RLgeV2Q+2BW1rp9aM/UAfjuX7kaKGCZqzd1sF7p9BJeifi7YE6pl
gtnZ7FWaE1vesUt9O/mOmMQrqBveD5rPuB3uFSP0h0OIP/YZUFpovZBwPopA
TqCVNxR05ubMYQAdBHdWUNouJPDIiv7bP0JNXYBjOKswrAG3mEdHay+xFnuk
L2ORHld0IQCZToiWP2/ig0KUSW3reCuNQ/r/3aFGspxgwZ6a+yPzzWvm+rBM
PtXlXaXnPr1FMGkW9GMWyzZ8aRuRQQcZh4Q8JoRYEcRK4OhaG57K2YVSlczO
aC/YtyMMDvTp6AVYhdk9f5Zc8RC/Am3jJK9bypY6+HQIxzvYomKscK0XkKkn
mc86yFDyy6WpX2y8mvXN72DvgXXXRY18Q2BTruyBosco8JQYkAKwipag9Y86
Qb0hdJo5IpEOQRkS7VrEojI/WHIb+OwEDINe2Yp8z68C+RO08ujeE5C2iN1p
1pPgwdgP+oq+0BpIILv+Uc2fnaDc7ce+tf9YC+z8kfky90frEBC4lz5elwSR
1+s7R/75k09eVXx04cp1qNP4DiRdaQW/Vc8d1i5rbAbn1btPidzwUbWWjo+5
m1cUGnlN3JjyqSmAvwQhPJP/39I3zHWVem1oQX4fGjtaUksJtm/4fZ/mMfHk
gmjkOMdJ9P/5KXotdyXFEQ0KcMw4w5/pjlzYonsJQuO8S/yehsDMuGASU89H
vEzWibONoiL7+ZnF8VZ/Jz5KnNHRomuptnmkcHaF/HoND314QTykkUGvNiev
SpXQIgCSZgj4IyEbIbTTM9+tNRVOoD+wgRmaYPjUTQ1JNB++TOFF8LhkrEyx
LzjUFeIrp70DwsAXICPVUnQ8dwFqq/QgqvhKFsxdH/Sd5ZzyeLRQpPGnKyjr
5AGHf2snPz2dC4nePYufJPteFL21+oKovpf9t77eDPo9RTPubYBwf1Q/UtSV
CVX6ZUAXn/0Ur6KIVkt+liZcZiqyhW/Q7NqMSV3s1yUwBPUPnYCHnWQIztrg
rs2okhYOBnB3iuWWtls8GDk/20bYvFtMXW/F3DYz4vRBoUI2aHhk+tuXxnaL
zCTyT4mpiGDtTFgXcn8d8/V0rdI8GgA7Fn56dV7aqLm1vbwNI2nxFxmRcW1j
KWQNRYaDx1c/3s4ro1Hm7AdhrzK9SB8tAK8peiZ7gPgPQb/R1xWqI238FyH0
oEh0LyY1Fi1hQuyVfxH2QSsZ1p1CMf5FeKfCM6deUhnppPYeZO3wv4JvtCZp
Phm5KbPVimoxNe7YFo75eueU0sd8gsr8K4clw97+uaBSZZs0eMPnvcdTlZth
tCStY9rN3mcvycfyQKR4UT6HD+psfkzYDOalSvMp+abVF/cJ7siVrG22S8T0
5zox2uBAB7zgiGTF9eAMTAyWE2fHilwPzH3GC8OGXsW0NT6TfXBWmT8asGwc
IzhMp+5rhqb9AHNEhwufmS853wOOHc1Eihg64Mf57dwn5Sjy2j6IH597P4EO
Y0QT2Ev6nA1V+zHATiLdcUbsbp1qa1aiB97MTjDOmTnZxsnmrzOE3h+dlaxC
q6xLjb+sm/HoieCKjijnZFXMoWFhICtM/d30sbJGUPSbnW8NkuIpl+a8ZamX
VkVWCS40NgYlNkoD6GCNl+mj1mAa0ptQh/ea0p5v+ii7+NzcwmkBQdlp95Yl
+UNkT4Cw4n1DfMPneP0bkXpbhzKkucIiXH/TLrO0pwFnb2PMZaxgsu/W3lZT
VjLssDhtLqpUXpRpmlnRNAuohlrBhUEWH5uiBwC+1YUmXKjbEd/rDCRwbrPc
/S2PnlnyhpEEEvS+D8y2h2zaLC8yq+cxC4IgiUjzl+cfRQA47JRrUXyN0vLu
AuNPC6jSQkk4es4o0+TpbN8oYVI6cqdHc20ajRYTpKyiBmDZrSa+XOfke45K
YCOKzk4q9j3McxJsheRfSFpEgfr6V8unsEa3RxyLeBIyOaOvgz7loIhf+ozy
BmouLQWA4Xkvn7T+8eQyF1R1hDHDZ5n+iT0/dHDdeijRnnCu6ye5DfvmySA/
rt/J96djgIpRfDCLmIP5iloyZfq8uV7g+DU6JfM88r8VtHT2BQw0UoaOKSU9
MX79Zp6jsc0rwnrSNARJpe49cUeCaRrBbeFd3GaqNNXrTWj7nlOyPrcbRro1
v5le4VkJaii1HJDN88ZKPDS7nos8k621HsVA3ZckbCvY2jPoY2ZIeFkYTJnd
HVa2w9K1IO7gHZIf3NqwmVX1XCu7WhNPGwTz8D7rC1/ggHS2HTgwrbpUcrT7
iZwRZNidG0wr5eFuNd7DHdaESNheeA4Qk8oP636I189mK9MlSRo4VVzW0e4a
dfZJuMq7WQ/AVwauvSnlgDNfhfX05bzWg8efXRk3OvGMwt7GdkDLtVqMzKp3
ZfiYQfvn1rIhii+QOx23pOmsnGn8ERAMlTQZVoSFjbrXcTUZpvfuF5sVe1RL
kX4Wbn0G/jEQpVkKy7b5xaKgJwg3PxQu/tlC5RxJ/OiADPUwLophK8UpEuzc
Iy/i9IG7kbwg3/KY0gL9F3qeNvShA4xwI7q4ek5TzGL4rfel86wpiDQA69/Y
AWxe1dLAka8FepXtOspvM8+o8G6YFUbWvYNT5xNhMSallK4yamHqmLx1sZNK
tupeUC2VAtY/XDMB4dW2d+zbb7niPodXHj+CNLa2F+DmzQ/E6+zQ5nGtbo4o
1OYExj/EUydVyq1ccYKbq1D8fnTlxoYP+vNkz9Xamw4uc3WHhbkuDbFaGOOl
WCuRE7qjJ+Q94d/VPICokDqVG1AmFhdZHwXUjTqEkqrua3mTdAAGJhfMvZtO
/oSefT5pigmTBWO2zXoXhqohQGnZWLouvpWtu5wouC6juE3cg1Lfwp/c25AI
1XNEk2EJHIEGb4TAJ9Lx8UqhrkXlSOlxoMqj97OBarykrlwh9f1vIPy5p+RL
v9nI3htKNqiNBap0AW9sKoLMkPGBfWNzfg0NZRmwUMiyAvcTwUvNX9NiPfMx
PTKW6XcABdwvN8WiOMty5roEqXEN7mVGNELxVGneOkGgYp586LuLqGJOQbFN
XG43LJWUrsap+nBTuqs0ED2JY//jR3un+MkcafiL0w3VchYxJ2Ggec4iaGYG
PShScU2vpeo39Vb3otws8h0euJkT+rapKNvwCSUnq4COw+HYEOb3fqGwAiVD
zCq8Gwh3FdVdaXLmJOd58Ec+B8ZemTlXOWlXS+hCWVkdIKIZ3TIEv2FYJfip
sZ72i2XaKdRySO/7ODQZ0E3FGJqlX7A/vySqdgtMh14GHHHtTRvGdh5cHV5p
9dLV2l9DqHq/DeQ+srUllQabZyS8aZc9/+hsC3fVU/HuiVhtdWMysx5PwPj1
/RGJKlUNA+CHWiQUmZG9F919CcFrwoET1gi/+D5P1f//Tq4ebMYTH+RYygSx
5My/5hIvLBs0SXSvKz7FF17/P0qQtFB+VNcCHgS5Fpeqt9VH4c4r2B+N9C/n
mMff1UK83QWNjn/WLBVS3zLt5KyotBMfMQQBcyc222FwteQ5ww+6nKpe+2nw
rU67zMWxiyWXWls4Rr0IZVO2IfumOea5jj/f/CbjAYkll4b7g6WmMsiYzN6f
bv0/7AAzvnamkUbgXaVJ5GMz2rLf43adAKbseaP/lzYbAOXyoUhIZyMJgJRH
OmyZE9/YZ0dYoJz1JWVy+SKOijvuvGSPgzgl8MV81zA5HPo5B3Un+wKI0Dqo
RlIOhNZwjfRle8L42fO5eIdRJB5eLNvyTR2Hd5L1u4OKK6/1eJcHEOzHJTeu
fPvzdqeWK78Dp2kECMtkBgNXtjaea8kV1Z1IePQ2kV6dYsU4nhmZSCGA2fsV
YJGXz2n2C1UI2lXvZz2bi0JV1kloAlbBNfsMjj5h7h4B/8E2GtAwP/r5dYXC
lh/prINGk3g5f5sogyqMd+xNHsoGmEPblwelh7h85AZOajr2wFB2rDtbSf94
rRnALwQuPTYwvOfSRmJoch0S8ACmA+4H1EUCcpxUkxxB767kPfzJSKWihluN
LI2Qnlzu/HMN/6ZqsslZubFE8jkEfrZg6xuOR1W0RcrwZtrVRZl3V4rDBlYV
U2EXG7rCio6c9NswNKyEwHwm0kgsvwT9I07ak6JXJSVRJcD1j2mYNKYL+lT9
tRr2yIyn7IRvYvvuzaZPc1WjWeJcPOxhortCmBiHIQBFoim0UnBWKJpja4De
2SdbOAfn+XWtq1yhAB/H6QXEWIaLcDx1QXc6jaqGg9ix0TxR2yfBooSzo1jg
4fp1UzYyGDqN76UWx3XTeAehRxzoJ19/FblUcBsYYvHue2t55BMUT4L3/2ee
c9GgJGd07xpk17fRyX0SHkbDB3tGfvK/mDrSS1y6B12/PmSB5IkRgrRJg/ZJ
F8BE9NKpaJudmFKgPDslvxQEdHS7sCaHsBw2i5VOTvaSzJ/u5NcMM5mOHccT
tq7YZOoF2RO8flvu8yK944TcYba/ZpRSumseDbUzzZNq3JKr3d9Q+PWYCTjl
iztsRJxt/env8G/3Zj+wFY6lT/FlNFC5vMQbKBud2Cph7qPAFjOYqyQJlg7S
vIG2yLyy+Fp6EsNn9mNAXXc5GSUjJ1y/wLSkKCqGZG3+OsqrPDZFCPm2cz/G
bDWIokO1xGIx6YMBS1DNaPh9auqWN/X2g/JIWVXAY+Ecs59fV9CfU9l3KdJJ
9lrbeUiP+Rb/BAWHqzthwpVdVUOJzvVJWiNJJdjnvXi21GxopurOyI24JSGT
shPp5QOWCoGrSKo2CKX3x7ibTHRSkZW0b1z+LGk/LzpAu1T1eNk3mleR+yQo
CiilV0Uas3lhzQBG/RLi6Aw4yiBMSAj8o981t7pDII5cWc+l8uESvREebAXJ
QB0z83Fz//5abCze3hf8QSnuAEhqQpNE0kvnmbtvMuyTntBFRbOx7uRuUL3W
SG6TdfkPZhNYDfG9u/iuV+WfdfCLQi9bj17jb1wzvPuMYxhqQenLN+rVH/rs
+h4tuQllMRmbZycSa6BUfUk9lj5akc6qJGhW38wzDLTe2GlRYElJYLzKaoGT
hgype+84er4l5HjpRfEQyu2jCBjMENIy5XNYUKw/5grNmTtgQftDyoh4UJvZ
zhbD9ZKhI4AAjESNRJvYVaKZz/rgqljY6bMUGpfWF1Ncc0I6PiN5+J4OKcFP
BGJpfySBn4Bim0P6IU/xLOWjWkVCHYD1NlISvneuHjv9aV5JBtlS+XeyzRhE
SQ4Kd/nFCJdPYZNFBvazQZCSZdxhNn0sp5MU1+0Vz+bYmw2MpElu8Z3fPAGW
hRZuliTQ6upF903JtGjhlO2Imud/WTWDeMcLA/s1eJRJdF0j/T0JWVxzgIs7
QncgohLyDyi9zEcJcCUMCYd8JiIf3AbTzbj6DzipsI2pMx8I0hS3iWcXZyA5
m3gVhxgmDHz7D5cdAQZyHi1LH4ovPIpdrNAfQarehzwJvbByPRnhBn9K14EV
1732FtDV3Wgmov4xaRkxuUmY4kVQOQ51QLxbDIp2+T9ooR3zsgHZ1UYyB8mJ
nZfkImxt2BLO1TlrL8TDV+NxUkVNhQDapqS8lmhWxuepER+SwJlK3JPAC3Kv
dG7oZ3ti8p7CHiJ+vtIPWA5U3gwlBKnPyZCd5R6iHsRsXcFlQqIjCtn+N7gS
acFuMLLo7aJQM503uXzAgO26t3xLUOYe+R0eSDkJEZMmDtVcxQgKg3d66aAN
b1cXJhmNGNHZ8xSjZemSbehrNPgSMesiEkJgI92g0jaahsfYOUloEQ3qkbaP
bfjmawbZVuzR/uuWR+mPsRSfx4YxqNhZ0oTO0Bj+jGGRvFHPmDRLlD3EUdqP
cYgZn1W54fyjHLfF1Tj8sXdjYF1a1p6S4jXDXfIOBpGg46MabnDV4SICgv9I
oYaxJcxG5QT4hxjbbdgkdeWbTO6svTpVkdOpJQKTHaPA0i6XJODolgGWhwJX
5onE1H9UtglVmitbmI1w9r87ad4LGYZ0AVLrbubHcvhiojzWyIB/r72AWg81
D1s6pZuQDPr2GF27UdEffj+2UVzWwNZ9fDThN+I78GseNbQPnygJTw2Ue8Mb
1ZhgrgRYohWeze1TgrnybaxGmWxC/tzCugvokCctr7AUgKR6KMeJEHazuD8a
UkQpoQfAvsJ6Lif2ibNUtZD5h3FK5wpLTFJm/aVv7WqB5+r0PCN/HE5NRvdw
g9LjfRZQEBalHbRZnicrk6ommRrB3Xfho9nCVSVrLu7ZORDgji8r6Gq91wb6
Fz+J+dOWeRR/5Nm/LEA0CMic6etl8cllRrSZ32Ij82vzhvEkfTkErenn3WUD
KZtrEVcLQlxyfH5ah+A5B+iuY+BFPgyuL42fnfg1fOl4Tl9Txsfqw7NRr472
EIhd+AXGMfxPANTqNhO79DjbLV0YxLxymlbpHDtQTe9p9I5TXdZdFCrgcXrm
wd4NQbWWg4qGSpPXrxEf+OSaCHsNNwc8d//tnAPlcy2JbzjTLBpceJZ9OTDB
PDiMstAHydtPzci0+w2NkcfMmrAsNNBKPBWKhPP6h4aZXJ3vKu/irGRw2OhD
Efyni7MSw4FKe6HkfZ+zeyMdezOb807yaMU3ITYC0k+ow6xFjtynwBdEmoXd
pgIpiKfbqaSNlZWFCfYpXUNT+x2IgzRDHTXp61dVFyne2PbDFcNNLoixSxoO
CWZWFZh8nalXpkBFS34eSAyhhPTrQvEENOT0P2Og89mNFWDFQme1ACa6Q+lk
bTADKvliYbArQ/m39WSmzvEX6GEdODBP93J2Bx2zm4VsNwR3Wab95kMz9Zr0
VILLyFfIyUIsgy27kp4D5NjD+4MCJl6cOqSqp/MAShmgux0EWz4DzBgJbQZ0
7Fa5RifOcuZ+q6GumD9JH3RXeKkkYaBikU/P8BiB/xi6u6QR90j2kMfQfKdm
dHBdO1ddNagyjZPqvqcG+39yc62RuMAT6KqpaZFMCSHjATSCLI703hFe6eia
AFvwsGNWVjVB9TTFwkuB7xfLcFiKTezglPco8728g3uMpTgRvB1C+lss39EO
+p3unYglQKcICklQ4Wk9vYoLP8QTerMIT2lZibdlCjTZnADubqCbFDTTJcvG
ii2DowMo5zhidvLV7vnpsf3BWmj6AvsCwpvLYL8pQu2if9QjDZCwBKPoAxL7
QKSDYZVy+q9nYdcQc9fAy5aUxVFwmIVKCHK3SJuEUpfC1Jf1Z+9oqikJWccS
YJ2nvWUvMzQkY0Bu1M3OGDT4Nscnf3EyZwOGPKTlacw8rRFBgLmULfh4KiD2
b6XHQYmFPccFtNGqKUplveZDCPKJNRbp+aIVpRCKgk7xgXYfT7GNjX0Dmph3
Em6sfFpM6aRy19Ke0gGnN+K7Qg6m7f4EDF6zGhFjYcYwaaRkvBFKlzpy30LJ
Xp76Oyvt5/1zWUbiqTQLhi4fQZ3sLhmC9QXDhWelEkScl0QxiINQnAYKY61x
IJ/hSYPzk6ADBT4YSTLlvuWFM3FFNdnviHqaPPY2yZBsM0iqdPOAgc464dai
owz30CcG7sAv4hdicaSjerLA57VwPWPUrN5d9cFEA7Gozbz550mu4lrTRhKQ
NMKdMGDmU+MHsyXsHYdwHJY3ykxtdNdYb5vGNi8KpxgkFtOjpBUtZocwUGCI
zwejU1imFBvA6dl2hIFZ+ozFHsxrxTJJMMw4PA+9x/otbAKrjTlB3yrujP9F
IjeTVKvdq+GBuYF1b1ShqSe43BpQbgJ5JTk3fmV0D4NZEBjs7QX/6gXQfGRS
vgK/PcyzhF8BzGg3FrprQpASmVp6cceRMOnxLGYIUWFjPRMCP+RoWQNKEN+u
vOj8Pcdq+nM1amE7xct9Pgp1XKYLXiIkHXK0guXygKsDDlrP3LC/YK3vHp/L
3MC4WWwElHMuTUyfHCHb4u3ywuquU1wypNtaHwOeSCzvCOwZPLsppNuPyzsk
yD4ubz9Popl46f4wsoqRwLMl26sGg0JYqwrujsQcnzroQLOkZIO48eXu2aJ5
e0+aLcL/81hQAFGS9l2Ap0G9edHcmCol8W40g49GSmla3+CtzEelyuMSJFRC
pYNS4we7eCLAjA5Dc/BvGF+NWSEBC+DmkmC0UZ6/nn6JP1SvrldQDJpaWynb
k8yC6SVhiMH6vkcrykET0j1j7CJoxNAjoOMz1LewX4CKn9+QiiMk01aksWng
mwZ1F/Xqr7uHI34KCG8chBHub7AAhrA/tY9bBPvL1EayUPDyaL2NIvZi389e
0vK3IdJ3bDun03THbyA/6oaZgq9kLgKunn9z6XdSWiqLVs+s9DW5eoGyg17l
nhL3sRhw9jXWzw0czxAyTnpOLDd0f37z/bD2NL34SHQr6GCZOOx2ByT6t/ou
OvX1VPIn6HpK4XhGBbU4ap1qLRlazNOipkFICdGJITGyEO9725r8gnZZ8Gmf
a77c07EU9DGqfi12lspgvvBxzRaefIfsPnfCol3q7+t6U2+TncNsJUbkXVa+
BR4yGYixMZhAAX8E+FiE0ErBNWV7LISdGI3YMOorVvVd45RDjGKAti9AFp+S
Bp4FuRFLKsD6FgwTrH3iq+fIi+7tOYooeX8eWH21W9KAPBTOsUoZRa0Ge1Bq
T1o2N9Hi5so03Fir/Pc7e4Kq5gec0e66aBxXszWeSnyZEv5Bd9yDAQNgRX56
Mfh1Ka/4Q8KJ2NtALECvLiFAU9VEYSLaYR+NdR4yKgftD6atpQ8wQpmG0a7d
RaX2fLE8evDkyD6OWgo16R+2VJNKc68JhpMiTijO6xci+4SIul1Rvwgieibf
a1C6F1SXVn6R9yvK1Nv1rb3eN+uyHDjXbj2QAh7OWPrjfSZlPg9vfN0l+S8S
fxbZOK7p0m1uFe+m3KtJP6nuU5vURx41znmy0Z5liR4nA0GeJ0k8PAz78Y0l
WRxEXkRhfrKNuZ5Wn2BpvIbfmiBueITOegIOqv0NgETC6RBuPWjr3rqiyT9j
Y3yB7SEQJKaq4oEpq+/4BfSDJku2XpkhWPl5LZRvIVGi5GEMGiRxSeshZD3z
ZRMgHs0WmOPy0qJH/aghSfwlbaxBrz3yxWXFawKKMfbD5/2VKXt5NkopAyHC
bMdQ/so6LOT093PWG2nMPAOi8dg3q0Fm1hoXBuQyI8wy1qMHypdzxKeEccMD
1iqaDem3Nc3JrjOvGjEymiXHM1R+5rZNCceNLOQd0e7tGjPvs5XwTIDGS8JI
fpuBEIRwDY+COHxGvg3CmwIX80ovV93d8/TNYsiEqJyuYnnrAGeCofexoRoG
yyq7E7IaUrR0fRNxWH7xrAXJwrZVCOngb8VZE7al2iAqRcocFmV0H/3KhJSy
PzxlmiNyXw15wgV3WEY/q2HsM1r3KGtwHoteK/WlBfTKi7vtT8T00Dmin/pa
JfnP4sAptXL/uyPAfOVrfY8c2XQruq7KB82x1PPI3tdakn9a8reQcPRI2Gtc
KgXXlqQWHKwExo2bqF7WncjHFmAGIHFD8A0cqGmXj96uuUpKivKpTSm+NwZp
43H6gsUaDR2+Rm5imNqJTAJ2FdWCgKk2zIMst9lfbGdFh8XeHtLilOFvWkC7
wpU5183UmqgJtEqEIrdJb2DXFfmoVe2GGjLniOy7ifHJ4T+3PUQgWl7BlvBP
GinCzpzEVGRG/FC/ai5/RH/wBSuc17/yFd51YQNh/rhaJNDqTfxmtqtaos6b
3mumBXxUe+6PzX1SmhSDrefnY2Vwy+uPYa2dlBTBtgv65NfhAyBSkg3xuSmD
NyHTmHsccIarWEkcS68MC4bDuJy5RQVIUaQPVJT/tE7v3CzvEHIMazvl8ibF
Qg7PJAaf80rSxTPEOvWCPW9Bb90TI2XOEIvSPGaiMXl8w/Xmx4MV4cPq2pVT
t1WJR89YeewX7xjz/2STosNUETiSrLalpX30/p3pM4AOqwwia2GWL28znzOy
pVxmqdHewKry/QZFBEBWHTWbKw0UzWAEgmfRDlB0ZTo9x7fy9u4yN1D895Fq
SG07FkFiTN623EJ684ZtEf5yQlVmfWFw42wRv1K2zk5AuH/DSDdQZ5TeHYLc
kgFC0ndJ4ssqv4LdBTs5WqUlAKsS9JB9dfC5yt7RRhm3LSc19WEpb8TTNSG3
VnVEJUhVzUgvmZh6qfWToc4fRN77tL1SypMxhBcC+pUrjUSng4W9rQWnbaci
MY7QMjOEBQrRfRSjBOnIrpDRgSPe5uhPcoEY0N/4L3PwtVtcKz4Zf94WLDl/
LlhM/SmAPp1kNQZ2A77y+JQdz7OQdjX3CFhmrp+uiWPFKYFmuNslFzNS/T7j
oa7vzcqxxQlDVNL7XvQbBM8b09XXeIGPx0KP8MqUt4ZlyqQH1WJg6I29v4OL
mMqdfHqGENy89PLqDfLX61wRmu4fzPxc24f1o2Mxp9XbG+ghTogTTiwaPRQZ
g7TLoWbMIZD0k04zl71MGSJ5MGtIzlJ9FGThF7Gjm+KqP4ZdJZyBSW0X0P/l
Se3SyTAFL6xIviaNltVHmPW/2+1rdY9ATzy0kgHZfH/IavkMOjfB0+VkKF0u
NPCg7fPkgj0ceZFW4dND2YnNuxTxMf5xZdHktyIDlu3qUd3/EfWTmbxugEbR
iYqBj9duo0O71rKRZ+swrnf8ldihCDT6dSZPN3GMFimtoLVfH9k1N/fI/Cw3
Sd7TlwR4+bsvtO9m8i/PIWHn0T8i/IrSxhtxZWnFrjWgodRjPndQZSNWFuth
5H+rpYLcEkCD7bsrSU9oWyRbz3Vsb4Qgi7rELjeJE69gfMaYKXqCk147SwQk
6aGwXZeWrR6JMdUykeCqeuwfQa7NMFhr4nFhKwTKnSfszBbkUUm1gaDJpLe1
weusAhWXR7XtaNlq9pSSvXQ1XpRj5KJGJhR6eNaJSStpaaovyNTKi8SYocOb
GJIyGu8JVwuaDIpefL4t2yjmdhUQ9g5u+dz6Qvocx+tSrDd35zLh5hdfVMT9
uKzmFArF0Pstwbbh4mOC3n58snHihZ8KqePUfdlTrmhqLELSDpJy3hArKT+o
PTe+VNrWuT7LRGJu5LVefSHcj9MtXZZNFIx01eI6lfsJlLYkmsJgrhddni2n
bCow0yXUpfJCKMkKb7SDbbJd5RR6od4RNp67R+n/dD5Z7K55aQ9wfve5DiNP
2sD5iC6EXXKQXKfYleaVVAE68vETk0BoAWdzTbve80t2JvMHO5eWo6SlMkOV
jefnFvfwYRGC0TAvvWXhXYvvuew4uai2lCghugvqsYYYJQuhRBvRHxltC2rf
482EiW+GzjPfOUpx9hWzM9gXrB6RfolXgtg+Y2lXEXMTQ4u+EzrrWgERHBnJ
r3qrIJgjRMtY9BnOGH+2KYa0i8U2CgQiuNz8V98k3n36PL567BPbnrcY/snX
xOH4dQKsQACkpqzynRhK+qT9NwIA4ovrGwRvB+D+dvyqxo7O8knMZTksz+XG
6El3jUUDKVdLYN6wbeo9iw8HcElQVKbO9eCrVLggt0MmdYpwfKeRBPE1zFl+
tYahrQ9KZkJh3xK5Bgtzm/aVRUnvyokpbOfByQXgulq0gr1Gn0bHfAULm6sS
u4pJSdDJOCNTxaZ1i2Aug1RaPfxeAkETAV04Q6f9FU3VOwilU3bxXhRhsHGp
URxKDD+Ja367quk0sP7vYP5KQ0ptNOFfXNy65E2Ipb9e5OqeztpODTUDLzSG
u8V5ecjy+T8b8gUXDaumvHLNc1/wkQlmK83ZPw/7XHLPirGEP0BQGpNij4rH
Yl1BokVlMADFneRBd+BhC/F3Fsel+l+G8tImQqGDz6XwD7YAaInWybl4UoKJ
oRDhCEplK9TCvEfyLOYy6BGu1r795+27eKs9uKWCkguaDQSHJBJm6Z0FbGZ9
VEFfLfi3ckCq1fL3Nc/dCtxftdY21/JG9JbxiHbu835256cKY047UdhQHJNZ
7fMHj1n6tL7irPEt5S8K2HxDOJ92YZmeqYv4HMG+vr1Kr9/aQIbPV4aLErGb
tedACecQCHARZOoL84EugflhyZcsdn4WT8KBLQbCdEvgtYjW3E/1wq6YN9ZA
RoZFhEqFgmypr2fx3y7UYd3upU3G51dc7XpSMvUjm+vsRGC17KN53hUoJovY
spV3h+NVk248KHM2hUIEsnJouChWpY1GhMtritKp5w04REEKKVOvVwGSFxmb
ce4q8uVCLusTAPqwcnVOliF5C4ZUFMiV7D6kQXWq6w6dvo87HjQi0pJDJtNM
CldrF7erwbu/lZjUytvCtbCUWhZhw+qcIeaqDjo+lqC8rO9q4CHqj+I9cEyV
YTJ8Ni76V+8i37IDNZOtFZzgCxmNYWVMMZEDy5cjW7oRsQ0Zq+Yty6QXO0Po
a1/w1R1SUfzWmsiIr8jAkXcTHbzWzDOD7W/MorO8dn4dGtCw3292rokayoC5
PFxxoXHUTXgzcG5bx1fJJvgoVNRtbvocWnjAbvvTrHPt0P5yDHrPWLBTm4jN
12u5LHo6WZUWrTlgVYLjBCN9z3rJTlVT1kWKoKREsQpObWw5goOnr9V6oyUY
4c0dg/BUOOVwhKKOA66xbUsIrcgNh9++rMPw+aUAYxyWO2puiQsk8YUbrT+X
V5/XocEPCZ5AWIee3hyWBucgQwIL7Fh295QRLX5QI/IJFfaHPlQRMV6BMMnU
jDA3DgIoGlSOOpNbwCiWrdHBLUrcGAK5Y0CCOunw87+lINCX2S4fHH4l2wRM
PMdrt9pa9I8lcA2mD6nzXzd8qEuRRYmhOmC+nVdT2JoRfOR3x6UdAQqH4Hld
IMjHoeXMMB2J/y7U9ve8vp/VTcpE3+N/4Khk+itLF8h0cP05T8/4knn/mo/0
bbfr4PkkuGfytwnwB31cLdZsOrklztrYWS/4sbaFFSNYPD70LLop8ldRk+hP
WLorKAUmI1VN1LM9K5r0z+5clh2WIwlhkKyPklxshxQASdW5tzfhW/IQ7w2d
0mbVOJfyrS8OvkP78biSpWYQ9V2bGP9hOwFd/AGHOO1BcS/94K/+UpqffZKr
U6mtWrR8VHvp3vL//BOKiZ+aX5I50M8fzTS5rHrFWt0BRDfw+cPaD1KmJZtC
+mAocuG4E8ZdjmTx7wc/Vj3iWHaiC7l2KZy+ATuuz8eC9+/mKsXR/y055UE7
vMqAFtTn8AoXY9mEFa+La6wB3REyV/B1bVGspVcDwM4iye09o7HbH0XbJTNY
WyaVasIJBevRiyLfqdTKTrJ/VVlhFD6bQofeC4pNSXNwfgc2BFUXfe409lmg
tn2iuIrlzLtYMUfNjXDb6FtBRlckMYH5CbtQc5n7dVY69vDesvtrk+AeO0cK
GBX1Hp/SyHligX/d5I+60tXdYjZYEQC0gchBFjMJoJQmb43qmrAccLTFGYRv
eEYQY48qKU0DD39/9fux2h96k2kdN/UaQd1TtSRUiuHoJoLO7u2NLgYnW2Gr
f4OHjx9npBpoxZIUhEfgfKQE6pN1ASGSd2OKx1y6Tj3aISI+lx7HHCfIXO1W
FYZhNqAK06CxFmUPD8+4fd7NyZfde5rTol3dpb2iF78KDN9LLWZCrDGcZsqQ
l39EeFWWFExKTh6OidrrnEaruR0sEH0HnzHmlc3fnOcsfXHSDmfz3Vh7sXaO
N0fUBjCZgm0yhGCMwlyNcdfYjj63zNRY6EBjJLo3XaBV9Q3w31XmT2q4Jfz+
gmhZSNGRcb2rKxfQlK85p+ILd7o8ZjWDNpOe+M+evQ3Sn9UeMF5Rn6Df/wUO
jVtXo4HS9Ifqd/U0IXRD9UTpJfaQY50WaCpaWMaqZdtHeOxoAnlZ3QDWLFqE
OAY/mwG+LQcjA6Bh7AvKjDS3+RCDkrzRw0l7SibRxJrqqGDjEzg3lbITZVmW
j8lLPGwIsU6+t8gtUWQIoGH+30j0SlApp3D/YFaNadgjVBJkbCviACcgVdf9
/5S+1dJg2URaNl/SKWYatnmF8yhZqtvuzA+pG23nWnkxgBD7JPdufmYRXFbh
AeMC4NEnlH9Ryje2lX38veAcE4Dgw5EfT4EJ90t16pNZeJVQuNcYKFLyUuo6
H4T94iS8J/zRCBotzLxc+98x3awiL7v7yl98YABzvRZ1do+BIN9OglQgEIRy
zTvPDK4zDELEDHMiuq0/hiGl/HnZf+n4smu9gni9rfdYnIfhKOhcCOK0vKVW
2XRVDKcfgPC6pQk6DBGjLx1hmLBI9ufrOMK2JLrF+tPHQOOK+VB57oRjyao3
Y1m7DgmmEg9YADBVtO3z6tkmiMnJkBW1dIshsgfnmHzCjVs5Kf0jLbmd5lfh
p/WACASRUTAJXe+DT3P4kX/9EqQ7icjYngyMkmnMnifaxNHCOVl5iNWdAHK9
Ag/hK03vp/B9FDVLhf03zQTlz5j8E2idEyrbbEsM22zbHDZzL5ATT+rG72y1
gFfrrE3ADR1vRDXTQCNurP8/qsUSIbB08xX43j0lbN6Wk4MoV6VlzObTyfh/
zDJ5wkOth18qH6xRp39pg0ybh4Mt/gMynWbVJ0JD6LO3w0JEDnaCU8uKKnI5
TJ8KukPo6V05uhtEQK2Fg6942LDlBrbk0PJ0E3YPugiYI0XNFWbJyWQKtbgo
8zaIBDkMYayDmJENHR3S+A7kgf/hvpyl37Z3J44a5HMNTExV2/k+4ODK8p3M
njf4ZKbpyuvbXQPf0+IaA7sN5sXyCUw+S+wuRRM5qxu7nsGsaInfG6kzvQHw
OKucJpCzHcf/QDWC3BKXzuv86hrAg22JI5VKIujyQsjhAUqr4H5G+54+lE6x
kH2ylgbj9iCF0Bde0UxANuDltEzv7pfvn7RHVBKtlSPYdnB17RD18jVjBx/W
+A3/3GhRETd5tGrZmDL7HQRNvAetjMdnaIrx0OYfd9ZbC3cM7sL1g8dT9nuU
3kcrzAdnqFdx3BYqRMfyCKLXDZlMUsbFafSOqlkZhZeQYYEx8siL8gu6KcQS
ocZbGlIEV8LgrEC5IexnDREsn17iiwRnvTFnZY4FfoNb5RL8nN2KNOGs57Jm
1AAaUz+DTbI4zU3pIj+PAvgZMcmbGMwTiDSDgcn+IsU9VhzU1uFAwRMPLAXx
JecdO3/lmjvunNUrNGz3/S1P6qhhqlNgnNU//i1SXvMuuNvIcfT8VryTgZfd
EVVgZLPV+qcSwRgW5zhBxgaFRGnAvxmfBgLXKEn/EnjqExospJn9onCx8WGm
gA9XarF6RalkG2FAQpALysJhUD8vsSsiCx9R+4lKUmTzuq8aGnSdrSwkpP7r
Yrg12l4GPZazB101gRswD0MHddIU8wbRGkW7Mk5LhtYGgUwPz8xywfxeCILi
NJ3gcFwvdXDfPU5ShwYE8lc2HN3y1aXsFu40sfprpg1eJ4n61vgMVg9nJWfy
57BHXViXaEPhfEyQsEelJ+pV08OC+RPm2ZOukBb5cn/WyIZnBwa4cnQrE5/U
lD2CdGSQda+tcDRSdfS6u7iBr2+dxsS5jfGTh34YvhbW+cOxLye4yHZyk65a
zrmqMuGfryyel1hOhAE5buRnTg9bD9nknVMvDilGksgY1cXjOF5HR5NRJ7Ud
yga2t6388N4aMOsZ7b7X4qUaMyhi+a7IqFmfR+edKikS6YOSDFy05UmllJlz
dZZzBpCs0mc5LTscSV+o/YrAEKLCk/nikSv+CzLsXLYwDto7UgSc14oSsmTg
NV5OYatbBcFV+gFakb3qr3nq2F8TAudLcGXJSFHZloufjAR3D/z9dl6uq9Nf
p+YxB7KAsP8MG8qF/YQVMStx1C1JZUHAq4WtWyAPwrnwM7CvRoSE2I0awSE9
IJUQv+9awT0UvNNVRcAGK0AKLYwbAeMi1I/zJnBRIY0KQd0TuT0hl+LFWt4k
w78BbQyw5Es2j/jD3OVqPtyIZsYDqJXcDQDUfJvLbMkW8FMW/BkqDYNsvnnz
oZtPS5Mb8OibTrt8X3d1dnItpeR14Y1ElWvFNUJzKvfEUQQc+R9DE/jP1Dqk
ZVZUT6oT3x99vOcQXDgAnRfY0tq8SAe8pzqaPQKvj2DjIkW0puCqz1zL1cza
M6DlJV57H5p2Z2Ao1gFQx/Xr9yA8Y6r/euWmCksMLDrlp81n9R3mN3DIhYEC
aVnPnEeHOYz2ur/csXNgbAhH3ZPCACm0VQ3eRAbhrPj9XwWj7/tk5X3FQ0l7
RTMqZxiFD4exNQb9C8IcJM1H7RTN8xeOSJP+4eODM+nLj1OohSZq1qJsinP0
qK//FKpJDuf353p6q4OtuaXoTXrQnyZwQxMvATIeL6dOI8XMhkZZMDTUV+2I
Zq/eWjbRtjDVMbVIeVYPeHjJaoMFhLE3D3jt0C7XtqacM4xrOv00Ftd0l3GS
AEv1jTNlWQoB0IdRZDy4zW+ueFXmdxklN2/PxNyEQyFkSNOOrfC85TuoEaM7
2De9sTdkf8Hn+jeXKkvr5Xm7LdYqiJwGyivSjEngw1R3edGKNwOb1+L8IUMt
JzeHxnRMKYjGHAeyS12lDJOV/qCAvTKynfmxXEhBOW8+i5iHfFVlMvxVOmsY
rINfay6hj8oZ0PwmUITAiF7ZcYRQWDaF25wfiSRka0sEIBk5Vi+CNzfQ0hF8
4BNjG6rT9s/UV72MboNsQGI/DLIyZ55hVx4Qj9tuT9h9wuEOaMPLZDOt4/cw
u6mRyz8VfVa0cwSAKtVxQVu3aYgiylj5bLavN4u2yP1UGom7BUebazwDFyIc
XbCZm3MKZXtP+rwaCxgAnK/0gcLBvJ9Fzote5DDc/wviQA7S5bnGSLZrz/Mw
+ESr4uyPy9mOjDm1NMzb7ZUiVYYjZDbraMydG9PREfEtSg36iiiM/dS+qNVR
3ScjLffJrI+VDVQ1HNUJ04epbpvMmqvwSYOvz3Y+F0mpzP5eQd31+wKrHtbv
ciMiYtRF7guHXe0vShWQMGub3trYkO3w0q8unrqJqc+x/2CFzbPXVxU1vrwL
QwOGdQCzBxe/4gs46xciib9rm4KbU478CSouKYXqoR59rmWVsnuFQUg43UVj
aRDa1Y6amzc52kA1u6hlSpHR9f0wwpgYlq32uzJIUun/+MXMj3R6El1GS0qJ
h69aKF5zTNlZbcD2SrKyWMCtKvKYyfoRKk/T3cuY9bjGtBV0pcX9NJjGdIVF
7fCKkcCOc8S/yE77OjbppJ834ozMZSH7qtsTvTgtKqmmbJdpA7jDpPRVOlcr
0jwOIOj0tLmeBg9Y5RT/DfXxdkRqBJEo+GGXkdrzBXzMVnqitEnBUqAxRX0g
2qnTXgnQv1tmKo4RV2WER+91kW31d74mVOMq0DyNXP9hdvq/sHvx6TDR4Xy3
kpG6UYf7aXsot81TSLisgSOXpDpfo0+xvy4Mhxv98wfjwhh1MwgUzkmoe2CG
yMaCDOyfv61sh8pYmUe8bvKgG/6r4VVDDnBiSJY98qbeNSUCEZCHC76ShY8Z
awdVyoXQx29E1j3B2HxQB5jYEDO3V2EP3TOcMTFQf9gQSJYDBkZ9Kl+GQ2Mu
rbJWcEFOkbcTCo+UvIMZyMtGk9Z8gA/fJ0X7UUN2nLrkbCH7iTgijV8l91Ih
fY4o6aT4uLArtosicqZxUEZfjlWL0eHIesdh5uO6YZUS830O8dzB8ZFOvsEc
k0IEyefauHO6Zn4Hk1vporP81tQk5Wu6ulFIvAyVm5SFY/AAYJjho1EsAbl1
T95jUrXoszbEkRym6n9Qjyac5nirc+1klhSy2H2PZErmEwitt+PKTCCgOjI2
i4MFU2WbPgmlDoB8rvG2djEWtmMYsDytP8ZP6UO8wqvaTz0ItDLdBoHgzi1t
ObGwlK0mWEQrWw3Tg4qhBniEdaIQ5xJr9HLN6/pjUSf0yjtd1cLQ/IsWLzD0
JRmV5TvhIoVspKA7LZm+No6+yPcKwYCB44xLIazKWZSWKs/AHgodZgkHGad5
TQr3bOk8+ZEq8n+EeHZIGkdOhXiPip1pogoVSJBSnJ501Jbpi3e3UQKpzlnu
eFmet3+tBKlkhlznMkQ05Y4Efaqm68VdMXQxfUZ8RMtJsNgQy8LWP9Frjy77
cT0jzyQ2GE0oRYDhEpopHePb91PtXaaoVua+fuOo4mOBmPotj+uTvEvCVmbH
ymaaz7DEfvt2i3USeaPgePEXdm0FlIssSbaZD4lXepfujxcFDqqUNrrpcoE7
hvsIhRzts3o7mNivinpbaauV8WJX3X47KxQyTgcy3IS8/ScxFChI0SplcVb+
3YmIZWGKuz5plQL/lfGiszsIrNd2c813R39TH7WFybDkByi7SsoF+rzuudft
y+f2rEeLA+xwPkysdl0zsFhMmDOf8hCmCSlGXnNnvp8OLQP4rqYlkfiyQIB0
Q8kwi/1M4kHwObUaySAmHPMGfva3yYMFG7uZOnn7rFujXeCm4UUVvrjfUk4V
Lv7jUUG9uuXMl87gH70N0avUDV1zmG6ceO+OmtHexRIQBmPyywBss+UIcPti
mREEznpPr/PeKarw1MbHffocGp7Mlw+CSjIdALIpfsv6rZD1mkqCnnPkJqzy
j/B88lG/5XRlOccpH0sruyGtdhTk5sOA11JTW6wmjUiiyqGxrDlF67X1y8qS
JENZaFZIuRD7weSzoxOTKCDXWhA0/fkSCOKw76BBU24CjOS47qQtaULXVpFk
VpUkk10/pAHDdnmR/KMRVPIpATC0mby2tbUCToRRwXtN+dReCU5SCvpTvSug
dR2OEYMfbWNIi9w0zWgQVUl9l65p48RBrkF9p14v0p+rNVVxsrxlWPIJNbiH
4VVGzD9pOJuvjzp6idMqMyvcqWk3DrFXZ+/+MySoekFm9ZljBQpGcresmEgy
wajofdoKyHcmthrAx0nL66tAzqGx+/qFHr3xhNL0RyvR9Yx2HcYvWNB3i/9/
hl0T3WPd7EtV9d6iJlmGfLopvHRvZiZrcotyVNLvV+XEPh4yUI/yNpyf7Krk
pmcBdOeEuc6eeNDtDS+un8+2uA/DRXLDcFLzHVZ4JIVfCzzdvNyxh6ktrX0l
istzl1xswc3x5jn1U0CpApwoEHDrteIehZAx1BU4+0OaNZ9IcMmynaW8n5zS
FcHK3he0MgtuPAFzoCuzkvDIc+m6p4UTOosN9K3O8FtQjUkUM49o2RL52A62
9QRU3cj6qsJMnhynJ3nmi+mluXbuFZjpC+Mc84jFdHfnENch69w3UwL66C3p
684jXKXJUAuHN6+9BgYv5VOnl3cSaQtiRv0PICRCYretjSrDQNqJnEMuhQar
DoDMZzUDa3zZ29XA99Gu86xDtQME8KSgzW2FTJmp8mmfFXSspUjPYXL5gfrc
jslKGJ+bVpgmJz/nFkfxFpJHPM/4WDYpCwkR8LCBx0roCk2z/fRwdsjWZEsR
JPav6XhRhKo3cy/4r8me3DuiEBs8MJqzh1BxLss1Y3t+iR14tlLMRBtiOEi0
zGLxfA37FkFbhO53+WJpBKiNSy1W55OuLiaL3dkmYSZCjH5pxKUMFIT+kd0c
oioTOsPxU1kB5v1i8pMAk6XPWKBPTJdRwGRgZCuCPFzSjhkRuunoRbns368s
pTRC+Nt/QvE398lt9Ll3rkv14+uEcsYufXpQ6fX1GScy07HfXK0jUEcZsvkF
iy9nTEJsgiJ0Oe82XTDxwXvms4kZeRa8dOYh4IRi7ci0GK+NF3H9/m3aw8PG
xhjSUPTqXsT3FAqpcorZStT4smymNsHWqbvufOlVp2pkK8Fp+n6SQfSsBIlg
wEnrqGRVAZaQo3Es6JeRDLOe4A+bXIhDxPjU4l2bkVabeHh98UNmq8q9pq36
msOAfHLN1r6Oy540NDkN01VC5UFVTkVQ/OWyX7SLgT9o1YY17T8078fqC12B
B0L8t1OAG049KqghQT6RHqw/I+7pASIq2lCA0TPPrZozpoPGCEVsBDy+5Vp5
ql+8agG7Wrn7FpIp3uHx4+sSD3RfNtsHRJ//uKReLUv5tQyvWA3MDJjQRic1
6GxvEth5MNUjmGCi8SfhpqO1I2mY5BPuB8eXn46WhtYDB7ZZz6UwmlViWFOx
a9uTjoEc4xbuzqjefz48CpB4MYpX7kpZS3+bPujzbn4AwTl+boPInTpxd9qT
2WccRcsU+9UdeuO2pPexo8bAKW+obkTwtHyF+6Kd4aGb4sdTkwCk7SoxcSpF
9Xm6Chj5fBqzAcrLtHpnRfKH2H2p1sqlL3OQrI5DsSZZUnkk264YYyyVlSRZ
3wKfpQzSUW0Jt1m9XeNK17dNwZiwy/ojWKjcL8fUcmX+szeoqk+KUjhzX9ON
6BEziVjdckAWAX4iBkN1tqvzuUb2oCaivuu2zyY/PiLDrj1yc3io+tnuVyFN
FcSEJNqj1M6qBHQCDtFLpsYSzgIs3QNQKgq2nUw1aBcWqS4/LftHFLGkAZTO
6d/Mj3fDa8Vkul2q+Ar6UHV6jJPA74MkLAeY8krS2hr8B4bZzs0ymE9yv3S6
/rE7PUVLTMeRv4QGfB3TW21JIVSFVL+ayNNdPyYsriXjRoB/nut16gREiybp
tnVugwvHLqVCA4Ko2v1NZFE9dGFBTYQ3Ys5GBdmB85m5cfts/03DBe6NAg4x
UnR63y4hszdVAwfMaJ5n2xXBzB5BcNUadhcvF9hNTUJk5izDz3RPIwu/l6cF
HSmavFIOlNBCnUbVKUy2LHawxL8EbnkVZIWwjBCZ2jjB+0lWf1UnVDHa5SSz
aFB+D2b6/B6bDEZF8SpQl47Gw+7BpVxT8mx3BEIiu2LSVsSsbNDjbEmBEfT8
C4hbILvDTowtz9so2hS44Jb1hh1Z0Ujssz7aetVkPVCxLRQQ+5wyhXKT7AeU
/irgNFt6r/hP9wFmOVUvIdEdKt24/GV4THlhDHs8aYEsEoZY3X41duCxY+cq
+aniuR3M2ItL2mWPuk+ydicmzBSYiOp4c0sYHI9mFD45/Lxu2ZyhVd2+Iqxq
Pz1GBHei+qJZLhrLvP+hVUEL7mg43EiY063cS8QufHXiRhz/lvtSJI60dPI0
acjna/WFIhcvVHyuCCekodEbOuhDsoa4NCi62imeXKByIjeM3RdyDXcAGZ5x
+llspwYCYf7srp1c1t0AQAr9+hBHJ2h6SSXFZyy0Xnc4/45b0pbCV5ckHGjp
wD1jTe2udyW1GGd+nduELmvtVEmmb43ml4WHGWl1I5ZGqQg8jUWmkRwPCHVe
p6PDfy5x25b/al80v+qf8cQ5XVImW6QVZdPsx7aQq/Fk4N0DPtqebPCBhKMc
HqZIYhfwrP5zlYQFAeqAZ6F97ZpSmT7/fXZDsXuq+V8+aEbNR64c6JuZDSFI
SaYAx/AAhxpOacOrwq7UWmw024oBFi7G5zebXv27WXYlslMWTZSIEkejz31+
nM2MlHJ6j62UFaaEYF2uzS4b6vOUQFKC4GhtHxcvij797hcJCiNK9VXMo8pb
dSxPSrG6gRc89fv3wJT0HloT3M4C652tAkLJtFQDBCuYu/nTlYcF91/1QvQu
tTm9fuPg4FeqCDZTifztfeKIdKXtRzz4aqTf+aqPnruprmtdoceSEqbEML4i
3Hm0dz/sc5Zaf1AkRMtiHH4BeYoW9KRLiyOdf9AUsoZISAJ9X+42Z/+94Eu7
ZGqpjhR4xUYIqWE6YmSdJqMJfckIh/FQ5nowMmHIL08irGGiaJdjglqC8RqY
lz7lhDZeez66liSefdVZgs0j6cqpMpLezp/c+1X8ymKIf+qDx6xIdkNNm8OR
xSJcVX40xaMOJQrnL1475U8TNne0ViRX5HS1vnSTJmmztCin+Mr0TdB8cwyE
K/lNf8L1CWy5gFeJVeV6biuKbGl6GTU5C59Aoy0eSRQypc73vd1qIZoc392H
yVaOOB1QlEAtx6ACMh7HNX4Y4+/IIpuzhXa5wup2D9DMnlKeRBndscWvDcNc
+xpD2bkAwA0lwJJxMstH0TWLB6nRxRKbhD3i1s7+aHzLfSbnIY3E29LvF9c8
T1Ii6NxrdJkNILlHTw55c9nDlDX4qxX6DltOAAsA8xnrBRvq4rCdaIFvHlpG
Na5t8a8Gm8Nn3PorvUMQ4n8Hj4lsai+Gczjwd/hMAEBOg+EECiT33T6SwSkS
BRn0/tIMXv3e3mCAG7sRgBnPuatgSeJ3mS9cqwfrPCzf5OgdX43ZFsRtGqXe
DFn1iH45qYEWvLe77F87ogyKwY+0+4XGWK+GcTjoPz9lZFXSMBqEe0iH07XS
Jup5QbvgADz8gGce8yjikzOEcVluRLRc8wVHHZqwLMwBlR0sW9wOW6gp4Tak
35QStGu04cUuRmnRlxcRDAgkHlc+Ecg/hUJ1vA42URtdOkZtzcHJkPU9D7Di
cVRtsViRJ1G+jMpRa8TRBJmwpA5dkanDAjRvUPjQ9zIXW3AVOKn/QeN0gnIj
BfNxnOWe6DgH7Tf6FXo47aKkZM0BYyvM45xb+/LK4k/aOQPwXHfzdhYW86of
H631WQEYXsNZr0Cqg2Ti+b1i5Wpz3y+oRH3+fBc3i8CfI9HxCe2fI/M3bDqB
Pkd0Rq+nEcu26VdkDShIHlprtFH9A9aJIcbpKEddo0ykK7ANAwzvh65dGdJi
iigeS/zDSaelqm7wQj/iQVyceZDUFzQ2GvlK6taglXqhfZNdzgweh0qSeoWu
TDq/aJq3nyRoAj6A0AB8bBbz/OSsGdRFPLfaokoFChK5CYuxzY92uRZ+zvla
hzkWBejxvfjyvJpEm7xTZ42Phhl117Fs7gHpJLKWVOMz9ao3w/uX3BpNRomh
ofyQfsHVo8TCmKL0Np7+UV1XuEdRj3IurSE/BTGLep6M97bCypbWLDzrlkjJ
2oKGw606oNnAnFx+G/b8R8k8km1hyTDS18RADsJHhntlPGJqhBEW/P+0aJA3
WjjqMF1wIkY1l8jkAhSR4yqEzBjCMRwYNFdRsvKrJ8f0HyGncwSzBklFB829
cHWsr2+CkkQ/4k46pCnFFXzBPC1g9wl8bg58I9TFzxxHh2Wp1DMazaRlGvBb
BDxQ2omu3xPMRJYVcNhuKmWE/xoul8bUYk+NZ/waFDlSH2DcHltkoyN+2Ulp
BurgE+QreADuAJE/kaZ/2js7MC4nmn7A2+TdyHIUAQYuOn9qu4d5rIUHEZFG
JtCaj8pBtouQAqRPXYOwYybe0jmZSDD2mQO7zEWHVAoJZtvCVHDZFQdYV+P4
sh4uPcwLB1eNhCpJUUoNPrqvA+jXXV/6Lgr7RsoJ1sHo+SZ1hp5NlkwzOMWD
rcpRM78drNWrLiwPmKxMlF2ANdrGwRsQlTtBCkfFwmDL7VIFHnlLKRlziICQ
PsEwLhuxgh7MYaGL+Q1a6YAzzjCLMliBxq95JPIMCfskFahNPtJLHbC5MAdM
53pE/A/IxqZVrDREHMtND9f8NTG5iNTJ8/i7nqyUHNs0rjLFkYTzOwpnh9JZ
4QvOX2HGzzDNubGeuar+mCObLF2R5zNNsRbCQQ6yirqID2Jpzj51uJw9u9nr
4ajp6uRgJYrOgNviTCn2ltJlEGBGiphotyUpe9JUtL0SNGoBCSufsWn/TBw+
Czp7aeWhFeI0xq/uDRZTzFW2d3OMCBgzVvMAoOMOW9tCitIveYsYx45CkI6H
31zcfhA7gg3U8sYg6HbDE/4XU8wcdYlc9+R3eDsoHt7I42qqyNxXA/N0X2Ga
SPv4wz74LWIObMeAyupnboMfmV7AzU8D4XGtaGA8clrK15CMbESoGB5BqYd0
z/EV8zovPOw/flEjAlfzu+UNc4jIifO4A8FVw4E919q6K6VJ6sf5RoeDz6e+
L8NUkAAxGgRGy4joyqB23iwTph9BIkn8uyU2jJl1NRuOG6dyFKoROizh90aX
CPczJrEh0Irk0O7EnzyElSDofIdMY6OCJvIN3cI4GQ8A29WUQ9WAqP+IgbQ4
E5kAakXOEPhLrJfxGjkfTgYxfRbhodXcHn+aUUF0FLEffOHNnNL9oSgtQYQP
nzbYRK4dUjSRv+pKE9sC/kfxQt9dWBeHyj/pL3szk4N2fg8Z4A+1UGjoZcVV
zSwEep2rwCnzIHbmxHeTTtiUjLufcertl44sLvx6rrWpZR1LeZLCTM0TYf9J
KkJCXey+/eAMJieP1yf4650aST2AIs+RlC/4JYyXcSO7qpO0woRh7SbjRX0j
elTCTtI/+rFwZw89wCgcvAFpkUwCRhbIjPHDzlxGb74gnZxr8oKItSFXmFVr
sBL4uI0XhJwJn/dPDmY8lPmdJ256zKX+03yqounYwNdwVdj/CfJG6SasjZ1/
mfsZTtoh++mWxOGxpmVUjOAQ/lUTFDZD+OIBI7LSFCCnRVpuUeiiAhsPFR2B
jIY3RtT6nJcYL4hOIH1PEj9n/vlNHUvsivTKCEBKMMyI5VkIrAUJFd7xllcV
5jZez673RHyQu79nlsZVTTZc9E1nls78W9VsbSdIRx3Kw3sh7J3xGlIwfH2M
FSo29XeNLVTzQGxXxjYYdWMZcvMLhn+KyHO3WgKuZZ6ip5XCCHrSdJHS03Fi
4NPId9V/Oj1mJo83HgTd47z9lwGXYaE7nSUbiMtbMHY6Oz7WMsqJmPeu4HOb
GeXA5Ar+Z7aWjuYb28xyctTz42ppuSAYPBdC1eVn738CF8COYE/UM2vpQ1a4
bYC2d5uaUjIdqV8bDEMkYWMcqn6BX0tcheFIN/vU6n/QMCRGD1axZCwk5fZw
c44Xp20dyV4bv54HCvc46ZiLOdmecaV4XjupTUz3U4XG0w8OoJCeGn3rh+qO
eOWda8pOzLkbecAiRYpZv1Q1lBNYeRN61IFrmkz1vKVOnkyCU+2Or7CbcxRp
A+1eOpQvjQahNnoZ+DSSeVJpKXoG67ZbLLPjpkS4d7w+ssQ/IvSREJfRNo1P
oC37ZRf1W0Skk7N6GnEsj8VMdxuxR3CwnmZe9eY3prZrsXjT5j7m1P/dGcvU
VLPgz4OKVA9msUym2JxMXIJwAp6zkVCeISoCNElZn5qBcWJ7hroD1XfUbG4W
QF841KHr443vfMsFoDBWv7WShCeP/CTGtoZsUzpHPVPrRYBDp6z+TfQW/X8a
Sl/Dp5Cj9wzF+0eVYyIdSsvol/jjh+NtAAPLvnaqO5WQ8UzXMfNj4HNPC4v8
U0OoPOCon1IF5ycRw8EvoFXpV8CeUmD+90iEhvmsW0NL1j/48zFzEDY8Aj1/
hgYWvcrUrUGi1VqKzJx6f44WUExOzTDYZqu3/bP91ARSpUYKvhcJZu7tWEhy
ZgFA7nrKfiGsysbn0wSP9+99qfRIhTHWJgU0WnSr+hH7QL9RIRM6OmVm9atk
BsKFk5F5ArPLQQTH922YxCoEiCUpr50Fj5fahGU7yn7xmcA3Np8Nt+Ae95EB
a7B1+h/opt2s4Wy/tgjffY+6TngDAM8FmXRBN+4kPHYSecTapoAPRHgJN2bS
WuvSTXrB7PCulkWgIvWax7MhTRQtzPahQHo5kyYFPbpngDgFpkKC7uHO4awX
oj6t9oORffSl3kYkPFkUhsAGPIAer0dt/489E6qrztInOC3GlFeGN6dDF2al
hE2wejom5toG4Xl2un9j2MLm6S+hiqoqBPvxier+YItmC/l9FoUDUvYsAEdf
UDZ43fe2q+mDkwLUd8d5QG62TVq/vcYlR/lvHekPClExJ5ea7FIB6NBF0bNG
aRUFLpTpJhQhz8g0OChT+vcfP5x2nVNk/RBr/g9mg4zo4T8G0fG1rdMKsW+J
S6SCUCIr4XU47KfHOVrilP1/jg/ggx1FJQp8CDuf6FjJJdwacXJ/jnegfnKC
U6kDKOu2nlOb+YYdTK+sntnUmiuMEWmfLWIMFdVOvddB3vNrV+J4+GhnK5F4
/PtY2KRxAJbYmsXLA7D7lxkwrt65eEstyBrEPCY1EDH9AVFG2qhDTuLiFE7U
2V4WmYgZeKps7spJf60V+WiZacJlcIK2o6ppdVPmHkxjJ3bCpFjko+3rojSM
+PdkiUxzoykKm+Q/xdpch7BWt8e8UvbdPIOyqaCwSZpNB49HOIH4ZWSDMonw
xR+kFPX0TqL4nek+vrwVBwWn3ORisWIFVCuGk+CZpB6fXrzZ92cjljbsp0QP
H/HZMydg3EeYelTAwwC0ePL0gVOPezTIy3MzWwLU+1kw0NBYKLvdYAhIIqhT
h95nB0Gf0cbegzO1RJF22k42Ue/SbrJ1rt/1kHeTxhPD66fnNfEKh1kFaapz
As/4pNnVSeAjQecUkhjPoNd7Up7iTJ8Zk5Pbto47UYhYlRucygQcSkck5JJn
1YLzaNhKq6ql21b6JEkHkwn4r+ByBcJuwXeTednxcUD5oGfb6sg/CMGwIZIS
GElruVmKQbMIUs+atyhFd6QrOK/3otWLR259EvS0snhSdloCvTyilOGIQk4A
YUr/EdVKXrLhIOCf+rgB2t96H0+kp4q97C+Z/p3cJHppCXM2FgQKVogh1PuK
Td5YjsTfeArj3RVUBqQ+0NWA5D3vvzmur8ousZvGRtuyyLhr8V/F2q/+GVw3
o/Gf2D2fM2Q2aDMKUtblRmmWmmypSo1LXE7Pj3I5ZufSLuibmfPhNZmS98Up
mf38eF/iFkUHe/PdgnWbtFVU5PM9up/AKVyxCyAxzzTWJfASIHNc4GFXeaxU
2IZnwTCPn3IuZPj4J24N5+sZpj9eF/+Jlpued4OgJSPi/704714h0oNEN8qS
Tjm6kjYhuiUtb5Vc6ewEU8PZtiEaLBcmyMRm1dipK3qwpdjUHBrI0VoPTcxl
ESaQB0aNait+/RdAUf0jfvwRQ8DvP91toQ1k0LDQ2tFR8dpvEHiNUYyHH65u
OX/zKVsnJ2zWuQjFh1Q9ymUHCQcA2HuMuKRIWSu8TqNt5ol7qh6Et+nR+6kM
RzA5FjXhPXY7R6imiYKSj6Q4l0lhgRG8QQ1XKU0Fd3MRrzovlmE+KuiTGlRo
KqVM06iGE2IJnAqpEK8KOIAyJgQTMs+iWWF0dzUb5P9FhZIqMJXNZ8N/aiVk
vNHqgrvnCmy/xiPlMZW5grwU8ky96YK9SciW2tLgjIaOAtkKaQnQodrjlyef
7tp1kJL/QS/AUBNsgFpJqvQ9d9eEciRVFbQ+d8RJmPtyQYsRxGPk2ffOysXJ
8AEIpVNgx5rx4W9GqjH15O0qgukaMv/HZvhyp+AiOOAHSjnVOWHGeeF48uh3
vKB/Kpv+QZeHoX2jai4QMIoOhHmw5Pm/r5NAeHx8DWGD1FUYa+MbjQSFbM8S
alRcpCciwSErOSx0cchsFtmBvSxfAhi5oRfAXM3HzicRS6pJ1HWmlqlkooIJ
e8GBrv2+eJ60XDZ2A5lmb3VTOQZkUXNFW7yRpymIYekUVsY9kk8+eGx5NCQW
U1DkCbHQUOv2PTDVa+ZKJXO9SMxWgxvf1CDPO1/GDzFLAEw+RGcDo+MLrZ/n
pIko1tLCMx/u30G9kM2DtcYzcpvmaJjZcdY6Z0rkBEIYrZr6oRKxKYQsDvl/
U4zWsQ0NNjSN/sv1DSaNIpTHOitRfiPjKx34hrmNctxbWSNmWzYgJMHACOw/
k79/SGgAm9pK/+7BRDj8tkk99kPTjS2J9flSjcpDPIEm9vtUQrevBYrKRiW1
5e626qJULR58qvo52FwdVsYYCWq3JGoI0Yls3ockF2muOwLsF3rW6k7hAJ8F
fHAxA5x/dNns0oed19POO79ISYZHjmFoOcJgKzODlcsJ4W0sgPOwuXPdjtYx
N79DZ0CFRmtir2Dv/fQvFhUqdHZ9vD91iWsw4AfJX+KRUVdoXLgKhOCv0Ron
8qib4rBAC6Q0zmZtUjm4XYhv8sepmlSu1WYCubexm+ElTtp5Wx6Vl52Pwbbr
Hs21/iN/zJQmgWwNCUK7guKVoKJrgSv0rkcT9uRgh/YDI5Qp4VDKsS/DU1Aj
V95ELgOkJa40FL9cwBE1f5qxgi8NJSMLImv4crJ4pq9qCJo4Wf8j5ElqALsV
76k9kHaNW8vL8E4BWoqtOvUxEOGU64NT38OPvy4H3CqP88z63DKqydbzsdrt
0OFDWnKKOPFV0dXNuE8al6TPaNJhKOLF1aT6nfs6upTjtaPxUhz09oawqj4F
2WieutUIxBbGBWVKRMo29YY0EHptjOgWYrEFsbEm5WywGL9tcZATuU8tJCLe
zmTt+EIlQFqq+RDf6tKM7CfHBwU43Wxp2bBnuWSczwAk3Yjc7cpDMynDf33l
LBNZwtKVy9HAIrGszaRTeO399d7NZCHtzfQJ1eFx/iN9+cJw9eVEkNQBZ+rD
kf5DjG58dtrXus9XS3Yn/ukw8Gi0ZDwZ5pE2rDjmEciN03Qul1jkwh8dcFxf
kIRC34m8hne63NadJvJja+SX7Z8nzTMSlfIwgxhiSnifAIn/KA0E+1lhCqJg
+RkfpNrkulbzY0LY5kEFRgA/jmzpHcU8rbTFWEVLoc1Zifu/uaDkpuDMV0ok
pmJifsTu2SsZbfq1kkx+hjBlUwVNO5BEDoq3WFtGfGTIzMZHLh7BePnkXveo
bBmV9XTcOcwUkN1rfkttm+8Ih1tYPBKQD0FTeApfNx+ZZqQTznXLfw4JlSM1
nbOguDOtfoqCwKSiyeN6/XJXnNdn8VT+vWSII9AptKkIRf8Hqr66pfhvnQ+b
mBzo+wW2oE7jkMmJHY8pKfHmPp8YVV/o2cltGHp/CdT6ZUhN2iJSCTg/O/dk
oBhnZItYp/QVy2nQD8oLkF6AIjROMniny/uZ1yc+7H/mJoKHujEUNoSqrzwp
0OEi/rR+uwUz7OQ0c4lYkpGTO8Jb2IIEMtUzARTfUkxZUrp3waw7tATfwr8b
kljeEewNE3hisAGIziaeQAxoNtvg83Oj1zGPOA/48hygjMtbYe6xhL+gCPWX
6WUa5/sYE/3MSWD+PPfFtWT+924FTFqt8csqSw3nWmnUkSPrULNgRuQTFW20
iBrfw+ir6Xx+FCj+hITZO8PYwf4gmwDbYUysIKv03Pw5seccyxdxjMrejp3V
EmER0omb7tdCrzewh5WAlhKxeZjUu3X7k+vXI580eOomtZGWdUaf9W4amRni
yaNfad1SUCwV+mGDAjYq+DfTvIRYcMA7TK37JMh/qmkUL72jXjtc2Ck4VHfy
4kX+lECE5Z9fHN7X+Zjujn2FTLlFQuRelKjU3NlNe9SEdIGOW8Y3QRQwRtmt
22UvzDmWBIaiB50QKODEGZ+2LUOZve5ktworMxv6BCInwjCON7fG/Sh3j3lv
3U7YTbFbvftdd4u/mC24ipTVjfpUIP4Y4ZkUBHbbocbmpvkqwhiFamxDlLAR
ysCkqlYfIkcK2D50bD0igmajpcSfvSlc1BgXDY0iaGsfMfQp214NPfwFveWb
rfeX416Z2616uL7ZUQnVXh7kMC60vrfK7g+pp1yDBT2vaXGvfOmLNordXl8e
Zn0y4bN4jseawi0P7BcR56fwCpM6/ZFdY/E9WmCh5rOidflRs8JXCqpYkNLX
WX2O/gdR/C5Vp09tAWhZdci03Xxo7bAK5wfxh1ygeGELzqvQ1txI718mKotq
MOGB9PCaWbBIpkl2KzD5fze44nWXV+SCH0a5NJ22A2XknHLX6Tgu3tRqgaP7
LbIoMlLEXRolvqGZkxjyhD16gVT7ZR5zUQwBKXTEBgfAxYp38yFb2cRfsyKN
UkZWZQyP/30zw4yF9YV2VMHlZiMsIaMoRDeK/w+aizB/lGkeC1dksvgWVa5z
wgRTQgNSYrwmGo5WYI2nDPWiZANeluE8FYweqrA/ADrZ9tNNtLz0V1q0E6D4
0MnV4JLLzqXA3Y39fdg+x1LnZ1keGWCjKPdGipquubdOroaqulyURCS3haQ4
4m0N8shk0Dej0/E8UdS47SgQhngDINGxOj93FnAbRm2+SrSt+sLXUcqhaxrh
/wRj7V7ZQRDHTZ9QN4narMUCa7v1Ng7HNNRFcpGq6Vk+xqesFet7LJto3dR2
RsvNhzoic0cJiA5Qa/9dX+o1sBItWRN55e9EcxPrD9s5axjeweMdBswdhfI7
Z7Jc+TD18gBnLVPtZSnJyQO5zA6n7ULB4N7dVNKx295hULgwpwIrGzX17Oh7
wEmyZU2o3oLQroh72QMlGFdS5L/mXZefspbGl6VQy3NWV3vfBRibzDJTkkdw
ETEsKOx2Nrnx6wOtoAoAxfosUiCgkdrbMDyAaUozj81zfUqEevTFVpNEork4
bDBtr5IlQXUG/sfNS7J6OjDAa8eV4fkB0c32T807GriuP5FF0P4d8l38BSK6
G7vlAEKp/VYRSeALBiT7ZX5yD8tGate3Exc9aeYdQoU6lrkWVGOrTRnosiQ8
NvqLbeXVX3rRMXVYfFwJgzrvkz8/SLT2073VMKVre4CdVp4DGl8kUCn7wnjj
XLQHh2pZwl/9C4bF99GMv69CA+ntGkaVL2ZX5GlkSbqkCm+k59rLTdTAZ3Ld
PXKKnCiZvmB2h8OuGJYMIUbwc/iBNrI9pzNL1pbF/zKe+HHCPQqxtFz5OHfG
Onm8TFF9xwTW8xM7trU3pDg0VyTrMoYC2e3oCyJTat6rvv71LlEEzVZzsd23
k9ligcXsMxIPcD9De1ixDLlGt07pkoNYTQi0VC7iSrM3y6akWGJfIbZIxJbQ
l/zDymzXTSLfHOoZI9Bx3mH92oizq5xvPww5IEqCnFv4mXaPVi1LmkXKSOF/
yXSmETvKzaTgFCtB4on+r0GN0swGRvno/SMf23XkUBHuJTK+LjwR8ibsHDuJ
M6+9yr2T5Gnj1lHFeWyuSjnZU1FhHZfJS4+RO9t793g3N4JICvSnsXOcCSAP
beJR0AaVCGH3ZHQLq/o5rkBVV7bsEDwId0Lb+F5uqfYB9q7oJ6Je0fcFqlZx
Gx73HNhJW+3tAjvM5UlBxmmpdkVVB1BeTHK710u0fURr5TKqCnrrLdGQKsSr
Q3gBv5QeJkaKZMiPGmTChJWrYdc1GnAXu4OYTUkKITbu1mHD6cea6XveP8CU
/1b+6j4qtWfnVPLPqGqWQ7s/IWpVBWElJF1sP6cUPlVOuiqxAEldoX5xH/jW
Ej3nxhZ6x29mC19L8WwDRlFiSNS14AhoIpjU0kKxJ5KVFbmJptuDkykytUds
X5Ec+y9NRoC3cNocCAQ1r6Fsxm4taQoc/+x4NzHobx9++4wRb6slG7WMdkNi
tbzejStDwxiGogaUcW1EYeRNXIRy+cZVHYirtDVPB+8FQONqPtkJuC9hNQ4Z
Jydif1Z1vGPiHVybHyZMdmxUz9dyPWj/4F3NsrUqq5eD84jLsDASe28o8ezY
y36Dw5bpapSQrciBJsys54G85r8vcDdI30XmKpMRK4h/poLqOAq13LXku9tQ
4D3LRjFKhU+mlg1OpjC4kFbCeIXcYquZlaieO097QAuqu+knijVDFmWCCM5f
wLzXBNV3a+dMYISqQ3HyDNwpoqTjzmKwR2GpF3za7n+/tU/nalbAQuzwSd3h
D5RVC//sHF5ftRuTii1yzj0g5STQ8pmNoUtGsYmAIa+igCr1iUgXrfba+HAY
nlpT5xqgd9KiNg8RBFVXhU6uzRqOViSFolFe8aRJCEQg4gNCDIZ2rt6m7MTm
mIhXyrU2r0CaHg2gTUh6F1FDDC8ZOy/ZojEPur4AGSTjL9Y3/Jjlc69SfaAH
8fWi0SjFe8hD7gcubkWskZIYNg3DEtBmXmoBLW71dlPR5X5b0VMabPBAWndF
NuS2FJOx4t32jk7lJ5JoLVsh+Ud9kksf2GWgrfxtGQqWg/nS4Wn4547q6l4e
xzjuYSuDE8pFC4icKYLNsD79XgCq3TADZs36z9v3z9wJkUnHQ+mGB/BfWheu
xhwMULOXBmSTwhhVUv10l/VsckQj7jzXKzJ7D3b6frqpM1fLOR2mrYYde9N0
lmBd53vtZm1hQ5rbOgilJq1lJbhSlRbn8J5h+mYBF5B1U0MmdG4+xa72VKVl
QBF41lot7xgiPW8xRe0E2d8r3IEoYOoI874laIvA5qA10VeOh+Cflnvq+by4
VZilcqsYGVpIgVRh30vUbVnuMRrDa4odyZ+uSTlJ0gLnw2QIYjYoo2qD6im3
7bGLQNkSNpYnn7s8EOH7s1DW0G+GqnaGdV57DOhtVbUwZOwBhhO/4D0RI1+i
jEDM9ssmP7OOF4cqsmHheg6gExPch8SxGxarcDZGOqPwJlXz65jGuhz0pTsO
IfvR6gtI1GKBVK+9q3pJFHt4XZY3CKDbiyCo5ZxYwEupY9JKCULKv1x31gzK
LNe5ie8KvIxMSLPY1WGgP8V3GS8s2WTNxj+p9SOEuTZsOWjVXfd1GzRUyoD1
DrGwICMe7CCQ6VJ4vVbsaqqgEWifdMPFYJPLiKAKbQFmgzyKNOKDxD+jMCqc
D+AvoNPCTF5DNY71R+k/SpgOt3/Ru7YdRzRQUuSwHHfR3++Yw/mp4oVXGc2+
lmlOZNs8DXQfRI4elojaGnp5eOWdJtPbGk4EM86ofH4AkW7/O17vSFsCQkYT
sbvBVJINiI5vrZQ9hWs7H7yz+aNW2jOnKPQhafjJlFiHJzA1wfE3Zj+EimiW
7EU4NnVPocWCnRn7vdwHBYiRh5+1KY7EstxOAQtGdJOR60Xztb/iovGZPXqg
LIA8IV1g+Hrj3w1xheeVlENHM0LJdR3S2qKiQv5n4gGe8JiMe0ED5VQjzXZg
j+sXDs9wsHUwQj8wG9yQ2HuiQ9pDEeVw3FlfUFaSs0svlSeZE//Xz+AqrpAZ
KjOn2v3mcgctQPN3pvhUYXg3TrT8wyCDFxta6vxJ6kBaq37uVkymoWPUxqoV
bE6MxyNWsbmQqvY2SoA+ryLXIcvtp/SdjnNm4Kz7BHNmyVJ/MvtythKmcy0L
JTf4KirPHY44O+iGBS4e6/AO1gbDk1mQ0HyM2v4RdQytvavyQnX9MDJuYCSe
6NhNiK6d+w7pRA/s74gDiem94amy25NQd4DPfQNc0wrRRJ0/WLFtuccDFWU6
352UiARcOBYj4gsGo/q9zOgelj4lwh/neAHh59R8jblfqGtq/I1v7pvQetub
MF1mX2gjpp62AmbaRR4Z2NrL8IrJQfFhfhOfqp2ca3O29Suoq8fZRuInVb/p
nlrWq7hdg/y/B59YJjSbZp3VogoFkhQ2u8vC5mlBNCWUNV6HLkzVAJXREyqC
RAlOtCD3J2VzBkgpJKNEGcZBI1ajdSDkLbM2kjIsUk1VQu6cl8h3Qkud6mWu
hcrEL/cmeYjFuHT5AD+AtRZjWBHeKbbngtez2Ip9NkAWXKmz6TqtKyOj2wDQ
YbfW5N6uePobXca9oseUNM+EL1BQRcGcbNbqLDiLZlES60a6XhgR4yP1W+P5
ONwvXw0E/UZT7lUeNc6GPZPfMwExGTyF89WPIZ4YacS7UbixF4lDNfxjTxiC
E63vxYN4tHMQThdFhyJYepZMqhDyXRbBhkTaY98/5Pyd9vP7zCU+EmHM0Zuf
SwAZWN5LugpsaWzdeP6pWIZPcljx8SO+3516GYYtkRDVLr3jLWMOY7V4WKeY
2hlB/3M0+0JZ7nUgTUHcfeu93M67DpVJuoxOB6pc/fONspgOoILOrse6Fmiy
8RlzOFFo/UzXNLRsWAAF5Idji14ywiUp08WVFWapuUH1gAtFJxwRN1aW1SZa
U9ishlFZSukkSviBwuq1eQFjF1Rkbizo+UAFXzIZG8l32cPAkPa/BUMalKZa
s41Q83mUoPQL9duXfWMqDuSvNdmeZa3kxtHiZ7svdMAG/JL0sw2WSsgwQcDu
yMznueKOzy9JdkLuHDPluOS4r6yOarkcegjdw6rXNXleVTfHXGppEmkKaom9
/imiM9aPL/UsU/4pN4s+vBopZKf2DSjjtDUQ+gRyrDCOl3Bxm1tu08iWlT/M
Q9JLzGWNBvEjWtrEHRwMSBfq20dBXZlfvdiZQ2fpBsddGzahuMOeJdaKQOir
Xxwdu55m+wctIzGPkIDevMRXkfvBFBbNXoigBlCGpMDbK9+d4LWKKmI2Nd1J
Y4d4C8Vm1DU8CKKIiZZlDEKXE419LSIMy2HatYmXwBRSR2qyeovsykG9Hnwk
GMl49HtFU7Ottje4fsLCpaDwPENkjf+Loud6Aqd+zxpx4v22I22ik5UN+OR5
YW75cNS9nyXl41WqzGCTfXS/Kja3BqFYRP/7/V/VACGEtvXDc1OqIt7wyJh2
EqAhI+QgRB/3JCFjf7CpkblvMO1gK6fRmVqC/B3yTtdIPm/agFt2kTrZzW40
e8/y/yLwhDCgwa3X3Gfs+7liC6AO0G9VYJ4pJtMzQnPoK3OWyc00ohWKfJWx
f8EXctjGW2zUYrXnkflU+Sy6RQWcMxTVoXN3x59MiiSXbPil81kGulsW7Mwj
l46Z07VUBkz9i5EkSDplIBAWzs/y1Zx2U12CqY87xk552CGBdRIP9gm9qg/l
R0Ktl/0bY17r80EftZKB4XNvrUzuQY0kkFz7MyVgB7XZnLyXpMVsvONceuKI
W0PESJxvEwuRcScYra0/Z5OorFJiTUBp/0yhms5I9sRhnaUjSVEa9xqYLwgQ
wITFk7PkSleN5dsgEV9K/xjbgSVPqMRf16gUMuZnvAoygDMQPa5eKSRNxRTy
tcSzXaZs3QvQWQoSb2dyNf8d7rkdrJd4bEghmugshunPARw6IlwD9uSy3P1Z
bd3wpi85/AVAE1LfbjP5xVCTy2+gIQaCwpSallM2eS+KXmlS7aCQRMtQ8z0r
aZKx6Rqdfk3AGJ+BPqpoxCfAypgesNbsrleU/Jr9Guu06jOZBQa2FN+6YU/w
WsnC0x+E8eL0rpeoWi9yLjpclUrYA9NHT7rpFavRh0aLvc+87G/UDngsaizV
4bfyAwlBiKPvxgNhHGg0O295xlkEZstgC+Bdu8+f0myEV1f1bLQoVpUjieLs
Nbfj3X3jS+XMPt6W8T4s0n2Xc+0xU7LK6GQgCfPfhJL3cdB3L8VP9/ukko4O
K/rQWfy5pbcKxU0uwfdH+Dy10UnIN6pWOUrIBn1K2O06AmyDAWfvRsOiJz7+
0yI1/imrFPsyPIlZZIlzMUjhbeO0iTXTUTgewkeXcXLO7ByvoNqm4HTpzDY9
aiZIjV/oXrbZf6fOeb4mj9vDinexkTaIgaIeRK6Oj/YVK99InDD67zg+DSek
CSs2ykhbPH2gpaeVpgyVQNdTO3e0emVp3dB6hWnCXYPxOgm3lgPVznJ9W3EJ
uzVIiza/gBFuZNy7Hqn6QfEd7amTQF74O54KEfOFPQvmGaeCKd6hA7ThiLdE
7WEVfwm0lwZWmz9o8krS3jBgyiC0k/65Y+Xp0JiU4seVMXr21CoQmqz0a3N6
wDVyzF6/eUNaiRw+WQSzYqJ8487vTYAq0kfyes+zEbvH9649gWP6sGVpgjS6
fPvshpEz0HXH7tePxhv7viS3JgHzEX3F8MtWFVNrkbaxuG5QxhaWbi9zKwlu
jBjOAaOCKpi43oNiAW8nTgisk66i4M1pME7o9IZukvaTBlCka7SUQ4UEu5Bv
1pKDgz4pNz7zaUDX5S9z/p+zumbva4WE6wwp2safR2t/YMMgNLwnojrz//9n
hypc7iW9cB+caOOTNEarf96S8oro3unqJI98XeJEvjxOnWsodl/NCb8PnkOL
qSk+AR6xFEnhHkMxq56m2mOaAC6ioXHiDT85hIum4hZbrLEvm8BBasH1mNrL
lzGidl7Eh/VzoU8ICkjM1wVqLEeyGVH0vv8QMc/2WNJx7BP25V5rzi76qXzi
75pj+B1bEYKK5wqcdJIauMltRvRe1VK/lLa9IO3KVHh6ei/mfm9pfQIZnyPA
UfgIOoRiG/CJUk10cNAycw5evLd3/yosiGdpNfbZWSqb+OBdHxY3eWEN5CX0
ZjFVjDQ8Vd9MHn2zHLIQhKZCU2ddXP798x1t04Ac2k2dpAiU1pv9Ds59t6sD
Y2GNUIknf2lV6eTP8zLbdDN17n4+fXLE4ZRSeigjKUA2DVxn8qBJrtaINo+q
9x74K91hOyfKr2hVIokAEGbGc8oAOah3MQ3lPL9ck0pqwJu58YIw3ahKrmrA
MaiDbeR5SBd3rUbCc43RLZY8JtOIlLm0U7X0khIpW6q1YrMGNlwhSLeaKN9T
DAt0FM+16Ya0G9k3koE08zu3Sw2hF4OoAt1+Ngzpy3j0ENZrDDdSyBp1Tp/y
B2zZujZShDYH1Uwqf0T3EcMMDIH4C729PPNa+hgC7496JL1m/6fGGPTUvzoR
oma3dTC4VhBH1BgDrgTDM3QqxOXaxxxl14wyRrVweEMfW/FaCMeAcpI1JCf4
LOgub1ndtdHZiF5Fm3mYxSMnqlsRMkWtAsd5x2uw1VfMAWCCWWG4RKUj9Muk
6/JcGfp2aFB7aLGvZx+DXqCBRN/tXGbT3p9wthXnGDGrtTS0fp4KSw/CaoD1
gV5TVUAmZwvq40fbas/FFuvmRJyuxXQZm3ncZNescr1JG+SbLtnT0gFQsM2f
f8hrv0XrUiRD8LedxuiquHxUkcUnynbW7Hzm0uF+5DU8sEuVFuT9MIMEBgN6
X2D2HNdNbTOVAkTPnZyZxAZA2EZn3TZ6gURwIcNkGDTF0VP+g9MN8m0uPTiH
Ghp2KJPQGat010ELR0JGw4bs/kpOt5YB2adWZys4Ydbm/lwGs86Qh8j0GqIs
xafkZlmMoecOhVB3WWpJ+pAcdUbSp6FLJR2e7+6dZXzBKSxv7fNU4+UOi4SJ
JLNTfZUgjSs3wx/eP55VUccz31c7WXzMBjgiliF6FEM1MVoOJcFYRose65P8
MBq11qSjgrvb9sVEoDiryaNSvhnTlKsibokkTSosKDo6peEePlqqtpw+xYvE
0vaDC9Mc1V/xsw5rSEszI4wrqz5kC/yUP5jcHCZkhJGGWffi5B5VoLydnfCP
NG2PVNEQSPXmMXrGSznDED91Zf7KsF/dpxBy0QFBmDk5k22JEiIzXUnTwLVu
ez9luuqcMp2qCrfeSy6VkYCPdvRcsRCU9SkipxQFcsz4QHzWMOHiCs5redfR
VFwC0CWid03DX/qDigcOGcTdm7NIXv8M/uEeRZ7dAIevkmCWPLDgS3f5ruv7
YYi7Ezh3ipMlz2xgBpRjPo3TQqgPfHksA8dxsll2SZMcp4EtZnKWH3mhKP4E
IUam2hkoZdYYvvQ/9v9hpplxEIF3w82YspNd1jFttUlaZA5gQCxOalWMvHk1
ELALjI4LCACP+H5gb4XWDzlGJJDyzwh0ZU5Jbgf4v46WAh+KwPvKvai6G54m
LQsQnVOyDLf7xXvMn+EvDbenvRoUwlAkhI62m3UGCwUbDHkeKTYfnwQKg5uB
U4LyrTBR/rv01wPt6XbECTYONsUiaQkW3OqTXD61uyPD3LsOhuXTC1HK6cx1
6UodItNgLAYnxQgO2THMWeEjq2mMDGqcvoHZn9+EPmPuN+7874jlx9zTs3Rn
ef2Wrr8IyNb80WRHKXcr/k/2WfoETIWulYOQa2mQsGx0iQoFwdjpAULvCUnk
hpLF17QCu/S0Y97r3nBa0HfPU6X7FX7kSMcx3C7llDsLFPm0TLd2VORwoOZC
mE8KZe3viSBDDPM7xbc5GfKOe+wx17sf3eRpYkCTLQjWt2x3YUhHZvac3oX9
KZVw9GToTBqRZYR2Uta/tXvDjyUYp8Gr4gzG1nY0huZ892EJ3sLzPgStQB8c
TqTWWcFhA7JMrC4DLRuZ3v3EL2+d/CBypt1yxq5szeCveX+GndMNOaEqfxSq
TEAidlrNCaCLhtXz4Sn0LQU6HP1IUyg3oO+8N69jGGEmkGmqrvpB7BsKXdcx
9h/YXnsOk8jyw66bsC2IaZvzet6AfgjxsfqlfHUW17SvH4dk6wTUUyNxVwlK
gHK5Hn/Uzrk+WNkaZ5MXBIi9CK140fw+DY5pFoxrimVw2V/aFfaqmMXsY9r7
Tecr997p1vZJFWUrpi9w0Rwg8yuK83Rxzj7MmcQ/CftatWRer/imcjyXM52u
iSrYnaHnL58L4OnoKREzcjZQqHpL24m+oy2Cb3lADWETM/nni7g1kJRl8wwT
HdGQNll90gllvGqQPrOH0Da9Xr+aJ8QaBJgUiom13E7xIqtENwmrWWZlbpj0
F3Or9zAINvitHqBN9LBR8461FQDOu53Hsg9uhHjk349tG3qnZlXVVr4Sz1K6
/Ds+4DLfLNQBK6gbbNCAn6W7PnjNko0i8cmPFtOhMMAKXqw2wIUfUDRlkJNp
FoCJhGMzhVjyoyiqFV5MgNtfQMbgt8IJP2i1eFpue0PIiupvgNGEoqFzfEFW
WR71vcsGHA27Ex4JHfKyXGO1S57YE9VsFHD2P692p6T7jOukgUIivQbDGM//
puU9RfKmB8/mEwINHeadx1ctbak8pbKG/pPpGu0FCa2fpMKx4Igsi++N72cr
6A8Q3mGLxg7ktbBmxUWuN2uVH9OsupJMdyhyYCRIV029kE0Url+gpAG1yxe6
pVM1ZwCIwDSrjuhq1WBRgPaT4hFcO2bV7wFtE9aszbk520sCt4yySESYwHYe
WQQVI5rne90Y+MMGcHcer7ey2qXk4xrTM+Idm5DA3X+pXRgxTOuWOZXXGNyW
PKTt/4qpNNza3f7h4pLq7912cjhqyzZVE1GqprfDBxu7sHw58fASScEn0137
PTf9vF5Nc2bzD24v40Np9CvW5lZ+2Zh3Jn7Rzy/x96RX0jp7ev/wqNfPpWMP
I0MpquKBM7UD+ApWS1VMk/l/y4PgprO3mISy4f003iUXb32TshkZXZJVkwsk
9nRZDGoAVnzHthy1PcIj2Sb9H8ZGTh3eXnT4FjIds104Pwj7tk97fyCky/RP
w/tWHZ1/MHpQA/Ynifmq7l8fjvrSR93G+dsY/zWv6pMH9AD91xlem0ReE1Zb
SH0mzt1+jcw2pay7ak2H/bqvnnMqWmQfDfzgM/Ngb8uyDrBzmcEtsvupoCld
nA5Q18wQh3Can5VhoieBUcY5qwpUopkePazWUe1PkU5YOUh6kB7Jhxj25DaM
UDVudvWpa6C/Bda0bqP8yd/uaHtTxXDCEe3dhmVu4YNHlsajX7TUUYUzr8xE
TMWVRaKsnSULqkQHzTuc1OmbwSmpzuPFZDpwuiPf1g4f/riXs8NXEAkwZbT6
UL5WKGfBmmH4PJ4VlUgZdI66vOfVXp6WaQj/ksOvlUSqLWPBUblmucahVFIP
L3cja8QBXryR6CHd6+oqkeYLtNXdvJRjCHfc/Z/+CTPFXT4sT7ltSZHJholr
U7/miQHaCP8fmEXNrIup0wEveGCwIK1KDcHQHlEnXMTEHxVHHDFhvDL3F3Nk
cNUry2/HiqL1c+xbV/dgK7c7Q0R6e/4bkmbn51HJmg23LbrVGz92e1KWazgm
HE5jEjFVgC9D+QnJIPjrr0WkvEkriRwXFsUts1VTSThMBbrLXxZ+PbqRqNXh
MhSXjQ7SUDzGem7i93+wKBq5PXVc5j7jG2D4k44JWHkHCaBaJ23YOUls4u/L
UuE+pKcIvW+yltDNrCBkbLyYwCh0tp0Q3LmSXH/0dEnRwygBpinrelquRu+l
3PtoKNnzImHW6Zc0r1EqRYlwEVq8vjt1Sa5j4lwPemiYRUViWkFx/PI5XC57
nVRYyDKj4cOu2glK3WO7+lmGiWWy/rEgN6N0rKxm/b4ZjANeTrSRYwUYBtEi
RyNMJ6v1Sm1gM0JcGLU3bgKf5O70OaGJ+ImA7u6ksOiIiCMZSxK3FbAQHxDW
YNUF4PM/T4obGc4eW6oahfac81pwipan44AG956LETwJndVhr0k3hUQsYX1h
NTiVE5idd2e7T6d1hsenJemRlAwJmD5wCwaufxY0JUzaLxGyh4JRMK0qhZlS
SbNcn3f+dMZJywCdrtRTPCDtf5paMdVZ5Ca9Z7FwHnLpo6Ue/uWgbJLQGeeB
xCjDNZWNJJagMIWM7Za71O4ryfvt0WMRXLmPTUuO1VO1L2uv6ULOyxx5dtwv
MLWCcxymot5VG6sAcoP1iQZALeQMfowdSrjv/+99ipXPL9zWi1WGLWCRes2j
UgE45VnSMU+569jJlnkOSmQfQMq/2F8Wj5NuHCPhbs0l1lBpOMPjY2BLAP3v
0AZdR/0DDo4rFP/aUVQIcf/VumnW+KdW2uhGLo0tbK+C3zPsWg/L3bhYVIAo
9kGQUsOBxT0uFs0Qx3ZJ4UufUpxK1fF8y81Mg7PkyuGcIBQn0bpd6kJsVIpq
Kizs5otWI92/C9ljCcV92VTcY7wVZqbzEdJ5DUItW2yqiiIEoL8hG/lfPcAi
twC89IvIG3vMGfqERyamaRHDjJv86cGc7izr7+e78P1mMxZPMj4qeLt5nXpU
oZVnsmlh/ZAqdBel0WZmBGHCaPPGJigHGWlMCS0Br6l1EBe3Mc8okfGDg8na
7NT4S+odTgXm5LTF5JWLg6J/SfxXKioaL5CUPs9GdQfK6QJKUaXp2B60pAhq
S2UjsOV5251jgqyvic86fz/FZg5OwmdRWxRvO6zgRndyYBkUAhE7NCsTPqDc
i2Xs8fNQoNR6TdT+wu28nIwaf9Bp/Ws84XOZ6s0KjXafydp2AgQRT/neVCXG
5xNzjbP/o8o9/OZJFxzs919vI6nufN17eGBitSQcuWufAQ/qSqaG9o+ZGNRN
0BEeQ49EwZMZPl/VTt+zkPkoyyiEUgOJVEdm10XNiQhD8k5CavzenCy9zFzf
GVjeKmoYXtH3WDWoDQ7lroZFX91JAbTJYOSuyiIlCn0TqFx/haBptvR9qdGh
MxHwdDtRFh/9NwrCfEs10/y/pK9mzpozzDTerLdp2ewwKK3Ak512yznEJ2T3
bdQjozggRxSZT1B4dunX8Rib4FgbeQHx9RRRXivQB0EXBnEwmuRkkNJrscoi
60CrU4RP5aXErh2TN7ZgPjFNC6N2AO8kZKF7Sg/nVzIsHOK3Iiq88f7qjQg5
A2hWlJ6byKPOd3L3yjb5T8LbfCtl9gITUV4wSzX/gIpIwP4ZOVDcFINGhmn+
e5AAw5X7e1OnHgR3HVKYieWyVoZPa+4/1LAQnpFTLy6RWuT57Vdi274dm0lr
1ytw00GuAPKAIxFHExUPs5aDF7oLjki7nTuEeSe1EE0SIVynrQFWPuRRVItL
DkNjhP+oR+X2ub8xxE1cuACELt0CNagTRiolvkuVeJ+562eqLkajwXeHBZ4f
tx3AVnzj94u5aWre3vmuHj7MvjcjK1ubgMx2Dqd6qD+nMS/XnoLNA2Dgy8xR
M2qqWHss6JoGG+xOBWIjQQtrKtsVQkXwidnqtfbiZe+lYHZtzieWceW5Yqt2
IKV710y5YSdlFxQ2J2snev3XA6MHQadMPGHjmpNONTAoTlIN4EoQHrvB+QY+
9FRxp4DV9k4zxYX4O/lqr2Le/ifCJ37zt62VKLYb/gy1znQSadfaC9Y3qTwx
1ZDGwcEr5mzzmha+9C4pa3CbnbAxFKAPt3r3kWlyIgLrfD7U+3eR+55GwZZe
gozLTVV0Sch0tAymKwsl/jh+30D95QfUNqW9x81EVrtSqcxdy0B6hhpb5zlb
s2XUC8iDwvF09JmlewbsGIx+0gwmPuLwpiaO6wFLcZ5VEwbg/0YPPFQgCJMT
KcrUcXRzrd/4mFeMK1d3uzqpTI7hxsa8rGAPBPomJk4wF1hvHc1SUIu1ZX5U
nz72yBY2Yn/3vGaNUSWk9dLhSkGqoEhX7xS3p2kkdolqJNnLzyaA6YAy3P7Q
/Y4grIAQ6eEk18RL5Z6cVVEEPLgkWMlb4/LGpOBuCQUW+qIUXNPicka5G8So
0MD/ab1ss8dD1LMUCT7kQYkxoV/8DpndUr20RHJe2jSxkt2jq/FNSxuzZDDY
ghkLHyCinURodHkPwMCOwXaMF950iOMsSTb7eHN+ZQRar4E9orzOBjyiVzsb
twkj2+eTrf0Zs3AMciK3set7ExHop3dSjTMhtAGEPgy4kI8YvixtQPc/4KgD
Smv94BDA9//TjgEmcjn7LqmIh1CUrNL9poBpbQopg0pzw+h/ZRUBs6tC9PGp
DJDjzZpFngGfmrh4vK8SxpncnCQTQY2OQ5wOfoXA/456QFG7p3nd+glriWeG
PL1lEom3pUcd4E/x/kOXdA/dfq9L2hhv9pKhjXDTV9EeE53XSr0uwVY7Yd/k
H6raDE5nLplerYERXQBm8HH8/aR4CHkP89+dU525akH2vKy5PNy/LGNk6nJi
jG0HWNhdOVFCf5vJBGvDCYnlHpcXlAdVZaxiJ1DFfBypdvAMTqrkbqnAhAq+
4dtuDSKgc4fGezOcQ1k6dDAhc1uJb2NDrZ/ImMMHlBChI3Ycq2iq4WH3w/cz
CAprWrlmeh7jkWn0YY9KAgNbfO2FFAmgGzwPu0ldj8RYqD8+NmdszelD2lzs
vsd4zPEtHtSq6JXzEV9dt4ACo5M9hXa32CSTlZomFlE/T/qQnghSWVrMQoZp
Wmj8nW4fAkbmewe5W0027D/yZCuBBs7QAy6srfOAbluBkRpAdXmElvRYHDi2
Ld+va009coclxHGKAstDhSlT20EJ3YsfgeXIB7fu92uae9n2HJjZzy0XslBM
iTGi1tjVVCnEeaItMTFgDwDREwBRxOjsjhMSuS3ROsVp+nUhLJKEy6y9mvw3
za4c/vA2G41hlkyx5OpnDPPizs1+gWu3tIA2miKJdoWPRjjlRyNykmUPJNHG
4xU9lUKd69RO6+05bwZOsCMDpx6Lat51r/avq1OshkVnh3TdlwK+yZDOQgv6
tb17FZJzTD8dgbzDB/AUy8K2I1UN5r/D8gYnbKogsoJy4iYV1QEFZpz7Ga9J
XQWJI45IVXOSk2q5rs8FuTF15BO2KV8NNyye3lsCdNjVJ2FpHy0R0NzSfy2f
rBNKv980G8XH1WOYQ21vZp7zkb92VgCcE/ixD79nWQN7XYXKKQhtk2CnQXao
tQ9fOzbQdXQA5tmJrhIRccJInK8FnZtUHvnkpPzTvucGO6+8t7ZHHsxYROpn
hEejTALPl3AGC3OYe9/7KPNwuHPuKzZLs4/pZGs6JXLcHwW6920vs+2gRqii
l45h1DouyslNlPhiMmz2eUFY4ihHqHyHUvL6FMYEkZN4+cVbEH3ABGyIpS8K
W25WWp0LtgfCE5rmy6S6ke8osZtzJHY97AEqbdQ2SuxraQ4WQZBAX4TN6gL6
CGvbQXbTOdgCXU3dmQqoAf5hXLqmmnnPF9/T5MJQ5Jfsf+ukjRilmHmCrM3n
bVHQcPgDDwA3okXbfAqdXmY/q2FOPr5dFQXO+7ogYmgSDS5hWRPbuyVlOFpY
lDIQ6VxXTlcndbyUnZ6DcSUVOrU28VwIE5Bf5+TskzEpmqOSLRTIJ7dNEIG4
AwPE3PscOEhWV38Zy9Dp3RGxV8KpqBI/SfWossJqAG2EtstlJi9zmnBYOFE1
mBvdgMMnQIUU2W9ymFi0/BcIzNIuwlw3ZZN4M2BYTqO3jxAtG3bn77Ejp7+A
c2EUIWrjLKHmFkQMrhgivcxl9zHD47AYZ2+bnUAWfa8vLQqpvKKu+bytuouA
efoOZekZKdcBGo3tdc8xW9hGIWeT3W0AbmZSPWuseLwORsHuR/3eZkixdAqf
qwRNv5uRZ8Lspjv45R+lZUDkDlmaZ8Y7PCLog6IqbR8FUo+rIuZi5G2PClvn
BJLug3LFZp7JzcLWP+eWxJuxdUDbQoGhJlqomRMO2l2FOtKR0BV+sjDB13xo
SCgr4RkLRdD4lp1zFy8+uTa+hYoFSy5QNs6TkmjxYhlRUU96bJAx7ce5nvxy
xYTxMBbh5HJ8sphPdI+D2A0s+BreMN/6Zt4oaKqaff471VUoHPPfhP2dn6jr
/oQhXa3AQQbuOMOk3kv3ExRsVQVj6dgdAcULnRK7Kl38ZQqp49dMiUqtnVpC
kGr4SJJWkZoalY6BcNvJ4FJXWxy9u+UVhx4pnY+3TpvaAMxnzQlDXjOYvPtX
qB7FyyGL9rfQ8lwCGFTZNkY1GDz01cPqFBUU4KenJe81FwxxjTTVqrZtl7cy
oTzENHUgKGVcWbF5YK/r2GX5U9jUOcDCLyqqHoK/DDShde5LBVqAkgYUeORR
3+fudeO1HBJIib6gpcLnWHpHjc8C3iaVgEAcNawWGwm3YM9zI1sPe+tqdVws
blO69KHxEifUSXkuH4CJskoxeM6KpQVL/i/UIrEZjuqGF//XTquVRCZ/bzUS
x+cGiMPlaITZFxUlRdzR74MPB5RRWgYHqLDWZRTqUvfcBEi99uaFqWkAucco
OGTD51g3mdjqbpRm4lP74X2PSFCyzDQM3TsiDHCBxwetMOwa57G9Rv2Mn78Y
uRptqVpt/FsuV9xXH/GfSjb4PConm+V5l9kAEv5A0wEJ8wWVopOFgXFI55KE
EljzFqO7HvvtsJP+jR4fFx4EcYA+vFJY0pTOXiK95/mnN/PYZLjqR0ILrsDx
sqtDmEoHzMZ+V6cHOtgFkaXZn5kbYJz0S0x6zrefswNZPoWrkLFLrFCh9InV
dGLKp1KMhufcN+OOy0DiYOSJHPZf/b3+Fk3TMyYvzo+pMLEqtxQPWQjBYkyZ
dvSDqFInRDJ/c76ENYTBnu/q++h+SbiB4caAwN8gkexMIHuZ78PpbgrCnguK
ZhW2IV305Beionj3Luu4CpIaT2bi7KcHIA3me9na476ZlBN4kmdBsM1b3Box
j2KJJBtj24YusfISgfZ9Ys2b/EjdZvmnT3Voh2kwyHd6tHBqN99dYmQE0oVF
1Hsj9CxxL0ivMYXiR727n9ApQkl2jI1MfNOvc5PC2TPI0yuKigeiBRIXEEfI
PYuJxylhBjE3HFcrbjFTrYIGw/wo36cQ7ZRqy7tet020MRubneqpBEbO09rD
90HlAvUSCkym/66r99QrML29xji485ixP77hA9NoeVGUPQTQ4PA5Oy7ljV1O
Vr7mUEENaIcwIcmOnEDeHObnCEML/d1HXyo/GnhG8pVQ4xnDbGQRBb9Yu8Tl
YY0K6lz1MaBXA2dzC64mQRTOaZfjW90wKCWGZ/2a5l7pkERLbpzchRx/qcCo
EMmavGxqgDFPQFQ+XpeVHYyFgVims10y9ueO0Vz2rRwtzSJo3dvrqUOxkJJy
gD7SEBplstJoCNLTwL9ru51RBXPlkvnaiBDi5KyUokK7vofuG/9Cze1shjIp
3Px+nmjTz3qH44OhP9i1mWwufjRcOQfC2jgh+mWgSgsAFKmJ9gNUsx84ujjY
ch8GByNDVCWOv8CbWVwrk43nl6c+ZYALYeOiqgxXtJcw3NgJa4iA5dJqRNqQ
O+QfzedhXvZ/92sw978FTo9iyrnL9ilMJZoed7m/nORJyqXWMPAEhDjpQghl
GxxBo6Ehi8VrXU/ehKD/Q+4dOJ1+lF0grP5dFOK6vGl6kF8IA1bV1zL3mbCn
D0PO1MRcNtImo+kidH4F7QVrF/NCKRB+oJ7DnHDZzQbHSR8pdrhTgKKbznAR
eVWhdJ96CQOdcxAUIeEmHg21Jxd9oHdUzipxPHT+ZmGsARwEFBFZGY9cx3HL
78QkdCzQm0Lipx/GPu2iaXxZaszFo2ui0xZZDFqWYTQb7+6n6OvoSf0w8rK+
GZFBo8tnPiSEiOiujYqtvKto5XMl3arv9AqW72DQ/3gMmBdC+HeD2hNUs41u
llXDYxBjwWqSh/NZlPvKIOYItLrMi+QJ3cJ3MY/U1UwzxghY5lrzAnXNCrPa
cyHH8sjHlK8RxTSjIuSXqxMk+3xnLqZn7aVjbTKOfnjgpe7sIijjCjVOUFYZ
2zMbvxT2HKR8s5hzfZQHg/4ofoA611+7IMYAFKqpiyt4AVgXU0Qzqo23m9Ap
qq0Ybtw4h8GE10Tp3fun0hzRwoLbEr+Z9b3n19zcrGWLAE7+1dKKZow/hNK3
/qgbn84umOPi902kEt6UYMkADV2Jd+f2QjwsOoCtBptTH9o6RHavtWOaY0ip
reo6mcACLnnjKYw1FFL0UID6HRhiNkYy6xbBqvU4nsOksOmuIGCsEhlLrQzK
6FP5MgVAs5Ergl1A9tYD0qVKqkH14ErlvyPfR/cg6NUPbcLIp/MpWJvEQlpB
vf+ndEqf/DqpvYFUMdUBbHJQRzcImSR4tfPnXH2HcpT42pHhQI7O+TVEPv0p
ILcQDamChROvfKF1i0RQKJrZUku/PVxhAnRij/sonXAYGZe3qI7hoDyxRcIJ
7L+BUneDRCtUHSEOGsLsnIKWhHsuH37w70K6PuzktLKNknhkOcYO8efkr0HI
OqsBf+AkwlzTXkpf1JV4LwYjA2mqufo4yD8caZP/5ah4qp2TD7wyeCFlJzJ0
I1Yn/k2QiLfE64ZkYPD6vMPAJbywq3MyCGUSf3WRmN7AjXC2EZdpI/xJevXX
MmCJ/Q+a1SHUvG0k0iQ1lhfEzNfI/lcWUs3uM0vb+sIPKMFttFiKSBDj0ECY
FarZfMXNMPy4VL7gH619Bmjzc3+44PL64lVDi25BZ6oPZAnU9VzTUpGKCZpM
AwM0XMdm+e4jjbgT2TCrABDxVzqWKOMMtT6VUCaFH4SahFEpAbzYmWSlQXss
hFMHhOupB3cPP30ncW/tcbhylAduF4BAntPEecqflzVK/IAcWMiLfJn5B0Ry
gOkpK06+RVxGeCumBB1VSswnUqcl5SQieo1nzIWwAdwkFi4TwBZnVgM/Xh0s
VrPpemZ2wiXXaFJ5UY98UpPxAhs0OTOuCWripMtw48nvQGveSDVIEmCbY4Kl
hU7Jo6IQlKuhJ+AJV27sgkkhRkZ701OBjqTXR0aJt92gsoeZNSILV7uxufDT
uDGxoIpZ3pZ5lbbnhaX0E+nwpsCjG4neptiuCUQIAnh0SXmrNzkgO9ZPzbjP
UY3pCXB+dux2HTb8g9Rr99lvXEvYV8HMBOF83RrFcKdksf84HUHsayA5j/K8
Fi0dWo9qxLTbFYJILi48F4SCNBNehctadou3J5+WI7IcMDKfJWIY0Ppd+BVu
q40vXJm7Rq4HJWLM5dlHeUrFiOcYACvEJ2SH7Ujyl7Cstgk/WwVP8PQs2rOA
xNFYRLN+RuJdsFIU7Sj7yGetqdEv0HjlvYuz5RD0G+YHJWe4FPtabz+vSXgq
ZPM555fHcdHZwqnuC3xFZEfZODMR0+BAYTmWTt6sotlnpL8wd4I/ipP4E730
+4PCrrGYCpIZdmSoFkv7k1X3NxIhfYepFozI9/5YKKa6RwF9QFtvnGrlVfmV
6OgPFy9R0uoAX+80Cm+Ye+NHbIbl9niq3iuMhxr07Znq1yeTLL/RZNk3hzts
S58heWYzC59BQSakNcqCNDGTxX38khdF7dvZn0bgliObdZoboPPJ3NbD1Mkq
QuLJpcksyfWw6jiyl+PfLUWg8AAhDr/yBWg2oLQewWvp0YKb+OPLizRGk6hN
RrKP4PmhqG1Ci0wxMw6wZt19BMHNqOaDxKMCaDDirLKAdFH5KGz4w4rro0Bf
nsGrelccInM9OqvE1gRaeIjTFmxaG3ek4Lz8FmhLvg9U/F5m3hXwwQ3XiB8t
sm/m06yZgcthFR+dzUU9UziGxyWEqM83tvoYmqwC67D1BPjvFSMzdJZBOKYP
J4geRgM9NV4qHwlQmvBe0TvySYGohGhMtEdWw6JSrAW6P3AXhAuEfrLJ7mh4
gpZXiegQVNFizcgCUoz9Arj3Je2gNZFxz2d3vvB23yZl/6rJsv2I8XiE44sg
ZvPo4D/jDt39KVF/Y2kdM/BHEYkKDn3piiqS0Vy0gHN5bbec6DGoDLQvPV7U
bDkSwgAcKUyNKVf5caVR8Qjkm71PABc9NJlPKocU/f1S1GWCmGWQ50vO0qiz
OXaGoEXw2FTl14S5ezdEACvB3O4TNJEM4b+pmlzvlYnj0H+TuuitUhJa8nv9
A0YHELs1MsEzpvNR7mplmUoMm21CaScdhAx6cNb2HNFkjOWl66UGDPeLz/ju
K+NgQoyNC/EsLTTQ0B/FFTaimpF8SBn8hqMtpQIqxlPW55YU/Fklrq3ts5ym
VNBVhh31Oy7uXiQ0jSHe3oaM+YKIGNbxZP8iLe/Wx8cYXf96WY16qRD7CCcg
ZuQgykXAJd3lJB8ty/QngDr5b4bVeklGjlHBc5SJS88e/MFL0R+Vdn5eANEo
s4wCJFedTY3uin7FnokjsD8LHS5q0S7HNVo6sCoJ8Cy1hkkkAnFS4spozlH0
D+F/5LbhlycW6LttVR6CAAJfAVUyGg0FzATfZODXqs7gTAJ14IS+h7G6eSBH
SfplR1sCJBox1RD+1LP9SjgiL0jFq3b9QE6/gWhNrsHY1ePeX8adiKOnSf5b
p+saEkoqhbp50whLge4f/Bg+0T6GBpVYTOxTnO9boRzKRiHMNbZLRBAbX6y0
7pFgRmpBYLzJu16AhaoOTNOKY3rsktU1eiULupYhMD8LVY3oHaBGKfuhoNgY
8E3NPJSep4EbGEGfqp2kzWdZP/SZ+4TOlTCgcUX0HrdIIP1AbxhNnUptELCj
gEXPEmk67sw0XSO5PiXMysrq+aaQ+ZoUHaYJA0KUtbsBvShj53tb6TAljpP0
hvNzBknZGlnHVYV9CB2Ne9rb6hGTVC8N7WWoOepA5tILJ8VpH4Ml3unFWY3q
Cvl8bFDdMhcnf0+gn5Ex5xPbTzhyZOYHZQqqInWK0M/gPEZt5itkEuNNd/9W
BW7PuuK/67N2IswDQNLEGcIDsr+vVEceXfVjQNMZcBWLKqNamUPFNWX8OyAQ
wrgkyx9MWmUYux7QAgGZgihVXPLxkf12yi9rpCF3UBS+2QaY4BYG/KVP85dF
1WFFLhz2FB9hyt8r/V/qr0MbT9VnNNMc7wy0jeCDLmQBJswX6YxUbyw5HMhm
34yUEcH5CdFU2yeoUt4SujDZc7n3KVkA+Z/SOxF51UzIGEgkuKdOOoC3TldL
7ySsHlX31RiNlDUzhrF4XTCLcnNublv5oPSUQmRBth9wZnDt3crXALcwP2Tx
AeKxfbbVSDEcB+otQwoPNmAXp3fiLhBD+CA2dZuo0ohe+jtt6Gf9ijyBHc1G
erdvP4r2VN8pYfCuKZ7XAFXX7g3CxbGhus4hLc2gQ4J6RFRa0dGg3NSY1J9U
eXxPCCzZnxTKktnmS2jZDCLoFBb9kEIVYKIM6uwnPGyEaGCXjlldDxKxKNIY
68yFa4zd0KMNnlOWzaX7H9MjkzDrgokKKddx3BpeHX+hcu2Ylog7oLwADOvJ
q4d9OSkEXrcTSyGTy9yAcAnLtZa/MrIdj4T2Cl/LmsXbrq1MuCGNOErmWk9S
9NxIrQe9BTMFccbxAeUZun8/elp6kkrXBzQMtIlR4zpASprehtj1s+roGwg6
ce00Nq95Ij5wFufBnSr63ZgYQJEBc9alRkZNwRXcRD4ZGBo1tsHs+z5S5zZ+
xxxz55+XF7ZnGDkoBWgrDGjCj7AYU9K+LonVr1bug0H1KZlD8TnpYy+tvC5j
rC8s4wljjvFbQTPWPn27Nrn6OM20zwFgJOCKVGpaRCxagAq4RjcbUV2viCB1
78rcts8fha9JD0hWWBsWraPaLpK5foS++WfExzJurPDNkb+xS+k5ZdqdJO8b
fbkCCapOcw1Bg3qbAXw+PckXfdxltPd54fz6BgU4tnFqsF3nCnL55JZ0n49Q
wXf4N+Oaj245F5FlivscbKOhhVP0N1aC5YOE4659rXsBpPe1OR7jLt99oa1n
Pz1TuujG2qeY9jTmkCXFc5cegkNugQ61YMXBG6mZLaGM3dEOrppAXbdasrmd
0YEv60gpIoATF8zEGzgva2BYj2ygiO+kPXAaQfwrmVV6GH6W1dx3m5cKszQO
8ox8RFyd6vZDHa5zuODRxErajJlHVmIlTB9qvHyLms1mTYYQdaFSPW4nsTRE
W8enIGkk3Pv+HaBfFGbBRzeajoBtjxXiIAneda94peO1ccCWXbU1kr0g7zI9
3bLw7OpDwIINrhSE6Uvll00TtCTU4RXHhhyF/kSh/hxKu4PVcbkBB604Q5wb
fau70tjEhGxm38G95oVJs0V5WIwpLQ4PJI/YLMqqlIpmUwnKiUyiTV1meiIk
S7jUwlOHUhRi1RJ6ujmptOx27Hgye/NfjlNVmb54Gc3F93LZDavvR3IKDCtW
FDDcrtGUfljkHVlcPpcMYxynqJhZWfXoBcQ+FbEqdfk1E/LpUpM0mYmo1+gR
pFQJeypj9iXSUHYuKgxXTTgtbtDQgGl0VJSyRPyXOHowhSg5gHbRbfrDlCd8
8OQwrOrdXqV//MCIaTA/NwouGpzyy7jVbH6MPU3QN41qGcNnefUFZlEAvujw
QBP5dTrCVguu6zhxLrWUwK8wEwfZBJ+AXrhin/hk0FMiU6PBzXoy5XVQn/nJ
5UYCgjgQqRHndheVJ0b5U6Bu2+qaOsS+OLrbzuNMEQPGH1dsCMSC20T5WVi1
kDwrxou84jPIE2d4bxrb09w7xbLR31GA6EfTBbWFlKPdMxqipy+cPYnsP+43
scsQxMIsgKcz/QebmrwOPxViuwtfEAFdIJzc/txgrSGXB1ijsAAHRToUrl1i
I2Xi1fRMkhnLyVhWpNClrPRGh3GIHVEejMxHbxnXgLxCsFR++/PXWOsc3o/L
76MqQKmoZ/qOwlsBq50POoTOg67uWi7VbStFlTOPnqKRb4nx+XPBQUj8IwiO
bRBGOa79G4h/0s3OyvloK8Bx1Il1D1nZe70cz1PePqvaSAOcqvC5vF3ZBB0R
V1zxl9bHFeEZ9R5qNWlNd6xe/Iruaz10bLV7IxJ6KKjotum3m43tw+j4QN8V
lSITqOXTJrv7LtzBMX/UnNk8KDxvwScYpT1Q0KqIX2I0fkt6geJ3s2125HM+
79x2WgdQjFnQ2d63/7wCIGP7LpHfpcvN+bauXJs4S+iUMvN+UM8/fyipf2pu
VExx1Piu24LtqmtLvBxnunGWtWKMEmtbjW1Rtb4mLsVkBqkybpg9IV974zlD
0//25Sxp6qI7gFokP2PnyB5h3YkJBcOELBJgk/VXjAaso5y9cne429VwIrtZ
Y8mKn+ErUqRVDZdx0WbHtXIpm6xBQdvWj2T58W8qm8fad3TEEgx1dhiegfj2
R1GE+J5KwjAQ+FYUBnbWgoiYYGOz4ckmzjpH1SOp9+1iWgUzHMOVQMEq9P9M
VuLtyjvlBOLpYxxm4CfA5QlCSaDkYAVqWRVlzFcPiAJbUHHcXvKr86+9TUvB
UTZVWsznOuLpUvFOO80qhWcsrEE+6paK5R1loANK/a7PvIbfuyoPlgRBFYB7
hngYy/XkeWJl5+M+HTzUhVLOyk2NsIKkg6cKcmcYMGPXI7mC6PFciMw1QnvJ
p58Ky5MNAS9KGEvlmMAz8AisB2yfOjRnoVPDtwHU8MTyf8i/Kg0Fm1/2djr6
4vKkGVTvcBM7l6Z0OqJ/K1OWtstgHEhpBRez0bkNAgQELCRBxUVN5zd3Ieeg
SFMeCQCV/zBc/T+H44a6m/Y9RZV4b/6cPJTKF0P9faR3KfYlXpm+v/R5/YH9
A0clLJn7PZ15JuYwvSG5URn7rhoQBSY5R0H8aUyU22dUUGU1Aec95yXjwYtK
PN1NLlDmDY1/F2jSe9XKjS3Xm12oKBXRa6patjecnqzus6ZVQDggp00P7KE4
bchFZZ0L/5nIdrzC3Xbn7mrInnASN3ZGnMIhTU6Jo4DfQVNCHt99RpNWexjU
d3zjhWWnrwWT6EPlAUk5NrwhdkEDndga3W8Lbo4TumLWHVRfn9myeaQZeh/s
rQA1zUGxMRiYKCOQDNcCfjyQDzaO7SdfKl1E1by2YtEMphm91zvs8iUhIf81
LCkL6C18J8s64rQoLCDiQTX4VzuOUhHT7DuX6JZYBnGYar6rj0BlPa6h23vg
WCU+IQIhm7KDC6WBTrHcAX82/nlY8DaGv5FKlKoDFyVeNFc6y3R3jwe1ymsx
yU6VPyVv/mnqaEqyxjNSxikd8RixOb26UyjNfytQ/ltE/tfL5L8M25WZ9Fbn
XDssigTu7sL6LY3r9wPx4KmaUdkP3ZEWBmA2Om2bn0GiOmd9IRrbGU6ZcoSy
4ZFfzhnkctgPY8mJjoG7FeOHvM4nsNZ9T1MP7jJCnee16jhyeUTtkc70sbyf
XdM+IVInyRGwnlatPHBI1x/KwEEBjLQT+b4VWONEX/nBzfZ6L0r4RCgs8bI6
W9ULt+vrx0m61cHyDz53vuJe9iLdYU6JcVPjyb8+U0qitqOWTCxX4FVr5iNr
I8uoWJxGChBjJ1eASrepgra5b26n7g4uG/F22YE9LcZWId7ukOGUUhrlJM62
pCfZYqw+ZVNZdgsghbEB02iuFehHqrJSj+FCOIIHffsow+NSsQqX42qWUqdV
qv0eHdmQAHNdDl1xH3aTo+gEfKqKtJWdKEQ8LQGM387mc91xyWtc+nWOw1r4
FbL5/l/e8gBqU5IqeNuHWzAgi5RbebILaT2XjSQLpwlrZ27vXQiQi1Z8ViJf
Y/627qXD3RI9x91SDon13Fgkj4toKbnrHJDqdEo7nWndyZ1WlGFnI/JVkmNx
nN+RVhut9Vu3ZnNtJlqMDNeOBfrxTPs19oxUA4zCIL8mer74RVV3ENT4U6fx
HYehRSUy8ZCfwiGDv3VPYFNbKJNlBPwf0MPQGzRq6RhQozu1XMNIfyU2g2Lk
cPMYuPdtMgDoCQdC3CBZH+wBFx/qA03MVQ6pZ9C8J66VQqbWoPuVYXwlWuBf
gtVOEkesQq7ZcxjuRoq1iczK+MINMEnyxAPIW6SrR8hMRWD0wDWhYukgF2Ah
R+W8ZdPWgsRp+EdHTD/z1yVzFZyuviROplTlcfb7N/9wRKyVqcgOk0pSg2Lb
RUpswN9I8W/AvNeWV08gE9J0ZKxgirdVQ01MiVSx+tejV7I/SbydWPZfibei
B/GLfDjOBTj2986vdehArZSNanF2gXqYO6lQEn7SE/ivPOKk8kUCDAIEO6eE
8F6sJ47wC/wRHwxFwVo/foA8f5G4oru8QtLT9uw0/XW3HQKY8TZLjJgtJlGV
RJrgRnjwwxLg527ZHdGWZyyFsinVfvGAvtLa73sBBivX74H8m6XASe3FZDls
waSUluGOM38cvGfofmYoEs46jEDyNEefwrhJwNxZQU9R1V0eq5vmWD+mtzgJ
oF1UocBTBqqUZGKe8bLOmoKR+Wqgt4l9WL0T1J1sABYz/HOEJRv4Bu550Lks
fJtnPwSpSTXi16Y9rcfD4QCljvbM2hyvDDxHyq/GwYO3ViI+VtcVXGx3kDSN
5puNWUD6zxEw3A8IynFgjF9C+BYAS7oPgJr5xXUSugk3dPNyyXDG1SIcd//0
I3ZouO+gkHbRjYyUGUodop1CmOmvOCiy49/stFycKmYAOeZxS25tymt6N0vJ
r7IJ/4rSoB67FTSbn1CwGq5Pptb8Ux/zvrcHZCBDmUPfQmWPWz6+wY1a5uGd
w7YIqf2JCWJKyN/xQp0BHRIo5myUTuZVilO1hWCMTU/yJRtU13GpbjHVGa1o
2LAZAmAnR7hmjvupwT7oUbqJiozGqXuTi/8g99V5B18q22cmEu37F8uxVXf4
huMN/WS6XvFiiZGA5ullFwv70jfsrAdEKUJYTIh6l1RoHAzn4aQGlsfJMDLS
xoa2jHqeTMwmFOjdzf6MSZxSODfgcBwzJLZUixkOK1E2VkvIGG3+J0Kc1aeL
nUhcXj6sYCRfF+gzdp6fbwrJlBlS/YJbZCJdLX4iN5WN6cwrPTgFnUh1FWj1
2adXSISANzFNXleXNgAs/XohotDVsji5kiGwE8tMKiIwOdEO8jr2RZfFHybU
gpjdIFDi1s3VXqp+psNRPxDMcamthtzHl9aK6WOhCWf9L82xU8DlU8Sdw/oE
HsRC6D/K89D7zETI1XcDHFOq1fD1is0rWr2CbLHvHqWzDA+/FlnwoDLuCLi5
qPSZ8z2/aFSXbc7ZdND6ivI42MIHdbbVuh79bmhS+Max0waIrnk6yVwWm1L8
7teCVKwRo3qU6hvfCjv89A3nrJWbT7ZjabYTm7BxLiPgEqX686+K7XFYbFsD
ckWaEovL6K2/SAl/vKtrXJA3rfn63M5NnrWY5NgF6GubQ2qvgDKuTf/T+pGe
gb8TIp9hEZVsiTuutqKsahdtbFexlKBsCWYye/UYkYYGqaiyPjJloduzS6yc
Y7WAn/71HenRm1vIZrRf6wBZJTh1KExOHs8HjpzrJ8x9sluUMVGb8cdHlPyG
H7j6k1Nt64FC9hjUIsq7eYECvzZTDLqBLEya+/hdCllk+A4TJYY3sRG+CiU5
FQigu7+YsEGHcHcCzZlhUbU+uB03cmO1YTr4SoMvU3bDtR1T71waPrIfXXYn
f2jFMs6E91rtTkJSCtuCM6z2560cvJjjRn4TMJ1e/W47q+mgbCgQQLruxKxM
h2RYKTYC6+7M+nUY86g8jVGJ3XVMKuao6u8qOjcK72Q9fyofchJHrd4fW1wl
WLKNHhK26+fhVNR0RqNNNBQf1LZR7rk3RK/8rmp4MD53ip2ByutwEkZLeFv2
kmpH6s0XvFb8yKrX04swXfT+44/ApJAIJZvxnIDgLhJliQd4s0GQk9vSeCLH
6pr9Wk/UHS7C2Nz/o3DF7EXAdvToaW0+cSaz1A5Tf6lWILd15j6hwJ1E3EyX
dSQhkFNKkQ7uGzPCDBrSzrr9NdsyleKc1iQuq9x1aC6q4SaAnOr4GE8/PkEW
1SsJ7E3vaN9Ymufvbp97/7mU4lwxaNWHJXa/zTqyZMdfg+6Rod0jlkKRJtGK
h9eQB4A2MUWsAqgEfEMSNo7WndrnagQjWHr/0ah12o46ivOLMMpq9se/YzTh
j0IAePyqJFuRiGmtY/iCOGiZXCuk8gh0Wys8q5AJnipsjLfN0Oue7Wip41D4
BMYNpgseIMyc8le04ocomMZdFbqNEXBGvr4+oZuxBL6Z9E76rULJxpTTifwR
9SYZARdpEamLVkHqIi8n4oMEgvzdfmN/uicQEm3XmyZgiPFEy1I15jY/VpC4
628MMF44nDmrAjQhtMrlr4VDlPfmTxp0Dg2sBpoihv6oAvU/U2/pIxAJMdR6
z1T5/nHsu1NFdUPGJm2RSsjf/zFBYtX3To/yBDjqGesa1D3lT2XPl6fAzW+B
GXAndPHXN1M5OI0BtH+PMC7ztwoE/Cn80D+fA2bRVGO1yQxH/aOLLh2B829J
3DvWZ1K6l42A/VWMjqOSqHvlo80wV3aulDDmpX3w6Uz+qat0qb80fGvZszHL
ZdgdjnNyrUgusgYuEMgfhJeEB6ymDgG0s6kYBYm4YAPjc0/ZngQZfZ8ymd6D
rlwUz7oHzUjtfHpu+D7/r1UZeoQeWiCi9KnolMQ5JuQrWvS4e+GdIZGDNqVy
tVXB6iedWVhWN4T+2RLnYsbRLHldph2IWaHGDu/wY9qjjteX2gQothe/aohR
rA2oyo8pP++X9NyZVYKtmH6mSTVnRYIIR8XMxQ/8il/u0ZWL039qRoYkjmlU
Nis5NrDkhudbpMRysVSEN1O8ud+/7eofTlCa7VzI5XIapfd7pJBzV3gQ1N08
cilDalMa6ou/HOd8IQ4I08vscxSsQKpoWpZo/PcCe8FbytdbDxY+FP3qJnkQ
WIOCNjewcxHow47xy3p5hlnpMMuJG5HUZyVhqyzyQDjK9Nh6Ptt00EgOkfwP
vuwahN+dx3z7SEh5meV4brIIaVzhHI21uqEJgFBzNgLiHuTOpSrn2C5mRLc8
bjB+oftdeahzFU0vaYB9BlHQwnYwI4p0M/mD+k4CaQkiGmB0QmyWRp2dgv0W
mzbncAd3GtIlTNzQh2kVfjfzF8SycC2SWuUs3NXycIgRjOZPS3yl5R7fMrsD
HyCmWI4hEim02G3MNkfJ6amFHqitm74ns1Mpxokqaxb5WKATd1vJ1LGrPfdV
41dDHAJ4yIFkOoD3AN9E1Dig2CRfCQNaX4bHEdDNkT673Ko2L59Q+6NE01bd
5EtrwflzLo3rW0fJPlafghU/u3Emc54iyE1No3vGTzN5le9ftCSUYEtiNJ6O
TvfFK9sEpRqxbsF09nn8PGc3XW+Lrt96nkyc6/PHlFmS30H5LGX8HuT2+ymK
dg9L/l4j9OGUG4kxfIXGwQ4XDMoxx7oE5IUtQ5M9hBxF/hZcBDVlkXrnOHQH
f1VL3EMGS5ZlfpQm71b8EYi8DbFpUZZ2ZAGtLQyynqF8eHiU0rXMWMaxAJvR
v2RYEb5Orcm6enQfvit8snaH8UBqhvTUG4r9VH/zK1MUH/NjgGxIjoV/wsCV
mrInUlJHXblnkl0nM8gyY3ERxPO92Q0f7JXSovkVsVWSKR+/VTqdcUZQR8YI
6yrS2D88jsceYbWlSO6Nr/HSslb8GYbEsiF6f0e/IOuxWjOaayMo8wUsrY9X
porUrPllWlnTPTOLsOCGAzDiNYbkp75slQfPJ8OSp85cyg38JGGlSWuZUit7
QH+WSyVOBWxk7bzF2OmkqHi8ag3/5IGep+GsnSVqUy8DToV5PjHD7obvw+y+
2RqDu8UfoC69AzkgqR/ntn86cL372yEY1sE7tWFle0fpCu9w1o1C3BW0bloT
/3ugiV2nyRE/Ot40cAUPfA6xAheByAfIyYtKG+UUECndESXrdeX5hjfd74A6
6dX4qShH0dRhCk9UFGDtqcnOrPbr9GSup0tPS7r2XgaZL1SXyCvKTcJbOy5h
sa8F6I7ncmn/WSLTCaHdbtd8RFpsCDO3THu22ZxcCK6/yNG/p2eq675/Sh7k
2YMPn+NWf7rn+OiIpS25M5CoBj3v+ObaAzwXG4US/OoNnvA0u5W4BEGaAKZd
kWMKAzrIj6QqfvtVba0/y5x4kKjmquxgDQltEZ5+poosQFJfdiDCWTcrQyqb
zZSuBHGZmLnt5J6FBP0k3mYfmLiCr3dSmQvIlakN5QnpgY+N84KyioSvA/m4
SVpjCsRDJko2A5Mosm+FAkfGlauw49FdUgnM/rU2ztRCgkUZoi0dvScpj5sx
GqvUQXS8+2U27D+Q3UebPiCYFW7Z6VGenZG8X4FczXiej/xJPe21BiIRcJ3S
zu5Rm4mqIkPtW0pm0zX0aWFl2/NtRJa/fjm/KvNxKft65nuNPncVavXhH++A
tPCnPlzXOZQtvmgSm40j14CLQcavNwMAPXF1z1+xtv2ZSk4MP3suTXaxe/I/
N3ZkGXHUnJn5ji6lfkSZd3EUVZbeupo4b2BMrAabnogxQFxXjgCqkdZugoYK
ULn2kdYoYm2zGdeSCZQIwiFzDj4a7Gz3FJn5pPA57aoWvEZ6dE5vk7kKPESN
2Km0BVcZCFBBIvAmkOJW1wrmGhK2B4+BT9ncitQ1+jiX7sD+wTX2aD+NEpBE
IHvZNIOBjMyKjeCIZacJVBKPdz+c36mqNid0noM/5u3Wr4xW1/wKqkrpqWmU
rdJB14MsPWw7W1DPH5RbRO//b+/C1bWBxjDIP+uKM6zOIYZA+cqxXawE6ybD
nlObwbTZqhC3GrSP0wwTwVNbAgI5v8tBB0VRkFxnJH6n2oZUuNnBwigKBMtd
zJo+HSkSyuj003MnvnmH2tvxbW7nQ9Zc12fFbLfccwPCsmVJm4+5oILUMJ7B
hCEu3PjpKGef5UzTVHO6tA9OHZD/zFY/c6NRjn6EpCkdvnMzNxnWWqgHpt4O
rbrCxYr5FDIQrwdJp530D4C6oQWmNI+2Cy1ouo6RlqCZ/uoRoAn1wUduGKwZ
kOPfMUmY/CI8tbg18owfJLdEWC87RYh8J9U385ehJHm7kpKYiphC6PDSvuFy
NadYsoRtXi9f+m4FLzhJd69ZziOsrBZVeIjSnDRYCwhAXY1HjRgurJ+5J4qo
Fyutm0HdZI//v7UJs5jdnKLm1IW9EM7tloJVtPYcaEVQNb189m+ronRJsoob
gHvg6YSkgfpfhETZ3XlNWDIKDbObSrxRY9ZCmvrd6FnWfUMY9iEkRM3FzQ0y
+cRLBl+fyGuH7nIHJSiAftt+go7Klf3geBzKWil2FXOT8wRursfB/FjMmLvq
j6RMRj8ho7yZD4AjNSAZfgDaQsVWKiWUD8uktnEmI0pZeVSxb9Zrvi6efYe5
RxRaNAJmtEP5N2GmmERLhM2UpLbLpeVV5eVPOyvh65ZKV0EIOC8temnNzRcW
jSoN8nS2DLVmhu+ByfephUnL5AKiz/Ke1vjl1E2L7BD4/bcKwF4SYlWaKTVq
EQvE76tqvoaH2LfkBpUd1z68l6/p3h3o787lzxZ7F5n1J7M4P9cE/hBr5Feo
FvXZjG3zzYKk4dNteSYPdGcGWDxSvQGstsR2OfmsIx2qY307nKqTz+ZIHTC9
AskoczGIQcqarrfsFxEWzoN9v6+U9x4IMBqY9Nq1jnCk43nWwR3uvGMZtoFw
bmwqhQ7KJjh+QBHKHPJTRNcUszu7QfjJRzTTwzHBgiR4apA0t+dFLQmCnrR+
lhU7dJDeLpMWDoIuBycIHh5x/RfKAZ2l45UcHJBWU9aD0Te/Bp70fvnsQ8aZ
BMFTBhkgy6CwJlwjEv6P5/Ub2Px7Gu069nejjedma6bXxjustaEHYgeNVsC7
ExB/TbXhu7PcJU9mgtKBt8xsYGRE845LlsmDBG+hOHHeEbsPbhrewVn3gjti
HtpzuMX3BRpW3mkFR1Kz+h9ffyaLwZbOoMsEajr6GGmojmLJXZIBaYz6jJaL
Tlx8Wd3vBTfeDwui4MxTJyPEHAwT1EwcCB4ivvJsKSe8mO6rd3CbzkyLxJYe
xroQmnr0rFpuDEPk/lT2BumFu6Se7+KKe5f0XAHTWWeDLBEmKnUi5PuihW8q
FZk9L9tZfVX61a/miGe1j86ttmD8A5vH3091eE6G6T97QAWMU67NJ/bGHahG
H14iAVbXGs3tQZBtBgFDEO3t2pdCow1IocfTWpZFUJE/XFe2TX7FjaZ+wmqk
LppuUY9F6zwngrIauww3X8jkuJXad8MQSwv+PnCiR+5jUJFExBd9fjUCZWup
vZ7tPW0aUmQVx0VvdvymxmhwITL7Fme1ZPHMxGWfSeb6EXBVcUntRbNIQZN/
/aEhxPFqq8towZ+PQC4qpAjn5Y8mDJ435vzSOgrJcG9YZ+USp7hTbv1965Bu
WIf1MZFuDUJkEeo8bpWP1g1+aMS2VrQvVwroSdnDM/A/90jnjyYSpdadRKhP
gw9IgMtTIhBx7KSYDzhrKEmmJgCAfGIQqXhyyvZwTEs102AlvZHkYHpiPWee
88gv7IIaYRLCDqxZ6/6L05a9lCXbL3+AvHrbDzLpuGve8Ynp73L/mbIx4VPf
v5jamrzpeE8RaLJeQIEPXqqn1eMc6DnpzLRkDDYgioiaqER8wr3VWdG27syU
ab3+j6iKVstjkB+9pHGO2hHfWla5ngvEh/74gG1M+5ZwKWDMrHtGPpWDdz+r
t02AN0a5FlydO9u0+stR0wu7KkYJ4M2Zx/UUbHOiElFZDw09AQ4zoKotMPGu
39ymt2Bm6oN6vLLP0UWIlbUgRCzHKzlPQj+mdNYJTBwyTC70R2twIrJceCPY
wBgFG9hXqN7/dIdQ47Gy77Ro3PQwIFlQgKrhIrCv8Y6WfaEFWnXZ1tcYSlcp
rd9HrCZGPlnHmdREWFI6YkQYL5VB0bmZV1q2h31QxKi1+eVW14gs8e2AUmI4
rPf8FShnfECaMzcpTJlUnVseMhL8r1wuzIqfFm/R6GcDneNQ4kClS3dLVX7q
4nLxU8RJMsJbd+HzLnSAE5MqwaYdeWdTn+xOvrVAmWaj5IMtb8dS2jBERVo+
EbdYD+ZFXvYxVXfg9XMcjRdM/6JKUmzsoMUymA52mDRmgs4ORIFhoZ67Feki
UtVXDsFWtj6KaKL+3S8L4aNaZi6kAauIyNKRdnzGBl0b5jPkkmFp98tB9fv0
kOIs/LUq9jSK8Ruyxjq1oYNyT4Tu4X/aBFGJmZzBCIijQ+JDfSeZs1lL0zv5
YklEfNTDRmqHhXX4iMRbW4hUky0XUeE4i3J9mWJP/Rg/1Qf/HR7skvM7mJ2W
sgEPPY9viW5sFw7RkEaJ8CvQWGobMOLr0uPdhUFLomfwzorYTrw6A3oyAegs
v7T+20wNkLAwN7of2eKHNK5p79/Zl9IIqcENszU8uUwl08hGk2aF2ZOwRKKe
iwyike35kS3hZPLSTJukHdAFDv4wL1/3v/ek3JaYTg2n20JohD9lqxOFFWxI
uZeDr/dDCop/wKW8f9kOXsoPV5h2yrd9DQNl5OCgQbzEEXgi8xRMWpuvRCRP
EyWTP28IqpXFfkfNk6c87K8QOffrU/xKwHh1K9uSXoqBOso+9XwTTiL2H9CI
ZMlNqZI39u5DjJ0J/rarPMv6unVo3jfooH0m3CmSOuePr/1jBCyttDZYIV8u
yNMjb9XdHCrolahXjtHAn1XzMbQhLgNUU97SZ3fHkARPPoEkbDx5tQSpNhkF
TcO137SDrr4Ntep+HtVVAhNKM9pQ26BbYjibBkfmJ06/nKu9EWlPz5VeVwbE
bdl/lQwVrzjdMPeMAOctJVgNE4OEIIkjOj6nMaa9nD/j5Jc20UpLOJlqHiAr
YHPJsw5aGTZ5gcrDS/n+3G2A/An37VySrWdtFJhBbQt/oL4rYY29ZKioooer
DW4QEpACjvOz0RA/lb/4NVbsvmCmXw0WrLBn1boxtYIiCbUV8uQam39EQsnl
y3CDwoDqJBSDhtC29zpVc/7XSXt10FocJwgFe6CWagfOnR2/uomrn/M9uGLo
jOhzjTcp7mC3DoiJlPwqktbKMxygVIAnELtg7/74eU1XwLcaB5fOhUi8i6wh
poBpf8K1HbGT/rkDQiq+34lTotPMwowN080Cx6WiNEgggC+NUJ01NB58w33O
H2MMKj/DYQ2qd4V1ou/3td6JJa/LgkJXONpV2hcRIUIlGOp+x+ccEpKqohFY
fXW4SuorzPVy7QZiY096yaF2zPBenRZxqKacQ2ovPr36WGwyROdt2cu2Gmzz
35xsSET5OsDXGZX0GaIkOO4tmLc5nt98vvOQL6efikrZCVDmzNkLjQ/W6699
O+zcPF5sovu3LIDF0B+n9q40ZHGCxC6EIFyCCzLAh2vJ4SToEhJp1UQsDepE
3rNsXMFVc6GmFt6J43lOB1go2qHn8cRes+q7YUlwJVYdkZbl3XAgbMiSkXWz
cd8xM1EGCvSsj+dZnFzCMK0QadL/jEcx/LbFlbMIohFCxplhDRiGxa0zDvlo
j8SfLULZ1Jigfhys98JBA2Rmp1zpxNvw4s6mmIjpeKP54+3vkN6NIV9uDXtq
L8vgjkvLiB8UT/CSikQBEVj/GmDO+Did7BdCyZiZ5LbOCQ1zo4uZ3n+9qrbE
oFxqHkg2vIXB1pciVK27RI+Bp8iO3JzKFPGwaqjO983pFElc75hdrOrCQM4h
ABdB4fHgxWr2YnVNzRRykJCaRZQpZA4kCgy6fzgDA3zAtEDldRRDc3ifo+cb
HggG+AFCQ/KK8AwjRiDvxrTG4qg09uRN1dFQH+bIfqLm2sjBTMW9YwpOq3z4
WRyEwKjtnu4JyAbeU7XTNmXDqfeNZDI1MeIJsocQCVn2wa/KVAUkliwn6wds
ea1bunlqKLy51gXa5gi5ISQVbJHQH/7jh+9ix3PFK3NmZdwcE2n7AUTKO3WX
LF/zq4sWg7Y3pwuznYRxyiEsJriwPid0ZpkO5vSaadE6aZaZqv3j0359tRC4
vtKOgTnYHvvWtodt4jQh0lPCLD0IRfa0v94tFmFmfLuBINvib3cM2XSSKyLC
Dqi7hPMndVZTtauH/A3g8JU4WZimV6VB3mAABMEeW7qdu6DIZO0TeOiF6hom
nHo7HwIpMtQyWy2utSluN01JYCHMaAseLyTuqZg2HwyR8x1JYQrwnZllsZGn
aHipNEN/gr4llKU3QGtlfLbyOSv45iEY3SX+wEfhvpcKZnPNtLvH3vSUPjnm
B+4YA2r9qUqmU/WvsNvvczdR8Mf4Jv3OVeQEDOmzbw/Q9gKjF4ANo716Ftfu
KTx7d7gGoZpCslVsq9Uzh9stY0NowAw0bWnO1ONI3/kR0FKZ2ZvK/YIPUqBn
CAlaydLC3uBVhf+IJgB+QDOgY0TBTufJgwLVE4t9GqNqthQJrHAWJML5WPbA
//V7KxWAI/Bg2VDgq6EhMHtM4KAA/g4hWA/WPaBa7py1FkHakmpXEUZLmSbw
Iu35wbZGJrA6cb3wB6O+jlnkY7G/KoxwJZn5/OjWe3vneQTstRVzy+zUDVoc
/YhusAbKpaTspusGpCBcLQOeEsCCdODhmGZ4TpF8s04992ZNlE3WveIkoh7V
DZ5BRXhaiTTY0oUJorlgWfH23sBYN6scQJWjYYiz/5g2xfAQpqE+j2Ftl2Oq
4JetxQm/ebRaMmGjRgugfy5NtzFaoFIaSqqK1LGWfNeZYwffALhLTDxDvaEy
nuVxMcJlqe2CIKZf68bEd9p3b9e1/X8jq9UwT4hbr8NgpsRNeY9eauv0IudZ
d2T5iyc99H/kPAXzWX3eqGxSW6zTUvTXlkKtqyJALZ/zZoZvgmMcqqugh3dO
yVS9Dr3rXM3Bk8mz7sUEPertIj5NcC9q/2SQzjUpd30hBkGUum7PLzSO3hOX
Q2xSLIuhY67Ttg2Idrl/5tNeBX3Aykqq1chPz1fF2q1MY4SDSApVY7rYLZHp
KqPsKA2nickKsSzicELhZYqQbTFostC29V4MQ+21nMgIVYblOFSYQ2QLGP7z
eOprfNW3oC1gv6IqoSdRuUebTpWXw8EfijXf8nD2TIfbHl6rRq6YjdM9I/Dc
SVbIbPUC4x+gHty+ymNzKuHSGDniACQ7+k1eO/C7YcreeM472cgWROHr3SW9
PKCgYohgtxpm7ezFq4+LYMt0eo1Doq/kF0wqk/L2kbuvT19AJB6YLdPKjCWD
dcfDa/vR+UnPshDRX+OEuluH6ZF9iyqT7Or6UtpxV1/gGeedLQsXJC3ul2ul
HSeOfAaZRwqjk/cfC0hMQjpWcDKabwvSQAT2UPcxyvhhrj0FJUhKcd9e0TWT
JQxgxrH921fnGm1RnzzY6yNq9IX1jYq8khjhuZwdPzohhUQ1zhEB5Fo2+Vyi
n9N45ngpNboHdRyl8nlioFYmoF4yEFTGlwp57ha8ucSqoYNybHVW4Fsv2t5X
LcW47MfY5Jt1qfMME+Up3tX5HEEwoyw+t1fnK7b0rF/0R60MXrdhYv1fGfEs
4M8DRKEb/1HM7DD0O7dNmxKz3sCx8Y5sXcS8F5x4PQSmToUaN/7Ujwqcvdjj
4Pc3V8lb0MXsTBckLWECp57mp6kkGn8vfX1K18EZ4/NhF0yAyvWVmu4FzJVw
CPBr1eRsVZv9LSBlgTXlbsqASG8sRFiPPBjIQXCzH5NCiSSPxmzJHimVObu7
QeaulzNVczU7O9/32RhadH8k/6MYl1wCAD9TT1mZJZMz14oQ9zxPdj417ij3
PqU3TThZLLJrvdrcqFFYy8aVtYFqkxHLPBQtmJ0FID1B6LzdblpFYesAU1vW
5K42+iZiSCj7um8BvAwKMRyZJQ/AH3MI/FdVPxJDvftWkYlAVAnmVVQkT52M
y4hDg9SPoil0Z0Ss7ThM+ffdsR93LvVpLzT0e0HJZE5dN3Q3KsdqT4sXJlIT
cgMy+H2pKvr412uW7KD315oKxCcTNlotT5/dF0+Yzovm8va0EkjgBqRwTvRF
8IyV6zQXy9u/0/eRkKFtb/soXRAbxlqnkK+iQmHnw38Mru8koO/99XMC92o/
/SMlACGxLVdPYHBtIpQ51rqYdoI9qWOR3dD/PoNVDrIlVTPpfB6RpCM5qcRd
k2hz6CsRS7QOx0HqJIVmqnCd9yLGNuYm/JO+1ggkZN162AuhNCH+TZHECZko
9PuK9qGlAgJgCAiDBr+PJ4DsPJknGoaTv69X3oDq3nkucMoNKc51vCw1GNqC
V0zDe7VX7+YjCCYiqOkLf3dSBTTh43acSNpuWHjqjTG0Me0ZtjZqPMpVbwB4
c8dcGDi5at3Y0jhKqeX3r7CPmrBiYdHEvufOMlGc/nlk7YP8zqcZTdax83ZC
U2G9a5+k26/X/VlD5HNsyPaxqrtin3+A81ajzFjc/BiyxENf+bysNmeXJFsg
H5skCVGBXl/iInS5vv+huXhmcW74A/m3DW+n6iavA7guFxqQU9jVu5oZqjBS
m2IlqLZ5bIXd80icZ3kK8v5gAmKM8dl/qWWEJ87xY616rjdCJQ/DzuylKtqd
ZLJCw492qHF+OQY77dbmtEMvhCbuBjstCnsxs8dmIgkqx2TYFSvnubj/CeDY
hLWeOzttc5LLvfWdfdfqLqAhb0uhq8nWjUhWp16WLq0B6w2xYFGHRaNjj/iq
QKMhVkluqU2S/ws9FNK6lYEuowWkOZZKCWsj+kxmkgKHM+7jHlAXWzZqcocU
UYckMXd7goTnxWwbxbj/X/p4Vp7obhjYgQ7YY7GWIFfoONrWmeS6eIDDBUtZ
7T6ZFoD1rjZ+s5dP1k+8r+HCf4FEIe48q8T5qred3aayVKh3dPBfZ/SSY6mr
ulRbStVFCRhwgSl/YhuP++t7XTPyHFdP4q4IMRP/6HqjaI7EezQnBaX74ee8
Q/8FmKGdmWgn5Iuifk5qxbXJmJwKBdOXRvUCJL/1dGrsbkrytYL9Ordv5QP6
4/UivOnGvGcDocVdg9i56IFFGDmoiNHmKRSB5KjOj+yFILqtePQ2UXs0vV8b
8uACzUxlANrgFcvQopx9ccExzbJOuAATv7QupEjlktcSRSpk06hSiCLPYKtU
hs0LY+uw99Io6RqEQnPmoVUU3KA4uLJcX06pQi6KL4EB2XTJC8/Uf69PIBmb
soB5AL+5oeF03sCxjMaao1KCM68beXCeRXTLNHwUgg7DYsqCPHKMOlBJBZvm
aRuTdt/zejzbO60sa3kkHvNx4yBg/G0cO5s1bP6LNGv2/otSKFsjPY+cWauX
eqoM5gE/SEX1g3VkB2CMk8053Ulg/m5wz8tV/5Ty/VrydDKETsV6TNV0nIwk
5QCRCIXtmyDWliTlhEI+d6a+wvK2lMtl/JzaekxXBUBQyt4j7rSyTdaD4jdi
t9DJYO0ElrPqTX4T/P7bgOePyyc8SHi3HBK5/uWmaD7z4NaNkDeed6GXeE+0
xQdUOBYA2pd/jv0BEoOU2YOgK9hHOXmqtYQYwKadVFSKGx093fiWI6/h6P7l
gAeJ8u32gBMM47WYFXKhfoC9xWkaGbvd3NpDAGkQCibI/hlKYbUP9jPQuf8P
ecmdhF02cbMFXWl0QcOOWXU6FYMhdSlZuWygEAeDDwY+Ixs/EKnbXqy6oXDh
/xnWGr3P6Do30+X2+wi7nTF/Ql8uvxfPDzfki7fYu+MaXqGjMJzUsJoVo75r
s/ANs5teo790/+js4DJwTbiUxV1UB95xG/Ua4Wl0rJARjf7a5pn/HbGFj11+
z1628Z3Kj7VJiiHkIW3gLTiPP0lw+hguKB+CxAv8D9h/aJKDAyXqx1wG9rpS
5WjzlaYuPBGt94AGacSXLPeNoLr1Gki2yuFFjFWNPPWQYzM87EfeZNB6NMiz
osSyBLaAjsCXhzUd7A/Rcmo+D0qz9cmXv5WnhUVN0R3NpL4smY17Wrt3YN+R
grzRuOUQXpLlnASIHfPPYO9XgtzzqsI5hGDe9LDKDdeH+hmmo8V+uLlwiQmw
WGRps4RwQewo//BlshE8XgZmHpZNfn9m8MaqnVDCwl19k+/2IGG/b+X89vck
UJaK5wk8olacesVrrVJc7+ZzNCoFFbn7mg8tMMkMnAv+2nYb2T1rQJ4D7I3p
K5/G1gCJ+4A5NZOxxyqdNiSOV9EwlEcfOMBioLwPO+ee95Ur0aj7r0hCFhek
5eo8xz6xXWwryqaUcXdUf41tPRdAl6AYuiNaCQoWqoIJWILNNLpSabbOjeyV
OTRSnAIyUWHaj081Dhpg8OXvzy6myigkX6R2aS7PxeQCUzjpFjXrhRcmyPNi
4ycljzm++ajtPpExkdvi/yILD6CsUv6juuMRQNVe6PAJsrloVqAqbqZ7nh2+
oNddAAalcbWeZjNn663kEWzQXDpAbP8/S//zOdUyRz+x0wPHT2kdP5WrRZdO
rmppTopFMgJp9bORxYwazINOIrCYwLPQt6MGJu71mvDI7KuRYSyYwU32iuPk
Qx7TPSFCeIWpU54YUpQkVZldeaII5dfBUALme7wKIG9fYfkbb+EZVng26NkA
Ksrm9ySW/XvyjZwKYmPerdRstUc8NGoFANsj7cEhZuaxx5JMQ0Z5bbgbQldf
TUfNcRztWhfTLxPqrK9nppBONogIKv6H7t3V/RkCtdSjQKWP+nrf2eS3IytB
EYsNFX+dUujMOp8UGwQh+FylMPWr/LUmzzTo2+EsuQkx89LgnWFd2WNENU0/
RM8j3pKGcaGZp06ocIV3i6zprqMKZlNu3LE2eR+7h81ip9ZZ9TIJlCp6GsnV
Bg6q4prvKtlp4j5AofMIRvdIPgs7fYGUYmm10xNY2jQpnHLzvbvE0l9fA+MH
ONOjr1EtkworC3Ap1UPEjZDbqqf60Grjq2vGXNsy075AlV1gB/rgMxhHCzN/
zOGC56tG1WuZGNvdmwxvGHCNLnspURELN/PBo1zccFZmSLwy20JQIi3vkMAU
v2WOsuxsqgLIckMYjbv6q6y/hlQ4r4UJGDmJCKl6dMhmgnysvafWAm7QaxHF
DV0epF8Jb5fyTaMX8vVq0+AVs6ypnlGyZlLJ8/h5a/6YOUXj2IVDwNOA5PDc
nFbR4NyT7TfpkPvOPNyb/TJwKtVP0PJDC8xZuEqqQq0YwCpgWOJg7C3SHBt0
LKSZQ5Lr95F4olcb3ZF9IwwLIHGZC+YjPcj/UO5OfhBjnjObq4sWIkrdeggi
J33GiUm/Vqg2ObAJ87z6WFrC4I+u4OaCchIqlDLyrHyP9I1ecZS3Y2Op89Xb
ylmyM4UE3CjnrXeyd/za53Y6UVeuRFNwK+Hd3TgrlkF0n3JXg6RJSu89tZkN
FvAIE2KtP6JtjpLqcWHSf7hBCKq5sZ5xeGgf61l6bK+ju3UC/s0P4ZDHKMCZ
OPfUXqZWwS5HhhumB/HeA2MyKoe4iSD6YR0l6Xy4erQ63GqhCZITyDxg8BrT
fyxEgRrNYY/3/6Pw3t0iklPz5Ic1ss5BOSQdS8ydonlGZxkTBHoheO4hvqh6
FsBdQ8Sw6waRl8Th7SIlBzfsWpz7xR4jtlbXjH1PKbBFWL/yNZngEkD4fo9h
Bebtv1+JfD8I5DZwoU3CIVHbKkD1dmCSAZaZ6r5GBkfR19iYQbMq5iC7en9E
449WSMEn4k83RQH5t2ssAvYC4GLx7YJfh4UekMnaA8NzABebWkP2sdukbyvI
eTFX1FiFZco5w0L52Uh81ciO4SV4Qr/bjr0h/mnJ275gQ+1fwgxCzO24bCgk
2/An2EYH2FR7ZDz138NvXHbdtEg8S63zrGHv00TRR/Au1dBmcq74T1tFlYX3
xZ/O9XLZAsq41wQ6fGBAGav0L2xwSiIUZ8b3sEOg9HdH+9BS8K/yYtyvYdL5
9lBSoPMumnTgIfWHvRPPJVHpxjx9mI/TK+CM7wX3PNker7gf6cEeZo8rRLEE
eZud08Ju8wGm3/ghAIayWIOpgCGZsUasD/sTD1gzhj408YCa5mOPRcMbmflj
9v55xYX/dLGLZcpNoeBiekjjY48S+RACIqyzLFY7JBL3MmYdSVkFz/xsSGUf
U5fN/fd1ydSsPELkNVJk+my1+x/tE4GwEMZyAkruKVm4lxcWAtssmEHrnsiJ
6IE0Yia4Na3ILFa5qdX5b4gX1HYhQS1jntRjMih/LWC1TDFQchi1gl6kZJRt
OQaiY41AZPF9Sl0/aKOj62Es7J8IgWCgKcOjFYCaGaFBOTGDma+iC8E4pVeg
5R0j1e3n+5kro98umlMsxKaVmKg5NoCUeuM1PdLmF/wkSP2pz1qdkW8/+zxS
1G3LCF4JzZihElZr67ovJ+U9zY1S3bsts0mjGQrnBHpT4voiSrUSTuCjU72W
YjwuM/Ad68+NuLPcjGQ+a82nnYgy0Xi3TwVX2Z7GwZ0m9xumgoi2XSxoDfC5
1IYngSY6HZd1a1T7Wg9U6URsiuaVaicMQCcQgohekXaTeHpYCOvnOkLKdVWA
1gXY7hmaeXsY2UJHlVnwzm7ddYtPslrh6OnoPMDl1W2STlQ5dYWOSlKrgFYW
0KdkoXEg0C4mfAg4Ne5Y6xYip8zezcZE+Dw4q14KjfJUM+4Uv6Xn93u0veQl
gynvwichSWFdnN+C06KcER7HdjeTf5PtwHjHN68dR2VKtWytYfmzbZ61JsU5
8FprY8SUI6kS1COZ2k5llHL87DWYLe1bXULadFOf9F7NvnGnKmOf4BC7tF4p
VHML9Tf1Rxc3pRiLvTcEReOKu5sETSM29I1VcpXmGWvsRmJvA189EJIo6G/d
+rMyOpmlfIFA3OrvIAQPlUuKWDCM46Tb9sRqyuw3Sd5rvoR3MduLP6fbwtp/
CI9A2g5714YV+t18bzVGZ/mm4s8lZtu8ptcHiyA8RLRwPJyY0JEc5XEi4YgZ
238agK9pUndtfO5+dsxDWArs5cGmIEjuOlU7VHlPOJqTMXIZiM3jCMkz2FOM
kMcxrB7qhAAHQLYxe8P/vhrjofMj307DfGlPeixH9tWw0joSoMKzvzgG8GF4
94EtrIiAU1W5EW+myLldZj4MdiGJ5dGy+N+VEKakggL46h7sSIMMATzKbxGm
0AjeMwiJrJoS3QkRolcCaZOoNeUoHJGUcyobO1gidDx4F/eFFtAV+a6q9Wxn
SivXWc4RUJCYU9TV67vGMjY70kYsTe3XZvS+vMyLF7jGlDNrRhK+zRiuc1K+
OXyVCj79o+koQqRxdrqj/92fkJJteU2vyN592AqyJKZZqnYTZa2CWORRdWIE
Le+deLACz2l87PShcQBwRNRbdjYfAmRNIiQFI/ijfPTKYj3Nxna1JolwMQRa
ogVusLviGD4K6rAnQfUz8BOqzfcqoQVyqYsQfAnI0Z3sw+XjKW/ZrIrv3oTS
079ax4HeXYPNXRBfi16mvlAdVDGPBJUXrhQQ5kQvxf0MQvxrjy32Bmx5Aya7
28UenmHPap0LrmYKbLFSXq51alvpuKsyJ44mIGekhtsrTqcPCOMtjFh6PHG1
Nu3qddzNRi7QTSsPavuZGCsbGyAMOqXiS+FVPPDL5oL4P+TZUmTKGXUKiNcD
d7NzfeGxIn8zmKEw5sqPj6QfBx2ZYHNbl81ghJz/tSQlCjx3yKKwVPsufcpG
f+eBMEhgIYUtegiXD0dOa1yQ9nd34TZkhMiSQ78WCeoZwZERUtaOwBrwEOnt
eMwmCeOfD+W4aaPyncsdEuRAnHikHAq5BOl60usdtFI9SLwBUnc2qvuQ6UON
sC5NY5heLbMI2Sl5f8qNg12V5o+P49fESAkU0/8YuWelbPg0CV/nd6y+4lIk
3aeuPsAKjY2oyrJXEMy3BAjGWCwDwFR62imxw/QqSlyeTF2HvuR7mUQZ5W6i
VdN4dz8gjrRkS9zY9vGJgxpN5Yobeqipno6FwTPY1ZE2JOKqN8jql3GOxlUz
/a1ywCFHHTMMaL0pxClcEmoNZuiRWm9ylRNFYUmo2eIPG2a32tSw5U6YbcQ3
em4rfcbkR8Tpifm8jh5Hb0mN6B8raWVpiBuM85uGqQlOlyg85DZ0eANd8Zmt
wjhSWsSBYVdzwbQDsv2lr7A82C8EJtWbH5gvVq98i8A2nsuXCe6cz4btWM/o
OoJSDkHGlDLDeGRcazwDHGE0teq0YooGmBCMtucOw6VAnR0IxH2I0JqfQkpc
obO170VzfjdKV3sP/dNJYZdg7L6a9g9Xmsp3UDRvXUnr5ztQAdK/yERa1hqO
9VeG8fgMX52cTfSfO0i2IjQE6xu3uYl+KZvxtPKLQmjRBP1vGHvleo0Y690k
aIM4TSg05gHkDIrVgihBAIjLmi3lPxbsLOnxmbGwyml8pVP5yOOE5Yqjo23A
JYyvnL5m3u1+Prd5kUMb7evlUOlXK3Xj963Ig/LB/WYEynrYD40dxz/lpd4U
5+DxuyxsUW/E0wmH0PiA79sZQ3UP1GMB49mIc0bpAtd7tUD9JJwI0nAHd+KJ
gBy/fvYI3Xbt7HJm19x5epllBiFTSrhneVVMVe4AHxbMaaRjHYEysWbSvOrN
/MBPc1/HPouiOwjLGWU/+RhOh212FgLyscfJHQgZL2t4Z7pm2VkNV3/FGqJT
wa8hO2icGlqHHTNHcvX50lYBjcyzkgzspxebpb5ZRoCgkmtvhsaugmoJVcFS
GUujsOB1MGa61JVTnl1gMB2BaUg7M/SxDQ1cbk6PvLN674wxgM9FM7F4fF6T
b/ZPVVPuUyR9dwdwm1igtUUdnFp/E2pyD+mEiaT3qk6Rri9jRYOkjC2z6d7h
j1AsshgJskuU+PpXvAkxTelcfWIV19pNWZt7eTcdJtg9+F0D0PPGMA2tznEo
eMADePUCBsxsYxyBB9fhUwaKnJ9nDJs+uV98y1GJCiP8CHqtJNoNVqx8O+jH
CSzHoltXYjydoLazgDt8si6J5jV2An85tuzaPi8pKK1gSBIsO3mF1LfovKja
qmd+stR3+lmZD9HF91hq7rboIHvOftNWY+zqw7jWjX6RciBfO3yRhV38ApXd
AwPOBe5D5kGInf3apH3aVCuPTZdwx27x9wKQ75uwLBiq1iBRu/G0F9cUuixt
xSbFhkMsE6G04mOZHHQBcsLmN+eEZZJgyS2i90Em1IbwUuL6iAsHH2b11yfl
IHaTRAfkVIfjEkOzw5oR5nrxyUH572HMjV6Bw2XPujbyZbFlqz2APCWUtiHE
vrxqxAZcJREHfnBUQwTCZBouVJ9JvagGcRKZ5gHBo2s6/ZSz6igE3ceR5AnW
7QvSbQPrm6+DFGpoP02Ky3DWy7o1/zFFZ4DtHjlODSy554ghY68OrY6/UknU
U/iRmhC7pgloHB9DbMeHStFki4dnjrFw/o0F1eYB/YDieFJRNoSHpUqjiSXy
b21CsU5LBM0HKKtD17pjE22HyNH6UHD0/J+BaaqgTCx5BEP1FB4oHPQalOAe
gyjg98nA5zJ3YOPPBRNps6pP9P3S32WKj73d92EEj9wFFvKNX2BSegLjf/D1
4K9fbR6FbHpkNRV1RXh5i3pzzT+2gCSBGP/MiJ4Jr0ixmSBpOcWzRDNX+fu2
3BT0N7WNFUbiukIsTnU66B2ZPGfFmI6kWe7iamkTwpdecQpLyuxINaWklnFe
h950jId56qtimMDoe8aahWty/VLBETkCiDSiJgwhOrvXPrfoB5tsya3cumYE
c+s2v4bNcBccHdqgDgO7vxHuhY2R1t3c0oGWWNqDNR+KmeUtHUSP5vOcuXK0
O3MdJrEzdMCzIRNyGTyESuLBnfB4Zkf+ayt54D6gSAufb62ahzLBIx2FfYXM
ReaPResymxc/OK4KNnj4nS0/Qt6MqCvKVjsyq/fwUBiTHUWw9oH/qRGiWUsS
XQYB8c2G4/fg5fvYAjkXpYQt0vYiiuZLdsa8MFZKyHe6OdxIKEedhlU4F/vx
dpNH4hxyvvJHha66xfVQ20e7eiHq/OAkRYMDWHVV1jtu4B1+s0qK4zAnOCOy
A+nKAYF0Eh14q4AzE71qZ/JK+JgcZIB8kjfB0tCz8BdZNs3OueW0JHzk9xvI
CpHeK6l45T+hEUfFTP+eNRXzAqgyQ76+Krq5KaE86HBL0+M/nAKN11x99AO5
rzl23NAo1u+UBu2EHhDB7QClFI81iNMLec2lhscFvv+ApQ43XUGIB2q6vmaj
k+NY8gaDoGnnO/JPxdgPw02Vox9yWZdBg0KQmKAuG9y0cy6+DhI+XUO2/Rmu
/+d7ZC8cdO0ENVCgPkoI8L+kJQa1MrhHfa7KyWM4vc/f8U0iHxMkHwHnuZN3
jDCQGZQ91tsE3GQPegySXFsiRY0e0zLhZMp+ynC1cViibbc1JTGh2Jqi1T/Q
ftA2m7FlvJWx9GyUMH31HEmj4sWlgAGM3twb50mEeKj/1vK8QMudPWz4MkKP
CQEH/uaG8evpACkRiGZ07eT7FLWK6ZpSg8e8jsgyduJv2rV7qQUStxFasWIj
cQDeINEWN0bCRAUZeMA25HyFyhyXc4lVY9n89GDinkSWNXPtzG5HXIzspAK/
qKAZfuNNmC39VXfu/ZBofn7ha4z30kDQMxK8jMrEW0dVuI3ySvVA5z8MMqPu
XvIhIPwan2e3bfVFoQMvEgK4mnKOyCF5lsk1n/BZChhlLO2xBYuK+aSYRTmJ
xdu68czd8aG2j4r+dGbz/sY7AovBtwLitMiFUaYbOBPQH8JIRi3R0tWnr41T
OujWKnLfHoQtkt9wqzsxfXKbl/XldRaiBDNFKa+UaLVXWWV+4M3O5C3ua6rF
x2qlvdhlzWB3KsgUW1h8z+BPAfCj/zZNs0aZ3FGonRWjowNog9/FXqCr46Gu
9Bs76+7tRtvtX/N0KxZK2AcolrzocSLhkD5wM4B+aglVSBSKR0rCv8o7cXlV
mHNjtLPwuP6z/tXcUWB4WwKI1NWxQ1X05NTiijfdLarEPo4FbvieEx52kfAn
jfDOIbFDWwIexYBb15vj4ryULM9j6aghBNozyKzwtjhxEclc6bXLgr4CxlUO
/4o6BF+PPYOAcLCJxC0JPdPlKSe/i2V403POfdYuNbwio3q1UzQpRF6RjoPr
DMC4JeutIffrHD7MBj3CugtqdIMbInC/UqOrC+4L0qVA3MuRhN7gGHg1W8u1
Nm6VXqLC+Z8gpl73F/uP+XsPJdYDNz75nuPOduxaM1u7vlD4w+gNhOM414sT
dFCaiu5IJs+ccHTF7/1xf6qiSMTswC8sCbuzId4oZDaE0GazPXCCscTo4W8+
A2maTXtM8w0MtC9kBRuDnyffFYcYEY8JJrusPZ71oPzX02orH2e/4+6gVEzU
HzYkrr5/WHdKvy53gSPzy3yjtknqc4F/NEPo8mLZWxaXxmfE+lJKiG2gsPB3
HX4GplwtW14QwvzwR8WM4sxFdNl8xxrNdHgW5Ur6pCCYn2tVGIx34fnWvp5o
zjw70ogrP7SASWVKuII1VuaCv38HxvQJlTkF597PoDblRvia+t0RmhkLhRZH
FTpLNLnwJbAuAYzLARmWvD8UccqM0RIlg8M0PesrBAre5F+ZdX6FDG3VdDzs
pksZCDeWDJS5yFtAEKv8D7TX8N1aFHBq4yEWHYTvQz9h+DdmAXp4kluzJe4K
q5FiqwROrJq9Jpvclty2denGrtLGNpQk3UAniO/myidpVyN047w+ys6eZmav
BFHAviiTNjXrEVSpMska7sahGJy1nthQw3dd6J2iqO8dWe5pFqCD/FzoDtOg
ym2+F51UUhFukeTCSjkUZaJC4uwHb2MSqjnPztCzbTNJh9qY9KBHzF710wKZ
cYXz4yErffT/+pOM6u389/iKgrl3CCytWThvXGu5QLpGHne7UPRW4DMYmBxR
ddQvZMFnJ40SMhPTotXVfVDmrN7e31vPhVsvoe1gROtMU7MeTP/xWkQcvs+q
cHargQMx6Ajeq5qZi8iyhwiHfZTU9xrNK8KsOss3DF/ydLgLaGv+2zsxNHz8
hF2NcR9Kd4lnOYcKEDq2fROVobnTweejSLorujZnpvpHyP4UWj39sgYzOy5G
3EwPeuJ1jZZ0ilwe71bL4/JQznQ8bRBQjRp+bTl50EUyRh/4Tr1FDKm6OvYO
bipMJL7ed/Z3xo347Rh3KdklCOfttUuQ0DPtOfEbR/4DbE0bK1XDaOWUzOrO
hlqSgb4myglKzUuVQ0v1lLWNjFHTG0oTEyV1FrFnUMapzWwLPwFsLsmXnica
mTGCnVxn+WN6JS6lDWZucj7LNUBdskJFweeYCQkyFZoTvQqTV8mOzakEC5lc
quWakcmVuGFvdfGqJZqyALd9Rxu7XRr7eN5OIlYFmbfaZOeh1+vKcozFoD5E
9/hHiSv2bRDiu4JQnglJc48gcHOK02jMRJJ6/i1b8FHfnm0h0rluNL+qFaZO
M0SZvwT6Zpb82Gwxzro8BD94nNlwKlZVWTv+uQvMn9JnwhT3AN1+ELm4vdxM
aU+3rU9eyr7gDOnu9fd6i04vMt2F0sAzaHMS/4ymKQ0NyQNI4jiQ8QQB3jQ/
pW08SyIByFw0YLKTQxdnX9lcVLfSUVKKRF9yjnMuUrlJ7ZKCrCvho5ymzx87
l+5mdgrOJDuklidlPCy+rvf9mVotLDZryueqNdjFLhWSz7VL384Bckzm0iot
GfxV4T4nH7qGoXhnlLvGxjYWs8pw4u5Lgs8XSimIounjvTXPlN0Ww9MlpUvP
MQSV7yRPE72gbC7kpehtMAAemSLnN63KakX5KMdDHRKe9tsqOZBdmyiI9AAb
s9zTAKnogDmKsJ9Mp1GT7zAnMZI5A9ZuqkkXQU+fLoICqyjZ1iXqFOhHvF42
boScjOYXh4E2DuYWqAq4iualy0Y9Fn9lfM+fixia87e3cd93opVeivZ+vs8/
Y2f3TIGXwL3HhFnSkEv8WqhS/spIeNZgYAEjdu6HVMgHVJyeBzOeX9+d5aKb
EtTqyBeIhCOGkma8rQWYu9LdAKD8Z8VAf81ShiMFE2BCcMfIQ5e5UBHqkmLh
3jqn3UnYj/nGgAW4dWRUS5gs5KvfK3/+Csz55A63LgnHpNYvNVZGGsh4cOwv
pMgYGFIzxXAnfiGv+fXTjmBJVufXku7jGddAyyczC9raZqRP2O1vOJ37Xkh2
6HjyAfu9ij2uJdrQUeKYgUepc5kwEivRwzB3Nc69j9vbJoJUsgvXsdwLqiWz
R5loT8PmzPXZM3XNXaqlKUN+ZgJKqEuVOLIFAxDcBdq43sEUMAk2/0ZD1n09
nswjxUGFuxNyxKx73D9LVqakLUOS14mMzofErXgP5+HxlIr9UAKxCzoSYwgj
ENsvI8vzkSj6CHxvdoArSVz196avR9/NAYsAKF+qPYFC4TEKqSxM0RWI1Yoj
agMBHvlAnXHHFC6wcPwytZzc7jA8HIbDmzMeTWdfFgL2TOl05D+uA5ks+jhR
YqE76eg1dq2+w76f4E0Q0Jfx1MoOrZeJZKI/+NsP6nJMd/9srXAIy37ueHOF
T9HZIJXRQdrvSZGjphjnWuREBuVTHayyRaEBySRvY57CPQh47kdNkI86tWUu
F+RH7+2LR6rywWe41Tf6BV7n+wn7GzBnp5YRLjmilpBizuq2VdfBUAVVZSQZ
b42sgmmv25zI8teq0pBsG9b9ASDc6L3vp0dvr84eGfaygTSqYgzfv2vZWExq
rkYhOoo2370+r46GXCAIf3V02xXDYTlLD7V2FuXk1jJDBEsSxAJnveLsbiMV
fp75SovnxnrD5tWn2z/D36fOjWvpd7e/Tu3SxZxyNKIKpcT/74T+RlIuC0Ah
afkfNc31ILj8eEpGpeirUyYTcmXr4pwCKu5BSNWlN5HhumIghO63pp5U+6fn
DhJQdsDHjhKbI1aZp0nD2CcHvncNBv/Pjspn6XOMZ+OuNP17MWs6Xqr/uSXI
qtg9mYl4goNex+89Pub/zRlx0YXRW058UmcamFtNWHa9H70P7Jn9/4YfsFTt
G1CtXuzeZDk18gUBO3bebBwO8owYLygsYZDyLv6krejWxBiI5zg3VcVejyYN
DufgUj5MdOO2h0xK1CqN3iCk4qvP6kWAZBvwGAyTqe3ST7/rtViU3ixuzayV
jGeUIgFx6VwxVn/+TjdHWdFSB4OJoq6Hvm1GnFAeX6i89j1nqJGNnUIpyV/7
yH3K+muCOFaxMeHqnNDRv3oKjYcls8ziDHDhd43aalK8DwXb31BHhN2s8tQs
tnYAyj5RPmYS7X+xHTIcb/3JtOjuE8l573IWNEubAfuXOe4ervAL9op8Z8uZ
K0QbsBUmjho5XUadCnMRa/ADMv8EbYCnuP6lgxz3WgbjZGfnMs5IkwHTHPQl
goXspazpMLUqi3g1q7mNHaq7PfzQeP1gg3ps50Rz4uEF2Lg7cWZDe0TA1eB5
m6WoLpbpCOXJCu4w7nl3TTco9phMh14GX6+xTGj8jZilDr/EULIHgNmPgCmF
Dk/AJufPxjk3WoZVq80AReGc4SADEKTIBpea0lomhzL+eokjkfi5FbK1jZh0
gxD5ATv3o8lJ+VFvYJM5eFNvwprn/cx5JXCCvZmBKgbWHXiB/IRGDt8MpnTD
kW0KsLv+tSxztpDNJmCe/y6jFxV4Jey44FdU2g6mwO6BXTClQ/JBafK/f3xy
fcV2wqbDwQgKMbO91gbYNkQIuu5BBlPu/xrmfxfs2wu3vhv1EGoWCkuc0sbJ
xnT51Sxdf6VJlj4MXv8yVK8OF6HcbYoCLifWUy2A6sO5L3fSMGDu3TnHL+Jh
3MuKdMh4ZjOxtJ4G70T5HM7/OQa3X3pmc9KPlTAQZ6EhWrcLMOPDxZUIKKTV
aQqP4yTrcZxwG6mFvw9Xc7k6vlWZYoB8KEcKpOTd5pqpKFN3KZJbF8n3HAQw
KDzHWTuPMK5NoOcL3C+RAnOqQas19voBbAFcCQJu1pQJSW4xdOJj9jfhODBt
dUTM/s8exsGWyAC3V5h/SQIzKVeOjWg1aggiBn/OgjiKJOvHivhztB5lgvr6
lIXs30Rubp/mmr6/sEw1FsNGgGegBfuFyIGZdhQnqRVPWuF2+mYS9PT8WlnH
xxTefm+XkSV3esL0WV+gVjyVSFYnk5QReBrrTN2S/dlJiTX8n7/wGPaUn5AW
BbzR29FmD6ZWQt/+2/RQd3dVy9IMwIn7eZLhvIpVgvgKv0/5D6oqp4y1PnIi
6E24QC3inxkrygAgbb7eCYT9kSXKVlRJjMfoP8/wCXiyXUXNeT3bEpiKttbP
Ya5RMytTBR1xw/ZlFALgJ5Gr/dwyUhBbub439xOZ6seY9S226EW1JVlQh2lJ
btzWH2Etq6Qfx70T6ibQcgTHK2UNnAqkGG4Y4L3Ff8v8UCTyOHjbnbhNWm63
T6CyVhOpuuAD43sviVxVQTgd86kxMqrU9/OySsmjQ7aB2V1ihCqQLyYCDQHC
BoxYLG0MlgyC72CSEA0FD+4lcnZ5HQ3miB5C/aEzLrxaJBt3qEoWp/lVMhYO
hmL9GCRTMsT5jImJXEL/qr73lKc15kmsh6qqlmqKzU3/c2RabsWJTPR2HROM
i5G9+0gjCTuNHounzqSTwfHfzZW63sjgda27FO8UPPYCQbYrPZO/vDAwOtHG
aWh9ExmGUSzLEP4/HiQYJPUSYuJcHK9muslxRcL1EnQZ2OpAApBbS0URegnZ
PpaHPqn2r6I4Wc7DKRZXE/14Iwr4fJeIWhgQkz3XJxgNSmHfYEcqXYb6adLX
bHE2Yyl3XxV5eUqhiLPlkIkgtId6TTpEIKSBjmTWMPIFECAC5z8bYq2QgViS
r5/ANPnDBshI7tvBOrU9y5PZfs1iwee8dR72dtxJFx9+lzd80cKn8cuDphyI
KioqglCZxC3CERyTPiAVbIIDVTrH7ZMoxelhbFIIyrGORkDO87gNfV3ffPou
Fflz+0u3SUgE4VG4LJsfDSUqDngrG0AYQnMHsRuE7kKl6XXAm+5DEzkGcdFq
jnP9NtGc+6hr6YRfAyo3+lXBWRMZ6auNEFEVitfQ6JMARR6N/2jy9bKnOVa1
QX4JhMJnmktZJYoqg040qYLvTcNCCa1HCkxW3SCPz8sh2sa8euPvqGhWWM5Y
eG04kJRD3pVdJIuDbujBKyg4PUOwBsqXJ1iOWhVhq4FJnC80c9r2p9UXIUhZ
spdewreYYCbGAhYHprgnTLhmlsknhhXo2DP31Gq0L3BLq3j99Ze0ZIy/8oCj
MpDA5H4ZmkP8BdFNvUgZcqAKJ28Iu3fMsFLwY21fl7L1vrMFRwqa2yAZefyc
Qi3W1sqS8b1+fY5CtNTEyJbOlaoamtbjSnChQzU4vkMIQDKK/gtA4fXyhT/4
x19DbaguPjtM1QIL7U542NbILxzMt0+0f2Y+u8Jqa2RZFbFQQ9MJwfYU2qqK
f8agrMo47Ik88LKETfbU62YrnPKpIdvPL2NQzIfgwtAgbarAz2e2OaIKHThl
80BAL//zlBkMMSL3VZoJ0C0QeBApZ9DQ1Xbwt+acpcOp1hllaEUxvATWr/px
H01Zx4upyAdKWwoZS9WgvMyc+1Kyj/nPnThPx+iVHhzxbbPW9LjupeoYtf9M
nAVacGdDkW9kDyZ3S7j+wNNO5xXCd+Lh6OCCOnWsQVKLZyjVglAp4GdvnYOU
k16K8+xONsNToxhOVFErlHl2eXpZoECLCb3iBpaEkync1TpQmrRjHXwYzLwz
Qs4W5p5IeR+sw5o98VNhjFpJmTtrQlwtmGFHALOo61gtdQPf24fxjRYinMiW
KkNMfpfC3N3ultsxoh+nO0518RVNWCk41fy+JBbX6dqcZPQrqP67Q+PRCX6P
qcyGsp/YY/GZs/OEHqN5wYCi5Mu66NbAwaK2CXMkSYuma1UDFncJ/ifSRZ/z
z9rRZs8PwtRJ3glK4AEFk8GoN34ffeKh29DWjzdt7DAjB0DgV9T2xVTnTMHE
7WnGw6YwUPt0iZGwffqW/cj1Q8wUXqxO6dQZhfDjSHXQk2dYHMo5KBRBzjmr
8+svPfo7LeDCAr7fXbIoLrRnWBpuvXY+85H2OFS5im26qWhDI/kvf+QlNbZw
S/Y3aZdzgPAzA79YfPHy0OfVmVIrxJQcMwhWIHxdqYkiRcErY8oGLc+GQl+R
uNxek7l8zGHSJBdAnFffCU+Dbu8PKNutc9oqEAuJ+r/NftDYPgDMBUmiI0V+
h+66euhjQFsfNEIvWDt7zjUSpAmorwP1q5xXo5G468de/yhXiZz13eNhlnW1
/AN5qN+lNQf1S1v4/+dHSXNKv4640YRcR/oaz4Mb7YyPzAvzTuh8oRjy4iAN
K06JwKOTbX5SUBTVmg4RKPgQYbt4R8KXIE4z8HN2iVy3pJCwwSHUetw7hDiX
2ZOcCNzZLxjdrPZy2fpJYxQC8jutVMwE4E9AO5DBXj1rfiD36ki6Rl9GQKe+
IgJPFAliR8wHCqaTB3nsDdqjzC6JjRwGA3IYPZ10Jrxyg1J/kMn8WRRwzjZx
GPioxIlpfeFB/EHrh3HPTT3XvDrnIWy5LitYI2CZGT5gIneEh7PzVCl6GjqS
vPzkBBJYDu0vEf/KgKY/m4FOuPwcjzFkPKBlafyZRAYr8tkP9xnSSdcbDiYd
WSoidif6VUDuruXVTcyw9n9xML9jmX7jFrTyOdMGdvr3wkZCoqAJilaUZ0zF
isdusJuYvPGQ3JOeCQLHOVhgGMq0j8NHnd1E/HGrH7K0tw1XET4jNFcEISXM
0PRtbiEhYV7MYIxHpIkvlVEqVs0ofVXFnZdmeJxYmirjHYdQFT/ULgNJX+tC
Cz4J8J1DtI/sK3PBb55XmhOyzheQx6K326YRYTKBaJFAsnrPFkIwR/vu+cnP
gYoqbPkCO3e87ew/86IC3C72+dipCB1GnEEALmIDicHMNlSX5dKxHT8nTsEY
/xaFsHs97KFZpWGMRQi19w6rGdlvgBU+nRE2q4HhGNPaI2EdWpUKMnpT4zMR
v4JDX/7nWuFR4kDgDLv4GbtpCyan9KE+gn8Zhh0Gy6PAg5l6aZ57rivrdMev
edRmmSHyt2nsgzds6V3JmUvMZHWHG+D88Zfd2ZG8MQJMfq+tliSjzGLfl//F
VIppSZZtosCUXwXKGQuFBPexxX6vyhBj8OQ4pcNSrRAZx6vP9geweZ4gbXPK
FT354RN1KfL/lYdhjZauxlAmHRALCewNBiHjveBidNTRAlNI2D51uKKBcVst
S1AQ9GGzmsyXn2z4PbjGoldPD779TZWJgBW0XbfvoILcPbeJ/SKC0/ueMXAq
KM5EfryYam/1CZrAek8yA6LXsSMdKdjVzegAGDJq8Q9bGywa3zV8yl88n1je
HGEdQHiu79wRl1WgPxhSlK21tjl+FKCNEppkyr05qOSurVd35v+3xXXM6XRK
B8S/KP2qVKNS5AjnFw36JnLOXcuL1I2grWV3XI5FwmxV7T13vVKLeToVoksP
h+rl0S+fHQbgFjEkEmisfo2D4S+rJvUyYKiSz5ny02G8TyEHan+QjIu7KIku
oDPd7EipnKIkokfmsxA9t03Hv1hkaFoI/lZ+zLPMkG9g4T4Rv3chUf1f4mpF
Rw+TRfCIebOpnuEhRjc5CVeA+5j+4H6IAWI1eIfg3pzu3YV6gTnlsDEqJYTF
4bIFbETx6fTVNxgzcwAbV2/YJuv/a1Rt39TbR/Xx8ydcvZk3jjFH//Rs14ha
Vj+gf9aY9o8oYmwdT76VT7N51SdfFPpA4Ee7p7JayYmfMJ5nA+17w0hegrxb
5fVHOAYmuZgvh1NmBdBEX09v/rPe720VXtyjqidr4Had88JRJl58BvMaMytH
B1HCIFuUjlyRf2c+vZI7KeoE8vP5blY/vfBnYsN0OuNEAXpE4gWZ6/pjMbDU
hPFowD8Wd21ofGT3qTMYsK5sdknRoVmJELfMnVkcZ3Y3Fsnak7IbqqWhx1HU
M3TSATXzDwjQSbK8LS9JvVxNazATNAonyV+BxcLxBiHvFsPEcAfQDrtXP6/O
fTolAQLf3brgefok/zNYxW5GiDC5sw1Z4A03g900LWXi+GH2L2osVzR1nkgB
voeew381akF7w5Uncwj595aRO6VTysPWTX3fRLbO3FKKnvAUap9xLCN5WLbR
FUGcTLl8/6iHbMn9jz9Bc2WME+vPO2UFvQtKrRxVFaDMAtfI2Y/zYsc0vLYe
6dNC+y6mxXEiizotiO2NhrOt71P5umakMkxO8HcvAddsNbp8TkTIdldEDlkO
QHI7zfyMYZHHZcwpr6bGJhgqnjOzUhuE4jQ5OX0e+usfN807VJmLBoNK5xh6
dKJXtwDRS8j5RzduZahyAghZSMrxnTUnrx9I0B7f7wFxeAIne4WKtDrPR7Ei
Buj0lBJEfV10GF6dfYja6oQSb+0Zj48heeBkrbG054oXATIwr9crK0+RtP2G
qUfh8IcAgxfQ2W11Y309EvHy2HY118QqJ60EejNpQ47nfSEsMv1iv9FoG3fx
G7KENe4B4Y9BCN5Zq+iWxRaAYCiI27r+gOTM3rYsxjuSSq9m1mo6XqvnysAP
W145nR7u40mxbB6Ge/6e4dKxjsg0jomREwqLwoiJ5V2DYsfF3usEB3M/tQT4
cOaCE+h4iLPN0ukYrhqSDIUTnaCK/DjstQuMOVSmhO2kceWrzCUJLnvbCpxI
nCJruXY6+UgTFqEK79mVh4qm+tkeIbIOpJZ6j78RXXtmuUj0tXrw3ZMYLAk+
2H/Lb8q+gLIIsWAc1pqKg98ufFgWLnalGc8RZGGBM9sL55IEM9Zs4xAoSiE+
lnemXvY6Pk7Rv+Mwa8mLD348hGhb3o/D4Uvov6ILuPhbPC7Tql/9gByjqsGV
7k3XLSIojrNDiF2b++9VtI+fuy76XYmieE+NJ0Qw8iPHfFov3BwQbN5Np+i+
1bWfNu6JiYGp4oONIYgqaRTuEgMqWrnQDeh6ojhe2rxmljTful06gYNl3YHD
sDbGtbt+pAKld4nbv4JrlERx25YcMkUD0iAOErFhCVjqUq2hUScOJxWvcltw
6lzfbWX/eEVOyCzewUR+GvLo1ncWVziHho5bhxrWYj3aT6gPVyYK2f8J6ez+
/n+4m7c42HoFQRKMYfQcyOiSoi6PNUIelGjisaG87ZQeMdGhZwp37Kkq3ij+
3SSVR7eMBAePk1c3i59qhpmT9Okx3/Bn+rF+0pH9YerSCH4a9TB6BkOIPzjx
8WT2y4On2uz4KpBMPGlF/VyOONykoIo+id2TFoDynebdZ45AXFZyBFNCCq32
/6YcU1IeK3DFEh9yxjrhvE4/49X6LuDVTokn0YS71/d8e2yKtO4rXJdjG09F
LKC9BuReoDhr1mKl2IguLVMRstdWdFbHz87ite9U0SCcEtmHjJjn9XnMYeX6
1+lQIoXLC3J2DZ6jhQ9JBu1Vr28BSFQEi68cBsNGJj+7CCTHlWi1PawdO+ry
o2khPtoucYYo8eoYmDel6AniMsK1QUHaz4QEq5HEF9DijSkcXzxsJwt3lC0Z
WCHZnX6eem1N9RpDArs1zwcp5hooDuZyYUUxGBkjdwxaQnIc+3L7MhjzE3kw
Da+BAxKYQ22dM6zP/Mb6oN4F3R1NQHwmSLu1ZfTeXavmhxT7ZHrOnRAcnSVw
qwmR+qMsiBPftMj8Y0buni9y5WuXXnkHVAu+BUwiKMslEJy7iDGEbXuQjWv6
DKxSRKTFD3N5WRv6bIekIot3TANQaBv+T2m7KyzwzvoNXDIAypKnB7jTkF9s
SH5sqsXbDPQugMBFSpyjChQu0IynCx0AI4QhPhG4zLbljjnCXb/SCwXxyFHL
BlrT7lgs3H5onobkGpUugkPRNlM1oH01AJ+8v0Hv0eG1tMxGmVQGiAwoO99h
QMAlG8PUFqi3kfW+9dWx0U0WKRlQqlscWsxytEozVatHAnBBFwpHGHOJOtpW
t3GTqcIr9jsnWV8ztt4PsvU5usCGuuBhEfMrJzXJVZsV087EIzBjwy/Il3We
sulN/TN5PXbz07zmQn6qQfGTvlP7AMjDtZpvwH4lAmDLRoZ8ux4DLPWCCrNb
z7l7+U3I6b3nCBd+QcG0FHFQVRPOUP4EswGy8zrw64iCDKjqkh6nRCd0KNPx
TFDT0n5d6AeyhyV67pfLtK+QUlBTNokVAt5oGkZNGcAShMYROciPR0VRHNHw
96vauVW3HrlEV+jbN+MkPGu2QYyk1YsDJm/g1u8TWo4spAWRcCN7OyHhkAF5
dH0v7114GF+3DfB8JZAMK0sgz+QnI4181oNUp2GZXFtBRR9ElNksZtJ2Jh4j
ia59Za3fsvmhEXIxUzqFGcEaU9MepnmZNyi6tXFByX2PW5/b3r35imNY4im0
83kGvGZVQqizxzkV4cJXhk5deG+yDb1zezPeLUMn+wp2eFD1iB1iUh7pERTV
kuQDAns7f8rWu3GajlAOtyDmgO4KQlGpb5Z7SpyJhcOriT8g8hHX/+P4c2sa
3efjvVyeLMKi3ueWC034nKouYcKpX6Zr/eipLHnE6pF+3UZRnO7rEJhkJ6/X
SzB8+jy3gH+WHNLt4cLNlHr2KodSiv7PgAKBdMaiNomXbWrN/Rj53B+4CdCp
Tj1tdUtYGzxbMUrs6qlODPILBSZk0CQ1u1jwR3r+BBghklgp3XwndALnkXN/
LtAA+v5vJHjGTIycMPbvM4YaSYpjN8dDfdVPZ09xP5YxRarfD3Jnsk+yLkjb
9FdNzQHy+2ZJZWyrx9GielfcOLhd8UXrzTnrUBh6L1E/hOHdEZWmhAShS7n8
3dj1w8R9oCnh8ZfgJkHoxuXO5YanpiyEBXmRBeg26JOZGexwbIiS2ku5iB+x
uRe39w0+1SP905zAMmliLc+FDnpSUfD6tWuhhSHZxUnpG/ucx/VSzS7YBzzv
mXmOuDHduop0Z84d7GMbA67MRiDxeKCYvOlUwckyAsLFtyxKHnvaRg5J/0gY
ITuyLwnghtUvalEuXe7szbCSBG9qczl+3mYeum5IsdAiLXcC1KDISwIoA8xJ
RDIlQEKZLiLBxcixJ3sS+B+AW+C+RP0c5IVwKDYcPOG3BC9pQp3UE6KO57XY
uq4A9x7QiMCSLfRrDz3ICkFvG2rHNdlM94cSA2wk/opxO61ZKUDz+JhLzIok
+g36Nm3j79l3cLhwJv27pX6prpVQSfn4uZJYTmacLumGN8eG1xa1egbkO6S3
MCG1TyDPnbGMohZumfSstUfaVVmh3su/YQXUKo0Ipp8wa5nAfT6N3psII72/
kCWuHVd0S9IsmQWe1seQFdJS42JfFcyYA25we+NJlj5UXID9RSZ1Sf2Stzww
sU7JUNoonS+kuGRkWht40I4wl0zJGpZvCY6sC+nxXzIkXV4cSbNWRiRn3ovF
B+gxW63si4e2nWMCZy2GUojDjsEsHjnbo0E/n/ROEFeihLjB3NRA96nnZldh
9+ONdgro/n9LFokzgS7XLPNnf1kIxHBxOoB0G3mTtn7zauhKOHf2US/7Ba6w
rCHYi3J7m36QUxFQAyx8JSyiZ/Fi19BqhpigdHTaV19adcUX1CaR4VD+VlB4
d3FSmitTflvBrNqLuW4sSIAZWJfEbgaKEvDiIvhFzCaes4MDPP3lpzoDtKO7
BOocst3J79qvTdkVg9VR08AU7rtGeGEdQXPtY1X0onQixnJ6lLdhdth4ZOG1
CamFPr0HKNHJ932jJMVQBYT7clb1tDIS28RJaPouhpWQdsCc0Fk8QN5685iC
ZR43vu9ty17KI4oUfN8d3ARUfDzmAzAB1fjISVP6zIrQTFY3+1Xb1GIW8ETV
prhzhr1a8Y3ukHR6O4daMLr1pag/VmdiqZRIfF8KeipAhU4aH8YYtl2J0E0N
Vl85amBxltQ4z/BzsKOpHxyAf9nl+WFywDduufUw8eqV+DGHPWu2T0Q8M4Kh
j2/ZJNumPON1pOf8Kb3/45PHiDwn17qm4hLzfadfNirwyYU6lt9GaPLiiM3y
FdewFgFgCjbeSQTKjVTgEaUS/fNSigekH9jSOa+/kVuLVvcdqoCWBGFgFSn7
/EPGeMJDwqydHBfSnmTq5ZLZ3CusBooqCkczOYPQV5/jY491PBDNvXfI3+J+
hZcftq5nBkVXFnzN9kbMKIqszst6tZtt3Lo+/dZcnQOgPiznOVbjbBFucith
SUdet9TR5aOlVJOUIi9CDKachYYlpr+61OENIYNGibi8URdaa/sdzeMVToUU
V1G9HlP7SND5kJ98Bzl5QAOWBRENKVT2w9aakB7VTmoZOvADIcX74G/3dm+U
Im2m31VCyPNZwHJxk75MCxlNWqbosokixcWDXOU/vmFtBOCP/tDxQTVLF2fm
+mW1vY8TyesLQuif/q+mtLfZVcENZAtSQt1KlcaA4gggcF/4IxCQQxmPetZv
Pz6XMf1rtWDl9svu48/7EwZLOG+GvewiYgM0uKOqroEziFXGlSRmbPOPo/CZ
ckH+1aOcOCVkCm3dihVduumS4qDfiBk2ANzQ5IMWOnjsgRY5+CHRBpjHyT92
Zzagj4CudLLwV0jt1tStm0eN8wMS3bmIVKTbga1YerJ/e0MOCEGgN4NGh8nS
5yIvyEIIM/A+nHaLsqoLta+t/MvjkjLG1zAw6n0UeDGlUOEjrghrpxY9TyB2
X4utcjmwY/XEfujhXAGs6nZpfZ0KkdUNVvT5TSVwspIhxLqKD0b3neMHRTix
L29eMpPvvwIJCTxe9Gbd2zOEOn9ldZ4UzsvoKcdKOW1pPrQZHYkzbvx4IY/T
P+iQV9KxzbQ7TSnKbkTP4413MdudLvfvqaVcVxqgo1IHrmDPSDtxOlQycXma
X4jc0YCybdhFafHaY2QSeq+hyAmaGaEEta0ZZmJ/4V8FOdLsRX+1ifPc6cln
c4N18PwAE7bdg0DaHgqkr+UI0/l1suIFIZYQKjTker7xYsrQDvLa/W9YRZLw
w39UyG9BxAC7pTvmtoy5HThQvY0jJ6pSf763P5ypk4t8IZyWdr3UD2R7dEjY
RVnjBwpU9H/jLSfJPRi/8C779INTDSOPoloeZHzV3p9iew7nhWqNxH2//rXz
XspBLyrJhx8U5sZBsKdWRw8KcX5C3qnzHQ1+uYy1q7zcKz44CtwXOI+QKwE8
uNJo+SpnN4xoqo334PUccoaWYLwL5G+/phKwOwlVarh4L+Xw3IWgK/3H07S/
+TN1dLZPzBBEqF9b2IIA7eJw2nTWvjdpQOJihpnMB7OcGfN62amUH08O+G0g
72Ss3xklYnZHmY6ZU1Z5VsyiU8SbdM4OjM0az6JzlUktK0if/pPyFm2ZOQhE
l6klsPu+/eSu13Y/yi/+qlqNjqDtsNTfCqhLJ5YENJrykv/oJNB4TuFkvfoT
LDEjzV7aaK9uFZfnQvpSOLDFfE/dE9UrPsZFlS9DtJp/9zvVPiVRCEUMVT22
fOvMW1k96Ry0AtucwH+GzfeQJzgTG34Oqtnw51NsBpih8Sltk8F0sMBTfQHd
cUJDJCUcSvFI4KLKXSyHf6Ecv/tCm9siFy5UAm1moj9chdXKlPGJdlF8OXQn
EO0ynI8y3SAu/OZl84KGd3wbg9afHx5xJ/AX54SIgh3kHBVWKwGnKfoWG3Ej
iAP+tf7TEL/gqXaXZPpo9XiX+6Oz5Dxe1GC/jYVi8qwL4SkbQU2/E9k6/d6r
1NnS4iwhk0fucGe5Mxb9qUZh7TnOGz76JKkRq4rYR6ZWVCc+YtaNDp+QV4Xe
90S8ZUGoVHu1OT0D0TCV+9+onHnYFF3p6dVhNZJkz1ic9WF6O+rB45UdoQuf
qQ0oh4Dkj0cdcMUIz4JwXRhh8px6rriz5cfyjj8KH7DxQKWhFHzPsnyT/8tz
Cfi1ikie1hnc+RHpub6pcZ3pDjp0CETegp0X2T03F/Np6HzJDe5Lsl3AxiCv
ojBDybFb9wjYKgTkU54Eo1nL8s7alwUrYQYCqZbPx3F1Ldt1ZjUKPxNQ82xq
5wtL4waBf1LwvuqjwAnnP5dWz9tpblVo4NuFaKWPH9voeG4NCb0rt7vnWJ0h
iuXKGrHAhScNHnKUWM3T1BW3/OJ1s6uf5On1IOlsue4A2HVt/eJb/Ea1Y4eV
ZhfTzbN3nU90ZP60mc2/t1I1y7yUASMws0EtNfbmdVF8JOweEljTXjMHkmAi
aO0HZK5po3omf5Uo2ywbCBRxxHG4j/FYtX0QmBnKNwn7/J46oX3ss5hzeEbs
7TWhUer2OFYGmqaaZjRp6zOQurRONgSoTyLAJWsMb76pc8C7tP8j46rwyyrr
o3347VLLomPM7JVmNuMw7gvKkY7Dc2TvNni2frbOT0You16Xos2ELVtYl8IA
kD2T838YpQODwTTOuneS4XrQufAznqj8FqxSKKQg/LxoH0cJnCLnzG16UYnX
7YO79bae558ebILSXdat+cfV8iKdCQNseGUwNiT3Mb+rG8z4sa8UtF9ef6nY
QJijcwvU5MDQCe8TQXXcplt15Rbx7ZWLOuDMF/zofBmGcNt7aFN3V+Bs6Kbv
c2M5OolFhSTC8MAiZeP5cpJ4i77VQY51g0NdvGwyVRWxk5zbArbrPa3DDqmu
KiSyDT9eUAYtkXej9MJ4WY/GBK9k2T4d21lL7I5jBEkUwjqz1Rf/Q35PrbkX
sWkebkJll7f/OxVs/TC72W/5qX1lT4i52OL1WNfCWeowyh1R7HZiZw/ed/zE
qT5qqWt82aSn+ToHNM6RGzZZLh2kwy+yXEltwJ2/VmVvcN+CTVRvaFkjmPA0
EdKxr/J8eGpknGa2yjQ7Q7qDWYysfhJ+ljo4f3FjZP6hn+AaCMTyY6G4OL48
aIMaC2u5Op8R+TuV2czP4ltmA5NNYAx+txRJ3wqT23XKzVM/DHxZcEEciztr
LLI+le5fy0fmC7vyGpU4rgBe6b6+Ia2K/0TKHb3GKHTlvk6/3bMxial+0TvD
LcadQ8Y+dBQTyFZvpDwh0dhtoG+4SpxtExwFx3j6VxDXCowPkLrtGU26mowM
z3l4ME5ZsySj3OfkoErK+frhnQEWh+Ob5Y8LvQOa51GaWjxUiWl8kQN4rNCb
ADArqLH2MQDCthlAM6NARU672+dWlBwciFaUDL2YiwNCBoIEpjKaSxFaZ+Y9
9iybNITa9ZZE/snMg6nYhc4wO47uKNoUbImfB1EvVkp+hlL5CICXM9c0IBNT
pcQskvsIEm1+xj+n1bvNKC1AGyt4UeDYNVSViaonjlWLRs9b15bt2G+V41By
zTsOoDSEWylDnr8mL+1P5mX737UkK2pZl9+ONESKE2/T3f9jXDtTmkG6Uep1
2E0GNdCSTHLuxpBpwNW1Jp7Ic/uvpQ/kGGt/hQZnFQa1jVE4eq4pAzjciBTW
BqFP79+cY1wMV6wKoxx0DlDfxZvSU6wK2qgFkUD3cNmwHglMcReS0pevSTLF
lRNPtRU2XPgzf2AUj0Atn7DTrvnU9A6o8h8m/daoU46206uhMrWBaYKrDyJt
jGfmZIUELXRH4zR45WUiA4OoLBNr0y5UBtMIZwSVNExaKf7WQlEgOw3fiIfM
IEgzfTePUXbXWs9QYsyWtYkgGBHC3Xd2ZvuSjNQrtkPEGAFs56B2Tygh+Zdc
jNUzAIZNt4uQKaP3ArXr+jvPZy84Ceu7s+kE7Y0kwU/3tyzKgNDCDGroWAth
IKLp8nc1s6lmaMY+AxoL2jFH1aTV2zxS8cYabU9hxwxDiUFtRBnkRi8eJDo4
dtnIL4nYqU+eXZ2vFoLggKNR9V2C4yaCQc3KjGa33vF769u+JH3HD2avvNCM
u4kPb9pP3vVJc2miunypDCCrGmZg7iaaXcenOo5Rr7W+C117F9xg8MzhlLKw
nibxupenDzeCTRjzmmJM56r34rV853xxEGdWgRc4HviDQjEIYavsv00P1M1n
h6kXBjkFooahS0qikU2CudwQreTLtMThazhc0fqqnec0bnKIlPg8Ollm21Yw
/6F1zU5b2DLZOvUcwXEWNDnCHl1Tjd2WEKh+StxMCSxllLq5hmv6v3BtsaPo
OiVEbowub9FePMHX8cPZF9Smk3eMFURgo2AWFMzJm8ULCv2toyKFxJdmNrTs
HIM1KDY4nAOMFbj42UZbSeJnvzqmaOClf7nGzO1pVnGFwmKzKsRVzlVp65hd
NjQQwkoCzC2iF7kJrmTzv5pIvwC8bEXo+ilzuDQT3D0H/GG/NO+Lw8EZitY6
7JW4VYW/AJJpLfjbHfud6+zLJm3d/9yzgECJnWrtih+7SzOX2KgI9VEhuFQ2
o0tZwzrM5LJwc+SFcaSatJSOwyJIKlqX7fCJVXTfI2QpARUZWUW1P1lwBaT9
RZWaotXUD6dS6wT8mTCyn2o6PcOhgPNGiMsYq3IZqib+NRFsaKt4hLXRqtCo
lk4p7Z81S98bH8AqKA7/KUzQsB95YHbpnz8zHKBlK17uA+gDZdtJxkkpdvPO
RBI9A1POXYCfBNlx126Pa1Fg0rILRxHnDkT7e8MLoZSw4JeKBNXJMzHCHknR
Vit/w3y2ekk7a7xybJiIT4ComMIJq1q08kTgoxHd7EoYC19uD4bEMmDKD7mL
dEb4ZEpWtoCOiiHigMvfJ7szGx628K52hxMVJo5rOiJXyqXb9xNrXwXncn92
V8pXaUn++5YYU917pVA72MJbzQjMlv7j5RyKvwjVhS1cBZ/nR1NXS9AwI0xR
DwGOhIWvHssdj3GUmDVcDRPKgfy+xK7BtsvBkAP1rkqdL++YYf3Hsn5ZTlIG
gKpBohDm2iXBT+4vtIfUHZcuKFDItPv1e3mXaDWbt9z2y/kaGUuNP7jnINXW
KIbwhY0a/dtPLzlXsmoZdDBJ0ook3ZP21CMl30L0auvxQovkJkdNxt3SpONT
BOgrRcR5T2cKf0VPYUL6lE7qqXIFGSEC6Eqe3tiTcVUofWd0kv8llZZYTE1V
mlcqjMOmfwVjg/Qc7MKk36DbFhtb6ULKGqpp+JNnGCy8bmYxRFWa1c2PLIsR
NkrxzsLcFGaKzvcA9FIMFpXxO+E/97hBE0fkZ7/Q15HSmwllA1GA9fOvYTT9
MgCNDIkZ4Y8R7JbGCD5auYJjZqczypzFcRcFR+oYBpL9+707dS/sddpe0eO4
YD+A4K7pvYuWRB6mKnHibqfm15nblfvGT15BOKlsv0twGuRcgyzRyxXEbVcf
2G7JIGGDyEwTmzl/Ef9cu10mfzA8MdNOARf+Q5DW5lliZO7Ic7AXya4sEp03
g+F7ZnLjwvILOYuFJy2xlulFJeAXYvtTvRCJAK80JUHVsJIZYjnLc8+DBzIi
iOk6HNelK5mR2Il9NiJl3k3EIQI9l42Cx692W9RqgiIclxnx/SZheFfhJbHM
ldv60btNEbplq0vrNd9AxkBRCm26xw/d2S/Ekw6JIvesVW3MV5tlDn7+NCs0
1XxOR9m+O9iDE9EaChYGlgenuRgo5PKsvUCNfTTZRgLWSiPOLgCSeiViPMFe
MXZjCyNvY4sOaMmohAZfPX/I5XazAhhlt2Stgxhr4liAMkLXpZYyKV+FX0Nh
SIFNoOoTT7ea4wt/LURv1RcY/gIjfTpyTX8JJ+I5EmqmXdPkY+mQF1mL3Czg
PzAnRilbrsWuq92OEZZOJE9/qCNhOoFnPzMdzwq9Ne8SDcGpnyN/+JZSYBPX
CRdHkpuiCMTYRfIMSYRpX5mw7ADHu4mxdpds7QhtcFQzPtehbPD6AMGAvbbK
H3cQalzxt7E5Yg6V5pa1YZCjoQjvj24VouSz+kOgWTlpVnwHSF5GLRAU+sOV
aFN56JV2MI7nyQRzZ4O6/ct7ObOmlu853NyhoHtB+gLUhf7P1pTwdQERATOg
/eBMBhovQmfFyy/BaCJAZp4THn2OE9Bf96XA4DQnCXmJjx+Vr9AkSBbbiDwK
McRTcloesp/QGnbvSaszRBPK9qg1QNYHnIzEm81Vdfgv1x6Mi1y8FDauM4Hl
Y6ulQ7zJHCY8ASDMVahffMHhBouvRKUfEIBjcqaTz1aWGmiFkcdzzaXwzePK
p3E0mgUCbF1xOJu5RuJOcxdECp00h7lruVm7Vo8Qv0+i7GZJ529YbpEbZQxr
no3DnZGQBt6AyFSX6wDX9PE3nwe2fgQ68Rj0AIwSBrWgNGvc1gmO+vhDanrN
nxY9oyw/vlZNM4/EihhnBB7xqrraPyEQ06/5jq1W3ei2XaK2nT/67ZZ2NLVU
nluEVl+LPCu7N/uEHpMESaBnOhpOYaKnBCsDISAswAxEFt39D8NuoZaWBSLr
5wNdf4X3RYHrhHKn0Kec5wN80GfW9H4LyZHsI0+kxG3EJflJE3FDnVoSgnDP
ooiTnEhUMj9QU27Z/w4Ur94a71M5EfHbyI9OB0lOcwMeQe0GSH8soThO9tGm
njT/wBDLAhdINPCFZDuSzZx/f0Qo0QgGHIBe3ZzKPboJ2nqlJOKeT8Lv/YmD
gCcyMCxyIDImJ10Puj8+uKK+/0ouO9da+zroFQE4X1iPz+Bd4QYJ9uuURDfC
RGyXCMGFCAssuXGdGRVmZEjBskUPc/JuGZR3X2JDOjUfpftweNcSTWtT9idE
qJ/RRHukiLm1zQQzGW+GKh7DnyY+8wT6vYezmWXpuQKbn2CTgKGZJlqujqMS
6CB8U0rxGXrNZY5jv9op2Pu45QhEABhbinXcRlhvR1obYWiUnmfpOR0pov/k
CGO2t1rl9k3VPfXccD1wpVNaVe7hZcKMoZazy4YnZ5wpttlipfj9/Iq3SQ1n
ipeAZgvM+PmbVJFJB/GehQqgU/tTSZYRN1Eb3qhYqfh/67XwuBDkwKhHtzMd
QByLFSR9wl7wlWdw850/O/SuDpGRvESr6NIl6KNOZ1AlhQQHA7eBrVidRkmj
UAq91/EI7S2wdubrL5W4BAXj/3zR+De3rRXx3V+teuYpJULWWeE/ulKgKn9F
3dDyoK24rCjm+Fjue4mlrTAvbsze6a2KjeA/BZ3u0ixbJz3q19xb5NE8/iJq
t6gti76+OTd1DxsvhfoFa1xUThYzRd+KCyR2/F5ByGh2sSqYsyvzOKFDyiCo
brLNl9g6WQqUnMS2oxnfj59mudnRuMDONX9PO0f81d7KUCLJ8exKYqgE8+Y/
CbEMshBCpQicQI0bnfymm8dYzSQhPMSzMCWYVZrycHpqJn0RLRDzFvTS4GIp
YZefttuxF3pJg4GCWgTkZ3shIDBynP+v+A0VkwK3ceqk6G15b6kBBrh+WaUd
XPFCLsqM1gQnQ6ZhJrh7dZglUh+LmgrL9gXf7GNWUCVLICquU70deQDujIue
tdzXrkmPrmYzNT1er3hIWr3G52bvnHTl0XxAij2G2RfcavPN1F5sADP7qdEB
le0aZpSZ9/v/0CzTacB3MkAQQIXPyVv3rHlRMHZ9rje1FuVjnfv1JyFuaPLv
GvczVRk4iL32ta/MrvThwcU0gYy6mIWjdNceil0gL3jYnHmt/jMHutX1rgrC
8XYBGVNee+PcC5JxhmE3DpNqjGPQqvivNdHRujiMRtPwfaJmUlVn0sBYGVXS
EQ3IxziznmC2D3jj0Gbo41B2tUXZFHzn6DTATs9y+HGwPvGl7ksPIJjtuaZZ
x9Oe/feQlkOv+gK/umyYOwJEBniXqnsdSdZurchx6iD4fcL899LVxaUmP+xe
kWujkvr97gpRFBD97eMhkhU+2Wka2amBQUsn1QpyhVxkcEaL2HyVtC1uBjDW
3/L9Zi29st1KvJS422Wzgvpqb6Hc3zvgMbeQreFPgu0uD8SMapnXNUsYJ9c6
duSam5CQ6APCy9fEldfktLeZN5p70Px48mIhPTzmpNh8Jo6azNAit+jwW/qw
X4LUoESiu4GSYm2llRwIBcrtbJ2ePu55CYLU6Kxjo+2oz3vsUWN6Aa6ilRq/
OfVPdd7dx4fmFYJgPqY8QK1Gja0jTGNl89ebwm6sG5v4Xr3lKqA/7+HO7wQt
f5i9LVoiAR6HRYOj1rI3K8+i08ZD37W7zqUxYzmqkPHdHyiiX/8IFMM2PzCh
9au4DWEWu5MLqraFCx3FMZQGSvSkRYn3KjiLsvAxxu3G4AkNejdUS+8UQQlO
ygCJ4xNVAj4YviGsTh4BIYTPxgpkVbE3GxpiDBmrG3+ruZnEEK5QcBTDosWp
pazkLQ+n6bw+yxlKYfiY2vpR758gex9t8S50h9G3vlbILa5kpQEZnSw3U04i
HRsCMEbal6n1nOegsRKirV3Scs/tRZxc+MWNDq5jSJeZ7Zpzjii7NbKANs8X
WiHZC4tJybqjqUR9VeUmifk5mkDV83hRJMJgFXDFxjqLnB2PaV8ZtSHxBm8S
YSDiYlUcPgrUpMgX34YrpTpaEpSZ9uIRHCVJ9mzs/vF7iSwknqRb9dAixoP+
b/lZAX6rU9ZttfroOmS+VETNc0gznex7pyZs/92/LPCllNUOXdvrAovGbDd6
maNQrDm1xHtIahBD+BBo2/bUHKYcNb5EH0vYyVBRhXdIaxbUKzeJ5Lz8KOVk
NQ3HDvl75SXn04pwqXfyrP0xxm6GjrrrvZ1XrtwEdpw6bIwhbkzuyUHGK8l5
oiV8RnZN5aKSFGgo2wmQrp07BjeSRd6eM9AUSULDN+iusOHrMHja0GCn5soq
LbJCquZv1108uy32E/AIxT4blFLPKweb+Nr5lM7/2lNLg69zfoLm7nmry1cu
tUwtChrdjZHbIsv1vI6pFL8weTjWyxUJrWGfqaUunKGFzaQm1wirvnmlX02a
uagocpMyVwgj9nmB8zOejD+hNlU506yKSv9MuRcvx/Fx3eQ04xLFXZqvLXfl
U60qOICiyCuXkZHQggyqQc8wUxwNhbMRJDOthd8q8bNt6dD59YiXcimUEHMz
cVoDGFubVCw+Zy4YHRLhPToS8lDAmZRoXWfSWBc/NIuT8g6p32m6s7QjLCOm
lzdp5HIlikcp1UYd/8RL/BfjoBWLJsvw+eA/FS5Vj2JvPI6BMOllgPYZ5tBs
MnJuDyLRaeugaC6Ip9WhEgy2mSkRHIGTItSQ5XRDBPBF0WoTqiux70qmblGb
YKDj8r9uLTMILWsqQ7cCV5YcAglQxWRnoUUb9oQAKzRyyIZQBltYmpfKM+LN
tp1hTTyUsQATNOHU1firBNRKaK+25fyBacgRJBnX5JqcTutbfRVaQy9Rmm+k
YLCbNRdCJe8ujUzXZkJ8wU5Nc8MCn82smy8bXazAae62phCv50cin7gEC7sH
SVEPX9iT1dKjsHtFTp7FV44lRi5KiLZisjnxTAN01/t1GMS7vL+KhdL6B8g8
8GqbV2Ne9PF0bN58BLpsUqUzWAAQvHC+0IvBdv0Innzc4i3ad9de62xdbWXg
PZHYn0vMPmJG6lRc+gdVlBnAfqpakEMkIIROAJ/NtjE/oqg8/7MSMbPNXE9C
UJ1M0hCdFBzy29ivX3UV811LF9fp8Z5VMgLmW9FiWTjSFbycVCGDIVCZpphV
b2oQVJKGlFZudvr7StEXAstBRuM3LD+oKPRPHzh7rXNqObbrUxmppN1k/rPl
ELzb8gum7NBgZUQlqBGTfzSaqSk8eu4nb5YWjpHrIPuaqkuQZPOwCiUyLEdA
YFcXMQnP/RbXShWGfHgTkQFWopyetxY0knbt65b0RA6RdtW0Q7mSxkoxAW4+
XQuhEK6sJEPE65gJhnHpbG/hABn2mStlUR2EwHGud6TSqEaB8eDiCmD0PHHm
7TLbu6fpalfWX9m89HzuHknGuON7RVEFLAw8F056usf5DmR/Z3YNL24hBEc5
jMYbPRmHSW7JCWk39Is71j25sblJ+R798GEhtxChmHAMtg+aAwhFQ+sWy6i+
ssM51f/YwJKvP1VzIHGFXJk8suSJe7LJdEpRGuwi+TQwrbhVrRFDPcitKR0l
sbxOj+lBiNalJ0eEv4pAXDzSDd5KnTEpawKQSdT7sxEnRH92pXHwU2j/EGZZ
ajsdvHRr5TdeCxMHJE/yCTGFkncYAcYDiv0yfUJ4qah6fUDXRhbbgzb4S2nE
2KyOOnTyMG74zSPMfBTmbz8lHAvXtYPsJ+MDJAuXJX83AK7ZdIm3PCymlR0O
CDp2EFngYp0lyUvXK5d+IXdBi5C3N2sCGR5yQlV4XzRfQ9T75dTE7ZAl5Kiz
Xw61nka66XBJiim52CYiSS8Qcgj/loFiFi7CBOSCf9aXcCs+760NrTOvMYd1
GLR+JyaQjri+Lai+f6kPk02t/QutztLUKrCxtfsR1dbS0TveZXDPCPMF30MX
XufD1VIa8gHy1fk6Lyhjr3aF5Js8THK2JdPfUKaWS+7VKq09vAkmoXARJMPt
XbOUzmi9TW1SABTdcqTSfTjJEgoZB7H4t06jXDm53KY6uycF+WwWgYdqJo6A
IU9u0BlHP0WW142L6CQunNTrMvk7SvjLS4+t79Q71x1akjC2rHlnhXOqQ+Xp
CQY/axbNIqtgswZ8zgL+LnAa/PGDNByT3aNkdIRNza4GP1qRGHo7FbzyPwxn
Nm8d1njJMvSY85OWRDq6ztnsXb/92Vbqz4c//N6juKKh0ZPrVRdZzea4wfni
3+2T6mImz9ifaQZl31v/myX2ukvYHzTsUFdDOPD1sS8+KlMS2QdHkiXCDCVv
igalnrXyxnJwYenVH04xBKV8bWeSJlfNTvZkRbIUq7ZFufnyeDGQU7EtjM79
kxbJl+EY6MxLZpPdxFCKwh5m9TNrDE9KAe89ZZExEDBiEJkutLmaPiE6GdxN
fVz6PqGNjPzW0ibLIcbEb3riAkg9QqSZjlpf0gdajrLvr9D0qC/WMrC8ES7m
+z/RbH4CQbCay/tfi/hGC4bNPbQe8C+ZTCt7352Dp5PvYwrzdLrJagD8/QLc
AvjhwNaicsxIfwQXMwZz8GimYIi/4/tHKTotdmFsJjfjKHdauYYuYGqInhik
4dcXBpngHpANo0JxYunnIrYUiR2KHCm8SpVbbgLcWunvUrTYGdWX8w+SX/6D
sag7W2FdugE8Fvtxbo7QZg93G4wm33hXA6PKIMxyOU+TZDcPjuaE8LJ/FBJo
r+q63hG8cHXzKMsFpSqqhhgVjn3ImlUl9LIeHcFvQt4ItHkBi+1yG7bZTQIf
uLde3JM6dShyYX9MzdSkfPaDn4ByoMG4S+5t2xY/jRlg8m5kuQ2q0RBcBYSl
Q0VYH+tKBBVvq6VPPy4k59xzk4Nn8Cb4zWV5Dzu+sLrrmUAZbHquecnt8mcd
7sJkiWFXQDIERh+ivc991BOR3n/RTH6Ce22Ejh2EVEF21OYDcNwYpXUlhtPY
M3T51mC4rWF8x9yufFXmIy4kO8V6z6ZnNoZe1p+CbTxMexDzv+vRWIuSLD0e
IJePr2b3tPwmOuQ+WQBM+ytenRTiUOKiCdYBRD0CAsR6nDrRnPOy702C3dOM
nf2i5JgRHpSwnoGD1A15/RLwhoJDJ43+70MFgcPez1mKA/gJeYcZfdzkNdDo
wcd0mfhYBebipy9JMdLeG1l4jXJ7YYEfDsukEpkVyrI9ah4nR+Nffk0ON74L
1nA8tDoYu7EKn9+rnINzzgIiOMYZ/WvqMYWmFC2ZrRKUEluq5pUKJu2NVOFT
G+LnN1AW/8y+tAIdqlie1dIG/ZczMli0kVuWutTOjVV3D16VMbnpUO5fdHIg
bWbYy4wqjJfuxNhNC1jIkexqxfm6NCo2q+C4/MhJmi/bv/H0YFqpEQQGO45y
NmyMYayXXvFt9qlaUF6cUS1mpwNg/95FoRWArjSrnva56RWBCpm2utgQs2Xm
MpwxgoSZRgAs5h8k5ToeHTbt8HSgmn7p+4uuyQPedQ/9saqumBE40hOLqCtC
AtA8L2Y1br6/umU/muVLxCyHC6+b32BtqGKoeZdDM+snuxCRMoJZIhEiQEQh
yiQER+ENekttl9WqymjdD4injiYmVE7PvUtWt+q/n+0+uyOv4YxcBAd8BQwO
h05vSWvWb7SAV5Lb4Z8R8ClY10ThXFj3vcSa2bJj/Ns8zO5xnJkZcDVueIIg
do5L/3Vb0D+JU14P9usSnXb1U2/ByisymPPsXDzQ2uhuHCouHcLg+KsYoAMl
dzlD58iu0sCqaYNsM4u7JnNVCt1HV74dFMAFABoN29fWBSqD+Sp0Xkik6Az9
gVqeEn4eJDF3cBzUqT1T/BLQTOCgQutajGY8Rpta1HxrophM5WncvsKa+ZKF
qcrzBj8Ner6fKdl0d2OlMjzyz32pAqfZc8Av8fN5Dx0dHq18/z/AhIgsg/nf
tBdQKsIuBM3JgjvS4zqu9cFlnaMiBrwT49tMdcM4opT1KFD4UigRdl+s/USx
Y4WQyKGC+Nf1pJr8uHddulZjTjTN1gP173wCkpMCW/jn2CjZBXVpf3bMUOAf
S5G/l4eV2bUhCfSq1RwVkOzANHCp2ReidMHT3uGi89UWhA3elJoQwvwd7d/u
B2lpG9NRlX4px53Vp66nPGvZSGTx0nKXuu0HvXRpVgOuA9Uhopqtz3ojvu2k
tXGMAZ3GmK8OfR66pig22yAGeffj3hzI2gvV8/BTCLnItj5ZwwQiI6JYveOt
Ko5HdIZO5ejTk/ZWsOZZGuvdVJ7kgFXecSvDxf0VKrGUy6pRCn4iM9q+rcWE
+ijLoeu8O4g4/p/wE3wA5duNaBRDnHA4TwYeXM8GO2YJbvv2Ie8nuX6XfvC0
jF7FWCJBomAcuU8hgRyoDrXGDRtvknvIkwp3XFpDlQqx/n6Ab1wBFlHC0LhC
ecQsYXwwbPmegpLX436y8sL5wu5D67VxecvyKD9+b1DCfqJhxReu3Y8i4eRl
Wkm4U5uneJSeQdK/ZPsMPhz6dn9INTUIv5xqR/n79k2YC4qkOw1h6qequO9o
PJtr5YkN2AfN6lecHVETlAfGhb+6j2e3Uc8qOTR8wuswMpI4gzcUqB5STofJ
Ioxm95tJW+1VBLBuhJiR6eAqgExhelxt9+b1dtpn6ECGNNirXVlPKhfe6BpL
UXTlHMEeTCsxO10MWSba+mzhoBuM8JM6pthokirqAnkvFz+cruv9K9BQPpWj
5Z714G7ke7hRlBJfgFH0ppvTAuTj13PvIXctzuiJrCCIXhN9Kd5ReqnNNvyU
OMDlm29pVv1YF9kI/BZcMu8PCTIQdzRwLn+AIFgDpKU3efZX4gPGS3bxgd4O
El/KiReQY6+WojJxvzD/5kzlWndrkSQg2qvOCF6Lh+BhRFWl5Oz4KoxDWLG7
JSa51sH/FGSvvWDqzGQQMMpBB1uD9h/CklDOATsTM2BzgPuh+LTcLRi5/G5g
xf14DOelPUJGhVPxoerR0wE0R+w963Djh2CMS50b3bfzBe1I+jTYUl02Qve9
gosm5c/+NibuXZrrIsA0KGiGj9LfcHkK77EtDEgeDG409PneMj8gnLWIRwfE
gbpL1EvgHncYysNVpea9krQAjm8C9/y8v2QXi/WZcnbMTAa9xR4/DnjnJ2aj
io/LbMpifRbQg15ex/ofT4Z/tIv26jRGBY0iSlpLvnjZaKHNrRcZgKuOGtsS
VBsk1TpnF39dVr5eM52E+LLIzEiry8bjm2m2deByOVJzocxvZcEZldYQ5qaX
Js5632QnR6Nm/oGGbDi1cniIBcpibr6lJNP6rt1StewVyqKHElwW3+jCRDEx
7Z96OJ/W13BczG0QR1NMoMmhLj9p8Au5sJTb1ljUylALrAocysGKTh4K38S9
SzVff33EpiUFn8WQMfVImcPuuBdObSpQV9oVLXeSAKG3InLsowRjiG567CAz
GCdOntVRF15WmqPQHxWlIgIPnqkSl60ayVEP9upuw5Eiji+2O0PgvKSRq2nN
5Fx7nX6Pm3cq2d6mk0dqrLBFDA5+HIFfIzffde2lYx5ZLcpW5sR5jeQ8mXxY
L20RPAg1JKJpL0VEFodJE0RaQU5A6kZUvJL4gUPsYwibSYn7PnEB+dcOT0oD
/yZDiKeQbMa/Hocg70Fy/3kH1PP8dnI5DN9UDdZ4gp2NQVrLuEiJQvLVyhDT
YuIrPycxuBXfBk3UsCzcyPQMY7ZrK/PUuFJv2B1O6UYJNdEU6R0A69G8VhBq
8YK4wkbGfQtDNE3WONe3g7lOJSL/bDt6xZAR105SxUszNy/NOEQEPrJqzMwp
1/bD+tcsJVWO0MxtvIbijc2HJu2laNiR2D/cvpXZ7zkmR/Xt38azzTY+cfPT
dJpQbjZUNo/9nMfw0Np+NXuglO+i5kpr7QY8mFuVZLUJgFbClweQ5ThlCKQ6
iMLGq8ntc+Mhkz3H04VmFUc//YeHFesvY2fr10uCHYfNTWruBHxZKHRyzOtZ
esN9AAbsTqvt6X5YiSAldwyNcQ0X+3yDwsxb3JAeBxbivG/nJiKHCVgr7NSa
LmHTuiQpV9GWTO4P0R3aG5DXQiY4pceRkTl0k1LNk5fZWEdU/pLU3+OSvQRk
E+W1h23DZtSttxnwslRWTcAhJDBWLx1QF8bJeYlDmqDMwsMjnU8zGsOW0vhp
w7pdTk9sU+hBhv/l+woE/2PZmF5LPopzSnqjzxOYbPvVmzxcq01dk5FMDvjO
/jy+5TVDzSOdmbMYz0XcxEOrm/7GfB4bkVgHdqKkb8fNMDW5YoGDJq+u3EwN
4/j65nCo0EDm9rabXBr7P/k12eDtELwzwqkg+EqEquDiX65TVl1sYC8yRFQN
RhYzhHzMZ29r6TkzPy233zNWKvqE+kBCVhH/uMggNCAQeQkc4Y6J8Uj94kXb
AiFCgch+dWhUu3K2wqurhq+aFdwV5ddif0bySjGBhbc2WMh7k6OAxAIJWT5k
tyfqkcuYRyabqHEpEccMJLugTfOU0eVX8yYhab0Bis9cbzrq+1+p/ZfPAXXM
8D1oIxSEClZyWgm7/xFMQMTwIEJRLjGjgGzFE/aVdFECDCeW3qonYcgK9U6Q
jyQ8U1u140bfQJaFWlfhEt6zDysZ3aWqCvv4CjEkvbuZ2Mj8OIoMkKPus13+
mtTSvq5wLXbzE1IXf+/m6AUNRXbj2FtYxd6MNVCRkWhb1IHGq5orQ32PX4Ud
+/djOEmsqP4mInehtOEqBXRnUinWM9TBreK1QoUsGlJRzz6Q9LtmalaadEWZ
99Twqe4GimrgFKBF4k8Jvuy3bIbs0+3gpjJVrm0XCvM63pijMspG5AjELBGI
33tGnfifl8Nxw9R0E/mkEqrROIxJ95Sbb3C/8vwgDKYJVcloKsn25mL2WWfq
rzi7jKv5j8xZQbjOqEkAzquKePgWUQdmiQ0qmn79RkitMyCWY7/RUBVUtIOn
5XMrBY4Ppu4BPad170U9+H+2FyBx9kUJ3fAR65U8I3MYdobfin2Drr4DOdm/
fCHPcfBMUfTr/joa2emxNZXVix4uSz6AVn4oSDlp+ymV3wki8PhMqUg8F4qF
gZd560qxjbDt4a7SEov1waOwqZmBHhLa+vEAYqfWTSfBHClYFAZU1vrI8LC/
kM3MDdJleUtEslHOa6T5/RfCnih+p0l7eWeRE2hL020L3mrr3QwzVqxPtCAy
gazmUrFEuq7VJ3d02BN6iiDphRJNvbc6fvefOCjPPY7wRFggTBr591+CVI1L
tkRVgf+0yPaBSSoiOAXII0f+SPhFLI3LTkI2vX5fZrICeVav2oQN9y+Erm9q
CgVuGNMx9oE2/vqimV/aZavggZUeA8pL2LHuMuiJdnrZdrPgC5V5z+X8qJoG
KUjpxLi27qJqRVuUCNKJ8uPlL5oDzmuGJXOdTgyb6F25xNeDUlVVH9JiP3jh
j5P0N7led8OqJzQWblMRw2ok92JEMosMF9lK7fquCjmtd8OEflk/dHv+Okmh
oEofJwg9EQ1ubSdLioawbK1Ek3kmBLD1mYE4hv5qmzfdLZ3NAtBfEm335Xpl
vf9PJ6TOWM4LtMyIOZ6MnIdaBUo7DUeoikUc+HtSHvzZhCsto/G1ezF2y515
IvvMYUfnb6VvGl89KLehqE3PXC2n+BJxdsp0VzOfVMK9LaUqzf9ggFEx3Ufl
ZNXQ5PGsOzJYMCNHYo/+s6leewZNr2zjSUcR6T6LEZ6vIeA9yNwgJfVAqn+8
9DvGktTdG27hxkLzqF2vqgSDiVaGuqibR5YaYt/5C+SZma5ykRbuJ1a+m6wU
d/aDzyd6rnYD2fJFdh5DhKHvvg2mpzYFHq5+gHZ+7RN0+ExRipTqoVdNJIib
0kuqQiryRr53oO2jw+ojZv5l6ZdLmHEMYvEki9IfGRMLvLq8oHmplifDX+BA
Y1N0LvcxGN5G3uLYkS6CNu4wxlHc3n/8dAY5bA1Qa7WHVNWsytvCyhWvsb5D
F7LCEhil5Eq0s3tJiVNkij7Gb92B6pPOgeChcNAR48vS0/VWfMT4EhuO1ur2
FcMMKXHLpHnhIeT+Lu0W1Dy02Uee4IDhc4jNehV51XMX4W4v8EaGLStsm/hF
8oz6z/a01L5NUwq1Leozlw0W3Vb/so8sFovv5P4BNdTPGuUgGl52jxYOodSq
8uZOLDe2G6N87uMrYNLMpqngFJPy9vTnvgVLtlD+bWFudr/WWHZu72xsDXzI
UPcP8sax+OvhteNs78khHoGGymnMb5Zs3aaYGdwc6VAsiRzFDPNXxyQv2dvJ
or8Y4IO+TVcoQ6vLw6ODu4XKwPclJnVYG5xyakPbSQUa+UfzyL/WQtXXNUqZ
VS7QS+9IIccy4i3l5hatblftTlOS43XxA8tcFAdKEnTDVzYTAqShaiiE4ZqR
jccLr4nSPgiISg14nO7OaWATlfdxVxncccH/M3dYAH7++BjXDXYhwje6+FRJ
xAjYZte3rNUbAZ9cZa3fzQNduHHfUuP6+czpgdypTZTeJEC5MCSb7Z57bXkX
BrGKS0TfNPc5Lx6Z3mIbpJaEdzJEcKFqBQFkyPhPq3nintDDEmalSnaAlZFG
nd8NvBd+5dQTmp5Xjsi+xjcN+CUU3YscI/dBE3MHGciVPHA+gOl0rL1uMBDq
ivZaTIvamSEjV32pVeuk5T1ohDiVurPzHGruktV1IJyxrX4e9/VfKfImNSFm
y/rbtV6n6Zw8cukUOSJqjoq236KHJm0wcTvYUOLfxNAC1jXw89nZ4VDrfH6j
bUa8alAP3SAlk//MKnU03C+VPUC4Xg+/rsLjRNtdPRwfCPrbliBMRGsEt4ZJ
ukIzNsXJQGRPhR54xj2PU05aRLYOPn3B81+t1EV6V4neZ1N7Mspo7wb61hKv
WZBlkh+QIq7njfjFo7mTTOm1Z2nBnc9Gj/5p9Z8Vh5sp3U//IMtVwSdvV+M2
u2MUnP4kqlpoPOmejNX7p9bCHh/41LVTz6Md8Cl34eQyELZVgaB5336fvFQQ
nuEy334747phhd0z8Kq0Ub1fQFBzThuPF0gNYhi6D2PKrO5t3x0QtVh8+fNY
0V8WaEq7vezQ8aabwVZcdf/SWK+Cc5Xz7DkfqxD+1lP0ebxWk3HYvXmVz1xe
4Fu+BexKsRuTyK97LjZOFjQ5dXRmFC4/wTC8iBy1MgPCTuogPOld4E6UlyqB
gOG+dWqhJghQJuu0FaSFyQYVXWACQ7cBedVuA5RzePKvEyz8L+ncOUXXzI9L
P8B7s54xIVMyZJDHMLpDyxrXHrC4Dkrq5YMH+xfyOQ5rJqESNb0CZUEADodj
5sPQQuhztN2nmQTl3g0Rss1SkLP4fWgbF/pHR1C+oL0MdIp/mL3ESUt7GUCM
jjr/6r0gAbomLmbDk4+V4i8lFeKLW5AP7YvWj+/wxek7Mc/aw4xqKqxkOQ2W
b7XRFqJbwWp/oyXy/ukPGg789Hq999bfebeikgCZX+qnuRPVxAOSiWpTSdOo
XZDfwiNYOdOTBUYz1ASlO3oxvdNQeRVl958+zSRj0o8Ubaka/GvKp3Mm4Gfj
gMBEXDGm1Mxv4eX4SWPyW4/d/ndFd+KwSF9M62XD0dl7qZSNkA7Kp+AUOBNW
Yre/GG3qk5zgFpB7gExDzq6SmudNWGuJYlBerjx8VnCdGVQDumSMDRI2R5lJ
IcaK+ge+E3Pe0Ky6p0bI6FeeMxst+zh9IlE90dLXT2SwLWE/FVBaL/eUBR7b
ToKKPrGOJCcvIARSrauw4Puko3huj4jkEhcu75sbWn/zMzWum6+Kuj01gXLS
NXY8o0n4Jcw7elWBu4Jvy+Jm6nQs4IVykrsxAdPUrQ63Iq3xSzk64j59X6ke
ClvICupM6n6gScOaradQ660/dZuXHUw/0GZyARNDsE6v7iPj2LA5cpAE54QF
ikZUlddMtge3ZvXzSJQSyjYGBCfiHchxtXDtGvCZ6DXHUsOagepejuPiEphd
UfBvKt++Hp12K8nE80lape5laf8/ihv0qLK8eXF444kXsjDCq/u0EPJWp96P
OF84oup7cz9E9oc4kSJmlkkXPsQ7EA5AqIrVfisdsxEchj1sSPGaMFccfC9j
deCo+GEbfQx1V9aWR+l5na/yvRiyGKhMYNbO4Zln7wup3AukIXp64Oiyc24k
1Pj98F2QFsb+ABeDb0fzec8nOIJXQUrl3Cm52/qnEmb+e5N7KP3ffhYe5DSm
D6OSNO7yL+Od+A54KBvrsw7kmqhZAz8z8ZmunooISwwpYFh9Ujb32S24MFwt
9gBnMYP0nTxHbMivfGO/fhIRnMrIlMMTvLx0FdD25BXEzBzsaPH4PreCK/MH
iCmlHAR2eZhweml8NXMsdTnpY+fnjHPZzxFPie49iqqxeL5btWfpVXjSRzDZ
BO8RmWodwv2E9OLmkc6i4aOcsOZB5O6qwG7u69REFquKJtaCs+zn+yZ6Iiyw
1X0ShKNkRHSZ4oaW7+teKCJk0byB1BgB/ZwabsrpZY+Vdv7WDCPblo1czTHH
tzIzOJalE1EqxLDJ6YTB02mR5sQKLjIzJRFEbTx5cYPwT3OGxsOEI3WoyfDO
GzOdwvXoCo33DGppNY3zfgppz/f+xDWU2LPFxRooE1m5+hLkP+aR9kdn66nv
f83G3yhvKJR6/Ys7OT8Kq0XP9I1p0653w4QDgnyniUvNfpXWGFNhU7traEtu
8gCIa+qAKIUFrc+0F1hAbMPJcfLUfLMLB5pzJmupqKZDWy6gUjeFT5KxUP/I
VAMjuphYk2fhIx7zmuX2eG6kg6s+tHeY7pPla29vr2AZIIC/Bt15DL/WFDNw
FyhNWwucbwqMrVxiB6d/tRpRiFqcKJAYj083cpu1dqX+d5mnxUOkHCGw3BOX
QjsCKgcCZ4aznV+u69s2icASIZfXHBm1kAkgZRdQ+nnnf2cPYsHaynlL4uqz
lTOpzBvt5sonVOmWwiC29srLkQLNzzWq3MJMyCiCukwy+tXVx1xzLfvYdxsY
A81fGa9+iy3oZSYrqlTyQfbe7hKBDCHi0++KKq4i1FPuDa2WbSbPPjw+PwBv
5Z1E5u0apbHHczecy0pHpqO8It6RVuzAOErSzmr4jrLnUrZ85sA+bTG4Eo+A
QuE/oUEFEFqUJllI9YolBEvUfgPxhwHtw647zpaTKq5VyIcWgKROANjzvl8O
QSeqY4QuVlLhS6vzIV+k7LJtiyl8UJGJf5FeTYjbSfbleRw8YRXLIhfSIbNE
yFgNPaXE7rN7aCmMqtqdm7hdXJKegg+GWGYZ+8Jytvvs/ML4nXsXL3NqNdRo
+SMjpdhKCT3nCOzZbGpiKD5YnspuvrQZXJud7gl4sDnJJKha2a3fM4a1BPS2
7r1TxztB1Iwycen5YjwCihNlltnFcn7Dske/IXU3KCUiUrdGlVvdKdFH6SU8
+ZcUeq1tTzw1UjK29wUS+NTZPkiJdnMDxlLnthU0WSXRhSDnwYXT13vSBHSu
lTc9b5GrRqI3Y6lc1w4jKPoKQu705aAMH0H4VvPWX1YdyM/VVUag41TF4GGP
OiQWK+whX6qrmYGkUupRMTU1yzT2vdrhQ/qKc/3CieTkOfe5cIXuSQbHlkPR
KtNFOvbHkEdRcunyC5NG5eb0Ui4Rs/0QXiimsrsTIhj+usyIsFAafc+/Wh6f
NzE14jJ8xNu2oNQFEm+6GU55wsDthBhQisLBXohWPfhUuABKyU8fursuqgvL
6FiONJicNPfBNPdt4DB+n1h55pIlxb8J4ms0lQXlvM9C0iWG69KB/gWzq0ft
reM2qp8CM+IzBG5NfHaZrmZvtt+mS20kiWbgqEgjxYTX1EmYR29mX+Awap1M
WE6osFccnp0ovDTx+/6wUwUWakOH86CU3rjpmJKZkGnjP/se7Ixgz0+BHsPA
wny2eyQt1xl63usoOIviTKED/CKUbCi9coXT64eBGNzyiZfwJw3D49ycq6WX
ibn9KbaWCl/aX2BNcsY88VJiAVFcXpeWLrW+8pgIsc0vFxqXXW/ijog521nd
Lnyl+CaSo+ShcP6SC0pwlaUmpTBlupJvxsT+iQBxa8cgvep0upGFs2ELrbru
xt7E8J1BaYtegIqin0/QII33DG1TgRw4DDs+GaTLMOFEHjJ0pkOpkq2e7J2w
XAoldQgRCOlTsUFoki3ZT5tvi79ActBqMq4m3gJgmJ+y9APE7i3DSuXj9JY8
jHpdYAVbInQXIzRVFa/HOL8ytiqjPvyqUkEfVnTIwH8cTJXLQ0JZ8Otu+1W6
nl8tqVooij2eIsYdggcA+vX3tpyybFiA0RgjNBABo8ntUuu9h/uxeeA/mTnb
Yu0tytGflghkuLzGb2Kpb2EfhFyIc5drwYcxuCB9csYeyZl3DQc/24qQ92Uy
bbmQ7lK/C0IKpbcudE9LjNmfC7X03TeAMA2xmo7UZHmaGcgBgg3Q0iPUgASh
ZgLfGp4smrkMKVCM0Nr/0uL9bXEaiu43LF0IDCAqDidlYn4u7IY0srdheGaC
F6ITco3CmeU1nsVsBQfAnrwTgEwOBlTIDe4RmLl+lTr2IW8G93TPtUwF6r0g
riwbje5rjypq6TfUpoOW74XNfMc3u8mKtABThpQXaDxRAWRcAlVj7rxB6NYu
9uOpCF8tOn3WoxdDW7et8lts+3iWmq0lwdP4UwdBxBlsuR/orqxuMgoDOfCy
jK3IIg6f5t+UFNQPHD4BNeL52u/QZZ5idt222Xg5JQ0PfkltS1dwXOwNvmXs
megB3ug5JCVwgLqMpSJhJAJzhsoA1DOxfgS7w7HSgScdM3i8eoX7sZkyiBEd
ctPs4jlYSvX1vTkVPg7ldjadOK5Ql/NLLkBkU57TIYuOZN5MAs6HwsWGBjhv
gSfSEBnG2i2nx0DyoelD4w2eWlzc7X65ppG9LW/FgI3CamEGDhYqBXyKVHMY
usUqDq5KD2lR35vRPNISyNyg9CMKydeUamPua67qf+kip9rEPPiLkY7R5fqp
7aAHh+3w0fqKyrDk8gbad8DK/qqWk+9MCODjdSEnYcq7cJ34dBp7oEKJt75z
/OyabBe5/Ii14NMiNik5D3irwRYdlOH3g0VrJ2CJdvul/AkuMLAO4jM2FSp3
5Oz8+r0QODLRAKkNsG0NXcsrkIjglnbgb2dxsjWqEaMTvjd23zdHya8KWedY
EwT1zQ9rRWg8DZCXdV1we2WVWUCLqp9gdnZTABoeGEtySHwDvOwVY15MM5jz
CWdDKBxPaGDUovwZDVCNc/Cu9dP+z78RVJi7+3DlNK/HkWp3v/vZ245QDtDF
duMqJ0/bHwwMwgPDpHGdP2BY0YU7gxQNPf5qh1tOtJxgW2319AgAxos4Ejbs
/+HrgsZ2/2grXaRKZobHnekLVV7dbcJD2b43kzy+NNU1D/Oi0pkYzxtys+gf
qgjOS+85YbWufhkMUKfntDChBIY22Om78Fzie8Uj/lGtpoNAeQ6Ze+epCdRd
w9LaZlcxYjWp1bgdFND/yU5YsHdD4HIT/lPQHFddO8o9JDc7LeVpQznqewRf
NwJY1yAVmj5pZkDZFhjshjqU4uC3qAKNd4P4/S2Wg+/u9dq0LUFDRr7GCWj4
N1rdSj6jhVcCNFuG4Ay78+QqBpr1m+Gh4RN53sMFfy3uKPHzdKuPq1uLItnQ
5Nz0/+eoKJT10NMjUilQorLhgKH1melDu8htdzil6GvjoNIUQDyQxMa/hlyI
l5QkxIRrpEU839dzDcK4KtFE6/sFAcuquIx5xhH+VaJmP9N9BZbDIIM1BXwj
HUHLZj9x5RTokb/IMLeoNsZ421FeUB9DrwUl4564kHlMes0VuGju8yJUt8Cx
RJT87WiI9g74Xszv5SiJfgiudGBUkRinxopRk/8kzRATbT2650LdQ78rC3cG
QP8kGNJVmaXpN/ZBmVJk2pm2ZxwROKlqvIXsbP/BGHHYNkXtKYgruDOllVZK
+RIG9o7OPPteLCkOu1uKwDNnXBM57hWhKqDakn+4/pzIP4XkTkAuh6NB7Ul6
QANVOKXMHzIylNjpcqrku0R/9erVcbXkQ0/l/MY6c+UPV579zlS3WxT6iKL/
SfETwYxUNaEXlh29HjXs72QSW8m2cWUpejgkO8qwe10rRSBOry+oVaeGJ3D2
oFCu/SF9uUrfoJwN+3W/aQdmQ9EW72e0jaseP9bpIdjosStJXY5V6fgfTD3S
PNVXQOSlH+Ns9Ox73+lQDtOzLcwbmG3T089x9CpvSoUzh54AsS9odeA+lIo9
fA2FvBLyTp9ljac33XRBEpyLVCn/KtGs5o1XxJYBYKwCaD1NCMnkH6yyu1JY
MyXR550Ey1gWNLxTZMZNb3dPL2O/i4+XaulIrhj6PiWZFBKMCl7Sh0jfsAWu
e89MTx8iTfK91DQmqm79Z9/oDXH0fdezPzr5mXpI1OCGlcawdOoC7csMCBWd
YBJhtkNNwUzgD0pJtbmYNOkCyk5R+M0BryD0ws3CpaW9L8LC9Tvt+0CWMA+A
3fgtt1mwHuzbr/5Vx3eEn05ks5GdYEqKYps1D4Ogcsg9qa74Mb5PS8YGd3Zu
S+U+KfqP3dA9WcrfSX3u+IGXshJaxSq9K3JtuU4CtD3QCWrQ26fbcJtFPwm0
NBsbEBS7zs0bowKfi2aFitYe8kIrNeKEeZBnOyCuUYSEtd/zAV6f909nrmXf
JNd5nNnbZnGglZla0aagjCJN0MTkeLAQZM7z5/H0Fy/s2ujjVnMrMrtMlrSI
Y+PJU8BKobvlOJY8+kxk2FArPhRpYNNHkdfmUxGyvC2eE676RBvYI2VGaG2R
f9s0aPkPM5KN7s3gWMMHVNPtjANbrgL1Qh+BFT2IcXJ/yZC+uSafp/rz5aHP
rsUr4opwmX5Htbw1b+Rj4NG1b20eLOuW2BcvQs8EViG1VCsNZ3K0bZ1YeGHX
4oXs9QSqh5ctnhqUWi4Q5joqK58QlNEC5ef/JZVUYhFGPBiJUaklJ1oGbd3H
VGcpq6Z+udE+S4P95F1qlZmcpGkmBw1zZ7wD/sDAIXfvwBulhYENmwLPj3Yf
7yKchQRJe99Q8hmfwe4XWD6HnaPkZwGky1KzTTY3Oc70v6SOwVJm5/EXJUxL
AzOxvL5Ax1e8OcctslzF0iYhfomtoGf/8dpVHth8IPNwMGeFW+45EhLp5h1c
PUTR97FT0/0BY/qdF/P27kN8ZPtIm+Sie34vQsk8XZz6apzkz5yilJRLWGeT
O/zR8pEkR96iaBdjBQtwBfGrs8mK8I18ORcHwh+e45jShL6G4EMycWyxbDc8
MAJFHDBkSlSyf2+bXdO71Pk74aZJC6IMKeYJrlKzBJqL+9wo2mWYXj1LM3xw
5lu4gygtTIgGKPdLt9YZPfRjYOLKStlNRmBJotjDvsYduOYNI81kwFM9X03Q
X9KRNT0xX8F0aBeI2N5vyStt19YRZwW5x4Ky7Dg5YYFgvDeAf5D6AxsdnMNj
M4ptKBvoR8dVUJBE07onmoh3B6us3cH7ABvQij+/Mg5Cl6Xeots83rrPBqsw
zuZofzoYyzkmHgcYq+OEeLlGCSRRkGfCT02nC6aXGsOcqtcboJHB/DKGBZi7
6NJ9Ym6YFIoauxCFT2UPWU8oI/yju5oV9eVWqObIx3p8ddsQO5mfKwTmJ7bP
9EZHqeSY6EjBsbAgkhF7oGzil7dCbxB1CXrrpGohsAxqjeEDbS4IK86li+68
ak7EwbPGOZVn/FbYAsCqrXdv2ZO0+dMEe6ndhGjg5J2hFAeqdOcOuN6cX651
wQYbSpRCQiIofTi0gHs2i6iicL7hJBGsLPo96q+LKC/atSmf1t4AarmkWdy1
P0D30rznuoRKRt6IaHyGH5+1LRjp1zAth8pLS6nJtuPlMh1mGzLUPcbKHd4A
HdXxXjqZN0ZOOENKdCRj7GU0A4O3RjtGU1ObtY9XA3LsjpDxFhzuWUVYofr5
bKRUS5ZNxWvVQqrowkXqms6WB6js4hgZjUmxwmwHZ74ffLIU4tweOevIQIdX
bpgAf7UFggyGn/+d9iKc50wQ0jvBict7DuWKD+GIxcvzaj3cvZmuvLEL4OS1
hKswvMFiRNNZ55VMBe7iUFy3hrmx888/iyBuZ/2VMgJV0pZmhShBzi/NJYVW
Lu8ia3AffTS/cL/JFH1+iC027G6hU6x+3P2voYo63kW3/HMeCXEJBeTjVbt5
+LUWYf8jPiuOLBBe4diDcoSCN4nGgF5eM7x8/9BjNTb+7VwodbrWZXzpq9YV
wS9ksw0W2lQhBGc2RddsiKA1mLC66QG62YvGBUXqOKP/I6TD+SBuGZprjKOF
b/ouBX9AeLogo5q1Dhd0x0VZHTtc4qVAWc8z49wvrr+jgLtyPrGOkc9jolaC
pVnhks1TM4bWhuvfoKyQFtpezS/moObU58Us0Glaf7XXKNrn0VD1dXW6J1lq
JtyVwc5UzQjQFQxzwpQDVDw+zdnA1NM51QR5ATz24WFO8IbMwQMJbWl2K90m
2z4ryMKz99AbR4byC2I381LC5XD3e35reJu/r4nM8zQwiP7l496C0baaI7Hp
HUXQWFf9p76qGKSdjVo68RVjIqj4t6fNniWJv1gmTYAQ9M+tL9xKcTTo3g6W
DmH4iamMlt52zEzkNPFxS7dAw8k4m5vaJdKyBGKd/c4kCliYvUchODSafV3z
BrNwROLnm1LMC4RCKpMNhA8YIqF3q2voAHLqzbEP6A6MtymvtQn0nknADw4j
7CI8e6SPdEUdSMHp+vl5izVaCloolitvh0OLrZYdP6gjKFKMajbIxx4afMRA
vkrCwaZ6EYDlsbFlSqvSKhPoA2lADIXuBycHfzw3NRrjLrkOrNj6B6nXb9Tp
EtEhPAlPN/fO1s9HrQ4KrHan6Bf8uigVKgiEgF8xZwarL9nYhxt4UwRm2LsT
/d9HKyZ4s+/zLgCiHrnpJUMnGWDN6jaS+bixCMUNCIFFvcDsQTDn5SRGIa/y
0rnSr+KDPUJdjEdVN7RAOujm+USMalXlJW3LuTpOwmY2XQvEYm72Yftzxr7c
CGyn7F7x6fuwYb/u2vEsRA+gIzSDlez/iynz8e5jbxCQQ44fiWQQuRqfGviz
6MWBXJkVlL2yVx9o+oI/HIGdWqkTyeRigz8u/RGfA57E51lB1rF1VkHOLD5g
5iKpR8kJ+gHSBn09L4kPeT+xMGwu5cdFwOUQjCA7Cdw9lxzDLyl16EzXXdGG
x7/yLLvBY4u+3YaRvoCEciyOHminpZAmIvi8djsEv4/4V4Lic5ul5aswmjI3
t7K/Dtk+13bKvqCJFJyT1hOS6gQegykMTZfGvirawK/r2mI96FhCB/tgdcSY
ImSHSz3vToBKO7GTsUaInaR58Ffvf/CHw8qJut96PyApzkcmw8vi/9oULiTn
NskdU9DgzG3wZVwapS+QaL2+/dAKSvbQSdVnyfN5jnkAyewZ6UdHTvOrZAzE
ThoNsgEGnZmiojHpF0ksd0TTM9SA0jQYQtxEFpHjnWPe12lO21jBdvBhvPu0
Cx9KqJUIbB0NO0sN44grc30axzYSwBgyHr/owH5SfIWUVdXet+P1t78M/dm6
e8sWqzl5K1t08Qrk+Teywh2iLgFptjN3dNHwRQ7eFj799SozIlBvnoHYibi1
0G+GaMO9wd9cDZ0f2NK+glPRuUyU3I++dW4PaKMK43koc2fASYjqNh/4IgGK
fy5jY2VHdH0rcZcXCI/g5sHHb+Gku+Y4IOk66JtHRIP+xP7KXzGEWZMKWhmG
XAeiJ7rO7pUG+Q6Q3Jkyl21Ath6BIi011KYLxkvAfy2gW6ENLV9e9c4ExRdw
P1I8zWdUPfa+uBFEM5xxp/o7zn0UKSLGNEKveMFxSrkqQYflAnXB4VfHX8n7
Swj+0bBm1rHWk8JhOdmY65gp8SPE+zS1RH8Y8htgjwX5OwqdABZwnl4DNaB6
HZOFVMvYXnYJNYDISclBi+0w/GQXO3Xg2mVkyrYK9QTSIORhJejzDBd8iC+z
LBv/keVQNorzoTOU5N71E+H7NZHX0kB82Qz0D4sfhZlnvOFKobDlKVUdkv0U
UXBNIPOqzf2QQmZyd5tFmzopmj69eUYKa4d/bDGRVtx98kyVJkMTWIkikRtQ
+Sm386IIiUFlNWlDcC+MzhwZKxNssP0JkzVrpQWF3ExR5se8Nxz1ZI2NCc8E
9bt84PfWH//w/goSbgY1TfoXFRiy1NJcah7pWA+YgiNZXs+SSz3D5yQ0gDF2
WOYeadwRNqKXvjCCRN3MczCXycjXTZKl1SDeqnk/kaYuPMqQHvHElQnPMXh5
xlKuI7wbXICggFZQ6wn81GbEAispO7N3lcWyyUaD9rTySt+xF6rOvtOaMrET
Lr9Hu4fHus03Gy61KTrvLjCHlLTUSwQvGqfhg49fdRQ8To1m0CtgAthIs4eO
iDqTmpbd4h0MtQoR8MlsHDECzHOF1Sw5LIR0ownNpSFNgAqCgPdUFYUw7gcQ
TKB/dQJkNnPIz8WQ7s3mRUJSTSS099qTy9exFvdBtfHVxSln0ivCuVb/qO8t
bjlmkoRwJ/oh4lvutrTLwk/3XFEE1EGIKfJoRq6pVx+TToZZS/SZHw37ivsi
9Us8AiZZM4Xel+3uaHpCCtQ9BxCq+5/4tD2TjbRp7wXfLGmaSC394eLxND3z
+9SErH+U2uwQLa2BHOHTPTkXvuWWpwD2LGBcQpknq/lap3aqx3J+CR4dzBsk
t0FUMyJor39ujuOyOBZXxiI1JLXEhUZt6549d8JmGJeLgnclaiZNjK2JHyWm
FYvxugX74HYJLm38r1j2eumQNdmSb6UfWMkKtfG5tbCBx8mqJm+8CjZ2gPCk
/paeapWGh8A5MiYlfORjZZQbQ0eS/1SSM9/JCarEhm/UoJfmi/16DDH7NeOf
iASN4qBuMMLur3o8TGXXvkNRXsX6E1Toly+88UOkhzC5aBNUxdvCcNI/4T/0
oKHOLWoXkroxhZY3HdxH47vqhNG+099emDY11YxHBWEuBd0XN+JAOnYXQYqK
F5KkRC6RBdynl5QJf7ReBunHBVpcePrNvT2BbYgBZ9dlGt9czewmW8lvD6Ua
1EIN5ClosmIr1iYgWinmj/zHGQzhXK+2KxCMK1mSfOC8l+kx++/oERJKvYrg
irH8u4PZkRR0zIS+ClbELpdJghd4vWU4GacJi3wjK+Fm16N8D9nyRo3NLf+D
xovzvu39BGsQKxLRGAofPgDY4Xabym4CkoappoGrNvEgYu9+PTYxNqLGfMWv
OBBDzxadd8Yet48fWvj0Ctqptse0NriX88CuzTP5sY8DlrKLrdFoFO4ifxdZ
LmXeO9bvC0JC4/kZJVPFc4i0gRnY04I06RkvjkVKtOdGiyYwIugDwnEE0cd3
kJIA5ebAFQ7Vo2Edgs6lzBG+nG5dmn1udyXbS+EMiL48qcsqgQq2ORZ+SGid
u/mlHjEbhJx4VQ/rNIKTr4Jgo81+mADgOGXZ8w/jIuEPAIGIf0SSP3oNOwt4
CDCuXIirHX99/jEHxX5IhtM8mkFIvF8d/rQBOXU54zVTczKnrZ7ecskXIFdb
ZGTqsk12lvoNwHZNC1qdrwa/pCR0JyxeprHitmEpyVukvGjnnw5W+hrniN2D
/wp9X8Z2HTPyJEXpBx01MzKSdx1BiXfxHhkRNidtis591h8EA6wH50/cjmol
xGRzGCiVl4LFE7pL9N3rGFbm8E4n16kbAYTnKn19CF8AKIH8ae1Z8OX+QSWB
CmyaEO1m4vNantkf9NAdlvCJpM8Yy/S88Y1cra0Hl4sbkoD9v0qVFVbf4Kvw
tcDi24jYD7S+Nb4j3KfJw8tpNQ88zklugxfi+h9b75jh2E+3jAQnPfaL59Y2
ov3lo9j4Qz8lWOLg0LR0cwFFiuFdk1ZTtCJtnZceYouHqyPAAqHyraG4xKwa
pn5S0Cm4Iz/ztG2TrsVguNuOIM0tTwVZqvc/Iu7kx5DkodShJ0/XYLo5T0cF
4rvjA1xENKW0JfiBVoutFk8ZgTnr1JQgiHrvNCRQ4zj2BIdfetZFzyVzzWIw
JUdsdNXTabEj4GfFe1Wp1mTIYC4BJ8xEVtFnyDUJ/JJxMrQqTiGRKJN03JZd
5KWi9HNOo11nj3sNuNek2u4RowrBj5g1p0ygahv+Omyfdpj4Ep78rFXTnuj4
iP3siw+fvpA9KmnFUVpJYE8gHo9YPw+efcbV0LJr/sv4YWV4RHNa4ggSlhft
71kKdk3muJUSSW9Sk/9BTpm1LcXWpdmeuVLquAtoVo5+99qtPrk1HWUepqoW
OKHomP0r6Hry1yB+ihvzoTnC+qvLirP3zl4fz3GftvejQHhH6Lqsx0rtIq+w
1PlOgITvjipYpsY1ym8krSYKfNVxn77FcV9eqHL2VpidjAZBMFcyR7lK44/m
gOZ/pJuHFv+bJoBH7WTY+s3d8Rpae/HEpVt3lxOu0jhd7X6tvUAsV1N4rZjp
2F9lkZdqtbzH8DF73Cm50QUcPPEOQQNNNNEMYovsc89WxbCVtNxsSux5bRAz
4FgO7IEZ/7DqegYhNm5cDXHTKLua3cDz1i3wUEsV9VICSQM85V3hRUjRnYYs
sxE8KAVUkWSXZ6fw6TKOx1vfUV92HP7KKqYlsvf6Vvx05G8IihV7xoDTgt4/
j3OVUhiZz7ZF2ZToYi+s1xWBak558QYIaOB4oaYrpaV3FTPwLBUnXCXrcJH7
KL+pgMuJZ4/ljlbXVySamxwkxXiqtkH57hIE71BiOjFg7sVSQpJhIjZeYLMu
buL534CXAwNwMC6zkhvDsJON7vCOzL67j93788w1MxvZ7NFr87tqiICbM9Kk
AfHOJHQINn+I2CLETkT321mZhpmJ8W++gUwXsLFVIdFPj+QvDthSBvgiphID
60ga+W3bi612wuHvidq5oEknzwkzCECjSb5GsmX0p5uUzJ90qxfXC7QTAMeE
x221LREtMa6reAICJ3twkLat0aJx/14NNTJ+8ZZOR7cJn5oj46SCa5KuD8pO
B3EX3vY+briB3zYRDzXYALlYwhKb5718jO5leORyHxQYDTIwZW44edvQTWQS
rYwoPM9prYg9saftZkqbR6TqCq/4jrlDnMuDQDUbzlAZwMHvI0Y4R1uVqWbk
ZYP96fpm2w8QrxVpFfWpl+9E6IjQ/FP1VUkthzPtFqQKykVIuiW1D/G85hYx
c4X+/GfWiSKeLFSZ+avP/OzQ+oTxfzT1G5z5/ptuM94jX3K/+ujyu5rvuhNL
t+E4uIGkzZ6whVYUdzTPtdtIZ8bEUc2ijAV1rEYpxVOcXe3Qgph39wW3VUWx
y90fqEkZbW/ADYjPlao5yUAYPIqNLmfplthIf11byPtJ3zP1BNmDtS8SRJG3
pxAa3Thp3+3LD+N/PgR0X+M6o56OznGJ1ChiDviumnKti2k+Sj8Vne4qygs/
wazpZh2z/37YloMa1W/g6uz3WHO0qvh3UTucXEJ/pER3wU1q5TUpooFTvw5z
5khL/sNyKIEBp3LBrZB3YtGke0LmMOfypC7VS9XwDx7UEx2tQbxRiRab7dbe
1arAqa5SlPvZ5Y/934ioiNOtyOBT03f4CjPt7FI66VpQgZO2ezYl1MxqLN1s
vq6Aim2gYcMu6yxpzaK7sSgx3+kUGqKeFOkYnvBEn6hamGkzoRABhvbO1EXg
5gcuwGGCYBIBI3fjNrk5KJzef05EgRTowv12APWi15LMkbkQbHFeuQz2QoPo
HvZYmDzQN3WTv+QXMvGN+zQlNnlugEc6csa+3XTR/8kVzeKYRUyS6qPukrWi
ZbX+JoTxPURnk+s43QVHwXHM9MrP0bH2tzWykOTelAUiTPJvnkOjz6Kx+ffi
wyFqI6UuYcbxfVFIhz17LuAE8jiu3NsSSZxDIfmq0MAG/1BT+T2E9uwIOiGP
/wYymrDznJPvYap2Q5yZR+e+MGArrJfniB26LJY2aziWkUGSKt8zkVn7gJYQ
9w0o4j/F1EIJHLubByZcQY4XWQTyl1IaZcgsIEaBxNg6VRK6pgIWEqbIQPbC
MuYu3Uzq2g+jlXnA0bCTZ+0t/naHHCg1FFIHwrXKvYo0x5M7mdVJ/nFZn2ou
WS/dSviqqW/RZIWrQS2M+2eddO0DQYvcIYVgxfz3g5GCfqLo36rhzYcMqZ5t
y4uNBuHChBvh7Deg9ah21d9eOBGljnHBtJP38wXwn0FNUyU2ZOfST5nTULSp
lQ4stdtvfXM1vfC0oG/+ILxGiQI3LAB7dywN7ycKbim6pyHsim//GhXRiwkB
O6rlhQEdGpGKbYEFTAN6d9+wGIGf/nZbJkWoo2DsLR5nQ8hPSQu/x34VQW3f
BrBtF0hSXCwraX4ivHWdaQsyNTXT3rJ0N/Oa5Wqe2eQ/cWlOkIIipigaFkfH
8nyHS1+sszru2eVbcGu6jEyB9kwAuqGFMhSBhpagVYeq3ahRdgvMD27WfdGf
8NDreaPdUqNtRYdnkkHZY0Gzf/EFQivX6cnoVW4ZWFwOjNEtRbSQK41uRthI
Juf2LnNMzowRgjpC3jX0aSrELNlRBqmTFL52OjqY4SNsC1kQEXL89YWvJfCJ
MdS7T7v6uHcWo28E9SrCsantmDkgsZcPWWXrGSIsvLTUsFhaNjYgsxWoIVxA
WHuHRz9XYlhpPoHI1h8Hq/mRxsrE4HCIPVgUYJWZthT393fHHmp6PREdJ9Tl
4oDdiUkfv8Y0QcJMmTmqzyS+fQAw6BdHBPtsyblaDcYyItcmIgE6oOyzob/w
5W7DkqTzWJ4mr7MZznf8u5a9q31C9+YuUeZIoEpzxDtg//FbCCTA8mnj2gOF
BBpfy+B5Q18Ff7wfLcgcHRn0lzh7eSTi78N4z8EDWtaV3ymDEFfW1s26lmT+
rbnPRzZ8CbLWjrI9cf1CDYaf9TjoA5iizWwGeHISwZ4sCOfm0ksZfGWxAZm+
KRCMcrm8Jr5EkF7y1+liq3QEr2tNTpzPYM50YH34uiEeYWqAymr56/CFO6fr
ChNm9ooHMd28n8MaY8+F0LuNP0iPt9upOPwjyoYU1enHlJ76Qxx/tGWB5wv0
SI+ZlaqsYWB+dXYs1KvPD+zDwRZzHIF73z8/lh2g4ocA53kirLdlrtQbC5Ji
i/5EU3O2lTB1XblCioNIxL39W6A1U+ibnKTdLeBhR0+Kjack0fLpuAXc+j2I
/nQO1r4mHtmszwZnI17eS45bRXbfXWBH3C93Cj5M/7GyWveYbF4kS4MSOEwE
DHFpgys8y8ln0VOvN7rNq2h6nBmT68gfTFR4TXCyXrYb3ePBJyNmfOKhbSzb
YFHoX8uRAJvISUPV8yI14ruJOW7719RbgITxPJmaXgi0TCDwSABt+ROCgs8u
i8Y7rlaEv6kvD0JAxrxeWv9hXD4vicEfgxOymzJgkJvlxPZvDvOY7W2xncPW
UzCab2830ZXr4fJRt0PR9JJYqs51fqSmsfXsWWX+xzRRWQoM3J6Pr6NlMAUr
c80Ethr6e789hjyppmSmz8tAIKPb7G9eWSMHNAhWkU03eHf5IXEQYAZ6eeXY
eKMptnhBa6ja2RJOyJkwM9Ik//HhYy08cIJHA7+4hTzthfPk5TKR0qfAiULZ
0vv2dcIN9G3g9iy97ywHf8mGRzjjQ3QJiX2ay49O9gNA0uVVR2KkssiEvIQz
6CINwEY+56Dp52fnR7nLgppg08X2NxNJrTLAkBGoZ4BzR6JqnTOWqzubp4aT
LxUIVYLTP8QRj1eNiDOmhnbnPWuVcSwKT8lVZiTY2gWtYlSr2R8aaz55tJ3D
0yyLL8g/gVP2QIcaUxmZ2Veez/UAKGmkwDfXdOGEBbMaFMPPixWCshzYnHDk
PI2NWEkGe6uPIrASBSME442LSISmWP+h4PAwYodZlP37t1fyrnmrxvy2JnwR
E98GDNJU89319o6BnO1kFIetrqCTgvQCAgLQf612qBRTlhyxqeeGvH9BBafF
SSPdduowtbxwuKQssWQelg3F5Jqeh3AoEpQuxSPYJF+Z9vE6v9SZFF5esFhT
Halc6rjmDedwIEwQw8MpqVzLxEQmICbiEpfEP2EsU7vivkXx0YnwfgugRcPE
a4xLOV/klxyRSnGEeettGN1oZT574hh5qS8YcXyufjzYTL6vCX8hIIHmfw6g
NgsznytjMD790EL79QDrYPn/X1FA45eikvAYa1GuJjPadAs6Nd3XlaI6CLr0
RFtK0VFVRzmVNztQuI4Nim3Qoh2/9VLUAPuEIOFedqHtjLDCBW6OOM9sL59s
ybok6Vj1L9Mu7/2DAaW7rY9LRTie1xf2DG+aEe1a7Q+G+UEQqwu+/Qrh4YBd
FnJTQcqG/4JpXpU2SERXdapun2a3lzjcZz1xCnW/D39TbGml5AsoA1PFB5Ba
SmqkBht0LJ4LH4+xTCNISUqhzWb70XZhYE67HCx4IygY9TK4Dohs40znEnlF
CZRC2/hcX5SPkCcgWNYSmyqzfqKmMOFNSvY3aqnVi8tK73ooV/ezSUT/gJbj
kCi9QQLYn5+BGA0Mi+VmdRk68tw1WjrYbloVtFk/PvqHEyrl03y+9BVj5zUx
ZLYz4i4R7CeYL3FjaAxXk0nLLWwAmB1gxfHJBn5lCLoyyV5PqeunRUrtZbSw
wl+zp9qQdSTXL5bnbw9VOnfOvdkeXvMjueCcPeiPBd+83oTRRRxN2uXndL23
cbBpKBmE0T4FQjBfMHDasdKGK3q5fpufklai4NcNwt9VtN2VE/aiJVoD4yqT
1rm7s6VUqcoqXVnRDt4welYd8QFUU+Z7nB/YWqvKxaPRdSGUVQoJ8g4VQs/1
yrqni5pvOoe/3YN/Ua2DQq2lKpFbuYmRgMEMit6/qUBJUfo5TguHHKFZ8nyS
35qBFP8IquikYFth7+fB/enqR9KBYvhDapMSld6O4dvmswsQYIVatI6Z7QXL
RAgSllpgnYSgTE5EBIC4Xu6Qrp9U6ib+ozcTb0BoAtqRQWorJ6obpPhC3OHt
WJxhiDQFRlJOJYCZbTtnOUXkFKtAmQwa5p2Q9chbptHfzfnzEgQto1UR8yYH
S7XoRYUoakzfdaB1hWOBlzbUhRhdaEXEjR1GzDzYuRFnhpPN25oAd3MU/Xlq
o65LD7zBFW8VFEg/dvvBOtKllrG53TYQVNPds1OowHp6/y0MZ5pFlHyX8vJP
F3UvJVLAfzCZ01TfkqCbAVlssQTbw/2AoT1Swxpo6Ztz+1aCoSjLLi42xvuy
u5lJMiHZasCQnYka2D2A4AhNzZU9cm8pY4nK53qcxPgxdSsbJ93CTwZZehbZ
npw4Q2Ia/O1jpMhL3uKEyNuZwOSAtmrKgvmDLYbL07VW22scod3O2ZvjwlNl
m9cxjPxQokCSmPmJUYU1sWckFzJqFOTv8D5ut7se9VLI3CGoOu0FDnCJefW8
N2uK1ingg7kyAS1Ls60JlyPonkl/QSQtPZPDgy+hOpOsNjiLHassmbK82Oqu
QXPDTkKFHCPhJrDmDLkNP76ULbFIcEePiC1OpZyKak0qx4ajLoE/QljcxBfK
OmStRtoeUTPk6Nk62bJxFLnc/CbCpSesQV63otJ0/4pw4wialu9vdZE3MxlY
LWv0Va+0n0JLzckaylK6DKbOh2IR0o4fi9PLxuZM1OHPqqreFLiEedBapnP2
EIHQCS5z97Oy4FJ6JCQB2kXoIxdh1kJXRcIG8rYxlirfkoyOiKsTny0u/rba
RhJn/tmpoTR5nEWtn+dXcQxFr6nEAg+jG60syFWhEl/lUQKcNsgK+DUXa8tC
g24Ccuu6W9V98U3Y5xA0sb2Tfpezru0dhz48GRUt1XFiGDhjjHvePR18Txly
TJb00IlzgscBJ+Ux1Spw8yuBLzhhvYFCIYJBeaxEwrbkzKtODxyOLCOm/RNk
cl1nHqoqGLNo4WIYaUWrEjm0UtFTEGIzc5dSlH5vrj+ZuOpoDiw+BfXgMfDz
LiV3Ya4b+XxkErRXKTcbmxtFQ8UclATeqXxQVe6jhfaGIAIJ4jgaKcA9YcrC
PL6qyRV6eJhHPqMzzRka+3z2nDP9kvwPtQ564PURnQG2CnWzYiUj2uVWkiM9
rSriDG5V7uE5F7wk74D1Z+axE3MfC0lpOYAHPGE6T6cQG4SC+EMRcCT6a8le
Eeu170OWdhjclV1QsvhGENhTW24z2weLNzGJgxqMIEuGDW5rfc/Xaay2QeUl
mRq+RpN60F959iBZSjkTC9npVohiSAlHqffjffy8cQHkPhKOZSJTuqu1/x0I
oc0vqSlW4GP/LCCOIOkLxntho15VyrxN+MkgaWwYXm/ygkjghDB40k2owRE2
ObSxTfNYr1RgwV9phy4ri2ph5aX8UhsjTub5dQ9QR7+TQngDPa7OwnW9ckz3
2Qdznvy1fw/yQK1rVUxensoWlt3x2kkg+D0HOWNzs6bbGSfNcfwbn5Tr2Dld
VDHU+UyuOBDchN6i0gb8oJo6vZouShq+VCdsBF55Yk7JFW0j+9GcPGF/jrC7
vrdZ2cZeW5/McXGKvIGMkAHFLvI41/wg71fm+g7lLMSrFvz1zGMFN/VXSf9x
SwfeTHOBjc3eh0SnorgFsaIF1RwXlGiNqGwU4NEu7hR2BuI3XOrlcQQlJ3Xn
jETCyhxj8oC1Z7owVTD83X4xBDxj1Xea5Z7pUWrWGXXCzEy7w4eUSbzsLgrB
g+yHV6jSY9cgH0h0gFLI225ZuTgsoRz2T+bsPFivJrl/dou3jPsULaxe+X1a
lZnJrAyq05Secg/o9Gf/BD7b2Co700+1IfiPVIoiaiwmpjvrXmgtLSBmmIts
8GbwOgP++XzMOzxRiI2FSjykc1nVh9GM+djSWP2GR27MiaeehhrvpNao/99j
CGj8eC9Qt/DqTFeIjeSfwceOXGYrhEt3sszcEKVzhXyubaEFRPB+KFT0L3mc
wBvIkGrI4iai+l75qy0jEt6mBTxMOPOsIJKP+mmMl29fXkMaTlq/eh40cA6g
d4AMRtouUWVbtngSLX8B14Wti3QGuVMVPKWugkU9674WbQt7UN46Z23BxT65
X1Smbk0yFF9uX16nOcu4lRw39PN1vM0eiEOZPY15YQiiRC26A6GNUkv5ILh8
L7L+7DtZSk84UYSXHazeh5Wok4RlDCA8XEk4dzYkbE5pELYPTOKpmnZWfr5Y
oQCAUAkQdB4W0l9UuDjo03tDirOSpMcEfHcDwhkr8GmXo4BkjSM8xKdLsEUJ
7Juu4gOIbQ07JQ6izRZSHdtgKrR7QER4jjN/NwfFjEgcsQgJ47mBMDIDvKRw
NioODiItNlRacAjWmhMCFbJqvZEfoGnytqqvs5GPx79Syp/XEqF3ePmQWTD8
froQLB5n+OzcEMz8jmS6c7+2ywuezBjA9xaA8Q4BK9q/d1+MrOu/7YhNlkN0
MuRJqd/GIuUsvLuU0nO28l1Ot3ygo29ZWtS5AOrKWHNAA+jP4MuKvbduPB5v
snsc1H02YsYurebg9G2nVcqeYF2a0gh9GnSP6n0D/A6dhpCBv03b3JVnu1k9
eofRrxfPyOzmMIU5DT3eqmJwI7xQcNxNa7GHbGaJ6aNI5ps3DmCz6w94lNAc
d04Q1Lvp10CF74H5YZzI8IWIRSZO1uKR7LcWDCucFJFAT5ThSMQiydrxi5cM
09Tq8t9gurDOMLZGWN/goQ1RW4R58+Mlhu4Iy5RsG8+tuSsRdFXvLDEjTNF8
0mF8SXqzJ2830goaYMyrwf13/qk+N6RGEyKw+6FNwT0JXUEycMN0mW7ewEUK
PxnSe6kGtGEvRw6N6IqF2kKFQzWRqq3A1nec7nYy1Jrcb33ArwJm2W4/YpV+
q5zT8oyHgQSpBcUPYLdFIQ+mWDRcRO/ZqShSh0zZxwT5EFOMjshxg9zEuA6S
HI4MzEHOWklvcRyJczs1xHvT7roPmL0fzvWSJ/aLdpNxL7pVHF8CH1h9UY3t
N46paVLvP2kDUmep9L2PkfnX3HdWvHGDeQXhxlTB9ZlUSPIRzJCyvlN/9fNE
TreRyfcZDrGQew0WBQZCNNyNZ8tI7VBIBe9pSv+wNFCFZ83bxz7PgKimMifJ
jFIkl/4oIrrr2dgPZYqqmV7Hl/2/asXcZTXczx0YOmwOXUOiKQQna99q5SRh
gzKxH5D04bAy0613HAJxYuLFznfkU2JK0SJcp1nXMTspBe0S/iZlK4l33rr/
CPFdFMvluLSFY8RGsNRlKW54y9SlMFVQZpSAWaWGqa4ihQ5EqR0Ya3pHF5g1
mqaD1dmc1KmHbZ9r1urAah7+S5Sv4F8l0hiYbheLP5qsyGPlrg4QqdbGky58
VNfbeH4anL2wT0SnEZolXi3qeAv+puWWrDwzbX5yR4uPvVqKdC8vx67Kbm/a
JxLSMLGldqxJeHiGH/xrpgShCYlI0ts2tz8zwtDNDnZIAhh3/jOdWLk1zPD2
yRYv4DxTGOakN5U5un6a3tPhgGt/cn9DLzSVQiN2u5YZdj3VrAmGtRI1j/qa
8m1iZGvobsmoKIo1qp1E0IK5C4NS2+w2SErkUGIVaX1a6HRpcGYXWXBq8Cn/
XYhxe0zjc0HSQAW9AIQE+4c1AErru+/p42psY10+MFi/kXqXHa3KSk8Frt6H
/8Q4XnYFhipTP++bDkPkiOORSWdxaBBkAcDmkAfeAuAdb2ejJtRRAjki59MO
MfyEVoznyhnujyNMl3mjWwAGgVA6p3LI93BC6TiGRgX4dKJYdk/8uG805GDf
1yOsAIjn/V1NTw2CVR9UNVXdGic+VsdYvyLWbJbqf9ypi6YWOKB+2AIAN6MJ
9ne8xB8+3OsCUvkx4PKLD9tOaDVfeu0cnpfQlPtgDP04SB7WkyCkrZKiPky6
h4ot5snVUMPKHQOcJ3jpi6766tiFlfBfY5UX9h2lwvY7ePihGZT5G7oXg4jb
lRXiFDPGxw/htrPteMcwRIwMz6ER6oSsHsSvDtqmrrlUH4Zx+zf+rEhZVPFV
L2g7eZb7RsQmnUbjX3Y08GriK+nuPefcq1lO9LW9EQh9BlyoSkuIkig8fdGj
tTu17JfyQZqq/M0y0LPNDyMQAMsUMBHI3eP5yTAMZ7xcj4aL03YCfSN4eQ1E
teQt+lQRmywKI2Opq4rI5u30igo8L56AgccHpKOv+FB2Niix1p5+V49OXhmx
Q13//YOvL3B3SljVPyjW6bfZ8Wwf4WNW2EC4roGa2wGSMHDDMz4rBGKFBJTj
YI0Z4EApmOBymWSd8Hmq5CbrKN8BEoBZt6E93aSCYizYvKbHF4a7x2n7EwJC
UiJsyKM/OYLDZiw31UbBRjjiXJGTZigbWhDPSeqRY9JT2gTmGD1RdzZTNXCP
keBDx+T/Bj5BUtqIU3+DE1C8aX4mxgkVGGl/kZ4SrnICwvOfvaRR9uueVRfq
f8MwNG68VwPLnSi+G33Renhrqp1fkeUnouguiuf36XhrzC1H2cyWQKzNADmm
f2MxTreknjh8/JZh5fSFArWHc46T0WNv0f3O68rUlEMI8f+YNhki0W6n0L5p
sTFw3Yoi7Fx2WInsmFqNgkknvPF9u1EEKv1QJ+FkGqcwBwC4btk9Jn0aHMz/
St7PG4FbvSPrh5uZDqtOs1OWOiGLzjHXdhcpV8DAR3cYD0Lz+beocmkmZocj
0FSHcZ6hFlsCICFHOEo7jIpL8gpw0gIsmFmxB6oL7yZFSokeETjYCBu4Rt4P
lbRlWFg4vJ2kH5+8eF58n3JWkG4X6/19Nj/FTEQC3Nn3kTg3gxtT/TYhiBBm
lXDdlx24p1pVkiWgHaUOK2jIRAqUIY8hP0qspbCSQb5udSWyp+fdxOoJs6ir
3TMP0CA1tm5H9X9RVxg7FpwnrtHhmtGYS+qdM+vKsIYcMwTQojYTcKPMgTJ7
tt2DdywbVF/vdFdTZrCRWRCCjEl99h52RfOuTFGQltuNFhnKTXmTutUGeHlM
iSKOsB+NG0pTlc0u8VlKq495Edz+0OHKSG0q3oygmymGRV/VtcE5aC3KWUJS
INcjqhrmzvqevTeW47MR1vN7nUDANm0knLNzG0j3gSYg/Dba+2gyQ598Efq2
krzGc7q/u8qOOfGqYrBMnNwJG2cW3HuXZGB84EhYRCajbK/RHb5YFcqP0cLt
P6JcfX9Mr/Zr3TO1ZFylj+RXG5q8bse/TZJPD/kX1k62UZA4bEOluTj0NgTh
+Dqq1DlN5C48x3EO+vYEBX2qGjB/zDbyXH/oEi9HAL/n31huAr9Yobmw2Wu4
up/mqcpZob1DfhxwxVHCU41Bz2DUx/1+RPFRQsXM1ToHvQGvBNYHegK0wgiD
Fkon0Yct6vcgQ+L24p1QkKlCLN+Jqss0l+pDltH5rs1n5rItBZd2rMRdSu1S
E4oVAxg0inYxtOKI5IHAvJlS9/blX8xXj8o6whmKjNAbZ5hJL+sR51ADA9JD
pgGd6A0q3pSW9yDtclU8hMbdM8pYLC76hVkpuDgXJgdY9yuHznpy8cBRGJTX
GCMMRpumv0IOtBXOxPli00jV7VWfPJFszWEAKZebr9CedvMnN8wFFygXCK3+
vhYtEv2jzRKbkbGrFA30AfwrSy5IkMIJxHnVBbn3UZdGPz/cHv2mjbztYx9n
hWEA0r1mcOnrtVhJtq/DsPyYqluR9fTPHIPEK5DcDtVhE3GPZvZFP+YrFwbz
pF5e/FWU8ofOiyr1u5LNg1R384ga7W7Xm60NVFFEfBzQg0PefllmFzn+ZbZg
NTqoWJ8ZZC9JxBWEGugwoG6xPpohqHW2dw0/usD0MeKy5/z7Atmut+YANxxK
Og879JQsTnc055mNCWSwEiNYK4ADgvrxBSgVMw6j8ViF04tMAplwIWiV5yas
IJT5/HmLohID5mSeU93GQ7/eg6QNB8WkA4l01ROqbe6+qka8IZkX7Oz6ZQu9
bZhXwRCWoThJL2EwtXp2N+cjCxtuy5emdS2dT/6s7CAg4cMXRXNfvVIf30cG
MdwiOh2X2kstBDzLJ3v5eXWB6FY0N3wXBpFI+P50H7PIEDx7vMGlgu9R/rd9
dxOWuQJQRE2Y59VI8lubUSD8ZgEmyBJ8OyCVikyHuqbUaVaoeflXYgvStlf+
bCi3RrEXhGAU9MzGbTyokiFtoLijzxeO8XrnxEZK4lSaCEJlexSdXgN+EGqc
JkEgPc3NMW4wF7BPsWumXxLwo8//54z6W/yeoyq+8t/5sHQoLAWAO/FUBrl8
B2nD2GtElhsa5YKHl2f8NMLxRY7X3rTcjo5ICn1zG/Fyr22iYmkC3hqiUrbJ
F9Ng3gFSzRdtCInDdRL8CY2atIYbHzQ0lcnv9lbhGQdojD1lUPH//N0vkhtP
J8Ol1L2pHsXMtV4aLUhYtsQtXDhGvw3xb4kSqW9bhDuXxgLWVDp+W402RqZz
K57FjFDQS1lh+MK6vVfhMcR0EOEcCjp0GOLb/L2/g8B26verZTrDGt/N+1DZ
ila+8VpugQAoCY+Wo2T6vaitZWXKDb6TbuzwQdDvDik7pIMLwR5Nc+UGeGjb
Q482WmhCN3NJYN38Dm0cwUiaiijgOsmYBx28KMQz/McPXwlx7XAh/jEbJ2e9
CvExmLShctm3eHKgix1gNVmAkcgCL5kHoLCrlpHZJM3HsUE/nSuRzynxV68W
O+ue/6MjMVm+WSTRdu+93M9/mpxg4H7QoLCt27+p/C5zGs0jqncufoQVZxnS
XD8TcVbSC7d7jhJvdTvCOOS93BIex6JGf0woC55rBlviPdH9Zs0Uy5EUk2Zz
ohL8MeMA6hAbwUvXIY0lfgG1QRMgBtwqZo09hHz0OELJmsThACk68bKuIEop
xngZuq9yolmm0MXjTVAro0nyPcBR8IKPct0Y9v1b4+ObytEcApdNPxS7dhtC
QmxiVT8S6nWtZqz8gP2tH0UWbrWuAf/6/ul+MDLTbx8ybQVs7Gwm5QJsyusU
GUHdCUrNagcDWEvg+VoBHV1sX21/4Dcss7BsquWUB7iZlKKZeF7Jxpjjwsk8
XhAfYYos1eEluDHHX+tqwwK60IOaPBF/Q6ZMeufJQBNJlvA6pZPHSzxZ20HE
3M4tK0dtSTG84Gx5Xhu9fnB997OoKUukZ7CLBCdcVXqrVIpahSRuT1KtxpdU
ZP1azxhMoEQX1zzktNgSoPzaz5JakXjio4BVHayUjafEIvAK5H2X/71Y4Pj/
Sxt1dh3qRj1EC6paYCMWrPFQKLOuEW8TlfVxToFNx5Y2pGvgrp2N3tfEHEcg
QqxRIhT0dbFEoXNsUWtuoFjXrJO5gmc9Z8pC68KQtwFIc6n5OavDUz2lI9Hv
9MMcyPHNHAqlyNYgG/FPdrsy9dsowFo6amjwLv22iZf88VQCMEGISpH+La7d
Qho6YNVVfe9etbVrTMpReLZ8+3WPcVX70Nw9rGu/XVckVI+b/HbM/fSA2Pi2
EWFGLYwFvCRQTeisDKURGCsOuF0U/ZB6BvprJXmkDabe67GacuOVlUldGn0J
bPJlO2e3SQ15K0QzixYiNI6AWEY41t687SXkMLN8CzlQWxgVZMjBnDqAaIQ4
5va8aOzfp8O48Fe1Vv+mdbXw2d7VT30vFLryUWuB/yktiBlmd8B0o94C8Vzg
BfCCTgP6z2MtGs2ySkfngKKmpoTw605ktF+fPWy6xifHflFdfho9xAKvBHyO
Y/l/VaQmhtMmM1PQ/X/O8WYOUJCkcCpbFFWWvT0KTwUE7EloH7fir6CvqdSs
NG6g1nLR2Oc09/s5z8U/VzWHRLp8rMdWHXMaL5yXYgVUd9QcMMz+ouow+8L3
ikj6UHeO9bEOnaMHAG6RbBPD+jx6/MKwjf73q96vYJiHi3so/Dl1xPBWb7xm
yXj+PjymzSxgRfrWgUythpXVFuKj0DqnxcIv2RPoygaHF86rq4RgiRW78/le
X4O74uJaJTrMl6gPCHTeuyqwr+k6/PO5J1GYxLqW44jUS85E0+Olm0jRTBJS
0sZk4S4vtMiuhmxZzYbwLjwxTLkzxPKEMEJG99GDV+dQ7eU6S3CXkZbawH7+
VZCdNVKJgNMKKq7G/c3C1vP9ISlGWIn1+HMzpoeOIuFD9omRVWljxmwszuw/
yvySn77fmDIVfTlOzT/+9bK8Yeah6uWjPIrk+u8ZZGZoJOlTvAgeyO7i6GaK
lNKvCWQNnJyTQ/J/gl+1NO3tBoOx/V1RkDlRBXeAv9wa6GvQON1lpewJ0Ps6
qp+JEDItNYJ0MRUPHjaDT6ztNqiwExJg1awue0gZSFV8jizspSYo4iWAUObI
E90A0RJrVmiK3PRmHD5D04xxuqN8zCMpUSQc/3yQGp/VUYL7iB5+8fJuiPbB
ON4RlM0PHyc87i1Tdi9wMQOTUIIGgyF9yLhx65y9kluHJKIDHhkNwm70jxfa
tFxS0jTCq+Ex4ot+98kVBrPGyLZDcztiognnm8IxHzvME4Q8mPvwvu31AhTg
QB3JpHvnhuVDxGOhsKAz53DsLhdJFDAkGBJ7t+g7/CTdc8vAgs84zbAVZepY
w85/0XW2Tq3DBx97LXw5uAxe2COlM/zPDrB74vrz3OcE9C0KP9qms+64sb6v
kLWWK99unmPVgypIWEl1N2AOk+mm52KhfcKr/Ks9bizT2a/H6eZlW8vKxywD
drVLBlnIze8ZJGIEsF1UoXPzu69Y/p/fk8FpFThX7kWY6T6OiDISMfHlBLU7
ZxTS2mfKMbIX2MZxOzwQdIgBp1nBydAqAABYFpmC/wv+UjwWvM1FKRwwM5Cc
H6xfY1j2YMG+hFqiIH39XU9Uc+ijMWsnmv6uAnnnfCdJDFnuwxBW7gyWiv1L
vuWPmfvTlT1U5upzp86s29scymE2ejpSOXLPdb/TxW4ufz8pKTXdKtAbl3Wv
OL1rVQKAbYAY1du43Bq39uJl09LdB8SpHK6nydiTDJkPKUnZB5BJstalxp4D
5Mx5lY1rKHQboiACvil2sz9O5iOMPye7HhH9EzlFeOsyiUz1eJkE0YRwk9EL
Pecs6nNJ8eOCiOJrKZoUjgO08b4EmG1fWTVFjbw7XhS02ESmRx209w1sr2yw
bBMj0VEauzhq+AsJZ1ec1/jtiPeetz+P/q9a4NtFq8/9g5jsX5+9OiHbS8Jh
2VfoNqgRPW+RN0saJrtndGpf7RADC/rWs63eMHM123j+f5i2MfJiKUC05dlj
xIneoNm6PnbFNDj2l78ftuyPQmLBwezUHXD9IJm0hWzr5uVNUzx8T8ZETsF5
zzhP4DC3xtjzOlGc6Qi/YOljeztsV+j0ylH4QGzzPlg6SjAuqM3UzgZtxH4G
7G8XuBwpnMGGyDvdc/duj927ZmW3HXHOLPwrwW1lifG8ekW8+jv8CKQU+Icy
OgxzXIpbmENPLOOV97mVgV+7Rzzt5B5flYdljmeG2VATQc+qz3Z664LwTnaj
XHAH/uhCR2V1Z1eMwpyzqW3vy2rCHWz3ySuVGsX3K/5NDLAlqFD672mbn8ha
45nukf2OCnpfExE069IilZQSKEYn5QICQCFfEpF/osQQTfRIaCbet0UzSS0q
Qk9THvRv6gfe+eYItBZVICjuALNNzzom+vlIUdQmFt9pHJ2imguQRgtVcG+i
aNWseSSmanIhjH/qsVCa6cgyFJB4GV8+LLs8NoacxP8eTLpVlWTQTZ9F4woB
CNlkzqvmi+4reiCw1u5cHXpfNN5UJjhBskVOizdfJ5muATc7HIUGA80m+THs
gqLPqS5/ezMfCNB4zroPXtxWaiDrEG8EzxTJWxb4bGzR4H/6O+mDArNC79CZ
PY5vS+cVkZzo6Il0jQWpBNvucY9UXDhlqTY4csHNovEb3JB9W1C2xj5lRLTC
mT30BBB7Y16fM/Ra/qr6U+dmmIXVAjWU68k8FvG8lZQXy82pk8gwBBjaNeWL
9EBAqLxSUfRnnBN8ZZJuPN1kU9RLnrzKDhYoLxWw6G4OerQICi5VsiK0RAEK
Hgg3+m2B9Q9VdNaHeE+MEVVKZBNwbsCQLU/h3gLKpZQ+Azm4s1lygtTyQyaH
JIHCimVibGeo/kfyYiSCPOrtdUDdHYRxx4OuEzwpJhFtbGCK/fAFHf9+LIQB
2QAa2jJEIIZcBRNTlwX80OwOHiE/OC5Oh9pDQe2232+z/5urV3ez+UjaiiHY
xCHBt82s0ldgK1vwR2zdxBGJmRnHlmChd3L5yZdR+bLMLTtbItm0fnNvUE5R
MlhAMMPOi5h7oewSA8bhAgEzVC0O313alPhgCBJvEXYMJwt/6s+UhCXg05d1
HowXJvLSI/qhEoNX0yDrxr/Y6gy2TiX11Ojo8RVrOvn4wpK31YHJeOBjvHpo
hEUfqTE3G5m9gsKb7ogVAGeQF91WSUWas24NVv4VK2DKf3KvaMi75Qhb+Ipr
tp6cSj5rYs08IN/R0xoidzQvcS0miFf8GcRD4T2l+yhPASIfwNfwi93CNbi6
5v36QSn+JQthiMK00jZL4gYs/JIIiyTsmHAUChwl9U5ep/85FdX1vyF/G225
xNCKhP6CcErsSLn8D+Xc7a+XskSJBUvIjYNP4LB+ti1csPLlSmgtxY9xuJ9n
MEjnP46p+9kYm5qPR8Dvh0eg0oPKKWjQKr+THbyMlsA1CTmKmRD9+d+Q/GyU
PW4eqtDJjxIloLKk2ptOQXDy+93mou4ej4t06Ph3zI7oUrIknejs4NllT/qZ
rx+c8JiO1eoeVu7FvGeS09VvyWxJE/cKvkCD4c+XTPzA9EYo34qD/jHlIii6
QMcDaW7QTnXrKeaCYYyuRyfoJ2bQFBPksy2onPlFN9RVGSrpqBAx8kwvdrO6
Q/uzUVN7LPxzispyPdogIg8mdMHDvDll2YeFOC0f0GTwNv7AhiwwEY27tjUw
Y3XvT1XYTdKelWLlHxltEyKBb0B+Jt4h5wpqupT7Xp7WEuIJqhcSOk4H5Xpp
VgS2YGbXlp4pTBMktkjRS8Y3P7P2jzbtXsHNQmJa+c7SChJ9Ak2ZTwq45vAv
672gkYc/Y6NIzUqvj73wMQGjjyQueJSW1BakX63KIUd1fM8rQ3hbtrRt7e3o
z8zcXhspTLyMEmjEtAN1e2N0CBLEA8pYOq5nBbRcAoQztG15UM6BC0dYuPKI
tnDc6b3Wgp9nE1v1Wol57A1a9rDlEBh5iT8/Z6/hWBh0UUrkXCjF91oExJct
s5GQFm63ctcKkuHDm3MZuGXkhs+IVbt+Bz+yYjoe37AUUkU+O1MK7F0cefwx
bUufMZaqXkUOP9RcPfTuslhT8kFKOD9gS2qWsFGul9ENur8PtudYQxAHYh6G
gRumQ1/x80/ETxxEuuYjt9R/hYCudNnUMChrL0H85YP6FFYb1dh6HXE29B8F
IZp+5Omp3s1fnn7fyRn45iO3M6w2Te2sjpehQ+wmoQPDqDG1Si1ltEElBC7b
+PxFJsVtCUQeSiBfLN1k+Hmqvwi9lkVXmkUvtuGBn6tmWIQ2dL4S0axhOm6k
epLzG/X74Gf5yO3XfsdYKmbD7DE/q+5YaAx1E80KfE8pEApr08/Au7hwzEe9
rnuhYb/11Q+ZaKXdWTOvgjXn1s+NQ84saXW5j+bKKu3NdWjjg9E8Wfwqkbqu
8kdauJkRFCqOh8kNKOoIYO4mZ1Q6s0mNHh9LylXftDYnhV62eC/yFLpvOmRc
z4rZzylsBpvpKJ54+c+h5bNa9u21sbQr9g1uF6tqHkt/3ggXx/botHw+IuVn
qa/n/L97BFcQOkqi1THUca8Uy6UY3OOuyFAtF9l2wR3P4nn+jxx4t6iJsb3q
4wTJAJpWeS8xSG0TJS4LiVLs7NiwSYUkK3vq7weB+3wYNgMZqKCNtxKFOZ7r
EN45IxPfNYnnSr3bHtK95ciBXj2BW/Pwl/uE/t1p+xq31RKAXILRb5UPWjXY
DnJo8r3NTMaCCFiTTer6GRBlt5NGM68t3WmN9QT6pd9aNt2C4EKVDYWuqmrq
6YrfyMUeTEEHtAjXvsh2gXjrzKf4dSuvkF4JeLJBGELLnGKGf0LT2226uVvQ
4hMcsZmVziqWNcHPsOQyMGkHqlDpWK1y44tmJCH/D7/prPKyDQ6WnYCCDdnB
dcgpAuJT2B6rHex9dGQvBuOMhcJpp3+I5EN90e80Anjz4xeHxTQs/O/XWzYH
5PVEThjD37Pz1VQJJizCAUrXMfanaBe13y6RRHi6ocwJY5E7Dmbic7GvMtMf
aLGewjSjKTxdHCmVfUWIGEWStUakvOW96aCq47OLKZiU7sGWj0U7BX66hPsI
Db3QbAmEzIDyfYAqrrXuHaUPBXQ8No8lYQtE20QeC5D7I58GiJhfr9OyYF7n
uURcc3l1RSRKkHA3e9d2f0NhzOSH967LBk4c1dZiDL1AS3wB9hpytPoIWfkB
E1cYc9rDAVACLp0Bclkhz7HGw3rrddunzJjfwbv0pbZfkfN+xMfFVT1NSzDv
8TwNx8k6XN9dV8uLRg9jkcFMsjhSwIOJ9XR6ev/C7f2WDUWSKYr7tOcd/p4H
LpCKLOz12x+VvMWQd+J4a6j0RclqHeqkSgsrmlr4Uu3ov8hVetsIQPQGVaXp
SIqZ8WSmjw/rtkiEKezS/s0ZztP9994Cdt36fXPCeA6IgXInVF8k0iGS5R46
Jo4nbfULwAdgsvErzg2O/qIU7WTFGOlwtoEb1bLuakcAZkOmNd7rf3oMe97R
c7XYrQkmYXJPtNmrF4IDnFdq715bnFaFptxOIs8h1Rz3A+WPNWQmOcJM76Gz
uq8kWNWYeHGI6btctsqbU9Y0fTWMn1wg2WK9A+G0smXK1tTukJpt/jwhO+r8
1lOcyNrTTGxmKMIYEOYGw8Xu86ZNHuSNkjv/QWuc39tnXkSuv9PriLW1EXKf
FBzziYvACNccudzxVXlegq7funlWkz+hDbtX3QIUQNYUoHOKAQkNfUQ0kcfQ
AjaBL9lzHh7mic9tl7cGldJ71D7E9/Q9sEs3P+aCapO4clkYvstXKAzuulaq
njs+UNUp+CvvC69UhZeJfb/nwe6g8WMPw3kJR0qgwg1hLsg9iroryDLpl9ik
Mn1Di+WLSUoSsI3Fhef51VxBX6hNynou0XG4ND1wqFfMUC7ua+nSdyNM3xn9
W3+rI3Ur54ZWSHzKLQGERZJYvys8F9jvPvrMGRDysGZw9P4udOLvzb0RqfBC
0tykn6KAOzxrqK+VBfVdAZvxzjlEnGtC4Wj9dpkXZ68t5ksLC38d20H8phCj
A8OrhxYEpEsyaY33M8oT8nGOwUKg1MEJX1/jTFEkayYUnAPkOs3cjJYYaGnN
OtWZlSMPt4mSsHmqtCdP2lY8VBx5PBsf1sQS2kRyLj4koWDH1Am6clHLmZZx
nbz0uz9coqW36Ww/N9phw/9vBUjXKJxQbWYaSKxndRMoxYi3VUgQRKsWngDH
LjXYYPqzcIa1b/E0Hl64vBw3hx4upoIxm4lXf9bpkLCgHVcGCYA3bKf0oght
IC0s0+hj9ntWOyJTxKK0cBISZMgJoGsi2dlIyuoFuPFoyqv6/lrCK18n7GsE
G8OVpFtgvnKIcuG3gDelsxuOR8VElWwZz9JdbzhgZe95stK6rFuV4d1v/SYY
BdTuDXCBVSf7VV0qE8EZpgz+bvNThoXe0CdJrv8eHKZDevzMEhFhYcg4mcoN
KheHjAMbY58yic3PW+Skf5OsfIJ3ShPnCK1JAp48mL2cq8CnzCRjstTjpnV5
3AEp52FDmuhu/rPdp1Rvn5JOxWNUdTbTtElnMY02KRhdut6CjSUZGxz2IvVL
WEf0iDM2V4bRcb40MzCyxVymFLRXPeyvvvneku+8pZpvSDSKm4raBaWwKGHF
qi6fRWj0UB87g5Qe/DXTnm3QQkkbNieYteb482ECr5nToABSqVgckCYaDaa3
jNRoXZHDVuGnh9s1EyjWUmg/fTe1UETL/L00T6UBRUlCp/wmINRgs9502lpH
A2tJVb2cZETuAyjclVHZ97hfC9clMgls30+IoQAzdvRA8N6qFLl04BCAOtJc
L1k/qg+A1SKkfsf0lsb7k6Lx3tcrQQ4sIEFkBjNl+4/y9GtHgYN4B7gYD7y7
JiRKqjwHH8w65DfH8wABp1HCxwyff+7KiKT0Yp7eEppXDCs44pd94V6kiiF2
quWAnZL8TtFfY3C1B9nKgtttNaMCMKcj7JbH+IDMElTRMT4Tjg8z1HMVyoJC
3fooLgg+aFr5sfRmydwXl54saWsBPT2YvOsCNA2nJ73Wb+C4/WVDR6V3/I94
OK9FUKF+PZfxsTnwgXMK0vgra8hTL4F6TAExab2ue1ndLtB9AxhpDVGdanjZ
AE6/EDPU3k/jPXvJVvZBBxk70RFVx8/NAqvndQ/MLnPkaxqOY30OqmFxVK9p
RNtU1j5my8oJFKaBAPEd5MIf9Vr5J45t+s63paLbp47wqJEZgVkBjK6eYeJt
o9F/81vR5X357SD7nbllJk+i8/upq2HM4s4qZ4vQirbTRH9Nuha1uFfVvXpn
qEGC4MgbDyXoyJrl9L+eXlMtoUhorBT+ijDRPOo6tb8N6ZnxTtcuD/9xSnEd
zOjBNwOqGjKT8/8bt2A2DeE28MH083R35vSpGctzhxd+JBz2G4K/t9nODI7e
NpzcSjIzChdQPFBA0i1GxIHXFRviXhSwa8/vKkA38+WLWap0vxW9akuJfdah
WtU2KEhiTg1iHn1i4c5Wilj+UBti0WaxH2B3BsrtmW9TqT0g65/UYxMjpais
aDgUFKlzKuCRxUauEhu5ICVcKrl1jiwoqJ7TKp8+zL9IIoO6oB6JeuH0MZ4E
329CvCglnM42Wy1FxoQxAYBJx3h7j6kM4VHtXmHbv4nIA3+GAs31ZLFI6tDb
DPGdouAgxwkx7gaoFRN28S8C4FOcfiDygIUTATCVODWk2rcBSnZPYnReRldY
TGOEKUNPPLYSTFLWjVVZWgPho8X+inTWWvz3/LHmtPgn8wcbKSBgFBLqONbM
mmisb2iLNRpsiAyKfjHm2nIvG8iLs84+vxhP5CHqNzRx9g9CKyanuB+qErZ/
N81ecYmdTQlK2MvPT/ZnoglnXDOOoCaUoNeJnOOR9YB/N+Eox+N6CFqU0S/N
fV/sKlqLWuwJ52rRCg/haTdqz7/0kAkzZe4DY1B4qGT4KOWgcuYesp00esq1
kPzXAoIpKkHwLseqEkJaxLMuKQf4Bui0CSDhnXDQrVYFXjBibQep05yvzG8f
hLNwHnaBZFIa/0FZTGgib2Pmj2yv8AIyt6aJXFUMDvZuCatkPISIfl6lJJzY
jovEj1d/0AyRE/YZO9vIyzVuQmah7EJc3txEAkJ4rx1gAMsj0rk7DImk0KA5
14hlPCwCNYxG3zoEpdYOaH/CHsRxiNLetVkbj87fsr7u/cMOfSJ5e2BEaNAP
Q+l8ylLd6O69MyL8qXZPDH/pGxixOOV5JH06nfUOdk+EXFq0tdpS2mWyM7nL
9DQn1ZCfVTuZqcRpkRKqnC22sN+jqmNI9uDj02wOvwcMaSTCnbdFsPVSv52b
N0JPY/UevDBZkbWtt3zluoSdE3TQ+IaqGT3bdzgwYyMwDhkzMOkfGT3Mm8xy
svo7Fplg7Nlfi/XQ3Vz45kZ6HNtudkXtaAtlMP0AHhnna6VAPhh75MLlySND
/meO6TWCr9izsqSdF+vgW9uWVEH8c4lepeAsg316fEQHkXNg724/otUR4jIw
bPTEwHHYPAFk5yMZ5U7oKF+Vims2kmK4ucPnAAo0TOWi+OelvrIb0t9Pc8gF
557iVKGRgXUdnUZpvxnZsqt+vYN700hsMkn8JeHXRTAoG/pDPwXOI263D6Sl
XxHxw3I8Sjn1bC8ZWMw1d5cJZCKJdsf1hlsb2olWsSy1f5xhjqCMg+9//Fg8
I2Gww74ZIEQO1lHAoXZ24On55o9QVVTgknsfd2Ngh4F9liU4ai/2m0+IHC1t
OGNv+7/yUR9lSdj/9piWgIt2HBsdTlZSD1DYVhWR6UygGGh2s5jZFVa2dSF2
givoY8Q5lwqLz45zTwBXaYs1f4O5OIL14MvPrRPDIArJKRQNIAjTHaJrdqZw
qH2vxCW3Vj0qaEiwjA+tyyNeIm1wBr8dCeMu/WIZ6xf/TR4objc9aj+212cI
Uybl3DRDmNVOG4Uj9agViDCR1zuGrYFEI3gHTurxt+JIQWVjNzfjryY9jqwt
kLd+BNGqbEiKWvFD1JyvnwuubE9kH9fc2UxNxZRwjB08oQNYdTq9qC1YVXkN
Hmd1FAdbF9EAgXQKseCYc0JJYEUSw0JxvVw+3loslmlQ0jy3YYzIn42WHrRN
368n2AuMnXoM/e84QY6a9asKb5Gr+bkNKw7zraKB8gANbQtTznt9XrSUVisF
/BbAf+G8t8WTV0dUVM+fUe1HQnrbeCxg0e8Z0VmZ/+BibAiXMf+bR1YNUYnt
Y8U/4gczib/jVP/SR7KGEwSOKcP62YwRjX5L4XEQxJ641uC6tIeRGUQFj3ZJ
4fJ51yFtjRFPpST+NF1TZODOhrGpa83jVhAr8kxHxgconOt1VzQcfKW+nm6n
2ngDS2BLCwWAXwvz8AVbuFGEni3gfLDTbdMHppJTrKid+l9bqtyf1cZ9x20E
UAAixQPe8YZEjKuazYLMWRIY4XBDFZcfcuoPSCZUi9XlZ2oKqaa404oQqbcW
hmW9gaa9frHmkkaO0dePY48ufv+JhPuHVF5B00Fl7jvNR8UY+NJcjnQVQeOx
VMLNd7LYrBeFnfriROArOd25tsE356bOTUl1IPrbSTsFOrc1czIowOrirG0B
ZOJL32ykN+StKTeSUhKSqJSuwi8AVQUfFiWDTa03PE8sik8Rade7wTkVhVpT
XiJhFRREWYFX4HTdth/MFqB9gz3a89Q791d5h0RvSM/r54+GkEaVPTxNa53J
9uruFX5X6mJdRAlbT3rAosAFZceyGp/8LbmnedEYQ63tm4eB+cbjXObuX6St
j48S7bGXRZBATDOC2+ku92aFowwAR0ahud/lLYv8JZ26gz34SkZJrre7BbOD
JFtUWmNsPAo3yB1lWI6k/iw2x/C/m2eTsbqcj+9SgZq3tjsBBMNWDM9qn34m
wtTV/qeW2etrML/HDRzbqWK7oeqGe1h4uf2q1wWywqKgmfjTd5ZjlFZSvk+F
GVTTq8JwndR9bNkSIpGGO8laDNICP0F6rzWyd+ZBKbYQ2RcJTRAgEHezHoEW
8HKnE5bxQEUEGusgoJY8gWWEWAlfAwajmf4w82dL95l+Rp1RP1u6N2KqdSG+
w8DE8UEaMZ2TEHCEQ9nM3m0UbK81tYJJWwG1k1ojZDnNSnboIaMgG2dQaLYn
S8+bIEUzj+IkSIK8jHcFIlS5rd2Pc099pdsfmO2s2k14//+KCWW3/3I1lwP+
G/Ic2bbPNXHp1nDilLyyOZBS/wSrCFtiri7Zf5WYlBl1WoWvHGKLCXSjjF1U
ZaY/jY7pbtfoNTDLJPZJI4VsJx7Vd9ZVqYMdlyo/CXt4OH4M9MdeRFveIKPv
f4F6fZ4adcITS6SeJ4rHp8ubZGaYlu6j9yPyJZJKckiXiJrMoxCzTaH2He+o
B8ugThcyyvEk8QszMZr5w5gK0sdt8mtkb0TlkT/oK9Bhsl8Aa9F458pBtrGb
fWyqwujt6GwnoqVgcpr91KH1GTDVI0tzZrhertebFRnbvJgEaCBGsb5BTDgY
QHYc9Zih6iOOlWQ+gQYuSjSVTigO1Tj4C76u+aCHzgBsDfSSvCmPqqDwhC9e
PztzcBy6QfdZ6QDsg31+Oe+ZQDUL/uCg5tY426uRJqOQKe+Y2a+PCqXRHtCT
crYgRgsgz84r2Fvem/nh8AlqQO3v+b1+DpixT2R7SUBw5zSM/tIu7aSwdRrZ
wvhqjD3/mb+jsBZW8iUMZ8o9ok8I7QuU+wA+GBc7/w7E3fCGiGA6tMKzXvpB
i+cgdvMwzT2TTOZuom5gzI+OSQl4+GvF/AUbhe2YVHbrDQJCaMWJNjHsegC8
zoyom1dett1tzFv72LUF0cSaYPlLO7aEWVDDmidCdUJ1hoJjlR2evT5tVUR6
YxQ7Gkoj31TJWR52k3Y6mgAgpXnbxb34amo/evVgrwigOOKrOrg0PNr0C1wE
wyaUiBwo/PFt/KcjuuyJ59nnAQ+bUdwXzKvB1b/Ba7+9cohLR+ObfjNxECdk
w4mWxOkRakdrNaXDYf2JaFZas5tZxrX4o9I2ekj4wc9odknpA8oBwJMag9Un
yamgzu+ha88xmfsxkr+uHS5so1TxCL19LFqLNTdhHyqs8mOx9gTokNKNro2X
9/dn7GURJ5YZEXNkx1lpGNhDHLnTMHvRn5/Zm3upPVHzMHru3/FBlvUIAPFL
/mn/bXi86kCuuivAIzKZ8CgLGgwLiVBln3HBuzk6Vixko02BW7RPDLLHzJMO
DMP+2N2F7kfnnBfgxGLpBLZG2nqIrdIum7CTf+EwXnZPqjcyfxUwjLgeBMw/
+L9ZjmQwRjyXpTy1Oa9EDW7SF/FB7OKZIrQjXRim7s3m5ChC+/Oqhzf6XyZh
wHkxnqBgOFGMHfPW+Pn2YGjDic7ClOgQA6hnp7JgZ/EZfOLlq/rOXDjln/2W
iyyn8SC3i4OCMSU6PqxdSODhzc/24BPPb1RS0+uebmY1lOaLbwQZjB3M20Ht
pTcuc61QKCi7eviDTqlHP6XyGchnUHyk3MXBwQ7Tbyys+5iIkSafxeCLADf/
RA3k0600CyfgTl6gwJOvpcS2iQ1UfNsV2AeWwdDFT0LS4xMG29tMgKD3SS4+
laHA9wQp5aHmSRvSyno0aZhxkk8gA1Y66ipmReIcOgjWact2EGU94Urt60w6
S7F2IcX2i8OgoFnK2XTeyMNX8K35uiDQzZtYN500blmcwIvQ3MlrDyOp50cS
KQRD4k6lgCohR79IbyNeVjzCC3X9z832uoanwt0Qe9y7E0zhJhb97wnbviFL
rxE5bzRJhRna4EODTZCo5DLHjjSn4C1V5umrnnil6mpASNeYdctW9pmyBFoH
C82Av+W4/U1QtslAkCuX3mA3ndKFnPws5CqUHXuRnYu4SoijIl3o+UNbIGRh
n8WmSwT8bbiJt3VadLiz5GYKRwcyz1wagqL9DJoRNQ0PTwGpptSCm3KgoGDA
3C5tEqB0lpek4NxcyINCJK7yHZyEab5Z2ZSR8H7ajoUcY9W12FRegynpKPJO
qWeGJaP2SGh71/8TrA/H7jQUmu5/oEBebxQG1MJz3BX2HiIOmCTiAoJAZCU2
tucEYXSj6hHKkbZQo+p+gqv7vWoG1HxBadY32UOF7318F2wW4ThUFPMCrAo6
BDEeZeEnmA1i85JCoSgrBmOxu+8yzB4a82xuJx4YR7zCQGVfZtSqYMaVaPDc
x7zlxyH+czAOTqnjOAnM/IpiXjE4+zYJsk33sEy3p9oeOfpC9eSwYeMb/Vfe
0Y5fN7Q0KGO4od49/jixFcXfpS8wEvVnTnK8ShiTo3AcEuvtRnkYMGbm1qiH
SXuU7DfojMUJ3Zi6+PQy55kL7TT1NlOld6kBe8CpcBTraOP2qz0ui+d4+TZX
0Y9lpcX1UO3rR6sKx2j/88A5smIRHeWcERaG6K54Ya8mYztKnU4alIhcXyT6
o42vo75GcEBhy8kxh2cYn8kOeM2FNGS0TsF/kueImUjxObQXxRss56xtH56D
gaHuoeIrdDQU8La+m3+RWVDNqT8oiKimDWcLfR9c3vN2by650RPSUrAS/M+g
k/Q0CdWQtJTjnXkqz+rs/1dXIom9+eUuDoGwxymVsSiAV4A5MANFBgJ3URIP
jhZQOHVtPyCnVqX3XqN5QdLqD/eIIxc1TRGoGwQh3uiDeIRmTa/jQE8PklDe
wBVE89NecTX/nR4KmukDgtNEQfWDHW618e6s/XXq6TWHw7wTvsu0IdKAGWQc
4yaG96P5IvOqSw2IZM2n2rksHPIy4hKgPpfjHfgcAPEYgd7HTE54sHHmmz0a
LjZ3w4ybb3PRWgWKUsM+bx7sZVEeghYa2yf+KWZa+rdM2SsCta9qCiNUgB5s
tVxNMVooWI/NroZQ3CKSeCdy8fy2NLsDsxZRJL1rwE0ThsyglL8FE+C12CFg
hQlwmTq6NaYbrhtcJ1WNrRhBQNtrQXi0KmELpVgMNSn5riw3xOH9+RuvjuUw
Wfbn30iKpNY8gIccLduGKwANVZBXNW/4Qipt+r9432UlWcuVsFU72dSTZ2zI
10Rm8vxnnzoZrJP6bHM7WLhhZwdGOaUBydOgIs0CRsedRYUZspvUwiViXQg6
GXzN9bLu054arrzjSgV7Z1j9ZIlXpOFa90AMD88zEMvOOS4HCvz4oqs/WUz6
SGquR4CbegPe8uthvviHnaIgh6KdU7Pxuph/DIovsDB5BuMN2yfzh4jskw2k
yw3PbQmHq7nMCRUHtVfE69JPiqN8K7AvJbUo3tGu1pr9lhNnhNMtLjd320O2
IuYfwn3H5mMB5si++OihmCFxvVDPKyF1DqOkQrKrMY5k5t79WuSlFYCRVcnt
92cToO74XfkTHLF85jY8xdNjrWGN5PDEZL1/JKNxi0VkA/y1RYBuX4sHAJfK
+Su/FgedoBSyxGG5HIu3bHB5WMnE/oFVkuVkgctNA3bhOFJD5sroCFXfmrcL
KY/TmorsY61Q2AyQn009NRgrqFzy4jaVmFOM3Zqx+c8selpUl4ueL0t5hWMC
Q0Ks1Ow05mnqEFRY0EJ7rHgadZK/OxXqGIF5pzIL1JzFGhua8jwDImwzlvN3
2lwNZ7qXdt40yNIZ5td1MsYirahzS40UPJLWEWp1sDiHJISW8j1nNDL3YO8m
zUiUEnflxasQ1Nh/xW08qKuP9BWhUl5ZlGNciDyP7e00+dgeYm4+pfIOPilH
PuFxdFwIWRaBYH2IOE+HgVfzXRDI6fC8BRrlcAw/7jx/rTI14VXHYmsWIjap
YbYSXbpoOQCC/TFJuJIFesQxdruWZnv5MweFIke19SDN+DuGwe/4K5TsZ9PY
LImZGSiInncXZjr0wGYVtIrRTTPTUU9XiDmxninbsVBg4TUWA2A697oiJoLw
IacLrykh/ytaY7k/C1XzpDCIIkCzrq8um8HgLQV+nP0irbDQ3EOrYI8w21yT
hoCYgHkD+59QucZQoXFaSKt2/JDP+X9S10eHMTvE/xU/fvbFCA4kgDfZ2yAM
Ee9Cukx3Jef3hnhCp6lCLoFxZk2FbTiuc15lmiwvo5fiVdR+KMZtUdaSblxd
uh4mcUsjbJXY5mMtgxsDnGX6NnO6CN2NPBivgPeDI4q1cNn+SsvvlVIzasCj
L9cNTLiCuOkkW8j2S/jvwHk0kxMsv/5hTxmqyNN+HTOfCx7isTIDIhNQmEpz
xw73+OnMXMQtVy4WwzRUsXCyPvVZF096UNqwWKB7pbHu1gWkeaaQAyWMFl75
+pwtLqLj/BVHW3tqfJ+DPKyInMsBAZy65L02cNe4l6llAVKnU+no/z32bu0k
A6aMsb0l+Fehyjv6oyN+pBgvspBGXK/yY+bjJKoe6S5lN9sn99kKS6o3JtUX
CBFlSwg31MGEIy3VOUlymQgOicUfwaqkthEmhHT7xVOiHSyKr73PmgEWu4PJ
/SGBThvkxNuwWEveJtZ+j3JP1/rsducZL26E+DNwbty+E/u8zNLNDTcrxZOq
RTDVMmXjOTG7v0idtq4y/GHzA+0CNraOFpg/9FM+6Y68jCm34O3L+xgtplOh
uYdiN6iUzO09ErlLG8LyIPqAK5MLGu2IDrnEBeUW1elKWdhgyuqb9YR+EmlU
T8e7Uh+geJNT0BpNLpD2DFgKki/Fr1dzNxqry7/Prgaur91tnfsbCFJt2BqP
tNzguJoVXr6x0nStDeScraonwZVLaJVC1+wAYmM1JVckmqOyYEXmgf+eX0iB
AM4q6JZ7GDObUTEDREn7kpToMqayPVt9wB5F+4uSTNKtkgU00T6qrA0I2c+c
K8/SbUqVuJ7hGbyp3/gJPrvagUpyKBmOAS1/jnZtWNcUW9UjIwC5mz+hTm1f
8zoW4KLKLjvkwjTx/4deZeIuUA8MKynPvrXHWlpFjwck3e2GM0NnYVuP8K15
AfdiIZ1DhK/vcRTn/dLNYKDHPL/kZTJAr/vhqVNLDSf2Qny0WRkFfAr6/oum
NHt6IYVr5H2MpCqgFmcFO13ihu+TVpUqJkaQADbTVCACQLq5Z7MnYqKt9FDf
/g/dS/0KzGZkPNiboFx9E27vhRwtmnWowp3TzlhryH3UuEsTF3cwuYwsg9z9
kC0ZoYlj+Kn7Cjbg+2dAcBeQfPmq4kdvW3yy5KLfuGc4e9m0Ms/f7euaSnos
VFmMPFoLBLP4Qk9v4Dtlw8/2WfA/+3WSBXsWAKs7LFCB/rd4ouPyZQoJiHaE
uUtQzmBfmEs95LM93bwKr9S55VZtJelvwEEQmWlTmnV8TSk4o7e2bCUiTEPn
uaAQSufTQvwjsTLq5OPLruc9qL4lResdKtZ2EOorYtvtc5dCT7bhbstpJeh0
lqkMWNH+dZr/YTzF/1AAut3zmHauXkFqWOIbWzCiqtGn1lt6ZUTw4yDCAsUx
Eh0tpf+P1OTJmopoQOgWw9hUhX4EtaXWiBnrvNv8VfVts1X86JG5XfH01XkB
X90RGlNgEy3VcNfRUTV9iIX4dSNsvM7wbiXLKoUpOF+3XC6A6Zk45xvLBh9u
5TBqZ2mElLISKY2fwbbNbI0QMxG/3jxHZx5b2t3QBdsbrCzLo82YQHF7F/kG
kz+9miG76mCRQ2xNc927TdCLMFMwYYj64an4O+y9Z7UoF2QGovWnXbJz5aOz
4r7wpaSWDfv2Y/ZO89mThXhzuwnR1UFH1pp/Kg/yAW5IK5Qwv8fM9VG9kdPa
7g+16Wf2wdFXD90iQ3Pm1MZCcUwIistC2FUuv5zw6sPMxzE7b3KEevQmTpKJ
w7o5/V5LO/I+RznkNh5UtlSvclDCEi/KDL0psXn+I0A7mS+OLL7F9a8Rd50z
5bA2xeYWauN6+Wz3MDZJ3PZXV8iQatRAdAQzk1NBownxB/ZkBVrrrShkVe0A
FP2EHyRFaAPCv7dhQ3A99yUaQFFAOETkQwVs88rsQA2zubb5LBM3pScHcLIH
zpyHyE2Ac/+dx7vS16915jw4GQguWzrPl/MVg8FNchOsPs+N8gBGcoFhlakI
fXLxkxx0ZctFNG5P/F/rqXFttJ+98JGvIFa9FBtJ6p7ViiurmjX7NjXol9cu
cAqpirBjrzlqhpJlM3LnI7mWBUUJVqoZyufnvN0m2VESRyE4xfJ4eYhCcJu0
GcQlmzgdlAdwL3tLZpd6B5pRZjT7dxdixC2HofGz7hhwGNjMUOwh6unFKvsz
zbmkNiS1qNmSh36rAV5ANlBPOqOI2Ernsi13Gym5DzgAkq8rUzp25U3KSRFv
OI1pyWMV7tFDGSfh4vljyed0gWdfAocx0MsNmQ9oaofmbYlxlRkgwU3scccB
9pZCttT+Zz+L5YEnY7fmC9Wl21RUnch6HxnoaRaRdsxnHI9/9QeCCr5r/RAV
CGRKCF64l20FLoFcsWd5VaWc8tdWpUZLvOtdo8T3rMslpf79sYWE7unJakKQ
wvnMXRSrp4uvjk7jTzAV1sNX0z8J3OSVg5ZLCLCLd4eih84CFwf0rIeq2QKm
1E1QlJjDyze8aj/L3B5sdseW5l45bAoHRe3YitFAeelDGoNP17AALLr7X7i9
HvARhPKJbC8iBI/Rvnrm+EC10avPgMiUSD9vFru00a+EUjM8dIOfvvBtuOUy
yXAsF5QhZ1eMsEjXIv3ScUX6mldtFUA9m/rC6ETycRK8LBLUN+TN3719uMys
S+bP04KwczEd5MpaEq/yY0HKrDngrU262PUr5D4ydfFygVTAelmdyIaA0KWM
+ww2nsZnxHUBNrE7vD6gzyA4gykCErGFmm8nMitbJXghZxUt/Y2ESjwZD0qC
YvfTF8xn+AM2tpS9QWUzTcFLshJ7W0w2Y4rdWatU5vQ+EbnMGnQKICH4LlWO
DYfp0At8aF0gkhUyijwdqVz3kKbP0A36VVeBUMfNQfgGuki0yNNSgoc3mGF9
t09pBVtRMqU7rVdg/SZpICy0LDR7v5x54UVKt99clhmc3cMQXa6jSP8kAMGp
ZxgNyp76c8HJMM+ebdm/D27ODTLFgnAotzUFF3/+CXZU7TxVbet7GboSWB9h
jKmUrmMtbUwWrCofaP2GcPnpweCHZkv2CmPcdpQ9c+2jLsZvOsgaoNcAXWw8
JE4De+cDWdNWiMTEokd2kxQb3/ELyi9ZSUY/YK3Gc0VwcbvUsstuiRrK1j+d
l2ZFS2rCUApfz2o+eD+KwKSGND2FVE2JpGnSWPQtvMLkszCKpwSW16O2bNU0
FOFxtxj/d5YkflZAmIBUDra/FIZ/gaZ5kxafMSBz0kTZWI3hviju4D2CDi6w
zd5V5YDwVIfFv7iGAQQ5ykxi8d2pmErxcc5AEgAryIih9yAn2QRrO9Cq268z
XzeyARa3G5Oozv5F/mvDKNJhvX9dnObhHwblu6VV6xjTSudlJXvQEuCsZgeQ
vW3CQNEYCH4z1T+T9Qv7WXabKb+vZpHS3GBCzrz/8b/x5qG9KTji6Tv/MI1+
kJ0sZCCM2VDWbHOZ3JAbWPd6C5p9w9fhKKRdq/yD4A+Fnxhb7pBT4cm+lxCy
U4ZqQrc25+MiY6Sf/1GGB37oJgdLejICNHQVvMuOO6kMFSNymuEDmsMEl+fT
OVXSQ7rXdv+hhPFYl0Z1UO65KUOAJL/YZRFjsGe/6u14JygeC3Q/zSRXpzFQ
/vz3Xl7gjB3RrbHnhhmW1pbbwsn8szBilVfdk/2Fjjg0zmNZ2LvjsbIGPLDd
STANB13cOKbio0zd8QBzzHC+0vargb99jmYB4qQIwOdBwXBknKNhzDg742lD
TBFqAJjZCCZ64/NksEeh8aTcu1Q6rbj1/qbqopGj200FJrHY2mqcuzvaniY9
ubNxqnAXy928hPDTwKVjGg0GeE4PxFe02zaXSVWwuSyPCWoXQe27BNSGOy07
X2mblLWnGfIyyxggcwJeDY4J+HuCbZTiEGDb+5taNgakxNlgZZGQQGP7DqdL
l1GD7gBG+Gf+d+RBdDN36AS1UUZWpgdCQkT3UjHLjkiktC5p6x94pz4Yi8I4
8uZ+x0dUf0d8/oiVtV1kqmgU8OwPsKUwUKHg2fUGXdayGXGugc2xiAHxdWfy
/Cp0M7iUP4QwCkIEFcxbcRJWwVNwHaPEgWB1ddfXN43GPiNmDgZU8i3IBiTF
W5Dr9EHxxb5vrBQO5rhILAPL5R1vOCf03e4b2HXy+WSfqfdYu+FabOs5JVTn
3fXRjrpLuBDZoaZk484dE/s2S50HyA/8cwTYGtRCDagqPPj+TsNxZXafyPiK
o1eHu3YLQrYofXY581fNSqHz35S4QUe26ZjvHnM7dLbac59/3n8UzdlvKYPg
N2yxNvsyuwEgaHIJQKphLaOp2KD4IjjHOR8FUDhXMEeIIMk0KPhb7qijbcRC
aSoKoDT/7dco2/kZxRoEopPphrDVGR1RA6ioSzJGXqI6GO55cnusydRM3KuI
RAAxNasfnrszZmWICvwrffXX+vEO3eLH+TZK3SVNomJMc+/MP/L82fmHtwpx
sT3DVxSZw6aoTHUs5VIfNx3wUChXcwvkFt9K8f1W90mFJhPl8uaup+1hkCEQ
73K4XBMfTxK1444rQ8qCpdRK607MQDQktoHLbOgHLF0Gqy37z20AH2SyC96r
lKB5GlQIfZ0rbu0dfflEH+o8CKljxUA6duPM1FxVk+zXbIiQbQVOGi8ZA02P
IdeRW36VPpWfpdtCLk2qP5/UUzs5gh1VBali4VWXS+jE5etgoX17/qrJ5nVH
//FWf9VoxiXHUw0JkQYla2T+wjvJlL/KrimfaZC0rQyClO354442yEljdrpQ
hNesCW8D+5vD/746FiVX+g4oDFUu+UgjFdPajAR76kEr2QPdxFVuNwR3V0no
BBeSlZt7FyuDt7C1YQFjW7Pr5/FrzeD43rOwf8dkg05DYePsRmB+742cNQzA
tEmJ1gKXfYAMEqmS2YkThZH0iK52D1S/TinKsF2vKq0gqNLPWiMo0OcPBJt5
tkpK+QACFOinmSjTDdcbdXYDCNIJrQ3zlUVQvg98HCSZhPlzKuCqsX2FQs4s
NOGj6hi3tj3SdXQl8tZLs00yAk4lcdgbryborZATQwdMqhSU4jJ+8Wp5u3ls
HTYmEWJqwoGcwfgUJqSa7nLwcG1HLmPPOxALFiZOoDqgdi6A5UkwdTpAaQBa
CDeGZYtiDCWGEp1YPsC8hDFnFCbat7OMrPYrFQImPEI2Dbp2bi1sP396h/r6
iW8IfQzJxujNJ/SODNthSQYGtE0fHZobLFM2nC5Z+C++lW6omtkJmQ7xss4r
aKttAiuuz/YlOaPgWweSdvyhqMMU7kb+LXQztZYbNU5Hq+rqLQlkrg5DIoxe
b7VeGFzCrqx5Qd4WqhGO2enImknq+rd62LE/0gyCTYhUDozLzsTPODcAcNSk
IH6aAMxJs+GgTk8XYDEHSYPr4ZzW+r3aNiD4TDVGSSsZyWkj5nn9R9I5V1lR
1sY/Xa7/Ls5TVuVDW+vUSWg/xH+kK1lwrFgGnyzJUnvSoRS/SnE2lLeHfpu3
NFnTYdi+BHHWWAhRm3DAiN34AqFwn5K9skQ4jq+DfC80Bdza/sOS8D3yFZzW
cCDGPfRfeLcBHpO0l94T46fYGlHahd9m/qQ3V3MJAYoEBHRZyWYaen/kqh4Y
m4mkmXO++S1neDvMyzvAmBTEmDqzYB77eABseMn++f5nV8gWdeFPqVP389Mn
VYkxdpiPxJ7j7Xw+6yGCIOdUzAZiL+8U1HIlZ2PAPxLemegoxzNioobqhF79
RItKT+0YG86RB1TxQEhTWOK79r4bhhEgRM/pveYwtLXi/1ik6frSXrUJpj/R
A37Feg2n/3IWmuXfdZHqqnGVz8YiIW6F1zhZkXcAtQa2NS68M+4wR0CXUBbR
WYHRxq6EkXYj9901snugcaJ0c49ZWaMvXM4XJJH0EOGlrWrJ0OaAEW8I4HRh
nONDG0v//QwTjgBeQ0ezXLhFQ/w3R5fg2nQ7gzM7FrKoij1+DM4iJeybL81M
L4shkFvAMATo9I2+2mfSicBpAcjB+SNTFpLPoYSHTXTRE1BmH5XL4JtKdPY+
/hpQlOJr+/wCnOLIkOXN6+Lx6UQE7w97sy4WPFSZXuRXas+FtI4N5AWU9lCR
lJk9CNoz33g4XMqScbPMY/Kx4eszuk5nMtITe0nn51k5c/06UbDH0UdxddPi
YD212agYn4V1z25BqwIsWHvPDLaHK4DDGFZNIpbUkuPBudUgD+kBienJJC1v
z1F0NvtojTp+5izwHZBeJo22YbrdofQ5MFMs4tezER7NRGayFmvQ12HKO/Qi
ybM8u1HXdvRT0oK8KLLVVAPYUol0w6CIGFTP5mlUqH3LeFPDTQL9NtRcn1HZ
Bbvcg3LI7j9mnLxk7VMNE/CaMEsvs9kxLxrgOWjvN8lNp9+RlcvUQh4N9ixT
G1/DyUsu2YfLXg+kA8804Mq+eH4uQysJKoDL3IHUWYGMyuGWje+tFLE8Ocsh
wZQdSnLe57+dj8gGsxgN+22aUaXqy0bbG3mAuNyxNh89/DZ8JxSnesVKS+bQ
wXLC3tApUgeUEJKBHyatsOdlkWCuOYN7Y0dnjsdtoulsTPQnL4lPEGEUrChM
/xmi8HxfbH5da7kQEt08CQgXlpuHN9h/s17OtLWEGX1aCr7AFt+zRnWjzotX
UY6BJiG9p6RL25seCSsSLC273MiChl4FEY/eDWg76xDkJeap4zyIFSGGbsEK
hV7pzqY+2TiP14yGzQBY9cdUAEhkKVmy2PoszchggAkLuKSrhPOEzqzCZav4
IvefOQ77ox+YhUFwLKiVEp4IKBPnqJ/fF6QtFN0lcHSjfEmrxXDxkCBeSpBx
09QwWzWCEVHIuahnD8frvNRQy0Oox1t0b8uw8NDxYojFvXRJDgAmcR+oNAay
VpUpaOCLv9rgAS+EkDG7+RHHu7hOzAQviyvVSg6JPPQdGYKqfcbQEslktveV
+JHSmnUZRWGvBo5eS/nyC1/V/XDQgnW6GD2fArGSmvDs9PHZ6I4zY7x0n0E1
Q7GKQ5UismAwQFkObU2GmhuGaozWxt2ggT8jwsb8762Gq3tr0qXBiHq12TRf
h7ytZqBHgiyVydvX6OPHbeyVIe9BlmBqUxwRUurzIPkT3oPQrPZXf+t4jfTq
CMUrtKKWuLZnRsOgIPMVRxojHA7mPHh4sxurFWldToPZdO8mxQni5OFPe6tR
qWxgXUf20i69BXTDTv3vHM9eRBmD9ZGlpHBttuIuOeDKVlzV71lQsA98uDVd
1xPKyMUbokngvMmgbm1cisaIWauMsxCwknI0OYlEnbed7CYhTE/bz3eMG830
E/k9V0eCZYugv4jBWP5wqBT4ZtYI+iWZi3LnCuMfi6AwFUR7d0O5JYP2YU+0
rNfCnF7SEt2A4w2vqxgswS2ILp3RmJKB8BHu8xZVXFcPDPRFvd6jau2FWKaG
zqYdJ+nCHZfAjx7QHXHQjTRgWFFS9iPHJVG41mlOtKR1u0jZnEmU/ytRYQgR
hsBajIdgV79r5hzXNdqZsIS/l4duH/342pfJypuCWPVJT+u8gR5VJ0v+b+4u
R5dZFZjTY0n8m8SFYukMWyZbrDBO1kLJLuSP/829fRQpigCKcxtgIoDi4mPk
fI4BCoTq95zJNuKh2p4MrxEfZjkwtHkOqYWl75wQ7iTQ0qoojWq0efuotyfx
7lQvK+ncyeAs6ViNpjJRsvoyy/ozrGJryVw9F6mfKry7+dKEHykQMcltf21S
PUXi/aByI8LsD4x2Kytv50zmLf9e5rarrnGml7lykBHXv2yXT9OkBB7cpFPn
1xJFkTAocvaKG2pCDJWVcYwXrIeT7UXNT0x6EAYLdaJhKGiVVR0+QzpYfjXp
T8jDEMTPiKYFLInueCf4cfzlCnITvWxN+FYbHKZD96FoYFlCYA6Wjr9f2VNQ
s4DvvsPZMbJyF/g3T7+4N/qV1rJxZR3vZvASPN6AE7r25d7nlPUBUZB4MU83
/JQWpbN4q2SVfokKham9vzWDLDUuUbpxBqNEx+ei+1KjnAwzuDJ9BxKaFeox
gg5aJZ55npwoTzqrtV6KfunsLHS/7mVyzGoNYZdYc7+LfHU6TYtQuP4YHnxw
4lEdBYVNEkPgujCmH73HR+sKofqUqK42YhNqHOANmXORC4/LbQW/BvgIQ4q0
F0ER18Q9chmJyncHMFG3bjWiVgjAL0RTSYo5cZnLWj/abYZr5M4Q6Y86BwMD
9OhX8w4yVIY7PCqQBp2ph4lBqQMcs3bZJvHKvIeN0uj8bRhek66GtNmDwbBb
ECIozA7g0jYp3SUokvz+6pQ9FfxZYOoid9f+abNgZH4l0YF/lI17psbz/aRA
UAfKnw+W6YUFplXsa9pfBoXuhiOZyV2I32OAOyEnPKfBwtShkjyq+LFzw0rA
zrOukhU3z9gctH8k1MUe8zxjunGmY6wGWvCg1aBmFeE5SHsMfZasXYRR/iJM
hsUWdv3+BJshAttsrp8lCHJsa+U1ygeYILrdC5cPwGx1MCf1l4EKaCLEf2kC
tsG5dGe4/QDnduE68kv2wlSwpQmgOTk+es8QaDveEx5JLtgb6f5I6Evl2NLa
xywz4iyPupu7w5RXjG8usftP2OSv6EiUu4/pFT9rSNlvlGE6NWPGQkTlUJN/
Ld8ysoaLiCKDNF49AyrCSqhazMZr/Bb6TvZjjkkhPGnmkrHukCfmwQlebOhr
WJMim/thPBxCHnj/32xOYnm5SMq/kPmHzsYOYgdRQeYixteqy85UKgOqNNAM
BZrEmDdvON3jqs0T10jf/l9oWqweMlEpVBzQVXahWKnv+CBKf7memiEnIlX6
n7VTBq/0oVfYxzsNMp1BIroGQjmLrMmJK+V+EZODVb8cCHL8xQqF5XsdYvVj
dUplpjxLobX2IW5y1DoU/eovNythG5XuPlFG5QaWJri5d4V6sL0kuB6iShXu
0EyU8Tb51qmWMNuTY5jpFGVKH6o3nE/+5r0R5rjiIcBdYv/CY4DLYW5Lbjpr
QGGkm+qyrum1KI4YzbbyyVqw5f2hi38L72IpChZWki9qRydGcHPFaF6Xd3Hl
wPNvB8beZ+y2NzrTwnGzvCsA8uj0gzd+oolYHcTtP0E8OrDaQKSDKF5VXAnj
YNsgnYYTV9UVuOdWoTe130hhBctCmFwKjrD9d2V8gSL32GcfeS4aDjtFARbh
EZpLJmyIiicDmwgGH2n/HWtj75dbjnAt9EjbZKW6jjsZO6CB4vgyMUk/fn7V
tvWdN+iqag5JSq0KtEBue9X6Fgx+LKIMDzU3tUn/2iBfSVHz4T/DB0qNIqZw
41yZ7tYbLS4/pJN9vuuXBkED+Q15OgeulM5dHZ6Ep2k4EGdjQrhjYZUsshAh
zFG1glmsJscqbFPnT/T0R13Rue/lhuGToE4OUBLCZQoFhdpf8EZ7a6ATCpWM
FFCNOQCvgYKeaEH0Npood4uXdqE1q+p7kE3Dp+yu9bxZj3O92VqC+KTGGER4
XPqqLI/NkFnVjmkHUEMkcGM+v0fmdk5mEtCDeGlLF/F6aZth2iaQSWV1CHMT
acoO01axtz/oOqryW+W/GG7ha+70Vcw3Ys7uIx6/APCeSWy7MjPKqu7hOEXb
EHB2Wg8ArHt5WtMnbOTTBi35PmCwKExt23bHwBKU+GvBAfJTVq+sCN7KpQpz
xZNnSCKfkpCZFctvCY/RJjbxR7KOl8rS/OtSiE8UxkljzGabgtLiu5A/yVJC
i+p5VaHqpXa7we8puAeDAkRR+7Q7DEnrf7ImvEdc3GCsWCKY2pahxFRms7IC
8KFgkRFRqX4RI8fZDteTH0jIXkSLiNreXsmPYuJebsWTLstR9bNKC0kq+Gvx
o3TJC6ZyKa8rLvOf2Bs69E1UezDYGxp4+fg4bJ/LcLuyaWawotaG7Gp4IS65
cTPenutEFEWjuPQKery3cL4q4llONespdevUMWOS/07VjPColWhmod90XKB8
j8uNjXBcbbHbjAU2y0yiIpDtUr1eeo96yMo1R8EGBXqmX1svSs1aDvUcYxKd
WSF6Yi3CUH1JPSeW/XuEBHuti7OhfYIxpK/mBDEBiSKWsLiSTiTXyLXoPrvm
vrF4M2jfLYnN7N2F9NGZl1rLju/iKojw9mm6VPlN/GR+Zttw6aaISm9UmmS/
B+rAmNRsntacr9vsZ4mMr7Rro+sH2xnBYpwNiRGgJnm8kBSDmmI3ETLK1VA5
Rbpzxl3SAX3Ow3aSbEiimkG1xgOFYnZTKtNzQixzldAtzuB+lspq4c3HNUwS
DKSABru4r9H1c0Z14JPR0SfOFEe2Rh00DdNSTrvzPYpKkcwUlwCJa1LjyPX5
V5WAzEXJYbQZ3oks7Uk1NZySNn1L4lXE57Gm2chyQfkLC1oYcV3e/9HdomR2
DEi2Q+fF9T1HOj0SWMhxcSvRk7Eu5/txLdLrGAqtgf6w3toka5MlaEwnb9tl
YNUzyYP9Vmg/5IKk7ekN7J/FooKAShTqsqAft2MAypkshmuhfBgjjIDEeNk+
3DStrp98iYpYa+g1cIamQNG2qh5EVF9vvLvAS6Ku0XdWqVPCWN6Fa1j8Y7jt
ju4Yv/LzOIutL6aApw6jGa6zboj9V71P/q8m8a+mNBOfF/wR+kIiTk5mNTTX
QH9J38+mVRdHQ/npTtBZsi84jxEPi+/puvKD1CFyCt5CwIELUFXV/iZ4Cj8H
hbAcFGAGiu61y/E9rFWMYQTkGFs8bIjtmcqMoAlm4heF7RpqNmcNrJXfwgPO
F9kP12qVNPPOsqIiv6d7hvCnNrGZ2qOUVylOx6aOlQCzZ85VodMw+zhmawyE
1i9tqT8KuyoiSdZuTXHX6TEx0sIrZy01g7XkXP1iZNQM1pLl9m2hIWE/wT4q
kNTA6Dv5lkjTb0EsyTmmrZmRllFuS3mcWQ+yNWO21tmktAUP53V3En08/jWO
W7/UML1vt+cLBXewRtqq0pUgEBtVcAR/+febMJKXQ9gwHdirWqxVK6VOtFTA
BdtYRi0qSsscu5Gf2Lwpjl0VI6aws8iNSbVBDE4QGVdlnS7FmPaywX2LUsiT
IUsYu+tVhg4WK7qCgU0QIHPrlsQkJqSCXbvDZ64KKB63QBaa34EH/caylLTy
kylzSI33/9125H70gaJDcqvBVTO7Zj+kdQw3hydAjBTugFBCRj1o0ZDaQXsr
nJab08vhyCk0Lw2eN+GVVKEJUDowINH9dHb6PrJL3NL5mGSI3xZyFdOEnj3r
647Fok5F3ayjIIDek7ahM9hRoMnqVnwUDhkqViKUs8rUaFxAv86No5R0qDv9
ZrbPcC75+iHXwJuULOCHCWpUQuMEZ2BRj8Xeqo3OPNbG+iSWpttNvA1L5uQW
kSY9QNt14PeJU/H7VcjsqbK6c9uZWRpygGnQLw1CHrx+ZlXOjQpzsFIDUPAY
bbXRGXIjBU486KUT+rhDl7rhjbk/rfsvHP+giSiwgHjhF/Cz1Kznf9tPqomv
CZvPQOrd1NKVhh7GpYoNA9Aj03p0kJ1ajkFVeY3kFwX/mQPMcVjjcYEx5oDX
gnkMtpueXb+kRA4mmP4CwaFFCfSbEYMdbba8SinnTQzPNNKmNpusTByvZX4F
4I+X9nhbqgt1M4mDjBLh/A+Py4AUu6dHqggFSSBxW2Ox09OedkrZD6UyJ0kq
9YU0L7bs+HLfuEOlYVANHmeWcZVNDTeXt4GG9TSYXh1AUP3Z6i4JuUxr7ukT
Rhv7BpzbO+yTvAIOttak6Zs28DqmoMDsVajKfb5QPfY3BM9dRKjcAmcmXsuC
AIS3hBYr0MZfGQ8OOyJHf4aye97oNbu6fswnYVgsQjSkXLhqCNN6Gdm/iNpP
gSsEbF9OQdI8gfDaAZ9ZS6fVjvuvUiwnILeOhHfpftO3OclQedoDixh6AVLH
LFxeC8Pv49l/tV5IyZise9vSQlNjxJQ2Ec3aJaz9Az0QFh2LORNGDYVJ1SPc
e9c0AdB+9gK6Yl9XBh/K07EsRr24EJlX8fwvUkPUVdRNXort8hHAIymEOIHV
az2FUFq/zcC74bclm0G7VrkW/iHhcTzmL3HhpTzC3EP3D/Ql72mi7Ew1Ty3Z
2i/54ZsbqbprDOt3j51QeJdExxFskCdvPieo484YJDnAEKZkbzdZr/bjJN3G
xf5/NUCqLwMHiLPVvLrvQ4tW1XfjhDe5Qkrr9JahjxoD5CnQ1v+SOEgBkUTS
HsYuiIhK5t/B/J26hoVqVUHVoni36fdSHYF9jLPFMdiRBdNwTMY/mOlmRLXh
IRp/bLHbLfx4et0vf0j2Waka9aFnNSIOkGQkcHBPBTMv3EIBjr6ATr0/Xeud
32xGXdPJHDNA754qJfcMtJjKcaqAfSwpbtLvs2NK6ln74vUToHNXK5z7QITZ
ZxUdpqLt8qkBFOtLfR3ZlYbUovF4Lx1cRFrTtddnRdS9rDHJ5lWlJGqbeQgH
/OkCsMniZ2v7kpl4yuzMfCOAbrL3KL7KJsYoD3tMkRNjapOLPBb2YZ/vwNoZ
NEEgzEKejFDRp5smQIWZuf69w20DsXwh5dsfFxkzZPAViv5PWog25V7hvRr7
o+33KbR+vvh7fuFKJoLSQdB70GJUacax8Tp5r2QM1KyB4wM93JX0cGxoSRW2
3Dux0U2E1tTz7CrQdCU3fKisDSsQOy1cz5ghg+h35j3jobERJe5bd+LIOqCi
19L9VDr7SNtlrWzA8/Z3PwM7DgknaLik1/4+CFRP/rbVmmavF2f+NqSGNjH6
2dzuf9vjaAx+dGfYVlOpFECIFtDZGIBQsgxBCWzB9TlK/3Oqu309tr328q7p
O+malogUmpAIPkAvzIqjhIZ0vUI7few0HiwL30UBi9f7FGZc7BPL7aECrc77
Ldgycm5P3GeDQhZ0wC9Ejf5M6bBXaHg7bEyChe6GGFIlb0KPli5k5G6O53Z2
ybEekVmysmtT9pH2GD3o8ObxGdnu7ZKfxd2k2tJVPbwmllnp32RGevaBAx1N
82hm0zo/D0MLUWIxV7Yno3fD7DErevYAa+zhv4813oumRAATPXAR6jeKiUmI
VvZDg2yzAFjYqb2ELh63vKbT4UW+T5jqcqqzBAVakqNK1tcpeIAA6EAUVdI6
XmYqW/IZ20cGAEklv9yH6YFf3Ghk/Stm2fcQ7CHOEh490rkYFB9pclaamkGl
DU7LyVzPP69qxl5c2ICQk/aeG/02R72DW4HQnBMpnzOPKnJiJhscRF1sl4/Y
/6PmqcEUAAcPXrr3fTaZsrAqXm7o/BF5/nqJcnUw5tV+gGe2xKtxfnpXOpiE
qsKuyyZd9dbDTkZl7lpafyP5uigi05PY3S7JKccM2sdGSVN6xTaXCpUqwINj
ok72eauzTFS6XP+8Xy4aOIkqdrZDXzCc1ygZ/XxtCOwl+6t4lECJiBIsH0PZ
grD7PeCVx1MY9hMeKzQArHBeltiDm2aZiXVyyWk3BYpAghjEFujNSft90dsY
7FpOTG61CgQA/eBXVy1sSaf93A+jDIuIzqt94ZysxrHK2dLYcMe8mjyfxZVE
ewj3lX0qgADKtrJL3rqXchGHccW7vXWneBlvjVIxPr4FOF1AeedDJo7WCHbn
J1ZnWmDG4mA4jka6u6TySE2YphZZuRr1pvZKThU3VWgERfX3gdhVnLP2koBL
zqnfmYqEBZDOlzX17qJybn4FZ9sTpDBDXtJoAKiNviHeqBDnLLO7PIY32/uE
4iiYLVcbflVXeFzn6fdxXLiolvitbrVfzMzmefcvs7qwVY+i1s162WghQR8c
VNjJnJAjRb76WwssvNW0FIlGWvAWy3odB71DJIA/q5MzYjfYeTVoha/2fV/P
q1dGadq3tht+TXlER6BgBNRrklarndJ+RwLNXxVmOSGlOwu/nhbMDRWndLYU
KfnAb8ghjUua7ecziUDfkWu3wCJd1VpzQT3gjo8Ue45z60IfVjkRxSbztk8M
/W5fnVF05CzYgym+rN9ZjyWZDIfOEG6vqi1tLUqFX7d0c30jQMhbnDZBLVfc
f3esak08EsxRV89jxPtJXDB4ren/XZObbCYrlryZSDkMD7R6sFUtZt4+z2Tf
vdni5ExSRvuvVnTi4rq1xa/QuASlwATfGKYKLuISomlBXgJJVHIa78OYnLys
EV31WsyFPP2cZ78XMmX0ARw4S+GJd/hw/kcbwK6qZEBrVBK3lulzBe6t35sx
WmMAQNX5oSCLgs5pUjG0IUuC0N3iJg+vH3UDCfbRFGtwfn3vCJFRpE8RkwuC
3h3zjINzU4xExUI8iujzuWv0Wyef5MrQ9HUYGfIpRgfkLmcLb8ActESYkkhm
TAPKq0QprOlpne+pMNcasLG71RTgjR/+Ks7q6WDZSGMCBeZFFvD9+EF8v29a
oohi5lb8amNUwZDCICgSUYUOSBZtefwmoEtFRLjl5hqA+FlraMSaAS8eTZE0
9CRCurODzHZp6yAEklG1/itK8oJCSCuGJiKy2Ovg/VYYcj/SYb8E3wkCs4tQ
rXYN2JekCzD8x4p9/CRgnqJ3ugQfR1zJGzRhFKHrfe3CCivBEeCbigwLzX1+
yI2gp9oI8awqiHVyXf4OixCRlijgswckFdzao/NolgfU7+PsoEt9O5r1ZIZg
O0trsotajNf9VCcR6VT2rCEIrntiyAqvQ1y1gqyxYO9w5ScOoLo/3wEyi7ny
6MAL0GDirfI8U981x63WeWZsIffPdC6t/SRjXU/dBRzF642cpYavkqMJ8UzQ
CCcKoYNkmzXhphyFm8IxRwUzysWMyAWcrMlW3vY8cPAsD0GSkPtfKMuPldDj
IfluNeoWfudVjE1J7OedYI97ZgFVCBKWavKVmZ9giA1WIGOQIoeNtn6RSnba
jF09rsmh4Hbkn2GqXzSLKLjFgsB6jakJZi9T+onUroC0jlamc2BBb8GXjJO4
dO7GjiiPZwktQQrKntF6rmujfcXdwGN9XESz6GJWj/WjQFCaIxjOVxzwQohk
EiU5MAj+8roKFOrsJgC6bchJcEUo4JsBIVd2CHCVU/JyyPuYPrF30bCy+R5w
IqGRv3hwAio94bdt/M6rHVwBhSCtQVWmqeGpGW8Fr3vtv2/oGCLa1xR2mRi9
utfzbBlk1cHHbA96NWlJ3sPuqzyxAGB6JvO/rNicL8Rvz5GV5EJi8Qypx3N0
gPUQBiXOWEZ5VRpUIJp/tDbw+CGylZ5Fyi5rgQESf/Cu5AihE3b9qEPoBOLk
g250KcoUebIK5BgYNaSP2ClbdCuVZKX6wzR6hvp2d97ovptVrbUmKP2kFUgg
ockUc1FKmjjd+BJDADhKJZjuJTz9C46U9ic9nk5Qdy5Zbb0aEODc9bWwhQu5
un02BgTnBHVeWfFSIW4+AvFOyZCGdwZMCVPHBJHGUQIQXsDxysmNZLvvUwYg
cMD1o6BcljszoYIi1g1G2KvL+v4FV55jjssslzgPRgr+/iFUY3MMx8KfKtvz
m5S3WoqVtRCEnCfEBwbKdtDP5B4jDQoRwFeMifdCXlDj1sm/pmcel1HpoOf/
5VjYoAp5l9UXLs80bya/nx4ssJbCUiNko0ikq99pdHKP3TIzyw6CLJDsVb6h
1EzzVAfa2BLNuyY28437qSe4Mh5JXUJUtAVq5A6wudwuhvOUYGhQJbiF/EqS
dKdPYQr0ay8AD/tWNoKDXIhE0jgB4UYhO0KBH/Q4O2RwLUN1Rgd6aCA+aLTG
SLk0L4bxvyGUe8ex6Cl9ysK33Y5bIHaPV+l8l0Wwt7PqZb0jLxumppF7NSvQ
plmOW8GuUGCuzrlV0EZx+hN3PqR8Sx4FGNCmtRKTfOfZB0E8RTbrYpPLawUc
zfrkQ8x0CFlDx7XzKmxjJNsdW/OUncH35sYXq16Vxkhd/VRS+Mk/RafD8vxg
5zTGX/0yibqwZ6dkV34DcSbKM8Lc75moZmC4jv5Qx+BT/cgooV5MhUDvh2Mb
FJBycOeGkzzDZvSbRwegUlLwrlZbDHeULgV/Wm3ZfLyBMNLzIk8kPQdS54Te
spty1eqPiepub+4XVONfQT7dM5g0yil/bN2DX2NMpJil4OS8MVkOURsD7R23
xVj/VFQmB4+KhBqml+P8CKG6T6uLy/z07h9jYzfqrnfr2MZ1sNlzw+xtZF1z
tQgFMVNKuAg8Nzgk4iWOoSUvIFCDK5OC4IHbWKnJwc4lM7bDvCGKsPKDQblN
q6WKyIA2TKeXyzjx8eubMYs+iPBtisuQ/XjFcWt6f7sldFNpw0C+4FCB61wx
Lw/x2XCmHGO2wNCKK2Yuznfe9FyXvwGlWLAaVkf3LfQgFKmysWU1WZGYvbED
xMArNTvvGdpbQiG0UefKKwSOaRyBZIzfJhXrqAxhE/nJzwdqAjX491bUp09U
Melx4Shm6c8VVbv+6jyPVALgdB2Hl7CCLXtTF9uF0Rf8qvzAye5J7Li3wgn9
YCateubYGAtNssNWoKh+qrttvwT9aHAu0zyuhfMyY6KQFfNMAvManvVCZp4J
DK9LzxsP+DqXJnMQTtSSQmLMopdg3oz2KSXfUvjgKSHciYF44iDy5zjyYyWR
70+im3UQIags6o7iAAUhQY2/YCFOT6NufT6TNIkagW+IboceBbtja1knkdbd
CGexibZ1XnRhMcOHoAOLF7879dtly4dEUEy2sCSWePPs3RgYyAN2M+kT6XFa
UNn919srffNS+/PvaMEeFifBT334uDWo88uchylTF19ajNHpr9Qva9XtJvPj
Mzx7+HVjAYlODbfQW9sYly/+3e/9PYQN42EI0YdooR+H4MZCrAz2/Zz2dgq+
h23uCGQl/LIYJs/XSBubRhRQaX5LZhu2AxBcx6uAuwcTNKrpIyG0Vgm6VqPA
inKMt66LsETF1ojavg3TznK+VmrYUtK5JcryrDICUzjaWbKGXwotv92OL/Nj
3oD2j1+zmJWhyuDq2CdCUxsqRzC1lYIjg6dk53hQwUJAPAVnedWNxTGpNdsA
MOq+e1K36cEPgNb0YltIFDa3aQLLqakidFWENnWUHE5Xn8qbdLjfcb78DQXM
AY1VY+ROV35mof68+HBTm5ABZ0YmV0hN5KndogTIjFfeLu009fuXvjZIUtg5
k3bhcXKUShOcHCuR2/hoo5HqxIqLfSsvnKHk/uR+XgVpyf+hyZOh/3A5Mzkz
jGPvOQoTa0tXshA1hDvGgJ9d0h8yELWW8MR4eMD7JYFD2X+wR9+4nGvKc0lR
3SPRHiT5+kbKEE47xQ38SwaKgfHA0d+IjbeL+YpwmV0vrshuJMnhlWGp3PHm
sRBUGFpc3PMvmcGHYmG8E3c+3SzV6WMNub+vSWYOcEjZA4xpnKLlr9ks79ab
fxB75AtkmTTWzxXLTU3UUYcdE30nhAoq9xUGT4QncvRgAmdYjwq2o53SfKbe
GPcQxZkKatBgGR2pJX464sNmooiDuhZEtR4zXuZ2ZbvUWCsMJXIF4OS4Ecs3
LKbOv7O7GXYeloR8HbkkNLXKt+lZsagM7CvBaaElgWYX4Gih1e2raMcw0Sya
ZW7ymHR2+sSTZf+Scyzx2KaPzPKgieou7yiu3KV7IiEIw0J8oGyx8yMtdtTX
VWIBnvRbGfgxIZABVBsM97EOaXyia0t5nnw4hMQr3dzdjPjF8m3S0QM06GAT
Vx/RJMR4ojxajNi1Y69vk2uIsJrwn5AFIMMTIubNSZisfcYzpwyaAD1GrY97
EsxCnUDL/IP5tFiREVDwfdAtDS0SqBrBOWNCWx5W7P8W/iYsi2AfBBf6l4mi
vT4xqk+F8JMszfdrly0Pngq0YNgZzwRHMhdWtm8PzMxbZ8lKV0XYmDpSpFYU
mCEwZyUKQo5LL5xW+h4jwIYkN6C9UWfENM03ajrAJfPZd95EtqKkac4HZonb
MJmhi1ufCs04M3cCbqu/a54Vha0VIegehkLK1h0eB97Woz8z/XMydb9+Svi2
uKBDZOehFwIf8/dAjtNia785H/S1rGbX3Y85jFSc9KqvwvZZXdAKPyc4V9KU
9+qca2uVUAos4JoFnotoMSsSRoInQMYnot07DKrPJxRw53hSxst5BeyIFiCg
ro82mLfA8ciWU/Ap3gBTL78vIhavFHTOt/00v1undEZrEKQpD8UJP196X+cu
USximKMze7f3muPmg+ZbDsmyYowFz8eo6JLj3kqGJQndBmv46ewb5aMggZFA
AhNHBu2MjrtRzZDQ0MEuWorQtcj9VssqFMuMEKXWcTHKTbUInTkqW11V6Ruq
0Rx3Gujfgs7zce14qRD9DWFIPgXtEJmKjGB+eUBe1X2+dgOlT/RsGcMpnv/R
wtvhFODBXHlVZwEHFOb9exeK/xMEfdtxLTevctaOB6OgoLhpQoD34lTRNxOl
jBIy/u5jqejf3J0quY3ozQ9u+vrDrUM4mEkSLeMpsP4+tcK8XJt60WXokYB2
ETnWdOrtRx9Cw9pcVruKgAOObSpMCuXC3rvAqeWTdxBhWCkSIDhc/msvfHb2
hFXlrCJL8yH+HsS9XSVV5xtirurmtftQP9rUocv7bN4c7tXmaMjLhgUX/cV7
jRzfT/Ks+XfnNryJsWcF2pyBvylHfzUymo+Llzq/oEupuB4mrS+RT0KWZOF0
2UkExSaVE/wLikUoeO1Qn/7fxWHEHyC1Lpz7mJB3nF60PjN7OKpi+65IM+sq
VD1MOu/BgicG7PDQz+zMU0vLTsuT8oMtX0e/h2xmVcZ2s99UXlwjKtjPtyGE
dD8K6c6JMEP237n5rYVLT8ypdIfPVh1wP4ahojnYCD+6H61Tllah/g7YYG8x
qpfRg/q6LMQqWD2FAQuW30dzGh/taytdBjv3AfvXZoik1kcXY1PiuEzdk0h/
gpzhE73PasBvfYvjaaKXShH/CxevL/Pc8v5nXXyufpxw12rTvVagr7kqGrxY
UNAPQ3R/usScYz+spA6re7THFdTerk5Az4Xl96DkwJogdZAQo3OkfAnKP6e/
tAvH30dVo68euzAYkIUR3RYzjimxNM189H5exSTIS5b4ocfEkXoo+jVp9cij
bCyy1L77MTtT/xqLWgodbg23P64/FJZrrjck5DDTIXE2GPrNPUrie96euKb1
OAjpMxK7UgMO0ZrDz658XiSaCzg/0txc5eumwTo3splBI4BfoDVdccNyQ8NZ
lAX8DDOU8V+qDbVx2gLsShz7EE05JPptJX49HJ2fiG1jP/ZhEBzDDtGMPGYN
MjHPG2KnwmMk6gtQU3Yi+Yxl6gtS/cGEJq1WCqGX5EcgytdQFweNjkNsAdW9
d0uXnkjic6TjP37PUb/vECakTCOzCcaJa7b9p5xrcvVQG7omrvIvo3HGvOHc
QG1ghVGlR3rHmFvbw8HQjgS38g3kj6SSRw3amfwZhZM8wkFueZOLoCIfT3EO
FECJNuX/2RzbSf7dCgRRckLiXSSY25oYgoGRLnV3aGL19p4r8iilSFVCM/8C
dvAIGvOSRgMD9qHjpXfL2t2WZ8EaOP+S4d36YsCvNoCdVU7GWx/0rMJQb9g4
t3/OGvmj8dYIFQ5WLtCPDRplOeTsd39l47Etjvj1UuYoPvPm9/1E+AytY2HW
5zUMZnqA5c8LHJV9JB7KffvgPt7Nfcs8mnymHlFDakXxIOPRAxatdTDRWO2o
xFFVAgt6Snd702ptqTlWcjyhRVpy+DnXLZF7LUFHYt/y0c2BNDFt8PsrTLTD
1RC/81dy+bcMSTx5lUuegNHrRCBsNrgK+nX9vdK30VR8PeAzGh/M9YKPa53K
k08MwM7ypvkQVa11OeIaOsl1lERPObV7yzzV7dObWhx5kLXFL1ss3nVvOW7o
PDwF71+hpom1BzYX6XrD34xa90x9VWV1zvK9BnjWhHjmGu/GnECu4iFEzpJ/
PUxv8Vvn3feEGz21TSXCXQSekmtnW/UCnt1xzVA2iLv/ZaO5oSNa0IvZJToK
/4mRf6WkT0AqQ98WEV6XBjMhjshqGNmFUdy+fVB9pfhCa3xq+pNnDSsb2dvD
YdLHih1gsGfp8QEMui6DUuLAr6ep0GObgKZBdflwo69ZlQTsypvYSsa4UA6u
jXqeyP+bsNFkAKWkYQv9O9e68iNtgSvnHA6cj61Ow5MUVufvVAprZIUfAB3a
/dyg8MnjHvWBm37hSdZMO/cXFqTWE+SHjrOiecumTMuBhB2h1n9WYwKf/z3u
4CtwwB7sna0NTk+0bJyz6uMmZ6abjQ2P2GyTtDkKvLgdNjP1y/WsgfrLKNcS
fGhDC3bv2jYBkg8cQg1hBMsX/70UN63opdBpVKLoku+DDmUuMrRXv5GRkLm4
nBn3j0t3JedPIwZStLVauDtRXUZfKcMFGfdEP7t4rrCmnGcqtbMzp/O0vCf2
jOE1qhz5rbTLQ/1MC49qDrzm7R6Z/Q52OgTRnDaKzYLu01FSaHWpUxJv+Siu
ts8R1JvXWqBrQM+4uvBDol/W13PQtxm5OGb5aRvs4n2qBCPjSD0QtPRs9Gb7
0/ILiz70YIB8tTObVZr/R4pdKRbDX8GMH6FB9dRt420xwW1/22EJPCBk7wbw
/JkeqhLUAH+6NphsgrLNCgmA8OJw0lkycmjzu6LO9QlXYR8rgdmWzIT8GR7q
04nFZaNMbpqi5hcOgdkGaBVhIIrtOhDl9o0vGnBq518XHPAcrq0Dv74cqB/d
FjVMV7Db/or54qM55bhTf+pumrmTrm9KGQIaZoWbDvsvh7hf/uB/wLzGYW0Q
BCil2WReU76vFRq3KZvtig2kJf3TJVBL5q/zzHcJ8CQE5y2Qd6RegLl5qeKj
UT5JWKhrZilASnCemdAoIA5Zx0dIy3PdPMbzBzhtg+rP9VwiBndeAu2y718H
YgjDWHMq9GLoqaw2h/yLipYDKfzaf3BjcMBS4zZqkTPlM5MYoRxNMAW1esOi
n9lYaskmtKMRuadZkA1b6OnWtjFcNYTwkXBfF2v4f3D6XUOWeZK2Qh/1nnjn
/rJcUclPeBtV3ODtRMDI3uyCgPUL0r15Pw+NLCYbtELMkd4Z00Xw7zcmOwzT
zyaOrijdvLU+gtvLKz++e37gD3GV4qPaUxyE/8fkDNZnbg7cFyklzyMijYAe
WmntFsMB/iPGoMo/Va8IGXIBkB0ma/jM7M+rGHYrtj3RRjJ+98+MnD1vRaGr
QIaLOUiAdLfVlIf+fk8O0AF8wS6yBOyhLm2BaayS6P9PzM7Xc4dgqiREFnHK
FbvOPtMkyqyzDvAScoIEOwh0t+r2LwPrIcSqtMxS3lIoEWJ9nYc8OvuzO8wt
a/WtKrNTTTd1KYFZScDqLcdnBW77Kb945hMEdeJuBT40yBf447NfPMXbjzdk
bzQVf3YShf/PyNyIffSs8FgNH47MgJnUiL2vNwKbP7VpKbNa50E5qTyhAkiE
xp9Wf+PIxR4b2/G/njIOUrNI+xRBb54MJKaNnlqnnWnIGs1qvdyxfhCZbLB/
ga6/LQ8EYXhasH0fZ80Bj7yVoQkJwWZPM1/puw6k4nsTyYREdAryzHcioWh6
PiwUKadddd44ktcH8qUROq2emkLCFd7f6REug9RaikemCEAdV+yEeXB/VcJi
HSa4StVOywlBxn4QvNAjOlWap/8SbJYG8zizb8EkY9Xebsyj5yZXbxlC9mf/
gi8yEyIomtpkzHzcKf3jhm33TM9XXD56FRGfdSkbmMcv7QHfqOWmKlYvTQF7
q9bInfq+yI1daQPLP97pjQ8o67uZ3XUiu63MpK05jRzaDHcsfEn0NFOTp5aP
MYeKvKo5gsZc0+tRaYKMMHJpw/JKzhT7FaWziaXRReyO/qhD5wb+GzgoaDgL
SA1Zke+80eB7iiSOCR+4FhgrwAuG15/ynLNbJc46BK1Skm/JXfJ+bZ30D8Yx
JJDZ+Up/r8h8O6wuen+luDOJu6Hy3oVpXwT7lrFkOHdqbYwq+ig4NW2dw+qQ
ubPr7j1Iwjsnit3jtNsMx69P6P8eQXIDtNYEP07GENQALjArm7wIiq5p7Bi1
nY3C99/tcBf9py4Hd+LxcC/Aac73xmW6N14Ftiw8/7XgZrY95zMZC56Ncn2C
QOq0BSUS4C6buzukXUiYVWIaxuEhTuUCbgSzUTEOp8urVx9GZnJ49Sgp+nGr
fhZkgVg2BHmssiEFKPQAFdIrEOik80hQXXB7AWEkbOko6bIc65TZshN4Wdav
GfxKSay5zAGkvMsv8dfUTc6POEwn0ledUEn3AGs7wES91cFk+UsHCyOhpiPF
BlsMwEYnYUb8k0fjwV+hPM1741ZhC7HYC8OjaYGvGXI+aHpCqk40Lx3JHKW/
XxaX8E2BPOJKtwQCqd+TN16K1g0Dci4oKhsuMIpojT55Xt2p+BvGfHjfi3Dk
ZdsTtqPvl4wtjgZWSmM8R9uxV5AU/n8G2dCt/OCQZDydqMNlVhNvB0OzcKzE
5Z1NPWZR2Bn8TZJanrUsMukmcfmu0fs6tuodXGds2PM9sGLJmdkcYRQKPP+M
b4VbZ83B3tBeRlRYZkbhEoGfLjaXhPPQggokUgX/AlebdgFr217um6OqM+za
IVP7WHiEe77b6WQAepTEuid9lcMGRIj5IGxYnThwEdbGnlfOkQJ6B4+U8cut
SdNE6sRA7enWgpSC2LFVeYytuxUZTugRHD1MXPiO/JUNLzJB5hA/rqjBioz5
4dTLBmOM4Chqc7YOcp4LhvLdRs/kXtQwvQMaqdNx9DKpIThomw/4uDQz8y8o
6ZUVKQAhjfNcXrG1Y/PbyufWm5a03af7AIl+zU1L5xd1X0cXLkhxTiMdy1FJ
yDDnWn5JFPIJcRI4/6/egz8JBHGyEPsaWIGpDPgBM9xazJZVUTy89aPMDJq7
rOvaZGfofXvblGyX1VDE/1DBhAoi4nbUkaQvE3nI36VuG2fmXQwKXdYURM6b
RYAcmOwd/SSbo5zVn48B0LCgbsVd0FbtTuoTP6Zw29hOh7TLHX5wXnO42B4+
7W2km2M4s0NH2n6XKhYI9gGUQI0WDiarlcRgZl3hmD83ws7MKftVZ9HvL8WD
zFNqMjkFPgoQMPwVaMaZJLxsT30m5NwzUmKH6r8b493L/1yziGrhMNkPGR4R
63TnXGCfv+wNE5AlXf4l15S5sPbWz06SyhpQ6y4NYQYyIfTN+aBsbsfldUQm
v8ZNAuc6a0Ulxphvghni2+oz6URpqEIKxWeGpSr4E7L95jNh9Nil5sEdvI9n
ng/HVc8Dy4KcGNq9AOm+YJAWYpDkCXZZpijAvpaarocIchzTam9i8FXo+E/q
fLfNqbwP3ae0queOHY4ek2Axr+frwMD15MJUOQcw2Ak2iqyKRGHx9ASISLqy
5uUQCPOobYkzSInoJmgMeTz78MwMDxh1aDYVKS0UPZydnB8YeYwX8TKebIki
fu7RVi6xgkLio+yAhQj9KnW6kUlZLV5qFpHv/OmfBNtneeTbaVeg2MXsxrrv
A1hBvQUrUFu9hHBKUNJPIaUHUHp5TFzckFq1UZVrlZoh1qaSeHzKarw8f3JB
GCKpuM8OJjTSrainNZMSaIzO4E6cGhi+zDe32CwxuOU/Tv+L6tiFddJ+Hpyc
l6mTjsIWEjJ4rUCFuFCexsMq+Wpvj/vB64ye8nWge/nC7tsJTuUxQxKnAXUC
zTVS41pOiMd2x3Bq8ARsJmu4aAh/07boIykAglZAr1sL+19oKlAQo/zmRfjx
hMPayKbGzdxOc89P3kOUFTwz+9BvMvzGbikeMinecZzYG9GA32GUQw/d97UY
yuGdGBZI/JPmJLlhZ7sKaY3JmNkVQXSDfiLxpGX1ztOogOZjEbT+0EdFZzQv
dLcbFRqAOwPmOkDjT/fVujXDaFLhYKfKhfsxAC0VXDe60O7hLO7DvwfKi7AT
OAWUAAU0kpOM6KnJ3kCMX35io7F+91gHByFEhcXzNPijX/i7KJPdz5tU3YGw
QVrijeAGBFUjGv2opGRYmAqNNnaZz0d80VsKSDzu9yLIJXTQOEp45hpWqrh1
4tszLG60n1Tdh8qH4yxjFRsxQKVU+INDc3xbkjlZram/pCkhc56pQ0y/wHSA
/4jI+vPQ30pP1qljeEja86jMx4fe2p+zqb19EJYzCRJFso6o7wBoiOk7FRIe
d8yeGIwr6+ulM6WW1Hk8TpEXVvXVWB1eIDvcXAvGGfKePGBJB6OMKmpAtxsN
fX3683pgj6GRbMSjCJUkJt9G1yDwwJqbudpQwSg36AxHS/s/EE9L1OlFbk4I
qMT4rg6nogy2JLyG0CTWAJKXfu0+pOoNVljoqLZJkX7J38qrDQ6DUrMuUC6V
PdmBPxu6rpnmWSkqRz98Ms2qiH/icO1UblMZx/J7F6siVum/40lauZlJqwkG
W4b2/FJPnsOFQFNDl/b1edCqVdugNHfsEzFfPtqDoU5RjI/s8Og4tzfPC6ff
cfgDW1flwuyk/Ia28Tt+/22YhSvWO6AGbhvFOeJOeb/cChLYfdB90pv1p2RJ
IUrp3WM+BuLad9IQRCWhf5Gibbgerr3eIxo0dQsTVSXIYZh4iBxGgKorWf4t
7wJoAKpjeFCkm5GsKSUeOZs5yAH/9vdb889sYFy1Bbs9Pu2a5CG3c8A3ju7w
9du40DJu/4WkRZy28BuZznvWddXDrunWmqqr/K+sHTHAXx4C3fM5Da/lmofk
3cykzPiXV67Xrj64s/ytnkRjCY6oJ6nvrPZJ7XIy8Ml52h5WwhmxaGs351fY
/d4GM9X/867BVAtxLXfmjR4SUUqFINossVJvW7OqvSLDBHj9zi7emSKXhddb
ZuqFt3EhTJjj6unDbd2GAjpZnzk57itzH5H0/K7oUYyUP1VK3aS7j2Itm0BF
UR1el0zrv95jrNepKcC9oWkgBhWpLbjgyh72qoItgKaQ8yIvmbj7Fi6hElg4
OIZvv2O+lh9PK0o5k+N8dnbecNy+k4EBzqtFs1iznxaFKCS89+wdF11VEf6/
KybR1vXDvvp0Bz/f9jKTrANY2tLEM8Z/zmvN7POzbVailOPF0tx97YtFWj5f
WmSzRrxqOZ6Hy7dJRotjQccZNp810FoB4wNnkL23Fha7aw+7e9iamjB3I2hY
l87jorGh69QrB24e6sCAQUeOv+7uv2JfAtQl6nwqZe2GnJxPitha6qTzrNwu
EQJYOJ1blGFZNedVLRjWyBKOW/nS4wwio8jxL/CQgqQU5TFk5cR6PohFpkm+
z0FxTj2FTlWN6e3XhDqRiCCKKz3FlGtRrJNp5SRIc2As48dLwCWxlrM3T622
u/86dg5t2xLafTxh59Px1VhuqKvED3LKMSVmxplkaZhVtYlk2JmUFr2z2ebI
HMmfZjiinGVWntDoe5r50doG7HytKeqSVEgIAP/9pmWZyQVbUXeCwOJu42Zv
FeQt5rYiquIkzcrUazcTJcF0MWZauWvX1XvrmeRrVD9G2XoD4ltBq1GN84Z3
CoWUBk8w6cpKc1cRZt+D6NEs40enQRwmASPuIUDJpZvtDyctuNTjc1FDAj8C
GPzn7pKL6klxueEnmb1VGmFJeEPVUcSVu43uxFRFBxR1daAs+93yrcZynEi3
Aqz7rl0WiSkYnScQK5WUVfElQAcVsHVkxFHMImeRM9tzAIDkF+MULUtOEwNF
j2nD8+RQHTGWVcH0gllfmpv04AW3HrVADo4c4yB/cWYo9CD4aJ8D/dJVOd0c
+LlTnGsJHXbhqapRkrQdeUU4ycoHovVaPXt83RQqupLFSR7EIHPAd4CJpnH9
/oN5nFhy21263am/DenOz04VYLOSB0gxbzNvjp4KIGaSAQ/UkClWGghb8frN
HSZaLqCJbZtZxe6KXa7TYp/+r8qM3FaTAZUq6/FMLf2HZjy5rgLY1O+a4Ebf
2rbJBjwhFJoRkGa9aBe+9i5tntPXs7uxRB2vpjWV7DQ+eRYiLi06jIkLDqel
Jxw8EHxlQv3t6SP2CLpkg1NGQopht1XEzFxWjjCkMj2HBfQpvVIPQ5KnixJV
5ysekxzPCZhUjilZQCTutIWQlLbjRVN5YLeNiMDyVgEIT5YS8B+PMBxHSM3c
JCjvw+eyQ8pd3KA+CPg1BoI2CCBHV7/5D9cwN7q0h2DGYbE9B4ZS0ARK3qP+
lhounRCX/d3/4uJucWxHWqGvv+jTBE0YHHNyFvaKGY2HVAmDbcWFUdK7k0T/
CpRyn1da0yngPGiWDXHTf3A9WKYP9TqqUj7Qcvu+V1Wk66k9FAFz2ekD0vLE
ZJwnbSsntOQbg6u933j/R+QGtsgwGQ6v6oy8o4ksqfNc+OpQM+Zw9CETUN3O
+exYa/adIDPqEFmP9HmhypGyU1wicLCg5kPFepQ6N8b4Stg3y3M/S/GTQIqt
tu0uZ46WBXZCS6cIu2z96ACsIEicYkr/a6931FoPBZPT7kpAcEl0+PltpCcC
CNefHDqBKM67BlA9x2s32fXwnEug3zuVvGp/XNViWeWtrX9Z0y7PEdr8qLoV
BI4Rs2uVjU1xfAj/Uc7OCxve5EibBLqxDDWb42p3yp651Iaa+1r5am+GtXnw
U3XtUMW2wUznEzX97QSYeA+5l+2juPgckAbpsWNi8URUQsAYGzQaOqr3Q15p
Sj9MH7odGR2QOaUOLmWEdu+B6eUO1Erz6/0N2rmJpsTEjwamWUcOfVpnrsQb
XTyDhUcrx7CrgI7dk/KW95G/taRVBcddGJjzP4EFyEl1iPsvJiMnb4AHGFBO
ARkjZU3Ga1T7VAXu0JI7jmWTYa8LTfcYlyTqRmLXhLUc4YMjHDl9dQihoqv+
5uU2PJsI35m2HcG7IYkYqTLZ2y36qepOY8vejt26U9HFiWMwweIU16zRAuGU
lUdh9Fd63I4WpxQJaDWWr5KVXOPy0qWDimuvmRhWgUe7pz5ENvOFuDsK6sLC
b+UxqOL4cERlprJ8YaD8A/3Yx6o8KkA7qcpkFamC8PMu4ecrqkr37/KN9DMi
cPUUstxOsdyu8E5lDdmCXGErmL5kn8aTUbDswgC/G9xQR35YlzkITD8Tf/+7
O3/2kDDLbaxDfkvfafcNPPCooKyZz35INKEBALerMobyRI99KHiV6DmAy50z
dOjmou9/MHAfRmIG6ZHUY7gfI0b/TTO2FJDJzWJr284Yw/VENmVXLM42xz9x
pwwP0d7bRwWZcxo7Ib+H7F4vbQsJmcJWC1Ob3ZZl/59Nfajnb3WAVkvqg4zW
giGhyjzZnxxiIviqRVOzR0/G1W5kCp4emPIYahWdP/sBOnUJ7U/lnR4C2xas
+r3B1pDu6HEVP4iLKj6vM6bCsYJ7+B5eJRWVWmeZzhEpZAysg9jB0XHEB6BD
qEBueUd/SAoESKpcX+TNOvi4pM7sm4SSUudH0sWhU9BSrTJMRCztraCLlxKk
l0hP1xcdiXvmqb6wph0sEOAQ7x/0fSUPJll3sqUo0S7vxJhEiAHvfEst6yr/
k9lAEwE3LvLvVz9CuNvWcriAuMBnB3Ibia6zYXgTExesf2fyFY+zebOCFlrW
oxdL+1dn4HuydQgStflaw8CNqZE5o98Hz8tsohV4kiW1bedFgNf6SwcdRi2W
Xkvi14ujWCkRJ8OR1V77VHeeLUopzTNllu9dR2RARFhmwwnXEQ3pRHJ3PiJx
7h439IyJxhEI3TRAiV05JqOOW9I+O5kTnoBF02ffq/CKZY19n+4mwIZenjVs
aa6F2d8wmgDUkJWuHIiyL0EHWVGNUheeH3Az2wWGAM/IskT9Pm8KhzWG418g
0vzapBmmX+MgW4Dqjjy6ZiU+4D6qR1t4mQlhrArwb+BO596cdJ7QFbvrdHFU
E1QChXWp4jhdS9HTbWmP5Rnq33oA9A6ATFRMpe+6Bd9VLYyDPRt1ohvZroIj
8yEeY5eV0ldUb+SSmdxPsWDymvDO7h5O/mWVUuxDGfpUr30Qaz/WZr9Mjly/
VqBgvTfZUWTKux5ipSVOtugPHY3oTPom0MvKXhlTwMkNu+mS/HzFjcbhSYKT
nqVyPQNWBbDUTQczu+5Y5rICamP8cdZsIjhb9dOWLjC1C1WMaUHy9Msawhct
v8UVle4BpYAM+wQ1RWDbriUyJrmgGiBEkgBc6CNX05Q9Atx8qIYrRAyopIWJ
7BS+bD5wZ5Tea329gkCNhqVc7tkTdm7pXvTQFM8iE+9ysn2GOgTjsyqcw+3e
++gO+L962oC4P4GEQ0C3WJhPCN9rv45lOeDavev+eOCIY2u1WfpcK0tfY8ij
5VQW0mZaqxjcMEEQD2e6klGG+2sqLvb95c9GiYAaFzLhB7WEK3WIOrZVex7u
qJQ4lfv5CFRUipcc/o9pxU9eG1qAxpiTMkYh1fcJKb06wt2RRm/2KPBuyqst
mNKEhI0GQ/cmH/EvuDop+AS8TFLEdygapREitaul1a9lLnZJsaUNhYprhJTM
OUpxDfzU4IYdimvyeMX2CfhNljsCbfRWrr3/d9AUVBYGnjhFXopzLSXwJdoj
XaZbUWS+0WXBpZwXUbIjJMI6Ibvxl7xSDFQOTTPu0UgCguJ7jjRPEy5F9K+q
kEpo5vHlRnZAILp72Tajz9lrMspp4GLK0ZDlBRCYYCzZ2ZWyKquJpts6oVui
87INIMv4ioFxFoNJIJ6ZQV08b6rFPES725yZmuW+uArxSBg6EEegOguxWaXa
cXDZvNSCHw7tHIa3t9XoNsJIzFa/R5Jxw4Lbnk/bGLGIGg/hZXCcIxbVRznD
QJ41gEM4lyjhFbtjnES45cdgnSdH9QT1Uk4Ot6yyhaIIdQbJaRwfv9IAEa1u
cAS9Qv7ZSYdWyTxFm3AND8PlBrA0VWD8xFwg5JXS/yVe7XjnBBXXVpHigVks
HZ8NS/a/NBm+bfjmnAS5xS3XosSsGbNsEIJh23E6lA/qVD2TWOqB/q1Dac0c
atSfCSdzc1D+8+e0zHktrtzgS54tWG5DJKu2Wi0vRwYN8qfd+HwDCv2I8+jl
eYKlFhRM6I7ExAfc/47Tar+WZgXFlW1SxQ/ZmYkliAO5fvsbN8EN2NUac+xc
UjCzPtZjkJMr5Iu4EFcv6RU5hkJ++l41FCqFwphLCIyNQcdxWOI2eKq0DPVy
R3+keNku9xkzxr00gjbtKQrWl54Jkgs6zblMwEpXv3LUrmPMYGhYA/aX6OvI
8xHtjdNhHyuXjnnjZztXJzrSv24IZb56ybhHdnFG/C9atqpMcpSAwGCfRYmG
BBWrwzR4jdVCglx0uCfnkWyEUGQuLIOLWivF0MHZBeTH4rEGFv3B/EciT4aR
JlIVeZnYjyzMKEz+zi43XqH3/0T5YlMPKVvgRaRhNXWGfloHPQPJELavz7zZ
p9NSn8UpY2bwGvfdwBk3RQx+YdP0bHLXrtH6Q1i6DcvTObQBLO0KcNPqGjHf
l+8n/psWCJsBu9EphlijwGHgelSV0IJPS0FgRkqJEKWTalnxFgOEenz3i8YZ
InFsBg/HM3xmSm1zXYlQUk+VXoxKV87s+yaf29G81M24+G1/5GdZ1B6QypxI
YA5+7BQiI8zcsAzn26rQXGMrzwJtmR2m0Aiw8Y5krZyvj1ygyiCXKYMeX5CJ
WYypHtKBk9HNdel6rHzTBq3RbpHC+8ZmX94mLDTyQFDjlOoSqOL3b6FXk8N+
20YkppIp/7NYl8T91Ct10M0iUH8si7rAQwGXMcTbPyDNfEVAVOvwUVNGsvbt
CptOCaYEtF5jG9kWJk74zNFbUV1eO3y5C4DRsBPdrFW6XXTWBdAJgsPqeDb7
e9LcA96sY3+mPah8NiWFgxviFpJ87RZjmu9BS8b/+3B1gaWBp/hv6HY5qH6e
lWJ+NQEzRVdS/OvIoGuUBoonxMcpueN3AWwbMbYX50hoiQY8YMpgsltFpk9h
c5fCyTVSEP0W0hlIFY37sVbbj3HvkzCoZGGTDKLA1yV/A7J1t5fOU5UfsAk9
xHS6/HMSJHxbEhJ9n9K/1mRR5n++ZcUCDNnUbm24OB5JpgxXcDKUr8EuTLxV
0odqdV32O9fT9otLzbtJMwIVsNjnhhOo6VJFDW8tLN3b7mwGdjO5cv0kTUaY
CZxf0jeYeN9lwAEsos5FeeMvMOHBsTXHTeky8E3NgPLPpVIq20v4pnNMuRNA
j3V5nZlc+in9VBXsX9ou7j6O1KP7V0343mlEEkT7Rdmuldz0cDsiqvGN5iW5
qawBXO0wb8kS8DLlrFrkAofUdwESoup4Hz4fKLUJsZsbbsiPayc2rCTJlrdO
ITwRPbxBUagT1K1qxqF0C8shmWKWTwIp2l17qihj38O7CumeRRBiWGoY3Bbo
LJjsbU4c8elp872ds38P7XXXG+ZNuha1wpZDEDUJLFVYdj8I+sFe4p9uqtuN
DTbq7aRjMrDsjL3PsbzHB8FaEllVEKPAt+HYeO+sFkMXXFPLHzlJXHxIfRgp
0wXlttUjvauPIKGm/8NkH8jnENaENmrZcGyjswrqm/iERGdnLOwgGT+tLxF9
4heN2aCn98xgKDKTGz58VoT8kI8CMH8tQluHMMXCTYBkpHU+0Ag7yAq9NTxi
qBLAElVfC2lsPHinGaWCQT1HynGggls4W/D2T8SNmWNCNlEYPmvHKxskvZ0o
btffCbiUPsKsJQtSfODRWrqaJuXt5nKu2TUNhijxAZy/Q2MBD4ok4QWZBo4n
QDZMFeJHRTZja8AUJc9JZ9qxpugEbyDqLcrlRecoAudH9u2rodpfMFgfbU4R
R3Zv8s5n+S6ber9oev9/lM0cpbxucsBDeyozh0G7AvXHvFFoa7Pka4mfCotI
qBX1czGfHcxmbGzzreClGY/PTx4HVwusQfye7jSYBP59Qo6pWceHs54RZLBU
UZUvkccBrq9HJKGukMZTmGE14heQRk38W6qUECz93yxAsKS/90JDRqKv7ltT
CK3Mjnc8L0x2bp2bTaljIvSBN3TyZZdCLdC1/xheRzOeylZ6yXGPrTM4ytb+
S/TYLVu3sJJN/qnZh92JR8YUNi1YtBuBFHnGZnpYSTsHBqwIZMkhvl0yb48o
9txaTHqQDwhgTz3SpGwouOyP31l63cTWnM8GWQowBsmTiORc/R9y+kkg183I
e58wFs6GTxeMi6fGg1vSzs3jd/Tj430PSiJLj8KSqyxnjFRl5BD1a9Hah2j1
4SYBYJJ7NoR4xoEbP+DJ2xShPOkdA4AjNWhGoHyjq14HiyoY1ivDBE73x6h7
H0F3n7yYdjqna2WOv93IyCyvf7rxFJcpiVbrVfUA6ORfNUXzUxGdaaF0C4tp
mLrJWtVu/ykpBh2+NuXP7geQG8IyEfn8tL1eVmZRDtNdmmxWWN4Lr6rqXEn+
6DeJGWr0rKVm+0GdVuFXeojHvMs7MRz2YUMFZlBBbHivV7hOO8K49xjCifRu
J8mYRdffCSz4dshXXuIC3SUJS94KzEO59jtsV0nC3WURncKLBfIDTBmIfKJL
MR/3NpmGCk0ythgdvwACCNIOh/J7Ooh3qqyFCMNCtI9rjU7lP6MxTYFb+6ww
Olzu0rMrn5c8wHoWEHY6wp281VPWZp65QIqwcNpgtsUVZUKKCiBxMM2G4YCo
ua3RFFKugsm7fE6sZgXV/B0CdPu1ptfcOgWKulso/eLrwFDgaVMyiCTBtqqB
Zsisvn5C6cBKSssyhMWU+nBg3FzmylQZsLPOFaFM90p1emY8WLhJ4E2A1QoO
QpaHVBxWlpoZ3GT7FM+wkHs+ecpi2gD8rMTcCxvJTd9gmcMehFtJiWOf5Lic
3lw3e2bZBL6sTJsIAoQVnFUUgzCmuI5nNeG1Mr3/3ZzT/PfY+KJxO+9nrw1a
fkUK/Im369rTWcO+trFzb5DFgTgzzCo9s4E9KOh6aLpNBqYSSY9ioHrV1bUs
1iRRV4AEdy7Og9yFdAsxtz8Cwoy8XhnqLCe60t4OgX5fM+GdBrqACrXBpXNO
4s43QZQd4MOVOzUT15Urdn3mABehtK6f/5RvmIMGKi9VV9ky5i/P9J/rAhY2
TsBEI/6B2/hQnxWBYeRvbKY9bBbXgmBVivOm3dfbCpx+Ze8Bcv5Sa5ybmW+K
YnXpAydcTJqtsvMydfBgCFSa9QuNfRzn17fsvmSykQJvn5wFTm0rQfd/iWjV
UVpGYNeQQb2M/EEqCJB+ifrzshJ08uFjylzGhOh5b3b9pRFT6HhSFE8X+7WK
jfYZ8ZWaa1J9hDKRDMF4AdJ4IgDYtN/+6ZSAn29/WV7WHqgMe04csiZIOvlf
WY/VIa+kR04jtbn4emKFAW9+IblEy6NFITw62KYaoe09G9Wci63jMot61ZfX
Ay/qlOdsG0fceGS6tLt/YlI2q6c1q3LquMdE3R89IrZxsJsX5A/TVJEFnR8d
N7+8/QO78HThuZbMWqo1kqUJyz9fkefhsFEj8oGpACT9fi4abG/4AynvdNVu
3P8aAayMMPq9jqc94Cntb9VTqTL7rdf95WVOFMfwp72Whu+mUDwHH2zRIfLN
e0B37lLoMAs7SbL0GBGJxVZ6qI/2cSlmlgwsLxZrF53GrXHtohKufq8SXsJY
ksEF0pDOmvykFl3cRCVsGNH0N/qwuYuILuGDMiu7MKQgO0MakOb/vDrm+3dO
bMMAF+Rwglq9HdEfU6/UpzNQSXlW6JvwvV+nok4S0tSxgsH6zlgB29lctvYz
wgrK8EJP4pOHs/V8zUmnDa7R1tVC6FJ/zRqtGr2J3mSrbDfNfSCDDRBfhcp7
S+oTkUBMiBV2r9WqSCGyEEpNGfOY8KvJ4NPP2lR5AeV4zv5IqLKytEXGf2Sv
z0pVJ90h7PbzFqJxjDI7+Hi2oaCVHyGWUKByxOWWTxt9wqalRox/Qv1JSHzk
qAXEBpz04v12DkukA7CoSuhS1MZIIQK/TiPCyRYRstk1ep3GjKys4PBt6sh3
ayBAiZmZCI7T/KK0GgO/B0SW2Wis+2GT5pKO7ZrJqkTMujA4SE29gzYBfDYY
WZmlf+LL2KqEgygzcZX/wFq8xJj0sS7IPqE8QDT+Ry/MNAnbXdsUzQAjq2wZ
3pJXnou4mK2oDvDrS6oGMmsKnSCk8Q6JtJfP8WTrdGfAgXqbafez0EPhoEDf
96eRNHipR50y41MMW3gmdHEUIouZM/ABYFr34P4+8bgwebtw9oDcdglWNYj1
wyTSO3dSV2cUh2/3N36rgFpgzBMtBFCMjsPRlq4isPzPqkPXbV0JYS5jG7EN
XidahF90zr/EPfxq1Ut3CCvJV2E+pyhMAeflEt0ahXhDmtGMIvkAatkMqLQi
xqCvDwiPA1SJmsa4bDjPpCw1Gidt/XLQ1CY7sUrRH8sXKn6SyH2zDfZTRABL
/gXB2hVhZhsjrKvjc/5GJDouPBCRUqAaXiO2fEdD4//awNIiShZryXiAogMI
IL2wVUftoesHcDhZUTIRT27Dk92IX3G63VvjNPUkrx9iACoK9GZFGBl3lRsh
ffatEmJPJgBb0AvsEJ+u5UGpZkgv6aNF9DOpM6J8XT9erbiaDYPgrqkAorWR
6xNxVTS5d3fegELEL9e/w8t8w7v4E8Fdok1I955TN87tFWeiou4/ooOnuvdQ
eH1s2yITYGrZIgcp66SaMFBQdYJxZNoMDVWyd6eYffUVSkxgx6YZLRlhyiSb
PJXPOvYxC1nHEq2A+alIMFSm1zs4DaTC9Xb6ytA45Xs7DxnzU1T6cXwcfuw4
qQ7pxqUzhJx0qxjK8N8/eYqJ/G0y+iHHwtJ6Et/NVVeNTytTmtS1WsKq2SQr
B2Cxz9m6ZoVsPJwHp+aEIFFPbQJ7MXRAV3lbItNHrUhiUG/Pf77kmNJf5et/
ikilJ1kaVNy6N+XwO/4BnT8rQJnO8S9CPio/S8VPUZH2HncAmKDqV9jznmIq
8qyCrW00GXtIlTMI67+0w2WvpyfU0ckc04X9DS7TtH73rGPrT7N4I0xuhQZ4
GoiCbF6PL1DUp7knUOjbf4nesfSaQp/ejJhfj9uzXWZFLQiVGh2O9THvpZ2m
xXnZT1QmL07c75/2K5LCXIa7peZkuD0hecwL2a+BZTX2c2q2GRRb6xGr4tNu
NdIfLHmvi+JFUBHF8ShiV/RuravytGnyhlOJpUlVWtjbaj9VsNp2weRUyz3M
DSiv2U/1nfClXJ8Q991/rdhod+UlSabE1/q6Ttsg37DHpLkHS61bhqK73HR0
Ez+S39BDFFAq+uxkeFeBCYR2xSVAxjGZHchj5RcHVDN1CUxiQeiWn/kazWzU
QQMSc6cog1gpEJrXNS3VZmaxyrD4WMwUbxXERp3bn3PjK0AZtPQKEw13oUNh
yzkzGPDpCXIucwya8PRsZQRl74XSqlVC8sqqCTycsQ7uGq6bPHkJMfoW1VI4
zaMo+RX0hCB63Ezyt/+5h0a2QhxYYMwn7Kb6+6hrMdli/Lr4k03tZsKwNVA+
Gqd7kgTzjg3OY4eAUxYBKDRxf1eqn64eidoOv2cnVzg5bTenqcBKAuXNlXLA
z3dAB2TFpMVRFaFO83h5UlqGW+EQ+17GTb4LLjbIJAXEXpsI9SQ4YIHWGNbB
RCBuydJerSzdIriNYWBYcgbyzIJoS48Ukt9kiP7gRTz6pN3Fc9PsfkWfbwao
C8G0lC354AL/iaeCb9dMoqQ1EKjx95zGNhgggUX8nzl9Ft31ccZyidch3v4n
pDvAQM4DcLKcemeX7+5X2mdLks/WGvtbJg0qNBVngnFV4WcERWpnzFPPaVD3
FeJ5YLoNcChZEHPAMOog6M/7tqKoor4/bAkoPaRsXLRZ5K8Dj69BofyFe2wD
sK/2XMpHRMt5YRDsTSXEPxn1PBC7mWBe35Xfi6QC3CqWOqZ/88fCuoSg/xqs
/rbnJigCU7V+CYr/vck4CgMIGUxA+n/53BJoBkWPIieRWr9DUpyzknKBGTrR
HeLwd8bzOjKSpKC7vMxt+YyI+oP9D4yJL6RAO+hK3GvI7BgcPftZES7rRB5+
tU7dAgUuCs/aPFMCUwKisnkkBH+eJqOr/+seQ3g9CgjkJL6k6QtolrXSIO5E
iu3/knKI6deO/gf6/5YcnsAUEWMhw0bsh3A72TUIpgWmlA5ZTVKUUIfCdaaF
RqqdFHbBSJbRWm3TUfYhiO/x2GZ+2H3xT51h+5Q8o8Py6BHcOyoKx91PYgvf
T7UIro3gqy23vAE2M5wbRXJU/Ynxsmjbm5dD5UXV1c/apaTSBmBfwFJ2EQpX
OEVNu5Ny37v3hDklfSz01wpuL/tS3a31Ov3i2wWCK1/+TAdhls3aiFXUTODA
3sLJ6thuNgcbPrVy7uSRgzWNvAYcEDJCO4467dMrPtVHyNYENLNaFcMteBLV
79XUfywkqOHaRg2zqWuWfI5MJKToB4wiFp3/NAZ/QHuAM4ygRfvub/H9mx50
gAwhRqrVLoYGL1EP3ij/86XPZ3XicxbnnAdBRXvGxyIySCOPluOIHhasBIop
rmRpnkBhkdgOTKOjJ80mxwD+lEbisXNLbE0545OmlGTHGaFH4Yy4KirYqaOw
ZkitWitkwfL/ha0waOh14W7UT4FgkRbQ4+VwUkfWvIRzoIzZY6ya2o1zNYDl
FExBWuen94EL94BKR3L4cw+cFsifAgag1gKS49xWGW+2wmZQ3IiKmZuh3Xhv
Th7wsIEXYa6yBa1fOuxug46d36Fql7gjyIhMM0hYhaSy6HC97RAVKq87B1Zz
K7nMenuRzF7uIbdYfdf+DxzhULwWAKPO2uzv40ALj1yR0rZmTGlFWl7K/hQP
4up0S20HDFDA15Gv/ckUNXdCsInXOOIcBb5EGcVsUgrwtT+MMvzb6H7+M3r8
FtN6ln7jrnki0Ztt1rPcSGZ30ORWgiOzMSe8W73MRqaFAiccRU7ubDeYHcyW
mrvcBqvaw//HTk5XtvcLzYxurJgU4KclWEfCibgtzxkwsLetkB+bTO1LVw2K
gjmZ/2bbk/Hv2EB2E2UAID5CbTo+eFzRUzlv6LOPqIDfWBmaRClQ6FptTwe1
Yy6jyFTooD3LB9l43nsafZUaB0jwMXGWhMoGjp5MYVLijGyt40YGt8G7ZNPN
8tPw65Hy7qCBW++uh5YsAOzdh3758zBrqTBIw9+FJ1XEXaMykA0t60lpKhT0
MbTOmw+OtGA3k+wF9LDCa2hmnLsj0juVOLqan/Zh5AI1T1HpGtwRgnFm3U5j
TWTV+rYGmJ3eFKtBJG89+YyTt6JueYh7ynWJ5tN57t14RoT7nebat8mGU+Ha
2FaBYA+Cjda1wKoqgX73ZBXPyI71tFTmz2EjjlYSsrcXbcSPDp34KwSasx/y
ni6zV9bTwMkMv26Oz5Zo7THbMlzDkp/Iu/OrfubGKrT419WOxyWqCubaHw8l
+mXy1FU94PCNNbsz7dHAI1rHrPlTeClNd9Of6EZNEuLCPmfo3iqKp/LEnwOP
4sYS9Rvh1N+bZIiZXd+VvFi5h7H8ixbuYApll9Fy1Kidbkc4h2h0F46+cLip
hEX873xYaw56kcTLH5fkzY3NGNE1VRxPPlLxjgbEohZ66pgAkhdnzpvFWoEp
mfB3Xi3fmdaImCf0xxbIN606fVnDPz5veu9Z+VQ31RL6a5mrG+5wel5guh7a
9yDuGT2fJRf3+dCWJYjKM21fUecMIjPoP4Qw1oOfHJn3un3PwWevA+PUzR2N
L6LqflczFfIQs9HrJLF4o0rRMRVivy0QkR5BIyDhlptg1UFbIXngDjZZ06Lk
xtA+kMusMJXWjmO4aGDeI7uAkyorsCbgIEHC/RIszMXvuKZDuVLlQfRuZDV2
3mQ6ONx5zDLWXttyP7YREcg36z73RF6381F2/imBtVvn9kKaTNgGygvnEdZN
ujZ0WDSCpZAlkfsIWNbUTa54H4PvPpWtgiBOmSxtwF8h5vs5OVmkeMQlBdaV
erNhSH4nofLDLHi0ga4U3GM/JgQPxj3WvDwB+SJLvxy9Fp8Anvy8Xf+opbGI
ZFIpzI5DMvVp7KmUJ8PekPXxVrdDS0K36vHrOmvSTbUEd/Wf4ahzzcHVVT8o
/sl3zPL5qrpjtwE2sarawbH8ch9wtINRRqmrQHdncL4Betl313qvBeCCBlbk
Ur91WAsH0hq7RzWeUu3H+r6fNQj/6OeeAKVs5eQOVfU1GjUpAQro+q3tl+3f
OxtLiZvNf6MJdH59Qv3aoZJ9xqHSPJ25hIHs7skDtLuNu5PTo5hyarl/YYSC
9sZELhrwmAar2zSv9WLPBB/0WDsWwpCcs0PRcmw6OiRLIDksJdrC6YTUncRL
b/Quo/s6ny49XoC7a/Nef9UXNLZ4I6e07Hb/46csuRZSHEg+H2+o2gE0jEXR
m+EKAeL7h/Oku2VSbLh20DiHigBjRxczhmKGJA9vE1YJEXbprpm2SGeZtC1u
oK6zzr00JtIP2vY5KOkRPUZmWNjaOd66+q/Sar/sGGtdLT8oTMwYqbHVNeUw
wgsIAGc3XtliR47gB/9zeialMWqlhB4jVAIwEdUGP7ncVuPshqnNxfrcj5Tn
ZYz4Zr81NDcsOm6NAlR2XcxZwbLeZ+8CYG9iP118HsTqZuBQplD8r5217kGN
/ovb6SIMQd87ZBJDcoqDKKvBdccl3qSz2/XSTXKuUNRoTfwoJe57moMCHKWm
YsfD+WLrtGU6Mn2MSR7ajNnJj8TRs9D/aPLoucixTcjPddwFNW6mHQPE9/bn
TNm45TUcMjZ3a0rJz+9Vv9yKwq+ZGhd1WkBjk3+PHUgjOgKc6ky95c4ONTlD
CdMdBijAQYsVVwcm2I44W0JWV0Ai4aLd54tlaA961JUk6Ho5/G0KnKFub9Vf
kW92Wki9RaCIqzV5vkJ94CdSVB37G2ilVOPRAvmBR+gVEMzanvFHSeW23fUe
x8RdzYAMJTUarRLpG1E7qRfL/U/+Afxy/FIroMoYogUjG1iJf3113F5gdfiq
9zKV/OLxJthuSqoStxmUH0vk1//Ot83rQSh8u5RPofA6tbqOyu4flx7ni62W
JLRPkCvRoffPchMsJLp84vhTeG5wB3TNVXZLWIS8O5qC1WsyiwfTJ4BOdvqg
a5zzJdXQ2zMkINtS0hlnIaim9US3YeVKN2qgIrzWG4hEDgmD7lWAz5iWQVUd
JJ/c062138TAzJNkg3WdaN5UY5Z+MTgqjWHB0xcFdC5nCGZmvxJARHBJx8JW
jBchyoR3apjA6tT7RQ+eixtQdqTkHS4gbQ4CkY9YaS6zkXBwIBRQNfsIbP9W
346dqjdVcJgrpaD6Xe9MNX6a/VpOnJ7i8B3kJrwnUaI4vkN5hjF6qhLzndvi
8DMSgBb/9Yx8eMYDiMomFOD/UFZ+eDrL5UeNt8VwRgtjJibYxziNnTFzXt+G
YbkfLODJEfH1l+4gXe5hS8LWYorpwgPcFBcsDyimjiBT8qi5t5SwFca1mgD9
uGskdlut7t7+y1Woxr+UYY/3Ku1k6BjjGYx+NZssGUpKUOGL4IE75DGBQQIg
dFjvQ+sA3ksWPJOZD/z1elfIdFdLTV0EDNH/gfGw1FG+P+dPoP0Sx2PN54qm
PVKgJnrJ/Omdts6HFsjlo1qL1IbKKnz4neAqIVMofG3nL7dT50KDLqUPvBTm
Fx0+W4n/cZZ+WMj/ASwUhGhKDXG935WViYcBp3FNRCORCJz3zEBhEIfB9Znj
hM7mLSz7O2RwMZx8ZKjL+U6+ca+dTB5WjCi1l2b5ECKApyQc5NS6B7ybJu7/
+K/w3RhuZL/SBkqkYsjHiWVk0/4bipfloIbOiB8cEu/dUKGGOSxpWjtkXafK
A6zoBMI40bCHNx0wnf2pZZEE6c2v7LW57ztFYBsLTPpiqMwbCjZjVmkNf2R6
vupW8Ckctt8H+SXENgsGH9b3A8mEWbgy9vl6QUAn8OHklxsIrbPWfRggBw2x
7L52sq1gZMMwE2aO4CQyYFL924Yi1pKyeh3g6hOZtOenF0PwDM3RkUPX+E86
b51qrMMD3MOwdJ9TKhLHxMk0fhdQbCOndoDQW49T3LrBxht9SFqDltBOml1j
MkBK6XEvS8hGPpnoxYMRHlGCB5QQfA7TBiUoBEHmdEo+4WTkpD0UrSMbY9V+
C8oMPB7AeGikMPPm0AD3AySU0M/0olbD6YDOE3ghO5uOGpgr6WusZfNfvUht
BUi5hPAcTCBdV689v5GVJiMX6hzsAuU9dBsMKmVPEuqjeDJq9wrfWAzWQLuA
kOlVDzP8F8CpqpbdicxzYXyeqASU4XvyBVlASRD9hDtqZPSRj5RbDrzL4bx5
/lkIOGCFBetEZNTuJWQ34prZujsliKMVYB0dV8LHwiZq4/doWRLVsnU8RoY5
05kWZduBa4QBLcpnfw+xI8Gx/1S2l9V3iJcDifP7NeJPWyw2QjfeFXrF9wUs
f9upVAibUF3ac72SUGJc+BcocE2uw9kZ/EtVWwLuEId+MJI0BFQUykaMoSbs
9vBGjEwJvM2TkLvNxMcDoTlEzuDhlEfymPB+k3w3NpqtOp/9wmuyk8PBmZdj
l0OS8HU3a3Rav55mXqIO4RDdgwQBSaV1TSGswBMLI2C2jn2CvmoYHTm10MPs
uY2Q4OK6R9GxmTPtH5/BqObmtWUeitXXPqoABxuJdSlWm66xvLiIS0c+nqoF
PHdq/KXIEyPLpG84DrkPPePc02PlHfdKJCX9VlohuPw5cEyc/ehT1bXaAAjp
yx3v8fd8kiT+qzt1B9hbYb6+oMgGQV1qg+HNTjxCieRLDA9nR6oPmGNcADkw
KD9NLbxSYeAz62gKbi29NKP/dIrarfmIpzIyKKlLo0I9s+oCwJcvWU5E3mSI
n6VrgpIRznetXtvuneZ9BX4giMMRbrd39eEFJqcg4rUOlVv4UMV8Ac9CZ1/8
9uRoWicl3j6PkI3Fsjwx69EbrdKTq96Yp9BImtJ2PaXe5XJwfpSHF/c2sPjj
UYfpsFB9bunIKfRNMoTdSrdLWE/dn7ybSlvg2HMDlQ220G7HBr2AKZq93pBO
QKG2J+imT8ZLMTLjHhpNlnU1tz0SIv1ZO12IxlLsNaBAa+N3ahBKVN+NF+B2
UJfd/o5HAWa3VFmRkcsNbjutKkBXRZx3vHnI57rW4D0fIMJj+tQxTl6zysD7
L0xjhXIzzn2VBNTxoN1m/nYIEvGLoPG8Vclt4UMjnasXq2yoMS2MY7DsV4Tg
7CATcCXXnyv9uf+lG5HuWNfbtw8voEL2IFUVFUnpHPxb9VMqB7GPLwlQU4/t
N0KhhSX29feO6ZimPs4qDbkN+RUevwreySjtzxd4XpNRyAZSNo5C1p7dp5xM
oyZufiiCdIH6o+HOddAq4YBNBSfiK6wIyFxda/6s+40sxjw3jqNVUbsFJDD5
tJ75thPw8NAZglV5fCKNNrdDjA//A9PjqPjJv+iyNAnnxF+rkBHvNlLCzPyv
juH6a8ROXkpMxm85ML2Oy41Kd6Ekfdk/50sgLkYU+sfIJk+w9H1NABZpAtVR
X5r9Wo9l5AZtYO2kc55R8CbXmxd4X9fKPOFvBkj/xjw5Kv2E2HrS2TjQa1B/
GOBeSfEcmRUEpWlZ7Kd0EVxOK6qRp4n3Ob7dfR0abRZAptMQg+CwoCOICtO/
ykCny3r97qQwOLNwAbzSg7yS9mwSE+V3RdJ0+M78D1h3tnyNFisWuJ639Bqe
mbrzK59FcS3Gn5aszNXrGE7pTtJWnwawVbQqtvyED8UvaYgqpXVjr9ZoJ9rJ
3nCWkU3S4FIVjjmNSYDV0EUQXeeGKDz27Vh4Yz64KrsLnQR097aaiHEgMNcr
G7F27o96Otiw29QRD25hs4vFCx7hB/2MOLqNZgwRCdidxhzXL3+Fr3sCQT0D
K+YQWdCgEWmGDDxzzyrBwlr+S9nWLQcGlWVAI/yDRPR55anCMsCRaF1Aol1r
EJtB1N1fql/q1GPXP9fn/6WvG3cQb+kktSZ5Oce0dNLIfzzKLlPDmDfgrmEF
HZGJdOYxS86L6BHfDuyCrvr5brvZhkGnEIW6Oq/LkmTKTiY6F4qrkT/25Emd
jlGyPQIBRkTBe5z8qgLCgeEAH8VAeFGIgh6h70n8roaM+cSBBBJNslElwya4
WoccP3Cuw/TADA2erQEYtYT/phMx76Ydc3fWiX1WffjhYFlgH92pKZASNWYd
33fGJfF280a22nfDuqM+Dc13Nv2m4SVsuFlgpCNlVVDhrgg2L1XlEaiyTdm5
n5/94REf3zi/hvA55e/mVkiaiLvgHxHLBHLylqrgP5mqWCXiWA8MIUzeBhbL
NGkyMsGpraxOD0/NKUVK/3bQXimO7IXfoZ+c3KuMXuS0pnapWdwvd6tUccXk
XTjoFUTdg7vA6+H2QvLx5cEncQfcq52UPgfH9m8yt4o75hpgpZ0pz4wKuJFv
XQpKKgCv9sVNbnRjHpOZqTLsO3wAokpoBNswvzZjd9rAJ+VDOhV+D//6LSzC
M0bFSfmZFpTxKkexvvjqYY6LfRx+siQUEpwU/QEZ6xig5BXShbMy21PjLxdd
8IVltSyoESMgo9vHx2Y0quPSZOFx9NU0M5ZvAG0P/3xj0EzdXrBunI7uTWqI
HNn+2cfAd2k6K7R+G4C8AQ4n9tcAkUs+ikViHpMu9BeQhAU4K0SNEUC3G9oi
TFwt+ntuvJ16xbYIepmN7guNg4kWQIJ2VfoK44l0ZZy112SGgYRGHE/eu1Mr
OVAfmI3CThaXXUrNIaz1zGPjNw8uDQgvBjhuQJmbokK8sd8M7zcPP8AAnVl7
5KytCWXMSeMB8QqrGdtM5YLMY3eBi8Un1DskF39k+SFeOmOZByArKm3NBN/c
dF/CZe1MUZiw8CBo8RN1MA/8i+jx1LxXcP2GtJRWZ2aLi2VLJdmw2RuFqvBq
bNKFedt1iRzoi9nWOE8CAu6YnVva9icUe657qHnBZ3iqKdRnKXWO44X/Mshe
7/dTut6uXm0KswRkw5HjrbCcm0P1wHK077SbA2DpdEVUzN75yJBmlh4biVdN
tkOxhE8Pqy7qT85zaJ/LWMCNRXquCVUm57nqYJFKEdldhIER9rkVJBRWxCAT
X/b6qDOxJHsvC0QHTKqke4qtidyXDwzjqVn4q3iZovjzyaIrXTY/SiKhs04e
9LoAZIUidZpsEbgmfvxzX/PhHtp2u6eT/m9GxamvFSps/DrbbAEniK7kZI5P
x7mr0tEYfxi7WsXNGjGwjWbH5wDt0LzkMgBDcGOlWIH1A6br5/NCFI7R+3EH
oY+Hos+uMV4gywk/sloYE8OSuTwS3LlauAGSOhVxQ8lcKqc37o9B23OGLloo
I/EZx7E3X378zS1Gd9qpv5V28J8B/SA1tERqc7QaqCamzYaBqL5LoOgNCEee
3+CXkRgqIJc8I81ycwQUYJJg8ZUcb6gj7DaPPS3ckTac66EBLHOBBkXGmXn5
KnT9oZbd1o87DjCS/AAQt3klFn3cWjlHbDJogcqgIBF8VKQIPuiw8kObmcGC
n7RnBJNncKlbM1ZGYbH3ES9xFKt+YqoN9IEVBnXATVWnW6+yqb0HDvjVc8N+
nx8phycrl6BvSKKwhhKUatKjqUxjtdgPOY3B6wKN8PsJhVmC2yQD7Al/4eiI
Wh5+P+L6top4Y+Zp0WhrroDYU04x4nRZ+u6mVfavM9fZuKOPKdQKWylKG+Vx
Yu3Sla99fJ4SaNuRNOhSJUtZPvZe5n367rOVkZKAEFK34QeNtxkUrdWP14NR
AzNMQi5xQF3OCFS5mMtU88qaBzxlb6Zr64zC7L9DKps3OlJSPJpeUZ7sXuMa
qKeiJ6mBg0bfqyLNSFsliB/hPHjIO8zPmcX9hsiy9Vu6DkCfZ0vqJgCS5UNb
3Gnx61xkbJyoMFwBnMNe2pcfdly8V7QhJpYjqMvEmKgi2aemSkQwcliznXnw
jUAJ3t44IPl/Ctboy3bPeugdvYbYvgVacvI7NLSo8aP7FXtxyglqVdOu/7/s
BTiwQprtECTItWHPXzDziEMWDSRDxC6OY+JciefEzWuq+vsuVj0uGQKh6riD
MUXiqiC5EoOrCzs/t2X90sPIBAFBqWJ2U3hTzKj+q0AEP8oOH6QWsjOeYHOU
w18PZme/qNrgY94mL9PaHiXNYIoT3Lw/l+9eOQGubeRsyznK4t1De1oVNcWH
N4LteB1ZFvUe1Fr1Rk9lnQJuADzIhl0akqaww3zl/Jl6N/yHlb6n8y+JSanG
1HSyNfXNUq8RXxl3qzMNMwMxkTRskADg24abxfnb8mBxhblbvkqEPkRlxZmt
k7BtcD0DMUkgIN5vWfDBYt67lcuL3E/jRNDyLwcxOuVR3KEkx2XU8MGKluvc
l6tsnQN9ScliKLiVtA+T5l3C0NW+AqcwxT+sP0ewuGUulOMk8OQyqU9A8/uz
LCVj15KGZHkx4w6eQk6e1od7LfgbYqDdRcdFsCIXcxt2pFN2G+T0rFsMbLcw
K6Huqt9BCCtAkLHuj53SRHvzFU9FVc7GPbgznLLMqSf74AM01DFWjuP80x8/
wOhs1/jJwMzfizdhtpEOYBCO++9umVifq4HdjIsMrBMuKTN6dfWBGTt4zOKu
Sg+I/5+84f6Ei/9UfOKFa/3zSnWuV7yoCVLPYDfG7JKiBsOn3HIDmW8OKH6A
+hwr81tGccV8Ywqojlbj34A0D7eR8cVwuIbF+5kWubk611SmCOVwH7lKtf2v
1nk2TBwd23rUBpPW/BvCi8X6wnPCo17vugLzz59wxuJHx29TP4rox394hZDX
ygI4jEW/vVGySwkuwBRgWz16V7QSpBDsH+f/E3AvLJhNCM3AlXbc0HLN3Jdh
5lZ+7ULLLG4Uc9HyTFmcKPampEi/pbEMJK0QQSEJkXirbYtMAwgPkmAIsF+L
dS4/TJNcMgDyR+ndUUVIwGLZoT7aLfW9rWfGdqIggEHPz0GxVOGJ2TAds/mz
C0Pwpt3kZnQer/bbIjCVY1Ybw8YjQeCK+q9ILPoQGjRWu6HVN1q6NcvdF5y/
fPwawBs6gIEx90RDRx7Wc18phDNp9fD6E4QdmUG/qBq9VKFAPC7KB1oICGDw
J+6vhLWV2U3LFierQi5MPgMerp0NC0pTyYYKMc4cSOC0L+KlH6zxd19Jjtb6
+ove6ov2UNBXPhy02zvgpoUTZW/FGEZ7XRdvgF9NagZMcktp0caEeFrJtdu7
hEdeVDn7vpjj636xteck4lZobrsiD+bCSo4gTdrLjlAXJ7cMIpzbRnPhq8Lm
vYOKb5gIEbfZPys+srIkguysvMJ7T84l39Grevfj3YdSOTAAw1PFi+itkXoX
9DtNCFBt4hAsMvMBvq7UM0XxOelqHgH4LkbKO402CK8/gnF12ZnCJxo+5tog
h8BLNuxgZlhYJFqMWCzKaCBs25gEZsraBhz0J0NUWf2ezpsvhXrLx1k9qr3o
ve2GiQ5S+jJ3Mq0VgUbFPJaxik5EZQqDPESyTQdcM7hmbS/JNiQdMpEKq1Lv
8Jcmi4+htmqdmEhA1/U5iRsFN+CwcbBSljwi5fCXYzocHZ+X9PYWfUKvSBJu
r5aLFpqI8bcQXxrUeFMDNohHyweh7ljxMb39bPxFqQVzlsotcK/VjGrVnsaP
0e74c1D+bqsAqqJMfIWtxZjyo3xrnw9m+/Iwznd4LjnRjp1b25sW723ct19T
19wfEdSKeQp7UYF0+g0vGv/1U2GilGO3Haw92zvr4RT7LiKuoLIkFJPZojRW
rQO6dFIiC/VskGihD8Gkr85LROP/DUO8YHLsEv3UCAO/7Y3LJVB3V1c7pQOc
6Qr/jE9WDwtcoKdqL5meQI6ZYDfXRWuGe3qPkp3DADYEk3tt7GcFym6ofybo
n/Hhw5F1L2xq4qDRndAPGHOT1KeUbjIuQCOcsUJMxfm/1UalTxmAmuVZlO3x
eBUyTriD+NZKY/eX/KqtlooN91ezavhEqAmoLoBjHGdoxSHwjK/f32c360Px
njoHhA7gzwmnWUqphsfnADZ1BbsBkrkO88tFRI1R4TZZWg0M7vsFrrUuIsn8
CAFeaYxCAguQ9pAX5+SWRIlBxY7+SXxj0p0IOGkeQ5N/fTLX80eXam2KRCGV
gkmeyPm2TjPJh8Ta/A3bdNoefuSrGsd5JTD6n9FyAo9VDyq/+EQJgIyTy3vw
NQ51B1VADxKVmSYjIxXz5My6PpccctMeLwZQFjJsUzwjWBkZRAPpXibq47z8
uKygtrttPusjkBiW1jZ6tdDs0LWMYEcnHT27G0FCgywixcNgOuPmIopWTE5V
miGcXaaA8f4IQWAUh/k8WpCfoGbQxdMDG6rmg3exUYx2UuJG6Q7jCh7V8YCH
aq3GoIB/Lci4uswcJcLuLV9MX4o6WcPnBS32jYLi8kHJsa8SXxeEg24y5OI5
kp6R0KgeqYfnUTB0/mWYrixyIIU6/YcGHcOvZbX/a3e4sfX/xo5bL4nxOw1o
QY1+00qscIXzJPE0sCWKkdGKkjb63Jpovj2lGFXNeGnPWMLwanHS+q0sM3Tt
YUr7WqgAp04C7Rcowve57EHNRdmKQE1J//1WzBr5CV3euVkhDMMhzHYkzpc3
Nk5zO+jPYQRYOQB2pXqCFW2jZssI+0U/3kOh6XLSB4qsGY5KeMqbV9xTFBH1
AmrH9Wsp+2Gb7qNBR0NgCABLrJtGKBj6wXsUDojtNl4dLNymgxHGNzgzON5R
CT38ap2aBqsZjlm9dW31PtSDavK4Fh/aPNmmLWcL16qslaWsE8sPCzDbgdze
+rZuZm3X+3dUCBS49GNZXTmol23Bv1hFdndkavWIN5GUuwWAUZfDnueQeEYg
GkDMXVffEgykw2aQhPsfIv/dvOH831+JqQM7Dfv/YxOYLJZWe15ssu0GxwDH
/pIcaMBzdmQ4VMKuZiW5dufAhFCkfpFIgm1679HOwxKdT6x1+aU6CTlzLd5S
uhbklr4n+j0Cn4PrbxMeIih6B4ED0e0Ufo5Dz9L5DMJCvT5Junz+32RStzs5
Sbt0Omo2f4f8N73jhU5G5HPR2LoAD1RHTGe+SrLP9GEn4dQfGVIDKW8FEKfF
Ti+sdRABWxoVdqrMs2bKIjT0kV8uElVXFrrhXbeE1zfWEFVzU30sbXENuw5D
Ti9dzzUZS/DnwHHwANaghISbqCQs7bNGHpa11sryU0hOAsga371vOWS11bms
wZTA1bjZOInBKSH7yLdXIaMv3y2GUEUtx9LMfV3q3x21Vn7lEPtJcZPLzbi7
XdpZfnTD8O/2UBBkK2OW3ROE7YQOVCLA3XxFjtjm8PgJgyemkoev/LTbY1Ku
c1HmoWQKkUZr1FIxJ7H80Au9C79CndRCk2cMoPF9Maxe3x2I5AsnqC9HEp0e
XYL+PTWRlw5VPD2FFpoBXW3F0H+HNXLP22VR5JaJfekHUvxtNihPRYuAjDAL
+c5hGkb2VaFMyUpyXD6CiOYdYmND3i5w52TaBBknkKW5YI78eShVuLnK/Pfb
wzczJ2Ax9isLNGfYEWSJB3Lb/km2tkEYTi+05FL5+4q0UzGWgJRwLB4gMpDP
VBOQjUywCgAjqHBu1sNSy4W3NdRqECdtJnWnO78YDCCFjWuWIBQEMLEtDxAp
T3mj7usiDMFLe5CYb1NCOOUrGHTuvYJpmqjq9K9mteMvfy00cNIo2NM1nh4i
XUNOLKUQf6fuQt7t4cPN0KqcdjvA1kNECIvn7RysqffEXQs8Tr6hRYIIJXD+
EnJPt2VeLqbkdoWWq7MVrLBQlVhIQzglHoc7JYWBtazb46NEmM8m3yW4UzOR
3x4ArL+RCm9mGTah1K2Q1jWRxXEwRq6qHw42Tz3bwmuI+iLJHvi9DKN+7oVV
vVB6Z6a6fWCTJVgaKspzxTHAEE8SJ7MO/Sei1JdIcCfjGIqfl7ztl7X0QnLj
9YqebPTX5J5QgYS7Q0nJhipTU9uUHbLE/zm1SEbxDDKHOljfWGg8J4hlHZr+
7b9IxkN+O4bdSJhWQuVVxPU+R53dgOZAHxGihJLtU5FONHT6fux6SxyXD7VP
BhOumXFr3AfvOGize2eMFRLGQIaS5ceieuXsQmIfZDtJ4Mio8jg1PseLdbWr
3h6iCe38eWiTZh5lpQhDZBPa3sbULLobaA8+YHv2wZu3vIn6E5jT/RSQMlbr
IdcmAraBxUXbStwSLkh7y8Pu7IvDi1LlhiQGS72F98Secy1FCeZCv1zG7F3L
5dK60GNZzDm4W28hdcf2QcZstls77jMl4HS1giUZF+BbXlY3xLA+B58Af7Uo
OMkSN9HkRFYiRYUO3V7Zbcmk1qqj8GYWtSer1mbN/Bj3stb0gV2mAX3ecgD8
lR/fZAt9uMS9rQMQ1lG0cremcGHzIYx4B9rnwz0TAGHclO2EDsTbccXIV2F6
wjyQ0N54/gpFYZMFVQ20h4v2nhN6mWqMMnkdirKIxAmAbnK2BMlza5orvxhz
QTCEz/0nheKqxFPotQwtcDjRd3oPlB+HqmpFsWL9OTMxqIaX2KcMxPA2HDCN
kFkYOewujEvTAq7RnH8b0aYiI9/DIaUCdaotmGB9mwe5fubJoQnmvybXyu/Y
YI0cAf8FJCrGutNsZBLFoQB4wGHM5n67/3cM12Rbjz0/yumayLcIFgU64NO7
pL/ZA4EF7VSCi2dq+XTwceVQ0NHzUSNZVA/5pF3rZ2pwEBTJjTFF3v+oC5c5
1Nr74qlRTqTYGSKqginuKQd/uBj1PxhkRBJWrpV/6zDur2r+IoVQqDDwnz3T
ymy2nCKYZB/Nbc/qWS84tk9oWq3BOuQgIJg6JsikFo5IKCateMnfSNJs0yST
98Egm4nRImrAdyVI7eW1lgEb51PVg9xjrWbTboY6+RXSnf3jC9pA+nOxEiSP
emm2aA+ThnCnh/eI4aobu88n75/k+TXNgslwkdlRX7hdL6Ekg8u++ek+mfp7
jCtrNv4XnqqISUEn1MWGjjdBPAusziG1L12Rcn5TTc41/HJ6n+z6U4tPaEtD
ubEOlAx25UcNMGC1VUBIu9w3Kd9sAYaTR6EOvfRVnZ3T3nBlIIPkhwc3Yqrn
y5hJPKxA69k67mMZ0Hk/Q85a+YAxar/SdAmxqeCoNADMWzZLorXCdTJBt1AD
fPphN4J9yxKVTmyZRwrzNrlClIhLkKJagFeYkqs8Dc9LQ+w4DtsMYOZRHzo6
17b6z7GRUtKksGvgKb3Z9l1X9x6Q/n45toWLjs8MLyInBTz331faP/f/2SGO
KX4e7URHHUyEG905Fl5xmgAj9cPfMIY+N8WV6el2Dw1R63JQ5nHNbz6ST/MP
5T+fXAsEWuDrlUMb6hoolayfvLDWBaW09aOovT2uGHt7M28HbpgSaVyKZP0a
47AbXTOBwwUo7O25PwGyGl1Ml9498jiNZs5s5wgQJYgYzZT3yciu0nXaQ25W
dfRu5LXUTyDnJnkydI8TKeghylDKsROekenyEcboTaheTgBGVKBz+mLFiOJr
AU2Ol3HnqRfD4ymDM1P+PTRb/+74IFzkN8f/nM/830AfCOsxHmcTn8g+sh1M
ItbyDpOCAFLPKQ5Szge4n3D0ogKWTZAVVXRRzqW/Pxpqziv3ofVqemG9JP/m
Q3N6N5/5VhNYQ92sTGduBimpxfMiz+sfxP3hjpn+OdnsAZmrNgr5tEGgbnfQ
ahMuYGuVWtavPiYwZuJZCimpVoPZY5G/cZsGIJPKsNtFCSFyiU9gtesxP5wQ
psafmHp+/g8KQKmXJpl0cUsbmNJOwwQgSSti5upnxTW/Mo48U/6jDG90ugZL
a029eH3xwDLzitNg5Jzg5ETZORWQ7DK8bQobMJ3YvA332x9oBqdW3AFbTYNe
GtTOljfVNNmW5ysjFlxKwNzLCtA3AJJFezG+59+fddAToTaqXQnCcthS3tNw
FsWBVu8htFIzs0VjUVHNjGJTzYXjLTLHtnuuOUU1NXOd4Bi0M3nufGjFlam0
Mibpep/g0707dFvjrqR2u9jpjCZtw2leHkEOHxhona8c63FehfzEt4O7Mv0x
EDRditCAlI+51KxwvHbViaq0+vny0Gc7P77t6Ha4wLwE61hKr+xDEnSyJtCG
tWgMzM/TLHKlFpRujqS+AdRWlLL2/R+BwFMjHRDZtFaVFBWN6bWReAEyGP4A
eJOglh0XXRjTwnWojVCeznEw0uI4rsVOOFM6lScZM3Lamxh2gLwygnlacGqO
I6Txuwa4Q/E8HpU9EUWaK8TpLXTZYrU9jIVd9qqOYGMQonzV5rDwcka2HJEC
BUIjR4RphklPzNW9Tge6Fu81QMNTvj7bCjUH8r1iWrpeAL7fReFPOo2pTUGd
9d4XqPflkMFHw86m66us+2FAL9WDhGRRv106wGh/4w7wP7rpm0gydo/GO/ny
f4KCjdA1zLGarnZp7DWGs8fMkwbAjHUQqi3J/HS8ozCrfPnpJnnePHOYFvUV
sgSub1IfxXqE7g7KFWoPzEN7/hbsdFniy54siw/LQqbhpnjd67IJDkx9Yjym
mH0cKYIQlw3j2XGU8phgcEwThtXyAhFlAD2+rV7gWPafRmoBkW2g222LJNHu
CQC1qSZMODSkN0V0Kz306iDrxyT0rw/B83N5HBvUCaDbOsCUVefZAWdCu0mv
iT9JqHM9/hdp+zR6Zzf+cH7s3h7HTM/7FvADyCB6hAMzuCOIYunp/ZXJHqCJ
p8ep8E5rlWA2AkxI+7yd1wpoSjopJ6RM/UHB0E94Ze3gPevowIbaTZ/Srcvn
rrV7GExTjGB4c5aR2Q4t5g7SCs6ISIrMhjLrd29IP9tItIuZTFLtqNAgkGl3
OUI/AOsSSwFpyQfET36YSHl01G3stjXXZBygYQktJFdToHRrN+OjDf3Io0GW
BMMP5YPQNorpnuoH4kmP9C2Cz3f+7tCSg4ESRJezUUFwa/XY/vVYokxCNp1D
Sl6dBzCy1RQL2FNNnTMR4cghFnrpH2/rvkaU3JL06NhPru7Juw0ZO5N3D43e
V6YR0HEUDb63dqzBcyTVVkZKccDvwBOcRDOmSKgNcqSFVx8C0O9rl/PcHlsk
evlhc99HHf+AmJ3jykVIIEKztGZvoPI65z5em2IDt5xLEk8up+YmSLD261sM
+T9HTB9lggHLmel3I7zI99q+g9RodCspxCPKvbU3ijq65PvXU6q6sXEV2cGA
wn0Ckiu2VJotBxTqiTnt47ITQKPYu+8P7CGE94T90B1oftyD5uLuCxP12EAA
UtVlPa5Yjf7t0LYmvxhX7VaVqA764WfCAKJRIjmUsI1BNRuZLuG9DZ1YRoje
IWySkP4H6BZvP7FoMiBGM97+XXlYUkvVXXW7Dj+pDq9vIwGHGy69aOjBGNys
rOh84M/GS0g5a9/T/doXnhEBWwutdjzWY4K+al6c4enVcb2I3J4UrBRm12XA
kvdO7AI/VMnljfFEdYRmyzbv+oyyde0o+o3FuIwhZB0cn5ouC0MIGgal7VGZ
gys89YQ1xQtZwHQw2N6PQJDxmlJ1sX3uioYcUcOXfwMMh5KC6VQU+q4U9evV
jmxoofFGvw4g68kozpGo+o9TAC8KgfAwqhtt69o1mrG+OR2B7qlibnGbfX55
LRSeYWdCeH2Z/QLykPRKRwP6PXGOiPO25pLAV/cliVPaeLVdFF4pvHaroOX5
iR1jyZqKrKDfR77ZRVOuQi6XLkW3eN1aG6cXviOWDjCRdLFHFKQ2WU6wL/YF
ZvIbSBJXzxnQdEzG/qkM8buipkXYfRvYQvFLXnwCx0J4tFuapnkeUT31V0CJ
sbcUtJ8VrV98YxesY+kori1iOMmiDU6Squ3fVlvQdWDV0YKB68tqYjCQ0p4Y
Xp1uFjXk5olAR88b8AUnYpGC3DJ7Ab6+5xIOASLOmI62i4HLM9+nW8MoS84R
2jUqPiJI1rasFHPYYppfJ6LHhpTNuZSaLlv4nAL1JpMSEFtPFkH7GCJwLSHa
tkERqiyZZrncv6BBnDvrS0JDpZFWJT3VQjpTOhctnG7jJPh2Y3mz/zxBOdgV
tzhpj/+OlTovhnTFMAYw4Z7IBxUuz8L2M9rcbsKtLgXtAjwbbOomQnwWyHep
GnBenlV9I4Rnez2YcSIUqOQBQr7cIJMa+e5hORs4E7BT3SucUc8hUc+KlWHY
aokl9vYafBKkyXidT79VIQT3ESPavKWzDdhNLevjh/X0ng+KoSLWM+o4I05e
Ak0llXPUZ++7TusaLRFAVduX0XN2WaXzsst/vjkswUmbuqTkbADXvtXKub+1
uxt+Gkke8Bvuhz2bm6jjM6BIMAHlSt/2NGSsRgFJW6NmqQbqdyo/pidtiSCb
NI0eQj8vHDmWKdMiUYAnEMNDuVmVK6JDNiKShJel4R0pcOWLDSPYpWS1aEo/
c1defgyUsiRCSTyoc7ARYCqXuREfSIZEWFRWCoTsh5XthFWwsdZ1rVc2XWJh
gXCSPTw6e30THCrd2r+UxbwlTPS5OP51XSrftpKp0x7o/MLlRJ780YbTkNiV
K4SGpulv+SSHvuqrYX5svx9fzTTvTSdPgcZF5mKcAztWocnkQ18iE7WmPL2j
Rj694jBzwzRp1S+zM5KRdFW5DMJZnerv5IMaZrKeolkU8dfIqvwnGKUgoEBr
P5PoxfzS83BQBWpVU4dCYuizJz38se7hog8BcnY/O1Rroi+QCmcx6yP0n3Qs
DnqilgeYRB45PDH7aO+b+NjIkYmNaDQjmOvAuCQ9erMe4+hpGXiJI/WKd06S
GXMjEK6NwDOafYWphtl/7xp+pXySuIemqzbBZ5gS22lMrg4//VLPfAOMUmZb
Q5TMMv6ipCTmByTWpl3jtE025lrYIAR1zLZKoUGRyNf1Ft15KEBcYxqQ6dXX
SbNDjggvpPcepczjbGp7TIvNufyyOpnYdIXTeju7RAPicyzkqYnj6yNu2EId
20l730LyKSJfDVB4BahS2OuxoA8kZxcHAJQ4FLvUQ5nc0I4PUK0kunoP6zNo
bS+jomtf+0rbUDqWvgnT+kBY7cPK2JrK+4HxogvS30eTEgAPkjwxRP4Ihz5/
t1tYsPsyZynsWaI9kZcZGhJfra0bV2zvURzCGktlJWxO7/qFrr24iLzNkh1O
Gaez3/48rGlwaG+bLF5rTG/IDKJmfcVPHZLoAKQhk1hWqkwfU9WsI5Pf1/lA
/Oz9D5x8ntob9wUXouvayYHy2s2AD9YapiZkddBqePK+Ojhr09P5nS6hloOh
t8YAsWAK3RhaOx6uzzNGoMlXikqp4D2m0B7NXrEZzdl9GRP2FKKQoUboYaFx
FhwOTmeJdNwP5Cds1sFsa+ktNmEppJ3jV6JCyCZNMscHTOsSjbmP/yzEiay9
dOnW5ZqpUwgMvIdacjDXtSSVYRdiDVLz6LBhYS8XEI7deAGepVx1iOTlmoEy
jVo84JijDjeT4g/QxBnmiwISqtRoqHHDbnPwETgJ49eW00kWrTMUn5oKEON0
n2VNZaj8wbMjgAbddNU1j3r3Ha8f45+yJhnYN60z1Qav8f9684DhKGiBnWpk
eXNafRo28/wtmX5/CB3MvcYPvIxgn3A+jSvTX46eTyH+BYgJShaUX29BwAU6
ncDgKzz51vD1+9usAgVeAhENuFcp6dauUFuio9FxRaGHre64gqpKyXAJ1x9j
cEbdS2YHZXRP4iiRRSns6bNj+Wcd6L6NPXDdxCrCHp4WaCYTykimZfxu3Ovc
o5cF7CoyanXS6Lgu5LMGigBdhHHZ2H1ud1qgrWd+VW1b3B6F6/jgXSDwzSwl
YrGhVhORb0ExtFF0dlHt1OGqgdZMMsgR/od+TfO4hRnXSZOXd6Vb28K2WizZ
cgaGH2hwoLuYO8FXwOX2n37wC1JUGuQTcyaxBW0IAHQ0dc7YCWjUM3MoX3Ku
1Ji2y3HG0yFyEJO3cI3pCCAaL2gPRcaQ2aLcydIt/vPhDt9ddxpPQurMtOuk
FMZVnvZrvNIw0vFHbz0FyRVfOlo2bZ4PrM8p+fucR1YTeZQ0iIduJAfIssCE
2z9VgY4JhGkFsEw/2hEybqqByfSeMUSo/xV3PtdS4V3H59hCj44t1FNXNq4E
BL7LZhSmAC2dSq6wKQ6l/t2cxOADHQrOuJMcFxtPok4aqdOeXLg5hLpA32J5
BiQKGZwatb05mducDUnPAPrtyh9yzSxCoutBZv9CmS9L35oiLn3OTpWqyp06
CdZ2FuhEh0Y9RV0TS8X3T7G8pvUEcQBbr7ShYR1tmN8t6FOQM4A4jcQg1bta
aFJuai/cNhQx6lftZexWy3IaDVKW7frvHZvM9peSguHtlKa6vAVA/uPtvoeM
eQjWrfwDMPn4mgAn+HFqlJC/eW4cBQJdfljGvsnfjRIgYtuHt5dsLLTO1XQW
BQgKP+sygqCvLpIdyHby6sksI9JMF+LpELYn0OerncMYBVJcf83fky2hiLqz
dU+h1Mc3xl47tvTuZhj158ekzeHxzHmzHaLMcyPNR5kFQU0NNSVAYGqqUAmu
EH9R8YxQPI4K4/5oyXBmx516PnwPyIBW/7p360nssmgb5mT6YQ1wTmko2Unl
VsjigJMX1kMlz53u25Zss8wtn+YVFT/mnytlZ9vbqBQhf8+Sx1jQf/tkMYam
Cmn6EfSGIRtnQ1sVC6yAb+MIw6TPQN07y3KXuK467lmi/Kwk8/+bFIbKPDKS
xzoubcm4Uag5mTuU6smbfjS2Sd1OAEs7WJ8UvCdMxuRPlX744j5C21yZy6SO
AV02DC4QmAyhBKGdduw0QodwmdLnJvMzvrMpDzTWIRceETxtBf6Bnav9FhJY
LpDtFA90fqzljpDZvLOLaGnlH9r5PBk3TBDU3+i6Obq8iuB0XVlplizwG+ye
TB7u2TXC1TYbr7CvOztAypKCbdM1M38aeDFBQlG8QnKQ1LLWSIcnTcPO/7b+
6mlDOOMcUwHBlwlY6w2JLairxJNzDTMgK9+GmrFxABxKNItSvKZXFlTFHtoU
9FEPUO3UaoSpZAXHcClbIhfNkL7geJNzFLSd+t2pwHWQqdYfW45drRDurXeq
NMGRPfSfzXypZMkBIUoXOjr3bLr3fcUJXTR7/hgMbusbGzvGyaqv3cIhftiw
xXlxfke/J1q/BeYluB00iOCIY94rwO3aNU7OdgTaFD0z94B+So+49D8D/hRu
6ybWUcoMiLD33TcvTmM1OEr2SVA/XI9rzrIyGCxFKGUaWkjiwkFZ/ZP8Wdha
G+HoPMZhb2LLehTYDT44hIdnSskz0HbY/2DDEzemV3AP/N/LzuTOY84sXPao
kGvohWXboIhYSFpdQu/zwxeSsNB2iMSLqxPjzljauRLyBAS9wvtCV74eEmO4
RfNYYCsmTH/E8bDSVXWzEZ8XaL3gazm/ywdR7xgsdpCEmaGnwReAIgGyCc2U
pwdvv7HfXV7s4ezc57z8Cxqlaop1PkAYORsTCgm9ZuPYxyMMTubzx+zxXf0b
pMnb62tcfGvLlPHvfwyjUxlw95oxJcdLXraGeuR7OQUdkko50ikToaIlVIh/
aEeSD/9QWQuky39Zt3Uvwa/q4V0d6PVZBkNbQyvpGZEF3HcqOnO41ihWJ+19
PLWiKwJAcch1Xs3ZkkYNr/Cp2tsJN+SveK2KPLKeGJBr63eQd/LqMYndGsTs
nFtr+EIbtztJOG8ue+Rg4Z0K1UPrKgoZSPYxsULlxmlyMsjkKacffP4fELJz
sdKaKRoUq6SYMpvrXIrd2CFM+32c/VZgiAfng9SnFV9uwdxfePivVJLyuaX8
sUaRyXGdu/ZEd+9yWkB2PKfWNFwzrEYMf5zYlw/M1gnYWIuHaHFFB5+QbW+d
R67U5Je8V734pVv8TJx4ILyRcnutks6CjpFMqlC/59IMV4Btg/CMZAfm3nsk
uDv1HP0day39uBkCfkE3oq/LV0nTYhHKNfIY23wzwdEyhFM8OSclX+5HPvNN
iFhsEHai+G3tREZTPMda4F/L+f7a1Z3BdCdpT9Tpfyng2ZxeRINGGcCDOh/5
yCecsK+6WWW9UNDvwe+esLZdCw9d2LbXFHh3FD0+fsTIF5owK9cXrzKXTfUG
+iohjA+velq81PP0Zv1VmHoiOCPELNcKdbXgRkxAaxNiG0EkGynr45wxItml
8Q9RJ4YlW1mtvq6sI/kIro0IKNT6OhdlgVmvMGsOEm/cYHtOhBpYJFg8hn06
5V/+OxnhneR16Xvwgo1UN4PPG5wsXWF9cDkhvnvo4HpFw95ogZEod57UsfeT
g3bNkQ7jJ4vToai+h8cG2jTj5+tiQEdWiW160+mwpOE02fwJxyPkDOhtNXRZ
yz3nv60BB7R3JZ1/LQQI9t8g9jbsjNHN9MlSlfxvEpjYb9a+mon954Nwn1mo
QlF8FpQVLcjxULeVtz6vi6xNCEmLXrxSvMfrpv/wbXCuXVY5dZF05RlcqxLa
jI7l52RgcckNA8oPVdh4LwASCKV0XEkR/1ElwV8dzCW2nmdjgvZrcIJkTbEO
5EtKqZ+BsXBVCbF8aC1CvU3UQVkDd9rS3fM8JR39gN4+xTd1ZlLFKsEVs7uZ
78I/u6eNfe8sayLlkO3CejQJlZ6L8Ekajc7QFnaBW/xhiGCIlWDKFDMnGw93
7J8Dci5CYVYhvI76qt8AS+6kynmKoF9mtNqGf6Joe7PL3anKQ5vOMhoTTFf3
xbYchVf2VVFg4qOylaKPb7WHUVg2/rmxANbhbwPoKZZtRGN+ae3E/OB1f+Rj
q7Wj99pJmRUnj1x7A77BmSI6yQGxp5UeIF6jtUkHA96MW2bnrPuJ2fl1zNr5
OAeHLmeAr36Yf7RbdfN5mjngfJ2/aUVEV/jDqq2dm6O7lliImojhnEK98a3B
9N+zZPnrvUgmZY6GUUjMR0HjFgIqXLThQAB8dZPxN3sK2fsvicjS3pF1l0Ek
8O9Y8tHp4oEklVmsheII7P1BY9mMcUWMSOOSAJof39q2SgCgcWwKv5O51hD+
JOgQpO3+9NBgAwK61rzT3G5D9DtHZ+7YEZfo/VyDTyI4X3EmUuN8pRoQKILg
aawbOIQfPIIm1CafiA6H17YOvdpcUC7lxkf6m5DYOJlbjT1y+7Ig/W14tw9x
S+loqWi3n6qLwSOrRq8PwuBzgtGuwIXuierxgf4UEXRedAy75qrPivdycF5A
O+GfAwZ6NDyMPST8HMvL8N1T3YfyMX2oevRL7bN39qMhSeuAaNm3QG0g7lut
qGSc9Ez4PYqpqGD9563Dmlxkshop8ciiDElzJW/GVazIQ7gWifk3o7qnb/bS
ASqwnuYRTy5kJnbFQe5bIj2b6rWQZBwxUucSCcHl8qlIuQm9J4zDma9CvxJC
jMfroqP181otizinX/zHbHc6v9n/dhHsuPef45ubrC4apRT+kxZ6G09NTFve
g/UW6h5LwwyiXz5ZLnt5DPZV5oV2bpK0r8/z0cW23FBrtMQnO1oWSdUHAVpU
Efs133EU17q1vwsTrJQaZ32sjn8juQJH9hhQ2Ff3X/Br47fPk2RgmIqu9oBr
fZHEEy/a9O+qGlKQssBAuuh4AJYyIAMbNZyL1abZpABRXr7OKaZIz8fVxoXz
5dJwE4IrEoOZfiZ4PAglSryxbvU9JLKgSHcR8Lamf9Z+iWgV93EqlGsuRIwF
MOuHrzWQaNTYIDasukOUw6bYOxySZv4WGhI4qFsmhFpiTG5lzSspSOFdTLNs
d3WGgdRbkDG8LCdRyS5Mlfrd78NLHtG4Q2DtMGLVe6RGzyfY6zhm0P+MCSGu
JR8rdR71Beam3CHt9Nxm+n8i31rgNglJf7BFCmQpaomLFQshI+5bukrZQZFg
sn6cgKWn57NFLmzdrjnFtMn/fqx9nHCA1m4EmYCGmNyniSQJppMjgifgJSo0
/PS+UZdhE46IU+Y37fMUx98/MTtOrx3C4wJqJrqdYeOmNSnjeQ+Em/sPHCw5
Rf3hbNJ9bfL4j53z0cNLqxrrznISr4UyrHGb3LCJPt8Hcn6EThjcuAmlo3oM
upwkqTrX2FGiNGnyXxiYIG53UF/UxJhq/0uXV9xp6dLzyxM/eOQ3Kl5YuBuF
Pkq3rGeu1mrYtyKC4IAVnJgwbpUL6Ep1sNBM5ig8LM95QkJEblSmYgt2FvC7
Fxe+pqt3em3t3bBgNyU4SvxU3tqa6JUQRNUWG58QB+jYGHfcJ2RiFTZ8lKsj
yPBCGlQgyUus2E4EdkQetA/7u4tyFsNnptvyJ7f00AvUmM3t5YOcs4giCZgQ
LuxYfcc5ObhBGc1CMofYINn8Hx+o+CWPc1Zd7PR1vasiOdB7WM5IozujX87h
CNH3VpqTqUX7ygh1uiu8az4Ob15pu7zBeYSh9u1XDwnG+BbuRJ55EkFUaDIF
Nq7zNUCYEwmhaX4BOquTC+xdt47VxjBdR0QuBibERYxtuHsUAdetsUbxOnNi
iLFoWIofRhP/sTh1yvejVBJcdVt/ddRhGmoQl+JcJGxGWyDUhXROwaS6dMDI
emDlGH+EqBX/2GWMw5v68Dt5Clumkz6A+gyFwO2YzsrdgjO2URK+lc7B/7Yc
sgK3fTVmeT/xW6tmDh823Kaf3q1u2aHG+cwBr6tdJgfsCjHQnIUeAMpibZg2
hzTkKvBNi4qVc1dKvFtawaoFw3oPSWmsKiLqh4X9PFVLt77VFDFumnJi2j50
nS0Ecrb969c0WIhNwDLZzEpScByDhsohquCzbJTz++ZIfqzNKs2l530tIMB8
ksHzB4oKfdNGsT77djaSHKVuF7CjAkFhpgXhMCox8ukBO6qDNGS4SyURqA2w
pEHDJbdS0gXY5jNnVJKjiq0Fx9uR85XJqMMU2D/BX6rLq+FVadB74hxxj+dz
YypyxcUZE4UEYD6FVa+f1s7EGTTE2GBXryo1E2Lq8y7WcZ7Xw8avAvDfyjWs
/FqUVnGpW71e/xUvHz11PB0g9mdzy7IYmwiUvMWgTuhS95Tg/5YW9PT0Jllx
nyRWMDQ9EI+VJThvR56OQ/N6N5KULwdJOqG+fzp5BXXYt4WAIPUQs7u/u1Pn
P+TZMAY4YqQv1GFnVg4FlOaAFpGE6/+RUrPL9xKQ3AMJjNFaTwK0IJdqe++N
uzMkLceiLI/AJkoQEN2+VxLsEV5X8W8V7NuhHvEkEIS8GoXfsuzJSho9qEAt
9OUJzxUt3Q7oWJkpxylxhWLfLIJMVYNRrj7UllOiATWlVEkXF/dsENLSO2ku
EfWdaEWxX5v9A0/FIn5Rvit+KYQDy9DkGyi0YXC3jwfLLgf184TxW8pOSGpf
u45eaOWSV8YOHSGjEL1jJNDcHLdYEgXcVYJ5rN6knHW9YT48zpFF8oojColH
4gHC1CF9KFsjKTdTlKKSk3gWSuguGkh4M2LxYJZMXZh/xAxutWYBW97WduRI
CtJf7HBpv+yiifBbDFMtBPCdi2S7a2wbaZoEki0hKW2SB3vo8/BZHLuRgEwf
/zVgCfurdFNk8YChBdgMNjvO59ejpq2YCrKutZcrsJunInsLsErMga6FpuJT
YfJvkHD7wOQqfwftb5JJqB434NubkgrrxPGB+r8mMQsSPGLYs4iMTbQk9kxc
hKyUuyXLQwTtKSZQCXCUrufQCt8HGAxyeIP3iSsJaVLFRwDjMuX/7npDrDCh
OLSmNM4pBI2llkW3JoJqbWSItw1F0Pz3ZUV4gUoENpdXRrmcOaN1jAOUSYoi
K8brSxx4n96QuZtMvyoWaKa2JX9qr+ZghMw3q05Csovt1eK+02uCKtsRMDId
G89wNUqBd+xgc9o+Lou1RMVO4D1OKyTJtrEjZL+L3cov+CKZGdZg05pAcNQj
8ykNFANZu9mZy1zc8WmIB5QoVa7VEX8Os9/Sdz14/+zhaVE3MCco5vUnN+ih
qi1azPIAidxBEIbgQgAlEHHG1xFs24UdWbk/zs7i5WIw2vmSvU/SgOWezTdF
HZeTreX5z2hO9xSDLwFenIJlEFAW6FBTD62+hg3HrDwEkxUq/9NLP8kW5tWo
beyWIo+Rtn/hi0cCbfdEJDYdRimwSUiYiCztHrN18B8B+2/6p2zkfiH3kIF4
ugtM1Wct49Tv23jD/o2LdkJvTj5MA9xp/4cpx36FWEruSw8bBbCdV+UG6wB3
gnScEc5jQ2iHXSKVE3ezNzhpr/vbAqwGIXjDK2TJGx4M9ax4Uw/6rhM4GbPz
IQgZ/tVjgmIRz95W64BOyqkoTXH8TuNdjSxi2Pmiwll46hCfZag9CYI/gwKI
fgRyeP9HWKDSa8v1qSa60R35K2IQqJdgdmLO9wHvP8rKRWIlcgewm9PIt8+E
Os0EWUW+BItIEJyd/xyyD/2Yc5RAHCwr3hDuuBXlx1aYFiIa7FVLrSyNHM/X
MwRcAOpDRL89rQsWaitllwIsKFWWDm3sk5K/1DLYewhaRsekjbHle9hZ9o2k
F1axGjnK3Q0BU1/ZnFdzQnW/s0snzutnIQuJkKQs1J63PnFqn8B+Y0PTdupG
VhCNefsMToBwlSK3Q2sJtQDiOGjV+eZf+JDbRXrVFoTNrsKRG8UNOgsMyLB9
2LXvV0XOAaBNnUM1s4FslaHx2wDS0bywqBLGlp94MFi22CoGZcnVyOjHPgYC
gnwIyhyvG3p5n2Y+77H5BI0tXYYAo5eKMQ53hVgvaskWCfaJ7CIKIAIkcQ9d
DrTEytEyu6Gk0USqaWTD/zDhjbOpwqWnUKC9BDwJd82Z1HO8/f94CaNFQQAr
hK1LpSnuSJz5U/TDhitonPdErfmvtRgYifnvtAlqzDWA3u6XK1G5RjasR+WQ
aydFFOxLceAiC1hg72zRD7aCMPM3lJaMKU/AZlOuGyIYIeEveemmzBdcASkQ
AsgIgmTomBBJtqp6JcL+2MNrawFIBmxWEH2it64ATmcEQYD0SM4IrhoGrYJN
XJrs+TiSVmW4LP3/tccUszqEZ95al/iBLmVOux2++4MoFsj+3dvDk3CjOQFN
eJYDsqRX5QdDOJwc1x5vf29kpRT3jSi5yWLguJ/lVJZ3Iro+56Jp6vQhGaYL
l+KWrwoffjoGGxO+EPkxvR0DFVG1ouiyYpssivpQ+E3uFgFzrPkGQ9itF0on
JbfFltqSRjIVlQ84Xwc35Qrg11Znwu78nSo7YWekTTSCg2dDK56VnM/19Zna
bsG0N54cWaGARb0biW8cAW+aQoeeNOHPXDdLxwXdd4UpK03h9yVfcsELlbsV
CPn6ZxEM4wYkmuv86w8z3fg197FIYWA5CJmkrvQ3pzVOP23u1wHcDONYWhBs
/HpACmIcQ/nHWAjmM+0gYSlBC0wz1GjvzBHKRjODiSnE4DzWJhEIrD2VmTpu
r9+3DdDebgpOBD6V0UuoDgIurdPrcBv1LFD3g/ZuJM6Q5v3wwuJPXnR4YTyK
yX8F3nxrkEJYTriDsGkqFfJy4jW8vHjgEO7WnZo57DTbfbVsal4s97MrO6K5
VwkBwPXRcYPr6ELMdDw76MKPA8D5SflvSCzRT0lsPzb3paymWILtmlUUP6q/
rD6JWAhJ+QeiuJQtEJwMS2kiIufLtVlU4nde/46sO3XOlZG0lA+5MgMSpvx6
ANGBPCibVPjpfMwA//0T71K8xyswQSnbz9/SWly3n1olhufZSLgOjyvZRw3y
v2FwVczoZuWFpvUHO8BsyoWrgwn/YsIFZrIMngvCdj0m4uk3n5DmheBiobGp
Sk67HFp9XHblJ1mkuzwuzE8Qlsk0sVMkaogKEV/S2zmGl5ycP1bACBnJXIHH
MlmzyNrNT+g/gpl2pf10C5EBweJHYGoXEDLU2diiMZefg1qOByfpKafASW43
bNqxOCdrvR+mLzkyNRAkJ7oqprcW8/DWU95ockoHICZDUXlrRdA8RB3xE8SY
c7i9IlNMZX3DHUSFpymq6JpBwdH/D3IPbCdeWj+xqjZfmJcG0gXWijiseriK
xiy5g61WMvcqKmbyYrvxAz/NdMTl2J+BftWBa5HsWCA6lwYG4bdwNIbLEVKG
unGBgv3AAa0Yz/FSli71lbUCQb1qi1rG+6UAxM3cG/FfdPIDhvpZkr0vGoFf
/g87H/+CifDAixLson2MmIZeTObTaUWadohMPhUSv0exb1d5DinGW/sSicTK
4Ju7xOlYsDch27lQCDFRoIe0IkKKf6F2rRtLgAjSY27XHw5vWYOq8YQaJMJM
IHRGEq95OrV9uLCSo4dXfeg74P8IhuR2uhncFMF9+dV4AaqHxduRQCROWxVT
CpNE9FrhZ09CTcOdWJWmVw1jVGRZ7ptXj5UWjqTppEj3ybsi5q/oNUm1J/BE
suD13OMIJg3Fa8N71FjzKlXLRWiJiL2eQc2zpKGkqKaEpK5dj6Ntastl2TmV
KJGTtTyfTcfx2gxvfn8Zq+1oLFb29AXAGEcee5efM8nF4l4dJMgs/G6ghuQD
3MQ9tSS8rJrPaDbnF6k5gCY/RUoR7PM5lV9FJJU2ZFRCH3WbNYcXF3zwVHue
NcHPWmY7PDpxlgkOYm+QbwOCms+tIfIu/+E3zHvapHlEWHE+1/7EcGATghU6
r6t03ej51GIzAS2d5BGFW1F0SKI2JhhwCvCNmjUsdU5TKb9Z7r0Kf6r32VX4
eg9tk9IkpqiV8h/7ohUoOvR4s6WjoyLBMY12m0FtNAMr5XyFQrJOAgJd8aoH
sWYXs3UjcFw6YuJDY7JYhxtSfBiwIKlX9PatUTZd2JbpJh2qymT8oC83a2BX
l5NbjjMpCQzQLo4821+sTQwflkXQWrLTXg2yR1PnJ7WBrLPKV1Bd91mI00vd
xsAC6pbDAklpogegQ+a2KVqy7H1eyUbptJswUbyZ5sW9ubdE8F0agSa5zMYi
AxJZDVGJ+nMg15/4mxscUiZK8WisBGoFkPW6FRTaHkpbu3bTsLnxfS6m2OYo
uIjdcbm7i6hKc+m8uD3Iqm3NoEdOTm4xmn9Eic6ycsKW6xKH5xYQEkIfKiVg
oBPUjfr1dfM2aL743v8CL1BejpJjjQ7lfPUCEqRWh50DRpPRlhsC4/Z/Zi4i
Mo3n5w54yEPxl01kLgtEUcsQNdR7DKkMXhP8gRMwzXg3BIsgLWsDb4bA+n6/
FKOSRJlDVb+Ct8yaBi87Hz37GYum1IKvUDyBUaHronGyum/Q8SR57FksSGg8
2fp39uttK6q9nTeIbZceUZm4NdizI+dcyvSlUduTOUkOeOemQvBCxPTJFyAo
ndeVkFr0MHZQL7T1Iv+1eCNPBNWtY9fEmfP7c5ShKnV1I41tDieZJPy96ub3
1Ep0xlbQVexy7fIzVbwWkf6zaW7xOMv8hGGZD26eyjo8AEdjymT2etoEA/0n
czYVM/mkmTRBLg25uUK6pBJMJmu5DQQAVGtb+O6PFYRfgQbuEoxhN4PdCRfL
nNrgVycwl+NFifvrHW7Ok7pjgPL0JkQ+iuRdvIUNxkshJqgT0IRY+V2CjPm4
WVdZbVCPPkU7z2FD3fA3rTKng5fEkwWG7oN6t81N8+9//edsrdHWt5rTuPX4
nYtXRAapbA0lB16MOqkIFLP0Y4nW8YNPWLs7EYXMUOwxVwtmExHhFsQZbkeE
6YXolJ1LqOqqXmPymzC94ARLXsYfuY2TeS9jS1cdGj3K6F92CgQ5UKdMZtIv
s42qUrb8jcHvtuIleTzUZ3XNr0i4mCFkJIWjfh6qzp9ORDDXy/baNQBc6z7A
+EwRDTNV5M/urZ29RSzcvoiNldQDuuSy2lSMBWm3zh3A7Uv5683y/irnlZ40
5LKnwVy+uS+2sZMNMwNA81SsIODviTR5hWr9fqzdC2Jw3oTajhsZzqMl9y4C
lkOp3C/r632WxvlpkQvTR9MkjdyxaxdqQImDH2LwKTAl8UKIztaA0jMTgu86
i6CMODCNCcrb98xDSt9QSX72GAf7Lku+E3u0FDRzwIuK+GiPpv9S8ReGpf+I
VswEu+yLIiTUgCRs5IiK6jG8CnIy6sIWN8ozKJsiVSBz08BWCTirHknJH22U
TSsWyfSFw4mRY4VBEBBMsGnMTLjxCJb88Jdi1vXjA5o5jD/e6CPC4fjulkEc
e8xufo36kFUtw74nq9gkuoHDWCTezXee00aaxKKcLkGlJBpRmqyhW/r8yrlh
gkBxhwYJ4Ja7xj0z0P8/yaezeS2SxFYNmwFi4FL1wW1pRnO5AUUwE22evGcp
zI+MAmynYuvFvI5AT+Rkkjw7xTQbw8JJfhB+i7pheoL7qNhmTGHldsBjTGyN
+G90bvltHV2/9+96mTWUIKzfdQU5A9NWiV4WlGqYknPz+w9hjsiruqBmZmy9
6FPx56keQVwzcNkuydDOgExmwgjcfTEE840C/AR7k2IFf1qbOZUYQmkgVp1Z
NS65aI73O4WLgLVc2d3J4dM8JPPbsQ2FJH7Q+kgynyb1g+5EStI1TdF5JSVO
gtI3pgS/t/GUqpjNQ8QttxUMyawES4njC1Gotf2YJymdF2lyV4g9PB4ilpMi
l0bCEVqJ7WabsUQTOtjN5lHmnla18R1bCnpd/SJLJxDT2gCoqOv9cNMyIxps
Zu6kOLGuls8waZl6xI/eLmtjuPcoO3cVy5uBIGFrykYlH9eH9JRoEhFTkNTG
os10qOjMFQrabmgOicksxw7yGnWNfSvz/cET56nmEB7fhGfF2ET4xunKn7HM
JRz1sU52dZgsQ/Kkcg1j0Qd/gggm+3n4GaGNP9XmrAsw6C8vpJ7NIrAqYAIz
PGZ54hXHyCCjfbKvdib7Ut2fYDiUkUAsR6Jnxd3eMVQ/LXVwsORZCkS17m8E
9ihkYSMgxEusH/heLeYpKEXWFR9+KYPZVvnhqIGH0H/cgf5UM/gGN4q3kA1i
68qVjV+uK8lkp5kNP8okbNxnxmxOJHT9bpW+yTppD1cmuCoJ7kep30l05D8v
CJz8EQk5J2lWQuNkuaIpdY0WjuEV+tROWoebuj9EQ3AjvOhdHC8z2N3AcNbc
DXcjurS7HsPtuQoLIcnLjQSUx710lpzhWVrCB+X80XxW1ShPTmD2VHoJvgXB
YuCn3LwuhMd6xfhnuCHU2KIfM9podjs8zpcnFP8Xl3KU1WZdh6soLY3ORmGm
T4hqgI7xKxS8Rrh71gCPz1g739RGEUA33lXkOSgC9J3UUKtv9N8kiLMDlQlC
jfa3tuJCT89K3spdAy2B56vVN88IVIur1yWt3Fq9g+ESpa3t6jlnxM8HYv4a
CBqa7CG/ui0CLp8wAO9bpk9PmMDenT/KQmYzC9ZdAhS+U02xgMXmp6BZEsPj
KlD4Rpp4cudDmihMomT9KcOEtm/nIRxPWwTD6oP3ypxSgrHCT7HoweB0Hkb/
Gcx4gvxKu+q+6brFM2daQuxQXkJd5/C63VR6B33gwdX/rpbDC32gGfMZqVGV
HK8VSANIyE3hJs8S7QvHoOBT+UuXPqXkzxFbABfINdnvSiLh0R4cjmWwtC5o
fHFE40AmWqxFHwah0X1AJ5FNTqzhaGsWngobPgyUdmoXUHPg3QF32V/eL2Xh
pDY3eTax/1YpN+biePTlldXoLN0p4mga4GrHe/lWbtz06EbwKWLn+TFSaPsu
PE2LK89BG7Zjdgdzz19QLYl//HEzf1CIRZCUMDM0pjCDeXEblwliUnwpymfr
GIoDa0DXLOKhwAgxckwPfA6+rhyE0/nLTBjilD8LSHtN4lnJXCg5H8//QAku
v7oraUGA1ArTLS9pZjvoe/URd2KO2hqHiqpivoiL9NNBQs5lqJjs4nJWHOAm
aWdTHrhPR0YRRD+yZPD7C5RI0XvoeAccpsgXMtgPxawBneA5isWpMbxQyirh
GDpygDXFOq8Su9zs701WyI2M5Ch9c1PdK4SJCIUN07tblk5aBFINIY462gQB
AZ3K9wpoEEzsn9e876/f2owBmtq8pwrDRa75qzdH+dQMkcN6DZCBN+RoqTBi
aUj5A24aZVOLq/GiL5bmn/lrL3fgab8qUBs+sbz1/vCLydfk06aYBDpIVOnL
s1cn6pk7/6K+qpOxfQyevCd1Uw8ALcFNAbJT6MbSflG1css4lZfSYNXVlrVl
9mCevtrgev4fR2m0gU7rgxGpTRLKJ8h/eL+7SyFP3fKQH0s5SfiRI07vU7WT
/kgldAkewNvtJRts0mpD/zxBtufFO5/WuRgTYqTXrHav63WLiSbJtUe7PVL8
gTzfnsfinx83vhpHnmSkPAJhwnAv9cSYsjeRKPj1KQCzbJo6ODihX+34ctIb
w1jupDUXgjY3+yn9wCou/++VuoS6awp8bhhlfUTOWtn0nu3T6ZgL5B0zR/mz
bSwWTzm0Naa3wuwJMkMvucOBmRZNU8WG7t+7MaZUwf34gbgybw7hcVe2KNuq
+/ruG9YhrkST7MOP9DLcGE8Pvh9IqsLSoV9yzsM+yuqkSB5d0R1XADgGjUP1
opwLEUbFsB9f/3n8yCSwWgeLieYnQkhsBKmwlRLqrf6AiJ4GoUwekIJn/gKv
24pOaYsdnHcH8ZD58gQA5D3qby+b7lEvpVap+1tWsDpk/h0F2jh+2Jllbif2
qIjPbVcryl5/7Bv7PTB2LLgn2i1BN1QxNur4siDZK6bl6H1DqKbtZxyUlRnr
IYF2ftHiK6O1VYdBxAyN3ziH0iLOxeazN49ni/s9JMqKpQJbj626+3dZWPlj
427Mka7XS6kvjEI1tyjK2qrTl12TbAIfPE6q2oKWtzvT5CgI1v2dN//eBxwL
lVazFwKJHakGvgaFr7Dh9kfRKP6jLY5G9XLgZw7YNBAPiKlSHD1kmGp5Wwi6
Tcv8KCEIjXbP8BcqMRTT13wMzr0i8iy6WvfpNAhV0GrUlds3fIVyIhh51YDP
opb/LxIL4F2xK85vQXtF/93/Okzob7ULushaaPhhq1DPbREaCVGoQx29ijFN
YQwqqhteS6IClKMCyQ0OeRVkZUoN/VfA/GyhDnXjvulf3mEY1e053QjIXXHs
NDl3Y8He1MoebrVCEI/fwOcpLsdJxKP7nD8q51LUNvk4DZF+6dH+0VqxMULI
kpGNLkMqRlfR2lZvc3mijCnNUJOwR4RNC2Fxlyq241Kiky5i24dd7XdBjQEt
uWQF8GbfIJ4cTHyUIU5+N8X2ln1V2B/DSj3DyEG+akrHutOdv/gVJDPobtM5
zoj9dHPZ61Sw8xWLD2BD46y8PzR4j2msgho0oIj4zlxPG5yxcOQu3CsX8U0o
VPRWuJdUAvKPa9UtJfPpDEhLLpZL58U9PNNw4S5dFRUT/N0Hqb9MNvxn0x2q
QN4jJqLAbiHRM3Uw9rbzmMOIPxH//2ROh0QKFzXRCL/pP9aO5ummVaFK8/R3
bCwZOmAZX8WDWqMLWBbQ11CFwf8vIeLg7Rn0Vf4ZnEImjvhsXMRbRqAqxHP8
fnR5ZkoPiQvhpTTfGv93Su2vvkwF8k9RHTEQgrw6X8WqH4tp5kb/BauUUM5C
UE0Yt7bnKl3cyjYwDhI6xWKgnJHDGbSS1pROAa8PelGTee9phHQOcztoBOHL
w/sBagdr1O4sqBjq1WRry2FU1KO4j4UzC7qxLMINpx7Q0WwUdh8o11z+Gzdy
GVMtLj87facspEIqcKZxqmYT82Ln17mRaV+fisCiTrazK7nbpERcEWCKbiol
qZGoMHSzmWhNmLuq+w36NJ65qCm2Cg+IK6sk7h1UnKhCgc1fYExm2BgQH8fG
4E2JRJQQ4g13iK02IZ9xt1Krxy0ytAiPNRgF+mL82C6Qa2an17JA1TYjFHvT
OvKssVMKtbfhr4TqXzyNNuGeMNHdPAf+ETQAfd/c8NGjlvN4l/ahtaV1Lj1u
A4WE9WZhSmqrAsFJzZy1a7hV8f/Q57AUaPpSEU/oohwzapcu6ITps34Ax7zg
2O8isP/X7/nMSVH0O31PSCVFIKk9YBUh4sNwLFcaHTIaY8tf5X80Ul66vpRk
hx+kui0fihjh8Le9usd9EXnnvq3TPG7Yo3AfFdrtgoBzMdvDHvI6sEfPm4Yo
zS5N5GeBaJEzGTrFJEH5wuvmZ+dC1G5IULnwXBHwX09jAjzMsBe3UBIr6nq6
55W2XZxROwcdV69y5S8WFzcGjBH/S7YTZ5vkQgk3bb9HFfG8qI6a91+AYSVL
SkElkUUh3Phy3UKRtzdEnbiBq4aZsFnypfD0r51fQ/JejchKLNDqO4xwgxUg
W5dhFUG8f0tJss7hqusN5B9BvzLePXygWz82SW0A+WlyGL5dYqFz91k8gT1A
wnZWsPv0xzWwMPVNTe6nwcYdsW0Jkhck+dPEX3SdLDPvTsGjBpdVUZ6uMO4Q
a1fm+dO1++/ugkYsH1oqI2VHfixmESSS+qLYH/lWaxXf7cz+O06ij25Ml+Md
ag8uQFdy9kkksElx2fvSfyGm1U2RVEiUYI60U3tK8C0CBajsQxRAzb5fT7n/
BlS0UG46HjjtkYjXBqubwup/BDBuxcha1KTaFOOuGTcoKFGXHUCyyKG2lobD
dYKyl+rhDEtB58CjD3fZMvseCrnb6gkgoJDoDqSvZ1je1ICX0NshczKyIyqQ
jo1wJAsfuK3LYrjfaesOdfaRviHr+to3MHr4/LagIzXRkwLaN0GqxAgnIqvj
2iRixYc8K8d/DzU52q8HPqOx2QDnLUDQ1DC48/NsxU3D7dRSC9kjnkI6CnXB
8t5Tdi0m8a4feeN8bYTvwHxVPkiXo+5FuBhxNALJsGjHfQgRuN/+bZSBn7HK
cbNAG6XxYt0ilTm2bU+hLkmQ9CCx/+YTa+O9cJGr1MHAvFO1q7p+UwHYeFfU
UQ9LYJnx3S6opW+l4vngdNAnABxxTG+oWRJRt5K8QZvrV/D4Gp6VlS45O0SL
+sHYbRAC5XFWcv9pmd/PVpYNMMrQvpwV/evkWNk7LIKg6FXwytAaQbl1ZEVb
YPYxvyPZCRpkhNoo78Rh9d9X3hteIifxe2wSc4yFfX7uTqDqX6xevEg4viqv
qFAeDwIIi+MGgZ5TYf2qQbkvo22nAoCBM8RZ4o7UVfr443nmhFu/64GJVVnE
EYJqkuq9Tl78FAOGhuPgjbcGqQRyRNh5GrlLUl/GO2Bc3YxReEiRSTgJJ8xj
2HFGxGhYrNfEKvKwqrR1+fW8cDnlAUqnYYQ2jWWqSu2AIo9TB5CEdeidETSA
9JtO91tUoM0Jrm4/grzeoAlXphuCTyvqgr9QodmcJFUXFnMI/cJnbwpvby4y
XE6n3IOAUdnVh+VhsEU8+Dh8YyoWPTKFsgvUgflB29AQlY7SFXJR3wc6uyDK
2yjqfDiNb0EObmsefZqJXn5I1eED56OydyvhdAjlh0s32hpqv4Cm6XStpLlN
5kbBB0EcdvYlrMI1ozMl11Q28c0YgbPd28DNyXId3rM4k3vVhtsPNupyCdyo
37h/ylNBgkWp8lFMXa8TxIF8LZjONrWsFLWdboJIPGwsw89yHJWF18CBHNln
aLW5AFGBTqpVzLJbcF886Kn9eYdflBgW0neRztT14bUHkCjPVok24zia5RyR
I8m5zyWRasUjVQwQNGa7mvrlnM1r+HQl77TZ6saq24k3Le6ja9n3pNn8yJeL
MTodBJIDTR5kb1ls1+7b1yE7wdq/fpeU0A95Kt8mnOGoprwLg3zna1A30Qgw
tKzX9KgBJRd8xCqr930btHSMoKPn7KKVsXc8LeUsI1CzPsgOCL5o+O4ZJtm5
+Y/Usm8h82uWCndehYNYobIeYwK355+z4xt2CC2opvAK6hfZI2wB1hUPUXcq
ZneBglav3UI/iEEFXGPO14evdVH5mYhADr5BMXRbIJLV7xrtOzSlRRJQcRSm
YAOZh9MEGPyr/9xHu9OsShJAgZVc4x00kYL91G1hS4aKhXdhQ23AtiVev9eG
ijbBm+udu4Vsqqpbx93bNWkcgfZvEnhNNsTSPdNLgcw2RkeGx6rX8kwm0+ju
v7pkGjDenPLaXgnbPILEQrVwSuclc6W2zJ+H1eX6GnwUWQx4sLx0dAnTvAUP
jbmErD6FkfslFf+6w/hmm4skq3Yct/KP1opvNtelj+4MXZTTxW0uyT1PicI1
eEXqLEfmYTDOLr5+TV341MpvMhNt0ZMN0LyeS0eL/zt8bI3R/m+G8IATeKj4
mDGwYtVsk1iZ5ULuUHygBaYIPcr7hXyLysfnxpOEh9aWgD1PBqoyUinXPkar
DFz/q9wghGyw2Nae6a6W1H+CpVmYHb0EhfpkeKLra9dXkUADfm8eeFg88LMw
QapX4EIGucnK60xNUPQ7iGB+SPZnSNgYmPtvMcAiYlRgMpzhLGZK5+bqFNBs
C0WHr6QHm45kzM5qQ6mJsSFE6YPDTbnr0eupXNVTQHISXKsFuWe+cyC8md7W
KEL9QmP21ItpA9KWbgg6kCXAZ6mUN6/UyvKObb4sqOL67eclFZzRWOGBcfrD
M4WliuyGyCxcT26DjOCdFTHd/bol7+0VPdOEk9oaIfqTIgS0dYgDXJXTceCJ
NMW4/ojERkuRrvYVHfmKOxXtOVDD3BDWTxIOHPotm2HiKoiLjm4/ZkrUuEaf
7WD51bkcnYZnSKubi+rc/rlrL4ovtf42iOZr/rkXyyiavtJDPWi5TPuX3TOA
1vuBSojC9bch8IBmHZX7Mnb0NSj8DTN6Ztgahw2IDHywtzxWb0VAsUbGqKDu
RDHXEksfvcem5uZNJWTsSLHsL7AzRWuy7DBe+iwwgGanTVJER7XviE3s/R7n
xsTnNvhWa4dAvoIrBTs+WtsgxJzl8fa9FTa3rE4/JYdIbTtG4clTwcMPS11G
VjDN2kWIhySInOvRe02Qo/z1B70Dof/OPHPVMA0+MwfasX+KLxSLYE4zM+bV
tpJ/g+5Hs5DYoP/8BsJWgpT9ahkzmzS1ruinGeTVpEDEp+7KR6h3p9Om9xDm
Zf7LprhPqA94pr0WCDbLKnwOQfAQKxntu8MNKO3fDa0kzdVHY8rZ9SzbovS2
1qReOT/UxZjF/wKamdlRgohyIzlZ3gwJMdtR5VOZ901plW9lXK1eSp4ride6
tM8ae0qjOu0qlZM+0SADdRjio5NM2kMTycY5XuXYdh+rAV74v2BUgrBPYLln
lXqEsp1yK6XUOAYc7HHMqL14N2/ohYR9HfJD/lkCRw2WE13JlC4dLHedvN+M
pElmpPe4wHB/jiFL9ueIFG4bC9ogvyCnjh/khfcnz/saR+MbOOz7y8uf6iG9
e0lME5Ksq49lmBA50zAywGrlbErF7zYkSF2LoG6h7SN59GnjcIykPlL1PJ6B
ugDKpXpR+DWanjl8G9tyVY5ZKDgcWU2C12A/XAaNCUrc8pwQu29wFfbNmlus
N7/0Hj2ikMdYawVoSfm3jtxN/vqiuZ9r7GD8z6BVamYDJk+SSo1rXlqzF6Z/
L1qdyOJgK3icsd961M4B1lFDAaH56zsmc+U9I7xVkzMnvGFUqYcdo0Z4xAm+
v5c7KbODGxCf5Th6ISMJEw4vjJiYWi5QFqAkaQhWQWQIurPNKomywcAkNNg9
iZZpYzk5AgBusWohSYeQjiDCn/gH5wDuEAOuvkI85IYlizpuEOCAN0cY9JzX
NK4E0bX+s5LqVaezhmYM8Atb/8EkhcsQtIra+bSnGWII8pI+tkWwmw334Kbq
9PQ5PeKaxCCO8gLdIVSkZdXq8yhC4mLLrmis823GyW0irXv8IxZeivUdZPA3
+j2CpsqZtoZzE2fRPvXAg1tw1FB0lEbaBq5lf+eev1JuZhNB2n11bzx2ClPJ
pu0IXLhmsBr1o5ts8J6eOIfiTM9KvIEdEfqam4Z44ARHI9tppjK1Z9KvcORE
VtyWvI6qb60NQQmlCH5Upms2pdCd4KF3picctwXsdmCiVdPDEPfdanDsvU87
3i9rwioB6pGZrkVP1jWyw29UduFtbmwUH+FT2ajiooRv/riO9k1n9SzeD6gB
i0S/LkG8D/cw/LujfmIB/6kzjb7++JhjWtXCcXbAkhtrkjFqTjWPjxcVTOzg
jCQOUT9c1JmLulH7/WKRlOiK6mkfXI7vAVh7zxg1DqsA6NOm86rt9vomXK1t
iZDIPpNS2YZT3nXQXDv9+5EPTSs5Eb0JaFOSI3ZlzxyUWItKxXseiMKHy4hU
lYFD8LQjgbz9eH2tCiqUTRhM++09JmEdSR3opn6QR1PE65Em2iT2G9XPr3qi
OeslzBzFawVFJhKJvCw68ljUjGVSAn+fGaZqPdvcl1WjiNWUgmeJzA6393mC
lQUphBO9fx3evp3XQ621YEX+ijXGE6BE5mMYrbuAbRKbqW2kIGkj8IT79Ven
+w5EiDhlf2g9rmababSqYjG4feRxJMn84ZO8dGoOkkHjltfIKIlHcLY8iIzM
oNp+/1cQbpf+uubekGGx08J15lAxFse0B1jF9wK3hVTx/S1c2kjfADIoJRjf
ona/kcJRzMR4a4oSXpdcPXFxrv4dua9DsknEwG7DZPq26vf3lgAXKJY9t1Az
0/jWkUqzKttFIXvHDmbtFWvVN0n0WGYIy40r7pAJIHThNmjpd+MoFjgnJXOp
z7lTE8eJbUMW7/pOuP1SixEi/QzMQzHlXZEk7WQoKgWOy86qg5Ihf9Q2QpDi
EjKENFxKl5gZxWdml0zgOtvYRSTjSVtQecbtCpUa5WEpURjDYP1A3kTPUCXn
BUc7XE4kgbZd91FXW7BriQbSEcMjpNrAj0cOLLC1aMJ/wbTeG/BBhZ96fDUH
uhuF2+drbbQQ+xQSaqF8xE21RHQz+MZblbfgmnZeFIg2JnE1fZEwioPGWFWN
YZxmc6vbBj8inlcxvU8us/uqraxHHMo7Sq3VG0zoxcW/tzu6rxDE752KAmvO
pJtefQyGAE7zne+q0NbtjrG4LVh2jeGCBmn2ISgSw4PH01GROOdYOrxTWAan
WRHZtzubfcFd3ug2ncaBNjXwNOie0dXjNVgQ8R9o9dtrmRAdwjU0OQr0nNUS
qaeI1r8er3tyiFk0yiAY8z6+qDLhOlHFyzZ2go2zwezO530tjn5dB6mptbrd
P2maIoUdroa2L6nMTD6llKt1dMvnO9MEJQj6LbmV+Hu2yKatzydiF+kqBkkf
O6x/n/pA9g+5wOkL5j/Hso1QWklmAdpVGRGj7E9yc7VxsptIO0q5fFC1r9qH
yrVxLUTuMg0iL3ef3irBxYPGcw0uzYqec/DdgUpUJdqcC9iCFa+3Cf7AP+mH
d5V+AxK8Y9+5SsI6udi0aRnyPwgxXpvbsOTrjk9mAM4CDcQkGZPRbY2QdJm7
wLjJA617sB6xzntmGDVrrraU/HCW/FnJ22YBnyvHNiw7lfSn1e3GqEFCdy6l
27+PZGVvzLsA6APD0+2v6kMGUAJgQ4IWMNShojy8434unuIWGCnXWAB2pKPi
hR/dIW+4z8wKuUcAJhfMfSF6egnlMONaTcSaJPNswbk3Nwx/ZA0uIV+FtzNc
XcdRvsROt/f1P9HgbjW070hyjDSzgu3jzb0siQw4Y55MbariOo2aUwJzMDHw
MyzNJgmjjCTWcZD+D8iIQJeVf+T0psoMMxFubnFrfPoC66b2KXA4sUGuu7w9
IWC42lYVuKNku7A8CUsk/4kqWQPR5wOQWeN9U3hzSV7j/ORr1LU9MOnsavtq
YSvV21sR9M46ttO8Y48YgLxZ8SwOTbqjINBwT12YylpbCvpQL29AL//6yhhG
uwi8au9Enw/56abvf0LFD9HJEhffMyLcgoT5cBjQhK6gfW+X4B9mBsSB3UpB
2GVmhufV4Oodk1QoUcAFhillP1zgP2+AUJcgGavL0oDvmUODIN9Mp9W/t2Of
UIXEN+O8c1rM/gpCxpiGfWAMnOg2OLvxDFiLXsjQ9B/dY8qyWBcJhxl6tZsf
hXT5a4UtuHzTX7t/14VH8ucPeBlMfHE6RAZUPZ+z3/swKq5fwUPG4y4fXfoi
JvScTWOqkfFsXhBo5mUvrdYSc1z9t6PyRSoT5D/BwsgWeuIE64xzKAAXbt+A
EWMw6LucI027tObUoo0rpEmdE+WbfWVvTecSjs62zjiDFtpN2l2JDYfiv1fz
WT8qm8jcwfCRee8GN8oMLW4wGsYsDnf8Xa3hAwxSM+OMIddW+mEqP/L1lNJs
wJgmUQjiPR+Zzvth5lDng+LFPBW/GRpVwdguMMNeiWlbtwIReiuv4UV7DYF9
bHHIlYOUkFgBbqY8EaTxagoSY/8x/lE6gUiIoKnAzMmslth1GPWdxaFl5aZZ
9FMUSPmI8dSqQ3fCtwQdZDtU+KNGnZYoCQ4Cw975ZegDSXOh4pSOMznPhBTi
CJ0UE/HAvx3KsfblN3Arusz20TfYkmOJGZx9y8vMHvQVkbd4hnU1z4HSd/Yk
smIbszkh0Ii7IjOAtVua4c0I9Fp9h7hxkXc1e9xB1CfOXnEOkx8Ao4BdCO/P
OwqJNw429nPsoPs+1w+cliJZc5Khv5CU4IF0YKQisE5MQDhEtPYpF66TSd+G
7A3pclTsiT9a0jF5KiHUQP5mFE13WY/bByiXL6n1BMi37TG+Tq4+1JbvA/iX
AuHt9sxiaNVO/uP25ySOv35Cxo9k1WTC4c04ZMm4oBcdal7joya3fhM1gfC6
E/j8Nk5fDxlY17Tlq1DD1jIa5VMurs526JfoGVFgvn4PaS+cYzRKHWc3MlMS
VIPxnY8hjB6n6eaHt3Re2CKAIiHBHK+4sprZtX7ErqUr+nG7e45H5I7Dm2vZ
O54hC5IksnRiwETQH9f+boEDs+OLhlRDqSgqQCifcy5fIx//kgj9vWmMHwMn
338V0arfALPL2AvNff0wTQLg9cd6+Tvqx5BYezitPKV1gqN8iGB8fSgSesY9
wjFdzgUfWzHb4hOenWFMWGPPeb+g5csZGjcN3XZYbAi6bD+BODbxC9G2WjHS
8gmuEBSst+47YkJtMddR/r3hum8I7jQup6R3aXgf5WX2PbMN5czHyfcErQ/J
fV2Z9FH4qrarPJhKVDtoM/di/lYG5cs00xJ0hOsl6JPJGnh5fS8u8luaxhJX
eEZDvjGpeVO6rSYRJ2R1H0CZRTH4KQsD8PUiIazTYHk3PUhFIJqLpdB7VqZR
KtOu+S/k1mFNkEPzCe98zzh46P/JO+sdpIXD7QqWEjkaYFsO6O4FNh++/M9R
4cMr8hHtf7wWGzI6eWnhLRON4OYbgJvgGmCWP7mq/1bPZLoHkFSAOx2UNQSf
Yb3nYcr1vuff7NkXNhfCpW4lleL1ZcdDsIW3XHS4oRMvQW8a5yycZojP7nrq
s93NbIuKlVAgqm029JuPtHXqPKKlmJxhSfXSRGJzW0S7LwpR4Php7+xUVM7v
IXgQSvEqJfMxVUAwnZKC8PDdfIpNuz57IxO2V6DIiIqyD5Q02/ReoDDcJx0G
ReFdSr74vSCJVU0h+rKqh/6NHjNYwXCXYxqgOobboZjq+40AZY32x9COOLzl
Z16bVIRSHmmmn0C8UlWNkL+Kz3w/ltQdRxOIUBzq5/SVimf19zROtNaJDIFz
ycTUE90hIeVjecuSbFb6DV13g1gE7eHKUOr+GifLfPXFlvkSLcCkJjudFKY0
5DkgUkxP1cTjakXkE61nur/zj5Dn3wZML4lz56g2JZ1aXKV/JmCnSGnpWd9J
/rA8f5wUawiEs7E6OWp7m4yok86Al9k3yiOa+mVY3Kay0eyokXBGOB7nmBLq
7LuxvcBPcoLCWUwicxlYOTNRFUny5qpRsx8fJ3gW03MmoQw1OWmiSOypP3nb
eFOmcXgEvJ91fzUowe1yxKTBWR5ClxYdCAuTRdxYq2El76DtCiwic3IqUvFJ
irdpWaFr4T7EAdjsn2I4nNRilc3o9fF2avNT53kmHfP19WrjOixITey+yI3q
OeG7dvIw5l4GXJC3NELRZFU+/4RpFH3iCXMfCpaL8VATRMS3Z+9+aRj+dDO0
KVtNhq2jWrxB80wJYWcsS7CkUQf14ZDbIqrhqxgT2tZVGzW/Yk2Zrc/7W9wK
OivbNWnkuAtwpzYKC59q097N5KXwalrSdLn9fqEMJdUbSHA0nKgZ9p2s25KU
DJgOPzI4J6g/rkK8o36H6GnlJ5neH7lbB24ZFXoIwSMNqC61Q+khF+GwbG27
/95gJVmTK+SDne74/Lhi/p64JqkF1Vjf7GbCigLg33Ru6wk9+vc3RXtBVyK/
PvyrRLjJlm22ftYErrIAXI1EdfQlndaFFGH/kxna52+W9ip4bSv6YS7yRsid
EiG/CLwoEg5HfwIBVULq9P5/defrsvZ+rFR0CQQJCPXZlFT3tJjCYEqvB8Ok
v1keneQiEyqAkcz2gGbKLs3kkzqQrJWQ4gLAFUVgSK8myfSf/R64x2zStST/
1KcvwgrdoXbN2AEIiJ9pSf8wAqgJGS6EcH7v/L2Wabj72epWxxJoQOsglBc1
zU7cm+DxOsnjoxZ5SCGnLW+H0alxNv44Jz54w4F7YdIzbGalhVVFMHxr+Qyz
TgqJOvzviXpJ/+HqLeKY/ilRvXeUOlNjdGtfIque1TUTXr4bAdWDwuDB5fUc
ntdv7/DkXH29kE9xIDNSrUACAHmY3fD9sbbUMuFMFFGxTqoCPgJwE97Pj/ad
1tVwZGrAiZHvDyByEETpAQP04yL4+NtX1vi+aUMWH8z+dRWAnFfHff4gMW/Y
QaXGh+rgxxm12fvBZHEe+o827qczuPJjwQHYr+6UhFXK1soDU1IAE0m9nM6B
1zHLFFhBPmUv9uMVwEt1UpbW0o7oYqJtW4ql+uAWw5StMXOiKi4HlCan+CXB
X1I/63IL+UBbFjKCcBk40JDdOzJti3exsaLES2LLw4Ex799cecGmAU0Jvbeo
KLfeYJj8CVkU2VwmHtny2hCMJxJig3f1/Hy9WNDPXK7jtI1EnE158HR4Nj/7
0SXveRjsecqhJrTc8rWQZd239tfyZsIrI8ZNhCWR71gGnBSbb8wSvWJyBItk
Nt/q/EU7+Ca/9nlIMAt/q3i6A6x5btBWb+LFDeStWO81vspaJou9jBN6Sdjf
eXcRGWhNj12yYMwlQ3jPAE/JPlNWQJHBhFhbGP2ofLYQoR28hONnbEKV+5TI
uUyT3FKMLqUJsa+l8Psx0/i7iaWlDipRrr9OFieV4k0+4FVUuA2ehR6Phc8H
wc7p/0dEuHKP2afK1LKN9trddxMW9eZVDnBgyA+eF7VUvPSItDTgYlQ95lHK
pz2A4JVYN6uuyQtEUfvRvDU++KJop0SqtgZeBm0B7hdG3AoLAf6TAFX3pDBf
J8+AwvTP+i0xHfKpw8p2Tks2C+4Sj2wBOeFCkoMxCte9u/LkzfDYdXmASzWX
ApekNfYHrb5j0Km/FudR6WoWsVtaEnNUbYtBKDMYY4FWKh4Lto8u8iByr1LX
mflHwTXs+Km9OPUldV92TswcBFSJkXwXAILbEk5wjhpmkUxdxW6/pYRXydfS
Jn9cRmZC+1LJbFstxSVsS7vD+3czEhk12KUQ+v4Bd7Mz3GX/l5HWiAZZkk00
xlRYEYyUKtygrUEOHiWi3l4JuLvnRCWx0dNbiG/Y6iIxaCqwYaeEw6Dhg1BT
f4GdPZvD+WHkir6KHQn95JL/azn5mu7AINxzPw6BY8xRVdcoy8+5VO0n4GDF
vZpJfEdLy4whehmqCyAW7sxHvZmuhcf/Fa2rvR10p4JCVgzHXKQ7UjpfzuzV
QNRZ8x3LgkJmIivyYlWSBdGg8ydhpe/HOtMA9KQrBywt2PlTMTc2ycy9KjmH
d2mCWueh57xJ8kSimgcSscF1qINErR474ifHD5+cXwyOQAIoefvtys9jOkmV
5YXdJLHIHGyDsJf2r+Hc1e2g/u9wbtdFy0LJnKDoy8oV+Hx+UD5Wj1Fj/HWi
UabLZs/vv3VhTptFpQ9v7yIo8S9HGhA862jFOxz5qfMElusYsO1Uxy6K5i6w
7Vbbp4afsP7gbCUgQjOFTa28cSYD6/6sfgLE3i3AwoQR5zXVoY1NnVvvij0O
ith+WZZa2UsPVRPQbJTfdwWwoMD8fOHOf+6RoC7paxIbdyZo3EuVGYaIZ8lB
FFbLnuvH/MtEBREIquo+oW0P3vkJZHAkqKeHMHrmOcah99aazx7EEyPE77hb
VGzZ8sr4DaNavQGZdPrR/htgklJESkFlgMeRZqXYWjDwohgNeuvJ7jVDmoJw
I7i7LJ08VTfqioVlAoR8I8d5c3P8mCEkR/C6Q+P2u95S9Sv0kfx2dTn/nbEB
F2FIij4fT5c3pJdyopFhadmL5MS5eWg2iC6ixy0E5Ndr+fZDGF/GY6JR3r4x
Ve1N9vq6C56MFtbgZWBYCOwzUHQLBtZPgeoUN4ux6iUnMe85jlkKHAXMImqB
o94tNN/RXHanJdKUN+Zxmom1t9bfcm0N7vynUniUJPG+UqbxFbvyVcQx+/bm
Sspfpo3Eu9p3Yx5OSsU8wzBY0PS3fGf3dCQT66W2VVKenwMFnaAy9vEWow8+
t0CAxWWa1t52JRRFyE/UM658k2pJPTklJyuUUTMIXyAMjQ72D4/XUnUzb1eY
2NbL6wldQhLeL1Xefh8uzs3Eblx/w7RtklJstD+Klm+T6ALFtiTgTWh2mmtR
A5iYn5kC8GcrbL8D5XGxZjZ9HedKaG1wmsZ5uku2EW+UvkkCbrZfnaWV17ZF
+j17GqQqhdJ+WOg88C20t9m+01++DOJE2U735JRsFwuyBmxvwXhbXIxEsqml
FVk4/V8WUn7AYmfbNCuDT4blZf8fDyOXBMPi+GKRFsb70h9c9xIJB8n4Ta6R
DwPTHMl8Yy8IpQXm0Ese89fzpU3Kvj6P8BguJTiGVoMR69XF/dNDb1YKZ4DC
TSoNKQViALIFf6EaGO8fqlpbvvV0FC8jJ899KeJz+xXcJ6vFUhvf+b5aZ3Vo
shJy9nl1oefGzUUr4AGk2xfrk88WBHpZFhugMjWvmePWkyfIAimVEAjxOgCh
WklmqINEm9uIJZ3bHxigWQnZNlKUasbnc07kZcvtsZHQ05ipAkAG4SFnc6Qx
msrTMdAKO50W31q8TwaFIjWP2JkEurhU5dSCa3SDo6gueTTkKjPJvm23XCoo
5Y2rMPRd/G+zH7o6AxezERwOqp+bfVFrcNhwgS8OSmMd4KxOK4tYpa91gJjM
wwg1+wlzC5OMAvaur8iKYf7nBrry7Y9l7B3cNzd/RBaf+ap2Na7lEldh8NCP
SwH3F6LORtVHlqCFOYQjMk7giD9txCA+ERmS7tTJvdnlrMgyyJKkY92tdVyW
ngOS5FWqvh6+Y6+WsS4mrQMntmVIjUaeHrWqIil5vfwq/tIzJUXCt69esI+2
u/dFkswnu1Acy/KCROohVjn6kKLvny8qG6LhdvMBcBRJ/BQKs3nylfly4Q+T
oTWHk1njPw2UxSGWg1v4Hr1b+8fpsJK6PRbLBjRJe9enuF7JxJGrbJi3+3+1
8K1hDzluYj0WSePqfvKjc8IJfdiAxgG32ahS/uBgjRX/Ek9TGcG0bmJgWF6j
z02usEGjiseMTKu7m6wqVjlhcjlx5xRHiokF1b/WHuAm6L506nQ02yBxuNyJ
lfI7Nv5aBRt8DoBzw1GLfFS1PcujIXIaNonXWDM8jVgEYML20fJGpHjcUry1
YUWa1wRzeEZAx5nRBdocPieYCJRKJ4rHiVqknzXA6QKACAUWb86P4naFYX4m
wO9T3AnKsqRDl7K3bySRW24NLsLBUyqc2LPVTTHD8QooJYo/sLcc7ARFswh7
miZr8SOVP4PXCi5bNPD9l1B5a4so8qNNs6/4ZBl8HoTN3iOU1YeslzqORWmA
CcRp2DHk/i7VqJkcYwW8ECArqrDzg+fS9kKE/fFb0OBSo1uY2XTzkWIJMhlk
6zNQvS/uAir5MSW6jqyCcve54exha8+XxF0TwNYrqaz3tUrTlZMMjSgbTFpt
yEcG+lzdOXJfnfJsEKUQgHM6Zu+Jh7TSl9E8Oq7ktAeHD97lKaWg8Bw4NNOW
+/Mhcj32DrwMkMoUf7ZFvAAux24hIJ+altWaG5BjvLPnQqNOi7hwIrs65kp+
ZecUA+D338qnLngQFlkz4Sq1H0kSY+Wg95GM2ODX4p6nbCl9l+OWXtnUVWTE
28hUa04LIq9dzL2RYJn2c9bw3SIbOGEC3K3hGHdZwXDQ2DL6ccU4vIrnM1ND
6zFtYbv3RYTrxzEUbxgaUNG5WlXWMIFQeYj8HCiLP5hjiQdfU74xBqLgz7t9
sKieH11+eVrusKVa8JPWZNcNA1a8kt0x6YayvhF4Q7N06RnRhSmPIs3s9+e7
G+nraOzTaJNJXsC3OM0RNXM3jBL1Xkgu+8CnB+GrAn12gyMCUNv5qnJIBZZS
vdVKzH9MKezPQ+HDWTtrpHx5NcdG5Fdxs0EnX6pUOnwZDNgSPWW6Gae7wvuV
dI9P8gPFsd3rgydMDBzK0/6YrcEHPq8BxH10m8HbXkDanNFrEE9SCw+HNYto
+A90tsK27t004eY98KkPbbsY4e0ItspaWHEsNfWtcXT0/Knxwki+rrrZ0hXU
d4e1C2xLVbkjZ2TxxWArA+X49kFVO2ZsK0Xf/IPUfTu/99Vtabeyrbpt1ka4
yuEddgVcsM/eshdhM7He1cvOHwpfocMEPynNHnOjk5Hei7+CbiTEVO4nTtcF
SXRhQ4HFPLE1qLC2QAKSiw3oVY6fKSYB4hKcOMoehCjjKWgFr+lneE8L1+KF
aQlipnoeUut1VCOD317rHfEcIdsldlHVkmt1xtLG575vH8Bku1T3UgpOj/Bj
KINT1h5GZQNQcpA1ooBmzM7lf6/J3rg5hinN9K8w85QevMcPjPnc+faQ40A1
Rm9HYvlXseIl6jmMuJdufY5XeQgWYXeEps/Y26YSd7FDvQjBMXSu1lPs+IEP
RazJ0lmSisBPiQsMNR9qaYBh20Kk7G4UIBVU7eWc9FQcRcJ2y533oHyt/RbW
sL26HLB/BKLp6XnX2XR/pMV9n8FkgHcyaDtL9tBRdd+ptq6B2dR+NYViyFjD
vjmOk4ppSzlk2Z7ETG7hnh5r9citL3iRDRauifcf4rDjO7Kmj22twbn+2x+N
am5rArrb+1IGw9cmE9I/CBub2e/zd+yyOG1eBANYs+Z3MmgBvYvXVQLcPP/y
4pUeh8RIy9EGvdgCwgq+ezICa9KTztpp2LkTefntQSkmXb7LrWLJfnJFA/cS
k2mSdamd+I4GCnR+WCCQHnDmB9AW7HxGTO6MlkibSb9dPS9oCY2Sa9/YUWKx
e27Enu+/YtuRZEW/71yqjy4V+RNckXGixMtDrT00dhV4xT/QrpI0zDdRkbBO
XznkPoMWz5WwYHlZ9V4tOiMyIOGbXGQbU7BrDtfo422n3MS9fG2rBhhppK7A
8NdG3cxeO1A+qomcKRevlJbJjBqfNZ7nkNsrY5Y7MtoCoyh163mLRLqQBGrG
XB3EyiE5d/Zif6ZMic38nx1w67Wth87AhJKNWbXF66roHvjL/UY4yzbRGcWP
awbS6oQavxj2z/VDhMhDMyBEwxyUZQH+gPE5b4o/cUXhJyS2eWa6NBIEXUGI
JFMN7yT+6yY1L1uX8DrdLQEc31RJV9C5q+TuhFdtrTvsKlWfspDL/eab72La
77WHFBHnRxZhO2mFJLVKEhRbw6LVRDNhtTn0ZLBlW/pdQgjrjq4XXFuwnAJJ
U8VbVf0KrleaF2Gk/AxIdMz8NIsY0O5B9+pHSlVZfepZZq8YMyQJdhklwgCV
/Pjonp4kGyGYlqRB5FU6XI7fx+CE3yS4krUMqr0XdsIERbPIr90DJITRqDjD
xp/dCXPerR2mzz9MqKiTmgmcYNhgswq7zTFKNz3a9GFfdPlCil2GpZu/JKWU
HI6kThgUNEhWEVYiolXNThtDFVmU9KPU18ylBbXcRR/mqqvAOtBUS7tCmeDV
uAon/RAXs2zfuax9f7/noabXZAl1htdOrTJDtEthdAO1+kQ/gqihewkW5UeU
OYAJO51nf3UaR9HD/6mo+Pl4DrnV4M0gFtEi0+xoICu98fx2/sE5p/UxO7z6
sImqFH+66WcbjjlSYQIEbvdu9C9biSL+PPQ1BoA+kO2MGR4MR4/L+4U01NCw
XJWaEySfrwptWCl6eJcp1XStR5eXIEREXi68NuanzKdO7kUNG7ChXJhRBFKX
aOe1wk0CIxLK4v+h7zLKoB497cZdAqsN/mWuxiWUvIbSCMXD38KCygZ+g2dN
E8z4o62hAPdnDkl/p6tsFoKNVS+11yoR2n01tv7alu6tRITt8p9wlNRSfTE8
G1lu6vIU0E3Lp5LfHqJAVw0Ic7nwa68ja8NtRuvQ04MmVSaZJc4GRs6Rlr8B
188cN+Fje6eMAG5JEmTlycrYBklTNQe01e/I6kuxj7d1QM/tr5pnIZA92LN3
LxG7M5TEHJyx3yV9NPNfdL1Gfh8vUak3gRdBW5p944jbHJulEQuvjLUkhQeA
xoDBPjKzRYZUlzPGSilEb6dCBJlj90gLu08FQJYQGW2+YnQF891af22IOTgY
V2zS82c2o4fWHIMgzqt7NF+vwj1XkQJ2JM/EOMOigh2iusj3xd4lAPTvkByn
PPr+sM4220aXz0vjuztOz9p1ZNBMt79ODf/YuaFYZ6wbX2hMhXQI8u2ECuiM
J26rxaT1Zf4ITrD98KmPb7p0gSKsMExICmV5IA47kGr66WVvEVj4jLvHaGKG
uEs0en2XL+EAEI3hReY4WXYBpPFYrhTuBLdQHndUfOSFh3FWhZ9nBV57Gq6l
+u81go6OM9KE6hBnvcWFYxXS+xQb+OgLIuGIJTXN3pythmSUGRqmrbXZBSZy
MotskQGzhthp+qetNIww6igAv6j5oE7w5QFtaJK6RsXOZF/Wn4BPJYVKmTqR
RGq0D8TerWkqiQHe/2tbv837twKN8Z7Bd1iWnXO9VheBmUmV2/FOJqYd70YU
OWmODulwPHft1ny22OlKQQgv+GqdRDzrIt0kXmsD/SlfpD1U2ajhNw0uDfMP
MRcvvT0EznRqYjZWwIKyvXd6KQ1+/UVd7QkQ2bedQQcrS1WLPlQBEpNTVFXt
FBfhozvUtH6iadLMu84sDPN9DpzT7yLwoRVxdlEqvMKukPXJ5WPcmOxgmU1P
zUg2pgUKZmV7q8c1dR1nuPKLjUbeWyOdyp69Hmngi1VPPGT49UCcp9MqDBhJ
UrlUMQvIemSXsOWvhqe1wDyFGo0KFUfXlAiZxp3E2dGRXk2ur1nRK2rbDzU1
nI8JnW9C8PyAdUQWEz+G3jojIitLmr7s2zPDwJaMyCkYZKYYQXO1VpfSrCqK
xIY9nnYRfu/6lKQxCoiK9HwP6p1OUkWlllW3haVWKq5hVuk9pLQm3vrAKLnd
f9sx0iWxkuvLfE2hOnZplGC4DFLzQZFFhDXlRsRD/ejR7/Y/wJuq0EtEHeBP
tdfwSSwxgOhqzHRSUR87la00R92Q+tv1MGF74ojebxIueqQRd3QRd7thHB8a
5Ru4UPkZ3tn+UmifC6hUA48XhAKtxrZuT8kHdzEybnprINSmOdPdFDFBGwcJ
SvbcR65g6Oxk0HOLpNnafImAin9mZgFhjqrnpOUsvzU1oyQrKKCeAdOPCZ0G
EjLJnH561dNDhDNzLJVUGPptAKu/CLviQ4G7uu94NkBc4jY8z1LGQOnoNyoC
xPBqGGbr2pm2iEbUvcl5KKzQ7/uaP3yAuF1U1htA4pa+5r8q5CJQnBnfjo1h
eu4OFwLHaGqW3yBGNmTklHhubegcrSd3fnbfMTrFfOlhX5+bvO0HfeXAsqy/
UW1/wc1wWkG/Q9wUHTCPYAfH65qXjiyPHI26Revl4+u6hyjVynuTL5CDcMwe
cOilF1/WHMflanyhCkOq5wbLpgWxsXWH2GEWMc85oxc0/UvX1cY7u+Osbgml
dX8SKVMatphLDsoCi0zrlFfcvaSH+IoGnNrtG3Cp8+mmuuMwF1suSC33oVxr
ilWnqf1i8K/I8hDgq593KsxrknsCGTmbSzwO22qvfrC5dFmufSm/Cg9j7X7P
ag0UURSgUl1zAb9oXZaQN62Md7uadrLiqYqfg8cyHl2qULqPKhJw+KVRkQWd
b+plsfTj68JWtEFG1dqUO1KTWC+aq1lgCbl9yfbJ5tuUPr/sqV9W6IUTCWgj
mSAJ0YQMWLtOdKsLzD3RPM0T9UXOBwH1Xv2iiQTuFrl8pXX4sR33A9Y1PUg+
uOxegb/VE9P5i6phBeBT7Tuw+p2JMSBgIh/mYv8+R+/7wHI+ADA+PopIRNMr
XgVVEkNMo1E4UkhXTuhpQ2U0HBUEK8NZbPXyh8cUDU6JuQIHxKZVjFUpEjdn
CLtT76E+oNPthBMWyMqNSfdCqRS1T/XTTHNjJRSiGkka9t6iQB7vzLs/8jYE
1JvJU8nXlcsA6cyy4XU2cL/+j8R5lK9MzwJz4FCEXwm1gPj1C9VKpHO/4Vfq
RdLRQnfUDTFFqEUKSBWRnoOr+WVMbxMJwOIMQaccZfNjmHJpMSjXCROocU8H
KTvd4dh1WoPgJ7Mau8KltTQO96OYIycrAHkxnqPGEb1BAwuaw7UCeI23hVwx
CP22Yr2B05Ykm9v7CCd7S8/S1xKdpdq2hOxRIHrpjyVOtmR92yGgGnMQ2EfP
Wxehte/TLpFxDRLjbluOuQSSW/M9BewrzGCTuEQo8dhIqy9t5EklqOuoFTTX
HHxsI+7LoyUWlp124YwFsPxPH5ajPnkuPPSGE2Oo7bnpBWTTCgqCVJ5jXrAn
Vps10K6TzVPlrsXxY1CuT603S4XkiA8vP9RNqk23MSc+f6v/r3kN13R9bhVS
cCqbxeamLw1NUDrAyE+wk34igsXcRp1A8AAafHzWHXCsHc1Pk8KZOjr4PuCT
WFpfqV3Wj9wH5EgVuGqqmL+DoD4nKUA5Hs5++yRVwYOeIgI5kp9kFS8xvYzd
9y4mOlrrX02hvgf3Mb8McJq1phZzdWbDcbFALFdhpSVSziA50CVPijlRBcMk
VVo4MkYyEsF0A514hg+9QirYdJh6nGblNj9c5fwJBPOJvXWCLjFC0uHO9LE/
GN1WLIOuI9A1rwttb8USzCnU0CMhkQY1J7QSZ8o5pTVatN9JBLatnA+xUDoB
op0hjdvU6pA0HxXNIiC8srdHo5JBDuxpJnxnk/GyKHQMGZuURoujK62hpIWK
8Hp8dv27YsLI3jFO6t3dEwqJBeu6SYZc4i2tv4UPHre1gPP9a7+fRreNMGqH
dpY3ZRa2WtCout50CsX2N/8/NuM4KxPDNc6DQsYv1Q0eUfNFRVARUTWBQ69X
ppi6s0Bvj0ckmwNxrpBuQH0cKVR4S9ZXQulJqb5aIMm/DM54bLClnmEkRsKx
8wLDL3ceUram3WKcz68ERUsG+wdUag56os/henBGKNAs5WCKt929DdUc9l5K
drEGul7m+UpQl3dVEKUBpweOiV63vXiY8Q7Z4vqN7dfgp2u8K/47EBMStKh/
ay+uyO+atfsBOzCqz3gSngwyXwmIa56thC1PGIvrZ4Ix2x3dL08YQ2383xRk
XtBAn1yTddaBODwLt5tpaA/NIPvBe2gnHPw4tSNjV4c7hUjtdjGnr6XkaW7u
gS1aviDz5nAPo9A3+UE8mMMd5fhMU6i7Yk0lKMxV1/KT3G85eCPHBpDrdW0G
sJz6cV+J2HwrX8d6ul7O9JUrQtvtzS4AF4eF8pCJpd5W95RO35nnQmX0Lghz
SyDtUsGO2PlMonq0T8S7p/3/IzVDLO/6ymV0QoPti1Bmw3fEeFd449yQ1t0t
IoqIwnMXNFf/1ws2vAva77QRHjr7oApWa+tVn002vf6vUWAb4iGKgtvcTADR
88bYXDXNvSojvar7jIPJmjsOiPBTxuKJU2pS5vlX96Q6WBB3bW6lJdbTO1It
enOYYnm+rU9bFe6QDC5hQ4z1zbR+DC6Mkx8VlS+H9mtmmO2i6Fde0Y3HzrF0
5X4QPQnyaEVq4FYYef7LA94M10TGQfyobErMwvUWBfMRktbWWEkOnvJLBsGt
G8MOUb5T3ClRRgX++j2dHLnz2Q9lpTnx4V6f4MHG+hyIZ+CX2llB6cKQ98i6
8LEE53Fe/JiiICKMrGhuD3ZjIQRl0o6EcP4IVVFazgBsGJVQ4vKfh/pK9tQS
WCm/qB2zu6NnGXII7xcUCLj+Iw9t/QVnrI35NtbZzPd/47ZIy5NGfkyUPnjE
KrpfisuyK5aPO++ubucV6wssdedqPG9qQSOvk4nWUbGav9vd0oezc2Lbptvx
+8BxASrk/iXqKkIaD1xmZ4G8u20ibAfWFfy3mYAweE+/f+H6V50PnNJh5Vp4
XJcXi9IXAlUd4vfhB6c7i78mppofE5QLowD6l4/ZCeQ3UtUGqfa51djQrPPb
WCOgw9ZUiyeBbMVe4TSIyXg+osGK2G38Axd8uomKcQBIYpBMpVrCX6QMTF4F
BG4TvUFZDDd/rL1+F80Kl0k4HDwoZh/gIxEWtTEIWzQiEJd7dpD8NXwwhk0a
QCaXi8A65ze2B2pAufXgasOVT2KR+Xe6imHsthOnCc85fOdsKDTuIshfeJRj
D6pGXFFGlyzIuHIjylfG1moqv9/evP1o38K4q9+PgmjFI6uDEnJ67CcJKuIh
bPDJJugJsBm5SFEJlZ+k++M4lohT6SPgLneE3Z0Fv4o7nP7xyBDufy13Sgmq
G/GeGlWADHpurpziJLFJmHIDj5a1nr9pYAVDUwIqNtSR+CanL+5Hvhdo6/yb
I4YwvzwQW3jd9yzRf9qXLPgiyKoHM4FZDyW2q/DaJzMyaqbO0VoEWPDW2aQH
cYqg6rsjV2+dhm6NKXiOX3jX4RdYTk9P4EMUo4bpssG1rcX43JifQ+pWmJip
uBs0qWckP9Q+3he6EHV5s1BdW6vxpMYEM8qqiP6MCZPVS6D9Q09zLpPDy3ZF
Y8XgnRAjLuUXNeyxycEzjZdJoCIu0rhVjamBtRAmAukdElPYFiRsm4jxjZxN
AwA6WRvzit1aqG3HWAoDhHzv0rHGGt0HMzot/AhcmjveBteaFYxSMqvo1cyR
5Uf63nokek9uhFAgbkoUngCx9sGCHN3H3Rg6trlkp1QCMfQyUwM65V6percy
cg89UIF6Puy3yePP4LERjdJSYnA5lfG5X8Plk+oV2Btoyb7nc5gtjtUCJQGY
dd1GhG/dwFZDhMGNtKndmvMqBdfy2aumFCt0uYZjIwN5uuCT2JjDMTTHSDyh
9nO8zJBXSmZVzqIcC5IR6ss9kNTOYaHV2XTQ+3Jz0VH6TF83HHVIIbVsLhwL
8ehHL1tRu8iYiqwVNzallqAAuJ1oF45KDwrtpDYadhQrhjEE2r+en4crBUYW
IJPFZuGY22QkjNRo8vZfmpwJoajysXlPaO4GRAdwwppD2lVgXVrQBKnxKanX
PHh0s9QGAKjq8K+sKx7RDx69cOjc4VhEaYDilrZmLc82vFeughMG7lraja8G
Ptw2ybiXZ/e3z4IRuEdInTZhZIoC2QzPV6vNeHAce2gA6w2LV9DCgYZPGr9u
N8l8zz6mTn6OIl6WyETtNOSu8dCuekw/RN/nGj7s0fOYPRcf3vo3MjA7qZqt
FyXIZShqPjs3h53pfYNe2n7RjOnyKnQCXM0UwhBrmy4luFf5mPG6LO+V4gnX
K5gAV6Yez3Ocrbm+aBWBCOFyHw3UA++bXxoo+7PDtpyH58kVcDqbbRb/rYMU
LQoKPcRu5WusVkJZt8NPTi8Um57tuaNEC6/pNn5PUS1IzUsAqLQY7PvSulYa
juOKdvB1d1vzs0Y44s0oefQn8oAYsKYyk7SryjVKVhCvUA8s4gamkPQfNWjg
StXUh3aTA0To/fqJsBI5nbedPvyVusNL0M19LY9FkxLJiObxh6ZIrpGwoDjf
7XNKO7ItbRciHZu5qH8bYcvQLfLlerLVp+1YEssvpEHeoQNOkHEvw8UyTZ8y
zu0fDyOjVIynBCcbBm6pRvVqmg7xAGXjq6TdYo8FBIPEgDpS9EvtRnHhq5dy
yaAu+tLOSEBZm4XcIyPvyq/XD+9VLQZ4ZTfZ8p1gGySgfUJOVDw6kQBr6t52
ABG7cZVaMUPptKfBl+DNt2aSn45tYBg5QVR7BreSBn4pDjSN+O+x6N+AQps5
s93HpddR0o0mb2PhoZtafMQw4RK6xRNp++msNX+rrdppqQmvaZWM6V6207lv
MMpaQiK/RG1N0cybFPIVRAkSNmr61/0SLbwVeKvsm2V4A1l36/PPb3lSaQEx
o3jWsQwCqyLPLoR7xq9iNjeSjO+h2mzuWIu6rucG1tX6XQQYM5cUmtXjnIZf
uHU6IfL/3Z+PP72/JlS57Bd0FbogjbN0Bp0hmAaCRvI8WEz8ZwqSxTApFPyT
J+OlBlP22pPTnjz4oTYUe0mNEwL3z/llpcXQVsA5ULzpDWgAa9PKARpdsPzw
WqG7iS2nw24dmRI7eKkZ9TjHqQDYt+FVmOLjIc9fNo1abLdRqEJxnaTzL5xG
FmqRzPPDWVIBw/HEn288dgHfREBa19kw5rdShqD7+8NepXfOE3TfrCm1sP32
Lq4ILLKvmaSK3rqApvWhni45mpzKoExOTCKaeA4H3AEk6bZvbVQ8caE+Q+Ke
XQUX2MhLbQlNzeoI4+l/2T6QLmoc1c0DEIpaDWdN2xOYvXnXSOBMYyp527Tc
rXIQXejGbNZhx3JUp67E7flT9FHk+Ua07SKcUms0nsWDeP1NTjP+Ene2KiYd
V1nj/gl4nAZju5PpCewoAfYjL2YqGGsyOhyzeQVVEpoS8aW0NRUedSrHIp5H
Ng0SDQCCIBVWsmVrtsbVS1Trg130e/65IO3XeOtpf4gTgUwzI9E03rv9ZUpv
VZdis2HCg7kzv/TX7g6DL4sLAOblky0IaUbx0rX8wVZTZxDgjGTBEN1NPT+Z
MorYybj1JA1EwzEJBTPffTDHODfFe9bnZvk6GedlWPwuOf84EJelcGAPVKwG
/PfPxYs7VwzYL4AABB5ev2ztI1P/reV7aDMmLnDzHjkIPGOC/1A2NjQ3eZiO
kf9yA37apeB469qU1rS4yo90MK+dDK6+lzAvMlUD7DDgUXfCITVFQ1wgulqo
aMw79MryUtXZE/6Bs+xXY58VJZUZhwmdhnuY7N8lVt4ru14cZzoBGnAcb7Zq
DIevDlIDjX9cZJX8G/JdR5duF0/OsgUYhmNfj4HCI0zgtsBFCr5pac9npUbo
mBca+lgfjEpoJGySNNGFqzV94AELh4nVtjltDpFUQ8gGuJuUBjh8305NDAwJ
RB+hBj+gSKMkhJ47kIgFR8CcqQcx8T8MpEDS1BkhStlmJhJgoxnHj7QE7yKg
0Kvv8mnLCHfq4voTb0b7alJj82hLGUiCz0ZORFfnjc2dvErpwnlc7dVha6Rx
70fyf4wdbR2++1bk1fu/tMIhus6fIyJXpSi3A4sLHmNuHB75UTGiPluUrgyI
8CMMieHD+J08gDnaFGrD4CxYGzrr2Nzw6eGzBTZnDjuq/NXVtVJYP+9JPGzK
O1ZPDnIHCLkhSBmpmahOkokWgPwZI+Xjl8J2wXfYJ6vCd2aEd7lOimue2zNU
2co2kRsYEdeoTPZAOAZOtqyqHwVJk5bGgCkuyFHbJM8jaWDNiw1+WGvNMRZ0
i6zQd0eaTTP7OzkhAamHpOB0irT7lzitKa2xbaU6rkzhqfvpZPOOFy+ZeHMy
DpuAGqDDNZHZuY6bQZjuilMITbu/43P5tJjnibeLS47SzKaoe+QIfbgFjrR2
mvssC7ir+nObpT/1GI1IvzZt/WpbOEQMXIZ9mHXNqCtQyBoB4wliYZUzxzsc
Pb8D89lW+oWB95NxpcERxma/yt94ymTJLIDXwz4ONZM8eQaZdl/KIXouUgLh
QoNJL7qUg4O6lla9IpJaGMKUW/rTrtE+rmvdGjBvshxkw9oiKtyigcWu9c8N
JcjzybPqbRWNA8S78DbWAvcfaiWCo0f3cjQjVW/hXj3kHZWqu8aEQ+aIsxIr
vQCgYemDa4QlTucBmd1YzbreVZyIyWyKNE+IRdRq4tfoVFS67BwVkO125Adt
53G1NPz/kIMItX8+kNEypx3rqpdm5VaMSVogm3WJeFMBy1e4Ml7A+E2/L1xk
cU3cpqelLDHEBU0GJyMsVUXf3QiYnasLMfYdveaSXt3PZoKgl7PmhU07C9d0
1H2Eh+AA33FpqQWx6nUZmeymSrHKmlym3x1ZwOUfA/cjTVDGkq9GCGfbDIpa
IIoAuskfq33SItuxQf99SajSEfABMKWQ/OX5lUcoeUWIHJJoQUqKW0xrI2Af
m2gu08ZOs0azSlOhYWM7EpniXLnhYTSrtLLwtYcS7cz07+XIcOgTALKuZ8Ml
LmzV9ri3oyf1NK3O2BqDKOwWngCy5ChNiSbvnnBt0fA5gh74p/JKgSCCZSDn
C6zJYDRCJwwBjM51wNQbDjWUAs6TlXdEgPD3HezM0RzTKssKfSZC2MnncmmZ
OxTqZ8Cbl2eUgzelxGPaqxz1vWGh7jx+ILrG3LDFu+t4R2Lctu9BcGAEbcFZ
fqC45c43WqCX3cHFW4ZLNxA6PZ1hYUWqY7B2yBMw71a1gOq4ycvT9PqBrnKK
MjQegkQ4LXu2GVvFOo5+0qm0ZuhVQHd99vQfV3D1+OFuljhzrYX5cjfHPBi6
hn16B5Q8FPT3hG+fWctfeB6ELhvgzc4wavIPFghLiWywl4KfY2sZL6GEVOq9
3IPPxrR5kIaVuLMHfPRTRA0iWgYTVfA3U/RoeG1RSw2H//9FM8PH9P65GXvg
xM9nV55AjCt8KidARQ/YckbGhKxkDXv5EG+igCWmso+FNv+ia/ukUUdpotIU
OgyMk7thoXEsXZQsEZ/H09JMciK4x8t+07D1uArREkEBOC/GzeivdWMvarD1
Jg1Wco3EAebtpC2ecQBngpHAK+VukuYTEbJofkKkJB6st2PhTCuxEe99Gyhl
ppuoP7XsNE9DYR1yPRHDnYMzXmKqgl7CmHO4gYjPIu0DwZA25zr25eIq5N+M
G3YKEvZ9k19C+eFlcvvEp2rnyt62gRL9/emJCzxLi2S3e1ZASm+nzCzxYZGJ
k7vTjmve+B1NoO5cr6uaKlU+YIA5GLYgyHyfjOOiDo7E6IUQH0EHr1OPhnD5
8JNfsFedOtFrHUUO6t3uDjcucFIdggi8nev+8Uw5a5kM+2qB93QsrNLuid5u
313X8EhHjeMY4lp5ZI0t5juG8U41jHHqI4h6sKSX/gr88wGx5QyrO50wIoTR
NuUWu4zSohGwVDecqgER6PYuStcNp9ocy2HtAg9NJvDGAFekkwNyDz4BCAE9
AsUdjrpnLet6rmf+sO16MDkcBNlEnPt385cMNIBGyL2wg4tYG5r1R2e3MZ71
SRTf0TTZw9BwofG5DzgIe+LgAqoJRZ90IRy7p6K303RCZI7QpTQo/tOquQZc
Qe8n1hR6NTJ7FBu3iRdZJSk6zG+IuLiDeWomzjpx550AOs76TIQOaspGNN+E
X5JrlxsGm9t6SrrohfWEvr5p4GzAOJVTmZBbyXD/SdjKCeUSxtMVxQmz8cWf
PH5e/t/w1MPHhFMqHO4zEkcEY8F0EhA5ITFSp8anKAixWIQc+ybcFEBzwXfb
gk0aX1CHEZ+DvDJMDRM0V5FsA0WoHYVrFcO+lBFh9Lrvt98auvgfTqWLPuqz
/sSUNZBi85e0FQf2Jvj/ZSU34kUYolooVdUP1r3Q0+bhS/rPC2xWn8AbQkT9
6rRhKvdFz7cdh30hJaFPbn2D0CwTw/aK0Rk0wG3mxbY5ZmxzvTTVtthJ3xiA
69WPFf61NvilkOQNsXDz5+cCtDyZWH8zgX62quJ4/+vtw3bKfePcexdpYlRC
MvofNMucwyOtoARltF2R3AGpK68yy/XoDzw9TG2cPndgzWAH2Q/OW0r9ry9S
U43ubkXypTplujegVevE85ogYE/CezdgSNjAsmoZ/CjxGycqzKgxn72WGDDg
A+lO9hvA52R99Zlm1s3l5cvpfOXxQQYi1wJZEOwbgiBJdiLoEhbx2piZtut9
pHG1lLf+kJd6PdQ/1lgaKG1u40Xi28HswjkYgNDwXi4Hj+ifoh4jfehzboGh
UKK/BstibZ3UpsM7WNTtkpM55b+827hqjGLqwNYaIv2E7tZ+TGHBJzr0CItV
6od35aFc5mBHPXRWfd33g+lrjc8Gv5p3Gzmj2CKTQVxkOJLKx+whpxomKdSX
IOwoc8r0YWz3le0hgsZzPendr/4DteFu+TjUJZRsy8plA6I/AVoVKQc7jNir
i25lWgxkkmr220jFmgbSW4vM5NNOJuQSGlIda8MLtyRiO7wp61xKzhORB3Cl
EeruRMEVVRU8cWFx4PBZTW7MVJNFF6eUxPDM9jUsgNywZBeYd9+rGSuCybMT
VxI8QpOwXFx8xpLRV1sVM/ueRjEEtCwrxGPCoWK2hr1B2y2AhZhlWhfyKjwV
w+KmLbE1FABuUJkol/H0vuCht+/u4kqk4o8xxNniH/TzENKiWY38sYM9oImL
VEsBHWzVqebvALhgQ5ssN0EyQCw4TW9vy5s47nbDvr4r52MK7kNvnuknVoMI
4Zp2B0tqcUnIyiH8x5VszyPkOpRhAPb3RYgsrjPeoKai2IbDVpD94xOswj9P
DhzMcZ8H5E2cX/E6/0on5DmLKXopiLvg2zqqvnHZRGBBFWapgXLOiIhiibOH
jwB5P/+nF4zW16ay73yGRpY7gikAPyvF0pdawn9YzHApj5ha3CfA/BvRd97N
aQSBngNzwWt0mV0J6BAJiJjQYu3HY3byR4myFKt8LGi/q6HXkpU8s4wUPCDu
L5biYBtz+XzL+yBF7Elt+E9HNEDRohKrI5ZBnNXh1OuT5Jd7w0YnzojI1AfA
xhijuzohM+OiNZVbPHSM18DSC6FfkgcROz6w03aAQDraJjTlY082mhrPqeNL
FDJvX5EAgxBmEXTefXa6Bimfqfn9Hvt445iHO75aNbvm9iD6/R4ZautA7auI
/ebJQi8gXBUp1cbhQciFrMthToeYpgN3aoY7JjykPcGRzqpYurKIstBvLo4U
cuK8+gBXyblhz3LkUNSeI05AqPUQYxIwwyGhQlS+BnIGO4Vm84+/pHcPNZvp
uYAqhg5UrWq/RdBc2LKD4ls/TXaBaB7L1/uL9TRI2tRwHsFqbofwZ4KyLGuz
xS4LDw/rGUhVmWw7DTfRrMGttftnG1siPRGflNZ9D5UeMPrujcQse9RASacb
p3fBDFtlzaHAFKLFHn/Dx8LUD8R1gPwAD9G8I/oVfJSJFOEckXrVV01uKLHY
/p7yQrwyPup/UFf3VaIaXzZMBrMKl/Mdmdhg5hCEylb1mN9u6SFdcVoLEV4w
enuVQZK6qoVts1/qgmuIP21rjzUTyv2KnWBGDJyV8hRpMHGPFVYtMid0n/GD
pNU249EhBFQbTvYlsHGRdCju5ryJpI4zF8xxe13y5WQ6eSsHTrOUxFgGz2/w
GujvfG6yTXCH6E+UHUd0KPQJTYDQtH3KbB+jXxrqDag0+zV25gE34ztDy86Y
xxrBy4TL/Ikkjri+z4L8EdL1opDR3WjBBDzJ6n6JdFA+7thzijFKAhixKnvY
5jsVKM3Udte2JzCw6FJNIcysOHMqfsFRS36BWcN4Obt3RnulZ4WnEAyjoUID
HirqdIESOSrTJ3SvBGRGCalKLfpo1d0edjsogBsZDkvA7CL7fAkrYN8UJLD4
xrvogSUfnyogv8xlxok1htNgxaBYNRGSrFaOREHR9JYZYiZMRNM4HzNbP/Jx
C7Es+tjET2HmaPTbhc6K0sBVxIMhcE7gG8dor8f/nZRF3wPmxBNvrSqCLT2+
vk1/pMwAq1C3lkQvBSqggX3Bt4bSQOlDzNuVWCIzGlxecZXEgahRWMFePCBl
Yg9j4q17qZHtGH9eXp55PPJnSuUx7hzdNLSVGCIEBZptbq/YbPvpL3PJCacx
c7nOr/jvhtuVMUUpzfX12zJX8JkSRbvMjrZWr2S0iknJztEExqG0M8n4tA6G
kkkeA8g0sEkDhpa5NeFwGJqulRA72EaisvEB23n56nYSQ8h6CFawiruCUTgq
T/OCPQPeExbwVDuoDy3t+D7lX4m+CafILZqLd0rsU25rUGF10Vo6Q0fPcHuF
uT+MQiPiQpr1t437F7d1+Tz9gd8YfMaUMJfe24VwXi121wGNLceH04xkZm1Z
4TIRH5QLw3IypRB4oD0UkFGLTyivaBoDGFMV5y/mu5regQDaqYQgoCmKvL2+
Hl5VFM5ls9lMhufkgOP2cBOp38QQaeuj6HDLEvK11rbGT8gcxCtogfwa6Ocz
8jHJ9QsNZOy7IGvAXhFYW5I4Qpt+GorYMmFNKJOz/JAYLg1UkZV2RgasomSf
VNAcucA4sUzy2s3VADte+R0MDHNV6bFb8jsGxHEjzY+B2ASViEgx1qDTBYk0
aN0mou9Jl4dny+N8u5b5c0NjLKQKbdEUky2tQwtJq/qBnbRfaJwFNuPEe9Cb
wPkgwQl7kMXno7dzhk/Kx0fkHZbo9AkxOaBLjXjcK8z12y6Jh1aAeh0nNxoX
eb2/4qD82UBFKwkyaK4NAxo6otlpboIxcyR59Gc5sIwg5Jg18gcLUIjcOwo5
TGB5Z4eIYjonUm/R9UuPLtapm8bEgLjiGugQlTYHyOk22F44yFAHuHN4ufEJ
dKJobiaclb6pBWe2wm0HO00E29JVomP/+q/yc47qwHC3y82M6X2bub8NSKva
Iu7TcaGSCDZL6Gk7EB2TeuWQ++LYY+BW6uKJfvnkufSMowWZ7Ke/GI7EI8oo
C0IIGvNurFtPX+hq3HQUSMxh6EpT5CNkwocgAJ3WEYMvJkUQhvSV7DknIwog
Fx78HQU4W1pQ9rHcp5XRFL+Wr0vpXSFJQsw18MhYZpQ3VpSUQh2hG9yScTkl
le8gKpc4wbavWEP41Dl17rV3+eWi5nnVDOi7vGxjJ2ANi6/jNOCH3CtTwDM8
Thu/xtjCyfCxDk9ET4j4TCMes1/kMy/G1HM8HnIMzYLhxjXhIOb/PdrATYyV
7wmUl484Lr6ZjoXMQE31sjcQI+eYbOv6zNaVqtCywVbnbC8v2oVcZLQdHZiR
crZ2GDGDkceTCJWPw4zS4Q1KJX/TG4OjNF8ELkJxNWVguPICd4c1HNh2dC2C
md4+H32XFISoEQDBOatQlY3sFRRnt2CWciAUI3llkzJIR6poptlvGLhjMX+F
4KRtor27ibveUPk0nekyihtR7mNZ86Ig8bAYo7k4sIYXbk/XEQoMWHyOZMrW
eVo05fV4SDlotp9xvWNBGO//60S6SEn/VuePExf1YrKUzSpJXA5egPXWDtSe
tu34akA+1XlXTaf45D2X7agimbPIJhb8ah/57PyxHdyXCqysghqy0f4yoouM
dqn0uu+SUb7CrhptIHfKdbJbU4GWsIQaWc5LPfMAgCmjuNrQLGOI8hBncBug
MMuD3T6afPbnSQb8cwDCrq/egRBuKC90ZhQ7mQ7zIXp/mhPN1gojl6z0j3tc
0dLWXFWrU2mvMzyHlTor51f5HsWu9hLAN3Gl7jmoYO0CYBN+aO45pccOsF8t
Uy/NBrhYI6/ADEbrR8usYjj65sJ5h5php9mnTIFfTKSkYHKgoPgjgRxiBTj5
UvWLinBBB3YmRrljkcX1w4wKYBJcphmZ/JKKSGrxW2yEDeBcgPkEL0QLrku8
4R6blPVagpj3esB/iVjsO4lWKCr91Wr9pGVXwUfcmlgx1Bo51RS/2kgi1Knd
NnlR2kOQxAFmSFLls3g09/YyxH+TG243OTILX2dWOhbSBeueHqNphG4fAEs5
eU1aa8kIp0a9N1YqWKL/js0/hcC8Sh2Y3gBafRlbQ5JYvQmzCfY3jVeFicvS
eVzAITbpOq4GLLFG0l9i5ieSlxpekbQnsTxd7SfJjcGnJreIETA1gv7+xv9Y
uiNyTOWzjmtX4oT51F39HDQ/5x1GRdGL1hY87tHm7N1MpGbcw4VL9xsbsMJW
gpPne84HrTwJWpbe9gRqjNO+BJUk7tcgSTCWimWaQ0ggN3hsJkWtLB32/2Md
ltSvq1Qtleb7f4Fng45uDqHoPqz20uJsnMJX3SPVWFdrxUGyNpsgixdcgaXv
GAsjC9ajCEmGNoQocfZtT+a52ukJhJ1H7CADpUSUv8dLrGBcmSAPVIWQo6A3
F0XvoJpAmQirz1Bm7JWICCszqxNAZ7seHkV6vLyF1ZDoakOQlD8TYhF/OJup
h0rOXtN48cT4D67WF8eaYrKpYxt+0HFURlBQhbI09acvgoSrojcUaxPLgpDr
GJXMatneHOW38nkv3JphnzD/zGe8GYZ6bWRvQ42IG7/PLujTAMTUKu5lriYm
AgpNFzZ1ly19qwRSVYwbdU75cq4rNf6lps0rQIEZovW9hJClI+mFY44VqMLL
VwWxcaChGSplRZI6WF5/Lfd4VzX/eKT938RdmUQ1nd2z8tssPvQny359gctV
5Tzp0+q93ZCknboR3XtC+ek7lTioxbPZdVYswpVo6e3hXUCLlaRCj1xkwKgK
K2nUEoWlvjTQmdtdVHbWdx4MlYzT9Ojy7DzVV9CUWl6+3itGgw2nNowTSPS1
JtD/DrfI2xPfjnnCaiGG7/14/z8WwnbhdNgRNkOmP0sGSxNCvvjuGIQTBpn3
Mh6vGKpI/7fvtXJIgirkDGJ+yCGQ2XBEWfLLkdbEU5VxfNe93QwvIjiTHQP2
aQMeKc8sJy+J92nLR+Xjr6r8M9UZHLu5nSgpYWKnuj2XG1GTi729KxDGWtFG
NgiD1UsYS9xy7TNac9+kQFThT9QsNV9r+KCPvtISlWrlD6EGPz6j3VZnprG7
IGtAYEury2Bd9xfTeSSNmnIo1CdJkc2N7FnX0Zcc1qdDUpEwFPqlEfiZCbbk
n3cj6jT2EWwTlwBMh5k9qQXslaSn6CjSlCtDYV9uccN1bUd2mbhGQ7Hv+dua
RNs+oOZNeRscfurhRwftIaBouep9T+E2UX31trQzw+zC0D8Kx4J/XSXr2QEK
1Ac3mOKs83Rl2wU9m+GlfQ8JBR0bBfHtk5jimQIA7HdbvXs6W1SM0h7JkLdc
f63301OKRyu+Nt23WlQWair1HRdifijfPKO66FE2n+95S31TczVb8q16ksJo
agfNdx2DJD0/EqCajE67EYSCGnpl5pXOT6lhZ4m28IdRAVVy4bxxpF547SEN
nekpEx4Orm9u45zxwILyi3BtLjrE/iupy4fT7f83RtIL5hqC1lEkXIeh1DEE
JE2xS7B54zJPzHYfI35RJYArPEgzOdvyXUyxKEgo1ydQACt2muxECUn1DMee
BgddxbqlOl/diYEcudQEyTL7N6WOszKdgSmqwxK1ZO0DTSRHAAncA+RQfc+N
NPb7zL7S4FIgygAygc8QVO7uWnqmjchJFBrI+zny5ZWZDVjCQGx6I0rXvLrI
W/aP462UMHt3U3vxpDAT4o6ZQo5vbVStfPivWpT+eL8DtFZe+vwo30+NzDp8
5leLEcJ13WFxbrKfFq0s7K4jMRAUXrnY9b7pYSIm73HbLkVcH3fiGRiAgGKK
W+Wqm1AW+4seK11UudaCa1rgJm1aStDEwxkQHnAEhNCG8bBiIw4QsvYYrlgr
70YNz8ds9K6bxkxe1QD94blBVYPseJ3diOb8JjqdmDFhycFkyb5pC85dL3rL
LGsy05eTKGXhKcN5ze+Pw3+adFEur3quQHtlRekJqgdgv5c7OsnftAN2kj+1
qeAt/6gxLLP2hjEngMBye8Ie1V30BRt8473ESWpBh7mAIOQu3dxnIAQEoYr3
hbA0GYiiiDUwiOhPeesd6F2vaApNX1I1OvUyNKVPMNd3dabdMGk1jGaGx7IA
va1SmprJVOAMuQSAHpKRkLdv/K92ZV19hd2RGCBooSW4pJqLUdFcb3HCdf7C
fVL9B+YNQD/C0M7THn/b3mV9LspSEP6ulljFxLIP+Zc2LPsOLtft5VjCw6RW
Sn/5eYAZL9zxLiqb8Lx0onXq7be6en5T+Aac0H9z6Ik5oNvsxBs8RH9KwPBR
fjAjEgK0vQzfNEhUB0Mt8k39ABfDZu+XtmVYlPcDcHSZlDc+pXquXLJe41w6
wy3UCuuIB6LGsDzAzILg94Mo05TjGlRV4GMnCd/VSDTBm4LbOntedNRaU/CC
Dl2oOLZBqkJI4I5GMAUq01+MC71JF/ilTLyQ12dB+U3GmwbePXUczEeYitLU
KLMj6DK5kmeenV6w0aFLvuldOlSi5orztUkLyRUAsd790N11FnKr7hTSCPAf
lmXPOLmxtrkq6HRWPWaQeCH8ZiZUMaPKac2FhKhC2uDKluT3les1tR3l3atC
N1BrXMY66etSd9ThAIqzSXkKZ4w0O+dIV8nS7EcBRt7c4Vv4URMTzhAV9DLf
6oPDjoKs5yqYwQy4OtASpoah+/qDhqUTQ3Cvov+qZED7fx9JoIWL7vKD6lum
/wBknwYumomGozRAPYeIigob9MItXDwnEk1BWpRqU7PeavIWV90/zJGL6yph
9IBuQ2Lybkkb5xovrVl6g4HTrKheVjPg4FEgersniMexLOpdflgUeSDbBt7A
UPpadiK1jHK9VkMsBdQiaxT3MEyRajIMMTuCigYgxOCSa7ezd8sn2c3cwedD
BVhAkIi2yWNQ1VShHIzSGfstSQqw4jY6VeLKT22h9xa4vDkxvJtXN5uokDrk
grOpWsl6DDaR50VeFR2BbqV8DUQ9wwYHNv9W9K73vezUuMhCf/nLYWuqvi75
RorNsQxaz2nYeeHy+MuVStJ4U9nlQOLwe4tYsTJiYwDo/kVF369GOBD4dCcu
e+hrEI4QiRZ0EnFGH/HDnEpa7grgK6EEXSGz5W7H+B152d/OxJsgQYPFeNx/
ZcVp2eP5SZNTcETHysFQeoGI8fVZM62iwvj8WQwlQKelC6xtrNrJyh+5qWa1
/Kt5qByhbQqmR+Wwyn2COUf0nwjrNFjm2+OE3EK3qDkY3YKNzvS/Wnx0Am/Q
skNR4P0t8nAMNLygMgNSzWLsnBX13ukbyjpmFku8sdqYk5Y5b4Xo28giJQJB
4OYTsSv5sHlupPZ2bs8MsHuxpFUTiUklwmwfsBEdDnxzgdcKO22M7fyuZxtJ
XsBnsTPfOu8SWPPhf2+jf5wRQ7cdXwC4RC7RZ5bA4adcGnJtqfC0lTXarWG7
3X1k7gFJEsYDIcf8nuc9Tvz0f8AuQdamQENWKPOmFEGErKGL+2H8DjppqRyl
L1vO2zax/Vo/4zUOpZLqGvVz4Ijg7ZcwwpOPu6vHuzPHv0miBysKq29B8l2X
xT0R+K6eSMuJoLKOig0Wt8Bek7CbLlH/b9hv2SmdAXLt+ioUQi+K2bMzxNYl
8Ae1xk3mePIAr+kG2I38IBhLHvv4PjQTtxlAP4SpytZ84/yuVAF5chR0U/7n
oIYDx3Q9Uqn1ExGh1LvfO/4a3SdTxcCQGeTmB4PrFaukJvXM3mOmCpf6k8sB
cVXx67pBYNZfrsHM/oc+auChmAk9sDdAkYasVWBb3Z1ddKW7Q6GJeALb6YxN
KZwOMb7t8CRT7kVbRh/urZLU5/EPffK1VcXT1qGbOJ4qwmwkqCtoswdmnoPr
TyrO1LcJ4/I3TqpM5F9tJIFtcHjhQmU2TxSEDPoeo7xJO1bDx62/Qk1UoZGC
t1FHhFxcyVD54ahnLSBBUqgAZM4qGWB+Cl2hLev4CG3EPvUvxofeJWDhN2r5
JKYwgqoGrI4bVNQUKzG50zYoP+B5hMUAzA4AvVd127WIZp9qfX6RNaMabTwA
hJ8cm2NZQtA5s/Xq9urOQ8V+KspAamCck8Dkwly7C3nt09Wa0puw3zD2ttkj
G2RNg1/F4EoLGSiBTHnOqlzc6ewTFv5TjJR5jK7WPwvwzLdvatzwXbTDVGhK
du2cdZgKBKz61wJkjxCDfrfr2tbPhGPX6TWGejpb3zr1mimOgWnrVI4ImQrM
qwBsPfJPcfu6z4mRMP6NX+WXK5rXs69hv4WrgECMCk+Fksg5lHpqyV0yhKYx
u695qsoWVwhJ8gjrGDqTYX8mOmFQ5uI8V/DEoslzKKWpM7OwOBmXIz9CeEm/
Ytiy7ZUgKXtgbhE02EwuR9CH+DLw54vc48odqjMQZTCeyyMV/UITWi2LQ301
uB1zVbAI1Z70nn0xT2bOUmGzUuriAOYqrNVlxaAW6FE5Ntg38S6SOOqi/f8D
BxhuTVCWTxzu8gKbSOuU7BQBXu0J5Md9B5WITD1gVulgA3dTQXx3MbH0yi3c
9GYwsVNddiQp5NwBL4kStncDNlAQqhR9T2bwfsaNqkwfmS4tDJN1izSEX6jw
tivF+MZFzlnAT4vBd1zTDmKmGXkNj2yA4WMvPvd5VbKVhA569qrn3XGY05Mf
6UfobL0WmAntjXKAi82HC4iCEZFQPCTIEFQPSkjGw8PkWBOghQOISRn6UTFW
rr1yb4YbNMYCAE/Cvna8wFaeaUW1/es3hBYA3JrgM1PpzjQBIyYVCbz3AWme
u3XLZotjzpb/Pjj55xyWjnf+qB0wEW68c/dHo3aNWDDMqDuRxUvsMXWFZpa3
2jCrMe1Vm8FJq+S11TZJHUqm+wMRaJ2v0vvqGUl2ij6++hI/sQFI8XUoywY2
uUqt1YVGzhiRZATYxC4FfjyCv38/Pd3MMD8YegTd1zGSN7XHfzFk7xkBP/PN
EMu53R4nS3V0X/7FGXOgKkwlqDVAe+M/nToMOgEb4Zb9X6o6byshUIiivm/2
SExiQOtIL5JlEAGUgXZvPsToUQf4fJeE16yjsWaE+WKy7wYNGbH1kuklIdxy
sFOOe9SnWCYA+FcenbOTIyO09NTmlab6rb+L0yLxHowPdmG6mnZ3akOouyVp
uAMYURYZnDY2mbQWgl5nB8zK8BrMgNo6vJnTqMCE7kthD2TeYzceSaqP0Llw
GAR42V2tmQT52fcfZV7vrvGFx1OKlf6Ye56slxwd8E2MdYTmZkPBQv/N5QUm
+h+jYp+sz0ONTqRWAeItEm/2GgaieXnH9iuuXxw5zxzn8EcYixsAQpMyRfZO
p2kqmYeM7hfFWJCBQy49afbn/SdSqGCWkUHOhrRUKRpaIp22pIvNz0XAAmIS
sR5b33epTiCxwDD92pf+iZDe0UWcZBPgiF+nJM4k1q5363ZPEXmur2ffEIok
cqH+nbjvjG0LUlETncFD8GN5I5T5i8i+S5KDFZaZz0ACORLXPfMmeSetDQOU
7ysYXe8Gwvjyf+jCjNKfQyZhAtW7lTLgGpO5sA98V8e//hUd9QDsfr3cxzYb
RNb7dFRVzb85bJzZ6QA3uHPUMaUsmzgfXU/wF1YSh51xTCD9e4iqaFzUF9Wz
gPgJk8K613DPd68KqP+P0s1fU+ozql4QxxrrCInxbcyvMs+ZBUn71R563LfO
0KpYUCBrH5FSm+PoC8861IlHKpCpw1wVlqPhwhqr9sA2ZX1WTWwX0XmCiEsa
mSwc+5n8RW7vdvXJ40qNudDXV9PMZobVV+ScdxOPfX0kaqqpbxGbp/nv3JxM
U14r2vzyGALy33eWzOCKcFFWe12hoIUkpl9jK20CMqF+uqImUtzG7hB89/3e
S/MmlE0FjAq5F1NtLZwdOOyWkjbIgbXGkWbdwCFONmFFnTBwQDLjaW1lV6Xo
jAR30SgPxfWvr4AMffYNyhjdqmw3/CrJzYA3MAXwDW1KSCjaT7ffXF8pqcQC
SiMROKMt2kORaXDF2UTyYlL10snhW2BMjdyLUECWwk0KBo62855Q3mijs75T
DzoflJmeZL4m0fhPOWg2N1cF/FxR+mE3E4+CkQTee+VOK3rFLs2KTukakD0S
yaNDF7fIfQRdio9WudOndWExQUSHVHrOhlyYmrG310E9ilqwdEDn5H7HKOyJ
Kq3OoBXD1AJMInGdm+C9AnkTYaP1DWJ4MjXgNEyfBoAjideh3gg1mLz0/Got
D2FXN4wUW3NLZ5Xyfix4uQZOmejlT4H5/L//nzhGV1Zrtboc+Vc8MG7Fwcb1
aMKKqciPRQOzc1smtd/wo4W+ltpo8yvwuRVWDW9RQeFvx1JfRV2OoSFc4trP
gUnBo0w4NPsYyk3hEZTY6KVAf7FOkpxDSglO+H62FrHiQGx2ePOEP6Fb239E
gLx14Sr9Mb/6+zaYe233tXB1GlZ1Zq1ENaK+/zxNDaucukdK8VPC+oduQhIh
ztejn/CGUIGeHPHtLb8HZa/cXZrsEcb1oWAF7OueOFRO/O/9bYssBeYgUJwu
WO/zK2EopTLgQrRbU4Tp+bpOHZ6VpJUER5NcW1O+3konbXp78OGnPianAwDD
r5UHVcJ6m4gOemcH2eSMPx9/ayQarSwolh6+YWnjai2xF+ID18AZ5h8Irxhm
dbbEftVjbE8hAub9xdQgIk13ISH5s+1hO5oQVGxkCQOy6mhAHmKxxR7Nn9xa
hcSn8VNqP67ADeyDuxQYj+AhXmjMgPkzfoT2gyYRQMAlvW2XvHVdTerRpWiS
xksG1QpYFR5CO8exh5t+xcvPR3ZmChr1XZoxlG61nfjiiEC5JfnGRTxgw/eH
4MyUWIcOYuQcMYJjZ2eOLG/npv0Oe8f4Eai2d2x0tpQTMXXZgoTK3H/AD3yW
F+wO78+Hzm4wxYyxm4nnyOHSLCjquELgsYgH2OG4scNErpgMbrtHJgAv3uim
lfDZm5OuQx7JiwkQEfurviEz9UTlcxDJmdDNk3Xk5C5M5q4Guqpr4hUOoUO7
JSV2qF1mjstO3e/JvX3UulraNCoCewLFxlo56sNqjwgX6j0R5gVMVO6Se5/K
Aspc+wvCMMx9JsFPyUrOBYr01snuMJvBLBqKiAillrGLvV3YPnhAUTEhs4Ey
2uWCzBuOWuNhVUfr66dazD5LpnE4KSSZhLnskEQ/v0r/U/1YD9kUn6pLDrhU
SqEfkbTkVIzVLKPCdecDhXFLakEflvOTDsGQQHo2FVsBjsD/2pMvuG8WH+1L
f9i9Z1zFvrLamXPjpWxLKegCOHa+PDYOELAZ4npKOXN9LprKyTfcdaHUDYsV
eVfBMXP4js8M5tphGsbxcoWwNZ+OmSqpGeb/OnEoZVmElBlEv72YpdAX2oZa
zgnP2jpHUXVb9NyVOIPFp98ufNpBEHPrdFgx9C7Dn/pKGDd06S2xy8zO/KIy
+Qe0KIMZKqkDzOpnv7Sb0/kDZbz/sJEZCruoeIkVH18WsHo649pbQT2roI6f
P/H46X9YdHlYetgJ30AGy0opWqdapokNDS6tkgxKFtsWWLIJDFpU0sKGmdZy
Zke/UlfLFOt6ljLWQ4sBWeBucLqkIman/kOM9XNgjpOP0gVtuUmHEbz2jlyq
MXK890oMNrprq5MXtSH/FfmXsi7ZO9wHHSNicIJJhdytsiyDCAbjWMJKjKB4
QSqIQD+zmchNw4/Gx08DJSB2J5aA6PwHph+/+mDkFvJ8lEVAGT/g9g6+cnb9
ELODMVYG5+toyiFf+CmfxmsSpFTLNmITYTrQrOEX9tlIzVltAQz3rn4GxEV9
j7K2MXlKW+V3RxhkhNplKQzAWjzZYv6nmX+RdwVyVZNA27niBu3CC3B34SNR
uSTPLqyBHs3y+yGlLz7VnIsm7ApMayy3ecpZrUSQnqRn/9/U9+MhQAEGHXm/
JmlmLSh+vmZapo+G3Wpskdrpb5/fxF3woFx3jp/wGo3p3tRniyX27DUGOWY1
qBNavncg1PvPaF7Sf6INbtPBg/Vf51rvbU4X8s6qe2ZSBZa2IN9ZvVwXgvoX
YiKvTqj4WCOsO0kcNR86Fy3cKiol6jLlyKfFYNomxcamWY94tapDY0eLY8Ti
Ljq3NnrqEM1X0kneX7rPhQtBU4L94GVpdLzLiW8tb6WlHX+9UW//Dg1NfYbP
C9K05MIdkkHOlrxjPzHmbt0onP9sNPiUV/GwOLEIzphmHtu7S6jU0snub9h2
9GFnrH/E6EtSVSbSvEsnU76F/JmYGZv54z/mCkOGvBrM/dZDirjNigtHWrT1
4PQC1GWpx8hucq+Ykogaouo5arTncXQ5mswE9VHBcAO9HLl14SwSDgLyup9T
dv5O6tjlG0e8Py52OhDncluk+Grenh9Zux/spIDogwHVSHTgs7MYUSBGAZvV
aQZ8syC1bSRlINWS+76rsV66D2NOGJGdgFv3R1wdePnoQTzZ46l6tMYttLv4
mCZ/WTQG/mUMet9EAswxGCZJWFccqfq9IwA/2LvOD5bEK2DWaDQlKTATF0K0
i+Y/T/9pCcFTUUzq7azuY3Sa/5LP/yEaKgeskuXLtEH+vm6DrD1Tz+pGSPwC
HVozvkbnFMO5UCOcbitANpQqXJp1pz/eyY9rcwGr3C+hb8Ngl65pnvaxbODv
s0569usY+BwCHRbRCiYqPCWscE+SoTRO2jRdi5gOjpSdZGQ/kqStDNpYjLTJ
mQbStTy9qZTIvL5AWSCySWPrWrOcOSD1BG0d/52JkvQUbODDDoT3fqLgBkow
/n5ssjHE7jPaJ7in9TL85fO88PFTgaRXPYkrmATkvUOP2701WXTVo/29+Bm7
xGpfWLMVuoUZjji5VCi7PE5TFwqf9nIixQSmUgSrfM0hK/+Tb4PO/zoqEQQP
UkMVq00pknZWA/+F2vzlyJ7WfX8cYJvr7UGZj7hLjLajz76uxkZxnHDsxBeE
UAlGdY9SKv5t02CSREcDUM9SfB/tPldoDbjLPeZY/2KkeVHlWDnDj/KNoAlw
QUWj/YmzbU5eIHpzxPxaDNOrPeW3so4ggq/RVGLHRWniBHq2QHBxdeYNRW6x
2y3Kld9MT+51cqrFgsDObm++5RqseSk7JB3U7q9pAcPdQx/C9UzRTpZ5Ulvh
iKu3SPI9RFqKwLPTBwb26OYLEdcfP3NrIxZpbWr3mQbJR+wOgxzzQKJ/BHw1
3nbwDdbIpoBa/9OIHJ8tWpBswoFOWm6h7mmuJGqwl2O0Oge90CFMUEOHVFzX
0Iqi5G4BbHd7oBDL4WMjBNksXvtDSxOWnLiMrX94IteHDPt0A7FWY+IGu2Jt
reeG40Y7uE+171hnQPF8b4TqWTxBakWmxrrjDTjB1ryWuWoMp23o+fxdW/pO
+14SllxoJ48/Ya2QtNK2+LCq1MR/QXt+ALOa9NvXpZunoJYz/MOs/EZ4DQCc
kPkZqyTuzDAH5Cd2Zzi6SZtkmIp28SnSgsm1WSRNaZcNiiQDw1gKTcFg0NN2
6aqaPYGeH1uhV3Gu6FOQ/wrc9hGe6wPRO/KWgenQYIDtkCeLjICtYDbwYn1N
VURkRGGN7HCq1BHaxkbl2xCe6Lh3gHtDL3o0dBeh4E/SAh7psL/Q9nz2UeGQ
KPoX1EB52dvs8SfIXmRSd5/htvq/3mOIvNQqDDZ8u3XtzGO3WH8ejHmlzRty
O+V1q2GNKHos9iUNrsPCoPGZgni2/K+iBsd6LZ0ZDhPycr0ApLb/tIks7bRO
u3yy7PLzcBSG9/uCgpo8KgbgoAvFSYuOY2PSUqU6A4q/oblChRID2Om/MwBl
Avxqi7/IR0yvh0HkaGoWGXgkSm5IHjSl5iMhtXrIpwTLe6WYYJ3b6ZyOpoNY
vR+b3KhMjzSzFwcO7C8teMOsfO7IFbsyrpEBYrWbilI3RRCVXB3Lo9yBi4ge
P6Yb435g/GN2BB8s9NF7lIK+0tXAE3B7bh/h62Z7Ys7wwy51QdMcQLeohWjw
OnqKEiB0us9P7iMUi+sVv8YxBRUH9Z6eicXcKQ5UV6miwZnNj2tQ6Z6bErid
tRQb0KbibY5TvtBxSLQ2E+2OLH+sCkzk4HJFYAqto8vMUtSM0OEsZhO8NGWU
+R96b7+oQHSyLk+xdoKjmyy+UD1bozZw+ArdwUZC9y1xmIUcrMJcOurfWEAY
zN8pnkQqaM78mNQIBiN59EZvNS2PcjNes5DsrfUdw8U3R41WpCeA+Bzq7gu5
i2b95ha+nnB4KYnrNdBPhW9ZDq7dfwxAb8ducVBa/AQ8ZO6mFqA5QugrVkIT
87yis2stgI35laRlilmgcZt81Ti5jtiClA725QL/78y4DkusYzdYpZjIeNJN
h5Gv8KqQb8wboDMVvwWLspLsPKLdAjp6DyX3Veo0eTndqU5w+Wo78/SJ5iX5
+0s0ZithkMY7X8As2MSospHHHOsYS7P6kWGXiBa2ChWLpGohjUKP5aP2OWt+
7yy/fortVpkpvmMGy3hafz+/LFQNBe2i9A/LNX9WiFC29V37NKvzes8BD3rK
jP9NV7V2Z/1J3PdyEsfiX2kdeBKKOdcpjwf8gGubLSJj8sHpGAIo9R8KZnG/
xRlcYaIkkaJNiPhfzFF9Myi8Zu9Eh/BffP6tA20L6L++yVQM56NaKzeqsKaV
O2eSMY01crhzerGqyTA6WtcCiPCwLB6xC81+QrDNFBT9JgjkqNKoK1SwNbVE
+ecKqG+U38grF2kLbDN1RAVyDg296/x7mxUOKmIjA7A55GL2/C1PF1yqmzfN
7w+mCb6fWjBb8V+k+VAadtK9ZDigLcztrBTM+X3LzYlZK2f8hg2nCogzm61g
bE0nynCsuu3Cmyrt1ly8Knnu9B2cPcFKfGxNkezNTNiQjrA7x5sbdPkgbjQC
nyTGgzDPsNAkp2XnLwc9QwMEncldhiQPfNHyFZYXOE6QMUFY/GTmiw83kwYY
EI6RPiCPi1POCxh9rG6dWFiqGO/j6Vn0TUskf78QktXeA/i1f/+MaXuztcfH
YxW/DFyI92wM2O5Fyyd2G7hqTZdhiMslN0uS6geNurvTY7qnjvimrwKvGTAc
D2Niu76QWIrfgSnZKIbuWF1UeH6jvtXLb2W6kSf08B105H3EgB6pMNn61pxo
YCfSbzhbPJkNbFfgH/TXhapQpcahd8Dlt6t0SVJZc52Wsz6A3jqlZl8Q/gm6
4M8RbmcgCfVh8DTn2sHOOgOyCj9lJpoC65MBOUK65QmfMCAkewjn/H+H+Qvh
jfL+L5zFjQhr8PcnL0+OO+679ea2Z6tSx/+HJBpuOBw7lzJul8PCcEyybme9
WIJB21OWEHwBgIIppGXli3NgSVbIQB/Zwca/sL2veVnqZQ7/Q8L0mC2kPqWD
37WwJzsT+iJgjLSXNBupbIxviFW2cQpk2lh6ATWk4Ya2eqYzTla3e2DMsQrN
W8QYqYNz6YyoJqK7sFWdeEt9Xq+/Z/avYmkEOyQLGwftOEbfTtTH7vt+2kVO
WO921eV/fPUs4ar7gawE3HRVnNU22uxTlcF0BXifz0utBXAa527S2dGpL7/Z
gtqNHm2fQbwNlv+NO1vNtkEcZPkrVxeekbq4hfHbt6nZTQM+o2/azpe8SgsY
XUmbAdLOTMGVDi/pbsPaB1bvo91wWgyIO2eyco7+kOv04l1t6bksfnzRGrnG
Q2LyFVmA5meoWSMZW/cNnlTQf2dtbKczSlTOOPCnLcvIfqV6aOkFedclp1Bf
q+60KKmUA9G0vaNJgrVc6zUTFMdtfKejU1tx5iMkraF543C1ctpjVg2azDzu
k7W5Uh3n/CVYg1D31E0e7Dn3+ZCJo1Veytje0P3lTFlVUZPTD6oJt1gTt7hR
qaX1PvbMR/IYUYfyNDJ7acr5nm8UKPf9LG67v8mCxb3kgWAhW1cxJ/03ecU4
HPyeuj8lpM0VdNoUhHg62qArlO4rh7Wc7SYEq7VW9D3+7MnSLsJn66sgbSF+
R0jP0q5LqUjg/Qye5X4IX93esL2OQ3Qssza/My7JY7ziAg24uep1MW7ahjNS
lSQ4qr+CK1zOlnuWeJaPEiN7Wkj1WFPz1R0sOA7hxMmPM/r+6HN8VGq9lIeF
YfVaIZg5gvaesODQjUZz2nd3gzH77qYJqBHsdr9D8Bg7lZssPb6zoJaSPnyy
EjDjZ3uwzma7R2Roiz+KCpeVdq2/X3n7S3SmugtjYC1ba0h31lNaI6XTTMV/
g2Jh9liHEEPsnbZO4JNOyoTychSjYMsjVGuNy7ZNYqShztU5cRxlvujQrE07
oIqm+tRabA1JPFeqE62dW/PLBjwmiqkB4YhHPCO6lv86ROulV/EJtR7mXK5G
N27ygBzPJF8bieuLrc6i8+FA58K1IpXJers60teYEYmlpMZAwCpdQhAcl3Qs
Jnff24hJhhWtDlUFmnwaj09XcowvsQCD2WWgzkxKWDh+92mQhfxTMIERPYcQ
/LKR3JDiJZL3dHfNotelRzIsjQOThFt+Dlc0ucOUIAuh2xKaSMSxo7MbUvVI
84dJITdm55TtPIIWpTeNz2S2PXnqKhXiwLMHEbqjs66155tl1iichvTOHt/5
9+SJmb+214VTuIzNZs2b7vwmj/BI5xxwSEJFoyOGWhbayiR//ijuFoyDRykh
ZZT4O1fwnKWAr18zD8/oXYOdcpxEFrI/+aJef5tMT9bVcVTyRSrBFZAIgGrj
sNqNpcN6A6cglExI7m0+vo/wZItk4Z8K6pGoEU3a1nXc/Fm0S1g0wBYdn2SX
V5RUmg6Je/B02EiIfFsWj55S60XlKbaQN0CrcWd3o5cymIwqVpecYZ+0lYaS
6eAp20saFuvxL7/NUOYtKgaXOHcx9IHm+7PiYYAhfW5W9ogKVOCiDHQD9Yn3
ve8+G0Ngk2A2XyZ6nduR/jdcD4DSMKOPxB9P30cdKAq7BKmiOqWZg6ktiyYF
sWuO8Vm1TaIR1DOPEEfhQ0GnlKNlWLaXrbIsh3Zfm6dR2mBaITMnFKbSuxOT
3AgDOVwVPjTgsEqSHpC/3nUJ+ZPJMFe++t9I67S37IYFZtrm+n75nJC566nb
fvQNPPlUtFQ/yBa5swdrGgYCS9i/E3N6BlW+wLfpT7R0z5qEHBz5r3gBd2uv
+MP/GARTVx1jDSvTUTox+1srigcgXaxZtCjjAz/+L3ZUQoMUU0gVGhA7Oppy
0W1fXVoHR0wFugDLVEaxjprNSadb4z4HbXV+7xeiUzd6/UQtVZyG+oIFbjIF
Beh5Ek41udQobZbwQfynVfoFnhJAn+7udUD8Dwggy9BYfi5zvTo2u/YuwaGO
0/8Pp9tDB4v8eZiIgzzoV3mY+mrqfa/fhSui09EEO0KPKokZxUNXeUPbBDKp
c+jG5PxQ+4+221i2qnqtva85J+Ccr8FVEr9sdmtOPrAfC88PTD1l1k0gIR+x
cgJOog3PYmRg+K+74GHytHTXylQcyYL5c4hDIeCB8OmOJnK27hn4UcXiQIoF
5sCCgRW+36OTxpZSUeqtsarAMeXuDb0su3um1rDRpFUh93uNK1weMIJ2cnx2
Iv9MiaYX23opkh7kbA648aOc54HuVygYm6/fOS04FoSIuhTfedXwIeIx0adv
DXNvB8uJ8etrW3wozgUnV9qow7sd+KfQOsgoyeJZpyqybzhB/ovz2hdwvxFh
Zda2S2lQyKhoWUb7nIRXBM/pQTwpkzFaZgj82XlnFbfgLzo4hlqZSZ8UPq59
zhUcDZyT7SpH4doMwnEELIKcogGuV/rdl+MDySJOrY4ljFNBPHpYFcydLfUy
RLPDrKUc/8tJirPJZI4a5iDY+rkLT06HO8/mT2Uj45xhp7nYtp5DgYLDlasY
fvPBz+d63IaFaLlzdnzaBUkB5oA+gGWFl6QCOLKYoevhojH+SVdI1e6krhIM
x1M/KK+UvWv1abndxdqrirqXfDIbgtWR8J37kFZow7neCylRp/mhU+WMAFKP
p6hs+m5Z5dKSMuf+zjFmEkAc6B0jOiJdwUmYdk3mUsfkNfxtS62rO1I1oFj/
CrEdJFSav9UDrCwyXuRWwrKd2PfBabV1isbfM5bJ2yXwlryG+lgFmu0Pbt4V
IkPD6ErvZ1udtj9XdOTZrkEFuOdQP6Z1RX/trni6V0ZZUbJyHZSpSJHEUgsg
J7eFHoCftx7TNpdL8HdmWFK2VLJ1546UJj1d/OoWG592mzPQop9PV/f6qAYG
NLovn1/+Nxo2usVpLpCAbJsPZF3fgMGqv/S7K3VScY4eTJlHOqkOCB4jCErb
TjdBnrANuiEuHeytfbJnt4Wx1u7jUgd7lGqik2/3Dx0EpSNdmYlZUgssRonE
FibssLvawsH9SxbNOrj3llCikbOdWIYoJarb61nb3Ye1Uz7VLT1R2l71C5+c
OvNHD/89Wnd8LGI+MtjIS99/uR+L7653kvQXrFvhAMGpuVGCOwNFMhxvRhch
BW22ssS201JoXjvJlIP4I2Vsr5wKqux4dhjpb+lZkbmyllVTd7I7y+oGQ76A
GQIsMnLwNFSurxnYsbQo5+FMJNwfqa8no+A7+/hrNqybiDCp9zvdsb84PKSu
Q4ov7belgTpR5Oq58hsj3ZL2KffdH3FC5qtURDRJ0e2xDuk2Egugwrq4okxO
Pb6N0dSDRwT6MLuGTUjxvg+LzrkBDwScR04DY72fuR/+p4W6ExcbVddZjGDl
0Kwgjj4DlwVPiG78cLnaQPZfzFqk4eSZayPoDYm2jXVLz1onu5BgZd/yCKeo
PXtpbh8XRYZVtGsiPm361Mv4py+KDa2/05EWaou/B4WlFuERTHA15h2LR4TR
2BCn6w3n8okPhkmNmEQ6oPwy2NjSzXJlU8ZmnfaO2kLBwhBBnb41g6pLXUTe
2FuKn9bRzmMNNfbqTW+6RI2JlTEnFd3IJ5Pp01UJGVLdKcDV5/MzOkYrN5rn
HIhPteQ4VhQKbuRH7aqECkRdehl3S/E6QRDJI5J72WWo+9WzeLfHjlEHsklr
U+5z6MesXiVEctWwcYr7p+tuoZtSqBjfm+3A9X8vxW4B/fOBO4WxHqSf+sKs
hpVBzakEw8D2VwnJokndhV1cDWmRezWqFAJXf2dW80xZfDOzB/mzNUCXdoC4
Crlw5ml3boV/2D+gwDt/HoS6/DO7KIorGEAhaq311GivjvQrZWM0OEPEs5RF
/7EqIROF/mOrVhUNl7EcZOaNgoAfQswfkBwBBpj/kicbHy7BmOrJjd+abIie
dn8G0W2NgXBnHztBQ8oFaOt8nz764HqbGo/Y82C+otO3OZnjbDuxLUZAkiaQ
/jC3gUIK3/aQxfog/gh394P85WtAJg4XNGucKbSILT7tebPPLEDufVkKPpem
RqsHmtR9VHwidL9HMpdr8g9robQf76MoMg8eVsMYclQwO/HBQZAWIJ1z4EJy
NnEbTRezEdU4y/mgVhjJWrxzFagg5i5dK0jlCu7Vwa8ERHTUUDSSZOqw+yn8
YDUlnly5MRiaBvJSW2/L4V7lWP928lJYv6/h/u1ps7FxBMHVw3e0ciDiQeH7
uUe0uOrrwEss4JZtciWxnHLSuE2ZmEIKw8FinUhBoaRx4PnMqjM0OJprjpTq
MG4zOTRn0apsPRv+FNvqq2rmn6FTacMBO1yeCfX5w85QezVFIBiLHxftxyBx
5HNRiiyGHm1ha+1kjF1QkMyS09p7sIFoggFPShvtx18vvFNaGWMWnAbUqI6I
q0odLcTHOpz1NJF+jy+Nee9L5oYYN5ibnDPTvxxMhi5UwKYuU+uLFAS05/tt
adybU12j3CPF+qBVYKZjvRWztqr2HmWlM0Qz0Uu4iIfTK0ldYss2dZvEnQda
TG5DqlkhiUpd3jt+lat33UwjlRjlNwL2jUAY+uwyN/SRH+pTjbmY14vHecSQ
0FlW16JG0/F+nARmS3KNko5h59oIlpJtcft0qTKQodBr0rCM3TUutccWKsW+
1/WdMIdX1PZ8jwSDC25G2DXMJCwYkmiexPoWnEJFefAvpNyVYPOBhrCw1l4C
MfhUEuo925kk9bIbxrkJiQ7Aqh9QMpKkzj+lQuiKUM2HP29Bp7dhW3Vun9x0
ihvH0pLee3snUbLKNHsJ4172kuuii3IGAvPUa/EMPKBejyxDPYj5+n4G7wAE
baRbyczd6ZJweGDEWt+C4y+Bip43nPfZ+9RhFxk/KEkS8xf0gJAaKHCj06+s
e6BdcqtQDuqUIUAShzVWEVaAR6Kcu0mMb82rjf3cOonalo337mX7PLtD2dmY
kGhR0CMneIdxcEsk0aGUbNqQJgAMMxq+vhimme6jBZwmvK2qmYXsKBryHpQt
aUN+oPS0WcDcRiWLUXeIXcQ5fS6U43h88z6LbxDWoeUKzis/jXLchwqGNpGe
IQZav41jopPkus8UMwLUY1c4rbx5tthqN4B+kMQvOk04VaSH1WO2n0IUBCvb
jP1THuCZsA/3QCri+M4I5Nw5YGepujmxO68CB98GZCgIOfUcMW4OrQJRAgm5
xTMwsmgk8AASAjIYAUkCppRgHuyHPndPd0kyLitGexvEqivfrBiC09luhDJ3
lnhLYnbkiduf8HQUaLFMx/i7/2WVWHcB3H38wzTMRZeBzuV9TloHKqo4igRo
VT2uwkTHh3Xb5vnrt/DzaqxOrrWXhvcGU7GQ8qTBYa4vuZNDPPDiVqFPbRb3
3NePsN8YNWV4N9hCQxw/I6ZqWBupK2QJyXBGlGHcjw3ZAhhTwqhvk7R2U+XH
VZPVh8O4o4niFw4Lra+v9oyzGqYmPri1d03IDGQ7El3YYM2FdAdYbaYgcgqn
ofljjnm6cMPqqX9MSiQqiISdVbSYnWv1gzygm7u9/cDlles7Du/LSGFAArX2
NfK89KQuC6ce7pyYOFZczQsE42rreBBgAQeK2DJQTfD6unX7b6WW2we/q70W
7Ax8QS46ClToJ75MyTT3v+a/UhAdzzI8ayuaMyYXDdb6y7gF+GMc27uKLBbG
EFclTzdE7FhGqWo51LZVGBWeoaH/dq2FQdf54JkU/0oV1E4jVTw4D8ruvYQi
VDYQNPpv2z8YQyBvQwEjoT49PZKsA7YiPHLGi6HLR301XeBn+w5SfIQVaRal
x2I706POYy56dPNsQEP4jNjdalQs4B+vUw6WGAMtBVXf4JKwDaZ7F0YPr3yd
V6iaxro/f2LLNl8IQcq5ltfJdXxWSio31tm/Jl+ovcCO4hi48WZ99NjBnSER
9mJnZHbM2yaSHbe6Eb53xAlOOrHiTyfhDdYxYRXWmAkTM2z9S8qcXNFhpnyo
/akCd3Jf7Qm8GJ9gH1mbNDKXtLLVAr7KZbPm1SYtCnjeHIWAzZTJU66rAlK1
MBDhoY8PUxGzJDn0Tl5sVDZALiHkD9nC1DwC8eMP390VncAMggXzZq2J2mUg
bt33tmXoOp+j2K6tZhrSTApiAVN66zDmebYNkr6MsduLzKUKlFlgPY5pw4i8
mUSYv7+75WGLyVhJgRsNwQ7E1BZ+v31OpzJXYTIGjleebwlj+pBviVCpcQND
3Z2Ch1mHTsvohOozOhb7r/g5G3VVpgHMmMbkiO+TVjKf6rP3QE0IB06QFvv8
UiTp8QBVj0til8pkn64dt7xz0RcRpPDU1syKY41mq+1qq0pa/S5l6J0kRvOh
7N5KML9DVPs2KlxcLNkVp31qO4oR+98col6wBi889sTRhhm5BC/ZgKxcZT1M
ThJ8gdxQYzBMPTxWNnqVPVZNSJa+IvEvK4cyrTMdeMYANt4wCsHGBlGLZqQF
XlaYtZwwTc9AHGpnYcDHlYWu94g3fQq6VeSGtIlv4i+z2Thdpqv1ZOlBgtmJ
FQQddj0SIVj+u5hDGNHIA7nqn9gxFpV8999QcnSj7czte/NK0zIVbiK7ZIv/
LEpsrwVtBb1zgYqiDlhwdUtWnP70IgFJR8d5TR1B2fdLp9S3cOjfVS0v35w6
qKYChDdK0XQ+AeuLK3iV+njxY9RmVXdW4ICrxbxewMX6Z6jPrE+l5e3mAxq8
d3XkVPjJIP/gACOeanD/XDr0dKlt77kXoWyX5gjQTaUftWeP2LVf0MG52v2+
/ZInbNFVstU1BHHLMFRw6bJt6V3CSZyHb4AwbibhOGWpXmezivtzv1+bOvPC
xAl6ZrOyP9FvPSVdLjQbNKbSXOGutrCfYCY1ChY9KzdQGZzXCvXEJeuRSdoz
F8Z8qu4cw3OMrvWaWNl1D6R4E0H/xzeW/K09sQL4xjI20sXO7IAR+wOFqnwl
pvohwgrQ4cnWPRmGJFqr6TsKGQMosOEWykG6SsQ3UzzwHLw9mrkTcyAqIHG+
Ey0rd6DtHKo80DpwmOIArcY4MW2NWuvOgge+zpbOLns41fGFhnt+sMarV2rx
x1yfIRXlfU2Q3K7OsBy4OGSDXC4abgj9f4pN+dxLz1tgx76QjtE5cchRL92A
MWLP8FA9ZJ+ce3sxXAFtBr6lP3RnjPGBHa0FZjGRMsLZ51Xo1RZclri/Uxvn
79dKrwFUyboMsPwT+3yYXmH/WUb+bgFFarzZKSUeXe7OJzLi6fbvF27xOeBh
jDJ6Sb90JH9j/R8rDLPeLpRhphNmqBRI6JHn6lhWAbejEK12pP/E3AGE+A87
y+S91Y6cvqyDLSJgYsf4kNYphop6+Wpwea9C6Qihg45PLEcunjv8sYXsvBgV
0a2ubujIj9CiCHpzxyP+bChybyyE3ZzXDFYY2/HLLIDG60yxoVWh64KErClw
UW+u4x06Hj/uc4sNiKB72WI26NJZfna8Fij3q+Xoh3AhQdbhLU8f+0qeoX5p
2ZC+732XUkpm2ScYcyH8qpc8MKAZEhZnaNNny++dQkDt639SZ8uc5bTKiE9I
OG442+Iw6xjtEARfgxQcy0EiBJIAWdrR52ZHf7DENBmcXpAHRooppTtEgeZF
VmrdvPXHl/sHIokU11IGqfqkMtCkgku0/RO+6WW2IrVuPuVevsbM4KQcgoBJ
odzjt6l2tVyAjcYccMWdVCFcENcVcuQqZHtLTin21AvpqVCMPgAmLmdGuX6D
JMD3YeU0/E4hAr0aluaW7jf5flFJi4OK1Wok5HElwhgFkZrAVevVzjE9Raly
QNq35N3DhO2MQez/vNI87anCNwCg5BoBKLgBxNjWyODiefAuMRbZYrlw1RtW
rCxvD5YQwzBzvnSTuWgtlL/g/lGGSqGXeaMvJNBNg29p5cELckPgKRHfW8Iz
YHNzahbBLZxRGBJA2FoAM1kstY/qH9RKuM/WN7uhrGXGEZZHjW79dJsBJrGG
UOyYK7ukchTrIP2FjpBJZq9Dmk9jqpBvsnKoOn5pgaxsE1dJtxBOYMWIlK/Y
d0OvDP5gtS3v1qfgKv/uarhUKOBMc7xxXHwFh/IPfhq6yYoYH6hTUMaKizn3
VrX0uZsXjDywYzqhIWTpkcnT2D25Hbk9icY5aJ1+EUTWYoZbU2mf3NqkSMnG
A3It7+OTelrWXZJ87wGNeN/EPEhlBXwWbzA0iDj7HsWg95XzyXbTeeAKmIp+
97efENFpQExSNK8GVNZOU1cWTHb5DAvMQVvQ7tXufe1gzjAv/xvxtGLgdzPu
asbcc0ZETdzwgYd4fS/nyxka1HXGuZzfkHPdOBJKRevZD01lUXQ0Txtv36DZ
3x2ZtNu2inrHWuhQ6OLcGG6lXdc34JgLyufkNyxtX65ty/A5IqXbNIVpfP4z
lGDV6Zlk9c1odvPKzynQDLOeOtzkmeY+qKDXWwdUKYGPSW6mKCFC3ZvTx0Cs
MCRI3E49pAOqbm9N6ZG5cuNp+vApgPP/YexUucZ9Ge6XzWZgU0i26M6N1NY9
sn/dcBaUNuit/zWRusULL3eFHS7VJN03Osap+cYpLUUHLxaEKtb8M4L3sq7D
esghOkLxBwKedAkgeN8AdcSP21vDN3O0ng8Fa/byNtCi01H/2NHzKhH04BKY
0glim/pMEYy67Cm+hWQgB/XREGwTU5B6E3Iz/LGernfEh4tBy3693VYbZ6OL
nqTrHOw2iSIY4CcEsUBSe/rtdqOAp4fwC7jHd2ScL6LETJbjqjHyFgLrz107
YQXCmR6CZiwTc0xZRo/5WXPMouYk6b8mjzLhaah+gbWSOqvCjC6hUlMEhr2/
TSmAwGoxL9X6gTqtgrzuwveSPuPW+G7RqIDwdZ6ylZu6XnCibaipr/6M4pnE
1yxw6f8r1S+yK0WDcIHXbsU3kg/1hPDSf21o1zupDTxHSoTD/eIN223m8cJY
yfFYSCTrAkzPHm6EB23qWbN1b3c8ty34GoAElBEkFhvSSGHuFQp2qSHDPgsQ
BO+LyiXb0EOqYf51js248m2Nd0UGZctIhNN930VwQSvaAbmNRC+hiLvSjjiE
JEesPkFMhLTLX2Y/0ua1+9a204HyOW3vECa1TxpnQn9wwOaEy+Yw2YoaEYiY
d1wXJj/2MOo3Jv+T76wkO+ea9AdDu8JMBETbqCGZd9w8WTOR8Exv/xKIGqRG
0DInYSV0m8VXWs++ch8lTxHsF+hFfnV6b6ChtWKJ8WMmGy1oIrrGNj1iYGnz
cOmw1+8JpSMPMEKlNwuUk3R0tWK5R6ijJ8IERRYOP9/k6bX1ms+Tutv2eznH
j1PXpYmZPW/DtuXZRYsCUxgI5dNNCbcPL+r0/eObq/NRALsvlDBdnALQXAV8
07LbUHXuTpP4HK2de1e5osxtFqkE1cZrthyXtveaKl2WSfUNVHxySwMoBZ5E
5yUtO2qSflJrSum6ZCeXoDvhE2IcHhBB6RTdM8A+fkfUSS3MFJarCB7K+oJb
x4WH4GC03rTW36Rlc26Y8nI3xeFJggIgsyqA1rtCIgZRkgJhGlPd04SPGLFn
PbyD0tfGehTV7LfX2l1gFp+HvyvOWfwM1Z4TMTOu4oXpft8GtyCbQnXimIG3
3n7Fe3fOTB8GB29fWOQ9MaDUsQ/O9ir/p029Mnl+jPBpti653PmJU/wIkP47
mFAZoQV3th4HH3sVeDXWnx8ukJ5zxtNKlGvR6ap8wxOSjHXDOPQf2rUjzll0
WcSVlP1pv6IJKLctiL5wufsuz6WQJl3zlL+tueU96FfsTWD7oUTesRvmqXV9
kE4IeUvau4fvHzasVkc1M6Y6cVivUc7Za/8xHc0xtHAmaLHzt6vuo5EWIueN
8aHmTMzWciM8MiCtKa1U144osiGt0+1702XSVNDhkTkp3q/oFjnfz10fhITA
HZu+8tvtl1mEiZ062ukhOcFjoc4smohCQ9m8TJn4jDodbB0Ln5bvmPR6O9l3
PMpeGk7qA2Eu1vpiiLc5f/6OgI8IY9cK41xdnRh+8xAjkW3iODsYl2AEv6Xq
QQmxYcHhFIs/BX7EqKpX6VSyEmNPwVQ4IqfQpZ3v1yodQWSu6CmlqbMtroD/
h2lo45lk3rknFa1R4I/duwmY4OBmz+uxD3QvJZ8tp/oKUyLWidwI2stQd77u
Pa+SWufdih1/W5Qj29hTpJTgH0w9DJDV4Yss6e45RBWUpYfyakGO9aYqa+I0
jvV+0avLlNDYsoW1Vcv8aHlpr0qnZa9prkXlKLmDVRQpRoQxnJgflhoPP8Rq
BaJ5eiOJLmA8ef55uvGuuJO2hGCTEF7rVThEUyjhVUGG+vtkEBZEH2QCpgJG
4qzUmerxCMUn5lEefEMgyH2pe0YaDGMawkC6GbZUkBzq0CpwxFpdHemIgr8v
mhYPy3j36Zsz+AJr3nG+XN3wOqqZB4qBIYcHWEReM0m79BH30mvBwPGQ4Nd3
lw+3SfTeUtfZxwQFT+D6tLVTp7A70ijeyKPveSfCPEN5jgfNCUdLTJXeTe4y
UGUljgKocGS5zFKUz42rbqF/Q8iiLGo5cPGwT1wUE04Bvm7pl79GSi2GsljB
vbo23+8erX3Zcuins5+lK2Rsjftpy7kZ+gJeKqP+W4GS3zFgMkXXVbCloXRa
wtnrhci3GPG8jl9t7Mw1bNMbejU5D3+ZASxqa4J4z0dscMVf/VkYPoK5BT2d
zeeg1ii6rzWdlna8arRHDI1P/gWV3DPeRm4+j8oAoIdzkYl8hi/6+Agf62XN
AJq7/hGy8R3LoR3qkGOEkosAEjl+F2isFGpcwWHJbQdtNslnytrkaP3RoSJM
1Vn8uYB/7jqCV8uFTBnZv9/oh1YNxSzSKRRqGZ4nWw0NarGOA33HegU9S+jz
C/ehpfVmiSl8atpgY/jIbD+Rzb3b/o/w47KZQfwSXdvUl+4NcvKjHT/3UQ2r
zk3+jpdiQJu7rCZMTfr71CEExyNBCODPTo7Xs/fePa31Y7op2m5YPxubOL1L
7x0KgCGDd0wxm5QNUGjJsfmDXDv2fE05mCFB30/H2APBdab8e305UxcPiMVP
Bv26xYDbIoERfh7gRTmqoVFDoJmKM21aZ/wTvgqBRZXa67RoVunY6A4LKsx6
3xeHLMIVojJVKKqKTUlHWgeKXcJ3vKo0luMLDcYAssuCwl77lFeTyf8zOxU0
PTRq9kWImbYvoQHIbLcXqhr7hOoECi333PDbwribi0T4u68vhYMgpSc07pD1
DNVb8gu/hB2JJhIDw6iH84seKQTGb+dbSVfvCv73SbOOKoI55dtLoKnAgXi1
1LvEvM/8KYxE6sjcm+hKazrOm2CBuvkH7CVw2jvF+s0sYrmF/yH2wE1SenSO
VvHuGuH9i5wn4PuPl24BJizZWKakE2NTNirEDqVoN5wChsGURmyU6VcKTTvT
TYmU+hjVr4L9xoPIoIoUpDTZoENvcKqCa24zzBvyw9zwsvy1GlpgHb7sIIeH
ExJTX6sMXPnHjkfrMF0DaWInwYKJaL12JpNYMYfGkmuBKzilKlLbkN6S1TRT
g4g9FF2exUIBthGX6jFqIHmAzfKdXbo9pPucHFISTFwr3etOMFrRzo1JK0It
rt0Gnh1VgoW0C6dDVoxtXkq6n96/9MMZhibKZahKX25vR+3fqfL2q1uYGvaJ
2FxIwGshPClunvh3dXzBoNMsI0iEzOoM5IFzOwrXLemvss9sKn+JzPl10Oh8
6OjQh7otZ1ws8IsvUM7ChGfC8juMA5IH21AndF20+Uk5tA2B0rA32yQoZ2BH
Ih7eWwVR+P+jsOJ+jdyGtvJea60Tvu/3gPZq7ewqJv83AvRD70qYun0k71Kq
AnXOFhVcVDowkcvy9NDR3jkSlyJj7U1ei9Gwv5jwSUCydQbzSTnPmzRVkrsQ
d6XeKbgKQNF225zZxq6dBnEZWYkC7xVTqCbQRbV1ZYLbYn7wEwtehP7VmEdm
524KkXc/Dy1UKXQICdUN7XFtlp+p9v4iJwU2UVjbwOHJ4vckU7kB08zbasYa
ZtldyB7dUa+TcO9NrCcJTCBzaCVsrrAQrJThO75Z1KxLFHqUFljq7fvFoHnD
zpOvLDZn+ks4G/dbuosGD66jnMUX7303rl6igrzBi5/1igYBFHwDOvOzOZFu
bJreuhfxteHvc6COKdpNO4zuzOsTW8lln68LLS19GS7I6dIOifcF/bcBfWa4
ttTZHOfRwTjeG944DmJfY3qswsFbmDJV16S+PJgsbkxdvFlcUFQimpgbncSV
/lNIqt1ay8ULeWrD8UkgtSaQmal5uhyB0iQgLG0VDb7VjHp7wu+i/CwLXzZm
3Vbndf5WeTpUnkrQJLTNcxXMKE24M47rzZJOHqJeQR2CMTgmAu8gb3oAFsqd
XeIpdn3z7yBRmon0T7rXjdrp53d4l+2eS/zBoytUL2arCtISgCDvWDcSNucT
wSfa359PA1PYdal0rrXPag2mZm3s+foMUu9EW/mxnBrXNVHjmnJxoGaHOQJG
ZqvEpd60x+d/imq2iGSKM5mvr8JVgPQxqomG6YoElAiMVbEHUH231AQGf4dB
dDwosuDeZsjAAidb/kRwnHuBSh/NU1K8rtCRgdkyIYa4xLy+QI7N+w7ZlxoT
9eiJogi5joXcHCJbHFCtSJBiNQL3fnFb4cPKZ2Eb1yVjipWpA+jcN2IpIQ14
HAjnmh9wYdE48eBdyCppsWMCSDln22wSU5osBrqFU+Kytn901oRKzumra1oV
Rvsk5vaKlvUnEkvsuO/LL/periugJhZpJtaGQOw4Wd71VW85vz3TBy4eux1Q
ysRggU4Sz6K911jWlM96nOuFHIdpn4djCV9cUoY01JKrev01zHpStNoVZkZF
p5tLAsQmMTclMIn+Gr4YmKpY9EyHFbOfR6+a/lmOF/fnzbFZ3XE+MvuQzNq5
n6HCbhPp6zv+hE0PL5fwdEGi+QhFRUghyO/bx7wMcJMyK+AaeKOjyGnccmrS
1OVnyLji5Vb4+73TbyWMrbeCr81uKfmgsij+AQxmvEj6Z6wx2IeHsEnQvxZ+
EwQxms3+in97qkSoSSkCPuazucmvlkvDpkT2yvbIC2rmNzbfLfRS5QY6qNqA
IT/LLoZyyp7xGlSfm6QVEPVMChxvBZCpFW4GtQ+kRpF0b0jqdlY2WbFPxnzA
Xcf+vCjkz5YpDADtFvDPy4inHvcik1H5G5I5jYhVD6uNiwPJ5Bhxy1/yYg6T
FBlmyWPJl9jkl8pQ5iHA8M41a+spqa59GhHGiqdjMCrdauLcbd9SdhYDQrnK
0jDkoAcr+HkLqOu5aGgQ9UgTUdtgYwGyugGYkRW60GXLb4Fo/q6+fZrNEmhC
0+mopjZBSWCVrnStqZEjZbEh0FzyB+Qa7SvIKHoKBT6+BFOwGNtSMfoLaoTO
MWp4Of/6pE1NrKZNwHsiEl1IIn6+anKYlzjERIXbTtGujHYEHA0zIkccR2qz
VFuwUJGjbAysSBhERcD0zMb3oiNz26qzMiOI+PLiFQNu8qXDqxvGh0hiLV+j
oVZEFhqZIVFaVPrpjg+eelg/Eau0PbLYhN24YcRLKasuvumJDL1NkLti7d5/
6YmV+ziN6KsQJqXwxe405d8jY2QP77BlkyPvRCqmoLE33KwYW/UId5VIkOwh
hprFXylfJ7ynoUTIc+oMn/ILX/hwuHYRqfevVPpRXs5dZUAaqwHsxvWJNk8I
zUzGbpOs52gzw5JwfBvr/VGP6eKijhB3Y1gagmtg5FVT/xXUBwXB/PW0G+CO
WpBYhVqso8QX+MI/ykLzjHuZZEGpccSJ/H3+HCem1om1X31n+yIq7gN1Vpv+
lapXLf6YvBqo1MahKnQApLEHUKYi6LcMYP2R9Vnnr3HHiXm30npOWrRZJpqv
fsxPPFNwiuFFh9HnvMLS/gqYQVCU+MRoM/7DLdanTCJyuA0jjhCjC22J3jeW
6XMm39Qj1aWfvAzV0Q5p9LJIJbnpk+7lgdl2eHfxF7x8EOeLzrALVpWvZQ3z
0Tw6OApnjcNqIN+VvSlYxXOyPWEw1ahLyUS7aiGvi8aU5EClaHeufH8T72uX
eW3o20nx+JgaMOhde4dSWiNiWbsAqP0jDGDDbGLUP1IhA0VrT9XuhABlOCm8
ZKCe8CSln17i/nKof5/s/1So1BUATQ91U3YRx2bduH82ss9CECHCKlkAmbmq
BQ4qzUwyLRPshhhymeAZ7/uy1tzj/m+6c3nAL7io7//u3D5Y/Pr7oFPePj+a
1sgry7b/so1ibt22eySN+GvtIDJyrTEIbwM0ygR14G971wDgDe7YwRDoGIRt
8/ywHW5jpDoklXkiz6M+eqCjXbBeT4vTkfSBsSLmBSJNx5xdFVKJQvdSib6L
/B5js4tP4KuajzVZIxIr1xgmkOgcxfNL8J6HdWf9PYV0vTQI72opR9cNHBDf
TKUtjk6lW04VTvvRBQkgDPoifbO4vciec8ZYhT8fuB9+oCNyBZG5dHhEKxjN
JndyIFuMt9wZa5YT//061S5W/1YC4Kq60XpDNrqWPo1URg9J0olhs0zBhxmp
dTWudVrM6pe8XNB30lf8v7VrnhpkZCSzlCOvgpW9xZLQ+J7uzJnw1CviEgEv
xZJFgCEEiapcFDnw4awI9xBbZtbiEW90oz7JFLKm+Tpfz2ewxLnLhct1C8M+
oiGBvMnkHI+rGd2TxnIFSRr61ncZG8crJoHoDWuhVKi67p5YiC13RjEHHer4
gpPTQrINkwj6/0LSAOmJ7PnnT2LTjRrqAzW6TRUSxFOou/jZXIfBEBgQsuHn
6AMk+6QWhnZfrrCHGGMvI7Ey12lo46ZvBgqZL4D4W4KbFz4pU9iZMj+HdWMD
iB7KP+yntNxNcp+HfrEg9rcUcWj86phnWlcD2C7EJJh80FPnBLirurvR1sdQ
gcnqJff6Ns25ZomjPMwy/Eey3KdA8BHGiMTmHGMQ+lhB6Z56p8SoYH1EFzrg
zdcI7sJ8tGQU3KbGUipAHIRxI8eOd5yAGxH1B9g/oglET66BwUGFXGDZ7fFK
vkOW4mgb+/Mg+ALetugPD2yJEgErHiifacdLfdmJN5jplfpvBW3FUB1ihKJH
wuwL1r5trfzXZJPwjHOTsDNROW7tEB9Uccc+5KHgHSQCebAvthn6YtdLU3B8
zp8baWpIwM65imLFY7dw7tPCLDF4mdMfAAxjeSh7jEZQDB5Eq48wbDS3o7ap
odl2C7nxzDvFw/00CnLIV71x6YYMOQoogvVTlfEmg4JPZQpZbcDpkrocoxpP
V3zO/88mPiKc/MLWYm88fRRRTsIlmN3Rkdw+AibZC/3wVTDA8FgLCvg1qo+E
eUHW6uMeZFCUPFavy4sdgulIIvd4q7b5zbb3TVsoDxeQAhWpL+gkFJgC0fQc
+bnrWmf51RcJGEM6WJIqcUryutmWTDN74cs1bG+nni7PPLfXVnEoKZF3sb6s
tCHgcAa+sLPLEK2dTFAqUQu5MZBD15qOWdmEo4wjV2ljV/69PqhVgjNJ+3WC
xuqFPsHfinCj9Yy6SIYVUd7ekQb7cVQ6rcXo/Ysu5dTPAKNFb06LS2HZXxgj
fLadADgwyt/+SNDH6YRzsKYOG0v7betEpwB59LahGS5g7RL9Gtpori+f7r8A
g3GWxAmWtKnZWaKqx16a2Dc2w01Jgxt6xQk157MfNtaZJWO02jWbjGJ7A79f
8OClG7mSCzU/NkLP6lVxa11YA+/rE+tzcdnsYYtYPro6BLIsZBQqvlb7K5wD
h3OZx3U36ES4LgIn/0z9ktGdw/9flgj+187JXQtxF3GoKZlgIaOtEsRXThRv
hw0d9UBBg9rJ8tQZUV+LE8BMXh1o/EDGqXazD4kxqL38Z2cC/DxwBPZcV0yo
7v38jP2HNsaHcJhM2hIlYav6PThrh5S8U004ZXxDcoo/9veknuKqGoMzPDWy
9SqRDkFrEVXJ9sZR7tiBU/aLNFbjuI/ZU8ci4r1Laf7tfzbLcwaUo15CwU7r
XItkATu6IofbbR8sBZjPLJJZFm31xibiluF9KnznLsdho7w1WD9xdgyqBHRD
2rnId2LZvVbTddNn373+JDoAxO9+CASI0E48+umX/5VucxOmRdmhaT912DNx
+56pjAUd2tC15zozBWfDGOlW+Lph9K+A6z7k0TDKV8p9ShOdhgi3XgV2nAhz
1qfuDz8GyGRHuqE9o4Um+Pcsy/wfBY6vEw4CeJwMu+1Vb+5kMM/XWKiAlwFq
KILvseF3dBG+fZPbGZqJQ4dDsC41dZ3Qym/2xs4nekh5yVjU5Nd+DhqqfSoX
kadV4tAW9Zt7o3/OvXEASOdfHQzGISLm8t7YUzdOZeGco0Pk4afG7cs/VYUK
zJoSOLtTR559CTljY5pi+IT8wT/mPXGV1rtkXGAjEV87MH7oxeZJv3+fjxYk
U74shetBbFIMKl3FIFlLSguFcA3xz5BvU8zL5X0G/8dIOz33nz9sCAx8UY4s
k4bTMZkti0SiezELaBhx9JywZXn82sJwi49bcqTztO/fFglg9wK1RXu5UOth
va9ZnKHq3xXTmknBEyp6dotHYMidLmq6rK7X/woRoQXTKOQMNXH0ClWa6ETz
2GGuzCDuiv7KbTxl8RBGrL2I0BNkhE2G5RaYKg4eW5Tk4GOMxsD/eq5UHP7I
Dtcq63EDvuhCV3pKZp5q6VXgT1rfX72qsIRxKsUcC7zSv/wvcWTebF6inPFU
e3OGr6VPdfnkF00v5r/ImobOiarc5fKEiFbCkMwr2IGYd1HZvgsxTr9csK+k
W9rPVusEUJ6BC7R5Z5VUxdWEssbS8pdr3YydcTFU4AGR8ZYMe24GVcWLYf+0
Te9FnuNh0c5BvQPA1D4vDZAATzsWRJqw6HVbFXzQ0BegTRrxP8z7T4/Bbhlu
au28ZhjeqviS1xu0Z7azVnKoKVjdHiCADP+nT4LfrRpd2dBJNjKx6+uSo4+W
umyZYZcgD8yik5oceE/Bm/7C+UNAA+p++GAtFpGpz03COv622pYSJew99oGf
2xfSmqUYF+UVyo+63GqN6RxO9QIAg8JyMW7TOhPfIagaB2WcsuFhF/hG3u6H
qynciyih+6cHKhxvIVVAa2KidZn8PHad3EmuwjkeXRyXfN9ncKoxXOALh+j7
3LeOOLGxKRwwgBXVICddmX8pe5357QjoqDExiO8iouIZzMs653+SfFNjI3SR
h7Uh22/Wr4mjEm6gZV8QX8RdQG6Ale6zWZX0Vcj4WKPzMGtCoSB8RteSxyVK
WIc6NEUebP673/BrtxHTx/K1T3W7IpZVr2LzSmlO8HFYkY/3yddXMRoMtBLd
TtOkVfB/uB69z7+p5BSRf+s1xaTmNL4vY6kWfkhVv2UDX9G6D+E+dtBb74Jy
NO+YoXj3kDZouUAsu/pCqWaPwtuqrF2Sn+8f+i26dA9nnGkSrcReyhvwznEw
qeAeCDnUxocCfnxWDxUmF0FwIPzeBoXCcqcb8tuRVpFCc/4ywGsvyuIlpHRU
iekLTUFvRmwpncqde/NT6LZ4vznIcJQU/GRPFd/+D+bt8bC6eifrW4i3EoGp
m+AbLJ2Y2fFhiNmIAPcUv4wkxqSKgD101iRpYB2MJ7visBMP9T7rPVO2qWm/
ZYCVLUcvNTwjzQM5C4teoIrOhWPq4kOfKN6W/v50vQXCwThKJBbkjFbrP0Tc
KYBKRfeD0339RqHvvOanx4D94IyHvwdgi5gm3Ctszt79ql380hGCJ0WDl15/
Og3Q9CqaH1zNNRShgL//iwzz3flQCI9NVCngXLhFUXaFBaWQb6qpAcEwrog9
hT+nrcolmjLqgDg3MW7zwohHmP6ly7iDL4+ygjBodFWdAtMUNu2/Ys5bXk4H
vrrAAF9z1tO14MoIJ/G1VwLwAHZKt4Sog7EiIcZ3cH9Nj+jezqkDHpsptE/4
/BVk5MbJBLUnN0Oy/8L83HObRW0mMiw/fLMZ6qA0AzeuWPIDtFjM9Iw2on45
19begApqeW47AoPqO2HT+iW8nmMC9BW2ZDM1vrINF0r3BzlJHAncauJEHXbx
v0cx4yUkBAjHU8E4IO1cfvya2SbdPxj3o/k/kmy4tY0W50yh5g5ETnWw7Kk/
jxDhs6MJ7E45H8oZW6g4RDynTzMB3csnRVEmrjc8VrLHxMsqio2kohkEMIBj
smzx8FmKgowxjDmRABzudLAYXW8bhfHDJu7VodTjdkWin9Kpazgf7ID7wr9S
Z3cdB2L8NP7xnGMyEk4ywlmlJjQaSUJoz8YDoZId+rCVAerlsz+ZarIHwUAT
lvAwlSMT7cRzWlQl0JiK5QN9ao+IB02A0MMyN4PDTO1Db3+9BWSI4QCpGLEg
c+Kcqx0aYr8cem1PXS0SkGSCl+XzXRQWPgnq52hxRSqu9hlKFXCtcDfV1xlV
NzH7jIFUWUGejBWpfisQFR/vcAtCfOKh/Ze88aoCZRyVGPvHPWgUrD2t1ufY
PXHaURsuxJIuBerMxCwwy42q8eBHu91/f4kiM/nVvWYuOxc/otbTnejw/SyO
9HFrEG2kjnqgzykknW0WhfBeEWHiehQ9Q8fkBOU3kMn9DmegA3hz1++cPejS
KJ3/ryYWrlq4TZhw6fAMgBHh1+GODyEdiCVrPKqCF989gDhPnkOC5R1eZHAS
zd5IZYyrkMpgWiTUL7CBJSun/eYndO+DMJyq+2HvfNxgVpXSeYEhQwo+ylUn
CbTLBrtwR8CLx7jIfxkuq7zxBu7k/YPnDZQ3oa1cf2qsZunsUMhBCtT5rk3W
IfSWYv22A4XIO+lxQVU8iqCsurVrwPN4VHohhLBb13hBVcoDccFYhIeFsLOC
Z6BInKnhpT+FZLkGd/QTriebzeiclN4hzdIURdwrAlc92dzVAFIexJsSideB
M110tIQuj1ub/ws57QsTooqZn20DhQ/fueXArfTMFYCTUgT9h56isbB8qlvF
427clLmJwMTPS95SGBsLx1QM9x+qOHwTTAA7FejRcS5OtKCeRX7ZNpJjuaM6
nVIovTrsIq/3h8ZBDTIAih+M/1ghs5amVxSGRb67cGXQFJKoHJ3oolJeTenH
QOPQi4KxlpnzVC1acRfNGMsAjt/kFvIgn4RsPnFgC4qlMR+k1krxiKyTlqUL
NvsW3+OFgOUuBHrgKczUcuqugE+cpG0oyJLbQf9njWtM4QPNaA0e56xvyFIr
SsOrF3o1Jz3jJ3GQsXwzR+YEComvjcQ6GxvXznZ7kRlC4Ujghxbz09/WIasF
CLiOZjDhZKiqkMro9xITjYmF9mQ0Yp+qNvao3/JsKsdd5l1Rfe1IlS4oUaA+
uuS73TX9vqiqiUI3PN/D7umqKjVUp2FzgvT5SYxc+CObLgEoFhxX93v9xmRg
07SoGy5jKPnacftxEHAis66BZAqzPjyI+Nuy7ik0Pq6Gpd1HH4rDwfoc5fwR
MmyI/3/NzSppKS0x9wB3Ui9lt0v38TvjWcimNvBvkiMZbo49UPMMAeaZaT1V
EjIV8dOfEn9vawn9Ptk7WP68MR5PF0e8IxJm0l0PB312nzXLQGUQ2QlLqFJS
0lLifDElYgS4E2bsN/09lIToG0tcSyQXT7h5XzPYcd6+HQbmadtEl9OStI3B
orQj4n3DBKeG1G2TUJZjLQbYXeW58rAp+otPn+x2zKgpMSBIfog7EpYDNdlc
Vk9i1BDjlXUzueUVNLR2L9CVLPTgiuIstp4HXkkw2vkJ/o/o8YyFaMmT7dGc
hWabZasJPF2krvF5FVPabDP8oUhWu776UqMwuuPOxLJUKnXH8M+mXnwZDsrA
dDDXwoJMHgzbgE234JYgvSALooDCwv+nbpnIIioi3IceUNaIDXhfALGnRn0J
RYT4GsnkU+BQp9uMneLRXE5PTTgd0RvbK0vKwVzGnxtxPcAXq17LYwBP5I7J
E4KopHYZ0RkhpX+6YJoqO+qhwEEvHnhdZBWnIuO4N/xAqccrHD+tyl9HabVN
F8EYlJ7GWAa0hHQahpyyCSTju3wy333kyLEoB8b8fN0Y06XEfjwsFsh9Ek72
OtX51X7c4wo6w1iXWDehxqYF1COkpfH2ggEU232OseZ0V8XSbw6WjROwy9lm
t7shzwikqAyESxkiYOY+Zxgb/rqIt2zXaskNzdken3hG455f1OR4BjmyvtJq
fovvSN+DTGlkuIiFvFLBHKrD5Cfe4WXGbWmOwsjeKgaGrSp/D0R0/enxJ66o
s0wenuMUqa76OUld0ozCYBgha0RKuEyY/2pNkyKGui+kAnIVagNuppomUBj7
gtRw/Aoo7xkryUuoitzmZTej24If6kCrpcmOLZR0cpyLt++wJR2HQhJNvWUj
RN5Gf4Ao9ncTX5oIorVEfytlCYE+nJ9SYAD64pmOmfvyTx6wvY9RUPNvJcY3
YBMP/37K/YtAS3ljgODubCEMojqthXOXXZcXdeJX4ex5uo/N+Lj+aG2p4c/Q
R2yKJ4wte5VREIsij59nLBHC29bD6nfZcf+vhvXJNA3lqZ2cY3tTlReH2ijC
88Yl7RjjIbegfEMS8KbrPM8ZBHldcopISUNb998EtKL690LcF4wu3kICRXkb
1QEpQtvqG+w3fuHDxz1P/0oJakWZe/QZcT/UM5fiq0l6R+F3FUIEpgaxsha8
ftUi6gsAQLmYxSNXOVABmA8eJ4SOKtF/g873vTPw07r/nAiq33rwa0/uu60Z
DzIceTnPW7CI8s/ech1IQJzSMxefedfLfctbyWRibV7N9YwI/ftygljGevnf
8kgRinBLwvE9GsSm1Lf+wz12B1iGtfDiovU8PZhQGgH5EKU3b/nm+IoODziA
ht1GyvoQOHLUS+s+l3jVO95Fjt4qwNjrOT8K2YqOiSARsGGku9lzLIqW4CCS
a9iU6OnU5SfK8aJU+ltq05+KRyGaThjDiK36lDAKzSnEgcR4ZVaLMZieBp2b
uCaylK+67JMvPb16+cbM6AqiuUUN0FZtwQ/TJSm92k0iwYT6q1qFgK7TJXuv
ZKa8seatstQOj2CUBbkKSN7dZRmDMGc6gX36eq0y88DDJS7JcffzzPyROH63
ve8LKJwlqqt9jKvIwFnVZHFvD2QUz7n5d1GEYOH/8VFRJ8R9G12ExAxBoQZG
rO5E9bKXB8JJ9kRMZdCwnWOYrnq8njVrt/V/dhoyVQ8CG2TivkquLR7WLRms
rK06MGA2hk3BjFGQ7Sq7acRLrIfnQn1zG25fZD7bJagMvhJR/c7ocXBeap5B
RZ//cMjsucjQRQr4rjxtBP1xJEIlbe5gK+o0e/nBG+3sbjdu/JTCDRVHo3Do
dRjwGMboNqGsVU5O7LO6ONtEJXUInXQ6SNufMhEv8ZLzOwtMfr7yRqDTk8cP
lzJIDRwHl0WMHX6K3jXlSsa4dKImTJniODT1AjmiheH0G2yKsE3vcaPqNLfr
4vhj3AEuQRSrAIUuPMYtm8WXmAZUJxQGeY13pC/u2V05xqvCI47kc6cxwR8c
UXmqBfdkaayMlB5HdGj2H59866XaNIWiDDPlTQbRElsm25ge6A7ka2uz5Kif
uf+Wem/uQw86+otYHlBDmh5/QtihxyKcX4js1EwsvrYduKglfnwXo2qHDwbJ
GaLNN6NGjQDbVutO+k2IMKnkjBLR/Ihr9kAtqW9gc2UzOFasqzM8kbCkvAWQ
l/VmI8qhiBa4uJycHCvbjLcGo4LPSYFzCbygjcw0DxYxBHCXHp1qFZZYntNk
AkEA0fLrg+Vj6R+R6scUZoeoOULKJhvqWKBseVHNKgqMqY9J1HZ19ij64Ive
rfN8uZgdZcsOy8UDcgXWfIxHbXHAv8UMCHqHvuM+eM84EsBszDJMAaYgc/9j
XR4V5B0OU/2VwqvgrRrsBr6Fn5mR342swJ1/mnnFV5XjunhBlIDfwOeuGid9
hoYOsP2qMyGzYs6QR7ZmkRnxfsQniYFHMMQFw3pZy/G8EIciDoL338clU7mL
bSWpiXGoDmLCteoaoEL0SZiKRRaOdIYEONWDTk9xQ36LBBeoUSP9LxBQZ/+E
uWKHBeEPKT1M+AEqDPxUxsFoA91zCkasqBQ06JkO9rKpVmnYHQc5SsKnDZ2j
K5gS1d4w+Vq9bZfhfGTsR1QDvnr7p0rUogOdgQ0n0ZA4Y43+MMKLn9vHoPOy
UKRccssvjoRYlUXTEb4YaxsLz//jikBve9/Q5sgHdSpnn0u5IKp/GXtzIP9A
cXGcoBwAE0lqOrYvV+ZM5Il2q9ypukgSY8ZFVNqX4DVfxBYVJtjBynltjvCD
P5QF2DjjMwuvBjTbUaCnrv4AS4LB+dDQXlLW4G+hCw7IRo1HTPET9RLS86Pz
ihSNpmqEbqqPdcYC4uUx36ro0aGlC/ANqYrzTo7KWyR9ZG0jIQ8y9Dn1reNa
XNN5OFcsqqcNkXlDgKz6RR78nkO1bjwphn8H4TJVboN2UwN92TXAh3lnTJZr
wgQpRaB/tteZjRNyicZxQK6ECislYlSdnzvgbXnDk/g2tEnD0C/TmhpHDoRf
OuWbTKnLVYiRHVkKXpvKcBpQwGeCH62xbQpurIQK6WlFYfoIIAbTeQGN7zJE
DoVTCa7PH8W/Kg3UCZFFSveIDmtQLV+KYOe0X9jSjdmGORotyJ93pYHNcOLi
hH++H2LEwcJGPRIi7JI74a1ln6jwcs/DgdwEiCdaDbOw0y/d8YfL+YJbR4ES
QK/gucy88X6BFjQ9j4uZZp6uLkeJ3k6KcR8c235bke83h2RqM8Oujx97Qi8z
rDrkLJ8oBpweKe/f3B1xHybhH7fZ9zo/MfqZNyNTHqCw+uAXd+ufTz2wFifc
zhazlxx9vYF0B6lbvJNsru3cnFaMDlmJSc9shzxnafE7VOUH1PZBimSrsLC/
ntRkUKEgdhy8cUikSUXJ8kclQFHSfEoemEQmh3p9QEDGSitzccJeoQDyKZ6s
ZIkETn3Ha2j3nOgyipMsjYvdtFMaUCWKOY4ycwKFLl20U9+0w+3EfEnAWNAc
WKzjcbarcHm5Y0tpl2JkJmORVjlEgxHcttZEAlHffgZpNFSnvBvSFO3ol4zc
q/q8PXMwcIl6Nx6wkKAHijU0VNFEbnxJi2APsdfqJEDz6S9IUjv0hwmrrQgJ
f5Pb+IP3OqL4+OH8+cekZt2JUkcJF/iShN5x1np6m90IyOtQdRN/vNvM4Qwh
IhVuteCH+FIGYIPIXhcN86vRb7+fjvvoJ2GiY/T/L/VY5CDRYVo8JRSs50t7
iXjSJQsW1hMz17t5iXT9kxnj42wiRJOJAFsLT6oBMU5phBZS23Xuhe50Xuma
lzlGg7MrqUuG19YExvDkMrI1IDx8f3BVvMf1UdkaAPxFYNNsM3zL7h9Ltxtu
7Yew0k9nHVgdxcCvCmlwAJPEKdZ+R4EX/OMEgCDHKndPTN+nQY/LsPPRq3we
nZ3ghgBjtaMVvulnpkcC+cQxqxVnO39pf1pFtIemvUKHUghz4hrjRWT/E20E
mHdj1ZAM/ReiVJmAVlQAmqy/9oZeRXQuaXlC0ePLQEdqTcckJq4oDDkyeJRc
8RQ6CsWf5moKUKGwFj1l4X8lNlHvhV5B/UBuIu+JSCX69+rhhZxKGTw+wwtg
5xJHY1VJNoImOAJf39jqjUCvBScsK3DBQyfjplZbOBH/SAb+EcqdG4K1rbpV
UpmQDPspFL/UZWUalf8OvmsQz1HUuLD5yDqg9eSSANkXfUtWvDN6QWZAUJUk
fl38QFbZSkSIcagvYI28o0SC1SuO8ilbTiGjkJ+UR9Qjgzqw8uLcBc6fu0Ji
qCrFaO9KW0p4vMBlvKjuK6GkbowhRh4frzqWa9D2CDOoyDtwH8qIPOHpp4uf
41p3RcAqF5J025ZO1XJn15rCkjU0ZVHbQJ10Bc8c84wVjYQLN2i8q/UGIolJ
Owt4tEzsKpylUcajaFzEoKMuLwTSyB0pFl/05+bUdBai9TvClCM8ssl/yT1E
mkcckKg8D2W5hDyNKjFkU7Zk9MJ9FGQ3OPsWmZu6VU8iTjZZa3iKEMxnL9Fm
LBCn8qa8eeMV7wpgXD6xaR0DUMaslHIcF+k5gBJ8PqvgLOP5I4bqaY4i20Zl
6OeCFuG0g27IKLzd6/bBe2gFUzmTnon4nuFnHFPyCrgblBStZDTXqIyisRv9
D12xesL1UFLvzxUXbqg3uZB/TFkchGhALfzy3/2DCaahByC3Rw2DQk5C5wo6
AAOwWO/5nWINKC3rmcPEEfdCZaI8D2mDEkvHjUJ7RjW/dSvZ1I6mYR/YSBI4
Z6zb6CcSVNohWF/0Za1V7Gp6ES6pOEB6VSLRPRCVM/GmDiZWyaRgdRrjPjY3
hcQR7SrxREYgwusnR+zFEEuudMDPZqdC69VvC/VqBTc1riW4pCVT0EeAbAba
7hKuW0MvGFVtCB6yGI6HR06nEP1+x5rmLSqTo7kywgUVwg+J0lP3AMIGl3hQ
C0djHxRzuCMnWaDGdrr8kKVIR7EYlh74r1kAW4EsoPJePi6qWxEwJ43wHPJ9
cQw5clmhCFn2pe7+7z7a3G2THTVvS2aGbI9D1KHDCRS891HAeRYgxNM8VIG2
k71V2tar84K/s8zdN0OWDrkpuMFAU4gAmknIaCd3sz9gejK53zjr8plMBlx8
sa+LjmhqAXoZ/x0CgNYUOkiDbhiVuF4RLKc+x7ALse6qTS0+dsKGx2P8TnTJ
E0TyadSk/Riynif3vxGVh8sdhkUAyb3bm1vHLe2wDKTuSOWLvIOKCZcPcxeJ
MmEjPpJZWjIFvLGN2GS6WmFVs+YQvHLUq0AJ5Z9P6CViHA4fcg+B9YUERWXe
S6Ck6zdfIUqRbtHsjmC+xlAjGFFIhV06PwLrFjiev1DRCwjSdUP3cVaKfZm8
ZLne+6kFfvef2xORUjTQ2754O6SU73lGtUHGHaO+1j4hEV6qQZ0F0BBos/gi
4pfkROamN2WVIxrcgGy4jInfFdwYlKU2jOaK1c8In05N63RBNYvarxP9VaRu
PV+6elbhwf05PYcsv79fgSahh7mDrMTWULs5Cb/pSCKgVSAorkazEU2QZJYq
EVoAPVoPx17nf5gF3zg8dXT2Dy2DmJ4inMDfqI0vI9WKWpmtzCtCztOdC+/9
T3Xn+pR0Ze6QJciECtDk+tr4SDRgaj1FjINdHZrmJ5XRreubMm46pPKUrZ3Y
XRyQmfJhYVZ7mdidVoqPelXTm9U1lVtVRWA8FjeMbVc7EW/Td94LfJUOU5O/
IVxND/aR5sASeUhxQAw+orNE2Et4kwOFPZTyY7Uwt6cdEpzJ4CFFFMjT8BOk
0GLL3HIj1TT/4+aA/bfofsCubp6jPYN8H7VmbfnPg6i3sLEgMa1JRbNvZZcf
RvryKbaWp9AMaxCsiy98GZHG7Mbw8U6AfO9IHX9rsC8EZckaVvIUspWc1o6d
kx5TSjNIMMOnnuDaRKz3yfBgPNaQJ5xJCK48pFO6unHcggkXXCZTxMzFEcY1
J/LjTjxLTL/iXJpZmMgw1fD175lX0t8ZVOdKxXuY67L2pJb4FFszmU2WoDHh
OOnXumFc2y6SFZjtfu3xbg1GnmqYps2CL2WucEI9gl4lJRGGgNnPg1TTSHxM
wQKKAVZmu1k+EVAbbN4v5Ssl47CAi3lVgUJaHADusJFY1AwcnRB3xijKV/r5
L3NR3aZUSW3tvmnFdCTIN1lzwmpHjKbur26lKJUpgLexvyW9aRv1RXTICC11
ohX6NUeQ2yQzJX8X5w2NZBb5tdj/TrnRYVr7QCZmWtlRM4v3qXDXGtktQ1tn
RwCsfZgZT6AWMcjwP6rC5+vjOwrFdB9VdU3yWj4Bh4s6HT2TyIGwvTwR7Wx9
kW30yV8kyb9dfWsJmIbksg1vUXN9y9XH17vanoK7+C0PuD81zqo4fWJmDiI6
6FoUF3o0Nx8b6o4o8m0YJJN2gwhYurEEw2eg6/FTyFUONxGSe8yEufr6joB7
tkAIUbJaVcFjUbtZOJRwghgMZReTSuWQ7gZlRvOX2AsdZo+AR/kwU9F/yuZZ
2IZBY3qXo2xfSWAhhVTPvEtuMOHJgf8FvFD+Sbr0DnABgaiuwStyJ4bXP2AR
LXJOjOSblh4Hpmi9tFNecvlJ/oeL0prMd3s+3oIjfdyqYH+rkj4HIjB9Wfa0
Pne/YyffdhDimp9Ge5w2sSiI6LRxKnBFIffJaSfI7vLwNpobSTjVixM7ShKR
eJ8K49vnYIW+KI4HLR3v732ohuFxr2l8fFJ3UrYdiFXcnihLX5utmeYJLCvx
2kJ/iLRdBBPCk03TNfyZ858xld2ma+kVTDjucaozdmTvn1dQDMewo1tOaiRi
VoUnfuweXBJ8aK0iYhDDvwTA8KtL1ipWTrGjhQzNxl+e8Sr13rtVhb1NEmDH
A5z4u7M4vsGIutHymIPFoYyG0IoRIjAvkX04T3Q2SISRPuUvz0dLSjivuF/i
NmKoFoCfRJkmtwhkY1S+GOd/gc6mEFGFqvuhg5y4QQy45GOfquh2C8tje2MD
sp/IxVYF3gVr/sx01QAkUVihox+ti7FLYEQUcfPGoZO0ZD9h4I86ASLD7a/H
eDWYdR93kPn98n/0MxnQe1WtW8El6xWCULYD9Avhu642knjBGWV0lNlcqGn7
msJ0ci24L0O3PaZ+vV6bZFCSQF9VIYx+8ydD5uqhTA/i206ayq0DsSyUxp4i
iKmapenVdyyFwGT716/o0YjAAYRLc5s9Xe8xbGSPVPKVFBuVLOPg5hU5vku9
ytooUK79bRub53wpxKWJuYArgwfGRFxZmsuvQn0z7d7YITFmwyiWGqqHReKm
AnYgaOV4hXEUjTtEEVpMjrCBKEqmjfLBQYj6NtTbwjTfkTPrR3g4so8vPmDu
BhK7yp7Zci6Qhzi/EkiCh1RdUwui18qamNO1mTd4ox2VcXQ/xpBd6Tv9D3d2
ZFr+AQlfnDIc79WtG5Mqdd3g4Iq8Ox++wwlwhJYSSOqXZbJBT8bgqqnzGZRW
gSCofPdoyv6LWF/yVKOFCpmQ3l5MJcPS2x3OjpuELSwDq9PC19thA5E8kdWQ
J2xb7j3WvNnP/LkLDy0XSxPzBjOXrSpNZ1YCKw7jgLElH1tBk1svF/3vEuYe
rtK0K3ZovPuYv0lKy3DYHcXjW4ePIswNdTdEfhrkBv/p1YUyHUm49fk6xvAS
rrSB0JKI3EoKlgkvVOxFrhcZb7CPdPPvgOLWI43Xjo1jaiiG6ZHeDXI5Ofao
QL92NcKx8xHzqfu44lMViOyKOc++GmEwt6hzznTXa24m/LXskjivqDB/sBjd
MAMpTdnOBirRt3ij48E1BrGA3l43ytIljmN3PsXNouV27utkaMvk7FSvQpO8
q+C3nSF21T5mqOWNSvN31e/piEFslD9o0PQJ8FzlAU7IYo1LOvpiA+QaNQxn
8JJUTyQy9P9/5SmaOlbiLcfu8dW+YDlVVY5VX85pz5djNYoR34aWuhUWxa6d
tLIdbuesyfs/wivkh2UyHTuVRvtPNZauSCNoVj5ZindkfodTqUN7qmRj2AUA
ircbo2WbaPrFm6t94xGOZxzPwiNoZNXHixw18w3sxjSDjQbhDgml6cne85Kb
iD1Bu3LcOhwINVku+8X0kZkjsbFVU1Va2WJDk5er2az6ZDiphCxGuVHMyGyC
QWKHjToZdzgV7TGBkSxfzDfmbaRp+ofXejn/lbteNghuwYSReyWZAhWFRsdI
ecpddTWmJ1TAolF/dJF42m9Psu0QBHypWMTP47kx5sBcFg6uPRXLgKJw36dX
15PEqoCdGfnAU4xwgM9pOXVXuhmCHMPoQFvvUYV0Q9+lHum3iXCgzBZY9mr6
LH9LXWMMgEjDZc8QCylHnnPGU4ZJ28TkTFyzbVtDOsOLTJMt0PLxAxLd+6WG
HHPBzi7Z764mrso69T1b7twkQjBY1ggQ1RL2Dbn3GfLiM3pEek/GOQ4VBfJu
8I+jfX2okZ+sFpA3QJJTyrn4FLkntcHs34uMuZ6U1g/S1h9/DYYWD1cj1hRk
M4ecsJOufZm0zAREHMsENLlGl7BpAYK5AhRfB2YBfQoDluERXsutx7RcTE80
pF+OHF0i8l9AjvC6coZ0f6V4eAYiQXuS/OWN26xzC+ilv+T2Ywmmgd//OomR
KPH3iDuvrNViw2NQVbjzl/2xIlsSaCT+WU0ylI1taFTOtYOX3+xhu3FE77K/
4UFK8virNflHjF7SNnJteNxmYpTW23chelSa5Hbn4UnGTxx81ESqSHcbNhHP
BHvj0elRCgrBDCfZp0DlvCv6bvE0cmtHSXLuK+M01h7rr+0LSS+v6R4H2Txw
Xm9HboqNYcLyMQFJbYq0lp1v4IbnIdftnL+RneHHtlrDeNLm0UnQsOsOhr4b
Qzoqa67z7fPro+xTglT+TFlnCud6XMYtsqLH4tjLNyGCxHv2SqnEgxB9zcWG
NKaxiTKfoLjq6B0dlIhIn5j0yfbpjkikWqcWgtumd64ViCiDf4PRfgu4Ks8e
jySvlBcdqFfb0HscB2P9rQuF8V2RrDIRNzbgMYYxRz/ajuxUm9AdOaLViLKo
UXMkojstZfKugAtzQxMICHY2zHjUzESGo6ko+b120rP5a+RRv/uEWaMywRw8
fDH7PkFUMpCRcaNqyn/nFXLQISkjYPfGneUpDSimHbqxfYQ99wjMhtHUcT1o
nqWYtt2HBnsJfZtYb37SI41k8h6EXseVfDhF/hiwSSqXVhY8C74PkKR0P0t9
9aUWbYGMApa/16unQVzt92Rs0i+5sb0qMp4Tpf7YsVxBhjoeLYQhmlDxfMCz
lrt8G19kyymtChqZ8yXhcemGpz7jGc74xP7EDDJY4A3yP6DnjCVSkXZulAyd
iECPHq7NyttKWeak8JUC+4MynGVoGGsiHE1bkBoc8tBLhNhKaNVfXWRWPR0u
tTqdBBb7HMRPt2x9zoxN+ry/Fb37q7e7k8gsoHR7DA7NZFfabBBh4JCFKLrL
ufZFeCnDtAYHQH4OZhnx3Ktv75kphVIL0AksV6SaQIlP4BCNjm6XH974KceE
OFecnJK43UNZG8hZ0REX+449y51Bj5KSsCCZ53I5Ww0hSyR+HVtlw8ac+c0k
8VP6LqLdNUqLh8Bx47f1PwzoLKyUgIPjeZ7nkicbUrEZ0oTDHG9fAhnEl5WV
yfaCv1FOFZrYBwRRjIQnCuGeMrJtXEc+5V2AVlCTRdsjXwT6+u4P+EeTDImb
APsFGcfyJfjrp7d9wGXcvHWPAJlIcejgc1XcPnFpDS0+bYHuZ4xrjIDzexOP
Oly47PKNyrGVcmrYTgY8WJKLwEjbtkqjnh/zq6muA8P0Vvt86SSW/48uc1jw
/ZeHm+foXll5x7XnKklP4/yP4j8QaDj3zhxedBKF7ny6V1fguEix3pQXcKyO
a91T3c0bhy0IZ4EoFx7xQg4eW+Vv4KGQT+3CAG0QZdZ3uY8prJTJxamwg0Y6
fS6v2Hs8UvTqfQEFYaPgICVqrjfH6uCKJ7o0KsT6OdZd2IngGkptDPimIbcd
2olZk0h5oPHFYX1gqrDBRZaV5vNRam+dEZAux6B/7olvtb4mBIG5zhfPZs5j
EBsJfxQE2GDlXEMOPc5iofEpbjYm2ED0oZWQDmLXcAcqJ4qH15SfpqXX0xYk
jp1Mjghj8ZHEokkY0XvWn098aO6rNaJHVV4H3iZ7eSQ4axv2S6pNIVeliHOl
wpwzfKTqUBsKEb6gJtB2SIDcu8cdlwKc7W6juIFxNzbsk5R3jZxBGmL2DhyY
TNxshRq32GJPrcPVFMZnw0uWZE/bahRWiW1HhBb5TO/bVcHFrT7nqUVDovjb
gXOGiUVgdfODmOQP1vurycZU9VxVjp3yonAVWdFS98bcI44c1K8HlL1TIMby
NSIwZczJPQzpm16jAA0KU7CwwI+r3Apqsjjx7jWopEE1PIlTEAfhjKkm/q/A
I3wDK0j3WLZgFn52S6GcWC/vtXtZEwVelNRCoTYpdxc9wEAH7RAmDWFJKekr
4Z/slN+6EQooZl68ltO7DP+SxUnNl3khWCw9cfJoc5YM6qRprmvEyw0zQCdU
9t4uGPLUu0MeGd2/kAeHiCKBvloorGanyORcQz4cJU8jlQnEFt+Ywom+2PIf
fAlo1P2j6Z5wngAoUeD4YdRx1R5cULfO+Z/j+ek/nVuhHKD5QmcVAPHaiByA
UbSZYcAsvC5XebehcZNggqZhG3VDraKS/YCRNlKI/JE5zkJ7nAn4OLzOy91z
7RoDD5qdmkZV9pYPrZUcHCOR0OZXMV8UN4UOWcFfj646KUqbL+VCVlpSlDL9
9cvN0sGZnETI7Zxm6PXI+c4sQLP4+SyHu+gucRGXZZa8fBlkNR3It0uEwt8W
jB1vg76Uxfbsp+t58RPVoltcykv7m+kctz1XUndTAZQ70cVHiEnFf93q94gu
d4xFoELP0QGftGnsCuk9+mAEvikBwNIvDPw4Y+h2JOUjpUrPq2EtrHLowLdj
k4yInim+e7Sw1RAOnEJsgVE3ej17vBlQoJ+IyInF6QoqYzIG9Wc912oMgMwU
zlMja6TB8Lquxb+Z+1Cez4szzJDHisRmeRHhBphKby5Kox5/a04i1BgMU2S6
1JMsEtIl7yTFN+rsHRiitMpPL9EUWW7D627nGWAjTMLtDE7JCXxPJE0LCngS
4QS0qMkrWzmRYHTx50Yh12XsX20MWTUPTLWG2sRtUv1Hy2DVutO9a9AsX1fy
2dTLzpigOtnbdNM633SFvhYaslVE/uDzr0VUpd6PFyaa1VWKAtyLFLgP1IUO
7o3rQFeyz25OzudMYCaM0A2GmZvIbKvyQkB2/uoqlvaBmP7IPF2eVu6h/Qf5
nERz0m11XPts2MSD0FJ25A6iH4eRH9ttJ+d3WN/upAXPyqwbLe6Ig/zIdToI
oANsJjm89Am9mMq/nmpfrsTXoqFq9ntayYbzHRF8iKPuNr8NfryGeEFJRRi0
wox4KvpOxGZnGMvaf2SxHi6hrCRjw6rg+Qxx3jjY0FkFDJDlj18NVPyzjmHP
Y1kbAVxOWD3rt8JpB+1jZ5cifHyybeSkOy1/ZrPvsZ80X6GyLT88cxkTW1ZZ
HbIYcUYlTKRq7SEj0qVkJA+0Xq5v5kdCofu8h60coQP9i3+SRnGeD8+uZfxP
uvP/G+39IM+CAehRIoiR5kl53O70Us7ZpQoDq/3qBdyKdnDAjYyD1iI55hov
HtBLtzwTiK/5WoThUVDULqQy8BvzBxkNC0JSp3EO4voFo2qOnRIfPJHozNNh
e2BsxF3ErkJJ3e26z9Bd3jOq4sPse5E/blUFudEjLXgwnQ2uDG0rsWf6mgAu
5gAX2JUm5LJp0DJHu6uy9wtF0hYelhFJgGSMX2hyS9W0z31FJKtBwecc3pmD
SCkCdOBYIhfXw6dZk2AjKtxciZE+vPlu1jC6xafd71uLZlzsn3nhxDW/UODw
n1xVauM/L/jz8X4jbFrkoB7swQ+GySqSHDtiAh8Vhnpwr+1tHloGK4Uk1pq9
9sbLQOrS00rUmbT4KwthCe3RdY9cqEMk7bpMpXAUegnxvh711XwRPx7NmHW9
pKPJb6R+dhDEt+mZ05qKEabINZ6K8xZRcVr4+s1rZgk+bpFcBcvBI+AMolz6
M8D9kE5OaN1FpgIBicM+HY6KfO17lRjHXY43BQW6jNgT8IeIS2o06P4Yh85L
OtGcFvprASEsOK2WB4UZDIAJv6sjXwYrvRuXd0Vevis9uj5oPVJ7YbChAiOj
sQnXdbWSUd57oUl58BLZnsDQkY+FDh6gwRvNw85Z4ELtGunRouKxbAowleVF
LxLGSDZOqGHj4EGVmzoVHRzEC00RfbywSSRckXKAAtwLcSdkyFAQXGTWt9oD
t0PUeogn9xwZiUB9vT1Tp+bmWtaarCL/M/F9e3d05fPLNXpvCe1iAyml9FSK
aI2qr1NPexx9VueaqQaN0KaN14/5zgWIcQbDjq24LLvNmWLRq+3PjqhnP+rt
GSkoMSn9oMcFYPYPMe785bxJvbAM5OOMwxXrNcnak0JgrePBPwviMWCAKNSh
RScPsqUWVdROQJCi1mK/kRsPzBveYhuqKFDGFGfejcmvwDMb7DbVkisaiqh3
AQOBfNWaIOTlKU8tY01PwKnEql4WuPjmk5QGf1NNx7bIlTqzE3G70Nz19Lb1
r0bMSieUyIj/Uww626t90JRPexst4s2OhTwPH8H1x6DKc//pDx3WqNCAXNQh
gG+J5K0HuW0Uvqk8eLMpOfIRw6igX6yf3Ws1czVSYOLleRDuuxEBouNEyC9s
sv4iXPQEF+KHYoQ/jlHLPcC5no1/Nc+mkVWtc+Ge2ZZlyznC9AuzvFQVSTAI
2zhTvDiQ1e0Iw9NZ81CLSi2ar+Nj/fqF5N61gO75oO/H56bONTuu4XG5mwrA
jPxHCENQ85/t64awrxXeX4Zpy8N3i3M4ds72gKrCvfvJeSzuBgsDcbblExtR
YfqsYU9X9JXZu08p3DR76jSN0AhUddsJy5KjBHs21/IJMlkLFtQXAH64M4Wq
HZ8spOdBS9mDKxzJM4+AWpaJFzkW6Oj1eYglrXBpLaLW4zoF1RlDZwwJpIlc
Or1OmLDbt9sy9SBOgrZ++iU3BBSui9Im5Qr1r2ardEyY/zfkG5K84aFWZMs8
/1IUzuDU6ePk/ONyFTSq69t6hca6sXqs3O564auJX/DXKUj7ucNt2ladBgGh
OGJuSYYyQKq1t3MwiWjUlvAzjtauRYMBXp0Ri+lLdViUbXwJQ0253qzekNOM
MduFcPyrekCXLNI8rV59iqXI2T+ly0X0vDVsp4KOECfzyPb8UvgZ/WYt828h
s4nKBFrVxOSAemUJfE5r7K8L816HXVKBad+y0mUEAokTFUCKItf+ciaLIYwQ
anHoV7bywO6eqQdXDXzkzEsS8q+ND144oc2rwByvoADdDlHquXqhoL1CPaUb
VnqdQOFebR231O0YtG05DpXFU7YV9kj01cM0PSYbrRU87fhbJFg8bWa1hDan
EJGqB6xBUcLgzWFKU5az6ioQ8LAUbbT7+KgsGXMnCG3UaM+66ptfAa/nRY+n
Olh8aXVSA6zlLrdtQFzz+iqRldpwHIhkxxKsUFug7wMpeHYpLGHWxGNaVHn5
4O2sptiSMGuXn54YLo/NAYFhOB/NK70FBcJnCrqu81i59jmYjQzf/JOiPavR
Qyd9gf8R9zcfzlnGHaQFMzgJdZ0oPVq39iUrx8Dnd6MLVhyBBvciog9NoT4g
8mdl0Ke1JjiUY3Q2qrYuf6FCLLDVPBMcQP1IAno8jansjTS1gD4+bhPakuYe
GQDDduSgpjmJHlOpKphFbh3nCa8zOOJIKDpUG6gifKtjtUzeH1W5i0OrDxRI
WiHi/4ln81V8UZwRyvzpfSuKTknmt87eOFMICPouqYtELlCloYPfaBUG36LE
26uFMFlsrRi5r3xvRfFmWn/gWdslRxdVqs5krpFiJREAnX1VtZMKuYBnR9kN
E/3bkhW6rokdlEEFLc5xT/gpGh9za67HIem/l34lGBlx33rfjM8hALkuPM/K
pW/LvF1kY5gKe2LqL9BlNppeAUKCpY746fJ67FNaVG0IDPSwoAd4XFK+n5WH
IruCnFyX3EB9c35EaQVYOEd8Kxe8tPbMBlnDKtwJedOjW2zu4bwIpU0I27HK
UWUqCz3ZFdvMiLSUd0Q/kys4cwWOdQ/7Ipp7g1c/OXsgKgwi2zT2OoaiAhgk
AXCio9WYJ1Mx/z24jvydUPQ64iNO5BOgYVh3E8/DOJc+0Y1mjLsTgw9qeXEN
h/VGBuXVwDLGpApd38YbE52v0mZG1cdq8glfkXYLZwIgmUyK3fLfyc9zNddl
8ejtexRkMxPnLdfnHRW1AC9N3QYQMjv8wh+GlMDc/BxBBhiPk4oeA4TbYw8H
xeXwJvo34SOWe64wzYaGudPwZNidtP085LF3LObB6tJue3NAeqIJfnJb+/2v
v/BtRC9boEVQFx2uQilqjfvUXXDcD1XeJGJ9+gHbAVCgBVhtkTyqk1h7txOt
3Zk+426YaKpwxEw9lsHL2hvr/eBy1qEx7Kcpt/JgeR8DRrQr9lJBhW+8/QzC
8HegoJ0drs8EVApbuMorwozOIe3njki0oBfeuZ75GiRARFw5yjY8XvrfaQLI
qTUGUXaktLI9zcKvPjXvvzUM0foLKO1AOBuFSsimZ+of8ECVd4n/tam6X8SS
ytXiWBasbyRAtEYxmJ07tSFTiQNrVGeJtaCloIZI1tSPzuAyZGkLur+6q4fi
Dx4P4f3h5/MsbYaDV1b5KkyfdgLuEU7aL54PD1HjYSVMcBlG5mvNv+y6yllr
xvoYdiXCkb0CiKTxPIaPPOo/orBY2ivF7gwRXMnqjsMvanE+Fl9dS1IqfN/A
qeBPOksXMTkDCPQBatxGyvX+sRIrtyfH+8Sigz7sF0niabDe6QK9GUN7SEHW
l743mX4MTsXqcEZhSaddhg6daLQrd3TA4htdDDb1KiOUQoTt75FxyZzib+N1
VIL/ujvEXjE1daNF1/hG6WIKG9ImbZivakkIDzVrtg01kJ1ZsI6RVDck2NIQ
G2cgaGy0M27wfJIgMl4Hv1AnXFCu4BWzkYX21U+iHgPmwyUMxYPbvbeRILtU
zTB+DcgHHhPK8AR5R3LfXQFgdab3akx1BTFd8D2WKITRHluvk6SNjXg8I+qm
NRHsdNmEq4mbpgNseg86cMeiCRymlodLNfW0WzZZjYmJd9UP2ba5sZ4ZlTZg
5IT8N4wCGbKVcpEU2odA0Ehvlq72F4ka1ViBMT2Rc4vSaH/uQpkhIF+6QdBM
kjrDy89Zu1n6ifHvplJGgB3w70uZHToJxCb8W8QppKVPvHaahV8lsaHLD5fw
VtAXvpYJe8JagUnqJ2IgwGc/cB0YZOBBybxLczt8QB2zv3/i8zo4OSNr8lxA
Dg1Qytu8pQvMAw+sf+WjUDeX9JxsBmlLmwy6ctqzfhIBTmIGfY3ZV0FI7HMC
o+Ls3zXFsMVnHAyKP/MOSv1+tUn2lMZw7QV4mInloHlgs2/VOK3/A5QVVj7n
2DKpv0+qxDzB7k4Xf53vNU6ql+3i6LOoJCcupmjLKMCF16qa8qZHchB2hBJf
uipjEAqaMnicSuf2lD8GAfSMbzwJAec4x6cVCVHOGYBQ8qhZuRhKWEUWqCw+
UaMIp6Wa1e+ASXKZNxnZJlps+jbzveXoGdlOdbgeEyaiZYAxHujuTyk5AMt6
lXqnjvUUhvCmErfZablQpGTvgjuTUsleNLzfPZfNEXGSF4EmQsntJvLCmWw+
OH9C0qdCLqMSmgsfCKILv3KjXqcB3Dm5uep4ddtC5BpFaXxdJtStp8mEtlp3
hyo56ET96F1tD+GRCo7WmW93YW+4XRxsU4Zm5c1P0p/6brtNaBWowdKTQg46
tyCvyQj2WEyBgiWKEtMWR46wdAdnZtJPcWBglLh8clJSAUgf3ees5MLnVyQo
adCurSIjZjLuFsRCbCzSKI3WMBoVGNRDiZMmL/bJxY0eTK2x3/4vR1reF6Ba
nyMsg6MXSPmlW292PGQ1+J2k85akriz6TME78FNhbzcoBd34yIhzE+7u6VL1
TngWMrO97w3fWc927iap+CYH37+mLjYsurc7Qp8cwEBKmpp62n3LukN6fLJG
1rdRR3MwDPQEFurSysfaRmu0ERJSHVBEm2aPRrKCEYtfuW054uc8kS4h7M9s
Y2dcx6Yqnt2iN/IvnSAIG3vIrupgSuRgsxwA+UOflwxeJs7R6ie30QcSAwwI
vmBm99S7WxTARbwnt+h+ohlXcdzVk+5ZHbOBOKd3/IOiH/hJWMSEGHCnskjq
nI7BYfWTpkaLgup18WiVRkG+IyoPB8Pq0+tMfL7OKfqqYvWcEpyY4l/wQFjK
r1huYQq00YvBcrkvOtyPHBNdPvks6rAOd/MqQBV/y++uHrl4uMHCQuA+Cu5b
men+szWK0kDY8DZSfoO+tOzmiVwkmNI/unBRemxvVn+bUVrlpxN3VHqXpi2c
eXfqAGM9Qf6FcJX5SN39QM+UDm/tnkpISRumcAIN6BTp2GzJZW9tCPF1wBS7
GgTErBMMai1+WXB5IxC7odZRjSMfzrRtzVklDtPK2G+v4RWcT79zhiQwprNs
0zptSQxcxZtd9fMPgvm7ro4GokcSknCcsq20FlV9UGh9vsAt/WtB1q14HDC/
SszuiLLR3VCUdZA3/3kTgnRWnXzPytLgDiP2gjPC+Ab81i/Kurorf+G3TZVF
ys0LffdgXRL9v+KZLoALnbktjN9qGS5k2YFm5y/y9R8Lh+fztEvvyHNmrMC7
gzC+UYTcwl0F9vdfStbNPdwspGfiJWVZcfk9+v/ZPwi5VE3/RcHGY8kRS+BI
8AOzc8hnCIUZVZP1Giv5ABghSJA67LBIXMv8akqQgBGQ7U82DuGKxsybEZJu
Sb19XaSUhURLAQ3OU3CqNCUjvEZiGNrQyBAkG2lziLz1LVM9w2PlgR0jrEtv
1MzPL/C/hi8iWhJq7j3kKMpBU8YBQBy5TzkBg5bkV4JJUz9VxGoc3dvlPcDG
tHn3xvU8CgJPesELNQg48IP1w7WmrvVznq6ofxsIxirlK/91IXNqr1dN2oQl
uOb04S10/c/KVJBqufI6wpHb2HllR6ZJ0dpUZ7loCcc5fCBI+NCGDkP57bMr
wFow28GXB7G3mbweKTBcFd2vefpXJhLApuw67UHoe72MCD9tDDmPOV5Mplpf
n0y3o33CT7Ji6TmkJcJzYffr525x5r8GIWW4mw22NWRHHLxKvsU28ByImHBW
WkO5mWpECE1xw//wKZ6d1f9xVQ2xuBmvdSs3rMNt+aXwK5RyxImh/MF6vRSk
KlovZuviSccANP/3y+pNR0jubrw2IPXL+JV2J6pw3+cE6NLrhML7YemSxNXt
vuu//Pys3Ib8Noc2X//TDK8L2Rm5CWNb+sU07U43d3wVp6hC//igvJfP93Du
r0blRVqw3utSZFGvyQhG6XfDF3DrmXhGdK2rE4v+re3ia5A3odnVfevBp90B
EvC+0xoMaaxtFRgLqYeS1KIZUvVPyCJFISgam9THO2DJchArI4TQHpokFtCn
IsN4tNhvUfmBAPVNufwos5+jBIIy9O+8KnkC9tabBMV0LQYQdN4ZPvqHR4ht
PlUBYfhpjoRCi5JZrodPXdv6cqQcNVTpOzljmBeHYgD6GA+lj0Et/FTpkTxR
Bcy3yIRQAIQ1XvlU9DV1NwZII5ovdKnfHEXW2Hb6tuTArMCIUWgnt/JB06Wl
1AZ6obuqMkbgncZ+oDSJRlP0BXF4meg1vzTIFD+tVfZS13RRqpcZ8/pBK9FL
CdqbMrolsGAw7/ld1OtZGIMOtQgwDmm0q8KrSXV2w2gCzUFvGJP7i3kVKaO1
zqvBjv4NkUO6GCEu3J+cfFg93ZNsn2ISw4ciq6CxVrHEL/eum3NtpO3XZuk5
25NWV9uWruz9rSw46wC4eozKsJExiKCsE4aEGl7bOLjYgnEmeyBaJPP5Gu03
kKa4QIbw2WmPmLeAr6Lip0OjHx/RVfmxJ8bLmxqz9fZ419yQ1Wdnb1rFZX/1
1bPfoeDKdqAAWetAOLiJ76b8vpzCzg0Ye/hqWCz3KWakgdD13nytx3jvUJwg
CheDHhDgnsSkoPlPf9d2gQxS993wNMrGy+lFPTq6Yqk0f00D/a8GznV0UPox
iL15TRRVn3PwZA5LGxDdpANSe8nGksI7HKGXT5XBCiYWI2o7dXnU0UgCNkgD
f/YZDDQb21L5ckvf4OKE+eyw3YFZLFvFcC0wVozOjB7dQbVjXBF9JPo/OR6E
2YsxWg+ZLd76t6cZeNon7rltblBGw+YLqIEfZ33lIdn9EwDqKSLZAk7RID00
sW14o0hdlTQgQua5rmNgr10azGBSrCcHZiQ3MNNSrSGjNN519+B9RXoibCln
mvGe4tHwWavEI1lx2eHHiuZFQTm8qkDQQJO4NdSGX5/CipqtupjUsm0oBrrC
JPYd2nTA2/wLOR3sK01mBGJBr6UtDmTrG/6rU7SW36rXgCptCF2g2cW3nYO3
q4ZlHmFTrklTcXPJUvEF56SfgKY+c+0YOO/MKQf3Li3Hmo6GlaaIkoQeRVgg
jOasPVcpjkcI6sveer0QoAbFKbPhPQjDd55LTp33Um4myV2YzoWWuH2stp3y
Twp7NDzW0ASFbLEgHDP+xpFhIpksIiIzhHtOxfvTNa+5QtdsiWO1/61VNZNl
rtSygTSVTWWSeRDsTnqB9KRPRFBinF4ip2rYPi9Rt7DKVCQ7x503sxe8qY3s
ymxYp3i2HbeiEOSwNsBnOtnLrl30BQCcOpkrw50a+5Rx4JP9uCaC1tZDsPfy
7MwcgJ5lqeD29hgE1tac4kPHZyDRqLECaf2nZWdziWJ1I3YusKYJy66d4lGz
t1Ici3JDe3JrxOmg9I444HMvWB+lSUceQq4s0Oxba74yvR08ij1DF/0WMlKT
gNU7rKb5zyu0FOWaTrDWfpF/xQ+l3ND0e2nCedDySBM6cONOhOO/Q5MYXPrS
bg7w5Zcxi+lAF+z5znH1ZDXYoW6MBZezMgoJ8I39P4Wc9xowAvOm+w727kNS
HoYTW21GsZ2nt4mO/rZNaMBOWLlaKChnbBjiH82+HBqSLxo54Mngg6t1eVBf
liYS9mtc34It0GZMTkKXCvRE7td9/VLFtsKXVMtJ3Ku967qKoRHXtWHEkLaM
1bWKNJvxA2ZmABkvV7ZVjL0mPvIQtQfQa6t0SnSe0vMqLkuCIMgPqgESMJWZ
m5+adAW1n6u2IMKxIWK6g0SNKrvYmE7ISuVgf5nf8HuJMVlSqLv5s8tJelhQ
Si4S57Qj91YUOUbyML6ZQ8N+dtdaXxcoidZYkd0QqFj8Y5bQMg4pWEyCUWqi
X21+2ro9/L/7sJmqfRZhpkboIxQvIGLI7s5wmCm6nK5mTJbGl6Dx60qfrSh3
N70B9UvUOziiv95yUJZjAEPDjyM6qxyTdvs+z2sFfD+Iy8uIgVEaPX1mBFsF
9AJzpq5jodeXaspry0w4TpMdIQmOGW9DUcx/l+aYq9O3nr3Smt76CbjsecyN
EYqE3+8vrMY6YDk8B0ZeTQ3MAyI+MVpiFof4jnygm/41+UctXpiT8+3g4ekj
rGIo7LH76FHWCZHnRId2nb5MH5hB1j5hLGAPNT3H4GZN2AVmZ667SXML/FOJ
baDn2Eso9GyPJGSD1MohuREOljidlGoM1kummcONVCGQ2GeL7xxl5CtHBpIL
87EBFpIoy2PpAv8YnvQYKQzbr8fIJ2+nFxd87+OI2O0oRNIQmBcQOUIMG6kR
nkcWEX3SXQv6STia7+QWKC5alG5hRsMvzhPvUaVqUbN3nlN+QMLFb7ix5wFU
vWkkhkemc9IgsWtaC4K5cAqbEntpxaQi6kSJECacyI+//4R5/4qnukKriot3
yC5mZssZKlXlXiCHOhJk/TbSujQ9RwmdVpnNVpJr9xN/ZS+ETT8UjTxSxLRU
W7giliyGeHO+HeFXqTEYEGwE90GVO8/y/Ewe1fLYHmb3ne+WdM0XhUE8Mpl/
t5BKpFHtqXYJNO8QyzS5M6TIUklMEyviARLesAaUtsbVIwNiYAE9uknliWzm
5Pvr3qOD960AbfpW9xYMUlifFlqotAI2/8xtCCS2Ux48tGMb7TyQsRHTqP/p
OOeV3iGDNQo3UzxPDGUmBhll8oGSzI73D/6ocl2FO7riu5x5mR2Y6ce7PeWX
tPnaF4zWEhxj2fzygZ/FbUQZIZb8/KZR5fVZ5lpd53o+aE7lWGKaYA3dc69a
L8boyVxeytIPj++S+k9uk6YKhxnQbi5kyo9tShB6agPXRtu+gZtFNylkL9c5
yWHUi2oDLHSEmKCjjwRii2LWLe9EUOmJmx3UZA/DjTGpjqOEWqPCEe6ySMl2
kbNZskNSfuBT0TEWy4TEg5aU+fJc/saZA731PIk09I+Oii6HegfIhJ+TC5JC
MZO0l8ODNldtRFg6pzcXGPFYQoIf7f2KAr5egcJLFCSxhvem2g8gdOyozGmM
rGk5VVLsa7THKCwzKzedYZlMRN+hQFW77T1pqv/PsNsbaE5XpGH24rNEglGI
SbHSuyuMXLHLtGdmNV2GOSBAy1A472QjJvPapdTuBIzfYakLfOn8p+ofvT2B
CroUGvB8bHKRMoz7cWguc9ovui+VKMQOG4N+LNHQI+k4FB5c0Nh+KQwlWaYx
tc0M5cdOLAwbeCSFGrQ5/h1GWKnEb9H1sF0vWiVpxIdWQdqdxDLXM9DaQhPi
jmi0e+3RkUQSlbngHLwqfOAvBn6pe2rRqBxPPMCouEE4QgDbaWxyGaWOhcNG
MYQ2bfIDDKN2cRpNDjiAG4XOyvmef/j8WJsacdc7FT9DZ8G1DUNtxpDDiQNk
XxRbVUHz1yPsBnhybecQ6fIcQbUaXLfJNkxwE9UciVRH5vBF3swYPsMSD2AT
2MbbDD0OL06tnSOlXI0jWMfI/KaVxHNlwEJ8y8R+n4spstI4LDE5coL2mAdv
5eOa7+CQyGdHy8P7orT1ubel98MKQZiSs8blcWxX4w8NdeovffZLCj9nVNBn
dxCfxEzCl45MySewJaWqmTUmwPcSQcQp/FpqBg4T649UY0qfunRn7N2PpsX7
M2syEVAeOBJWeqVwARjn2Y/vD8CcDpEiJC9bkLH9mHrrb/LfZmCgCAn39YU5
uhu2Wns2UEMOOgsFWGcPbDRrV+iHNHOFrRPxmpmbUZBwJDidSZ8OYSn/2vsw
fGxicAmOpJKWLOZdj0z7wxrYfrPYDopWOkK+5oTcdUQUJh4S0VriBoJKdmnl
wAARLp+7VxPJJJmce1cGXHxc9NTsii9uu6LF13hrN50QyoZcKQ8d9w0WV2gQ
gr67muV5TwbpVDJm5TLTkl4Gn2h7P+gMIsr6gdSmZy0FNRcBid6+ZUHi6pdC
Mv4Hahu8/VuhDWUQLVoSoSQxV80mKavmJjOOqSCUrzVkzUiK+bjyryf/dvQk
xMU9Ra6TKSc3iInYDygYhAaxWsWKK4KZ5yiag3Y3fVVYZRcvrmgGWNMQp2dI
xB0OMQdoh1X3ssLrSfp8oGTUzcnuY/dmFSOnF8EWNuI4irdnyWE6ODWRfCgv
yJyrMOa1ry4K26dmsCEAMvqAFBIwdTSP2NmRWP3a5nZ57pWW75/v7EIpEiFn
5c+29+LyvOhV6II22iqxA+PG29+WHAj8512Uq7hCPY/kqq/T7WDgxz/jP8AL
L7lZHOxo617Uu01Ro0wa31GokxfZFvODWcyajn0cZb4rWikH0U0LMtDTXSdo
tRol07tkqY/1ZnGNqC2UrH5yChGPvf+l4et8X/ZHw9af3RBaM/kwl/SCZ9Ee
q04BukEaV38WcZKY274+93r3pLTGjfXz/QSmQ36ka5O38AhlWp9APLgePE9B
IKnrFQvsiaEcfwJdoHZskNpuhprUpeg+1wqgbBvjNTNiV+7omB5BW4q5Iln8
2r/z+48pXpnJeHiDJ+0yv//VjF/mCvKGDy49WGXzkptlqvB4dXX98LGhQ/68
H3ecJ9iK8MtgXCJf+Lt3aLnyoj6vcmgKCsudAyI3SKdy/flvVrvC0u8AF9lp
8RuGDBaQr1zhXhTqLf8nrT8BD83GtyVyj/NmCq8rfzWy8UIS9XhOsI0lht9R
xnSwiTNgzSYC3NnRJPYMOSyJlFG4t1xAe8+Erfs4E8jDUhQOgvDqTX2sM8+U
rhWtMlfEvDGBf0YBUbhFQnuPkBhm+WGyMCyWBbH0JkIcwGb6vBgxiTofijWO
hKkk65owLSBaSRHcqsgqPBXJMJ+XnaS+aV1EBujWKD4qNvzbQ3cmBrp3OR12
qp8sYLGb4hhSZ/29NDpNTcA1gs407yy+HOa3v4DEQtddC9pLzk6JSRvbjtDt
o7lQ1ggOGXWC3a4G2b+d1EbiVwgIEUBGtA6plZk7pLHYQ6ZxbVQMxt2GNy4Y
K6SSELsVSFystMFC//MCEBwebmPvKrDICf/ckqpiXMue61ICuFQAYyS4gbJ1
zIPaefQGv2zYUqJWKXWb6X/7IYM4+i64bJoSuv989jdRghFrYgfAQb6jX2R5
iM02vOB190BoQ79d4RvAwwLAe99yWpMeHtw7f0wfewu0yEZWfwvPk/EwZ8um
k9PRk9ngi/YAlUT+ud2SuAOte7q1hK74HO0v8MpUHbTV+uC8YOurh/acJTza
l36U87NQAfN8ZBv4mkpl2WPKmCGgWqhVoU4Ih/mB9UzHKKIIscHHHZn6R5tY
bqo4I88RDPMy+1N7frNukna3IZTRX5+qgdln6jdGTL/+NfFbrt55y4fskciU
sNVHP5K5uDj525t+GGzkM4B3O2PNz9JxDkBD5/GbS/hB9eEJA9vV0jprYHlt
wA1PHvpU8gYCZSMau6nTvgfC1zL8+05ZSd9gL9NxtNh5J+djceI0sWCBm8ji
0A6jM6zOsFAErYFwz0Y6DmbXSiQNP4q6BKDlKjOpbH/u6duM96aKE5BhRP9b
UFMEsNuoiifnNOlCWZDG+kfbZDBj7X9FTZBr341whNGbt0j5f21JWR4cXqkM
DtA0F1THX8ldpjnrDbb7/gkY4UDHCku7OG8yY4brk7g4OYyOLf/kN/9Xe6/A
H90iQGdjauyB5Ok6Dvyi1gJjfeKBWbr5lz9wnvDmnHEo8EiIicN+8qfwyIHE
lfXSeiF3eob06bythwM5ICSGIUoossMSvyxwBvzuWwaJNi6pIu9pAWbePkID
qbwghZmb09L5MoZCnIMFcwavrE8V4PjScYCUquYDdr+IzzVUC67eIbeW+nNy
D7oBBkQ3RdGJpdcwlfueEv/kePPn2cvUpRCAMyuUbjAo45Vyj4hL0yrtoR0v
YxZvGbEYiDeV07CacIK41/kluRPt1YIsGSNtNNBt8iABeHtNu3+PKABV+xxo
+Vci/JRSf2U3Kv972BT0pkSqL7I4SKZ7qV70ELBOxABKgdNWetXqq7lj41SU
SNXXNeT8Blsodu1JHA1hhPqH5N3LaeM8Fvnw9sv2xR3EXKglT8zIlI8V7e0J
5q3zd4WwUpn51lfw/BdWMwBg7NafJHnhyFhN3Mk1F/jhJs6SbW9zFL+EVdV4
sAJ72zZ1TF3AeEHJGU6/q7c7OnKLI07TWYQyeHKy4V8mho5zheYlF3LaUiPC
zmRBRl1Wx3PxtzO+f/F/No+/FSgJByag/DU/dDK4dG8id6qVImiU6nBtzYr8
rhlyAYQu2k/EVnPpt4MXeXR5R1vaaL9NQ1EWmHUniMwr4D5H/BXvvqNKERyR
mbRFOeyC3nktQk7O0Y1X0SAGJ0Xe4zsOgmig5fHc87bSmIApmlZfBb/AnlEQ
+H+l5f+2dMS3U1MyNgtMjj9+ho8aTAN/Jy5aFw4FjjU6IoZs00IuYzdFNgrr
ALQ2Aa3OZAU8NFT0PX8N+N7hvLzty49c6xKa/4boc4jPedFR0WFFvF8WTlNj
1nSbwfMVXwcrKI3aAZblT/OVf2kRYh4//FRQpzpw3yaRDw22OEtkNoBar7fk
qHTQ834VNU+UR0SanU8uCWqLnnMuH7UqjWjh6j8bZJcLQTAXGxpcfEiXTUwb
cu5s59c9BNo77KfkRQjZj9dP0EFa1z2Te19GVbg3Ljj5MBpCLdqMsrd1GSk/
0SxSZEe1e05Rv34Vpk4CtXS+aSv++YY76pco9YfPI7hvSTIddzOHNibxSa9A
tstAKCJPCfmAYN5Oad3GEy5U1h94dfQOWzGueHOrO4GR4Ehl+khz7HcyQQoS
TjvfwJRciKy1Hot/nm+Uyd4lirUcNgB1w7nunsoC8IkYBA0X6XEVpUaerZLH
nmryA9dJ919wbXlxb9X9tCz+ILef/6OlooBM8Pyn41PnlytVXiZNEUEJ7tjt
ieI30wEXYN2B+H43y74tRw7e56vahsIj3itxaiK4nWECp34UZLVMOFhZS0VN
Tas6YYV8R+lDrSQIXmHrltWW1f1znXAJ5Gc+k4SFBh/0nEGqHFNIEk+PM8Ur
sWURhU/PjGIuOn98BHxohW9QqMuCQt9j7J7L5XzoLQcPiWfpOFdcs6avb29o
kO6EMvUkZ1FeP6lkJs0UbZ5Z1ZExqNNUVU4eWzMgf/osLCi85w4JEMCmev+z
g86zm/NNGUoZ5ZFgFAtVoHs7dBq1VF/w4VeeQptHCHNqDF0nIuNHdqtXAK0V
ub9T+saDPU2J0iItnc1Q8o+seU/6Dv7MsRy3sSaN5Ii2jC0PfjHxP8YbIytp
DG3gVlN3HIjNOiYpil578jXz+F3x3lYuB6x3CwSF7iQanZpC+0hM6LLirsBa
MiAZCjYu+BUbpkJOM0MqeZAuCb0HAGYTT1w29GcMFLjStG5Jhl5XJAk+/Hg9
VK44kx/q/2KWE15cGikfJ0I0P5/yP5CfAfAhJf4j/dnBnmrjV/ypQ8aKeLtz
Fv2WO/MilCMhVkeciUv7lui9DkJYOZytLUDSQyWSArUw8afCDRa9meEWMwMG
Oczy1cGhRxA2usRX3IoqAUCywwJBq123OG1mSqc/AWNHQPULbA8MwfF0lcFN
BD0GF1A1Ws9YBxJfyWY7OtePBD3obpbd/Ls7zRrYUHOl7/SO6Rne5WRnVHI0
KWA1z/JPEQwGWKo9NnIDxW+iFTiu6iZ9nnpnLEHiVZh8QTGoQMbcy5wWfWyj
RXG2h3X22crKWO2alYZjrzZWnXkKhKc9LVMxajK3Pgu8pFIV5JV1Zhk75end
K+JYhRZMzvxyArKOkSYj9McXJ6Y/LQf3xwLeTuqWHx/pDLMBk7q4OtLB8+vN
L+zJOEFzL94Itb6Z0AR/732bfXhF8MPayDUK8ZBXPfUXKDfSUKvY1+DwN73c
ku0JGqRETUT7ThqYmVxCdauEZkJW9ULw1NzvHS1b2PiFYFhZ8c2EfnnzGokd
xW/qSmnCjJbzh0emsVZ2tSavJveFxnMiIjiP1V5Ka4HYbXRxEBIIoH9RviHE
8XC5Z/3m3hdbSq94VyCAf4gf+bbxXAtitf10czCBMH6tGzKSBlxK3Yj9B11r
XJSUJZnWSeGyfTmS9e/+rU4D+S/L5t24g8bxnLKiinWqD6tq2i03IwFsG1PB
06w56oZvGh7t/HhlnNIZKeH23ppMPxf06eBLq5x1nrjJrU0t4vxEg/Z3FHkh
ZlYC/0zXH3Z0L7/eMCHzVvXLGDocPJhQsh22OgYBx7kJji1YhtyWiDCHtp/H
sQ3OAER9Mf0y4i8Sxc7gtDPcxdMlXuu6KTie0TJz3JFTSqSokYuKx713X8h/
ch/Uw19X3bTcVPe4rJFXymtU34p/zIp2UthJkk5MAThpvz9szAA2bT0sX30d
8HO1SB6Ciom1XPFrhcUyJ3WcNoePBV6UZQbOdw8l6gSvsBL+1FCe3ym38/7n
2h53sL/R78YZjXd04w012U3GX3cLByJ+M/CXMdKusce1EGosGI3Xi45tk9sn
96UNasRHkAUS0qQwlQzWFQyt6cMdC+JDLUl4/9BdnKkObvILxVIIsbkP3C43
kb9odlw/f7ZV/Glh8LJkmhgGcfC9ps4Z34X6GDFtMhECrmNvB3C2CFE4dU9p
Jl1qwNB9/H0OADeAHXoKDWxw+/oB6Qpst8K1ZZsSZQwL8LKHRkpT+BprUfi6
Zjd+6OMq6R1fUuA+o+VN3Ewqz5U4FULlWdbKe+ku+qZuh0VCoeXdedMAvPx0
7H9kA3jlGvWBOGZbY3vTnujWS0eYnRwPPhlx9YWgzGqWrPKZk52ieAMR9dFD
f2CfZN4X+pd7JQ0C79RMRDm613AFfdPrPVR7qREtXzPUDNvfrqciviK0wTjp
5IL3JyOOIag/vIUPh3c55zoHrJMpLBFm1joWQxQsvN1nZ/kH+1e5Y6BMk0Cs
xeJe8aNAUHAXMQqtYGSbvzOWhtHY55XYpPoJXnTNI8VkY/qThhppmvJGmxpT
glUobGRa+1+0ZXAzPhZ6ptoeIbcoXO5lQ0o40ui9+z+/hmReqyKmqPXMyZdx
D4bBGdnECKNhN0ieto9Nu/12dqwXD/wNBMIM3RnoY7uJhM3MaTmJ1O9yUBTi
BThbFOGTT6oxhn4a0jwDm53qoVS6/g9ZklZ+BVBhuCUszPdyLTQ5CLZUsbHI
DRza+NI3etNhHQAg1SZegQTH1ydxXu6u4r9TTjrSvKpwtuBwuy1BH5iSHefn
OAh5WvjnEnOtpO2vS/eEwV2XMk++u3ZDshaCf8SrI9F8QJxyFZBPpGD5Slna
PZ9f93QkhhLsWnn21Wq9tT1n0/gDcgujXdNnM/NwHZYUL6RyrYI3ke2ErMmZ
zbQ+xaN8QkrSmB1ScLhD5sWSDVmhk5sWLDGHu1j0UJPnoh7mlYNlnM66i2ES
cuaRUmJ2068kqdbd2QOT7wn9V2BC9hNhIxoSmihKz40fgxyJpAUfDbtZQv1W
MK69EAf4b6Wwdqw1fBz5EFB/HWs6hgUdJ1OerE9jyAaeB4MRxpA+1ajWrfxe
J4Oc5eobS3POu964yySQpr2mSLCvtjrSRfHddIgtPphWpAIKg1Kz5c0muClg
9a5r01va9PkXd2YIKiJFiqQ/HiQz+hGsuPpiN5xDd6Gz0diQmghHmPmYuHjc
f40oK7BDpCcmE2mWnV9DQ6vodE2/Iby5jRyq6xvnSmkQUrq2XiJ341Ahk7DP
VbUxQYGVePXXFkPrdDyPZLAZM81c7pwzdV7nlSaGL1WUmekGMA8L0X9U5Mwp
13TZ+0bPp/tUYYVRMi6hWWafnvfyIeLmUoIY9XkPDkz7iLb2A2CBsIr7GZxC
kUsP7g9eN6L/qNrUZJMluASnLhB75AKm9GlUUFa4uHcDx7URcFyXOWhyoYzI
Woj0ADmVw4RjYl+PEd5nBuCgTDYNimnRt9STWVTn8K0Lp0bpWNCgj2RPYlMe
Yr7aPPgx8uGYuKxf/wpyQ3fwpPE8+6QTNlrSNfHH9YXb0jBdzw6MnU4byIyy
eJuvCM+pO9YmSFLKyRsBg9Xf5Q0IWKk9yKfp5XBBE+DHEp2wBFZNRIiJgbPg
mRVUy7yx3CuVEX2VKezrxUGTQwcxZJIEMpkgX+YtijlmNliFw7f6ExTuo3kT
3c2/jZqIe4mt9eqKmrbzX4gYYElQFZyXn6Ek2DlxRKHR4x2upCZe/QNZepCs
J/rpY/GIeuxXi3W7WnR/yD/rG8Y25+0026ZDnpbTIXxwSoN3f8N14yVJDQPf
8IKDFdlCjEBPycSiJ/FDWYMXGlifx54JxVcQzhoL8b+szXlsOOtJkl6dT+7q
YLPvPRAO17LfEg0IY7C6SBPyuh4+Gc6t+Bn0iFIblJB0RkurgKmbQzYnni+C
oHTE/bM1visE1CNCSIgpf4/rtDM49DNqHL1DKOyTBsN1R8sL8U9UGL08Qa7b
HlxYj/KzBDI6Au4ZZIN0byR/6d4MTIVsUJA6Q2xxYziM6aJKsW8niGdHLCbo
Jy+w7Sb9PbYozEWsRD7mg9RKMfUjh3IjxAuQ0R4TCJI4Br5yJXdZg7L/iIXS
ViSFmPGWovXl5nTceTTftYjEZCmpN/HvvRN8f/MSz0esNRMDiiC5yGhsBbUq
h8zvLr20pWwoUIsoJlXAtNv4iBWarmcGjde8eUTVhd3v/fJpQn4Aa4Rd4DN8
l70c8SDGxi30fvraaPe+Xck6oSfOvfwroBQYFhw6BJ8Z22yyx2H7EEXsyc1I
yKv/78SwZgINho0zKnxmv/6OhhPpbm/4C1S9ixlF0yPoY8bMRUFqYhI594ch
nUAH+NcQ/fI6rXTuTnEOihX3CwqBcwclNAxn+J/EZnQKooO5g1maqB0+nt/R
neImJ3VHiQXnL/3vPcdnC7WlS8Am0ZlAvBOBNwAlQYmn2VyA8g3FCwYFTZAI
zOVNE4ADSTnpuwPFGuPEga83X4Ay09s5gyZQ/s/ki4khwSPcnxWN3w0jQtEQ
hbWJabubOzxBmvhsj/ljYZu8RUXt+FfsPQGIKUoBkc7ph36jwGRdAHquVcha
TRJYPwNALHmJydgAyY3Ja5a7mGo6fu96qJVhiHoVoS/6gEBJuAUA0tiZjO4R
+THcM+w8cYDICLzd7ZymJ9N2KhF6DOGvMdmNMWHBf0C95pBLXXz5gp0dm5tj
L056fd/d1JCTjEaI3Rao4hJvsWY1eNtDaoaX5yh9cI9Luxq4eRDdb4oA/bal
55o1ENg+7lPjqh4F5GY5nyJNiORxMqjR5BdtNO+OTySjzW/IOfdBQolI2SeU
HoLYzNasE8OKzgoem3c+UjTmclDVpE9guYxfesiHFzbvlCd1G/BGatTu7BNL
LyihFMdgKgUN3z91PtjRP6tbhuXMEWB7lf5lEKmSFxRbebzeI7BaONYYqmPm
MISN6ne8B4JfhoI0VHRNnI2QUwl0UoGErcW40x62eDKn/5UaW3l03PS+bOJG
oHOat0dEu81NqLnJVoJ+q0AgzNSKSvSb9d9d+N900q9cK80zVa4Jq2FE/gHz
GuC5ikPPwASOeG+zkUGqYjgnPwUvDtBsaULJeEdHhZ8yiAbKLIJRqnvo24pf
BTAIo11Uv426EV6C/Vp0dGcS3szLwDvtdGb7czxjMjh8btr2h7ejXg5WuclN
UA9Ul/WeQSOReQHilwYqkS7aKzcmmeXeOOg5fuyrvV4GqijixW+TH69N3i+K
bwjambVnuUoNcmwl/JGylO0L2SIZy3BX+aLbB7/kgdS2BOSbx1zNw6A5ulcf
8dNNLzf+LfI4O7/G1txtZ2oUjFzI84sOOyCa7m7Wf8NZVFJdxVi2wKi5FTzu
NQLhD3ZURE6WgbiNnhJNUBYvr2Mf0vkBhmTvln3WbmvDKiyEUnmCNQP8kslL
7YS7hHFcHbzLFvy1UOn+0qUnRNlahSi4R8xwMBb6wzXsh2fQQmZxQK39sfqT
8chQvdWa4c7D1WOgqzqxHm1pqw/ZWUyIMd1Zbp4Lm4waSjkKxEzOmha0cbLs
Oa7SePI0FQiPDNKo6hXNfABWC381Sk2JThtK5T72yJfaAAy5Zz6AVoEq9J6D
35MZSaOojZNSriS1Yb4DLmx5No2qvzO3KSY56ATLWxi/nXf8ka2rcBGIKSdO
BNLYFL6j1/ILditJCv0DbrkKUED3Lmtd83+0Nl1KZ8cAFTwSVpQsMLlD5wQX
4kGKcimFK0feWPTjLiTqRFqPJ0TcZdvRCiHdf6i86DOXVzqSpPUt+D5YD04e
vtIGADHtgm6ooE3hIH7X52dh00jCS7F1yAm5qHHyFBDygR8/hvvHTkCORNB7
E3upMDpWtxl7l8if3FA379V/klkCfMw6lBqY5nstx5aEp2cfT6qyGFa7LLLv
7G9WSJcmaL2LPv02m1JxwU/EKH4hD9LAY7n4DBSg0bC9LjkDZ3u7mhTc0N28
QMEqTUh7mwGUhCnnzZ+pZL0whMDxZT3ZmHYIIRxqWeyFN9IkKKadX7tNua8e
qesYcPlkNtrMdYpKf+qybDvuzz1FPppitdi+6nBh5WTC/IMazb9mscaM/W0z
T9nw1Ph+044ldgBJlHnrH2bWIgVEzmx+SUK6UGqkKqI9mxKpzx01u9H1B4hW
GNpaoESSzhzCCL/4ZpZ8svDtVZXO0dWbJau+AMvQSMlePS8usparL7N6Dyuf
RzJr5FsLmt6EJBNeWoSQzem3WsqjETNRR0viuOdvaLWrgbMeR+z+FqHsBeOv
syoGgBlbhwcFJbVN0LRDmTn7TTC0aLj2BjYkJyaL3gQqwod382L8D/TEf/x0
b5xHP8mv8rt+I2GXuxi8oDukBfxqk0Z+imeESfmWW60UdcmSRp4rryU69c98
Zh/sARzG/Ja/8VcWOZsL6wOaq31tt1Qa6jTh5HdLOGr5J/O0A9jnsvm1HXv9
xORKr7HRvurPdZ7l/a0SjVjdz4m57ZOTs2XLWQqzUqr9xVGNFZqBzKRKxOTZ
WxYqSUrED7uaSeOs5N5ilxXQ1fVWEjpVII3AsI2C6GhBlhAMcOTYgOoMR6Vf
qLcVmzdJEoplgA6ILNKXE4OO7nMwThb+UK+nuLn41RK/NAWQSsKE+dr3nDmz
00kktYwFFLAR5ORp7WqBZBdopWQ2yrD+qDuB6C9A3QsJuOecfJsZh8ERiikc
tCfySLGNjU+ZZk0nnGXmstjvNbS8GeT5xenYHroyhu6dzFcdQ+9usveZsAQ3
3weqFHryVVSSe5CULM+4idha7TVOa+j5Orrv/g5wVtY8O4UwPDMcblHQNP2F
lL+90QZg92A/6QQM3eyX2czdk+iKPLDyiUZULduGtcT7azUcIKORGkZuXiQE
QlBvterXLH7kbtutREwYIaBF/6pYf4MpPRMct+KsKbsNhN5EZ0B/M6Mt99q0
UQMR3j6WpfYtKv4WRdD6IlZDzBbjl4PdwjcdyrBY/rT7xcO53dZcaUl8L3aD
igEIynGeHSMxQr+6jFzw4dSS/AxowjSuBach1wCZw9UvWEAeyFoRk0LmWhro
rD2ct6dStbFw0tRNt25/DW5PeLnNnLmlcNLKaeAljppY1p5IKuJ89kCXCYrV
FP7vLx90WzZINzQS0K1i8c/j7C+SnqMcFVMttaiRrGgnEUPozR6KI7uI9Uub
TzAT6ZT6iZ8S63dzmfiTW1ZZUeFnBy+2QxJTcm8xTKV9vQUL7m5ppHISw5ZN
XG3w4qS6rEF1hseY5iyINJ6h4bk1w6keKfSlMHSCMLiMHozQtW/vN8jt8wrd
psaIbg7TN+C5KDgEzS1ZM0w357xfhDrt1liqF7aEIVs6ZfWhyMPGdMd4LqDz
/bnzUStdjbvv8aKJU60M4HXPXqnobbkHLsnrDuwJOOgX2OYH27g8DRR09KG8
8DR0oRDGkVr2aToh3WhdhFuyuRnaKLylJ46y3u1vAQ+k2qywwpI+yx0q2o5K
bn8qauzRqwp+Ud0FydjzSgf2XvdM2g4KAI8r/2pLmxC7xBvourAOd9hJE0wz
OCYMyEXK/DitsxeFALNd0XHGox3IdpUknruBKvKgyFcv1Iv68Iub77njKCdD
UefrT0LBmyw5ehCcnAt6gjw0oPvh/wuaR3ohHAtp99ww/15ad2oCbGYHOlHy
OEwmX4LWb7ll+r2QGhhF/bglHpnUJwR8wCOFI5bSgAy4Gct2sQXZciEA+v0k
55VvVT4Lou5ycd896g7aO9MKqV/D/LjDoDUB0bx09a9hh9T+tkJxvTbGhMtk
5rXWBKKAf7sts02wAIt+dkUAZWBkaagpmixvJqbiiwaCXyEN1D16ypZTtq2m
47CuCQ/V0BqlTXuGuc296HcCBBUMTgHnIJCweEIMO6S04lJ+ng/Q4Cfgblz3
hYQoP/X4KpTY/SSgzOY8271bvviUWp/OznFSoUPYq8mJDjTyDD4L5ayvkaQa
tfR4rQz1mbodr+YLD0hWQX0nqLhbbSog0xYm1ZvksYp0H+7n4h99N8XNwxjs
Au5Qsc6i908qC6wrgg6HQ61MfRqV8Qy4AaEEBltMO8wV8uxAN1vmrDGoZs6p
U4b0Std7Xx7D0lJo8zPvuXLzLl3VvrLFYKiQp4GZAS0WkJQS/ufl8OF/HZT5
eAi7+zJlhXyFFkWiLFgBw8Z1hFZ+eb4wiN9GzdJ6Uj48Xk9A3fusKUEkHnDP
6tdyVXq7uFXbD/IHRrHAHvc29XyLr7uayMrp6218wYrZ9L0jb6TpEWrR1b5k
zXMkZ2M9vMDo6YbXYh1Hto66uc6PBgDZN32uL3CPAPEnEOEZ91TPU/VfdeIh
8uJZQxKmRmoirz1eq35k9ABloC7xyA1PmnzN5+yzMc558krURaXwhT1asDLV
Cr5eSg+dOfr1T4cIDsrfQKvap5qxT/erCkcnMi8qa7j2/zzny+KDrDOtZhIb
kwsycg4Uu4BimHMLze7LqRxNdaR7nZdfX/+xJsPKGt+C9ZylY83Hvf4+n61C
aK2QzPjjLe1xBHANetiYb/YLYEi57zaa3VubDKPs3TxWtvhlwlsPX1LrdH7B
QKO90ilNL6tWiN5ONnleC3Ip45d3dLDezjPwx2P7PspHstPDle20f8rqaid/
lF1PgfhNqoix29HQXw7WwcUfA40riSF7+IAeHNihQPFtLlHO1VKRIsai+CBx
sf37o73hNYp3zmL+J4O82RltvtBUYlDnThdZf0FOZWM7hKQZepv4ePIxj/Kw
bK3pSBB5+ltaTniMvESeIxdUQa+1b8HNYt46fcCfH/OxOopJpL3yyWfn7xsS
nPDLGehqR2UUPyAslJujN07Cc7gcdPgfcLgZi0t5C8PqNHmsAuymW35knoNh
dIo+V4fTQd2GJQhw4tKW9/Q6JBiICY8sRLxDyhVBhX+QJfWJKvHSIxqBF6D8
FfYkBN2tDPCzBgcMv4XI02giB7ODg6F++iG/tfIS+aHNkg3SlF+ZvR9Cg/2o
hUTO81gxddcVDGowum1Oa8Hth3BtvgMkS/bY5JTdHmtU28PSK611AJjgpKmx
7+1VzFTpSShjwtbCJ739Ns7d5+Z2ijQ8z2XfEA5PG8vseStLY15dKEHtyQlB
JIIes3eScRMc0+g7N90wIBCtDUPcdGpoInTTQYtdnJXGig3b7MLttujwSa1K
z80U5ViYFCaBUIOiQXhQTj3ppZZNlcrlDZ0j0JRhCaftB3qxCXnQqMTkkTV/
KGIwP6X9F3DknxG8+S8eFTUWVANKF0p0tytxTDuI31Ktoz7R4bChRt5YWGWc
fim6GPRrY2x6q0wAS7AflxO+HjCrNdbvfVxPJ7Jz0WL3ohBzBpXs+E3SrMDT
ipU4hEt6mfCO78xaSi1yjHoZbOJxKxCAFwldsYzXXKmN7ZXqeOZDQ7bJMxtF
3RjtcFu8gt9H3DhF8u1/DfpBvq0CmqOn3z/BUoIbwhgpsf/S/XlTwMgbjrMk
gZYrNzeajuXPyKQYpbQTKwTCF7B4k/vqtwjcypvyyIpWYaY1OmUpysrU/4Lj
qouNW2lF5t+C4Tm7c5Ncv6RNJTNRs/vnsbn588sqbC2eQI2VESC8Z5NRO75k
m+r5ShN2+wmnQx1IpzGRr4deExUBuzyX4gY5rEcAporQpzsod71bZlf1lMgU
3TlvNO4VY3N4m3nUpLFFKZOsiav/rBkgtcy72lkYS3YODlctPF4a8OnYHt6M
Gnfbu/uul+So7QBFpMgvFLPkFit44k7pwoXKT9YoZcVA62Hdxdbbet+2lZLt
ixBzDs4CkzmXFeeP3c2jC82S+apMkw4lrUj87PGWbCLo4wfPqURIlrc2v97o
5Wzi8ZRuvHiivJdPpStPqNsUfGqE2yOBy4wqntljwibZVS2QnTpB8wYIciwe
19tu7/0neJjUD0oWQFzbI56soucgJ90MnHT/mkLYTT4iweVQLyfIOhgWz/2i
c4pekotnU08RL73XVoCqE2jErO223kp1fq6WzO9rRAYPKkg2T0YVrK23WalE
cu1HmNfhIE19YeM8P5+7dsEBbO/wW0zwgJsgGetilj8yu8XeH5mNJoOPzZvV
PySgd1Yjsys4sKY1gHLlbfnpKZ/sksteUfKzF0wxf9oQRPVh0qPnV1rHyHfM
3z4/e/UK7u4EPBH49NggyUvbqJ+Goajinq5zju7JFM/4c+W1FQUM+GvoTuyI
SYQJ58MKHKAK1kOcwzHDWWCgDeRs8N8hrHFZtUwAm4fy8hqQa0f7y1h+L09H
zlcWIYtJoK6GBO+5pYliNeXDtT+ZKFb8haYQS8z/4X78Wpb2JKn4i9IiaQed
Zk4Yzjf0l04oFeXJt3sMaoyl7+aQGClPS//9nbTyDivDKRioV0lZYW3NlVXv
Rbi/eF7wezNIAGrTQzmmr5ELaSo7MA5+aqeSATcCU3dasI44TUlRpM3sleTQ
srzCbQztR1w2FKIuDtvrZD+EOzNBJRsVokmfbQo7CcIBQzLgiMS0qYQf6wc8
uQrydoWnTBC1x6nO6GpThcbQxutEX8R/LrxfDNqXuEZMPNwZkNA4h8TQADTs
08JPKmO4QDb+Hp3GwBpMAh1EX4IetRXz3kdHyFVdD0mUfY29v0nma6podzqZ
CdsKG9BvbMMWtd5KcArIxYZqDzuKxOi9onIW1eG1dp5yTHQdDRVM+0XanN+F
EfG/LfkSnkyAOpow3zBCkbTSuBpN5k18WmOc+H9Nm6b316upn2QbVj8MNVYA
27qvW3fQyeMc5ySs781uQ7rFhorKSPPNswRwe6J7oqjiyx+Jvzqp3sYKMYse
xzVikuiMeDeaVkTTslDoD2OJew9mMVaFMJJp5ojYQObn3C8huJtFcHjfk8AX
+/lbPhSrO948dfgNRks9yop85WfaQLpWy7XVvsKqEzDUi9QI8NgwyOpIJhN+
9oJ7foPn0L1HCXSHoKMcl6EURrdClSwgnZD1l1QZvsKrZZQUpfaRKMjGH2HD
t4MFpIbQqzV5I5n64dXq6B/Lf5cjZaAGW02Lv/KEuCDFEhKQVqZMxCRlD3iI
zuksujXnkiU6rJPVCZTrDTH0RP0CboUJOIDXz880KwyjW+Jh1vd1YQPdjwBA
jNiVr0fBQqZU/m6uPPWWxP6cY8Yvvx6LOMtzx5VVzsWYyq56ryCrtZzEB9eu
h8Zc+FrOTFYv0mQz7ve22H3y20oJ/e+ZtVDc4pJaHJgiAjqopVb8iF0mmRz6
pFvpl300wLHdZwQiLr7YNCiWjkx5BSrcNR0aNDexEZOKhl58vorDPPIX0pTa
sDEEcFhr6ADNmL/7pzi2/DrDy0YKQ3b81YTsMGAXasFwT1QSRY6206sn0Mke
NefOP7vVqig9kz0pykE/IA1O6UE1Kg37weSTZ9PxiUsK769IMqWYKfbr2VDn
Piz3yCZrwEYdtxhr88J0V5Kc91MVQmBb9zEMhhg/ofRWS97S6ELZFuUijKTA
cy3BtLB8STzB9KpHX3OKjH0mOb0LEq/2EQDaDAZ17b2c8c6jSOn4arhL/d1T
nCE+Dnu441Zfq6ecITTqdcnsqSfP2OivrfuJGKgcEohVkdP2qElHDZvT6a4a
k+XYrfH03yDb5E2YY+ssFopOLOeHxDPSK5NkL+5+/IxlTXskrXTEV/QyuqBB
pjuc6R/aVN0s2OcuOoylf3lHilDV7eao361ewFCf6UHq0/7u0mb2RztAi7iC
sDOyOLvIwd0OXtKOerdVpjwsAu9G+EqIukWfXgM7XrpiOEaxvssAu6tkAkrb
mOoDTU59mthiuhdsuJHkV5rC3Y3ZPhiznGtyUxWi8sujqAV/WfvicC1VpgdA
G1GeF+NcZXDuXduv5PjnrdYhuWWTvYxybTQIM49Ec2MvsxmDkysBP7FQ2exF
aOzQHkEPCmTU8O8wG7DPxNzf6PAVFM/ApwSJac+pHtDXRc4M4h68zmcXgzul
ThBBfqQg3TbnrfWw4mVRvFDgFQa+neo5XIA/y+L1lIzmAdWleLHNqQrRBrjy
6OXm7N4hnR2ZHELtWhaxdyv+3rkTGVeOVePxDYocmtv/9AMjqpgtVyfzbCcO
Sri9esspk+aI4yKkCJOXukgvn6v6RxRnbxTqozYLfMOsPQlNhoxltzk7xEEZ
UMPHJ3f2VA5N4+mp0N9YtwbgBCPV0Dksj4HUU6JUuEGiULV1ukq+hfXgnfhu
iFApVJPJA10ulENcuvxWtTT/JdCn2oI4ZeTX8yvBqYAs7hjtOr5fWmxitUp9
MaNyQAOUZl2hOySqFBPE+ZLxPgzuuhRwOUmpIeljIID+DjGPb2Q+6QukTpMb
+LlxcYI8amJunukTa0u6LmzCACLRokVgL5QHm4NYp3s4ox7y7c9Ge5Tp6Mrt
eS1PIxvf0vTkrcPj90MAIFgljc2mczTZ6MvNcfh9ENcXNEMlNRRk7veO0OhR
5UAa/FwaydjRdpbfsZLzfApgEDP/6PJ7yZHM4ztHLla3ZQURauztFU5frs8L
LCgDlfqtSQSy1A3ykiTmdERS+LhKaAl6zuvPnV+jG29GRc7PPcge4W1OB6qG
4dTXMVyfLqjw4gby0cUXnEs0DE4MVJyXpo3I2kkvHIvkLa8O79t7XTRm/vM3
PRl+4xZCTYGflFBRKPjFCV2EUPRS31MlX9vkdgLQ7VtK+NAQF8CgPcq0Jir/
LWLnhvfb6BHXSZqphQjzd3vi8Gf4g1k3cRj8ynGM+rllyu0ydMbGELTb/Acp
+tOtxWZzloZ3u+BfsQ1OnyrxqUPJ5wjdsxLn5t8JvCXqJLuhfi6tDGYoKuhQ
8jaHe3LgykydH0lnv91Ru+cCuqQ3z6CAdAt2HLv+dPVWgYtYxpTvYlsjmyXM
LeJscikfpWCq0BmHvj2+SaCkEhqL4iLWbqDNQBaVVwU4mmTfKVBQsqiN/6sW
fq5pDYLJNqJXEbjksucUIKcfBOSjWDNPdZ5Xndyz5fMcEhv6suHBTKF+bAcG
tGZPqyhIJdkgZkJbcOnVc7+OxDdeS66He8zlnA/42potQDE4QUliJzciMcdz
3sKWTuaESKZEGMp+75Dl8boF/FwADYloE7M1sCydUZfbfCRTpJUIDlHRQupE
hCnUDPpPr4yqdGWpLGjCyGi5zTjFKpbUi/VgkwTW+kLboQJQkYUGIsnPz962
pPBflc79Bdj+KokrLk11WjOMTKEuXpCMDQFkikSmZEiDQLHRgHmwlZy+XHb0
b4QAlUc17FU+wO8/0XNhyUUfUVROHgXSMGU2Mjuz+lu46FDKufFeSJtgf3C9
4RsTvS/33YDHFp0ubjuwtwcYcR6jhSFDzJYBQE0EDkjHX+tFipcZIUm9oD0F
CMomsSOW/mNN4IcpVbYfz71p8UytoWGp4xB8hxiqbRj4yUW9qwP3oHurCuNK
5fYSPWnu8uJa2/5/ppfocS2kajiDfQ6RYKypea/DvO/jkw7v+Nq3My01htsd
GJFffTffbxtedNjFvSBqzCTvzUcrhKH0ozxi6WPJN/vLMylNqABx7q2otbxN
54X4IK8T5TrxkMNnFFxZ6rEAff8u4rZED0GcbNrh+bDR21l9IJrlmcDRmThT
rgrfj69Bgrd/b8nc/e7VeIcU2AIOs9lQ/5L313KzWxNWKyOjdsqQWOJTUOOz
LpPZ2A5CerjmJYxq3TuDNvNbhtuxTntOh/gzSIRsy/jaoRNgl9RLFhOn20PW
ySRN3MiKYCUJR9eA3OK2o4HV88pLmF1hkncoCOnXzjKRMPwFyTO2Sb9kM1Dt
Tkm5QRC2UJ9+4boLigBK1jPpJhtu8HrQB2Xa00SpTQat64BAz0JfmtX+l02C
TQ9S15O2kO7Ykv6flETcSJiBcx+vSkBM4JWjHap0N397QCaYH7rBm21VuMSB
lXDl6b0dy+4Z79LEAkDY7kqihhppGyR94OsvmXYPOE2FMlajpHlhj9W41KqS
YdwxZf8Iy9ZB+JyPizCH98K9EOfoc+KwU5eBVDLYc5zs0nN25rrPNL+EZiD0
K2kEwyUP/Ncw8XqcNuVgMycH+cwNKJL3abp5pI9mrWQEgaWS6+GgIb+HjpH8
+gHKvAiokmoUZnkAGME83OCS4tk5VN5jk6IXmdkhaNEARrzJeQXh/l5dKbzk
AsGBxozFz+wctS1QZo+lws46kYwZB+Ou+pIBqJtrC5Olw8xoyC009mpHvew3
wpKr8iImJEbWPvz5OMD6R+ypCn2Sb5MOw7UVtdPNJM9NA78veMG02GY2Lg6J
fi5IqrFt7kf9+m1nDOMA7D3ujcaDvQeXsHjpTuSF3LKWlCcIZEfSYw2bWeiZ
LP7bFpDq8zqcScJL2QxLIKGB6BJVslH3xA/M/MpYCr2Rbjfzf2ecXwdV59ve
9ae3JMknaVxU+3yVSu9Jws+BLMmXfSD1rbCRXb2HXANCFAa0UboNhRjLcfqb
SSty7CsanKtq8q/yV0O9qRknlOixvycumlAQSWweDkOfnm/qULs0ozjRPrnx
oCCVeGnHKte5YRWssFQbYeDjsKxstj+qvb+6idMn6Qc1IUgLat7BxErrx5ZI
ZWMt3wj7MtR1PH4xm9O80vHOYQMiBybz2N7HB9nkF99pAvOb7xqrkZeMo5tP
tiZXfBMJ5PgZs8Eh8FJfCf8An45P+2M6qd75da+Ttakh7iYBT7uwtgnb2cMN
4Ejh8QNfKJmftaOJInp17GlxPBRGaIXhnRpyLScbrUjpMOBOLG/FLRIqpz8+
M7b+nA6G5r3c6SLyoS/Trs9qf9FtudC1vf8YYTbevOfzOPL74uFYWqDM6kDt
N6g4yc2zfhso4mB3EIRixdBmexGjinX7arv5yiJd/mNZOSn5cldKABxw4SFP
5sd4yLhMyw/z+vHP8m7Qcq3fqjaA4vjXE7b6Dzrn22Ue7/CdN/pk2sPWEreA
a31HI5pFWHa2646385k1cYIda97vqjU1goW+LPfl7hzZN+aqVGXw7EqWruqT
p8/c4ro/Hp9nMKNE2p9yucjxSLH7B4Ivw9XEsFwyXZe/xD/euDUTmznTujyu
2QBkNb34ODMclGoiEhceHgdNYamm0cIZvkmsEb9Bnpa+EdRB5PeuhGU8hT7q
5aKpGuN+UZ/Pe6UVPV5qevaPPqu56t4qRbc+FzSP0F4IRounzE8oGtIWo9Qa
NnQNA1sbSSaQRIxqaMM2DCHKEYv/lGU/eQr81XovQhS0Nx1hycYysfLRpl27
B4zCl6y5idq8Pu3hn3JTHxuRtPIhVa8kH7NntdFHrPXPrhizh5HeywMSH2cg
30bt5N6gvpBZpT0nEt8/qmPpjT6OMypyBomaaB0jGtGk7K6shLNrZzzRXgUS
1DVBCHkeZX700lFACfp4mX3o6PnmaemMT07mmXfh7xcst25F7vnGpeEetaf6
edB9oxMXetTAEf3JeiQTT23aIOyVvItIAjslKfbiiQ/KPx0/X92IiASa34jZ
sRQIj2olH9cnJebbEQGAwE4ERwkOh7rTkWOvJ+FYl66860NVG+Lke0vNp8g/
1klU+khMEtr3gTZiGbuC//3WiF0ldn26DCrB2wmQ1EF0JI1kqlxoCZ0nydt3
Ghij2C5y/3umbCQwc9rqcsNdYHRqKhbOLqlDWs9N7H5R7ecl9exLgFxjejeu
2UYwSGFOEXsk2z5oUYSsLwXM6iWCb46rKLTPyb4raiIPydPmiYVsnJEWuXum
dIJpS+TOZ57CROxn3JuPoHisG5SvNVE8iQxFFsWrN9UN7VOSGkIeDNsI+l/W
B1bJIWwbPAgoLxmaw/bzzt1cXhzz2+lnj8j+QX2VWiT8SyKPbSq1Mh9/JDCs
AT7DXcA8gzQpebjBiQ9Cw/lHXot3GjUkyP8CogJhw2Dr28nl4GR94XPsEdGT
PBuIXjCG1r5nN7QnsZBpvywzuHeDaZgO2K6gje871R4UuD4oGWs6nhY5Yasj
IqtffEEQcaBD+E4eBvD9GIKyezfr0VvbdkCFX2lkmEKddCtQVZLpN3ungyZG
4+xsYvyGaQTpIESZ70tU7owUtd7VpySFI7sD/CZqHYB+pWXweyeQKuN/WBZH
IObh+/uM3xD1WBwFM1OlRDxPjBBd1i4o0fblq0NXhZzV3G4wWxg6RvfRem86
YNr7AK6jjKv8GU79kSvp1Z2mYAisJ9hR64HuFFs4/+k71egwLR9bsXKa3YM7
PMw0VQzTD3nM/kiNNFyk68JzfIw6BowtODlT63hKxeGTEcAe3Pq8WoBseUI+
G7QKJx9FDSYQbvyeMWt3Qnked0bk+Fq85oDWHanDflZXSAxx3neo4KcYV6fM
vzlK5ARmvckaIQlLNlIn504LGYC1TnEY6rjzvP03eiZ9/GdRjTGdyXNmfYr1
UymkWWr3vgw3T9fbb1X11WTGpJpaZpZwOEwgokim43B0VzkvMHAtzNIFywYB
HESZswcs9cY5i/05v6sN3QjkHlu+HVb0cOezE2YotNh0JUFZd3/YQp+GuYzR
VEDzFqtETbr8UI7cbBhS2/o3UhrXcaaLZqYg+xEB3IUckRDHs4l3cD6dS75f
BsBlCo4J4dtnlx5Lriy0tAcpK+nSSEEuOMpTgyx5V5bDtdZNaFiaYZq7BPe2
hg2FcJt/71ivVSPM9AkPmuoa6WPZ/hqMk7gD3B6is145KqxmTPeH4NdZgjIE
MoQp5XWeT6xoXNcO2i2eKIt1nGVLTuyVzjIPRq4XTAe9XaTNzNaQS9aMl3eF
2YC7GogPrANNdcyC4ZNFBexnmXYSiYMuycpCpPSq7HmRnH77rnBOT6wtFkCQ
SLLxhCCyNxyyA/JMVdGIwNv0Wc2/873mWTIJBeFsLceXj4qhM6SlopBGYKCN
lu+Xy/hLkEZAudO1TGCrCestT3n1Zd6y5hSWbqr+cnHDglw4yNsNyqN9AaVI
qD/Zc7/8AXJBVQoRzuEot4T/rmjRM+i8U1DrT+J/5znSBAe8EC+B1atuhn56
ZIkFeULjv6P2c9CiPHYdLtrydudv/zteVxCaPBNbLuWetpT0vRFSbt2LoKpj
pd/AlBf0yAuaiyzb63j9uMR9uDSkoCSku+OiQi2AfWkFPbky9TTdEi5VOJgS
xTLKIiNrG3xGQKlH6BZxWaeOy1Z8YEk6aceCquPvtHnaWtsblooitR8+W4LC
/eK3aYMIYajgBohOu+Vv9TbPb/pJY4bM9ZONAA+vh3J/joOTeuONzfAvwr6o
HfgNSri69W3F0hr7pC00TFL5ERGThZEfhfC6QEqEOeDwmPjoNPh800h/k4v5
RfSCJg4BtmCRvPhIzuxjSSoStQkQeRifxKZXpwXt1PpX9Do90E5OQH4oxuTO
oV1arZ1YmKgC1Y7W0cIp0LrZsgQPlRd3IV21HagpHsjQPkQsERcbMocrEsuX
VOvFTB30bio/v9xjpe/BX5b6xebJsKvyDnvo5N2Kyfh9Bbf8XhtDZZ49p0un
TTHo+TWWtP/8frHAkvXCct/X7vjMl8qCCH2rvNtRqdL5kVMtQLtv3E0n2MNQ
3Ur7t7FKEl1Sx6c7t8EAymejoCEmk6oUf3Xn1eZVzdQtF5FT2P5GEO4tFGuU
TA9f1cTMNX4mTwFPMA/8332cc7BipAR1Gce9vlKyQ3A8mGaaI4eeVGBTKYLx
yxjp3bz+02lzS5BAqRH60R0KICIYC8vFE+gJmHjXwhP8gZMnBHPpxojk8Rqk
F2USBhV6lMzksh7GmWpYAKKLENZe4/ztI6/p6cUURZIbT5PwfbT5HsrFqqdl
Q8jE99gS4I5qE9PY7BXo2Dt7kScPsH6+nO756MnJ/OtyyjgCkFxIeaBkAiWf
lxnB1CAcojnucdrx0hwlUFDgzmsCSBsQtDvJQweiNuvQo/9oZbKZVEmDDP0K
lQA2uuAWTdvkm6GphV5qYqZvyKuRWLKdDABbkVSjFBertINs38qQh6puvjhn
vsMMu9aDfdymi3ESZ+qs17JwlpMVWrbnmHwvssXW26F4e/e8a2FbbP9zFL/k
jPCCUZ1U6eb/8ss0B7Wo5QUGhX/XQkj5bS8LS2r5y+3VlWltlEq+wACSzbBq
mGJXWCDlgng/eZd60oSC37F021MbRqae8eRCYjw9yKuPEzuU4YbLZGmRzhmr
hjoqoFsv1g3Gn87JOIl/hnAcfcVk08D11efKSoWgmexEWSXVIZnaVDvQj03b
r+4ob4G6eJowIuaf1HVxPgDDQZ1UhzRbkyNXHKlTyfK87nAiZ5EeUH/gJzDY
VL/0fvbrMlvZb5VM7sWxAgyR4D9HE3Dm+iGWv8Fq56TaY/XLMCzdA0vrIYCh
p5p6ZGngdQmltMSYGnwB2z2ZshQQC32oWSXpa3E6CjMBfhocUE9tCfVlEU0X
ZnbqOFcte+Koujv2PIIB+ncw0lMZD/GmZ7bWzhBI7iRLWxiO58/Dm+8w0/QE
QKy5yBV9Em038Asa79I7Lyv6MaSJRJ86I8f3gZy2iQTxbu2uVs+5uiNrctuG
D6plVZctcFY3uUBB44EprVEeQtKv+Dpsjdxwb5lIf7nvH7xcpeSjGUOX7Bm9
HfhYF52m6WtPY+U2+EYg0ANqfSSXS5oRJ7yaYPNCX21EtRvQctSru4WQYg76
18txMr6aJqsn0Ezcquk/5IrCkZiu2zzcNj4l3XLcLF6uyNXOxBEKhuzH3GdO
pBjvLxZncloMXdhGuN1qlN2fZnawFjJ+c+yfmvHOZoAndV212WRI2GmKk9Hm
rCdPOt0unt5tEJ1A+NYjmHDc0kNSjiTtBv95W6mMAsxQjTvRAcV77QxbSSFX
vXl96g3Y7YgfDjwQRbkra2fBqZdl830llvMNwd7xP/zSb+w0oIj4A+m8zNVq
uUdipZmgr8kRm0ld+8DRGF9xTG/YGfDr2MvQn7DcjM/ENMaR1mZHU+4nGmAN
1ndP/fo44dysB3m3/86uEyWqe6PBMKsc0XguCaHYvuueWOT3WFTbqCMWiMwt
MTstRyhv5m3ua70df8FYAn+WzNLB3F47z3Dbrr++IFJKiciFnsm4iq3hwwnC
3UI1NzI5EnGP9HwPCvI7reHJKb9kkDZIq8G+rITS0oKw0P/KXG/A64glpXiX
J7Dl/o93zieeQK1EXoxyDr5KqGvPKdTzudumaDZxG9tW0sNJz/sBpYMwZpVp
wcaHe6GAMPmWCFynuEPZOPIUB1dWWvW2mu35+z8YTdSh1e7Ij1l2bJuTuvm1
Enr1Rv24zFYXo6GvHEHXF1Ffb5p8GCJXry9Ozh45R4uZMsr2tNBKzjFMyvft
X4UbVtOz49Ey71PUecLf1r5VBXDrqyCVa+f1y8ppEW/QyPyUdUpIDY2mawEj
/uybIf03Lfc2DPY1KmAXzPEfW/TiHV+NI1MSsudva7IjfsIBcmZ8QVTgqVoU
C8okwnWh8uM+ufOZxgaNJ726MPznyeIyS1BuV2P/FRTAFhbMHzffM4Kv0Bxf
Am24AcBIr6ac7y0xC3jHFGatpuIEFUfduzgiGnj4ucUT1/oSZW0WN4xEV3aw
s2zcbPBkHvGjnr64jf9HFuKicD+zottGCMDJ4hx6qn4R1BIvt8gXuNMjWajM
RwBT/O1TSCZBjT3A9d7BMZMecvnWyLdGAb3qeCRsSGooCvJMppm2B2U9OSCE
4TTaf7a/8uEOTpZDbniZ0kRtonVS/tHCPgIX4PdM96FpAn6o8+8UVwhGEfhQ
Xmcax5NSDuG/ZX9W66+ZhqHQRrVOWH4wTk18/OZyaELkscoW4fRMDe3mlZJ9
ri1UDoYA3K2YX2e5Hxu00UC7ZRa2NqeKcquEEBcMPLo/OT9833h0L9VApQ5P
IyYCA2E1TTvgyMUiNLWMG/cTwuH+4V9t/A0EPMPOSAlV2B6GnA7uIXk6bbFv
kl6EGCkDJntnKzVHlLsdzsulMYcvunwjTA7WXyaSFqYh86QkdgyZ3FUmtkXF
1QvWmGQ7590Pj0kx2xAWtguNQW9jnX9cxt+ejbVwLxZAHVBqtY88q+t+QvVi
JOwW02SdY1WGZv8QOcVuFfbhGoB8yWCFJQ6ZiNYlBwU8W3O12YSB1gwwN+jM
xMuLQxAgC415JkQWsxcf4dak1oYzf0vCEP818wMBlDPwsTRzwAk37n9CVDzA
qLF04XShcMM0giCViX60YiKX1OXD2uIiZrbtYgWyQtHRC861Pu4gJ/oslYR5
VA59yS15qLIZYvkt/tQ0KxYMB6QsGMnMQUewMuKf8BIcqRXS2EzM0gRx/l+u
UzXOmX2Zzr0WzSzwcrhpv/SoODBP2CvXuYi17AHFcq2nHHLoOYGH9Zx6LhZn
T68X+MYmanPwJesiwL2/rPWETH1nUPdzFjScbgkgxL72y/U+CNC7v4uj/8IW
l09hPJkS1B8B55sVgVxyFSPN26N+e8DC9wtTh5wMq/SW3u5SHBzSfAWDywRv
n6FAj+YGv6lyrzOjq96QTA5cuqa/SHGVeFU9p1K2v8jf6yXL/7aYCNXfjwX7
My+J9589Z5hwyQizzQIGZX8DCVHAXpuhjvF2dQhIUMFa6hczKz4gSk38AWyf
ilqMFLY2SkUDfPFXe1v1mrT7/iDk/jo5IGSuWe30LTi8c+/ji9OM8sGlqiAP
NLDICJOYQ/bur7znLONGPE+pTGogg8dLe+zVSDzYMuC2lEcBHSpvSRU14KFU
L6wlei4+TtoCnf2A5b4drGU0lzHTg9WGtwxRQ3GnjXJF05M+NM2PDeR/azWJ
AGbYYKpz2m1Afw9JmM3Vtin/8Q4eIEz8Aowjfpf6+ZqR+TTFO8n/VMw1Wa/p
zor6rNNY50/aaOVTePDoCHjSgHu8eBfpU8gipaXwC1W9wE2W/tQMlj3zjeEA
AocIBjb70+h4i6waLivUGkegtM8DiPYln1Uq81UhO+ET6lceYFfzNVMjLFpQ
DgRTFpc9vjDLJ9Cu0uaRV5JRtFpO9hH7AbS6T3pejhF2gTc4SRzghoTXguok
jdVuPwu8j2XCKC8nFigQgt+BQMfdDKOnzyOw8M6AdRPQIscv8sBr4xXdu8qC
U7PN1hzWIXLBC1wPtIolnpU8jIIi8eXs7hmk887P3v5ybzHXQLI+LovGS4Hs
0tM7CoaATQNiS01qrPmHjghsOtRDPM9mPok3n0luQAzlTO6QpXZXBkakbTtM
eYiPHuCyVkqEcc+0wmqzDuZ4YjH3zcNZ9hek7HBe+z9PbLTw59KtyTAGo0Zp
C0XndXkXrLUBpu2K6jJekO6hNbO7JUXvf0VXy5BNCrkGZZOBUrPrsozEf2IF
YtM1/gqUWGnuTNvn4kjxai+qjQ9yVwfmpisR48GPUtA4hqeNJCmjUHP9vDQx
cWFzraddzOSxRQI0tb7vwwTLpV6/WyvihRpnvARKwiFBzPzqfTlMX/PJ3uiD
M+Hn/yPQ/V8LdpHYaJ/ohSbtXEDXZnt5VIsjdxK4iKQvHWoVcklGBS+FuT6V
avg8gIrssvSJ79CdeW/qdf/R+ROzpF+y/8dB+q/effy7RonbTpmjtP8OUrrf
9wE9/pbiPiU62r0OsPsp+Oo/v/KBArsgRJxM/IXmtP23APXO2AY2LIiuQ/Ph
ZuO2wCpkrDoMmtvVGDHRZxSOSrp10xCK51sv5xYr3j3Qnc22evWch/qGFUmb
vZyG1V/q3hnfVCPSOKV77zOK5YDllYeOSXafegMNLdvnpGI1IaHc4E/qSrsX
i7kDTjl18U7R1h8LbDUIT2r2/fRF61Fk5QaetjVOXLGwryTMxwY0nSVCXkC+
ABlXIhmAjOJ3VzYnQy4fCWeWWL+ZYFA98RaXsrUEd5aaHSe7LEm0RkcoSgfM
R/EmQVoFtDDxU3HYeWCzt0+yZb65l4t6pzFKDDd5SNllyWuqZQFaR3f4vb09
/eYpeGAvGSiqU8qkigTTk7lcIjruXsjj3FujbElOnCefH1SEEVn3Dck0cnJv
tILbeN50qtWDBzqmljxXbH5ufXAJJtetLDp2LpB6JQJ50C/9aiwgQgSe+B+H
0dFa2XQtVLqnM5eYy+yjLMkKNjd/XQLICGc+jMWoTTok/nrWlTS4U0AFp1tQ
4GSOy9a5k2lltJcz01xUu9PYR8LyNqmK9pF9L7ctwM007Sg5LQyhhc5S60Ce
Y1t88Ict/I2iY0AX1SBVzvAygNF8JyseTyT5aPcW3s+ZMdMM7ngxVGo4aVew
ZEaX80Ty6rEbKD7CP1Y2sKg8KxKhiaLuJiUZIRxLzPGcGVrqQesVQ3CDAQ2B
F10oPYLkxUwqfF9Awhhf7P/jWcJDbENffOY6bplAz4GYiFQVNrHsgad+lLN0
elrihOQ8fkx7vAedKADaGg10MZ13R8dktBT1T4DD446LBFjQwGM+OXvekUgZ
ZFMwa2H+ZGiKZ79zr0lDrbc4+YGQvspqGTc5Tcg5llyzNyJAcSV+5pp3swoM
Wrj3UaLSMnkCc2/95MsqnhIl6V5dDgEMu7yR8Y+PW1KfAVkh1bg3xBX2EF0h
8ki5NO9FizUqkGvOC/t27845IgIHGPrcVy5lGqQ8odAABk4Ay85Ye/wxUOsm
3GHRb85wuxXnSs2fx7RNFPRB+LH3dnHUSHDhFbvnwLM5Kw16CzGKEFXIRjNB
bAgy5iDQVAXjCu/UA//OMc/EvdbLkDBqZazd62odU+ic2E2JE5FSJwj+AVBn
ITHgFdrxSHaVoToxsJ3yHmiJTRz0U0wPeGUb51Y4Ie0MDbL5XLNWIZmqfjks
qv+g0w8pFxkqAmWlHjT9VdtcTpF9cjohynrnY8HbaeqhT/Lr5AJaUxjIsTC6
97OGDWrOgArBgo17FriWeR02YyetZW9DlQUnOUwzkjHxMU+18qkiNWQGLFzc
ob253+Bd2Ry9WNr47ErYDjxblgBTSdXszMCSVMtLGf2yAqKvEcEBD+k9YQMh
GZ5rYcMdInNl0wm0Lis0W/wl5mFJDQhaSt60hpaB01Xj47YjYcG4KaIs9deH
qaS/8ULx/XIwszsupga1OymMrtxyF3oFwUkBDmw/+Q7iLeaUxtOiCRFtlyPb
aPrNjOiXte/qjt5Ol2oYPo2MBsIbighthzjeNenFLgTE2X9kk/3LrAuuYjsZ
z2/fznDae7EKZH6IntfC7OkzSEhap7KFQvUmuCyrh3NwfpvtUDEecSkjxdkX
hueRd0jZi1au3TMSQyw0onqmDQ1fcqXGnr0cCxTnMh4VUbkCEq50vo33xJea
8qea5F5j7WAdK+mMMrXGnaBfYSarTNnw9/8pRbulvSxBmaWIAPQnuu+JztEI
OFo4/WahrAeFppIr3zOJcKahV/pmZa0JU4HYk3LL/81SCapMOAJRNcpMYEBN
TPElKEWkizMlz8OxPTxg78uKWAwP0fJLv/PmMy1gRKsdEAtnu8eiH3LBl84c
+j2kdeXaJ9aoAX10wRglt+4mnUli9Rjq6XqrTQlfgplHFmlRG89QZwEBwHzo
wiqKCbunn+ahQymUYOopDR6G9VD+PAlKvQCGlBjthkhZMbSnRJrH56ZvUHTq
d+MpQgrTIyGipddVy6UcshM4jcQ1FXOVuiDeA6Ug7yB60RjahU3k8looG/VS
PKHV21Tk9+majr/gnS/xg67DnIKfrzt9q6wak+vFeUpe35KustIBEvZF+orR
tAYVEFsbgn3XtNyc9mLn1RP2lctNKbyhLyjqXznvfayB3QrIKZnQTg2HcbDv
lKJm8DlLWRSTN4gTpvFy+kQ13ZZtVrbh+zAvT1YPRfH2nu4XHJ75Bnpr7peo
BTpT29bjsZYK9GQ1LKkywmh5K2oaV2iUV8VnimydXf1UlkXUdOhnatLtIDu3
R+ASNbV11BdEHyPvwr8iZUg2gwTfFagYcd1oQpgqsxM2M/jwNK4hIprgrM0s
pcf5DYjYDV40dIyCf7nh7L8PhbcBCMv0krQbV4olWZd+JzPkGx+tktmHVDAf
yTYUfFJozsm5yaY8ZKtcHmWPIf6C3KsxduJBVwDsnIFJ7bUEq6c97Kp5h6BG
neWS6TEzOxxni1czx9RN+4JUesOgR6Cixb//llh5D3PNyb0lRR0lCSoTc/dx
3R0smts4bsbHDaupwvXPHF6Jsxv6enBCWV6l9fxRV6UOPMn3XW6nubYcqqmb
B2CT3Op8zuTXSsHopUBl3omqCC6U/Out8aWyzsKjHn+94q5PU3XT3TD3S/zl
qgI2QpAwUUf9HtLF2dfqOmFMBHoVcP3cmt3f5CvbU3BemQUEAAV/nCXqxm2o
3wXrAEvcfTaXJycbB1SBcT22k9MtLMk7MfFn2uNtR3aV4S/UN4VWGvoemKSr
6m4xvTLcQKaKpmMckVbNorxryIUXwHKGigrAvBOqiOQyhjAMFTX2jqewv6xo
sD8EPvXrUkoZ3+CnuJNBYIs2fmjYpcPZl+gzO8QfUeZbfzhN3BRq1Ou+ptmf
mNYZ1tbR1UCjY9JY6YRFyiFI3HFmYVMkw8dEW79AmBho9CRyKh4vvoRySTN2
AaqPX//duFmsGkSJucoV5MifP+w7Bqn5Sp41MLgRwLwIrLNv1vEIP8jvbgQJ
IBRpBl4Bcnvv7hQJIxUJHQeYH/d4PYsTMusMbQafKd99zBQ0uxULhZIak/PU
v6TZ4Q9dWKouVr4fJX2OIJZIKmx8+mRxoQG5+VdTGzgbTFx4NTpZD6Ym4kGH
N5yxKuMA7cR2QU3i14uZudZtMNVHXj02wSukd0xaIHtGy+1d4ybrI0sLMRRu
bNu7A4Nwhh2zVwYmBkt7PxvbYJjNyZZLdPSIBA9RbcrDn3808+sDOC3ndjtE
IQtyfTgNw+Z21BdSQYrWqpu7q5F9tnDgiCh4cFgubkcK3uKTizW/EQDfwJ0u
qRgAk1HMrjS1Lg340Qs5q33kr+tSyhw0NjVTKDkY56MXzfgtV3OXYj4/JbxX
puVAq9yjyB788DbJ55OfbPgIhK2VBz0cSUuTQckUZRHT32FtUjXkbIeiOWjY
/BW7oHRAZFogx1g0Q2mJMieO8LfG6oqH7rhV55we2A7bHAj7nCtZYFad6mhM
NVnp2Xd9ni4lBWGDZTrHW7xYhagUUqyq3BGwtA2cJxDSzMT+hQZBoud3eTKg
JoCZhVfkL6dIawtMspiP/b/jYfaSpJ+euihc0LfGVN1hVInaxkvXeX3Bo1P/
jI24uS+vLDXmX+eXK0hNb+c18X+mepFh8ncO5pl4JlojB6LeYoW3urzsrnNg
lyNpVqP6Hn33YdYo3K/to7bl0rPnnSc7ZYXOFRAuH6PdYBdXMpBp0TPkRQcJ
rlfCXxh/WXMC7rPpHjeyaHJQcr5F/FzpgUe5CNw3gcyYTW+GdmDrN30F4Aor
Y4q0GG8OqkSVImoobFqRgYPQXKuhdFz/XoFXMuodx+GiopPEhhGelBJCMBgy
VQIs5dd+unoslDUMbY2mhageNcBZ1UEhUSuAXHq9YSvMmsT6SvCU4YkHoEs7
GMPmktRKvNY5oT0XKFMZIXkd8tLrtl8pm6SVmuD6my2ZKHitedvkIB2Rb6jx
uvsLwVUB8lIlgdFgEHSD9twm2drPlySRu80k5bLlxu3mcYtP0oGPMPw5LZOj
CsQgJN+eSnqIEpDi/PuREEzjBNGVmDAYlA6MsppCIfZ25KBQ1XTUKV1KF/lq
dPjiVCwQSmvXJizLOkdIveqzgHqyDq5u5D9npYdD0dcj9WMqAbfIPEGNiEQn
xzkM6NuKOuvFsOwZtcW1IwCdOdQCwoXtc0Uu2fjHA8vVyhd3Jp11bd7MA9VX
1gfS6jFxzyO09PitI7MLg4rwOiqZgSSHhG84VByrQZiol0PEp+/JMwfll+Yt
ITz8oxtGGp+cLooG0lRh7bWVUzfESVlvZyyjgVL4cgoYmJM7IMuLWmuj8OlP
LWasa6PuG3z8LNs26xpZB5wZGL4adZIhXqbJiMK91fYnfuhkL+KpT05KOfmS
IrF9cJa0/5wSip0hxFe+DpVpecukMDzDre9RhE9CqvS42G2b/zhc53ys4Dou
F7zOeXPpdNj2BpIv3qyWRtnPDg4Qau2iy7rmOOrYq8nLilBZPvsXwbrJU/Rx
AdHDtId8o/IzMV09/rOwunCoQMiPtvu1t06ggPw/ISkvXzHuyHNmSSzpKtyi
9E9StbcgbPePSL2AU5omKS5CoC/GJH4Ji9vVUCGD6WgGZWwnGDuluQmlmwy3
KzyfVp4xT3zqCY8OxqIGE+jj+9RBNqRQFX7U/EexmyJXjyJ+vlwKw31ddgj3
WWsub/AQ39T0dvicJ1BZgAZ4SHZiai6RPOeCfCJTFhWMH6wkGvl/jSp1ZKly
S00W+HfnzRFPbvPqk6eMuRiMozhOd1+RPFJpkQLHg9BOlDPfHK1tkKVdxSO6
Epek45y+1Xr2un4CotTZuzpYEIvZipxkFihdjnkKE/KOGmJ7hnL6hD3N6b9U
TltGLAdk/mcS3wrNUbN4hoSUYdBH0IPyPxbiRyHJBkhBuUPCEdOhTZl9cS6W
4BhXTMR89H4FCmOZTvMEwWLmx+G3V1kXJuC7rdZJpotqMkXn2DRTfdoeGS2E
f9wCxHJ/JNslqeQulICgnhf/EK8LdlEcNzHz6FtaLiK8VnGg5UxHf8AdsZ+8
kuz4JuA4LehJdKtJGibL+SUWDZ0TOM2t/ZGTk+9nKK9HnwdPUplqFZFR5aHe
r7Aq0DLjG9+alzrvY2jDYB8biZgQSlHudx6RK4yQDm7mRlriabv1KK8SfzU2
eqxee3ZMJXP6v+Mikcq8cTA+/PX9SePV4HztyXoupcYm8lyjjyra4GjyZ37P
htomnMuVd2909y4DCEMFfygu27JOPld9NalS/4+asGvEM5HjTWZN3M9U6kZ0
W4Yia/fUpkWl/MM7fERXbVdWUC7q5imM4NjHJ8xWWoLRj/t+hPgd+ZRXcRun
v44/4KKAZ0rSUcWoO851baaJS534LNar2+5NsZThXb612ymirbup/O+uhq1t
BptJBGRIaefaBv9PVkAqmhxScOAT/GondTru5oSzfU1SzfneG59YtOZ5IDvG
BRXyz9OHx4lflrREYTOGMPQw5PvP3a6f3rMXk7Ba71rbdUlpekhmj3hPQYwX
NwUtYEKutvItC6pWPM7tE+nMm+uEG2hgX3ZOv2dVsRx9qAl6fwgdxEn5XwsD
/1b3EdJVRxepUbLllduXeoox5SWMJVzeWIORTSB/hbzCGJOPGdaA/zeLFLb7
dWXQXl9qnQwpGesJ/AgWgkLIF+B7+HyV9AbtlyzKJHNMIJ3BjPKjhExYf9tW
vcujefiIz5J+HaVTNhoCrvnbvneBzPNW8N4QSsx1sfbLH3OaVpUidw8qlTOH
eDhfJ6rm6xvRwuRZ3YiyAUDA+F4SHIQQdNzd3H4/hCrSAldzlsJ/2zB6KwEa
WXjY3JB4713VyM3Km95gLZWI3WdsWsCYZ+qJLGe3PlQ8izcmw9H1Co8hj5d7
lylOSyW9iQzrCaapgWYphgvfTNIpZGiuJSk+OlOnUEkCHg9B5V7yC/5vkpX2
eDDOK4eVW+636nUFUoC8Zit6riPlhbqD/qWerPYujNle3hEvFzODBlIww+fv
QkxKcjPxFsIwV5rpaoDIIZl9ZPNkuJNQYNVDCsnDcx3PCYmvv7MqM5JbXJsX
d+jIhLn823OjQVF3JsdhkmdFHX2AUO4yrn/MfGnM1yqrHMH9t5wh5WOGRcMn
1OwcjSQJshFFUwhTzdFDIVtJV+nzRHYtuLF2SJPEDsKVUMIb1RQ7/mJIdsou
UarWJdLN13SK+eNWj9KKxRPQGfB6o3YKzync737/pPtVV9EUjS+IhKpWsCqv
6ZHJO5ojyYw++w/sL6kbQlXs7bauK9FFYQFvQukpJ8NUC5M2p+k4gebSmnBv
FGtMfCQGlS+cABPK/jkX4jOWU6QpwSBLqMbfCkBhSGqgpySBL3+ac6TbAY0U
SHSaGmB9r1Fj+SLPoEt8FCEBp/zM+UHPi7hisWIifGHPhfxawa5HflU37VZe
WaXnAFFXaL96QS2WCrb0csqUBsJ97QCNngh0As4+eJcHxizFlbuPgesYLwxT
wQIa1+xwDDEpuXypyusBTux8iRHfN7+ptO4REdCHmeStvpTIg4uSHba5lD50
2ZVmpA4qucIG+/RFINfenBV0GDAqcBytBojTHxvV8cRwhWIwaI5pcBhhUuWt
PpUj4UAfIf5Yb9iCbsyVdi2gl1ISik7erT9xfQXu90mSimJUulSdAsuSt0ZV
Oq4ZqWtg0802JZ4hnS5EH5fd8rfCNp9OIfFelw8DCXOcUTl4EU2LyKny6q7m
lDlhURRFqxM8B35tHNkb9fMnehUoOu32CEEmBC/pMNe6xiu9cpVZJlyt5I1K
O+a9VYMzd8rSvsmtAaFVK7p2gNIvYveUiSzii39jVRYbisjge0ZAV2L/1ipy
zKvvZwKZU+wbe3mhFZRVhi4yleGomyu2Waj/xzpVhGpgXOh/1hljJDpgjfzm
LX+xYh8n7hTGS1A9qIgJWRuF4FAHg0lP630B9PjFQ9B5E1SrbO9rbY38844E
xeezX62sIrOiYnuCCVVqPQQPMPf3lHpnZgov2bhVct6lZvOhvXSmVhuN5RHe
InBnoYWvkJoBL+p36UKM+6Lwc3B2g1Bbi0yau2FRFkRQSuaGzLNl6dWu397S
udWa1r9yt0iwOcwabtc646CpWbqJ0tTOrvLf5Qf/GVeDGo1iLl2JBjZzGI7Z
f42dco+coM5f5nO5jGT5SqKKoAF0GoPYx0GJiXBNEH7dUIN2gibexD2y2/dE
c6fEPxZV4oAlG4G7MPM+kZtN7ULgo/e6CBdBbLLItbRYCp3ngnmhfK7j65fa
gPomZfe9ST/4W+T1ngMnSeMTIjEO2pUrv3/Y9r38uP4wPhW1lwFpiDKF3wH7
jOkjvcvoU8uCAzg/Lz33qt7NorCpvSZEczudThTU2C1+1Ej6r0iAen/Ccv5m
G19YQaTmIcL8kuYPbHAEpPQpHUNjRliOLJV251bFJ0Fbn1UoUZyCegjcvP8P
EikHXnrGvzkaMIbZP0oUptc3X0ZYmowIHCLq3lYfpLz3pcsxhut3asa3QBCN
WRtitHQurq8hNby/Amt1kg2tkk9IMLizvosQAUVk83+aufFBzmww/iQz08Ye
Fo/NkTq8SzA0ubI/X8AvIEba8NpXQinQUUjtGYsqg5mgaMT0niiUeJpYdNcQ
qQsXvVk/LQX5fS9Tp7q59C+ApFDvbl/KFowFgGzs+IqXun5z/9YX/RMVErcl
2t/7TaoKIUUYHQh+fCyFnkKAmPhPrUd/sdo2LAsgKQ4c0uiX/qZWleoqAvLH
IiAvYj8vBpv0KnEjzk6dDSbCpd5ND1xdnuGsCHO8stJGboOOLlSRXukiy2mz
ckpVWJCvpABSZfeXmfUFyuDx8ABfoXajUraSwyI6mROvN6jmstFwGTxp/aP0
N9zBL6qR8fbCsyVB0M+zJC9yceWV+9sqYZQkHhewpKhGVeIbmrOOc6GxyNzy
fVlvWbCTQTeVpvo5wIDoYhMRy1YbWZ1u02Ukcrkz0VcBCs3X96ejM6iaOhu0
04TC6M+fPn7jaWuUcD97MM7sB2B7FAfQAymjecvBZA/h6FKkBd59t3k7d736
56tXrC4P3pw4+6nLEp9SUAL2bYdfwzCyH3Dg2TAW7ABWB07k3f3aHM5jo7Y/
xn446B8edVqapysKsPrbXMt4plh5N0W8+PAM28fg10dWRLSGBjgzAm4h9459
NGhhosxiBuHj2udBzhDZhx9u3P6UbXTtTwEJMU9OlXYW1n/PHBqwgWAn/skm
xPugB2bpgxlmPQXj5C583amfJjSC/i+UEhBNfM2xqJPJ4uWKrL/283bRlrUY
F3sa8+iav46fiXS5EVYsegW54qfXUO9ZmKDa+/mfSmEiMYjCg514IsKMBYY/
CDE5/hAP+WP3BfkfI/rxcKjioffZrOlpNVGTA2MtpAplwRzYhvU9dRrxmkhf
EL6WLxF5hKUBDj7bpz0Ltxz57/g7IyKehMGFeMddKNST1IUKuXAPwwHF8wcF
QrmStBXoBoDkjtldFh3x7DENUI9ZjmIgf6W0PCX+hpSSvYRYQRsm/ndIeBsq
EHLHY0TRmSx3Mb1DYbKdq6e//k5XH5gno4g6oF5cVCFcnueyh1iCdjIMXWGp
G6Hi0SfVr38OqcSq4/kaCzENwVAKFB62U1/t7VvIMUWOCWlOox2cgEg+PDd6
x6W+rP5tIEhzxK0LgU3WoaSnEKMRuInUNmRPk9pzah1aGcWSgQpx38k/5R/S
ZRfFiRfZgWWpAkzHfIVnCZkJ6KPkvUYWHbJLGksH3BcsWG5ejsnowzSc5bVR
zTMMTfC052sdkGFu4Qm8cfDzSLw2d2hB4GJSAcUaAMlUQ/tOrnqycpNJ3klM
y4LP01rSUuPTJnuplfBFxS+ZUUz4u+/6MN9M+zJUJgO5NL1e77DwLzJorN96
hgEfTLmmn3dz4HgoX9bRe8dR110lLuSyU+oLuk7BHBFqG4koAhJLecJxiyy5
pJmg/ZDeLtsbDpfZgUP7737Pep1cHi4+yMYQgS8t1NpzPgFCBBZnGxZ1hmbb
RdcxN6TD/gq+uuAO8vfTnRUPhrL44W7RSpNxvCHNxr6j5jA+swqn3iyt7tC4
YLq5yvUR8YxbJPXYSVX451+TxyJfszuHOSPnoC0U286rHx5qbIl0qE8m4cfn
C2cqYCzBz8cUY7SYuDTHUAYWZtNIEY/O0PzX07MhxpveYYFuqj6ygENYjLdo
pEK2djptCtRhIYyLgWEiBMNpKhPKA7i0lo1DW+fm/WSN3SFo7npW7KWg8erR
JyM25LAfr/+1klXz5G3UBwy2kD0Og6M0SPe9ERfUqDvpPK3EH2yp0KOoqgCx
9vBhEbXHIL6dSxVshre/vi+GhVICDBcIncP9YnO3aP3p+Eeysb4a/F9Pqqs/
URd2641ylcF/wKveYfZ3fElNOBD4Du52AEduKiGcoCGLSip8/HfCAMoVWsgF
8KZolPi/AohgTbGX9lcWBVDqkkdL6+IwMEdEnqMOZVk4AVuj28sC9jZDPZBJ
b63t27JaQCkuEenIMXSZ1DVNDypJHErnqLoJX9y0M2v0XOVMGpEpFs5UY8EC
a7xD6UThYxCmcMT5H5z2qPGDJaoXb+2VSVGJNuJOayQ3/+LmNeO9OLKMAN39
iUbFb3oia9cqnNXB75wL0T56QuyK6DBpAdFv5g1ntPO87h/zEeoGY5e6+Jxq
u4HhzIjAexrmPhJeccWcgFSCCwjOURhD3i1/EhTc5WkoQmDogal/sjqoR5I3
d9w5XEfXQ/A6ddZ8ULwfKimeZVPjnQI032A3RBc9C1QcLEFOqRoqj6gRUB8m
CiQ2NFmtAGjdZFbyzlNKpBBWmogqvshKg9UHiVAlPkiFFiHhjFJK3dRlrQHo
gHUEJmvXtq6t0oDRughdfSlHxDBeNQm5cfnUhhX8JoRgVkatJABRxE802+cm
KbfqAlSC4OhcxnSwq2g+JOZlt3ER/D+tHpOxaoYU5n/XmTEdAazd/h2WPMoS
FBFacY5cSkkD/TtnLxqQZ3ag/vwPQ1ARgGt2GVRUvwAT2DettJZ7FLwmFWPT
7yFFtPiGNppLiTdJSbpJNLEWLjkigbRaLtVas0PqZjr6v+7iIAhygc6Q0xEf
oOsr6W1GMtRgzlnH2wQ4ZO4hGsXbnJH+0a3W7IlcXxBAt/36Oy+SiL7Pkf2z
6uvwYmUV69BjyQQlZnMbxXKmhuKL5jpV4+u5AgSmVE8PaJ5t+KM37ynD6EtF
gs8tfUQWBIZ9tWqKedXN4oSUcuGfEZb1EO+RqRo0N1R7qT8HXkUQosMckh3x
M5qdSJ4ZResVXYYsoSTdWxINykJWX93MFgVuTdaA1FwEg09W8/wubX7N51Ml
/vjLMiTsSYPTAPocIJymR+aLQNAc5SgyKwZo3XQUV8SXH15kp4b3oTi6Ip/9
aHrzzuE9Ws1cD517fNbtbNVuSeV2rYIUgzkDhm2shvBbHP9d6DoNBofam3OO
leV9eXvzQ0AM6dao4w/bxx/lU9+NOweglTGo+SbFyn4e3/LkyeTBJPFbnCuh
qwnm0TYSMgyh7083X8EmxLNQ1ZBvOaruUZwgGx00Nm2MKKN4RW2g23rA6I5X
29Ay451XVMWeb0L88yAL7BJQxy6d5SLr7gqe2b1H0y3dWXmKGa4JjBzckOOr
f62OjX1yCQe3h/OiUP9Wp3LCv+NYjvfYmj1fg+LMVS6ZJjS1EMiabqIQJux9
8+czAeV+DM0yPmr6eaoCZbV//pJRdfIoys9YW0En9Oq2QGDCHfF1sBsgmJts
kXcmRHlrmarYhNLHYhNy13KlgGSRJo3Nzzf7gNS40HSeOWt+ZG+UywmdiAod
QcY37eBpl6HbCgmg3LAJq6WEcnO1EnYQsRQK+LKl1pvxwoXzkXYqlL6HhWts
IGslj3dQxCXfbQx+SXtCueuCPcT1IN3+7fCWfrzLTNVZJc9AcrB1HisIsHru
D5P4+yaYiFuSY4opFW+82x29WiBxScxonzJG9YLHyEJXCTbIsRmcmJwGo2Dl
bUkfH0J5Mj3/wH9fgPKFcSDgHe5Q4gJ2VPBnIKhen0+ar/WPSf/2kk3oap62
8Q+jKo6fZsrl+0+OkbyIHtPE9hD7gH6xH7hgYIsqmc/+s67v62Vhg53b0c2d
dyAxtKwKp59L9XQKs7ZtqYcjbm+K3k3F8OV58ORSNQPe9khQAfFm+0RBvrBe
VhxJfuErgTHItdXqLm89gOUEIMsc4H4q8u2byzsLPaV+zQain99HtFaoSx1y
ln8EA6GxcW2f9yYiOvObbaFQqJBknkcMjWioQctInaO3Vw8JRwnqsKXGTVDY
d8g9p+r9uzIG4sHrvbSR2FImAXmxZxH4vNA9Qz9LL03M2+UbzFOScAe01ISB
j4WjKpneOYLuKu6t1XDuAmCLLefI9XsWkMriZRwJrF0ba9kQSIX4esTBu03i
R6UD2qGDVo6EpYNGRNIzEoUgfRGnIuyc5KxAD+uZfn9y8PwP+X13XJBLUFTq
tF5tkdAmRaEhDwu7ekdFyO15K0kRwYy7OvTMAcj5cdpg8wjTCAKa9TUk9o/n
fRKTs9uJN3jskpDCbjR+UkujSxETVs+AmJ6hk/A+1GJhYucc2VrW39rK3BTm
HA5ItiDCN86DPzA/CjXgjbffJBkg3ueTJsV2/iT/XjdgZRxrGmEPmpFcnvIk
K0EMzRbiVdID1xEk3DCthxJYff72j+b2F9YELfuXruK7tvmDPKBlROcAk4eU
46FPxGkGIwMTb+9rCDL8EcEf6w6++eZ6EmRVYTOvFt7/dOml5/ZdvgImJZdR
hKIOWno7MV1pMHE20jHD+x6h50PiU5XSBnmOCpKDf0SquqFjTuV79a2No/Fm
thiGuDt3iXhR5tVHkIHU31imCvCtD5ubnsn7zRX1BQt+omIKGKV43jZiQuCB
xVW604uVJQMz3YzlviuylswfRjEALvYBZDmJPLoYKGRLFfM4Rgvu7SXmgAmR
obcZx54/i7AGEidDcqIvi3Ox5T0Xct9v+CDxO52LFPhUCpO0ofT3JP91q1wq
ARmPTOxxQ+Uj/ei4idwaAUbc+DxoA8Lc24msn86uY/OKsEhQrLk+2Nkm0yPA
9+hThudEmTaI1RC0VwRFWsRWqs1tGraZHmrGnxX1PIwBhrL0CRBMExYm6Xxr
joc7VATBKypNtPFWSd4gpVoF0MjBDz4Uox7vjsbyRemun01Itqcb1kPCY5uF
EHPdmP+cNchCQLG2+vBSXDmdQmiv9cTHWw0ZzSiUQeTgOkA/LnvsKWYWDCkF
/42n9NcY/rBzBvhbi6g124+CQffNAlsj/uD9Xv+fKpwhrttnTWcfoNsu/T2t
Su6dSnAsDTYUIEwA5Kg1EPZJElds4e/5WAXMS3DetAlLDwhjiIWLXnQUObhz
vmKFZvsYetyEX9MFz89eRFJ+yqoTxKf7WShRlkyZF50Lrfwp1xgNDSpr6FqG
pMw8NSIzCbQw3dbFOCJ476zSAq3Sv4PaLNLhiZl9lzk7H8twqajbeEsI1x9U
IQHrYLZ2tTgF8NrDzO+Z9cVtpFgpaXaEHL5Rv+TWbXtGOG3yYaaDRJrhEiHJ
MAcV01B/fzvf8LaXhpEr14Kka8ptuzt9sHJIZIyEEhg+/W8iCzDlci3zOiSr
lg31V8ZcmxezHR7+NmCN/CuKH45/AzKDSv1xM/vTMajiRKXdkwCRQWDAKYcL
ZxbAY3iWkg8YOJ/Fkl7xBVbJdnMa8MgRA0/HDgWZSfHIm/FG53h02D+bzMmQ
kCMdYQ4GGbdJiE2nzgT4Az3EO/mLr6tj/78vuHRJgJSiRkBIih9h5pBSBFih
9rNVGQmYxC1EvSfodLTq6vvCq96P0G8YVvCMEiYl9vo+R0fi3fXl0MlABxuX
6iUN8uiU8R7zaLKBaZDmdmo8EYY1I008PsaTVlkLJC0H0DDoIp0tNdQeBdeD
KA30uuE9L1G9s40FoAWGl7S/24yZ7+pQd7H4VGYZyMCvIt4ylZhI5MQj1PiK
W1wmxr6XS+1UDzCXTDpzmiXhD3wOIW3EjDzFOQG5Fc9bbfoN6HyN1rChAXTb
Ro1zDZ/rhWxD/TyIKdZnRF/qz0B1Qb72RVdIyRLVWSt4za9aAF1/f3zjOV+W
9X+UYqjIeuKL1kILUHkhDiMgZl+tJGlzp0Pq2XQxA3b28i6yNxZLh07Z2DFh
8qIiMhYpAt9va6OjvacRXqynbLo5IDU2Ox5Nj6WYMu9vDXqzYzG3cOjyxEfw
wxK/1rbEkN3ogA157eZEZ4+GDVZyc+Wnz66nqyNHv3LzZGOpshpnI0KdWVCR
pcb4kM4FkfS3CbQDGQzcyXGSj6lUwWJ/mqroko8lGbS/T7ANX4CQLkl/6a06
kI6Wkdo9IMeLWkM7mWZbp7ldMpfTDiXYwTW7rjIDWDnh6ono7ba7dGIIHxvC
k6LNAGaOx3IizdiyvZAojZo0yr4rUXSN5RuHERckSL4Ou351Dm2s4NTXSQau
wFgvSaoLxCBZkyuZFUarh2APs0Wm7rqX2pqbJIu+OvpB9fiugI12dRFIoLP0
y8GYSMFrPIXrbsmri0wvSBk0RKq/+Kep7IebCbR0aasg0Q4pDNIG1PI7T0zX
A78jvGA3gvqYHzyEoDfAZH8iPv+eCvVbmqhu+9qSlb6LzlgozvtdJzT/bqFv
IJz2FnZ7egbgxRrDweAtfRxci+pV/lQ+I7PCEu94aVN0+X5TUOfJfPO+sFQK
hU1gqZqHdCmDet2m/QhfsfLHwY5/euGFGpmcuE1Gv2v7FjPHWpfJkg8VRaTD
25Pnpy9LIKyhfDxEEBr/UUYyqQ8rxsnXxVgsQFDf/wkcYwqOFcGLtvdVC2Q/
Naa4N0xY2VoAAEBRDrw7izw2genKtXmIRKH9nBtnHDGELYEQPf17hv7n8cB6
iGDIck7b9pg9bxxNGEf6BT5HJS1+Kxt4+E8edLgfVqQl6Wir6TIUhjbPSyWo
Ny7J4eq6+rOIjNYBiS52VKmvVlCmv4k6xi9LYnDyDC5C1a0HGYbaSy1ZJjPh
sL1tOsP1zOv9mp4bnJ4Ah7amagyEw5DjFC/JPap2+IvVQ1OFXsGF/YXkEb1C
yLvm0vMBUKxy48QfUFtUBJUD/KQ2F6H4d4/np2b0JcN4KCxkiH8ekg0qySPK
P7Z0V8d2pDFEbI+UyQX7fUAN0y8WGXhpN0lRFp0jT44GPbS4uH7TB0VsR6DQ
1/07vLW1bSRXJ8IFpU78Q+WJGgqXrfwUpU6e/HQdZIexuoPUdXkmQJFp/t4Q
XTGuhjgSA+k0VHCA2QlErTjDhhlpJDR48G9kcnThGPSnnE2aXWFV5j/Xi0kq
R+0FUrtqSJju8UV3Re2JMq0GssroTvmw57eck2GCsMN6jQKZ1rUTFelLbByI
d9qnkgCDj8NZJXBWERmbM0XJ725YOjqxniKdrtTqGUaFl63AsaXyqSpjPT60
YuaCJoG38nvoNYokMxdBftZyT1nh0iabiAKnvRlEJfDbMKMgB3BtR8VQGDpa
qTZswIviP65Jn5E2s3Jwhbwq4mZxNXS+c9eFpiuFMwOi70CS1O9nwB3O+Vvk
d/m4+h2XtKKN8K0J0U80MxWtr7bfHOzdG1Dd/BvR9bZ8MYnk5BL7oRMDkQAI
q6YPe0k4Sc81VaXkF+BZMmzVwxn5S+Oocl0/pEwROqW8sgoCYUYwj7JYvHUs
F+JtmBFnb5niF4jgSIYwbdAUm/lQbkBf0+DVxsTdggAousaDbWBDDPbJ3LUt
1LW6IkUPcPQ/gm1fjVa71z9zFi7raqnioCOzyRjSpvR4g2CJHOeDH7VSgRLH
bzae/r1LG7KUdT5y5dekRFtqka+v+d7rl6ZGwNTHyD9KFJZ9jbHY1lutMGJq
C2Vpmarc/Oirl649ZD+nwpR4s5GSIctWZg9paETd05rgolPva+thYwBAy6WJ
BbY3HX3j57rJX4ulQB+JDQTGWL+TFiS5Eq5jwHxNeLfRmxQiooI9KsnGeS4K
fhD/+gNImGOpmSAMGB8Ghf/Db2B5pSvXWWuRVnOToN/DEu/mxGcQILVJYRVo
KM7FMqc2Il8NtIF35FFfwDxrlJNw5nl3ko1B5tizpUY2T5DtIH+ANJcVf/iB
DA0wwwmWNow2b8Py+cjoij5TUu5qIvm+tLG8aXKQiobi4jbGknlgrD94Skvq
0aJdEt0/eH21WExdW1A5HyC7pKfY/PJeNacwb5uXrJO1+hFn2kdzJuvJjp20
Cn+dVr4CV9WcPIGMco/qP7819k0Gnb//iriJwzeeuTGmY2GlVqryK6Hyz+le
m/rH0gw3ktCtx1FEJEODtZUl+vsi5zQltpndXoNUePUfxh237szBGz6Okif9
rdm06d2ICzqvNxy17OmA+LgDKGbtpCSlDkqrzH7eHG9xcEugHde6lGe5SyfC
bM7nIeZGf7BzKZu/5H078Kn1yv8aAM8qiMB9BJqiMEK1TvIJb08bbsAqlCOw
j3qAcGyMcalngMf2gqKUD9Zbw3KC6nWtv38Bx7BjV6kAzcMdinC1rswjpoXi
gGyY7EYfQlX0/+IGRAKOXeIxkXIHRwMOL2E2Gkf5e1moNsiV3cmd8BIQzE+C
JvaiWzuwMnbjRQSGXgMWnlX3TERAHCm0QtHEPaB5h6xbRkmbwSWtyACCbbPT
keLLMAVgj56FxLOH87f4CP0Q7Ly7TVKpF1UoL2VQ8aI5zP5iPmqV0r3et+b9
9n7dpMmYLSQ8P+SGLss8gHjGeAeZwMTGrsnbOzlywHCFkiBGGVE0aRHv1h2q
CtG0fIbGAyQlv8oUS9xGWSsrGhU/E5qEOM0+PArNjoj1skcbfpj6SQJ1dVdd
BthsunevFwKQ67UvMc+hk1Bf+97MsiReFq5Nsrry67o3wdzHdIeb8/rLZvFK
43rN8g5lY10DVTqv88hUHHkf0N9hsLt7K3O0KulYEO4OeEZAmI4KzaPN9Y1m
7IjFcSOSVQQMaZRmLI5+3h5lOOQi+bV9r34t3OKFjMcAQWUX3QidHB4S0Pm6
3EsrKtbsDOjeFrsJPEgBZw5yL9iaqsySfKZBbZcbc2w/lqmU8EyxuA1rcwBX
r+KBZFHcmbOYkLLiN0ceO4L254Xy+zaU7P3HfNalrhBUiBKYOfMPNldB6Lkv
BTh+oOwnz733qjg7sItzyxO8tdkfB7uA/887lFkk8Puu6jAfZwoSGUsUxSXi
KmlFoD13NxTr+RHY7f+G6jcBf5ApPF//D9ayn+RAk+liEjE78e4mT3qZ7tLR
ZIiQ/FVWtY8LJpqx5C3+GhaJzcp/2MlMBeemwEuxWPgc6Cx/UXxLg9NwjPsj
M+l2rxu9bGM4dcGdp4B1NX1/Y9fqrsbmJNtfpFL0Pbv4SV29WQ0E7zJ69kaQ
rYsiTa5FEJZNxXEmujBIeLMsrd+4qzILUslWpeS1zI2ya/n2KDAcq4TD1N+O
DWsKBsRwZnDq6TXOhqzDRKmdUdsKonxT8EgaTuIsXfcA9DumUj3Euym7fKVM
lloTxXobu8PRrrNMNoVocQgCpUYvjebj2pZHdyW8pzjx24/J4NXPDzYJIrEY
woTQYLUP9RHD/Bynlts4YztEiGuGDpglcZONrt76LhGb+FD7e1oMXDruWBUz
pBmtnxIkn8/uLfZAaFk7x2y2CIWtdNFOWIHzSnnBipa4AHDPtIBHMqXPYe0S
An3w/fDJ7UZgbLPrWj6D3oIzi41kYRx08+dJ9fdM1DTcAAb8gy5CMuFeSzU2
WmsHb8tmpGmZQeVak7yfPHDIp91SkACFZ4QePxXI58pabNeECPww+E3SImem
EM/DkcqH6cP478v3+VQqvHmw0GoDM75pb4fcpdrquHWBhNbKMxtxmlfG1qYt
KJFsY6xVHna3N7WMJR+s1VOuzdXIzSrqXjCoRZg4vsi4DyBkCOOAPkQ3BsUT
5TZWJPMpdequTabep5KtkMzpGokoqoGHkMSvF8cqHeFB1ssvCh9f3jbgssu5
oGhVOQbZ7KV2045KVf+D8QxP9Buv5yajW/uC5aq0BVPj0FPwU4cFTDs6UUTF
yRCG7x2jjg+DxDcl3HGixI1lRdyU8n3HhYbsoOMg+cGwbFQ/BxXIAmLhGFsv
UI08Asq+4pfBd0B4hAXUAI5cWSRmcfPg8Yk/zxP/UKT7drS1ZosZDHIzyEiI
dES8TgoLPzxw1B+YQ1SxajISxuU6+dVQWGmht5cYeqSNDt7bSNXrM9Dhmd5z
RMkO/Lvd8MV/W8aOUHfzyo3ydF8hI3o4NsTjCNllT0E90tr6RrJ9I8d+m4Od
mqRm5ozMQ2UCvZpb/wN8MiytEN3VdkaeuPU+jNgixlRsg7DxxIr+OI3NnzBu
eBxDKmoG1ZTgkhU4RjYt+Nqn4PDtYMrxCpUWlEM+XJ9titMrJm9xQu4Diii6
Oa735+SwsZAaPC0JrlqeAGIktoJh6LBb7CGOEvqIXhenetV8lnsjjYGf1328
+AWTkbBnwP3mjMvndO6B7zgW4trlaWf2pKxvk05rgen3g4NbFpo+RNDb9cIH
1m+cfVuGwlR2j5EKHzdQ9GyR36m4hOe1fImTG/BAjCzVs1qQID0a46dZpFhG
/Im3w2CcT5jrOMdXpX8txGOEF3IF0JVV00EhneHEtjhJW1OzBgBD/85wOv7/
BzdDyVnpxgG1oVEjX6Tw5bue9Ega42ucERIDa8QwBKeH00tXcC+bUWoBUQmK
yEgkGBcdPUws2Cj3KAYt2txdzSOOgxzoAJRGuk86VocZHgZNDxC7LVEThBYq
yGTEpezWRHF6DzV7qF2jLRoXOrFeUhu6UUtvLyTjaDr+5Q4DiYHHg6oQXOiQ
FVROHO2fYR5T6/3okXvSR99y2o7Y2BjyNuPtFpcYyZl5J2MFxCXvaPtjCXv4
KLNzXBw/8zMrLvy/YzpcbWZoUBnXjryLCYEpwvWQYrudo73e9LQbfSb4uVyq
gzI9dKCQWAmk7/5GVKeHM4THskye18s8s3J0/sPWJqaXI2X347eotavawyqm
XeHpYjsOFXaOb529FuRIw3nzJGDEv8Gte7+8raDS7Wm8WfD6Nxtj5qU/Q32i
osWqPuoQFIcLls37tL39HRI0dBqgCULX+ru4ObQQ2YjKjuh4i6FcuKf9kHit
tO2G+d3pB9coZuYnlTnv85jm5RCaVlxYXf0ex2TVKMo+Oz/uO+OGkEQfIEtD
B1uKGR3zyyUSDtuFJsA7kAj6cAkPTCJ0lptAIa6O5I5wyNSR+j6ufYUtHKpa
ITP1RhtQcgQWxGS+86vBWpG69dMl5W/iYBzPisS+GZnZ+TAyY1wsBM/+Bdg0
Z9vYSEBlqRztAYXPos4WKDVdh/PxtOcYzQDRa+cjz+cGCKpia820fpRwQlAj
2+K5RAMW8otg8+1qoQ/HKba0N+4Ig9yaBfiOXTE8F6ltSuP+KBz+dAwGS1EQ
NQZmEqgPaA2OMuCivERaLmYAUKol8uYnWZnC4Jc5ZoXjeUgDhiHgexCAfeVE
juGnmvpLi3g4sHnUolejthBHhLsEbekM9tKjByagrrZYdvfsp1p+eNZnGWV5
ryJyAT/i7rZrinamEhXJXwPPuckzqcK33Zj67kPV8vKVbs7UkYthssQFLw+T
ACuBPfFVsC4ZlUjvrfU5sLPZ9qHOF3PJGyvNWS2n0Ac6IAlBKQQ+fDAAKt2a
opYGOVDp9Ry5RFiFAMO7lD+Z9L73VCuK8B9+O+uDiQ6QUq8BimJJHAXxj2JO
DMKocgHfhN3BN6wT7G2NodLcYZ1azyxb0kwqOzIEFTQ1uZQgCiKZxLLt3UPW
aeVijCxSy/WG4tYhtHjD0Rjfw6jXKcjB8OsJnqTmITpGdj/cSxxcy7dtLs7G
X8dEi6xMiBsRLfqglyXaM868nYfGiECybmhg/sPQtQzlrPuMW1DQWYAQKl6I
buhHEJTE4CVAKDQGLfeU8axbeQR8MeJozkxTUF3Lv3YoFozT+KgnLIPiWFYo
8Gr9uUPthXwwf4ixQXGBWOrlhiFgU0aqD+/LasGnK3lNVSFft713aQ/rEZR5
/5m4oOo0CsegeSPkWJqIEhGlMt7CibKW0atTqF3HSJ17deH/q3lQ6nYDJ25c
WijEuoVu3nODYjS0sD6fpSDQ5gtQ0EqW8GRNIJ8jMpGJthxDBvylux/sRs7x
xFRhPKK14d+EVG+LqzUSAQaVPAs/hYdm6Wt5pfFYGcx16OnGxVtN0vppSlwJ
EoJA4h4pIV3o2hz7+TwWj2RLONhFrp46aZdUzhNEvx+snO58qHdDuDK8gaTN
WkoHrm1fDkx/OfRE4WrgRB7Eo0wGcVNge+XvpbCsk3q++yDKJYA+3tt91LAr
1r/bJwYFfzEqtxOruElREXX393UHjHflw/4UMxWZEUbDNFgartZoDh+SXTKs
FYH1wY7JgfHayigkaETagl7EED1/C9Wt3FAWXIvOXPXchMgyxpwHy2kGpFv8
VZMAcP3OmN+v8fH0bcola6xt/pJpkxepk//1u9YKxPnbLW4EUVziGYLUDt/f
s3g8+W9jILnmPHC3FECHcL1R2G2+LgmLQaW3bolLHU2oYsBR++QxmMb5TT/a
m9estNNfCzkJpMXxq+h1y7S7KoDvr2qcmIvgOK8oII/OMaWfIs033MQNVcjg
sXZBwy65Kozr0sqXxoq3koQuP5jhV5vWyGMcsiC1mNo9HaxEtvrbWCwhJOSu
vAte0CEi0sNRIMgjZWN2dNh0uzJKaTbXcVkiki0seokeXa3iVj8qp7OUDcVD
jsgOJyvaGUm/J50L3JuzSXH6m9qigrZK6dwlC2iMgCNVqHOYP53Nde8ZTVOg
oJHB9ejEq0Xq3hcaARRkgwpWYy32d+scE6TMReOMya0wPn7qD+hJDeBvH3Lx
yml+0rQ7WB3OGlxWQTQ5xrNFWslKbcGqcsWnYedEwPW/cbeGsMedQDOJQTzj
iYAjDqMTECBgl3upDAztT1BAboQVT/ki7M0Rv8/rM06fYWX4SHV283hX+Bn3
2r2pjekX1yV0g2OLvg7xDYsjB0CLa13VIUmcud5QtWDC0eoMstnq7dUFzmNH
1w8ndKMJSJ+XaOls76d3zIQx4SIz7GKezsNOO4lhbuhKUG6Fhg86CngnwRQQ
bsOL6fvjp+cRp1XAXVRz0a/tkZVKVdvZIYMvt2wQtTw2+8bm8R/W0QSQNkpa
Bkx0Dnna/bSdBwUNVKo1DqtqiqRQSQoof4qr9ieI3oZhsERJ175Cu8dVqBYv
FlTIwkkqapIz+LslSFbdfE7QCONdnHVmjZf3ujE9GXhMsteLN/NqkXbMVKyq
xNqnMtwRabO6sxlrAiHRhFQErNaX4REDX4l9VuqykBG0w7pCXDQR9cOldKqO
RdA5dlJrpEvUm38W4uSzkgLqK4PsPmO882KpLL9l1JklDXYJV45b3xb4Uz5n
Gymfs2PNX6DH17755wAENseSUrK86yD3NL67KbukDSiVHu2gFRo1LIz0qGDe
Ep+5lUhAcT75mqR531019x5sH1xVQ3xJkju0TvznFXqxzMS9fM/xmDHddrcV
hlWZGZ5O4Z7sPIIgVmYr52P+hvXyMSO/fClS/qCbcxMmLJ3Fk+vs9S2tPaDQ
BM8bA2QuLT7/VReeSDY0RVdebUKTfLRdaoCNh3XZy7rAEXYPrJi9AWibQoB6
8LFHS/ElFe9zRqq3ubaysMPjYZAYAIhcLBY27XFd7vpQ4yHzx9/l7uzkVc4u
kPuh+DUf61/g9nn85na2wStzwk7Ma2ZNUBlhzotxpGr+/1El24YzsF5Bq08w
JZ34ypgMacsnnaS9KdZh5GUUBMXOW0d6LB91CH3DaZW+oLCDgwJKU/Ab7LfW
TiThsPqMWiNFq5J6Z96W+npkdnXOmD5EpDdmXD8pYVVOK3WFStuginETO5e5
LEYfKpsL+Htic/0NUy2u9Jbt8pGKBNzRCeg4XYaLIBj/O6LU/a68PaUfp3kD
I4Vjn9aAMLFOKsZQFGBvxPyGtSZjez7vIAHlmmKAvMa0Hl/Gq/R2uPlPiarp
vJJ8J8FEQArb0t+l9bRutuSsSDzYHNfd1mJJqfTrwzpHW6htYKzh1wHJJXtK
8ng4dq1Jq8o6+v2rQ7fFzwsCd44Floj64RdRFnTiuoVhSQyiVjL8nb57NW3g
iWPuoVoFxK4zfgK8naiC8tUe8QPSe70Jt/eIhGWo9ZceyPFBtkR7hfSvmZ29
xOjknWbE6lvaujEUBDvfDc0olh6kC4CCmFkJzKqocTk0pPU3AhElP36E7uIH
JpwJ/WtmQGDWLMmcWY/8EeZ8WXxSGHmwVVxnbCl9Co2Rh9Qnc6yxJXJY3ajJ
fJEKwVX1dqnwO/wmcRDa3x3hsMCgyk7f/SXVaMqDrm3KREXYyLQF/hiZM0ls
GKtIJX1RNaJVCchkqYJvu5zdherLR3iTt8O9KdGGVm7BeKf56yII86F/NCMV
lzoyIMlM8Uy40ohJLTnMfT6GV6SaI7Qd6Iz1o0I2xWjS/lBQzk7QjqKpemh1
G8O28Ep4yNBX89eWq2RDbDfUOYOwYVjZLVfVq5MpsCnOBO4jziH2Gyuo6HJ6
+asBgQEU8wv4E+qodQXWCnUL1usUI09WYoMP4jpE570X0BsIXU22kNek7MTq
BgqjUYn7tZJY8hhKSAUpPDn66ZVTBTIleuNBAMb9RGx3ONwX+kuPOhop/IGN
YhOM86dqKMn8yEwni4eo1eVeDhO/b4DnG024eMyRWyX9GtIYWCcNqwIMFsHT
AMeph9j9c2soRN/5GA2NzW08j6Fd+1MEwSt0LBDah3ueO4OHbjy2qtdfZkT8
Vj+ucbQGDjg/rh9NPzS39DKcFJH9tdZthY3gU236AAkzzilX5qit7OUWFSdj
qr88csyhJGhf65D6LW9OuIes4RoP149DEv5rC9rGaiaJAF+y/r7rlDUdktwq
Mn8B4kYdEyo6fZaBIUzqRpI/Ah+mQRAa5bCFNSUs1X2YAQMDvU/xOH8365YI
yGDDTRejQhPUZkLgpftcPnUIedeq9D8SFvxmL5yoSbmBwqrcdj1gA0GPYJdH
KDJryoyQ4chqKhGqmO8eTM419nEKyo+w0C7/66W68ExQRQ+Ss2Fcz3tf0/nQ
pvOXQ7h0a4ug//uUiI52FyrKZ2rV8vI3xezWc1Ma7rdeVj/XjbHYsAymIc+0
UfbvfL0/hNuItuQjpzZhVJHQZ7SsJFgSGqPgc/Ue+cl296IlNbzqHnpN96Ci
wH5u2BwHvQbNe1mYa//aJUeDGShvCZdGo+wWsRLxT+L9APSaWkgAtOHhKLxv
5ZFO9YTSF/SguzA6RSeZCcpH/iaYoRUiIeMVTZNfdefc7F79ZESqqPlP7WlK
cbAKVFM/wV1D7/n9duXTqmMxTtwVBA6DlT1aJlMTrpX7Hxjk4cpYm7VyKvkV
kWA3T6fxgjqKYbFHOPmutRVkQuI6z4yM1RkvKoMqtRCnFk8aaQv9jY/sKh4H
bDFtAjrg/b33o9271RGts4aaGC0bDTQQkixOcpFvtqRy8uE6QLJ+g7bSES6f
Op3lFHorDRdEzhgc1xgTy3FgwaPE+vBzky38maKlinY6jxLtqi/pEojUnHm7
ChZBLDpCuMtgIKgThYtT9cPLrhlSgFoqo0kLCIsdH+6KMy+Mdhq2ACXm0b0d
xQxX76XSk+7JRGj+cqyziG5vZAqBI04gj1Nf8K0f6k0NyMCn6ddAJEtfIaLA
za0friys7ObvKA0WCBlLHLf23PvT4ZRnKxc6n3pEKaz5k9q2UUhkgSmhWm5j
kkXBOYetD8MWpgg0b2mjpQW+/DGFwM0XKsJ3c3UYlX9sXe6lGhDVMYZVJ+3b
JOZCEndMgVZODF0T7tboD1OBe8dNMwKrAwO3qSbTkKbJCWzjM1OVZbfHncNX
NaDHZgOeCnZKrIRIJoHa/vL/7RMPkaQVy4J19bJYqmZ1e5yVBt5r9daEoOAo
ZXvn4lFXjVB6cZFpXkp58c8BAh/JzAUt8YEipjTJxX/rZLgMiDtfzl9f34pO
BRd95xbEyQ+Mtp4qoo/YBTVNhs71lNgbWoaGFXtCp61scfw4wDRb0Xf+Lmv0
G93CLSI+108fYoYlgybaosica9UG+6lhp1HQygKhvU+JT+im909c3MFZr6Ga
sEsN0lcO0mio4BUytevYvLkBkXuAnrLn86zBGRXEK20SInIZF+ptMfh+FZv4
5tJWjk1mlJQud2L8MRWQTLBLrM0v47EM9BCTnOa/UClcnai32jyB9kMgd9Rg
M4h0+3T8Yrr+lIyDcSfx7iavvxU1sed8mKYMGJ+g137MkScijxMkqNevyxkk
WnMRK5W/HkBtJ1Ft6c4oXtusGF5FbQZSUgvCXOVvFVpW/kHO92uqbRb4MAgu
vXNZCrD9bgwIR3L0pIYL66LXEVuH5kGXYMDcqromHgyDUYYIy2GOoUTitKfg
uZgUTfTowqTY/yqElTHRhbxo+ad/USkP74798JNqNiUgGmkyXhWRhUPssGLl
T0FhfyQ9DjxexRukqN2eVP6dXFMLNURvQjv7+GBgtt/XDB68tmgWNpQ+42hf
Jfnp+7LutqTjdyEoGPhXPbM/XCLYp7zrovr2Jmi3MxlLx0YFVCcU3l4HRVyp
NAvqxY+3Si6RJ2M/6XaU53FhnCcRVhVzIqmKjdYG50cSRtXj0LlEaSZPyt+H
7AcboJgXJ+7HawkD9YiHD6nX3u+0PIt4uXJC4W6SZQoOFYaFvt22ppWGYBo8
RgOU4Y/9a61Vb98ht87LifBdRGm8465taSsa+nPU0wLyDW9a9h2DI2owwMu+
PPe2Y34BSOGvPQHFoBCz9D6MErBNFyX+i5mGHCWLO38/OdDyXnEk7Gid71zG
5AigC7a60SnNcUJiRRn4AXWSZr7jH77SBp2lv8odcEF/QBSHUS2WBJAL8cYE
iIa6Law+JsaoPUhfEWpuZ5gxQsp54wjys2Nm3gmR4sGenM4zTFLrNK4iG0BW
OBaRH8kfnpJFplybCZ2bnZTYm+2u/cJWenQhgEUMNOo8S0t0ALhl7syCb/Nn
yys5uxC/+v3xbPhILoqhCnPqR7Gi5NRZb/CTzsh6XcawEOTN4E4GtuXRt7qN
mJ0ZPgUF4rtsn1z1tzWdgsnVLpCsXx+WrJF8NpZPTdMxyB+i0eKU8q09vp5E
y68cBsGwWeeotQfE04TXmSkJ4/HwJDMBwpw5UL7wTYx3ZaCUeFoZ19x+Qt4y
9NkIsGt7waf8ZSSVYy6Ip7VA6FyzXmhOTXYzT5Lx7N0a35Vp0CDKFBK2rUJj
My0v8ggBkossa514GVS6wRiY5UdfgrQ59SkSB8Tm2+XRMXv03eTBqMeR4K7s
mWkoEF9pLGi+/xky4V40jp5zwxzaPU5hpSn8U2vgc3uTqP8P7cd4O+zScJE6
5E2YzaSp49POjsyXF+RPvavVMRqfmgqat/r8zrWyDyuvl0ctYj6fdRcinon9
uPSgp0nZPut/q7W3ewAeinQvTyr6Adzndy68cL8g3/Nrm/V9dzvrhu8Nm/89
8548SkCJ8H7q3PuaFQIa4cuRvlU9GWMEq9gHgtFAFEw3qc1P4h736q3CFNcl
T8ZHnSkT3Ssn6uCnUZmmxE/xtypfDJYNk+Use35nGM+X439qgmP45B/qs6IP
uWj0wW6wwZ0+vfZGvVf8oxfMxORTs2/mLdW21gCp1A9rlKs+pfAt0A3CuSuI
jZvPvjUI2UB+zzMy9CkwnOV/EMpX856+bRVqEvXkN/hU/p8Cd0a+G09X6NDQ
vasHVB2LCAo1X10kcObqbqDFMm8+WfG1JNOmrQW1/gU/moosmswBUj9ZNKq2
/t/ifwdQYDURsZdZNnpIJ7rTnZL3o8rAEUJe2Btx7Wl+UlTeXid/dDrI2mOv
hi1Brxkl+5BnQvUEpQy+0NEp3RYwfJsAuRbzStAmRqOo0jA8B0yjMPPD6Cb2
Y/OAhSMpUbCWSHsnxBDUIZcgSUhQc5O4FixEgqM69HCWucBwsRqt4NBGGfnK
19YF9Hz+rgflfYdMjua9o8CdysgkVbus0LzySkIyNvRM0ZODeZe0ahuMOQOB
SOi2V3cqdvcbGKRxUhHIFUgKX6CGaKvjLBUsaMVE+ZrK2JpUqMoS7i+ql2+E
5ZedzB32ynxchNGdbULB8JR/eJDt/7K6rmBLWPDGdLRHKPw2qcF4QCZgh2kO
1K+6oXWMWYIsgVNK3XT76sqJeEWJBuMIHAapjRrScTJlTBinuOc1vUA7CfP8
we5D1RnkaPY1HioaPosnesligqXTDJhOjrah22M878+lquIIXpC6iCg0F6ZO
Nl4Info3vTGJkWMPfX7OEF95ITWRqa+jCiViKYcVsMWv/hrlEkgOAGYJmXZM
iEoTBps9AqyBQOMJd6lMVA5yNUk453Fgj2VB18i0ZD3ek1ZDaGIuZ8dRufla
3ZV6LfS1/rwvDV46MEnWySj8qynLqd1Q70K9r7/o7dcm3vv44wYMhH4EOsFX
SXVk6WOU2BJKxjYT+7d0CxkHHXIvbspBIQ6jjgw3BSAUB59Pzpq2V18BMOyy
xDkso2k6sU1XlrwK8vlpoeUZq+cZfNcbbtDwf51iqxKraVfRJ4fMhVForu48
s7o7lN9xVYHMer1NyI+c4pggkCjKupI2zPZ8eEmxyvstLC3bw4mXJGAe9rjx
s6iL2WAAqHUpF+74RxPQ3KbWJVyny7AuaxmfsU2k9fjuW7+HzNZxyvY8nwuF
IJEr4WiO90f1jt7NEyNnoGG1HMTpVCiLxD4p2TnPVWpe285/hK5WZVB/PkGZ
dhS48+IoyET8hqrZBBRafoCVQ7YtYAnXFeitzjczF0Jp5fZf2gOGVGXbCQ5l
87kHKz5BkGXEaq2IC2PucKeQB8lheqZg/G/2aM3vfETC1+HI/ZqOwVI3JQ/Z
kK+2gbWaIK3Q4An6UYIVRXxqRtl6vPIqM7erfECnchz2MH85YIRweNqEfiDV
5QqMsIki+GCZRVhppeR6811HhkGtPc3K8z1zlyF5Ntd9nAfwpMw/rYDMx49E
AOSxFx3zUBQm/1FR5NOPKHkfOr4FoqAx5C4Xq3vRKxFfPlNlIz1rw3XlOJwV
sJ0TZnb+1bhw0ztdFe1QrJWIUrO5oRAwoRJz9OCKtVYO+TlQtaieMT/jseBV
81gCf5JmB5swwdf7kYaldq9sK/wE+9W7IBlM2QTee1qEpN/fu6FQaagiFZov
1ux4mmv3zEgC4L+6ARE2pkCMzaQ6hSelWu59CjiVm8d1eSSb3wWPW6nZakKz
ESwjzSnS/otnkrBzqfvY1ms8aXUEWpvhU3zx65R9PPPaiH8yJhffu6PGv7Xi
A1ZDtpNRC8qT6YGVwRDgdZ2QRLx6brov2AX2WELwrb2jRHXLvwdSgXIIWf0p
UnqEbqsNJOMRLx0e2cOkIyfl9T+Zhwh8RVTd6ytmBnapwIYBVHLntXBtwuPa
JIWgl57peHUNNyLvPWg7VI9gujpEnhDXet7SlU7CngBNflFcy5t3smwunzIz
9E07gtV2NFW8dWclSO4UDLKahgHzfZ4xEI7M4P8EXQkekQ+vnBnUzG5X3cVk
h1PQPu+gvG18kRy1M9sd+gJ6E5vmz28U7Gvabphp4ZDinQr6hPTJ71E1YXmG
bzYqZ6jQygBq53b4Nyt3bwqXUbyTpL9gnicX64cVttEUeWfy80/QGRPh7YX6
pfFxnCSuyMTsrFaQDN59mgzpf7rRXTZqs42YDpo1OvBvu9r/eogn+aij0JWa
U6FyEMWSt5acscl4OcMdsRvMenkyJYH+QeQhFCg4942sfp4AEl9JhVXU2/uq
gAnQTXagohc6QDPuhjf+Nj1t+AoB0/N+059T2pAutbyxh3LJRzfGprcvM3KV
9hyUXWMrQchZsn1Vq7GEjTstloaHbPvKqzZjHLPNBzsNecAkWp+d7eaGh9+a
O/y4679n6DDI4rrerwaZFd10LDgc5Fb2q5FeBVaTVodjZSADyi9xP2a+DdEw
r3TdN26eDzGRZZJMNPeD7FqZOGw7nW1i16uhats7jWtBwfMbvrRG9+Ecs/BQ
KkCipOi1Oi0iUdATw53cP8sNJ8Ouilh3JVWLewKeaEcqFNzqTRrMeoaqdgTI
q6Z9jaUxGo9XJEnwkXSB94PoTpQNqGHKzvkoISMIg2jJ0doB3e+7fpd5JvaH
jWi7oOn4+i8tMsxVzGocmPV254JaSL0DkJ2jY7HQdB/vtmsIGnk8C28EmgeK
kuXveFNxWK1IVN7oOob2+xKdOFnQp0sxSHGBf2jTrtXifa595d0cn7MPEqgX
bRXPPKwf+H1XsAjjUBfTg8BRmsgXWi12p8hk9JQmoGACDFsMGr5qLvVjTI6i
sO06eAr3QBnfCB3QO19bevdg1/DUNzepq68IvDposzMTUuClq2GehzkiJZ96
snQMVXq+XdadpM0O9NDTIABoazdchR0ykGK2aeRyWJmcmTW8fIJrnfVdUvpg
SXJobcqX5bFzeuygoRhzjCaqSVqTfV4mdNkRJcbEH1WCALjyW0N0jKl2PCIl
8FpOtSw7gw3TfguVfSyuBpa4LR/jIQuq/Hy53E6M+VJ6VEC97gpihu/MFmnY
ld6MLXbzymvVOdbgcbYdx5nBjmJag/qmXqo39UohIBpQe4kXSyyqTuMGiigQ
0OBmMyZca88zrGjbyZL9OZ+wcj4HPaAU+xihOsqHwNJLok7zqbtwO+Dyq8GE
+D3UooxI3N+dH0gLj4Txs0r9eWq3CMvxhRjc60tJXG0MF3ZBqziB2jYwQIL8
VzH2cRr3tpbLdUY534KHJ7FuXQqBFZkB7Q4lAsl6E5ugSuvSRtcLwM0RRLSl
nMwW3qZy5FXQ8u3LhhHhgFxbiJgZsegh7amM5cN45Bdzu1kWZqPT+luxA9y0
3T2QG7gCBNixagUBluOOZog4I5Be8yaa6bL8Dko+C4oXJZwuXpmLjE9I9wgm
JSYoBI6nN+FA9+tfPpF8H1ZyUPGdvAJfI+LwxUKs9cIwjx9dHmJUb+X/s9M0
setmMTUjRE5CUNKhr3MOWJjcQZZJK/UGAz9MjjbDqOl+l0WRXgVSvEoVKFQj
vpQBzLMFBoUW0BWUcmD/qlw/zdJa2TQkpxcoHDF3lY3DFtDV5FhW58qbnkzb
R8FXQ1O9mLSoEwVw0Fgaw+T4miC9PisjirG1lM0pA1OYe1tnX+74NiIvvF3j
XcLHwkRNlJGyh8EahIW4HYAFto6a2C6ssPWeQbx0hHCH1j1L1ttOYfNJRrK5
ZXfflLpR0iSa7bqAdc75hkWN0CwOP/Ji8/ISFjB2FIySFgWONN/IxnUW8sNO
B0aMBLCpjql44oufoUHWYh21n7/n/MSymXuBCDzjSzg09ehsqUvEnvNKAxk5
g8kKP+SFgXJZPPoWswLlKIzNrXRaodWCAlRLM6/BbUT1NQtSpeB9NPa7GNvK
FI0dTJRDkkZGneT7mls4LSJyKnPUKDnxXnd0H06m72yqnG37KitLbOMosGUJ
/nuqhv0pLRwlMBalpWsBaKUzqF4CB6N/rufTwaHg/0OTEoJtR4nJlo3r7deS
932qMsGGuqctF50zdgbkGETcKYxfl/BtsDrReUvyLcTebl3VcA2jN6/Q6FBT
VUKHNDz++bP4bWRYvjpygIb2uZRbwdCGVn7wHAt/TQ16Yaboa46IYR0e0sZI
fMlCj2izsFclV0lX6OyWz2OAAwkdgGJ762kYHLyemAVT3bZkUmyYcBQrE9k0
hgVMifYSSjrDHt7bDwc2WAEEfR/K5Z1I27KHxXhlPuLLW2wgtPrxREIs24eY
HPa1UAf4ZmM7TYeQgrs2/6bMNQfiXbwcjFSwX5mFCDXea7rJMzZohM+os5YM
EECcY9zoFggG2dg0YtoVh+stzeCdew1xs7z2ClFzX2xpIC60A0vlAKEAVINT
aEQ3XM7xzovT2PYUBW3jnAzUr8TmHSuQUwlkU+Kp/D5WpCgax3wr1r/YpEU+
wcoIvSX9OzJu0iUMx5ysqWSVtbsdr7ksJcyQQvujt+/H2scK+xgZqIlid7xT
YMMiGtf5Oi3ooWSgFM37ksM3oASMwDF3h8ai9mRNjmunKowpfSs0zIU8S0Pa
huemUXmttj8OeqhA661zcYVxyR8hG23Zs8tbGHV9NffvhXyTJx6wKgL5P9/5
BFyABWmoqi+/hjG3ec+rpxodqDeYdCM1eu6LdYtF+oo8J/w+5t68chOUNYSP
wt3roy/6IcG4xNGV7J758IQ2q+6OKV+PJVw86frUZxo5N61ETwzAsIGrj4SS
8GPnweHZ+uVQo0ZLj3w86RoNepZkzdRSo4LmIzBh4frKT4pTMnPRHAGKns4B
p53icsm40XXOCssE+Vvg6lu+wY64hwRReX8gBJbscE3lO18/6njZZCWXO85Y
ntF4Ez7HhBIjDRkxc5vcEpNid/Y67x+PjfTxtXR3Djoa+wVKoVlLI6uDBy++
hXgNa1CnrgeQFX+ZybvjMIcwFQg/Fhtm1SQorYklkX+VC3Cfpu4+qGc9w9vd
AjoiHxo88KdZj4i3ASoYN8yItU/DUyE/qBNxA2Qfl+LENzlcTDhf5u9Sbg2T
gEOCV74g3bzVXHxnubsCNYSptCeiVSBFIdfvl/337djS7JXdtKQpRKHSwiwa
t/omvFtaPfkUUJa0g7WkFl3Et4iqKvNqPOhvKIxPHcbn3vdb4cPVUXiQEa/A
IzJUZoohiLeP5kNMwFEpasH+9tQMCdLLqY18Hj7LT42T1CoF8tOR2hjdvXy/
6easijGc0mjrxY1TW61D/UdlEr99hiP7nKQPaNqfLLFPwhhIA7hwzY8db25m
836Hl4qAsc0RakwRpCd1Kk6IDGVq4CDT0a0rrJn0J7oTgCbcYa2cCrMNfpKy
JaFno4+1LtKIqLGfASQBkjkaC0FcgzSqY3MGGT/V9/sxL91fGb/1V1aO87wo
87GUQT6RSF1HQ4urhUugtbh+FZeQea9hL88wb+b0hRXbWHcwjBhK9KuAZear
L45XTgI9DBMp6TNSRi5B42eNiiYdrvgYg2Tm51PN/22fE6r69maXDGpRQ2dF
t43nKw4PokNo5xhJ0JFttL3ekK7quVPCQWIPFCTP2q6HeRpSUqAKwoyFPB2G
f6hrXmOVcojtaTAW16Hup00U4xQc5WaEaCcibxVgwJllpPgd/dLrwxmTozz7
b3/76UfH4CwNutBJHxToDckkoSgUvk99fjzFk8CKD5aOhoaWAtbdMUCy5FiH
FqsB3QPLTwm/Q8IiyKonfBBugrKRox96qHYyhlCpQi698C04bLdLrIVhgSh2
1RuGzj5Ol/lbQT/bSh2Fysiwj8jxvtoAahMIMP7xpBr+/4FqDhV9+imyXaOF
0vdo31Yb796K1h2mAxY9IUNC6zArxav2tERqA/GoGJ2gUQnsmgZHEG0nqUnA
vQVAiarDox0NPuy2RyVY2niuJkU/fBWI29vLptYjePAGmrgBwDIdO5rnlaUl
flI8ggQwNfEWb4RSK+Im8O3T3E0indD8A4hkFfLLNVpEWBN4TjRlmFwO7yaJ
ZrVZdCr30uqns7fRv9l9WhNfrmYB9LXu3PCVHSq6njoRIRllrJKls5wLThXt
6m0QpXqeAXFZnYXpsSbLOEtQY68UHZsZZAL3Oi16oANv2z1KiuAxwXcf3Oi1
ILmONmzeyqtPCy+eZxA2iaAqKXu8jtk/paLWATK2enml2mxiHI6WfNOjNvrI
SDIuW4zmTYADUdfstLMaw4OnFkvac4qQqyz7jlmh5A+nRHtTl2IX56kVUzKL
x4RiSKFUXKUTlRiBAaHnlOi4WwAbeKWz5knZM6dsZc89tIo/nSQJdErrmYwq
NCLSFjlPQb/ZGrXsSHDNm+0LlCKYe34aRjMnQFpg3fNNVDoyF2xjESUCn2NF
Aj5xeO5pplNTFblDHM91cPv5Ct0ZFatOZ6fckszXq0VPrdMbalna4sukktVt
wud0zEQ+AQDaUDmPAJatHmbxBXTvJ1tw1b8KXrIqBaM77iWPNzjcY3UWv28x
LCXqGki/32kgAXXkOOhG8n4lXWgq1uNrMmTYmiosVeh3OL5pz9was918RYVI
5VBVDAmH9Pfdqkag1DyunlviIXExcoRNCk1deDsIKayQT4IMKw8tf5fIRoVM
H9yORrKBv9z9nH4aitRlCXdLQYqE28NxxJZDxHDw1WwYXW9bFzk47jjeltH5
4nkCdhdd5aWkGc3w1yH0uYVnfk+pMuV66/O1sXbo4zrvrLD/BLr6E6ufXCIv
NAtDO6sI15S12u//oNJtoi2qT67uFyVTU5JeZ58jtdRd2hxyFuyTgHUnMRnC
lnTliA5sfApTbGUaWC4eJ4UtnkRwY6zspko7R2rCJcSQcxUdxDd6NHzaeIIJ
7n4fpQEO+S8uT65us3rNAaTk0S9gm/eaTRums7eGZqI22ZZvDUJ4eBHNhQpi
lvjVyBt3EYwQmtfSKJRydPawiqLZHN/pQ/DLovOc6dtCdtisjM3yHtxZuRO8
TkEhWnuL5Eth+h/JAeul1DBWJZGRrrZpKVuKZ/GxPBVN7u1vvm7QMtk4fhs/
RN5z3PEgVp2tmRABvq7hXiH7d0v+vf+UOhFAnqixfXkqRUR4HDcgb8In5ENr
dMk+fUU0zOobpWr54yRjsb6aqJKc61aqZLj8iDYldhf1oRkUvZ91b3tXc3F3
C7HhjbAtS50bJwLjpjUyZ3OOmN7ByR579/C9E0UyaGvttqU5T7EvEs/Hu7ni
FZ1PuNAUQnDQw+T5M/4bZljWR8GJKWYKkfWzSj87D8LzSIhoZNR/CHjva+I9
OB8z10Ja6bmZ+NHYnVe9kXxsCAsLDaqhzZsMV29FR0C9XmKwVgqeFMxLDz8C
FJWpIkZoGK1bo6RcMU1kDfMUgfOciJawirk8x+R00SWfhKgMo/bJuYJpMi6m
js3XMLP/fprfDaad3Orgpf8zBuo5UZo4Dr/kQXRf1/wkGD7arlBuPG1i3eDn
dX/sGFVPlpmCYwudEzsoSdycNxSk0FhTjActwMExHs4WbW9wv3lle7RO30Dx
brpjxjS/so+TlZkGSLDHsYLToKOoj8jfpEQsS/eHxxSInsseKttkmjf5VFdZ
GA8HcIUcF4IbFcKAGEceAoCPuwBx1XaSajVFJesyRfT1b20a3A8xkcs9CuRP
m1NFGokOWF/pQUG7/p891esVwqHHj/vihicI0n5rMygccuTgvI/k3B4wyGr2
b1J+OP99wmHHqIAbROAFzOtv/ll2lhOo6BAh2pn+kuCqjSlsGOJEiAp7xy2q
WYXnMNIqbYtjp4tBtVY1JRXo01UeE+ACe0fo+uRa8o7zRieETifozqtPVzQQ
oejWumxc3gMfSaPlw9l/GoM3Sr3UNJxtblZVdGnj2ohnTNviwPFoD6T/lAcn
x4cjzEMDS5xIQHkxEOn429JmcV64f/kDb4pxyq5MaShBB8uGTWlpIHL9DKmE
+KSDNGGfwrRdt9uXa8MXO1azbxiIjE9QmChYp0WDBVcDJC0iH4iW+Owoj91J
InqsfudsYRLFIgNFup20lsmhUJZweQejnJjMOO4DlGqJA6xiUGjFW1GWt1Jk
CwKIiOm7RwkjqRXel+9obknR/V0lSyN+hpm2kBvKrC1fAjORwjMHhrFip07y
WyDxkXc/FKFfrO83TNtPr+v+JXCbwD2oZxVw0RPwW7KZmg3JG9K3WaU4S2TR
yipyR/tVPAwnGDXl31q/prgLyNErYw8hJ9BXyrYuOdwqKXJbY+c/m7clzO4k
hCBHmFKUHswwi0fd8kyP2DDMNgtopJTxoX2AAAqNktB0wfjY74TDu1WcfF72
16vWu5STQpYm7tC70h+yZf5XodzTndZfbe6fDdo/L7ZeQdBNijaIrnmb/NEg
jj9Z8MOAw99UJm9ZYm6dz+2NRVdjuf+nUq3n/rDLAGMRawIAV+EwSSt4OBGq
fziL9fSqMl2onZvcsXvT+UlrrwntnZkLMKjdO8rUdwI1oThF67PX7QivwEZJ
vZQnO/Am74wHwssi9OpiQSFgBf6Mgz3qFlahanS/+LdBHBk6/knSkiNztqgm
7TZhd5VnByg/l8e4+z3tbQc1zG2y9wFok+3xAmf39UBc/wY2hfHRBHosZgiA
nsjRUxQtgLnDU/glSrG28rXZbT93UrLNVhkOfjYPlhy66EdWt9wxx3CkBGfD
zQdjCWwWskSIaqYrfR+giEr9wQRZ/zFrkQgAgfYeZn9OGov4BF/Je9wiN0CP
hcGLgL1aXlsY1CJvSgu0FDrxHjyCYHCqr7Mbr0ElkPg1vPQNkEGE1ieJczsh
k0JEheFhG4qkWWW0i5ry7ZMY1VdBo/2aDaTMhXNP8GhCrAcBDbnUlUMhAyIc
6nARulZnChXJnk+AoplAeQQs+/Qm/iuexSjJtnNWEdvvEMRZ2vN79OCl9lkR
L8L2eY5W7Q9tWnBvpJSSh33Ri4I0eTI90FJdy/H2OeDiKR0/262DrN2jK2G2
d6jBgnJEJMuNcWExQ+ZU2RbDmYHSHNtBvMkXPQL+J8MDxAq88IPuaWDPPze0
AQ1TJIDQN28nwuKpJuyHQz9Eb0VGHzQmyKixL2IDHJ7bUswcClFG/X/JF/ym
8G6AudeUwMWLgBYG2VBvEU0gETtQaW1vbFAhyYYpeZihNGyNaNiQxskuHjWT
ti2Xv6oR0+cWlicoiLjogFRNM4rCJSlOk7bVSxU8hD0mIUUJi98KKKIk8aMy
uKph8pkLNMxHKUyIlClNlb8NpF4xVkBEenp6UhzatVHQQnog9JoLte/VT4DM
mLXC/P2Fd8dEYYwBYlEtQhS6IZTxBPlbxKt6AA1jgPRg3gdeY3PIYqA9dFxT
iQoNR0vLpA2dYYLC+74fUaZZCPuhlLxtgF4oIYFs/s8ZivPYQGYz86I+wvp9
VeuB1dZeUkXDzuBNR7Uxm5BZtN326/1c+GudAa25Fiz3v4cn4KB6hh0QNcsn
8h+HE9SXJBsJzSDxbhJPVn77wTctj3PzRpB32zMRlq6gv8lcMPVQtwB5tb7p
soGCKBsPIa9tEy6m8lmmjK64djVykpS7FQ3XmcWcQWo49vTWI3znBCaqPO64
bSqFrv/c8A7cfRO3cyx77DpkBfxbKhZlCSZ9WsvZZgDs2YGY44tQZWKsIp+S
USRyL1qfBb3+4ETT558s9c0ze2Cv4JzIZ+BOLAun9te8itLM8AUX3rqqytbr
dsOY+Gtgss/e1uZj1rWb+iE7vIy5ElzhzjcgO0xtM9adEsIi3FTcCxOBU+BS
a3Cb/IwPaO/oGK2pMWOo7W/QTSFmF92MYJbzGQYAH3WDyUnuWcUEJQ92W3Mr
/+ptKy63iJttVtPbP6mSBDyYUXEWYeea7/SQ9JXViqjLbtrj7gV2QY04X2y4
vIsJ5A0W0OtgPSEVUupLwbzgGEU0NqUJdwisK/kq4WQwTnhesT9rSWX3kVtD
f3wBLTVmxbdWBDBLU9HQXnSIiOnam62NrtNebFaagGa3jSnD5GBblK3wwODK
0W6uAelwej1o4D5xjxMhbO99qPmOnp0l4RJapoO6HJqQx+EfnDA14ohuAI5m
zvsrmrXgVXZfLsocFSTuTxdFVreegkUb1V4rW6dVpZKZM+akcNOL7jhSaaIN
mQQASjgbcpekND81PDc01Ex8CUdchXsVooUkwUZD7Xw3bMYTBnFrKiyBmdbJ
IMAfKBC7NJ/hIre2gPHd791tPStMkdwnMOB4gJ3EVZ41AaNek5lDlZzBKryY
FWQ62gDS1RyqDdeGCM5m3Uc9sh9Cd1D7YeF3rcpxoFRhgWJiLBQgGOdUu2+P
UgURzlBXZy+dNOUj9eivqHYrqdTOBvKTADidp+C+p98WZc/9OOHQk5Lxf3ct
8wqrAzaNSiFUFfaMUnTjPcrjiffJsk2q3ow/zFCapQPfPBfmm/+9FRl7Bi1D
ekKVB02+/exj4rMN5xG03bZlp7YhBGJOJhPJNGkOHFSU9fmab1yaLSINN7/P
Z58VGRid++pjsE1v1iRfjOhY5xalCVdQnAlxRzfsueumQexiOb2fjN4DxgJ8
WtEi/DL+QSPYKOYWex52DnafGKWBkCsQaMYvVjiIMXDca6qEtLZQ7KryOUam
hHjigkuRvNgltw6Lo2Ogd6EThqbLwEq9+3yUtACjRP64R3wnha691efEtJXH
B7ZdETgHKBhfQ3klG0MitkFc/17I8wc+kMwcR+4aUuBjYlgk5y5Tcx8Ko1Qq
A0DsHQkVSBas6fPuwBCC/KAJx4akasnjZoJPh41DUrXxz7NlCk20VOKKx13L
n7BR/6+fcmJWZC/6co28qGbpbiB/Jro6D9e3FMd5wLFKN6/76Fu5GS8UgYDn
8uW5ox5GUxffDQeexJPvLN5pVrXpAui1A9U5z0JU+MwMIulBn5LilsNE+nVr
OuMx8Y8iVCJfqo+RNvDLAr6RbV3d6yW+zh74q+jC33flRljsO5CeBUPrYfc5
vtSEyyGWMmPWXkItsJkzZ1JtlRu7hGRPIMnl86AKOQeEHaNbcyDMNCE/b+xw
TS8Z6Lu8SRxTrxeVrsF5rLB3xOQUSDuFzG1L8KWknr4zICk7G3SoypR5g2fa
juZsbCyCzbYPWhYP3M1fJsKr2aLySGzQLzSHRccLynhy48a6Ne3+ndqjArxv
enYiRomQRMNPsXn88yR6R/9XMyRMv4YwMkx/OC4aOAFn4Mwc/VlENtFwQurb
VH+ZXa/EXeGv/pYTjSL5irIDiNwP6OtLJLgjvfPCYWCVBzaX7gY4OWH4pk43
NzcjPpmypLzr6b6aikD31K6y9bh86woCxPpVlDXMhIOb7qXvkLO2Y8fpRbnQ
TR/dhj40OkYHgNjG66OFTBSB/SvjvA/UdaMvw6e/EYa4+3BTDk0eRM2kC6YM
RkIiNMiV0sKlfy8XdJ2YoQ/iDKWErRX1JKNNRADU7oUlPVWRhiB16XjG2sXk
7a9+egug8W7MuQCanRnqa6sZi15ercALLhTpeSUs7aqoKHhQqIFRa5i3euFS
UegGAxAiBKtqZSFVl2uTnYEFVEANJSRpC7NM51rmbRXWo+2K5iabUWNcX+w1
Kwv1uN0R8N7I6WBfYuAv+5VdwOm6WO5LqHQSKNnAzUUdGXtMs0PRIjLZtHUM
19qdKSaEAsE4P7alS3cQFXmYlJ/CMLcIiWrFAKh8+zLLihihBwdkZic6JaK8
pBJCyTT5dNb0/RhAHcOOOQwJsJHqwNjDikOOgPDQkEcUzianXpK0rB2QXcJo
yC4SvMR1ULD6J9GB5o3agP0aOmXNmMyPVGM2Mxi6002u3kCpcMV272zvIlQG
C9BorEDEq1hITJtXtSLf8aZIPurfltyuV9H1mI2tgrk/99koqPERf6hkUFG8
H4azwXnAbVisW+Y44fplCofv8Nyp9wddRtelnwFMnaTCSOsjYEoPSd2LL18H
JbXR01oJzAlzCpaUGdo4BFb+lBsmvDfV+4bfzcLZJbUPMGlkwwOCnQbgCPfN
kYp7Aji86D+Q5ng5V9VmsoMNv0Nt263exe3dGbR50GP+jlYnyGZ6vKoup7KZ
7to8pN+4J44TIGq0t+cNgWULRSAAkCE/uCDYDtCOURlL3WSSWGtyWOuakh3w
hmoqEYtmgzkl615173l/TGe0lDP9btyUxmf5hNFOwvxqjXkT5D37R4GUKvOB
+/Esgkia71uccl/cYRdlsxDyJzPvB3HKEsr//BM3GaBni6xk+2xslv3nKdR9
wUX/QuCH2P5itSOeboDVPEhy34+2sJZBDt+4cAq/nBcQKAbQrNteDrQ5my5H
f/Fi9bIJXdChXBPtO6OSU3FAZQ16XbPtS3cZN/0YvWu2XoqYx6C74+f9J4Yi
Uq0tsWRdGDPbCzJc0rS5UZqACyFgicbGE5/u9yyB6uYQ8N1CUpsqcsdbmIvO
9t2jtCdtWd7+8VkxsQzpXEsBr/jZsJXz4V+KIj2axipp3RqW5v3f0xWmxQZe
1AOd8njHsT6Euh4FXcYiuQpjbqwX7qAGXiXfYFbpSiZx7pzVTL1hL193hh0n
/aTCQLvHfC1rKEcM2yrBrzba/q9xB0E4fjNgbh9g7EQMSbkgjgevCeyt/v3h
adKDanwvaad7+XMQClPeR1RpMsOLK0McIcp60B2ByOB3vobLGLeT/naTzkSK
FC/Wr1YhSwOdk+D4RdoDpa6IftBoW0zBBs/bv5sy3pOGsur4BONQlla3rckT
g7k92iFXonLMdygG3cCe2a0sxGVx5qS1Ak/whg+E0gvkQGLFXcYr9UMU0Djm
AH2WURD0vOarb38mSMv/znPFt85yp6YIg98Hq5kItmo0CFcaBWZTxBkanpMo
ouheXKrDa6F+6h3M2itikge4Jac3W01fJ9iW2p7B8g0jqIjSqaCdL+KsfIu7
jpPETq77hCb/b0Xzjq+CqGYLzj2G4mKFlBgcDPekIACB2Dqcb0/HiGE6NaGF
VbA+xU6RxmHa20DW7Tq/jUFoZxyZlIlnXuVVfsgNsyyWSB03xuVcp/STb50y
vDlE1p7l9OZAToDQ1blEFaDiXrAIXRKYP7NIt4CmIH/HZESGzVNLyKsCxcNR
N1DblgSJ7lNhoGq3SpmH3kXTkgQKLLlD89b1qCjlih28Ph5sHNWl/zp9N2Wu
1EmXXlvh9a4ppvjPZB3n0XCWMBNxTCfLuT4Q7cbWrh2CfabdUydS8rS63Ccm
JC+vueQxk3/n4VkuHeDCYmDYcxfk6UXTGEDVQbDRKGNVbrhQPq5FS9mS2kO8
bh7U4X59i51i9cl02DB0xxQUvRHsWzy/MFhoDgz47sHpGk+l9NpqTyyPcjnS
fdOvNsu1msQL6z1l0q/xXuja85vcJhU5ZsPvHPxl3X1oqztVCjKB90ZtQ2p6
3V6mG57VTRU4zykyvRjNJ44HkMHXW0xAnRCnSRqPaKk3tRbnLOtU9LAGtRNF
cP7lyRJxM+zFxH+Bh4QrzdGguY28wqBYNNprHGyU34TWvePo3r3hApcNU8YO
4/Y/lDIcNEObt4FPHtDwss3jfTzLILpQpxw5rjPiU9mKhjTtWJVo90DqpPx8
6+egFwYC55e5Md7dDCB95xYM09ZgyKXmovUX7VBuNuLpDGR5zdRRTKjQT1Oi
bB/uCkhB6QEpqfanaeBRJTjK9NLgGxNheVVyUXfBoElrwAYVYHYSTxfvavHz
3HnWyqHEndI2te99s9iyHC8r/QVbLxqqJIJs+Cqdq30/OTqM07Ja0LUebI6U
M31GMhNumJpznEmgE/ZU/yYbqZCGetPSqrLznWD4ajxZ98D6Qxq99Bg0s93F
je2cIXwKkq1NDnXFwL9kgGoB4C1TJHmAjPHeh9AYLHW7yk9SYxtLv/tiqeZ2
tiDAteAIo6KjERKer5Q0c9boQ9p3lpQLwwFqeAyyg2LXmjF0N2E7jCudIXsO
B6JxMVEN2BEMOUKd3hJ8A2mGy4XsXB+XVR4NrQlFBQE08/cVlh4TBAdLYqKc
ScZoYdHpcvAxQlT/PjbJRt+wv3eeHghBHn3wdAYyojKKZb9dWajKq/gaw/Tx
iLyMMIBvPuMDEIH8U77m/qQkkIENqXLNFlFU9p8pI/R0cVoMTyCMH3/mmZBC
9qC+EM4yB1zawwxXb1jKCsdbskXNUvXcyUiS2HLAbbxDRTtRgCwL3Qvo87tn
JPT3pRarA9MVgzDnj6qCwhMQ6nt9rrG1aC0dRI1qAfITR61AuO7fB7X6LIWp
WgXE0Ze9oqoskHS9q24gCQFJkKTMUBA4N9D2iTnvDFRgxsqvllAE9gdRAvqi
CPbNyp5Ibj0OVym66r8Js9lsWgkDuPUVmEkNHoRsPhHabqauBzzzkJd0oQr0
XMYyV3hDk0PzfGvvOMFbS42oPiw3A2PqUERLaNm7VMLY5793gl6VzbvL0ABr
fPVlxeG7z8cCmSW5Oj/OEovSh17qHEcwfVNquia5nPTGks8srW8zpIoWlgWR
3tuklrTAsWA1cTCWz0CvpzXA7YVfZjINe7/rK48UKHduVeRNNg/HF5RE/K3b
t0k+6NVDfkGVp2pNv/ZNrDGhxFbxi4FKdgEueLHdw780AVxdV/6hbejQf1al
jYlIZzwFBr4bU9Xq06J7SqTYpYkKgOvFbRnUBCin9C1DBw9QW5LAYSY8cRhz
8k5//EGgO4Oc+iTNaOCSIfm10JcGm987UScac8/yVE3pSWQGGNIvdJBTcSps
AryY+JZYhAYjG+IWa+cts51SjCD1312Yy9PXIm9JO7iGO+tGJcTvPijPrGk4
LV+FzNWv5FnfthWZzF7dblU53IJbqUhOLjeLniSphqGLM8a/FuMSWIJluKKQ
oEniZKkRevTA+DmXgCsloKFeGh38Kkk6zjyjvuFe0OO+03teFdaBgafHOB4/
6hNWGBmGkM6vVtCXml2rWtoYJFtqGSzHRWFa326FkpJyxHWBAIoZHAK7hTnm
dndYvY8sMKNQ3zkWslJdJniIkcwrL1GkhevZeGUPIbcAVNBR6CVDplFYul0n
HshWtU0Au4eIQxPJBknyLgS0z/lW8oRvNH1XYROoLt8+FstR36UkcpRSaG0z
0yz+/L7eSIPFpxB4Gix2L8dJne4xBUOkwpLkJSWasr1ELWebxbQADMvEaKrj
V2QVtGsHfJq+cdxpiG4/knZPx0rHjzoHh3dwmm49fOuGau3gH1QImShW7FF5
Lfdw6r5d+CLMtY1SeUax8RAFc9BUNm+fbcF0kmImr0ekX4FPuHLd0TAUBFCC
jW+BgKs+rN7F5b7h6sQecAoC8AEBLpQUtTRfp8vTsg7vzITkKqyKeJNyEMp9
zW8EXIB0Pj0gPr2Yg8S/a+GTKe/umvvXmlSUV5T3wiCSAlBdYhZ31YNfol0X
CzRrV0iVTbWa5GYBfYipqGPeF1wKi3S/9EqU8BKkhHMwJrRE60o2rnIQoCSC
sLoZmhX3UwDgwvLvK2iL1+bOe2igQGWdeeZ0+4B0ArbTvIdseIZ4yuNzKPcF
2GSScJ+ZeyYnyV8paYQJtwHcuO3SalIytDHRmW/IZUomSYHH5TEDKFcWGOmX
wRI/0miFqZmKDOAxJ9QPhh6HhGhu0DlaJ/4COlULfTPEtkWMFJ/94/TjDpW+
DETL5jVNmPehdRr3Bxd4J3KEULQuFBCrTsv/tpn5QBSr/8sWmQKmvHI3RtdM
GK9mKiEnsLpQEFTkg01hi718NU2TymWiZwOwZMqeGMpDIK2yNRwAYRjoXx9e
z8OzFAFUcYyNjxpJgM5tMaaUA09EpmqOnUgIEPq7L7ChF/pfczqG85L5YFyA
k5EWkO85K5aW9faZnt+lDLyLAKvAaOsMx+n1ilD4So7jxLuOvGUQkach1ysw
CbaZ5So/oBQaVDGgXuWtXguubLWdFLVcwLyOYXGGSjewEwoFgmrHO9TdUY/F
xyRBEbgnOhOxyqaJ3K+yqZRPmDIS78qJMD72y/2MfMaIL0Qh6YlScxT90whJ
8iMpXA+tl852KtdOY4fbG1Ax43G5IpodI71Jx5C0CIUTIvQxVHtuXrATK63Q
YL+WZd3kMufhycuddnUxDqlJbSQxFX6axj+Ull/WL+9/j0ohjqIfUnWtMsz+
lfmhhoq7GweqgYf4Ik0OLKOMX5q8xB2Iby/3VxZD1v9uYoi3HHcoVGUt5e2A
Y70qaRbqPbQVGtAxojeLmiW26GLZ85+7xq+N6PfAj9FTH77BYWZ0B4A5zo9R
JJA8qerofGykMhpfxA1SgZREt4x/tMVA9oYczSWwCY4sBszFxKnytllLohFX
s4iy5NNEqWcYdRm59BMTlSpLRnKoWuAm7Dmd+DMuvI7LbuPn/uxiR23G1bpI
6Ln/mLF9DHYF51Cx8I0Gj3dhOxpbL+ZgCXiunXg/PakNUeNkzjxDdJu91tHn
BWZoYH72sY6xBeUD3ngjoMLp8aAwryrIDbHN2L0ke8BWAeLs/TEtfXW77qiT
6CQiQ4lOjp0d9MT0oWAjyQErRA9N/H7KyBH3VEIZr4y1TE4LkkJeSkOIalEl
PGrvnxUOXdtbELptWaCRrQlJNIFVfVrUNeu5FlGjOrz5FkzlhUqAw+tTRlMf
mW7WzDLR1ZfLSEUreSNH53FC57QwedEGdAECVqyvPPpfPVtDsHGO+Tzx+b+1
YEeHyHhJ5juxvDeMb2/DNLf1e3RsJLHwYefCM/tS2bOM0Lr6dP8+B1Q1pA/y
enRBYcPMcONU7gjzT00ksum/VTZw16s/anCNFVc2MCMX/wxSEjgUSdIoWyXa
7aQOyH2DEr2XzGe6XAcxhvVuEBKa/jkhYFDi6bGbtMyW96VimN3vOQQI+MNl
OAGheIWkQwbuKKqCFj5mM0NzUsGfk0uPBptD5EiQa2JlBlZRw+VZjgmAsNZX
TJu456TFZthHzvsfXXJwnjbRFpRsSLAkn7v0uynlzc7k//ayW6uJ/uXfp+VF
ZBEASxSLMBYoedBKmXQfSyedOsN6PfjCIduAdwWcQudZMZGXZPX/KlNUYq1n
7Ct2qYNVCb2VjliHoiOT/SDnKo9G/7P3VS49//k1wRuPshnt1D8g6qdK8Z3m
gONCJSxFaS8L2X8hwQXU+0flaHo586iau9BQYmHYikR/Y9kg8DRS1NW84p06
f94mWUnU5Ohl/GqWNGkRyxiYgblvLcAORggneJQA23/t+UgK16+siI0k1668
opXGTGsBwU7FaEWNvmlpFbDCEzazbULj0lNbszQr/TtKyVqpDTZBeAWiYVV5
0tVOcVCXsfAjFIVrpJc5R/tQJXw3fecRph+24NO2lizGCX/90ZuUmIOIgQTr
8Ns1i+EGMvT1AwM08m6QYC0W/+YvvbLdgudf+LzRxA3lApHne1F0yULFwRiT
HFHMww+Jm2kausanRjqJE4dtfQFc5oDgj5Q+Ofom8wS8TzGIByHDrdullvRH
0yFbqEsYqKl6va+S7aeYgUla2Q9GdRVMXWgoxbUKd3rBFhQwJC8suG1QRFa7
5swdpBjI3JtBkXQGjq1U/Kex+omWSdeCKdoO4cSqXbNIdj5KF29TuWDwiK9H
ZXNH0yQVgTW4dOViFs+LyQt5lOTcKDCqaxmwNg18EJFSrorTYO8vMF08Oncy
aaCpcIg2Ec6u/fTtMOAS+mL4pBDbxAKRmOdi7UygSgUiAileIb0TskdF+Upf
pjxIGVqhbhPGJtUNdYQf7TQ+J3Qbz5t4AgPSjeL3+4xeb9NBiJ2G4tiQU2Af
N4heLQJtRtwPcUJwQgp2Urxd6k7yeSk+5+N0BIEWOrA+rTgLr8CS9SITruOr
dE2a6G75mTSIhelUHK1xNf/+sYSxaJenkJGo3wFRCUMiDeGAwlKPepZfcIof
gcPsXCN1ZMW7gZittEByOAibg/XXylUtoEFZ0LYJoZ+9gmoTRb0LHynmlY/K
Vqo+IvAfBLT1vQeT/x6feVhEqR/raIIqwQY8BgzjiYgcNzQrXW1/xnUe1EiT
SslB2/CGteauipO9pdRf+wMoviBxO3UL+1iJWEYeKb5Xo9ENHSO/9VhZ3ZYB
vIE2NfE19yA9AIkjcNvE9GAwxZaUldOo2xRwNMpZKwx3DDOvDjh6sTGbdtW4
dJy34CAirAbFdFsAk4JyMFwRnJh3IF9qtpwoyc2kUqtRDDUvAZ9SsGMqizp0
TIFFSKJEtyQd2F20WcXFB7MIAyhzYtN1p8OdJt57kQ8ektvUKlQa2O8GiDva
WvLp/3n8WtKEbFhchLAywF1tT868ZpvfW8sP9ymaTMDhxt2ji9QxsK6RNTRI
EgAZgUS1VSIRRoB+I5R1JIhi47SgHpG7FgFrVyE+8ys8G5BKMpWhCgT3oVUV
AfILSNiNuaMxSQJhMu60MQcNUjkg7lsE7Lru5+Iq11fAYQ/vh/zCKg+kT76x
eGCNaaJ9ZrLabvMHRd61S7zkI5QzwCjTPmGMdWQdEoNQg8Zpvg6hAPFPzuhW
m1Ztna4Khcm75HIQ/qsfKzLe78N+YtggH5oeIhN5aWKTUsZBwMmD551VdhDg
B5BrBkIpfcldWlSzmQmoa8pfy3s9wO0f5CfS3ZRMk4dcSrqznsdTj98i8Mo6
gRM2KJCcX3D6l8jb1fJbsyP8Zo8cWB7on2tnuPqJxJFgQUTZabtownpnoiEG
Xi/ax58mw0CDJVVkHGl+2WpZM+8C/BSdKEcamZ4yksDsSzoAfal0aWH8ePV2
dMQeQGcpZXC32pZMbUDLF8lxT8jzwueM4kRIBlB92pqf2oQ+IXY59gDwxwB2
Akh9B9Kz5DjBeN9Lb3YZzVt4YODIRcDSPQLBeQ4OoPCYxmb69HWXeVqTcH9X
EuvW9zfukFibof73ipjYIT+MMNwfesYGCeYFlPQ6V4LlB8aX8CVkUpXa8Xhf
SFHpt12sPTFYKAC+cNKJXIqYBom632Md8v9wp5AxYoYIBtWBpmFyTQC3qrzE
YkO2v974GJ7clzEDlNsMiSNcyOt3X54XXdUGLormx/Yy9EF/yfpAMcvNxomM
au3f8Swx0OqDYzH/xTfxac6NKoNi5PZyhXl+oyMP78y7I1QAii8A5xCiNNmx
fQtZAg52YKgXA40mC0d46w/A6vN6+Ri+xk8JaZTEM8FXHu0gPnHCkALZYQsA
krSrcNZMq1jqE4+D1eQxSfp7raYOEqtrLmHNDtEVkV/0nRWX7f/NrgGD25iR
TVTMGXekG/w1URjsf9P7PM/L40YDtpgHzQan/Z8qB1cNQjEZsEtrW54CpTO+
QfHSFjsTiKv0lma9hVshekvl10EiVs5Q9PWTo0KuGLLE8CCSBlKN7nuZYJbe
5MYB5QjKwenbCbCHcjGEOcZef2Im1Tcfxq9G/gu6dN4q7Zp1whBx8uX8D2i3
wuHndSKI3egqXkVAZMNiGWHj1BELKVvTs7mVfLbY4a2wNAYs5m3LxId1nVEW
VzwzqYCcTWOwHTzMyDnaBYCyn2xaZUMi65Z3SXHmm3DhLXoKSS9A1HWtHEvH
F8M2fhPCiqBtrHYP24p3Fdlc0TAfXHK4+pikyu77KjsOiBP/sVTjOU+xG/47
EID4NKTyFh12hNKfUaYMvny1uPxeDDTVhELvYz7vOxYTnfPF38B3ECgHeJEh
ca74ogkK9Nm77CZpPrwrL+ht72+DJ3LF/5f4KihabDiYK45Sh+msL9alPrT4
BSCCZfvqrkAfm7l+XwlUuHjmqIo41urjjdKCZQGmB5/tG4bZsftZdrffXCSd
iX6UlsIAm4pHDUodi3kSKp70zsQgUDJHFVd+VAhTZkd+exgFUq0ncoiSqJVc
hFO+ftPlWBYpctHC8QBb6QG/uxhni9AQVa5wV/OJmaV7t4wnXopbG/SRtSvT
OklDRHByQn6B0p6scExZuLqco3lYSDrR2/sA4M8Yi1Z8gDasWVxdUNnIyrXU
QJdUQ9m+38V6oUQL3NV5SMKiX6FZyBTQ4xpQQcYo++i9n1gMrSFS6MbfjZUQ
Tbeato+0pB3hsUGn/uk2zhE78tZX8mZuECgu8K0OUMS9WQmYeAKH957OC3jV
Kq1S0nov8zB90i+RPti7pry4ycjzudQRyhoeg7TFFNqx3dvoo2HpN28mAejC
MMDFaFw+RdpAiCAVAcKDPecwGlHuyIOBwqCmnUu82TGWAWKZ+RAtzkSJwAzd
GxMCaYPRxed0kxDFqgh9qRB+ceCJ1xMBsPQkAhyz6fgdRT8l+3PWK6GDOtIc
PRbtOu6zs86n7SoBYwwjxa0rfyp6QuThwOYqHYy6u+vjQCc4PbxhZwSECi5j
F7Hsd1qh9+TB0gNYohc+xlXWRMfZQNge+l1T4HLDgUMRXX7L05PL+DfIqzjV
gTRFismtv1NRCFGu4avHN8nA2cwy18YCY9egAurXNtj/mp7R2BH7xds4+S6p
/v/XKIWh8M7rpCqACXxLHhvsKQMqVcYSuTnBWHT4uOy63U+f4slQBhqXkd0C
2U53k/Js4Lg98p303AqXxLz3TMG52HzWOAu6FM4VDpYw/6Kh33VZZXeqSiUJ
DR/rIekescGQ3CpfpYJ36MuqkQlB3zjVSDT5vONeunW9/0jOhQYZx6V+1BRq
3BhJZVQVmwbwgQ8CVDcoRuhJpppoXo43FNR+iHG1VAq4HuFw50PTX2TL3MWr
9ysXJGfUBT6sl3i6TkygiKQh0qVwYgoQlrONFI4zP5AJ0dwYoZ73Y6o6pvqc
QI5NB5gwb0SM9ERIigzhqcfZJwywLX+9oFWQShnCGfeNUYBW4ls8JdRw1K+G
PW+xXMSM/f51lAsH/COHgAi7QI1FbgD9JOUlN9hjLPBLV2ppC8zmyEBYlAaY
OKF8SqB+ry1hAlrnDUmCI4m539xRMAsZQQVqhgR1HHVu8MiLC6+YUty6SC+H
NIY33femHnnWP2W0oUQL4xQUntd4tz/aF/gJYK+5JxszD5WH8MV1/XsofXok
E3i/yxks/8jH6QtrNYZQVs76WJARq3lk4KK7mH1JmY9l8/oDmIKo4d8MsZph
Kajdfn0fSD/oB1agEWK2AwQjXirF6XfE0YbLqNcL841UTCIxOHrcXKC8y73u
MwgvbhRhQniWidy1nwWh1/cENcueHLKuFKBb8WoGeBFzv48wzERof3HeXV+q
mRuaWhTjeaAQpanvBW17VINZZmGfE2TOBQsnEm4+7PM+uayTYTK/4TYgYXsD
9aytYSadFHQd3NjMeEQjrqHbeykLB0HGFBg1VnApbhDcApsYA5OtKzeOdvV4
ZYKASPcJsWtinTmwun3mTe3TL5zO9gJO+udR50wMMLBWcqvwmnCuOIyXcklQ
Xe50X2kjzKXZarG56PlV+KB9OaRzGe7lN/O/2r9kXHmzr79NaSYZOsH7FOmt
UIvsMD8OCBPvwe+sH+aMNmipB/tQDxqeGFjB/cWR+g6mMrrzQDBQoQsfSpDT
EwiWJnegUqWO3ZBaXuWjMAQlTrlJTI1bln/lPykSk57p9kVd4vaAYI7RzwhY
lM9oahKcn2wC3GtUDqqUTugs17t7vodxKuedYUTD1cghYDq3UHRvabbq1qIk
Baec+BcKT/qv4JhKjpRsRNx5DRD5SuPxh+BSAlOG/p7ijzW02vC7b65XpiAG
jeqibYzQuy9iAUVV5JpLJVkTvP7mGEiM59bN9SJ1dF1KxsQCBY4sWAdSD6dd
nfY/ger8uik2imf/14t5FOtaCZWrHLDAt2QMBEeRgRoETIIaE4KaqWqn9es3
aIv5hQnbXT5S8Ae9snpqCw5fYfF6gqtQHP4TdeJZSghsjfUO/tWhWV3fZJEB
sEz/2iFGooYFcTUrXVekuC/LTiwqEsaKg207FKa9S88OWCxwZSyDRGLeQSOw
ealSuSU1n+bWcLfvdV1kXOyA3AVQyXr6O3tFvsQ0ffi5IWUyGgj7gFRC/23r
oeEbWpQY/hEdRxayLvGqN2Jl209Oo7KWa5t2bUnSrDOT8xB5cl0TPydawBkd
JEV+Ot4f/WlsT4049vlBmDVZDwbMl1kbE2sD8whFyz9RsYu/LHlpwsk6hItj
XlnFJnp9yV2onsswDyC2Q9ye1LJ3Zum6mt1MwEGOq+e+uC24qIoEOJR1qKJG
UOBIZyzqLT+qTN3cbxxrme1wWPx/qHeQnYeZJfNF4ldIhN6WsGoSpqyd77H1
9g8JBVa7LWirvak/4bmUSZw0jzwbtNs5bDIVuz+FQ6nXp3a0iEkC/xjQd1Tf
Yl/3U0dRBlwrZhFAPEQOdZsPqBINMrhv9zw1WyKSv/+43ANTj7FF7mxjyxzU
uzFI3KwWVbdaE0UBMgiEFbkkN5zQ8s1XmcRalYSifQ3FybtKTBAgXucamse2
g2uVxgAmPUgJBRXuyE/244heVVEVfTj9VuN+hU8IzKkMtAyvBfH1T01iFj61
ysz8zJhBhDdnemgTsnvoge0gJ4lCceVd/mWLtQFKjfYqgrAits37oQyqmAwE
scexTN51u1t665SdjcInfRnzkn/GhwnWgBMd8Mig97JP9IX3C/Qh5N7YQKEv
FJtD2Q+zPhFqpxCJSv6QG1k2EcXMaf6CeCnZ3MG+TFlplVLuoNqIX7kFhPco
FVtbikutuOWdf4wRRacF3Rxo3lT7juHyta+qDEJMbY5SM55QSjKwXcgzHibp
5xx6HxLMXNShSr7fbEx97O1HwM5pKlXWI8VfdECKOo7RusCKW1YIrUuzohyH
fc+9TmalmZWEnlGa7JRp6BS+JXQEH0AWaq00YNqenL5lgG/odZh8iu4CPLCF
lzvPzbjhtNeAmQijK5agwqMuaU9MuUUcJHRNOS9baUyjuRhuK493CDvqPtDP
rwVoQopeKbgZes1tnekgddQMsntBHN1s21SYBEfcx75VD84BKNSN9w8SoSHn
tiFk76E6V3QJ0doy8UADE3WHSmc1sObGu8CrLVXKHK0pFscKqAnl+wla0vXQ
GyQvSOWloDBSxrciieuHbGTrdACEv+3fjpwdfLb0P3lbJhyYyIiPsFE0HV/0
94ckRnaKahOH50iDjou72Uywgd9UdTPQt3Ap+hwpenblA7kGPD/5YzV2tiNV
+kKC5nvPpnO7apTc8j863BElOcWCRSeFRP3cQyGugg14pLh1eX3+A+aQvXku
dqy51rT3T8WQrzVhVEjflqpjYxrK3gG85A/reXWUPdXW/xELDfjCcoYLxq4+
lZt8TXeZdMUTYS4rkngVEi9HExL+9XCgpWayYd0+zZg1pm+VWMgLcry9CGrM
ltsQ30YlDO1rM2WmJhqQc5RAqHsson/zAM13Rl8CThjGxxjdxsqOIFUzUYWd
fs9h2OJLrtB587wums6BukZwwtDRwnX6Dk9qe9ruAiDCgJk6urrRBM0WU+ng
SphgsiG5SJpAcgUJ3kk/azNtVtZPbroMbne6CLptknZ8wkPGFRy9kZae1Ynk
VtGd8dOKMzE46LrSWRol2tOpKIhn0L4YGEYmll5A1Gd3e1CqywflbxXkyld8
7DMtUUNxOuzwrtCJK70CB3mFWuY+QAdLgXg3z52KhPjMmaNr/bKvDyyO7pTP
uXkKtCMihkTlj2Ae88PRKp02ZLHXRoNyCLM4vPKdHjPzerQkl1NVHbL/FINR
/RB2c2+XLBpMR4eraMNAqpt6lPGEbDk1Tt9XeWsaB12X6mI/0QaCCvksxB3S
dVBL/EUGG6Ocrc+9ZtCZ7G1w9GLcXEEL/OCgWVyprcK9Hn9y5QmuEl1cshOc
e1s2t0Ds/rN9MQ7PmHxYonPJUyK5+WebBYyyNwfC2WAHgCv+Eg3s4KWgMcAK
BybjHbiEa61UB43SGEl2nOoJcsIB73GRUYRXw9Zukgut4eJRme2r78Un4EoG
6O2IE7AQ2xs65jXt23CQb6DwFqKr9nXnLU+MfaNfHohMO9O5BQmi2u9R/csk
UjeoHM5jlR4T/14MZ+n7uwDh+DkIEHlOhZiyK9BR9i59zJvHIV5TFK5QsXF0
uUogXZxmsBluBYYJfPQ7npcrFArQ4SGvs8zpdLM9q4a9rYxuwyjumU52CpNe
UbUzVsfdrG42J6NY2e4ZJHGUpjC8NAl2Pec1NZVsAJBd4bIhho9d60yjn0hk
z0JSOTNfOwYIdBj1LL/FCrIjIXEsp4HwRn9y54OC6tW5Ml9PgGlL5t/0bWWm
2TAyoGtV1G+Pg6r5X7JrdAPeHDUeEkFwT05kTO5Xfj8/Grlt6EKueRurgAjT
bDsaMXGuQkY/sznx3J1TjimKBG6o8UjNN4Og5+zwrNdrJonbR9UbsauHHQym
ykhVNePTtU6BixtsGku/k4Tr+nkIsHO31PaIe6cAY13KP7Yfsip7KZMnCpBd
4dhtnBPsQDkTzBLY6sHHhAE2UkgAstYcin0ISvH3SYHWLBbl+OxNnUf4ZKVj
bnDJQUXvHLFgQVxo1HstpJyWamh8F656HIzmlNggSKeuvlXfU2SDUTPDxqe6
7dkFRxwBW6Zif6+Q6eiNvh0VTzMxU3c2ABb0/npn2JCAeQw+v0Oa0d9XKh/f
IPLDv1BcHZLwLOgWV9/D3o0XF4ler/tSVq95/St7JUCAmcehgUJk+ttJArBL
6dwFL/de1rpbC75fSb2C6bdNqWw6lZex+aWBDxCv51yBfDckJ49Lk9xkOHcM
epMiuGUjLC+b8SodqxOQ88cWFVjEjFcUd2LAQZnKH9Xlr2iE/7lu2t4n1c7L
hfjbsikHq1SgqVZpBZOso8zsqeJrB2+Qkwy7PFiiTRYPiNNjFNaHskXJzDwk
LMafFBie6dhWD5VFaGZnIht5QaxgRcCZGklqqbGv2QknFS0Z+lavXfvtYpQ3
prUxfQYjkOes31BuDUxMVHoCNl+kMSDtxShtDCEUrtZJD4cGwOzhQtjrD2vT
DatxqleaXM2eYlhl4YzfY9QUlHRWkMijO3zZRzozRBJJiMPS6kRles9Ye608
udJqV6Vz1nIpiuPLcikADdVukkE6iAWKJR83jb+NAqXYFr1+wWnPyqjZyDTJ
IVqfK6NwPRIOKiSogndc2FcLipFjkM7L/UCUiFck5ku7lLRxuWRray9LZ+5h
BviZu+E01yKabk2CvQuo3nT5ZWQ1rJX3T1YLj5BpXHp+jRrAhryWa90SXQMk
8sN7II6tU1M92SFJyAQ4/DjCd3onsCpKdVlI8nd1fxLuaXk/XIc6nbGFoGYQ
1aDQkJvcy31e44BPB7ZHE+KZk+qHRYZH+O0YJQKK5pkPy4tcLmgAQxjdGDLU
j/CXcSnZlMxNRVFlODAT5a7SF4vxjdrv6pCb2f2kHG0de21hr9Dz61qjp1r7
PZwNQPrbvT3MKZCmAt+2NAyvr3en/P6qXjYYG6xeTmobjYeEqQWdpZtZN2sX
Y0ebSNWl3XlWNaC4+J7BFtGkhpwD5SQ2XqcPV72HQciGaPZBb7qkLTrTSlP9
PgJr9n2gEcwyhT1KbSWfwA80+As5PS9P6633k0wNiO+w17d4xDvkPCzBpkp9
mvPFUcVABph6LHfBJ0zWSHV9Vm+jkFnufoTdbMr9GUBcH8OdwXRgY2WgtcUV
T81/Gf7vFkNQDwiW85a98cLl3b06/97nYXPymZd50xtyeijcAaZ00qDX8FZj
sR2CQ+mkq4ZJq/5XSPvZZjleTEcLdnH6XvEBrG0EPdL7/BF69jkWmrcQbtMT
A0pHmKSODkgs2GADU/lDgz74IrCm+/EqLJwjyWABA3m+t0twK+tYYb9aQv/p
4WWIwUtjtKYtPfV01zmyMLkCb693HduPcasu672q17wvRS9CUxCm/+kiwqaS
AM1cXWLnlJuD7Qw+LIEBBF0N7OtwiV7bkKZkuFtEU9WA2m/7b+9vL0DuDNU/
Tel7m5VH2BCHQccSR5KrQroqhNYCNguqqeMWLvMJNcA4AwtoCoouqYCDkLD6
sqnAEHIAzHSnLJaSrEpLmiZDrxlKR+BpKPGLu6FMAVBfbewLr3+LwJmGzmZE
w7OVW0gUZ9B2J2ilVrHd0/OaqVQn9TVFfSBwALHC6+KoK8XhxP/smyrhIxPy
fqBwv7ykEzwMBFLJNB2ZaMrXOmhf3SF3d5douOzWuVj9+1+CMyfJEtT2eXKV
MtqJMkir+UoId3DICjFUjb+IW3fYSlLPxLQjnNZ4AkeYOovo2tvovzOmR7ys
ITG02zXF5LeNahopYnlph4RaN4goB+BHgWEkfejHgJbixiGs1fsrlxQyq7Xo
Oprsfikk7pwNXlZifhOv6aceURXVaKr77/2y8mFb3W4hoOHGpm3pYsB5EAwp
NMkBrq5olH6a4FTqL5P3fF8euemcc8MS43xQVJjihA4EOCeJ790VAWhRf2oP
ZV+vH4EcuzUHv7cNsuL1KZRMCBNRTwoj7SSygyGY9l9CM0deq/Ttc0ncFq0H
LYqZbFORk+eEcvFMQ+vAjeepdfmj0DT2o7guwxMTgN5OfGRXEyZeWTkiVlJI
Hza+BINK+ZcR46PZpMSDdzvOh0XwzL+e/DZCZxys2qUAiZs9Dn04L/T/dvue
D53FWfQL1A+nkHgqRlJKVLl+9/RopQ9juPNOk+6WRUh4VOkJkwi5nDEfo+0Y
S578TfQ83ni5Cuql5fXwOXIdF4vr6qv7VZEHzYPaeEpQ8LgeFxwdPkwh6c9a
bBMFAO7yERS2NHAuQAJvrmFx0JmbSI0M01oaDeUSlc8Qb96BHhPPqEhBYpPe
F+nTZYJsxCcqF7k2ygbwWhRXv+DQV4OQFYRGSWOKyaN6qlkAjjcG3plBUtWj
vYuLvK3sBATQWD+SesBlGcqdjVdvC/PeTu1rGeOC8Jtcz2k6MP+DkAabX/gz
gmLsY8ROoG+3Z+5BWyeX6HLfGTi7KGiGwd2JJJyMSm1q2Iqq0vxig7IJXzM9
Dk1vRssXeelzglxg00FrczI9yQf5YBNKTDYPWpTb5J7OUtSaCX04WJFdoCci
RRSpPG62ciA7Nre5uIL0WOmz/z0fOqwI3g8DxCbJ/XXYsgTOv/WBQmkqcVuc
ISjbykxbfONujg23O+41Fm77+McWRoms8ZlVo0SDhFQXS3PzHZ1SmG1c95Rk
srCn3MvcngTEaiTTDC5hTQFKAgU+gkbqB0dHJnVgbXfMNCitLK/rMq7l8aBJ
g7aM8+9qIMxH5zGjYowO/0RCzYwjiYLC84mK/USg0O6hdW9XrCHyt4ag0wfj
04cRLL6m7giZpYsNn1ODQqd0CUfhxSvKr+ZA3kvSX8x3c9Au7wgGhKDxG0MC
FbHHJV92SX/KThJziZG+H/bGOFF0JokQJRTLmXSA0S4hRSRJIKzRdBkrArbJ
sLnlhyaJ/urdGQaFc3+Vr50ubD7Poi+RchVdT83G+lZJdhXSosz4mo0pzD/J
HGcs0nQxYWnCy8bfqH0Yr5vp9Tb5e9pZSnJlnkGRXbjywggtW+njaGOdG1nj
AHkbZAYxf6ub24B6aICQ2nvMrEB9o6dOxmfw40E7mSkrHbaxt0BjM4bBXKvo
ncb7zpU8LGwA4MsGq/3VnqEeFy/uQm+FZO0UDV+mxeZvbVki0rySB0kHLEX7
47IUWJYslXukXzB1yL4bF568WCTevC1Q+NgsMo7+4zMGRAokZWoxYP3Of+Ex
QujkRtlmPxgEkA50Dcq5KRYj3mg1YGSj8PSzQbdgC+0O8W6wDxpqNm32wakq
ba/l7KtHkgHC3sETN1hJZ03JlUyn70L2E0VSUGYSFJXcGRkaNo6CPswohYhn
Cjl7xfLlLmhN92d7VqGDoKDm+H9OifhExf5Gi1Pm2xtdVgs8DU/HkOUkPMMp
/trnn3cyoitO8y6Tq5CAyJ+da8WfJa2+hEdGMYzaJIMaEhYuHPjQ2tQ1x/Rl
xlgcInlHbEseQ/F1EWRppeCcfMnUX/txW60JQS6qHYyjERO9oVMI9W4aObYj
bu5zDTvRtvqPLshzVURqAi+tlp5KZnm4gzLMAkO0WV8Tta5ZFI/CGKJV6f+L
cIy1J5Ik7VmfiWgkdehlvkH6s5Te+AOyicLYVE0KVErTrbVPMJFpDRsapFBs
phJTgwHtCBftUBfeJrmKytMPsm+qU/GDmTCWwb4PqXBfxSZh9zIjiti4rl71
Xp6OU9CUoEX2SuuMFPVsGrVg4lzuUQuB5WWFpcuiH5FtDVa5nNqnb6KC8f3J
1TjWwWMeZwkiiU2Gp6zTZpABNJga/mSpxk8v74XMCuYgBaONp7CfOeYFJSaI
FVCq0+eGfzy40anCSfVqkJWsF8PHR+HehBumkekaa7YJ4AUWxWwuxPEtkjtD
uO/kUxpIwMVPU3XBg2moRYzaPgknLsTo6Nw42/XTpG7zyjNnCERwmhUnYX0r
ax0oVFpwRCoRP1KHjdgrX1LzbHMi+9A0PMbHn6X/PVyEqzwVf18FAzpw5bNO
Cb4VuH24nTwzXAr/CUXg9u3uZKFBq0/rhb6Rp7IzH6rJKNQba3B3uMUFiQ+7
b+VbTJ05Nqx+bnuLS1mmMVhsySUnYtYbGDXaJOK7/XyUFJA4KSLbqRfvcggN
URjYoV7lyAOhVU0tEDLW78+8GRMlabgYwBwkk7cK9WgA5J81YgCu+Jr/bbCX
te6LCUBZBeWwZxNLwHNXbURDp9msmzvgZiPVTUUjzCahIxL/lR5bXOgZWFzB
ItDxi4teTTvoCowmwNpD00awJ1PDvU9hIsKaKcom4/zY85wijnbHW3SmQnDF
z0h2Feu2s8zpMi7i7WbYHz3G38dByztHfyT51rt1SmkU7varQejwCezovQFL
GdLI0h13fEyk9NOXyiSLOf+9snBRgFgQIG87KDRyWA/ji8EmAgfjSXz/XiMw
VsPxykRtlyOZC1n7RGPCYNF9GBdphDOXvf48T335NVjZZKvIytoBI/qFfnGQ
yWqrWPtpvy5aAIpHFHUdhG93zSTHLwV8cmbeP+htrvKWWqclLTU1ZCKHnQG7
G6GT+TYexlvjDXh8Awf+Q2YADuPHAf6H5OhWEpOAfC7B5yz/DftOYCVVmvJZ
A35hSXBTbP74rzwCLlzM6uk+XbCMFQxIiZl4OsPjaqzVGbRkBsKcTgFslIu6
IdfUwnwmbADp/DxeGH3zWMxWsXLYnOxyUKy28LohG9f8qeYoCvALdaECBK0v
J2OKiB13ah++ZARiGU56o65OULI77nZ7HqEUXYHVmzOjeaF+BL5M1WahI4+X
c5P/FIseKcvi8lSLEsuMw+5HYFK/W0JYpWHRVjnpJVXu9W3SlJz1T3wk8vt6
G1KicnKSMMNZCNK3xVPrhyQKauSTT/LQnh1mCL0UQvag3Sg/5ce9FrbdTSP+
iODAIxqVaGglPECwDeFWEazk/yLNbTpf9d0faf45MFZoLvNPw+Pu7nKSE7xH
YR81RjI2ei00GG//ySpOPXDudN5cDQXkm6kdJGtQVkdvDM6TY5w8crNT07ce
uWj1VLH0gx/AkrVMy4Lw+OqsQoM0wei82kRy7ZIL83SLovWNUjYHJ3a7n9F8
qoEvizmQGVn+hHZUTSTYJXLwkCVvUd8+F/AHbVdaYWoOk/mP0O07knE9rOQ1
CeTtT8oDxs7FEULFE9LEPk4NH8WPo0vREG+6dKyVMT41skqzCGy8nqrbbL1E
XN+UWU+VojtfxarDII5DDaWQSSoS31TpKQjYkvZ4eZ/uszGYmUg0sbYl64mS
5CyIbzMJrxE1G/AcYcWhV83YTlg7tD3FwBgfu2xMH/iNjDzvcTmtx7Zkce8Q
hMPXtXDHc0zMnJ1qtS5qp6e6V4/3y1wsGRbNmxm1WF3SsI+wr0vOvjFsAGpA
+wUYxuzzAx0WRMCXnSGe3VYcOn9bk+8IDyQMDlUzl8J4wFpb8MLzmEZa4fQf
681lRsdgdAqqSghNHZ43kJmgByZZX0o3MmbDD62SPGIHjhjJBO/0excdAkXV
VByK6H9FizJt3KPdAvwZVtloSDM+CoInSWUyxM8KBu82LzkAHzWi5wery23s
+a8dL4iXaOJ9jLxOFSw+mev5K1vQ0n9lKHg1S1aXt6ilEpK5F/V21YVuHnEA
CLpTZ0w/c4QBBSbYbK+rDWr6G3ggvAab2ieM92bboW/OJDYVuec8aRkjvVZU
CGZKsCI5lxAHd7/8CgKt7lf+rATCLJEzv4tSd1aCLLTTq3xGO2yhnC1X0lin
PDNKLKHPZVhH4E61RT0uA3YvrfT3IousDQCljktCOD9Hm8X3otrXFaf54pvZ
Y4v5F1R7TGzXY9HOxojesIYhLQINXnDsXpD5Vmp0BvYuhe7ctXrpwtwoRnKH
Sdtp2/eghpBAMUVXZ0v0Zhbxyn9l81xBOLnnNg07OyMyh2hk5tLwwQ4i4ms3
R4DFYOwZ9eubqvqI2qeTxTKyS5dIR4XzX+NoB7LZ5FdH8MOs9GQQEPHJdg+l
q8tNM91xxFEd9sDXnXCBtYpfTw3C5TXo9uB4LBp5sWwMDZHJzWtkMEJs+iXg
Udzr/BbS2hMYCGxmjo0uJwxz7qPGL9X2jlFZoJy3H+nadzE4ojiMwNUqG11y
1DJw4sHAty2VF3JSoskVKvJHcDtQc0SMfuIanJpA5WXN4iNeadv3dEEXqinM
/Fum0Gr3MEyd+ZIWhZKpjMKvlmwwJaKDuwZlIf7yCFBEGp9C8dLzOxKMJsOx
gBG4bueoPqEa3ns9lamVCCln8PBna+aF5UDXaqK3R8M5FPBF2g5ucOl6WFZx
MX5RWGV2dXXYkru7wNd9g1FhBxtGKXDZKlTPu20jClUNu9Cudd8a+u6Iig8Z
gux1o/sWn3d6iHAf1qvzZKAYFbyrGY0N4sVuluhbf09/H6VQzMXSOA6ti5tT
JjQNvJAZtGW8EwQMTgIsTqq/iOMMKM87uiMBB2iRhhlxIG/PJDFkAt5YbYd8
kwwqVy7IfP1KSJOhDRwRBogOKFUdCndiYux4OpJOI+JBLrdTLXd1R53wqCrD
y6/FTRIYtLOqGI7m5uGTtwLrlfAQ/gsXTDoQotSKB3gx/WY3jwbrfyqiKsyQ
KvX50WwqOklCi3WOw7lqNkBBn5zqxX2RguetQovSQG+r2cyxwqCo3sm7UY3S
6adNJ1Ia32zdnIV6LHWPI9l1jaw+P6whzOiR4p96dXxnuH0Am9NymWEErLbH
4ww69OjRxb233zaQal6bh/Qhg+P44a7GNqU8kjJdRjyMgBrHleeAvvO2NK7E
l5EVk5WmJE62HoJXLW+G0SzB72XSurEjK9RPBgrt1hqoTKMlEcS4swcXqowq
KCbL0Awl3fMNRyHUVD22E76RMdzFAjY9VGt9gMwrJPKmVaAZtEPw5AgcUofd
HslWkAs/x+KGoiD2RwqVYxMOef1+u+GIt0WlI5aJrDMVUb3CI+8yOxwXLwvn
9vCEbcNGMj7tnGwl3DpluOOAm203UMpDfttMlBlg12UYkL0qViXPwMlZ7V40
v25ziJcsLw08L8TCLpr6p8urwKpioWqR3UeirljInxSzt37ofocNH6Lr8UPJ
RYQQyNMa2jqEmqAnhjgJaKQ0DQcT1RmJBqOULIsuKqd4huqVlizrOh69taab
FV+CyhxA0I9gKKi8gW66Y+vc80ALM82OkfcO38cRFzS29IqSawrGGIbBU4mp
lh2rn2f6wja00hehJvChdSL82nTOLMcmww2yOjmhgi0u2BPGoGsCx2bOGWhZ
WjoJSeiBFZuYoWcO95winWJ47x9kQKjafwZvsTYg4PlT3EVJWe89/iYoVcBw
SqRqGoxQeF7pQGKpZS7NSQN7zjB0AVtEbwjRan4sr20ug+f4+6CrVDyRb8B5
ZhcuZfhgVMu4eduAPAiH+W+nJPStl+KKQ95RTMOb0Gxy4z3Fz9Amwa++eiYy
Z/yiV0RTg1pLSYzRRzveeR7dCITQnnCzlPUbR6hjjXcTza02gzurs1zFZ1t0
d5ioHreS93hYG3sRiytXlJ/Xmf+JPOwTwM5FAxpmHHyCa/b0r8x0KIAvPtfT
4KXPPZVPeMNbvKuWidHl+YrTKvcSVYpTmQBKJ+bulYt2chqVoCaLbqVrjIDz
tf/uhZeYt1AW9qumqLtGF1hM98qiG5zX+PGgGp/32p8UJUXr7c+QW4SXSFDt
O8L/I92RxQpFZI8qwpDOf4ATSoYM5mfrChO2WW44XlhCSMtYXEF0ABMnO266
EBAbBl8hbePsMFaUraiUukvFUWcTOJEy7fnZbVY4wDOmuleUoMW3sNVj4E5o
tDrnsx4zV938udpaH0tK9Nl3W9RbRZXm+4XnnOkAg/Xyj/FUkRP7W4g0JuUN
BkIXUMM4I9H/zy69mM+du4lsr1t63Xqc9xRU4ic3rlntHPFtg2xjuJ6Qs1a5
5JDu83D13g/YT8Yq4w5W2i1ts/DqQHGx2Ki8M7ZHoeHabPUFP7Xt9tv8nyH2
M9Sc/j0R5trB3vO4vhPx8Rp3Ss0PZwxkO19V6E3qOEQ/mGdr/JGuc1I0Bl4H
S6qhA67XMBgISdn58K9fujVUfLmGqJrxewH6s8L09lgyXg+8t/FJXAIJj68o
w0xTwnhJYV/ph9Qz/6F2yT10gWyFEnazx9oWXmmT4toH4ndDAdxwfdsSkF44
Z+mT2cpkHaj20kiGGTjrqw+ThfIfjgRJWS6pZh0RsU1PklZNsDjgrEYPD0Hf
WFWeNwgVgRRgRkAUZVbq5lBPcDjOnolLub+2TRj7qM3Xn9i+McRKs0gRmtSV
9y+3rhNiOsyO8znKFLI9hOJObprinU0V2Cn3OgeEhUC+12RQOa9WsW8T4SzL
/YlVtmPc7aI0I/Ya5exHbQpmvSV0ODb6WnF8eTR0nvRIfO8miDfaBR09b15O
mFmkRvJQy57W8G0ziv5BrwPWgN86fGzqOU12lc/CmdiL84y7vSWsXQc+Q0H8
vKw1Zx+7BQvmQevLeIcbkrA/CYEErv2CjVMja0ebbM3iXN9WomYsl63mgRJ9
kHWXq/5aLey3+03hFZ0et3Ci5fc0picHgqGNqcDRZg56/oGgUu04dYfP9wOV
Q7q1R2PjHKnTfR3beIR3TrNRuX+cuwpgCs5muI0a+ZHTh08ZBlCP3Kmt7Szm
iwZO9UM+0ekDnXM8sILf1+JMz6glCv0hjRkIiergSTJW5TxFiS16JAm2Kbuj
BX1zXnfoITfw4k3RBwNNUITbeid53MIVljgIoPHPtYSoCXM2/hGfCz3ZdDIE
WLTrPwLYSYQDuM1AJ9cF2EDZ6+yT1tkvhnKfJ0qP7qARr6BXna5ZK1PLGgGo
GbabooJIcnS/jI7yCGlmxPYGutsowlOP4emOi6dzJ85Na6MmlpSTrYVCRuRv
vAoyz4Uve0WP44Y9otWNclVS8MkX51lJF9TZvcNylUdUYpsznfbj2/RAnUA4
zQien3FKScNN58koRuy+TuRmIvRAG5PSBp5gYyS84ghtYvo5K5DWTSdf4osY
ikIVbE2svcTX9qEPJTISJuWNFu0+V8EwiCMwzA+CR9hr/DkQ0chIW9gDHW/T
q+DOOHgsMPKvTMZrlZIluPSAD14mDoDNk/uoLktfI55gBBM8ejrK7dNe0Uja
jbBcn3hXHwhgcWXmBBfZWmTh/eH/PrTnl6FTuY+cjBfVRWUeEWjwO3dSPNER
kziUg3d766wA0xxFc9DVNBJy+56E2Hsznhxy6PCMqvK7oLROwuWPh2QAoS7R
WF9IRImz7w2ipJqKLPdlMAn6AocfjdMcusa+UVF3IZOWvsOOcsRyOmI88ODP
3RDdrjgqTK5EEn6JRwVZOHWMHZJo2cAtcbd6DONeUiy80nWTUzORszkVwNMo
peZoxBbmuCxwXxRgeKfafgL7iZlQxZVsXzzVr2Qo3gpXMczZfIkg74irDdsw
lkKUXE1vxQ9IhmumJ03JfM49JXB5ChBrkvgCzj3oFLDAyVB2AuM4tBJhsT4B
GsGMojZPRxTwZdrgiVrJ4tR8HPPDktBUv9i9xPWpKdw3DmA2XXgRpnzxrRty
PEUW106NPxt5XPqjeYggZLcO4B01RDiA7B8WPyyWa2mvQtFioHw12HF91iSn
0ux1RLWunrzH79XhvRanp7M0TQ0JFAzzKsJ5Q65/D5jSO8lfmUo4Cz7mZyge
SE1dlD2ym73XUKBDca0GWYB0dAILa+EWJS7nTTyUrgGeIiaGCAr0GSWcGrDE
NTYv5HsOKG2QvDy6VlO0FPIWqUj8hCnHs09PH8t1AppMTAblmQBcxNFjoVru
8RWqgGEE5lyRwdaHOZHqmRzJgC9AZZKjOPmVNXQbHscDV1PzWO7kqzyIIhu5
DkbjjPsDSglfl1Ob7KFqT4Xama5R/lhjwy82DyLh+/mEOlBLiPxI/vT70f4U
qHYrfPFDoashCEpSoUXOgqy1VC6L62ng6qcpieB2E6tAQxGpiwSxB0UkSfpe
VltJGvJGGBMtK5tuwxH8wakVLreEgppDHQ+kMtCPL2eRK0uc4o0uZPHg6IEF
F/byIru/tS6jaYonmKZN6wYxPaD1oMHGzXGssptvMkFcsTEGZOINKw4Dc0oH
Ypp+as+pu6N4POwP53j4qx3NEou8p4Guo5sTpAReFhsH1oKprJbWHitQIEOI
Jr3eI+KVx1/4KO7t3cJJEBI9oFCtXhfvwdZ8VebI5hcQgpPBOeQlxi1wl/eC
hOP6AoLspQRXv6Ea9lMIV6L7dl4hEM6dwwX00nRbrGZsCHK/DKB/bs0pkzCt
guaMk1CEjWaGx/k5ix/qQkoYUUUKQJBJlKPN0Thm3TmKRfXeaXAN90EqD9FT
Ro1WUlo5z8/Kz75+n32N3VhULlYxTbPFR44ggMAcDji4FzpJ66pxcIif4BG3
MXUexC2fnEEJ7yyk4LsN8LNnarPdf8Cv4WqLAegmDTjTMp4+77+mFn/eCBAG
vEulWmXWDDQdJF7Kft+G0zGM150tWW/jb3bW8/2O9CfvLRLbsAnEnYegL1ho
3ySPuVbEvpnmn9MwqFMjwnENb2Lljfx7KWIwjQrMQaL4KoBHVTs/47AqaD79
TsnlcwL/XSoQWo7MuXUhTIAvKJttF+VWSW5q1QTAwnbCOjZae3JhzO//+Hum
cPXZxNIOJkVUjUkzfb5xdvH78EHLJhb9zXcosy3GMn0eStc+PGaOtybDieIo
L8iji0XcYbK/GkBi0BLqLDxySz+slOj9D7L/MpebWpVDII71A8JbUI9de3WO
NCg77GdcpFbUxef+D8O9NNSHYNcFB6//uD9DfkbY2yTK9aLNCFdLfOE/+Igw
FTxyGohMEhGF0JBIpW5Pz4ARfE8o09m0HYkZegY/Qc854tQfjb8YrzxSAi+r
ziVYQIeo50VcpKuNE5V9308FMRMBCtUJLGeN9AlTe10d65zrzBfU/8N+3Y5d
Me7mBCBmOB9uYPVq0KMKvdztpk+qM+8QZUa9CZEVMXMMWv4PInHgLwi89YPx
sW3YZs9qUU4lTmA8c7y/K/ATF+Jc/HMEPbceZhVn4nx9oE0AOzTf9ZFep1o8
8XaRCvfYh/dx2c67BLwfMNRp0z0H4SDQHqTtzCA5ldStstcVQB02uLa4xsO6
1m7FJh0Ld0w7TkzsiEr5bKU2vTm1OErq7o6tQ99/74OM3rG3xQpu9XluT/we
cGd4CwhvEwdQOVf66eutqWhw2SpJXtFB1qAbFe6MqJF6FOZ/sauLaval3V6i
zY4IEYcStyhgB3arGjsoTw6iftgUmozb4rnXV4H191EQ2Z1q4JTagGO5J15u
NImC2QBp2FuyeyU/rTvH69zUVB9d8XT/VcIGuHt82F8SnasIpxTaetvTQtJI
+BpG2vrUV+bHae0X+Z+uvfWvjh1WYVrPe3KTElVFaGY79Y3CgynMvU2vrFr+
OOCGBjxs7hK0fez+WVltUxOrbQJwLCd0CvqlDYULPtTS36ZREVn/0agsKePj
pEa4mT7FvQoT4z/krYZcDJbjJArRktGvSEFPD9Ufjni2nfmESJ5M+R6sooVE
3IqJFu3j3qdtCoitC8VqNdWIMEJzoNSVL9VlWrqgFdrXss4/b58FjWrcpoYL
Wj0++8a/fDRgGTFXuKmrjTZO6O6CFyAapUTlWbmxrW11fWno766yJKsDXBFo
C03AwzHNmm0ZmY32AfB0wUThEBYFJ5LODF7rcfbWnNyJBt+B+w7jSvVEIWTv
HJE/xK3e8+3O7lPtXmn0eSFhKaqv+zDhPzuuPXJho7jrSESbqrHSeFskX9zE
urx4bObVo1RdMv+U+UW/WCJODQ/goqA+b0rFkvBxd3Qd+DS4HHZ4UpNSRtNm
SSlBwJZD753GX2Torsbiv6M8E1VJ9uTBrXTtmUxcFdhhVmf4aaEu4prDEoHx
H7GU/DcA2lIyXmB1cFPo+n4ZvV1mb318hmkYycMVGK+82CtO82se9VjZ3hlH
+vp3xUBZMMW1Kp8orGWgGkG63qLr7mbCvagi2T76veeLiuxKKXKDftE+RjrY
OKhyZ4dbyAygmRTd2XjXIjb8FmBOxf46kgh4hhQ4YaEU7CVmAmrfAcQ7TMYH
iaGcb5UHpElLaCZGNV2AJYLCaoaX7KzDO6OMCxVf+9autwVTKbLNcf2uhi9y
rh/iBF01b/iRab0Z8WdXquiXP2bSP41HOSV7zJAEXRIvaJGsk1trw3yYtuMo
4iILETQRIOXQVYvg4VT0VRk1z8BLmOwfr0SNW8OT2z2RKP7pesxm/mugsLov
7FhARi2rSKSwgNBrcYMiKsyjLJ3VSdcz/CrV2KLirg+xSNVT3tepwpXoluge
Ic/RmxC5ZL70hayBwt8NvSYrCxgDV2FiC5EKEkN6mbODQNSAfaPnD5dE+2Sf
u6byj31bPcYhxmhJBkprIpHOV4AT5b5ihOM2q9LR8kKD9ojjTtwwzrMfObVi
czjERMkTFtgr7/X/O3jm5XcZFpZ5kyZTV9fomOjN5GRmHs5KQIBYz8r9b+Mj
7SLjxmPGiKQYMSfsE7ROzallSJeBO27VQERGLNcS+y12Ys0jdMXZd4CMKaDI
AGZqoPOq6aRK32+OR6D93+d98LFwi0RHB15jPgt2hDlB68bt5JaEwDsRrPS9
GpiIQU0xari3uDhrxkg1q3fHyI8s4Rc5ULpG9Bfr9Gfw5UNbG1cMGfI7/qpz
X3N+2ID6ScCA2N34k6BWG/yoFRBC/s2YoVVQiDJ3803yrj7RbsojmRmilYfz
j5pCwcklDwNI9L/d1I9SHfDCIwdNIYh0Avmfsf9drST8wGnV9td6Ubt6EnQD
OFSS7kWmtWOVEGT+lysyU93RnpJQbt1WfsR0NloOuUmJxzO4paJUfRUug0ew
v1oh1FHiHTG7l47Ai7Fl/2Hd75gV0a2FlMiFgxciGI2jwhJ7D/5ku1tjWU6s
W7VCBorhg/lOI3GtngqDFt0Ms4vhHkSVSJxGTJZHltDlRYq3s+wXOMcYMfo0
HQJanCH7TFpzzhtcXcssscbmSVaosO2U9st2upP/+rrIs3oRNwrRwoWL3uXT
LU3meSu84+Uk5vMkYL6BfczNLhx8uZgliVFVa1JICoow44C4rCKE184GQy6M
pIn4wKjnVefoSd7bzj7ec6uT9pLzzrvagDWgJeV7Gxs72Pj8Q0Ppxn7k0xsr
/q2nDopwWyo4LwW4Z38aINJ9OpBo3R0aI3n6woKkyOMc0xYL5MQr9WDLIJTA
81VzDVfbMsWKiwZjzvkpm4z2uV7stnUWcuV7BU9YoFiCJ9sZB2OcI01+9ZwJ
5tTDvLygso5h6RrNFBXOaXSXqDt9YDbP5YnNmuk5qLTNLXelEzBbglAgIPkm
fi3tR11AkkAZmfF8g6IcZOIdBhQjaoF7YaSQh4QtA8osm27ngC7l+KLDVMJX
uXgzHI3cH1PChN0u+6SeTzAb078wR8JSSUnx8vdZKQt4MCTVSfLH01hSQFzv
sFcqeeh5fbk+IKKGgb/OQyFqo/JWu+CpuoLBgZyIzSNNHGF01ZJkyrhvCLCr
MScgssQN4V1vT0u+SoQmHyWsmjpouvrlBLrDTUWvG+qPmdNTDnSdrYn+g63L
CqbwXGn59bCD/yv6l5MXYSVpqGFQ/GNWBRyhfuP6GzMDSy4Btp22y91FPUjH
qeVCk3X3FSoJdO7HKH3zzMf6USeW82Y7pQbHAQfX9Mri2kNuQRkGxEG9b2pQ
yTw5ahutjgDnnciRfFC4hiqv2ZDi55fYayifrSA5ZXsYYwQMEB1KJbngvRiU
fWbKIQ8QkgXDphZTyR8m8rwpEPFrUagYlWilJ6nkvbpFhDoJIvPv8fl0frrO
ZECuD1o37EYmCO3TpN9Fv0MFPHNYbkI4xKeF9atXms2epumZZHHP1HUJ+Mqx
Gb5FTosdHX2p40so7RpMb3OgSSs2WNQxkpIeuYDZHh7sEA5G2gqTh6be+7B/
PBZUXBWlXoWl9P3HAqCVFZXoLckCkuM5H42Ok9FOjAz8gTQ8ACMks/8e3ywy
IwvJdplzAijQoaRRv4QfFuKd6YPFSM+TxUR6sd3mZUn9kh4OBywFtqgbwZ5O
BPXmWB2wbRQayOdsgiXSpplp0LJY+78VaHQlowTe7bK1VSBt0ILIc+bCLeHD
4/wLOpny7WziU+W/2MMwoHsLJRTCMMUrgKrLpDnkM1ebjE0fOJs43TIJisOH
i/yNn8BDy5tSW7fgxqPjJ04cW5qcpw7DtPQMDr3uGXFm5JTTPXiRfnIsJg1h
1UTq2X4Wfy1pbVUvTs98c16ezpTjk9H0/vJ4MdZr4qr54v+ANaL+0ElXS+n1
Sq7kH7OnOkE9mZpiyqGrj0OPTdvPHnEhCIrUXvOVet01AW8lqfVfMSpuwflp
qnWCvCZwHO3bXsHVeD73AOUFj8oF0J0VjWhIjRzot4qI9hvAV6tDyZoVpQ5D
cZVjiIAVa7UqIU5HSH2hkc12k+w+PdzqCSB6LKlMniAo6IiGpfj7964aJigC
LrCv5MKrVuAP+87C63yd+Xn48YsXCjBpFg2JjjQCxAAi0bng+O1uN/6qI6w3
be5PBIpg7y5cZuTiThKIrtAUdvMNgUIYz2pJfzLrlp9v74ifJjG8AcqUZxdO
xW7I74Bpu9Ns+5aANaNTt7D4iTQE6n1eyB6aQGXkRmQdhi7KiEgyylNA+0cS
WOhp8foKbNUkrL0dtbJwf5pcjds9LBa6hsKrNSw6nVD4FjOW7owAl4BG44KU
OTD8otSQhQmPfEUCh3Qu4dpvbcMvnE4mlsgcoXYiGda471gawYZsYevVMZKp
ReQSeQ8bQdGjNBxWCEHjy/phMIFGCtMpYpq890qedG+nCMbrbuag1d6Iysh2
fpcelZZehmoa9afR4UKBWBvJl0o+/umKsSibhIcbHnpHWcJbLNAvA8cP8l7d
tjg2FiwVLUbWinJVlbWFKllef9BK4F2brYQDlbk+eQaNem2NtvVnY4HGFalG
snkBdDGLEqJ925Y3ZL8wQRoPomO9hj+L2NYXmBlxGOP+S3bMTgXJJulJTyNt
IWzLTcFYymMnk/mP4EhIPsnxwjAh4yDEfX9o2/bjf8MkPdR4c3NeV/WEhaMf
bBMJkT4F04h1E7qThk6PUFVAkUeQD6VxtRpwjnAIVL3dg3zzA/IKt7ru/xQu
w03aRI9qTCYgu2gpgvn2eW+vCo0f/kgi0sKQ11aQ1Gi89+/XL8jN5SRTAO5R
jSlUtfANATAONbH13elrE5PMcCr+3r2HAuaAF3ed7uuDheDj9BOalCCacZ+A
f7/k5T7aTxMUuetvN+E0sor100PCGOXxq7odzsj0odtcxVNNe2fUuG4aqEwh
sjIbWBirqUYcTnab4lGSOSRqavkxs0m/pY0IBAobbXHCunecASoagK143XNh
wS0EUsQLJDGZ97sD5Y7wWfxuGaUKzghf0UaE2l//rj+tjpbYPkVWISx53sbE
ULV/Lv74VcN1uGpSOBbdKMxq+dm3tU8PGByJEf7PkT+xStZeCQXoNknaaeJN
Pv1yG2D2gIxlwPNldm/gKQ90c/r2cgfi3oT504jLf3G9Gi7blYvk8PWw9mI8
mVErghrqMboSfCervctSGE/ESJ5+0C0lET6cY56DfwnPLkcRFszacSnPdhT8
s6UTHwHZt+LmOjCLjMxoMaBU28LwTdtg8WXqan2RSwhqMQJUu56l0o6xrqNo
Aub4GwqEuCCk9EgWrvwqt3uYeSsglenRPOekcDhaj2Z6aBVS0BmtjYCmZn1S
0O5xuYpBK1nzXqgubt2K92qVXBdomNE9Ymi1f1pchnQqBG8t8h49Ndmcf0qo
8hiRG7VYt15d51nX3QTLc/OEsOSpBl6U4hzaCbjzY1EnG4i4OAGeCU+NzvoR
aNWTRQGVUwmx2g7KeQ/WKs76FPQt8jKxapsv1K8o3/1sPphZ0NMZgYG47YMW
zMj2go5Lpu8W5JLzE3SktYQJt4lvcuPkv4IMjrtE7PD8EoBrgry8Hwcv8wgq
0PLTON/QzxH65aTbZKAJoQehIuqJdWvPZeCe5DdjjRu0xtnNSQrGtW0TOH/O
Eo69BHTi18lKxTWaROEd3lP8wacSiGZps8OTfbqFCR8qKw4D6SbLq+AtVoEX
VbXFMB/aFS4UrGHejlvH9Wl7txqZRndJd+qN43z6i4Thtq3LGYhHD5tZoLx4
8OQtW0RACcaHTvAZkyEE7BAdi2CaWhx+NRg8rD7jJLMvxyFF7r2AfrBalF4s
1SxQXxJ5x+IbNnaS8FurGlWPEr6rWUwfex+VVONCX/bilVaLLZR2wRGJ3kd8
TQ4PXQsPbIF1dzSzpOrMHPUTIsBK2ug9JhfJUekXvju2ilwMzm3N8nt2pr+p
ZhOeEP7+ULEZgAehwfUvS28Z+GlOvx+YlMi1liRd5gMt06ZrsRqY5RD0LKBa
i/WHv6g72YqE9ExPP55fz4mqIxTCJst6IUvAj4gT5qEemNvj3U/LPegQCrsy
eACpqpfGrAPyaKZCxt/wuGLzf8s8Rz0OXZYGQPNRjb6cDha4s2GRFvEHVX9M
tgysv7bGXcF/CyAoxHGC4l9yZMkSuKgGklXr1zL93r/LFlqxJGVy75xlkbjn
uaBvnsj4wfR0uWjm8UYgPy/rqvYIu2LupglDjUs8fiRxKwDn4oaputDFHiir
7aoHxQocXnASTE6JC5Uvt0sxQ8Kl+v9YtGCkumSlCLRlvmDkgcXiG5HruMRX
bguZhEiyVR02xrEyU+4WR7/CPyRlA9ItVHDu9XKWEbXb0n42axHqSKeroDbH
Pq/J+8kbq/8mDfG4zMI/MCCr2FisRUsI2Ynt/GNalCNKUSUq9Pp1FZBiLi03
hvv4LXGrf1bul7jrEvymRjNrOc9qrinGc7pMRAZhpwc6hDzz3v261jOu7RM1
pK07D5vkB+ERFR4rY33iIkG2pqU0oQi5AuNmnRYGttSV4NHB3sf3JDIqB3k/
cb9fLkx6Af8v7DgNo7ZAr1elyh8v4+nJFvJ9INXKFex64gv+WjGlwvKtdE6U
qa3eWztoA3ff3tb4MVVxDR3MxdUk7Xn6S/6x+3SyOP2UO0ScBZi1WP4U3Nfy
Oi+a3Hkx6AVPJvOtLnQrMTSKKEtixKijpPQ7punwM976dsDaXsGFeCiubhwe
esatjTT1sKXC/41fiQIIhu/AkbYUF4XkWe7ULeT2OkUP1bJLDJkLGyj1gP8b
Rv1MCS6xaS3z2pLgrQfOg0OnBsXFHsnRLUmcN/Zjpj0L3XRJ9XEeTndQIlDF
IZ7njwctCBJzLMHXDCpCGBlYKFy0uwlXcQzjwszFWiCF5vs5ct0ykZ9I4Fne
SeAoJGUmYPmbNoDH3odhAt9ElCdCBC+kl1jvkl/DHtjhWzcweDAB66FS0oCS
TCP/7hhifeQ2/8DoWOhEIfyGBjzFJEIbeVvxrM69l3KIYTJ6zKqKUJ1iH5lD
kGpEQXqd2P2c9dTZWGqit63cxk1cxvLfUG0RxQk2EUsxhMyJ8TncoxchyW5y
nd9+AW8j1+dGNXF3mQ8ZL6gFESjtQ99SeSqkaq9bImgbO2/vZPemiZB1J78C
oQkgJWUfNgZMjeI6Pa7cIIkvuPRNSJQhRuNZ2w1K4IPef/6OGO6VQ40aL/jf
BaBeJF9Sa1wKkZ1IMQ4C90vzXEkqjZw49ZquKv/QHR21gHAvn8k3CTZu232x
FJIqrEfk+ODuJOKU9ATCCDonfEzizw9l6BxUJD9fgewzf+8wxMr+yjWnG9ia
bI+yk7zA1Vvwl9JjAdOIy+zqQlC1bA1gR5nQZFfdQQj2pny51eG6ZRfiuuQ7
dOQpjb643VtnMfVOkwspJ9wVm1QyWhBKX2e3fPtC2SzXoW0kX+/FZJETbDxp
WiP6/3ZDJC1OqDs6Kt71iP/SR6welR6M8jAb7qbBT9OTnEJUkudaeC7uLjyJ
Bn/Ji81/dKhIk+J7DZDlYIleuFmqrXhyUS33vVPuTj2eV0FgUxl4nADvbav3
NJ1M9f5dzRSmHwaxN1cnDF33zCzUkkIORJLGfU5hEgf9EvnHnes2ZNP2kA1A
dM65QpHVf7rZSlZdkqZ9qxrmSoAdf3wljZaLwAVCoCSGU9LTSNzRFSy7KacF
ryCxY6+9ZldczSQPZ0N9c9JtQQCYxcKJ5ZZpULYC/WUqJLHzj9A4ihzG/PVX
smXMhm8S3iXohH545je4os1W/CYg1ylXc9lWOylAjbFhZSJpleyIh3Zwa/Ac
LX9IKDVX3nMAFOfIkRVAg1+OT0Cz67+hth8N8dfN1CwAUvg1gVXKVpfFL4dv
FZpAPthM3ts98CxMNxY2sAtO+RojYylci8+zHKxJ1dTEWwsD2//24j5lii7X
J5gyaFI1IbjNPwBJVix8JWAEGxtdm1rPfla2M0BcwHe0CxpIWweUesXLEV7X
b+WOQadV7isQVTqU3kA8NLQVXBqsrehIdOVu78uMOlmBy9zEh3puntI/AWoe
roSP6Z7Jb5uPK1Curqgn30cmhVtpFvzKnfnFu61JE6iHWtCLN1O8cBXrLdMw
LDs/jNXSAkfhebGEJJ+AWyIWbbrRfR03LuXjZf+yzvsKHcD9fZQtruYMEyPw
+fMKJnlRDdy8rO3x61wVX6jYSXxEQozDz5ThgF5Q3rqIHsjmo+c9mbXOTYeC
BVJD7Kn25l8uDdOUfNnSNipiOtqPwzEk4UHUVQY+Kv+gq1tvWYvSfx19RqqD
Nv1D/peGsF7/drFcnH04FIC8acyXhBoDoTo7aHWmHLTjc5rzUVrlC6Zw36Hj
mochmF5ZUSm9nY8W+o4q+HkFHmdxIdf70Bn9fA6uc5EyMcEHVdQjEeUKgTpq
0DmAiNuhx3L6gXkPmIauXfGuBSAX2KzN7lNPqeAxXO4ElhfctFP6yO9cUr15
5NmJNiJTMgICaAgcvdXKTX23afx9ZTn2Zea8/Dc+q4x/MoB34GlXYjv6suiL
olRZ+LeHipGU4/1kX2BfYkTPHfCgQhB5ETPbGPR/H5JMq9M3yMLj4JeBjt1o
BgAK6bK0Z3SpU3YZagohHUU59D0dnpfOqoror+kBHpFeb3Xbm3JNyM2C32pF
015ObpBhqqnPOcyrS8t23Hw9Y7aDqW5Zhx5vY2mc6ruX1wzGoX/8zsATYvr8
O6II+B4AFzJWqs3KQuK6smSdRpCdkFFoI4qcSjlHADRcsD5Wyo7ws94+VLGK
AyFbj6sJHKVWkkn5qTrnKYaNTo4dKfGboUxzsWr7zLqIEK74hX1Nks4KRqNj
8NNQyoibTWJvMaGfU6qbfq5M9Prj2WuS4CldgUYIMpm7eKc+tE2751Ghe95/
nBx/ugObSkanIWTgzugiMcs7QoQdGNzVHnJp5O2YQf8lV56O89rXeqmUGzLU
gypr8q3g1jJM6Yw+TfkSWHn+Cy2EEEouUHdLRffUxBZGUMZPDMs8cMpner9O
rZ+bR5rZKGWOchVIEcD0P+UyimpLPTJRDbQoAFTbz00Ftl+2rCtNcGBXWFkH
6gIDP4Y7+/LbcDTn6muiaGE9nGsRFmmE3oMbbVE2AKk3S852gjqfmS8lICG7
IgTy033CFY9hZDKpoU7LAu8YlnitLUlSKjI5aQHQPWiSoDvFAmUjUbmfb8Ei
nh5p8DIdknpCElCYQmSMUUNXbFPj5RAsFl+GZLtAeDhynFectwDC908s/A1K
lucazNOQKf7av5moibSseKwp+nxi1ebMX9hEge3qW0gT7N9dfuFQcwdYjqiO
P7maRIcqU+a+PMmTMtJ94pKaEdxmjgsReHD27r+RcJ+CPKEI8dtkI3glfH3A
y6nw9cuS6q4fVg1oDCktAsrdRORUBBUzvcY+V8IF5Rr2sIYqdHaN2xHgEFM3
CQtIHFl8dwN0L1MKTtWsOdvOe0RjYyJaUXWlVfk1AiKul7ZFnpjJHNtO0hti
H5MQ6mTMfReSwqcWBUAim0RAT9mcSiHXS5DWd2q2ve9PkNunohwJztNDaKVi
wGt2ionCsuotL1rvKUqgQUa/FtsSAmk9r/dmBnE0CQDngB4LyvOAps2dR/1m
rUIU2Sz5SjSWIpzY9/zBN/1gRnsP0672GkrOT6mQMJYUOA3sEDnk48/TfY7T
UlyOpiKWj69e/yA6SUgzEgV/T5Yg07vgOprw5YNJ6/qn5NI983qnvBlGQX1w
fy4ULdky/ZNdLQKu7q63y/xZAIDBe5PnJ9uZxu/kwZBSo5PWRtI63SnxLFRq
VQqt0iChJKMB67Gg1kArIGfH3VccVEgxdnxDOz9PUSCR4Q9m+1lJLr25sX7o
VCu03Gd7WN8pDIaF4+I9sLAigMFsw775EP/bBjAZ+mme2kOD5Mu5GvOuzI28
RxtUhFwe6O96fEgxq8e0RyIBoDAuhN4vLcGqtNtxL5QcQ470g1CI0mE/JIiV
yScatoCU3UfjGx7uhcRg8VsYP4sEklDhfLweKM2462j2isiYwnTJW+kBaQM2
bi+ubLw1xHsGB8Uk2D9+jjIQPzRzzwrnjK9XUF9B7cUKgBc656FIeJGvREDf
NUyKofQfzTgDk6130H8THJtCT1eOuMfJm2r0sE0wI4oTsRYHsL4x9tueOeeq
dW+BKuB4FEm3eK5VNxZnwG9WzYeAV6P6Ka3IYtW3blL7xo24+p1vf9zOWmR3
wv3EGS+3QhR488m59WGV8n21bot4hK8zaZVhaWzumcPCTEUN9EbfGmGDpRRb
BnJxgOpeqnBWAtQWBgCsVdYNDKorSpaGEN2EC76K1Vz4MJH/9tfY9IJXprfo
fUJGYFI7QlGOH7hESuHZ/IX8FN9bQi6ATjJ35KQ2Dr3ch/aWM8LZJ2fJOwax
cVpqGjaffePEbvip761JKpSKVMarVu19mSMTBRz192Ynew96527fF7ZikFLc
O9cvhE/VBi34tTpxfBPJ1qTWOjShcS+2VSMRwtyxndfcg8KXqv1agG9QZItG
R4b9MzdC6soxQJFBVGGIr8eEzL8EQxE86ybhygK+lMz9Zo2qykmchnY85bIY
qOpf7e3xY1xLcnCHVNjFld6NGsRraOEWAFz5FDl2BlllQOcPc9wT05I2lb/9
tXePyvmrxp3llJXGFsem/CnpuBW5zofDTDtzCR4YdAChnB5aNDdWQ7OfVaar
Bzm6cMCKGA7i64ugs82MuZ6jSqUgiJautP9RhM2yU20A720kFxU9p+07yofR
aET4w5tqpKBdoTTp+AGxFedJlqNzQUziLVztcE0yPGERKgMn+PvTLsNOmEix
HXNnxVXLfSAowitOn4M/g9f0r6gzg0pg9tPpRQjW2slSQbIEIC8svYPBEI3+
kkqZq+DbXUuyRV9s9Yy+LuSRZBvXQhNSY5dMvlIyctGAnGMO8SxNWAJ7LG1u
5UczWtOgbtnZTnd92qQ5EYzWi26VSx1tZoHkWThRCQl/59gsoLB1Km7az+ru
K1Tf2l87ktUEkJG9dSXbCORu8/eeM2YAeyt6+ekdXSAk8LMtViUXnF4lAAge
WOLmQjh3VyLmSpXf6L3YzEwCdjrEngksLBOIfL2cwq5PWBnAZF7XN+FnO8G7
YvQOX+Ke8yzp26RrBFzuNOwBPojc5lnuPO2v1C9FyeQgF3NqK+UNJQ9tqjmA
YwZx+xyqaKjn83rjUWRfTdDnWUWbZgRre581zrvPMfQQIKpz6I6uYJLOO94O
bX9rhchOCs9Du1USPyn44G/P4542tVLVH/RSSC5Sxr0WyK1XHO7yvEV4BiiY
gXHE0kjFOKfmwy1QCprYlqF57eU6wJ3Nai6gldV/asm7+MTRvUcXe7FwKF+a
eE/3F/wcZ70SfU01F8O8x5QmZJAmRcCatZqMus+9DhwsV9mCfAOhaCxItf9I
i+/0bizNzNrL/i16AiFPxt/GmTGVVccrZyS6aD3RtBOoLe866hGEqy/RK6RI
p4f2swjji3WkMEKAGYP1qZj4VQdBAt1nPtR7uAHpnPY2Odh+YwfI1/94BI0e
BWVeR15ZPR3hB7nfydWN/MWbAgIjhkQ+kgfj1BJW1WI//nTk3pKIgWxBDweW
jvGZgY0Ru2pUDNDOzKmI3cZDOjNGiSqVjKpj7tArhVeBU0MgakiNs5LLTfIq
ZesZ1YZzZZXtzt+/l0p9BwzfcbrQ5NWi8Ai/ipiUPrlGmLPX3hjew6R0z7zv
jaEUrsrMQrWD4gwukAA1uon7RVfJRrIqefFKZ4pJhX5g/3SNBvVhQFUt9ID+
7UOHl3Lef7BUIIGN6JAmWdh3CygGowj9ZlEP0FtdeZNtAevR3DgJsxt3xsm7
6oBwpTDhWRMwgQXgZiSm8hmI4wX9ExDg4BN5WymKxpWMHnHip9nIdp+g7IJp
ANSCFvQTbgLYtnBhFcjVAA1AqUGUq5Egef+XgTvjc99mQUtBypKnuUa/EjED
pKNPV/NnIQJNggh9mnsRcIFDkCjIpaygyImaqmgVLRvnbX/4Ri/zMbSLqwos
B6KNcPqolGwTFaAZeuLRREjUPg1goXzxQV28ZZ+u/Zf3KJwt8fHMcFVcnAH5
whBg/5KsfoP/iPl8+C+mn30Z/Sq8CmHPEaXQ/fF/V44CoNcZa0iuLBKiPfyn
LoCdVveoQmxDx7mIpdS+GKUJ1Zza6PsHab+42+FqxezGIOLG3PWGCPE8r0ny
bThv9q4z1dM0/ZZyCa+lJx2inRjyKVklupySvhZOaUDlxMBM7laySuMeRkw5
MLNW3TGloW+IOdz/F/v8/ThChydkd2lASP9cwAQkRvzMIY09bTPngzkgCKfl
2KB2LwM2QrNYoWu0cZFXZBOTHf29eC7Qysi9riQ/NJlAR31otDbRE34f2DKO
6YpoRzrdtzgW5NW+RAw+XaHz/K4fP9bZA/U/Hcros7sgkleHtMUIE4AhW50i
lW7niAoOxWhayW7LTWGIRJSO7l9yEKJ9Rr2c6NpvdhDu2/vPY+fJEUmbW8G0
FtBRQaliHtewj1Dach/FULlnfN8PTCcfZNPWnvn1PGceFP4xgcmgNnneCdcz
40MO8PCkiinRJZpU1BteIEj+o3rL9PRgH2NKZYCkR9LCRkUR8gLEEP5AmIgI
IWf2d26sAWdnkkh1IvyplYiSL6k9uNstmmq9z2GlmV8CILBKgj+Vkv+Qgi9t
lTORnOKxjs6l/PsSVpZmPiQCb3orSyT4khpnDz7gc+4lw8+s85kuSus2UDVB
kS9uhBzEniAVCeiGqGuHmRuLdD/kwD+Eti5OPm2Ge4kmSRd6HeqqlU9FZ7Uu
mYqSL3FfJO5btvO4aWMRx18BdhUnEQzPiTRCghQ3uSju40ESUV+fkvQCClvf
XBlKKDupczAA+n8DrBs25RPfWzoTIYH/TU5MbiitvVppBibrLC5DcVrXsD0K
HxEMsatGu5zt6MPvhTKhk/aykSzFoRNvKSK131gII85hu182/h4npnW64ZnT
FT0ta/6BKBG2MEom5JK7TKxBiPOb0H4h9qIXPbyjhWbdl6lqL3jlUs2B4QoT
FZA0ni+iyxx0bbxi9hYV6hAXBdNI/s/2pKJSUG0eoeQsGE7kdMW6HSJG7pyj
kB2MKLbT9R+02jYqDYJymHxkD9uaRwrNo2NZUZG3Miqsm4YqBKjiNUZBWPZa
W66S44OUsFRI9aFoVWf366Eqt3MGHedTX3PPi+kXqawgeO+l4C6rhNuufsN7
06vU5hRN69/W8tLQ9b+M2ZUJcjzZDHe/4BE/UqDu5PAZRQ7xljirdynR5AIJ
x7krdq7wg3qeoQ4QwvZDzhDDJgSkySfCMf/7tsx5ovEZLOrWhN3a0SHv2o0J
uhZ9Y8szf08I0N4dSWNU1Y0vE8mVjgdrfE2MWH+189j/tyaTeQc5rBoy9Xir
mR6laX2b4Gbs3Ncatb8HvCNzOTy5HosVVU36SBmyyf9Zq5sP6kO3b+maudLX
+4wnra/dviXNIaF3Jirjjg/JKVsCzdMNSK4DghlsdmSj1POQzHSl4NQGrCAb
pjLFGqpFRogCtiYonp4IZh9UhkcldOZ68y696zq69iX2BFmuenuDbKi3GSJd
52oKn30CTWOAVv9RAZ6JreNpaH2xVTf4itHfNC91oBSmoZjxvwF51CJWe5+r
8IGRe5NxWKxfT4IAKws8ltrdxTuX1j1VS+UQGcJz5GWj/oeTOyaG7836+rP6
WEGDHfqCzZbF2QEuEY+01z/kyS1Ti9VQtbVzg+71g6CL9w4AipRoLwtccxWq
Z0s6hFXYea0ubsIH6hmrkoPU0q0YlYGrbzcT9A5McLnkIHtFK2+FivesGali
kDt0qNdmSKBR+4Kefw/IpNKddFfZP6+xAnNTyvE4NNEHVDJTMUL9jLIGw7cm
wuAPeLjwm8OOyTHMifJ/Pd+cgLdHSzXe+WrNMSpVl5ljhFHickFxkwfIkuRC
90+4UXX8FrACQ2V57ipy1zWnDeqkl67RjDT3G2xjlCevs6DT34xS6/DV/vKx
3+UylZRue0COZcNiB/UoWztq+ElODQO/4M9ZHS0s4H2Uwz8qUanlW/SeaeIV
bmfkzBZTwV0pbp1sGQc2i5RCK5wxty2THIOxIz+VEbFmpkZ4ru03a4fUTrt7
mI4aipM3YwOAEElMbOIO7mRBzXmVJbjoeT3upg1SfG5Fi/qjvuf8vl9yTFu/
5Et7dzZvpw4qQfEFwdISxxFJFqF7YJXQfGD9M3FhtnH831g4Yz2tGHFVGndL
SHpLbdmG4zr0SbZ2YobkxnXHRs3yMeA4jpbDh0cKa4rad1St7XAdtMP3hnrn
kYSezEJdYDknj0j/CqukhA1rpKamB8/v/aUsbYeqlnbdmTzMisws+b8xdEPO
mAnVH6TyqsTldq+XZr6T40nYG30nwBP/zpnacvl0mTb3oBS/aWNYmrXM6JME
MBw0MwXBiO+qCXx17UEfgx22hokLihknpGxhcwShBFGm0GiGFgRvaZ8jrswW
JaLwwJxH6DXsv2OnZyHk0sIr214KJjjFrCou9+7o/DlAYT9oRE0Dyx7X1FsG
tk4ShJEv6/CVJcvCMN3ppgqKolqIgIrIlhdRzkmy6i1A3A4Phvz6miBVJDU5
I0SHvig4C2NPwBLSvcvvKOvm5cOrSQKk9L7wPB8mg/pczu3f/Pp8xiXmWpZI
4/zpDt0YB/C4zbDa2iM37fYtYujoQLToZbfrNkRmZ0ML0+6X5TbRWSeZhyPt
umPigvuwT8XnEpuWVQSpbO3jtPfEY12vJA3VcXdlbL1Y1KGnFrh5XvF+YYtZ
F9hAa2TDppn8L+taDFiWZsfqhZoMyRTkQUxsLruMLZQ2TG2AfTkV3Jf2+kMt
W3AOofZ7Zr6KKGfUUtCWcnkgztIeXeSSuL5lILoewzuXPc+jF08cuVGO2YHH
FTat+FUGGCp+IAuW/eZX9/IRaNmzAVuIsLbjJlwiGyNOynF/bHHjVbh4AnCf
TiLizm05pxvmFiO1w8a8So68302VFVJKaPMa3rg/3Mj0m5YVNcNYTSCGuERo
oRB6NixuNb6l2ih7NLFFx8qmd3jZgvsJWW9LIf5mcIp+46okaNjTq0Rkn8bi
C7XxFFOWPHhIrr5OJYNAL/KjdgL41nL3AsgbctsDV658tYa5/J2VPCv9P0JD
5xs0HbB6iS+b/jyaAciKCLWopVGZktKdxCKK/oRC9phtwT5d66xdVT9CU9LE
DBeKgK1AXFbiyNQoJxMfLiEaNEvdZyoRhPqVaUkcWkCrNskf68ZKuYByWBbe
MjWeOjihtZxmspotHz8TM1zVGh17B60SfiU9Ll5JGhGRgV4Ai+urHK22xG0H
NC0kUZV55mJXnsxd+kUUqxPoJYvPXUueJcd8ltwY4dfjQKBm3Uc3Jx4K+lz0
/VS/xBV7JmecU/Eze49reUL/WVqwSO0uQfGyPjoRc/19v1k9hdxFZ+9z6DLH
/0mBc473Bf4E+bmStAVMpD8ILTrmIRGXfqU3yTOHN8uQJ6iOYT5Zymrh7rWO
e287ES6T7oGCtc3R/sNNRLQJFHjBQzFMRYdw++PG6JOJemQzDVBH0tCyZy4B
GFv3v1phPRMsiryIroMyt4NjDNNOKdatCvqyaZZNoYNCcU7W0yvWZ7TwLbGb
tuHtshlwuHeOJ8OVJ/pRHYNvyg7uiOtx27BscooHh9+vMj1zctrUCgaU5r7Y
/IEaNFGJK3JNWfV38IdpbPXqNqVz7B6TuVQofmBBAx9pAmU/9YcsIUuJON6R
4V3vYQ/wLOVJZ232S0ttD0h+gmfo77ZDcCsHO8zWfXfelaQTqvDlZd/kbA84
ws0GJrOF4lkIqUrRmWqDCah0Da1xkvDGKgefFY7o5qDEexwBvpjFnMVxd7nX
1qBr8storbX2ECg0sRnMxdd1LDTn5aywoqh2xyIfrby7QtzLmaQRv/5Wl4vm
qXBG5CfOBKivLKlfjv5AvQwVV8MCWN1n+F12ZptDCiuwj7KOv7IRezWqTVLE
47qq0r6KTYWHm3DZwa5SDFpOBSg3QQSQ8RyvQOY6RVWVUSPquOuzV5WzuzYW
aGprC2EHJt6/KCWxdku+FriBABGQv5Gvln9SWBselZLt4hjKiIRLcG+fr5er
tjjhP5UUsiY6iQW2y5EDKJ6cLeBNWp5inwK22ZBBXzaiBXf76Ft4urDB4Om2
ViUtV//Qe5iVpJF8q6zpUOFdifkFaHve8xexJBBmcWcU7uOcD21Kvc/F/C4W
9kcqwUmZdtwIYEP/jmQXFRcnM7gNwo5ReFeK7BLy4m5O7kPsgeT8hn5zUQq4
D1NMiC4B09xeG29HcnnXTJtvkBoZzp7p47S7hSii9CcZdrGAgCz4fB4wmsxb
0JalwFIYkmhb81xv7drSyveVFGrJKqExRGkpVyQfe6UUYIdcY32VFKb+DR5o
hzBbQnl/lDup8/lD4/9rVPGs/NiSjUrxjY4Vq+I1aKz7qGVTDn5vE3PwteA/
A8fTwu/SuuQGRLaRF3O4p/b0iN1xwLRzylJJVe0ISV/6H2MguCUD4wP1U2Wq
Fo93l00kH4F6HEQiG86RQdiulJoRAaBGisZ49ZpigKqzcXs+hpUQzKa6oGUl
/2XUkgh1k3Lcabbf0GxZIzeT9tXFJtfzsewFwoSaCB6aeDXDWIicbUwfK6Tt
uh4H+eGnzKGMJhmUi8Zz3soVvGynAizgH2HdLDy0tNnf7bkNbi6MJSKJvGkn
raIrK2dpc91SSY4p5iCM/G6e17x/3zh5gbBnLEbAYFjL5mRxS2jhMLnXWIhh
npikwM2JXvdnEfKEi1/uGWCPGtw2ehJbG8ZrNUqesgCTRCfP4PW/FLptPVPm
qmscpeRvSmbqDMvxplyinIy8rzGV3YwiAMr6Pob4TzbhAE54rER6uyeHYib3
MLY1hmHpfM+ybnYFcMnnGZ5qDmMnCypc2caeM7bF9TXUgSl5nYpo1uabIJvn
+ZV0iQeQ40ID3S2WezPbzR24E3v5w48nrMdvJGyaIgeTLGR4Jlgav5Ib5rcL
HXpeI9Z0d39w7eYEni/sfJjrKzbVz7UDvUZzA6RUykpgYWWPX8QYq4LzY+YJ
fSob9JhOuUFqGacGSGqd05j7QNNJp/G0sz018VejB4IoERHxx680W32vpV2Q
H8n1mofMWS3XwSDQnH5vAAdUwwT6gp8bK1tzeHxdPzopPnphzaK4ZV2JciHb
dz4vRxW6qsCIvYv8IVUC5GjODeRNclnw1fOTTy8jAZJZ2B0B0+sPTACcmX3g
T1fsHu+W0IMJiCVQEFJWBrPZCBpngS9mWF+IWsL2+lfn+FV3C24vUGacIub+
nUVh6fTG3lwgoFOfDD0ANBEg7xQqASjbV+QsrcgPPKT1HkSlcEsI5wHg9Q4V
19TL4ke+xBYvudKbTakMVYwkkTaPp7CgRApF+HYFpPtirF7vhLu3JTwpuI9x
UvJUxYp8d7BN8JDPt1zMYTaR8jhin3bT7xdiwQK6AHL6+8n8l7NaXPiAevmB
KYRxYtrjUfi4z3MosvPwB4kgHHhUWVWvGBXrG+Kuo3tR69nEPcXaNUZ1rKCR
gvCrYbzrphdbVpInWY96kxP3VbQaAjXuGK+bugspyNg4LcYtsDklWC3yBa0G
uCyZdCIVlQLNaMkSBjTzVkut9GlkasEcDLnSaVGjPfmzfhDy/Kk4g4nXnK5n
dY5Aoreib+k/3vplcP5tcNebIx6Tt815qJXGI8SRTdmm+ex5h2EwcH9Jkpcg
UoOsi1VkGuZiqfVopW43CGCGmkLKfbvnHOek/Q75g0RzSt5SC00UwzLb6BC9
80+zY2WB1Aj1a+aBy2MiokUgwt/UHuDDF7L3KbvyRkiUVw2NYl1Ncz9bYn4Y
SXG0+zd4/Rc8ieuPwzR3IRIJJcIpv9r3bvVCeVQ8SOZ0gult+l7xVSESxAAK
iJEZGNSwllSqiVbxBRux7XsYIqPLwaMWlsC7AbEVp7Q6utWyytXcVSPZs86T
s7OOBZLmdqVRdoKNRqGfQrYyOQQe4qwbVxY2IbDS6JxyNBrP+AZ80X2ZOUpG
b/V2WUdLdqE7RV7JWfnX06eio8v4icw0Y0pXTbmnDfvITD0aSqz38X8t5Ar1
VOP66drYcRRTuRcmlbeFDbdcwKaK/gYGAoAlCN4iIvuWgd3TVDiOf6sy8hy+
2uks8vMv3t9OToX9/Lm1XedKelCJZy1LtZiSiJcLdvN/ZTMdM18ar3s19vMu
sdqnksLCtQYlSD41GsP6MgVtuGj9VzJiEXESPH+wZ757ecffhWKnwYybkYAs
M64pmCZtMk3BIa889p4RhlUt8V3KhiPahIhsZNbNAHPnP69lsgibTBFVzM7E
zCWlN9cbJ8H75JkqWh3h+dEaSNTqP30L2hYpZ/8cth8RQJPB4oXCKZ59vHG5
QOeW3A0fHUlVyPDsQFuT25JVGcHQxuZ7MLgndH7WCthYG6f1TmD9T0icNGEr
S4uacq/OCfHRu50VAM19u2CmID9IWVjvwf4FhyfIF8t6Ilp3+xSk8mssK8al
QUaHCxFCF++sav/wrtYWYH3GTFPAlvQYhfm0QPtc/cmlZqMOyU+A5TKcpQFC
OZI65Zeow61ognH2wWdImg95ms44muF2dhk+ohbJny2laFs07ycLhHTZWq8p
srrkId/TzHFzKRM1IpgittHUfXtcDYMb6kFGYUGQSwnzmEw+LPArdX6/OMUi
dzdHZ3Wr6a/N2pH7wX8mxS4Aih6BGnM468xI9G7sA2zForpo3DKQ1oUBwa6r
sp96bkzn9fl4+wjvdsGhIM+XjcOk/JREEIJWNtgyfmNiRDCT2HN3fdvR7Mqi
IN1m8uGUj8BzTNNV89wPRSOmtHCDMqCe4A3fMwi7TQZB7CrYKceT++xmPKqg
d0p1bevgQF1sA28pCmCHjGVXe6KnjlPQOfw1TjywfQxtJEAC9Zvem30fRMjk
7QBgLfy9+CEyVnHxU14v1X5Ik3m/EyGBaGJKmziv8YApwLDbqjIQXKdwtL26
ikSHoY60JQ3go4MVsMf/XRWN1Y696sDAWk1PlaqR+m7R5yRLiHVLyxC+fF/+
5m48WcrxQ13uYHt3q+06rnRRWQAaIWAufEMcyKF55ZZtVelnu8A8jKwU19zv
7eeMNtY7n1LGAxIoWBYjKVRdMkRRe6+mSB6uhlKEL2/CN/vLIWRlpd5g6PxB
MIgtLbrPF7fsp5ZfpmTiNPIqiI5Z2xd9nMEytBerE6wBGpM+3ZrvwHnMJnmR
8ytHlD79Ubg1wTmei0yu23KKjQqzf452PqgUsbYBqSKeU2Z09nxj3mBG1Ou/
XgH/EtPanWx1UtpJh3Go2LRmEiiLLMmxlZM2SD459mdVhlxU6y+FPJXzu12G
2otszCKSL+poz+9YX1sPGYErRaP6iZEwIIvKzPwqGesP6Xs/wspqxVo+qMIS
/4lAf4wweTlve4PzOD1FD0w5OQP9y2DA1fJI7jI5Spy2rrbfLqCG1o7ZWcNX
EdSAih9QK0cTMGscGJMllTLD3ir707vB1MHRyNTdHEggxe7T2/94ViTUQl50
Ctdd4lIuiLC+M4mSwIXBwGMfHPkc5o8fIrwzDulwKPwMh5I4PvAiCBUgr+XO
ck36Sw/CmHSm4sTkVYrCZKj9zFrTMJe+pgiWIS7Nx7Guh5hSMyDxS+H9buEZ
dbc70VhUoXAb780sAZCcok3lalJKDma/aB/MWtADpJSxQthACxylNaCvTFvE
sTMpR/YwNCIx78OKWcRxhMFBUTX0EZbm8Izgb1pSjhTON6KctpZAKJETFGwZ
fmLKu95ENhBQ3+6J4QGBDzdcfyZtie4f/B/u+RcwQGHAhVPdFjyi5ao5NyNS
8jv+bg3s2ivCLf1Q4EbNU+fS2f22HbrzH8PkOpmYlEhuh8C5nVIruGvcRPNZ
QipprN/MFBp+OUqG9X8ialyXEzc06M1M0UdFjZabcc5n3y2dGmb6QDrpDsAJ
7WzChw3l5WQne4tAGELZ63gH7mRU11sykp9FgsQfrFl4GSQFbOC0qwLouDzi
tjXOZhIud6dXKoCcRjxWAUwQDjtZpXKryo917sOSok+qSHNVSasip9dli9qp
l+PbuM+1A5fSsI2QAQQ6PSM70sLjVp24p4z0vhNfypNDT5IoE0aG3qtqIKcF
60ccWvu4Y+2ApmO+H3AjGzxhdq2WAtXOlFAzbX+kBMUlk2SYmIrRU2i/0JpE
3k3bbWC85OAURd0Q/OXTDOlyK9IQIeVpJ54/liYDIOFYN4M/xELidA5Uq9cS
t1KvfJ5aZ50tjG1e4+26cRNy2+ci7TqvA1ciTlzjDfo2xGioVCk6EAvY99Ug
umitb5xoJDxny186w3e3NHvq35oPwekt5KeQL8KF9VYIVl1Sk8xciiIK6Ztf
2G9dE2zAoezm4PZh+Vm843WZGzB01VJUmNQNosnu/3Ihay3SQrqWrOY4yiI1
+xISlTEyZUvHo2D4xrcJfy5mEf5KUCuyHNWEF7D0V0RtoBU8/+G1puWijyga
BfppoDEL/n862kN4tSC2F68zz/8ipYvUjdhHl6J+tXydAsfTqwozK2LaL2M1
k9VLQ3q1GApjiFDbakrrEvjm4N1OB+85FNjvjmGlEWiUrZ41igKLQzAngMoJ
DsO6sjUPUaHPcNyd98o1XfYXpupdHrdLoMJQKnHirWwjRlF9OL0ZvSFRc6Ap
cmg/r6V4nBbiOGXzkSiJ05ja1reR1ocLwEXkc8iBsLn0rmQp2Jj7RK8qvTTp
cLk6nXb58IGZW7HeXWCVfy2wyGUUrB6RBO6Rz18/qcOSEDX9MiMIo+i99pK4
Ar9FbOdC1/kigpq28WxGmeDaD/2OQJh9BjPzZMYOE4R6sawuC5mQWlsNqGek
qy619o5yNDRzS7e+As17WokgtWngwOJ8RJxeh5+Fjue8FjRAif5k45hItYew
LW6myqVVjeTDPfLHzADNhJYg8uV5Yy1AFfewvTeq8KNnJ4l9deo+ssJEi6+j
FXzsYsGykfeMIOydeOdVVjL9J15Joa4iurBbOwGJfjp+9XombYyYC0KzvrF6
tdyIq8LSM1e9ls2rp7saEabYZQeXu8D4csOAp24hXUJiPSzDufTjSaz7qG8L
rKzu2+7okALf7pnzhRl4uFwAKvCNpxqUL7+9Pghye96nWugXdL6j9M8YQXrS
mdSAmq/LO1w+PcCqihhRfi+sJdxRSIIx6e98iXSFv2g080jGKPiNDb8M0sdT
NwJFTho3RHpbnt7KJrutXorydUzXHUUEVw9FR4j8r459WeOZBsZwbsyxNDMR
qfAQlkUQeo+DiOyaxenYuBwt4lB26cNQEFQNkbK562HjrxgY07iQP6wNLavp
fyq0vX2LInWhOSD9XKDRifQpPCWf8aLEhWsT4o/ZbMAM72qhtkmQQF9x6pRm
3oT1pMBaqeYPxWH9JRsa9lWiOEXyC7LVXQ3w2fBdW/8TTN/DvwvINYCBdx4j
b96cE9sSkLYjzejiz2Ck7IvJVGPtr6CIuPkxlvtfIRlOV9FUAauC+G6+uf+x
IWXmDZOlf8XUJ5yxQ4h5eLdWVn7jvYmT5dwhoriwD404F5feUwi5GYPOMBoy
wbXMFXPb0+6Udx4HiIm1HWc8Md2hC8y/ZKcsFR2nHKGCaoylceSG5uBilimx
+rKr4l5mM7U77I6lm5CbZ8fTLglSUZtKn0Ht1bViiA91SIKYTn6o3rebFLoq
a5nOkWX80qNNkiCIwfOpbVu1UeiPUbKCvdhDOkmpFYzwSNAKSJQttaENPU64
8N8qL23Lq/f4MWEexpbyQ17UrehW6FlwCc3AwGqomv1Zp6Sl9ILo5sJtFT8n
0TXxwLGj/GhR8Z/uFWqYpRC7phIrMjgNrALHD5o+aGjNg4VKmSMPpUpLwrCO
+glBCICCd6NisDSFG4qU/0XvqG0o6OUl4Qh50N2OBQs32J6Uabi9AIKvhPZ6
dtJy1/fdKv3wu1AxQ/xqCCVVNRCwLqOByk3W5vpFn/5co/2/gxYdBSL3iV0Y
Kh36+U5YH5vHtl8t49mqIm4DSizZancEN0bHGo5H+X3ZOT9smlkbROLCu9JL
r+busYJ5jtVrQKuXDg+sNVuXmz4VeA8QTpATI46Tx6b+vB6OZpGx/LDbGDB0
i68V6ACUYWvhu+F98Acg+tyzEF8842ymZlsXb9r2ZAj2R9uatmKgiFgh/qGm
ADd9PbK8MhrM5c+cHxPgl6KUkW+SgAZcs8BLf9S1B6tNWJnKlo5aIIZ1q+6d
x1CNfni0tufhKRmo+9lRtiuqLd6CMxGWV/J1g45pR4zIkyrqbgYgqRXgQvOD
0qkcGsmCOaeaE4LPIO7AmHIqDyu0H7tP0j56oNug+8fh3fuPocCmKdfOxJrX
fCmcTb4PKxdU2aZgmEWZaR7TabozyKufepYON/ooNH/aLJmU/LCMY01eVSUm
uisOApHkNKKER7iLWqUR0AOmWU2xhpN4YjK0GRKlEm+lXkrKUmm4lZK2HYKD
ybLpRcbHg4TngvvlVkFy+mKTdLPzEOBnGnNTVjrDMa6EvOglW2L7kUS0883V
MNZQrDAb4CmUfdvZJ/w/P6wk4XX1BV1uKBOgOgmawl2wtNCFmAgILhLQ2Wuw
2cHrfAEwFJIUt6pwiyMTnYA55dL8cuNAYOnSdbXnWWWJsHspueWMttLaoPT5
cukMvVJdQxGYtgUmmFazd0MxbhIZa+tvsemRV9TIKRzqwfnzsofMoNJ7JC6K
6/OxqE30j9s4FsIeHruTfVMuBD4Xoe32ZTWiDdF/UA84aJmXj00RGRqlvLF9
0DsSA/O/0V0gVvJBJmWhRoRrGbQ5W+UWc+sZVn3gSBeNti+mVilTC/rbye80
O/qp8b0wR1zHSHXPhgcUk4E4iNbYB2NAu2NkCrEnFmuD2grNn2OiGkzMBssY
GF/bOk+ZEKWmMQcVReW2JhDVvR+Gk7+fWiOK70Cgq89FsNWZZKsrWOhNaE6M
x41HCxWiCPGCUcc7WldUdPBD7xEypiAxiJOGqq1h6dbYzKYbmJTM3Wu2eTTV
7HdUUvR7HcWmfyJp1ztL2E3vpxVOlPl1z+1t+WxVAEs6vjJYTF7KxqnYdqOa
QwIwfge2pgW9Q9dcAO9zeSsKLfZxq44eWDhrWPK20jipDMP2O9WjQfRZ1WRt
Fsq7OjOQuzL149PPw/9dGTWJzs1Pd4ThBIYa78IrG/VrVZjGfpWKmvdvDL6N
+TCMuMsZneaIXt8E1glegOl2C4SZsPW8Wh90Wau2l8XJ8KKMdsjxrfopN3WW
2qLKZgxd3spsflE0giM17TDCFM55lZhS+YOkk78Oy4nfylET1+vf3OpOcPSJ
sE78ATxX2DSMI4Yjyh+ppRPCS4oBpFOe4fE8u78hD2dfsOoYQf3JvOINy9eJ
Gxml9dwGdOK+eg7lZJqNVKnLdJ2ge0B/8FZrvjVxBFc9zrqwAPwoJUKUK1jj
oa0D95TCRFqD4SRCA3JuMIjdyQhsKw7U4kvMa00Q2Q6e+JYIcOHvb6aGThv8
0kERVBeEMvMSzh+IrNwp3ODWvPcOPLcAWnwJkQsNDVvP6/hlJLII9BW36kCw
+XvzPecsK54VldarXrzAZFq6wTTOEG5s8ns0lx7NBW2zZlwvAt9vMViI04yH
UR9kRqZl0S+v22raCBbGR514RewDl3Yl9Uyekk7VUPY9bNw7mxB3gsJvvJJC
EwdvzfS/LxCqGPb8O0uv5rUbgIhj3CAWgkjN6x3gKQjJix5B+nbZ/oBfSka9
aRpxFSNTIU/YhOvFyfbe0OE0wRBmjSQoweffkIkffiFZX+cHBD4DOuB60dcJ
BMAU2za7AF4sXcZPxtVvQ9aQskO8oN25BIaX5vT1t6fMzdvGfDmr/J8tTbF6
j3ZOtjIQIWbijwo9Zon3Y3atiFpIitwdDbfOexrb9DrD/0v1s857gir42Vp0
OXaG9dNg6JidPvrnvTNO/37pZm5kTpDU3Vk/XKRz2OXuuSc6YK6WdLWB8mMT
iAbaLto+1HyOf0puuNIvufuyRdYB1KokCs33PNKSJd/XlMZSpGIRspm4zDc1
2JQP1CHSrT8KWLhW0bxtScA9sw2R3KctAv8lRKE+vNqol9r4RrJbDH6vonkF
NpZ+Mh+PWGNv2H55/eIkjrmg0KN9d5Og+I51G9htD3WSja7tSs2oOWKV20WP
bPPX/PPKLbgUljPAJ5QnO5zs1a/CUqaAKvWcLI0JKoxOTtamogPf7vk/eRtT
JtneEkaUmxR+JVirxAAMyXYvkZ0LSTQsu7zjYwQFpOnbAB/d1LcX2slwjrMx
v3oeasOZX9pmneVHbOJQxX1i3OHlh7zEm6JobudboS3WJI1wJGaaog6Jq5E0
ZqSIuFCGc8o8sIiyJeudVEvuirmB9zGjq3VH89horaTd4T1J5xwqAOJqeu5s
BvP1z3p/rlQfc6coSP0VRkk1Y9ejsEhY/hoJiytN0pTgbZOCnY/+T1lCI6Wb
7kpkorQEVH1VLwJCGQjMfnGvATWw+ekRB4+yhjQa3/ZHYmknyWn2yaIhFdxH
kqmBW/9ueanLoz7CT5N8icmDMMxAhHOXm+wTli1scQlnAKudEgm5snvEiWDW
Q2ACDoBkC1bRfucQYfmKoH5VT9ZL6mwZ+RI4+/GD5SAvHAMVGRWuy9yXMLJ2
5lFPOYki7WeASvBkd2tGGl4phyyTTZ9O7MrZNFCCnGZQtU+RmPqquVC4ILqV
8rZ4wrJHEp6RIMXVzcSI+b/qFnZYvacD7gsYeppVEbrz94orlGgERRL85fbU
Lx2BQgnhNAt27KDX6t9MkoRNgJ0o2jte6dw5mwfYdv1z+mTk0BocVOvq1ZQB
jdZIWSlFzQ6Bi0QFDttSiUUCFRFDHfnr3619iOexZ5VevVd40qSE3Mzfml2F
URcwUEmGa01+fK9J3wM85uoQk6Svplnnb/VWPXe9xzveMyI3ZvWvxhoYaa+T
5dNAJ7wWZzHiLa1eU2uRu4ztR8UfV2cL+uRFMtOwIistxvTElrX7fTbZwJTj
Bn+y99uDllgCAIhj23hdbc0ye5Lt9cHNbYbxzgNA+lOkiXK3EuF8MkD/N0SF
RhatbtsNXVl/x4zwrcjQ2vzplEP+eaYmO1cjeqgkF3F9eTafFLrX4CYgAXxb
pqouiKuJnogTzdpDcvCwk+3DemwAy2C9XMV/0FjJkWJFhGwx3enwyvR6vPvS
Xn01f43x8H4NUw4c0aVWywjFUvUocrtsIYWXblKoxJT4bsgGWtD/Le90Vk+T
4YinSPoAxg5jtdimVEcWjwdropS/kOrmVlLRR48K91zZSjXikYcgPiWcocIB
LMngwIJHCIjiZdNtBgNLsXwOBZ4bgnSARZMvxDkFC5FXqK0Jge3E6s7sibuA
qE1warWOjj4TsDniuQAZciC9oA8yqWrjSW46ThIp+3jBScM+2VlvBXA4igLU
7e6w1xnXBi+rgtwucJo4LluwWmPzt1wYm7yEWq9eBXT5NXXGPKNRRxI8mDun
dpCkdI3dPjPS9/JqR6w9yf4Z9cuII4MzXMRM9sYvkpnKVnBmcFi25MShvm6r
5P4u9PFy9rFgRwUfpzJTD0elnEiYr6RWYHSIxLmPSHiMl4rIc0l69nck0eoU
0j2/cJi7Z6i+pZ5vw2+LGjQ5ii13v3pwaPhLFI8P2L0za3979UoCtknPaxl5
CbzPt+pJqRKbmnk2JQkpKNlC9/TehylUNtfcezNjxbSNvd5ffPEilNdHAeW2
erQSS+tgHJflLEdFgNz/rN9+GY8y1VxEh3qBU+oUeqbSY3jhK6wOXLKwVLeA
3271jj4u9hL5gFfIXZtwAYTava4CtQ1wVuYUB9XyY3t7ydCHW4ftLvDE/Tlj
Z3+iDvgMyBtY4ZeR1wdxlxvG1/fttSTOdpbLMibtMthlqHH4bozyHcrLkq7S
HUX/I3XVX8VM8U5sRTY9hNPTFDWtrWCUh0iW5WJ4GbwJjbfoWjxLUUEe+AsC
mibW5naUIys+odVuQi5MT7wUVrQZVQZrvuoINXW11NGa7XaImq0Vtk6qAViG
Ln7xJTuXRDlcV2ltgnqUz2zAz3q5RlAqiYRbxjkTsqLWvZcsgzH6bWlw4qDk
TOW7hVaEh2RXxD6Z9vr4GpgL8gUIbBEF/y8hDZVKUkhyg02FblGz29QsXxce
tdaqWRyvS85ZoDcbsLUvALy/T3eukztlFg8akqHGTpYXwUb71Z9M8UhLMBLS
J46T4ZO8X3YGOV6uwQQM7r+xyBuaU6GnmdCvKQgxQ4h7MyyNvzwGM0YwJxfq
YLqGDgCZAX4siB6OqfyueudOJz2wv2KqYUIMXsIAcFYUhq9xJ8eoFrmU7Tuz
sFP16BEDOXepodmJvOBfpWi1EBTYRFNhuuNDll8Jnj1WfblZDfIn1Gl/kC35
nx3F1XnjcQzl58pSqJhI42zpW5DUkivzyiOFzl+anIPq6B0Aw+UwKJbe6wfj
vYjMfo667dlpa+CdpzvROHuhoBsD4/GRylkqevnmS90cGeDBGnxztrRLK3et
0oBepL9MgzoOk+vriunmhmALTOITIVCIodcndWn3bNW7H28KBDi/hNeZQBjE
mQ2gdlnat06g7fckkWP/qgi5WiBNqU/8ZqdcVwAmect3M2zacEKuNTiNlWwg
AtDqjelv1Vk0/tEidH2nUSRbhUIDh4g5uchB6pjWjjoUFiY7Dye+JgSDVJ2x
VKsbMX/BF1xrPRqwE9aiOuXyokigc4SnY8msv7Z3j+kaaQJVcWgsADUzTel5
gd3QYG1Rn5LIdjqiBEyQGIaSq8MXhkEZStraTyFmynkX8WPOUT2R/yFGwwV4
FpkyscDiu/yItqF12Vbngu0Ndzrxlm7EqW+hdTt2ITwtRAYTfwMBH4b+kbQF
RLzoNF7LMnS9VynmhquiFfOOAo20pL961JCM82jFJMW6bzFSL4FxJyii3QNf
Z2x9YhC3x64TazPMV3sx2Btqz1TnVjsFhv0OSLodC7rxYTGR7JLR7OA00tLf
ZMdFxTQkPHE/tU2vCOPG7CNw456kduUW0vkENyOF1pZ3w72MyY+SuaI6iwph
wVqIbwfGjS/zMLvmnJgmBK/RDaSzZ11+KI8Snaas/cuN2AemYBhZkI8G6d5D
RCEKdWxeGDdxJCCuLPQ8gaW7SIIZkNNgWCJQRggw8DzyUIRPMbfddewMkLbQ
d4TDPYFyekM2lu7jvzvQYMaxlAMo80ODCGm4oOYFqvhifIEAHYa+ATDMhMLo
RT5Q+wKid45/g2xvf48zXNot39fwBILmy2/he9MDJG/sDmcIYtDknm8qJ/Yu
PbgAAdxxc+M4tgVqzrTFeduh+hXl79XQf6SSjXyfB0r0BwlwCFNP2A6FJuqs
IsE2Rw/hX1HPL5QGHcR+9baDrrLA2qpr6cxENgqpDt/U9KDI+TG5dEiqGBC7
l0GYt4QqluASRf8RvXwyzCjufhqNycr7yTbqeJYOLgurqQhD8CDX+OuJ96Mj
KoXvYNRjMvSge4pNOyq8hjWjlLJ8fxoGzVHzYK8jxfVhkL5c2k3bBoAx7jpd
4zxQP27SUFqUqE2YYYd5wbb40rGS97IgKv/jhetslKSOcuI27G6VihLLAB+u
HCVu+4K3Hep5O9pObrb687ZTzVF5N/ys/YjEMtL/3T1RtEQKY/sWFiGxyxw/
E4Hij+9oCj+F2K0suggPGuZcvm4dlb316wCyNMwjkjK0j79rkJUj97/mKVDJ
XWQwEiSlDxWwfKPBK/Nf9zMFCY1of0a0QIm3UoGRURQzvcmT9kbugkDV72ni
3DLi+mg/SLyFtY93FGucJ0RnJklp/WQAEHFtZbhic1JEgdaFhWT5hkzfbZAr
cLoeA7NjGCHfKWpe16a/00NTQYmdHe6WBp6ZH4BmK2/2c5eZ1Cpe9kV0zEJ9
HhPv8M0RuWlO+aFOHKZZZ+E0nhSypwadM6iswo71xL/WVu+Jw1qU5btPDUdt
TAGaeffD6x18bLH6hMQzmA0XuEMvJyu79bpFUj4C9+M8W57KlA4Zz35fig/L
1eCaqLcEDPnj3cjOZ0EM6qVqtC1aOJPJ+PVRNsg5BJKpgSeE7V8jV7OKfZSc
EyxFTLcRPirS1tHkRQaWuufDk0rULs/jMQ9MPij5vxZj1c3lVxWy2m1dVApC
q84+bhGhGV0t1kdbC/XTT/sWQxnhCyFh2i7yLW8YheU4ETXfs0d/rea0b1O9
5mh8HO1y1uj1Cfeb+w7nB7MZNrwJrLowT8KuKeY9EQSWdpuuxSVQsOIl6udF
UIZ38Rhvezn6R06UHmgk8ecFxhD58yaFhicbbqUFzZUfowfBrLD+e4jfwa5u
uC9RlgQw/+h4QAnMcOx5gyJ0opMG4kOE6+eHfA1LScVUXXqOczrUNPuEKo4O
SrZeYbUb0YA+rmaAnFYQedzwAF/eA6gQsHkXHO7P0edB5Rlw7/D0wCKZb6aX
PsK3SBe0bWnLNEZtTeyLcnurqhTp6CwCjN18bUeNCedefJcpCaVORZKFsZ39
vowXfDm0ua12Lc1KHOVSytJgVbavWk+MhwLtIajTs6J1Vpeaef7rU+yRQ0wR
fJO1vpq/gffUngoEr5p5dX6ZSDk7H//7MnN09EGRbCpKgtgtzxkhg0PX+Oi5
0J3X+rfpUwubjbkdkP/Ay10V7QWQJG7sh3PTaO2SSeDaudsz8EITEU0x/Lsl
XRg4Csu0c5w3vUDMTfv5FXJD3CKnFo1xfrfUHmiDMLD1DZ2GM2ZD4PB2xpGF
oxrARflBGXILpCevuWI303RX7XW8mOJv2OpAmyFjWdrjiis9Jd+5RyotbY7R
mJfqvNo9mTfr3ztLx4iaUfs1VT/RIt9HFGQu4CmB979GhhG0n9wf7DjNf5U5
61Ra8DcvvUA14j1CVx6PalY4roKUsUQV24d/k1txICGY8uSnVDILqRlkdOKN
xU5nV5YLVVwkZ8yF/sWs9t5Gbs6xdoRpNfXQNRP3xBhFl54uahr0MfKedDWo
27NQ+TOiAZHKYtdq0UVOZRMdiS1oncxvsT2m/3onvPkoam1G2CEwV7L4qcj+
efXG0nfOJIleS5vv3LouiHCQdETc1Qe/HBvAhMc/rNAmadeFwg1rFyCyq0Lf
KxCZsSUflRyIevqyLWsO5T+7Dgq32fR+EOcVa3fVf/G6iQS7i5llYsrZ5b7h
vZIhfYt4QuZYvWBVAhTQ+HSjs0egNcDcdfr4/M8CPfvChEpzRB7hNLDdNe0m
DnArZc8qEEnLzSMBL1eZQStT2iJYCuY9bKi1O5hLd4LoTX3YhOTC+tffQYEL
ZkoDDhi7FEwBpnMqsUe4PeKEHhGAZB2T8y0FxddtnIX7obl6hf+QjWrKymzl
YvzRQdNTWxsm/Y2D8FcFpimiv6W9pKxiY6jj5kQ5B1/4KFmVDZMIBfjLwLXk
FJ6zpiQhS+qJnWWODLC54G0GJvFvdzYf8+EMKPz7UJIgSk/TMqf1MgUZAD/N
jFVie/4SMzBGba5fB/fgaA9VXmMeGCoc31a3O8zh3h1nWhX0i+KREF9qPlNw
LBobqVox0R+DGOzv9c1VkrG0M5aKMt3+Z0L2dwUfL+4udS+a7VjcQVxfOjlP
J+5BcEsZAdBa7fcHGI+RKBCcLto1Mk8rnAxIMlafCg1pW3D/MJ7eHCeD+OqZ
988tu/4BPnmmx+xjnZbwbF7FqRPeb7sn8RZqDPJEkSosgorMp1hWpXjzIZEl
o6DzHzYSure+WJEvv3kstwewNxBxwnPb/kvALHlyf7mz+RZUVO8T/+Os5Y00
X2jTxXjaUhnsZs3ra/lozLCjCvIUi17padQLWJ3ilOBV1m3CD9CNTCKzwDhu
itDUL/xp1ZqTZ8U8k3U51llMXHsUWWwjkk8H2xAr0bj+39D2VytITZYzYJwD
ujUs6vmu5ky5KRb+PXDNR8ZE1zgWVi/ACmpCppya/fVe/8qyGAXb44KcfJNX
IwAy5Gvxkqgpc+rNw61wQ50Lo9nv5+DKCJIzAHJP62huzVUgMKs/AO8SW1gh
SSrKB/Mqy7w8Hwl3dNCwVdW+LmRB/xAJrXAFS4YvmH3jho1yh8LukJrFYJy5
1Cad1ci2CRupLzlwkoLbMtiuCMAB9yWvElv7qlzXnyxVAKWXyz+nZBt5YWkk
T2tmVEjKQN3sYRcj76NIiAcLhnmIYojOVaH/G3FES7weuXO90/EeibIeKX58
osp4qSg54zMubBHouNxC3VptRHfe3hbFJ+A6sOqJhen9iLr8eY76klSkmzXN
xbGVOEspSNeH7uvSZ7e0VuuMWxoFh0GlMUmydAxzb8V37fhS8n3WD4Y8thlH
W0E/DdrJc+Wb1UZN7W7Qi98+qlHh47vCisTjp63SCoRNnyHk6e/wttVttrpX
QpjDj62rYmCdLyS2WK0c1cQlRNPxQoZrmZ/lcdbuxYDHZL2sPCvfNBF8Avo2
mt4xZ2z5qulIXlwNCNRSGDgRP3D+jOf54kQ195lnqfOiZ+fYVswdulB/Jhw9
fx7EQ1gePw7nwyDoBvMVdzRF3ELrOK/++Wu/tQ7VqxJ9koe35dVeDOL8c9t6
GyQB5mJRUczWxOa5zNOvw+Ecmz0nZwL+daNkrKcD6tGuWakWqDSPij2/pAXP
bXdQHIMFVb7L2yvzR1VItZMrZMhJmw/5Y4aBxVXB2IL4qLmkvPToR71dCX6l
sawM/y0H9t08cJKmLulVk035Y/QDx1NYRglb8XNn1YQb/KwtVb016nICnjS2
/5ENW6nVAbv/PzjexODU3YGLGcPf/OAzYbDfCEkx23DFnahBd2pJHssn24TO
vhcX811+CVK1T77T3sBy3bQQK0dPbzg5iQxwbpWkC4b9s0N046pyCuhBjFkU
DhvyuBaysCM7e9jheiZGZn2QTEnytwKxEmiNgJmynf97OWO7MTzpRmYdAisB
/lHkL9vPaItUcptfmscD3k2UAiDiTBiRuHPnfH4KdaH2Bxrjg79OE0wdiX8r
q0Db2R5gkDWmm6yI1QxreW/nIF2zk4dSBReubJwOaBix8kKm1gxd/TaRvsB6
wJ18klWESgO2YrnhqYYuBvxhoNHYh16VhdEgMPLPI3s5TIoZfPOoO/A903vV
3+YZ5WR49eTk8lVIUEkV5oVU1xenOYI2Vmdy//jTvSyU/dd4eCOgXZKA6k9e
GQNIfPo33pptVPiTmLHvq9zqi+qdfpz1NZgeTmNpczB73qD6J0OZ6z3aopQQ
3jyQawL3HdGlj8RksiV/CwX9LUggUpcPgKt4KqGSjptd8lhUPpp12vKgvLXe
X3OQizyshO5/m9TW0KPvhR4tinC8msC/aDSmN89dWWi+sqQ2UfbtrMOD4Qyq
8pA6BKkgsbnTm1UwudRKRZAaLkgkzZZX2bV6w4ir+CsvtlnUZNPvo9/+bwzC
zKagF/WhETxqkKu8o0H7BbslXdqpmEaSbNUl5SoY3TUkA/VB9zamND3Bd6k3
/2CJlf0HPT9J7WaD9Nylhgvrxh+hCJX9T32Ct7t81mBkiBv6dc9G9Ek9tZOU
YLTCu9XVwR8ACotWiDry4clPsNbbQM6Rd+g7uzgVgynw4Ew9GAIYb70PeZK2
m6jQ77q2HwENuPCJhk9RESve4xBh8MqzNwj2PLavNQukggEplfP7PFXhrraV
eWwDFUDYNqCiBvqRxpkt4RFe5cI09vvEV6YXqOCr5sHEGQrqvQVXiEPiroxU
ikRFrKIuvLWqhChlhTl76eqZjayci55kFrfASo/hE8PN7KN/hhp776UGrl0y
+fwWnM0j+Cz2IlcuyI0g6rw+IKsCF2PdUhRhIM9K14lPt4U5HiY0V94ZFUVK
u7MYFVi3ZO481MDfEfvR1Ax/67vNLNpIbmWsCUXrOj3CUPNhOgSKOI/aLzgN
cGmzOpvstaIbrH7Q64rgXrM9RTim8jeWEg0Btfs0aa3g2feLIZJhU7ZEq/sw
EPHJDkgPGV+Uy5WcVbfPevVXsA1GLbAgToQ3DEEkQFbifIYUAFHs29z4msDt
+NEOljvohauPiQ0HHDufFQ/jnSYcXxxQhbLRADP8vx7DVwzv7gF9dif/qPut
4QXeJELXu4AcM8+cWKwEIExVcG4bL2f1H7FlZ4Ab/YcAIANnJkIjLsceUKTf
K5NmWwJqWWQtKvo1rpme4goy/bCDhVn/lhS7oYh/C2scfIDVz/OIad/JjWu5
ps5881rTHG/QAc111FKvnUmNNQ93DQh7A5hP3nmKQlvTO4DrQifEhdlypOVZ
/9K7xdfeo2CWgD4H+ANhWYXaPOOgwqthrUWk+yiy7rZ55Ch/Rpwk7e3Ozq/D
j1UMDxonMwv86/QNVrvWFoqOZxipkusnDQNxsPSo7N7lEO2U1qoUdsYznGbU
xPILigozWnmTDeBzz0vwflA740ISp9IYKqba0ih3QeX9RZ1m/DLo0azlJuPA
qT8efIMF0fansoBjgJpyfGYwdNP1rsyG57OPq+Gt6vdNMVUfUvpSA3elbkgN
/e5R/JHC3nEhKNmoOHGh4sC9x33GdjwMCMNqTKaUo9gycwKyWzS9zj/X4tvC
WXAKw4mG9S2ZB4gvO1sKcwU90a4QHFo2We8Z0+Qdf2o9TN7u802FZ12hgrZ9
nor5X1NtMNi/fUS1nDNM1npLtfJR5FDQuQg5KtmOcmcoeXc9CU3PerRh4LUB
xnvU1eUNNKFSt9KpaCnUCkRwQ3S0PQc4dcH9Gqi43X7GUpEPg1EEG0M9xW/F
SZnmVwx6eo9Ektf01pnG3p/+Wi7Y8Ol+29RPwmt6XWihQ5+0n7rq+LbePorM
84b2m4RGankYaYCdFP1NCciTKNrkJEI8GJv+MIN0o11h3BLAYjpkG21i3Uf6
MtWFelV5Zz2ZpjbBlXRS9Oi5fu3p4RGkRivw9eMlRcJPdTGEGIfmmwGpfb00
VUPTQRZ8BwWwNSM/3GrBEb8zYWZuqg45UxRMc4uNCPGeFoqRdd41DV4lLuhz
KMsN0n9pdvTvlNxa0EUtUxiRCC/vR/T+kQIhej+TRu4r9zHG4mDAQREy8Vzl
FIHgnO2LQxWxvrG8HKgc+RxPftb/CzZDxV6V/+S8KrIRuf4tp5JTSAgQhMQP
GndOnK1ybmxdyF8XMpJaYnKsvx8uGg6RtctKpA5UUXsoHwBHuMmcWEyIlXhC
LU02Z0gA4LygjtVPGCmyM4liXI7TwWrzTYYvwcM+cwEeXJ6wp63h3WKV1crN
mDl1zDJfMyQ7N4BLX8WvHgBoCAzbLArx4XlPFxxaRR4CadAxAvtKtEf/f4S2
ucWGk+XMu99IV8XK9hMma/AXalbd9jC2fFL/x7yKK3TprbHadulP2evL5v9u
rVzVdPCRWdK3eQDwMXklURTcZf8S/XiXxJora3PD+j+fr/4jCOE4FUtkBu/3
EEBbr7M1RtG1HMdBH09siOHA8XaAf2gcMbhLs83AMF/hdrLnMtUr8kd9Ljf8
+ujj2KUw5TujqVvO6Hf7MA7jk4/RrDdxEg3eV5N9oW5DCLdr46sa+8A+dvbq
a6Ue+I7qCmtdD0a/TKDJqKKGE5aynrC6k5d7N+u4cXf2f6Io8VvoZB1rDP8A
T5q2AuTjNI4FjTAeJUpk0N6Ol6T/ks5STDYMTFGUgbht1KIBy4syUkD4YQaV
g21e/GD16zfHEYYkdMDzRqLTLTUv4YZ97G4jYDrhJe6D5dGnqVlJSxxyQFol
tZ6XVIDnBFKbBRj6NqeOzTe8FseXKvpXhDqfwImvkHAcAHNlIbIBnxinSiuW
IehQa8TLxH270jm4jdmmlgOhUqpzxWVwSPRn8UVgJOVBvqX6ofPcCo2cdkLy
Chov4BunznfiG/DP1mI1BEJ7UmGkmbMOD+LxT5H9w/bV98FHLbHtdyXfc1c7
ZuH5eq8K8JZWEox+bI2GT4OKoIU9A9PlfDROMD5uInlH1JU1gg3tkE+5ZeZ6
E8yK4+3txBmlDWkeUCjxBcWg3vne9QZOyAqaxTSgI3t6BxP/4jK06S3eSK60
98juBm0WR7MpSizi4LoDT7HDcVmzIh5kG6Se3J6em4e3nKJWpyv5i+Nf2p1B
xgas4A+aJCXbQW2kO1Xufo/hG3LuJ0fdSTt7wfS08+hZ4BnsIb0u396kpSDt
IEo+p5K2RmzSlw/33gGYoFuT5ZEDu9PpAWr2XHZSLyZWuZL1IgowZFdBM3cg
SIA7cSbxvFZcJeOiNBvR1me+WigrhdCbEchFTnz8jQ8Eyl3pXpG+hcbLLD4U
SMv4NODYoGypFKZKa/A4mbuVbqTqCZbc93YNDtOHy/m0dq2y4NULVkGNKVRq
yScNO+g/B/g843HdbFIgRJHJpZ1Gm4ic5EufrSAaRoBghFN4+BszUdRLyFNH
qjk7rmDRstw2bQ5YiVQTy6RR/HDxX7HiOHfNZr/CvZgKGFUlIGhDQ22akxsx
onM9sC7i71pZuUVdpEAte9jfgh6t8thVCLODmUbUO8S9N2KfdaMYsQLxprf/
UDb1SoFtO/AMd10b93FINdiwrmuHmMDwI+PDeu//tS69637GjArIoR5a429h
CNG5rCyOIpHiiOfMWIe0sLV1k+Wtls3Z8tjr2OF2vNBY11uqcFoUw/1GqCSo
gXKDoqzivgJVTXDcxrNG/fEhR9hPTsfdY1ICGevuIoUp3m8z6YjsG789t6pi
D/+MY6voXdu4MKrnEfPaqe2paekoVyIk/PRdC/2eu1oThLYy2BZ0bQMNGm5V
UpyDL2qphmE8CAM/PaZWnMgcxzhb/fXZaibES94XgsmRWtnRHp02sMNQuHjh
ESU0xndSaJaqkF8hiDe1vxfTJwVgfn8HpABWfIBFZcj3ECCH+oLXjjuSlKEi
xk03b/mcMPs7nmYuvpVXw1iYTQEBfwmu1xCLll86E9PoAkgQwp/FWQlKbEg5
vGhFmFL6EYUQfqy1VP85oppVLhSvreUBSSwcECQYQ/tDX5PHsu6UcUipXe0x
6UcMVWn7sGBjfSObW/hNwKtfykILuPbTtT50Iyz8w/hUzv1/v4CZ4TqEXZVA
Otnbb64s86RRBDk6EuCFU45+jWd7v7ek/7ki6a0nEzUTj0N9tk4NySPR42dq
xUJgnr4Hdo0kHC9F9lKN4fkKEVPTw4ZKr2ILOKSGDQbxxaw3WV2Uso5ViB8h
6uscSxXlEX6v2Hh9KS98XwNdOMuKHHtaSR2IuRaAQ6DM17gNvrXJJcsGJx1Y
aDFRiBmZtXndr6ZmJIXjk4UmoEdD+CUs5A3Tr43QOAk0sROyn0rLVwXNK86W
r2v3PSMuxVoEjU3uxGJ8SVuyzP/Kz70TGB3sWlzdRjR0eUFj6sSOql+htYs8
UlVar4j4waiGtn9IfhpPW68XEjXLhq5eGciJiaxs/02PW0FiwYG6oEEYR3B4
LNsXq0ZPSh9yta0+wftZDQP8cT+1N9OqTl5k/ZaH+TQQsC72pDlUoD/3bwn5
MugbERa0L4w9LYsKJ6v/AYyU5PhCU4RkRcFgPosaN+upHSJ60YIOZq80UHFP
0pFb0tzgXWmu3XX2ZeV/EWNuY94H68rHVBMmI2I6RaqLMMwylWRxDDZcDVN/
3GzYhEkaWsskCMjVL9YqZxZHO/Gu7K8Onu564PQPc/fmdqyIo/quuJsgU+ry
DAJXZoJwpXoq7IwcuEY4oWadbLAKYWoBAKGXg7EC7sP+GNcIXAC+ukgmXRQy
W28vI1FEtn8/oYwaWhRNlBBCNm3isyIFC7kCpcC9N2bp3sNZz02RTB4hNW39
8weSNtVxWdKLhJekD6c8z7US8F1fqJ/yMwAz5UZL52/03wXRDtE2I7AygRKS
uSOkG8hSmG74M2F6sZJ9wr5peWjr878emp3aHEuF9bDOQKo4oV3XjbMMvdc6
upqGhPScRH6eE7whPLItVO+PSX50wpeH6aqihmPYzs6Onl821Jx+AWyG3aw7
BxTAe7lBEMAqwfonMb2bXShdjKPoIOmwIcR3EPZzGt8SAeAU1kuLhax0Oij5
6gNdnyiQhveccuzTiGYkJK8CDeJLah15y6ynD2j1VMrAPZH5ZzzMJfKJzbJi
Uy9+DyaYY6lMDUCBOMswlwBFbqEJTsEgRUnBZ+IfdwY6EvRWypzu8Ql8YSfv
52w5PiyMD+Mnp6pKYTZkbTB/2fOPPhi2xPMUm9upiGJe2OAftmYd3EgNDnVI
rxn4IE1N6FM28ea3f5SCmFwL1OTHCbe1cHgvxc+5K7eCTIJbaIAo1My3t8k4
PAUEOpYcjb7cqZOcup7A0QzOLrOCYpUCm5xl6In7ShdX0ikBXAoTR69GOEmv
j5GsmnQfxBOh3n258YyUdTQfxPt+AuSCjlAOuyuHRKPN2CXcFl69VHBVNpMB
s6UI4IXnJ5HJvLiQUXL3MSbJcKl+g7BnPjhbpS5EzILowwGBUDNK8qiVGPv6
MVyZwmazjp/Y4oJvtiTDstUgLDPU3w48qBpPN+hrkKPfgompeQRHtUpfHPPJ
sPD+DzceARApjzvDUahnD0SlbkyBkBMYR2CQ2bzfuw7lB7LRDT6yw5LfR9rk
aUU89BV01ITmHgMi6q50UYTicuf2SKqmqhq2do6JYogFc5aGCJ7DmWu5Fzsr
xT9sHjR6QNpTqQa1SBq5HWt5KkdJRG2fKxMNgoqRPBqsWqA+k21qJIcg6BZJ
0bbGxwTHqH4p5v9id8M+Qoc5Eg1gvARfO7oPIO355cfl/FrUS/KqXU+TwvJ0
tWO36cqRgR7GA/zyh1vXFkJnJI+kPLQKrklxwRbJQiR1FrKr/Y00fqRtHzRJ
L33iEb/xSYG1EuNfUYQmIK3ngYdo8CEdf8jWZM+4+0aVtvre3xv4p1K+lqIm
iW/5WBls+59YR2402WCu79V0/Bh3BeYHKDnkCnvSJhII1I8nLBihnWCetQmT
O8WPr1dQ8MzrEVjdyAIjBUefjNM03CnMeeVhEuiPxqr4bc2NduS4aKLAA+jv
TB3OuPHZNpI6VtePpiX+gqrTG6tCf4scMgNWNLhIG5+Q2MB5SXt8kFCXmWmQ
M1tIQE7Uo/E9tsinn+f9nnJbz0YAZztWO+hDDouXdCHbVxitiGsMFEbe+p5F
AVrbXM/9NpYcoX8qEotQTAmm2dbHVU5gmXuiiFqBEE5GrdJrIN5Y8fhF653g
8mN9LTsBzKXfwZPezlGWmV/PUHu29bPK2o4IarO3ZXcAKHkAYusWTkqpxHE2
vaSvb2uTdQfjX4V5bQadsKhl080uq6F1Qv/pRqHZvLlAiUcC9eJ8suN8cNqX
t7uCjxnoKYtAlTd2nEYvA7XEMsm2dNkP19wDGWhj38I3t2bnDm5bEthckza1
i67G/mc5e23A9Io9L2YIVWSM49hA5OY5Jw2vsU165LnUfYUN6fAMwrcmwGeO
dUn9ADBqM+R/QxCmU+exsaw8hXbTWIQL+XP3ZinVbeScl7d1GXVQ9NnjD+fw
NCcEzvcBxA5R/kd3Xu7l9Kic/g1h3eoBpO/lZZR+R64rO9Yy5RpsPaWfFArg
31kbqanT+HTTGF+0jbz7TX0UwnoWkJrEfl5UbtuLlkhivMv8ACoFiJvm8mHw
1cUCigdO3Wk2RTyQ1LOhZMuVzMucqWL7YUUp+EsDiOr1cEmOu8dM+tzijoAD
SxUmkiYN8vUChuh5Z9nySTJVsShjBE/EXuR1sY6GjYdnV/TRgydhmU2nw0nI
+JwTwhnj7Ks0F8drQMW3VEuZQelbVGbFIbDcULwl85Q3qVJ8QO5RhR5zAj+G
cHcgRKkpNhDOERRlsu3dVXyGF0mZ+EfdokQHDjzieIlCp3DJyVH5bffjK9po
NSfZdk1TIqaYlYZScwnwlP1DdTuxMEHRtk9/obU7b5W+BCQQEvXv9DVG1ERJ
qhKlbbrdM0+ICl9rpQafhEfEAZNMYPQIAzHUFVMBTRS2eX4AcV7dnieGwh5d
zurDIJgWjOdq3S5uQd7+rEFXjwAR0FLeJ5sK8IVbs3MMsZSl41h9CwfN9lzU
ZpRV1rM1q7bbaUJDkLHFnH3umLpL28Nb+3j+uqQyuEt1+qgtfJx1DB9l3KzC
gv9TMJ1dIxxjTyBbRjOhqq6D3dztBWzVK11ZhAxaXJDMmYO92LekvBOPgMqF
Nc9oeKCRE5TLXH9jhT4rjojnErK8on33nGdWjFAu3rmsQ+dAHUegttSP+HpR
F4Sb0Q4rgHGv+v5EUsNH1BoiFYGU5GSd+r5m7Dep+nZJJXPDvcPuPIx0zYln
u7SYFSEGWVtt9XZeTts1lsonLuFS3iliwG5lkU97UDlLzmjL3xF2uIFg7jE2
UECdOCopYZeBorRUfozBQ+UCWUpkPBE+tnRL6Vt432CKUnvVoeQObRou8nBj
M8G1RyG6fK3H+hzhWNHP1ZTel30erRBo/ySKTY9MjgCRVbuticZ5V4m8wNtI
HRPe8lBGKG1I1MXaGrir1dkgYKpTjgEWMhb2KxbWBDCMqHNfGJ0x+CnS8oUU
zFGofLJALbfPCW8Kj2qGYYlIMgfY5mKEiH24qQvyY1CEvVaESAgCHBdFcYlY
Xj9mlK/8qTUiB7/klRB8EkSeCF2UsCExUNFcHx0fIT8B4hQpcHVjrte04CLy
oboU2+N113Py+5GjRJPpW3ncqTsHdeS7CxiGbN1uvrbQM9Me6S/1atsH2kyk
2ujLc5+DZdv9wxUyxmjT5cEWK0WTI5C1t3rwa/HnVsc5GHUbKLBWWzN2HATU
g/ktqAlEIs5gwY2BceoX5mzdwDwVPKPsc9t/TaU3Kzsh3JujpaHWgmZo1+7x
Gnuqx7Alwj8lL/xTF982YxtqyLKbjXcXoGxsR0rh6IIvgawXjaTcFmwgVPE/
UFVHOxPuY8oz+GR/K7KM6/3fd5Fypag5UQljIZT0CtKLrKOoVVsetVm004gw
irMyY20X8BFGfQSEcBi9U+A7bammbNr9sf79K2fhBZrQqTnbLgHzESj4vRQs
KeQXEtirXVERMjjLwb+EFjZmBGOyepz2SusoVMKnnfqtYljSVotj2Uc1M568
B3zW0qkNPa8z1u3vn7pGA2M3nz0MamuQCFH5P5R6MOMXoZzCir+2kQ51TduW
mN4bvRxag9rr8X71QKgnU8lS/zwsdj4dl58ApA/pv0pC7YJPzXlZbMdXUol+
oxsG34RW1VQxSX2mYVChu3GV/OqdR9pbEZwUV1AXdKYPukDPMOBR6FSqf4TB
rDlzVus5y7SnPYnIt7npUwHLXSJ9+KyK0JfqH5CPnsAiA3FKr5ViPgPLF3l3
zDtESTERkLecf/AxXUHaU4NT3ry12KP1OSmXlopdZvmX3WPkxRCpZ5GJDiBh
L5g3Ii6mnK930m1f1qqpNQW0zXOFvuy8cQuGCH3z8IPxKLS1IXReiIVNhkg7
DiTJTF2l1Axj9vOlrHTquC0IWPpPJcR3ZY8BNpojN0Y90r89tkDNtqHqHm48
eQDRAARcBVbJ5Saxb28EG6amSKoiId4z4HVrFoo4bE0+wSK+Qdu1mWs4tzSL
1ztZs77zrK7iOlfCBQ4A86wwlMo6Yp9gTiWKkJ56j1l3GHxk4gST4F5l8lsD
BUFcUMWIn5xKGU2Wu3T8Hl7TB/8GcJO10LWqhA7Oa5/NWu4UIDx9Q5t39951
eAy++8YNQ84CXHcf/5zTPeqp+OgLUUKTg/sGc8nKzD11MX5DDUy6LDI+3Dsx
evItAx1eD9c9ekLc8ux5Q7yj3kmvb7kjyPvG3u326qlkYuZVkewB2fFlb6H2
nz2qfJ9EdagWM9wUM19oiit8VynSzxE6hNh3VifoV6/Bn0yDyqFHVN2Y9uDM
SHwS+vBnmel8g8RfSpyZbx6Ag8RuIlQYOi1g2fzdkkbtsVupD8VFaDLkNF9L
5GVemqTWjjP3ZaSJP1W0PVOdeCzvDE+DMJayXB3+5a2mzFy+eWXilpdovJey
F+Iuqq+2/uAzWQzuNOIcPGU+lceMC+gtgMIbMs3oD39JShihRIbrB9k2SZBS
s2/3WRMi2yqY4AU3T7A2D4PNm2L8VHlq1k2CAXLdh4czmeJJQIex21vek1MY
mLC0y6sRahm37vd87lFoI/czzO9i/+A7PkMrBIjavq4pENv/St8vp53NBqcf
udoWvZ9kFJ11EO7cpP7uqXfIDCAMwiMKyywmMOpQHAXLV6A0ttePZKJs3lUU
K5QAyqVYkHpBzSDBq5wxWokgcKuT5XVfbhvdUrOQxNBVPZiwQTMM33UUYDSq
rv+7EmrlfpY9+R1UnC7RBHRWj6+iRpjBZQqEDQnC5E/W6U8o0YM7eXamnO4b
cBjNKXrYjhWP81c+gBJbufCCIvXZJonZsCy4grK+CWPvNXWtDnuwgq2qNxHM
F7EcyeUpc8F9O3ZK2HB+apL4EJ4955YP6eEwUD+tvWy6dQ9a63jHHy2ZLOxT
OkJdTrhDXGYfdpI3i2itbJW/ASU8b09T1FzAFuITjRjjiqAAOshJ2Rt1hwMx
EtKVJUmLjdony+2I9v2izj8xZOnS7EU5ilxUSvfKQkFjUUThU0s3t/MFL8t8
AeGjsdHWui+Bo089Y8iEGm3ZmiE+t33M0DYTX3a6Am43Mp3uKqQVAgVUiNFf
Pfv0s5X3VqLJtGdWoAL9UuAjkXL7/bF33QDU9SoviSEAhVoyjqgc5HQD/WsJ
yU7QYCsCjruwgpemqV5W4HPxO0bw3GJd9IwOw55tCmpT8R0/WtADhYiAyxLK
AM5Pe4rxxFaHqWPMtfgQeVq5HLZPVt9jz2eQ9rdRPeKAsGHaS2SIO9tTCiZg
xp2gZAwT+PZ7JwPGGcpaRndgon0oGlMIBIzmQSdO4RhQsQGtt7WKufwAh9aa
lDfU0nA9dNPVhYcDGRbVOanEG9APuWNQMIrgq2GXXI6yOk4P9CKsIsamat+Z
xru4cl4nzJ+co/Mu045/lS01XqYO3FO1hn8P2+gk7QCQ/lFWjaOEeS+3egsv
CWUkWeFQX6dF+aZoUsq5FiQmrxXD2NypPArJGZlBv9jS7kX+O1usYqqy7xxg
ka/nYhYPnLmbw3ov96RJBbNTS1qIpBuQOBazwo8Toi2zDgEoi5EtmTstB0Zo
ehIBGv5tPSEBRdqePuFex7fzGv9eFXZyHbi8cSn2nDQxzs4QLkrfRZOyhvnQ
C2JMqZiHJYXuDo9FVqM/VdIjqNIFdLnsL1gHDUEDSLAeTSYg0GgiYeEjvxO1
6k5YzbhTJpGfOcH4EYGrNOvgNcIdOjDBpiIFlkupg8PsTwQ9UiEO/2rI0vKf
rT9xzTDDV/90/3ZrwjKB5jL4QWkewD//highZlFszEM0KaQweXXmsrFKsS1o
r5yFH6cZJ7E+RjQ7B9hHwCyyMNf3bbWtCHrPuDr2Yj32g0Mw9s2WPtkRN9RO
g2xRd0CIRGysNqgm5KkXHVS75h4yHys9EyA7G7oyrF0EB++gnw3QtjhcTuCr
giA14yaEI3f1AljusFzBunri+FmjDbgb0PY647GsgbWtvvj9Y9dBp/GF6X2i
3MlO9xBvLK9B0ibURsSA1rfB68OJDDr+3F9plKGzJSSYZlDSSe7kULQKnMq1
VSBaiTnjxIDALALuqhLE1eVQhqH+gWX8mrolulYwgxlEgiiA15s3cW9u44h6
UAzvLS0pcpHNVYQmpoNMefIl+7Qr564Vhp3ZUXKv/jMxH/fgza1T+hjw8udm
ThkARAWZTeDonR50Iwczehek5OgjCQx8bJjdJr5CoJQWHTfz+2Q1ei4XKqCv
sivoCxgyFTK8RPxHewWoUWXz8QGXLQ6HZ77+yknBAMrI4RyQ23ndYmseYn2L
5W37GjLDAVctaBDu6vJk3wFB/RX+uxtXo9OHr9Mc/vYWF3MM9POo9pmOQo/G
+AZ5SyRpdv+SGvFqpjC3z6k7HsY0lfsDRlfIuJuieEcHqk4aHu9lLYsQG1wA
d9knQeOYiWqUD/mbDf1V4uCw6BL5cO89yM+2JaaX5Wbzu/RD/bFLvawqO4jT
eTRqn5Ldp5zRqj2XBBBA9eMRDuiOUErhJw1SEsKiu3TlTBffBHnR99oCBo+b
WHzAIGgwvf3O6da99FvNf+GckptIpo/PWy42yH2ucNWS+amrLXzfnoo0/Wyi
1mb3FaKF3YSM5kh/+zvpyN7l7v7bu7AZSd1DUW7ulZexoaX+AtMEF/gPxtlb
fEReF/INL6quj9GuuepUb8U1SbjtDSqbzmRAeiARi1LL5NcpRkxl1QSNNbru
gGllqYPt08pjmQsbY30WE+dgMn5HD/zV2VuRNtbqP3Q1+UZf65XiT9Jh1El4
UtL1wM+vECTaSf64jtp4xqgovH4o4SLf+SGY1W0+idATgy0KxBL8v2jsGzFT
Qwrz3iE2rf47sTqG7WT/jruzXVEyHzOa8zEUgxroI1q2SGL8J0AvVG2x4cCs
7rw7Yku/ucRqgHmUDan0v1Xd5F80VrQ8LXlAJfFEhU381AnVfKq0Qs+ciMh4
PjjmSIJIKsnYEYgQ12GmdZ3oCRT7cc5x8kk/j061X1v06AgnV8MJm/qCXBZS
IANvUw+lzamEC3miOp3IBqEYx0PwFOvvCcxD3WtEKAT2VfGWhayJPDbuk1cN
8AXBQ2MIzMuWFajpFsCmGsBN2iHr9pNAhpGj3XeGGSgBhBXBKq0G1pweczLq
+F18INKP+1r6uRGXzvXC+mZWYaInzQxtj/BiwW57ISl8VtTjztpjnc34+Fuj
iPpV239nzizndJrc3Afy/j+XQgeWR0myZLUpIGWKNbPGTLcrEZHfXr9V3DBH
WQIWfVaCzDd7Gy+qUDeYpTB4bbioVo9IZQMB2SS9x1Otvo+z3H/EI0PZSj6+
aEXagjcXz+VyFBp7K5znonvBk7UFur7E69z3N/erzeLH7V+4P1B/4S5H1dy4
XUNH/FyTg7RHuEnY3lqmVKbdfdWq5ecK0t7CiSit507Vc42LOoIQbNg6i82w
dW0QzjbUWYx8oKOK0DyRZcT6292CTOEGWCMLKAXZQ2VuLGLH/6Ncsp3cw2bW
/BqhsGpsxslFbf8/1VQpueq+8fPargPYURk2Ilsslj5kZ94UrhSNtssSFBAD
KLY9DFDKsyiRjbWTSOfURifz/7EupiDe8JPm2fETvBkoc2hP7JntkbmYs4ou
6Hmhpksev6vug5uV29JJ/4FvYglnWPobAuGCWdQ4MQQj8Fok+xcV6+SQ/QUj
s/tBRO4rvQhCyWEplwgi8iBILFLIJy9T97hCSoa96kj7T6a2/6N+5v66Y08S
rzK9I1RJqPrhkLK0aqyWUlcAY0hWfxR98mkvz8FHOv+55uNF5MTiMqgferfr
sfV+/bFc/qg4Ciq1lQfe68s6gt8GqOSWMohDChLI9HWUQI0d7zHySc8iGeuC
gvla87Zfrvun/ljAS0v98K8KLlBlvvUYcTxC7YA9xa0jco/CaJHU9Na31tMy
e+qIru9794h3V8SuPhOKHEeweP9Jm6AjtDbwy45NU4bNUE7kt7ADbARgoMjx
wQIi9nTt4OyVz6GZZ1/TdsmXELstuFL1eiKEUBYslW89mbz75yiAIuxAiD0M
opdWsitvv9zWHGhc48xiG1VTVguiJO4wZKiH+9HcxPUF+0kTdu1dRhlorppa
h8fg9u1bQ6jADa7UCElBCKGVrkWOrrPCPRn9BvU8ZUdTPalqxbh94etFzfnR
xWh0NOj5uk87sv551zD/mtLIughl0/vBXG6ivNOgYc/qIT1HKv9kqw/CpH2J
mCuMriX+SdJfYT2nNmHF1FHjXzSwsSM5UQNMyu/ik2nFfnPFrQnOUJqd0qLb
nh+uIOrucjXOf7SO4ECv15zaFjB+MelrQ2Qj2ItwFKj7sv8BBkT6arh1w+Cp
C/KaqST5u8a5+G87JDzXdMS7P4wlVgN/RylYvVI4Xfbqa13VMkpL1lUA5SS2
PzyjF23JiELYIuNuKjXbnKHbhp1R27Szzn74iT957uVAI3XUNwUM2MGNmPeO
86FIZ3OJ6bfwgj/nsDyAWOEKapHErzDC5UmiM4lMl/P8cYA4Gjx5BQK+cP7X
sBqu6lq1AceX6hAnZOLKhUxjIC+i3ax2pMu+bLpfs3gp6wsk30VSdU8JSl7h
yxRHAhwX/XWQ4f3d1Vg0SEGCRvjI9D3svnw1OcnJwZL5XYvk1DhPMVesIprb
0jWbtkc+fDJC6Hy++mt8811qWgHqJsFy9gsIBhWY6ZLRTiyYA7l8bdbQXnwq
I2DqUmYAH5sYk+nbo5mAxyeH/c7KE4GM361JUIAdMmO671u2B5B4yNDF+48x
8RKbKTR/mT/cRSo4kQZdXJ0AhuXuM/LNGwLp+yQHsZIWUugtAiR4NIl923aj
MUBA0wcntsxkTAyE5KxarM/sZoSkc2kEg9JP7tRTFb+z6jCTi832VuS+cGzj
DdaI5bUzFaEIMqoFnku+e8ZRx99MdgH/dCzqXts7l64qcAPxpkhQdFwwDd5F
N84Z6SAbNLYSupU69INMScQWNGESuL2asQC420uzMC9MthMbcq/sl6xhFy6n
/UQTgRHwRatLGtXRSYYEQFijFP6Vdb2B+YcEK4MTOThEfffWobSdYFpqaQXF
HWv4Yz9/ak2/I/25ZM6dIStycurLvQSJ34r3MEVCr3TJCbag5iK8V+9Mqyjg
/6QViHX1GOzeSFwrbAc3LNN+1vjWiNSgPxkIOi5Zd/MKdzJ6ypgCX/6an/O6
w47s+4sYNRxQPcmzf/+CemVc4E64WCoL0j+7I0Kmyy9VZAD8Tv/LUGq6oLZk
L16kDlPewRDiXjHvsyl8SKLYL/G/0W/cVxzBmuIxcFSrxHy8Xw7vl75hFgrL
E2m/5N1IhRpJoCVE69pRBlwSC/3RJvjKUzmvNU21JT+KmBRu/ghHMXC59WJe
P4iP6YXEdlb7MoRAJzJ4pAub6DO7CKhzTNOeNdQUn66twTBa+uB7Zw3u557I
xxClMQA90j/dVKcbKurJSnAHsCrkrlbwEUG2jzpD5YuXB7THxNDvZexD5ZJ2
0zLf5uOSifz4JJ60iw+/whPhoxIijGxeVd3ZdXQKGzfeP2H+kjgNMy+prSR3
OEaKgBLmZrgDR/EnsUO/y0/uBongRGPTfo26B62aCTKDseG8EJS1OWh6v5uU
9hB+nzXo9elg9KURpFoIDUwwI9adfPez21ARS0m3wnb2watcEbFC2jcF0g0c
y9HwYknyCGGfmreFH+xjup5AVZU2fdWAD+PX25SWnZ1960HLaI9zzg3QLPvo
bJSeQ/T437b4rJUAttYKL8qHikVYYXrhaf8S41H45hXcFUssb4KjflqmINcE
kKLyNmgqH6AClB8q15pDTHe03TtHlErMndiZlD8cBIlRYYsK8rDK8rx4bD9D
kBw3yhkZIS0HoU3pGmI1X4nCoZAMMS9zdHWRAK8tXcM0/bSDavQBsqKrsAb7
j6xOLbaWik2nPMjmWwjNy7jNtTedZwfsQnBqsMvwfxvdt6BMwPLg7cOC7qws
daTaXV0XDmwR8VdJbPlJQAP0AI7kikE5FW/31aStzx8/CDO6ZepaTnGJG6J7
7aN3o7L9MgWfheCE6OQccKHXi0jpEUwjIuxku4jEFLOcOGolaBi1TfypdlHx
vRS9K+IK4PJevTiGsQlutPKZ+Z7Dk+LLf8+yKExo0gEX7M09JPBNSEU77hSv
QvSVBMO4vQoGAlzEYyUSVDFB1pTFvzIovGs3XZhjgXcUJSx6cpkJpIvvhao9
a8XniAl5jwmjfCQUUfRFvjsno5UHoVWnFKHH+h9zln7ozl/tqIbii962fPcR
UJKMckEEBJgoCr2j1tiwxPZkhXQPrI9mfrdHXjQkY4goq6d+YBfnV0GBUHgQ
fGCygA5NL8THuXuIezVvTMul9uAvUg+umxBZOrNwFAvvZ6Dgg9OFrLCV95iP
zQ0potVh4Hk7dlGbvbgYnkcOaLi4jDDvZpW4Ui5cBltNamV6UllYbVUQnSNi
8TNIbcVKC2kMbG31WaZEEzbRisKhtvFHAyorhM01PJQkt8vwJVp7TAIaitEJ
sbevK40FFgyeO/+8ZrbSW9J5WNa48A/iYCY+gf1if5SQ29qJ97B39Qclyepq
XGMKhVhvDhb6g4Xx7Mf3uxW2J916OE7EvLsgCsxBrjwIVoBW6g8yE9QSeYJN
0nNCHut5VRI/PfITuHFcsRMMZfrZ/mPLBZiIOgx3EPqqyF3gOwJP9gYl9QO2
2Oui6zQ63KJngDDHc1y5vVqFfWQWSaJU6PG3NlS5atmCPm9Vg3bCrzT653/g
iHmP5056x9Piso2SAgdVqQvP6OLb5nnLDUQ5Ss87xzY+2VCjxo6Q0bQPvlkD
cZuRHqbPV0+Ymed4HpIAJcpMtLr3uW0ekVx4R/WrPDiIa6rPGLrjYNS8Vtol
2ZGH4dULK2Ir8Hq7y/+fZ/MzD2rvtSIvFnksPqu0ffBRjVe+szcqS0fjOMoY
+JUFhvITGEqojzz+HNTkOBSJ0fEubhswNCQn7+seDo+zcgFY+yZTpbRLAOOi
MYway4uCcfGWm3uLFyZx4SfeBW2V87oIBQwhmDMk1dHeaGaVO253dszcGqKS
LsmY+lFg7lw5eZCKo5AVlBAukDN1Zzl+gGDde2+gUMFViM3EyW9gcyTrSrSN
YjCDyeShYg43xvog1eXYFVTYi9eoUj+eXAAnFNdIlNGigSSsRnLi6WGdepWT
92hl+KfNPELBWu4IxHdnGMjU3Yue0HLw14xDjZsH+mIUl0Vgz+2rFAQb2NSm
1PRVhLh9cT+PttJR3w9y6brFxjeFIWQ3Z1O1NUJTZmPiTgr35/oU1f7nnxLr
80miTzj3Ptx//NheUXDekwaLkuZ0fflpbkdC/6r2RoqQ2waTmlZcCBLDgcFp
wXSJgOVdbh3FfbiJwLeTgnyMk5y8/uSBrhijLpO7SnvE8D2EFXjqBEFWZRID
h4TEOYfBA2XmMkCJI+zVOKT1sqY2JD34Vt47V4rnERYt3CqV20LHs58n76B/
kXfveZpttzjDFc0fqUmlJwzurg5LkG2oiJYW/R1ok1EN5eL6vTDyZST8lzQ5
NmfUed7hBfFpd1EEbtEKOGgyGreP853F+jq+J4Ypzbtzuao5Adva4BBuq3/+
48y9kzcMpm21NYHoRH8nf04G25M+OShLzDlDW0wDOSMpf8ZpyBiNkt7mKXjj
horCyd5ZEPwT3uBLjQS9f/KepuTUDDsTMiGaF8I5OfrTqXgV5UQQ1aVwU/f+
8a8TC7nEp3kRi28cDp6UADKKnpEunxwfvH2qZJTqGVGde6Po/QlFkSATdiRT
TQrmRFvMYbfGBNglAUhLJyK3KDYvuE9JL+UfVMBM0Nl+cjCGN0L8D+jXW+vG
KKq42exQvf/MCDP+W2dUSQkaQKjU0uvhxh/cQD+PxMvYowm0XDiEqRFOrafO
IskIUdorLtuVz++wHX1zDdaNeFzfqziO4cHAQK34I0zmWcpzaK/LmRx2mOSV
ZpD1X6DQOYZ0R/7KWteQiXwPneSKB+Ogpyz0OSqDm6daObtDp4fCyx9MzK9Q
P4gDxzSzn7mxA3IPCfrHg7E6Urk12zxpFmjeGqwe5EwC1HsCQQ106vtob1xn
tqTt0M6lldGoZHlL8pFOaEdHYOxzD+KygVItsLFNPi85LrH2v68a93XGQcp9
D25OQO3n8/xkHEq+XuyWS8VhMRmPo6mMzr94M0XoGjnY6l5kcUjk7OXjbbob
NGgRQpHc28r7scqH2UlXB50ezane/es09sfDbU/PZmJxOzs6AYjgl6EEEGGc
ZVjNOqfa5qcFmYtIEW8TT2hiyVHoiA4fr8HljiTZOCZld1cRWyKHLxKHqd+J
KGTO5tSzoPbDafEA8JvBRNwb+JKEOBNYcBzfFsq2An09v7g64oF3GotEcsqk
ATRb6kHD4EmldCY/7Np88eIwdPt6f8GVNT0Um3sx6yOwztEj6f/C4vd2kKYA
mocXp8a//a7QTEtJWCwZZatP8SkBPjdLcdivtHin7UAAVIAiOghBsZ21aOtO
Rxzg9zkCuoyfD+R/QDzprwai7HRhsffL7JeIRmLQps6oGhw02rVSxAorxmfp
y8x8sGlTdlk+vXHODmfWN6bPzNhswh/xAp9B7BLR/lDPgmzpeOdShnV5msxi
f/6pFEDkD/25UohoX57a8jLjEwD2QU+56AQ9R/WDISCWqrbRG5KvJX5a8QtE
95hRVvHENr7U3Jw/IrPpWEQJbVYRJZU9IUBvRi1VU+IYnXpiSb0f40u0W7ZI
t+2PPooPR//oFRAMSZhmvOx6LkVYJryoj1VbTjxqO6lwYMx2435GTeFTgvI8
s9qx8K+q7l1Sjbq8FTRWLd0lbUB1q7AxvMuZAZB5USe17ef9n4BE07Z5bLFA
G7xZhNvfhpxkVVCtyeFC7rRDbAeXUPs/dl4ZyI4okNoB/Jga30DeS48BxtvK
+9I3i7AGv3H1wipvE2N35Gq8Kroqh7ina6YKdWzumTfIL4ux9cFo1rVvlza0
7jWVnU3Knkiqlg6CmO5ujAn9KlYbNnza7KTPJqqn+8UxAv/T0BXXtSn6uDFJ
MwYqU94JIZZd2FDz4q+BRmOIz4xQYFTjmtpv8xb3GSjafO7ezUH2QMEvKzpI
BqEz4lb49t0iFOFj3hj5SJaTT7f1mMBx1LsefkHItluutuDYyOMvvzT2Pnek
cu0PZfhpflLrQbkMpAebyXlsILe8g2BxmGurQ1ISlRLCeyzsa2pNH8ZbwaWy
c/PcwcuI9D0jtDJCcKDqQDG9PJzMErKntkgCGmuUDn/3fkTElwR9vYECpFN4
I0qOlYyINWZrVLDrq/puwxXvDgcln4l0MBumXsPFJi8dO9bycb/rsZ8JBXcC
Jym03vfTjuL/Njl9olax8W88r/EtLpen7GDuk3DwKgPClb6V+RexnQHafhnq
+aGUnbUf9ddL3Pby1+T4emM5K3u+Q0XMv9PHk5bbngsIUdbGnJv8qx/rht5m
IAiLrFbVT0SBJeKtKFnfUMhJtCuFmRyGKh4A8R5pOxwSTermMvCYYECDvQBT
zXOCx2SIdYFkd1UAVUUYg8vGWpeGHui6KGZfY4D4seEpisZPL75265WTD8cq
r0bTEBY8EzRhHdul5KJw+u18Rm/Ppk31qLpc6Tls7+4SSZcEgRYeblqPhC3U
GMeoqMo8xzx6MRPdmpvenrjR2dLRBXAb0oAFX18pu7GlK5EgFLI40CQG/k+P
EL5p5h8fK3LFOserpXFIokwbcVOzxctPLdLFB4NBaeRUJ4X10OA9zXEhQK7A
1+1Vu/SDtWk+Sy88Ao2TiY2CjAa/l8A5AP6ZYNCod0fVNe28uXaicWSZ4TsI
F+qrXH+t5uPp6CvSfA96GLx1LONPZ36pLVUKpgD05gIQurACuoihqn1JU5fj
rmKggZre3aoFtELsDg5pL1Z5p9ufIxqIpTYQYD5/3w/DCxnGZzQaxVWvcGjS
9PeAqHjf1WNMjiVdWqz8yRu5rT7yh1FdjAr+Ye73734fXbJHz1C82GJ8D+nu
l+AWV5UTiFVwUJMY13PELcZ3hDbXUrnr3MyqRrm6xubkdeS813GKHArwoTA1
jz0iy1h9WAcpBPKKASDDrvAJl/FR3crN7bHZSa61AtNFc1V0cPx4xndwpBp3
FxwWMXHRf9KMSxIT0wFzVFZlyGlDk+9chPjgKvZ5tGIUOGUp4MNvxuknhCPv
KHfYap8C45+MiViZEsYxxgQ+rsXaAXJfPCigGdHrsewv8Vqr8msU7H0/bpAe
/XUXUZYvSKwkMjIblEGK3apavORy66uLdJp/unn9Row0JheYdqsWFH12YjnB
Y4uBt0MqaL50CuERqGnSThCSHf1scn7N3GnGqFauX6udCjVy/ifYk0/3fLfA
u3iYA5LIoz01b+A6Mlj6OCMF8v9pERzOshmNnCNwoySvOK6IATJMYQQv1t76
m9ejlIHdNG8kj2G8U2bUy1Jq8veE+M0iSnZjeCH1/A70hjYm0dz4nTOO/Zv+
ZLdl/1y4UXGCERp0l3L93IvE0HZNHhPqAltOCvEptA53GG05lKq0n0CdoCJk
uCU629xUVyrzGRmi7KdAxmc02uIy2Tz7Q1VJqkSFaldKzp8rcZ9vRrhcT04u
dV+Y14aMmrpQ/9csLeOyIlCuDBoN4GKv0uWJiMAob6ih9DE3FmVHmcZ/MfAv
gbBq3m5OLLj+omArMBeLsRumvBH86lJrgIm12E+tG9y0yiyaqOPNGt6rsoV7
0ZL+KEGrKB2z4BvdZw9RwRLXu8MPHD3rnO/ID9S7C0kj+A2pdHhxLbC4pEhl
OgxlQTBr+oBmdC+lW8gWoyI3vOiqEqj+k0jUY4ZCYzeF5BhZvsES8Rg6OIsx
7MtVbOSVwhElEotKxD2zrE/C0+z4MQ5v4M+qcPI8n9Uv0lmZzLwyJ7ArLcJX
sOR8RtXfV9KAv+4cQTYXI8Ov75tdyY2J6HWioNnyK0m1WBGozXlcF4CqgS8+
yYKFqaIPDXHG4AyVJOLIKww5zj6UrESUMrkiuZRwP28ncPdzOJqOpl6fZaty
j2OyXqVX6OJK3Y9w6Goy9MhvkaU1cA+jqQYSGm++lZaaUSgzrwQfEjtx/ETI
LgG2eKjPvEF4aYUcOpN5TqcRtdjev0QMF70e9wOxaEtMrItuDcXBy4zvv88U
WW+Dpg/mjwq+7LDDebeeQN5DQ6J3aQIgjIwoCMLWu4PG55q8w1ISxS7hkqWh
Qq9VUqRbuDpPGVe97hAqNVFicteVtZECyh9ykKTOa6LiTZb94Oht9t7EwrII
yIRHPENUoHXl4oT0vZI6ZPBATQfHTdaC9hZVpCaOAC1oVnkcHtzD6jZF3Nva
SpPrVbXia3PG0g2c3b51Fs4W9ucnb4hwWlCgLNe8jc6zZvtUHt+rAx76lV8E
8JlIzVhBjvRfOm89EPTvZSt9M5lTIGrtd+Glr/o3lMxLQy5kDF74Fh4Ub6y6
xbvxA7vpEsV/JjECbZtcNpwRZsrC/54aCSbmNvqM4x3od5C+kbLzjY0rM0Oh
VUtFIj2o4rFmuVrp5iLHeX1J/R+jJdPq1fUn/ShguakA8KSoiPe4RxJH0j4n
OMwo9OyBAwV1OoeFSGfgm4LRD/U3h/mQU84rs4hgFlwupGhgihWZB0gcrcuT
K3IgwlcQ/6SEQbXXxryjEpoKKtZSjQhlbcpY/TAfzlcc7shONEAuA2L3mrEG
Pu4vYgweP8sp2Yc5jLTKyT5AcvQRvzBn/5t9+pja+Tykep07UdUIpQWnjMQr
1pdiKP/EHfqipAVVgVXDEePDxJLvrpYhcGGryRDh2av4OiT4KJdPy87zYYll
cwUrqUj1WnG1Fk/WGLXejdkEPGcpV+oLc7MMxaBxXt12h8GFBpRcnB3IIO9q
j9Uxfc354AIYd3wguJE2/6qMylmVjSVfJ31xL3+G8RN+CMxIlnESPfjzT31s
bEqxQum8sly9zIQZo9CX1TOyje5Bi+bTJ+s7RvDvy0xcmxxcGkn8qyY203Uc
4gcYdY7Ajp0D1QEn5/wwm9KVJIejzQIC8/ZyPkQwC0P3mhKqWGgQGN8GsYuB
3r4EsAlfPfaJrHmKhSxro01b02sPxgbYqRrK59dQZTKZHcMxsHDVDfc5wWXL
t0mqcP6tclZGJSYHn45CG1PgkXwpG9VBMjfWIvSvCpiI2bMD8qS4BnTHBnPg
L7BE9a13OzgnHfTq6/lc2XSaUIJfE+SujHdSp1Z60ozi53ARKvVbeJt5RpP7
xHaOhKIZS330o/Cre111PcOWNlub7tM3cO308uJZw9AEhvbmBzfCCqR8Za+q
vPAmsz5+zGJshpcjOntGC8AnOJLy0cKIkiTpILIM1aDPvmWR1H7opJrk9neL
cmiDZnqTjF8Ul9fc40iDu8jYQB/m1V+fn9pckk8LW0BYAvv3WUnKqknAAKPW
eExnBPmPaQt9IVfnZbEsVP7ixtFXD+a9iQN6VDYg9R7DByatd2S9rr+AZFyd
geRBIXPS2fBHtfpIW20heOOl4yvCl3nU4uuWPDJ3mcRj3eP9AzaPGyLoBOpH
4aMI3NnjUCSuD/DMpcQgv4IJ/FA/1DpxXwQhcQFS0RIZc6mSStn2ExrLdp/j
Y3M0oefX6qFRUHs7Zaxo/s+IIWsPpzAkuwB784bnUrwrbL5XAx+rlUCT/UHV
tvF1z7BW8Z4BvovhLgegXSa6wdQFB/tbQsztgZuy1nbHFGFmPwsTnbtc/Dnh
asjXa9rKMkZYplOrLeIfyapoPU2W44l6OEADZhG26HLdq1ruZAvaCsa3EilX
fqPsS7R/kXmErx7dbe32SlJin86fXk3zf16Ry2KPpONzgGbGCGxTBcDyipY6
SweEfdAzlX8A8GFPh2ikzGEFpwvDND6rlvpBQhxxJtELDrUc68YSEf5RZ/4a
+9Jbf/PKOxtXSUaXHnh0ZQ9ZyT4cj7JMdG8hnnAKtnKqYlM/Vd2ZOlKgp5e1
4bWofV+qXMCtIpzlthiabOAGzoXnZYHbXGpm1vt1uXD8wavdUE0A+GUjUzjc
+12tXl7Lz+S3Ez7gcuAs1jwvschu0AiVxh8poPQHtNrXJqlVuJ9q1qgLXh6P
nz6xYh/BbH1oTEjOxsyQJ40/bqdoRmbjZ8qXsMb3kzXlMWsOzYDuzj3zfr4a
m+V0Xx2RNdOh/ZLS7JyusZEwBuCUt7R/cqG8qkKiglJ/IrNL87iwmPPo6o0n
YfmGcgktYbVU4uGSXMuJ5bIbg6SKCkcJCxvsL/jqeDVtGADyAdYAIyZJjyRR
rGdyd//pzSQGihVwIQaXgpn0AvqhpXaiYNsDy6rH73F5/lZLDStoZOPrHCaq
/Av6xkVkbwyiQftwVMquUygVFOpB3Vo6b38wdz3iG15xQ8ZkLR1+R79tsW/C
84cmsarbf8idBU66pwwzKITQtff6PAinICwSOpAimpVdWSaRWr27WT71Uyuw
k1nDlx0yxkGryJr0rz/bubof0tRIv27uieujyIm/0W82EV/CL6Am1aMXNqf7
VLKTWJ9sMR3lGoK/DWlsv1puBN06mea27QZRe5SNNoLPHnu64xeKiatRvwrX
O1D2gjxWcahwnaFDYhGh2R5+APglAnvHoybOBwro0XxUEJgZTZXxQXtO9aql
KmBx8GjLpmxvbPh5AJSqZFviYlccELs+oC9ZxXsvJaCfXP5lQcNvelx3vt4u
NM5WU0ZrujQXbOAzxBCS/zb2KIGlSIXSkUqVudN0wgA7QAPbOVLJ4GqWAjFT
siMaNPyCcsTwYoLHv/RYwUnE62+aJ7vpIQgNXtQrdYkbxXnYYcyltxQXbMYT
U9WEuWIwGedKJqFaoeLB0e8xrIBB8H9kVL4EtrSRqgsqWnvLIlqSthEDNGe1
6ug+5OT3nd7NKyJaFb4CUqLy1+qjvNn90aVFyzEV1eTugFkdF2tHltCmGuiQ
G8queBgRxZrHDmgKXcWooxVRsmYcOPRo7FP5cQd2MDUvrPmf/wTrNQggAbPD
U5Bt/eYzSAUpwPTriw91yrxuSzN5ZdTK/DTztFyH62NYcTp0WVa6YlhSutwc
hq8UzQaLsqVrP8IrfzkTobCol6ADyaiahs90s9WnFBa9CKagM4/bwSED790B
fIJIZ08kzT1owX2cea2qtNT/aQavXm0Y7LXQ3tZSNBxVJPsfluwrtqyHGGlc
tQxoe09/0nhftS5pfCMVWrRWPc+QElOoWsCnYazPBolHCrj6hAhXH9Q1ghsL
W2JvBVRsFVTIKhQK63Fwq+0SbjPXV0pQnUiPIgh1VoMxpi+FyIVOQeGZUDTK
6ZUyrTJgDuXTeYRsbVLzJMTAEkCdvVfvWNJmIhfGfX3f2tMP7S3q+ZMShZIY
t47KwCImRa22eTID5qz6wirYqQovV3Gy6qlsUdbOMMFb6AHVxqZyqrEy2Se3
M6ng8q15/GbTTt3r6Kov752nBaVoYjMlh5stXqNsXlitVG1PzulaGQnElamP
ZwTF5pIuKmQR8A9ez8YXCb0PldnKOqT7hEKVjnB/HOrrtkDWi+nI3F78Woan
09i2AZ1vgypTxaBxheoXvchQwvco5MKSzCCd+z7qHo0gB9hE+S4fGvF0yTTQ
QJJVg5VfXL3Z0X8b2Kjdkjufw6KvrKi+bo0FK7PexL49kidw1k2WC8yAPiis
BCSJ0v/nJzRFrsDcO/kgfiRzq8MAWX5ZVyazr+nfW2YQwqIEOaGmUjBp8cpQ
C7GnRUGsFa7CCQlO7/oSerAawQTUhJAYkJS6tNABZRNWfjAH25I7KK2RHGhq
EtY97pNMCVbtPwJo32E1wc8HXLwl3dTDuw372BdxlR04GsSeODeo2yA07Xuu
/ZtosIHysIoONLKJo7ckT9xydBH2aeulG+tR0M0X27lNPZoEYPBR8Eb6qgqq
uwADNIODePIZzA7Q1nm4hp5LtSuVgMrrua1Njzxs9P+kyMm+fjblRvgy8g94
CJkCXd81CbnRFsTKCIJozSQuTRzXVnoLUyyhpbemaQBo+jmYfNPjzQo7hWdw
8kFVSu+CvksDaB/5DVCQ4IDzO2gQbH80djL70vc1UcLfJO3su1Ahs5iUFulX
rVeLTR1uj2MkfAZtgSnwWub1Ep0s8ZwOsZfVRniIfAvcCvQeu/NjTtI6JBv/
S3vqs38odUezR4EAAgweEXoS3E9AwGXulW2HU94C6E5CvqnHyb72Gq3hxVTY
8i0dr1QzTVpkaUeicp9XbuqI6V12u2zp1khUOQQLNdPHDOmF+D23KJ5z3UJx
tFUQpfHXQhGBEqdq3W7ACeDZUeMfPLndeJ+c+MQ4SXbwxRJmGxoYzZoydyo2
9RuDROH6clC9cBRf/rc1T/+UR2V+zz1veJ93Wo3la432+GiR1/7LFuaS+EjW
W0Qs4/hJb6v118c4VTQ8SqDH2CwcGP61c0frcm9XStJE96Clitms/6fY0OhG
kBiP+nzGRPN/SoxYYa5/mipOmdrNABXZVH0ZT7npthj1vFM6UPKSYAagvUeh
ONNVjEzQ3fCkUVNGu6zX2PBbg6Rqm5sAXaep8zw1ZcASpAsLWubX1700IrqP
B8JhVND+kk9Cocycm8yCACj5lwaJaYUWq8WJ0XSXZ3cuxturFzCMYet2zKWK
Eb/20lfs+Jm6ch/dtj2GD7W9Mnb0RPd0BfCrNk3Zdnh9Em0IKg05uf+SeJwK
/HI0rrTMvzuqgCDnzdrw3IpjEvO1nfZ0ASgHUSkIvOtA9RRp7KjhDTWGmjOS
A7lvio3dVzR3m1RnCTyUG1zorP6cD/j4jGIRU27eQte4F3zdjIqoIeSRtGUB
7lKXGQfpl4/I7ATHEkFraEKy2Q8Kf++c0ZJBHV4qBs+oYYFHsPmMe5g16F6F
6j8a4NceU8gB4tkiXmBkXsrhJCi1GZtm6SkIHfK4wYOS7G9VFcmmtOD3CLTy
Dpt/3QeHmNLHJUa/8q0Xa7PYFWZDaSYsOBrgjS0C35wWA10zCSO7KMc0oFDh
F0HDeEE2WGGop45mrFAY+XbsqaVWrhqIxCYw/btKUJCQmub2PV5+rUuPsPKE
WTobL+HKuACKhAgO5nweKOyO/nGsh4fFULTLKauKQ4Qk/n6zatB6NJraHATk
hMKgMLrM1+vjUmIVY/JDNfjj+cOm/6WRnOFIAgGTofK9ShMVnznLXdy0hcAO
GEOWE0K6BYJgDMsoC27FSaDJ7zFuBpbczNTJKfl1vDVdCbHCqIKuo9qz5xbQ
c1tfD7yBgZbchDvIOcLR4Vv24d3JsRoAeogKwmBMJxkzgm2pNsZ+CNtt7nfi
Cxc66iq08C1gA6jhu3/Dq324OtZw27VcTth0xJIgbERm/HeyJc9fnC7b8PWV
5MGs+SNTK9hXdtGrF8BUCkrAd+JDNamNSEaySGE9MgxB6JTtKisI/lJA4dyC
owL0cLw9eyzBYxrOSMvMpUHD6pwuH2BJmezazpnCfPk5U0KVeRE0ZhkcdA9M
fQOOdtozEpVXxa6tClNy9KWxlX89b8TpYfxs1jIrQqyBGnNAQNypzcyq0oU3
TfhubMChQmm/ghMXp0AcFlIpwOktdSApFW39NLsIQSr4epz+2KukcKpFtQJZ
7e2CG+FTBq3XfDynYuQRJtcjq6tbGTpWIAwqx1ztwM562dG6K103qUiCzUfV
G6YuRGuQ9TFAExCQ117k5wMeuzGAhfhM82Ll9YxLSi8llgPpv9XmZu0KinFe
K76aK6VFx+9Jxtj7YINBIJGiWUAJ5JwtW2wAytZP5RTd2+8EQnlT1QV7kEsf
HfAtT3sGiBO75iCj5vBkwRuHUr1x9ctJYCg45oHlMpswW19fVmc/g0bJ+gbf
dMSOtQqMuoeeBx3QEoc6nlEw5R45QBy1PyMlz7GJW99UWW3Nf7FuQDuCvOgb
bddPdD5YxGyIEAh2J5pUGVA9K2wOr9/PmrtaLIDnhQOwbuiaIHG4A5VBTmec
xp6br5YXP2H/9QraY2XBYnXeKiZbHtRqLVRjILP6RrgcCVaIN5zLtwUwiHr1
jaEDAO9slly/89RNHIjLgTKep9knqZoXK1+4na1HPqL8pTy9OhdAYzjn+s0D
pGe8K7vlafJMJ1J7EU/N/OSIkM1/f3olBWTEHiMqrmd8uGWp2ZkTjRabQiUv
jWkxAP7cbM67WKqOld390nQ9THr/NnQbzRTQ7EW3Z8o8w1LKHe4EWstF3KAH
XHj1IG6GPf8fpaSiuGGfYPFEqgh5V1/mNkC4GwMfbytBPSlWvE8ZY38chTPC
KJEQn04b+XEZjRvxZog+qybLB8/3JZLfkEWWAAdMLVAILbghi6YmLvT4g4PD
XmB+MrCfh2WPIoGyKtTc5oaCzJtSr9Cmvi8HZ2NG/NDx3C2U6q/RDtrlPQx0
pUrCTa8rEw9DO8FBoNbRanmM9ucm/uGCRnKfEn8fFzv8QE/BJrdAa2FiauvO
9ZBi1JZwraSMGOwb/aCumfcBRP5PYn9wG9rq2lKDY6ssnVn0fQ3lURZlk297
RvVI6rpWjSV6n/BshuzQ4z2dwyHkcElH7Z7O/3nrd93yhfk36m4CD2llHjOJ
6fjn1Q/t4+2CEZB/vIx4aq6urHAADDUCXfa1bJtGHYqE28LVFofByWBQ0Uik
T1NON9KtvCZXSjGdzEJHcloM5YL72tT7GfteEOSa5nlZ9+gByKy6vV1f9yIm
NICFjoWnAm127luJQ/dSuB8yU0zqHJINMHHDnsvREk2yFS/JSKVXo9bB8G9/
2qlo48b9eTOwdaHkkhZyX2oqTpxayRI7nk+MPHN44dPRpUZAMGG+AKllxqrr
e+Jrt0GSwCB1G9DadTXcMlys30hewVj/qOZiZFmvlGarBYQosZO1PF3jgvv8
580uMOZUVtq3cIJ29xMqw4nqjD7jpt96x8J/5DaVX8WwSiRj60b+d6u0Nieh
vG+kLkkv/q1szVjBUM80k5VPKs2qvgTmaZTkF4ncw33MQt7z7/kY+zTjK/1p
NaQzueLyIcovYzeG3uzAvTLcI372f1gaXJXZMENWFx8lSllt166DKYHQVeKE
bq5OXigg1/zy59xaHObxq6/eUoStkIKqS+ClcQpTLa5gI6Ebh+VXYHAuvuxW
RHMDaTmxqRfDCJSUyZjiHMI0oF96tH2NF8rM2txa4huBE3LcyIHzm/n7glL9
WZInAQfwdLJk/NZmlHaE6tjNev/rINxl8V5SFqHPY6cxr4hhQ0DjlHq/i4ar
gurGWBw8E9bQa5pfJx9Cu6fSDADX3YpIOVquRL2xQoHceVUt/Re/G472p/eR
F3CbqSYtxrKbl792z45ZBrQS8QxAK1PYUCzpwb/5aAMpJ7FMcFtkPoTxOG0Z
To5djAc+qG+P6DQgqk1bZ95Et+IqVlXE/NZZIXhnOOFf14zjkZP5ZKJqABj9
tW/ga8/KiH267XuNQB9E5JLxIOmCfaP6D8Cb7d0jWLSwwHm2gYvzto+zINa1
UEUG+bIpTZW7Xma/tJ3RCVl4Uz/hMklBMbNU0tN0G/EN7x9QGc6vGTqIjA6p
b5CW3XwmEOMjnJ5Zx6zXGZ705hy+85tNXlg5/qVNARErd2E0KaZ3+LMRkGWp
tCAc8OO36zZLUG4nRVvreFP/SulUriAhS3jRo/9aGgFUxJ2mxebbVKZDceJT
ZQ7lc/Kgk2zl8bekQZ+4A/ZvUHFU1qqZfDaXCWYWWV0ap5Vg0Ckjwdu1qw3n
U28KSXPpV+61WW/WrdjMNFD1EOFAEWQyo402ZrjNeQbHx7wlL1YsVxcZsmk3
Bn1nuRrtipLEKmBFkRXA9TYJTi3xosVt3nrlsDsklCfqihb2PVtAnx8KYMJp
sfl+JeMRRT6Wg+cNbhj2BBrsdVYiYXfLRX2kXATQ16EFvBE7Nc5M0skT/dgM
j6tSQBHBH0QVMQzJizs9mpNFe9sRxwiq4p2dLxlJfSc6MfMBEsq88ZYnFTi5
5FJ/8biPsRjBqFcZKL/P2cmfbuocKWJWm/BhXAI6AhRFRUqZJSdgIImMXAXu
g7FG9GLwpNQ+08abzTxcWwySQcxewAApecy+ajzypSaSZDqS69GBZAGLnl2k
W1yJj5GR6WTSW8n1KWgtefZa0br/ag6qfhCtaIMLXHlhMv8ZqqtHoTUFyXrU
qhNizyTAkadwd2TYC2Fp/T1pePipmM4Ye9Qgxlf5bG13k22cH3ufxwBw+iqn
+u9qEPs0fmWZq0KM0Z4bnp5me4p+EE5I+TDVlsqpZGZIaoNAtUBQzXQl6i3b
aG9xMRbyUa4Wun0iybi5rtHzeaM1+CFqy01NzGdYvOuXRjXvqXSEXaiY4mWh
Tpd8imrt0t4giKsn79WPBkGmQ9UJVyPqKC/vdQQ40NZMEgD5KCNbu95QNIL7
u3IhHbYw2Zn8kTQ0nWxteUkS1q7cwAdzzvFjn46f0I7AiMBZLBTWKhcyaHPU
52/pJue1gC1JlDDAMAxPQ+0pxqimCrss4AGYJiqjIH5SNSmXAI6A72ukmzAx
VKrLz41Vg5A6STT9Ev0r1r+CwxVymEonflpmUI3494oDusT3l+rDk4yiLjfY
Frtidju94saJZdST3yxsRnLGAjAT57kzBB/3lLyplmLgHKBLfzdTwogHAV/5
QF/vYn771Zwm90mjxnU0xUy9BjA/N2Uomq6HQaxuRblC+p1aiv6MnZ5mPjr+
Ma0BXOSu9PVRhtRaG335oOUuKEbY9vpz2r+ENDUuDCJtZdyIOeE2DqmLcoIl
14HCi8G24p6YzpkKPLKBal0+wUakd+As10kOxPpoCuQTL3pcfsiE+rE7QvK1
627GpPHozUMfUvP1XfTYwtd8H8KCjWjL/zrWPMREnNt6GBSI+6BH+Z5l5f4k
kwSM7Jgp0WkjZRgYTAJxY0YtQH0gsyIvLchm6Is2FI0STBHH/yLwDC+nIHkV
aqdFV7Bpu0b0iJGfmHCGY61foBiktB5BwKYNX6D4czZrl0+l3QstcaZJ+Bwk
9/x2+TfGJs5lvSq1KVdjE4Qo5mPmFJ4XZ9vUzV0aGo2jWHpzpcgCAo+AGIBr
ayZof9BOMNiTT6sgcdyrTClOSKVg8r2t409p84M2C8nuTJ0IyU40Fe2HlIAC
666OvA5rp+/qwoy2GwBZQwQ7afl+xp6H86jUkExERPwb26M8O05mVvrKtQVB
hIizgAzKhtB46j8gpLm1fkUPSceC6aPxtilGAeX9qJliRnIoH10YAhmd8nuV
APGNv8ZQGbV9IBP7a0wQYAB861sA+gXDPUFR4mf5pYsWGIlpfXFvH/G1s9kb
8tvHxjZPr4eZJ+h6JaOWSXeA06807VYnJ2r2JWVZxacgQnhcyZPGV2YkPh5S
t3KztROk3m2tSUGbF79EPWNvsi5gShPGFxI+drW229KZX1+3k5cfaeRDOqgY
rAhODyQNZqLJDSSv6KYG5USiP3oPFS9GhU/5zIokw98nZdr7o72tEQMzBN1M
xqHpAekYuceQhcrYdUCvivVu7JWVUaevkinCO6Hmm+EBUrkTBx3deE4QGbeg
I1eUvct+lUNV82C0WaqOz3emqlLG/dgBIyE7kqdnWqMt5TRe2nk8mwTUUfvS
D8PhjvvapT2ijvcjUU11ztT0ZuoV/qcb5lFDJ+ovailGty+C75CMDTApb6DZ
bjF0LN6FTT0CjxI26EAkT/OOewVUtBpL8SF15y6QIrokBcZ42+BKjZgM98rf
lE63TYN5nA/Cp5yp4t9JCvPOduGxrCHb6fVfClvKTj8tv/Y3dObkGFnYY5Rc
iIHP4o8RXYUKnwW7Cl8Aw1kXI/AKXA0HSHW0QGBlVDUXybneD44frRYWw5ge
qQ4skbz+xfGH9YMUOwmZLJXj7scsF5GxD9UBX23nbhlJ8nAJMDA7Fuu9ZLs8
z5ZjrjODm60vwhV0fa3OYOv6JheB292/jxEJdhPCW86H1DoIVTJOVDzcXf1s
mAMVvOXNztioBRHJh4cyCairAQRhlnnQC+wXrNL7zw1B9amyutH6ciKjGvi2
3awHp4h2FiYFBcI4MCdeSAXZF4krT593czGscLLAVlnwLn0Y0fWbCXS5r2s5
0MLQpJV/Mkp/iUIl6NuRb087o4RyChH7nsWLBQDLHlWI5EdiJ5ZKiPb8glp2
Ngt9iFvZJ73FsW5i1tiW9SyrUUY1Wq1RVtf/EUjuz+TRqmHGjTGT5kKsNgkC
Tfxf+i5RvbUeiQxVSL2aRQP1UsM2Yp2Viilqi5gLKRs3KqahD6yXayTHTl4U
NZeuxBmruiD+lptADGAsJ+AVJzwUxGOrO8QhxtGxhcI50nEDs6S3t+t5oGNK
OJ2oMMAtw90lAGw9tAoCwHRzmNRJf9dS+Bb5en2xTs5sCZadMAcdSXxCs11c
zhxCu5lYDsED3mIUQOVdw+ZZHFbwJTGlK3yumOtd059jbsr88x5JSF3t60rL
vzSmmadlbXs+a+FPoyPNJBJtBdWTltqFozBuer4+0OYUxLncQfWI3UWoLCXA
Qjd6lGwY+kRWaOjCy5/jr8qOGTqFJCb3h3GMhC+TPUFVLvB6vPr4/pHnLMVz
O4UTMo2u8yXJN+PLbYICHJxv0uk3ZrrCVTqcZ/ibVuWhirnXJJKGjGaELxz9
psKkO0cuaRZBurm5xteQ7BQJGOk/KTQmnT+hN+6+jPWrSa0K+yPv1nSUi9L/
Yn3XCLBUk5G647XYEda13yhYkvTIbhzhPwIVQont7eQzKjToCy5p4ImgcafK
7nZswDQ67cG2/9ad0HydRg7xqPyZaCZecTvCVzKIobm9yYSgUNgqbib7bQtF
MGOUbLp01Dl1j6FSSb6yaNnxDzK1LuTr25lkn9DaakdmZjXNYBPnSTplJUo4
DlfDH0FiKbsxyICaTno+HaqODX645N1buqFgaqQ+1gy50mA3l1vAPfk97o6M
qT2NyPTxMIdo50uKRCnNNm9CLWo35xcjGpCo+QQHujsp5G8yOS10PJ3cTORb
mz16vCf4TDELL/WaCB+zDM973Hs+NMLarj7MsuM6rnozpUILuyHSDrHOBn9Z
p/s6JUa5qn+tool2gceyc5SG0kjaEWg6XB2e1b84v2kIPXJt3VEO/lxFJfEw
OjS4A3aJypc09W6c/RKhtTBmLy17itpFg7LE/rd7omyDbTU67W3Emrc8BepW
rPhQZh7ugqI4/UcyTWrmdI2CvALD0YDVPkMaHTJkO+3iJ3gYp8DE6ju/ueed
Jo8XMq78Ugfd4FoG6JMFtT/cXTM/7XmvpqBWnpvq6mu9Kaf2AgebaHi8bRZ6
DzEqOmKYOkrOC4KYUkvk5huBl2w4OntxlchQr5lleUWEZWHdIiA+qmVed6aV
4m/puoL5OP3a2HG3gY88lOt89Vy2KdvDdQTu1ALtvtGbE21pvlALF3GaZfiJ
+yWoRF6WR76jQb5tGwAkzNB1mTaGH/bPcDaH4Aj4dTL+ifPP0O4KzWV3DxTI
mfZMl4miMCyz1c3sOFRUZWFInZzryBhcXquGGU17t51F0z18JMMI8KDGcnyL
O48Sdm7UvHKQC0OEMakn8bhrKQ6rzT3gwFvPzemjR7/PQunsAxrl/qieKVw7
kChTCzTKXdRIhmbFq6FK3LgN3rzQCh3gdUTkIxR4p4rs4q23pDYwGBVDNn5t
RBNYz0OTo8FwJzkgIrcxSjNKPjyEhANaGZA0rMR1ZHytEPDueRaA7jE0fM29
X6U78ydeCPP1zzek5Xiy++G4HyY/am6pJCRyRXEeapsehvi3wIvt6ZxIpLt0
XwiaREcreii5RP33n2dsEtM5sm0OA7pco708XjXync4USCd9m3qOeINa7fhR
ZkN7pbNlk1EgKXCZGDh6iBc5y2rqCvHK83x1DcCL5hoi1OaYGsAIB8QH7sdt
ze4tSK1eMJ7Sv4SlnGC78bLRqDpoo0w6kZm/twEOiGMUxLvqZ91sjPUP7s2y
DMB3tXYjF4K/MeWPjahJB9cdskptd2SdfeQsQTa9fokuBY+g07/V2eyuy2Or
Q+c8RGUxHRzgIZFyrGHILmM83eiNUYRyJbA2zPIW78Fe07iJ0dNmP0z1C6am
WPbCqFef/ctdeRMyKtMpksjIy9wcO2KhZbQGeSCeUm4tVmr/WTUqmAfqYD5J
k/3O4cbF7lCgIjgmI4kUFRCnw+Uo2amLj57kXQBvhkNScgoMr++850K2NMRB
h60t4Z9owZ0T/Urj496ueSA0RCRx80kTkObtO3Hlj+ekAQuxa48JKh+0c5Tx
WGUE/g79iF7S0VXKjfDDvLOftqvBlnGCQytIWGcXXqIhb/lXr9T6Rikq9se9
rC//nn+YcHxyx5JHiiFiJQmmSVm5SE8ogpTbDu2y1FfrkZEufcKuGJU9Wl+F
BvqJVq819ITo3Z/UIZMvw4eRb0eDC6zALo9ien+O+VNjuoyfp3+of49ju7ya
98VfL1bncVJW5ZD5rzaoJZvN3os8oBFE6/gAUpE6agnyiq1XLMBx60gUJYRS
23quN+DTLEVOxoXbFQFUgNLdxL4HJaaoPLgJbo6btrm6ROsAOCEWUQWA7OwY
CKTcytx+gcWYOywE0ulvy4qwyJInq7FQzfZJKYyfM7BsSUVkKPFoAcXnWkYF
jgupHbzGyJhzZaFG+uM+pXeKjJ811BXvHOz7bvsfjimOASyNDcJLVnVdz8YX
BHaXPyrKzN1846O6icSU44CyCOtOlDNSnJp0HUA95pbBEGCHDFlGn9xBCKlY
kbea21f4yhxYx0LZpfFrT9f5hA0guHrBdgeKZ6esvUcEN1ha8aC0lx4iaezr
ElVkcSXdd6l6zezonnOoCXXQqevmVk/TayPbwrVYOddTn4fGltZYIr0IuI0g
EaLMKGWbB32CnrJOhW90vHYFRuQd16SZAy1RdvWetGOGuyi9+SaULanfajjp
BeceGkkKykR7Qg5vvhgrrnPN+H7IBHOShRd9Yt26+b8P/NcGCrlvaoZOvh7s
gRMzlSh4+i9zpyzK6xmOTHsmn5+dUS46+Uggqeu1J4Rf0tEMDBcmWzMFHQc7
4GlwEV4IW/OPhxVHiofA+RgG/GLTl9nKXqHxC8K61X9e4h25I120S4MLMsIV
dc/XM99a6I9nAObtZ0Jn4YFLkpyMb6dq405iQROqbTfzIIUt1dHozJJIFOw5
cG9QtzcohClGxYyaViUir6sZwy2WG3FsC1dYM0Yqo1NVUkKtr+zvwaBZxCZi
zNF0zZEZHmgcasjQhq8tFmnV4gq89J1BRbSY5QTJwZXYgSI7INvqx5ndeiph
JW33w+lo1kbltMM70O5qHlwLhrVk30NX3H/iIz+XegHdrsAVvasNWWoE235z
KsI9wQQOW1jYcrr3kEcRczsJCXdJ8oWPRqwDBzB1lP8wrhWiB3lQ/oAdzbhU
ShZGyBexNeUgfaeeAgA7OpWDgLa6hPWgiPaxilokqPZdYcN8VGJrf+eip0Xq
rVFdla87aFIa7fHzlNDXGNWjGrNSOnXdtquOFcsAjXFlLy3r/yUrdIAQpJ5I
HsXR1plpDQ9sqq1hYbM4M9GKttySABUhIgDa47V5AAHNC4WjdduFaTTS6h9R
yowsbrhxWgLqASLk58EOTxdCLcQBzcakDPhusg6BcvEnNsTY0cgXJ6ieb+s2
UUlCOvnmKQ6E4pSpldOgOzcpOfE3L6rBX1J3W7utfDgmdXa7AD7YmtVO0VnU
zhWvFrXHqDTx9RL97wkjYnAN7NkJ+0lshu7aXYVPL75ZbmEuXbY9KGjLomhA
gq4kAzn1SvxXZn2ICz+ymw/0KbRL3wzPkQIysR7tXn+CNwLoSj4DMCVlZgEu
tpYoChboQs1qcGssk9RzidN3tHo1h0DG2oYQCvWIRVyVEp4PxYPuwLrJ+OCE
lOIScbnYflE7ZY7e7n79RzoBftHEWEeCC5xBEW5vznOyyTbrKVtFFy5jSHhz
W0O0QnReGNc9iQsEGejdFGkS8UlcsDnSnicVVsNW6lX+lzwiBnUOxPgJfcZM
cDGKZVmhHDrpqmW//SYPWTcILvxnUrIfX4zii+E1b8Cv8Qkq6CE0mXjKB1F2
dxH1yAXyIpLcwCB+QikHxJf2qe+TZ+LorZK08DvPpMh0GrypxPoLthIK7tz0
IToXiS52EjjcOxMJ0wNMBTR5OvJrRJtEb4jjwVZoqbqaZjPVTYUd6X1Y0/vg
bgBbip9+0Wmqz5R5MDu7LSRdzdn1B9IDS6VeCZdMevJBsnfz2HbQp8iOSViV
Cy+5DyfxwhaAM6gMuCh9xSubG2qil3XLJtJt49T1SjLT/7SKajqKbm7GZMpw
xtxAXzP+uspzqjvedk/LXmNfaScAUd8tF5lOrLcvJ+HzTDNwsBbaV2/aAN2L
h7gnR7K70064Pr8GeY/EGqCgtfs87C/WjF33hawyaW7OZB6oDxRtFQ3HaWKK
65uyUSv+Z6Gfv/zkoh2iO2fGU2ejmAhgwqJfBDBxONJx1+V6HyR/EsZf592f
+670aS4p73Gm/E4b0VosCZY4jpiH/JbZ5nr63g9Y5T4FwzgKEyLu6GzNSh4Y
2duZVXjtARJLWD8xbPfUrK5O2jQlnjeG2sfZWFWAb2iADEgxDhkWOSadOuZI
zsUo4xEWLDG5Gx7DYC4mEvtsLRWGDo1lbwki+N9J3zJ3nhGNc4txA/CH16Cu
SyXtjVereJR7DlBUBvz+a+0gTOpcSPEybG23jKFYhSmK7rQVGhIvGy/KIA4o
RVufe/s9uzkaYiqjdAZNtVMuUmgUtiwT1Y/znBb7zSGvH3AEuSO80b3QKF0Y
lyC+JprPTA70sov+05XLeTgnflLYvmT8F/kHq39SkJh6IjZfkCEeeUMIK882
eRFOEkP1pMeTsLe6UlMe3x9U4ymKrsZTi7am5n0oFqBO5xoDG8KhLRp4TIBf
i9XvZQAJY759MOScyp3jcZt3Z8dWF778sE4lnKngT9cDWaCM/DPzHZ3zLjPt
gfPbhe/LNoUS84KjWlj61/5FF7nfDfAbDSmnc8eTxVeOCPw9bO28kYRZte87
I2glhObCBMG4H/h+qsCoS1a6gMXw9FbDkN3WIvc8blcn0rWbkz/VO1FF3YDZ
6pL5QnWRYmLXt6tzdS2lL5mvFxNOavNR7xBAuy2Bk4afM0r2gMkUrae/DMFB
Zajw/WWq135NdyH+KUcImO9H7nQI6plHwjf4x3tfaNpKqxKKgCFowAF/fKY5
aBQ+Wscv2NDjVnJfE2LqBEGccH2U2b765zmnSmoadl/YJQVzFgJoFZ+YmfGn
rRWvnxFCg3vGsd7U2u2M/4WYPfyPbhsoOJa7Jd91zseSHeyt+CBTvl9AUCeQ
tV+2oOlzQ/1b+kn0xO8xgExVaU86ZZUfUeJ06zOvoRN7ngJkugFtdCYGFVyM
tXolHr2NI4AOUkO1jj9+ps+f0GELc40KMO4DQKThZXaXuHJ3G/e92HOImwBB
hP4PmGsDF0P/yhJ84CfQx7HemKh5O/MEbgtwKIWWB4JCWhCEYodYKfjpASt7
ZGsoKSYKPEOUsc/fJ6Wb7l+IwrKkv1jaSqMjW09LTyBFi1EJF2+gFSGQxsXb
/LSZFw3GrFU5iBm6lQ7SlxJhoCFNlwbfOLC8z9z9y4pV41xnLNvDiN8NMNWR
uhRYImtab2TeYPIDFZfjivR4Tx3SlV4IvoKWV/PuYEwcyh6eyOn9axe6FrAy
q+fNk0T7ysCEKduGLRb6aWzYM+0m4WWxJExiXSuL8oDWtJgCvGJJO+sM4cdH
Qo8yA5iFbf3KS92yznsESC6Zqeoq34lSYYf4LIZH/IXfPHXxOC5Hs7AppQul
jMg62m60s+QddnwQ6nwBFuoQEMnQI3wyIo/uRQ75ekdiniYYar2z7k5kQhJJ
PpcQUH8ddF20UJOnxZsgzMyDxUuTpNNQuIMoELM4OztGKRyqYsYGxpTBXl+V
4jcBWDuqE5nu8IW7aryiuKp3OidxXl9apGydmnb12hTQa7X6DKXlwQHBUbjp
nKvIGKWxahlG8en4/Wm9iNzE6eGwrlJ02jQVunkYUhhfcprNNPDx3FVorYuV
nBigVpDFV6YU5qEd3SH0Xk0qm3dJWYIr6iKjWMupqGCFOxwgRkMPYExKf3Bj
x7gonIJ8wFDwPm1kTPfrslyiDUALiM/4zk2a7fG65CCmkTgkiT3RvoCDZGWX
PW4+OWzHvmVA98OqExK0r9w3j2uSg+Qp4hPq6uskI8bm6qDOEAMKpwpSH4yc
2SWQVPSpDih1cQ5P/y8ne2im/Bdmxzmbwqc/HiJe7yKI86CvmCvX7bTxt56c
XOsFYPJhUetBZW7uTsJYXktP0YHXrGtzDrF4L873irtl1mjlOQw6USyDX7AA
21bBlTEcSe7Nee7HEQuOV3R4p2J0LD/dlofUr4Jiofx2lNKfw+NkUK86DQrH
DabO91JrHFYE6trm07/nsxlHZEpZQSYZz2673JbcDkFzwidVOsmI9f/FgGIQ
euGUHBHYXEytWxYW6OBItghU2nB7BHnNLLlc3sXOY2rmEATqUFWD7iaZSUNg
9vnyMsueWU6dRj5Xb6TZ1SmmNax9x8VmKjzR+N0OIOuEqd4XcMV3XDIWw6Pu
uTdSrkSonb5aGypi8F9+LvSy3C1sI6IoUBYAaqsuctOZmWIFNa7QePrgJSUE
9mV2pGRTRXANilqwGrFYZeE9ZkQGj81hRts5Zfg/2+KunOnTomcSv39tmcmH
9tik8VFVyczci1tnO81GbuZ85GEkt0WhbKZ0PaNo1YQI9L6U2Osy+SqPycv4
8FxlXpHPBXSnWLxwCxwQSDKj7aBSwOqYyC0v1L1FrGqHioLQW4d3cSA+BWIN
omIV8pmK6de/mHA8pxwUyxk34N99qSunX2ZtlWGZ9mN6fk52iQMmCthMMUVr
J1TFY5l/udzu6HqOM6Ok2CdYxv0cKOKfMCn8YHOvnL8/Y1LDqxJu1xy47Hqo
yBwk4SdR6u4Zkfqux/NX9KAi8FYeBBvNYSFsnIJeTIdtYgEQ6EzVJhVzN7Jn
VULgFjqgz5/8jnoFajCG4PEzGLVdbAPKa4JYq2KxngJqCyG3Ma4RssAma1Uw
Vl8HuiUOBrQ5LM55xes1VObnVgadN5qX7zT4zIg96rOVvPYbpBT44hoLU1Lj
pBoCxlhAW0GD8X8CjDIkrjpFsr452BEf61n7uemEDJE6mwp0YfYpWqeAuaWC
IJdtNe2xhsTsIcTj3bJ0egkkMoJzoDItGx1NkPFuBH73yR3EymYv5Y+4cLZK
cZ3K9W//eAjq39OdUUmiASeQh/yI1nsL7hPBSjuEdf6jTREFW9JDTOZiEkLS
jvofK3Sla/G68YIzsk+tEp00WgARaknAjPDjbsh/dFXspJM+RzbiUuo1LC3g
TZn85J0z5/zemNlp2tfKZNY+f3UNubY1JWtcKmANLeI2eHjNKTDMXBYR6Z+p
n80bnPQT2JNouepwsPaYeEnfgyBAdQSHMXZTWlPx7Ssaw3D13H3TM+VE72Dk
LsHDU6yHxOIjd/XoD+kESflrnFYNnU8CXIDAQsXIiz9lSP8epXhd0fKE0H7S
Maiqrn/FKZmVpMb5qt4GPcPVP0i5mP+lcJCP84XPe8EOUPJQiMe3vwAFPMul
e47oWJrBu6gw8g+B4o8V6Hn072OFSqonsFyEWHS2+KsGf1MbQQjdhShZDS46
ZfN7uev7jjbA/UGlrC5cnzQrpQsan/uOvrfKRTNQQIr5Hq1I5H46mh5pQKi6
uIuZE1TKXgxI4/755xZX8ih8m1/+uubWRuz3nu/gzHtXdGRx1KkZV1ue9PBa
d0LJUz25616AJ+h6D4bpuWTeyFAsWfFOuK1DLjzuiRQ3bqgJyUlzaBgDZ/kf
1DjNctI5lO3q/6kVOnKGVhdSzlbumWiFyzQ6k+68DXUJ9kytvDYyZzgAood+
/6aw1j1j28gx4VLc6FoLjKEtdWZ/YGmK1+XD9A3q12t/R+KMq55TxdxVlfYA
utIB8nj+J9835WtNx2Mn0pCVUj0SGBATmkHgXmttWNbm4dy3v0YdfVJ95/3L
5J8HMnSCpHWYBgCevLLGq5l8077+bD/fh6i710en/V8yOfL4ETgxGpbsJGuq
PFBdstdweTLtJk0ENE3D5uZtYsUTHUVo9iID1i0CNBRwS9WONnz8b3oeD94p
pXbIuWZhIuw1UYO5saN8og8I3vfsttYKC7yhk6y8LNgCIdtGuQ3A30eojhme
5utXTVwV3Dt6zL+IDnBL/BiVm6gqf8oH0+pLXuNtNzD0stv0ImzpbBCeC8S9
vSeMR9YvoObcOPskZ1QB03ZgeRZBLY1WLgWpKlB3lhK1Bso/aGLpAEmqaPZ7
oCqGoO1vQk4AEnsyArYdj9pLb11nOamy3S34ayWlndrgCOLM0al91UHlU7Mk
kgKL4+Sw53DPC/RQJgvRegefdNlit/IHVOJ7PmmV+P0zZS29hnPnQ5WS5cyq
b1k6sJplLHXNnYHxAzsfIXeCAgZmQYxcEmDviC6zp85qZNbedM2gC7rPC3ZT
CrFagTLUNKZyCfRwI1NBEOY+NYC1E4sz93bLC++vmcfHB58beY39Zzaxstx4
jYE0pfuKJ0pY4wNpm6I6MCUIBqY1Aq968ypGfPCrJ4qQj1f+qMN3rjhUl0t9
nfrbRhV7KLU7HoT5zySaRgNF1P6E3YPft725l52TViqDkoa24s3ok3LV861I
3kVLgMMWh4r/XsALYUbKyfJN8xoeCQ2CiClaUrZyJIn2uPSCir4uYrRzWVx0
vveQkjiITmLfVaoq1+IooES17Vh+LBXgnuLQjz93m4QtSd2ylJW+GIxz7i9y
0eP2+a7TTskalou4qgnLPGzh6arRP1c1Tm21F+QAen0btKyRhO+f5cFOfmbk
k04NV2RMu4euSofLpaTYrngrZZDta2yv/pYwDLDLAoL73RfwxzuXOXrFHnKM
/NRDcD3unfFwoPYYW0lv49LDK7rDnwL1EXaFFVC/0IgzEbpb7NLrdPuEiUkD
MhyzBqdj3szh/X97RAWr1RK6BokFE1QxdMbK3Wt0bxGIjjT29NayBxXuUfwz
6/Oe4ttdjK8cCDRUN4imdhXQTwqRBPIOgus+xlqwpTetwsiksoSCg9kjuDZi
/DxZhvDX7m4Slxd/tQ8Kl3htpqpfEes1mRG9gR4XuvhjMQRUmg8NuBcDz4SA
y9jG6kP/7xc21j+U3nhAcZHBHQVyeVYCROI1gNDkP3WaHFKHB7QrDM6Q+e8d
C2YSOdua6CVimto0H3oFuxBxorTSmnruEFRruZbnWXrdlC1Mx5b6oraxrzH1
Q9oo3ayVhv1jkjBsJQiezcx1DiD0vissCFPFG8v1YdDNIuIlJ6vNTA8Fiuus
5jA1hzZIEt2D4zs0pSZXcwyDdvwefhfHvBnMVWj0NfGW9emaVKlVf/R+bujN
1MdOFXrZTStjt8cM/6HWxHym5gYeFnunh6vjpp4Tl6gA9IrvCY1ZzrNQyeDx
AAA/rWyYCPltEFO/CuAKgWWC8PHSuGeyQKu27xQj8Lf8o6xTvbVqk/PuMsw/
DvXqOpzF1LrHs1ykq34lHJ6c3G/8KlYrbJ1BFKZB+9+mcA+IehHn7zaaJWEv
TO785SJ/jX9mKUzyQzQZkdIZdRKUdcmZAqHKcxFfH+Q3CwqvZiG7pTOx/O4p
rsiG9yd3At3aU9RoTLrrQQAENYMKBiCqIWcdR542IUqS8JHFpFIpY/ahwnhX
FqSGTtRMuyR00QzfPLe6kNhCMfwzuptMieCL10DDAJQZTW5btwtoeAKxa+ap
e9JfbvzxmK/mtoKFlgABcRHwZc+JfwohB35HHg0TvNDO4qozDQ9pVGKSWmz9
5+0AzyPe9AWDzahrDYr4MOHZvXRCVyqESYAhiaAsqrGpowWE7Whk9dKWcNU0
SJBBE23DFtVUPasC9kdU1l/950z0nvYmyNrhZyEry+JRtyI46Kt4j1ah6kYI
J1aE5FFPllI+M9P+Orbuh09R4yAxNEbS6G5P54Gh/Nd81ywWeUJP8i3tEI51
9ch7qBzIsdY28jkMYHkpsf2wTCBmcPCxsqbJ9XeAKWP6QsPVjNpD1Bym7/pE
LzIF/zf6Fg9qi6AHawvwSbkS3H7Mrg6HlSIhf09ycqxXnmGNnmrSPleGP9rt
MgXmCw/WJ79tJIp31TNsS05jhxjkxL4nkrzQwPsQCVgVU/IrlTehbEFHkBlY
WNBUvzfxuD4OunNyC3eOx1rOp6FZaBJruuFv3cCX4OXkwI3TbA1mEOsHzBwc
mfw0Y9puQqHlUf96wEReOcUQAgtosx53peQFWIZ7qBzbFUOj2LlR4cIbYk+5
YZKQ1lydlbv5mOXx8JyhbaJPkMxmv6Denv9LphovHV8ZRTcMXoLzem+XHVPr
/XR7QimuvYFoN0JjmCyReGrIM8QkK50KycGi2XfLCBiJzzxUwT5gxsnyNUFn
2e/zho9w1qD8dqL9jr0UlnsRrIU9WrdT9XGbPSWF6/dIAqmSqDXTn8bKX4YR
XZYLHOLiroTJL7IckbuP3BORlExlcZ/MIfdvytRNUzyT6MqQPJGdwSgEM6W4
iePq6r3+neCLYau3BYLGyHRA0GnMkpZU6RtMtWAxHhBkz1jWRkj9Q8Bckcsd
DemkoFEY+7fO2Tfmdtc8N7ip4/sJm1WmvdPzpOz5x01SUQGvOCK+iwIv9eUT
Ca8Makm+3QYARgg9caIh94/apgg7zOGBKx1+161LZV+HDuZrSQgiK8jHtMMT
smxDOYuq4c0cUhFL8Q047fGw5MBfCYa+gHO1sAVdOmAZbeDhSgQaOP/m6I43
MAoEcIEul178GZesGeh1cmOSWwAnj0ay4yTRv3xcbK9iA+LYRRBI+DORlU59
TjNS3nNoqyqDnE/19mRcwxr/IPdCeIZwioCtrFA8G6kcqRFFPAv3FcfWjn4/
vSHvYKgAuHuNz//AxJmOgdUcaqPIPl9BVP4MMAP5ZM07HrB2l1rhJbSQq3m7
0QoW9G7ezaP1Z516IDl1ckGj1evqxr/hq9vOAqy6OONUhtE3gtPd0pnKWSDG
HFiubUZiQmjUnjIzjs1ytAjneJkszQiEt6wMK1lv1CDmuHj75EWXW6EB5iv3
HuCEDjb2PFFDb4+aTzXC07hb304YLTirmh/SeP4XhH5WdhxiOsEN/6FZwxaJ
iF2DHwwy6j2qi3ydzFlvRQW9di4qAIjjx8Ol2djxx+YDuU0GQan6zGvb6Ika
EvE2pzER6ObemXozy/bRQd3qQ/2cRX4nfvIXYD6dyIOzVoHAWggIFv124wVw
ZttxSv0yK+Zj4Mf+Vrn2n+icOHguSwKCRyB4v8G757dth9SspoSSuigY2Wr0
2bO63tc6sNMeXbG80CD3sk3ShmFHmEEXoHqBI8vqaIPDyqJJQ75GUBj4lRaY
kgvLnm4Zo2J3p3w41LMv4ccxDuIc5n8Dwb0E2/UV5CyTYY5bzzvZQUvWjf7G
KIyIZig3963ktKJU7uaPx4xwl6rR2OAc6zdcuN94IXmcik1q0vZmUqZTXqOn
KP5a5oyd1v0br8eF95AcqsoYPh5IUKaudYs4tx6mLBy0+KoEKcxM7b1hgMCk
u6/fUTlSicYzqqno+1anlFsJ7TQTwB0/i5GnUeWyhfL6bJmfpPvaCYEMmMQB
yYpvnSV9pHMtxCi1p5+B3EiGtyGG+9a0Spc4xfQEvT4JDAYX3te+AXPWSPh6
DrvCiMbnAIZU0odpmqPzsyCKe5vl+egQHixQqn+MgsHd+By0jnNX8iOiENAE
FHvVcMRlq1pjQZxoiXcAve/kAmAOENKZzJFdzdjntEwPQgK8hCRIrHmC3+e2
OiPrfYSiXHC2KRofatM+d2uEvftB/HlELEEACNOiVTNhRbQVhoZSJ1YByT4d
tt3M/cKyvEo4iZF07AcVG3jXVEO/zn4f0dtX252utRHflADMLBxpfMPzgZCd
gz7KTFtJkms0Z0c0m9cQNQU/4zkxylFbJsOAYT0/KNYxdbmUemVdv8ciRIG4
78w1dQ0bDHTF7mP42G+vCRDHIdHyzdcaUYwyCSlMXyh0KgMgetQQeGgbIP7d
HMBl+JXiQmUeMLGKK5q7Gmt0esxSXSKiPbVirZW8f6UkNUDfqXsGr+2k8WVK
rUReei8zQfBu7H/InVBJcutTOk4Q9UYh0KmWRj0p3YtkYRXt5gatfDdyLGKm
o/9eJsOtllKsOM2pMd0ti8Uc1l/mUCXPrFVvuG3jtUmIgX/2Of2xL8M0Ok/U
M58V3VvNt6LOLF9lESEKQxSzjbzKZWihuHJJSKIV6TP8A9fu+2Q40h+l712v
MnIp3dWK9ZcYfXHinWkCV7wNiXA5evBnjl1YblJpVtNfEY+C3J4FLPXrdc22
Xb6lwsydQRDDI0uJVzwdxp03QZj5C3SnjBGeAfqmMliX+LtxCC8Y6WTzUCGL
r/HWlM09XWEmnH0T7B88q7NH7G05ORQsJ3Xg2odEA/1xK8erFwNhwNFMlmfc
uaYlP2zp9yeeuvIGa2bubj3QnBGYeo+/EkeSe5LoUgV2IDFvd4XjNhvwaYb/
sH8FgrxvYCLL7yMhCC9h53eV8/WTA14v9NaBuqzczUILIRv64e12eR4Pkojl
f7nDO6+kwwyVg+6Oa+D42aUIvckc2C6INpOJ1cdM9agpL3lnap0sQMXE6DMV
TJ/Gk2Q/coECcftvaYswwSRam7inoETTT+rMacB34dHthHj9Z6qVnCPvtRpP
ZJ/KgDpMwKVqwOHA4ihnL3o2uhxzLunnj3ErEKg16N5HPyRQHTWAADB1brQl
5Dm9yX0IuFvldxTxtcfXr3jtsj/h3X5zOTy1L8IpJsVYCs+GTyFsd09y27sW
WTkPNGDu/2TBvO5HglnovukSZD7XYn795BoiADcl9rYosHwfEcU7Q/xWSw+G
DxL8kg+JJ0z/xirOSo9tYJMPlmqaxw7k6KotXjyFIA6Xq1F2UXhDWC0UekXO
mJgWsPTGYkGG095gHbkLATV0OL+1SK2cjoKadkSnvzrL23RWN4iMqc+RLFPb
TF2VB6AyA1WQreDCFkJaEDx1Mj9W2oklnxwXjRvdVF4XImvpjt1KM2K4DNIa
WYyJ2DP2f59MCHvtR0m6Ej9CD2HwYFNP7icMQe/JQ4qK4OHUaD++gJLSLUBG
cAfE3t5CpBuFZ5RazCeG8x37hOpGaTjBRZgP1EfryiIiQIzMAtRWw8RGZt2F
W7SdlRzECvXKJ7ecPq2wKEZc0JmEZytmMH1k47lkm6DdGtcm/J4jRHIlKdSb
4TRSaTY2tCZMlgQoRv92cXZT1h6U+Qfjv4EkqYrAjwI3t1caLl1VZbE4fHN/
Mex/sltvaX+JwWQgCOHlbz6beZjYOIIO3K59lqbWiY+ikJMGAkTnASaJHRsI
ZVHnLAjr2zmmbSFL+a9wwp4HeYjvP4U0GURFgK0Lziy/5YfM7Ew5iZBooBrI
dnYOK1UjWnm6XVpAv9i8NvCg1T5uz8o40+dD/BsKYwDMlNUvHD7T5iXQN27b
Ie1qpWE5phqsOFiyJteHtCQEiI2I/qOCNxwcMUJPaJCpGOPyX9XPRzhsjk8C
WB9wqibxqngPH83R6E2n8YwcxHyDl/kkEmV9tP3OfaNa6JhlOupgOE8e0gry
3/CgobXnE9+khYt31G+GVrjBdsOLTsEiBWfaS/oq8SPzRLamfAgMTKMXi/jO
vDv7TrKmuDdpxBuBHc9mGsLts3VZpeQc9nnIqAiqSOkLE1zxhEcuVatyUoUl
9wEKGIKVN69GNKD2lHOS1JQ16kjcwO1N07D/Jq6KEXqiIw8FfO+QlGOEpX5d
jyoIIk9D9G3gDGGOfMxssiXeReEQJjh0KlsHnlfHu5jHROfcCwEMcFuT16NK
WNSk3soztzUJ+dArzC8r8FzRVybE4Bb1MdNJL1Dw/RXcJ9s+dijqhUBYcSXx
90aoJmCrJMmxoVJqhv5fSzp+ZONj3l+mDEZ2UA6iKhKHsgChAvUpAzdOEbdF
OI5BC08YU/hOPAqTS9HNImt3zJH/LBh6b84XDvn9Bi87NZyMTMGlSj9GEU40
FEaK/bj6tVM8ibiib1V0F79dst1WMKI2neK8a09dOtgP+yhIzX/3+SJEe0zE
tqUzLouRvsxsLYbnUD2MqhcT/dF9PDwg1JHx447IdE/Kxdfi8FrVivDht+Wr
tcdHHYJoH2ayd4iz2q7Kbeinad+SQyfXZczBIpEI0YQoCQD+3rzLtCWMhx59
QA3jtBoKuX8Z88jD9HoO5pEVJnhvUA1bfbiS7cs2ZDW/WJMBbUt9sB6Dl9Xx
HbB5mGIROljsP9Uc6QZttBZVLOOJVskKuHzdHFAdQOttqL9c/YCTthjKyL6j
ZgR5MaUezBxDP4GIW7/ZaYpmnGQpqM4lGA9Gf/AHqx8yWYvFdVXdcxoR3uKa
7nlLCgsJWnTqcoZMJolvfH7s5EFRmv6/JF5degUXPWi9egwxZioJ6BAO52MX
duynYeYDlWup6Eh97HvAEru+NXDOmGAdsTC2yja3EyFPTdi4if1MaBjxYSFX
IG0W2TN+9wbluYOwKIWdrHQX//DVMDWsYi0RBardREfi7pSn4g0WqVO5Kblt
61I1X/8iZidbRtuQ3gFHagI7vvh8aEXD0cQUbfCLh/0YBnVqAeJj+GGTHnXi
2b9wgSg0QMLNaaKFI0Fvp3stbY5fAZzTxTOXjLRRBPgMOUSE7oFdoWO5TpVw
z7F1TUnKUixl9RQ4jFs7mjcursfthglMtOD6zZ4atnqlxqG6HkbY6ZRwbckk
TTdTxTJ8+iq577EyGhsPmWPfUPxSEYYm83wahTplKQVhS6eUlSONxCcegTax
nSRr+NR+vXtF6A8IjpG5+QDwsUmATD7dp/biJjchZ65rfVnU4OM13swxQvVD
NhvmHET0wkdr0mF4q9jS85avOpGdd6KN8E9Auooo1jy2ngyqiy+/PgTvzWn2
ls+EdLnfj34onnT794v7VdWB0OE+cQTdStD0GIlHG1kPew57XtUdOnetMFaO
JBD/G2O79+pE6yFWN5YBluJ/QKKJIlM0ZlvjAVsZdAyiPNtCo8kpboi13ZsW
8hUJtB9fptdgqaMSuOMxJ8ov6KndKdhAFd3aq3sbjhmSDPWvMsXBldGoU2/e
45nqfzE5N1OKLzz6GCUanspE4iypuJgOCsAI71Dl4zdEow0yQkfjpvudSnpb
zMiPltL9Ch3go6PuUfnGXrYHuvKAs8uoaLToH31CBOkc1K+Okn7fjM7rXDRN
g7w1pZZMvMlnZ25H+ZdCeAInCL2A3BsOuWEP4VVIu8KEN78uEof4HTpxqH5e
ssOLo/L580qJWVjRmtkdg37BN0wOmExLTxcP2R2ME3cpvCXDVQHh7l0sjsNE
C9Wwd8id9P+lZfntRxdHJ6AKIsJJgTEx2BjtLhh2NHI7mBLVWgH2mzgVdm1v
D4L3/FBnSynSs4XmmfVrcq9EQBR6XuA1CWPs3ErozFzimFdA0/cfjHV+0eJL
6GwwbKCMbjeVYn9klb+NsX5lxld/29UUWV3EYXqazkfRnjw/5KMC/AjtiGDX
kQrdcC2GC+tSIhGc0TTQVA+XK9QVZ4ndB4s/kTait7OIFelUVC0jmVgOPex4
uvlUm/MM5qaFt19WCLFOlJ4rxMZcKEu6dDOrQfBz15ON/AHoUeL6qH83ISQ3
poGLa1Ki8223qmDsfd4dAeMwxpuGRJBWxuaFW5rXed8Hrxlk6MNcxYZhNurN
MKMdufypRXDNInD8iFaq8XiiFXkhmwBhKyatsCzzh0xyCp3BVWKfL/k7dj37
lPLCkGz9YtnClTviRsN5SDsf4OqwF7m4AsvhnE2p8WQ1IYVswZF/80s9neC+
mwJPbsAvRhgIaTjhMx52hbtTfZV3ySr/71185EP/T8/Iw7m2y7ps8DrZ0FMA
YrU1SRZoT5Fh1xoM2UbWCF7cQqU/omsk2juSmuiaAWKSxcnNhpOI5VUwRLPR
5GPcIQuB2nZm2miO4UoU8sIrR4vHPPZS1QBnCX+cDGdx+Qf3ohQ8ayjNfoIx
T+eKSoEqpEnytvZN40cRzPZYmWxwNPPnmRAt3IFaUF41olQvGZhp0byEL4//
LnB+GbrmG3K6QYDP5+WeiVf4VpBNOqa/5to6xoJli/YgqV/NYl/YsDAOiLlE
zQu3ohdPhra2V591eNuWtXt7deDQRfZ6HhMqc8MwY3TTR4IEuNEMVk3p5BCZ
XiRph1W4VEK4LasE/xaY2lSIRa+isUCt0E0N57CwTsa3fuRjE1trAqOMl3d8
reZA7t5MbjrP33c+EQQxqAj4peiDAJl9a3LwT+iGQWHVN4CrmtXKvnG9JmQw
tPWOV0z9Wc33uw9ZTaqmG2rJgGPgivQGVo8KITdUjuFpspe0C0/zTBLb1Z3v
1jaDbcsJmoSXUHhf6GTrSMrnu3OM00AM6Kj3XZMKe7ak+9UwQtmeRDRHYDMy
HiAx5JrwybgsTdnSi3xFr2gsm9ktFRQCT4t/WXGpusWig5DDMfN4PlXDpol4
bL0ukBScjy3KxKWrTWWDi+vFrlnl7spw1qKrhZE8HdHhEUIyeVx6nRi8OMwY
rLwGorSb3fZCQQ/3w6rnCDKYI5Bm4QRlcBKwHyvQS7zj/KIj4IAy0pI6QSJm
A1ySzMEy4MXKlVzQUj4oEG0GiHBE0mzeJuFDYVwuiGBPOh9Mb1vZachg+gDu
pNIKxEMh3v8rZZgMPM4eucC95sSTcF4uP0/MIGHkHIylIAvkKrHYnRHmRDCA
84BsP28tQLSOp+NtvszWl+IyjVPQ0Nm40bkVieNaYclurj3VJb86AZrcz8tx
mOHwCi9MWMRM9s6tVEAXFIdJJrPTtFwrTEl31gOKkCU2xIcgNz9JtUm6q/oc
X6/4ZyPB2WMxNV1kxl8rNjAJvLm/nT+y4yrHxDUZr3b9SUfTX9mYbaf1KO7p
N+CvT+XLh0/bTsvA1KDNCRo3IoOE30KCD3MXaAilougo1fe/vcRAwpQB17Pu
X8/QB5i6CWzlV0AvqWZLoNt6+CbMzvKqWrThWP4NA5W5vYSakSCe09diyw+/
7cvJTYeu0Sv988iKR7A8v6D/kwgSlC8B1oHgpsZ44nZX1nVNfYYf5rGBTAX+
JYWGePexV8g2OfQYRy8dlUl1ksWLzKb/LZFXNbkFS8BFplp7q7dkybpeuAKg
WXFbFPqj9I/nHB2+aj5kN86q3tixHWy78cLbceCxTyBygRzoLcnWW+ytZjqG
uBsl6Fe+vSrwMhJ7Fsd/yiOc3dFztygfQjLBMezxU7OfdHosxYdJvHeiIUcg
LKKRaoQkgWNsARqWtbPj1OulfSl9NYeWtxnQhC3wB8W7XsIZFC3eSwqIt16j
ujicHl06bjWxQhMJxdHvBRm468BdpdB0/M4FPQ0Pevm7/gEtBuxfFjd/HDRX
Hdr9LD6zI2iKdrYlATznMLn2afBqNBx3k+V57adhSi5+q4SBNX3+UVr3PU0g
zo2/DhWMKWlHvhgGZSjfBdo9jp7a1uYSf6E7R7ilrhXPaQi1sQ8zBZaX3bSA
iF1hDXbnOihjDygWSQollnP1+TwJkg7lYSB0UjB7ekSYlD7Kjy1di0n23yNI
D/bfa6j+dhxTNdt6e79myf4o14GXpQNUzZf9OU1F9XcMO5YaUHRPV7txabLN
LiQsQY2bHdfQtj13ZNIjdc8tCM4biDs0c76IQa+xZDXbEAHcl0T7PbTqWSSh
8s7/e/n+dRP0J8LjgpoqnMbFdiiyenh8rBrsP7OB8T11+ZbC43z6G/EHUJOl
znmnOD78qlzLwcC2No7fmb18qC12N/HlEtVssHCRZrUfzNbKaQ/PMaC52S5L
khqcPi3nuOXBlbX1mZkK4i2R+q1/syi+R98rSfC877DIc63GngqPUL/tjjV0
Go+MswGceKjCVZTIYmqBgiPRxZ7ygmdGVaqNalfq1yjOrZQTRrFMKlbQVG6n
TEte3SP/Labz5UyOJWBcYYmV3lcwizJrlgC53y4sWLNM9AqW0r6t/rg9H0P6
iXF1zy7hzvnzF+bg/yirFl6BnJHkrnANMX5jzwntUh9B531+S14YRGw9CqMt
8MI8Y4N1X+Yq7B1IhubssxuKt654+pkMhSkexKZGU3aFTjHpw/rQLqR5h8iq
ZH/dLbWG451ZloMo3eHqq/uZTqOWLjqfGb7Zlju11nry5PIzTEmVdFJWsHS/
jwJKI/KP9p2kXLomhICymtRvIjgDrIX1qb7dHBwd05xHvO//uT7ElKxDFWsA
EVae426P5fQr0eiJeiFREh+cMAwAv+O9fxE5BgPtwh999PFRl8kw2H+5fupq
FcudTXoz+QfwZ8CwcqEqOTrsODbiSULg985Fdn+JpTAUvId2f7L0NU9p/czE
/XAyVTZDhKtXnWYcdrIUfVmM5r3XmdXZ2RLJAFBg029MV1Gcn2jWnWoRuDTV
4tiiiOFttyE6H5eLT6x79ML0eF2fy1nEgBKySBrYNUVgNMMDwcSu1PCUSZnK
pdLs8dCng5+yFx7iPDq4DnNmB2/FtYZhnND988UFuMN8NGk3fh7IdQl4/Qm6
phfP8cY8vnhiPCXbcl0HWLQjajIY1iC5lCxyPAw3IielC4BXGR4zdTXDBpf+
VAYoL8x2LuZOhnz5dB4bVVaeoUonS/EvX2ATh1WGA6sbF6nI9FetwKiN9B+u
QjD42+LvNNgh0OSpxmZ9PmOP0VPtBfjR48LIOVlQw/poGLGfN7iZeUffxdRt
1QW8KheBYO3dvOWWpbpUYRPQ3O9xcdw2zgwQ0R/DFjgFQrVnZb1p/3JW8y+V
u764dGx6+qwU/Vzms0weCG1Mis/S1KFiCkf5NxoShQ8I7IKmu9cA5eRacpG/
BWIvGLJIaT4Xea00wUTqFu1H0yYJ6wFWDzU4/Ful9uZqLZzyEYzLaD+2HMXU
lP3ofrxaFgRXEByhO55oZfhIKDyrxLW5xhlfB3oQImcb3B/0hNlcrUfuE1vg
ugffdTKp8jXVWEhavP8cUltCwsnmi/H6sQG0woEMOvYKMeQEdg4el0HntPzU
uaRLNS4F/TkZ8PcvmNUDtmk4FpBHSRJq2na5SYPVBDWiNNbHAnLI9+vPPVnK
mKEtYNFTqxtqvpK37eNdxL1kw0BRtyj53KDvsMV1aLx4BrbJvTVNGNMshws7
QJy0ix/Z7bB59ZIdYkDk2d64+M6Qt3Zk4R/385OtO5TeMrVkD1ZCDt+T7Za9
8IwuPBKZoSdpy6wtVcNcUh0gk8ScgD7U63ol5/kYziIEBEdFZfV+a1ESebGz
/4cOwMFGbY0mzgyJP4CySlL9MylFBiv98hLOvyBL3AmzjEaWtHKh1hfxi3lS
X3BA6eoJZgmS9JzgI3IA3//aWuDYgyZrb9V4dcGNwtOAlX7jPNq14m9ZkGHc
y+sZVw+OOisUva5OOd1mGVRwjujTxp1WdNFnFw/rLfcwTAVueXmsrghl3Rbh
MUcpZXiQUgZajMu3d4zYEXT+pd/4yL2tGrciSUXAbjNF9wjH6NNIW77828KP
gL2frTqEUJxWCvnXW7w5xfGahFmHUWrblEClYALJuXR8FFIfqTeZMxFzwUaR
VY5dCmnlCL75QPZDnLM5ZqQ0IqN0EEZGlPAXIpdnIInFLdDBpOEVfvgRFQfI
hpKleij396Favy1DrBAZYMze1ebUHN5xoU0USD5nBryd4sBg16yXiej1UCoA
Y2+gCisph6Ju3KneSlqaNHgd8rQe9VowUGXRCF7mLF5QT2EtWTPug0aUtnXw
qM9r8SH/phWj7g4p5GhtTiqfGkKj0RIZU7l9mJJH5iMKlZdolRqnGMYOfhBk
gXKCJKFDSnMt5vKTZ59KRlaYQlN0MtsXbPzKWoXCJFmtK2RY4IMIrIPgS+c+
Q8+OJRA4hnpHUzXGJBhUp1KkPUrcXwCZv/CtYVKz2R9P8HPKLkHRQjQ2ffez
eD8HD/Axk7JPOjmn4fiAGwdBdunxDmOg4C/6QVGkp9ZgNuD2UDMzaoh5IKAM
qMEKmheohd4U2UiYJnrNVwoj+RMZ9Y0Ruo+qXucBLFRc8fpTR3qd/EcnVwNv
uEkHpiqLb8937AIAbYreZPbXU85/50IT458sIqmntb5QIefk7RWueQEywUCZ
pOWDRs5Hu6/RXQHJ3Nmm9QegVlIGC8LZ8S64VWPoR57jdlhe7JCGlB1EaGUW
LGi4QtYyh6bicVdcoW+/YPVWhoSZ16U4pQtzqGwwQVrMCzzNf7BZVw2hCWm5
2TehJo6euL0jVaWnvMdr5iLsd7RG6ylcDQYwZveZ/74/FEPFLEyezPKiZZU0
XRLy5v4qNpJZLgZzXJ2IpO0jfVd7yTAmnPJ46CwT9pLlB8VJLKMujmCLwAG3
4Enoqvix7VkIF0SiXZ+1fN0LaU9kIp12PqDEssO4V97XukTVoEbFTcwCYw50
MLsYPxXhm/lLQc1AZGqdwqxE83yIizw8KcLorUJmNgg+DyvwqpOeHGMl7V14
iQCjK9k7x7O00HfYIX9uX1R69NMvyMWzqB4Bb+FYTW78TgpEZzZWpphLnK0G
LLDsuTif3nWmx9O5fDVrP3ov33nSucaMn0UuG9CTGpwfnPSvX44NdiPw/DRQ
O3VqBBSTzQu7BHX0ImRpBl3u+u9EE83niEmgovV3cxf4qxE0acvaTPxF0MBk
uPFtTMrmHht1gU5Eyrqkie8tB7/s+8NN0JfiafVnRNnHCkl7Ymonx7ADw7Tm
Y+IbAsQGL2/KNy1UzszFpV0Szg2XYcf/RWAGYzKu58YFqMnuZyZHNESRIsFV
1mjaWkSME6XKCMQdKm8FBbP5CdaKe7bFy/Or4/UeVKv0/nbsOrRM/LCVi2Ey
XJfRRMFVec4+xU56QyElfZQ4NBxOmt2nii6SEMfALXa69J7YKf774HriH/8/
7AA3bu0DdU75EsfqKU2fJArB7Ml6YHSFPCL4NPHiHFsKdqTiaxMMGk4k6lBt
4pDMo8KHuYdf8jNsqD9lmoPYC1G5yCtkH1EDTcKIchYiJOK+h2kf1UAO/W53
mP/tjg53NKXfhYUaKj6l+hepeFJ4ExFiswvCOxDm4KYReUjZPXlMiyjwYef3
MzgVbXksvQGT5tYIErFhK87aBWtWek1mZjQPpjaODCH3mDVh96wYnX7Xd8cd
fKewDtX10YJrPwvpy9/VvovovhrJ7P7VXK35aIC2JBsEdUL7lC3ETCUlY0FW
Vc62TABDj7ZLon3hBCVw8Hg5bdkT4VuBV4cZ5eLBoRtO69go7iyueNTFznMY
Rn2lJZSP0O6nvQm+dMB/d90jpNmm0vPFs1IYSeHtQa31/AeKyiHB5YpRWGQU
IyC+5ZNHT9n/BUk/QC5ECQd/1OOBTHIgTOdf0EfV9ruM8QJfsdb5l7YEIUOA
9lGc3C7iyjuw68BDLSoB6CS9a9Qv2Zps9UVYxe4++H93wO4MpRFpOYRznulC
L/miLqI1bKCBS/whEzviXKNvCTs/QV0sqJOlsB8hcs0SgmyJo5I0EwzMA468
EIzcOQrcecRcekEfC4XKIDZrDwrWPQg+XVsxJxeRVjxSzTzlbfRTXiUhAFIL
wKNR7VRTtVwuEh0cjFZ23i/v39fw0yrcJ4wYf0F1FvKBkKUfe/4haNyg3MoG
uz0mKFFjcxNdTLpCme0OTG2QDpuIGz6Jt6BhQQzgxxKnCFVwFd+d41Lj8vmh
S+Vk6vGgR4WGJ9sVrpz+ZOEVq2+jF9jSwByZeHeiq5ccYTpKoZhMflCuDRqO
8lhfFHJoG0GrCWQgW910Ody03CHRhiTWC4+jt1e9MXdtoQngOYrvyczuiOqU
2slx3i2otfd4EXCBX7o4GD2i04K/bjyVnXOjGNdkDnd1Ce08zDbv78LQDBzF
HtfFZatZ2SF3WrzoajlYYoSHm3wRxQ8IpXvj4Irnqxdnmql+ueQTZqIx+MiI
x9NVFEK5DOtA05auGIF3KLS7nDELwm1GLklUz2ExvceCRqlhwn4TQ7HglViB
XXGCBOFwAb0GePbG++w7w2YG9hfZQ6SMDTwFAt66JLfOpt8vwAcDDz2YOWy6
rd086YDmThxCftf9Y+i+Z2W/ULJl/OFIugU4FsJmAv0mzwmAUoKkis4jWoSd
4xoyGRZbChEO3QV2HyH+BfN+MP+DHj3L0RlESM6FLJx5faiRk4/4HRYee/XL
9/FfdZZSBg300b99QoVq29AQkJ/AJ54JhKW9fAjcna7TyJ63HMmgnhNlI1aB
n00jqJ5F1veT7WZk84lvzl69MoAgwSYo6qeIjhRDBfVr21HTXzG8hG0YQw6Q
JTc1850NxSIdjKIxP0yKYQvL5OfB3l7HcuwqzziYz5fWoRp7U5vdcaHABts6
ydqckz/OrWSZqZUC2QwNaZ8eUWaa/OUmt4XCQYlmcsKfBqU7qcV5NrEL+qqQ
KlKlWaOhArjQlR8oCOHwtTzGBtRjaF0ekaFZT5Lt+NAx1F48sVGshp9MNnOQ
Ga1aTF2//9jqiWXKWhQJUxtdif0cAYCHuXa1TbJxtoMPD7S0/W47tJYxtfD4
INqOnwCZa9P6NpHNsWHa1JjCyMFxKbAK7jtmXY4TOx+DA1CKrnTMxPnHAZ5r
q/KYHEIlQ9zotk9/4wd6tMhSqwqYApkO/jKuKDwEhZxWCzRDVxX77MdxweU4
YQaaqNU0+9a0D6RQJ1+BT+RszPiml2pswI4tGmoPC0h88rN9YKvJHsCv5jWN
1t8000Aq4xkSKiQFK1r84nKkCR5jLtfXjzEc+iPOLl+WY93MUGdqnLNWkllF
1EbAA/6dKkwf6LoMMycna4IJ6P+h4bTLFGVhY8md/1KfiOlBU98fPON2tccL
4BpD9c6Pf+NoldXPzJqBOMZJRvKDSxQKQ/Rcbr82K/7+e+pnYCWnGOj93xBZ
9+6NxeXLu73Lh973LvWCpDXFWCzlXllwsaT2tGhy/kS/lNc77mQNJWLlqjY7
CS6kwWx4l62xuRTAMrDRNN2HPanzZTv4fJvs5aI/oYpsMezaSmFNzm19zZDv
/EiXoaz9qKzb1dLJlTD1xuMiaeKpFhiXTLDSiqxR55u+xc0940UtjKIzB0dz
t0FDxAPuF7EkwjCJ++WygtqerHqd8Vrw7nWbpRkMU/NUuvZlFCDsL6Xr2Or6
wlYMhfljy7Zym0PHlcEVe52W4lj8dTtOYwox/SF1GnF6vDLXMTqmqiLKovkl
bIF+kEEKdCDnTfmDMUBrYPmmVTyrfLvuqTzxskTSFrveqrpoXugikAQ5+soA
iheQOln/8VzCiYGKutXzEM0g22hCPD7/RWqS0iZL8T16FC4sIkPRmOdw+TJ5
PtdXc6OCh2sCSSjcyeNSSumfrsyCv4qdKhT0a8cHH1MS9Kw3c9+M0GBUeX7Z
FTaUdiPnbiFej7ZinLzrH3W1yWAjvrbaB1jIaPYVv+1OFeRFFKi5GWchY7CW
5tY3nZvZejBR4rBPS0uouvqeyktmc6w2rdWwkibrjH1+GMfnoe+ZMEx80XGz
ldhT8rwuWqecH8ckHiyq3ab9CdxqD9f5dB/U9hIykYRUYp9/Pve1BK0srcXH
9XvWJN50v3KJuQ5hBhx+jXRiRMqGZ3595h9gfDPouJp6iS6LxPAO3LsbJ60L
dv3TgkjkvwC7r5kRLqgZTbpPYZ2qAnvDXSkfmMng2fQmC9RoWTFgxIStAmBA
wZu/m8ilLg+sMBluBuhgY0u8+91YQLxfbPsipcG0a3J8hp8EFshwGUpZ5ilG
N1h+3HU+qt0OzJPdgOnCAhx5ueKezenISNfcuxhuaLUOxZVzs0/3GtsGEUk3
MD4AAT9ggq8SrlKLijlsu0fpyoYW4uw26euVf4fF6/fNTqJJEWTbOquV6vXe
MMr6kLUxCs3VEcoLRZCSMmkaHgJmB2WHJ7ZLL2KDlJaDXNlscszYvoDd+tQq
0oDr/ayRjZCJ9gRLTUyGtGY8re0za9eYahnOQfibE0NHvvgs4ylPYAz+ExJ7
Z2DqBirrVDQKHeoIU61kiPldbDd6m0v+ShI7xz9Kyxc3WBkzclaavesNGHPt
c5dgdI5+w263Mz8u+uQr4nhowt6f/Vw5b9BWDwPA20UuR1NFAe5OdHsUZmJ5
QQ9EPfk2MxfpCws9GH+fSNa14W6FA9iyHOcLwC8t8GYCEFU0CAJKbQAQzGdy
qvPyOjULUDIDCiOrhHg1sMRYUqDwhd22uTtKoNLQS+hkEqXeKkJVLQHz1EqC
e+EH9womZpwkRUyL+MYKSSvuZ52TnN3Qkw4ZZn//R5I7M1Juf7XrPVzNth5m
NT7AKPKsnOKYB2+ER2VbpTB/jeLQB2q6WVFOhVGIiWGcFqYSEewXC3gWEB13
mu7P6KSLnyIz/MDGWd0GfmmJMcOf/YKcYzsIiHA6cFvraoQKBZyOcnofq2zI
6F+AccfUe/m+7UiJDaSrz2DWByFkQXk0xsAcR9a+L4/344Fay6J6KWKTaoUc
BYpNirQI0W/Wx+X8/NY+TT4R3ycQphLqbEownx65GAynlWfHDedH5kCmQlRR
fT6RJsO736kbrn8sSgfb+OKCQ20yacurjM0skbRdnn40mOrS/QuUK3zFSoCh
KTvtZHpbmOSM5FutVM38hm/0YVOJepMX0/RVpEbq0v7bAmgSwMpB9tlNqF3v
GjEQLg0XdPTWxchLzoeFvSzIO0B1SaAzGQqI5DaVJqNRwRLsREsgP6dz0Qq/
l3iGN/VwLgW9reAfgKzLXQgzfbEKSiSl3hYTgEfmFi7h1oR3q/QaaXnTzH01
gRGR4lhqq8StiHaoy7JtHUu7CNtP0NbbMABpP1iz8U+A9NgF+4aPY+jp+oRu
jhP0aS1aW0rkLVTe5NGvvU5H0Tt1X1h19kJ5/FvJrj9VykoMmsdPPN5p748/
HSAEKB1ms4o7kCWMEuXpKLvtYEUieZH2zupGKcU5gfFupNOhIkO1inxTosxT
dVgJtkd2caBeRp6GX1t9Fjh5edSuVVESiUOKcz/JLQlJ6QeCz77j9GIZkrj4
1YY/bUU1OYJ1mPq9DQ1Xmr5QR4Og0EIrKjwjQP0klJ7Ex0oGJb2+SH8IlNhW
BzORtRJlRyb/FFHbHb7jiRQIaxDkfMNcm6bu0RLcG5hq7320l33kWA1eidUs
NJ0Om9q4VlT2LAYVjFsUOzzV2nFG4vtKSj7PUat0V5+XYcft4HAl7HbkAzUQ
B6G64HwaFk4Bt/3xhq+zpTKr9qID0wW1CmpnH37KPE5wlizIbflXoHkQBUli
kPtJZaBdrJC1xUShbLZob6LRfhW28Cl3/1TXYR9I0wMEMVIpxYogUNeaQmaI
sTVUsQvmwwzFC0W+jCiViH5xJd+D63FZrSp3t0CIJZG4MEMqC18JbkZ5lieQ
zcfgpQYO/jrmUZN5YvUVqEAfIAq2UaL0JxgJUYpaRiFWWxjRO+5Z9WGRRXqq
TUtoGS/j4hRmT+FRxOGS28NAFmxFPJ9tzboFpSQP3IH6o11ZPt9tzZBhNQSk
77KDsVCjh2imjmy8pyCitr/8vKehcJs2dANNy2C3oKpTBhiWWeIHQ/eDdryx
K6pVheBV8661TPBBzAp1/z+VNX+rewn8cXrCfJfTOEXiu0GMf9xyjU7qxchW
8i6UTxrz/SEOjuMW1AFjyk6JrY/1p6B/iJVkHLeVNL/qliYBE8wh/yvvgAyT
8A3hP7Sr6R2qPf6EI9xT+UjEvOYJxGsJlZlWp4NsVhQO8VUSjt6ogSuxzG3M
+SE5+Be+KYRYgTMn4EEFSb0a8Eg1fiqKYExt/jdcOqAenB14UsP2LkvbNIoe
qLcJGP4NdXbo4+HB9lOkkN0m6Ez8h56KbR6WXVpPY3HN1SwIubVZk/MEjlmv
7sAAekZZPlX9XIUg6/0W3QsGlf5BPyv8kMLh3zj/NAGe+CAOwf/i9pgImvfu
kSgw5exF0DEZyQgaOdOdVLPIfi0jWVXApFAB0gmzuCNXQ6tLvxVJGkeBbp7/
EmDHdFnXaQIQk1Xj7Rt2qxwjlbyHEPFKcE2HWI0Q5+hWDCSB3WttVOUHwWFp
1n9pueQBX+kzYJ7hOBC8MKySNeO1tv62uwSn6ud5m67obRrwIuJ08s8ddzsY
z8kLtnCwK7sQYy89ujmOOl6mY0ZmqUNsX3FJInKw1L6pey1l6PXGqkf7Pul0
ffzIVVaydGbM+xqA0PzNC+RRw5GRPTXweKw2VM2YW9jFTWJVZNwyESc2TfxN
gX6p1cT2SuXncw2+xgFY+znapax5hA++th+V5E58f2BOpIrpabg8LtmFCSIs
XdcnpTOslqC+8ETGsQOppUYaCSKhbwruvX1c/JGVY7xGG7RsHSDP06pG1BAp
0DB+e5K8olh33EtdaCd5X6Zfuvm0F/n8XOqOy5MltP9Wo5p90rQUffqMO7Rn
rScHrdvJdnkDdYdhxZYUncMMVyIWlxm97OhHRK7m8iVKnHgmhk2bOSKN+bzq
JNYt1hPHQobK6NDoh3NLekg5anqvUTT8mskltQ6WJv4E4PmS1b6ofuP8Chdo
stCVgXX/5lQ7JxsxbibrH6VGBqLQoy+IScASKAaBY6ss1N3XHfDdTuu8xZIn
IIpT2XP2aNjgDp+PJN9W2PW17XzaX1GswtYhJCcCSc8C1bkj2BLfyCmIe1NZ
rO+BuhQybMsPxl8JhbmWM5j27bdCXtPhiHKIji4+q355CEnH67ZKnd4iaf1u
oSKj8Z0GftNvxwd1mXuSX6thgHDFC4kdveO/QxCSDR7mETFyo5etF0x17g9Z
AvhUw5FacH1YvemycAtpbFpazc/qxgwEHKPt6loNyhu7cH9hUJpTO2mjC7BI
Ls8m/iqLhUu16sNORV5lSQPdd+H7GsH0uu2n+XiHy/T9yyS5fZepGWj59CjW
K7dqeevu0bU4nVrrz3UIYV/89xpIffB5myY5GqrpNqfivkfJfCOi6Iqkv/Sp
CXCmQbV2RExvnKFLf9pgQ8c81/XP00/2/MhtVFscO6eIeulIE440txDcYKyb
XhaTWnbjpcyE7GzaMKF85fy1ixd0D97MHkJB6hjisB/t9zVci0RuIIIXseO8
UMIhsCCeKHpBfvLDlCoTIzeHz6akvj8e1n88Fw/Li+DR1IvHVL1lTEQS2Zri
Hja/ixuAA1rEldZSwEcGPtVkbtRmag/xMAFM9HffefcP5JU+Sld3kN1TPDHW
UXRkT8nbdL1Ti3b0JvipAmVo8XaxLGXglgcgtkb0aWgjiZl9GCBH8hJHMY9D
tLZAQwfF5fhyUpstBT/jQDpRNwb9uV7vbzEQOLgzIdoP+a13ryt1ujT7+FnY
akhQgbD8FRs543XuFlraD1DJoHrh9Fx4rWO+9xSXct0O37n4B1wNHOVAj5tn
RIiAZ1sRyvDgDm/QHdeDGl+lcmt38IXTdOV/bxqScdlGmQC1ce+4pizz9iAY
/3v+iQ5h/WG1Z9UOCAi4ThqKo3/h4V9+8Qcsz9bxcwf9K/zXT8MkTX4IkEWc
ehrUqZ76l9u8n/se7fWQ5aFPM7gTEnuY5b2pPlbVPexJD7l/lThvGeUW7TRN
1rSs8cR/Ax9FsyOKAs5zxjZhMirnHaaVtEn3phGIhZx4XtzPrj1OWGhJpzpD
6KwvjNQcoSO7Z4gdeoXriSJTPtfiyRJwqv1Pg2oLWY5iegX6It9JLLevNuhf
ET8LFWIU6lnDJ0yvoBJM0vStIQhJcI2ixj4Hp4/MbQ/pRCTQEcNjDrAf4tEb
4+jV6g3uS802/7mUKYGJOKFO0BaafqWaB97weHw/alf15sKJwYxwL+oKIX4v
wzDxGaeKSIKFqPTkLzuSgsLSg6yur+j3V1RIvqnkh/jkNgLFIk4MQARFJjW5
b252msatGRFZIeQYgN0fHJhftjGXW0wO2nVwT9AdD9fyMRbeA16MUOWsHg2h
HVTSMVG2/7Tyc9f6mgYRm4OdCdxFIdoOd+gTkRA+P0FX+YKthPE5dv9RvNRK
xxb/4qWqMr35qwHSR3xmqUnxWlH0h8JQUQkkUmCL7Lh+qCLt4C9cuuYifWyf
GElFuN5fEBbHfLnIl6/vJpf2EPs2CDBT81Pp6Jm2XtK2F9VY4/RWq0Rpp2/B
3irlPge+jS6phZUC6RYfx7zoYLHVaKF090RI357o9izd14Euhpy01I9dojli
bjXMCbGP28upyWYiAtbedPAGLvxw5Xk0KF8p5T2yx1T40tOEeU5j5ZoFo6bE
a0IQZkESmuCEeV9QXlNWjEeVTmFwrUKg1OcDi3DQEkGx/i011fFUT1atyRlZ
sm2zTgz7Mf03NVGE3wq+C0GsYKvD7Y3qSeubPp1+i5r+NzDXR4hC9Eq8CGk4
ARbx3cKeh84T8cASwk/obAvm1SMjoZkOq9zPMTWW+I+6R+nxwdT9iwljMEMP
Tjq2FGQ1GqzvQy92TNdGXVQRzfaHuiE9rKWe6LLQorkYqNuoM7ypZtLTT8PN
1YiX26WRrTNxG/KYRNYpYwLMhc4rgzl1WIyt1bwMYzNXqG6AHHlW3S8YCyWm
AOFSchuGfTuqeFURQT79QE0P/+cKyFh1Mqfvi8hTntK8V2HF4M5VJPNQnA5l
a6SxZbY+A9t2ak6Wr3DaB5lX+RiaYIUvnWkFN2jq6qNBOO+fyzO4UMSMhGu2
Fs3c0qxhn/CEFZOtHN92x9IjOLmwX6oHy5ac/6XcIbwqscRquIAh0IR43fmp
BjRohU5c8wj1Z/Wmpx7CXTNoiG5hlFZGnDNJsPvZnwWEiC4bvTHafcaNpg0d
1ynDpunKLVUO9MdFgMtdAER6b3jC/e0BGlbjpbAk3i6XVKP/EtS93VE1T896
U6MtE9Avf2WF0TQ9sVLndd1Qo5PB9hasEJTj5V4Y6GxdWaHe42Ukcmh5homI
dj0cNlIb81PZ9TM5Oibqvwq3XiYBAxBqn/oED7M6mNuIQRo7WZNoL4gicg/8
C7+ITbzIDBf3rAxD3xnmZNLX512DArFaPGimu5pHlguyqsMmcYtWgNR7rqaF
+CZWnGYG8SZw1EUU7P3Ukv9gb+ve2nGqgd4Ko4nGNmRLGiXtNNdGkcLnEw9W
doxeYyZAnur2/ESUqPVqiKbOD3To4aEL7jX2S1Ke/tTzDphdp7DRWJqX0UCK
WR9bhW0Q4TtX5BckEKQGa72vYmnrVPcgZ8E4/arLrXjuh/uMPlvSGwPjKAM8
z2LerPHuDjZrD595d/kUhZJxE2lrgcWbsXQk0rI9sR12L3Da5y8E7bLlcvi0
3R7TdtzOFq4z3JmwVIlZoR6vsPIyMmGetXKvrOzCCqOv19F1C8Df4WDx8+gN
uKxduMRdcFkzFESwbnTZlZYY1JvRfn8PZBnZXMTCkqHvLjFnjhpIT5ZEuP3B
Ibvj69paThxh9GlHd3DtyKbYPd+TkfBaKTK+xrbjd730uZhz+xPvsZsK5g+n
iKtlq6MPGBztUe3Dks93+Y6o5JvTqBmq2+KLOeT8lfOtvnBXXhVe60PPYkLW
wgPgnm5fJ1Q0eBQBfsuNgHwnB5J+x3F7ioNpZBrjW4GkMxAA3utAh0OwEjgm
93y0pVCZSQiGqLK7orqimh8BbgUMRDHEudoY5uNYaQg3zVdi+FKNHZWVLyqj
PrY5EfdcPCGtRWS6lV6n0sc+JlXaBha2EtCnAQVZnyH7vUwrdX15lmdXlGUj
V/5gQxnHsy/viEw4NqZNXOKidHlAxYLyREEGRLgJEZTswQgaoZWMyfHNr0DQ
vLZyimgLLdkxknE57/E595ClnE499yBhhaVJuVRLjhg3uBr2FI48RZ/EGWGC
ujOugXLo4wZjXqZTtyCMpDa+zh0zj6zhQjUmzqNW4sU99rMvBY80Si/7bsR4
2Sm6YcdkPU6OKf1ElTk5Ao+xcNkgkAbzDUvadgpTbrnvHgec/nKkZVhr3rWf
bmTq548+/u3cWcHQmNM8T4i734LZSHTZI3yJmpDMLgUm9yMU7OIUfOy+vc8y
ijBBv0HeTIpo00xkvqcNAu4cL5Ce1lrEw8s1fXThTsG79swXd3mWM4K01xXJ
ZWq9zEwR7y0qd9DKysalGlQkWP77a3+MFJJ8u37pzine8xnzlT4en3Ab5r+p
ZKrhWrfRnfuw5bWWt4UqH6GK5YSJMVEBsNbwIV78xX1wVM74fCdW0Bko+NMS
gO8Lrl9tQ8Ah7Zkw+Pugpw+BsukJXNNQmi6LzhFiqLKM16sdUJ9auo8Go6r9
WfMzmd9zU/szzJ5dJI2twK/2xcfqi5iobPELHZ/92T3VG9jr+0kuQCvUF4Dd
Z5mS5wJiHpZHbzd3YiBdtiPKxQhJVP7OWSWiRM9t220RC6yixEUwc0JkEsHF
btaGrK1C+pmbm3SmGhoBE5mhk/DKHHwrFPIT9mrZrCougiN8CCYllem9u4oL
fu7AQTn41Z/CvuXpde2H4MEb8BGztuCntUxtI2VtY3lhEOJRdJs1rhP3TDAq
95j6BhNFltrjxRadxEWjZvF+JVspQ7WPOxFhac/Mu848lz/hS6HM0MUfO8SM
iKkJQDKmnYZu2jh1fuRkYPOLzYWahnKbso8INfEBKcUNPb2RQLY8zxBl/AeX
Jo9iNMOl0M0UK73exT56p8h7aYazxphVWDihsjJLS4iE90p/uSssfaILTSt4
ITElg6M+YqbO1R0K8n5Q2X+RT1U5IXJtPF08FizS4myE+hR6K+9mVMEz112c
107aZpBDfPXpxZTZzK59pk8dbMenGoQM5C+VpLwXtkD2EEMq9sO9M0j7Fr5Y
RipDHfIuJPHQuGX1lRQ4nibMkFMinfCZBGupPxhfXgmUQokQkycdjkvmKVbv
e0fp/A3kphcOs/fvRTkAmNaL8u+CEJkMlr8HnV9kwoLt2+PUNXmb9f4EnT3O
v1SJAEpndQLyxP+HaWZ9z8fhP78t9o9x2zOfy4WKOEXV4+EJlS/TchPxyand
3Zf58X8lF7XeKGkyaM4OFZIPDy7pTqOQ8EmHtVG97hrtpKf9B/RPaG5ZIxXX
8+qna2u3SqidolyLDrBQo708vBd9sUaUusvUxQAiMRwtaGk/y7DTc9bJEFUl
5Jv8ETl5TpajRtFQhlAAeNgW98xW5BISzcC5oMZ/EinsR5MxB9KVyFTxggBo
vlKPfaLd2r6JkihJHodFpBz9dTYmXNMEM11lih7IB7BmdT3uBArgVNMzWnfX
5WUIg0LFlxsD0sibRnmplk64+b784OSL/nvRuR5bx6idBdkIeMJ2v0GY87m7
Z3DWabdHdq8ywrsAjBiJva2DPpHvyMyrhDXATcaLxqS4ClgF73e1gyK8pi35
Nsj9c5/XO0oWv9aamiwSxZueTmYPA3uEiQ1l1ryilTH++3RViEeRwkNXgyhf
oSnFOl19efHohExc7ZL4iufElFy7mZW1B76W7QmNLzymTAyf9hy/vjSjJwBQ
q5FURA0r+Rlv5kLWOeHx2MThDIsKRjI5AC1Fp0UJzlaUDNrI9MYLbUofGMhx
IzHzBGKfbRRqV2Ww7pXa5BpVHHtDajLtY5jHNQ/HO8X9AKVouVvvvtmRazOw
cDBNNVhc/v0hmcePMec+LE3InV0O7XiDd3E3JfnWzHlFdUBfjqgRcTzH23QW
3KSld3OJDnsx0APN+dGJdfmGhxY06nj/cRGhKKBV+8+97SWAi/nwY+KmzDMN
mqYq35hXMPF7QLGbgblCTTCcFUQXXu9kIRbUody09+Xz6T4WoTs9IRASc9+J
SkbeVEeBo5dj3f1Q0JAwubQlBwftpAgVqoepArhtQGuE/i6NCpimdBBgUaBe
Aig8mpaOw4ukfbQ1rf1jM98WHlFPEie6J2dmbd+UIkkNjBWcuJCvzVecoBZ+
gMDmPAXZoBM1NzBe2Nr95uZqG2MGx7u4jooXR0vD4WE7SvDiybeE7uU3npRQ
aFGCA83oDvzRV+nNHWgnI8IsbqcKaxl23K0/9mX8f/ZnkSdDBL5q5Sp/Mpqb
yoMtHafu2hkrtz3BVhCMxAxmn8sFwJi8NTn85ppKV0U2fWvXzidZyIkJPKtv
mV3pMr+1m3bzN0MQEcF+V+ByFzxJZNfcVyPdD057bCc3d+rVCQPAkk3pebNp
n2KU1/6F7dgwq7QBb+Pl4DxbHgXQZwA87GO3VDFPpWVJiAY1vfu05RTcBNw/
UM4Fm4GBGnfbgM4al1vzFjyAZLdabpbpc6t0cFbE0FyU/MfsfF/CMm9PTkOO
JXHFCGNFpyyoY9H7g/VxV4jT4wAPdQ6aAQvK8Ud0Omf410t3tvDXP/GNrnt4
YX2YWwQPuxv9jzqxZp2/B28QXFaNM5bztXM2ya5/DzGPayTVqrqo9lm2uHoo
Sohu0Qeazw7iQ2msFt05xj9o2XwGogGI2ZLLhBrOWlyiqU45aiYyXO9H9vH4
p0eFrMXSgDgM9ZC9zPbUr3Rf3ofLp6SoogdEdJdD+7eLvYPOd3wnKs1wS3Ou
jyn0pqp0gSNfiIe4AEGM1N0wEx4a1fHUgJNOsDh+2O+/DDtMZ+HC/WwWFe5h
nHFcslDGeTkF+6y0q3s224QRIDLx1HC4xeH8dst+EcoD+oJl74E2LVnkLHEE
3fHHB+g5rRiRnzcGy8uLJK7r7dlpV2JoD6bQXzmlLhbS+vTN3SiNrIBCjwrY
2HcvXDFHbWoMShpQuiHtOWcBWlYi/0IY7EHdrPko1FvPgMn1k65cfqJBck2T
qR8YWhvd5QGMu5StXAiHO4p2GU83/BNYHKDT+AsyM55VYJ1l8UwzUspiHu3S
fDWiP0SelQXlHpFYwro50XgwxfLpAZocdxk/uRaSqqJ41mAPFsJSwxRUUDVY
Mk3qLGfAQv2XPTSJP1Zow4GOLTgg7+TT/koI5zN637RnR8Zwxg43s8BoYPnu
iodUb30/888XyzLOkDYh+2exKJjY34erGkSQy8vIxNMu0/dzOwUMkAByTNUt
0EDhKJLb1PgmugizksO/Szszp7Ab9CKxYAGCDfg5QWbgfuS2via9lmg5i0qk
DZC5rdQzjqi7R+BZY8O/qHbBcQP1wZ/in2fSpVUYizdRQNGPmUBGEKrKyosQ
yPsE49Ern8EaMl4vbBJRjuTPnxH2E6YDe3mayCQoi74fzElTqtmamymhcCX+
vvsix3+tH6P2V8opWgEzN9fIyuhgTKZBMCM1VKKp97mpq73udsrVzfA5FAPt
o9L/bjfcQpMFJWLvzyEh+F4XWQAYlWqbUQGiIuEfP+/UnWzVxMX+lFyRd8lc
wqa/A4w+eBWr7iJBb/GBVjTGPx4OyP7BeQqJ48Asa3+1MSRutQNlQtbTAwSH
vAq0w2QhV40yuygPgp2pkywILOl3WLs2rY7OKTr+Y7xPBCYLpKgyZ8Y/XvwU
3IXPSODSk1zf+5MzI81UcKNhoJPdClG4gCOv//JA6oDplSez7tBdl1/feGVj
ZY3HcXj6kGsPnADxYCBVJZnqvJY2D6t3XKgaMHRUX4nW5IfELJR3cTfbH9gr
Z3kRxRPNsR1TZg7F7bqhx2Cm099GwD0TmhkTo9TDqW+t5yca5yUCLgq6juHS
F0iUI8sEo3RB+iyI4vqyk1dSKH/6VBl1/hgQip0z4+aw6maySzQi/TQ18Ljw
YVWqlTdiKj/wcNNjHU9LytuV6RURJ6bWf/V4nGGzSmj4pBlqDvAlkUiyfOj9
xAW0eiNakXSSZVzzivYr/DdRHx7os5FPDdzXteRY1D1+yl/WDTKB8sZNCFmV
U+ZOCEBDXKAR/4+INj4hJ26DlowhOrVvwXZvcjcRyuxyS5o0CsXFD2pI0r/9
67NQwJN98XvUxLy9rEzteqmuzhgk5NK0YICFQnNwuCoAWBwigZPfmxnFJOgh
S+s//wBtgkulbG3mdtZyTpDDXnqigvVGuj/sPbLt28kRMLqa+Fit808Zs3+f
dk6G9QM1XtFO5sX+9bYn//5Bl5cH5EUSg+Dv3sgdf3TCZ8o6SImmmvLMat4G
SF2/R5oxxHGIEZ4EuAn/YPdi8ST1zI61n1t2GacpsbAKk5kEWjvsDG5MrN8R
HU06YW5yv0Pwnrz1d1NlzJy5vF7GizpDJVQCcKasUkIRGfgTq5a0mjsDhPqB
7EHJPahSxgclZtAlxm7xZrwQ2joGtO+X4FY7EYBd2+R5TCZjbhcfbMvKyon6
8/7qAIUCpJebM3n9gyGkjqBXxd/PnthAIFALkGMJaCbEjtXMZqtovBzZDCzT
5mxjcYBCSkoxRDdrP5OwLCJWabIKQpFMnn+NLrqgHxTVs1/nVz48BTPKy6dz
I7gKOfZ111eRysgGABrs6t2wRYHpkSEx1In1VDlZEOOjHhyQUxbDCDtWQ5aG
oz0o6yBZv/IYhhih0CHqPFpWCTmFIWT6AVPo0WbspDQZb+QTnzmVbF54135j
YvGAK7J8zuPdvKNnOA82YOXoWu8wXAwLHpqeJhOvoB+oT3hEuG8XKXdB/OUS
4IQzyyrOXcuMgok+ySbRRw7pdkjHPktQzDvOtzNmAc3VcNudte/d+IgUwQ/2
enxje8061sI0vOz49bbElT4C6xvF5JZ+F/kqXQMvRqSFEG7f5Urgwrf80Fad
uEDreTxDStPteG31Hlc0UFMBxtWnUGfalxEM4oH5ohLYMzTymN4Ch1Efeisc
/vZRQnfzylhAvCni3G1gwa9sILWItQygUktJPtNAat3ZRZDHWMgKyjAfXl8d
dCmFBlQIZuPBr+onCm0aqrUCd94c7VE6tX69QWyLLoQ5PKkhsaO2DEbsuJLi
lORUDbeiYS3rsA5kaooS7yci2N6w0+iJzgNcoY8yQQR0CJd1erDHFpp6j/+9
oYfyNj61ZWwm8TyoDzjjjPF1Aj9nUgl7f4Cqrctl9UTogd/Ow4bZpOGgXQCQ
Xr6Iv7r3rQyKCuePBicTI2aoO+gYMAomcptggp3HgV8hX9Q8Pa9JgNYHslfX
Q98Q/7S/Ude/H6C4W9uBavfS1Tf7HPgmO5Wl9BUp3DuR1IvkF0YSXHPrw0Qg
w2+xQt5U4MPkv6UAOh6fAiK1BbV6SRpnAwE+6//FQ52/xbH1ixwpJa9fr2nk
yMaDDj4Uhd+jk3gkuusaVnsn8f7bkdMgMylICoLYYxM7hWTRlMhtj9dnNJk2
jD/2FnDdp0+YYT0qrI8nPHBnBr+BudQTFVfL7Z1VMlKHmKUR0ZswoOvmcQzt
PS2C3QUvQt21lJ5I1h9zQvdISQcOVwIAcZKNPX7qJXl3uy7QDcm3H4pfnUEG
aBFjHZXlx05BEP5ekn8NwD7U9KVZAjSRwHcmdCFshNLcuf7LOQi+miyuY1UT
veTEsnbp/LwBaFi05pdpg+A9s+Xkww8gxXqqJNfFMQ4vqH517K+04KonAnxH
5glO3wNnjQ7MyUbZxQEzE7shpaa3PZ2RPYxFpfFrI1y5cVs2QWp8lcPRfCnT
AQP9ACRsdQFGK46VDbRY1GUgBiWCNIb39f7I9wLHF/qUDt5A4Qgyb0aiK46z
6JfEVcXBjY+JLoOJcVkbwJScKxD1mi5hAEwNN4QLbHq0KhAwKv32dbkZmGwp
7f93PxFKOn9nHT56+MM97eutwdmarZ/1w8OAZGWwRrs+vEMu+/6dz90A4deD
wlXFRdAr0MJy86xsIDHcIPcgCnxXz740yceB40RV506hmWK6QnoMn3AnCoF1
c+17juX5DRbswpRvdFJJuxgrA8URYHy23Xgu55Ky60Uf7AHtYExuuzVttXqO
uiaYELRY9cEOtb0zH1npipE4joNUlMlCm6KiGuNOxnZvO8k0N8+hu8/h6jU/
Nwn7WK90JqtYD/LT+6kWHBYP5UV9fDzRNymtRBl1hLuRnNwCQIN5UWvzrCe3
Y0/v62FhaKO2Bo+BeEVTI68E1uGB4HrclmI7nnGN6LjuZDoprsUG1Dp6lhmk
nXb48aK2mKojUOCUd3EJhKA6xfS15CyIFK3/rCgckfVqHmQhCjISB5g0C+7S
Wl0CvuU0g4aOVnS05vp7gvUzHVqgDFeTQXM68dXXYv71keYGpajCR7L0Wvgl
2MZV5Jd/BRBDm0O4zQwkwHmLnzrFtFVZrPxpAkYxtV1ZHvubfnKu0UHjYzTb
VOqM7Q4A8pAuO1uvMwXYa8URSprI5Wz5VcAx4H9YQ3LY6MFLkGk6Ym4yOLnn
YIJSScve3E9zSlYCGDuCXnmIye7QBUWPDqDMzcc2lC8O9eHYkSDbKuCHXMys
1Od421tM7z2f40CFjfcbzyzh/r+YUFnGzxVRmtA7l3iET6OX5VIUvDBIu5nZ
gCjzzuowvUKmmHSHtTt1AtmolhmjgHO46QXz66RVDdUrKsPbeMH58SFpCkvW
BMN7PkUoSjvDP+fOAMWisbnE/9l6/IwkJd+l4QaK6VelEd2TTDIeFWMJMzsp
2JJ/5L9g2Ukos2FydwPv8xRZSw5EI6/am5FwZ0MUvFo6hw2XMlOEfnc4llnV
NTym39ZV3slLJA6q0hmoCf3cg7xZubB7RgnvbB12cjJr5Bbuv4Z0TfTtZmvc
Do3MRKiAXFS57sici5GCg8FCAvI/NLb9iM5xzl8lOs0pDbjyCNna6VEnSHvZ
xs/kEB/wX2XWKMMnX3H+EPmuElj3z87Wt1b1gGCRamceFSGlLGCV6XEywglt
NyU0ir9gDElozRwVhx9tp6+HMrTpcQuDyFUochkcLpADB5PyyoPK6mEc3wuC
JyIdcsrE0zWkut6HSgvFJ9R/MZk5T7x+uX9aM8qB0kLij85teKW3OQPuZqYe
xQ71zjXHS4+4cexIVELY9Vf4lbVTiIsGLtBwjzXoJUqhSd5DZHfxVCbJdK9M
17NsaKOV4RXbaxZfAqeMX39OCfwzek3h3j+ITwb02yQYaSgwUdZll2FLUT3H
dW6SXTAggmk6TDgDx7GyuVEqIuHRnndnYjgmHxiov9uKyLrEO+t2c0jRhdZ8
RFm57FRC9Kq/FN7kEc40ZA+DbAyfqocbX7tyMVx62CyK1cPZrjNQhXCAZ6Ml
Wh6k9KB5C20zQTEHIEqkH9vjN3FCBN7wOZ0z9TynEDSqT2Zq9kLrCNxUvbSJ
3NTh1SQubbLwS48spxqB5ZZqHbJB3O/OKidjiUblvgXiPa4zec5pJ8kzL1nw
Cgks0HScMkXw77Tj2CrI+mit8xoDlpU6WwiQpK1v1AGW2+inqEqO7+RgOrVv
bWNY8G+8pV4jamuS0GTzQKh+Txf7K+6vzXCVswpKk2vh49Qfe99z3BMr8CYl
KcJrb4/FS/EogZNK3Z8kQ7yGKosXj8SQX4NM1cZcJX2MnLr24ZTG2Lb/4Luo
dJpwmUSbpaTCv2JNHMAsDVEdMFprwixc0ZcdPnC3WTPTCDVasHy+TniADPuN
AtYEZ6SbFgHyLKv33uNUpWXSbITTenhDcdmL0dWmcLjKu60QlRMP+5rm1a2Z
EKnENDp0B3+RV79dnDQXxZZeXsudBAc+XtKL3lFensIh9a/diLK6qhLOZ6oC
JCKwPIolDcIBMm0GIP6fx+mp+ih8AubluYjWOAEottDfzdKby0CQ9LJgcy/S
iNBca97Uav8l5xoyzFqRqz0KWtm7l4ICDywd4hcZNGJ5dSVIRJxYmIFukmdy
SQLbjvb4FipiiYHuo0SrYWYUlDC0c6LX27UH40i5EQ3sjnefdh6a9h5E03XP
GSTlP+f4UORcqykNRvZfYLmkJa/2CBW2qJ56Nb6YkNZKyMAJ8jtPFfOl9FMc
daq+/FV5fGesBxyPsa8q/rpVWJziicGLJ4aneWCxPsGI2/hFdqEpdA1yLwHs
rDJnZC+M5ec8Gb1GhLnRRCSV8WwiRbBZ4LdxieotXMOaWQsZl5GDD3I0vIRe
Rrhd5F4fBYpUZTWFZlvwS6lR5JNDcZOCZ4wTuceFHeQjEcNlQ41Aig5ha4D8
RmjS1q5cM4pxihd4usqO4iZFdGJ0T1cMahE3kLqxfQYxC/ZLM4vdTkzHFMH7
/COyTaT7Dp/x6ZB+qMVKTNUiTrSrtbZYXSeB0C2pIP4YuNWfXBNy3+48SuPQ
wXPVTlJ/SzgIy+y5VXDL+XMZpgv2Ubmvp15KQldlFVgN+3XibUOoyElhOmTO
S7wF/8k66rQdjqxnQK+r7/GMsC8xyJkgsvDJ1kdXZbhByXE17cn38XifssVR
8J4wH/qOAUwQB5q3XDUmcpBXQAlCD/KV7EWzmQaE7NO0DYL5Ttia6VKAU3+u
y1iL0HQUwYjb71gXW9xu9vQX2DD1IOwNumGtWcx0uSjeNMR4MsFAz9mcwzyQ
9Hgf3lqARiyXjz2896YgYHvOyf8YlZaCh1EruPwcZ0B4Y0pfcKDyZEYKTB/S
kfgzWFBkO05oQi8ar5lDhsHuR7YoaF8oFqBIGlJ69ohj8fRvVrSP4RFD/P7L
dtfl4raYbOli2+LCgD/oiAtX3Ha0iN3OBwFv0Tc7RBFpuLlIG5jqJ4hm2HtK
BmESB6r05qz/RUdgmmdOkDmQD5mPnm/4Cn1KV00BUPKhdx28nVb96fz3w5xp
IhwnU4H1hM36LpB9YR8rWhGhJVTJHh8sUbZP2BDP++kEEBGSRL3qYI2qXieM
YTXOXBXfaaSElTSGHKytqVnuzfNj+IWfqfw9sp2CQ3O9SnLoQs+cpr6huDBW
IY9Mr9BcnWEATk0qB+ufIhaJoD4JY2eIlfwbgBpKQcSKseKtT4B9nKZibcmD
25ZTrhcdpyYy40fDe0hG4OBWntU3t357qZ3AMC1ufMkzAo1BEK+dZ1x+8nAJ
9M4+6tnH+gwwiRx9YijVhnXA9YN9MMB9dHie5RLGuwRwGvHuVbh2UIlB/UbH
uZprEwt8DSQSI+lo/+ln7jF7/NKzMwh1PCGLKLLgL9tg/ha3TFB7rUgNjVjA
pg52jF38jvwQLB/0yaMvpUxdCyUJmFA5m5oUdBxngQsphxIJ9nCcNmrFKF03
hONta8uFZ488LskJaz6SfhSZlyLRCk7RAdzeqPb+g4o4ItO/vwg/MIo7s4Io
jCRVo2kMjuARVSRldGFbs8OnFrz5+d27994ntSUd4I34xbXXOzY2Zob5od73
XjQe8ofVQVY30/lL/rD0yG/m8zXVlsoAgRn1gNSQe5rQFHIk0kPSmA3Gc7eB
HuCraQ5fX+ho5bseo2BeJ30xYHq90rrvOsUqJPnvG1ZL22CSrAcuZDMhNUFS
/n78twl+ZHQeoRw+fb28QJfZtnzSUbFsGK08jO3Cvvt+eHYGvLKwwRANBbXX
qja3qQrxt2Ca8dn7/sXI/56wD2la3kzlQRGFSNUbKNRZGcepa4rJEBgwH+3J
NqCLtSH6m6Gm+W1VkNrY7sYdU9Hk9zGvl5KClQx0mU2iPBEraAaH8I/xU1TA
EvDGyEXHYVj62smUOdhQ4F6Gadq5EBapOqV7laHrS05/TAp0QP1iGV1JDYKY
Tcnyv95bUuvYlMJ/yhvhr6WsrEhO2U20CCS3GH5wYPA0t3Atzpq+qAXw7HQV
6R6vZ987jbmXlQU0f8rfw0gDg1JKp9FjlXpXEd6qhKA0TR1iNHgsUxvPo0Iq
XEhDGvAb47FGLc2lzWQOYToaPnngU5VYFY4q0pzHa871O45EBSynrwE0J+tl
ENHgjssrmkMfQ7wukSSzPPUtYnig8Bg8FpU5sl8Rltxq+aYv3/LghWC51pIK
kZdiW3s1oZDUGdhLJGp8BE2xDIe9Lg4Cjd1w8zoFR8K26/zcJ96CbKWXA2Ho
I+eGDcg1rCV8QxotjSuWsxvIe/wk+2FhRwP40n0Z/7sVgo7VfR8D4F56CTaC
ArQG5NdFvn/M6eUShmA9ZQWgkLuIZ6DmwnJ5zl9/m39p+l92fVPIxbEl4RwE
wEwHadg0blsf7dLNrKl+4qCtt2s0DTAUYU8wwl+dhQA1ACzwa/2mRV1cXgpk
E4zeXBQyQYQvsx6nvR4EwJ0yBsWrtT41J9qf32fW99bU7K6JwyYNQZ80PIAY
YiX2hzyPnjaTpdCeEVtX185HOfpOtvBUZJTzThJwScXunKOl75VPqnmwVGoE
IF+lkBOzoVvMAozLJZ+uuCMyMveqpLojrPy6wYfaQtO2xJrSfPA0+p6Fhf1U
mPzfKWZExOYY1rGfWz5ZxjRsa+dY/VasfxLNK4y8+75NMrTJkRkGASj+0HTE
lvZQFD5p35l33jz5Sh3EniMojz+11VBBRApvCxA0YVtJ8zlnAkEFGECRr4IO
ce29hnoaD7H2OcOfivkNjLqu7/vzdMYu8t7LQG9WzS0mma87dNX9UbGdvaOg
L54CFBAOBxUX7+KmaE73iJakViI5EDt8HDvxVGB695bS8Aeg5DbrPk+03zx7
Tf8cUnDDjtnDrIGotra9z/vrAIr3ogbecAsgeJOT3w00CCFab4SQdyPgNQb4
wTfnLbuWNqnH55Tovssik2eul/XLy5gh8SFCpE+0ANgmWlyj/GevXTNAjhWN
g/9SnZt6WYef6kCP8D7k9LmfVOGfZ1JL6fq+eJX858fDCiZJ8dm7Rg5JA4/z
qVufxSyesJpOjloB0Lma4V70NZ3WSGhqCau2po0gCczImYxvK7xOwsTb6Dlp
IKAeKMJX3tWV20y6UiiPnTcJv6SEUnIAmzeoHztnEkx/9wKpr8A7e5ILz900
IxEvm6E10axJH97M+hRxBH+ooK22pHaFYmpDRUpYwoX3xfQodn+uB34LJ9oi
PqwsPDevYdVwqjY/IfZ0TDypQ9fYS2qAsqCMWg5ex+96GCWYznaH0pjFCbAM
gZDiN8jla3OS5Rfo720bC7KTCTXwmmuRysR18tv4K/alztHr5Gr1IvlZW6XG
MZB8yprbNO+ri7wn2tSu1HoYzoGDLcfSW5RqsjhKZzAbLWBI7Vg5TwS6Z/vV
kQF5eLXR+2sHEJzoOj6eWxh59BQKaD9va/nKr/RLrLUc6zfR3yh6t4csVq1/
i/ZAxTjbfIx46AvQgrMizJ/C1xbUQbGmkg/kOQ/1ZMCnOFRFQ8ETTOlDemTH
pmlhQxxDX5lyYI1vHNu+BoAjuWQ/ZggfCXmqd7b1tr/k/2jsfXrriG4m2Xq5
0TtDz3o/v06Z64zeHpjS8Mt+2Z9QsBLDzcIQqyqvIAmG0cKRHcWe4PPvnLyn
HYjs0xpCO/Lc4cHoX6wcboMBWGWhJkss2wwd5Ft1mGPTA5SEEDS727wLXatK
dxZX7V2ubmuFunDQawHoAkeEbOnsPZhqf6aqiLdhrpEOVS7EJMbFmdDRa1nJ
G+qAFqofqEGg51eHXzNRW+5c7KI7Wh5T6EI7Es9JlVUpAbyqlA1ngtaUFaHF
vyfkloY08IqdtCveBuXbzYsEZJOaTo2hIHbzDndcE/jniKbyvjz1HCnKI92+
iFcBBQ+qcTdX3Vpbiz7SgZtIZn0FHXIsWtvPIPxZrc+VAZppvHO8678ERx33
Pve43r4JtqyYWVXvxCF/qrU9SIrnydMtrBBO75Gq0ijUGEc4/OGk1mK3Anj+
IntKV+YBf+NKvxRDfggx7FSRwcZB++mqDEYI1JVljX48JLViKLSU3GB5QELj
wkyCFk6kbIdIiYfANL35Pt7gv4x+jPNcErWxMs9BLaKoZcI2GQfi5+dyEzNa
sXJehv24jSMBVCx2RcWf90tVK+1h28tORwsthYP7mn5D6/yruELUbI3OK4iq
T+TVZiom6J39jWVnXw9ByrytVqghn1AVUr9U/H8dMjJFwUaycH0DLfpBkSQW
WyrhLW7/Raj1Acy1cZXWP+ojGDWiD9QrLUvMDSRaqbmDS0aEgb+Y+PFpTlrp
Es/oajPzB+ke+5SWSaV6YEJ33Ckfkl5k/IitQ9TX/0akEGv6FhCCY8oqpCVL
aQqY+eTqzKcEuUGmQ3HVaoJEGPbefoCcz37BjMeBzc/G0y8BF5MpCcn9QwMh
j40QEtUH4+XZ+pWK7QLN+q0Ue9Kf8iJh+3pOQXaAOT0RugyPkTLeVqC09drZ
zhb7XBIEjYdras0FgeGhheiU50J3M9QIzRM12DCnITxczrp25pafXaul+9wd
DBkKLLDwFGEmOL7+oJYRBPWA59Hcqy0oL257W/Un8QtM1KO3yYcOSmqtpx+J
zu+/jRby+c3jsqGQD0Y/du5xK2pPI2G6IYM1GPGGfvdc/0l8N3PPBIgj3pfJ
r7YZLqIYN7LXF02Bbt/EiKZKSTMj5fGEAEkR0B9uVorr2Xpj/ojMq6pWtuLu
7Rfz23Sz8Q6j2GaXLq2MZFqvTEmguy23J/ELUiFa4jsOV6N/zyJrKC8wTfj0
X3WRhSP0NWSAxTdqcJcfG1HxFjAfX1tPg5ltmTTVxWE08YSXgEdWq7DoUX5N
7MRPaaLUicN7po2AuDJ3xnbUpuh5iDM95gRiqclLH739bioo/p34Wi8HwQoY
GzdX7yS3tW+IN+cta7cwqU3kQykL41WSbiwoJHvzhARDD977f8dwrSOVPOA5
3qb8/1dG9gmTwUNQhpYLFJjZDnwnUngsezwGFWhVSzLqhFBvzdGPQJg86aJA
2vRULQHVZlARvbeZ00fkMjyf7N9Rtr/eCiQIN3kOp5A4Unwo5HvyKNyN+zBD
OYb1Rb58RvMTU1ZOxceuDZJlnOO0/GuPtk+dVZaj8fEcdqOiXS2WlktoJDpZ
O2KA7BNlNCcfwz/auMyXeiGAJdvZ0P7g77DPO4bUNcyoh6V2i5Ni+QQh+8sq
UlIPsxywSwFbO2wwci7Sx4jD3PgQD0OM3hz37Pcyj/EXXMzTitaZb4+teY/G
4ck2VhfshgohafHIoYWUHnLeWKFdfjHirVwSaueT0bpuNuoScO1nV36D4NsC
L7rdld13Vl18hAO9Mk2PHOlfRMP5tyhQCrseRkHlZqsGmYD8Y8npUZNeuvoW
RBSzrDRzfoKoTIJ8UOiYLzeoYYu1mePihhYvsYjy/MtyeiBI/I6zhF1R97vv
uNjqRJBvrlhYXy3HhqBlORbgrplMAd1sJKYyhPVw2ntEY8VsKWCz/SNWiyiw
Bprq10pxptMAp+jAc4JrQ086rydZZI8usltEihDCVdsyGxPt7SqRLs8NDkwX
HjWRiauyIGtYOIJ6mKD2hCnGpe8Y+EHtlZUYo+gRG6zhEDc8Xy7kkNKwEG9/
4TRP2UsSciPzbLw7fRpBGB6oO7wyHhJCBKXnEospHCaLhbr5UTURATxXwTAA
Yidv1YCuM8UF8FeIgSAWw/QQ5yPkjMa53zcuIOZfHdPo3mg09sToWx4P4Wdl
HvF62kNmPQew34YrFZGbBFEvWGOUXtSmbbX3vUSHNntpGV+FE+RFrJpKND6V
Ah3MIE1g7cl7Sgtbi002+kkKUrjg+RGkRX6Xrw4MHYK/XE9xoggpOiIQLSPv
8BtcmfFIQ5Pt9F2Cq1tGFKNyYLZqUIOVB9vmeVwaaUdkm3qe6+4Q7RMAW9nM
B/RcPJj0kT7UE55/pXAwKjMgWKRewumMEbQF3pC3twNNAGHeeztRFeyp7wHW
m4n2UiwCCnnYuSEalv0aoJq8FklHDG6kuTyB/qpZIy7y6pn+sqF1/U2TA622
LJUC3NEYGL3LLNo7dcmjdkdfY4wSbOCftcMxtMZ2lpiLFcA8Q47gbW0aNKSF
Qvcu+Kg9FKY11z2ab6bUxpwRWJKf+BssP35lKqW80gOM36liAGrk8EVXz6AS
dKzdrkhR979U1tXRf2ff4/pKh1XMov5lDinc03KwYorMh5k0kpSDNtfs9Inl
xh3ChpLdct4nbH1lrs17vaZrCvh/OVOTOmXAYrVV00yVf3AoLkjcwJxxCgwm
W1uwl2qynU2n9lF/rNPqx/2sTccYxTMGufyFYKrzbVh5D172D3AywwQRLxkN
GrbszP8jiOnTf4W065kUYHd/hOgGg0FUNwvbBDOWyk1SFpXbHpn45iiFhlWm
OqFTP0wHc86ZquJOe4Ah6CBhN60GvjsllmxYDO0Gdn5xRZNAspd4p0tJGWMd
12OJOtqbDbuSwLEa78nlrDjRzIrj858U3tM035mow5pTo4rYqNWzn3g8Qcei
5zm4nbfMaKfWLd/B6mikANZghABKukXWUmhf/RbqE3jqfb1+zkFoOd5CbR9r
Mel+RYZDN9CU4SPvgaoE85F7E6XCI8IiKSNX8PTNBldP3c08bqVe/YDN/ToB
xDIp7rbWXgIY68YPsmHnloa7gmQ4KsZGQYN2No3z75tcu+YKaYU8fLVpqFok
ZPf1ElCbjmh3dNu3bx9rkL724tb2NpubD9Zj5bJuAe+VXgmwzSG8T4Dwn7p+
DlZmSnHH4QMV8H6d2H1f13wzjcGke5JPeoMyt4Wq9n59OXtZaPQ8dXTDuRqU
mcx4BmcfXnBH4oRJdSZc9UOzSmfKUa/x615TCpSUONrn1JJnTJtjL+1++iHO
tTJMS5aOzSvdpbb4ifbRmH1nSdtTEwUjNkWR+NNvqv4ETd/hf1sDikuP9q3z
H0lR5kdrVNc4lwj4pWeWRKHYCXDcNqie0Qdrp7ZsCoXj3cx03pyhljtIOxI6
hIIZgiuL5iwgxOG8ieXQaQl1R3s85QpmGG2HUjP6hOjqQVzcbMdmg5xLR2XJ
/80BYHbDsWHCdLr7Uf+UJHJlrjTYSz7PEoLbx2/hP43joIoZknDPBRvPUdjD
jXfAQdsUVJXx8rZ09aL+fMRHtHvN6Vbtu6gzegEmC/08SAyIwu31Horb5F5T
pe/Ngf2TYL4kJ030C++Hcdp4QC9L9ApV4xLkMK8iO1I/z0HBfwNpg39aQGrG
s32+oRb/KRpg4k68n4xl0yPUNDILuVWsPAAX/YFqVm6iOb7KfcBGCvIbH8+p
5bZhE7BLZNhhEHE2zM3hvaQSXVlQKt1bBdgMn5yghQgyoxmAmSFmxLD5g26h
cwZGoSqxv2pOBcN16Q44tcbcne/hZE01hTGAmTg7UmlS/Z1zIsB8a0KDAP7x
VSIMI537fdz4k/4xwJNYr2/DouWuFI6vWn1UTp7Fdz8F0F/FNfIILarFhQDl
hOPt/Tb85sIWNxi/Dn5qzxEjKL013dXxBchaMOtE9a1JowSXO6o2n8uZql3h
v8vaZUcyiBV1Ec305oDypClmYc+fDnmBZz1X9aWk0rXcxwMDwLZVMY28RHGC
e8bF9nxvFprh7dpj1qaDOYXUTiYhVeXn/v8ZQ8LQpkv31gNVHtG03mtBdL4A
Ha+zz1SZo77OeJSMpWccWs8DORTMV3RH6bDFu0VEezh7g6PaR6h16yuXoLMX
fRAbfW6JbhA3rVs8TjFdECnxENAdhNh9fiabec4n+aBKQf1J9l0rse8wX2p3
g4Ikd1M4NXKMTrM05yWyLfaeyJmJeBf0EYcS6mwOjk8n1RZuKCm+PYuAWT8E
mayQbGcHjALFwIcm4oXEXQKUbXITkG5W5PDB8AgJfMmgd44yzzCSh1IdkWed
ls+9bhcr6xIydnM8zWo5zndUM0qLiZPfcxmVyfIgDpDPe8gnN5aYbeBAIHaL
fQEQzagurkPsEdgcJjVfhb0HqcHCq1yU6kiA6cXiMuRvRaAQgtHu04jNBMPi
X0zmNWZjni/165rhNkSjHmvXNPchH1kXhP2Rlj/tr3gO3ngc6RrSqFB7g1ZX
o2teJZKaywxoRGtCi/ifA4RZXijVaspZyGEoiNzc61+TPbTzOy0CrwKVqOBZ
0TRngXtoaQiP+lCaXKa1ROnmbYmtMiK8ZiQq4Yg87Cb979m5BAZ6yXxl6Pht
g5hP8A8OZ9hiyPou6d/cWs4YEMO4Oct03c1p3BBWt7I1BeEEL4AFEBOaqUij
xOY33XztfaC8HkKMe9pJ95Sim8caEP+UTn2Fqg5sY1URH2Mj0jpwNAVTCcEK
L7M0hFPDWw1ciNET3lDN9MN29jRbp1KEqJZRhcjbgqwgmGNBL5jmE07SUzni
I3T19Cz1nKHXlDkXKJeAkMC87HarrYQa6QZkZf2jioSneD1mqWeaSRtF/L83
0bANoq0gtcDwP26dO+0hRw/NVweT80m6JoluCkBdDmHEK/5ZyfhWVi42BdTr
r/8FbTaQnnTsqVxIU18+wiz9+XLKV93VHZGd2Anflah9w9ArN5g4FjFZKLT/
bpnfwIjkpI6ZcwJoiOMheB1/T+9vV9XqAfpwqXkN5C8FJGesZmRvzH+HFHIF
8BhTHL96j+Xl1oJ9AWzWRFoNSUU52lcT57lbvuny3IheQ+M1/YwYKrQ5umVu
lRPESM8+KPH2EMq+QzPXzk85I0rBkkvsBKPGRr0P8rtGfLIG23LpzMecdzT8
PGZee7PN6Ia+4v5NsLv5hL0mPl8GPkTJk1TUSuo3t2ihWuBLDtWAwSbEIL1y
Cxf/KVX1LkNTC9Q2tbq+UscHNVAHul3RhuX4ZmSlliK9IOTGCc1f71Du05zk
Z8+swd6iUNhkcvh4gaDu6y741vpLACx4KTjJb2Y5zGCtIPkTf3eAiljUmGR3
Tv+LfgkOmZc5ExdVwQXg4J9DE2wyNxABdrsHUTLyS+aOB0cshLsQWcSoqcUp
dKhWukkKrT21YJ2fI9tFOq35Ex6XnrX/UiERpr8PLWYmedVLc1BUGqDqxTyS
FtOqWdpdTk2RAsxy/OJBI/3OTVYXWO/u5QA6y/zqi8eApVAwJogan8oWgbbL
bs+Ic8AcUU6t6XwiAON9q9Dg07bQKJoa7GPJceCrOEu3Ps9YGarBV8opyahE
5LosozmswS4KCMZ0tWh/fICSsmAoJLufvSWsrox5/9lONMhOIVOSb1JL+Ngu
q23YfPfSEA5d3RGwcAA6/9MetDwrbNOrQn0z6JKUfJnt1kgA7tlhuh+vwqg6
tdttiqFAnkOyvaIoduVMkVh3qJU15X0efe9AQPjI3zSU3G90Chew2YrUpxRt
zpS2zzNNfWCQHPvgMI/smxEKmEI/chXnUHNlrbOsgsOirEqPAu1ZNLQFfLg9
0iCqkln1MZ4IxHGXRQ8xQmfEFbOFwf1y57oFITG7Rn97pJvNRwCCX9yK2rvj
uhKZgUV4lG3Zo8DqYr3nbaYfTdDMny+gneMHtGWW74rQFdc9kKCnG+x7LLrs
AOpmMtX6bwJuYvE9B4YqqdKsRDoDtu+5123ONK0TKoBJBaofmh9nPns1Rftq
V9QqAXqrEVkiIBRAOZjJGKsDZNl8JjcOImBLGEuqnMls3UlFNYSx5hiAAt9r
iHuL/5dMNoqqEBLq2v3jRQYGkKK1oQ5u5qYB8PU4rs0e0e1z1k7t7oN1nFyr
QOa2juTTzBP97cmKXxlhtFnfVwVmteMeDK6xqTUDnP+bmy7zsPr32aAbONXZ
3P7bhq8yBL+IQSoxsCDQ/KgYGMsCecKfb2MRi/2CdhI4wtbIPJ4vC/YmyCem
EDULmvAWJuXBu2IGeS088wQq2tqRpLQFE/p3j1mbvJ/LWhYAFvFzxW1WQjZI
hXOkDANIqUodSTePPpSGiHEth6fLgwexDQQBmMQucmQ0NsDer9YMssjZmQdt
a5gly3K7tcg3edRdWqo2fIxXTgYMewmXvBh7677CnSIIjLcy283WNSjbf/TD
42nmAR3SOhMvMLU+6HFAKA7ZqhkDc30DlT/CvCKuhHgsUMwDThinpubJY5KH
h9ctzaYHff6IR+VfjkfVrZRJUKgrY2sPjqdPRemZK0Z8fCCDMHC5k5qEuOzg
bTQI2GKfdrA3mk4x4tWZvR2CbPxIUkZBVMf5HasDHLaEvcQVKmzeD0EpZzmw
bjv32M51eT/u/WIvbrmbYj4XxZNPfWC2mpcckARtdYpU78+IDvNe11xIQF0K
4EVm9er0bY5ww0FQ701Zx+y6AP032W06K/4HAK+2xfIaICqVSqC6rUHe4fp5
DIVPkyrCTg3DDhuzUhH743Er47SlKBTYq1Z0ogyR5bG0x4nRzH+84h8k1jkY
uEtSX0f9t7VNHRasQ90LQwIpFM1IuvvbFqUdLBPFimWkkH6zecUHF77J6Zc5
VoBTskluqJ1VlIR7IZZeDtYtMxNSPpZqMWtA9GMb/uqZEd9E8m04BVUVslWe
yvFU+771MclXcr4otEUOmOJFYc8pwkYZlSKRBrrP7gNJ9gSuz6CxmdqJkxhU
TUFYQ1xU8CiDfMKZGYTcGKXbGZ5I/Z/gFwntOLjJivLIF7zuy4DYHe8Mt41p
1uFDjE+eQKtQ87QRA5wim9JiJ6Zhp5VySNKNTz1DtG4z/wx/xlkdlDPMa80x
cgqYPWz3WaHQqiomyTOdm0xhhhhfLvKe0WeRWubtACramnt8FSEqfWLcj1rm
e7Cxnpkopsm5x/kJK+KHI//TUcuLMrvKKjYnUuUpQDb9FRJPllyoVdkLnMvx
sLO4o2myIQR4cQ/wO6yfOv0mhQlNacCcaF0Z9+4RB0PjsAWbaActKucd0IoY
ZWh4WkqR9s4yad/KdxzRkWLjl1M0UTWNQRlMI80Dd/1M2VQ4Q3TOARf8Yy5c
9taTxAsWDsF/FKwwYXhZfebvHg3e7/Z0ZCaMqaipxsUL0lqydtXFT08AIRnR
YUDg7ZI1Ems323lstJ4j+vLTUS8iFjBp0qOgoy4zU+/6Ke8Ry8VeicvJhK8P
KZYjfaygKIPd2RBOf8UbsUUSUrGzXxRrEsx1SCQoPSqlvGHIzo44YZtfHCse
WbM2gKmkrCHd7Y3tlVeZsRTtP/dqgEfRG5ounIF0oY7DegQx9MyBbLiBpW4S
HVjwiRDQ6EBiEMa5Kk5QhVFwHajWCu9Y7SmCTyOPQRYBqQPwyv9C7qjuxUTj
yfxKm38dE1b/LRQ095wrGMx+ISfRwKuaYfOFEWNs2ZDPSDgd9aZCa04Mz+yK
HnNOIPty+q4K2uu5wgTgCuluUYXzyp3D4wPDpYkXNstrYGgIsp5zRaDuItjj
zgMVe0oOXGmja/Nj+hCjsypbpFHieEUE7kwY2yCpS+Trf0RLrZ4WZiriPXLo
4cztkzyyD0JMJP33ikV3002ffiiW0NX/6kSINSzgVVC/1Jw+JbdLq3GZG6Bm
ohYrIDVczSGE16bXRitnYKDUnO3mZtJ96YyyEkYkWkujLwG24zsPSGizJd7j
wlM/SV2B/Q8st+ZJj0xE1wR9ZMtFyZejeJghOpSBtEavWqx9aNQhM3Ms9ERE
QvDt7nGB8wIA7nT7hwsuInE3cvOMXhGNqrwYV4bx1vHtnKrhMSocE6qtLv/m
6E1krw/EtC13ZcJQofn/IPNv/j/EjmNSKNmVuXRKw16+3zJeb8fKn6sL2R3W
sTHHMvjZnBtxxNiwi7FT1XEn2jVvIrbjJGn7WC82LvMH6CZIF+opC5ss/OVB
HkmWveDwe6SQl3IZ0Q97j9cTsMqTVCEACxatazeYQq1LQgfgrYjfAnQlqfi1
PhXSQzJXCCguNbaongHZaP9s9ZxzTd1LxD8NcYXwGjHNVP+55Wc73lBcylpv
cmz5M1G3o1xLm5ZIQyrnOyxKiVJ2rtaXzDFDnM/km/XHUgTsQL5y5zVXvmXF
Rpwam/FJ6NoLUismnwxHPzTqV/7opqc264N/ctoexI8XPvvew/2EYs6+jTxH
mQRFVNGX7CwLXXVlZxesCqVdFJECTajX+Gak1oNpFCtFReAwzEEq3VbvrUK2
SW4fLLLJwh/UnEJDaycmea52Dya/lrWa2ce72r/iYPFi+1dKdrVBJGB1oV22
gFwtDyqURTkPe9/sVZcnnYtKE2c/DDxE+idJrliUEuE26O+7XCNYXNjxUWsS
MO6m5R8XKbntbNKFx5YxebrF60RKf7aNB20TRQCVSZ3HzeODGsGcN48QkKw/
OlxlnP74FYRSSj+l2tVBKjvhdKN90lQVQSzEFYikuPK30KJ2YlV97OGsGe7h
DEOl/As++tJnFyVwfKjbJiBMC7+mh4tmStE7ZG5+a7qyOsFZrbcH0hJ77xN1
07nZ8v4r4YrzP1cQcIzx1g2X1oKbFy8mNInBn+4xSnC71TcpecWRBHFnLR0U
Df8g5P7yIXsgjrfGqu6LU5kK/PsOS76nWXCLL7inGVmR5qzlh6EJfHAINmRm
DrrJmRVucFY311beSHVXlOsEhs1bfV+EgRzWM4stOaFpv38GOnRoVPtjU+um
pFq/164W4vSEpJNMu4qwDQUqYJtzDXbyFLSONCPzFv7i3iOdJGahB6oaSPqO
9HWA1GQjZ9czGGLtK2jlise1XC7NRdtJPdxQhBOHqp1XC1mAQ1Sf1Xp+IC3a
zaOtkIDVECvJv6qtv1Iqx+aXBUSVm0iycBfA87ZdFVd9Qduek21ol7dGpgoD
KMUTq64wv3v1xuMajZWQwzZ7wxSNxrvypu+5GAijqylC2lnpi+3I9G7yyXQh
yRE1Jh5l1y6/3VDCLZXnsu6f7QFuNCyjgrqE81PfQviJ6BNAQVvmCfgn7NoW
rXVMmr9NC+ClLy6onAG+gaTUKZxUCzJGJl2XFxYjcM0w2Ti1E/sfidTLOyB5
aXgVpoP5O4IHzypNV78nzWG6JEyn5iF9tzkmQseFVl1lnrvIJCij8m/EeAUt
jJl7buETldNwK0PyqByokrc+jfeghJZX27orC3kJHpmGM5ucg62MW/HtJjcA
s10n0LlcPdantkKC1C9p+42gY/16Q9JNZsRgUhLHxXeFmeOfP6Z1tln6AvyO
YZz7wZMgLoqXsD48P0xbHwVCO9S6WAxO3J/jsnxiMnUf3/BTFWotg59/yG/n
KeCseGSyqrl3z+memU9C29g/UK+HKdCk9MCds4XNG1Z8+DbOcLoPSJI+haD7
ykdt2dB+ertSbM0NjKzjQCfKUJS5TTIOnCldxE/wm+2lziUFQzlcKG957Kgk
qLuHsi5IbuDChLXUTYZuUn87TIUh1kujkz9njRhkx/9rNbggfEgj/zNjm6F1
dt0hA7CazQL6rILhwx3Dpxcg1vY9A8X0sBgygq2FfOJ84ANDiXGbrnaYi4sN
QlfQ6S1NxcUcg63hUyIcH7ChKNUINyXo0pLiga+vxCbsGE8AVHQNRA2tvZ07
CYLG+LNqpk0nIlRWlmD2xZ7k5tYsh1/3N6MJ/ZL/Ec5fcdbLrmgwV0hqsEey
zVxwLUScUSu7U1O49DnKoVdHKH9DW2pwM7LtMe3h69au1dOIqkueujgTcOP2
8rwDXEWctX7fMTRUpOcHGGkkjr0267licAB8NE7rpBQj3eMvXcM/mdlhDnM9
Og6+yBoJRymBg5YLOIlOdBQc/wZJlFeook5BLWgVvyZy17Oa6noJ9vWIo4u0
q2rd+NjiOja4huID0MVL+GhbBU5N7RnHC46Qx4ZEZ3nKuGijSwkVvB7iAQQ0
dCRlJOJGVJqh1eoFnyjhG8BQHq4JyKHXdaCoK06BISbinSVYu3ngJdzRIycF
UbZ7WRAy6GyqEU4dbRVfD1X9stvE7u75StmxRCfr/9IFMqrvO0qtVhBIxnCN
vnSqnKwaF0iSTw/iOR391h1htJea34yu+q+w0wXzfONJuEfHFO7/CjDOH20r
vM49b8ruV/wLRRGjcMu9BHbDNS18i/qEbWOnpsK9xwETQIxjk4zaCO0RebtD
kjHOU4TtWUs0laTLmXSNoZuHxJA0wNHcdt84Tz3ELRwGV2VmvcJCYQnisk9N
qk7H285YKWINO6yiDbwt0ymDMssBmvP8X1yekQBvBdXhpwvIK5ApizDrz5xG
QOXRNtvdeCdzLBbd8dfFTBHLEMwhRecN0W81mZqK2xnarFVsr8PJm+obixJh
ZZhpFk/IvBSYG+ccPgS1cjR7Vj9e2qEhkzvrC4T1ahdLP8zgTnG65rgngthC
yVRoILVU0b26m7rfUhliXzMb4cvDgrOk3uBwcTdRDJn4K5JVAP3fYsPSfumM
oX2T66lClB/hhonXJ8dWYA5OxYTEGm53mfLhFUJITyjPRlVcSyvWHscxgCaz
+lv9lr0LOf0WeyLVv5MqzS92MqLORyWbpTppHv/wRrpE4MNhhQcwUJd8NAr3
vYgVDK25V+sKS9nKlaawesT3VqdI8YKpik5804r4BhEeMiuIVzCpfT7j8gq7
L7iUyIjLQCvYdzt8fR3/eQghnLjba33BlTOdnOHHlkZb3zMDNqAmW778wtIV
cXhgHmSM045UrF/BCuUGppK3N1pg1daBpX2s7qpT06pMQo9wRA5yZCY4xnF/
lcFsuzXMEUH/N7s//1k5/i/02UkYDKBk28SoEnovkguYUdMnlHUgosCTtRvv
umDm9k16jsklLiDl3H6/y7/V4nUoxS+rAGS0BrBrPhdhg0DapAImzM6RxCRP
E7QaVzoXm0+IVIRbQmsrfudms7qsPPZnUPWiZ0/BifjGWBPXt1zow5M/mmGn
0Ip5ytQ3eKR9Acjouok1zYBZ4XSWenyJX+b9Nq2cABBOeAlI6AaQMsf7zUC/
o5Aeu2pcwtwuNGK8ByPfDnJKzHaC9zZHfBEnX1HMuW6df7Ejw6tttoYzhBSh
JrJA54XLy+ZGOrYDlNmC/6R5X3qtylVKXv29CF+QR/REQWAyWbj361r0ou/7
D2ZwOCuuQI6nU2lOLjEXfxK89gtYrMwBs11Q1wKz+BgQ8iPykbcE604T3yum
RxLkVjntGYUkcbMACul3JezA0kpygXb3LMtxgPSRkPBXuYeHazjMO8kvPlZ+
sTcskQyusA2610JZLthV8oyRAa9NMoHZKs8d2FB3bNv3RWzvZlMZXqJ3zKaC
1cvpjpkxnVxhSXcxEMXDuf21vVs8Vtx97i2JvhDE5PGX+HOwpbg0eZQ0jpmq
Id+WaIv5aW1VRnYwznds66rnOPYiWhu4dCBOH8wT29SpJ3ZfNOOCa2ercKbg
PavBkyPT+BvEV13beS4LOU70+c6/4EEzqrvp4ryUKcI+L0jrMwHTDo5+Rwcb
pyOM1+AGv2v7zxQ40wfKpYPx6fWlOpFixY2hxEBxC1602tt3LbP4YWmVW+YH
TXU4qBZC8BJwaIY16BFgn7FC6of++tdXUqct6hFXcTOKhv7wO5iKtBxB9y0V
NSvPx0FKjvueEVhyc1iNO1PqtlIVCZEfpZp1RB6MJkMCknHxUkhzmISoRRcb
nxYb2N675ezzibGrpPYberlL0IymDeXtTMivPCOi/yCQB0aWM52ntiNnJykF
Adc/mvcF2820uNR1ERKUmaCwSQnp/LQqn6gYmpjZRvBKN7KvqEw+SuXgxvR7
om9vuogQR9uzMkaAt0k8P5tzo/XqLHStWg13/CJgS72xZhoYXSNHRMQx+Q7F
aaC+VFWuZ38RVCuUstTF8Wgr33x6NPJEBVyyfO10iESJg/Ey9m2jXkXZXea8
Y7U45S4hkK8uGZqYPq4afBrYcGHt2aCSWsCC/xRs1WaiqbfRU+z9DfrXEuLH
7hBomEssqIJyl4Lkrgzroxyn5tKn/C7/sauYSlBPEhtQZukai7ieuhDkmwDu
etowElvdUrEQX9VL9/hrEgC7koWG+YrhOfyYl/vwxpkdGwFDhbsfeWYH3RvA
j8lxp4sEVDiQlpw2ow8eaa6Y9DDVCnobn1WTID0jjKVkt+rPCHJXahdJzbGM
rqMrNE7Ae8tbL0AGo3DN5IQfiZMMkzrHPQCWgMgnXYi0qPsZafnrisSR4YW8
oFC9FWfQkmITZxvTwbz1m+nZ8876VeVQ1H7vh+DT7AovwKyinUqC4h7AzsyB
sPlhm323fMnrTHm7ngkfOY0GBiEaIu4GQ2bTvfsW2Ue/XpSd4uvdMMb9lB6P
7kBJbrvz0prjXoZ25ugpKjxCSMzKK/rdrW3uGQTKVZNGz2TIsf29Bu3GNK0A
qtPIrrcwgoRpGLPXL2i5tN8i/DbDRixoOxeJ3+JJ0LZdJ3rYmqG5XQa1yTMF
BC7Z4ILgiT055vQSMbipXp8UYjZLnp4Q6/TREbBw8NA7JSHu3sO/YO3JEhUt
K3TSxleXvgV6F+xD2Ggn8ZpC8cQI+Cor6GdFs3Nfc6ERzzmBeC8KFFQx5lI5
1aPxdF8LeEFzX3dh1LHfmZc2pJnMpncLZGjt/mZaiQJnpUzY3Wl1lvd0lKgM
KVlBQulVz80GftmwiAXL3OJ7LuzsCArZtyHGujv14siWgmIFq5FNJqQ9/nNb
mGLzxv6kqCaGrH5/aOPXKKfpc0ZeI1k4cPRMM71ETmnfv8d+53QfWNDdVoKj
Dgs+nRraAz0rOek323xDpLloyOQTJAM92Gfdz/N/6Ip2CgTfwohVCLFSg+7k
m2tUsrnr2UY1j07cWronT0+Jr92n+ZfJdIjybWf2Tr8zknYmeU03RKBQ2nN6
Nw/lJG+9kGpDimCymIX2kGjsH5xAds77RRcpIaIqkp+K49lh21Zk9WKHc8Kv
/hmh2H0m0yjihrMrUntsiv1RjvdxRZtcE887whuVXjX7XdhNqeVP1wc2weDR
NMQYc/YO+N15nylcYvLj8/Zm4X1MTniEmzBW8C53BshuAwLuNWVbHcYOi3V2
QN0UL41IQnyKSscPjYfM5KleO5gU5ko5I7i1GdqOwjvflii2oc1TI7mz8VKq
s2Es96eCMdsOG0HmIiTkIKUMTbOt5tgGPrjPVzL89+maKGyxGmNmN0Yzl+4p
qZY1GVz2bedINpeGGJA2A9+IsHZ3Rn9szPBX8ax1t0xzlxBerZomAbD0JQ5A
YOPhjbC43t+c8tko+/xlIt+KJxc9SpIshzMqToDoqMPZGi9WWwDemNGHEhsm
thqsLKT/m/6KEoQdMthvlcbrsGvYqE4hccbfDklCwutxSqVzzHa2VVjKcj6Z
vun40rptMMPDSvjFDbe5pXs4m3rE/Cjv6PIMo5xTC7HAaMlbtK/xqtqX5pUO
K1UF+Rno80pLPkL8tnVfOTEOL24WbIzcR0ABZKgwQDDBzNI18G53hkk1dBTA
WbYtUmlVnAG2IB4OzKc3WUHKNdI+PWHTPEPKdZrYco7pQ8zmhqldjXsZ4nsT
hJ4D7m2iKZkP45hNMLsW9y1L3HOY9FTIvR/diSio7VcFY3EbiynLDhC4oQa+
H8Mgk/wFezyKZ+OUJDaUmYI14mcQy9o1xRXjli+ce2drQNSBnTEbNvnio7+2
eAR9uuQ1qz/4TlQU1j5NsvHX36KYpt2a+5hI2DD/eRzf19JaC/YtWSpi0Rpx
ZLy4eurImaYA7tnCoNlfYBp4IpYq4dSJSOrNW5uKTgDH6jhFcRppE58OWsGC
nQu2vFttV7oveBNAvEKsGvDGcRLe7VIm1F+Chru/QpzBxhyfA0LPPhcp3QPF
wogperRsK635+bTPB5hAVYzDKM+f4OLJqX6bG9reBkwjsi8b+7h+S0udihEm
o+wq4UG57/0Q2Z/4FXES9PtYP0yzsrpzXBZ2idKM0+8Ua2iXdSWQs9d4Sg94
tmkzMxso/MwKo3SosffJtn5GZfXEGBJMGJ1LPS8tbizE1D1uZD/QGpytRKGm
XFSY7beNGKoN2yqNWSBJA+dmWKrQxCFou2WY5+5Vci8HIeOJ2TItNe5BYkQ6
m2OUT9vlVdnDT6Knv39PgiWiFrdWGbrL5ZVEzc1aNI5IqsI/w5IT5Vmm4b1y
gsTzziFk+OQ0cHItefieAJCbrdjEkRXTwQVew50DA69dnABpF89395N+h5W3
OF43Erojo4ZMIKMSRpAHxu+GMWybzBk7ap32Xlwb9+dQXp0keaTN7rYTgBES
ssCiZ6dj01VatLJCdgmzqPVfdNsEpZv69T4Y0EzW7CjxdA16vrMcr90/x4HA
sRivMjyle/aXsouc8lWKRPHzzIZLdOQo14HDvGum0ioDPkLx3hdLt6zxVjgN
86UYVp6SAVxnTCrCZNsAoxAFLR6mDjT03EAeaDtcB/pFukOCdnlSlzcPs5HI
UO6fEAWWEYv8pEN56WjsqZLQQQ504okhGtbG3ZzNr+oCwb4kuf7gg+EbsJT2
1bewYaIKoS6TrAyfdbm3WewACQ9lCku5bCKPEIKzahiespfFQYg0EiIpvOhr
VLy17PvpJv/jZOaKHniOVuKEk2ZbCnOZ4ur7RxJ7GFvSXEoiPCXph0kJIA+6
+455bNcZCnCyDA0zafqWzOU5vQbx+xMuzHfyhKEiGpJxju5IVOa8tEYvKU6V
F7Eql0JBzKJm4wLeEYK0umAaSrNXwo4uC/qtWvo+XXhcCLLQL/xl1M49kbvj
TZYP/bCrEc+FxpJnFQxF4PkRb0L/3TcYghOyw3qzTNPr/QXK4RaUY2dLSkoz
aeka5h6sR/jwjE+VTFjxePmSxMzPMTwXBRannNzOzG46UOLg/K43zj5s6bx0
tai13Un8bSkHMAaB/O5Ize+90UskmfP0gAjAB8zMZqfjr6p4eOjjHpHbBxfR
Xr07LKAdX+L3+ybWDsPkil8gybLMfRpK4pY7QU6doUQ2H07Z2qSp03Qm6+T9
48s7G1kUFN0WFMEUP/E30lW3gJeuHjqKhaRMdsQgf+n2QsM/RkuuoQc7Mo5D
+yfCoDlBMK9mXj+3zgPeTZ7rHU+L/QT0hHF3XiVIllzFUfP8pWR83imb8doW
TqtOjO8En/8PvMM7u69JNO9jCsv4PVHIsGI1RYMz1TNRpayyjA/Te8qUfXUe
oOUueYGzJ2AWaMv24/+Lp0TVLzsulLQgL1XLSPU5LWrxDL7JLSOKrUW8/18e
suuHV0IR0pHMYNlcCHPp6/BMvUL+LYPq1G41J8d6LlIkeGTP873lBd/uYkTp
Rhzh1/8pkwuYJDMJyZxfIwTuq1no554WialnJcR0l/vbPcw8Uz+q6w3npN5S
uY+fa7A+094ONgPFRwfQDUQn8MywdgpFgPn4ljtLI3yOlPE7/C/DECu5j4oR
1W8Z+DWym50SowuaX5UgeFh7pQywZ4d+iKrRA24drmggjNbroUq5nghiSs94
N0RaU0qSZ5MujICYdmNNT1FvD2r6c6nYPxIbPI1nDm5eqq0Uh+AszSm7W/mv
JX4qQlSk0OgyIl2+YDrfgpyI0AsOP8Z+BZXlncKVbv3cU5H8Pd88aSOJU9P0
2wlH9Qire9O3I5GsE71GzY0dQGEXyoKrj6sw/8j94jYSlKUq+Ey+33SVLskK
0ii12rDvmUnL22f4Wm2P9DTtcHy2u4RARXquzm4sULCmDzMVmlaC6SLr3M5x
gWhQsWdmwUmAkmVIy31A/gDGKImrpgsnZnPWkZsXXDayVvdKNTzdnUn8oKC5
ctpeSSqYdJFnpgpbVk/w8oG3IPRjYQuuGIYSuQquUBHZCEZWWDpSW21nA5PE
GbL8WJLCG3y2gpjyKJDYTMxYEoH22Cqoz9PvcmyK/olOv7L48t+e6YSISHnM
thsUIQS+KYl5ebDiQaZ8RnOjPM/xKzXY1Lrkl5WHo/IWKRgqKeH2+gYXk2VC
yfn2VoGH3xE+K3CC1EGOd6cMyBNm8YHAKbxevFEDgjld5SFdAWCiWTAuoYW/
YDP8nSripN+Fbu/VATcVE4+WKpsPEYyQ1GjNlsU5img4au1fK4p735mtSzNF
hBoUD6ogerm2NVutlCGCJBEd6HmqAWRMh7PQQmuiD97hJ7ujzq5RPrwHy47J
6bXmZaEPgEK/wad710xUe8pp0dgSu3y5UccmpBFhrEbgTdyLpOHYPe/72SRd
g7boOMAHKI7fNdfLFuI5hthfyVsZnZdC0PocHS726q602BNUUnYyVmyPo3AV
/gc+xu7n1Y8u8kUh1J2cKjzPEmzbaw7LXkx2fx78Q6Liy7wyBTt4LTgDof4M
8zJsVz94wda+jsJkCgw93NFQXexrKid3LFFLSs4PMDZb/pNC7jGeXbTGkdWG
519eMOuBresFgZqtorTWAEs/FFqRq4ZZ+mccDVgPWjF2v5Br0qPy1SaE+bKt
yTsWimAnVAM9bToMf9sHFt9fwXRMAqCKc8RG/fJ4UR2vHLRvtDe7W+K1CGxy
KKmsxLrCtbQJrSMmF7yU7JVn3AT4ILkaMNGIchRaoIyOO5/2483BRR9QqD7n
1ZX8Wc1Ezs6VoS1BcDjkjhf0YvOMgnq1UJsQZSqllag8fiaFdYcw6DmS0zkB
YqeORF3HOl64ML3i4vw2zJuiVJc99oQA6sHzlZkYTgJMODAYAXxInOvWrvwc
ZpxVBtSxbi37v8A4KkHrkpTNSKJ8HyIEkZdTr8BBkHJEXqcWTxINv+hR7GuG
5vcHIS+xsru/EMQBcrLaN7V79S/k0jXfBDs8XnxrvL1l4Ri8BdhJS/qEBYes
x3mzewklFPRqydL+TjThYZpMHPs+sczflTO6xWW64MrxuHfWMdi7CuXbPnxH
mdRMWnwoBQDHB1V9qoqhra2tOUFNgUa/K+vezIGbEfCfBMPtJY6/qFX6Ro24
N1GkgI6v7/pQ7IBip8sokd28gynLzVMrP9UZM8GiSflqUr9YEZRPpDHXLuE5
xlAKZIULJ4buIknjqLX0R6TgJY3IcmjEAkkGXq4q/CjSFROG3dTt8puc/UYJ
MtHVI0qK5lnHBmhwp5RiOn75cuJ7apmUbm+hnbkJhxdjr3YEVCST6MPaJyjr
kgUKZ8rhIAIavjRBCQ81TaySA7INhIWvr2kNQ/UJ9CqubgWnkAKczXE9oZcp
RRWv2weOKUF4Vm6q1OzscMT4qd+K1FgFSfe7nsMv0iYYyscw7iUqfZDNm7kT
SfovtI3JedAZjjyrh5ZYGRDOys3AwjMY5J7vJJ/Yf0Yi821LG5pcRwX+mUSh
tz6he2HeqHZJPDppG82mMkQp4aegGWuz06QuiBqLTagbMsMUELQUU8S1V0kI
B36hhR/rKdDxxccmc5JJMUedAAG/ZM5QrGKaTnyQzwEnsO+AZyywOnW1qbwK
WJAueLATONK6aY26mU4NsQsoiAz+OoZPENVYZ4NKuRbQuMFSFcCA5YZHfUKJ
DQP0z8WLzyjp1TGJV/VB38s3luBkoDPyDe/9nvI10gANy5BbzQtecoPbPXLE
1ZHeNpxjwjgdBEJXzmLDjecyWcPyd2twtrcxVg/xZBcf5L2ZMW/51cROr2E2
aCVO3TnXvq+5b0dbhArjx2rC67Al+eyRuPdQ1AUx/b9KSNW4RX6CXes6vuHY
mkS8nDMIFW6VYE0s3P5Ul+qaFWpaotx8M59I1hKnqpul/+ycwnyxHVltwAlu
Uv4rksNQvhVoCpjNYI5wlG0XFubPEWF/h2ftDMGFNnELgUY+QWsGg8KmzQen
FqUDb9RD4sznTiILLxqH4u6A9RNlMjZKKdSXX4nLl7pC5PaVNAi9WYDiH/fE
tHJT8ZNm7oU4+m+Ub8fUc3TppgHFFIZ0+/Nxf/o4ficucUBa2P+f7mQLHZX1
r4xAWYlLoVwMqARNHoBA64VpUci6pym8M5p9KvURMWdvXhwhX7ViToXUpXGn
NBcm9hPrr/wWwF8zh7ksg6EXiMPRtfnhqOmX9TwG2cVlj2DOp+xd3/SyJves
YyAX6+YSrHjx+IlMVqQN3Ag+rL82p3eG2uWKlQOp8SJ6cJbKKkIdRu8Q1E5Q
WBeJ3wo5BMmdT2WudrclWYDwRfzca7vg/mQnA29Ug3MvKInFmi5w9LchSsl1
JrDUDHcr7ctQAc71qS6Z8Psqyl52ezFsi0dNsn778u1wdL1UX/Ysqf061rlK
QLi/0Y2lgRGGlN9Kts2qWecb1y+EL9kbs2ETdXYf06SBmoctSjUqUctOpEDB
BlMFzh1PhTdagB4ucGav/fMQsLu9XUSoGL0YKwOBSWNrGnp4WbiXABizY/3Y
xjAx4yMPFV75gZqe+rMJUHK57aAa+TlyLsg1x+yhHDQieX+QEXuyya3H8a7L
lEVscLJFrV4J+/9A8sQgsRsSwMFZ5yjhF50b1cjgvK/5WeWXoR0u0bweBdNM
yT+T6dcms06NCUSXYBwf8RqbPGdfcwQBNo7oS1ZgDrv9hjOpNIT26LgUUQNF
7OaIzwf/6Y6o85jHbz55YUL3bS6AsT1ZOWwTlUQD+teKM37s+4EayZlTSzLv
CONdLwoup/osxbHLQJ4K6+aCv7VIAJE0sqa22+4llydpfrXYDyR97mVXDp3j
Ixa4u+RFo17/OsBhnHRs8yQLoRJqns4261OpYdy5Jc6vUh6C3Wc0Sf78j1jB
8gSEYvSv0vy5mI7BQCbhUNL0HQghnsIgKLdtiH/xgRfguk/AiaOEtTIG9CCO
xPU8sHrG6KrC4CpkOjHraHjilIrwWuPgb8PmhOVazFUM9wp1LicrpzeyVqNe
FxOiJzYLswWaIthzlWIjTnSs4pbXPtNFDcFg73m8N4mUdWh/Ly3j6uv2Vi4O
XMEs5vOo5KNqe+bLQ0urLfScgQ9Ls9Ahf2NQ32YziJ1lHbwO0zvD6YtVdFCk
JPY4PVJOwSy4ZsttAemDQBWv934V1CZcXcD7j6KKLQseFoOxlcPjP9OnNOsV
uj82XxcnZc+sCA4pU0JynShrNcQ2FArsI/1X1qgHbCdJlLaM7QmAIr6Oxyvm
0soyAdOLgGDgL1kIX+SP4OSufgCaTIXZ9Mhocekepbpqk8vcafIGlBr/+u5R
Ql+XeTXhGGF2IcspfXEWXrHxP4DkJRohXbUraF+hQaf02T02FJ6PkR0e4gWI
SozW/lqUV+M17W3k4Q3adK8QP+zRxwXSirbWdk4MvYV3ZEeu0iwzeSQCMqUg
o/VZ/XrC051FdqF3aQlu+VEnpzNcKZpAnj4E3oYMlpl6k7xjD1vS5V+niNhx
uUhaDRV4sxHsFPDfhL4EXiB1SZBcI+jKhuxHWB1X5m66bnmWls56Y1H0tb4Q
o1YlcPXKdgB54jXLMTE9NkrMGldeLcMvYytmlWH5e140YDEoyNhKZvA3wx4/
E4ZKwlDCUfmhb3aNgX9vfyXbQjQmeQSmal4VSe9bD1IbUfPUxv/XnHIYKjXx
351BMwpB+dIbZnTSVDheYFLs5u4NtMsz+P/Hbyuzsmus/sFGbyxQ2oX5bctX
VDFI4n1ZsoMpPhhQWFasnEysMHo0fas3plhwwKjfQIVaHrRD6lSnn9Y0iQnC
BjwRibnz76sb/rfiFkB/mrfVxY83zYMhkRMJMUeTJ6M3RvMd83RTdTXYLl6T
NEGJjCoWRNHlGE0VoWVI0Sh/7ofKKq/CftgCHK/aWvFufWJAQ81yAcb9uJ1c
151rtAYeWVzkB8hDd63C00yLVh2wEa5HSeCUpXrhXnNjZcZ/656aM5iyyOEV
l2R+7YKEQh/9S5fBzoB7p2uESBkc8txtJMJJ4wjwHVJsXIKkvCl1ga+c/eFN
ArZM7QqfTvL5W8JekkkyhtnuLMub1zJ0vNK+i2YorQiEMDQiVw1xw3IkrrTm
CZkCNzwBpzH8jnsNBWrB+7+1PY4ktQTFWXZCK5oB6794TQThuGIno45UzuzM
cuJ4dnoouD8SdWWvBOnezAFOVT8yjEy0Jd0YTKNXvJX+A2ugRTFJzFQYgg4j
AGmfiosWOXbHTKXK+iHNNmvA+/fDFJX0xu4j7Mbui2NU3DLN0svM6LY/aQ95
JlFuW2ZPu9AW+TQa4Bs8Rg56pmECYAh3DGDiek9huPcXrYYjmpJudr2G6XyC
PZfuHQj/p/E6yoLy7YFC8QFEZA1fvY0havVGbZAbkr6Lln4LhHSjqk/b+lYz
50nFivshfQK4XJa3D1ZJvG4AHK3cwyI9J0KaSiJmwuz0y55FvXXHTanHFOIw
QMw8ZVrlcyPMyaByVWlpjEL/sXl72//ViG2ObDylUmTWFKptmyjXIH+P0Q20
BnCSQ3AO/I51etfhN2Io4GpAVQBDljRXBQ/2KAK12QOdrjAwJdOXhNDseG8Z
b2KDnyciDN02UxDUoZyIfV+Af6XK+iSnQgCkFszrUk7zoO1TQEgt0s59crZx
old3WtGkh8KrOpK2tHEcUTykWsZfYZjLiNmq9zZYzeQmMBgwhwHXlHeCIJBL
x1lj9g5FWrO2D4Lu2yUZdS5Eure20eJ7vp97ncgIDdfjDy6x3mic+7TULiBJ
+s9AVcbGkoaHAJl2ZKkyJg4Xpdgd1GB3J9VuHlrnUMD0/4VAZlB1xXps2mOf
VvcwCOImJ+tncfMCgkhuWTuWJvcnSMi1D7BlJ1gsLCZ5frUecl5rNIwZJ1AP
rFYVOMawTIBBSuP+PbdArfv5myV7Ko6f0srt/UYzDRNBb5RVPaIbve0A0Mde
cYcpq03+tLfIA2zOlvjwVGblyv9OR2b7nfEb+F7RIyFRBcyGvU0YD/xZ2cNB
eZm6RrDHF4BY4iSaLQksUO0SpqXl2Vr8WjnL87gJvhvjNE/IKpxduNdNSEWt
QY/Wp47lV9DXBz5s3lj3gaPEkEqxgI0PmrnfTZz2wJ2xUCyjOqn4InBJIZEH
aNlInfskCqmkw3ngOgUBYWmbw+kt7pCptm0Cw1qf8ySdSZYjptTcW5lOesxD
0t7UesgsA2IfvTJC3dDG34ZNylaKwK3p0lz88W3hanvOaIWte3+9WB+4rVLB
yNOPG/5y3FUCIQbJNXS3RNu0Zt3ol2zL86tzGA31k6whhU0BQNe50XhJe3ED
C8fUoPsj/OyB29F/74iirt71LzsFO3SRf+6010/yaoMgvSfk61uS1zZz8fPh
CYiF2K6efGQxxCnJ0XoMkxwY3zitTF7/RmszFW5klZ4CkF6lAYBs4z3Nsu0F
8feCEyTIZCCy7jEyWRJ/HDRwos+VEJGAX1rFD/tRVJJ+954Y6Qnb2BLbHYOC
JB2cR3MGdxggQ21VeBG9/Dnz/zHPJ+0nkcOiwjuMZJpiM6AcZ6pYMJWi4LFD
7AcCw6GO30MTVMh4094mADSFVI6I8IVr8ElHjqdoZi+IMrtWD6y80V7tfx7i
52Wg4CTqZKEQR+ZV5A4TSlpjA6m6n4PsZgp/GiDOp1pBBlDq2OzCvdiQP5qk
/vmazO0aKhg7sCR3JZy8i1/GQU87GndiWiavkYDcIqNkX/BLTLtBmnp4Re3P
wXC0XYWi60n1HRWRGvcWpFns6aOXQOB7RCjv9xwP+yPSjweL+uAmrkoOzxIR
AqpyoT5bVAiqbd8qBnK7OtxHwdokUj8QwAw3ZYh/sG5unY0qNi6zARBq2Jpu
sCex0SeO076VUCLzDXuN93vBSw0b/OYgJm6VWN+qwjKgMDQVE2xfP3qKyf+6
ACS2DFQkyHzmp1aTWXz8tFe/qsJfWKsyivnNfiKR2u+T/nVqYl9VXR7R9uUn
ZDOfWqKOteTABCSYuLpFwpV/LhLds00uikxqc6dxpbP0wcylJb9CUQRJkL4x
spG1Mec3KFKWTD/53rrzpX0vZJMEylobK970vLP2tl4UcdpvTV+FDPJ46Ipl
FYAWbUZy9lZPQHeeJe5mcDj9h5kRHI7qtVQpJosJuI7SvYfe2TaYeLPoFqbt
Xxcx7p6qmzcLJ2DlHvX+9wCpJo3QMYdnUMtrzo24VqtGklNUYG01GAVMBB5K
Q4QPiTOep8abn0AlWqcu37xptNP68ulpmjL5tc6JiyLdWewV+jfdL44mvhAg
d+87T6acqa5PLFnPjQVRqREKcCqc7fmAwL5MnAJw+gHiwZFEqIBKvmxWvG4l
m7zPNuYk9fnu9FkzvSZ39048Q5kCX5MyAwpq1pHbPJDNC3fRJB8kPCAr8y3b
Eu64clPxao5YXevnCWon9PEG6cJWzMLQ9/hPVrf+oQOPXvIC/Smx//14OExk
tjcC4AxtGxmBj1zH5ygXDn+pcF129cwNFINJm2mS++1V+uwffm8AzOgeIXxW
LQe13m7f/IRKg1woT7EaDAXNFuSMTQwvDwM6h+5WsNfwCfvVLczP3BHnyEdL
TsSPpf8c3a3+VV/sHGPU1yOOTPW9L3zsTiC9bwYOQeZvKaR51V3bQj4B26FN
4GUgx9hMnB7QPI0S6xp354+lWqG8SMHfymEpXcU04IslII7I3piE03FTI+VH
u1W+VNEu5VmrnO5uhBRAGMalGg1EAyL963tBHzs7xL47eHPUP0+r2EQ6f4cn
GgAyvxw5A0h4MOIwSimjXeKaCUSSSc/ITEc5x7sDQfXe5k46HHTPnIZBg7zs
q0fHS9JxqGrDhBfK0r0n5FeRWaeyWzADaGJVHdqjhWJ7UFijzE3vpP54ou/4
CrDWmP7K64uxvk7ldSC1SznFrHWEr+UyldsGq1mYcqFOe/TbxVtgnu9Mx1o+
HpGHJv+7KWFBsLo/nnAC+WE1C9j0hrIxPB8aawM2TOI3NXRvd6bfFfpNPS5A
kZYQ1PjkxenWc9s/GOXv6RV17lSOtGpPxni44CIe8tHC0T5oh15VU4EPQK57
3jN9+8zpjIvubV4r0lmv4ws7L4lE83t5a8kb9Touv5VgxkNqLh6dcMCl1fUl
J/evhWxJKa3B+U41oGvtpfip9xA735AUE2OkqdOWQVtLoADCsrSGVEAXzFB0
itLqwhU7FbtcunRI/Jeu5k5OWX8U2D4J8rhBQyoYJ9OtK3mQvkjWSoPYSYIA
BLRqLm0wuLBnWnPLh7qPY++vQSbjFxEAAJc9ZvHlL2LzWMK8xlf8zViixdTr
3mFmV8CygmubfslvJHMcKD5j5N74v8azfKKdsPMTijcQd2P3MiUmLBXfBzWP
4hKoxg1aaHkTdtKQr5JAI0BwjMlxEoIooTLI2++EkuEykjhUBOi2SeAjq9iI
3DoP6rjsXUhWBqMdmbnbtTkP73D2vsm0wtfjF75U5uebSvJjUHnJJ0KrIJI3
AjnU6L1h8ilj0r1YdMYqlVPlWyWR2b91aMXlGy7B6twnnKEXUBbhAO7mFR1T
S4fL3sPUBqV/GbpAVI1czKx7h3IuIpL8HI/OxJ5KCzHxygijBNitXUxIwYBs
47Eaq1vMfKjF0NhZLv0tK42/zKmI9N5vS2MU0gH5G0/uGcaFSFX5R3b655ZY
OgpppgzGYGIg1bfPTZi1z/i3jbF4Tx3lf0mABxEYkGxKVbUL9MKjgcciLBFJ
cFDmFrrhXcsZH4cJh+HNU0pgwDXEz8rpCyabaatCLzztS71hcz99wPWD9b1m
ldW1RWLJwXaYwwKscdZsJ4qd7Cu9Un3UDEj5dvftsnRTQyQ/99Ut0l1tFh+7
PLfyFJfUOP/5CP33jmUnYRbBayMUy2yUQofiJ806xLhr5BPWtRddaIfeK68t
ho+cFLS/3Pd7H6Mj2ezjrr/NPMNLBFNH0HDjMZ5G966XfU8EPFY5SSQt+usX
po8G4cZSvCpqQF/g+css1dHnENQQajbqCEIU2IMhlSf88B+KZFWrTFphVR2b
QwMZjhKRPDIuh2h2ZSSrgS3bqZrszu41J/yLCokQ1Qgsq+qXTBVs3KOfsleX
DTxt1YBpWBTCxah2iauy83s0dqTK+9D5YVPLT/3Lu6imzjfTMxIBhHvfC3sK
g5EyfuWsjdySrybqqcoEGq8jw29EqUVIHRBLlsBLwEYDxXMgMbuQSBGop9+I
O6Y8HI6xUoGX0bsXU3OUkciZkkjfcOqKq4zQdaI80xX8/5asIKkiv/HNDnmG
YsCev1bNYG/HYGlvNtwGqlI5GxLZTAD7yUR+xnzXQpYg2o0/AMmNxQ15addb
HxijS5Clqhnmx0o0x60ru82jXuzdJdXoeGmE7kfz1s5IVhenk8TAsSLEGZMS
8oD59E0MGwedszmKvkAkYj0xSdctSxj0BgJzpzxgbtQ62qD6yc8f6tbJP3lR
9ZewToQ4p5SnbJViwZC5Bk1vYhn090137NVvxL2SYQuqzKnmUUAe4XHbnC0e
EXHw8CmKyr+2/lURmkx34nfMOxgu5BwQeGW3GVd+ss5U6NWy4S6oqtXgC5rw
tr3uX+k6xRGCProm0np+a9mwBOYsAbi/Ksa9BcqZlPjtf97XE8X1p3t75x99
V0bwc8SrS5WFe310TLaIbwVR2aIbke47wuv1z9AGwUYEyq+blkWxuPA6klWA
1fKYgjsq+97VPXDHk37wBb0gHndl5cUHo5Pl/Po9GLFAkavDFMZcIiUKCelX
tEF40d7naOGkPTe99Ix3z5Ifsh2m8hVozUnAgl2Wq3NMFw8zbBiJLsywwuWF
xP+LvAInt9BSyIY/y0Iow80rvUY0FSwEnWAgKHeqGT/ZQy4jjWGjnWk33gpM
NeMfMK3X+Q5W1jyig7YlSt+bo6cQcPPRXe2UkUKPg7tk106cpjgIxRm6uLAd
JHss3ZjANez5ABA86E1F070tUDUUdzwUpFFHgUx2FMECuRP/ZJu72wvYcx4y
H3fxpsAJ3YGDCWLZOCsT3ghZ2pbL9XK/hLUA20BBHDmKQ9Y7SR2DqI/mrdog
DzPPK8zouKh75z2273Dq4SR+MoErow69RPXgZZVgdBVelrAMeJ7odtsGdUuh
YJJxlBoc6q89Nj/xoSWu0SXxSRoJXIG1Wi53tkOWXatS/EG8FraV6GjcdNcK
dM6jG+Q7Uo95/XfkqVLcrbHXjfNLYmDtBtmd9d+M2MNkKJwP3uYClZPLDL7J
uufCSB25xdSM3YmGYGew5ExNRBPHvXuYjglKb4dAG8oyxX0RE5hrt15U6wIf
aXhxYlB9vR5gihdZQkBzOgXnOiqg/341TKX9AOr/jn1GoS+83estTU0yJpo3
YyuyfB7pET5uzWOeB3hGo1TlKlzSNugQsqVx7XBCyBYuTBtDPQqqB7SAWacb
HuHA0cbcIwlUK1DDXaVG2KQbxoeTGAr1zsihmoed0OUExVcMx3dlZtYCAB8u
j+N6GZfXXtMd4hHL65/PwU7VM07L5PesiVTxY3P4ZXk/Fx11tMu6C/EmSvkK
enLLN8gRT9NDF6TA3REd318VfR2fhOcX1K46eTm33UKl4LgxlfrKzDiQtt8V
zaNJrETmXbQEf289RhfHGw8dKtT/00lCBy10OLk8+YhxAvgrGh09JS8hYgZ1
9F1zF3Lg4LZvEk842vBFDHaqesTAgacbN+IykipPEjhrReaUs6hW7a/riom1
5URxofH/0u6buvVJj5zFO2M1lOLO+EteaUSVEPQbyTYD7oF1H548Jk5+AwiZ
u4IMB4VjHwNzO2L3s3MxG3FEENPLU5Vhy6ConUU059tqYjDG/hG4OjQ2Qi72
FqieVT/KUcUU5zVY9NIA3CUDwdrEv25TgiscrbBqd4vBDrI1hsI6HdAM0dj3
K/GsCTIT68N1Iv0SE3gjbeMwYCU11bP4ttgU+72VmlPWQim2DrgiFFwhUkvk
U+enIpCAqYbExp959tcbjGDbb4ea+IfrNyWNOiwE86mSVJISXRGBSr5TDSzg
aRXBwJ6c1EgFoNcZMZwt57CybLgrTq8k88CoHt0cAIC1LMFSue3tViQOxdE3
cPCeBIXsH5pLWuuxGdoeE+Sd0mY/HaM3bFotFshK1RoVi6yq5o2O4bIt2VtZ
bKxCDtTnK5VQtUWTh7xE108bsPZ0xNRWMIGn90nPisUnSBLaguRoCTzlCLj/
qsxxJtQOWD6VnQoX5lXrvXHuSUG1ORgPl/Xqif0le9GD0AsGs99EXNS7RKYO
9vwEf4UEpyINGF8w2sxsTG7HatQN75/62z1RVLxAfxqdSlUEU6jliGXV4paF
zfXLSKcxB6ivxngxgrX/JxCrnmM+PeRg99fl8I0g8coroNZb6qxlcn7YOv/W
knLgcUqU6ELiLXCLu6G2b2gIx9Td5DQz1xZH0JDJXZPiO8sD2kXRSnwtlXtq
0iWwWANDl01LBAafNayfZhlHz+83CdpYB4s0UfysmebRkjMyQWCPTDzLvOu8
ZREbGMc1gt+GjrKRJ5XRKYg4xfMXIa9IcNHL+zWqM9/5p3EI0iCewj3lNrJL
F1xov6rcs6nDzsCjsCMizMOy/t/XDNSd0IbpGHPw7IXgHk0WJ6veSl/WRSA3
4n0RjdiYu74ZMc2nlFUkOmDUxVlWnnrGLnrgS29+4qXK+v0UagCk/oe1BmcC
PpXlrp97d4urhkkDqIXka0J/+6CUKb4puyJONNH5AS9mE05NcbvpQcrYeCh/
XvHBhD6LFcfmnfmQovk3slBdjvd05o+Xe5XIwGvyWNRTJ1dmyyH+cmel7HLE
ugN53BeaQWrvZuLol4VdQX3KmwFwq83Sf7iHM8rIb5cOyE1Gg4BkWhEOCcg7
jjavyOBppfbTQD5O/3trp6sNdtiSCAUe5jw9AtP0RSg5Sb4S0PXhi4yvlP73
MMrZYxhI2ozQ5GLMQRcfR2wsfIz7bMy4BdDcsBpG96iNBxCOoj8xA2R07Yk+
XHT1KDap/hBdxNYrEldpMTJELm8+o1yZI3dwklxoc3bzrQq+sLF5Rabk+Z2I
RjfmBqvIUU3dE+rsuLXkSI4QD4Tx6wWq3qkga/VTTysQ9+YFjtfbLErjQfAw
niTK6L9VOT4dL8Htop/Z7lBMl7H8uCfDlrLtsbwq+NXfS+3jOi4TZmaVO097
+z470bPgv2nsXpAZELpR0z2r/4nJfChRNzU45lkWCuZUR2nyrlV2ktJDb0uK
JeX9Fuj13NL8ICCURoUSrCNN+GxdAVSmeB/MISNbdEbFLKK0VKq9Gz3Af26V
Itv+glJPexVRe2I7nOeWrf2mgKAWe+KysY0oMFtMpo6kFKUoYefTYv5UzRcU
Pz+5G/6MmFxdrslj9UjMQ2EWagAwGeVodGz2OZWFgcws5F6fsG0/pAKTe8bc
OM6envffXiU3xFG9594wtcPkUiwlsd8J+lgPlG3BK+BTfUxyKv+FZlqy4jMX
TKxeNmQYKXxkWyUJXjzkpJWnnqM4cNddW31f1+ScZXsLAmCCuud4bq5M/f2U
wR416nvS65F1DAizyhxV0eGS4qAzugZyQVbTXCZWja+yzgNsbOg68FROwbub
M5ukAHY3f0xvQxGasydHROjLQ3d6AEcLTf3V+JpH+SFUTRzqzNuuiYNAS7S5
lmi22vHMjxEkkjfp/LpUzCO0e4/QyZBoHN5h7uhIPGhBnG11oEKI84HtN9sD
KI6fDcWAZ39EPmXJWHFDpMeaDb9z0GcvgpfJWQ8+SqPW32eh170lEr/kZc0z
S53X/KGqI0Bjqr46XwAzZ2JvM9cavITXfUJ7WGdK7U0EjFV+Me8YPUYpLkxX
3KygHo+2XhaIistT7m9skkYWDB6tQgmzS4K28//zDzzdzXg0/vdZ1iX/CiOw
IYS3XCkS3ndeg9Pp6U8Nzh8MhTkl2pdhoJh+ijy/EgNm9p0wMZAuQlJH0bWf
VXaU+pROa+8UW2o7+0goAwu6X8CWjn/OmQytMUnpFFeDju7tgJuxgwrfmb+H
2s+1Ylji9KnIY+uPoQQqmjb0nfSqThrJwJuPxRSX43AgjrT/K+4hdgPCJ/AS
oaYgD8iitE9PAk0/Q7r9+upJcPnzBOaGZ9dmaQ5jKxTAuAY622GtfWQUH3uD
sZyZn00bCw42cTib9l4c4eZDSFZbDunbNP0QVFLiPAFss9LtyJ8Y61fSFmOf
bvDfzTtZzi4KjdZvjQduvd6a8oHCa1lLL07LDK6X6RqMjzbdQIIS0dW6eOqa
VVgBZ26rl8pEj4MqCf5ybn+XPu766AJ63iFxQSUCfWURa877UvC/qoWUlTM/
5ueQ39KjMTc5ZzfnBa1neuSWAzUvxrfjYcn8rdzQDbvufNiHRYS+Szh9xLmV
h0hd2ChLpJwXf4kxYfFUf4NqnAljDgMvHcYhVd2BG8ZJ3JnsuRMchnnTLb/n
KTVqKNSrMZPR9FJSshTA69khlnsfwwXnxvJWH3zVBWg/5pJCbmqFuza9D9+j
XDdywTU9Gzau+4FIMrg9FQYmQbQj5cn47lIukCVdzbK8eAc5Kcxwa6RDsoGG
lhucUINLYUfOXk++FTUywEzFnEZ1oR2hDrNVsoPxMlh1h0Cz1kDiUrnK6HP+
QLsQVTLcXWqcB8igKX2UEkScQJncJ8BtePXjAbTgEBHxzbBoBjIDfcGnJKb5
kTtL86BCYb32iZyAE783iValv7OPQSc28dR2+XGLtQQm7M5RxrorwCQe0Ttg
NypDbPCUKJ7JXEchnEO9/KWcNc3OwEVLLz5U6jwE+J2NpD0jASw7F1/7MJWx
EKIJX0u+r/9FW8JlU5NYJcpvh4a+AfM4Y6gbHb+47oc+Hb2l027SVVVuy8hj
TOkuQXSrXQde7OJwA1ctJmYueTfK8vJMn1VYj4Z3jfTfQTDREsvmGqedXdnq
UH+ZbKwHwe2dvVTjTHWfPLvlRG0BPmv+9u7UB/ltDm/gndQasQeZMDBm5kJ4
bDN/FxYtp12BF3w8B35wWAjFBvqcdJIfPpqPk61k7sDSgydi72fe6II4JUwc
cK85dmPbkkbxVCYxUZolwGy3yq3Gaw9UNJ0wMCq/orze6j+mMfz+VGyG11FR
z2Emw3xLYGJlRJMPAXHSE09fAZ4SVIGq5Gv3XRuqy/8H4fX5zlFLwy6CuIPd
LGIt18Dmy18f8SpjHIrjidsTYF1mW1ZGOjD/KT7vDFeo/IrCMFRSxgFdLJHJ
S4uVnCBYRceDBZfm0x0uTL6Jl0/XnAptGzJ7YljDoDIZjBE/oDrGXnYQr4Xp
Nn8dqluKgyq2JvQxUFNn1GCMWqg2zgEb4Q3KfntDH0pR0MGdY0AHz+UARaiM
fRYnZ6pLrp+ZCNk2cwhPTNNY4lWCUy8ibK1/fPGvfgtnBEpgqORHgQDoEL1L
8TJNyoMsI4w5RIlECU5VV0JPSDpzMPHRb/j3KbZjhKi+uRsD4VCg2kKLNore
nwaMVPEdD/uoLwqn8pLP+wTs1sqZPoFWulc89hUAOx0FC4opjPoWyH4RbVFZ
sZ2mMzzQ2EoHgm03hCzELFOTubksTP/xVm8UzArbMJKE3geq/TyyRKaNn+eE
XDmV1B6uFv6cgRvTt54IxBaGchiNCnIvUPYh3A4yNLa34MFbuHjpIw3YagYM
2hksD/7m8fbX0N1hXbnnqVzvqOVaLzNuOz4KBz7kU42af+q91QSMD/SXpFAZ
jEGn5FyDgCEGUC+L5paHkvv+mh5b2sKgIpoX718CZ7lzPJWGfnnU4/GA5YMW
TuUbc1TeotBtsWooNVUOGT9Vnz+vSk/pKeW1Q4naq85xVDpGcjE0xTyVa24p
l2DQXTcrSiy8lNHOx0rwrxKCmTPPAPcAvu2eQKEaLM8uhJ7ITtsqX+rkCQJs
6WrriDmAQty9s7NxPHnI6Qt1EGDN2u2qLH3WzDAQc9JQSmAOehZNBRIXG/sE
/W9f5TYi8lzq4rm+o/W6TSWC41EoN1IgwPWY2CbNCvDyNZdHEuBpfvWLPsXI
gbtbkNJ6lBammRcoKbsNBii09D/zMHJh+W8JZ/WT71+kHlsMSi5umxZAE83f
clNqEB96OFf4yHI+ABAn19B8fP0D/yFqd9f8l41wOIbRZ0YxfFnN2y2BHQUf
RvXoTz7RXGnlWR42/xXsBrMsRO++LylhhfBWO+VGCClUakCgPZVyGltQr4yh
mFe9zGi+Qdztlo99z2ncSsyCV8lR7UeTbtgoWcFIWcuXlDPDF66vqPGQyAKc
G+/xcm4NsaxXF6Ycp+MobA2D0X8ft+zVYBr6cjYS2CSR2rgJ/rH7DETa7uQf
DhewOV8G4zRMpc+vmA1rmuW6kbQiaQPzILNQ6SuX+XYB5Va60R/qb+vn6a78
2AJaQJNloMxEZpwV6Vj8j/WkZOue8aq6rZGVffGnbv9YNJ4mpIonQSJ9go3b
RxvRKVkeYs5mtSVCjlnJZuv21ZlJBtANeYnnx9x9IMqG8Y5w0EIWHS7ZDOXT
7OkrwQ5CLniV10aKduVFO+W/url73jwwkugf2CmYjeAfWIylgHg1jLmHCFa3
8emneSYodnoTAxx2K1GRTjBNmnplWh1/F9d2L6/qI48lAuN8VyecbhRW6v8w
M+zNmNoeNJYIRbGb9Wv43ezvupDMUJt7BgZBvq42XVNC2ox7yrcyHHV/XFm5
67qWoBQqb4BlJs3D19rjCigKfY8ICJxxwa4szhdAYaTAL3UYo+kUO7ZuLrZh
fvlgz6HsD9cxbBSo5FKGsVmLMdQWxzwdk6bKurzXXEHjdue7AiU7IZMRbRFS
ALGm4Js+Gsv2hc63iM7TKV8SVsT9ASNbhK2tIHySUVhkzIKADfodcbiStFNm
c+qFQkWDK/T0Wg4t5tdzqSfEo8FJkbV+zntjedZadpyvvohHhotvhdZ0T5pe
203DEZna76mKgNebxEGC8KUD2CWJgEQT7aYx/HADDmGrKRrmTOi7DAkq5kDM
1OOVJgLzimI3Is7Xhp7bzb2nZ8RAPfLEP++/lflkqJGKirHgyWikumFcIC/N
HGZJkc9Yqv9+MXRQcwlhaFYvU2HbNeH0c2/J+b9K+2lMJUJwNFgdfN7gx/oq
+GPpdQiqtssDODp+YQBav6EdvqVpYDL1RN/HEUt1XYBjl67NDdTZ1+2zCzOK
d3htLcCJpEqbBD7DOsLk93spqUXAEFZSg8oWfJcP9uW/7agRr4YVIgl+aKnC
PR1PjN7m2C3PDsWFRQqEvy0Aw8F3U1AIagQi5vVK4jmpAiVU64h9oVoh0kTZ
xJV582EI6ue1wOtT1LPQW13ZlzGy3bW+5gq01iiFosxo6whOdHCwhSCI85Ux
Wcq3E7by9wgXZK1uFX5/SCFKzGxkuhVFolYNVLSMj3NcLhHeGh5tjZXFBNV/
XUS2YC8qHSiTP7pKAnbYVa3o4GGwzQndQP9R9oDj3SZ/RLS8hJVp5A92JcLL
PeKI1cnfZyfTN2oajxWLV9p/iA/K+CEPi+IKvvcBM1H5xbB9qlDBftaTDNtQ
eRoAdWLwfisU64pyu0d8jZB9hW6r73EUEmA7vOGjvNAz5pUlM8Sz6jBxrbSv
vJIrEEyIsjzmsRFLA8fv1iVfBYbL3TeMzbxcgaSuIRkcNn8/kUZKy3Mj7b5M
G+Ck7838CTFIveXQ5VssQtrR+D1BcD7WZlRDE3pq1xs7BxJ2A4y+pRHq+Ka2
x9JP2sOgHnEpcKJMsgYWjRy2dpyQGz0L5qQujkPXRmEFFdRu9e3EHA48ag9l
hXcyjRcX05vUVag4MIlsfdpBlwt+3l8P1FSS7PFRqdGwqH3q2Fgtdu21VbXa
GgPWHqD5cQkiOlgq+Zmlgf+MNc6u1+RjvGe2LfNY1LFBlQPuxqfS3xJULG4W
Y9nhehIHP+sDQUPSDIUGV9RUKtiBpUOFPXBhst64G1ulHYBFLvVkota1SY8x
6loFVCefyzIesqtr1XCVrXmyjU3hzXOGUPTd05CHHlqV4HWVUTRwMt4NF9Dy
mrPalxgr1YPHBQ9bM6U1pFGu6JAlRdKQnKNwV77HsyDwykvPceijmLFg9XNp
MbGP1A2pLpFoZux7qvryyl+7gHVIy6jr85A48gx2DKRhDAABTg5Nnh/vr4vy
91mYNF+zj3Mn1290lH9ZbwivDIcCp2R/d72SwCcXaRSNt5LcGB51pvyR3J8I
iw22VRWeyEUpzyD9fcBIRIsBVMkH3CLaCtOrR+gj3L5rJ9QwqV3x6vbVdH4x
bnt9PWm0K69md+TQftoIl6pUu1joXZ0KRkjCyA4E/xqVdCKMOgR+mTqBlLCw
z7a56vKwZ5UIXWb5l6KUqQWHY/FpXpmxprhzyw4pXzbf3mjtgJCjDwX/LQS3
YlTckq++pqj/f3skIFttWrw6zhbCUYyrAKu14MSJRlBV6iYMtLeMhn8LRnFC
TQLDNhnKLCZLS28WECLpsaJrxB+02hfy+r8QTg+z33gverGCEJFedB4tPFU2
tKM6njk4Z2Jc+9aKoiS3NOq/S/cweorPisJXzg6YOOjAvzXaEzqVoIkhP+oO
b/AvwYs2ZHx5cP15YT43CRLzmA4DoPN1yvBFYk3hMvt6ciBGWf2DuN/VDytN
W/2tlMwPY+nIKv1v3kj0j6NvfKv0LfYqo2BS5oo8DYnk6qUy93RngnqJpbjY
/9fH/xySFa3hufAfFEPBha+9khzbdUBcZhqH9PYZgoOKyWvQaEA8tGmhXvzz
ACZlSXFWOBIJLmJhaZvg05Q7WcVXskydAuZ2vazMkSHdux/3w0OZzZj2OmFu
YUIKu90mW+koanxQQX21AAqek63fqYweMFsW4F8s1BS9VK3BC5t/ohdHB80G
N7T8j2sYyeKq0/7DOTA9UB0gbPc3GbCidaKHCYComHvz6uR51OsGfVwGgXTe
Fhmm+F9Rg5SpVGf9BCj/it4YPptJnxqeHAp2Oub52WCqJQWHp9lwzINhzngy
rwIG/Or1p5YzbqetCzkk7eXJu27Eu4IgdLXfBc1XdbbagHO1HSvA8YumXqFn
Ow9QrrSyzHSpALhSPs+SbgiwFqOZGCGfyWWtsOl6opdkG3uVvifsMLCVnjag
YpoKqDMsGhYS1YauJSMfTcAu5kRaPaBOSG9g9PQDlRuSP9jAt4AyXa3cX+V+
xonAFA36ojJfpKRDxu/zY3lRo9haRNFi+ihMdDOh9gy+C3mo7HtmPufOCN65
m/UYFy82rNCy0vkv5/YnZ8KC3zuJMiO2FLRy0WcuZlDxHoEW+H77cEJwzq0P
qk2D2kNTARGOEXeWETYcBEamC0lJ3tIq99mjToSyPseaLATcgRCjt1hnTKmS
zpfky/qLKg49zZp2hzrqWIhkWio6XkTR4cngpLym1FDzkC4Ty0qdihheznzL
j/50uIRyPxX/WNXEcYMmcMN0hK/k8O7gN5kZOQsQ847B7ILSl6M7DD8YSO0k
QqIG+Izu+3sW280pWWUJSya50Wfz3yY0WTm7TXctvbyQ1WLzi/qoQoyxg3XQ
9WDuXh/3w02uhE/0Cb1u/2db7ICAeWyVBvgS7MNqi3LFNTyZKjxQRYrzPNEr
NQsnkHmZrffxIvsVr/hjiB2mcqPYAdtCPu7FgWFSYgV9bzdHeNT+CvySFE5E
Y54yCVK2h/5+eSpv/Q1NHGZ3GS13xsMkk5dPnsrdcXj+B6uErNN192XZArsV
t25bOlIuA24nzUZ0HLiC+JziHi13MlvZDapf6IaxET6/b9Sr+r/cgFrUvPru
3KOQ0e0880333Edjzq/NUM2DvndKPsCaOl5TcH7+bwjVRW1DsUqh2sDqmODi
hxAN05svneBqCHumzZHUHi7gG4MQOxcLfVPD7b+mSYz7z3l8lVXz1FH3ZnKw
u4bvCqZBhARK6jmjVYxVsE2VQRvRePW/UuMqabBKSB3U5WE7NaV9nxhxI2W9
qsgfXwHz8/pl49mrHdzuoyJZRiinU5tjoE2kH9+gZpC1heP12/tLpV9vAvrE
cw0LYvnJGYKe5mQBF8aZA0CE4FScphzB0KNx4LINgG5EWoPKCfXjzRYUd2o4
UJhIXDruG1WYr/2wbLtezV1Xjmarcw1ZT2ZgrJ6X8qwba1z8M/V1MO+9nP7u
rwcaPzNdwR7UFLQFwG2YKLb/N8qex9WJla2QqbaEc5RJUee5S98z8460SqGW
HIPQmf0xqo22kszGxTjfYQ6xOZS5iWBewObBWI3UxIo5lehpzRnx/2IO1UUc
4HP+sGbs8C8LA2EwAhZafJkWaEi2gi/5i/mKoJt+69vz0UtbwOatUQgfgSir
ajrGyPDoJwtp32T3LEcllS3WzTO1w89YWkjV2PA15ujwy5jAbwQ8sxo/72s9
kDfD9Sert/KVXAEjoWRg36U2jPpso/nTR0nqr0C+efC7MuxZQmgkGByJW9Su
gM3L9BCYZ2hlg0vl83AsmJcUvQuKKALDf9M9HZgH8FBMXv/maAZYhbupPvWI
I5n31tZEQleIXwoKHGNWfjh3IJXhi0f1qh/AdJfpvJPT77eGI+WXEu2vaXKo
CEkpaYTbSV6W9IM5lCIFy9ikUzXIc+0kAmNTm4OxGUK+l8eDyO9scHxqprCN
mFymD9oOiOzDg9qzLXgROfF9DDOScQO8LEy3WDStcY7xgQufRq3/47jd052Z
07ZJwEXih+hpb9s8+QRlH2aW5HrU+RO5XDNO9EqXDV6ptl6NG4753WOkK1hl
6uSqM/fvML3cnaXa9EIAMgFGuqBy6ARtcLo2A/bHwsMkf6Fv0KZejKA9/BDS
a3rOc2fqMm9NwyDF1FFVAhS83GK7Uy6Czhc4ro/m86AVaR9H+R2bPRGrbPsT
9GrLrZtC6JZ+GTAAi1pJiX3TkxXGaExfZzxqDa1+C/sXXjZGeqeJCt2ik+If
FQUZkyccmOPwgR/6XJ4XrUlS2rwYA8JheZUE8aLOewA7g/AHa3PNcoW0rawZ
svFEjYqbjspgN54nWZCoLAxYEjCcQljDHEkv/nFVCKQuahhRFwkVk+hPW9kX
E1KKFLrhgauTnBzTvtlyC4nNDm5u2bxh/3upL/P22Xl5DV7D/P543mKznLXY
KpiR1UWmHAUZbtLoM8auAybwebhIQ4QVQ9sbX3BHFJCFr2Nx/fQrj2dMjGQz
woSEBpaCoNZ4dUHjaFtj1J/KTIc6kjoQndYxyOdxa2P+tsgRgCVTxrrhkTL1
nBQwW6eyOnU0y4cG1wsZ1YoSJbB+9ndHxBX6xHpqL9b53vEFR/zumGaQ1veM
d9i1rC0RIr1al7/k6TEU6CYLupINMB/oUyJ1jVoHwNakEHU+4NU5uyerCUCt
/LjUGb2DzzVGO1Ssl8SKIOYhARi85R5KVqNImoa4tyv9lqlDtRoaAc2lKg0h
nZ4uNSpkepuBMha244InzH6DuJ0B/RECtfsidOcbtPu7t0Yw2gn86loxyni1
eNWJ+Byf6QeaLR7nZCip+br2/vDiwvHss4QEr6fZjF6mZO9xhFMyptOg9oc/
cZS0ZRJSVksJHbUP1U0mNPWjxHS95M3Vd//5oXE2gXJwMmN+BRLF2AX0oY3k
4tBWQsLU98JHhsm1bJRw/KkFxx30HLj0GjtAf9nwXP3hNXpOrlNcSAJYZ9Gt
AjNGjkk94Xl3SPBbJnzBgy+9LTw1/arOwA3sPKKbBxEtc2PVXv2INLx5QfAG
9ca6BrHLqGjBDzqsSZR/eQwyS0g8qtREMA4OfjzPmGFj/dpeNGr3uA7UKX1O
0PR0muQgWApILhX6sA9py59NozxanSERlFycJMJnAZwIJiXwDPomnx0dGJje
ROK69utgIHpoHCcwl9kpjxEMCLEh5vaVcss8wr+ZU6vFm9EfBIptqoRXuWuc
84QdFxshsdZBKuRmR+l460yGOJ+ZEZRqWjGOPZcFQUQAP51PP05WjHzebeiz
Iv0I5mP+GFaO71iDBuAjdOLqq6WlVQtZWbR01TFUvxZxZdE2auCFyI5g+KFt
WuKIgAwfuspsohANhl4Ejf99FP6/hO7q3HR7edbvVaKLCOPSCC4RDt7soj75
1Qa146zQoaoCItSviJvOcWLkKpo3fD+uo5GEiVGCyjvLd2VEKvDI6dywADD9
Ivnuy3hgX/6p+a9kluw2rdKzjZlMgxHbTs380bw7Xewd27pjf5Oz+muyGBAt
wpUsDf3CiZRAXYE62sIwPaG2qdbjU+x58rCVKX78QXnvcztP7IT1E5jX6BUE
BleY2hNJxIp1s8k6HRdmhC3cid6B1+CJMGeenQxPzz+gP1Ti9URoDBNDG7UQ
XaF0efjfcDpYq7ZPH0nYnIjjT0/zYjT47EvhcYv512Lpr4LfEVVWn35rq3V0
jqIlvMWHQRHc+ckUj+/pqdsq3tQKdVbyGRR12/tSsaEIlkVAM43LXvVWutRf
1agtMwcqnXjAPDg6fbOr4t1oyorgLUnwcWqdB8jzOrsxo65GD24uxykBBRHA
w6D02wq6+praWTuLCn+DJ/S+o4zYKI0ooIG1JnqL23dZ9Nu0RS7QLW1y/Aum
q9xtuQVr1cNhQ8vlygGjzXCQY4Fid77ojZJRtI9XrqK3wEmQfar2+BhY4tsN
z6yGazTNLnf/SFFXMEc/WHKNheuIqYsbgGl6q6YXp8kDqRCs/EtJAf067r3S
r1ToTwYHFBTgNbLSxne9InnZ4WpxmHBTTGFxdfAYdpZSGW/Sl6S2GeSKQ/S+
/v8tbVfheJ9eNxHTreh2HmdNVaHOBz3uwsDA9uVYAjYQhN13Uk5M2mtaW/Ey
CAUfHQWXYTasCVEOPFSwTVijutOEaTnLn4RnhPoLm+h4kqVQIFd8rnF4YrpZ
eFu706tUZj0TAENcRWERNqQdpemg0/5dM74aPf+rKz1FeQ+BY2Tebt4OIrhJ
B5Uc/VbBCUe+awTCEoiUzeKOhXkvFI47UtfC5fhH0cmRU5JIVg9hzQLfhY2u
FRVwYBuqNCjiGSCFXBrVF2uZisgWGDYDJjrHG53VL/ZbP2JccwW7toqSVrm6
Y7sfNPi5oCEjHBFNfSbcI3jm33nuy5+uRV2sTor8q/00THcLF8j4bmXZMi5+
wb8E6IGH13egTuDhVL74ukK4oemq/tyFRwLXHNP8wmJ6FDp9+MY9IWkzRMR5
CBRYXuTFYMnCtz6pLo5VC7rMJcA1D3m7oiX9fdBHI7/UX40tLRoz54oMBUct
Lbi2dZMu447tIrOsGUUHTM1f5jB039JUS9YO5B+GDbf4dBPuoPz0IRad/dQA
+SXcNpleKS4Nm8hrNCGp/O/WuZkepV12GsHcskswnucFq1bzUw4CmKJVNZjr
La9cyzlAdjmBa/jyOZ0Bb/HbYjPW9aVdES/aKA6so7b8Y8WchlQDyAdQpPpt
UmUhOaWUDxdM+lPQO8L1hN8gsR3MOyszVzNoNMZdJTZEVCNR/YGafxFaFKVG
MlQ/ioVGAdJ0fUWtgnKkEXVVPjupts1ie2QMG2NRxZaEJqyt7SSWUIXpP1bg
45TgwTucbEZfS7eDo4wmEPWkUBuecuR8QMM3Mt/HBL/zW6C0em8241CL+o7P
mxP0UTDaRxbhNjTTMX0wBeQpqDvcmRNStt5Gy5eB6ObNviy0Dz1y54o7g2Y7
rUw4xoAQcmvFIAhkyNDA2zPua4cRSs8OqGl1z6tBlr/hYWv8/TFdmXaCww7n
bjhkZQGM4O/M5uJNwsetOKHcZJ/nJz4eInFn1r7EsbhkQDA67unojKP+yBJ6
8BKnoWc7t6tuBRG6zjkUUOIpWcdax8yolkNLDrXwkLz5oi5gI8yQGGjIbQdA
RcMg/fYPUUX/Bbu3thqTy24wTe0ITzZnv2zfBlVOfKKrrekechhkyvVWlMRK
m3SE6Or+GuzAASHVANN6lyVYr/OBC3SfS4epINfQZn3hsLrAw+2vbn7Ymi1O
UABPC1aMpzFMTyY7frYd5sCjcARdMVJBRFk2xej1NVy6g3pWpcsy5uRqEX24
4//eG6YzyYxSeSks4e+2JLqwznrMx3mSYEE8MqQ23NrynbOH1hn6zdKrVwRa
DXSMstJacBswZ/NlSivv1q0U8r9X5hZi8wYvZ1i5oNWi8Cw4Z4f8OjkDEy0r
K6EZynKH2b/XzvUXb/fUCX9/PkmYWuaKDfZlv9m/znVMmsxVlEgONYAZmM/v
IaOLfdDdVAmmdbJ5uaoZuULl8Z9HL45POAtR5Tm54ptRJ8duSv9fVokRDhr8
NnVKoy6WYCgAJg+3YaJvhtjVreHp0lu9mzjkEL87/b9PjDPUix61H6T0hCyb
hGjDrZFzUGCs/jX8h101OpFzFsJIzdQUG646f5qi5XUX9sxSkCAVrP1Qayw6
TyXlrnZsFsmstt1KFY3F345+qg2XGgnVFHLqh04pkhqG1dP32IaKLqxd9FCw
mtAxCQhGRCOMYJoi5RJWnqy7jY9if5GVqapSs5PwYf3nzi+Q2bls9PccHWS5
D6MihXG+RWFG3JrsOD82+38DW9+Y1Y1W9h6IJdvdVHIMZp25X8FTOb2rTDYN
yn2xoF5FJxIhxwlcE/MNx2i0R9ismHfD0r6yVSQSc0lt3VBr+HCZAZ2lL4p1
RbfZRWVYdgVLQydMTGtf4/wCavS30QjpIDF21iIPUH9gMVyH3BzateXKPCRF
8VIjLaGjJvNhyPtTZfsc/6+gcvzXGOMmbMowqm2PrTRuzJS64CW8BCPv2k8d
1e8wTmjH8RN2+7HCdbCwasMgNAGAHjkF+ne01YpAkLdcUSTVXGgDaLwDelVl
NXTmWajxbfG97KNCRDseH9RPitAYNdtj1VC2mi2Ta/nSXTcn5MHKk5Ngjbby
jctg8Uaely6ilJWjUsQwYdU3LhcFCooFYt/U7nIMBSGAgQvIGXj6PRRktTuY
0QFv4YOCJueU8bV4C/bRWRsyQgZDcPauvchbGHju547sVmAHwOdbyBQwccNn
Dqvdj0Hhdw1kyCSKQkD0ubIEPi5CvkOrD+YXNSLS5ykpp0gyvmgnaaIu3sM/
3vUwVZNeY95kcMfE8sARSWzlwP9MHpOcoZB089TXwMWbdINcVfQQA8HkuRII
rl3RfelHo/1Sy8avM8GjXbjx9Em1LQ4dyhJtrDqZUbefu3kriPZxYxb5Cp4O
AQzGTu6ZjlFjkaG5MMCPeF5Cegl4T88NCkuLcypp1vdREfRu5720Eu9w6lzu
MkGtr5e+RXPHcvhiqQS/FxdO1nG1wk0Mz11fYBnlW6IYL5Ptyw285r8j64cJ
0AgpVPDSbQMWQWt+hjpk7C8L4K919qAzGt9H0fG/pR7dNbhl7WFHRg9ydj9q
zIlcgSeMl1y7idwldM4EdA+eOS5QyguVmsMtvrk14kmG/t+nAr1haZkz/FJX
qG3v06v/CLdIIS6v1CP2D4Bp+SJvEk+mWD4LO02vEGpLGlSA/K50uxX1XiK+
56Zxr50ihEs+3RJV+0/r0T+cElbvkFehcW13ktxwqIHBzZ1ttyspTsujUC8J
DY+A8MtMQq40tmt6nKWiypsCoXnp+VcgEf8W2H0ehoQ2Ucti7Czt03L5obCR
3k45698YNILLhbNkQKFhsjCAH9SdW0wWvMV5MR4yKJPuR0LChQ+9aLswND6R
NvQuFtuqgPBWwjy1x5GC3u8wmxVKwDhaSHTCPOktaHVtL2MF+XQrQ0A6h7HL
vTP1sEgoWArplzvGTeHrfAXIumkHWEFCHPjEP1a8Q8HVAqoTv55lXIpa/F2x
XWb+FkP0K7+ycRBkK3cpIfNfHlKomlF0mejJziExib++3dBjw0zxPGJ8WqXA
NZDeMheZ4EQfQMjkbj42V/342XIRA1UlzFa+pmPKarOL0El7tdcUgXKbQbc3
9MHFvbrzhML7cM5JN8HDPZV+I9erefEkK05Yrl2eq/6jotewzDuULF/B0haO
rLXih8qsYvjAbnCayNMJzG54EBMXAvlmnzgPqzY+YMpJSz2Fmodc+37ugYji
14YNht1f9RPyCZ2faZEcustuy/Fe/mPiK/vksyTyTobx7x82zNuAYKwicxX+
xtnjFH8DGO78eVpFa5KRnfJM3mIF3AI/0I6FDA0voRe0OZ3Th/0foBtGTebU
ixXuOFiawr5pAVhDEG11LQOQJfJYX3BupBLANUSp5Ivt/IAIEyw5lFWeeEN7
rvCf3wS631ClfpAI/XH3vquBdMC+0Cmvg4TbrG0I/mWFlPmVkAAmSAl3gWAx
OdgddPYI4JFiHj/K5DV3ozV9JCzgG8zCHYRV8qN3r0t6p68BVxDFsohiRhS0
9TRlUurpEA5m1+m5L6WwPTR9NAqmI3dirJ5ZCE0vPAU+hwBdq3+rHajis47+
Nf5kfonw3RUg268mLP781JXO/RvomNzPOlkf1c49lG/TPheJy5XIcpZ9C/VK
ohrLFFonOsbjq5Jf38Y7yfgp1OJYlKcyhIPjdbJkeDb5JsRV1wC5skMy8cEy
7fiQGyp3di+IHa1kyDA+hLmLsfGvWWJGf90YKHw67osghkY75kUZ5jbYkzOK
wI6GUyD8UID8BM4faVDgFfwzZgavhGNcWq+OZk4kO7r6MrRwZxiopq3Eh6or
p/LzGd84LorbrZuLnv8dNcxDL9W3mWQmtytXCSSfxXEI4x5J4na+3Mafp0eB
oUMFZxbZeRP0JrBSVpib4YwWWdJVLiRC/KkDZZXjQwUuHsmxO5x25LczNkMh
dxrf1yJs48GZkQorNuEdD7Ixte/3XKozV8rl7s9gL4I6RkA11rgJrEwMVttC
Klx6fhcjb8C8x9PCD0ac+udu7AeSgGsLQpSwxUFHLny8pqn/PSEv8vJYwPtM
1cu5qCNJ1ruogomNN/cfI0EYB9D8LccjVqAxEy2OgLihMkTuzrxP/JfhTfDu
XI91j2i9M+OpfQdpFYLobelhusMkM0n+i2rS7yL2Kh3j1QDIBfI6j9gZtxcm
2e44niEq4VeqTU6CohXtjlxaDTcSjtjyTw7n4llL3hUjZgcKvXtkntGjGCNU
i1Om53lMbxoK6VJi6pz8YpdvhBP+6SOyk3vu8amxU9wpaWzAk5Jc35sJLciR
vHCXNpKPSBhRkZacEGJO3cW4+EBUFfhAytZNn93HuwDIJ7QjCZjrQPXyIoeW
nkG9V/2UVz/BT/bXfjaZlFzkQtTpz3W1rH51ykIMRu6I/Ou97PNYlT8BOoGI
5ZANE+wnxP48t1wSZgLTK3OOeBReIFyd413+VTsoXaUCuHaGhUqTjGCrTBwp
uKfmSoBHiZsLlHn/8BVY6J10oqishPbATR3clJhRZd732iiR7VO5pFh6A6vp
nypSe1mTkBgMcY48JHdf4P1oG9sKZPBK/3h+vztbwLcn4X2jANfAH2gWvJdm
DobtC+zE9FoLYCMpmqb+zu9CWRDbADro1oW2uUGJrut7hedErozteYF1OI1I
8SE4o5wj+WbR5fzRuinyWIeGvAwOykomZtSABxeS+sQAI4VUZBMDApPT1PB6
ZcFjqjzYlecxV7KpABvOBj/2PPjjF+vu1O8m/jxo0d5+/FJdiBRJGJePHaDN
+3jCO5DjmycNrnFMHYVT7bTOLAIKJ14yETvWSRAzyKtr4AoO/ZG0rX7OcgrD
LAI/DwYpj8i3+EnuwXu1rKr1is6bW6NF2CBSNwAKNDGaOxdBOrH3r3eNNhXl
eEoO9nvlW58AOKozZHuNEmK/hyewJAvzK3O3BYyHqpn+DMC5V8CsGMHhwg6x
o7lTrg//Rpheu+un/NP8D1JvATC0dbGC8uXRz9sC6dJ+mQvzvc2LM2KqFvaM
NyxGjyoLjsAB5MRdYLMIoneKnVy7Ra1dauW8YksID7dKN0B0Ky6prAXWaH3G
EgtUKwxZbTcrpUs7fsefnMkS4Cm3tEpXI1xnlsaiJF2YxaxfZeMM4G/Umi5o
fxKSmaOJpISY3Lc3Bap4YzkkW2A4mGH0gw6gh92qrs/l9ZhCrzwdjsUI8lxG
lMnm1gKzaCqJxpNf6VEpTjhENCqoRC6hfjmukBK1o5HvQiukkwML4BiH3SwI
c9xA8AwZnkZzSPhkmV1hfgaqfb8Pcn26P8GtGPmfkL3AcwwBZdmgUBL4pCyG
x0YKDT+eeo8yKd3CHCBNXuongiF4vNBX0OpXHjgK8X5BV8qTzo7PzNCgDwD3
cw4SS6NUohH1Qm+YCY6ZyXEp/pk2VjOv4Fq7NyWqdotpmxU6gNcr/QeFm7W0
HEGsLGoWSLbt/P2oHHp2qWZHO+SpY3jX1c7vYRE7utfBwJ4gTQGMii0i9eAt
UPr7AfNNxtX5owJkFpwTzEH+yL27B9P0EciOATvv7pgFwaK2B06tuba/G/BK
fU6ckFEJgr/mabduQjyxec4FYyCt6n6+gzNXmfJZ0QxE9vvVyPMrYWyw5VH6
aobOeMzQw2BfHvK0SRELHT99Cfin8wyzlaAg4HzF7rGAugnoqXCztzF8DY4r
Ea8JPskowV5mmz20aKUgsr6oRntPHu4P1l4MZnwy8UOtYRgB6ruvuJMM08fe
XkRMny3wSM+/4upube6c0V3lLimFQUN7VrOu9BvNCx3YVg5mLA5qHS5XJv3x
FF7NfwYLDTEKYInthK4a7fsi6/+lEuppyfqtkjj7jeZ0hW3hiZjXX5IYwQVT
w1/gHyWWVmArE0zE0EH8Oewdn6sMBrf+A03Mt95ebBD2GQZMof1FAyj0yeAC
gep8t+gU9T+sWHd/rJg2DgE1CBIMnsLW+n0s7PTWuV2Fa0Uuecy4FifgBv3q
MIeigoJcpOrhpQxuaxYmZfCm+jEXNsgt8XhVbMQNWxJgdSlE1vnPBjGMI9eD
E2GIzI5V8mXi807PAPygq1PRCiPLun89gINGMsqjxnrPHJ23eqDJyXMwpjXM
u9ehZbwrMvmqbxnyLB0v0S7JXxsSGI1F+QQ/h7EhB9+pSnmwn7O+R8OIYxlw
W8A5APY68cY+zMucOmYPwu+jwTp9D7lq+Dvd+/hA6BiY/knAjoLWA0Y14BNN
WW4AtgtWE98WdbotvRkdSQmvKsEmIjYq8RWLa3geAPNEukRaUB5p1jE2zZvo
neZS8+NtNbuDfKDFCwn+ZIOk3QFj2b0rgqgclkNzCvpyHMVgGNW8pRxnC8nl
z3gL0bGW9CH1fssBKltLlBrWp3nIKKFWR6b53P8bfp5Gx0+uw4u1ag5IoNNO
Sv+xwR0hUDwWcXzuhWl7qgZkeL02aIGwac+PW4Cc7yhx99Hwl9wwVu92/h7D
QciPRBp88Oy1nDqI0OZEt5A+mT2O2StC9DnJ5eonzzscAn9f9nzi3o02AGnB
kPZYJOztQWomNEm+jKWGvP0N2E+9JP2dmdegqAVrbJyQysaumqi83Wb+eZ6J
NR7g3RSaEYD6EMPW9DgJG88v3WxiNAFmvWHMXHlKIN0DvR9cV8b7Yar5WTOM
mC4zJ9dnfNDI0FT82q2ueisJhIB0cJKGK7d/SONvhhFGFNYM0/F6msd4k/yY
K8lpdjYXrZDVvcWQsLyfTbCPiQvWisiodknrUYRZoSeAlTTrkInMaqjpXZep
YYxcnOGLWfIk1/UF1rpT/B8h3E0k2G31tCOYnIp3QPvWxsZutN75toSRGnFj
eew0CogOOLNaapoX7SIaQ+FMvK1NXaoZo1/BVbcFYeDJrZB2nSoUQgBkIyaC
7I2JZ4/t2NndDIOxxGyi7jP+C+qPNQuAD4UyLBRLiBLVtmB0LjJKHX6RIuyg
jbBF//PytlYt4xbgKnpifOZQLpxl9hE4dwELEbQPc6kXlo2heItyXTwneCrt
i9JOaDdMb82/zhwaIQsl47co2NZ3lYtnaDBzJta/oN3aRa/APJUnuhBhSVN8
+ph0Og7+XndvOCia6vzu4x7Tvd1LcZOH5nsr7y/J9KmZkTsoMa+aRCIGPGId
H+TYvkdgzts1+R1VsKXS4psu6F5wTz0m1LHgNniGJuvzRYl6ZiJGsdyMTRmk
kyZnnOVAZdIRpai3ipmjbRaBqzqIwykw3JGM5H0IgRYGAWFjKR9nxZMhaUyt
/OeBR63/QEpwNuWwJ3a5dNHpUMbA8EcvT6rrcxZB+n8GhKpoMcjvRhq24tJV
NNokoIFE//39iw2OCeuMZCaRfjoyWimJASYLpmokI3DC8bgjQ5xZm0ntIJ1x
W43cwewn1rLCmz6is5jFpXwojL5/FLlRfOGnx8qGveh7ZxdnzU2DDbbDOBcV
sXNADq2JJeLQ5Uy4ZmTqSPVuLpy9WgrWeGy4gspIKamrXAgjoPYRU7WUURZI
d2MDAtLohWmmsrmxK4svVTd2W+2+FAqZ6gySzWU2eu8uwII87OjbiV+8Tkgn
mDsjQZE/pleMfhEvo3ap4IRoEUxzVrieTjdfAv1Sm21WCF44YAvN+0GMK4lm
VZvfiCCYiT/PG7wnaPooTKstJ6ql+6hqb5dpHl/WVb4kAKtbjsjI01KnjV2g
tIMpG/axB1Ad8awF0ApI68rc5RYGQpfAkJpBRY8Qh3OrAQdZ4JjcEWcKpBI7
3FZTPFcrQBGJRxiZZ4BmbxD6lQLtvyM/qZIw3gNNcvs5QSsmF5aakV12xFr7
bOU+FBIpC7MKen+TAZbHdf7Yn67lfJoLD3Ccb9z/YgQRfRkCyFihTwJ+6jI+
COJYszc8AIQe+MB5Ub0jhS71EPq6pZX1D+NHuSWleh0FW8P7KCv95oH71S9S
luv93B6iHOB+hco5wWFFXf1bJcbiIeJeILR6k/pzgjHBkRan/Xh1XWk9Gs+7
PWJ16q4p5lk4B2ODX8Uh0mIDZZCzo5ePz40nppsbl/+Nucf71EVitDD+d+rM
nzXf/gADpPqkZapUqdEWV6PTYNrgM366M9i03ttAZiP0pZDhCTVxzg6G6G8a
gfET2+c9W/tOBQhlWvYHOz4ycm4S0rVK7BlierKUWu3skpI3WFNI3ipWIYhS
ddQdAaxyl7c6ej6Ojqq7NQeOFgK9jzd7qySFkS3LTE6liPiDMOjoQ3dtjJ7D
NrdNq+NtmsnF78p1xV4vr2jF6PrcPu/Uk3t3Ax1H1xEDXUsTTmiyt0woMdgJ
t6DBFt3peSRCXdLDQSVB6+q4jlCQKHknFjYWiLzuJe74DM8ZNu27dLZvxa/v
eeQRPoCP7FW4nA4r2tb0bTyuKu7NvNFPsC1pmlBtHOTAksqxuwHJyV0ANJT6
deU7kryy03LafZpjCnkjyox1wgjlJCc703Ff7JdUHsx8srOFo4OI+tRDzd0O
VXTUUHtmPG+GifMIG4ydbOtOsBIFa9KZs4cFzr2ZNgBs2waWzAAQUpl9vN3X
0K/tlI2hxwQFviJsnQm3ztArZCHHaCRcXZhom7GqaPKWwyMasbEzvLePjQNf
v0XCDsY1nvkrY3mia0EVBCWUs/XPixL/6Nnin0SVgZvAdiGbPtsUKF649VUf
+mmED1SsUkELlF7Ws0zfHcwukWkxCJxe+v7GR3QMposf0k+FN1NSt3xPJ6IO
EciPX+39n3tPjTga0u14djYmXFfFquV2NZwNSf0HAY7JKAPlMBj/YmzrZpsF
Cy4E5kmMuIBGQPNRzk5xGncR1AyxzHzjCj9RfB5fwieihSne1UDfKnQEj0vm
ECXuEZjh5dW3zlr69WcvQpTzXm8qAzNVxC6UYec1vRGX83zUUBTnQ2rIh4nG
b648BByJI0jExffWSTmVz7Rzn7tx051dWSHg6/KBXN7LSDIVugqj75LdvcxB
MpNFZOLIq2gsXFLpuyEdTlpNPJSVgJCF9S/l1zi9JUhxZcxExEXm5KcecGys
OzFB8q7X1c1COClBu8BRcmvS545X/Dxzf/HNC1oX/rPl12K+e/rqK80A0pMV
gWF7mtWy5mZb1x13u6j6ZNmQskTrfeWjLXKOiPz6FDAZOWWQAdJl2d1rVVhr
T5Xz3+lMXt26IeGcy6x3M2JywmlkgCmCmiZfWYKw9QmB8xQK3BBvCoFGb6Lk
tPdfUEWAfFfpUYmKYYtRgK91lfmyjlzhQOetOgWgUS403XAN4V6s1MgO8dPd
e035EYz17a+Wp2BMlNeX5cVJ5mUThIsiaAkTaDbx+sBzyE9/uVA6sNGH9UO8
CguFUBIg2DcKOiW7NeQAbsr2/SYV6nTeOtLdYb9L/yrqRSQVoYfXwXfW0Rxz
aTEAU7kMRZa5dU1eBjwpx0GS8OTPc6PzfzQOwHAGyzY0yvP/Q3k/Ri8w2jP7
aKPAxP38gM+iazka6210MEAUoez9H2tVDMfscBBiPj2/xmmVTW7DoKRr/opA
OLmESQAh+4prdpqogYfEYQzhGHkoyrSbiYGHqINE6PeH2Hk1THivXpKkYdgD
dHoaTP/Z+XZDq6TmkUH6kuIJTWsU4WNPAIo3MAl9T6XJP442dNLO//UjNYmp
CSEXs44AvjkO1zXvB2YZQSOjqtIWjRMBAasdoWAajzHkB8t7ZJdyWQYY59Ya
WrTTFPB6fax6hyVyZxc5b/HrlRfQFc9RHGv+kSs+56qRIMD7m9BBfEpLm0W9
5l0WvQTACo/SWmhKxVSCbpArPlV1TwCMnKUxLD3laVimmmAdVOqn6fE0clxX
vgUfEHFCwF+3WBtNw+BquprMBZFTLkP0qGVH3f9Cl/VBgpIyjNWMndHxg1Fo
qSZ6Nbc1pwYkmZmUPEY25XP5jOdchGti3lpFGCBC8qTPc0xeZRzll/SHbela
f2uAM6uolJCGkeUX5rGNzN7ywh2B9uFwsjj1Qtp+Y8nuu4iHG48gwh6Y2Fbw
/nw4jlAGdsYq/gnqVrxFU715I1KJEhZkF3eRZyYSZnBGqFW9dpcDaiUWdGbU
YTqZTNXjb0FLybECf6IWOOag7DH35DPwwtKRtWdw6Q77tyOa2YHg0Lh1pPQx
dkhz2WxDhLaIG+Mtj7Etv0mAfSRLoKjqNPtITJyxiOuPR8FAd2IXy+p9nJfn
azrloNtWWWfK+F/1ph8eIg6wNzsPgh+LK49ejIKOfuXYhGTXx9ULeYbTaFQU
wkq+bVzhuT4j8B6rHiLyRzA+qF81WK67t/DAKc9A1NOqyoIPJmyEpUPpuOSu
vWeE/57Ebr4KdJWEBIY1t7fjWki6Mau/AUYdqlyyx9tsExM08Rga+vnHa9+N
Uwkw5vE92d8ANbOKHTW2lU4atJeXcUbZZEQ9Mww5O0F2C/zhNZBj0K51ojTo
qw8y0BvTzO56HYSGMQhbmtZTnqYqfTTzABpG9/gJXWh+rlo7CnMEJZ5FxYWY
j0G49HCF328Hu6ixFMXY5mqOpYbElP32LAlh45eNoFN+IrojM4bmD5yaTC6x
BDtHWzJ/0jABWbwh/XqoEiDsISZJS9Zhr3op5f4GdlLSkiIIh1sw5ifspB8W
2UEAEaPy3djugLOfDNkYQNtygInJYKSKdTfoeN3CHM3JLDBbwrasasqRm8L+
q3H73uqAtiyQJxxWp6oRM6bZ77yqAPIpjXmIhdBEod+Gq9E7qZdto9FO4pvW
wxN4wRNQYuHF3jGpRnMhohsynnXZLZs2+Bpsl01gPy3KdxNvKIjiYUS4K5JD
PTW12bR/SPiVZlNDV8sJ+GW4wKOlcsY3uIOC+KGhSEG9SfZO7/14PjHQgBaA
IEfNDqx5LfX54Oy3gee4rZ6AWFeVm5F5WS13J7eCTyoL8PK1iNjUs2Jxm2eL
NghHNxAxmUkXGw8aKCvkxXnPCHauWp5b2KC2RKkJc1cw5JaBmXaIDPGZRIef
abag1P6Q3a5Ls+pXFGbdsmEW2Fe1AJbm991E2iFopVg2mwUgQYOat1VGc7nj
DzfPugRMz6BmgDeaLjWER9rwB3m2EqIqKLmuZ1Ql0stSmpUOYhuSqDg95rHe
W+USQDL/GIM4ASCQk2XyweR7jVcPgSd+AIts7SyOzT2FTVtnh7QS5LIzhaWM
/1TwPdpylGfp2nnoQs7HhdHhIdsx9/r7YCuRNGV8mKejRi1UnJJo67vWy6zn
5MhCnRK9c9LdHWAUZi7s0O2qrp2MX9BXRpf6mzmoGgwi7Jiv5sJ+p16L/sSS
K74qU5It1LFtS8qzQkCzOvSsUp5S+WIfjoOC97CCM1AYApgwv6kjJWKOk+z3
ct5xQzHQA+TXpBZmdCFkfGrCIV7BumOgBELi636mlk6eyx6WrhySG0yq7ha9
oynoVjSbV/2vxNDtcFi73z1PKZhRtweTY2S09/EsQ0OpLHJjNlSsxnsLIgKi
a49GTDDf0Ue5ZZtDmLSt+vNacu7B4b5ANx5zP6ZlKKUSY9vxNlsGwfvoc2y8
VwFR6QlX+vJMPoXh3DSHOFJgPsEowCwBz7BTl8bUdA05pji/DTlIgtCPpih6
J6+qotd60JpMUTcWiDgeFtD91+MTf6fUo71vFrVS9XeZAfx8EmKUKeuchb2l
G1vGxQJyz5XZO5HlqY6WzXzG1Y+K+6a5J06xJ4dwc7LRqHtxvLW0zPDYxbjk
MZiTwoNFlbKP5XrEAA6ulhUPi8aKHxzvjt+2C+owOameVHXSmLTfV8FCeXM5
ht8M/T3BIlBfU2CpxdGnnZ106IPtdWxJKaneth74UYfs8Dx1gTs+9T2F0Whi
VpMokZbAsoRR9tYUbRP4Ns3Uv+NUdykdR83eTJ1f7y8X9k8V9yl3MMorB93m
uIqR4BRnkFpKwTsshv5RkYT/O62N8FLtljnRuPRwlBah2n7K4wgoxz0RKcxV
LME7KQ93CmedOxNPhBfBNg94JKbDIHlO1mpfG0u5b7tLr6jiJEu/q3XiNasE
HG+ROWom3Gonxo1Tqe4Ts6WIAtHMfnvy96yus6MXTSQCnIRMlDx1g6UlGnBJ
LB9XSmgwFq+3/gqKEhVwP56u5ABehDHKnGTQOMOvNrBgDMActOEzkZzUTTvQ
8rrbomXIAlIxRBIryQOYGcpRKAK3k4rwqznk89gfuYzQyxkGYpm7H+/M24JI
qelIjCEm+wQjulI7+y7NXFw6cyedjD/YsgBDDXH81sx3SIl3/vpn/WtyioXs
o1Movrm4jlSAF0hoLfYrMHqWh+/dFbsP4UBCe44xIl4eaBbZ0XDkJwAtTkg9
J9fqW0QN2xC3hfuv82fjOwC4Im70xi1Qohx8zhzM/tsP1RVpsgudP2q8IfFd
wb3Tjdyn/i2x/wxllFOaA3V30rl/fGtj8QTTQ95mcixWPxNnE75yw/t7+BpZ
4QWoGnupSpv052RSOKQeU5/uVnS5ifZGTVdAnpaviZSlz15QknIxXjlrHRkP
NziL9y49fRURZWW2f23G99srkr1oVYK8SOWIVgyFJRUB3xb9Y1SFEKqBPg2p
sPviYC1qoSujBvGwUg2f3f8XN+p5a27epXGgr6kvE442DheIHzUOe+n5HXF8
K9XwC/oDUK7FXEn3AATF0t2g3UKGB+6ayemfeep0uYgxWqy6p6pysKk6gb8V
H2zCQ0D+HVBrSWq4zAoYl/JkVOgMkYFZc2B5AE1U9RuATcHwQywbJggEZ9Bl
1yv42s7dKs/TxSgr9+FiP9EqPyVvFPCtfz98KVeVKgVQdrlg1XKcvRB0bbQS
DaSq2ajDASS3Bn9bBVXHyqa9nkTszb5G++G8bwupSmuIJF+tYFrYdNarkKJq
ml078WPRK47aO827ddrfVsaVVWYf6ndv5LfvyTkGWslK2AU7ppuvpAEtMOBi
91o9BlqDSNKi+a71ZEWnK9uhHLjUc3Btp50B1C12SnOBr+QndeiyC4znO53F
u/0HZ5SixqkSH2EZeqBUBkVbh1Y7pVHRjgNQPXlEjz6qP79MO1U6wVgtrCj1
q/hAmUB3ltBKEv9IZsQC2RG2BYdeevq/AK/YWpEKYzK5dLToB7MkwQ+j7Eyj
IW454/pbHKrT3KJ4rLfdWsdglKfIoXcJHl2q6JqE1Zi0+RRSnboaMwRoIIS9
BqHZ2YdFyzbUVJ5JDmD0GqHJrkAZccMPa8zNYx/gSfwuLcNKFAhW2xfUsmS+
Q/DBXb92Z+1t3Tamu7o9KUS8+7a4zPKsVaGs4a7cZ5Br0OkkV5eNlhxZh4zz
zbJdbaCes/RKoPxE1hgFG5mUG/B+7oPCBSJIXLMqO92yze7xZLT2YWK4smqO
4zn/YoaMLAS+91lHF0sJuaGJ+/QAv4To3IhhBWEh6LlZ1Pwo20olwaxrz+2J
5HGPzxqATRIqTB0ZCGYIptQlwroDmlimFkyMMti8FbFB5MyUmR3ofgEp+lwf
F76LO/SUMdpbppupgIZ7234TAaAyNG43HVbXwtB7a/mSNYViyjK/PUOmU1Re
u4FGcUXxVsovGJYRjzHmEY8bwTiM5rzP8E+jHxNerJ277CBjWQH6VIprJWD2
xKNZfdZbiezwnea/cc8ETwRtRkyKPDrO5N1wkcbhWvYw7PvzFGWYeXLswWzD
pUMhy1ZuI378+YL1x5qE8GqUU35zS4nhMwLclabeM9ettiQl6IRCwQYVG7xW
hKgk2ooEg4Q7JO1DP/1q0WlO0JljQdZb09CmJvbHpIRu88zpEJ+veoNxTV8Z
a31bRzrsnBl486arjzgCbZO5BmlZowtlWT9KowM6lF7E1su5OjexcYwOQgKL
I/Zi6cV6i8tfI+HuLoBaGva/4fZDPvsf6J6lBEdKdjFoCJP6fV+9uHezaIYg
CgxS9PAD8ytuXdE+OsjvYQ3RzmewEGyAMVRA7OMIdiamX3TtwZJd1nF8cf4N
dlQVqYsjVbGV/VxZkgezsEV+WF6PsXcWQi/izmw4+Vo2w+XOgbgEYVfd1zPY
AYPC2GtC6C1zaz79kIgn49eE28sqjQQznIIMqq6Dc554NsJDkUQuX/fMR1T6
NGWNLuO3CWBpv5ewm4xAjrx5B7OPLJPg5i5B6aKsljGDuTBzyJgReixjPPn+
6PFaEajgNxb5s4dZhmhFRf7AVwW1o0q8446zGm15AS0nTePBd8HmdZFlAEzp
nAKPCWVeackanwy5evaQ/aAGdoKjPUlp7Ozol8QNpJeiN1UJDSn9cBd9qfwb
JmS9w9duYlQVlialXejUkPzTttRDVZ3if//z7hDv0XjpchDEX+kp1OAK50KP
sGvCxZVC4cq/3ortdrF2Y3u+aOkpF9t35trExNk9SU6xoSW+6j3svjv+ETq+
tmjrVZdFbAhupZ7JZl4jP6d5NAjsj9vhuiJ3OUhx3NANck30BCHDvhBfvscC
sI8Evt0mCmhO5iCTGvpgPwPetqwARuaD6EcSIPe4SpnG+HoyjWmZDlVTCk0+
Mog4ezyMlNrfE6ral6Merqz1WqKH2IW6Ov8TEqwORUJy4t9KDoQ4sNueY87Q
NN2SFgR8t84UoexioJyrr++PSB1fKdLU5dhVP+LaaDvO5p4QrQVpM9G1CmPf
1CtVVZOS/t4OZLobZRtgSlC+IYT42KrVQF7vHamtrTgTBjrZidX/irQzAkyT
uzyBOSppkjr7dN6SRf6UchHu+w6J1yCgQ73Pk5Kxw5CybAx1MpU4DJpljrdU
RxBc7vi5dUHM3orFXp744wNDQQuLxNLlVTQo6e4Fnt9mO54YIU2uQDF1AA6P
jVjfLbIsMfxFLpj7WBW8Jb2SmyrwuGXUj9PJJ05yK3EHfKCQfyRU0QyXO/8r
sOIqlyxwpBb9REOVfCXuwLK2xU2sNJvZai936d/K23+j3VOrk8XWxGGwGVC6
hd8ETeh7YHL++bChlTvbbhLSLCIf1vVUbL6WIehSfMHQRDOF3SkmsZWXonBT
d2ZeVkhaAUTPrPRWYQcTX3yju+eiM95/1S0acsEzY2GCV7xcMNVVR0QopGg0
J1YZSn4pJFFPP+N/z393/s1/D3g+SI0HKBNZmqyZuURGqo+Ea6diLm2V4eMK
1xpwrXGMPrF8AXluflaI2EVqogQ9euS3l+soL+GdVOPhXimBiqQw76Wgtx+O
gj0ju29szSnjUkD5/K1k4u5pTI38RXBVVUF/g/00MHASGM2oZslVI9RBJBx0
hUFmxuaKpilnJetTjIrAqGp6IZgtJs/hrmYg2GK5AbtOqF8nQCXuotKlQ4f8
mupOQpAUdqWjGGMSFUAYkae2hwGea+LgVZJ84J5TY4xUdXafqQCtJbe5VHdA
r5tWPaqrRcB6S5B6o4r4CDTQPU21CP5N9IMwbUtcQNo/oJkhrwmP6Ud5Qj4q
NfhgrikPu463R3Y92T89W5/A6j3pZQptwcD4ikl/ENHNrt4A2kR3f7ZMaG+F
hnb7aQdSqt1WYksLUCF1ksJLrYDgLDToApZhfh1+ZGKCOKL+78NC4+nWROIz
szC1qhbBJ54zz+fwkzYQwDyF9OutWIBjPUuQtfhe0dtIf77VSPJjzNfm/vme
4Ak7vkDWwLYh+/ntbVXizUd/dvWT2xywXqEErHlBljFfprKwyR+I5gzI/WvH
pUKxgvHTPY80sk+uecWTcrVp4tcNplqb6sEulzBSEfYBXlPr/tYFBgB8OgYg
ltNrfiqcsHH7VdqghSfltXCgd/ch7IhV6hLPE2vCoeEPZImyhNQdQ9tz2yFI
w701dNar/ZVxpKjri/sehMGLw7eR6wDTIhTgA84vqZ3LAxN7zE9ZJGbhBd/g
NRXOj0p7OGXrByfvGOwhEgNfX3+bHlybKNR7C6Hjc9vkXiaiODaYn4YAcS63
o7VjamrN7Jfi3WIB5sA5f46zqjd0jzB3i33LtEkAQGRWTZTmKzERtrEAqYb2
9CDqIiYfVrOcAxdGf1/t0opO1g/2KIEeFuI1QDs/InOzMD4GzSnoOkQZ39Xg
qnwOXM6CfODZJeehdgiDRX/B3N8437mghY6KLO/IEg+x8JHvZBXzwcfAnTCm
10ZKKqcJDp0va5OnBuVHYz0bjg/rhq741Lt/pwcNh4MBHzvwHXZ5cALMx1jh
in5yf1Acfj+NRTJAK1+MDI2FoWYmVxkc7u2V7moKuLb1DkpswL2LtmfgMmYB
JeN3h3/upXdXwmJ0ZZ8V9907LuRtmQj5PjkA4ASbd2PN4Z6Nx/3MKzcSGHqR
zds0LAuRQ6fSaynFmQUdihHVtvVH7hThbWk/upBa6VDjiq/RLt+LHEH3zQ/Z
CGPB1amz1/lsDgC1P3FKkpPq6y1fLtaywuIF37K5bzuDhhWZuAE2fK6CgdHq
51gXig806oy4lL9v13tPXGWpoiTLgL+YjwXDThnEbENiPubGSwN6RbxSEv1w
0x+Z6cxbscInRf0fr8gVZlw7LJzxTn1EixM+szIwzsRxZiUgAKvtsFZZT6sQ
wrqA/Xuuwsqo5pzIsMFO1E4REME/fjr9Mm2eVNOqP4X39ew63l4DlZZfBnZp
mSR7DG3c0OGOVFiORTbd6CSS7HJ+UXGJKKDSEZJg6+eZYrsQwnMLfX085WUB
GGJCLxPih39+XHLTGSkck4+p+v7P3eubEMZOKJUYc3wrCrk2Rpn0JgghMmVz
fM96Um3NClDf0HW15yUVPwXCHXfA8HSX30Q0mJwriQu0rqV8d9Ww+Z/JEAxy
eo9Qrd8rQDVuHvC4l/u6CEwc/uhivnlKLx0hN8udMNJSNbfqFXtpzR5QS7LQ
ob2Y432hGt3vv+4Qlk0UjC8CAkmWkvsnGu9GJQuT0KlpDpykuozZep1P7/oI
0rLiqiDj6U6D2KbMPNv/hkJPF0/LIxMZxfDit+mTjeuBi+0A9KG1jzat+xLf
ngQEuv97cB9fUZuQP7KBE5r2fZ7BGLsTtuyw1rJkpFZxhtX3uKV/BerPqtKk
hEGw5Q4W47JOVIqRStfzt+nCo/kXVrG5cJejpX5CaS26Zv9Ka56ZnT3f7n3K
k7t8bWHaeMH6V1EtcgeS5wXGsU5/Dbgc16j6nsiqJbvWijW/8YgyYcEaL1oh
q5M76eGDfB05qeDQ6Eof9o1zDiEfEN4/GCWsQ8tGlx/O68YkbxUsVJkhhDLb
skILjR3z1SMeBKageGKFJsvxjlUpfrkIRzrMTVz6RkuxuutbKJYtK2OIRG0D
7s8x8XrgawZfWi1uUc69eusBdDZH/aXs5LY+pvPnT+v27KdbpgiK3cvmEqT7
4G7tTzPlKr2cxwJmZpRqCSHPctxDiRz9ncSoVympC6mPfz53apSrikRF/lTY
9y+yF2770yPc2Qlk5wMp2ebRBetLG8RIlweL2gDsI6N9DgInyXfqeOi7zW91
9lmgFnEZFtBmwb5k6270jpMdnTRfGpYfpNCwqRqnrWygvGWa/g6d388RelYt
Udeb5J/Bqi9uhcrO6926buU8sVl9KlhoIGFDHIRj6RZ4HsxWlQNDaJtd8OPb
Bu1u9ljzOip3z0npGmieiIGuHtnEGDP+kIZj5Fs82VIJcZepdd5czaaLn/yO
i/NdB4Um3MM2SE3xYJieEZjupyk3VKLxTIib36EfX+5YykXG5jQy6A2soklD
tdSyv5dwchr/5gtrzFPF0P6BxzpfYFJLjbj49GlwJLQxsapFyZj/Tg8D+cAc
tCsfjDBdPPxZaKWbCEB/UXKlIp7+3AwSam+AKYVH/FGT9lGRVJGMpkY5T5On
VgFMNOXKxYm+XpjHBzsfNc6pJTtU8L3wuYcr0QopENxGnZoMVmkZi01dsP5y
IIkKOMXPd9m5IUqmt62LtFlBSxho2UK3+xyMYAr53jFOw81v9MT2gSlW5jr8
MCl3t5/aehGb2xEZtjeski/auFfJnLYDyhuzS/rsu7IhLUmgAKkb7RJC31GP
JbuZCrc5whcp/nifdDBbKpNUPHKZNFAZALacmh5rgC6buC+Wwj43XJPZ66Ey
bKenaxa61dZRWT+hJ1K+gbukyv/eGAavDV0GiMtLDWx839lIn62KMpNBaYba
6mqzr+eMNEG6L6dI0S8SfW8fg5MyI60UncMFpSqulMCAiq5SLtgX8WgyfM1f
wC2bveaUobv+aAuLgzUjpwS497HhkiZ877CqJPw1T0eA5FTRHCBleFqLVUsN
8gO3+r94aWv55m7vphgBl2HBidB0usv61wLlCc+w3qqkzKb5VBjs0zkQXVC/
jgYWH9xur1ox8xIiTjkH+aIxxJCKN8LMo6/KQeG3i0LYWNmnCrMTBp4Piuqb
XyVLyKSgDG5wLMzHtyTOVeo7We/fsUZ5pGSNmgWLqiY7I3Z0IzGD59rV7E0k
suNTMBqlZ4GeFCuuoMP3aXQOcoCbsLc4loe/4LWEHYLpWofL9Z0cn5DZfBQ/
ksr6no+uhUHOz3Kqf4BmaX56FjX3LQqdK2aV1wop39PmK8mrmvEzv+05AZ54
J0j3+RuSXy/EV9i5TLc8Za0I8yMFyqsKgdwiIBpmUHyY00Z6s9l4HQuhNpIK
hXnOfkYDOL7RUc0pTx3tuii4bIsUSs0rAt/rfs/kFc6GLf1PPk9h+6IXrPel
N/Q+3EF4p0cFV9GR1zDRQzf9+GDmrr5cH5Rkkai5FF/FjmRSmXGlnsXfAq3f
rr8DdZDmBJWhO/uaeJMEe8y02Lblo8u7//QwTOm7at61Ah7jHhmuzj0qB+jq
oGUluaO4gSrw9a+Dc+EjZpW+DvhfGA8Tc787iWZ38DLtl4bIbpQ1Sj+6DYIs
JG7BUdXRXjDFfiGVBLjMcmF02o1amCVy2NnqYZHRz1jxidKnvLM7TMXCkl/z
RsecT+p5ut9VKL8jNHvW/y1Yv8zOd1ygtv9mdox0cqz8OU1LJp31oEG3DOXp
lF2UYrUeMqNeIJOeX5DGKPWbm1jhopfwV3+TdN5gHT5l9tUxLSomUa1uCcdG
XZCvBG3pfYiYcaZNWZuTMiDDpztGOqLr1xJZt7hB7T0iww+UWH/zHB5g1biB
+YbGsUofz+Uy3SW9ugzUUkFtV3BxKyDPXPUirNdxEYLZOamVFIUhOqudG4xX
OyGMOUP6b/OOyDb3SIihUkhhz11LyvkYkLHhxnqpzau83hqAx4Zqy9RGsV38
4fMQoaybqL1+ovIwY8h+PapLtlMFXbpXoyTQkOF5be7E/Nf7DVGrm2ENmA0g
w6TKEzrJEMXtb8HTOLMP0cYzRLJJ88At+mdRu8qafDeApkXCKf4C8Ay0iXMw
ZrAUiuz+KNT7NDNzqrEz01G+/PqOBgl2MJc0k0fmWLDq9R/VnmqpcBMw7GSQ
UMBJP4+eSGLvjAGvLfTzx5CR2zrj08nK0yqcK+K5XHIHbU+ivt3oyRPMJT5N
0wYhen9Yu6rRpQomkUR5/1TJjLeVcgSdUEj9bh3Yqik2Wm0iwSUYvVM7sMj3
PJCZFJngsBqunooYHbwMRSfHS3ptIv19nnQWpxrG+UFKOEcr+DwJJ18ycGRu
kW1C+uQYXbAUu7LJZzvZdR3VYZp5u4lzeyPKgLwPJOvy2lEy95aTDT4PgLRU
UIxg0gRr9aEAkNXeUK47LJUsNEGJUtETHDMPwIfTeGJHnjpeXyIPxaSSnvl5
vzI97/gZxGUM59Fg2uoD8l9BfB0xaluCbuuVMdtDDWwyf4crP+fG5UUSJ7f+
Mmf8HIfgc3UB7LXzX3hAb0pyvxxl1tfghNCjIRBB398Do1CtnQnmiQAEk/qJ
qQ5Im4M8QMK5MJ2QINueJhQ/Xn7C9WUq8ci0Ib4PgntWRtv8n6wXdGZ6/rTy
Vtj30xTxTDSaGsTQFmXdfnaRJ56VmR8qRXFIvhOFWnn7s5GkkUj0y08GdBCn
mwOdfMJYQr3SgPSRVsYj8zHZX83pGSt1UGdouz9omUl8GZrutW0IkitsE2HD
bi1HK0jX6NOhXo1+ohE+/A6vzNrIeN+brXdfMCBkpp5ieER8B1Z97gg4VqLD
EIap5rOalD6y9oQHXKgeDyIZsRIy+MxjnDLRbZxXBmO3m9rK6clvG3RPyW8X
HgC8EHZIpk1PxHfMha2b+a4k1VqM6JNubIA11wfvPnuKd2QfGJhOAa8GKzwZ
pJY05MrdmkKbbJd7K/rhAX6UHcG7q4KtOg/HjttMbXHP7pR3T6vNf7iF/nwQ
VIcmSGpFyGf3iOpQKa23l33VRftFr5iwa5amHOyjt+0d/UBN/FP2aRmSs9VI
sLXocLzOyX5taJKuEtbHA8PptNDz5FLxJBIZ2jP/dAvsldMd8iVSDCmBJn1K
GWMEg4CmSvOsVqFD2SroIiA3NwTrKy+tYSxQNFmM02VyE3LXQvwWp2tGtmhG
g1C2qRUJaweNHM7Lnut/zFSSPY23fNtKC1TZl5ly2W52147h4HvXWXzD1tsa
iE3iUMo+TExNpJ8/ODz+xKgrCT9xebDOn88GOShD8JaSr3LF0/P74YnzuJxQ
H8x1Vbie6SGw8ni/WfVsGAh7xmRTvyZWXi53GZYE592CjN1NTkGkrphgpg8h
3WtrdzBUBAoDYS5rAxZtXgAfmEmFJhfJoN22DWSjns3Mwi93alNgdiEYfnCZ
s/1hpJfoepwi/ogEUGf1pczicYvYRnnaMPrOKevzite6BKpv8kW+a9KvIjJN
3JfNMtqsnWQe4nOuVfc6T2/gyRYqJ5Vc2vSqJez1iQUhxzhFttW39pYjWQ0R
00tt9o1dh/zCpTgEWzddOIJgaX99DgXzSJBXLSFnOf6xHI7I6eIuBo8WQWAG
y3rvRbDelUG9ajnVY3cg4Gq2qIx49TNEVXW0gH0kP0nsBk4znSqTcmJ25KVe
GXpbub1xKv5Sm9JZBDoVRW1aeoJnieY6y3iEVMqRcFbzr17Oti6X1BnMcfEr
wN4R8mZ0KUWtGYUuZdsG6LoPDHopuni8Hst91FSkJdjl2FHQvQfoGlhbnPHq
3oPtt5L7VvH12VQpo7GV1yGSpn4MblspBOFMkm1tTPrI4TOGKI4FqA4TYwsa
cEfa13cjiDOpyLvhoQ3GLJtBZ2xPbkT2dxZk+ArwctLXBaoXBqeNRoldiJsx
5F6vkjk51M/QLfBXPGtU43OrDV5X9D979HBxJ9BDy8/PJUW5iLUxU7pcGLIs
Ct2Zy5d7CTaqBxPwdmJK50YYWkyNtCwgi7Ys9mSumjgZRC5+NLYbMI+bMJTh
Pj1bLfJE9BTEn7B/BR8sUk38OQdiVP3UBRbffCio+HB7ulCZuxYR83Jf1Ush
3jREZngLdCgla5bSb/CfJ0KR1+pllJ8u9NlCTOqh/BlJ3w54IiIuQx4mKyzR
RozH1CSwsNHfAhjO+wVC4LJzcBfZ5sfWG3k51/oBXRf85fG0KYx9D1pQbiPZ
Hp2V10lIJTUOrxXxhJQY2FbokJ3SQpQEwtYA5mwrk5UvgBwJkyvZxy8ppApI
Mlw4E6HiSzBXdS9iE8Wi61P4t2VXW8oyfKBqgDaIE63ySCxpBM6y/Y7ciMdk
8V9HNYKxDW2Pm/r+TtjAzgkfObJXAL2NYYjwKwEPuXDNiMLV1yl8mzBVLd+y
rPaEhQ8xu9RmsekHbAiEJ4C7afX7L1HJ9sZzF4Mus8C/WIybbiX2J7lO4Dy2
5mIFFZLuJWswhB4wIykKjMWXih36chTt1YI2rXzSUbDzUMVAweDaqbbrbpbs
hjWUXUIMa8EXWyFm5LKyR0pzSnDdk4k/r4+E7qFa6/C7Trb8QRYSkyYNk5e+
dqYbiwiTdFaSkdNQGDZrudqMXHQ4J2SkBJL3iUqwHaJW89qetM2D1oXWU55M
th7H488+L+A30+ugytZDdVg4DXEYXzkprg53EwBuQ/Ue/Sc9r23Yb50Gitbg
dYi5Np0cOXm0FsjgI8z3N/QTdlZC33FXx3n7mpLRQk20csi2Fo56+s2RrFQP
15jsqNUccJr2hhWph5x4L8JTcH+YlWRaABWq+Nw1rn4RIGhLHElSNefvYr4c
A8koTCwLJiBNFGD9oBuaQMjr2uDGOrgqZUZ/1m3vQj3enWTripNC8Y0sWP6V
EFwCfNhPRl6QLrJMJnShdMz4KNWvfLucD89tjBe5akU2w91yTzoC3q42jGRK
LWHDiXW87zVDsoy1fKHIH8jfSkQi7nGZhUEHAFH8IiN3BvEiM7wDuVZ2o1Vl
G2WBBPbSJSuGQrQVgrusaCVKMdPCzGu3fyfmHoXCgUcOZ1g6t3STIpKCJrLp
4Q/KU2qhhd5ZqeXVXsUO62OTm4upcq+VCvZN5tE5XZsHBiGaJZcbKypzsKIT
YS5904HxCDTvPMwR4dUkXeRV9LdF6kMYvZlsLYwuCt2O/L6IIZblaBXMrsuY
Y2wQLzvg3LHfh5XdZ+DIzhOBKpJxHdOGw8woUw8zcMtoGMxvaWVBO20ZMahZ
7Uerugz4lACp8/TgicYwIovMWPrBYZcnnS5u+DTyj/lcPzH1+vKQBd4jIFUF
ImVXtYr3HgmR1zDujOd7p2Eei8losAjuOr9sSWWGyFoGCUM2Af1qgYuzW8VD
GmSkJu/khWnPV3zJQsgOaynyYNWR889FFZX6LlfssSnYeS9ixTdxL57kcbso
5spR1kpGr1lh96I7CUWetz7treph4orhMaQ7lcUFV/3i3ViVIEIOPIE55yAK
fLC+DWp/84w0jtsJ1SY1uPrqO7NqR6vWjBKZr003OhDOEPRHluvV/L1df/6d
7PgzZhb1G+qFCbNv190qOu0czgsHHMFXdz1LHQ/PWnldb/J8MKoWXMwIW6JN
HhdJwSltuho5WE3cEvX1WXv2lDgQC51mHafooOjSnes7Sy1p0g1eGT8r33tP
hTHzLKGL2njLrg5KIqweA/F8i8RZfiJGGc1MGRUvYT0lNCj8NtGJyQ9KCyK9
w9Bge0ovWpyRqOXj0d+RABs4/goATYLDl68SSew7M/KS+fJdEPWEi31IGyoc
v0Yq0mK6zeSXe+P42cD8hO20/zHcGO12d7v1rGiLGEi3UMcnEADPcsWv6+Bj
QhMit8kBi/Ngt+qCoPLakn3dCaDcMMHNKpvq8P57SeI9bhhZn6EZ/EoEF8qN
wYR37koXAMCI7I8/vkySfX/yU/N0z1VlojHgBB7AxXkodPjFwO/Uf9EasbHQ
YVi798OtTTbC7nccNK0oqXGaITpG2wToK1AQS/S5BLveUD2RL2xcWG4RmMUs
4KsBtzZspz3STUPRWHiCUc1jLxDZrTSDxFK+hjxRAfG9i13CcfaAVlSz7iZ0
foVgHMwVfMLdL9HXzd54btO2DwTKvFImT42dVJQ950Xh9ihIf/m2JkKKP1s+
hamxo3bsOmJolTfe7fMHMnlLAOTkZef/pJ2R15hDGiPQiIZrTfxqV0dQk8XR
7kfbXZMYggjGCRAeNxIg/nJgEoH/ks9oQs3kfdqhn4LHYEeuZCnDObDS/4V1
Bq63PJdjn8vGDAYV3gcPAu+YwwfB1jpLImh3EGdJwQGkQJxCBQ65J+2Zx8Y1
CUQVLUZS+zy89BcrMA5XkKImYzPhaz4BxrZ8P1pHvDLkjARWStUaqmzGArdt
RFVqJ51lO8g5OKT0m7HVFAQfokv84bHrsixSXulcIqVh6SUiFrK7gran6jon
N4miNyyiotUsfs2LCM8WLZ/CtdOse6BYmTvQ5S4zTVdlkbcSzcrj6frAd+Fa
puV8gd8MzVcc2rVEgmrmqX1GvNE0uf17xFavwpxp+QdvVIEHMLcLxwS07JfG
A3J3FpRfU6tPHvZI3XuGawN639SZ+UugqssUqwPANsjMmuxX71kA19kINYx9
LYrViR47HTysOCku4D2wA08K9NKAVu9s0613kDnEa+8EbWpwuLUb11QbLtBr
xaEiYBRHJ2IWRrnVSgN0eIHgWuAXKnHu5LQW8ruKQqyQfebptaeqMa6CZMGO
K2zoyCxt5DxSBjqsJ7bSEA9mWeUTjEw3H4ufAooHONW8upDi+QU5YgQL+ROC
Oty4rD3gqY/sYwQo3vijLidb+49xXUVS1SpHEXlvQp5oAuCFDdx7jb5Qqy8h
9LaNHZEk100FntRbLxq8b79KRrbUltRUK+LG40CFGZHW3ScRQ1NO0JRXOqXk
la6IApNxLM5WdYzosq4xUixGNhweiaNRTPeqmVHLHAvd7oX+PJYLXzPn6foR
DM8JDKQu1yULCzPMt3Ir+bVUnUTi2vw5i/fSzh2JLGfU0ryfpSXvSWo3BtHw
hOePMzLwqRkpwOXIkyplaEz5o7eOofP4QmkvOkuziLcIFGAAi3/gLyHBovGq
0NiMPmIuYetpNtsChmKIYBtiohMo1td06uZoaPsiW+In26/6ikpcfIxyTrTM
QRsvzplbW41biJHqlCBQzwHoEGmKi/9zTmI+B323FcXrgOjGhYSUPD6m+1lT
1VPMm2mX1e5Ip7mWDzP7jLtBSnb8D+/iZPvtlWNESBpNn0mhwn9YBUk1hTDL
QtB8IWLpDRB5WBxiDqH/gaHNeYqsG7bvPRVwsajnfC2YSTDddGxi0t9SleuE
0fxLv7URWv23KN2huOziDKr8k+rr8AzRzyNlIY5by09z40nuQEEgm327yaIT
Lh7NA1LcR/OSZwXe4YJgkb/lZhJF0MwDWi6TvlM7N6FoUvC9X+s8tpbEwg/g
VwUrbXoAJcxiM0I6MEPLY24hzD4fPHW+4s+qX1bHEeC6zEaN7GJz28BreHz6
oMLjNSdK2Ru31wmiUWipmFx7Zvmx89XUtL1Ak4AONrk1vaPsACaLM4DoVmua
zdvBzY0I6P/FjCplklaXhvBY00ruGLcaqnI9zd9MfFIecXVw2NnWySyUTqwT
a7zYCNUvwMMpoO/sccqIifm4cEwLvaJcmBvjOG9Beyy1M9vnk+1cce/JcvH5
ML6I1Hct+yssSQA+WBrHO6PXLDAtaDQqJ6w7mLboJxqDtLByK63mKmhYxBkv
rDERSQhsmfWdHv0ousCHDGycErDVjb119X/Hd20/O6fyTU5SZ8gHIwWBT5K2
NLWgWqUQWAEqwGwnw23XTZxfQwrfWcHFt8XUc8P1SgAwXEs/nePCoyz9vysq
lYl4D6lY/evg4qLYeHeduM1GlNpMRFFiYCoXZv1NeHLhKSKA7ri93m4aCFIL
BqToOr0LDkB5s6EEyRJ1+7lS8PhD8Az/40qLdsLtPZy0Tx8N5zCa806wdZE9
nOK4XfO66gy7UYY7A8uAhfKR1kIDaytjTHk8T+rVGF4NGobuKuqt/Tbaj5ry
geBH8Ul+DcI9GisNjJ13qErkZ7iQyxwn0vAXdBnf5RrOEXW/kQB2PjhMZxYQ
WbiGMijt0ykzpiNo6q6qSVFm3kQ9On669opKKJwgjgEAnJvcF45mGOULItc0
mTh1JYPnlwkOo1L0VwW/l+MYuD7lPpgq8v5KbnxfPu/GSu6FF3y1FTpV2ie7
8KHmjDEaVbdnacQSQrlV2L4shngHWQDx7pwz/zqq4cVaysu65zCNAzVoC/6f
J8NpzUm1srlQUzXOXjvUzGIovyCp7bVjKsSsKbrs3fyAhzHI8Ibt6wcuMmxV
bkDpJ2LeBFYxUUFbY47vrk0kj69pMq20eR8M1C4bYSYKw5L19m2hki2i0HJB
qyG2fYCX/iBMTq3jWoFxdFJwMmCy87LASqQaimWwfvb3pPJDy12KaOztV+nC
EtIRlG0mIBpDJy5uFQ6TeqmCKZZ/f9eA5pJTc5s5BbAwpTMfXaC95x9x5Jdr
M9qrR/ICeVeBpK8pIzHaz9l82eurkZ+P1mhCB3+IZ3WS7bjtLAPGSeHhJ9Iv
IRyI10eKEi1Dq7s1FlvmZj6TLeAaUd2G43fDyWPqGv723O6X4r/A0m89fbPz
gK0Vtf2+YdAJebZQs0X/mkt9BNBo3IZ5jwt5G6HoIAZBVojNxezCTSTtGo+B
82ctag6J7PZl1vOL5BQHXK3r+6zlmeBP6+vjfv4C2ePWApNUTROS4Ue3BlPD
qKdYnso/5w+BdnT/1zxki4xqFcxhn5zkbkgt1RabM5BKEy9Wy8jG99ovO4Mr
wwgbzUFe/SCvqjFphOg6fGCrm78WnouGu8R4a+uHYxlzPfz7bxsSagbw68dE
nacqtly1QMOGDNoHXyfO/2vPcr0qlVCLFhCRxKrHkhQNTAc/z73n9PUHeHSz
4RYYUvq26MpcMtFZHLWAwhqfp/peRnflpdOEJ1RCbUM5YaGu247wIP7RuUOi
qpRPyki0rlT5F5hhWNGtp9rBU65zehkSQzN3JuqiRaGE8g9lOEfksSs6a3O6
AjIYL/O0nSj7ShHc03dEK8BfygwGU5hyrw1HXcanYGO2GgZ9cu282yAIVP9w
vbfo2yTit/znzllOwiDYael0heaAS4C0lM60qBLw+SeG1mHpV2O3bYKwomLT
mMDs5ptQvciV2GUj4EmHkHCTeEs3jZZ1gz7XQGgafIvDns0cC6eOcFUbJuDP
R1koWcrXyo+EtScK8g0SM0XATDK/XRFR7W8PsEq1b3M78lz+0XmF2VGHb6Bf
qZAL1kmNqpadHgF3SgpPK/EhbWRE385htwd+Bprm67Irco56Fy7HuOS7lZG7
BLeJF+y14cmvDWFWbtr72OoVHejJUEsiNZoSUNOGI2lTgI/uvQykcJnL7GAg
oEkAVAhcv89Z9GBMkt/LnpRXcD635SqVS+t9CHtvDl3XJSCzysEBQWkbs9pV
33Z3wV4tU+Mw9n4cbh1mpkUl9s+ZCki0+U/kBjPilYn85xNi8m6/SaF+ZoNc
kpJ5qu1NqF5xUnIQ62dnJFBqQPMOpXHmEWC0Q4xU1JAIN7x0VIBpsaLyadeY
PTa8ZrDwJBgHuDUUycv1qcnUngyvxep5U23KAEu9VQ48sWFCwRDmCrgIq8i/
t38MFwtxBTBNknnzXoWgrSV4jedU66HfY8SxdhwsOUh9DNmW66mrpgt6+PUP
esCqHLZT9GpnX33OjhBm2ptqbWMFhcVyeCzZpEjSW4EMpryI682EV5Wp8viV
gA4f2RhKUB9uz0JiqZgdV77VhpJeaachNql5ekBeHEyptRfT5BOPlxAB53SP
0nkCYM2vacgkwzZgFIwhie8ylynR4NKZdu6k3ELa/+ohNQuhfrAN4kc+8afJ
61MXc+KB3oYRXhuUw42/JVN7tOHuO9I1ngASY1vZskghXPCEzUkZ95uj1RYr
7J5MQQBu34rngdBHSgPhFqxE60t7jUWS23spz2JwLx7miTyHEK+iXotgxo+D
6AEB3y4MeB+kE3zarp8hRAh4XElXtX3cTYyPyz6uz+4VbX9U6XI09AhWOAt8
DCVOYx+bV0yNYhq3aqWvlXFf33sjrJTN0GyQ8R05BY6t5uhB3DrGh3Epplhq
/AFs66JRTjSXy0t0qfIHRuDQJ0jOgP1EQ67Sr6O4cq8R2IUh8qiIf6tV7/pP
cdkhSicONTdoO5raaWPH9zJcEP6EI4XQV1p2hKQGLbi0PsDwtGzJOTAmdb5/
e784o8GgZwFW9VGGqdjl8sKMp8rdf2YLew/sr4ipZwGPeBFlwiAXdGwXBhZa
rrHLxqRNuFuz793pbbOD0MbccTmaXfUFmnI+WSVaR+MuWqDfc7KuF5u36/fA
06+rQZT7EqyghkfpBYLcSx+lLXo5diEmfSlCiCMGOHw3kESmEnuaI17qoWfB
tSHutGo8XkmlvxzEuGRX4GmR2gAfJXwqZaRrH/SxDjM17mbOqhks+b6eJdYn
OFrU1POzA3Vv4g8fLBvygoOy6MUNU5nhvYp3AhZ/y6RaCwPBw6Pjgmlrw45U
3TdRAvvFKwz46G3u/FOcsAfl7bW4g4t+OUsKZ4ROAZ44YzaSFs8GKhF+QDbO
jQWxupiVDqJkHRQC1wfQRbwsKizGwfhYCe1ppR5z8y/0le20m4bOk4BqmdjY
ncb/8mD6fIs1tozdHFWpIjw5SAZhmbOCIvlu1/+tUIhV1G/ky58fElW778bq
/zH3saFwwrisFIG/VP2pP9IxsncpwXdpMNLYAYB6q3Nl70tinpMQwrgqw09M
+znOubrDo9zDHqtk6bTJD2Eerooi03OrH4rjhEvu/5iX5KAj8Ydi2HO9CwOC
GWvfgqRIVUDlwg0LtIftCxLkd/qV5KXGBr73Gwd2RSYoEfFnC0soxQa4PXmL
yu2joUA19FE3dvGAQmgil6dpFB6JbN6fBDXrgXgY7ukaSRHaRO9QhQ0S34K8
TxBzXqtzLWAKs+CAJHbYXCv/dsxSasr5zsucPxRBbfRpwlZod+t1yqzXOiVt
6p5R4fwWHqC2RneVB4Jwxnn/05NU6Y8QeDxDsiJebgKbd00mxsMzDN0KmmMs
ZM3YNizgnYUZ2tRb9wwuTS9xsPD2NRDeEx+iPMkVDxUxOd5e8YK5qlNzH9KJ
S0VRq31iE5xDQiDIkFqhibxMArx7ci0uqvcWJolMF0XU8MNeVWl0iVdpH/Ww
J3NSe5kEtV7RYmDTI2mrwHBKpRaJMiLgKjF9Fvp95hxV+CtCnwUnQB1Tk0zu
M4BVe4Yj/b0XU8aula/Np1rK7+nMUJcDBqEg4bBq7hNIVcmlzucidEcjFTZP
mJ9F8p8JOzOw/yDAmXDIEgPHzHrLR3TNmjPMgiGjTrzvvWvW4AbYfRSQNnFZ
D6LP0dn2QsP8lARqixCn69z1VHhsNaAb1d+pUzYX5imTyr+hW1dS5o9b+8J0
TwEnievarlwTR2FBBkeQPIgxcCWaD1io0csd5hFKQFW3x8eQZpMJ67VOpyT7
nN2YfbxaQIf31wt2gtSPasjJ7yO5ELaAvzOPeL0yFydkmzb36AZATImzZeie
OaaS6I2QaGA36sQH0D55aMMVIxpDN7975iPe+efsKDnHX7rdtjKMtiTebe97
uzj4I0aQC6clT6s48F/G2VwtgdaWwINRtesFrt00aKb+sltz92jLK36NUpRA
xpL0AGsPN/n0TaaJI9Q6ANY8mLdhc44e0J6IVVpJKKlYCN/MLR8vTkOG41OO
vmE4SFbif/L4pJE/fM85bYIrtFZujTxnX86ADLDvlNcvZozOtVytGQ4EEI8g
wwNdNb5Wsdsp/NgHMSOF3SQ/qifQO4R3jHJlB+3mq+JQBQyrgbQrzrZ0aG5T
OEl6gQw8FJokeyQDN09cgN4Ncf+P5A8RLr3hg9iVwCbXfG77eZLuLvp2fpjO
U2Mto8xooErCC7fu/RwcnJoWaEYuCVQd6t9BVC50hLp5MnDOKCuq0q1thIiL
6EbD0LoBpFfaaGPGZT2pHJFflA5y68V3E11Teun98C25vW+0Y7VY6nL/Nt1k
BVa7C/KQfwrZ23LtT5jC7T9hQlGNlGEAsFjVhfXSD75A9rmElElYSXIhLmE3
6JI7JfbU2xObuozuASRnPq/LPws0Z23P99ZYoA9C9RmxZ2jUDgSAu0uKbNGS
ueW4Df2P3mJ7My2qYjg26B4S7x1wnez9pPMzZ/3nUcid2aW13qD9oHKxfNET
lHSMnyE5UYAQpiRXX7Aj40BT6Rm6w5PuZiwSBtT/Lm9Rr4BdQUk563Km+/D+
sjv7y23ry6IBr/xBqFPZugV0Wm4iZFU/p2IuwDgMyiSDtbZTba6yPDOOJidc
l+WlFzbQmSd0IHVQYW7tMPmcUlGgqXuL0BSo6wemdW0qNYKsW6es9G2fL9n/
o8vEWRRC01bqq73RHDVtZ+rF3o1PMqCzNnVvi945Bh04tQrPsIOyFODbTYNr
i1FqX2aqYnhKl1Ec0Q7/rAIdhSWuHSvYvq5kl8dyPS9dKSb/qzPi5afK7nAJ
XwU763qgjR3LQZn/itz0nNSRwe4JSWMWhUY9+uOEv78VIn6tXq2FqJ+4xWXs
W6+P+iB6itprr9rLgoBOrfnVdkQcu/xiS9UE2RT+dGJMJ56CNMKk1FISdsdy
4ZG3O1JsF2YtK/aDHF/8wKI093W/wt6P0NBdgmLrf1Hq5RkrZCYTRJvVkGvB
oXZAzyS+kYVyILnAOsD7ELbGAr5l6rbtsi+gmgOrvH0kXLVXxnjDrbmyRoQt
FJcovq/bNdM+PslG7ADK/Q84hq2wkxdffV/aFqN80efCgyv8Ez6PDcBSG5Ik
GQmKvUA9S6/Vymj+vsVMILj59F5Mjf80flnLVmQqCLDFy9rjSNajMmAeAhAH
erCs0/lcylqwNex3xDArPB9MQimkB+awXj+2ckg2EvEog5Q3j+jRs6s1h7AC
jh2yIOU5W04ONxiE52VEOLO2adrJ7HeZs4MlUT45aHKSQjop4rtgFJNf4T2P
x/d9CrVHiNry/Tvhim0bfKVhHyxAPKCp/8kBg4pIGcMuo1zel8no1kDuPQSH
lMB5JckAALxfZ+5f/oab0bDKPuEJEuoaYYhzGkSvO3IpwEAkui77ROndH2Vt
fk8ScHMMU27vsCyoh6PJLWLj2e7V4pj7N/asCHgSDZYEcBIvvFjUrBfbiR9g
DwYtZi/xla9gxasXy40tFrlRSu6SoR1fobCP6u9udcBTN8U3cLP6LYpTsEBv
4N1mlLOhB/JRQ1BpjtKxOLEzGM6AGbBvcn/g+UODgdfyCcRQK0QDGiBtJ73g
wnCpqohCwJf1WmjOh4e6BATBSp6cogwPLZ7Hy5jpIjUf8faxR9Y5NEAbp0c3
rOj4xz/mfVmrOmwzGAURz/y12FsfZh3Z7RVwbQc3GgYOhXnYylMLKhHElObK
Xb1fQQ+Vv0KbBP5a9eouHZzLeeWlPCDcFQzmDP2DTsSsZUwUxXPx7YqLKmpL
X9lirsN2Qxc8ISYgYrQf8joOS390xZZ3V6VCAL3L+xiDCyowIqMRM+hmyBt6
rkh5m+VcnMvnjTprXVQGdqVDViWUyEnOER8nrih0nYVkDchJXIEVdnM59m7r
TD5GlKW9X84DTZCjSawzSOQ4Hr75ZMqIiG31rlRYYhyTvh84Sx0Ft4V0sulG
7BENeztHWnctltYGbAYwdYq5/+W7/7hh4OHtaqAn4jYLWwv4SEhthfPUgKIs
02eesov+bj4g4qvAHdBAnbAUxiZpf1tvgYoCtlfwT79ekOj89v2qrhAP9Bcy
/18qtWs5dWB2pAYpy9bymP/gb8DlifXQzU/haZFmeKBk6UI29dxvrV/A4nHW
SLri58PuARxB8XTgCrZWcO38krcPjwJT2kaVkxwzTIzGawpvbaOvJclNoJ6t
DizDZtMo6Q+XURBN7LYrKtm2RaL7r+SzEIQGunT6UAW5ibsAUJGt0yc40AXS
bpAZIPH9R4roRDA24qg9dj3BypseLOcUEjBF5X1gB7pNXVfAgKq/4GD9Z3t3
P04ZLK6pWM/P842Wu8PvzR57flsEqB1/JBdMzPeFNEEmq3SVg9A3R71MdtPQ
7BeIOZmvr/xQ3d6lE34pr/hKgKdYPoOzJpf7i0WSyGIBgSzef0fiUPQ4+IJN
g3dKBCkhjhYlrKL19KcEqsUOt4IFu094RPvIhvwslfqp4tMb1/poOZB8mRW0
oPFYpIIfTbNtJdLizImbjnAakR9vGeiUxSO8imDWKGns7NJys7HRmD44NOFq
2JPghHYRl/YgAmOpjgpyHWvPrgx5wV6ZWB48tq/w6KwHgfx1hEZmMfdjbayM
lHs1l7QbFA6VATYSpQjej2IaUt47SpXoaOH456R2nvDb8SHs11secEnzQ/iF
mZed7czyrsx8tEGFiEBu5WXkLtvrjDHuSYBYFlEa0c8UbAxF7n4jLE4aqZr8
QfLanuMSZSfZUDJhcYY4yfACFKO1fbYLi31MnjBNY+WVGfQVq9XzIb9OYF+G
flP1Gi8icFbS7VnCfDBV7xVtaIS3bXatkO/b9e8zj0R2/H/noDCGol6bwonr
WSA6LYCFrHNBHoJfiJeYPk7CaevF8WWqBUPAGWOkPRJPHUzGaAZUaAqrSX5C
GxIGyKiSStoFpo7kQfUjagvqXkpF0S5RIqzgpqpe6zGjfoP7Lo6qGGX/lDxK
0Wmn1bwdtUDzMp0BN+ZzAAkqU5GY40SOz9RkAuXjTMcRzFo8IF8fbyL2TArX
vNmJcvqu1triqjmgoLS6O//uav+84kANgW7GmFjseQ/bh97CTfZSQnvzm2Cu
zYH6KfakBotF79wWRR57AwOoTLBki2Hv+C+kR+ezZjLq0b7+Ylxc6mcmpUwN
VXyOPpFsRG7r06SINt83N7Mofd24SPznueoEQvuB30Pw4VY8hZO+9AfwSC4o
iQU+i40cfRLC7Z1uI6fwiUrq0oLsF+W2FTSq1FDLAkm0u1MSUSnfr9STwn01
hsnrXZBtztZ3+uIZ7zsKsfgTx9PqshP2vDE8wZxFjfIqkWmiOcEBcuqtqN3o
kojXBph7B8aIDFx7ilJHoH7PVZP4Mod/oR54uGri+r+Qmx1KwHPIGYFov9b4
SpCN/WVeRtPBH/j3/6yYM+4n6dkt5TrTjXIKg+2RYKK12IZctuTL5SbLtyGh
Ti3dTcvJCLidxBK95GPolLvwGZPYtrqp80XPOBZo8GSAmCgtuxd0nqJBLbPf
o2B6wW1z21cL5zN5FMFe52SfqP5nrbqZ/+PhLKolQymYqNWAgNF9iYZK5q1Y
dU7oiowMvp0FGokqfy/gJC+7nUW1bGYNa+9vw2oAEQBmW39dw5GoHoS8pyp8
PiRBbqhAQuQ7dhY9je3NJP5w1TmMfuQOjEe3ss1NBOzjqEJhuxKr1/8ySnGh
eYC4JeZ1PhOvV0/Uzr4iJBNUQP4959Zwa8fIdfiTEinKGYcADrr0xvzvNY6D
1lJi5gGt0+FDfN1nVhubJsU+BgVvHL7BXFwXlYdok78A3yej3vD6ahkYRHi1
J93+1gkvxjR4KuIrwRZFWIFvAIsYSVcmLAiYUPBwF19MhkNNaeZxdHoYAWaA
9DbolaUtwH57XM5bxDQBtDsQSQjQpdEaBzC07Yu6NeiNS0syp5Q/vQ3+5TGQ
JV5FUjmwySyw3xLaslSOhc1hnDTUx5x1AdVgBrjUx8LmQJONw5+1+mRvlrSK
3hCGEiDwwWyS5zwdYfMesHoJiTFgSwLVE70IGy8NDc+fNsLaHRCSTIqprZVc
CMfEs+MkzCcRoxAtuH6tg7ygINqcQthtuajHI75OWEYTETkMrwAdY87NyM60
kftR78VZ6x8TM3QyexSI6cMrWBVjf8VBfjqdKviUx/uHjhywkzqCqpNTVRGg
duhwhgJW9kTgquekS+HgdRKoA5plcdght+rRUKPBFMgqXYG8WMeDkmrD9FRE
B6nuo8Xa2RXioWl8TqqFwScZ5Tnf6TNwEUWM9I3vRWbg3ghW6zmpmJfuwII4
ojTM+5ZCEuUbEC4YeT0fM1LYsb+Id3QadprBaj4A4ZfN/lpG9tpwu2oRmsy9
O1+wHi6WYC3lcC4Z/JvXRVPMdDr/6s+sshK1R6a0ZGlq4BqmgnSV9WP66vA2
CL4XJWN5VRQJJMXw5gI/+7ussxhrG0hYjXI3glsiRyRq1doqR1ddUUVdPmNJ
/ByTzCLmYRQJIeoe3BknrASTjyTahpE8qUKHLX47sRsKirwgAvzeQLbmfL9h
s0wqDhr4fNLwzyfcwV+6aRp5SeBZPjKb3NlJYA+Jo4gIyB0o1n9y+zPq9C3j
jcnAfCVqphDWwUHM+ghuiCuqbv1un6jELCiVA356kLbzTbHE+O5QA3BMF+P8
JiSDf5lzMACSBZtk5o8ziuRTRH8R7vBdfGEcauRlYv1N9+yxxQi8d6t8Izc/
2UXR44m700t+kaNs5Lu+Y21b1UKO10cA8ZlWLNCTYYrzZP16T50btCOrpFC1
VHCpZ5wQp2JxGdZALEiQ7kXFKAguCvMYajN3K9QukBD9tZxHPxk6XPvvBvWQ
ipPj2Fc6UHgngrts0AWkzineTtr7XjPEYj+bpdYeV7cY+1tvSMIaV4nZ0bk9
BA77cpaScoklQ0yg4kHFaSRhhDQxzdxnwijxI3SeDr2yvC6uldEqfPXuei4d
TWpbC8Uz7d8+Av3MtiZd1o0vVMyO2xcqAaJgHnloE066rw5Tr6qKkpU82Klm
DQ3Uf5rlz/eoCHDBIUaI47Qp+rRrcBWpd/RE2k+3PPEdaRJd9OZpEhniu852
p2+Wu6nKAMsJ6GE7h7XuLcGvX99Dg/xlX6k/BE008u4NP8BxBHV1C103oCY7
wnQfwnEoFyy0FjhWRqL7JgUuRXSCgkXf3Jiue22ABgXtN5bB1UmvT6DMzaeA
RXKCmnTg1VN9IryLztEERQl4K1lgZa3o8y4iP3bZkZw8OIhN7OJFTF2IK//f
xJC/kcVlzNoJCSgMZRzy5bS0xOW+z1KoEzokjNGAh4jp21HXji90cZyzCtZh
+Nn6abSYf4kuRzVT+LS373kIfKo9zNL0rw/VqOE8yj5dGx2x2+QvcDdenMtj
U/ywi20cS+1Y5iMI4IEMpWrqc7eXdGRgqQaI2kUf+uvMz8VbBg18BZp+O8ih
qJY+2tKGBiYjva3w/kkWOPKMDSeQATPydLNgblRCsHKzu+9tdlKEB1uMTF41
MK+hS6suDsN3T2L3AymKWrzLxvKfvhrx1CueMz2hODniWDd2pVD3mmrfStcG
MC45M4b7GCR4RswFpFClQoZDMP2Eaw5qLQRAciDJs36jpb7QVg9YqzRn5r3f
8Y55E7mfb6PsSXOQGIo8WTMtE11hwZndTMD6ALM1yjI+eqhp/FUwKp3BXboY
uHoIz6gMVh65hkShCGATLRsurRuCIjqfF/v5yJXtN1sJUsDx8Ir+6Vznc9lp
sDm/pskvJpEU5NV4RLQJwLlxbooxY1sOxKcVs4fee+Wr8iaO4ozpOWKtk4n2
8XhLWA3RDCEvHKEBxTnro7Sw8c+c8oNT2CqEHDvEn2jRcmQymoFbsLM/V1Qh
aavlPWFtdh64esxPCB3OS8kvx/jNcXclNooc6O0fqI3grBTvmdcTFvyYYMaJ
hsN42LMUGFb+DmiMaRc5ShlHmHNYgP3oYk2bk9UfvK6ihwuEu2FQzgkUQK6o
I9ZYlIIUuX+U5AuzQxsNB8ebasRMfJcqrYS96VyHq+yyn5vnngCU6lkirZ24
cdXO+Heothzby059iLpyg45dmx4T5+8GVBVZsoF+G743tHbuwh81z01+ycuq
uGiXTc9OeCpEYzHnc+H+eoamxm0iyxkBEB565n7y8tyNV/KFz27P7QDJE8IR
Tg7o7ca2uUR/1xYJa/+8x8FRWroEPuKcfwCE1p1zA4Q4zMOdU6oNVWBghr2S
uQ4VtSdV/VIXJzS510FYA81HHyxCEjqnAOnfLUa+r7Kwa4D4mvFOf+MI0xmX
A2gEXLDfkAAL7YzkoltbrT5Z7ifrsrimTNWn0/i3poIWLWibuDquG/HgWdgo
RCYR1sr/qmV34wvGHy/10mJgfnD8A1QwnD/aH41Eq7jHGLAQoC4z/J26Z6Ht
NHCCOuVjk2uKCXJHV24AKuTivgv/rYY8HGtXu6eR+tAglRXBT1tE4v6bHYv9
1gya+x1918eX6fk9ISkKQQKfKht2QT4YCYTEz3g6M6ckP46cxiXN3TUmQsWO
eZ/uQKq63gX4rJ3J0jQdrPuLuFPyHKays2wPX1EVVf2GK3Emem8hUuYcIU4v
g8vjQoPN3cNsK4x9GePSNx/7hd5y04sKbFWgCb8ISFOMK3iCaph+dDZQl667
8K05JCWJvRQyb3/eXD+dz2CBSAqhUMM8TvQZtGQ1+6+DqNCkL0FJXQCG/FYH
uPb4saL1J5iHTjk6DpzmHL0zkCGjq7HdmoB3xtd1rgyOTsamBNDxmwxkf/sT
27jQH/ljjuWkr0/rBogJKQR7T7G1VheS5Mq0bVHieiIOk0tpFZ0oFnTYyx3S
qbB7YAg+8dMP8rpTOKU9394axjCm2KUr6/PhLIlooaanZoBYxcwdAr2tb764
fMp+8B3BrGslQN4YNG6YY0Adg0Vj13FNXvifpxaQKqOSsBcUeh1CNt+OLxE4
iT+FuaEtF88LHSnjbAlwnUXh4km5AqpJTURj7nD20eSt2vE1V6qT/qTWgkan
x5ix78YiqPRHtVR7dUY+JYt/cYxiTD35kMOOJlGZ0OYQsY6aXW8GaRmgbORg
K2Kk2AMTyl74rHtlqh69HTpI9aOU5Tp+4jwn0zuoFAMglxLOiu6Uj3HIID89
T9oMRVjLoeSkkJWzMziWaUShhzppQ3SglKZb6uR3Sbg0iggE+RdkXvRgiv4r
jL1S6z5IP+J9qBc+0DurPy+ZszEliOl3NDKAQ/vDj7h9+OYIVBL9eviIRVgJ
+RaRTp9TD9OCSYW92ufldWKLUSB3faR/WpUKwwE9/vC4t/Sxy3G/Lb7ekmQH
2Csr0ZdMLvwnARlJoycyqS2Q2hMkBIYpRlDu8k7k9F5MgzsXJG1UGPsXz2jm
WO7PoYW8Q9+YorYaUPZ2RM6EMSrQ0/YQ8D2mkc6UoROJzNpF0/DvhIcEfr8T
Dk8vF0KNv9m8cCYmuEwdhyP9Ym/8edqU/eeLD7iS4M1G5fqQ3qzOXgSwb1TE
pq559+ywGSjp9SVEdIgMHOes5K+matsvT8MQoduTJQWfSYc+Wa/7Po3Itdr+
IV9D+7i/ulIvGnOap+KJgRkgJQ6xwIiF60Pu2r3ffmH5090ThH2+b/zFUxLw
qBgC7MNSCp9u+i8p97aDC1w600arFbjWo+LxX0DbJuajVfJQesKRb8zeJzcj
PFb6RU0REiz9rmvshE0rBs4OyhSBW8sCSZ8FvAWS7QcI9pMwtTfSvm+bKBwJ
Fs0VO1/qPgFBL5vnjWSTL0Za2XWEPLRYPK60BUzt1aA8I+s/HCh7JeohE+PE
gpPWfn4bZpWL3K7Yq86NVZt6xPTO9Ps8qMvL2GxelZYflNerEuUVaJRfeQxb
P2bdmHIoxyVq8AZsVkXJ650MGHkmIcM9uH7hlYWXIx5GN10b53VZEHowx8aM
oxc23CsILr/a2OAD4/MMzS4B9XT/xE5a/+qEolDlpFh1NHc26+PngvfJOs9P
EEP/JP/2l/eIBE9H1DcSJWAFJDqp2oH7gIiuvmFG+AKuVp8bOOnAERXhs37l
oWsFNZBAOeBqBSXF5PAExdTsYGMxl90pyipHz7QekDTBfzuN3fWT1rK1jBri
8H8kB40AFCIAbADDgKPFD/xJtztwT717h8dTolZFuPk/7EB/QqCFMC+FQe/3
85qvAUqAVwgDDzhwmykiCNMfhN4Dt78OWNRhIlPgGOW00gfrTA+HgvuXfebq
09MVUaQizJx5TEmzi84gXhxzi29sIkJpLevClWWx/tZgFpgD43dtBimefCuJ
QS/D1rLYD3ajM6qRT2YFB+p7hRkxpb6HJ5chg5azFec7yIGnDyNud1TgJc9s
K7UPdBX3J8il4Tg3AjpRLpWLj01dh7yDncEzMBoxIxhKb49Myj2A4C12iO1w
pw5SsFaqw56MtRjAwlv208MlRBReAjdzW57TnifY65q9pMmjPYeuS9IKRb/j
Vw26yya7piGXIK3wZomhdqV4X0MelG137cGgbcH5nQdxRQKPdUn4hbEM5IU4
s/tDehTiBkXAPjK7KehTBqpeGelJvznYJiXl2tRHROMwZwRq0x5U6KYmQbDn
NZH3lhb6DJ9pqJwOQOWOkNTLREB7qka2ZgWPC0mveni9IAdifcJ4E0Zk7b/L
b1t/+dyPs18xO9n9tqK7qvXef5eA1bCpmbnMUZONwbKH8dHRlVCqYQby47px
X7o+kKf0JCoXiP9HY4mfFUDU6D3yn+Kk/zm7E7K1OIrj+j25EZw1RTTI1J5q
n9DNfNBlDth74Ou0vkmyFW3Gv1rU2I0B5YMTcPxmEdcjVKAK1vofZiY2pXcT
8eDc1X1IHwaMgReYk/5jEgraVsF5BAMwgfhLjFaUWMAc/dblMS1Q8T0xbN/a
Sb+8a/LWkXzcdJuV/rGuYCmS655v4D0HwODVZxul1Gs4cgRmLA2aFP/Q8sEV
KZcpH6BwDVxjKY+xrZ6eFlejRkTQgUQZ0w15iP082upOFzuQPve263gJt2Fl
eSM3jAFcFZFe9hwV1TgH7RI66a8L7Kj4rFCbPD7HF8+y1thwpxdEmkNks2QM
Cs4Pd/I3HSsMduqxo4xNeTo7Au4vHlW1nRCSGCdTKJAEyc1hSgBqyJHVZCIp
KKDOyHT24KY1fm8qLy94FGrQflIN5cL5j7zejJpMFFp0ndHzSr5SvoHbFwVF
Q9JIFg7INxATww/qOhXVdR+21kJ/ZBr2C2oyT+aobzgQy7cFtMODoLHY8yIM
W1cNmqCHxjE8gfazp30CdKK3+RuW338cijT0ZTYelbA7G0nCpTO89t02aTez
UX+ZnzSsYISAJngqnN5XyNbkWjlkHwxGJTqvOvx29AyF7thH+TVZS+l+aa5C
k74TR0MampGcNOROf6TkbDGG1gleqe2K9Rt9yg0IYAySb91nl/xtaBBEDF9L
4gGxN3N+z1yk0pMhVRPxQLDLhp24ohtbEZQqsLlogHMitU80Jpic94HPFlev
xyuJcQzpkYCFzR1cnSFroUcFUmZ2ouBeIp79Lj70TMP3gmfD2Gg6eakgzGPq
Je6GkJoo3KSzryPo7mkEH1U89S8o9lk8wP+BqPfSlnO7hgScPaM8xz4b99Be
4W1ZiUkgJZwsUYRn4TGm17CPgEUmaDmv1t2DW2Do7Sf2OJPGmKR21G+f7p3p
I0LL4sJTJV9pxZnlB0aHLT0yvFMUGcenxNu0j4pfdJoqQE3N4vySY2vI0mHA
wtraC9lFWLy2294+FgP+4Ic9XGOo2AuEDgbJXqi3o8WOqd6j3R4UV6g6tqra
E0qF1lAuOBSB1urCnhwIWq3vD1HakRTLRn8CHSJNFBu0jbw4pTarqFKhlBwl
a1HwwQyLthnuYzzorNlCFifBP/gY47atM46lGQsKR1DX3QyJ6EJPAyYFG41J
aeS1pok9lZe6VHvTHbLQ5nNP4tUjWD8l5jTZXOkkRoN0+Fh0tTABCLXdJfWt
65omtrFA96hWvNjnsFlCGCpT8ARaJ7II8h4Lt8z53CMHdhCnmO9PeHFbKBMv
Q8bg0qDU5Fdfs992OJHupXVn1cftPDyceRRxrjUGfqwnfOQY7DN+nvjnMm2q
iUiUzHAuh3/T/kkQ2DtUUD2FtLK5YBj32puFE9FGfIhaKEw78QpRpEmHLymS
0j2k2WsT91tkgWwviwsLtUrFNHaWWxJlC88ogT//1+jEhkgB2bvGbtslw40/
DBeqpv+QGXqZU5Mr84wnz/jWXIBjaBzWiK3Dq/RuEIAg4vMMNCaKW0m0aQ2r
uRzYJwYNBICMif0gPA9F8e6VF88X3yyKAlsO9vyOSwQshS2s/rskjeNy4xL8
sExBcmTdJnXGwBcITW7u1gnYU8ZPoA9lhb/QB1rRLGkUaJDonauYedsWlBK2
nP/oNmEnuPlnjGL8Kxa1mdYfx4sb7LqY4Mzq5YOpD44h03hmbxe4m0gb+VyO
RCx+ktkz61X5OA37Nmz21HUdez0/iK6/eZ4eAAumdeVl1CdzS3yY+jJaG7/g
60Tl2F0Clqqb+6zdJMj5epZXL5RXQdZ1rnIveaXRcmd7SH3cO+cPsqt/sw5/
po5PNTJi8l9vm6V7gX79yrgvrLed0e5FxA8knLIkAIigFwM+93beL+U5LiAm
9479JkqX4k8r34a2W4MHY1UKCN7ammLfe9wtktxf9eYWWm2f5v2luWgrSy9b
1uUfI2A9uVYEp0nNFpILZ0zsR8WxBiAKcfNQTbP5spT4NEI5RPIS4q2vHZ6I
S/1nV/qwh8MTFCE4feKZNmAMFPxF4t6cXJQrkgI9eAerW8id7Ze25vcpGYQt
CvzzaN9+EcRwt5dZsIJKhuqm374rhntPtYo3KdwQKasbHxcWiSFpxpIww6Gt
YTPr21bp27iK4M6gHIX5b4lfzdij2x9so2TsJtKghh/rSQ/EiirVfUtLV7XT
ZmWkdnl5CC3WLRa5ruo5EGCSjlPmGmcvV12VB3M7kZcrc+u/y2AZl/4Af/vr
1P0y0j3sFckoTfAUss2NQv0AZUwW7Os4Uzsty0OMq+2jTx1fP4VUDwVf8LRU
+MVjUYmte13UkjDn6PllX2iPx6PRTSKtEGfgoAexOGlnUXbnC52O+9fVC0rX
jHzMPMOJngrrekLx3fTXYWbGbZiSmqR600e2R1oG5qpwnajccunlDLxahsYd
QfZEon0yXydGWS2qtYBUNl2X73/O5hZmmml34FxWkz6n+RyatR4ogXt15Z37
ljGkaC+pUKzyHb+2UjdfQcmA9mTU5aQvLhxSJacGJBb7fdBIuNVXyiJpyqsL
cKP43Cr6UvLTWJocFw7R7ycNEMuBptuLr+OWS4ZacJTYfb/KY0pQdUVQyyw4
KEs5SQvCtofZt6xsS2Qvpdyg71ZzhcKvpraw6cao1/dcrjbv3YbMbnArlnE5
zoEkGnmqaq374OSva/qWjY5gi/2C5XSsh9x7dPMgUctRmQ6noID1YPIHi0tg
+kYUnpFSj/pvkmVqrcFgORjk5RyQhXgcqp17dtCTqesL95tGYzVYZnnRdTIe
1VhY98nvnoKOzGg3D+AbXoAhh/uDMFO0cOTeePMlbfNYjq9m53LiGdroAg0O
YNdxZhinJigDsZLIFOnQdLHC/+IIeq8wRSN4fItH2dr51a1UgVA+b+FLT5+Y
isfhRZKap6jVI0GfpMOuh5YMM/7VVTFn/ZUr5YU5QnYwyPPUbxkx16wZkf93
OqfpTM16k7lmFwaka9NXbinNoMyocbiYe6MUhkr0hDNbJAxQwO/emwk5tWH8
nouCw9jtyoHBsdGpHeovT2uYed/FpTbflGpdrHExlLjdBiEPgxvGAN2L6xMo
FLapZLS9SHTqPlfDAkRmu68V/L/VaA9/7O55AqDNGFprwawYY2ksWCX6ipL+
IRc26CeNkjI3sT46+X0H4iO1sBDT9sSt25cxzd5YWTDvQ5eH6y3KzTfyjsN+
dJwuDIdK1FutARGETYMYcfoI9QyfwsNj41LSuHdiPJZEfSL9QJ/sagbo/KpH
B4racuSva40zpfSNGp0DV3KzegmfFy8zOwFsStqDwT3e4YHVUV6NmQtkyIBA
hpotsZY3fkjPjHr+0yao0FZAdX9woVIEmSEiJ8dJ4xgBSM3EQXQl/PWxXUZP
NNVH1iPgyPWyEByKfQOufHw/3Qedi9nNC3406d4aSsTBSftz1kmHS5/OyD35
mocBBCccHlL+jT80bGmWvoV6dncX1F4hnAl52mYz6A4iID+ciW1CIaen8lRi
GcWBjxrT0tErkU0vv0Qf2s5kbypSkWpO6ERJ0o70eD2IPOEvBOpubqsaah4t
Fm134Cut3o4omaFtA1JTwpI4Az0iNsjBjPKUAEtwNEOlMium35UrybxbxjQa
BA0Pcxb8d9ZTMMm/tF1myjAHk1OjTyOAjMjpkk9xJEgh/vSwtpxoHHkt6El+
cQJCMOdKNONQ8ZtoC/m7iu43ssskTIasq6x9IVPFfGRp/qYEgA3YM431dJeK
lqADAkxNmAKsCSHaRznRc8jgKTZhOlp1BoUWHuZtTuPkT4WiI51rupkOFiTb
tKmsx40tyExl/epeZw1GvEk9wChvhoxbBIlBIFMmd55Q5E3QFXSOQ6eQVQPZ
jbuVpRdge8n0IJ0/l7ZCx6V2dhoNeXuaKxKQxUocnYt4iiHna/N7NqqFCvmZ
KwfSftef+i55Wc/zckG2CbQDKJrE3qQDhkw2TQSsTLmVpv6nx0MPRnpX/8OC
CFOkNPTCv9Apr0RLlBxvOQMNNnHu1ntZT1HnLDxE09bay3D6LY+5C1AewMwx
LexqQfTeqR9W3xMdaTebNTKmqUNRYkcoUMMIddLcBb797ed01X4noOzbx0ZP
qQ3Vaj+jAL9bhalXpOadE6+0qYSqpRe5EQFPRjfMrpTYQrIgfVnsMH/ZX+KV
YA6+oK83WS/3q/m9k3cCY1iqdXzp20+YYzNuDek1IbDHUA3cicEPeQNSeQKc
z28khUh7ZPuktdEEbZnXxzh1M0c4kiHYWQ4cqFURZkcr4fqRB43oFoQyTIPk
b8FfipJWoQSWRias+T5mKUBS3L3KkfWStgQ9LKYcYIBb0r5Y7NfzA7HHQXVE
KVlnp7xymOr1Vl1jwry5ygg3oMvqSfy9gsAVy2JLSvAkRLqfm2avTJqMw2Mz
BgWy6xJmkcmU8OwVRrpoQTy5NNJO/mjLBjAaDix3ghr3Gc1vx4Fa34xHDEPp
BhE+p2ac7CQowS5s9sfzyvKeIqtIrbDaxkEXClahxnUM5bWayHFkBaouP/TW
ct9HTBKxtqP8CaX7yHtvGH7Wp9iGqFP6S2xjb9tQLWciNR41m8Xd7UXsaXF9
dp4/mKXKXC1utHYrgLFkHzBO0acV1v8FbMdKITD2b7XFk9dyphrGjkrbiL53
777/yUMuApg4ehi5QjWaA4a/Oy+KfA2uUoFkEjkeuIaygkAAWkWr/zwsTH64
sOGnTsQXMzYKFlwzrRQLlKOYYnVZwBs419MgEGi7+NFvS8i07EEWWzJ1oOu4
5pe7rdiNJDPiMwdkHAcgL3tl1GY969rl8DWavXTO3LBwIYbvHnF4q91X4DtK
3YocokMjoTa2PI6D4kIr2aBj8c/amKIDXOvQk/E0aCTUG/gw4GBoZvJZE8zV
4swrA7bmyHHY0kgASfF9sAZ+rTzASDh66NHjXHQPPldzWV6hsHwt2RjC+kMI
I/ZUsozu0fLNj2clWz3ORzKNwf1oSmDGCkc0RWjYqHEW8t4ceVttLrXU1ZIU
vibnckPNNhXIDbAuAuTknIh1Sg15BruzaRBViGzUY5TMscsCpsaaNYdT4xx2
DKHx/UobssGuRXHrK6FufG/E2T8b87r1YpKmVAfhDGDIQGgQ8kZ/CPbReEVh
toQ6jPsJaIuJqbf7+xTiQ87dhS/0pbqhngruJzPvYD2ntlVOr+B6rk5FRKBm
V6vMa+Ii5Bn3KFrgUo8eEovzUR6IuQG0J2j8A1kzcLCk8ALrZInYR6sRI4qG
QbHBhlYk76VBPlDH9NHvDD8vUnbUhABXzK72nJ0DyK3AwMSJO6Cn1DtN6B2f
9PmI8n6pMtYB9yIZ4p1k4NPHSvzfYZkvYCjXUzXM/0DmAqLTM0VGCXUVWGxp
Ax64+jrbQaXq1A5YQzTwTCFGoXah9TY81IyQQeJzk5dp312TAGlw0aG0iq7r
Tpay7TBHls3FjwJtQFa8wUaaHGtKydtfkJoV/rV5fQDIWYVXMOCKzenVb1+9
0SrLDcjjIX67/0/PB1rQzlmYHX6jmTlvWy46FPzYkOdg1xZ1DtNwSAaNCWR9
YcKa9pa6+Ce5EqTTn3rnIzFkuUiRZeHznhH3/svl6kqmLoHsFEk0iJuHHbVy
/3mr0R7UlGASQXzQNTKbRdhCnUn3sGEnNQFumcmWFrGcM4/eWTkWZdvbNuxa
vVwyIjarHVJbbIZPHWa/XcbzI0uSGgPphIRRCIXZ/U1VQhaBWNaj8zjnWpF+
sLSZ6uFNCXAanB2I5DwGItKiHLR1LG8PRLEDA5t3ImVzI81UK58GyGEZRQvA
ABaj0jXspE1rPuGZir3zFoL4xKTQaExBLiHdK9VS0l9NewJgRRjT4TdAdplj
/D2Ua4oCdAouP1T4FxAk7fDp0MMODiU4UNkPZiMWJO6TEKEhfX1V/zttMprg
aIX2i38ai5/ko29XjhOtS1XfENFDxW/Mic2GXIZ4srB85r3L7rWuUa+XEiuw
TYo7WxKOTGYe7n818dzYntRenAnkY+tns0oLycvqJUIIId7iEfT9xWlnE3fm
9VAD6Cu+T0fffWpc0Phyze++6n2vRN2zmbnXLa2lyzub04LL3K86G6h6Fr8q
kJF85VQEYaDkZ8HaWjpiS1JoGHnrkoBI6X1G24MhtT5n/Fgb5xhc/5ZqJwWD
tRuhfTR0nbemCrdRLF1V9wGxD9wyYwdPl+mx2jlSdX84tjsaACTYLInv0AeG
mEG6FeZ6RW24qHuOZTzLL6D4X+/pkrErdkLvY3GxSUYcOxVxLf1OqcgC1JOh
e4J0aoWVdAPc6qGKN5j2BQWofzd+YlNFJZqhUy3G8a9riPnpz5Yr3QpO7PMA
0kiQf5Tzwu7Ony5zW8YT9EV47n86K6bi3MSFcm8qIZCjgCgSweUDml3yhrqE
KzqyyJyyTl9HcqL16qWW1PD1bEqA7ILMtUKU7NfKGzYue4eO7sYK15TxSDMY
mXDFHZHarsXczkcd2Qv3lw9LP1UlUzMhthuDxPUp8xEgriwbVKoI57eHaOV0
vSA3uKrhdm9yEM7dL/UOczIRH7G7ZqW6UpKAd6R6wiNRmvlUQJBv4aYXkmPO
SwP6R1gb+PRcNO9quwn7CqQ0G9HTH86AwzGKi84BhqCk/3xY2GopcGecUWa3
h02+UGjmWD77f0oCSxIOQtZSNxUPnHmAsRaVqH0d6a16fLLeEtdZtHs2QRbR
sKEQ09TfH1htimvWtw9l3gfR1PEoY/F2cKDNntPs1SVAyda/61wLbkXFZr9y
2tU/MSKUJF2ywbq992GJpLKNj4dQ9lvx7i5TdoiN08VW8fOv2a93d0x6sLZb
ITPevjq5PhibHlPTSqnYI/dUeLQCSef8NGjKI/gZ4URmi4yGu0Bt4IKamt6H
mfRMM67eAgFGZmC/C4lIYcKpQwG8ir4EeqMZBbGb1Z3F/eI614iQ8nSwh9Gh
QeC+4Ap7eRlksYMltehiTvO4bdrZbQQI1Br/VWDyRKIRsWMBBir0HUo8YfAa
uKyy5/7lkzibsGu869QYtIP6H/wWsi8JUSVmsafLd5W05xPKPUYeqbi2CLam
pfrQcuPizNo0WRfMUHEwPDWo3TvdDVrOQk1fsea2vIyQbKFr12eTVd+6ciWG
zuGTWsxGoFazoFk0MP/0TZQdwHsSG0KnchBeh8dGc6Fi2ZM9ZhbEUbv4XLIv
wN0j244VMbRGS1Yzs5kGsfjRze7wxuGFBvDl3/91A2PQu13DC03wHBHaj/zj
62ASohkPtm1YVd1ycWH4eQywudYILcctkcqc+EDkeyF0AqA5977vcinfUNLR
2KY7ywE6MFJKeRt5/nBqw41lyZWSExuBBluHJFVu3wCvODdj5lLI5TrTZCnp
77HyGjDMmuWwtPXq2KRvxG/6H29f7U/UMYjeQJV/3StqjZ1XtZAoKFBs6RdM
AvICyCWdmrW6GQ+GzgUaliHr3WUtYk+wqiBCNKsSfV7qF4KZ+kHdwnS8VDLU
H1R3ZAmT/tIhYw5O1gSLWjUdpJlGAxW1HWpJnTkXKSI23/plZHGq8/GSxNks
oCxxF95dIgnqrdU0NbuLL0XjSGXEw+bzseDKfVeyIpheyC4lDQiDtNtOgpdB
XU2rzopBr56oMjNUK5t4BH1P0SOSRSFxU3my+L0uIvgol3Arr9ekT1+eU0Lz
iMQVwlsZh/1TXJ/0h7KXbkcNK9TMv+MjSUssok2HYoYzMd5vVUU+5CcOe2Nz
D6t0MRLM7GLKHyWefW//aRjCcAc9zyHZ9Fp+ZJmptiJbQ2Itcmv7KUdVJYqV
9umU9yBbTdlpswyzP93uwpzRQSSM8WMAJk0vQfjyXGuySUQQZgRnXCsReNHG
FM4T3Hn+JALW2L7WLqFa7Zhs+U8+eJojDYjmWNM/mvxvIpCX6IiqYwgacUoZ
2pK8oRj6rNyXa0BGdpGEGjNvXXaLqCrGwb6UNzU5XCH7p8h3Num74X0KY+Oo
+aa1Huz1l9Ake+QGvQYNUwQIWgVCO8d450lYSA8S4GZdNiR8VW3IOcjMWmuP
Dyjple/L8E9AObp5R/T59oXDnMm6bOaCTy9J8KXWfYntXxkv/LiGG5aAizfo
qQWQLuECkPJtXw4p8C4zj8W0eeVDp9tONAg08zYS+Q3INC0QW/aY4E+1KXpF
w0aTxQumHSRiE122txUOEWpFFTZhtcTfQgDzVctvKbxUGLy7fdlroMdcyMu7
40aLLWr2lHq2OJiYyW/uaeUn9rFZ5owkE0deaMY0BF17D9/RqmdVWsZP96PA
32F/noBvVHmd/xBpU1uwDl+umL4wrG4D39Po3zUM35plFXca1GxLs67g8vv1
ueNdWtCug6c5u7DE+ofxEupvjJ4qKL5KMQzm4jR8xjKCXfdFT7ebkMu7ozZP
B4r0fYDF/LpMuGcZahwpMfS6fpjx/MfYA7543B16EoOTp0gHJVeaGOGHXUMo
SQSsrrKo/PmtP9yPbIAJT5Pf5QDSkjKxjd+O7D6kcDrAT/UXC8S2lz0gz3QL
V8VTRwk5g650R+I0SLyAn0mn2aV/+noQhSa1UiVGMNfueI/ARJFMgwa0XoVh
odLBiuwLBuesrGFT/lZgGZD8R4ReHzXujrVpyX2EJUyi+fJmcQivifprEf/z
ado/vhTCiRRTc5KOAYsHLtEsm3B7leV2dVuoPUbV2L1Gc9T3lf9MD4j4c8kr
ZU3L7vzmB3C9WOv6gNcIHoEH4URKBgORnXzhE95emgpcAk4UySPU9S+NG1rN
9+I20KUOo8dHx0bxG8lw9oBBmFEnVfdG31gQZB7uRp2KsAf7vg/XYlaYWqgi
OHoVa4jwzsAWhTbtCarbFFC3BAvPlhSNotHgXwGHP+ZHEv4NfGuMckZEq2iO
eYhxiySWDKxW8ti40fvhRnDA6GhJy6xpHiwfSe5tuveQLhX9XYBKxsiDmend
ipOWnI++E7PQzCAt3iUl2UCmb2OFZUevbCAdkom18/djJEhJlYR/qTnkwIcl
hPW6EA7rrrtWAuPIJvu28virLsWFp/7rQDpmZCWx0cajQ3AACqI4otKzZzV5
c+5xZACATiv2NP2wet+puAgsmz6FBysdWuBVgWcXXH0nSSPJF1LAq8LZbUxY
Xmf+Y55pwYpElJM0j6u7pjFfU9yRXij7RLJsbg7kRX1FNAtQefqqTBR5FZZp
C9emo7DVxgvmA+ZCRLYzllsRgKyrhdUu55w+aOWWRpWNK0cb5iki7XORsbUe
PSbIigwgpQ+JnUUfwrPPREV02q2AefCOEntM/Js0g3jk7CkltgNhkl+BRUKt
o624sL82uJZlFR7m3P94yYPq6XR7NykxZRXKD8MD3fATGotuxFpAiyh8a1i4
zfI1rPIOtut2pzumqbXbD+BffTFCGUd+H9NwV5LzS0fSOCnOTHmSzuwIUVfn
NGbNycFUOJPIe+vHV9cNu00lEVogZBhyFcXI/X5jEMrA5+Jf2QwS2B5C2gJJ
L6w9Mlf+a9QE1WPeiFTJKBXRhj/kd3sLMqZHoMNtoDB/h3cAfhJKTBRF2J/3
sCI9Fk1xei7mQEkROPv99d4ZVQ7vjKTktjcTuZlakwhnf7+LrgDf3FqeYXeY
RQt7jfGpGbOO3UyglWJlvh+KevNx/fCK/ZCYURpGnC+sCUno0tbs3SME8IS+
pFqZdSEySGxntKRAiwdeAnErGamirE0CH1T5ISVHdHoYhvLS2GgJJQlHnufp
TeUX4wtvqmKWCO4eLw0NurEPEqEQTjNA0yh1w4dbAwK1rNgsCCt3F9+VBXkK
GlnmcPvv/160nyPGKD+15PTTATgK2snklBQsJ3pJatOAccIzvbznIMXLfzkG
Tj1xFYSIBTsfOKLpdwayk/g9DriDoI90W/VJnnD8zbeC7yTHZOjGqQzoJfgB
p6xciNACbZ4zKD7U6vkvPwEvJ8SINLaw3qNtVqApKSyXB0OMzkKYt6fTWJbo
kRDB5PYWkbKWOh4rxNdo3LCe9+pQ9dwmXi3lwo5UXDyV2S83WlILsgCB6Vou
xACJUkHqUUhbco2G6HIkk96Z6KSsikNFaqInAfWl9dOo8gbFOGdXnbTPVi/Q
qgC7Cez8OMbIqAjJi1UCWVJT0fu+wJvivJEigt2w3tVb82l9RoruGLNTz//n
rtpN36wn6bVo5eTYZ2JJxJ92UqRFV/OjpC70y3IA7JAPYyIkTG72xdxvnXV6
r+kh+gGg9CwFo+0H+m75CEURenHHiyqqMB0rnrXp6u3ZhLyxtwIFQpTDr432
xVH23y10/R1l51Z7iHFvH2DkksI9otR/dQfqlWmy7UDzNC643RZ07zbSdwFU
2Z28vTWkrJ3DUDJ/Ax6jMndS5np4ktXkPi+KEc4SuaG5xPnsHnYnhF0XOaz5
ZKNIxs6vvO4PkEBii9/x9xx4T6gIbwRoVTLIRPn2YNKrYk1jdxjz0gimouWe
J905pmlbRxf1saSlGIL+y6vUTWQQkK//FgLfI3dqPBBRs4P39OesuGGAuvG/
sQ61ItbSE2ZyCr+i/lpEm8XNpwRoEth1eY69p3lEjBewKSasoUTJPLAeVTIn
J7Lscie0nG0QROAq1j7FW2B7X9ZHDgQ8IOyfNesh9dOsTFrVTpRZwJHn7fj/
o6RLLX9CYs7QwXo8dVYal5dqjqvqBqpcPAmmSUmMWC0eMqK3aZktKfdm/v+n
capGbt76LV+zqky9lA2nAF9Ylow8mR5HObeV615CbC3sOxoQ5dP/4IEvIhUs
pQRj2NjZ3YUaCXlMZhYOJrhllBqdgX7ORS+tv5+RFiM2HYknP6uqW9icfPdx
wwp1I5jrV1T1SvmUl8nyVGVgeM5N8Ga4Ro0P6KQ7OrruKQZp5lAnn8hXcjub
SgStBwHy/vhnowzCF0nWTVaTM+BK4mYSlY7pvsv2gOcAXpmt9sA8QzZxP0Xf
8lXtWIlXjMfhvFL2ib+iBtrYSzzCn6dzWu4ru5y0SLR1BpwkaOd5t2zUzCmy
6ejGLBE7l8yoE+/D3BVkmtpncHMzpxpJp4JsJJCIV0CFps7AiL3sy6uQ3Jq2
4wF98Wx3hRWMs2cXkJcU7V5bdkOpspCMBfGM9FBfHA1QJEc9pbl/KWXuab05
pLqH0HW7J5QwGLc0lQNZj30ND2A2Xn9P8xuIUYsT8V9WnzWsZq4t9lzYv5Qy
nYEXTikB9jsgxWfAoy/mGW2ubr/kmyYqqZfTrarJ/OO32TjqVcJPAbu0f9xr
UvoWTb0s8pLJWeeOy6HtIuoZhcI1fOFeDZ5qDOIhJmCji0jrCn9RLjiX01XQ
gUqzGqtA857XJktarA4obkDplaRCNpRSrROXdO+9RYGwV4cS59fyehCjPxbz
/ZOaIYWk0qAlWicjXm9cwM5cJDmvCqDPepAbVMDIFeL8w4aqr6gzdawK5Ah8
BJtyXoSwpfPH1ZsTM1UM8T5mJCFxnABvjBpXyKpGz8P/7LNjE5MgcyVVq82X
5umyeApgOHuPPk6QFEogAbxKyUDF22gD+4bQGkzJ3xfgnpqcm9vk3aymRoLD
9doFYyFawwJl+nEZ3L+UK7Tbia/Erp1pSUf9f8u6HRbmqqmEblQPA+z3aeBk
U2N978hEVtbw8HK7VUECdDZigkuQ5bLg6sgvkHT/Z5CrBR3XaKecfe3bXXsb
+t8MeoEMT+mjA8qGr2IBAgQgdyHbfBuhMKgQSz3maYw/Y+oFGVt3fym0Zq5b
zdQmxiSkhd+9HactpnczDYe6GutjAOGRUs5ekPE4mP8slLWQyeqbFSwasE/H
skBIsT2vWjIaVkGUodTl45Z2U0Zub4Z8eAg1WCsVmHGZlEZNisItM+MdtCf4
+k9D+OSvrNU5UTXlijun6Sb28g23x7SNAqWafuGc/db772vRWie/2/HRK7vS
ZtsUKqU5xgRrCiKw7X4PMmnc/s+Ta9sZNv8Zz3sfUfHO0Ny4MDvom9OGCfx0
m/YZUZ3xlO0EcQa2VIsITP3OrVjFaIuT2yXriW1r2ypHEO8+ertapblIxm5u
BFZGOcjRAzjMKo47p45sLYalLeJj7GDXX3L9PdjFfrlJSWWrKAJfkSSzhDOc
IsE/VAUsFoVWL6MMtABe0qQgVPbLlf67i0kGX4m1U0k15fyY250387Ve/cmp
nGoR7TiJbU4Sn1MHV+yejehjEZoaqlc9+aTc/eJg29mrUTpUyd8cIzqCcl3M
9qYztBGj0vHTGjX9HoXUWOJUU2dIirFn5G9tOXpKsVAOvBA7rvApp92dpyel
7mXEHHRl/1iYmFBYmUQrbD+txMJ5veXj4fjqhPns6y9/0Frlfq1h8GE4iidN
cwuVZQbkB++lI6BFIE1ZYqWtq4uyEiAZOVdLGxklFW9AJTTg9D6d5IrJDooL
By/VHAJ7+awBcHumHWXe+QjJyJ8lfuLaFNTfGwJJ4wfB4ga9qU2VHCslEzxr
/v0FiQaVDUSKWxGrawOAhZeEKgexyNJSjNwrfO5Ps+grlBYRQjnNRI5Danha
FnPVdVx1Gcs7GOcyC/dak4AeWcqAvOyWJf9fihVC97+6AVSi14Zzyej0CFtg
rtp16+8A7wDPVURJpP2MdHGj2gM3BwScgEEWse7rRj1XJRkbcXJ1153Wrjw4
9afJjadlltvOTYtOL4oAcAGCsayyAA3/mncnCwBRLaNPZ8XREms6oHcxzquN
+vAc/prHwMS5mW/G7olX4thHXWXZaRFDLWlluMv0jcu13V6JKQ3xNfC99NQG
nQKBHGDaIDNRqiVjd+hGnxc2n90EVl0YNs9sFbz3Wt83ZDJyAl4ipTqx4LCs
yAU9kDnx1J85Zg03FRL8BRfFUCM5PC6itWg4jJbL5CYSiNXvpo+zF3nYJ1kC
MxykWq1QUsHaq1aS3sXHh2nAX/d8lPxTMEBJDhfxTJy+NJUJGy6JxMIS9BF3
XfDw+2QVWf0gTQUC5RgRZU4WNBrOdwl8/dB5VTTCUp0a3kmDM+Tcog5o4nUZ
BtbVT6VkgvADqMs3ikJJW2qzWnr0lBC/b3esRyTjQ2dP/AZ2U+FXkdd41kuL
PSuGyzonh+MDYCDHRdG64xQqaqgywFPSqpKgYWiO+QaEiW6qesCZaafhJNQD
7VZgx7/X4T99y4/cwXAaEmssqL9BbPzE8U6IT1oVxCazs67OtxYAiDzx74rS
c0Io0dHxGWehEnheAOO54n/2cf/odkEP4Y0KZRfug+q1xbS5/+G77HKvJaZD
2kcTkvX+1sS+rHB+zyfRySLr2AAAltNPzrYrpdm5/iJAnx+hPqNRpIx+vSJK
ZitnMVU3VR/YkAgmxBqTQD2qVNtSAgXt7lzb+ZW/Fy6xyecjYVik/jnw2JsW
zoWb5JoKHFKQcvHdRjae/pQf7+jbxgc1PP8pMr4C6QHEVkmWXbAzuu3zj+57
FJye1+/nrviwA3vLe2f0X7RxKzB071XqwJaXoBuhLaLQz/0z8dUw6+3utSis
Y0xtb1B4gBQ2++GstpT/mtKCLH/S3HNrimia7kMa7/esM0bCWaOyZFRPl76M
JjaBbSgcPU6ebMfdS7wq1dHsppOA8Q+AQcgQJBTIkWU44hmiPl6QeTsf6nW1
vcsg6dPFrl3T4QV3FInSBI7Ix0ywHko/bTPwXDwSsYHFc99g3Ut9P+LIcjct
mQQE0v4EkPFRcKWjrE/P/JK85KDRl4cs5wtNo5qQpwah5TRRHeqFlS6rAD/B
DZ8jySMFiM91A4VQZ2qc8VYpXcBsp+tdlaldRor8eU6qVMwMqIPZyO1qbR04
tOEjCMiaPjF/9eVhvKOpEm1RB3zyTfXSzup56ZAgEOmFFbIzGdsgkvxIu5Um
Jj1/58nHs/l5W0xbummc+qzOhp0j2nsMbXmzUr0qaZ8QGRIvsUgp+5LJFmfy
Up1Vb/UkGaaog678dvwih6NTP7PwTzM4qny3F7fhkv1MegC0B/qzBCMS5opj
DcFwI4EMd6wP646pc43Zinka17Fq+/5sVYYMYZPmBF3klrOw5ACwmnYIDDk2
6oXHWwm8Xd6n+TYCVeXCZkDX2CVpJYEMFLRWhI7k06xJStdBVUc7+/Pwp1KN
uKsHCZkPaMa51lZFyf7hQFZEtAt7bAzZ75M13LuPON3vCAzxTISWKO7q/hmw
PCpiSMI1b0KRhs39l5iovPjMp+4NvV4i6SFuN60szAZw05NT/SdcMRGxv41Y
OpAtjYc0neEdw+mGurkbyjix3oI9CoOqBqsPO2qo+w3p6ZMSOKcmNhgNKHGr
VsKPJsmWAGxhqQ1UZ7brlrI4s5zu6CNRqLWmUTbG9KUmTMGrzoLNMzeQXuzj
dQGptFthxWNBWm48nJBE+a4BeFKqpKKwW/vyTKprw6bFyqj9Mh375q+UZ3Ld
MTNN2hrXtXKkW3g7lAU4jHse/q6rsGFTrRKhYXosywcvIvv109i93d2FW5pe
n0DL4XW55WUpUQN7jXPdCN/q6UI3Neptr0u2z3YqMI+BeXuoSSpXE+dbRgvc
y4S+/pp86W4GILpljgaSrmlz7AURWrR42LGVwkvwFerQZIpm9AJ3V4xoGbtW
uJrgTvdgGQzNHx5aHFuH6/uKR5NJ/CdcCB2j5r7/WH9l9aEHlYMktKselGOu
jWMrbEk/5oGyb+NSZqU7CB4Etg0/8lLjeTBbqOvYiXnX0nF4R5RAqqhu6VTl
7JHHHkK6kqoGuENr1iQbu9e5/QDAN6QcE8C0BWu3A79SOEcnPM02JgN4f/l1
FhDQokVy+1vFqoYiPh/yFTaGpAg+5e5FuL6KLWW0vWUb3Tfk9sG2+x0Jv1CU
WUpXqY0tydPsiEPKn8TjM+OhG8rlU8mb0Kv/aj+PA2bwBTXsP4A2Llj/2q3/
jslilXg683zyJD2RGX64+HtVECYmgGmAogtbd+nqoCke3IJvZqcT4fjRJqht
L9Rnyc8zJCWQYCqfFVZCrstov6o2SLtkWF1T4qddnITaBN6C48rrRG3VXoL3
xtgNE1usqmOQe54+uRj9iQeEuc2SbNzg/ITh3M89k6RJhUbfxYCjsLpooS3N
wbFnpn0B7XVX6isN6NBc2IWZ279HYb4X0edl1JvFfov/V8H5KkDEtJgMfXZO
dDPeQ8JZbd+snZia3k4CXUtbLSykdbWwqvpV0574kw2FL8igYVj0TtjQ9Vzf
50TEpgAChY3cOfLyyOmvYsYNUUQn+yCqomH/jP4vSQsB+OGxfYEE0Ws6ywSz
0Li7Z7wFtUCZClerwwKIlqauGHc+Rdz/lHX7Pf35g3FlEJlUfSuwSJRO8qqz
6tn9P1XvF2S6zldcD3XIJbJa+Vetbu8kjyzV7694RNE6/DKL9PtFrL1xP1ni
ZfxZjR6u6ZCiFefqSrFSCyvQj7/OsY1qcuR+nVeE9zwUk5f38/pTURP2pFZ0
J7VTN/SOI7RHz3mP8Vnt/V83iAgVapBGgZ3fx7j6P0a+wxls4+aAEIgWf8gd
OlP+z7m9IjZbSr822RJ6137BiNsycLZioPpv1F29DI23XVsRWF7t+RC8vMd1
A5ZVKttbiOKbP5sPlDjkGyVlUf/2mwW8JaJs59zipexKsc8ahhwbe96AAOXQ
4qUvMEUSYvtxVHne6+QzvRe9Gf8LWk0O/IXFguI6xCD3RDLbMFJJcAoudcUe
FHboFnx8XWhSyf2FcRUAJFJElKbWfidi6YvwiYyHaU8XrRCLWSjRnui4VTOt
CvZ7P+OA/gh0h/yybpeoxkbFIrPmTfSgFCnN39SM18llD4dOSJNrY42KBceY
CyUCRDcZnTdkhhuW2R7frzQP81TOv0/GOeLkviS7DJ5PZ4TQ6PJLkj6+tsuR
0+aYPkxxWTLMOYUTfUyGuoYiTA66skf+Gzt738SKLn2uf/ZvVnagUG6Ra2Fq
AhTXLVcVvfRAd/WK94EGHr1zQg6Z0kZqlXXK7pHtc5W7QvK6JsJJTW/qNzHB
dB14vax6l4/JDM2bGno3CXn+IwO0J1nikdmS1dkbfK2FcaJmOAgNHpttyET1
RiOdQDtokOOrEDvt5CffnC5tK+xT3mnWR/H7AB8tiwmYANKvHPQOGEqPhg8x
7ZcMigb2hdDLCVd7EB+Alhpg3ukaW+SyB/anHUtZ58MmP5lAg71HBTiYpS4A
e3A6SIWouDz2Y+mVk3phHT3rvhXE98A2fQNRCNR0DCuxBPUVI8SbkaEgNEFF
/F2dvC79NyDOm+Gfs1h7Zkls+kSERng5YPpndik26SsGKcffSFsRnAXb0QbD
WvuezsnNABbss35TUguWTkMnhqhrPpvfVkRdC6OHRygkcRcOmmfyzWEhdKuM
S+PGb4SOWg4mjW4yTOHDfC7nxF4CeiD9jATzSmKWumn5zcm/X0K+y8vQGSw9
xNo3thjAOm8SYl/vIikrB3V6ia6bSJQZO1kkUmMUxbuxHtjBlrnMZEXeWxCh
XU1vykyIvZKktYVFpg8/niZo0AmPnKZCAEmQ1KC2RrygDuiWGpnnA/BoYXSo
VdSzureE9ZXEp8tFxtRrQQOo8NeZSjMlPvlWbIaAk8lOp/MGSjgFO1N02FnQ
2Bnzyz94deuVzwrYjgG6bESGnOf4y124mMAC9xbtdLhfJLGtm3TD23qIdKzU
m3SUAhdp6+YO789sTy/E836Y9rakuh4WhWDuot1elTcpWutEyZYHx/n0JPeL
m7s+bqxeI6wIBi8/uTk3uhlF2P8fp7rLKA5FW2o5gmceJ4Xti5rcWBUQgOha
xjxj+8CmxajbyW7i92MDwbnD9nKfjYqs3Tx/Jv/t6TgYeTMGGLpq2Jjy5BLa
6AMgkm0gdQMx0UPW3V1WGaJkaLHQhRkxqdGDOOjB/AwYyPOb5BanBnS08rLk
hQ7jN1sB8hELYWPUENjj+TS+aUl8S/W6EYmFTECi3Dvx8UOIg/uKrxoa/RJ2
wO+TWMguI74xcthykX6nTOUHijHhmhO3g4dKyE9/JHJ1MkAQvihUYARjISC5
HbVidSpXV4X4uf20DWbHYOGF2OO1Z7F7xN60Jz7rKEUl1Bqjt9QnDl50iQjo
US3ruunGuHkBo3iGZh2+sitbjMMIDFN/6MJxoTL0fn4ILeDo+6IjvzYiqYQL
ysg/HZ9/k6yT+5Grjco2uMBOFZ3n0hU18G5UTiaf1LLGnDPKnxORlDn08wOv
uecMPnnDHy4HEwxXuRozrXeQqJ5JYWAfoqBT+LzED5nKKeYxEhkP+WDtnyh9
463s63GZbkpEPnEIh/3mJR2CBwESYdYDH2e3cRBJOXOdyzdyf6dzdpHilT3V
f429SvrVNTsMTMRBdS0rxZADacC2ZqFRL8GXNzHU2ZYN8SrmzTACQxBQDG8e
hHg6wzsZXV/3GESBPB4eAWd6U5vZ+Xh82yDH8j95KBOjRdjxTArmMtHwsmz+
72E4mHUXajy99BcaajnJLdqhUqCaeAZYPtoJbfGtGp2x9i2OMWlZw0M+Jlf5
AEVeWAFJnak83Y+QUSaviQcgNYHI253SsnH3lHtv4QZ+DTaAm55vk4Ubk1h7
m6U+039jGHvxhNJGcUOhKcqPhHQfGoBSHrRyKGG4OIOSNpOnxowNyXdztyft
HZXO7jlSsUH6qTIP9/TNU77g36ElLxjGyWYzlmmWS5890YD5IVyUto77I24z
agWsqHhRD6PwPXg7DCyU9FUk76XziSWiUkVT76T3NdVpJ869efb43RfWrHbl
3hotRzPQD2DGwfoO/2jzAbI/m8D0rqr8xJ7E5b6Ut43+1Fd62tG0huFZjBDg
aKciav8WWY7qk9aVzZIF8WYEkQmTVi+P36nSfxsEA5Q/EZKfmir3uaSuimfO
4gJt8xUpfsh1hUpMLu5W+CZgbh/3bh3qvLRDDWel7xEGouhZXUF8MbgNafJN
TqziUP0QuskAojywSwrKbSq1mfykpDRRl4egrpidX22gchHk2RxKEv9NEvSL
oCfaLpD7RvVl+H2bqDXxBZFdHzKbIOv/3Egm8LENF2jbJhpuvYHOoObab0lv
9l6xOJVoLIx6WTpDuMrsIAeEig9EloRJtDqtd5001TSb5EEfgC6yRY2q0rBU
vxC+Bg70Wv2fHfEvdY6Z78fANP6BxwogkafzG3sZ18xm7GGSQRIHmp3r/83I
IUdDigEwrOlsPaiAdqlwI54F9aN/S0LqMtcvLapXXxf8N8o9SPT61/S08Zjt
hZb+SoMsywXTtuxpWitlcyWulRnhV0Oos9oK7tJuPJEOCELchi5QHujxfNjz
KujzPjbOde2F6u/UGNG0PZ2sBBmF6iurhBiLVXakj3P3N4NM27+QKLz/fUmy
jOi8lLCBiwE2/lHKxl9CfdD0aAK0wbHKoJCtrUldBu5M7jRmwiuqzmo+FRWW
6nXba+bHROjLHYnqC6d+SdD07Iz6nO7f50V7jSLrUgt+V1JnyI93QYfPdln4
zgbREsGxzHCfWs2BIa2JH7sCXXDWGBI888kfrs5ymRpAtYfvEvTt1AJig7hX
3v5qHw7bXmF0ofdiwZ4F3cC0KHF4o0dGiE0B5MjLQOpaIc7aHaAo6GRFKaQd
q1Wqn0RJYlnvlJsTK5YKkwhcwAFGB7MA8Mk/wYROPCLvJonolW7EEGlGNp0D
h29tPci9vyCgIpZ1yPIhrlFp3RvIwT2W6j8Rl/9xcmqSPlQOvp7whDLwOFUi
grTJJiq+mHgrzdHx1p9XT2sTFu7QoFgIjo66OslUNLPuDz1MwtaLA/3/Eu0h
QQpRssCis8puEaXYW/ZPDsjG8LIrrHWiYhHhVNvKRt36hkDiaDXe17y/Jcgb
MkvPJUzhklSqxyY87IKpqqCejPXH1UVaPw0erdi+ni6K4nEvOQRuA7zt0TL5
6cB1ylC00xhW+TS7TVE8/72UCQWrbxoFL79fMbGLNB9+4YJRY5dK5xGhkmiJ
WUhdKFU6fBfboXT1kLGiEqV7qbo1rCZywvPV73GCsl4/fb0RFKYqE9BJstkN
09YblBuSFM0TE2b86GeG/K8EDdK/OFfLAQDSTWa6n9ygIDgYPVB4B2b917hJ
fsMvSL9IE2O2x7nOeX8dbsk4VMN7rdIeOMNW8UTNMo2/w2EhfPLrCuF2w2ER
rf5z9WX8vZZe4rE4F4jp4RP1kfWhrrfRwmkEUAdLvPlqK62Ik/bSExkpisUn
K59QSPP+FzTpxe5P1xSM1ZWiqCcFMBSiomhSa3GuCgvwj14UyZq2luokCuhc
MS5FUEnczzBxhSB++3V2F63nssE1Qeir5+MfLhK2E5BKhFwDYWVjAltNtPJt
A89HEmYYFZI2dDfPt6vWyl9+PAnA0wkMguRQO9RSOBw1ZCj9Le8+cDh9B/ul
IieuYDReMX6ubVwizRpc0pRYol9KWs8v5TowZ2+SAYWvOfkGsDuoHmfoTrnT
BPwlr8AcxKkYovCFtaZYnscQzynfe7r7f8HKQXszPPgRelzZxSFnuFP0jTb2
A9nlr+UV7VQx3AkT2J350hv32gaeWfpn3Vu+qT4ExYA4emmFGzw7wgdimXfx
ZXJrZas3HPD/X6yemQa5XH5a7NajsAbwiIBelF28OU9tpCS0yV8JvXGmA649
WbBf6enSdpXKeGHKek8deihwcoHx6RVCgUvXs6rpjU/yjxn01SOfTrOT/3x5
xvKw27vaJRt5fkAlmdK8UgbgPo8HhE52VdQPS0s9WHLkX/5zpkVwgZudRLBD
hwKIVDiXy5HgTabsfa2CcAPtJkinT/+cr2FW2wLcmKvLDh2F2N4fqSA6qmG+
/Ik0l5tJkGYghhIfApP5v4l0SjiEBljbX9YmaCuV6S6I05OXmJ7m93goMNXt
fds61xj/OF4bnVohyKLtQeOjYQBI818QN8+FhsAb2A5dUNueF9zcuVTDvAb0
gwvBg6VGDr9d7t2llFAFeoxzb1uJ0/ezsKab0LGeyr4jMO7IKC9EbVvoFEqU
cbzS+AaOTCG4vy2nAM5outGUKjUXza5qaA5ZWrq568zcxLd5Iw8BxeR57+mi
24JfKbV7U4f/g356hM0+6yL5vzhwpSTMs/I2I08UQhR95ild8qa3lYO+ZbzP
d9cI1XfWegkUnhCqXtSIjDyVX9vdEUTiQ0aImxty/JdfrNAulevFgM4KZZCT
5qf3PIoC31CU7S3RIw8BpUosRZvIED1uDfeDcuSFdfWDBtI50SLdSwt/3cIs
buKhFHLPHwjx6ZvDj4bOCnN2akXYy5d86C4uvPKGSoXVqRvhil4+bxPA7vxC
bd+qj+NwU+h2Gq5h6qLOJUp1se7jkouJgLWeXoTKcsTtd/kND4MsPn92ymtl
uZHsX1/B7oInZT2YioydWhRaI8cn8kqqIXpmTSLrbE0yKXbbC6ChxJujtfxY
XM0+t41BqOJ+wRJ5iJwmdjZ75lLP8pPPpMu3o32MyrD0fV0r2Q/Dgb9yawpl
hdqfRbNiZ4n+sR0PH3XkyrQnVF6VPMP6wPf8ILlhu4F+WT6ydx1MpSO2hHCM
m3h/GXEFKqkBY+pcG/yRIobnGe3Zg8hPGpL5eeXrDMVnQNXthqIE+tzCD276
KoeytzXmNgsjOW/JaynkpLdaz+BGC26ker5zXSSx7cQzz3morUDy0LtiwUNZ
yFcncBDBdZnpg5dSF3qZlZ3gM7E/BR9Aoa823gsVCY0aAxzm/t2zE0JbvHpH
Zsd41rT+QtRhVxfq2kzYv380lMbO8El+cA5Yaq4vfQEyS6WwK14EGGSMTYwF
AFQMz3Q6TdctT6ZaR8HsGMP6oo9xT1LmEzazEoHKyd6csIjCvvpkJz2yKUqe
Z/iMacChdPGZlJdtrQBbpHi8f0kuemuVVFUt4BpCUaIZCXMwQhQ89Fb2nD/b
DPAQzfytOhD0pOBZNLtMiU5+iylrEDN+actKKo9LiUw6WloP7qETyduc7ult
Ke9DMO1qxBdDDpMV3foXjG7Drbe8R5WvG9DcLMb/OmmBpBS8ld4/btSiNULW
BQXeGzfbdxpYx6Ys1QteWu53xAu8h5+XHibXlyH0OMkrR+f6Tl1uD8+VIIh8
ipUoA//IJCxPG+7rrqW8wpy/2fUEYyBj9EpryP/KvItRG+mtidZQykpKhFv4
i0FA8aVRdhmcKSFcMuS97ukBFA8rUyvGvNv7l5OezDXa7AT1H1o1xEj8zUa/
b0CbotifGqHtmIJynj3KZCgmtGOfZtL5NHh8bDiE0+tSAl90x8lLRZ0YiJ2t
DSO4Z8zwzYIc8t2KAJKW18iUYMSLh2RqjQlAsiom/DpvI15KoxtsvAWAAwf9
9T/Blj5xQ3SXusyeyjvEhQTNnJbHFhUeOgyCyHVQbFamnu5ABC65qML9lSgc
xKrlI6sdHr7avqpoTYYdBl44XfbsSq8vFir6/AOwyLDyDd7uG23giQ90RIIo
08ng1gt++IkhNnDJgapOZio2PtvYmVZU4vgvJBAdkXIhg0otV4/92+04WC4l
vNSwbW7HeQFvIkaNmKt+w945FRwNpADSbP3erNT3rMC59lkUaGU06mpL3ooj
ImJB1En02ioU4SbXSa3NZpmQ6M6KArORtnJnfCrhN8uiNL5NdvqCJ3nD72qE
grbhaht5hEtbsQftMoOFa+1pc+KQGt9f3fbeKNdUbCpBGiqjzOqgbo2QdsW0
bn4v5LzPTb1F76MX9WdB/A/+QN0UE2pW/u8eH36/tJlnVF/Si+N+n3yey0gs
C9WlhH1jhaCu6Qac/c6wkzBmOo6JhV8fJ0MVNNX6NamOlJVKzdkn8YhGTJO3
MeplYnZtCdfRHsd5CE6/INdFnTHPRv+5aX/2F/Z43knpxeRdC8cNuGyWSXDz
6lUeHfZzlY8xmuY6gwHLWV/N4FFSJcGdTtJrZZX9vQPr6XVM8RQqfNK/3oyg
DVkAxp8HNqGNm6AYsuKYpq6tTuYLeN03XqtPjRZz+D7W9qw05v7FQ0zHgs8W
MckXEVcv0E8s60yp+rkbH8bScNR4GFbQVE8JdFtjk6s+bMR8sBpOuRKimC/N
7cLeEs9zuZg4SCMb2IHK/Yv6gsZJ9qNU1bt7nhsQSfp8ZVAiJL7994nJ1VJx
LiwGK/K+hvWRPyUOfkuBDSsjLgr8+zGES+/hMb9Ex6PzVmFPRzmQjOCR5dL5
fkWzGeGdQIFEvlHXhe9ZBW8vkhDIj8FD9D3C0PB6fCSpnQg4ra6Q6xwhVqlT
JSewznWGw0q5tvvSq7F+AT7TE9vhsA+EU1dITrm1LgUBSMyzUJ3XEIQx7Wm9
mw9dJasmIKEQzAxwa4uRvC0KEA73xLbx+8CixFTFkPn2YnJ0pEiPrpRMDyCa
gufZal33NVOuZ8HYF2IF6m5EUrKIa+xj9dMdKhWDdJTTmqfl3wHagG4vZmsK
I2APCx0ya5pk+1+FgdiP2xhomufWKqeKCu6UgGqoxlXa12h72rbDKeBw8Fsj
WYIiuWjiWMhEKrMXbuWcwnl6AhazusJd5F/HSrfBDpC3fRM3zvUYgqS6Xai1
HvwWZ5Tmt1CFaH/1UMcVPvi331mc6Hau6aUODuHvyd1GeglVBFIMSz94Pqro
cZTqAH1XsKf/B+EieRl9elX74gEUlqvunEX4Y5cSK3myDstwc3KZ9h50jMiY
KAddCGk3hoaU3JfkClUj1Hgw8nkfnnMKR2g/YsHM4mriyUV6YjU/7PBkYjTc
OdtT16azHOj4Vm5OTI7wp0+8/5aC2kgqVBXx9gHIoqB7vCfayR6q4ewaeyGd
aBdgBV6CLwpMMxdsvIduEEgtsk5hM/BpfjXWYlZlDykutQgjpE79/LS0RFce
7/kvyc5S7ZmV2gnMhit17pQQug3iCRAyagev5BVZPu5AS/OUPvz212fQ+PUk
3T/22HWeDKokd5ffsuunyy+G2iui6DDjwxa/I0gAMjz+aD48S/p04ZfWLjY4
ReR/jpKN5ey2TFIVC2wLQdB5S/sZyBNglo3ip0bpYw/0XVh9JgWkX6WvlO2B
bOSPYzg4HPY5EAS53uMk02eh+x8IUCqGg5YbCU3vUHcXlaNrVGBJyJ4ovk62
1iaxflMEsSM9qXZiWLv09J537cWDD4/AV0rhmJgRJbRYAdQy327CgKlVvVxZ
5gsOqlDybo1iqzMA1TzMH5s82JyDFj53QrCNCu9pjKBC3X8rFdF4EpAfPlPz
O3qGrkxByMnJUkQ6JbGFuB48CI/kBc62oXms90PU28YwtRNxgAujVX1Ur+c/
L3Q/t4VgAGZWdD2Hz1SAQ3Tnhr0x8sTY5XNAzGvCMWzZ3SdS4PCpdhqfUkFQ
Namr03Syg8f/Tk5fGlnEcDKaMz9UDl8WK9Qw+VIGy8zN9jQlIu2mOAHUBc1+
xZYADbsh7AU7yuT1QpmQt/pOaXFb9KcIdp5ahyfWIIqyitSGKU7YLXqQ8lFp
FQJ4D/Zquvn/uN27Sd4qrsuVJIKAsCx7DtmwI5a4rYrTpOhvoa0qB+fbqNai
BXGS7rmcPwyfE618gEKg2otuZ93RYTIii1Y74CjDePB/QygIkia8kbfhetcY
m1kj/pgVHuZ+2u34SvvD436L1YExTaJGY1FQgIRhTyH3llauq+SOrmzMyk0w
aPMQ1g4BI1Sc6nUDfB35aT152LJQxdJ/VzkxhLiBTDD213DE2M8Gg42trMIg
nrfUnUWXGLyAXrodiv8yQzOlSKFiaN1u4SjW64peuE50hzdjfzB3+7Clok+p
vKVwgpLpQfXqNc4kBBV/w5Kg6gonwmF+JQPIpctkagbCRDHv0lraCx2AF78C
hWFXx4R3tqX8oEFx0G/DZvVQJqTpD1Ec+rdHindRcZ7G7i3jxexqPhca63jB
llcFgts9WYIAeL1T1UMXnvY7Jl0FjuEt0PgQ/PxKlLbXPp2lTm2LFWEM32gD
Za+4YgdkQtUg6jaF3xMu5SAaPtZxdZ/o+rioKOPqjrmOyiXaaS9fjjSBvqXh
Xujd9bPebisCHuHOp+TEt873q0xH4FQ44XaAyU0tE7V4aShIAjlCi7KJn7d0
GhtN7tDLXdQ2AwH0UZ92eI5zd4aAWeGTnejW5M/jgOkFDWjKa1rVxuRm7f5t
ylMH+NZURTlbXB3H6NxG17hCPsyVpCK9Bg0XGkP2XSf5QNpf4NoHecUXoWsN
xeQ/b+x6r3QvAI6WRjfuXXg/WI0O2awW29CUirSawm2cS/AnYh52SiWQNNO7
Cr3B2FiMS6gys1NOdvdqPA/ExJgdzjRE+0lBwRYXCtjmAhSmtwFU4wf6QIf8
EU3lK819zx5Mqio0d5Yl7aJ+cAl+lHqBembm+VxOd8ZmMBFtCcDL6ITr81Tg
wjPv6gAUt8Iuo/AbyNKknaM3nZHXLy7Uykivg5fv7MDP1EOXuw28hX6KjZtU
SOPsRKcadxCLGx2yuSdVnIwHYdkQsoPylakUTvYGEoGUY8qU/uTZ1etkvXXs
rGAi011G40t9IhLEheHZDn2l5Na4LVZn3GYgkv6cEZiB7LF1LLoYSvDFKi0c
ZqMd0gouET1slZuNqnrOjk9UW8EYLHBYaLONTc7YKHTGxsRsPXz19Iy11LVr
4ShCLFhxRcmqvggdYGcM72Eh8f1CN7RZwyRL8Lr9TWawit+k3e05YDzic7S2
ziW/jBDhtw/2+NGXIPW/U8MpC031hIYM5vJrGZuWcJc3TIt0rIlOlBpVaV60
QaGtuVs5UasdbGnHPNNxpgBRfppv+gYf1jebVtWO0JHKtxjGfNZ3IhWOQkVD
wW3NrfrrAUAjZSFwy/To7nu5ULjq7s/9LW4FOZWsHqrkvTlfcPK3hkW5crPL
kNZ1PKOE5g1tZRnd16NyWZoiuDuuYe2aAI+nXVuinKpVzyH9KtNJ59R7xKHs
vcliZ5mVL6/7NO6BYpn3OFSDwsdu888E9DWm4LekFaNb2H9C0sGvSXGkpyrT
eo0Rzv2lCrzgOjyWi6xX2EJ+yq1OkGJ1tdd4hxWjO+wkAPkMS3BwpiT7X8WG
5P2GD+7kWhyaxwfcZclwTZnPF3UOwCjzuVLE1XptfGE89tm52HDN1wwgEr00
icu6+dIA7ZTGWsvxt8+oyUzKkgwKVM0GopTO7gYeelAuXqCu9CqBc/aU3W7U
a7MSVJlNN4gnAC8WcIdQLdxVHT2QsBdXRL5G2gzJba2mi17ZSlG0F/nH/a08
YeNjamZSScI2YWWbRVMxlHx12DLH5EZ8PpEOFJxq6D/R8BMQWTr2OoCwGTDH
tnv+wrZ3VBFmA+AhN63ywJZLc7ym24ZkO6gBBsYzYzIA9jYl7LffZDhrzu1U
9eQgcxnZzJsjt2OTYbSb1R382UPQYNO47k1GItBAJR7QlUHP4dNll6OkaS53
5WcUPhbSIjEqu6LcWzdrNZo6VaqvV66PhLi7Pv3L1hBCrPBicrjtyYIWDutG
W4+f6VtEnpFGsd3fjXunL1ESphvpbWPhmtz4XK7SzQmKCDrDAFXBmz/cCelr
Fh0CnMzBzunYM32mlTiawM09MSytSOSakl6Dsu6gM51532hjskJZtFU7bFZX
5CN1YHKKw+4nR9RvUM8LBVbjwQjKW5rHD+1ySyOpGNupOCdyCOqLezBxGrEL
j9KG9YXTau0Ndpb5tyOamqpOwniZg7pCD0Mdcv0kcjkZoV3ljGASG/mFnVKr
FBgZEY/stg8ujGgt47wRZm7ZejGixh7BxKm+JIX0oKsXcimf9nafNcVI07k1
6qeoVJQ99pc65vldZD0Ar9uhhz3GP4RV0jmM/8vew2UlIemql4s4rtEz7AMl
UFnM4B+1WYo7dFMkQx24YuUbAwTsOpw/o3viSZYSySBDVfWT2MioirFJoCxT
p1uX7NxUAAU1t7Pk5YOYnIh2AhUPkf+ne3D0+PqUqP6I8P2BP8jkuGNB5Y2W
X1qxlyfGLpJlvebhP62PYtraVqfszs8tlRnZV4u1aSlaVb081UZjFriSwrav
c0KWcomKDyUMDa6lxKRMWh/zt3+ew/KIXoHqCVA0DyNAxj60n+954UMSpU9j
YtAyJH9vgFVE8FXfLyTHI3ZwTY1c1wFntIKfvyB5oL9maq0tLKdEiCnlwsfb
m2Pg8o/w12DtcqflBnQ5SSjyFjh1nIbsj3iY6FboD1z34r0K3WQE7H3tVfMc
RTXd2AxE18U5E5fkLP/vRbsktmvx9qpA/RtZJWn6lTsn748Z5Emd3EedLXFy
cVDXzEFsAw5j6TpTuDOZYdOrkgULL0i365Z+EFpEFJOLAYbBPfQ4vbVClEiC
ATdmTTx5bCthTr5fU2Iavk/ShFvQmpQQORJRI2FbeyhhXV/XMxDi6Wzqt8vs
FORlmll+FWiD5p6Q3tzTb5eqESMZyAt6Bo0XLEG6PkK8pgIqpK1OiRpXjiNJ
MkeQxBafRmJL8/dZlYeRpuSUCzWsMfW7lbSTi5hoI0zfdtT9OKbJO+vDfXlT
8egRllaZ/UvPxwf0ZcV1gZoTvB82D569k4Foty9bH7XQ+QUXLC7z0x5Qu1s+
lsPfECzH9kw/f3D4yBT/t2mVK1TJTgwEtCcGBwJpLzsXeF7knRKgA31gAZAA
WnyKGx13s2gbbXLcJs/GDnMY9RprfQNwi9hqWaMaWYjm/acm19fG2TboWzuW
jbIKq3iP49ZnWHoM5gfBDn1KhqmjdXBXnFj69AotNSyDznWNeIRkAm3V2HaB
qsJRhl3rL4Emd9zFAW1OGjXaL8p7YuyHnxDrryfLO6okyLIKR7Q2PW5aKoSV
TVSnewKaHDLyZM80e9rLkQ40/HNRK4XhSU8t0gAw4w3yil5civ2lbHSwNTiA
7sGeul04SSxALtRbYC6Re9BEZtCh9VwGSW5j57hWwQfF98VwmdZOjNY8aNLD
SKkdQa/WJBvzyyILr5WLq+BG3rxepw9IidI/lAHkR5+hcRWhezRVvNuOT1NT
GjBY6HSEVSl/SMSmj9l05DUIVqdrFZMbWaxpMQLkvf/SS369akA/+wMXZC2N
P0NoNFtaHLatPhV3iO7kvY8LtQN0EJO05PIRAg0uvvccIsw0HvuIZhSNS9mT
TTro13RkGslq7gu/iFSrERa7e1ZsSrEL6b0MZiZC+ywkQ5TIT+dgRCDvPxNb
M6MusIl0hrzi73LllYT+k8wkJwzP2vnlJPHOhxeLxLVIyjs+ONoO7N4P43iR
5Ya6hd7KXJGO6OpHPUzEs+3RTNlnDfUAluSiaRx+GTOu2fmy9ydBatZC9f9B
VIFhl781BhsIgX7xUSYH74lfI4F4IuEKv0x1L/yAe6pMfsJbOw1D82CUSnlQ
6CWxKe0RstmjCpcb+PblzGXTzFi0hT4Gg++tajF3mG8Lq6M0TVcPE2bZQNII
kBz80mKya99TQil02oyc8MqpIkQruKs7b6FORFSn/W3MM2ZUhwGafh7dqVn0
Mn6yGQAtWAQJZ4DC8wSpMD0/PXqlgAhHGJAJ6ja0JoTnsju/KwIU0786nhBO
uOqkYzsKCzFt0W8id6fxE4L0AbVJ1n5dvxud4f0N7zRGF9jlAmNxCajCl2Dx
ZnJrZjTF1OoYZynAJ1JgK4DR8fK5opgWsRmqK3FccJWUInlDaQL6Hbb746zB
MCa+YDasAzziDM4rNrvBHPVuwK8nuLyR32rrrfUneNFg2DymSwTQl1JS3omd
lYpKcdeHB3/ztvHstcfEjhup955qHhvJ3wuekAGwqgTLl+x6b9TpC3smFfpa
UmXbIzja8y9m01BsQgIDnWc2/5GckFIMWlG85r9Uj4wRyEgntocGbvGLmZcl
zU95ShXeD8Txmxl0a5PW4TKuu9iiS6ia7sl45tXTPX7rRQ2ezTneNXhMFCsc
/s8IYlKuk2D1ztg3HYeb1tWXQcX3jy8Ot+zJF0O4UeOmDzfez+Yz2qcEdYpa
/Ct+VusB6yqmW/LwGVC0YRAbTHXRv+fxKR/l3718EELT2Ag0K5bXK3mIVJHJ
xpq7rjjHTTRQaD8LQv5JlHTLKWSCIuFvL2MIA4arANd243wCaRSbN5qxO9ea
6GzMycH/khbuJWPzUQOUNq1X9cnEncsaa09i/ibAfULF1IPT/Kz38xE9rg3t
7GdVGMj330yyhJ7tHD3NWsYF9hT62SZ2a9SpSLrJtK3eYFB3x91PjJapLqGM
7FVlKzU16xgpgvRS36Qwtmb4EkmcLpS5dYnAXaIHvBjSRZnT6yVS3ARVRlEd
vC+cOIdB1OkcZfeSvHuVRFFeguaNsEcCwBSb3Xsp/9XE2RGmBXNwawikhtx3
emTi2gR13cZ2kxTcD9z1K0nsdBvOdU0WIrm0I1IP0mtJyQxP7CIGJj3lnRy1
A82aXH4+nCn6Po0z+QZWZekY2LOWYpvMyHCK2cuHdEXiQNM7BnAZ0OVhaD4Y
xtu5dMXwPNpgq/aIScTGjKmdMYsTMzeoyNvJYIuDfOyTyF2HNjnV+rBbAafa
EusjaItkTXl1L2anMfuTV/4h/d6DasSbAfrzZATtnhpaCzsUiFC1TiwRknU7
RsozZq8eT7pX9GbBtAk68my/a2gZ3fzgmXmOnJVtHXdVSMDK8A0E/XlIkH3q
dUdB5gPJazwVE+tJxd4gELvLm6GO54u0QijV9Kqc0CvNb0vLC7eTtpnnrDJv
DanO+0Nff2ECfBjiIn83NmuQheqlQn9u2h6Y/U71NCLxAcFB8ZBeW4uhA6zW
ZGvqM8nH/hGmkrSNlT0QA/VImh5TdqRYA3TURzwpFdqHeqGyry4Tho4XMXcH
2ait+iB4ajQ7r5GjWOfB4dMkeNMw5tgFsyla/muLTk/4DAG/kyrWOipvNcbR
/SKOcuVbKqVDbwGSXScV4N1/wmWqMGufc0G8q7C6EBAp2XVOSf/2OFDpSrU1
Lt72BhQfxjwITnI65gk5MztpjbA2Y0oPUCO95ZJSABjdd+SKI+2yncjIS45k
hRdbcXhnD/H8UHB13lZBMNw+Et/vOZAb6t1CnMdB9dYP+vl4saMrNdvBPD1y
lWPq565A/giZjPAsjADA3s8aArllaBlL9fi2GbiM72Xcm8PqP7EuC9IGe3Ap
D+VzT2vlu5c/ZFXvrH6AlU6wTsbzEXRuewHjEJ5B35UuQYzEFtMI5oMyxlm0
b9BetXCaT+mNcph7HGMKKU6BNpdsuy3mD2ZxUr1e6N4sWP4GrgmbmA0Qv+jv
XYAXw6b/KnKtPTVdXgoVNO90q7cGBIc9jnHt9yWlkS+IWCE+3C7OVse0TScu
wZCeuXH3NWYyrJVJ4VGzoNfHqikOq31x4iLmAJ2YK4HmbZXb4N7buoyWYnAX
/uHPIiJ0m8KaZFcHjMiHGHz8Gve+EScFiES7gZPUN6ae8vBjKJSN5ZyVepdE
nlx1qDPUUW8z9BRDjOJskzvgbn7Ae/FbwSOldAP+wlAn3b9y0MDD+7MavBks
bSH2Ta86eDWZzN//IUHSCdVnzTCLm9I1uSYphkyaT7jm7lAZ1KYh/Ex+Edhd
W5E9S+pSjFyvCudKDYSXMX/dHHExeMp4V0PwL06DWZatdN3QmWmTYQLjMlbg
HYx1QyaCUwGLrH6RNEKaVbZlyLNrUsWGDxzGtgHXUIjFuBEevqmrHuQim8HU
mywWM+DlMJAkV3411CiBisNY9zep19xBIq9LI88kSfpAJML7cqYfKAdkURKS
DYPeUM4yzJiMVeMDbW/dT3HYHi+gHMiCr4z4TbIv8O+XGEvcFa8nKiB52YrT
vrsZrclX30DhVdAt8AJrAOj78nAx77Krx6yG6MwWqNg4Lg+PKmILR4CzENge
qqxNTTChBa10lotPHSVo5OIO1ftw+H+s6rP08gZ1p3/BK3sfevhSLdEcNF+H
CjWJHu+wsosANwfDKz1CLRw+7xCFqIHjfyo9RXHPZd2nPvftvJxkR4S0GVC9
QMpMf8gaPULhk7aOOtj7pzIQZ6Xw69PyafgyUlVX2pJ5D4KKTNqfXtgw4ccE
zMfgIe19TXpBUX2VL8IqEoNo96xkcXLF0RcdvGCidZduWI/CATF0PEFnKAvs
SXH3Rlu7LJb9ciIFdVOZltzrbKHs+SSyCcNQ3p6gOLr1nvGT4bC7M+aFKN/g
vR1SfeNXWCZ3XUQ98q8uhrNRpnb2yFF36f23Edrsr7ILBIC3Ip1cF+E3vuEY
ocgrNKiMDefBnxC0JZaoZAksC7l4PbNy4MG2aMc6Km6t30TAYGWASPnSzs7A
dlAvD1GUyfqu+KVna4riXMYw2W+c8JY1kmasx4vqVXy2M9Ye+pS81CpJg4aP
iE1qcIIAAPt3zahOI7nsTjahbEUM2ROy1nAn/nBdHi2FemJWF/Ay4F8PR3oj
9gfKTErHKEQO39FJrdYJaYiEqpW90NkIjrUi8qp4pVqYpXI0t5u5wSuhXNl6
ZNFGs6VlMHB5hxel968Eec1X1PtsIBpt0wnHgja3MhnMuPwKfkdJfow6MSKQ
oNVFQu00iHUlXvFKwtB1b1m66BvKOnS0RvPG+7EizUUu0WTZ6BFXltwHSzJi
Zo71VCE4h7zhhNWF+cf0YA1Fix2Qy7Q5PfQgkXFvshfgsbaAfT6mzit8FdEc
3lLe81k513c+OaRfbB9WzHz6m8PdRG/4QtKwWQs70nbUOulAnbHqJBQaph6X
zofsE3dMhFAxD9+SqHx3pFvjTbnutxR2sBd6QbY8sfrxFj75SmqE7KT2zjZv
C4lye/pVMfDse3C9t0RCF74RP6Qv85AHvkPp2csGQowD9jo7JYydxqd8EX3v
qGHMSaSVSBL6a3X0bRPge3JMgv1wCuCXoVQaX2aP1/HTvPTxteJRG8UQDAwV
x8gvCUgRVH3iBQ9+Ie6lopMX8KUMDaD7IZsA7klo471pzSizPqvtV0CZb2yl
2tqYobxKGSnWukmQBLwMqHPHyrj+qb4PMq7eaos/zIvJJYrIYbkX9PdKKe1K
QjsBrec9PSH6pqWsukli8rtWjAx4wp4x/++txhE7/dm2HrCxix+eUSUtt2tY
IF3p6jyPXj0+jnsF6AYkkije5DrpdCKxm2JGwMDQojMLfIbtEbQEYqiGNMcJ
poBJZugN1hKttYCVJmnYGKaWiO0vm/68LJ+8W5DNODhvrXOVCou/ZLy10Am6
ALjF/v1duIadkRONBVWN+tzQKYLO4jZnYqAUedRSPhW9qKH5O6g5uainu/cz
qbFV7BACEF06zxYpubgxS2QHXYxz2CRVOk/EpWbzs1kB1nYbqTgzjxPUWoOJ
kwp8PWwUwRzOzcQGuzQf5STHI3fZ6MiB1gH3WTcHN8p8skYM3+zjHdeFbgLw
ALVAK4Yhf+V/r900cEtXt2qbKS6n4MDXYLP9kFXm8icgpaPO8C4oMDInq+OP
kb3xa/MIWKkC/lcLkguY6YoS08bHQj8E8gp3Vkx5bY83hKxTp1sZhNDm3k3P
arFIDkmi83k4UZ3iSOhUUTfeH8F9CH6wlxkJfGUG37orWOQb+K60dqiskg6Q
hFw6C6GZWeH8abTqJRG2V3uYuFiMs8R3K0o5jVg8rV9oc8hyKfhyEeetM4HD
5vgIIKT6vptySR/nFUWNMZav0fFFpKVmKRJrbPqXkcDYDmPYxphpGnt7VXCx
d3bm9aX4pF9UXIT6rSqg4iVpI0YTmHWpD4yCCw7qxNSYn/Hn+2VWY0dms9D2
Ja50ANljrSWTocuhMXFdtBsx41zWbgjh9STx69KPkJ2nSXZ9h+rZHf3z0Unf
P19bPfWny4WB9BRrr690na/jHJ4Ue3p1N4PGgfBFTPKLjCH+8oaGg94rz6Nf
LeAZg+1+lVm3uIr4euk+EIjk5eGuUBT/kV9puqQTGBmunmGBxN66aNggYIbU
O2HN3QPq/l/hntn8BvKTCgoqfxOTCWJ7eF3KAEK4tzcGBdoxbQmgHq83ZE4p
QeAYeYkJKCHV52kn8CDFZtr/bPglUhk00+tiWeDkVtHY3aLnBsz0El0x164T
v7IL4CUCYK0zm3ngWffTxCPhU+eHj67AIvN5JlpdMB2Umby47mXfN/iLGob1
DuFHwAnXAUFt9I/INfldkY7McrY9AxdSrQWB8VuOtPz7DnpeugOqWMWyYoYy
s3nt1RNBuNAp+woXTZO33BzDF9h9bCXtGgG3IUDwshDGJ09n9CV2PlyWQN2H
7Gqp2bneuDVLffZqIwJojfPKNavV7t/UXBmCnjUGhVuKa6SiOFLhI8e3Gp+w
dGfycK0TV2Xq/heerakGWK3kTIwH/UBEVQIgRm/JntGnrcijk2/H2jmf60yI
2wTv2IsutOEDpP9vqVRACiWXQ3RfT2RdsvpWLxLZ94q9WYD6ErmF+Sek26YT
9g4cbL94D1W0AIiZw8P7RhSCjBV3oGvH/247TfgOj4+LGDATVbn/lT1FUUhD
/vxm4khbkUMrAJ6D79apUhVeP24sQyk6tfDP08a/ScqHU5TRdZxnkwxgBxIK
SFCZoPoyVRklulq8iaiUNza3gN4yb6mJ1NbbUI6/bv4Jr3BAozpaNo9dEBcP
gCKBgO8ayoRL4V2lp2Ru4vQ8legwaXhh6SLz9BRKPXYF8GB779YgmIv4bzxE
cnIt2bs2pGvAPSTl5QC7u+FNBwawVOOd4m2kngSj982QZd2llYQCX6Grk/80
b2cBZp2N67RpT5+x2lQMrEFVcI/fXvOEr85qwKkQRbOVCgEFeSqcUJuYRaWA
0a0fnorY/Yw5QmMFDdjDX7qHmAudkuliupDABS0EPLINK8A1hI28xrqHBsQJ
QpdSAMZgk2EirNxDF9JlwSFntI1q4nNiZuBD5JBgTVDDhfDsjHaXVq7B+P+0
V4qUqKHSxX6mZ9vQp6V0MH1wZ2ySny+9Z070Ia03MaqMv0ZUgVr51n2wTfjP
EOh0QF6czz4FWbWrbc7kusK5LaVBT2cduGh41+GLJ/k/4GwrlHgRWHJQtyUj
l+YaCqk/i/qDXimftmnW+GWObOo+y+Qqis+eaa5Vjd8HAYNMcSrnMLHOr9ce
o7moum/ZFLzqvMSHc0nEOfU1XS+NdUuDMvuUJVRJronuSsoPnq5yA8DvwPZk
lykVDuDDbvUEFrMHX17QHmezCnvN11Loc4Z8XN8aLKOvO5YB2Fj4GMGrxYvl
9mmsNxj7eEqQhTzNchydpKbEMmGkIOKXAg9NlQ6qrPH+7DV3VHJ76wMasi86
pfYjTllXglzNeIcLbxPo3EiANfOybPeALt+GN/RBXFSLYJXndejPnYAkWFxv
Da6KzFp1oeg4zI0qoK7HcXbC9y5SCog30Z2X27bziOYmpfrMbpbTqyomEjsl
JBvboqqYqbHuCLTwRf4n1IcBSh/BOSTIvthlICBSWYjQguQTSOiQjAKjQ+b6
nH/RRK/9dYK+8IULsKmdh/37chiw0opiPOGG2z/ldpMMYCtruqsHPbMIxhz/
CaOYZCpu9BgrQHQv3I01popDoLWpGdmd0blzaIhVycAouE7ola5Sig1SDhwt
PspX37hH7Ksrsz4VOhJrdaOm26/g+1lRZpahnJimoFMfm/7SlqOmmAL71sVZ
BGMbvz4/NXTAnhT4i+E5SxHSmbERj8P+UUoeDJKlf5R88sOrrQ1juKtdkaGr
U0+q55PV+e/poC15E+jlANbyhqQfHxz/FOd/u4iL2hkWWOHAzUjtorF2juxN
xEKE3SV1vHLv3M1/75B1rMbxlqK3OKiOnfxVM737KhSVq5pwQcSH0OX4P/lR
ni5BlO5s8fDgSG4r2pu3H3hfAgnqED/SA7uCHHTz0MLU3XIwOPSKyeTLAjsc
HQSq/dOs80ne5frmIGkvFazt5gGtEtx9ZIMaMy6HXqz79hMqDCp0PDqDLaNN
/HHrNyvXRAgxcw6WZ7KSN5lKt6KWddOfkbIvRRIzLxqPPWTzHEeHreuGjE1G
pBtqIN371A3+gSx/Z02356exK6LAmYw9+0Q+WZnVreDpR5dHb3gweq0eozUq
JOqDVb97PRiVq0yUyIDSX8rQQgyOIxk+uW6RlW4kBpZKMJRe9rp2Xe/3iOMS
QAP0Kj+f3bQcZFyQ46cme0g2O21zXES/9Sim0+u9PLrF2/znnamCXGyOldLa
tTsfk4rlt2wm1bLdEn50VqDlrIQKYh+qBHxkaLb+4+jDEOgtepebwNnd+Me9
8oWYXiy6nqw+FaTXszenRxK6IKZzWjm8ihKitCmx/UGllezcxc4m7EqGuP6P
SCnV9V0ZAWkKZ54YK+5hpzxs86mW/h61Fd5ZNBnfzFXGYlShiRIRRb1aXzI9
515NBSlJtjbIWJ2P/L6NTpleQR1mIe/Xavtomi9cnDK5THIx1LiweIMkF0JQ
NQpO3M78PpD8kCSP+S9gu/J5WfHLSK47SzaSmuFrPOlSsffBTDLX8HIQzE0e
pSG9/7c/iIVq86B7aw77dboZpl6DuykrcMMux6DcKfXYodIy/EPZs2AmG1h2
PZOwf9yg/ltduUHDzKmvVwAjMOEX5uPiYfcRLY1r2P8dq2LjzuocPERTTF49
yJvuseU+dP9sWskT7dESoXOBJhBZlmOLp6ACa2MQO+OmbN1aKJ8TYQ8X1wrT
FnHT85PJ2J2XTVXmzBx12uul7NE37LGUU8BN5YWVPFFbVL9YH6T74hxAGDbO
g5SvmL/0jJ3wfrYitwD3XsrthhT+XgKFhXoWjko20WASBLFXjaaU5lg6d2qX
eOzJcdgvZUTQztwfzOEXXhNS7tlHdjU321q37/UK7brVnqzG9EyERPAAqrTC
Xi/H0JQGAIH8jweQY5snMKayxo4s8PDukAZ6EBuRDcnRlvsgr2IFQdXnATWl
y4jVsfUz0aGYjwTULBn1RCdp19brZmDeau95si6l9tKkJo9OE9dUjoLSjEbS
hBa7w55EAfwdhJF4xBK+zgcXW9ydZ7Y08jcg4W8sAhqlEK9kRBCljaHf10wa
briaQPVR6TWdYkIKUhuwL+p71fuRO8PbEJzuLQuQ066/IRatt4cI2+E2yltO
ba8612fQj/b+DosbJInnL6J1VGaHCsshetWP0jNvs9llr7J7/4ySSJ2bsfPR
oWP3YBYOOOScML6KAXjMiFlbx8Mu06IJQVVfMRg8lV637lEgIQucs3epEV15
PtKdEWNS2Jt+GzHR6WOhUuLY4U6EYUoZm9UhsgjgqcTj93BnsJXsr0/du9rJ
n4+tbvCMCVUFBtgkDVdyp7LnLkjc0St/z/HOjqebOSPfUTCvaI81kNI0zGnZ
HgmS2xcbOkXS5D0Cf3bzu/ZPhHwIe8722+di5BCvRU+cK/uNXYo5Z8Ty1NYk
AmwE7pKccz9yACczoBzCQ+xPq62Nd9xlAHqarxleQm7M4S/IkjvXa34Vdw3p
h41BBkTEuhGP4CpyIvPL17cJZVG/gPaSEswOZrqeBHq929uwbxG7fGm1+9Dv
WSpr0Xk2tInFBoH1V+sB+IDioLFvxt4z19xvKz2a5c7i7Ck9Lgpm/JQNaH4a
jbY6LlfBTh30Ml9xKIMMN2VpZvkK1RxPTErlxonu9j/LSc5JyKb/Zq2GHrZz
lha6Jy9GW/OWmH84e99yXHTx1nuuaD98goYVlL5bQtgabUKT5CNpjJGoeIN5
r431du11FsUaM8WKO2Q1nO3PByPVLRwmcZ/1snHte/8x/ES7fL4bgMVVJZDV
fnWSsiRx3ZBGsmETjTiAUsFVUV/e7TpVFLx8YXk14/malR3VL4LFvflGefHA
A1GnojPSvAPnTQ9Mzsjlh29n3Bs12+fDP2jefehuurW19+H5ANU4ompIT3Yh
WJLv8zCgMQgjh6zUJ/fRDuVoINvvkl2f+GMbA8YWUOw+UyERXQZE1QpBeZfB
6SxctMgIILq4EkePVTL8pVIjJvcOcOYwz1JTWFFGzLE/gNueEBwWcgMqPwiw
HI3wHoJgUerTej9caHj9+KDDfcTM6zC4LwiB8HUK2V+h16I65BHBcLugAI+p
7obRrhLS/AwrgToayJ8UTGzImOOXPjo0sWcFc+lPopnhsOErFFnikA0soPfd
0FHn59ZpT7SnmgZFPf69Ju2Whi/Sjr1aBayXsIzcA63O1F80QCOvNvbYjA2H
mOopnBH98PfrlbIgv0abcnX135YCyJyPrrhRaBgPse9WKJE5H3CBSeEkKCbw
CiOa1R5B4NsjCoULf7AzabkRz0XDfEPVCZ83qzfd5CiaVNTtAuXkTlGqbuG0
AC2K0C6HC0q1pR5c3A/Lzyx+mj73uED7/U37ilZA6j9GpvmXlWzlqVW3wGrZ
EkCmfooNe8+4ThXSW+cPFNA6JX6UFOv6myEmr6D4+Hv77Ebw4tWfsYYQFGn7
VMT+RJO4Obn40gLOCMKv+Qo/wZdFre3QgLS24WP9Mu2p+S3po06wR6uG8KSN
RLA8IdYotFQhsGgrVe4reSO3E2MYs3psVt95m5WcwOyPu+3fCeh5vp6ukBtL
+fZchSBiU58r/eB1cLOps09nC2zbFf3ampxuvfQda0YcaUqZsqHbW1XV5GMm
AZMvO9J4dJac8FTQOFqjT4chCEPFW31VXt0ZLT8yZGjBQUvmew96hAWEsIdy
L1woOKQ4ccaBPHbWd/OWJThIFe0ECvt/OFUpKAhR5nU+9aHwkR5xkpAWbcQ9
ZqqW55H3D29IaHoW6eHwnuNpy0KiPUtRhuOhEG2kJRQtekunbSSD3jzOmrmq
vNi2ybpuexTTSrHMt5fFteMZBc2inwd+RyxtwrSpdw4rvcCODHM5uZ28Qmns
MqzkxUSAYGWxsEKJWAFEnwsCIfVqIse0zINLkzAq26zhoMoJ57z+u8ErXTgB
rM3lGCXMZBSH3+V8lUIY4mocIDiDgOcHuMIoc+dMh+q4jea2KJDlxte18hFu
I0n3Mqv9jn/DLws6mWzVpwDTaPeQ3Fpgv5hYMyIBRx6Ky85Z8M9uRWweWwkn
RVTpkygk4zpXGoDwO0FRJtwIt80iVJmAStL4/LNkYXkns8ykSicU2KkRg/Lz
dGXTLgquFeahke37+FZZ3HU6t/pNV8ydzW9U3FRB8AzjqL38xZSXXwaBgMpj
+JadvxfnwSbyHmZvbRMYRTwtJ5Hf+K+8zow/pUgXsNFc7YfF8GgHfmAYKRnA
N88JuSHd0Ql5AmlIGvP+au8JIVVQU1Px2+THZZaZFr1mcG7PhsvkdSfG/RCf
mkF+NyT3lJvyx3quslXA+5MoaMikYGTEcwMJL3L1LsTZOuAhlDCYYwdk10+T
brkP9qBHrzq6ffxk9w8ejrl6U9PSCaOOi3DWRQ9w+F8q5LWIiThkkqFPXauJ
3Wk6RVT9KH5qybmafKwmkWLnzk8JYBZ3etd1QNzhSjvKFloTguWFlc8OzMNf
o5gohYLk7mi2Vo+bqXZV4yEe2v6l/pHiaWMzfWZwTYkj8O3EMq8z13matbxr
ZzVHYnVZhB0yoXQdNLB6Mz/sWel4O+Ymqvr6H8AgVDOeD0a93MQC1tcrsv7J
qNopuFBK/ssCX4fTKS3aQBOR8Cjr5AjmLKVBfPN0GGmfCbPRjtjTAWOnh1PH
jbUtDaJz2h8jMMC4jrAcxYKJWwtQ4T6I/uasyooEgbkidl/TWSBTTyMFsi0+
UOK9yGX0kPaGLrGlL1hICIdQOKSMjGUB7jP0N1ZvoR+of0CwLpUuiStclKhb
kc49xUxkQW4MYkXKazIoShwWc9th0uTH3h5GUdZVs4/FXt8WJjjKvitBU8zB
+fyAvz8NGk7WGy+nscWbGgUS72/ZJgvRK9qnyJTMgEyVsULiZvyh/5M4QBSH
Eery6/+45BBJa8Fx3wxgzPjJy+2eacEQKy+myT7iqj1ZPsfu/mlNT4SsdYt6
O806R/3PRfGW1wX4JHSPQUW/WE/B4Zcz4cifMjhGX+pz+mLDVt3bRKfFblaJ
CbYynNgeTE4U+mFZYgB2hyF7vTgl8FV0n8GXL4mAt+fSZWcuSsPi4371L2M5
ZjzIK7X38hFf364U3nw6+MoZGIYH+DWkR0ZByO/pjqjaGzFGQxQOJ5mHaBp8
JoMmRARDuktSZP3AAlhws5PC6nWaR3lzAnGVeaRlvb8h2WBi/GqkFpY7VVfc
2Rugi4z6Nt4/7QMBnVSC2yw5IsGRIbzzDxphHnEBgUALTY95R2Y0po2sKQtV
KWSjFm0c3vaQIZaSh7Rl92Z8rXop/wivHj7hEV11rBxSkPW/otmUqnUk8cTw
CxVNFZQj3heFu6AWme5Z1VZ/3z75TwqzLAcDgOWftLgb0oVaoEdRMpCDyXH+
zPe8TSE6byc/P3odukyA+W6NK9HQGrWiiVkCwMqSv/R6Ocq933uDcGjA8GCf
8fjBxrHs0UwXqzXNe+O7uzYNpn9BDJGuC7q7jjpc4tOwPi/PzSmdV/tXSqck
3NSnrnu7kSdXVw5G2vw+wfltyJ7A8p91VLmcdFHroKW0u+dIo+c8u13EWDw6
7bN15VZ2xsJG2jz+h3tnyJxXLxAqDaVMfxYvedsNwSy6P9RJaIFxP7lHASuq
ZdpcE/Buv+ApxannvlIjPQS0pK6sHiqSn88dRQBCdR9hBRtJqS9xCKEd1dOA
3EaLtV8VocGbYW+HbSLRfn3s7q0lQBO5FYt70D4Z2+X3BvxIBKnw0v/PO8+1
JOUqJCjXuD8RiPPvogn48nns6DvO2ulFwBuwwzPDM6qxasU0zIs63UxD0b92
PUcfJW7lA9jWFM90/pXGFh7XOzMzBqcC5+FSN/U6ginKqNjx9cL1mV+130WL
71SL4hlptrNsMkt8o0TRrWxSrtWF2s3JfmvoH8EKmdPS6fER3qwGbaLI8pUr
gzDzGcHscAZzIUx7jUm/k6JByiRCYO+lD4IKRHU0wMTHufUXGRIu+jYcEcfE
eekmFLuscwb1+NQD9wU4020/ZvK3ELemI7ktuO0QoVsFBiiLU7P+NOQamSlX
5uELWQtOxS5w+7ywggwuQx5lT3K8CWs8QrV4CVesaLnpQ900nDc8U1Lb3ztM
Tfs4eGV1GqQAiidop4gM0gly7yDvbLVTe19ctBvNIfIjdJRMyJ/lA6Ls7n7I
NHyZlgHZzEi1lRMzqTYSvD++tUaFSvVs8UqaBoMs+h+dT4G969ekFBYlVi83
6ZPL0WXqgr+APpHHTfru+2HPk0g8RjZoMVYFxb70LHNHH0OnvUiLRdL2G1mv
wq5Axq0EadGj2qaozWCFNt58gnxb5IT70klVyGihGVZLK7B+qWV+CjQjiBgw
dN5Q5b9sPbm4uoTtBvpeaFwJRmKptZvuUmUucWulwoa3LYz78wpBELLZACk/
Ub3uoNcRy6GBWe0/8Xz4Au4IwFJSt5vkY/kFpH7TRCmEUDWL9A7K3vGAI+Ho
D/iBSn0z+/Gk6DAjo+LcZHcxj0n82VakiqJK6alj3/8ab4WCVvVOh+6Nu1EM
ei2hwgehMnTGf5lI2qNAM9A32Cr5gYdwVohMBZJoDotNvWnObHtYRwD0ZEoP
gwE3bQWcSR9ufy/zuY8wCY58xhNn0L/R8gHsCR/O44O1hPvKu/n3KOAqzE+5
/0vscckh/PP1009Nbw+u6EO2+n6eAgjeptpsSHr1ZCwBh40/MfVIIOA+3PTE
33U/Xs/P8GR4T652awREE/I5HRvTGD5TZ6j8KuhNRsal2t06Ixi3yPgT5rD4
4XzANBFFCQG+rWE49BFwCjbcYo/Bq8wQAhETT6dNWOp1wVs55Dvuz9cTbxwc
YfTefFwTFvafttvng6sspwNQOtX0YGCGZPFvJjbfjEQFy4n86vwfFiIrW3fN
X6O5dk1MGr1YoGtpSDNGzRZAZG2Im2G9Iv9KWtGA9A58v1Y5E8qcvUWWDIir
AHDfTFgxQ5FpsIGaNAdAKT0xJ1u4WspzXEMT7dBgVnT+DhEHz8FIS/gps8lM
wq4T0axp8rWUiGDPdB+5BxRoBwP4Vn6XqHJWDvB3qzA5dMiNaDKXvc2eHpVc
NcaFjN321HR1Plb/i/KMZmdB2HqpHfF1m8V44J99JrZQg8A/c5DIHtNQd2xE
lFpvTRZ8EyhNyhxPCKcOgUsDr1qxzhmIEUZZlNmEMrMmL9PFz+wn+eoDE28p
sQndY/2/hge0wquCsiDEUo8lPVQeQCdrjjUCk8hv54nf37pfKnGoYWjAQ59Z
TSkX+TBdkr5gCSNO0RusWPsOHwnmRVw/zOn0EC30PCUoHI9fWSMJ5SF6xdTQ
fjPS3Ds68RdJeLDmg1IrKewFCRiebxJ4sV23B1B8CLVB+YyUlLNiIRAK6A9M
Ixc/N0pcxYi1dcgKKU/pOK4xda1ccbbZzQLW/kCxU8GV6U4dDf6xNLNs/n4D
rP55zToPwwkERTTe87BqhnLL0zubBCDnr0uAGu1A3qd5JYq67rZUcLbcNddK
2X2dd4AFSeYpEbFHtveQW6wUJ5tnxz0EkFLXUs3NIZsXECnFkKeTpPZ9b1wY
SHjA4neL/knRVrxVfipycCIgnE5Twt8r1AX/s03ut8K3qfH82sm4lZx59rbO
Qkkil8ivRivkR3xktJ7CI1jlGaRRPwmMrlq6R5pZbhvmDoOt/kxgHqcoP0jJ
f7BYypc9iBGahMCBES4ih4iS4msoBdWH+6aByEGM1DyfJgngz5KhVCY7XeMH
knETHqlQrQsebIhl4pSMuk5Xouad5CGk9MOkWh879A3c1LdJTI5rKi4tKT9s
Z/T+DQviIQf4RqQYRPcu2Dx+At9vomV2bWO0TNKUHHUhqsEuw6MygajFB7xL
Uzju14BZnYi8f5AfdZru+5gRaJYnuQLTqaFuu8O14txuXyQNWuh7UBoAKXzd
x58QJSXJ+HicjExiME12qLYa0aXedbGKSWlNuvMp13bb7E7Zl3BDk6Am5OIQ
hJ7eQIYz+S/IIqMhoL5Z6c+DTI9qszKzEM4XzWXlOkwBgx10wrLmpFS4zRt0
96fxTTuJKoExL6m8OBz40B/3x6X1A8+gcL8vH/mh5LpohVdJ8U++Bw/YaTss
vQ64ngzO68MtIiUEbaBhA2DgfaAh2auVdTmgoATRrEVfVohuXfoC+Jxssp9L
pWLAhSe53IAmQDIGmxulKkHgmzb04Pyd8pxuJQfW81Ehk6JvqTclazJBzkD1
AC/0QdPMCfPcfHTbdIUAiy87r1hF48aHS1K6xM7AZ2gRM8a1aymI9CPwkyUN
uHeTYd025wBtR6V8PIeWIWhm8/U9T2CnKHXgjMKaxGs9Ugi3Ogvav2/7Zo1l
I/cEjdr+4cziVrAcqKrnEzefx++4tWqMIdP4Dni2o4diqcLJrd0NtlErNGch
GzsAjmYi31cgepMMp2uaF2lfZ1jwc4LEP1GAsOP2MwdF93zmUHUNIoXObZEH
mL/Qqbqk1Zb2hWn/kfLjLRL1rZEAgXbhlTtjpY3YA7/QuxOCqI8/grkHn1Zz
dBaZirShvH7Lf50LpJNfE8jAIaqYzu6/6ASzU1Fo1yj9gp3THYgFrL+sY2IL
5bGu1IcddNywZwEZUFf4dIPdZrVIYcAqdHuuNn2K7pk++iQFY7/lZbZg1GRU
TYvPwy0p0oScrV07j46cX1UF3iu7zYOKJyEYVTEyw2wCz64q427hsbbXgoAG
PpU17J3EeCg3DxtAyWjy1BP7ZFROsqyqcEoRxAeQlqGMAMSwuwsjGWSNvb3B
7ZVzthHwb2rCvPEom5DwIaTh+9VCzOHTOJE1V70EPFUp5U/bKk0D4V5pi4D1
CIDpmI8ebJ04mxFHe1nY1yb1+XPMhsLtBlXuKEVCgYzQ2vhFsuWdRgKzZmLH
BZVeJaXRlr787huDQhgDE76qgR5dgVstaIu71UwHZuhO0zwRaAtM1AILmUPU
7oORdwiaYyuWCab3yW91RojrWvgbK398ntRAI8IAdCqBeb6uuB52q4v4UTZQ
TLaBawNx5xKrC1O+N9bD3fqPg9VaserlP5agnsG287vEhzhZInU8VwGrO4iU
LPbm64Al0qE/mE7sLSrG8o6HaTi/iB87dML9eBPhOTn0O1aXeHGRz+05/f1e
ZR2yTKQOW9oCpfXJS7EljvJC4sWUYeIjwrW8KIBD/qZCnXCzneG5JKJ+jleu
OZ963QCLjDQAy+mJ8KHUfEl+KP6DE3+w1e7//yOHwc9nQqar0ocm/t5WK31X
c/ANAH6hB7cS1vtBjuPtrynY3qhYhjpEYQRXwvMaVAR5Y4r2eSQXPxHpJWqI
3KgeQq9yQHiKMD0YRpVZtFxEf8DSZb+RxLPNshD9mvA02hMDLgu/m7dYLn5p
FnBunimMGhMzQoxCuasqN1TBOaGDQ3p6wmmcNQwSkGLQudCx778lJr8Mc+2j
Y7bphBp3nsUvmgrjBOMpZfIdTiYi8n5hfa666U0U5gDMTAoL5eGixhxrQ9Cg
34EKGEO8xyJrwPqPvA2mgNrFEI2ySIYXk641g8g+8IwtFIVpz4RhuQMGhOhd
5vKDeZ2MPSDSa4iVs/RSW68iZW/nazVjk3m1kJINJ4Jn6XRrV9Y2kgwQcZLG
Pwku+3jahlhUPu1NV/NlZkHQYUHoOgyQYbOHQz1Hlhj63/D/mubZwU3p5QI9
/G+pg69tsknTumTY8tYRinPMoR7apbF2sv2kMqmYnSAlfpeNowkZv6ry6LqN
3GdEN1TLX4W9Atvd3hCDungbu9n1wbYMe44dbyn5WU359LDdCmxSammSyfer
q8HO8+/YsGs/9wfg+L3a7osq2k3KeO2aWiRtk+kxLpDPzpI2/IKCg+3B9ZsZ
TP8TAm/FA8ubiGjEPwqct4cx9wKOkhzrz5zVBrzL4Z0pLgOJkTlYHYkNcWOi
0VtvCxOsxkiCJWUlP7tHy0PC1+Y3LRgYBdFxNPBZHbmRlNt+VVAJDWGO3zzL
9TNN7b0HAQB9vuPlwcDgm8CHwAV4UvarByWAaorhqtHwwEQ5fvmhq/ZAhydE
ip1HIEW2+ytZlM+UwdZJiIohsuooyXVxlS0x2v5TrAM3+7d4jR0Dvor24oAs
rBtueg7J1q+dIwSWe9wJX3pelTa2AnayG1w/tSil+JvmMAFjjP2X1lLMR5a5
xQQtPK/vWnY1AWbyy4xAeUf88Q+SzQdp7WESQnlsH8ITG/I6DG15+5qviA3Z
r/g89XXlT+Ob2pl65WVZ5RwT/+W2MjXBoFAJn2XYu7t1NCpGvpmyruLsdBDA
gkMT3Wzd8SKZZDtohFD7t2RFeWHoMLMzt4oUxS97hwXYoBbaB8Pb5zAHZWQ4
6wKTlpYfL3ONLmqw0akejcoGCa10oq8sGDf9kwnPDZty7YIgQwJ8FgZaR74g
4dcH6yU+JTX/xFjHjSQWMWsQjG5titE6mLisVe9vRdYFxPIU42pKoSiN/ahn
mrnXWkt1fltOuPEDIdoiNaWHqEObgfJp1UyONqhs/kGI9OHIPG3j/Lo6ipRd
crjj7vde95Dws+bNaBtPanfVXOofggZSQpavZPRD3TSvE9HrGZXAHJ7wo799
pB2aDzPlWVo1/uzO1JLSmIe63dwxTyy820R66W+POWt0c9I/jiF9XI9HGMGx
tt5bqava514hX+XBvG/bRw8JW1x9SqtbGDRsmgHI/lP6CAHZb0KGbzbhjahs
GmTgT96R2FnJoUqdnliXXKyLxkI7ENllwfxwpT7YZbJ6W0sVpnJYDAFLzbAC
0JgT0SCu+jUCk5suZBBf6f1Fo2VzVjzJdPtPVEirlmmO1jppljgOqN+j7QXV
gbTTDMBOnB9qTFb4Tjnni2oYMjR8fZJ18qLW5V1cbr0H9AH6/j1GwpSX3xQJ
X1h4ZRTX3sb0hbOUoQ2QmEz/kEg6klfgChapIB/5O9miW0GkONRl1AqKOML8
HTi8n/mlTQ9BJ9qHEwQoLU4VP82aSNMc5DmcNGk9uhiSJiK1AV0feVKi0OXI
AerzvAes8ik06i72HiulUQEfHE9uPYxRzhKF3/FhaIU9Nzn1Sep1mVEfyj7Y
5HN0CR3SYnbl+Seih7tB6J7dyTzi5o3MtDcngvvxzEdpa6I3TAlKzGyag96F
kB0yQkrfJX9rbmwbAsfh1JRvrSUt25/S6ujtZcjYugQnMJTg2Emj7c1OB9Lh
ai8dzBjC7FT5uZDX5U31DxGUCshO1kRUyflxQG/YSCKHNAHWOg+p5AZaZ1d9
rdnZ+RGHtNhpeU55DLEnClMNoGnNuM8ayBjvvoVpZiINwcdChiUUiRndfrNP
m0c+K8tCPkM6rqH6WVprWk6SSZBHjxz23tdk2sXyzAk7jOR46tkLpbsdGsmx
76hrEcuOVmI0WRnbKRPXDHiW/gCHqlT+dqkM717vjO/mKh9sijlDOsdLOYuq
TnoJnzAsfrc6AZVD5NIppQzP8KY0rktVCrSQcyBU2mfdLp39PwnU4eZ+YF/x
UdLt0/hkhj3f6dZoc+QEr8XTP/tmEgCYAQPffkhRuTghGkjpxzgwGKPKYHSP
UD0guT53sc3mJuZ5jSNzW1/Ro8gwmqlb5EdNAT5hFb254yf0oNpGSrRnfJTm
3QR4YFNrJm7cn/zhYAf7L3oafcPEfqyOGS7KqKsah2Nu3U1TWefWOd+zmr5M
A9/Na7RqLnchWjMf/7O27EdLhQPRoqFMNMttdwF0BmFVWvFQq0mwuwbUHu08
H9H8F96Gm2APa60kI5zNyriHADu3iwZXG+3QyVZ6A0F0B8bgSDhTFqcUEa5h
15fXC3Mzww6JtKX9e4HePkp5x39TvhO0whgUQKKa4rgJsmZ9406Txe+LDO4/
eWcKwhCkDi4gXiHQK9Tp9y5w2Lhojy7WiqcZ9zGCduy/zwE+3yvAhYHCfVHu
MGxUzfFSfCTpubQcp80dvP+2erPO+1vEJoB52iQYYc7HNhdb4gYWqlE5oLHV
RCVXCkIftqhc+US9yCbj8Fq2RUbVn5IdnzQxMkJ+q41Fbj01CeTktjomHBam
YFsFQjnLwzlm0uggKcLWAdH3TkiNrRfNPEttwLAWv5OM+hrAWpEj3gky/fFc
P9YGULzN8Ah+qqBKMnlSPEA3z7JK/PQQITLFN5ii6Kswq8kRZUgDU7o3U+rx
52e/kzsKA5NW2dVFAuN+hcdOlPcYZhimQ3/NQ8Gz5niOkMBdc5DBmMmuVW7g
EVELhDzhERh4xOLYsSwzrE+COo6Q8aR/R1lB0Fg4nSMb/QDK5RwkqHjQmzFp
pPRFAmkKEwCuCWRM6l9ptRJuupU0CDARH4oSHHa3PJcb5uGoW+BXHFs9CxMp
poA/j43dudq5qLeRgRMHhUg46YFMDbwiRZ7azZPdgagrY2bB0GPfannHC5tN
bHtsQnprYa2x/uDsxUtx0vAUD5z+dg2Svpt1O2iKyjdpec0SimAkPXAhNw+6
kW0JXDIz0MhZc6kgb+gHY68PLPqCHEWkALwyckx+VyTtV4+AGY8siYypJMnR
6/9A8L56TK5vjTD28ii5YxQ/uPjAL3O5Ab+/wkZHsy+k5XVw33oh0aySTRpQ
rrsAWoMWdoc3dM6LILW8CXUvqKf4+eBnA26miBn3WAgwQkvnxDN16XyoCMGA
xK3X8R38N1f+WaU0ngHYYttb6Sa8N+vZv0O0F7XPdPFSCTy9bDHO2hdenIrD
jgwfyxw//dLfN4rwjjQFlWdynYZCZD/Q116VMM16/ZcV0UjWq0zHvlV2+B+M
VS+QCFPub92lxavzf2JFhi+o3ZEbr138tLBRJL71aRsSpqzCXQHADnoX0XxS
IpCRRj+7umwIHHQxtu+dvbJXr7p7k/cVZ9jkCu0SksZdU0+PS2A0sLgzWDZb
dO4xK2jmFiCeNm5HW7hBXZFJtPFpuXU5/8oSmoGoHy+R9zhWQv9sJfvmgslP
5MmCKuPVTO+ye7yjFQNXpLJVMGaBQgdkSaFtZLeZypZwwjlZzvrqqDxG9qU3
LyN/yXCIXheMs4RPIUdkhteF2sUHX00JQyLuFF0WTBOk5ORUC4Dn4Ecq3oT1
TC2z5AJkIWZurabwRVQb1741DboECdRv539IU96cjCnHDpEk2ibG5jM6oLuB
FpQPp0g9tzdzNw1rVb+Btw5sLHNheBkAgYVSdbl0dRYDfCjHdYIHSDxvl7Sy
Rwfrj8e7w+h3JESToxI1OA7KmP9o6UHLInA9S9pSivkdJlZsXQ9Mk516RVqz
cp52KKy55vC0q8AHlnvJqidk8F2kCOLNH+9KjjukyCK8kir3phMnVQ8t9LXm
Q75EpdvHWEVsyhEDCuvukKeldORnh/fUAjNXYmConlEj4po+OxrZqKBj/dgi
KLRhtT4zfXVIelt4TBkbmz368HLXHRArGKX0WzFaA2sw3LHx89oIcO7eLVMY
z9GK3ngpp8glkWdWR4XssoLBAuFSBLDeVoLJcGOnF1CWr+NRkaUWr1ffxWu0
Ju7g9NiAlF0rjH69u84zz6IXRIXMnnJtLQfUmZ6Vjl+FEofnOCYhRVhEgocq
se4XWcRi5EGA3r2duXpitTr0rk1+NJihpuBBvIqKxmjGMSefyoxIkvaZTUtV
Wvdk71DxYi55O9TexNZQxvSiu8krJtKBh6iM/UvEI/kHe8IZjZoqPMmOiq0B
iIfYpLNYJPCtuqZRXoIC7c6uXsFAJdPeRESssBcbJLc/zXkT2n4HnJ+IfNu6
3x2+EBZUfqGAI64fcS3naCFHeC42P8+Vwhjq4lF/zyaJptNY6CxcoeOut5KK
Nt+nRBIs3Ng/3WFzcXO+DjwrCEsfJaOYHtcEC8J+9xavw304N6qywIMrUF33
8GVzT0rkmaGt3n+YHTq6Wm9NSLxrQUkg78cBSVArUK3lcVaGHkf70L59MAN/
hhIbLiAWwjILl7U8U/tj93j67Bxdhli+cykguqGceRRVlcg9bWPm2TOcXfM9
8hk9OlZimEZTmQDqFuwgMo+J7zGoyAizZrtMwwfHuhIE6qkGClqtf3DsgykC
M4Y4GCOno3TcP6dd1CC3hEvd1c1ik/W+1kE8rfuzpxiDhkguyn6ddXzjZtcH
24rmTwQsSyLy6JcCB2eqzuv1H+HjflEdsdEMayK/AiuE//+e82aduuQNyocN
7Ub9mB5l3CRVkBAXFRF6haczOv5nTCu94AfjlOuSVisyGfl2YZLqZt9sc2f7
M+vlb9fMHGwCe8RtpKdCbRnMDxjYM9+iwdplbNOPE/tVnGfW0Qk0y+7XuXPW
GkH3zQBS8m5jJqlxs0M6Ln5OXVZQ0eb0tZpUpntNopc99NT6ZH4ixHQsxXmI
PXscka9Ga0Mx5+UyQNFfnCpsezkcy/HK+AKUrIGJYFJQAHh9I356FXqcSDnH
6iy3wfNSXSzbi1QDaGFcVRER/TU/NlAvJc14BOYd/WtPhWkM0aLZVVmQ7xwi
Pr9rRJzg+ocPdrJ61kMMRdHUkq8QGabGQscZ0TBmv1Q1h6j6DBr0MzS6xLRn
LzMavCRBikCHdXjBWGNJTIRdo/Iz1TelUsHwnUEHv69cESTMoFqtsGqpV+np
s6DW6tf4Mvrvnedpl3vFqXbkwkE9eIznqFTYmQG+ErA1IfWCAhPZX5KGbIue
X+WxLyzaJO/jzZrtz1bh7jnM/iUZ1FG5Cz/5fqgHlmr+ZA4SYUqeGLtqoSL1
idebkQQ3ud3Uux1tgRMm3FjeSFgLJuglbA3WmLJHTQVM0KMU1Z4W5Nz5je3m
SIED38nSV+lyUCXu9EZSdq2VgRrAUZY1ZW+clP9UUIOuwlTvabQrqzjHoLXx
H/60AZG+43bCG5sjswz4gxGfk8pSNTjxuSZI0XWQgchMlCh2csSVfRtTZeiX
ZLCvJpLICvGcw9wS31KBbAEYYa/bxym/rrOfSU/7D69wKDAzINrLBypku3KA
hS3iGSltpRXMT3qIxpFljlwQJVfk2/SLKHlgFsXSr+I91+bAUoikxgj75dYf
zEwHghNkRFqhBm1Lzr97hKoTU4/QnKUoazwR+GH2fOFydBDxcqpFCDa4GkXZ
oBMu0uKHvSeZMPs4yQ5i/++PoSRk/FhDq2X+5AcrbQiDfc6shWmDIw+yCi78
Hk4yaYMdgp7Hupx44vNtC4iEWcPljM/Juw3mfsfMq6S4IDnM5d3444l/QUAM
hXbXFrk2IQXV5u4wNbtlaiVW6gf3dM1qltgF93ohKEO2PuNYp4tLyYCjFzBU
Kj91KWhI9T8aJXj3j65UNbmJB+mE/OJvFzsdrDDokUkqZbhdq5VF08sppt5l
a3CIA1sEa94BD88Bji8Rw6JLtgEloEgbeQ5G78JaaPc4WxWh+0O34qOCIbWx
CsaTK4g9MOWordca/WwvEqlzqfZ7x7TpOeLrVcK3+9Qs99H8wcOHsWkJfVA1
3lnsFVPh95PKdxhZH0CUlNHptutrFw2ZZYDwOB9vJZXyl0OCF6jUI5OLPMG6
GAR9iBdF0sUHZ6EgWclNhJrxSzWpnwn71ivnLpnKyU1VzNWiGQtTCBe4oMF+
xp7AdJ02xy4IiyoSznb3TXfa4qHXRuM9NfIJsKuN8f9VWKITawelstJTux4d
31wJw6i3sCLoCrLOkpuWB75zcycsQ/rLvqaGB0sb4CBmxGTlZrGkdZfGBAfg
gP9mjbqII1Irg0wkjYJ+/tptOycZw8MGxvFU91h0aJpq31HdIPrjpBGADCn3
BIEjw3t8p+EglQ6jkQrezpy2A3i5IvEf6WST29sEAZF57jhRsicJpELXCBaC
oBu2zssbpOlBKKEXWvt+TZkXj++CUhL7Nur12+WU8ButV+AW325xhOSWDW9v
MMlIu0+STtfm+mc3d4PgBSMRemYngCkWdbpUZpUSJBFazBTQr4mOPbvHybFu
OqtD+M61U3yLCJvPYrZMh8EkQRNJ4R8HYMvRatxH/3AP6123FSAi6h/N3G5U
jL6MFP72uCvUDx23M3GjsKhL2Zutl4MjhT75K1M/dquUsXQMZnVL9TzAydiB
1WlfieConPxOZihy63dVxj/kqGdd47j66v9J3uK8eypWuTkSQ9XWiLiVmQx3
bE4zT8Pce/VaFIeqRvHAnUXGX47eaRPq1i6t1qPYglhVjhfHyqbHrD5Qt72U
sW4Poze7f8DRe24GraxNZnD1WWeN0Fq83E5Th+I/LVt5PAQD/1Q8Hr8/v0x0
LeRjyJrmm+q7ysiblWGR1S6XlYCo970OUadV5Q1h8xSlAT3jGJwgrlrLQjrh
J6x7aC5+d+3kCOIctNCRV2X64e7ME9EO9jmz3kZPwH5O/JcmXutF61ZR2X7h
AURxHsTca5R70sFLpHw4p42iUcrDojCyZRfMniD0ZJp9rvMimcEOQPwS/GWt
6E2IaKLGvU/jWAXs6GK4gmTIqc71yPyqP+WwX3FTjM171XTuD6LEqyxprBxd
euISsA4oce4WrRx/gJdhV5vT5vALC/2Hr9JN98lCsBcpR67NUhYRgWQQAIBR
c3qMJh/ZQzWQs2fJsYWtOxKxdRvq0fnSs72nLnqy5lHV6wFq5Yzv/nZ0eFHZ
x1yVVgeyhNFsfuSMcitFKAPU2WTtc0MFTykfErV+0ynp4avCdlYvzZNH5eJE
DFDxq8sxBAJQU08JjRH2zACjinGX6dbt3mBnloSIlEQVrbNxk6SnmM1rYCQl
9Yc7gtCiLNEuSjXbHjJrDUOhh8dKvLuphSYse1jjyH0oatnvETUKgkSCQxGb
oEQCcJwnES+IHMHf/EREJoNBC+629wf0CH/ObGZjcz4nk95+canBdhzkSCK0
UqW16sRPlJMm5SwCL6veJQfx8LEY3myOww98MFeyU69O4YzcYhmBQZQ3496j
+DNH7amnUWj2ejJ4sTeep3v6yksKlXex5FVPd0dGxNLt1ts4FbODfZ7gdRXr
sucfHFN1fHlp20h/fRSh4hAV64EnHnEBIVx4WSBppgtU0uVcTGx6ADVwLTta
BundLQV/0Sp/3BVFxjtJUfHhTNGA0dX2yAxe2g97YPOT7mu7M0dn2PvxeQDN
hB5JoQbvW+qDD4z2L5tD86XoFmueNNu52cV9gmHliig19/yNAlbPw0YIASLa
qDHP6jMJi2e4Pcci8tJ8eUFr3Mm6a7lnlS3LC8qozZVqeahpfsuRd03cvyy5
nXCFBOJNaAxQS9WvTkXVf9AYDveFSsu7CkNSEl/gg/HAuboVeEwZ/2WMJ0eE
RajF/TBOPRCisxLM/ms+giwk99VT3tfN4Ff3c0VwJ8+wO2zhj+DMgEVfdOcK
sVCgVACCeNSKsIGSRlqMUq9vqE+YBJUxiEZWsBtwEnk/ePWcdCSrQ6nIjdms
clOZXz/Ac5DfIqGnLl/knjaHhYMUg2nHKP0p3hNP71DWc9Uc/Rkmxsh3mJwR
wNPaLgNYPMgXnhcAsCagnJfwvT10Kk3ENSyBjYgR0TPSHwaf9zCVljvC/E34
GUloEexe6xbAW1ct6nW0+ggtikWS4PxT1FAr13U+aqPBJo8bo1PRzDXBIT5Q
7elzXpRrfWYo2VkKw4zoeipf0vm414vmVImIyV7IrD3kM80mOGLlu+zxn1d1
jHP/ni7T7FS7K6pakhnSOjMnPfY8uJbPaiVDEC65X4tai89/2SkNk+pKxIml
ThO9ROW4zl0ar0cGRwrHG5UOLtd608p/p8RLgwAItCJewp51E0UXQpArr8m0
Ceytxqi8hXWO5QaULfKr7YtVr6+A/PWEW6ogs+UCXA6sKc5Ubf++iLtUfrzJ
OdHJnymPqQWQ42bnRsDhPxRwwVLX0VFVzb3yZI1CvgFDe8wqv2s6LoYmT3sq
E5qhNrDlmLXGIfaxs3UamuvfLJ8i7K1W4k2RT/YNW+ltuVuPvWvIz++JS7Y1
5uNYaWV80l8RkYIh3u9pwEL+bnnfy1nh1ebkhKzJFdvpU7xkA6HyyCYfZGRx
OwgLQ7BjvQRJeBbNQzIUtiBtrcScnlOri+0WXP0d70NI9ASTyxc95bShwspC
wUb7wgtRyhi/tlEJir0RJe8hcJlpg8FQn+K1uz8uHN337ouqKNnsj8ws3I7J
2qG801IumHZGyo1pTWWt6fMVfHtVKkYBo07gtc/hQ4F7rvA503VYv7aPqOxj
WDf/SpVhRGvMeoUaosl8P/IXbdvjqMsI1LV41yn+UfwJrWzA37c5xlaHALhl
d2bw5wfywkykhiFoTR8HclXI3EQuSCSJJZysHDlMiGmDfwn2teaYoQggJLbu
xjw7yuwR6dGesHgLrbKSHmHCUE6V778KFYZn5z79IbgWHYpOPRMNUYwZcLyi
JX6vYyzAQsb38pNd6B0of1ePNa+HQZsxNO+dc4e2nXty8Yw1Mdbm5Vbzt6+8
IovAdNWHQ0wEM3nJxGjxbOTIFUpkI5s4QPnUFustoJ7VoWfl/sSGrgxfGGPb
JKvtum/uZkNyfPjuKkq4PZMkdXbhuUTZFwwWC+i4Ymta65S4Id0hpaUuSU9t
g++5gCLAmKwGNb6LIy3Zh2TGTYGXUa3XDCfEtNJR/eEz4SNbkMbuv6CyyFey
An80mbzh3Yy0bVahls5hlNLefMlSjlA5kUhP4JpbI9a3nYIX8BW/AEBHq5W9
A4ao3VRxW3wgV7daD+9U5ahf2WpHfcjzTruOBk2Uad50FMT+IQW7V0v+kILU
bUgl2yfWKao1CfGIPw8YElZqzYVJjtfSf+OSgH+19qeMl1KSwSJ89w4FOzHh
1BErwaxf6Zg8M7vmNvggEkegiC3tIVRFFEYup625ML/fX86mUTFW92TipSiC
HDN1Oz/0oTWSFKthZdwavVdnmJ4HDpLY3PE5encrd8p/+gkKK1qJDty9Qn4n
zJGkdKtefgWpupNLrbCpooB+W6EjNgNYAX9TfIL5YzS0Gvi8xrirmXWTNkXF
MjYqJkeEuELBvhE3yxQtuubbW/NpTTnQy9kR888uqDM57eAmiIpxwPQl/Wny
z+SKXJbI9JQ2Sh1lnmA+Ad3FKCUmyvVhl/Pr5KKfGCMRsGH8Z2Ub692qSq8y
uTioTsbNo61mOh2scO1O+Tdc1VttAbWK5GzuHF9MqK+bFY3qPMfcXVT+r/7Z
fOs15xzT5Kx4Fr8buQ/5a/DZFPxAvydoAerc9nKI1URAQORikfSh9PnhEcrC
xAHGggDC5aRn6aFm0C0bBQ827Da3y2pfajj4SWVnh/xTTjMYlVsLY8uAFKiw
jVwr2g+0IxC4TXmSCNscbS+zHwFiWAzie+Otjx+NHvr4vgQohNkZwYbzHaN4
f3ZInh3MbcdfhbWWgrZYDVadNBFviy1fLdxELI6eunFzvQwoRQYA+b4bVolj
c+jjhVUkaP5dKKQ9LGUXUiZHwWsvdHGTpv52bV3kB0M3rHGXgwxnPuAWmXox
ibBW9QD2+/YZ8KpuPiwwwtdYru2BpcA5rfrOS/UZNTBZ9ivkLNYLm9Jr+QUW
SVQkmJ/zAjBpdfkiybRU8F4KwwR2oBBbg+A7HgQrTdurzBjCoYgaTBDgR45Y
Pp/x5CMI8Uzx6o6j1nWVCKhogN7TIPDx9/JIYCUf6YqNFFUXAE5iHTLGhUzT
AublJh4qE9iBHcE7vdOiDMnmfA0c2QX3rZEHYUHOUHQVQFB4kEn4sfieRnM4
bkewpRWaYj9YRNMaErDJiEaevUsFQMtmYUsassBwYvd+1lzw3v6EF4OAo+Qr
CAY0gX54WLbElOIsA5SWh/DbK6p5XBJfXkP3y89/zX25Z46VVvvnzzAaQg5Y
LiwTa4judPNTwnYy8Ge7N1rA9ERXU72kmbeNXWcJd3x1G6NGLlEd3iVxz6T8
LNS07lgp0xmutzYFReuf5bCKHclvE2Ht+fyY2/XPhQehBt8V4FYihSyBRwtc
laF2A9VDLU+RC0XhznNfDqrETZa9pfAOhkVNTqGUWD8SVVXIdcwi+ZC+YPff
3f4OvTLIgB7XZxIHbEba966Un2RCH7MQV0ospy9u3yNh83Y6h27kc2nNNj10
xEX4YMofCXNkENM+NGUnc+mCHLiTvDx5L6nzJ1vHtt3YRIlfATPUq5xsvaet
l3WHvRweqfEY+zk3IYi95Htf/WyeWu4zjXk6t9rp7fdeM10JczNrIyBxqwZU
T4FT/Cn1Lba76KXXcrwDTp0O3d0GbfF5LHyexWGUeozUNSLsbbxtJHsRLoij
bzF5yRQZecBTdfsUcrBFXPuyNO+w80C/tFljXnNIb7N3pv9Fb7rlFnzZsxd2
Ty2gT/qwjCVpwfw6c6nrHuiINzVaIPkiUsWJluZzcE0VhbWTigWjadE2dzT6
rcyyHG/KeTShWkLd5n7uXLOqJCVD0fbxd5oTV/YavwA6WG2me0REU2zECv/j
JtUzODhehQzf0hUpWcsRb8i1007YPx0NpdQ/THYKyZPXFi9DBPRNLJF1RWpn
jAAvP7cnEG3U1RE/PjeZ0KDrpWIKvFd33mtB73lvt5w4zM+z6AhIZOLrw55L
kYv3pwzYjHZ2OuNvI48f1dUh4lhLJS9ZnrPkaUASs1E+Yl7+yFLKT+4Znjl7
f+NWtoU6LfkgH655d/WnrkECf5GOHEF2rnvyORApXemCTWnyfc7dyYzoJsKo
KpBMUom8Bk38oS56J4qbwa96iU5jiV90/FzEbCA31xfL5/8T4paRVAzgmFfe
mLyxZ7wyeDWwFYp+jvMZGKEFlDcF0hQHJHE6OY10aoJyAeQWE+3izuYq+l7d
wFbO+ExiyG7bZdfb267jkjHY6YNArN7CA2w7DWMcQCizyzXP4tjvaVFKYOmb
t9nkmlQeSufPwG97yNKHEZZvvasSixIRv7CSI2+sPgiE5pEgEOFNe8OMZG7y
Qz4BxmXMFkRYMGKtWkEbCOtapC3sF7fMLG0Rds7qREWIFgukhvLjFEUR/nNS
FHMeQt671GnHlFFE++JzT43wE+evdd8GrDaXBIN2D+L26GbBbabdS3PZDd5a
WCESyo3GcL8dBjMNToHYexvtxXoYx09gWau+c85oduaPCRU3wuxXdtzpYxr1
1IqdQMPapRs8zMLsnAHL/Q5LkB5L4y7Zxlww5bww4IkXi//fLY2EticMIGkj
VKLhsyLcVzo2TuZsGl1MtuKfvbg+o72N5P21uMqdNFFUXvu3JARnwsoQlHq/
asNbcswhhiP1ADQ7DrLiPnusxvu2KOAxEiWxe1it7cDTi7IN6VcTmHxM8X62
/LKMG93N2u0/cntX3I+2kdxXG5cXS7wWCnpch71k4I/yxpVBqGde9keEWXxo
a6l8V9Y8Fcip+IAV6/5BNkpDa8SAe26pc8yQi93sLFzkBGUAnAksNghlwLQS
xTtnG+qaqbuoSA973HxUBoE6w7fA+bt/fkhbTBcgFw8UUjC9akvKK8dwcAFo
nLtl4FvBYib234Rfm8P5717JDLmXg4qLL81N+auQnOmLdQhEkZ7uSSQY4o0F
bnDtcolCx6z7StVh67NlsR9A4ymODgEQ3+vhtVjaP86+/OEsXbFuN8puMOab
YXHTDmVj7Y1YvOgeVusBAstEVc6l3wDU22Hfq7rTPggfgnEY93B7GZaCLF9l
wo+jndpIJcAHC/oABharL83/F3Hg1BQYdJebGCzpJ5m4Z7Ndhoa+oReOjD1g
b1zB8Vlh5GZNyBTG/VfsBwUvp/kcxryFzHBEC6+AlIFZoJLxCHAj96crSrkF
43kumuRhdN+Kt6xooIeCbl9HCKqNtj+LhKcj0WB90p2xHQW4YoLAugu2g+bh
QC6QdRMgAtPkq038ZuUxh3ZZP06mmEUs3weVYgJ1tz9S8lTLRePJOt1uv40C
Ss4s/DeT6BUh9LsjNZVewtrbNXmBDnO9h/fhCMtRav0UkzkdJKjAJdR+mL9A
Y2LhNrpOIGmXN4aYhrhbmXNFdQjLmfXSRS43rfkNDrhcHo4Tr+y0N4VaTqVJ
CeJm4Stwix8Fa/MW7Vs0yxMpS88zK9+LVYaz1DDRws2ifiHJ9N4IWjsflV+H
SllSeJ8h8QmBHyvM6DdapmoP4uSjcJNou6DuR0X4cuCD0ZR8GAwFZH+DQ5ED
MMPKLYTI7FOhGkxuT7A2KpgnqtiTGsjECJGAsn9XOMbPwEBOSzEnkyECzIMt
XALwkRhYLhSzPdpxlmXIEiM8XKAvQiEhPGKLNLP17xQdqzjq2ZqZZqiNWECQ
m3sSoBuQJ9hAwj/KGqdQzdL58Yg2sl/iEYyaCWqDLSshbDFZq6XmvSf3r0ge
S43cPuBAFTZLyBUEvuCXWH/cU4WhnM0NpgI+nJi0xqomMMu0kfZpCghNDyFG
AphfXko3bXcRvKHlmxdpaTIIm4Q+K1lU8xgZZGnpJ1VNP9auITDKjZLk7Op6
UYuYFcp4k+tHhqKhpO8VQ9Khla+O4WWg5U0J+g4a47h29XHnbEmTKul2VOWv
TG+o5lK9qds0ho+f5hI33S0d0y/AmBCxPSQpq2lG9tunHK5DwvOItgidWyO1
hg/adf2J3bBLUSLi6Dk82zpRFZS74EfaZ9q5/AiAIoj1sDkJLrqYvQFiokb2
H087ryo7hk4Dlbk8NoJcLIoRdWiq+k3tebjUecp6w9eso+Omc8qzSyJEQ8+F
bV7Y6DbYMo7c68atTOAmOrOAxIhnZcIsP1qrgmVL24E4atFPgRg3RdAJIRfG
rox9NzyIlGn9ejRZXNknMKvcoJvbhLE7w+O0A4CeOov1B8bR0sOKwu6bmp75
EA54ueUd8zZkDv7TYeaFMFQ/inld9fgaP4yV7IB1tRQnug/VSVk5emyn7kCh
+DcEaDRn3A0VtyIY1U1j+SHmf0fGHlQHQFECy+8w80FhfnfR0m5yy9xTv1zL
7VjKYkEy10CUKFKLc2P1IGjkgFut2+ZK6PR5nxZe+GWsk1rm424AhzendSLD
IjE6Pcawg5Yogv7fkjzO+ZXKZ77qhXi5QYjcRI2IQ6fyr4T5BE+tNvaOomJw
B7m0V2xOEEjfkFJjqCSZ8KPK9aJfkpgT9datUa0twxXcaxbO+7tDhhniOvyI
1rEl8uLdC8d6XwRgVze9+uGsusgf3J+2tulYwKwPdCVlK3PjqUPx7NtjRgmN
scIFPVLme7sJVOUHqygjYOAFsaAx0lU3bkwjYn8neATk0OPxLy7qYP1y/fIj
eQrLU4MnOPnu4PhCm0o4aTInnz/l8szjk7jX0yvmM7ZhGSNyZQcJnnltbRMu
cYOGBsAJUX1IsraOjQVGrV53W4sG9qXfa5BL32piY3AIlpb4fcDlCqOTkIuS
j0C1RfN3JS4L1mqlKBfYl67M+HDLiOAB+OnhLxVVYZntWjWiyST0KIvOJCtP
n9LNfvITXcv/slqAqBGYpe1G1Nni5QUguQTPJJL1HsJzSwqsextRb7yI+Ka0
GNegrHNs6kOiFVKcizC+l5R3Erz3iWhiXPJDGHYy8dePbsMnGr7mp4Kp/Fbb
O5X6WjVhZDHM0zwwlEi55HBRAOc7NipC8Mk7RfQtxoh/VRpNn1DAgqW3hqSQ
rd5W4gptCt6idGZ2PqEzXmSRfgVz40KZ6DFjj9jsO2s6UMJprhdvZdHrKohf
yuKBEMZqgTuJVzzLx+5+bKy6UKzPf0zST0OYg1l3Rf0n79EJi+Lrp4jXLxQY
ErARuPSshWJRg/MRARjkJSTWUz96Fk+Sma/S/ywymMJNhrI/1vvtDAV9/lZf
3wHESJx9Og/Vjg71BbnX5pIDt85DGdUXNCYuCILAw8syqDCNdYnnHlY1VXQ1
zjAzPw8+0x/hWqsOEsjEjFVq+/oGLxTWcVhwE4Z890fmOh3fx+hdkEjSaCKY
IkumFRD5Ol+i1djudpqa7JLM6LXSYeQPl4csykncidRWv8ZFutU5S+r2OUZu
3Q3hqxgXn22Q6XOgeVVLANVb6pwie5OkziW0BH3JycRo8ENS71QP/J5gQy46
MZ1uMY+q8DN9BKT+iXaJp5dy2g3OgLDW1YmouYUlSmxTlZf37jE4HfXwDjHE
lcpM2EnmoayVwxELbv1177UX0s5daS3hR5ruGbtjVsTqdf1Fd1PKcO/i6bH3
IQv+VeCr6cPHeOoAiv/W65Px/wMx/Xv/XVe3UjytV8abeCSBWi1Yay3Egx3D
zvOVEAmoe3nHKd3OLEimQolO0nsiVz+jhpSNA4Ir8m7bPsO6GnzAwA/gUCLJ
DO1zrsr72TY1HaGtvVzfOg9OaTVBvJrU6knOVUDIxRQFrzaxYeRQquG498uu
Po5LYF4n2NC8vSjeVNFsJtOSZ2Q9vxalT/+uSaxp8Z9XM4xruqIEHC/g8vr2
96odohTpii0QqHBpONQZEHAUNEOdxr6NrarCthAo8gRBfVIfI7LPEnaEVoBw
HC9mnRfcbqb9zpAcRqT5zHLc+Wcf0yJm9UL7akGYervTvI8oTmRzKKWtZToF
n17QxdLHdq2jp6BOGot0/2Iv+oBldNZlwnkTy3pANj32ppW1Auq/jSaspXBr
7SnqTUKn0283aeyap+1E1FF9xVGYtTes2lMqAOw2IdBJNoifrQhxaqdHH3EP
RDGZeCuc9ESkQcAajZA3PgUIiUdpNqjDKjIKOt21nPv0M8Ht7hIuHxK3WX1N
CyY202irfibkcJ6Gr3ao94eQnjyCWKYlZ8905+cTZgCKfx8fJPBFTn8HMlIW
AM5XGKKU2ZaHZzt1PR32WmmQy87kwFcwHPs2i5bWG5c9GnNjocXfkid/r5Fm
mjezHBB0TXLC81EFWhwbEc9etIjzUkEjpyxrlAd6IJtgGl3IGUzwIeZTIOus
Hl0MmxqLnAe+UFpQrdlEPdFi7tUOHJppTgDh0Fr5TIANSRKJ9ZzAx34SrNBt
XRN/MQJiWbOiJ8yaoNQrApoRj+xFjz/x4kLTjECCPQv5QqxQZ5rhodnlEMMI
LljN0FW7T6n94RfHBGlcqJjsAa+sNztMII4zvDpW7dCbgd9HAjkCYOlzWQEa
0d2lwGRuAsE8CDFj6VVi4Pw0nQYBoLa7JK7+iOsa1NJmWHZn7qNI6ed9tAt1
lH4GMwKxToWzDCtOG7mKhR2y+0C1/sBSINiLU5i9wPNT/2NJNgkVQZAc6KHp
B/BOILMZ1b7oWBGK5sE10jho4Jz6CUNRWXzAd7cotRvePqAZTwPLiUY65m70
xAJ8nFpZ4asoLKlm36uvlNE6a3Pm1ysS2dnzwOruqiTYduUOMPzNxYDzMd6u
KHxfA2R7Tq7DGWEp+c1SBY2dB3Cyc9yQyDgwoGvGVYyjnVukQGu5t6PMBSUR
pgVTcCzVVdgixX0Xo8BzZdxsV3/6vInh8N5f2PHsS7PIQm5OTAET5U9rGrd3
Tw/rCrdjJdyK+PqtjOSbzQuuieymsIogjtpOzr5nTfiwLAOeL67n9YubcQON
LwdQvPCUmgrKZK+nYLhz2B586NdX8ZEMChlh1cNzpWMnH+iQRJMY1YRIDuYb
gMF9Sf+7jleBZSUxl0Z7ns7NNwERtDIWtsX/qXBjXzamirsNW2LBCpR6dn+w
m0GuKqP+aHjOTwlQTShZvfJ/q2xajET3UwVJELXk7xkz7krXPsL/KiIfGq6p
qwOxKaDek6PEeJaT79LR045EYHKJHCRxXB4fZ+dS1pEUMxSZdSrStrV8qpMn
iQSo3XqpRWKh6RjDOCSmgc0k5bkZCGdM3TF88ybFkNCfOhB0tIu6ABwN1DMI
WWMHzvKtEhfkeWLD3Vl4HPkhaK0JyDu/csllfpAiBi4vVXqbFuwpbw/ZOMtg
cbdbec+Oq1OkgmYiIOokdHPZU9J0tg2wAlMSev3W5g6IYgECh2KAwlX3Bbmf
ZLWReQHSoEBXYpvi5TB3A+45DuzSJ3Ewuvla96RP5kTYo0JsBstloc3IFTaq
u58mzQy/6BRqwTLT8dh+/X0lGdGVsFgCYBIeRGqZYUW9aVvMJWFYGOwKQevh
S+KR/Rd+I3H6BWPKewl9Tp/zSeoHTEN9MC2UOrTQgtHe/0M1mAbbcvjt5jsI
mJlwoRbQEW9QEFObsXMeydGbdTtDkbTaYl0wd2xVAsnxqe4Un071XwdnQ5dW
kESyiCcsZZh4AWKuttmYN8RPEU1iOD+vupgc1Z9r75YV7aelEJxpnq1Assh4
bKnfEcS2nE2WT7cNy20f6+tceE5XUns2AOQHJQVrBETxpv7XDgtE2Z8Mgz3u
Q1wHYM1tlh2kk3d8X9gOz28vdlutyevPZC+G5UPIgBDtQVLuF+ZaOhbVGqTa
RLW3VMqUi6Vqf7vIqbwMEM4TDuEnDQ4xNR8hm0AGgD1Xn6zurnnZWciJGpPV
PjJVsLZ40FqcL/PD/XU5u6jCVjMk8w91UDHUxAVPxW0rIWn4m13dtnlXYgLk
h8HCpS7Wh2rRbkBcIvJ8aWM9KsV+JqtbYphfCnqDt/AmDstQR8lC5MaDqYj3
igpUVe1nM0wBbB0oYV2nthD3RRYo9C67j/y7P1bEmTwEyu8Mv8Pae5yE5jTx
BZi0hEhtvDdeslHBliJlw1OygfAiXdhwpc1LnvyQ09TpBXEeGgtxKU1uAqGh
A++y/bIZpfcJfKzm10Wz0MbJxUxoLxa3k+Kzuq2CXVLvsOKZNoK+UNR1Mr+5
intZxc5GYNyBmh1BNYscTZM4TcUGM5Vnn79s3x5cLp/XSOO0eAw+OXdPNaMQ
yELi76f+TOcevUgV+KoqmcTHTYmZykODy698Uiavd8sdjVHcarZfUul1fO9S
Js40jx/+N/fmJHB8RtHy6i/ywPCXkhPBgP+K5AepAd2FTli+ShF1ZlAtAyni
OvTq/cykPwdCbtIquNxkv2QRNKsSQ+cRwgTfKn5reu5OjbWeAWBQMNSk8JVo
F4rNdqyNPXHmsnUXDQYd0RD6faQ+JADbr1xzADnicqg0wx9Sg/YHP2f5rhbu
NtY4G34fesU2YnNQt0h7dDnQlov8SjpiYtx1Y2HQ6KUNxVjPrXwQSFJW71ux
xTMyGevmmSDX7QF63eDIQ2yvlbFA0L2n5Wy0zaFGVS0NpVtT4/HIeCjENBuZ
1hPAsX/oaxkWmv1rXTzNj9XoH8p/E3l587i+JvoJH0GBrvw7voLDuVB/hAPP
CLUCgyRR7EQqaM6xaKOGdFf2n7gkM52wHkNznshR0lps0rAUgW+qiEGPT03K
hlUnHJHs+x6Jc2KtEKjP+DGoqOs2wb8H40cKBYL67qaf7SwHqud9icafqyxp
DXhEnSyNnXoVxQBUY5h/lY3wRhlt7PhzcsH+pB3ft9hZYO0xo/zkzkDo9wK9
rcnakRmcWVulF1U5LJEBYU2Om/CMMCnLb79AB+fAOztRZBMMpdBa5ioCFq89
d8wmXW1hJ8Ik8Hskq9t94iI61jvwiodsa1Q2eB0SH28t/rbGdVaTaRGgD2Cc
xd18waDX4pd7eh/SnTVIImSyahtD3gSuOQu52jnTh99gRkY1AMM0Rgu0KT/N
LUxeCI7+AdRMlYa7TrWTg+06w4LL/YpQ3SEkoh/ngsagMuEE9rCb9aULq3d8
5xfvyagJOYg2vm2XG43HSQe74xCSB1YOcOVKdNP2LB1Cn78IsshUun3MgHYl
Zkd6ELxZ6gmFAZePIlAjbEcLTS9+drdSdZUEda13P+gkvMASdAWWBj1guOKR
S0YNYMVt0SQgNEg6qb6QAgDP/nt/qoZ3ep88XHLUIjCur49c0Ie02R3avXxA
OyKFYjdNv5hcVPa3R1AR8GIgGnTTttSZZHJaIJmgARrl+m3xEwP+iBq+W9/9
rFEDDuoEzSocfnVGJ8HZ03V355OAZKyvfK3LF0WS2LoeLj1/yVxDxcNLm6HB
OZzpNYsjjFZeZtl+CCMeGCoN5I6Q8tOTYnazH20upE01bTPC+9lYZsQBmjNs
ZSJW1Z2sUZqFIbIxbBSEINXnzVtCuYQx0dsQnWrubewzzwlTdv2VZizF6vpC
TlYp7o4NAjGKYD9ZwoI0Xmf4BuVYzP5w2Ge2D6/4W3iuDvu2sIgjskXvSXfy
cSUZKAnkfFLWOZrB9hECpVH+/fEq0DqsTb4OShBWgCmw2BIBVkUchGcg1+2G
62injWB9ZztdsRoHYfbQ6b/wh7UKrB2P9VS88k/i+Hg1/OE+kCUBkaVXrYAZ
3TFpiHzrcpho905lw7FzlRSzroX7P5Fy5Gqg39tspM0YPWbpaotut8BcF8Sm
TM2Eru6mHwGSmRQWPHuhZnhNqSOcXTTSvFLQZq9dT52enkuJRJQI8etxFZ6S
o68o30NT4t9DX6ARCYLxXaGmHs2DUuOc4feRQDffk2nErTfXilzZ6xFqueqi
wordJJtp/SR9jhQZ5eWmXPyDFpct7ilRFQ2Es0dc55glgIkOZJ4St4vpAxgp
zEbi96is0WiQWJC4va+KWhRcaAebwECrJ0n7Oig0RBuRvh+m6KsyPic+SB93
38mxBD6+44IMGnQ8mAZwCV/02Rv7ImZSD4gVGEFVOXTxdsjfYQ5KkS9YlfaA
tdlpta1r9vQaw1fCkPGgqquhVnznQOgNx7EE0VAqcPnFcj9gWYF2ZJsLXIc/
Lj6QO7n3MWUlaAytNIu0f/CPuD72ha9bAGlbWSqZJCy5BUfm318gF6d6+3Av
NtgI2BLXBZTuNjS9Hoyy7w+OmolezJw7KMznURB+gx/nFnt7x9AI+o55tu5I
DNpDi7veMxsvho+rBcAvmIeEBZRSFPvNyZyWNKcDJc6PSfqJTPyf8f4UH0oK
W3MFMjPUmX0zLj0eGx8SvmSILEZVrTS6bc4mO5JjwCUaBZv4SZdQagPQh7CN
I5nR5SNAI1KHiIkikqK2I6reNk8DH0nphrXwQfMpT6AXPTbkXTO8nooy8JIl
Zq0XcOI4hLX/zcYyO3hj6EbzOA7cB1HSr0GSg96iilkBU13BXSKwCAL0kkV2
xUIl879ZkSXLATZfTm/NqkKIdpOogxsbCOcnz4isRRJk4kEQYpBV+UpS3shM
bQF4ASPiq+k2uTcEbEjQzHOxbAFg1C/n6HAuaUEgHQ8gsLEIVWQ1de36KoSZ
YbJfwtGNKB5Jpg3R56KzFWNO64giLU/Cx21eQpnF6Xx39MyHD0QAVxa7dP7B
wfx2I9Y1/P6kAE/sEuojUEWnWfogbxYmGXF6IjnUOPZpsrpqPbBhqxRG0xzm
sYJSTGOM2vPt8IxyEAoIJbAnD8Egrog75HKhD2s+S3+tREGUJddjWht4DIGs
CdZi4e8ieJVzTEOkYd1rzJQCzibQDu36yja6/XLElK6e4wmJPDfgpFWefIu4
s0DQTEPgnEnM5DDJ0GLCHgT3kaFbEGX9J89wT1z3FIN504YgebNtLM1D9D8Q
ZtKnNu9tZb3eLI0CczTxGIOHKDQq1owOua+Po8VQ3Jf22sDv78Wf9V/7jcZ1
lv9I44zJjjsqNHeAl6b1yn5/Ye3JzBTiNZG6OQnTB5w9nE45S67HLrzNv3Bn
Od0sYo89Oa5vzZQFm6qUPojw01D/fxsV4k0RAFnFXay32Kv+4qdD/MKsBCYr
lsQTiFh6c2Xs/1tuLrN7wnUSkxLPAdf6PBrOnovteWLRz1Qkk7qNfHgKNmvO
B8EGMTyafxgw32FCJgH/HLnMW0+cQkTj/mIgRxR966SBFbZEc8zRLXeCC4kJ
FMurUHnHqVz6b/mbtf7TxRVC4hBABHtbwIiXlqbVuN8fODil2a6n0jfrLBaj
BU/KIVamqHg+Hmt37V7BAm1izhlor4ByG9Mc5ILcYDLRUVZTOhm35fdXh42c
FK9hoizc0AQnMKenBGpHv9uXoIZLTf3fnlBBIVAwYUPpXPT6hm3XEYfDefc7
lS2v6bSrBUD5JZ85dAoIGe2aax4+o0cSCf33R0VhNMfxSUnZJEvdgnUHCW+2
kSkqrBBfMvJqSnbYcs0xcqOuKIsxf/jXuRzLiP15J1hR7AQJiByKJ5Zep9gH
08llsriG35kq+rQzz77AjYkv2K6TGVs5ahKi4D/Ykzg9zJj3qIStCw7FOYZj
bZ5MVYyIIhisD5LF7viuEGaww7Melim7QJfYLgawJWGPsVbF7Dj2/qVU71Mg
PjloLN6TH0JbSnNI3fsZ+I6ckt4pdFCsRv0y8eRSvg+FJoUUVjM7dTWBmHI1
QgvEr4qO37H8LXPFrWKnSVxAx+MkVQCobDztJpCMmITkjWBTvKS4S/XBvowa
elgClk5mkqH8K6O9Be2l6zW2RjT1HqjDJrqgnB822SYsNeO2MX/FlNlgpBHr
RnRJznTyJu49Kv0AIwRwqVGp+N7taxAKDDj+GPQGhfRDlp5ial5wOU6tp9tZ
0gvw6N+0n/u+Y1EWsbAt2z/KeWbdxh5xOK00COCe1qP33+6fRBIbaQU/RUfh
pBzBGveY3EwxuXk/0oWaa+tpXnpidYge9JSFzaLQPFEmPqdLiFj1SzXE4kFs
UUS2OUL6sy9D8hqNQm9Uoeicj2ymEZnqVHMLkerd4fl9Zo7W+JwtnC3iW8Nz
2h9u+b9Rd4hUkBBfEw6lVjtn+4dQT+QTmsdxj2HErXZKJIiiVbV9DnxW9BCD
figvlLs/1UjNJDpqlSj1mHzejNP+fpG8IbZIMyAxUGdZU/3JsSi/uXzc+jkW
Ua+95fkIx/Np7wQd9lgLoCIj3eMo8yry0LgH4GCenegoP8CzQ+129OpiGbL/
FEOlPhegyz1EFJY2tP4VvH1ptE+fjkf5ez33Nsan9Jch50L+AyXrCYwaBFfV
zZcGXWr2ELw0RkPRZuQWEKdZ5v+N4WIprS0g+2ifE4LqQNK3ngtXGEQzMa55
Xp6sFmlTP1nsdiMbpZVR1LZ24+mknZ4HwHExpsLE1LmChuPrT0sg7gHLDkA6
NkVWO3l5zrJjnNLKiRF4wbPQYCIVKT7rxrnu0yw3qCjNLOTPWtgV7IKnJC0U
nyafsJSLpX1gVEGJgkcOFmbwu2qRdABUGvADs9DvQfd13Km+XyqHRQB+iUO5
EjJToV/LmKTXefQLbIEXuNQ1zvf8uPq1z1KjQVBXdsrlxTYorkyYakf93cgq
AEhrWa9zFfKZnnLwgnWj88SsZaewE9ZtgU47ZXX1XmQxhD/NwYVpVRMdzztE
fTX04uF4hXtjfuiab4UVpeBqU3k7xNvrXS+kaTZ09UQjeBGEqWJ7ro4voEWa
TFwqp1QVXbSdWMBcWXTu/y7L0Zh1JrAG5vibVFJ9/r91z+Of3wCgR8P9JXqA
D/JeQVkEYP6pzK6EGrarHtMeRKWIDIKFO7w/wXohJ7soUn8Vdd/sx5/NBXHj
OsvpfRKc5AO5OK8CPCudnFuvvLTu3q0qfosAOhharsbGKRsPit+09U+xM1jm
sjgmb8+CmP485NddSU6hdTK9n+9T2fCcN8o4OgcnvV8xfNYK3H4S9At9BSMh
6/x6G+k0tggk/Z9NvVfKyGZOSs3xe+EwyT2TLin7QqL2n0OkPdOq0ntd2Q+v
y/RiqJ3UVl3IE2pQGSUzqVyGiov40suK0X8qZLZ6/0xr0RLAdjrO64loNep/
gR5LJCeeJdCShBKSG5XJx3rfTwMg1kDr4N2Hg+InIYvg6WH4fD5xhhXjtVlc
VO/aubkzHQPbOZSiW5Ui2ZZGOASnSHE8f+zGMsdlvsh2WO0VBIYSSheJpbCT
pe8hLt92YkoRjBZPcNfOEzzYLatidXnlx04JYPQjCIgQpIxvUEkuefci+lWM
03W0uS/OXmM66HFpl7jO+WZcNhIujulql/WczppjvHM7n12ODuRunqCle9Wj
SxI/FJiTkgrxHWHHxX6VhyZmYcQpROrne6C9E6McxIb4evn8sPlHPT19Oh4+
S9N5LENPucI0KvOdWSeBmg96UWMdeqkNQohMAa/XI4TlQM4/GhFzZSFO1GRS
a7hZy+sBxGA2Jl8YOUEDP9Qbmvbus2ykUVYA/M+jHoTyXYetDXLKnGs771e4
ytN5b8EHl2QazBKcDmLpylDXIIw3qa5Iu3aUAqV4JUOqofre0VCYzmEKSPk1
+x6ul8UVjZN8gOhVm320YRwhJB0MzaQi0Z5JbTRHlhkbPGd2qcM557zhJf83
nWlQJ06jTbY4VxeDqinEyAHjr40DPLAzdzKr8+2pw8tWIus0eLfukT+1iRLm
OKSbuxrHQenVw3sP6FfeSapcsl9NJVi6ERBenTH8ES4GhWxapPXsUdWhSUcl
azqX1rgzmFnSYhRo+riq6pBkhERYCrFGniSODI8ZZU3FhyVd28ZAeBqUs0lN
DyLNbGZCN+K+xWzPHcSHl5721syfifI/gdT14KIe2nCVAkNbnBI9IlovDtcQ
5J0fCGUN6azPFNaZjBAbA4SwAnJSptmbE+WVvjthAqF66lxRnIV0ZNh4YhhD
XCiZk4HQ+lohd1msxbR2LXTA2dmEWvInFMoFH2I0pWwvi0mqhIeHKdzeygR4
egK1owzYn1VRals/G2gskzGx0g4mYgxbb3eAKT+E5czkTFeXrbE2Dw9Fkf3f
FBHnwfu7ME4HicEupXVwxPNWyEnlFuuFi8+qVmA58qa0FU63cdIhVm7TqUCU
OJ/OL/1lcGjn/mC9xYOCOH8KEOBby7vrWm+1oTf4UnI6tYlYQ4Cp+oi0b62T
2EBDwauMrUxIKhbeTfxINKuFunU1Hqm0HHigjYJJoig6ud9DvkqNLNO286TT
wPPbplKY8UIHOQcjomrpITdzVjKibwNaqkEh6IxQDkKE2b1YgSUEOU06JYQL
975tYLY0BGwJyje+3e4MW3FYbPGc8yM2ekRC+Oi8Io0OIS2dPvAklcs4m3N7
YgUCQO3VL88xmkynTSFI1D2iiEadrmtNYJSA4K3xc4OXLLrNXEfav/d/CjSa
YODjQCgH9/k4fKzrQrOgZ0gB+1RUN10ShF6O9ITDlSqBAJ5x3qN9kgSHdrnb
4BJG2Ev4ozVHyVKl3Ptp/qzI1FEFIxrOlb7BtpqLd+pyVLA/URSAQFeGIjjk
+0LUiWnBgqUa1aW3U5h7xQiFR9bwUJGsCwqj/enJGiqqT9IwLttvOBsrSIfG
WYZlcBsp24t18LG4m4UeWHQgxfShW6Qeiv/2BRo7zf7gRQVp4eKEKLmt888i
+bjZTPK95C6CbGYfSHbCCltT78kw1ehOCTBRYT9nT+qFst8PIRDSXOeIZaqU
x9SSxTkoZrKH8uy8SLy0waczU/b0UqhgFHCvuByZ6orIZPdZXDaVQ6dWbK64
zwN72Sg3ATmB/4s9rlGU1kRbvufVAv4KAR8dNJJfGm0ZJZr34ZGN4iRggEOV
uVPJb2xAjvhQ6elhAO2rkHECWlwZSxeIw0vsLUodQyTaNSv8k5ySRV3rfwGd
2+MCwV5OVXDAh+hld0+Brc57crN5cxCjm7TOuDk9ohqxc0e4KrWvQDqkGGCn
KKpxWjSOd8KF+2co1YsQ/bqxLfJt/SnlLtm7fzf7GgiclgP+zMHLvW0vwswm
XINlwSoq7qvMmxyG0Bl0hNalNlUpjscDiNgla27SF2HMj2IIcXDN5TFRRLCD
HAVxDZ/O3NzkCiwWmfcD4M83bAQeE4Vo23p6z/cXXHJOibu09tOZtn1BGhQz
EVVsqjRhJlW+LAJLkI3+TaRVak+Ho2g2FyrNTgTxeWgD/pbTSJNJ604V7n5f
XdRSye++21yle+LMYVYI+OYCru7IR+OB+yrziDaIP4mkdoKK2tLOpvkOtwyw
LXZel0rxcnzIFbJmt17vZbT8ZG1fYpGSwbTjktrBoI0p7KU+1mR/okKVJd4A
qWiREWVMQRAM6WAc1ABEzIiVtMhOwH/uDj8t3XVGnKFBWhvm2HAKZWN1Yshq
wFXvIhcKasrgTw64b9Xx2t/8OHhezor/YBWXn//bTcuhmM8VP0eQnhdTQ3Dr
sDMqzD4WxRWz7115T1YcHHhWa56+efz/IwEiwaJkhX8oYq2UA2L5yV5Tf+im
58s79sciyIilg6A1qw7kkWTWCIEVvmWDRvvBZpXUbATHpKJlr3pLFdZHE6aG
C2vyFg3wXg9yQ8WlkKR6MyZ6srjJXtBlkIK806RFTr6SivEZRxig30JlMeKo
KJvl5AgRKXOWvprDOiaQxFqko2e83antrbYS08yJcU7m8TKNNzw9SND/rwB+
YLEFc7uklaYAeuSkz8sKQ8mkj18NyJaNbZ9NQ8Ms9tb1hiWMiQCD1PRvfh0h
c9n/Z/Pi5NWjlTdQYch4eRklGF7e9UeIdPkekR/vKJ4p3Vi++12vH6fzucDZ
UObaohUaAg/CM0UTIl6C2hPGExHXEj8eJD8FxuXHk7quBW2Kwc0/LOsAchTn
VvOU0Ef8vXL7DqULyx3lSGD+rvaxNlvRPwnxHetMFG5EO2EMAHI7cXfHAGxv
y9L0H/wQOMBstr/d8qZGfg3O4ZFwHlwGkiVqgDD44sxPW1PR8VwPtyu4sbhA
sFRmD7+cq5ahsiLYwFQdJAum+xLIFBqHoeLwDAoJYDuC/JVdCjE0OtSGVdxa
NvSNyLKl9+hg/XuT7PMpS77SBFcrwoRpHvWVdewh3LxhkIIovhINIkYxTswE
lkaauMJHzyQqGDBuOr5z1tyU5r3D3DcFAxHtNVT5BeRwhuaZlNertaB/6wBQ
ZMME77CR3AK7sl7SMq2fmXOdNh9EMdGC+EF6G14FwwklKiNjVwiOzk8lKDmA
qnF1s3cNlK7HVeVLCmfzXcaH5bHgDB9kJgAmgD/TR2p9L5d0zbh7gwsjGP8B
oAsoALEeocyOhD6p8CZ7eQKaCSa9rBZdsWnkAqUM6E9rvEnbBaMd16Eobk+P
i3u2lsin/wARU9zfNkYw8ihj8CScI4oGlZELQyqojln/liIX0yNJtNhZUNBs
7T8sWRAujA8UTYWgADW8xBwvfMbq2Aki+/pjFse0qabMbxXEgQUb9cW/S/WB
qwXgnAUg8bU8OXDNqFe7LwEzy97UNYHTg5Wu8M25Qw4CjVql2Xyojb16Xs6b
IuhKOmYc3SmRkt7+nelZ9RUDwaVi+cGyiKgr7irLjMaElnqw/6JGOu27pG06
q+OEoDea3WJOntwcw1W0OR1h4ocwEEz08rgcI9M8zTzE7PrwWhHlvL52glw9
iSOz/ZZhuCy+tKYqN3pVUo0WhajQb3U6gGIB9ym70mRigJFivxsYXjFS3xsF
1ZfWRTeB6ynKJ3XiULrLlaEJOR8VfZTycVX0MdyMWPA8pfFVZbo+IguUGVkZ
lrn8VvgiNkCW8iAn9PKaMqWJVL3Sd7mj22G7OsTfEcqaPYvaTEPUT1CUJq81
ks/sA+es8EtoFwcX7XGa+xCqXkduXMBuGKV++z988Z5b4FKlz+g0qqkZFNT6
2rbuDvafU0PmVGTSJC1TuXMKYIum5dXf0YmF7zXAHZdWA3yl1T2r7nIWB3Jo
sBPoSEz26X3T83KKvWTJ/XVUII4+KinLn0TYAEWgjh0K4ZoX5Ywj0+OZkVt9
gkv8i/O3Q5Lix5CJKGhMVB66t6p0y60KfybNeWNDa/Q1r/HdD9yXlJOGafwp
M8sQYD5++kUdU+37kbTcIQgnQNNQu1gTFqF7GBF6fzjwlpSeDJAOZtNlzTXa
gvysL9IMHmRl54Ta2ZUaHqo7DL51cGhb0YS63lBUlWRQQWJwmseR6Qo5XFNr
uXswWNHfMC0+XZxVk2zzKlxxQb/WdX9PaOlWfdyI8uxx93fkJU5gecv1G2Px
H8ZHX5cm7c8Uyp+ZMXKo4IuO9N6IYn/ENudrlxQP+6qy1VbwsA186DsOTDe4
2ZBDxAzU5+M/VqyZXgaWA0Nl//QnH+YRIiBSEHSkCdN+mkbTsiwHdGBswiib
Cfn83+OnsrTvCZngVaCDct4Nu5+KoouBS3igckNCp7iLsOfsyv4E1/v+XDvg
z5bTqGzacBpDLtS+7AAw/fS1JaY6W5W8Wjeby4FlhhGdpdDcVTosIm2qFXEX
Dyei8ftb37q6nBt4borZYtRYseqjitlbRcXmIL8A0RRNsdG8LXQG5AvKSSin
m8It28o2alwzAN08hovvcOARspl0TSFgRRsPNq8kTujOoYWU3amLE5KdrZMJ
T0cdgsJ5Sz6uPFwaCkKZyemIkX6yG8AkK3uqaYFZztUYOF8mfqOM0JAMhvGn
yzvQOiecXgTwrMmnZheOROgsGlSZMe6GypNoWGDaqpU7hDGCTQgLObV4cMV6
QKjaXUqKKw24VqWTOOexDmtV1Vzk5GPyYByxi0DBSCr8duyIlJ6DXpUtK6z1
KFHI6t+2/yOwP3wLoOuMnuDf1KFLRU/166I0tKWza0NYfdxtY7Ljr0O0OxN2
YcvW6XtpCSdzJkAba/S2XNXCo/UoQT8uD8f4Nhe53Oev4WM1PibR2bmelfCj
I1aQNaTpnNNEA62StHt+s+2/PP1dqf9KgbJ7Gga7K8joDrPZWRm1tAsd1By5
JqyGigwixlmP0OR2uGX+8ZHd30jeZ17pGWtQarY71UmNTS+Omi5UGXrqzklM
2RbbeofYFXpgAynYoo18DZacS1AltbL+EMZPPYaqsZGQ3sZgZOTkhv3WiQv3
IbKyapNjBEz2zA2cAVwUWIow8eGD5fxMUStvgQuGNZJnRL4Wx75ZwhS2+ejz
jfYK688X6J1AgKojaj7UJdvK9mUEyvMGpEVGDAOVppC9zD/AjAIlPCimiK1/
ofhpwtyqU6Z9oT1XaLBBIeY2j4KHR+uGSmOXAZpC3TLEDdJ0cJ5rL77sXoJ/
Ruc2TGewqPTDBfuTkCbiP1rusGEXSz5XoZEeeIbNLGrqxhJU0Fd8t1sMGWCC
+aeGP/0GJhGfo+LBDgzeocU6rfGX/9usyLR8joS/qy9jcfHET0ttnLgN1b3N
qpc/iO3KawURiV+3l0851BvMQueiJcS2sXmyIXktW/+E2JikRoTP11hZbU8l
aVnTTASjBvpwa1xTR5nDjoiN4vUJldDJNzEPacWFHR4yiQfrEnOiqqsG54w3
3B/tfyTeMSKixqgc1BBorhG63i6IgO4avGQAnzOHgY22yEjDNtJHv6/InjNd
NKxUGNl1JlMhINZfU7C8QFhJRNklvPSHlQVu5Np+083rAqKyPAMgzTwBYIhK
Zpur5Ky/cjYjFUDjVJwi1MHDtG5EeA/zTXTRxX7Cl2G2OQ5Zc6X/rzOJIFsH
J69P61ANcNlXOGXy3vIz5ZnXjV6EVHYFpDFzynEmBZLXNwgAEEXcSjcLJIQU
q+WfPACuo3OsnkywndwharU3Co0trjfGhPE1wqyj2t0bnWMD1VFr55GJdtNN
SpiVzqIAZdweDDWnkGm1gLdWCbMKCJFCDdcwUWlsK01L0Rxxy8ddwGFfT+WM
hYFY7V7PoeO1tQpLOuDtvnsTKt0cYqRqj2hL1ghWNtEYhBQioF/EeJPPTA05
VxAdPxN54t0i3aatlRCgoG/0Vs5re+VdYmnneFy40Mm8Bll8e2oCgW34fwos
ggqIgVnoD2sqn1J2BJYNgt9leku9Ssr2zh4e6r7kpD+jCnDMBAVR5bp/CKKC
M1V+S6nmRE++CEoHyaTYTfI8SkLEWhkcgNKq6wGC2lsu18Z0Ss4bEXlh0kKT
2/v5TPqT10Q0nPg1mB0exQYgh+KHFDswRxD4tMdVr6ehqaYfJWLXSOLvod5+
x7QIllYmtXGpooR37D5TZkVnkpFNv/pWJHVCvDQ/JLGeNGvKhngZE6n+YITC
Q2yF5ld09K0tmjyJso3DAc5xFidkkZ7XgMGr9YM1iop2wGMGy30m7TArCUAv
lLAkBm1nPaYocG2Fx+YES6Pd5c2k8LRtxHbDzaCeDFajEKFbDpD7Hr60+465
NI26+9arLBF7U/6sYFSrGvQEtPQoY0gXAfOCjkd0F512IFAadbCYiAf8Qj7S
Ip0MoRKaK6piRI7lP2rgYe6RR1xdgqQH7ee9e8BxyVmnTBRb7GUo+SlGuHQi
ptCmvREsjjOubRUmo4UbsefJPYZdJTLCZkhbTuwfYHxqJNo7it6b0iAw4RtC
Sb4CkToZ6mXw5YmaOSE5El+avzTkT8zK+HFYkjdcjdR4wzHd3DYiGnB74VcZ
JRDLivz4/UUlXZEh9tNV3LaCxfITe3LQ2tFt4ntgmHtxuey/dSrrnGFTVsUh
clu1rPsC7uIal7SEsLcDZtUIcgt9iPVby8YhITHCS/lmsELIWG7KUIokqOUT
DpVjtJONScDgc1FDNIZkqcawZPpaVO4F4B9DjrR1kQqfXB5VsbxeJLYR5dGr
+sZJKCb/GWN8pwhpIxbjmDGRpkpMKIytbCWdxXyFtVZ7wruij4h4biC1lyXp
kkws8ILNQypdegu0VdPZPN3CcUMHZlBlZVS6cT2Y6CiX2Zo4Fk7D5RiDyLVj
g54C2pCcWuKLZwA04n3S0p6M2AsN5ja9aJhMxWMy/MnPjjyuMvWOTy0AMCrE
Tj8932TdA8pGGTzHYMXClzTnNa0ydjinIdLKMKJkBaLmBNFNpU1RtX3Iy115
snO465NrG8xFrHA1nb1INjd+cklz90x3PDhV0Xr+g+G7nFdjmx9ZtO2Odfiu
IVSRskJUbHvqWPeerAwyO9R/pdGFNfpKWUDHr8lICFgQdMWvoSyGoDnV+dG1
jeSbvpiQt/tPKAhVlHCPQ92MvP/Y1xtvxIbyUttdMcdj93pHGY6rS1owtZr0
HzNtXplYGLBqfq89myq6fHoZAUTaDKSqT0u7tkh+J9e0s9Qe4IGsWykEw2GB
D1pfrmVNcJjPS3yDh54iDp/kOy9HZfIgSphPrLi5wIfJjfDm76to31q8qkiH
6iCkdLZTfcDnQAN17lhUNTOb1MnEOROuy5izukn1+GugOvhK1XbLBWCheHPx
FEhpJ6mqKuIWFDNjxVm3f+g9sF0fxVnPzHkeeSVr+H0aeDi6dPPZwa0bpMw8
Wil+GenJMAYx6R5LE09mDF6suMedIk7InV9am9dwL3yrNuP6b/lPQZd2E3Js
ZJPqECM1Pn5KSoiI36sI61MM4ncMcr+WXWSz28teUthd8EZNomBEyKc4qn+w
CwcMucByM8TeoTYAHJspPuhpTZ/zrt4sD9t9ZVTo52kh5MhnATSz8YJa0bTl
/23GEaKBjj8f9X1SMagfBb27J7A0uNQrI/qkSiT5L5CFHRDim7HXHpi738pI
7DE+duMOMyZlZsfCRkiQfE2d0FNo8ljzWoESc6oz2oC/gQtO9ihu8F0LBkvY
xnYo84u8L71h7UB4PrCFkJJ6GS4a3GnGHA349OtQhGchcWTVzQoV1JpS6rQ3
zqIAZw3UzQdU0fT/8+4rx0scnOLK0dkiz7xwyNPLloixkGxEY90RC2A4cLPK
hALbwCuVzqQbF/aoNjfEt0Op0RtemMcuba5tNXH3czIctourr9qvaZIZBvXb
mIuBb6uedID6HuPZMEDzxETIWSgCYLIY1G6oARX9fvLAfKbIwfZqI1bqQZZn
/113mOvk54ykhvFns3VyrEnx1RIBA+UXmlKXTgFttXikE4xZO3yK8zxVrP69
FOvRpGBuKmCqsWi22zQvsDJYZHt70MJounfpgBZ6nFgXi3H3tH4D4cTEf3tJ
VYVI5blrIOIXrQmKFkCrIcR+qUrheUy3B3les16RWlCEC1fL6JZqG+Tmep9u
IvaJsX6uUXUubXhOwnKvzO5gOPJuG30vX7jpP9GqoCEt3gv8d1Lhe4W4so12
uW35DekCYPhkXwC4y//xDwqlbdcKzAj98NriY5HirHyt2nrsi514fF+Jc9N8
AGc5Od640MdliBgm5qYx/WE2g0llik5KWfXp3jswSf77j3dIVcmGPhP/v3zr
zc9LYsd4/4ml9c0eo8bRkHC7zfRyPvrY0xHUV7S2WGCnh2Eh8uWJXFNNb+y1
WeMnHpuuqmJJJ93RzdAMm7WvXy6SLMtpHPCGocEMQ/O7ROoj6A1bX52EIDhd
QX7tdj/r8jniloPwclgIixNdXq54tsWVxGk+3jGobi6ft+Ggmcvld415L4+Z
7XKXbvc3IBuSVTH7cXXF4mMmK2bqoXrmFmOGV3gyxgMi01zqcShRTt4IGtow
MikcMmchg8byTm/pf9Q1c2I7mUyrqhRW3EJb61OWCRAquEXBMPbbCXjLHvle
ta/FSewtGpr6syZdyKGBZUZz4nnl92I1ZTqQ9b6VuMwPkE3vdxntczTov10X
8y0WCidZ/XOMDYBHYcn07o7C8fzR6gs2raR9GoU1XdO0DmOrnNza6+DJdX7K
v+Jd5u+fuY3eBFKcyJejR6udA/I6m76VUYN3j/EX+VwyJye4Y9rmh4hgSL7g
5Iq5tOyPaEn72ciEC/mjOtULK8y0swZc9gHL5yrP4ZPeiDPe40qLtyVuR2Bz
N+wtot9AX8xoKSkYOMDEAA7yDZ+qHY8np3iYVtTVgJ4ggbEGorP6EJ9ofWZ0
juNT2GwQ0iNjtu35wdeGuVhFj9r0XU7plf42k8awTIieX+gVqwQ/yQT0mYO/
bYIcB/Yxht15k7cJCmoy+7sZqUJAPb/RgkASe5eUFu+dwk+uS1jP0qN+5aza
GdBg8fRyVH5fLrgrFybFAXsXFZCT4rrztAsUVb4lqWSKhtCkDnFDF9RQgqTZ
p9LsJX9nUMvntW5Ro/S87+9kMspSr9cGm0qHaOiJmJTT9YaiK6Pli624Qpeo
JVQfyX1GLP4cUVwOJFl6FkPt8SJLYoTJUrCGZuKBMcf8gTpP95SQaWremDeW
PNVfCF1P4zSNg19xSky+IRGsbOebp7XdX4lUpAoLTay0CfXzvdA9M0IwrcaS
EdgbamWNPtPQakBP8HOZ9Bvl0QIBlIl2FIqmjKVz5To+LiRwOGRLRxfATi7f
4D15DbPJCbAcYq+68S99B566vFYrduZHyeq4aBZiVHoF63UeJe/Mg0NnIPKl
JsngjtiMPJFq713gmjviZpa0gc3Uyai4XmxvqUQWACtKNKPzMjruwFXcAHuF
7K4H0XIpGC2yZ5eNn5uoQpeQ1tDRDg5rW6qB+TqLOCe+k8W1TQAB9oF6IVCR
3B0vwm1A06HuyQ7daNAb0gO5QVUQOECj9YAOIoSmlR1RcPEI7UtWDnpoIBqs
cScu0iOX8T5Z1RsV3IT/mWWx056FQRrcgf/bhHouTcdkUeseI+uvfG0TcQs7
RiTOQFRikxTQRX66dJQNXJ4Z9MGxFcsU5F7UWVm36OTjoGvGfO9q5tIMYI8z
caPkVTj68liaLjnGuvhqIQU4IFjPtxqltMnS9LWcHkeQyIZ+RUFxMcx9gkLf
vjCqXbKednJxAXAsi2MpEbxl6d9Fw7BOiJMcZbirftMqxRHKBBqbe1vRYucX
FFdaKPhM4SDyZ2u90DpPaAKtU7HIWH6szGtgkt2LacxiXp0csjEiUr3WG6sE
EwiOWy9gt+VVvZIJVMnyi3lbtuAN2YTD9Hwvuw8LSI77HhZLAWOo53eqmYSR
Hy6oynf7TM/WUb1b+VncOyPk1jlG5j33K3LD8qOc6nsHMgNbXEIoFZm+fwUI
2MYF91j81IWtQwBhI6KS619I/88D+yZMCRJL2rJuvIGAIwnSvJzDi8yj858y
fDfC7vX+NKPolyBrgnldkDtcfQ+BInkkX0A8KFWU0KI/e8qSurdUfzjrZUjO
eLKPhb5F6sveDZuqDqd0BQkN88v5mtpxKf5R3RLHtzw2+qHTyqOSECzPMuo4
HLrq3ICAbXumwUggRtowUfzp1jcAfP9nniWiyn2QUCKQZbfwc7gmNUN0DArc
gBEk8xgqBn9lUbOGgdi6eF6zMdNoAfj2+XPDbrdSyJhyQQ9zkwZIamwI/3e5
P1NsDoQDoW8/VeUAYdfcUgLLlJsTap47Q7AQLp7NPFC5CnSIBjCoeTLGKgD3
Bri0lYF1Zc09YkoMZEvtlRKbezm1SwiSVfc/aHfEfbg+RC034dptZdT3bN9e
yMrM5LoJ5iN6QRamM60pXVz+t/U5rOW4I1jy5Ec+imTrt7ESSxAvs61y1nLe
zeXk0HAJAwn1SpGv5+zc4AnmCxAHDfSjCj9+BVvsZfcx4lozWARpw9yBl7e9
UtFiFCPgtkrzzpujTCcZWslmthRharZ/ScqZ3viBPWH9Pg6IDRDrFI/U5SNx
HW6XRExMbNtrUULl/7CddxLX0cExDrRr27JMGHzd1BcFvHZHWR23TNL6TOd5
JJeboB7Xztg3HKnuScRz2EAonn0Z23fo23YDwxqjgmAFd1fvJemdBhiUQY9N
NR37W3X5io4+iQuunSjQtlZf9a3swFWL95CJrdw4XEMzfaYaNdigASwgz5gc
skcTndy19FzAUJFfqdR+yRJR9b0GHmNVjG3ouBNlzl5tDif1f21KHJfKUBz7
O6XIYYHFbk6GqL0ymTNB5mw4xxO1qcPWAHPoZQlUw7s/iWcsUdzt9zdV0dCp
Y4Y/ioS2bDQ0tUxtL2iGx3yE0JMV5TKwsJ2boMMXUsTgc12TfPI+ArsI/ZtG
Qp91qmxeAX2f0lDt7EGmx5LQdW7kMKDjkgpOLEv8jekBIMapZF7pAzWsfTN6
4p15ieQeJpfXLo6I3ZSPb0ImwToRDjjgsx/tKSgWuD9duNfH4VMPbL1BAPHG
m/NtRfltpbWIklcg+mY4Xvyscrae7GBszU5orNkC7VZ98QkU4yM/Dx9PqKRl
C1FgyDcZCLmbHcVH1aRRakCoBKAY6R0H/mPkw2zuhZq4iq+rbczzxlrLtsTg
zoUJIRy48zzhd0Ym63XAsqfGNr3fCYkmn0P4gy6RVcaa07xlO3eVw+s11nu+
MuF4WtWbMrSg21qDLfOSpzqDurye5Sp95Td7M92rc99JtKLbnkg0lib6fwlP
Obs2ubdoXpbdDfh0EEKTZWrAOi4Kp8YzqIHw01pqAL536raHw9f3SANLFClw
VjpeS7j0gujEPC552siEnaSuhVRXBUGhEr39Se0qDGI/frdep2S+2wMESrpN
mTrfN1PoElI94qFc58uKCx6oauwJLYrw39bjWU9E3nVABOErxvzHj5b5rCBL
lwgJ0aHuNPsdZV9l+KBxPFJNswWwJERVfkx62gRs5jer6f0znClU2cj8N6gT
qnpvbkwxFZTIs9G2nHmx+1jFZ++nFNeB/VCxDZ5k97LUTclKA8qksJIyMhwY
ECoGq+3NwNZmSH0lRMJGBu8Idamu4AymWOBTaJPQjwrWoGUtunwr/LDOoU/Q
KRqq5MKKH+8wQ1ypqWHpys5BKKfEttmSlYc44/tSUgVXf609PLsc23hX2tjl
JzMKAI4D4aF2+7ca6fC1b43KtXs+4b8YOKZU5cKnj140MbTGBupkwr9br7Tk
ZgbPQURQxkfV2k60cdFaN8CDoAL5QgUj0NyiS3ipBGlcBaJIDrjBNRT2OcdO
wnVV5GQtmKDrUbcrX9rtLawYqQ6vqcx0gQIkmNhvyJcOJfau0dkXh91HPpbx
x45LU0J61SHz3uKUAsLSxcvaCxGm98H14HjqakTVc7iRgfSexDR05istePmh
WyeS1/q7loDHwfg8UbEIhIRhjN0VqpI6po3wGjV099dS1H30N2Dm3sJX4P1J
1pb7xtGygeZ3tpZo7ngx6f4evJlOVnbLbIpxcZbusA6IhvUj2aln1TO1KDZm
5lvrfKf5JpdcrF/bM1iZtJUkLbMpZ220VMoXQaMGLYZR5pn+hqKE7rYUHUpX
+r6aFOqAYl+z8Wjrs46ZnXp2Xy/Gobdm6/MdhCDTlLwtP+6MchPRv7x1M0tj
8KMzv4Zyx1tY83UvVEqBn5iiXzu2plwjIS92ZJbCpbWklZ2mFAg342XDUydn
zlkuTMXfmO79NMyp6OTmZ3/qoSNXGfOfoR9krUaGZck5ICTfjjSm8VSYWOUX
gC3rhAbLb2NZ5uwcjQKD3C/A9wafXZuCzjA/qdmlQec2dNZceXICBhNpg6Dt
QukdHmBfCE+38ESkIGNAhjQkTw7ZfCzMsB2USJLIsdrccIj8L0P/wnNdrQto
RmNcJQq4gHl+LJe9TCfMLgzpgT0MaY1WE+soZ1iIwzx09Wq1aXZ923dUaRpM
npfRpgMXgCq+di/e9Cqsft0TA8ZVSlbPB6lk3f+KxvjOuLP5Vf7ZA+ioaB12
1fRzujNXAT7txiE05YseqfCE7QO2y2jvQOWet2sNOYLTvpTLPNKod0upFBrz
4+Eg32nJHOGrF911l4emPdDhFDJHmR+2IFxc5ElaL51XNUMsU6spRJZnrcyZ
m4SZwh3S8k/w6xue4kAs1aMc1pa36brHW8ocCQ3ZKYCxmvYAjMfqv4IOFx/Z
6PLBhVG+3f8nvxPCvBTqT6Hlf0p5V4GcwY9gzxaruVm6zCBhesnrVl2pzAgX
14tsB4RjNoWgnHyrfKGoors5EPSm5+9TGJWjPCHwnYdCV02bFsvBEGdhADNg
mW8d44VSlWsJUgGN5OZa45aU36Y8f/qdjisn992arBS1Jr5dQ4GsV2eHcPdA
r4X++aaLFQArSODd9Z/Bzw27Eper/U5qWiyZynC9htj45oEY8YTVF3vcQfhu
wdwoNuPCjer9kZLqBxPE+kL/wy9Evs1O2JFY8bAZkQpZUfxIPqAw1ucUZIeJ
oc8a/ucq5P65KSgrQ104ltcvRaqHR6azfxV5hCvPzskcuDJKkGZ2sCgHgIQG
gMx+5nAtFuMzeMxg8BUznzs0vDwGiYaDwnMVghf6A8TjaKqIz2RmMDLQsxZZ
AVhsDs57GDVK8JImUXfG8hgmAe0r/yWfApEMq1ZutHrUIoJnkQChGzy+2EFp
lXCsFmZR1YnOa5+YqaF23XUm9WER1cPCVkMTIFEUgr4aULtaJnNYCUCQmYQi
XiEY8MyDSHaZN54T50pJAmbzjzqLyKtCrUZfM4tZEOG21OkJ5K/h41ilyi/J
bO54TAdYrPzWlOxi0hpQ2HZExDQtgIamNmtqPtHC43mBG6fhpweTnjVBJBGD
2q9IIvMKoiVhgfqjzcnwxP+rOlFiDibCKJRMRNExfJemR3xX/w78thkGGNOU
ceneCdgGqvbphxfzCSPD9/zHw8jcWEsurBVesbiO7U5KQ4PCXT3/UjQZwgCT
bhqHeeM8dGaZWZpt/755u/Nn6BaovWu6TiFjl6RqS7o5lbfzBusM2UfssGe+
GIKVVM9BGpePzXUfJvXvcYqrHulRLer+7sbHhxPrcPFqWm2TnpIFL4MWm8Lf
uU+5yz72Sjj2EV1LQ/K+yHfgnHK1qJ8KWD0fWZdM+qAqTMTxZ0g5XC28kkLf
oFrgzsF81YtQa6QZyp0rQoSWxfY3QcZcB5+Y3Uxt+dYrT0Nolm78tDKHDvuS
jLk9GXMdgCMAEoDbmVKnhyTayfNpr5Y5+IMweagEpb94bk8IKEcI47u72U7e
jTjs6zmCa2MR5yYTJnF8HBwNhJfAKo45JBszk/uHlMRvEcxheYjMfT+xX76u
Qh5L+NO8QQQOzhLTFxk7W6ahloPqzTE2CpaFyNa7pqp2Td4i656LUBp0yEwx
+tq7fCrS9AfCuC53XUmjif5eBuDEEQx0rZnFYanrbhWi6GTRrLSAe00vFlTO
cPPLVGsL1G0+VBGGR5dj4hP//0eVQdJARZDkw1umPuppwbGm+LU/BgrcPIvM
B24boxL0yyVwAIEW//iyGgrG5awN8J3XmxwZPEpNLftYj19/nZjGo39PIaSM
/Nii/1Rck+4NFrfv9B8jpMCWVHu4G+Pm+XQCg7rO3yjqxyMxGyk4u7WQxEiX
tLAzxBT47wBN9uFbs9spQN5D8N+BquwldLHKprVEPc0JywH5bfedvLw8RzMn
00OsvtKsDC1SHzgQZndLfDBUGSBqrdxgYsFVgPgf81x0k9MMwIZIxLB1h9xR
jwhpQ5ESCCrNxxvz0laJyaiMScdaiEogEMZQDtCyICNWcGxVH0nX3/XGwKfk
eYEFn73WtKRhsn1xkgzbJPBMgm7N+XS+vU68CShy08lfkKr+5ergvGuyKLEw
b5050l9QlyxQupQl1H400MNnpLeHXcHNR/hn8ec4siWW+AwQdILjsoG+W44A
cv+9ooosXOke8552CbbstvMMCJwXpslNyJ4MPqkd+dKUT6JWOoOxbDXzLpWD
McpoTCuuGZq2ZYBhx9F/hnhADPWr0UQ5LEYvVw0K+hegFqzdOot0m6sfu6GQ
p8mris6etpiVKf/pyx81f0COcCqqFHoLO3rqT7t3gakbAwoiHk6enHHeZf5Z
jGIaG7HOS3q1jVL8kqKrk6CGWoqpcT/M0pRJOy4B/9pjpInbDV3z+NG7vun6
pOihHl6iRwU2MzKbhHe0DP9uuYiOKJ36C1GI5ebff3lqD3iZW0ykDl/SU5Ej
SCP9S7xBVp+CZBV181jpwtO3fQ81uH0sI/pFkrM5OKBIiesjWSnGEqwZKLGR
7bOiXRSDYGsfUpCU6yFONl5RTxhw28nDGe6sK/kcDTqPSHgHeYreoUS8+IqP
3yhMAKS6kIHtEMm+zUjtzxHRmuQFHjFmbd5ay7xWsYsbZl5zvwWAb84L1N21
1k+dzg8GBEUv5hJKHiaALVjrRSMtAueQa+vGgUZII/h4NOEaWWRr5yD6lXRr
Yjv9LDJvaIhGOnwrLNUpygmE6qVQftSiSO3aeJ/pwlZW+3giukhkUlu7yDVp
KQMsxSM7KZYaPjFMuSYPsiHp7PIVDIMUx7y5EIGlCJ5X8/gedV3x6QD0Z5N3
MCFwEPEguAN5GVQP4Rg8ACDEG8InvohVMUOP/jnr/jz6FnoceqEM3XVMFKlG
sC8UcHVKxI7eFNNweX20QI6a7aFFLzbpeJUZkLRbtw0T8r3nhP/alszkLSIA
uzPVkIEcB0gw8cAXZWwUeRdQX6n8ub33B9q9xh0vlnH4wlZDJZUxsA1i1yrg
ImJiybpJruc8TXWaArTUGNQuXNVtbdGFAb/MoJv1fwKI+Dx4wlNkEsCKL5po
PHDL0ZV5dn8TPWYRMm8QocXMzm5ii496g9XKWZxq5lNS7hcdAggLXE3ZdWCU
FBUB6KuL9+Is0IrKN7rypvwVUnrPK2I7rVkahqVsz9m2LHV1eFvxDFWNW91p
gYkTVe2cAxGNOkp4F3BD0L0NH00Nj+v6oW7BLWkl04dC+abfE9WMrasrkGor
69xgdVj/P5aLsNMVb5Ne2vSI8brmvXLxcerh+NsiY64oEZFp7Xh0qDa0VlVJ
lkc8COWvH6Z/FuQf+v6z9XkbRLS7sZTq/vMubsoZWkLQnACniLI2REj7waix
lSLr4LjJYto7G1ToLkZtZ7H8igDKJUf6F1Gl8x27APf7zIGKAtE0dbR89mP/
r+ltLnMcfDoCQ5xSUcwpjFNgxiA2OrCPpUGI5E3HgEUidYmJAJVtDOMfEO8w
JWJjePoENRpEOBa26TeoNaLuT/9egRClblrw4Chaf1mGELlUXJk9CoLumFVw
IAtBQHiXj/fmUM7u4WMqQdWy27mSv/DsHOvQdtuAYYBf4dYGWyaWLsKDOytd
fKT50Od9k6nCr5ZGABSnl4boeYq1ypzUIzXtqFQHISg1NEtEay/7DDCp6tkH
iFPxSdWJ6ZzETriW/dRzbGIw3wzFkccRKPCxdDQV4NIzpoEYajIku0Wg54Y1
gRixTSIDzEI7xAB6gr5LS/uAS5IHdveT3e6yG2wwyl/wp/NmWMztKNGoBC7z
AX28eJMV6gBusTazpqgQsD/xOim/8OpriRUrhe3mVGRg+kEcF4fx4YBwQwxc
7rl098Wp2fgYRgS7btFmyFIupzJr4KluGrnMXNkJ5mWrhZuopJ5LgJ6v6yvD
i0HtahuNPKlcLW0/yGdsKhR5o1UU53DurZ49pWr45w7eWyM52wl8HAuEdz82
6JtiUTgmQpM6/aigKADwzNWyzJMiGLQRzJlq50VcMTjFDAut4WDgKdtTzoX+
ytxgT3p6ZKQ+BQP7Z8OsgN8T38BHueH3CQH3Yqt+N9bkuypQN/O0IH94/Rm6
8CtrMiOt8JjAKL4pNMhhkn6s63bB6zwza3lvwPe3vmD/4DSJQPZAt6P0TO7h
vu9JyAbhvoe4pyt5WiKESiRT4YG9RYLsJrQwcnsbrMHb2Pyih3gA6CJGNvKT
wDgfdkdQ0ltaftbHDbmQ+pTuP2Aw2Ce2nQAlMu0t8X8LaHl7UURRpUWxm5gu
N8nrb5e4Wtyk6woLmRFOdKjgydAunUEkNg2Irzqs/TEP0T3DDrQ07MUcjbNb
nrhT3O1hVn83G+6jXBwX9eVJCBFKbiPVY3ANM01Fp3hPJ9isS8JYlltUDVBa
HEdUxwY6h6QGkOOCLp5cp2WRTxIAob8z40Ih42s9jA0m/waUbAZY1EBnIc/A
D/3s5Nt2PrjXccnkB5ktuL/EDQlH8iRmDjn7XGLDdX78TOQrsCX9k/jj5Qx/
ZUmv9RGm1J3xIgxLwyb9XMr11ZrlskuyAT0eNCgKRgl0YCPLBQymZkJpTh/6
JN1rfOPuj9Oyv71CPlIK+1Ud+IMFer4o6P2V/gaD86UGP55Py5m7Ca2mMFU1
HfVvVd7OjsflXPZXYHaNNuHuZ6hCM5uHaH44f4xMmiAe4D5K90xJfh615Rr3
zoVIQ2nmJpLfQe86XOCF8HEZwGNYU41GUJzYPVz3x4nVoTbb+Q3nhatmpsU1
ys/qUB5/4JRqFHFzlT2TayNBuV4mx4yVuvVxCvJaLVANKb66iCuhEgQlJ4wV
i0dt6Hm6g0VynQ80cXcvH266nSrigL5FbQWjyDYMGvKCvObacO0FK5msfqMR
MsMo9EiZAMnh5sW7nu1PmoTB6kDWKsYLjxIBkPE1LvECKCDtd6KaFXfY8+Uc
MsZu0sUyQ1iz6byekBAi3sUUZAFbVsgJ4hHj3Q9avIzlxx4s5bULZxat7pGx
hXxGvODkjvneJauE8NMYsAAwCkA0lroCVQ55iwCT8USjdGZek8yRneFRvKMr
boNZAaEMJI67t4gWAKWxNhI34ZTcxRT8eVx2oXTfNc8wUzTCxnetteLVClEg
VtkMkQymLH27KFyyjkoSIxBqt424sp81XMS1kfWrbEuWAvFEHUwgOQUeorxO
t6kgoPH32QDSswFr1ZFtyzSIx5/91jEcNEWWitiwq/XiSlfDrCDGHNY+qb+9
VwmWgx9VlC7chasYyOM/N/RyvLXdbzZb1RRQLxVBfqrhDET4uQRB4VzMgbE6
uQt+LTpb16c7rjOKfnhLiTzhfJEBKdW2aEWXhsWnVoDWvrgluwayQoruWFoU
NrEKC17tZtbzf2f7Kz/2aqQWyGAoPTMZGwO3wFwcg3C3HpkuvoC1zP5ISfGV
7Lxq1nX/ESm1Mhuj5batIdCD64W+vpTbPHWerIHrMkde6x+aaMXdi+NMDP6W
l/ncMzNkvEDecn97ga1ZzLy/1k+VkxtBtgkWK/bJ4leltOqWpvGBz4ugS+sW
x0miUxFaiQUttU8FSpA0g9Y67qr7w5OfDSvgRkk41vapDr7ihrszlmqXWUwx
HjA0McH7MX9GHHhhAj1CITDPKTK2qDupuaJXO1+hQcgjntZaSXGf/jTgvBcY
ekPMbhuuU25x00ixxC6JO7gQbMzUGPs/i0+XgFw4SDb44eodGrqzWXrhQ95s
rwW72GxL57hhurtQ/eUZJU7D6dtOp+9A0OB0Q8fJ6o5Q47kTfPK3ZYNPzi5g
u/gfNPDK8caAqJ4+GXmXf4FABgXMo/w7UxZk3aenJEikClt1Ls88bQvM+ubp
KPjDdT3E2HkBO72CLnKFi8NfC4emQ5fWBkbW5bB8L/xV+ZONQ5KvNuT/K5It
Yn9Te3p34R+9hKbs5Adew1LuLxxBloEvFORetC2mykqTebCf6aN2Ylmqzg+c
y3TvDQlV539tg8oGZsiJhvdEjAFW9u1rivEn7plTaFF9edbFBFoV6wuX2E6z
2Qzn+hLFUERZpBZKEulZbyahwr1Fo/pGzxNE24SYYNw6Ap+MeTnoRFLZTUlN
ns7b3dgUf0axQN6Fe37lhSxtZzd42nUGiSYZ9WTZeHuHlJWc1yBNDb030SXq
WoJWX4sObH7mVXFAJGj4GutMbgD2d5j42AfEfDf7w8gKGmduVGYEXJSdad3X
jQ/Di7LW9RV4Q8kFTZ9XdUP+vFFlH3w5aKir8OATslGMvSQFOASiFaPpthTt
bVix6dh0FHqquTgCWLwPagP0tfcUyJtNDquoS4afrvIUgOdcB4g2AFPqEyhF
6FCHdRXgGBqi/geFmJsHrlauZfT9cOqmtl8RSx2OFUvkuBAy18CJwZ8LZQJR
kb/1Wgzy5Kt4s/dT3koXPwBbtFfMGhNNvCHLfhXt0OW9KOiHI56E+Oj/Xvng
C2S36B8hH2i4v0iaNO3Ecrutfh5YHZgFf6BdAKk+vFJUXAoMapQJWes3H4P5
cqbzekHVfjOO2cOcQIvyz3aV18emJQlPQzdD7MgB0xMjPJuWzma5GsOWhLAP
ZTRmVnB1ArMPpbfMh/N4G/fs5I9+ck/oy9FydCGU3Y3YnlCXw79PosBaCCm2
km1tuXA9RbvqpvGMECC10aAv2TY28P8wRNP3P7Gk70HHdkM84pv3rCNKM888
03U0HTGsxii/ajA5rvjIqf3n1dSbJmfZKquNq3E2sdB0i2jgpa178PlA+I8a
mmuw2jgAeu/hxFID+3Uqm/95aAVSA/imYFi/rzYhSW/Jutk5SVJIEshlMl9h
lPBYy+YOzKHfpqINmmasTUzrRL/2w/zEJEPjPs8PGHZF9wGObwoCs5UgSUc5
Gb6bXK0eoe6NQCL6L1dODxGdbzjpmZlt93SEFkDcylramMiYMZacktPEe/Gp
qrdORhafW6s5uL9clzTKIy6q1EolgR676KTNoueivZgjmQD5Lhg0sZ6Uci5f
nNKrxUSUSBFPt1iDOt6xLQlaB/DhZ9qlIs/I9VIBrzncV1Ezeqx6puOQu1dj
ZTWvB9tdxrE/40QdG1gqTzbCQojxp/NuyJ7hD6QjbGRmX+De/PONBYt878jn
MvtszYmHcGlPLk6D8p1DQm829qaOTvM0m4qDuMDO6CCszAR+xLeNay/r8QoP
S4bzb91jSm1EVvxTGKXSXs5I+TIQPFPp/XKROplO0QPbdnSkzLkKDIfgoUxQ
iQRaE1edRX/R/ZD0RXjwSN9gTbnG9ksOV886iwe0GF4JQKpyq1lV2CatxCAy
TlwNBgzQdC33Tr3ixgwhDiwa7w992IPfi7mPHFtu6THBsddZF0escwk8/Jq6
5UBOr/x+p0LZSZr0T2Vjse/SW42NCol/XKZ8L1QKhWHoGfBQPG/Zx4nME1+z
Ea+q56NER793FQghqD/Z8fu6yePehrZ1kzDzz2reDz5xuHv7U9zdqIIGmtuf
YBEVmrX1d2yjiaZ9wyAZQQQuPk9nF/euJBI9+12eCzIAOufD++kvCsR4nA+T
DUUjdVlW4G5WbaQA4tsRXiIZxYGNygTQJNTm59RFd54G9wpfxu9f2oNjLZve
XxrzWST4H8fAkxWQG91roV3chpnfrQmGnlysCP6tyyX5xBv3IMXapvvjdHtK
Q/NY8tI/dUfO5sDTa+Bu4GzHbvUSWYQCwZhI5h8zEVwPvJ1t4mZW933dTGmc
smyt+uZPVIK83Kg05+fSj1U/7HnW3Eim7m6jgJ75fgj7hFIImizQ+Rj4qSVU
VsiZKbGASqvIlDL6Ys+3aZK79wW+D4Wcgn4MaU+Txwq9uujdoRWqXgzzFM1m
jL3RenmWx0gdU00+s2nkP94FEYkCMXkTQwgRasAE/sNmMDrsUE0TyjZJjQwe
sUyW1z50eSmo1wwQNyK3Jrs6dwAcaYh7Bml5xxMe0ejl+/TsMoR8aUWZ9APg
XBX84MFF44DfTqiJm0RrdhWIJ8WuPokwx5sOdc9sC680icHyKQGBq3n8q3xk
Xf0i9TXRxCqw3f1wZZ3oRVynlM1kOMZiKlW3OYXn8ZpfSiez6weRx1TBFRfM
Da8w4txiEOiQZsdiAqxFUzT4fanAxyYVBAU7jQspiv2r9Gw5e3wNbkmc0J1l
sCJkAuPtIT1sE7haec05EUsjKX6EVA6vF/22Ir8wmCxaCOJ7VNUN7zvxrIBv
QZuNOeCtTd3gJuxOh79J8v6m/YaTa1BiUyTf+SyD9hFZONPXXrBJkFUUcuja
yuPexuYbjKYrt7NAQ2jYNVW3SUkn4ZT27T0aFxT8Y/KUQNx4RQwLmgFSjyfS
dhqiA6JwUN4UO3nW40yD0Lsuhmkx+Bi92sIM/RFihuEFbHSX3PgRdJkjA4o1
YfJw0pepz/Z6ebLkGYjePzRMbtKD583xNoBB3pjRSULrc+x0IkxnWk77Ckwm
QTXrOBnOD8buUKMfnqjDNMfPEsOBcI4DbD4Q+4GRkBbD3+/+WdvejncYsIRq
6GDr6diPKKGdAkb+QWg/Ee3EhdxC9JKOjtouc632LrfSaiM/INN7GT/wiDTT
af+4Cohq+AxaYTH23X57peaKmdsiC3BDDzfNWe+UtoipdvZDNYo0O3oA7rqH
/S2dnt/uGo53hD42eBuOF4EVtJ2H2hTBJWhO2KKELE4a+TCUDy9qi1KKrf5h
5uXQeuVsr+v1mige/K3wEYqwPWZEMtkSEEWitgYRGGC1TIoftaFS5yQIgZTT
m9Qu5AfV7tpGyoZI/DfRYApHu/t/7halUXrqbRIiEN7g/l1QLRXlVMzudkyN
COT8K28CUTCQEVhAqm2I1JCU998kj9FbI7zlDTIstvc6jsAL5x13JJui7iVe
5CQ1H73nsA+cORtDHmUcY1wynXyT1mLJ4EjPmgcWVqDmOemPPtvPRadHfhWA
Ty0X5XlXg62+7JvUhCRVRInoz+HVjnBWphPx0wJNZ035Ws5i5QLC+f3xnLMr
kSvMk+wh/ecXNQtukL7EZRkjmOHjN/dmUJdByhNjBaRMk5P/5s4F72vXm2DR
KnHClVm2ehVTJ4MSE82taxA5WfW4DTjrYo6hspKy6pAM/UsQ4HFROwCDX0W4
0srsGbndbDpsIb/Bk5uyAA20kUQRx5npjgqzcmgntmr9AMmcSy+1DJ9+avlY
HyIRLYCxkdrMzGXPhxSb6ICSLzf5E5EJXavqtufV3t3iPJw/RY2v/bw3SUby
R/PxD/SuZCV1odpN/8XKo/YVGcJlQ0PIZ28/T3m1Vnrxw/MuqfAD4LWPXNu2
/MVlx2u5+8r/+6EKNuJGG7u8aLEjc86tnXNcUphT9z73Ye48+CM96FWSQkE4
YAp3e7w0VdiybiDmQEYwG9c5RNgUgv03MP8XEX7FOygNhtTEvavMs6BXi7pj
Q39ItdA4Ri9bQOGEgakqI3iBHlezRPFHa1gqhYfsuhte6BF//omMhdJ0abHV
l26UW7F0KLNrvKEiGc06v77a08TYKkOUvZ/AAhqtwlxImhOgdbcNhomqoDvG
2KNhHS1UO65ga4ovWugRztoYLwMAGK2JhzaQmY/nNNREyI70UrIH5Ls9dQMC
uapuYAuXmd/rF0P6W7wfoB7RYlyEiiR1beyRkoaflULl2ACFTaWI6sN1NgCn
kJ0FMwTrTFY1WvDiN+KhclcgDHtJLHcDIDeHf9GE9zdtTghHcnADXeWex17X
drqhI1Dnn8exl6UBQlH1iMP78KXkWNebhaj60gwgNnsgO+8LCvxV2sLMn2Si
/qcTbvKBD/YTJ5iM8rZDuDR1agLNSQBAbOctekacynHiDXKalcHqfoVhcuWz
e0XQvzfKuKjiznGUnzsFG1hIw6Oy5QS/FwwEdGPIrYz9dC6Zp9fe35WS0Fvj
eDs9HOZhoOvPTGHXMA2U2x+a2wJZWbKkot+36VWvCL6GC3iL7qtguXK9afsU
JLlncy3IIonyjww322Q03XgBK2nARXI2OHNVd2tdKxzyycGjK/vRR4ed+IIT
djd+9FVjLCbXcA8bzs4sPIRGHVgSL0wehFH6O/7sK2uDZb/fa+xnGJWEhkZK
dV9b4g6ohGrM8wYkJFyqLy+sAtswBY/MOA+yBykV700Sq7hCYTJtpbxloGW5
0nL91q2keQtB7GlZ/1VLIThhVwquGNSw5hQi+SzujA3rGmLSpZL1HDmQ8AYp
JrrOMmDeEXUodg4qQSeyl05kgg0momECZUpcE7X8j+bSEy3iBJEjy5ultutd
KoachWDoWCfQtuy10A3OPIRXsahGE1M/vpQGHY8rxM8RYeJ05s00xo7mOFQ/
4UsXltMqVYKzgabYgB9rbjBbOenLRGreFBppugkC0SLkAueLhPBAWsRMOnNI
EbpC5YNjziJWS3fPE0wbh1GHYYcS1uwHixVmhGhvgRuL0bJJ9tQqwHcxFzoY
+UKmTrilO6LlU/U4/oSOZ081xafFV1E6ZIMjZNRUtGBbOAYsSIganRAsNc2Z
G1+cjzKWnn2bdMKfVixOAar+hj3GazTWlSnNvupHTsZumHEhXYHwY/bWhiOg
aF7y4r9fzgA1TdvP3hmcXbRTWj4RbOhT9DTrkYcs2HaonZx5aUHbnyifBBEB
PEw9ZJ25AmcADTPrxRNd1h90LD0jG6TW5mNL5ASaj5yuLeKHvIRpTNjp6iSR
GKQKK6MTEiYxx5PpTVdtY8G3aMmGvixNNUzULHqHmVB0TV5y99T0vCmN8sn8
2G32esWSNj75sMVEc/9Pttnycyv/gR/dV3W9tNVoR+TMGKDhd9+Af+Y5BPfZ
8+Qt7Y5i+pD/N9Xqp1ueMVmRXSkTCNxiwQ/ZuCiAziTZpizCtAyq1kbvSAzc
QBOmuhxDkcjSSyKj0ahnZHNIO/wQID2U/1Io7F3hPAhgLKWrVhE5UeJ5EgWc
w5yhSxSa+3DgLv4KR9R8algLhUQdd44ZNdVJId8W1K6k35H5CAp5tGQ2QU3L
+rdN6zfCpWAB7IRACxgob35/TPJ4CrN2zNdgyRRSonTeNwZfid0T6jOuQ7sv
JF572w7H8yXfWgHhJk/GUlgOknstPssloIY83iUteWEo55NUlLZKE1ReB/in
OBABjBJYfQC65F7lJbwqU8zpAJLIEQokMVg/4Z3IZlQLMScA6uVKmi+sPiUp
rUGJDYU2Up3r4SeaO+GRvqkn6nXYNcT9DbqBqbW0ndWUEGWLGWcYoetmiCB4
NfPQPqaJoIhR4IEXgJ/JVw5OG5/hzva8/TBnV1KLd58QvaknC3YWB8q0ynKX
dWpXqFtKjy0WJojVbVWc+a9cqrW2km0cu4EYeFcmTsyZ6eYm42Sk5AkCzWls
O5iJNJt1u/mW0W2LvhsqV5j3X3wTxRA2TFTlBDcwOV4iF7AGW8MgUVeOT1AB
qqu5pbfiAQ/LtFga2k+bcngCojLiei+ahBAjRu+gcvtQuH25T+m9sFq49cvx
YsQnCS/cDGcyKbUClEkXX0WotsfD1DFIive+HFlFNPuu7k7QnuM7Bl1qjwwl
c/B8Eps1gMI6HiLx2mlRf9l4vBDKJKOAF7WrPEnq+UWTUq9A/Ccm4FWTt2vK
wuE7M1d4eCojxaZtFy1Ip4aOCbI01MeSZIv6wuphsrG/fBU8lY3gL4x/9emv
6sqBFtUMLzgRVctQJleDYujMVi73k0Q6ziKGusrYzrdloDEZ5b5lNioGPuwT
OYdrKvXiyTDQLr1iO1TNp+A906ThxgM+RgjvC8AepwTwEVzB3DzhkMCFCQpp
YKvvaEqWz30udyg8TqiGcwWCk0PsqFcRmhJw1G3FkeMNtPKtM16SkB/+mTEh
70rQu5hnV8gXhDQYnE/y851PDUTCBUywJLrcDSoj0+HccR4r2IrgRsthN+yf
AUQcNtAZtOrwhJBbK/GAmYkTJfI8PtTcVORSBCkk2G+/7jvjizfYztvEI1pY
ibzc0G0rKmbWHbDIzadmkLvqU+ncsWe2QHOIfIcIoEfbYN4tDctWpPpo2pCT
gDd8Yn0pA7ii3quPsRFVSkQo94v6HqtDIDh48PMOcavgeDUs+SxdNjI1JjRc
eYhMD5xP7CLq5cl3sboZFOK4JGTlbYMy+GQG/wvKy/kRMCfyxpOQ2EuH95Ai
mraLKVGs+Q5iATTqSGjrjdVDpz9DTHVCQeG1nWXDNMmdk5Q6xVBNjpVprgZ3
TLkuQZWge47R+qVPC/37lepzKLB8RBeN6C+vb/M4zgIMuA3YHDgHhZsWPlDW
SizVvFLyXCy4gOgGc6T23JI4HwxecWiCoY49ayQ31zlfjOJV5Dn3gCUfOPnB
iVZx+plWqd9LNYlkpMQuVGI1fXIDgaL5KN5gu/HwyGUh58FCFVmVwXeLzHOm
7YKXStLlLQG72g9OEzIabOkfmkRLy1hFT7za86upzGE1IvSeOP2ftgpauJqT
GMsLpzqXya4YTO58Urb2ewAmbtluGRH8Nr3CKNptbhCrGYB0dwyYAb1H914w
O4szUzppNoiw6trKm1PmO7csNsRhHXERu87onCYN4icuFL3MlfgHWJyp4EV3
lMByCb03YwMkjBTctxPGSprDOjTPJ5slNHEW9mqo4kxtWcNLcqZ/gRuXxRlM
kCcBbNF5RNyK3Z9zMdS+8wj/e3d8uQne9MO+E8nx2HdP1baSjwdIHrwKLkF+
nJ9zXcqEO6Zqh0eEk/WhMaY9d34R8QHHMw4a/M1cne3/F2l9zo1OGIpo7p5S
pEcl5gJZqjicNtrzQgWeiygAbte6q1U0IOOIqgqRxjYqaLyCISxI2CDqmVOY
poixzzLzP5lxMFKZefSzg2hhb8I7oXINARHOUYFxnBY1KKfwjT+QRDf77anM
BxbcOZqYHrM7w2kss2hSBWgLGW3CyJRh3IQMMpG/5oFzettEK7ulWgPmbvfT
JBp0YffSeWalwyqM7IAtTPTOSHUW1EdYV88pC+hcC11CDSE2mTx+YufR7cx2
AzzBCZdIiDcSOX8oPfexo4DekBeLk2xuEhYP2BSZdsGa1QlSB8U35jvxT89T
D4Ok4EuGtM1i8Jo+WvusEsu34k2CTLDKRODjL38RVeaDEGwZkgdH2F64sWrq
5NV1O7xChWU537AavqtpCoiqQR35MPfH3A66j/VOA7SJHAKArtw6IJAZlwKL
5SRHcNhqh9qM7bQIx1HncS5AM6qRF8RLzl07XC5kaSz7S4usz7T3YkgFyUiz
xnTsa8/fRMusrRGt+B/+6CXF4ANO6/hiUSSTKUJOjQmDc2S+HkkkoNrgqH+t
cO+FjOqcyQOj5DLJNhjM6gyFPwbaYxB7qoJ6Marw8cwgrtcOcfJrgF8mMMVh
4XDQIL6j2Gaafin8uW0SJ4Lq+7TsFoPrU7/RFZgJHhXlsBCzuFkRQTK5N+7Y
EXaHsxlZimK71PUB8nlZOWPLCLWaeiT0aSUwytNtHV1T9CVhsWgZRUhjxfkl
M2egIaZ0ckr7uI3YRy6FWemHe5pvr2Xiijt0uuuECUkAHN7U7biYIgFO1AZn
UAMwk657uebxKBl1c1zoNXpiHaeJOHUYmhmHbc5SgTbR1gldrHrM0fOGdfTS
qp002eEm727DZn8a5hrWTaV4SwlP+cj1YgEhe8zj6fhQ/db1v1kKvT5J1emj
2whAIleTEe+8sDprzhOzABlAqEkb03OK7F/B4Wf/atUvuSB1kbZZqIBHhRq7
EpoiXXGqm5BuE8cHESmi88BiJCCS3gbds1A4AobOSxiVawnM+CGviiybJH6G
c/rmC6YdEXn7+8DCpF1gVcsBHnUIcK96+YiWUYtLptp0+D6czvNtK2b0RJ3z
zCRXNDgHPN+5KP8qXt4C73jCnJ3ZifZUaVKtV/Bqoi5Fj4FlikrtjUHXexSE
hAOrYZ8FDF/ZC9uNBaNJy5VuMXs8rGlTYO7yYL13Zq6kGS/wevq5LK48KcbN
S+y8OhfNuALL1GpnrPHLcn/hi9ptrwbdUg1WNQgf3zTzBoYo4uRkNyDW9Log
h1u7sQ+dhrjqk0oJIGqxfAKdGcReRtsXLMxgW4l6e+O+MIGCU1E7hdsPosOO
6TYpXqt0KAuPAQm+RWAeBlZEK4mBFfJKt1YUZfRRCHoN1+wZI2+zPbkHDC/T
fRoOYkv0FUdql10EdBkE0BQxPXQ/ycC0vucxZDRbObiVMOJjYluOyRhFbDlR
d9p/ttUItI7tDmvlmKrvUt8YfQqS6TS2gVjyQ+/5QEZNuPN81uCxCa3Rv244
zWc4ffrzs/HkWVvfsUT9B6uLMWC6j3LGs9rOfc3+jjFYLeGsHT2dBjrCZRfq
i/r5mv9hVsaZ/WpIiUSs0p16JPoh/5lJTJuZ4jO6rGboewJAD7WL0CTPLOuh
YtYpzrNk7Apm/lcpld7xNlSlTYHbNAK0t4LWO1/I6tkgRUpvJFGZ6lBBVtZO
Fe6n25eY5kI8xwTEp9dXyyGIdSdDZ6J1pIrDVgnc8irGG1fCb1jaNX/oHef/
56pqr1rVfZLtuVH4Q1LfVtxVuRzKgr1utCbHF0Ybywas+jVccAxg2qOOFIo1
Eq+SlnIXU7qDGnU9WZuM3u/It2YkzIjOtsO5SkcUxN0NVCzOdA0KB2Aap1wv
/yTMVhnvPVlQU10ZdsKi0lU5+aBFVcCWQ1vuUcOPzDl3GJjsnXBNl0cQDMwi
WDMWC7cuYirT23CL9TBsFTw7POoKcZPi6q3fmI+5EH5qtDYtxGiVAXfxBkuO
CaiJk4r167GmBY+PblOtDA/fkdbCuj6iswhqY/7qqvhmjY2RqNRgeekkg/ju
IKDwzXg695OeGVRqCGjxooXCfC5gRp04bZco5Qn0JUdu19OrKw5385VJJTGp
0CDbk4+dvyLiKXOgazQ6UzKxU/xkbcTZ5WAxIIZtLkTOlUgRa6XTC0Rqy0hd
lTzCRBfbRenFuoU1AqK3H+hOQORp2UKCNiVde/QNtES+0gdvbDSOdTezqw/P
khTfi3ezCage9aXTqYy4bE3RTBGpGYWT10EFIaq7XFRGCYN0w90tei6CFTeu
6RQpIiKg/1GrsI04ednyfrZUqXLfbguUCxr3wW4piy2WZcFFPi35T5mq7gYD
WxZSR7jjSeW5ydL9IciFlFIfELbOm8CcMWpnrcB6VNsavCDTUhcWM+LDAGDr
Qg/CwmhbDwvaWbwVRnUh8JnMds9E+z5eT1196emJ99wtbgluZY/YzL7XkmLC
p0iUWIYGF4DJpDy3rftPbywjoQLBOTu/gdtLgwmJEtcqsN/LF6OO9EWuDUid
AQK90+Sy0d4GwLrJDX7A6vXtJFLirGH1EID7JYGVJGMD3FIPO1Kpk707G9bn
DuvPhunc74bu7aOGMVMTTr48w3KjWK6H/6TX/Z+g0h3/yp42+fXctrjdImPE
MkMm9+zuRHPjjHHX8uN2YM8UdLNhbO2Uh9xq3jt4+oSXkpw25SCLLRmOk6jZ
Fb2JYifbBXduJSm5MbUx6pqnLiG8L6vRsj5qR94sE4nVR0F2WRafj7bijnHM
ePunfGLJyHMmvAiZFB1khmwHP5a1AlJQt/8JgABEsxmBHBecgE5Ui90EHt/V
8v08OwbX5R1cv3svL/tZpRg8OhWKY2hAaX1yD4rs+zuk/6nQVuj74fgOvIus
uwJSTKfzLaqsn1fXbC3uXthuKcCtaAZ4VqW4Zhi+d2aTO8lAXKOjrBpO+hUG
LP6nSr6gbA6qsbLETdcxN3Ss4xJUZT7e9xYHNCqHY20gJdQuNzZo17eCrKH/
mFPV3pZEDb464hwXdUPK372O5/ICVpWQvcl6AQ9gfP3ZkTdtQShnLSdjRTZA
lWyB0xTokGmK659An60QCOJEknOpElobBuITtlu3ha/4yPZQZLQ9DuyDvaOB
tffTn6YTDqxfMWHhlC5xxAk98YL7eSm40eHOu/OR5OxkuFY7OASeW+Y62Nj5
e/XCH+u7EO34W+zC7bRz8GR67FNDiYZ14LFZ521y3BOhnvEzxEuy+rw/NPjW
hz0+V2XxfIS82hXXgzMgDFU07cEYSdLv7SRu9M65KbSiNcv7/ohXrEWo48Lf
iw2BgZoU+T2BAzXyxKpsRKiI9x+IaHTtkiOFUd7nQMU+iTophPO/3Cbaq2Uw
yxMvrZTW7sxljQ9Q6YE1FfPJJHoq56YZYmPxkGIMZArjO6+hAfMjtYoJXBZE
EYy4wZh3Ep8pddpTF4mMO2reX0mz0Y6t7aXbGvSOX+W7fGV7s8wF7sOF8x/U
j8pOmzXU6OtdUakYacqqLPKHvAz5ozCsNdOFC1+c6F6XabZOnIH0hyt18s84
qQTw3xa+3VMMySm6HB5sThkVDnLJq+ov7jbsmpCv5DECFZt0GgEW7riam6yK
JsC6mCUz1NAy0cQ9+LwQGBVZOBSfxrAJhDGSxOYlQIG1t01aHID2n2rXpeVr
fOc+/hNr5kR0O6kJ8JRjWroy3lp5n0X/FBZFWjdznQGuruJiFl8XKOzqOP2a
qhEEWZnCu+73I+zP6Sto6gJm4NQlfscYEqDjB+cltnneqgsaQTPYusC6rFur
+0tQOEwUF3N3VHJCLNQyIJ2s/cuU5TMBHhnVnsQi3SbXoZN24jyBigMRoMeb
9egYRmT+EhpkhAoJAbRZiYNTM/j2aL6QWbXQeEXZ+BUG2DS6GhMXmjq2TVUh
tIlHojYyCUtC4lnFwTOWxJF9BpRldg1WZ7UUrn0S+6IgUgJNpfgRKKkB6A5S
aJPx0eW2rKauJX4EbICT9CMNd+ccZYHKFj3lmWs92l2sCiycL0xIVetYFvkF
nT5Yku6nQn402AGALSfnNiMw4Ca0yFI5fflLbVYpR+G9Ud49Jyj1HA3Ljawz
AQVqLd58/BOM2ziFat/Iv8IoKTWg400M6rzxZUrl9dBkXZa4mXCIwal3FmjK
n9ohcLNDzhj7yXCNV/3VGOSjs8RQXrmkdgzCI5g+4lzIqoncmII9m0JzSucm
Uwutyer3prsOjXVBEQ3VvLvSoF+TNGInIlZw6aDQrzrStTd0cqbrZb3JxUgc
HdYbuaPj9aIusYS/yN3JXFwMU7gKz2M4qow85gIda4/6HD4dFOI37J1hj5OU
0wBHqQ0dHNxQdwihwtYl7q/wM81xFv/Ovp0tYa/2KcZ7jPRiifU09s5Jecf9
CN6HWt4HjmoaNhQmD29W90eR+T5YgCkd3+QoJFZk5m5jf1W7yue0krUTGWnP
c7JZsQ/FCO8H5PhGD7oJUMc9DtYBMNmgEtjr5uHfRw7pzIOeZ7gtEEv5FEV8
46i51x8LBuDm593M3/N6vy0nuq68Z+BbWBMjCwMjlpxkjsQ1W5bpRS0fk3le
V8+qXkG9cP57xSxmyYxZX8s9Wq4ch4JIEUsqO+NMttJPkxZGZL9qlIBIGL5f
3rSs32sWaM/I1JDfuhsAr8EH25ZWVkra7tMkoCUC1X5lmPmNuU8nynfgXDsu
iFM/WzCku+SzMIFmDsb7XRweGNpFp3X7fbtST1qWVHY3EEIsLjT+PTR1iItd
Hbbokxf7EPT7eUlmmwbdiRE7an/iccW2ebwT8lHCwsWxLvyK+7H8kDmn5RIS
1Ei/Qf2wXzV5dN1aLB+j//RUrs8KZkPSD1+Md1GdRp/ff9/kHDVoOwVjIv8l
z4crsPWmu+B9MDJ3kHtf1wswyXohrFWoKdhY3bL2yXekkc/62iPgbrFPrFD6
0LvLagQNeUankCLsPAOFgi2ORo8oVMJyzt5j3hNLu64VROXtC7QAjnQJ3kXK
x93DRckH9qgqKCtB+SOPdPvW0mG5T5OpZYreC4Dm/dqaAMQz/oJQSlRSODrl
a1+tAv6SpCP1mYekqDu2znJC1Be72u+vYnN0PjSCX0Ho5eAlQsyPIf+5HJNL
MzJT4ClBy4UXsViAkVBEXWAf3Jt851JJfzSlPLK9/+3U4VLQ/4uqbQt0zCXU
xVW/HkQZz4Gy3cVAVpnN4Q/2gxNdKGQnQbkXEnQUWl4Qeg/rCGVZ1TDZEO3H
PK0D4WCQveA7Trn36VSE28uBGlAhgLfyRD4Po043FUqzCe5tf+SBc3fA7KD9
8WXs4IGjY3F2q1BIhXM9A7dSKlBae4HyVHvZpgZvW2c897cT7azhfJ3P11Tz
coV4oUqTJa2PWqe23W4pupXrvH9k0UCDWj5tumBwK4UbIAmvif3dUr9afU3J
k1AcnUBTwX/UJabVGePVTmO2lRzZs8ltiFul3pNpqTTLY8eg0QdR3v5zh3oh
Jqszte4DPFw2DMYutG9V1ArlU3tSwQrAurk3do6G7BDoqBEF29sq9REnN0v4
r17J/q/YExrTJH+ZAF0dPTNPsad+fxeqdJsdYYbTjEn1GUwPKCvMLPlwNlJe
w3ItZGLQ6x+a9info+/vf1wCPNocXL7lJFAoFZRHSF7S3fdK4RckzM/bOXSn
WspJatKYPzkoMWDPJamsU2m0iVmN17MgAxVSWWjHJ3ryM/nVdLfmcgP5VJ6J
9md8Bpl6Y3pHO2b8gXmXoAwyhwdVxH3aO8ECWxpGD+cbryZh8sCW5ROI9ZF2
EP/eTMgPu67kym7CAHgauMFulf6yt7th9B6ZYWOrROteXLeL5Q7Le2Z3v0Rx
CEaAAXKf/EXZFD99QgZkkgcmSo3n859jNkUhpYUMcOxJU/80Q0nkxf23BJUm
BaRFRcMluwHkeVyojw+R/MdkJqh1FPAjtlvtu5b+fPlT7SfOSDBSWNomDj+P
pijxe69pstSqv8RfJjjRjJnI0DkpMDYs+cdQ3e9RxsvnnflCiU0yGu5fHaDI
Kb+d4MCcK1Aij1jRhbyMOY/7rR0pd178B5OZVBdqosm0OycYl+6niLAi0mAB
q0ieDaO5OSQX4eeAlCCtFr7vto1/v6lM9//LsyuzlpO1wQ2Qh/tg0SLAq0jb
sdYMFb1Lm/K/97ROJrKJqNhILzMpfxYqlirKVXpkW1FT0w7FF6xLugU1EPOb
EauATcjBzwdSO7+1YxFKC8s2PY9GWRQZFfOSi+mLI0MnClDQO+QZvCt9zGm3
MxgIH4oz34bt1aIlJnrlqzZdN3Q7dATy+RFtEoSrj1dUlYv58Mbt0v7u5GsV
dxubjoIb1gvdvJF1zMd72fLP0rvg29PslIDnKKU0MZgU8RBduh/l9oGgHgG8
xV/JzjGm9UdxRdBl3lwMufOGubMfI7mItWXVvGJyRnb0Xsl0aNIMmZoUVDu0
w2XRP4e6jN8pbcfMocUJtJubVgupChnauoZyeod1Oh4+nPoqXlBB5nnsjV9a
2qZK2cEYvV2zet7YtXv5RsswZ9VYIcbuxVYUYcW1r37pLd4ZSQpoteU0pV/7
wbpzeoGW0j4uPsWS7iK7GoldqNcpAwsN/S6SX69ThPNQhsOWZIjjv7olCBck
Bz8RHuswVyblXzXXitFBuN7kiq3MONKuxMiQ5bhl9XHB0bcCEz5oKlVt/XH8
hZkU2ZPFAIRFQmEgevtR9eY2qlK+YzKRDm5UcLMvfHfc2/+pKacmtkkG35X2
7TUTqMtS3ObYugCCkyxsx1H52Ev7/u1p2S9tzioP28pvwlARUYw2lHV6QnD7
aHDb9VMK/7xvF8k2emJ2nLSZeaJaCVDMtrFAW9qy4JnasGbQzvC99T3A7rxe
F5TcQ2s8rUf1fHwq+heQ76Fx6rsSf+uiwbd37WV1abXBDVSgKZgz9DuZVzhF
l+A3Dlw9R0Qt0lsaeykZf4SQpdOU/LXe+eRkjr+sDK3mU/3z71X4Ermj3dNc
K07nN7P/Yvvfcyhr0gxL6U80+t3UP7XrmehDOGJDyCWsKpHriVyMaqGHgunb
lV9RcAWqW3eyIfoNWxGJ2Jk8yvi/qhw9yKBYuwXYJe/LM0agPJtmuG/WPjYu
mg3LcCuOc0CS9MYLrr51FQWYGzuvQGMl2opK9ij543MoILMkfdVesF5/N2QZ
KLkn2i3e0WVftrIvxm0ATkJrl7PvxW1QYWT3BoSryYBKFkiK5jvyW6ehN2iM
Hwx5SDbiZbjANlYT1RUlSdy3lmPUyHczpEijax3voaAQyVkPctwiC5V2+qwr
spYZW61x2rbEn1qs0MHcQhvD7MWv2T8rJ4zaUeyQo5uvGttwNXUOqbdiarn1
lcLUGlJZqhJQvp6WK+9wX3oaK+JHP1M32hmlz5aeB1suTZso4sZ4oc6tGTXi
MBe8o3i54Iy52xSlGeP3A10Tol0wBMvfpeI/DB3VdPkF2aoq+4wY7C6qfYQG
/fscoV1AxWZkPbeQeUqtYaDV2fsRTLCvSYSS/KYRbXDz4XSmW/QD/VpSkSB8
os9Nk5gcEmCxYZjv4hIXkdVsgWFi0D7H32EJ9Amjf5kUBek8DKS8Qbt9FDis
j1ZKKVIviMFvCtGOY1imeppA3Qh6LytlybLdbgejcklsb9NGbfCYfQE8sPKM
slh4ZKyJBHxCdbeBxRycfIaSMirftOdBfiZkcq2WBDjS7yUjkO0X2LQPWzQD
ncNeItEHIdSTIB/109KlmRbkcxpENPKt4UK1bQ4NsVHU6QSLDdinIOeVDZSO
XC6igS1NEN0Q4ocSWsIxwi1CMmG02XP3TlB8ah6xCg9tVVEenOCxXtFtuRP2
WdVtyrw4byoIk72zIGwA7ILxerZGeui8q62JJPtxWrNkKNOylsXYpkeySMo/
xlpZXq0chGsEVKPbXSW03zfOOifdTWLJQ7sVtWNnElqo8QWFI8L/BrA2ygMd
OJlk9sPyplnRWIAeBPFhhYFxh8WODRRJhMz/vS+B7i39jRX+jmqJA7X+9Oeo
xmKqbMZA7A0M7qDdzqjnjl4eG8iSY9nhy/2Dw15N85xEujERVBrCw0AlzZr1
C+HUUhlTCJGpJpmRgBXfm6iYL7fqxU5EUPswtApCflZd0qIrDqi3wWDC7krp
4Ab96HaV05xKBpZa/4TUnQ19H8apzD7PtlZEIHEED83ZlN/oxhSqRCLpNNoW
XknWoEx41NcnyeybXyVysqTENE3I7ZEerK20T/tbYxBzqE83CCmYDqMgWuUL
+27df7FYb5obEHwZnqUVMZUEAiw4nHqbgXxWK2i7rpDKhYOqNfvGGpJkT1OS
dhBjMH85WbjDBLqsHOWkBUyD5Q4lXZu9WS3AIQ5GTenunyMjETSMLDVDuqeb
ZmA9R1MxXhe9X1+F8snSU3Cy0WnUc1b69veeoGEs1y/8b09pligotBH31txi
cUviCHbNnWwC2wTo7Am0gUIPzw4s5lfh4RywDm8Y/XomkJeTPWfL9YgHgBz7
QTaMOLCrrfHf5WzgFKFPZZd+1MSjjSflKI4F41UJJgwmZIFrriJDCSuUHb7e
CTrKjMhX1AkqYGOend+CcumkKfSvAaeFhldgmVDx32614fd4nf4d83/g6axh
eByKISy7O85rH8/qLtxtHhKtY3HyNBCYi40lA7CwN5Y2GmE5WYDoPKuu9zNd
bJnOXm4aQHg2IEgM6EUJ0sELAI387gq2lqfeJpG6XjHi3B7EztYu/S3VFS3T
rqaoNp9muAxGCRkwxkYvGyVouofSDWv00dnNibOm1ytyXGf8cfbXwjJj5lfl
PujPQP8rBHXUNkaA7ZV79U4UJVNh4iun/j4sFVez9YMKnM8dTFBTKXWM4QCm
dhR5ghiSSoCCeLA+yEsnZ+i/mAbTFHO69pQYV4qBrQdKXqN7PslwvuIJrPGt
96Yuc1ds2FjpTY3rivpIOkAkubDPL2a56WL79yLLf+BknJBl5VfDhZHNvC2I
fbYLf/kmzFS2jdTt2BFaNh7VbjxiHjYoxFKRheP0rfRpdK2JknqO2RlMgEHV
1GOn/lvTlRhwFXbUOcnFf7DTizLFoooai3mxaMdtVTw4jIUjisVVbSuyHnuH
23oWv9qnk5fOUGJdOG2PRwz/pkmhen+iQsvrWtMA4sdRuI2Btjnzp2Bll2dq
3lH5eeiHO2c0gh7D4xk/cISsVU5Bvv7RxPjJsaASK9C0hlRQnAflhxbhTgnZ
nyOttd7gcLmJ992mIgaaEr0E7F7QxVqufburwU+CbRGni2hEoR/9IjDnjlmc
jIos/z4aaMXkjxrrnHJ8oyfcoE5c52KLbQIX1Dgua6PtHivn/iwxgweMaroo
bHP4SJEr733Wmhg65sUbh2oEK/cytK8XDTPkBwNXZjZXXMR3fl0Czwt+HM+Q
vtUxRbV2ZHc+7kOcJ8FihOYZhUJUrO/epRhh7dtDSQhgU3g2Sy7ou1wT69Wt
Iw848yrXmca8o8y9DhPYWVLFENHR4Ya1eblaJvrm8xAw5l4ejLcqcjzjgnVa
fdUltTVtuBccgD/eH7laig6akV1NnKdmOXHQdjUKIwtPVomZpy5+GJFDQ5B8
SIcyBBFC8WhVKMb6LPuUi+AgsPo3peZ6BvjXpxrsZIU5jLhdaP8Lvy29Dvul
zwbo9JSpW+H8WJwqp47wgTPZbr8nRSwXZtiYz2pp7fwclxe+RINvB9BceB7S
/IOWFlv8+rVXJ2YBXwquked7lWFE9F3uNcDb+3mTY8FT/2eeDMnTsZo5bOQ7
Py8v6LrmBHUfTmcVvr960/yArMpGelquOXqYSLIL+vnDhUGPlHpatcLN7D9j
mnzJrM4td5JBG9Nj+j1uv4ea+enLoopE9zHJM+4RjTKc3i6kpZNragXaoMV4
sbWrCdVHl3UECYUQvWurZq3AKYjYYCCBQClEoc9AO5PQVYD2hbVzUO3j4mM5
pjyF93pXiGKXofX58qEz8qMslNrpfBmKNRHZfTR9k78a0yEDEM/O4+y3Ve6/
1USDDQNtf6ejkLh1//DzBQJZ6VY43iRKg8cmdiB10YTjkdrvoCsQgGCtt5PF
p9hcs0+oZ+11VFYALlTuxbQ+eKvz3rupmcX+pXEAICuiAq5rQeIQn8aDmY0A
yP22HtjONg6wXDQyxgeqe/8GCmiLgIauoJC43CeBnTB7oh1babf1HDvuYnfg
FALZ60eXkiwWf/QzDSC/GW4oUaZO9ZJqmqRwY90adjSZJRbOV3FWmqYKGugn
NLn21YVkJ7MGYWB6fKTB5KzKxhRWSgwAa4Z/P0jKpJZy5thAtWRgeOTZbDLK
C0Vi/9u80y4JVx7pn976wc3kGXG+8Pv3JgSHnX5zr+/Xn7YLJYC69KiqoEbV
sC30LXiskSdCthVWim2xjk7ocgYZY3DfpaBc5PvnPJNGlpbdIvdbkp4liOwn
IuknZDVPwdziboVEUdsC2f4f9HlCQ2Fjmblv8IW1IOVaszcJ0bwBPYQ76vfU
NR6dQNGfQpCBowcOzvwFtgOgMZX7y8VCg2pB9wrfpBmVqyO2iVhpH5Z85j9x
T3nIlNmod381+AgrANcIsaofs1fhsKiFAIKSt2/5X6sf8DU+9sQF4FDYO8zk
wdh25MtNAc/pK9JEn6c3k5Vo8p+lt+ChyRSwXtFuGQgDqGF6PLQzPpnhRV/D
xhSOHxxjeXgWZO0TJg+r69RnmkQtwqjpcJHz4IjP5g+vbKTsFZolvSD950nf
P/o+qnhctIaEmSCRkppaZ6DqirY8aliCsw9I314vVvMwa0IrR+S776XnfOV0
0UK4DiQOMvd4NrS2OYq7lt8nXoqLnSHmN02XN5P5l197nAb3Fb77DbFyosSh
IL+l5R755dmv9Rc0gWo8MN4uoIYeHT3vOu7V3VPAkWIea8CmnaUtqQOiD9eV
hp+XfMijkOpHCNoHfc5/I7B1+xr8sFAQi4EixidBmHV9Z7jCQ4sKrjxXGyxZ
H/l1vXXMsrALJjFHnO8diVx6xf+NQx35qoOfQaV1NptpCGmnu3s2tXlE0lgl
p58x7cugXZhHTASGJVrLGMZRvaI58HYYp8hwX5wH1cHPvrU1Vd2BINQABP4y
kZSk/ynMXioDSGicZd+T7CAbs82puECHL9ZLn7u5bVOemVLB/azdznAtXqUz
A0RD3xXIc/sXlOYDgikOV65IYdPRh0gmE4wJPDuweIt91GZ2qnXAs8RP290U
JENoHM9eyW3VOdfp8/GeOFxPWlXU+0CSjk3bOl8aiYztGFbaEq9BpGH+DI9P
gNnjkU6xlrRaPBw/Oq+dG7vDzm0kkPd43jJcptQIm5Tf8EF7MBwODehwRUrq
LduFQXEA+Do9ql8q8rKB/CT4QPpAuuOzXbVE93Wi1hFwGKFSqOmjpa3Pk9ju
Z8rZus99vHYIrLSBnXGH/PRAvNzNnAj2NQCJFLcaTtTTzHqpdRwFOg+ZrkKL
2tL/ymusNckEp07Prfpm3yXyCtSgDGnuIsWU6+SBAVdNo119DsR/zzL4mAeg
uCjQN9hy8Gt7Zt5oWfndGNXAQAGqK7aoutV8DKAayYr8blhCDi7SSqOWlObV
fpR4QGQplKzfPz7pYeBFw7QIFmA/CArl9A7zCno4prJIv8Qc+/VDv29Dg7A3
pPbaWi9hv0GpJRLeJmOLMzuSK97EoN7+lrkLu5tRNwPLeOErStySmVdSFtXr
ZA5C7ALnjyBdVUvBrkVTTm6REW7BMV8eZ7AlRp/p9uF0N9PVvt4lJIFGMHFg
glV+rtFgojE6edyG5WZcsQw50McR0Epum951GUZ31JAMd6SRnfsFA9oAu0NR
G1i6VLQWXY7zdEMG34Vy0KQgilsiNmh5o2bf9dLO4I+AJooPhTmWqaemjMc0
fhM5OiYcjHLHYw/RTs4TOvxMyZEX2zRPcpF790g2xqeHdb2UIMEiIh3/fxby
2kJ43tXNgFfAsaffhA3zOcs7nAPYjtAZH8x5CGvQ8st2jHZDaM0Kg8CdYZOk
qgLewlJ4A5Q4u0V+odV7kOi3JKSqmxE1yb2GxR7vf7JG7CFnu4SXVngFmzt9
4ky0sDAHuwPXspC9k/AlPnWbMLUoGU8QO19BrazPV+aIEDpWm29zX6Hfulen
aomzQtmOybZMSBRKDZEUjdVCD7KtadbeXtpx6BW6E+fotva6B4Ol7hIdPQeT
uP5WpO7g6bq8oGmvSYRlzeYdRJ399fcCFIz0uJLOOiZEAUVuifPPpBkU8/Pe
yC07y1HlaMA1Icldw1AWXzqvi9oD/qUIdzcjGfVwTaWkxMThmORo2GuTbW9H
GFQy+PpYFyJNzvAszoWA2vNsmTVRNTy/wW7CCc3ePsLM8G93883V3EUeAmnh
pvml14a+3bRZOrxdIBtIXFuZqMtWI1SaEaueZeUMkTVZR+wziBNSjg0bh+Bq
2zKPqRk6vYkRYSQwU/kNzsbRgpBFWLnuIaaD6v+MSx+T1DTPxDASCZiolO4b
6Ofl0EYFMHY6vLWmsn9QTVZ62E41gBQW0yWxnf02j4Nfgnqn/OHyJ60AKKbg
niW4/2JA5VNajLp7V7Xx8NyCEdYENzzsS8N3gQr5azmrJVxXo449kGR0BuLZ
oLuHdFysRFeC593FwXrzFt0OdmYVYZWJylXmO8efICxg6/2j/3j4KpZ30LdV
n2KVvM9wdANmf39RHnFyUylxClYDJmmiOK2pdQ9zB3WFHy85KIbFtmaRpXT5
ctB0dGtBRk7165fgIbHCX/V2/QreMG+s24v6ZiRAkxqY8UZYLxJiVWYvZzrr
NwG6Jg4v1pZ+OhV84aTu94u53BUeU5AUGs+MtCeOYllqHWOHvqaKOjqBeaOJ
Qmbg3Xyf+q6mArmUEDIfG4DVluL2BdMqyx6bXYWdY7j33lPPg5ftfDiGK+E5
vXF34NjPLQye+9e2hxMxd6aOFRZ10STb8fRAL8U6vJpdKLyGGCXAWZColNAt
XvLV1bCz435p/EHNDSGJBQr1Gam/xa6av3vznqtykERm2Q1FaDKGaHfUbO4W
HrOkdZZ4LfmD5OIVgkrjweJafDXGBuIvD3PgaHJ/d5tFfEyrbwH5vnbGtyqu
DOUX/Xmb9K6hPydMiLZ81cWnH4DqqPhqUw0zQM5l1TZSFg33NsEG3VWC6SrX
SNOcD+gWfP+05ecdtXDSf4PRJVvRR/crZdI7O70753J8l8Ff2PVwGADofTte
2kVNbGDavko39xyOlY356Cflq+fBCG3FLwgQk3AqzuU+D3KhdSF3wkSp5h9t
vNSZA1LjMAJqTkAOJodoBmwQTXi75jrIVlU3hpyige16uYmnyx8dV2rmrKQC
4ZpQtS/9oUhwfaeQfu2f2beA8Obhs7ma17SYUnkMGSFAzb67ZgHCmQ+Far6b
+gj4MAPdvCvdHNa+m2fGLOA4oo60jIspFJtnF/4pr7v9UkaQsA0Wf88Y4lkR
2N6UoCcBELCKQSSQlE6fUhV82W1/O51eLnbFr8/AYzHuD8rL+Ul8qiwi0SEU
NXECI3PEzzAJzf5hO3xQtdtnf9hd1s7w0VfdTiDfwan10W7c3/F0b/OJBT5M
CgeTgvtdwQlsPfEbT0us1jxU8m8xa4vJHziyaWnobsIyULh+0p6yIH4jtD4w
TQ2TTaK+/LIprGK9YPyBQD7S03RI8Ndm3uf7UqtVaGz1yLAQ2B+XUipp9FlE
tL5ok8hDi8p43W3A5h20bfzYbdG8OMtPc4dj4VD0rkZYoVtqdm2VFEH/wdxC
2TRjp2m+S44OfYZ1Ea+GaR37tgb+PVkC5EpQDds7LjGB7OP5774yus50N4eo
4GRIK7sDp+SJc9F40Q6/WdCQMkM3MSZQDpOxbSMIeHw/2XcQ8W+gOU9qkI6E
JsCjomMqBrZEldFeNLphYfKEiXDunlLVRVAuITMAQnMq2KDa9snrWv+T9m8h
zbvauda+apNAeOekiM6ym0v47Jp9tIXiuzKnpXDe4iG6n0hjI1LTsKJU2YGM
45u8UC3kevrHz2WMRFZulrh1e4IqTyUlmYLZegEddb6F8raw+YankDiNKHIy
6lDbPIN03ItSa6mLnsVrKHRkNzqm6dLtUTcvrBhm5Gipxcxyc5DZdVKU+NqY
hdR26IfzooSBIczLEkdKvXRlqh00HXGqqkrc5Fo3ELybT9eSdJaSMM1pp/1u
12j1BhV2lNNcyur9VuBDymm1kIZpmX8OTGBiTxHX8qV58+3agoDROTKG5H1v
UC4PsPvF2MJwSw8YQ0OgqcSKJT+r9VVte5lXVbP8OHNR3dOShmh+xJB28RGK
cjUu2LBz+zs8HQumoqQtGRclVbhQLrvU4/elsHVT+r2oHvi7FYDxZ8UFS0N6
17951/17c/b2LnmFRkiJsHO8TybX2s7TMTbAv9MmCI0VM+gsG4LaLUnmv2qQ
VJ8Gzbud12IG+kUIDzlA3yp+P2TClWNnp3PKFwyPKCtJeDhbKWYymSDKT+tt
olYs77pHJAAKF4EroLEwYoFhC6s01oyrHLdtikz6aac3yuDFkJBiMdG9oe8t
OVnYyEzTlwmPUXFzSlnX+iGy4X9iduiepI3ru4U5miqyyZte2tUum4I1TfOz
0/p7z/BUX0yNTbm14c2NbDCz0FCs1L3NTV8FXuF5aPAqN4NDfBQpn6IQNZrB
DQOxABP1XGBZcS5ySi0L9AveZFvaZTK51ZmFp8h+mSCSE4AVtJa+Ni7LzFo2
aRT4hwzy3R7rjEVQRoC2j+ZJpD+lEms7LQxUHLO0qFRclSqjgJDMc1rKGT3/
VMaiDqRTnBa6LVod1YbPd+VeTZWq2D5kqKMbclYgoJESmp8xGIir5YuTwBo7
xdKRYksV/IoAhxZ3g89wI9Q+IMXjLyVDKzWb151pVzozmMKuMm5CksTGhqcU
OcQWK4NrVwIcWNTbEU/masNmHglORZny1NHen/r0QMtiHewutjKoqRf39/az
UzPFRqKVAPdJWMvEDpNdBFPfmXmmhMPU0SLulI8oo9ertGvx/R0NpNRlf3oM
BFlwWeOiz+t/tlRjccd/hAteioZtEuyi0GqMXx2ix3Q7HEYIdvQvL0jg3Zt8
HhYHp9N4JBHzPL8Uh6G7hnmrrVDuGneQZafTKyw8MqZP/7Os91O47gcFUWYN
awDlijgMw8QccjiLKIujhU3kfl/Zw8WI2NgYyKdelCPWZHNsLGMiU4Bs231U
sigdGZrZT5fTRZSRwuWx8Li0MZOCggJZUVe1gtpLM4cPWClvkPmSxu6q5Uvy
nZ+ry8DXQQ4EUmY9ABO8uBy7QdTEJCyLhrsxMx0jCIY+6f8hcNIuJtKn+wk0
0Qmx7v5+f08GLIBvtQZnj3UeJ3gj2gpRaY9zYw2FEbgLZNTTb0DZZ2wwWi0I
M01CeAUrA8Oegg/Ft9y2qNL4xTyQOjXl3XKkYR9PqYNSet82/njT8lP9BGlx
JvfHHOOoOQGZ67drsQhoR5TeBLeNr5G22paR3LI6vdYjV0UQwW+Tmm9oWYhn
dYnZyhhg+Gz35v1KkCx8N/BLRE5TeyH/c5hM/IHI2tIQdppvSFKzCuINafPP
ckA+EYZJMe3Zx1uOzgyR1hl84V32RF9y02TxTuJANE+aPURpQ+MiXd5k4ZqN
iE/Xg0ghV+Q4avYqbIF8SZ5Co/mbA+N6pAc3CR47KEouWZkvybCUujNWPqNr
k/0KJ8Ex0DgDWCjUQwtJlCjXvCz7rRejqGPcnB2X3aTRuPdj7EfkseaIHv/4
9UL99FCb23tHiEyHmosdvu8LjZcMNbIpyrOZolC2RCxzM2iDX6tymy1t4rv9
tOKQJAbckuVEWnDijwF/XUESBbpp86cQX41NhvrAJd63twTDBrwR0/iGwH62
T1gBFwB2OgZlBrbpEQV+X2oSVaNdtJNk/MRWtTkOhREEDPPRDpEu3MaYCWaw
JemlZgzf0x9TZE8QFnRGVXypRv8NvWfLH7jK9cWiYZpsDqbfL36BqfQrpYkR
Z85uG79GJSNNRuelcJfC4yL7OCtRS/3Y1PF/DPNwdd0W6RyAq/4zPK0hq1nr
ENIgv002vT5ZiTPnZiANv01UzdwQauArViu+7dKOHB9cZ1EFbbNekaE03COw
LQwYwlmoP/z8OfqDFx7TpMeLFfVJVT3Ow2c6mlwY13smQD/uae5XM/LcCDmx
PCqvTP1vgt/HBVIgBj9nAHIXvt3HAQWV0a0fQOjc5fQy5wxIibz06GHMciud
m5kvobn+e2hvOTbacTlNlfw2qLBTRdjAJbYB53svSwg9o8oBuMMg0kLWhiyd
e42y90MDtmzavasnpsRqcSS3S48/sKDNn/25q3t1qJ6vCU4baAFHaRT0mrRZ
D3KXdCe/j60TlOXIjBtj6CXlBsGDrMo/ADkbLgwxUgLy8nDK5YXsAqpEcPVO
wngDkVDbKgTtH4QQjfhxNmvScTseXb22lzqRWb/jYQz2C8oAlUw3lZGJPMcP
yoYEMkbrZ/UGHXgj52BE8usGnGOwQOFcigUG2ZoNPv73BKIceSWtsrr39OrN
yTBiAEuD7udgov5Xw5LpWpatSmpCS7ZozKnjxCxzmxSDkWKrmYULW91Ol3i/
l/t4gUsUDb5hIIbzDFkgvt8o6IuQ5Fh1AhutT4z/CNRvqkrehiyyWmzuIrIF
TbCkeOoCdYXXwIsKbPnqVVgG8BtadQ/aX6SGfj8tunoJE4rrv7/XAPB4cxv1
OdEx7g36ac4BkzX3AUSRaQwmglH3GsPHqunCvafe4KgDxaGFdXfXejteagqq
Ja4yMnGqx98XG60zw67qQdUpTWzHvDpvX6cX5oBl3UWxQK09zpwFnRglOaYo
jPQPDORcsHegAyc94ojSn5HmXDZ1TbZJfSNZKgNjWbafI1Xyj5TyY+JHz5dV
yIe2KDzgpsCZz1Usx94787fl/YVDRP2IeGrr83N9dZEUqvC+5reOaVGeT2YW
FGvQS97fumjzxJHH5jH+NPjFG6hw5bBF5tJzsN99daoccMUL+fMxAoGhhvdc
7qvkeZTqy1uisrlJhkh3S9bh5ZrcQo+awx/9rtTO04l3xFlHXclUxQwYjIZ7
y3uOi+b0NWlsgvHZhcnoHW7UF5iCoLrM/dCrUBo4FDbGgUf9GAfx8BQomZbg
tva4d8mHeVotOXkowVUetGHeeGB+t1kV90CTEhGiUlpMhA9ZRnqB6ETAZJSz
0sI6iqcbp+zPby3ndoMAnZYoJN1DOirMytgRXjIJy4fHh+s5OEqgVyJpzwYn
ov/7cJcZD7MpBD3oZ6E8esyMXSLNDRoq/Tdg9Mkg6TyeEbeepqaSeNpaXg22
53COMqyZXQAuUCf4kxek2qoXhpkoMtNp4fAgiGkORvDM5motZ35Iep7yhxw+
Nmq8ZGM88YyRYISc/BqYHZNV1XMCp9t2tj53Q1Cbv2eUjL7ZnCH+BYOEFblQ
T1m7yOQcZbwap6nBNNMwBQJzFhV7Vxn1Am4DiacJYQFfg8Xsx9F6Supyk6KF
4T3WXa7rlwBl+TReaLaxf+B+SG+ZIfA88v3//T/4gRbitBDbIeY/FZ04uINJ
+AqimfcKsqhvk3nJ5xiezw9ozU3eiqUGX1GeWFr17I5ezDdyNMw3X16l6D7X
+2ZKRYwnDlHTIZ7kOVx3EtFWd/7XXM/o+Qmuc9/wDhDGrqG6/yob8kdX9+Jk
MJznVbX//73tQcyyW000sp3cQ/lJSK7eq6KAbl6v/16vXp8uujCx9J3dpdZ7
VELim0Fxr5EQOzTagCq7ooV4eR5pMePtWOA6KrgcaaedsXIB01zuhePp/WAl
IvapB9TwlDCGfGdqpl4yLTffZRNIhDeaP6jMn4tdiPgOGfEO6j5p0uQRTSc9
8h89KHVpK3Vpc1B7+puzQ7Juap7XINFUW3wRMNScKRw1NdQ2M4hGGau0vCfk
+E+WIOzaOswzCgn0gAGrsCFEj/rv6iTeelcU+2JYIm/O63EYvxZIGIHKVl1E
o1jODExE8FBOdJmek3NUaVeNhhTNK4Zj3IIvTrEcat5TEVIUn9JRXGgYBMhO
0RRXwrQEjQOx+IfG98UYGPtBMN0iscdvEhyTF1EUInc6gb3F73Mv+0QsHNrt
xYgZ+oJLrFMuAxN77GDpu1cSw2C8eAoA4p5PNIJ50TYeH7NauV0k20u6g1rx
51NzqdqzrLld5XoTZqnWMeXh4OVeeaMhlUN6gc8pu+ew811HNai/YWah5tLN
SWO1PWmIXLyJImfjs3lmZ/L20R9ok55DeH3ACaadY7Kuavwmc5Rvnx7W0wj+
JdkfZ5f+YMn5qtVCtxwyX83KJGZLMQqYtc4pktbspH12bDtutgfnUnGs/vG1
G1xekevKVZMoKiWv67dKdtfN8IZS7dvplQpL/EUunb2praxdPbEOX1KtB3TF
9zY27exKJ/dJ7Mu0SfWkNwdPTZcJIB0TrdiKEHmai7XrUy3lViPBIL0z+TEu
83uz7dxdN/5uKLAaVBitjzU7Kh6T0g5vAhqkU2x2Qk5kidW2e7N9q9Cuj5rT
rXt1KoV8O74HRB0bRth9Ro1c+NE84vPDrnIjFTYdR5lYEoZS4eA8IyZ3ed7r
bXSnFfX5P1t2sIxlbzz16EpjvsUXuUompCIo98K6SIGoAsLg7NQ3QvrhVqSU
6Btfajz87ZqvZo4HZ+6E5XAA5UUbAQagZABUchM+SN2D1M7NDpl9mnJAoxJx
eglKxGDQdajW6dOIr85LZ9aT8laR0LW+QTv0ge1E/UAddMPoilBIlD9xasPS
f55H0Q4D6sDCydFh7qU9duwoSYdAXIZnVIxXi5cwHdQgdVW/sQ2BahH2eThk
CLAGQlopOXIbDLmZno/jpUNAJbad5mf081anPR3nnfAekmqIs2oNR0Bd6hUR
gREUMMzBtdvMQ3lr9rG8R/Z7PfHD5kW1tQk6fduPtMFogXLIiwOUXBGJeG52
a/9wwSgZp4YQZP7bD3w/NmY5KEG5coJSlPLvLg3q9EKEWUbOa98slgfJjszE
1XBte43lILtUVgoPUQVTVYqIx9HP98QPygtXEfQ/8cOBrnDnKSDKR6TUQkvu
a+sMcQm6KJ16zMtAC1IbFwKuIlI8CIWy3xKAHhDwvWcyb+grP0N2NmjF9VeQ
LEkbVVskCvYfU5gGuv6aHTrHP5rrbfv969h5gYwP/Cv+HrmZK0mAOb/WTu8G
7OKcr/Qy5fhXpuIwC6u6+n7FXWH0gyWtHCg5UuarX8BAGtnootDd5GFkRWdm
MicCdhCgsErPE0gzqwSklo2SaqbOg8IxRSNNz9/z5TnGiD+xsgjGvUJLKQp1
fMOv8eTWskQAiv1Z14i8xJ6/cJ4Mfu2Iaesb1cQFO86L27EHNM0vMopFKSnB
9NYmQjmUgKMgsgkyVZq6u0I1S4yP3yWPvuBt6NAEOXBC1Xs0J3V9tSIS0c45
ch3rfZ33NJ7wvZXe2qQ3X6a1XdoA8LxyEJ9acFuLblKD0aHcX1BsFnfsnMxb
8UvGstCIkhe1GPDgbbRirB217ADaDnyYTsnZHNC+HT/8owenfTj4iQJRZPp3
3CCQUkitOeVTH9o8ywPbVmFRTrd6uDLK/yQ2qWAJZrMLultjsQHaFHOKwQA8
yPhbm75hjkF2NgCcL0DRV1vWqjJc4N1IXkwmycqtumji6njNWJP8jo2UwxGa
fKb1wu6ve+7PHAbudrwioq9YfhFL1Vk1G7kKVqPLQqgz74jxILmtoqpTNIdD
N9vLkKbGOrQb857BSTnu7Eb709DeroSTHEZDnQOEF64qdH7adiSASMEOwhts
NosBgOnB2t/LDvI5hwnFxAT3c6r9HBwwRFY0ndxRIgxR278fXaHqFCWSz6dZ
QNi2Ho89S3mL29GUSeDZmGxmy3FIIHZiaFqfsTVsGkETfB6o6UC14kuVHM2j
OOn1lmtXHnerV4WyTwDlFG7kmrZRzte/ZwyPsqOVTyCG+HLOmY4cA37q4tss
u6D7MboN/ly7x8d6ewkt6+nUIIyW5daKXgREHOvgP6aXb58M4xlYxTLJKSdY
+6ocwAJ27uPdJDWWCuUjQ/Vugd5AWmyUCPvuh+VVfC2HPgE886gknNLK11Yq
T/lgChhtx2aCF6dU9bysNIRWcApUj2CqGt/nIIKVMUnHnjPg08486EK5BN0Q
jAXEr2RXsD+NviiQUPWT19cNDHIr9ZScYMB0v283RpAbcsJVcWiM+IrZhSw9
jK5jSkGxxH7CX9O+5rmOw3++T06+hM0qbuqZNBSN1X4zHH/n9Q7R9vjgnyWv
d3WdJlPMp9DUuKnNlG8MY5KzRdRQyki4+0n2+SU1h6JjxMnzl/bflVUx2NBG
PqLotjiWI/qiA4DI+uZp6zH4epuKgq8UdxF+1+6DSRkB2+4atC979nnVvhf5
D2V2sMp1utxz9RgioRivOC81T2N4E879lhwSNPT/rhjJi9iEuaGZ+ocCx/Ly
qLsHMu953ZtEijjzVMaSVk3NEDJnw2tfpy5c7pDqoL3a0r/L04gVQwnehQWE
fu00YMoRl09tXJYqmGdxpSdbuH0GGwAyzHAcDfTTqVfXnHiRAM5Gb1C8Yo4F
QY+bYADeTz+kv9gFrKfCBF0T13eoYUTx/t8KwNRtwgS9JfGabYa52nQEPuTt
cClW72KOfBEX6enuSQQmPzzo/v1scppn1saRfnEooHPCfs4u8Q0Wh/3sOguh
QEr9wTE9+v9yhlCyAQUyKhEVnqkPiX8uXv+dkOVacicRjK2VdQcB4Y8paDbQ
AOWsWe3OHeiZuN/LZ0OxrBqs8WuynDymKvqo0VmGS5AtwAKThqoDwEMCl+eG
hxh1gAgzFaign+SzhtCYMhTvCfTn7kQK6zsQnTfzwmL2FyYhBxuW+A7gSdXf
o9Nu+Oywki3IwKSCWkm4ZHz56PV67IRcx0F9euTMlgt27qSQX5tBNDEEaILG
/hS7SyVW8UZDze+pkxFvlxeaswhOLWV6GeSFVjeeAjvC7QtO4D6qKAfvdIdo
3VjFhx1dHce2ix+5c5VzzlaoszOVUA/Yv37T8jW9P1TkrIM5GOIf95jyTPYK
RBQYwOlYusu7o9y2hSppWpxEhl9+X6QbftRdLfbjy/XgqK+k3ec9cPKwIlw6
bO+KNKA9NdAV5tPVwj0DcdfQi9bPOy+wmNfC0gf0Bfs218ZV6QIm7ManmXrM
WWdzcMAyEm5dtt5YVghTgUXqT9H+M7obkcLyZ7SDtXEFvxQ0ACy+vFIjK/cc
Wgt+H5kNtvNm55lhKPGbI0+H1LRWI5ToxTtaCspv/sx0Jsk6DKS/w/fRUXRb
+08PgS0YfulYBlpS8+lxojG13oYwuT2d7BmYVRG+A+2CJIQgmpjslVA441Rq
qrfOEVJBHm2zf1zgo3IEutmNwTzmInKDnv7uy5ygJpM9Bp8DMd6/TcgHt5A4
rf7B3Te127UAARp0x5jN4snA132NNq1HmXjuaEc0WD5wDSOPyKw2aG251W1O
g+qti9WEas06O+R9BVWcleohaJkk/yHBMvQLgJvVi05NIoyXgHjP3yLZXio2
gk+g+08nztozs0tT9u7gekThRFiJAHVkzl6Y77WhEWWHuc+Op6Hj9naE27cl
rNwrPGFHRRSp+KPAxXt6ieP/KS1zEH589iSzvmD+fWhL41aRROFYLnRsMvDn
ZaBFFjqFTdk+f/Wgpyri3Y4vyAF1sv6Lz5K323p058h3Ef0d1uXbRfjgXe3T
mFCxvDNxoo3cGrkUG1JKg1SZHsMhnf/1VGGW+kzP8CVkHoOTPR4S/WctV597
s4eRXHM8m0UI9RqdQ5K1PLY0YoNr2qzPgmHeoA0cQzmNSKR8jjM79aZ+2nhP
kO7utjztBnVeazuko2j5vx2yONVRdjwI1gf9a8gC/qsNqyI5RLnOerNijj6j
ZJJe86eltMp7NF7c/sQPgbKBA4SxUubzUDL9k8q7c6eLsAC8O+sYx4/PnRgM
DIJmgmgJDbfaOgLPZ1cEYTpNPuBN20LAFbClC6y+UoYihlknMyrOBOqk+U+y
2K2j2LG8WpySEuj9tLcNz6YCdc4FtMO2S1Z+PyeJvG3QSiq6nBn414u9C/iC
fNRifW6nx4cX+anDtV1cnI1xC5qNXEDcOpEI3S+c7YpAv+JHDBAdZNgBC73q
8gjUgah04+QcKXCGw7wnfz4aaN9YCVehkWXxnYeOLKdqlT4IN7JxIapn8otO
dQToIyD64TECN/3eO14Z2GIzZCPTfbV4g6izlqeG3NHAgnW6fwboznFjeVAs
4r/E4uwhwPbmJnwyOVMKTjHFrMJFyuxeDU0QKVqK+miM5twtq2wm9Cg2V1rb
Lz5EA2/EHFy8MCFHYHAFm/DuR9aOYkscHhf8iWelUni1jv/sAobKBKJJ4EyF
lO6Pkv3524KKaRB0AcFNsF7WF2GQFJYGJIGh0oXJqIc10FwySz9/PBqN0q+p
t/EVBmaGnqUVIxNNNzJN3Q8hV7HTWq9rS9t07lJWzry36surdvZ7IWyJFzYa
JcKIds12fAXx1H4dO9dG7BwZ19w0koqzGc9FTNNmW233Fpp3ckjMgnR8IUGh
g5up9ghiiTjLVDTF5ZRgQ4f4XI7mMb/f2JfGzHIlK6xAzm3EdMoO3OlOyDNd
Txdz9JxEWa/aXKJWnfHqM1yRF6PLMiSj9gB6ZuKbmKbdial0pLmP9W7/d3dv
PwXNojxpYWZwPZ/ygyXzyNykeVTjXbTcwG7OKlmIuij5SJeiK/EN1L3UygQQ
yfGnpdGI95vlDLsTRb36eTfWUWGFuSzsd3+lCNKIELoKVS4hofS7tQ9HaFdg
HdJhSCmL0IcMsVlhCXUpV0gt0Qz9RzACzUiwiktuNGCDrJSOKVamdnOURt8I
3SyY88uxP79h+uozSbZODOqduHepy0FHk4zVyPguG1DArfOH6dAOfNO+SK6S
oxtChIE+QhjuxURGym636e3AIcuGZMtzL8d4AyaLwqBUGA7S0seonczq5hMo
vqIixetek4O1YQqFsfM/uJDIiwIgJxJVvc3pkryl3AsAc8K5MM6luOhdjRV2
1KYA6zWLGD+MXGG4HTO3DcmCCr9OjG1yAipL3wNHXMAtRiITL9WeHLPfqzAr
O33xFOTf6aIH3iLEYPkbOBUdOuZ5cLpYG/4jGiIK6muZnVhay6X+qDHQ8LE3
+BB5PfU8cslIMjeSMsOMXCNWOJAu5c1+8d0x9/Qr9CZsJ4D4ILJQlHwkHn5p
ys59BmqSCzQxarhU3lyVpVD/w35mVibN8mZHHM/RcGEBZnYVXcpS9N5wQMCj
xHbYWTPWgWMrgSuPqMw6Zdc+Xd6w68BxJA869S06KNlmF7urDrqyUaPmq8iC
NdgluaghuhWpughCMJNo2Zbsk1D0gxh85xqf3iGgqELSqZ9YWEHICzcPcSkM
teqlKk9BzH0fdDcId5vzmCncpkk8FF1IhBobZ6gaMrBG1kaNUPPnbZr54VcM
+ZssYNBnomyhQXJdwaEMq9tyTaqX9n76VMoQap6tCCq7Tw/whrwaWsc0oT9r
oF8Wb5UoGKHwJViXzXi5/yQhx5UPUkRGGM7mkAh9DXOqwUlXjAu4byP2yWNj
2Z6HsCC04qAVDxZ8e2YJnnpPFehJicP+lSAn2m49RZpViJMF2wML/Bi4yqN0
BJGFz960iiP4DDfK8VB7m1u8mnjCisJifD9cHYDEnibMATm4UlYUHlhy9Vzw
GJ/45jfqcKUzOZyDRUYTr3rSSi7tfk4s+f9+Vp8lRPNQ7gUkRlx7OPzCoLD2
BZQ8QF/rVOT4DdOyDmjg/175daHfGC87AQ3AhDFyl4RRKIxlzNvnAefejs3u
hUHSGF/l5bUBgH0qyA6kswwUqatLlqXg0CySdigJglaER9HQdAKssLk1d0c4
QDfN3koHqpj24N3UMbgkpxLnuxX7ALCDG5PeuQ+efU0Lz1502BmmFuDykexO
ImuH9RP3zwdadvmmtrHHso9qzE3ufIUN0i7RNEIMW1K3sdVaKuQaljRLSuuN
EvYlPhvFliIOLNy5SjpMVZmhxOXcLWfRVB1yAmyyZx5L31knhpxHu5CzrGu0
ewwNx1uFzzhDrCE9cHfFgPVv2Vr2yqTqLvfpH2UEgswHMvwjY3y6VYfbtbdx
KungwRhh+n+ihenCb8kD9ah4YdjX7Pc1vWZS/XbPyF2ggkJvpstQFZ/huHCB
nxqEupMixdOPWxHGp9SmGQ5G3qaJcDq13Oxi6J/KmfXT9EuFeYhB+T0woBDL
oN7l9Z9B3ZAsLOps/nNWtxZnROBZcb9oIg1v2PaT17QKEz0KrpiWbrvh/4DL
CHGIJmSQLfQawQKkr++Y7tqzY+g0BJFmSd436eRGHlj6UMwifexMWi/cggZJ
EEwkvQykC5D4Ns6Klj4JWlh/Be4QIopclblOnSDq6FANuibxJPDcV5gqPKla
MLyLAXjvxXeDttmG4cZZvXzxkmbMMxgTqPZxlKzI/w8Z0wQYOAF2J2hqj9yX
HLtPCdVKNl8qcWVTCWDNvOlZy+GAi16N1pVERLQOLZL+TtLPaKoKL3SeAaCl
TE+bEQ1KEUzwRerWVJX5wr/xEesMs4L+C4dnYzjlplhdieZ+FD25e7NBRpSf
RUo+9GN5CLe356Wl5X2bXwOdZGHvqX2G6+HYJ7KUT9pO8D0ydgtZS+ARZAPg
rBczxgfqEONoVBTsyojpTTlCFaMl0lixfYxTGzCj5kw549pbd7NrNMTXUGU0
X+qwlTHw+thrhFwkiBTtB/7V6RUmxOPkavSVkhLfabIMDWgpdrSBPTEsUgvS
nZ8hZACOTUz6MQ41aEmJ2kr/JpI+lhiTzA1Wk5BJiDeJXggTiaQPL6SCAEv7
1N1mQ0f8w5ZSv44JD7Bg9TnYZREkboih/U+5jFdCCg3ik4zqhbC4JxCTCjif
7Sbd1bfUznXuHKt7eaQMi3lLhTx4BPXynX5h2CcXauTQUHQu5pojlUPNOSui
lZLh2M30mYvPve9zarBUynNnV30b9fXtSGhV+JisaipQbG8Anfz6C4xzhMmd
82bWP7dUBx0ASLjYklpb1x9GtWWx+XVK4jnrtG+OQdUwFio8TQqzGeIHKB93
x76gtUVMWYlSdY3ivC4/HXOlyGb/y6bJg8z49C2WzXn+KG1vAK3HHAFJhziE
yx+NN3+ebQ5lXfOtmMaR4KQQkTrVdUhIEVbdGPmFqODfkHtpaW6iWegMnPMw
Q28KQxi/+s1xoiqCZ79aGJghSvg75tcLbci7Y3LhSCCOIsFzreMShUclvHPr
bRn+spdZAaTaqp33orltckXxkGKRi6G1ja7xIMwgiMAccDqjxrshjRRGG1em
FMkMGgGcUQF07CBy8bZTlT/KXmfeyMaQ+zuYiKkyHztdJJUoW0wSv0ohryXO
KmsEQkaEAqp6Ok+YVkrtUAAF09G1fvqjriCcLFDSfLRhueFhBh3OqLMB0S0e
Xmdv5lLGMSPwrDD19ky2o4oQ73tn5ZllJ+8BXRSsuiPTd9y5KJYHW3EZpfn3
x3chXqwZCxmQ2o8FNrxHyA6MxlumP/zFDv+Q63oaI/B/4yK5yOmwI60jbPOE
S/Cv4zj9lDj47+xfUaAJvRPPQG1K+stt20uA9oA/Qrydk4c4ITcMra1e2if0
2I9ZTrcYNrZOtJgnAycV3N8grsP07IyW1jV+U5TY+AAnm/iPQ4Y0YsI8T+pb
JYlj1SdjAK7u4EduhfldpmolKYx3oubWnFCM+kvDYR11Dog2cJJz4ub2fTlx
WBUJpQMhz40PwUk1zIeTbg5mRl7EKdk8fG4831vcbzPbvPdGMgKkxX0dv6DL
uDVexWoS7lkiBIJZ2nmVgnATe9aDkKiE6wbizMYs3zYpoD0yikgN4Cr71uV2
f/8YCjsvw4slruuSSqwRqxt0jMEERtPiKLtZebQtfWE4sS7tikAggDrG+hYP
H1eXuGx7I+m84WhZetBlFVvq/I0E4lGLofoeZXWzSTCjQUaL5BG4Px9DNHB2
V0geUnlxtNhyBWr0/YaeRqRI2iqOaPfhoowGlxZP62oSNP/GTmkUHS0JlBTb
mvvha+75H4HhMtyZnK+xQjkzJXgfGwgyG+Khy64f4XJi3c8lMriGC2r0MzeM
b17SPw32nHpqz6h0Dx0iqtfTZh64eVj0HYzSelY37m7BzfaxYsaRRj6bp7C4
zJS5vzf3NPPxascK+rF0ZGoPou4H2jQ3Vb7gDd2xB2idsHem7TI5uD81NQkk
qLMaSHexJe+D/T+xdF7cclQX7uS8e1s+ApAmEtfnsjQNLWEgeiLn89JFsOFs
7TD3LueqrT+Zn+MPy2eHQwfADjfPAB/zX1BJIk/IGEQqgxQwKlKpybX9hdZK
BxOEJgCMMkeEtA9LAs6V6QTawS+91T3rl8a1J7cBsuoVIkaD0WrOR3FSGTAM
qyCiIFGfGwcIkgwKj+dW9GdsauESqt7O4JyK0lzMD5o2WwFmm2Azvf6Dcq/K
iOYpgn+CBeTdYJD35wlVzXdwd5U9eESrlywdJe4GpuxGkbMrkqjis76LkX8c
82y1qFiH86EZYkHmzH9DSK0ZLfH1y8J2dFwUsu9Wr8UMPE4k9dz1fMCbvq8w
k0ka3lU39IqLLrLXXNoCj54IUT/kvR/ZCEaqY3/SV7stnoqW7voml/n0alZg
6CfXhp53Pzlq0vStOmu4bI1gNAI95r3JOojrdDSCQqtTIoPphGDR7bA1itD5
rKCZ7oE+hdxtOA+ZLkurFel+XNw37oPYVlPkiwq2YgJjHEu1prnHyRCVIFg9
Xf7IqXbhAKNg9jfSPO0RqR9g5PiNorKdlsVLW0qYv+M2jb7T4w8qbee974pS
M3QMM88m/HuEUOFoQNaFrom9lA93PR/tuq8OdNtN9K+pKLFwDgyWOgLcCXyH
5mBpuECRHKLsdLtvTnSACJdo3Oi9EwkTGBbDRLGdBpOC4DhJ8BmIwwufNXU0
ZHpR1bpDhBh5Jsr2XMIOSePQljS+sPpOGS+fE7xCHXzsvD5GGGYRuiSGstrG
STiFH6RzPfvTHKLui5k3UlVj2HCh9C1TqhEjqe2/t1FSk73XVHHOhfYHkLXw
cFjZQfIaU5v/DYXCsET1ZUGaSC74Mx93toA4TrawrPVCjHnJlGWTMzbVl9N5
i2TUNoIWN1yEOKwGUii9Rsin06pnhjRBQs58+QsRnP3RdVgFISr2F3sadfut
xE6sfXem82eUjWlHWascrTuAXosrLswKNepmWAcRF5/YGDqHVPEf87RlZVma
iqHQpDeeqGmyrkK432OLHRrfqxC3zOwEaYsmcDep8EXtD7LRFENR56yQ+HS5
UEsIbizzzwP7s9B38V24t9iRx21FQBlN71UEY1bgyc1fg4PdDdFHcaPnLlYJ
Jn62AbJGJerMo2NGsAl6rkhD9pIVmzdLHHjGyub7ytM1Cu+k11CXdC9gajMW
brEBOHVc+zi7k/Fwk03F+aYEHEKpVpKMvsOhvDECbjhC5GXrCFNXv0CZZr7H
pP3ehT6MiVoJzbkkWCM1/k/yocmjHu4G4UicTNOtKRT5O6KiiLmb7g7ULH/f
jbCTUB4jNXNEjcGvfz7vmFe5TmRJrsU1Ee1J+88pPqE0NJaeJ/cKyAdqxARs
F9ZD2nSlu+QX2LE32yL9sxzF9OMyyH3u60hX9zYe13io5UBXvuINg0fLd+r9
f59OhkqQ++1666pHCQW0yD2CE9FEMWxfRnR3JVP3Um9dtRXxzDwwOxcMHzpQ
V/z1QXu+VSyhm80rTiPU77UdhOZQ8nJQ5uqjtk/ufTDVJb3AFKYXIHwP0o55
NJgevW6NoxRkOTjGsY2blel/KYDHOgVyLyxsMjOG3inhkfwKk6N/rmMoFIE0
JvPnfgZR9VSlS0QFA6US7rYeUPCsSfO91zP0WNbuVf/5Xgpu6o69oj42T/Mn
DrSJkvXpxYJwuo6vmtgKGtw2Hin7gJ7HKikYZlmbYPucdSjI4uKh/14k0OfY
QLAKnsmQZ0KW7GUhhhKMIl1RckKMqE/2wQF8qJnT4WKCmHDO3TzXMVnneilP
VMuEUK5czqmmbWNMp0n5oFQmXTlvW2JcemDzgIKde1OnXo8XHWlhQnZT6Oe8
Bj0v4SlNnKfQxi4ciiDjpkm9HrISYB3gFzFnvFi7jfEX/3IIolmXsk5fZz9J
oqllzn1RYoaYYqolRjqqcyS/1/KCv0ibk16Tdku3uu2CXAU9tyZujGKVTL1H
NW6MObXH1zE106y4EYCCVzp4kYkrWlzX6RQK3viMCK8+e7/Usv723lhkjq6g
X/w1bdZVQFhCAtad406jVr/9yXwX5ryO3woFT2kVAnSZwstXOhCZZsI5CAwh
gH3q2cXVs3LfkcJCQm9q0sJk4Qxf31rOucjj3Y6H2SNAlhLu/2II9VcaUiEJ
rTeJGffymWl0uP9VlgMuQLRwfAz/N+MU+LHzzAJN9ULCo6zlKOUapCBaJZra
u+dwGCErs+Gg6tWPZtWZ3gHLZPbQHvRkKG97w4N0Y73MdsVqRl3aYykf083a
VLcewKyajrz9Lb8j2SKSViq3rQOVmQ9aVNYDN4PHJQjiy+qpM1B44YEt/6i2
d8iaaDeMP2DrMiT/UafNATcs9Uu8rbFj4Cj2x3Vw6UWm1+qqT+1cb8U7avs3
OWJLWrEmPdb/BRf9iDxuKWQV9oRZF669yVRiX9ngCiCQfNR2Ip5v3+jJ2cnR
GcAQo+e0rIGTIZKoGhhshn4HwuHwdZ+MWM3994ZC10AcImZNpZokGFsL3yjY
Uzn1MwmT6XUHhfXhB//wJ9f1/CIBrJkqDK5ia1JhFX3bGmcj3MT/teKUUSW8
/nQwlNUQpGMBBzabIcfsaTWP9xJ4WSSSqE8YUjHTuG8s16aHsPr4c9z1dhsW
G7zJFxke6O7k8nvlyIaERUY6w+zg5kVNRKfEXsrRy4ko3GJ22f5M4kVI8Ubu
XbOQIQtYMB5WM1ZN5or9S2W/EQHEKFzhV/0FOjUoY6Ot24YURwPt00Phz7f/
VsDvP82xo6gGcUVym6s6Zr29+DzgbyqF05vEBh5JYAnnCifiYnJWtKnVVmfd
P5ExER1Rn/LMXBQdyoviagOH9BEJ4fHhCX6M2D3tYGrlYFMVei3b69zMNtj1
1ilLVt73v4YChW3wcC/BzW5M0E38wFHFTPDFjiRzwafuxS4sdonERqN+FGG6
6Rxr4+bd32R0HCjX6HzyQN2aUty7o7qHPu07nhyDqm5/1EnOl+XQ3mubhhtr
hG50xSV9PtKvuCl7ol4TDfQlgLCFE6XhdQDNYTHKdB3jrpE0az8nsN5dowuW
JUOAWN5mYuWILkd/1L1hMK4943XKvVd5+ll2JjT/gU5zqs9bhZ8mnigLF2/q
e1xTQISBadj4p0rMSPqx7Jq5bp09hWDqjzONiuPeT552mdI3jxsGMuRjObWh
+LvTIrsN3GKIfyQcxY2S7fPBFmhypK1Y2M00YCDYhR+mYNBOBzZ6F8daGJcc
m38Vhb0ReHhAs9SalJfMXyrKs8R063VwcZS42yLS1+PZ1j6U4L+HkSS4yAuT
aIUz3OsDZv5rUo4FUEyZpn0sLN2Hc4/wbf2pxV7RBVdCiVlkgv4aePR+53cz
67vrfdfuqYvjzB6BfeTTkA6z50xESpF/4ctSvxDHPWvqST676v0eqQodnTI2
iQU1XxRTmSVoMP0C7ciekH7Qqn29boBVb5Rbyd8iEvBOpc7uO9oROq16wRyx
7swq7KYr9SZEZIh1U7fVNMGeL6ZH4FjlMbOucoDZglgTXccSh5LdnCJvlvm8
mjdsFNEjfg9m2Kgte3KlwiW7ciQGXfnt73GbN49be62HAXu6OMbotlBDvtNK
HVHelysZsQE7QoNS79B+7WiQ2bpxnHbQP8yUZVcqGhtEMHrHviALx2IOCcmy
1ZEnYvXohzNAQZb4d6qXoz9q8GZSQbCtqV4VRk1SmKi4MEkBHa6sYPkhs3FA
5ygu4zgmejtzoH+ktif8ZLLE8hDPaXmgkDk/CDlWJ395uNX+KuhhnIC/lXTI
fb40QNwJ5c0OsE/XlbrkHPY6mHjOmqt74JuxdqhzUhywxzOHhCUMt7OSSn3t
jVVTHpqhsP6tzCp8gwC6n5RjeFtNiGuMehlu+F4Yycw631yRADTAsWgTUgMS
Qspf51q99PCAvr3sf6oXewlM6bk6f0cl0UL+H7ByTjzCCZft38tNei8iDVnF
o0W4L0R1HfSFv3BTz0YteeTVMZg2BYj07d7Gpx8BKWyBBT1osihHC2BoVddL
Bxce6LqjXQ3xnHfnlRGzoY7U/WQxrRAwWQGJxcD0s2Q3yDQEXrM418Pw6MuS
XDqiH63e/omiHxVX0cNz/acO6XDfpEEyIxFcDvZ4G9XhHApWJC8bGQ+iSEO9
1cLC2Y+UWc/owEb1Wp8MS9XUaLkX2TWayhKoo+HvHsQjYqw1yFqG5NaPYFiA
09jgOHwKn+J79MTK7yYLsz6v5D9aNgQaxA0fQ/lcnNVfVwTHyd+4nqEq0yyc
IZIgXpWlV/HgTEzP0yZECvOFlBp1nbtHDdaMVhTWNMHTI9JEzq4OwZ62rcdQ
JtsZw4TmpoLljsFsFAfJWC52iWURtGuK0OI6RGvrER2Xmde6vd2rDfehPkMS
zzNA4fuWm6+0F/y1x3A2cquqWisHZQGxWmPHbxcfe4ECJ789XzZGrnby9KA7
NABeYnAAd+nvJynSZ+0xXaTSOmH+6vLKCG8wwVNDDRuckLlIIxQ4H6uARc8A
4iiJ61cwebPwTxtPPu44sNt68gdSpY3gt9qqDtkP6MUxgYRXUdVJFOE921A3
CzEN42tifwCt5pq/48OBOZHjWYx0bXL1RfxSGWuASnI6k0pGivBe2oEEVXaS
HGgYMrtdeM7pq4TOKlhnyvgELuctfMFB9Y3PVadvs0YGuK+yTyRgYoKlUByY
8kF1luvHiRaWx4Mk+TtFZ+bZ1gV1Ru5Nr/u4nmVCLtqUGfboWOvh7UV4sxb+
muiYmvnTPPHupXuEYzxUxk91AnqTaO812QrKsbs1wOFhkWSl0u6jTfJ6MyaD
wPx1FB4+M4vmVHWFKFETx/DWjDpJ6X+y2T4abu+M5jJmjAmsHbPLbDsL59Vy
NflHOIliOLMfsdE6CBXhInAN7QWeFfg0SmyHNm9F1PE6/+mpc7Cltm0cWTlV
ef+a20ZsKUrcZ4wLJumPPpeQOKljgEGMASBEDvG6upfSGPyg7B901AoM0XqW
DFxEpiPsBX4osxRcIrLmTlVl5j701L+ov4tOAk21/zIX8OWrWiHWMN7PtlwQ
uzTPEE2QBQRnYun7zaSCArZtbEE6URqjYuGVdG04KaQ7nwv/caB+VZn/UaEz
UJ0k7K5ClNlVBo+yjKXVDU6xu1YU6E4l8g/efJ9u+FpQobkp1pKq0rQ9BOug
Wo0EO84g73ZdziL5nHduG9ghEFsQJoSu4rTRY+7VacJ3P8hbUp4DvYCrrqu5
CWy6zxxEU/w+TX8ugGWWmCrdxo+oOx+9cIHnzScyRuUZ0lSxHCvFzJwhQFCa
qZJvyEBFxtmTytLMggVrpmFmwQfig+lm/qX3w6QS9xR8hkq5XdtHKALhE5tR
R8lIFAkIlbSbYZipPH1g8yfOEYKZoNymWS/M3S5qupPgOMg9ktm2ohpXI57s
mD2yJrFozDV+Q7TN8TxQPx+aLQAVxrFXAgsRhglEIN8eip47qWy0HvENgFS0
+dXAYwHJCU9R3xXj0jInJwjP/3ZRKi08UeJSWGLMTSQYG2nZ3QgFKsgikmzw
5alzVVsRxJxqtqoeayq2CSJQf9o8YJWGxayb208SKHAanLZzfsqRht4fvtmP
ZMDRPSoPuWMs10CxxgILNxCmADP88nwOiebse8pTnqBviLaCROeKWVg56esi
q6dWn+NNyrP1/397q09PBEgpAwXCTOACAHBXtYJ3TLLoQa7DzwvIi/WFaYOM
73nRDZEJPQBDpv2ed4wAY3zxb4aMOemDC5NlyU8eEE278GtVPB2zRAwx/q9i
tPddrtZ55XSIdCvmtBZvmDumCnBdoUfVTdYqIj1krGs3LMnIzyuVpuzQzcA4
k6PHQfzlb2hZ/3UuNK2W64RA/wO83uPmBRUfR9WijoGsIoRHyX6geOo0ChPR
mAjYY2emNSYe65GjAkt71CpF8gMadqDlsFkbg4UnPETuod5B6bb4YRNU+KNV
+SdRlKkE8CSKd1i06moguls/CLOf37jmrtJY0wskKgxnvqVgBKbiNbmW6rNj
ZgbGQ+MVBVdJ6L1XTGSIxBeDuhfcxB4BAiMMomO+xQI76FgyhCWs49T+IuUK
xHD8rGxImOsmv8ddYmCE2eD8l4z2B+q40M0QEg7Hve9+txUXHsAwEG6o1rvc
aI3Uot2M+qbVpbHirfYMZkKvO3sILgZloDAQqe4wtNML49zmSYfQrMZ7jzI6
x60NJWdTc+VtP2+iqvC7r6PQ/HSTUMUtSnlGWvEiabFftVEGn8wxNeWfVuEq
lVA9iLapa/WAljxO+rF/PDbLTsaUbC+rMPEZwtgFLFIRNyIXxrJ9eu0dNye0
ctEsq4b50eah1Fv9u0PcslTc4kR/7q2bPh+AMcau2eXuN3hysmILoZgm7Mys
mKsPGi0lr8dYDXXqsqfL4Kv73CqqIA/iR9JqyE/QcvGG0kN9ozvBQFQUBr9c
diMNMJRqyzQgP/1oek7FnRX/wvqRI9hSbaO/3SRpd4PZjKGh/Qis+Z7rfEcO
Jfhz5Wy5TLRNbbZlamFDlrZ3pZwgjsGOXI6FyKEBs/30Ppfn9p08XdPKUeYc
2RRYTOPYb8d+N3bwtS4Dn7HAVNKe1c5kySMCparu+yEok4QjcpNapHHyzAej
1p3Cgblf6WxCREjx7upe6I5KZ5x+vS/BQFnvCjF5I8j6ZwNs8l/N7KnrsTEv
BaNrPGh87w7EJeTnpCsnmfWjDi0jpwKrxUlWMmSdZCEf5Il1SJ1X5P4OL9tD
7BpClzh4+05vZKo1WyTWG5fHPkpMoNF4NwlbO5J84ibvVmHUPaRsoQY5GAP2
G93c0fni/HzD2NRAcakaveJEse8l5JnuTt5GaG6iK20sKLGKb+admnLYd4kR
ljL/jcNuCM0x+HvH5PiPAT/NHnNdwvpxmkVQA7DGzQVo0HMg5m360wUV83Yh
W7SMYU6t2qt7G1kKbebV91gwo6y+NFOmPsKzUup0q32/o9wP7Gl6P1tI6I7/
9Z5XuKuAYUQk9cQBHRSuH9zJ9LrHd8eWqBfrF5uNlnIY8vnDBoG2OtRUj4Uy
v3tdPRizaaZZSb2mfpZkL3Wev7X+w6Kx/rnZ9nb68L9+cTXl2Qf/3IoIjv8o
1eNODg8tdscFonNRlYauRyRdR0ggCYLLUV+Vn23hw0Z5hLFyLvh/HjTdgr0O
BmDMZC3O/TkHma/7PE7RFljCjdvHjKRTTfZPi5iEfCrVLTWhJNbvCBlGVSz1
xZZELZOmkHjcut6l/ljDNCeLecoWd4gJj/eTyaFW2W3i1hLCyR2zdgU1HyfV
ACcKfuZcO6TXexws5ay0oHl+CRqxI9AdvanjcddCoF9OidR5c9YIrlDWO4Cu
ZMctyTbWv6HGy7s02Wzl6hqjgJlJJhEZVZNhUGjQPQ6iz9QBRbL2xlPF3H+x
dqLg1D+F1zUFt4cvEf3W2DTYFuENy/jE4tyQu5tHrKtz7djj3ssR2eF4pcga
0Z9hs8DSfDAYWDnAuRL/lxwqaHHoZa7GxFS+QXSqcHSF5o2UofMEOtJokQBi
0GWsCt+2YzIOXRMc/zfjhyp3O99FKsSLMJa9lH/Y2TDURSoLiCNACn+8jcDz
cOKOMPS38MZazki8Mq+NdoZQY53DSCcn1efrGKZlE0iXOTQZy03X24RzdjHQ
4v0tJEtSi6inv7O4Ifh2oDYIn59iujnYzw9wZL1TloelPK9qiFPMp5AMEhvr
Hc7p5G0W718ypbvDPTtA4EW/SBNmisyVFdJJANYv28DmiVPYSBPb5vYZnThX
99I1KV9OlVDPYW8qDwBmKUOaWM9eRIJEjreKDgfcnpWWGOen5QKC9COPLdhV
p5e8IQPGj6CKsEyqXVdzEWpadBhVvmdbw/ZEu1gnRTLlwzNJvcT3EvI/Biu4
un4+HMz3GwgPeIS91lEHa2uRqfE1skMsdi3+klgFhBGhtmNDSuZyo8HpZV0o
Tv23fDuaHI15jXRDtn/yHkcyjKcW6HrsW2hHX+kvQexbmJcm2FqfMqYur2Gp
pasts3XMJiji2vfm2QtkIFbmkHLAeBkZetX9YWCMh+iHZw2RUA6zNBvLp/do
BCDWV6JRDAz7lN1Xwck31x1rC9WuSVsB9IaRnrAmNQdq8RSRBLxaLISYr5iT
9i3szuzz1slgof+IVHd0UQKLUWqbPcCbh3Z/Eou3UiRHres1Sx2pg1tqnEiN
V5RvMfI3wER+OLYelCXHyosG3ilrjoQJ3lEDXMg8p033rATdX2NY7EtVVySc
yr5QPXCS0u9CQpBiYtYGF2UGkQu4CmUML9qHm2ogV36i0JncsFSp61tm3xGK
6Ro9e4PkaS1nXqBUKPiqgIYckBJRfHUP8AAHA6QQRnegLvXAAIGdU1sdqyG8
bGnBpVknF4eWKnqD+hoyh16O02xkBmnfbAivqJZR/7qWGM5PMmOw9+/s3Cl1
tif12SWSm6z4T0SgLoZbfeNwoLFHFQ6Cx5n3LV35ljKH/nqzeINDQAUnAClj
dJylI8r8RH0dcgd2W7GAiL53GrAdNlK79oYYXRzcHSN2S+V/S3j4xZkRORgV
vpG3m+M4fg1WVZoDeE/LqSEPxViZw6QsFf3YPswoIZprJSvRdX6kQKHbAzm4
3zkNtHZ7hWWLFST/tUCgpgmuYYxnWlDlc+OSKQCO+fla7557r3B34ey1VYvZ
MckRdSW/KDBiFsX0NxJ/XOzmwUt8XCsxntr19ZoAs/t9vM7T0WnAkfyg4/Iv
Sp7DukRcn6FKEq0gnuV9gqR1IcmO/DGs2uPmr9SmbECs5w/mcfuN9Yg9dNnp
U+cnppaPmqIlS9qzP4X2x3Ptd3xZBhjsAUuTnZVCpBG2Oa6M1hbUS7XMSX2c
iIZuD0Qgk9TbnLSnucIX5t64zu/So1HgGRSxxsB+v1fmjOy/4VIP/oUccb64
aoLAqRsQPWmKe/VcOq2sw8KsUm5T386aBqXfcPtXke9OEOgv8rodKC2uddSG
Ol/d2z4/7vw7QLxsN3sX1QBljVxuQT6yslpMlve6ERoHWNZm+G56OQFmvj61
meu/VJkwViLjOMSEyZGAVYF7B+Z9P1h851RSAK+J8ZOv77OaUIbJxGs7UDi8
986nwZvrd84clVYwgbpD/klaw6DYUiQUYGf+hlkMlCHjxGB9HBvYWh4AtAyc
u6X63oaU9VtZ/YToUQx6PJQFNgHe1KuraSkhO20Y/FSMbOEyJPXEW/mvsUws
kBtm3PXp0mO6q87hYWj5kaidNUMuuHcZaEPjf904iX9DuLaCLfyKAI2XR3DZ
O45aTwlvQg31HXCcpsULAO3qD9uAs9xMA1JevrxYxy4Y+lMA5ClNn80V6I/f
ovZc6UCy8wTRy3adwsCCgpUGekmiFXUPz/DIRlLMZkXiOW0aGrs5nDkwp5yt
mgVaH67TXghUgEUh591yJazOzR5Q3z/+St6oB6U2CYB/ZJkLt3WSo9z4ZBEy
IJ+h2JSNitmx5PgdcfN9CYTybESQtPNiZkeiy+/nFIjVHtb2FzN2EZC8m/MX
MKrcf9IZYiX2xmKSs1bzGZgqqR9L60FsRPVLXdcDodq33Ck2+45acY3iIqq8
oImfmSjUL63WNIKru+Q4h/7QhJPiFJRHkNF1rCjn7x35cyPDlPVz4TZBaIQF
oXO7nLuo89K1OaSNHfLCOwjLtDSDmNzupt8syQ9IK+v0Gy5qeau3R2dPwNg1
kiUzemrSnArqc3S53hGQV1Mdao58y/6CnBUjXNZOA4ftgUq6+UpBwQVEbsVD
88HOZjaLHSEs22ghdiI7HdizvjNQxa3UWe8aGxfN+R8fTKPuoSwLIGEXYOvS
2C0ymNrTXS8SzB5V/hwAwfXPqthblNSwf1c0W6/ju/HtMXE3fH9O60F9RscM
C3Vf7bChAI1kgcYhQkdxZu2m3B+isDeiXdsJcy29BJIlwx/T1fNx9ryoEeab
Jsx24MdNAGizUFm+HVt/E5auVdqeBa4GeAEzEYHdaqYHkbAgn8L8CVurW8Fw
EpMG2DLPVfXHNpRubi+TzIhGjIm2yR79Xs+8Ax3Dlun9OflpgCTkv3BVwMVh
AunyPMYGlzBcWPMoMd5IHki1AwPtWCMT05qHvUnlJZ3edg4jjroGJdua2xwE
7aJGDpBD+jBl+bTfGn4suPVGdbfBf5mMSFAZus732dZ16RVEzzhH4cqTQk0K
KpWylmcjVBiRx97VvQD6+szS38locbIxf+7XyE1PBZFLq7AhwyzsAjZ7sXXc
oGI3GFXPCe+yZFvIpFo9/ugZx7KNWbBLScA5F0ZNK1RW1k0Pi1phGGjvMAat
cDrFQziVMoDNS3Ab0fqammJabE6vwXCBygG8Fb5yOMnQLJPKPH8tbeZjHRd6
U/Jb1sT4y6eaB2tFgA1raPHduQt3uhZI/mxyF1PQpswyyZkAxkVCjRdbg7eJ
airPGd+Gl61+765hwp4wJd73TtGG4viG5H6y/aO0Ha+9Vu5W8CiU0Cs7zqvd
d9dH22b+734C+KJCD73cjNmjlynsGUHOY5OEuslufaI4HdfhTgxun0ZXm3Qh
2K3c6Yt4JNz75QWtI6p7pKXwuHl3aBrDFUJeXrgCbELhF4zjrcgciCMbdJ2g
NYLqlFtOXQjHpBsoPhBlJPgcAm53acjxnUve5hI/x0JP/SyszaSBHsKHRjyh
bj2Dlh9Ba5BFJNhSqydxCmw66dTZ1licU6NBEBC4AszUe7P6NfP9K9Qk5J2e
BB6ocQ2pQ0S2X/DEL7sQhziik2mRu6jx41B7/wMDxElroJY0jfhSucNrm29T
5UHP3udZ25c/NMag3T5DG/WmIG6QoCVK5zljcRS9zlf7uU7FARV31XGt/lWh
iJ5uaEiBMi4lRFvL3kThealYy33mEu3G3ouYOXZCiemAvN2j7qqCfqE30y9I
uVeM/gRqvPXvSqWujlWDF/r5wQwCiCptFLYP4j6WCzimraHuZ6WTHzBoF0fm
EmRU2J/8ONjhd9KhnSpBin1io2b8yOe2htsM8ClDSSRMwxdDG/0dE6k9Wjnd
TiaWUqUYcN+ONp2fHHZS5eOWLny8URY5TB8OcDSerXBraFUF+31EOU+6NAhG
Ln6a8Cij/phlYYZyoKikcBcNJJWWLAG0acqEeVamtr/mOO4GuPtMr0XaHCTR
O+lSqQTPnQSKfrUPvXdbOydkSOSX7JQZbv8AP8UI53VYDmQK9giHwTWb4suB
pbiEt/3ih/BkDPcTs2x6uHwkRwTPdPw5OOOnA6a3DP9tLL+bHzLofenACS8Y
dYN9pfIthColniyyEvT29O//L5SDKldWMHLNmRcOUxmAQJI6ZHGDDtoFquv4
AosgRlyYsFDMAGGGHTYuHlO0K9tTbxYMWsCPihevzm9p8txJAzOIpwt15Hzn
xn02oldq1cBVRjpo85yB4WNYwRs45pAoDHRIH+nZv/7k+cwm7W1Y7Sk7IChF
7MAq7hCGhEYFT5/vetuoU3z+AREPSS8C8qTJzpbM5ZvKwHfQhOiD/jrCiLjQ
kibQZhbOcxHl1+vbRylxhqvlxZPddMGESWYQo9DFAQSRubBH2poYgSEqE/Bi
Nktba2Mfiz4VJEnskTtNwACIHP6I/p5lz60QXDQLjd7hnPsWHL/DT6/Px4m6
UbUha4SqmqcFkI2PXNwj0Twm+TBNl85whZ3ytfCF8buwORk2vF1AkWnItF3W
aVahzH87NnwL0iXU/mRbq7IahQQpTUW5pnrhleynYREQzriKxN7MBdVKX3WV
2Arbqa2nVg75jIMfWYV+U7wOk4ijIxVeaStB83ZBwFuepvOWtFJlHfsy5wrE
ElmBu0SrbJh3LK+xDR41jwm1zLsRq1yRFfra1KQeaNsMH64QpOa6bq8Osy53
jVhQZc1pJr5HhpmZ/I0Z0d5h/fxWXhqYUmZcHUvneoSHhXEJYzRAlAJaogCJ
VI/jI8GDClai1VWGbP/RVnLUooOJyrU4K37E+eqkwHRdAbEXT1x35eUC2miW
EXhOJJZxOKr+ubmDX+xdYfb9ztyBKYSyFBfVXO6/DmLfCoGEaa6xq1W8A19J
OWmsfOQdhPbHGPWAysFA5yJfSmX2hpt6VmbaPgzviHcsYtiDg+4A3mnqX+mH
JMJ97Je1xVOwFA/fP6z90Bc4BRTBV1fnhDJZvtL4xBj6eJYwWzDoKUDpcegW
k9l409UpJGqwVp33u8lboixtKA238uW+ul87a2oE15phUvHPX70xrFE7uwTz
xwOXt7gOCHqtQyzx2/CTztXmu+uPFmpRlEEiVuHfT8P71jad2bxL5uNQ5Zez
4H9d2h2id/zw+/XtoGzaP9Kbpu5HwmriAcwPw9F3WYph/YdA2GYt5Z22H2Pr
xO9KTEygTG8SYKeuNyHZexx0d++PIekiN8V+1F5PIkn0ZeETM/qxgSEX1Kd+
x2uBJKWSw1cfwlzXWef+mshf2CVYigKT+0LNN67rqDA20tLltdACgq4NXVGn
EaulHrYKEK3i+s9uQV0rqDCQ6CJGE1dHVc3FJ2wosCKLdvqkG7fE/bW9rJMZ
cuck9I+ksy8xsaNyvOfGqKK59CTmonV4WeMqbNvgvs9WxOZA2p4tef/oq+RZ
+wNOIhKVlYt+8ClKfOd8sg4T4iqZhtlrTYi3aF8r85aSNqZXXbOJHTBR1Xjl
iBD7FhFtjEuYssNdZ+oBMjQIfw7KgGxY8spCeU0+jOuwGDVK+2Xe549/loYf
tt8Yy1IUeqcT5ixPgWIgorao3BPwMZnQBLfQ/E29B+j5NVofWl5DAlpeFU+E
RG0MxvTIP1BEXkdR+Ga9C5JqSl2xPgsJxC8JKHlIct2s3+VUHNDDcLB5IQlL
oO/oMgwauK+lRDFXF9H414dBuEMd5zMVg2NCrqI1FNemELGrnPYaZYRn7ftG
ugpQgdlMBnOR5z9kNEHzW+bCdcWTnyxI8zISGKLA4BjsGKQyhBJDYvZwCZHS
teRCtZbUc+bIe3bJ+dg6+iBAyLhMMHJO3lttpZ6HylAR+XvTt0tK9S8kGfgQ
kAfzMed+3Pkf3LG58xHgXtuKCojTfW+SMMfbd0G/D6mSmY4njU5sRG5xtRBS
8m8t+9Yj1PUbhTSyc1n9ExteDxXAd8GmIQDMtA0Jud05JsBcNpbVuoNJLzOE
mlhBVBLaQavPBlTL47mU07jO3LtpPZp2vtObAr/dL+Gt0xh1K1BT5FLqfhFL
/U0aSSVWmLribJ0ADKEKuy2jiuy+GmKzEE484UOfpN7ay38TgLTSD9bHVLNp
2Rm1ySnaO2DW/iVCDdkUsYgwDb0mB5++t6Kt3BB/FzNq8qGnEh1nfgKzOU5c
VbfAoS3fR7FfWbKNdqnD0gfZvjumsWYBKUUVjj+PT7524mY0EP57U50FLYdf
1uxHy4Agl2uPZlJXJvdJ3iBAv4583hFh2zYC9lvs7TRfjRmfjIJ25k8mZNUw
Iqk9V1uY4hADV26tI0secXr0OhNO7CLUOIfr4h8X4P2X7b44lv4hfiz5+1Zv
CTG3PJ5MfG1rGlyEoQTIaB9Rh0XXDZokSfcGbcZmG2u6yh7tWI5uw2R0AwlJ
7nPjnJte4qXboj/z5Zbe1lXIjq1zDrOIFEedkM6VpPvpHdgYouHnRNdpAubf
IFnTl5+PXGmF6uXgrT+kB+rO5HDAOgPbALT56mKD9AKcRXS1cJBNdalqnkc4
EP2LvSwtHhfw0FWygIhkp8zB+kdq/qdm4chZC9rUzgErVZkP2l7FiKmwpAj4
eNtxJWjXmcN97Dhf1ESJdSbCzyGCmupJrVZoFQtpbS0i7qBJQnGrtK7wIzhc
S34magkMrsRCZxUlPHYeV3UDHbexBQCAOYTkHhvVLao0rlIBbuYbFDVIlGHl
5NSXwfGbmV2sdpnmtscAb1jTEs5DnZmA6jkAnfmseDC07PvuYd4xwHlQtNn8
HhC50NNS4BntZAo4eOZkJWAY6XOcIx0l1xIwGEw/Y3JwRdnR8fVnOwcXdagN
VoKc7XMRlJOP6StjwY86PyWR1QwyxxK0avr6UKGL/XhHm6qG8sV4O0ZLNSgp
Fq+4eqaO1lKVBJ/JqS9VyqwRRxgpsFPY6DcJn2eBQCeRBWunsCKV9h5M6B7i
uQT4ucN1OlNUuYp86fzLHf7zV71+nKwCwV86dOtJsqh/+O7SNJ2hvp8bRiWd
6JHqSrQgAfyxmOjgDBnZbOxbdHIhSgEwTOLZwtNbaq/b1MERiteOCfJU8qzy
3k3Xj8O2mVZovyyVnSXBca4G8q+xkYzFaKEuMcJXbL3cwqQWAa4UFzYElQcQ
Gt/7KeAXjxh9vKLNjoGJAe0S99WEYkqEMFNVTPNM1dULsnxW08uVkDP6vG0d
HAMFX8gHLt3aw8sImBVjsHM4KoLuyehJScoh5otppkSHxbGXFK+BxnyxKh/3
HuvFlJNYzaZ8RFBW+HXlNoIJsWg5eTNI7Awv6d5V/v8m19VgJZOX3R4u2WAt
kWj6CfJBq38XXdC4+32QbTlMk8S/VQ+RtpBSkZrKspsSR03D7whKjjLqbnqs
2HwNukwU3VDh2+sLvumqfyxyAT7+i0vrcfYDUcFgsHuQu38eEBT8lrZ1yPFY
YbrbE11VnDOgZpEs8tAZ6pigMNGqA/IW6+dlDsHSiR5HJxm+8oSSeqcdndFd
89jLKQsEABMfKTb5JoblC2Z7Koe/su0AuT8GahG11F/5ChkAGRkOYpUMSPt6
STgSsh9C0JVETJIUvzzFDPJo0NUuq0IMqxOQvXFoAfdw85PiPTvUSjKs/VnQ
S+W5cQot1L78mT9FTzOr9ppTof6HmRkxjLxiUueBPmsWD0f0/cfDl5UzxYtK
E+mj592yJqt4ELRsDPPlyqQn715I0xdHM1GliG3pmK2L+40pcerAaabu49yo
eRZjEcTxUXCwWsqAh/B5wpkhENHwM+YS00mR388WnxGe9qxFOA6BvNsB5geE
3zLZwJtpoO1tWQZH8hbg9Lb2IesgNdrvpdtP1Sjx6jQydEp21M8AZ7u34YMK
YTOZGDAT/EasIKcoZuj9snC5fP5GQIKPcg6Vxv30CS4R7YhvuIafskQZyRsq
fQ/Zym4eophp/OL5FdivO8pun8Yb76r9IOOSVgoeQyJeHaUiaG24/x6dmJmB
essjuCuESrVtDC62+XCAE+YEEgBPxaLrrju6IXEefoVjpYScBXyKS6imR7pG
devlVq1JcPin6HXS88T7kmCJCUy8d/ChWmwI3lLNMnEvJqOEhGJ1YkJ7W7GC
RY0jB8wfo+xzV7Yi2nF9Hcg6Bo9EXFg+JL9Z7DOmz7oCnvdzcUPROu+a9s0Y
Pi0vqkOOPE9/UrKo124IVeR1fIjleimK6dqovGYM0xvdBEm7tL1M+IWdbtIA
N/lTEfBLVehwhYmObAuecdFztgqbivpWSSpfh7S6XXW1ySfMC4Thx7rC5voM
0aUwwpc57mwxzoF3a7h0d+5/U6HpVjgC4z/Y8J1MEepxo6VF9DH69IB39OcD
YA7b304m+9O72ndKe1kxsNRJvEs4ermgWqGxJPwKhcwaBx9Prr/G5LCCrRD6
p5RNf74qr20lmSE9+ispqJ22dmz+ZzyprhyUamNCwPytXaT2/xZyJwcY/wAu
69tAFzCKV3Z8VKlUaz2F4DVnrH6zl6l0nIcoTgi8OkCV7eiuiCYeyOkWMWiU
lKSq652B18LJEQqvbPTrz79HKuKU3QbBgvpZik4KBCPVrgqeCgZhnw2L0LXP
E/Rxv82qNz6PHDc2ko9FRw13PlVfl2+xZZzpXeUl8LaGi6HaRVXT9ERJU+64
zbgtpj0eCMkzoNkYYIC9DjF/L+QJ95ZlrYakq8kng0/2CkN7mwIcl9RlAWQ2
IRcai7aj3C5swR+xzccP0/QHTLqF97e84KzhNGdfpvAub5dFW+q4yJ9kPk1h
2H7LzAc7BtRcVwmWNLYZAsWJdUKCkdHQkLWM9TvW4Tqk6OmVhhWiG40GZnJN
lco/OZsFlQSwNWIaUtit3RM2iG6UPkWyud9LQFeGjbotsT6cPMYPwLm3866O
Wzu2qLE+rBQNh1TQ5TfZ0z62gOMRDl5r8it0k+Rit18F/UNk9a2jFWgB5PsI
6vog21EzHBug5IW2ky+HcTFsVxhJdvuIs3NMXiXvasjFGWoj0dUQSP1ZElqz
Au1dAOnXGCsW0DTbuEbh6b4PGzKGTtQrbMXJwg4/z8kFO238Big9zK4DrS6P
iQxx48DPY8yCDCJ8H84Hb9qZ3vZjW4TomBia/FLGXePQsxED0rUCAQQBOnQy
GH7lSTykp+PLsqXOKFIneo3vzoB/gchso9WbqC9zsLiKz5uPirJXu44yHTx6
Vm13eKZpMrfLm9LNoDOIEg9QoRxu8rDmMIYo5A5O+pqr3D9Pnqubmq6DtoM9
aCHrLd9DIyAsF9iPqWm22JAkRnt50b9D+LjfXUvjabgVdOVQNtR0ppFV4Qzk
r+t4BY2Thk7Bl7f6HUxCtFtABcbe3ZmuHOo2jI4uStS4A5yAmFzIawBWkJ+3
bhyPa4bigV+jT3NI5r1fZqmWRZqYEg1FZmlhnZ11XH73leTxDONOcNCDf8jK
d/9vzJVWuOxs8OyBiuPdL5cCNzJSAK3BH//9H0xD0uwr6sqxj+kbirddXlvK
PUtBe4YA8HKHGACxc3mJd68vzbxPsROGsWIwxIYSsapMhl2f/BVoksqeiuBV
mIZqV64kJQoCaHP7FksEfpysAriaW9rzNtogn/X4dYI7IOCuWUXpomFYV6Lt
z160+K6PpMqLpq+4LiU5OZaoLRfqWqFI528EBUxbGSKUwvgC3iKGDAgsTcOm
Ifyv2Na9Zr9O+AEdLdK9+9rVNQCJeS9h+wd5Wh2zxHAQFNKZLOxAd3jHiLe0
hhjGcBe70Go6Xj+Gga3AiZNqq3KYJfk97X0tUwwXuGEY1iHDqJ8YJaAsr/3d
FG6Nhgnz7eGOR9JlxhCLewPGMTHJOF6ttbPjes90654y8be8Udj3v0opws7b
uKQLU4xtRIXTS1dd2WihjTnV7fBix+2i5zhzQPxpiarivfwYhnyR9NZTvRN6
PH/CBVCS5RpLLifkF7JRIbv5M875T6KxNwh6uxEI9sck51lzHJwUcljoP0I4
fJ1RqoNga0i/ZtH5pJF2Mql90b2NrbdXb/8X51Y73ogcOnlfizEEwJC2ECFN
iiHEEgetrsilrYxbwiWpdNv++nn87NOkhhkjtmXdV/NHSZc0Vs3wSsZFDY5x
8MZi2ncrk9DAme1EPqxJ6SU7JwEl2hYNQcKYF/jhi+P7QL6ClIsZXfCAQYvC
uqN+Mhvc8rO0t5EvQoJdT3R9UpWcRugWr7D7HUaIC63uM3J/Tt49x6J8spAF
lgMgp8F4aOrbbZE7Ewi/IReqS72iMXNGuZ6aw+xoICFs3+afabh26mGIyKPl
3aOlRwi5J7Ep4FpnIRUH4ZLBF1cjXf8/rkUFUuHE3HfXrU8AypfFqk7zZBVr
pD6axSWH7v2427ygOnYTgi3i3TdwW+WNakN2PoR54lh2WmgH15/YL6v6rVkb
NKDJ2Q71fBlnFQScg+MZSsz65U/qJv1Yu1Kcrvdcal4fRMu2Hwxd1+8iUM7B
JhkWGuk/DSojeIIEQ3qalyns8U4qKoD2mFnIC/GmXSbRHu3bolek1uPPvj/m
i77G6mtSZwFxkdEGFXk6V/cpnBE9/06KdwRkfuXw8PYXGs2TncqzNnCM9yRz
LF/quY36JfRE8Tg+cw9Wv0gpVeAeHO3ABMg2mmda6Hv8kqS98UoMg5KBA3Kz
W7EkPxsYO13LCFAaBnRKCl3tlvSvNOqLcpWo5dgAUkjY3UujxiSh4m0xYcYx
2t+FvuIS6g40UNM6/gC50ZULWrL8qdm6s/ROomlXwxOsCCtf3uJubyfFaHDE
9FBXxlo11FwKBUAi7kC8yeBMLzq0k/bj4hrx+MBcnKqDi53yPGfTYQSKnQuH
OIswvDUIhp3haF39VcKCd4l+DgpaRCLCoNjlrvNDhc8FMCP8SnDu6FRhIDlj
IPBzUhBQ4Abz8ffL23i9MoIwHPWCc/DQ3qcgKKgrcpMUE665unza3AfwkCjD
1iNkWXXKsyQhVyQRxiZw6Bg1USxAAqQsObUeKT8JJNNkQKeOczt+hfh4G6wC
Mo9uEXJD4wOng/kmiJRQTWrKr9y+7t8pFOjwEJaOce9DqbBAoSTAhYU7Hn0p
+3mLc3H/C/rMI+jNFKMdrdAp01kUq20L4XolhlEtzDbTqTg1S/ea2uEunk/t
ZQxFO4o+q4+blKLd+bmUfrBLJ29/CIqIo6XhSIQzyls/eIdvYaw0xL4x0qGH
zcmhYxlf5NALm2My0L+Papm9wZUkNBt8c7WBJ29cUVKr+qL9ld0Wi8kFa2jk
/u0Wr42OnNX+fIDAar8RqOnFMeKzNXUQ9V/bs4UUYtTPVQcJscVDvavWkjfW
wvTV0b7Qfb1mHhaO2Xu3p+X+ekkV/Z17gNSOyr/kx9yMCe43XmrLBtdYmDzc
Iwnj+qEqUeZ1pyhagWYgzz99ruibK5+TtvuP5X+cNhs9W6OkYytAISVktpUi
7Zn6vEPrihbrUjEjxoNoS2OanlODMyD+E0dxgD8yPxjj1iBakZOsNzOtQjg9
dwzREnWZiAsK/bmlbGRXNjRgj1mnZiW5SAJhnCc8cfFUh3JJokoVtXRjngjO
4qQrRyUJ7FRWI1uKqqHjCRQArOnitkDGSD/yr8VCeHG/18SArHWbHBbueX7w
Qa/tPINDW6EBSqxzO1vP54RMXuO+ALUR0clBAO13vJq3X5DC7MDOHNKX8z8y
3yaLLDcjC1RjKCHLtcOEDYRxKors6TyLJd/vcOVsNNK4KlOEPpj5VdE55lY0
JwEVL3UHlP6zXQbBGqdmk6zwFMG74EiwNyxXVb3QMfQz7wj6f5wEbkuQtf7i
WIchhXM5aETDPOHyO9/kBRSCDIV3MFrDvxCWoR5PiPcq7Yj7aqoB8mh9rYeP
JiGfdwhED5CQTbwNeL8CORb7+elWfMtBh+L3sJVhR3+JP4fVGJd4MDduMyik
de0RRTBCnG8E0QbuNsRx7clMmLzH8sr1WNc1kYDjw771BoroHzCWdDYrS7QD
UjEATjzX0DloTCLXRVDeahRVR1wUNQGwApoIcyOmF2/hWV4IL4M78DQhkBmK
vGUqJGocGoImbQg0u9flkgbGRhmcgoiOlYtHsm/5K6oSoYvRCRP5OZAGTHKr
/Nxzp3UEahZRQzOKTD3UYMHLKFSK555I/C2OpB7OtpxL7kRndXs4+UawxObI
hAfvP+ctjVYGc2G0KtEj2vW94leE14935bUCvxeIBNuQfYoUcLiVjPLRoeMJ
ErHZmhut2p1m0zg5UoT5CyKMUoUE+q+DdWeEY7KUeDyWBe8IeLnmKSZV1gfC
ufo6VPFg7gv5eUnewe1L223mdxBhcnGPsYDyjarOcwTkHRg0TzMszwdrxGlY
gRZKwPuYpsHCtokyAr82jKH3EyvnqZthWWg2VyFt6Qe+5yRrOKhhC02tCH18
sWlkWwfHR1mYNylRJMR+sgpb2wKLCuQv+XSoh7eDrL2kHQLq90ak5chNXqTQ
60+eQYWFHJjPqR49V45j1MlW9ZKU5dT5v0Cxmqx+NnPJQmM0j9ocvFJScyXQ
jtUVp0aW19oHqbxvWMPj8yI3p0Zisu0LCcMKyF/7NTTt1AotiNxKw36SgJbw
qpFbXc1TS4G5zQfqbNN5mULjdzk7/Aub9Ug4LJ0Wqk5m3z6PLQXQK2PvfxRS
BqQh2Tu2ZBoQhkrbYWa31KmE+m9BKioTOfywlUhwcoCIVC0EGixJRYy406Q2
hSmMlLSIq4RRsF9psksPSWlFvSpu79YIehttLTvGu6El0QvN2Or/H81O4SZL
mfISsqx15CuCKeu2KDCdSECcINsZVvBrc/uw/WtRRdc0VPwbObUSDGLdJrLF
IbAnZ26VCzQTQhHKTRN15Y/lTmy4pk2lCMRvqT9rhGW9h3nyrqBI3MoQ1YOa
TqB3jVc3c5ZPVIJF26RtkSOQP+OLw6HjKpC5pyaExvhQC8ZbpMnvXAL/xvDO
aB8kx2Vc76sePfs7o+cRa+5DsTde/3F3s0z3xCKUSUqC8PyBcs4EEBqqJPuo
OxLZVBz6U8AnIHlTSLFT6Ci+IqbxrkH1oC0v9XUnb+c2FtUk3HoNXBh49Kd3
qnpZ63+wm8zLPCIlid5UAdbt7d37L7N6Ezvta+1fnbT33sFcjDSUOPnLsAbQ
Nfl4/60Y9RtNG0rNtBT4vBNPW/EOxjgMKaAgQp3T4i7lf++nYm31iJGAGBFU
yOo7kCy7/sF0ZHOYo4PuTElHLmJfNvVAiFZ6TtuD69ZAkfsl/tcFPV9mB5OV
bVKki9FtCVj9w1cVmDxpbDtxkiIr+NLAanHleUNJOEH/opegnJYIWcLp3LkV
2RWtI2tKXW3sG5DWWiubGE1CnKpho9pYKYmVDfslUPRJ/+/k4mWuoFHLlsyq
bDkfVA1Ejqz/MSvvpVE4k4Zu2xIA5sxCoC+6ArQNB3hdyf98W7pLla5s5u09
VoqFBBsAULrM82TNADrA3nsW1kraJbmcASpYTSmnfwBxNwSJkQ9R2RWgDDtV
fjkrrr0oHP2wxh8voptW2eX6D4p8ORLxfIz33PGWlmyKor3xvoVbeUWAnQvY
kfnA36EKm6d+RItARe9aJzehpjgkj1TqJqGV1TQAzFedf5GE/FFj01UsGdXM
tdP2ErY0fh0g8onlx2pIgOK/GO2TGlqC5zH+nq1mXncjqXY2vK3DdhE+e108
bkwNd3oDvVJN8rg0grd0n6D/GIOTow+i7dwYqE8jyrsYW5/3PqRwDHUHD5sx
wynTg7hj3VxPoF8YeFBZ+jU1568l0oL/TvoliH+mnfV0nFWMM7Tz41Cqp0qu
cTWl7t7tupJf1TIAUWiZAr7qWFwaNiwB8BtdaO7thfZivtonlHz7mxHViD/t
8n6yf5No5b/J1RwhbXFP3SUzb97OTx3sYunw4Cqg7wDt9jbcR1VjranLRRcZ
Ww0Hnf078TFmsfRSKsPUMtW0fUa3KHeUrkg2M5V7bPEiFJJV/gpDsL2gOkL8
uSTkZS8JrUS0U9jIW9WHMOeZhwnU/OQI7ngb+uzHMCoLiVtw66fonPxDB7CB
og1N+A+YkxFs5FN43Aw7R5TDVsGjYeq8PCZcnekeSFyT2CCGG05xHMFVC3ww
gz1fgM99M0bNoBHlMLgiJsg/XfX2NvEw52CWe6zyS0bUYfg9xmy6zEgUm/t1
g4hWACBz4M/+J52U0ZcMf/vgo7ljjRq8WO9+EdSn3qiyGkiE12zextDEYsQO
eA5Tkfl0kOclG/qy1tVPcYZ6Sqy8aTa2VwY0qMGTP4t845Zii9g1YyMnVW+j
R3AS/GUXHV1/l6/vfw5xtCXlVLPCIE9htc/gMnTXVnYkM2iGaXH7mzdF6gam
5yvkN6Hu+KclglwOVpxy4mEE7+/Sn95GR9oHwNqv7dmaRbzLdDIaqrPMOqdw
53UyUyixPsFd0JpzsduHG7zrLY4PLBPknTPP+bLHKHzzQyTSfN1a7mWTi818
NvfLu7PErX2NOMhHBuzQDQO17rIksc5XZfl8TvrlaRwigb0M7Z1HFs5R9CV+
iEd+J4Xqvnr5OeBLO7I+f2CwFsSXV4x7cnPb4OH/zM1ULQifjnFDB/bNQDfj
HJzZKSNT+5wWk/yu25Rn3rvxAznMPT9rp1+3ENuSaPgvnQCgP+qApDhSUKV+
OqGz/JAJHTJeBaw8OSOeVuhrQuNee/Yw3QQKlBu2PCVooH146WZIPXxweSih
V4XjMLZDJ6hQIRggi3hctk2cv00zABpyEJAIQrCsZm81AEJAg0yGv8NCKX8T
zqH7/Udy8QmC+EoNXk+AYesunzxl/St4FxVbVY0Wl+tjVHj3bVqsuuTQd5Ft
+X2mzt3lLI+HEZOL4xnqysmH4vtV3YJc9/XeGP1d/CtyCPIIRn55Vkf9mfi4
xa9FBOtJM3l19lRcn/6JRr0RqETzZR1JodJrv0GZLmYftZqb/Td6V0aeNF+D
K6ynNsIoOjz5n/gN62gbfhJXwL6+3JW0saw4OsWFABEmtlU74tb8FXps5RWu
DTsv0wQiN7FstEYpwkE6RYPoYFwcilTW8qa3mnIVZXM8d8iAhsBAQHuudeWs
biWtZMWBgT6D8lOuzkaAPo8dvBwLiW7cT9po5Pgds9jOmAN6gJHNOf5dAArP
hggeVGst6RB/0p5jSsBenqbz/ypBXlCj8FaRnlVarX5ay4XueBW6iSBDsDHI
oNCxVj6OILKNrj7U2M4K+QCSN87yPKN7neTnOL6CNDtSEljVZgY8nzGmb3A8
sP09/prn2QyQRvwoF2sbtruhY4rkJz1K5YdHK+EZGTEfmJYr650Loo2Rj6H3
/ZwJ8ZBbLqVvAsh5uO5xzhm2NKgfBNadzDmNjT8+iobasGugBHGpygfWeQBQ
vToGFLvRFLPL4wONaPUYKCv1B4r4nJeB6i9fk45KlwCIAjIALfmXZ/I79b4u
stwtBZT47IabhZ4f6gKHiTGeNPOf6ZJ4LRkoaZpj3dlFnx2yIZ09xWDdZ6OZ
el3wOpW6zpR6FwFcg33lsAOibVyqUtMZtAHwdrwwnFOpVaLeE2NfKbwHQjB2
RQ+gfScBt23l1lITPdfm9+J2F93VBX+wFhfhaVniej+51Bqa9hdxqZj2h6Q1
6EY5L8Y6CzZ8qoOrHrBEWVF8QX0lux7yiC3la0+KbQhoPm8zICZRMUcu7Am+
hPe2eHB5PmlahyEuh/54Lc8J0FnFpu1oS92Gt71Agi6kSjlWKs8W+HDDcMmg
TJAgJr1vx2ToyjO+4J+c9JIODLfUuEWlXnPJToqYiI7Oo4OM2KC6kJPSjJmt
MlCEVUEtF9cN1vqJ/bBZPQnHBQAf0FW1s64Tbjqo358xqVtHGVQuVB0Be/qz
I/Hl17nfCeTb3m+07mM2sO6z/GqGgxb1U4KSlNM1xVIiT7v/TikpqA5IC8lt
hL6/J06vvR3cUyZCq/owJdAfoOg6/74yR5kFR79N+EYprEmFmLWm2+KZNl4m
6zcJVMZvZYX2/dz4xT2TcB8PSismplrYwutE4hCj9Ut4jcHn2WQ78hnQ1yY7
bcs32otNPp5yg0ry7mTtgzaw2OoGxA4LhNQdI5/PGy9Jot6JjMLOgGanHX10
TvHp3xxJ8irrqdYeFeG66YmtSOFdBZ9nlmeEBMQiQhBSStY8z4VqSY+vJXNQ
dGNFmKUo2O7k+4+j+H7nqEk7KuVaxdMlJD80RPOfLX0bMIX7eMz9YVUW1plX
ERg5OgeQ4hOysjXZZBn6CvCLb1EmIO4USUyjoa9fV7Tssl9YbUCZhvJRiY9O
/VYxhd0sisifhiGao740Xj1dg5/zLdcZ7r1FmZWbK3P7Sk5HrPxWOVXan9Ax
udYYxIGEEkSR851JzClgKufGMrgdgcncNNhvayqWW+MafQb1EtjTDv4EBOt5
XmsJGWKlZLNB/eWkuBQtoqxEP0O2tJA9VdhVxVkqOApmcL8ojY/bkhgAdsWK
zSyVhm8wbXMcf9ntnR7TcEUNnwG17HyOnZzaRpeiLYxIb6eBFLZCh3E0dV4X
5hmdMIRy918Efid+KTpdWRK1o8kIyxSez0fnPaCWw8pPiiK+ykJNJuLa2jgW
L8PwoR4u94VjPNNa0ERn8hraWD7+fBX8gJYCyPCxvovieg8mZg029faXsjjP
bB7K9JCnQ3+8mW1/m1mjvu95LJyao5XYWKkKarxqT5mqvcBtpujNCUQsXuXg
keQ43ZaLxPmVzLCchiDfgOwcV+fwbrLzdZPYPVdF9byzCE69He27aIGGqgvt
A93U5+2/eWOSoUJdtPkCKVMd1PLy/1mtXKVuOXDUJqibZ2g6dHSVn5IdAtEy
OwWkv/xM2xE7xnt2AYeRGN86ZwInhfRlPLCJCh1VzbQdySm0t8Qbjrr1LIfb
LRc28mcfnw83VprqvWxeAi6F8JAOfALH2LkY8OzKcG5zkQJ2Gt1xQbASGk3i
hMtmDMWBe1sZTQ7KH2ZBaaZ5LybwCJR9ZbtpnUyEITqeDnyEs5ZXHg/T2Xbr
FFPMj0EUgCc/dFXsTvGU3Z3E86ELQ4Gtjp4hW0En/oZYKoD2pwOguF3bTKPs
QNix0DXHpbljJ7CyP/1I8hNesQ0k+/fLTxhRjNYWA3WILL3T74tW5T7UaF8t
MZz/gRXn0esKvoCzrWuRQLXRiqi/AMRuFMfpuZb+2zO3rzx9toGstRQMx0HN
rpjvrzlrqAE+v0iUfjtCKE7NXjpiu/sFptEiXsMTPmPPilcAfEXhjwo9P1GA
FTyNXiAA5Bz5NnOrTdZS7/bvF+944bhwMqglZXgj9SEkm6VF5Pjp/b3uA1wf
v3A9K1K1ZEEHVFcYH/xx4rucpzVvYGGhKfwdFhWQd4i8rcq20V/09atXhrCc
AFFiKQ0Ryat1JdVvC1CXN0maJIzd53zL8uQ1rYsS3qDI4IMY8dpynJm58M2b
qEQzqwNEM/dwHOnw/FpF+uNtz9vrfoGISSnT1jhJWk8ZXGhcv1lwa/iTFlC8
IdX0vpxy6f92kH1MLQGZVdYDsvDvnGsdkJCi8yaTuy5XoNCkHMT8DQgbihys
jJxjNwga0b9nq8DD4upCMombSTNcCKqwi7yzZZ51a/XS2/uRjb+/w20BVAG4
5OYBKKCidSJMS8H9gp5YuiJmz2jFrcdrEQA22NZP34baXSUhFnb0QRvUQ8wC
SuZqGYejlhM2l7RjsF3Bg88DLQlTRW2JfejoG1sDvAXNjYhLWi5KKFoJ64wl
tN8Nc1EBuHuq8L/dhXaw6sIOfLSIzWFMOJLWr8tHqaKGvGfc+auyaTlhvlWv
h6k3wwfsxL0oh9teiYrpNpjk6pExNKcKFXVMcTCVuzVi7UhzwNjSlUhOsxmC
aEnGwthVknlP3hbCFlg4OdoHlPJROteVmzEbUzc0+DiH5jWcX2nMZHwUiJyk
Qs69igCP25lFs07clMlY+IDJ/07zEzXlBYB9T36LKNlb4jTf7Sbw9sJBnl9b
gRFEJEzj24g1fwWonhEo2xhP4iDMBWW8CNukGQ5tI3LCtOI+qLHb4+PIdWky
KO21FU0zHKJoJVE687ZjNPdy3LU7McYc28dA+d60XPinN5AWB115QeFeRpxR
tj86jzxhfCFPxPfRotzq+CCHCalStDGZ4KIzpxm7iAHpTyHK3QpBNUVwOd6o
PeMtsJkMwajeewKTllEzXXiP7tVAnkr/atoKZbN8KN+/kk2hsELn/CzQeMfM
FuGgbAKvVK0mUc5/fVq5URub/ZzizZZdJ1jfN7JfWF5FXDHj+6prQ1/FfQYJ
AvQ8nSe/HcQV+QJ8Pe7EpfHYVgrtK9WQJY7QU4HG+YQR9gMBvuljFYS5FF6j
ZHluNUnK5ewxIPS1BgFvg3qubclFjrdZAjBQQHBvf7hPEti2svJdYmf1iSdv
Lsv3caK51B3zUZ73eioPxDJu28H/NlgvwNzlnnC8sHyha6FcZUP3XqNHypm6
/dfLU0Sr/mQspBZE2X32Do5+LlSPJwXye39HKSHH0P7LzWXIUsraIvu9mWXi
49NFrIJBm8tVFtRZuwuNmiHR6sZb6mpUh3xAEqf1iDYFr8sXuBih+IEibBkb
8kxZ62/NFTNpJgOhVknZGs5YgePS67md9JrPPvHtWC8sGF9iYz64ATIzHJZq
JoQ61SsoOlRVW3g8pjVOXXJ+a3Pbbbtpn36lsqbckq9YIeVNwAKfTzlW8gKe
ISJ5ISJVIzClsdqp4Z2N3k9Co9PGD893JzMFCaEiGtdqOIVMRzn5d5tzU983
2O8dd4vtJjb3q0vDcIIXUELHx6kEy1vvmifY4cXSQxEAFNIskAy10/fD8cbQ
rq3hCf1t/U62JkdE//dO3sSRXfWoPVp2MduuFCPguW76lUrkeXsSA6OMESaJ
wsN2FroCla3VZdHQ0MpORFiviGGtAQJsrKk0Q3LwBpzVFbdZbGqYpKcNvNbf
y/mbow4FaMBqnDO3PHskuV1JSsme5ZKeZrrZ+N86BRZDksH8ivfF6+/uNMyK
/XwL9YxlguCm9KrwRbdUVUdOH5cFkH7AP+1ti7jREwbU0L2PNHzVBdHWRHzZ
yTOnVunlqSQdYNeO2W+dbjylpM97jbWmwBGYbrKHaInU7ABCxQN6qUlJ5zkn
sgqsPPennJaXKPOYjpALtCONMUf7GMnJy2KN3wTeOLvMK6WyiC+q74VVQges
gsTTpUqEQYcvqwHN8nXghwNXmQcS1eV69Bblng0hBFkXsLMi5WoaqJl4aPVs
hYQryGKOg4GNa4j2NdG7To9CXVpyWh2lg6LG9/HTlzv5AZ2AvyXDVXA2mMW5
zCvY+R7ouSKcGKM8xPLvXioetBcCAXz2JINAfRzCnBvG+5X8pGmX7uucl+Pn
rQl4uR1vbh/mxmrfRXXC2an1JW14s8MSx5cb3e3txMENEi6m22guCZ2J7Z2o
aScDqQoMvbS56OiWAQfaHd+kCqF50kE15gw32+PukVHx8onPjxjXn7W1z0wD
QPgwrtef2n819xSl4rDvEoXviROkt1smDcKvQ5x6gIO8vFjzH2Fv0QQ5ZASs
1pPsP/7AARkP+hlgiVd5AP7xeEU8G5cWuuSmmRIm/zRBaq/2cwk6eNDsZKUI
bB9uI/n4CbUo3OAwH8aw25/B4ROFHdyIkM/CLIaBjW1HXz4BQ4OJSmRgm+e/
nGN+aZ3/JEmtgXFgm5uycv3XUy8+rTepgdRVY1CYOXtjDPqjUU+xWPi7ejcr
e5UbnFN3+Eff/qt3xvO3x7Y9i8188MBag+rTg7my0QRgAE0oq2qzZBD2k6Lm
f+zGzOz/BvO8ZIjbxZ21j6LoN/uZu6S1sziLvrd1jJNqAO74ybyI185e6LIR
RmGZ+/tlQ/mqdOks+AgnOzZT+jRkUwdo5ajy/fMOltDuTYgTaDDlUSfVoti7
gkIhIvAn6CqCdf7Vy2liFevmDiHhk2v4QuKNIFp9wmzrHC497LRQm/5fwXtW
TxsKCBrOJ3CUPz/PGTETu92VP8RacIGeoluXygfmgxj0dUkpIjSpWmJs/HG3
Sisok33ZdciJIxfv/VvUOAVecYTSMT/CaJZdNmjkxE5mafKKDNtKy5fOb96h
bnfuMX47Owij71FTmGQ+F+Ncu0yXD80vNYrj9eeW1vt6QJMFIIY40+fO8LPN
z2PT7JnRfsk4Ca9damewNF+ePDvUxra4QEBCCEE7Miv8a9sjCTTen0C6ykH5
w6zgGNdM5rxCzFAHVEAdSZzY/TzKQYJ6Mcmt1fO6yGEg0IawivL/6GImq0EB
fPSmSlyclu9AMQkufBlL/TAwhVwr4UEOFP2v2zKLEy3HRd93OoUwWjtQ8qBw
IgOBCmvbUOyYjvJZuKSr4jDk9Kfi6C4Umo/h9Jz+rQn3gTvhaF5OEpj5hxck
rPPZwV1FPkh9hVeL0bRH1HQVLTl0Uz1l1aU+uzYdK+kAX1Oibp2MBv4NLP/O
cYT9kJ6mgb1VomaZBf6/0AfWBAfW1FZwWvxwl2bdf1Lj9SyoH5azvg9psnZL
PW1Ww8dWhm7KJ7jlJRlSDJNKurQTb+XKRrATHnAw6atqs/4SLOKxfJrp+rhj
XbeTYCgoLPSB/OWw16pj98jD3oOXUToNksuz1MXpXMgEH5/swEGcaM3lI4wW
XgzzOky31QHqjrp2xYZilz8ZyxOT/xIaVjf0x/m1i13mFUBcMcWM8o24bWTf
n7SlZdbZ3zH/YbyoyQXPwX4OyUKevloO8MgUHGVIw8kIxfFOYMl1+e0RIyNo
cjNRjyZJQ7tEGiVPpGtCbCifuwU/QLakzJ+QIew4iRWFAn/+a8wLMrl+mHl6
QNg5y4FPXfp87abgHTVvu+TYjpPXY9le1HwFB/seC6Jj1vZwKvNqHBnurF1S
Qvw31E7d2pfWwO8nLDVHH0rZ5ci+y7GTttKPVrDUT93fjqicuer50PQ+7D+R
jro1LLb4rvcDx1iaYpZUPYhDxKpfBZ+7XiwIVi31sAClvYEqLPui7UG01/Wz
wXtK46tubb6cxpdPLLf1/edkezMcM4xTQsaoRn8QlnS8JhPpdtzS3LNR/opt
PlVCg2LkteCs/T3OHLcIaLlOpZO9yhWvNxB3X2f3nbBTvAkQpSvIxaIYWRWT
VIz6CdHgZrkvm1WpmzmqNnI4OqMMlOeRo1Ujq9EP+dmaEDcXpBhWumAFCvAZ
/EgWWsg+jZNHIP65XLz1XPfMIap6McN26WaGtKy5yPSs3SGPfv9aKPjUdizp
0xTWASpTQGnkcZFJ5NfDdFrP7TPDv4UiYtz4NduLsjr8NtFs1M0/PFx/QdhW
aEQpfo5nk2F4UybgMqyydkCQjzPrjUU+58+5dxrsFTvHvHGviDwdEDYmFz/D
S+8ji0rGKqlvibi+8y8oBU7SqDrdybnuHhYnFn1qhdxPjTaYO8g//G+VQvPx
Q3B6uCba3XV6/USfExWBgs3Q/WFloHW8dqd/VNEtM6zMt3BCZ1vyJX6hnkDQ
AfBEunK7dt5NhaBLG+gwa8tguM+10mDzMny5GVmNXULLwOaUKJmnUzOkc8TU
r+IP6vngdmPUshLrn2ysX7zLuXVd+RSfm0BVf+kxGHTh1iMcc6jTTuuAOeHI
mpRnM0pmJmB4NyRDwcauFE/bU9LPMaAbW42Am6G65Tb0wTkcGD2sgQx7+3nA
T3lLsSmxKBVNAhMPq42bo1S6aGkBlOqOE1IgOwBanw5SZ3OFg3vQ9g6M16t+
KTrxjvgRZhXdVMPvLWqbsvYr1NlU+eGVw6nbPZwS4KHRq1eOcJ55aoeg6zow
YJLYWllFIwixUMxc8ayOmbcL4MAS48hG2Ba93PXrbsR4EF+36aX1c0NUbRH4
8wmGGy1QzhAwDKiB3FbmcFmpml/C34k2PVZl0bjcOugFpJpTkyKOCdBqRBu6
vUyyN3CLRC9flzpv8rUlAHDNIGqL7xySnUd1NEawW3rC/Yia1loBm7uzUxsU
Xr7FBEAxz04ZfAN0GPQmAaMAQtCt6vNWZVcTcHDhcJnzwKcvoRDU9TTWJaTq
06cvLGWxOVjESu/E032of7M8wSgpZVUWQkh32fXjKqpPd48h2yNmEp1NeTQ0
MtmRhh/3+0DAPEplkMyOipyW22juAY+c8Op6+Z4zY04MZXXEJqmaHuyF8XcN
IgeFNi4dgN0vqx9uzi78xa4NMWtiB5C4PoYrllMvbhkGQDAhkprvERU2NVNy
WepTkup08NBJ/XLdAI5XEnlq80+SRghek2+Cujc5XBDMAF79L+A7D4wziQjW
Wxheakbcz6huWw8Zj/5+vPmxGcPPoZOd0oPxdUcWYWNDMAu1EKa/R//b8MHf
0aaDRQPSvB0wWcosOWX4zV66APVhBhyagCr1U1K4UnGJQO+PX7PLNHkf9Nth
u0tgoFqAJke9trMOKAiPiREtBhKvgvyS3xLOsk9LbpoGEtC8UrKR4PvYFzfK
iqdOTSSJCvqbFWJMRm/3cINJQrp8gboED8HGPLtAWa/VBGWTbAGvNG50VLf/
JhrbouZuJ7ToCH4yFkqWhd9muBuXhZZViyZ61kDGKiZ0mfrnhxP1RSCqhjOW
DBkJhSBsTbM6rFAHwlGyQD6pgm9PqUf8NbVXnqA2LdQv/nYePJIjleOWZtZl
UNBqVEEbiGr9dXTTAcZM9wM3ZMJs6L0Aerwq+HNXJQWdKZw673fXycr8TnAE
KeIuXwSsrcHAQ2WEsyVg5nos098CrujaftXojXdGGfV3pjQmVZXhIxs4wV2P
NUtek35539b6i9d6LmyVjDcmf7WpquFYavKDzzwAbmWHZEHZz5OKHTS52uSz
9F1DfTGcz4lbqVbQArYLFjqhIlpzgA3X0TPbbyIxykysOF9zNe0mvGGNWApv
PqoSyLe7QTSFqbMp/3rHNumv3eGFj1IKjQPCNyQxLpGKLBFWI1GswEYsxCMW
IH3UVwMHoRkGUplcNqA+aTtK6gGhB6h+JSehlZwHqg+zIxpzKgWjIP+rI7S/
jtDhOQ15xc0Gl1HwcxlsxK9/kMJr5FCUSPxceNWGKPo0BWkA3zb/i4J2I5Ji
tG1q8IAmCJreJ2zf2O529YVlQFD9fk95VdOoN5AlFyC0JaV61nxAy7Wloy8e
pnOwN+BhTXorfHOGHS8Rz4b/2ve8rqj25dSjFNjFrJFfuynPqwIxbd5uuFDk
vmUP7EX4yw/qFkh6VfNSFtJZErpl6LoqLx8ycEA+IpjI9Mwb4CMP4yz3jkL9
f5Mm9jBod6UX1XUY4F76wMGrqKkolzhWsYPR3cvYAYQUVvq4n4HZZecmw+j1
N/kxDving5RgxYJFirHg4rKSVB6IESGdb4xSMxy0ujW9iob4jDzvNYWFXz1t
DEvchBxP91q+PMDHeefp9lhKC52sZvgaN2SPePql/mk02klWMt/jRx9nR5t5
sCkpvIt4FuYrB9TtCF6NeDhl1zgzZrM8kHDPHQI1lPZKGNBMCZZl+f/dgImu
33MdSCaR6b3S051KOTFoQ+pZV+/Be3MS4KlSUnfh5ZS/n5skXeeQ+UXbU23P
WH0EVRqkkPhE+RzXA1O9iXyG+R8D92tIdTp3HJlXZN2+VuoioqbNYDw63mo9
tZY6o51SCScOJAPCYVwh+07roQSd6DS9b5etUVNN/9RDXyTZzvniz49a+oLs
NHC9a4hL1Uw6yNiSZw9fbmZ/jPDLMWr+CnDel2eQcdkCRFMcIoV2b25EmDUY
K5pa42rBudah+aDLOn7Ek0Z1eOlgbAw/WIuOChrp0YbLaQb0QlWScV+1L5bl
iyBrjFfOsI1CQhWXbPtAPNyK87i096cTjr02gT5cOI4gsg2A1RYpsojht9yN
zvlmB0G1/svBKsAl5qeU9aPeik0bb+yBrWY4E3WvZeZ7MbZmUf8bfc/X2iVk
v71q0ao0XP+46Op2HfT4ERALHZGpwSQvN/JNBQgNIyTrVDhF42U3dZab/mAe
q1iJPCzmc/OyhOvYQjvZHVyQNakR0yZt+zCc/9qgu568i90nGUYn+EsB7Cny
nNjIx5inEdj6qS371pE3UGMmfCBFdILtSeqWaWHj2V3Sv5179wdSTclZ8oJh
f2IEofh3+rZ7Dx1bs9rIxRANkDKgcy0F8gX9G/qNTYl6R6WnM+gY2OADvAI9
+XD1McyVvJbCQLzmtDlQS2ooHz8YnVFoK12qipr4TZ85Ns+6qHSqAL79shjL
ujIfBy7X1my96gbvbM3bvzGGONBtwPToGyV7I/cfhoFSYjOVvQwXqZVlEaaG
paNLZZoA/EWjFr2uESYBc8qEKenLb0XQC6Cs4a9E/mJ5KMnHbruI0mIcXF8B
RzXKv/on+Hiv1DHfi4zbv7w6r5w05YDKrXHLBJBe9xH47dKnycuZ8xRaZTby
HmTu/nsTd9RY5A2kRThBGm2e6AqEvzgHUHTGXMAd+bZJ51NrzH0fRL3xC+zh
NALNLvmtSanXDZxsNwpOdBgY7iDPpOZeMKTN/L6XqqrYHljuLonchTWSST+i
k3gqeNd50vRMSUSKZZ0hYql0qIP8GjliExRLXRDFHROPeQmwLQ41t4djE3ub
bCCa5ZkYlXUCaqeiOvUce9Yrt49sd8sLLpYW8pfs07PTMeChUtyL6A3Yh1EW
0Y7cAXdMMrjGYUHASzm2HhrDx3Zd2ZF+2s+thIQCiDh5x9DcxcP0YSPvEZ16
Cy9VvhQfVxGUiW65DRfD7rymXBLmW6/q411eb6QXjumOo20qZzTn95D7wtRU
X43DBzzghYx120QSe6oHSb0WAPd/SKt2SbchbLKeaGYljmqLaaQeKIj8POQp
b+Aqdh2I6kfzs7uom1KoG6wpS2R4TEnPpEESsgkL1MPGiae6ZIhwU5xi5L+5
foCFw6ShHTkIGpKwhqVJpoUm7+GLZ7YQm8y24oCfVLSzcch3ORIOCe6RMiMI
Biorc2kC3ZTZ9CYUg1nipOPAt6LV8PJZYkQhiXtwlDty98lHBkZPJQmP9xxW
H9PgyNzCXPXxB2tiVThmHiEm0HPz3BVpqeq86w9PJVEJ25VHd8P4CQ33qCt4
kg59GVprGLCVYuCzCblj70CtA7mtw5CFuyqTxq7UEDteV/1DuCL44aaJQgli
V6R7ZP40uGW3dJJwxV7Q1kLdwcMoxf4RGBvUuhhJNDUg69nJgoYWqK3ZzAz9
RdxFD6EC+t8v5ajY/gkMDHAWI+sWDzvFwkqfeB9F0qwh8KnEkMzPmeUlSxMB
zmaNxRHZ4jopZj7EIwsHAQjx2wUxIZuMLOmI/b0XKcMZEShOFumAULOSpkLP
94vedvSNYdGobKVzkaS98/+kD+gob6b99Su7G+QF+bVvperoYAHYLWLAvAPA
RN3tmlNJEuBfpk9q53YDGlGxrQ/TIPjUU0lsWNv4AsCvlEN6ASktjZ40xOGx
sRoMeQVD8jQrC3I88cscrrW/YG+oidN6W6H2LR7DMteZRlMjOSn6HOEm4iC9
iQr42ZKf/xIWGGVoB9XqOz/kaPKdSh9Hnvn2ZP5K7zSGzK/PhQhEjT3JlPwg
xaSfT4kOmzOF/jNIPOmtdOVZnO1YKei9BQYiNzgPh0XQv39H0DtTi8cYeYRA
2c4+JYKHz2emeGLrf7FEV3RTGBL7UOxSlT/gQDIYasRUOxAkqqiF9KeN0ruc
85CgSftBAmpQi3HcP6o/rINxxsHlcyuBtUDmz8fHV5fehlK/KS3xf/mDkQH/
8fTs6mDHZzsu282IFFYfcoHkw7U1aWg6/Us0dNmSmB32VQoDl5Vuk+fTPewn
OCEj5js4MI+eMjqjPCKOhJnELP1AZ1GUfvE85dQ88pdnNCyLJJINgPIZSqRs
bSuBvLZrkDa9m5F4hkwsZSoFAFA+DG3L38jxKtCFCHyx/gtlt1Z0D5p1batL
Jl6nqr5WLOAi9i49Ygh3wTnClPXXEBgd7gm/KoJAQCwNqemppG7pQ8DJejHL
mu1TtNrxgLm15QuIV1IrJL6M+Enim/Vj2+dNcLK02Q6Wwu2R4MNLKV64sOmS
2bXXIUMsM2SOqhRy7QyQOk6rdOXOMRicCoi3OoxotHhjbPHNX/+cug9NK9Sf
B0l9YB3iyIJ1G65a//P8PPQZZUz74DlxYgh38GVIphgRZjOBuf3zEOWwxd4O
lsTThF+kDIatAfYD/TVySWn+32wGxBzFf4oXD7Bl/4EfEAnP34/GYgzKOQcl
VD0yJgDMirae2mmeHokxw530pSXgORND/R5rPe9pW7Wlle9kODADvy1EcHWU
t0UG9pwlxU5OFGAZaIrc88W1pqg8nAWDUq8f74uC+a1O9Undm8W7/rrjWOb/
t+LstECpcR7xRRY426Zn9q8E63jYhraN2vMalEBCFb+2Zzv+BB1yQjVA8lwe
Qff5wn7L5Q5Hf21zj3FWrt/AyR+2OyYVIt1tG/j/lowvVzPl/vzGjQ1pvyl5
xa0C6/nrI5+ERyr0V4jB9etXbcfDvRKrCRpgxiId+6km2OH3OTxDjJVFJBT6
OOoOGVR2ddhfVrHVl77KsgpVWJRsqB22OKX91IxQR/cAGKDAxgm6QBF52Fgz
V54xwlNiZr6Za5EHMzCJFyyV+QZsiY45EegP1jWYmqPafLzZfPF3DsCkSWsp
oAzskIX1I9oJ4qz2GrBevmlnCMkgJDECVxT4jZ7iX6fuMwTl9Zhj78RIrEJV
rSOLQtlCfwwCa0lRc4+pRfP9Lzu4k13i2CjeGnhgrCjq2BAFIMnNBrpYsej2
Bi6O+nBFJNrseqfKCsR9Sp5xqRQVhFZMU7Nls6fQNVLQHK4Q4N3b28wpOHkC
pSm2xAgrtb4kpvFJnUgK9cS990KiGN8R8cvngVWwDeFakuDIO++Gpa9Nbjrw
wyLMfY5J8kyAuij/MV0qUKq+/CO5iLe+A4RInlMBtt08FuXZHZJZ1GwcLdbj
0gtImv8nK2QlrX8uCiF2gSZj9Y5d+wnLEJMTgTt2bEtvXx1gGgeI4snPJEGv
v6mZOH2Q/TnwOXCI49ZcFU+hn4E+xj0N/q+aO5qMVzv8R0iERtM7CDsvHvky
Zd5WMEIVDU/ipKDs+2GaMM1oktzvcGaLR/00yBaJdONvjqjO/9Cw3VFxcuUq
7Fb5noibenqasnTq5/Tp8mVhSYcnYyaLKDh5KVNKqpuKddJ40hpOPsPfbdRV
6wAagvpoNpos9jlSqoaWObFfquB4Ae/IJ8BdW4+RNCN4uRRsFeRePrxScN66
8zYkvVD9Kimg27dS6DXyLUirBp0UFTtwe5lQB82F3Ipr049F4TsJlDitWFJr
apX8HVXhwQpjd8GTBlG97dJgIV5RInt90xZJSYaDYNCdMi/wjr36EgqSX16z
k+bDmcU479zBpdldy7nZx8JFGvHo4nMH7NIaIq7UJ+9ZL94TixutiIEKudeA
hVLQ9ed3aBhOg+1TDHvYBqO3dGfov2URh9KXd5ssuEEUm0cU3IxSm/nRY7j9
ebIrzO2KQoQ/FChnr2cpKaLYTtgo03IxRxxS04myT9hUTXbgmqp4n7QhRk2Y
U5dl4m7J87MHCgl5dmIQ3gBYvjjHHzg2rmEw6WI9rO3A7ZdXJaJqK9M+E+r7
C4YlrkLyOI8Z27UJkaMcfqyB8W9cY++RtePofVTZkK/JiR91CJkaVzfKaCKV
0UqN1IOD7s/8tFSzkVLPjDLAH6aIPEewlLe7OD1m6j8RdMyzFJK+/BQHOB75
3L9YV8P+R+dAOzpJDXchog+XcNFhAv0SnGQ2LwgoVXtzmujctjZMB7AN5rLf
f0iwyK+RTtbzKegnV5pJJYYuG1flhD2tP6/l2OKBXVxpXmJ6Ow3uj613Jquv
lbFNgd/7SEZGUad4i1K9cnv1b0kvqm6EwNXVJlCf9eBjOtjuvln2Y3J39nSb
7cMWd6ORTutK7YeZCtvfpfUN5UA9mOSwztKSbtaSmSBljZR5GLUdb8ZDi70r
jXLNVfbWrYWWEagMWyAC9OPNHVab63VAxP2b8iHadLw9q9T0BhxIZtwjcoTi
4I98levBmnwJ7s3bvrxgeWqjpRYeYWEpHiV0o8M4pW2Uk7VPLZR7Oh3hla78
m1s4aLBnoEbr27Cnkjs/71f9J7bnar002qwg9JE1tfwby/voGJMYXQ3+QGo+
XkqhE8GpCF6Ct7p7on+u6c6PX6pFYfaDS6hmQkafWL26IBTVndqX7DQNnCGn
gfGbp54nD3EDzrQtz7xL/d7OJ+2ibqTS8P2Fayav8mnvAYMb/dXpL46KQwmm
7BVYgAS6Hc/mHCkijbjogossTYWGaZM+EWBgkSb5VnVXMhgNCTAWI+bQd3My
N3o09g5kYc21P7rwmIG9dX6peSpKEyjcT+h9XB+QxE3gbnx+ts+Z2gzV3WZe
gsD2KCAxVgKUI6BRaizbK0bwmWGYtY3GAUgmXPy+l11N5IAc6LJHPipMZR/I
ZfjdYHIAIKwGdsgYAh4czI2VrmdhL/dirBhdNhnS24PwTkAWye9evTY9P3NF
0JtLYjZZ5qMzUo5G9IkyBzd/PHuKTTxa7onEuem0eFCvgdhLrN6WEJdl16ph
1AucWv+xLlBJwRv7IS7pSC78XcJ4cieA4tg5LTSjZD0VS44QyFgfcD9nOAhl
eOhAfcKUU7I/Kl/3hQ30iVzWcjKNt7LU+iUaAuC/wctWFuOmFex4AVjul0sV
NHWaCv5fKGCftK6CSU74frAXEF+7Xyk1jMmIFPZhgekhzRss5FjoOcFgW6ZR
fMSjlP6kvm4hY002Ao1aHZWZm0p1nCQjZSNESCcNcQ7sr35EHHvLXeTgtPwf
3mO2ph5GMbjMAajAR+neFadpqsVOBGUXHLudFQ4UPMNKTebqno2wCWksVGkO
YKInnJP8aKutoeINjvLbMRvKlOLugYHj0Pra0ukiR+ilnosvf/JT6Zb2NAWx
J5XGs1rIcw6KGlCR+X7N7xXioKM6q1K7fK94g6EKoMBHJb1TPdEOyfrxPj0L
+4mJM8fw/0n+7TrQE8IN+0E+T35BRcRDigPbhhoKiJQ3yTbNTVkr1ZQ8PrmO
0g/R0DBTFaD0JMQqUQMNTEAIpG4iZ3N1L9qDilB++4ubFistIbOLrhYfkUrN
/0blN1az/1xoh4YKIvadnMckbbLm9/fOyJqOLfMwKY/E0EMgol7XU93IQaC+
eIwBDe/9QrBylOleXJTlSUfxpFMPERSrmZS+djcpxd25lcWltXAags9f4S32
bldIKyaJNxcYOeVd1Ag6EDYO5DN2rTUuDPVliFMKGiqm554KFr/MjKyp/VbA
FzKQgsF9l8ag4bcr2i1dR7RQUOwHtJUb31/FDXUX5iyMGBmTFYI0nC623B16
RNUXXzeuPDrmR6Pf08/uyj+P7jTEk3wT3SCYw6e2hL3D2Za6hxVtNuKx5eit
XURb04uOQM9f6bZMpc8zNg1z1DhRK29LNfNiP1hf+ZIZuCqvWRWxEXmHjubn
8R0iOKpGsMBaMU1iGMpPW8WpHM2w32TFjNoE5XBmGFACyGjIYBy84M4FVzN7
5WpbzsR0vnTzVe1Dbgqz3NKLFmjUcWU5+qTdckJNXnVUQiHw4uG2FGMTg0xX
pMUEpZGSzfoe9a2nMaM8stA9BgHDdtJwdVZZw10NND7SC17+5qDlvgogKNBu
jGWwMG2tUlRhB0SnMoVHYs/TqjMaxLdGSADmnxZDPhhpKchCTrkt6z5LBxj0
iRyMGj4EqXHx4PGOl/W6lbQOb40Lhg1AKRWW4pkuryLobAUVIQ5WqPEi8+Le
VjCdgmVe1g8xitcIYISzq76tpFJBZ99eUud6FK/ZcsFeTa/tJBfNBWOmY/z/
i8hkS2S5ouyZjPfrCX4HMp1BN2SjtQy4yj+bw49o4ZLeln+0bOX2+UIPoYz/
ql7zD4ZkX2Y0+YzqGiOH10y8+uQBPZ+O78zH8iDRAIQoPMxIizYKJYEjncms
amBep/VxD8WyN6I+reh2xHvFWY8qbCdmCqTCkcdXs9F0Dw/A+wIF4xGCyNVH
l5dfiiTtHqYRTTUSC5lZbcyDdmQ/ShIb5YDpzjPKrUEIOsfN8cJv2YZWbECK
jV2Y/3W635pT3MWvufpTYI7l+mn7d6mU1EDdHwlFEv8G3qw81Sh8HsJqnIah
Es4Y6YE1idLFsu/GabD+HkzOBC/RvTGrWKZfz6AboQGs49K9iV6DEkG/lQC8
Tfvqt9U56gcfEtriRdHLwBH6vDJdwkLI8/gGA468pfSQn82H2FKB9KG31gCb
90SVVRehUMenONRxYLOVtbVoVWh1g1RyG/c5r2J8UpS8nJkAO1cCfn/0I7DK
oLr+Po4l6CdBiv6XniACGQKimP6TonupzcCMSvSqpbvKxadXJ2MFDf5Fzon7
u4GrZASjH+5JutLLBVSot+kECwOL09W3zsDqcY2X0yuLcukw6migSo/R+4UA
UFjntEdu+2UJtiwAY0hu8fePFHABVmwC5MhTPKgmjRdwdcep67qf+nxiN6Ox
o/knU5aeNnxt/7BaVD9yuAzIcFGl4pju0ILOjJA9Aule7l2HTutwXZ12bYMj
MhHniDyAarX3jDqnjbSbSQ1wRdE9Om09c6kvMNzQHxC3SI5y0UoZ+goBTa4v
kBBPpmtnaZNN15dY8ov8wfA7kpadprndte7Bf1O5BTVf/Wnda/pERfR/5jS0
Y9SGhhuAc4/eudVM6IC5UatVL6bnEN03oHVa/SopPUR/8qrnfHo4UINZK7WT
2XSHgESKRkYWnJLoUJcphbrg3lFGUw4lBp/k39r3QgCxFh3ibmnylaxxoAgq
aHZjyMJXtdzsgtIoJPrgse+BbUaehZ9TjaA2JLxQcwSE2yssNvcS0lo0gcg2
wtduR+5PZ/64ytOW5aqyj2DU70MbeZHzqRAtQB2PZeosgIBOZ0B2zbRtmkRc
F/i5u5bDQnMeKrYtJhLVqL+C3KDCMZZ7g1Ie7ydukQhfSBvWngMRLsFM7e8N
LvJeFrg3UQKqchkEge1fF0iZhFsE5We/8azm9RVNS/655nt8txiJdSTZ++x4
lHk+G7y9tgqqYn4TYxvYLhKZqRaAffzKYP4SsZOOviNNiBksqIJIdCSY0LZm
6VIQHxOuRiURK8pYWk/ufdi148YYc1VWXqSulMCNcW8h7CR0a7NhPOOz+Psc
6i0Ty55kKfyi1UiLaY30j7wEWpLcmnCUmv7q1uzWUBy7vDf2IShW0wrr5Vsg
D4w+GFEE0UzO5SO4yX3w7oxlHeEIZ659dq8p+D99NlDbsIuSvi7GY7pczWMc
kK52ETT8lovcy8ARmqXRuj//ZDj6SW8TrCBagav6nHp/f3GWHb5yhmdSm0QB
i+e3eO8lczbnkyexgmYuLbrq/lm1Xyq02RWkntTlFtiPyE4xBSdupMAa2ge+
qcSDlkEjYpQpKLjNHrzMwZXLWGtvOpTrXULfYcrv5ymiKRHU+EHjxYPg7afJ
WER7QfsVh57qTR7pDl0zVBL5/qkHl1ByaqsV2S+jPeLfxrb3DqnCBXcMO8ZU
Kup+jOhhMHYnSAiLDqElLVBEeRGkXxmfBYVrONTz4oefYvNtxOxnA4QqJRVk
xEOQwxrwbhS1r+m+svTsqoUNBRWe2H+H+b5iwkICUGWVEZV8En7CzeB/MQYg
KobqOfbj9rdatzNfyl7bjdxFufvbXFTyniKvThE2QVYGG8HmGR2SldI3jqUx
4830gesNK0wq6xFkmSWY4vORBtVmCO08xomDGZSmOlc++wIWb7iOBvGRb29/
2FYUl68uHd0JSDEuVkjrT+LDecoYfYGYgQ1x9pDG4BJPCUHUnaKwh7J6KOwb
lplHgdymvd1mLWDZ7bwhK4sieSjp/TwaOoXCzCO/agY9pcU08nQHPFM/SuUp
1aSJCe/Im4k/eDEcghwCsnoHqza+bkrC+7AKGy0WyfphPePKVdxaDB5gRbn2
RWAPylJ6g/Cl+CAEiCiJtmgLp+cm9VPHtHsiQRNVyhyPzNLguepiZm3BIrWf
OPcK2HhZoMN8LvCUddn4Lj1DXgvX2k+iaRgAoHLEZbFt5vN9dVE+uFiiY84Y
6dE0ow/sY/rlpqy6ZLfy5wCmbtXmKAjSpI8hSY1U659zawo3/VEr+qtFPsvg
Y5eNW5KSRqh5I+DvfsrYZBpiRzSZYvREQv23My9pVnVrZs6RiiQ+GrtA5Zjl
Y6WXUm8nXefMtmZwpvylU8SIxkh3/TSDsujsPnxTgPeaO987qRjThO5Q1VmC
lmx0B1/BWKKib9r57hmwrnJnChWLPcSmTvFtBjH3i7Ghs+kbmD4vY68juSWG
5uxfP4rmVv3rhtpSxonJfB04R9TxAbcyrC/lj9yWE3wW67X7KYGQrZtcUMaW
F9q9DEJ13bQAsUFfjIFz4qN6lv3S09MOvCVoNFVkUk+DlGyg1E9rg79EF9Ob
ollun32sFFvLx719dVxncxiwTUAGMibWs55x6uAiBr0EBW03MJPwL8yWxOe9
URpd5xljwzceI6QNtel/QXbrlLSNgEW+8LPSE7lsbMi0TkgxDwaZRUpZ7tBW
WLZyAW8TJFCUW7hhH66XnPCABOhNjbjywNZvBftGMV316K8rGWvIB0n2AsN9
hu3fPj2/4KN3GZG5p+Z33Z581DfjlS0j3MugzmBMW0TN+Bm9SPrCVanhBzw/
XZpJv+tpm7lNNz7Im5Q7UUZ8AZApeihjnKE6m4haoOgCNPKXEFfoG2D0nCbX
ykBZeGIHgjBz+URnxfKkIJ23SD+3jkHcT702jjqB2dgoUGLpt1dqj1PAGXwQ
/LR3sNOlB3HhCPcAWJ4GAzHR7lqzqg7BgWe/zp9fjm14isfnAlqbBxXEv+aq
r/vVXXtwGBVdZRTbkvus4zHZFwY5BxEuE+BMOzmeAHF5AFY0wKhNxwOOwZ07
nDUS7XOXKyCXJ3G82RvxnAbNXcGDw0J6N+qFFqBKWJhuJlHnWTO6A52IeeFE
xMJUz9DYcMs6K7w6Sajn7OKZlwBPGv6VJn9xoL0YEN9tgF3IK5Ojw8ZR7UxK
kCEUupfINpksejNZ+h8PJyB4/6hUa6JHEP/Pr757u4s5oFIBjKfOIXjlIMjo
t8VCf3YGIvg4kSheSEXnrubcTSEq5tFQrv0waDjvqXCbcluPYffOZPXmF/SS
tqkzz5EG0r7Hvmtw7EBOqcIXcaoSa6fLcwQYQXL/lkHN4hkLRbn2mOrYI775
TkwDGI0oTT/cCu0+KrLV7hKYWn8XiOK+J1aoOqhtaZrG1motGP+q2Bztjc/L
xw7HzUWBz2G8NODNqwvvgnkuXNY33CTIwcYft2At0HUFhdzj9ENEXAjRPGgo
K2VCWK1qGBQKkPnyuZFwu7lyTkjwrs1lTKn4zF0HQHJPwijrv7JUnMMshhUf
6v0lSSfY7nayvzXHpKe1lv9mzJqmSLGeC5h5mjKVbthCH7RUa323FirUpCwl
/3THvFvlGGay9nk2HKSigH+j0j+oal4l0rZPwpNu3YIrE2x/hD+DCl6Uhvrx
ywnvu5byKaHpbospCqE9l1Tcfiq6APJpyw6F5O2t/0AWPtmdGMheHq69JM6u
TUogEdcJrdurR3GUeswVpKdpQbJixfiCD3LsvmiQ0awbxZ9fCXd4xvy2O+Fu
94rGw/ZiCTrulVgkP6CdAmxWFQoEp7ilSS+i5z1MToEyI4x6KYA9L8g9amF2
uQtGt1+x9sGpMXntF5KC68yx/PkL4XcUxOdExJDAhKtzzl8b4TXpRJk2YfVW
lH5Dzm06Yf0Y5aOrWNhbXpXdY9l5oW2sDwsL8UAVxrf7EE0sP62DxXQ6RAnG
OGnOsg/jJUdiBmamLpvTA9VG3Xo3XpT5eop/8ZTPWS3zcrm8HxIhG3XdGMke
aREISOVcBjTKV6pZ+NPcse427Cnh9v4lJeAOHJ2E++ppvQG0JDR36hVw+wKp
q0jPPYsSK7faXUEJXlANjC8wQZ02ZFfN7a6BoRTyGUxU2BW/fxSZCh2fWIUR
v6myYVFfTvfmvtM+ZHx/5drFRN+l8XHpF3yis5wOOyuT58+b1didExiYn1Ug
5Fnc7KVlXCqqHEPZ+WSLBx9wLejscryFCcMSBFZ0v1vhdJGHmRUQn+hUOgls
5I8K2clZ9SXJXI9WYcfdR9lbeJD5v8UxtkO4QSDdrTrQdgDkIddfHnVKEeFj
USpDYAHjZ1BV/Zyf0IdKqhAGYpLjzKAcJm65Eby8L0/jMd0cYnYwC0x+3Uj8
KckiY5t2At08wlOIRWbvvRt22mBLFNWM10+5MA+gFNDbbfKlpmry4d6oLlYH
q/+82Rm8uNqiWLDWXg/0K7FUJSa54xeNLv7vQ8/JyycfT0iP3kmgyeldmcvS
soVlyTjs1rgpEMlPhz/8VRgXkgsfysjbg8/rNcJ3uomQxRb6eBOBMQ5U+Dz6
482xyC514vMXXOukAcRS5WFJz0PY+OzYP/+n/Aah0CR1DOwyWqrwdUH7C0dM
e22uhjhJmx+etD34j8BGSRT9iWX8/0Yz5ip9frZAiE55H0aZmMJDP9YfXeWD
jdoBVvL29f04IyK4aGVPmHdhM429Kxa1BDdR2uzLI47XydiqGnYcK4XfYeRZ
d/mH5zp0e1Teq32a2dvaCPJQSSuzWLPP3mo3tH91yO9nmbJSQSsDVskAH0Kq
0D+vYZb9a0Kwk/x1FoRwFsvVhG2qFoxVttyHIYaejqjvh9BFyHzaUfl17nI+
hcDOZauL5JSRYlkpOrmKjT7aNlc8AAD8lF/67+5oYcwpL/y9OmK2hYhJh5PF
W2YT6+6SWWS2IGgXqQcHXZKPY2wUC7UQWRPtsGS0ybyHGVJlXPOglZ3XQE4h
O2VWpBWf1mmWSCKpsVHbM5cvq6W1PTzLItDmqIbMShb5/trhLkK4DNcDt/g/
wlS6eIaoyz53aEs9Do/r0O6JV8rQwvIdSbzrTww1AG/iqP7tU8BmRPECJzOG
Gi+IVuRCkzHt8Mm+jIAwsfrOfeh4xOOu9ur40HrPcE39vlTYp1kcFHuIyS/C
f04csckh4GCErzwaIXaBwl9ScmVlgL8NnKpjvQ73mbCbXFti/nFBtu3Hl7D9
tDH5F2gCJAagqbzj0axBjafrGBr70C53DsuDrUvx3PmBBbgdhVXt34Bi1NSy
noL1GH3RSgMCyJoS8FVrg/WSbIXsvkYC4dNLxOj5HnlJNoXcDaVplWM4G/qT
Y7ePPkDUER0L7Ef5oRp8ZSjiyuFANf4P+ENilqBVw+TKOpXQjYanW3Mct4g1
Ybpt2nu9HO6ylvVF2s58RgTdXAy9OnU6cOyW/4Dj62HGu7WSgJS9c9hhU+D+
AiyUxbWZAw6EUe7GJkgNPWZmvzwkMKr9+Gxnkyg6BB94gnh6pL42G0Zkgf8t
D2v0YCag5aP79rZqQ2+ZR+whDoYn25weHsyfFBrcAbQTq8kXkLm1C5MSwlVL
099g3P7dUPRcY5+O3V0bbb22SHHZL3UFwJYJsI6mc1BwLDnGJ70ZlG2R+oze
ZJGM+xvbiwiQb6G0ezmo0yOq7hs9u3ISBDCa46UTaLUqAYV3KhCFBkcZtgA7
DMznCMQEsKGQhAHX/rL0800oisADQCEi6tG7qlG37rTIvmjskorx8R1iJZfm
LZ1yGr98xSWbFPMlnriN+CkbzyoJD0Qwoss8N8/O26fEqOU0CzBQq4RdpBc/
RhbTM4bJExbKu/Uxt3qhz5dMyhAnBKzPUcrNQzLZ1YwnUeG59hQMCCArRoxh
6B18PgPyo0Wb6+ALLUfXUX27mT7CuKFzZh4IRRllPJrogJke/V0RvaLRYpEn
JG0CnUi3dH/bBwEh2mNZOCte0UiDS22ebKiFr9nSKBMeqdmjPkJQVU798iab
wx/29U8ALUOs/5Ok6jAXBb/hbgSnpIiJQNHMRLJEFl+ZKwvttJdAZ7N86TlE
tTFzYKvZs1cSPyHWhE9vTLhsVIey4OJgVwuR1VZi0YMup9qOqPC34yv5rgdG
lK1X9ToK/VqMCrfq5HaRlnaDcktMlMMcZPHAE/wjmDcFlQv0WAOtauDl+d0z
UunNz2eSKRLpecnoqx8dmPh0q7EgaPcPzWfZ1ARG0NFgHfYKxmmnxKEuCGf/
dNUKqGvyWI7FYfvFXaWMbeiIID5DQAPLisvZXFF6YOv+O6WINGbi1F0QhGaf
tBAgli/AANrH4I+4GwWQcrjknJr7sk75jBLe158rBlFEOtqrYf4pXK2InzFC
wIPeQ1RESsbGLwaBjtDDPRg9x6W0Y2Qc9TYXHOSfonho6p9S3wuiyE4SIJu7
dqy85RapSEkkTOVWl28KGxymbjSAKviWlLjdfSENrmcV1pD9PfLONy5MVHNG
4N5QVd0+HRwmQftZK/H81/C1oFDVPKUY0fbYgE5Oi+v9+ORVoTYRy0q1Vi1V
o6TLi1Rw+ya904hgCdXx66KlLFDxr5dP3tI+V7C/JqRdF3GABW+ZC0QcLa4h
v8V2IxIaOgFzevT7sEEyYRcc/afxZtTQONYhvWr9tlktV/sn5QHuzneSjMa8
MejHY0kjpeIoQ8Cpsxf1OGXOIBEr2u4FOlhXarZJ1urI0ZR1GPKdds0ON+OZ
z2N74nsFN6KOTEE8GSMyK9En/OcADUvgbiQzRM7N+XNSwL8woEBIHUhc/sPb
dCAh4QzBhnpjITXNEnvJVP7Fq2Ns+LX9H6btmsSIFJkDLrw7bhJC1UwtNzcH
W31lNDQaUY/Au6nStyB3So+a13ejJyQha+SmQi6mBV84mGBif72gNrlBT5fb
8EnKD8M5BC8YasxF96TCMgkjy3uMaKhTZuH88YB3M137IZoAQHmnGixz2iII
LF9hWrK9GMUXAwh6aityw2Th4YbtPmvBZHZTlK0sdXskVQg6wj0gAgVFH1b3
jP9YpTApR6N5BheA4MjPoh32cQqYAKlY3+nU+gyVyO+ARJfIt/npFwF7pq1v
h45y5W9gUVdUL5m6QsmBBnhUpr+oZCzrQtCqAfrh+IS17Cf4yPSeid5pETdb
gMXCViDvOg5BIP1UIVI9MTSnNWfF9dvmgjuK7gduAgH84m4sJK00wo6eVCK/
pynzdP0q5r6R7BKUcm0CtfdI54b/gEToCfOji4ulG+N1TkwVcHadHEMzI9yC
BcdWI152aYX+SiY2a+DlXQxdMkbSEfEqDaKQSwmb7gko5DduY1gL2nGV9MBX
zOpI2OijWcESSaREJR6ZSwnHJWxl0KG0s37yuzIQTeiARCMnSjxvVzTfkE77
lSKCMUw09E4RguNTf7nCTWd6lkpz78UNAlSD+wuSfbinmHq3OR+tSsrabGv3
ENmbwm1askaIl1blOxMciMLgmf9+vihvp1FyATw+kJF5bg2DC5/jlbKUVTpm
xdqDeNrQlrJvhuxH2gqw0e4/NZXRsNz1nQluew2rSGmgcJ7a4LJlF/NPXbFa
XDgejGOEFWokt1NTk6MV4vUYlpeLIjU64sDH3PN7hJgZ/zv7CnhOKPeqQEfv
IkTPBXIOZ/7KgyiVI8La2YkRhBvdjLrSb2AtsEA4TLvcONbFGS4uKHSzk1zO
zlf/vNtstIL/4GUIBMv3GNQsGsDi4IV75TRlZ0NjxWZUrj1bgAcoPuOlTcOA
+Z9zLBAcE6t+eLmDVicE0SULkWDjgu5LbHEFSnG54KwM3fIOD1lhO/DQcXaU
f0zcD6Hz3KfG7wQfx96MXYvxGKyg2jJx5Ccn1xfweyfs1ztWwYJymk/HlDJh
4t93P/aoMaO71alLI5M2fl/s38vhSZImJj35P0ht9Z0EDbBZuwo0uaiC7vS+
1I/RghPdxysZnATp09tHZuB6onebMpKe1S/l4n7uoNvTwCqi99E8QcVuTFTE
+5/6RTElLQiUhamqABvvnluakZgdJxQ30bQOA40LGeuhaDX8hhHt0k4erNm3
SJDlXHzy1Gin+KS9ADbaYu+wY1S56/xaJHD52STXNFYtuQdVY3YkiUjG6cDY
O/o1LX9c5Avso4mZMpuedH/4iOAaWJZbZRBsf8Zau8B8+rO0Us8FDXID7iPj
S5LmJRFG991hBTz40QWX07o5Tmbt3hjLIB4CQtUz8Do3lQtWjaCNPGqTS3gv
/68WofMZ3q4W2UqBChccG4g89/GCvux1wC7lcVhB0Rgs6zfnFSXshDf76Kyr
UDm/eDi/vTUcolqRW5AheJ7OweRM6GODTIYNc2FJOoSqXAOLGGVwy4qgIR5y
msY8hGH8T29BM37Vbllxghc3xT9NOf8x+Wx4sCYrLXp5SmVin2TNvCM88C27
Byqd3fbmSDSEm9PJUjq9gb9iKdUshrHSe/9FAcPVnAsltAhxi/Nrfd2usHf7
34Hnyj+TpgI+HbBrjyOqywEP4g8CuVQaWj7hN4nzG4bBm8jlqDEWbtA98WjO
+4w6I+gGxVykrLrKsLjBOcxL5EoWW7f4bEbp0BAZv5PbJDOuBF3Q2jwCsGyj
/r6RQD7H94lQ+YyxRP67cKA0pp7/3NGVGgdtANJR6eMeKiPth7OguFafEeMV
+9/92WQODNIgwn6MbPOfeMcYXPEBRnj/7Dlsmi5pq5vgTDSNBKI31gJBSFgN
vdgfdDmikd999uatBpM/7b/IixcqCmNlUtEURi7l3gLwEZpqogg8mRarjFml
4jTJonoToGlXzVU9adJPBZ2RGsRYkwP7mB5StaBMP37E5adoqBTXnFNJA7sF
bU4Xv66efl2ctXpINcmCsYrR1pWZNJdZrQa3W+tlghjun6Taa5bqG5D5jTv6
fMjIp/fLUbbIB3owThP1ImECCLfGBN74JHXm/HBxNWslV+qwZ2Ypa50PDUHY
COlY9OOqIgIgLOtVulIZS3VRSfJgcZJp0c1+eUdgygPlY/OrO15NlH4v5ZZS
u+/k43F7hNCAb6WoyeJYt23l62VN2By7+/0B7Ir2copPbXXAxPM8cgws0qh7
AxawM1yTNasH8u7m0Xml20hkG8dU2DQqUfaAG2EFESWqdIo3fRYmu35sdOtv
qtRhI9Wd2mJ0tMs9cYtVuqSRezsTAto4zSqvYA0rLQvbYSMnahhXAivV0CBW
yMIhx5RXWG8Fy8ozob8zwi/XPryUyRp/VtZ1bqdXR+qOtG39sIGSTHIjrjCc
imCTPOt07rcmEuYKN5nyfTzh7yZcUB/cqfyBqlCy8ieoeFoWt0pj4vEGdWC6
wMKpQBAfNAQzNf5oZQfIggtP3LvVJTim17QoLqmsNGQLN4XmHGCPk2oNWo8C
hMWIscTysLsxx+Jvvv6Xjmj0Vhdyp8VRVNRqaYKxQEh2dCmc3qGZdVXe5Kju
rQsAE4KNgi+ZTfAl1zRtmERnWdt1RVsxT/jBUuT8Q95UWr+1XHNvoCi/cQE/
wXpHN45+fNU3ahTNTGbOhEMTDxk8nQbxzOoZIB0pMF38gzyZm3j2Km7pOC8G
q0bOMHypI2urgHohR9DS/M6CsdyG2H0jaxLnkpOlv69QenQ1hkut9MCrNXVX
spZQ9lKpe7uRCBUSHbmXJrvtbs7ptnFrq4dAqsmMMCpviRAYlmN6IeHUJSqy
Ixsy91lbAe6PPRx26rUA0Gn3JkAKXpzIrOb0wTkXe83uqOcAaUcE6FzYHJ2y
AbmWecdLqEVf6GTXaNl96vUUUbBmCXr6pCaQu3K6dT3dWUgjzGa93y04xm3q
+KG2jDPGXnBR6JWiBFy1bRIL81THWrhV3wNtT5AOqn4vFVcykJR66YhLFYNM
Xc+cX71HEbJ9V92Q4kAqHMaVy4W6dG7gOkgdVqQceBt7l18uqBtXXeoP63OI
vcQoNXxU48HEMsK7l80QEhO3wHaE/fMHFBU9OO0rGcnRNnfVT7+12S5FdwpA
7YA766P0KT4EOTF1omLm8PCY0XbcCa8ZXHd0q3tEHuv/0a63+5eZEj80pnd+
pCIgT7G+ZvuciZ3tsSybN3cQy0Caup8l+Re/UN5RWc3QvZyEA+RF1n1pJmgH
Ppr+9e39pCzQ2wBbDzeCfNfFWFZHRDK0q+pensJQNBo/EGMkgylxqxyjB7rm
0gERYX2zI/h58POGZX7xZDfyAAgqKtfhA/2TiXlQGzWdMJPg9S/QIxxag4m0
58L+eh+rH+SWFk1sqvUShJqJ84/L7FL4W1HFz5hJOYK7tXDiQSfg2zTuTjjm
UBuzbW7rjJjRt3/WzcfrHQih0TdQzurnhX12pOJQpgEGoqTdJ4UP9vx/DMuW
t0VSX5DUgkj0KaYJUiri8Pwzxto4KINLZMCIzqX1bLSuPH78RXbRIBKkPwEg
XwmPfzLWCm02kyGgxI3s4rNgcHFpwtTObwt5ci+QXaFpkdroPzTS7kAPNvNn
bekVZwe65j3iFGkSZpct8c46Pg4VwFF14OwS9zFKxz97e2rXuUyXIpz4hSDU
P9c/5YTkOUX8zt86Nx3D1Fh1YP2qXP+nRZCDhxIkI7tEOxTnjapYipTbCyOS
j5t0B78rMe404ViYCjZ7wEjFBWpkrUHnLZ8QDv1CYg+HuKzLfHbhRg89TRBp
FVjPf6rcSa3u5/5wpD9ZhYqHGNKGSrPC20/4Xr9HDV7yDlPdWQNaxL6xC1/x
j0w37T1zkX37efbA5yB/OROKMVX3VjDwBuo8+TfYSwPXhetdfWUxy2SB+VNF
RdDNLeakmT7iU9VGjYLQ48fHn6YnccGGkxr2xYxvvAZTGOHtHDt7ASOGkpLb
OxO61ibyPsly9iEG4V2AineAg411/eDAlH0VMGYnxPUC7+Pp+eMtfNECofvd
CbUhIBFsiBATWtaSm7LsmEYDAkajS5FVs0TpFuVLIdbmjV+a9E9fOdlyV+of
DBxQmI5r9oMuMvMKfwjhBfiamzKZsYZq5h2Lp564X7j6JQyvBtP6INBcGTf3
rPkgqWI3XWpPeVbfmtkr40HX67SAV34L9oTuDTV7wCEmDP54d9+xtyA6TsNy
T31ekHoWuKfJHFkhKsXOQ2d2AzH3JWj2adSMH+uLaALbqMiWy4i7n1Pr7Djh
Q7I+Acry9ng3yJZU0/Fu0UC15At7zrE55uQoe07/3G6F8vdoxdEgxyF/evyL
P5tYYtQ2eLxpo3P5cj0VQRApLXByOer5HpeVo9HIsIjsiiL9+P8RZSeLPAaR
Cdnp1rpKRaas0DQX2bhSO6rXKoYu6cif9cVn37wpPJ2eXR5GV2ZlBxmA8PzD
4aZHjZM0unYZ9Hoyy5+Ff1OEisZ5VWkvyYy+OwCGRPIXbocGLg/hADYSClPb
p0nvh8LG42rnj5Ehgnj95mogFM1yf9u0PJb3QFF03gQiofAuIeEqqAC/Xazv
AL8Wx6JHrrgaDudt9aMgAVIUsbNBQPUZCQZengwySEXk/5ImJQUaa7pwbfU6
oLI+XudmH6oY3eu5U359F7E26fPF0/b2iS0FcxbhOqXf4vO/scZ9tAMdoTgS
0E05qSjzLijDvayaQaVPRYQTiQLAJb9DY/Ogyj5lMI0GvcAPMJr/q6hkdsBs
xHKugtNMMyB57oBJ29Mi1FWiCqkfIM+lkDfSfAmjuF1BZmHVw9di1plyrlov
AKmy5SEOxgre8JkJxkmNAXF0xrzpcnEP98xvEzbng8swPU/7c1xxGyp3z8jO
AnihEmiTEyEDtzjIxiSYZ+/S9R1R/8mM7kzjH8H5pvWeiOYY3O1K8vYE9kc7
OpU7X1l82+3itVGwv42sLdd0goXdISfrjoCEyLwm5ft5GMbr/BW5yRpGW1If
RWs5Tizy6tM8bzYx8NdiAbFswP3MVn2mNW2ZQSIOClUw78AZJXcrXkqjKF9W
xVEiU08j5z1W8kc9PUm05VcW4BhhHr6tM8sag0DqETpU8r+CVjWJ+27II1wj
8lOGcJTHcG7V2DvOCv7sNX40Uu83i/3RP68GuhIkRsXkQTgHM4ErRjqLWqdF
WPufsC5da7TQpv3mb7G6sXW3gW12YtavBjEsjcxHiU5kInz639KMC5M8p/DS
LkPdwmzWiufQ7vuK5JVHDtGRjr2RvJXUXK5wAe+pt7DI1RsJJ7sWbGrinh/I
UKA5/4ZXu27Pepsc4DDbSWnm/v4R/TW1RKkM23pNuTOmcAEIzfT0jELEQZ6F
EBX93/woN6l8YW5nPDX4nZjQHixLNe0fgPfZxFmpnkHX/TzENPGjtuJaKZ9E
GSXfEkh7VVc3pV07CAy2+0jB5dusEL2oD82mbBUXfnxKfhcO+vxvryiZla0F
UcL3ClN+eyxg9PDTwVpT1fDXPI2EfJacX+7qnmZSHUhyUV+iduDghCWqfB6z
Vh/MYmDfmIuykGA5snhZTayJ8XRQp9Up+7Hjsl4pVFbg306mnIlXfX8CZE6f
Pj0omVhrjyDwsMvtbLejXO3RdXL/Sd/cDOeZz8i0omgvCAPnIBUxD0W9uGGG
x882u/NQ83/erIJZIlSqNeDwvtwIAGdci8S5hO8jeqzddoSpiSvOkzFspMog
B18/lM38cCMyvKLbtTCvCHspxTlVuMOo4HM5Vmd9DTYdU88Nb/4AemrWCpmO
vlLdb+34H2mePsCLXYVfvFM+HOTMVk+xRJbKaMLCcBWrcwBe9ozLbsO+m8bp
6avDSog1HFjsVZur5nihjdddO3fXhmgL6dYzkgs+98Qgib0YTO+FYbCaj0O9
Jfd0wpnlOv9nDw0LpeTFfFZSuPD5+niSJ4/vJuddeXTkHxkqPZQGqZ1Et6xL
D0wS4MFv3fsn55M22KUdMwuF7bUIhQW7G9gQcQ9BCOryZ7cPksb9/FSv4tAr
6RnwFhfvJWFDKCQ9/9hXsDp5PhPyzpBLOA0yySLC+TAZLzwmVPJo8jRWAX+l
8YYQ73NvJteaWG5sJkuqK9/UHz0Rb65OiysYHkZVjB8dueBirSLR1EGodkGh
bKLwNO/INlId7ro62w4J3f/Ifqp29ABiNDjXPwLVUD6vzPLVnfgjPmmp5+CS
z+lp5QHYwXpNQ1F9AqOrAIrI+0HMts5z4DQDYQ6rRRK9/gDGvCRiOdT4TGSv
kAtkHtiLHMsmKkG+JXHIILyOUJCMJSajQgnLhHoy71DVj+5F5OGjklzqmCUK
7AytZaqpqkquYkN7Kx/YwBDlnF6AogXRQ4yJ97FMrxIoXW9oROzf23L2gQ71
yn5qaRYV1kkdHuqrqb+wvuq3gCH7dTJ+wEsGQOXaFJTfn7+qoQxb61ZEiU4d
Bu6oq2fB7nNnkLVdwBHAf1PkEsX7j+4mDD3MqsqpYXRLa1s5jKVLdlO/Bxrh
8LJm/LJB3psd5ouZ0aUMGfIsQsdOSntOl6GQLe8x+NkRuCRTlT12gYkNPN5Y
OiUQmrL8/fFSFFXGAoMrXnmqPLhtDZgXXz+kYb/5dJzpeJZkOJgBQjfOPzAS
WbYb+4tdILwN7042uxFa9YqqxsTwHierbuipVtrsmRdlJPiPJaaPMM93lCyX
X8qeiwsSqJAcgI4KU+6fFykSgMvWO59ozYInuxLxxkrql0Dl/FvyLlK5zYqJ
qKgnxxx9DG7E5ut5dBe/f2A/V19tD2fpEssbk2LHj/LxBIp8FrY9oBOf50YS
mzbzyt8Va/jqdSYm0GvABPRYwUKWJ/vfcebiR84Re4+ceg3v4cbv1tVS7aOl
3crYlP8UYVB2DLprJDAzeotL0C3nmlYc5tdGEoNpbvFQ+J5GVmCeBxGTiYmM
9lL5HkvST+FdybiZmXr1hb4gl+11dizUCVBAsPRwKWb/GgcSzGf6BRlC4CRm
WbbTgoZ1gUqkfv8Z1K0v72Lwo+l5k9GTLaldc0C4w5Q3nKfyNNlMyHn/v2OF
H1j65xUhJC0cWs5yUBK4OOTYeBY+3GBA18CktYc/sKqiKPx2JfTfNJEq6pu8
E/IzqqX1XE1sxKqKJMInK52UtNSP5+I2NMC9a9LIboeH7GfZIfjoLxNsMAY8
0lEZcXrBdC9MAI2sWuwYMHO/Lr1uB9XoZtxTbeyHHW3eVFhY4d8y1MkWYZ/A
nh9Iz4QlAcRPzylRYKITZDHUlsD3ruOmBxE2K+jO5nkOC4QCi7pZmiqueW4P
f7frlO+59qA8AbEZB86wK35c6oVJOqmTK5xP8kd6E2pP6rfqX/l16lT6DvR5
ZH1l7Mo2359VTwhBaIuw46LniRSAAa2XR9Cc5qeC1V7j8IWxU3t8nvkySD73
6HDSsh7FofNe2KZxthPxdTcxI/Pv8FQnGKJhDhWbgW/9qgi8XHJyatVTJgpC
pr6ScbolKihLPPyBWKzzmJG2/kJ7pzk3NcOlKcIvQnsPrrvojQ15rL2qCFd6
4JPjV9h13elD1dZ06IpsNimFhhWPxLuvwXEKGoHKRSd5bRkgdzKqaL0QLPMm
EYj4q0d7fn1hKuh/BKl4QUQ24QWGtuuuD7m+LkvkvZOKNgfQvafZFD3vUtQY
L3nUhLjjqt/B0oJCC2U8JrBXMWYv+r+9/PxuD5zcVwt2pAWO+WBWNMiMn9jA
E9cMRQ+zDe+BZhuJYrCSoEKRiY/IHARJFaI/mWq6kt4X8pwn75TvXcWzuNug
VrliAVzFr2RtleMfGYee5BvHpz/KCG/5Nicj3zG5gN6uy1C+c7XCojGKhwLd
aIP5eJvJb9Gi/pBmFaXToF6biOtTg/hIaMFZS7pe6+grrkN/kEMyKW43sXBo
AA+Q1k5yVcG+UaK0Aq4z1Ma4DbtQypkXwY2N79z6qAK4n2Pojbi9EdTA8DBe
j85zzXQaZpJivWnG/3JAgheBl2hynw2i0Dz4jxIMn4zZFVNh6ngrN+3QwFi6
9iKe7c1+qGwAzAcRloNsUaEjcn9+J+9rwBNM52wE4Vofk7QIhqitEwtDh7jh
uSZF8yIs6/DH4iQluCQjyK/jk8zSf/ul9lPpL+qU6Tu9wNF5ZMxx1g45Us8X
ej378RJCnvJD1rpv/wNlOxphJHFgcP8JxmT9NPTnNhPCWBpG8teE2PBAvVL9
fTFT8rU5JxHfyEXk1ftyCg4XolS1Mb6Un8kFBBiU1Dg0BLGCPDLkVawHlU2A
4vt+dXt5dUYyac+jJyX5RiN/URrqj1kCunJATFaqG3p/nWvL8e2fLiMzjxA7
8HA/54683zS/+1Lz1W5iMYknuQuij7nFGRUVSjQc1FNXrkMXALeGMq1DIJL4
TjE67IoGYopetJ08WcJQg5s576oO0QbjrEk8xtsyf7G0YBRl4Lpe70vyZI4w
y8mkYidVtH/r6g9Yt+PZg+Si8ccFeL5797K15CjWZ4fsn89ijVZ70qBr79IJ
dTDpYlqCOTaucjSiYQUs6owiyk7d1z02c4MCovL4RSw9CqXxGTgfhCzSqIA0
jmqfCwNrH9ysktdqWfMUWeWETJV/mpNKwIaLniRverZeqMFAKrMc5UG/8gZa
GKVQdESYE9k2g1RDsajD/hWfJkEYX0lLZ4sDp7PrqebRGTI8ShhSriI8+EU7
Df+KiAmTRoIUjXeW96eUjdK9OXym6sWTo+pNdoNiL7J7Y4CohJF49rDReWtj
UjhjaHvI3ybEtvV8NueLXMWQgZIDX3BD1ijzAtvzxyGsWD7d/7uiopMqFEwY
D8Ys48tHgIZHhbaUhOXKa3aF3A5nOVvnp7hgt8VSLtGAXnYcTRkY7e3mndEn
v2oV8eahfyl6zUYyJ7wliZOwjreU/md1JJoiNsuCFzHvVzmUGVtQG2eNb7WC
rPyUGWLkGwMXmeSUWPGpVcMnOYF06/zzeWnWggGRhaafvtzFRQr61g4tWhRU
DwvuGBSKsFCMHD+IT/xzyTPGMgqw/xPJQcQIZRVjY8wC5inrRTMk1vEHIKMz
1Zzqi5pEE7Cp8tYPlx5qsdiGk3fFQYXW0aIaNY6YN401Ebw3FFp0vPtGbMTB
fZXXm0oKoUgd9eHN8l/T/z4wM++OWuzJvqJncPgSUptmXskqCj3g1UvFwQq/
oXETipPUyxiopV4yrpMULekOFLWEqfjXdEmudXhJQdqfjpznWEdPxooY6OEO
slIH0IN3HRDwH2e47rr17PPTnLdTPyevhNGaG9ZLMiYo8f0MEVTBOGIaUKHm
z9IQyxUO4A5yEpA//i5TnkI08msQKka/V/veeFHa3Evp4XHNSQLnv03sgjkN
OAcavufmJNnpTpD4LBpURBU1aaZVtoTW4EUWP1hooqFCa79xb0B1mt/g7+Kh
LEgdk+NjtOrWd/wSxGr1nyer7S6nyAw+5G3fELrkG3ie5CjWGBfu0DpDe3yM
gGFSlU9XqacsS68n9OIHc/8N4EviGEsmcvUQEyIaUNCCOcl+V9Kzo5hOVxhb
yl/T/2JKmI9X/xxJcUWUh2RF2FJdbdwzO4ZckO+k0VXNUrUMk8bggOcvNFmU
vTpHpv91aNqSKC6zZ4ShW2BkzHLaOfaL7jkM8NQUB1yZPfNv2e791bAFoJ4q
2CQ7/KK4m2tAfyU5b0R8iO2L3u5t0DPUfE7JLI8oP66UyVt7RNUraBYIjCsO
kWns0beKttwo8mjnWvD9SRkBBDL/bJJ108MZmbm0rxKY19FPNklqNcgChHky
l9c6zkSFwnJvDGHA9vWD8gt4HEP5Mw7DxXDcKO7miquQ/ec6irVz03wWfSQv
NAQ96s8ow1M4ALeAqe0uk9CM9f8a7AOMPv/EKIXGI+4Trn6BZVXM8SXA3SlP
EFlla1x/aHkn2Gdl4haZHujmL6E+UUMrL7rj53ebrnhjfGk3+nyz1VX+mM/u
FDUpuSBjMoVpXSbkoe4ZFQD1WkkW48z6zP7jT3my+wSkgw33m7dfHkrYR5DV
nyagc25MY31xlJNcUVrP949o7XJrjdi8HSJYvF3TpKele9N9TqBqzZfZfyDl
1VHTkJtBqGmWJ5vldwla5JixuOqgL9DpSW9kB+yPfBVy6p+TgW9ipDqktkFD
BGlvz97KCwXOFX7kebwaxlqNp8tXlawC2Mq/HKDmb0hM3jhtOGhFsmEzSeLu
P5zFj+EB9++xGtwp8sBFOanvWyxDKbEuTKoKHCQolzmAEKQKvguZ9aOzAux2
XRgmxNUnPrYNWUd+NWlHzfOcq+aAla+8dPNlnI5SusOcPKQeRB01wLwQe6dm
15l4XFJ6KRG0TdrL8aq/rkgPSy67KPYW0Y07xHW2S3VbMXReqLt/Z1CRuUXs
Q7ziiaiQnxjsGYswJm5lApFg4GiitKvhTTCx9lFPtraYnhIlQffGAubOqju+
A5q2zDHNh6sGqGjriYamYuTQkT0r+aigi36sa/OcTZ6CZVgpH/NcOEMfnvzL
tCCJjFetjLCFqKB7SdUtVuS/mLpsIAg4DoxilESUZ96oTh+W9eGP6eWjzB8d
L3mjml947Wbg6FyueLiYVs72VtIVcrmYDHzh+I+bBUhPl/l2Y2Ji8ksK9AD9
zA63H7h6qLYi/8l2nLeDTI7VtIrM9CZ7MQT7VVN7/qlUWB3dP9+LwMOVJOKV
MjFb+2QO185B0as/5p5DFCo8nYv1EnuASb86RAEvZ6cymyXifQ4qXPMdGqTQ
lQu5/1gmD+xknm/C3oM1LIdZZGLilCfPH5T6IJMu9ZIyLORB4G1depXvpJE2
wjcRtaCxTp4mWKX/LEDYaiUMrNjhgTXW8sinyQUMTu8ET5kiuKZNotyMyKEQ
nm/FscAfJZ/u2LIoHhqm3pU+lOn4J/rD47z/JQYpZVleOEW7j7uel3qqyipZ
lmeA38AIev8LsxhbVDC2LsKYltE7s1mXIRMFVuV/hVGaR0xsXnn1m7mRSsUx
WluA56QUUC+BuleJQFvi+6ynM5DbRF+YevbTMOhkbHJGUdea1Rycbd7RrTDU
dV/yfmNxZIbqAU2iHlLAPjKDrUxunkIvaZfnOJAg8RAXPVbpCnZJ6pjMcvTZ
B9SfWH3gSR5kePndRk3oiFl+93hZS7Rj1QsD8/8nJFl25G+u19lR5HBh2+/u
XjZLavVAOFwqlwLM32Un9buO8QUisRPjtLd6YGQ3xdUrKqhMQcf8A2AOFSY/
VQAlKPG2w8B36ci01unnvHWGM4WJcLhjwP60UTH4iyhEHBExJVe1X9RiZ+MY
4qx0v357K2lX7USzKo/gKchYGC/jTfaxCnpqB4wxwnmRJrzlyhrMmIQlP/8+
lksnzBdQpUdqyvYcEx8YgsQkcMBiGyy89OowQdnu11QucnSG65CD5Q2Jd9IW
66qwvSbrEfP96GyccwCquYL9qIjPTi/UOHRrR50OemDcYWJGzEsx/EruoKkF
5VmyCULSfgw5ner6OJpI7FWgjrGT4KVIVhrNffqHQSRThby48gRR1gZX/UbJ
k4EPiQTtWcNDZGEuEAofRFjCjNeSSiT0PdxwApc2nLKpmeRnIAmaG30F/X4G
g04wcrMbQpPh8843QnyzwNI5K+pJvyDTymhRmYfqPRn6mzkCTiljUX4U1PLr
7ziNKtOWK3FMJcWZjE8ImwmudY735Ks3AF1jB1P9fwY/q20nDkvPzOVoK767
YyF1jEMtBOvl+Z7FdPtPEw8voxfBhjhQ/Zhh/Ayc+y1yUCfibRmqqYkVUNTe
sBDbnxWql1fR5umFYPDYoo1RBBoeY+p2Eyz1taJx75s4zR8myF4WgD4rR8KG
WAJnsU7rrkCDIg3/YL5ulx0Y7zHJyVmvMO/+Gcxi2jeOBlQN6byZNtCawhrj
aA7B+AIOYLd9RPVDPv6tb6P27CzP6vkI/TNi7D68fSOyJMpEObdLYMnRJUcg
vsIcUp7m2CuhkEGvDVu2lZXzPc5ZEl8h3x/2Ww6FZ5LNMANtrDXc6onDJ5WX
aPDXFBkr5YVxszdSTmmXRpr3tLuoeD219ZduS3guYfh06OqLUcBNWe06O3dM
lFDT+rHhjn4JKuVpQJPMbHLhGJ+Ih4sdcHEVeiygQDexgmaOxzOsDRnWma0z
ahDGk+ktjQmIZe4w3tAn7uc+n/6Qi+Y62rUDW6XPMpSLdgNYkUr61gJEPbQR
5x+Vi0Fd16rAIrcqgcQs3qdBhGfpRLPxSOCt8ND9YE2EaPQ94X/Bg/wRcT1p
iTIEdBuXfk+a+bv1l89R/Wu3n9JzbbpsYi2kEyjRWBheY7DqpheFZoJuGp4X
Ux6WO+PTOxnkGegzA4Vbk2tLVDnVLgklcRmshlXyUUqGjbyIJpVibevhSOQY
/o1J2ZO3Hms7E1Dlu2cpwsRCwEWXHW+1qOuVoWwToQ94PzAjcvy8bkmXaXXx
QKziNS2Rec/30f2T1JoGv4KHciTMXlet50t0EDGCCz2TlokUqiRioGMpVNfW
n4uNjmSS6uXeNhV8lXZwt0EVOQk1Ro+2Vb70EAXvOnqD5RUT25D7G8qtvKqi
BfI0+3FtsCEneo+tG9V+cCCAHe1x+BzPt2P5bxwAnEIRatqxcADwcLdWveTW
qsuBcV00HrTM1q7GzdXPiiYEMN+vRq+5zmlcnmFKISZRMes3y/hRfH8iWWJG
POggM+mWOusZztwiOakXPyaIEvgE1ik2JuCYRcA5S1A2rotJ0+gGGnH8zbQP
3fnrJHY1MiJW2luE/S5ExokiJ94nbeQ2i8tF0D89ysaYF13W6cG9lG4hLQ1X
uUVVFV03hcHju+Fx9phuiMVGob4rMSVPLT4SVPuD5hgmRUoVZVe9c1n2nxHI
8wwnQ6znlkGB6ILk77cy/LlNMbk713BmJkEJrR+QCw2MnClgHOrLfLtt9e9A
mPaLIEgGdOI6F2Zp62G9qRyVzGvQBwaawuKawCt53JfHEm3QVjsPIIYH2u60
BJhsqTmfpV/gusxcW/cH44y/ktMZQ3ysGogyQH/RnwyZT+wmkPRrSQ9mgkIQ
wzhveoR+J6gnICwvnmW9QGbW42ra2fusFp6Zt5BQC6Y/+8rphCtbIMuilpya
yuw8XpJZM9v5vZPQlG35kwb6IWYUUn9ndVbFHq/cLAvtSuhwXHRzl8kop85K
EK95tdOIfndevVTn8UM2UKUPwkf4GW6kLYzYg5EfkxNucl1lrSmNv28rPW/o
0sF8TLCEzBuaCl0nxQ2LLr3ko1Em8RzG2+4BcVr5g6H6h1CUpCt3o189LGCR
0CmPWKvtWvZV/gQCTKtfEkANYdQ9y80hLFHlZT7RaGz8MorlhQSgeIKwuUrR
Q2jFQsW6VZByFnecE1UkoBSL/1RSHi1NMTdOzqXF873zOISLfpYJu0Vz4Qbd
9l+sY955EUi3OND45scE1TgKRkBB2dPNQaS5YXz70qx7eby+ifpNHDCnG27u
xnKQNmdMNMNarp2F/V5AmEF5wRQJdZfbXyeq9LwYWyxfWwq7XTCn0iCWSoKp
EUG4kNA0dRcpaP/3r1GGunnT1bhRMKQPdM2FnPmEi6vzNF4H8nK9TvOfKrCJ
gQy6eDL9P3h4NQLR637Ea5xkdU8KCArbWFcGLxCe4NA+LjdZYQWTXZqmlvYS
FvY2Yo8ipHgI5NiO0KMLDcdAgeMICzYl16L9KJ+jrUDhb2aAWXAmU/hgl8us
ZbNpzv7HWDaq8xoyK+rtCWLxxc5Dj77P6Ar7IlDRtRe1Wr9D1tcFykJYGyK7
3ucDVPh80F4T3SfT3PBVqOzmhlV64foDrMWHdrSCR2t31uEbw3WhrAhMMOhS
MvP85soi0IHQdIXY2pkdhCOa1wPUBX/UTf5V7Z/okgKUQJErQ4fN2kC+8oUL
MhAUVWtIpjH5NqW4pI856vt+5NlVC8qljKsndreP8nwPHy+UHtwVyhc7VFaR
iGe6r4NbqXRYtrYfj8K6w7J/+gn0FNGAidIlX4+chOIZWJU8AwvzGsCV1G7F
je9T1+wAuscw3koXNB6PpJRcwzc9ZVG8y8UsA2O9CBy3ku7awbFHRPTgn8mD
xMN22SK79LCZ/brPHZzOK9ZnklxM+ZEvzvlyZu6PESUOZqzlxQh5YpEOLoLz
QCF/ZMMpjwvmPhI1SDfVLAMo4z0qI3RXE9kKNRWWZprQmZ56vbbjCATrFSmY
uW5aZ1Kq+eht2ZuDFGrQlI1MhVLJv6869QnLWDT/YkWaXgg5TVJJQfFqTWnQ
0qPH5mfoB3o4tRkU6c4ZVNwX8rTmfPNshYyyOu6t7C3sHYBf/j/PZho6nvN/
BRGXe2VsqLT8ce+TwvveCL72hCZiF+pVyd03sf+Hxf14nnUnHSztWIMyQkJJ
mFHVhxTe81SZY9J5ufhUYyLoczWFndi2EjAvdqkv1kXMqXHn0B9KPxZYZjDR
Y5mu3b+rkWdkbc+WbUl63gWdtmA+rdBQrzxg52apsb+xYGAQ+yCjWYLpprEd
9taNkWXymxBZ6leH8lB6f89thVzG2DNi5UBuouaeGu54APJ/aws4Lf+JPb6J
JoU89F+dzj+2stBijXOFEQIkdKkmBkKStAiHfQtk+OHJGkGsF+y7WBM4BJ97
nQvHLpo6+iiypSfSLW4XayUOgwVuQ0mHRGfcxr3vR3ErquQHpfQEbAQ+LaSv
Anr7CnXRkWvl5OWU67+scmXhPWelaHBFVUxhV3AEf3J7M5crXiYh1n4O3EHs
StTFnNjWI+Fi1MM4fktYsvBZ+GP1nYaiJFZJWtqDxl86DRla/1A+XrCJ9R4F
InBwr3c0UpN72Vz6gbGrhcqkB7L7bNhEgu3z88ieBbr+13wl8ZJ7g+pQ7u0H
3s9Rr9RzzLxwddbIx6EB251ZgMg64n49BkOgmw3AGRe3aXUpXNkLYAXHCngn
ugv8qX1r1QrRrpLB1OkIGxg3HG9khU0LgblCereNpIs/OklSslNei0dLxmEg
WMQyGGIlKLYRmI5AmbWi1VY8tphcJ4lmc+sldmijeKNLj2+iAnT32G0OyWoy
A3vKU9t+SHQt6sIueO7HKvexP86E9vrLqA0lW1Sr3yIn+qnfPedeQ5e0k3in
tuTL/WpzBKxH2APMLw9lpQGEvcM3vZcaI7VhXDdQ20hBJHr0DN0WLJilHNBy
J9vJTI7zfZtksuqCF8hltI2PyKkYefY72VQVzjuKiUSSYyPDgLOe8HPqkUVw
/1iMUhl/1VW0mF5/MildwOJ8d6yIGIi/OIxnfQ/aDPwdyCi8Bk1b6193z0ec
8zliJ5+Z9D5V2gmVKCUXEi/b2BZRZzkxliVtudMvABgvAIPtqcp3dVN6TjSl
No4W3QaNVix3jmAbQNQDtl8wuPVtuo5JrnQPJYM5hd8jNDA8Ez/KTfNKGeSa
7I22IyQr5crbYMelAUaQqchXOLXOFU2F6TsBO7pnFbCqiwVfAlBEBxpfCNrd
qSy5afVm3B0fHR+qoGw/twf3cwqxEBW3T+orCXVgw+uYGH6GkZmBQbEzJhEc
WSqLc4DPkT3yqQWS6HyBPd7pvsilcFB7fAXFSnhdQcp9Dbvr0ovQv9XZ7ihL
JhBKBoq4ARRAnTwmP9WnuMoqlz+DikfmegGrdRvg44E2+7T+yG3W8TTJOX/k
WE2b0Fa7CcLLW0LfKEdNk2+J8rTqY4eQ4W5ss79+HOBQ9JrnOw+UXjmFMbWS
avMW/OO9Jmd3Ttys8ULzyI64AOpV6jVWzrw0McisQ9nldGaOOAcCU3xSX93T
Pfc7eoo4vIVia014lC912HUDAoBVGkf4udcTEGb0ShjhyVZUie4xNgseXYcs
c5bcTPs+BS/mVYcMDlhWGPWuOGaXBVjUy6tIOqqZHitBZCVHOkOWbATy4Mtu
fG0MMVJVAEG+MNbCVrIGYHpZB71kwY3xOSn+MmD1VvcEm4opDH0AuqGBIv+Q
/eBEszhh4wkEpP6CFISkYGkmeURgbMcNtBtWEuB8b6arMyjs+7mYcPl/bini
FFjjGtDlkk+10LpMIJppkuS6rdd8zyBcUsUdeJLQspeAV/eHKxGpNgU1qbVx
gJ7HluFEtD3/M3E0Ilz7hrxDLjWMivys5xrW0yMMTinBoMscL0Mj+ORHnEVx
XGwaWV9E083AByeKvxs0upF2Rudw8VvLavY+rXNkBNOz1pQYJ5Vghqnmt3/z
yVj9iHwis1bOx5vpoHcIEzvFzAXH1jGWHeB8tTjiSIremDFB3cbEdSH5tcN9
tfgBSAPWfPnz+794amTsQfZdbgoTf/Lo/1VSCJU3fcyy2X9CTQ8F8M2Diuat
bJYfBD16HJe+F2GnMskQMQzgpARhEug7oX5+bOmL64vJppOmv/VZJkHB9qIS
JLI/nA1NI3Vx6gNluWDM4k67Zrnvv5R+Ykz9NM1VOYtDdJ1hc5fRQ1UxDQdc
EbTzCyuVTHlfQWOs4oSa7DPfwKG8S/A5Ydv7u/D4JlvrAeK1xR/cyOlUdeMz
hg00N4LxssNxeUU00fO8FTcXYePpLXewgQmTJBingVd6Ddb5iem1XlHhSlc7
EpmTiHfg1fwpwML5ZjQyoQVu+SU2FFIwRFwPYlggsw6QOG181upC0J2EILPV
Mu3feP4GaTEi6fbRQ5apMiKdXkjwSIJb35zyR6qBExvvoPpuOHuKOr6GfvFt
hHxq7bzK/3jPG5wRs719vK0hMltpbd7YFH4QAkyNvm4zC0nDPK/2d59xAUC5
O4aePNU3tkHDI67esQwf0WPB17XqY4h7iRMqMm2tpt7VRjuiS3EJGEzHbu4G
HPmHck5AGZvafbWicbbiwwrc8OzRvV9CvBt75bV55mLLsZTh6+Eq2vC+oJxl
fcfAXlM8MGF2wg0Ms146+adkVzifariJlfLjwxLZp+Hib3ePtrBQbggvNEhe
UGerLdf4liH5zEaklEpXwu+6UmT01QsNegNfQXtLkKcVs0yXdivwFKVdtMXI
AE5W1hsIGQrHmmprWkpj+6Zj5ugNKKZ2OeQJt60ICi0X+BtqWAn3kjYFkCXg
6TYMVZ2U3GntgADiib5XUpdTM6gnbWtdJr6D0OuhYC2Vf/EFfpzBUOhKBmLx
uJedaYCU2QjN8Kkps8BUrtl+L9gbjC7UFesKx70kOCA2z/tzu0YBZpeQPwga
T1KP4Ww61d6eJLLdcOkcfT6HvEV7bwu8t9UbcIWg8zkIzMd9eel3vvUo29tV
PhLUxrAxFT7fvdjKufnOOAogMWpwy03D15rfZj232ZGFo0KnQ1l/lMQDwfS3
FVk8zEFTCHBohntj1uz/6D1AnRbl7VBwzVlYx6Oux5aN2BbO1zJyy2nRFZ2/
IEJ0kEH6oA8rRuyyoSBqZ+s8WnIgnQF2B8QVcATb+50xwgBlL54cfXifkzME
ta+xCFzVO8VnMoj97mr32KkLrH/zVGkytAoWQ/WAsiMa9PbJn+OG9mOn/lLU
ExUxQR8IdBRGEYEqWy5HXIV9lheDuzIuBR8pjp4FU2s6MIqdp3bdLhQuj60R
UGyqAch6GTKLabHtyjbWzn70wxuci2VFBzjDvSIk+T6NvDziDBsnAt8Q69WL
InP3GDDasfVtvGTekJNEbSwisOh3/esGbXlrTWAXv6I5NPJeDtKXKHKZMrj0
4q+wmlH82fflzEjG5r/IrQmr3dcjn0zj9Gx+yWtI6G1eW6KjLDeIjstMwjUl
uOsvUUQMognEP0HbHyq007El9pA/jXDJ7d320CDarMfAc/wwgyfCCfXd/oJv
XI0leZChqQmO835SS7/ZvvRuQr9ihpSjsvx05G7odaJ37tKLGD0KDpDS0eIK
xuEkWsTHcgY3MmRD99Iquc47CnrCoGoRhP77V/Dlx7QLUqQkC6OOVZHj5Zjx
3BFQP9YM0eO1x9ZGn+FDwZcuYpQS5qvJm+wti7Y6GPnI0VrZVgFdWdJLaLd3
g3DWI4LSCdep/nC22cleacHAodpssk9xh0eI3DDNL8sqcfF/2AQaZab3TJtp
lX4Z7SV0HQVfkM6sWr8UaWQvrGQ3oLUkt5iqEUkniLmuiT6ZTFUa5Km4Nehs
ljoSQA3jAdFTHTV4gWELtM2wH4U6HGpftSLDTmHrX+wwHWZUg/8BCTI5IwNG
YGXyQ6HCg2f8BxnjoJkWQy9VSwMJ9l92xf3aeWOJ2vOYHyZ2hPU9lDIpi4eh
5JfvXrTCnU6vCYbWnUeq4UsUHuQLYlpfpJ6+3lq9vFhVUpe2XavMBUone0ip
ZzyvBQxSISAZvPUdw09/f0urDwMrRagxxYvAG0EnPbvcJBHp1/PR5F6rQAwU
LeC72cR9lFpcqbwfY2Qq5WydVq+lxNums303e3Kz7FJTMWLhNNI59Yvaokol
cxbXPLg6xfsveNmz+0j79wYdqT41G6WQoqI0h8qW0RW3wM3AciFlKRa3oTJ7
ugFWO3ngQCe9b+OTFRmCKgE5A/m2bvOhk5gAYWl0cYFEKzS3W8D/HyLbfssH
A8nN9vnSGByMvx5KibtRRqLiHskAsx5sIEIU5qzE+pz7PMpy1xF+o+Iroks1
wIji1KG4hUuIdtUiq8ijJzkYgvccVmZAZwXJiGzjFhfEI0RlYj68jspFlWdG
y1vhwiKSyInLNyRMgBWnEhzL+MWbYyjGn+wog/pMtKLA++folTtIBMipNO5P
MLMDmKmGMRe48+Hr+QaXRUjrmL3oEtVANy7Yge1bbH/xSH/T412Xy+wCCNHl
REgfDVcURu/SeWNFAQkGd4TM0QERibk8NOgsMPGJit49G6NSMx51TabyRMX0
XiQUOwJYFJJ6YVucFsMYSzoIqxL/U3QigZm8J+re9CqKy1k9iJJBk6vhk651
0/L5mf1kwM5JCMmJRgQfEAVVXUHliNZpZh+htbveonMw+DUsPEAotkt+bh/h
D4N82wpLGOb8sXVK2inyYzYterJYsseePOxgNGtRo/5oSqjlnIvwEceljDLf
efNuFTXDEq6NGRyLRF9OHv4f96mpBiyYDv63K/GTh0JbTQqmEjoJUbmzapST
xlyTjJ9vdJHpRQsPJP/Bq/D0VijESuaZGL/7Pm8d3t3uYzUOEiSWYjr6S3KA
UT6DWyKQDnGWM+OihYnPTIec5yJn+YDmw/vSpuMx/+injmmDbwLPsOWV24xI
nmbpN0gC+TvMmrjjyqyAg+oSaXc+armtGQ8lXyJd7yWYapp/j0tVyJjLFSn/
d85K6ggO92LXUk9XTz1GkObDqE1bdcQtms7c+RdTHLLzOdKHqNcDmKCavLvE
D8dVeRmhkdrJ/HrMHPjaUNAU33E5fdeRmMNsXw6Zvn85RAEhSA0SSwdmiiQi
ZFhyo2ZEIVyCd3LrfW+Vxs+3nEDAJO50WBugJ3aYDO+MAgSNB13JkEDVl7Xx
584I1MWoi6opWLZWthV9n+E7gffv5KwSRYKQEJhcRw58ui2tyQ0qRAfM3WKm
/RQ9SihR8hmeZ/m/VbXaE8P29O1RzQPJ7gLB+fCusLXBK9f8bEcUYWOPZaHI
+0fIiP60OVZhaxzoMQofoXS27OB7EEnls/Btrdvbq4JIC21hF7Atg0qH5VMV
9c1wJHQOJXDY350S7jxNT12hg/fAk0BEUdYw5jOwfL5XiHCB7aaO+TZXsF5s
yW3Ed6umnZnHurGdk7V2OtqlYbCJ3q13rejLmE6OW4K5+nUoEHEF0GVznK56
HDwJq0QLyG0a5Oi6g/ipY00WxnkvL4d8FeXSR2eT8wyuv8PWYesLgF/YpW27
SKYkfbVVtoULSZ9dq4m9NpQitbr6XFFlp8YS5jXwdu+s2Nhv+dTdybp3xzxV
qtzVY9DFBvrYmKu39DxahVC3JPARsdQTrwMJK3iafa875qEyQ9rupZRC+RSe
ciC3MKjiHz758b9G3JDtzq38ZCz3UcUBmbwqytgoJn0nl3ydYacRK+P7Two6
zKPr2lQyUNpEqvGY7rtlkAHnpk0iDk9HI1kmFdk/nndlPdan8aVclTbbNeCG
DGbzV0mKOvguofrtIgUaUfbCl1wxxfp/oD7kiACkCpM2v0VXBoBWDeHQarVt
4OdHNOefAoXjyklJxDixDm/sqb2XvlAlUsIi/Hf8WTWsmq+lQoqqb2dVQvBc
3+MYbmk7+bXTbEGI+5qd8P0a6a30gEELDpkAik96JluVFKoaEuth4+et9j0i
PquhFuP+EttU2ZRnIeTnZXVo7r2HIm3qZ66Vw7DXg6nt08nM4/E0rJawlEoW
7X8cTGxJeKlafsvD9aEcyf6bdDqiDyKSatM/U1cMbaI5MeyjbJi04ekUdnAe
E7zh2ctvMsecaOyCa66j867Xrsz/Q/9ncvc/2qEMA7wGUr/1/TmdFgnik0j0
WXrPtdtON7Bj3Zb1n84on9wDV4GFOgZCgDZWm3Gm3lCsf/fezdn8Xh77ZmUr
n2V38Wpay3Wmf3ZHWl0UUDEMvy/1hbJ4h1xWpeKTFZlHmIjAeAspZSpulDsX
uT2nRMxaaCnjpQTp9AdxlisydaNqo1Jxmq6QChuRiWggvYdyiF8ojxaA5DVF
Q1HaaxwXgxBibNCJxG4bRtriSBas2HQ7GqWlNLqbauy3sMCWsXyDfiwAhcpY
l2/KhQ/nYme6lyrXTHQrhLxNquZjmA/EiYgIVRbD1AcG3b3oMoafaBBn/rU2
iJ6A4YjZgGBxRAWC3TCCmRmrjlUhHDzb+CpKJ5k278RcdqkipszyulhM/8pq
FZJecK9u6S6IJgkBMZJIwad1ZmOzRYkGYDjBMx5uVTbg1Is/t0Vfa4V7Oawb
its0puQhJyzE1wX7SVtWuAhmm0SRGnKg4MFaOGD6//GIYsRl4YdS8A5vxfqD
0yRhPGy6X3fQ1kAI+5YhXEL86YlEpf2yhYhZnznJVKCqqwOyZLxLKI0C6CVG
OsDPiOZ2Z0lf0H4hn+jm2crxm/M7OISMNfZKm6zUxJCWwkwsrkT4lKeNY6VB
XTRHqcuvy8n9sni9DNgBIOiuWIupqimv3LSum1W5HGLmY3vcNSeynhnjw9XE
GgYv5dTNKt5cVZ9UyhhFynhaJ/7u77Tv8nHWD/focGYoGZzmF8d3HidOoEng
tfZqT7khohyxIG4qbzpCHb+/lN8rKZQv3nYuaJ+a1mGAykg2WiZE12sN4qDk
Z4I+T4vnCkNDRga3/P/23BM7VODW6k7z1fDS92SsVvdLxtw++OrS3m0K9dB5
rLqJh8oNAgX6krRMrpPENMNh03vy6ASYw2y9lzKmB9WIlX061BnTkGolBtzH
GdmWRF3KEPhb+NmSceORG7lpokiPTXPnI9dSbNdaJheQr+orUVmlfPKE0coW
JsAERpP5sUpWZIB+0XKk15bdMeaFo1o+6zzsZiKHIK4S5bexhmtvL6rGNUjS
ogIHPFLRFJxYd/BuemhxSI+b67V973R+dJ3Ss1WywJe474G8XnHTfE/fSiJ8
jAmJypjyIdRcTJFYueL8nEUPQ0e/HoANFWaFIK+UF4zY88n2Zqki/EZ2rp0o
RMZY4q6SLjDIzyJVOboHh93HA/+/1mXNpR9Fjo48Dj60yEO9N5aBaVo3nqFX
gYSReJozgUVwoQF9pR8yEWUVpwP1PaulwW53F6ZpUzig8kNRG9L+P7e3krKT
/+3OOBoYD2lsQtma/rB4mfpcuKQ5xtYL+fwWCunuTwkJASkDB5fpIJO3fgbh
jUJ940d08gew2Dq9cOMYvSiRyZv8SjWk+JA+ZkaQDEM4/d/In00YnjMihWlK
LMf7Hmq+xprAAcCG4JBme3RcefOIrprrxCSIphHR5LiL03B5kPUdIRAAhUd0
FU67sebngFpqE2lXAbG/9p34FDeb0irkcyVS30e4xcoTfvSiMmekjYTwMqbe
pgdzt4rxKMXKLve7RRafLCq9mTKXhgMGBnqgEKvJ4RiLOT280pZo5FjKnyI1
l3IvtwExVtyuvT31GDQNophMdx/sKqJLn1VVzUFAyZhCbPXzSVllcMrAl7bz
aNR7QLy6WQZy6BbVSSypK75aURiXkSn3x9OkXzhzq34D0n+EdoSpjPjtvf81
dihsTf9BQtldgOpofRnTH5c1wTvdpwH260YdpYx461C/KKCcANAvMaCKrmrW
aO5cIq5zGj0ulgjC3f2/FjCQpz4aDbCZmsgW8/cYDZwXJoiq86X4Od1GOhzm
wsumFFMqTWwYA+BXgy+EAtmTnQCGeT58NmCXN1CanEFnBfD0GTSNyyDvlhnt
L6jFcDCGpUwrLDxLhshYSG6hIBY/JAfwJlFlzvjZTFgq2hM6wkpIVo8oi9KS
sGU1kUJIsq1o3TSbE4KpOx6F/aelpmf4XBKQ/x+KwRTUN4acJ+HeoaWDMa7O
9r7L7PYCrqJTysyJhuqVXQ/q2A9ZSWp307UfDKecog33dr3EvfVXJ0uYkGqt
1AemvSxkGkN1Y66A7ZCun/rUjTWJfPFfXsEEXhpVU+5NOdcxHyKoOuUEztlm
4FULgIb6c4EL+8PcTivjFZ5wUjGKmW/8fDF/eqFw230xHPLdyFtsQFyebm5X
Fc2SgAjVuaE0sISYZDLjD/BqH/adCc3hjgNtFeGiAmCUqgcae2YYX1amdYnr
HP9SRhzQuqhB/ijUL2rkRTYXsGhFdYgv4Lc1qj4iOVSh0TFWeVPCinP2r//o
d0QbunB/5I977zuHNgga+xBrfXdFvGZd8d7tZU4EvAUhffO6J2v0+F1w9egT
KXmQdFnaQgjXRVCGj0Av13YkM7oSWC780EGHqFeYkSkGmtbA6z5vymRBBQYz
P5fT2Q9/E4tuYHcnlH4q1BY6yYrCfciur589OZX5Fp1+qtgthuAsZ222xZG/
50qEJOlyKM0Kdq+2B9h1BMGHtKG/SJ0n1DzSI7PeLU/gaW4r224n/0xbkZqL
DUEIdWWwUpN8Nkn9pzhtejdp9bsZeakjc1zfI9bznTrvS1Q7y7PNNEDkNBll
EVqvOmZY1k01Ld615AmwCIcbTqeVCJ3SadNlJqw4g/q0JSGqVp4xr3ZzFvRj
2gIhNWk2EVQDEUtLVjiEEz3QNIUAdNojcXSOKDofeQSOy3ZIRtE3/jBocg76
e+9fug7+YpAHNf4ytfeq4vx289z82dedbDIL6AYa+FJHil1SeQD5pxjw3pGJ
cCOcgcKevshNcPjT+INv0HaqZ46PMvqNHd2gqhYSJ1t+WqnRcpWyzyMz04vb
DbSxJqM76hx728aKKnhok0z3M70Kbl2d4/j92B1SDwWCyggdwudZ0NWSz1B/
mxvqihPZ+KChjlPO52ELe33DrWp7nac0G6ZHQpYID3/u2AfRluDgDT/sHG3V
JdX9THMrsvXXNy/6ahGvjYLA5AJA4oR5va58N2i3lRIKoGJJq1rWKCzK+QXW
RtCbRqP0MVIs9YQaSmkjfB5cQwjOk+jaUdcnyVvFXcx9IVcBrGJBuZEAkaN2
ulGr7DphYJRpMAwmuY5SIaciZSWi5EJflHHGaN6O50UQKgPAXNKeBpdkjGdf
CK3wnYdfvXZoZJ3wSKzqIgWX7CnEUS8WSug91f/fuLZumj4l33Bfvd3cVPMl
03rjGGCImG0gQTrUZoXGd3DcE1pfc4U77N1AMr8CDbMP3Qo4FKDsUnfIzPhx
1jt075BJZpVcmkXVf15xrsKpB8PrST2i0ww8SxXezROlP9uqSVfKR5qi6l5s
xk0WpAl1ShB3Tq85wXTe6wDVyMADaJbXRDVkize54SaCDvRxxDY1Lpll61pl
w8UfpAZ1MGUWZR2bhJqyFiABMX6qLvHDnt10D7aTtRcer6ljxcBBz9LN8/VG
7mkWf/w83XAmZwk3ZcZib4b/kBOrMviT36Lg/uRp4yrrvOrRiinrtguuGCzV
Iq2t5AHFL0UlHMsa/Tz+BA/9o0THHZfcMdPPFVE1Hi4NatiCW73JzhrPD6qx
jLZjinc5+FJUQHzwUvYcKhd4e2L9cl0/XkIrhsj4tZy9UI1j4+8j4JVrEyuI
OFkyvmodudryAu+x9AfGdh+G6Oz6O6lNzVukpa5LYe4FJMQwpSfJl4BsRgGy
7PGH5NndtV6Hmvl6exXu6L/FSHHQNnbjIgfBN4d337NPXh7pRFkZgwernDP3
Gzv9EO6CuHl2pExrceDoZV5jS7q0wnOryBGJ7QFtkAu2aaVz5BlKBGFh1WBR
ZFNNZNl6fqZM0sZexWdpVsjbHlASLzezfn3MbAwQkvVX80fXIPIWG5IiRIS/
iCCeAyspFP4GUlRiHE5n2KNDGGkSTAz5A4pGzm78uL30c5fXdURRUtOdjTAL
NsHmrgo7OdALnbsNNhvSHLTVnV9GEaMmM1tLRlDKPv3vUyExruE7BSvi9NRt
xppAXffikZq7zzKTYOU1J72lbN/6QPgsWo+PuaHW3txboMa103pXlN2VJcIV
G9u3qFHkfXIB7UfeVVRYRhkclLgAbSjKQKgqrApp7uhVhr8BWwb1q9L2OUNF
aj0tCxBk4xqyq/cY6H/0Xm6AAHsM8fjYgGQbX481H0hnDJZZb/8xOxqzby36
QuTi9YKZ4uBaHuBUSSL1pB2KHOMONrfJkRh7NLtOodOPNuE8QJH2YjnxyvoP
CGPp8vRwIxp+dkbwdpZiDemT+OD5PCiYOr1y+RRKB+O8wGS3W6COYMNuaqcE
vOmBvk2fjSiuk7OE6ou4EvLu4UjsWX1sdAELXmD90DXZCdQRIxYFYR8Va26f
Vptu95pEZ4ztklWha07BwiapinA9jAmsL5AhKiNlzoR7//fqrKxqlN/TsV9E
C9KfvEijsaD5m2lilZ7W9Lc84Jka62cVvsu8I2vLAs65CzCjl25O252SytKO
pJKe5XZcJyZunt1OcUVeLMzRP5nMoSanz06UQWZ4klLG14bTdvahkgJKm/qj
+IsJ2BraWmti414y9bEqe6gZ4jKkxMSg0pq3R9Ylf/GoiQdbLJBH1cpZ2Nkl
OkbFYR14HlX8lSD1ZJCG4t830TU/Az4F5diPiVPEMcb6EqsfhHxTvhkJK7k6
8EK2vu8KwfVJe3sq2eKv2eUeW/GZyjRzykMEmglUrTFGZ26ee6oa4zQYBW6B
Ydg4Fa9qhniDhvygh47LUyZ5V7FVnAOIjVaKMcHMyKs5223ax5aRBp47rabR
FRHDaeMk0w6Qimb7dqNLBQiDC43BWgTjZbvgxkyqNSLLhDb+ZBq1O5QyltrG
gHDuWjvvXcrcDQg25U2hRMXY39bhMT4iWQKcDEuOAjnKDdrLgzciFx7AQXih
A5RDsh9RaWPXn4mIXYac1Ad5Ud+j9FCcQFA9wfMvZjhqPOB7pRcnBzZdgBnA
Fb32iosM5C4LF9P5udS+QabbXL2bn4MrVUo74P2shH//9pFspj/1LtcSHe6S
xNUEDX5x6XgABGyT7YpSqnm9B1oRQhIfZeHricT4EueTU0p3as5qpDcB2Jnl
AZnZLuF0WfbulHnUjwr2smYeX4XZAcfUjlFbnvMUo3Bo8Vw4aCwRZ2J84ZFE
4gKzaI8klMlJpJRSDwDzsDRlyvbbeZ4RR7D35o+SBRuAWjUc7yuKhFQNHKXV
jsiuvpLg7lbaDSAJ0TUbNox2MRAFnlJCQ/B+3fbeBD6vx6oZ62Ht/Zav51e8
6GNWtWUBwRYmRyCdnxaXTTfgPAkesCcstQcQpF7DZB7609yaI/879XW1Gnln
i4fR4Y2NUBb18aC40wJyyhdL8aPPA6a8xEBQyFMaoSF4M7F4JHoeHcpjIkXP
xsFj6dv+2Dgizk/qdnonNlmRnAsoFojNtzxzMIQB/OfXtkNPf3d9ZHGf+PVp
uSt8ArbM885BDGac3qZxgqeifHIDbx6L/uOoNGUr64+/ipxI+U+g8GL7CX07
3QJQiJ4v+RF2lVL+qtey8z7J7V7lKqI8Z5cvg5Iy34hs7C9F1XSbe+MxkrTW
n2rJzd3GszV79L6E07HOIO2DPfY5TkQzl/C+9UyVAbllFl19/e8fZ0wIve9R
YcOIx8kEgzj96dauZMb0V0nNWqmUmCapZk2DJfRuMVC2AAsYHqhMeyApZBay
dttL1DILgnVjuP5YoJVnJ8FieOqt1n4Z/XR3yExcENj9DIXAxs4jkvPV+8u2
+j3+tVPgHEHppB/e6tSov/Zk/wQY02gQInHVtxkMqnwtqzMxRWeyMyhPuFhO
QyaVnnvlB75r7cKkXaJhKH6JDm2R/mvb1eCq4VJ2wPKP7gBTuyKZdEH1NkeW
PIRdD8AFuRJDCX0ppR8JcyUaXBgSiFUkWGw2SH0caU53+0PdD/fidS7iIxxg
6wYC7NvUv/jjuDXGoS6eK5Gf15P9ebEBj4bH687/5xQZ+/yA6I38xo2EJTGv
iNoiWnaqoxcrkkytLeNcbwJG4HygBHHLBgU44SbRdB8ZoErfBlPyIttk/uoQ
fLqjy2T3ZYJ15YKwAzOL/MTunha3nNBEfsm1oN5GURhDjODIlNI6Oxxk67q2
Ldx1m8IOTMGGi9C5Xjv8F7Ubwax59RiSJKGxVpEZqzwR8LIq2vORCYEQO6tY
RYshx6kbkvGvo/gKOCCZ8jw3FIiIl3IwX6EMQuwp4aYDkRaQge+298uf5Y9N
M0E6oDseCzkvJOHfReVIRqA4AzApWmRPEYMMjX7n32vJ17SbEkv3aHO93cFJ
DtBebSiUW6tOI9MDE5NpKnKJNTIChYQ/bnelNN1VNv7abJLMJC7TLTVTTaoB
Q0jZb64ggMAhqS/jTgHv8JZhBNkVfanuBv5bAfbOe/5Kxy/OnrsrZJnAPPIa
q8AVP7/1YpMaprRaPI14KWanbbYrmBYNcjHTL5uq/+J0TCs2gre/PJw9XYoR
qmNs1vRyweRswGIYP+HojN4ANdGQ9TBJBQpdJ4YIega6IndNovy2clfw94vb
jieYN/DKFIf/cQNRyS4bzUO0z70FFC8U4ut7GVyZuFfFXdsawqHAENhPB4Ol
EAxx18mielS5Xm7cGN8P+jZd5nzkDK0BwftLK1JWM7RyjAslkVbjRp6p7Bv9
5aRS/9Pdij4IB4FRBFeuic1goDYKW9PpC9vm4fnq9PIMo9/viKffpxDX3ZEG
83jK7RbN0aTUg2ACfNJUJSQgfFbycnLc0koR0PmDGvuv684TjYG7pGnZHxlb
B1HXzQtJdQqWH8BE2FjIbdaIWzYrDxjHtnbUA7Fb8mC51LNdSAjshImurwt3
kiBknM8y57UaK/OnFPzrLB6NFR0kjd7MU+PpE6pD/A7S6C2jr2Gf8UYYo80k
yi0E06KoGpNlLeKWssuAEQKaYfr3EaEEMUUfkIbM3mmnqAPg8ud69xWzlpuY
WEpQy8kQTLdGzY1nFzG44j1w54Fv9nDTH9NZVYBaB7GszayqdpjPiG9kuB0D
1WPEGItH2dw4zkrq9dWg/YbyN/B2ZZ6lXZFAxJK/I9AJu6SK5CzgPFrvN3V3
28TIZNh5ZpjvSjNpUP+kGO8PAS5AT8fustgqwnY9/xkQprzk0DncRDQR6Czz
Bs9SxnN5zks/RmlFVLOHcudNh6hErkgQCAQ50GSxkFh91VIeyb+0U6rLLh5q
0QMPmFxiaxcPN8Br4DKWpEHd2NfNNbAs1fYT3EBbaKY+wESB3au15iaPfjg2
V5qoR5rj9h6TuyBaQntP5jcHr0zSkrHklakJzBqm1kcpbUohOyPXx5Sh16kk
a3bjruHNAZmYXHIVJM3CZwUiEA0vpy/xlke9Ly6Sm9lXPrMVqxU2bSUCZcHJ
Go+PW/44O2JJFAE0U6PCYqT+mX5DTZQc/uC7z0Jtgm/YdtB820TxT6BULsv5
R3OraFLXod9mNDVrJ1TluGjtigizBmLz3FDDvClzwSqbb6heqTmNvSVkkfnb
eyeSnL76THvxFAVVtoLEilDp34UAW9N7Pu+4uBWRqPFZemZu/iadiarz26aX
qmROFI/9a6HLk0UlkHSTEP+z/D7/8fu7tEcWuAwIJsDBx+fzRIu/GSfsv35h
J8zV4m7HzyLToEJpc2/0W7NbE7nhzDz1dZZ2DgclVkO2vEHoiI2iiVdIrYkw
Q8BsMPM7ck3RhyMXAfv0R2Him6IvDbE3/Vzq0ofKi8iNFOzXrrEICCN8+eD9
eXuEmWWur+SBIbmQwIK6Bhd7xrsApewgdIwSLAOjBxvTKIbjIp3mZhcBasDI
r0nsnzjFXz8vC/qt98NiXfgi4I94As66Ag+VaGhQKmw/N8pzXR+IAk9YHIFU
Xn5u8obig3tsGBsLW4J6IQoRmD2SPUjeyGOr14N48TaL2GUa/FSW6PzihMIX
tUGt2fkGOPGSKsDgBCls9yFFuj4z90Nvq3MFTn1nQ6Zg3mi2gxgFTxxh89rv
L658NjeluhDTLWTSKaCIF5KBfX+iSLb4c3Yh9J2KHdjw1dXq/yCutduRyddL
4zWqPfGDg4NMdTmTzu7HJBi2GEISaUlIOU6gbF+y/F4ovgxDPHr4i7zM1ai5
VL6Lp5hVHPHiR6PLm5okCfYvVEjGy9MZhTN9h8iRmL9bEmfdupBK8Au0dqzE
+zlkE2+K3oVUtnu+6bO11yeYDYUG+fMwwezjCoBynzbDTHbwPv3UeANBwQx1
ZZU3X1L+vlNCPABCURQ6AOoWTvhing6Ck4HG2kgtlsqqFXc2j66YJ+uaLayD
XinKYWEYIhLsKnWiYnkNEr353QEi76UtbUqjEAbTSaHqLbAo9z18+Khf05A1
PAJs9y/vw0sgmACL4De8CiW+9GTvPU4vYAw6IZq2z/auYaOtNNnykA71mU5W
y3eGaSTmgifG12h3ImOyobDIW4Dae5ZYS2tZnsdmizOCU/qTG9Jusz3/l/XH
Rm7Q+rcAd/iT52gfc8iYTK3lWXVYPHyX7DStSTALdqHMHwC+CrFFcjrcjPU9
QXEil0/gOY+7XvTSGTORvHAk6H7FEm0Ri8tQoLXAmj+VPt8IE+lpGyfJ3LWf
FrmNQK7P5NliY2bLDNBhkQ+jLsQv1p2gf2Zh1Gjo278f6bcyquoTENNHpste
9cqouEKdiKnwesF66tEpsmpd4UOt2scP+jqqDWQBQICC0utqnnMUDw0rMa3T
TA2fiQh1qSpDBtacDoCmWMP5tRngaaUGLO2xS2bA8NJp//govYZ32beg3qpV
wizSMQtVgTdYhMfEs4OdJUA3NGqcO72bwe9pxWUV7741qm+GuvJx1oKnWK+y
TgFQcBvlcjlr+4mqSkOrKJNt/8PbF8om7tAArQo6FseErgSDrFR3ce04XN2v
Bm3JUI0qNVgQbqBU9/B6LBY1Hx8UfLWvpB5PHX/By3arNJ39L2C84Kc3huvK
Zqxey3K82LqaOFe5pEkUOgs80PrdZiWnIKy5ty3nxw83VJM1DpT4gITrPlyw
sUi89GD7N8R4NULoQGMNYOAF9dkwIpAtRPVvryNmKrWTq2SuRl6vJR46d4xi
3KSLEQkIqXHVMG5d1UCsiKUv2xI8axCURDceFI/zC4lBgmmS+ww7TJoIFBYG
qIkQ1l5+2KKoX3FC0YTjLnBVIBAVf+ZfDgjoV5ym4Iup3ZRhZPNbOoKHFTPa
A0HXfQwp7dlVwArHq6lwem5T899TTz30hGP5q5uQ1P1hHoc0vQWFF9epqgUf
EqMXsOybAqMU2PW5qXJPDTPfGqrfmhRF8+0NMtnjGc1p7BxMfid5s/YRlCed
7duVux3UbaoakwT94KA15dYBXAStkZYgQxUlSWLLjzpsNACUR34QCLxjobBW
hsatKHlntLHrJ4+VieQIQhgcHclB9hyTOQ6Ur0xtNKt7Bk7lfVjl2IuVgvU6
dx7jULUk/Lxs+E8O+AMDOSaw1WQ7crFwk13ImK7JkgLjbqia4i8It1eDUtWb
m6JkWM6zK7YlGkWu6DnivtQidmHGOPHJh+C/h/vYaC07tGoGRfBrsOKe6x04
O4HPIPcFSS7Zf/uAaPqXSoh0K+9jcufaTOaDovCOC53GIBLMrr3SAMkkla4u
lMQh4LcCwHhieVO97gJVQPt187qPqes/po8WeSKLCLh30xpm3Xc5X4d65zkZ
FQV0/OPhg9wR0st5WLjNPUUZZsLSROV2EcjvmNJYG4l7iBpiX8uUahZsIX8S
g21G6NQPlixodMG5Azts8yY73w3xsOolqXoOtsAUnh4RW4CKKXee+HgWoB39
NIl3ZFrKtHmBDKCxcODrp8VLtCYcSj8I8aidEM/+/uc0G2a97Orw1TlGczc/
GWMIz+0ZgYwvfJhh/R2wMJRi/62vq32mh4t9zeJN8DhsDtctmRtd4O/3+YND
W+RdyvXW+cs67C6vCBQP7TpGuAfXEGXpOMllJg/1NYMOl4NFjKvWnRIusrE8
1QaaHvfD06ZY2He4wnCHQqyAA3KhqJ3rKZFKCWcMjXBzj3U8Ztkp+fHp1T/a
XEUbtmr0obpjnIjoJ2nsr+4snRPVcJU8dp7kC4KVMI+Z7mAFSg56NB1ZGOAE
/+wUAWn19n3HSklv6kwNqxCfX0YHS9J5b2c+EM5xjKR3lukI8wcxXkQqprbU
KXzmKVpfZc7w7lZ228MmYmW2ZtinrFd0dm+3knIYkjybarZOE6qxviAtOSjP
BJH2YVtHFdSga5SyTu46+RxRnC4N74pLO1gEF9Gk3uhGUKjiTjCsg4NGJG5s
eSIe8Fybf7xqwPb4G2q8elPaBOSwpws0S7SlJtF3znC0kgOJEwpc45cEhPEi
rt03F3u2/djAbtVEhFfC55Wl8kSSvE6T9hksxy7CTqIvzS4ASgeSqWsV0DOt
ipciHRzQ9NqXE67m+RTU1ggWkXNbdC60GVZ9Ge0DSsfY60mpB7LfGJA2EJTs
AtYWRyFzzmjIX/nS0jmYbF7kEZy4L/fvX6dIwukTRQ89SCSacM9Cevhis61x
ht1ZhAgwXGI+x3gEcRx1jvheGDlJS1MgDxYa9JktxTxrsc6snS5yF1rQphJN
2Me0RwsZxocPjzuDgxh9iiTjWnF8ueS+omzFDjZK4UoRJYjIVY1E4mnVOj5j
gR+DBkiSx3z4vFHUDV4+r/Y+9zJjgDTbKCfP8uj0I3TD5NATW96eBCR2tDZs
Bkxuy2MZ2cjZCv8z1hllOyGIbH1bMfXajjS7ylSJ/kiMTRPv3jspWcEkirbp
SpPUusLICfzEvlXfp9iCN6KKlSmrg00aMOa6CR5JDLLrn2S49+bgbXUbAgiX
eQvyR0w3o/oGMzF6HvFSiZVrEyNuVA7Cce4eYBo/0xM8B1+hRxsu/ter2Ocf
nomTiDJDWkpoHtBLqm/QHaRlkDmF1GAfmjhXwUMD5v7Kfz+fxKtPTJ4uTYnv
XNzL9xNgaAFb2VXZWnaba17CgZiir0b0ilQB/IRG1dYX8MwuZCKguoFUly+Z
OkQ/jHEbXqH7pnUIeSOInQndApCNYhbyfw3/OLwFZqqHO6grKYzYuevC/8Bz
WVc59HV8q3h3/2cYKlKh0C28xLLf6DUv5jyKGgQnu4fS42zdqa16swssMKTU
lV1lRtcerMqgBDCKozg5f6ylifNdg7T+BjI6HZJ4u+r2hKcBwj3UWft7SZ/j
uKSYYTrHpARtbtNb0p4C/fs3NbtgKdhNU2Uo/pWjJmxR3Sa+P+332TCau5BI
9GJzk7HtZBz2i5qtYQ19oXkkolLUey3zEjF+d+V7cS/x4hSCrwUZtmclry0N
F9bQ04gtmkktY1/2YEGmhRnx1msw8Zyfhdfn7KSZsGyueseSRTE2TytdTkLJ
3mK41oVX39cIUNKEDwPdjiJRifT0/OrP6QjDQUkxsXCTWxpZ+Vgr5Bz+nLoq
l27ltv/mphD/15Y14PL6+yRUtov5CiZJcCtXExGcoKFiATd+gKx/mrsMNQcG
or6widEsJwVRZg5h646BzeSULiI7/LePClL4v1Kt2/fWckW5ogIzYKuv8brG
MsdpOavWlXdpMEYj0zHrH7vYewUCDoqHzj5U1DzCnWshpl8fZlFU/N3TFcS1
/Pw6pL+GyJfLK1UUVwoRftMIeXY9Io1rlb6MSoivD8tS5UYZrrpG9YZlHkCc
aK6JD5ewS1WhN0kv9tRJg1FAI0y+JQeWH+UNlXPIXZSfeAbNuqpa5te/i2gK
6RNU52ZEFb2SdBuQ8fQGo1XfptvtfG7RxcaBCotUr45+CBvgYZEjMQFQ+NZX
PG1Z+gFVGvnUvbS+9iDmBj2OdfeusEow3moC4rYZzbXgmVA1zhWQjbuDnDtX
h40/SKM7Re3il1Cj2OA0cm/ZZQNPS6VGvFCLNYbnu1K7GNKsLl5mqGe1AGuq
Ztdjs0oS20XZL1fQMfUK/ObrM/3UMrpnaaf/gNJEBQ/FI6tmYMPBCWTm/rxu
L5cSbbL4TPoSOPQF7mPJRxOCOkLJ3KHtSXo57llWFWvUjDbAkk6x/WIj+qIp
cvKjQTWLvzuOVR9zg4bogCdZFxR+tYXOhiN1hbOgK/PzvziDuYDO3EE/lMsm
9PpTL8I8qsqnww82Gz8+LEz/JsCaK2WrQ4a4lpZp6RiJNqPqza5d7qg0tZWX
nb526FPQJSnJOrK/255jILoT8M02Ik4fNbt5JY6AJ5XBYpVFKO690gIaZbDA
xg5oJMGZhV42fH3Vj9/TADM/7d/31reWlL18CrUWJgqiHuDptXhjiP+CeQdw
YSrzLXBbnH6PUGYc4yAE2GdNKul9KqzOkcHoEYLDiZLKj2PQYBtalPohcTGJ
qeNw75f7zCpKCdB7m5K+0Q+Kv2VjU2/ebn7+uvwUjdj7oCwY3kTC7GSOYn5R
nwLRTNI6KZ8QS6P7K+y0lC8PP1v48yuH8TcMH+/H2i/rCg+qGCCbN7RBxfwR
OjUY6SwIBne2R/BTcLWorNfn1VWKMTmLKdyZwyRl3+CjGvcif6B956UzUcs2
V0rQMcgfOhI8lnXdj81tucrUCKQ3h/MOo0/ZMDpyTkrQBMjGvSwL42DfyZLg
xxhMot/2q517y4/RE8g5OmRkh4jkwdUOsHa7KE/JZC7xoxiXVPxkdoq/UVWM
zfrv6O7DygQ1PdxcpX77zOw9bM9O8v9B6PgzHuusGteQWHLb91TI6J4G1mza
5bdFERFkFtm4kIhTLu8xU2g1awR1Tg2PhvAPJnhmF0C47e994DpaJymKJmZP
ymz2QR9RFGtAPQsYX5LzU4aZG6qYTWJuQ88vkTDFEfDblU95sSYRShhZ+zcr
1V4tFDiv4kq5YlNuaas4UJBQqnRf3nylLMxkZlcesXlcUynUxLkZ0OguMart
gWUIsrcUyjDEvNYZAKzz+fRHmth/a/vnQ/xnIgZfv8JxVpWvpxWjRZDKBUXb
lpJU6IXpwb54QeD6jDucnx/YmUB9svPeQ7jiDMvpg7U/QqWJnOfBZ2folhUO
yCjjaRIAAl5mEEBMOX++2f/mFkgj89N1+lWuNtydGkRULKXltfbvR/WvB1yb
fACSbkz0EdsS75/WgNvIIlTg5HK3OzoIkpXPGQHTLXgDgtx3kwfl/mMxjZoE
+oNIV90Ln8ebC4wl00pJ4PBxb64+f4S61bcRB699CQ04PmHOpL3DB21OUk+A
jQGDw4zlznAatTxuYV679SIaQvPegFp5/y7XGkWTpmLE5rFHrhCr9s1I5tph
boLEvid1zmuaWQtrYk7Xr/G9TwpTA9nq3ou/tHer7kkfpk7LTWrvdposU2M7
k6qC0JF54axzkMAIrqNFFwzy5YGk4ghoNq4e0tH7R1gzFDLoBELwPyi+a6am
3k/VoWZJx5kOAeQumMp94ZkdOiDZTePsKffguV06EMcYRWEqGx24A/dMXD11
7Jfe/jYyt6aJWNoxo6Nh4/XktxZrkgpxzBeEk6iPKaMbRYJFkpPkzGVkxXUf
eR9VXVP2brp8h6ENpG/l8ifWow0XOiW+dMALRQ0dNT+NN7dSTcwSo1FCPqVJ
90i/D6M906427TXf6a7A7I+5KwrOzah3b3uH5l6uUC4EGLOJ6xwjSsymRzAW
JSUXrU0a7MD6+wKn2zTfSUs35VkhT3LDiSltAcxNlbKrjNjxOI9Ld8LcRruv
vjGzm3BAZQMocT7uV6mNKZdNbU2CAxky0yAqvOmITUk49I3oyEgsGfwY1Xn4
ezPumAlfjQ8con3pVbxejxnqDYuCoTZEjE83b9PTR6ttJFocx4NkrfgYsbkM
7l5n5TLx9C8nHnEKucbuXGFoDKkWpJM81XoVpzBVJer9z3ekXptOjBSmA4qA
zK82oupLy4W61e14MzCO3QNNV18HPYeH1RmfNTBsWcRcfCqHl3IBaIihaENc
SFehffqyokZkbTMPR/cwKxQ5jmy8C5Kst/iCOyCbFUWLrGb8iSPsd95g9+qm
kXIQQGlSv8vgQPnlgyYqSk22yjQQhg+rOA9Y4xv29RSclZ8qnbhwAZR/FsJ2
yiOu09JfisT3bU7BJmOJdbUOCtapoESXuyhTlogejx7PRQaeTWsbbBzapkcD
sIo+CEt1TRrrJ5N4rwUwXQ4CYEGYJ26wpPL4sCmQOhCn0EaeF4NXBSLuvdmL
8IP/k2kmokeRiE7HjGif5SG6yGubyuUmVALUKoJFgy1OmV6QC8rboBmSSnku
Lwa9wmIA9Vv7XT3DwJDiWQuxnS2pwobIEKMylracfae36YnTkbuuSkxTqEhv
s/qemPPEDjQwvcfTZLqe0xB6EP03T/ujHOvIV3w62/EvztPtXe6LvrgXrFcH
DsTG2RZjnZmnygI1wlR04W+bpJScaYcqB9hNiJHwytywJnklrGs60QFHIKLP
W4db5Cjv9rAOOmCg1wTqKfg5rWxZ6vEFaTWJyTPKsIDGQw90v4bhUstIEXt2
SPUScbVSvyFzOXnG6VOIUNKfVy3a4gEHww/AnwmSK+Ob3xYURZ9Gn2Mrefbd
wMRGQEYM6b0xIAxu/LekcGAcSDQKAbqFNlLOviDuXc4kwbdOU6X72Y1RLIff
NvN0sR5LRHQrVNPuY94IRdxWbJuWw8qC1mBxcrMoUT6ZAiKpjU7Al/CFBO3t
2+wiJ103OXqQ7vB8zRlWWt7LO7ZXpkPlUSh+dHhnmgIyvW081wjQ/NdmlNhe
5QXIMMcLo8N3wZ9sf52ZyFFb91WG4bki+m7xcbEue6XCF0T/SF3QsDRV0TAA
Fa2X5ARiEF0lYx4odMSoNsyA8hNS6hJrhEaMEkrYCWm3v6ioYNai1hOjXfih
4CLv7Zbuw9IROQW7Mvb1Feod77W72nRNffy7hJyTULVxRYv13t/6YvHoQfbG
QKfVI1n3dgAR1H6tUNVxUveDR8etI4QeBmqxTmn2p6hJdf6GecpRxF9KkW38
9E5vdulr6J0KRK1prprJgbstZiTKx4Kgv5plleuYE+eebqRDqElBkuF6k5oE
bElNdb/aElW97DwTbOntDpdXOgu/FRHmcqFlGwobe9NaENQEFo6k74A9RGaM
92soufU/m9rG97YQ/AyOqU33MlrhpdbudtM7LZdRtmmD4CDLAKAfvEUGnZxG
VapuwjTgkHNiWgsWZZmv/Peb9lbmjTQ/TS+VfaheAa4qbdZg2axxxZ2asDZz
QrEaDLoF9895+elHHU1QRo7lTI/H4/8bFWC+2Og+F/oEg4+KQoJ8fP9WT7HV
lQDySYLVuAgI2l/JkmmjTC5UirPQw8fZr9LFQrpZjcDM5i78svU1WT7XC7Py
QTfU3EZMtybQZP6Kd8kQB1E2T8HwZhdEz5QVCZFXEij5U2Jas3M5WuoDFBNF
x2YTiHqHFulq0QTc+bk0E/RqwqM6fivVoha4nUdBiAtgKmgcXiiQrJ7QXB7C
6dV8E3CvAGEfpNVUvdg5fPAHxq2DjImujbenUFmN+bsCKwx5R46X5dFctyEJ
B+0wlEisQ73hjLGd4q1Xd4xOmOgn+CqTALXkYu9dpT46biBfXQqMGaAY5l4X
cjFmXjXtmGoIlU6fBBnNjN+LWJK0k8rXYgFKwc80QQ/bY7hM6SAhwyMLZPyY
zt+n6JpBxiAMzN6poaHVLxqpAeJ+sjbv/O7QuVBZTZtayF7sNrjeES/8W4w5
2gbaVGcMEUxDWpcV5WGf+192ITRV7sg2BJ6+emTW1eRH3Z2xAeC9s98gAtIf
dYCbQNk7SY1sqiTl6wV1Cm5aO2jeYCmyH1zSAr8vox3SY9SSzMM0U0oP92wE
gL04IcMQnMDQrK6e4zi2s90/Fu+8aZ52dPtXI8Nf57X0kEs7mNxQVcPLWwmU
5SikYAPA2rikE1hlao5/LtocONqlm81uKTaS/jcZcWT9IPndk05ydFjx93al
GTGebHUcjLOQyuJ1fY/LOs5kWHEEaAiRp+R6evUYLEfr2aLK+iFFaUAjHOns
yjejh7NweUFfZ4cr6k/yf7vFxKKDIKGAltmkfIhMVzaMTurACmggKDdIA2jB
JMiAiDCC/5r0RBXmSFsGmqP4Z4DG5xxe3dx+whShZN0FR7X1phx7F1x4A/2d
dWt082yM7/S1ZVBado7yrlCgp5RU3I8Lc8ns4SmfxfIhO6kMQIs3vlBZawm2
Bo6OpVRdD3KZ+2/d53MBTsAepGodW+v/B8TAwjrN01M//F0Ebaormt667byx
AeAMd+TL7JA7tXsUT0CbdiLOaJcZuFWXPHehgGGVUnXM502SpPnr+c2JXJbD
nykWmSvnMdWN4MjnZUfGQIVkHh9RNVFMlpjoJt+YpuTpZTsSlXUfxZ3o2Eqv
dLi4fxDh05IM5Xh5OcGotHv4hRf1St5XnQhpkDEHl02u9lYkBXCSNdyc2+dT
848AXn4f0PQwIsPf1bZRLf4fRvQ5O16DoevJDER2P3vXu2ez6Nv8YLrcReLU
H3Ttf98abGR0G+q+aklE4SvIi+81pDS84N9Lr2h8fYBFDGNKCEtoVKLCl7gx
S+QOVrrzKCKAl0E/XnfqSUffls3ZjEwD10pRIfM0Ehi/VfcxU8VqahNo13/g
YgZvYa7qdxobBH5p+CFgN7UK0vrtHjEjSmxmGi5Vx1L3q1p6jySGEQIoOoAL
6cd5wI0ssu56CHWaotdXCoIfn+7UzQYsK6IBXKgrbz7c0c1/paAS4oVUkDfV
zqwEuyw3PFd/mkOC6tB2433cpc8gUyhqpeyMjKe9Dbi+TYgsHowzaVlLSLMZ
LHU7/oztbMTBg9IGnMVH/Fqgc00HG2xMT0L5ukWyxvhdyTSorC6o9oJYV6xe
KKj/2IyE8vHu6zKLgRSjF1k5aPvZOd7e/6sgORAcqqpr4CfxV2pwpbGpy9Yi
A12qWHCO9wTgoG8M53ZTMdVU4Csx4a4PofieEmzfytYEh7f8y7DO9kCExIZb
SnPGyvZLQkOPzQg62iKs7Del0P+cHtvsSxSk0RNw/0QOq9JewBb1wM4eZmpP
RWLfnqt3VQxwSI0NNaZEhHyRFkZNWSARvFD3sij0ii9gZ3nTLoXVTG62CEqd
RHjna0X4y1LgS2VoXXQ0cK/bYjJjlkA7Z+kSiettxC5RUJMfFw47GPkFime3
1Vv4CxV0c48QQtWYvWhRUVkLy2I8GZwOXqM2uj0xNgke8yO2ayDpqGJUumed
kmBk21t6M3JEX1mmi1dzmkz/liP/Enw5TC0KNe4wCoFjV5p1Uh5P/+QwYY/r
pUqQtgnV+ihFgmJm75Wt+al4v7H3IECznEO0LbnAKV9CDGjtE+/RbU0xf/KD
cxsgYPp9NXXS/leRDtSMn9IO0BRfwltJkDmSg0NXoQzaQXze7NbynC1Bzywg
9Cnk29duMIXMdVzQglMJ+yajZGM3R2+m30CvzWAq/VwvuHXtW7jcUBCAIUpp
Ugh0TDwp2gPG3RXQvRx9sGvbKj9V3L7Zv7Ib2hzQBjgheCDH6DrJO4sFXlEP
rDctCYtO/5bTIfeyfjsqA9dQTguQMtlKvH0NLSF5ngvxbUGWXzNWgdfLPfJ+
aZtGHejbChDgrHIygR9TJcIdfW6HxrgtqlIajl8AhZ6A2uQymeS7PAR55pKH
nqzm9cchBDv6lES3U5esq3q/+LKpg7JJHjH7y+brHIfuiNz7bchPnPyOcrcX
vfvwbd65++MuEiFoJhblubp7tGxk1itPtJdZBWeLkqBLz0GLldWxFZE6MTXO
IiWQX8SzyFguz7p4v9FqjCQO93Lj41AI75H/jjpI6kxFLfxtdDFkNZGFS7Hq
3ECuVm98M7mGe/2/QypkBdHOCvwpLu5GuISHGv4g/ybBFR/fvQVmgvkVi5rR
L1AX/vinBWXVpApC1/HxnaLj3sRtBptAQUMegu/+m4jLIpIlMCMoV2lxqEYx
NAJfb5wuurQlvzwMEyTk+N9A2IlgX+cIUZWADQRvTPKh9181zwepjv1yf/+2
4fL/NJajezTWj2kskkdL70JrPi0tSEfnWg+wqHKw2i4eldPvHEba/z185h3m
jFjVlHZoUb7T5AqHVv8ZrRbKWTEA/+pcJmOPjXHBe773paClVpXgvI/yZ84v
P4CbeZSCmFihQw1q9RdOd0EpZx3hPz4XWj54rMpnqCuHv7DHEyppkWpOItmP
RDjrmQU5fd9J7y12T5dRkKGSNT6RNUGNoutvdfax4fp/0EnS3nViklEwbYfL
P92PdHUT+Bv11YrYYe2ahgN9PDepn53m+8dIKx6eCRfHTTROeUJK9zS9hDFu
UpkpNd9N0j9MPr/V+Vbmq5W0NqfVFDVW5uzfoxXsw4plhjx0dkI1baMX5RhS
rIb/D8LdTsMRjeWV2gH9qYK1aGd29wlxDLROhQ37Jnwl35sYajFkiFT9nSyK
deECH6jBzY6Nd3PhuEoHIwb7qa990LXibhRmtceP0Ug1KOYLn6XXKOjR+/cx
C0jUAr1IZzT3+gMaeXa3Vm29jBKvHDfFCNRSXPgRIAxHnB+CS8N09x7b2D1e
iI/4zLrhj8gIQ2d6INKRKrFKoAa+ksX6EqRqe0A+g9CHyyrP5VMBtOcHKXVD
cVlJ8fgmqPm/O5Vukxt9CfUhL9YsTiE5IKXXKZpDRV8sQXj6Whnpl8pilOYO
dc0yhRja4hmPhhCOEmIASepgqZV2CqETF9ml4+klLXwC5h//xYRE5apZTBnh
SzNPyYaRhxz0XQCk4syuIlPRAG/ufNU18mcTTYS+f96NM3vt55dNWEq7ALcZ
xvmYGfDaTFQ6awkzX3SGAioq4M0gOK0cACh3eePcsA6e3hhYAYQVfA0pi054
fHV3X2jRVYka4BztDpr6RB/klfnaFA8UFLjPns4cqOFhqgem5iaKa9VeMioQ
k6lKZI7Xx/nLXBQ6QXZB+/wfMVV9J0eI7dMig6Z+/Gf/4fM+p9RDXtWiTM8v
NBPN2Fwix6njl3rfWf5xlja9hmxU7CZrv9gC2GlD755rMUlpl4iWb6XhtGNL
qDs0FyC1S/iGjaW8vtf/jQQqbbhBCEIYeSC89rq2E/jNBHxo8qudZI3zp8Em
NYavwpb8SU/6+HMzLemPcNLgDJAsVi6OoSOxk6jH8NVv28UF6UqmwN59zC6G
72/SEovPg/CsBTcWMnic3K2WEKK3cUX5S8jNFo1sEW3argOlZxR0dYBfK3wC
0rifzg/1orEZ7Kb/H2aYxSx96xCMEvXhEDUelg1sdETuHPnxcls18aAErHLO
NqwymDw7LXUzZJyvHEPB+yREcUa9dhnuzz4G1DIOYwi9bG678jw8quVfYQqt
v5JCV6OlLdrp5Z+a+yDTn/3IlU3fwpnB4+O3qeLW2K5opXXl93RtTw03ZGoQ
Y8zCDJXR8V2iBFuKOAH4ua8+ILwp1MECq6Yg1TGihzV2Rh2ykJFTWmhhd1EA
28cmQnc5y58kr6nh1NQMz+6r+vvlPzNoyg2yFF41TEcvG08w1f83rGnZqnUb
bZ0iJRHYL3PsY06ulQdzYi72vv9l58ShVNnzQEsAq/IYLbuPs9vXugSARxtw
eE5F4UMKwfQwDu5xGQid/OolLZKxU5ABGb7BxgtiAiXtkJ81qMvfrHUVKY7h
kTtTVBlrhLPTlakofOlALVQVXgYJZkH6Dz8bGj6KkD34YmJ5mWYJiqQhLF2N
OimG2PMCvF1XfpDX8tV37T01L1IIqJbOgMHohvQRihY5rh9PuSWkBWUJUTxS
2LW7cTpsv2kMpotb4aGiTQMZ6luZBpDrHOEw4uvPqSCsZfKJwLKgw4pjcZly
7bDhWuPzXyY0a0PtQ4TYX+I6q4UGirIn/FeDz2wxFF6BS6Z6rGIrr6sGoT+c
jvK7GzSIfz607zpkBwfH8r5sYK7AIU10aFqTYdLtGjjGGWEJw0VIgOehTRTy
+vxvzgyRhZc/thCdh7zgelphIJYDTcwI7+NIosftD+V0f2YMR7dejjMEOXA5
ZdxglmcTG8ssC67ZEy960q9eA0bPM/OVrNPQr/bNjiTVlYBtyDkuTal7DeDe
NjCRDKVWeqDWfikgTpo65SBUksA2x+JCDxqXgWDXvnGa5j/AYqydNmc8Z6jQ
A85THkiplXjm8Mp9kXbDXxgj6roNar4cmx5P8z1l4c7Q6xvxI8ZpnKyf95k+
al0weAuCC54b5zRS+IutvKEeJzpTKYjTzijfYfzK9io0Bmf5+etBk4nnUGkR
RGuT/0iOVFrQdf0RS98cBoXxzcnBNNP1KepL9f05ny7H18Cblp6ifbd7XnM6
CGHbwH7VXt/W9teEig2xw4Cv1gJOsHSXiMDbG7ao3a/s4RghmS3e0oAi/ZQv
6J5qpVgIgmGDnsKs2lwsjMSY74gxPGD4x2HH/1jaQlwp26sNb0xfCIXsui2f
jZZxwkGuXapr/nG9OLIxdM+1shsBgJNfIWSCSzN/+hi+TlABnVItT84oQwnJ
vpXNy9GvPA5R5UepKxy0UNgMRM66qnsPxtz5t+EhB90Mrw+Kr41ghpfQ3fid
qVg/vp5Q/webBRmNhUFb0TQiLOz00DepcbfbwMsgGyZBvqfX38pqHpCspbfR
YokKRptJDkPtMrRjFp2MjzAqHdnDKOhlZ+urxYtLIYgPQj6MMFn+1u8H3+GK
xE1QcuHLUDk3LC7TzS2EhJHIGD3GPx0iUH5y9ZRpKFWDWuXE3a6wplx3Emqs
l28la0d6Ei/cwP9yQ83SeZWzvAOrA0y9oEIcpM2TK0uogrKer58NB9r3AoGQ
bCErDy/WYQhqnszqklm69I25ZRK4UeTziwUtBE1J1zWPj9Yh9SdOwEe1kJKU
p7vqsfmG61mHAKxF1jn9iS7iTNJrm6VV4POYwqDwPvgO/ChjVzUXp0ViACrB
xTvOzLQ169DYdhheUUWYvjZOi7eRVG+jUAVDsn0KeFgK8ttI4RszAfqpAmDr
4Mp0xQWQqf8xVTdhnpmeZAaW3WWgL3p+1vCG06c1euIwsa+7xq6ZpfoYG6Cf
ajWX897QZVdsHEQvgC3h1pXykYxv1YpNgiLP+tpg6U6FrUW14VTcOAmBIgh+
y4dKdaBljTfKNC2LvPrhBOmLvHAxdWoLb1jwQuHJOFHZTMgDtGpT0MxDq31V
KXdF1zsFy9jwaEc2FmyX9sfwHv04ElyXUtQ2gT4xyFR6g9BRG4KitowynyRi
mlHmUkqqXBzJv3teAaxBs1wRdbb1C7A+4exp+/qL1pxYrPUIlvG2DQJ/1Fa2
f9rMGSXsrkuXMl8JitHMcK1bFKbfpoPZlQd1Hf7NBjYKO/+ZNPI77Bx4sfIm
NIJfbBvh2UQqjlv6kCcEt/1AIZLNEbKD5/Zv307LpFriUcuo7djtRt8r9jyK
IUpfiE9rMGDjjkRkfHG614m2WSiQ4fqikgUVyExUk9zb4Sm1BRoMoEy0vM61
HW4ovF2IbuZR/L+VO/uGtnJLDeU43akohFHVYWOOdL6WiOjP+26GNfaqaO5M
sOEk6nAZGrw8LC5OyOrOMI6XQHID/Q7fg/oU+tJVffMElf9j593ckrR+nluC
H7zZLT6PoOicKyA4ptpvaHEkrij9APwTjAoS67tVt8viYP8Zz13XnfyQ5ubM
265WuyKUVf/erlQ/Kj886wER5if5dtzI59fgDl/WrsmaQw4iMWsAACL0hX4b
PWFsX+G1ojZcJBKovYj+BT3CT1aacevprIuhDu2K/fuuX59E4+P6DMdpd5Mp
LRz6DTT62K5We/T3z2AnBQmddvVAeoGXa9K7DUGBM7bhmk41g/oPYeb8sHnm
QZlj8PQZ9IH0uRGNa5wg1oKNFYC5r60tMdfEWX1c3Wj0hJL0EO9b6I2k93di
ohv9I4o6HhytFOW/wpBzcQCfo94z+ZGjj7oGkylrOqbydREv7t2shti6+0GD
ipQELPJPrS3l+QIAjn2M8bxzK25PhVqceC0DMwlaCpYi3XSsXP3cvhp3iVhU
2z6rfEGSa5Kk31c5v1O43aveY7mG3DB+WE8J13cpDeQUC+P+Jl4DvfF7HwNF
0yQR28QW728oG9lRvfXEQrykSAbZyRihEwnn/7DUVT9jO5jU2EuNaki5TVgk
TY/4n6zik87TDLufg4ZuHYlOcuYwfSC0yEvx/YV/J3K+9djSWEYHxtdqPNjx
dFynCUmYf6LM3+fA4Yoi8ilcxbeJxY5b75EOZHp2EPs8GsnwZbpwx9Z0ie1Q
Cjxzj408Rf2naSvpdZcBkCnDBbAsPKT1BZh4t2Uqf7MWnSo6TgEKpHwRTjxy
62M+hG2fpKF7npJYv9gILnH7O9sXFRiN3ci7RUUJ06nCPkY9/maljKWi3fhI
Eaz657rRdqLLe9Imwq22brRoedwsz1frIuAQNvtW94gtJvfenZJSEuaRbhW4
3B2DpOkv1vZYIJIBT/h36fQI7vegixLK6P5PMXKCjjFj5sS2qgQqVIiv4bKY
NogXTS8uXP5LUdBdUi8+DD0Sd2hLviYlbBmHnYlmJecdwtVIFkd6e5h+Ivyk
47t6SqwtDvSnMSCYVXjgWln+107+I7ENw6UuJPZ9EXEnSa0pmf+P1d9fOyi5
sDuLOWCw/kSRPyA9LInUc1OnkryfvelXZbaRSSBzc2DYvzuyS00rV3ME3XAs
Z6ELBt9GW7ntN7UU0auPJNGCMWNjzOWWRmcy5UEgdGHzY8Ljn8VHK2c0tlz0
N8P2sQOdk6weGPYcgXETvsp+Q3MF7kfuHW9hTLYu0b8rmYLyHEz5Tkgxy7GP
cOPZNETeXTv93iyMjZNtooBcKn/3BPavxt0iXx+f+uBUCdJoH24mkfWTGZzJ
0WIABbpnXOEdXv6gd7QRBzN/bIuU6B7xsDoaY+QxwME0jhMarobaLztgq6Ez
SoinvFlVFIJjVgDuZFbgKXOF9Mv+jp47QjO5WQEA96wzxVHEsXkRR3x5kEg6
EOLvTzROjNffzW1l1x03VLK4SvblgiqPP6WZqWQWHAQkVP1dnuUEnTuVO/K6
fertYs1n/vf3hbWrptMQIznVyv3MnSBspRK3sFT+5xtLanHeuMcYWqGTWhDR
zPSZ3v+LXG5mT/poALxsvrYt10gPsELRiaYG4BTydqaQSNXIbkCeZke5M3JV
Kb74JVM38E/TlvQriiijcZenN0RoswsEttXkOnjmS5ym068EzcaKpEfHn8C1
RE6y934SAIOr31k8nuDZsKdw3bXTByelPVFRyUfghhr2fKAWsXjQQjMjziYF
RXuJl8C8fzpz6jqGY0Fy/UigqDVvTrrp8BaXlBHiWYZTOoO1xs71XfOLYIoH
D0kZPYu8ukBQ6UoH2g5tjZsNkkvhJuLCXoDALOJo8NODC906rfkD55HPlCLO
OeZqdjM2enqYoLX4h8U/TASTFrUtK2FnIf/Np30sCfrbFWcbeB+OskYjFG+p
oIf9L05GWJB5OC/8sTCbPzyZFmKH3hix8DPPOQOkzcQqHpP4Lm1HduzbN8cR
hLtNKoNlkLyvhrWNrD8ob8utkNde736DLCoR945+uWjhI4SXabp0ieogeDCA
XCmLIu9vI1PR/yjLL3E3pzJo6Mp0YRUSEidFUFuzeQh6b89E/+mLFcd+YDhK
9FrfPaGYmTX85x8WF9h1nBfrNXwPlu2acrDh+hrhe7vGRbTF4PF9xegTWi7P
PrzJ+WT1HGuXDdcuWdIKnWfLDSQDElR3W0TX3ikd+SH5rbXR9Ds+rHINk53G
+yy419W1Gm+loGWrMNXJ9gAcgWhBg2rxH7m3Wr7IoM2vc9JUIgjeYr3yHvXN
ZkvdvMIH9JoTFpp8yfCEsS6dMwJeXR1UZcMfVjBS69pFnWxE0l47odmkM9J6
XGA3ZcfphFQvRXOZar2DSpSTK8Oa0p1P34tgIQm9uvnp329Kb3jTwPbAb97a
2woQFyzyeRByVm170kFA92VaZAcQ5i6pERw7O7FxnujtLrp8vBTCt7Ob38U3
hDC55nCVe4aOsHaOic10Y7jN3PEDUtXu0QM5DUFHz6nLXDs2S+AI1bz+2sf8
1NyGGq3K+BOErlqHJDJeobM3K/DUwiFRC3eotxW1tQ0vmvNaHvGH4gM25sWc
L6wcKswIts1JgEqbb1UUohibTTrKzoah75E4/OILaOcrqJ4omX9L2YnX32P2
FHABC2q65bPajs7jq/IRH8aAcO7XESxuUIv31EIXWK5BcMRN/yFaXgkNSShP
76Dt7Lv7i2AX3Ebk7LF46N2N/O+eMIviuSGspj+AAgXLDRF2SgIXbRIDev/E
Yc2VRb66gTFkGTU1H1WdLJy0BbYIlcx8uRNpuAK9o+WN3axeHVtSQE2k9VZq
aJpNYwOVoUdy6tjJc+OXZkBvrqmt66q+gB2lhnh8BsizSpWzRuiTdn6tI8Vt
eridbjELNSFVvPZit9hCwLfgmT9EloKtKrUU1C6QOJUqFs/PeI48zVtqN+WU
MfbMZ0+/rL0aX3Sh4jVq6XsIrFAsS/pNcd7r6z2d9KycGWvCZiIjHosDlj3o
3MCTWUvtW+omgi/vwE2ar+c72qUm2m5A0eLcio+78EAqeU8sV1iajzK5iGHv
Qyhj4EcaMRx3nRIoit2LkSc1z668K+1DCEY1m0q1Y0iEwnSbEfKtsQFUr4uh
x3bmPxpInayRdqeryKHZNDz8HKC+4TYFtdGRSVCZBopx17u7hytfLdoT2jpn
v21vjReeV1Liz6ynVtcqItKscxxqsId7k/WP8Px0NwDbGwW7iALG6NekDOUN
rwaxrqtVL+Git2Z81OZ4r+YlOcsQSfG1MfaI6g4r/Ch/iR5zYjRFBQ4VsWWq
99Nqm3yq7xECZIlo027th+LEKx700q7xrP0gI/rdSA5J+z/W8inheEMsYLBP
wQ/HMdmvWN2gCl5eTwq/GgKAxSH1459o69zZ7TbVp8d0rz3QU//+ZayiLVp0
nH/CikCTAQvGQyvJMUJ6HWe/Ia04W6O+mDa3a+GAjBm0xbKLiNN8Xiv5TLTE
rQ1qGCvZ1YRCY//7ZHmSp5mmwTtXlkzOa/AeydV1iM9xyPIsMPOw5t+dsfVo
BvohnBfbi/oLwY7pnhjBjJduNl9vSCrXx5AiGDrU9EofQsFYSeIjWEhfuZ7I
/JRUYKU8GPTDOl1jQjOVxRCfDrclU09qROSs5GPKP8+xNVETdvBFuapLybhq
3yCSV3EB1g2fIcQvCKmyWYjuCaDP0uxaXnHr5Hsm2BZaI8FyR3K8pPKbarnc
xUfeIRiwTqKsTMubsoftJsubt8YRkYXWGnZajYa+XuQiRk9ji33mVBX6x+Ra
uoX00QiPEhfqIxbeINPwL0cqk1fTV5PAUerxpBxpc5QVBFGeElsuurBFjWlc
FDya+J++yR0ntLjnOcFn0SiSmt14ErKVjYSQBInNQg3Rnr3ZtaDYEEyq8ECm
UmWGvht8S29Pn1fyT7puXksEuzs6VH/fINvRLaOniqeb6dCkJP9P0iwMHVUr
xp4M7YFljuB6JIZZT1svWb30ndkqzEI58iSnawYJF0uXrDxiGvZ8yCmCPCYR
7eLv2d5YD1AKoztLta1EMEJ9CkR6GoauXP9i2BjLfbrQX7q77ZoA85qn4kKx
IywpS/wNzAgSy8ZXJYdxJUt54LoVF7mENUj49knP3RqMbaZSbuKzkOemBuGl
fp58+xuLnejVKFwY6ovM1W8VVDBdkEqHd0wiX5s6jzIiUVUM5uQGNtNpRhzA
HZ1+4Rfy6dQhjmb2CyPdkK/9O38dpNV60gSAwj5BRlSHj0w8bvLB9zgv1XLe
XWNE3QyGdXnFD+4puh6z9p2UVe7mJkRuzweopaOEGI36iSmRr2uKNZluzU9I
NAS37nj2mBvuTaiSzSqW5YY3ZUHdTnFhPIA1jrD10PpGRRG53tkMEsvksSe8
JQyCAV2lSBMVx2jbkGxYcfcmQcarmurD94N7tYljbmE02HFzV50MG5lDv/6y
ATrGfYpIDZfkRItwasIU3tLfuj9Fg2p/MYWB+ZyzWW+bXOgocUZlhMcccTS8
wVCK5V4X6mykJuuaOZ6LNtC1Uu6gGgjnGzFHPdKlPqitfweIjvQMx8GFKAlM
0hiliimG2W2/QijolJby8y4a5dkQIL5fDxDe6S/hDUTeANTvBmjmiMeG03Bc
DkQz9Amii9m471T4g6J4nrHVW1tnsHg094ty2UfoUVZqbxEwTowtbCfwJewf
d9fohzaShv7UVUshy/P7f6/85oWM0SAvYteaHz71tE0pUkxc9S8gCiJp4hmd
3s9veHkAM+sw3AOfCgiQnLhKcI5jp/CTKPgd2IHmwG+PO9YyO3uHz3T76xiJ
whb5o/FbQZWY4dJXGhmkVr+C7oVJDRVByYucv4DvR6E5fjzS9ogy33ZUzRdt
we7NMsLb8pYEQKDKCij7a27y7vMa3FeWqVMyRUxk1ZQQL0K3FMjAucfTCvGY
HTuuLUDhAvY8WkKTFCyGm2Ty0dpBnceFQiugi6n+Ks/wdN6bPBmS/FX2XMkj
DwQs5FiQkkAFci5ZhnE99tOa88of3XYo5sWRrZ7zTtxsi+hm+qh2I0au4OxB
xZGy+dyxLs/VGPjqsjo6219ahl8bUv+qxA9kiMxaiWhv9qkuHdlnzysHA/ZP
NKLG8ZJDhLChWM7Y9GsLr+szJ1x7LKfUMK3tmwIZrmadnzW+EEr6UKjCbtyR
tF8gu/amIddDiHU2PpHBSLAmAPlb62GYUPTWTeBO12KbNl7lfupr6hjKoB9Z
jsSDKFKGOlLG8UZ5QzgRK+BSf5tgWhWobc9bJ9CMXWCQ3gAotlHoiAw5Xdj5
pb5h9O5U3hWh0nCDHD088v4FcPP6QwRxgFrlRIdderNEVhRnegciTSWCap6x
jHf8r2b/AM1ByXkQi15YYkZgXQumcIXEvsYFF3kBVGSLpyW9TZn/TOfVtoxG
xrU0fjXgPPqXbSCxuNmqqgejhNLr17SNnvUAFV6Nj3c0hbJDHI1tuIEjSB7F
t+aDmpBF/Fx1/zCIVED1+JuV+xaR5SoudrTn+CVIWHDJmTO3ZYawKbX9EiOA
ARZGr6FOSs2FEfZQMsdLy02CTXQ7hhoGvsxpzMyPLEJfInkxqLgTcrOAKVCz
NhOn8m0OJZIAnt6H7VYiT3YfjtwIZG77uXvJgeC6+gNZO+RElriZz7Vk7IKg
/lPZY7KkaUFt0hNbrscur5U+/yix+ChmpxWBK6FOfZHDuJy82f7eHHe9StPn
LFRsPV8hRoz52U9XKMwLGfWP48MDq/W/NcB+f1K1xSzUHUc8CTOhZgW6P5XJ
bYGf7o0zRbaGWenxbtwfBUee7ENEgHPeTxnzLRCnj2XQyCwyJkkcHHWXJmox
DiV4fgbSpXhqQazvJcpo1+pg8u1gUfY7qbE0VPWETxCkzPcebByvqCrZsxxD
4WdQGMdv7UzonvamXdsgvWtdCGDy/VPi42t1SwhC2Sjfx3B3yacLfIFJqfjW
8eLGmTESm0mXd7PHcqsyu/7JkwqJ52v+rJCwJx2Op4eWx++EyXm5U5eqUGZ8
aPFSirk3riLhJl4eLP9Br/6oWhG1VIwi33bx3391IgnaZ2qeg0bSRALkYHX1
VYJMWodqsdyhjiNCvvoytBw3HUxOCbwNrZExLJQpxd9CWasvaqge5Dl7zrNZ
oKCrFW28uoZOmK8dZ08nAVbjbe6zC55OkD+xPhuwyscthN7NNtSvkYgEf9Gt
0Necaoe+Lw+3dXUXvGfeAm90gvCGH/yECYoqtDZ61d1oIGQvx0W8tZsUX8YG
wQYGeBJzkUS3UhZdwggETCQ0U3mfYFAkS1Sbw7zHVM76KG4mvlvRGo3PT0LL
yAI72IZt2dYUpGs6RV6X5q9D9r7AeVQHCRor9b/FDIOnAj7ouaAzUqtbBXQa
Fekr0bWDE0khQSgI7MpwmApP69XdOY7EEAB38zhNW9dCTVEJz2QaiKSd6yQg
4wcUgWEI2DLzCVpc8f+0oRp8oURdGtk0DIGxurXos4aI1X6rOGq57Mzhf/xy
y+nO1459sETc1TQONNZALOsqouNAMtJmzF1zor+qKphW6DpJQE7fvFf3fm++
YHFGKxuYwmGa9f9sPw11ULkPDO81S6M4j50mLUm27kL3B3HGMMFFr60cHNRj
B3xF6LJp+jRCIAaEkv2TGiD0/fFHBaB24HzBXxICgOxvMMdnXBS3P9vjoyyp
87ppxGRrkdCbBWjnXqdgJxuQGyV/SZADQv8z/DcvXFGDA/AhFEWCiuXBrX7F
G1ulduqlBSvwT9z5YiiNMRDQD+6ILxB6VfsN2JxbsBQziG2z/cZ/qTCT7Hwe
9iAoPyXpntzjOLN7xy9PAtm7UTQ/X9vJsLLA8l5gWXmRmVXdw41qeiyxzUft
TqrvK7S0XqGijQPzzSVt+n2G71X8U09/2vvT/+dt4raasB0myFDawD7tKUaP
maWh4IMNYVWjzFXh8yqGWkIr0X9kQYqndcPi/fqu37lIyV0zm1s9RfiCBsDb
UgX9lcCAVx73jasDG7iVAGL5d5pbSJQ+wDpEIHN22jdw46pcn7lO6VjU+g9R
0Hrvi3TWgnkD6COcTOUduDjdiMrNTDfFFogIphaAnbSP27BJGYxuLTrvv5kC
OmcSFOMFaKmEsT9xcyd26apzDMlRgKheWNUaGl0clu0D5VICloIMVnp3Zz01
Low+mo/qQZvmk8SFL4hMQ0imU3Bupp6sMZJpzM40iW37b66lmvCp9SyQy0sM
X7uV1Hr18NvgIv7IDRgeNQDPTWU/bDdCaqWqKod2iKHlWTCArayuGJHnG+EI
tsDhv7PmkKRgx0zyyQD2Z0pf53evD/8mx/mZPy2gKN18+ehRigIID1xLbxI+
i1ePtxDLq72LpRRLZC2WAgpuR/NalI2RN2Siyg+xH7uACiZmQxD0Urq1XByZ
6oA+729YsOnoW3P0Sx7u31tm2qwDo5aXmoDtFnMJxMeioXlPK2TEZz+Q0nBD
6atnJxMOdnS29VyvJ2BrZfrBy6YkM2tcSzJrCDBchgCupEjB2rLqqsH3a6m3
ALAyifmes19WVXqXZd4cjD3YXz3dWP1bobtTnyXYee+ZjxiiE2FRbU+vxBVe
zyyJwiiyNk+DF1x6KB6BxwpFfDUqc0tKdP9Uo3ybdvVCunWmqr/bCGbV1LOe
3RFW1TpMwKRHFyfpqlfl+WiiXUkMzLCSh0YR9VZRNTqNSaJrzPLVlXQd/c18
R3KJHBOIgJKRESnCMstjXtGUkifKGIBfqekLSBCnhXkyZzlQ6Xkuz8F3nBSz
QO0XLoa9P1BzpoLSB8n3OVM1TCeFvokkbVQKdrwRCGNxLAkQOkl6a8jXnKar
n2d6HqUDdKeJQakTF8yKNzD661rW4fPetSgEXS0XeG6JFP1FKlTQffNeOI2O
i3T9FgwP0Gwsj8QHAu7CqKoS1rMHl8NVbhG8jfHkTEyXArkj9MoOTCyqsSVT
Rnap1HP2FezKx6LdDt6OKfN4Ez3xuDUMJppKcvaOP1iBoLIdByrZbJf2ThBK
ZOE9MqQ8vU+Pvks+X5PMc30RZW2nCP7z5iisYsC5AI+u2q+1Rb8ygECd2Z6G
BscYwLypJ3GMZso2Ea24H7EjDArI3h0DnWNo7mG8B5sMWCswqlnPyGVusRy2
NZWnndywlqlbHuUSYyp5+CGzGxXn8Q7B4wtRt4P7Zm2jE06Ebst3xKgMx0/w
wU8X9GocHWo3YPiLwtNr3sbSybcBHSAoRpOOqc/i2KbZqiRFrFwF1qv8SpIw
XZr+9S761/z42/4zAPOiNJd4Jcot7hFhPBejwk+bgG3GulT+eBQmlv/fbGco
Oj1Xs0nNnUTfUM2N+4UC93l8UZwxvpYXIYSSxejouAiLRwZjLeGUgBfAQXbl
/cXCkA3ibkbAWiunS+JNdxEO2RnoQmMQVaTR8JW8KxNlC4NSHqpWoAgMXc9B
60yE09PBjMp8/NOdWK+MiaBISjf1WwDkPdI1+DeNsF+7jbTCv2fnGt9esQST
nOGFK3jcPQtLISrJ487R+f1gLj03IxtiFNe+cRqKEurOUgOkV1uCFBG8cqOl
m5JqI8PGn692tzjc8xKCjj1FDt+qgOdNwQ45eHJsybHR5shp6ov94Hal7Tvc
cv6GgU2Lk7fXeg1yHCm0DXPcHhBOBOVVDwKLM3ZX4qcxHmAwTKLOPQF7EGij
/hXZat956VVmEK6GrzKSY15hBOzcPKpKdycy74cLRMttrqhquP5l/NdMvB+1
DjxlxGBMgtT3f3WR2qMSnIQSOBYqXloeQjD1jn98cNd4KjL7qp6O40/LsHTl
HE0Yxw+HA4KY9cq3ZFQVvIytugAHbYejRHgyxjToyoWRRlZx6QuGgjwzmc3c
bDRc/YEp0MCuSuCRbJz/bpg5I6SGWuqDhk11cb3xTqwWmRRjw538R3Mf2rB1
IPr24NsVcYjWsih7NBRmNamB/8ZPnbgW27u6jEbXOvUZNYklnJLIYxWl84CB
rF9eWUQcffmPRiqaHwshVGFJPPVZsS2vMIULiNPDFYskU6NP76pmmE3V16Gr
kyGycOIlS3TPldWJZZFzoPkXr22Dih/FYJ3l+o21GdmMds+CHDewhuUnISWO
oddQXMdzf+hOJqopSpxJMW+H2AuwQLyu4MYytkYbMnZfd8WXba+UtLx0ynhf
h3yquvDsf8nPob0IaHNMBq878e7zDcGT6ltLu2ktG2oSlqlC+AEByUcSNpnb
uV2JNZvQO1yF46QZT22X37wuPmSlr76b/8YMcDzVvENdqGT1biANDmdviM1X
lJL2uTfsLYb8rE84JTJ9DfJ642xpFLE7Tn5FfU6+kldWPxNJiOMoZUSqkaZa
oFpK+lp3GNEbJNqJfqgG/raN6UeHSjoDcOmVQp1oArUcxo7oik0F717Hafm6
qNRHlLYHJ2WQJS04Ir0KxjMdPPwEyz/EZlZbw7ZLjy03K3GGn7u4oY+nZUYf
jgXEVQgxd7xDP7sBppK1GwFUc6UBT3Nhx+xJ6acwfIiUUfN0Je/2FXt+oFsu
XDP2Z4oSppqa2/Ufvhvd2hyVBKBwggGjcxQRo9grTdjor7Cz5s2qAg96hCqU
qI01+uwU0fMMlAo+6Gkb02bS2epO26PAQHpkrycwGvxf0BoFNPMLwJV0vbPk
luZCg+bhd6QP28ry59RGlWmLH2+vBSfDQ5xg2nyQT2ESr24nJNvpElhu4hSP
qGhoyAnrhJKMNL10uhTGls108IRa/Tx+OuNQtXJlr8dDdmbmA5Z8cICHeRwm
3gWyafNVL0IjQG6uoHFcnDNZgkEMrFpxyHP15FjiaAhesFIWR2DPgapSsaXc
ZPsA4Risdw/FlqXcwqIzE8uzdJAqVxg0PB7M/SxsCUYgFwXBJgmzX+De8Hwj
49qfkWO3IHrmhoh2VliB4r148V1we/X7rr4KNFrn2oCUn4RrcAp6pPInq5lE
IyCL2CRyEfsFCtpADRKMUZTJtkKoSTTj8j7Rv8/O4qDTbaU7jNdNYZeoG2dg
ymZLgei0vnzzvDr7N9wXuHEO0MSO6wP0Usb8DqOHSXd8lhDzLtOEcT/espkX
nRcukMtUE5xlZNqUX5D5OG5c7u+FIl7cpYqUvGCwPzanyisCR50zKKMID1UF
IIBDMIhaGipdGox39AGl86IAf7uKtbM3Qcj5JpldPTDvgog58vYLHudWv//v
gwkphx/oCCKWw9wza8rBSvT73l9Lp0P5NQjGOKpLYzjXwPqDHK+N+L+K/Uvi
FnX8QbCLcDWp1Q1yljU21S7gVsO69YeJu9UWxtkC3idCja/hn+9g+jcTwb8K
sKLOBtUzM5gqYJvGGearoPDcFDqMm1avAVP/xq35yHzMOG5+dkHlKUU0Rwwm
yg3wzweYH3lJT1q19jzW73WiAejeOjAaNWSeKrVRBIjXcPTQnPZmrIeE8kGz
odPKi7YKTudiB3w/r2rGf6ZO0smnlqt1eQ0dsOXFSXLU4uqToVlJFgvo03qc
8tMcTHR8iI+wmXr72EaADjr+03/9RKKqKo/uzLyknLZmrHTjHCmIgSLUE8jk
pjINshCeEuDJWrHpg9783BonVQr2fJkO9ekJ4T0W0qkk+O6CcxSPLL/VMARq
qgRQ51hRttGl8Jug+fgOtWLWtzvBkjiy3771CcikxhC7SODf6LHuFahYng5Q
c8umdlVk2axrLSM/dsNec101KylnScnbwTCRFrOVoMwAvEJQQ4QTeOgSXLeZ
dlmfc6ejYqBBmQmkZgEwDt06aHVhJx9WEbBmZqXnruJZvwwdL6F2hynWsway
bHFKFE2BfWLPH9t7Et0Pbp6TXWkCtMbAy4ak+xzY2c2QwFT5z7f7Aw8tyH8x
bkj/zo6bKUfm6Q/xvfL9uqq9P1lpRZbMvazjGhoLWIOxxIc0pyj7qXDo34W5
0O5BTMYtzDd4tG1ZsG4fi48Xp1W0xIb4U5vHHRJqvFMR5lGpTpiVxd2e39Bi
GII5T556qdK0je8QKj43dqm8s9XrEiDnx2qNgAepNPZ8dD19tS3dB1l6RQ0R
5dqKnVziZBse7dwpw1uUutvOFsxgD0lZeks1/+HtWtWJdB7vcE4EwNHjOtSF
nIfIUJK75TIsan21zgNwEEK/BRXaEwSYIXvK/B+NLjQJe+3xD0zghlyk7rGH
T3CsfPdEFNMUMkK8KgNai7dwlQO9jEsAOr5sZWFhjBqCcphNwhnOLAhkrhWV
jdbgkZhZx168XStJNltoLc+g2NsOoRtd7NramMrw96OGXWkbI8MnyoabdbA8
e7blQn3Kzq36HWYuxpqzqRMTnEm9OiVPx3aU4auxUlNXiyZDd7V2Trvg2l0P
hc8CID/JxjO4rlyFnv+NLYf4F5mRfoAdrDKxUOcWHnky5T1e01IOKbJMDqkN
VahncrdPRgFRMETDHJ4NGP8lcXi38R7e4ZLpqXw0ICs+J5b23foA3zZRzNCF
MIb69RLJbGLUS7Q3YcLlDWBVO46OVW80bAuu9ByVHKaoQ4fU7+yym0BbSmrc
ZZ/t3NwE+oDu7zY61DHctQg2K3uogodDu9KRyzEn4jjr0HZFriJ709WvR250
W39u7HcFwnp2YKaXCavsfe7xHmbzj+UkgdTYzUhSGOzFht6g6hD0sscQwFCb
Xq4vJn3bgb1YE3EmhAq3GFaaFeKHVonAGHucaseTWOKDkE35LokIXOHrd69Z
+FmSJ3yJ/n1Y4bVr+oZHPIDy6skyT+wgfmR49SE3pljUHQouSvHNiYS8L/9u
yIRiKlSXwkwc/o/Nn76x/WSNpgWgn40E6wIY7NE0d/8EUlfyv+qg2a5gWSof
KcgItxv/+HVpg4cOkE7qr3hIA5k97lCUJEXpqnkXhKs8XtT6F+Qau1os1XJN
5WBD999dWJ6w2QIsgdYxl8NRlAXJpZmfEkBYPEwKOBhGBeBWBEjWNKU5lJsy
y5T2N21BkAp5q9gbdqNBON4N8fEI+eHVWVc3grYjJoqP5+CIQCrh2yXOCa30
xg6SOrMiwox0SEYhFTPo00NpFVhlcjxfKvoJ5zIXN5Akjs2VCOX5x2VSpOi6
zQCU2W/kX/ttpp5MRjhfSsuWCT9lLMADTnns59aNv2P9cU8yfot1ODivWlWw
ShxlNxjsjfOyViofDdQdj05x2Gt/shCUCrAsufmOsOrQvUE4JT/gzDUxCBrr
Q3z0EM3iyYeuQCdGzpTf35Dsr4nJmt0y8wLfPhktAAhLTttcNc4ceqgejuoR
JvF0d690t29CxP7cOUvN/Q8HHpaAFiuJVHWg5TtxtBkpXo2QTtcri+JOokEP
3Nlt9Yto2o9VNz3IpQ/zSIuGCmEpMcgKu0POF4sn3ai1t53grSzn643IASAP
Nat3yTow2484EIS5Fq0LXTYdME8NJr8wD/hXvES+rFyg8MDSZZ7I3iR/uu/l
5Z6R2PG4N5WcgJYwqqgrxGX7aLyEcQ9GNl3YJeaLqKrG7L0Ljcx+pSHiFoPe
XrkKy5r3rSNdsqLhIeM016pPVkOizT6P66fDXvHnXhw8+bewHt1HY6WF28Ke
3GsKmNYj69beSU0rW8KxHwhFq4Goo/SeRv7+mGK6mEhPCnth4v7kTD4fUPIm
fDDdi3K42OGON0x1Q+oY0jP9hB5CfPayX2k3FdTZEiHvGEd/I1PpaFhwDaH4
lgNsyZiDn5ZOHBjNNkjp/6h70xCTRZqWADkvsnhb2oqIghkZf09+LidsyyIK
UO82+hP4IZqNeTGA4XzQG5oTsOxRNE1kayh8jXmo9KPztrnKYWIwJw/DKgwh
kHAcO1b5Y4wsMVb9VmPsPf9qc7EOf8cGD5ORtfbFq19LrlniTriqrmEZDoZD
kLkNyD/X5OVzhx4X1Op4S+V/YP7hhvEYkaDG3nGFG9sX37zEEsHXr8YVbd1n
szZG5DTnxkUjHJQ17LbV9+VYUZYtUqT1b3ckB1lqaavOJqcy3pxrUiFd62Q6
AHL+pmZvYWwpmMo/DqsaYb3CiVwv+DXo4XhgculKaDV74OiRt/JI0BGYbNcQ
VpGdyhYT6Lz65c1SDAhFxUSE2GVoygtqSkgjuXaR03/2LxeBGgAQMu3SvYBx
7PIClZXgCRksQSGHAKTaDeQLMnXlWpDF6JmGmBppA+oJFPIqHhUxQAIOW75k
/MomYQ4fPoqT77sXQ65sbo/J8mYQk931anZRo/hBzS289jE72IY2qJjS1j1z
cCBgAIxy3q9t5LQBoBD7t13bg/Xdz3meYHfg8a68W0V1lBRGfb3QfzSUEvDL
M8crCH2dh0cD9R7oUXfaw8ooervxeQ+P2pzDfYsJL+1k7U9co9Au6tJ3FrA3
rYmWBo8MB/OynUvOYNak9d1/s6xgMdTATllJTPTf/fbN/o7OsFUBp+NgMoxd
e5AnxK6vdI/6S0mWb01nTMlFUxoSmmIu4Kln64gkKaTQRZkm0bF+sKpmBbyP
YFm/L6RX4AWARsX9wyjKBxd8irSAS1PuTmqg7ITk0yM1AOvRL22ExtEq54EA
7b/6BLDK/vS3E4PoBzSazZ0lKgdq2w9NZxvVSsYI8XwmaExpEnMMBpKiilSy
YRlH7HUwV5T3fL5H3YvcR1ky/zuzhcpVdzVGbVFmEMYZPPK8PF6EVoX9S5Kv
GR00Yn1EKl0wsThgCT6YB0sCf/9w1OEJJUIVOvX+gqLpTHcLkj74TPDjF5N5
GZIgXbdLD5pVh74pbrVJGY/y4a9wylN0mJMkGZlmOYXhS89qsxT9QEj2Md2p
/SDkvzipvRKij4wb36sWRdCiRtAJVUY9/yaEMsLVU3lpSwaBrF4jZzSa6sBJ
4qyk/EJgawNQAVwXHcP3Y41SEFxWyKuqeDT1ThrxDlyyhhipWT0Foyz7vCI7
kpnJZ9mlG+sdsBnAXKbcTS5QykmNWCYZXll0zRzxv3akphrq6J71LlXqTmVh
4BlVOPxvjk7HEgO9YWfzt4e3mnWPjAIh+g5kVH7618L8qRgUgFqPFts2euau
DDkEH5xRZzaOb0q/+6i65JlElz86xrC1npw35waVaCSfRCfQXMg1999aalWM
otIZyCW/HyU75zNfBNQeA5sgADG+yGxRYzry/Ff3jT1862ig3fg6QQMvfRNj
zyM7gcGNEIdq7RwDIZXtGIagX2hngqK9ab0a979etNbSkAm9u9ndkPx9j3KR
ahOZcScbwU0f+pgSnGHCwbraJ2LM0T/yxgt50xrgbgRr+qZtOLj8s5OmiNve
E7Xc2XkglZnGgoVWtWzmmMnaoTPbuStaLy6VuEmcjSOJ3PSYDNx4d+E9p1ri
Uo5kp6o9tmJdBTwNsLPQoi+mff5f+eUY0QBbeQLshRg5KSt4HG45ACFZA+hN
WYbEW7YMiGHKV5O4FfMWAK9cc//TVAR7oJLrgBbw9FeihokJiX9Hl0CJQQVn
IIMzu69Q61dHRLPxz/Nr0UUaD0ruUBNbJNCMui9r262vrm/QQqacpmI0hFrJ
3fqvHEJTD6Ha/pgm87+t5MaNJj0Db8sTsCqESPSog4LPjocGXKXeIuoi3KQ6
54Cr42B/a7cwO8zXMYq8eXFcs2t7scVjlQgB0lUMeDs+3vbKQ8WPMlUMvC3/
fak/sJ/xmEemLrhhdyLOluvWmsdrjRZ7ouhugpQlhcESGp2qhQ5ZtpQTouQm
qaZ+P0zblIOG0cRX1hvulkrz9A7En58B5ilZ94QSx1AA0y1fnH7eO8A4XIhi
B50ZCMyOGRhoAljG1Ypsc/+A2oEI0eGIA3w8eW2ugDKbNNvvrdXDzIf1Dhei
lZV++dOP3AaBT8PqlRceBUUPF0+ZZR5F/g2JGqjburo7Y/8eQUg1Ap/gWc/t
84tsrCNyc0Mc/abQBqWdCmyG8XLnX6kPppVtgnm6+PHxDMBy7D8i8/ZC4Q/Q
m3tRkWmjUs0cHh0+e0RPH8rmbdfiQYeHFw2/VuRP0zuQgjJCYB9Mv6yC5qiO
FIsdAwkk0t+2XffzFs1Qss76st8+C0cUtUGp25VJVsYN6jYKO/etnDlcbZVz
S2G8tZzyg3AUmj2N8vpf+z+Ylr1dg5uRaStMsjCDsJYnxWS7ACeM49Ej4WSD
LSfOz2ZJW5E+RwQDOubCf0BSI/kRLbQsnQ7Np2cSpoZEu9siFJ+rPS3XMkj+
ykg9DrD2TiBQct6TeSVav8On64cAKmZ3DyO3pyeJwIDQsBnCQ5X1kBaCZyeG
sRXmIkNdKyRUeCRX33KIsmH7/dPiss1HGr4nWoLSqqZ9Li9knrjjM3mDlE09
sSedWvLxDhMnRCpq0tpCPnQq0aIoOp5pWbhbbRJEEwYxfxK1jw0Y0fR2xnXq
o7hz3nKKjo3ttfdwE0AAj8afX4ckwxZ1CBKaKaPOE6LAa8YdXN5Rd/I/ikzo
LvTM8dniPphai9ad6xzETI5Suv63EhHTGesHB8EsnKlQTIS/gc+iyeQRFS14
4DY2YXvw3gOfnEo/Z41Onil7H7lsOKkDmitlOPlUXzmymTK4XVxVJjoK1/he
bK0cWOqDFD0GOWSCAs95n9yDthc8FasJlBiGFd+cTNjGBcQyd6yJOD3ktb4X
2lrWvzd8/DSKkU36uzxCLEW+XrKqn81GdyOzGQQmztVPZ0oa317ZvSz7DYJz
Bv3dtlLeSAKTx9YnR401Xdc5SPoLtrP0ZozzDk+vDF0zo7CUNOe9ohw/xfLP
yY5DJN44YvTjCQ3R2OZ4woyeuGZ9uU2XmFIiUKprdWkKUGC48yMN0T8w0y7F
UZTkOcIpD2Mtzs73g7zwcfsnNxPyaVEFcXWyTiHmfYrrGuZwOOXDaplg3Uuk
9cdLnj9h5fFu72AdYuBokKQW3gWWbuiDXpDP7Tq0KKg3f09oQlEgY+7m6jCL
BvSwDNbuDmMz7fKnauga03I0TyxyZEbKLDHqmJVwJHZItOQtCO0HyfRZMrnr
fqly/Ajhudv4ExPyZaHHvsOyLSOynKRKxpQe9CCt66/NjRA4ow2C+fzy+Ag5
U/BF/z5wukYhZEtKWz9khtWon5NgPh4NVmR0S3Z+BnJ5c9u2WtANeFUNodVB
jPTO1IM5DGrC+Vq3FuItNSkXrhfB/VKa+nmVi01pXe/pamXS64o9mtMb57a3
uJtB/JmmWpo1Jvuuqfm/E9YnOcjjoSlH5JyMxt0wBjh5GOEljBBX/7ghbD1k
4jVkGOU3UV0HnglKjbNAZ8pgoTvRKOx0iDPpsLvr3Btclp/ehw2fbeK+XUkg
4rLa6rCD3H67qSg9kxws117dHqn2cFoKIHX+vsXAHNxoHFIRXbbpt1DsoylJ
leTpXCQgFCC249Qx1dlgk6B6rscBstb1Nj4ZNn78oG0zetyOfRfvqGcah2OZ
+F5QkWmn8Ig2A8afd0GjTzi1lQlvyfHwmpOkw43x8CFzh9IMLuVUuB5pjRH9
TeFuiVIKFmPksFRRMtfOMrvb9MVMXiz/cyhtlyNRYPQ4/RCQCWpKuC3rcDqj
wxqJ+Eb8Ag2yat2cCrt4eCiqY7wCe8V2yFssITo/Bm1on5G8o6oSFKftubzw
4+CdG/T9o41KWUkVvRDJ6O0QlLZHHUBy+0CdXT7n+MbvDjcTqJJ9YzcNsE7i
w4lm/NlIwRVXA/hMNZZkkO5Kdu9dR7xOvBZEgMqOmbkp8HVk6sAhZ17B7K3q
sMi18/8N3j4GLqbHwNnBoFC8Ur5rBxH5aocPHs6pAAmMP6mlykOOVBL16q0d
d2eo4v+YHjj5WFE7GJwtZ+a+vXYRyXNfd7JJH0hOXYwpb5ODwFUAIOm145f5
CWZUSCpanQwF3aWSLs4TFQbJ9P5ds3im9YrUWaRwlVtfwyS7BKqT8hn17CcV
9uThPM5Ck6NoEqtdfEhDOs1m+pk3mDdSBEApu9ZD6Yz3Y2Seoa201nq8tB6D
npNHgWDYeoqyKr3x/uhM+D/n+97LZ0n8po0FfALCrkzo45VkIzZGMOvQHGGN
kM2Py2zQAlefs95vkMmzIRQpiOtSM94PUhGO9BWWx3EixFbcI5pZGGWmbCFv
mCqQwWgbSoDMiN3+JjvGfAx7NHc4LndyEJYHdkcDUCAMT+NKd2T+tiiY1a6j
E6u29ZdmvO8UaDvjrhhr8zOYnGeo2ZL4jzhuNR07iCaDGClfm2fCSw1XAcnk
QPss+WB82r9VYKhstihgcboEazyHSmWTs5qqNVMJ43Tqhu4EBtjLQNQZ8kOt
NR9jfyICZI9pECilnMWEmUQ/AIu7dS0M89q2OC0CrQ4aHO3akEx7XKNo45pm
fBCTOiOPIGoafK4WkZNeToe6NbSOm5gnK+QLjoTd9+p+pyOkNAFkC8rky+89
8bx/6E2Zv2zDQs30ZHgPymVuqXuQHvQ7hn2JVqAiEuZOhfV03BQ5K54KbCKp
PbHjxk9efd+QNBsjQpiZeF9UJhEKejb22YHhehGwNpP3cyn6zAjj4NIh4xnm
eaAffh+ZtQQslJ9BcDWnTeGnviZbcxQusu12Zpmr7AVbF7NdSHFgX6QK/XqG
V6gPW0+qi9ATFZkOOQXzkztjvfvFkUiFDkpex1JovcxuikrZpTyECPgdA46q
PnixWLShjHuPo8gOofO9g8ExVMtKAayPy/JOSImvCSoPaBYVk1OmG9xA8LSA
ufnOzKlrVce58fX/lhOL/NPPhqetTBwCDcR75pTFXd3hAuRT0b/g7usxjpaN
s/Ft2jv+gW9w0/r0Hhdb94Mf9NF4n94gSAb/nTdA0nvI14Fap33Ct7Wpwcss
VBFbV65Z3wqTX8C81+KTUFR6D2wX+2aEwYbJIIcu6pIyNUaU+ImT31oO29/Z
E/fvcdnzo+DBUtceoJUQL7WxjZjdJVzvqhXr2+gO1QsUyJJOrHAFK9UnuWgm
ydrF8SIkzPn/sDyDSqQ4MJ8FcLO7tvkrEOieGRq6VskTjpGuvzP0ALz7MNH9
XGtd16yF1q9o3ouCMlxpfVZ+AZXoZANU17EP7cSGvK6BcDKFmQNhO3KHodRl
z4HRa6YErl6+hn++k2DIovm5ercxxxJPzloJw0R3OtTPUKyqtdroh/yb5pk6
Tlm+h23lUSp0WQgsAk/caLK+OwXQ1V0ZvtH5MCtFllH/yy3gM4HAA4PtRF2U
llsOg8NcK24wRmoY34kwH/ufb8iH6xZeVnZLSH6cb5HJKfGKzBOxlEmcqapg
gLKQLFSVGfPzP23EuqjUPski8QrNkma/9NIDCT90LBc63pMZKaH4Q066xeT9
sImhFnYFFPXnDney4dsyMkshqzh273gW1akARQKaVo+CLwyj8xDxPHSVkbi8
eFl6rcRCjVjsdtZyaXi1nT/XOy8c9ust0ecXFJcjjAgpsG6hYwn6xxMLRkv3
WUxgM1pe54CudPvNvs0l7n3hODMslM/AGtDqESdu5YtR5Sh2NYGAXv5ZYXZ8
IAcn1Vd3KGbdxzSkNqU41wsl9XROCWCwtP30zSFa7bFvD1LNeCrtfyTss/fa
ZO69LhFEJN95fg0DPtNgNBqHPhhlHXRdcq2so9TRiobSyfXdo039BwJf6AEu
HKuxkHnDISXUAOm6PsBhJF4BDyizYpTBY8G+pr/BWjEHuOGvv67z4MMdRyZ7
wJj5JCeQNX10tiIZaPci/LCUGXtyZwzUPjdWX8irIRuCT6oCSyBlZjdnsJc/
uoCAJ5EBYhX2EDZ5STjb7DHQOGtoHxP6fV891jHXqMea6Z81o2HTYDYLefzN
0If6KdF+DJCuhxqwACV6Cn5c8C5rNbtcJX9VLJOGXXUFJqQIWNapKNkrkn0Q
1HP3IVms4LAOLGiwPq3SIGBrcyKNrRWNMYhZovqHVCD/I+I3Es7qFzImKPGK
o9U1daes5tm0afl66QLd9T2aoIno9q9u9vLVe0Uq1fZvkfnSLlRvybuACJ8b
mTe7fvM2xOuqb+iSncOVavCSs4uIVeWz8lzqqqGZV6yvdeW8f+E/fq4Ucaxj
U3lu1PWEC8rJQoBWBOBrQj6C9dnUOZDPUuvwgA0aoz3mXaisf+jTB3XT9V1K
lUgpuwOAdAlL3B0Vv3eEIaqg/kelhZtgYZTtPJGqn9whmqrGaDNbC8iDH+Af
07QsFsdlpbM1LGhGekuhS6fgGY2jnv3Xq1N/mPBnJMRTeSjllaz0tsSIGeZF
kGkMgkU3UKbwOxmFYeKyJyfQM5o5wpZq59WD1AJ7gwNwye3h4V9rnkCaegOc
iUtwB5epNI9fPV3jH1kUaEjXLzVIpk61YxJDsut6862QQVE+PGmtQZAjpTVR
O70E+5Gp/wxWQDsxIaAAMT3aF2uFmJHcNQ76NooD3DbujmwKtFzewU4fT7Wv
zb1wXLAlEV40jqtCvfmJo0tlXlw8H3Tvs4mjXY/sx9s+0HgZxQkAgiL85mgs
71ydeNhwYMaOMDxN7rzNwQ4ITichPkwL0BvNPTUV1p6lYRugHkNAanFYXeh/
EJtSRLYD/Z1qKyDJ1yBvhJ45d1J/0TFGk4OcUt5xnTCojFeMDNIXA0Lla6Ld
CbMeUZZBoNry2PYwSYXfUB03Jaa/HVTtSjLyIzaV4mwARMhxG2iHBZqmcp1d
yJVsm4TMw5GOvrS65ejbWpSshM5aBimS/SS002YZ2wyNq3reDlaAjoNYo2TY
2Gei3FAnMTLf8EBtIFiGQU8Ynd+P7803+tyeUrsXSy+OvUMw69JqyVznwE/4
oKuXX/ozvrflMdX7WqFOgVK4ffOyNjFdTMZ7DNbyimj0iEQSr/orZKwtoUVp
BTagrwnkdMWHhxvWgVghQM1aCcdrQd8xzNB6vFScgi9OUeOwRZMaJiutHl4d
4O3qe6nZJ0IcxBotGbOdWy7PcAUsddI7TRqVvhSMrS4YmsiXOdnIaiTpi0tD
iCEef+eVoxr+MRRroIs19ebuSTkmZMa2k+wnWxGxIUg3rUCA03fxaqXtZ6kQ
/7WhoYcnbRm9L74pFFzb0trqRaxnTTZRWO+7Y+bAww4UxhshrjYgt+EprNaz
M/1fyM1yONzTHobN8HctVMMwuquVU9dYMqW4kV5DEcUL+9ystqn5I+HzNMdj
YoAZO4V7sGL3nJT8G4wNW+FeIuEPXLHArbm/3JaJrRFybnZNxYV3X3Ibzc4J
qbqp1enYK5rIVQoM5Pv+lKCHzyXotLXHjj9XLySM5gisdmP+1SmvQVTa0Osp
ahicHroA6g+bqnrg+OuGRFZFfhw71q0Py56mS1qKNFKv3YWVIX7+/gMpbriC
zb1lekR++uiXzKINjLq/jjwpJ9T61sPsrYIJxutV+wDzDD6fRLxNtxjNd12R
FYqSX73MLYc0Rzf8DG9S0oevO4NkIAxz9XNKhiGBIratNOQ28jk0CxC0pedj
+W352ejH9lcHqa6BEXd5JaChrecSMTv6xNfh5xVi4kKVsXrWI5hqi65kaIIR
AZK7Hzuxs+I/NVWh7sali3FlQ7uQ6yxFixW8HCgqfBC6sNG8RqhgiDXxYjNt
uB2SILn3HokRaBPqMW+fc2idiWLdcdwrx/2rvXTQ5EnKMwfgllFfFl1ePS4j
vx1Ybe2SLM1LcBzm4MYoTh7Zpr1+tdrHPoTYZiBVmA+/J6S9Saynx7fJhxhZ
4PfkHK1MXvKglTrWeD1MEaLVtIz09r07cvBs5J345eGodhnbtjbXPhFRBx2G
ugrjjA0q7oe1Z12u50uhGONT8PfIDfEx3zDR3VqFx5JeQkodyn+l7Oj9oLdU
TtvI5ikIoN38Hjpz3hkIr1i/H7dkQ2B84liutLwD4DSvRkiwPw1TaI9t/DdZ
LhK+QbZR0HTvBpTejlyb8tgdOC8FbBgDVau6WKDIo6cOb0T+bdJJ2jzpVi1R
fwrtAbmN3vyLwFhEKUpkdnJLzHLvdRvt8mhBAJgmAMS4rHbHbKzVHtzEo1Qv
J8YyaIS9ShbRoXRJsV2UFKZtsSr8iigrm54e61JpYR1aCL+9ZjDi64fJFOO5
11IRl3bBn1ZMgVZ+GhlcNPavpLXaYdOcQSV6q0sE668qBfLxExwvJ9MyrwKL
2H36ahRz2f2Jjy2E83f78WzKBTyjoC/AJAunoTsamacrf1n5ShLN1/Prp6KB
wSbbfjNFqK8QmW4tR7WB6Y/eCt+tN7gDy/dYC8dqnwRs4Tq0H2aEBwnoHHpN
rC4S+pSWHuuuBZe6nER52AlZ8yUhVZz65BrMHxmldmM2KJlxn4b+YeBRwiz1
xOz5EzoHiGeZsQZXxcArn6wTC8uM1YK24vnvakPM6S15ZGhKxPJ7gkG+cyC4
UcEVElvmFDLIdRZ6ykm8iCxoVNxkdfPY9EbDR+WwGEviRTPDH50SilAXsdJm
ApSxzjfGfJiF+zdhI2Z0ZUzH0mupkDIZwHjucFTFspMgZRPsg04AxmbaLmJD
cN8Cm8ow06SnpaEu9pTft+BOttD36OS2UJTUhLPToQkjo30Y0FTx63mu4eW6
0d9zz+9U8PbNd9CEy8nq0L7Np6V8FEwt5gfoVzUZbm07CDWc8b7RG2P3aQ+u
KcSEQng98jUNOtgSuay54hWJuh2MkroTWADra0lveDpjUiKyEZGeY1eh/EVk
3sRRfYZPS3hwggZnYsJgh5WYvCDU12CQu1uud/UykO8kmiNpDL0pztbErH6w
QmSjrXI3lt4vKEfGujQYV78r3F2q5DKmv8khkYlYJbQfxH0ZElfET9urQh+w
GfUZyuGduxMSX8jeg3JTxw/DSM6jvVxJE3hqnYU24UKBv5pBFSn+qmXpPpbP
rV7cL8xmbXTKdiHTsD9Ubw2bmiG01IyzeFIsRKr0c9OsUiVwSSYhSaXfYdMa
5TdJ06cYh6Zu2PEGaT5LeMUVgiQu8QFMq7Lo7DEYxn9yz9I/PZcQ/mDJNw7V
Qzn2Qmm15Vrbpuqa3Ugnx9m4sNkkRbD+J9TcS8iYT2jXCsAjkMGfkOda9i9A
vQjwQeJwwNFG43kEqTnNiemDhObdGYPD/Az9zPNBgN52sx2v8CGp56d4YSMu
NpfgeqG0Qj8VRgPu7Od4kZ6SffGu1j2gBauNEpGCATlZ8BSGvC6op3APOCXl
gFTw1VTTFAxzDkoct0nzJNg/nexqBVzQpb6cMxmSQOnIN+Oujp7n4MUwKFuw
08HFuHV0mkSKXYWXe5iqSpQnX2jQOO8GjZ4cFA5CBWtqIWTOmP+PgsrUh9+o
DBI6srIdBOElyU1CARkd3gVHOePn9lci37F8lyM/peOmP0Ys2IRQ9qVP/nzQ
rK1gAbHTaMpiA2f63Rp/6TddoO6apFqBKFTmSfCuDd5gs0gdO/hlu8s/p7GG
pUtfWfnifGR+v/KrGd5/HpTzQMVTZhgmZ0ThUYHKBYNP8Cuhy+ROXvdRhrYR
6dJjypfrNgJohA0fCDprk193WiP6B+7w+CyAkT0qjuPN5acSpnff96SffSbH
GYYCFfhVtPNoM8pdndWNMRPC90Ncld9Q4wO/lE9r7GPeQfPEXzJhBwkAEvo/
v/WsrwEUDPgFWKGqB++CKJmuXehPMk4GEA7X4nkmMqTe+h9isbZy5TMbqMwH
NcyX4ZeX8gld6+taK32R8VrfIDxd6isOeXEW+pbUzKC17OPXCf6V3ji6JT2o
GLba9y21k9mXCEx5xvX1qpEDZHDnDDSUY8YzR3Fz6JE6Yf3VBhGBXRUixS81
gtuAKuogCRlZ8EwhV+0U1PUAGTdnRZtAIME7WGPTMYD6aNB26BAp9kDITPX8
pqgJUECNGDuU+kF26d+0trNUcW5u/BbYqNEqo7PPLMmAmT6g07mmmeFXWM26
lOM+fSEytW/r4WG7QqoNiT/4Spb4n1WILh0zo/i3yRlfl2epc/Ty/q/zLy+Z
4wSyBVvmP+5gwjvC/PfX35qCeBROVOG7YbAxWMNncV4saIO8P8l9ceOpcx0Z
py6UulohYxF5YxqRnGAqsOLqKHjZcgyU6ojlena39QKYYHrYCzcpTcFt2lm1
K8U31efp5WDJxHy1B9MZQS752JNurq96TKRTBbCoNZdHEtpykNmJwTuzQfkO
2V0RwdjZ3H0aXbTIvqQnDAxesoHa+X8iqCCb22mAyhJaSNCpW9xtaje6pxyr
VG1/kfgi4BZv4ZJr5Rvw/0DchRRKKeHWxWYx5yfK3yiM0oKxINbyY4Ugsgrk
GyfYqoW+4WMWvss/F6K7aqXuzWvTHGtF8jY13OTsGD/TsAvtBllZ2oFePcPS
AXT5+QvkS/RvfXyDP5CubUo34ihxBQRmxZNUnFl/fyhBCH6yBmHgNYTvFWdd
UB3SCIffJb/zMjQtkiidGW8mT1CUgjuLF28HMdIFlXL9Sm5a0fk6mCdxTGmh
RwXhU+r2mw0985MKRWDUzxJ54z8mMjsZbmgFlZrNHHXn3ms02c+QPLh3yZUi
UnH0QbTrXY6jNatOqM6NKgS7mawV7nlEX1CusVoHbIddXTpkTQa4QHp/oxdn
D/cOT7Kcfly3ccFwdG3dZ3szyyOCxRtI62LkILz20Rth99Hfpiad0zvSq4GV
C61pKdQiAn8IpQNAlbzdAw250KUYvXGMcsr5V88ORu7kkaHswdz/HdjCzO8T
fsPU67ZVHXwWsr98nqM+gc+JckEkBOJYoPn3M//Ztz1Bkwyvv+vTYeQBioCP
0boNDeROlsQPe5ani1wWcLW9tnBx+5BnBR7UirB+lgFeVbdfyQw7a47n5bLw
P/6pBF5FzW+N6J7A1gHELRnMZd2Q9naQldidHpZ1O//TDIluix7aJXGeb8Tx
GgC7P+Uc0P/aBqXUcPK0HJqeEOv6v9TfRkLBbBxfHJToB43w9ltz/rzZ+sQX
RsX3mS7KAmZA0J4drg38I2efVjEGctAEdJLe6YlD7jUm+f1/f1eW+K+HOZUx
efePqzChtSkc3lgcaxRG9SXf+/3JHUKFJr11YOQSnBnANCbyyIOsaY1+zzyM
9MCISyKMTa1KB/7pVRwQnC9yf3svXgByv4Xo+T7vJDZQLI6MiaEXdyuwuLdm
ZUuOk7RWDvUV+jUZUG3UChKEZYRNehMOhkFicfebsdRN+Mvu40hRwV7s+ne4
z9BG2cMHfZX1k726GLp97alzkzrE7CESwNCaC4x6/6vEqi8BcamIjdyLd/kC
tYzQFpccoMDIQydT5k/wpLgbq+TAEnPSO8g8OOm3Yu2JYRpJZ19YFG5vItnm
UIYOv8c7NSwF0iT8VnbnrkLkZJVOrW/HBgHYhVy0ZZhvyYoNw+w9GP3qaaN6
0Z2P68cB+P4hnfujbELuBZyIz/as4ts+73ffUJYssmrLFAmQwwr1dqUZYplc
B/ZBc+wtxPynVMEhqZVhPPRKDjeSc8fqdQBc3WId3mSMdkPh9sjSeZvjNHy5
SfsqalN1uVbIRq5u3zeDrX5X5qe/xlI36JhjQJU5xB/Rd4/mzC3iqk0Psq7p
3xCHehn6l9pkfFYsbSC8ll3wOQpTvhAV1YE3xqIYJrCNCdRrnWK2reny+E/z
vfyNeUWiZeqmgN3FfZu0HPqvqDXuxqDQTpD0qq2QSZQQ7XVCIZEwssEOSzlo
wWwQNVCUTQNWru1/RgccvwazUsEEOA/UCOl8lytLwR9nMLTHb9oZKe73t1FX
JF/np2QoEsroElyHFEsghDGITtOoFOLBHHdrMRtSsOyzw/xotjVjYIqHNWvc
iXH107CZvvvvnF/8cyM4hO6b3xCbPEsy0edisJGc2aYAW1uP0HjYJQ7QhY8k
bX/edq2GeqS5xgmHFPwR/DKEGykY11qN6lLpCQsRNyn6iEsWOXxrV6rPXlVj
G9SQn+vRJsWf8o6UHl6mGPTUZaGP476bhvhQu/k1dUjzWs4FLPOBuslplV6y
o2ztOZ3eHjwfeoAuXl7iuMtxy41TRY2XDUhKq+54PCyfhEfnsq3KWnQK8jUO
3uCTJsaFL7zQfJxGN5yzOkd2BLsyHENsT+b+dQD2Gq2tsKVF7AXNcu3ekxgO
5lDZ8QS2fx6gSCdiLdaSzVpMnYf5p+y6GyvH+4jSgMPrVIlf249mIa1KxUeH
S6cZPfENkChjOok9mGetsnXIFA8mJR8+2ePczt8zY7Y9XNBwzg5B4E0VJRCd
sy5w9JATwry+JwHxjz6ny68dTNvbAhcS0cwzLvaGyJbckWr2O/7JjWgcsWMe
kzc/Q10ZdXoa5O+CJvBDSFnfxY/JXVuZ7nISlgkvkplOJMFLWemTBjzBFVMg
jig7t/+oeRiqR1LeYJLVMFFb5eXzLr93hpGbjRgH1oNVCAI5dGjV5Y+bBSma
dLkVcEy90hReiE0Lr+9w5xKrOi4cA7uMs6/kFKYGTx18szSTduK/+EjrQLUt
HTpF+x2ghO2SjCPhCvYwH7ir7EOIf/aTVwMBr8LrjPCOfBNN9CRiDahfhDJI
UNBV4/z/H2KKQviQE900dX+wYQ6/qFKqXDI08QfKENnvZTXjXOMCdFETvC8w
dKIzMPtDuMqsPrg5iKv9UlQKTUWIvkNsiYnds4PSiMC0cJkP/guqBH1gCevR
uR1MUB04AUUsgEA4wc/OSnh+XP19NEp00xeuzFLgkqnyZHK51D+ciTVqyGhR
lOcsxEDjNsFrWVM05RI9b8OWpGYpYuJ1W39o4SCsAvFORgsS7rLPng03Ka+u
zwLwyKqS9a3I05IEQE77/sVYlOx2X4diEBqwOObTCUvfb4v/as+bVP/F+lxn
Fd45da+GMUKbnwbNVJS73ek2nY9xSvGGBVIfOPEg5e/zu/JzQn9sYJcS4H8t
vpzc4K6RaiEswkoh8SJdFXJfrbMaaU69R7VvG4VBALOgpdcJFjNVzx6ecBv+
SoO14Z48c224sN5Y/jdBYePY/U+KN58v5s22iaRZEDHyEXbffwD3AUa2V4KA
2sPkh9LCDoo50s2JGQaoGnV32YiUBypjuNsbd6+XcRif994mbzduCpXS+YYN
UEzjSyMsEypl0qEIJsYO+Nd6SxmFttYeLOiLBZ8F40SN7VYRVorA9HMo7dfB
Su9E4xmmhNMBBh3SpOt1+st3Xch7rlJigJmgyacBS43TqwSwpcwrxbjghOQ9
+Ov/18mubnOuEKGW9l6zE7llF45TJwT8/NsTuRYa5vv+iAIbzgnni0D1iNW5
LeOlRa79Ks0qsMnCJ9L/UAUp5rL2AEQ8iubhVc4X6P5fZ5WRyF6heiIWZNGi
R8hnX7AdYoRYEy8aB3n4MYOuVGQZRTJ/H7XYVdtOpdLBOZkzb6q3UCMbndjr
dG542Qfzh2e/BpqXns2aluLHE6zkdYIjJA8zAvY8nBY+aK0fL28WgbfpbPJD
dt4m+99BkYNWqkHfwh4BC3Nx9uR7ZPtytCCHLDxkrQSQVbXqObuzZ8F/zVwr
jcEmEwYJCxOAKdMKePB3HjFZ04V1G4pLVn//RKNKt6wRdHovfllF+9x+vmi/
GXaztoBFpf+pEOpswEf2QDWtsEAThTCb3CtchmqtcMG7eD0nf0wgTYY/9vRq
n00KM16ckstxsSR27We6UjqBYlvOHiafTDsCEq9auKDjo27XH6PEElQWIC6z
VTAiP7AIuFFn3GhzW3gNg3JCqclq4+6Ei9nMUcTzd3qdoEsSi4RE0yTdPn3s
BzQpsJTd2GORyM0um6TSxCjbwUiIe8fzZe3umKVGTdU+BbYOXbgQiQA8GCWV
ZzUe9FT3UaX102oLJFWSnrEZDtiFIob76nOajBfrLpnv1XJyQuLCgB1wmdXv
fzD1Z6MEgenYiwFCK4IzUZv66u82lzTMHFFSuJ0yOmTEFo66sMDUpyGq81TP
gnl5+u9DbZtwqCEk/KZgDIgQwmvuhTN7qf8uzOyKf1GtkxcoyeojIBVG6AJb
Jd1eOO3uPArP6U0/OJF0/5Tuy3Uw5LRgrWhqiSxyTQL/zTEJDYAPDgAjMMJR
sqU6RMrW0urscMchhOp/00BUYZIizjz13OWOaXG7+o2+D7zry9+dZm7UORp1
P8P5iQ1Z2dEThsglab2VVoNaYxBQ6s+M+ZLXR1Y361MmS7KErBvD4LMyWtuf
y3i6WclLTTGhi3AmE8p2yKz9OWwkVJhIvxfi0G2QIj3CY3WIkj1j1kV6ci0Z
d4I2bq3cUvN27dFA0R/KR5+7MOfdy9x6vio3PmbelMwQbjCZaVcrIv1eciN0
cXcvnge9dbVpMUOTJQaIj4IJ9rOpLK/f0RQhWLw/eBVX3f+dfkusvf9E2InR
W0caI7Np1EvLuvmm9bsmE9Nayb0qxwbC0V8MCsTHydBXr1A0F5Hd9oPcBIsH
E5gTDJnbEbRrzdyp8koZHywkqymFCo0WA8rPh5Sj40g6GLO7xIRsEKEBGLXM
cDM4pEhuK9AGbOz7m9ylPMxaR0plLj5Ozy+mcPaDUNQMOWnxkxCqtPE9yCQ6
D/+ZGn7LfHwC7GSuDPBtW2v46owexEhNRjjYhRT0cYaYQoT+R+YO/6ePMAIa
nzKfT2Vh52H+6amGjzwimkI8jovejC3wFjQ54Nxkt725ig7bTBPeYroRiNy1
AQCV5Gu2aw2qHEwYGWuE1rFIxdC5bTu1pNVkxb2wLRAyWzRuvu+BK7Kj1BXg
1FvT7PguEm4E+yUBcV5629Ulbqy6+n4E+RIHgvibfmTNTNSgrDqzDv8vWtMG
1f7qZuWmRpupvLRRVVs8zpJXT7ybDuvCJxxuDK9U22q/r81rUJXQlAkHnqRk
+xIUF0YRmJr+BGIG+/fcUZCNfVYKfuvd9MKrRHQC/Hnony78/iTcbbzEdA1a
JXhSyHl/QBULBb5mfbozCkmOBaFigZjqLiALFM+TgBb5iDgPRAIYtYw4hSUl
Z5ft0m0Wm0SGiJY4Z1RlzVhsLP9ijYwQQqP+nv0iSaOIi3qfvajKGfi2mbY6
JuO84Qp8/3yBVnRM2Dl4Agh0ukaeb+2aT6HC7mi7vxHu2aNM32lh07+01RCq
7zDt4ypSkAMM0PPxxzDeWB0kcmXa3xJTCKppq8e633xq8oqjm8jiiIuI4nGp
3KPrrFjxryPtfae7e85XETJbMS7VYrIoLjDCRfvJ36gylKk50uagvhq9ZFBR
hN0qXvVNXiiNd+4LXsNcfIAn1OgNvLZIAfgje5b71PTF0kVHwsNxoW5A3Ti2
UemBw1Emw+YitBeJgB8ExpO+VveWZwUPgKltfWb+BZANP1XZvdXNNstwfeop
3AChZjrgePNwdJkXdcgHBjLxYaVILIUQPEPsEC2tIsxJFoXavAF7g4ALoPpe
kjzCcWY7I4LZyM3c5SxyAs4843297rLrM10OnhredB4YRFa+k/j0So70+ZZ+
V2uML2VBKWlS2vVY4wMEAq4bPvCHPTrKYLHFwm8ZQRkqTs0Eier58lHB9mwd
iAG50RhoyAuOU8X0ljAuRCNmr8hjAlzrvJhd5gohicCyIumIAgepJ9FKIxlN
pVFrU1OdhQ+xzE9koczV79uJPA3/4ktEQzFya9//tMrNUJBZZwOqzirWeBGz
Sm76WU3yo4FU6McIKoWX1ejHoXB2bMhY0ix3TkbNjwf+XOF5s0r8B2lx/g94
VBNTLqN/V25uHTF1UpXw5ucSYkEEGjHjBPZGXypALaRkbCeiXkizqaHH0noK
J4ptjLEaEIePwr5Cn/0OtMeFbrgo8GkmUccUvcCYF+kNSijmNOtBTVnFzTsH
USvfHz7OHPQ+YtuD1s+yCGUlm8L14q96NpAq2YJJXo9NWj8PXPoeD2Jckw61
lExpFULtV7yP0giOfBTw05coP9Dj7buV5LI50ZgZcc0sGWVTdlITUY3KrZuC
3yuqE+9J3u5J6B00n/LCWqlvLuUz743UtrGSzEAKdFI8yP+cfayzCERlQmML
maNd7sVJSIdPSfIX/4Wl5NJhje7KObRQkN3AdHVLcyduOr1SZvDxzXhey2um
jnu9wx2t3i87Q99yYm6jIexBZkGzHGj58TbC+eRyKSnPdLLo4zr5w7rXGPnv
eqmOEPu9yRlqSAFHHzAzuB3/duDNqTLBHemS6tKxtA4/rhz2e06FDAJPwrEn
KblhbMxjqatuiBFWoFo3glFup7IOeRqV4KxjvTEa51sU7zmf1qw7Sm5+b7am
0c2Y2NqL81+0aHanzi4cL7gXSV/35Oy7+3yZJP6/zvH0orwcoq8tdo4HrTlX
p/7/hKZ6UTQOd2OAcXbUsCYKsnOXoMGOXv9WvkK72RiPAMWb2tJtg/uxgf1P
UgFVbwgtv5DV8NWSNAc0IXJut7mhAkim7xGO9HGK4pL2i1kp547HapmNy68W
3NqjvJK4xkuus69asg3NusxzMarq5yWJSEb5tyJ5lzpEUfyocM9/bcL3rCeQ
rea9K0LmLlGkR5zhXvXdfY6E4WsIhwz2AobuM1xN9lqYt6AW5MNuWMSoTrTo
wOD9E+9zIq4y9SQINXCwEJiJIDI9KS7ZIE33p/iqIBL5/H+xwY3e+lxH3la9
PS7wsb3P46l+QXLjOuyjVhcBKIXKCkl1WqJJoNKGwMhoetc6T1zxUvOiuE5I
53PFGyEPZ62PYUkS///6olVdGweo8wWBrBF5VLLj7a2ukSerg7jJY9f2OeA2
f9gKa3wZe0Ibt0/Oi8a5MWtzsQd+kVLo41qrc6bAjIjC6ligf0+eMlV86Xsf
12Z4hXmGNJMlPNAzfZqrP08Su3pydGZ8shEGANrFpTeRMzFQ/AcksUT7jjnk
uRj7BEcqr31nBgGyRUIZ/+i8nZ7cz4WV7wAbBv+tf2jIoaef+NOQNbkBpD8R
hs6yIWHnSSBAGbs4hhmpEd7AB4YXlP/6hgOtxJz42YhUiQ5XglPrKf0O3ie6
ZN1U9a9HagvMGngLz7LFAJ3xE+JBC++qC2I1NLDbSH1Px7zokfcgNyH4z6/W
zdOzHV8IpFQzuyQ6l1/4fLpUWbefIb/eZXdc9KLz9x+B0aO2XeiBpX8RW5ra
3lXCCq+t00jrh6LnM9uWzeq2H81HIJ9s9Or+VEKGKM5ixMnWHDh2Iql/vhZo
TcYUTJBOXEvPem1+QPNjXO2TQnDPj+jM5j46QBmQT5TkiT2U+ES+l/YCKtFN
z5Gne1E9DlZVRB/fZKz0PIpqegtPjViNAcS+AaJlyOkuuiK1HmTWKTDySgJr
dz+/sfsWJW6MN+FiCqjvni7hg/moVlXrJGkhhu7X8QMm8sI1tiZ3BM7wdtRU
UkBxKmjGav8h96DRA9z0I8Vi5ny8RCvGb95JWYwRaCjihmRxdZFDghdB0P13
6eBDAgTCmOKv9sC0shT5bkbmUkqjWv9Z/JOhXUZ4IaSvKNsZgpBqT8I1Ex0q
gzEGAe9qEyg0IIeS4dpJLQdEa8/Tazw8Iy/5ePdy4hWCHss7FvRr2j+3B2KJ
vgaPlJy5ijUZRxtQ5kT467qlIgad0z01WBk9NUqENZRRLD7SlWWuzIUJIGk1
k4fKMXkOQx1To/DGPyBiZvrG1FTpnRRff7AYr1E6ZsxokxhVOc1ZDyZj4i5k
A5WRu8w9sZRE7WOltoaG0YCvY0C5KKXBME2AfPT0guR7nN5SqEA+oVdslj/z
Erz2Vl7CnBqCAg9puIyfvyx8mXSU2DnGhDo7KuasGxTGuCpdBBiSMUBGrzgb
9n/JuuDZDjHePtsZCDx7CLxPl5UlVhAprR+3O48Ay9tIgt/VSmbCCHDy6sK6
EHITC++zy9aQAjwZLeeDAmO+nI7RtQmSCKdqsXTBNIbytflHTIPo4xP3am1F
5ckSsDv6c2Ct7jBPq9fbm1Tf8kwJ0nwGCeZx1I2Y+ZAfqy5/8cC24op4rs8N
s3ctLxziTsjkQkjk0Afq8I2OEqeQQPhkc7O9g4fZpQFg7LjmoCZAkTwQGKTh
/2dCYB3nULbkoshl2O1LtP2ri6ohNuhgUiupkJuvvaXxtuZISvoMnN6MXyNP
sC1PflDY+Zw/NLc/fP5wi1mY2m8qzC/vXbVl3vvXTU82kI+naHV3ByP2dkyY
RpbAEv/1WucLmwimSq/48MmEiaeteeZdRjYXy+dxbos9U4CBxcd1HXAHQsgH
ujW7K2TjRya0XbGTt0u81EH8IlIhCKJaG+1D+KkjL7WctzP85UlLHUOHpGey
8GX+kzQU+GjvM2At37vZj7Z4MNub48Xt+6N5ZR16iDeSqPjE2BOcyfEXUUZy
EhFsMI1G6mYCbb4HqoGbYejq7pfSXZVEWZuerlnKXshnRUFbOkOqBe9kpmif
3+uEA+EX2uNyD6hWalru3GZzjrF/yqiyyJDnDYU8oWBFBUvqIA6OcK6Kcj/N
D6xlBL7Yv7XATzir+MnwQ72uvbQzjTybn5FA+sHmcnBtesgCK/v5xWdtapM/
9fgzqvlaWEB9HnqtyCb/TVMY2sHGDQjPHc5VRWHz74USX0ZgqQo3nX7yrY0v
r1OOfPHvGOFY+4+25l0o6tka6P6gso86NXRtMcM0LkxWEgym+yAhDDRNdFR4
NN481NEZPOvy5WLw5T4yxww0mnDzSfMgTt3iHwBNjQ+tPM6FE5qiNa2ERfhT
zCQfebcPjSJWcPkOHmC715Vk2HZFd+isFsJiwgf9xHuEdmochHdw+MK4BBi3
SPwOA/WchdA2+nMs0YbTmf8TMUJzRRp2gC0Mc2osdI1YN//wLaGunR5kXBSB
Uog/+E3NUUI/OI0j+ZaKM08WHbFrhotgjbgOAKAk3jIPOXVOL8XYBZGkCfzl
vBMwslU0x6sXv1v+JOu1dx8u+HHcp6jm8WwmhfVT1xXtSmj6sHKZYksQEVXH
xMcEWiBQn1XqCoUey0lHssDjyMrJk+88Hzy1z0k6bDTzCBlOQSP9lFLzX6Ng
8rAPxIJO8VEfWEAIFvB9GV+PVspn2FETeh3mJX+2juEHgpwAu6gRBJyaJKoC
G2XPRrwjVxxW7ebgpYL3+7dPtBSozdJ5OOIzZnXfyH8PzwT0XTGuOKzisCX/
AIf8jIDL9T41XAHMez1DNME9K0c2kNbpXrT0/SrginyajGDEvT6nt1NjR+zm
d04DMSgCxQczLUKFuadfDYE0STkmVxJ2l9d1Uan5V4Sz3hk9z8EC4WZweyz1
PZv2/fxdPW/9KqRlBddgLfRE5n31PsYSo3Plkm9F9hLXQHUEtV8nbpyAmDM3
eSjJT7C0hnWX0HrOA/TONmbCMxcbW9zWSixbu89z3ebih6GPcegOriEjTInU
bPwLOZ5ra2aU+cuLSAoyD1sa5unIg4fXDQvpQasrH+oM3R5bfzc38ED7rjy0
yHSYUfh9sHjjNwSIRXDeZFMaRq7MIEVJSl9mfTVyweu206QembynLy7a+hpX
+b6HfeH1XKSbAXRtXil2JZdgFV5jZ65tr9xtXYtfw6DQDXidlkokS9DamO93
Ra/VljLAZSX4xhwTZSU+0LRubAH6lKtIaQsp51D/EdsOh2K6PYEik5iJpCgW
Si/bfMP6rBKuz/8Vht28BKXXZpj+DRjAoePnnuL3YipSdu9o+lwNLCdOt5N9
45tk6aHSDFBRescGXqoTH4AUUckOSHwsRlfTNZOohROguUEpds/kt1mWsoh6
+jVRsyRHKr0swJDqOWJFpS0E+WuEnj0xwLbBqg+EbPNQpjlU9YvYMudJSNBg
5fxWQlqcUb+3T4IqB8EQh4jjiSY0tZqPbHSp6uuUYNH1MADNQQBSLAJd3oZ7
aiMVUHMlaGCWvPVmF66yZl53drnQcUnkx1yjqs3lKCXKhcNYRXVvQwMSZAtM
5J6DztS0gk8e+hi0fWUx0v04zWGtwrL3fyFm4rM3B5oB8cR6qIxuyJgpNPgo
N0kzyxRQbeJnbt3yj13yYXS8lUfUy3nubXT5UmpfSXyzlvXKBJcOL1brs1qG
WAoaNm1rd0VUmsjECcrYTvFhhplT+rBlu+bVuAVXnB3c7ozZZymJuvMKYDMq
0X2jQlZUocZcOzDN+umT7xhuG8UcDyg/Bvyu/I/8WSiUIp7tMLorytFskjez
CAfEAAbAy6IMjHUq3Ilc7uzLK9CCZG7NSZtL+sBBehsBCQV0CHbVae9+ldCu
JBTSUiAdN/ntxJP5FO6Ai3p/f5XBpz3dwlaTh46f1t8Pb0W5dFkalOvESteh
m4AUTpKhz32WQBjiujxTFVuRCCSONSRAC6XEX2I1jXtymH7wdZ3Pj8dxJTID
1LyiUoYeeN4Il39jJV6R9AXEQ+Utlbn6jD/ZwDooLZQ/YL1IkbHEuC8pQWQT
VN2q0O8WTApNgOnk/hSVvbqPQNpbLs1bYtpfXRTE3W8/pKO+dRgGCDTJC4cH
1v1/81Zz13YsWbOuHFwwtQJbY3QrXQKGev+qeJYvChyDhvD4bIdXODrLimXQ
lwhV6m4sxyWKCKXwMbMUDcBSmYARxDC031ASyzktLGiWtu6QLGz85ov0zk05
crtGSSueRP9gDm0MwtZNvPeRrV1JV+eP8Zk0NVZBZdG1XrQqmGi+iWCMFQe4
I3lOxbGk0C87+PtRqbrWU2HyXboEUgTr24OHl30PkukkeB6VXFwqU4CycjSy
/18LrEaLVmlLPlZmHNANkdfe7Ua5kENRxjLvmBfcU5DfUGbFJD8+rUpoBwTy
4C0/iKXd0IfFzH5eIiWvOa5mzppjwDjniyZWAAx+fe5OBW6Q5g2H3jHUkqEN
p/FVnKlYEpzRt3VFT8GNhdaC5KZVbd1o8KCRq4WPNLFLv82VSc6i+6WnCbHi
Hn2QPlG3JnGHEtEVqxfYz7w1pgt2B9n021ttu3E482m3D94yBv21AIW8Pvr6
JMrTELw7jVCEv7JqWCO49MFaPIcZQQmgDD38xId2+2qfsWfJUX9Fr/BKq3VS
+cP2jjlAzpKw8vPEn/TXtQmJh2CdukE06KLdXUX9lgavgOSlPR3fgbNEbtpu
JmmZAu4Z4//OBzq7MjVPbxjBt73SpWhn5XKmmWCGk/ubZUaaATx8Cg2jlf6f
N1CcaZ/cu3xmTXx9kZM9EfOrRmZLuU3V3jaoYas4QpsyzmJDaHEG35sQxV9y
JssWX5aMj9LExtT0cv0Esos0fhJ9wwhjMG/ONoi1zN7VsqVwbnxQv1iz0hVg
CIfmePSuttBNLRQCa072ZSHJ6k2halQf9r3EKwlwJFsOVdnlZHZoNRjI57Y4
ri0tJN0iexl6HIH6YujSphW5B6eMeDXHcGP3n39hf0RArUjIhApymGj9u9Pg
H1ugUWKJ0n5jCyO7BXSrE82/2tPbk2qr3shyooRxMn93A5wTrMLS+/QjdhGO
OTCEfRghFmJNLKYUhtuVAPHbvlO0QXWuBPVgvFQMQ1151aY67l16n1tO9ONl
joUWysE6dHsR8tuL/iy0fAVr2m6/Pt4QyV/OjMHkt1gH1aVICwHr8ELVyHVf
xl/pob0655rib60Pw1Q52E3OJv8aRf5kg2KGppbWPX966x4ihzLqo+mUseq5
k8QnOISHAkBbqgvQLwBV6hnL9Qm3NyDkGYcdkQeE3HXpt0xjKxycHSQjG9an
jtEGIx9MD0z/dIZ8TVfcJBF6l7sgGCQtWC9NY2hD9+56Igaa+3dSTi/FC84M
xaBD7DOYD6uudECLuGOaZVve8leR3vfERjBOUrpyUSIEEHKGaA8EDkndGsrn
DdK4DVLLyh2ytEz8soRucOxX6fxR59ICeLW7GwGO1Tbmiea4BJ4rLbN76TF6
DtEo1pxHR4tVaIJZGmtb/uliG62FjL8REGJLq6lSSwVIzIjQyOf/KLKO8BaJ
AP5cM2C6muJuu914RWwuaTGRhKi+iEIQlQpvlM/dc+CTtkzS6dWa9Ei7kg+Q
Pz+oCXLjf3o179Ve06r+JudxL88r1Bp09nASnVRVV19h7EjvFryup0Ci8+Gh
Qan15v+O2bskcm+pEiYOZBLpdJryrPJ8aloIo399hkjU1vAx/D1jrVr4da6R
PGGUEC7Ke7mRLLhwY1JnTcbkyDdtInKS6txePQxHYMMXeWHoSVqPyy+PGi2L
TxwRVNbDL0Dfs4YahQyx6Xs0Z+zHygDmsT6JmAruwGhUgbpytfSyh/G2OviL
xUByjvmMWGI9+YTLbrGcqjhqcNNMNtp5WAKmfhykmK2mkc5F5dpFGdOy1BBZ
Uwp9B0SiUeSklkkqecZbi20Vdx74UJwF5W/EJaXx6LDjwOn+Gy3S6hMWaKbc
IIgyFDjxU4QgDdhtP01I/V1ikrKebIZdXkti2083CLAmyNDXK6YYHacpl+ic
Y+vGn70I1Q4VnrBSEci4tyd3hwjXz6/jIbAGHAaW5rZL5suL9Las2/YNz07F
n4Xk6GU1pA9/8IO7/eXx+z3BBvlYXxAZcZeEoQpRqRImteF3Bx6vIDRB8B7B
3koOf3Cb5yQ2QzQeK+hpqcrZhfoqv6KC/+LJZV3LARyGA2ep+myxXUXi+/VT
nrO21M7AKlkimLis/1hu4bDifFasGKsgVIKs4096mLlyMUIPn28m8bVZzWje
qRAspDmbQ8Mos+6d7weYAH7FBXoR+nIQkn+sI5GBEeqWtmAT7vJlF7nxDIOO
kQsz0abk9IX2luz9XMF4oFF62Cm8Kli0l9dQ84ub2xT26OHq15V68x6Lz9N4
dvXGa6MDfSNTNc+LN/NJDMd+imjK+Kv2o+POM0LB7h/0ZtAaKYosjQybyVV0
0v9ZCJdR8qNpW2tVJakn60CAG1LUuQz1bDnQVvfvdHZdTK/5Yg8NfDOBoCQR
lRgoqXYcn1ll0N7IC2w04X+GxpIejylHzjICjehe5XUsuplrq/lATIY1pHgT
UCkS5X4Kw64LvXpHsXlTSxwxD8CS1cUBM1twcqsuLBS7A7HU7s5+HUp88KZc
J83PDR7dlQ8Jk9zZQar7ZesqgWm7mLpoPG/+C0pxzg5tqvCG3Wvk3sYxMebf
XifaX8oSN2eCx5U9apqkrHI1lTgfgMuu5VF7y+kinZd20evnQf+dIdb2EP7t
sXUiIzbIDxw6ENwT+bS2qC6yhv71qyaSn3mJuCG+V3ON5pGtGf6WD/Sxg3Ct
CARFoTIaq4U0TDFwGwgd/BKlVcwM7Ksy3B+9pcCkECkYxar+qDz2FTcHpiGp
lOdlHaOgPV5P2nZl56BInUZf3FcgyVyXxofLZpT6PLE0kRWU/eDUHIxUhWsu
bnH+Kpm5OQM4AvN0AaDA7KcbxonZhpReSFhxN5XEM8j3RQtdF9C67L5x/vYq
UYugxNlOzkvIX4CjWgpiyrrRGW6ed2RbakBzigDW6d1i9iQGDbBaNLOMcpLv
Kuf2qLA9a1+Fq7nl1LZfsVbwW+z3Um1NqllweKBY7DlrbsAHjn+iXY3tiQ0d
44I6gn3lzUh/bMHizZr2vp8tlrR2MgGUVoMTVJym5j2u98OBI4Uz5QIPSUVl
kGCDIuTtpc0Ko9M44dFHsKnmXzMZCkZYgRA5ZvRM2ROKka2BBU2ykTtRyF7f
lUAT9jtawAl7bc50g3XZ4JMFkCBLQBVDwuobNsN+AIcLq4Lx8f/Z+qTcNP4U
3b3g/Pb6zrCCw7tAlMbE787mFl98m78rbE1PhsN4V/XkS1qzdJji3vieLvEC
FIWGcxgfaA7eUEaVzUIDQrY9eWsJ88wB0UsWXOkqqfh1LCMLlaNbYtG+giXb
KhGfIWw5thatM+U/sbFpA7F4F80uUwVTdKSq6SZPFT+4VyCSz1vrxaG6+0zt
+xVjWNKmFexCuVQqoByoPm6Dnt9pexwOla6iOnhsEdw3zC1b6rY8qe10lXUr
aKZoEDa/0MYRoQbCya+/plpPzCwNe0X5B/Knb/ormPdc4jFMbgtpykxcwa2+
0In3esROprnjGfYEuw4sNxNQeE1zzhRQv16aAmfm8CwuRKc4WTkSreVq6aaK
A4wg6bmuIkr2SWtJ87RrAHsDL07O3aLbdk4q+Sngc0RxONi4VXcW5lF96yda
KVyn8+VHr74kILlJbAN9FJHaSTKifb1bmqzOqyAM4ciYeHOKWGEfAQeqWt78
hRuUXd+EMOt70ePzZx9Juh6U3WhIm2kjeeIKgdkxOKsk0XVLxKNlLqUUDXn8
BbDOfNxA7sMUvSauJHrEk6Ejw/P9E9V+w9rt2xbxznTawvJAVdzJNDtUYwGH
6VRrRTx1Cl0dLY3DbG9XYbaCvXas6xo5GkEr17a5JcBGE/HfYBxx8kouqD08
I8vPTlc/qNyv8dxgHntFeWVnke8B7CXPJsdog5Q8mXEcRecyV5kQMVIP/WJp
F63KO2ae8dXpejvvQQSLcNpczCBdYMv17RnjeD3HtJk3SQV/DV4a/Yph1kxz
j1oFMwAtzBWx7EPdWS6MJ3p9AreLla4e6hKo1dubkFyuwkQyQB619Sax9+RB
au5AlqUi/IJR0JxRXJEHGRfflNe5L2Qh3guwLTT6UISGevfWyESDs8pUTgxG
/QeoAOLQvPQNVoIreKN6pTfoQ5tYwpBrmjinrnjhHESIA/nce1Qj4Ju0hWHm
UCFOHzfNROCeUdbh94mw+BhK82rQO+tiQykzEYMYtg2rbsS8+wdPLGtm/WV7
+fl7T9h5Ku2N7dfbpohah9tkUrArsfhm0x07LyvrKq8NfrXkZ+CQ41bcjK60
w/WPNbBv43TnF/45ufm2+IJvF7gcBo1szqrCyuH7daRfvXipZQzRoRqRiD5v
avyBatZQ9uJcihmVDtJz8kiA83vk5ZkNaX93Yf1ASDNCLnnWC5uBB1xwn0qz
7iqZHJJsbeODWgmkGN4Bf9/pkZmOxBJcy6eOMxSHPv5w5D1fQFNUVJXI8g78
tX4Te6hr/+18lJnl1+8OLH+jLy/r+Rmgmm1XNWKm/RA0CgTX1mmcxwMcRibY
zcEJvHcq9U96CiW/7lPXVJV+MnQEKmSJ74yEvwq8gPoYn/zP0tNDEz8VUhst
cmWuvj2X5maQkk4mQ03MykI+MBPEmPMMPCw5bPkfL20X2hjH4XLXQmlhcaIR
yFhTk/ObLT7kIM3OJrp+wpxrLaBFcJP72um93BkoIdUm2vg4vCaWuXe4TKUA
GGGDzntMGEydXrBkp9U/FPZ4KRSgtUUCrc3tZSqU99VM9mxIpYmojuRxWbhm
TK2EKPFZDg5MwhVUKvW7oV3FDc4O7ePeMnMBgoxctawFJnkbrVxLaMPewABI
Sprv3GOVhT518Zr2fId8y4Jl9FfBr/h9f9mNv1GisNWEcBPIzboELom0fPeI
iXDJo2AUYTlhKLezcEdNjNNP4WAtY8loZ0oFAjN9bsp2DLFgMA7/3rIGfQ1R
itpKOsmbJPntfk6fQI0r2G3sPWL2l0dtC5+25UfyNFljGmel1j8yE/PSFuRd
2PmDxmAwX2OmXC3PqEfBC6HPHJ9KkHxzCHZf7Kx0XRpXoGchnrTVvJm3l37x
s+Z9ZYgAYbEAcJFV3k93yHt1jLzEMs/1URA7MOqjOWIEY5vssKlOYNO3Xy24
h0aUSIZ/dhN9SzoviZPBO2FK3ETzWrsX/0fWVKrIuT12HWmNmstTaUFyDh7J
Uw2c2G/YZ4rIqm2+iE7dRRCIe2/KWPYOMTGzvApB8Ll3Uxh7RmdaCNczTot6
9OBzL1QXnpH4SRVCnsuazAY+tkNQoq2fsYZlgpDh+ACaOE0ycHJ/Y/AyZb/v
UqhASddh6iopZjUuzFvdkcYRDRXm+afPWswEyRg3BOBbwaPNhTdG7OSx0/vf
2+sl7fexShIRTCKKIZfWBiOZGh79MiPuZDjp0C+Ujv8PLz1bojD0NrrJFRrM
krkVrBgm9VbriWJgLuOa73/wnNpeg+3gz5SQyswTjj5pk2ZPe0XdI0ah62yJ
PkRg7rBWr6EEEguwA8gBhXxlBL5sjHKdjYtZ9NObiqP+oLD+stJRuiEPtJaI
eWZpAgf55skTuY5orlDHMAz8ZNbJp+fZ/F+uoiHu4tjoMfqKhE2bMPQUL4BF
s6tfglUuT3ZjSRlZCHHLXiWFd7wTllhs8urHeWYmxGY8nYL6X7lwfo43x70h
zicN0QoTDoFZIH0A0Cy8l9EqGZ4ZC3BqUWGFyJnocG+QsAPUCcQ+huaZ7Tfu
hb+IxGDGH3I5S+iLItp5wQNKuESef0An8LSsYsvAty2MKzxC9eOK2H01StN/
mzKi2IaUy9KRK8tkrBG0ZPzVRdyNpQwKHiGZRp5sT3HbX2wC4Lj7CwDtPvYA
R/C58/lZM850k5BLzY4YILexckfvHM8pGkeWj+k0SUVha/9qGbJmIMgDR1pg
0Pbb0rS+15ZReCQJhAhvPy49y//2q1ukbcCg+g23Y2lzodzxAjzpNZKhLJlT
BRpudAW56F1K91pUh3RusSoGzo4jfvRxqevp0qe3CuEd1JPUdcPDrTbXWi6Y
s3eufwXKteiHfLOQmaNRKE1fhResok6kEDEPhdKjxB+o44eC7W0qdSpqXLqC
fZrA7sUGhv8LKMRANZcY1MG2gWrS2e1/eDI23d6O/T4ZwqIKF1oo+0MXdqNv
ifA+3nS6isgfOvg61XhwF9d24Echks399QyRsroh6l8pqx5XHQLuS5Z/K+cO
8WDSPTXKnnMAG7xDY4LF8XJslv6IIQT+GVb8dD+yUfUmVBzi9DsiELqVmHTI
EULa3Wg/jR0MgEL4iFFPKnVqtGgzWVBtAbwVQYVLKwiaYaiS6u2/ncG3irWT
S6mH9zr2srhxx0ekAxKqELUpVMwPO84B/CbebYTKqG6P7ihWcqWdtGOAPCgS
aeoC+IOGCIAOvlFBw+YFXSe7XvO46v22gk62EuqWR3G/Xl0A12dEYekTAz8J
N7r6jflmgei7nwG+KzMvY/wktH5HxkkYvnbUEQtHtBm+m6JK6b3w5W5uIAV3
Yu3DK/JJ+LBj9+Xk1pZuU5u6rP2itj0h9U1r/eVtvWOM3DceONZKIWq+1fFi
mNHTKwDaABpRusAn53VfO7Z9XGbNCuHYyxJeLiOnHoFK2h952N5qzXWr9NlA
ZzSSqXfDCeQAd1oCCNeytMHgsxzkU3G2nLgePQqKcYLzZlomvnVi0zgYAbCG
1K1onF/1gQkDMAm+oX0D6V3dSJf3R3iQErWKxDkQIHsE9N18O3IUN8/3SMSy
aux6HmU4FIHBwx6XkOamrSw1boi2HdEdfEZ4MEOzLXArHlkHUqBrtEbgC30P
NOvwRl2ZIH63G4f024ZgrSiPs54l7R6ppg4owsaoLy3gI9TxFimKFoV6v8aj
1oyKHB7xz1V+w3dMp+hJPZFrM5c4D6P/bC8L8ulMmtDtq8WdQMB84UMmBmzO
a2jlziuWbfI0xY1SN9mIetqNBvWsvjn4Jx/YfqSE3zh/7UyCeZ2O22RGn4jI
425ODZy0HqzhaWNoz4n3Mb4Mo8UVts+txeajy7xKf5CDD/qLrnb3SqKzrzj4
HknbeKJh7c+DjSljPyX6cvCV37h05bR9OoQ5wR9ztGfsTKP/qbGMv+dQ73gh
SgT9Yh1Ssp+RekCaJLXR9XvYYsT/SdWXL17Eqm+xHMZIX5dm72B9KMErzd5a
hgFRwv8iVfp8smlPAnfiHiq4qKjTNDKO2oYahZ+ni0cf/GePVT5XYFM/vv/z
M9ePEniG6lzznQlmpYnFwzzPh+n9kfmIlCQFYXNx6mVGDzuiehirH5N357wo
bugvtWYza3B2/tp1yF0Q0jfa64S2aaAM2P1gFLj7dwS6VvtQRLRgLcx0FbuR
2eISqku8nuaPRLXIVcQ2UuGFnOmJTGvjsBtVh6G6aYMiT4HraQ722LpAexHZ
7WQRqRMNujY+I2DhcQgPyNkAytBKyEbI0wvEsR6U/STaAAmSsRZzLPmvC0ug
SjI8Wkv34Sx3vX/c8TQirTXHyVs6JFc2uCrEH2qF7XB48yD4bxiVG839bCau
D0B9Dxy/RP0cMQHgwU8+ofHEeDyCC4KKMjn9u0KQpZoZdq5tRSiZC8R9R6je
Ub+SIrHo1Vw91inkClEUHr6j0dMhLPTq6B46Cbb0WcDZzhpESlqy4Ihj/m0f
fqeVHUjXi7nneqSn/uaXfIZfxjjou1gmCewth8zD69mnDBRiOGltC5PZ0K8r
RPSeXrAm9VmQyqHLGEVYrE5WfsFqW7SbsX20DH9RgzCwm02YntRmNianATB+
rl6rGAdRUzjnfufQ25STliW4haBmbWN/PuBcL/8Iccqyn0jkFcRxxMP/V/o+
eo2R5E2UdBCUdZA5QijgYpWNU4nGRkoPEzv9H0JgXaWpthuTz1OElJTK2D16
fuvCZJpbZIaEY7DrUbZJRAn52w2ntP5DtA1HwD6Qs6l7VVkyRgOFJ4hHKOME
nakSk4NFqNTANSpHPGMQIpnIwiYtF2lvjlfB0ZXD4PCbJdJlPvs+S8+2Rd1p
xGUUUHXg1gqvMPwqzbLk5BNnBTCzynH54usEcs+2qXxN9mN9a6WZYtv3ElhN
stbjqGjXIOJed2VqF/ksHPep/bW8xCFJMPJ4BAeeKBiflQDMe5EPxp0snlEI
AdNQuLszSPfqzlLUyg+7PenJr/TkoH3H7zbj8fEMcfCfdzu6pj7qhiGfK0Bw
ptDPzrqu/0q9ofbn+gW4/T26iI0743wtaUcoiOQeM2In3Hv9m9UHjJSuk7Af
U6OvXtO1wJtM+Pjejof3jA7d1R1ZD78q7uF5Alr5EUnSNmpxPKapIloyo81I
29DN1KVnLjo0nuAl1z144o59OjtR4TtZd+qGUyaULQAqDhYAIyBOklzop8xt
rLgn6T8aC8m1ADB7CwjhfI/T0dbnTvPeD84/4pnBAM7msXB7IbC6VmZg3vwC
tM+ILukP4gnxwt2FmyZujKE8t/GzLBx/UaTFUM1mXOmRDYseK1qIZkdW5PtA
KpKQV5gj7ohPc9mWwlViWDiYGB7wnFVjI+ln4BfNGAoLmPm1HXDna7CRzYPe
2putX9zQCQpk98CVsVaQvweglVj7Gq88QvQSmLu6o1TmS7Pk6oUjRYrnJe21
VinCePQklqq9Kj1uwWVGc8EJaprZRxK4RjyuSC+/RhD8GGfx0VOare5GTwPx
Dsy6X2wkEGmfzwfa8a2upyyFcj11trp3QKxQDh7lxDWwNc87bprPfnu/5YKw
jS7Jx+HY8ww/Rq+Dpf7azqH1/wVOzGw2mx2uUK1i5WB28liSeal1P6fbKNLq
hxRKWqJQb+aSx5hRoIbiwuVOKD7XASY/Sm2S4fKhXNOpKZTGSoyj9qaYqxoC
QHvdeNIwr2/UcllIRTicj7tok9kzfbIqmpe4Ep0GF2VdCPjY2W0taktssjwL
gf0FQ0ug7XWedbNDYCbE2Z7GWCwJBOYR6DZacLXOLM0F4tdU4ssKlsTMoqyF
XgvZtThgajkYnGFM7ogAiFJgo6dix5/TCTPYWNesjCGw3szzll0T8V+xuspa
1DfMdv7fszD9Y6eRwIAj5QoKjw/JU9JkLGgFUJqzPnQqjWInBdcDXjPYwb1g
N+yK7c5O+uHBhMS21u0Fft4JxoEyskDfOpTN2WB5cltP03ka0oEtpu270O41
06AUj49Y4neRZf0xEZOYKIkN3LC09GnmnXmRajr489/aTF+mDRaQDn8CAATk
9MdOZDWTtzeeM+iFQyYaMxvL2SwXGzJquKpy/594GKjSWL/v9gonuxZXwGyp
kKZL1KWhmeQFuyYrqwYmSR7k2g2hp/YIdJAnWbgqY4hNCVoxKYkf+4k/1D6q
VaY6rKRUmNskt2RjieNmCoZ9r5ZYbrPT/WHaNwpetPPNMGGztzQly2cywRJK
QDv6SzXri1sZY7SbIVlq+2xw+gcB70xqIw9GvLAQOi0E6bsTHn+h5npN0fcI
nl9iK8ts39rtzmCq9XNa1E/5rgh8JeXYSLZCY6LkPzNo8+FEjWQJQ3d82QKJ
9JGw7OQsheLvBZm+xr8MGwpVakQNeOMAaPogd9RN7EuwtGARm/R++JYyZc00
X/kzKbxVA1OHKAkti5iDKIVMorUlIa6h8R2IYUD0DglDNfMylXn6CrUE4lCH
zzxC2P1iYue5y+HX5N0s/RmXjl0JVbYcIvZ8aFkC3wcnlCy2zvXPepga+wMz
GMVEmvp4GsfxsCsFzckicDqo0jDZ9fG6ITQakIC4nSzJl/0tjYMV1DQoNlOI
LT7O7oZsuK4o5QaZy7JXemjiaFoMCr4b0l0Sxy7Ub2JVwyzOaueSPf+Q/++D
/vaJJu1dC212UWEPAhSHG+FKgTRF37Vz5ohCR5ZCIlATts5qRB3cJE+Fkra2
iyU+oWdlAWea+9VSFpldKy41hAT4gXfOREmNf/aj3y1AWmRIdFKDO37QBAnO
2NKTiLlWYvO9MPXW8R/Fw1t8IVl5c+/5e78btpVJH7MGbwp8uFKbaWcasCSL
qNF7+6g7T164RSQMzWISVzuaaqjWy7wEfiiOikO2ovMUABZW0jXI6CIAKmiP
Qqs81GwQbYwM04gpnxWtfiGm1RxsEYjCwA6eeobgcbOeLQr5khGBRnPeMpap
EgQojxlvEieZ8A2/6vVQR/HpY1cHKC/oe0vmTl1YiSEpKd1BoMLQQ+zn3++4
2WLqCeX/eBxlk912gjXX6UPh6fa2eLgXIrZz0dSWY0LZfN7rwMLHH3UZUmdr
SC3P2hphJo7gbOl+RZOLdRdGdROE+1xzHVz9YFGbwJYhK5Db/ySy3BJnzB8m
RcLj7uGupLg/NEDyaaOUORNnWwO5a5+fh/AuY7Wi+7tpAF/tJnDedZIggWUQ
TUlxRW+ThKOifwnf6QL6HklF4MNp053DhKNQWFoLj4Anlb9rosFUp35urLWy
tCO6vV07fYJF9bobmcF/wrpuH6lds6mI6ds2QvB/JBOQ6Ml2L6P5GbH8SJeR
ytJvpFdrUoOCakXTZFy9GpkgxlI/fnKJaVYHsKH6K3FTTCN0eyOq3eb49Tb7
r+V1eNs+bXGR9GYllpSgbFNIX70nS5m0lBUJmjBJon2QELBB5mpC5z0lgtzE
ud702r6y5CmqyCUO6lIYGvvu/4XKyjU8km1cluK1FNvOZMIqTE9sskxdqu6D
O0Yx07HRGZ6C7omugmsp3J7SBXMfIXaJGWN4EJo6KrqEMCF9LeOcUuCEBtC+
qtxMTtf3CAqomHmK3uBjLqTSDUzd9IFUVRRf6PS7Jw1ouNuUxhh0c41ThFs8
s8tvEz7hv9cEkVsmhcqPwVNGPaN6YyuggOIJGE235J2ijPhX6QgMw+R3V1kN
nM6soHhGT3M8JtJcLYl1FWDd8+V+65TQ1+B74LWn0a4R/dl96e2Sf1ML0Yl2
bsv0f82dPEbuQZxIV4ZZFnybyRyYFLE6w+vrwNDNBFji+4LHtG9uWdVeO49k
7H0SJaotO1c6E7CyAK1CDaY2n39wl4tyXTyGWxJt6D6rhIUiRNaRkoI0lYkG
DGDOi4CpDsHUc0emRhCt6SH8X3v8X7Br8mvt3BFOBtvFFWswl9v+Qia+KlxG
5iPa4Vz6Kbc/TrP8U6Tb6CIqGjh2prCzCK+zgxd645psqXcMRIfbZlc0pnZ+
3Hj/P/PGhlDHh600f0KdVf4T6xz7B+INtLSsuHAKNZ1bHy3mjik5d3V0IwBG
lP+ev1GZdbnSAAt7G+4YjKCEp0skYBarWRbdhyoooVYfeQq/kgZlfsyK5BNg
8cB6bS7jWIMveVI8gBpFeAZuXF5ip95NobSxFgkyZCZnKbCXtdH4sO1SeVGE
vd9YVBrc5LSGFKaZCiQukge0p7xympuinJmXnoLUf3b9zfKdGlrnsSd7dYUy
XqCYyMkosRBPTb5NdPrVuaPTsfg9pXmFJKH+7jHBVNgEFdo8zwA6g2e6Ad2p
Igg7G4DZDwMhk30uNJBJvme1LqaRFUr6xQqT5w/kiEAbTAJIJ4OGYrrY06Wh
hwR2TgJxnAyjuowdNTwhpo0X1EaALEzONz4K5h6Cy2oHrMh8XFKhbYKBySTy
YqOMGmPFJZWVL4UC5rp7mIzEZiqhr245pxADpZQRMgwE3CSWoelDk+vyxpRC
yLIDmTbipt+YyIg7KKiHWtJ4JAiqSyuLFF+dnrkV5ae3tb3JBVZ9/30osQfJ
sT0EB2udnA5ZFTZYiBKgRy6oUcKJT3/5NHW0fyTok8kQoI7y/h/z2IDaQVye
D1mx01sLSI/HpMZkp8EtiKOPb72AkxbKbufzux3e0AEsOaXQGKFVVlgTo2zu
1LkA55ZEvZBK7SZTyHtuSXUhBkXEMkIXMQX2psOfDp6y5GxJkQ/8iDAqdyBG
hrxihwtx4dq10s5IjXq5NouH1sag9gAcKdqG+O7gsq+5RwdBZ+QC7yjHyNDE
rv95jabxqw4M5q84pW34SuzVgZMjYFdiSMPbhvQ1Rn1qWO1NAJd3D/o9zZ2V
7VJrRL7XRLxGrhSn8zP8nMe3eYr/vqWXlzdXC6usp/Q9Mb2BWqSCkU4jkgjt
rb6M4xXNfy3ob1mJSvoFWCzEO/67q/f2uCk76fDCksfASt8yHEt6+sySPxva
ebezJK5BCPRktLwoe5m/FCFbJiv9Xkbe7Pslf+Kh36kalIyVkly5P0yH1ASA
CwRbWpDqAkr/NSIC+phdXfMzmZiqtymBG00wW854nImhm1/VO54TMYXCo5J5
8rY0iSyos0rYyelXLowE21Kj6qtaDd0hXS41IaJMtG6N008wdjd6Jc0l5e4D
9xG51Tm3+rz3BVql9sxVvoE+fQgsXBm/OVXRHSInO99Vj9WTt2904NctEfp1
jFI4SHaISc2LS4THoUPrLkCPxi6IcSyNRxOGo4iO4pYa0w7WCl8NMN1Y4mzf
u1ioM8jqRNV4Eu1IGQx3oPlQSoB6eF07SAnyHOncFUkgNgUntuA9Tc5vxPAd
o2+U/KfFvbfz7r1I0MujMFNbDCvJ4l15KcwSy0S75eByJSI+t0tGWKvbSWHX
lqeouBZskQLk+Ow7gIoC1hQzW1HPPn7mSDKK7Ldl1xu588PVlOd5NTVAMGJv
DTHT0RB7+kyX5jfDs17OTfAkcEEPK7J0jWYvMXzW2XZEPzkcPHnm+jJLOZb7
CUQ2LbMrj8IB51rmmbnLrOJsLwDlTj+Enpox1V3pagToBkcGqtJOI8uvvODo
e7QSe5M7z5jeowxhJN+Tr3DHD6dz+IGcmxS+FsJsov0ccwf3md1aaazqPE6V
P7hwuI9K+UWCoQYynJlR5TDqyrFajN8fV5znmgOe8NDxi8CD1Ecr1cpAcin0
mTtayicHvt5nvzq8aOWVnlci80fta84b0/DDvzC+05BrQKT5T4ou6sikqlvR
VNGKM+NE73CDixNWOkHMLyukPh1I7BZI7usYcZc3jYDDfkQgE67ipLENG3+5
2gFRH0Jn8iN+LtPB5l3Tna7dlY7W1/j6oAAHaKfSG1yf17A8vSyHsnDu/CTx
QOd+87NAGhAhWua4fr45rGnH5E07STqK7Df6laZt+Jnx7p+h6KEL4uXqrW1/
+3RpXN62E/gswfl3dKbBVdmKDZzHr3ckZ3n9RA7YKK0qUze5IOAjhgAly+Gj
cTk1IorsE6YltpyRpsUMHy898wvU2u0Lr47zR6QUqzWbsuKzNHFsl0Pli7ge
31wexuewhfjLBLu5HFH32PDlpqtQXH4qufMsfRjoI/iVhli+uPN5hmxlQnX0
rDT1oOyivFtu14D1/yH0ceNfU6nqXpFF3Z5e3uElZnjY9UWgK2T5tMX7MWlO
PM/W2VYWExpnSDTqgPxHLM9RUawLTlNYRukft+3710UsvHATxP/iqsTTw85P
8WCHIchHU0WIjtCZOMxI4yS3eKHBKmIRoNWVR0azQkzBQil6S3RruA2mEWuS
0xOm/1MZVlFH4s8j7I/5CzUc1lRxm6G53Wsob9F09d/M81npPC2EfuHebCIc
VOUCuXUUsXSsmu+ZkuWC30Ueokp1FDEUxusnSV2Jc4+zofvLMY7SBpJA59IP
lYXeB8hyfBfkGaEW2JYKGZErkRAaDxC75ACG7eO7q2lwSO1iwOcARHu+hDpZ
OUrybY91dAAN05duqPuLa2IyPiura3FwyFbvvxRXZ/lEUasRSzViVRPR3fk+
jr8h8H4YqekNTqU63D/UuDW6DUoDWDrqsijbHp1nAHc4kpMJ8qrHpl0LaSJ6
JwYxCQMOQXakeDdsj7JGbx662rSkzBoTaC+zDvvbKt9iO8uftQg1r6Iq+ePL
qvQ5LOdLDvr1cfKhHK+wix3jI6Zchg8/1LWvFR06ngSsdNIE2771x1AKUORk
hiF4a0XzcRua/tcUeQrDQPZRv+bigOz/lztPawpstR3WOtoXiDlaT7BRecmn
0iUgjMX1N+3OcfwO63HQ+yJKaYK4MciWb1qF/n876XSFNEsaMBmk5sG6HHDO
FscQ+Ewo+VBm0s2dEvJLtfl7WaBMibgl6qaHhjI+JHkcPTr/ZmVOMA1ycLbg
Sl8cGRKW/nsIkaDPUirDdG+H8+I9jQku/X+ucAFDZF8Pj/PwQZWAPF/6ajXS
GlTuwmV8MnrT3tUzk7WB/rzDwRt+SIfbxPMCz11dhwRvm7/Alglh4giWpJ0r
MKAxiuGPjtcds8+AoVt+qwbJ6kinBWCrM6qxMecdgjbSDhhvw8VXn+hg0mal
49j2/awg6KM0HYHjrxItjdZKPxhSJohWjqTrxUqKp4uvx5DqrZBD6dxDNzAS
0wVLYHqBsXJpjqMk8WP/FnP2FCdv1iWW4MHOgt3Q75MfgP/dsjKOqEn1wA5R
rgkofFiHXtS/SLCNWxm/EZCPex0WF0TzvHJ3KUpgGy9dv3p92m5N+ztrNmML
lxV3tDkxhN7/9f9vCgqWbMcZSoqTHtOKTTiLhJEJwQECw02p/r3tyezUPkE5
rXk4P3Khoqk4nq8cqWqD4fyHpd/+5dhb1zEXOUZyfoXcKgxS4VjNHlehzJk8
u+iU+lpEjrIf7a0YNUmA1Coa3XxaD9YMzhWhKWLwJTpgIdxpRcjMBuB9BHjE
Ae6Szk8HX+6N5i7q1X6SAQaggGSMU8fQQm21wO9IVvO/dWEm2kE61Kn9zB8O
P4lpECiS1mPbGHNO+OV59osgBx25NtAJj1q/qDbjm/kPnvkoX4KoQ6lermkH
LSShksXVRSdr/F2Qp9X1HeUnj/W3NiYXVysBoCtX8hT758n22JjvdpphcKRf
eHNvhvbkkKKkfOwsqxq3E0mdnRynKBX+/pdpCgine78oQoZ28YbODo++UC2o
D98Aa8yd8ex5/t43j9pmymJXqAwKUx4b8wqh3yfEla4O8M8v3YMMvkobWLUd
jTl/TNVtN/bfcKkIizoij+LhQfZydWcFxAmKseDhkIz7yqgt5ynSUQtw/re1
yI6saaFQ3ZH3tuWdvTwT2Rr5CBN37h0u8Z8k5l7u8VVK0XFMrvFEJMZxepP4
+5mTn+VIBM+ujaCl5x1R3ox2sD+v7wMzKhwSmZbLtwW2/lnzpGydpdnkZPMO
ZmxyvjNz6L2cXwfdk1p38qSKuwUcCMLEGktTbL9SJdYvhMHjh3pzPj0BPuYF
gNncpvLXcHInLmqcLdzL4ZM1mhBMS+N8kP7Otm18CmAHG/cJMQEeQ9UPl/q1
8PHu2PT84hO8P29xKHESckEDraqRc+tWFfnlDw2UKYMPOry6gwsrupvE+Tu0
qD8m0+gTraE1C+86lequcmGPg7IzoJefq65n3ieTeVE3btzsvB0+OuzE3O5y
zpUSRAH7akg0L8x2kL57Y0/8/6iYlGdPwvBTTqLzt2ipsCOW4pVq5KriL81m
yyj29de+mEjt3oBkhBYGhPszy3VouAOn/CCh4ii+R5sTEMo1yQbVNMP9fxY3
YMQP/EvDq7+N/OlibG/IvgW173PGlGuFjzk1jbgSzO7udCqi96HIiDYh87Sp
yuYn1kJ6dAAQnlmbGCjQm56G0fpKG4lXmXoCGC2tGZ5OcxZuVZD2TIJ5NGHt
NSDm/DwJga57VYXyXOWeXMjQgosEmAadk/uY23Qm3lugAcs5OgIxIuu8q8Zg
aJ2K8uY5HzZGGZBovjQKET2r3ROLoDnsoQxrkTHG8VaYYEYkyrYXGsTpAG08
Qrze0emFqmjUFOGW5r3FbjL/HJOaHt5nu+y/WxqY6dGkngKxDE/TqcdfDpkZ
lvKvV3IBK7CWDlgqjxi4UXkVEWdVDsriPBRaVno0zXe8YXUTQmxWhp5itzZy
sKvRHOkBh5GzCaEac0twrWp4LelnY12Kb3UkVUQN2tKjzaEakTrXOgJxVN7v
ZoF4lG7n/Yz8MEt+zKdTq1D/mzxLgCV17693vr+vEIBFsx+tLabklu/xtwVl
R69xl/9Et1G/4QCP1WXNYmjf0ahPBfFTAvNsSXIqBvidcICmFORQUcPXFDTM
VDZBClWAb7c7HA5npDKy3/W9OrWzx09nR9XoysqhW+3h+I71SMZRxawlB49U
a66NclBXhvDB75wuaLpJOV25bm6FP8NzT8Wa8iuG5YCs7Xhh31XaPWB8/ss8
c+TLUa3D7RM5y9G8nzQ39YdfWWyuAJu4ZcWjrL5OvdueCpQGtpthQPSOMjvQ
RUTuFdKwFGmBXdCOOT5eZJ3afwUMIEH5/TFgRbveSM9hrcK+U7u1vuju2cQD
HOhRunlYMIg54LwtmBY2jOybRlE9ZZjV/iXH6GnF2pd7MrEXxtxUDQNd9eAa
mDan7A02khSCF2tL+1iiu37ItiYvr5FDHK2LZYcEVByP/bW+8D2MapszODsx
8IPB99rx5peWgJXmGqRt6NlGDXUS0SP+Wqt7yLOT2p91BRB0KwgfW7zC8HgV
zbzMotlb3YjxChfzCbLvj8GpeWgO3At7WowBkWy3Uuv0rvfCP9SiuRoo6WBn
pSh2k9tBNwfyP4tN27bQmelcTGh4WATNvpyXIPVmPVibOdyPFX6rLlptwxEF
wmChX1j3+dSIk1q9jgzJmJuN6p6H3RvVhkdvJ5VMjuLEzRhGM/KpHln6veBo
eE0P/hznxzLmWUa6cYF8jC9bDPGgaLwbasZxjyQdv/xAlHWBJqz5zXtw0IS0
QB6RMe10QVAjO4oFF3wTipmR7kUN2QXfYRDTfX3eFYM0SqwvqDXd3fIH/tGc
qaLwWspeza+Kd8P/NfAmI2JCgcJ5GzV8VCcpPE3Maei66WxSRcXr/A+H0+BG
qEyTpJSlRIMoySQe+2v5Xh+MSxxLtkS3z/xzd728Vp9q3F51jQUFSVgjpU02
y9m20I1LYDSIn/z40Y1rHDZihsy8mKNVUkKGM67ylWv2wxmaeYNMvV5EtIQQ
bggiOVJQGU4HNPMFGHvGDM3s8Hgda2apKC8R1Vtec42nMfUqIQcLMSuq9HdM
4xJ64XsBLWV4/4Vow/e9gC75v6iJQstiRHbwO1eR2alEMDQFpxkZInRghT2l
bTFDaWy3NTFmis0LGer/ZTg437e/w8FTdfOFsF8gzlgxkRBBS5FTKcYFwn8J
P3lVzmSV6ItStvFhpYT4gPvnd9nj0bfb4B+PcvOldckACXlaUUQFIxitxPjr
Zrs5onVBC/jy6unN97aCzBOR1by01Bxc6lhb/4tpUc9h2cRAHFUXiqHQRnAT
FuiF82OnI+i0AegxU5adOx5w61gUANVyVAFONi7ORqn9wKMmEa6h85G09n53
MyAnxg+5k52v1gWwg5pl431OATZfOWEfLYbQp7EEapkpdIiD37qCq4OLVdN9
Y1gTGYGUZ2hqb63EDeNIqzB14gYEPbTJpLGkksif5llRbrQ9uBIsbJFdw79Z
Kpfj07H6DdkoTxmd6YQtA5N8APSwpOGhbi5ZE3Y+UrsJoFsM1cUYqTzh9Yet
b+9CfK0aP2GMzCadYmQ7goOY2e8V0AW8QO8b7HLTS47Kvbk+x5gvwVhqdgGE
z86DyrDIe75H1B8pOdcTu0XHt1KbpRnXj3et/dckniwIxOPiEnnstICke0cJ
9n8cywRtoytyF5WV0bU/26ptJiOanP9+1v1o4xH9oC67JYK0RQNJHnNguM+W
KF2oYv2Aq0QOtE0KFCB5+BQ+bOpU3vBOx0keLkhKo2ZlJtz0VQ96ZnXPsfhQ
RXpQHlqXjGUqh06Dbr3Io0KoU/p8A2NAXxukxlcvAJO618/1VEOpXaUrVBjj
KqTSjhSZihWyj3GyhywW001jQNkVWz7Qt7L94HOSB5BnHKWbeWuf1GNauB52
oM+FujLe11+mmddCYZbZ6Cm+GujqSmDya5OYX1Zl0YeOBVPOKlB2nJQvBSN7
wbbuEN2tmOjWPIhBUnUzj5k64nc171W1PcAFjw01MEhSD7rvyXweintJ6aGG
PRXZ5+0yP61Dwe37nb09MWETDBV8V9AYlgN8VwPnjR+/569fe/iOG9sioJoO
rBwKXNOXGA+cwHvFTVn81RDsxkmO701ANG74HMIAk/Q8TyL0I1cv2s5o9Ev9
BGlYsyhNKvRWXTKMZ2e2f5lKTmCZOPmbNQl/oycWXiVt15CSbQhLHZ8J+Wi2
sr8JarzRwjD/sKWt6xjQ81957912Fpqd01mf5bDCUZf9EKpSP3p4V++IWmxj
Kcs7i0B0T27Ja57MpdHOAHCiAp+dkKjyzqTChxs9RV4jdYshmOgaA1dRtV0x
ZXGAIdQMukEzNcEMr8jcLkvhpXAehGzlx+VPVlAfr4lpgMcKOh+B6XMWdEH8
y/K4Y+Qi18Cb1CDWwPYfh5ykZQtNS2hE/t7hSFIhf/b8GWKNeXAtfAwn4Xpw
3cn2DFV3o1RFvPbDWXUImumChaKqRQ9IwApPmfUy39bkJJWPDPMmoII397I8
IBpIInSZAzUg8DDaWMFaoUBhQGjDouo4T5OQkAydjt2YK0m805W7tobozbS4
AEQkywCclT8G0s0JcrV+siw2NqQEL3gOEwzSUmHPOqMwSTXfIPOa6W46/DYQ
hNcWLKHps/osi0B3z8uoxEWCEn4gQh56oTH+fg/WqqpmibssYTrfsW0Hfok+
S+zbluZGYac8rK7ygO8Qx4L43j9kJ2X3buGRZAWrzBMJM7zJobuRe/vhzBUN
TXfHDquA58c+eABiobINBxdWn2VcgYzdqhw7UBCL0qVBOXRaLyOLQMNxcXTS
H5HFsnzEJUl2o78dx4Wi3dLCXAtsfQII4RuTFDuT5vWm3/NrdwBSn/gNxcfk
koDNYfkWMWLzOzfo9b65ztwTT1l8G0AnWENx1B9eRYQeX44mn8zsgC63sfzf
KTrRioeY+GP2lcu8UEbsKO0pwI3GB3W7hWsGc0wauZ8LJn12FyhR0s5J4wM4
nqluRpE4HJ4D7DKcPU3nEyEDDdvHnpZtEmGWs9QNR8GadPPEpsPOnILq95x1
T72fZgnH4PDWbc6FLyP46gzEoqEbXLCXdlbVHKfswh7JsCQ6Ib48XcvDlMKP
o/SNjNZBtsELcyFv5c0wBfQUmWsUaaVGNObvOnHQYnXs9ntftptOU4pSQO1U
P83m2t7C8ULNU+VYXVEZPaDXIxL2R9YWkeJxYE603TYQgysV/vg+GZYVyZOf
rO81MMNzA6cMKOKsoj943K6OYRyoz21LaP7JX4LRCIlcFE3UTN5pIKM4zU5i
m0OCWDH26owHJGe2zHJe7btaW4vBIoAECg3QY2+UfMb1rLO5NuJsDMWs7VBy
t9aX4aOaRZi2TW+e0sT9qIidITexfW55VS61wgxggqt8JXic/Ux89eDaniiQ
M1tm8QZIpBQqJjMJY/ES6vttjhQa8h0x7wRDvhWbGv7iRmbnoiENeIDn9YF8
YE0KeYVzcLaF8jwwkzer3X1f9f3zVBOuc0+Q4nZhHBKgBqj5q92pfJcOWnUc
WXP6BN3ZWh6MUEjqc9qjyqfe/NM2RpDZN9Oa5VLBDS7u7P60MG5Nls/XlOPX
Sr6eRGnmOWS5JBf19LOocddybwOEditq/Qdv809O+w6i6rrfpZMlCGa2UOC1
hVCc2nyCxNwt2aoaXrG6Pb93XzZ266aYIMjsVRR5sHnU7y0vFdeowMTQRzVi
Eupz3QRSDbTI8to7cBNGFi6nONWuaAPR+rqAtc7SHGm3BpwQOdwmZUz5P51B
5fEXItS1DWLbpiI83aB6CbaXzCyj7G4/48rhSa4RiLf3yzFkeDkrysJyX/CG
lUXoqJgdWNUQYM7v5mq/6Z8tsQkXzcG8RxrMovYom90wZJdkQlCX0EWkQCmo
v7VnW0pyw206/0XvCw8gDGO6OsNAuAAakHA+sr9czI3r3GGGSN31V1iD0Iah
+G6LcbBhHdfWyLrqEnVzzWHZjcA3nnIKWKNBqAqGpJiHbJwUT5dlPPNdJRa2
ZyjobcDCbFIdqBx26H21jbZJsO1hL3OFx4Ex3D69FI3QycBJRe+WFRzd+nMv
c5zVAzTZXfdGpcQvglMCd2UTEXPtRSSyqcFm42b9/5KR/AyJthL4cfHGy+fW
n/A2j2loyg0TlKnRwLBq5sWNINnugAuNKSjOPlmr+pE26VocOE7zIefROOqi
ynDSe3f3r1CbtBBqmU2QkqPDXhNKCnFghNDfTKTvdW0NuMeaT8UDAZxVtzYb
BH9Szcinp8sW/TiaKEpObO+vBfqnQSOp+0ETkUEVsPlZhoSeHNJpExWyr1EE
nsJbaVB/RAhCGwU7+MMAiI++9w3TTgysRyIH5sg6NxDlQGbOra9RgnYCKE0B
DkYUpo1KNvgUNVCW6ZVDoEBrgcOaBV/QoIudnxGGZNijCucu7ZET6pL9FW8u
XkkutrSmJa2bent0zT7B9INEeM3yBdu/Zi/lu8lhMdVU72MsYSP6EOlXNcBA
fR4CE7YGf6IqyIwbcnv5gdM5OECzAZJNO99swYdNioigMCSsMQHS7tXJiKx4
0PYpn3rw5DE6S8z/dNL94lAKyStajrH/GQmZ9lmYaAMmnhH+x0KvHvinPz5f
OIs1RhkFimSvE5OXYLPgVoyblCB0kfl63i0LuHEe1RLst+MbyLAx58460vZr
HtqRWhVqYIdu/MdtSzTFrY6BAHQaTZ5UawwoRN7hwI/PineUM24Ob5qsMOvb
J64qZFzIYgjwH8H4PZXBBDRBiy8B+SPAowcM34W3nUjou6OZiksVIxc64YWx
ysswM8L72ceVzKGwDZrzW/tlhA53YXfd1dEbJk323qXTDrWv7ywyvGezSJcg
Dz2xgheaC9voPy+OZ43jtmVrev16MR2s+iILMgmNGNrQxr689E1CO+XsYCE1
ECKimTSr7+ekPvpxLSeJBQqHL+MsOTicl/SN+ALvh6hZCHha5UFg8pwFr196
Ist3MNtl9lsfZxyk0Iqs1HqQ4Aw50ZHmm7WK2BpVw4sgkRSyZ7L5mcw7iANx
hdF5jDpG0l3RfTAunACOEhaNSj1NZf51HkKhNuUM+o9SzPQjZk0NEqdvwJ6h
ttpm1qU2IdJy+GG4Xht+cNoiZAS9t2wwNaUG8dF1Z3MGsJj+HaLvhFr6yqsL
37MwRmKAEafk0jdOyix2q6z+inkA+Nu/eL0g7t3cSgOxUTObyp3lP7oBFXoK
WYAt+dtL4uRKex9evmQxK0T/YXTvhhN60qIEUW7ECf9pF3rGWBPTa1iwp0ba
04rqNkRXK+Lhp5vWBOKdVq3wGK+rW4aH7nAa8J2ZbPIMAm4+JUcpmMTmpjH2
vZa3IHPKm3/VcliooJQX16FrsEV3Sj7hqxQd1DZAVaTBKPjorwKEcVz5Hc1c
kOgXDl3RI12AkK+iTSqtsAipFYG5DxHux65yUrdf7fRCRQAnMelgcBMGrm2p
Sg+dfArA+/MRuobAyMf05QUudA/LZRs6PKecXCpg+SMXnpLyEEBN2tNJ10NE
gJ8MbjE9sTfTVo+4mX8JRc9MRrBGS6ya+XvICkeBGaXAPFNUXiIFGGqmS/9t
y3Uh3r7Ntx62aSfPglL7SsrewYmwmDgt9HbrUJePy9aBNKUhNG99W7yLj74x
4fUKCvY7YlMBZMoMOWNYyNVINLrQOIZGQ9B1iayqkEl0CEq2xR5eq21NHjdN
lj/SO4kTZ22AJoY/O8p5kim754EmQx63AfVg6uirjA925rmA7dDkUP4skMAm
fvj6C0ZhNRtacGBgATKPbtuW3PMQaARd0NlgsuNRsMR0oboG0kF1di79V+h7
yxLSyqQ2MckEkuiMQCnRjgcA+IbB5NH5lWSBektXih+giVOjgF7M7+esek8j
zqQyldEeYBN3gq78+ROlddk4jzOdOgJhgcQCVlnGtO5Sq7crmznDGetC8Aln
sIGUvW85UKmfjLeLvvPf4RPRCjAg9a5ZcGg5RLIc2O522jZtaKVC1hsIyAoC
P7VWvK1GR3M7/RXb8BcPc2UryLtiPJAd3JO48kqSIvUjzaO5VZlMkX7vsFrK
yr3CiAPf3jl5Fu2Qp+RA2IaQP+QVLfQVn+BybWL6ajWx1oJykUkKH5b4Qqck
ByT0Rq/sZwOTat/5RC26XBVICUEUDrVa6vLmDjxEfaZ1GlWF6apBdvLVmr5L
IH+2GCEX8+/hZR9N2E1QKMCgG2gCiLo9W8sYHiLisUmD3EsY+VbUS++DZlhm
vsVBCH3erOt+IS9M56/Io8SBOu12rvnBq9ZfPgHFpeyJl+w00jCsu9dL49KK
Ix3tAMgeRMULqaMQvmIfTv6J9YbmToLN8dF6tQ1QicETl2UbhKw0d7sKXzal
fxmtUYFUIKA4uolX5kmmFVSKb86li7XAUAaKzDvGe+kBgfgKhSrjVJ8ZHCzB
pNvs4N0zmlebLlsuxXAGlviPTmospY2wNEe5TPG4nAqs0CeMmlHWh0Jppkt6
+Gw9hBQ6OcW67uTWnCm5Yl5CuZF+4/FSxsddk9OLOhz0wbbr1WBldMDhTyKL
CKBqCIVeaaI6lTUNHMCzihOtFBgW8UaBNK7AC59YSMMDnwQy21XSto306tjx
Jo/61BANcX5mRqkHIC4y+NWlQXwBc/5yqLA1mrMXRfwRwRMGootVmXMRa4+N
/3VGniHPxWc/bpcNXycnHWfnttC9HCite+OQFttpe8KphJkRFZiIkGmEvlio
xdnX6CVg11aH2e66X27bT+OdZBlGyxZAmItEd1Pv/t+6bYEU2tYpbEQdLLcZ
onDaySAopNtK6jOuKFlZoZcFG/aJxIUnHtG49cBJswIADQ2loomQb/o7g/yP
Lho4yue55SnMAXtQvj8Sg12qHbIZn+kUDcqTwUnabWpNio8avAxhi6idJusv
zJ9sZHIjn0OSxzhLNgKw/q8ZQmkEmSeIDTDLWp4Hv2IZfNXM0XJLaUrGjMal
0byVSuvvGPufT7tETUQJdtLbtw0EfR4b8Z2zdLdHFr5BwtAbrdN0TZOdG3s1
vCubmj/0MX8zkSg1YfObpDI9+qP+uZd8RFpisr7fy51gzPG8nkGOtGIi4SOw
HXE/ubGzYN/JEXcL6GhfL8DjT79GjAkqJzzLBSiWTJ/Ot6mlGJ1ns4YOLuoy
zSBAnJNGBdTXLpJXAp7rRc4+VqO3GFH5zVRMyn/kyWIGRGUljyevcEbxyr33
f2BXkLEqZlGSo2gbsx41Z596CR7Vdp2Oaz6a8H2ktrHuJx4EjuVDvh5pL63a
BE4u8kv+ipx4WzqaKxenTmogD+P1TBVreTqxtclW4sRHTx77pe/l0AOHZsq7
yYaeonn1Hjp4PSj/h+RE4/2CTg0UP8nPg9FFfWqfDCxIGqgqiMaDxnC1ZPqr
K6nbOs6R8c1cxlTpSUcIdYt/IMOiWUpPMx8qHqebApDOLmdFpiK1XaAzP2Q5
+JSNAwWu+ttL0uUfg7TsrwCfie6fL8XnbUMJJvji50esq6lYNx1X0rmlGCJH
72rYVOe/099deM5Ckl8lhHwXZBt3JVAl9TRfjJ/Oe/5rYEFzeT2RuemqzyWb
pe+AWZwX1hU4mEndwGGTgzbX7n3x3dtUkdccSJeK5JoKHt1OnGbtWx1BK52u
wwNr/buHWpX96Z1zIoGTdR1TZSE27ozfl6nKpOuTVb+2Rr14BMA9PTNOmK83
EieW1A2pnzDIBTpXO4DblEGpmWd1MR8tv9BAYCHtqGpGVxxcQJmIXIPguuVd
erl/M4D/Di5+TbhStfb4bxDHTSLRSTyO4WcV5qBFriOhwqp5dNLspXf2+UfU
U64g5eo5Z5SQ9Ix8Jq6VnsYttF1TB6WB4xmLNtpktYidA7zisgS77Olphk9l
go/EOis7eg5cTp3AWP0F8bz+r4kWrjFMfkJYj6pyOiD4qVHuR5gMs1SQ7nU7
49Gkf0tC26GxaB/BEmQK9Qqh1cYqAqhpYU9j0fHArBSDYmmARfVnY4u+XdyM
+9XiQdDLnIT8kUD0JLLTvfBI5fVvIRZghKZngoqi9Ldlr2LygrV4YHJZNWh5
ZM5mGqMIiFuK4vp1MaeE6BKZZ/0oHWzRBVc+ixBUlWCZLuIBs5a8sqIo9mn8
M6eDV31rB9gjbMgY0fb3d/sIKf8tu0ONZ1XMA944BH8V/fLtjZ9OYG0D6BJ1
gFeCB0uhNeS4qMhbTSFzoGG7FcOJbmbrTFDq8lBMiDik+dm5+JnXl+AT39Ch
QaIWcU//3iPnysHcfnECQcTnFckM04fVpeZlpAI+sbf0hicfOnk6tOoj09sg
OlyORqdUbtUOiUGgFDQCjMEK4OVtBduxz10s6Xk8DhPdU0P83xrHy3wkEFS2
ItQ+qIXjPtKI593OP8YxhBaJLPTIS+O8/H1sVhLtAG/hn5Cmf8w3pG4plQON
mVVNZ3D63NZOFKc2PMWgzb9YXFaHiasIr9PthcTAIObBhUWEm04OL9f9prV5
669s0TZKJgDausIRiX9AfeH7t93IqARFH6f9jdKTF4DOCUZpQWAeQyvXy5Oz
UPpV4xY2dX0v+84XLaU4g5AfTZZriQzYb0FgZuBNq4CAzkyEInfnkEdgH85p
NujS3Hf8bJz1okKZ32540/F2gx/Je6ktHK5ZIZyE1WEhQLTN6D6i6pHL/nU+
VWmShFeXWT55EJqORujEjhqfO+AKwOE5iBq0lFSxP9g9y2mlh4SXRRQAQyfS
wmryJ6N5fRRrwz9AZ25nxvoFpBxQgZHMo8CliAlq7ZPIr3kiC9NStLTSIVMP
102vwbttBpP4NR2KIOmaHYf4sSyE2G6seekI1v0qptTL7brRLuAW4yU00fNQ
gqbHXGa4Rkaf7Puty7nS+XJHgx02tysqoWCLbhnkUGPNpCRBISypgXWMSbGc
kq6H+k4HU1ChRHjsDW8yAwjn86CBebbt/z2BMAkvRX6LLuBWblJtPim1Gc/M
KTh7owTDLqtWSj+V63UIpIh57SiBKGyVFznAkRamMPGE4t4CZ3WbwJp7MqHM
Q1crHCP5CaajMe3EGraf3F9FsD3Pj0imaHw3THYRpjAZCovKAREml0HMIdLz
RmXx3kEYvvOv9yU9giUtf8sRbJL3p8VZpfvhvhkPgG5fgG7bzLymCcRzOLLB
ODK/1NBSzEyYiB7OIE7LfUYlONNRRZEcCeob7uXI6KnddUhOtiguJyHFMBW3
YZ0JGibNCYVJgY7t8Ukod8Kg3e0sLNZffYP0Sn9X4ahA71bP2wzqKNL/byPB
0rHpvgjJt0CpV61gx5cURf9qEcltZ/XciSnw+ZzBEhtDd9xzn3Jzgt64ldkA
38J/t+JEBBq9QfgYeir2DTkhLEXQ+SG1NmJSKGXZ2ZF3vRFV/GFiZGaievjk
N9UFvqgfsxTEL5brkSGOv5pRC5Y/vovhVZAXyHaKidST0fywwiEoP4l9KuMz
nanqH/n1Qroo23QRnc6uIu89lbjfndbTqtrxpP0ZzKI42oZSgfjICTlYanVx
38MqaDQBxi5hx+o8xMJpLmTSK9/4UF4NIRMhsfvGrM5zukDF3JfDOG0SgVqf
AjJBUjECoTK2PesAdRN1Tp/fhsCqqDhBJ57Y3IiY9ghjKPcIihYQTM7/9GZw
EODfmBsWh1VpJcr7kxQ5Aly+OrpZoQvJWqKR6m/TXg7StKtv20M90PvfhrJJ
aLn1lWXkGmrVSOaNYrhPJsY1LoAG0K4JTnPhlxSdb38kzXp8/qmCOqnvnv7g
3ATrsLTYpEy4XvTnEP9kREzUyV2BpWd88TEh5pTQ2fxbgsnE76/KaAEYF+a8
eRW89y9N1qPFkk7zsvb1w5l8LTpST1edFdH+iHYLknwPmkqlcjR//KbN2UhV
nJ+q+GrbIy4U2Pb50yKkZi0BSp9zPZT0UVD+WyopQe705wbfTKVh+YkQnNqL
ADyRYjZXbIYyWqRWm5wk4fVha1p1lu+zSuUT3LMzZdLfppeHvrPdPaK1JNQn
7KQ4aOph/XKbDVUIQcFJ4N6PWzhZWvkVjgmXRBlN8gVJKbHX+eGqQjJdmXon
3AVtQSeM21OFBsVNqQgh2djeIA2gZeCuZJrW2tJTXtQKmgv5f2URO8L52WfL
8lQTGk3qH5sPPWLgax5VOWAI3QyCQIzsaAT7XAzqw2PG4/Fjydl5tTKaatoy
h1z99aldyZtseTB+Trc5vDrJ6sHEWnrWuslIKcdZ7MBY6uj7kQwlkV1XZ4N8
3gnNGc14RwDkP1QQQPcOzWRlj6OZC2IUpUZNhjQmhQsBcpJTEgFkEwsAHssH
O1Bpoy4EI91cVX37HaJ9J2dLILHauik5wrx7PjkHS6HWY6+i+V6OoR/Lk+L3
3fhiwcTcI+0lnFpppm49T3iZNBx9gzNA0/sW1zFVo7ZDNhJN/WIlCme/fzxA
YjNq+mrWL2sTC3801ySWnM8bjnBvCHLODkBeauLjGmsyXoim3DKHVHKc81W6
FiEs83IPOqe1ox6WPPgCgOlE9hi7jVbC3qILVMdAOYR8EqXOL56v4EDjaFfn
vcR+LkAPau40Sr8Bi1BKCPMF3u97E5xAQCQV/L65pbwjP+cP00G6cBAESXW5
jq4sDUmeEqZp5cvdUZW55uLV5a181s9Pu55VzYFDti4Epl8yF6CmflnViR01
HMqMaVviv23jd0s3L2RGdwe8iDCyrnbA9IMTBQg8fKxYIrDNAuoDrQgoPMVC
D8LCquPuUpZl1AG8YnEOrzzYJY4NOSqhn1X9IMdbCn23UA5UW8pV92kch8TM
cq9F7LmGHxQAp8q+ekF4OgsLthZxiOa9AVh2jOmwYmB1vY3/tMrZ96wQeeb/
o2K+pPX0Z81WrHtyq/Nv/lJSSt4vAhSVPzVooPOwNPc5YZFjAwAFCtwooafA
31C+n2Q2OKzny+OwjLbhVRZADDqYzJePZsPeQwmBDPbwZsjg0x0QQ+xWhORB
KdCZuOk0gsO7hCI1on68mpnNBp6lqwWFQJOABPymYluAe5tZSRdGEBJwo46L
ZwCItPcfR4Ue0fb0e2gYRpOiupy+0DQvZknxM7yr70zL1TogIA4g4JyG9oV9
ulmraVdGnGzpQTPgXNMAHMw4e9qeqcmn84R3ZNCu2UfyXOP0Mj8WElR/8FYr
2Fgt4GjW8Cjv5hdkYaEWAe9w3usc8f+6Xev/DFhxGt0KtSji7/tTQ2UELgl9
0Hp5+d3zPK6Div3RJ9tDoF+XhEN6/j6WPRMoXEA2PfD/xjSaej05nZFoFGAs
h2hUpDnaTwSiMvOfbdzdLa/bS4uH469JTcNTQMEsHBhehU2cr04w0AOh650z
WHSd2vauV4Wd3cMSyP6JHNk/NMKbyPQjBNNYz7vD8F9tcPkSG8g5YVH4LCIE
nPkyuW1E8raFTQ/X9WbOdG8Pz5L13dqwojOuD1J5R6goB+kNy66PUvGdCTL8
RnEVDU+fLlTdgdYnywIK4d6PO5L/QdlipFVe8wYdjMY5yJiKudgnr/OnjCSu
pSKJku3H+LFGBnSwwPnO/qo2e4D7wjpwm6tK6jC+A589X3cZKG2k/FoX8N4O
JhV6KYC9aq9/nscdOfQ8pxw+P3scGjwKXWFG2ulvIlF8BzrJnDSQPSdHsqgC
qOntzuhEGWBs9KpqrvluZ9I0FpJ2RN7ocYmdrWDYvlIY6ZfY93l9LPCH3EjU
so5RmkjLAyKSBmLlkapx+Q00miRJMJVHAuLxa8AdmQfBA+81y/2Om6QXEoPQ
pcptJHKsXqbSrwNXMBdw1O2b+QlKQAf1Ov3SVyvqOHoUKYrEJqdmWnIjSE9N
poe0zhX4A9LHOx/DSHmecHqVV5Ki4Ld0dO7Py/MeQ513IoXhgOW6vGZmcdDB
TA41TBGyc+y2ZXAdcbaFQ1K85vtXp5w2GDFp+nmF3rQzCAZYHIi2E++Rrtur
SKPs2bEWeTRM492Td6Im2s4Z6pd+3BySFJR5zfYUgJkZXXx+oNVhYnoZg0Jc
GAnaSsMqmWgXZ04+hMKowz6z3JJ7Y9D6P7L0i5dpgD2ktBQ2xLqLgqLO5bDl
2IRKp7et3voOxBXJ4lFAQtYnlOrV94rDXxo/eazAFWBZ/Z6hazRD2ncOFzZT
5n8PgejPTPRidwaLvOuFEisjUnL8aYTAIvc49w8dMMQkli+G7TRqcNsmb80T
pWFxnabZ2Ojx+G4J7/E/DbXsrcBrC8KB9O5l9rZO/ZAdH5q9Wyj/g8t+yW5s
4qoPwd3bEibf3khTbZ9b0iceid8NsU7hYaiIYU3q6D/IhYEaSnJ6O2yEJ9nb
n/YvtVhw1pw5wfWQ6gp9QLPsMvr3h0Iyogtzo3fiK7OLth6Oi+XO8CECmV/u
64a7sL2AzEX0x1EN5DBQu4kuYkk62cgaUifsOOinvwMupx0vdhUXHGdVc1OD
3F3nl6AYd38cVgNj0Tpy4T3X/d2x+/JZQFFRBA7FB91QTD1TUj8934JqKlOu
28cDh44fw+qNjxnI0XGdgAJoTT7DKj5FdXzpSpepMO7o6v8fJLTDdfyzTEv/
ssjZIpERvNhGKaz7KsOIl1lyJ62aoFdvRdTCvPIN0+PE/dmqDxCWOPw/GV6W
P4upbi2mlF7l6RIlvT36Ze6kvn3T7jB27OQ3St4OQz3uvqmno3l5A39RKdb7
giLY6ZdlGGKOGiRwLn1HSJ3iUUGvZDZ1Kybe+lAgwrTfosg3W6e3oUDOdGDA
XOBqkv2XkRxj6Qo2silU6tuQImw5vpLY7y/ud5ZuUj6CfDJAhw7qN7bBxHzg
MrWZ3DGsWYAaq7hdOUb/DjDjYLvz49x01rdJl0FyyPhFzIga1mDu2btYIsOR
9UUrKZWGQ81pNeF8nOck7g313uYWZh0rFP9UQiZoNSYzxATBtMZnxs3AGSry
5FyjR6qn0zZua13FAP2EpD3EpoQBojz/26NLp7vgMPG2vUd16Gn8cce34mP/
VcTjF8UOxESWXbxQ00bXzww2+uT/i05iApa1g+8vqiw9HBuXI4PBNTgv7XVI
nwWX2QE34Nb9HepRQsGJeKv326fu4ei+A/VZ1Ug5o1JidIX71h8a33pTKTb1
SEmVziJdax4lh3muli1Uiy6ZmEUDuElYZDlk6PH8/pT6MhPzIykhpQeooI8T
8jFGlYsSSBzg9VdP/e3urhEsQDqV3ryapqyKTaXA3X1o+YSKvMG4Le9oTVu9
GJkIhABIp2fBSsTW7VWWE9Ei5IpVpXSXPAPNsEnNpJQDO/DY8WrPVqBWkfq5
XErfHqhtnUjIZ04Man8dpRBS1KURGNLG6hOX2V4r7QeL5f0ECjZIcydXcU57
vLays96cFBBXxWXe12gjewVZcZDYqVw8o9L5nLtrkAy1NFqGtJnXvE/BqVDf
Kkdxp6L4Oh4Ld6Kdx0tj1Fp2dCC7PtXyzmCrx/vdVX9pblGsxMgRPZyGMv4A
10kAp2dqVkQlE7tZjddyPy8VNxY3gT+odRhpz2DvhpfmheAeR4vX1MELL5ky
A4PCVlApLozpDA8BCD50U7x6GDCtB10mRvP821P30pF3fcPp2Tv2+B558GDa
TBp3MLbkG2X60uIOJrrGKOIMFb/UlLXPHPUakXUNB/XW1NcyJcWMJz0aT6dU
gQPDKz3nrjH3inrKukRUyC1ByOTPqdivkhF2v7F35UuyMNyP9SGz8Yr9DG3M
CfGvEJJtS7XtuZUMzApTWnzQfHwZ+9dZtqjPREJbfIgIGhFmZHwA3cnQZk0p
8w2Asg487ve5wViDPo57M5of6+DFbXhaP6+FrI2NrFf5yxzYxioS7uTBYmfh
OkBc8+y5kyz2S2klRBaM5cvSikkcIGU/+WgnVa0XQopVY7C1Q4ODCK/JkOkN
aviqJU1cu8cUvw/5+w6o2w01aMSu1P8u2u50FoLxdqCY5Jd+nY03KeFiX8pF
W6weyy04Rq4ymsyjvUwnCSQYDNCl5iEuZXuwWsmgCauZy16ipSJYhTWZ8pGV
bE7sSgeRCuU/8VUD25fS0iGxp9qsD6FUGeeNO3IveTBsUSsdxnYWbASZRxPf
I8B/cPL+r6WrqHRhtCb1ndSgD0erGQc1x6tynFPwhAT3sppuW2EDFPnQGuCD
DUcIJXhiwmNJM6sn2Mz8u9O/gPl9kosqq1x6oQEp4t2KEfy2+te5MvqAMNk3
vLfKu+XI/lGgLSBXRmbVNnv9kOq4dvdRiNiR3Muy8coZnNMKglUK1HL/S2h2
5AC+Hj2ve8MwK2662saep85UcNo/6TTx9lxTgdY7cXD5GBWwZCshaY3Li1eP
bLh+SDzuNY0k9xZHNR8LwPkAHJXiXuO84iY6OUNhfTr566VZMd4MB51VweNh
ObKznKWoX1E50cW5nqzlcP7ygUsPNln6S8WTkhlPDUBmqDMVepI9jZU+M4LN
3JMEcb7avOcTO4Arapd48aVLVDJsij5oiwng4lSfZRf2CDFCfD6X5e8V0RE5
N6ieVH/AgcRF1B8izmPK9NAJPPKUBb+IwxUPDdBdRO8UdgRNu9KRzU/m35q7
6uAJauF5rbVvYaVHwiMeZ3LB5s9E80c/m8Ei9B8MBud7J8n1TE4A147AwRbD
Th8jJdPtQ71IJa4Kh0Cm/+QXTcY476p1IXlqq3uUaja7M5kaFpWvN6xdCQDX
GqBKIx2Cedza3Infwkvi8L41iueG+eIfMdMaWXbtRP0jUSh5Xw5IJdy8swpH
gfCeLO2T1gAaAeTZVYRY8f591C8x0odvjbb1I7HHgPKvof/ZmgYUx/brS6wT
Pf7VNIH+Fu3SQ46nUhtwyesCxPvcdDCo1EIbRdAR9DIo0KPR7ffArHOYaOUx
pRBYVHF7Olop74T/3qC9KeFPz3df7lcust0rMJ8a0Ab8rSdK/YgblFHbrBQC
37mpD0MizpLbyrBBJei0t1IPuLtJYc/037IK03D3ofng4GFkSDr/bN9MRl5X
hqXy+nX96XD5nh8vOst1B3EKt9GEad2SKWLBHTAmRwXdVvRH70YbdSxTpzcU
0z3nRjcBUdw+Iy7vaLT2D58s1ZsVrqW2B2nejbF6rw6Ez3nuggR7O+uo1p7w
I0pABVv1LadKuNCnYxDO0MiQBhvOKb+UWUIauYINZWB0TZZtQJGLm0EgbxFW
+pwYYz3UGCPs+9vMgnmN+25uL5Ol7CwFR5DslQeHxyxAyuZo5KrbjgLjEdf7
fCsDifqDsrF3GxjdzSzx0zaSV+woATtSIiqE9eJ1nlVsPMIOoVmZUdD3zBAL
Rz87FjP/bABonlYrt3St5RYJkac2GvjVtJyXCxLzK8Hbri54g0QMnsESGoME
7UcJHyuN1ABwnCnM1AwUfSTtHrroZTS/crG4fon0LQTi1cS+C+FpB5atmaqg
FCB106ofnXy1aP1m3izNsJhC8ZsIQbOtfyPSs3/VMq/R7HJVZtgtE6kPhrWq
0SGOQvfz01GIgRHpriGCzjjPF0dZDH0/5x3He6Jk2cOov6qN3kwCtqrGFXVr
OArawKwXQJrP3PufhAfLhb2COzF8TP0rJzxIaiK5rkshPftKbVQ3y3jWalMh
mLtj9jz2bGs5Ex4A6W5VtKYOtIfqPaDvMKAKoUps6e81JWAAsw2shVzWycCG
Enobg6f+zfvqef49yutOlDjhvIpTNx417AOpZbuP0EYgtxmAzsvh9XCjy3hg
oWVfBzC1flMQ3MhLwv+ZtHZkLhmbqxvgTuSYBHq76nLb2ff96Oe5EvswLdUd
Dj1ldqC8Bqk7kh5CReOjDgyqL+PIl9Unv5ArZSGB8cKiolzrW0u9hOJgp1X1
aDfYEv4N+zolvbUWkfrZueKmYNab/B7IIFfXO39el5ZKFlN7i+1tYi7AdbV7
3vM9jEJ3ykGHF/39BduEBObR/bpEX5IYlN1AyR4VVLF7KGaYiuoVnp6yrm+/
lpaxatGLQJzPQJoFyGxDh4R915PixsmF9phG3Qpz6BDyyYDx/nN8wTQ1o6p9
0Q670Es345NdABYk1PHQkuDDdPdZZfKwf4RUXWGr3z+gmicbpZq28kRlhPqN
fucHBkVqJf9BhXtizqCrXan+UOVAR78Gwr4rAAs5ae7PnNfIFQizR/twdBjp
lc/Y5QjUVGamOtomAFBbMDzIPGN7zLMadJp2zjHe7GQvNCKL2wvZ16IqRYEZ
VHvU/mSFR1WKw1tSUEHr0vKV8QF+umVKcxgu53IyOLvNLsHOtlX38Hto6Epp
5sp/ki60LYRgrVP76s/oeaG+R6iaEJE3kKBLjKbmd0D1e4ZlbfOHf6WTJ/Nk
ZkucPg8KP7gyb4xTGnXYI1+dMRhvSANBPF/VtfyYnD38VdxmbGa7bC8Voc6t
r0G+neGeXVn9nSREdi/PD0Feu/Q4MSjouXALaWloVjbXYmyn29YSPYpg4BHA
BXddsz41BODEniAOs/cW0etYyFFQ7sLUyMjBHxMlfTgzTaCRHe9ivcOMfCpL
dN6EuIYPPIFJ0PrZpidrmkgSHu03ogs0Bhr1/tG8p8qtsIbe8GSLxymnrULs
3ybnaDGqEZDzNtkRBRLqLC4sx7zZJckNAwuosCt69/+1IbmK5ORofVpdUDjb
RmwUt0hQDe1t/k3AfJjs7zKZj4Mycq1+g4IC+ESPMLFDHmEvModTpENzmrF4
E5i2bI+LLVx2MuqAwwBo8TUaqeKemZ2VhJij+nORCf3ToGKTiVGzAV0ASxnR
SQ5AI6Y6+MzUznLtKqS0CPtq8r5J5cuCmlf/9haKuof3C37KXdgE6Hh3WIn9
ODzjUIRL+fcdaxg5IPBvYgpebF+al1Uqf3sqgZE7yKtTA3R/hI7bEt1w4yJf
nYRENPID/XnsJcIZ26C0dYT2RZANwVtaHsZbNhEjYfVgLiDvyA01Fp74GZ7q
pKPH/xEoo4TjUMq8MgU7k+Wrcmcz7m4LKzwoZsoKFyFgxVzfOM+8W1ttX69G
WLJpFF7/yBpe+Vydyi32zUJcOtI0twe0cMgKIXCeg99A6zQ3aXR8YsF4YxPW
bvpY2WsD4D3CEXWyud1W8kqhhGMhU46w+FzUXwBr6KrEqyy+XcsahYIqdaBO
L7yCLz4JXerOIp9mzJ3f71Zn2sDxD7Ca40ASg9fyupXSk4leLRUWFOB9m9V0
Y17rMoOhEVZJllsIkCkLQge2yaGcWzlfzVs36MRv3X1Enf+XSZ+pv8UfYWHT
mCE5I1yGbFr8ZayaosDkWYXwYdkLmRBIXeP0iSlITbVht4Le+TTyMKKaqzpM
HEaDAqsN6UTnl6KhcrGHRSt/TXbr3faBriFxZtkCe6oYjKpervcEl5NixmMx
3bpQyyzxu6jEfFZjUL1+pVg6eKSABbRJMTg3llVYa5A5SeHk6MwL6qpzr0h1
nFdQLRL5Y6QtmqRUTLZUh0vGY1uOZPQwFljFE2u9LH5VsUfsdk0SXu0oUDlK
NMUaWENSPneU1I+Gpm7ihbpkqoyJyvn2xmLn1qKShM4vbvk6JRAbenDJd9Q2
DYNSgw0xqpaHyppXXdBPDjQUi2gXaF3QwhT2o4eVMNt+/6Eoo3+ZXgHfP1Ex
yhzlAhKCeGgsslHG71T5hcQJM1c+qGbWyPC79BZ9heuzAOaIvuierWBi21nl
0sJxI+KW8jL6OypQodT/rRmfQiMMmgwEenbFQ7hg1ZFtp6/Pt2Hz3YtoVSs4
5MXCLLBoccaqbRqcFdhWP0kw28eeebhYM1ndChwcwQ/AhVgx2JbjfOxTxOVm
dG6uTrCpNIDbM9ihm6ktA3UFAhGjQ3xpcQ1qbuJyMeHMT2XP2fGwf87xo4hj
WV7N/QjAArRu9yKDKNSVwL/ZFvAAdBGZPhdHgV4xOkabt1M4oIZggllVxLy/
I6Y9KShj/ZviqfR5h+D381TxqIdN61f0VzDV8/zi6sRoS4wZBDgioudMVI+h
OqI6C0HkFMIS1wZc2kvwIpb7qWTo6fSi/B2SAeo3LAkKHoUcnf7vWe0Rpr7Z
06ws+0URc/+jA+OqrXnTt3CqXZmqI6A8Dz/aUZ5raA8jt1hH8JGbSpMuPJoi
g1oxxXCmxMQkEyf0IaGfRUoTllFILoOu50x40PHgAdJM/Hq4kLo857qgnZrV
gJB1rIL8xsER3O9fusC6supDPBCExlfFoP3iylJwGDf/IdJdqzM2373bMXcG
NjiO0PXstnbZrCIaQPj1e+cTOFwvIcULuGj407zaSXcUsna7VgP3SQXAeaxK
8rM7VVKK3pobShO0fad12MDIoKjk5UNkUHbTZKOuryqBrm25jW0fYA8RtbuC
X6gOxm/rnssKr80Ft7fnWxUM3JdxNGlaiBzwp1I6wynPY6AS5R8XS4U0tAUD
zj3davwjkxU4I51l62ltTR/T0VpWx6x2PKZNekv3kKMWiX2JulgSvWQsV0tO
9QuyNJ44WIvweU0SVr14DLYymBouGNI/9p3N8r270faWH4bdP2Wbs0BnTRMF
EPMTs3IGXUsvYJYZ6aCZV8fBuygejAGPW2B/Nmc086pg+MuwIPpnDAVODLon
q1uVa2EnTjYCtA7hbt7sRQiA8DDfRsF0aihsAYGEAMr0WkRNEupqXE2d3obO
EwdwNnsA+rpp1OzfPoNf+IDUQAfkPzXPuTpsdI/kvFkIx1ism/WvhwZm8yMt
9VtvrljqQVAmGs1JBLXpMs15t4j8NwtTnDbZ9T03/NIYzjDyVcrTymM0us/I
3935jCS4QpvUD+1RUal/GF2Fb5UiAqDs9hySljKaZVRhAEbiUv2nz8ZnhQG5
XivQGTZQyiOGXqPXNWz6b1OLLPtiNS/wOox5E8m2JzSjbGMvE7GsnfAgqp0z
I3YZyR/xcc77GqdtKIacsRxHdzdfWEVeG76SeuX+Jd0WUyHMTZ4DOLRV+0Xy
t4Z9LQ8eGyUJN9uSsS3Hsy79S8k36z20y4xXA/oRQ6l55dBSRyaKoecKxhIK
h9RE+be4bV0388YmKKBqKXD6lpgG/p/Oz/k+f2DDtsmW/AvWVgcBLsRvUrR0
BLv95BlVPH/sfKTmpduvHSwTdJuvh6EFiG3EZsFM80uTB0NMNZgNQsQ4NKV/
dmXdiHdM/NbwUQTkZHhhEKwIeaR9VToGP9PSvasoMo5kwoshmBOzr+HFqCOP
0rfKzzOEW8GornBeeleQqoybb030yoswNOLfEfu75xjgxgJNt1zwIIn3vGZn
Edgf3yF/C74CANN2zBMyFZnK6y7WWObFne2qMz2HPvD0I2djhrU/f8Im53Gb
KwoWj7K/7nWGsV+5UVdHUjF6fEaFL9L+HLhMVzhPp01KW+PRsk69JG+pTFxy
9jSxMZUp45kbBdYWOWn5iN0BFvyvYlOqi0ahXDpoLzyjnIiRj3Dx5AM5KqGM
8RDkDRbahV16/hv5/MuXfJXPmZx4db1yewmVXaHD9i3Wukil4L/H/8z25If/
SlA20hrFNJWHR6yWwy3RyIKAVJ0UPG9Nztlg6RXhxu6Z1K1QoSvaIRtrCgtj
gSCbUhxBK6QHbr8UdjHHMCaX4PFwtlQa4ZtOym428J5XEZAp7arUcTtJxCeX
WWQB44j1vuLz7X+c8BroNQp9Wg7xwLS8Jc0D0f4siGKWvO3q0DMf63KhhSYU
g7najCPvfqgkN+F0UiVUEQxeMxfXl02jfeiZvSBVDwDEMDd2x1qwYKkPm/uv
9lIRyb1RmPGe8k0USIY8lRm1ODCepIy77q2Qyt31pBUMHFMMm3ezKDLscnHo
pq2IsvY4FANp/7u8Uas+LP0SSh8aDx2iWU5qSOHHVyI87a97O/76ig2om2I9
3QCBkqv2sJ4NtvUEdfkoCyxWha0aWQ4v0df+arb9B8THpNyN+UA4MGCDcGrC
vgbuXjoJ1m36HG2VOz5RkSTi0/L0RIqEN56FaVMxbjwaH0z/KrjtLyKcjVgT
LbfNRpXGzSQ8Q8aJSaUYrCoReF2BjU7qrB5jbpQCViDpxv3N1zjk4RvTC/Sr
19x87L2XmoUGSzPfwhg7LuEVtYlrL+2embXGzUrr/Sum5SdjToh8DMuI0b7/
vvn9EGUGdjB6vUgJBSC3YAxN5mkPUekLFZe2IHfcHoF3JLegBMUOI2Kr/m1p
UZ/O4j3WpWmiVWO1zCi7GnTCOIvn3xvro0F3mR+P0JXtiuQpwWgb2uk6hi8m
/57sbO/Gw23B2klI2Z8EucvheoPYFUQqgL+yY1zyL3hBzIFzNmYC4jljTjoC
hxrJkLRVN2hfxb742ZGj9GWXtlVL46TJDjIFzbVOOvj8fQ03ax3h/lrK+8KO
GgNiM1ysITUGBGGJABUWyJNOYAdSVVTrMfvpxggCC6ZHYagIdYBakRDem5e5
ynijrIT5UqAy5bNEjvv6NdVMBQKHDUKFtaNeokdQ5r3PVo4YtWWIOJF3/9RH
a/UQTLlYGs24jNtGqJlrdbXMMd2esPK2ES1we3s4WlyrdKVgYheETMCSpyL8
IvkIi9L16gf9JKmZoo0X19ENQTA+hl88nVhNfQRonKXSzswjSErW2Z9uYRQO
TG5qF3J0N2b6V8CNgU02WLnD92x+wZ1IgVWgFCXi8aLyyORguJIY0uPIm03v
g7Mltj+jb7zBHXwlsmHdZrq+87ElLA8gjp9QbZhcOLdMRBQu2WTi1KF9bRY/
AevaEImGF0IhawskV2wj5xyQCID9sgtBnz4f9RpkFGTnIPlnwqLBJdf0GjEj
c4Xs3K0V8tFdtoboE1iXtVgnEHOa2df1prqQxU5E6td9+JTYgpeFUnUG0Rl/
+NFP3I3vcCUgaPwGSsiGv9ptH+u5cz89tmjHP824n8X8b7lMyk6IdgBW71zO
ZPfAQTII5TaV1OLFvrdWD418i2O1jxipHgn0X5KJaIlx7sr3QO52Abq8hkwc
Mj5SFM9lvpmeH0aJ59iY89B1rSdMTfKIKKF98Ggj8iloIhhVKeooWuRTMIXJ
JnIpDM1llIFLrAJ+qX12KGVUjzyOKXel1yuVZrTjHd6g959dJr1sO+6WOgM9
6r9Zorq5/xLuDRNlDVzYqodO1Vvm6I59pmdRpyVH2YswQ08g7Rus0HteC1Kb
aNYpW1NUJFwH6C1GSYn7/q1qZhj5TyxIVMvpZW91YLgWrSYkzih8OGqth6SY
u2GVTewFBVINCtne43ZroAeancfzReAPexCZ/l5AQKRnsbWn8lW6PUuGc8sh
zKkPTLqWTJnS6D3uQuIDkWmeQbNpk8SnHu1hEy9Ygbx4sFms9uopOlenDpiW
wiS+RnbtN5qg1VAUmRe4wm2uO+2oMonm3jpLFcZWWv6mWlkbZTwBJPZOkCQu
uRmnAfi9TStA9HvmHZ21RrqEh02NeQUUSxHANQk3Q/Jqs97Ln/ZvXvNcI0+I
oJI8enwFDvPj1y8wbtGZKKAlV+yDGNh7liKjIHq+TxdqnlcayiODLMAwEeE1
tswdMz4pRbqXtFKHo0TYOpj8WFxzz8sZCXroUUgUtHAFUjCUPOmijGLIvu3U
E1wRVdFFQckg4OrkhAZ91ekx2IYHLBnULI4LYICCfKhv0EXtY4OosuHhvwD7
VW1rTlFtoJIVPOuVgvFwe9aGs+74/YdD+UnXtMlqb268avrUrNbQZ7WMVyK6
P0NPEVN8QFLByLV4l21nsYlNSeSnOFK6orTtXAD+QOIMXjdRq5CdCFGOV/r3
O2tzoLeu0Hhsf8sGqmniQyrdRd/ehDdI+eDCySDkxZcZN+Rk+Tz6qSKzuIK5
2/qPyDwkC95/lPTaEmJeeSSFGvQXrbNGBgCk4WxJqjEOBIGNN6ZoCySf1ikq
NjM53OEQAnJm11XpqZACHJl1KH0N4hqAdv269jm/hzNussRxIF8mIJB10XtL
ozLikXCnPpLs0fbr1/R1H8B1ZYa9wuJNyHeXBOJNn2Jnr+DjjXqyaVPesbGY
EAAJBTmKXkMtnXhWeKwtdra7oSg+B1+N5VXPP/GTJUXufCYSc1gprFMhsbHJ
FJoGGElxtmSqeQSqmxbeSpCyDtmiaiHpILk2PSeBOVJM5Fpcq8GEcAgbbrC0
tLA6yGQFW2QpQRHZcnpG4bL1bVsvXbNhhaTy9B/czoBnjQciVyMid8j/j//w
iGX+dSjJUT4tLItPqM7eGQsfG6zKmFHfA06Qei7qb0zWheNrPA44snHbQ+U4
ZabGnSEtf/Rees8uqSBkFKOw4O0Lrjt3geU7ZPL0A8K72ykOp3217H4T2AW4
bLCPwtS5EM5pKwjz7Ais0EYJk2ST64C563I6nT8M+MVXb1hqseSzDgwULann
hxbjjXspc5hTBwL7hTuZX5ccteVRFjk1Zu6PNwtrMTEFfml3fBTC0S301SCt
y/4tpHn4CKo56OMP6mW8PI0Zr3gBNQ4l0IbMmtS9SqSAAZSLKBy5OrC2b2u8
dnPHCqTXXNQuNz1QVg5yAmIuhEPewnp8DFh/K7FgV8D7jdYrH/a5ga/XWh9w
i/uIbeIMK2ChYgmepBHbZpZ7zDZSMe7ihHmDSp2O1wsmoWeFzeB5cklOfzkF
h4m6nBENGplhfie7n6x6vgHght6fsZCpkiqUvtptiAFVPY4m/s9F5o64kwuj
WJio/39HJ8Z3N5/qP2kfT9jrZDKJYHRu9Dgm/YPZC/ChjrWwxd3OecDxkQNT
QbHi7llFccN4JcL//6+g3tqYYW1lE2Gjw2tD6fpHDYuVZhozlpH+JXFT4qcb
AgJoAF0yvUUbH3fbC3W27408fMRWmnZKKtgUYACef1c585MkiSp5Qfjylded
6pi3BTphWvMKu6NRxaZuuP0lbxtPF4cyM/Cfm1zOivve6R33/hOK+RWPse1b
UkwcPvCfgNhpp1i7PDITlLWgnGoskB+8AA3vSub5+cv/dWg/OyLCVkocQmeX
u1QGZYi1yZzYtfP6Hu1dTh1Vp60oyVDDh7uwg0YFzKNPrt0BOSWmRZmgt5Vx
PG5B/H89qLndWGr/ZZThGhiEdL9DXlmY9MXyNs+hZVip/k6QeGhZf9UdOvEb
Npbpa0fZC/8VrWCyXvXT2YMeE9WwYWQYOOwVPSxGZWi1OYvnLX0Lbw9eJ8q+
ao3MYas0ejujk6keK8kvioEpjQ2qDUudsUpsVAYoq5QLzfK8OymESRwaMvU0
PXvRmWUPQjmPgojTMfxpeC/1GBCt/eJqnQHcEnLE5Kh3+yceya6igXdrbwLG
cnfQYVbqUKUE/nAKXWlnUnaxSG6N46WmKJg06U7SinHL0pfMyybWsBeXIiaL
VQaeocgTZrvmco39x+WTjMTvEcOIL9dK54b1Yjd3mCfpkdYyW9cCYfWcLw2u
VS8oOb8U2w3NlCCI16pY3Y/kwI3rHPyL0Vb6WdvtfvNrj3TZ6Aag61+hckLe
zgbcISq3vfS1nks/9yTuhj/PNmcK+n77OPlvaOCTRSryjhLtWNoVJCGa3B2A
KGhwCJClP+BH1PM/CIQzooNEexIkAAOFSfGILhrEFGAjcA4XN8sG9XLbcEd8
NyoxXWRe6yeGw1xYmrW9vxVUyW3rDk8isdSQgSxW2QN/7MF3XAjkvlreHiWE
9PigeDauDzeUEDNJeUTs2XVJXNk3rhlLaNF9amAHF+UgsfDfopjanh59cTPU
Lzc7yjp2MDhQ0Xyr/ZlVktxxMHviAQmWRJo+3UELHAEl+8vnNch2Bx0HaRYY
kvf34OErcoeV69UXC+usC5GdXvMXQwMFNgnMUpqHVraFtvrb0Caz+K2Ar+wq
F9rHswU0yzJNtJX5yqBbJw6WBcYF28z/RGNbeawzypDMsIFy0usDMwSVrA0H
EKCuFqu9KOo7mctwGqcP8Z62mFUD99ZWGWSPZfSNCE+WYYcxrdLyX4Q6yNmC
5n7a/cskn6jzXrVY0U6E//MHxMaUeeAaIoVGTT4gyvzHFvaXS/O/J9V4E8ua
01FDdwACOtAU4Y72P66iLHp6GFbQ+KjYMxI1qbMourr7myQQ8AN8mzIUADq4
gZmwQz9/0GD672Y61ESkuL5EHtayyGAXYfX6Uccw7oHc4sq2pX3Hxs7zm3U2
bPBQu7FdfgN7RHe4J6BThS0riWJduG6vk9BHtkhOUAE9WZpTnYsuRZKaVuoV
8SyUfhGn0+rRxuUtJQVkYxBPWqbrcLGV4VFPROOmwBJ2XxWljwzRfDvE7tp1
GKmii48unLTNfHnO2TTdOP0rbU+8szvXljAJXoIsFBpvG28gUAJboJwYFrsT
IYbxxGqWpUadmWq6JW9Z53+KEj0G5uo4HQOR/VTSAuAogBlLlcopXWyxjKjc
an5IZfuNOcZd9LL+V6pxMSBuVga2U7Kv1d7KeWEvELfzNRe3F7Ej+iJzeS+V
Tr8plJgfsCuJeGu605/a7Qhi8EJ6TahhIi60jqJO4+PCSENJb3nuATxKum/h
qTODml1Wo+L2FPHwi9eZZ93TYkU19WDi//wzLKRxbhe8wM71m0r3Cs01veCC
xE8xa5ZOrr/Y1Qoo+NH+AbNj0/nx2T44nXUQxdiG8CC7h5mqq80fFpzyqsHb
c8+Ets31kS4GqiMDgWDjy25pf+6GtTJlBiGsYp28jX4ehl+OZcnbjRCh0wnG
hWZ03kNvMyPjwjo+d0b5N4aUWqqELQImMyB6quvNc2CD95L3M+xRkUtwEXyG
cHihRa9+j/KVhjVQhEcDwM5tobVQ3G2Agby8VzqM6h4XPitVn9GbNsj0nQSQ
OfgCIvziaZkaIEQGBb6ZMr8btGv+mAdnXDaMjhmwhn5eqP6ZUFjraL2853Uf
b2I0uuKZ+Fh8EAgtxSUcGG5Eb1yAoq/vfGjG8IQ8M32ttNcPRsrohdtg9orx
kVJClvtLwg4a5IEyBMcn6IH90F3hxPpOYWNdO18VVcGBj6bcEIy3BjHUycUv
XCQpih4Nk+WNolf2nio+gdRQGtXfq9WMiQpS3Y/d8LWhC7aTt+takc12YZsR
QV9SaHHUsFWiSrL7TRtR2pZj0uuli6vW3NTJsd+8zJV6vEHIb4fx15dsOLzU
8q1kGLAhpYknpXhxW7qDts7xusjljQOv4Q2BWTW0nc1B/X+lrmHS64awh6tr
j6l5PrN4o3STDJxmmZBUnMCUTjeKxlv6dvsWAV53ICneJUig5eX3HRgi0tjT
UIrmoGjeWd3jLMXcxzxxmlNAZwbXvfxVVqjAAl6EDVfmmy2wyM9NYam+gzJt
C9OVd1cf6ZvG+pi8W75bCRqaP6k1Rs41uRblInIRwVM4PhsRouq7BVqC58se
8ZrNI5v88iF1sJoc+Mlvb5OoalSok7xTVkR6XXUPqHwaRNrznE6rHErDaztf
7Irg0LEr+Z/RQcM1eiEpj/ILeolTMh30aXRR8FEHPr+382eUmAYTYtkR/Ynp
a5bWY5rW1OX4yvdXuakZCYaVL5qy3GMmB8WaIx+b4RPP+RObFGboZxr9OewK
7y1/iNhLEnehDsIuTv4Mo3KHPTC6qmJqfXyx+4NA+pjESbSX2Vvd3JLRgvm+
yrdv/XhLEIDtegzVbGCiqe9BAyqJrzmxMAstOGMTnksrRQWv4Rfx+KjVBNvE
hPL5VwTKlhSStEclU7bZpqChEEBZafCDaRU47hnSpFEMr2JRxcTlvFiN2w34
mHjFimpRiftoIMoHCZJlnwC1NGZJF/H59v/9J6GsxcHjO9Dc263CHFpdU6hB
N/g+PdHQefRrV4e3ZCu420/UsWbnHDfruHIK+optUyybUomcVCFJ9pAUa+Wn
dWlTPjwdjHUc3VqpLa4mJtIHsNTlx9k8oFr+vTagi3r3KCfGMsw2+RWWbOI5
4Te5kzr887eMWtTuCzhAh0/oJrnv1g/moUyHEQ3Eee8j7IpVQAAWHFvNNtoB
3A0DkSpMGEsktKIWnpWLKIVJtBuN4dN17vaTscdiQzYC9RYQhcbqjcsjSA6a
3SmtAnaNRcIZioMSkCLBV8WucKrXuCsXfmTlG6zroQWna9WiH6gtnbIPX91L
mHeNjPuorsZirdx0vkLuNr2ipLTDLHRNGBbuId7NsYOi6Mf2l6fCjuo+7i4T
UoGpk2yfqWwBAk+z9f4NApVnJ8ttQNe6dZ2O/4Ji/RtIhkQPDPH14Kz6Hzpf
LHagaCgyhtghbGnWvOWiu/lQHBwp2bzCDqmozsQrZUxW3b7koN6+QHpg0avw
2TdUDEtqH9uMcqXRGqSNSsJDGnKyWWRw/sVZaVapVZ7KpczuVDR33P/B3Qhj
xxADBkDAFb1pfgSsjZ7+LYcVcuqWS6pxxvQe7T7QfF7WxU71Sz54iwku1d/0
Y9FbTsX9qlZvk6TI1DStk+CKPtKEBvaogJBUcyt7KXADNOKLAug1hRUn/lc8
i1oucneTroXJGQpAEGFPR2b9jvOyP1hsef9/BHDl0Kys2VEEV4P6mkbkvN52
rTvTESW0pjOXE3QhrXN4GZiqn5tv1HXIGDPAjUJvOXjZOVW+HjmwpTXTuaHk
HRga/ugu3Z3dWv/Jxu9A3DItsnwTKau8/qg5msz7sbwb9wkbbrTiULOxkgFA
QU+gfoGEVUr9ZS4wp9clNShzSjl6Qx8Ry5LqVrltFbF3tTOzBAs5WlQ435fZ
oYbsk9bldPESqpmLZjhgLg6htCDfo8MilpmCz7xT8G3i4hFJpoBCJrS3TxwV
FCztdPjqT31EgR60cRMejqpFnTr0JEHDMS5oY1CQa3NpzG9C8ylwarN1vVeI
i5exsz0HmQQAgsiH/jHl1pyBVF0ff9bOT37rCPkmaaU4TLEjF0SnpWncH6yI
KXDEIV8GRJCAzm232zNZPSWCa4NMGPgfOSCXt7wdpovIe7F1sbFgC06tQEpM
WXNCQLkmuyD1UmEpacwFEz0qC+1a6trGEEI3EY/nlcZDyWDbT5b6OtE+xtlx
aRuiE8ffq7k+clp+dmxQwT9N76p2RExMYZNvhL1jDoqYLqFzPNLIUfH7d61q
oAXIbihBAte7fne2/gev3RBEWIv4++ohl0dqK+/fthPzk1cqCgNdm9gAiEge
P9KVo3vDY7oI8QHcM8d47G6YkXo82nA/mS3En3puDh7AhhvzJ8npVNu20vgL
+0g8sM0iK7Rrf7HGvKkisoOwETeqv2t+tfXne/L1BGRf37sQ4NhgI+d6a6V8
WnkVdzhwtlVLwus7Fo+l18yVVwPHOfkEV6Yk51rs2gf6t10L75O47WbsBEsH
xMNszervAFltOs7OM6Th8IM0hgcRka71rg7JBBkfIqmz7pxvHS2Y+M9d3K3C
nirWw4TwRk3gUuKxYt7/benqvUMlamXkEzd8y3mLnA/Ilv3+yxwMQ0w0PJwF
FRfsP2XDzwqyck9roZeIcZo7BeND3WrZovlHjNml64/cyt5yw2nwD9+8LGFu
puQG6ow6mwarNLP6VDrKghWUdk0lPrzhf1XVq7sPXbUYJlgjVrpihaLVTSbh
YGeaO+kTBxVDmnBoprCIW4/acuHeAJYVGV+YJKGG5ci7l2pdHyNspNJP66Oh
Mn1yAS5qRuxE90E8rhvKl9u8KglgWpnyWaIIRtz9aJNDrN70sGOSkHK8SFVV
DsdDYnmu+75sHbmb7AnxsnGByTn8EYvltZUBke5pnSN9/AKpt0IrFhCqah/G
DGF63OFDz5iyb7aTeSwRCIG/tooRZo2kmweN4UMiq8YVcBTlB0ugn1paEWzo
1Pb5SO5XYeYt+f5SiWscBblHiXRpdNIbxzz3IhP08iLquNUXNlseevyPsvTN
noyw3UAYLupFv7/QmNEGcbr1dXDz6odV9i7xiRJNuBw1I6OAB5YGUYN9OUlD
E0xW53JUoTP3cIiTL25wWKSjpZRVlFQ9e9eC5e/qbNjTM+bpQYMOyS65KAjx
Wjg4fsBYpBqdBnUiWShFbepBGEGeKbQaS1rE4XiMLRGoJ8U6Z+gLOjD+rzSp
+rpnjNTxNejJywT6o87zAjD/6W1RCTM3sHzUJe1kCboEP7/bus08AkZPxRG+
i/j0U++s67FirGwx3K4WgrG+4ikZ0MzK/KvBK3ARas6Xz48T2BmFokWJXwBI
B7YVSonTGPmQDgvGxREHDUHxRmh5/paEDMts8KjFbu1ZIIo4QxPXdBwe1g/A
XRLiLMmKyDL0PyXIbTF9KWur1DONx9s8VL869ikT6w9zWUnMhYOxkO6HayEA
Quc+DoiC6BKk/yPXlw9/64vXbK1Pk3cvlq38kQKCP5GH2XD4sATV/i9fHbiH
iwGVP57N60I+06Tkur4yGUKdvAxdwVl82YMg1kFWXxcdycH21XZ6+o230SBv
m+s6NX+aCirc9sEUX77apXLQIHd1ITUp3GB/vSRAc4BFflrwz65f8UmtgCqs
3D39Urb/DBFsKx0MUBdTtPal53HQZHfcV56MVb7lnNNZVYx9G2IVwCIOyWud
CJyxmx+XXn0BR5KOZFLWnjutsVqa3jLXOZ1LdGcS0HE0gxL6tyDEge5x1JaT
cdg/hp5UeP3dDcdQOAOg/ShUqn/0+xsMc7oE839EL9W1DNf/snrDgdqbfIWG
Kj9eIl0ARbaMc9RQPvDv8RhqJfmgnS1v59G8A88RSuqnxsZfbpZ/tP5DqtDy
8wJpq967DmLgkWx21MF9ORrm5WJrft0q9xPrmNeQmze+b/Esf0R4PQR4YQzG
9FDNvhnoOV0qqZmjoNiAjJF71hP9CsonULiBAi2irj4vTKDqvybA9CTKMGdM
jbhvNsxGbU1u5bZt6yLNSgE7H76Pao20nbsxC8L3PTtm3INmAWlJpa2iDE5e
HE5FQiz/VlSy/MeZDtAmFZ+wA1DYc2Rr39BMEE4JnQNHh6dtVyS78GUrdPv1
uQRes853qfl1jRjHRBU5kuOONWlNmEr7Ubo+PsWIr9V0BxhUxNbatrcUNKXw
TF6aHzbdzczizzewGpEkiif7HMKv9GYWZugk1KJfE2NwqmDqZhDfAUnj2r+q
ZLfUyzsgU2On5uuwNzTyV80QrxLoJbQH97sCTSTD+WR+AeAsOHqJhBULf9u5
sMxgh+URJsCokTvGUdnu7lleiP3OVea0f31z9NkdKpAeFsPTF27o3r+egxFt
lsvPLGVIrhc3nqgTer3zYX/Pfwum40Mlf/EEPMJNu52/hjNtmCdYigvzrV4p
sArSWoKRK6MK6yB/gJHs3pCV8KFEcVWbAij3mI0xCDzcZdLAPcirboWW+Ncw
MsXXedRBee9nAMC1f273yyXPEYUvxJGk/O+DDyC3E0Wo8HC0adBkmFnQDwhk
i2tNFdtq0A9YnVElYRU+02cFMKS+KKt/4ydSngttdaGLzdJ70DrkyKUxGScm
zsWyolF9J/lnIH18djO7KeHt7bCNtqVHE2Ub5hu1IMf7vWa3kOGMx4E7Zqyq
tBWtjPbT6Hf0k5lXQlK2fdR3XC1M/XiP5NHUVdYx9ncjwB70Mv8C1fTCqGu9
ikqOzwLIh42oMx7gaBV0aJ/S4FkA+XTMjzq3RalMQ7jbC0O2Q/fLcnum9+EF
WryoSapHaIiEH5+uPv6zbXqmcnMGvdLabj/qpRtsYIBZqf+RogqqUft+jndU
N+WktpAtHoxwk8EqW+2Eg3Axdb3XcCX686LHSNsOmVruoWPor7vG8y5wFxev
SWC8UmIbMNhLQXi+PTE6pnHbeVIzutqwmx8DZ09DlgjMV7fwk+0ECtHHb2fP
w/8u64+k5W8UmrnzPkCdVl5OJ1TREA4u12+cbMFb3pmd70q59Nq7wNcQZz+O
QLzT9tRK8G0IC3wF+PSml41LcARTCPwiPgP/RF8CLpQVAtdj1i+agpiMlWWg
kOUsx0gmnOKtSdRbi5hJO8GOlueoSS2YdCfE/koifZwOrJl3xjIosh57vlbA
Un66RRpK7XMvOnBwVXot/s7SQXHktGcpgYDohGQ330EFbVmu2BaEF2bPuTgT
DjbxgYtmTxDtsydxrOIevHG3xjA05Xx0Uj/1lqMgqmx5+QI9KJnx3Fhpc1PL
X8bIXUx5qFKj0Z7csLVsIZBh38+20LwNAWNq2QOl0MCcI790oEdnM/bYiElp
BZmGB8b13qJHxa/BO1OlH5Z5dqvXXsnhjLJzBMFE8fHWeimm55ffNiBxPIN2
sU7dpj5yEDE89aPgfNn9FHGH4w9X0b6cPDeMseCsfon5yOupLaZ6256ia+gV
k5hwUvU/5YXTLWy4dvyzQv/BLZu+QPUvp30UEVVIo4Y9cJvaXikumVGfjoXO
rADQNyhQx635lrem8kmJLE22AMxeLHvHpeCmWFVwORRfj9L/eK5HVVEHV0OD
Pnt/J55jJc38RVBl3QCHGFHmwX6+gVm7DJwfs3ciENpS1KQvoLAh3Xpqd3PL
VxZrMMQLzgRSPqfuz3XIC/RKGYdtOF9uo33gb5BLFN4TLyb7xhng1jYFBS8p
pAnGKMx3+4rTsMusSw0LgEsXPQeO1ayVbEOg953f9d/ywHggowVuUa3C/IHG
oCMy0iRErKYieygzlGZJ1aZx1rZqTBugbrbNhOwLPVLlyO/Ay4147ddTsg4B
jsiBM9l6z2Pa+ZTQaxGp5WswwOeWu73O6gEd85WKyphp3EbBp667kQ0R9v0u
9BKfliOborhhUfJHmnZrTU9LaufO2xx/4fbx5fQGSa7lwVUUGQABTPI8Mvp+
jZ5kXwNuR303ri1Pw1ulGMHxEMx8KSyffzFs2SBJwk9z+S7EgB+iAq1ZkA0M
4zbA4UpeIfaT0lLHuzxq/vswi5fwn1bcI+HGhCK4od59xUqd66xRWK1bcKRX
Ru9846mlqK6U3AqlWK50//R+teY/Oxyy5iHlV3GQf4I6VCJZVXo4O0SqJstj
nkbF3j2k6liCL84KMQh+6bwczqHLWDyVhggBGgyZm/kAUFhwz33AYYKJMQKn
Dae29sbAva295x7Cr3Wuu1ZsUqZpSvMNx/O6NiFp61viCxwJ42fFp2xlSAEt
ct2dAjP+Xj1hwuro09tOEe4x5HH+92Kfp3gF11t2/IxOWaKv3H+4CTQVQLTt
ZhQR+uXxrwBlNV5iqvPjbBCHzjw2h50Qn2ogsoXFzqCz/9S7O/o8yYwOeFoi
KYWfBNjaSPXEKJI2vhkvKD6zBZHJFKfd0QU1d1l8TZVyDFWUiMSe3J/vd5R+
RVpLxj4XMgdWDRwD1MXWWuUmNlgs7Jl9aM6I9P6BCjTHlIvCrcTcHJqR62wb
GKAUKjqKNHxlzt6kDjONdPeOdzKbB+5zxRQxiNH2cZTcFAt1bi9A+1+YY1T4
oHfQGtd0HTEscFkhSn7o4EXDcTByXaUyvA3yHD2yUEYBO5FVBCmdcRs7Ocqx
X2xTAiGdL/r+oBStVeM0ENbiRcVviGWgNQ1XAYneVE9D5HOCC9CUYZw+JY1b
KW3TCPAeKxGiVINgn2ehi1TFZenZkPou+Vrp49FWs5u/U1ibW38AbqZB5uYN
1x/WLv5McyCxlD/A4l/nN4HZexBZUhnkyPp+xQR/uR1MGCjPmiNxggx8C5F5
fkY4xT0QcwbiPU3T0NcKnu9D+EL8GmjN2guAl2i/nlIkZ8qaP7c+S0L3/vhZ
DL4MdYrjLHzG3hmxHDOKP/TtvM7OMjerkDFMlSD4s3ekTJGcXz1DtoG7v1lO
F6hIwYe1qDERgrmGdW5JMKYsJugd+pB2xjSlfobEqL1PEuUn4bkymHFz3d+e
aWvV9Ev7ogzZR5/BGj3fLqxPi0IY96GnsiOcwvcDwKddV6FvS4LF3VItpPu8
tNCJhd8/QoAKV5aA+zyOj5vPxaJGzhu9fZDco6X4tkzner8QyN0fsypIVzaH
zVAG16ykuSc31HgFwTXpchE/NF96f9kO+YMkAgNgTW2LZh+qdY7aylWpwdET
dGN1p1PCF1HJhmhq2G2oScXI0p5da4jwqCrNWVrG8ukCvI8Yd5uvo8QUlqG4
/CdmsQsuV0K+LNJpkbjQ0VKUXTl2Ujb9dyCuiR6iQYr5M0IixPTWCoIC3kMm
Prg+TkpoLpPFUlPseunrbGuM+aOfBxGDc+KQA3czWXJ581jadby7RR0PtVAA
KVVNEVMhkn3MaG/rn8rgf9EF5N70ngRP8FzvNEN4r7q2rIkDeyyWNhCAkbk3
HAPjtQwk3VPAxgZgyUQA68jeGDRe7lo3DGGLH/4DKRfGXeaza//Vj5BHnplC
93Ul6Idll7sSQVvkEl/z2XaoRCkQG3aYNJ+WbQs9Fqy6v3hO8JJRMVTMTIjb
uwvKHRCRgpruBYi2nFfMs0mItW5PRvk74KBxcDhOGD2cYw5JMxqB/Z9BTows
waLwYbE83uQY8N71Ikjm3awIPAZYbTOVeHIaltPx5pe792D2Bkp83IixHUNS
gq7hGMlgt37XTy3Po5XqjR9ZZUSSwW0b7qB22jfQoH9LfUI+it+Ffq0vtyFC
4+pPFUn20PhrBh/K2x+dXVGry5T2ctME7fCFRfEx7zDmAeoHz2zy9XjjLGWw
YAXtKffL5LHGOombq+FwSkahl2fsXlO9ZLxmyBn+rCyoJHIRhLBNgwb2LuXT
13mVen6XYYoIezvjY1wYXLIWvYhCbCJ6ZyQXXWfy79nFmMbkWSaUhhEe6j7+
08AoeiBCxTC0HbwU/oNX/kbo4I778KgBiagera7zRlDHtdavaZ/XsD7EhLxi
eQox0nb4JpPFlVnnxLCPJUKPm8HVDY0FszxXdPYBvhnLBVPifnvmrwrmYS0e
0CHkSDzDlrpCH+oZOt3hIw8EWzY7k0P9n2zbSO3icEGzElFaNggPXuhTzt/Z
Kdm0ZiP/XHr9b/CPWChP75FF8cvGMOAu+6kGa4sNVe2imqQnHxPxp0uPfYhy
6Fdtx8VRba9fix17r7WDlBtp3EyrAA2vX1oxXGMGN+iDRCl7PG72FWtR9aCH
1e/eq2yvhZLVayyFSHXgphGV8PRzmf+ZdpNlPq39ZCoRTuPRiCQGqYeoTfEd
WmbbCnTMyHcyRO+sO/ZbMdsfhhFwuIbz/3bh3DiJvIcm90mHWW/Z3xhN6UfW
9FBINzuR5y2RfmAL9uwD+nsKlp6IkPP+dyROsQeuMAb9l0jbuwqQF5KWQQ/I
rB204LWOyYDjJbVWd3yVRYYXO7OCJ6y43A+zjGr/+5Tp34/kLGR8U0nEfRiS
cF7BecdkYsxz4epMAqL3PQAaISqyXNp9J4CEcxsrqAmiaLelkevmj3Dh+Dei
P5wnfFKljTIgWZergi9xfPj4A8Nq4+eWzAtv9zU3Y8CTHtjUhuOPtdnXvEfp
heO2PrnxkgVAtWxoM1Q+Eg468AOEA74LZdi8UQyEU6U0mK4AzMYQuCfSoAZ2
kTDbVlbsOleq3qgQujQ6cg5kacYQjCSTjmMGY1Ol0tOAJmt+SHwElFKoUGzp
1piB7aYZ60cgnrwuKAx7jhqKDM1aSthxeSKgiyCJz4Rj2nOkgQvErjZSgjQA
LsA6BJm9IgIU0JFim5zJSus78nXuLLG1gN3mj6sXvgCnlNQWOgxQlZJzwt77
f7nTJT3mKRSgIdcX6Qb9Dy28cBtNoGrKdHV/Zo/RXmGnqMgrr8hcjezr11Gt
NTgUmvmevd5HZaPxJIymsXaB9/qcKtOcwHokEAT0o2NX7EuZApkdw8+ChZFk
WitaWj7q3D7sIwPqW58NVE5ZdJSEWCu/r2u6APdCsJ/eh1x0X6H/ZbxRLPgU
h2iY3enrssSVlMMLlsbaTD1ZMQDk+iqEx2SgUXo3KlHwrBgaBgtttuQd2QlK
CkR95SzNrMp8Uiohk+pVcKJWyx886aLSIHYQ8teGIwSTm2s2dKDHFhCV1F+f
IWjpPTQGS0T+42XsDGluWmtGrLw+z3sUiQyvsFyU8NJf5GMcYCuRtyW5Mw4w
epjN/+Ps0YNWafjMi3WSoepgWQoejSx21fvGUW5YQznGJVVGksN8AyBm33a+
7wYkk7/wjHDd7J4NZcGvcISOGd9LaCgqNDil+gmqGMQ6D9qNOR3TgYn4Tlrc
puY9+jIzy3E7BY0u87Ab/EzeRQxCSqOV3ytBk0PFe5ok4nejB/9UenzaNL9y
NO+Qvrqp69D7l2o/QnGpB4Ea95Fx01+JCLncm9gbuYV9IK9sGwJK+actw75K
wF2PVwTjQ57KCwjjkRWIVDIC3DphBa+K22BHjmO5Ijpbpo9QPrHUDDV8O7rn
me4qQacbo3MHemInKTN86q2JbwGjQ4CI4D9CcYYhBSlyp9cxJ9sOWBFLbR9N
Tl8zWatMLWRqaIoxzDrymQ8t1MiPE8ZrtNJpZJS0Qhwy38YBcIS2LKlDeXJP
t3AeSei/C5FAjh4Sz/yVDxmi9/gKddnodCzpD8d2qKYXjzK2FCptbOymCIrB
ucOE+9P697eW8Ssb6poh9Fm3YA0MaspK2/k/xmvgyol18xVygqQTqNK1FWND
dn7TJDgMNBKVUWExysI3h9GQywfl5amaMs467BiN8HtyFYNLp8wrX36/8pge
dvmrm/CcqTlwKmo4hlSDmtAZKBMdlp0Gy7aAavX/3Fo5U80cD1Cx4xxiNFSM
8RTfRw7YQCJ8tdbTEah97Nl7E4MCnSrvHtcs/iWSWhWh9IK+slYPfaEYEKcW
UorROtduzNLiN99EQR5mhhskPyzQnaUMYXbb/KeCb9nG4N3gq9p/yKye+1uC
HWaHwFooIm4ARO3DT8HXrwG3xTGallcYLKhdWuQJJv2vcN9DOzf0e8kr+MJ1
pRqfhSw0YniyYYlosqddjuW02IQmDmwuiWTtipKKbYxnEyJ3iFHmhMfQ0KA7
cfzJv2OzILoWcwLgdutPDyU5zevrehyiI0I0KJFg70X+ArqqFYkfHnUlq2gS
MrqCPOXxFY3pOPFkbjiGuYY/Dhzc67V+htUawnfh48hmtrtRwmGU16MAF6ie
O1x076f+uk4t5Z8rXp/6wLkRSNtyvp1cHQHqvyNsvSKPQUDwEV6o2ImQjfay
QscGWfFB9OaNXSc0zzJF9p6oNPmezJxaTY8qqNJgaki4LDNx6LIILCy3jq0e
DcbGla8EdNDZ2Inz6bbRuii/s/vYQgZj0HGeCxIZTfMKKBZCdwEjNmKaNVuW
yTzIIdUAxC7bHZoTZS02PiXPk5t0T5efasAg6ZMo8TLI+xzpyfxE+rndkmLN
aRBqlNm2pTkAbbC26Rzx0IbBJcwY2rmw0sk6YgSVvaiUilyi7xj97NuwkE6r
+XtqyI2aLI34Rv+EKkWLCltHnUD2KNLXDO3cRkNFpFdmtswkP5QY7Rg1hE6L
H9jrabypqdIgqjmRYcRNY1oDtG3I8UPYjsG9+HUSzEeQbsCdfedTE84D0AsS
p27tUHkNBUtCPQ/TdxwecuNsqZsMJh5eGMWSDBFzF2ZQvoweHsFvQX936K0H
W9NUGZT6qqhednOh1KtpRSEaVVl+T0x6ioqS2do0LtsxlK6uTnDF1uaETFel
ePgNlQyURlIgnwSjz10H4dZcCb0+UPnHGdXU5OUy7KJrxe9SoQb2TUmZAoIH
z32zu/UgdhZuS+QpCO/HXrKYORXPDlOevgOq9pas985De8JpPawYW/u2ZnVu
LjPi2H4b4Q3VwimDNFWbBzT02ZEFGJKrGHQ/uq6ttTP2RSRVa1w0oU9uTPKj
MkaM9THom1pyEybnNadT+MsUckolBWs9FdtUeR8SHvbaYoW6KgzLZWgsqiQV
LATOc8P8wNZ5km+0JMO8l3QsycopI0CGGEHBHRY9cz+Lnmy3/JZDJf5x8Qzx
RFkj4VlslJc4tr6D1WbxG5awn42yoeRDj6RWNg5tS6XJ6AI45uISgAppBNJ+
PJTbktFI2Cbvj7XRwJdDyw7N2w0clTUv2L16ed4MwQry1dJetQciRLcmJTRP
fjrqhCTmktdbSbDYDADMJvqys/r3y9ZZdq+EgSVkEqxd+3QOcOscqUFZ6US+
+3al/Dv7zFRJBcwOsKtTXVIfHhX1lU2OpyQh0/crZW2GBVGJmT0DSVsHjs26
xojH+xuevhTiltQoAwO00yjh6KZncxza1I4NHU4gbV4fbG0CxebEn2TXzBvE
et19rYeN0e55PhM8+qFCAQ9UTTsuP71/d9kPGbULtau6rFnqfTDCONqWCq2e
6Z59hq99Nfhif4TqXdze0rhGSyK+u0bVxQK8lLQpeHuk07weR/PoObM74OKw
4GaSkjRxNTsbRwA9KKf7WX0zFi/3yFbfsD1JrvRk+OR9FyEPX6Z3zs7jqXnf
5/otcoaE4+gi9ZZFQmyMYLL4QnE7AXIRXSnuGy8EOxHCSAZKVtszK6Y6vw2v
7cuaiEIgN51lzNvZOaF7aeexoE88R+IhhXSjr1aAXSkcn2SWcxBw0vyC9oAu
RAKD7qNgBm256+zb6ksFa8ZZzY4tzcYvUWbUywFh0ycoJWOrFIQOE3JY/gg5
ERk0mYWPIcBtUORkC2gcGoHnkUmr6A06CdQ/GWPXmEOL4XRTnTDLU5TlM4jQ
Rqu7Ip8LSBYBUWsi5m2SLCFpJLO8s8Z4Tu1x7iN2IdnW0kavBS1rAdVBIw6f
m1pMrXiRXSYt78330QvzNSw/NTxhYqBItrkbwAvcbnVRcr378hA+YO9UH9Fc
LzSX1imsJyJKeilmS38aWwRy7++0e3fXVGIYdEXv8zf/iT2Zu8RTYqXgxhJ8
J81fiMFLrHcCLd/DfdmTWd1PMkkIiqCV5//OF7WfXL3XM7mAx13wOS30oOdG
cSe6knFR1taqqm9FNzM98DhmZ725qwcDpJGHs//6aUZ7Cb77f+h7BapwxG0m
L/JSICkelITovI732K15gMMVNTKYZMqNIxXv3am1aFr1lnoTKEt6MvYG9ka/
kdvUisGu33J7asjOnI9ZoR+LkghyhwrROZhzTYwFLzZpha8U2NLaWQoap/pj
bTdcluRig3cuz2YZtFUqRNx0IwHaISST/t/ZlkPtPC9pFuhFkB2hWRjNgMRc
2nS2SbNtu/+3s75nFX+unMTv/F6RIOTBSlMtlrOAaZm4tpi61mIclIC7UCRn
hTLOf4bGIBjnHcW/uzs+CR0eFrxzqK3OdB5fSNKc/B7JvKl4mBgvT78CN5J0
wRl+kLqn38c7TvrNDba0eXPg2xIlWgde5yuGRKfDjVxxw/4Emo8WD6H3IeP4
s34b4eiYQh6ngldAZ9bC97+ZkkTGZ33lhuGeXMzg+tJEX1oktoTxpFlXXO1J
YQe4UQC05hO4V6kDIxxJlX3PvShLP9yxpIn6zF0fGt/U/ZemyO1LE6vQn+Pw
QqeaMogxF061pF45mRz25gw8OHAHURzOc9yAk4vP2WdFNQZt8xMmSu/i/AmX
ba4H4/DTiZ5r8DfgynyGbnvygD2iV0B76GliBYLss62ple+Pz8QZKxy4BsoB
ytHBuHezD+ezZ2+KkX170riGMhwdGHREgMJP/3BDlKkt4Ib2g7TlYmzvKszM
1pOfuKSZn/ms6JfAxgrj/iSMeFqeYhAaWj98gk+CeBFMx4adaBZQs4dGCqI+
4oUH771mh3sHV5PBtDOZTanP/HGrRZru3xuOdjXwTbcHtqziPJvxLdXGNB5/
2duvZlQ9Fi+ZMMcuaDOZvxvPXlr0CSzTzUOO8KBHhcg6dLnVtBd3vYo5TE8U
aEkmMCmdaptgU8SLgY0lafeI7BFBQqYVhmJLeswXs/izjFBFcnHMX+L92S3X
thi2jT55hxsglxA38aM9S3n6MlXXCZTB9vdQ2SVN/DfyAHt0vlthFg9J3uI6
BcdlBgkJlDU/M++kGxME12wMlFhK8Apw3TWCmqH629IAYp6PndgS4H8hWNLG
/5C4BiFBrlLUP185q9acyKubMhzYqiN5rRYnvPSfvTjzkMpm+mfEk1P26scD
C1Z0ZExrQsMZrUt94uRkhroaZrNLJw+fp2XF6x5bpWGNbVLIHZM2uI/GtGyk
VyGmMRDZLB7V+b4fX2gcyDRL7sd7fyzM4VfAhOWJJ6zfT/K9mRKDbB2JPGYP
oBvhYsJNHSh0aL5OwxDodf4NjkxRASBdCTjCMBat8sNdsKjz6ltH3qfGS2Vy
NcykFnOJivrLaW8Ggkr+70jEka4khe0plZv6+J4Wse6gAVJw5fEAblJL8q2H
WcB9cTh5ZIAgDIMJkqDxRU31I7k3Y7aJyg2P7Fhrsarxx6s1p6GykOoR/wX0
EImxt4WllHZ6IAn4Ek5d0lt4C71tt8v2qaZ9HO7Pige4khw3IU5IU+HxE6WG
L2vhk2AtKKDoYWDvfdM+nexGEZ4EFt6dY/iev2ILN2p4Uanyn1LBpWGFmF/Y
5Z55Zc3aJUCWsR+hwgkn4WJ8oHhnHasuBci9w/eqyWTJ8jd6+dGLa2jWFViH
k/6v7KDoXhsyDK8sbFDaZrtcmmCpGAbB/yTlLIbdaE6RROuOaIh+knMr10SY
tLf3ER2XjSGXbljxDdueqtcspYrAN7e1XN2tZKVLAMlkXBUmIlXyH1kPN9bs
KFw0P1TCYfayDbEs468HZloYef/SYPcph5Hp10m57q8xuR/6IhHjTdw9c5ea
y6yGRnBUA66tQfK6+AOCKubcxJhKTwhlRNu8JBbqAZNexb+qcsikg5KrrzHL
6Kww5n+bNbeT0vRyRtvCXpbRElbSV4cjgZPSXZVZ2b6XenkWl7VWzuUsUPR0
ykqKKfQrZm3pZ59o/sMCCNU29jKqyW4xOnIw3Op+x8dX6gSZTtgM14GRUEiO
3Oz1PXjvTEk5aJMIbuFDYGJ0GN9Hd5hgySA+CsE3nG7tAmnYChpHGhc6CDQc
fmd3NKfa/tfkCfCDcvyir2lE+ZzfSsLc5UV/F1X1Qs7Vg9XUQKb/CivwSCe2
M5I9+13bjh+E3Xcvw8wY7I7YL+7OAkF62jZNvRXTHeGVVyorACuyLnwEplaR
ME0wpM5qp3XG1qevpsVIbMHogMhrdzFo2m4PzDH79LJDIzWxqwaZl3CTIXpU
kO9Ud0XjmPPOpiDFXXlBvFQWMEHBBq6is7z8/xt6i3b5h46L7wp13fpEsRGl
+ZID21Q3A+JZNZULvH/uzd8eKfzdowkYMhaR1WS+/OxKuGIZKs75jz3nxvcA
9exGS/w7P+fB/km8eXxfAmkuqs/R7UbbfwIqq3KwTcf6YkT3o2kKan4Zo3VE
F3Bs9taX4TgcZPqnAEZQpTDXv081EY/6TC8xrWWJkyGec5OjBVbRtP35SgDT
nxNBHRcXhutJ02EMlPj+yawmK7VXSbfTAdgfRd199BbKVjjGHH+RzqF/7dNT
uy7EBcRBUPYiSdqYzZX74iWrB9k6xonU6J8/e9ZhHHLsk4TkyVFDKFYXAiSw
+lym+7vFAQkwgIWbl04UhCVqm9gal9Kgsc+u3+TR42gi1xme7P44OL+rAWyj
PB6fSOp7vblCBk9fFQ+6NLNc7MlL6FoUyHmB7PDNpG2KkIRjjrMpeN1e+QDM
zByvrdRla4I+MP9+lMqppvkcVgEo5vs5o6nqDwR2cI+w2tSgkVnmUFkuj0+e
mz6yv2DajbpTRxjsQJW2ZlmUj97z3CintYyapwC3JXN0ddgV9tVO6FFRbp1L
u3Tk+F6YGKxPbVUXeBw+RN0GSLdljuYaOzDLQOvi4SZdfSlVrvmB7IkgG4iD
WbxSO16sG56wx5BkTfQmbBhoKFsA81lWsjbRI+bFuEWy940aVdxtg/RSYozq
5Ay9FV7eRMPDBd7IRLR2evMAJAN2gbhs9qQUexLA63ep3OtWER0D9KGCGAr8
WFlkkbQc1asGcHn2RM5SJ5ThMdLjQLV8E+1mGkmdvRT6ygrsIywJb55AZ+EK
q7YOt/ZYdDnoYwlXATrCJ1FO8K8LxOdgUXhEFcbBKuEjTKjL1+Etjx9Qj90l
hp5Twutda0z9mfThY00/qX/CdhN00xBh8Ev0bHjEV5u1D9GapaU9Hrp8YtQL
uzdz4bsW1UR2rqucjyIxsdKyrCjqdajqEp3ddRHtxfkzLlndsRNfet+0VRPR
3HhAmy3dOaIlF3jMYtGQX/kjzXjMt4jdinhV6NrNunr7VF43KT6wOYSg6oxq
fS18PnUYCVWVNSL4pNJAJhPTQa8o0YXDnt68yI6T9qOW25xXxWHHNmXxYGxK
iRh9sXBE5rCSwBOD8pUuD7mmvuxBIsfs+DPeflvEl7qbAdbHKXqC4FOXA9Cv
A+GgSz5G2x3bmxjKw2az/DyYVrW/9w0b74R8ute77yVvjZ03yYhjR2lfD5SW
C7QdpMPWOtpva8qrECdVAvom3wZtvhvxwjNRjKFTx9/Q5wXP5C/Mhsb3XWf+
fYSbM0xwkqPHW7V7wee4UjDkPepvlzAxo/X8PLkFctHi7HDeQpZ278NKkY1T
0rMXbXMmXF+4eOS1o0Xd8eQBbhT8V5DJMUg0368r7SJrcz1+RC1D6HaCXaBW
njKAV2M7X4e2lVoe4lpHovqfcLliQIbrjtS+F16hdHE1IBX3KNIUi/PAxo60
xceALJAapJbhnxfGcspcc6Q6yPavObMd3QpY532iO7rbJOkcj6nMHPyd5AOH
sYlDCxg+dWKntoyk/POVOa/JIuTOVYWnWbxYws8I8PKREe6SMihiYsCUIkoe
exAE3PGvUS6kwWFfw/YsYmoDQYrm1Zmjj163px4MV8Yo6WoIlZqFeyo4djRI
J+IBBHR1mFQqgH8e0Om++ad1zVFqMrs98pQ/qp74k8UktjC6FrhVX/zScHX3
yJv8JdOaQ+UBlDtJUrnwC3Pzp36Eb6tQCP/RIrvevEL9IvI1D5gUR3ifGGv8
F9oAsv3Wus7wumn13atpYcAb77ztKMxFwsVvCFQRAnuKrPZrxpwpjwi4Q+z7
5lQ4vq5Eu7hWl4uMU+YENJ4PPkHzcPU/WZXgfsJo5rLP++UgZEL5y10tu/DF
fYleQFwrta4i09VYJdTn0IcbUnidgWu4Z23URh+Bjs1GKJG6EScpR8ehW2UG
nuwf90DjQ089hSoHNOxLESHCAM+Rq46T32TlNo10ePvPGULRygiTRMdk6pP/
945zmuHCrezmI05b/Uwn8wK1wYHs8s9DbizeVt1hOTPb8pov95MZCxwD0+ft
d8oCEp54gAqmxWKKNteQOPyWo/ufppZQwC0nTokzuqNALjRR0wMRV2WYqNUI
E8j5S/JwFA0tpEmGEkb+VLrInQ/BRB2gJxoxLftJWD96xgsexWLW2Q25BI4U
Ea77FZ9Yyd98DwmvZpjjA0UKgtUo+SB02jy6CIsSrbv/YeGabO2cNIPcqvOx
Cn1YzE9oCC+BNXY/OPOYxhdyu4oUyYsApEAj3zU0MhYL7CGA3p6hnbrRGTxY
mMfrplQndYoBrKq5pAaq9IJR5EKf0trnikyYw6AHJ1mrj3ARbalb69JTVBKI
YmhZMCKJtVAyykW59mUBiWtEoLcpOIEXbCYmH3LJi0Fu4pqzRPCOSLFp1C/4
QiHqIRjCj1RecxBp7Yyw6L2RZoCsDLUukdha4McYq6q7BZk5F05SLze1XA7H
TKZ1e9r0MaGqr2CI/iCkEIURDFM3fmgskigi90WgDe7M5/mU94xOQ8rvhNln
tni6PCbLzJwhnFshWAEa36OR/EwONAQDtCGotDp1882uBKBgED6xUIplsThe
Lw+KCIULEwrkRM17gcwYKgEcEXkCYGYhPXLwXSIiMHhFtDZPLMKvvugumpam
Q3sheZ/sE4r+tnVH5sF6ihBIvTXptXQ1aXySlD9UPxxLewjX9ci442iFPGLC
PeS8mkk+pxJg4PnMU2vuODzx6B6EeDPbUtZnMhHomuQ5gTDULjZTrgVtFgNp
jZ/CDf3+UVmo0jCHKotWJPjzgShCwtSFA2qWLWP0YYZYQPPCNyRNqUTqSUJE
7hPvVvMHnM9TYO01etlYZGZAO26A/bYA0JrGPrKMBV9KqNn8ipM04l5e59wN
V/bbq1qa06MuNs8wQnFITzSVoo3QVFsaebwKT1dONEDi5wTJJvGUiyea59fV
kAB1JQMi2o7ZB+0GwNMMKp7IA5tAwmIW2l2IGszll74+qMaX/XYQj/ZuV4mR
Wp0U+PsrzfeVzotod6rzITXFL1rDNdEPBcbKEnawwz7dsaFel1Y0LBJ3jRWL
V7ny+CXCcWCmVycUNkvDLiQlYAOvsqsZCYYcnoM0drmbzc2cHqzyKWkvajC7
UvUpGgutTF9CjoVnRFIRJQ+diDiwD+KyTruC+uNK+5Z9URnzXEIX0RCLAKO+
jcv2g8KK4ZVAsLB0wVPbPEIgLWykWReMPfRJPhlND9AirHYe83EF4MvdPBUL
haI6RMmWfKN9Xq5fCOFgRPkU6LqgOrySzOA/vQSfkoNkkfZlchA5VRlr5Tny
v4aMO0/pfBGt829iTdCfLmeTxjzJnpP3J6oxGSp+fwwD34R2Hx9Vou8QmuW0
ZPOBMGVNbX70DguqmirIYApXOHAPjurX1ckGx3aMlRpxiAgImpw3p7WoZAJo
V0GxBN5Mw/n1VhkvpLBY4gRoQ+fl7D2HyNlCNYxfBXRf5i89cIHtCP8mMg2i
YHFi+6IAXVzlVPHoaR2V2JABhCAo+2RwAMyjvJFzZ9YxhAjaE0tSkDG1aw0+
4fe+pM72srcxxKxBljTRlT9ZrlDnbFmAXJ8Ouj4UYyid2RvHQf0xb95cceP8
GU0lT9E1dJiICrVGMzStlPogjxfTp+JQyOmrSGmtyhom9pEVrIRMrWjmL/YN
PdE9WVObzWtGtOrcn3AOxkZg0H8MPc/EvyqHvqe6H1OlDfKk3AMmyLK3b6WS
oSJ1otrnPvcCr15lieGb/Oj4X1jM9px+VKRM8NTrrJOJGhYrXotx5Zg1JoXO
SYP9oAFmHsoSP57xTdyASLKvMHxD954zWcUMvhR78V9XmoVJUosDLskEneW+
iYdWfbxHp9MvxXUck3f7MMs00P8ZBodfvJxcXP8Tdu38t2HInZOcHm6a33AP
hIfsSljfQ2qkfRKgF35YeVoKUP9HU7pcPbEIuFsl/2wsjhaIv6Pn2+8JgefU
9Q6orNNDgrL0wI4crKruNrv12fK5eDDaJzBIv+5IkBc9j/uVmmT/zrJzlil5
urfLDvEuwEvh6Trmj4CQ/fTDsH3epdUrZVDkgO2OoHQbEadusBXIHKBP4stW
qoFA+QT6kL+EvLog33TBrUTBsl8NZhVApzMOf1eZ7vVE/u/jiAyXGeCNH6r8
q2lHX51ediV7zwQFRHJ0M+1QKtLmiwTcCFkWS5EUL/TAk5EUaILwN4GBSI0X
hA4yVlOT6QblcSinhGo4aUUAKyJ2qnr0wdwtD5SJNNd4FPLvUYsXoJvAA6DX
pPxa6R/E5BBODZ/H4ckIbFZWlxP3h5CcBONh6eNR6x9qVVIbI8/WbJ/2AEt8
ta2Z8ngQvFmojvApMWm4Pgbj1xgdblX11mFCW9Cjo35PJXTq5zlHu7+Aq1e4
PzA00rEY4k03MCgMZYvd3wJmNIIM/qaMqhRarziehIy+G5FQeOuxp9k/dyCK
B7PbQCYy1HEa+ba4Iefdu1MF6YvipwK6Dx68iVVjfaWZqxon0iGro5QKBHXC
45Vqf3tLIk9ItW7w6B2+hqeKaChUfet88bjH14eSxxVxjqqslVMQvXMQYVuF
qf/1uGc99nn0WNGuyErugu+DdzQYQPuH7/v57231SunwCeuE21lQCBdMoJz9
gBjPDn1qeHYBCzbq5662Sh2EnBzSzjyN8RTXlUGJ/KA8BrDsXYPUONvaxrVr
fA4s49fkg690eUEMF11juEYkzDrFMslW+i7PrfO1xWJo1qcL96PDBn+QssOH
h1o442YoIZiXIbKN//TA2KVYudZiuP7dS1pYDr6padnnybOl2/b5R/nvQaE5
AQzwcVuVfIbqvJtsLwmO1urAs3qoYHcSUrObjJr65iBjCzMEJ0jgM3kmtuXh
pRFzofm+bxtOrnjecrucPrIa3Lvpfi6yz0uy+TKGqw5KLYTpba7Wbg5TvXPS
kqySNShzJg/a+oDI4ik4dDYGMBseNyUZ02GUiwukxB+aettv5KNBMdFc3kkO
LkWJG+wWxo4pdSVjjYTo9abLt/NGjzFn3QNhqKZF5KE7Jaoz46PfzHvqRJwo
sl7n/bsHenSiJ20prs+FmDDiXlc/hw9bOmMMRP1xWuXBbngiz5NM4KkEpZv5
SmWrAGXlAbnnFNAY6dZWafcCV5xYictfD5KvWfxMWAoyKonjNjSAx1w/g2RV
ocbWWDqDsYT0QB3Z3yfceQd+CxB+EjkpEmbRdwOCgK2ok8FU3Na6q/uKFyma
l95AcesnEV43mautgoAKMfKyBubADbPTFxQ2vQR1u7bRgYeCzyeewgguHC8D
9uwzpdSISGRsix+frUioRSI33VLtn5Fafkag0BNvMojoIS+eJ/1PfdgGmO2H
fimmnxj8urRKjnEj4QO1clSL0Nl6Xs5UMWsJgapdTeiFgdA/qop+7MrqHxa7
w9zNP+xBKVipAu/UH1I52kD9uLzHNujytMKwsWch47oZmqs5/pZuTkstOtkk
Er+C7vr/FohwnKxcV4ukt+SDWGA7rRCpNP8cGS7Ex2qPH6nsAUFnw0dCOLfu
pKipigBbac+9jSxqiDHjmpImeSnPEDLGSzFt8zfzq9Iz3oC2kgnoh5Rtv+nT
vnHd1dLMYk7gIqpbuJrUZZOFGE7lmINn15CGUtLM0sFuKaN/R7fy4KUIbHYd
0JOPnZc/im/ARS3W+0bxVYKaXr//br34LHCI2zD5ALhSA2nz3iwLPgy4/43v
yS0//P8FEoFIrMzBbJV1mHJcHxwq4aVG3hXdi71YlRkt4TMArwApBntMaQz1
mwV1lNkk1hQStXYJyyvJYW2DCj/yf9yv/QX9iE8sOsyt3508/Aydzf9hJSgW
7Kt8XTGwPNJcZRlx52vSSUEAMCYp2vnDmOApZ4p6kRoX1GjEfHf5p5BeEa9G
4qzRMdmM6a5xiIcAboiq2kBzh/gaO4VQIpJSDsawxWx26JhZ4z/NsAVUkFaB
UDh0Avg4TQHZMQRJR2sr9yyciMzcjtpulN4HiR78S6hfj5WvMrcaupMK3iCE
Y6NqDiA5dEJXZ9UbeEWyCMZ8nT/SzdYQMmNvDIYcCFlSTtfaIUGAdPcCLqCP
h5pJGgSPkGNozHcUK+m8ccWJvdn9/rjYwiiDv5CyExSabktU0FhJ1ifVMALd
3bNEj2eawI2yRf7/OpH3Go/kRXT5eTj/+/7VSjbb8Gvw12j6Cd4CamB6sZXK
Mz9+NUzxgQuuKhso6ltznT6BSxbwbLxBbZGMgf6qH9SZ/P2Uo5dpjC95Cl6P
uTgxBcUk2BjNWjstVvPQwZnfE6K2K2zw0i/XeZad4lGU8P5SPkSLj1P1EJWD
gV5EnbLNGF8euWXNbxcFb5gCKGQRULqA0OZ+forZdvXU5weTOv0fdAeWiOez
QXLuyUtGVd1CqIG6tbi8fzrbs+ZJIr7fRJ7NQxsQHwZQJDIDR3LPpjyoFM1o
MeUvF6Gv2SBP1TB1beisHxghhfQq1pdEypcHIy+Z1L+RF99WkJtmNoeWL41M
CwZBdUXjidBxM5XYvWB4CRP9GZxDOEL0OAsYJYeQwW3t6oYjetYdtg7sSov0
zvKZAe8V2nUa6Z90HJ7t6Jhxmmz3J6fiaw1tT5ZSY+t64cQHjAZT5wwBXDdr
VPiOYo/HiI54fdFf6iVqVUV45kPoXfO+iJLDcnH1opRovX+Q6BxKNukT+AKb
8VY4opFGncsgaxScgq9Tdw+qXb8v7tOyWAxhbXvLKyz0DHHVfM7kx0ScJdF5
6qHV+yjybyXzRPaf0CtMjiSHJ8kv5d9FAUomf3cAk2v8/yMGkRIXhT29j1zQ
LdQYsWmL2KIB2gcaNQK35SJYVke9e68MTA/tc+EXFkIXGAbioKeJ+Na9BWm1
C5z5KDuWL4fY97XIq5lBn0EmdU914Gnz6F/bpFr65GiTW8M5J3EZ68sKhk/N
RSn1IyPcYaZsGMagdFyU0hRUIXIWuSzb1pNsswnyvyzefRc3UU7Cw+7pJtUC
dGXtyoLJPVwiXbN5EENiUi6dspfcqFsqnibmx+1bZMpQPdLYkafATJoJ6L+v
gDqBYYG6FeSfbEqvklqbEQ4YcGSrwljkvD4YpdczEqMbizLpFX/cc2BPrXGr
cddswOalxb8x7LLCyPpB68p/jBgCrYV5Bz/VfxDon9wjRbjMddoAuLIThtan
bI7bP9uTRDSyc/eX5uGSAEKp1u/XE/MXl30MDNeDwN/WktjQn3Jx67tdOJU2
qysApSZrNjFWWbQ1zCCL+24+7XHYOlsQS7eBCBBaKmuQAa4Fd0Gf4gLxAVsP
bm04pOPzd2JSsNU61VKs5CmkM6q/Q7Z8gVbEK7ogJJGjJp05yLS/YmiropA9
FEh9zIUcog4VOmwE+cp+iZ5khGQYHEGobvIL7L//M0o36V1pzRmsKbjePojo
mWyK09bZkBlXnyfz8USH5pPUCgDT0AhQN6fbVbH7vQQzNIfKlsbKhlS06WMO
FJLne5i2pBPtxvxgfNDtBumtjtsYFFDg6lN8nxUWvZMKnj1ThTrowtBhcwQ1
leRed5rl6UkFstnvF1iwfA1tt6P/VEQDLOBc9RGtkWaFkjFXgIK74jycdeNA
a4UbCPk8kaWyjtFFW+n1D8voEB+tt99KP6OyzS9ykNir0SYqGCs5KEbekQjs
zEUBNqN8qyZ8k4AoVwKX2WsVzO7dllombPxr3oh1o+Fe5mp4Yp0AWiK3Ed+4
JSs15KRh2vwvEYAqQ56pFHBGRNkmJLkjOnHMrcNhu1WpPhnGs25UOELqjizs
f8HxWlIgvW+HwHKZDScsJ20xAxJhUJXFq4oZjb3Ebh+oaPqxQ51eaDwiaWA9
Fhat1W6mGS8rSg9oR50EXsEuuWEHsOTw4W9LVuTzFwVVMoffm++pANCNzz8Z
RXW5TFQKubTy/Nh2+ujg0QC9R7UkRAid2TJpiXy1HnpCbWvTdfAhG0CiomEH
fu3kFGcSpuqW8RN3ZBf3KEEisVs+oH4SZaXLlVIUkDfzAj6nxT81vlLVWar6
2nQSqvLoMOWh+7Eel3mSfAIxiGCsBYY6qbC9QhmUIrClHCEXdD0o5v6X/U3y
ne/fVf+NPPsA1JDJrb4SP4xl92X4Z1LUnxb/qdrBcWY6+rTTwWi4lPc7YTlO
IS219utcBoZw5+Mbe08MDar92EPxISXUAEOJQQ4N4ZwO6vk2IdRXIAkEy71T
gzeyxf5MCGZvzpxQPfSgJtRpBXpjU/HnLk6Rxx9F7A0/Hb6VQ0q7hkttj8Bm
PcJwzk0feEec/leksY9RGmXHmIkeVDvVkNQIQBhOBSaAPjcP2mRgY4c97oKL
a/U3HAgoQad78sH/uk/tHkJgiR/JSeppozEKUmH9l8uTSlhszYu7CcqAXdau
Z2RmTccbrhrA+3tyocML5xd0r/PsrtHykUHSphaXgvck9Cajq8sBjTTjICsd
zEdxKlYzcrWRTUyQMXehTJY6sFCw+jROjZJVDp3LO2/qGE13XoqIsd6zay8C
WgdzRQ+D8qT2TVosL2l5i5LWNtVYAbbGlxj0cdbmDEv9BnnUZSe5ZdV+kyLr
00wqntI2DRuASmdT+B3hFxyrGSu08z+ATncjBfL6gzmu99+VffjZFNyZk+WX
hj9OqkCuJYoJh9XRLrVVM5TuGzcYWGeeLMjTLiZ2+lcka847h2tkam9rxAcZ
gxyh8T2Fyyy0pMzCgMtEHr28/wa2o5hfWt/ziVf2RjK83s4fIbWCsp8RKkOZ
hlaw8D7by8Ajm74dUZrZzHx15i6/zHOpHKIUla1pND23/NTXoCAix99WeAoI
hAR94N4OKzfRs1g80IbRatjDdRzzkDlmdZegykGHnq0URN0mZIhj1OIJnQiO
mIhei/RMHKvjeCqCDA2tfF6+vZ2dE+R7l1BFop6AH2PFQ6s84iDQmbRNYTGb
Wr3q3tgIcaNX1HpvKEJqdmYb0T7ibZteHVeiajpO+A7RVEnDlpkbWTRs/SDu
IDoqM1TwsozWl5eT1Q3WZQVMCyyq3LVBlnc2fBDsYjRIwquLOKY/Jd1TXc2i
fH264Jl0pNszJbWmQkfL0Z1SwZIKuKFWka6478pfjNCv+e41RylhKs3CBNGq
I1n1qQIbN3C3pCxnvbAPRj8WJSlRl4RfdwAXhn+Q7K+KVkv18HWpTP8JwBkQ
ckIB5MGjhWPH9UQv+0TI2VbP1deAycDcssg96fCbxyLx8EcSlDM7yzzaFRJl
hdCKAO/lhas/0hlsxIMuF0unJmpANB3nsjTgZLfur2hlVYkV9WvKUIcPzmMx
IPC2n1um1nGD63R4jxbZU0b0DPMa0TDhYNremj3mm7+fhcFR+Kjg7qtyJ6eB
T1FUBaE0vfKVAymi3ItPH1jxNA9cSVnyUoOefOgEtbBVvnheOFSE3jIJVW7c
vDA91kTaFWP0PpkF3lHX3DRthfiyogD2Y3fyLezyharUS9EH1sNKlhWFP2ig
qox23Z+OjS9MwAWUaJSbc4f67UHKKL2hrtUFtvkdBwrCQ4j5zT84u5zbFx7i
Vk3yzj64MvgRf2Gy81QgntGtWk6zF2qdgjDOrDJr1aYktP9CzVpELRg1UuHd
kFK7i0e8Ehd3ONAIHPhfMmpqUVDSSDWYkF12qwy/kmaYmvxOAlTIZz0vFnyo
56D5WpimfIdJ0vcWVN+jHddFtNsBhUri0B//IedHWm9xG9xOuYgdtfEjhjix
HV4qpEbZcTrlnm8tqe1ORKJUKK1YP8GjBOFFkIPy72zGh6Pn+CRYBa1w4fyz
ZT2TtscRLOQG17+29SOH1wBYG/SDf7BWE+javHTe5QGMvME7nB2Dc7dX/O2R
WfsH8hx3VtQ0siyyeAaMBVAcSnyIkN09Cfk/0vVcg8CCdaeICmJIJbL9A6mY
tyR3qaLqstqUzgVKuorE/K6yDUdLJDOK/a1HYIABh9w7WTJNBfZZULdqBHId
21S4sWVYBDRIeX4L/lUD1bct32DtCd0O+IEhaKcdng9EexMmjs8WU/fgSdvj
53ry66qVvhY9/7R7a8O3FmEEVZqfvFmO27G6yFGYWZjrQLppm3Au4rjLTTlC
ABdawGLEP7lrcX7Rvs2/JeB3E7qx7cIFkzbRdSEPknZuVicVK+Lm/Cn+7Y63
ZS80KEBZqjJdrhcmC96XFZ6jLl9aNr3kHwv5dz/0eQrB+dp7yGtZaj0MmkCB
Tsxb+FX1GnQsaBwv8H9iHqP9+XiVNuBIKu2WyudJRYY/FvV35u9WgxaQ1OWc
O4VMq6SICIM09GI9v3ELQtIVEbb0FZHpgNTpNzXthqsfHZ38Y+ROFVrnlxSt
mBxgcXO9EOaKdtMR2Tv010ZUEqDyg4DJR9yAfOeBj0AbgQ3DgxURcUZUUvGb
bC5R0lDd2SnnO4KyLnB/lZ7h2GI/Eyj1CW5azjIttKii3mjrUBbdxjC0ZrG4
8wKGxQINmKNG6zQq9ZvzEuYL2yXaF/JX/we1iNal946GMen3he31rqSW/HrH
L4aHg2Rg01/AzfpZEFNIQf2vVtO2bDEv4064EeEXRW2tyq+paUlCDElETwu6
K7WhSJkxStGuO9diihpfvn5HNcaCpvgHoVmNxC2m/Tl+uYC/0GaQCsAi0u+2
3RzC+MwKSIuDbazFj3JYuFWyN8/5vW3P1PxUmg4vvv3+R+u1+2vTZbVSZS/l
4B4Azo5yZ+gi0tt30hyPREJyO+QV0qcV5IT5hF0XKd8zKpU80RhcjhUd8V9z
wgzfzQyFTggNe7F5GHX9VIxvX8jrXb7U04DLGmoCykJclw2+3QgNhSi9VM6a
X08W0ginDfoKhu/v+BEr7RzHwdA2ZosuBUuzL0ZqnCx94JWkDZrJ6khpyj4H
SULgqtkp6Jm7j2dIncqozSd2fvFCRYJB6qUjszXJNKQ9Z06FERbQzio2HLzn
X0jpTuXP7cthSbwaFxRatUioCv8wSNrvoba/IupygbZAWKbj5XkmfxDLDS7F
j61trlF5/+n5ZPwbf0GDbjvMfST4tZ7E/KcrIugYhWVgAHy76nSLWdRX083F
QkQEDUPk4FXfEUoJq76Kowh6pi6rPn3nxXVksh7DtDHq8r/RMF4O8f/tyVop
AKx2URW98re8ckBvve9g9UvA1nYdjmIzv0d/LqiTz9FMFmCrnKqiMAi0Shi+
s4rbbnY/cNhgNKXPk54izk/1ch1nBqcHrTqQtvj1nlwX2VNcp4b+NM8ijMiV
rYbOzvTA6dAR3NBuavLNJVC9pzk2Qo0GdkQvjoOPrFd9JsOij703H7xNmdrL
+7R2owDQTAXmn4gmqUL+6AVnmN6JZGHrXfvOyYmaepJ8Jw3FgASsr6/uPgmf
28D9aAmv5+cCQQmtHSWg2MSZ+hVj7pcxiceb3Y7sxjhJtm5OwPBaUqV3/RPP
8mTyfGYGyq1dj0OMA0HTsSKxqvOjOLiIa/K2wzmzDNZdtZgYKEaOR8b59LPm
zV7TiZQktHrNUex5SYuKRwSd8JIhqj6+YmqLx0Rs8hTKU08Rzuk4LLqXhjp6
IgVBDA4O1fXbmoIR3+I0JJ5ZX23Q8e/FTtqAFNdqVh+cHG+mowv1pA+1a8ri
gmLAYqw8f2a0+pev8KVVgWhZaFu19us3yGJBOsq0tJofVmCvi+vDsGHc2eqP
9LZCgTV8yCFZE9+r0uBdNOdYqiyJOVD2ahtV51+6Md9MU8EhZSUHPDz+lcXa
6wScvsqFzh0l+MsahjG/3u0eVQ4Kxr1FyscsH9M7VKMyFf+Jht2nnhCYCImL
bZiRNJD71KYsMYxLiMSb+yuLneZCoGtUvwdomufjFKZIo59rEdIt3fntFgy7
J7cZ1S6sNTL/oVRoy9gy+oQkdwJIutsy93bNBS6NKs7RXq7jFlPOm7S/k2CC
O5Dh0i/ag/Or/RrwiWREws7GXf6PqMtNEN26mT8GnqLkCzknXBznhQy4VTGJ
yqletYsksRoasoptipbCAA9m+rgpHyQU0q9wdbo4hkazliVfMizX3QNUkxxK
zlRwVolvNIjyvkjShmVjMKCl+/AemjVTWaEkgZ4Cicibtwh49rgOPAYtYjYB
6C4AaQ1MLyEQy75Wp/AF430MkuG3SBi9goQ9XIn3jsY/kudOPOHoArTC+XZO
INZaWR6PuYge9AYoDKv5Gea656kluv/XBdRhYl5DudeYPbgd1EDG+HL92ndv
7+DxYWtDxd7zZJcqlKRKuYJRzx/4KR41aLOKV7sx3xy9v18m0cY2YmxdaXIu
aEKR2mYNZF7+wdQ4wcS6NZUd65gm/ySsseeqH5wnHttC/JIbnP9q9G9IrxDq
JwilHHek2W0clOewnZPa3Qlk0OxX/4Ib/23KEUmu/Jy1OBOfAHdj20ShHLcs
gkSZ1xHFLgDn10mnKTC9wI9rKT/QbXP5f6nXDPEcHxliWmDqXxtV+xOp7hQ/
sIhp2oNThyatxGtPEYyA/zCWRdJhg9wIjVjAEbh1Gqhc7Mwwesa1AIJFhgcN
0oNxJ7dmSMyre/cxM2v1RqX2msJzkgRn6FAK2/DXG/K4Atf0oAunVfd/KKqJ
ZVUOyldFkCVet9uB5NQDpXcoTyz9T62K4Ge00+F0KaCp4stAEycEjKT7DkSY
u+eh2SeCivEPQF2MJRaNV4BIbrfHAY9849zJhKXWH7Wvryoi2y8G7OHeo2kS
+S9NzXxnzsK/+BsVAK5badmY8EE8lMh/HwXuN9vsMmhdWT5cjqwMHucxkAJc
hAPS/u0nD43vka7JOxXYz2jAywJMhIF9J8OjcZPB28yuoWkOy10XBif/maTJ
GZqfJ8b8xBBdGcD/djZTDnRrIjt+rxYKEmRfXE08j+FH7qmV67JeoJOAM6K9
MSKiaOSmb69pbjdl6XiROImwsgXHvKAxrf8F/ZGyHHXUL4IEp1NCE3uJ2U0C
X6is1xNsTXdXXEry8T7v+CERE0y0h0ujCqDu0HPTCdKX+b2QMMOuUPRxwh+A
QKux5+aeMfk9jgDh1UT4nN1WbLeKWcNuH8yKGuPFprzGoy7xp+jQA1R0UFlo
vx+nQxGh5BatfmeeOXrbhV+8dX0NEiYoZroiujRGVtugGDS5DoAyq1fi2sXb
jP7NlizjweI74ymEx+kPhllcqGQMvR7QYFOJKe9knsmgWV4R16wmKNdFZFMS
H4wWJWEQ1tMgp6jaBp4jS9x4LiS2DfR+9d6hgNXFV35oQvCIuTVeE1yCmhbl
Y1l1H3/uyETZNKfhH3Y66OJbEzia7J4NmFUjHvtwicLKgijYdy0DN+/UwKY6
YYRg3d7MIIo0i3qUeBMAFBED+9YC14DUV7l95oqInuKFVSfEi2lRAgPnFY7O
onBEW9bXf7RvdNFPWYsUePCA3twPNYqOZ+Ul4ycVutAJ/u1EqTSydL9aAIjV
FV2LYmu/ASmpuUPWiF3V35fzwYGUYEbyPJV6Mko09xN45WZcdsCvZQ4yvjzz
5lC/U/r1P1yyYkNix4wrlxhQlnbNZ1pJ8CPjY4DdytYQURnz5TT1ZvImEYLV
W1SR5tIeLOwR0R/TtNKGPJTc0EyEcLcaZUVC0eD/7AaEkYPvrYklxcVzcySR
aJMCbXdp1UQJ4kXPar9rCRbXHJ+QjaShnXHCFq4LMgodCMzFvYHCamNmMBOc
Fi2WpD9Q12n4+ylWheyFQNfaU1pkXvt2w4CqblWSrIOzdDe/Y24A20DJUfqk
c5iQWa7PX7vAIGCQ3ni+vWdwUIUTIzc9DhorpfkGtIMGPiEmbQcNdt3tzvb8
E5naagqIM5R6ITmxuJmNliI6GecKbwrLcd3ku+I8Ob5dwHmTYoLttS0Ej9Kq
ObM0ARt9Nu4zaGpLcqy9Uz+xGkQ/SRygD2lP8A+JNAvN6DPt78R72TT0wRlz
3jGiy2XAcvqPLW9GGAoAk+84ywF/tKYozZkpydtY1c+D45gUO7GKpsN+735x
wcbNLxhZF5I/kq8NcAJFqS44igmTzd+nmiie7muh1t7m541ncQp4vyz8YYSJ
jloAzjWPTPiZxhI9vZD7Xik/sPia2Z67tG8ekw0AS5RQLxJM0k4awqyp04wb
i2LGc54sAxzwqo1y9IkJM8PeR9bRimOnYLtl6ID20sfftoo3MBSKJtUxQolD
gA07LFBhKFGgSmey9jbbWNJOKSj/ricIvzx5s8plNTiJPFhMrGDWzIvnxzxo
JsLeZ9wVzYT/AayWZ1QMW+ohsoSr4Gu8rexep0x1TWuNsGGscwrSMrNXl5z+
wN5kyGxVIwaDn8IuKUG8yV4Owfsb674Ch28LRUvMhrSbA+s3s6a6CdFXgi93
4nenJCbvgn0AvjF+hzT6yDkT4PAehGU28n8ZvbOVCK6dVpJLCZfrhc5mGl3l
DZeQfFy+f9+40vWr+YXueX2d/pamWGwuPxynyFB8pH809Gf1831glvmEMhmU
VvMLn4DmnAaiHhjGCVpdfZmbdyFBygHnrjfazvZxNYY3oMZXZo5AbTdtiMU3
ox2xB+kW2XVEu1PaXWFqwwwfJmwXz+qah+l7woalWEC1p5LvxnWxLq6w3RLv
mERPhnnyreslBZleEXkxI4Im1YbjaWroN/75EP6MgUp+sa7nwf6tfmJuZEnj
n2X8XR3H65npk9HluBmZcYHsipuKuW8eJxC5LdTMgXcBpZZ8PyySuX8Jv8pG
3zw0xNqklenR5BPf09msRlnJ54cbBYIg9/2ZGAbFlYZLyQ6piCOK0KH/yj8i
8FF1nlZi0KgtcAdI9pBGvoIqdKf8HBWRtPv6aAKaEPGqBO+KlGKLxfcvDOt6
jYtW5ZtPpeSOqDsZOCWViCa2/NZIs7ynm2f/hQRsI4/EZou03kc17qU/BN8U
SIEzK1v9YH9BvTGIG+16d1yUcwVdLmwr2GYx1TdIu9VvjnuHbBoTAgLNm8ni
PqlfOUnyD/EfVzBQkZggS7eCZ3JLh/3DDCdFL7Ca9b703QJLyZ5afvkExtHh
E4SKmf5yoESV4ocDBGp4fhrU4n8imRRii4IgA+r+b4rcOsG9vdjqXKiUv79e
uRWHqgwNFCSSvfBzQT/8Z9MuL32awzum078KlCxWB5yIN5//fzlwOwJDHI6s
XltiQFn+jXCc86GbIDDR5Li5Esx8csJvk3Z30F4VyXYQeNxq68stcsnZ8rt6
ZrfVnpHcHIIiPp9rDj2zaN33HpHq6pCSzmDUKN2g0x5o/JjrTqvpTlZ2imli
F5GvFBHMM+HMFiZOGcSUDTBwwxCPrGgQqrDLsnqxcLowOMcyWdOKwV2r6eCv
8QvZypw4W/DuaCE5kbc+cGnpNq6/T1g54WxpqHEbu4jhdggVvZPCizYaIvKf
mnPxnItJBOevuGU13ggppTQdUZtA4pAxj8/codUsKv5h+isAISNB4sPpBl0Z
0yQ3BKpRzs4Sgq3EY1S57g4vDiQrKbZnruIOAXDMS461yRtrOZ62TysoXkIa
UjOdB50qNAA4mzKA+jizWneaQMOwBGP3Q1dI4YcWa64PPGdCvvycu4AtETWS
CQjYClwzUYfOx5uP5guNGLYYXlIieM5iY1Jb72KvvCzYelGJAQH4Jr7Zh0mY
AbSGku/cfL5yyaFesWA8wgs4Bp/FwNGnAu82HBEi4CIClhr1YLiS8+wUs9Yu
nekKawbQBZ+V36K8mWd6/M1pg2JqdMWBRdUR2j587+CJ7LMIlnELVuyHAKFj
Skw9o5uxRSI0cc/POesib/Fm40bh2Tb6UodXTruuLxZclvqz3fkC8QirJIXu
ibzAiBGEN/xn8T32/FDAJ0qzYbXGgQGVhd3m6FK8Mcgzri6NeUwZH/DurwS+
Eh2O1uwpDURoS5v3g/30qvrljGAXt8scVn/mxF/g0rrAtdDuoDDEMfdQBmjl
SKgSGlA1lN27jzZHf5JX/g+V3ihTZ0dRiWtrpcSL/2ciDagaKkkR6DPDAevi
dQTeayXCiHXz2HoqH3OFTLEktqbfVTFc1iMP3nZVJqDW/ejEL/bRXJQN/DhZ
R2Of/Dpqfy3xrbvb+5N5uJjjW81OVQs+quaNg78BOqzPUNBsXjv6XDEstKHS
I67Smf/M+eN0ioS3UrzAW1h1M9SkhAnsCkqqjW6aU9heiKbmXLZkht0wVJPT
vSIlwjF+NJ3z1Z/Jpodx3e4nP7rrVa695t7OeIxrjdHj8YHoYvcn34TYWd7+
BrANMUgQ7RAqtixw/4URaoIg1OfrISH9MkpCDaXGtDeykEc2i386A/QdKK5E
dIOtPq4apVCytkyRoFfmo+cfrVxHORU4hfMaF+g4e0MX8OP+qdSurRA8jkFA
rwTeCY4KoqJTPG14d/WIxzq9F8JGMaXoaBt2/6fYo6GbCSYEaVEeKGDp8I7g
cyDS+tYLjD/V6S0uuFnBsOHZkpvmJhnCmLAfUnkwwtF2uXvHlZ28nUzmk7nl
sM8HzdEpAlVC1qEF2RvWF/EBJBz+qN+h0byIAuut7IbNxoSdRZAiAwZiqSiZ
SEDScMByJ3hSYEOunqb11DU8DqD12HLsoUcAavF+22F2rwHWHNCfHYjMObs8
Bz9efO/W9QU5voqqYrMzCh/IHEzSL7wEyAkxqQp/Ad2aR2MfQ03x5NrKM4Uz
x5Z1zaFbIOiOGUPn9Dm0UNI6zDP2riuiWSy7tYODSWRcr9jdfqM7YuXh8smH
rlV52ZUyRmeqSfkWtsuO2mzQcG+uwpbBSkD6OGiOmFWhJ1QQOlgegdyOEOpc
HBlbqi6CUAab9p5EHdtt6eqGHOzGFzNh4s60s3FrDn5FhjSieremqjwxifJI
J4FvdQytSyB1e+HZ1DzNxcICGQ4W9qXEMio+zXY1tHNVfwyfrW0u1Ew8Adr7
WAiPsLN1kK75NyetY4UFZ9DpO41jyXhtW7oIds8aTm5ignwj78YtHxaa/KNg
J1d3EHEZMbww7qnBu/gG6vSevyJ9jyvnSHB8Ch1GEogdKe3dY6NebeFAIl0l
gfNRshMOMstn59eU15LYrleIg+6hh5UUCMO+RHLnac5HlDjC/p0kmOVH4KsW
Y0DTj8rQ5Y+Vaycu3fJp0WYfx7/gBW68eDb1t6/XV8lFTGnBlpV0kcnUXCo6
5Uj4Y0jTcjhmlRXW7JOyLQHnWzUIGLrDpX5NnAtSSa/3gEwLF3NIvr2cwS6o
VCQvXxoa6k+ielUdQkQzxlt8KaRQIMU1hsFUc7+jLOBy+4UOZ1DwtdAgK0rP
IY6MymGucjtoqAQVgiAZPde8ja1DFDRvtD9jJgKoLxgDmvSxh3DiODQ7kGrg
FHUp6mKPf9eIZwHzI23nNB+rIYvh+uF+IqqKtl4OMIgcucPObH/4ZJxNDM6Y
+p9wIANeLCz95gUZ59oAodVaTFKtrOrFV70o9kUGtDTBGXHwnGbA08rDR1Th
zLSCmNIu+mCJczY9RBgQlVJ28uwWBMx7l1J90uPMHiHWQheyXNjC2YgJCBHO
p2sVrFhBtN5cTxT0EGFdM5yLcKL8j9FhCRUia40C1R+lVWyaQ0F7GauSK5FK
NLXaTxTZ2F8oQNMI3M49TBIZWxJuEbzbiVC/retprcfUVVZPDqN4BjbN7Ano
ADA2tkctjFJENY7B10I9tbp4R2k+VJzsp6OY1aCATUn7qBhmLDfM9C9a3rBY
4bxzO+a6oeHFDfcfich1ICYtXUHDual3KSDzRslKZHy7Y5of4L90yNvQCZ9g
EEj0vzQ2kU0zhv0LwB2BAUqDLcGYpRmVF6o0a+/Gg54k0kBbVKSW7tRhknCO
ylWWV2ghg0L7cgSndCAoAPVWNh0QAdpoUvUIzLCyObkmZRsZgnyPYveMAp2o
+XepkumID3z/qtwK1dfyvPhQexkLSakBPG/8fRoI32reCd4u1pPt/V6R5EK/
XhTfG10G8fQuii9A57zwpbxjbXm7quoW+xEZXh7DqDuqrh3oVtZyo6z1fRDS
mbsKHo+KdmX/Qfuje1CjeYpgpI8fI7j5/bSJkTtMVQA6pCeaJm+MWr3iiZ7D
pMqrEL5hJklDnrOyDU3kFHliX6KGYDpw3H2QSSQYvJo9lxx9dMbwyG5WvhIK
wYdA80pwJA1ssetRm8DJ16cM4S7ovfqpY5trbcKxehnI/s+s6gOqX9iKruuH
ewVo1oWEEj3/R42/jwdpTkmGEB85fExCO4A4cn/8DR1UIXCBKngtDOjxAlLe
DpXK/G1eljqnjwOBvJbmLD9Qh3FESyaBl0Q/7rDQqmDRhcJ5M+axIXPE6rfX
HZpI5TCsyIHXLG5dtmUW1cWxvnKCzgV49i0+mgJ/vsFuYIVJkOmv/UJMMH0e
D2ps1WP6+f4+WBustYpdxDJyQzy/eEa5HVQ7/bNyy7dcc0NBbNeg6nnxGhmZ
K/5s+lUzYOjDlkDg+8h3Yov//AKt3qcOK6ePFR4VzGcsfwSwxFKzFLDevow5
W/sjrrnGSTJIwr+LozB8EFV56AOopNmy3y52NBSSotQe+QWKh/39DbTHB+sG
QTYyTI3r07qyy32+3SQC9CUjN37e5xmHgjyRR9XCQ7+r95j27pKcWsJ21C2P
CvZp8GwXduxOk1aee0QahnQVy9spJGuW0UV1M9kChDsg6piY6VjZZoN0lx4q
nn9OZfpdYNJVa1afrn+8xv/b61tK57qRp14UKWZ6lsoH7/GkXNAfrYi0mSIg
9Cy8gokvOpgT+eUO8wH2G6OsQOUmV6SSScBciWIMZnhUK28XIQO437UrUxqG
3ozCxVphWYA0bXX2GzDr+NS9DkKiwVT3l4C+JxI+p9GOnJqtoquAsINzPLRA
j3lMlTgOeIoZeWYFETR5NtF6xN2RoaEfFgPBMselI83AMNJQsYJfjqfIaujU
kt1EAG25InfYImkWMVt0lywOU7u44AESUzn3zKfv4NnBap0BFLAomktLvjqb
CQLUnKM7RCqfI65uCc9vVS1jcQ3uORDCs9E/SLxe2S6jdOTuM36Lb1TwIfxS
LYqOBUSK4RbhZDWVNqMCA60+NEACsLgOAgz1XhmuzMtIqy29fGegcZrsdjxS
EyJ+vyrcT4uD9BEu53KaQtZY91nBLpikAnuGbUhihk7q68OS/M91Eq+qEoXX
oA2/weCz9aFXLXIPDlqdXRrj8QTojaDboW2hHBJ1uZMAqDBEZRutbruJEdpK
AiZqSJoYIkRp5QwLqmlZQN5mRbrxXnAWZo6AWACPjfmuBldycHOyRB4mAr+i
36eTbQcVj7uV+LO2XheK4EZXMOcYciUPuZaY7z1Elhj/wAiI45Hr7W0g+AEN
nTz6/6b9bTZ/A/QngxDCNHQtyQ3P4kQgT3AaJSnbwIi4ei89aiXSv7o6xNP3
MiZJj/lVbe0UWNtmOJnkO09s+AHcswbFXWoYNHppf/7oma3w3RfRn0vOnPcY
guXSngWzXX53oq3hfeRRBcgfztiTbguSW0AeS6k/I+AWGy8VSCYtDLs9dbZe
dz11+gFsvKjk5+lBXS2Njc8zdNF7JW9CsWZGGPKdiucK9O9yfOrj4jM+lCdP
4xqfou0JvO0jNyUFnxLXy3PHfsdBJHg12SNOsuq5cTXOO8QSyCLyOZv3slFH
TSpscRbuwJH5NcvSKuQx/22pEXzJFCwGu1daPyADCMTNuk0EnyBGbfgwReAf
+thewdZihiXCN6K8m0eibALJBN/rTDBwvdR4++4E/dUloHRoGsbg+dM4rNQ4
z2cnUct87rUgMs91X0Cz43cGM6B0aDz6OYJc/xe/+KVA+dahsCi+/SNBF060
0GaZ3HciX4z4OQsMU9rEvfkgFHZoRl2zKsX9lG9EqxLomppI4feqpcFSomtI
98opo1d/0jCEhmp3juahNhIIivafbYAyRrNMAMChGCnLJN9KGwtstgFsUz5q
a4uZHhuZCxfqChLVPTzp+v31nhezHGwzhJUR8ksQChsKcLo0zp2Ri0ApP/WG
jafdphDH5skFM+7MNYWNohbggtckhpqPgVWHHV05g0vmnQp8A/keJq9z+jvW
x7Ene39MADBg2h3/OZDsoBYzutCLxduAqJNqYdM8vOJCjg1KUl3iHnQ3AisW
7iVlQdT4BAI9Si1u+SbQudpL7CXsICpqRlbm2FTSkwaaceK5rSww78riNpGL
EGzcc33sbx3m8M+FvDWl39SQxfg9HgTli3bPHrsIVRyM1Lz0gyCwjLwNkhCL
hZucJcV3L28orC2VWsdwva3Zo5IZjiqKyA1dInjeMVrZVZv7FG2donCvnYU4
K9ah870Iyc0G8WyBT+jy+HpNLiNHlvmzlK9qcuVuWRsZi+6o8BjVf8spL6uV
jIjLWss4iyUQ7/8Ju2jIZErzJ5vEsYJwrWkrXuQb+4pmbAC7z7P4mFojL6Kv
+nIzp8JbVrtkKMfuh0tSBj1PYTdAtlvltJZSXvZf3o5hFUsKLTKYFFxXUJUl
SnYrVM4rwF6O2B/bPp95+DBA8HtM1dif/LyRrPRF0fLi6Uy7Svr/drTvzsPe
EUlgEIa/KTTNhfjbi0z56zOh251+sARVRLjYK7Yh/iSqOzFqi652JjYvXOtg
lugqzmWV8HwrzzPA/xM2p8ufAOUieeFKuvrKYaYB8fpKGBDcmK9WF4c6ljb+
SZN/ZM+ETlJKqaRlqkd9mDZM/mhYod3d0d1Q9lzYUpeqftLeeRLDQkW+CBTo
tVNneJTUZaXzv/TZonxwN5cvoyj9IkUHL3/h+IldeuC2D6wZojZxDs3znkMW
q/fesRZBeAmOg8bsn29RXvOaQJvrhgghaZFhuj4sngq0Hwk/A0DHg4HU9dK8
DMDN5yfuqmPOS7H+8fnmu+KUp5QaNeDvhDEE6YwrtB8ERPNeQ6Q/5khzxXhr
NBBkWPOoU4Sx4bmaMP+KP3KEOt/QWboSO/f7d1W5rUNEcr3M0/PQzUD4xKK1
jObsZ1Mi6io+WFF6q/F1ATW2ey8nc81RgcJKd4PdeKgWimSPGZgVPC7iJ3od
39RLuOan9ufvwFUz6j4PdvCd07+xoG6lzo+t2iEACRt9uD+jLdEJmnslTHVA
/ahMgOgTiz8x1qfHrhjAN9w4aegXzrsVsgvZycqhgJv7Ex1VSIvVtVN+D2+7
I2rOa0r1fssCUMCwHDj9iJAaPmrz8YFMf0W5OhvwOiWDFcy/mAJ1HoSCZtyH
t1j+FHVOomk+vjrRRIr+GTXlAIEhO8lDqtwmH6TCJUySRfwCtQZnj3pR453n
OKJ4RMsk9ryFrMQP09Gqhxp4ML764FIOQl6qcr6HRJIgOGiiqyd7zAh1Jqp5
DQj/nYGcXyCJnPMvjEXKqRuZmpdSq+ouDfybhcqMiWB+ar6+jbf1qrm1zk6B
jHifaz6EFi8NylKNZdl7ThefekgvuLNQTd2siGq5oLVETJwS5RcSiMHzaeF8
aaTqT0McRf/yN6twdP08z/+gVWgCSaDy/M4NUJTnyJJwFLPWn4LQtMTrDjL/
GxxT+W19S5s90JsH3IEWIidaMVLJ/V8mn3SyBWGnmz9jCMJcRXLaYYGhrNUu
9SESlGAQ7rH6ijVoXzMTySQb7FQDr8/+TItc3mGtwKpz90ISVDW0N1YSmiNV
BR9kRrjMpXRDgGSvwbMwvuJv+JrhhlKkcVblmA+OWLLTNBVJ/wezEVHJfAO2
sEF33UDNgYnHHujzSdH6WELEQ1i2CAYkt2hzrK3Wrrj3wB6z1NWvufjhC49P
GR+WxsnJKp/u2s5IeyweVs22IZNpuJItAMV+bYZMtYi1d3vIcsmHChxM45nr
C7j7TJTQFnLw+q1zQDyC9RD/2AWvyk9GAUu+TjAHr79k1yY5+Esz9GlEBfgQ
rDzUxtsM+zp4ClQsCRrlTZ8+gqoojZ7UN6OlFuuKd65HpkO8XWyogrHEBWLG
XhYeuAuwkCN/uAnUsC+7DsQuxrq5Mz9blyYpG7KhMB+S1xB0FncPOqiItOpj
YUaPOeObErDx2oIc/7s8dQmSXZKkaKP7pPLAJ0UUa0PtE2Ssfq671RwuSQJG
zBx4sH6a7ueZ/NF8L64Cpd9V8ra03GV5HQuIpkXEfoSHn7ON/RddFfRX2VYx
ErZcnyZAKpiq68BaQyZB1FtGsUot5t7XgaDpJIPIKd+gI2WhcE1C6XdKF0ro
ZvZUjG6yRG9DQh7sOGqv3EVdGb5JbBGUjqOcejARdyaV1cl9eUZV5MNAOZ8m
/MI+zXlg4RjOq2vcSgXUTJXZzbGqNnbftCMstGb8oNtSUBH4Zwej0LfI8+Ys
N2iOH3eb1sMH2D40xnLJT0qce1oWhyFUU3xOlKq48QBX34TlneX9++5A5D7I
G01/TM7xGjKqj1l/WNLBr9vMHmhZE4TuSw3OFS+NPhtj/h471mq2MqeJGJk+
SWOQa+gxqMdxfvuO4KL+PVldWrT8kfJPZr4bEoMJfdhsOizxaQwwwNHHLW80
fap37GQSdvwHVYs0s8TzEiTSPQZBDUAznoL+ELYcoyvmgZskFlrWZp5UrQ67
51QivoG66yPBzVSCn329QoiYbb3C+REc5EN1yTCKOHz/hMfVRUGodAOZ766X
K8jQ7TlECK4AXjyujwKaHzttJ+RahOHpO9C/M+veOn705cKdk0CBy4sYFdq5
/sUykW252hJFo8AE98GdLno/WlTa3ydbBcbe/vwlQSi+aEupA0l2akJLO1xv
SZwEm6UmpU9cHNwwB4PKXlWfgXlHggI0Br8GAGGYWYcjF0RUNW08KNb8TQH2
lv/g+ZM/bNUeJIjs8YOU1DcEj4+WEjvTvIOxG70bdIGmGSXVqaLlJ0gmoIWA
yiFGVuNwKeZ5ApxVLf6p1M/NAwCC2u/sFytKfueve4GRE2lT2mljqNVP1M3f
jHund84xrXr9+Jc7fK5XUyDvtu8bt0lywZlu/wG/MaFkCJ1sFqJBwe/McPdZ
9qF7tqTJ4y1i/X5dpSNUmNpjLMpMOez/NERB+elREFgy6ipORnFhmYsxVIRq
mmJyvdo79vQ/aajEviT6Mm8UQb0ifqE7rE9tSxsnPEBB0TRS3om3mNX0QXHC
0ii41G99nAx3NZVVY/1erUk1yg5sz6MwRMmCHcQzN/Fjl9ZvH9Xdch+qPfvn
u6yShTlGu4KDxVfSghvfRDqLDhdN4laE/oJR9uuSnQ+IjbxIiafxPZCQxVdV
EIjKDNphzyW2lMJ84YqUIJyqjhEt35NbGmVcTli7SHJgrjFccl6zDxsmI34D
sFVLkiCZ8Nwon7wwB69IHb4LOKXT4ycvRnkRiGh3OFyyOXrgDNF/cHPW8dUW
AhWygvM4WGjwtdu/XeIZuzoBzdU8Yps0mI3p3nmjifv8wO9M1yrSfCACFgiU
4N30DvCVCB8KVGW3aZfbkfjUQ3wx9lE4Y8xrV+vNkETwZQzxv3xuWO3Uo8hC
/ZNN2xtfpCLYg91mC7w2UXEkM2ZfbLmC4EGoKmRWgpse3R3yarHTqYXAh4Z+
agtcz59qsIBMcumu8KSRASOKLmIdzXPnfgju8Si86J2cbMLYXR36SI8AoE5G
dlQN6aBMYIxB42NNcHhobnE0yLZhdtan1zFsHmxNr2Xqa6qxDD0Y7yGATcRv
p3GDhNaigEYn54htrRw1GVBc5nvoA4MZWTTelVgk8aSdMY21oD0txLAIdO7y
qpXuPKp/YU7hvlQ3kdEBiavuNKlPmTB1lBB21ZvuElKqrkcl9HDwrbs4Bhlk
Bdm859k8r5yQvVz/BhscqrJOWhHwvkFYgJv/JiQstdKIWjJVqGZUsPO5R4MO
YiJBlj2JLpeZtqI2E81CBTmLVqZVAL1N4+Vcs2xSGWp4CURWwWloz+L8HIkK
ToxFOTjjcIIyL8UMr5d8yf3v/7b4E90JbR/GEkQ2/TWr1OrlbAdZe0J6nLKL
2XTraifct0p4d711XoxO47MyaX33N41RdXE2YPs8LstlGWHyti8tTdfOszkp
Iemr27E8OcKP7iam7zaDcrVDqQcE18+CrumMnlgbX8AM3t6NoIZFpC4Qq3g6
pqCxOFLtUEpWOZI+KMl/W2EcPg1gMb7Iwp64qSdXeb9YESeYHQTa54O3OYrG
8Yi4/a8NWztDz+ZaXOrdXAOXWC7hxn0OCM7NDMC0JiTgYjp3M4mRj4atin28
QVBxs7nDcZTpYHLJmExzLJi+Z+iusCgCA2zTHpY3ZmAift6klBt9azcgAdjl
M5z41hF6H1rNAL29STE9evWldneTEwMp3q1N5aabE6PUhtqzLtAM63PZtRY/
pNLNosY9XOCivNfhxeHJq6IDp9SBYcyvn97CFzt/Zq5xUtSVmSkGmIllXwpK
Vc906II9BYBqtcG5wK3JlX18ZMoOORKY+9ivxRqqha1A/VWrZjtH1PoqvvDg
Q4LkB3T6QH0qIJlbjuba0xkPh1e97zwBpOesmVTr+zBWc8qDVGn3f3jNETjv
2f7WG6A9yOxJM3uf00eTwCwum0UVM5fPQF86Cq8A6ydCCu4W5+zF5HCd4tkt
QBVyDwAOlssRfplxgvG9WzIQugpjUKAGyvp65AcqScftKikXFAOaik9FuxKl
uxXw+2ORY8PUYxfVBtnCz4eWogZevHh8wTGrn6Gjgs36RgUprV4KfgueCwtm
nvanVzIs+SqNlogmk/+MKhMR42W8OtaCId34SiPVL+Y9jmYD7hDM4eRfwlhP
B5nJaws8XWAcJ3apHSQm6OqITUsOvZGb9nVRTHRVIT9NLC8ch6sCygII6cmT
F9JPM8kG3VaBe3FvuKAoWzCYOU3T3MYZMoPUhmO7/p7e2jjJSFDS0SVPE0QU
VZbgavDD003VfkuJoT1OHXbs6S4TltFr0Pol5krETyzAlam75x+wVSrNS+q4
HizhMin5umXt02AwA1Jm+8LqTXkl//Har6lOjkdl3QBrWmiTY9qYjVVgnKSn
LLahb4RUFh6dZ2PvNdVaO2zJwrPyBBi492kUTLGGoYkKnaGCmlKqcCifmNc5
Xl2lrLouQ7eVBD/zqyyPqVHU35DGrGcU8n5s/xSlNVAJD7YxOdklXVKZpeJG
Fgx1G3HYJcRrzA1Iq97MG6FzWkaZC2OEcL+H+YxW6DV1V+ji26khtG7WrOZa
gR+ln1njIiHLjFJWsmoHD038BbMDVvvrQDaxU9Z27eDMZaWivCSzdDturzpD
snuFr7gbwfa9u6H9fhgPQMNlD4lLT+fhD2bVrBLesYHVU9+GigLQArwYPzao
HEloB4LbmD8CGWNjA+5W1+tL99BM6CCNsBc3FHy5rlzTRPoUXy/7KjSxwo2+
2zmojluPqlqDV4UgL+YfNIxK4UoxxJBk1lbxIyw1XPY+C+hkmZm2rU44shxL
VFDT+gRdphLLZ7bd3aeXcOyd7dzDFHDRI2v4//8YfX6/WMEamJMK4x+ZTBEF
nuHGm0gSy0K9UQU5rcjtGsIKTR/6ewj2st6tzlkXlzxm4AmVLdZauJnQWxtV
guk9rn/tqdCX15tfx9ZwnjkEd7Ct9VqiK3ZSa/zg5jKIO4bROV/dD5PQRDnY
WKzR7aeCLEUbos/NmyXDolhE74gr5SI7EL3jvSiWlBYoJ5nN1CrS+rALa3Ce
Qx/QVHXCnIMv2E6PST4q8UXJ5M6oBipX4L0+o9rxd7XFBYW73X+TFSsHGrDU
99JnqXbzEuH61C/WfIQaITl9m1/BWlM7FtKVwgU7Lwr9KEvxBISZeaY5vMpw
YLmGNLxYMA4Cqc75SkFF0gjc/HQOcIpRRSb9W5w5mAQl2RM/VlsQQD6EB9ei
mfdGGBUj3ZVjcz8JWwmGuj0bycC2EgGBAF6ZJpQNxWYUWeMGxTefzxB1kkq3
bjhtFXNINbqxMOTPclEPqwshxrIADXS6fiR/fZxobcH0n+pLT2Pf1BujdnBU
MDbu3h6Veqt6Bo4AVoWsl4OgFNcYAJJaxU4/MXdxtrdUziVsYNzMQ/VFFQM0
9rg/NQVZJCR4gjux7WRgxzoTndrTLssdBHMlufBNM2XKFwFh+i0+l1X1nKUK
N1/+IM/tLx/+k6hf5Qcq7fO4xeusOF9TgG+nJHSH3KNx5fWi8cPJ8E98kC+x
cs0JsNoRA9kE2mTI1H7dkjepy/Gdlgy61TiXl3qvPmMBGNnXLnAbxUXviP02
DIgtnZlkKHM8S2i8clsncFSQOP8FvBg/w17tdCifBHvsMyIQF6ePIlADbLBE
TCRB3wCG3pB+4i8nHzm5hda9c0gsK3cUrvw0cYDdryfCk7eXqxnfpMepU45w
g5cdRNKtpfXpTQVzF1E6eJWzRWIDOlD+iL0W1cqA7MfNiHzOaMvSGyOHJ9g9
3tQM0c6EsosZjl9peTSMaydwrZjMEOIUH8DnkmoEtsxih+ZEJyMVlcpPUrnV
CukHLYb2NIqhDKasbIRduhlTgtTKAKHkaP6fp3dHrU36IE+s9OX4+DxL968t
TJ8EmDb00iFeIAUmKVhMOsZi3KuFbcLl/40QfdEyNMqQCaJeXcUGWxgRAypP
+DLR7VErD/iY6RUzU/3O3Q++s20fLYY0Bg+3h5HhJpn47lGSrSlfUmdMKg4+
X5yNg03DbkTnfA25t9pKkd/mx7ouT/OSkUT9/RgESzsud4jnLFalOlJ4k4Sd
6Otck/7LLs7c107a8a1k0JNX7nKQrzQ5jEu6bKRdjzXys4ej6cyEHOL6X/GD
63ndn5P/tdJETgPgWgiyDVpgNp8gf3EFWKn46afdHllDR2vI0IsPOPHw9Jsa
B1pf2Ys9LgQoyFH1+4lhxqNML93IixyJWsnGptClEyvYae0glxlFi9rYXEM+
7SCLPxMKzMsbT4sdXoAjOptKKjbD5I6k4IGyTuNfPjYmvpGzltUiB5eLUZOA
CdAIJuqjPovmiuU+/LY9pNynCg7OrHeHv3c8VA6ODG58oKmjqPhEfau1RoEs
kQn87awwfp7GohsiOOjbbscJiPtP9m5SaourjtBPgTxQLFFY4Em68LTybClm
cCy5/QCCVFMz1x7t0rbpnCvCIdNzJKzrDjfyfHyCfIxE4a/4xnGP1GCbeWmn
n6L7nDTojq4fwVhMoePkqQHIZGlRpOpjY89Ave3KEtipno75aWsUuqzs8Tff
p1agqQkeazZjFAgerd3CKh2hW9G0IF1yHhYLEkGIn99O7o1JCeZH+H6baXzk
NOhI0PCLjrkeHZeU/2diDtLsotNZ8bmk46FHIi9hUD84RvfwDIoGUNWPpfH0
WC2hxp/Kn8X7s5Dm2tMuFZplasyXSKLdVelHKLepld4foq47wXs+f0FVi0TM
vYvhPx0BClcdZr6k0nrPRbIrED2r/0UNnheN7+/NvYCh7ZbYKjcZnNEN3vZx
0WoLjE5ehXzbhsX6cCy8DCrpPsRxOImsf+dJrjF5N7+GY45apwBxWXVo/nhI
zE0iaRgadCaaHyPj8o+t0YfOeEX9qoU3xusT/df9jBqrROTImnLnflhGN8R5
eLBwUOlhvtn8zfUK9GNqkwoafR/9q8sKVMhz2+GB7CbUYhEXl8vDBuyF21E7
q3yrMLjcditt73ZQW2NOfRHmMpgX/GO5yP1of4VKPZ5KyqZWBFpZWSi7r4xV
EuQaoSB3/4aX6lA+fjCBRhtWOH6Y44ecFAcfZ14205EbB5/ZTEiqNJN+/2wL
DbMABnzgS3L6pe5WX8KWedwvDHymWYyr8T67SYHmUPDtsD74G6Jl2ObGtk5f
J8i3jSrL1QXnWBQWZBm5r0qHmjC2eYdW7aXYY5vRpIW7SJqz3HjXlmrKClZg
xVHebJpPgzvFdkpfTbuDp7lBm7EIVMT11KRcRH3Vq947fIYVWkl1xgugl0YC
SuWgj0SsOx9dBDY4jm5Sg5HDhr8594wJmtDwQV60/U+lDQmxNMwrMcnnxSun
ALBLy3nEYzwBQWgsymNsphpwd+bq8q3KgKiHwq7+cQePch7O3LzBeJHIm+Tb
j+rgMeewyVSwaXvs67nUPSXqexjkVh5OIkVGd50gjtarptojMlVjiSg3uctu
vOCZR84wlRI/sbht7Gsa1PomeuHEKqy4PdJ5WZHNFJMWevO4Qxo3obV2H8db
cajACobiTKbbzrIoypLVSRLE/Fc2iyUEn5Qy1QM0zqXWNRr6TQ2oMMkuU87+
onAvWhpl3m2hddY7dBGj3hGCko9zi3qFO4+eU4LlyslDqq07rKeH1iJ+9QBo
8bqDRgOM9vyakTIDWC+vq7xPPfIVm9wY+BYR/dqBYcChGzk7pya0M5DcmdDF
lpQRR55QxrhG9UdECUE2uPafDUWoa6rKK8SNWagCo9QmXICGOAlwyQalYTK7
aS/uGKzenMQhLFlYzBKRchX2tHtT9Q6QoKjcuhFQG8qrP9USTYL9n7PPH281
1yjdJBXlqPfkZMd9Uz71LYN8gOrwJnX0v862WEljECD2kkNs5pb9rLdNqOGl
htBFhQmjEtzr4hXIJj9c6Xyddzkgcu6oQ3S4dahHV/xJYMxXvNP9Eo3FPumM
hk8MW3P6DPe3s/kpI2gyW0DP0sk9ztH4UbbLGFq4IKKrD8lL9MENkCsskfg9
Ic7ZkKrtvF0FFaOYZetBVXU4nW8iGxRFr46/AQ6TDzn1U0jqcjuhOf1ZvIIq
ecDC/osUdu7GiBu7L6+fc5ipZKS9ysFfGAz5lWgsRL5e8Vsey/G9CBk8DpS9
5B8EFjkSfspxyfxxAOoWbBWDPC+1aKyTvM/Y6U8jp4YSvOD1pHBxj0VZ9DZp
8abF+k9h4wTDMxf2G+vwxJ11n4KBu0npM+Z6RLeVFeUFPnaa9cLPCx4z1AD1
qqwTUZSYO5FoE7uB7lP3stueGOfUqcJTnUgdZtaXPAQZYrcidyePjDPupP1V
Vg1MKFpVH9qGcj3VOTsuh7MxMwQXc4HWqg5VJmctOv0G4wg1VnMZNhRIMI40
ginjJCfN1bTQmCZKFTxEmcZUFfof4prBY0N2U268zfodfWLklJADy8fcrc8B
rFajkCcjY3PzSU9Vj76j988yAcJI4IuQM+ri2AYduPGKV4dqiECOqRbgD/0+
zQXu42Skn0jJeDNZqpYnBSndqCEu7K4rD73m+eFV0R1hElQjSBO0WZI5nSnE
RAqFB6aaN5bY68iGLFZWY6OykVMqXZPB2A0TXNvGhg+xhrESC0Ne0jT75Xmi
uqF+iWfeHLSfco23N39JZDtox/c1pmtZ/dbvePRzv2IeilEliblkl32QhCF+
TST2+7T+Mt/OBJr3ElBPHZPoE2MdS0cVnIwBLYFlHm+GJMr0oqhSOPZPJw+t
r7o9H2yTJa7Gu/kR47BfXWZgjkJYbXnrg2r34VwEVWsB95jlUQrdfV0z++oX
y77Tf7bKB28iCI+3cilyDg8c+dFd8+ImxE0ri8IF2H3eVWMA/gjpNZZYkSWJ
BUwk9KL4tdifB35tReXho5eyia1OLFW5F9mNBw69VG7A+tIuxntIfJCO/RWa
qfMu/3hzuyW2nKdawTDdLmgld336ipl5knFWTgxLHuUtp5lNwQPaP8QW/ZDW
zVseRDeTqFFSld8aaNtatA8FHEwwQ4jgonOBLxxg29MWjQMLRnx3NYkNbGQN
qT2BfnBNEzy+FHFdAmDLavpcfAfruR2ttU8h/ZSUK0L4ocIv9TfG1n4cj4ev
0akO8bp6x/15GMNZbfoTNykn4/zgoLG/18WJwx9NwuuuyI/VoLzvmGFVFpDd
ONxQve5Rnpa4nAZnkOkR3/jCyt7+romkQHffhDRo/pP1ljzUYtxIyIj3+ym2
gFlSYb9j+Ip0594T4q5Vkp0twapL8g/stXAppxiik0+iBANPIi+WqLEvF9Hm
eOVn/7oPbX3ymUyJ3nrz3C4jikzRg4/oe4zCOQa/k7reZrQzmoLiE4C/B+nO
g1ahORWcOVMTHoFx+xEqmOzp12ujas/t5YAfMTMgCrEPfaDNui+GaGHSf1tq
4GmQ1kiu8ndcLEWpilWMzKjR+fZUPCliPt8V7QLQ1zmnGA0BxKEBnFXcD0U7
P3uQRl2Kvh5FlwTRUiHfkuRqSMEvlWpC9W5Svg2eN9/iTZFIJ4cr4i7qoveK
AWM4QseOHiBhIDWbL1IMO+zEid8bKgCU9/x7ceTXaYIm6ilXZIO55Ej+AU9U
BO9eXzR2x1qoqfsoNGwGSvocU1o90FKnVjUyIOyMXE2uNBeBL/9qfP+Zu4M4
tpT4JiGpAunhkr965lNG3fKA0ABI1RRCBRM7q/tnLu+jfxvakm2l/WZhuU6h
x1vrd0joEzhqyId69B8fPchrrXfKG8Z4634MMsihIvvbsxHozfraDdz2Dh+z
Bs0e+ntd2XI1viX7JH+u4+kcQWJ24bio7kBNDIu6tHju9ucE+iieeDioZwGM
jgEubppgBIiBLJZEOEYBv4z8EXB4xV1EYan/vX0f8+xp3Pn9V18/4uawIRie
C15qljkal3/lE0lrovyYzhldPA7D83IlS+E37EGcxxnAvWWP599KA7Qw5EQb
Gd4hgl4OmiItRX4rzqNUxoCRl3u/XSPNKE0yp9jZ6CYbX5VDN0fTz3Wu1v7p
aOPdp4bpADGva0Q46eefAzPKMvLwIsO89wdjeJtE4nfXowWhcvlclSs7xS4W
3NcNKkIjQ9Rwj2ZEH/h1oJ062l2gz6WO3X5FMwN+FPu3bI0GfjxKSzmXcb3T
47dPNpTkriIoCiWzsDtjeyeo2ATk5t8NCq4GQ8IrBKsi5OuYnhsxKuOU8Zsl
yqZv61u1OyT9PUF+8kN59FhcRQKEGCUnmI6bWPm38dcDn6CisuGGEsq+Rb6g
uhwtfUYz9LwYIVPw8e8zZouu+46ZngmpoOZkxZRB7cNMMx+/n8DmMxBrx5g2
0skbcS4AJhsDz6XIfjWLFp09ClItVcEvX7/ZJomQnnNKOVw3kp6F1bPX5xmW
2v8s7EcpXoYHIqWr9W2ThoYFs+nT6qiVrOiG7CMuNo+t5HRJJ5xE0mvEUVVl
Rg36fkEEV+jvLI8umZtpODNFKnRrkdT0TDIDYV70LZuG7xncHKGhZsPlygbN
jNZTrU7CByqj5io1ioHvwTzS/MIfX83aPa1qkKJ2XFVlC8BPCxL369BPMeHW
mZZKjc3DtIkDVHCU7JIpThSbxFiYKHn5TYroxP9dqPkQ0HJ3EhDHXCwzZnVi
Tw5dmsvn7xeeZWvEdpYItHs/DfNlvechFaG8Z9NST15YH8M4AVl2mV3i7C6c
ksqnAWTySltIGzKkmG6XqWOm+P+Aa+M35tiDf0RjW+T8LNx4711pIe0c2esD
OCWVq7bMPnwICaCwVnVd0zXURb05Q7uTXPPwJR3spU84j/JrzI/vSiw3SapA
DriBKsCfhnDic/nCg4Irln8/HhPgoo3BzrVLNwQZ0QdeYyzOeHBVnz1oX/hn
voORoLgDmBc5M5w2i3yWOBRud5y7lFL0k+pysHu1MmftOewmjuswuMnE08OL
U7cWFtuQvfYmqz800rVGHxOZv426MsxAlKlLSarmQWq/WO5nSfak5RkiKEIs
AnQkc3+t40K8/1Ea0BH8LWH/Qw//ZO6aF0hNCQfk6xpvePgnnNxm/cilgMTO
i8Y7YKbbyQciw1NPkPgbPOq3ByLTBRgylDu/El3y+nRPvnOsWQ+mHxMO8M+Y
5Bv+fI3lNjN2GUknCFdRUioInpHBeOeorCy1qq5MbUby4wd5Uebg0fB6ls0M
AExKceq/4coYCQThtpfg0RQsHZmVZ4VDoX4C9ZfuA6K0SjyjbA337BBB7qLX
nx2giMhxRNJ8gVs+2JfjiLgSS7vWi3q5dhA7cp8Y1P8vYDGHMo61B65uFOeu
vsWUWgECzEvG9BYdqJhsF0s+3pmmc25z3DFrR7QKYYXMpRm7b+niIjh37h+Z
P6edXE5RzaGQrrJhOiVrCBgzBVRO2BKQfF4jngu8HCQYmP82meQ8uu5YTfiQ
jaXOllkzfUsLyqHwIXIj/+vkdF6Dwu/pRhGNGN78nB1hXmiOgAO39CXfggev
p68fxh2KlSdjCZBHIMy15PIsF19F3IThIvBUXUnCh8a2DpuDvMY3i1bGf1zk
KSpg3wkXpAA+z7pqPCaxwXW7/NYqKO4jV7L/NERHs+jBK4zCEBrtervAKlxQ
u/XoxRq5txKYcM+X0NwaWSt8U4sCMFX6/cM+pUhRdegqgjOkvh2Q0B4DNEqU
Hj7JkmwLVWMBrtptotr8yr9qwBJujZAmXXjC9TzVobdQu+S6UvkLrpY9Yx9r
mOmIAN/3COX7Z6j+FGs3++bBHlw4kA4/HyAKYYe1YKTlHhhDyheWHCeOqN75
cVjWJ998euH2GHHpsSJD3SPgV+8k2OCGIA5y2A21qWi2JAJR/zSdxqQN+l0y
yeTa7Av5bUoqntm7hyGbBXrttEiYhSuN7YMjrpDzNnjLvA8qspZuSGPgKKmZ
VT68eTt9Zn7h0TQgjQQ1QQ6FIKY7DhkzFZOsf/M+lfeoMG7M5PCVmPslbaUs
bTOtxwQhNWtPy2EbafCtPugJSOpLmw2pXnbdoPYkDc8Jy63qE0z7IbKvEOjw
kydzu/2s40/07hfAWLKhbb3IAHABz1varoxd78S6RvmAe3ooQq8AsBJcFAnt
4QdE96TKpTdN+zA69ImGhpYPodCGnVbsHvn6ooQdYSRVYhY1q6v3+HxzrUfa
5auz6oXVgQ+869dZGKFwCAJ/zJglzXvOYGMJWxYZgABEgUIsf8MuPNi0Cl9j
hzuGY6iBbpxn0VWC8QULv8zCpaXb+gvg6BV9XktTZF91HDpWpnULRcNmJ6ld
m87jWHEl7aa064hfioB5AxvHlnAjNHVTeLIYY8P1LmNJ+4+TawDfzv12WKPz
gkwknS00teFwMY3bw4BiLs1J3jSo6uKaUf8ZFs0k0x4GunhN4bEkBRS73w1u
SGHm83+ToKA4/QnvNBZMwi+fV6ZsQTzA+r3plHa/2RWnUHh90zZ5hDMCNXjZ
HYCDb9Yu9l9E0u4wERjVe/SAXyMcxCUMiMaebcsSyrAOwIzeWjR9bZqvatZg
Ji/Nmeab+xb/8jkpxkeGZUXV9QDE3iyuoOVqpgTEYAtLhGN/EpbyYxd3rWgo
VWxR5kAbVIGpFxRbQKeCNef28JI4C+lUlR31l8FpvGvSIu2qmrqylBRoPXGg
40wO6weCxTEn7y9q3D0HLhqdH98mhCcbXfMY13rmPSO77JjLx+6wJh4AcLdP
Ya7x9KBMybp7ByjXsPsB+yuzz6YcmBNQXh0L95jTk9GtNkrtSG1SL2QL0zr7
ld82Q5XdZZImcBonF4LtTnwGbsZxMvh0niRtzQthOVm9aImOlerC2xP8ZgZS
ClU3YOQQm52JgpKQs11jwTsomVaGwthHLVqTC4ljmZ3CbsqUQEsAVF/koi7/
G7CjlNV4jd/divFLI1SuwyzSUHD6kit/6bWXVTbYN7x9dNGcVVlGlsyW6cn1
xkuU2DmAWc0GBUjs66m+ASOCneCIm3gkc5Apr3gHVV/FiYdcfsboB7QzyW1G
rLPmRI3L4eG58tDIYPJtj7a9fdVR6LaHkB079U6ScPFLH0i4enFLcDQJQqZ1
d3dtjIdqB+wLRODdJIS+bJ/j4sVlvZPJ3VRxnbkbHqpiQUUDhubaO4eAkfml
xm/K3y9khnzixCbhc4g6DwHjFHVRx6x7CU97tp2XluBlOyg1iNQdKnFYKVs3
/2XEBAPygDfTinprd6JhC7P5q7sm+ygq2/e0CU+Te1+6Wq/SriHh8zRXUt/N
sQ8Kv31ZWOlPQC/xhKnFAx+ottrmYyMvWTLKTqdjVaJRDkhvEoEfNjNz6Xbn
PIA0ds97loMYvRC4lLAZkmgcKS/Vps3gXogvAPjDm8I+4PJt4mK2p+2MML4P
QNP9f1XGF2ti4nvibv1P9hu4phEMaaw2azsjuVkBh7OHzMhK+zkEWR55qbEz
b3nVEhAtwEydVr1ZDyNqcwW8EZ5bgaV6LDhAS8dQ4ib5VJaGNZX/mLUChDL7
Qj36WICLrbu/kv3Tl2atCZd7yL5ZxaIEoczmjgtQMJOjh+va1vV+5zWQIOpC
bl8VrcOhr48OiIfSxh0ejUWlZ8/7pKFkcvylQDQDZQSgsvXEgoPdsH/lLNrH
TbSHWAVNyo1KsPoMyexrcr4WGWI5JnN+TvXdWFSBn49gfsYjJz18OglZzykj
+aECWasQucd1LZ0ARiiyS7AmTCBAHVIyDPCobgJJkzgvDRViWVvy0Rqpnq1Y
eiNutkQoqotsN9IdEXbgr9HvClaGxGqV4CtiKGnbij1qdZaNbGLcxSO6ZONK
9rtfabzpC74e35RtzOHMEwAxkFf2EKCtyndeTm+Ms6fqef6JlBkm+UctYp73
tQBfSbYXuX0nqBm7LNM4YyVV7k3xSFDSFxZY2i/zlI2xfpx74Io+9WyAARWv
giMLYmG29uRtIY3dBCM2rOW+o/DrS2S4eZ3qoUY8AVoAVfAejGeRIEcg6jeq
BjkxIxPS5PJLGb/xMQcnoRGw8tljTpYDdKZl02szUIaySVZa1aU316Tgg5Sv
B1IjXXmc+01LCYnFSGyu2DF3B9MhKqPGoMv1rpjuTdpuJVYS08nXAC8hZj5c
dTe8ejkEHYUs9mtZFyqEvdAOgOKU+2PiYcnrxy+lGYEzBw6gNd1DmjuGkW8L
h0Z4pF/u6q878QnRgF4A0v4LkxwJS2nNzVibmKvlWuuCCHI2A7UHVehN/z88
QaGleXP3aasLNA6stfSKb9IpmHeUbNBLGBIzhhURQw1tOJR33fzEAXLsBgn7
AlNvQD9tJU1eF7Ys4k3++R2aLDnTGpJXzOoTkMWQiW6cmCFXb7YOoBj+U1xs
cdz7D4TSl8lPkjmTvym4kXrgsYWoL0WnBjpjy3zuKSnZSm61m3SrPsLSwUIB
6BrBQL5KFqnTpZRBiVoFjCf9lqb/RU96hAXuVpXFnN8cwYL3rXaw078FYXc1
pzYFqD02o6JCvyUqoXXD/fxAC1g/Enl8/XfCdjKwUYZP9rfGdyVEr5wZW9vT
IoWgoVg3K+Wp4CgE2+1zc/rt3MrS5W3biAPfLevHegi0wD8Ds7ZA5CAo6VOa
AXA2rOr5osZp9zr5MVNJutZ6JFeql8VbyyfBDKuaWUExkNKpUnUHgJHBSGWb
/XeMf1ylrE735WwYSrjjYYNs13RKtGMp8zvrsh00iSMOBaiqOcDQO7OgCvxL
TuqE7SFDNFd+ndhY4ppAE68uK2p/ZATkvYFxpxUWslubi4CX6BhGIkb5D4u1
Jh60mcbwSywiiHzy6HjRgKVqyN+bXGaJkZ/uikIwRqAeDJTC3OWLAzkcs4hr
ssJnp7QBtq/cb2t5DziwiBfjPEAGl5cxzMOW7b4zkINAGTDoIwpvVuOCsSyL
TiID+JrpIUlGcp5Dqm8BZ9KGFBQKPoxZoplAkSdE8UA1CvG4cUrIDyFh8j6/
3hL1LXWIourfoFT/kqMlcHYtD4vYCdvWlhTqEVWGyP2zpHlGlEFfDHmJeoVQ
dhIT73tGJxVr2+FUJQTLZlCIDQEL4Ju8fI/NLndsmztKjSTA3cPi9qAcFjvp
aT9/nbQkdHOTKLLiJF7eMIhU130ePKupZylD5zYQAQDrYoE4Cfp7Sy96zyzz
qAmbIOcCrm27V/U3MQ0E+NhOU6Pl3JfQ+uXJSwgLTRVGAr+dbtOugc2m4PlX
b5tDHbL7hGFZgVLkCD5C1FxfKnB6GNHGx18dFhyJpiOBOV/hUa9yWkx6hVUh
/eifNEbGqrmbTP4k5sO3/ar3S7974udLK07PZA+Ye8q6hrEsgm4S+Ot++0GN
rmrpo1Xauka7oaa+zHbPDmI9qBjbUTcPPCS+MM/BTgojtYEKeKtvGI1CkAaw
uidkZAhUuiCbQcx6MZqgz/IU+lAYmxDKmm6dSOdVPIZQCygwJQaHcMrHD8O9
pr6eU5pIE523v4LZ3I8Sb9Q1eZt2IvwnEfSXoXqoUFL3S62TiedpelqrH6+4
ln1RxCV9Bzx7KhgqXFLBaTK6rqUBfxsK+pPareltHLjAf1vfOFaZLrPMFR/K
6CemUyumpyEe/+xrR7VXUzNn9uWjzgI6UHFqI15KxSeRuF+0OZdTV03NlQSa
fvvxwuwOApLdK01H7wlu+XoZCrBtm8hZWM1sHMveBaojZCQ0eRFfFdTI8b85
9ms/hNtg7rTGN/38NpOPLgFiP2ZVjA7mW0XsFGVLL11Pf8+p2SwDvKC+6bMp
5gBjd6lMT/pUQSstFA1al3c87qCfNq/lvsWdIGs1UqL+HpwFz8kzp6cl36Xg
Vcsqfa9FCWNneiNGx2wjwx0Hc9K0khiHheJNW94rlqeiaCNbL/6OgKMzRDOR
ioTXA5bpuwnp+KzCPSesNCl3MJGoEv3aknUCkgAx83CRkq8/pRQG/JWZtMIu
XCR2Ud+09O16d+8s/rYq9n94bMleNKlXYECiatChoBDLTqXxVY81KGS5YYs7
aPuuafsS2wgC45sD6A2TKg0tG0sJ+VItXtzsmhdY8OLi0s0qoMwMDMNIrzYD
dESEOQwn7BGOS80YvyqcPDryCy3ySsUFRmBlehOLvzAABRGVi6NLP3iihUZV
GKHuCcZj60a8Tj2c98EAbhEx6HaWMGQ3l+3smNfVNEB7WoIGsv2g9kJgn/tb
RbXGq6iOxWimQXILGDuo2ofNu4QPPwvQRqlw9N9wkBESjO/MCpjRgtnHy/TI
9WKXnc4yNGCmL4LAsmz3+nTefzaINpJYhIWnzKT67pXlJOUZuFxl8vQEDltl
iU4zFLf1HOx7XN484uTiIo1gStkX2+8O0NbScMMglc4WA1Bqoj3atNmKCC76
h7GEdUm9hV+MMke2xKCX0msoLZZluj+ybT49SjbXVGNFknJvFpoB7qQEVDe9
A6HZ5QKavgO+rH5WY79f2cxmhx+cPn8xwuWHQF3lzXPFpYBH5sSfolBgfg6D
3Ve3vd1GY0UTUXDnlDCJJnRtqcWbhaz3bvVzr+hUV78O8QXCdvScSvV0xCg2
WAgAahsam+ZvsKwN+m6MpuxeEcIz9/6GUm6czcnRbI3qSjkvj5U+OVGNC3yS
mbdy4EN9EXsrbZEjutX6LzO1VyImVNWchInY7vdVlvPRL+bhibU/IzNMkajS
EmTpQcyCyEsiUy0LtQsANL+0aBlha+7RX7Zmhp64Ys8jjfajvfQdbauRzlkN
bsI4JNtwCg4s/koU1kI5prohiKwoRtPk7NxXRXmxrUyBPTrrVL/1lpH7F8xE
GJgaYAJupVwSx6A4t3CzKr9Prw85GeFNwFPhMb+54e8+4k2gyKehy9+RLa6T
5a2oqkPEkut1BqZnrrzXeydFWaKvqaJSeKU6V/7jCPCnrCvJr9PtcEZac32+
2ZWAZ8uXgKMGah5Ohodsm8th8un3PguXqUk9FiopXSSUeiXSDXRlrxu9pJje
FQKx5wlWL+QynWI2RODZvO5/yq+OvP6lK9pO/HGJP2VEFJFv4cWTWU9kUAgz
QBsSMO1qYNs1zVNsUMO5OGDTn0dsEfRPRInz9VvXLeCctE7htvlyaD3v068D
z7jc5RVjmnhmcNsEytdnV65Jx5w3bd90B9ixN8xm8vmBVjL/UG0FqCUb7nA3
3fShmFNVUbaMwnQhBagkeL1i11+Rz4NN6LvVw6hhFN85Vk3QZYrIHsHX9Oko
puMjEndq21n0utF04lHCIP18MbrKNwNBcjf3rsJq4XEfrJbin+icjUFfXM80
J8f6Oew6rklVtR96rl8vQOtG7JnjPSWrW9lu1W8X6rbMzoOG7wD6JNc2fze1
XrfqLmPgN1PT53sVKPg2zfqop5MbYP5e7fVqx/qE0HdQyGkc+O8BXDp93Lp0
UIHFChw+tQkqCesj1lQkK5L+89EgXTU2heONEzV4mcaVMgcYGPmzsaV/xQZF
HlOtcpqgPlbo/mVxCJVRyhpblePo0aXSS8UvkFVG1djjjZaWH8CpjgKYIKXs
o8JHSf6qhTZoA/jTVLU/2YDUZerQQWrF8XzflDIWRJMgBJUwKdK/dSIFOuYO
4uNJPLeJPgNp/Jt36HQNmvQHrqLfNSk90zf49rvYB4d/PHcS4lMx1AGQ3d3u
wbRUlFajRXY5S+YJ2HhU+AIl3Dq7cmJ4ChDqBuhIKHKvNYe5BNNQq2aG5wxx
tQX7ITOGVURuMRquJWF9j391soNhsCZ+E6A5atONy1qQP2skh9samGHyJNqS
CwzGvjCBrVgeGQ/zmP1nxKs+g+lSua2GJsSpkqpJKD4UCaD773CuI2p1+4g9
xlKaICYrIvs9Cmf9uwiLIWTPKyMxQYefb3XdmVB+RqVqJPW2MI9fNbC7p10N
w173ukTnTJQAJ5/NRkz6+M6k2Qo6pTyop4AjQ9P7H+Ev42EYB3uuqyOAKcjx
Jfe6VLkBBdTArQ6sJqVwOs8nUH9GW5rYQHS9OVfm8TcsfDTsCIjZH727tozm
A5CJDQCOp4xTmFhRPkAJNGxpk6XJLRcUaiiRgQaVhX6hv3mkH7Gq0i1B0YMx
h/Gq65Wr2h1m/EcFOsvJVamFNheejo+8uFSSDBOQE9CYSZ1bMSQ5tZpFxbxX
bBgrCC4MXn1UhiDlWfZcWLkyombYyb5lYZCSmh118jYhhj+2EYKa8ibsG7U1
+kHG7xac22eV/tmJsaRkx5bIu3TTkTLQo7YwxjUK/JB5O5iJeOQpU33Cw88t
nab/guBchtBwTNVxntscN37FZ3QZ1/dUIKEdwgvMblddve2WwlRL9Fqni7nh
eAD987E47JC0Up7bo7LvWEhmA+eUcwqeZscHuCD0GSobaGcwFoonllE1gUbh
u9gyIUpgp0KEKqGzphc26KlqI/kFABeGeJd9jVfKLMfSOy0lSL26Iqni/OM3
e9+PpPB3yeoe4/YK0yR16hZrFqAdmHGVdzhAlIaZ8Jc2MukqD0s7zXqSSNVI
FrVZOrGI+O81620sy2/YkzKCFRT6NzUMvwVettF32cQIX6iZirFnNSp6vMn7
H7a0hSC02vhEskh8CAARh/cUg717ntO6TS8IDfQY1LiKuzbBzSpKE4y0jjjQ
pquO0jYbLYBiF5HcDjmaoQCC0uVPlmVLIF31X3UaVh1Z5V9/b9VQagIzDZJm
Gu1HxjzAlgUsL0Kce2kiGFCAs29SV98EWa/fedB3WJGB9wS1ulndX7fRR2uu
h16MBnGAkrDfy5VNQSH6Yffo2luTAj3iVC4E/CohqnjsIEI/EKbAlHE5lrXw
M0pR0fhC2nnrbUR/Fklsait0BX4RztvAcd+kXBWys6gXzoeNKLyILDvDX08t
N3fRLjJ5ogDeIfZET/obUQDjMMwR2qoSHbFFqX9UjbmaGMsKTfXd2c/9Jgyu
sqMPsUe4eBZFnsLo02eVNhyWQNCE+G4ILl3XyKu5lOY1us3SXKZw0vfyPpn6
D8qzJQ/dTlc0Y2GozRNtSItejIrHX0U1gM9KF6NSKJPIR1u5N3ArMjqgCtgo
3+Q1Lu5cyYwSfEj/+i2BRlJizzLsBNUvQRw8ISB2Td23caR01Qe/9hcKCSGe
hf47Bj5fGanC7Dz2dsK8yzESNtv28Boa5qgSdhKy4g2K06hh9K5WK4wMk4RJ
U6+ujJz9OMfdVuV1pCLwAo/HqoYCUINYHwovTBjvnYYvCIX8NqNpe4rqaIMw
a4YpWifsfbgbVOPbCPnHjltriDQiDnEBxSTTriED+oLmMx9kXEo5it/0EISn
XoeZk2reufVqbqmhPeWks2zSs/tHEO1nTBC3lvgLKSvvxrPBuw/O4fC6YSSL
SXzBni7OFPsVwmctZWUsnCXeq/0P+bJv29hNqK60MlFD2Nf7z+AHaszIj+Pu
BrwBO7yQOqJ/lCp1JlNCREuJiZHGTvJ5lWvRX3hX4jrm2xMewGIWVIv8m7Mm
pSWv0r6c77GAe3npFOW8FLBbPj+ePBcHMeOhdEHSpcOdPPlRvDrYQGyVZeH8
hygjakhD3LSmT+y/pJTrTFq0AyzylY4rZ22z0kMm4agBcI8elGMR4E5D2xU7
xK80quUUsDwwV3U6Wm7Iwv1qRdv0RPCWMGGs7PmePEjfdYlLgyTrJsIBP47K
E09bwL1V004DPQ+oqa2G2FAHF4z/OGv4oJY5ua0GhmjFFr6JbHEQqh6dl0Dn
8JegUT5Bn1JVhTG0kGGZQNq/Wbmf7omaqJHtsCnTY+w0l2dI38GJIfk28M1E
+mJTUSBttXzprjW3mah+3dEtSPhCc6C2wZd52UpxXiE8r2ZLvRy/XOWHgtoP
XgHjr1px7I2RY4fy2zoBiEhKcS4JXqKBOA2GK2v2/vVCwod0XGH/Ctx4veVY
E4uQr1VU3W82gwBXtzHhpBzx4EedtYR4pvGgrrXof+sntJLJ5H+46+720ecg
YA/KFrVq+nc6Du5tJJtU+25Bp1Oyg9UpeBq8qNt1HW+NwO6+5DPps5W+TuXp
gBgt/VGzP8x4RSAgttdV7TWSNc5b1PSuvI7FtH6aW/zBBTq9wZf9hvKNLm8Y
gCs39uC2LoDFzVs+O/J0xV/CMpkwrbi3QtM5mpMQkubM88ehFNTa/3ZhfFW8
VLrsLjMf8UoL5MYc197T9OVwZ5zK4VkZapqhA5pqsXw3Xhh48BC4LW4+sB9P
AY9jzABq3hD/MKnQtHPH84hfpqr6D1l+dOc/nBofVzbVfZlYi0rsZ53LoZQp
NWQ1N5GYAj3gx4J3GPijUnBDIpJ+JleM7tYU4DjowI3JM2wAJIzJOuejVNoS
u1jXc0eBQfMsoNFJniXvX7ctp1bRVCLO4Vb203RLQ1ESj9X0NXeNAnbm/N6K
rcyN0M3xw2voB0EhCCtmOGSzSRYaA0XELGhylC3F8b9IjWRftahsCHXaOGi9
hEWbqe3S1JLddLxzyNFXrzOBzmCzVqAg63+RuNB9bdX/Y7ra6nmGeSZhFFXm
FLX3KiZwb3G6jStjcjimxfkrpj9iInYg9kMpi6Xan+DoUNcrqQcKQm/vZsCZ
l99g/WRQqMM9HoekuCirUMykCxCkNDjBZc5CdN7OPr+CnERIBkhYV9gIYREz
M97ctZp+oAy2jUxdReyaeYVLBf7ZHGChkeSMA+Z4xEEUKcWP8ir8d0UJtyYH
VTk61GGsb1C7jxjymC3ItazrlecrTtx1SYXsNtV+ooVs1jqk9wNfYUi1kjeE
Ll5Yn/jHBNbU2Vp65U3T7EoxlE62skdi9DPzIkLRXVjsUtcEPZYx/MlDAf4O
4PlZuwU5uZqa+I7SqjjiNR6di9QUhGd/ZrwtB35zeHWTbcCiHVRv/XOz9SZ7
e9dKZ9Mgntg25B9aYDNrTMUkQM9bDBgUHwopMigkNQoFuJpPv8LA+Sc89DlA
Wn4QRQPaWhiOIKTryf5lc/cV/8ylrWOGgD1XqRTZMCOmvViynUqpWHpTuhbI
CgY4iIwwdRj9+qGc4LiVOQNONgvSDYSKNJRp6iGlDo75GTGMR/PIICDj6lpC
HVcb2pReUiyvvSI6gkVuVXLFur1GSzKvwDKZRoiDjevxsR8eWJJ76yZ8VKEW
JRTV8g51S1NFBU39CZAdfetuOhCUtlpRzZbvdi+w43m27dKH5Kui2O7uJe0J
XWLkXqreKx4QtoazwwaEAFMP4Ls9HeWCx9qCXk65EEsSOBxjpG+xlYUPihWZ
893zCK79u349s+f3v+XZ9zuhOgCEQyRjCFblLo1mj/BeqlpnU4ltyOJKikwC
5Pvev/jV8lo6w/00RWl48lZva581lC1OmxUHPnMC2hGkZfGrw9vKQyrPg6ZK
cNj5G8lsX0R0R+m3vjKUGqyM5+R5GaOGyADz1xGL0XE0y916nw83xkFomIV3
oituea4KR1NOAu260xOzbB1IzcLxn5S3Kh4CWBWl/QcOFUWpM11+V/lpI5CC
rvpyxfN8WzvJXB+H7zccLWfCPDA1Fdu73EhaxxIm91AOPN16K/P6tRrnK7NR
TMpsJEpw7xDZus4Pryfc10qpPt/vUjtoezWIr5ihCVbIU2OjynoBA5amZIHe
xvpybv357eWZQmufNSBNvOsKVNkXKIcGSZ0W/VA/g1hmu0ABYEazu/649DXe
OSUqglwLyFjjlnS8lJx5NYe8M/8RG5PbwKk4Vi7K1jZYMTIBgxLmv07olYOf
gnOdxxEQjqkFf5XwPM8Ancnwsx591pQSshKwiyPBqa/dofWIAMHAg0JEoy/Y
8yFCL3EK4E1TRpu778Q9eo0aqaBl9vbT0aKJaJShYKHfinq6BrFOX4D2VOK8
IQF1+Q2sjt0mDFlEomWqtHZQJlr3C02UblK9rjDEFUommDhryCSAkyu2LFWu
Y2y4D1cqHWi8+d5Ttvo6lY67rSVEEZeTYV7SYBHMHAXFRoDs/D94cvvuscdp
sg/djf/GJsFAc1ecQcBiovovqSC+h2iezeKd8IhhFg7UssDucEnQnB0qsNT0
PIeqITAkSo4opixsjyPPgniK5YOaAdPBYqqkhtfKfKKrGTKpLRQ0eVirlLNV
xOf116JNgWCDprWp0GAvdLV1J0QE/CSwUM7rAkc9TICyv6yoedfgnzLjbl/l
AiQUxqsW8I0bVbAWQYf4HyfTzwq7ml4BOoS7NS7Vp/5NXUAvWamYRRKRaM3T
j2Pg3cu1J8aYNc8jIzTcJ8VsteChrw9/f2pfvdCCmngdhhL1pG7RsP3E/+9A
V/ikQkmB/JC2VtOj1e0MkSfS0eaPB9dEvXpCdONIFpct8LOkwpOI7lYGtxuS
Z/KiU0ozqp9qurHnOqSiIaI1nO7XGNUaqvrGdfd6aQWmyRr4LrCCp6llRyy9
OgSlidGJiHZDY1WNsQyKvcOyy80pvzmbidey7xRYHBQL1uk06Xebi9BbhSwz
8VS7YG3+3McXAHibcY8wIccJy2vz0VwtCOL9U57kZ6Ea3YVSpNkUAp4jl331
+Hy97V3FjipCxuGyTdrMWtaat9C1Immiq2m1AU0PkkdPPFZsLuopiUXm5rP3
yspSn88d9YHXn8xm87bzwqtvfIhi4vc2wW4EGuc26w714KVL/QlTGTX4dJfq
GwS73kY96Ehu58MiTzpPawbYoEwFgsrqXsbZR3FPt+1byKxTPPp6r2hP08si
RmiBqjb8A2WUPfFma/SLhtcNvoA/F2DZBrxWX8Ty4BBvCdju2EsC+ZYehdTB
d5pt1D1+/l6wbBIRYjKu4hii269OKWWmb0NzWHcaBmkX8EjWezEoEIWj62qz
8D09ccOKRb0hSua5oray4gHs5ET/OXnzbNovFwdrTgQVhzS0ZBjl5EUV2H9g
zhL1bJyh2r2Lnvid0X94vvlRAsbyoGSV5Lf9TscBSmiUtMu1wZN2WNKwuvfE
rL/gUKWaIislXXgmp73Q5xEh3ySs12XlYd7CFEXXKSJvrr8bM/RHisMV0Fpy
+f/uWEQ4DKkXjQKGOTKAjggoqRTgtvm/AYucdabdNmS2Jp2lVVNP7DkF0g+n
+fCQZzrp6zun8y6ca4K8j3/GSXnrnE7kU2JKRDrT3WvzP3I3JXyLpn769jLz
MAr2gBdgRz23ivefrZLXHm3Ilsmne7IrOxhyD6OPVVDWvh0fhWB3cDTiNAW0
LzxjXyB/jCfUDawSLAwQQw0+CGShII4Dz9hUyDgRtgTkqh03k5wvAmVMZBUB
YfoJ4ax1UncfVtnSPehqparqr9fsAkTDkEm+E6qfW0BO+TRmtGk1SFwINR0p
UFaQkAEYk24qCe1inBzN8dI3LbjX+pzLS65shV8xEJACvJfB0rY+P68Cng+R
AQQkMahbw6bKqaBYHYSAlHRV/ACSOaBETVP4lQnsA9I0SsUDf47qxb3q0kUD
2AqgZngyuau+tsQTox/n6pvWuJgDK/syW0okYMp0oAbHDxRcFb0r2VGU/9rp
QKXfrvgtqaKOJUHSczVGK3jTe/MnIY97iEfXh6V4MGOuCvbbAHcnXj32ml76
7eAFi93cistaSQw4c2q+qkk5bC+Q4I77Hi8kh8FhXR20IennJIYh74qxDVRI
CbbUaAeN3ssrSMAm3Z+lgYq4IMFByyoYaQftGApUPgsQUq++uJ/h2zLUUho/
nkrYZ3RgMfM9utHDMbfnz2r3Xu3qG3XMY6POrCvT0Vt0j1JhT0t2zzVcDSll
vh3YfpdxGUnZjfjlAo8xr0xHoWOu9bDfMc/991X1egTB+XaPuk31/xReAsD4
/DFDV20rJxbLJIxQlWcOdyG84ibVJQfafkZXTkUU6nxs/7WHtPn3qjYyaOTi
W/53b9gKeFpPYhE9VfdMQtbnmcFP/RtUYcUfHRoG4rZm4yNXTLZ49RdjFCbA
rLVfFvLYSO04Zcj7eyJAzSUs86eTeGkMbyOcSoUckatWjRbx//66wKnMH0t3
pEv0T4ovRD1aNC0ImRvZDjNkyKSsloOTKeI4F3kmZdA4RV1xBTl+MWJ86MeS
7O/vY8h0SUfAwhZS8Pn7SXZW4hI5qOTLQtam3tTJGFz3fVE8ESycz+JiA3XX
HCPoyPeOo2UqaAhAnc2Hffg+fW66BorfHVqf1NwG1kJ0+j2s1nVx8A3zYin6
BxEL4m5HrKk4ArPxa7TZ1am+DZHYT5HEbcN486c/Xt4iik/0r2NAOoUAPbnL
zJpJeP+maAuIA9fQMKyjLWx03KcwRTE75KgCYVhAHVAVH0B4JIHv1LBPfNwz
UcDpuhx2SJRfM9+FHAN5ZubF4WvM2dNwPc86GQbksxCCpNk/ImfPnzDbvVBU
CmAJN15h6V0khvo+1ib6sh0/RqKFTMzWU6Mi23gKFVwt4+s+srmEc/YlA4GF
foGEcQ/oQWF7tXcOV9bhFkT8MzNlxE8lIGW9Grv/svFHHCq33BNQuafafv0Q
sXl10Kv2z19lEbCnHYNvc3fuAfSPPFmCmC9RL0OT941mU5P4cEvk/HZFsK/N
Hnz8onbbum9pEXK3S7ZFdsEBL+1rGTwnlO0zvjXaqQ58J7fU18MhscosHUt5
6PrToxdn3LsqvQhAerPr9rcPBVY1Ms6jIWs5dFNfGwq5S4cyRoRVsmyoDbXU
qtt4E+MQ2jjcm/OwwOkBXGOPBtCV8FacAlACOpWBAlKsNjevBUjUx8vZQB2K
wvZ4wQ6zY1sulb0NmbJBdqtInf1dtHAW9UTnjFW3rjcbAP8pB65PjItZ3T+K
lwOVrrdrM97ff+Ky0C1nqlYQepYtuQvF3OAMTBw2W0eAVRO+jNeD6F9geW+K
EtRuPCaZ3Y9Zmjeom4/eJVIlYwmKJapT7Yx4QPxBHwExiU5T3ICoAAKhz5Y/
Tv+NmW18Kcct04VtpSWo3KZk4V8hrL7Et6nEMvvGvBz7OBPLNBROi/U51JZK
2CT1mPMnIiT0OquRpDc19Pnvi5IE+gw6w1vbzQtLdoBn/zx+om23ZCaRHi8C
RpfxYCdjaqo1vFT350HD1gQOHRhv1wjUF+4o1ho4mlDlWdSDc9mQFnQbgnAT
2VZ6AqcXOOkmuEVhbPb9K9DggqzfWBtwj0eSPByetsGi+ZaHfIvpUc/FJBXw
8+HuuUuIDUCPQne25CmeYRisr7o7pksN4Dk8VVdA5I7myztR6WQa1Jb7k+6y
jcapLSZgA6zJay+aQqyKPhQW1edRdKEWzhWLuXk9zj3S/fDTdtwE1tb0314/
p1IyPbXs5aCO3scIdMpaLw/uzfwoGxY7BJethbdznkL/EeBVfgl6IkK15dF/
F4wsZOm8ckMzWWty5LWhfztn2RZ1iX4zijgJUkuQKjEb6N9fmO/8newP2bzD
uyhHUnEVYmq7Ve+X8br0cWinCtY0pX5PAHr4kLz7UY0Hz70Pj4l9Y1Pc+Aas
vGF3lOI00bjduAPc11cYaOdXeMJ3nZyn7vEf3WMVCX8UFqf2803jAFxpF5F9
qrE6lyP3ZIN/Ta5yPwsOp6BOqZbND553d2BH8DeTL1RhFEosQyoK505EfCut
YFPL0my8kWmyuc5dJHx+4oiE6Pgb+gx7NTipfvC/a7IaXCJvXSa47oY95CC6
QffB5pc3e3J71FyggH3YVtmofqIJoCBm0e4QVDV/F6HyOggqNnrtRT9GyHmG
GKsTT4kPNut/l3yalkezbNwr0tTBzIqiSPSOb3Lj76Ibl8+sruj3IcpNwtWy
IVDZ3YalpmckL6j5k0eLpIqwGqkb3dBJOan96Bsa6H1jK0MapZVVr8UJUz+L
3By9h+BLy4igDshz2QFJ+vroSBBUQjMUWXcpOdch4jDPO2qAgqyw8sOFF4Vf
jbBinJ798C8/oDA74O3cezQxJhuHGFyoKvndv4RvaZa13WVIkyICEbDfjZMZ
Zn96wsFgyd3IinRgPE9jBU09ujhyl/yG7LbaEiAm9gBXo511SBCTlutlL8Rq
l8TucS7nunCKq+wj2J70wSqWZiDtB7gPmZhWh+BrAX2+L2hNyMnIYgrGJH/v
hQx6ECirgT1oGz149+GQnj1pVbb81Yxk5137m2QYgl1lUeHZinmnMG21TA8t
GH5WtykfKeLU9k1npSV1WelXxTPRVeS/RldsJfqpqrGJi6p9aT3jBfKpU1Ti
EGml3ib7t31Lw2LwwRYDhX6ZUDjEx3U/DWkSSxfBq2kS8hazFT4yISN//3t8
GBpiVzHTp1F9xFNbclloaLwnr8/p6LDLF4wFbbZI2Mq5UG7Xea3LxJGx5J9B
wiGose3KjolVpDIcRahsWP80lumn2REfk9CNz/R4bOZqtnGfwx5NtZ6EKeNZ
J4hiN+xcFKZXX2UoAFG+0eTrOs7bkKjfX1/we2JNUKBV0OEC1QQNZbwHfb8N
B12pKJURnHMkhTpFZYy9gPiLUePs07Wws4LoN700NDtliaNGaB3lQDbFBl2B
Cpx1XRVVIWFAveZXYL69fPDK8LuBZKDcUVQtU2v9ZiMNdgctGdh+7Qo25rq2
TQ1nuudH7cacfVwHk1UO7UJymmFqk+O1eO/HnNOLIAB8MoX47qSLtUPXd8Yd
XkNSKHolPZSV3jYY0l/21lfJIsYi48UOg9n4f2y2E4ffy6pLPLAA9UPA4FZ1
mn3favgGN5nzyWrkgARX43lv1hOkvgd/tFZNe1CRD1Q+VUSKT+WM+hTa/8+l
An1dHce2cuMcmyhQSjwtjBrFWd+zgEF5GsWCMY0fCpic39NyQsn6KDSxdsVs
D6LVpamw+UlKcaNCgBZD2//ipf7bkMywHhZsjBjkyt0JNVh06X+7YLieFlo1
Exh5lNTrXKGDyaO7+0aJPVfoYv2K+C1Lvmp2/IBYYVQvChJMmxi5Re6csps7
SO08ZGhnabVh8FtALutyGXb/YdhniOTolN8NGAYwtxpoYdJQAbAAWFEJ8tE1
Bq8NnE699Bg5Toe9HEK5QKgMyGmXai2Jz8ocn+zf8vZm7RXNQKNGs0mM8yza
iKhJ+WMcHNc1MTI/FT7JpbNjGQU+ACGNlmV6wD8H1i9O/oiToMLj4X37gXls
sXdMXn20nVb1hdcDjhmzFGmmCdtTO0houm5kPF/PxrFZKfjUPfYmAB6gCsV5
zfneg6Qt9azbutDOModYfTFHiGrobQ4YN+RtTRAGgKV0cq0l6uY6rWtEcGAe
6tvWSoFpUdhwqIXNZEMexT8fBmTpqpT7utvTfM63npiG0NaBmsxWZ1aQMFee
o6KmMnPzLB4GHW+7sGBknkm0dJHl02oYWKw2o6ZRNAV4ki5jzB5EyMGO/R1a
qTvVy8Ns5jqmZVAyc4PJJHkzwRLgDf8K+bsCTxwhUuTeQWod9r3AA2E/5PYz
hoFaSRvowE/V9SUwRP3msUZpMU5K8WijmMDG0qFXE11igTDhr42hbaxgAHa2
vEbbHmmiAVWD2czTo098Vp+RbNFvcPbNM6yybtU7Yz/t9onhz6TUW574GtWI
5nNdxIrA2bS3wvFle2klrmgkYIaRakn0kJqwT6Jx35kUrQTKrvUcOFjuXC2w
Nz88y+vzh7MmTkj8eiBP8kvnrQ03PtuB2cRM2S+JHQ6i8KQcev5TuL88rPP8
INTZxYpn82OUjThYNhYB9YZrJfUwO6/XcLwJK+/7eduQqCxNdU+9hOvpm0CK
cOQMNCHsMXEbJIg9hjVPj+y0lsu8wWYrs5AzUigF76UFSbpW/VCA7MAOmIWH
mtL5UE/nUz3Hp0A4FAXahRvfzHW023aLWgayTRKEay3Z39rNC2+CNcJVL/Rh
TueY6pUwEIwyj3uzYVYaFZn4RxFRMp9Imr+1IvzNW0/wa9jm6lU6eUrJmKEK
aNwjBpOlapGRfBub925t2V1owQ1AQybHY1X4zr7bZY3wsEH836sy50iPXO5S
HwoQJ1voPjDtMKZfrAaiXda6RcZZOnLOFqFseM/BUTVUKrYjJnNHkeI52uS0
Y60goNTC98m97aSRKje/JILPbiY0mNiN1PZkQzyvzFPwJTvpW7w+trZBsUPw
0hEp/v08Z+rHjnUEbvI6q+xcapWSk8cijgYrrTTd3AixotuEmnwQvtYgciZm
RpNcyzlq04R3fgb9GEQYhAVfh6YljVSVb9GPD+GmbfDiXPqlJ2hiDheKzQIF
V66bsANlvzOgFk7RdZaTZkIKSmaHSyHztXJiecQNofN0gq1EJREpiZY8woX9
uFur/H2UtIYA0p3z/kv4BL3tdY58+U7SFZ7A8/1MR/EhG27jwSariZNdA7SD
QOk4yoq+FM5o2ZOKnuvkVMXkHzVm75NrNhyhyVR8OaQPcgKphBcoZ3lRZc2V
qTWQpUL9Z2uJz4am71LVcf/1xYSWq+ZxgusZcZ7/Jzoe4TdxuDbjsEJZmc3+
8au3Js9G8q/YqEhqcyoKkUvk8GYqJL4ySZZf2Raf6A0wIfMywZJyueAqo7EP
6eSP2YmkGN0XZHUP44JO2coMAngMG9V/9pAGfqA30Q1LratAwV+n9EPRr2lC
tG/SIt+WY/SkUlVuWDpuYt1S+KraaME4oV3efhNhcRxcfoAlrWBg2UusryoQ
TY3e+208x2PksBvy5xGETN66ejIHjCybCHEFTtQwHkM9LlRWEOfqNx0ydyFb
OTaen+7RK6npb7W6QUmbK9Pu2NsJk33J3ajG6SJVkeDuEfdrZkQLXImz0hEK
KNw/UEEAu9V51juOCzfQqqY3/BPEbmKhJNOY6/QYRejaM2pN7mWoSo4VvM4i
Igl7jZcg5N8JBDUBVdHT32uPt7AR1ryV8iKDu5dzGyIFTkQ+aUp471rvjHSU
X3RFbr/ln4/fuI/0fGwYPPcPkXo/S+VdWit47EFy0TYuNbFDBEqdpdi6pe8B
pHNNIqs4UeKlKPy45pih+YiJWJaE1A1eJS5EtsBR2cuJ5+Q+aoWZDaottp+r
hUymPhHEwoX2FMeziUs6aGBe9PVXv52xAMHup3QtDLjUJylmJHQA8qs60cqK
5dHNIrVD3679r18/mCRwipU9Gl5CnvNULId9AfAJjRqlPxasaXyZPuKJb+E1
Tw6S4RgcFnr8xGqtIa1rTK6zPiC8l6Y4GbhlMGI+SO2unDkvyIQcenFZ2heP
z0CI6tTB686gvMo8BMmcaVqzWQiylqMbRI6FuPiWo9nTAcDZSSCpfdc65e97
TtTqZQWc9RCfdDLvqXe+In3Lr2+Xugumt1j0ixczidncrp4JJojC7rON3WiM
mGUKtZ/Tez64w6JQ20mAIUZieCNzNZRD5s/sjKxWu7e6LDgZWCOKoo7KBQpZ
yHtsgBvEqKzJB3KsjZv8S8DEqPrzdzDd3Nmrdx+ONEBGNQl6xyBRHmR8UKGl
iqCIXX6CaiANOHX4N9Oq+TJ9lwKh2cWQTYWBKWCvK3ViZjPd5gnRx+OTwe0P
nYHDh9PXkcZS9TXXRF3XXDBVdkq0xCGM56Mwaxa8UJdNlUaQQpKP16Km0TJZ
GPqyaGN6NCISK6lznpNlzgZyXvdUMGsxDxl0mOC7+cglJk/rseCwbK73HqXm
mms6pLTcEcfDRbeeFA1zuQtgnhOcwo2ZzElVzgH0/5iS+5MeR4Jzo66+Mhmi
cFmA7Y6Ivue0ZmwlGzIWW5YIgFaY7zfOreG9eODbBfvmkEd3OGYe1jxXAycU
EkDHUiuTfWl7gkrWh02hm2ei4ENXxDiE+Z8O0Vhq2euGpo80zSqYKu9xThDm
1xL8q0mTFVGIhQZzZ6RYgirK/XKuCwXAllFQEUwQ5fGZ5eBKtmhCbBXr3IHC
zOGIZJGUooYN6Gaa9KaWKkModVuQP6XD0z3qOuqoBrV+JvMYT4w6LwUVtrSP
F43PhUa1mIhMPNFZVntAaHuu9lfT5kgaljzWZiM2V04yOPpX3AE2YQar6Z9g
glnZBsjrlKatiZZAkTYSW2lA27MrcIzkP5wGn6x5TCctWk8EnxoynjF72kXl
/DEjAsYpZFKCkjd1RLdOvr0nfgQSut87MOeE6CvxAw6AjL8CUoSq7++REd67
MHpggeToCu2UCvCMOCEs9msIf1XJY5Z11dXpEt45RuRKJYixv3Ewk9YM+UQK
T5eJk/IMagxZQ0mv145sc0DAExzS6yyP2FmQx6G9AmYP+4wFPi6rva3Nw/hd
DQqTPAH/cFTRPUq+0713RvhXUQkDFHkoNocPe+he3D4zT6oinBhDMksOGXhf
Tm8Y8FN2BuZWrnbAS8MxrSPNQZ5L7ivkdBY8ZkzuLscqRE2ICWtjDu0Y4Z+s
TVe7Oba7Ily0DvdNT7sjSyBq5j6PzrXthipQJ2xP8ooXGwJ/y5Nq+t58htlH
wGRRBuOVPMyV0h2BTIoT9lMfIALjZj5adKMPDTHtq/YGXT1RrH9PXxDD3Jw/
vjnKjaGr1/GdMW2wHG1WnvVccKREhn+IFkCfsirO8BqVe8K5Iqou31WJb4Vd
DnUoczk1G/PCOPb2VjYkiBxRwhYSc0XYIxGD5KlYCixQdlBuP5c3XDkxCsio
GVhkrxpKMgPCvf4RJk6llvzqYL00NVBzCOTyoJuLmVtG3WpaKXrGZVgf9soq
wCL9gsvr3yC9HxPa2UeDLkqvIXCfL+c3yOERXsYwvDGqDjV4D9Z0wgFBWx5M
syhY4NYU8Yn+T80CToGsyoozIgg1Frr50tmha4bPEV2GnYJjSbwk+2r/MWPu
kKPXisfiIlvFYTwqK+0VuAArzhp2yOUXG6Zu72GxS7qX9NGd81Ce5AgYwOPd
hbNxQJyT1TodwDMxisiaTJKjuYFJO6+MbE55ZlQZfpViK7D3wAiOr8VeQ832
Ns6eouXdjv1iuSg2hfDv8p6BLrvVHZR0aXlASZE2hVFoxjVBbl8HhNa2Uc3K
cqA1RHy/nr7lN7D4VcsPkpuipfp5Qb+NPWk9C+nOry1Hw/WE74Gf+5p24ltD
JhA5j2vEqeg4tQ67BfGQfzG2yXnVJGU32zt+sVrXsZfXpLmh7LLn6Dn8x28z
eCF3pM5D5N1OTSicNHX8LQgR1Whw6x/j3eKXyksC+521Gcs8N+FLNBFgrRbw
LWnB+WZW1t2+u0xGXrP3ZUyVY1UFq5OGxHA0H5KWWOS504zPUaMMByJkSfME
t7XFJ3zgn/yk0h9+KYyo4D736nTdSVCDALEaimz4c6/TYX4J9UER+cyrxFio
YCDixR9xQth1wqTn/BJS1XQoSewi8XjrPF22eWt+EPi4vXG0brXREG0jSfWY
ovkUnk564wFKDxkUc9Az2AQNW6WnnUG/oiitdX1UDtXx49PVTQUl5Wb+JFct
0dzDgCuMMzZ8gapbQlObu6fuFogsxSMKLA/od+S2m6a1zmmVROm0LwhNbV3W
5QRDR34Vzd+nANST+2VBU0Z1ReiDKJDgyS66WcrI1+Od/E+TRXqpkwjH7kbE
7fXYv/obODzbfVzwXM05aZr/wZkeJjurfbaG1Bsu44xQ8pit0QnVZCyIbzla
Hssq5+v4c+VG0B9Haq1HH9NSBUyNxDl0cqbcuNizbw4AjjpO8t19UsaBqvf+
+WkcQQxdkj/U+WBXM6c5zeVFR4p6AhTbB9LgET3xIilo64+W9xp99ygD5bhf
ZhMesLvvB1FpWwsbNVLpIZ8z+gHik/6E4yJgXk6zA6Q6+VLopI6zN5xBbBuP
d/9bDV4jLOZ/wdKt2g03eXNiDfteiWYQrWNBBZBRu3CeCDtwpB1lo1U6k252
aHNjkY2INEjwLlR0jc674RQ6rE2UHu3QDwLJnMCwSviI9slvbBYwIvG4AaqV
+LKStbeb5NF/+FNYbXQjbpBQxyrTc2P2izKbsVe0dx+XiEKldP7wO4OqBZ1G
k1tcN0yTrf0Cj+rhQMKlMDh7q2f+e2QkCL4QifLNLhlKKbgRfP3q8LSxx2gk
z6DhKe2D48C62aAA6KsTD5MvqTkbung+2o2uNSmDvpuG1Lyf6CZgx6bX4Mz3
Jt6FtevVKrNO7Q39BVcbrX3rvcaUwQCInoShi8FFOPGrRyaqBOsZ8JMPFPWM
EGjch9fAWLX95jMl6a6pDXBWynA9DMJkD6O9U5lo2d6IKfGSzImRApEfLTqS
/2OrgyVXO8cfsDL1v7OXPW/aBGYv6H3kJVpiZD/xN6LqMR0reRc6avJnwN6l
vougI/hRGY/HIE0SHKvtXhNmnmU890dpWtfB4dm1R5qGML02mr4Sxcj20nll
jju3AKMGotK8b3rEpoxlKTLdy11iwIz9M0lhKQtsbskPwr4KSD2Q4m1Z5109
XAH9wk1Tc9dyp7UPygOtFshZTj/EQvANJBDXPVRoeKljdMXR1VHxhR5m51Hy
EHmJqmAgAu3GL1elhLlx+/WIeilqtS8uooXepCFwWlwsvUXCf5aNapDni8KK
1XkL1KSGVwxm5ctZb+a843e2t4hrTEZR0SMpgWw38X4WGuXXsJLEUjt33hYy
hLMu0VODp8awnYnwFCaJ5EnLP5lj/CnK1ZbXD0xkx/WG9BTpliBJSt6debHM
iE9VKrK666ms9/4nCLNPCBTvIwsJi5WuftDDaTH1bBrhMm/oowMoML2AEgdi
FTkh/6gXgf6YboHmv4oz3bb2nXyLgL0PNW3QHCMVC8XYwfAVPnjIs4fws5dl
Tk8lyXab1yUyyyRpwFoQs6ZVLnA9xS6nHxMOUmxcbQsRLceHmYztPwfQa3YB
tiuSjUCnivURmJoN+nU1uB6jdCXqmREnlzbSuWyo1V6xczFn1LL2GBHYDikl
MSQf69r9V9Wo3o8ZZ1vQwiTHZdCCIvGFog5ptNQsVskBxECrw4Fcwpl+IGwO
TfmVFzcLGRPL89iX+ic32Gt0OZUQBo92jRd2VIH8E74onF0JEfltBEJY0djE
loUN29krmrXt9Hh98MMKz0TloV5vIrkT6R6YTK6/RBofWL01g5W2KRjY0ug8
EGQWJRGiA6ZqP+Dhdrq3S/4X+oGJVvzUdi8VKrQKwDBFHODfdKzgdoztAplV
EkBybvSO1Wb8FdrRXExjSJNr2DN93j8BBQH+lIijHq+LClacg5pcqy/HtUc1
7r3CzUTcpUlnHSeug8auxdYq98zJglpWCAxRi6UB/0p70yZd1SHyv98/BaZ6
bLpkSl7OFQT6piE/gv4dP2AKWv4CMeW4AUZinsxh48fmf4nsGBjbfqRdI0fQ
xMzZ9k1KdsBKqonrKQOuv/WMRt0rZDHZ+GQ3eh4wXsJNEsdPYeOUrmhyRVaV
qcoCsCT/2hIudMdnXyM9bulUp+Btm3CTHhWEm3Ji6PetU5+Q7OyPf36sKeaS
75zvTvuyvzFDiMCy2sF7+MXQDmaHLDaHrM7RSa5KGM9nPZNA/sDDZj+/8w3y
U512jR3RpY5uDrOczXRxC+SiMt4PnvimL+W+iRMY8DFzxftpnZ37k8FCHBBe
4g7Pi0Bfm9NNqlyZnZr/066GLN3BO2Ic48UQDl4Ctaj7tCB7eauITjCkilrl
pZ8/jPrbdseny/1Bga94EeiH11BOqF10L1Y0y90lhglcoV4TMpl5uLppUOe2
uJJj5rP0mlUXTCM5UGumGYdFIO/WdbhfF0C9Ykzik6syUe49ZnxWBeXNyf6W
X3CCGlbwM/W0FNMzN72OdImOUDXRv4oEfdKyRvMtza8Bv5+Bysll2P1yfSgB
rWsXkWRenJvzrxw1xTLKZiafoDKtJwT3oZltClKZ+Cer3em2M7cjUC8OplRD
OllfSBd6digflGmfJyjtemdkiezuOOfLiCrHm5PXK1Twbt+Ui+L+AexES4rV
iabZvwicw+MW89/Ohnj29GKBAkepYlgmCJ77KKoQRf/3m0TEfyKeCPs9ut/C
5BEGKUBk1Uwuu+epkTtPHWmG+AFRRjPFhO84i64xFU+2SJMo9es9xjzWzReV
KzCqatkGEZyEbz6YrL/+aGIpUtlcxXTgFa9BRDy7HHI+GPTnphFwU88K6IFL
BH68RWEr3MK7PoC3opHhRA2LC8MhWs442MZeV/60vlEXO2vjOPyZxydSsZWL
+f/wDqdfgswSAYwhswDwnUCJafkJM7vXFVEZHGVKXyPj1vJf/qaxyPT8OaOl
YKoJN995+fF1bzBfh+WSAwv6XmyeFGNut39sWljQh2VDcHuxAypataz7Ge1O
FfGx2GBdn98tZJNy8T6mPQgd0bilQXSD1eIWJuNGWtBmVgDJIwb+UYCUfa+8
q2ZZko2nNn78MyREzNUeudAZWL6cVQP6Mp6UNU/Io0tL1UypkdU1ZR5IAsAz
Mz4tIZDJGb6XupeK6znh99Zxh3l9YjFmCXYjFJfviAkjEi1mC6tcdyYh+xNh
Dvh6XOtuX9GC7JdZe7ckBdg4n1gUR6SsmDZ7l/YLQjp5UAHbarCiSZlBPENO
tUhaMitfShRfiNEh/om49+hT9MQEHP1ABIjWBiWBKPdbChLNXb8lr3I7Fad+
MskVmFCdxiGB63F6/M8mmEYZPSFEcyUT9EQu6CQTBjQyXXCQ/e1SHDlZiQ6i
T5EEeg8PtNJUywOm/xwWtTfrzoLSNiYW0rTAciIUkusgDTy/Js6XUIrSppWz
686t6d5TsGKSuhU7eF9hL3aUkkp7FGoUsBi7I5fjdxzhX71ZpGCE+80sUvW9
4h3qNBdUR3+cY46sJCJJuaMITZeKM0Od3Y/BpPdepThLccxUFbJqIpPsWJHO
OwFncX+lPdT6/QBc0qwfzwbenpgle7dT38tpjGJyLF8RJMVRFsNSX9wOJ7ja
pzX6Xd0L1aGQQ2H9kNCKn1YJQ4J2D2gtZgLxY/4hd9PJgulFU+UOa2t7VpWd
AD/T5edMUZeDcYh6V1LCjLsTRofpV2S7L2cazsLYfFaLjcI+n+beEwtS+q1D
FCweqinr/6JhCgr/lVCWCvCQV1cm8RitlL/W2d4DCFPgutJC0Sqdv74G68KC
4ka5Gojx4wcP1tDbsMFCeRRX/LsNkWdNmlpzbbgnXK8bqs9NVhNGS9EnMoEZ
Gi9tHPwtDfYFPwUr6+EEPLogTE3l0LgpcaDIbQg7DxXno1xxAvmgV3R+Kzs2
B/rRaXnelsC7Mq1T2a8036l7UTOLXH1EaWpAbVoKkzHipZejvtLfXQxkfiyY
uHpgiuCO6em8deDl2bXx91z3bntzdagpEi1izkNmTUpt3EM0Z/gb50400P5T
BwyBG8Vp4PpWjxnPfl6s1djh75dTgIIpkJ9HOz9oSSiXHF83I9ezKy+qdN0h
c2dDJwze4hGOdFAZruugKnoS+Ofuf0mY5RM3we1Swkabz6saDE99FKHrx3ea
e4pWxbzxUJBWDlY6kR30Dvw1RbFokX//9JLFebmoWuoMg3J44Rc0uMs/U64t
BA7SkAqWXWKKJH1X3SCcNjVQIAFpxxLeZig2K46iIMAnScOuo9XpY19+LKVg
qR6Q+F48WN6wtv93pX1FAga4YSAu2iIyhO1tfhJuBZeu1hP9N1d9ayvF7nb5
qCcAnOFOmEZn3XfHyNWOVwzgut83AO8H1aO9mJ9CUt7TNAELZgyX80sMcHL+
uCFmnL0pYwX0BMtklm3vyfTRXI25jJdRa56s7XCU2Vor7TyRVjZJgEbBeM9D
FDkGYZ8zSe5vBlyvEh5JgcJdN969UK1d3HAshWXd4Qw3miELZuDip9dkaMJP
aobRx0lRpKxblRAyDANBdYsUXaI6EpAnKpt4OTTRreHscQNKa7gxzR82nmIO
vgPrhqvFrdwyToJVbaCnADN8T2kUPCcZfyuLgIk0R9NSWuKL/MvT310ih3hA
shzKu2DyfC7aVd9IQ0oz5CeqbdUemegiNd/Eklu/IJebp+mk52+6enoUylzb
10UbnmBLK27yJQeLXKh/7IxGr3wigK1N721i1SJu3fQHs4vmuMsx0t52Llsc
2RntqQ18hs6SHJOF0ahD6JE1sQHcT45MzVtDyKXcuq/+CyBrZRvt0uuHrZjI
HhpNv+sTQV6rfzwxg+9z31sIRa9Jpl6baWOGMEaFYVOkR1FjxJAZY9DXg+MZ
8VzXARa+gmIVwV2XrcTxIX7WnS2DN7/Vf8VUmLNsJi83yocuNmYyEpt9dh5i
9/wlnGyQewnfMhfYQMpMn2xZSRA7VsWDbwor5e0qTrKf1o0YXULSp7vvdxwW
BdgE/C1hgwvAX/fy9tLZrEmwFNWsd6W/+Hs0u88br0KLiHd/fKM9Z7QbShgt
6JKMApxECWyY/RdGvnoNNh9yShJzhqhD9n5KKws2am2os7vIiO22+F/Mojvo
nhTkko3pK/DBlQPibUiAxfU2xRYLdXTGzGuzMTHHdBWDPOpwv+Mu5nDMF5ow
LxS9phFmreUptgH6xP5E4SEqjzZl4sRNrjInYmXNxzho9BHArOuZFTJLZMYV
b3puvPIHkAgJ8QyquuCX+LAoN3ZExxE98MQr5nBKnGK2zaeB/NaqXwUAAVbd
dZNBKRRsvRLigt14owW34mIJ+ODe7D9/gxMqwIkFNw6U9MgFFonFlOAoWf9F
mnDXTs0x8w6m9M0ihxkOPCHW5HwxxH/8zw1aP7y2ZQZdk7Czo/LtcvFMEZnB
yXjqDTQfbosPGWFYIYP5fZMx9BEWOqyBGftz8jjsm9MItvaunSOYuLDDvQ8T
RDENVvYShmEYvV9J3Rwq3mUP8m/7+dXi/3HFwmJzx2SitMyIw8hYlLCjeK+k
HpkQrlAj6CTMuEgcdnZS4OeZAIBtfMH4+LI41c7iTyQgpXqWTgKGWXBKprpJ
jZ04gN1FdZ+oc4wt3ndTdscahCRKhVzw6rdBXyuU5ARiBqq7HReNj5L0f4dv
wYysHIrT9NnWdLCtbKrDkqou8y8114Lq3lo3Y/0fyR9aXJevBRfD1UWkvBiL
jMmKuCuJnHn1oSMIB67VtdVRmO5/alG0XA9ThFaE3qOnv0DWVKzuWBbj8UiO
fr5SSxEhQrA/Cc0ZkYHfjSH7OT2uOxZf7Qh71vwNnVjtqlLH6sVdVrAH54nR
NUNoj0hnFbz+JD86eoso1Zu49EJuU7uRXik98SMt4Nf3F6mj4Qx8zHlYpxzI
M5BhOzBgTQ5xxa5byW7NfIh/olVE2i5oy+q3ugN3zD20n7cgzFnK219RHXT8
SFr2IbuuQAOkulDPcgdfjaBO/MGX3QqPUP2wXu/GGeqQTTRPudJTTN7DVOUD
7dGjnEnVjZUE9ShNjtdCdrum5PAe2Cg26wsw9Lu56TfybtxoP4IDG1GhjWyv
mHEhEyLkVdSbYMGdyqKeaILm9nDfRAINJbun/mEXmf9VX3t9je22aJWy3Vwn
mJfa2WoPpZN6JrhfGWAnE5Zi9y5MTUE+q9y3IWeUgfYVhf5hY74PVhNui6cu
QoekosipITs90Vb+YihQkCDXOHhUDX/HydVO+3rDjZ4BZzH4sDm2Hk/BAP1l
DpL5xTiFQQC/4xIRSLzQM0e4QwdEBdJabm6E+alQXI6LlNOAZRHgln1Ly3A+
OtYfYjhe1v9foNa22w0KkAX9q8MDqJndkO2nBj+I9LlNrpBOTznwXGQPEe1j
zNRZ/vYQb+WEgIFMMNq0m5N25rP1EpB/B1EvD3+rCKII/i6CsaeNTwGXxg/f
Fb6q2X357/M8Lw9Gt30ocYDFnyf6OD+2UWY8H0FMUD6cDxBuL+sf4WL3zT0u
ITFAS2m4w50JqXYdDmPqG7TJiDRhEEoqv9igKsN7FvDh305jLbRoSZftlit8
f2m1fOHpO6eHJwfiixIGzqo9kKKd6tVT7vVAYGuOnu2QkWRVEPTXOtNC4agG
YOoAkfIMs7zZ+EtbE0xOtoHV7OAW6Ubbx3fCQkrDy4hWdl+6K91z+0GSZppv
sPkpRLZDgiBzemsq109lxEMtuMsnOD5jkuxcqtvXoQ0jkvJNmbzdByqeAsSx
n5ZU1X1YxO1dgqgZ7qoigVtPu6IHY3pu9V7+/St5ACBMeRBut8zM0IAA+3nJ
jGysMTaM0eJAoLMK6kLInKRhOhmTDEYIeCiq4HsGW7d+U6NWHb8md4nvHYjq
S5TYyXv3hZ6HwCm3H6bXnodU4N/OROxCZ6iqW6BZxaIF6VM11Uyph2gjQbsh
9Fnw7sIDVxfYgHe5sAsJMhV0RjI212dPrOW6kgT8Jv7Y3WePpxD7Z2P+/vLH
iHpSltiHP6jkVPrqHYNnS7S6y3UQg9NCaNexmuw0nIaN9tKbJZXKR8eEN6pi
tFUur9/8lMQhPRz4T8mwVdP1wzLqgzVcRNiUKpSRn3j5wvaqGtW/90+h3Ubn
T9bDp+foko0wIjnY/uwJVBEez+rXol/Bw1v4Mo3Gzr4VeZmtIuofrhpvTsSb
QHyMy8E3JdICd8p/pKm3H5u7bvzFKrd6oZNHS/mwiOqOffOokHu/S2JA4Hs2
yMSoQOBJ+2v6hqdaEMrCAQqWwdVX2WhAVLN3SwtPWUjD8kTe/pQ7gK3ZEfA8
8KKyJGlaUUnVF0Af9iSSjUB681q9H6KzmERnYuOBIRenq8ahhhPxROjCC2X6
c4ec+IcRiLkvB2E9g8e+TPDGMwyQZZxLQxsrob6aOlzq5hwZA66pSMqyIuxF
7ShKtgZ7ibaPZJcrwCSvrNdCZOAMnBgaKw9KNimVkDX/Ip1sLydwM6fOAdrx
AT/ZxmNh5M+FzTO6r0Va2hcuAr6MN3zSDD2dI+OwmtqP8fl48bYSHpANsgMd
xcoCuxDXHeLaBA6oxel8LcHHwvYvs9/PQ8LRz/1mGGBbxQ1IcQS83bh+oNpO
RP3lFcS0Zalnj4DfCUKVkXcn+PHcVrwBHGLwlEP9ATxB28d6snPLwqqXgtdz
hJT7R4k8MrF6Obx3wYMF9FYynuYX6fCRdwEussSTW5KRBya+KDV13nfPzU95
3fuhENMxxB4xvHlnkKXSB7FuThHyJI6B+kjXVgE8N9IviSb4e+w3Vs29hiC/
psa+5TUJ9QsME6lSN2jaljuj/+tu5AV6AIlIEkfK0nyQG1jGJOUZAFeDYjev
hNKYMukpc+ErxHiPqOAaS0kLAyIqeaHdVsZyCxmwzgLPPUs6ZP1PSk/ExjZh
8JdHx69HXFvRb68vsMVQvcf1Rm2UveyoR4UOMATe4pC51Ly+sMhRoUw+3BRR
xK+xKHB0K7yX8uGFml2Acz3Nt78xeLjexP62nutx/yCysl63d7pNGsV4ppWG
b/B1p4/l+uB9dkiwlUGDlelNa01lfwnSIVEmpvIgZVt5rzNXv1CMaVeV3Mvh
gWjMSo9F+M3J0zaZbrLHQX+Bca8H+ljmRmMXoRfDS17DpZoFVF7AKk1L8rLr
MWXtktZe5P40jIgKcyBp75XkEzTk4CfWjrpopezPARqtdYrCFxeiR33ujDAV
tJm0IJTFqQVFUaZt3rfJm/3zfvMlphgbh2N2qtmkGNpWQBCHs2vbultdvzDP
+qOaNeTW+sCnG6QRjtgy1wLLgGka5owH9bPZYDUXHPeD+hsTQg5H/0DZ5bWO
PRCRCpSDwYdE34sbtn4z61vqHRMbOgep/lfw5ZiseeZbw91zrXC9hY4IIcp9
tanoiQ62rjwi9jGuU46JUrPxQUQNtublJNPoDzaFUcWzh0l2cAnK42RBbUxJ
aljhGgx2KrQY62SV/r3Uvu+SpIdHyPqFBHhbKuU1GiZfAZf7kRJgovWBamsR
yYMoWGPAfFKZsCBAtNhr4SFAKGdJ7oLh86R7DcE7hlvgnrULlOUsXE+8SdTu
z27wQX3rcHmPRN6Y1c3t+szzyQ8DWn4kRafXB1Zdu4HSRCeP4gaxp83Hn3kh
9lV5/TrVbJfAqpPWv/lBczx3R1StZeAxDGAz71BfP8UXxkFyX4uCHp9ZAdaH
8CQgdYMycifPTHPjwg+CkSrGdw4pcp4sSXz+S+WHhMZp/VsHCguLfl859j4N
/iwoiFz73+sQ9s5P3QY2dgGXcCBzpWD7a5nB1AIsetR82dAyiKMpNAVRVP2D
vQijlfKI1Jey7WDD5ldc2aAhSLZOpgWq6/Hog0p9S4rht+zasPmX9nnTTTpB
FzPFDnBxkSBeTwZhwDgGQKtgR7oHP1ZsfIc8GpeyEnl6F93spRE3Ihz5Ojae
Mm9rPj5JvAclROTEhXHFR3/YtB8Swi9xj7rum8b05o0KwyScbQekOOJhemAX
7mhuxt5GU2xVb6EK1Jp7/cDYgcg6gRzevJRKE5TVkvtEDTdlzyjYpquhdfMo
V2S5f1uDcb2M+J0DE4uxYhGDmyKRyrqk9w2fc64Dr178yaHS+tXAor7X0hSn
FSXdxc/L0nFwj0q+f9A5XvntEbNDsAlOWTbOXOvRAepouJwV5l0zfdQoa85r
Ho7AkV0Y31JSFtkNVLd0MWuSH7Qr6TZbI0RCaEkL1mIciLRtyBajWpeQ9Fa3
sn3R5Ip7GjSWVVVxLb1KgVY9v/tY/weyekTdBypCVbVMX+KYMEbVuBUGm6TD
YwZBo3l7PqL74NH62z0ub/gU2Dye1XYT5Fc34zjnIMhRJcMf8cDXmVdpc8Fl
r0sU4qoLsDa2Vuw6paJrBe1f/6gOT0MyTBp72CMAb+r5ggRbdIW6VTDF3bNM
2G8/1GD4UE2VakoIOLkrYVZ6zHWHmenwa412LdWT/o+tPX9RdMPzOrSTcHpK
s+LslMI3vnwzMiSKVU47uHUct+GRBDmerz3vhM+bU+Xu4gByq0Ema9W2KQ5X
+ielhizhaD4lukuBkHsG3jdZJHsSJlyW0rjgR3MDmBEJeQ2x446VzuGjARvt
nC9hcaO69fohNIoDEUyMXmoshhlws+pM0yisYyc007l85/ra0pg1XATg+TOR
I5R64juLSAsLssn5eRXiNrGslTbYEnjWWP6vSzqdejFAehNkxTPGgw+sXpVF
JG+K9DzpKdDqJHXpeg1xUHMyX/EjI8GmdAmgiOauS9gotuKCTqiadxWCEpTz
Q7aeIwiWCj6EOsYKz4r6dVvfA/HV6eK8vC27EFObsq9OJfsh5y4nVk0t0WUa
kzhvLxWOy4CuSvL11LiUNdWy+1U2KWW6wyEHohlhmhWS7juuj0UTs8Js3p9H
3r/5cAT0BlQCcvECrA8jmzpsLS6NCLC4MEE6fMJTn1eVK75HjIEWRBVFBdjO
ZHkVcF52JHHSQgnXvt3avaA+joHlM33d85XweZeHuLu2pEoKKAyLUDp9MEr1
l0DN8FM+OpG6A9V04u7+np0qxyhB0YzJQDBm/L5tT6hkSgun//fTUR3TC2n/
B41HtR8QwEojlaQpMVuYEzjHghApGdMan9ny4iyapcPhjhSuCcIKzXujAT8u
O/rOgeRlqf6cowJuEVEx1e4hd7RHkoQnOYqiXewlFxSDAcd881oQZ7Wg8rqf
tPyHunZnY7f46DyIhBb6PSjm5+YcB8YBazfG6PZNiDgQVOQcG9wS6r/JlxAC
iNoNMz33Wvwrr6FpV1jy4bbC2ncFYHfvpeGI3HxbQc88MlldN/JrP0e7aDi5
yjQdtpWBWmUSwFfaEXo78PnavVc8+fIZxnVgNF0dZLXh/oSimhIBAYgdDWlc
lK54F4u62kswK4JvXJwF0H5LVNAaGJEEqqlI5ywFvKe0LkmpMcp6lYe7ALp5
nEj9cBc0HQeVF0RufzoWYrIw6n+twDUoETafxEBodQTj29HQyvF4dnIyd77d
rLQgY5ljGlrBZqzk8vIv9QQ1m7+92I7Jkb/LswHh7rz9XwuKznEX780Esjrc
o36tCdJnjiL5ENq0unywjxDiqcCvggd+B9Y+tUx4Fj3natEPELngp70zoGXv
Zl/RBgyi1RrnQULoX9J6N76pn2MNwMs90jHAWhYdmq93Fhuj5SwNBDgXbRKy
S3ig+rlx5TiAz9r3o+5I9jlYWLl+3Mj5LW/jBEdxykt/LY7fZ8N39egaExGM
LFyjSH3zBc76FW0uCxPHUrz7MZx/ZqAsj5sxLM2kTToCcnqy4YBZ/SFCZYQ5
SAYdZOk7Ceb/c1RRWUqZjXnYyt3Nsvh/IVrnC9iKrvs0BbRE9feYpW4vAvvD
fWRin+Qc7J0H+OIZTeZHXxv3ziG3sYv+FzfKQe1d7J7Z+wf1H72VDPBKrm7d
+ugyESFhmIoJtRUWKmeEQ5XYK7DS/kzNZN0t0lCidPtzVrcQEbCyRMLJbVY2
SCnfW1B65tvY/sW91DURQGmTihnxcYXT284Lxe/8zrDaDYCwCZQnEwXU9osM
3iS+25rzvFVqxrAoZ9CQczm9hT5df2QWyRr6zmBK5iW0H0Yj0wCcuBSqcqir
Ys12H7KNfosFyZaRzHz8Smm8lHDLTp1orOm2cckJoia+nL2wuObt1kVxtzce
2YTCeduStzC5Qjk5BHl2d9rAosuF1dwpxRFTx7NjejBBj3M7p+JBiIJRvdc6
EwTVi6hCE1Wc37rH5Gh/nTj4m+UsDbHoKC2qPZqhjIIA3roJETtqA+7dlWep
jPkIhPmhCrFIOiDvmFBf2mCeQ8ROUSfELOA/1K/rcE6hI0zbmbkTrJuZzUvm
kywy0wt5oQ4sqreUJvbXVYipyrba8b32J2b5zixziGfZ3Qg0Nh2GxBKVzu7m
KxyFI47qtKtqTMcevTpc0DKa0YuVC8PuiFSyenVsXv6F9seyyzLIe3nCchyZ
oQ6AjjefoHCGML7izsH1sYGW6lXcBfsAbHvILJyEFPl5/Qg4chorIkXIwQEp
AQpC1YdcV+2jWn4JplkMrxZ7dfS+8KDhtY9HpeDDzu4HswaQgYHOo/qlDl54
dGTCzzSIZzu6n7D5wZqI6kBDPVUhGxDuotJOWANWKu7YNbxOD+iHqSZ5FeGf
NN1q8L3EpZ9oLMLfnywV3U8lzryTlxYPLOtTCSacHQIcsKjtloLJ3+iX2jIV
Gj66uuQRCl60WU8ghx7EGunyKev3WEQQZEYXc/goNq0uXHwQ54r09hpWGVl/
dWiA4n9Mhw2HQkqOm49K6yVs7LqfK+XsIxxDDCP51Bbz47YP/dUK54P7bXjG
uk2uVx6ufK+MxSmCe1gg/xlG1AILtEpotQD1bKV479WRUZLuYGGhAtNZGXhT
Uw6aQ7mkOo2iQpysHG4sgJICRUJOJK/2vacLdOeleyRCHeDCG755U+ekJg9Y
Aa1yBvitDSOAOuTKFaTdeCluKLiQz0+s+AOQ6NEzjZ75UjRlrjBknO7b6/dC
mI8I/sACRqQRkC4Jr+//b5JYeU8qZu5JiudCUqCaW7H8D77ZroG2jP+vJJvb
2moeyZAbJczw1CLi0OAdboKYNkNiD1VKlL79nzaRwLSdYmrCL6noCpn4qloU
yykoWWvtCFeOOMbxe/4U21WPvqwFcwQMj6jQ+RIRqSg+jDhVj4+OgjOsdRRc
3P1+G3giziD+txyoGJp77KV6g9BgR5OWNHFC82ssRXwGi/s+SnNI8/beP4Ng
plXmv0hvhhiiSO3sGnelfUa/TI4yhn6s04sruVfDgQcx3seC1QDyTdUMt5f7
Hy6ZvBavG5ALZVm2UlvY6J9oFl/tPW12qZoXGkWgv54km59UC/bIzKvUQ2If
bW9CFkYldh43haYE6evg+93NwDHFYMoGGmu2Jx9WUGmsBTNu54ejgVRmKxef
NQqZi/LtclmriiacyG4rxnLB/PKgVa9GQAFIx4HIa38IqTE1oVAWkpFIqcEm
N1/HvFSxvA/C8LjsBmWzHl+Z0RjB3QD/Ag2Ho6rvuzaMfeq6suBnS77stDtK
B7rNAd07/ktnNgea0Dj//M3rHRaM+kHDXnkkbGeqfDfgBA1wDMlzDcJfl5fm
8b0EWUJPi3BlY9ck1at99ksdaH4WRHj3oJmMvepVraGzGtuX3odz+xLIx8YK
P+YJPEPzziWG4KzTnF72l8r3+VTyMkLIdyZcNT3Q49NDeWwUQF/BTSi3idxQ
lU0ycocQPLFw2SiR6IBIBLnB8R6XSW97Wu6xn+6GTIrjlvwlGXi+WRPUImHs
hbfR1PRj4pQn5dpV+aToNd1Gl27P2EhvVn9v6fXh6UC9f4H0/CF58MZhsFhD
kms57txiNlgcC1x9g6fyg4Sai/GyTfPJYQKnapCU5RI+7S2ayj4N+KZmlroS
T+1upTVn8uI+orjIDexIR8fRgQoF7P+VDeyGc0QAxHN+wWaGk8IItbSYt1J8
4F7rVDZyJFw+yH/O2/QrE5py+2ISdmNboxvR0JaiiOqf3W7ZRFt901H3JwLf
1L64Qi96l5MICANDsqeU6fEGTGdwo2zcyVjIIhkXVxPBg2koAAhSO8bDGCHT
wxgX3kMY1T9wfgwJo9FPIlPJ3Vb9qkOkOM0yC7symdTFhBQblOgOIfkD/UE6
9ElZeoQ6PHKWEqV63nqANAm6r3SbIQTttlQpcf+jiJri5ijMcxE34x3MmZPE
yCSpMj3nnN4qDHLgq8XSL5I29bYcQYRleAEyLoMTS83EULEIJvdWetNxjuWF
Fu0PJEDtR7ZBZUClEvORoqZsQCI5/lDkyG6ngXKiUEoh704GJYT+C2jh57Ow
mj1tusRr0IEToEUcj2G1s5gbYwkpzUX4Xkv/+DdsWFF+yttUHga1lTqdipv8
kKTsOHXrjQxCI33GNlbQ+i/pA36emsbD9XBH2O/grPCIfi9vAtwrfp9soscV
+kZ1sfQz4skPvOMmiDbLLgRjYcKrQ3Y3tqJEp4rQCLkBBYGDgsJzUt5OyBij
+lJ3mUTdkmeSvYLAr6aPDdlnVLDSWlrKowyIeBI35S2BBTIS6/vNTPex5Xm8
ticBGEtidC+KvA+3NUvaeiSSZFFn88xQOj69NDs3g2/cBtqF6lQMEU0bjkxi
vzhsA7bZyAq15kfa+aAEI33STxtYxy51RRr8+ybnfXGrMa7KtrFZx55wUkx0
5doVIADBk5ncFBi72oso7ios9+8anc0pKtKj7PzRLUVez23r2vcIc9H9a8in
2F239wDYJghtgljXvHiDzg1wrx8+K7CcUg4VPlxxJ5ZGZO9hPoZV2HqE9Qti
JKIzbq9IYwVu0n0C07q0eF/DD7bI2CG4AYYmDpjulO7z1XaAv/ffyJtrsiuS
8lIPGIQU0iwtgxx8mLMg6wWIl5XoskME3p1gGUNYQaMWqjJp/ap6XaN6K08i
mvW18DXJn0X2T3lpj41BJayWTQpXdpvW9amLUHHjhd4ZyyJDJVPTY/praWg0
MvkadXO5y2Loj2Vf0smewjvGScNIe3vimg05tREeIsAEKaWvxGJzRJB2/jNu
vCmJEzDfhpjexS43Bvv1gEVHICT6JfaG/bLO9utdO4KwDYKF2tKLxj83sP01
fcG3bag5fCj58G/Gb89HH2dPc6KmpvunGQiMt0HdoqUm/U/LYSJIjzMXBCj2
OAI7ynSeGPNLEHDx3TrH8sJ1FALhRHrKpgW9kx4cxrp3sZNBO6KeC5L0M4bq
myYUmb68DaZEUrG27FnrcZPaub09f3SkYuMWiYovoGTbys5qojYNuafzwS5k
El9iV0fV1iaeTiUfDozwBgLKbtowZll+moSAbuKcEWdszBdBlmtRmnmNZXRQ
uu2b5dX0rr1wj0IPExxakqSIy/8xZDZqI0LUX42R1Z0BWdgEcxcUlEpouRt/
3EWhrRWvdehQQw5XUNrvJBASQGzfonoi/KenXv8Pl/pCIyloV/PvUmf15QLQ
w9wakft5FdRdLfcM9OKFBf62LpT64BAIPugdbuFPrYzWn0u+QjDr0wz6iLMU
ZyWlrH5Y2/llXzYDfqfIum6fmKV98UFvCmLpkUkey9mdlHFccrtbbRl0V4mX
jJX8/w11p2pytLAAQ6azN2kfBnFcO872O1PgZHgbKHumZI4zixdjOOp85+A8
9k22RkiBBsSvoFj3yxbNvJ/HY/kmjo2RuiQTf73Hpn0knLbFQ1n+vw82fclJ
rCnf0Pf3Gwb9bzXA4g+YP4TyBdCDGFzJzRQjtH9pKrDHvxGQ7wCn/9f9bEO+
OKUvsiwgcbGLTlJ19CgfYetT/zB5vjrHy15KVK4h1wvzldPiJ3ZXf6yo+Fzi
6NFgqCAreSypFtHv2jnJ3SEUg9vGnQj0DBGWrLBIHaXIaX2ba9GUZ/Lt4Mx9
dtSsMFHUXDhqHqToTu34NkkX2++9zLz1P1zJaQNsbqtwDOwQhtKysGHO8BTK
xNEkb6k2iX6oWK8awyHntTbRkZmg47BHA/+xtHK7edDkliR25qqDVZaSMh78
E39sZ3OuRLhwPLu2FHZYSm2sitU3FsR3rfqIgyRUaDkPIWVANljvCQGwVH3M
6lTxnRV+g7Uw6/Ab5DuXKWa8yG0wXBz3ImKjyrVNS68G3G0HnMlg2BYzURdG
jYkCPbkuAepp4W+I10EW5knyZBpbXj7oKAfTSUoqyGgbJtIYo98bqAyBN1cw
JKNslwJ7oZ+tOnU/wtfaxtgtTJRwu+SpWUSaBhxIUNl/OIWVBZg4KKxsXamy
ACLp9i13mJhHcElyAtcvuTseFa3JZa/tke9+yYcXvL0KEbAnRwBu0rbqLe4t
BgeQy34rhK+Pl3iWRXwUnmCFI3S4WTvPy4E6xqxtE/bSKiOD7c987/n+qamq
KRokT/CJn6XggehbWZMIdn8IBEvnYUZlsA1TiVFvQUUAQOVxML/VLiEzGdJI
nQZs81LdRR6ZFzj7YL+XRfDHgCHzvdW0U0KzCj2jw/WLD5l/hAygxdeZc3vX
27/rfaA4nj4JDjFny7VJUzfIMbqDfdVN2G1QE1igpvc5/6rNkHic+NsVIQv9
fQX34/2rqyyfLYMYWpNRw0b+zz2DqbLiz4rRXZwhEP7pXNYicru1nt+BOi6U
aEnuqd0RMbz7rS9WBSU3hB61E9pCo5Tttc4L7hKozZ/rchb3bN8qtSK4OU2J
DZSISCl3EGbY4NUEB+6PN8sURqEtmVou2u6pEVkxGOpV/O5kTrpN15C1h5xl
Ke9mPcizVluWrLm2WXyWZl9vCO5tKeTYVanRMDiz/xMTfdkfFeVhFbeUHSpI
EQToUVrY+HJV52ODT7MXhmtapkVqN4eZEZGycbGuOGF1uZ8lO/u6obG/rOLG
vyIZpUJd/POlfWcGNzUDsKbQ1SKCP+APVIY3O2KQbVyI2yhV6yilRdcsUQYO
3lBP30UtqaD3dyP5dh0nP6Pnn6YjLz3S8NsrDkoDr4YYOBVUj1yBR+VhYP9W
kEkFnPEFNur3ZYLbMWAhhdwsBakWtEtIb2nIyw510DpbylyImXLmzQCOn5ms
vkoNHLXeCqhj5eZGsvHQSsPVC2oCH12wAtd08TX/yjzRzuFxN3qZyB35q/cz
Nby7n0PAvDRbOaOEtuINV1nqHULFS9/uWwB334ULf2IwQzX4/uOOIx1OctQt
FfrVQhVo1/KxUpRtEuCjl7feo7+TFZwMi4n7+M2bVw+sXHbx0+M7nkn+KR+V
pzK2han+ZSN4R0jQS+oxeVgFJMEfbOoyJOwGB3eyvM9SwZTgglkoCO2lNcLW
Deh4JkuEuY6QwPLBHC0iZtKil1I/TgYiqRcDc5PRluatLytp36azLhHmKdy4
B4WGCP6+KRan8mVLrsIHquILUlbisMltpl45jwK10kXVrqE0lyPSKycb66ai
qJ69lkC/MILTzTClM1vjBRiQbILxUxjKgHbTcgaAGbA5KGnEgyaTKF0o7tPq
yGCw+JAK0MD4lu1P51yhTCGn1P7Pruus83HudAGC4uVP4p4QSPUnF8lytuXa
a/+UAGg3UoqyruNQHBFPm1/exqXIToJ4/9laAgJpjzmJ+I/NxW4ag9ACmhlD
I1EzN/rUHGETyYJ0ykIn5lxidibDtW96QO0IUUkhrLX4clBCBEHpcYo1ea7p
snsxKqI5m9MXInRUnOsgBLH/OS1jN5ywr93yczp25ZM95noHuNdMjjitJ7aL
UprknsIefNNXowfAkoZYZpJrp5rjiT8ZIC2+fxvlKoF34KmbStlqMHHhCHw6
DkUVyNudyPnbX3zJmNfXRvJsWQNTwKvck6Nr1k2SlGXj2uisnPlMwKAfyudb
/xZatxA2mi7zw/tn0d3mdRbvZI+asnNUVFzvk+535Fch6gSBB1sKMScY4CVj
QOvB/Z3WJfc2L/SnDJEM/Wl4jo3jqW0WKMrEy3WdSwyRM5mBQnAWp6t0DSFM
zF3+YOyyVB8DQGhV7oGruxDzbgnrCfC48SxsfiIIDxOkkDAzZPe3C32Xe/Pn
kuF/g/0/FAT96uisNLBb7CaZWYTMgShTPYc6exUB4Mq7wAIn6CBXaA9jEBtM
dRkYXHCwSEiJyJbDf5DLpvJ3tgk/wi96/CG0DRIdkcO4O04PjnTAcTgCrPjt
LDbg2vja7mCjr/h8WYS0V75n23pVVt8/SW2d0300q5QLHJCbRTpQFp8qtZtT
O3KwASguwVLNTbeTITqlgpHUhjVpX7ESbwrhSbPbwQY1RwQTEdilXz/nFxTj
4HqpiaBqs3KHQ8yGT1qJpnaoKCRdg+xWe8Khqd4cqcrMbNqWXyzQDp2+KUXT
eVrhcGI2pskd8d+QL8yyhv3JtaA/Fumzby76K4fluDAwbIiGcpMUwbfh251q
xMNORLgKPju8yHnITehjpBLOm8bebtFFHTeiTmIuus6VgtLtcZTU2nhI/kDP
n54eeNmuFkxvlghJKzobCxbJ+l+/QzswTIkIwP6sMBPFRc9DxLl0qIh4NpWb
FMdj94jkOWOOmrHN/nYVMBHcErxxif+2vUhkBTlCfv4IePl1AGpaVbmuNsWV
tm4xysll3I42AuxDD5LQMkiRLC9Mzwju0xQcMhQrR0iOxpPu732eCbPT8+Pd
WHeIJuODpq1Vpw4vPOAGA6lUndOOLmBzcIU1H9t+1bZQXQUkmhdLvgha/coT
2gLaHVyUsFMCgVJ2JjgvSh32ClvFCrZyc/rBi8jRjS/nhi2JJOlnVocmwLY1
3pU9VrIhFapk7lsSxf7F1k+0ptqETJUtq8/f/+PgM3/c15m4n32tP1xeVxAB
YzYDLiQCfwlyNdyS2c390AuF/PSql0U3qaZIAOFxQDd8dwTK6+DuE4wpeTnp
ZQ3aQtl+r8F5TUFHLkzl84GmU7IAn7GX16T8J56ah+VcTy382D1/lFN8jG9c
KR22XCgkTNU+FCTmP1PhQG6/naN4g1X/sIh1Msg5LVwLYIBmTYvHirmlIxsL
WbpSEZk8eyvodAFuwOaOLmv0R/RsVpHjbi9n8WCB9rhroIZeTFJUyvOZ0K15
WXPzzVsJVtJjikKe3kw9CW2qMBTt6gMXKnLF5pHHzgY7M13VhxdUt99TahKh
OQddEsYREaToY7Sl+mbZTbb2MJ7zO7bYVZWjJBp1Rf1qLy1Bc5+n0DIAA2t5
gLFYO7+Ma8zhiuNQDZhr/pe92bg6TKMkDl0Bz0CKJdzC38wAxUqnZPe0oJBI
TulF0BhJOkVfdOV9B+gtVYvsQ4vKrjkI89L/HdddQvtjvyC8DRl3CrJ9kig0
ZhfZmEtXzl9G4l6Gi0RU0yN7mBjfimtbKFpFtMtDrI/k8P7h3cB2C8nDr9vP
t4bxGYNvBowzvfSkhd9neIH6vxKWxyRtUCc44nF8KLMS8qDXz4LLq76AwfJq
6l7iBm/pVeMiYLBivXZi4co/tovLP1jmXTVkZ88HF7G3PYTyF63jy1zP2Le4
UMT9d7rNdudtHJ23xiwR0vB9hmmadwXzdwUh4S4x6wkMMxjehpplWGKr09Al
89Y9Pabt3/weEti9+6qR8wGu8raaKH1z+VJeNBNoCBLhJv02J8j/6+ncMdyx
x9MeEI3TetVBd1iw5PWfydFg4AxVAK1CUnpwKC0C6S5IfOD1ZFy1LQdElbET
QxRZefWXPlv/oP2aEH4AQDRJsVn+kBvy+b0ZJFsD+0+09f8VsLg5pgcs1Iau
PQPMVdSeRtlGwzzL4+WHCIX48qiuJ8y0qvEt/TN+r3edMoUc40NlPC8V+AVb
Vqo+7QnYYfzzz7tZ//GkwUrIsE1AIbAmFyIBvcaczCuh1oj2FJnLL3WZpDic
bH7oUWEpoYbI7tSWiI1henT3Po9iIDxZC2Dv9eblQqC1SfqolcnpcuIkQDdw
lKhNThLeSYnAonmspThMCGrj+HVy2UkTWQctZqMSdBildNQwiX5SHvufQq74
C1RnqvACBbtRr5FYhlsaRfqyfaZy20DBwkN3iQkULo/s4r04cnv597egwczb
vedOudckOrLqtojaHi0Z1lwifhzU/KC+W0fjJQmOt1Ayjeu/pUH/oGNcMebh
AFi+qjyE1ucPIzsOdP/d3GyR2qC9sI8uBVUrOK1wNMubWkeNhgtY5dTMipLS
hGLX5pLEeRGcHDkXirRulcW+3Izq9A/h1kaExnQVWLVXTb+0NoiZOn4ccXvv
eDPQSMSLbqg7lVUBp9/6oPVMEa9DVHa58zNIXvkPpJpgRh5v3wD7qjzWKN/p
8jH20+Rf9DsF+ypsCayyBQ2Yv/3d7fLpGZJn6v6fRkyLs6KDqNuWPD6PQkzL
dxG6nd+gTsJvGJ/x1PbfLyO9syoGrDjO3j0JE5MkTPt1oBHaDX0O+qZAo7x6
orBmQwqnBIGjLhT75tqT2pg6x488yw3O3YGleYYHE3wovdnb3UnDV4Wg6Sdg
0JzqBfvqloO3AzeR0YZ6fnWjSEO66qRVp9Dn9Q36HWVDQwVLYJwqgYENztTo
Le86LjP37xF5FOPZ5g0fFj9z331flFoNqbk2M0mxlthgBV3oamTCJQIPklVe
AFWklf5p3SETz65CACEvvCVk9o4RPtyK+tD+/S5eX3jyErOXM40QVRZzQin7
r/3cssOLAArcvi8P1qftPyiqTfyoX7lveYXZYuw8SMHRzkSUCg0i/d9W96lH
WflLvFcaP+VZyGikzTUHeiIWdRiu94eKGSqKrdQSov5/cZa8VzFoVQpd9xVK
XVutxijZ2MYGpQsq7BfAcwpPeIWGmOgrw6/Zekpo6HR/cHIWc46tTcKXMfXK
LE7aweWZrqZ70/y2OFglypmq9D/q22mTJPVGu0e/MocCUsMhxg4Dn6de3Y4b
nqxCGPMTMgnLQdfpLwsTcB8rkw7AYK3uH/ALVrxcJLckc9VFk8Z58Ci/5FuQ
kKmbA/6RA3sr93NmaVuXK4evwpQmTyOf1ri8z+1+xO8vltwNX66IoLLaZU2b
C0xfjHGb21cn0mbxMbrRWSyaczPxBxfdyApQlRFeSgM4bsvj1Gz8wgG+bj1I
jiyOsh9c2owjKEYX9lOmifJZMf+zYBNsH8ElBesjJBBaMPY7pVZ8rA8gKTkO
LaGy2hllgyHiWtT8FpmPXZAQNHbigQscyPXzDhLfThOEEUnSkhOb/E1HtR8V
DKjlGJKGPKpuW3wobXHxZvAzruSWLx6MAkZovqTAakfn7MLXU4Ly6Zb9gfR3
kF8dMeADdu0nxcASjH6yLcDj6NIxTSnEDBHM7B/Xtaf/6tdrqqYGH+gVVTH5
OtifowNEOdvob9dc16ekpNOUpZ+tnirA6PoZkuABSbizUIssFwYYK9Hw1Ynp
5f6VbaiboTPBzXQHoegqdvEvxINz5SLM0uNjdDKh/wp/QKgax+Di/CxlQAj8
wStHiobttHOR1Vcl1dtOmDRc+969PNNvu0GI5mYh2e3nWzsy++rXeWEkOm/s
jPUS6l0dD9IHgrG3ZofDvCqHHYxNxXFkTY8YRq4o5/fmwRo910CNiFCJRr5/
axWKLSpZTOBTCJkhBFgF35apss/yljLj3hqvFOwMA9JL3h/3iE1dNm9JM/2v
HYdkZleKcxjK9KatFctscubxeSGEMtisYUZum998XaW2/gwqRpDutB9V46nU
5g9jXwQwGT4cwT746iix5thsISclRHb9/cWKsCLWAltgNrbCOqGgg3anrEW6
rjVM8niiVpueDvt1tCpNXIdu2YmhN9JMEGu/dsj9KOG+0p8QRjtOfgID9SOL
aONn1INaHqU+bHqnYqbGmLAqmPZvu3eKK504GyWwXymrhKxoOOwczhvzbfHU
bqaB4x6cSKghDhF1c9TCE5BC9aoTolmq7gTMcxyUdAkS6kUrdbmKZsU8sCNo
8nleSVJb76+wtCQArNpDwauUVhWWRKyQ4PaBRw2dXiF93WakWblOGsHUZ3kO
7f8MvPIwu6j4pK1GBh4NIFGLTHsGJs6Ksz8MNAMq/y4sxSz82wN5aRmHXr3j
8Hk/YiRq1Ovr4639hoxTCBgmS/HvK//qJN5jFTrDE6qQoKM+LejpfFJ3bGxE
uKZ5PMi16u4z7znkRdhf7RhqYlim4ccHNfDQdUGOR9S2n3HtEv4os0papF22
c/hLyR5Ly2dkrp8jgIMGmW1arHZNUrrxK7rjmIPW/9fi5KjDwH7BUErzLabZ
i9ccMi4FxBEy47Aog5lY8nwvBgkO8OkjSfG63EKXwqbsIrleJVZUBCqQcD/c
IzIiEyyiPzx2yEHDo9aM1fSStMWoS3MOHg7p/q7WXVhmWbeiqwyUA2znOV8n
5JzRYSUhNRwsKKMBJeqO2tCBD3OF393SIRTYk0f1bilrOe7YAmcIH6e/9u1Z
qLt8wQY5QIP5n/UsYdHhHQgYn+f2QKHMqRZ/Rwiv+WiWjWYGQhLjaVp+Dxgl
bF7v5ydA57Z6hQyRcdwCyQ+iSBHCcUpSzDn6pS9pq3mqLZCV6d4bGmm9pSWr
clk1WBRWpVwmGpPeGGUPHyHy/3Atq9tGj99iQfL7YO8vXpAjzCDZd1AdmjQQ
O1mkNSHT8Y/cGaCkAXAXruAfCATTflCuyuXzvuS0kx+ye6aEV8Ci4mITjFk/
tTI93sdMrqjsAqa963FCqNNr5O4iVnwpB6P/RfkZ3myamfOryRFvkM1M6Zak
nZWWgaRO8RH1RyH63BXOlcZPUpOgdkbsQkRY3Qbvyrk70OwiJHGLulOQuX86
kWYz3jG3IKnqwuELcKPhq/WeKxlVjyf2o0rnHZ2XfetWPAF7cnTn5e0shxi7
BbClZimwnrL0JXHYKt/Yr0k7VgHjyiDwUtbycN9GSPsBmgXN1YF4/3qk2On6
bMWf7Z+HGPn/gJ+esydtUvD6o7V8DtJfoTLQt7KUPCraLBX/AQ3JwSAaB3FD
AXNXm1yhfRc3Uz6vYxLl6XGaT4jqMKGNgkGQ/gbPSnlLZ5kPfr45EuELc6KT
kigsQ1Gge5365O4BW34XMTwm13X+8imamEjbNLyr1OMtV7qD19xc8cDDTTKx
D1NqBsvtNpwFqot/qcjRWjiLGfgp6ciQFmDjQlJLLXyKmuAmhVCqEpUuJi2e
GtggOMOEZCk4OXQPlSNBF+xgtaDq3ghBCerz4gJLn+YzYrI3R5cVk2qnZ3m3
2VhivNy+wCI+MgE+Ty01+hrf0l0w1s1DTiX0Lp66NLIA3R5I+tGmFnJoD118
LPV59YXJ7BZB61FB3bPTLUvd3piSL/7+6q8Pyv6244sLxSS/KZmJe8tRe/Gs
ACy+xFlSwRuCQiNqwH9w2Zz5rF9a0q0+psnJ/udVlBNRUjsaKzgUV2BrGtY0
SC1VgpRxBP7bnBPCvI20m5bK0TFyp+05Q0cnYrONSD5p4cgJnQXD4MuJFQ4S
YcgzILDhsBmvpXsA+uhEkAM8zvs/FpgB0+7R7tHVsRaPJo/ZqpU3TS+RCpGb
jYm8aDFdiwgoOnd6NOCbhNFDdbszfuB8OKm5c0Xjpd5Crl1fEkU1CCEXfKOp
2vUTX7lXUwTCj9VjcCXt+1Mtg2CEIjVV6Qv44P9n5ois21ilApnLmgzG0xVS
tHsJqjT2wMdIrrqmCtfBb6NwzRotwoC5hyFGU+NjOxOUKeHYtY0M+a/MuzHW
Oyq253ykYosmZ4WXcloThdLHtSlbgvn4V2lQNPdxrFDY9TAX17wTK4/2EnxF
NFcF3HOzLqAOUliqJhSOiifsPboM/auxQMIquYSs93mKaPmF1t87vm8F7wgF
RjfF/EIwBRY2mOlq/ItyJPUk1ym6I8Fh47W76Gm7jCb6P0+RlE/H199kiOw7
SXLkOxatTkCc19+04LIf/FZpB1sOqZay5CTZOK5GIpDUeIHnQFQWEMx11Wto
jP4ugs+FX+1I7bnF+I20hXCu1wKNZ2dUReIMKBF4LXmBEJXzVFnXEV49J7Uq
u9MQFDTioQ4WyUPMfNE80CYCoECQ73BO70nGVJBDegoaZWyqU89GNkOKNNMx
8n6sZxIPaeIG5bqy3UdwOfL2LtnwAWMdkozqK4uIx+u7DfJt/wQ1Ul+kqlxZ
THai2WopLGsLtDg3TM8U4WCEF5m1UBD7wKV2vjb9AuArp6fzOiCy+AzWJN4B
BZ/rsTRI7qHR53fYnifrSn0y/3dzmq5pB7CHW10yPH64NzUzv8HPhlEVYdHL
l6JsgsNHkXodfdH6y9f9GwUOb2LQbuiJNbexCK8Pz0CbZTX+22i4VhPHk3p3
iDU8xOeZXkvYrPl07WusWOoN9Mogyv7JuPMeISQ9FxdnMr18Ho8KDJ5HAcyc
AkF8zxElj8YjjzLa7pd94xIdUAkR5Cdwj+KLtEYDxrb/IZQIKsyNyQFj0A2X
EbxwThEJsCxz1mVrk/Gej9IAxCZZgjK0yo2D/XNtn9N7Jz8qkuBDHasINyfl
vmMK32+LRaeAk6Z2QGTR2YvGoCHoBq9pEzyKhcZvIvOV1P4CWsUMfcspNT7k
YbprjHQSjNzK37ktw1z650EGdO/24ra10Dd11gv/MZLjP5EFe/gnWIsZlw08
5Sbf7JgOnDOvAKJTfmV/kl+vJTO4fW3xgn87sJmc9oU/LWfIm0geVasmbHvm
OyYZSKJa6FyFjoCW9JpR8RHxcse+MWLcRUaqcNViuz/C35dk6g4XKexbjRMp
RMQDCBNl67MLHEioWliG9C2Em/fxLyP663gXX9Nb9Ce96ct3zrcKdrSoCJX7
9Kqf58btVWCSEg3kl9Kj+2bx8gpI/APB++4kzY4fLX14NFyHoVg7Puei0yXW
6ZXu0dFy9rbP4FtmvGbbmduy0qobfZvFWkgEIXcsS4TsD1CeP33bZioHmtew
ROK5UvJJEuYyaa3cCc2bfo7t+CxngLyObdqswOufRzUFgVikVQpV2ts3Waa6
M3rEv3YHGLNQ+DEyXzU2TKI2bGOvRlUusbxZcFHiCbpE2niwjBP5EYieFjeE
8f13WuBRWK1huVdbQSCS0/C6eu7XZbzs4qa7x8G5beChWlqGkckSi25A7rJm
FhIye/d9JBNqRx2m3KnJSwD9BNQOGMl15jP3B/1VDtj7vYB9q1cUy1B77rWV
gM7hwY78GHYZfhoJzKOhcvML3sCZNXTrDrhMsECDi8Qx723Zx0RnMuLz4cCW
NrY0IrQxwXthAFAT2tBmSE9mTuo+BJZ2neoO7wC71aDOAiyB+8Hiv4xW7/uc
DF1rGqfDO2RO4S+dt0QLOk3dsdmwl2AOu+TJcTkVGaAQetAFXuFuuAvRR29S
g+EJxT//++HTohrldF5Djppn228ILe3GHULVKhV976GHrZGbZnHtPGay2aIL
cwPYh/zFo86/SzbovSmcZ8eamjOlFXphfl4xkn2G3G8HmUigGiVGNs/l8bxN
oH2tMk63SXeWMYwQgAN3BX/qaUzAZXZWoDVJAHCZo/ObTuAcWBAp4J8x8PFq
AiNDbr8v9ru8SHU5s7ggJNFOdAgxahDrq86WG179l3yt0nlvGlneVQvIk/WR
Vim1WTL/EZQIXYcwGMx8mx2pLfhVFqafnRqY6lgXcye2Gt3jEy0YOVB0ym/F
06WkjuxZc7o4f1Fdg2n3VpoP74VIvOGkCkylRk29pvFwrYGyfDkWENPXojw0
AqzCiFVheLGhSkjGUkUKLeLWFoQPnTyIK4Wr6o9hG9g7H8xeFzKEGF2gQcAt
5SF9679tU2gW8/2P6QQvHLQm9eI1qXP3tFm2mGKhLz9O5xxIar8W22ywn8Ni
muWXtZDl5autDAPNS/qEFRrcgKZKtoba2tsK8NVMfDS3QJwYdBCn+U/rcRaf
osS1AIhPHiNfRtMdCZWByRuLTQJ+uYhKv16RPDpwRqnJ7w5UgZwieIk/yVx+
scjJKxladbLv+Kjx5ZJGgGJHcPR3aJj5XABCHjscExZ70aCow7fU/v2wtD5u
m2hQ2kZtQNygkeFVvHf/N4pvnRCeZET+wlKX61ua8PPh2hdPZWwdFlroXQVx
U+QQg9WKptB6Z4bX0DfC3Q6q+Xun86ewT5SdmVyfUBQFdksqXDfTFl2EwcJ0
6+dbh6Tf7e6kpN9C3CjgYyNEm4yNHH12M6fPCxXF6HwrIsmkP0wonA6SxQFJ
JUwW9UkAW4kyl9HN1L7BSK2YbWB0FJQQZWJ0a8xLDEaeqYO4Bm71/Ti/x5MW
yAYxmdKpINbTfPAkkwit0VMrmpYE49OOzcs4YwlDcc7JVOqJVNZK1fOwORFV
IqQwIC73VhMlslYqXku2hf/DL1FgQItLbRobjfb3dosOaQGZMtGdUrpXY8No
uxefWp2HUHsEmOcW0kFphEQdBHI95qEUWJ0EvSSC8U3oUhP2z2t5ViSwyctl
RBEaTr18PjayHeXUU8w+XraTcL2l+Ot0ZeR2bTEahSUNOHFvsqgPpFnP3j9B
Gkckmf00JU8Fhi3FlZz6spjgEpn61nOOZKfQCYg/2yz1sDRw/BsqUbdLzckZ
b1COV/i7oVZiQrpdIgNua6HRiRbkgFP9bznJFAxat83kcmt55bx42Jh3QHku
0MWJFzdxsK+MciF+jKut1IcLl/TY+jtbL31xBxrmNPPhQK7Q0nKaTQPw2M00
rhN7bkvLyIGvY60M1aw+MFffdcDnCHYTA/yZMg95s2HD25bjiS1kMAW6ysMx
jOcN4qG8ol1ZK93/Kah1bAT5rM78vzOD1hOYDRIE/bp5EwrR2QxBfS11RSG1
JocyqfIGWNDHaBGW7ySAMVapOgQJqk3fHYf41wI1VXb8OfMK+FLpVo3NBLCM
jacWuKuNTCWwOWW0jcXXl9wLGSnyJ64btmVZPXdcPtOy0Nf4kc21HBTJe6jg
5Syvym2/275CQW3iM9Lv4S0B4CjpSb7ow6UfQhSd6pl6HuL95N/ypymEaYzq
Xd7s4xNvjliahSaVptV5B6knBudWJF1TnTJ5ZTtADeT9TzPpxz2OhoRZklLU
JDxL+74C8O4YR8Aa9wwCOMApZgqqVkpGtPQhMWOPynEytCTWlqLB/toLxUGY
NzqVAjXuLNgJeRdXfe6ErLIRZr41K8DCO7U3EDKcNrMxEm9fQc7oT685HSke
WZGkdyUufvZMMU8ME2MKa62W0+Q4kEeJ9K3e1P/u0Ot30UrFAeQrK4CKAO8c
Wwt5V3NkUVAslnFVF3Qy9pGxKQMV9dzE6ImajQ+ZVlaCkcSvTrX4fVWmF5sn
SvrP4n2HnvLvjlkLR4uGsoy/7yqy08vTZBRVGnu2kVfO6Ap34anttv/zuwpX
sSFuPtxNIkDZXXe7EM5nKov0hgExgwOPwkRgf85S00w25Lle0Szv3OezB4ec
i+XjU1OqiKpHN3M3DIOYQY6QbGWyiqdcwuF4HZFH/5svNbDXWS7MrUsEg5N9
4OymwuExNxXhSJqessN/SCjsco5gBuU63jquNckOd+7sooiDl47+nR/syTMx
OXN+YRqbiygA1H+9ATze+49/Aq+Sa7FWp6FlsOuKp4ip605PYeke5T+3y/zQ
S2rIyEKxfFVxef2BjOkydYXk3VS7rTopUF9bbuwfMYUE+IZoTMdlCO1+Ld3M
3SY1PqZirDmbZagqQTczaNveJ5siLCS5H54pOdzOFm95LX3Pj+IhGn5guHl8
5rycJS19WXBaY2o3m4OrQF6KTu1V65tYb79/aY0cimVmM7fHbQUfq2qEyCdd
2/lee2BVvryrAqJdsC42pCp85r/u86WojIfpfCSUWr9qk2kzKW7dg8z/G16O
+cuSsC6UEWRaD7/DasNkyhk24KSCJktbsBL49e9kAgAsTEGDWFhb+H9cKhpT
8e+LQQfVK8KwPHIZiuWs5srl02aHbAV5wK5iKWlpfUgLwyMgprQeD23vAIvn
qrM66v2NX11U29d5Jjh2U6zX6p5/FaTtObGX58v0WiJhFclfJBJkw2OJjsll
dgwd9CEMZ+cFe2NQhI4BOzHBvHEJI6Ta+fgB8NcVir9elXD17S8UJC7plJdV
NIde04y2huvawCk2NBsSbQzO5PrnYaiVE9asxjg4fynMvV/NB2+wDJIaklhB
amWFCGgOF1tocDzD8qaV97vN7JGJdJVihSb4v+ENfIdYWTb/tcij9eUbkL4T
tb1gkFX4/vBjZwbpco1yjMYPfhMeuWJZ6v75yKL9GDREYOP/n6InwfGAOGvv
OpArLk/xM8y4lxRjoOrQ1Bp1ddqZJmxNhgAMe703ooR1n0BZrurLhZGtYsv3
79BpUqIQUM0CuuPpEdVFAE1IMudB6YdxIMzLVtGyKHrwJ/UgUKB0Ct58U+ro
K+Xjd356yBBrdTLrE1x+DNulxgOLb002obU0vcj50rNXYvobDCbq0HFvape+
kq7bnrw8PINMAGO604Wd/iEK0nYwAwNcvQLVwSABhHBN+FM+IwRVyyo7XYlL
C/HZwVTX5mw8Olxujy2ChDLSNrc8VDf66udGUgeffHPUKW/xfn2wuaZq+aYT
MRSEBRc0fcR8trMfwGPjckkaWao0Q7F726vuGrRjQDU+QG04wcvJ/31WLF18
fC9EXOji6+0F8RXEIzCg8mxkv8nYEDedbFmFKUPslCEE5oH+f9QL/hGzG1Ip
WcFfZz+IMOlZu3pKB8YGcjZu7SQQJPTH1WQgPl5rrNzz803ViIyadcZPDBL7
3AJiZa3UHqHeE8x5EUmhAYYndvraihEV6Lkf0q3balqb4PB0vd7x2N9yctOJ
fXiJgLeCQAuNr3OvNhwo+xuxx2mai+R5TjibvE5K7kXQhgJGC5CXv6p614ji
phxh/4vLYsZI7NMUSqBmNT1RNebuwpMKUGsBT5lxqL1ZP3I3/BSXvnkY5pdj
evjV3I35Jcnjrr357t1raBDI2i8Q1W99j2u/0wqLGSnBkiKMEVaLf50/QAwL
LEQZ3hTOfaw2n9nPf7864jWPK0x9Bye/hu0G2uh7tk+FCmOWaOJJT5owEkC4
7hhBY2/8Sglf84ijm5pSyU57fufAJKuBuODw1Iy3AYwV5HQiq9xtO45UmSKB
KCRocjlcc4M8PpJjhUrGJNm28sqaoDg26arvEXqydOnTvqXO3s9oI93TQ0sR
Pw3l2oBT8UZNUGpdpQ8a5G67h9/y7IgXCST+06frs5STKdChWzWMavRfOxTH
0K1YeMNXylpprFHdoie33d2rTuiiVuQBn9U4GI4BjK0UeJSdRNCjD06yjBaH
sf6mh+xbW961xkL18RtXBGqxbxJnMNz1pGsaQi1jWd3Lc4RhHNmxFWeoVHrY
X7nSgcaqAeHE6a5hMEYuD9DIBcyVScVlwBfUEz3d6d1ZEWZf1dtVkCPESomx
DLffzxOODS5urWzEaPzxb3CUJxyjnkoOXZ3440Ko/U3+xiGrKKz3dVI5iH3d
jUOlAzGZiGTdoQeuwsY5VDI2YjPE6b1KPmcPSPtcApv/j4UkB6oBY7JImZ3Z
m+sOxB4F1KNjJddn3eYf+rI8ffwI7HG2q+BZIG4IjeTFLMPD/w2yr19Xg/0b
K684Nza1jFBLPLz/AF6RfiS++ddfYHwJ61NVHPRYYvOcakYgpVhX4NUn6Jot
I8BqhhCbOb8xdTo8gTJ4rckUXx+SF+wpjUG2fwmUEwEdOM6Y7OkUxJqhE7a0
pnHt3zqC9L2BzX2eYoQg4buY1BMlQwlU3benjCDqBwZygC1/5Ebso5xsywxL
hiIdaEucOgZ2ILogcYN7eDm0GTsPP0TInlV6o0yug/0gx6ZrYMIPeGDPUCFp
EhgwKkF4ioRnpuadjVDYrCBSu/LFnR1DrLTzxTPv1DTUg6jkJxo9xLyvGK1d
WJ4CpTWfCEb0YiAsijXXXiY38HxQeIKf70yIe0P7sZhi4eawPTnFSUc9CcPP
+mtDZBzBCcdNDPfw52jq4o86IabEYO3EGzGzGqVGm1pK/+Ai+iXDGTkH+eki
h3qJz42QnPmgh3GLdiz2ZbQvW7MWzHAa02wFvhEPx/hhkDrrXp9Sne8I3jk/
PoYISVxXoW71iYaOx/f/6USTiGLkML6RdDvVhV51vkCEKQhwdiKHAA0SSXAK
e0ImkLri5VghOmS/l2A3prumuxefwjChdxiAoQbWBr7oNpkboIzGBqVk57pY
mqukX/+Co/uQr1N0GAAMCXWUFbFt9K1hpeGKrzlPIABSg0a0GdMaSoh6F+/Q
pDfe7V2u3S8RRW3RI+RVdhuhd41NjdaBY5r1pStmzgLrcaVPkGpiCozMoqA9
WTVxc5FSw87HPb02Apk7YVxJuJK2zXx3mJusMAVExBL6PKMIoNV6vByDVqRE
aIWEI/EUO6lBNmYi6Dm61Nttx9o0nzFvZfjZwValMTGTCsP3W4+VTbc+VxXV
bxAzKzJTugjHApg1VcKQnsas4ivr0mIuVhME0Y01O/eYdwtN6/AD4If34SXr
7JP+hHQtj/ltneQztu++i3jPh+ujpYBHSwXQRFmlbcvc4m1NAgbHOlhJM7vL
T363dCIvMs9Vr/z1q5W0oFwQPwZ8gAIkeUimywwdsnFjBesPf1mL2+8M4UNc
EfstRHXD5Dp5ST5+UaqBN7+lnwCq1HxG1TD60FaDe/Vtd4p+kF90CoH3Nk/7
UiO2FEwrtkqpX1vdBVbB6yizE2fYusgIpljpbnI1ImxknmwhtNLw5a+lHh8I
LgP4ARZIsEhckPeBl7hkjEDQta3w6L4A+VQQJS3JSJtm400JXbnLTQx+KT1C
ac4Il1Q6nwfmeiX73Fd5yV7AWz1kYAcOj8fON4h9gDT5rzGkJeyb4ovmzalU
fna7ZUFLzgvtqyXpQh4kb2evvqnnuuo3x4XPa2XZmZWCrxS8pp/OGXllJy5Z
keazzq6K0UgwAtUaER4QCgUpxCPh2F2GwxGrMn/IZn263a5KrowN+aIrdGMJ
79FWUR0BccOMW2AIDvKw8nTWS7Fdf2nvwY/ExmINxK8W0qwCtnHQ6jkSlT+U
oLN88EfnfSJLUS3BZ9CZmBcqmkGdZ6Om5wA+QwAltMiXoeQ1TVpMhc9SSCLA
5Vaq7ddA8dX9GzYmSzdPEGx6Zg4RVHBONV3RflBeWlu1nhABVNVXlWszxf1x
dzFSqbQ5R10jMDc2oSv7w4WUY8hgWqT/TmOgX+SvjzYSddHJPL/QFqi6WvKT
G9LHDInXVLEBqeyCSCTEv9b5gjkgym3KFX6vTA9wkNuhgBXlyPiwKTzMcYYR
EzZn9v90wo5muAesq0oNChJPXRFezQ+WCub9C1CXsSe5pQwm6g3K/sKmPxfw
yv5u0ikaJtUdcpn1Fsi1DejyUFeJXD2RhAq9RlQ36ovcXjPaMKm5xDqkDjnB
BwA2S6uHjRWOt35TuOSUckdDi7mXIiE20ScPlibYYK9UQe5CDGGPv2oJ21h6
IqdXuaeGk/ljBcucwQToPsrP/f+ONu318j+YRKXtulfr3y2a71C0CWI8hTSc
jbXojrvKfDZZFwUS4O59keotIeOAw1M02otwwpvp8eZPpBOZ1rdhX51/3JWK
7YHzLd+2W6CBs5QxsbiapN1oGAGNDSC4MBbeXucU8R45PJP0urTMAJYnhn3D
nRYKs7IhKd9ZN73+PLDaYkiEiBoih6NXBIWWjGUCH9ayx/kPdDEZJxRXcGe2
B1wkx/+Icu6CCvb1a3pO6O13AtgqabysON5JGgiU7I6YM/Y/8v7cZM/SyVNM
mnoS3UNlw5hwRm6tw/hp48gNk3OunVgFtSjFZdM+Iv19nVv8cQiGijmtC/Kt
LfDulM8MrmyT5MXoLrxKio60hXLeCSLoRu6R6uvb3wDs/3Hpwv+WqvRYZv1T
zOEex+6eSkjjaUPfN28uGu02XaQnc5OSmnSKP0zsXrBWkz7ISfDFrQe7Cn39
KgUHLCGxmZKktXAgp3G6esKhAVOBU+Q9sa+PbeoN7WlceIrINAi5/yKgUL/c
L8Yw2eo9twHG/mI6vnpe3x5iQdKcFy7D0k0K3mL2DhllrA0BzDBzvQI1ClHi
KBmzutm1QYR0hil2S90tmf87xjmvkP2UETvRstJgrN5n5GMVYGRIRNZHgPcA
YC/Y2hxvOkNu3GQEuAYkdUKdjWWN+q/klaUfqh+Hr/ckzef9EeZMPLpPaaMZ
eY/f+EE/nnvI1lG+MYr5lcLb74UNciLyxp4S8PODTtuUfVwR1DK8qgKIcrfB
zPjbzgMDgRRW7PZoCgYPb0jZn7CLTkVUqVQ+ktzWAZRo4ZIoaz3cZTaDiZ1B
T+vhRbMJwqU7VH+Bk4rudOHigVuCb/Xd399vP6DNxrTqGQDru88jrsjz8g4S
JOR5cOJ4xdKj5nqKmCCaVIKQ7q27FAG1tyEet0nssfgDTArlyZw06PC/hZfi
RtQajjw//S0E6fEJ/W3/EptjVxkk0xc82c8DM6ecWepmspUMivRhCCzE7JaA
t2FLwn0MC31j+XFTdPH3fes6xm/PjE3lq0Oh3tGLzpONRXCIhVEcTRbX+m+E
iuUo499XN+ZSptmkSu7RUb71Hs+dfj+5/yly5m0EF1QhKxosnsHbEE7e1z+b
NdnTgY7BCpUhEHbrNTeWJ9zwSpfk1DfnlNm0/oi3lZa6t34llZ1jZDxR2zkG
9S3R7eRkGXevmPs6iH9DqQuMLv5rPtLKlbFsEI4y+IjKWKh0orHWSBJdzt77
faa9zWgXxrMNsm7YkTvY/bts+LgHlMYdt0qGobulZR3Kf9CWY7l9gmRm8n9O
cRZwvSP7QAgAHFaMfpRY27sV2NqKUDEdeT8n8RIhNeB+FpJA+2YtEZsnhQyf
BUPtA1snhBsDeZ4m0n1J+bnZ7pkq6X/qlgIjG8j1kaj8Pm5NQMUKWOKd+IWN
H/o0xWGkdKrnDBVlzGAWEIBsZA3JCU3tmDAmMUegb1qky249y4pXDCnP0gxy
y3+SlkR1XPAKwflU8xX47s0k9YZ+BhkxRO3yb8XpbA5WE7S5q0dCcGyNiCnn
9LjA9T1OXCh8KO+E9OFPPabPEBUeAvjha3uJf1TZD7fB8dYlhGRxCHvNrJjk
Bi7KBl/9CjlgzbthWBOIexYqcv2AXbvyNO+DOB7Y93ifIXvsEZVqAuyc0ABf
dyR1+k+fto0o1H42Rfn2qNxbmPKA+9Ao3CU5ZXn7hFPHpNsEgJmilWFlzkao
aeWegOoGFq8rZh7E76VJN/BsMT79LOk5J/nAvBqzY6jLkQKw5iyf2Q/CPxiN
MpXe3kkZp/yW9hy7dfMlNx46SD5pcvWd5amcsTs3FbZ0E15ZIqJx/JJNUwRm
sxC6j6NEUYDUKMWCO7MVQcHgY6ReKcHbRYH1JAHr1ORc4PVxAoHVnmxvImt8
B7nzuU5+YC5gQoq4n15Ts4K3QEUgX3kIQmVDWk/2E3LH/SvZkjnc4LGn9zsg
Cxr3C08uegjl34rH6PVEPQanOhU4wCrmV0hVUInZVNK9DNVS1i+u7KUMIZIf
x/B40HC0TMo0H/z5UqGGCVmyJpUTcTC+Bcvpti3W/chrvx5SHj86oz4YWV/s
iWx5qwP3Srn/6GJznn/JCHAzuPpa+XytqezFCPR/GjjQsmW/FNrXBQTg/piP
ttqXKRIDH4LyJZMhAX1g5x9nwDDlWqZL381z9OvyT0AbIUT3kbVSs11ViBz3
3ikjjFpnLKPWXF8ju1kQcxZW9LHQyV/ivl+DlV8sjcdoOTwAcuZL3B+x+jVT
Db6pU1Pw6yA1FIyvnl/Shp2bMtI6GwH8L6JRJ05pKkMYrZ1ovvytvr6FMNHG
YZYllUgI3tiMVQgZId2cFHLDnGfQqjXoVlZxWiqKqaavVqXxeMVY/ed9ymog
+DqPHLHWL83zwmnwzoqMB6+mu4LberM6IkuSlzs7rl2nGT5hu0KEIixdOMJp
rkSfcY63aYHqjFbWvFISUrPlpKz+J20ILfMGzG6khnbcqHGgPOTDMoNggcgh
X6tGlCrvjjoCv8DXbtsQOq8WH8oxpM8Nk1i70wit6vSU9Rp7umLoHshiYEHf
UTWNETPWiThdVwd+1dTkDqCMPJu2aH2AtuySa3II0wErgu8nSD2FPB1vpG9+
NKNK8WYst5v478Qas6FfPkdmrZ4ghCtzBavrFeR6s/ZGgvY1646yORR5yTXy
+3FwKhwnv6zLyB7FpJL8+nlTp8IPAARP3eLr8nBSydUKDyDrbzMpLDuJC7W6
c8WP7RuAAslY6Y1ihqmJbwzan5u8/AFsJ6vDI0kTgnSrKeteinF0IYmdq3BW
Sz2XgmUeJ7Zcqe0KFALcL3KXn2VOkUHdQ3l35087rflcPaeqkdu7fjS6F+kG
7D3id3txU2fCUh1smVOcU1RNywgiNl+uVkf/ppP7xNHlU84XI1RlqZj80bzA
6fAOPJNjwCdEVch9LMFr9itD/MLe5ObZOpZa5UgfYNQfwGnWQ9a1Iezu53NP
8ZKG4l4+Zdqj2gvX8hX9zvxhoqFI0jlrxodYtX0AuGbOYoNjE0DzAK2b8mXN
uxYtO6aoWOcKSjAErMX1KvSHpFv+uG64ya7fs4VVhaMfFpkzCWrlSXJZ7kHY
/tgif2diYJ2om9tHMQm4Vol3jYPoUvKNeZWqNcUSgEMJw7jWA5XOeR6q3KQV
/16T9T6wWD14t6kSatFDtrWHVoG6hBdzG/b050NJWGn/OGu3OQQvquaURdTI
X5H/FVkHTC0wjB+/hni5z8wwik+lovuMRk3RnRW9fHo2QlWdZ4wrJhTRFB0r
+uY7vsjXie0gGjNTrPEzOykQMhpWGgylLxt17+iedxONHbsjplyoH8JCiLzq
5FcjcuxuydK1Smiety2kswO/32niowa5YiUuIzTz+TsvBF9G8pz6MhymWERj
4Djx5YporfZMlGVUrvZHAPGGmj3XXFEAe4fy6dGNcguwlewGwmCnZTzNYIww
+NmD6x3QrWs0pNIHmNrlUz5NrKqxIRRGMG/dQB2pA5sWQ/f4Y556vyJZVqnm
P83eDjazusIxIUp13ybKVec6lvoVz9bokxCC2tw9pMdUlYmtnvVOgDowK+ev
GrZx3xx4cDtF1iqCLFiNs/Thsrw8ye0I5wjP2wqO+a/EWA8Y80jT77BlEGaQ
sqYjM5ak9GnKMcjknfPWcQCxcojis7w+svLu9f98WQZdxdZPIwlRoSfvOEh0
3t6L4uiHT2Ae4UJVTl995HdHE+H3Fb0h3uBAWi+jTATuWAx3BTXdNYDOibtX
krBoPHn1ezG8IC8SwjZnHI7+31MhfIU+xkCTmqpbufZgk1WbOS2c3rtCrhhi
ntqG88QXKl9IcchrHg455++0zfGRMHihZuP5+tV3WgYsB0tSK4kWGz+S5p71
cKbHw6i4R3yuGwYALanwkrSOoK0fR5JCYlkPr3NgMSQlavbQMZXq4ul67LJ+
O1nLBC1UQRIFJ0V5fsDyzu681odRkQB2g75gbd89IVyN86wZ4l5TvPHAJOjQ
QFPRWJpzqfYSD+W1jwsQMQq7eqwVNLX1blrzvayFBdxTdaOyChxHZ+jh/J8q
Br0evPC/7vLfTrbw7bqIxesr0i2kM9t0M8ZXzr2r18PAm+bfCbBjLC4YJnR9
tgO3vJylTorXenucRdDtGTvs239THId8NYOqY4629SK38dFpZWhkLZS/vWFg
DOVmj2+Vct65FbV2InrT6iI+5NmKM+RhXXw8L8cmRPzjcrQc1CXFKmpgXuss
ogByYgCP6UYPmKJLq8nJE5XW9WkXrYlnxPN+UF7EFkwm935DhMtA7dj70T2u
y5gK9vGX6IyRpJZyz2SlaGcJ7Pvcl2p2UNbNEZS3jq3TldVC3YNN9fvJVXjX
LpDrGH2pRutrnfwPvazlrq1Vah4w/7FZkrmcHTzCs6NmaEDN8iZ+AfodmrHM
MKJDWm4nqngvnjVon0vDR5p8rcZXzOnDehq7yVKe+C0lrhmElry2vdVw/+hR
fWkmpkFD9VtLED81HQxBalphpJjfhXuRdvHZU0+RA4xjtjKGm5tpVDhTZSwy
RlOWfsD+VLC+VqSRzZbVdsqSdT/t7yDG7Di5nYJA5QYukvzyRJvHkYm10REN
GBEET/bDzGRS/iaP/+2dNK/E8cBLirmwIddRILi8f0410DIQhPryNCDCFtM2
VWEBX7FmpNcc80r7lmSpM4gw57cpMTHc3xGwUP4JxRnkwGkKbUdTKXuvWXwZ
TF5eLjZ5BMu/2g2N1p5LPRwHrlYzjk8ptzMie1wSlgkQh+MKSeRhXaocgOCj
KDOQ3JqJG+pCekTc0JzvWxWQ6ONfMOIh9AxxTyqchGE9k+ACSpeC9uRE6WcQ
poatYfCvd6LAgiPYwORyAkp6Db0An7Xz5qv41Z/dTJyItGe7tH9bP2LSk8Ir
r/YpK+3Me48KR2h/hp9G/fYNEOmybY/BWFVXhXLLtPV61UfrEm4brdug67hO
j5tstsJI6eHiCT/JGka8XBywIb7no/qWrJEWrLFfGFnQbHtzffRcU4Losph4
axXfBfngnYG/vtyK2mf3W6+Z/yiWn/mj3/tnI02cvbxjwq94P0ejoPOms4sV
r3mbflUG2dNmYPszw5f30dUa+2MPx6DeReOvTr9frDKIInHTGLcHxz3LEnBH
4u9R25+igZS+8fIJ5qBQJaLR3/nNYwgYnngVAvm/H1nKcSmtKhxYrw03QTJR
IkC3qv7rc5jxRm3fhtTdsnwAOv95k70uPmWmYYKZa+gZZmHwV8qQu+HNaIPy
zZ6WCwZaZX5j8sQKWujxHhDLBU4NSQavxlJaRyC4hbM2vUmDUPM+wtLmDX3w
fPQ1t8h9GzMhDOQed6YkTNnU0lbK07Ugbk3N5sd/bStShIw/Mr0fb7WdY5M8
g99nIEDnPA7+R6q+2yB2ed0omsuMzk5DR701Z/DO/8a9gSjd8fIjxuxRPZDj
UCcl/liQ53s/2gnDFrmn1YElTat9p3FUAnivkjVe0ora/bei0v1D6NPp9+jd
haVQbemTvcxQYPQLokJj+kkyNm4LbMRfYIukSTTlZKFYbrB/ujoxeNTqgogZ
CxCRDlNL7D6hjvobzOUpXJol88KaQBDetPLBRv7v26XwGRMZ/RGRoihNrTyv
Jfn1aLykxvb6in5h6khg3ZgEx0wdJyK0wZd+WCvJMn4iiDxp1rAQdhCgtfEK
PYCtgzCekbRw5v4+xUaRvnbYmdiJUbTU6wYu4KibQ98ROi+6SDmmkK7TvzOY
uHYRAlB2NLb8y9IetPfUnjOBz0LsOaZQXOM8pbu4Yb5CCmKzpIVUyS7bozJE
KhtdN3tMVcxnIYyB9HEnNITaQ1zk+pOkdbjAQ3DydqBYKtNtiKdV1C7yY9wm
h7i4hdHjMMutuvqjlpo+GKRnHzGd0UnYwZ+N9YvFeXSD5ahJIlzbFe4Ntn3a
UgQSV600IXNt8ziA0rXkWFJvG8cJ3g310Bk0hqCcBMEcUak/muF3Ejv/N76V
WmmzoSqyu+lH8G0FcefY5+t+jKQO1yLK2Nmnvb/mNTD5yN91DnPTLeUFceG8
kz8ZJg5f8PApL0yUYxF1kSkXKD5frk9pCODUeTcIIo9dbRMospdXJ4H7DPZD
FvReTMB7P21wYAn8UsrfxIIdS5ZfOiiP8eFdJJPN6rYlYPvfY55rTDCHwB7O
f7W5J/Bl9lcoyemNbWjt5LV8KLD63yuAnaJHx+t7y4SEo5wo9MVeBC/RzIY9
RqE15WoTVsDzntRf6nEtfGmQt1BN8Mv5crjzt+bAWHwMcagiHWXVYRqypqzN
YAy8LHo+hZPnvnSQA2EwuGHhDXHryvMv2QhGq1zYrV1U9TOMbOXrxqfREXak
PDMEUfZUbXxupPAU1SjgMCu2Of+twZeyz+WyFn9dmP8uPxoiXY6sSjFyO33V
5eBlXvf0SYcjcmVpj8OhNDsgMirFLDgi1iXRSUEpHEzDpUr4jt6JERLBWi1x
Gm1FC4ClsCjbVHWKsCFH84vu6P9uObccQ0mKmktW2JUNapZhn/lvs6lemWBA
wkoCAFIL8pZwX5oZA6rVm3CUUg9xVMT3QOKzcrka1VGOQq+dPGd0j23PBKpv
mRm/cEmdNzwf3HuARyyITYkAo6Zo5Fw6sPdDNV3hkuENNjOaqqLjIFWmEZxJ
xJ7sm02UESQaNTW59YaxUyQ+u14iOzIz14CRjb/y1EiJYNpyIsrBhQV9NPqx
HBiHRvXkJwDQMy/j3a4SYrapJyPep3tSuQFcVMOEXJj2b6srXHoQ4Hw7qRCj
6DY9ZljAj/gOMIGYzg+HYHu3HPd2f62NaawrMPxJcQwCi65401HJt4b02oSr
NGXbJV0ushQKUjWQI9Em+tfXUZ8qvLxDB+qnyHtT56H7WIK6wGrrlIS4Dq3B
L2NE+Bb/6djLdnQOmGOEMgqAaGRuE31468cYpAoGLCvTjhpHm0iCFnBbbzvG
1YS1VYnMoO0PJRsGss12QZj4JjX5lGY7xoUXkuAqe+pv6bGw0Ntr8WqP4754
+TjVBZixm0J/ThaQpSPlel5FPofjA0USwwFELbfNUXAeI/IH3lslvbKcM82H
9OB8jjhtuGPXNDblWVingN0gVOsxgD/CbTVnOS9wI0cyVR/dUrIPiBX70TN6
6rXXiVMlPVjMqmCzfHhV3t14Yhh1EwcTSpmYPZ5X/uR/FaEuYbk+QyNnTa7b
7BspagT+NoUBiqNBkGVerZjamxs8cApeECSZNx37idp6gZQMZnZiU9vd6Jk/
0sx/wYitgP5v007Q2t4G2GzteMcJiY+GgTrG77hFw94NVWntn6NLZxaAj/8u
Xzvu5wQcDnN1JBXnFO92XnzodXt0kDQI3vY7ohA8L7/ybnexzYevbPpgYs3k
Ps2VVJjcjuyd8WdFHuflxr3dmRIQiP8p7fgIvY9GKKapirFwyzfk8fy4HZQH
zL1xFrrwt6CyaIHbNy3uqJJ3qND68sYiDszZ3F6eytnE/BlyZww4r6iPa1a1
/EkCm7iv6rpMfqekxYJVnymzWyEWXLtxVb5G8VZ0BgkcW5b8TIH/qpXiVdi+
IszxTYMmUnN9y1qB9VPot0oTvbeGI/S6nD7aqzZPrktfZgLjmpUSSG9quXmi
O6zZTsaR37AxewYxV2HenMFwDrMTGqBtjP3bH7cYW/wsND6wDEhYLWZdph1X
Ef5kZGVHqEUd9jJ6+UC2E45OLnQ9kJaNjveAKqPfljJd/j/vlg5rsk+W5AbR
RNvwYW2OW7v4Y7r4ImZefo8FQts9Gv603VQ2R7hbBE9rVu8AL9utrsrvL6QS
t3xx/0NjucrKiFu0yg8mYz3MFjTxgxTs0UJVSluIRzQJxEJieBOpeMjD7dUK
cDphxIIKifdSvcbYqK2KcEDHMneR8i9RrxD/yznEdwGaXGco8sJLCrYySKH9
vG9qciWEwiTtfOyNzwSPx5sA8iFRuCxSOW/o1V7aD+qDUCKQ/1lkELufY2ph
/jyPQ9LtbMbgnCv1jvytG3I+ZDoMVpXzzSfL+H/gZ44KHmJ+kM8Zo7PMjXW4
/+xdlOl2bPrMsXVfhjbSXk6ceRaYaye8eza4PVEVhpWyzI8ytsfhWMR+1IfX
RCgPLy+8Cvbe9z02eOU2ZMsqVYJ4+L1JSMczzzjq9MPTg0jyzK8Io/CNBij2
dhiVAM5umAHIGJjtO8SFzVD33ZO6ykzDo9upGVHrl08SQ4CqlulkZKUcpRz8
/iWuz8HmDVL1XY03qo8l0CNqWLPidJFTNXU5s/wQ62FlZ8KgDlErwwtdFOQS
ijAQtyMA0F6LB5yWJiOXnfcAVT5xqm81hslwEGq9w8hJhVJRMQR/wDBG8av3
dxrAhBYH2w6j84V9QJQUmP7sKdbL9H136yrHMe0F8APOlXFkZ9bi8+RIfD5p
/onzNWZ2FeR8EEtsUWhAtkdzLvuMbGcKnJVWBV64RRbg+LPXcfGnIEsrBUK4
/9OaMoKrA/WirzJGiKgqWTuSG4+ONIcaXvNO7CGpKBY9tJTQCrK7aZscsLw4
OFZAXgQNYFWi2TNkWyoPyJmSy1pt2blPQ+ziF3RM4MY3J7I346QsXwuoy01j
LY2LrWAb3PdjVVPpl3u024Fe6xk69sCmwK4tgmdbDWgWPW9YRrqk+Oo9AYTC
8kLbJlYm9ojLXmGmpYw+kPw65UkQO7oR4UFLlWRzGvBN1GF77Sry7uVr1Z92
geemoqvol6/N5yD5Nda1/b33OfrWkdyP4EfKhee1GTTD01whjCpGATH4VgYz
3gSisAQLDmOKz7hJCHB6p5L90CkdO21EwszI73uTwuvkTVLcM6WPG4yELrOz
9zYghbVCIJhyQDBYOBRtXxAYgyQcgLTMyHT4zS9U9qez0ty4OE4t/zbm8nES
x1rPnJfFLCVZ+2FBdW8xBEEsF9sK5yTUDUflD+/nYiIuw7eM7hcOzITyu1x0
aa9c6x9OCwAkfWaIRLok6RYt+Bx6x5Xuqjlfgou9C8n8sDW6xSMB1IoWXxWm
6SHSYG2ln2VqLoQroYIWx3fXmczEOGdUv0lmv6VZrAheQ3I8tEEVg7c+DPFL
DFDc+ybEuricCr/mS2MVw0TY6hnV+ULqxU4AbIn1W6I6q/nbfK/BXg7jKwbF
bYc7yTale7WoECQQkBx/jd9+Rbz7g+N8l2WNCjpGV04ZTpI1JYwxBa1wV8s0
rbOJK1bP8vJaDghO9bjIdWac5VpjN0MU5za+UlTnZoRKz8OmrvCa8SlXSaqC
jaeBSqikFhMkJzoYoytp08xrcHHeqqjVIcx1PcyBBu+q9vyKGLeYvph7AjZr
4uybCaZmM3lONSeugbAE3wF3DgvrPReYMXYYdrNpsILWbYGumtFGSFG9YkXu
cbc8IOGHLjpX8NKBe8QD7GBnGYQTfrgBTMygcUFoFDRy04/Ii/TM33eM3Ya/
Diks6cc2rSd32/djC4mxDyOHbYvVYwFv27aDzjvVieDGZdOW8Xbjfkogt2R3
g1ASMzuABiFr5i6tCJg+zlRwe6MoXEwCl7j+ILn4Rpkk++PJYhwpnNiD7CLw
0qRPkn9+9yI5dhUPlYA/m11kdzrCO5hUFfV5qY4KSfx8GhTuRXo0u8ZkL4da
4wQmvhj8SmySuhf2huW/djC8wWhpC0wrnRoeqRzy7Jtd43z6t0NwBWuk87oK
rxz/zuc/g+Uo3vm5hcqe0JP0eHibaSDP2kquPAI8WmOIH6IkjUrLxIxq78zl
4IrcJe7N8+rJJ/s56FogaWfl+S5oZryrILZJQxYQEmL9n3skd9Asm3K1dmRS
/ph719rfU0gawjJAjmtp7471VDnZorSpJTAlRKnSb+uGAWh6GG/D3jbavZih
N2uh0t9lqVuko3VZCX8Bt32dCfLcvDYF3pYXusWpTfXpm8iQ/OK4d9rZJOjR
Bx+Q72dOtrULvC4Dqwe+PQIM3xBx79umj6jcpwVfNLUedETj0xDRmhd/NUgw
yxXYEo5DT+f1B/t9jEdLQStz0RBcx02TLrLyu+IP+FKP4auEDpihOwF6xapH
BLYrtXf2C3+Yd7l3qcog+iyUZCtUzAKBBiMvTiZnLPI4ijqhKAw1eYzoS8lB
7Jz5FXFNN2EPWCOWPsEO5m5tITzooAZsNQ/Ba09OTl0XxQMzDKY2fSiRP/oO
O5T+x2ny2wHzJIZ5F/vEHLRHNde1G79RInLgDLvlF0tjmI5p6IyCaugzkGPH
gV8J2ni4KuYqn8NDaUPdQZnJ5ShKJjKTGxpOK/YsuXT1JMIQTLhoTL6bT38F
7gxdIQdrfWznCHyUpSqSn2RXdqF+tvyE8aHNdqVqxHQm8aJ/X4CBic19E4xO
xSSCQJVZw3F2ABk0UEkxgpDHo8zrLL18cZ0hkKqUYbGwKxXdpcEZ2ka40D5t
LFohSsdK8mjbarK10YYPiehcxFQjJKtockE1u32idfcVggwqOMQN32d00TL3
316cUGAGlBLZqEMTVPZSTcO64ox/eRmUs39RvCDctr0IBOx63kIRNUYFfPsU
dx/wbzmSw077oRaQ+v+ynKm2D98QFbCm1d0Z9kwr6JWy5qpFaUEMsNhZIHqk
b1/OCfgBsuy1rVrE5EV6hFi6u9v37zPlgHznfa/ptJY/aOR1P2nhEk+4FpVb
SMQnNQJeENvEESv6L12fF3sd+/zVNLBI6jZnRxr8bgbzTzhVR88bryxW+7bZ
ozPt14PQIB4MeAALRlHoPF+yrwYnk5M1XsNZSFa+7BJ3bEoHK3NsqeU1TlQb
KsWLH1O3VvB/hMtzdna7xwlGPVUimbGtiy0T9gIYjY6ki2zWb6SCa9+H0pJz
jFvrccwRTC2iWr3Mwv+64acD7YMljyQo5JlTcdIyjLLkkbiyqhzkPSricjzs
2XEDDRgvVJV/i8WM74MxQfdur6hjBSNbgtdNgAuwIgCWBiZ5d8l4tTj3jSpJ
Le8a5USVVTqdJFhQUgkXTFL9w/3guuJlnszPu99rvBvaCxwvE9uZ5HCMqKyc
LH+ucwWvdayks1+LBmUVPlo5J4ejMi8qparwSlTGVa43CjochshLhPryOxgC
sW/VLo2+ym39+AP24DEGXMDy16e3CwmdANvJZo5HGz2d2JHq+/9j8wyU55k+
kqNMIPGt/SeO2eGgFmwPyFYdY0w6V5yH196YmGYWsixXCb+ooppKeQauV10l
lKDChsidXsqLYJXjcVbXlaoRPpahtbln0it5HaxJ54Zz79TBTTByAfmf59pv
C170EZya+a+F1AHk/rdCmic9Ka0a1miuxAnRjMB4IpJ6I7NWqi2v8riQSwJb
OjxSg8jBIYZBmZWPGIpzRBZgPa1Bb6D1Ann4wPOrR1RrjEdIj4K6EaMBOx2C
ViQCyiza87bd60BOBvsHgVJEVJBT9CXWs9FxMVDYKelXUWttG2k06FSxm8ej
dwIft7qOxIbeMld2UFzyCTMoU0yLF/+mhcyBxRZ8GyUe2ebAr8OuHmg1XTH6
qdByLhsB6hRj5wo7PWwbZRj/aHxxTBhljo2QyGWzOQJXs/yfL+rsn15jS23q
Z+nC+fjJ6rLT+O6meWAWmcoaf8ZOGeN2U1v9HSbRZscaEDCao2pHM0iDSEeD
UnmjT6/QfCmgtwwWw9wUIHjqKbjTDOZ+VC+RqFqzZ7w2ouecUlK3paB0tzyr
xgTpSYwfL3T+Wo1OqEc3OuvDhjaiNGPU2GeL/bisBpwkfdybhR7yHx3PcaxA
LQH4yfLUnP1P9vi8CtwaAadcC6w8kRnfo9CoSqFqDp+kayR1+Z2bkXsM8Jrt
4SBMYqSzGoAJavALmU+Zs5AiFbaHeRiXh6nKT1bF9mdAR5NCTQgX0HLZ5Csx
+D9KpCZvr3KrmDN+d5I4CXZuhy9aUE9aQRXZpVjvZyK5AZVqduDxOVBarDUz
qcBuHktVD4pCs2WIOcsn43l7uq66ZMT6Vbgzov2hDBWcxc5SB3YSF8Zv5CHf
NGETQbK7TbjEtkpW+y0BWbagSj/T/znByIerxBwCN4dcUVpisahBRGnfwfgG
nvBPOUFfzivYUQJx01GyvQnKNroMVIqClrjZ4l4ck8fDBuLlnZE+hTueYxGT
A4zF/MFA9i3+0ZlN9hTcVoZtRb9+B4TbLPg/A4DuAKC2jAJCzgZ257dAbw7C
geyISCeCtAjbldYacaYunNi0z0aSTJaQkZb8gk1QCDiO5i8pTfAkrId0jGhG
gC4DBumEJhl6X6pu8R3cDwJ06yP7T6WLfHTHN1s1yNEEeEuyJmKe4rj7w0FA
i/SFTf8sR8WDdSv+Uf0k2RtnWzntQ2SeJYnymeAfsODTAU4FoZ11mMoxg9o6
3ACYGlq6cafybOT1bSVvcihxUKomymYGT5RNgwaAfeHu6uLbER3SvaOq8vD2
K//tvZSunJH5gGY+h6nISn3T7gKrp4V7eGSTKCMfs1/2HXWHkt2QWCFksqWb
g31tmsbZx+/DDofeyLfZWXJFs2C9+0QFdNHxpOZ7mhtPotSJkGbekxMGN2lT
HMsBZAp/wUvNs0J07s1ctDmbBJXQMAd3prdN7Q1Iph+0NWVmQmJKOLwAwSEo
nprXZVNzvw/A1P+0slC61nFAgEOm3MBz5GEVmzxwFCs8yeg7cH5eoppVWPEk
IGsK16MKnuzXKNDcHGmBcNIGTBQht5uEujPrkYfWKuNxCwwqEZh6ww9rlFaS
S2QHuZtmlkZoOyNhLK1ELySYltSt+GmH4lwZ1yWdXyQ9eL4eySwiS99CKFNJ
1QwLVcUXORi9UBiDAVXVZkq+5QmJs8F6vh5QtjYnVd4IUHW6w3UEbZFcA497
mvx2a64ZxJ6jZhHXBQtcNZZvLGbwLwK50umz+Ut/f/gYzB/wVAarSMR7h8Mz
P0Scv55AUTW3RMfKOBKwjMRncKMdBXYeskIii3TTKcDav0FPGAXB2q37hObj
Sidw+cO06KDZHAqUnktMxSCMU0ZQCmUKtDPpj4fzc1s+GESw36zy5+Rm8S1v
a3pwr8WxA8q6psGQ3PUhr46ILpGmmSK+ifRej2smpJJ3rTphi1wW01RB0i1O
t5dSJf96FoXhlidsX067Z3B7IaH+ddEjkN8WhGbNAm3VARFOHA3y9LSpoV+7
dnptpRHy4xGrx55iu0veyMcfxC8N4oD8LAPYQB2kR9Z3JiuMETusH10IQtEh
ByOjyIvASQdMnCapjE1TteX3boCxB/hb++R1bHexouVvJKX5qP9foj0V/bru
5/qszNbUpZaWp9HxQF//99ihNtIGeg8K7fIuBthxGgTfxUeo7p5Wh+gGbaFK
OLAS11f2U/p/vmIK+udYudajqQ37F0Bo/tj5YUqQatRyk2hWL6utykEZyZdE
OhBwSsdnqUR/eApqcQRfYEFxJQMGnUyB8AyZIYXOggbDM2xQyP4My//4Z5WG
yQSCWHvD5TBmjWqolXl1IUoEbKQ+vvYXTpPa+oyRCLuEw9OLIUrSY1mWeZmP
Iq8Vxa+aqt9vnLEGGCc4OFTBLFLhD5ie0DJPmI27M9KFXtbwjwTPViok6Bui
0yV0MawMTcJA7CQh/FaDMTUJNIa6wRCAbAEMUhHcifqD1qAS+3QtLeHNbI5O
4u34ymqgx1uNnb0WmZMd/nA/gfWVGe//ygwdbvxd5D5CqJ6C41APpQq8PJVl
RjvZNv2MItftaxyt1EPu165Nqb3RpjpJU2LdsmG0Tg2GV+5QfqtKgt4z/gUv
jk0W5sCUiFkz7J+uxmETLCjaOZPf/wAPCrDSmjEajsyVOQHI1YfrIsvjrKuG
oBU66M+P+VEdbVE+RRM7Qgs0w2bPmNl4gt1WQshXqb6mvYTrUDExbl2LaHRu
BBvH4DvKrMZn7yUqJvRkRPGrtcRHj/bmVHu8uVMm6xBsHV6HC4rIWg4dRTaI
MvdAZFuEFQ1a+P9TszrTAJbPS8Nl0ZEaOaclhyuDwAJwzZrtUVtxUH8HL5u3
a01hhxr6qNRlrS+dRp+9okS9MheJcH+9LwfErr7Pd7FAYpIOuOuhBaYSzue0
W5+hWJ2CZPnJOXXfeq5MS+GlFk9OaY+MUX6w0vTmCaB9DivbAebycIA/+azn
mJfYYMvZmQT0oARPXXucJi2yZfI9NF3Pi43zVFgPGHdT+924G7psobOGbehP
xpfh06gOmAx9G0UqwiLZZdJYK3kqk0w3Fbc1C3da2DLx2mLLN0v4mLiwYJr8
lvB+bKqCt+r7EW5zDhbI/SBxwqCUNL2k+BsMnPXC63EYhyz2KHy6hXMFlrVT
YB+mp0PrlKFC88hHHRh7Ha6auYsXzd83vQIc+iUWsVUCDPe5XLp/MNCIXMXv
PCwHSY5oHxIpHog61lt+L+yN7+Xq/2/KGylEdjIzb/eFid54rNJKF5XKvmeT
MIsAnJGmkjjnabYU/gu91NmncM+Fgyd30MUwrgqpP6FYxGle8uvrValddVOp
MKGGOwUCeagXFQZMx3tIz7z7t8HgMqJO8MrR1yfj8IeqdJ9w4ZQBTenNzsh8
g8rfHB/2igCYaWcHV3Z8K1YoaWH0tHLn5Fj9GO8zJgqXxFObpPvHwXzRQS/c
ypOcflnxFJqsc5jHe7lTXa6arMTn1sA3W96gNRM4/c+XiJEZSOFiH6yhC3CS
yBeqJUwfPmilqgUdhNPcrCl8pMjIY6pxiXtiDOnpbcHT1kQO0JQrtHtCE/aM
a9wyMWdhTYAbqttSr21R6d+q58c0BI6E6UMLXsknRIgiuwLOe242duBV7jie
EUIw7GzpHTcOg5h9/n2g+i7XjtdIpYK1hxAQY6ui41flAhT8PG3T1fl6r4bo
qQc/t77HTKs3rWcGJyYdbx8k8ONxNSYDbPPW061/tuYeWZMq7MJspOy9C7Jg
0rl8QvGVBVZQ88VuJeqZYU0PSYP+OyEonF0bJToT2W7QrC+Ma9fTRwm/tlu7
Jgs7Q7fYBjvPh9OBz6dnQklB2rDMTK+/cgE0sBcbiQp11xMNes4Txa8vWeXm
nDYkasQJUsADK+v0NZUQK8axjaC7cGlgoN6XMf0DX3r33v6tx9s3coYUvGpr
kEcfdx0ob+vOv31rms1DDtd9TAPaY4y0xw939nvdFtmSPPIEWP6MebpPuFtf
vljjT4aIuKE+NTio78tBo5XGYDl1Rt9NJCq/wv7yRjuEl7xOTUl1CusE0Xo6
NyCzcBcz5EtoZApbsOpMkxB4eP4fTVEnEZ35jjWJrSQ/VN+4QjsCEoz2eXtI
2T7+cS9aQnQ7Gvh7KBfRU1n9UseQ0YUZDGC8hHJ0e4Iw4kgBUQw9g2nllxRm
qZ/UfEvl4JBxlVQgOcMVfII4GA9suCQY2G17SOn2Wn6vKXegXjRmWzv8akhR
2sc8TWIrK+J/GH5rN2hp+ds8NIp24+AE2vVzuTMX499CF0MSy4wOOKdVR5BK
xLkwJFsk5DPiCWrId8neHN9L9P1i6a8LQVWSKaVa08A6mREJpl1p0CVPPZIU
Ip66iIUJrAFu7kqQIlgNoXnrutUXjhB/PZmxaD2y4hTGdnIc9gJ4FNMuj+je
TiOzLiyGe4HyMOuUnCP/7OlkhmibQkMS5eSZwNsZ1bjE7902/l/1pnrJJQD5
NjwAZHiXdjJwa0/MyZIpWZLae9gKPsT2X5oKXbyPgSlhONAHvsCNpp3HzAnV
YfCUcHmLjHokztUZv49NMY2BydGsm6zNW9BjdiLuc1IWu6DTDNd230BvBQnA
ewaFPcfjFFZ1Vi3bb6tVbFumgwIgJ1SKalzVdAmSKoBMp/kHVYa5vJfHRPDC
WIAiKpljCKIiSYpFdPWO31ZAvbT3qspojpp6dbdPOKx2X32670YmiP2UbMdp
YlbdTPx/x3lVDXeo9CjP007Zu44fW/gNXO8LUSSyKX8NT+CkVjmJ1cY8KcAg
nhgWzQzzU3gpyN0dAR3+4ZOgsRYpwAZzzTQo2eQFjSSixpCDg7fNAsiA52Uq
jiQJk8qStb1v0GCN3VLOgJkFVtT7O51iFZRajscz8kUPcqcTTfjebzNwOoDy
cQtXUhUPvOAd/KDejFLExj3NoEIH0a9hsH+UOttPL6XYnHbjZU59FJcCs5qz
h9hLsugGjr6eQIdwGScZdzeePnKM5I86Hnak2aDAUkRXPloxIE/e5LhlIlSE
zcsv/K09oeIHrIkjKIctbu9R16Y7VtJ7F2z175PPKwQqRLy7h3O45EH7vxom
kji6bZ08CZ+O8fH2RK29sEj+NR5Bi3FhwCnLWdD/y2NlSbN69vzSA8ZcR/41
/qCDaREv+tINBnmNa734z7k1orN09JWShbpj8qjBuyXPQyCz269kkCThy8Iw
0ZAOSuFUVShCHcn/qiTN+5GbIqifEOrwUWyBQKkRIdLkg8G02Jh8hyUC3M6D
Z8XJ0VjyE6iTsXN26embTyeT9PopySZ9OvfVQVc5rVx78uZFQ4OztyNLSKRM
TVWQcEZiAx09ZrMhYf/muyK7cxUm0ttf/KsaFaSNUz7v8A1K6l665dPl6QLC
AgHYtw9LeiwTtx2H4Vb/3r8GMicitRq7I1MA9DYGMqpLE68FiU+XQg2usluB
cb3l+/Cd5UUpXPMDedQ70bc0fJ2OkSDE17TehYNJG8FBiagXuaTKfgz3hwJr
n5PB+gBMxPtzgBTscZQwzApWJGxWU+baO19DGPvoa+UNSkU2ZTXx/wsIF0HC
cHdWt4NkbVQwkPJJZRVf2uHYNuSriB6D2HNQZkgjO4mXTWdymZqIk8MwZGxF
CzBwVvf8kcedufj14YeD+dtHlfT9K97/iDzfDtBVZUqOy3nynSQEOEd3ZSaR
LMMNlZAJq9pMDVn8xX7jP9hv/lRcgCvQpe5QCcqAuZoDZ6iSgepBb1Hh9oCk
KI7Wsgpatj/W8K2nhvkKYpx1TunyWqS8jDrvoZo7f5Mhj/BrAZCoTL2T/rUp
hX9vHxFOxOyH9Q+RXWrpCDzRoUczzbxt/UTiPZiwiI9vUJNzZ1JYNtMbkg3n
QsUOqXcDD26MhifQqO/mZuJ83jxJFel0Rx4CXSIQToUawj6OANS/YQVPU82w
zQNyj5KwlQ/QXh8R1kqk4tc8e5h7FYgB92LkNuDFVZewhpCoLBiCxe+sWmaC
sKDuE2oLPtq3ugdVxQo11at/sS3C6dpUU+G0FuOEYNSQyrfTi7Ymga0syBJ2
iLlU0azCcuAy5ZZnh34hg+LFLMLIe+QogopbDbrilgGXwAZG22wMFfb91B2Q
bm+c2fxLIcmbIso1sKh1U1bXAmSva91BkG5BZesAqRV8ggkwzbPH3GiE4amV
7QCzWn2rNDzFWrcnC+ef96KgDxprtYgHcaUyQ1/xTPDCCMqpJpz0QEzYFtTK
KOiiG6qxT1y5ONaJYg1c79jJ0rP0lWuEpDyOUKRV90sL738FduSW1iIIrIHN
UBDUI4jm7/0E7bq+j+2WDxFdPDsfV2tdzi7M7C1/HMGPkQUEAiCAnrYqeCnq
acVCmFzu7StYB/HPYCifUNVl/jB2nwhBg7DBrVCgK3GJTZKgKOqrNH1xnaOF
mQINA3FI+3Zi62nBiP6n61lWYL/2P1G8wyBgjDLT+rs5+GStohgKrvXAkBrZ
NesLlzaUrCInyXo2BjdhmZw8JnxCFHuG7zPbw+olY8SrOKCjaj6a81dVTkVf
gh42bSIUvBUN8cLwHdYgdgXVDhXldXplqqh4er9PHtJ45Od1SsFv0TMTlOFT
s6LMTwc0uBSh1WZRjawE+SHtVq+jGlbWlj6xcAKwbBJ3QpOjINkd5WX+6Ago
MXbj3cErSomxAduXd4vwi+7dxJ8c0CsWZvP7zRAYtmk9gIdmaEY0gR2OEwe6
VbX7BGP8F24Yv3F2uTGHhtPOuNazdZkBaZ1yopluYEdZjQvJUVEsFzVEamka
pudjtFu4h+E5jBEkW39z0pd1C0R3tvteIaB8l6XTw/J/WMjV9GpFiLBIsCNP
UXk/O4cwKnyoORyxzn0+vxzdCGLe0jYY79Zgvd2p+JSILuAzb/jWGGihbwgO
XeYemMeoKhpDZq7g4cspxeJwxNZZp8p4nfzQHdkDVuC/r2e5yx8t1gymbfzv
QGkKZvcYAWaiP0VmgBkVHPSsIk93zMoVPGfSEfb/7teGff8teqvz+ikRvGKo
bFezcJEn4DqjCaH//MvYLPkuwMQmmSlTZmtiwE5Ia4NBvfDDx0bCZEylRTKv
C02tSlWgvkOfatG2ZBC8w8lv8GgEj0HNFYxpN76ZlGa0qmipm7fIuQYg0Dot
NdolyRQ+zWZBx1xCp89j3g299I38U+Nh6xF6uXJ+ZBTcXcW3QywVpSMjlf0W
BHJojJ9t9qSF4dshfx3GotlsPXcPDtIleuUsS5c+5QKURoB2f9VBvtShnjj2
iBBniOpuVQCmWA8AoNMOwPFMttnqbT/cqsGc88Uwn1HK0KhgG6OZMtwBA607
V1kXtnHz9Be45FOeF6CiEQrGh6DHxsM0N37UrztUKLlGJLK7JmzjFRQOpVBc
hKQsNtVSqO2mX3HE33onOPjKrDvuHnFM25sUIT6wnFa/oPHTT38PDg4YF4Mg
D+hpj+eiyn/tRahVskhT1R1UyCEqMEGTeGt6j2md4Rhl7+j4UBM44SOaK2EW
MeEx4Qi2+WCVM395bHrLjXC1Gyr7R+3YbshW/jkhxLTgZQeQT59u8T/NHkOd
b6Q6sgJefykjnMccswmGUdbWChws3mJHRr8c2RPHQyBeJiRz4bggH7K8jI6v
fuTKx+sC+O9JWaDmBEoUqNGIzyzzJeKo28ICa3vv9Gr8bB3e5msgCC/rb35J
h7KZSCR9DKHlRxIUgZ/35UcgBv+uGrdVgkR7gtY851TSMWPQfvdJaApVZHwJ
vlvof+Ji/SmciPfK0rfkQR0PDozDqgpnx5FymeSVAXFwsYrfdKjtnHDGjIY6
hXKWdbduzsXGpuGXg5JcyOWcUuBPO0ZPtGGwU793XEsqd+KJpy8GtOFK0pXq
FGihSrEFhxiMG9UkzbCavCBmib6pL9zGLHCSDJa/6lBZk1dCljKj4fEf5xz6
AXDWTZkBLinG59H7vh9BRC3ZKJ8XG8/zOjqUZ6QCYtYfcq9lek48tcPJ6eP/
jIWx2Dam/+fT3qrFAzsVLVGOGPsFmbQe2HlsMQBG5hDinhF+QqZpAk2C6jji
52UF/71t7V3CBHzlctMPX9WSa2kpiRp2SoByjjbkQFpchzqLEVG2DIe4uWDi
3X8PjFh+CeR8P8NPo3Cuh72Cd4IwaI+7jHOkezunHorKPSaD+gSLkVYTH1Yk
iscPr1EZx18HDGyDrYW+MzqoRoXbQiUBAqBdIoKzqHmcWqoC1UUygwLTdAr1
0gX2RzrMhw/vbzmId1DNSaZrXbRlR6mwjBqwxjFg3blIamQeT7Ycspa4+1rX
RQhj4oUxKESuBnzuy/4upgOuHulaPGC9S3aOi9jzs51TT5ncckNhzoGubZ7u
iaUB4Dh9Lnv0OaMxujb/139QiOjUSlEek76+hbO+/6dQY1m8XPVQRuBTIPM4
kENhc1zcYCQNRRLs42bNoIFE52CLGAZHmCp7m5CtoHPyo3Vn83gWYYOGidvj
HrDdd/7d1jOlvacQfOntb9Nj1TTu1qjyPO0pl2WK5/xmpVxy5gmUxnboREiv
o+ruyTsA0gECfmd7CVQHUX3NMOE4q+I9s3oPRg9WPRJUSU/mVD9yf3XOTr2M
8yLjahSmgOqU30q032a6zcTrnzOjD7NHMbgCv2t7rZXAW+eWbfT3xZ9yKOCA
usFqfJKiZfBWJqDeQU0ZohaRPSqrXgjB+fBtX8phWJec0JuS61ONwkC4SrJx
IuJSNaSmUWWd7P6+zQ3+GglBbfifwD535f+6Z1zOJsLPa3sg/iOmzP22Jwp7
ONRAlv7GgyNbioS408c0j8Ua54G5l9VI70bZI3fLU09pvYxvEg3fgLFkNYtU
N2iBMjIfhONHhgcKusFZoLpQ8Ym72P+62lRbS+JV8lRqoEkI13wwdBp9rOBk
zZTqGjGum/jK5sUHBUJYSSNz3LbN9i3nrDypFAgAS8hmxuPh3GE/OhMsjr9c
d61rb9GoHIy4tnV/PLC/N9WMp4qUeKbVhvV5DFWIx9X2lYDA/MJEFUxrwH0s
QDljmK+GiFLS5GW+Q7ZmNrV85T3cGhyvOsVBbJdD3x2FIzfix5DM1S+BbGIZ
UoewSJHD4S2guJFqHt+SxnzyH18n/u4kZd1z67JveZs5E4m3CIanyULxb+6I
Jk/KHnFUsPIBj1BJwFdl3z/T+oIjwvMe1M3cEHdARD4O6E20Ngh8nUOr1PRn
SCTv7sT7VBCCbulMsF0+DY1ktuXNUKvE7Wr6XPRvfSDy+hXh2q9t9lrNDNUf
qdon5uopzVhWhVImyMgyaNG4QeB5CnsI7R3X6N+Dm39BAdQtOwnswBHMABHH
GmfQHHMuW1fff7f2fKjRGnipi0UOrYVl3g3y8/eaGsqil6HqIK5ordz+Vb04
qYE7H71Ch586+i3UCaOGYWwmTWgabgVkYU8DcmByiPJKPpsjcY/wZ1JDJoC3
YnF7HVNq8+KRNnyxMFiCGrBKXX9kHxDrDg/x/tyap8irarTf/OuEijd/E9QA
VI1EYq8ZjTeF9kPIlP9PhsgwbNfa61mKXwwpJkVQdsQbwxJnbUgfleGfgbII
FGcdrJvMk79mTQ4zDPDMjnLXZlVGOR8RJIYpokq2ZHQ2D/uUOAq+E/Dr1iO5
tEr+aLl/idCClLY+y+36ZoAI5e5dV9vLEedEbUagQWEnp3z3QQH1LtSldtmz
VIY2GNgujqyW/XYCWZSOvyyKwX7WwCUPfGWc9ABOPigj4ujSok4VTEjRFqs0
Urkc10QSPDHPAlP9n0fasHL7MNrwMoisXatGdR5R8WxhzjBDQEKDz7aBTPiY
0zEmk9XBNAJhoDoi352J1J8F1lBHTe1XxfRD/FeLR/ADOIQo5KIjfwxDZ7NG
/Qg/J1UHEmJndbRRejk62dkNwAujDk7YYu9TEW1wmCdjpyr6ivpaRt6ogfJl
Nxpaeb9CuJ1SaJXTUFruI8EflT5/cLY+SP/LZB7LSDoA7NxUv2kLDMdqsFrp
u4P/h/YtXL4au58IeT/fg+/Adq+FP1KNX9dWLbV66nmTks7GfmDQ8zzbCZA4
zUH4YBgrGXAtfBCSTNlnHoN6qvFwbaYD23+wK3QJ1XFu7BWkeWjwSRuk1PN3
akioEmwzigsceL7o876KvW7KT4Xr17YKlmZux8wSUw4NRJdBPOTTempG/0Hq
jwmkqueg3vyKYckIXCqpnAuTvJ1bvU/4OP579c3ZxjYKKDvVB/sOOCmb5yMr
q6pxYnAk8ZFtbDMVQtiOtBLyxdZN7LtrbMgsXCf8xDG9yVL2xMnKhU/IkUtm
eoRi/QnHmBmvPoH49uPVPw2UzirN+Q+655+rsoENCypLp2RAs7LXQw+nB2r0
d8OglYVh0zcmcB0sfy/iYvQ6W6wRFXab8GOktn/QpnVOH69Gg5iU/e0QKrQx
NAwmFbuG6JrQmKpafQBYwzQ52vu+QAbRY+e4BGemY4i3SxoHnSIm7j4b+8rU
cX59EkkfoFh5EgP77A9G3Tcb4aG59gLID67qwFHvs7tFqAtzNeh8dNuESUdI
UGvghg4do1hjvrHVZ3hpN9KhoiDN+j0yZP5mbBvZwpzYj3xPIVZcPVsQ7uts
e69wcDoa1GxqJgrvyIrjMIpyG8UL6HPMoP01OD8L6DO1uJGo8gjTNM18/9+8
2xGqBCZQ9Mw4auxAPfR6r4gY1AlNulNxuT/Dz2m+fze0whG01XFdYXe8wQsW
nj4XuSFHHMqjA3+6O+JIPBCeZG8m/UZ66+ztEUHUIEA5rjRQ6WtXYWC/lyiL
r0Y9G8NfPtA7wW4dFjyGmqfCd7abgtTddQQZm+Uql2UpCk4FNbmtQubziKJm
+EVtfJCpZyPjpCL+ECqvojA21UdO7A8v4Q7vYEgnYPgPADYtjCvXKSFt0wm4
qGvzkwDOCcjX6WP7RS0HOoYPzZCZM+A7WywSyykiLLAicVZ3FKiOgrAWQHTo
2uBrtmA4hnp5j3y/ZyWxdgnpYLfPVK7kwMH771Q9D4xm7H5/ol1uVsABvdqe
yOBaE/ehqFYLPIaXU43EQ08rhPLlv9rLBVMuPjC7bWZt6gxnrsOBUejNBYCE
eoOf0afZRxKVNZbfYC30pITEIhENxio94G7Ezed1G0rig+pDUYhYpHpOZW+c
muJiR+lwhSg92GHAis1tAVEj1PINKZoVCnM8M4tJbwJBEjVerSDgWg+pBqw+
ispeNotqquMZsmC3PL5ihINknl7MObHBfefo+FPFKnizF67/V3WW3KFI+WzZ
yOVNNYdPmlZkXlVZ4+ySkoDXt+2CcDJQzitmHZrh8A3UqKG2L+2VpF0YyfSO
lKjwt72Wa2quFkD1cql5FpUiH2dZdQg8DuUcHgUOBt8S5VilYDjTJQgVFUV9
5Z+ouirJTetxbkkbCTDWScH2TKme5GCFobFlJdjib1o1cMmPVTEsKf9BmaJw
c9Meq02uGADySJr5neoXJEbptj+63Ay1BsPjG12XDfXDOb4seip7NsOzymcU
+XtWNcHpAogP12QcF/xe4TgKBWuXSdkPkUNpBxgBQGe2vmzDTb4WpN9dNnSC
IZ8ug5GkBXJeOmcJA3T5pKLB0DgzuWg3I9pIfZ66vC1WpIr5/SgsvizUs4N2
57FjlV+jQKBRHonsKxGt9uDB+5BhXn5N2P1ksKXad7cyNR65kb/sMAjVZjbm
sT97hVlv0u0/wiE7ZEx367LvIqIpyt3U/9tnleApTDgu2KiP8U6hgVS5/0i6
VOtxLbO1l0q8cjN8nB9UqOC5vmy2wCVZ68WipK62pNFxG3ovq67uwqqKl9NC
yXpYoUt84ZxDJI2jr1cDaJIUJxwoxvjfKIx+P3A3N350KAjHyNeGpQ4BSCJD
mJSuNSVbcNcTKTBL/UJZNiZiMKR4T4zTAZFrSNG8hOKls3zXxdy5cQR4YvPu
fTjCfnSsQVXsazk4Gb6igJORTWPrUhKHIg4r5BpiGjdau5F9lazjXjVzlQUm
IyEMphvDTo1ySDlHnlh+izJ5OKomkwD66JBARAv4yC/j1lgzS5b5Tk1gnETF
KmlTHI0i6/zd9LHmIOF1bREt3u+NCCDlQ0ddtdH/647phvtKjY+QcQiQIETZ
MeiUzWi+zA4QcugWQYLM2LWCKfnPy5daEZEiG/4lwEjyw9/3kgX6gnxcImtB
/+vlbinRsWF3QlxzGkvPLIB1QQEpWN154mUIbLq4CD6EzELH0DqogEThIGi+
QnNQEgEpHfBF8kgJg6qaL7EuUSHVFyipJVoK5k5o7tvuRx5rrJ7GdpJeRupZ
5wQ8NhZDK1ZJZriZv1sEi/OGBl//UpgrNIKn3nwgBYlTiqYJeZebNoCYJH9a
uJz4bZb/qD6fG7PqVRAT1Cd8s6M2+hYiiYAdnwbyCAs87kcg0dL0z4+7T/eI
nHAKin9Cd+6CghQCGMgztWE3bNFKV0pc5ALanQtoeVopSHGm5tT/g5ppHpZK
DTJK4fj1tf7o4O3SNMqitSgOuajyQiKCoDzeVgrmMuoh0sqNeBTEDCN0U8a7
OvNEk6Hk+6uGQjXjb58M1i0LRXJB+Mf4n6QCRMTOkBa0WaPPCOGMbXMeY+Ok
M72lCGxsRfWy6P+MMk8qU3Dw0i7lLuoJURDoeuTBESILxk7MifRdzZ0ESLag
ScNyfybMim12Ogn9Q/JQ+qdlAtDfQWG+59umOtkQ5qsEzTz4Km+QvGz4PNZC
Fl0Uu5Rox6Iwp9KAN49i2ImkKOjvkSZ8M/KthJUuPkI5ixRt/KDWm2J2o8RI
y/U9ci3K5DiNAE2WHEG5vHGgVOkqHE6MUaH6tWGbz4QtsLP4dWewOFQjdOko
XHKW8/NRrWe0RAiOoiuSS+0Mz02R6iJWr1kWUBP3HCg+to0L3zIRRLD/9p0B
/noP9fNbYhg9uEnwCB4y7L4T2x0VPGGahqg8PibBXPEzwg1oaOQFuCu8b60I
fyed/3RYCq2t19RjjMZqygqOz8Ij4y43VCox/gAzJsGX1VjzY9xX5mc6v8ug
+I1IrRd7NrzGcuKG59XyyEq/gH6oHmH34zbArFM088IJW87M0byvqUwx/3rv
K7j1dQla8l+tozt3dA3Za4zp7JXMMiU1H+WPv0rpSaqumlnj7Q3JQxc9Bgm+
rppjEz2LLl49DNfiegJ/Rupeuf+6MwDnfeobrc7/m13RuFqXvGDZ7gOo7eC1
OsLSlRUO0I+3xhrTlWd0jLed2zXo5Jmq0E+cHRSe7hOfAuZlKrQel+XOJ8Fs
NHx+n25nB/qjIdosTbJgOm3QiKTpRIyfpefxY4hVyuFTE2LgnKWtUi7iwT+F
vcFh7llJw94JlaYYZTRAp47FI4QI3EDMUl+DwsaxfCWxm5CV7VCYBF7GT7SH
Dl1FFeVi2n1uTkGKBND239Y6Elk+cI/P6XwN/h14VxHwM1YU799EWRO0mo/4
uajFYcJAh9g7/VgNFqZPJkhvVTsQ68omEMHXvdg/Zhvhj9a3ob2oV8PophYI
vSEUDMF+6/++2ahU/ORVcMBtPTMmPyi9CF8xTQHaIsPxHzPjntD47aWfOZq+
18+fFfb6LxgT1eQPwvAOFpsg1w6rojqEmc/yjRUSPLJn+i4qowBLKXOttUVz
6SXl2j3q3burwR6MALJfcTbappT51OfcgO6lyoCqIZ4pCRoTHc4Zi86Uqf5b
kYXOjrEwBpkvYuNUFfHV2n09Ykrmrm9f2PjzMcW5JFU3hh8Jur0/tCpJp/4F
jNGa8XlkLXHY48qRr+E9ypB30IsIyyzziMLqq9oZsHifpO9E/BcnoNyay7bI
6asJZLMfOGeFhIeweALtxsGuJFqWXT7Vwe7B2JyHuV+SA08vwDZP/3WacqI1
8ky9gVoXOb7hvYO3d1ThMyWv/2I0xJJ0UfS7F14aFzGKKNoii6OiHGcV4bpu
wHcm37LFkz90tm9RZstAZnW7qIC5j8vFEMVi8pqzm6EfjwM3idYO64WqX5c4
CJkBbumEpfMhzBl2gFHyKC5QmSQrFnVRmXR2fOuIIxgUhtXGkIKqEdFMSyXO
mGmCvTqMeEfC2xn/b3rYA+eS/2m6wIFvXFJdpueEoy82aoGxOXpmkH/0PB3v
RMunCSO0Y0oczGRm/QwlNXBeejBYDmc9RPXpEp2/bbvGuwtSuvNTd1Z+zU5F
APQwJ86pnKR8Zjd47YyAuUzlImOEu8xh7PD8CQ/QeW6jZtR7fRdEgOzWJL1K
aG1nGEXpqcYg5lwMpX2SDFKtouXXnPl99X1MZAxnHth3M6wOAEy4gNqsf4VG
/SxOTMX8Oz9nw+1UYxEQlOj+hdBQdinrzrkuVyFDHJ29IGgm1sRxjnDgD8ER
zHOEkEwwsZBFWwSAxZ7yfLwP60QngeKElnx2lOMvAHKRpqxj1FmLOHFo04OU
1SuXrqM8JBXEjKDJLHeScU2iUD08XdPy3w0AJIL1rHY5qUOX3nHoKn+LMAZm
+f9MUKKdhJXL6hi6sjkxTkeiMVOMeCHKthONnIivDXsJOzpeUHmgesVjScyx
EkJMSCDbmVfknBL8KTE/8xi4SqcHUl8DVn/g8BPrypPrynlc3mkOhAgxvt8A
9Qk6yjyJLjrl2X+A5tOUb1gBNV6FglNkxuBtT3InCvAeUBHC47xsGOrwAgK8
NVLbzSkKQJ5yUChu+SsyDputas8wH75tN/CKhOMn2Et6LjlHiKSswF5YgIfC
NpA6Q7w4NsfAv6YmalJnOhAgCX0gUWbmsqOhSxdNbg8xdiSscQkPpVqnRjJi
t1mRNeWwR+GD29tU2BsEco3MK+JHPPq2k6+vJcKkWOAPNqzu+tea+n26jg+R
uyRkoNFaCnC/Y5hHkJF1IIMHBw/KH7lR+OodhC2pDBdymoaVivtdgdcNkKmd
7pLg2tpzns3NwqnmsrfGsNnHvNLaQzVak9k11rm5WFApUDWrqA0i30J8vh7T
phaeAx5Z6KfYApZMvC7azQh2tR+qfhzxEWzsPyAB/I0RbfF7P2Rg6WOwcpya
gFJzDXdxUn7DH1sPvqdEv3PZCD+G6BbsbJQ0Qg3+aVMas6Knz0UiOOKy3emI
sT1VyJObDomKGl3MDTXPtNhtx0I4cL+rRd0DvmtmSuQJQJP6dXAB8dWhvDom
vt2O+JZwmqf+6HnDgPT/jVNruLMfR/WMOw768fCvg0rUPwDiFSNH2FpwNxdN
yj8xmI8e1AdTI0fVcAxq+vHew93/5us73g80867AV1mqlpKG0P6DOgFLSgAJ
EoDptGbhMqPMnz5pJ0pX/B5NvTXFFd2q3clPQ54NO3EGK4QfCFVWr9T8JMYB
RryROVIhj6e/F+mwQqzzav16knJZLeNmjXjtmFxkmbLsAWpoJfeKaqbjX1K+
GQ7JvmqCtp3iCI8eYuFGWi5tIQfbGBiaBpKmfk3YfEBX3a2yEXmbH8zjLn2Z
gL6O7hacOdCmYbRKjlFF13BAO6eL3FYmT/elTMILZdQmnbEiOATb7IhGf8pq
KsmePo16uFAxFcyFMr7XJ1RffOFu4JoKWaHN9ERCBb7u4DtW3HuB9j4eCdkd
dBFxO8M3zK7XRE/PthPd6rE54hzx8o/iyASOLj/tGGzNMEaASsZ2gs8iBBHn
vjM97eSGt/rVhmzxiKPqXVfgfU10wG3dJM0xDWdKY4Xst0CCkMiGvZLb0BvI
kkxY5OGkW4rmpvgjeuqtR3bgQisGndFmd1reYNowQsyTaxQskx/8J5p7H/VZ
fTHWfvOrA2QfJTzdFIChIgIEiMpSyK+T9D1zSnJK9Idq7OgkZlXdLfxUc1Y4
weMyag0msCAHSFBa3ukCWHCbRiwoSMB0DBPGZ4belYpnfAfMoTq9Uv/G0X6Y
eofLrCs97nkRoDixS2nM74gLw4CU9i8ydbQ9ytgh1tRlotJQbrUPouFJnxdu
iKpQuxaMt3xy6bXxEn2oHaneKOnVe7lmEZHSYs2L1KpDLyvTqHDL6M5ig5hl
Xr8tdM9FUFGz39DKC1eBqejhpn4giojRYs5ZDKdRBX/VX/aqWFcLFYbYb6KU
loZbEcCYNG3rUotoq0JBV58bvROlq7Dcqtq1/XoOhWAWNaf0/ORNXUJ9FhCp
DhkdwJ9+hl3Qx/UtO7tzQ3rYA2sluPCjsEejeOcLEw1Tv10doRNNFH8zlQq7
s73uDmJF3XjCM5wTmsrZvqVz6/4vq7e91s76Sb+Bu6xD+lHR1u2C6tnxakEX
yBMQ7X+0/NnF6I8H8kUj/9agt96uZ1A3tW7IKPuKyWMGXMy7L70/r4szuCte
rTGhw8QoxkeSLSPSYSy80DMmC8HmZE7IN2XPQHS5a6P0ggF5qE1eqHoMTGX8
ELDSfUQdgp66WLa6JdxRbVdO7kPQrFcRyqIIl1QUxt5o1W21PHFOBdMKCVSt
gCzvVVBnSiebnYOMulsYJcpUhCCKa/LGpDNYiYx1rXoYnhf5nHo7mS4Oy/kU
UHihrhy1TdMCoTbtkoP2IVS7G+LOxwhNAuiP2F6sl4568ApmHd+5OKUZrtG6
lgOJKrBQdw2XplVt4HW2uE7g4+UPeuzRxO9bIC9CAG4ka8SmsMflwG+eXZ/I
mQbeNQ7R4NgKxnmdlbSYAEwGjUYACF+sriUYuX7YPPLsSDeAR/oBwdpGCZkF
oiuywdnPHVNM2lYIIRzqIRw63+lc6M+C0VaB2+uG01BQ4F6dWM5QKSQXMZhM
6OBvV7/zDs8yhp8AA8O195/Wi0EDYtidqvYdqOU8NtoK+XmRFpL+d5r+XbGb
nLxPmHbX33wsuLewqXp+K7D02S8Ud+jY0vkeweQICFuGEyhwBXF02sUWENKZ
UXCpZ9YEsf/mxYlC666cFgiXG0SyC8xyWieyfPNKeR4AL8CTagVKxcx5vq94
jVQOIKJdaFAmQeh2bdYKgjaXfn+DW6NgutLEu7OxfVB5TCkTyCehx2m9AjP1
5yKCrPqVCCtavpEhTXXijvDk9FPObwa8kgQ9OIpPIV3e+RfZ28hUy5iRN5Qn
nPWNA75G+G/wIVQMwiONWGqNcOvyE5+aCtDSyquOtXZe1KaTrVgpakAlfY5K
3ve1KVL47WHzc0cY+ta1Hc33uCtUuqojsnb4K2e7/kOGa4TCDsTojbhv1Eoa
RXnWKwvsbmU2LbP6z1o5tqw4nJHvsy9f7Z1clADyPlX6/ocRtldMOrRD39g3
mjVPWAspwW7ENRyZCBP7W5fs1Oa4eDpG2+iYm7FrlwS3uwImC2XqGtR8IEHP
Xo6A1AG24hed0nWMnaRVAMT1ka0jR0hllZWiSYHIJbo0ADsLzn5D/0x5cXlU
OTgqhScr0D0Wg3SXEJkRASJ9iObDIce2V3PU+/99rBaqSkbkx07h1/5bLKe+
yKfT9O/aUh/3cCGw1Rukow3sdsj21Ol0Ec0pDiSduM374FdCoxlixxkthPIo
5q3FsGBFUws9ZVpErTdtUYorEoXz+g3aKs0JbLuoys/dVokIj614aFX5+oo4
uHRqKuwo8MC47QaQzrPrtGrMDqyEyE3+kz4UHHPU1Giwk25y3SZQedI79iV3
J0ZXWY5Vb8O4n3XZI64ILOgodtb3k8Chb11iy6O+dWGJDcmKcVMmf/D5/6X1
BWmmdN0BnAHU7RzzdIhHVeiA14g36dNNtuofuuXoAOWdJyKjDt7KnGQZ58d0
I1w3D0EVy+TWg518vrV3+baw9mc7szquFE7EiTvsIOaXII9ZwUPu8HLaGv5R
eLSQ8TftlTSBoHOukHTaOX9jyQXWMjrpU4UBaegacche0RgwMBX+mlgiV5nZ
bDL9fHFbFOWtmF/AhgYNvn3u7L7dcMZPdkzhwEWjV5tQB6bWDDXMTqEoxwgW
Ph0oRenShl8QpWf+xV3mFlKmkTKDa1/qZBMpLm9ykPEZwoD27RMv9eOGrkTq
2bnCt+zgko8WGQJOi4K+qNOl3fm7/KWFyQhNDDGfrnYU+Ad+8pkSuvdKuxRQ
R+z8Ys0Qq7C+rmBPQbcnr0nXpTWUYOZiWMx8oBkGHWSp/0pwtWT9heGbZUXT
fIkGna07lI3NEQNmZ1fPBtH5dOY3EZSJrhbFLh34yb7kkhygMTaGmfq9djaX
z+uS2kceKuJBjyb7M88B0E587Z7wSjIbVbCIzcvXF2e0UtosAukcB0n7i6iW
4mbZRSBRELBzlwU87J3AZSB7/u7V3n3zeV2O4IXCZCZQdFYOuQ9j/AQu7qZp
jatUtNPXkVXtR8fF9OZzJTrA3LNdcCxwjOGdoEXwB4uAByjYiBetFX+mOywI
hTCSvMA+B2rv6x9sW5MLdoPC6aeWvb/H++esEaqkjmfDLodl5UJldh9xfjdC
lSIQLvx9JCzoUyYspKnzX10fLijxqTM5/Ww2NCqS8JdmUix9pbThywVNRbTy
Id0OtHwMXbN8WRLrKRXOHF6jojCMVK0cU9fj9DHpK3MA6tp5mBbhYfb+0ZKU
m0CKxExWy/tp055Eyk1EF7CvqL1vcfEaM74/TiniENzbhCUntG8sBUzlowKj
a88g4ldjxAY/p8uJzI6n1Qumx+jeEIiS0pOKh0qsxM7lNVk7e3Ar7Z13d0Fo
upUR3zBPHnznvd8OjLn7LnMqa0cUUSeCnAf1vZVW2R2wi87AMT9wVRLlXM3z
xEGXXHD5g2xowJvH7CAcU9wmkMcY8fQcV7bnoi6wW+Q1LJN6KBhVKcpsyQe0
tI4hCcFAHuAQUXufn1RRypgkdTsizru7X2eu+tF0Eoo0XHWJ+46xuR3CYtv9
NlKMkBVa5ruFxtNdMNledoGWY5lbXBduke+wnydN5rZsB8mPyqUNYYmLexPr
eGzEJwGLCucnFSJlfwk+7Hz/GaICx5i8j5ZWHtQKaCfTIuKXRs2tS9T5a7GF
A4X34L1lh0XlBg1uELdxWdbq8m7OvB2Hw8j4vNcm4NoDy6I7PClp8nt2C7gI
JchIlxVogP0kfCXKLLYsZ6IMg1F/6vbe1q1XbXTXET8nv9XTGoVX+w5HUfTO
JNHpgnyevGbfoiLhsz8r3WHJ9uOq11vWW8M09ZqYQAP6MnAY15KNE/gHjWhK
wf5Y9NXc/xad0khbAjSCyCPZChN0DBcex7+saWuQb/VYXrn+J9jEoHm5Bs5i
e/Df/PSBZGtdCnAZ5d2WJf2LcTYfdfFt5tT9O8VBsfgJocrFjPsOePX4JFob
YeEqfX9Zer6i1qgHViYXJQQgn628wsvNE6DWZZ1VlkQV49JOA3sTgSzl4oP3
caUY7yW59Ro6LSE/+crjDXxxxjnl/XJRg7+98VHnqnux8e1OPw9ZGHAMwNSf
KLYdgPW8o2AKp2foRtd151VrnVKN4q1fao8tPLSUakneKoRKwMxvDIKv2y7p
saUEWujxSzrpqOdttt9Wue9wZJY/P8xY1kzKjOfncNIUkbvZLvP8VJQRkO8J
gpV3FI94i/zf2/ABWlpDfUbSXbc42MNf1jVW1SG0xo23Dbc/JO9siQZu587w
fA/Z02LTRfj7h8HnuvVYSyri6z0vARnx6HDPJ+EbEWEI7bffLDHZ4BK158Lh
pDDvBmUfBlhDUztwmDyGBJjqF5jru4n7miOABVjVttY/MLAXk2PEOFvwrhJr
hK3iywhhZAbPd7ScMfAlc04O0jdlAIJ4IQJ/i1I90alL5pSvt5bb0/C9VDxz
UlMW6zZnr5jG4rpwVETAJzxpRUtO4PjY6qgSrVCH1YU04Ga6ZrnFcCBHKGJ4
x0v+1Omo9Z6iBI/Izmbn2t64qWDJM5GpsgN/ADz+gQDxoZSbO+fsveVtfrz7
8rwLXhJd/ZVUGl6ZpavkbdPiO2GbgAD3IX0opLNrEcsrjOrnHwSJV7uZGMCH
OhThRa2hic5+l7zBgASjFpIoCi7FREUVkDAE6dKFxYZEiXczUoTDRdFoDZro
ZEbJARsZ7jiOLjZwP4BCsdJmGcLTzE9nUMeoDvj2OwR6AI3YWyHovFBJlUrE
Ms0gS8gd2ctZ/QzUWz+zhMb8d05rfW05mFZUpJHPwSIyEsJFyKl8fAT+hHLb
eDSe+S0l59kKP4+DKIk/h9mZxKIj+yhgFgcT6ROPtZ2/4x32Iqepi6dFVJ1/
b4HwqkjaZvHaFRpRy94kjxyTJyfBo/suIh6vI9EglhuNK6lKjmv2p5HxSTqV
ZswgQsPTgxODehrqjsFzCZYFoVT/XYHjlvBmwc3JbzFZE135dyL+7wvkZgoa
bbWiSrgR8dQRsrNOVAlmCVWUb0IndwIOCUjpVyZnO6EANu2UlPKqYR1/tMb0
hFpd61E4mdLi+NIZQe8Ca9YiSDqZmbJETtFtFlr3qqaa1lM0PZOvqdGTQf0c
rSXzdw4PhchucrrxQqATxl2emGCf3AawLcTNJQIpsoGu4H6d8+eqUGZmO4Xr
yd0BbvktPi8o4vTVgpkgY8PflVNMB/zCoVfSlENpyN90Z8gVXL79z1XovpmP
Fiun774/1cAp20tvvACS9aVdSy1jHLC1LMVPDilQcva2owZOFOG+oV7L9HHb
Ire7kx4mfJcn9z1A/kHXIIBcUAtzGvz8uogebyzIN1QHnblU1qewC2vPcb84
i5UJnKBnj3nnQ2uIuUq8TBkeq45uRQzb5XwMHJiLoKd6ZHvvwhqC/IBVHUKu
Yl4PngKRwip01CD9MqifnjPFrmuq0GRBu+0O9ZvMlKjMr0KPOXTaCpn22IQq
DlnANthjjZoZOa4f5upaXtK6Z/KQ84fZJwX47ZgzSJD5qr6T8VJiZFIL3rMl
n4SI+Bk2saB4bpcgRzPQ2ZGOT3M2dzsGNNwFFxFDqapITeTE8oqyqOECcecp
DI9UPalTUESsIzM7FHM8xIDRYbqDNLiv1xi8XSQqKHbz19T+9YERDXsDwhWi
brSregwmNCo6XCmwIINaESlXk5vI8K43QINvKC+15u2FWNRgPLKCxCViWMc2
ZGIvXhkvdRL9SNnh+3Z0UtzARu7QOpXxNSUfZ8xjSb9+TjO2Wjw9kxyLQkYw
nH60KywzyQ9SPN2orNxIugvLHsy1nl1ULaFj9FaOouz9qH0pqnnswy0atbNU
nYnOme+lUGvHQ6Gwz6bsUlz/eCHodCbfrmQFywgixWTomzRjCnnFZ/f5VzwL
InSBTJs0j7rBWw0d1ge+paRs/RmijZonrEGcWfv05ZmE3k1uQLEY8K7f6Ue2
AfV65mMay0Qgzl7z1Hib6UPgJl8B6BOpxJI5ADAHhDmO3hD60Z2S/jO7sL0g
iMOdFNOFAJ1HdISfaAmkXiQrBZJlCtWH6fVP+vmrsQcbVieC3qGoA/VfHXcL
tHBXqn0MFOPujeaU6NV+07XTt3phnPtDl9OfNw0vd5qnCsOk5aVLKg6+dXUD
c1S92Roup6IzFCH/+wgC0rENqYuX58qVG8WozkfFBZzkQELoKFnCLyxrwYYs
sK75NgX8hWtyGLIe8b1hNo5DQ6hI7qhUyHELDKi0F0hE5BAv9ZVfDnfxmNLX
uNaCoPSQkgqgMTAGUnLdp6NdlpbbL6w0CJLIKoYjA2uznuk882yxB0gXuFke
25uu5l8tTw831xopzRG6TxVh53BcNC6ss88imcnO8oejYgUUi6hw/1RYPXP1
F9l+3qNs1jqzvyoKO4TQ0I0Is2V7n+AbCtbuv7AwgI+E9EKlCyGECgMvYiHW
POZR6bCFl2NGBVfsdmCGWdxDZNgUR13Gy76NTxX2GjJijfforD0kI7PyATZW
QhCAVWR8wAJXwuT9ZsqRIsrE3lAyY02ggxO/RaELaclxlh6UkZduFnBIUGK5
m4G/81bzcAz854Xg5Oj8wONXcjnRjMPk3D2Eu1s7SucFfa+AuiFQXmjuhnKh
/bwwEOHnv2dQCkDFeb/A+syfQ5zNqForZINTYxbqAp+VzbhLPh0MQhgrqEhs
hSxQP+K7AegDa72Pl+tq/jTG/IquNXO+rNxJPvStmwkwvtFWMneems3986Hz
okwFwZBW16mc33EfyNdpV/ahNmEkcW5bFJStyqFtSJnAWoGaq+5KrRJ4w+7y
FBVbPFy99H0QHrVhBRTwNbkqOiwak3CTh29OTPOD6iWde8KqBcLMVMfceLUj
N+tQVS1nQYpIegLTd2WWcEaKIIs1gO87nWHylSTVf0cVIsroXQHznSBo60h1
XAPkYVwmGTuwQh3Pj7bUnEa1/FKLuZCGiDLi4RtOOljidW5TVsGYd0Fyhlt6
uSoB+67d1kJ4QMYrxlStqRIZxx4gJc6XkBlsWCUmMzPkh6X5vu7pehbfsIeS
clxoCIyHLMcb7uJS1Q6o6CJnAWnmsppiDcXQuzhYU/6rSDOvHmJzk0OYN5oh
PFxSWXlFwd85dj1dqsaiL/JET+lgfsto05aCBL8h0JBR2i5zKnTwXdaSlKYG
n/RVJTinhOhoIjfreX/fXk1Gu/2Lx1yXuTTcnylJHScsmBia+S9wks8GJZ/u
EtS81PWTpu5gCJLwVZePH61F9OF1d9jlYylk/4aE3WrSqXtyhTRSK16j76y9
pNFBG3P88KnQJk/mER/w4xGztxDf2PQSLDEwoLCNTT1COGwutuqLSj0gM8s3
UtATXeftcGzhTaRJxclJnN5PXMG7xeEdQslM53f1B72BeUIqqE69iC8jCDU7
p2c8J4gY8HpQiOs7giKHZNlkk8wQm4uY7r1UITPzcID5BKmuCNHIlTPVjGCp
AguQaUhzuLSCXURbR1jU7x8rJDqvPj87Xwx/Byc09iRnbvoApsbV8IQGZGrC
IX+M3O4VCCAwMlGU/+14Q1ZCVLGjSiJY9D/OmwGFiohQf4ofBsoCcBQ9CweT
GAEz3WxzXOC0qp16AbPvCucyleuJKQwjuUO/JKBye3g7zY7XbraiF+sTIYbt
yRHvJZoh7Nk15VYpks0CtXnO6hv6Dl6hkhHzJvFny8Gmb218GyTutPfi5LRz
X7ydU28RvK3h9j/lHGX4la2CRLnr6VywrUnrpnMkODvZvukKRU35p6yWo6SI
XQVfusxNYhLZX0f88hYC7EjBiHpIivTMPBfAOd4wQ5WBMm+xkdO2pUgueQnA
Vtb/Bw+/Xtfu2nCFFOjJ03OA3opu9kzxRUNrR85mjAHn0dWXgsgXU87NScS9
2GdgWuK7q7HEd55L1vQxk7aS6lQ6jA+6tMUk8SF546AgG3LWyeLgElse5vbF
eQ0hl5cTEviW0aeE0hiTiFt4DT9RoqwLBmbALorhEnd3eQ0lPHlGaCdIt+tM
m/MykA69UZQkTrSL+5D9mK/wXEmBeNpwWR1amtCcl0S7lB4hayXMjHdy4TZD
H5XJVKC2BQsg6kHU9yxEhdTtlz5cUfLcQDJpbsdG8RzznXwJSHl4wq5WmUzs
GzNOXuF17yI8qOQix030qs3Uy6TWMJcacS6QzUWH7trqZMPNSdt9jswboBxq
R14eK9AbR1CoD66bbU3VqlQeM6Na3ZcpuB8ph4+gSpD0v3NzMKxKsBl8UI6G
I3oFeqZdjEgWdxXpmQtMZhoj8kAiqGZyP5jMPMbMs5Hm5Ptn1+KDbDLNzKD7
7XdiENX1b7+iFwaG7GmJgKpMFB+JiVRPogpv8Z8DlHxNhq3IMY87ksHpELT4
WeyasTmdqayB2HSbhMegRZbVxd26YA20+cJNoMshfgutmrp0eO+vmp8aPvPa
q0p/6c8nv8nN3N5JbMMbfNeb0fFSnie5O7NI16FBiqbpFt1kzWEj0cfej5+O
i6IgyTBCvcNkZ0+V4AtSF3hjNYQEJWfWnM6p/P8NK/l9zXP8lfERjVRhZhyO
wTMadQwiIi77lASWvUoJFet7j4QrxmX/5ApElXZFHJUWs+VJNzPo12wzPzVF
WRUy7IP0NOrubpa/FcRjeUFVNky3UCNt9tMcQl3PE7XerfB7Mexs7UKlI5kE
oC75tta1kInIKVZeYvJHO8y69LMyq4xLeFYBzUUl2WAiQlgkzqZcO1RhOkP4
Ah+tFxnD461D0PUlGZSdYoRCOGYWoJCF/5g9kIZ2Ry2l6IvYYDmggvkBFZvq
I9einQ+vjwTTec57+fNOw/LVyv20CeZZOBWYV0FtrXl/syIK7fIeJYg/bw4p
Y0clP8aA3B/XiVfes+MDxFpACUHsfbMdPlOaHb6x5a/WUfmihPtbrthkZ+FO
4EBeWWHLKfv8Hsc486CKNy+pwcOl8RUHeR/fbfXMloFFH3C2t2g+zWKOLBjR
XEdlZa3j7Ywqq3lifUNExRzsbh3j75u2xf7tcDhdkSoRu5zR5GmQum6gd9ne
BfUIBlNTCxnZASadMPqVI/mDlAEtdSXU6Z9HhwGZwO8vhXoz3nR3cQAbOWWN
7kqREoMjht3uFH6PmzIVc+UuCeUlfWyaSXy25a+YoF57nasI4pHGVuCxMFFT
6oGwlmgjFAKa57goItr/OztJw47B2vmTQO1kAIRnBfWY+d8vVpRF2kixUGMV
0Llp4wpa5IdOArM9Ikol7085w7PQgc3HCeyEZc/5R6MDquj01Y7EW6FRDtiF
d0227OSgVFN6HExFKEXkb02coRWjSJSre9LwlPP2Wk4CM+rkl8oq63MVWgCi
zeGFy844NznP329xfP7dIXnMB7dOdqcQzuO/xsZXU06N1/5a9dkMik0XDwED
LY9S1c8g6DdD4aJCFEDFjWCjI8sVmJ8l/w9EIcoSWlcg+NEoYH2KRphB5GUD
q+20FgKOjnhUf+2oseb5T7Pux7yi3HiUqvqls+rtE92rONFI+3J1pOXTCzQp
YixHTsi4d0QAcr+B7Dyf7KZHmKTUS27m1Apm2Cf+robsPCWRknN9MVjru+J0
fsI/rJGhDHy8lX+g6Yf8el9GQSGOq0RnujrtWDZDlkkpuHepILETETGLacj9
I+k++WiGX1g/FMOnBm29BAWl4hYe5HNw/cbvTmaPxUjj81CY7B1THtnqLWek
wjnhkSXdy6830Ee39FDfVXmu376QEYtbIoyIEVWAUCDz26DPM/N0R+8n4+yy
g61EFjdS34CBJ66lL1MYCCwPMlPVfHSXjaaYVkQIktCvVFr8p4jf81leo2tW
5aFchRbICbI/KWCW8CtA16PpgvdR0oJacByXPrj7FDdEtdi21pFx5QbC4nB5
x/E/l9vL9zGdQ9yT2JXm5jctNLWwN6ZGDpTf+IIAiMiHhxOjRrICSWCbTIb4
lfsvvtys+m5/7fj9FomQmczBWsFiaM3mHZcqMBfegE7WLXwnCO1NMTOErjS4
4UBiE5k8C3MBOtfsA6ptTp6SGBTWkpikr81DC2s8SXarMppwLwt60LKGRVNi
JsqKcJ8+ARzngk+z27Y3mXnOijKCX4Xo4GCwjLB5lYV2tJS1UmJOg41Hqzgf
SHYRAW4d8hSdAeZUP/38f+GaYLrwU1NoRIC8RBsIbFlxQNtkZ/ceL3J6i1Gh
wop20pxc9PfZnlyElFM9QG315optuXD9jEctB1m8HUqxRJwSBsTB9Qt5RYiX
/ziefGWjXLbP70R2PyPyFisZYBj4obAS5RGaRw61Ukxt1OQjHQ+u2NyuRjwV
8CpZLqdto7iJ548R73kUjaDA0tSWXgZmGku+SBYU+n8lwhMx+VTdZupHEten
JOiCbaak5q3MVWuoqN5qSmlael6osjYIe2QvSAtXlG9xI611adJ5ydInWLzD
w6qfxrcjlfBt/jdxjgFl0N2LAm1c2Ngy84X1VUmV/bbl2QlcGVddXsb9kdyL
NJaKjY+FrMehUMPikj6YkOLUGvoZJr7O5QI3W/BQoeJu8scTwirXLfnuvNH6
RBDDsBV4ciwdMah90H+aS5BMkoHkG2v2TKhtD6CKNLUCQfopSzxcjnAgb6Pm
b4Gd9pte64luNc7JLGxRpdT3jxegqrqg8FT92Fou63YzeCC92xbvs/or44ut
fFN30iI570pMnbzS6vnAj+aQnXPTbk1ei64FajQxn9C+1SYwV1wxUFeB5RZB
Ff1bN6UQC6mCoo5gdvhhU6I5W+I8/6DGQm82N5OUwbpXAcO7d57bhXg8zV6e
RF8gFNDC4xP33gp6WuLVLkM6f5hysRPp8hT/87SqfUU0O+2Jpp2vpKFldi3z
jZN1b5ICQmiaxQv7bVg2snZO1JGu6kUaTGuqlondXgUUx0GfhLVFJidg2OSm
EtRh0eHTs1zP3xJY7PhOEvFaKhoHLkgzq6S9NHetalUmE3FmJscxWVVwZQoN
4RxE7P4aR8toSR9ycrbT0byr6ms1ROOKt1fgUz43PcPoGC532OXpSQGIBV8+
R10q7EGXlefoLOXFsEvn+BAs8syosuiNLgBltRZHzHZtPnmPl3KFo8Io1ysW
TPWy09lu543v5k35YqkaOKKwdNdPPHVkE5vpmmvWpk+0wkYzDoQGA7mi6PDU
nVPm/luRyjZQYT/FTDNAr6gvQP9ORFiWt5NLmYuZOdWhoc9DPuCO4dI5sT5W
inZ3FkEGZ1VLmVoZ5duGX75a1HK2nqDfYTwWTXeB46AKFld8yji1xARKZICd
wj1kO17m7C8XXAM4tpa7cB1V+MV0QUf+RxUt3rFPhTe/sK68PDN+UaOVEcdt
6XWntnbNAntI0NkrRMgwJ8BUt++m4HAlLYT/fDlvt/uLkJcNPKbCRLWL8+hz
eCPHslQrLrKVSPMC8/p31hV0kAeCAePECRgZrozAYrj++koSc0Hw/4rIg2Qr
/v1cKvG+AXn0sx6WjaNqyGiH+wt0S2mDUHXX9lsySnn8TgHRWPh7YS3ipJMi
N8zf72yPXvgtARitIsXquEgO9e1cXXetHkztyvI+lwRZ5NWht8CoVJipwttg
FM+x/DNv81gJPFvw3KqpkArooSErvSGvkxprBAgOT1LnVpsul/q/VPSlfc6A
584WMBce4ueQWoP+4Iptt5gQpdaLvNJYuZNR7O8zD5z2JyA9PTzNHhwwZ6TV
+zWkFTDQ6rKUYrr0g62YQ/pgkYLCp6sM6dq2ocxSq0eSeRpufavfnkBupb+l
bGKbdSATkRrdzZ+g7RrUVLCuIDqL8yV78vnSYAnTRgpcJxe+nHH2KU24sL+9
P+/mgjkaLoWFh810ycBNxIw0HH8uhmSY2aH6B7Rt815dLt+JP4Iq+UYFo61d
CqnMvo4Og5og9Cb7h0QWTOxy5HUBlSJ+TJmfXozelyrg4FfOhghdvU/gsLS0
Bs/SpVMbUfdOjCS69eY5JSwUCqnIg5p8UH7tl6c+ehyrZLJEseOF2bRF6V+g
k/gtafJ4+XM0k0rA6ZB4dtzzWEK4n0k+TsPRJzYvy6mDYTjdo4m8hWtGl7G5
FdEXQYC9X+2PS1GmRJBTxOkXlP+VbKc1D/2FnZecDUH0nMtriTdK7/+azBwZ
CD56Frm8tt05ccVZSIOr7LQra14QsNlB8RAf1OR9ndP1qLsYrgJDc7YBZ0++
f084t2tIwVzxsfnSdX71It4Sbf7oIm0P458Iz0oUn3i7uyGjfmw+VS6T+7Sr
6du6o1YVywvzzGa366AEwPzH84fDYdtSVYNYixS5d8XQaG1HaX+aTXF9cR1a
woyusUXkuLqdgJGgpEJbkoeEsIZyMQ8P5iWXMFKjdWVARwF3UFf78dcrccc7
7ygcL+3LJak2gSShPsQmmXpcP5F46Ehn9lpFNkeqcnuQuMMu+7ju2iU5Wav+
AxLqTQmE8MoqtwIEUxjGY0Mg1HErHVhYH725AZ50PKscAR89KsuAeZdFbUrT
rapibc9FOEPFoEw7L4ijDlckTZCoWGo/7InnAI7yVxvhamlr96u9pvjoGUZg
/v9AM3MRI+5k0lKKTK8kN1U+ZY2889n7Ugugo2Pr/vnJ4OxKaFZUqjEog9yl
kIGSvfpc3caUnWDa+0Eebas2FiXOhEqbi13Rx7w9qcYnQ3HwBPlhTkfntx4u
UF6UU3i9ilVUWyifR0QGi6c2nyinXwdhA6jepfptQBMT/gH40O1yqmyr1PJe
jik9z5VeQYrHy5E6WEMdUYcq5vSLUoBe9mTWMvt8OaqPSiph6XX2bP0EwTep
hVsvtNKAdPEf6cgywLoKJ36k99LHfaESSA28fA6LDhF0wc4a6r+SvmaD+k7/
x2yt/mDa90BylauettHG5bzt/CVWqZzy4noocqPEpEn+Bpdjc+KEueYvjaFK
agERPaTP++sWv2bZncNe7uG9W5dfeOjWZlhBOozyKBttK1Zesv9PrBapWBCF
rM0v8RYkTDSIPol+NoCQ/ZQqUUUvRSGBRwUT+VVxEE2ZBPylxePfFBgq9oxl
MtxXSN+3GQ7WyMei6rzmboFts8e+FgHn+kHW0j3Ns1zEe7J1x7w4rn3Eyxjv
7adegxngWSteoVDF2wnkJ3qZSoBMnROwiY1R2VYy7zTvAgYiwB7ZQmjVwgOE
NEEtYjxncUAyn3ehCaaHQVJmjyuYdhHE1PhaQjoMT9zqOERgJhdnPwla7unb
1GgsuU9YyW0j/92B4qfWvFZBmEXaeMwwIbjqPt6NRjRg0+8GpXWcKgSJtGrY
xYaQcDfs7yw+loiV+n0kM4fdpE/3SkIoCa+xbWPUkBzxyt1hJXlnwDLy/zlJ
RefbmQcGNDT7JexsEBoS6NVBCBw9YmI1QjqhGxegFJl4RFDcFlE49BnpsuKa
pysy2GvvzR9H9MfKIto3jL8aEjNqrnHP5MLtUS7S9H8LyZyUFS3Db5WgEYuo
opCNoRjrxA1o1QxxN/lIO5HdzTf2/WA7oh83J662MyYTgHIyb7ftr/yNtLAK
9QXaYnLhCJaBbAXxwar8P1XBE481hlmIGc07ZYziMir2ABTonzq9pqRM+8gI
1XwWb56s8ox6Wpt29FGU41jwCUOsnuYZlTjjgjCqHhamMirEfo+9Lq9dWlAk
MyEw+/7sTilzTa5euTe0/4peiNpsSxkeavkcMyQUHtW2p8GN+XHB/+bcKL8E
FBvQpk8b/fNm//0rnfxjbdNX/jHkozfq/O0zb/FMwEhPpPL6w6hW1YG2SXvw
uCTZbKwWo8fiVafrJHUkg8hRscs2zFRACE/8TSMZ1PwW6WIaZO8obXk7+uQQ
MplJaR0MS5bxeTvhEyfMChrqdSzBgSPgNQJ0grJfVMW/ZP4OadYEko/iO7cs
31OHKkzpShDqpD1Yoeu/N4zDIqGaSpA+kzNtxqwt83qqfDNjSpM/xd8teWb/
5ZH7p8d/wKaWYHOvPcd7Q/l8waxKsrGi+T/EhhD83vqsc63GRpkGaphO/Ov2
ms7X9a4RPRBVcBMD1qTyVPOkJ1SmbmraX/ZWc3dCqJ7oHrxFkQcPhhfbl7QD
u6HSjF7wxMrnC1AalqcSuHpQYagyNCgIJQ/eR/UhGdnmR4QMjndIGGh5h7rS
kV4XJlFtTwz7s/v9+v0RNmELRwjzWhKNq/XvvcpVNUsl0oabOyqjlYJWbJEP
DqEK1xz05NuMFTq3rfI5uNGwGyeQbuDkZNOTqxpLCHSvCWv4aVO/3BM9aabS
7EVrE7NbxurW6nNyDFu69MrGCzdBXa7bj5FYdGO18hZo6jBcKXEEqH+IcIsH
3/ycdMDSW36kYiIZrmzL9BIGEz9yk9+fCJ4OygUC6vVQVdX5u29N470NPtER
36d5hTlaQ0IExUR+d5omFrMqoa1NXCXRt4LD/2zZ3KeqdI4cMl3e10TiUiEQ
AbPiZe1F89MkdBAAsj1KsXXFp4uHO9rW9xsswVXGY28bea4lWw4YdQ+E6qT+
NXnK8ykEAkUCfuNMaapUC/ditzj23hbUX0U/g4yn0pva5U/Luas+xXxv2vTz
KIkfoROmV4/DXV4Xbfz0XB6jtmUTxrP5zrlh+AWhrFHvvqaS6FGAtN5wzqy5
0Av0w4xoa/8a8AHIdCuSGXl6CsZeDKEA51dq2TyHHrzKaE/atd9eyoIE7QHa
MVY5BUA3xW9lcjS1ToHYoxdn2OGOW7fsKbIiCKPR3biZIaaM0jDM6S7Us0L4
KTIr0cItyUJMlmf1q7ETQf28AAbz/ihXyIfiRHthIBHwK3yEEWr3Bqs8IFG7
6eSMg0IXrkeflHLlMjD3f2z65F2YF0z/I4OAhMKVlcuAczudgcmY7Q9kjh05
45zSmbQlvymA2AqBiA4LAN/YwPby67EDK0tNCLaUH5FP4VpfD6nfjfJ5crWt
aB6j8rMPpk8AP2CYu3gca1OEi1zID7z45bKWJxeYhQMOgjc9lbY2m1/k7fiK
5kBhScwUyYMpT2XZddOmnBqrFoUXj4+SG/tuHyFk4uvPHUOmscKIzFDh8Bji
wOcWhKGox0TJeGatENyp07a/xI1FvjVF5TYn/AhX28MnoF9+xMwG1WNYsurz
9uNZJQ38ZQ1KC1yXduZytnC5TRbd3nPIn0Ws27UNrWfW4IcYRSElEA4xooCh
kBFGRSp+dP1p591CydgwDuyxsWaNDZnSoBL9EqEzM/IcQecqCp1GMPCgUUCY
xRYEP1YBYdpM8xRtHgtPDzEjVjtfq/760xaZ5c2VhWi2oDhD9gOvXPKdN33v
RvOJxx6qtTolTYqiywU0jra8075E5lxg/+zhR1W3JIgH5yyt8jwwQWydRc+b
+ITpos+TzSuyCuoXlU90Y4X2nBU06ED7z8Ua8oA55fSAlw80jzb+jnHZU0fI
JBue5tShJfJDCx8OTi9IaR753Tm/xqPZXopC5NOGXL0joqNujw8Jfj3krD7Q
5OkUVlpku8ApchuH/310+frZE1wfkti7FWJVVJ2ri2+UcA2b0IvjDYFvFHEA
GaAF+IIwSWZR69KkTQkSl6YNRtEK4jM6y33wQ4mfcPtzQSDlmJ9t8o8WVCrC
Ag6NSiPaiUAhf5eGbYqUugZ7MsytZDTN4HCZgG9ixJM9OH39be7WceEekxbi
3aLyVjUaEv9jSEzsqNKunAl4yh+3bBbbsUycDBj0jfCSlp9BD2Qdgjvs19wx
nV2g660q32wIAK/yeW9gU/Hbx6cmTwMczBFIbgZhsiVZjLJ/1SKVBm/M366o
GR3lAP7bokI7HHg0VbQTv7m6X8E8nAXSgPI3Ycb5pZj55qIMxyFnt92somS8
7yEDrWiFPB0hZKC1XHY3HWA0VUfcBsXt2BODdYXvAVSIxFDHU/7zvQoD33Wb
C2qtCmuJCF6QdVb3KM/4MK5Xq+FigyDAp7SgFY5Qoz3CXbgpzwnzCRUh3Sc3
YS2wyVp0KQ0f8MwtQF1WeNviYcqEYBLTlIuZ9j3OW5J9XtN/kwy8PlpQ68s7
aO39MN2bMSEK+BlgzlwixQKvCdK++mScG0C2NSgbsZftsjdsmS+tXTlPiff3
Fs+IkqIY7sEcj5QRfbMepSEwSaLG+JTWHGpXmaANDASyyfdMSCOAf+VV031F
7XGyiK967iER/t5BcsX3YbAxMcD9trbQq0f5ua57KIOkh8ZM87Rgk9FE3rSv
d/w7N8VkqaHnTleDAgYkvK2Ydqr32e6/mIkjDDz4SCqwbQ2jqNDrtCCQBWav
h0cry7sQ2XhG+RrilP8rxsigz0pYI+m/YXZbPMDl41vEE3cRVGdUyRGIUWVj
oqGMmAI7vrHwTx5FuDoyxIeVc3XiTmrOfVgH346Vqr4L2dZ7tPcx5vbVCzyI
wbBhUo/gko9jDtP+Aj6RiZSJm/jtu82r6EXkulBSXRAiifvPpN0mR90GLF4L
D18BNOwKp46X54YcwepWe4/USxtRrPG1cqd91kAhG9QCCRSKRRL4kYmVkqZc
7nwwk6Ccffp5chLM4JrMCgVUkEsV2y4IuOXocaRvBauoicgnyjHW2QMwzGZh
q2mxdRkMV+xhE6yKugNOrubH/SgAwrohfYyGdYD4Ijr/6H/XGSgHh35WGzgW
plAwbv6rAtWKeokuW466goZJqg/h7OgwAzbwL5tkpQb63kV7PyLptqb4bg08
ego4TVARI6p1Hp0l/PSUR9VGKK5W/O1yuBvOpY9OCOw1zHbfvKcTXHg3UMzp
AsJKi9SYoh95HCDVsGqBhVYqqzLfrO4UhR3S4/H0+xlLPH/fAfYldd+NDj0H
iCFd+dsDabTBJ+uhSQo87WqzStTB4dqQjaWBG6LeFl4kAbEtaWsNSlSvW8bD
kIrOEJ9OX+KiZVxbxmnEkddnxEZtf1vY/NYFJ88U1AwlkkYjHzsjPxJ4M8sk
b6ymd5p9/Ca9JFFNBYanuCmAH4t8dokWrQPCjZ3uoKw6jdP4vcqLcLInht1Y
KlLFYkO7Z2rFjC6IfZxy2fnC96lIrhu5l38LzigGTiBGum1tLdFaeReZGLVs
2hjT9va1NWWFQdUX+qWPKTgBPb6jtQzvXgIml6mYgMl4KOMHnxY+oHmWwRtx
B9ggv6DYLcCBOSTg4alcDw5xm/NShpYa5g4DSnwy/ej2tNGuTB9WbA149bL1
DBEv0C9t/tCtUvnKKs5phDpi/MYVMn0LCVE19hr5+VoHaykJsOy89kSbbsKs
l2BODLFEufYv8jxqc4ujlO3kRIRrQVSXlWtUWjF5DtvV3tvQbL70GupORNGN
Di4Q+BGwgCGLxXQ6DCDGBvroIsNLu1iZlWEpSHWpC5Im76ofix/m6ouKm9FH
tfS1x/GIn1BAJXSC9PbjyEgau6yN1ZNfQ5UYRCVjrgjq0uh9Sg/qBifTGOow
jqDOahw8pWv6+7Y8b3mFd7kabaMAfKfoy+/SDA93IWqVud5GvBq+58n197ms
wJ4j8tNqIbtmM7UBTlHAyVhErKciIN41ER7w4WUjOzMYOkT3uIuxPopb/4oh
dycj2zM87+p3TMsdPDrriZm/0jIJ6egQgwiS1wMiLYKSd2OGjz2zctwwif3K
MuSW1L2fIv4b/nDTz0+yMf++jvKoeFJB1DuPyALa/CDGie8v4Z4jnE2Bbqxh
nNfEv7DUhENwegLaYojxJ6rRoloTQBaDTemGyBvIcHkefsYEIjNMDIVpZpYU
n7y/Ncn8gvfbQHARoqCSlfwvtevsLf1neJt6mR2Kdb8BpqgS9l4Y9oYDbTgC
VyWUtuLER5nGguId8CmtbRn0slGNZ8BmV0m4Ahkqh+28Y1D3j3dmlzqfgyBQ
zpo20Ng3cnr9EXm+wPwVttbGABzD3QAL02AdqqIlHqbYD+c+w6nvvnmExdJo
NRpmuNZQY0WF4dO2xVPNffxsVHuGGbxmOboK+JsW6WC77bX568B60hshKfuD
4KlRBH+aSyxLbYzSAaxHs/WFbAU1SHebqYHZpKe64kxv3NKmoeQlWmUe3Nat
4fpZ9pFp25rShDE22gF8s/zsmZvTuSc3VJmNYclM+fRjTAqSgqHIUTMjl/ue
V8rAapb28Krt3gf906O+cZ/hgHUJrND6sCx1/Ab0rvP2BlV/4h7xgsrOCEjz
vXIOpx0rVwMSZ0qDSMWeyN1DBKOQko/QLG+MvmHy/MnG/ZqfBTUB3o4tvjYV
hsEYk5JwIxEZA+OS+xAG2oDTSw+tEnCRFcajwbOknFrWlZsQqk8PASHx8gIZ
69Z2AKeIlnzWvGZhLhk1xnLHmVQCZq73G40q9aFMXojpXRK8PjiEoDEJSAHP
PkdEEYcz2tlKRTlv9CyzTEk11JgasSH8v+SW5M8+ApnSM8vFFdzdiWz88mvt
bdH/rFbYwckXynw6ztpP37IOs8Y2HYy5U6GO6Iqsk5amAVt9ar9/zH8dB8hj
rRQa7yBCqAJXYmFtbbMSvQuTQtk6WpISJKoZQ3kGit3qGgN14hKOKHMtb+zZ
VM4suhsGklTIIGYLoXaZi1Ac2iU7n4xTld3DOG+Mf5P4n+JSjsCrIXOnfzey
vxoxeq4c6Xiqo8XdWMvSPJZep1MWVcF/LHKiJTg+T/R3ni373Zt/E2wWxgIN
tttW1NjKi252U5CQ3DDj+u24GcgFTG9JTUFgC2rx3SuUxtCGfKNUyFZEah3j
aFb7Tg/w2yEX60bxr40v2bU4eY3koL1VZow/rmQ7tOqPZXksQLnSlUOkV8jK
sPDkA0lhhSn8xOUBdjmTuffEfBfLvpjTXcs5DATNi+pRjK0dmuaC4xULYEWb
nbj+qp2BcAnZmEooiT1JYMyZ4nAw5XIGQ5A61x4Sc0/Ob/9noOs/f9Cx8P3q
87O0WBqrvijhm31v0m2gMvTtCzJu29kKKjQqRV+WubYI8raUGxLpiMHmVcld
wBXrnk4eDyainBImI+jYpelHq86YHQinmDbIcBBpPpQdpGa2RZ4me18evEP9
wqDJqtBMhzJXYjQL8Sz+xTroGAaljcaR8iE16+hnqw1FxD5u7qkV2kzuv2O7
yTPH71+DB84yP3zY9t6G/0Gn4vnJW+mkHMLsh49EMWqMjsEixoP+A8VH60g5
zeKlV3YrBsmgBGaDbQQQ971wkFERxvA3g4mVsVg+JWaXHLZwqZT0InGmIY7j
Fi9Jr4OC7fOAuSp4OaouuZUDcal6gfoDO2n3kZxqcA1sJ1XZuv6bQhNppeQw
Dp4jRICnLOz0NmtUhqnuOaCA4SU78Fe1GGCmgwMYFoW+Aq7DEvd3X/DIm8Lq
yqdpfabgxAU7bUyd8pLYZj1iig4LLkZhXLjat05TFOWDnsfmvy8CuGbMkXf0
5EfeVTEhdMsARoZvopgMGR1z+BMiQHn7jsI83psxEsnPJnTAfV5f9qNG02PB
2EEqKkh4hkcdoYZfy63NABtYUDgon/xdELEUCGz4/HarhVKEjEDJoz7LQKRL
QPWJfssdtcVNgzHmmoOQfVwfDeYyfK4ra5KoH2MNv34N/Yu2/VJdHaWDzLCV
XVt6lKgT+tYiDj6DhycaV74BK+EKQyD2yYxvCOiPXhADeAU3uCuN9DxNJY/l
gznrRmkNNk1B0lRoDQswakgC0zUKGEvnWxxRxKLQGgSl/TzgtMEkLdNqHyVS
g63Ee7d7ksxw09HQig/ROVzHxXdXcyJErKbUDDgLvYDdnpF5PaWR9RCYm+um
SIKJuEQThotbpuuXH4GwYZ9HsyKq0hyqtV/dGPQPUR0sz71EGSuXTgrBXuE/
8osJ5nCA5/Mg2DlXu4VtjsQJjF51W/c1q3iIQD3mlpST7pgE1uSu49yMmBns
Kwr1EXPuc7xWjphMbooiJkOv2lTizlih2LAjwW86W6KFNNEgexev8/CeYEK1
bHi2rew58WnP4mIZa83A2+z0OU4IuTIs0SMnyzgjJJ5BrJ24tCWr82sy8IO4
ctZPSXdEFGiC4KDAhEuj3+4k19CqfF5yFiGTky6yrwfd9ILEzkkwf4R+6aaM
RU/wc/aKKibri/FXNZ7fihpDFYXAnRfBqtcxzOqYGyfHTY46K+Il9u3BB6eM
xX0nfnLWDmOl2ME5D2GN014/2HjXZsJMGAraQgW733nvmigd9UK8f9ZjFozc
yXfwDf62qr9ilctompT9zgID61PmfV/YC98eEznQwxl+LGs+xh90C+OdzUxv
Vft8JoYF9tS7JgWsQeQYrLf8msHF5ntNTw5Sl2R+36I7nkdwZlExC1x+31GI
F+7pBd/lizuQYAkfEZLyQlsYrEEDmijcfUwze3AAF0+a0xsDeshVdnWrKO+d
uyjwaIcTWRZNwnqlhmD32+/sr8LBTI6OBfOBQz/WuipfCQ0bquBSbC+8beU5
uwrznLLnY4xFZrZkt6npDkTpxjb0rBgI8sJzXpng0lIYnd/Jq4KmbPE5m43K
HfWXLTWdhHP62hJmcZntwJiDJdWaku6FSgMw3BBWMWXcWAsFn+A+enNhSUpr
P+XpkgzhricRAmxiYhxL6JWObagMVSlG/IqERw2K05mQmGvqm3rc3HzKW5yv
WcNfH0r1YoKvaIyBmHdbQXUtjHXMSto4SAp8w8vJWUOB6hbI4eas5hwXMH27
3opI82cChmcgGKCuCQ0yjbsKUI5YZhs7OEAg+K3tZ5gWr36NSViampJYnR6w
iGOLkOIJWSZnL6S5RS5b0+RDrdIZQyWfZHhHkRUnZjwLvlLmUBQf/hl/HBlQ
JlSO0/3h0dPtcFV82xtPs9O2j0XRAAl2cyJGUR2CioOMY1ery8qwcAEpmbFQ
Vs+DEY+khQ6XnyhdZBBdaKO1S42bVY5Pya8wbr7dw/C/y6VdI2R29wmxMIgU
cnnvyI4RgrNqRt3B+mj0kiaG4TzYn4NVPj2G9JAg40PG53KwtCUY8G1bLzt6
oGUbbiAa+VibY+8ouPrVNQrPfigOffD+Z+4IfeUZ3weDdqAbDbKzGgJ8B3lf
l/lzdaMGrkZRt7pcTtTI05oePlSEHp8uUgbeTtrNQxC64qWK9N5uv1iAYZ8p
P7ccuG8nYgCc6lJuSD5+jOPaF84qCdDemVoM/rWPu7qIJwkRNmQpl7mGVXQN
5cK277tKj1gzceYFxBGFZ6dD5UVplP7KUJUdI1pOkU/Fk4aa2p/ztZOGx7wQ
v++7dcp10vGhdg2gKcp5gIGUQwTeEocc+7Mh4M0kQZNaxnjO6BJkZzx3LsZG
Xy6/0QSkKeZgK7gqWVmqjwFrFLghrhOCMYVol4rKQam0BCxx/eLt3asu6Vn8
b2H1qYG6+udOHfpCYR6KFy/Iq7ekW1RCygh/Wb+Jm3YwwA0kIrXhZPHdOzyW
BddojZtYA1sd5JL8obU4T2rnCwyWhISkyrD4KPZPQMYehAaJzz2Nkgc+FuPn
2J8W3vBcVSc1tLsY4TLrPV8qgApQ/s+gPb0cevs3rLERLKyTe2Gc367XFn0+
/bPIQ5OblZbKaTHP+Suo0+YbgBslFo0lrUDJZNtUBm/uWdrUnR4nB5VCppjN
zR18Yd9gzowII0dLddm62TQmDAlGU+Kckkld8qmwhYhYBvJmpkCbukD5pfRW
JMHl+Y7zxiw7CIh9Qj59cKkvZ8+r+mrDPEDEFRIQnHkGtZWH/iausv9ijLp2
7gfL4EkXZbnvdrKrtw1p0+AvZK4l78ZomX1S9hnmYuX/c7ZONffLKIz6uqO/
D8u9P3SAky275dV9zkXUfOdPdk9X7WYK/I3VxhGsmFj1QlEflnbGEZKe10+f
jIpQ/3ov0L3ip6YAPvYOqw/toSblUf9ZLDJ3gHi0APQxYiXH73afNM2LjGOU
QU3a2qxVoAMsmHAkjgN0sMq6i8U/X8yKAs46FIm2TG8i4j+7iCI93R8QO+XK
n7JsVxNgtrN3GSkFTykJwW8a1SRnn9/fBAmWWIvjxGquF+hhzF6hWLT1bB8l
bdt3kswxl8CySn8OzDOBysdujcv2HydS5YUAbYVGko+kXU73v4abcea3CvtW
6MAXBuqLySE0uE3RwHCxIpJn4rKNquiWRfpb054tg1bM37Sddqlqb4FYP/1g
YxU8Get2u2smZ1X7jhmjjuJz74ejrPo/evX7Zvb7pzg7y3JCAfdUHwyW1N7i
uB8iotPoBAMmPYkM3v6tCWg/oYq/5jfQafCBUmQxiz2ziPp7ISs3L/7W7cDZ
N/5KV37IrW7Gjn5LZOLulVGPIDnQ9MUcArkpdzBRCQlquwOaOvduhkyhdckK
dVJD1r86T5kL6y5df3KhnTJQ+5xF3mlBjYGeqf1IIphHJLYbBDiCZpVpmtRk
NtrlxIR8UB7Etf+2eNjtRcFE5VHlctnDkFrhUpyrL3hwit35tUKXar4YZK6x
k0ffXzusZ0/7majRZOMm9J4jdewady2/CyJb59LM+ttWkZd3VDvOIM1T4FNV
O1sWUJNcRkxqWVCN6Izku55Ct/fU0oVXaiSgVWv4JvQNgbMgruNO1Y5xO4Hl
rxceTrUofhUm+SZBwGxfF6sFscJpEsKsNLrjaX4eUwOTQuNPItRXA08/RYVs
XFZNl+hubgLo3PBrKEgLs9o+gOCnoYiiv0rSdDE0aHIovVvStrH6UV9Da1vk
iNR2bNY16otWpDH3yAxlnc1m+247RZ9mf9il5FSlxOI65wfeg/1esx3fge6E
/6AZh6O0FVV+mkRQxo5mTBu8lZ+EiWCcp6jvkNBZQ04Ru51dDAUo2PPZc7VT
o2PvhxGDYau5bfhgWC9W12T9DzgAs4jeQzpAhhm9jJx1AF6680TxKUdSMkcq
G8YidiM4xvwzLfroYiF+e986RSBFqwqZ+ZJdwsUdq2w7RkjlJ8+iIvfYu4bP
jc33ocn8BQQm3ymWHJZey5bcDhAbF9zF07CUTOQWjqcf1zo8ZwJo5Dp5z974
+RmQPKdgd3wTbudoN7qDZpk+DNlBAMvdFNWHianr2RT2EECwZ7GVFNynJGLo
aPJ/L/vMw0Ij3u+korJ5u538pnBjp6l7x274+p9XTxOe0AvJ43Hke10WkHoM
xzEPcd2y6GxADQoELiYP0HoUl6xCrubDirDcHPKvuN37lGvPvCwgqR2gWYJR
e/CZBSsA42FxnUphQtHS1y3uBJ51yY6MuB+CkKU+GeY/cPGJe4XD16tKfdyx
odIBa5HAE051Hd8tjNf83c33FFc9n3mE4AIAFC6ewtfqAzsUFE82MWBctjmG
F7Rx30RndFn+2VhNScQTavipCT6sqinWfzzQLODNZuboqjkc/egbQyomyAJo
yTaaXzz0wXeaNL06F2i3THkvcr9c1z63whB/V1zCXSp8c9gVBHUSd0vtkxop
/Sq/BFiaWA0viZFQRNtU4V4+doUUokcrzbCKxMjbxzIHMkgkkrIlOqlhV4HB
apNth6BEL5k4+k7Wv8iURKMIX7e9Q4tpFFngbZCuIXIceHTePL5RjA9qcxfq
q6KqGOqqFXNowZDPlkpMOtxj6NCi0zU3Hq8Xmx0efRjglcXC0DWg+o7JXoAF
yWZbqIPF2spRmxBc2IxcRg8zG1IV0hvXHHyqrsI8nLCsohImFDKfyZF9Gyjb
9vdwQyrdfRWL6O7IQjLIfFBibse7cMWq1LZPd3xTMEW2DU4Z67Hoy2Cnfb+t
ZaU6Wjb5XpQjL6i+tVlv7NUcQK64CG8eiykuseMaWVxGdjAItRBXlDbQdB9w
nyTSowu4OD0IGnw6rgvB5OKMonalI0dBokD5WIUybIk/Pj+AW0Al3OER0LHd
EFKgZ228zg39s0ODRloZNR+8c62OCvQXdoZOdedNcxxypLYxbz78ceeqcMle
5NCsjSTTrX5CTXbADuk4bRLQgf4xTj6f1UBhOBsnwSuzrSSAVEIhXa0JzlwA
FE6Zepzugjir427AdkMi/Hicv9KDLCpwN6Pnizbm9CmDCoq4YMXiAOhhYBmc
594J94V7AXKSSvo3u8mBCXpKoOOTQacVRQ68l2PQNMS81jRkG47yOuItvzDr
t7EDQO5JbkvY6FXUO/mcne+F5N3qUrCP+WWCv5o/QTP1f4amikWvfV3bDzox
CvR/ejQ4WZ7ZZah/Dk5t5iyrM52Sur5ueuVDAZ845H+paNVAAingaLPcarV7
jB2B2HnTwCvOP+WmAg7jcgzrA9V2dVZLOIqzS3iqrcUryPX0CDUceR6ZTA5a
hgLzyL4FenNDcwLDmVYH19wCdZkEGbG7HqNN5jukKkItSJXGVD/I1NiHE8xl
3QICZaGJ0lVI1baHG1rlQvsVHUKT+TqKsc1aB8sLdb1lVdflIkXSITpJwGgC
F0dYqbacffh2Y2GbwQmU/IaYmn5pHQ8joKxBJhKt4Q3gmiwA6mxOv/V15IZO
nE7i3BD+rOn6mp9YcrA/lU3KWzw5IU1NIYk3DSzEO5KSThgwfsmIDmEeNDou
JEx+G1BsIff4A0d+S8w4ELY8IB3Q098WlsI6AD4vSYiNdbI5L8+SzExs01nO
kCx8EFrKAzjaoqyjLEHx8INkgHaPXuPb0guxkQrlFk3vDoBQ10p+Iwji6l7s
772oDHBFjOJ08MFg3Eqj3qO0I8Xc+dcxdXprSXXWUL+9fIdRTPeF40a5DcEu
5bmdY8jPGm+Rq5IDL4H2GJaqmXXa6+3QZBIbOfmWAKGIuFQt5GDT9zM2qcYm
v+z/gDclreG+g3H2iAi8hhjNMTBlLLdYnHERi64cD3nEY1qIrLvibJoRgjTu
nV8wmxet9WOgWbgX12sGjVhH8vBS0Gy5GramO7y61tWDc+dMBDgYmuasIY2l
Am1aqPAxHKFCVwfm+yKu6ntl/iyxLfkn1SLiICwsdJjwii6Oc1f/CgFExjLF
iKLtajzB8CFd2/Dvt1LUJVvj0VFY2cQU8F4hkJ7uvCgl7UgOVduWMSgk9fZt
5yPIMDPo+JGPm1jzhcaikPFhkmP72L6Ng7EWp7qBheqPbPfQhg/KregePors
ywaVIuf538bHurpwfjUcfzRGY53eBFMODn1e/7y4fCK6oRZEZSciJU57nkpb
aHa+c+GmHur6ozdJE96vZkNTsvRKYPUdqQzXNT0M2YeLFso7Ux8bgwWVHvZ5
r1mR56pyss77mYz7PMCBYi/kLs6XBOxhtpRj2hPsDzalNSowlXj/y1W/AJ5Q
RDv20E/AgqAmW8eBKokKyFyu37cJojJJqACRvlOkWZREggHEQWhs+NfkMQtm
QdLg/2iAYsNbbMMyBUulABhCqom1fBAav4UlZSkCyxT371pqxs4RxjqJewj5
SIaYzsj0RRMp4UMzMw7JjWOdEdmu6jLCWbhoXpdTgYmGCogDqHC2QuZdZ9Mk
bFrAQElqH/l18IUaITxewvikNEbl6vYBjBBE2lvOWHY2luH5YFkhs/JvtSLu
eTp4UvuzfkCh42+9Vuiq/jxZIClSINrQCqYdxoajdXpbYkpgsNvzIVTOp+EK
BOoKP8yjXGIAKRJqI7WRoB7g455y3NwDwBkx33gwp7B+mShhF5AvKqkHqJon
2TgAg/rcQEbaKSlSmeYxRtDff3eeCOXfYP604RsDF/IGxlO4dgi9kU3SaP2Y
X+o9/n8FzQ2j73975afDXVSlPQRiLEjqoR26Zbjmv7xjh/mqdNLPkgNWJJ71
hN3GYcW0dj8d0Upy665OQo1tDVwQFX2NSwbjlX5OrXDZdFdNn7WZUs9zhzU4
ac4GwwAEZatwx3SV4Iyq/FPRv4HREupenc71ptW2KV0neihWlnFB6IPx/hlC
FukjfR00LB4fBsg/M7S7mLlfr3OvrwoCaM1HWcvl2QOUPZRvNaE2P+0IvS65
jbkGIEqzRXu1HVg7L2i9uemVaSd51ac8ZLfXUuFj/3JV2dq7pbV4A1kxniuj
TDgR8uBnpFZXZnF8dbp1s0QGDjf/w9DxqjLBXbP9Yj6J6i2rbqMWB+O/G1bB
Uz2tHNFLyQFgZNyBAi9LNZYVkcF6UHuTuFGZgzdvZOYgEd72NnD/aZs+cmSh
jT0KzrjjIp2bphRek1hhp0lAG1p5Yp5+JiqqXv3k6S2hRBOe7DS/hjm7v5FE
A+VmpSaC8OXLFI8viBC+VwtPQ4alOcv4f1D+t7H1adPTkJsfOGlKOeDey/fm
+hzqssD10FCzgaRqCjFR32LDT1FxKc46SgXrzRJGqAG+dXdq9GKZgRZ3UonN
fN+4pam4JDJoW8Afr7lqitSAdomlq17z6Q7Qq7FtioLl2geZzLLu0Klo0W0t
tpnU81sBPKaftjd+bAt5JEHZpT0BJSBdVTfeImX+T5UuTndLW+3QMQOxSJp4
Uy2RpYcN10hDaSXllCal3vFkBYMGN3MgFgMli4aoarV0kXuqE6UHV8co6OG9
P/tLAO3zX0gBL/9m+9lBSmUAmkX6HAIbJSukYwotT3q6P4s9YIt73a38u6Sc
YtC/xCaUhi3jdOY3N2pUyvRuknu65HYvgpvYwTAqJweF1LAu82O5ZgPDifQg
uNpTSroUn5xwUFPmCxTfkfmoICgY8TTx04c831k/OSdPAryMCG6ICehGmEzO
dYTgZlMGjiWqPw1Vvk59jVGW0yjuSN34FQqFkrP9amFBaPVZ+9PUmQ1vi1oh
H4lOngPrAsGaXMif0MvqzSS2pE7v9+wMQNhqR5EAJz/1yg+nlRtj9vxSp8l/
PdGSLnfSC8XL3V8AcqNXz5k34WOKEE4whQFMFLLyQwh4rOzovH6OYhTV5Cuq
sP7Js3uOwCfWLfQ1UIFjw+LmftEYpuRkwcx4dXcZfVj+Ld23IQ/X4Uu15sRQ
2tcdDE8tTtGOuIXpzvkX3wg8U2OeW+dPvnmTq8I5xOD4V8PiksaTFGk6sjjo
Tgbvk2kjB1BGgBxUGcsATUvg/Cl30YzxHfe9mMp72V8DqlbhuOoxNBbdB/3U
2Ha/of9sB07gy/ESYUqgm0tNridRNwO8bGAklPZGTFqdAO0vxOX4UukKe+TT
LVOpI7uxB5yFzj+SrXTAB0J83dXZPGxsUdbBx2Olfx9WtIv6Px5QHgBU1lPw
j9IRSyBiGPAxDIIKzft0HlckSmr7NGNGYFD2Z953cG0oeidVEIjlX7zdaO5y
eFIaNZidBbWASBc/Tcy2vmlsvV8ZL1gPnUzu53NsyJT8voDl6GaIBUM3ea84
vxsM7mCB/FCxHLwLyuf6yjwOVkrWzqafX/ihLguWZs1zlNGyqCckRBawKzIt
8znEBcM133f86biPhr6nmmK1NDv3fMeQmTCqdP85EXu1k2gNykBjKH9Me2qE
q2HlObIkW3pbLIquu42G4BV2CdL0kr+Ns38Oa16awlPOJ+Q9SQV0TAJXDEp4
eAUvkYwrFxOq8hrtMxXoMF2MLUGPIoyYJ0zFepLaqIsb7ugYWVBr8gc1jBdi
+oeX+Mw3OoXpmUTYRcOlHcy9n/ldLMqw/jBa5HWjVLTj9QXS1bx8cApLxxnw
mRE3hW6Qq+MgjMqG37fMxUM0kSISp9CATqV0Rmm8pzf89rCbPCLAAVFC0V55
OGpy2ojhp3xJ8tsj5/QArHk/0FRLuADPYReVCkNAj5iIiNSsZhUpo6jC2nlV
NzmoOL/4WxEARBaf/HdRMeGSBixyOUrtZQP3zdJ6Bd47d4XV070/o8CA7YH0
AHMKkelsEHmpy34R7vCabCMoQ3ZExPvOqZ4uzf7PePZ2kV9M46l8R+HDFu7E
KAkz6X4hj+VaG5xaypMkcPN4bL+oOuU23DRKzHD2HWWDqUhNjs71XLomS4+s
mRir0VQuWGdQqNWamDWtwo12Ak4P7bChdMRCHTWIhoAxh51TQGI2dppC1VXN
RIdjusisiXYTugtICkz0HDwP0rrLuZkR0Fw/7UaOPsWyjJe3Q08xoAFTT8Xv
wAqGn0DoP5+bL65FwGHvCe6YBen93oBhR4oXZkeUM1DLnXtX1VXBJ/LG+KIi
sk4o2N2EjyKeFxNC8hdXOKUTOIrt2vk/fHaV2c1s2cyqxh6wtWU0+Gm5Zmpr
3pzmjwLixB0gp4KHCPCiee9GS5kQBLysGPbp3N+T2vC8H+P52eo6AGWHNXwU
oWpgd5FfscH9CXzfM7/Ja4woYLaGnVHwWUSH/2Bs8llTrS3bVuBmg3Z0bt2W
xJQ7mccale21CrvD6H7PfW/51FLmu+jHnLN+OJAUm/zWvGY5Tka17OC07guD
gLWCEeUTtkDeJhkRA4ZgnutpiaZrMAGV/vajzKwbY04bWU04Lyqf56C7ox7T
Ovai6uoYjlSL7ddvcVZ1g4eOUbt0asGotS/houzikUAi5qi/SNQAxC7OrNdo
RjdIAT4SRCuCkloopVN/uHKLRn3Ffsjc3kJsM3e8miby7SIrinayVPcNvXGv
nVMGJwI6VShq7/mZ6/sqgEB1sGsn5r0Q830Hdo4SOkZR0NoZq8sxnciyXjyu
XgzkMcwEh7Y0BfP9rBKgsDfdBz8rmFGk2Iw59Tur+YV4MFy281UAP5NC6Y61
tnQSsJ+j07hPLyPCt3nXZcUHrXgkn84bYgTYBFE2meAhrgemZTwE6DaqtkUL
6oCXWnM0/YXr43mUN4sFgnyfOooHGmU/wgepfSqB4JJQc6o+FtTJ8L4mIq9b
HbhTUOJaQNgG9yiBNWP3aur5UopVCjVLyZbY0vHGeSFiEU4tnQGa4zteeHqu
ig6jN/0rDpzrrqjAp9+wJootlZoQdfmubpOxUtmGcOYVwWqcwKF9uPVFeVQV
aj8xMD2nV8XmVd2z6xBdBDOfdB2usUj1QP1lRSJRhBPv4XKTCvBQO7GeWKEt
HOwKCZ7C6BKu5GiHwA7Pe7luZ4DYULDR4YICEXr0au3iH4Dft8l23ueyUuc8
8FqoMJXpF5zea3W+6fukHBL1+E/yUqA+xMhBPKoa7fpKYOSB2x70X0vV9DVQ
D4foe9NOdpUEgcg86IW589xsxXNFTLdZwt0770ICr6PMN70eOxNlrbTa+uQY
q/vc7aVyktToQ3jfKOCRqr/ZJFmSwPywd6o0A1Qf3O0bRKLPUEYxLDRDS7X/
+m5vczIU59SgduSfBHJ5vbjsM6PDPHZ3qw1jquOuq/H7XpMHW7enSm/b9CEo
yoKlbxc3LHPpDRa7Q761GayUwyjOhgsE+Wpti0qcsMy0bg0H0gbphybs4YFc
qzfde2A7vR61V0LZCTIyihFk8bhYpr2TWjDiVEKpQ6AdhhGZA0Zmv/wxnveE
F3mjNZlJEZx8t0mzF3cS7n76XqcXvIWCMjXFtwWoKtsuDuQeKLdYC2Lom7uM
svB4tkLjGptdoWA6ROC7ESt63DO67hoFh+qRhjNX5yEuI8G3HsGsX4Q6kfHZ
OKfMJZL0wq0DMki7w8fsG5pdGTY6W9PsMf3NWJyrE83tKWb1TYgI5PkKnmf2
rTKiXyvyyGdORGpCKuCEXNglCyVePRfFo5DILIxl0VFdWVdZUFmZbkWDWJGt
MesJOWAb4okTskExdDX8FKdmeGp9aRInsDBF1KyLREv84budrr3Duuy0Acvt
lSDpjoMNAdbqoFPYzHhnGarnEoP+d0rREbgwVe2KXQuMkteqETuy9SCAz8S1
m2AB+XT97kCiJnavox3Ws6bqJgZJ7kUfIxANgEr0z5pCsUQav7FlBFUYCGW5
EzfaVxiz0ec2zpX3JcGh6ofbJXxDWXD/W6R5YAHg1vnQcxKM5sVJbRwFoBRQ
+0ItqK8q+eDtx7QeBT+xOkp/WBMagXG1w6JVB73qyCXNNV4+85d/aMGTC6Gt
QrxLEZID4N4DgFm3p2jnsxDcGQR0dt4P2ZQUt/1wHKntSLhJmCcf0ASs6bWx
cLV4FTTLMf3o1CjskEoirBDcrjBFfAj/EM4Hm50gsFCjXUDNDlneE1A/OFuy
1LanU5ok6L1NmcLTDRH50BhljqgNEpjA7rKbhYHl73GXUvGOl3uX/9sTo2D2
mbUXahYj4MMR1UwuEXN+AqsqTTp4s/I94bO7Bj9u4Zi9Wnww4LUiEAftSrlU
QAc1F7dx/ll1n39T7B1y/Cpb37dphijjkUXxTi94ldw4YdwNLvzvpgzWa45V
rcViPj0tWSur1jW6/YsqA58s32Fnd+oNuiszXCRUmaoRvU9gGFZfu8XXmK4L
SMLqn0RgK4d42W9ImTJy6mBkKlTjGWYUrOjTe1Hhu+VYboDzCO1P9d0YFQMw
B+2ukRJZhkv/pPcpfVlgTkVwN00zUvbW1FDAAYNLY+9crk2l38SzghWb0g5G
Vk1vF07ZawL6tyo1+46Fp8w8HCmdSfKytXd47P3RVjvMH/lsi56GDRa3Alqy
mU68WQ3icswy+DAfEcMaDUzow+KpIQbjXKsuKbo/IGjIFoq8bHPY4BM9QkdV
ZwAZQ5szIQus4bv5jF9oBD94s7DlRY1L4noGA/ElSYqwcrZd9GadDQ2V/2Ey
dJ4XB6Yka4Q8fUuroqwoXlxUn/gn0BFcVfjrnZCqbwpnm3iDyYPM1F8PqLZ/
mpy/SIT0XH/dHEHx6gP9gm27ZZPi67BGuM3DH3fzXX26jzSdJfGdvO1Ctbma
6Q2Hx+aehoBB23ZcVx0XjlGC1tywo4f2BPBHAWSpSGDKWUlvsalkbeNw9p+z
tACR12KiY4CFyRtwPIuwAEFxF8dmtV1rRu2spCqXXC4tnEN6aVYjEyFF0dCH
/Nq7hbhvut7AwsxUi/H8DMgmvyI6ufRO+EijCPCBzzracw/A3+7w685iYF2o
eqSXsN+XEGUaiBb1ifTmNJ9rXQAhGEQKTqkH7j/x2ET7dYSiTxsOY9gPjqSL
wIv9FxhU9LJDVSqLmW802jEOc5t1IYhzNkpaByJOxw+dcFbpLRslPdVFg2/p
I/9Nhn2gnqTRWLfwHYnoTJDNCX48oRFK+QrTRf+1vKyGzUJmuMyk29qZrGUA
vDie4aUpQF/1gAGiQ3SAZR+2d/O4uUb3StiqqhapSj72ow6E0JcD+QYddvfZ
PAO5dx90R81lcELUHeHAqSsMV1BaXvyomWjHRl1Dmwye/5Curtnk2VOZ5WHz
/hZyFjixF+9gZj9YNK7Izn+qBMlyYsmaxAg4NXDoVQgSsdvJhi8WTpESNent
QmFw1+VmZtT9FNrXSLyGugOcIprpj4Lienw/tnP5BxbZH3aQsax5USEtiD1c
ha/L/C9fm1wG9+T3CZJfcZ/e32559eG6bg8x0wg//F5xbdTKw7wJd5GsiUxI
s7gE+Tm50tJRiC40S1r0IpVgSH6OFWmev2moVx8aJwfkruFdSY3Q+MJQMQ8a
VL2/l0Il+olV47qsCSbfMzUMt9I+EbSXTjLepqUZcCOagAnngndCQqrHtdVY
7LE1HOTu5nbGw/NG7rQDqiYMfUZyCKLMFh5LignVvBrlhtlaeU5Cl3+tDajG
gCKLHS6bBKXaI/sN3T3VRyCv31p15Mj12NG6pHVE98cvOXL6mjjsNUzGkCUp
3f5bsssGnAjq1s8nyNNE5LAmTlPN6ahZY9Sa3bTDUf0ep1m/FmTDvPaPSbNc
iqWcQESwbYICW2QtSLUNhtkO/p9eRj1hO14wHfHvlF9XNdYRuk6zuKwOWWmC
8A+B3zqAEfCzh4q+H3sP7fjPoebqY1GQPZqDPkcn7OvltK701lccetX3SgGi
Toxg/G966ScWKjr7M+oAED1n1iXDtgsnRp0nA61VlL6BQ6WIVoPhIwvH9yvQ
HEBcVF/MrhaOODyr4yA7dDhHQa9hQLCWl6EeSSH6wtf3jzclBTSUAShO8KvG
nfB0W7rPwo778AQxQ0l6ZO+RFiWPI5TlmzPEYCJvN/Es3d38rXsLol4zIe7t
ThDOGF+XQxEfFvBjI9XM9LAX374GboaJrGMUli5wPHTwuE+exhSE53Ba127Q
qDlJNrbpD74Au5Xu/Q24lkQRFw5qxS+4d4Gb8x5rZ0Ejp55JRfMx1X4Fjl4r
9CRle3PF/ollUK5XpznlmoHq50BIZ7TnqGY+oF9/ekpXDHCwj75tXz5Gs/lw
isbdjSLyMjjZVlZnidqVBG4OzKISoXjlzh5w3rWg1jooZFia2Ci0rs81WSCA
8ixpAMLhvMyzA0zEAe1sicgG4DJ9ZH4tHqBrtmMcnyejMC+meL9IYoPYZH1+
hr5l9d2JyvV+wDaHR0iZdIUb1v7W3jZCUgPCa8GtRf97Z87Rk7gMwuAYMLGC
QBSb9+8V1Wx59YHwqTHhApd9AuXB5ZeFY1DNtXicVJcyv9wdVuNQwcDN4qi3
gHhD8hleJCLAjB49J8BSGBVawVq67wv3gVcrMYBXZfKbUqNsdx8CwuWdDsu/
5vkXr/nPHRUUqLxikTY5XHo9Nm4mjs03OkKjzzvZEyk4NT/8GNMjLGpIQTaq
0rfFFcMkKivQDabySxE+zZfc3xuKjzok55Pjh2mSZXv/zdf1vUqNr36r6xTw
8r1ThICy4LaAw9GrbRPGWxgqYav0r37SrP4kCgoL+L9qWN6Vgw3mRuHdfrrZ
QBrUc+ObJv98NFluBnM1QbyNMwHOuFxiQawNvGzV2faMYRK7GtQzCueLvlQZ
0dZYScr7MGgALiLyuhlp4LMbA0lB+8q1H+OH7HeaN6RtbmV/XYIqx+cnQ6xy
xctOJq00yn/mxtNRfmslcWh3UPI4Gf/5eg/xRcfWxuZCa/+vzIqcSL3Elg+5
bXw/Co5Ehr2GZEBTkfFRHhvp2GoDfEvTiNLxL2vRBE+Ay7HBUrBx3hudGP77
/poffzJVQMg6xopYhEfVnpg7FJkG36EhV5QbJSUtnaN3XHbS5q3ibYUxm/5s
Z1ViDX+CGR6/qSgWd0OfSa8qMDccj8Qhh8FbqxKdQqEbIux+2Frw/WL4cTLg
ftPdUmsr9OOtUiXW3b4mqnaEt8vacthRR4ryrnVrPiYg1pdNLfnkvN6ISajR
rDppHpowljHAvYDMHwSik7fvw3Hv72f59NKXwlG2C4C/au8Uw7zIuYNcOOql
Da3+oPVazcT8hMsYglAy2NM0zJbsvfSWiGcuhuQ/L/+3Dee++FqTO4RldhDL
Jf1kdhKb/62jc2Me7Nh4oSROgKhjMtnFEUPqpTiQwp3MmbN44nieLYZRKGdZ
kkPHenkUGwloNiyHWyGmyhdmEg9G6jU0Bth975d0H30G+BubKxsGwWEHssmr
r8Rp9Jm3Ptvmo9c2ko4IkL84cLkLN6ivDnqEB27zDe/Acbb4Qpg7EJUVWQHH
PH4bGgtM52uofXNEnTnK8Lv927LFIi8/Q5LYbQUpQex7OMMUa+D1LOFjrbuM
U01HjzSinftUZu8H1YP6mX3TfaF5V+MHIkeSEggRXXf7/H5M4oP8wCsqf+WS
KF6IsJN1QRXDdnbAmhOIAgSj5STM/VgUHXy3oPVqixtVTgJ/UBhcArqmycoV
dANW+MmznR8Neip3Z4ee8ZLL8/SrSiaK8JDTQ/oKsEkl063pzUa11/l5pOCm
WV3rchnizcaobtJD/s78ai61GjgDrhcNx3G9UuAn9nODzxIZ7lf7Mzzxljr/
2C/s8ZG1MTNfm+L1NWUcoI4X2oj9el9G6VsoriplqIU0tGQEfmslLLyjMGzG
uhGRV7i83HMS1YPXORoQoFQf7AfSzxrDfBbdW6ILWTIyejeyXs4W8uSnK83K
CeoaeibyTieYBV+TEkL8jRR1plIsDixVjcaLGOrrCGiYvzQLsCtHg3ntqKKF
0mokXkv226sL9FEtLRNSN0bwnXs4SRBd2DtaZXAW5Vw61HZObVNqlMtUgSI+
I9RPeQZNS4bYu+KGefhMsNgMRI+xXwuFePT1gqLEnNVZas7hsx26qdFbxxsp
21lwKXgCTGhn3q56qPd/kV0sw80Np21EozWQYMjljBehff5amHyx/iLML1w1
+3bC9lKF74gzBj2l26bLxnwvFwYhZpaLe+V6TV1DvcfIYvquBd0xCU72EbRH
cROK5JohJap0as1NrfY+KbCU4SxcsiEGSiqu6eTNfH7dyJ5rd14JR0a5N2Mu
qumzQ0uscK/hVVHPmLSLnyzkDK11NgbsCzJjpYTrg49plFxCFkp+C9s7Brsd
2RWtcy7diHMVszit3FNKjlIuVbH7MYyfg5TdIpyNNnPaE4E2i7Dk6iqPmqWm
QEhf2vwlHrXWk8D3JtwkGf7XchuLydhBWOOBEq2ZSAlC3JwIjfdSJT6Btxaa
KHY/LNcA8uyK2z+HJYZDO/rgbLmP5kzryNEmcECHF7Dwl/lJsSi+yGcVw8VF
uO4p523E1rfm335TArisiCgPWMxmvqi89eo7+UWDNoHbgQYmswwG3/iZ+H49
jLiqVyV5d0bBTkMT5QU46yrmxRxZmq2FOxzIwh2oRf+RALRl3cjFUlOb83O3
sVlv85pwOQmpIOO4oD62jWTNsIn1Rr4Cj/cryOy4oF5dUlRakzzrrXAmRFgK
WxG/Oo7SLCbxyB6BD0izkNnf4fs++wMzgNF4J3195MjX1hSFdWDVIsozj4xV
AurFwkU3YlnA9k4LEsnGwypmZK2X7uaXwpxBow/Ij3EfyR80um4RD7/KdoxE
IfPMwfOUFcyo/w4f8LZCJSOjEfbxpwNUh+ryS4g2+3zYsAXnZL3OchkzVwZr
T5NV8Gjfp7bJgDId6J7JzeS2y2hur9iNixU3U5akQb037uva3fDMHGnI0qzl
X0LDAIORy2YPU4em2KLSMYtSsuFmp//jme6L7NsQBmtFOHnaFsaPZTScoWVr
+oYGpfT7Y2Zcl3r9R4RpLgI2rvnqigPOe8hb3jP7HrdUD/JxrBnwMI9ZSBKf
M1vIzUf2KW8yTYuBWBa1g06SdCM53CzgIE6jyj3oGycHywjCr/f/lnYRYpaO
QKfAVNFmypuII/QVVFe0+y0lvZAZ229Uz0wMvzzG32MNmSP6jiuHQ0Dz5ieD
XfQ1pKnn2Fu6u0rIuriWYCMrVX4wAWdsMVhsHcuNgTTS5tGi0rtEMrNo0Y+c
VX4djKFCUchFEpWBVbf6DNK6uLi+m9jBifxHCIZekznbCHp6uCesOSS20SGT
2QtSXuq6eFkqt9P4Dp3kmVu029+3CjXJqI0AbmFa/cRFXfCBaW772Q1mLtma
4X3Eiwu/5BQdQnNn9uMiNnC+XknEW64v+LXK/6EbDO+IqVoVeXKgbZ/OKZbK
wAayBso8CZdQYWX8vOkRmIwcm1IxmvQPwshXAyDXZsw4RfwRQ2CaJv9cvu0q
OyYYVYXofC2R7Kp+QA1Ntb1dX/FJgJmMq43vHO/BSQy3EskvRCU2x1a+xX6q
FSwroFzgFp2Mv2tcb7Rq5U7HR90+cBYLppd1YPCklZsg/9Q/84teqcWIvGIk
GqH7C1sjW+D5ztoTCEnrOmPrfo2AGmwBd4GrVxae6Ct0CccYpbCN8kP6d3Sp
zVQjvCDR5Zm6LCL4ZeewMjPzEOsL0Znl8FcyeAqi84DQrBmWQ/SXNewFFQmS
bLKfJzsok7ZhzxuVV3MZDEobNTUC9smuKqdcjgYU65MPqWyZXyso1drpL6KO
Eq+mXEdarQ/vbML69SO4EAe4MP2ckp/+R944cDgIsDluS5OvGHpY2ekrX+rH
YV6uaUCcEuAXgQBf+4r45ZhDC8nS6SNShaLCd0JgsKSc6mKHhDgAyCipT/C3
hzVtAKuG68GiLL4vt8JXkGgV1MLSlcWHnvFVoaqx1SjbNxLgwWL6lPfMBIgy
OJLP8VxsfE/Ix9IgxnOOGLXCq9zbKO4OrCzcKl2FiWeUWcfMX9OTZqRrNzki
Z6U1FUAPds8Jg16aqmhCvwYZRumxtd/jmT9xO8UHh/xFKhw48j0PB8pCz4rM
+JgzFnZWsF+GdglD6WCSXJBHqR6TmdrkVdougUu1PwuzeGUxWWTRzxmn6MST
qdQWOPn0q4X81gKXkCxoaMxHFZ6udouLMqyZxBlYgp8UqmAYY+k/8VjAVxxU
oxVycuSUWlEQo4rBhg0RrPjeTXpWeoEGwhd8a9DS1zuvDkETd9INC+cWszwX
bN2+avuMashbm80XwBvYkhd1JKR3auIeXoLdudvIyLQAaWw4TJdu8aKYIXm9
hPGR7TwRiZDVTqFTXgRvFZHigH8ii5r7oYGIeiOtRwRwQZjnx1rMF1wH6hnB
DJOHb/GwurUgnEzyjmsAeXIm4OUxTilZ8wUkAfTygr4f46rywoQ+qm7+DsBg
Ou1eztiWpV/5l6qu68SHG2Sjhr7CYD3UzMfI8icggX2paILih2ZDKjWH/vL6
c6dvf34wtQpqoD5sPr8+wn/Ni4SPIEx1sGB1xBlno9oRddv9I1wTM+6Bq5zL
7fCW4n+O62cTiESCiXQ4M8PfdRN2cVcDsVRLKCBL6v98Veu3aXwP+WHT3IY0
+FCRcVuJz1qQk9H8zHqi/4VtdHDUbHKpZzJL0BtXWZGNM5EkwL4lxQxFDR0v
nCZWYYlJQctS60dEjPoq+htLusVbQTuZ4J4Hin6e7J0gPawURQRKXnKSQhtT
CQEBrT7CVTO8P6y3n152Sqh1Ej9zK0PPH8vdhr7SEtHHsf4N2li50NMugaYS
xrX2+1D4+CICvtDMxNdMN75mbr09LUJiNXkg0HVTDnY7/Y1e8QXJEOr1XsTt
EG54FJQyul709ETWQygMKtAcI/Q/Y/LVXevdpV8cJsNcJxSgK9+wMpicqV37
r3U2rxcFdETi9W4QiV3yw9eFYZFd/B7+tF6Rx/Lc3nNDTffg9rS2llTmRo/7
rSjPFbapqwlfehZivosTpJfdsFl7dqP6jHeR6svu0SlXo3XtxKkLLf4QI9cO
SbpUzo8ntySjkQViqwA6mucnBV/MFhCno+T1g7cGbmx8U0cO5I7BcNPr+M1X
z8vUGZZJq53J9aCB5rVi7pbwGnItqcipFRfr7c+3oiZWjnPxVaKkFF3sYzpi
mbJGu6JmPrruzRr2BGF3oup/OqfIEGfrVZARqeityGtEVLksW2bF9jPx/UHT
v0BcNUYWsHRFGXkU+HXRkn0vWSZvKtYk3o0rk9o9SAL19Ch0f77HsYsSAdSE
ESu86ojHS1fqXYsyBrxQvf5njcaMPxow9oZqkGyERTXFiNvSyA/LabZqWzMi
GUphwWh4dC/M7jr2PMWHWC4ZTvvFAPBsGzpWaHmfQMvxboDwnlfRuMc7mEmG
wH7LbckSJnvz77EHOvSIZTtRjtCQiJgKYQd7ANsvlD2E/Uv57EPiHdpAdrsm
v9jtmQH7EJvkAvE1t617h58gcPRuOMkUVHjPr9rEOY0NDal5QzerKS2zfqBp
VXELIrKcOFE4xH7fx1MynTvqsDG7PEHfPnvw9AYFyPeMBkgtxJzkP+GFah5y
RyvO+5nLwJ+QTjAEve2cXdn0qJLaTK+AozaxndI2uEA5TCQ0mi83+3gtqNbV
1IYEyU43HdQmR6/T2VMtt82JfiCaCyuWi5hV33+eK4USIyrp2LbntmQz89DZ
ArziEcneYM+ry4eHUrve0xZnyVovKYRyWy1gKwmv3PIuCDVwGde8A3UQR+AJ
PnOdWGYE7oqh3y/4NkSjZodtihYIS3dciPbsSK/1dIoB2fEcP5ex2X/3W55j
ambkdqM3xbWbhn6I354qPxoYHYjgFJCT2PwtWAXV7Kxvr06M9Xt+diNEl09Z
6KVYj3xIFmKTdjaPdDvzT44IqnO+vsTMrBlZ6d7sllmjXQ2tsGrirbUzmtdO
PJa7vlyfTJ54qdkTY6oba7O5P6wpVKmMJWhXsDCcX1IHds9YsR5go6e+su43
oTbafHPDJyrgOZrqr3QO8t/5SVfuMNzggn2qWSueWMSxoYItbLnvNq0tsHl/
Yw/0UUIPCo1qES0Pt84RSLI7IwtjXMNlz7SCw9Rqw9UdsUeVEIT0QFmD6cxn
3Xij86SR5DW6t/XZ+qdiFzHfqS048dLS5gMmtxIX8KrDIYEmSLbDSBBEK/6E
K79P53yufTbKu96B/BaM3kAz4QpXm+AaZrz0WW97pcaK5OPPs1wYbmpAOOYo
2Lz+4xjCclt3TPBsOsV/D3pzWCanPgjASl7X5iCyCKdDUIvNso50GKeHmwL5
DmX0T4xR8IkEAp+fjcfmVrUlQfcLji1MjF3cbfjwl0t6uwl2y/yGuhc7gJv4
WQcj5O8HQyRCPjCCUSfWTfLWa5zF+AjV0ZTZzd6CxuPxuETrYLxgiFCA6Kif
DD9nEE5TVaTgKghvjShXndtDqtN+DsrDlARc4a04dMGHuIJKSfJ5sJeCXGk4
KRLICLauMHegbrjz4Ktnih4SyGmxwRpHXA80hVan/JuSxP1fqCp3hFwt7mS1
/ooy4A7N6vs1ybBD+agPqXNFT6YmjwLPc5jcHVSUshZ876iPexhadmkX+cOQ
3mffvHJguGMVUbfQ1zlYG2Vl3badFyaoq3MWjtQeDnKPgHwT7RRrs+mMunkL
wU9NYhfy6gov1zj2j0GCDMmvz+5xaiYrL4W/FV68KPAd9STIti0Nty40LzTl
/ikO+CwNgVvzJWubLFAjfnv1lyXuKGoof5aVbbJ9vYZfif6N1Fnc+4dDyEob
+4gM/Ey7pPe7GtwSt0NVUCnQ6Q/jt/aZhefnQpm/plqOHhXaD0TgJWWl2jV/
5U+vYtaKXQqXYH7V+tiGEGyKQUKBWGSO+aIba+6BH+aqteVF6JeTEKXLaN8J
wwiUnwv2ZWb4eR+T5M0rHURN9xr5ua7wO6BdUsSYa7V5KZRnfyiFrR2wAfvd
cG0b53Q6AkJFYBZ9bff1AqiEZeGC02cd3BUS4lHME6ZUeUouHWkb7j5JrS3P
IhIhXGMF0uUnBkNSQmNC8DYNBeDXeVv6zIFCsrQIvlL0xGewNTlBjF6p7ai2
FhIBTj2uiKJHdA+UL8Ht1PMqyFNHoDcSgzS6v8uPmyaVmj2u0ueD53QpUblJ
FouRRVQR2w05BSBt4NirCd9bSkY8x8QKml4KTL+kGa97SjNGl6okPPHQ6q+/
O2e+A3HBxBw2a/496PNgTSA8E4pfb7/TMmbJCUGGxmygzdsoF//XPDRL6Pa4
34bTQp7jIwqwkyBvgZ1mifyi8N+XlRI3wuqjChIWB0Qi00qj4LBwfnHkcaY8
WQqra39eTrPaga1Zo8CgTKc9Bb4YUUQ0qTKGgcJaUY8goPX2oU+SlaU4bqee
3ymMEyJ3uHvS8Loz/vnfuIOKoykqqxcliWdBuCnxjvw6Vk4zeU7zguuwd86S
+IxMP13A8Q4csxd4lzlQQ9HGi01yj8mxAQzGwOplcNV6q4g+yU3M4FuiFNHD
pCGnP/wK2w6hxw26nKL9ez3hFdF+igZk+rm9BDC2ej6VoOukFuNtESzimawV
cn0NCxagT7RD8g0+LWd57vCydN2I9IpvMvWRBwsciqPKdjXyIZS+lHdo0y+Y
H+fDR1DJB9duPRDxi++9OY8i2E7e60dGDtm92raSvtDXEIa8PA8fovhFwcbS
/pCU5+bSkIrCA/pFkC+xYGqfn8Olq+2jzb+J8SjlcVl09JgHoETXu94JzsIa
twvI8RveeowsiEzwjwUVcZZNKIewr2/2XhE9SCHmivzM89OvnHOZ1at3nu7V
+3CcNXZOy70q/jZ6Y4WEry8oe/aUegPZiEsbqn3+VDsM2Zg0e4i9daASnRkO
L/SVfM2WbxizVs9MBOQ0DTb/Cy2DRlU/s6PYsynJnfWEGeWPpUtmWhOR3OXv
tFbiLOBszjXgTHlDphDiKaS60J54wrLvr4n2zh3BuimHapp07w+VCzb6liJS
lkuUsZsMhMe7fPysmlQ4gSBPlFVZl6XzstONWexUIjA6LSSjHGmE03uXBPZw
6VJDLYkMNkOQMrxNADEnRk0oBoqlToRtkqG7ceogN4H/QAnAWFdb14EStNGL
LLyKfPlOQfcW0hIOR7AI3dNiM/P94ZD9qqoSHpaGZP8kMNBC9wuwtcQS6lPa
h/bXUjMQfEI/6iriTMnqQj+wJjlQvAhyTeqmXdjZnL4ERxNxJ3SR1b51SWkD
wc7MSH7ZM2yYB1s218lsG+IsK2M5escbBmNQ+54Y6nyXWGHV4TVUdwv1A9fq
Rwg29KA1B5WtpGM/vZpVtMMaI7lW5wkIEwj9pKpFb3DUbOa8wI2vKFdaQ5ZQ
RVbCjl8mXFZ1q8y5D8Nr61Z6YDsVKDEgaaa/aOZPSEcuaXgLvYUwgF3JuLRe
r1mEUOkAhuGx1GiuwZnddo23Q5LoHoc/OIcw3c7os0tcp//P1UTzBG9eLMV9
ej5BfulouIBHkCYeDs86ZzpMoPqh5NOKyAGFLJGaDjr/KYWlyRa/oxJjPLy3
sM0bt0iHvvuRajJAB6vfTeOJozij71HaBT6Bdcu6OtDF4eyxpx/8yrUWN3lo
VyEUATnRlODdcUPvM5mqcMtRUhTGNttfV8wKp+FBotNEYyPYsPqweF28zOW2
ChTbUi87jfcXH3VRQT3iR8sDCB6kUI7P1XyGtAcNase69lkKTXCRDSjr0vID
ZQPUPHY8+dXfRU3R0wovJf+h4TZTi7sV7xyEHEwhbGMNnTGB6IS2Tvv/y8Zf
acorQfnaywRqS4psjSx7fqA/ebU/c3I9x0zjAb80dhgaR2dPRymbixz5XCRY
U3rtonegip6NiKgYK5jIQMT7+5tevfa/2MAmRnn82aK2snbIuFsJEGgV1YXY
LBG8qaGYfOFAeNUjSkhdmCayJQUChaHCkCNdUl5VZwNBcIYTxPpG+zz6+lYy
PCxx85Q7Gj9aLgycsTVYn8SsyW8tbuS0ku7HhnQRSsab7aufW10lrsEtu4L0
evG+QlMqHk7eNmueSF3bBvJ3bUWe82IrGNcbJMvaFj25keLUvMhKI/SsN5UV
Ew3qrlAe2X5+RzEX4i91wQIkskhyhHBTJfsa/+OGbY5MHu5g+Cx3cPQ9nSjC
I9D+sOqnUJof2Mc33jTZQ/ClOZRb9hwhMwrttIFy6Gw0FgcKiVTT2nxmoe6M
4gUQkh4uZ05gDrCzCO5nNQ1ut7cHW3fSUMOP5CUqPnqxGFY67UshrD54jxMV
vuU+MOQfhESW67nP74Ou3e3AM8qu9PWjEqkvQume/X7xm7U/DbIZocpYJrWO
BcS6YLeOwx4GOtNRZGEl1/gaZM3tIXO8RlN3j1VcoRl6jUpIMdhRQsTgYodm
wC/mrlvN/Ir4yqM1Tevb6UALEchWHLATtBQxMwi1kf67gaJdqIJzxHdLI7RJ
wPTHVFTi4VoB7kzPIuXu8RAKpVjacfQ9uS0VanfcYbUgnMCSBTdmKnXUIt+5
uESejakN75o0wMRVhfG7aHRAUNM4guzIaTTRxDassSdYIqbFvcDAmTyh9ofA
qurycjt1aFQ8NxEMM8QhxrYzHlT7uURSX20uQ3rBN0mwc66/DC9FouZ5IQC1
OvSb0YUy06i5i9+hWzc1lmoDT0kEnZwJV5cWTGZlEWsNXTXGPRdGfGrMlrxM
TrQxyDFH+9I0ECsjOQ+oijsKd396lYySprSLdmcBVg2iaO7tbk38wwWEymzS
Blv9c0jgnp2HkMkezcQ8M27DPDn2cgt5qhRqk+OC1ZSDQNDkOyiCz1vQCECZ
psMgIDLeLMIQNXwxR6FnixMuTEikICrHq2w8Vlzol1+6JRb0Jkn8H2xjlVMk
wrO8izkiyh0A4DLixaUX9nq/bgRHuwBt4vfiwvxNptXw9V5zchmet9Izju4q
srVnjs8XjA4f/pSirYBQ8aIaqzqs7KCg8D9LXTUD5Pjh/faxlmeWfu6/MPcI
hEF07nxUVhz/CosIyiPWl6LlZsk1rU1QJlVj6MUcbIDdo+A8iWazlc0pGLD3
3EtpBoBl3Eagm33FyX+z8emOYJr5O+cMoYAMj6vOyvc0Jv6OEG00ZLqz4aYX
59gIPJOEhtgaH0mnvWnMp8RqpR+FgW28nIsT7zbjcD4Mt+6gXMuJeTpabaHm
SHgXiqLyhavVXx8GSjvVtJZf66jMOU7H5HoFsgAmfcO98NyjWlg4oo5NEeUv
MzN1f6BKi9JtOd0yCjQ2GlHN8L1E6/twOUur1FYtbDowud/jSA/zrwC32H3U
/d77o3kEb5RbJPx+ZA4LHxEphaaUjHdLlTXhG/dxEXOUZmE8TxJc4SoCf8u/
FLJbeqPB79S1Nuj2Pp0asIN1yzn9Ips67/g3YjGbtbEUR6lBckJ54W0n5J6f
UkOOL3Osths8vuS3LsjqKPvVyGffH0vdCl/NWolu74jCt/ESFAwyydnRiw37
3oDn1WLImx0+2WknmsmD9f+FQX2ywjJD+cWusBvmH0pZu6cAOJbPk4pVOttV
1VPrCOWR3qkqAqWWkEp2Kck0GvhD6rtE4GEyfT0JJ4PIkuT1sldWNfNDBR1V
VPKdIucYhn3HllVpZhp/Cehlbcw3fVqG0v/Ahr+RaB4QD/L5Tkk1j8P7Bl+k
MVjE7V/92dW05LecSluQTK7b0/P5xNI8UDbJHjhGX22THhDUPCNNwDEclnik
8OKoGP4sKknFIJu/i2hYvVXv1Sc3mmhXFsD2+aUad650CHv13b3BWALno71t
rbrd9HQQpyPQmVQroBZZ8fJTPjO0ev9gjRTLYv3mpf0chp6b45xEzRJplPSy
scH5yTxn2hGojE9Bf6Bx5iw1oahron55C4ntCDClKwIgSqfOhHfa6S5PbbN8
mvWKcV88olM/GCzkOzimqJsr2ELGF3A87/8qvR8FypiYZz76sZw50JZqPtk5
lteYU4ays4jB0tPxyZ/C0p92C/4KT9gMrVM7yyev6PzuQN3GzR2ugbx5JcUx
ayWuFbejQqSVZbV52DAI20lnqBSbAL9uITE+MHWfeN4sKaSHrSkeEtgzwZ6+
F5DDK6KAamWATOxNxqrPR3JQHna8gY05Pm/K1ZgZA7gSQsl6I46CXFR9KhWG
cazpnd135ld2SyyFYyJ3Y9MkH5hsHpn/9huvzBTGbw3gfUksiRi3SrVYl3ev
yIWuoxjYEvjH024ejojIvRqh2zic++nvNJvPqeUxWqxuYd+LdnWFW8ybm5FF
MqzcBydriXBsWUVa1I6KDCOpIqsXRe9996NCCdm0zxUZi/3x58T9pSp/UN2D
8c6FuebNl3xcvyTLIpSd3C3oOsOlXpFJNXqeSpSURDngSE2m4tVBXS1trOWp
iyf2o9Z1jmp8n6XrMb3l10hnw7zkgSAu9F6wBPUJNtPhvIpza8nZjVRxOOs8
wAzfe9B7mjzhX1c7/OAKDg87BI4EkSevq0Sg6iwmXhA9EZEfiWYmrP8/haZh
twLUmyPg+5c9N/GbkAax+btNv+LkOhg6lYuW/6VAXi91toEcL2Hvz0YWFVkI
4Fkm/cbhFVvU7G8x06LJHS8Tf6zJB0zCNk961DaXoCQrH+D0dN3J/CA0NWTF
cDsvAn1fIhxbC/j/0eW2g7UN+IjnW4Oa+HlV1BQ04R0HpIz8k0DP0/wOqpLK
iqV35YI2pVLS6friZJmMEtySUYiBslmfDBVURdtXUAKSLw5jx8b54AvBeghA
KMZd746yr5IC5PZMnlBlgTPlw9DlVJ7qwqXV3o1ZysHWeLe5SBQzvi/91Ut0
VMIYHQ8FQm0pfa4Kft1ZZXEBiaB0W2FpIEs45NPhey/h18iCzG/b1FpCZAeQ
0RxHTrWKb492lu8rFrH42a8pppL5ql1Uz84XMwdHrkvkYNBGuADVxUBr623Z
4XapbUfjniB4qxyPkQT5hJAGi/1Hp77VU4Lq5VlwTnSyZv5FGG7gSOwS3WWG
TGEYwIDohWBpTjzsXFU9/CdniGFeyZbRLlWWsh3ee7jZZDGHxznDlFR2PvSt
ba8EO2zkxUSSLkgGpEM9LVsCMitB/PIKXVDXJwnsiDu008xBfV3VtvnBHUXM
q+jjmv1biYwepVrF72SaP31aUDmyUu29a8e016+r6enNC+ludF/Xe5CwG+GT
8hwvkr1wRLUPOt7swhVoCdNmLz+M6s0eqaBvFHm5Twm8uSZbroFINactnUQq
v3LsGnqwELvUXJJUnPCtQTFEcxMlDf41AMICoRx3H+JZf+IVM3wTrMslQRVL
2cDLpRjySUQ/7QJyauzSqxwROjis4INK8A/UVdE73b2bRpB3jgfbVRVyuAkw
73RQ6FJPKWy/V71pVsSm2zz7eJKc00vwibpopTK/CHIMt3k5NXfdGG9qRW9N
j+aJhUdzw8ESTS5nagm833wgyIXfRYUwdwLOE8/SXt2BlHxNyGxwkN4oS0Vc
GghSJQJBHNybmdtq08RUoCfawQ1/VNLDGbgBbr62S4ZfJ7c71XbABBdMMZJN
AEqxP7/hbyUnry+GuEI7RjnDQpQq4BrWod7vfN04OHiZsxNK+RGScXkVRB4P
YJKSAFLEq8/SkIOjwUxkAHdTbJUWobzveEvSLxAT2+Jnt7MoD/sMwr6B9xw1
5jIXT2lYsuzeP12GHYOYoXqNF5H9JazlOCJUHCsgCaRrO+EqWPq6D5TemY5m
wD9KEz7RZc5CmnMqpC6tKVazrdbT0i96rI3qfw4RwDlTEZ9Bz3HXORQiM5Wy
eQNIj8U47BlhsB2rtR4NjX645bk3cfxWDmhOYZQNUkxMjF/Dp+dx3KYXtqqo
CU/96Mdpue0TAwR0bzd+NEstWGa/v1ql5bwZMjO6+rWzhZe/8d9U5AMf8UK2
Onz6n9z0Jc+rGtJzVcHROOERucNLmc2X3pkeZer91To26owxML3TKJzceTNo
TdVMu5k+brJXxDwx1oYh+ss6LbrZwd0HN2lYL9AQH6J17FtHT4qRDbaYNc4a
4u36xdRcnelzg2a0/SiFpIYqtPPEEY2r5bVsZplZMlqmLSM7AYxNvvUaTF71
EOZZJoSXVtmt08s4IUpump2+XCfY4I9lRObcQBcYyZkDcWRGEdCR4/aGmMKB
m9I2wUPufsqSKY1WfQNys8cMLGU+9ohLTiwDnjvTLXUfcrLZfjNJe/7k8clR
N9VmHw4L0SZhTS4cwvcQebtIw5AK406TMIHgZrww9t1l7Vkh520zFzM4v57N
ePzPcA8DCPVwe9QwYAqxrgoWa5DPYNYrGAUMjDNXnS+8U6psQCj+5xc0tmLo
zUnFt8a7B+VqWlEd9SJqoXgsk+cA6NeTlPTuQHs9Ze8kelIRfNCrVKEmvg7q
KRC4y4X9BCrv+V/BBGq5486kDBclG179J4DFwZfpkE1NNuYr8JtaarNbIpjD
lfppLJW5CnqbbdCRXdQzxIIqXwhq+fB792ic/LJdTB6T691n0wKIGhjCWhSL
5Ak8tGI66miqSFPsyuOCrTT7JquuIfiXi1y7aB+ZG/kqPZwhNpzw3LuUyqte
vjKzeZcpF0HrpGf7asogeTG5AEi6tFPnr/1Y+8HwWE1nRTTyaU8j6OIe9rM2
gQL2GjtabB84JfaFEbHlf0TbOchaUogy/pdCvEbHf6VfFoZfqPgj2Xh0gNHw
WNG8fl7bUehUTtpbmJOHdzvMfG/1ZUgRpxQkHPXssqfQJ0cWAwihG3XPfP+7
g8ojCAt70zahiRE/xp2SHl3pAnJgXOgnPDfTTovtYUi/GvqjmV3vs5kS+Q0O
uX1plSIIeYVmVpOvZjsiAoNOTnphmK0EXt1X177jLldIGz+LIk42sRREwuC0
plmCyULoTgNKakeYlI3uAvP0Vb4CPiKbtaTNDra1TE4wFjaAycnBElJi4Q8r
k5OW/QA0ElWVWQAug4JR5o8O0dsFJBiCBnjbcAohL5QVQw4U003OSDOnmMhS
nvRdPvrEoENfecR2YhNyoHb0tEJiAX0VLrrIM+3SNoFJX+7zMUTcxuFkaMxz
d+qByem8mweEdeZN4eMgOYWs7LYQJUpSjWFks9yNLfDPjp+S4klPphMaGsqB
270ETxvai5sj/jtCeS+ZKwlYyjDyXBEbc7ocEg+tG2mYo7VrUmFv+kzjhLsB
YBYEWFTpTy+1wjimwk2VT+YX8T8p+p5OQhz8ZTkCejd0TQ4AvjbiT382rq4K
iSMQIJoFZZ8pIpoXxDaApN899O0QJ0XY4LynViW/6x0FduTbW5sLEk+88EWy
TQU70HbgYkNY90ORYD2AjL2NJuVsoGJ/kOrf4zPo9cVoA6oPnqhLjkYSzYdK
3F9rawuB4Tzkq3yUvl2tv/CuZvM6aaY+KNQxrBpsHtA9onuEXylCCZK3HwNg
ox9UtEaSReiW3Qy6MbJc7Q/1n8bqMEQxdPh+7cfvW0Q/whN/BvYt8L6SGVAL
PgGRdxWb6wNUS5k+OKTqgi6a15ASticIYBNI1rfiX6gKBfIh9npYMYf1edwI
e8nH1fUlpAZByxHT2EPLy0vpF4KX7vwQefrf4wM9sRE0UDzpICT8g2LAQkPr
QaLRd1EZd8agwSo3uHaP6xCUuO1nz3f2rZ+NnZ33X/mgJZNi+T0p9l8QICqa
WS3SLC9xs9L6EOfsNb92iPt88P1aDQnkJqtaXxJwVDSMNqnaEmMfYvgYuler
vBpCnRVE+enuJ2vqZNslvyOiUMg8J5EGztP9+J+Z3OM25AgTujbOscdzIRnq
GkKQMX2EMXJZeXgihfAuLLMoGJHW1cv6NolRGV1zYS+FbiiVjvhmApY1wXrB
qxzh+8pdxiwrL+3njrhO/+XGo0G9QfIBc0+WIBHYiVw5bQ+rOAKIl++cmeA0
a2vsR454XqMdtSQHYN+XUxPgFI8z8r8JtXdCMw6bUxQTnXbwRRIC+UEwXq29
Rz9f4CbN/H4vkTBriEINRjHQhWvfY5CPtjtHizvO1jrVCJFlTOGyODlpajE9
0uRoufcSIfLar2X2xyrJv01tpdUsXtVzR22wO+gLl2Z8IxSIAaM4qUfM+aZY
OO6wobVfbm1vSBwoIky482aOeoI5c3/rjSMaannizkCn6cdJIzVIvH8eLgOj
KrWUYMix7P4NnmlOdii7gboavpwdKQi50kZ6CAljJ6W4OwRncXRl3Np76nwe
LFEmX7H26k+Eji07q6T8EhIMS6LRB39Bl4SaLv4mMwouq+5ogSzaiiSDFiIZ
8yRaSuyaJVfNwn65aeY08WWAS2STYtQyE3A82xf5djIgGE1E4GCb4V6Ky1LN
8tYuhm4fdR1LWZoAFX5P6jrMiuZ3hv4IioswRU+BqbHNGXcMNe2x/cXhvUYQ
zXh5pdRzlHnF2YUMbmY7BK04hJkCtOAtKQLUcGSKzIL+kjGo2lwWZ7ZE/Vi7
cBMirhB2k69tlfeKEMo157RvKSRE7P7jEB3iGLMARGtZ+TZUdVDdWgwgdOCf
XKTutmEpHM+sVyNVynTwa0NlIPJbK7DoOvCRSqUx1SFblyb0Wx3lCRqVqjzD
TUuQcQckmZ3qnIhQ/bskR0K8IbM14yXIuQcqOrnXhxro1KO0ifk7wFrVAd9B
JgVI/ngv+AT6VAYOvU2O/LxvemV/lmJC64vEFOcqI5UZ9yM/qSAd8O3W7/hu
jrmbyJGVqEbOWXI8O1/VU70fztaiDwvcvTWppS1o9vqHjQtkDTJJE/AKR2jB
DnKrQlFou+U66FWClqxpyJm0kqBhz6pI8xqgvsiS8OGyr64ZHJXZuVlmEe4p
w518uUfpKn+28qmOqiu0wLbxgMEH4JNGOyyy5cePqP396t7qoSVHXLpGVWaj
ROpZpcYhTZB/+1x3gLKWyfIUAtnFRAWmvnx34+Dac/9IxL4e9HVMnYpPgjLW
BZDriTvGfWca0NmsumGouhufw/tGUw7oVSmYpgqdkhriZNo+udbKQnb3DfRw
yZN7EN2VxEVdXOM2qy7t2bLoW+11Dn+ylJDH3p9kcr1qE1guMzGTZUgr6gL8
ox7ElgTv4lLJcB3nep/fPMvZakRsDwszGILxOVCfwMXBGvuCMFokZ5jvgIDd
VE01vp8FJxl5iK68UEr/HLer0tBTpDksTHuVblrf2deDY9BUjGDeqrJ1W2PF
MdzCl5FIhdpCyUY9Mz81HxC8AoIdj9H3+Xg4ljk/sIXq6EPquOM2khc/wWLh
L17qjB4sNnAFtJCNx11FqStt49brGSc9STBSmLdgZofyZYhpr+dMk4hqBS/P
6g6xg4wPe7B9bae/sIkvZIqA3w7rbeM8I9o9E6no2d4vwF/HUdO2re4FyOAQ
qfrJ6inOT7Yr/bT2aHan9oSUt8sR8+EcyfWiGXDzSCGs3QhIc0BoAZw1grJH
mf1OJr/ijvQfm6hdLBAt+UMVjfNagc7DZ5bgiunAqTTv1brhdmoIclhP02WQ
Ntpoq9dOccBdGSzJ+caVzHMoUxzLBq0C+KFxUCmNINn3JjFmUHKqV9XioqCJ
/1DEQ59CiCRokZmBFcwT08b20MDTW5DN1PPojcmOTRypoorz7TlB1vCuEaeh
XzLOzxvWLbVe6BYIjDqxu9czQQJs9m8b4Yd+JNfYYaIrMLV+HSW8JFA8hMWB
1udquJrmqT1b0JITMZ3EHXH/AhEc5MqFUKI6ytskGy2KJqNywCGLKun94RuO
IDAovQunt9J76lWbBk9oSErHGYJG8zmsAkNvpbpezI1NRyliYuTVKvMNOo3v
VdhlspwY7njqVB+3o7LBrntQb7SGypGGB6KCIcJYyIlAPczKHHsooj/j8wQ1
wUXMnQRpo8NXVBSeIe+mPCP8pDKTVXKWXc3UGtidvhraz97q6+wmtTlOga24
3OE2jw7BnUrAsqsAMCCMMFmaUGNgdvwGEK+Xu78RUHUrvAJ/zdhJxJ6o5oCx
Hk3lHZhuckWuOYA2f78vhU2A/wUH95SscQIkb/Ax9QuWSMRilHp/lWj7vCut
DqL88SoCZksFvDzKeO83vBMGqFnzHdGbMhwyM+wD2yMJ+rtkgPZBdwpeKl+w
T8aVEfcxSZh8NDvzijwUNQL0EJaVttAHVSZGeo1zg6BlVEp1BErKibzcWPma
dAMLO/4k6IxK1P9k4t6/vxVE2ZVduDQ80GVoesPAou57gFsna4QQ0PcIKsl9
cn5AbW7OelSh3SCn+EKk+oj7GQ8fVdgLHsYCtv0WlIBpTkdU7JABR5Cy/Wtl
Tq+0cP+TSBH2UE9Ys10aMY657OsYQJFT+0BAmCfnlMFZlLzHaFR4se1M9HQX
w+xwnOoXYPEUt6xCfnM4aY9tMQF48hQ+1viAypB9hS3/aYe42wKw/LYJYFMz
3Cmf/zuCqJG9xPOtgtuarSha/zW92q76C1IH7L2nciPstpC3bJtlERyayIzA
iiOAE6AtCdZ7MI2sUP23IRUlumifmW0BOiSJ3lTY0YvZk3AIFoAFprvYYQxs
kVFjWEjoG6ror85E4BxcmTAUnRs5NqAbUcBIkmfGZh7r6QTkdTQjCwmopA1C
7zQHgD3751DNaK8oYQZDjTpqpd0/uIGyZnsZfvutg6+/Frqfs9qzTvaYNULV
uVvIprKbX90FoFrATU3Zi6znercG7eM8UeI136E65yEMVu4Y/C+AiF22Z5q2
JmApoQ7SIzRiGyw6EyziS/GZMNbAqCPehTNuqJvfmGettEEDgsh+lvUeRSTY
iR6HMqt0GXbFmdaSn5zw2aENSFEdUSm318keb8OlQDqzVGbQZRm+EVSqt4aD
iG1A2EcBit9DnT3vrIr7VKPijEMtzMoLY4M9l6ndEuARktfaG4s9JcWTEykE
Bg6Umo7X7gcGi0Wg+Su2tW5jRmBOQkIr60eguAaDgMghUgaQGzBSJW/vi4yp
GA3JZAa1WKVwKVzoBrvR0T6bW0J9PxYy9ejRni7DVwWQPH/jTmvQ9BF6gnw3
z8JcLkuTqZRqrcmpZJEaXEJGnaXe4wpx6i5n81/L4XKLGpYWERfRfc3t1lvm
CLp7C8pxwAYFgXTnHfJQsrU/ze82enRF1bQnm9/qPgvZ4/1ABg17+Qm/XXep
SIsyZHMymSjJtdQFycdn8RXChXy8Y2x8uIWSISZ/CJ1bE/k09plzUx8emMnQ
yzeztC2n2awC+KhZ+ULpW/H3+4MQ9Mm6Ay+Pl+dvfTUHlrm3uv1NlLgSpTJC
eTaYE6QUWXitVFFVW1BBnJAO2FZ5t3+KaDfNzbWyWeNSgh4mmj1t9i+qm6IN
p9i1lGsZE6JGlVUT4G3vY8Rq4kS4u20oKq9EBm0Bgri/DlCEns4/FrMycipZ
XPnUcla79YLCyPt0dbjQ+7wKoO4a0LQPDRV++WswBh5Sp7aE/Bz0toBNBDzS
nkFedHYeHoSdsI9ATOkv//FOjpYCEpIMJrgkzzl5AgX3+YKK5t0jNZoZrXAx
7KuQAvLXOgIEr9usKjnad2iCdeFcucheh73BkmJm6njZorRky28oNvzutQh0
cqdrcAxgaKpHn9Y6wk5f94RO8fYo+ZM9rY/gQtJEzGwgvYSEPyQrjbBlmKa5
EWGNflPN7GKONtF8r19pqW2w9DHNcsoocBk2C1MBrO0V/j8DcujjFQpRbYKn
9WEc8amt/WIPqmcXBq1laUMppJOecbFuWt6NbWhfnvNLL5L2ToUG3098+09a
HTtQpcwlAuwptwDi01p+/NY/Vqm5fFAD4ANk7O1ev7W5jvlxpmKZWdDberfi
KMLh28wcC9iNO+Yu+QuM7uAiHFKgmYT9wdygFOVImU7NcyGa72Txzh+naVm3
DetXOIQvlmothfFPtvTg9M/1xHUND6NlW/YndwVEo6HpnSbXgZ8euIVYStYb
jbZ+mY1k76kFWPbRVKCAxuqOPwymCoUruF8+00/YJtqg5qUcceRyOLQVTQCn
TiZ8IMhEnCjpJ1GgMy5Kr/Ey8QUNOE0ZIR2imnCxAL8/gTJQgFjmHKpUTx+r
D9CUANManZTKmnaJE0ZwUQ8Qgb2aNbfAZPYggWR8+nrpCeRgI3hz+27OWsDs
j+3x92z1rN6IJGS4644yySn7la0jOtCa7lq7TU7NWyssG3uyqNe8MK+sx26+
IwBpwnd7iBE4hEHchhKwkRMuC3fTK4ctYengzyglxlh8e9f+vAXCqjb3bhaS
Pc0k6nner3HlqFQZxqpQp9SKtmIy+BXrwsKzjKv281+gfjLl2lRairupM/km
xHgm2zBBAeVJ0yMeGltF4sm/gtr0KuNQHUfEa03rRCw7yKK2Fb7Tj/P9Nka6
kwkw3OGXFB4w8ChgvZS1G8f1BM9ym+opMvdz+mFrlUuLItSy4UaACWxDb8g7
g547/NjzItxjxvw4cEzinMZNZE4rvnsNDwLRUvmfuX9pwSpG1AYvFCYTxgl/
TCR2CWGaXsuIkd9MbuM9T6QoWfEYLy1YD7qHJ0miYrBfTUeUGFifHJpfwbwW
SkCRoLWNNEQ8FCLCEkIgnr0wdfO8w453hCg8IDjYcI8GfAd3UXqjzhmu8Vde
bJLKvdIF3RRzQph1gFbfz8yff0AGM55gTHdSYpY5Yr+KbkDeaSEVcKVFBucr
uT3aa8V459DSvdU/u/Wf0/LEfLq+60SOLUL5CKJPP6uQSfcIoBP9YO1uEBDW
NOHVjVLRfd+sdoP0zm947fZS6Xs27/zMMjbSELyD34x/z7aOUG0627LoE1j0
Ra4nn5/jYfQzQqYT1+7Vu3BzvpznfvP+7jMWhcVEL+wYgWNs0tIvmM31sqLN
9MSzVasuz21wLpJJolUuM4FxId7agaVnadUME4VDjFbH1W2/HRny2+uD+ea4
/PWZtiwg3krRj3EITXjTj2u6QykZucSM6y9Yd+IWjPXo0zedB8PF7K+pI51T
zN9Kw/9f4RDBaTu7/1SktmSp5NlvWzzbE6ZBGbgF7SRXi1P6ogfUnlcHvdw1
trbJjKikVKUABYE4cGbbndZFRou/UmxyR29h89yHTwk2gTj1RxC0P9+QHcd3
7ralpjpo5gsv0G4zi5vmBi9Y9ac318OIsgXpbtQlDjUN7Kxd2eC7bhJh+QsQ
9e5R0sWPrWZEz+xoqzg7/39MBUMd0waz621j0ewCKkabCQNFoACus+Mo8RLx
EsivWTgzKgiJM/2gUtU89qCL5st9pj2qS/4oj9eqzs2JZvzNNsFgEWqIVS/I
52UvRup5HaP2Z3SQgZU/G9Iq8LAK8+trC4jAj2UtfM8mdhPxbvuJkFC3Q+G8
qCbdotLPkL1CUM35AyDlk1a+GeEz3Yd0K3Bw7mAltuO+xZabZfrIgqyYQLaE
svE1FbKUtU+S2vpIXTIGecuU26/x11e5uzsYajN+dFVz6CDbA3unFFjsi+Db
dTbP2Gfrzm5E3LrFwneYXonz7IZidD7nxpPDO0syEEE1XcX3mUOFoQHY/eGB
1Qx6C22znt8SxVDwpf0Xfhc5r0HVat+JzsTWSv1354vckeOJe/om/MheYA6u
rCnDZ/8E61re9yAV3jYM2Ua0ytIJmW3c/N6w6/BZfDttV/s4ZG4FPJCV4BQ1
HaPDHn5SaP6B33owKXji8Yb18Q2gr86PQMyPUAmE/C0DYCK9ALdEvUUY58RK
cbl0UFouazUDq4zBpMvm4nQvpcnR+Yfc0EU552Rt729dKNX7tuPRJhH1K/sZ
Mc5wWke+C2qLCwhJPqWZ8o9a4JSKfSFgomDG1FN/OLAvRCfOIqX2DVnyek7s
Ut6tfCFGTrNuukxP8BZ6OFUYGR8eyE74SIvaNBg2H4E09SCh21iQ3erc7Qy0
fXtc3NCeRECD4D2uyn0ZhB0QRGBQgVLAKEpyTuVqN1wVb9mKadMTbzzvYAxm
R+k7tBtPhgpvfCJQ+0v13XBHHHXlfiUO2i9lREafsjefkTZ60Mg2f8ydi6kT
IqwYwL4p37Vf3Goa10/fus7SOkfBrk5S+G2lyVzHdIpUx02bfn5jDdNqxxLI
BQR+I5dTmJbDawl6XEDxFS30rO02ZU7D3T0CDOMyhq1cKyZa8jG8VX8qP0eI
uDV1IZUkguEJ3LrsI/3NOvtYPUKSpdboTP+4caHsg8tuzjT9gHCV1lJzcPvA
YuYHVSRnJrSKvtCuWYbVOmEauOBf+KpOEplImr+7nMigX9laIMumyRT9AMkm
4hQcBx77eKU7chE3pBv78W9reDvZhO4N4zjIFbN8gKU41N/3fdAat/hCbduW
50RBHqw57BSFiJOzoeVPHQp7mEWPTw4OtsgzO2d3VtQvDWZD9cCxzMKWRB/4
QX7SIDazJH1QyCbds3uFsE3gMxb6clWR9aleWyJqewLAze0Qnn/fcQx13gV4
FFboYtOJKNYLcaCtOGhLapNIEBzXgsHtkOpoP4IYU3mT4uxtqZwTrfaTMq8L
q/sbnKGgcHoD0Pt2IX9+ZAI8Crsw/fCupkdkA05ed7507WwRAvaKhgOyz6ZA
1u2PgrWUOwq2DHMgynkU+Xe3M9ylFL0BYPPSw6eUIzcW2SqLmOHd/uIxipVx
jHfDd3g8qejrBH7Fa48ZOstOkM9MkzaIjqJG51ILt1xW0b42IZ6B+HX/tCGR
WYs2O78ZzhsNnR1yAMAguDn+H9W82JAko4qC8gb3h4S61PMTb3TffX0yEsQD
ah0gcG0Qg7U6UbTz/3Hua5bmCLGfLqMgtDyBxDUIAHv30SnQMIkHFSOqB3Vp
UaIlAoh0+bR37gnMMkazsc0qU+Bh1+CnvM3T3coD7p6fmj3PrDNVD29YKi47
kww7C0sj/8fAkOBlCTozZrIC4kZUzerm38V2oBSPLnbLAC90nScV8ouk5wh9
UsotRxRO7JZzfqibX4j83khJ78IAjuvFo5bkAOukkDGHuVtQtTjXsghddW/s
fmWn5yvTT3Txo2xC3H4sUjWg3DGZvX3rVaPS3ydrJsiGkJvWyi2trq2x3I7h
hIngulsitA6Uu9zJsIIrtk2Ed/FryewowxfoZnTJuBhDi0GkMHbwcfCBAD52
KOlVwUNxfK9sGpQQ6Dn63c8+CVrNy9YluYWevT+VEkGalZtvutXOqwpYTWhy
vjQV6lWz5+zc2lMQLDa9NySEj+61lAolAzlCjLka1QuHZJPd+nfEtbUcf6Lp
aurTZ3w0ea9QxsELRd29GceeYi2vF8TSqVZnX60Zwva1xB851Rv2inMs++hm
TV2R7Zyo0bsAdSLy0JvnVrs4DlD74Y+OwY+vSKV6Lwcy8UnKIgZ1Trgqnbt+
752PLOchzKRHOgu7OAK4xCxOUf8blHQ/ipJKPx6GVN2eIi5B04BvgViXZwwV
8hk8ZOPrdEGJZ1AuPmgo798CbJaLTjpghyEY1IwtTRaUh6sA3QgTqnBKyYHa
z8OikgsNOyCVVXOh+dhXCAarMgpIcTq/EJ79+Z2LbMFhyS2LQHrYGpobKa3P
sjcL7xWwzrnGVmVR5vnLx85I3zHvSiO653ric4oIPl8A5nEzjHSk2ktwDzT4
qgHwwnCDE3rxEWnQYGlE0W0MOqUjaP2mEN2ZunO0g6zO+f8mTnuilhUyi0mH
1ewuc7HA5zSOsrIYYD6LKMrorrNiRk3VbP2/aXBR1CsCX5t5vFDh0MM/475O
akLBhEQybIHJzyNb1jXBpPu7qo9Ux7fDRLGw4qbNEVGfgy6hkZGztG47O062
Bxg5hHUypvcoXZtDzH2hvYTwRLkrijjsHZslaHltzKMox/NJqDtQkjDC/opb
hxI6PVF3bpZejm9O0uCcQEZdZiKea1b2PSLV2Gxo/Or7qGOmlCZJYnEIqyqm
kXGnivOQLYGMkxytgjxIvufDtZySygoYJjUpQjqgRrDtAQZ1c+aMWBISJA6+
g2oxU+sJyyhAW8UsCykFlT9b2Yu7eGIYFj+z2QAlAex+b1CyPysDazv784F0
IBNDyj5X8983LdIUWCdeTKjLETq+fSMlhVojBFXAz+VkjLa1UnWqcwQlmk6K
l6EpSzp3+7SUmzF2u8fD8r6eV2s/7+zBKHd1nznS6rRQtN63iv8HCKJx9cBM
5m6cJTNKUN/0ez8tIWkblkUhtoa2NQYBUeT/GFV99hWD2iPlVXZMgp4rpEpC
KE3tMW9Dtbn0usShh6Ds5DiHi+WZcjYZYltjLkYoh9jgXnzBv/TwvaW4ns2q
38ZGlE8vEL7oGpS1+1BhnyGPGl5AJ+N3DIv+SK/+KtcjBUZ1gOrfbhyHfbjP
RDCA/0NLhIgS0sA0nxZTjCttWwdlBAGDkHr1CTLLPd0oiWvr9CVOLtCr9XyB
g8jCjQOqkX2iNnWyYD79yccPvvR5pkkBqzewSmc1H/WDMQLSsmVd/lUtkK1g
MhVBiw1ZncVfRwJ5pyYyVYJbOLjELJ6CHIafrwGd4s3k0qrFkJE+6pDtGJXw
sKl/7ta/AqpUVNOXe0tOLCXPMMnBeTe7hfnsXhrxb+7hB8GvVkKMxjyhiAaU
c2yqSAhab7BkAgzfQeKpgf+pyH31x5c4qLqU2sknZ2VgjcNXD1ubjh2q+vQi
+q0Pd348tbFn7lCFF7NqqJkf55MNTWoT4jOMy4Kn/eOm0rB3BqL7wjUYD2Wc
ZC+6uhEpH7Ki/ywXl2c/NFCbK6iXQGZfZMvEba4ZwQ/jwjAteIALnY2CivUE
aT5d7GBIVlaMjtMUdfWPgvl+0vUH1cv6Nvh9cbX1ZOPCrRQyIvdiqM6ICCCZ
fJg8Ko+e4jnD8gU1mzdYc5lovUmtL/7PsxExBIM0ZKtM9fNDr7/6LzzoL3Uc
7Rdzh7NDgk0LsNUhkFQ+sxmA51iX3dqLOE1dTu3GuntRyHCXwnxCKuffKThH
uKHW4Mo9Newd1iiUpj479GfzBQIOcYKvCy/ay8CT11fglJ2nd4KNy9GJMY+Q
KgbjGcnlJO8NeUpQMs53FPCFF/vOb8lRbd0hAKiVUbF0bFFw6Z/oY1oJMxsV
g78tSq0HMoUh7fuCp0c8ewFOyFx4UA8Un3LTPT9a7eZdA/LGVMHc7oyYmw9B
RISr5NIhZs0N77ywkkWQkVBfdOdCpEVlKqOmMWYD2TIjtrQ5NQKa2zTEa1ez
tB41SAyEDVaCCj0uqYsMGfLhn2eQAHvq1CQS8aHQ/Gvdfqb7fkH3RFER6e+L
RqDtjpB6b+o+TZnxm+mIyQecNGBeu6YMiHV0rka/9BtHMth7wzqacnztRkfF
3JI+898Jk/fvzoIcqiwJQOXL5DV2FBg5o7t+Xgo38f4n0fSpz2n5pNHfsWzB
VzsjAgt/ZXlgKvBVcHEF7vBUuLi06zK9F7Fmq93y8g71bkT8W6G/9rKpUIPt
R79LcBTkIh3QT8XJd1t8haTCjq0zdnU0KuDJNXmE/e8avnsIcKRDqdu8mEfU
bddEzfQ7yZaCJCXb20WgrdUZ0DMpGNJRqA8HPJ1rStjyonosyOCQcJXCUZzu
hF76bxNcGeoSsF0PKKPy72pW7TiPEWovjqsZyKhnpZDRr/wvX8J2yxICKja1
GvrW2wzELph9ITH4/MD3SiiQ3RjN7els98kkszT1yjPeqGN93WeEzJ9FCy0S
TcS2Hl0ReHgE5m60WD+sIQMCJ/sHsIw9WfHiKcHfMJneGPNTFuT6wBQzmjjm
cD1T478U4Y6178/0yE/Gln+VwxlTw9FMmRWofXrVguu11PWEcHdN0VWAkxxJ
rDQchShPczClRZ13KgcLd8QdTwbOFdKEuoLJrdsIy3t/XH0KIHWRrWn7BjIb
8Ijh99q6bhMKrCKotCdM1BEjyodfhRdN4BSPeVrmYYVKfl6itOF6K/cT78NZ
F4at0QsCv0K+MX0lJBImmT1xXIUyHIKAS1N7Tz3pSvBn3wxdxngKIKBrDF4p
W580zJFhecjCaIR2WyocSQrNfymj8ACvFzKztIVeZTBqj96JAtgh+JxV5w8U
GKQoV1LiK9GCAmXt529kNhAzp11LtD7wjoQc30a/N6zeeR3xD0QD4V2yXkAo
CYTZEMwmKc231QCw/l3NwVi0m484SCjP3AJlBDJUnz8qij1pI6LTvqtTdZOq
RMvjwTnVfeGDPisEP9SWdfKAWfu8N1cJKT25l7t9NjHtGhO2n7NIrJfA+2t5
kcmmAT+BrJu6p2R5XCCT+/ruSN5PWlHS2Sk4a6Esp2TEev7x6nfnRL2rGA3v
f1x9fBSLkvvE8mB6DIOCPtO7JGEdz7pSs/+yEWr6sMOEBZ0p6hsgb7W3gsao
YhaH2gPT/jfBpyjADb+vYDUI2JlprEtWqJICAIL+zpmcQGSaYb6N7vkmQcFo
z9rWqEaOg9pnl30z8ypHtg00YGIa20ldpfRlucvG1n0R3OZMWv3HXxYQ7gy7
AsWwhp1/beiI4ya3M6OdYUhiDotsfHBwcDZSUn/scu/zRVX+2OkA6dm7qajx
aribxgEr1aNYnAe650pypH8xZZQdIqr9barjnBWzhNiXPxKVCxVsMwBhVwsW
xesXnBzXrqIu7m11nDGHAJL4vLv8fzsGJoBkVRNEJg1QUqfWAF7Kdl6r4QK4
K8ni0Sk9pYaHeAT6JFlu/ZRo/Bss9zVJfncw5VfP8cQ9riZxCIhGUhkmYGLv
LJs0SdEEyfHonZSk4XRA/8/DV8jsLAo6mUkIBlPvpqKf9aEi8ql39cpv845y
vk4dL3ZwxFBTycTvkFS2XQ2k7Cq/xVPcOTMCbGngjRK3LtujEiZiTIjq5q9I
5fSq9Y99i5EhSrFupkqidyJ/V6eQIEw0PF95FLRPdVz1skER6zs022botfFK
0QLUny672ELhRvohLPdn1i9xEa9ZrJ88yOKmjAI7yHIxx6f1or49ccg1nbIB
2xoIcH6SrIsn0QueNzMJpWHNcNYlREeV0LQijti9bgLXYAic6B1O4YG5+w7y
07KMS0AXUzVTrZokU/aQgjbBibGxTiHw1FHmdEg/EX3GI1KfkxK9g/whlmLs
YJrnaJUGC6MvGADGrEzO5Ok4gK4htypzofZW4omJSgvOAra6be16MfZv/A4l
o16rNUKUUrzEbWf+VUaxbpYQiCMuNvWBsiaNUqCvFHCTxsvL7Y12qJc7HyM8
53Xf12l9YHNOj7GqfvdQSsFgjia2ahuCJVSD8duPIb0YweewhmIuL/dVMUZJ
g/njX6hdOOuN/7DMfXvSxLuSuNvPWVW+gvuEHELM9XfLDKeAQBgga2rZqrOE
Y6m6LT4mknnk3rCDm+2FXyEk+BHBA8X2v951OJgLzQlPCRXju6u8TddL4kpS
ltX58JBmw7/nEA9jYuWx1NeueG1LPYWKT6weMH1TLG79F1PYX/OMeB2GcJjv
KTChlPNZYZ4kZRnofmTRK0yIfGVM1h+R77nmZF2X43ry+fsJ6Ls2/UNFWAz5
rPEhLWCZ1jtAU7YbChLTXygmrjBxIhVwANlvCvnb44RZtRFaYjpLKqSy+nYH
3lAZb2rQgzmd4b9P1aJBzUTSHgP1L7BCF4LwP7VCU/mi5UJrNFF/DBxRFaV+
zB0bA9OcR0zlqRYVEHi/Xd456mnGcrMkPisCBjwc6gFYHfwdPFl279WYaAEy
bk+ExHAEQmNcKfHbxRU+aHV07KnB0bb3mx8MGfOHn+yeCHdKXLYRBKV0VtE2
YSQuqA77T2eql/EYymTmSMNi5YMXEvB/oZ45bVQuijtib2OVxMHr7NFFiV86
Hr8Eze16kfi1HWo2+cIVVfKxgQ5kdeg7wnJF7WcJ7JDynO0F7hdVBrArZbBQ
SRT7fC4ZbkfaRa6+sCBLGbvH9kUfJ6ZzfEA3UbNE7X41GlN/JCl1kwUZEGkR
m+X/rAAVwLBgcJ5jshNA01Ao+maxdYlaXv+G91WeOwrw4GiVv1Ri3QMlvfqi
8/Y1rxVZOG0/t2iXNjCsj62eCxKuzv8v659LqyCDymiReNRliIsN7dT5FSN2
2s1KCKSchokIa+m3lXHwopDr7tlRYq2YM7wKakMcOCTBwZXirLDzt4CG4Tr5
nE3DLzbex4MS90Tt76MBEAV3bOVxSXDZvE/zral5+xLKI5p8QgFfqGtt1ugI
7aj4B41oeOlE9HuM3jO16BNgGe+LV9Gi7FU8SL0N0RsVTY75wq2Oi0PCekQx
Hhs9GCdxSJNZoBDqHvO24Z0zze5jpQTm5i+2Qcs4jQJH0LF6DUu9jEGB9I9G
Xh9rljVP0Vplpw78ujXjAORkOgDCsNa0687jCpHbCJD8dreefoliqTXRJxVv
Rh/SMUZlp8M+m+pN2pwluOUbALzxEXcUYTCyOLA4XpzKmByWFVKe4QFeGUtE
0z5QDhPfV0utFbCypGag5RxpMSwEnj942akCoDU7FTASHcW51F0lZNnjT8cM
o1ReI1tKmSFP04cRvZi3xts+wGzoXHIUNpQIpoDTDJsX94C+ou0YXONl75qE
21OvT/l/GYmOk6d49g93znh7xfsco31tRSfZyFhEfKK+7/GWY61/4+Rr+2lR
NtNmf9WaTvXU3Zy0Aoncriz00zPc7uMn3ovIwN+kwMvpdSkPjSofQ459bhEG
R7mKd8djE34Gb+WNvg3vOSMF2z86eqPGkAEwSwZQOhZYsSpIPS4yyRaeixsw
Ca8VMqbL9SVZnksRPkUYDxWqPLU8A+2Wnh/mlPrlJ5SRHeyI9LC209K4XN9d
/xBil6b5lW6ot5mCHGdAH2COAg19vyZSWFklciS7FY25CSVqcZV4lEqr6hxr
lVURazQRy0clqvkqctjvd515QU/K9Nvv1vDNdBT5OHMx20vmj+H2cLCJHKj2
9j7JdsKkjs3MXG9Kwyt1xdF68wSj4IGs1BtrThTwT1XwEx/LbtAozDyqBgWB
q2eQassukr5ky7MHwN12YVv+AUYB6y9FC2zGCRmRAGbZ5JQTOTHVB7Tc5WaC
OYZeOvHsqrqcJXydVisba6GB0voggJu1PkaJdmkA9q7IeHXBb2CheucOSxMO
nK7/JGmUhZu8sYu94QlBHzBSTAV6myT0ZbxgnhzpXiFlrw1+GSr19latdWDK
GJXX/ProUpK/VvTxlXGqKsS77iC9Ig95l2dVGNpkhwUfjMRyKIGqoJwhLkL5
u6wKKceRFLacWIKL7p6KyhWM6qfCzcSFRp0NDTmLw0w+d86tjN3smklqEebn
YCKURKYJ0QId5zw3orUAYjlNUmztrqNwWTZdAWFopw979+hFuBHjJlNKgrOT
UcRbEOco/12Z8Iwflv9dft5vZAJCmCyrIOgqTBrjopVfrTgyUurM3YzHd4Ye
SNHfS22y3QlM9rnn/FpxuVCNohrn4OkKL66sFrVcgv4+DUlCbJQJyib6Pr6n
LbLaajwvqMX3vlm/WoR0EMJP2IhSUBzWSns7SQ7khEN5e7DczkEVWltZ5w1O
2gckMSYuzitB4x6OjGqHg/ohOLOlZuyDWtusKZ9P0BzKzDL73fb0njG+/FoB
ayDXXyN2C2zCCz7NZXeCIsQily9+wDOxj41OUwEvzqikMR2dmy0TVfQJ/I3b
BaE/JlzNLE6VwPbQ22LsMAYrXpDv96NH4gFUlXvCi9Z54qSK4pt2jP8krndB
CbPy53KV26iMUCt76ok6ooN+7j6NM1mDC9xnXA1SCZsGt01NDzcnGuY1Iock
Mocm00IICGOkIkIfQYD3/NTaqjoSCT+N9ts1xbBhZckib+gSUusDbOmzzxdc
UjtxV589QH1B7WjNr8msNwRHl/K0KuSK3nqwpBw0XiCeaYgIfSbPtkRk4ZDa
mw7nWqYJ1odX3qR35NEKlenDO37nqIFl5SCkl0SXmn3MLzLUJUb29iI+53Fu
HXUi7BWDYqgunFj2zRIE8qNLvPmHxCKnGm2kp0/FCjWEuPG4PqcoMVr6rCgx
jeuS6be7pbWxCpzfksrND+B7fjmDM1UxTOZjcySFms2xgQKK0Fr+XUaujNlZ
EVW8afKQdwCwF1ysi+z3gO7CmPjP/+INfyTo90OQ2WHwCB7dDJj7Jk0Ab5kj
FNi8PtzLzslh5rlmY4WJrfd8yAtgNdf18U/h/OPXnTAXpx9NKTc92VVNlX6O
HQjrWx8qUhgDSslpUbiujeWBLpxLzm90Uwik99H3Y9uY+5w+vy5hlamWYPEo
3CcS/olZCUz44CJlEpKyN8bFKZOohJTLjXVIQQNEMOrhrwtljh6qSuELnqzh
QGKVTN+ypHa/L7xTgBYhkYx29kS8ZigL0D+TDxw/qSdXVg+fS3U5hKGY1Izm
ev2KkeMGL5qGm9MO6JIWmjszLGxp8EAFmjPARKgx6zVyl54gmjN4JJ7Oyg8K
vN4Xvk/2LMm++R1ZqTZShI3Hzq8eMk8IZQuRimv+NUvoSgAnXHpsJsRBmzv/
N3Gn3XPgK2wR9lVGiuNyWtNf9ofiOaP/+ZYFq2xp0Qw0QO48m5ildIboXM8B
g3IC99up76VuI9TQeOZ2eJuUM0lgt/1OJLFseS/YIKnjrGUia7KD0J9GZxBV
T+iLUVX4D9AEVI3pR8g/NXBcY454RUc+oL005DZhQY0abKlkkJQqyPeejgDz
z39jCxdCZ9x7/aWLJJyfb65kp08rP5o+S0XYV+i1tAR1J+P9bcAu1OaLtCBf
rbm01U3IiBYJlvOcIaLfH4hCj6KBqGHQwK89sczDyV9QCY+e2bvFygYHz7+m
N9boRT6Ge4FG67/vA/ZIkF9AZGYgL3kiv97MGUVGEISuUYGm536ra+utRBjA
/UtCFfxh8fQOYln8Vfs9HQMGkADX46hOEy6HOADn79lQGuNLFZlOT3U7gb5A
wWeLiagr37alKWRAcJkpBtiJWo/0sYYi7tSnTF8Zp9wBSvC3TEcjG3GzdvQg
mL4tWNDZqhY8uy6rqOxg9jsk4km2JLx048iQ6OmX5aPUcGHV84hvWhZ53VGS
7IPYRrW7HfxwKnCBZNj3uqkc5kJyNjziDlt2pPAu4p3ZdXAHJHxChl3NSFbI
iRssu3novcRqU2Rit4bYZCcLGmXUrPw6p4D9ga0iEE5iWc/mBROuusAiPydM
Aqs7HGcp0ATlV6L2yMFvTy3KyHFJqC2sjzMdG/rMrkWMa0unvc2QRrjUHFU9
tsR1HSRAwVh9I7wbPc5WTAwM1MA4A7sMt6DJ7p78KKHGAAO+4Ca1w4KRZJkK
xI150FyyEydCzrAi+nOlhHT30auolJD6t/8x409fyk1prbE8PIj+wRO0CV1u
3WONn+ZwCK5yonFnezeOvk0OZn2q0xNBihoOa+UaZM9QeiM+AevBGKCbogON
ZU7M5aHh25o0rVxechv0wl2FDum/vocP7eBqxHZl8dQbcFTqiU4GXUJoHSH6
qh/lj1UTB77rH5d3Rs3J18fW5eqNmsXK5eRxl1UHguxLYBSJMHQCWZdEj1tU
JWgohjlNPrB61vcxXrdbDC6F3TfwUcAk7F76N77ku7b8itzB/GS537eaNUIp
uWOy8YMBa4PIzQkYTV5Z2UT8txLQMdiCZ++oCGFw4qcZYxuhiIa79v3/aUAp
HOcuD2tP78VXq4KLD/SwjdtdD7rtAqf/hB5IkNUABA86UvHM0cA/HXujfM4I
nyNs7lbYF+B6xuWEwVRWKT0qCf98ofesuZWAFSlwh/2entBljV5bJb9Ukmq9
MZTnPbW5XxBD0lRsG7QH09ZG7tH0hl5yGztw5r2ykviSnMsRanHbWBGrlHZ1
vyZ2TsWOekZ29f0gKXteE3ZCoJzpejaocQ6pu7ysagFfNKlDlfUgOrQqwwE+
kR+JAggBQ2rmL26t7vCnwEtQKK2ZJc85ChB0sUAJQzzRVk/wEXPXo+H7sFUW
S+tnSGZkxLph+0mxpx6c8FdIcBB1Qp7nHi4NAuh2YRL2Z2v5VkNA+wxutQ1I
ZMRoVZzAyQ5kTeZLSX4wKOXDtRE6/zfCg0wrRD4ksQyl4SXx+UYC8eiyDrmx
o4ovGvX+WjG6W3SNtz+Q4xISDySgkm7qQJrA6mm+xyOzGxZYfObgn84GAi8u
yeDGjQOAlavmr67wzV9wx/+9m6R6JtXwyz3gN7rmwnKOyq8EHaE+0ewMWQir
+ho1Sihj+/o1hGkzaorGyJFoLnmEdUttgdVMhB+KHWZpWxr9mgVCW/G7+xVn
pivEaGs2SQuR0Hx/BLAFGE2u/flv/Ba03MK7g63BM0lI4bsUedK95tmKuCK6
3HHFmqetrzfLtkbzgi/aZFE3imLu8QXRDLRUcesfSEpQh+YSS8uyd7loqrD3
KCN3NhsP5/qYVhxQNM2/e+G2WOjY8j/4FGzUBmQVkr8ekg6QVYrrmNy6idtC
AS2nOztllFN9hxxGl6QL6NNlGEPNt4wUcHUwosCPv6S4YweCec7y/adpEwp8
s+wNX5JzDeI8YXBacl+prFWr7zvQljLbgcQkV++NBBSzLSuQN5CHLH0Tgutq
DOPSBHeuO+lVnk5g+6smtj3IHUbz7TvfzE8N+i2nbEVvZJWvFWQjQB0v/Id/
l2dy6LWdb0PKQKF4OybQTyi8YKM1ZnqaxZ5dlG04Ign5Md8S1uh7iit857G7
mAWCUivHvzyY3tD+VA2Sjptbcj7EfqPGsjbKaSa4KWtdnani80m9WzM0E5Rs
JO+RPQ/VvFIbo4KZFzrf6WbQW+mGu6CQTHSO9LnHFRu5o0e6W5BUiuPtPd1E
NiC2xhRkXM/O0GFqBF3xKviIeawxQ6iKueuqcmvsKaLdaGMUq0yebyTRMX4Z
dUjm05prl0OhoQHZ75UEhOxieZ3YqqnAUWvXk1ulxp6fKxSXCaYjN5sSUv5Y
3F7xVjSuGD1Ml5YRuVkqrGdJneDKx6KdWu06EQ/vP3vnNVPDzHIsBBfKQPFP
IOxWeA/D309hd1yMSv5v52UuS/f9bEzuWku6A9+H37ksqBE+lBnnzdWzhdp8
Ek5fQBMcXxdlztBp6yTYIOMB4kHiWckZvW5B72iBXepryP92XUX1PTjqUgtq
3KFvkwGqNfyqX2QRYyy/L5S0SJ7N31zbP7hcHIBVObW5cNdp0OB/Raff7veK
6RYZPHLgsDBOmfgdTDr5mg983hm1uVYTSpOxn0DQqNzZ0RvgS6BBgKOfDrbH
AgGfmafSRN/u6cP1/6DWzVR/0254f63E06W59Ctpv3Ot5J758SjEWHeNOUfr
nI4RkIKhjzAxUvR7YyHCtRfDLM6+/1IjzG0H1ajpM0PNfASkrdrvKwpDEk9k
4R4MpXkC90XuvKrT+PJ6PdeRA2liwryC2Y39FNjnmKXzhFpTHHpj8OiI7EAJ
6y9Tdy/NNHpAu6It5UqlTq00DT/HpN9IoCZS+tQbwgy3dXeyL+SCXVDnRVgG
nBFYiCVQP0u4BWYoOZYavVmRbM+Hq2mZgC4oDtJgjrsJpxbLAeydvrLet131
5IPVyavv7DCvSAPOSdc1vTyVAMEDQuu3kmepoRzK3Ca7+1hBZ9X/pcg1nPdM
Hi/TKzelepyQLmpwcACFVvKWUuOa0w6zw00iTLCdYiHlVI4U8P87K1OVwDyl
NSNAXUOYOI7owtkUrjAvqtKAsaGx0Ug+S4Z4GGQtm6k3XqM8DkSuGme8kNbF
kNQkTDuPNP3eZQqIE9yFZsV2NiHfZR3WVoxPp9x4BGOWj5QljaeBoTUaU457
+immS3RmsdxQbhM2yqoGR2hKMCyNxyrMc7kmVSF32UUSU2WP6sfRyOUJNoxQ
VSnbDm7B6zbt74UjPRHGTyjdK1W34Q58slUAwcoOIOTxlhPfpAFXEL2VAAtf
ZsxisckvFnPU0s1ikfHWwl+EMXyZzEwE9HNcCPc+R22IHsog4/o7SmODlcfP
86y4Ia9zzNPegT3qYeWZ88ISAZumiwc09vgHym8X8u9E9/LtCqBP+TtEDL8f
aRcmld23DlN4juWaGKKkWO3oTnR8Zsm9URUM/yBWHxxY89RhNEfmfp+0LsIF
VoMcrOmMGKow1wfVHFWPlJEx4JtJVasR6izoIcopYgDK7lhW3W4rGXd2jqPS
GyGKQrAYPfJ8/M9/b7bVbM89+wZPQ/2J1vA/K2W69jG29BRMb5cPTDdhPteg
NPXKMz7qJkVIQUojn4QIOhbS4lh9BY5t5VF14MBMqbva1n7ycMlNSV6XjRcN
bj76WrTsLAiWmu+cafhSFzIAv/IxwXNFUHW6YkpxwrPhKnwrdl+q3D8xiOJN
aA9Y8yh4l8gcI/ZnN/7GDvANjV+xT5wJOtJxQByDrbMthaKyzwdH/evdQQ0D
HRbSzDblvy+2uwYfBnTaz20f8LSjoLdqCiYuPvk8mpHIHLlm6sxZzwjU5bJ6
5WgSDspGeSuykmc8Zzd8Ho04YhG8yZpHIhTN5ef2EGqlktJXephlaVYjdLN5
4M8GX5PRo+7hau+IzCOQUXBufbE+bhnEVrW8o14QGIxBeF2G9Z5h5l7gv0n0
WpKa25tWOYweMNpfrJ9zLWtaBkU7FNXNmiqkqlFXe42L+uYg6FJVFl/6M/Kb
UIshpG6Bw3qgS3Rsu53j9K0MR6HTKwLHM176KVZkbhXJ2LDSW8cJ4RDUutIR
FVmHH7I1VZotvwZzkvVruGhQEMfLMIeIBLYMlBxLBhFSj6+gsRhaiZGK6VHn
jPs4acHjnPV4TngsZUfLxvsnJka5kFpxQIUNfCQg6FKIGa8y2p4AavQIle34
YHS+0oh6617nAOgT9ZwkRk2hJCMChPHNJObOirR7TES7YpPjiq1zEnxfp9bA
98AJjoNhkrsFIMupW7F11Ehivyf+84OgTXzYSVdS+hb99236vKInJ//bmTlj
mZYCpVu0dq+32IF02iSVmIHsnrZPzEWyjKXqu+3/kYekcv5CX4iz54vFOYFU
n2/lmnSsrQfVxUm9y/N7Wg+7Z6msNQY1LL1a2lSVsEG7OPyFddEKaAw4uNoo
0s+dUgg3e0Z/gQ3YxuiYNPI51FE5GCloii5R3e+Wj1MHOD0PtFGFxim66qoW
N8Ismin0VIwPFU+ybUW3Mt0N0Jet+PnPjdW7fgkbUrdBBNR2N0+g9S3coDSH
hhDGe7eSdZGqWG++h+sJPA9q37P1LiS+9WLY/iZ5sxDjwClGiWLuOWj4ed3n
lyJOwBdVoq8fjEoFkl4k7XeD5aM6VhMTo9Y0xre+ozBG2igxBBD7T4Ic4QAH
wHY64pg20DJ/TB6VXu4h6hl9RMwi16kKSCgNPZrcml5f0Hg7jc/ycYtykCOA
lfSmrtg6LU2xhhO7mySwxadjjCZ6+Zc/fU46KO9N+TlVsC626Jd7n6kwYz43
xccfwTaCLZyjqP/Gx30zc3RNtTh0RPqCsfm5h770vxhotQQZtr1FGCsys6g9
96MnFZHli3IXU9XpI+/7FgMyCa1PTvMZctqELHYbgS56Cs7UDMO7fBKtUX9X
THhL+7Oils/QhdozNAmCTki9HTdEuxloq7199smk/+rD5deBd6xmHyQnN4Eb
CsO8eZKZV75kqg7v91jEpt9cZTyESpOIgZlcltJBQprp/x4XZyS0Rq3NbOBJ
xR+3gv2/qty+A59tr+//Qv51ARcGIo5YlK+nvnTxGmRuc2EMzcYQGR+gWI9+
XRFjSf+uhLMmM7boa4YRXzzVi2orVl4/E49Wfk0uDhXuejgZYCj202KSHHX4
D4P9DeyJcw+sPukKhkwi6MSkmW9LW1LlBKEqIaBVN7Mo7TY3rermSun1j/wR
mL+oCaXWkqqjF71wYYG3ATvw7AF5qve1uZ9SL7JYLJyrWwPxgiH+TFF12Lzq
Pe52b++InlZ8Ug1xcDJXM3wpH8KxzHmggE27D9rYv4oNdvVzDcWbiR+ow8Zl
BshkSsJAE86hii7afI8SF77wfa0ZgY2x+zlJlqd0e3p1BByWiOTaqLkHVanx
FHe0YoBSUPBP6hTM5G8r1twoReU/SzUUuxtYO7rKsj7HJ6MXB0kg86WSioTb
oR3CRLdqased/Ta2tAzdQzP3gtYyAm17GQA6UJL1EOPCpdlVxn8MKZrPAqX8
PVogPtSsq/54589bFdszZAOS1F+ivjDjx3LXM3m/ljMnf/+qKIBJTtAHhVrS
7UcSiwuvyIluITJI1Ve/51Da/hBFrw8mOZn8e3qvhyGFESjiJXjJjort3B2S
URZMDXNdXYnaaqIO5v91CpvkCUr1E/CyGJZv3hwR7y0TyURs0dtfH7t555ZU
ikNTz2vxm9u4Go34ijjPGe+P+CImPJQ45FNxGbv6RtcpnYWb9QCTvQBVALao
7JIHwBqoSzhSHzvA/8A6RIQFsgMo2YHgM5E/lpKkDtsdcwO4hz5P89sq1dhE
mEKzS4eh2s7g3F88TWFn2mFrcQvfmrlgTaqHzHICaH8qP8N+PZzVBxbZWlaG
gxy6rqFCn2vrS5+mTJKTpzkmj092z/K1fVVSdcfgzR6/smyTwKrArI6RizT3
01fgcdo8ijjMS/aSBtV9xPt7gC9FwMXSMK6NPkqPGj/CBhisVuxvBQTrkSFt
n3daK4Xr4dfsUq1EO0l85JGsnPdQg19KVgijOMkWU0c+PRt2/ExD22Umtk2X
BLqoDYjyscLoBjkFiYT7VmV7/fXRl3nD2++TGXmUoBylCWpgZXiGhsyj3/6Q
hXi8QkBQCpX+jNoT4O38zMqXZwbNbgbx1Lwq+ineGjNfJRsztNRTXFdvuTkB
RvtmlBjtn2wc69Yw9mDy0rKrLs6/XWf61KX/e6ZqS/zl5JlnlV3kcUHmB2Xx
U5a29fyii35hkpjFVNoeNYl1rF1FWy8omIM5S8dFNNZKUKEVmRwsDOFqWteo
tjyGPBTpACabFmFOU6nQJgAqiyxvtfOZiz+gmyDMHYlNguYzb86CeZ23YHpc
iEC04w2ZinR+9bq0FExnCqhJqKojz0dr71HnWhskUcs7UFQQiopObyBoN+0m
lCctU4xj89iq9LiW1mJY/ABH1ZPdWtSVldwAEcTevNSxRSHa77TWE+bzKxJj
Ydth0JU/+awHMmlZ0+gwUGxBgzPW25zhT9rampNXH670atTTbzIVjRCnckNh
HPFWqHD4OCK26FLrT1I30AWGWjWno53kA30VKsAAQ9Fw//L1tzGJVwkGxXwJ
SJCIB3hZYoxABltN2Zd1Y3+TWxM0U129ex3AzQrHeaIElT2tRHezM/sK6pR7
g1tl7vK+TT8uiWQD2iKGlymT4g8WWTzjt3E/HUB5j9DgAbXHG3T4DEfQqzM5
iEA/hrjCRry7PlnWSlg8c7s/FxxW8bKp1WyBAMq0nQCBnj7J191oiJhtvFp2
0rHkkkyWnDizOTtLWhTmxLzOyGJG8EBwYmbdASJrM1489/k6YOeHDi4zoFSt
Jzb7AkCPaxhQcqhx+YO/OwU2zZq0oW76do63fIlPuIjpi+MCsqZQG8BiikaJ
5+eJMzXTgOgTPVhu7WiEPEmNZWkEPYugCRepyMghz1G4C7IEByJ077+iq28U
C4VBTl9tj3M4TP/6ugv/Tz0PiV3miZduocPAPTTHKkc7JnMsi3LAh15AVpCI
SP60Ax1DaobOkVzDMmeKNdpX3os7egWHRLAS8A+q8AePazoXc2GRzJcGR1cb
BDR4U9EOPIZgnJY7B7KixsqFh5mVqKnUdcVPgr7ml1qM2DTMC1aIITMzc4BL
LGyKVrHOr2XBTlHLtvlHPZ09YGqL7jtkKfJlZ6XQd+1NlpatCjsOWc0+2MPD
2l75vO2mZAXCl+UK0YGj3jd+iJ1aA3hlVJrqHel/BNrpLGEBL2cwxtSOK7SO
NykKBvvAv8MxTHPZ9puCmsTbMjtJFaQMLAjFIZN94AYmFUDs400du0HS2t0w
xqe/4/zdl3/WlXtTDFNMOdNxsTpM3WkOOMA4PjKAn5oykpt4H2+ZXFw+xri3
u/kLX45rB4wAdZsKUDnlHM/NRXpsD52sH933/9Z90VVM+EMQXxmM9riwsh48
VLNx7TzypYk8fE3APX7FjFWlg1JmfyRufEOzhW3Cp5NrPBf7lazvHuz1utzP
J2c46pr4Gw2TFPwOqzDkZf3EDeiEOPJ/qwhg4mE4IJSd9j447sd/sTSbEwY2
8DOVWbF2bYhwgFgaB1KqeTDrKFJ3/84WZ1fHuCXco5+gyCYMVzjBPvm6A7at
ZgTqJrPQxChYkw2Aj0u8IvzniNwuzpJGGI22Zdanyj1WkiwO3wkb/lKHJCvT
laUjI5TSJI8i7NLv9TWWioJWQ+Kv1MfAaLnLkCUhGNK4lCLqOks5cbZC/HOz
AAKbHlrw9R7CtbLScjNt/jhDWJcnJ88ONjFA1OEuedk9AcTn2Kw91BoSjknX
SA4fsmELrGztW8mJ4x4ArwtrtfCnREE5+KfmVohZMYZaOVsY8ldHlevzOGCM
7mgeF2ioOAa/XkpOvO9jpQ9qa4mPf+hqRa2lGAulALZCcmhcFTadL+v0oaDj
cHfBN/Eq7CRA66UyotxuzS8URhjPv3M8nZaGtFMPW7e0ggPXSwe/A3IQWUEI
D6JZR7SKSAO3hUhRy9BnUEwzzlC9nrul4rjLs2xCCAw2SeJOMn1bf50yI3bR
gJJFw2ummOb/HsNFkMaRr1RUqIc6WsCeNs+/lLiO5a+1t4hmRPLfWkjjeV8k
ypE73myjF8DyC15xdeWXU841eUfEthY4IBQQLULjHCk8de0pwA98XttKukj9
KwIBx4m6dkME3fTxiGIefe9phGCzHntOklVs5CbB1hHJD9l7+RuWbAJzZ2d1
WHzpDLK/xRYBYoOG355YC3ScEBYylw7yZ48Amt7+OLbPl82kqZ7vR0xiCAiv
Gko1ogGXc3oKhzND9AiIR3qJrhOfWv1CxBsr35PmO5Qgzn8oiX0VcWi7lGeN
IYfjdnIgNjDhLPWM8QnLs757t6qvLHYdl3gZjT8ZonXsk/jqNzmrvWXpI+Rw
LJpw7XSNa+wFUsO7RJBd6TJlWvNGtjpxJvwg3/ebRceRveOBvYOgiWCzrew7
60X1k9l8KFrkJPApneb2NleN8Ab3asWoVjt1bn0ugfdIIaxOupl4lf+Eqsri
1/ftZa+WFE2F/ajWswWq2c7FW1VbfVUonsEvipmHSIjxLNulEhv2x13mh0XO
l42TQF9LrY+jdeY4jNKCw6KwvEFCLoUYD0oWaBrXSq5ewwqmgScmEgTgxUbz
glK+6o572ojzMQi4jkqlFnf87qsFOyKTB7Mudon4XPZLrBLwXIQ7wLbEYEoF
a17/wWECwII13wIMbmDbrixEvIvNUuzKndPxPRiFvmK1vkpckBiZ1V8Etakj
OfxalVOHvgMM2wesF6l+urLgW833J+2uDmAg4gFsVShgG0qur7y1rKuChg1o
xjGaMMZ4FRz687ogLLlygCKBjAypyBxrgD4pPKqZZoTHrFDZ+aICjOLdEnJA
CTaKmndZ5pMlG9g1bfivFMDxmA2zqhCxi43J52LBt+DLTnTF8xGgyIXoBjYM
GX5Eq30H2KCnPiqqzIK5Vq+pksMuYmVi5iPN7AD2RBGmQ1LWHSYU58wZLjZD
wP1Y0YfWUboTOQgAWvrCVYdVUnGoLfOYZ3gdNhHPiW6X9y4fWTWaBG1kBSNw
9YgswEXYQ/7OH8AKBPELub76wZKAeiWsGcGqAVimmWRMWUULbxS4Ix9B2s4L
7zJfOgS+6Pr2nq58wRE/tpTO41NJabPYlLEwclivQ70k3/ejjUXPET5V9UTM
dTYTTmHmdyRt0jGGbZGeWSIZNU8n9kxD0YDbXy4XTx8MzUZtA0ouobkH6twD
wSPJq4wKvd8GutQ9IybNSJB8SQhq476H6ZdWtWTVd/aEcl6XbfO7tsblFadC
BIpmDZSKIlDm70u7Lq/P1kHArYgv7wHXbBnp43Z/KnwCLVZDouNChrHxsCZU
S0aoR71XJif1SPxRoEySiiamelaY6D9mpVbv1oEZvVRmAtcWCkkntmF7KGKT
TgyYb72zCVH3Zxm8n681MOq7A0lLKI4oEX8rGuuDVkJ1rO/X+eZYzczv1Ulr
/lsX0Tn1Hvj0hwdvNWjQDzS2VBt4lvMCRPaIkVtwlfUOYeqTd5OqMF2Sf5oH
UZU4Uer7f5774+JzOlw2xFCQ6jFnFzw1trgobOLClE1FyKUBDYXVk3mJn0dd
nSiMElxTO9bx88kyF9mYxVfny5IITjIBvIfMeZPR+in1ilPgW0wbJ4NCZgij
u2llBPy5RRNKgk1nS62rLue7K1Pcrersl/Femix4I/JxuxXJXvSWkdRBkD/b
ts8Edp7pmEstcrcezXMRjpXRMYmYy+MxLp62gpgL4oTIpbYSA9nYbpd0/Eii
od6lHBLoriobFT06Dqdhu23sO7bIGH0Y5p49cgVA///KgttzwEACkxPrx0xp
WCmKq2cGAmxTfCoLRHcfBGztjvbxD7+4r+l7IFERq+XiLlVgA6UCuZuOG077
fg01aZafx/pnSPAvzJkr0erJZBeAeabm/9ISFc1H/X0Qjg82MDwppRm7Ni/5
SL9SAV06nTLVrf8lt4Hatz86xs17zdiQQtK+O4mIC8N5Oqm+8h/PrKyUldRJ
cKoHR3o4x/yqTCY3+91T1S5JeRpkhEY44LWms6EY2j9+irYgQBZGGGbfgYjl
Sq5L1ECe0wdB00Tqb5ZnMl9R6iRRwPrPQLo8ckZcWjoks2B+btqwWvVDVtyi
uYIOtcyqEaaW0XA4JjvXegZfoyjct/wWSaT2/TZXw/3VLi0B0mvsVg+AmO9b
+9sl1xMfeZwUcAEXRsSJXjRxL7kwdySRw9be3QyngSiq7bkp7SMxsVE6yyhB
axH8q5+LRGk0xWVijG8CuBDuOzXAfvqFt7YYlbf36rTHia4gpsic8T6b5pTb
ObAwtMgTt5CEXaXpCBNWCAPKAIAoOfh2V2Lgo28Tup+6q6357WJYwWbfx6dY
lj7ZHxsywyh5iKcmQTcdpe7Nw8orpp4lug/cXjmpFB/A2zkAMgRaTCWswq7T
p3F7TOXRJDJKntmnotDifs7oZ3giX6hwNhV50UzbeBHxWtcadADyxolUg59R
SdoqZMjs0pGhm8fzKXZV3BnvDBzyY/xKSMg8TIXZip8TPKwLCX/vOOIdxt7H
658FCEDe2WoPyROwuIPSikSGSYRPubLL7P+WO535a2G1yXjhx3BSRgRSY9Vn
FVPAKFX0BlG9ubiGL/PCV750rAT8gDPEU99XNDhiVJSEs0EJ2CMfP2+Bffo0
kSWnadr/jSGRV12M/86sLAM1KlnbK2WeFUGxv6YpLleLWQQVskSqMfGQHB8B
cv1TFk27pMWxdRxp76nvk4AnKx7XQsla/nWuy0OK8t21Naz8k53FEBD/wVAo
yl+/YMqmDu6OhXkTaOq8J1sSdYFJqao8OXJMy7cLEO+jedYhVD7oLgaFFess
BeHUx5weazUfF4OYlViHTrkUBA9abcBlTjzZVf5VzAEL2YaUzLhbw8I+9ZWf
E3cWfGwl0Y/L6xY9Kday7iysKq+46tIcZe0XMi02jWDuXg8krhZcDli16YFr
3PljO9x4XkaFT7zqnX6TytAO2jU7dokBFaIZWfnzaZvj6/0avtHT499tjG08
VHQTafMLdGf9aLEfRiMZSjvoFAOVlX4U7CF0aLZHtmclWBjXb3yDFBnYxIGV
6z9s8OyIHxtxicWVnn67zU+HBWgdaud+XsavP6LurBdN+LPWwmIlocRwdFc0
spKMbv51OOZskbO1R/tXRUtskPMS5xVZg2ewNZvrFSskedrlBsNTuQtbjd7X
T651NlteuK75jkGHWKRPfs1l0R0C/tnjUZbauDPCcUK7hPG6iRQQsL0PB7RU
hKo3SEnSM0fI0h4ozsZIQMsKprbFAw/BSM/4sxOc0A/Clvcs5MOupEZjygfp
tFBVqwGDSXmSbwQj458/AUJrmJMllsOzzxkyqBrBd9WY/p56VjVYgYX0pERl
cpuVDA/zS8j2KSe6Ssh6NLUrBzMC6XUyk9T6gnq8V07pRTXuBZOmDyzeZRQn
x7VkuF0iFgmtfxNmvy0yF+QVw4aZq1J6uuRgB4I+69WiG4A4nRcO4iEJtoJb
bJ84xjALMbz+ZvgKf1ny+TP88oSzm3d5VRA747TodzsIp8m+5kxukxtSc3Lf
AubeLNB35424iTbM/UJU+2z6XnNvQEUtydgX/UlV+E/3t9Gk3nJWnfT/VW5L
yc3GyfQq/WLAspQcbPoxMCR+oGkI6Xj4EdouRLSgwnQGPtl2fBVY4KMn9Ffv
vTencMUyyWALOl8vA6/AyufK5ExQew9dz+2tXdQKOB8dgOGE7SKxBG8Lqk4u
VBsqe1BRs05rQUIytK6so4AW5kE1z+I0hhreRcOFPvYfn7POUlc3cJW9ZFjb
NYpfh6fg4TKxw0lUWMxwPUh2xi/gDTBWcpz9cZkB0oLNEEMe2FWpbzeXHqty
CDrqX6dYRXMwK67nAM2Fypv132RjCco0NQB1g32kI5fh1jlbgAkdF0/MyPuC
HyLKM/CTbC3VbH52JxwEQj5KECBSb3DEegDE/CfUtXygB++0ugVf+sL5Jykf
3ca2juIWE5/tQbkdqgQuNIcqWnfF2oF6iwNMBxDnaTvUaOsPLryyBrLgt6BM
H2T+VKKemP1uqRvDSPwp0sWTgNzY3RE4OXONaHybsQCsJJKd/KCv0Dv8gkcv
et939MDXJ3RdRFgI0Zh4Bt0UUOSJrmuO/34QfHb8jvN/mPFmNkxsP9ySUkQ1
dP2k5nfRWW8oZkzp8IpP2Y4mn33Hug7qNtGU5rAcja96atwDzKTW0x8qtB4p
O0JIA5kpVf4DwvR39A3A8eu/x76Cdxmwogmgi4SZDeJ/gThH7jOqvsyW6hJP
7aJDQQ0drDa/1kjkipPoQKltxJbZTgdhW6ijmb4xizPBAyBCir4TcZCmCD9z
cXtv1qfIRrNJswfsHPS0i4rVVnbV3muSRStRx4YB9t5rTYm21MaZCwIy3w/c
XHIcfuVoP6/oZo+clBSuuSqks6YG9KotRyh4aetXZYIEaJiFSP4xjKPjG1qH
KS1PDjPZjm+XBrFPGrYOR5/U6CWTXnw4zD2d8EfBW42+00dAaXpiy7VLGOLz
B3wf06ZKgkFtlusvTxusN6VBhl9rkhri//V9XBHcJBFFzjhQwQ7rsD6dH/lf
Kq/VNDqrTQgAP7ei3e3VSWtoAkWWH7Ae0fJjqMBKyJETJQzab/z3+yzT+8Pi
mJRBUwWkUB53jkZy3ivPFR7ixWnuDUZJAU3rO0NBjvftBUqEpqPonS3P0whA
yAdsdgoWYLPbnHYi+TvMETLoVrp6wjn7mmdxnhdRqwClGmf5N6bX0GkpWz+d
c7rhqCv8NUYPCMwgEmEaeL1GV+qtzHSlX5uLWll157B1CvguhIEsSJpfqvQr
D3hwmQv/QnhCa+oz2/1+DM9Y6m5c0v31aySkM7dtA7kDiKDsxSPY0ikVD3uJ
5FmZovtdT7ddLsiOOG9B7AF+SQBqfGRMWDKDk+udYG4Ab8fVPJOC+BzQVxIr
ncSWw9ts2lnP+HZM772F2E4uL2LEQHkKrEYlvzxQgBFWFscTruprXkOHbIal
U2lHrI1VY37ty2JX64xFqii5zZ27txsQbQPVTwwJctzBiXdKHqtYVb0XPWL5
0yey3Lcps5+tKYKAIszZIxlRcbapU1Q6LDOCVJy2rkMAYmMm8epO1hXCqAcD
fttwuqw8sqq22wAGL+5Uqes4/cgFjUxLDFzUkK9zSVXlv7vkip5GXvf/Lonr
ZfczqFBIkRye7DxBEzCpJSbQiJgP/Mqh+bXiH5HO7amRJWY/uS1j48M+URMR
e1GFgYGzbmNfcJZ3OTGKylqWanc3XO0YFdAdEZa3KVkEVgSONkXeEAi4Dj1W
yGRTXtgutmWH2MoYMSQ38looMg7sp9sxbaxR110IW2NDApnakg2untWDn6rV
kVuebRMD6Q3mZm3oHHnZtcYacDpjOwOtxxh/q2TMldLWcVlRJF/+noPVj6nD
AFY4uqpKCLdqsP9ZGRP1xRqjQlxNmTGP6N5T6uP/m8u/lYDjNmWLy+/tDBcF
v2rF8Xgomv/DBecxakw1rPTpxHi5P6RWfI7kmpF931tO5YuJo8Yd8eXSxNPB
d0QbTwPG+dt8bzJsX6RmHgXne7ioU23YDmpTzOH0xbvBiTHiY26Suedd1lEB
qRYK9WTyYvYADwgBLTrF5pA2oH8lflTk2ErdKsQodQs/m3ynHEP8ipCp/zBK
gf3dr3DBitYaMwXa5ZKJbk1XkAhRGfoKHXdl2mOwq+NXXv8ltd1BJEAqX6vf
JORp+k1VY2GbS8/ScbZ/Jfe+UwVwW/9MYzHUWGEp9hv5FbeNME6VTQU45XuE
GPCR8LMh9oue47pRMUo4K8hyxqfIVYqNoUof8MMyW3u7WRPL25bIAIS9tn6h
5276nkXfA/XZsjdqTp91/YhvjCbLP4IcbXhvsEz3P8/FA2LYcMGALGzthNjd
68spz7OJnIxWQKo+AU6izvoOWjB6l6D+U1IG9aJo+9fKJRotmnoTEYUDv/oj
dAYfai+iGtfIoBfsRhBVjXh/JvzZzzuLUDi+3ArXUqXIZSTJWMa3SQJ/b/PF
UDNiAEEP1aXTciVcbzqzzoj6mZh6yhWSis/jT+qfSX7S3BcQyz5iMs8XFGSB
ZRYbiPSMXNWlAoW+Ki10okQa54OJ/gkXJGZjZSAMuA74Pp8SmoAIIlAVB8fH
DVL2PeDQODaWmAO9zNY7TH40HOI/AKk7L/61psTWJwVcW8rVfKHrT56mcd96
+y23jko7qUVKt0q8RfOMz5i0RW2n8Hhy8R28i2JlcAAbFSH7Z6duPvmCcNMz
bZYJA3z9K1TVc364zhDyD1JkaTFzAS5e6NqCELx/6Va14k+QdFucYIJDf6hM
bJv7eMo+PQLmd8sT3ndx0+mV0AUoDU2HICVN5mkkaPGjw0FUsRiq1B/QL27c
NoT6+VFPGCvXDz0m5K7Uy8SodnMBcLEQxQ1Lok7tPOtmPO12L3vrEDL4KMwV
gfgsJK+BTx3nz6WqaGhrDcCHUHOSErtukl+eNs3T2w16JA6MCY9UxGe6Ak9l
TZMOy3kzwyuMlldYh1xOPQVABL1OIg/PPWOeMxaqq92wMRHm4ZXFaRvaXGg+
k/T3tm03Qf3hmOtY97y+/W9ewgmuel/h24f++p/+hWdY8ytxp0Fb4Edn7YQK
jizAZjJ7jpEttiUfOgUbmafRWf5VljHC1bqMwpWUezcirYrfdic5gsHnmHR/
59MWt5yztDIT9v7xCRPXsELMyDodQSoQnV4OzyGuQhroj9fPeOEhX8iIVmB2
6kBh+n+OSMtjQSv/iz99z5cWyUSH+mypioVLNAeMvs1trE9zOairtO/LIllP
oztSWZgcI639dz3tSuvgEbnB/qKWnQUcswUlcxGZiDrLLqPAB+mJ4U7uznIH
O2eRmUOreHgIyrTyV3E1xFT1pVwEiBj7L1OwGwUd4xKk3sNkvXAhVhjuWcsh
o3KxBA8iMzqBhg+GGzkgGBkmkR19Dq5OZcyepvMWBHhmBCe4ptnqB5RY8wtM
CqRbnpcPTmGNpkYCOV1ZAuI6h4p47TZlrXuCBmKKmla9Hi2++HhOAwPuzLg5
qXfjirWLDuSwPT4G6hN+kofCbFDdhj1isysdKPh5PZBWviYgvc5n/5GFcdLl
97jS/pv2S6tjpc7CZbdd6R7tA3yf1tMh6THd3+G3iB992mwgYb9ClHCklTsg
shgEIA0MKAQo1uNKO9ol26Pn272TuLF+UI7sFCIsyEN/O7pGyBFYsiopdlXJ
uCv98Tmagsip9qhqg9zviudBp4CGHT5W6QkfCgmjXJRqG8LUemcJB9gJhvpD
GPp48Cbqw0K0gFffeKWIP+BEPsVqI7xjhXSau3M9+/51RJYmcYsE9bjw4gOc
fl+ZEy4K7J0VTlCmckE5eGGDu7F+9ybCrACfKByIFUlzdALVx1AW5X5dw+un
W0u73kndzXJ/pFj9frH2C8pm3u0HmoAS2T9tPJdaGAh0J/F6nXGHMM3pwEwa
aeoZzkjDFZsTxpDjEmtrMUw/X9X50qA7+ugKMQJ12f2cv++GDzg95+RatW21
FyGbKA/yZcjtmuPLTEhMg5qOUOe3mHWRU1v/LJ1UfSdLqHo8+rijC8wiwrA8
OtO/SCwPTIHDWzaMKaJQ9F/sN1o8qn5AHsj74iE/R2UJrDWVMQpo6VsHjYOI
4KQ+yFqRVfWpCMc/RwnRYZjTfjIecMUpxz5v3YYNJAiYwqyGV2g47iYRcdai
E8v3PXj9n7qnY6neAHKq7ug506z9MDo7JgMT69J/AyBf9KRbaMWR64N+EvGT
/GsuwBjIR07TtAHZB5Zj4fSk2dHIugGNYfk8Jwum+QyHCmTsMPS45IpFiG04
8B4cPMoovab+arJyESD9qye7HgQa0VAP1Qn+lAKkPhzSolr5TQoka8RnVQWx
LUIDw6l4MgA87Qa/Kb46Idd1sk4v3G9Gufd81ZZ5eRpYqcw6Akb17YJxC7Ri
AKgt7xTCYek+Wm7j0wcJZUGvYlcrmFIPAn1Ge5HVLvpfkWAMLdrHIMj+XxBA
nHZL7xvEPWAY7AQcvD/W5JTk50b0hByheSAFCIfN3QJkN4n0p3mmNWwtLmnF
0ihqJ2+ER37W9WPJvSQ0zJpjIBjYiHzujd0j5Z/94mynea6lompS5CWGJ+W0
L9vUA1bgwUPX5vsfpdPkMgE1D59nqDTp+gp39ETRESiVL48k034iZmpVTVeJ
K7tq+r7r+p2lhvWO5cyChWw88aEE4er6Jh1bpmv8OnXeDrdNJj13xu02xTrp
mPHpIAj9Ieh7tfS/Kpe59ECEhgjKiZGEF+9ANbcL5wQvpgoPlT+rnJhzZlAW
lY7ZxdwYs3DvBOlLF/vz4iIvdPnsRtauY4F9imKJ25WalDOecusyqFx73tmF
Dt4t4tbqWiQ6zIz6I8N6fxfdAfIogrRWz8gBwQIFYpquqs4qB7kSxrXYVWaI
b2RXUrmt9LLQ6HpHHVAJYhHK7/u6ntH2wof3cUBBuDC9akrdhZ8BskZjtDfn
k3DJ8rdTwsso+31/0162o7PIGgvSkekb+Dnqyd+xSM36u3HNxwXvWwiY0Cf2
//AhRXK+XfWVLBX73pcsDHgSCkVzNyF7QT77H74vnTTqqEMOwuNPliyQcHfG
TgKHU9/yYg9xSCrMyf6t8jIVzevwdJDDqzwWscMVdTx6GlSbYsuPec9q3yZG
qaiNx4kt8fH7LUTqYDEx8CQqHGOwV32z6uWBpdnyTu7m1fdmpir9oDVfJ3JY
NNciDpowVHbjtJ56n/0SKiafZFcBwu8TUVsjoKEfgSmwXrJMF1Uo4SUkr5Tn
Cra3cdR/IBO21/ZVYugYN4g3jVAmahD9prvMoxOkVaqDod82nMmvn+PwOeQL
QQuTXb0FNU/gk0vASEumxg4xWNkd3/0YJ0J3KCAVRtzz02GRK3dkWbk4AlCU
mnPItBKrzkNE0QdV8eSOLisTQvrfanb80cnQ4WyA5UuUp6cQ7cwjpNP5tNTA
Wh57WG5Tmi/U0MY/VzjainNQBliquB2khEJSyzquEM0KcKRBqwHIjUe8DA+v
eNTTGSoTzauhy0Y40Q1gdugpUK4FvSKtDwJMcKME7iweYU8yyuAUOdKAQxTS
Y/4qBIN3Ml0Gly0+zeDsyUNWUeWpxLaKC//ETr2wk6xk32HE/nA/pFlRh+dV
bJ4L5g79tOjoCiurnvHDClXaF1hUvCbyxbYLLdzAnV0lFWKh7hypmCcpFbRf
gdmZdZtSPlUg9OFKLJQmNoOjlCcA3NFnjOZDXi8nZFHMsYFfJCas1NmnDHk6
2li8aD9QN6GRI8WEVlpyb7qx/2fTpk2H1DIFjwlXnUTRhQkQNOTwaT/DUYGx
B6NHsF35z/X83fp2ylT5QQbmNuIa3IFXCcImssKMU1Yh/dBteG9dNws0XTxo
CmmSdCkSDigA1SBJ1xPc4S4Pfrx3b9iCrtJPWaqwPJURaXS7Sa5sgzYfV0vD
n21OiFGQKgVCxfHOvNQQ5IjfRU4OHm+nHrO3dmK6yAVI2daOKzDRgVidndwK
x55JbE7OzvSn4ECA+CQyNJFy7kecb4AAjUNJvw0h+TFOo8C87XmfS2KQ9A0O
UK/OgGaABriivPE4ToTEBh712TLo9exfy5QLIAO5rAsyzcRVs8HZLFuRd1fp
gi+/3NsITSQ5iOXrNqjrA/obfsg+nZyWZW4cMiospPepQk55fZvfXpngF+0X
aej0LcXYEm9+oLg29RQThqVjWtEHhe8EqB+2iN74ESAejOhVliUX/oVBsnSG
NOZyoIspn983xJHuO/tX9IvH+efIpyy1838s0eeWygtbdYSZXbOkviJ0+cvS
by2QEL2GCxa68SPvJk6NdiqABbOGGUvgV+DU4HEL3NxZkyBTk12Vv3Oxf+/N
GDHe3oJbbjh6dSZf2qH2mJ8/z9uhIawErRRVGVXJEKNKHmRxZOttjs36PnTZ
GzymV/51guXkrtNbLUWa+6J/ekQL4dn461wpU9xWGqqIYBkQU3Vr1sEXS6wK
zTxD6nYN1gC3PYS6kONAcIPt1MrCM8O6leew38HRcd82oV3VccRtsxYXu8f6
VGiML2uaaQBkXC1IG5MRBnMRwEizLGOae+7Muxzvtg4mRJj3Fw39Ta9qBUwk
hxq/Oe5DSJN0t7VF/1J/MxYKRE+aZn6ALAKWOG/019Vg5ARpuEy6Cz6wYTie
QvlxBcNrYAnr25kyBn5KKBdTdmPNHCrnCyTsJ05JrF1B1BT7yBiG97gC9XAQ
SlbwGiASvoIN8jPdFjaYmaCkRnhjyYCkwGrux0Lus31KYgZ6KEzvBgZMwUre
MKrJdn3tAYR8qDmwekW6cKE3OQ73pmZ9bS/wL8I3kt7lDGCQz3klI+eHrjco
fN+ISpBITC0DhXBrQdzooz55dCJ4ZXoD7NM/URCzNaQeMutWpEN3TdGvndKa
wj1tuft6JsowhiVJ/GB4YE2f402M6nF47Uax3jGBtN5H73DR2Yll6Eok6kFF
g6aD/8oH9uOwAB4hw6xhXCP6mcx0MUcsIWipldFwdOZNzqkXeU5B6+idmIie
vmpms2OSY4eh3zmXGki3AOzwvLDoB1uBUANdwSIAL/A2bNDo5hGh+BDjZOnp
pTPNJ/behS4IsD744WGfUj82jP+V9i+gy9dv2mhQCKwiEzClpzkAOiy2f7gn
WOxmtz9/QrQZriVJte0Ge1xzZcVrwZJl04N1fixHpR8rTvvwzxoH5WP3hh2s
lr+Oe5SQ11bxwGkJVxH2BAa8i9NquKX8EyIRoLwD+7dIFL6VgKbIDCXU862M
kXPyrBe3f8R7QSWYgR0FdIcttmKBk13YuVARXbiFw9PUn+CU9ez3XRlaez+o
UlnyUMzbw/DCMYNHcIS3hVi6vG44LvxtXY2OFVVkHwfi+nkXzlaFjH+SULBe
QqBDWy046neG9MqeC21PWOKWhZNrQrOvsF0loaxmUWaLMl/a/Ih2gXJG4VVb
rN8V4JQ8P3nvsvB8RoclEy6c1L8mH53ZbVxMIDN5l9GIQQr8q6TUZ2cXr8Ky
fox3DxtxVIW7Q+g2lAIR+w2th11m7F3ELpuGndsljqG39Oe8fTgJUb6yrVZP
RDGPVBvh0oWEylGYsg/s3knL04KM8ndZWsCSd11vUeuihRUwO5yIKl8H70S/
XlpThS43Qkwvl2pjybTu5zcqGkNCLvud+IYg+ZFkqkS76Qz+e1iRWCX3HxGT
wpUtv+lXDSQ00+0vpZcC0ap8ahznfoGIghIty6ePyv4l8owyNmHxGlrz5QWs
X829KpBeZrYAllUJ6Emv8vM1/dtQ5/MqsSP1A6uwm8gdbRSkjr6yMkxi1HoS
PA3Z2WkBPTkZKW74XVPki78rpe1KqhaTK2JU5jcMBplU3/k1bSV9nBFaQEco
27mdVuJsjLVx+/1muISYXmFkfC/n2dW3VIQllqkcunD8ogPO/Xm+BkMr2rce
zjxiFLEGvum9XRcfIQS9/n2WqRF/fu/BghJxt+5H8V/cNv/vGWzOCphdXTGl
Gp33Kf48UNjSbylpBrJvK9hl4QemOyD9B9SyWNc9Trpjsz2GP4GmJuVrACMa
X8IIqqiY2j0sAG25BdgXPqQ0tEHt2DCBSldd0KTx1yfeOZ7s+z0DK7q2VsM1
6gq4TXtHaY96wcQXoy0mOTZRVuGZwNfAan+oUISwCqMY4e0Rxx4Q+XIdGWE3
vvFMXqP5BWC/yViyfuY77k318N0/14fYHE1/wH1mN+/5bmIAuPm/+uX18TcU
SZe9AH7xs7JbneeJl4hM5CVr7qZPMO3vKOVe/CsGbSrhRYhGTHerFswVA2LC
hzGoFS0ckAdlqpGp8JD/snymB4cW/rOBuY4bAAPrMTmXAaxVTFZIkgUyioYR
w9MvTo1gDRiFTmMY0bXq6e0Ae9WnTwsgu/54vkoFKettT7xC1kyidTetKH56
pVlGsCx9FEhTZyPHlW8xv2/1cMUMggsvtSiJSuyFDvJCpk6e/0CEYQ06CcVS
XnMPMMTGCgliyh/S7xr3O+DW8agcqGHmzz2LjFXl3p+8ri4aDRMzCFjLCIrm
LHWnroJOJfpV9i1qBADOO+KQPPrbjB5SgEEImC16tX9zPOuxN4z7xP16ULZ2
t3LgaVkI4MYOVJqyoUx3NqRrIj25EwuaJ8kwrcV6EBjCSisbzTNWMSWDtdMX
k/Y8zE+Icujw0U1pUgFqXEdsdYmpzt4aBSAJQtTMf8hOnHrPYL9NcFkAfdi4
MrhVL24kxygWPqc3v/8ciCqshYtWcK98lRrqq8OwOvGiooQWYNjbadNx2s0a
b2ha8LJn1kKdILTFG3WCO2aZv40fQj7I4B4Z7/1dmT/VaGrJRTXPWjNlzgZs
Szht7RQNNhUTOj1lE0gb9YpVDBa/QjKyR0/alOTZV+dmTE1RAxjiB58WgJP/
MJkJVCxAUKC/X0goWQ47voUxLKe3fHtZDj00wOEKIz91iJ2CJGFkUKHoxSjK
H8v8BUoMw2OMMEgmASl/LlY2mORSog7h/3x4Wtxt85fYm4XNSIIVTqTMM0g5
U0A50F5uVOgnnVKQQK81197Wku16tZ7tRzA9e3TJdw9SMFz0N3AiTtiD6U0o
5IWMQqdPHBKR/Vk5xGaRrM3na+TN10EwLPRcONRmx7vICa9KGog7yI460nza
JkjRTri8i38tTGyeP64kTwKtYloVNSMNVHGmS02NGeMgWnTRxlBxMUrklPnN
I8Dmua1dE3l1BQYUZH0R27cP76W/SkCSVDM+cif2+josUOBRJPI3fxWfj01P
PdBneoNDPZ8d92bxV+Ic1zI9AdMNNEHUmBPa8HAHEj9YPKP65zZvW2FUDahU
eFeqigQZ5YjK2x1AqBpYFrZSJYmu3g6LEUIDueh6n8AC3CBHSk0TMD21voGj
csJ02OymqaJ4JfyWu55S0oeYwQQbePrT3tmbBKczctYussD0CabYi87d0ng7
/So7bF3V/UdCZHTHgxegsi41+kYnVuFDpfkVIyHCgnFiOAcF+5kVTg4yQSjl
Gw2ABQqdRntyz81T6Su1u0wjofzigFnMbP3mJ48W6mb3PTPi2CTy1Cxpocrh
Pph2ObVASt2MDxw7bPdwcSWirr9P6FctazGas3Ze/cvfeTCfsKAd68NDDcSs
87HVMmSkG81nk6G/unaR1Ld31tFs7g/2WqtQh2TpbvGm+dtxKj/cedgU88qd
VJ5Kfp1awPv5FJlv+eXaqNoQ3ZlKctxG+ptnlEcSb6kQLWPtyitrylB2vJ5B
feleHBH7Qpr+LvrzkznDxr6lb7fJ1AqiHX/KGOn5CEyvhKGK8yMegGgZ5gLa
p/tGRNhK69BEH1YaaRBWrmP3nMs/KYegFe/pZllc1AWptLomUgSnmDVbG+WZ
swHMxUjiZ1I2YONGpaWRQ8JY1miNqmct5Kfk9WPyoLoVKOBBUMd3Q1oTulXN
2sh48Wx6XT4q0id6A748jscAEmFbccfOvVoaZj4lCrvPvox9kNUbJ3B7bv92
2iTYui8XveJLq9B3oAMtgyAbLKMyLyyHS/apU6Dora6fHlQ1UvkhxWpAstUy
UrEaHNvTCprBxB4E705hmL5IRWMBkIAYiEs4MMPq70FjJ9r16DvdBfC0sjv5
fdqzXhh9aaytNPWdmG7SJG+bZBn6kHlDygrvoTAiP+NQDMHNr8Tyfo4TfBwW
aqyYZTRGg6JMXoFcat1SjO+QlP09Q9DF3+KGOOM6/uAtGvL/uoOsj2OvxsOn
oPgCtJGYwJGtNwhRqjr6ndOXHubt382QRZpwGwle6xwqKjf90R0kzk44Ovbb
yRmG4ioG6RDlbgaEVQaOaCwZyUX2dmp1DgE1xzVzsOA0aet4nA3L7HR34aw+
aj7S5xzS495M27FFX+LbEi5G9GYGYH+AdATXLexLYWpfrks4cRnwjYIwZPmY
kjD3B05fEFdzr5afQi5j8b3qyHnOlt8pli1gV9i4n1SBm9t8jCPnxQR6YabP
3rkr2aaMtZtMcOpJ2+D0g4oHR5LQUK6U7rtAKrCCGbYgyYjUABNoeS42mBfr
59nLfwz9j00GIhMu3Y7S1W/sDcPSHkuor8A5PV/KynwMaa0Z9M0S2rCDa16U
nwpKH59mgi5NJNj5BW5Eb/Vu0yXacY0ZuFfQMtkrQK8TxLdw2eWV2jZBj+Ky
EoYyWIMoko74IyFLObR8qc2FGEqRiUeN09L6Vau+YxlbjSS9hVR+AG+i7NR7
dMGFua1lhoxYjJeAu3RevNTFH+6N+zbCxEoKQnf0fJYwqxLORGQDEAye5Vmi
7nuXky7O4ABAl+flBoUouHkVM7NleVX9om7D5z5eD8+waiHY2xnm+jibB/u1
gRWmU5432D2VF+P3Fc/c98ZDtIUk+HUXHdSOD90yjxHsfGUujKb5gDE9W4DA
ExjXgKFWy6/mILZsakvBtjKnMyNvr3lNOAvmVjUFdCE0Bap9EiZDVMKXtxnT
xckdZS7L2qJoeLG9QqdM2qV4/L1PuysSD42QKicpAAq76TJTkC0tHHf2ighz
1MbUMt7iQMeZNwf2d6t7K0Jp5ILH3lDRxJRomNU9ATHPVicjx7fEtGyudPfk
Ywd/Nj4QuF56BBVvP1Y0GV2HYJ1wyb2hzvPmtDgK6hDZL7CEXenbTlxdhFE2
8nFAErgoCscPjrHyhZyoV1wb3O2NffIsOcVkRuxL9EHRe+ZYW9sSWTB4Gu9m
ZBMlgbMBheWQORZSJSdFOLUeOjWaL5PTiAyfAa5oBaLBNpCX7jUsitEucW7L
5xnG4RQfm45bISGxaHB9ZsGCC5sD47Dz2VM3CISbfw1nF8BngOMJpNW21nFC
FF1PSA19qJbme+URvzjsernYqTxn5u7ZcaVfvF7KOU4eIzq0sOagpLJakflt
avNd6lTbIzj7cPZWe4dPQnFVTY9JvCzYqXB5mPowdEkYHQYFNVG2q/mrBReN
s9VWCqHfn+JONc6+zTOonYC4JIyeT83UIu23/Tz8Tepiu8NErLQROA/PLBLl
xO1/PrfZ5FEnN3v8UmNAUnJwQcfzdnOX11et05LyFYpCbUElXUadPMptaIns
3ZdbRuBA1soMecAmhBC8hQ/OEqjuyGG+geETU7XmPhuoPcMCzIh2L4VW4OG0
318MuutM8O+OOkVumdAU/43UCjRWugdvqaeo6swPFj8M4437juSGdeJ3nyB7
EWZ4BjsHgvA55BP0IOnwnD0V8TpfwlVzjQFFohpEOe9iZ1TmxiG0aLU3c03W
v3V3Uo94NZDM5+6biKSmdymmBIQli3b8oiU3DpynnRtU24VsadxUCWthsqw0
NfbuBlSnl0LcvjQT9M44cGom6YV/MtIQMn4Rjd8XSS9RCbjg2m1iAfHSV7II
K13qcmtEXftnKryPUbptGSW8Abis8Guf1mUaebGZ3rpCx0U66feayvie7I0w
4qpxlJkdAUznEJABoXZoVz5dC1zo5rFFzs5bFuQgrxypGCv52phHI3rI64eO
9aNKcpQ8NlNsCbbOmY/QpB7BvadDNjzYDSl/1PRhUDqzAKlovIQXV1fyzZwz
EWH3q/2vAoWGrp6K+LsABtzdGDM3Eu+HMJkH7apzNGgRf4NzmujOACjm6Kvs
yl3ioGaULCEarW0r/UdfjpyWER3X63QKsMdRuD3g4k7T8rDKO4sYnWNwucev
Nbh9+PWYSIq38PaZObFnB3s9MCNJdRbQEhBdCwTmAdkaoSZRekZFXFGqzweD
2vt+zTSodt0zZAb8/DubvdCF8WWpz/MkGcF0lZ5Mkq1FZI+aAe7uYBUG4chY
gSQIRB+ctj9W7zYnQTvmKcZsADRIjLKa35ci/gyA6R8wkCAJ2PyFvgH++mE6
oCktUKhCRVjW/JFCq1W7LmuJ9JSJG8bcxM/83iihXG11Rok7J5jQYbukmPtd
qmNR4JXCnowI1Q2XA5z+o3HF29Au7o9sNHej2OB8zXD+U0PEdC4qwPp4vdmj
IJeCvTUgwcoGHDPZZlaFOxdeoQ9YnG7Y+r0olmeWQW+d00XuU8AUgXtwYizl
OPItKGaIw988Whh1mk2PBdPFYzkV3yeODhA9flvAS/6ffztaA0nnO4HmGLVY
AO+43mLGdolFuyYS7GBrq06UB92Zo4OYzRs24Emh0dUU77KGFaLY6Y7u8ocP
hatfjlDo/sMt79xv4If3wVzWBSAQccsbDSpqxIwuRSGlQOhdsnfMn4P9MnWL
TJgh6XAlCbtXdV3hrFLADkCgE9pyH4Ki5lnGZFyOv3JMb7FYbB3I3hpAPaNF
pJ9Kx2pmv1vRusdcNhxOT3NJbgIVlwGr3V8Yvv0W+nGoqxD+2p6xi36NCuId
7mgoO4TMHq4PHY5a8kFhtjUfjYEpvBnULywv5cjWeU9bhYM5uiOt1xYlPC0a
YImih7bzjEXm8cXEZqVPLX+C12EOoq+pDbZKWwgeYYQSjG/pr5eNbZS/5A47
Nz/fW5hnRenTcJTx4rYyDcbsPpVZ4qpFRVPsaLd+qldqN4cLz+rIsoCBud9+
cpq7yyjbJEW7p21ZEFzcNmPIujNs8qL439KRhnrJHISNNhk1SC6uJNufKxt4
11PnfY8/gIro092j3U99DxWj6uD45BJokv37UsghhDj2wjKFrLmMa5Sl71lk
ODkYyd/Zp7PGGgaVizNX5tOa+TLfqz5yKNk28h2ckm/cmjuEeIak7xVQ1pst
+iMdyMnw77/+lmLCIbbtPTgjzulCfcKujI52HLjnJn2aE0eMyzfSqQJt+sKR
b6mAruRnehT6PpZl74mJqRvZrOTaprJvg7nwILRUfJk2CYTkd7cfi4YqLNYr
t3A8spHDCLVwqwwy+dJuXUonuJiDqJRbkyJcRlaOEsxNo6M2mg/+rQCLMKh7
KSyhYBRKExbQMTU8T44lBJISM9JVJBzP9BinOxOVmhW2M9faQ424xQXD42X/
w9AvZvEnsu0Z7ESjxuV5jo9uskD6IA6a91Z/LqDzNl7ajerPhMN4P58zFxpW
AXbDjtebkKMCVepBGEIWMEm1W+LnGRe0wxrXYZFZ2qxTgESJu7HukuOUiLhN
NkvK6mXQlaTG40fTXm5ftSfLt921M6vopRTFoV/6KPOYOd65qj/JVWgk/HK+
4wOmnlyQevrAclUHYo+UO5zV039yKxnUbfFK1tzjeQIl6bxSs+p8Eb2Ryfvv
79axoxtyujMbN8NTDIM/vIZtkhGecm5Et5mGexqVIzHl4OwU6y6MAesPM1yv
HUW0NYfjF3cioF/kQ7VjRDKkADIHA1GclTm6Q2etgxtvGQ1arWlXvTct0FMI
/N7OGtY7Oj+v3UfqX+peh55qISb4HYpiEI82xtfQ2+29UL9wHvryTQYHWkIZ
QFzYwAqQLgMKMdunAbnHTgAZHyi6IfXfQcv615eTQQ2Fig6mdmauagpvdjk/
oJ8BbM+gwtTabM+IEfIUKxbciYeZADzv1QKelGKxc1BKLokx8JpfDPZYzLuJ
iA8EbDecEcmAOLyy/zn7zABh+eV+4V21bV2jXWG3eKfayomsFMNsfXmJ2QEv
v5Xoav5EGLAGTTDOLSU1VdQztLoJhOLmE8t/WFOCaMvtWzYhGa87aN8v2k4v
y1kNZfJlOrgr8vDiqDFp8ptoqs7OtsomOpoJFxzJEp8eRlGtPIZl3goJ6RBz
pXEOCED5YRa3TofAt54SGpWfKupPaX45G1NzGIXqsiPLzmf6iMb+UQwNxIxv
hdkM5Uoro8D0L4trRTQQLvZ96C5upTBeil4eR0ScfhvFC/Y1AEuOLzqGygVE
+915CYvlQFB9DMqVyh3qb9WHjFKRSjjXkl+7UD9CHCYMpcSkmZX7cOfaovdw
Fmnp22YmDacPG05QbrIIJIa0JDViAtk4js+lzfykNKG0uq+e6w5UukOPEznn
l/bh7WrB7NTkllkoeWYBajk4BdeoubKuEWlvM89SzUUKNSli3mELWKr+6z4m
41RTx4ZU8ndWnwVZvy3+bQRMXlLR0QPRELCYY7zR++EpzEws+jg6juRiIazM
T1jHE5fdibAEKYZ+o9wsbxXzqhsh26upSS7H+4legq2512xgYlgdOhLo6E/c
ke2epFhRxQCKPVSsHj3lwDjmE9JVtizX1JEcNIhLSr+2SKTG4pn/z0dsPOWt
9VD6JtXBMB3Z2VokWmTqW9jXm1EnmIBW9LuKsuBq27sx1cxpyckaMF2Cs0qs
k3Do538G37eQN3kypzvhLCJy4WO1/oMhPsHskArA4+0G2BWtvT6Be93LDorY
ij/Nl2Q0QVb75KMzZZwN2pWksqMtFMZtK0+BTx0Uw9nEeyKnHFcpX0662zz/
m9Z1gTUETpdD3UGXY+uudQCljPpZpM7KFbX5i7aAwwfViYWgai3OlnX3vb1u
qiY1fidY32QtGYj8TBF7b/5fjpVBIMxZZbP7frHgCqGntx2cGocTpa7A7Lyg
rxRFopkyP10wXNxW0Ide1nQRlh4eqARcdsqkJ6VSW2iVkKE/kwE9W4JaCEDW
LEgmDK+6ISsogA8RwUkkeuHMhanp5wxaU7DUqOFebrkBGchhy0qd7kUdwH6f
gg+/86wQkmFLf0Lc3z1ytAU+1Ye4JEWX9lex9HBjLLrKbPKIdgdKrNb3U07d
7M0D6LiisGZDjoeS3xhA3X3bvwlAlkDLpd8c+4GzVHjlAbCNnts65R0sBHq9
a9JmzqC8EIocJR4a/utYdPBisQHR6EsMvDavJxzlDGguux6AoQS6KOQFMAZq
l07WKbVjaUVHMcJdl0MiHJF+/Rn5gPuYbqMwhG8yWm2THU6qYZc6D+giqkb2
LoPdY980QDXG+Jsj8Q+SmdNpUhFiA4c/qHo/Y7ZjfNusfc7v7zWDTW1ftSll
HgCtva+JgOly2bAGYAYIdLQ/K6yAnJW5T1aZ8KdQmP8eONdW16kInzVPOcGu
G8tMjACSpIdV3EMyDYXDIlglYrMDDjpmRtG5HRGbee26V3DhN+LtMbyCPbz2
2DnGeBzcT279QoIwbqPSG/NSszobG1ppQv230dYagmhH0leYyBCxbJHVIJ3g
W+DumQcS08PxnSzlx+QPzEs0jrHXtMwELApR16YaZBDj8zZZfQJNo3pC/ybu
vZ3QLooftMD8mpUqPlDvq1KiJ/E9/4m36XBGKbfdH9xiRzXDTQdsLCoTq/9c
U50iWzJt18WL2JYBVdHD4qZ4/M3jX1GAC0s+PM+A5Q1IKIYJzXarJSZSZCRG
AoUN8n3jO+arLOECcC1iwZtLxBiqgmbw8iXKJshTLoxz4ojWxkk3zFhQNKsr
CDEbYtLFjIwLKfKBqQ9nhLWXSwXZOOswN2uvCJEa7zREvBZjTlGmamyPwNtl
aBAZFeT4OE51dCCoYuv9b/RPrb6NJCARyf7kK8EVCIY4r63indF5R961x1Tk
NYst178dgDypoL2glhcfHVKuJfZrge7X2lhRoUcbpX69thutvwxxcGSYCBkD
DCiCfZb0EwgzFoygnEbztu/lYYFgpr7yiF4TByKowp617pXp/rE93RXzoqJv
ifmtRY+Z5syZLWJM+h/7nujqxlwzeC2SdAcRKgrAVs81zb3U07rE/IIEb41T
7f2z8Z/NyXvjf++RzzRLzFwnIbqvGc5rhinOrJ9QJGPRHmlPSvWlL9in3puy
jYj6IZfP++uXoAFqo3ia02Jem6uGn9V4ypihW1XjV0RiIJH8alxkye1k0gd3
YPDr239xop3VPpYrPdZzhlXF4cAGYGu3XN0yio2h3Y6CEOrfYaf6AYbD+Ait
J27yCEQobCOWdpgew2F7s6DJJJt4jEm8uAMTxs+LetrBM22oaT1uSW3P5cAY
wa5xlLJPOdXjoyrSrxiq4M1TViXrvEu1pOs/m3y9X/UlOxDWCIOT5m3nG525
kYzqooyyaoWcwD0Y/F2y6863VklJ3n6IBB9EdCbVuiCaXCjCsQsOjhLceQJu
E7iKJPwza51XJ2YE9rv+Cl/XYl2e5wIoUEVPiegbnBlTtIMn0VE1gSmWg0/4
bfpp+yu4qOctOLXDlmZOkx4QwZC3HT5tGeDOx2HxH114HpzeYgKZfEJ2L2Rh
qIk95sK5BKHCDWrtEXqVmsIJjZA0+F7MlaK9nmYusxLghHNSR5oxhEOnA5r0
cKCeGJ0KKgmIkU1BQVnFTZAVY1ofaXx1DxnY/ZYNxCZES6V4wf0rVMadvNb8
PfUlJ560q495BG77C/Q6f0MfkPOLuw5amI3DsIDa6+cDt5qDmx8QLFAQP5Po
Fz9YlnKvlVRpFqvdpmlMwFKLh1QMf1BdqerF/XFg3eKZFjwFNTTzg03YbUld
I9XqkCLQWqyPRRjAI8kck/n3EBWEUoD2mani9KlNxtRx7Qp9Pjy/zVIh+kin
t5aNGoYCFLU+bpSx6M0J+Qp2NIL9pfEVzHi1dKnCj0z/zifC20zjyncKUpKj
1ZCS9qgBAzlKoG4S103Zaput21l+lEllNGOoqGdU5YeBPVuKZNBkcnR7068M
wgpI752z/BW4yLt9jykNKlzEkedXuU3oCWaRCnAqLld8AAYsR/u4oOF6pYrU
WaNVdbyRCkygmtrcwcv5UftmQN7uUJ/NYvyaDY6g5uyXMxpXHGrXzKUhAtdK
VhbAMhYtphrb8lBNrw+vOI3RnnoInfIqh6q+FjcjK5k+Ivhd8zg8DSeI0p/V
qo8GAIChn+0w+eFeNgNFUffx5FbkVyQB21ynMRSMfVz9QthxzvOCUEnPQL60
MxKvGyvFTLICsJAk92tH9Ak04GEZOVuMz+Nk8pFOJO/wPQUe2wHXyehfaBOI
dZCrNR+5S1GU245obsPHJX01oaZISIJFWs+dieDdBfxXfHf/QR5Zlh7L38MN
km1IoOH/JSekseHFwr+T/uUNPz4+vDMBlXAR01zNh3fil/W8/8AYMP80WZj+
BJbuVKMCX8+ofvpOYO5YySxNasIkR7uo4U3v6kimZql5Qj19ala9kJyc/BLU
7+M/8lRpOkg8Qk0EdQAxCRxpxIN2tyheoIuRcLd6ZEGDLckBISDo4rDWyQ8e
qGf4Hh4wypmzB4uncxDaBQR2NmEHmgLewTnFNBNxzL6BW/Dwm/VwMv9uoMXs
S8Iu6LzfZvcVMvH9Z1dEEv4IbJliA0tpTi1K0Fd2uiNXIMPmmsZqsAtFbAEl
SELLKWfX7unbn/wRv48RSxgRm6cNIK9m1MwdpAsB/u6YOt0njiixlEjough7
VV2rhPqmEy5irUkAR3owvjD9CtxL1npnBU8P0/wNM81oYNogar9orcPK6lqk
YkLTKQ4ReXW0Es+ytL9VFIbulMO28gBetllLAAuYxQe/u26PaHQks5gx9/po
ifTHCpiSxr0L7eBKLcJBpkKR+vYGOtbpNZ3AfwJWOuT5192V7EAuH2UFqy8N
sImBNl8Bw/aweA1kh2u9Dgu5Otyu342kEmxbmYX0f/DgX+J4C/zZGzU9xEUQ
Afs9h3CQagF228oVtIe2FcW5JnTmV8cwUpwTt0imbi1qkOQfdpuXB/x1Lr5W
0OoUJlBl+qFeu3fgmTArB9yNkK+Bj0LdY7MD8KKXwtGRxomWTXzRhALhTzFB
lQLxHZQyc/SacttyeRn0Lm/bFCf+Wk9Dh0d8i5F7PNtoN4Hjp1kP2RkP++BS
FhQbkX34gIbcd1Q0E9TKpQFMWp+Cv2Z4E03u+cCT9MvyL0ap6D+53Sfwrov2
I19yRVXG06m8AA4guokGRVYoON8M4p3x8EXblq3MsUUjG9zfaBdPdYqBd5uf
poUa9GqQ6MRqx8bn4e80epdxsgOABnwT4J0UxyU1HNNRux6iD7krHN2ETeMx
JltuEJb3oTDdg+znICuWclUJaWUVKPzB5+tgmlS1xOZo1dDy3lo/DyxM4XS/
CT3yQgSpgyUyAzdtHXlUl/DuYWZt+jS4Ws9PRI2P0XTPtvlDrQDXTIzmxDgZ
plczq1M7F9vGyASYwQbko2V/VKLg8E0GxhajI7yzFZXLUC7uCHuHpJqyTSlH
PQuOHDDzViQuWXyfgOzenu+FnjRR3f6X4vBrqWS1jca0fltP0+KGdXxlFDEb
o2y3h7Xuw5QuEp+Bk4zPz6Shoxa0U2ZitreA/INyX9MBqbnH9IkMPLkUgLPG
xkgZTOYm3xdNbYlQRNSDIvasbiKL1E7QyBGDjDqo5EwvchbuEnejLLCJF7bD
AP3aI3PCrEf5K8uQXeYxyC8HU/2rTJQODMuwfBYkCDX/7ziFes2bgu1nP2a7
iQ2BjsXdbTL4tyhdhrWdMWw32aWhD2OEhCbqQzsNr8SrXhCL2vtrovT5LbJW
PpRkOjSGZ5TnUW++/udos+Wv/qCJSl9o0pqI0Nvl+iykSMaHsyk7ndgFlQcf
J1BdmWXeEU/l0RTv2jvpRCc1xeHhNS494uqvOQaFfXIyF2pBB4XsE6UzYvlj
oU+pmEf3Jxopx+/q9d+fS/1UfhG3z8zxNnwLJBV67XqTuLajmL9QoSeK0ArC
64a8i9q2W/ajdbGmjvFIONcEB3+KBoFEoTzHwWzyOpTRY4cQTGTlWcmi4Kxd
NsR7AvhSFNn9g9l/KpQ1IxyNxyGIgPWEGWplRAWSMfdqjz4gYFV91x5agzdq
lttvCDj7m9G6ncvXj7/w0rNFvuLka4z8hdGQ4URhKpP7mYW7lWimfXth1FeA
1tmNhosTlngU1tD3Wu6pzyL2YwZxtnIeJgePCiHn4j0GrTnMFh4kGli7VCJk
h1KKLq661fxytdr5ZPf4MCZmKH/zPuBc9qrdtqECgxgLuMNeUvkuHPPpnzWo
DmGOuRreGc+e/to7xMGjuLMTv0J+2ps1Xm90c7kl2VJVe7Re23N+gmKgM7Lm
6ohcW0UO3qB081e9GFyqB8eCjt55kTndtihJKF5CB3JEltvDp7wsKHS4PDFM
gc+37yu//Tdud8JpKjwkS+ZSFKXz3QKypZV6OtxiwASLUldWch6en7ltEKtW
nqoH4+F8j88kkjTSf6vTG/qHSSctLnbkWEo+pVNo8+81r8wYplMMBUpTRhJh
J6JmAvTrX92HeA4TtULCECntjdSPe1Ar6wYtXzEqpP0fKMSKWdH6av7xeY0y
LWSUcqqh6apUDe39Pi9nGauCu6u6ItoM0A3BGt7ENz3UhP1rYXRRip8MW+4N
KaBG4jS2IJhjElenaEiDCWRvoe2cFaS5w3Zd4bBc3K+v/npzJ0asuXlsempv
AtC4+6ErHic6OqCuiNKPZqAHiIOQT9yStTuNPmOwoVlUUP6+Xrr6iT2gREoZ
jm4+4IRnMfQJ9fbt9S1hlJbQGU3Li8eyEVqLZ0HsHSLvroaGDsH87XJjb6Dy
U5GjGVJWv34esW6MYDq1z/1iEGN3nJJzRvUEseKA96rf/GoRJTWwe3G7VDiD
Rg7I5enNp2drjdbsJklcK77tZ3UaxS/gnZ5A8TKAYVUW34KWOTozJ3mT/q+i
6+qatSWvNorjsEHEoxFX5TDFa1/KgsoVZYhpWgTr4CMHyrcGT1dxxNRiCbKD
BL214JPFrNbqfsy6Fn9l1fdGd7r0xbEJXSEt4s1hED0RSLvzf5DRovczjNRm
qtLS/2McnrZ/OxGPjf3ePYHCQOXcuJJWOj2T6D0BduCdUlhmRa1X6LH/oM1e
/iPIj3qyFUtZiZrXpxLI2Ed2sOjPLurlBjneS0PhmOqk+DAihOTQpVfaaXqO
Wj82wZ/u63UUc1FXOC/xHjRAwo+LUpctdkpcs/6XftDqDDFPA6fkbjbHmQWh
WzYbSBaFdRwX1vnOl3pf18v2gLtDLGizz2I3qyHG4AnfhPVF8UtfNffXa7Rq
dFtSfjttQqwuT2IWSGVQH9XHT91qKAG0NJ9FCB1RDytkBaEXEiQ73A8YEcBl
adwzVr7Mv7atim2Yx0YBLbjN25w9wibOcUKWyDwjss+z3bFDapjpk6Op3Q7I
/LQZuHliHlH9l9Go1DkgI/wlbBRHNhR7wDkWgG4rH0Yb9WEFfCzIhzuIsa3o
rUCOQj9Emb4hKbQ1B7JDFfn9PjVwpGA866/Gdat3mOfxJBrB5La7ayDmaa+B
YplwAJmh2Cl7DGDNPPrrW7VxxMpr0OVfldFy0RAAiP4JzRJCRHFU68/+/FET
Qt1Y894sDc9ZMx72dMR5k03k6d4LGNlyX3MYKHCuMiTn0VjQJqu7GZ7wOMEH
ZmRGgSO9GVE67AlwdJm7MTLommYvMU0rGDHSUjLLJ/ZiC/xBQLYToxaC9HVC
ryJLcG9icEz9aC9LWusoOIZU/WuwdEEJAtoJR79FKP0cRsJMhkJqrpOZ4qPb
bzm3gIKnYGIZORKYUvC/vSo1YZYKMny7saA27Qml35I1XYjifDYPT4LB+D59
u503ZexT67Lq2QGw8b33fleSUbsjFpHbVIqBIUu5UWkC1wXYDUDg32BOvBJ5
bxkq5FBwVWXKbOF+c29benh1hkU8yWuP0Fx9k7D1NmMYsq6ryczfpwYFFz/Z
gkbM6WOU/3IMyIPz18EwH5kj5eg8gGYOmqEy02r+YAxs+C7xn0EkzohOx+LJ
wYOJR/5VtzH4d+7zas6Pz496njtKYXC4RBuYcqMs8pmwOHrwBTBtSiXLXRji
GGJWNKsZ/6dkhdSBQUv96IBDzb3VY9S0rB+L/YL+EJhel2Ud6y19+bJw/ysQ
FecF04gz7ZgL0fy7l/0704Aqms8Av+1O/6MHHdcZZ64WVe4cdqc96hjop3tt
vlzfNYPe7aYOlrl67Z2hZigPfEEMkxVt1MQhsJ8gAOXjXIAatrZsA7BKKN1C
Tk78Wz3GwTadbyUh7OZNKM1qWo6gV6s2ucd+iYFO6QgXkYyxRdAc1RA160tB
QlhabKGVbtHsdRIoqiyBaD7EoM6QH2mEn6C2n1pTSfclK2ENguaJWicHDX5i
YYZuH679sDTz4cZ/7oI+6tkQyf5Uq2WUdE7ZMXmouCfixuCnpCuYY5SwOUcr
l8KEQ0lvXKJLY1Rh+pldKwqBkH7VDGHfi7cybEFczcvyZiSC7bmoNbk9RiIt
ubfWKEnpaR5WXgkaCb3Hmqv8cTtme08ick1xZX9k74dOkWhCkAWdX98WNStB
9ELfWGEZJ4/um1QdIbe1b6uk1GsPujGmd2qObsGessPm8D5v/UVpIQUX0JBS
Q5otSsxA2dVG/FjYKIdPfb9u6x/BQm2O7HsEJSOPVJbex4AZjRBz0pJ27p0p
k8XToUr5o0/Qt3TKehMK/6nvsLFgRvxXOHApYJSwP+t7UKHLL47sVBuBWjQA
j8PTNikCAt8shgeDRiy4b2DNs5inTux2WRk8MHhgiUV6cje4j1PZ0l8QWKaP
Xc76d9XLhao07mNlMclQ5irr/qXHriNeLYLLR0MeRthmf8SnqWj9ViuFYHMj
FNaHv9WAIK61y9cxlHGwBYCWdHqstoJEc0pG4UcovkUgcl0xxnWExUg4tIuT
YbrDdU40sUP91DKFoo48VeBjM+h2yIDFmxb1Yxr3EXUjPhwMGHlfBx3XVkAq
zvEIlgt9/UZohcWsZ8qmVtmUbpJD5DuWGchLxwE3NgdIosEKRfDfFILfQtF/
6Gc97Zp3RJ8KYqN502oyJuFSxiqAApkomcITX1YDjCEf/+MtsxLVAAj80k2t
g5d/y3VCyMKNPXW0Qz4AOD0xV8tY/XEBUr6dAutr6v8gJpy+2p/0CNVr8c8X
dgnCkm3tDX7e4kMv+uzJlrg3KkqqJ+THSaMrXrXVlVxF7EE47oigSuTCKZZ7
tWfciFT8MQzxy3R8u3KsGEfRyO7wcab/N5aJWLWtVVGyQWAhhTTe7jrno7vL
S6Yy2YrQUfx/9xQMa1aQ5mPHDVyYhEHs5ZjWTul1zaEiI6p4RqXlIxvnZ8di
25KhYhljxmt9oAGCZ6ZrlyzH6Axq/wH+BRWGhKrrl2KmGjCAqP+GIzBTGWr/
UG1rrq9ZTMPZGUKmPtbovFb4IJZhEREj/+cxFPHFUIzy34b67PbU3bBOL5m4
aHEUBoh9msoTi821YEOOswsNsB/uEG0Me9/yllw6ax2k+M+hT4e25RzZDSOC
zJnBdIVuDXgWNhiqJOSrjgde07vft6zRhKbtnaz6qKrjWrKeVAnhy1YfWa1T
EDw6GwbQ0MKMuACYeHsbBmvgRDEcjeTumpkM9Q9Hc6LXJ4zvlABqhLq8SQeZ
GioakuwKkYJWkxUf1qsN+qcQMCI6ORdqIHhv9JNGM91jl2pXMgeT1UUs1qB8
VrXpjOwOzYu2lCJTSroDNGNEPHuUSI9Zm9tovzmm2REvrR+uJiMUhONTdH2W
HRaNu55vSn9NXBf/sAPiLNDIufawdbf7iYLceyMXOiF8TP16DhTa1L7vCGhR
oTPqD593rG1qNGKkpyLMaxjwknOqFxKKdib9IUiJsEBPrD1dU0sGfEOYE9sG
cprD/Lz5mH5s9wrZkJ4P6yQaYyUjsF5VqTRVANJlAweVvbDsLmycCkbpq7p7
G3E1pDcyO/YLUz0xMEwO0nGBYgCnTQTdGKx2sQDJjIBaaYhZwevEyv0cTltn
ISopGSZImK46ZGyAz+iBVo54c1xG1cYwk3Pcx8ILbmRzURVtSgkKv3LP5FHU
haYC8aKpOG6i/jeAVzm0HZ7Nfsm+S2ZOSiKxUHOrQ/aYPEFHHadwkn0EwQ/N
Swo8sNDsOzdICkZ3fbgpMIpv07MyApPTOQq3g2NeDNidzx+TIu9QS8KrJig+
mpYVLzqEWF1qUxZsZlmVZuYUTOAwmNuTheiJMZFnygiFGi49oOZUfx5+fiLj
zZlMnG2ZKCOBH3+cRihcr79+KuvaZFaHXrCiBdNBdXldcMQBnKKmj1Y8NiLu
CLoA1bvI8bkfozJFjzjBcQiCkbOOdRtDiitTNJ2pEkI7SCxSWBaR9xRhLtmL
1kfp3bfY8m36m4I7VGZheelNB6TieTRBbhGR2s9WvxaHz76CtOhD4Wsk73iw
P735tFTlCEIjg/TDdb3LmAdbNnykhsb8CwPxDN3lnavxEVGjc1Nx3GluRUk/
IJNfdGyFU2vgiUuOacGeC/7mNbVfPNzUcB06dePWiOWmSVPHgDOOcJFmBYDx
ALYM7bzWcUHZVA9TZQzHXzzieYpWObBC2zrw0cFFk93RD71QqegeYeDJkBNj
vBhyytV5wFwt3I/FsTrkBaabYduuw0sJGrdoyxJxrbvOSd3eKYCx2UYFYSQD
Wa/CDrCDd2OV7qepDM6CCov7YBztYyjfW4BNBgkW8vZUalsHA9uV62BhUm7I
gjldmEaG8gSqErvjUxVTBvRV4dhZ+2nwjaJs7qra+DoazOremh/kd24hpyOa
ctVcQM537GlCY7A31V437jMYhNJ5D8O9V86KTA/e4ZyRQTxZ9f3CcYEhKLw7
tssELyi0jXJaQA23uuxEfzQshG2P+2xNnGwN4uZoLXxuzxMes9UOMeu9GPrf
3M2HTqD/IOIazwHIzEI5eeaaWZLQ/QU9MjOSqf0xCSCSUOLLDyzMhUf7oc0Y
oUu281g8Jir6u8xRlSVMQIop5zoKZA5N+OSw5+JK6JR8nvG0oRu2M1fnlMTK
xOXm9N7nwsLDZ/3d0OyctiZsZsAFOGHzE/QuAC3thtx/5slhhwPLZm3YvORa
o/doVH3qDkA01c8DiW1zOYm9lKzqK2ls/2xapbKB06UbZHIHVcRx9e2KGJgl
gcQKWSXdLSdCgGDr2UtRe7bR45azdOLCewb4ys/+waSzUYtrxsh8akKpeCXm
VFwcDSS+d5aOAswOemmXg5P+QEn3nvnr/MPLokCoFMSrKy9rsRK5j8/2kjv0
UHUl9CcvJ5QCod4hdBkAopDeowqazEJtusbXguJLqrlvNQrGz1Wk3ufWyr9V
cCS53Wpwi0iY0axwoeGoq7UTq5TllmBkpZ96aD6lB/Qq3zO/1TK15HQ9lrEI
kEzErqIrekyyJUE41bH3Hns8I/uij5jarskkMka/TF4TY/a0P4oZRIzDUCbf
j55E4MnatbIE+mKkWuJLus1dr1/oNlV8ncMqGip080VEy4IxDEAkb3yA/tM/
u9ie6J6jCu4BwYIJsk7KFPOMT1I8pnxOiCxHOPrW0z5Bvswlt3y/cFQdpIo4
ZllL4uipLUpacurqUtJwXm02DAQlUb7az6khPE+Ov+iavj4k+dbpzPH/Joe1
qy1D9N1bFnj63awPzrSZqyFkj0LYSdwrzZnWBjj6K3H2cd7GCfauN17al0U6
KtAZoghkwg7tRzGaqh0361TurQIocDgr3Tz/ATqe9fIOLcy/u1THx1/d65cw
BdY5EW3DoCnvpQLfZhosbV5xgXi+kUAtTSPif/bFYaCtIcRJGV09rh1TSUfO
UbXfHmHaz36CJufuzl5swq2RV6rVhFNmJTrxF9bW+dfN8nYprl6cZSqROVO6
/dFrbKCGUtmcuT13kCdirdDb2yp2C3p5nf5DweOX3Yo2kda+6wkXJv9R958Y
VH7Wcixch2TqwTg67snkuC3dJl2H76Lz5HucCDb6466W8uKLr8J0dH9F3bak
YcolsZjx+Dj5Np0BHGst2Ap/Kx7oYlq9mPZwBxJGVw6YmlxCPGoC6rXVEgPv
G0jQFDfT3szpBzcfbSZPRI/LEWNxPoY2TzysqUClgoC2QEEwV9TRacEPnI5g
IRvFNujki6VK/cAqn6WwsM0YfbqTvENOKY+PBvCVEV4hAAVpIP65YgFPHSFw
4TXKwbw4t2c+YPC65NQdgxdqdOGFWI30vJg1IBLLeJKtQu4I1zXiafuTCA0Y
OtSxKbCsxBPDC6G+JTkjcUmxXABvN0RgEOlQvMAqvF+ODKZzBxS0kAn00gNf
p3pYOzo0p6vbI1//YJnIhu+hz2fozQPlXVudvpxhrHuqsny58PJvWqZs3YAV
B7fmrv6OxIhwd2FPS2i1Kmfb9ttAhpPCvrErh2INSOWqkSu1QVUIKzb0KiqU
OncK9ETCK1uNMEbLdfBTTi0/WHJ1zU7paJ20tsm0AyDD/AfuMRA8IlqvayM1
O1xhs5BwkL9UPa8vfRxFFNpFXsfa1hKeedMEuGeHYouqw5Z4Fg3fEvSBzS0F
lS8GI5A70+t4fVxOSurQT+G/erWcEQdlmWW66LE+nbN1y5uLKIIWFZv62LxW
B9EOhwGTvgG/xlSn/E+dtyF2pGUm7PV7wJwJfk6T8JjOB0QrLUB30SNOt1PB
VYmEm9Dzl0m0wrSDTtyS91Krb2vQjkvyxmXZDgcHIlFCocxXvSXM6+eNb9D1
GmPMlVCP+La3GqRTYkUTrpr5CClVsPEgSQvbKCZ8DR+0VYj+Zxw/oGjvgtXD
0mEgQFI5rV4BRApmCwxCKLyGFzC9lRNbPB7Wq5goS986c0980+vPusEavxqj
Sf+5OOFi3QYnAL7UAa03bgoaJCJvildLyDSgv8hOZBo7WPI1eKI72+fDxAHJ
wgz/8mePkOpgqtv1ZyXmVBFzW65uy7cWN/BzBuD7q0XGvFgGxGMa7Z8z1OTX
VR1nFHGjbFxU9PwGbLzAR6MCpIDBpo34oXCUWgWmOpewCW2vMB0hyn0Q6KnN
4FOq9x4L7UvCEsasiYoEhe3WRpyl+xVezwWQXyfWFkaOwC97zsDfdhpO6Jy5
NkWIvNO0gywOTDZCa+2Q0EOGbPjCLkrk/Ivij09MfOoG/fBBn0u8zPMoY6TD
tFTTMcU0fUlQmBs5Leli+oEiGYJYqqbioldMFEkJq1cZQeA7LiMg3FWjhyUR
0+trQKWb2706jyU5qnhJXKt2FW+GTFm/kzu+XhzzPUhQ3SNmYtp8neIvLEpU
tkkBZPDK07PPp6Fvw3Dc7H3fmFpHB+i11RIOmH11u7Y8yFMbHHF924+8R2pt
04ykL0K+SvAcFg15Jd9qYkF2t2q6FkOU3sJ00dDcUlSh76Rr9cm9HsS3QntC
sng7zA4MiNHemjJQcm+KKVxPqfu28ZrBEOOP9V7DYByoqyLOBBUM5hpL3HDt
Fmk/n0Bcb9P3G0L4OH4WPR5wd0fJbLyA8ryg1wUjduu7YcIDxWIu+gRNfwnK
vKhIRaWB0SHP6sy7xu+i/Pap6Gb/1OyMV2tW5O+xLAiQsozKFmF9rsWMgq1E
43LsfQqqpayV4qTkKVkqge8yOgmx/nAS5w/PIjz9xff3y+EfWF9d8k4GCMWg
s1g8/4JQkKUPeXa1AEgDLK3mLn5s1dAxE0x4UcNCiECyNrlu709eaRR0O1R8
1xVulApVWuVchF5Nm2uvELZQzrcBC5yeZH4bPkxy/578X/Vcop0WH9y8JuH0
VFEjadHTNWvaknCPXMV5qzOM5cF5W1PI2a8cjQPHD4+XdeHumvvkhz8ddsRv
nMjgu3Jnh3vNCkVPfuSYqqCT1IP6tlNcMWOTY1i2O4zoJSRcUqOXtk+DOvO7
gWPZOqYCOkJ8825xhnU53jydaZZ19J9z6qlcasstgX7DDXAGqZVvQkNMPnGE
aJhEhqZSXnCC2OOQJUwE20FMxpf4kbv44vp4sifbLRuWsAkrb2UEJGexAa/9
tgNB+WY0E1+n0JRMc8o1qK6yUhCpyvj3BGaE9qtlEB0Wso0wZ0ATbPXnhP+k
DAfZe1WTXAKKcAwHWxB2i0WJ8OAp8BSrs7dmTLZoHBEmpdL1p+8mweC202wJ
MSoJwNPIVSxFoi5qOIg2AY/tCb0QJPXcCWkRRLZr2BuuGw/ZtKwA775RyNxW
4/mEC3qF7qA6SKTjQhDf+XILIBJIVKOgRJjAVrDVBh1XMUE1zJ5fYNiO0fm9
Hjtw67i4cnTViHJiMUYqOY5qVkd9l0WHkeHHwavuqCBSQz2cl1GRPVPK4gg7
H+Y+1p9sFL7mV61WvOEJseQvcLo8bEDWaVJGTAp9p7nF49ndUZGLo3ruyP0B
4kZFHsoWqpQz0thI5s2FKLixu6cbEAD/Cek1rqnNydxhzRArJnEoTWLisjZM
qB1YCti9ipIxfpJhx/mTZ/5AcXzD+ng6S4cemYUAxnDf1EYpWI0Qlcegq15g
e/O4tIfCqVGJlaa83JVyrTHDPfAprHKKqS/qDwolRbQdW5RorhtPL8+oU1zd
LEQHsiq5eyLuMgLpSbxwJ9YwRGBnM0TwIUZa0q4B248iJdiHZfCyCiDOqKdA
2t+hyExeU9hPo8Z4Hb1KD9FdIMR8nRvq8vui4qamdhELbsXT01QhujG8/uvM
4G4w7E0iuxTj6gvDyvFmk3NQbDnX9JLXeda2RzacE+lhllExQjH3V8KRd+GH
0m/adD9QXsDzGMU/UK6in8Hia8VSYi94yw6MhaTLVDgjOC1eBBENnj1s0gZ+
l6WrJhD5Tv+go5Ybg0u/UF2CFiOC29Uzjrn3YjKpURi7V9MVFk2bTZ6/iURD
Yls/Sqto7eGufOiC6KZNxAxdX8c19GBkwt6K9XzAsSzGq6fnx/Y+3vRAhIqY
WqO0lPPg8+0zFy/aaXOtdtsdcI1nLMqK3zk38uYnU0BmoWfesDl+7b6kQ8/X
78GPsmDhvk3gr+2lhCWKEJ0K/yfhQTvLZcRl9OdsOl0rVN+rKY3jHn0hsgWx
g+4U8wOLobbL2aOOcgbrmlvPulaj+pBaifXtUUDiAHewtzJqsQrcb9THRkac
nep3b7qGL6ynmwEKzzN9dXk+cUgm0Y2rnok2TcvB3GhkQw6pa7EVm5WoXUuY
FuAzB1XuoR9M5Cy6FoX8KUxZgXXCkKYe9/M6ugAU33oOgWLGYmcUkGlxXnCI
ggMBnN3uB8ngwJGn/OTg3hbqrMvIJU6iAthAP8PQA5fYpfL5H2z/NTTNTc2q
6Yzhfyp3qyNl4Ar/8KisXbrsPDoedl4QOyYc2dyPc5G5eRSv3DFK1u1r7oY+
gzsVtWYV0SfUAgZC3pmec+JPAzA9R7HwXt7EYsQDos0yK0x6xarGejCP6f8R
RwMVOFvsxoxokOWPmCfMyU59T2kjZTfyl4S1QQPkPafD8jHMObv7Z0uKwI/u
t+DNRYfx5jIxLYXJ0JPPsqDoqi6M+NWEdPJ3pxLmWGOB1Drf0bJbSzIwlAbN
QUHVMdTfPxfxONhEXLSDo2iXzI5CNozCS7849ZblX3FSn6UfTX9+vos6DnRO
RQbSGWZC8nBVmycacoEe9nNbLoJz6N5MtcviKhwRqq9LwzjedQ7xtkmOVf86
T3KcaWcvouRVBVy/QCeG57TqwwKFgEt7Z3Z6v/S+sAy8uTyaWfpigsnyw2t9
LwV2uuRPHre+eUl8CvYPalkwQBtjjGSREs9q5NqytFDFmjrpir4D0XK9mTpA
VGp04ZebZbdfcSd9D2Kf7wsOILzJdCXXmuqlxrPlO8aFvWGHPGorpQRn/IOX
9mBvKYpE35aASFgt4y5aSUc2g3jqlmGbLvr6s4WDncTXuL6M/OsjJILE7y8j
nqkMgH3bpKViBhGPtaRRu4BUuq0kV0SF4+bpVJck6VlhtVWS8205IHBo5QPl
Vow9VxxZR7CbF81izx6FT8CKWqzquhFTFCYrLpexLMLr93is84uQ1d2qxZVd
qwr6U5qtEmT6z47HS3rog8JfneOSV98aPYmWlSeYOF2zzoVv+3Z6ywhcvGjH
usdj1lozlvJ4esC5YcN8+MfB0smBEV5ZntJrU2Xnn7yET0RG3Nf2cdthkcBU
lK8Y4/gsQwNB9tqrnDS1Sv4NqXgyQcT1nApvzcE3I3amjoxRRe4yzRSkU3Vc
oF37IGfk0aZGziAblYksx8rQJUwTH0fYwfEostUjybh7AiCKVqyMHApjdKLd
4EzXh6fvWC2/Cf1F0tRtOb/py5U26X9pncVhH+RvUbd57OEPTfEk0EZZkcza
yResBkqCyuGUE/WRCLss/il3PSxmUgwiW9JqspGsA10CSc4e8x7x9JSPGyzO
nV4PCNmNJnq/JY9IXjexALHlQEP4lBQ+W8Th8837ymjOc4slUPE1SOERKmaf
qCAay8yawrdZsFt+5TfBXI8JKZlDFQfPkRHECQJ1tDr8353Hvq3GdlhperHJ
r1ujd4L4a4omXSzLffKSzqD19O+oMHC5mSJP+qxgfDyI3RTQqSjvQPk9vaVC
BLzL6b7zJLmIUZCWoZ0xVx5+3gPfrEmd+GQaR51Qwod+ix/reWxNwbSfs0R2
zZTGgAGXq+w83VtDGx9Bre4qdggNfiMYIh3OtXrqRvBEwfjLl1iAY5VcYwYw
nAdk4sTJokJl+OzBRa4Z7KkoyTgR6ty2sPvAQM5pEKVunVuMwl7dBrEIIH7N
AsiTioWMddzhj8sXDfJocXbtQbHS53NtenxY3Z/Xe+4v2CqT12sZuDFV+NUu
kN/XyqPqtiDA+3newd/16ZvUWiw/b7awsNd6m7BzFq5oxwayHQnBhNGTB5wa
2uiMPrAuN1vcVh1tWWxWuJ/fD1g/csemV9//cddp0Nl10y2jR7+zvyWWY9W8
hd4bBO8ZUxPqg4pC14wC9o2GblhVj1Qni9m8nE4lwi4Kecfc9F3Tt6Vq5GqA
oCXbu6Nb89jLjqbM278dIeI60fhiOBfM+Wy53NV0r2M31KWMp+E2zN1WUDg3
e8878lHJlLdIa9009Gv1I8soXgJhRdiCftbYYNptTqcN2NEXPs5oPV0bIv3z
eWr2UqIuPKN7CV/+46ypJVQDYvjDlBiZzByhqcWDPrwahvcNi8gLkTh9mcWl
XCY0T2RdlWCWz5jKowHUS82PdHpd6c050r1HQlzQT7GTnkPL0SkX5c3cpXOx
+ZJpAheAle1jcu+MJemBsB56nu2/9pv5UUjaTtPd6RnF283fv4AOPq0e2Di3
JMkrY9zWKee8g9etUmP8L4Ql2k29hyfMKiGHYBtVx3peY5yi5FflyG6LNd08
sYBsu9Wc6B/z3G38nx/EogdP3Hs03SVU8+Ui7sqGE4dRIocTALH1/vlA0297
z6Kp3FvYOBWruzD61q/YrqnE6ofejU5YvnPHkH6UW9AmsveC3OL25Wx8yt/I
+AzMkcKOT174Tz69fmqA8rCK0wC/5ipr/acgNy2dytMyJV8lLVSLfm5EEMTQ
ZzTgImf/Hu+zIA08YiVQT9RG7wXYJCTOZWhDOjO8DQZuGPxo/5YdXuLyhLvC
MbH9WCybEGHSda916V+t+2r4vJiAq/GUz2hkPXTk1XIqUXct+Zx/iIp+ofS3
+SwbAU0YPYhT3Oei49YFqddm9Q5MQ2KvYo5TPO0TZFNAMLYMXzeNKTtbwZEm
wdGyQJke5G3+vKCShXpqg28KmoZn+PJ/7oReF7IZqfj/DV1mmxkxT4BD1Gub
BpFL5VeuZkXg2Lqtu6ejrvUfWO/xhoVpH/KXYV77HZy6Pt+vG7h1EDEwXYKW
vRIqTOtbgf8zcaFSdMZahBOsJ5/YX3lDWsDbyvmiPokWf91PknU3bb69fdAn
aRrWR16mIjvN0ILqsGtgLBg7zZrcSg1MqXEXpYdGcgzLS4obtOdl9cvQQKW5
bRo+4fCr86mfTwYJrTofSUrRosILV2QgCX6RmJa19yL0bb4kqIg1vB+8tOb5
QUs3pnYMIai2DU0ctzkCuhGCXDk+mr1xBFUs7JMECXshGlOH58wttgPIxTed
cEq1K4KXZjYoK7ZSC3qepD4rz5tZ9ii9hLTepOB4FOEH7hPs4K1jpMafFdUx
BQ98L1NsVgc28ylc/3mhlNnDT5ir+f/zACE4tm0Byf2t+jUq7absK6pocBft
H+jGUbVbsiYXGx3YNfCcNCY+ySrpENq6Z1PkSdB9ec2iflKzE7l6akTlA43E
d/OwrMjD3VVILdTWq8CgEkiQURl0FTbPSSVa+FB/JHktCD4n0krcoVaoFijB
l2b/PuVRTQyWDtE5MTQbnRNKVaFYrsfeLYYWrajIxq8epYCP9haD3H3mJADN
tclegq/bGZJjX77NXVirfkQfEWS1EkNijYH8Ru+xeNPR9M/rtgZYnmiAM3Wh
HVnCC75vocL+FsVXcTa+UFHSUGveWjiO5yc6+AbSJaxspS75VIRDPFo9aYOf
PT5hxFsSXUWDrY0+f20yKtvzUwz1Iv9hOwCyRBMmEIHZvEG8HRssPz3tNdBV
rM+e5xiICAt9UWdx0bESiiQy1Xvx5dHeni80DRwLvdCE1baCisByLFoUrzVE
AD1njiq6H8jjsvNtgdWhd6v5SxVsIL2cBUrR7dhMDnwErdaVE+fTqe2hj/vM
AUiK+FI9ReZVpHJH0le/O/qZBg5GTT5m87112zeW32RVHVZ/xRqOdz3GvZp6
sD6ykswXdmRrr+P3OzErSchCIpW/pfHCMe7RmNFwciT0OUq4tO1tp2XbIpap
hTFjjyaYCq6vWB0CjDci7Bd1z/xLhW2+5q+Y9d18iRxHbtLAXC495AZYOXZG
4VTMSobE2QzAEgdB5aRdCWzwcyfaL7Y+I6nQIo+z7PB21S2N0YJdaJE6GDIX
amxgT0syeMJiAdbhfLRvkKbbVQewr7ddzQFusMJtXfHKhw3KWIjgQrPDTZZm
zCviWhz+dPV5MlN4c26JTynuYYErHTx35Ix2SHPRL9eg2vgCWeC4RCyWLWcJ
hDMB1yODChOzWNw6Vud8r4H/Z0LZbx8/f93ENDhUnABU1Sn+ctfet2GB5r97
LliJL4T3rprwSwAcbzwwrCbyTYiBkybHsjrE/th2y3uYFqvrxLeydST0//3a
nktE4IWf+qcLf1XzjLtrB8kGPpKjdaTTCsiOgGpjWA+lKykSah5gVtvVG4cU
iHPpb+FJUffOVLW27OVqPA+z+yxVqWKuG1HtMdq/98/Kcp43nUEjQIKb0p6W
7C1LIspW0KQ/UL7C5YgExyCeelH42ojJhpLlKz8trM4fTMDDFKxxyfS1mzAI
/0+eY17vbHjDv3JLYcfgymGnXCl+YMirf+zB6nJoqW9CIPvb+7GUahcgFWqf
QkK1in3LU6hPfG0SlKpwlWAsdam2i3EgphvYbEubQUT9DMJLaEuVqcBB6n10
xTTBtdJf3CezmkciJ+G1FAu+G78Vr2f3hjHLq7M5lTAzhoLk24Z2B0hFimuP
0CqqScs4NRUc5J4PCSWBKzF1M9mXTWtDkRfFTWyLTu1Pkcpv71+dnYwXQRgY
sNyyua3nd4bQ1ccDshGW/mej1yWa83bp6RVibvnYMvqS4UzuwQSqM2IAKo/d
c/vX2+eAPmf2YcFHkM1pBX6pj7ipxJiZHJDNXH7MEdYXU02tHmKl6rAHbcsz
VTqBUs4LxPPt6nhl5JsqXWAVsnYXFkBmCSlfWRh3fJLOwtTuyABztVDBectb
rMS5tP+10qmgYW6DjTY0f9Xj3SlHO1xeVkN5VeAeBK28zUJ9ZG2hV4TnwAqs
q//CC+bSOFit+QNOSqSpBAzWgTfGP8ALtJqeU/TPZo1VA3tM9bRtdQnLqsn6
sNIO98ecNW5Skn8Htun+/09pf84V/jE23/qjhbxo/kLibDOvXqcRRXA1R9nv
mbShov0fFkcTECkyGM/gBnYsgjT+CtPLjXGtPW5L6B4Bm9BpsgqS6/PmuR77
ivQNY5W7H7ac0LGUNar2nVUOkgfF24kgoCoajRjJDD3JtT0mFOahpli33fi6
Vc8jC2rpN66CV42STJkUJ1m5sRPY3AUZ7o45VaSmE+iTqKSO4hLCREDsiAzD
bqPCoIqvH0JJhbvaYQu4LVD58xOGt3uO+8NFB0zqt3RIf38zxljI0pGOjhkM
Li23IfnFO8zh+WVxbmuUJl/Q1A40N8gxfR5f+K4KrNEaeM88KdA0S2EQ/SWf
B6FzEvRm4BFcUkx0YcLZPWjTGbXSuTITfrY+CU4BcPdXKoaSbX1cEf7f/+Fd
Nei/wKBGbXcb72hEWPZ9a7YlRTWemLkD1PTEtdaljlAlgbP4gdDZWb4qNnYs
9maSCfb6y9cQJkSr3vlRMjxh+4m5U7Z0841gyPKpCJjzyzWxGQodbSUM2F7a
L+inoN2YYnZPlxaLaUX1LyIHmkf3MXHUQWWjB8rRb7PKU4DNu0kLrQixWZ78
4Cso3ave0m9wSPyoxlnn9YSecM9RcYWR6OUel8M6yTmjgFtQJ0oqScNbl593
y488Na6fbrNLDp6IB6t99HD8QU34YpxHmPP1tikIwxgCff9kRgkkyfsSqXAq
d4ACHijpD0ZKuSgaM2B+KnDe7fOV04H+EkBfVs55LZO39/T6DQ0iYth6sKWk
qVIrk9PxgxN2HtTbhvza241VEarWeo4ZOHR0TJNvA1yaSTrYbgpzfCKVzgRU
M8GtoXA26gFTq4SWnFimqb9FPC0LAXY4FeDLTXP/ros3TtZgUtR+6SxaSh99
rdc+v4Jy/dcV/giK04QUTK1JSuLUE0Zsbcg1QUc5ShnvsD+2bPqHY/Fm4DlU
C7eiEHLDfrsNoJgtOAp1Mqewxc6FVBnQx1WMOt3NxGfrOpRf5N15OrUEth0S
ZGb4CnWspH4KDro2q2cLskBlWI1r88D8Ij9voXE+G0QR2+u0Kl14l92Mgjlw
dwatQhUGT69LbIXw9rd6T9mGRqT2tZ9KuwXsvATNBF0lZX2WtAFjDlAQhiJX
d0BoQikA3oEmkbV6hxqCdvru0I5PREYQdLfFn7yi6ldszChbHI6W7NGQAeZ/
HdrVZ4LldLpkVa7VHwvTgyodzbTeDFr/HfqO4BMYrnHPVECbi1aQDacEwlhY
s2VvFwY+6TYUTIBJ0QQqbKaEnDAH53nn6YQwPBikeo8HfF57e2AAsUk8B7xw
//Mg8c2BAtHFrX5XY0s8XGt33SLSaZo5IqlgoTGUa2WaOzK2mLimmZQZNiVU
+iqUUBQcUZznA7+smFxnjjylgojrP+pw6ZfmJCyfWizGCTcZ3wUTDx5cEOHU
3LHbdlqIdPIMo2rh3l396m92hIvDKszeZPdedQKYyrxz1Z8hiK/Eqw2a4uFG
i8hksZnVOc3i5oax2nBiiNll7JOi2tB4/X4AuB7UbiG3HTiXmW8qpQIVjb/G
M4jAOtF/spGzsk991cOq8cV5YHrsABRmwPa/lA95fRKoXztNMgF6EVewmeow
W9Q8qLKvdQtitzde8tw6MzdZYzT7OQbYaaF2wNBrM1Hxqv6w4Q6U2lk/Zy7c
ydZ22asmasLXr+7s0H7XwBTeTeVlxQV+5VsjjR62qgDiz5HFNOW0DNlJEgv0
0haDpB5pOuOLlJ0SAYRCSne8HYOQi5HKCVl1LTi0PAEJu+7dLyfBbIYQWmJb
q8kmMtkPh6eacFiY2KuamKVNb7QdG/TzyybW0nGB+D1F2Hlaxfx7RPxSumnk
vuQ2PP5k/ybQHcbmQWmBU70pHy+gx7YeZ2GiWgf/SZWaBaQ6KZ8iucfrLXhk
ljtnJdR3LXRds3hT2n2eoEF+lhl6HnG0To7/xAPiYrgI0T5Y2fWpeQxroRk3
ZxJ2+KjYVB5wk1/EzSSuxs11TPXf5Jov2ltRATBZJciTZYESAo1rpMnyk87v
TI1Rvlf5OQgHq6pGGPfFUEun3cwqeQ5H3kIkQk1mBdrvCFTmh7NZFiVw2ppT
iX+revSKXQr1G3kIvdlbq4YGS/SHXPcaQFC8nreKAHJs2yTcRWrAgKziGIj+
2m3xu5ZDLLSy8Ny+N0XaF+0TDJMs8D9RshmodnbpTYaEJF7+5mCD73opRtQY
MXYD30frTX8q7Nasvzp2+RMXDeOpDP+4cXpr68rpgovpRgP52uAkGojt9+iC
0+djOmPjDuo/RdymmZ38GRWkQNuTmdD64VBH9XiF0NJSaj09iwEr+ZSfs847
XPm24ISfIvXoxe6J5pxvs/l/u9MboAtgcC89OOAUkSABoOea0vBPIGlsAkJ/
/wGokmHjon6J7g1mDFep3sL+1sJ78Jl7iDrk5fDW0Yf1toVLm0WarRxWNQ2z
y9JmPzyx/jhG3wDWwUkLXr+7KWVQeTcrIcL8x8XbMEyeeCat/TtSN3GlkVaw
99PLZwJb5zrxi0xihv9KxS50aTkp0rUzK7JBHAkp+c4MyQLhy97rj3lqNYOy
Yijic3D/HX23KenpmV0m8/+x8RzdoqUdgnhE2u+DkuiAQDIkiRAM2em7GECL
Tpr4wbyY7B90+lyceJwiTJRHxhA6O1R4B4QWNg/unwG7KyM3z3cLRGrvJQDI
8bH8eLmnSwwEpKObPOCJ8ga0jVnuy2WrupD9JZTr44UzWy1lu2BH43Al6UOJ
enFh/hW7AH0dSAIjJSJ+lqNgelv3ca5c6J5eUTYvMfqFmScurZ/tcHP1we6l
ZP2a6MIktboOrzbuTXiz7ecxZYNhX7LcsbcvlWGk50Ym9Y3PBHR87Z/hI1Vz
15Ma1EwkdnUHVyAp6OaV8xS/ejNeuWkoMSmefXfx2xA9UywJXwNRLKjTZQ2z
IqTGOzTkDMn9FPwBnD3BfQpPhAl6S7MLhohAA2/oVaY6oOMYcC3m40kwLmlY
cUcggkNBj3NBaLNrEMJtZHKHnHiywVUDZCPK5SuPVCPKgnKntxkOjzkXcfO0
ezCqoY/qA36aHbnzNckHuIPRvNkKQAxSPwQgktma69KQu68Q3OXOO9xSGgil
jr1mpWm9NMnv1WFwQlv7Zpr/hPqQyNlcXU81YIkiZ0rwXokw/7OqEvQ/ANRQ
ynFxTWaJJjeo/mvOG2mercwyZIOk9qXOYsnpEev80/iniiTROy+fLeO296pz
Xf6EueuatRcGz8mBV9oKDqaPYnPLlR7yp6l18kBobavhsfw4wzHW9U8VuAXs
ZNMXcZ9+uaOJjgbjpvlsLWAUYEgDd03GbLeOarCnrs0Qz8sB4Mi3xLwTy0MU
lXj93T1+gGRvht6snObwNcOxJhTyvGw9ZI0j3fR87VNo0e8wMEcDS4tQ4TwB
PxmPPT+RsJyy+wGZCD4LlZh6e6HdkNbawosTdeCKn/A0OWI6bZi3g3WlO0aM
korkIpMwTPTR4Qa7ODIzSENXmYRb6oXx7LsCu8K4BQl2uopH+iIzQLkKzbkB
OYIUfY+KdkYhW0BsO/ach3aHDAoYwfT1iKvYUugQjLo23zqUtu+Dp5B3Z3MN
gtEXayrUy6KjI+7PHbvLQgEvQl4Nk11lU5CITG8NO5AiXXs6m1xHg8naY8uQ
o0CoHYGLPFRp/atche5IZuIbHjBaiEj22ud5Jsv7k/vG3SHifrJlI8cbA8SR
9Pm4esJcUHOlzDArv0VstWWI95oxjB8KhFyA/2C555T4DUJdrVjGGtu2KJgq
gRHCZ9kMTTFWxzvXKYemE9SBa43NQXBb0WVdd38GhWnVQeoGYwOZpS/PqN6q
Iowiopd0jgrs1YnyDkNGtJcIlL3GNGfpESj6X1K7/IHqgygb7f3423ubtDOS
ziPvzSCVSTkOyCqd/y85gsisjgy64mVY2Mxf0t89x++GlTcsvnzvsfteOPK9
HSPeaLxWgtgBgy5O2vbsq495NnH7q35SpnvaECT2CAjV75kCcZZD03v5DLlh
r76EAlZDkUslKphsI9zi/z5Zx/7Xxd3F5xIxF4Ec0K7fdIhcjqIC4rFFSN/v
pCj7AH5e0PfXXbEO6AQtckf7s32tvladZSsNvHL1A4qbxLN6juzTHBaCWW7q
iJkGwnPDt/h5ehLrFZqefbLsVSsLPraZtfotZSlKlf1Sv4fMW2uoNL+t9wn0
sHCmH6VLgw1qPq/1hZjRIvvL8RJMtQk3lnQJmqjn7LzBps/r+v0teNcNTLlK
a+ZGfEGgtyYePzHl5Fh7pXPlYDKh03+BPr5BZ0GYjD5qftt8aNaKAD+zlX20
DoONJG6mdIirtGvkqHEGRi6+g8c9Iaj4ssYT5lO447n97Kba4m+7gXXp4bgc
kUpAWjE7HFR7KB1ZtyEaoGiVM+N4cXE2AalDH7xR9VWE9ADowPm3OFp2xJLN
uIgnmJbQ2jaRM31SjeY8sVZWURyjFlOUGOeaV8wgfbeKkcJNdd+CIZTVn+oC
V0WsETz6pKvXhyq1oeefqCdAoC8SF6uCMf8TwMMlsadYe2SZU3Q0UrX3IvQd
5ftnHkKggoEBpZESWrSSdAMKTGNXNcwcPkInrMsEJ7qV6V/Z/qadABqZJKRO
wPtcn+1Jlm0eccTzaKkV7g0rIoMTi5PUAIshyH9LnCQewNT8OrvCzYRRrbSo
NGwOEGTos2Kh5XxDs9DdpTypU9oSyZXOU4HqkHVdFYAf1fklYF7Krp53A+3P
E04RwrPlPaNVfUPRIK0xubnrvTVOiEIEXLaHwZRySEMPq2SYJ6F9rqfIvM0+
GBvjTsotJnczKhCd5F8Zi71sahdowEehSNfuc6uAuy5y8HTTwdE8nOxsBRWp
S406xtAVrsJM4mAaADHev3+HWNQgGuva2GHVNpS0DYCk46e76XCGgDTL8USw
BaMrB4SgNQHoZWoYRukfjJWzFH2SA5i9vVe7ckq2uL/tQmI2sLT5nQlXYscj
uj1Qlo0SjbkfIw5KDNwbviyhccTcLf61QAaMEtss/PdYb51uVwioFPCnDZRr
5UlNm4fd42soBviBa4D1QLAjBep04aFhzalyP5URNFXWtmKpBj9A3gEuBFTe
g8eX1ZQLoX6ybVL7oqXmPrTZ7jTLS0Bg3936ees17anbx1nzSHeFc9pQHNUR
5S/5h5mlsK8juQjn5K60t6Fb78VE3pJHRcyEqp1KwX8CndiiA89qcb1TG7pQ
Ktv1xGAcyU4UUNPc25STs9WLoKdXAfN08w1UB8s0qqd+cg3xpoNT58oB3g1V
00rB2CafRm6jRTWAWfn++CIRky12cNBn4oIwEe2b2IXegRssK4uK1/KoW29h
+ut7R1Mg7raNfclbCwx+dOeZi94jLmu1NpeIANaLMSX5gVa0IH0rEB4Ylzgx
GYabkWisYmHmN0+g9/MuYk58yOXAoVoXrd3qvnvAfZQBP9O8liUgZ85u1a1q
esPQaMaG4LNd91vwC/kWf6GJshpWI3gQ3eialuyDuBRpWJkGK77zgvtR+7u7
JN4zLzvZkX2W0EXqTT3CBJ602tSioQXwxdRB4IGm5Mm6EDZ4u99AfUdsokOG
ncYq/5M09I3RSNP++3ngzM35nYOsEmUQgSdy+eNSpEyvqOwrzNzjy0IlTah1
McW7nRL74GJnYzG+GTKD91OVmb+iIDOhLiGUT0zBKlm1sI1NZcb+kXbLV30S
q9t7FU4d/NNMMiW4BHFAoxb/JGKcYlaQkBTM09FbqHbQc+mWEfYeA6nFv0O4
G8eRIp3tuNYdi48oWLAavmZLMTOnC6rIBuC60ZhSi6Srr3udnFtlKFvc4O7T
zzVqECgebTdcdJ7q8to64CtSRwzpqfXjXlw3oOv6ctd5i56z2qRDF2zpnz0B
dbNllGh+5Ezonfvg0LNX7K9ChmvAS2irDvKDiNuiqD1QPZfUG+FzrJRZLpL2
8LpQhkXz0K9lbuwItC8eKO2/yeTTJgPcqGlH0vUic+IO9SNXSkH6PB6VjISn
fcVsh8rAyQlXdGu8oOW5Zxp32Q16e9WAxiP3sg4znEff75TDhnFEJMNm8fAq
2XDhsp1pm3glN1BV1go70FkVkqKBHgpJpHqz+qvJH5CO0MCWpG85im+ZPLgO
wrNRYgyzJbOfdHJ5584CrFay8VkXi68577yfmGw8U2+UgTH+z5dttaoxXhcq
0iz5uMpivuuQ6FzsZ3agd6h6avzNq/WaE3NXIkudmJW9m4Jz3bFl5g8hjmnx
ZwbkENuYgFH8tQ/3qlAXdDzZ1BJsr0PHwt+4f5XIg8F66uA8SXyj+ZfRWzfr
khajMvYEKhPVWJlH/0n7zNlrnXgr4TdtIh+U+OHRtB1bTs2u/MaCYgJ606U6
rBIJqoF7epc1ZUMN7XNO5nsRALYTCQYntCCSWRTGFLLd/glyrQfBa+zKT6YZ
ikhp9YRiGCVpOxQMhTqtgyzsAfCc1OywZxmo36CeAA/9DJOL0B8vxZM8+flA
A4x3Jmx3A0XBJ0/tffm3+ucFvvKR7agTTtw9niOjGWUlktz4VBTnqNm3GaHx
DMmVc6aEyxHyWd+azA1oZobqhbq+HA62OrehTYl20k0ysGxDzc+07YqzU73t
gi3cBUlyEX6PkEZ8o9SB+5A3+2469ftEHQuGiWusRX2vvpRfUohDojcYiM2e
zhzvtXUQ7v0OjPK9kRf9UBtx/g/nPuX1Pi7gw6a+bnL2NeYKF6tpz9BsBxYH
usj79ne0h7oKxJD4il6OmqZmMGAY0uG93wZ6777wI0kcmZ4a4qNxGkk9c+97
6byw2bbNNmyrakEmt4yDSoOgBYQDeGcc+giiThSqyQqPZS0CYiNR1U+Mn5rX
Ho9Z/4esdI5XbreLZrvrZv+TQabi09eyosTpO4z3F/ZUAVo5B6C3z1Yaj6IA
z6TkybG0919oc1cTz2xPYBEvSTE9hzAdPxtjIsUGST46tEsCpNKBBtFUWZuk
dePI24g51E1Hfv3Tia4qLY8GRWyWVnSrKz3nk1q5dlAoyQyLH6dT/h/7rchg
VEA7neOv4mHbATgMhduIeFsVWxPjdS9uiyJNCmOHDSdpxjLvCaNSQ2hcfeHg
e5Fn2ypxumC4pXXdsX/ja4+TTD5h9JcqqiUr0DHe6vCwEDWfFkkxebdgFljP
/YP1lVm1TBoDFY9J3zKF3tTTAkV73CoIwUI9VhIt3MtIa+qWus+7NFFtXGTj
9CxLjuX7K3EsN1aQMaWc+G3QbqbGI1BP5tLzkLI/RAzYm/jQllyJjIwXk5/F
1hYvxobP8vAuVLgmaLpc2dNg3AQ1rKXkqSk6PhACDweda09bzSq+nJcNndc1
hGQOwu/15U4RKqEJQJvnX2qEDOBOGPvRN5aUX/FgaSFkOmSy84lPd3C5bElM
87gyMDcqcwe4saBWnOduWPhI0edBZ7Gkozm+TBfn6kUnjI/7Xlv5Riy1khPU
kmzfXNtTS5vh0VEST6HHI+IHFRdWV8FQHhVxqDpAl0UoVeJ/7VwRh7gsrZm/
XxeHuTy+CgzZPl0OIR9sUZ7fFMDGbt8yiDJ1A/QAti21fpBoiy96KCYiNn3P
6l9SmvF7PuiC+ljhPi0gZGBB6wsd7iiL8WUjwTDBlNUx/1SrdKJXsiXfVCdv
FFPHmZfTWBs2olBumamdFSx+OModGovpz9IcbrwpzP8M5LxayriLTwVliffH
rPbBb/GOeP/GAR18fisaHUHpOop1CmO3ArXuIiiP8Js38Eka+DUCcGYBT8ns
JaqUACEpx3MeNUzlaolgezNX5e/ZqraWKkzB9TZi8h4RpubdTzxJX0a777Wf
7+8kELTtAMbTk18a2K8z3NIvsqg6JYp4ZBG/feyImnDHZ256WrDRjz4Yi+7v
B+OwhsYK0CawbK2tPzK1v0Cz6vzr4FwoWCPVEoZgxuGNiLBulXmsLKC+0VJ+
dKz49q5WXC0PHODNm735IdS3yxXavLDOUmCGdxC7C6DaGGGMh6ac/p4AWZMG
T+vbgN4QT3p7/Hn07t8iOgsWuMkTrXOj4RzrzXWFeWjIj3+IgpaLGQra7lU4
lM7mEwzqSzFBLUVC7JXL2TfpJmmgYjTmxxdYKA0Gh8S85MUXAjaYcB0eDn5W
Ew/uubEhT7LGE4/Ol+169fX7Xa8B6517dc2SEh4jobTsD0UjH3PMEnrjspi/
0gzLymIkpW2Z48Y5MdUxRiaFkuzZWzwyM/bNBt94VzUAw9v+2dHx1B+F/lTx
FOPUs33e7Ty8hH45xrJpZM/rRBOpUU6caVyk6p/rhBd3ITKIqpk3kL98OZ9F
s7f0dQSBDowaZRySlYMlx85Hde3ZtZpDykps4tvevZIPWCPukba73KYLhfKR
Y84bA6AkMxvFdiVXwhzUzmcvUh6Zqvb3nGrtSbwOq6KGAozuv7nuHlS+iU2a
XNdewtZPLMuCuNeBajaocQgz346Za5gJhN36A4Zt3ktpIFQxqrZKHlwnq/qC
DiMptio0Y3hfPOZO+kRwTnggk6bQC8VznLAPUfSV7Ak08wH/bz0RhlsHXt8K
Hh58bNb/h01Prdg9fadPhXJLsFJ9a4K4RKTufOklr5cnEamLvaj79YD0um+k
DNWpCRc6gqq9ZBZb/19s9uvMcOwmJofCwuw2R7IQR3eIT/XWGbF9bCh1u86g
VY9MedNsrmXBx0cDrr6pVspJOehrtRAO2m+uVZud5lN9CQOkMvcmt4m1bZor
rneuPjamn2RNItNLxgrbD+aC2MMV6hH6TOcyF2Ajr6EV0PwfnaksNIhE/Rsl
N4DxitZmpstmz45Yb9UrXNCYYjBZfKYoVsb5jxx8gz+EsBiO143yWbRy2u98
PjdPKhntqVPapE0RANjKCT0arGHEWzwmuAoqq0rkOOJfMSmlw4OXVdQc7+c6
USidoWyzag+MH1X5XmKIE8w+UW56eQtOcDOvKrvw+a2jtDwFPQT3cyUU2OTn
9n90chIoT53I271+D7UCi5TVvq+/heyDySLykwR0wF1MY+IyInObAsdxscRj
/5iA397KHJ9wBBez8/lDDdWcitRDF+zuAMARVS18rcV3hbGvs6HFrMk60Us0
GbAcA3UGLHK6QxpsCvAKFWgFHaidXjv4FYWXCISzEs6Z/0Ry370l6LenbwMw
44Tr9nKWld1I77JyEOD8KeL0MsDninte1WOMG1N5SE18AX36co+6cHsCVBOf
DUJgguU/j+3Pnac1+hIbIB2jrjyU34p5Cth9zjjnukEdQm6QG94PIA3HfdzK
IH1vIZ31H9cwccc2O/FYwOXLfQlyiMoGxf7eEuAU+KT1JfwYGyvywfE0fYsQ
bH6kXrwV56wsLAYjc3GwHtmBVPYvNVzCpoJ4C8/WFYxYMVu4l/I/CzHLiOaB
S/GJa3luwBR7lzS9ZN8o48n62TBURQ0BF8MIjPH2jAGqczD3p2DBQLgR6MuA
5HWRvIME+n7z04vKzSXW2kpkvTAv7skODBkzq5L1e2TR1E+ec4EifSLC6s7k
cnLqPMAiRfqE81UBSYfAnsajt/At7RwJoSl+os51nQ1DTRRiAVXR/1VIzDtm
z8mzSHSxh7U/AzmngJVuE0b/KAUj6mSIRpbzpBgFtN4YoTyDMGIpXZZNJOJi
WlCH1Y1cY4NdXO2K7XOdhyobfcpoE01HUtjAnv6l3vPKPuQGyMoIXP3Gan4E
QXVsjAOSFvGmZm9EWKpL344cnyALLyaS7HUUpk+bDEM1IqeDxn6tvPhsYkEb
4VaojosBcHlKmU2Bh/iQMvnrmteCTcXwHYhcyvZHv2t7jQ76+ZDgnf7oZTyw
5ji7QAyBUZZMUhAxKmNZdf0V1w7vQEdXW1WlSbYtZNMDwWTCATWURYrbiG4J
3ahlNgWxiCR4HhP6YqfftdSsTocCzLwyWlRkj3agxaTLPN4uN3n7z8IBWDph
0n1XIs/bNgNYWoUoZarnBIErQ42vnFp6x1CsW9Jv0OxpjDaSFHnYolgydAKe
tYruelPV550k5bZChWVTYzw+VPqeTJB6ZNATlOGXTF/Davz1rTX7to5AkWns
eVZ/jup4M2q8Y5q6HSply1hIAIJZ2Nl0eeY8cf8GqHI+aIHMsVkywx226uan
YIEjoD0zODVF4ZeAzRopc6H3uDnNDbhjZ+Gt+pyGgjuLvwdTvcpM00d04LqO
r4t5VOUkVKdt0a5oGYC6dR83oyWi4MH7QkHo+umoINveTZ5XoDg5Q/YJxN5R
zbU+pdnoB4/FEi03Qgm4F017VOoYjpIN7oZHkV88hdIckQIHjlz4Xsf8ozE3
3zmciXLjgelmFCPeILEqkmJnPTz4Wk2CsVJP4KBZ4ZPXh+48KYxxAmiwUszi
mqZZBqsOwtPG0snWfhDXBqy5ZmDCa29E3DNAQGP0F31QDY6Em9euZo6+ytx7
bFP8sVRdwodSms21PUiOIi0jkg3xKj27IyummB4jfox7Q5VPsjdWicOTXJ/X
fXbcRQm4GURMeQG97UlZVX+OjMf47KFpfkQ/iEWV7CT7JEic9OX+G2ofSoY9
nN16H/UH4NUxMpHCcbTEzSXYHT7EW/0Batxs/uVele8Q9yWE9LVW9c0UJqfh
ytbvocKLJ7J9LQCyTD4O6yuOCFIv+shJamDF6A1XZ/WCtqzU5TIh9Miu1tG0
3xxPnOTzSu8sw4pRNQ9YtQWHK7UrvdTJ53goWeWnbHdVyrB8DdDbA9/hRYVL
FUp+seYAPN6qwUwPqV3LXRpWgaOId4myMrPhoPIDp19jHuT5k3mNQlPTyw9j
acrbkuMSFI1YwIOxpLn3DRLg60x3qcWFX7IrxwS6kDnXwxl8UGyYdMjpgS7i
7B4gUJSemQu9RILIVOOTC1XLsdONCiNg995UQxrFOuiWe3XSw9bK60tmm9ZT
Qipvce0KBZJuVNI9hNJjGmsO1poFYp2dMT7FsN8Alh1F321Bcps2U3Eic8pg
agXQq3kUVHVJDGpmaYcWSU4s7Gn0dWF4/DYC2KIF/sKCr5KlbYoA9nCK4RHD
GD6vvzmfxjiIpv6C2ekWXgHOnIcDFYoxwTcqauQp4slOt2rjVk165nHY9XYH
4cW3Y4QqK6784deWcRvrk8/qx/Y2fV5gpTUv2ObW00cenaZ+oEt1KGlCs7vE
B0AH2FrwHYkcuLT/ZYP+janrpNyJQdejCfYIMAIVa4YOfNR1CPw/rdnXSd19
Hvkkt2JQ2BXVertam2jjL5LWnm2sIdIS/thdWQiewk+rSEflYcXPyPYVMiKr
ApGN5PTISTHOtzQD2LAiaBaiBMY+EM0lfbrCJ66aQWwXQ5L2OS9cdILqS75D
NFWTeVyDHrNkJ2TNrG+JALyBgjObrRg8QMkNvpNNNj8uSledptxMtUIl+qyG
8iwNHhwjkVwoh9Tkv2nO6risC11FAJoxwj5gTxJoN+KdYwIHn4pbpjukLQJm
jKEFeyaUwr+m3cs+PqHFz/rX82lSukszUCoqAwXXd+uJmK+i58xAK95zTYLK
xn/h4vi2/ZxdGmOqdpbzRsrHMA0z8+Px9at5xTITg0skVClq8lyS42MW48mM
i4tLtc4q6uS7Zt1JiyLbgx8LWIK0aP6c+c1msP1swXCn8QJGkaU0PhURfuTX
9iBkPQFddad3vYb1TEX7bpnReQus5DQKQDxOEH/saqqf/v+3OZ28/5gWwDW5
Vv+8MFmOqw9bIsoVg1KXqJydDETgpktWnmyqopLd5TLebOcElYg9v0eYn0ty
KypvJqn/5bzk8q/9Rr/2QxUXTIIEXu+SjXBY8a6fyz7noJRyVcNwRgM5kDn9
4VX2hc9cDxK9gP+uYyPqdbr2nB2VuDm0N8vY3uMSH8h8pLJsIjt023QUs5IX
Oy07WJdYCtCfZd/zjTO1QcsgLLgC+83rSYNM21ltIJN/xLYrCx8gbfZTrKIS
rLyakGGD5Z6xErjN3ZXnxproZ2kr5/B/6S3Z7/fwU4cjPquOaFivF1HGmdtA
ha7eC12M7OePwZ1MuN/l3FDrfdimsjFyFz22pA6d0TJrmlo4CzRX6Wo9Hxmy
Axn6Yy0fXrVJlThrCwG+z2nQQW08mP8Vdx6EtuKPw2IobLkOdFvKVpLfBaTr
C2dPQoJ0mEIZmzI2PyjaGH6mVI/5R9mRQD4l9wExhChS8Ew5MQ0iXGRy9zEq
pSUeV/+XONrsrkE9tOktO+hlrmO5p3En/03TK4hGKLcvBIk0SqGCUhwXuzyp
yN42PuewIZqQxjyz3QNn5eHFGo5kY0mcnBRo/Eq0CiGgGLCQ0I9JxgNTgzNK
Y1XwU7KMVTyRf8zmsrmt25W1ieQnj6fQP2rC74mVAT6Uti/DDbPEX4Ze0YWT
1/Lw2i9oRW8FNonoIFrwTZAGbxFR74+lXpIOrGC0AXL8r1uYdSnY1ntKjWu7
J4PrCVUVl8AxIe4uAGKaVeKpv5tzf8R+JcJbsTN78VYBKP7J4kk6Q/cE0M+t
bGDVuPjjjvH0sKna0GnCFSeb3JQ6NfyAQaherSM/mZHW2H9w7X6E7K9yvpfG
IxVTBcaZm8xke/MToC/mDuJeL85kVdC6PzZPV4tc9rCENI0DKps2lHDDHvx4
bj7hwt/eO0Ljs4MYZ/E9U21wpjzRwoqjE7cNIiH+t/kPK+hsCXzs0jtNnvvo
u+1yqJFtYIT66Y/jxcImMLmN1es1pnhxO0T/gb7Myr+xTE77qL/qqPPts2d9
PIOPhzaY12wjIXA2ify5R4MDsIAjtOXNFvVdpxmd7EdzgNVjFhC/PtmhUbWZ
qXJbKLWVyoZZgOln8jNVZM6qRbHjhrkgJ7QU8M11fSR+lRvp4t9OaNnvx+68
88EOtk/hNAJuEUmmAP77TB8R4zlfD31D+klOWab/RkMDF4PpHWMt2NiK20I4
qNrw0NWZfgusJQnisrFQ/lAtYGiJz/p4K7R1kACKcNaJNgrx6EpVTzsk22vR
AQmevMprECsYYNm77CCtRlgpFuzSndn9Bj/8QcFnUM7N7e9LV8M1L5L22BRK
MkSYtvxmlR6/20mlCsc+5ZrDvsDNHSPEYuoMzsyiR557jDQJ6pasKnUr8lbt
q5B8/kzxi/pQqQNgc8d4Aucddo17Ax0+ksSc2f0FA92eMD/rRSe0dIrZmctZ
g5Aym3u/FPrFiR6AzjbGon05gme2kPsPPTpiBF9d0mv6yjIOqSt5ugdiae0w
dq87qOT6KNWQE5J5LqkmdyBN9DJ9BRC8wxc9jnh8WVA4nUfDFCmuiZWvXXjk
YExpVvQyP65dV9YmSWAHi3P/rwx5QjQROZoAJVLAkYfHFNVXldbUus3NG0an
mD2bfm8CYWexYlWfO8M+jbnaMLAcY/gVB7hEBaJCcXyKJ7Ei+PHTn8mx0+Mw
k4f3A9Oq1Le3T33jE2rGoTjpPgbD3joYs5W8l731rzmDoKWT3hxmK7/Ysczo
+ND/1pFDKmxJkiGxBaGESsRXw3W9lxQzXg0VOQArwMORaHcSWM0EjprLb7qZ
zPITMF/KkFCUWk9QPiMsJ6RTmzJaoiy+V1w7BLMLWR0xROBMULQ6s7M2sktT
ulg6dCDTbpbtAjVFoU1o2skwEoDQKs8GIhj7Q7CNXNAU/5ICGSerJTkbxU7+
YvFyfAg7EWK1oPMJECxYt19n/gndTO3AYmOzo2XqvbXwIipPDtDl+hs8SbYj
WHAfJtw/tih8XtHcjCGC0eLM2jvxPxZIQxHfP6IemjXqTrcvGduKzBajzqxH
RF2B/b0r+mKeb04Xc5QPXJ3h61BG0qvNaPZCiHCuQY0KaznC52LSKAjddqM5
1wyBlwnLEoxxlKnIv0RcFsxlM0oJTBnZ8ywDVwjgReEBBhzZaAOVscS5oJuz
8TDE+4pL5rqURNNO3G1ue75tVEpNi8ma7almtSROzte94DIqi5tQfMvEEFTu
ZIE/SteQF72AQq6Nvc7kQKbHXwoJKgkg1vMP7zHxyc44TecG/z5CKL1mFWPr
+cBcvz7gtwpVni/nDTOEJWz+I73ounVkDvl1Mmmif2h4/KCRRqhK/CrjSd2Z
AVUvwl2fSL1QDISbhadLP6PJZnKYC+IlSN7AUeIPwbCsFAZ/zC5VRVpzUjlz
Daa0PCfwdjxTu3pXu06tGjgkDzykf+3gryDy+i6eGt3AMB/ssHMchH7AIYJr
clc0oItlHr4+bLavCy9GAshz1WkkPNJwOo3beAXzRjDuseOHn5Ix4B1W+bin
cVYMfbFKovxYuzff+hkug0DcbKrYqosLm9vtSe2gUtC+4CghEsGc2K7LK6HT
OJQ6oHOV/3IyIXm8Lexnma3CJuiq9mj9xAby7xkJhpQeDzZ+ULvaLqeOykg0
uwUldtldaYWb5bKyAHW6qL78IlSty3p5iAdFuYWc9f2bpeya/7M7B3kDV3dG
R2d0cFVy9nUXyF0z6A8DmNZJ+o/egXxA6w6swusuV80NXy8WQ1OL0/K+0RKe
V0TdYT/FuLu7sBGhAfVW7zQi+G7sz/VA0MCMGPopoy05oJrq+aU04vi/i5Yb
Sav721cbVlmo0dzfBgxzcQdtDzxzu7od38hw2jLYXJMMWY0NCOrqf8uH3q3q
8Sd4TF0YZTA8cHCf8Q3vKJRgVZ6oIwxS2sLJxffF7VKKPgh87kSd5JumsW9I
/oUjYRJ9zbfo6mABEYiDsyFLLSMQiPn366qPTwuxOkiBYk3YhwltGe/x5KTM
rNPI67eoIjvNnxQk5z1whzE85einxGy9KlRpSnenX2Yl6yl4sbeOk/nKPpdj
vpUfA1PPMMObeIzu8ecCxXTzty/nwrJzarqLTIiFZts2yG8//B51YucPzzR0
iqzKVf40vi1Hf8florksXow2+tvO6llWM88uY7ftaue61zxmQj1nup+VwKNG
3z7ekvnuGb+JFb1aNe+gmhcsAzORXTYV+UonYrr8juEF52tm2WaKEWXL1+s0
WhkXPZ9mOE3bnmMbxHoFbD2nEEYkUqHZk1yRCWScJzVFSAV5NPloJjkhmgde
d5iOFfzksjk/7vEe7M1SQOZLTTqrwkEWVy9IWKsPyZBnjYWUIkXu1zc4fh9L
RqR8znh0YAwtI8lz8lAumcw10GQHjoUawNQ451segXrWAgCjTIffnK4hZ3wr
gI5Tqu9MAFvU2nm8DHKkJZQsPTIQ8gFnJpIsps0Xsesn2RLTNsO1t8NOyc2V
O1llaHwtZ1DS9mOYt+bWmDJ1E0eWRU0G5+bxlOvEE7Hej3OVAM2ueJ4HLpiq
1lMkfIGY0wtwV/Kc0YbSVlKUS+OHnlmHgGGLeeksEfmDMZc5ZbZi7uBOf3yS
IQ4CUGtJSFPYRauTvm9jaFsx45gWJD5JLOFCp2t2WyGqN8jzm8/SRTaBgqxs
VLdYN5YvH6BYwBF3XLQWucPy81Dzr16bGG69DIr230Frj4Qi+coFRIrUMDtn
4qP5EwrfmgB/2OM+PouCidJtIDPe+8nFHohXfeC8jkXxtwRnQ06iNJrfwtsJ
Ic2KoMj2UUGqcGWvZ5L+mVWhyb2ABdlt5BDjPfrMw/9x0OcTolOQUu6U+nW+
8dYsNlAic9hiucvUl9336YYdexOwGGnJVmvbjhSQuzAm2Nz3eYdmsoCL2KQ4
K+xvX0Eo7nU7/L1akr/q6HBkKP6Z1bRicCIOCQGXwEn3ScIgGCBcm2sluwHp
sBZxe/S3dva47oCqgfswe9/WllZWCzwdHl7xwueMg7tom/tBhkX4zqJnw+4e
WQ2vvgXpcZypX/YuaKThVcvH0tbls+xNEhqFQIFYWhOS9KUhQiNyR37aGOcF
0v8c9h7r/1lTY+1XVpxlCO3OI+GzXex6D8u0d8ELPCDm7rzVpk0+5WbbWgQL
IVafFoHjlgwUzP4dAm/QC7RAxzE3X+Elrmpz0qxvLehXl8NYItBXp1gHaH0Q
jhBwfQ2WSH5vn8SWqOSC8syr+y7GK0ovWjsOksDrk7uoOSI4PI4kATHPvv6Q
IHsaDO7pbPkkf5INcRKcZsxYFwBx4dF8mjwAvZ7bLA28XUXP27SQLM3lt3jL
JNLMxWca5DEj/Wv2eBLjwFSZCefmUp7/dGGAJsCBeDPmqYfWwUqteindAYJk
4zYxW90SZB4quHuuvvazj4cz8vk6fusYSuaUdMOgyTPC8+sRnZY6PR7zZxp/
wEo882uYHl4WL2ubNxQMwmKlcX8FHKY2VqAwXJH96ibPaZZhXvDpTCT9vxMN
FdzDClH8UxX5iiXHNvOEPAC/y6zK4d/1eqNRfLTnhXIalS4gRKpzqIcZHlir
Pd+XlyL3ZhRgypXgWEzHW04bnAN0bh/j9lns0b8vgpnOrSMuerPMNULF2voH
JxAZrIa9Jd8V9djhQ8pzTA1/wm1x3yES/+PzdXqz6Q2OBjiaZC7gpbQ0f8AW
t+IJL9fzM5P/0PmENTu/sC8XxCrl1xw/jVbuvAnd2dz+JVjFRbl44ctSPX9k
dF1B3CPKpsHot72bPURDyikcOY8wRZmr71CmZylfXMIyZwGLtMioj4KxMpWN
bhvYKOrUA0cteZWA69Zl0Pac8GWBC1cQoUuOR5xctsTnOT7kZsbwVJLVul83
TCMsFObkQH+R9suMrCWdKOso/yRChdVsZMGUrJxnoVMz/tvWVomFOjLhdWTC
GcaGHZtXSH293/uxgd7MyhCu2dyrBl6xv01PiUduYoDzF4thjsgD9bCkWPde
wzi1OjYlfG4BE+geTLYhF8fyDrP3/aEYCT4LS+FPgxIlqMa7TUPEyzm5toTi
qiNfM8JDwV22zOQ1guhw9l8k5rMEsrBAyBki/LKhOZkK5mClhTJI2lSeP6yw
vJNx5MRyCWTvQWuK4FLElRSu2Wj6vCWn+kphET4qTdA6tLKNMvSMJ3ISinOx
jbvLO5qiGRIlqp01vngVRxcAJD6qP7GxNWb5/ubViJuiCUZFvo9tU6/Zhlhn
wq4nKUt3AWNsofyqg5hAS+O2bSn3EGf7a9IQK8VOZKt0mL8Bsomld1UrOBsc
+tRiAMpbCaRTXbF7QhwJlwW6K43Fhp5uN8HCD22SVLWwgyJGVRD+duc0fnM6
5R75IgaQv3+CByc4zpMUMuiEW1o2gkgjH+eKj+XQ8YbOVvfV/nRUfNQaaiH9
xemFlV7h/Tyn7thh1/wqVc5WVNsRSnv7BEUZkFZzQb1YA5+v8KlWUGTvu0YC
Z3BDNpxfeiSOY0cfdH37ay2VqjiR90E8tGVZEq3MACd//cxgudbValYl26NO
3O8rVjvlqIW4ie/N6bEbRLYW5Mbn4yenkoQJlDsZuZEQdnMDMvrzhQ/BwoZK
okupyXLznuxkr0vjcu7AuYuxOkfa+RCFoUBL1UhXPtYK8Ik0dFglMtCLAvqG
37hmO8D2VclC6kWahXg8Pbao1B0gMDX6+fhUBguqu6/zvv+Ovv14WbgJZlOk
Uo4f1qfcUZoiTJfkb4MeXj/6WcZRHxXrLkMptrFmUBb6VqyBcN9OuBVkQC+w
Ahi76q8Q/ZTiW2LHIqea7x1Q7Z3agzo38hUE0xS6Ynpb7E7/vQmHoKmZRHwW
tYDiANj8MHda53xrOZ4YN8jDymooTumCsF/jAab1PsWciS+3BCnfokVOLwq/
A59nNs+r5nEvkeTWrKPLVMWG8myU9s3Uqe1twMDkOpvb8H/mN0Dn9EOc1BWX
dDqz5btrM4K/v6hpKreulBX9KmH4dxinGYECRqYgJ1BvfD3qHMCb7bAFpUA4
CTVwXrMrRjd9y1y7lq0+WXb5RkVWYvT7LAQl4od9a93zAvX6i1CJ5WpxZAyS
GyQU0Vs31kvv490A/6DP0z/peItd2QyameJ+XRYcpytVdqRKsA7w11vZkQoH
2EcdULkAzF0NnOwB/TN7XY6qpPE4H9ltbXIWZqjMHZwteR2r3OPTSc2JLAMW
hM0OCdzE0Y7YICKvVo9W7Pskt6bTthJXeFPFzcGq83qkzy/AfLxY2rCIlcGf
6DvY9w+wAtVtfnTfboWPj1jUwcRPDT0WbLanbEtY/Q+PZEIo9GLG6IhcBK9K
Wet+sUMshUTv6hUQtXJVoWl2fHJMji9Z3Ub/QJ/M58ZSYNJp8dCY7eCOvKAs
FX9GFr3znvJCJ3APa/jpJeb2A7QUr/qS2S2hEIHNFTLgalnf47EqEKsdrGUb
YZATpmn2EgWs53Mm6n3jPjw0Bq0b3EsEBoaxqVJXYjtyAb4S3aG3lQ/UgG8G
5ebyUuI95nQ9v3OptPzMM3bNIwvhSm5h0RfR5qregECdGhsP9t9KWkroY1SU
NNzcxsq+/dPwhPqM+GWluxMmILTudinJOLHyZQTCk+CJi5QWNQ4vCO0a64/D
cpacCSyD9ZwtIc6uRp+LYU79ArwdsvOZFat6GrHbdXQzWOTfzBk/Fs1F2Kl5
csI3IHn2VyrjrDIbexE1BR27zMYPb5212IgMZEeP8Xui6cVNgPjhr3GVJE9g
54nSnZGmPDCszWTABL0gamgErPo2ljGDcZBdcmvVoo/y+k2JDHv+lzZd7Izw
FuUQ+SiSCgNYJcxB6BTyhMAtC123wLJUubtssdYZKgVs6rgvnmqUj47VA+aG
5pKmZeTqMOScKbB6XY7MzSTkAlXhCMRshfj+PfOuiYJuYUv2PdbINXu7urTq
XxjjZUfQJEJpPOYObcOzslQDs21bo9/k0hzOFuFpgNjY3+5YYyENHHWwoWVK
8zqx0+Q0l/6IvnQ6+7mF+fvnU2ak/7Hrj/vQdMUYGkjayABT/yaiRnAb7sYg
ExHvx+1t2iw/uoo0PF+Rh5potq0UxCuI9THD6XJNlA6kma7/15YWdIr2okzB
bGRloTuDXa+fhtK1lQ+VRn2DO+H8tGfLBewCdt5yLZud/BKcRhYcGPZzIzja
iQsvY/1o9A5i9X6is4UItBoFHCFpPPqrZp9X/QIEbuLQHZQCywKq+jfTOpQY
sJuys41TctWsCYYbNZwHL4NT+hyjdvJlOKRfqRcpRO6Dp2EA8Chcuf1vdVKc
6M9H/CdOg9AECHhCRxCg8ub2NVlSlDD1hZmNtJGbtpiM8tg7Cj6e2gizqT4w
MSSCCXtV5cp4fpOsXrw8WJHOej2JyGde6zlCsyGsNim8JLqM4G36SEEK5nur
qrcwTz7EI8vJu9/LFTTkiCpMn0gSv1yGxUEhXm0XrvmZMfL00TmaGx1MWY9P
P52PomJI96kzlF7Xzp+h5soTG6zG5ujx6wsV3BKNy1hDgbAzqXQ5BhsjQJVv
Xey975QgFiKwajBCGurxpeSG23Dzp5fbkX2MetoWNwTpi9eP2EgebQ79Ktl6
yJ8tnT814YaxDk7zs6QW6PxA9LCoyx5hbPxyewPkx+O2zFoRzzsUTjRKgWuL
4KmK4gKE3WD45Kubd4R+DzoUX5blKD6qvQ0aYJ6fDSMWIAr3MymoMSFd4yvG
ngqurw4fxBxMTeaDRuOj0SNhX7PeRTD6HqMsP/zxhDcoQkR0o5A7oQjbPnK8
WnKmZH0h3jUw7Si7BOjth8E+2xyYhl1F841rk+E5DJpz0ejSQ0gj71UfZrrL
lnH1DFB7TY2QwlqcaNe7RcejYyITpfsEJt0mjG2wgyMzKiTgfxb73CAxaWXv
rSdb362xIOxBEgNi/IYMejnmPWcKm01wHhK2DikHAcaqVvxnUYpVGIZgRTm7
PjPXrdV6e07nrJBp5P5jvRQLv49bNZWdViN6g6FeGHX1pP6vFge3Udqvr6qs
jo3lGm8cAlRQCORbHAUp7twBUSAf+cReKDL9aoOgJwnnu4bt04uNI8v/XOra
TARsWPV1LyMqXjQlm8LCSlRYC8KXUTZNZbpmVHpEBFt/8zNvlnSMK+vUvVFy
dOPwJkOmBP2a/vaREoj/7PrrhT+PAo4l2qBdM5fD874rWVBxQpDpDkYzbnIg
vHyfSxZYWfyAvoGxuFs1yQ3IiCJh3pWBvcND/WqowVc0+mVNi3fQJfBfaJOY
n9vk4hPkOppi+hl6QWTFSUP+N6P/T9CwqvekxIfi3DCNiJXnc0+UEajQch77
jPSTG++X8WrsJzqAevJ0YA9K+cebQSyFasLYgL08tInYVO4nMsn79q0ep1Fh
Q1uwOoUua2Qq1DTQqYlC6E92W4H/cp2FlBQNXq/W/WZIQRfGZHDFhSrBebBU
qw8SoeJs9GVMDU4mtoaSWjskihQcp/rrL5S0iYWM4ezcMYeas/868Fxx5pax
0urm7Q8plMYGcLa7qIciI5ic3EXm5egYQhZ5b5Pp2vZp848VdQs86li/ziw0
WXTvSG+xjoFlyKy5Z0arUR3ay6dD1s0H4MHZd389aRMg1/Ja2fLh7c8eYgE1
rSYko9IgtipWToaOg9+p/lbfywLeCFkkuyRUmhp80Bx0TgVJ0p9uPm/XaL9K
tJkHHVfRKf4++ECVUVoJITZAsy2b3bCbOS9LQgcEdImZ9rDmDJNwt6Ll4VcT
0yQueCvKG3dqca8/ZDv9l0WltroHteuJ7qtNfsnddtDHzXZf3xwLINvEK74q
skyFYsbRkM8cgdpFYasNVFiOiXHXAokCFsCsyBlyK/OJFc0ICNSlGXtZjkUr
MlVpSWK4UODKL3ABfe0LtLwgcdIw0J+tPCyEUCHd/v+SAPzBX683XSwrdPUI
w2U257hAIfbj/92yU/NDl+4zWnvJlfIG5E/mrno19z0zFrYfMAG/mEUWTPg0
K3xM9nOC9D7egljcgN/u7c8pU8nG06Sg0v0iDUi5sWMjMJAV3CGXeYiA6zxq
zJqwGcJ+yaHLObWwZJBninMXluoufCG7eb/4fzD7MbgZoykXZ+5lYZ36i//6
Zah7doElboFybmPJbspz97NvnX7yDPZ3ecUUHnG7AY8DVVcuHK5YmcIJ+BLG
WrxTug62aqCFCgrcHa2Djy1qvXBnju1KTWMu2uHFj/RrZXSpMa46kq0qZh0A
m0qZPUNk3/ZG93zrAIbYLs+RgtdthQnmyxXXv4UHKebh+dTXtmx3o0sZvGpM
sHgg61qpRjCAioj6xRMywV3bVuMi6Evi4FCj0E4wXppxfqLewy2x4t2ZM8k8
oXapgsFE1Fl5KN+H2rjDYH7u+D+wG0vy+wOZPNO2uY6DqY36e+/bvrg7re1Y
fnsXCPehPVeh+AQazi0vMTHgblDT+MxnX9PVtHp5Lyn5rZWBBFXuItka+1zM
tOzGaSwvGK9t7xNcxZ5JJ0VCg/dRvX9TklVq4DKkv1r+EhICEF+T/3Ni4fuJ
NuvQDGGOz7JnyxPgY7MpZnGuii2gQP7m8Ulx8h6KuFDgj2k8MGKdsVSJSl7k
/TkosmMTvaT0Lwp+WtKBhnIEtt8XyfrNWNUKfcETb2SpEZ0zvpd4FnY2040T
WAzWjqFe4Xy1bpXBTCQ94jOjOpl8nyKhaqwQzCeVWatTHewcLnax8ZXbU8Sx
mvDy9pcNmTERcEbQDxQ6JUk6NdItXrtEZyS2fSR92ebCKPUl9aqJvVhekWhx
3xIYCoOAORIT8/zO75s+ebt5IPLeht7td+tmFZlcdg9Oj4Jgkpf7vtf2iGoH
SLAa95Mx76iJtM6svd9oQfLJsEyqsFoZH6nFhdmCNjB3skJZu2e2aO1ntZbz
qohluUaIGCo7lp9zVd0pzU/nsw0xrnPT9KbwPEqMT7znlNAvoe832QMsGMsr
2GbJKsDPSvfuEUd5gHaMYafj/C+NI8KQ6A+ezJ2ADxqmQBwdMVD0s6BUBY7o
pWgxB50exx8bFKVCnXGJ+GTNeEDleDF999RS1Q20jDNSCV24a1TCjDra2tnO
ORwXrBfoE/FI+evvuz3v3aMSDG7rumtxef05eL154qU8+CZ6UoSvs2P04y1h
IfmGjnDsVzflbE2X6PPrMQmwGd0lj/oHWxocqrUUTuJ1YaQC2pIzois8kVpf
QPeRGDRDQiUcivK+oB5t+chXndKL81TJqaDXZd4UFskcSVxsGWrO6fQW6g/a
xDHascgMzKop1H2karbz3oc+730HRkCjwcQjASnGEJfLP42NKW6r7sqTXQ1M
394cH8cYLfboVy3QT1OFVtk4PzbZYJI1bSCILgsxlhqy6X84lng2oPXqGvIx
3clHve4P6Xg89HzkhxXcZHNafTXy+D/rQfEaNHZwq6IzjVro+99bWFhDu9Jr
3o1+1c3/P+IKfoeqUBoPslPqbZdrrF94UOJGh7MbrM0A36+Fik0MCH+H9n/8
+GQig4bcxqzPbHeui0oimDbjmHuzYMecYzmAgAX8cc9R+KQawCaToUMerI8H
AkZfQFG6P/+2+6XCAk33PIdcfNofhvspHudRPbnkjKRqnQuex1JIZblJlKC1
IsDUezRom1KXB6A5CTLUjvDWN0o7cZqe0/i/1V5l+0PPTCjLaMjNR90rz3Vx
lXKDXSPB5Q72UUOxPZZfd/pNSnVtZYhEwoSQyxsn+46N3KMmp7QI7K/CtGoX
nA8CzOVoLIlnmawvPEt73Ut869XPWRmsUvVYeeNR26wdbp0QAsqBRstfutMf
s+R54Rfo3IpZfYu7Xn1k9OOwenGZ8qdQN9wMHpWYhww9wpX8AiKt6zh5sMMt
1afNamZGSEdSAAVQPeLAlReiSaPxJoKJkdkjUr0cgb7R/w1ByUnK6sIB1dTI
IiQAYXl0dNIOOkNykAXXNuoaH2RXvfXXCw35bHoPJVDh5J1HeNCIn+mqjlXS
j4HuMkJ/aKf1P0uQA/a++3+RjnelQhbeqjcCSNbLj7eM6WeP/I4+8+NVkTSX
+o5R5nEY2Y+YjRsePWNqkdlz6WtYt1B3Zo0ovqq/Cf91D9E8LUZQlzjCPW6t
hlgs+XH35RYXWFXIcLpc7MV0XGAWvXoJcS9znxHCJdhYTbcb8I8ublnGtl8t
4ufFfftmCCh7bDym2BCsfQg5EN0cNbeyZPVXHrqim88EN62bwgrTZ+OtrCMs
XycSb6R4XoK5t7fzjNqfZmJKun4J9gT0aPM6ljKC9dr/5FrZv0l0h3D+TuPC
BYl2+XmtTLgwPAsPCy17tD8RCpz/EMl5/DZbhURYtCkRx4nH+OJ7th57cdaY
Ain1ItZmz7GUnGVv6O97UYI3Jg1Ik5LlH84xOqNy7/KmCzKKheOm9lm3FjTF
qellV/dAcDef14fJt/orWJVreefhSqDbjcz1AiD6iQq96K/SlpI6EVXnTTrM
6dmWY7m/nb6B8Nv+EfBi9TdfrhkdHtSdhyu/zpVCs0NMxW83S28E8ZhPdhlV
z0Hr/75fWow4ftAcJcH2nQuqFnUDDxTfGnyI9r5Dm3rfCjaqkPYUF0NN/YuR
LQoQeESeGPDR6RKC1hJ/Mgmpzy80yEEiZD2t7uIB9YRVzLzEDHqcXw6WaBAg
xCR0kZ+763Tg70OrycjZRRwzGkTIvOWe6kTxcocIag8lVzrjaQiXXZl4g7xB
DqMKlY6JgBeIh/VELxIJVUu7Pwi69FgjgmsAtv9ruMdhiGbbvKoQHPkkPLZh
vFrRjW1TCt7JNVEdhvLZm/mDORzMPmX8lVUD1U6xTrvy2ecg9C9zl+xXCiDN
IZ0gAEVK5QbGvNJE04MK7gvocEvLA+DpAZoiAsML7+lGW3XDDk0IXhod2WTZ
+F/mOAlVC20B6UZ+a3NqYW38fr+2mM5lGOtl4qX92iUdZznzlj8aVx+4nduO
2n+trk4I5O4Iw8epjDlE9VyMxznYBDwtmiMSBEC4nCJeqy9snUBzz65/M8dr
s2BD9GLxIHIXHRHcg7SBTEPCi8GegI567YBLaVN4yB0WuX2Lc2Dn677tu6Fc
aZE0ytErLIxLcnx7EDPKj2D+Q1w1evTQNWZljsG527i6T3/NsCEkxGIPJPQg
ND5rP2F0FKcFV5K3dPWBccuVu3ftkyHrYnMQuV3XjAyy+3wuq0tCcseaVATA
kQSk5JNZxh6EhnnoqGIkyVs7jRT1mVdjazuMP+K7fCTHjUSivabizo+7vGWG
o6qZXhQdPaD/JtAdoDTzBsA1ia1N6NxbFjZrv5blz89NgiP2A1pkdZgjdpo4
bLo0+M0hGE1e8chji2g8IVcLD7lsw3A6VVXV0U9RasajmxLl8E1VMgC3NMvY
nqwMu4VYhSHTFSNgTspZLwolyZxQ9DOtoLMslxYP8OmfLp5rqiZTh8Yji7iu
XE7V8udaoQgb4vJOks8xrZh3Yv/N5ax5DYFRD3J5qSUHUAy7WpCODK25niky
/y23g6vUaSkmkC3uMgHLi4+inuMv0tuSHdcp3U8CGhugkP1np0e091G2uz/3
rL8BDGF4PX7N+WAP43WJrcEze7d0boGCALbMRkh3n1cis5MszbYju3KVrbYQ
PFXzE/GJbinSdoBq05bSvNowcue8cu3bh+lYrrIlYRc9C2rfOkQ3Nbg5wF8r
c4ij+5n4VyxlxLVYOKkGfRaamGb6hc4lz8qFfapGHrrI3N9vSRWzq/5HpZ1u
1bEiiw9CfPCuyNX0MVOg/DV8lEs8VnaD+JrjHXRlRsZcWRolZa7uSwpC0Q8A
wi71E9OEnGntFZ8NbMQGYNA2l2Vldy8F98lRnyFPVjn8oyAr6wwZfPpUTg+l
AzxFrumiWr5ureEZ2Mkwp1kOLnJbaDn58bIoDVVJHvaPeoAU1SwWUAov+PXx
i3DkUzZgs3hgeIiiOdKszjg445XAIx+Ka5QzqYw8kmKFCdhkFEt+BdFHoKrc
wCWN/uTfsZn5d4rzxm498PfnXJrS5yiuy/SOfv7cBm1dymyWw5HCRYhraYAL
Vyx8naeNUrk6GcD2F93zzqQnCmdu+H92QWjOOnsnC5AgsvksVHLSyd+HuK0M
Mq5btqTGTAuu+aOA2dpA/iUGMCntb3tl/qUWhq/YJKW9rxHOGWmkSPNXTuyw
suQHfBg9jRF2sVP0zwdngQboYKYrb0fDFo2tAXv9o0PyIrdtgkkAeuE1/Nsb
uCdysTq3AuT6jZ1rUWwONlmRUL5My7m2S9VZYQ7HYopkEaO0VL9KE4qdZtie
HvXTq6AsPvG9Bg7vMXXH2nZ2rbBIUGtlVeGcwkhbGdluNxcGw6Ywm1NdzrWJ
3Q0wfD25/pHvnQfdMS6craCpa+qgx8fQ85vNUIalVv2/8d2CEPaCDLBDMnuI
2SB3NLnlZ3zMiB2REKRKegNeP0/oMayQ1Era5SnY/YW9vS/gbtd6DrLPzxr6
Wi2EATzYTs6ZbCVvFQ2DywY/0NMEoRI1Qk9bDU2md83F8jweiWDh5qW+Xs+r
bU2+VM1V/ibLoUDrT2sx+4uwXDKRY08bNk45CfYbKVSDcs1apikV7Q+IL17Z
zwx3hQuZ0Qgwwk6mQFmmAsK6q2TpraG96wxgf7zgeiByYofy/nMwjMNbZ2tT
MLxjEjQEqS1g5b+FoxVCjhj2//+xzNOJZPEjRrH4O0qf0EsNWuxkOK8bFchF
0iBTo0/R9PE5eFsxvpjdHT9SUaAT1jI69zAviT9TI1YHLQQChN1viA8m7SWj
dO5hmY5tSq8ehfVmojhCz4b6S5nuGuN4nkKryzoNBbKT7iiHnmUGazy+MKbV
TVe8+wgud3vyk8nzvQeZQ5l/Bq92k3Lmvs/le8UCCz/upD8UM0pxFwt2GdRe
aHxIiS/EDGVvlp094AC5DXeKcwCMwIBCeVxiAqY7Osdztip/pHzOh0/i5khp
c2ZySfyxLw8BgzP/ZGi1caJ315K7jbnmMwp/vqO+9ismii3Nw3Hud0mJWNbG
YWhiyzg3UpO3/Ww93XPL2D33d2c1oKH0DCzQGan3aX8Ge86mMcyE1q36xTY1
UQDSgdyiFkbF1TPpQDWe1i3GZ6eYWgDzSuxX0AXUXgXSPnMyYfB2Y7HxjRtO
XUFUlQFAv6G5pNAbVya3nAQ0Tm6J17wMsh6voqNednU8LXScGN+ePBCIgXI5
nQ+QClYqU4ZEzZyuA/HwY2Hia0sJs5ivrSh0zHIU1e2bYCrOG0UfO2izhGfD
rAZw993VH0M5p0l/jtUKL/cZAhn0epHiqMdMHBmur3AX4dKORRO/PVCeJcRe
9oTLs0J8lnr5FkXfGOQJ48yLYeSZxU3rlK9J53KSsJKthI6qC4FjvOPBIAHO
ryktpEHlAu9tDn2UhlgFstazxEKunv9kgaYK7uYft6r7KcbgsniM2Y6+52RE
Ra0lSmFVyak212/OkuHpN31X8av+oJoFzB6toh1fz75eWaMcNOoyp5bBc9Cm
qsr1NDinu3y8rxuA3LY0YuuG/XvLQTLR0Nt3wFbWrGN678ruJpqzp7AjB7ZZ
hGArGMbYjmwQJcF7Bv0nrYwuUhnqUIQmAOI1dPSzVb+4bwW8HW6zJrhqG972
Sqbpu/KeK/XUMDp2hOiHXIfR8xbADMZtvjrbzzfhmIru2IjyM9pigzzqLmDJ
rbh7JSmxgfBgFEf14GT1DNns36unDkLOwHbVTqtHQ8/DBxXmnN7FdQDDJO9d
2LdW5zLsCiRLcJmzacDeBWiAmT4+Yt6VdboMJYHaO8rYrz+7+sskoEps/RkS
tijdZp/tYET4L5ol2f9qEWC0sUNi2WpFdjjrbS1Nho87ReW446pFOr7vSm69
Ez6Un2gII83CfVBk7jnENt0WYhxxUml/Bd1ZlAtr1UoD6K57WPqBs0RYBpeQ
64tOA8l09EHgrZ+RcGbo9rfeIE8K5Zy3vf4d29y3RkXXzkvgQVjnXnb7C5HK
gBoSzzzCJRWnyR576dN9s1Si6bfRTnKrjXZ4tuy/xexT0ZAg6o4Ge8MXcyB2
1giKPFVeFR/SKTa9Y4R+Y7J0dp13jxW5HP7mL106G01uqzzH+e9QONMPBt6S
pWrUsGJ640w4Rb72WkW9uBCYyGOZqOV2/0HmkOjdaGyG+b/dP4kqCuzzKxjz
Hy9wORU3oJMlm/mMUz7Cqp8jmVY/cPxJq5XtUUW1CGbZfiwQMFev99rDFaTH
HcDmLDfl7uv0GSsokeW8h+jA8zsOGSZjQly+Yf4XWzHd2ZwYe0z4Pfnkt9MK
oAKOWkqF/tGfD4GnTZEnU2sJHjYSVHkYEBScASpZb/VO6X7QjUStgJnHyQO4
tut93TA6bEZE75myt/xI7fSNqmv0MXnZwkMcw6QLSJF4M+KQKVLFYxHEUih1
dRVh0/jyjVNo1BWokjV6dTKQ2ATncUWYn2G4uThV5mHyETJV96iGxC4bKuFQ
VEBIiqDVut8MWVIuJAIjqHdr1szbfGwJ913U5EvSMfTg6wYwJF7Wyu75H6UW
zowQqyc8JbFpd+cqYyp9bh1sywV1NfztWdbymtieqjT46AeJKf2VlQZApe6D
8sOr65G+xEy/a2p14nXzOU/0Xp+wOkYm8r6JyOjJf0Y3WgcqxT2nkOV1rrIY
EbGTRH8XaDuzN8gx4u5vftFM3zS8ddKp6ozuaLnHT46YEZwffZKfx7OovH3N
SX438IU2dxWSUTgB0CUl8Qzj0aJ5jgK6x66RmC0wY0E8/K5UYo6los0hgK/L
B0vItC0XiboYMv2aKAXh+88kfDjEoFlAcryQqi9quz/vvxOmOCYQiqRKBZG4
4zCDBB2SF4K3R+lLbBXLw/uT+ccdGdDWFfvsbIbeL1SBmeGI9w4NTljkBQQU
8zW2lLAoQoirCXl08NriTkaXARZkxrfj7ZVxoIYGvnYvakYpgeOHnUVPo8C2
KKrTCKw5dHBdvukQ9VPsFbDStfFB7S+6OvvcqE+t7IFQ7kcAjDORykASZM1j
/vaWOk1tVpYzFpbNyemLBfAXVTawlVH77BbU7JNLYsVXdntYgr6Vv4b3cZLC
m4sl4zkyLXQ7Knbr1bdlsKFuPeWpqUEz8tQvuXsGv4uUs2Zhes4C9BgSX/VI
XtWqdPIcqgPaW+Lt5ha5EOU1VnTo6nPB9FHrAdfYgL5gkc9hQQRWkAA29bMc
9ftnQLLvTlWHgmJNrS5vPztLD9s7n8fLoA3YVyuMi+3rhHULoi0Xm5u7hlg0
0dRkyOhDNogvVnvKo0r/FDXotul9BH9OgPRHMrNZsFnfo0obP05gWfnPHyrg
HSovfv/XiEDDdtrHmcOyN3cnrJ5Hy0J2Bn2mYuro+/dqpp8MUFtgyBmMbPWd
UgOjQ3qFoEo7Ap9mFiUjPY58BfYJir/knEQf/ddw/bUVinOsyytNBtOpxOKC
DrW+RVbAmm+W61croeocTsn4lMmGzOLPteQ2+RkdWE+WmFiqyF2lXf+QyrjZ
2ykpkI1U8W9QQdcF9ZckVVIsWqPMl1fRg1XUIdILvLLOLvkCzW96d38VPoCp
mmUw8zYAvpie/Cfh3B8Y/4VIufSctYqZSD3fVpphqp5ijQeMQOyHjQ8CEwK6
jrUK2XKhKPlsdNwfXFk2HNLLATFndr7y2UyVBNY//bXjcXpQawgpqquXPcHo
fHhGJKl6osYhz76tCe8/lQD2iWXh0AbiDulMucDmYaRdlgmkxmFC4Lkyv8U7
chg4HSMZ7yOO28S5JIShNBd2PvB5JltrEF0qtosyySr/zY1e1rjRLJM+j+nA
YN0mvDDSZlU3x6kFnvXmuB4kLnOX4HQ+lWt/2vFoD2G6YBDNIJOj8+55RFxD
Fg/VkSiZu518fPbkzTFAW0WVEPWMIgKV7+7xd9RC/fsyjdl27dpbuFn9+TBs
f23EodSUpi4JnucMqQj0Wr/WC8x+yI3pK5dcT0vGGenU886SJcy1ffEIHBZn
AlEXnAjYy5/rUeaxkMKV7ue83wmjJ2kmXWNBj9PVmx5ixrpEE14UfElbeajO
VLSzr1io8hl4kB1ed6qwEPjgmGDEmY32fsjLi2OS9pH1U4Ta3jxxrUKRxH0y
L50e/3cIBx6emevx2gjbfj4cB1OR05Qu01/cb9fXrxmhWXqDanKEku7lqMMc
2PaUxBXzdYGNG7L1SISDc54//ManbE14peDI+65lvktdImMZnMooBCSpLIrx
L5PYfCyzBd+CuVL9BzP6TJUGsJvKECQkG5iNaYmyGytISez2TlrWebmbMh+k
PyhANcpB9Yu1Htg7nh/AdZ6TgMscOzRzWVHVSs96TZReuKbRyXogWzYbHIz8
A30FHXIhlYypZ+dFQyp1Jw+JHVyQW0uktyETnuWbYnXuVIyQaa1lb4+eGnn8
KDqRb+ZeWnWkFAMcTkZOPfwddCSkZssXU0HJ5bqZULT6T9Gx4M3ado2URMzj
P04HKtNKOupQLIpe3/5o3ZJLWzDkDga2zP5ClgYy+EcHFqyTSv3k0ebF9Ln0
VtkNDWpZRJ9yWiLlaRT+hX+0nqTYYJmoMZJMbPIfK9lDM8hIMGCsSvxD7Fv0
XjWm+ud0ewOPOsa2VL5d+tIiNjrGwFeXb4QBMZVeD/67BLLKUoeiTWURbcY0
Z6IhLfCiePn7xq4n6VnM6neHOa19KoN8Ic6iI+EpdX4ECpuKADooPEuSflEN
CLp2eHJNtk/qNw5wY4I9Gd9GkaZSKqqD0XIzhW7ZD9D4Oh9Y4hLOOHXJnPqB
5cvjm+qMJMfl/sm7IQ26IRdWulyJA/bpuOrzi2Ign4qgFUdmsptwdEwXH158
JGY2EjKh6seXEw5PYmWwBiHj5FLB4v1TeD2a7in24XQCqrsWudl5J/seZ2U7
Pmg1kRS1bL0Qk3Ba79k9fUCexmkaZHjnkStvR1Jw35DuoOGQO0OBlUB6fJ+o
dhxalBu4kqf4QnfKuclbQRAa4XR/TIku9xu4kvgsABCx8cWhXs1imP1Tledh
ML1x6C9p1t57r76jCzjpCNIS61o2vvV76SPomOgMj5KPD9nguEZuGD508z08
ay6YL6hai6NUb0JRrLGgKaKyrlQquvsWVLVrmQaxvgAIW/iP0yX9azb2RMb1
WzLeUDsehfI0UCgJcepcBZTFMwuoi8qqsNrnfUyq3rXL64nRnYQ9nRYvdHzY
BrKo9PnPce8drpwgWw/ZtLLWq6A5cXJzT3sr35Y8vQYSotg3nOutTZGBUc+1
sa2itCBwR7KVmy3TmYewFEsnORY4etDpeI8s6anX9+bcCI61Y8UuzQsl38mw
amNqdCxZWQECmqkEGit4rFCMa7wLxtwHLGNM2nP4WKr2GVZqBXCG9bvfts+H
zhopQGbrINM+HQJHrGMa39iK/CQv2rppDame+dPb7rb9wE1ddboGVbzoCMmB
s4x08/4q5cQfhmIW8TfKJN/KSLLgAPnosvdEJ/CyGASwExr2eRnHsAWg0X9o
VMNUFH53vLD4F1+U6ABvGt4FXDTIZDpwYaCCdXZ1pg8CKJBX115w2mmWJdth
JlrP0eh/ljRi+LXQnqLmZJr1LNqkh7WbLUHjYAhGxADfsopxb0HkKEAWV8IR
DpvQSUYZlVnXF9RHkhby+GG54Hx+qUlj62v8UZYse4Gcxj6iRnJazkOgOfw9
7V96b4AM5CK2/wFB7WD5Gp4pTcWuLTWEAviwjzB7QgdofNC5JWzJ0GbzCiO+
brCTCRco6lAkeuBbHET0yDv+k8liW2czxmh2KmhA3MQiG1NtOIjkwOGcQ3Uh
0JGjMlr5If1NX+QbsWXMXvSdAuT2Jlkz5WdUHOOx9BnIYUUKKubs4gDezPMb
q+ULFOiXlg7dQi0X9xpcLSWnSf+0ZMPEDZ9mIzsciRxlhDedXbM1euw5vlxn
a5sEYKX2zC2UBebaQoJfybCf1TItC+6EVn6QMhUGUNKKc/FTLzSaZO4gVI6l
Zct2lIiL5hG4eonUZCr/ZyjFxP4QSm7XZKuZG22r6bu2uWXyRgYXL4sqpq0v
Fkla8Bt46WXDpQi3r/SCRSya8/QWBJzVxWCYyM88793AFvplPKCmE1OXelJS
7CN/Zw07Y68YSHcVxtXSRkiJuXhb0eTudcx4XLnHawXcmBfEx1agcDY17a5K
5O+9uG4e7BUJ9jY304SfNmux4BtAqWBkrkukx0akliKmZz1QoXFrMIdNO4s0
eiXR7O1iAnGQx3GxV8uSyCr7HHYiK9qJl7ejS15MHHtay+Zu09v9E8jTJ93m
VhEIixldIC1Zn6P1njr2FwJJvtEk+qlrheLKAh9gz97VGe7beGwvToepOwYF
DsniroSCp7DkMG7f1E9A+4sevHuN7PrjWQ1M5Pklt+3A+hDdVVu2/dDTKfVQ
LKP2/FgkwXS6anhB9S1xG6pMt1TrYr9m9owh829oIcIuuTj6YopdNmDqMfjf
Ikg3KNAIzyr4JGrg9TcEQVMrlNqvJ5rPAan8j8kc/3AK/c3H4seeF3JFJGrq
7icHM/Lsyw4ALSMpOFf0uBqhb8wEFBUkbeekQCfdo2SYU7n3V6ctuIZSEooA
CQs9HoIAyt5ODyVqoTuuHC71NbrOFWfmtnv0uf05p0WUfwJSph91b8UR0SLL
W0hiUI1YK2iixQGMHji03XhaXK7uTW6krbFR1KurUkS6a/BO2t8iSgqYWJEI
rgzWtW8+KZd7V+UwoR21W64GbBCV8pb+upoTnstrpJwvsD5Ebu7j2lfnOaSR
hJ9DvBzXyrBTEV4lbx2ABDJyUF1VrwgPfvP+/r8TQIQ5TZ5iK1Gg4lzDE7rL
qUuWAfj9h7h0zzrIRoNw1vHqwL6u27RRlHmxYMfpYeiTbqrNxiuG8aToURuQ
e7A5aTPCThgQcNGVVOVLFupuLBAQdMxeyZzBo5AR8kH5Ni+32ureUxbaTLs0
vHnNuuL/sAU5doFs0mnrogU3hACuVxjIkJjlKuq/BqXaX9dkHiNnq/SU0bCW
QrmDaA1+eqb4wvh5oPmzC0TPOHnDeeVM6oCCnpm1J1+bclwbJVosytpDChOt
ilqz8HKbBJVJnNLHMy6guBQ+etMPBsRtquRYWpGOTS/ySA8roeAqzE18lGs3
cInBmLcmMgjSvRIj1sloK60cbt/hb/W4Mw5QrJyii2ys8+7CdV6LX16+d/iP
V02otl2qKzwzQ/yNk6A3kRgXHaW+7sHZOJgZxuqo8BwBcSytcGxCZc0Ptrj5
eiGRid+34PWj2VX7SF8DdpeHfwdrPUTlI/1BtgdJNThJ3KwobDOayAoE+6Ft
Qv+oeMesxFuKL9a59NWIpWZfxe66lU1ufTvTN9v72jjhOGuIZnqxAHyWUooc
ld53cwPB3az/drJFPZzecHPGVdJuB9rgRSZQ5zAOPcFxSwysDvo68js+wSwa
DBBMMBHipd4XJM9ADgH2HSSuvXCW/WvvuIyiNnKmTIyyvH4nGU0zeEfUoiOv
ZeCyZbqC/YgTZ/aFFTdbCdWajsLkny7RrjJjl69WY6lS/GfVGYWVkz3PER+k
0n/TVZC7NRyFfM8GWpNzENpnGAnTzLEV/caLFqVMBP9tqxkcVO/0uB5ZQtoL
BN+lhpipyi90090ole8IThdq/gDqQo2+L1YTN3C6gJ9rZecuQnKHhPNDBElq
0zH8U/pTdDMwz1vVaCjeceXlOo5V01HfEL6ntfhzdSMUpnQJmhoAk4URqzKe
Jz7Hs5RfFy+FR7lbR5BUcupvU9NJFFUrZtMQ/QIvjpNN1M4Xkc+8UpC+B8t4
+4P+feLgxc/PImiLidvurPt9C8qIc68087VWCIHmtmEEGtT5XqigXr+tfAXO
yzFJdUyJqfM3JLGZUkpooYsR9EO6hW7j8Jd465lnKChlLo4OGuRz7qIVNxEx
2JZ+fr4CDWIh9Ljwum8yxeX+x/ssuyZpKe2z4IeudlnpK1HzGbGhs8v6I98v
CaezsJgCoBj8RzAdK84bpBOut95UUyXHB1opHQJ+BqsroQFcoulBksG+l5HY
lQRbvSXtWuJNFVfLX9/PQfjv1OMZvdert308nHWVSvGIOpjJBKF4R+Aj82Ej
BiGpxtxMboUH7OjTribxzf8RIzquIAwUpJ9pG+Wfw5ECpxV4QnNfJXLuOTMW
COs4ovDulhqKVmNxr95ksH7DZKTKeQNpSTypzHFL2udco2VWo1THc/fvDzae
QkogOhdKX/cuRG235tg06Ya2uVHwnildvW29b58Fej8WNbz70c3gSA8mLBY5
MCpOk6lD0/QQ19i1QlWpZGeCLw0NLUNM50Vf40VbUo0PU6rjyzBl40EBQBNi
gvRA6UlpX8BEo/qK2MTGXBE8ItLJwsShKM4kvHyJG84v+cullv5MB5w/8fd+
m6CjJ3BNQoipthHOKgNrYKokSvpP5O/p0JVFRSSDNpiRge8VFl80fVVS6FIl
2T3GviQYlZO5fXIVyf55LNRbWrHl+HR4MtzrRBwrPn6lsPyV53TKx6vJtHes
d+Ts9cjurBW2ot4ylFOQaJmU8t+3/ib2NDVQTWrKgEtMMnmh5UNgfoNhMMPC
sUyGMbU7ZYbmNHbVDBamVlxd1LZTtxhyiqKiWM2fBCJC9n4DvKLccr2YxMUr
7zpXpD9h4IbUHvBP7SivMoKmZYXZCKwDFCygEgRmRxMjdgJeX7zZk1GrpGHk
Jr6E+Gezb4uBdwj4MlOHTYC5RdkA6cyXLuGsihgz3VojqI/jRTBOXUuAmGCH
taIrE16qIBxq1dhH9b+kWdfOrzHrQNjOGfZYJNfxn8DUhPD4+FrVRRvWLcOB
a8ocO3px/ndeufakTH8Tl7BoqKxJBfsKJGFGglimp7i9odu2J19GfgLQc6QF
VKl5+FHyr80WM6vhlnzzx6YGiih85+JpDlq7TQymF3bOYZmQPujTSvJcmhkd
gd40JLqL+tFQ92JZGRSK70jnuwzJepPuxoEk5TFkHXowFvRbCUbcU1E5oXRG
0hCHWVyBt9GT0W9A5A3XnS5dMn2+skwHuhipWr43aQA95G3X2nEtbXadW6RV
NRev2IEegsCBcGwVD4GM4oUD3Y9g3ubCgjwGJM3E7oM0dzRLIrQLUe/t+9dz
xFOlC8tXp4PjcR5kcTgXAaovoBa8XC40ojI6vHvA6t1rymnW4e5GQk4O+Oxg
iSDesVWB38BBBjXICoelSUWtDT7D31igfKcDvqzqVHnreYHw/CRe5s+J51BL
yjmWTLmuTz8Evg4j30O4F6WCp3vKCKGrGq35rKnsWcQwOE/T5KY3nH1kqEsG
FQQqCet9Ztc5+pAiOd5xCUypSqxI/jLWp7C5GlsxEOHxK/tHsww6/4WA48CB
fcaTGwNB/3Bdb85YTssZIp5d42ZC0rYuVKHx80nvdCAtnp+5Wrg3RYinyewS
D0tLONC928K0yTabNnsQGHGNNG19AAOhkJ6YL19US8on5rBfPOZMapD6rUMR
zRE76wmsttqxLd+JrfuzjizbCVelmV7YuQrIYVSATgrWKSBsE0+NuLVryB0s
zlFQs2usDpfq8toV1diKy//qQyGvrLzZ7XjR2lDNzDNp38VPJ2M5PM0qz8mV
03djIynhmqmGMzWEy95K8lDv+sMbKoJVjw/I+EEbhA0Api7TlfYl+CkJV4lK
ZwwSLcKuY4gmasRcNfczDEO3r99wwbgkbCdEq8uJJCPVj8Jct9URVzhGObR7
Na6EAPfvBgM+uQjLcahk19hS7sESGauAdXXuH60hojQabNRCTrt6TDuGWBXF
fGMDETw6h5yBMDiu1qVuuvhl0TvAZMMK3tHIS9na8RT+VUB2FUqyH4E+S6YW
6xXKSYdnTiQmB9RJPBmVZC2favZENwyzi3zDgNJ/Cr+YIMBOyj2g77oZm/l5
PfOUbw5XGuH8QhBpIp6gdTwRh9CvUVRC6ybTSmSmIsKyOn8p97k5DDvZghfl
oIdJRqfaHrGAa7Xz9RP8OsW3tHtXJmMVuVr1LoK1Tx6ZIBYsXmFqmYfr8R88
mb1Jhf+u/Rpbdte10AtiVGbDvLBgru64czTUKGUZZMl+TEaOWLPrTdAQNyta
cOp/zwsiH3bgMZqBNQL8Lxxnb05MShNOuLCIUDXv7Kjq4wVYu9UlqiuPqTST
r5SN/7PeU8P2b1TXCk746VOYwHck7XMnNg2eYjviDJdsqLuZDDO7oOjfQrzl
oieUES7Qb5gsQQUQCNf7CplGoiMNgaS5V6TWBhuQFMrfZTzdmw/OqZVu1gTr
drS8WQ2W12+8CGxCu7abH5h7WcS2T0IPCPPKSo9OcTbP1MDpudlEJvUIZTXR
6Hv2lZ3KkAwWZHD5CRa1HmGGa3G4wSdLOU9gzGYn9Tdtiw4VisQ5GEzDLCYU
fPMd7CHVCkIOEbDVCAtHYbfzyUmkHHlYPwmlzwQMkHlIJ+T/KlY6En4O9PaR
5rH8lH/nYFluwOOvY0YdCu2kfMUbglOgtfbZVkQjg4dDThuAWUKs/h/lJ9Jq
cMaV/ttM/98tEpBqP3ChCQC4/QxyY9AfFv9M3erXzaQsJP20XSjpQLHiUnRl
AsPq9Xwzv92WXSHTXQRBIlKtywJQ2+ZINTVBpW+Q7jV++N+iZR3hLT7epUwS
5zrOBZc+fJHMZ09XblfV5y1uEZaCuoN5fXyEZ9YbB+WFaF8NATkisYBabhzr
0fKwEEUpYKadghc1yDS0byzfnW3f/cpkDtXe/NFafNH3Wpa9U3rl1qIvjxaK
GQ4bOCeSvs895Cf3HFb3z+gl2jhFCqDcc6USp5IzxYudSqrQNpxUy4XbU5cI
BEvnYMyGNbZztHymIFpG76KyoLYwWmSvTq7+jrXxcTeK0iuTS/zGiembHaiE
PBU8USWc67c2kpPHdDKLA173UvYqcJ3mrgydKj6y1LUWeRX/6M9U6M/LneKp
oEk3L8ZeYEOq2fNeGG80oEIqZGeRHdDSXJCe6DnhHgwvrHx8KlNII2RQ43AF
hX9ZOZT85mNV+zle9Q7A21vqbPkqtJ98QHS+S76E1bwhFcAE0U6dvbuJ4ElS
0T1QF9g2G9wyvpyU3G0kAOWg/P+BvlDzgtqK9hLpnDkFUmeo25zCfceo4MCF
et/K96dmZJ7ZYAE4hiMgU7MQdVkhpYEn/etDaR/G7UcqfBM/pBhS4MQJ5Kxv
QAKuvmAZYYGFz1PHXauKZQ71Lbh2IICfADXyy2Iq75Y+GePw2OqLsDwITpau
/JcGlosQ1yyEZ0+uNDUnJ9JnXTgOPXqUJ4fdsWiyikKsenm2tSSQR2h9A4sd
G1la9K2tjxcfpb9ACPFnE1+JhX6QkxbO5s7TqTVnse3eA4N7UmVAST5ZztFV
uNTQYXcF2tgitT3pdtqhH8AaLGY2jK/zrpvglc5g/96+X1i0h2D+2egmNVGj
bjTjLbUbqTuyC30U30hxGK79p+uFVBZw+nlEdp0UKTW1qpq9jrKDOxGG+OVv
s9J5m3m9/94ePcIi/sRVW5xrquDbhw8XdkU4iBd3NH+mpI6vyOJK1xzUyBSr
cshjauVd2hLIRF+y1WK2zFOMhTE8ssx3/wS5pbv+O/pd5KH0ma8lurZn8NZS
GQmK7b4fllZyZziDiqjtlYm2pTBCr675e0Y70ptBzeR20kIRLBCXmO0B6ug3
krAbLvfNBR0iD3+tU80FuPDSCsDwGE9JOsw5+Cq177Fip9OarQT4OjiIm80E
FIJtN1Kl4heM0tGrX//7/eU8hAqRrLksfZAaBncEMIqLEisjuxI+crSjHkqm
VPFC6oXSfutpn0hoINDRzEuvFhiPuUA1+k/MpXPKRlG0UXoz6nyzTpr8fulF
0vUu7P9Gi++ZYAbxV/hIX5yhEhCbb3/ymvEF26VWJlK6H3C+8dqw7Glfc14f
RFD1DFmqlpz+V1ZMLc17TYilnHy22lPqXDs59qvfCibvEZ8Ieugr/aCImuAk
12osRj+hWqomwA4nr+wSN4UBLGRwhoUvke/5BerBgNJS4Xw+MhIanJY5xPCa
UFlu9jtKyfG+GooZDaKP3EYXa1Q1Xqc8tA6n8MHU6Sr4+HDZkPhljAQicxZT
DmhkgYDvlCUp7HXsuJwOChUB6+8yN2ESoUYrsjPZ4CJPL8JXcE/ZZ3FnPd9H
BdUshbtCB3byydjHhSTAqzvMX1ZItH3ZCwPc2KIiz9FRCZ8njf01unsn/5SK
EGPiFCVXUQ/za2JmWRAFjH7VCvKPYLNhJVFYnHUmAIvrQNwuktO4mbXtLj3Q
grVgHv3WkinRZIBQmUzDubXIl23B1Snj5CH/IFhG5cHsWroe5nRkTvCDHmaW
u1nSYGwYDZP8bVEaX0ulJ8TNI2mavCGrb5Hlf+7vtU8pCnK67g27hMBcih3B
3TkS63/81/xhJ3Iy0I4jCMuxjLzWNNvRl+nB2609qwUYnh0ZyHAxTLDelDhd
dui6/YFi777NyBGUDrvNG5qo64IxTufacVZCgdnSfRBjZGCUb8ASFQuK6l68
MC/BFiPeyruWxc8VmdrpYxsYwXKf8RNUnh2U5VJ6yg6MJ7AlMG53krZv9MBd
N4798e1eLW+BvxlpyJU4rqdEmUk2i9cj2N0LgrvRQYdmeRL4a7da61ckqQ9c
I4tLevtEjhGIE37oVBYP8tg3H6M4Z5a0Ntfuc+Syc3YIQVhMQVLZ1V6IbNtw
s9zLc0y1x6itvnmF24j0TKNM3lWOiwL3CxkVczyPsmlfluYm1k7YSeDa3Cmv
LeLAektOdEuYLZBozBbOGlDwEB9YLM/gS8kO08YgtovEY3V4E2pD9426Hy4k
2s/0nVpDZWcYFF7fbkRVSImYsZdrY41WFuvcjcNfY0ActKKrQ+S2InDf06xw
/OJRBVxY2TOJ3u/13rD0V+sjW1eNzwcOJApfSEFv3nz9/uqvzABm5DVkxP6M
THsTAetBkCCS9mGCeeZJmUNnNOkKdCkoTc+8xkrhsauq2L6JRRBLSTV8IH3x
SurdeKUg3m4RBYpjzTMlT/AyRfhbdZSRhtyx87WIlV5BFvTB6TRICBMnL5MV
w68KfJOjEp2H0GSZMUh11FUHll2R/0qg8aRT8gT2XFMIiC4JMt4afH6hqxOE
xnvVtnqIdj/ACftY5gwjIGYRgs8sR1zNLmwnp0Dw+GCPcozkjUlLLGie3p9L
vnCqFCzNf5PXk/D4og8VQBV+kxeLuwl4ZMC50z3PdCe8mz3Lblj3KtOQtSAT
jrYIrSBreW91opP78UIKpJkgYz75YshhHi3oJi2bZDXVCFpVQedWZnoOwk2Z
tfCwRyuYgjzWwt/lS0ptygIy1oaqC+6TnAF1Dx/F+Qw03JHlbjgGo27vw2qw
6cKp4xPDSC/Bt6d3FZWr4yYnIJ/AZE6vIPLLa3GeG9OvOnlFGU9iDmmpM1yc
+kG00KubEAvvqrh0GP5UWjL0sCCplNGmSBfcWQcOvy1sEHxZVFNF+wHr4Jkr
VPNa1/+rSGCP81p0hJ+h3LP+hUYUGvwp8ftpdfnwbadozb3992aKSyilVeTj
nH8FkwWB0mh+kfIav++1aiemDcEnZC5bqEeEb77iSwvxN4CKzOQoIEYe744P
4CfxfDZFCIq7JemO7XDmzlcS6E8HDFUucjTvnkEj2aWAPJt4ivWbqG40TOed
d/qUomx3wYCsancox4Csk4xZkMpE9lc4MGVBSkEPo0QqFRcyKjrVOK4Sfcfe
5E935IXBd83bKJ4OaUzh4BCCnuLLaFtCijafCgZZhgwPS1QdFAaHDjYc/ZVT
DOIf+ga4f2Y3VR/BN3LaLcD7kAk3rJFylNe73Z8pgtvFIKggQuT+3xIv0kcM
SgsrXGmk+HIoRzz4wuRLLYtY1eMBCIUnu17ZnZJQ2kZ+7s+HjzVT6xKJMVhu
OJIYhDZMvPpa1IOwTEdxbZp87tiQZIQJwrFPNo/RwP3xM9TSAee7hwiPOl8p
+hvdPKzkmHq7orEmJ9rtYxBoDVBECLM+hACJoFCmw4pZIGqbb9vgF946WVQV
qPdiLpmDjpwMRm1392yj4rvVnmFgWnVLCOAU5FmW0+56fZJqdyp+9tBGnear
LB8VhCY985mbwaDPTHhatHbly0JCJoSCLBOXwmZgFTuMerjW+UpxQF/p+ta4
PQOIvhCAq2sayEBwA77+OGImDbcWCHJQoXPjk28W5tFRhpjDoZsWugnQapka
7Gvt8Wzs4dkEyt4prCsf+Y3Cy5A0WPYuSvIZorObg1xg4C5icAneedyAlWZG
irPvlrwaPY+dxMk6cRu7vCa5Bjj12EzkWEStFKd/E2Uhs00n0LJ44r8YKe/a
O0Ndc5Fu1V6jhKIHqkL+hW1aN69N8LMJMhaJ3/lZPg+PBQbgb+D5Mey70q7y
N4LpNwLOKX4YRiuYrqad55TMfSTp2vOFXjsYwGm89aL+UOYrih+MlejdmA7+
7LbhzMZqu/KZeF5FYJWNq4/AExTMvTtJ35XaQ8FUB1XcrEpCqd6AKYvtNAUo
J1z58/HEP6MoToM6AukgY8pQJnXaUcslfI5qzaZQ5jpXQQV41IHi5TlR3OPY
cHPfFvHLk5Wj+BiNDpIJnX0aTqVA0b7MILL8lFu0lqi+9gPKkKbAWV1yPoG+
LNcNnbGRov+ht4ESW8iU0T8uhqdUJpm4uyytYV4fub6gahZzJEgf2seBDmni
VeZmIRO9166tVAnvlnP4M3V+CnemNAcH9QcvIEmBq/gGGyGjdtwwpOdb0p8r
zZ7DMma59z/UoH6yG0Dp4bAsk+tFWpkoL+d+gakvUD0FJ8LBFB3JJ+f8Z4RP
BbkChFXqQF2+6tuBcbfQYVqHzbF+NkfWTIdqvWJ1+tWmq85IIQu294xWxHXX
k9PhrgoAq8/6mSRvppG2ueozp06VgW6vnv181FNNL5EUuxyVCfw+fQpzMq8g
4+tmdMcbpNVvzopBivUtIlaM60oj4K+Y55w7Q4hScxKYf22lVoYroYA7Usp9
i2MyGX9p9W9Oi3TNJGTTxsKKE+p51cMNw3M6Nwq14lbweaFFAdr/LCXfLVPz
kKj/SGUYPuMh2Cd1KJF4EVbD+aN8at3kBiywPInrBkRuGf+XwpONuMg9ZtLn
YtJjVtmA0rAN3QfSNPcfq8ruRUjc+C7v1AEPwlPlPTbg3fNL8B8jJBJ1vICI
/5CpviAtNslomxPNJyuGzKj+eHtYB2TL7USyYryhMylysXRHf0JXVb7gw7Rt
Euf0Mtgt+D901R3fSRBEPUye5X6/t4vXKZC0lHVFtgXGHiimKO1Hwc93XdFF
GAqsDH9X4OPXeRam8YPPqQBAw1wMrl1zMv0/i15Wv26qJfJtaEtKZXmMHKcT
sVj4yqcIEAMFrg7G3BTHzun32QmSw/CLYy9s9rC0ISZfs5WcDK1nuOZBmUge
/ohHS2QbRmmBMQE97YTH0W4v3m9ptvXR3soIsW1PMl75Qq7untF1MU5ERJdc
zY/sEM1lwDx7j14a5N8cZ9RItw9cr72Bq9EwJtMGEmF/gB2AW0F5Y5leE38A
vT1RqtCFHNuW18Xn6ndWxzIIr7QyGJoRTrrGvIzoL+dsYOQrzLY87+OsZAb2
1dg9XueShkGEmoryCZ0j38DHlfFNZU0AIkfglRz7Bn3jJXQz+5/jiOEzNWIx
uwuX/ajwUiWeF1PdztDnNK1HMTIseTaP0sKCWvGDtGU96ayo8jCCZApDAEZG
xCM1cwFygCGEFoC1r1o0sxZIUiQgFFdP4xNwsWC1qTksASrd0rUr54/1LTJq
QTpQjfQJgPogCwIkARzsHVAHJdpB7hQnQfJ4gy28U8ohIUAx7q3+KkU2irG0
x1NBZT+S0OocKpBBFDlxj8svIkGXJ8sgXgmxvqpFYce7xt3eLV0ISk/koqmY
1kyvaaisVI1MJORdkRdGwO10Whcu+HkdPIC18CV40bNQf2VajtKMZf3p91j0
QLL7LsBTAFMvIp4GkdG7LEYPRvY149kGqyThA+ePSwb3mN8qpOUFhOuCJcDP
+A4B49QFGIAvXNaSoVFptnYgdj/h1ZEawu/AKY3CTSLGMPfvsqwxbyoeaxEI
liRm4C8m0AbzkrSsov5rqd7THz2t8Pqh2or90tiXoefJrLshsfU1/g1zVgqp
7xKT15Cvvgl6OnNK0KVHpm8YnqgsRqatbegDLSi29IpxibTiNbTRGca010DH
lLdiD8xIkcNjnuSgejO9sByW06Vg2zuhVVZe9sZ3Vt2BuM220E+T3UJYt2ds
MT87uMPXV8MhoCnR6atiy/WgGXEpTW5mmg4arULZb13tiXLXEKV/rjOKu993
iOVKytwp0koAQ3CbYfBwe/O+vM2IruluYtpwujmudxuGTcQ033m8OC3Bzefa
moz5Gr7jpvF2yVeymFBrnDF6lq+phiwASPLXhh63jT5HeimuYF/nusdqiI88
HTpjFMPBKtsrhg0LkExm6KPjJKAYVIVq2Id6YtDIQ7OIDLjddkMrzCAzBOh0
+6kfZwSaFirVGwVitojT/TbqqbmU1F5ON/eb2L+eU1rXhSiLJlIC5tBZT9Nu
xHrJdjznvIx0gaMsLWBfKk5aNyNez1HeX6pF0bulxKxQEqlV9kX+Cq1MQItq
b/l7XoxCUinRRr5+efa/UjmJSFYdy8RIMCRIxny58yJlXhj1nMWyLV/an0yv
lgWybwCRJzu5tMgWDl7sBJqt7sG8kBGOHxGyKln68OMNvs3bs7/gcVjG+kDz
4LEEY5EYZZ67NlqOJDVHDt51BZ349sKz+95+3CdWaRZESor47M94cm7XfDle
q0v5kKTQirQ8e2PoACmFZte4y0AKNefGbF8o2fladahcyyhoY+wDcnOM0i3V
clJ63gYnmWAj9YGhZRibpf3pcy+kTC7tGxS1KWTlrAYUsJR31S6eAl8IoeXc
2+Tan/MWYEUvGhcP0xl4RZXp0PDmSMmPqEVdPpBPBauyOSIB/zZDWbsfhCP4
vmeUZsSV8aO6bPG5sFzK8j8ZVg/3cr4ilZ4ZED9H0n5ymYXjcKNOK95TLbAh
8fz81rG1kLxPlhHgDZj0RGM7LZw/77V54goF72fsf8rfOQZPipELm1880OMf
TW9cNdbd3q2Y7oYNkWuQT+nzoy678aj1r0nE22z8z0K0YwrZbQNn4FSNoOCG
HEOczCOcvvaMALHHry6qPp3pO4ce+f8g/qhRQAVAqQ8xTv/v3fMBRcats0cU
r6B3YWlpVvmaH2J/BgDugIBtF5BLB50riB79Sp+ZFtco3uP8x+/EuF9TFvmv
b9Go+IyblfAF4V76AYLxX/Z2Bn07R5mdwfWo7C5WQEtIf5rpgd4Bj5/VB5A9
w8/eLLTOHtcpSR2ugnOvzPsnPNnW4RTF9Od7DYqRzr7x9VvyI24l5unA6iUn
yo4Nj2NzoAgBTgbL8hUKjESKAISUffGH4JalDIaZu8aosqhVAfvA6dvXqikL
Eq5yyHnUhBTNje2PoyCrznTiGFEfGUp/nBzwXL2FLSY7oq5i0qeVlLc0P901
xYlJ+Er+INNe/27WVcS5JqeUy6PcsruPRmOXqiX088NpbfoBOjW4znuTXxvR
bsNJX2dzRzenzP8JgiPAYr4l8BaMAd+NAkrfngBlmFGkJqC5EZoty80lw2P9
1Inb8X/uqVVfMsSVnlTySrBsrr6KPQ0+b2fNn1YMYTFUyyW4uxjtFVDKYfmQ
sqMETNVlzqHX0u8dO/SQj8rkBi251r4xHBKVFQIKvyVTq0Xha6JNraVV42Oe
qo1zvDtoAIy55FO6JJZQxO+uIMupylpAnUowut8tDbqLqO/Rma77nUElZQ13
5bBcZqhL0s1VlOPsIF4+Eblo+kp21yFiUwq2cA1ZMAArOeF2KwvOSwZ49CdB
T2Nx6GBwfs1AKgSjg03SJS43N9PKv4k9vOc5RHy/We7mwlweK4GMyLGM/Qpf
tzK/vJETxpaT3Vqqsn9xKFLqj2Yq8iUu/gk0daSayHn327JtQaR0+vTzxFCN
nfhkFkKT3aJ1mAyJHkWHEoi3SUdSxnegS2FLovkx8dShvghVhjxWJwwCQ13p
IwzlvpIhMhY6N5YpcENOBHs9Q8vDpvij52dXya7/Msf+oR8z1orU/LTHK1jS
f0wnnUfjToViChpcaZkWcxcF9bp7HwghsPYgimIzd3mE1JJDxTA2kpwvkHFS
4048JYgyuVEROdColMigHAfHYZMYXn1JHVZynyLp1o7kfIDYNCB0KKHfLC8x
KQ9ddATWMi/Rtuyd6rVBndyz3RaKKcnluj2B5dHR3YXmgsGL5yDfUncsFrt2
n1KwjagvJoFhLooN/odLjyIh+B/9flAvU5/+ZlePQ/x02Kah71Ob4TfX6Fwm
X1aINjBPLyuGdI7xXUyZWYuUBKrHUbU0U/3RLG75QUzn3+4JKedRb5+ZX+yq
22WKFwHPhl6pSUgg1sPH2EpULln9gFdgktPnqP77s3cvYfWGWJU39yqpAxfZ
ryjF2v1YieVcDmAOx/3V8e2M6xTmXHKBBktM8xneLWZbzFrDP7PWYSWkh8q/
9E7TaFVefdYi1mPfxfOW5t1Dl012UWphOLyxGk5t75QunWaE4camYz4I6PuX
FRBzkqwea2yq/pX089bs2to4cudETYM/oJserzP1TSnX0vzzZO1hqH7ouF1B
a9IKPhxSU7JVlEyhUKzh8fXuSAHszlBx04x0zE3VJT4kvFfSEvQZbE0dZIdv
7pz0qr75feum1RKQFagWVmIXqI8oejSDVjnRp6zHesRhuDdPC0j1dfcYYKED
U+gsBID/e0gP4rYQ8WtYKoP6DlgHZWZ3M8wKu7iXw4mkK8b8zSyxsAxhw46b
V2rOeD8ZwPNIApQrHN4MArp+Qzcwy+la1oqP5F++2VJgpBIBYplxGRnYaPJ7
YkiUqgur81OC71FbN3YHZFZTVFXD/UdbsVHWPnY6vBLSZ5OPoUPKDJcllilM
2mOQOWPuRc002OSy9T8Extj8S8iS5lcLtKuAUpRE5jgHWaoYiyFw72earVZ3
SfXsWvSi0/KmKqNKrV42aW1GlPe3/GjOViFjl0aQzxx2Ktq55s/rpaViyKHL
T9An9kPXHmjUGXPK9H70ppG+o3T2ZQRaM5Kk8kTHPMDrSTrXBisbajD7U3al
EwE6gQ+8IAcPWxLiV7P4Km6gbMIUEMO8AFktWSTouzt1B8JJT92sxjLUYV1w
QKfMlkVWhjJ3hcXH6jQFaIYac6AyL4KmowcJFnoMptHgXEVE0LZKGYMymTzP
AMlCD1FaQHzBZJ5WoPQ0fM/ky/81QgysM150j7VfVkWOuwjUg4Byizb8XbCV
uA12o+ri2ugxmal04TrK8lWaKr5gUNlI+O+y1biWe1MLzwTPFwCIB7E/9qjb
/Tcg12yNHPMCzXSwKUQ3J5UGxeWKwvG4U5m7y6GmJVGX93gwCDnDwXip6PYT
JG/hWcAnba2nBciliYG16qu4P+VQbrECQ1Z6QodR4N8ldPIAUSKVnjb5556K
vg4TwP+Sj4iki8qcXBibNTReub2MY9sC6Tkk6HKum3n1GyU+lc8438zH66/2
A807kBgXZnm7jgFx0IyZW9DBVlUoH637Z85Ap3u98Ws22gQ6GsX8xNFioQ0a
mHC2s/sHDDE/XUYFDG/QSrHKsXDO2B1fQOdaWqx0mIXLlXsMbyGf09DeG9QS
fOtoolvAowg3JJVZbVkDEVputDRxGOM4N6vJT00G4iVnoEYTpQRNHAhuNQ4G
ALjVHXfWSJWUz6iaL5S/oAwJ5QqeuCy5srrAZKVsOM6WqT8V9xXsQaQyinKF
mrJ0rNQjzqcK+x8jRoN7Hm7hWX7rs5volv3i17mCihWJ0WNVoR7dmkF9A3Dr
v3Gz753aXkoAugyINgVKZLg9vcriesf9pJmHjCGFDzWYJVbAUlCGMsZscw7m
IfoHehBiBk9rx41Koi4oiXwc4ZJ0u6CYM+b/4It1cLgJzumWJodkIaAaOztm
KnVVY9q0CrAAFbTL6ht1Z3qcdSH7+RgMh+1tKYkD2YPbW6+4cyGJxXVOFDrN
JCh3Qg+skZot874jDlDJPRSyS0SBK0T83YVWyMYkbsCxbTXGcfeNilZ71+t+
/ynLbdegbcklHfZG117p15eTBnN7+xOefwQRk1l6gew80RZdPXVX4vM+vj+6
CALb7a7FuAC+eUYGbkiUE+LmBMVtJvJm0CmUllNcS2soY9raOPU4127PTQDH
an5pFr1ju1+DCuBv2PFLDiOXSfS0YWhC3eAb5leJY6CyRHOzVz4W+3dGMuNE
Li02Cm9DpvCl9fwrZP7RnqmMVYt5ASIKGU6L+oV52imZrYao71e+okbqlvrg
jpItfKv9RorUExhvtQ5XZ8360P4Y3RDbjZQ/RgWuLxw1SXT5B2fqGHR60crx
bhUAnxFqHYjDrDPfvwDW+VGMOb7hDBXkoQm7qbu02Ruzu46e6DCzSFv3xaXs
5s5X/xrZ0CohkT+TL5vojljHcteEKMh+w7d7bed+lDif+OZHVXUXkuM88DTu
/TFSbRBcCJGpIWzWcWDN+x7X1vlbuLK+5XaQ0F5po6//bqS3bMdDubdgWRpg
fo9hHHPsUmbsn9TB/19lD+tUG8PaTHe7m7ezI1I6HbFWVKsSezw2lBMcR6Jl
QnhBvnt2ZBSM9GHEK8q37eAJtbc+0MVGBCFNGWHFICpn5QBlCerhn+5IM1Kp
GEzAfJwKSBsonw/IWELTYN2KYMm2xlvl60JhUNF6lzezPnvC9ovJv/NdaFwg
/C/gmQ+XCcATwAXs7NVzjt3XDJcbLihr9oN2yOL34GQIbJcus7Qyu7gtsz2j
auv1BAcZdCd0Qlcln8vAkKp/tn8Gm5RNcHzI/4JV81oM3pPWb+Crk/N2LPQl
2ZRCb2ulV7lfm0hX+my3/aj7wKwt0CyrTb3yDsy7DrMvmlWUSDN+1Wm5+AxA
/PM/qL4fX54qldxqX4kNhImer1EJu5ixoxYwxV9kzTFdWIW1lqKGRptLWkVW
rSGwDIay4fUqQ5/mx8rRji42XFNihu5whLetsIiLaSUI7VgtS4qo/S3HxVBi
HxQjmc0DLnQWj63lFQb4ev8WCGtkAIeHLVbqfmJ7wjbphyNddInCsCaoUaZE
22/eC+43Lvsd/SFP0aei3i64EZ+v540ye+KcAba3/gFreRuM/TylPzL7mb9N
SVnPy4O4WQJXdPuuPZwOsPVc3pXzjUERf0JtCQUWk3Zm1Fx+RGkd7R97WYSy
sf73nt+N7vLZt4NNtnVSDLIOBt/HP9BqRKA7f6H91+RrbGzE4d3/qC2V0WfR
S3dSWIXj3kIEBr5DgwDfKnArsdPwREPCuvwcKzuLVLV1KjNOqq1UWYYaio3b
QCihq43R462QFwoPsIWSzAbq3cArk2jGRV7R9vAOmByNI6TKQIFc4C7lnMQ8
/2MtuQXY5QbtCDbN1HsjwZnBcE2eNKFb4n78ZCXYnh1Yuvj7vsCxQfPDZjR9
026/7xtZl7LgF3UJzwcHxIdXSp4ZF4b9D+o8C04lnKeBoouF79gjLYEFjU/L
xJh4z9UrvYOseZV+VmIBRwxBZdeglZz907qMR6W16luM1v9+REbR2a6Nt7w1
XZ3A9olt4bUKW6vi19TAeG/K4+SLPt1FTW8kfaLIKq/12VTbCx471O3uL7Sf
uKHZjhC5lM39yP/f3/rQ5j0NjtB4+gyLF2a7bA4SStkp4ZnBuKQd6igySFJB
YyelRNE9qa2+uwjfQ1QJzhhH20wIuFrG9BaWrGm4wreXuZXhan38c9NCnr7J
XxAnwm01GpYA2MFtzonYOElFe0CZNX5usAvBuceCX0ETFVcTvELMl3CBR0Gz
HyrtZT/tIyuABmKPwmMaKo0KYHoO783pwBXoooBbURsAhKuVVAgHR2+Vu+4k
mCYTJIMinZM7M6gVhDr9OvzUW0AiZ/CR850ujAoJI0nr7w+HpMRuxd8Se3IB
8IINSPP0a/BGCcZ9EloFhAwLun0mBeAeT4bfHwHWxzbIuQphBula6icmrKuA
GjCO01hleIf6oDA4W2fbh81HsaBHS+KPgFFXFcl1jmPXch7tVdKkeF65DW/x
653P9emE7Q9ZfQAbHoVkrx0vP+4NRFkvBb6uqgqw+XB0xPU5WfYdQdvJjqE6
u5vSaK5y9mdV1a7xM3zKPY4jeXIIQp2gm8ANt4hHZpmD0UcvQcNCjEXJyBJ8
r/WBlzs3Of0z6cwy7SUtX+IT1xdPXNX/qTdHYs8XbVAQrJ0B3HYez41qMtFQ
NW/DLvAySL44EPycD9yGlV6g+FrQIlxQYaa6dgAWnVQcvRYqS4JZ2RRsCI+T
neuxJKn/U2UTOZF3qxjRhS5fj+Vb1n0QqrQab5XiGK84MluY/cDkBv/XNeXy
cZm/fIo1qIGfvxsoIcmBjpKSNDikIS/D+2cxtRvbKFUvXwSUHZAN/3zzQfPX
v7mqloEKssdYKv5EvHS8yW5MKKlZeFXwl/QNjOnqwHDvLPhIPK5LA67PynzJ
I5JWfUQi/P9zeH2ZRDtKWFILD0bDs/nI4wRLvkIhGOfAdI8CtCqGQrYfPWgu
pvkLLhIks7k5X3vNbW6ChiOyNdjDikBneTpo09AtUKTvMy2kuu40uac8CZBu
h3dN0seT0nlaDDpX59rBhnQl4q7gMyYYowqWnF9AssqjtMBnLq/7YHSshd62
E7AqeOVCU/yIBhNPcYRJ+z+6uxsJQWW+WMwZTfSFFSk12THmlhNYy7MP0nt7
Pakxm7TYmNYM0YyGEgyVnrNqiePhAuMzHnQGL3V8k9jBv+Tg9I4Y8GS6hcWl
N6Y/wm4dOqS+xT5VJl/1sDcrdTACbM4IMTlfvVDOuYO6/N4RY4ozmi7RzFAo
rcQjk/7IoWhcpK1PXXu3IA+OHbb/mN3r8DQs0MMc0HDBpu7HnFdY3ewukZ9Z
F0FAfeyAHZm1P0blTcexn0H5tEbkJobmYGVdGzUyCftHSACUtOB66mYP6wO+
HeqE/IzWMId+A6YaXAtptB9DfQBm+v1zoUyngEm6NI+kfLh7ZB/UQtLyvt6G
h4ZZWy+GdluljZ1lkqpTqHvFa245aht6rYKGfoYxp1eB6YAd6pB8g5wtMRB+
ZmM9GjL3Jzod3GYadVFoTCxM077nfmy8jIu0GPTWrLVNSlU7hIy0YlYghUaB
W2W/bz7yrjBRkwWpWQSGSaLwixzDMX/a0MNxE/pTt7+zk34kAR7utvKC7LbG
Kqffr9bgRuzEElkNtoareRZar13wWDHzaEvhlpMwIe9mukI6e2lKrE2IIC+M
RZWsl2cqvlcLMdqbwI6LbFtz56PAPptc0SLLWavnouB3OE+X6tbo34pxpSyd
N6VJ/57vLNo5D9/n5svjdZl6+lNuWZaiRSCQ62Uk4AUsqR1En4iEhMQvbErw
s8ytCVw0xepujEmLmPnwgmqGV+6Wxo18MNhJHZRiP8D2v72oBVAHmURQoaPt
DX2y1ikvYh2cGA56PMt7gpZu6nYt16KiY12CXBl/Q8Ty5Q9iLNIbm20aK7Po
6v9yRdytHVwKkXckygK8bRVbVWNdby5c3UPxRwm0FA3QFqiIQO8ANZguVDKD
sn/IOiBxIL1HKW3b95lcrX2lOKP9HIWGFsGXiA1C16lGIg2W0cooFx0aQFyZ
vgSYiR0CXAMMg8iOXKxfENvBzTwWgoyWhvNtkc52OKPhLamR7f96QaHxLQ8u
cU50F4xfwR0RE1zoUZeC6ODTLS+zymyZODUZdO9AFGxJMkrr8L0qJ5lvXaqz
lPFYS+7Xea4P6YkYihViIsnJMZwD5EVNO557Z+5cwR9gjmGPE/naLVKgMKNO
nOqqWb27KH258i2EZowrT2NHHJ6o4MUQY1I25LY1+KBKA5kSJfl98Iwt31mF
Rnck0BWYjfwUKzfBBcWwPXQcDsSy12gRtUn/xckVtLskUsXPDFKUiDGYSK7r
q2NbgaemGA71L49ZVgr1LBhYwu/f8tIFVuTuBIQKW5nrqppmK1UEggo9hvfp
NTlj9ZIvDdKyqFQp0l8JYrknFjhVaa9CD2sQ/2jD6rfefFZHWLyIu/JHUInv
pXMTxCbjPTiLnQ31Qmw7XImIhYIMDGrm/rJdY6I3D8mbpsASi8XI5XQ6rsoM
PAxQFoWBBlwVsP3vbyvOeEj0gwHVb8K93FOI2mzHJT1MSYiQTR+RvOjvv6p+
Ew1vvkQoZ7JZiP3krvBmLEnam3g9D3OQl4EJE7WgkTA4yRyOxvVP6kaU2qKi
yl1RCpeCUNUEjXbBJb/cLEMex862hkFdXBnAYYq4GxAYjIechnqw9nq8NJrM
yMIRMITI7dEgAAFlvcwxn+C01h7v4RmAZrCPyIoTXAuXSaGlEQo5X/ySrsJy
+ITmTfWvkjk92jr8mceNvtTzP85+5RyiELzkuVGp3TSDfOrisFR14XJHPO3/
UxX7XRAPlDUwUP/f5DvVK3czCbi4mTFahpVNa3KCJg5zH05p20F14SbzGVND
JZSgqA8J6x1MswPvWSslzowNWf1xhmPDNTXo7t8M1EVeQBykxhabt3PpKrP7
YQnKz431+lXJaVb6IL7vF2Aa0lWdmuI4bWPr9nhNv9VxiswQMBcXg1EsUEAr
iW+/KBmhPWeDh8HL0z46Z82Bs/TiN/Da3eAvysjfacbU0LNman1km2BoVVss
Ga9590RIrcSAEaIzLyVdzn3PJZ9ag45H9Nj4YAquBNy9FUsNmkl540SumE8W
gqS5v9zH+48WMNxx0ETVA3vr/KbfNR+pohJ+2iltfzp+Q5lsf/h89zOg6oIJ
3Yjf1Y688e05R3X/qIEtNrU1Z1z/WbVv9kGJy/IBXcAylK8yj4xDVWuG64hu
MSjFSKTpV1WzvmdAhA/+THjVJZ4bMGeAObUO1beVSLcAshJ181+6qFMYErC+
XPHf+0nR8IKKpq6HqVGxUK5i+qmzHl2wtiTZ95TrNECmnHAna/ObHi3HLB/4
D74vcr0dbCvCgUiQPYyHWMkNN1E40eWrEGLLflPna2D/7OyMFaQ+1mBvDBrd
4UAwKFYrOZJgca/S9DLfmR395ItEx5fWTt1rjsvD/YCn5K/iji4uuzvk+DpW
xf5Vr16sfT7XOy4SG3rwvZUhUM0akmVSHajxwzD8Slk5sJizcYh+MudJqUIv
OgyFVmuwva1cZ1JXyxwGo29L5SvWWsyNhV/rVFZ7N/c9naE/XL4wRu0pS58V
bDXi1KwjkS6mX5u5HAf55JRI+btLhni9vZpAHewjGn1Am6SirdHSt3WgDTUi
EaSr6aScaCoX2PmNUqSnZdrkTMgxCiWFMl9hDbDHnrmYZAZ/CAqz4E/ZrvaL
KqBJnrCuWjyZEaGLQLwHinxZjLC5ZHMfgLqCXehYTEOCM87VK79fBZ0iJBAl
X2rZ2un84vo2SKG9gQGF1idi7yGpLUOkOACXeD6yCajOhDWDN2otVIVVEYUP
np003GQwfEXfWcxlxX8BJtRIPm3qpMsESPQ8d7cqRxQcKnfDeQB55GaVeQlW
M7bhaOW40MFa8oHvrP/sP1EeDhUHF4uByi2d+lGproKnTkXeOA5tLzY8VFzr
pXxkKAB1iorpM8T9WY02sGQTHe3JO7On7xt3bFdL//Wv8mMy5MyjhINNUwIz
y7bjXwDCzBmFMSegyCsQUg+KxJd2baFbOgiohXAFMYn/VTUcAtDKd/FmNIJZ
RUak4Bnvmsx+62UC8e9MQ7wl/AmPDpv3A0119gSRbvWDXiz9jupv6OQpZ/3k
ncs+tek5Jt0mNruMYBccMDyif1rN350acbrZz8lJXA0Mm7LMHp5LcmPzng0+
u2QL4Ws/oT6NxhKa8awGV9O7h/QB/eH01W+m7RjKajq4kuLm1YPMEr9eS3zY
9BsRWsqpqHQ1DgCn3QgpJKbGfnaqAk+hE7ZaEWR9TLihdSs3bFZYN6fgCbYu
YgF8BmPhM1/sNmJsbLFE7ivpZ2mvxRRRZz/P+psD6sPFJfDU4zR1lCI0PHKh
L04Svkl1U2tuOTvuL7pNdeiNsqmRqm0ckGnKoLeo8RkYpafA8qylaiiJpKbV
PoBZRvA42EgCKe8niwrorfQKLVd81cst9GO3S5tZ5oDy8Z/KQD4p2GfWPRSW
gVZLFZOSeOBivw4ble52xMfTv8b8uSXhpVBKJJVIaXtfkQDPkNafTH19paMr
ZXZTUGFwQjIS64/AxgjNWIKaTbqpc1jqy2CB98jR9R+zsKpbOmdJzs3KuEQA
8J5Fm7/6n+JGWYXkCuX2WT0+bFXgSBB6r/viTgx3MAsttWyraJaV+XAznkbb
CClPKlW4opbyqLN+Zh49/f3EJMjhnxYByMOceY1szs3lL39RgrZUkiPfJ/G3
ico/0TjNGZG7/SnJmvC7S1vcf7FFyQ8viYpq297B0ANiMB5k1JTEtB30G2Ev
T8pwaiwsIL/fqXHyDfEpHzMBRheFlcQgJqxAKLoDiWBEx8QWp4P8oUwXws7t
Wq2NykxapALApdguQQgMHCG8x5CIrIOKdakLNRu1iaunxgm3F8gKU+hk94lG
/dln11ad9AwXR/yM7mkhcyBFKLb7Oxdpz6yv8B+Gx26AA26+A8drroFdQGSa
G+pZMd+JL4/XL7I8K3VbNFhz+e+/xaSdK2PCjbZdyxmdUw7NkVCK5ee3Iyk0
oBknD2sRBfLcs+mqNMN9JwhFkPnFc5wPSTNZva3D0bz+1Irv6xO7/w+HED+N
KT0zGRX01iyF4TslIbleDcte8GC2USjsdwcKOoC46TCYxqqzlGzPQ3HCZgod
TXQ8tzVTvJa640bK2v12aISVk9erShKgIvVY68z0XmSTmRnnshqh9L+uG2nA
E23Y9+Kpx0PdH13207bFzlY47EtF1gyh0bFDCLQrtGIyA604pzsT9jeriIRb
XrsQJU0yeXo5EpEfiPlcxZr6EfCu5eC0RkCtLF8hUg0+rsrQ0srr+JsZ4k/r
3sw0dVYXlfrQMc0tffBNOhn/3M8jmOub8ETZbUZbez7c6UR65sRValWPMHFh
dh1U4gvWZfQWo8nJnIMm2tkKzC+ezD8OuIEcqRFZQB2Iy9WrBZ6TiF9Z2cfE
EaWiqjIT8Q196LFgDbf6TuPCWz4v41FE2lHCbOL1k8M10hMK3nfpHjky00wH
CKf1cb36E1o4xCW1kUFUzsTNILXj0i01w9mV7WR2yg8Svch6bOfxNBx44pUr
5PqiGyYJ8oxezbni9l6oVP7nbf39NK+GI38fp9QOgAyAVAswY27g4zct6ysa
LljOa0r/TE4OBF2ZeK3sC3XRrmK+Zw78v3kDhrHadyqqEYDUeg1RSxZtfZEN
DmgwZQO2icX+EG4GrgMRcVL5mrngM+VQJRn5ME9mHLXRCYrHNvHmbXhFXpvN
13QmTx9nsO2XX/9bbTGHk9xxj5W1Tb8fcVZg9Dd+dzdrpyEzqoI6jvJ3fonH
pMM1RHOdOftsfDXrqxqwOpnijthagkz3GrxHHfYRH57y/fJG9MsGb1tylm24
F4MJlwobDra2vo0IPqWzE9cQoMsXqVQivMNFZenxkLlnzn90vyDKKqPIydYb
sXDNqH1bplJgn6JVkaBB3AgQHKA6k8hAX5CzqbkeTv+ov0+4DlBzeSrxOGaz
T9h86r+wCTVSwhXkeKA/mqPkVdGpL9PFkmzR53NeZW7mbCpcJkS6X4ngXrEN
sYicX4ysdl9dEmUla4tsTCWWr4AXNZsj3ClbPUfPNGD6R5NpdyFQMGDF2HHb
VE+W2ozW66Fc4156OGnHlItaco1/uevnomT96YGE4RcTUqWXGzglLTBdAXdQ
XQym7d/A6i+D0yJZsSO5sfRR9CzKufD1JV/VOiolC0XLva+Bi+LMKAxpIKp9
IpbNLWhisZo7zI1ylr0+y01+0G1jatGyqGRh6BSZnsmuSxRHEKpzs1QDnIHJ
JII9z10N3dRXi+wtNQYXLgKsY9/tqsnjB/NzQcBYsPSIoPUKQBmDxY8wUlPE
rDYzRZYS07OlVcHdOSXnrHjcDUk2JOgmhFCZtiEDtiGz7xsIm/jmA+CpOlFp
K82gJNJZyqj/VvxlPdT/cOTVkF46d+q+6jPs+FFzbaiKwmkgmACZginjWneV
Y1RhRNaJ3yg46tCTKnWlktxkr7YeLPvRNVqW3bu6xHJy0NT5rCHIWrMtLgcX
SypMHBdOi5BPmXo5zVXwTaUr/myqzUI2LjOEueqLmhxWpklBHjf1Tzrj/eXi
13OvPJmWf5+LSF/M+WCGkr6UHg9IEUXTqf2c+iS0rtMiJMLjUph+DNda5CCw
lpRulBWXr6x0vWpbucDijPFBD06tnJJhTuk5OsHNkpK1jmAR4WcLdKpBEJDf
xWAHOlHiUADbqetm8c29+ltZS/Uq2FoX13gW8k1pI4PT5H2PyCiqWfo7oeJA
FAaTrsgzaVH4gyjXhyOy8jIWjXnDdorQ398ay2RTjRlXQQr4DKVIIaLCS0f5
+oOEaOVKcu3ffuE2W/oKDW/HvuigYd5dTl40o/kc+t/pBSphORS4+jqgr3d7
I0bzNHer2bfgz/yxPIzcJwVYz+o14WQ1ZvfnxP46e0SqlhJSW41Cy1ZrFtVm
IKYNx2EPzwHRXLr8bfTnBHZs7gs7vdsKHF8hyNxYvX/Ij2rYhLSl5FASyQlU
8BWM16bydhX8JgdJKUkY4YPZnUt+H7QlpIfwyfO0rGP3oTmqFHj2rHFIN4zX
krLBO4osUj96RdU6UN9b0HoyvbZ6laosoueiQlVMi8H+ZGItW8W/vKyyUfYK
tzXjLSdlIziW1pM+hi3MT6Tnjg2U7D0SEPLYLHoznevDj63+43Y5xyaPb2l8
13L2r7SK5ak0GIB5LyJD9VDJ+OBzoyb0LnjSn6AUoMQE+Tkt7PY3DycYkZH6
t8L+lXIMjvG1Z0oDVTC8MkE7eJ3Q8osCyWuYRx3ZS3qlK6PBCLzw+vsydhv3
7uOCE/NUDLQYbrR17E0ChJVLOnhvgHGG2MrzA5LgHsR7ud8QlEKQ0FXjwYbd
m0tfmqKA4Ra6SrbgQZmeUYT890uUp3VH/HiI9clnLsdTjdkTRRVeRc6aPpfm
0tOdYxauAz2Lxx5vwMgPvYNlzaX27p4HEosYWiq0q/VZvjYvdlhs3VR7PlK5
GP8i/wOLI1XZpQQm9mxakgTIP4GeBLLgTxUUTOlAygIc02fB6wx69jVb5DFa
YtMvC0IxZ5QUkVyYfPfch5H1WKxlq3C914DhzDNoA62bJG5Hx6Tj09AWHtYV
6Lu8+lArgjZWdmL0JUFC+7AF7/+xBqYutIRe6SN7/zfflHAKK1awo5eAbtiq
aXWiy0sEGMGr6sKb1v/0O2wte4hdGjbn+L4LzAoLFDqO2eb0KP3qi+vO5F+j
rqL33P30ZKJ1L0y54l282hVsKfeadc+38fwwfrvBSheKjI2fURJSLOdqRFOI
0mzRAb+120s6Tw2pW5eFCOSrasxbUSAfFnEw8aAsr+oxBykCS0JFZ6dFDjcO
waHH97P0NCPGhOuTBF383IA4f+YUspXVhrHkLbG0PK2LHWoG6+YSsF3Khtf5
8invnEQEQ6yNp3Nyk5VxjQ5l9TG8oIuFc881pDdLIYgKLZIXXsW2PurU43f6
ku4gPe3hwVk8cA/aywW5Le6S8APIDFIkHzDn6wJ72cdK/17sv2OGoTFfz1dx
m4Xf5bJXQoOlWVi/lQTU/DuXx0G4BY4Qu7V8OIP8lpwR7KzV5cF5rkLe6p+q
NfLFJhNDMhZxME+hoAUXyMgpw3EDVlPANKJ6JahBbgVBt6NhIuNXvGxYzYeV
3B2MOSqkW00LYvhJK7oCv10CMP2PRftqLHpI6gMiLZZWjmcWyt0UGv4NSV3e
YMAYYjSgxIjMz3/GaDoYbEYwWyO3Tk5YbM6vriWb2YoBo2UfuE2ZDhrDZPX2
LDQx5QvrTzEYWjWv7On707pTo9QF/iguxzni09iW0BF8mfKGNEuTi2ryiyqi
Mw8k9Y/gNPNuZj+beMtxh95tJjZBZSw4g3u1bl9NKmENdhl8KfzduJJoloFq
99t69IL9tsP5t/rDrvx+u8mcNE7kKZenToA55OHFXSHJJqrk6hglA99iYuQF
eBvQhc5tIOwn5d82vGJR+QnBmZito1jw1GNe5nC8HevoNEwL6SH1QlrbTU31
zhBWo0q46y314p1SIT3xuDK+3Bbw0Csltu3JRkiqsNmO2Ir6G4vJGXYrrAFC
93KS7O2XRnTAxLCJVMVCaD/hDlwHal4mxVZRIVl46cNR5HEM9zPEo7LvzvM+
q0hwydSvnDjXJn9FCvUb/1Jo8hdrRUICh8rgFpPGo8h4MgSZi079lR0VzCsH
u4o8KcC/6A7bfzhaebseHrunVF/5/xNrD7gjNUIu4+aLVrWY5GU2hK5R9vKw
CM4JTPBw68cXOqRuybjtgNcs5WjpXyRJcSI0NRzLFflFcR0h45QQztKvNA59
oQUbOR7A0DiNaEFwgFFEWm1gB7wUNTSevM9jkoFLCrZ8/JhatA3g4nOnaEwu
gSVCalTshMztxEq+V3W+yeByRm3WxGxlIBooWgKKmPGjseYVNIy2YokCIOXP
FtV3k+Qp7ExxEgP99BH+vc385YxeACKMco+5OQ5iVtfwHLQQg3/25EQ9tZKP
5R+pQyINzlpZhdhciz5fCYDp9RAsx4iabp4mMUAbFWZq6czaF/zBBXY67HID
fkdbtLcMal+phs5WJsywE2JycVHcCRS84/A8Y894lZsnbKfmqOdtgTI8F17k
RhRlR79p6h2NBWOYwff7SUg44fwXO6M+Hg9Lys48vvyTJP1eud9Ak7qpkkGf
rVNxgm7Wrn6YrRhbzBLENQWWPd2G6OTAPqkurW4yi4N+2BYBKdXoT1CKbi2Z
ocy8w9ggAU0G6NkI52gBkWDxrT2JdwHAqAQT7b8MRrleyHR5TywCnB62ah2k
s1g3RYjQjTwP6m5gklLhgH/ms+MTZX2owdkUgR3r/oJGLWThQdxYKuGebWB0
o8DWhAI54QWh2FPF/IyIDOkCEtVFdUnHUWC4jCOvwqBfkgzU9O+YN/nqN/nQ
1eNMjmXYvp5USSeN+XklnoUzjXwZhmpnYJVW6CjIfBk88MvkXocbYGCD6uRl
G17cwDF81tE0MSIDux0R2Hms1sZUwquhOhHpzfQY129mBgCeMPXReVp0g2u5
ksQsXK2ycuF2EvP5/yphzeux2j94F7S6DD7o5jC7wIuLTNn2BY0CSHSmHiRc
SQZLaZtETzkh782uuYa33EWvor9Yi6A1mXnTCktq/ERX5OUSlwIu69p+2fvb
jl6hxZtBdjuhGBXZVbFL1sVsgLrYTV5uJC0RCnBfIPOdagqtBOafGJW/qUuS
yiG/qHV+aUkGKV+PGYdmjxGudkZgZ+thefT4Fee68NRjmWWwRR43sYR8L9zm
kQYOn3BcK8Ah/CU2eTvXIepW0I+UxhGcHQqGQUnRnJxbx2uNC91E5xxJo2BN
NuHWFZBs5hWFOsT0D5P8hAfP7/Gg+jSd6RxJdLAZwPSqEBM3lYyX8zD2EjIt
czly6uSu0uiStDk7W5oo+uganR4k43B/nVEUN80uhw22zEoRoBvS+JGwqdQs
bwja40FOo62aa5nZWnGYTIOR1F9l3yrj1BaFBNlMHGAZvOh5bvR5UiwVOtsV
POGSSqY25F67VfNOMfeeJ+eSDQ0j3eSMCpulQkllxw1DxA4+JSPLUVkAPWw9
8cMtiXO7qRCINpMEv5xjILJvx6vH4fB3+n2NQeKLOr9USlFa3JX2c98cHZvQ
rIJVP1HVDzvRllncxRWq3SWxtZrY+5zII6mZEzhnoN97ZRG3bcUqjiEx34m5
QrwMBU1pgz4DIeocf1Av9MHhuU3wQfLKSe3CP6/LvakepHO1Ey+48gmzJ8DZ
k1/AbiY6mxVGFcxKfccq074AIqEVLmBAn+ggoZNFrk64XjGVnxwPxwBjXHqh
NmmPuAdDXEn7TQMqL0H4bB/UgvfiHaXvbWDUDteh2yBSuGNSqcdfvdnBtVC/
LDB/CfYtSdv8a6G+pCFatvmhF1s/mVoyQGwSyyEQu0DN026C0tRHSH6ntIKt
cHUPXUhdobKFjcTQpCZdtG//Yvqo9vl6jnlafGfQjEouKfahhlsROYSrtNHK
RViHy+3bnaX5es4GgshvbbZ8ZATVwYAoXzDHuVmssnIvOZjke/Jtiq0WiaeY
pjA45g58Uwu0E07iKmVDrvWYERSogFNem0u6AAEsPOqSwLt5ik4oJZ0ogfTr
lh6+ZpSnhTDD+5qd1KwvaLjGd8MtR7NuScgF5g257b1ci5L4SwXMdlN2E4JO
vWEePmV/RBiGqtTv9EZnL070E1FsrSh8sim474XZLA2b8XZYmqf2OEjiEzdN
/xc7bvarLfO0hVo7JCmngDyATgR2kwcs7HpqdyVxYXprnhXIu+Fal1vVatHP
NMAytJlIwtch/jQAiJOoae8p5W8Iae3HdfXQoCGPJxW6WKgHpunS4ndqB3rG
nvDquOO/lMpxJpAT4K1yi4zhob83WHBXhc9V6e1cIf1+Ex7BJlMUs8phFBNk
K3k5DCSg7QkEfuhMGCyao01+fzRw6+m63rrmHefagx2z0n+rVQWn5+NGORpp
l6lrWEO7b8wRaT3zqE9WIyHTBBwyIjxDN83o0oSx+aFB2Gi5GOfNKFNo3VLn
mezPjEi3eiXktcBIzWLJLXW+/YLMtK2MEstVPAnaU72hwN8UFkTDDglyfGUO
hrXAkuY1zNCxcNip+On9RTAzdPYIlkFHtL3V84AwQVsSYLhFtfHSWdTJr9T/
mh0+nFfVKNa63WzmRmTXCZaVfHI9YNJmtrTCRL1eg3+FtkuLumTirAb+S7SF
YKOK9B1+QwhabdSKuNS1c4JiL7wcic1U1W6wChse5EUau05ufKy3sugIQQJ/
S8ZLBOpIMah5A4uUaDNXvv3nJ/kwbfuefzLDRAjzAqWWRtlAiPYTuf+EJIEe
YHQ1DFubbjHKWVUOgo2rS34j4Bzmx1fsoESmQYlHHyDf4XHWRpAAFAruJLE3
jQ/Hf0uQNvkwu8ilNBy9tlJk6utl9TUa/D48rqUj+/UOdFgg3bhot1mQYEJF
dixFF1O5T9VbhDV7/rdUm58DySLjbdUQVeysczlDANoJEK+rSYuftBPh4Tny
FXmPqOlNaIhrG+ZdKvqPFhAGFYpp2Geb3Zw9umFjA16zLNPawm/6cz3IGCkN
aXQ6zNIcMsG5xTISmjBsTYS9S5hni5NsoqnYYlwjGWtao4tUHrJX5T3h+zP9
xYC/dAviXTidzBZWpGuw3RO1JiJkqMdfvTQsxmdalLbBqzJlwotoV4X2IqTr
LogjwLPDH+ariDdh1FICga26/1/HMXUAUqCTsN4vgARS+jyOp5nJ+9LmObxP
KXTruVi/s074ZROpiI+K13NUqT2cnb+DUsAJ1cxzdl4xk5RfSxbrje5oiW/O
nSsjMxtvfDe0YYXngzufWFhuKngIbgYAMAQHhE7Wf+bJldOzgszxQfDFrMVr
HPrzOccDjcwh8e+MkUH/Uyf3NYBpkbkywtRuoFY1XJNXW7ycAGDGfW1hI4i+
hW+9Y8xPoDGajMPkqqbcaUSLMS7bQ7ERJP40ObHypXpIpXuqj4jQqbdUC2Kn
T5ntO1RiSiuuQrFXmBsXhmrIV2ZbWhD1fqrayRdS2vjhYNmoiqz1jU/su67a
q0yBySdsgP0p7A+A8ZYTPxRu6P4MWCD5LP6sMlTdcVOfijSdyHmmIXq3FO+j
g5YJLMuCJ2InbPwFImNR24gOXRAwdozh4CS4KPB0DxFTUpnZLn4Pg4/RYvCp
Um2nhdTuYxXXCINCV9o260B/+3ru0jmqbfgA/KbTFmg1/5l1eNlDaQo9apVf
gyTqUV+oI8jKsT6U/CxBmzk0RfeWH9mlNLoZW0iIPIkfoYPXcCyxDcMJvQit
DpTF7hY/0mkqwdaPiJp0N/2kqlCc8kxT93jM6G+altHlBaUClw+VhLNlrrlT
4l35iRiB7/mm7J3VT+kCczJco83WOLeDOdrwKFBeHsGG25ioH6uOyDowvQX1
U2Z58etF74ylQlb0qU2GJwaudFRCROw2ktdBkNoleAXFriLskOLIyjCauXP2
xeOoBEItVdUabCOTdGegM2568wr7vAlcwle6wEmTL8qbapIbUf7uTUKMZENk
/o+hCqtLkxJlYJOuOPP8zwGv2ugjJb6JgpjPuTRHdKZhP8rY6uWGHxR8u09S
O7f/wS9GgJbOYCSOKSzppVWPKSs2AUl0kai0oijMT3xjF7G6jXg7Q1t0/npv
6dv4IJpEqEe4qIbkkuQmwZi9pJ2umrDZ2BNwCVr9Hjb7xGc7CJYM2CSbjk2F
RCpXqEzmLFoQpQKq8x6NX/ZsGk50x8F5dPGdZmdl9ZDP/5fAiFY6dBNMo95k
zdKi58H75AVHPETl2VtBAHTrq3eKm9kb5gl9fqD/TH17JugD9JCJvVsJseTX
f81mR49jOgVFKJTKEXBAzBgGBh2CnX5voogo5U1yGIHdV11ofdnAsbg7e7pD
VWMb+Gc9ddWAU2zU4C+Q14sklOJOgsDWwYi0mI1rrkubrKGzcBq9ddW6qyv3
Y5AsMYG63Itf5iY8XXUiapb8YI5TGT5LnEn51PDSC/95sWAjpHNfXN6PnlEZ
6NeeEQIhoB8tq2IWo3C6hM2RGqGwOYI4h5Qm3Y/ywHipDZvwj9qRuw+5NOTA
MJ+3ffBaVXLj2LFMybrShRnfmFJy01jEKImU3gihGKq8ZRYgKFqqq0XQzYRF
YnOuF9ZYVo4omZxTKIHT4h6lrFc875RpQYk4u2zw2NA4XELT6zQOAVYgCz3z
0jYVNAFwzEi7zAX8btMtM/Sd0qc0dcMlj97hhFbvcj9WbJ5i14LdabCTXAPf
/MYUXzV91/Kh3+jq1aykZRPecZvI0LgKS2VvaG40NKFTRunpNYSIyYbfW6pW
0B7cTXeK03TQhFRplLdgrd6ZI8lYgVo0jDixigrrE420SMo/2RqihKyPs1IK
Jo5WkHTmiUKfldMkWlOjWNi8zJAwDcqey5F+PzmEiZlTwXjvkTovb7OqLOXT
HMsd0ImDv5i+bgH5jB1P0VnG6ulg/8FbCFxrGR8F+H6COEzykMVCCr0+7uQD
I5rDUlMKQocG+scs8ATFQYzldIOQB5No4gigrZP7ZjUVOeDw8PCM1TpS+Ix0
3lSbjRDTNtilGcMa5PYVyuA9Gn7Q86+UAiMPckFngOwuAGfHpsqYZZGiwPaP
EMCHsufpzPMdBPA3NXXkZgVbXJ2FgUJo4LDgUKzf7Tmk21l5c76rS6V7NsdI
TJnBbTY2JNUlip5uJjOTTpqHELh7I9sEEF+mTPPVnDxtE4dJ+yZE/As5Nn4J
c0InXmh23rovFp5+AxUPEJfvMuPkYGXVYZwFQ6Xf2xgS8mPskYhDLuO9GEFR
rEiUHOIkTt+K2wXm2sqAsaXgcuNc6oSioRd+xxeu1yclmIAKlR7iWU+nFy3D
TyzvXa4qG4/i4JOmycTKTYL9A3t5eilUzU+d0EQ3ANAQI/ZUaou+MAdf1iKk
Y7y6xrKw+/ggJcDOyQmzwcNoBej/IfIVK0dhQYghE+Ihuq2stqCzuoNMmr6f
iOgOJuKTBu4Tu8gioKCopu8GirU5UlGa/qFoBIsbGweAVYoacIQWu3GkiHGQ
hdOHx0Zw0bhcq3MW/2Yexb6GYhyXs+IPFEje/vl4bIzpzZLLB1FsOXD08vq0
npE2W0aFJ17wbte2yadX3O9WHWF/NBi4M8ezMmET0J3GXqc5gG7NR5s4e2MW
YL+MBUQH6QqLPcXn3On70qqKifAprr47uerWRhv6ufbSfGpaZUMSBn0NkqcY
SgRcPmjCdgu5bt8Zf2IEUNTh4ugWfSEnkeMnEVaOd3p7v14hiRNmxVA6jYba
KTPx7EYPD30n4ue/5IvhTZzGu7w1Em/YUSmOg3R1baRcVtQTprJqsJr2m9cd
7Ir1l/snCFq29ku9ayq+qC8OE2Jf5wjyqA7/d/l31ujT2JxHpnr2CH3cMWmy
YcW/ZUFe29V1OqLxrQx38z/GgJZzW2h9+ao98rvcK7ayxunt7Ne+Xb6gSCDw
cGDgDSQD/qRp0b4cmTIK8+/pEGIbzUj/x8M1INMP/z5FNwTKQ6n20606oREp
AKtJY5JFedpQuBJMjp7/rdKWsoSiJTM8Wm7jXhr4oKfvZWzIwp8BbRmNoOt6
Ps8gtiQMkVlqMkS/EVYR8NAwnSpQXVVPbKvpAVwh1Jnzmi6WrMefx4wb3TRc
mJo/LdVZF7OjdPH6MfIGSUUTbvD8AhgHPpHK2EB4s182viCibkl71QBSse0W
wKZaIHXNI3wO8Z1ozhiAbE+kT3sOJd7tOVkJhx/khWVsqotk4V4hhShhSo5O
lCfSRWfbywAYjz6WND00/HUJXyLNj9N67tbnK4w9YVnPvHjhYBwIQPRPcnyJ
moHqgpl6idhHt7cBYgleyAat7kxww2iP9R5IRKyWbqYE2O0+M9QD8Z1xM2Mk
9WbZnlLge2kQduW9ZLrNIvCJVM4UB1MKmw9DtyeLZNTre8d2axXOiZ4/KZxR
aQ4VSBXG7qA2rSJBghWa8l/wl1ioYTuERSlA7Ll/B36oPGY6NMf6Y4Rcsk/2
/JFD0b69CXDY7SDQmZIvpb5WaX/D1wTQhdjIjyYGBOTj0iM5l5DyBTcv7CXp
kbu4LgxB9uj0nEISM/M9d2kar5MiP8S1Qfbc4S1G8GNjlfIms8zfpdcnBEA5
GnqfC/JDKIf97qwrTf+Yt8BnBPkGdS3lcDNQoFldddwfsPEc+wDarANWiKnV
rxa6ZrwI6TnaxKXCJOf+pa2rGDNjnm4XTPBseYmRNzF1BBV9OpvCJEs5jZnr
lvQeVCBd8uDsNcwYr9LpgzZEN0tiUsCH2Pv6ME3v96Q2pqvS/sXSlImRrmmP
MrCAEG5a0Ecdtk+NKx752BhvqN8Wg52ngyQJMJDu9mD5/0J7DX15FuJNTnBh
f9vJBLQXae9HlMk1vl5+Wag1U1qg2wTdMc78cED4simQQVDUMpKEoRHN8kuL
DjhlbrePU9hGPpBxkaB8CCyvYWJBRdH/Bp461LK0ZIEZRMn5zd5VqxbvB3Xi
SNha6OC1i9/JLKaYzsXy6j/VExA76hK3jC4jh1K8BnsgxY23DmGZcMtjNqcq
ktm4LyVA/13STRHjjPwZt0WFes+oNPy/gmUKGwvraSdtGb/MDb5oUymTT84g
nNCn+IIab5ZmM9I37orpkNKYLiksRnC9ABQBhb5nDJsGkALDWoRBkH+ekZ1p
ZLW8a/On7WMmw8edsRRmW14tSQFnFukTWpW9w8oS9Li3PV7fNeJH25FH0b8Y
crR6eDQuKhdOAYzD0cK1ZlzpdcVqeaRORP+U6mKmc67wB98nnANzfN+e0ci0
k+cbY9mt6w0JtC2mxHE/SXu5yzB0aBxTzV0hLjLCPsckab3iB5lqvBOL51+i
73ElFMEtqtlu62te407AUuJkT0Kwi6UQt3GiKqyLwIaIyq3mdh7VsQbuMwje
67IqZGK3eYbB5TsIUtdjgn/UxBu4Q77c3rpa3yCwbrxEbshfFDF1Pv5wP/Zh
QHNrfdnk5A0MIM7wauYVNheoA1RKbUmvyK6TYXTbpWfYUEX3SMqGBEfO/hDz
GprOjdClrTfvJ46ftYM6JlLDJT7mIQ/KqAP4NFUAXEK+bUGhPHwfzNmThL+H
WLYnBUNwrIi2MukMQR0tX59b/I7nBP0/HAq3I25m3jTWYQ7YTwXFEhSRtjIw
14dvXaEq9o8QwXIWAYPf/eOzDsJNFOq6DkkRq41opgLrX9cb4jFdop2v7DFy
u9E2JsjURvBvo3xJkaS0+z/nBpISTVEpsOU16sYabZ8kbTnuCl1WN+TuTocc
gbgx3NrT45sn36j0Ga/s/27OIIZfrUZntivTCKGxuGpxWnmkvdOZRskaM7Xo
5OpbrMFDpYS3Fj+qY5EF7sW3RfNDihKUNSCN+cgxSwRlNzRCB5/C9Wo4ZG1R
C9Tr7Nw38x24210TlveiTYevybCBtadgJviogNiFDdpksDXCPrQctVFkfipY
gfxkUJ2c+6NvtCUxoPiJ5UTabppCuuTIN0X7PTutys0r6de9u2bNCcScYmcz
csZV/SmfsaLU5/nuEZCbN8kRyXrR8OHyFyLaqUfCNviDM3iirf2hlS7DErrU
ZO5smTuou3eLz2E8gAwHLuerE2yIK/oPV2jUL3Tfq0q+316vlK3Pzumn/Y0Q
cpNDjag8kIH1OTZM5xke5DHW6a1EL+dQjoQZ1rO4kocxkr46XZ6/pSfR/ECp
rBmnPB/GHhFIPxIiLcMxIzEPRKtKCB57WOD4EFi//iIL5kFyBxeCkxlSOlQ7
kJLssLM3vLOso26y6cX84ZK0ZYNj8qZrhJosgtacGPOOw64Pr3rpNTpI5qlR
SJV+l/e3/Comq5SZ+547WuTfD1M2jkuhvS+dCPkKmqAsAEc9c3gibarrepjr
Vmgt1gUNJ7xrpAVcRfuRKL30HC0FPLbrbTaux069i5GDWOaSKhBUQxz1wuJX
Zs9HO++bJi02TRhslsk/ErDUBpbyizZAdcHem7PQYY0NsbvnrQcDrf/Zzgbs
thVKozWkch5ulofw2kDp5RfJ/JhoXObe7SBUKDLUWWzm2b61Nk96BLPSr+/h
WPwdVsB/K2SxCFzNPOKug+de0Zh0zNYbNWDlrZD3ldK9wyeW11TUd1spe4Ic
YaHU3piLAjGmg4LSnPGnC+qvnY+AEhMpKUpu4pV9L1AHU09gJzy0PhPVpPTC
I5AAD7rrrTIYiLnN6cCuWQAr8CsurGCiaILLX7HmopFe1BDRqig49NIdUSWY
v4fXSvmVy9toAtuzTXSgGGx+XSnfgkebXKD1trNWlOukL+ctvlgc0X2guHgV
KQz6Uh7c4bRsZlepIVrnMe9pwYYpr3PttbznGa1e30/lchXbGwsEw5wPOw99
kk+Lovg8Iz6HSKAXcNV46qInS/E2H20kaYKh3cK517jnhTetmXQgfZebX6V1
RsbuEQa8aa7+KLsEi4Yb3wt7WiX8pqAWMouBq/IJCpF0ZEjE2gFIVUFyCX2c
iM1J/0E48qONSn1kNg4qk9kz1HZIGTbx59bm2owGM56Rl2JfXZ9bH8LV3Uxj
pkGJfJ5nKPrTYi/eCXyb5j/g8HkmhCZ0/VVO/ksTy74jBlWF5zpCBAiuN+TS
0KO4B7UyuiBrp/cNz9W0Q/FrlUOj6uFG2HQX81a+//P8cm+GzvpjZkCtOeJH
5f4PIFe7bOiIRO+6VlMUecIREEo6x6t0Cu+z5aZgL7zoXALpB+Xr7VemHwii
V0KrQS59OCA7vQ3H1ZKxVxzVg81Mo4RhVtnzWzUsIhgNjanMLq2NiC9Rp/Di
yi3v5EHPGg58oP1G5q5rS7cRqEmbRq3loxiGHVp7yTOMSImjKSCD2Xky7QAq
PMoEaoAEXO+djkmVdHAUQUloHS6PyIC0jxFUDngDsEdRa6tWTHzV+7ATWIAT
eEJ6iStVqOkHbKfg4Ky0+OHCwrhxw7oE457Z57ERPpFjsU6ImNiELJArwn26
9nJ07VWcKsZ2b8j/GcMfHtv56l5AGg281VR/PnHnmD7SG1dtrnO92kqrY+Wz
GQ5LlwKspW0DSv2DckgRl/sLABaggIuSCMZtgpqCeE4r0febDOQHisl2MyHb
cIpeWeYSYaywJeMe3VHn0yYB5EwYkxyc6mQoV4fztjZvdATvnMxklowxtZt7
IKC3xXSiV00lIQRvnjruQJ35IiVxFWXWkREG4oE33afvMXHjGjzIpjsLL6Zk
t5lKEEuOtq/yF8C+IfY4K1LqjhHE1/zeJeU1JAVjtcO30l3a9yVu2P/1vl6g
LMBxzmgR8ThGUv2WuVyJaBTwhJpF2t/jEc6lj9onAYEFumH9FPjdtm/spbWS
wpXYxTYGcr+yYrzDJnjbUKiwwUpVSyg09tlYz/shtBI2NDKHSGhzrYMMoKny
qVoJ5QYMI/yoMLCtRlG+M5lUoPrYlgXcQPcN1GFtu4+n8sYxht8NoZJSho9x
IGSoj9UsvZLUTv3ILRWgKHiSeyamHHI5/PbIwk1m1X0qOPT0nmoTVqpsO+UG
b0d/I0krde16sgRG4iVITS1+Ds3ug3eHD3lqL0rnyj5VRpm2UQYQSCYtgY8l
C6S1lEI1lGzx5J7jjkTGaEDCoGeN2s2NL8PhZvTS4OegG0a+OI6W/NKQi2cg
xEWd/RK5qutn6RYDL+teORT4/pe9JFm3GwbiaBpcDNyeNwjlhZAvwnwP1vq3
JVhUQpTHFteln7S8UePJFcpLOPX2e4C6bOdcuAXvM92j8Ofu88aowBt+VGGU
jWuJ8FhBeLbsawA4kbVsyK/fD6GgLbXV/q3E5rU4CIFvXLY8eZ7BLSf2zELy
HACLzDQKYr2EcbHO+zzO4FL9wiMQYEjSPt/Azo1LiF7ohYfqRhSydnHy8cNv
BSxKkGv7jNHmoB78f8QS4WTmvCitwBB2qsC3QZQhUM9/14mBlzw5KZUmshJ0
z0BDGamyOiFsCrzdS1wtfiO157z0wI3KgwSNb2/uMMe0G7+EXYGTIo/RwXPK
UhsekQHH19bSUV+u5/OibuYW9zA6ipr+is6uUD41ZTSJqkEruWuLZPjWoKHO
31LcXghOxiKtgPbyGbt2ieIY5L48QbsdXwj1aVykU5lV9AXaHRYRYLXHh3LI
n2BLccBJ+sEqbEJXguqf8MuuV5kw2ZIRDUTEzDyK/07ltmhbcKf3Oh7u3Nze
ftdxd/dToAnMgaJ6Xsl8ShVi339w5KC4C70QfnID07YyD91wgc4/ytOr43AC
XaJ5QT2tMCOfZGfieL8s9kzOvn6qAkWK7zrFayGSsKTBhJIDys6aGXdS57hq
xKxc3CFgXGdpqPQx9tVh9ahLLgt62oZHOdOswV8xIu8n4+OVbayRb/MjbaR8
mr5hu+ys/iRLejfA4+LJMtTcraRU5FCTXXtKSEbzXk+LY7GOKYbOlO68ZVx+
MvlNby7SsX4S0BwwltRYmdBZ+Guws66aPWcz5nSTHIoHKFH3wDlgeq3BY+mj
a6/oxw8sdpZc3JwQHHM8iaQ60+ArM7XVEHsG2vsjP9hkNghK/IX02WefexZ4
YdJLq0J+ZzFBROJg7lrTDbdWrrRdeflyE3qP8KHitLkw6ok1qWcFcPT0+PIb
ut+IjJgHHFV3nU4cqFURkL4slL9oCio+IthaIIa+J7L3sG0rSg84W8RCB6xL
K6dEI+5utpUHlMxcQ3ifnCoZYKCUPupIuKLGeF28umJAtCEUWoZ91uH4s2R8
ZuHkvZpVgBgD38zf/6rXT4o0VbLmAuKSIQtL5GjQUL7fSEmQz38TOZn0N//H
/j+Pkmnvcs7TwgHs2A97S++kke86cvMKnpeI++oxqBJ7xcbTUikmjiD828Gd
htTy0TmyuRAvHGoUfHuXFzmCWH20ZTRQ9Vgo/XHqt1l4kiXnqgbLgrcNH7Gy
JIcW1jaQ/ege3f784q1c23zGHAkj4DFBBzKSe85+/VGXTocx0mymIu6Ku4ZQ
DYqeFu+pBRHfrnrybNGF2gu9d52lWEJb6gkkOXwr7ZjE7zErncdjCD7jqIOz
FFme/iMEcxuIeOYLkgjNzgLzewXyP43y/CQex6d8VKWo9qcergPjpx0QeXmV
gcL6DV+qJUtr6ulv7Nd6MlDNh5Z73WJzA+9aB2GnIFujEHAIqlLRRRwSBd+X
Bn4y8r0VW+3/8DBajazlARqBKw0gPkfw8VorInim/sRIfuxIzILdElgNJYkb
lGDoM8TXU3IBI5TPRQScOZ26WnN2G00DUkSwW+hA6lq8RNrQHMeQnQFfC+Ui
T6BKdpd7z936cxuJukDs1ae4S6ity+Dmys1czbZxm7NFThtrzUApJ3WZGbRJ
LflXxRYTTAAi7l97/h3baRwy6X5s3d1H1X3C3mwKEl9ES3FYNxQvJc6tW1Jb
PFrWZl835+Do9c4TKvDxjDCNaqzrmZjIZddyFxAdAdwz5hQVPb5le2dfdxOF
vqBQhSMhiY6ryn36V+WAp6yVyA4bPhF7SZLGV06nhDQIwYX3fIrON8AiQ4Pj
Psnxh/+zIv69Ach4k3lra2vSEVGVOUV/OhJ6BPQ4dBp4/mdBQyjl8u/Zkd2M
A8gmNTFgSmO095q5k8G4+rpb/mTRSjjr8ZUgN7IlvzufAPaj4xohXDyOIEzh
soQOhNPSxoHJf0RbPrIhwxrYISWr4WtOY381sFRCcIIyXqEIewSo5kLL5hoy
CZ5JqdscmO5IPdbsurIw4nBW+VSNZtIUY8m1RK77pWstxGpiG9w6PH++rvh0
j/xwMshor5kRLwcVPlaKQC253A1HmHc2MyuAdITdQhk161yWKAY66Q+OdPKs
kw0xfl/ufEED/vUzC3CT+kqFQ2kcBSvaY2oOFs8KzhhY10i3tTo4rkvB8IjR
o3joBQOHTUbubwLLY2J5C+tRFssaTIkc5t+CLfdsBsA+Dan2VJ7SAqBhVfWb
53r5KtCrCJi8mCKFlXVAqMpX7yQMsf9Bg3kwwxGgWm9zZsnqEYPdY1h7rgzm
Pw8ydGn289tP36uZ2KmLRHMOZW/i6escOAxS44bioX5eBZZlmSBq4PzxHiw4
CeJZo4s8Kmo3+ZQC4EMStkOvoBZkemtA7Z5Y4D1bvFUEsqb9CrVZjxU0oSLO
BjjDguYJffcZvuh/qOmEqs0A/FdnU8u9baOZ+jS0xs995YlRxI9DMOdUkfGx
d+evzCoHxgJhOhXpdWw98PHUGfDgXAtB/Cod5cZV8WOaslfH0/kOzgF29fdR
teRytUVDUQW42L8NCPo30ia7dsnO5abFVRPWZtw3iZdQvmx062r8XKgmDioW
rL6RGDe9PDpcbU9spDK5oaeu46oCUrxa7Xm8IVV/9QAYUF36eb9f4931LUfi
AFWDO7vxXQmGJe8Zb7YOh0rfTWv181BVV2yfVagU5IGQWNeR0Mw8rEN3e/4P
3xq3jJBAateKzjcRtI7ROTezjUxH2CxrKDrKPwFKcaaRaeehxbfc7jfE1MGf
djgRuHyyHkjcmeoS8hmgvauJXuAXhPk3pF+DwjlQC25s+G2jR6fw0XD8pb6E
XXPm5QQwy9PBeZzJCqEOFS1epWBqJpuBFH9eTLXDiuOW6r32IA03FJ7kYmJs
q9GM2gxCLflMElrCioN+hhVY6DgLreg1NCV7oNPfrXcizDtpF6nJPKJg8rEU
JZr5AA8WfuKBp4kzHSwK3OB737FFa6mD5NRU2racx2svBksIl2H4TfHO4jeQ
SU/R6Irlsm/5cim2Q01b8J0V7q+/NuArb1uYC1Kj6mUCN6LQ+QxnEr5fOf+f
fbYkTG6kodDB61BTzIBEy7gjilOAjbHe+FWTZ6JxMsFHbispnz0zQLehWcWC
kqW/dwCUYTbtGFpJzv7tqjF2UY5UU+pvS2CprxY+F2HwI09n4mAAcNsHDvqi
FHxdgyHr6qw1S8TaYCNhjSyah70xTBfUgSifXORsFixE4QJzEf/NaFguFMjG
Mbwv0Iik2r+lT+AdDyPgcqoaFqn3vcEc9YgsuMT/u2ZfwrpLuUkKc9fKt0dl
ZQu0jflOiRLX+V02CF1/YM5NpYsgS6JXQvTUJKYJmpTE4aIIxVdf+akISKRW
H31KxxjAky0zQViKUPbZEyS67ZYNEvwYrZzpvEoMCoFnAWXNT16xIvU/tnn5
Wrb68CIZdAnaO+NtZFOtOs4pxPmrvf0BokRxVCyt5Qb902D5NyPGODg+akXQ
zTH7k/E3gg+vHxGTuvz0hNBx+zGd5lmm6OknQULs2Mi1/pJYlvfP6+h+f6zT
l5rPOxT0OPapLwHWVm17OBtyKzKHFb0OxIpJlCD4YZJQpcURBQPiuHhOmqDb
EfqBuHKjUOVJHD/osmG5ujGB3W/twvsAPaS4/ivA6uZQOLbhsxX52FQ+lSyp
nrCfB4MP54hZAgaQA4PSbJ68tYJMtL+7/sShAi3MAYDz1ReACnBxDpoGw/Cp
oRIGMOVMN37DLyoYyqi1rPIF2hRO+E7tPKUFmAVIOzW+aBNwo+w3C1ZAGj8X
OdBlg7Tvn4P4jXa/iZJo6KgQb/prDhBWoj95ximoqG1UckrxcaSO3EjqUczO
1PSY2aPzXgtbo8pWClOFdDCr7vRIDCpA5XR9xlrxD9VCYCuM7/dEVIZRUMyr
E11Q0Y6NS1MRQ6mdZPqItGSDZ+6gH2GoVe0GdxdqlpLBlvuY+5VoZeAu47ZP
MbnVMFPRjtM1oEdCipT2iygGc7Mpcj90dKY2xIPtA4rJtNZOGF+8bLWJfsPo
86zDdAhyU1/ScBok4VrrofBxv4O/ldet7PORRSAFZFkCIwYvzXJquo5SAswv
W2O2BlNeGt/ql5dKuLyiPI/iLlZ/w2NV+XgN9yVFnjJfCNMze6CA3XLWhOBU
FXsf8fye7blMX88JR0eYWGSg251lQOhllNoxYHldmyPXzWQc9ef498XYy0IG
t19Usur6EtMlrBVs+XKav82qSqL0HYvgcNOpbv0sx6L6/Cjlv2xYv5RUJtDJ
OfMzFvYG+SPYE+lWSQyg438z6PJJkr4F1V5FLYzywdSXdCd6Yv7w0KMewNAx
rcw4lffP+huB836UaT/wEORjdruIMJZyX2mT9gfx8V1AIrIO/wJQdHsKvlOu
bojAQQD9E3WrT6pSAYwpmjC9OKBlPDOtDibHGZtQKGlX7bp6x/YFbQLPUd/e
2RqTKQwW2ozCYFoG0SpPr9IbwD3D+am4s3GWPLxYrr23TZUrJNnz6umTH2me
VitkpU074EaNLHYzH8XOBHLUD3hN/B5Y3fRDQJL5K2E7ShZJLai0FWTH4VCT
eSBfdVhoVZ1+oZM08R3bAcZcZiYiC0h2Q8H14kbnT1WAsD7j6iAwBdUGMqRW
hFqsIIhgB0+uCPN3rdpSKpgc3AVzywsZlgDUqm6JbDPJXj9bUJgvQVJPl89h
NBtv4I6prKQWo3Gz4vzcooGt2wdQrhH0SxvcFkYg0jZho6eni05mPgW0Exde
kvYTwbPou+gBqzRXAeJY+SwoyLOpEW5HfZUBqmhOjDmJGmHqwGaF67sZFjRz
orJQobFAf6cC9lhlCxXgDgqw739ndPCt6Z9dty4uhnG2JFvvnwXTalPuYe4A
nTwNiTDaPJkEQkquK+8cfv4QnL6erOGu5/9bAGt7x8tGyC+6CHwDj18undZK
RPr9u9OpCZh/UrC0Cv+OF5JZ08MVig2q12V7WIvytlD0/4KdHQs/ugQAZMfJ
CC+YmfKaTZb/IAZC8IdiLlQemt3RVcpRDcbM6MFxUKAKW8ss5rAn4YmWqGSG
VeSgoB46QDYPfd2xDaAvjJAwsaubdayyZywwd5noIBcKsMP0jzXrhRgIe/Sl
yXkwsTuIU7xtJJn2gMG1ZPCRzjJkdhd7NO5kRZcmbXug+Au9UtQGbzaTr5DI
cFEWkO3tJJbOQ+E7BOzsvGEOm26EbGA2T8w4Rao8rIJEyLi+fxf74nqsKo6x
i+HCGAS0B2AtV/qZJ8ghQiWEh5quqb0WOlwPkXTvBmznPFWQYbgTGwLGqvwq
5hRhd0qbtuSVXNyWzXIxuHkYc1RrDL8lkpNXLMOi+emzOSn3SmkMCOGIyxjP
YQQqXuE3GLlOhbGOuvmyAn+sBcQ8+dqbxS0delw3GdaSa/nDNJdFBJKpxaBX
bv3TYmpBni+2eSzv1/fgEL94z4IkG7xoAtWeBaJEN/VqC/AkIv56gh3oIEf7
PrjoCEEQtjP2kfdEvsjRgwQ5FwaPLKEwwSBwgCZoiiem3UCK3TBOQkKxWX5h
36Nlv86xGum6+15ofvKS0JPihGay1WtA63B7v03yI58zezpcUqXNSk2k/E1H
UAg9nGyUZT+uLGQNyB1TXV5EHjzut9pRjRgs6nU2UAyeW1vnaZT7C4XhRzSb
TmrxSxySjOv4/u+gGr6mmq/E4RmonvSM+cJgChcVHHhWTozEBnu9Z8LTOOvB
7XNsrxnPI17EJGvgk2B1icEBO4P5jyUVFNeOXbYZu3Y/DnBgQorhns2lJRRu
l0WHGC6/d+effuUhxFIvpMG+QTXVHDL2LONbzwPcdY8LfZJKQT8fRg0xb+UT
uAfy4Wr7wwyctnqyE9sgitkMFrLAaaR/ELn4IS17gvWDAFJjsEEcHzA72zCf
ILuQjqbYw660TzWbn59UinDDlXcbP71omFoN1t+3BLQxZ1vy7TRM84XY9zk/
6AqTQMklPtC1+kCErwQWlW/hDPWbtIYurMcU5zInKi0fMfLWX8N/BLDggoMo
p5oDMS3h0oKmieYg+8nB7nxXY5nGFWbYVue2og4Ce0euwKCw4/BLm4muleou
qzaQo6lsKmAs4naQFg3Sp7aXnjV2yvrPB6q8BlmMzPt9GdbT1JXyfiA8Gk39
P5PzC9bcILMITrOv7iMyy1jPhpvzyHH2sVy2mAIGnxEa+wqD/QFZt+W8EafK
mUBjT+R6zhEZLupPLCkNJpKCvMS60n/XJdbJNyllgM6jRzVKb7gmhVZG0zoq
lVaY5qsTSfCbB7cw5zYr073kgepdp0gzZgg67aBMRRExzlwtiagdqCilACy5
QFZZ2NVZGIRDjoEjbvEtOm3GCcax09W/jGfy55I9JzffwzilnNz2H/nv7omM
ikqq5e+bAhoLcSICWMCF8dPKO4hvfCP2f6vfOOmSAMXCojrWdMpYUzCDmmzJ
XpqDXWghdwy3cyc18Yn9zwkpq4ysRt1K/pLywT5lcz1sJSIsAzE3hA/8QjXl
Zzm6Lf8xm+1Ul+gUNsi73+VyaumBAuwKL6UkaCheU3sEDxfKxm7yZ2xCV9tc
T10GW7dvIsKKOfA6Hu43GGA+yGVmRv2xouD2uwb8+DAwpN7SHVeevgbPkf0g
voaXrbnS95fVxmMDZq646oE0nul9m+qfC2Czd4HjMLyBmH+Ti1GY+UKaiUrF
cMHX38n+BV0BECunrRFywQ7sRh6f/5I/xsrCYAtqhItE0c2Fb/EKqd6RR7xq
eoTr96vngNtsUbOq/1e9RlLu4Jzc/FfOKnvwi6JTHWIYjRv595w2Iv9Ij4mW
Dmiga9FEvXgueK1B3Y175o49XR/YhpeRVrwHHepO97Tg8AHlHRqTTTXuKmcg
ssOzhMRibVv77OEak47lYqZOWCFxOzLCQEXUWkH69Aio4PO+iRO2XmllRYIi
SagNJ1KSYuTAv443rVrN9+gv1GSWp8GR7vk55/dDfKsLbvYK+Kr5XgJKPbya
ZKMPPsGdWeraJJAvgWLmXybD4scsW09/JlsNsjK2sWaoBXMPK6aZHXZ9eYg7
7jj0SkODgQsLjLGnpTlcil8LRKvUJBKw2alatogVtDClT3wnVtYkVGy+xaCa
SzaTYN4msfKeyOkvFWKl03YrecFPIqiafMRBoTHpPlZq/gcCoxH93RYrQRwm
h5kSeJ0J4hGpzPgDpcqlDoBji+uZimn7gLMJWwNb3LgbzmBHpURQnbS9InSU
WaCig4kNAbUvV5S/izLlnjAcVK9tAOyNW6H8zboGEdg5UbjFkFrkGLKMacIK
qwlfm/kdl2V4MNVAeu8Car/7Wa2ABLB6r80vYHasSFz+5e4l0TSrpMkUUra7
kbW5MiLqxTViexIOXZg2N4LMm0Pt1EgssY5d1xftsKLRHj+4lx/FUrl9h6Oc
VCcw4MEuKLA/+ejeQyRN9JZT8fxV/Fi4PQ99j3tF5EuE3IUA2NJiiITiqt5r
pdenuCD7gdp8Hw17TDUR9ZegKq620knkcSqiCwmU4tthb8tSxk6OVgbZy66X
buQF1v7/kcNE5uMFdKUqPXdNn0QpdVqNzSmFuDoTDxSlUfk4o77z7bXZ/JGZ
J9fRv4t3SRLAEjCXtO2sEN5LEFrkDZk8ghZoMFU1lI+hnjQO/RsVmaHWt/WQ
Orr/SuNlGOzKSG/BEsH35EE9ZcJuD3yoMxXH6bVVmJDXyN/zPDeINpEHHLGS
1+p9At9ezhhNmNl2tIEtJt8tR+0u1a1isxogApKODtTkjZRhGEjZMl3/ywpD
mA+Q+Izh8xdnszptdoaNJ83wAnQ5bfTg37cxh6lCueaiQ6L/FzlaxZTjpmj6
kkVnafS/j8EqlaA9sYoNm5mKK+zpXTz0iNSX9ZlXl9KnNoQv8k8BzcsZPmTR
p8rWmJNoRylt2JmPUyJoY+Ac+0jjUwfswHrEMDDMAs+0lrCJbyFnRcLfDTtv
60xAfxj+f4qIlb4Gxwbi6a3Ab1w16pyK/9ZB/PTNMkUy+cP7HEDs6vq/zjnI
BYY2b6PNxsBmA9mWUebrirAu+5YKT3w3BXhgXoj3uepQV0IbHpy5fd9EBNDD
BPFObsN24wdzTx5lGQpzlAna4/7dE8Ru09+x1wSpiwr/IlEQ88Nwx9bodw46
1w15MrYkOHCDXssayC0y2MwwLqfgwMUtEs5iT5lzu3iSb3/NgmX7SW+4QmG7
w1h09fad9uS6FKHG8XHd7G6kyEjGToCUtG7e7D9vzfkdyTvWOfDHmATJZBaR
5mpoa3YbltpZmYAxBXAp1XZztQyeqi6Iv/uIye6gWVAr2KI1y1+JTbLJH7bR
g4uaxIh9PUOAMDlHHu6VlDty05eBsj2EZo2qT9QP9cH2a0bQ6f2m/M1c/8HN
HSD2W2JmlMRLechdr1hZYDZvyjHFtf1EEP//Nh4AS4JFmOCiEKLC0QChhH8t
zU3f+5Un6nQLUlp2BwZI+BiNCK5+pAFZkFJPKI8wu1RiIQLXkHG31rvHmB/x
Fx0RQZ+BosJQCD1hJMArunyrvsEee+mebIYLIwoSjCVmyVkEmREWgLf5senD
01IIydByxHywUpOThzSZmkK2WZtjJbl7qZ25EBXgSZC8PEqpTeEyzqowxA6A
23x43lLIdxES+dYVQ6mdjoknp6VffzvntLA+I0YgEBHXzPhMLaT3R97qb1jh
lFmYfTaeZ2rNRbb9hd2Y47HNAIyWSuxcB0yCAorWtCQr1T7fD/KJgMeyw4np
dc4c8F+inbpRlQIWNg6FMrKEoOpUz7ybISJUj0I3t8kSASmoZhF1AIS7zcO7
3BrzTiTZviTBHhXuTttBBo85DfQySS7GLDZx2dW5iDRI3yZDarYx86Jq41EQ
rDr+uctBeUw/bii4OW4XsYHjrGqCEKReFHoB6T61iY7ZGOM00DzlCSwPvc5Z
DncbHaeIrPHGRxt1cjnr1LXR6qJIXFYn6klhWCOLxnWXKLtsO9UHJWQ0PZ5q
5doZbq4G13ad7mtuHY1vlEsutXbFFiDRVGVi+XteJvL2Rxdp/v1uaAJnaflV
lEK8oWXJc1rcnz8XxCcdobW/DuIHVxABq7XMr8mnCduS6Og/pZWQczGJH2/+
dR2B4EZRMqpnwOpdl9o9vt0fMER7Obs6erX5liVIGDWAgNwtYlBFwVL62gTz
YEWDhuIuTs8qs/YVS4a4n4LgNwxyW2hAVLZ527zhB66MLWzLKToYvzTlA9N7
Cq5fGrIrAKL+6hPe7Bt8fvV5bC56OKMkUq3c6JNqcqTqrI2+4D6rKmtfNYqU
TTBcIplFB8sGp1PFC9n7UNnwOCelSfrqwrB8hY/cnqPINxQyix9Z4gm6Hemb
YdzNMC+ZN4VWBscRYwdznAQLXhjIqEnrX2PxVQU1gc6JVN08ukcKXKR8zgoe
TH5uxCqVf/HU+qI9KtUfDpisxfVV+ubWuv63ZC4ZQfBeZANESs7O8/YfNfkQ
csdoHPf91tQbzggZ+wH+Ix4a352No0RmQXDvTOY1XwEw4PvHga87vZYNHQuB
YAJvYQZhZqWoKjA3vB5lBg47vbLpJWpjCCVBHYTP+3jrM4Pu4d6JDp83eKPc
yJidBbgrzjmdeJCpKZLJ3UMxydbnGPKBTfJmnwbA6e3OuHvKEoA+LIhf5X5S
hA/KKO7/mlKeHUBGqvQXCbbREjPBxvslKWCBF5YxBsk4+Dcp6xbPU4FuJQ9w
iyVuKiyq/SJbQ+fM3zHI6Que2zhgGcmmk9CYafvkDLBKNGq4OvzNPGlO/O8/
jskUhXsydIXZgmt6mDQcPX6dSXvcQ2zupR+/AcugzVyoAVVNJgNW9vPP4Z5k
gr4a92pcf5XPwhI6ll5cy+kKM08getao1fI+YjAylunQw+XlHymJiYJtpgLq
TsxVn8+9k5luHX8yAtf6xAs6Su2hQOnAFsj65BQ1wGkl1kaUpZ5lfGTxeYeB
jaVhLuNsgtLJKSYh/E6EJdTh9PNw7Dul6eY+eEa/4VtgbYYro7hN1BfNjhau
ytVTJ/tTvQjF0egj772Q5yq+8WunVb8mAermkHC8kFD6oRHcy9Hj671nmUg2
kw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6ATGE/T0bVbvPXLEVqwpHDa3bbbQyDAW2QwplvQeo3mTCptwPKl3Wwvvi7HyQCUFHjQUfE9IIVSGeeY/AWohCK8iIpOqVpjhoTdvz0UC1ne9cXTUpHscHBl1seqXwaKbKiHt8RHmLERHRiO323md1wa6ANzuE0y3jCV8aXCkqn+S8vTlj3Rk0w+6rLUSW0hNZOiYs7xjcXvKYslqkx90zAScchDLHRpZ98/RtSB0du/1LwIRV8huUnrvrKvxvMgeAk3RaE2+k4NZkW0fzpXBKjnJ+ca34CjfUupVOuvuPAsrJzpw8AWjq/BW4/I5TfiFy8KzrJeYLEXDBwhm7oRHFJyf0/QmmecY20ej+UOlqahImMTM9ElSqS8mgS0RzJqVZCBXhDf2lqVot3TKsS3Ngy7Bmf1ljMSW2Yv8a4YRpm50Iijl43gr/otD3UHiXu1T9NdZUV8/3Ih4okviOr4yiBgw0tBi2kYKpJ5HwFP39WZPh2PuHHtem3mVmsCguXQSBJgEpKrqo3tBv60q8W+FdXhqKmfv5x00DNQvrsrZXk7mJOWb0z9qgPJqfNYnd3lR9HVY3lJLDCg/SRhevn9Lk9kQ5sAxc9u68q5aVphw1L1NQ9T5vEInklwiGmdlqdyF3foib3Irvorh1UB3KveV83jOfgykmVuRPKoy8Iod8kE4HLzkt5g/MGPENVNrn+KZFl7eN9enTdpa/EkXiW1/tMcTEknARD5wZNa9NUNawuoaZswe+LwEMcRDj/4IwQY30WWqlxDcqD0mZ5VHesKmiYT"
`endif