// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
shyuHrIQ8/eKxcXZTL96bZWK8KAmcQZSAWw9JRpbITAkP0ejpGXLrbib7pS5
tzBQb+SXE8qKUJXnZjnImJMcr+E3Kf6arXi5JlXdSVVu5a3WBsMW9Fl7ZJTs
AAE0gBSElhCWBMKB1V0nNWJGJuHMv0vlQBgZJ0VL21UkxWpnVFsZn/rZUDhB
Pa2tPUJzdzpmZj3ejTJCVZsb2kTb45hEKDTytOID3gTK4adeZcTfxF1y9Uqv
yGltJlEv7SwKwQv1I5Z8d4mOn1pqcD9A4awQa+GJcxszN1fzFmxSaJoWecDY
oiL0gPsMlgF5jrjv2dvIRbXlyv0m7Nv/0tOZw/Qxgw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R7tml8Y/2DsaKlE1sxJKIjj+S+8vmQxNlFAHtz1d8+PbODpXhO/h4EAchIRX
YUWj6Zm86+sf3BUvbFdW1lo/pPL1Uvz8joSURWtgRP7zGRNBifoIvTyb10Mj
kfTcsu6IYt+c4A7UlJENHyzbxWNort1K3p2AsOqf1xw3ZVXJBubkGzVsOdaV
2vFhaSvYHjMzsJrJWecNJOJ96lukA3XSO6j7LUmVVcUlYMYVD69FazY4xhSF
1lORrG51Ixa9SuUwFmsps10xC5ztZr7Aq2JwVt/l9RflKEaM/SowZqenWZX5
G8+LlcHn0NqOLJ2Lf+R6sF1soQvMl2k2OfeS3dqDWQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C91yA0C+EMZcGPQN02lylCR6Pocy3nNbaJLj3sn/tmw5lrW3i17vG2shTFdu
Z/dUZrEscaVsMzo6tPuYGx/HAjNo961g2Qu9W+TVceBo+0DsFB3mxyTDbMWs
UqUXDk0cFBcmiCwqEnCjgAUaB84DJ2nHOfBLkQgR/Lc5ATqJKSmGBRUegnzD
gpAbjIELQYREXzEO2KXX+Us5f85RjpMT4ZEH5PgbltuYACeUtBg6PVtzcOrE
sjxtNTUVdvDGDy6ltP5KLcR5SZAUcL9LC4d5kedjlzaPSvUFgzZDfuQP8F7g
KADc5OfvhSbtTi+4wSqT4Kdz5hkWio/gvAglcMYG8Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R+ZEMMmPWt6glaro6UAb3C8jBoVOyp0bYrhmcoZszbzZK6vZ6xbp2f5keVCL
iue2Ft6D06TgeqxGngfUVMPo39nPCJ1Xj5+MXqw6Ue0EN+734JVeUrZpfmlb
RlN1ZMh/aNLC6OZVElXKNR19TSd43QU1Z2T2v7JIcd122r31571Xmb0sRdCD
EvYWHTA5ENdbpHmXhDPR4YO+U084rvUmJiUWX+LmyvsliEOxjY/ufvO5aOCZ
We/dUru8bQbfV6lYnCn/g7XxTBDDi1B2SHEqsnajA9XPDmxcVA+WVZX3cMgP
bIsNIH6PAjxhWlbTQ8CARykSi/IEwuepR+cjB9zyWQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fwYf/aDNzM63nV/taCT/DW3Zaq0pHY+EZZuMQKTPxwphiXkpnTri6bOkCsvp
V5yJVF3Klau5a/TRstNNUHBEhSjQYJhGoaphu5/eQIZ+joBrHq7iKrmD+COi
AP5edQoq//M9URAbz+n4mfdJalAeDuLdArXsGmEbA/nL7rcb/o8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hOyBIhmlYp7ldOb+i9g7oxzGLixHN59bXJ6qQMyji6+v2im5JmmRVggVevfA
8NrisTuSmCt/OC4djODPci8h7yALNdsGjQ9gpGe4k8KP/wYWjNLLjSPlNIH8
tEJ+QBYXh5qJ24vyAkvBosftH3tl+wJr5dqTrZ1V5JMxUKZIFxBZS4wCqXMF
w8oRF/J8ZTKqjKqk2FpYzn5WS22kTTRtO60XMi4SZL3RjMf3UxYoGG4Ar7f1
QEiOWbYUZtdw4Qn32FlQOJmi+OODyFR7nwP5M56wVXj8WZcVa633HLFTKtPN
+cyWFCqD0yOA1Eoqep0ShJKdkQnyRMvoSmG4PpUsekNy1Q0/SPE7vF4atfbu
dzhubWJBPcKrAexq/Es2INnrRZx7c0+QkuFplKkfHZtpCL5eT3/MxmPYCLUV
jXcwuEEyGRTmyFYEfK9xrEENseVK1ceuCjdXAirycpU3eYfTOKsUpsfqL8/s
9RRmhjjYqd7iSRnI4Pw4B9akAMc5hpgR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jNn0aXgWFOCupJudAe84IUwwfXzq9Hc+oYVHHdDtnRlsNYsv7gbdbuDLO9IO
aQBOQVjgTAFMByCfz0WyP5Zd50Osvuqa1Ao2vrRJj95mwtGzSHNovAlYWXAJ
w4hztXL6ACubW21vv2NN4W+Cb9dUAWgsOwXMbADJ8u88djEHSP4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nr0JPi8EG7YooR/22d2NCdo0/w7XYmtWABCZ+Viz4P6nAM6pGfde0KkLKWUg
njJfhH4aTF//dO0J+Uk4m11q8EiCgOwe7bn+6dXj0317JyJjKNWYCG7jZ/wI
JwEhVDPkbgNxgC0CZC2HblqAFGKnns3m4m0YS9mvcYOR/6DPvww=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 206208)
`pragma protect data_block
vbNBs60ksFK8aUEpqDqFppl6OJewnHsdms8C/+lOq1EIaqZ1xe/lpAMSbx+t
GkFjXHPLlNBgh9e6iisiYmOmTuqLO9KGU1SDd22B+o03DxjEiyiGS9EkROZA
fArtpufHs52Izdnxgn37KgGnf7ugrreaKHlrxmriaJAISfKybdVbpqQhOy3P
5gIlso+xbudqymOKWzB4kp1HRtpVDHgdliRvDSPvf///l7BTWbrQwN71Ksml
GOZ+BnJ2b0SVxo8+pkQYDDA64Hvvc968Nhwj2Q8gOrwFybI+2uP5KJmv0N7a
KxkG0zQ1EjWVQ6XezKwEdu1Yyvq6j8gMcqLEBVUrYM1KpkasaK/zOsRdYVJR
vwPkj10IbMBgXknrsHrP6n0MYpf6xxoIw0d9Pn74u+QLL262kWuszG7raaO8
JK1FpbVjQ2s5CPu5ZcysP0dFN+GBFhlWVcji2+inUa8/BN9/SwpPRvCN6hmF
s68o/8po4U7+WW3w9o2MilWQQP57Sd8NxkbWJCnkN/Gx0yMZbWXSRp97Necu
mAHaYY0DkqCt0RR1WKPKu+ZZqcBB+jOPvi444VrwzF5Y1/aUWQhYDoqHI3fO
ir1idoiHx+AnukJU/VQv4pH23wyzLk1pTueEth1UOk7jm/Ku1obyaLfmNpMJ
MMfjDh69REomGJhPTQJZWwafWjmxhp5ySdXsNj7udFdl5n4SSZzaOxEmT+Lq
OGnd+CaiRRmlF+QxcGAtZQogR6AY9BasGZ/dU+d80uJeDmea0XDVsioOl0OV
QyKG/bjHDhKij3O2vklzf88+oqb+7jQzeipwaOW3MuN3LA5Cw91E6MSqS37S
6WewlodrAeCyvb7492UJFWQBQco6MDzB+85L8I7c42lQ8NpEUWjTZQv8G3WW
jiMFBwUulM9p6Jaiut9SX4PNw19WXJOslFionV0eMX5GHJthHj34ULnYHuzG
jeEkl8VnME9+hotWf5vqkVufwnbIOnuTrgtU3VP5fiHY7Lm6BmCI4zzMdoVc
hmsNhtrNi2+JWuCfOB392huZFy2ptNj2hv1xi5CF5Ipd3Zv1MiQJQhn5R+Th
CUfiNoQEqFG4A8y2tmqkBZY1AklwRWRrtD7vnnBT/nPtSe/AvYBvk6LKT6AX
Swle2fiBw/LHW6dC8XnGV5+mmeSU8BAfe7wrM+J3isc9JbPeBuRrV8TtHfUe
TSyGuvKPLO20pzgZ3qu9DYmagsaC8gLtvtPdvhRJ+6qvuVaUEQlZLl+M1eJf
tWIRSEo09CABv9O+9H8P3PDLeUHB7tcIRmxviTzoBSJxKaYjkSxHFTppRoeq
M0DkilSgokalt+e8up6LUKHtyvMLIMRXbIGFXvz6/B4M64tPb+ezlN+8l/sH
vK2bNcsR1+PnfHeFrMyZIJ/gQYxuW4PPFullWwA7vFUr8yPKcObwK6zqQ5hN
kFsMDom7zYCZywOkd8cpil9cLHJmr/Wsrj+XYmyIm8BsYAUF6n+o4xMwies0
jCvpegYy/pw8sdgbBeACbeDjdKqdQg4qBFn/LVJSGQb7yZXA4RxvYTOjT+RV
cs3eYTyngtlu0NzwzKg++Jxg97wKNXlmkNfz3tJ3CCugLfwxFqE/ExOj6MLs
6zIHP4s9H2fO/auWQL4h1q4OTeXHSGqhxH0RWdjL00VWnENZKQ1TnLAjGLRS
l+srTX1IJhS2UMLf0PoQeGfyNU/s/BSQv5wtuLR4kROQb4sVJZM0dzDswKI9
70iXm32p2K4YCYsDoQI+qp71BbZdY6+5TlAn/jCxfqVDgnEFDwwk46+4W58p
TnL5N2BMlMZ4b8G546LhpF9bXoWNzckXwAQ7XDAzRBRiIxOBynBTarfXyc4w
Y2vTBO76sVAL2GV0w9pkEhoDqFYQCSQUBUm/uUoEmkK7eH09AddZBvbXIOJl
sXMmwo1ajtCNl4wUxRb5V/zTddveRXOMAVHtW7Cfh+d7jIURPp2l7311AhNC
GP4a+V2JgRan6fFS2lcBfuyrXT/o21+Eg76/Jv/O34kfRMluMXCeUE64bIFm
5YIyHEe6Jz3sej1TW5BWQ1WvYi0ORcp12dq0r7qZNJDW3NTtMuXlWmNR02UI
vZtmIyDJ/X7x94I54/lrQGHvNO8imWUJkCX1uUC3Y2QXhSCIO1S7kndaj9Ca
QVO0Rne9uwH81thdk7r5m/UsOmQXaBs2bNdWP0I9yeVGyMF5D5CmYG7wuf/t
WxM2kA35Im9PgUeEP8LsPbrd8iCGz6dHCZyO7OJOBv0Q5Vvc1hBoY6aP+9vf
hVMPEDGHhVwjYA3O4bRQUjEu1JnIEqPGIGcCT/BOCW6F3Adp1C7vgoNERIMf
uXaPrvkBoenDZfX3aMzmfwTy/XJatDpYaMFOEhI+qMxVAOnHZOac1cRGKWbz
vy2LjkzjTH6A0agH99w9aGs/Jm3wQen4CXK8nh603eHp8uEcmKUhB63YeTWJ
lxqGIDt7kj4/qqypBT9n8Y/KFwQfaq/FMJRnurjcyOd3pXwwmeLZA1pxfPe9
X6Brgup2+atpkq0P/2Et+iqMNta4fRL5DZwIXue184KPw7yPzzehHUSyIxIv
iF/GjMMWEimkZ2Va+W8BP12gD8/MMh/C88tcwdW2Sqyg1bXTziB3bc1c4Pon
jo62UkY2JcwE7qat17UEsLi9XKsfJ92WXYNJ6z63m7/XNDCg+RMgeT8hIX7B
UaaKqNFOFv2HXbJZle3o1jxAcnfxGq4vO02+0OrZLUM6DfOzmGVQlbw1tKPz
OTjja+KqyclXn4XPq997VZ5Orh60G/f+mpr3vLyrV4pDmJee2dUdLQ5A4il7
iPHS2RqvehQTsaHV+pM5Ch9l/hvgxg7MGp3wuWUr0pEyWBxI0qpoZhPr9Hm5
1iqgZkgVu3Wzq8/euMRImfUdxu3oqpkRhBp6o0CbDwa0A6FEI8b338qgdjZB
nNvbYW3BGMAHAjKSTx27Wh0CyWcGIz0hXr0NL/BFMN8BFhFX6eoQza5T6W+s
5VAAo2UD4OEQd4FVxLomLmz5UM9EOeXDdXfnjt8pZXahe5rgwGZnC5Bh53Iv
TCsq+V++p8iC8uZfM5M+ijhO3zqRS0TTIVkR7Rp1BS0Y6neMOelM+8FRyD1i
F0kIR5uj/BFJ5HB9DZDselhy5LvoRs/KY9DLU3QIq2rT1zVINifZ2DBqSpPk
Jz8H8NIRxMM5RKzzkzyy/52oc29df7uCTkmeKzFUY8ODThMEpfs1nj1AZVEu
9Q/QMaviw+2ImoGAuLpaQ2eCwZccGWD2BhUiHCs3XaZQxgEHCFX13bzj29UP
hmfjBndeJAQJF0IIF+Eoez+U320XvWmr6dONcBIxT1PqNhHmLFij/sftAv6x
dFwF09LNF7GuDShl4dHCDoqCblrWRu76d2ZD9lShwLnkuL8VbBdD/TWhebNU
Cl12ShBPpqdYfHr1nPz2meb8v6oWwgTWv1Crc6KSG0o45j7E5xXa9QihyzoM
Xr888276aigHoilUaQU1MRAhr/1WZs0l8DEl7V6QrH9egc16kQAi5CG6GK3W
Uc7KnIeSBP0CYo9b5cz6hPLYa7552lhVgCZMpQG/doldl0p+0EZHwXR7uFaN
Nm9wXmT2GSV/iMI1NEyPP+sY4JSnSheiDtxnEYlPR1jQJxXsssgaPL+hDWWw
lnIYy2LEbF6SaDI1Jd6TLBLJsNCSDQaTyVydLCcU2Ugp1mD2WPraPszJPzyh
nXAO8mvGuhmqO/P1cfaNl0PNDpGAjbHr++tH/fHAsvQr2NhQvrf47uIc+//d
w9N+t/o6En0LgMAx6W7xGMKKgREjkrIWBOYyATW9kwN3FtbTf715TbMh9jq9
yGQJyGflfh21cjpLqUjrNZnKytZrJdbtbrO8RcCciujixNx2bvu3rSftvMP+
2AxVgZNaYXEIbxvjfY87ep5rjugaM+NQ2ZSIf24EtCHbU2BYjUMjrnJCa6Pf
15/WY/LoyD62yCOBA+rK/fkB9apTZ5EHYHh7T4siMos31QAitRkGG3pnt6I3
eUlozH9ZnL4p746SWhBfjucaRV9DR/jFd7td4jT66kGMdeZstBjumg78OnF7
yFryJ5oF+e0zPIhyJiYp7VbW/RMEDIr4w4xHAS+j5KNj/nZqx4uRytguz0lB
FkJA9NmMKzp/wl1lTucBONMayrQpAG2C6pGDbgoymd288euM2X/RRfBqzzQZ
s3gT+WxtFFcODjKgGfD8io+HWHq1Xo5h5moHg1HBM0TdHyeoKdNuj5N30A5u
W1b7wEUJVAYKFqfK1ZK+D7QlNIWv0I1ZpBE7v8k1NyQOw8qvFRQn2YMM9Pbm
aAjIjjj1eh90/Oh7bU4vHoYdyHNW86qHktdUsuWyLAJslofv+kXIkBVrMVVM
KNIqyDbOq+yLvEluKiuNeUOPFilj757UKOQRl3I6TrTbp681V/Sm+8Snz8CB
nKM28fty8wLwPZ2kMVbNiJrGquXqHxleDvleWbmAj6Uk+iTouCf1pA7XDtWP
2Z3IKnvaqJOYes/WTNjkPFEjn7CUOAdS+gz1I4rwBoYRxVoQ1cmEjpri8XGv
vqLmVwTyeNjJOi1OyyARagQgALtxQwCbfUhi2I+b91/4FoFOOO930gfxnIz6
arC1PJ6heBAXKUsPtKEFhxC2g04HhaLGcT7ATJOcgp8uZrQxT2gKwzGb6gwP
xp7O+aCGzTwBqdOCTCiTLyNSFXGgH6MsQfXbZ6o0iCXqrMoIMBLkfS3jJosp
whB6mI/Jx6/quSRQ7tYkyyUSZrTDiIoGYR4PcMpshUVwqJzCuRQFezqVc4xN
/AiNxnYmBp0Sjjh/wUux9tzHCZCJsKCo9rSnvuh1lfuQeC6zysxK6jRbeH9I
Z20nNf99hS45y7CfIrv4xHAVRX7lWE1ClugE9NOC5P0uJbXCtQ4LgVpkpCKe
5AdPDqCqDWMSnwW/QpWKWPcsnlFHtZJbRtn+OpH2IV8T8dDd9ZQhlqixWA8y
w7XHuHNUZJ+JkbMaCX9/5FWsMkOFP5YKGsTi72lR0KO2vZF1rIzl9X43J2bN
copQv5RInOfmBMDByPkJEaBWhEW+zifmjyqpN6Ua/4bDdsK52bYy0Zta7u9c
rC59IrJ8D6l8bZV4NDOkUhYuPwGZdyP2+UUgazY0j90Pva7q9lKh4Ys/kJix
QUJJSecntnFRSkOlSEIEIqMvAkc0HB/S1tDCz5U0f9wK6L/HbzlgWkknjZyx
DQna1/8ycZromKZLu5tCd2Lo2PFQRX+Jo6xekujFHdt0mFQS3qwBVmikqQKK
zPn1HMczWgmCxFPjpwL14s5jFCs6zXSTNZ8s+7EsMtyxj9HQPM56N46ahs0f
mAuusjuM18qHB6pVP6lL4VJpmcvaMAo8jsnT2I56d9H21WCSWhnEFKBzDJXf
nWoQLWn8NkGdElukEhj2CjHyD4J5KmvginiW0qbUHxsdv/hgFdiL+II9FIfk
zwghEBsmmLYanF6ROvdISxE90XdzBngxVekbpa7dEaJCWcThoaBNfiztAOyv
BVT6tvZSivkNQXm8vyitEEee2X+E0kaqg6r8o2AcMncLzoT6OM3UzmgrY1t7
vYSoF7pS2mOHgGbGW4GD1L+f1G8Vn/r3pA4TccXysIqrmQvP5x/mHc6ZNGcW
QjqP9io4E+5v2GqiPQFLpp882AWWnRt0xP0tEnd4Pzu2A1ndchzeKXCkYKsk
wBOEKoGY9T4XmGP3yQnSvyCxdjER4rv4NRdLg+ZiLLE/nGmCSSLi/t6qIJkF
yz74z8D3MUfBW7hP0sJLG4K2C8iRlyEKoSpJBMoMlOwan5rKubv8GFjwHq7Z
ZDiXWyx+Le/GXGHMqoJ5LZ/VohKMWHUQkXORhleaYisvLFTRgD91evLzM19t
b2tqrMFBtrSKui258if8ltrUi0E3v2Egtr8pPIfriCxmDUhK0bLKwf302FS3
VB/yOTTFWWjHFlzvoQk8cviCyW2Jd1F40nLvqt3sjeh3+sSlSl4J02m8qjSI
5Qh9jA2cNEDBcoauBWlqY/D6bU4FeZyRPr8wAtnzeIrctb9RMek7bRhp0CWh
bsvTG0+4viY/OL0QrP5fXg8V8aDEb4sq4YGJQCjMmQ1eWFfdr7OSj9pcd2Xo
VjX04jWoPhPMeGse35t0jVTcyHzV3u/HBJXRcS6LAZXq2DDejqagsM99CUix
HmKrkZlKxCCBrdVBsFCNXLtSkBEeze407CGAKM2gK/mr5+bABU3FLyvtluE+
HqOPXbnY3NtDKC/Uw5S5TFg2252opCYra3khWqZSmjFSBHZjYDYPLSyQxJZ5
naHNvZ8y4U80N/Sbxab9okeO3L13aKKVjone6MKaiN3aAuOC+GMbbChxvB1m
l6Y8WmS09AAyQbae6lvrLaP82SO5+rKh5BPU4+vM0W1nx/6FddBuYqyjHcPO
GyWNdMa0DZ+cVO6sSrgxnT6A1FCg4AfYwgolwjgxK0D5lO3mwZvRwjpvpQK+
0ZmsfcApB5F6H38EdFgyJH65uYvM81HNJ0bHteUU/E7wyPajB0YOxB0+RbLZ
0U/OrFVrS0/R3IdLFVaMk6LBel544i+usfRPZKWWczZFroFc2RNLj/bLTM0x
MakQk+qi4ZRrEoTdEMp37sPWsIXbO+W4XqAyUtgnKw9u4V1QRaoOlKxCevsE
vI/oCuZ9P9Y8ciIHMaY2JnsyF6QDijpsA9L6DDogTf6EEO6bS9Qgv/XLb4JU
HpGzqD7OTAeyOhZt6k75l6xQRYjBDyf9VNuN3U0s1X5vH4vMt5HGdPGTOR7x
oAuRHmCPzG1QdH4S8i/GPsNqgcqoG9kI5gzepfhO3G4pdz4XWmdJSdZV7Xmh
t2jzOFGkJBx4CQNm+32KJeIhgTtZfNYSAy72PxBB9dKB1g6nnh/QV8SIxWZ5
u4F9rMUBKIAv0uMj2+nWxV9Q8xTwh/vzZzpjVAFTwbiJSwL+7a7I7w7ebd+r
C4kZw04aUCrl7TKWipIuhaAAsJM1vhAz3EKkDxe/srJZxFjNhSWEDnaWQU76
JI7IDEMaNRbHvg6h298nyxFDK0DVRFVm8bvS2SXKE8syDaCmqHavx8O5pgHT
xvyfo9MRjii/cSiag3QCrhTPREz3/yb3c8SomHbxIbZLY2NKJx6ScTJqjMKQ
sm4KYcseYvBxPceJWN+vfiiteonFM0INanfPY99rwX7eo7LPkp3ZWlosGjNu
VMC/r4BGquG/47wqQn5zcRG0r2muXV0CJFsLR+kAGvqUgQbrYbKS5MkN5EgM
CDrS0pyuPgveqKEAhSGTrFpeu5RB4F5HUxk759n1K1MvcnbHyvSlEiLh66yd
zFfNgWbDyaNBkxbJw8KY1TZMdXS5wuKCGhO7/ZpXiSb8a1+qOM8c/JFu/VwD
Os9WXEYiHvm5SdzCyZnyRZyuYspCJ0J0W8IJZQpQFsUWustXIjLtemXBX6L2
wD/FdLhcBAMzfyOf+JqFwCpLK2NbAADal3hLggqC6nnsX9+hRPUYtaWtNFrl
n7xwt3iWts0sFfWCS2C9Mq4263lHey4vW+206czZEIk8BSfgbAddxI5PSMLZ
YSpwYv/y6t/ry5QCKYU7GCdI/L/uGMrVYS7W1gbmPqFIo9/7/oPE0JPGdvfP
3/CFFpwLFo+E9SjgQXbw7TDhUXGjz5j1cTauwBd81ZKFnAx9MBAWRiDHBQxu
AurCjJhqoNG8sw27zABUlIRIXEBb9qzc1nK7WAOrC78b6PWMDqad7ZDVuBp5
la8oy9eVEPFiMwo3+zaA4mQq4e+aBFAUZC53I+EpWg99m1n/Yiu0fVxkd1ky
0COc/9IpHc7t9lfdxfpxDfWC84u81yMeJo0eaD0b4yCZzGRIqZDpY0GhzMrK
rHRXk6o+dzGoRiwsrUn28gS6M8h1XUQs5WlhPZwZQ+az5OOZ8LmGmQSXMr7L
Kou15jnS4M8mHCLsX/4Hm5U2ABM5yVYu7Pt2/h4YXKC8T8cYRLUNCUCKQHfG
+KTARNkY6yzWeH4yf3wPQBNjjaBgDTK0NoLWyYzWJJ2ysRzBZQHthddOk+U/
fUVrfCW8LKp0yN/CJAtboPX6KC2x6aT6s6FPU8sLTt5DZ86hluhTVJ8y8Id/
NqMSvKbEQFGQQINc1ULCi2oG6E/G6yD8qrbUEvMJ72NTky50AfETn2dVbFK9
vdS6GR7HXoQHipUDESZdkg69d5IO9DsIJJmFm/yLKkSid8k8pRdzDWn8dNvv
sV+hldGvOFf1Bnn03ZAf+mIsUyLKV3mGkq0TuLddOYwZ+fbWTZYnKbiHyNZ+
WBB226TE3rAxEIpCILlKS+93m743oR2yQ1AcSjn4QjQ3dSmCHixnBaRnRovE
aBHSqCGXX09q7gcANacZMX0uoDZTTssidJZbTdQ3Hl1p6MpwdhNcKJd5vzRE
vssP81AP3bN0gEvhEcGPH9uLuGKGj3ZRjeT3jkcWHok/Rk0ttETEXQkd3y4N
xWvHChd4M6eDDTNetC5LXubm28bg923hiUcwhCGq3pWx9mQE2m/I+1C11Kqg
pdH3niFLvW1pL/6iL1MisvsbfW1ZauNg7Vhnb7aNVqKh8MOfL66WLyTcxh2z
tDQILFipYgMUIdRBvVr2sCAVG8EzBjTcKMW2vn1T1kPfaHHCTE/k6ZKeh179
X0P99FAlGs7M1EuhQOzLrH0o7oUcmETGhsr3Xux1ziPI7u5TUw/0+LjUJ3HL
72FDpg7cDBaM2o8CPu7n8A7xTWTanJVpNOniPPXemBEI28sk1NmKGlIeYSlL
AL7j7nfZ/Y6WxLwOcF9ff/TWJtqmq4SpoTQKYaGCJYK27yHPGptv0Hg3VN+r
v+Fi0gGKDKFELfXv2zM2Hw7z5VuNhUHg5XC81dKlg/Bek0VEdJKJ7zg0qFwC
bweUnco3vZVmSBaYvQXfglrQIDccPXxxhMKbh9mHNYAx6qP4yYTS03JeeObb
JeWu3VnyuYWaBVzW9Nw811b6inefw+zJYFal5Ceum9gPaQntSOTu9XRq7mfK
1yvQWBy0mtzUGS5mdlRfv0iCJUQnZyM7mG6bSWdtxpwNrubUj4g/b4hoq3KQ
yJ/l1j+rtQofVg//QZeR7E047rHxD/hU2CVAjHSYPoVuYVqIS7th/534MM9W
sEUTZqEhczFwY+IZlPzmLyHBPFpZe3sU3SCi6tQDNZUUOIGw10GB6IvBz7/7
x9p2g0nU3a6Hd+xRFSRPPQVjbtmTGChbefeXKvDPo2AUzY7Eae5thTX0/9Dt
NA87vKbazV75JOrXzi6DD3WZVed79HfeA75ktNgk4V3CQc013G/8T9tZZNWb
vrbSW16pz3OXw7FgEDn/cXQQp9oGCrDNYzZGdd28cWCF5vaQpJqfrvrZvriz
GmcDNJI4LCksWn3URmMgclkjTYty3V/FsuMR1nBZxIl0Cc5U6rkIHNZarJ/y
SjOXYElC5E2qSyCUGKUzxhT2otwXDgQMHK7UP1q1VA9zCUcCmlUzAcUGucIs
B8TAP62TyXC0z0fsZvw0VO+VE2z4ItklAVEBxGUr3WYSwv7rEzch++RJVGQd
sijR63doo+wU2P8ZHZf0uTeyOf2ROIGwdnw4fEs+AM32rcDZm8ret0zi9DOk
Epetsza9KgwMBDXLJuxkHSH1zI7iQEGLwBv8pLeP3uNgU6QGhpY1sqar7uE1
D1vLbHsK5ZKvmyU0Y9vonCoS6oo7IdvttOBm7zb//8bfktFkJTB4+gmBkana
fa9lxCMH2soOaoDdhxQ7lxaFVsnrH/ebIRk2chC0kGT2+zzsib5sdI5xD5Le
oHVy6vhY6q11oNXUbPqVXSS6OqzqkhD72y74gsGpqZZbCUzne6ZBCKcwlwpw
gnE7BlnXUZAOT9jcdD2HplE/aPCM3n8FOHslANB/tJtGYX7QXjmj7S6eCNnJ
QIzohns4Vz9b15SHGfCESlWTMOJopvpA3XOwJV5g5NP3OLxGIVncpldKOUWN
dJ+yLuzvvhmYzzvEM+z89s9LGpZSTdwV483YQ3Ty3npaSdZ5gfhzOUf0muzA
iuvraPTJPmWXy1gf3wHODO1AeFlaQxyPYRoNO3dVPNgsXxpijdb4nTagc2Zz
waP0KztgUkkarGd1CdqlWLYwFLXUaFXc/oXIYmIHwp/Xg9ZFZ3jTxgCWUxbQ
NblCkrnsH9zs2h664mqT8AA7U3LmxssmbJltIn/pmT9DWVWvdzWGjMRt4139
2i2nkUE1xzFRSbfPg7CjEDBWklohhd8J30AHFGegOMJUmb/rPDQrfRyS72RD
0n119CpLdoXAig/a+couZhULxL4DgsoP0jG6osydyGRcnHJucMFkHzKnwLU5
K20nqECb02etrIGmyyDuG3hP2cE61aXBrmCIw6dTlLCEVfGayVGbQUaeYdXm
itxGijc4XrIO3WIomXZM7BW6vv3/at1/xOlkhPsIDFPEnR7NenTJcV3yMe7x
LuKAPAYArwqcWZfdhqr4AnT5xF/TaW7OnA6mjTL4POJz/GAWG4k8E9i8ThU8
60uuDbWPyYY4aViFy6piuJXw1qSIzVKGuWDBPndiPTRYeby+DcfHj98UflEV
ci4+/eT/Sk+60RU/83LDhJhB0jBFScPX2omEp82EO4cCPevxusAD0iMQgncD
0gcJJzhVRed7kPUjsa7pwtF3izk1JYeWnAAdNpde+J5VH+YeyoWnrBeb8jvt
lNUiF+il5hSNRL9u7MR9qPV2Dugsnx9M3n3fL245SZ6MNDtDlW/OaVJcR5vG
cp0h5AHuDZg1CKmFd3OLnfQMwmDqHF0Bb1L/dUbjnf2rTZCsUIKM0nBgFiwL
uLTnFOTpvan4g+d0nJDsJ94PUnbEwz5I83qXZq1rQFeCv5KkumLIrIRi1Vf5
eo3TWtxbxdYy6/y9tNfKvufLvbPsS0CPZPNKIE3W2VTXsRMvh0NyC2ExmFO+
Un52YsS3KkOvqXIr+kamUz1WcR1sL7iwM1gJOKZOpXN3WpuoYdQTVyu1vdnV
uLfXHU7g6D75wEqpLSV8DKwNGA3QcsJVOlUuRf8pHqJUTE6nf56pxLTNqdC/
5Ms7PNLZ1SrdwrCT9K+cbBbmKBQgzLN32T2Z3beIcOpueuot+D9VpUi87vcR
S7KlcR4gP1tcRyni+tLbRWUiGvdFf3yJUirNs5niv+mVYnn97hqPsqLfjVUa
8jJK6pclRty2tyoFfQy1eamPcF/h8NLUhUva3ncrysl4rP54xd1RiGZGrHeO
28LkHIdPEDiPK3mBJz7+pjEXREACe5zAakzpm+Z5oCy5G1WqD8Mumii8UgFn
DQ0tt5bPm9t0SYeCLYl5dXMbKQNxGinqD2xH8NTwXw4A9ieN74msj1pfWdJG
9rXYfEg87GkqQUUFtuYylOD/wNqlc9DDlmcxMumLZUXVC0fb3y6ATPEmBTaZ
aX1Kvyo253aqiTQLcYbEV/+vHbabl74QXbVg/hfJS9Ih+eOD5TsKg68xqihn
PY7N4LKx9/UNzRUE9NB7IualDEv1QJP2D4h4R7mTmYqwGRsxXEQBzqJ8/XQp
YiRH+zCqZc39scwrLmmNYSmqrNoLsfni7ZAfDtPx3Q9/VPK2VtfrPCYOvGau
VR1L+4IkJFihY/+GyphTpfRitgXGQ91K7P2eKKNgVXlBu73XcLzuJAAQNWNl
4UZJi6mJhWxJsrl4GgEx+g9lFkm+95evgrZNzr/b8vMWlw+v206NuDyGAAvq
/XkWGQDjojSTcFquZqV2crOKlaZdy4ECWtmYsc1ORsQIS90HS5tYoUvHZ1H2
/XPqf75WKDNdEtzzPM1FDCU6p3bGBeedvjbdfnfducNYOdj59F3af87UQ0Vm
63gziHY4lp5RWe7Pr+az/5l0sJ+xkjrbhYutC7emmKHH8IcMZCNVyNYyFKjE
WldUGto3/wAeUbGhfyDY1LJPHRe+OYjgCDxAdwz3PpFwf4KNuF3aeak9R+Bx
kxlYmNRY0NG3mt29ba40yF6wYCe0aU2Q7NNEUn/UkCasWKnt3I6mDFKa95NT
qTAW4pcWoMm6wasqTijTnwtWTT0/WZV6N52nPcgrrqQ3fU8A6iK/U+0ukrop
3A53JILvdMfrSVrjmqNH+ywlTLRN+cg2xfkV5ra3xk4ZcO7yy3NLPVnJXjWr
+qE3emtHEG3mHNzSaRLNjTOwoVzv00sQRpR7JtjqjF616DGugD+D7AYx7Ch0
WZ3B1N8otFj1exHxia1Fyp6SHBQrn9TJCsWjyvqTN5QoUqqFIhf40wlxaVRO
i7Ur6WYUghZYSQx1tEiQ3ljrKtDfh0rMC/5wSTQPJkASxCcPQpGAbcG6P+rW
0DstelKXKq5qjQ+dPOS6yDuduW3Ep76U5HRgGYoozEzYhF60tIofvPZ4fMti
orVHn1KHF8LRfUdq+2300PzBbuuF/wq3vFI0htgydW6oWUNHUREHpZkaLIZg
/S4Hq1Sbuu/thDIu+PKrCkPYtvkmHVJcJtYjHxPLTefRQlFbuTqJVcr/JbP+
FR0orEPYZPX4EA+EMTXmukkPZlHm6mmF87i8LDOWuZSAGm4Di0o0OtWCkhec
ueB/oKIWoDMEyL0TpIDGjmqD89tWKKKFBPtFH731n+I4hFunrXRqIPLoDOFN
k3TjqnbuuOJMgfEp6+LBFtJYWltt0hbLP0TgwSCSqExohbZzmMvDnsP1FabD
h84jfE7xCTMoNQpmc85Jk6H3G9asoyPNDOyCzkOne/DmAVrIw9M0F+5szskg
Od6WzdzGWy5kmyzt3EY2D2vZpTMGjjDE94szcFDUXFeVwFSVIZK4ooL1doVY
w+lzjJ5Z55lg7KzJbwDT9iBZfzGy+P+CgbRTPobYqzhZLVcYQSygMBBv1VdV
+2XiCSpYN1TAlfoBzaTWZA+YnloPhWjsVR4AMNX1bkNK9PByOD4Aefs7suDs
dM6hzCVVIU79LJlgtBQ8+ssDCLBZgE0Y1gvvcG2iUgm8o0hDB7JQx1/LhFzi
uM07EQcqjmnV9NzqMW7ActDTYfymASCTuovzjcWeq9LlYZ4bxNydZMbRWIA9
9Sc2wqw7NPKUxiinKh1d689NO8MMXEpoP+swPgia/aPSDceWNYVulBBmB4je
tssw/JP5ecL0XepnmQeVPmvfy/4kZnI1CW0DOyZ7BLQnxrG8hzXu3cZz2nFw
8TCMwgqIRNXQt3JU9iMd/PhGYHCHhmHAPvTGS/fVqH0ZdMjAyDb7vHPWvUWo
2LfGQANphcpxuv1YUZsNm8ptCkZrt2cfZ8dRnRxYf4VzZk87P2HpZJHZahZj
MCGtWQTx6/XaZmZAY64fpq7cVkrmMcFCyrnSh0V7tfrXFSgcJPkv46UhMAO9
0XZ5gWVXDcycLe66PJuhdBhO9Zk778RbffiVv7NZ4CarKTAm/JY9KZzAv1nC
etH+5bUCCe5Q+GI8+XeJVIh5RUj+tRqw1Te/E7OA8a3TPx25fNJdcMLN+KyN
0Ft2bBrECYCEKiipWCurblD/O74Cfpol+JYXlG+NMh/hhhv2Ade9gkMSKMO/
cCes03VAcdfJdzlqaftSxmd0m9IsB5Gb/+pQefBYdsyanJQhCxS/+Mzxle5B
wttaogdRhpH2IuFSKLDqm7ON0vaS2GyvbU/pUlOmQf2ypikciBfha6DDWcba
QHE5nKH1wEUogg8hZTqMvmXaYPghAWE9xSd1SSzWUv5IGp5wzbQv499sgpHo
0RxRT9flMy/kS3tRg9Rzmlnp1sZ0HIP97ZiXqpgsnZOCsn38Q93ZGNKhV4EG
Yh7eyaLorxoDMUMXMu5ZpqBnsOni6MMWyJk11+B51t9mrq5Mu5+ue5ROFpa9
DOvW4HX/tV3erS0J3hi0ynmPlad4TNmcBoQcx95SFOYEFIca69k0CkpgZqbD
88ZNX4yIjQvMw9d4gMktqvkCTwMVeq9+qJ36O4ja3k0JtZw9eRTSy8+dgaBR
XfuyLaCQRqqBAs8a+womZJ13umBoy2Ahc5DfmAL3CjGxgJZD3K0A8gAquO+G
fDL7++LEiSE5vR1P+mB9VFTD8qWHELPpWlpgiaVl92aiKuSlDDsJub26bCXS
nWveBJboDwKyGesk7xmcRlMR2CloXqw0Po80Xi7BLfpAPMGnme4wYmK80oj3
RQj/ZuEIqCq0XI+7CS693I7wO658N/tMet2WVd/ADEunZNniuJQZrBg+gPCl
IiRo/U0N+xIu9ulsXlIPjnqoKrbWoHDQ5qBUu46lad2Xc4VvtFgM0YfTu52t
yzxe9vKclFk4VXQ9BH6GZ0B4Q49RCUCnzSlOah5DiZtk/P2O2EQAzk6/eXzC
0l5KgPSMjx8byXVav7q0G9Zq1EvUeKejHpgY2D0Abne7gdniq6sMJMIYGPOC
5k9mqWkyYjzRdMbO7oQ4Mie4XPSLALdzBFf1dI1U8UqhD/9Ukr9WPHWoagok
RUC0wCcbSmWS9YYt4/FbK8AjEMDw8l5S3XEHzZrv9tbZRnuW5bHb2rZEnUAB
ysAsn5dHo5JywuMRrUDOQyrIZbwkEUCI23GW+GFQe4I3rUgmV/7VBup3tNGE
aownBLezt+zwk3CZBBkGU3U06PmFK4j0wa8dwfRYDxnvCAltJnDnFvHmCtDa
+3GBiHbvRQFRNyo8V8LobfRNDytkKSlLw8T2Nsbr/2K3kjqTyOKo/uAdfX5q
3f5fZbiPVZ54TxVKaicyi272KlylrcQjwjaDFLg5BLrXrEpmQzjNQALYEoEu
6U+OJYcdQbWkyFDtp9VlHJSb5OBbOG43+nVoZn/CqUJseEjeNFZ/bCaKeumM
qk864qiU2/z3mtYt20nK/VUyW4R82MVoGkl1jc+2Syxn60z+iFbdoVQv9HLh
9jRD8jyri3NBWOqwcdgpYKrHwVKjQGduFdFB/Kvsk3nugSpDLxpuv762Rx3Q
4t7tkMeOYYxv3JcurR20ciLxMwkAzZWiuuvWBLUNdP5BiUnkXf+32ho5jm6o
huXJ5BmxCrWjkMMId6lEIokd4RTKl2jDj2qarawvmWkPQKKvCnedwEVkfbgV
Ab/nTzSlIhOx81SfQyrQ/U16heos5bNEpgd5B59kTusrlhjiJI+smaPotkG/
WeQegt4sO+lvNDHfRa2JRcQ7daD+d06RdriAmYUZA+eAKqzWhNpMSE6X0Am4
4ds/XZPbCdo9zM7thEbIjoDWRXL2Wf8tsvFxB16PO0bzcVhR8gLeR6oTjLnN
RdqhRYt/kh27foRKkndk5Yco//Nvhq8svESGFXLadcr9BmDq85qViAeauGL6
9aypwxO71oDeoka9Da30FFjG/Q2YDvJg1AQBLGJ4SeTprW0bSeSb8kEtEtx+
ewMpSoa5JJRO2LZozFYfrPC6OuM4XJPCwi1MfsdbN3xAdyqkpwNIjoUowv4a
g7xzoQefNzd+NpY9iWoaz47M/EgNG6pe4yT+nbu1kg3nij0OsRuFKnJRp6EL
+COHdHZVkWus57Bx0+EZkTnJCqPfBxisCxRo9PV4hWXkcKnN3sEPmcghBtkA
ItVCzoNocP38CuWriJOwRgrNxpIHFd76kP08fdKw3MTWCCM2YAPzBNVF+YRA
cn6a6BmM+hE/XB+/iRPyEM9ROiWTcx8gJLhMjVrx9uB5evzU85xtYhkZFeSg
8XvCDukwvo2JXepiYj03LDPf5RKuW4s3I0aSfrCtQ9CQ77XciLwrMrK6gYbT
ww6SrN+QBz4eeZo2tT40paIvi2Sz0SoiMs7DtAZOhGYPZX+SXO8V7CP5HVWB
5s49R6jskcQZstQPxSPgC5Py/9bDTaQc37cF7WPBj9K9IqQ5e9iafg5uANlh
mU5w/cd/y6IRVe0DLSDoawxCZq6VO2tvcdJNCrp5bhGIKiJuVmqZ8R/evXKm
5Tt2WAcKmtOmcq367uPqc+SXUwkkq06D3HgaKVwE1svt9oXL+SjOMnhE8Naa
2HEHq4vsnnkPcgGR63mrhwXj5l/bugvSzyREHmw/6wTxvvNvP1uPOgx26ZWF
DepFgsb2TerXPooTmXykjSoSxmr0d/+JYBO4ZE0D2QcyAUmUEqVqEI7XckaB
RRQAH3LpX+bXiyZotXp0uLv/6sdJiZ0cnlyECZbrVzH07Ti+jh6XiitPYLgF
rRMvZ+H1S1FAOeRnp0VcbEXzG5py81TDauES14bVSdBj03aGJ2JsAlUPm8y2
YWpD+R/IJyqhdPaR7lOsGQ6B0IoS4rQVvLfmi6GV09jisgJDWnVNoFXTBhSE
fmSLGyi6kMXbp4Sb7o1rjlcFd8ZULxCW71EsQ6I9Ef+TMk8AUgnFc/ZrCaxV
I26jL19NYf/0dS/pTcfZnV7/SCj5jncwkeHvUgkQekJJFGr39nxCqs9u7AaY
G8BSyIwvwH0XZvHdwGtPOch3WrVMWej7zEQUagv3EzMZ9ne/WWnEePRwt5i5
qsKd+qUnkKG3FtlUIXojv3vAgRxji8FtwVfTCs43RJEXJIPcZGeEIqHgrSgw
OZ2pmJR209izRe8KbXeWFoDB6WRGK5OP8Xu+EzOGUA1VaK3EhZ8W791nowb3
qnRFfDPd1AO7wKaVtQiMlPLFLoidVwgZ/OaEUWnJKIYZ4wN4/S/Lg+j+1Zoi
QS/ncGY+bQl2/Yn3uAdKxGWsn9SUzPqPee7TU7jv3aRMdVKQUKx6k8aXw5Ha
0+L6vJZj24PGnspLggj2HYEPy+J2NZDfspWL242cBk6Kn/hjB4cNUEx4VI6C
v6KVQThQzC878imFNNI+ggt6jU0p3X8ZIWv+J+OGPo2+INS7UQ26xRuGtX2H
BDiKJCxdlig36DjMKYiEGf4c6AuE5IxdvtpuWyYwX5d26xCgpWOuZsquMCvL
+Ut9mZq5aQ4EM/ESfDSzOKwIX55QCgwm0STSGSs834R1XX8/uIual53+lckW
QM5CEOr3IUBBkt+TmPftoieosE6ma+eQchkxK5Y106y2Q5mmeeio8iAP0jHY
mt4X2DPOzR2M0MIruRsrzAp7BeJICEZpzcS/aUDlPwib/RF40pJh0vPUuV9A
nl3ZtXnWZ8X89fcRY0cad4cFa43HlTnT+KcX5tojOrm/mHqPEwtC3Kn2oYAU
3+U1oBTIVghNd2OltI5U4YIZK5d6ce8e21VGrBlsyo4Qu17xAdpq7+3PaMEx
xQVpzIO25PdYxKeuTqhbrxXqO4acPzwnCLvoedoVtYe9jBBE4kw6E5M0N9+M
MBy8GV1+OvoOsRq+1KsfvNOah04rHv6p4KYjcmDQMNap487NMgrxGxlbzAKI
P5DmyeWrFzn6EO6rsZvjzFsHo4KC9HCKOEBxIt8p9Z6Vf5DWk0PFWKm0ggbA
iHONb4FthUItayj1yOm80FaM7S037IQQKLKaQnphvXxE30/nUbyusEEoJstz
y/ty+oFPfsqCHDLrvnQrIzvFmPnTuIJvUaVVRLe+mFNye48TNiyhsPZKLsWf
H9CXjrjhKQu6daj4ExsPYE/4XGSmTGg9Uv71E81F7XEir4fY7p/viwNzKgHS
fi0Ts/KSZ4O6y0Hw6VbQj+dlHwJGZsZyUksRHddMXFO9hzNONOmrZuajBwlM
KCUyz4Gb5GrFIIxgwv/qthZhkzVmuD+RMDaOPA61QSjGMGRJjqYpBe5bJ8xv
6kMgxVOwEcWN+jekdE4B8+pCfr7Bfot7JHvKDmKTadpHsSvWgLQb5CUyAlVl
psaAK5J+f0nSTYYV4a1tuKJoqAm8ABDc6sNo6BzruYQjbFUslRhmOAk6ouYy
dIYpDrDU1wLhplAgtJmiUBr6TiUO5YNYiUTAFfTNCVi8vQ46IShhtuUxqcOa
H4H4qh/DhPNSumnnWOEfGpA47JqYgxqHTYLMQ0m5tXhrJcTqeK7jM8DoUAwU
+lEmuE4YPyt6TZ5aI6eR2HwzZxnZR8u1JG7oTVaut9qCobFqy9g1BHreQWwX
A6aqu1IPwji9skTKNpJNC/c+B4tIHnpEJoGlF38G81HqXosX8B00bs0n4AjO
BvlWiIqYpofC3qoH/wPM8w0NeZToCsMtocTWum9O+sRdmxD6dvQiYP/gTe7U
Ppkjhe3Rl5IEDzikqE/+Ck5OxQS9EBKgvYYXmnyy+lDjBQ2k6Eke4+qAutLU
OeTU3sDdJhLJHGWWsbQc9aub1tW0tl6c1GscrQeuV5Q6SS/Fhj2q5ewCsHYz
SxXMuxpJCSm+BoJlZMzmsbwUenaD47y4t/x2gphtkX7THiQwDzHG6t0FOLbV
0GOi5OvwY5/FVhEVTWPXewv+467TYcyVJOmZRjVkZji6nbUS2cGnKi17GVFK
xKEIt5w/rLczVktEqjplu6oqI+kZ7EvKRVST67JOQAKVoiCqvAR6lkfHeoxl
5+oisdnzRLp3WxUqnBkp7ziYp8hC92qeqgRe11c+upoYuqH3ZzmwMf6WXwA+
PBYBrqNAV4J2URsHOpMGHnzDoj2ApqJrS7c1UAR9ozTqDm+DloiIAZSg6KBq
Y0eGta9BrUlJMpJ7pXJYI+U1Y/JbhB/OuT/pCuHQSwK83Qeqcrt5mUU4WU73
sZD0p4XucLWXyfAx7kELV9OZ3BaOE/WzHzqrdvHNGwXNyM5yWzzMgpMTCptw
xD9cS1zGvLH/F+Y1H3Z8goKE3dESTEqlklOPkyRQW7Upie92ithMPAXMnyIL
odxFlUB9p+NLOuaGlusMWhnxWe+l5zfzodVrL9hd+F4Fd0QFzLvTeR4F81o6
P6HyXCaXaXsH/cyzkmrOvJe0MvEqV0ly85ZsXQN/TTMUjclfGlFocDhIX7dT
JzXbHMMKLA1vp2eB8W9tRNFX5xj+GXqm2hjlP7qVDiauSe6+WTHifnePWmND
YZptaw2pH6e79m6ggGli2K3KDMezwWPwc17gCy8OpAZqh0uvbMrP2LzmxfYv
R+VdGLj0MNoyKzUunQlVJdOH1avV12xdnESj+94ka5NQGSsO6o+V3HsfK6dk
c9lwh25IZDLK7GfmMpZyVjL63LAQal3rixdyiODiWuRBQNpe3h3PPx3LvhKl
SoGg1BVgLra4cLKezQrc1TFrCEMGT5OJBqkfFKjcJclodTqpnhi4w0iWeTAx
FCwTNr1jS5S8+EItQr2awdjj/XrTIKqtr/mHHdPfCaH4iaaZZBwy9jtEl823
pvvD916eASpw5v6vbv2Ya+r6nnIYEa67IbuvDPsSoL76GaOzB6s636FnLlGc
IKGzvPnOzDUOoUupyjxmDx1SBt2+xbtrwJriOcPGnKv/KdpCGA0NaMj9aq0k
Jles18e9RHmrAPxCwLL+cUI0qr3BSJgcmkvVjjOd7ernFz8o2xfyO8u07Hf7
uBuXXCSQ5OaM4RRm6l2vOVM0OprmbBDkOoV2i5+e7J4H/k0E6QlC+BzmpwFE
XyvvnPXg8Yt9ZuRfjd1wycJj2noZQVamzz49H0ReYdkrt0ASlOwwfJbxRw/5
D+pPFr0wmaFSRg2O+VfjOnBlg3fUdI4GmFRjpCzxq+NDoJuoj4F6F9RvER4U
nLCoxMGkiByrYn8wb7HfaDyaWhmh5bb03zFRvkku/00KNqyeTOa9AEbSOET4
un0bSwa8dRZEZUJo/EqYm6PiKtJbV9auw0KwOG3rZDmHENj1RfVfR8/5nWIO
xvmKs3z9GK6Affy1WHG8Ey5NLOHr/aTXQH+bqdulr7yePH+MTlgl7YhQ6km0
z/YE28CR0YD0WuNUVCSEZvA29Y6zfUAdmqTftAFQoIVfaDKj4CDeary2CgvM
Ly9W+3ui+6CoFVPECV6dAsAPkHMrckuAyay67yigHZKs0Lm3ExJO7+ImYl8a
HE/sd9hufFc0IeUZ49dmH52uxel7wWSP8125OXXptOEVQUpGIwcCG92mzF0E
tpa0oGWH86xC0X2NJjH+++gAs4zMKaS83eeWYnrgqnV9LlV4Al5d8i0vgctO
NGJjGwWZCGdsXUcGn4WkpDpSrRGv4RkY6mEtP3a7ZCVkiNq+Pna16ZP+X1Ut
bcN7rP3/hzZyxM1DyIgEvroEKXAMGrLPK9sy6+8ODDI9/Dgqsue6hXM0wFJS
3hcaW6wqoHttaDVN30wRoZHv/7g/wEqoTLi/58/j2YbchecIq3KK4zZcprEN
4yr7iTt8+94ckl+btEbtT1LqpDcllfTRho6bo//yezRguJW9c3XoHGxBddFy
+auUXSxl2eU7d2J1l0A7WYYRnb6q5H4XJ7KIQqpuOQethVvpwMLn6ulzvGWK
b72Qdm5GsTR5f2m/JjufxE4iee5qtLTEZshXn3uc8Jlz5Wi6lDwaPZEqmYWR
5Shik2W3PyAGFDvIcmQFPlmFyRPoT6dDCGfok/oFvuZTrHBMocTXZ4p67z7M
5JAyxeNmJmVN0PmGrDk5tLv5C9i5copf1ToW8FfizsnMiI20DPJwNZS9G7PY
UorYlHI6FwZpHTdy9+G+WftTMGpaEnlh8DMi8m3gA9Ze7HtX4q/A3stc4wXS
QB4ofjs85Bfw0snX6A6GgacxpJB0JXOJjZpqp2mXze0wv11YB5UVGHKijIBw
b9E0eskgzMBwjLBjlHD8EGn7vQ3TODpQBKwFbjDxfNICklYYBX5xFcc3AY6G
B+mdwcAxXfz6EakF+U2kG39j7mXt4ZfGxZNYHFUR2ceYFSV/COylauD2Y4sa
7rrk3P6WLP5Wa3HgIFpNfYSMQJ5C/VGmKPx2vO5TPeZePKCa17ENXIKOUdfC
fp4kBxvspGfulJjlXxHkB20VEl4tZZOvJ4S83SAHran7DVYfOxdRcb78fh52
6vLNv3GhCTmkspNAtsGIxlZRYLwiO2+tTZfnQ64j6IzZ6qhMw4P7n4ng4zPC
MGA8oCzRf6aGvAY+4a9f772dy6rFtLEU+hhlfEsDhL4OjKJ36PzzpM48v1cW
lVmrGUm5YbbYeW9btVGUcl5UnZy53JLwArf0SFp3zp+AdYJsHUTNXw4ticjI
D9zycIGbZHfc6fQWY7vQufJqToupJlEIec00+QRuP0qcau9OiH+UnPpx1EpH
9TKk2jiB8JQskw7AHIk+4usLroYGTvo8aaiqCwxrReb4mTXApku+LKqj6gPU
ECgQvzkWIXWRF5gKw5b3BmCCGKi6qxXJb6wcrpWxp7xGAqt3PmqTiyrYHknE
ShfUA81Lr6aW2Uvby7GAbuloTOpSaSTor+EEOQgeyj0fxiIy9qA5v0oTw1HP
ZmZ28JIXnpJhRKUq7QcVCg5f8bN5i8efISBkhuQxL+QOY42AkFNjkq0n5deU
107M3q/gdvRmGTX/5cHoTzGJB5sIN9xDOsFT2MR72V89gqQpN+WDw3lllngw
k6K2g5jK7y15Jt1kkfI3rwV1q9AWpUW2DpqXm6MAkTSsW3+vTsCe3MDlbf6r
ncUBdlGY4TkFZfTUyV6fe6x8rpPkgEXxEHnhyx51FekyAIKg4WsYfGEU9ZME
d2E1zPb3LV/GgGPH7M1jy6oNPmHzg/4KK4jwLYlDxuNUbEaTn7TqZlRb2aXj
ZSt/p96FOlm5+3oZtZkF8LieeRwiXKtLiF3ipAjom6KXwlx4A/FBYFnJ+18m
7P3f8Pz3UJ/I1df125MF6K54ESzPpYnb0CB9YgvONPNi9dFRqUuR5wW+gwPT
HeMLIdfjA2hNRNju62F6UiPzSTDW5FCBYA6vnrA5CGFhIpbttrn7KBvFXvZd
N2vf+FQXXegNV+M0I6DKmnJn6fjNn6b9DjB/s9cYz08zqjsEU7yYHZBgBACd
vfhtxmI/nqV3Qd4VaL2oCajpsiSwQJxxT7L3wXdWmO0regPkm1kIhzpm1OqQ
0cQJbSTA7DnTrB7SHx5kmZ0GTexDXfxVscWIcCkP/fkCGEa9brWfNNiDgsBy
ENITqDpDMQDXO8d4XWJ00gjP9IYkqp9x/tIilL2zY3EDKw6Nw2Km2VUzgnah
serhy3GFuxh28xTbSMPzfrFTyrc/UAbZ1cNzBajSRSmMtbgPamdkKspslmIX
y3hb1m5jIkFtBL0D6mOfdzxhP4w9ZpJbrmWg0RFAIS/plPY5df+rT+IACFwK
5V+cR1NfxuvvfvfXlCeT6ODqUdDdg1tpjTfWyt1H9PNpDDV+ZwvOYkFHy3IA
817HMqzrbYiJoMmfmZS5r+I43MVcNCKFTSspTQ+QSgf7ZHPACw5gr0qBvaBx
g9B87cGbfINJxakMmvhmfphlwo+8EuQOBReWx1ysSi4CP3Mw8eIiPhi2ipnL
LmeeQ+uP+fjb+dnUrAI7gBn3kxvM0PP5rYzv8UjMHfE9Vhncic/sgPqVc/j1
kj3UHESpKLqikNt37knp4J0IC+GOxSlS+vCXQtsDMGzui5tYdVQR6zjPivXo
rRS3DPpeoWhnKb3YkZRcx8vCrYidAYk+bxafxN7WnbfC39+xP2WO4vKHSToa
25Km9mAM3aletxLV87cdOISyryy4ryP5FJtQhmhu5wiUbgAFST1ho049wR6E
WvYsUx9+xQynWMVV6yZ4hvMaqOD6cDazKycMlHygzrGeQJq0FFTn1XF80oAA
aSNDNaKssZeKA+w/wqCzHZ4gJ8BGYP2gndK9o0nP13cXyuXxw2ohid+F3U1S
MP6qYBbplM0ppkW3h/soNC1JyrLvdiwqUv1gSQNmIZ/kr67xoBhsCmnfNlVk
Fi6G0903yqa5zL8/VhoDPeCXsRUMrPluaakrIngddRmym16kNOW99B4PN/gV
gv7MuXk/IilmthPnJ4cVE9g5T0IQjoQs6pmDDcRhzzlLbJL0jBLDGKUPDAxX
jt9PcnnGoU0xDhfbzPw/5EG1H6c/81JrO4OtP+8f6N4XrJJ/CoIwhFbkq9wk
xQ4TwzQqKwspDwhiFHFOcpowlXhlloFZEYdB9hsFwhijp7Z/yCYpJGO87mXP
2A3q9U7wN6NU9Kdl5WL6/YGRS8qBbTOYpB6rcVDTjhpF5wYmikpbaY+2zJrE
SGaIFDNQm/jwp6o2lMhSp7zjRVdLLy/pZsvxitovNQaBxwKlEEQP8qeAsCXF
gX8TdpQExuU+rLRc7XgW+cQNW4zQBXmuAGPzDzMaSFtgFxFKwrkckJN8ENh1
wx+F19yGwUqGyWHQJsEMwDrXf2nx+ivO3sr+rIXwh4CufRyB5Zvdj/MMniFJ
6Yhq3wZP/E91FkfdH79EpwDrGT0ByTnSEQYhSSgKSBHGETN5ITQrKYNwqmzk
tFyJmKKEEwwcVQJn1yPRdiCyZGsR7UldbE/uQdmcWNmVbFM8OpgqPezaMtEy
RoQP9XYpJy7ygJQc7ozOlHX31LLJsLF1uDW43f+vmuyRenYt8c1obt3YFyKB
ojvqncuw5pCBYZ4frzH0eOAtx9RUkiOOj3uD0U+tehkljR5K4n71IqUMcy21
X2A0NfIJGlKYHjyQJRfp3F+0ln33bgWGeBU9bMF4v1JpNcDE8XQixXvo2VBT
KispnLuEnuSaX6vgzdUw+ssKrHR3HoYvqEcQWd1vWjhLCVJkCAnlukgsSr42
pAykF4kt1Vw47pP3Sudp9Mc1YpN5cNK1xG0KAxhwbpmOHBUphf9rkDUd2qj3
yTIrsrCXcyfhaxctOijTOwqBKw0rek9NjZfjFnNFBLamuaRe3aRPsVwsbvzV
mOMg1BgEbhk10KYYH5VaGWMFQARJ1KVC6V5mSFfvIAK2Y6owYAcng2g3SX5+
dLzJgI2rh7R4MHO58/vpyRWC+posCUyK3vNiTwmTaUkUC9EepfuLAVuEaeYZ
L3/OuHCuN8u8MQ7aw283r/t8yt4G9R46gOmB5I/B+ItDf4/PMoKTOX5vcZmX
IviPniw0f/2jvSpFwnNlIP19F2pg6yOacBRANZIuw6HN9OO4UuN2HeruZeIR
F7bJZmUUH9GLIiUEyQWu8jAXkVDOFsqvwRZaH9ElMhdzLjHDnopod2avtKPu
EdMs1nY/DoxN/5guUXj0lCE6Gxw0wcaQRvkX7suxV9ChTwkWS8bLv/BHTdFC
R0DgUIKvZN/OoUi7KzNeGnxGJZqD+k6BTXxnv/9fm1zj45QjeETVje9Co/A0
4rqWn5JRgrS+/Ucm/6/IrANAyJ2X5g1H+She5+adw83cSN2z37hkd9Ej5J4O
6dNG6bmPQYUDuQrG8sOCF+2kC9DArrBSfeLO0fs+CygpOSGHUOUqerL7Cde2
4EEmlsdQMp4T1x7eLfwsPai1ho4L/YZw/0jiCsNWgqnWvzBB0sbKJAMk36D9
sucwJGNB8OLr1doZ7ZlqEgV5kf5R7BLK+8/W4ctcUzeENopuE6ssCrUpyLjR
H7+vyumhq8Ib8PJ+HkO9oRPYNmv/h/BOzcf4+rOPTsf1aySSCm5PMkPcLUxE
HQQ/WWVdUpto6PFbeHWsaiCBmW5Q+OGoD1Na0OcPDkeGKVX1CrwH8fT5iCVz
51kBkpT5ZznU1yZRPpMc+5UdNog/IWVuKKEAibSMBKkW3YpYN1AMPxw8u9D7
OXs2QebM3+Sd1VfiZ2DU2BApH3aDhoGKzRb8iGjYLSPnUf3yHIS6qkCZFZlV
8WrOEmOkZx30JVX2JxyizxrUS/nBBVnwuAzprOsZD0FtOQUILY/th0jU8TKp
/K5dYLV3RMV9wjjQKevhZ4bKTFjB18ucOwscfa/HrxiAn3sjI8D1o66lm6S0
WgNeNa9H0r+P/uuOxK93VpWcLkuLukcm06byRxqwQ7JEXx8Kkhamw4WfwV/j
/TOul1Zg2rXW96ajnb1K7ZdYlt4uaUYHvzeAVgRxBBeCdskV96cIGHHMJ94K
PjnIq++cP6YW//wyhSwgkx5cwaww6nHvKrKUpOgzUTdtEHNArQqL0aSvDhmG
pekJkhvUbVE69P7shR8wAoBBldydnGjKbYpDTpctbr7fBc3sHSxYt0Ds27Wb
8TpfWQvVcfLp6R66Apk0TkmRGBFx3Sp8qaq2rQwAAGjPv2z1351JA0VOZGuX
PlTuCYqnWpmya5un5NUnriZVyEfyXuLWTn9R/3fdxuv6PmuMOfBaDAml9En9
9o+/nRai6Aq8NloYjXDCnAlrnXfRfcXU0vvZsxEYsvpno2a5evDnQBjIdRA7
Lo4tAYatjDBrdSQt95qOPfUpvgHZHawyUazY9WRuLO/+OB88Yt4xQq9/0iut
qJ+UusrB9RKBk9Y3cmBBuUmsMXateK3GGwxyVSDrNm6S78nOMc7w1h3H5EGV
mE9fKSRWPG6lfP92E0rWPL9VTTdg4fcZroZIRQNgzPyVGfUUc3t+42qewo37
1WKfUWiox14rgPoutXDDUakb5Qt32vm0Rdt5z4MWSRN52RdYE7z+s3jkUnGQ
Yk6qIQRBZhZVW0GgSNXEZVoYBVx/EaAiJwoP2VnZdFKN7/R+iA2HQ2g1FUqa
08n82ZHg3N8nood5bHVzPf4xxQ1zD53q/7UMu6BUGGuDtwCpwuhEtsuYJRf3
uPl2pEHSC+MLHFV9dlhi3XoKUjXKVGVBowHlZ4SoFSJe4PL8Qnqbm3waRpT9
nHo7eS2Zx5c2KWrgy9XdySEFBf8xxifZJ243iAMmsIcP3LrbPlaBaNHfN5oC
H5UT9PXAIJa9opAdMskutqE4CQr8ItxJOWn09vdQQbwvU1uvc0DoKa97dVhK
gGuQd8sbI8+3nLjhN5f4LEnQsChN2FQgMyfeQYVBXXq50c9tGsQ64laZnZ35
f0FVkPYw78w7WsAoNtfuVdkCUJyNgvbkxx6Rgti9HbmAVVwl94EfLsRVWlva
nHtZWg3THyvJH3x91Z8T1s20vqphwrLEhUSJATsbcJwcOh1gIH3Lv16vGCwP
S2drAiFPbanlP/Q6750lqusO5jj4O6LLzQIi2xwgsDFjEjMBU2rzJR5zAZ2L
kXGmmJuafvRhvIwGk/WegmDZeIXHdWQyq9b0xTBR7JvGmMNb62bwSBpt99YA
O293W3dutUB9+aKfJe6Dw+Vg5R12Eogw8LKLmwRPXcWMHIh+j5y87+cfvK2l
lDxdIWjTUd6QKa0TWOugx63mU5QF5aHfqPKyi57Xv6Xw0ynGoKDsG4ohWuWG
cTWi/aTFw1fIdEdfoCMUt+X6hqOCasc6KEaOUTWUkfY7+XGb/LkZ3rTsRuCD
5tqLlGCHrpETKTzV3zpazdzEWr4vDYSRBsaNejOupwQJWcRZy8z0C8lOsotR
0diwGYw+kCT8BTngfcHp7Bu8sA4WdJDkuqmzE8au5ybu1rBpVxXe8/HKDG5A
TDeb9nLPZUoaa765ZvjtEgejc2Xb/h2dntJw8uqfa73m9IFWG8Q/k1ceGfg7
RUj38IqLFjTMUPKsN7kH6/iwBD7dMAFmy21yohMR9ZpmYZqo5Oq3pGh67g5o
YsClb6Lhx5adfR1WA5DXWnKeoIuf95dtcxLKiW+0z18Gw60CccPvwq21Lcgv
MI+28eOzIZ0/+mQ1Ghkoe5UkYPnXC04OFQwxR9/8HKu+2FJB8verfr/uV9wu
0C4yUKc7I/awjEjwetjK8qQJGTRoq1hE9W7XXcV22FjnZZZx5rJ6zxno43zf
HlIK+c16N11yM6URL46ewOTxAA/4ysK9hUhiKv+H721JiGCnyaymcANlhjcV
rTODfJt7hamYQ011tlviM66uw0D80dZuNjdjdOpzlN5PemOhBxqQoGVDSD8p
U3HVQLPC22/NPwE5IHuTRhuES0G4M4F0tyFiwtbJbBD5HnOSkCx25WC2cLW6
LE3dBZYlQz0wqLxZvt8FZwAScJIKOXr97XLbO35jLCbpo9PAgcApS37Oo10i
bbIYPYO93DOUcbhd0TKTqF9Ud9EWnFfER5Uwd5FQEwe78+MS3/J+Mrb7RKnq
fHL/dCOZmy2dYMBlzFDUtk4H2HMDOBzkHx/DEDGxBNP/rpRyQOtjJFVnxmnU
HOqndhtnLWz8wIjJy+6Y+lPhDM3vboCYpm3uoAeDIe6U4H32SQjfWEGhqhN9
QtpVve/izegC7ch8NeFNE/xsYbTGjnNdrAEdX64LGRk3/cZDI0r5+XOxgmfK
ZnPCjw0KkBAKtWzDmn7CVUyGdVdv/nhBTq5e583xCERpwdgz+llcZUFg6ZVU
7eca6w8/woV/YlXkLgOcgdpPDfWLN2wyEOT0aTXbLVimix8xgnIwms98BX3E
ilZRjwNlZ+q2y3wByIWzPhrvrmcOGYan/8NssVWbOJ1prfuk04RveCi3Fn+k
wACWPmlLlHxgL3a4VvmzbTMyVxfWpKRsfKaLjXiIBfDVIy/6diI5ISPm4AQF
T7x9jsowll0f5u3kPY9NkL/J3SdVdIf3eSGZEvNumH4gusua2tyUhH/1S13E
gc0a2Tw7A7+I+tZM69ifzZUXGQo9UAXIIU1vBl0185ZoosU925toSn3jB/it
O7NUlFZxl3KkfwVuYaw7qMDVN5vEnvmVAcBvxDsPtyZRAGVdHz8NPI2nIfH8
y3znkzLsxb3TqMioqkBnRgms7JPTPhgeb5tZzvnOxivf8uWAlb99jCWgEy1B
2gx8OeoGmtEse77l+HrLZ9s5ZJqWW+omFOVkrKUABVcmkkdSxTTKIzFSe3zk
PfN4xjplHQPGhdIcVoDIrI0pPZthHvUWlUBxfYHPMCTCQLXGScKYHe4iHOWN
4NZ15trVVKBp0ogRW0lHbKAc6If3Zc7iMILBRDgFzfgSCO2ynJaRXQfGFAWb
5cT8GbV1RcJEOSDeU9zsfWMXnvck9T51DO5gFvcF53pUgI7K3KyiRgDS/9I7
ftfpduOfXeDxKsNxi0OknIUEggWZPFs4EZAuHCDwyA30WDNZET97iZCipIo4
irbM5U0+rlG/1pUbHQCeYD+8SpbnOJlTxXaUvXMc06wH79ExFfr0a2hJZmdy
UV4Aj0h77Yto4DgmM8jnJZsZSpKIJf93mMXeSv8DVWq6bBzsXkGyV59NCtnm
ITqhOIWQjbHCHxW25c5MteLxVOxp6jGGrtCzh6R/MYjFaD881jG9APcOYnVM
lM/H4qzW6Nhq3qPzaFO7JpJvMtwpa8sgZ5U+aigl6lKsZ+jrbS3fi7+OiyQt
SE5W3ZmIkRY/PLJQWH2qQBKHppERq/u1Up6oBXyhsaX5cKs0D3eRbjXRDeXY
OCRvIghnOT4ixpUjdngYgJMhg0bFN/FE/HfumddcCo3VP/09391bgmoUL2Mv
PJgEAuUX07OzKuAoKsbRlLx3isexMPkRBNVfIu6V76nOe0cyz8XF+CDn0gKq
YC4TeuL6q6ZmkDaH1KtnQhWIqoHwxf1bE+/j9lwe9KiZngMPHG2Cv4P6oE05
K6FkmN663DFe0fMLqDmet98iKNoTLIgoLtbhl2O3jBVo5M5nUyjPO5BCpuP5
p2/orvHGfaakpZ4F7vj1vGLKTsY8Ir2V7JnQuIF8ngRtjoMhwU2gP7FQTa0g
t6PHrMVjqqjlQSLqWrWPXVIHnRiolzRF3acOrLHwc4xHmg58ekBeiH3R6nm1
6jkNIvFx1RdkNtnbfV7qZrxCLYSpMc58bylBKkUg97/qWLcCGQNN+mq2Kdqa
PjtV7iUOMftCjaNYA5KJMq0fPceEsgb/2IywvImLNpwe4UyBxJeWFdF0ohw6
qt5DZ/Cg/uwQX6bkVQtBga112b068LE9pglqE4NUNviAaP0aChprYrhhAJ8r
8x4B35BLzRZfHrXmzZDdDiKr1jbUVPUyMs0VLubdWNUBRZtZCPt8+V3r3r8q
OYtfe60ScT4ljzOt+4egbUQ+7HEUePPgTOfruoFTnb1SktwEelV+Xm8Uapme
IRvtfTFE5yDwqu/lKEHgutMN4iW2O87rjVxKbU8AsfVqev+jD4oy2DlT9wga
aU9j5UsEa+5kCIzvFvQuhTuOWGWu77kb2huySl73am1T6dW6uQfOtcorsSqj
mNb+KItnBesuKUD9DoC8Atn6Fp4qCigxCt47Jnwf5JBC/88dX2EvtnLobc99
B+E4P7QUOs+SW9dB72MAiRj9pCB7KyBOTVpg3mtXLZxeY/xKvGJK3dT2cBzN
JF4UpbC+dOpM2QEO3YGDzFO4ZkjeTuOxSuOzIhitPYW2akAUrnWTZpI1orzA
QY/McXmvDKe+oNkqWk4y1xvxHDTj0t1U5r7kGvu4lrg1AId/clfJod8ojxer
9by+WTXOa64hlZ26VdhayPFbvvzoZunsE2cLAZDFtwWCPyUYui1ugEZY18PZ
79Yhr68bp4PuxRR0tUd6dqr9v17RdazFM3lR6SMAypt9Vqt6rzXTluSQCw8u
eaUHA0x6aJlZon7i3LX4Xb+QRwYsUP/YlbB/SF+heuQW3iUzD4kWBCEABOuk
QhawkTRtNpPxNUbB46eq+17/EAQ83VaRJZx925+03M6X8atJ4yF9oBogYQbE
vBYs0Z2ozboBIKOPJ0/pA/D3kZ2BXuWfWqDhZGrMR8KD53qwRGvZMozmbIOc
ioF6s2WdCc4MzCWkX3RBok8jE7k2e0NWIWFzxki3m3ZWDwoJfL/PsCusshz6
YQZUAfzcBVoP0qNP1s/ybRmcGwAEStagcEDE+1X35nc5OvrwOPy1sYV26ybJ
OLfHi+vDXsFVrGyclqWY7Po4cQQiYDPoTzSejnOXKxUApxMLHHYEuo/S1yJp
Namh9emFKUgvyzqhPfbwkK2TgfAoBGMjcI+S2pAovrSbsHJzYahhQg5dhGKp
hrIYGjyjPBNuahM5HQ6FXArFNBQY8FrRS5FRnsij631/UDdM9B/7XSdoqSKJ
+uN8yALF4f15jmwE+3WCks6CfLDPglEb0cWIc85OmkQadbPcjefnc8DR+h3P
Y5ZmFxUFRiRo53x0Qotuh+1ny0lLqD71oxTrunm+weCv39NhMQaA0KB+tDZs
t1clLS98MtYbKZFqzmttWRkpl+93f+3Si0j1eMf2sKc3NSeaicZ/Ka4kqgtw
3RNwxWLT8BdwQQPMzUUvEgYIq9z9U2DidvrSKZmeM2lxJKHl0SxXNluM89me
vddSjue3yo3FZqQ5pbmomEUaU5ZXIA4MsJe+aXUxVXKlft3+fwzGXEVtrPwf
fzKWR1YRJfGx0oEw/rLeFxnEMKmUbU8iUtuX8HwFEuKCSOV+DXh2wolB0xZy
QNVeSbZpzE9ZD97cTzfBGI3LUFtP/8rKvpJaMAlQF5y1EcorzBYnKojmuVZ5
pQyjgen1f93Db7OSAUIhsmmWE/XHK8UCV3xG/T68xDG0mEoDK6P/6nyF1TRK
9F0UM1p8bO/vTNwsCEGt9g3MESB8ZMfm98Oy3Hq/7hTGk/q3O8LpiFf+kwK7
5AtOkhMC1Q3/PITUykEqMgQkeZMr3HxuH2Tb99vQB+VqjYO5AAkMVwUW7hTp
oYKbxQRIa+8vlvo6Bz1YDMI2DrbM7vi42RUfsi85WKSpi/Fr964HbdkfuHQs
cgEAw1FryxonuNCysoevUbp661o4UodnY0EkpiOxHVEoyTgCx9p5nzy3okoI
qo6XbWpqzZQyrUCqOfOB/rgvfQ8ASzlH4cnEO1KiGgJ3tdH4fPaH2sQ1h75W
HCKE8346fcahcQAf3Zbj5VDSNCBxd+TWzOAZLfeXRb6alnrqiJM6TQiTelhP
v2/mkzMGsmZfjxOpqookoO4zpWp8o+1GA7bS8MZXS+fXtXhbZLpVRnDa95fu
H+DwyKsTqeBxJH/wZYWyKwVzPNj2r0vYmSMZb/T+VS5EuIoHPBQua0DSNxr9
kT8YeAD6kBPq+4wwLf9w/aXUrTUDCcZRyvBMBtkw+bbhyrWai+vafrxxbVVl
Hdia2Lm/3TBsRxDwwFBEwARoovcOw9JJdCNWOzDjIDYP5YXmZcO8Mp9WAg7o
iyhUQxtRKN9gCzBK6X0tSDu36+0spMkT4LVyVQAnlAPNVOh2Oug4KuDho8zQ
uFuI+KuIbpfoCWmnagbBLs2i0+09VRk7jeapVKBnSuTlanGkvvwaBYs3ZycP
ny9wbKfAjvW24w6vg8GZQEIwtsavjIzDDem/Y8TdK83zX+WliHRTAp8D005s
djVEIXR+Dcw2sy2/05JiVnT0Cwc7LFIWOGgfeUhjDvfmZCPJIApc+zBorkhp
bcmixqyDSrCDGpvp4eMfplB0df5zQSG5qPERaKAfU0BQQaoeWGk11+eeDncX
oTBk7O5cDtIuiQBFmIm4UXBZwi9OEYyQuxigTrMK83cooYalCl6MqlLG+H1x
4LnYTp7CA26l6bqFZSQ0ItI/vIJ5JpNygyNv94zuLhQ10/C3u+AnuDqBKYaN
PMsHv6Bd0UQsWh9BXcbhpudd6+ajTglnh9LnBiKH5DOojZZ/6/aIonqDhTqP
xmFJuRnBqt9JGcp7N3CBqCyVcDJ9YP3nh561VJW8PZWFKGxu5tftj6KgJkfK
1Qmzpmz8LK6JeasGko77s8j3H/xlNPwWkAMyn6wO+Ho1OgxrBIBiGAlMfoqN
6ICa8D0Yd8y4dYXIhP1FAshHXStmXC0VBOEmGQnUy63wUhBB+IikMvg4WVsg
9pxRhMioKemIeEznTC7VlVeUpRf210CJIk0UElJtDhOByTPdLyNTR20x+xzF
c74/Vh3wUpq5qTZRgyXy+DdTwJkRumQEtFYzDr0Xw1bs6m9Ye9QpACo71Gbe
rZS75ebOl9ecTG6NezfcbZ5g6+efbBIPzekAqKrFRWEh64+rZspOd+ebQjG+
yw7Y0aJRn/PqtXikBKtoeDpiN+ZkaUFA1WiVOjp9Y6MkD3Nt/csLiZbdiixO
KlfjqoY9u1FPjhjUYduAxVnZl20Ed9VehO5t2FXkKGiAaG+59iEylkUC9/CR
mmGcE87FLjeX/q/BxhJ/wkkA04FI8fI6HQCSVQFfj6nZuPKtLRb2E99EGEVU
H0xsuDzRQki60mjgyUkv4bdmQo7nX/XJ4K7eeA1CcCow4aCWxCW3zhmJJSIq
tbdeVj2OIKGswIyRUHOHsUPRJqK8QQw0sNDQ6GUpeCNwYIS9MP2Uti9Yho4t
/KZf6B4Cvf3TW8w5SZnu2Yixi2kA+zL4riDB3pcrkZaywKYCkXAVsRXzxUR0
o3py2CIOb27NLbfD/FLNcsVDVeQFxZdrTULL79j2PQmMk9rz37eOwR2takXh
IU+uz3G1Bx/cDQT0QglqDqWjViZFWKpWpAK+IhH/pLCI2B5zqb2X3Jeiq0DF
BPv6E6GRSF8XeNBjM14RdmsUmTdjcQquvsRp6Jy+BstfX4EoWF7XK8giB5Ze
7+ce+vUuu7Si9+/Bd/hYonFIsg/P+FsW2UPOJ/bmroUU7uCp7T9bteTRvTSQ
zzvh8iNVBlf7vptv+tC+UkA/LeV5ahFw/0Asfm0QVOQQB0pnzEXEZZuoaVMP
tL+wb7Mp+uijLwKbzBagUi58sYLmrPJC6AMRP2aABLLuA4es+7FTC5CesHhv
3kJ8HlJpbfLX60SySJJKZcJpexOn2qlQke1YSOJ8WGfUbo/jxvIPhPnJDpXW
/K2zZkqBTpvN98W5SPWASC6o6bocoxkE3iyH0hXhGCZXuRcyADmDBasnYJJh
qjBQOZ6nSTV7VZQ2z+X0Kf1/TpspssiFSYVLjtNCShtg+douqiAPTvGyVzro
zhe6A+FrDNe+9a46VmFjAx2TTktkjGhIZk3dyhXooZZpE5bMBIBaXcBHNIZr
QEHNCIGoKXiVU6D8qBUBZ3e6sMxdOmbK1ilt1CIrtiN+6ceu7PyfbXo6NrMa
R/CSMBkyL2XGc/kkQ0KZObhxf+5ZswXoThQA1SxTxNLGda3ynAaVChwpYQVD
U2Am2OE1PqoStHbgqaLmamY8rsaG5N7DMSNqfXR+OVmONfjDW2nqhET5A+gD
vRcN3qiPJHEJ4a+hzalX/sZuBQCjg4xsWIHQpeym0jLdL8Dvc4/AYHqI95Aw
8iJrzMxfYWtXs9nduyr7l/HYTlZ0PCrlK+uYv0gg28rBCdiX8Z+jwl93n4lE
il0ZCiMjHLkODKx7DdergQkzdsuAiwl17C3BYkwNQjp1zHufFcbCwS2wTP89
4woUEUQ1x27rxyUdtCq4UmY7FB3RH1ad39fKCmdPGsr7UMITf5xsYNQ+nMlM
rwiQNC4OWjO3CkaC1qGCWnfqbCb8h22VlgRrBZEngCqoNht+uczqwgd7HSjz
rHAcRM5U1Ume0uMCCKl4MButo2sffru+vttCsIQUivrtD0cTFjrfQ+m8kEii
ugOTDYQoAzJVTp/hwc9gU2eNOt5NmtQSo/6zltpOB13TOhX/WQK4o76yIykJ
IH7gZ3ZLiG4Ke9p9HHAjjfVtg1yL/9PCrLIKbZYE66mvvL5KN1IIsjWTRZmY
dR9RnjJ/qlWUoPkITRGYWAxyEhDozsEz25buzIFpPpDGzK7C4NrWQDLFWOux
Z4BkpqWlYM5B+TOj9NhY9mHWtZ1V70zGsZB5ea/hR9Y1ZXYzggXrCYTDcGy4
9vHKvXWXmPxJpqOs0AOSMWqaDMbHfgyQYBPS66kA3oSJIOEKl/VjV3etNgQi
5lS5Q6ROiPHQcecli/TXmbm4yK0Ep3eXdnPsOK2RcayHK+34PT2AfoItKpna
MWgNAf21P1KvbKHsEcV0wO52ZBuA9ORxnBsumvXdqrmJ9TT3z/reHHVxAj4F
cHKuoEqvIIPTcpQ5vLRV7hNlPE9nIQXNRKN3U2v4+2nlaMFK38QEYRYg81Rh
AK1zuZa62qJtWfXU+xFLLN0y22lX05akp3IB2OLZkPqYArG8qVt90iJnGdkP
FGl3rWq+buhimqzZt8T8fMxGOw5QuM26go3soYvpF2YWlc42KHi7P1JBtez2
hE14+W20tIHdeZxF0XlHANH14fCKDWGZrx0uMZDvp8xcpbjwOfbzjM4GLz0W
E4ke0wgDIeNwH0gOxplUx4hB9X/+JNald8wvIRMrDOQOY5g33tr/mky+6icy
g8ANQ/ZEPjZl5UrQFe6dVoMpbpLUNQlHWa4yd0/X+GAo2zObtv9trvcBoN7L
jU1sYjfitn+jNXj2DIbveMbFh66lG0PfOWWev/sE6OcWherVbWdDFcmvOsok
cwM47q9M5pdMRCf382KIgL+RbI8lK5Bdvwgn+T4ieDYtMHOk2dGZ6J/e8w8q
xvgVbZg/qdEOZqrnD0O7zR90OWlkZVBpuQk2oMq7W/Yb1Gq18byxc2PDwdPp
bxXKdowEi3BiQLdHMAzMycZ6tTtouTiE0zze4TuZogxBZCPUdNQ6Ph7d6for
254imz44gCvL6CBxB12ttPvVS9N3aZAmjPLgpmlXWAF1AZiHnNt8Hwd2yBbr
/arwbcpXc9eorShQced5n0ALs8VLcHtBBEVe7rzZlxsunirGYEmROeCbAS5T
zAGr3hUc6o5MEcfe6k1/xjXWnF0ojSoCnWuqN4out4tEDeXT6Po1t9lIRYGR
9ykTDRCYNmJF4j854+9K6SJDDOh9xfzpNBGPgoht0RmDHvwIyuZq54XhzC19
dTgY8knyp8G7E+4mJOb0Bpfwk5HfmwRoUyiVRtNzos4G4bJKI+gcG3DuFgrE
FWzY8oM6dKx5PoBMQbEETYU9QkcZs2fnRNPn3PXu9yUeemkl4s4XpIjCUF2w
zCSImDxWe0oJppcG94ubCEQe6ZNw2zLIQ5NEwbn/mZOTo/DdgE9PZxSP3RvD
bW9nlSuVVuc6H123aLyr2ooB55NrMJHlpkMGnTTGVoFx+jDvS4nthaYLs0Sh
R3469jXSSSvHZMhkqlGUtOIzyST2SYXj2Fl0m8dY7Fm3AViJRE9v7xT5WM6I
eQ6DIXXQnsfRW7umBNVkpOmaUKlehZPuuNWjbe1IDQFVaXT1ILlJS0YPRCps
3wanpSFWTucLDRm+j6ICRpjLXlhofrkqcsn8Axte0nQq4ifvaJCfzYIS55oF
UAH4UFXpQrq4SsaZxdfjLDWS40r4sAbjnTUE34UJATYimXbkffzOKw1+Dfp8
9bcGzpKROGnTJjOH86X2iIRmi5euGHfieiC/tjqR8WgBsSswhTABTuBRTISI
r+TyimUQU6A5S/Z3tkJAz6v3DApDZDpgedVKCiyJlf2lIyAGrxkDAAlVJywz
RbFRDMEBiAdfRzgAi8LIeGM+uotDxoqmfs1Hz0b7Oe9UrbDhbxlp/NmOE0I+
Jp+d6jXFPobxLl9SMT4/D9Mwk9Qe/53YlQTW7RGP3fCrF5tDnIvPsGBrBibT
z/x+qbd8+Bz4O1ckvCKHLhTwd9WrPdniUb4GcY5GsGwxWSPyqAiu1yqagIwl
EaF6R/Be5NKqtRzqLvwRaBAqGTJc3QSUeBbu5wpE17RTnbYSHuwNmbvasPr/
PZHV4AReh7pc/gjmy2jbZCXWaa1hMNZtXelBk9+4Qlil9o8WgVwgeYXYdgPl
XONaoTUdtfnjqsCr3zRP67Qc0Ld6C+y1fsym4f3CSE7foAWxOPgQmnJscLAU
KuJGwRCKddJElW4ZLf+dZtKbooewtPwoVRg9VqVsK97T4NI/qlE9CP7Smjw8
FuVRIxWpDQLol7Zy9kEm8ewOZMMnsAjAMYENiah+uy3LVJcZEErrqyRgTwWA
a/6CTOOrErZxN14prgJL4b2amUWJr4s4nuOg5mR3lQz/mu4qmPOSAn5TiNBL
uZzZhK8SAsvdxSq8KE5zX2nHmru2Nvz6OFFnAeL36YNw4nkPHBvgFsfpGNGM
f6EiFGsfJQpWmQhBFrEFdUtICF6Whfz26hSujuCa9hEjK9WcZW+6pn+15tac
cisMYIQRw5Cq0Mj7p3aMSF35z+T5q3a8NdD2rrvqCxyjMo1p8W3hJyM0NbbF
CIp+zBlwutl8vGWxvQJCa01oaEv+Pwi90ne0fg+EuGhycdsAcC2wx77aRo4y
iwB8UtpDWeUqidUlQH+dg7rbl201czzICcDFZX7Ch92EgGswNW0C4HKDkU7i
q4cnl76g1h5JD/Fsx2iMPss/2SI1SxdfugAhuzDK5J/XA5snoSgvxzZury2s
gfe07FoqXSEr7jqKsjDllrsxUOyN9ylX/xHZajJXFXxCaG5YXVNK7Jx14xcJ
qEqoSjGX01CkNhN8AP/q8gwMUGQ/+uNQNI81JY/IzNCRy927JODhtCyeECK1
LV2aW3bBe7mJxBJ7R9mVJg+hnKEbICaZX0sxET+m9MrbjcoQcXl1DDXp2cKV
upjqPH2O7VPtiUfJnATPzrGOzqAInO1DC35B4EK7XhHY4HggBhSFgJrXhJ/S
/b7munSk3dPwqCfj/1X+UybC04bsCWKxnIsgv3wgaIicKzjePSRka5bhfQhY
DQzfXi4AyiXd0B4ilEungZ91XLuktIFvgX7WnUIKTjE+2z6BTxk2vqTP2VtY
j6MK8UzqrF3qjbRgrb+/9KUBeGH4BNgUjASXUrW3aupMYqwp/lm5uFtPNt0A
WTXhFDXZ7rDf1lwlff5QIXvIbXsqVeWuPhemp7YtKNtbjRrPnsr4t8f8oPTy
N2VSbwsV2k/e0ruB1JPT2WgkQCNB1sX+03I+eLDODutC9wQADiXpjgXwHTMo
A8uEqmOWnuxolrtkR8XluZzCD9CWmKzEXcvs5isYqbQ/4Nz87sbTaVwMUSVe
0RK9fCn+1oyyJJoskTWTNZBKcsSjsYadexz3J7+tuEbEsgGyLh7yS7vsxV+k
qnVY5kOejYXZOGfBcpECyN7Bl5MKpOnQf758t+DnUd0LAdn5geZtyfFncCG+
/iWEA5vhnf98RpcssbhcHDI29qPp4dXleDFEcmueYzqNQQOoI32e2OpnQNDq
aLxAKlrNPHSgntbDL8SwA5sDpLCXKabug7Bvd5p/JqrtckyICLZyGrs4CkA+
zrsDVziB9xwIL1JylmgCYl5B14GvKAqRYVXUj3Wvjn85gEf8xA+byKT87PiF
Dik8XBGrNBjyIrg2YWQVBbvg5JGjX3zo2Qw9cgOSH92t57wfqFYn0hwkFGli
I2b+kZ8sCPzUGCydOohY9Jr7reXeSU1IX58Z0nFil6ZixLPWnEwyKr/COCgX
DuulI8vJTjXG2/i2vBEAlWQIJqIgOzDkwmpvowOZfNIkIkd5JmItE3Vu7VP5
B5PTQsCxJMaNBvhizgzZBCtl/CcckVdt+/6d4k8pXD6hABqgNM1+atIEqdLN
HU2qmk6aA5HagVmdzx1Lvv45V47H/hQDukPce9U2xoh96WHcLrD4nwEECpL/
Z/w2WfoL5ZvpVwazwa/0pO4SZkgdwafEIWPTggnwadZHgKUi7aAZe7GZHKIC
xVvw+6n2m4EOrtDd6bVG/uiLq9e9q6/RHGQKEAOebY1m+zjrGOHYqtbRDtOh
BWosTo3rXoca4JFzwTcCs/LbK0SYu9dDbcKs37dtlor8/mDoyn9vH6lVzEN+
AuG89mKdTxUXVT4gGug6ofr94UJY0PK8JdcFUn0JZiQX8bktDd3AuKMYKf7M
/n+3+zjxQpWGAAwnIZp4q0nPTxJ6KiZqPSLcUtwCADh5rJ+cNCVfklpKiW2e
WiIg+d2c5NciKnr4uslrHFMM8ma3FmWKgMOk2Y4OJ0zPwwnxVKo0wtIzRSIq
DfSNJaN76lK526cfIQ4JoTmevhkK7tYp897MTgtYUA94bSmsl4RqM3tpXnv2
5N+P+tvUDridOb1JxsFOtgDUVdNcE+JUtDzK4Ls6fqZXTwdTF7AHr34u1Lfl
HWWBRYJ8xfr+RiSHnX4r5YMNuGXivH74O+TJCrA2hW/2koTFoqL5FO99Rx08
Lg//W9UqHSniZHvi0Mrid2+eyWkV+1v24eJtdww6/aPkmrCH/gEixJpFZJH7
7Ok/A6hxGZfd7WyuzVc/BWZxJkuhY4fhM/akh3Kyl8H6Ea3PL7ghSIX3chaY
FT0z55Jwe2itJkJKbXHJOwP31vCMz6uM8gGZx+2ZsPE2zRnGx2uNRg2qMN9f
8yNRahoyf8UtxboGY0EkjVe12yBuHgfH6zIWk2Q6evbDhPkugsK5R9Cd+HF3
SfpSVG0LxkmSuMvFSgQ9Ovv2ixZ/S7RWYg9/oQLx8X9375vM5e7gMNQDWm6h
WcMPJc5nLgn7vNRYvOzO0vrnIXgGddLrXJpCq8LAcMp5FOUDN7oOD+UbFtxl
GhKT8+/8li4q9EtvIy0S+k5jMAH5dwlIYBy6ATRmjWBLq4zTAyxru6nZl7Z7
MjTy4FJrY1CY6Ovtxv4cdaK8UUIKVAgCuvEwCgbBoJl8RnqXc4SoEGRYDC+P
orOP+UFqg+vsw8khpGVDZNUZOVwQMNMSwbSYmZcK5/ec0sdAUunj2+g3r7YS
NEpo9NGzeTsarZhG4ifYEMrlBXsivJXwimFULQtuQ1S5kjBULR62BdnqOknQ
pCVza+usmgn3RZMHYIfZA+egcPrjUMgcOA1QSkSo1m7Z+x1YNEyD0zhnAjQK
ms1fXEbwXkyUt9saGgmlDNbXRs93Yr36kqi1cHR5duTkX/AOZziAfZrk1hes
0fhcCvuBkJr7hbYhDTmCSuv/iHrWqE/KeytcGZQRVE2gBmYI3zBc38y7xyQi
/7I54B5zUMCfnuZr1FbS1DrttUykl9rcuDzgcfn5zSpqf5XTeclC1VuToho9
3+YCzG2zwO+S8U7wGE6BVeHD18pWIE5+EQ5SdwqAOZbPMilhQH7ERrT8XY83
u0aVGPUcHKNo0gelcadVS8U3Rf2eKfyG/nranVL1Jh+89q0Wlxl++EenZj/y
9HnPfoy3yEAVMGX/yTgiQemJh0TDZfNvHNpcQOzPPd3Ht4mEaUiBgVjajR1N
0Ej6SJmZeJM/6APtwOecALe6sNiv2Od38G8LvrtWPjXYhIvtUOwlFpHHGPCA
JgtAhLfxQ/vWeIJBSybv+ZC7tw136jQUfEe7p+vnf86h3W5C3JmEVwz63CkY
1VgMNMGhParIKKpL9WbEoDfZzEMYBrE9j1CoLYfaj5Pmk/eVq8UAtL6GZ4y/
n/TkyYlI63e+wurIWRlqxLeA/zIc1BOAjWkVo8RYIKeOtPeM+PQdiJuGMaYe
u8EtV2vGfeYTIhYRei6zI+VNI2vaymmYwH4JHFUhx3Z1oIA3Icqrury0+AbZ
KG/W3wCLPFVkOslS9gin4bZc7/UcDTV62OF1yQzXePJhT3TJ6uscsvUfZ36M
lIcSGyVPKrsaYK30HcpqrIQ66RH737V1WDGKIFMhdlFEY24JDhKiKAzEFDBd
BS8kr4tosR42sSktfi99set1K2agqe+YRB8qNRGXoxSl++1arJkFhYlM6ACg
tMZftuZemXYDO0dSZDB9rue05eGH+Sjn5Mnc89IMwbMYSZb3GdKoc0RdKjh+
PvKRMbPn7k76OYSHeWpp4y/EYtUyZl6Mtq6ErVUFVeBspozDSY5QLpPfgkmT
5zf7kgkqKifB5ryJ/lVM0S+bimsuXwHrgyqbijivSqSYPWPBUdnaP534kQSA
4OjtxJJMwGJICsEMz8HF2LOvpQyATLbt+G5tJDQl+ch7H47gmowUoMB6pEoB
OBoVsan11tPuok/abydgbX+39fgmRmpcAVZu4Q3B8i2mHegCyQpLIu5sEXGP
qJk1Gk3hRuqeuJVDAittBNNatTaj4kxHQWZWMfpw9nMky/5kAW3n2cVW33a6
35vx5umFsRqydJECtG46xqQOxXzV7MEdt3kBDYx02Ye4o25edfzM/NjGrWWe
IjEoBAlfUXPIfc3I5CWW2C5/4acc3SObO/rJ4Vl93wlsBWFt6QHEBc2JSpv0
PNdcYfBF1m/e6TawkESvUuBC4TIM2Eh0T+qOJTrNUZQ+zw5Gs07riHYkCuVk
sEDh01xiDZaloxxUkZ5dbLLZ0+hCNvGLMmFhZPzMRDnhc9xV83AJhNhjyqE2
QLAkqL7KnuztXG/HyhKQRvdfEsy0D6KuewPCKshXyUKKDXHWZ7zz+is0qw5Y
FYe+Q78JPnnZBRqAmUd03KTbSrODdGPRr5bXfrum+F+qwvtw/OF/EVGxuhBp
15GL3V3zwnnh4YZMyLOD3qvT2G6jmKOTOQleMdtc5/NS9pdeVILrJ3c/zGA/
82FAVcEq0PAWEmVNhO3Y/PUAxTIHvthW7wRQDAej6H/gIAH4AjE4Pziwl68J
xl0uyt89SqW6egdUpMc9e92cLLH0AdCWDttAmg9wa1Y+GDHyxAen1ucpHgTz
GLg7SXJ8PtUIVgum/IwaEfkHvi49UbItJhpZwDL5KSs/FtinR0vUE0P7dibL
600dGvR2aMbkfWsys8TfOyLBVrhxlwHWdTOnZS2MOHYuc0+qGeAcxoInJQSk
qwFM0bkETv1ZnAM6ZuFtLGPCzgX+1LlTdQ3xrBpDyL4p5rw1UQqgysnY7XfX
rtBqm8akOrF8qHOtoPwEQCHNxBKV34FWkjT2ql6WN5sydwFv704lTDwYPom/
Zi2hpHCUj03Jd16KCFPFXLIPfwOp478qGXVzMAAhOHogNHCru4w58LDlxh3n
/5FLLrLS0bY7DZCiavQ22bLaG6kzx7yVi6mpv6/JzOdtRQTf0z0d2S1lbL0M
sHVTdwXwqfnK9pnxTB6xfqIxZnVnrtt+dWKPShEbD+f/blz4FPpu7NXGom1K
SDjVpAAVFiIR2VWlstQ+gOoF9g+X1YeVFduc2B9bELbAsCrpaJauzuQq7Hjb
+wM/IEmz0gphGyw53eLygfZy6hnFy1ebcJIbbEZgBc/ylBrQC8ULwGp1MW6O
d0QOtvAb/EOgXPDt52BCzRrQU6Ph9gEevy/IusMpZRCNDyE2Cw3LlHBGrPYj
yW93fCKxnyovHPCmtgifoHgvpSA8ZSoNXKrQJ1v/4thKaqJgT5p59y0zoh4l
73A27tZ7c04JQZP1TbOQUC+Tl/6z28Py7TY6WNOk8vDCXzBXokeldygy4+SI
9/hj6P3J3IeEfmYuyS1qGh0zVykkG0AG39Cd9u0aHVapE2MxgUMjqUbixF4j
G89kXcedjKu+swYEl4uxSjCr5i81O+b+o8PFsDXP52AKz2DMnDk62T0JWzA8
Pm++Fj5Pd0RzqRK1HApBU4j57sQ+G8R3knZ2XWx23vKbwJkloDlLVhWRiqq1
WpJne2sNqRyzt3BfUL6P2wtaGe3PL1UjsoTpPi7lCj5x0wBVvIrUeqPmD6NB
jqwu8ei84v6CXfSSlJF+Ys5ZnS+MwLJucCAamy66UUWb56bFmCzbwxtdEnyv
JxmfOuhqt6Kx41f4nVB/aGYXKZYDpsQGI5QaiaNsgYh6zUFmCBbFK5jPNdUl
2A4U+9zmQIIT+Ngagar1+Gh4/9e0wjxVWiZ/dj/XfG1pNeK1d9sSuQ95MKb8
5XnXShunWmw2QvFt1eSf/RUXhBobLnFy+3r9GjKl4XRRpUgNMaKGJdh9uPCk
a9UgpuBT70nQM5fuIUDezlHrtmbu85d5i94+miDKwXTpySoQJt37eApKAvCQ
LzHnowETFeH6++580bfEwjOs2ArCKG3yZ+TwMgVMWWOfDXfYrZK3j8T0r0FL
1cQV2cF5d9ZQ5bG2hA7nH0keMWIIXbMdrofc5b4FgaF3RQcQV0DClZ/MmrPs
wdTKL9cqU72ZvZaFyvnXX0t3M3jA/ZxpfodB2MHLDFSvTBmagtD1AY8cGnGg
gacvkahmyu7nZi9w1xqHrpQl0QyhfSN3DMnczKKzZ0jmdTNCOkLKDLcv1guj
DGL9739Im+ZMYMEHhoz4wIxFTlz2OY93tt3At3FOT73/tzWK4XlFMANwl6Bo
/uVE+TLt7E916co3bm2A6I0ftNBMTgITsEQcZwJFwog/UXfAEa35LrafRcSK
HqpS/RKHYFGozpRkv/yAvO2Y7aacNBcV+iq8XqHGpMOnNq6/orX5zMKNI/xg
+/K4aODcXcM6eQW92dZwINR3iEQ+jmzVhfRc1UPI/cB6U8RUqGmg1MB/jFjU
1MtuSjAAJohNDGqGPz4qFoqXZBh7TKUSaYHa6cnW2YfmLY41kBdSp/x/Or3a
dgeQhIKMPace5Lw5UuKZ7mdve/U2qFO9IZRt/lw39N3GXZrXqPMIfoXZlzI9
8DVRcM3u7n0VsyAVTwIPXe9JpfWJ4Vo791pJle+2vzSYKoxlHA49BgX66d4p
7Qrcmqw5+pq8gxO/rviVrwaV6jjr7UOco6G2TZsyCKr+M3XaBIwKQbseUZMZ
Hu65oysn+6polrBZEQ0nld1oFqODrwNUL1aIPWc8zhYP+n1A53187QK2Ng+a
UNXYpoF9uvFjCFaMirtdsG1cWQA4mwg6CwyV7uA2dSq9011kaTqpCCmSNrbX
0BMcRBsP7S5Lfn9ghU+d8BN8KiVjGnlUq74+4qzbQ2a7lYx+Gc3TebXdZtbX
GS3IeMHG+uEuDkigugBuCz4x2ix3XGJ8c5jxXY5CkACV93iETvVqFkDanLtl
sdoxupKZwqHd81Vf/7WRuWEYvrEl0gedsIXw5pkyed9f9epo8NF067s0oY3T
821HL+FrigyO9yY9geliFSxMqESd1L32W1IMVdlC5aYHIEc7torNmJS/PUJv
rhudqGyykddfAsXUoM4fd9/GIWBTkPZzfWo2BgqrJXxIvZ6rJGWOqNxBEsKs
LLxb3KLIpr7M7+MknkwT8PzaxyS1o6T4uIeTXIdIqK6s86RIurfJsJ0m4M+o
ZWvrVCZBjNUcCEim3VL0cv4UKtNxmScIklyxB+Tdycgoi5t4gTso8RDG4k1Z
lnId1Hs9erq+T0uYdmx5WbrbaQztpgzHO0KFpKAUblbAVcLrGYUULNkQmMeH
zFOwrcIRTjadI2ghADpMkGX566jjysoX3NJciZau3F51Czpr6eoDVVJGjMKm
Nf8AjReT8JLpWw607TksUZ1hcILbj/s/+tncqmdLdj1RL9c1PgBVdHBpACN3
ToGitBPOH4QvyRqgav/FQGRN/w0J2iGVujnRgJxjSpZLCjLJho7WflNnXq4H
iI+ohpgsh8YU8m1jOUJTfp194ILjx55MgJGAojiA2WfeXIKqReGXiuYjusBN
7jXo3vtMpvfaFvO7n/cGAoRlpuqOK2SYNJOYVJ1ZBgHdy/stnoeV6ACZQekj
nUrAM7q3/8cwEPb6Tia1GOh+tHI3xyHnrohtcwA1cRvGk4ggNVNfth0R7vqB
m0qA8vwZA28lknb4x2oLxw5ajIGT2me8J/ltQIJQ1AZBGfS2WSF95I+zlMdi
h6EZmTgh+uwacoRJvS9lurf+jWkkIuPugSuRhWmOr5Wx6uQ8N7iLNgliDdoV
YRN84bzc0RwR6YMrcuT02y23ZsVv2NmY5IALS8PESjtBU43JffRooMUCHO87
n5KRiU4xOEXeI+oD3kJy5kI2Gmr0NEn1gwYqABLGyVtqr0Z3SP4tYrl26CY3
vuj0PfJzulFZloIAGg389kEmjWO5SxQ5H4MMzMD7nqsW07SsE1w0mn4mMbiR
5Zx10EHGuXFJjw9XFzDb3eeYgUhfMeH9IxprDSAoCYGXIsJSPdjtXTHic9NG
+mNA4ZyD+QvC7hP7jp+CBQXUrhQyBWcrvMT3gxrgQwqnraUzzAbgUAcLGWEH
hwaG2THautuPTgidZkK4GqcE608Lg6X6ZZx0ZR92aO5pcmp5B79P7ZZNyV63
iSN2Dl1/esjLPPn7m5CWy3Pzg112psmNLGWzeZLatR1oj0T6NOKgK4K4DRvS
2pHpb6kq+56SDolb6aZi427CyOb9wQUCcLDOLD2J+Gh+Cq3QwBT9BUli8/ih
SMDTPVEaftfLaVlV7PFB0/+/F713Lt72LM86nABg6DDg+tRQYFVajUFaybjW
yVsHwhBQVshPCoj9uS5bJpaCAit4RVpKEnegFByFPKDVxQ2ulm+mOmATev0y
qbLN9S/K0wAtkZqb41xh6ucUbCNFOQKLkH8il6RabGE+oxCyH1wyGPByd3Ur
nToS1oE0FjbNzoxskiqBGmBNgJfnxFpbVMcxIp2H4x5PUaButiN2HBOrxNP8
+PncCe4haJpfRSw/Gz7iKGyOsBLJ1D77JxenpyTwTit6so6jI+T7DpSq0o88
DP0HlX3lYfPHJLNyCj1ZdUh/uRuIoCmGtpARgPNEUsSrMa1tV2B3VhnpfVnu
DYLJR0NlqyZlwRefcVRYRsd/JrxQmtvj80wukIJwzAdkh3C69cImBWwKwUnD
ksjAjB2jrKA2hUqxN5Ya4tJeAfX6z1/LM1M897x5hd6kTR75Ch4czbQ3A7ZU
0TGl97GFUT5B+aiIIttivh0/KFMCpVGO/M7Qr0Fj3XYEpmzXj0eLMUGQOxpb
Qpt1mBZZXx/0l6LHGqbjjq4u5bjAIqHvHu72P/4/58vH1UNUbA4FBgODszQ6
67BPqOxttHFCJft1vgEzbbWLabelfanzmPaUIfxvwkWiLvBGDcllCk8rY3uD
ToiNZqyKIhZTZqdXEn6pBJ5LvNi9UmmGLNmQp6T9f5C6FOaJ9XDV/KytDMe8
SQaGq4QJGIuJbva/WvFeXELJI1ZGgSkoR+p1nqj31TWWujo4VSAm9rgaRFzW
SV4Bj9TaxjVlaAJYQlN1H/iRrDMKvEPTgyn32R/OG5blfFUJIpt6qBWeRXcM
5zDjHXmHwEAEnKLd+RV5j/kI5a5s8Dp8HzSjPTkCRcwq5V8IG+EO/3J9nh6+
zeWP38I+6dOaMSTAkx+4BHYk9uogzpUHKWnsLCKtr7tLh44kWarLariCBWJj
y0bFwrghQXVobW7hH44M45Hb1zoAyDbU4w5gqqLoWngXBaTV9rRC2ED2Sw/w
GurH8oSg8sWyt5JX4UaRqIj6TNVvxJdX42OeqJpBdOaK5r0CPF+a2fnW45Lb
Fy9NTaxDOaxIRVGO95DLXPAM5NcFlb6JHDg+sBgnOMD9lcyTScB9rzhDXesB
iyyw17rPJwN3LorUAWCQnfbAfX82G9djJKWCZCtr1tHitynGn3x1S1zG+zdL
rP2HTX+ngZu8/XBQcRloaRCtMrWOBGfZbtvKyGM3cn77FAJHE4P/peiTPjmy
QKB6MxsPYZ074aEs/XY8OSGTPNy+zggob3/hfKAySZ6E9f9y328t2ZE5duay
vlocLHYNaTRMUhLCOtSYpuPNsnEjg/17nbggGeHMQv6A5v8SwkuDGoIji4O8
7/eOOjjtdGoZA/UEKRZKWDUBsAdRBz2ow/pJrb3/L5u3bPPjZl8PtgEE90JW
R8U9Q5fcUkFAaIcw6PiArHt7l4UnvE6mwTdardtgJ11tWzUgb8u0hmqhzrdD
hSjDyXmJySM468f/XhfMjkyBr0x3hPbgGMZVz778A4p1h47ufQHcLLZ1dtIi
L7sv9l/d32nwquMOQmxR2xf0oVAEpu679Z3vH0dBBFLxGAsGyUB3QUnJkhiw
U7UzIcG9hr1jlLMCmjmqRHCYIlZGsT8ZwNIYzEeETn6CT3kac3aLUEpn7s4K
3w8A9M0UnZq9lXPQKSPa1rxgd88vxM61KL0BCkxiuj29tSf+R3jyrmG0jV4S
u7BprI7Q0ENeXUhaNniBGpr6I7EOa25lB+EmZnSJAm7zMvoOvUMK2Bg0Emjg
9Lg6gxDVH/XjCRUHmxrbAIUMb7BfsU+EejDl3XOTXbPmjwKatjp+gvmcSOz6
AVGzsq3Wtri68hWJDFjeerYCeaGYs2/za/5gMQWIhTAW5LF3QsnFTzzGFf3u
WcWykhgKHDjvScxHfqhGErjXaYAL/RNpqgsZiiEJreXacFAZL/r1w5RrwwCI
o+LMpTJO/W08W+qtEe/1A6tvUSDAzC4CiRoXSbAeixyd3ukRbVeFya6X4Yws
gTz1pMFdrB14s+L+wCPB0aFnUXcvVBT1lSPJPf+xXLnEba80nLPErVPoOVS2
5J53BPsuHCukT+eLIdRHZUE5tTE+CwKP/kX5Gv0Iq6/Qvgt9Fa1fBjSFjp9G
RPhrJqSNRJAq5npHupqL6TRA3xjQ0lf9/BdddlCTAd8/2bjIBD8rQzvMc5jC
V1+6cK5Iw4F8d/CY7owKbAxlMM3bmZNvncVvMEmRI/Y7eJbK26srhjlxSz6O
Omvlsf4/P1eV8rvuNF9pA2qPEf2d0m4VUGaVeo+E8B/Kqym9zq9/CeIiOLtR
xEROV5M72OLmFaW+IHr7dPIrlJgSGPh/MIsOirrt9LKGG9HLVqsmMQnItw2Q
09cAeUE9Qk7d5yZ/KR7WWb8gqa7OpC+pn9735QzSMZsg48b6Bd3qUVAbi73o
/1Jj7G4ZdunHHmiGuHst0deVYlVHPhlhoI9rl7k7K/MnW7bWxQK40Jc/Knn9
48dBOk10I/HFF2rylApnONR/hqu/8/iYA+IsF7EjsBAemn7gRFXJwNQc15+6
w/s1R2S+n2DbVflmY7I0pKWKJS0nm2762puhIMyR18zspLwYoDcDs0mDJB/P
oxH3FrzVy8PVmUxldJ2CIkNBgEqP58a+ZnCWO29X4H88MQiFo9ERmhKENn6E
25EVVsWTkxg7R+GSu0rwBj1BF70N+Lb7fO0ET/jOYqZyf3KTqkZ1JbfJlvn6
a2hZq0wjU64vY06P30xYkE/1WcAw/D0IuPyGo573eCFVXTU0zKslKe2HTdbW
2iF/KzUDZSlX45D+F3hsSpMulSWgqFHrPxbRVbUS9JgyhHsejwtD/DNt9gfy
AlcSG6o7LfLsdVGqMz2e1NkJ5FXZBiEXJaLNnekCJKJRYEgw68KB1JvWFUtD
OaqlmPtEpXAgO/m5kxxZjhtEqd9M8+wR4z2uglK2W11BIVZaXtABeUwsEdJE
qnVHi+znaABP2f4pgybG6RpRte6GU8pAotKnFKi9wZelwfY5jYqLL2CBOysT
cljgMDpvt+MaVy0S9YqaN20IhOB7ywz54rtQAtVjiE56K/tos8/4h1Ypoqdr
YaBOgDAbe+7Symlp8VbJLoMTOx2Z8BRNacTw3A/q1b34UZA9Fizqq4AaWhQ6
UzeAt9yMFyAZblbCOv1pSKjyOVfQfhKuyCaPBnRTFuCQ0CRH824Y08oqKzJ1
gPVhYlzdlOJ6Ch8dnMKCgF0f1CyGIhFbXHafVe7RG0FlZamAEGfppGjIMtUU
O3+Wh4m5pBJeykjm1oylmsLpGg70vpnh+a0cdpo2IOLioj7d2jQCeLibTqwn
0zFCImG2Hw2C1qD4YcDwYTt3RYmfo+RQiBFgkgNYlo+2QBRt+3V+05HrnzBB
qR5x9FOq4OpY0RG83d+ooCQ5skH/KA074nrXvrh5pflh4DeAWVgu46JNDivv
S6KI06AyWUcBBMs1KF9Yq5MflQ/MWYpBIgZFMNNjdAJ6s6Th3zMJtUIgU/X6
+hW9OyDSjteUeELffi1APZCRrz1+TNAJZomH/OaB9W5pIYvfeK2zi5BhKkWP
TNeE8/sOzOmVkEzeMifn0FEmq4VQmR4bxXO/CIBHFeDILAIjaaI3U3RTtvxi
P9vcFBpOngx4LRRTHAlGSDM5J3Ew7VGF5xq5QCXLFvJXMfTg6imEC1HX+9wp
t70c8uq3RdH9Ewgiln84eUTLm6MjCXcVX1qLlF+gvwFyeqWaDQF5UE021BaM
/2Kzln7Fj11/3c7tyRHJcyasNt+ia8wxBcdIg09FZj0m3xbN0FxZara+jeKV
edc4LftgTit3oQoT9muzlR2AsAJvGDiA45MvX2TTJ2FswlxHjpJnyYwA7SZy
KwLiJAeX98g9T6GbFfRgTc4LgXWEr1lCM64jhoXhRk3GmrQ3SYjwjg+yDC/s
1JoJmvyIcJJYWyOuXEPFrnDnzQoS1dohr1g726OPinzTPV1XaNuBwt0By2Hv
XTqM6KGGe+x9V+dPUVtuI1E2dWzRdEAa1HjxaDT1hz8Dwhp9hIH/Nv3w2S4P
KDmyJ2Ajm9Q8dO9PAOEyqwg2Fnb7qpoYLLRZXrPerk3zvqOQJ/mQKz+vihjE
Ow+CtXpG32I5ffGmmiMwzvBdTEGDC5qaXJXJr1SJCsyV7NcuZIlSRrIbSMng
j3OAwQDrKIBS3C3LmsenRnjf3hBVwfDBEfFECFa56bg4ut+m1pOn8lMd+tE1
Sj+62l5ukHs2SM/zGcrSVFEJM2JAcOdeBTiI7W0kkVKQhC1cm4xk+9qfgG/h
/tWcFNzMU3zM/rZrVFq4Dok4+icoUCEMOZjXdlwFLIZQCeBZRBT0I6hKYBjm
esPMwT2dPmosGxxvillWbNPGiaqDDx8WcKBhftvJKUDJMyE/t1+sQHS1mDXz
IDEfBwo+WE0bPfK+27evAhgLOZunQyx2P9yOt9LcQXJJieIanqA6TDmGsj21
/mYtEudAjd0FLamJFDeNQuULhwR5gcyVcY6waXbrQrTY9xENyGIoiDWoz8pf
npGlPxiWN+xr+m1/AKkudzkW0RvU/O2TLxdlLoaE5FK5rpdJ/rxqR+8BTAfj
sFfFp9mFMQTwiHOVUE6b9fvm+rCEvLzIWVvFtfGa7geSPrjFQoqGRPOjCSxX
+sklGFzmNgi+hQqY/hcc/5H3ci4Z2GljN1Km2ms/IHVmfwTosdG6Rn6LTLAR
MLhT53IKgdAZVpXweBkUjsMvTF33E0z10Nv7X2koorbYEPtR9FlCXb4x/8QY
02Tm+7YAwZSWhNpgyhPMi6VaMEUu4hyc+N4pjcuZW3wcafO83/NtwAwBGMOA
axr4CKgWWQJ+4+vIDCPA6lAiVyQn4ABPfAONISlxDNignUyoqLx674bhq66k
BbhaybeyH2NvYghfhmtpBXtUCwu9CMa0mamr3PAisnMmS8iMJHcslSdMBSfu
LYuJJSCjazxmX37MGkUZr9riyJyRF67Ckd08k9XZsu8o8OKJenG911pzJZAs
l4cEvBpx/Ry01K3NfEkK1EIqqEFHOGtcWjBeH+SzMsMtyZPYMX9aDsRmDic5
HjDki6vMn6Edl/fy6Ks9s0iCLovwlZZkSxWdmB7RSTspMWEA8SQa44Oa2fhv
RNQTxae4g+l33/teAYSUPkWLVun2z3vkthjLad814GYzb2TmPtZL+ODbJrJa
UIXK+ONIsOjfUI7WXUxPwNsouHk4JeH+p4hZv8rJ9b7BEpV7wFM4woTSLArR
pklmTFw4uYKjefQ3uF52GZwpOPxN25ViKn84SPfBAHsWn6u0xgPUNpicHjop
+D19/Azwhgwr0UkXTOvMO62vH196kcGZcWjaiWXohcmVqzNoq423zc6Te9Kf
/ME93O0lIuz+B/c9Slwpg7lEEc3aIrdbNN6zMUJToz/+NMbf+VzsCnHnehRB
oXVBzVZnhYPVM8Vfwkxssg0Y4OvQ+JQ/H5/Uyh2FswVvuwt37Z3X5aBVrQZ9
uHi2DoymofHRCuODX+TKsA3Hk2F2+WXhhF1VdQyukqqMG+tzpy00Z/F2ivT3
uMJoveBsd2FM9CwE6k7QGi7lZlTOwKlO12ShEMAqLu5CPpRcxpymOdML5NtI
Shm0IMjrMHB7HdcmHZKtw/nQDb7PlZf7i4G5Z4s3Q4+q6xwTWzVoUpUc1vs+
8teAgD371kgaYAcbE4LFDXdd1Ikkh/tBK3QSaFc8Wy2eEQjbFoAxQnzmZclQ
VlP5CTD6LOGFV+57cB/SWtkh4fAGUgZpLR/IQNcks3jJT4JzSJqahxUC0gLk
ef3SHwA2ijc9iL18r7+5MZ0ZVSe9rpT2WbYosX4MnTu1/a6qERvjpWjv1B+H
cX9+fSqojylQV2lTTF0xfRfBsj2cVWdXYptWcXvdLivuxfraPE0yk8AUdLst
k1mgqOQ4xGcULGiV/nWSvJrxcOKEXY2e5DFfC1xIWpMKCOYz1SybcJIoOQpW
Tlz5MmKcJya8Wc44kZwyQm9ogvVsy6TXfPCUmiTV/DAcTqDTO5AuzFLdpvRg
N9DYXy5CQJdG1SzN1fZjePBDfnMgmrmzww0WbgbDxyGjuC9NiGSoSaSgJTeg
O4rAhmGYC0okzC3EXR0v223AUALP/EsLu+gF4mrt34OHtkkky//49x/0ICbh
h2zwlFUvnwREBvebFyKnQjhimhDz0urVnFjrt495ZDcGxeM4D+Q9bInuWeEd
kXcOWbennspOq2fjoMt5zEPskexYsSqErtuz6Ssv/utHtcLaDbPgicVn34vI
viACnma5Gisw9X8YAvTdLc3UIUT6lPp4wAWO2bSHgkI5PNsLD1vLM0idJX1I
WtqzkFN4t1OtB4B1jpNrh3BJXJy7QAyk1cusPdXyXhFomrG9W0kImVzw5QQZ
GIeLRn7IBA78MzAt0vlVoCktcLqQeQnkAOTm4t8yO5tFJvxWO233FDCCQ3tH
mi8T7eK/UTbwpA3dpY6yn4zghzcoKKBscBOkOAUTnow4PvGXHi4WWMOKNkX8
rt+3e/7yEJp3z6f9WwpJ/pTvJiqF4Y5qzg+aef3H6gug8r0uikegBaHpvGy8
15J1K3HlSM42vOeY3RhECKijKA7y3aGijnXSkgCm2lwI0hKgH3LARfYLg1pn
bS+QimmO7iVrbNE/oBM4e0HoMIBvHZzTKrB/6mpMMuvFeOrF9izydbe8T68F
InqESZz1qBKumsPkAQZj4lEUs/3mZAOyakdqU3M4SQ5PFl8CYUreFdudJL4w
QG2mGAZoIsIwbGQak/fTyY5P9uzSN005iuV8x+6TZxmZ/QKJk0wth6tott/2
dsJEjaZsHSk/va4VZaOYELgg1YFltv65W0rCTOpevjGMSUKqvdhB6uM2ttsc
Nu/6F8fpFT23RMsdiEu39Vv+fHvdf0vJlOFTGtpPAuHZdYhbDcoG+NUJw+Ih
KsSFf7LtP5ug1spChEd4C8Y7FZ1oO2zjivUvWAXAy1+75Pd607O9cg2xFJDf
5uO4j7a2ugCcFrTJWph9ocZtiiVHjuclq7Mci9UwYFky4vAMuZl7MAYreduT
FQKtx4WO2SAa7+cvPm7O17bHEpSKMiEX/BBXRR0vUsxMJLhmzPVWa+fJ5wc7
dNqPC8PpvqjsxxESoW568W2jgllPo+f0wbFW6+NW0AmcjJyOAPY9qcMl5aHv
7lVjP9c5Hv+85JW+Gu0JU3OC9Y6kZPpkUZ7yCSm8pshyGZeDbDCuxmfSxdS4
wACoyq3Wm6bHAi8LrShFnvJgDC2fpsxtzrve1Gz6rSVenuX+lu2lBnPZuQ57
zQxOojp/y1WQGDh2BQDHjXpJ8ZfbzoSqeLpz2Lfbup4ty3BX/HcSIQttU0zW
d87nxbF6sJiisYQ5bEuB288aPn5WzdjYS99Tiw/PeUphgVelo0KxYG72/BTy
JRM3QOGNOSbOTXX6zEzYui/pvaZ0CBsC/VkhIPaG7ImajO/B2uPlngbWOB4p
IM3aPnSRNPzhS5FhIh3eFda9uXcF4r44B7Muhkg6PNRx8JGnJlXaG5uy25qZ
nUGDprH0cyy3o0m7cUpVczjlHad+3ttKhWR/tURKXkYjarYnZNKrj+KYMlTr
as+RxQ0pvlq/GfXGjg8AaMNzKFcPR8ns9vXFLJkxshKekI1BHR2qYrHEiB5x
m4dxUR5Gt4K6Ah2hGeJuVcNs+ebaTWVNxFmSIZVwOVefIR4v+AZWDjUXW3zD
fosscI5R7OgfWOaEnZwb4fdjF7GbrhWePay8Cmn2IcveAmbCJ9KZSI8zF2rN
dvNpQAAh218Z2yJ4xqwjVNjVrCojTn0zoGhy9czteKQcGbWpS3AxrC30avic
NQO+i3WjDB3cyxqxFIg0cQyemFmRPDbeqtriHdw92KkLGhx2MKYekEHkianE
eX3SUjCIzNdFH/LIxGObV0ETrbyw5jX2iqStNX96lm/XtIClPsWkHxjqOwHl
kPOgmiCE2fDvptQm+MHPZxszAhDm4DorK0scNzDATpSULZgpRtAtyvmHdriT
D2rpvpPRvisza3R1Jva7X0nK9TLIFqxDK4kinie6bWr9xeUWMDie2zCjRv/2
lUardp7m3r0qol/XRxEYZeKCcYZlXCQEafRVxFlflcjkXFjlCERz+hO4IIuF
cmz5Cx0YaudL9xh5fKZVnvmy+dSimpxGhh8G/q70XjG0SHpC1DTtuZnwdwbz
pF+UKEuLVN0w1dXRD1SjBfLKSJH1zVCXVDafeZJR1UsiPxPjN5aAhXpOr7bf
X+hwkq6pu9PhizisryJl/nIfBPn0qLG1/eDDkEiQPZY0R1Rde4p+WtmFH3zp
14TtOX2lpHQUWk+hDLrEqwieAW3u2TBfnGak9YpaLW7g3hYEZHFTr8SvcFdr
MEZ/Vf6+tW/8Bwiadvlu0PtQANCe2Q16VVOHkw2c1k+hxDi71jVXiR+RzCrC
ynhTtGdluvRqN1o2cz3BjOGO6LSyfULJPZQ3MC3TaPJ+Yi8gUpVje44IIrge
mR28QnojZDG3BJzxAlHQrGJQ43VT4L1JUdwEOCzmzoByxOtVG3CRn85D49W3
531BXhWBDgdaUNUigfNEEK9a9lvYCy4E2CDg4ZRuSZ847jLfGO1KVO2LIOSj
8LrOox1FgX9nQoTzLlCVjFSGJyM2kkqeOmtcIdOSIDDMVRTx3Nj+dHqb4Ocw
f9G6sBcFiJEFfZ+IseNJB1ZY59zkgz1QPFhy1dsu0v8WWhcauX/tf+3q7Z+j
0fly1EUK34J9u8hMPu95fRJHnjpBqOTTu9hB3VDd6hY56QO773rPZrUsrj0j
/GfMdu31MHhyPtBza5owNhPxvC6plpoxsQuoiAr8MvPCdsEvL78eQiCkpzXk
S5mbQguecFRgauzuybT77bMJmjLotUdZEhTjtZqxHjov7okxkgUy9UDRl1+N
m7oDbEha16cg2DO1l54tl9hIvE4jxDfcg6vMrIEED0GxxBbTJiwVP9nuDMNS
BEHcFAnzUbzCwjb5qrlx4DLuLTuiUIzZhdv06nuG5t9iUwLm1HQZz3qj492m
fiA1sQ5gxC6muxdd9Ve3ZdRWs7r71KnnYZWCUOWjw3bJcjFGgI19yLIVzP4W
8a8ySHjf+vbKEre3tz5pS0VONS8i7+Hx320pW88IKc8tEY4V44sLj4bRBEdl
ejoiEZaGRzp9Ts1zxxh8hm+OuojWHDcQUfpAIiDIiZ84OWvdM3KSOudqAi8q
YUVz9pnwpJp7FZmMKaT3UdkrNk5M8/h9h2R9wtxtQheeg42f8sSkmFYlCBAK
/8agjz48inhUYrmsYclGurN/SpCsfEF4AOdj5scywiG0MUT1TC0h49izquaD
bP9uHyD143tZYGsDuc275T/o4tOsovkFrqP8EIn8Tks8q6PLQslMTWOOBuaD
Y4gIvmpyxaIr/YX1dDDicKK4IR2WC5pSojEy3z8X6TEGo5H6NOZYsn//H4/Q
DEV/vek1v2F2/uIlk643gOfusK94MxWoYm7BoLqjOtHk/WTLea1L8BCfCL10
IHn008KCPowa78WEUabfFh1huLruIDYXPbe5IGtRIzGCJPaUWCIYHo9tvNd8
mq52KQN13UqyWkjvjeY226gA2ebZ8fKr08Nm1CUrCCRe0faIMc4DwSVldhGJ
mmPd0vpBI5f79ICP7hESbZsxwgoo2kdUPd7fs/AfaxD1Ybph5U3zhEWe8zrt
USepYEdQwEtiQ4MwWMOGl0iuRnWq9P8BIDmTRFf0C/qMduu/pIizguBJTG5X
ifEnT/DUTsEZjv6A7z8+NcLqEsjnNJ8kzUiBxIAo0wn4TiJPaAdqgS2ULGGe
cCphV+vvWz/QG5I44Me4WAUyPxP9Y39vKXbBLXsiefupRCyY3blqb8BHn0XD
ZJRXr5fd6iM5FOuVgkQVqMD8VFhd7nWGWEAv7WLGA5h8TnP5xu7IsId+Cu5K
KyYR4alW3pA0kwEVMO55gBM2r1VAh993GHNVecurDQw+usdBVoNfnkl8xTMy
Zsgsn5JUvUUFzAzFJThJhgSoLZowEYX/UoCVsGJa1BQH/yGRG2TaXVl0s40o
gBzVZi2O57FtSg3DTWKPXN/SsA1PL3/zAhyBEe2HRfJrZ9foKfhNbqs3ysID
HYzcSeJkpeEUvYbvvyP0bJfHYo87O10hLgpHkzu44GVCN71as9YZCAGUwOgh
vfQDfywV6F347Kgw/7iSHpSZouWyxctrUNtyLoGz0yXjl3qDMovkrumTU3iq
eygigu9wL5dc/Yb5A42ofDYVaw1LkODFluSoo0Gts7PI/qUJT1DqWMZXjdXv
uDXp1iMaT+leYcV+7mJlEqLZSnuFm0A0L6tp2Ydrf22WJdh7TjfWrW77E4zU
hAtxrxlDuq5aE8vf4xgihKN4ELdd7ZUnrwF/tLKXBEoZfX8cy0/cExF1sG6/
yOIg4cO8LT97XTfqLb9W3PR9E6Ge3gqlxRsqc/5FjBqp+hCpTG6sWXVpBuzy
ftsLqcQupEdtkH0/CfHXnJjDdMR+hGY6bki4ObscXDU3ghXuCBpcIULU9w8I
2yDDYAsvoLO4Ce7pSOYjPlNhtmZADklJZLMycCbRMBP2TRe9gHTm7YkkZk3b
kHgJDKIY9i5KNZbzWU+I0+xQAz4HCzrZTCc+O30CNi/w/6tGGbP2Q0TSh3/C
oiP9j51R4zGr2Xpu8xidyJzvCFy9FOC6cwMtWC4nk6TZcbQfjthJzGdY2Cpu
ya92GmW6ounh7gXlXrkZbeUosqAqxZF9MtZ0k1bZqz5enYDGJR22+4kaONFe
2FgzZ6nUlN75kDXBoO0hTA3m/YwWfkQD5WXB/TVPyasW+TXhLUaFsd+KSCBq
zdg/sa+PLNTTyyZt1AT8bf5GcUoI41NiFz1l2qYCXowoIKeI+eTKvkQV7/Ot
gnYDjoNKtqeSUfqK3SDz6hPXZlU73tclnmEULuWrvw5w4TK78z7llXHC7LH9
hzA/RcVOeBHX9jXW38ZeHaI/osgH5330y2xKkp8T3ybAZWSwO4J/hNrBJB1Y
VN3ifRT8+RTiD99coeB2PviDUv7WVT4Qgvlmths/yAo/b9PidI/Ab+ZHOYb/
QUolBHJTgXnSHkD15rgIEHJv/F6PjzMW6vVRddpoKwwmBFKm/7/WkUHsZNzC
48f1siz3Fkq1V9dOR+5tY/xQLjlk8sSWFy4io+ccczsL8jwUChyvNSkVTfMd
B13OphBNUVhNIUpGsYVPN4CNMQG3UX0pyBWppdDLv7hmNRsJidJNk/ZYbs4G
wt1RvXucEcld19F/GpZqEM/G629DOGuhilyFErF7k71oNRDgvFrE83hvMTKR
pUMvaGLY3jCRbfHgjHroRcCCrqKE2jl/ectvG7FGhBcDPNDhSLAI+FzpecJA
tOSwJ4K9HPf3h0p+udoRkbdte0UoqgzuVNzxMvZX2QQ7PgXtF70WEZ6AGqN0
PzYpYwYi+aqi8nPLIOSG72eWOwfBbXtL3ElD8rme8vs5ao6fInAk9X3siF9c
3DLzeDA8etK47TLGCaJI3EJCs++JVHeBqLcFGbEXi8sDPO4tOiRD7bCxfpRD
C44td4pF1HPqhLeiQl/FDrHUm/r2mK0HkO8SOj4zFI47Wd6mAJnHKCQoUWFg
2MLYMuo/kzn5+z5+7v7pru45+3PE7LxTJCXWwX3cCofQGHfqifPqT0x4QVrA
fwPWj01DdzOaRCVqoaqdYYzm9+JWAbt8aWBmDjhcU5O071HATnDdZx1wWRNA
ysVV6lTmQJyZUex9uJ1HhnnCted/te7oCGvkXhVoOfOODzsKyo/S2uSFxAvf
ohHRddbfcYiSKOGQCX0fvm3nZSpbAo4jAaX4xcLNW96Q3mixC3fy8jWQuM93
ALvtlTjlpVatpUyDURxqjogJj/IHrvHv9QYpsP2IxQt7hP4VDaWkbom4V+Tp
42fdZLRQIUR6OVeEXUSETJxPyw1ZPA5LGPlh/FtcMROG2fY2ttzWGNpWVHw/
U8zPWPoicyZasXgbxwMNUz7+Gh1r3qOGAh3dF02xYQjMAWBnqmbZcNaMHcTy
WBfZmOa2c/11bTEPbRjhjoQmficT/VVvXjIOoYIIfYqxb77D8koMuLnKbqf7
m+HvK4rKFpc8mnEaLzmAiTBa/INraEQM+Dooyja3xMeweevxAplp1dSxHonN
jt3fIfWc98h+BuSp5ur6mc+HLJPC2gAhfkaWNehK+5hx9Z6A1J2X6NX1zQee
wzAN6z1dLNKYWjAzpAaGOvwjIAk/+3GU0uVpj7pBEqQ2deVCefLog8NmKPHo
yPTVd3Eym9TriHc4cbFTlmvNwFkoK3Wy4wj2sP85793uI+zwSezcWqYu2H/Q
2m/OZJaLlDU6YTQcm8WQ75D0SIq3ZO102Jpd7Icenr0jTkGGY/LpHwScQMir
RwC+USw+KaszhpAwhw981PWrpSwy2JlTqt1FaRevCx26JawDaH/xFQgRT7Hm
Tp2hQMdbUU5xwLQz6yWBrwyDwbdSrBngjx4ZHhMlNH+gdpTlFkQHHpAMOtKW
YRsJnx1kUQF2sMjfZOUZvNmyLp42FXZ+zoh9ZdTQHUyVUHBpt3cS9RIgF9h9
GzdSPjB9TdCupsIrnUvpalUBopM3r1reSpUdZH87Vk6how0Tw+eJapwnt6NY
8J6LAoXWosJX3es7N6uGFb3riESxxwKFBW+XZTHwuvkBScmGOjPyNeyIQf4/
yEkv2xLhjoX+ySy2OQctvc5FBJ3+9+VNrfGTC3FzLDhECpooFypyBOaZcaZy
Fuuikaak3U8MkeHjW96csQqZhqETSLhc3Z4XoM4Za8nw/JGXVFhWG9GUoDYm
406W8A3dZ+LV2Pvij9uTG/XOEjPjhgE+6t1rLfOb6eNvmzdFMtBMinM8iryw
D/RI344j8rZbo2aJvnFpib8fOnDWCKPgiXep0TVs+6ZpSjxIhBz4X81iDScf
Ok34XsXv0k3GJIec2wXZBh43qkLi5Vavg+qKtIKu69nrNeOZ2nOeSyft1vH/
gnJ/UO3w9kXIq2pBMmOH379ib5lFIu5JVN7zY16/XodrNaAMEMa+J2VMi3Fd
xq6XHRdame1EISbdH9f1czqLEN31+iQZyBMXUev93ZmCiJyr7RE8VbqWlsAO
u+dvnr6qRh+qE9kOkLaaFyIbVfBWFGRvgwWCkRehMvYhMqVmAq2rv88mBu0F
g3fSyOtIzEHnUFgkaY+Bl3qcJMAGISze/MeGs4WsbTyKcIXW53qpl6O3hly8
49w7Ww2kKkHXhKR/DYT0VDmGNVrdMu1Ec1mCf7I3Hdz7lMsbb3rt191LNlld
YBUvdMYQt6H9ONy8rXs0dgcBdVsQcjnhvRUOVYDN2hXVEFl+eCMAJiTdLnJR
XywLFaXJJdHBD+aEUNmtzMPj2z7BIohmToobfxnxeFDhsJE9w7Z4BA8OAhmF
buZ/35X/mADj4Px/qHiLNb5eyLJrhOkG1SBoRIUcBjMkDdri6yH/4Yx0E6WM
qM0HWZlx+XDd1SKs/sDCDCKgtpEACVo9DMqsmHuyvSCebSGoEK9uS1kxwF4u
OJTJxor0mDyiOA6LoNJzmzSOV0BlP9SZEIIccQAw+xFUYyj0saDQw7auCXQE
RBxWlPOayvKcKd85i9OQlrOmBeSsbzCRDtWXS2IyLr45l2klSc+DHHxJ6GAV
W/XdhC2tVxl2ozBI2Wj5VGzXr12wwHVckhCjlcpoa9VcnEPxIBPYwFMHd7rc
aR4/tcVDqfrHttkUnSzohS8DweEZ494rJ7ODDiggeYi7Ilu9DmGWFiepaT4d
1dSq6RpyWDQrmTldSx6FVBbvCoMJpnbuYVYpXJMr1Jwb0WjTHh2ZvVvJ2ZWQ
gBvST1U0puF3HK1c2fhlnnFRSX4WzTLUQT4gzZKLUtidgP7Ho6kngNLDN0UG
3dqrP1EFuNVFWizHgTQ2eIQ99XszCgn7F8EfC24QL1k0TWS80fHYYg+LQxEC
F3Babrt6mSRrfMqYea8k/SxMZ+kJ7UxpbL+GFWMOovVLnYGxjIwiHtjpNvu9
5G25Xqlv917+Im+NiDrSciLQzWKbjVTYrnIPPO9X3Hq5F9+dMJuidfs2Uo0W
y2WSENQhMalFLRHfZnSgUs2Uit9fHY+QUDhRFjSvOuUe3Ko6+H8Urj5Fkm64
sgUPQSGox1hvsbQHEwvBn0pvp0/hc4hKGbq2+Wi/BAXQQYbzzFJMKBIoL51x
AiGkrcPH8KSJ03eYjMrOdlGpNskWMl6YC93/KJa11f/HueP5ZBNZcHtJ4+8k
u4Xfub0tFpB6F5ntNn7LZe+8zovl90Rb4+6NbAULpvlecaIe3Sd8GKnlQuAS
/kKKIVW09guNIE2mvh97h8xYpuMDr2lKjCMJLI5NwbIZ9sBkqj0MyFXA64UX
CQe/bu+p/c4qiDSAwK8rbq3dDBKpyqvm37U5Xqb3vREZxf6kKyKiWRABBFCw
edeZ7vrSrt98Mjl5+wZ4jpkxBeRB5zDnuIKXxv3oMAD8GG0pFRu4fC+fc4lT
IuHipxR9sCqzkrh2HdtN818X6ejIWzh8HtV1SyVwcBxHbkjkkWkQQwXlpv08
8OgER0eyDToSa+ACF8OqCBQpCUV+2fflOQKl7P1JsutajaYYYTm+iuWM8rMt
pGxCYUAo0cYwSY2tOTyuDgzN+YeaUc4GVitYIflzsisXecibSRg1FVpoqIbC
0rxUKlrZMpShzbWeV5OA0ED8s6KYNIDvV4tSEVarvQssfgQMkiRByugw9KFL
lDhoR8h5F0F2tQrU/GcL8GhPn+j85sajunChgvdXD08VI5HY/7RV/kaIQT5R
dXdKaZJnFXEnXnOJjCJtE3KPXTVJ7e0gGtuG+iLcSAhExxCRiJW0Mj0FsDyn
czZ8vpxUJLMOO1/D44e/+mtUjV6j6wk70lkGGae9fYQn1vKr4Z6yC57bRUqY
B2VpeJ+vG5xQLd+QzEVEiCha2P43E+wm4amSgGJCJ57VfDG8yBzKBSqlc84g
fs8pL/JEN88heIAG1oA6I0NdfxZWi8iCiqQ7hUPqW/77BW6B2n58+6OrlqtQ
MGPcoSCZU2G2fuwIenVAHcKIXOZ/kueGFnRuvuDXi14IlavXpFBc11dnBI6M
autIh+SRBN9Zj6ww2vLSqtMkIRQw0D/3Fe4+bWRVJ93V5FqsSQnJQRGx2rej
QS/OlblZz5w3//1LncJ/bWNaiyt+RctkofSmbZ/m4HFCD+FGdD+iscG1HmCZ
8CYt7pHOpT+G9zJeBCShWxYODe3Mjvsy+sFj+xE6fXAWoWGLw68GpjsMm5Vo
W+vSMpxd6f50QXCdp47/0iT37emU33+Fl5N91pVnxLw7GdlJPnS0ivunc62p
pELrAh16m6JC7tIAD/xeI0fjSZjNAYW272+Qkr0PKSbmgfsLMhE0SbTjnRHy
HtaqUkhKehmcuvYZMWkZ9+m8Kpxz3YRAi/OHU/IOCDQuVj1CmtqyoN6VyCDo
KviwR3lrMwjQoj0rDZEBtj8fRmLYYsCljureAQBDLZMBZKZDJ5OEGRYs8Af7
kMRZn0jnjhpOAA+//FSYsEOJneY+wui/QuihZcbdKgxuuuzg9GDg+HRnvEKU
nnu/ON9JxR5O4vXzvToGz1KHwFr+HrXRdOD2VfGdnIhSkwyTG87U6hr49Uks
zD6NgjEOuUxWsb2YlwrHwi5y4uhX0qOZAdqejfjoS1iBPcUPxy8Pi75uA6un
fwZOD7RLq+FBJ1lcYoYi4HgUBhBesbZxH6n1eBD6jUJsAIVdGcMfrMj/iP+3
pwELjsCah2IEirLAPceNByC73N73QfdQ+hYKV1HvtO6OpW0zeV9d9EI4Rq0D
g8dR11d0SYqzGXCQPo8u7E7xwPJVxxjz3FGBYBJ0W0j7sL8T6KO/mwz/kadf
dmSwBOzOIMA9UGcZthdxj3y+T4/bZg+DJIqSKeeYsU4eBf07x9OePwb40E2K
kucWVccJMAYhDNKzS/cx8iPXpZaBVYlXciJBJiRX7QNE9/TzrWFPQTvbCUZT
Rx+4LdGvOGXeh14CvR+R0vX7NPvy6nkk041d+NQFAPE0p38nfX0+Wyws+Enq
MkNLqQs7/pv4eFzoI23QGkzTd5DqzuO0EXBKgjnQ0Uz7d9w2vqla1uaGHNAD
kZVsgmvaA1bxvyViGq5YDF2/35tlQNPz7IsNeWe84vUA557+75QjqqJJAwZn
IAAdPW6JFCg5K85viRs+RT2v2vXIzbZPxt9hDxE92gD083suwpKjAcQLEPHB
NhlQ0MANBDLO9+a2a4nCiI27A4aMiW8/5dXD30gFcdyVL47n0xyN9SB1hcoZ
oXxp5m7MUL5mPRKXcpU0H7cwVTJnKkWXdLYcp5FssV7qEpMtrLS85am+Kaxa
N3tku06J6EiDD/8CZ1n9E+Kwdmc00spjecQBg9s1SSN37bP4PAegUsi+gtXY
NGQrF4xP/MjnRoudihW9QzG6MY9y5jNK5Z1Pb+bEKZppXt8OIkqMVDEDxLoD
pHw3I3XfdO2JC8KRUmgbHcDTPwwB1IfqPmY3gWURFHZN8jDZD8hHDV2CDRMN
sxsYzDlroppCqU8/FatQxDpUItxDzDiWsbEWNnsZsVln5Nh4zu0u0bio5ixG
5R/lJGuAuII1R0ba2uORVQsrgMzOvSNLkqsjpbNXJNUeNFsEbwbuB3E1mK2N
vPurXc3g9hDOOkKRDfb0dwsrMWtp7+QwVQH8Q9RVflZBGmBFoAOBKIsGU9xN
B7VkzS4C540pdLCQ6gJGVvO3AUEqv5ZR0hthbJCWpENv9zSz9fj1v/tZozMF
TNW499HA2h9KP1IxSM4nPWz+gI+IEaF/Qng9eoT2k3KbBfbXcRMvL937YYrD
XuQfPbNky2/jMtOhX/dba1LnhiUbj4yDEr2ZKQBsbXb4Cs7oOafY/kMIlnyA
hBt8rofdWtqFv5Tc1JISOL0ZV0VGoA18wctcQcacIhfyc6CsRRXDQBSt4Pfu
zZgU+nTKUUAUj1vV65NfPhGu0Q62mUvGCJSry+TMxlvEwaxGTCo8O7Dtv8f/
Xe7qsuD9qOHdnQnzLpZTzClRTnQI7rtmXidZR1BwCW7aG5gqph329FxUiMdZ
TCWvLec4VSmG/FceTgktgDhXvykTftdMT90MSpKP3gpCshfE5ro/aOXvkcZ+
Ypl3D/NoCtAiEibIEt/MP9S+arNIRqRiOoP9LInJ2fxWuF+2TWUMiZZXOhET
DnPOyst15Y0NzIO0OYU3ZOtBYnWTSFEhArmosmaf7RoHeleCOFwvMqtGsLVM
LUUYEZYoQ5ThpgJLDzY0gJlwEn2OTLzZ8Mf58rcdnbZcrWrgUE5oHOUK/7u+
nYr6/uzfv9MZ9mcoLnxszNlvrUTMtLemb9U7mIGhJYnLsuXbHJETESASuUbW
HdkIrXAlWv7zjParZ49oTkt5ms+ow1Lsj+5+6qs8AxqCTTJTCYYlFmLWpJZg
rWbLTSJXBpOLPJ97qB75y3Pk11AqmQRZLX7dh8Ps1iw+DG16c15BDJdykFe8
y2WNiPhLirdnxcc4I9yRyyeSPBJ1tsbwVctPz2zrvtVGZ+V/ibWUUo8egdcH
47u+jlMqvihnt3K1RYPtQHaVzkbq0CEVUbb05nXfTN+U/YKVStVY3yECEXF1
aqe2vX0LHyHtACqTBKfojZ7svgs8JvkXvjh3GINKVwxXA7qzjhHsOXiajn8O
jk6NuwGTWHnTj3UwmfhTRYxCSutfjUu7nJDgCC3qM/a84I1tF0dT3H3eCfVL
CV746R2L/nSOlpPpAGGFvyOREEr4cPgz5w3k1jiQeKVEwnFzFWKx11yFChcQ
rqAept+4fFLYDOVeWAcouTNzIFilSKc80jv5ZPoxqNPikXHjLXSJczso6WUA
vwsOGQD6ag+oO3J+0KJ/7F8ZjhjM9tyLsEc8m3Yyu4uaBpqI9CXYKuPK6NrZ
IYGEhpYOwu1AoUAefRryxEtb5NGEflSZOMT9X6SIsm8K4zyzC4ufPoxnerYZ
jwMQyBaplpkoHVcYc19zRhpgzoF9Ukj7KrKVbAMaNabjaVlUHDgxBCu6qPiZ
2UNKNFROakHsd5vkB75sU0YkOw08PWMpGgSB56xCxChaJbygFTcuamBGN4/z
muRI3N+gumDexBGvkJlz0Baf/nY2GadpN2ZTkbY66JKaHbVyhOpReoBBce7k
0ba2HHmQg2zzjhFG0hkLr5Je5RFAnEN4iSyNh1YWlFyqL44SvbTsUDtEDodV
xJoITozcTGSiyM4rkSShiOvfBBzta+hzfX8vC5XW/0ZzM0eGFtbkcN1jlRPf
Aviesx08eqP9jQxSsbr9yADVUrPqoyZTuu6YYDHJk1Sblpog5QJ8faZTOVFO
tVsyGuTHTKdhxFhk0zUwMCqO1MC7NN6JKZQRjkFzZOpxax+K+uIfPTfXqmaC
G3+7gp3jEmqreM1qIV3ZppTvYZjvVCmTUBiDgNmncistOjJWnAZSbbwStKQU
46GsjCL7zusbRTYkZ06zBHWJe89V2i9S9zv5BRYJI/I0S8b2xvhaElOlAnNm
c7EwHykUNddug4QfpdXayoYmq7bTxbuYfyInPo8l3a31cXM4HaqDFfJ3rbpM
pL5fZbCZqBA7qY38gQoA7llXxQdofRUnJepv1h7gRZf/Gue/a05S8kMK98ao
ezhXynveL1hfSMH+XAv6URY2m3Mr3foog/sQnopeYgj5XONDLgd2umi0uYev
EHTaXmtXPMQOhnsXHOjdrzKbnp7nfe1/K6Zgepy8XWNSXWbWTLbG3IJ49Hk3
GS2ahubAZ7Ws1EKcnI5701mwjuPtmlBH0dPQllxVUH1Bnud0BBDhY2XvYK8/
MtR43hqmyP/XLQuPkUyIF3ey2dbj7hGjL/KvDfXBCxX/tR7gy9PiWuC7w9a4
Hg8oV07EBoY6iBZR8wELf37Wc1fY0VyOj3axIoJ0Du+zPEQwWqBFO8yT//WZ
QSjSXSU+G/bY2MRbj8RUJTXHjfZxvgLsTY06eQHYO/sphbIUfrBYPSysRVYn
rniSOKaTrk/ar+U/Tp1YB8s7GkZCLINKGsqiMh02b1DtiYKJ5hVWxfg/8LS8
VNB5dCYKnaTS4FM6SQhV8/2XNpijzRVw26c8t9E8G/ELg4cYRyTtOMZHi/ty
VlEFHNKXn9mcxqeMKmopPvg+fojIG9SRwj8RZk0/mC/zipSrDuCdrfH2GiKH
MgRszlM6RGPUJRBWvQEBPVCf098TTQWt91QpZMkAAofeRNTzIfLHhJeAh2hW
UzP1TjU0Ud3BFid0VgZYipA1NWVGJu5V5aKhF4JMS9U8A3i97CwuWiBZY7H3
CinsZImJqbd/ftkGDqS8/StGHsjRFvVsXbvC0WWuuAilGiNdsthUeVhO6KP2
yXKH+Ip7tNvvIGEiYFjTexdEC0LpDH6vN6M0JtGId+9guIc0bg7I8DbD7vIf
UN3vvT8xAwL3FBq4MrhWU7aygASMvqX9DEAtWD2PI/CstrsmcBjxpHodvkdz
/Whgg4nAhgnTkiGo6idOVFJrKBBVDRwKILdtbspJRQDpVBgYAhbVq3jvWOpF
pPTeJS7MOWnIBCuBqY97PXMyb6XniOilG3FR3ICK4phusfp4/PssxnRQdp6+
rHsKE1u0Ob4BsAJpD6XpJrNgllgGSZqGhPyONahWLwat/t08FgsH9o20ao8B
2t6NjB0DnIvfc4vdmVqktyptE4/B9kAxL/PfEhGOhqhjIfE1jMl5ulWJoQN9
fkA/LwP38GS3jS4hUKxNDNI7WBOgcqjOyzirIQX6ji+r1IUDRJvUynVCMd/X
9zaloaML2V3OS+6/pIoAfy/kDj7Y/7gH8CFTpwecSwf6UFQy9xidFyUsAmgn
mA/QvCGhZ7PMYY18zNCz2hw6yAE84MjMYy0BdBd6ZuWqS/bag1aw/3815F9H
WIQ7vS5+Wmx/NFntIWDTH8G5kH0ntz5A3yYFtafuLunUrn7+09g39R00hlDL
Skw4DAcOvfUeRu5T2ZpqgELCTrk2ILNDDK5ytFTsoyxKjd9WfjoqgRrNrUk/
1a+mrHJZKiKUF2Eq83qOJuRcv2Ir95ZTUweYYMShU2knd4FZRfj0k+JrFYot
w5bgacHF0bIuV/EYScOcPuRO3h/xVVJf0sdWo1l27pr3RZhr/q+3iW8tcY27
NtuSUmbMt0BvBsPVrkqsUv1pw4ljEoKo8SipIqzVJSnjJ52gIT9enHPWxiWK
EntIFZzCHQRWRrZRwGAYhd3/274oOdjUhUpWV0IrLiVAalm6Cy+VszdrB57r
CUg9RkcZucC3pZJswhn6UCRIULh4AeBDlIIQ5w4pJIsJVqhituy8o9utxnGP
rGchT+c6knSYkKBoCR3UED+yPNDb1GrUyuJC5h+HUWCag4sZQTTSn9IJ+B9e
hORRVXtXpSSfDDG79Sigdot4pCtg6Ioc0JGVwzPcDF/DKzm5sDtVyzHqE0YE
L8SSR13kmaZeQBiyYmbT46xjCZUXZD8szl1jUC5eWt8GGIvKjgjOHXgvj0U7
gYUrX8DB7KXUhHJ5agrsyPRxh34Q1bL20apRNjUiqHxXcve3vGhU994T/Oqc
kZLxI56mvMCenYSHBOGeAf1SOGeLALYsNj6GHGl3o775j2jv8s+SW4VwGwz2
vclOUwqpupRjrkLWM3j0WfFYvj/mD4W+VlrBW5sjerFkrj5t7exJvHw64bNk
aTrnwP75tW9DWb96C5ppbz5jPv4lDOYpQx/SOHfRsWOyUf7hlRoRHO1nTawo
Gejsuk90ggYydE8OwnO/gG2yqX5ei0V2fU9KmGlj9sa+5oDoYFtxj3ndvgaM
D4TIlJYgUuGobgsQ3OyQBmhoA0MbSemyK1cinB3unJpDkqqQsg0covLvRP8p
e1a0qO/T6cTGg4eoAaJc4X0wdZbdv7FliU2ie2CkPgAJMHc0gNkAcK4SC0Gw
yS6Z5KMGWkkYXOXkwuQ4bo1P62CrL8NZM5hIO7h24E3Qija1JcigmpplPMhq
7IdJKdJuZsXLT4Xj7PTy8psV+VAEMF72wGehDNxgBW8KwgF6/kHzY1KBtrjJ
lKSkIXdd4q2EmiLGFIjyqDCydg95Rf5LWm03ZJZgXSw+hG9aMNl7m1uiUSei
QLTEHBcvKaloyfHux6jEuF1aj1a3WYtTmN4+tW2bsr39sShYpWf7MaoFEdPt
jjDOqC6M9H+9qchCSnvJ/ZjkZ66AmUERSQ39MhQnOyNoHBWeIa5N2jZF40Qd
laZeRnlYWedrUGFZIc8A3rZ2MooFoM1fhO1LAfVV5XRMdhWs4uvmVJpU7WzV
EeGr2qwLMJTbv2YCNAs4dpqdH1Xu0PeN0hJuc9xrKY0xYdHDJ89C1nWF+BPK
495ZgQUG7N93laxns3e5y9enab9eABzWRCnwlcYM6/tZbmrNF3WqkzAN+Aua
6tQMc0aU3E7Zv+e70RObCWRoZWltZ+rhM/+6T7rR/EZvjOrjPco+OElvKzFn
XDeCHP2X/eRv0L9eSQ1TnAPi4NnQqlYh8oLtgmODlHlko+dNLJppYtQqF1wz
mLlltaevucMgT2Ymri/dIz2NwkSj4m4YZG/zvvtArtZ5okntj/1N7MZR5COr
OGz+7gR9WhTmuVW4pdDsiXq1bXw9Ldv02z4aFneFWi183ZS1USYRrwTaJEgW
7vzTxOj71e7daEePsFhxRcgPaWbJgVTGJj2jEutdWzgqI5rzfNbvb873fFX+
16GDF96zLbE9zQwSC7pqdQ98pzOxJIX92wviWvWV8L9+cMh8IWpJVEJ4hd/u
Xns21RFmldL7CsHkyNxF1wNiMXcmLNz+RBFHqA1x2ESrXaSFBW/Te2s/y0qi
JF8o6kVj75Vd1IWtG1qyFEt1KMH0CaamQnq/ijfFC/1qibThqbPbOQNO0CQ9
2wHz43ANsQuXJk5rxF3DbNB9je1tLJsQApEeZNghtz4MbGWHtprUP3k7TTAo
lOvU6GbmbVt5+RSVQh5sWbMeK585b54evLDZubcPrFeaZhEGqNFlywk5YVpY
+RxPW5iw16Yl6cNP5EzVDS+RW588YYmk0JVODODRCvwlqKCj7m9f54xC0YpR
S0nPYr+RpYdVQ2LU+Coxyt38Xv+mPCyvvCnCYDbtQGa6A4BMImV68SHBJhs/
FZZRtxeWvdQSt17v4UPr/ajn3nNEuMDCgNj3oeDWqBkWl2nBclxgLWW96sx6
6JbwLFDVsT0BPM5yZuOpd0gByHKQkI+YCJBwMT0Hdf4rCGLad8weAm4vCk/Y
HOkCzGRx/4TadntlTDvcsEtrvQeRtisvqYaVEQ1DTyf8Dr2T+mVKuwZo124M
NOBIyS2p/WLgV24qrnxL8rVVAppQwtY0Thi8QepVsVzk6JVgWFJK0gZXPpE7
xU/b331zHXdIUQLzCQrVhPyc3pSp7Z7FAcAGQstQTlduIbFx6YvjHCdkjSh6
R5KzQYsxe16YezcGjwuZCOWC2ceIQawk5hMsCgV0XwzepP0brlZzNQoLf17w
w1S2kTGppscnHy5YSPvcGjzcKtrYwQ0/ZlyRnFidrhDq47PHGqv4tFpnjPFa
LoaFSewqSx4clpPMamSZD/v8z94GH9N5ZUScHEGSyuXOQ/Dvx0YOn00RCyk7
74IleSKYRHwrDoWc9FNhMF7jjMyce3raydWWAxAq3mIYMQArkh5StH1FBHRH
yaEGJuwCyyIogEyEDC7VCFMd4aYcb3SXsqqC1ySIhld5LRML/TJA+I7zvY5f
FqaUIzlz2gzbzbbbZWDW7fdw7ElvyG98OCBimpPMcywYktApheirkeJYiDna
WFY7GJray0bIP1cEKW4BCs4p6PyPHM3+re7J7idhlsYGLv+EGLL8PzdzVXcN
vkJ3nEYbpa/lEzOTQGxuyjliDKCfBv0UEqgUviImzV++AQCX9ELk4See66tS
hCmef4LeMTHYBwplMJBvIRPaWCrrBR9K+SsMN7U7ANsfB66LQyLoRuo7IOSl
0pffaV3TFaw8O9eZUj2+sfrLo81DwSrth2mLrpwClam4ZJVSLrBwX6MikhfM
f4Bm1x1rHazaK/ljJJ3hwuHU23f+7qkCZSum36ut+1iAM5RnKDUUicwo00sq
gI2bxImV5pwyTsy3uAXLY+8n2fD2yr/QvfLv91x7oB7PERWYVWke8JXtmxQv
z11sLrcnij2tQeLBcRwjYi8Fut9dGKhjBDflmaS7jrclCHTS7aIl984giL51
aK5hTZuAhKEJcvkQ10GAkCaoarZoAXbekqk/8r+GZGvHLEBFx+sFzva7i0G+
UqDom3GazLKbEzGZpBN+4qTaotcXqGGkkffHbOHpA3T4wv9jp2CgqsLw3/FV
bAXH1t03cRYOGZfW0PDErcbzZ0S2ftpaecoOWlrJmRNUIDachxg+aH4LvkHH
EHotKbeeBVPNOjK+uiXYn9zDc2AGYqENRIcjlp19VFXZWmr/RCyBHud96Zar
zhWsGvdURTpWYlhW80cqYQ4up9SPBTX6jU0qHl3CTJz1Vxqlw2Kbcz+knDY1
MB2QPuYmZ1arxbwaVth0OzcR6YBpjlS094qa4eiRQXTk1IWxtP8+SSTQvzTZ
Os9g1BHkVLga9MqPP8/10vZ9l2LetovxCyVNbcFlN89ZdASSJT8Sza5UsZ3M
iTo+nX0Cu2pzpI+0fsHUxLq5eIj7mxEieqCLD2NwlHkz+Wu9gVoLi5TMitge
Vt92NxZ5vR59n+doYSFerBhWNDy3e1ZBikQEIPW8YCZ+RQtXpNhhe4To3rBC
U5omzTxDV2uiv9vhPSQ3EAxcLWla275ejXcOYKzDDSf7IP0d/anHCtcgv8gD
t5B0fvFuANjweQ91f3RjLamlSLKfaHFd3kP/Nqt7vB+lB6AEwgX7C74i4M8s
E/qfoBpHKR2cR+hPAojs9wUkwN9Sayx1qzxn9+eohMUZzeu4fH5dEKZksd7o
6gFCuXXOSgEtPAbaLEqkjU6EBWLbvxVZ0wvv01mWu5pqazCPvz3luXe5NwbL
zXGkHiCObpVbodoR7pNpo+NtCYwuq2b8Xf2mY29wc1Wp+4KPZoY9frqxHfln
JZj2miRYhdMibWGE2M2XVvOV4nWv11XK71aX6wvZnps5TafF73I1TI0VvyIo
C5fMWuvavs0D4WWVekLxZgD+diUEdAObqdj+yUodCZLGppBM+ljD5BkuXFUi
VFqcTtn49T14NViVzKtpxMny6qE4zWY1aFPiC9Y1mv4mXi6+HwMFVUXW4c2q
32rgRWFVY5MtWo0DUKFnHENXhvTiK4rUl0a/6tSBmmtRUpD5gR9N3Ru8nyDu
Uwh09RQrU1a7zkwyZVaXRVEQHvGisK53sNXAdR1vxR9siOI3F4B5wXaO0nyz
eQRQTssJeWTaFSoVRfjqoXLvoyvV3iOuVXXhBt5LTFL4svqv5kWHrhlyZ7Iy
H/r8V0fBbEUw0g2XfXACksJfQDZLVGZt6FprR8yiwYgqjkFcyxLHpRv2rpgP
Kk7Jl+o/OGOTHiFZYZyqDeD4yAcWJtiOKNEbUBXMcycGxfAK5kfroakO9eQA
iPOqzXutzgdJrQEdDru/8gKq2l8eaWxsko38DmN/VbgxX9CHNKBa7+BRb1Zk
O1yOHlQ0wuvtIY08Lk2OUSxOhOBAXulq9RwkKbkFHOE81dnaj85Jxvm/z2wa
JSo0s3Bc6Zqxi5Rccjy1OsW1LBOZP9cTaSvlS0YFoy+CHv9qF4bC6OJ1x63+
C6K0ckREdIJscTJSCbUtSb1dtCQMJAUa51oPO6bEgPvNFxjPO8ghO27qBZm8
8A6ZFTWqzPcMAAbWxDOtTJKlqjFA1sLm2NoMjTqRwfe6o8OltPnwc2VvCGFG
whZIq1PZjRymc3Wc/8Xnx5nMVZEdV3uICUspciQ+SF8IkzGG1kfzT9Pxv/yX
vFcQc2ph1R4wZMnE9u1M6BHNCx1qNXR7Z8Koeu9oQr1expK5oJOfCHSxxHA5
8DxfpqqPwdQydPUBpCKLyFVDbUIbwbR0F9dNlWgaS3qG26OVl4IC6aZ7rTKX
i+uQhG1xi/F6JKFu2nbToXz4cf2ywohOZ1h19kyOpXQ2WgmEAxekflwPa9AS
qeqJMnVma3562Zq0OyT1TbB+D18QsbKZQ3OWhuZWAmwm7NG2UgCpbUWNuzTm
wSbLTAvvGuTVKuP3jszaKogyHzzsCtD0rAHeUZuAU3H3y7q8tfcozc0HAWhU
zbKh5rtXThj4P9/Fz4xLJ3nue1Hag8mjK0hrLzYcbukYjeP6AQq1Z/c3XiOZ
n1Go4FNkovlU/vpixnLem7VOotnoQH6iXnB+M4U6uDsdAlcF4qPC1bnOtBY8
xHO8lnB0RxiaPoVMfVMzAfIML6DPeioS6Dug+UUn8B/Um+d8zviIHmaKv5hD
ZuMHnGM/QBKWbCSOFNMzYq8Co74NzLFqz65+CNvTAoXccodkNNKWD94msoZ3
8l2M1uBWvFZ7rHOEdfrfJWT1dCuC+x+4WkfGB4iK0LNYIqXxVCOBMpB4w3LW
fYrU3xbm7Lx3pINs87Jq/YfhJKBsLor/UWhQsR0NyV5e0igMHjllnf3bDUxg
VC4gSnbCxcC9P99D7nTONge7FFcfEJBWJeVcP4WBBuWYE/OZp5jW0eKw77vb
MWi3eQXzVp9yC6OzKgaIt4sLuoU98mHgLElUwwSv0mXtrT2VZNsYDrotA4ip
Ns1kgEQAm+KFcII/DG5J73CY5HCQsCVv3rkHQyXmYg9CsA3VBcHPOyV5cqcC
sz5esvtPXwkC6c5QHF3QHp0+5qO4xcNJz28nSI+o1p49DEK+j4v42f3j1M80
Fq/ukj2Pg5/vBNdRNW8dCkmMYAzEevMKxIV5ptbV3Cx22piO4Vc7l44Y3E3M
VhjZBdyHvCYLpemGW+HlEK6D6uYeM6avkGrJwK2tfKmS7vOIPt8fUHqE0fqC
ipmpVD+FFZ9TxP9mxAd03W77nz6M7n1QPbG5Rh4EWtAvKrarGIDwqToWlonF
UoqzW/SDMdAaNdpc+Q/5c/2UjGlrZg1GZSoH4w2szyFFtN5j3v5xEc87XXN6
jyK4rfOjsBqp6z0AVBYYty4FNxMNJf72inBqyYnLqlvkphNeffeswy2xk9ex
2tbk7vCy8zUgy5cmWVihzibFr5D9TqR+iSvhoXMICb9A+DGmTUaYn83NJrw/
5YhZJrx/2lXf/gpFoi+Np3mWgwI5DYA5+DL5fI+pCyYrO5WtN3Uf5Cm+Vgh9
MgtwLaxn2gjzLj/TKOd4guZYrEz1vIRdV+J7Xjx4go2vFJZvFXwVePDWUfOS
n4HG6FZ7K65Ghu7KCY/nUo2E+8ZMBGWPlA+2qLi/e/UH/oW7q9AV0T1rmYou
5eQF9nWwQhdal3Cj6MPQ+0kmxqJ6oXAhUhgvI0bRmof4yemRtqS7p2LztBnW
uun8Z5QnahvK8jA8BpkprDiUpFQxGza+KU/r1JXc+0luOLK0gPh8vfCTVZJm
OjpnFAHtdfzlEmxureSuf6p1Ght0YxCS//TiBKCSHW00gGRZq28MOhMfjDK0
lGxqRYpVjjN4v7lEtjDG9IzJ2xnThnJqIpjP/hc6+gZ9uuS5P8WwGkUuphV5
N2AikvEwddJZWSi6hr59bQrQs/JhyiYmpETSL/VJDxmjhK8bO5vzamGyfPdL
K5HbvFX19k3snWe7rOZR4dteCvGGHIFJ8XAPCxvkpJ2+QhImJUsnR/35TChB
Z2Nlp53RfwJC6+R5DaVkx7nrrX7554Clivft9kf7NZwqdVXRFaM+gjePDg66
1pn8+HFrjxZ/RIAwJXbPIrzJKbF9LLWvXu8QAtYxqlZCqcfMLyJezF4PHIMz
/MxSm4mY1/dYNHVNATPGOOBV3G+zyqeYP4iYW0Kzy//VJ8sHs7nncgQewm2a
55EwCv0jkRgTGgh2gV8h+hGQiZg++DI6QQiWDHAFosVpzKQ0qiQtME3CGFNp
8J7SvSnA9wUv0pt48wdx4+JNnoQtDIRq8L7Dq8UWCA21RUg37W0T2TCzhEdY
8mMpAmPzoURRjrWPlqss5pE660gb4txHvxM5KbtZtRFeI4JzC4Kx1hnn1vii
kuVYFSdQjYECcWOolcOZJf8JiSx1/nHmPdoksywG+GFzICajFzGqSR/HEy8I
47jNTKJwBVSgpHxmA5J0wCwcMLDrriodX4G6uAou+Vv/k1QTb5AdaFWuHhl5
I17Rmkzd+pHskkX/2tdph9KHTABS6VNLQiH2UtwmX/puf2nHCFmbKAb0Y5XK
8ou6sQzu9Bo/bRTWK47MoIA5qpYBq3mRSxbfaWqbv2X1BSpHTQx8t6hrrv0B
sny26jtncp7trSYku/Qv9W0m53AQvzvcWemWI3eXMhecAkDfsKDh3OvOzlzY
SxJsUFEps3Hes3C6WB2bUEL/nCRXUy5bGDaObBDhMOjB9HIhTJpwFjgbjpq8
ir+REIzUav0TrAw8DFEizVekCpgKAKNh8LEjGnJH2TJ+7XvCnMd0vuqmIpAA
G6kLHvrFZAjejWE9MuMcsDbSSE7X38jgSuPKSOR2sQ22ZVfZQgHasJkdoeQ6
yb3Vh9SonA7TwpxaSlizeE5iDVjFlEBloBKKgOVPHgBstm6XVAjGQj4aMkEw
6iTXlmzA0k/9Xkyx1o3rOr2vo4R5NMpEP+xrANrMQI0pPGHp/zpTTHhQHPwc
22sX9Gb7f80MgClyeJCohC6sA/rH9y+q/R4w8pbdGjxi67Jb/6UlkR8bD2Kt
KU5iLPsf011RglPWjid1mOaZ3e62yS+VxZHErsaY9i9hPbvs6zfi5Eee8D0g
6oNNlIm4oNcQO1rsyardCRyzMsx5ed50hqY/d8oWpaGsewkqyTMFoh1xBjhk
zYFMHfooo01Xnt/bTsEFJ5JbXC6Lav5W5H8fr5cU9jLcnJ/uRtXN+Nm7v55Z
Z172vQHstW/SRnSXB3dVOiGQY9qO4LbQ3MwkQ6NiI4mPHe4A9WJz2eGcauEg
UL/KJzqHwb3+NHbGnkfbaX+nHF//ocTzhck3EgBFtnmxAb1lmG+63f2MFtX2
6Le0uBiKTNhE5dl9Xrpv7BTol4zW+YDfLzuHUSwe+/2iLbp4Q4qQI0mb02UL
4b1dEg3H67Cd5UiTxgBbxxexv4cYseucuhH6FEQtwhw4QXVo3kGLPIo17L7c
rpNXzpSkD4weRRXlXbawn4nq7r1TogrMrYdTbyT8wlWFnwHWedr5WYnIXT0J
6JR3nKs0SsKZqH8T70GNPDvzpVOA2lgOVI5jD0E521L8YL7nFMZHAgx9Dwzv
zMJ9C8GbwriccBPrmUuz5qYF66TCuaUAtOWPy0cJTxtQd6N6f7dl6TKN8XL4
n8r4kyjXeqx9T0udQhj1W5NuZNIT2/0A2Uc6F9KphbwPwHDVzR67Ly7fehKF
yBDkGcj8H5zsb62x8/hmNxnJNYRTRmTx5FUnY71l7s89TZIdTgy6X/eoTUsQ
0jsnHy6N5ktQQeqPzMsiVjuzNz+BNxdnJtdwLcj3jaQQjVd6CTDB/7qTV99P
yLt3ncxGFjLuqP+yiMI3QZJfyP8spB/SEhqavFTOSsQexDqs0Bt30UESKfX4
x2O5bl+WlA8WtRKuv9CYw10t/nV/6rKkaNeX7BzieqRjvUPACJP3Gs14bRNq
/IGFgmZD6TKROd4cO8i8J8/yOBOCJy9/zgGQHcdunLapGc0gV9JnWqt6EMAE
vrPczk7quHf5iuosRvrMh2mtopy4xJCdIosLFTM1+PUgphv6i6hVXFG22nON
nDou10V8NuqVAc3YVmJM2Ps0B6iKDd7KjYnzfzf5lb9vgYaxshlL402m2RAS
AQklFc98tg9lHMZ887Q+UpSDRAU4FUi1rQOdf9twg69r4D2zwbA3Tm7lQxK2
HVg704dZEfkEAshT6+JgQMA8yXstHwJC9o+1ChmLlXkY/gqRBV18dmp9IHj9
cQZoeenG8E7BTZ/kl3XF4IKxmqvk2DtJ+v0Gdh1oP/N1aeC/984+StXp/yTN
9EOLHxcoiQ2DGdz3cmB2byG/9LNa4eh0J+9S4zfESnHKzct9Wpjl9dxXURWk
A+4VsaszlwCiktTh8K1gjYz2h+ftCWDPvnq0dGbGpnXV4PUNykYAlnoDShhT
9c2eANkXktog7eiylgCC5oXcePVo4Qqt/cJyiXcjShH6JVUOUfQ+fxZM2SwK
GExW1z/v7VG22vmY0ibZDx9inwLeA1MFb+Ii4b94JbILCuXENwzngbxd6pr5
91D3tw7PgA1Cu3wRWgvI4UwrbRHJfzEmmLHmtC/P694N0sy18S+Kf4f1Te5n
rb8bF47FDbpz7WPN6N5XrBlfh3bvpAlu/wGB5mOSC9sitY0XCB0SgIjAws34
7iFQANA4fyBmysNscXTMRHk903fAt0LOnstDkl1qwwestPPHHEQQl7hM9Dnc
Aq9wiSzyMDCBfrtMIE41y9Fbb2GDYodjlPCmg7S3hZKbr4Iitx7ouamLoxyZ
nnPP46k36Hneg8C1B136tISYYWL05degwoQXzZBRCDZF3kSo7hGf8UEtKtYJ
8M4pVeO2Xx5OXAOQwypRwNtC4bAnOxvVJCIQnXe+MxYZu/SVEbCuG4AqfAEQ
OmTXNO2mj8DvfBSjNgRNUtBdrr3KxvpG3Qs6btqltnHGlju4hQd5xvPuHLJZ
bqdkkEDuDdTSY83ad+CGf/MkMngjBGCttiToIiiiOJ7aT34RODZdP8HcaHlp
quENPrYKad88eKhoe7d2a80NFhT64LU+1Su5tv+dtWki+wUny2Hp8VEsT8LU
L74YxJKwV/tmM5BhjXSY9cR7Akq7XuINlHa5jd9f5b3zqdnbVpTg/Zpo/BYp
AzfvzgiyvpwnmO+LSD5lXVTMyyBN1511cNtY3MXH+/Jl+ZPgS5xcUCyBWA5s
IlBdSwO7KemVId355cXgzUlvcZUpNEaG4PW0NZRunhI61M+JIJwVU/2fRFqS
jDMSu60JsykCQmYYyVMLtDWoD5eG+GbcuGVcS/mtMb57n33MjzSA1CwhvXXY
mj0ijnHWlYk+yd/OtVJE/zSf4sPfReLcWbJBHAsLc5fR0FRsrPhVGvneEbNG
UDJHT5DI2iuxamS15wGL1O4cFiJrxifNn2weyf8Tlym46ko/iS4cwREnMcRB
Shv/29KYcKSsdiDnMOwVmPEZop8aBaCGG2peP96M3GvCG522uiYNSKiJxXka
u7IfEQvwrhlxApuNmyAXEbnZmkGc5WMm1otKuI/2mflSHINyTz2hFZa+I00L
V9thskXUV8FZzRNcmhB66K0aypTm4scLkvQ2htUUAngOJrGklVNfymPvxDFq
tRe8A7k/JZd206DnTC4IFROOtwM3I3MRilwtWiKN+xdorowqvuQnKaeNAEap
HX3+y3uD0inZPThpU2fhr/CZso+ILZAQljvF2cGatQjTIR0aJ/FWEo3QreE1
2ngq9jDCr08qTLsGk3nqvpv3EiymR/Qvp0MKhESFxm2TDymQSCm0ndPRj85i
pw5y8uBaWk/nIbRuD6tNOOXyaXW7J/gYptbTVP+kVFTFtIJpaE7gave+4vt0
9LkP1qz7gJwqdwpzZWpotnNGayU5lbV0zO8p47YoSy6IC9ZoM43+nn6/8QMz
5WEi6DoZdXBQyFCgtl5YVvCtO9bSeHhKwi1CRMvfXRo/EGF9eSwowI89H9IY
TyMYjjhKEMSIunC9pkmDBx7no65TQcg5DdVP+cT3+pO+xliaAGruA+JfnJvB
O3N0G/GI5HABHbYkf/jjhcDhiYXUKDya0C8mFio95Apdvfzcy6VIuu4Cqq36
kHpk3c6T2Waj8wuBwQcvIFUiEKM88q8XvffQSqcmScyfQoy9DHM0uvWOTZhJ
IsdGSe5r3U1IWFw0oqIcfioOMsHZqoQcNguS3fP99DkmDy2BtYhHhXZCTO3J
BG4NzVVUDI4p63myMeeCEsAhSskKy81uRVeT/BExPxKRXdWmpn0MDtwYScW3
QNqXENFW3w4q3DVabV8Clc5EpT5FhoA+v8YyXoM5SNZdyj6AGOkU5je/7SXB
bR/Ej+SjGgGmI1nn9OVCfMiuMjYaVNbBaMb3ErbC0ReMu+wzu6KMBaQjSXIH
vqzAvumfk2UqLd9X3dlyBkdV0OlyCnPPrTgzBr2O9yTms5dphUGyAissdW9O
h7Lr/OcwujtAl2h0bp2T/0i4aBO7XSD8AD/PSaolkrfIuoGvB6/J6TOKQqCQ
2pa6+NaEH6c5EHcOfCa7oNYDcbJq1WXEmkx0Bqy2FxlA7oADmg7O8xCp7o2O
jzij34ajUrFZzTd5Q7PWQ4cRr6MnADhozewdPvC8Vso8kso4aC2vk5PYStqU
H1DbS9LjccdtGFSr1OoL458uTx6AWXol/nLa4VTtzta4YDBAwmqio421xrwD
e+qdfaz6vqAjP+bc60FFnG6dBcPiU2uJlgZmdie21ieIZ2ho5LbVxdq0SWLk
lVouRoTmMQjWh/1bKpuOeL28PzfqX3ZgQbnBVf0hZ1uMcGqD0AK35kvaTd3E
6itxVeYiYec9Gse1fkeHLB+LHlg002vtPG5WcRDlPCdji/bS+qifmnzKYEhl
UbhrRAn3rWNEqXpfviX4YghG2T42KAaM9pjySNEwrap6x+3WaWYMXV4FhzAN
kYxNfGQEXnaq7lxJx/CTIdETyWEiTm5kzwAXBXv2UxMP/+oxIrmHMRgL93Ca
JrGt4nhDyT+uUQXVSXZh78OLnIBon9z+VxXGL/ScmmVC+Q4DGzFR2jbjMDeG
pQpqWKsDEb4ky0hSNtSY3clKV3mUqPJG6oLLuSUmp245S8Yy+A9r99SFiZkk
OHchMBlygBygtB8IUz+SRK2YBwCDFup4mnTONRByIu8YJNbVLhb50XY+U03g
ZFoT+93bVtk4byL8zi+C6lCRwyuOlBhUJbm3t2xK1USDrlpqRM4wVkkiUs3G
0bha39x2yvtBXbZoctNvCl/RJS+5KTz09ng7FVaFCAShGRkjiI0dy76fTdiC
iRLpSbnJ5As7Xt7JHC81ibz7Uyk4t1gsXSZNZ386P8T69CT7GcOGxFDRwSxU
4Lob2lFIGHJnomRsD55upKioaF41nP2/HLMX0CwhR0JL2Qiklbu0OSxzQA4Z
2skimSgLuiRhRDkRTBSrulQzV/jk36GCebMcqy9Li4DOSnrrORzbxptAP8GB
oZEAnib2Fj+SC0a2XAoEL0ED/YfliRFA1fNTBYxPcgq0diSZb6rKaXF0aTd1
v/dXpLhUPBn/rWwKBrCmF4nPDQXEdFKVFMjPj0nIwNaW00NUdq3zodZtO4og
GLJMBHUCvB2dNfSM1R1eYzmA2OtBR+j/Wd9qsU4hrwwdL6/+EdDc6TirmbGm
+LjYsufVRNrPVs+ANmlU/e4AauTSXKhY3y3opbbx7UVT56hJoX25P1okyjKl
bHHxlr3s5WkRd68lKvsbW8TlQbxeY5iXWfKvjEDxfee7Wq7qV0/tidYUvguj
RqDfHA8cQN3LSvIaTp0W404sdk+VzyIiqv23eLWXiaFUUvsxLou7f5ZHdDYK
ZH7DYo/EDOqKpzRni+9L+ADBlngXMhupPnmFsCmHnLOZpljz1febJffLQ8mI
s07EMfcFuCahM6mUMzQtXMi3oAt3MdsIfgXbW9zEknEoOSo2DX4/B1DiqWXI
ja1xB8hruEgqadHogajnCaakZJo33uJNr1vc9fnPbHWcGE2mo4DZaAgSKba7
7qYH+izlEgwS35cvt39114rgyu+8m+q4A37sg2b25ao9/vF2t5za9NDGNjP6
SrlUFxjefD2lXYd9q/UDID7Cxx7nXGQZ5nffCX2cKRL1pzje8ZH+7UBtmSP6
fM21+/m7S45Q9euR/elhwNjN8aaVKKwT6OxxB5sit8dZhkQROy/nmklLLMD/
Oufrny0QtF48BvS+Ir24A67sH8nQi8EG7ZVMyLfc/WNL4zq4VtFEEx/6ea85
/w4ckjuCBdG/J0I9TYjX5FaEFqQnnuEVQbM41M3BIdGnFNDWBzaSZHYK870i
BE2EW0oxbl+/0r9UzSp3ctpkyVbxUL/fPPRrBZ08DpQmQUX9Oe8Go6QHL2wR
Vpe82+++MeZ9i69xp5s/njJ37g2Ch8FLDMnsLd29C2wJ2mz7qI54sVYsc+HX
kb7RI21LKm2G/wfnuYKM/47xK4HfSFxxwSUY66mhoz38FEaRmpw/8J4nmpRc
BU25gbpvjKzlUyAFXbajJUT49YuG0yBO/XHQqEm0BRoMBl8DVfZiRQRFkz+p
xYDIyTZadu0jzZC7r5YO/o49qEMWRYxB+olZGQklIFQY4hTp+8fdnTb43XuB
9eH3sXq1jEGyPEF7mt1VnO/FkAIZrmwRj0UcAm6AP+pMn3HdplmAdG4DXEKN
ME4yRcN8lD99UEyoOWTrks+zDHFfZ+NxBLnOdx46qWAMGVAZan2pwvPXG7Jx
GLW79wqaI7SC35k8UargCO2P3sjl12SML4JJSxAOngobWGjtLFgSx1Rtgr79
j+dzefwPk+DCsBVV9FLY7YYCIS2Cmr5p3Plxv92mK98xl8NHP1FXgrWGhqxM
Ocd63jz3h+TM9pKdFpA+z0FKi3LeH1+WEX3Ch/2oK65rIIqFDUlFRKc6mupO
3X6WFP/V9jX4jKPgNshyRwweRSaTbvWsW6wRJCbdI27JnQfNJ38ykAnWIySB
mkFyQ0Xat8EWpFy8ohkyYhd0mf4pAATyUKL1FlLHnI4QjcDoes6byd2wiE48
VqhrEvwrD2jioNEJZbnxVzrlW0tfDL7PG0wMmSWcFa0vM9XXhOzqHBiOHF2Z
vMygGpeYLAzDFckLWXAhonMDfXgIDbFJudNC66e5OjnnbHEI0UY1Y3ntgyx1
y8fnkK3nUAVvF8/WhOp4rcQRoCDgXFNcs39WqyR4aveNlNAyTVhGVRuHrWbh
CGgUZLa3/XCgWeLVMxqn5yMTo8JOKGyP5LeEDsc/15IrJgwz90tVI6cTJHWN
Zih/8slVVb4i6Fd8P57jCmnYagU4JC6XISnoJGEQtOQq4VjpAPn+0wfbPybD
RND80S1/NWs8LJ3YFdybkzXun+OflO/FA/kjYYKKhllScNBtCNrn0myd/zK5
3G5G/l2PizLOYMATbP8QMYPdbiSghRQ5kXFMMRrHHeEuBoHqJbYpPYq0oQFi
xLKW/0ORNSuAR6Y//pEp6UrkSKiJxT4PBKDMMSL8Nxah+X3LnY1VhPvtAy62
LMwHWB+igGsF50Szsce/53I08XrdxOO6OjxLlAbAHh8vWSv4sPYRYQZY3S2z
E4VwGoevfMJ7agE2u/tE4oEEPW9DegWbG2npOxEp7kfaOmxzATccCrIuyaak
+OqU/LYI7hA892fF7H8u7VCsfCSfuVdPkfidTEaIuulwABBSqOsFbrV0pBZ7
y8541bI1Gvw8pCkpVhebiz9Wr4z2/bOuKrEcgHcXsmQwENhqWvUfHshpv2lI
v3rb3nuAn6yaNROVGPDb3b/emlMm+h2t0h3LeSB3mmEw3VR0nzr4dDu6urUk
RaAVE3/9miyoGphlQzDidsAdrziZ3I70/WgSEyc/Yvugnmm/BPqD2LLQhh4y
D+vztC8hgU53e6VVyxaVBxm/Z0SLtO4a0S0QQcrpUGljiwsV5nJeJjMUiKn2
Q0nyl5rx949+3by5qA5kaUNBljlEsaFnPaIqUHMeqGX79f9VxQhQ0vTU5kaJ
cVhB/Oo6jZf65oy+wLGikEiFVv1iwlAjcPvzqVj0wfU1fcjfWGM26wHEBQfq
AqX8BYPVUZsBz5quN8fXp64vqIas+VDNXChYQgEzy++Xlwotk/Omxv6dfHMx
BrHEXZj+MCCVM3UhrBnOcaG6TNlyg6vzbfluI2VNY3w0eSQSGmVKZTGn25pW
MFMlD45JGLFOAxCIo6rIQ+UR/s9jvPWQ9Js2M0G7NHUxdzJYKfrhJm5kx9yq
IIIFjuPJeX/OuuFcCKfwUGTGXHAu5I5KaAN5bKEmCJC8aomLBElNskQJWm1w
RMQeMVsNBxlW0FGQLPxy6hqmN1gh7z51uIz8riyAgqQkxBkVy3E4Zw2xQydy
6QZ7XB7FSu9vFB+DOPlVlc8MJxFnJsq156H4bAKyqTCSpI4s0iQqxvjw7RO6
Ii5dLxJbOmfbfKrfnTiPkjSkZZ/zCKAYKUbtqfloabjZa/zfaGRogTOko1mF
MDolWBSsBSE9nlvVjpcIgSP8rh+Tyop/W0FQymQ2KxgL4r3EBFKwjnF7alYe
eyTi01+Bk3z8yzd+fGWWvwD41oMburNCuxfSR0T1p2lVTuWa+/tDs+l2v9y2
vETN1Bcz+uOLEt5AaT9O3/2OaQClfDIg2wznxehRcelgCE3gSlqxRh8iguBw
ivnIO0JqGyZ2qpLdrqNK4bJhUPK3iugGKVh4hPXj6E9SrFYp+jPgthwovpbY
FTYXAeJroZkAOr2wdi7t/RSPqQkPei+SB1K8fQZYhWj+tNuuMOOHtWwEuz/I
/rQRM7QnEyz6UHwzoVHLK49FwR3xdvSHdbzgJC8oyiCjLz66qf0hiI/7KzT0
Ai/5rq2PmNKZrBF3G1KHcmHNI8eWk0x+NtgTAG4Jbg1+UEHUiqvSDKeD8lxa
SZnJ8foiZwTEGwoXLN+Oh7P+jumWO5/Pmu+g7wQYUkOgIMupE5ziCTXEZx+S
NMZdLnjsGRo2Tml/glSscPem51XmWDSDKg7bF52uu8CO0+GJq1kwFvIjwUMI
w7sJFi7yJIFXIOBLi8shF94bN0P51NwdV2KvRVOstDtwYhPeXOibst4hDS/0
nibnCDT234O0xmqFaTbDfL+LfCAchK6PijPlGI9Q4liCawrpyZ/KgVj/qW8k
n3RL/E/uTDSa6oqZN8raHH1riKCHvB0J6wZxFGNc+/pYchPhebPQc92zFme7
VTJ21Rk7ErMj/wf3B6KwVPik4+OEYsn4tonBVeNZD/eIsiSnuAvnSgKXUEaG
wOlftNw3TGFhAfeV/VoS8VDPEDdVDJD6p0x55Mys3NlrYMmYqNv+JwBlH5dl
E0xkIxFwa/qJaNnPaGvRCUrOXiW56LY7sHaGUfVLHMkvOTAd7dq9gnoN9Pbx
On+T+HXXapQK6tfsj96gQCVAstUifiLS6SrmIvKgdfPlu80JsIuZ8FS5pE3J
o5nCe+neZJy1gVD3ennPM+71o1RrmNYo7RFtr5NEHmjCBkX8xv07RHJ1PqyC
NG3eLgYSBNrU2U569WsMMVY+ermS8Fg75UmKl3fozwVWvvSyhf9uFS4K6Vhg
x0fz2G5zns0AyPFljIKB01oIEW+UF4m/Lj7710xBrVd0n9n17PPyPO4PgH+8
6SbvzOf/7KdxnwNL4rmTiWSzp9tjVG2NHNr5mxxLPTLAVvmzH87PyM7QyBPL
YnSFYfRguOAk9jvEhheNJePxDEfmoEiJk4GXIj3lZIlvjtrK0eN2bgvp9fe0
4qSL11TUU81c07goXuLzCKUXcuLPzJ5PmriBQQdPF8a0CJg0UMFu7h3mN10p
AIJ5l1j8q2m8Ve/CGN2nPLTnvzPDd84ijOWQGHicWzLKlRRSDG/rtb2WIen9
akZOULtSM0XWgDVQahHcHhhE2+XW0+B/BGp3Wjtq5iLqFmYVPD84iZIaoFhq
/omK4biH81BQ6q91cIytQmaRMJgfMi733OFY9MpLs9hubyC45q2lzAVTpCWr
B3gWFIt3xRr949S+jwPtMyjBRe7mFwyac1zeA5p+WKfG/wb2hRt4bk5f5loZ
Bdg+DpPJKuGshnAbyqH+yqBWFpEAx+SWCDl8j/jJ4U6/i32ktFPzGcOufWBN
/bsr1iGwktkTMWIBw+itxrM+JzHtWu5MtLaJs6KjOytSb6knCyDTzOvGKDtj
VAxLYDiM3y3tyDzatj+9DbZPIBzuiEH7bupp8IEhzmA5j2ZnkPaVPBkgTYCY
xLM5Wr2E5UbeX2vsYTb83Y5SkvSpxvLv/WMxbAnxUAFROoGoHF18Tag+8UsR
ZfaSVoMiv2Ge5JkTvND708I2dMo46pbQTCNJngz+vqrj9gXtMUwnb1qsvyL/
S29I2s4bERm/1FQX05k16WKwRXHIPxmshkoF6KakNg8Jfwaniw6TXgzNJUh+
GoA/zCunhdgoX6rh0aoJuhsxGazLEkGaS9PY5kTPqWMVCC9CCL25KIfFYmYg
RX0N+OlPC/AtMvgE4OnVPmS+zw/elFtTcWydDRkIA/yvbcK1DMnYn82YZ66d
GrW8GF5/QlhFTr2bSAQLY/Mjc8/xtRv3tExEyk4ecNZ2MsSzzvFTNJX0AenC
Nejc9aL+amnZxVHrM4jbZy2BaSua/moiTPBDoYx7EBr7oLcT3uMPtYn8T2tK
NZbX9X78nlDiIW8BHgjAayJSRW/2kEnuL2Y9sDz3TEWT0gC4Uxtw98OIek43
vUklv3FrkTFTbkG0QTqKi/eA4+GTwCUp4V/CevKiBGUShvwshP3M88Bfy0i6
OKblo5RMJCO4fq5t8UNrF7im2VmoG2P63z0kxp1cBbhDsu00aFfKlLbqn4D+
FCMQLy2UCb4BM68f7D4sJh8knAt+YV8j7AwOiizx/EWLJy3d4V9FMcBUtm2X
QCHjAkOi6K8/xRChm0Qs0uMXFLINMcCL8l8YzPQm6XnhrVreNA71dX5W6x49
sjxDZBAJIM3U8oIUhBDJm9FHdrnvTxxVkViPRads0tt8Cc9ltIZJ2rP7t3pp
Mmusvi4G3Z08yydeB+6tVqxWx688j7TIOh7EZcIY+1NA1cUjGSgSvXixT5ac
/sJrxCIPldOoaYC+mFPrqo050YmuUWV8DCGdEBchghAMnRjDaRZ9eDY+lnQe
wigkxKrwW6nFlWjVf/qtO5XFcMZSlN/T4Q4zExxbbjjZc1CrQle3prg83c0F
dnENAHN269gBtNDCW6sm7GGBdOoNJbGV0p5qSfoYqiIKeAwk7ZynUgRcgMIj
OcKAwknpXNCSu8kgqC23I18B6jB5HachGXwRthzctYo5w+ckZ25zezG0an1B
dPDjEgAQLbpWVPxqlFZBo00dt20rJ/nUkzqQt3qWxsX+Sx8ae26R6m6A6HMb
weiX2ieGxFPCBqScQ6ZtB5TWOW/Udo3OrYVuoTswnb5FNm7ntHhEBo7g5/pw
kwE57SiIvIVa5peIwZFD8yZPUD3KN8pNyunVE1uPD6J7gtN9n3bkd3hv5MqX
9ZSOJw4TbjU43swLPrwBfo7w43+eYryahp67u9G106Q5Kn1qKjJBYN9b8hiM
UEt4ViU8dyLsJ6dTJPkOh1ht/ddIfiPdczS/pdvN+RLbDCDVEEKe2uIgoPCG
MeMyjMh/2qMmPAceZeUmN03IH6wadP2tLqOpJ2/MVuhD+N3ZZO+Q0SwJTS3g
kyxg528XEC0J2Sj6bGBafB3Bb5tqDUBcAhT9bh8JSYWrHCDBGhzM2IWESdwK
QQ7vF1JRLR4Vs24i4Oy7ZZ8y0jino5SCxz5S2N5xo9ZJePCBDI9RY/SfvO9h
/R1yjnxaLdQ3nWh8MiuTOMuck51kUPhsXKFebWu+ksz++TAbbNHQXZ1K5uBR
3QIjRBKYdYhte8Oc9aZQU4ZSChCkyplW7PBoQjN9luVt+QDyPa+AS4asFvPw
PSbnPwAz7pzVU1TUAQu3zDvFnASfkaFlwVBEXfWxF4b9NG4BmLuzdejKgbT+
6RSn67obien29Jik+RcZ8pm5ypd0UKzlhxyrJHwh/n6lJNhai2yQ3W+/SXR4
PmOazumt792mfAXX9KwpmlNDQB5z0Z2hc+esdiQsW8039dPhcA+u8LG4ypDS
B1vGIrbbUZNobIceMol0rn+Ss/xu+ojtVAbm1vlPTnJ4z0+V+ttU04PirT1U
RThq7paN1TWBpDoUiTqLIB3ByWhcwzytUCWTS8BsLa/69rHKfi3hEbPj8ega
XIIi3KlEb4h2EOwR2/HDkkyvBWHoD77kh6alKjm8Cwl50prLIGwOv4Zd1UOG
0WLlOV2zGub6dP6LWX8la1kSAvZo8BvoY8dWl78ga0rLtD8OkZUckK6SpYRt
P3Sr8PaZhwCE1Ajc5eCRjRFI7jvWU/MqyHHUOmEHdKUvcPneP7f5Q2Y/6OkO
ZmqiwJ5Vs8Lobq1f/JzBTh0ePYceF/rGXRDfpmF8LjDQki8fEHEVrpU8ObYM
d9EFRUkVFLSHBYumY3wUbvTjbIWqh12MGmEe3YaiHfXam5J+BhoYnztAwoDq
MAofc6N2i4oInVxVIdRPWp0Lai8iNl/aVeU8AmyED62HLs6xIXGbMDYXJZv7
A4QVVqQ7jLXfz8kcc83ui5MariWJykmoKGlyMGSkT8dtjc/8EV6tW2u+bjJ6
CkUM/EVtQBJL7ODMXJSBp40Jbe1ZcAXYQpcHrEG/Xt13IEdcWnW7TVGBD6gp
Ekb/IlaRD9823r1iFy6inUaZdAf4jwwXlpJAkfHsUVCMHfMWkhlCsQhtjgdI
b7y0WnN5ZfkCu+fTM5pkCzkQ6mcX3ZSvqZ/5KuBs8elZ+ZJ5Z9ykCFNow3s9
6G7px2ob8RtxjpEHWaXp/LveFZswBSiwSVIMIl17qb2NniR2AWdyX+M0Lmnm
gRpUNmyduh/QgcxYRgz7hIpsAmqDsqBWjbW5nMH1n7FPxtY3WNfWyngrhNuu
gFzReyrfIYckid8EzyqHb9AJjlk89tSxu2nj0z2jPBGoKdciNfFVOQTKA8/Y
en/9b7mGG0XOtgDO7XmvsFHtCkMHmocwd7ykVNqrN22f/m9wT5PQmLbrx+Zg
C44WRQKwuqKVT1Btyn1QniJyf2ztI3Ct92EjAoTY55KXYyWW9EI3UbgCaENb
ehtjvdNZ9SZXrQGvbOFbVAovSXsUFYnZe8Wn+kDDFhReBJ9ZVb+akTWGBW0O
J6Li4TwjT1TWf1dC8KvYoY/9bspLX7lzGhUIc6TEXXZCkY5rS8Cgc9mh8IyZ
quDBc3ttmwLv0rFvSAXco8o9c6dihmNovkHk7fcvD7QWJtPEDu3gIeHoMT72
45UQ/mH+TTJk340TfXeGi8teIUxwIwGFbLGPYxVN5gOiaYSvEaW8uiZ9fond
W9DN05VAr0vLsCPSuyksw8LnDJkWauNqCUnd8xN9btoAZT19iZyeuYmMVgp1
AGC/HG1PGEsJXUM9a06X2ZyvY5ybxfM80FCEODkwTZ20VRPoKzLP/r7GVhlZ
eiAJm5rdXiX5ipSgKD+sG4T5fQXYHzX1hEmFekF9ha1E68K2MrehkgfODu5U
rQg2PV5dl1gLh18uZOFHbLVTPNuGuuOtpfQ+Q3AX+hgaBii9c0fhMDC2+Peb
zYP+W8I7AOHKqrIKVFhpyO8n39wO1+vTiH7jtkpAl8angwAED6/4ISX5g6+V
gssPHKtd9xntBK9dqL5kUxws7jChDRNl0wjRKIXn1Upr5FVW3rkc+RZWMxzC
zxrUWLpwFlWizRUh3K8+RdBIacuTEi81SWCJ6882iI0JgM6utZs/5eANQH2d
hq8ZziuvUWFty2X7QnWxyfaZfV4lwr/GB+OfvPS7KTwq22degXXlnnljszUG
qwVuctw2HOIeeC8g4vU5x7srtCspve94cXn2t6t1IOD3KDxq+Ul8Ux4Q3PlY
Hy75oLCTDXaN71lattIqBEfpr8u3yk4zvCCqDzpPq8ICeBxemphGDT/JLKN1
VnfR+oOe7slOAOAe6kC7XIEq1ZzDAwUm+ap3zRTSPVsFa6HQl2sVaSctknf+
/yKBo5r3II4J4r3CAQg+JYYWIIqoEB/RK33a1QQ3hnjgYeq6JtkM5TH6E1tj
UwHgvU180TobagSI/jNdEVKLUHEVbW0EVZDVutBJ25Hs78KYbHhLwfqGNMyn
LvpBhVJ9F5TVDv7B4iBX+Mvpvfo7CJ7fdQdBtvVht2tS7JcrZSsCHHv4F/Pr
aN7o1VsRQNNDKLJHb3E8FaSWs7XiYVHsf8qISw7cGKv8Mn8jEye44nbdd2YT
sG9krb7O/ee6C9ikQExebhg4WzH0QCJEQt32zLT6r4Jv+eRHs+rPyX3ILZd8
CgQjw2OQl8ZUoHaXZdHscPnqLfSlqe9vIObkB45M7N0bh1a0bcSqQ+FA/L5s
m+Rczd9Z1dfbDX0eQ/5Am7VxhPqzckHVSwhHJxjASei6/PAhWevsz+wSSwO1
gabe9Ydknl1LuxPi22tyuCgBcRjJQQ+7yUnttHfBPXspHJ33HVc3+07/LgtU
wnc7P7pLfvTc6KQ/fRh0AfMiPz0/Dih8hOjHE6PE2NVglV7/RXsPeOtEDhmd
xZjjXvzhFqKG/A0Oc/XBKllA1J545pVq9GTeHwT42kmLAUPZcJnfBuqVk85Q
i/bfoDaqfrTokUlZTgyM2uzF/sVOrtCHzpE44TlWiAVPg0RYnJd2xnlCdBDA
qKj3KHld5ZQBsQGpygiY4Rcv41762bXIbXbCJmIkG68Lj862l6jA2dV1KddO
esSjnglhg7xGK+ErmlbMtGz8MPGZgYxuEze6SgZN3z0TqAvLcElyucGEMT8l
6P0C9E2wwrAbGF8E+Khd4wT7aHt6P/73t91Ct53kg7wd+Ui5FtumsHF0m6R2
nEqe/KnSdqxBWqfAZ10mtpvvMBtsAr7hq//cQGsfJm1Ac+txKoyV0BDP90Te
Uew6Kn/JPexmGuQFhRYl6UicSS2+xEbJC2n8q6U9kOoZ9VERHeRCO/rCKixS
d1N70QLc/eCzqOtj9JgAepdmTBVenW1eAT7SI2SOXkjelfdGMclxkg+mD5F3
FKex35CUMx/EPB9bjX++r7CwJD6ERIVsd31U7pUtfsBr97OyLBi3za3wSsFX
tdx7c/zWEkHmNuKYQJOdNG5/ddwfdA/d8OJRJPwnQ7rqO57diajbSoMS/dCb
YKUpS2EUfpjDx3rcsFV5pxhrZ7ZapjhHv0hLGceKHYIk/dMgc7ASAFpBbUuj
9FAqAtaCr2AZ1fIL6kRhZm4GwHlDJzEv1A+KIx/mDvLVzgdCk3sji8UXuyDt
IDsijlXrrXGY2UPULyYbMivSEPJoDhSxQ54hotGzf8NgiGDUuOW4Ec44K40K
0tltGeA2pl2fJ2Aay3RietsoUqJuso/mFnUJTt9C6d1gOPyRrEomxpJX8oJE
2OxejBdtvpFpYJY3Kysty+kI67b9xhpFSfM1iAA/99oy7qVKLd8HKGSRLmCb
Le1bY4eoziHKV3a6fuXrY2bf1Qk2b9OIsfM0mhDqkaA9B/4aszeFToiuXggb
u9TTsQYqoDv6b+GCf+e+mECORgEULZaDF18b1cSeM4yr8UQzolScHXvefmsY
t+jAdXZFXqrNVH04UxiK5/u+BI23FiZn4AOJPWJacyfboGSah3SORXZniwj1
1saxLwhDQJd2jgeDjKM3msWSuLsYJ1bSXKNi6ZcLg8lzurB/oZgXtRa7IMLU
1qdqBxlHsFmfuRq7/dG1X1c22xIqIn57aCW10l1hoWSjOCXOY2z54tvKQmZg
6YyyYXGsfS7BF+FxdDAd3FmPu+M16H/2jh/6PYZskMqpPIaTzXlYbySbYkEq
tqZBTUheCpuI2e4NWdzRTfDjNejBHjI+IyErVAJp8+sMoQpI/b6PKG8397P+
o7wE1vZMz/2dbcbCAnF8wVNdCKgUDf3R3lLKLiaPuMd/KKP0s7UIStTutuNz
0OkxzCNVnd5I70TUMe/25RQDAsyd7PV/GuDY0p39OovrMescCDxYmtDHstoL
wkjmvuKkNKk3yO9YFCr1fp0GOX+Eu87HTfAJ/4TqeDaqx4TNIpa9olC/LBA+
O9ItcBxLUJYVUtx6KFZkksOKzwFlH16NXFKyZ3k6jl9nmBtYzLg6QylXH5gU
p1DKwr8fAp6+x4XyOhsS6iDbrjTgPnGWU5QyXE14wn/zzB8/zG513IMNqRbw
l6NBlfXqiNtbJxGMl3zINeruY90p+ibW2iaVk+3JBBzZ9DUr9XP3WB+zvDaZ
u+8nN1EL9EQq+PLwun1BOVZiN1MYKYgbDtQTS/9/GLY2J75hSuDju+DDEOUW
9UUQsNCv0lax9fj7LsKicMTCLUCXhIsAqu+48+rz9+pRkWESBYXlcdioQPq4
N8GZusfDonfokzIRcwxC7/6IhPP68wKXJeFAbDJ3iYQ0NgJEVDmF2nA8CZ1N
Guiblgke+BWAmgfN7CidzR8GpLKgemAgdXP62nVZo7LIvPLK9gXm3jKSQYGE
fP2brf9FCMp5c7Ur05pEDlASKHLjbQMfcvFFLxIxnrsoYf7GemHiMWofBZEw
mhU2ZUSMUhiDVKYy6sbValHZiqhqsvngG9cRV+SRhJMD9BT88/UgdOpLxXhf
JhGgYSjD6JGBKjMbGhmtgEnTvBSGeaInRpO8+H/62WEBmAdCi5DfA0CtVYcn
orpZBHplEbxPdTXfXH705XABf2n9UPrl/NhqOZ0MbsKSSfmmXWfvd4BamEXe
HS41NfLnhIPMXcJDTGVVUxW4Z6rIVd1WQzV7NpjxY+rSQ/FlKu1e5IP3+EPM
0ENLjA5irXOZdV4Dr3wi+F5aaZKHgfNLqPEuocMgHG/n9gc+MzAyV63rrK22
1LIw2SeBu/ZaaX4AeT+K7eVykweCn0o9TgMcxiytHhcDl0jWgveIl5N7dTnT
vvL75PwSDfzeIa7Qa+DdlKkMxawcQwcgPzdw7AUHSMMdUhxKygPygmzEURZV
ozEaphyEod3pLpfYB7xHXkAP6GX5kPkl5u24cB9WpPBTRKM0UrMIeyh1zPi0
RGppjfqHoYqwtLLXGTsU8EjgPWCBCSg4Jym+oHtedn7EFPR9YXi+Qhg2cawD
I9GBekxkbPWyGbt+ivpxkYBLdQ2hGAkljcx+H964lsyhQAPGYceUn+6eDiFy
3dJfcDZAM0Z+qUQCbZ4csAxKPn9y+BYwZ8r2Ko9G3Gg+zHKCia0iSifdBQVS
Ma7UljyAVPU8sxLXv9iaeZwgXv4EGHFzlMgPJt9m9ZN2Ml6bdcdbKJwWV2BY
iepLvcpIq8VQ7RWyqXe7ilJaQQfcD+2mDHSGRHMchRITs3lLR2aqFwrgrYPW
6o3byvQpsK+C6vqWTQuSZG7KFhmBJ255f0FgOAZywAj/agaxrDr34xMawMmf
BxUUgzQD1oYV9oLBaTmRV91uk/DGivGYzeI8o6rOuZ5WW0NnlUmKQ2NYIN46
1wgw+6KZl1Y+EK+laS4lTtTOUW1C2Syqc4mKQWBNTslE7zrBF7LCC3HO1UgS
OlCfiKDWSgJUuvOD3UmDIQanU12vDeL8+P2IxZgvFp4dYAer/Nw+1uCu9Y3x
MQ8OnVcVGI01Dv+ym3Nu//CmD7fCt3LA2qfD6enIAfB9FUhjm1qaKr4ucSsj
gSPmgSR0BO4slSUGNOciVMZ3KTZRd6o95uU82jwm3dhJZpfcp6Ku+OrhJtq4
dgZoj91BqGGa0IvdtQ8/MItZjWTj99qqRkezB8Ed6iJGDOLlAzLe9f+eGjOA
tUm1BZcUxlpd9Fo2qa9n5itKtEIE6D6Uoh1luZ9Fdx+5Xd/r5A07/05Pa0o1
EknmCBlpUgJ3gyWI4qAoGmquI8CbtYmFy/mC9DKluAr8sKIm4NhTVwPeRCDW
LdHbhE6vyVe2LxIa/ddexo/OUxmzaMPEzVO9EAlFWmxbPmsC8YZLZh2Wbyt2
vPsV3U8FD6tYMu+WLH2JLsXDV7JVzNlOqAmORi9p1rR/TYDQ4DTy33RuwzuF
MbZbfw5kwaG/haroa5zGq1DLqRcohnNVwEUba/+XMRHnQgAmxmOGjU0+wgQC
BLpFGSIe1y7X1ZX0aqAt7AeFxVEZwjaQIO8oNutv7G/R6oPaPbS72sgyhp/J
Cx0EUI+Nhb3HrqUkVyR/uBXOutoVMs1eqUoa5fJTej3KQAxsTAJ+IDuPepLh
HX80xYwas1+Z6VozuAbqdIAolcdfk/RffWfB/U58ohPyZPTnJ0prppXzaAta
GDZUhIQ6kzVbQbeWqezqvJNwaxjQaKia2StH9CRLl1I5TEugS2aFKDgjDcrR
9nyoiCtLH17fXajOWClHX+sjWziN1aCQocv6SDupgTh9Uc944vLJuadNUfbQ
Fvh38bnM3Uy25tvkI5k7LZCA0ToThrjq2PCZ43s0MQGUxRTXMMRtzzhhFUJ0
7vNM5a31/guW61h0KDMLiLOJ9qNmB7bxNCznP5/BEzlSqjELC6xniMsJik1W
TEDr2mS1L45ib+QdgvmZMrrvscikeysTP9uPFACStOaDkw9zQsg0adSs+di6
COxibbpd0XQvCvOL9vd2RZr+2WeEgSHXofIFKvlcDAo4ilH4GtXSWVnP58rX
hHR5MQ4kNBj3IgFxMkn55y+U8UdbAXq7QYPOe9wiTGky0Yh84kPpjjbQZA86
0ZfhXn+nISNG1DZpMe9GuvxQuwzPeQNOUcEVaPM6wLp7LzTGUNpqPqKxb5dp
T0hGEw2Cv6C9G6mxVDCJvJBKgVEGrrbwbrPlEk9X8uXUNZjMbxHmvBsNJIN8
70mhzSl6q0AIftGwXIrUFr9JKlnecapiEYaSa3DGF8P6MMs4xLy3+fJa1pjw
cobzfSY74orSb82bx+IbPSCkoQZYJza3vFxBC4We9auzbvGl3QAt1HFg5zs1
Gmq7bES0BVAhq4r1u3HZUkh2wAXLkWs8RFvGcNiOeoWmWw7IvG3sic5eWxIi
hItvmLKKG4fBLym6gwPPIuUESs/nIlBnXcHF37HQv0KRcgJVDWvujzz7OUxV
MS34KygiAZOHSPCwTTxtc10gy2nPv27sed7fAuX0ZJJXwMxJLZ6LZ3/Avtpu
LxwGu+p/RNlHnD54QcZKMJx/YoeBQ28DtRhnkxXn9hgBbO+k7k1np+mHoxLl
ao05A9NhScgsf+MGR04ZFq1ImYCfhidYhODrZI4hRxgi6h9xEUTpyTtNtgUb
8O5VJJ08xi4wNZC5ohUV7d0PdiuVwg5NCuaav3ASEfq/VffZD1GJg8sFeMnY
YebgCmMGKu4tnh/+ouAVpIfPLKkAofHm2/splAkNxdTW6D9cme7Dxbq/7aRO
WIny/YIv+mbz8A0Z+DxLwWFvZvtTKX65jH1VcpUdCWfE18o7TEYE9QLDMc4P
mKN2DQIhfqUYSZbgxhQoh6iD8HE9oMfnwLXjE5ZuVkZAVsdB9hvIuM/q/PpB
IG3E4GFIhhzJ9AezfYGz9bgTVFTzTUacY2UugetxnwB7ZjkBVtAMbpCTlwBc
geNZ3XPUVD4udgCxvv3nYR+aqLq+5ceQG6VCgNDZH8oeiQHYw4Gd2e6wOGZR
0HjxmxQ4LJnrTN/nXyEjQSgsoAjHMRoXLXyeE4yXRAzIDHY3/N39Km2fUgdO
DeDSKF3BzqiZ0SjTM9P5Y3YVHEpB8Imf+GPd5ywPYLB2R5Ndf4mOeoTe1p/T
blGCQHCI2sUJ1/giaMXHYnIjA54iSLGNnBA4PNc88iukfzZB3xfI0FC2lyGT
5ayc0OjDJEnMVxhc8QTMJVrz9yoq3/Xpl0SxJeF7CuCSciWs9Rw9DSkYMRwX
it6+eqgKYRSzTYSoQKczaGY6f4UoLsSYJ3SaDAzJEqyGqEqb7HE8fK1QoSCj
q7vV6fCvd8go2wChL4fZ1aFIV4w1PKk5zm8iRYn7cTz73OSbOboEpOYcyJT5
sXUdEjg+qA2Bup57deIsJSRDEhVA7eNraMNq8KkFq+HtQKH0c0YOT9W/vHxV
tC6uhI3Mr7BtPQatRMhVjM8yMMdsJFFgA9yvZ85sWq4O63OxRHv8pbSWlLUB
bXf0BXe03cs0pk3l7KZIjE+oGM2U4bxWsDPAaIOp2zRnH5QHBX/tTAXr7LzU
YsM5I4TjYzOuVuckude1tH2Tg+yTbDXTo177MXmotlLYD0PWsEUIHiIvlv8B
XwJ2O1Tr3cn/xsL1jKPzb1JcyPoIZsVrJD7iUp5V70/9Pf868liezLSa363T
kNChUoKIc2pyrCnZ1wM9Oa7YC0JIjODN1Jt4M0RM484SROpbqODfHkmH45dF
iqMKueKhRZcjdNy634swf0DE5zT8ImjnDgWjlkJMrcFL6P8vzDr8/cmHPZO4
FmceMIp2n4KjMxaNyJMgwNxp8stmLk4X44wxzeQHplGkMET9bf6Ig5IhjQoi
qw9opTZhpdlzdDMcnjKBSbXCX3Y0oofxnB7ByPyvyxlbwtzmILCj1gf0ihNb
E5ZFr7M4YPb3GlGKfWnJemHCuWuie9Vh8oaL2nN3R6IMvqNjkdM5EfxsLZR7
wZqZmGABySC+eHCgZqjY77/5wL06bwzRgH04x/o348a9EJNE4QP08DNsPiGi
dcSmkQ5+2ryet4JYspj8QTeCrlWh+T10sVlNyr7zLd4Cvfv2V9wVvDBSplLn
99Th1iaAYgrTlRI1VGoNeFdYhxebRX3zZzlkqzFjUaBJETW+jGqxtWhnmVKN
x8BZ90HKoRojvXcwdMHwwSJx8dCT/RoAiH79qLdrejI/Gkg3nr/3xfDW9APv
mT+jS/lGW6EwdfsT00vWdpa54aAwZj+dmHwdX/MyHbMebMvZGoDw5S8SRMBb
YoMxi+R3CmGE7O2TDa0Nh5kwBYiuHB5fhlKE1Ka45mrgHrRkCcL62kss2QOx
Hftl9OCNb00d4w72XMV5EBmAI4PaQgoAKDjp3DU8Lmk7IiR9mGpzqmOXQ1Im
F1t1+ZRQxGkGfZuD9qWjf99GJWn0JufJ+454oiBFwIhSHVOGoyqQTslIKBZ4
KsI+6OBYnhBRK2A/UtUTNPwzdQluH7AEBbXj7GMBfoPynFj5ZJ3h0WbuGBLl
w1Pec5FjKa/uDQmlBfHehTTREYJyWGYViWayQp5dpcIMzpARLSwqjM3VFbiQ
6vawLESvR5MJ+3UdIKPGZLp4Xq+KcYF08fyeLTGOKjiGvrsnk4dFZd3bRzX5
54LH+6V+1JpGv7nF2v2C/Ovix4h0cMJOWN5TUfMqf8wz+TRTXNX5HlPZENdm
qODTIqU56MBZHAS1vitblddKwXhsih450yaqCP+TWYRIh4f6zgkLb/D11/ap
XYkrG7pnNN2P6uohfkcSNE6MKOmnlNr9dgZBeFJhf3LtAkf2EJ7QdV4vpv+R
QzxxxcwOT7543jyebuau+YcnZnZJKodFzYOtPIdvbXMyP6tg7Xvdp2H1vyKs
UsiMP83mRGqC7uPieoiiOjL6uLtYWeHFqkeCQ+E2DpIz7Rxyrf2mlOfiqUeg
oBHdOPfQWfKkdLswC8AQyR+2ivfqQ42v+qd8drCSh9bpjgLUbDklVymtLi9M
EOXDZN/zJZ6oncrBVBXwWxxEI6ovvvtw4aidRLRZFFlK+j0pQfCbw7E72QM/
Vwy60R4P9QFrB0aMjjmoWiCM1DIPkkDB9ALz0Ic9gzlGksLPox8+rXmpLDVP
WBXawuZzee/Gz9s24/KkV0fE8XAI+qe4q1v0wTr6eSDZ3F9SPnrMdC099vQt
ZoayyKpTRdaibGSJ5AcCjOMPFhce5LzWXS6dWvNB7hQpNqoNHiJUpr/6WVii
UsIQsogV6oKvdBuRpvAm0rnYlhuoiVnUMGxOxfS5K4C7I1E3ldsYbJckWt5/
x35YBIDfd27xXHHwX4ZqK2fnQ5TufyXMs6D585mWsZhwbgFSAyl5dyavYo9J
X8smMApthEx2YxndqZSAqaHPZCLPkZ3rIWIdsOfzEPKC/0iy6CtlAByu6XvF
1k3vs7l6r7yWCVxviMmQDi86PX2oNaZNudoK0nzoKSVPtsgQ5GoYna/PyPvx
YkVqmlxxz/UF1cxyAsNM3msClwCoyIILhB3MsG7IfA/+hSFyt7G8MlcQhs0N
NrZPrstOPA3BwsKz0upNzyOQmEdkwsI4izb5Wtl4hWbbj5MDosbl/meB7oyF
Juwmyss0XECN6VAnh7SK1vwmQ0VmLHZjWYgDlYW158HwXr/bf6MKiM/+Heaq
mUckaVBp00x5HeB7gYq69Sq7BlQ7HVPcHlcHER0vkm1ipT9H5NmzdZKsRwOK
eowwQnCsJel0M6sAYFrz4w0ZifwVQwYSkvgStL+wYBhMCz/sEax1iA9HpIxg
ShBuIVbiRVIJGDr8HwebdCOWeOiauXHvMQnfDJET9Yq8OhIknDIx/YBPI106
BzhkDUmKrLjrWiOgdzQJOXeAsBmL0AMe8mCG3r/8irO3re1AlLBuOdLZ+oIt
fOOcu7A4+xO8yUiJQYWUCyA8ucVDengucgs/rOEDZVhJr/0OpVuzvJjqx3tt
EwmPUtwi6xasLLnjg9BkqIVbquA5eVY7qbWqaQ5sll0cOQIn/cYjN23GWdAV
4zEexWH873KctEF/tWQtNPeJevWjo/qM/RRfD7qKaz2jZo/p6Mq/fEz1WZwz
925PQErh+Ldw/4Ojt8eX7K+Q1R4x4tTUQbAf5sZxMGQW4ZdLnoHX8gfB038g
6UWeZ9iSoJ6W5SuFz7DtFARL9j5v2aSNqPWbyCTXYvlU2JgCqFP1pj5CWM0m
Hfg2ip/jqWgEwIBHG9ejLALjejjMpArbGx7VssETdtOuNKw5tgl4mzNCUc6q
51BIBvUVqCnlTcJFDpzpDHZO0hFNbjYCyOmzYfDWMPs2KHquz54FDZDG+j/9
FdWlTA9G/C1x8Uz+pFX+dCyBh3AmRaYVNOjhBKYDvh0QAqW40esn6MvpA6od
gpF+3D9Mg8+xsHvoe6DMrFCZCSdY4mow+E3zK8GbJeclBYgD0SDc2OYaofkT
0DWjvpvo4xY6RffN8oNOD10Ixjit2qWoxBTkLnkIosjmU81MSsZeNY0aLCPz
rrsJz9wODKc7Cs3ddG4SuzDl9/Y5LD0mNK9qxzUDv/eTj4iqI0Gudh/UOERr
LrM+nbC3BOwNyENMjhBfnb1IBW4gqHTD7KtUDVE7ZJpYO+WJfnw0zQXOZ41R
kFYazeKZV6oUD+yYGjrYg6ZQ9n8nIfjFZe7EKRCiRIuzXsgKkS9ChYOjOvze
qp1zz9B4+giabWbqjAE3m+amllg7sc6Zaps5QjB8Musza8oNb7uYc8Mkg3zk
ZSnwEQlov0N9ku11J4qbsWBzuDYj9j3XjOmf+KqseLnpR4Rf+Wq5mu5bqwZQ
bZSY7+n2muT1zYRl7UHmJepfIAAe49qrqUs0ohdFuRwJPajc+i0WKcxW0d17
Xdy3V/POY9TzLTAGB2DIvxeeSwEjCRVjgz02ntWaHx6GpG0pj76fKFusb9oT
iRHBknWg6Hh8cUN8AYPFfmN3KdwDqo1yaTpBJnJnsaK9pdtwHa4kNLhqCYE+
d8Q1CaqbsSfnrvJ8etNGgz4xMlcKxNNXBRhR2wCs1+ukfuHacCglFXfahV/Y
tbB3LwCSIZ1EqvdPDeQzDQNTw9vPH8BDl1PyscTFJ7ARpDlJxuROGMBTwGCu
eZKAYKTOSiBu2WbPsAtUmSF3Yjiv5xneJtQUlMaM5cR9A1oEuDGcuW07TGX+
Io0NEpLaTTfikZqGJHsq0TKKR2ZbEQ8mbP/jnpRtSOvO8OMioPrzoREZ14nY
W86IayeH5RYO9/x2c+zQgurJyfsI1qVmBvsYjyhthkrOHrKEUoNvSoaoKHAI
mva4nVrttqhfBVNkgqkUjynUEUR8kQnZfsbKIM/+K+R6j/J+FEt7gR3hL/V1
fc4HCKe/VhAEVX5JulGYjF1zQvmyi0kjpChMcWCnju4ntTHLZmzGoiuvPXj5
TivERTsn6FVgmEdxpdsV7mV+bezcX/vWhicv8RcDg0gbh8DrZFuI2s9arDxw
fnZCoYM7JEu0bYZRnGRusJk0KeYuGMg6DnbdOZruD9Vr7tjzLwhbVYREG9Jn
nhoX+gTfRiqKPVl8FX1n3g5mdjAQF1EjQTpsUy+L4FqOxpPOLYlkro5wMYhk
85X9SfamMZm+yez3Y2m+sCFUSuEqQ6ZyxftSzUx5PKjG5cmHSajvBSWoifER
CrErMCRhwRK44QAOxQqeelbnyREeGgszlULq+Krmwwm1ncmsGpwNcnCDZeaF
9bZt8VaifrsRdpSFsN4QOu4/JSpxEqDnOZZSXxdHyaJpmx6hy9uJR3qWjE4H
wWDN7Q8WVBn6Z0oUK+DpL2svlGbiF7sS38hkZX7/x2mYIcwGBybwobNWEyr6
nAR863NgIicLpUpqB36JZy8iiwnvI5gOASCbjDecqg8bAa1FZXfhAgh2bTbc
vNrCU+D+7l7dU2atIDJuS/+OefDa05k3d7FcsvhIxkwClcGtcxUZDQ2mJMBq
aMtTrU1dSOOJ6gJUmPi9PgHKyUm3VChnFo79WR46IqH+tJSukMcM2G4K6eHD
0shJdMc3JIoRL9hGbtu9ooBr19i5Hd+UjJ4dQKwCvJk5bpXlxDHb62b10yxy
ZhYNDm/Kt9EYXuIE370f2MnNKotuJwdiaYIqEfyLVxstEGleEaIXVW25B7bc
7yZkoK8MAmpVfIpfiDH5mCCwZ4X1LGbAZYHZEHEXCGYZtXul/G07UzF0rT2u
o1Z/sY9z5jW0f5+Aua1E8WRvITShIyVnLt1Y6ytiVHjyn14jr4u0ovuze1jt
vUCzSEMfCcJYudnPZoPKu/nM+04C3YlcXMR5TXWLZ/VpKK0P26RCeaaAQTXu
YyP0agbwxn7INQaAoC71Y+itpAZvrxODnCIH2LYrbId6yoCZsd9qAg0I+sHJ
7RWKAZMJ8VphWO/bbYZXrdkuHYMeHDt3hIEoFxh+9RB/C53jO5GdLcRiKvJS
yQAoAdecGBjYcbP8uWoxKftXvtxrA7aldc6rC8juJE5bn+FejOtlFSwj6fcQ
Nk38GjODq3GW0QeAFZPdyiYuFJfC1V1SWfeonUs7Y86DWrA/vQv0dC3LUB2a
HR8krEeQXYYB0ZUBOqSLMaXhCjitfTirWu1hjpXDQ0Lk1ndgh12S/ZGL20QZ
QSFAhWKssogJqPo+IofPqnIV1GJHKoCXiQ8KyOT3EF1FJNkrCFvpKCcawY2I
aK8Ey33CCAT/9cOxD7DLvWsoJ1D4QDWioBKv3u2+aU/WwCplNXbG+vBd/Dac
WtUSxKVJJu27yIWWlqkr0GOPGieKC9qOqfpYaAb4T0y8RnZ7TVfOW+/DY7/6
oD+OCPxntywwIMehwk/WmwngybdkWz6hxgWCozY6YS00StDly7bKIODT7SbI
jMFGT1lDZfXtf02QO5afijvn8Kb1ud5F0GE2CP/M1+PhzcIOC6S8ghOp/6fY
dUiLEWEgpUn8QsVIfXlTjurgq8WrXDv+dYNw5xKGxMV8MKEFx9sOkoHbzcMr
1Xi1EKxWkKPXbiea7a4fmqRxdSR3Mv6x4+Em8+p95S8emuHdGnJ/AKPKe4AM
SwHVtBIYWLvCAwlj3gaecDWVwUG9gl+4AbogY/9axrHqYLwvosi4IwBo9zsz
gauQ9lLk1PDfsRltKScfkJaKdqdlHvFwuPsKq2WiHSdSIQP356hekFDfNakY
MmhbbfPuqZjsJE2eTW5RUg2eD3AY0j/3i1FiJFbUrszLn5LCjTCg0pHqjipo
mPD7HovyeJpOiUwghk+AulR/unsAeZtUBEJLRXD3s63/0p5gJhNL5YIWYCLT
qU7HGLLJ/mjRXq2gQ4ciwtLh3qq6ApfMVFy5Qhh8rlywvn3kPEwrtDb9DOKP
otoRYUy7AUogCFYW1drpkAWsp6vjhnimL6JK3G/SRh2CGurFe8UuEAwqvVAO
ERlO07lFqIz1eVZ3+UwWQam9Fz+EDC0vYUT8Eb9y0+JrHazite1Lf/Q5sqVZ
1GU1G0SH2aWSSk/yhEnJgMVePOR7qpvLduXCTxSXy7ZJlQzQbBvSAho7FKmL
UpeAELy1IAeqG7E7YcQwJyGnkGDQtkoTskH7dm4J2Gwbw2Fcth3VIu/bqG2R
4+gSGrjt1LveX5PmHo3/FDISDxwLnvwSSDMGlyLHlUA3UHBZNaOBbiisHobE
wjmPiATW60d69FbO446pkZFCgTfN0f7FFHnbmaAiC2RKooGsGjts1GiKPvQp
OA3G69cWNxM7d3Y0Q6GfzmKCjsifbJvlyuVqVMCjiYLNtt1VYHMS/CKYLm2n
zsnAj9b8PpNJ8vnIRCMbb5bPyqTLXt69cs8pw/kvKDkrbUYhany//3j3O81a
Zw5wZTdqkmNaouKfam+eWD0Q/fXfP66xPZXpUMKr69BRLFQRz0V/ZRO6y8n2
gMWvlobqAyZuBh5OyEwLCjhfGGxf9pHAzkYiYHKoFm+7qM/8V4F9ZvjYWklc
LPH7FYgg+AHeOdmwVYKWyZpg3rU3k9TWnboGtchfnmhS9k563wkuFIvyAKAT
1lXlsRdBu+k6V7iw0hCY+JeTfRDJZciMDoEanE01rw+J22/lSWuRPTsfjBh7
nSfYlR3Y+cQgC1gK4GhHfeCAO/v02pOjPBdDZpMVuxGxoL8u4XrT7m7xSsg/
Vr453uceOObJzBE/9XwhMCVua6CxIZsZcdDyMDsFwVEBGUCk/GIMJpCsYHJg
/dv8Ol1k0+gbnnCUx5qXaoJ0mUCSwASV7Ex52+oRGKRqQXp8d7GdrJqboD7M
RCI/bfN8ZBYxMqFV0r7DMeMEDnigvCkyVZ+HmGf5WIXSUjdP+yVKSmKaNoes
8v8ziRbtJHsYucssrwmFeBwNrMsjKJ5zrzFHhSMiOgVwZN7tKUdXVF45BTXQ
wY4CEDKmONPk5Wip9+3k+dI1YCcs5C1vikGcR7FwOyHHk6YdtIwtcTKaEuKf
KI3T9xB5e1IKNI1CH+HyjWAvpYPPyejp5EY7KqMS8PqWOLCFKKrkDKSbF1yB
u/tKKP+r51U0jinT/RdsjmjhtdfvLDvVnHqx8S+dtNY4o5OJL2xqHhhAiSyG
K2h+GW04CMoheWhIOpfYsUWLE6ibMZpNAHDW2T1EwmxvQWimyN3D64MaGBu2
pG+XZr0G2r1RkRO6+7aHz1cWqIuhvCiER2L7ETlJhbjV0gotZnKnord1y3uU
24jf1TYJvH8qxgO1+0fImKa/dxE/0d0p3rGtKC6Z4ph9NaEZQyP3jKfzVnXi
7oSr0p0YUX+enth449VWP06a0v8N70mjcUqaxS/IjcCRrSCZZ+RThZUpMnfc
EIFr8CFTklKiEPyTbggwadI+cRDtO9f0exvAah8zDfbHc5QVI2bAMZHFL1wB
1S1jMJU79EcChgNdoPIv+AgfEFy02g341uPreQnYm/mRXRJiow1d9+B+WWiu
XccdWpHWU8iLIIARIaKEJq6OZeNFKbLWGFbwxG2mi4HpAGVcQQm3KEBmOhi3
jBvj6AcyEefjdPCq+QS7JSDeLwCUqmIDxTLqdzi74PUK9wNUJon2w4Z5ACil
Z7EOOE6SRSp6+KP0g+EVA0tmEVya1KCPr02bfmGULVfUQmm1yc2mhbkYrWe/
OmS30vIkXCo5nbfrWQZiyOYhPhOLe2pYQhv+tqKyEWtPvU7mXH+TilBnTUhf
ulh0tAOOsYJG5Y9prtHN4B3C3l3VZ3gffomu4Q65t0O7OYv3fdro4icNrtuq
BcycqJFIPg3H/JKXE+acQV4E9MMSQCgiGhnvvEZEdBZM8POxWkPe+/g6pL68
UgMRvpuI6VHo1Rom5HhQ1G6ivRTOs/JQBjhI60WpygvoKzkDjXGMGjJF1slT
iY6exNetKEpSmtRv1VPavngt+1MAap/OMyyPwUJl5JxgykFU6OVSFKqL3E61
pWHEe+vMEOo8F3Cq206+CYOfQCguoue8D7eVXq0uZhsnYdjjwEmS3ffMF7TU
Rya3/uMlUhKrP9cmsoYhNeSOIexgpEA/vry5zyEIuY2NxYg/B2jY2Gh0MgsR
HfS0psN5aZf/ZCy+X4ieLuUflgcwm/uX7mbNTfPWBN1Tcm0qK3ZnRVu1a6K2
E0J8vOTrIrm1m/ciqrHpzezCzhkDYIuxgiIOyL0Das7QimuImwKvzI7uY0IV
qEPII3VnfEM23BH13xVz1KyGZdl/JQBaPIWIrWgyxzcNu+kZ5x22kITesp0H
cPsvBSXkvcOT1kJRpc8VNoCe4TzvRWTwieY4DZBTn295OD0oHgTqXp2zLzCs
I+IoDLUBVHRXYkYMu0EjP6E+ibJRVbC/swdv0uaGbkzDQftlS69TypLtouPK
Yb+D6O5uBDYQ3jgmvggEoMUBj8Ts6tod7hKX8lbZDf9KRZeymzV8IHT6cx27
AuV4b7ObIdwayCzLiQqc6DyojGItS2oDx6t54iNhk1gluc4sCI2UkZk8032r
OJ1kuq6TmwGQfV73VqlpQA5N+ohf92U7Jl3p1qGijEGO9RFdJQe/liFHH/Kc
NqsI0VA2i9jpQohlw7cU7rMW3DyMoDBdy+TnjBx9JoZ/7jD1OpR6m+qD6rPZ
I4JXYvOIRAr+AD0xKySamPrPVqPcdi0AMCIuFuIFmfDS2DWIlnDsO1nwygYz
XcfOS014iy+J0nvRcCgJ0YW4d6j3yXpFMRdYhZ1i4XIPx+Zh4jMFH64TsM8S
47pJXbtkuyDdVflnygpnCriNtHHXI8q0FDYPSiBGJhGngKpoGvwnFskOuH6R
7/yHgb71W1QskbJi+GAWOAnkt9xGP66HrN5nwtJ+7raiC4Wots/0Zx9c88p7
ah0VVVQStq0DpnBkw/qmYUdQA7o208kmRCfnbufOTis4xu/C/yqto2EJ73lB
1VTd2uyTaq4c1KVFc7Ha3XA2uW3yFprMF8ftWIXi1FNvZklEih0ZHBR9r/mK
337e91qLxGoHIiRwJyTiM9S+pKCYKODrjICQC7QH9KRxwTahEYJ6atgm586F
1IIKHv2nUbelNhsHww7HcXTsq+JgYVAyFO30gJcPlgl2pcmBrrLWzRAyWOyD
ubNoCP9Q8k3Zi9LtJOQ4aJY1wMsrZ08LxCx/KfdUkrZYBCuBBOWCbMami6Cc
kPqcQKH9Z9DkgeUlwnU0JXINOE80vrEqr4tcjlJYp5u6uYSChkgfSliNJFMU
x0nHiBIKq5KlzbmpioV+mlAtMIekrAoLakqx8BcYldlYcZ/SNjqswGRUF+dm
a6dxRvnblqpSitmCDWFr7lmwwtGE+HsZWIqAsxR7Mj52UybFG61vFp2Q/rXX
qkINonHVxVeanlLw2GqcbHquK8UA+u8Avmrp7i0bsCnt0fSEVHnTPQFUHABp
ofwB6NLBr4UagmYylc2fMGonSfbCyhReDfO8C4c4xR6HpNo3V2n4RexAzSG2
edfdlBRbYXNpzfXoRgaBLcwtR4fSq05bX4I9HDUbvsq2OkOHJYqwrI7eQeXc
jCdEfwXq/AIFZhwPN8+i9rprlFYotBqdQeGQKrY3FsTiHjgXRqHa+LglEM9D
ALbtgJX6k3Isq8bo0AmKjTw5Mdi1rl7gvXeNZUSy4wvGYdQNqd3HWi/S2A4+
IMnht/ziq/POkJWiStPW+e0lQcGe/luetKjXFkmbG2i1mjPGex9oqK00w6Zs
WhyKfz7f+qk+bj+U764YbQBDua6zkm79brRqLcCrOGvYRNZ2tXGALKbmb+R5
T/CQW5ea3wD6LqloGpqmdmm0PYtXQmdvmCgaagdI8IEdxKDOcy3f0VzgePHZ
TwhdybSR8LAAaS9kHplN9KkWvgORM7vowMAMm1TufBGTj8czz7Z/MEuYWPH7
2inaC88XdJjm1BxE9f8fcowyUvIKyMrXTUC9q4jbwtENcf0myKfRmAImTQeM
lzvxazS8oHkOCjEPI3BAlAF9+0MHWDzkLopEGv+vKG5XpZ0htDJkIz7quten
8nlRJ3p51jOKc2ytMtitSs3YJa9QlOesEiDNLbhQ6MS/MTDaMjkxknQgRUpM
UJb3cASFZzjfvux3SH0AeOw915z/NbAOQ0AzHse+FtcZO6ZsfSdDBzFOKr1T
ulZhHogzskvCMj82maokcf/28BsbPJMequSape7ckz9IcjDyzNixPIwpRIH0
68wQVu7IH1TrWZbMq5ii2TMTwdu1I6EjfDfLr/ELcdH1VWheNod4+TVJbn9L
cVxsh7Ud8VB3JJD+Giy1QUBNDKRD23EPY17ewqrCP5YTESMxcT3+xgU/VgZL
aivGNJc/JKK9gVvNdFa6wRy/U2CpSCUThBjai5jy70d/7+V3AEpcBNXB/cGE
eHuIvekJArHxan0ceK+4KVk6DIBsnFIp5amXZhmzrYFx6aooyU+I/FXLYD/f
McwsBr4FPTSBjjVbY28z77gH/rMpig6DBa2v+pjXiVudg1CAQzRK+CzmC7EZ
0FcKl5Xj2iD2fG75ne9L/euiFYLNxNtedO8BxPhZiZ5oCBxMCRiXvKTTZ19C
akLXcxLUHfm1qP/CWraSApJ1epdRlIZFFbOZNsPcqHq54F+N1pJkikWCJ+dA
0FxTCDV71DngQ9YAkrssup8g+HTr0CSlhSD/GPFDiywJNl8H1BofBiOy80Ee
x6i3gCo3X97vBlqIp09PMwiz7GiNHsqTDUewoXFRKIlRqOE3XEjsfd3ZQoYc
73aOPcmPEbcDyUK/KCGzB7oWQ2jtguQ2O+3Wm894XqpkYiOqbh8CGdbjPWn0
rNk7EbA+YPZdS+3ZzZoXBXFxjZmDlWFkJzNAhWBezqx+4suE+93p/HUG295P
1HgGJdkoEsMARM2mugQPC3ZdFmGiOj02GBUMcKGrwesIk9U1OT8/CxI+lMZA
VCmJ/JbnmLngjfbkNOhHxw9WS6SoYK8JK4VKC9Pd5UlNEiItGnl8tmJBJCGH
n6WzBVcuYXON8reXlNYyipKMEde6g29JAefG6wUKLPLk6COy0OOQv0w1tK5S
WgXzcRUTXhtm+6e2epDXk4M/9PghlXjvdAnUiAh+QhDeBGPUy3PwnPmD95pK
jhOyWuDeQ3rEBRpUwTDLLGhia67O4Ct5kKwZ9U6rUXrlSrlfC1xQAX7Qd0FA
AXxUC4LlWUjcpvcebbxix3G++H4zZVvd72xvNmd40vrIURdj66zAUdV0BwwC
eow3d96NV6eIW62LhuN+xeck5W+ZpapAWSIzMtMmMFVQkCa8YP2rzPiK37N9
A49O+fQfBf97Seetjoa0l8CKmMouhfnw04MCLrJUdItEQHA+sx6xOVkL1WNG
WOj8WqRlmAhukvg+FWtl8YoaZKOls/p1vIy5MeiRz3uwQsIIP+ddBCHtl/dI
JPrS2oTJqZZuRZsvufRuB6/AoSJwKTsFcCIxtQanVwHuABbXTzr33wI92gaS
qMR60PE2IcCjvZ755raEkx3PuW7aeWXiqEsZFk/jv46dQ+Pu7O2Sm8NKH8XW
svAWbPak0uAuqzhxpQQDxbg2f4GExXsh4hm03OGqxKialCv8PjDpN+/IUatp
Bd6n0tj9GyOQOZxZfMXiaBivGpkDeG4iN2XcmAs9dliGAcSSSGuZfI0ksPOr
A1J4PAYP6TZDXECmW/C8R7qWUX0wMt3kl08bkkvzTXKPCvgcyLuZ18PN8HL+
345piaHDbrhbfGFuK8A3IkSCG1KQZlqKXn0mW/pAhG3DHFqYGQ9o46ucEA1B
wSGLFX+7Arde//Ak3aYPLWUq2itASkB5Mki+MOd/u+LexPGpv9NL2yvyiF8W
Dg323Z1F9etpdKR9tIpIra0pB7N7j66Rp48eiOfV1CeIOx4ZvOt5bG7YhvFj
Fm3jyWPgQv0dCr5XfLETooGkh7z+YhpJvq0HF7SoTL77Wj9oCfMydRDWIGhZ
T6oDPeFVhQ/RWpX1aaE4FZmt9Qv9iIr1hWXxKn0TqB9cpPdf7/2KMSEhvn22
XquVjtokIdKcmY2QOY5ZX3uieKtjUB7l13Jvqghpe/eeuoZodOdcKbqLJ35i
YzO4vYA1qdE/NFAERouNP39joND8PVs3EjwK8ejQTp8t7XJqfiUilA/AfI/w
SpE72dAvyxkN+BbjhpkjYyH2SjgzCcydYcafolLpUeH+V8/9zN4QM7+/ocGG
kptH71JY6GKFCe6hKa2iAt98yur2iZwCQBv8kNuPaugT5AyzlUdCc0Q4biSC
icxkT5d7pO+PTPk4cjctyeSB/ugwkkLKGL9wp1CzbqoSxv8D8mL/H+gJSAIt
/GT5LfJbJFrPIkkuBFBDNZPiD0n9MdMllCCDJNzF+7O6uR1CLi/7Jkm5ooXJ
Cq9K/FCb13eRfTDzArQONbUHFF3OINa5XP3StROIgMq8DghkPtZdC+zeT2To
q86T8Q5FEGcL9oT/BmfII6gyUHr/cvp3am6vRN8nVFFLE+noJdLgvJbF5QL+
9vDq7R+8mhBAclzk0Tiw/WjaCkZZXpxxr18Oc+TQhisxmmsbPk64th15iGjt
L4LvpwrFfJsIup3bvweOUxz0bPybU8UKeLecg5hFQRWgqWgy+NAI8NTzyXar
x80rKe9pF0c5pTuGfv5HawFl8ES47dTo1ISBtMXTrnbI0i2W3AatooGzH6xj
v9Bt9U5RO7M21EE+WPg5K3yOzzy8+zzKU+IJLOQboITZMV/FVTRYdptaRPq3
9NoabbJVZXLCcPwCftTvxiVjRZnYDDHruUy1KQ9ywR33IcH9CMlcEa2fxsSn
fizMBqSiHvBUMx5/C7LZPG8fW9q6/QgGa+/TUmXWcvEeHZupjdx/ZR9c9HF7
I1x3Xd7SqWN18TfM4gxa0FKB9sX1xVHXj0JThz8ln1KqVGvBLMM/RM7/PTCi
iLn+un6uYjBLJ3P4sMLcap+Khiitf+TX+OpMHteVKkYhlJYq5cQw+LpNP46a
GiI8g2CAaYiQ4WkPufa4ngJCa/XPI2ZpgMAdTtnKa7SBwiUI1z0gqKQ7v+7v
vvIBuXqTLW6RngALaxUt/t2rsNd2abo+g00ICc7z1UopsU32kIKnYVuSt86c
TyR0+YHnJxDP/KZnmbcq+FLXz8HUXnRBKnJAi3s7VcRolPZdI8dvI7T8W/G8
o+U8auibAcgzv04vJIw0Izx7oxPzPY0wHNqULoYYB4YyFV7qyYwgU321LAWQ
LPWyOnUUUIsKLrjdn1werQRlpskigre5cE3fQkR6kVNjzsBYKD5JJH2KAD87
9KN7Av8jLs4jg+Gqit8ZeJqqgglA43nNumy5Qg5xBlGwBvFfulG5YbYBn8fe
bVVNHYXwwG04fdgmTA9l/u0CVxmU0X76xPj+hKkoTQZfvP0VmX/qSPpU0Z9a
lwGG32bMilfzlUf10BooYBFCxRVApk4VX+8Da8xv4yTVdr7lRzZBwNvB2KxT
vsPZLxWF8xn3QGINwk3qIlnEvMWL9FDhY/Bzpl5Cag71MWC60GLr24et2HQy
hsm1H+n+tuFL4xO2AWoTEDqXKoeYSEyisnkFn5kRlCjoJn4E3Ej5Fit9Z1hm
A4SZptnYtz/zY5Z4vIdhGqO7ASEmMrvDaJHONlnO508Op7A6c/XhSIpaW9Nu
yQhDrD+Wf7dUwdPQJfGMdcCXsOLXv5ToIxufiL/E/GL8fnbgFBKeWbFXp2sf
CVWw9Q1MKApa2E9anAIY4L50GvXb4vCW8rYOaMofqJQw4Uxdrc1uGa/WyUL7
q7JPsvY9Raft+MFqP8wVj3KPlqGToHNOLi9wHyPC25PswVcUGthOO7IwmpKe
OT/jF73kEKQ0yFHEdBtOyYYmGMl3SYiaTPOB0lzAlyHoY+iJ8gv/On7YKuQJ
xizSTNpnW2BbdGcf0sbJP0SYYCNl989xYS8oi6uD7uT7VnkypyELJ+PB/+8u
F2TOoQmpyBLiCxf7JmBPaNYd53VtiAMrZszaU/3YUnlEFXrG/YtI/DN4npw7
ELuZt/uDuhmzZzo6Xh89EY7yGXOqKRQMep5+hUZ4fkY2g2YVLVNc01q0Gan7
7mGXzMLZE7T8Qk5d22qTtOT0Au6QWTPAtak2/f3DmPC9kp3yLnVwyM73hwR+
LaOOhpBzsDtn3/BNno2dMU12JZLzwdKYCs0adl49Ty6R4j0ISZ2H3N842nGc
Ex0huALX7kotSYHDfQwuNpTIky3DILpYUoY0cM7VpHlRtrloMfPqzcg2k+3y
XPUkZ3fWYEAxyn/nt947j8CAGS7HQRkqmcJG2JReXfQwlwsji4BAFSzaCjH4
MM8QMHuYtTNmF1MfEw59NUQ0kr9LLBZlXWDAwG5JAUlcOkMNQ/a9Jdmk/7r2
Y45a6pRSvtzvigsqbc3Br8t146c6n/2+YZ69vunT2kFEa4qv9Wob9V8ewZVi
qN1+bob6opNKGCmIt//z6NfEq39+6Xa4atG9T9UjG9IY48KZxUUco43Tak3+
nobS6yV/h+jhCis2fg00058ygvj+iGDx7nGrXy9L5en6SvGzyXkQ/kDkL959
nuxHrnFwDXGnsEZH6oPzDbBehNcveFDf3rmcYlD5nOOiLDl6ujz4WG6uPlu3
JA1R0g2K5C/YEaLMlT0HAPXnqe998W6g27KYpLc9pIm6LeYHpwDnRTAt9QUf
fVJIf47TmPZOQjmQlPjTjeSmXQt5h593l0HPtyR+ZAZKhpNiuAOvyi8l3rol
bLCwjqSslaWlrFRsEyFHvam+wXh+LbQacYVpxbKuRk2NfdX4EPhNfCJrQjf/
yfc+YpYhjJqyhhok8NzGMmrAdLpHzZb+GZKl3Lv1dYAMlvaTMpseFeRnHhRh
XwaXihBXEC8gs6Tg2k+apA3HqMUGsp1T5AiJWN5CUifqX6x8OcoQtogwkvOM
dqd2Q3vFAadw/SIKaJWmupQZWrg8xTuLhI25raXyNo3c8dV/IFnK6xpt2R/A
zcDoPHy8VpDR9ry5CmjN96VQ0W4eFIomfqA8ZVgMeiR6ir9MwyjRNwPHgy0l
Lg+LqABjGrylWch9vd9KLoFdmrBy57u6EpDTvwHudDlmeEdE+x+pHCM70OzX
BRX6NYPuPzZNjLpomCMuwM4fP9+nPHAa1hhG3mw1G+tmedaV7GWAPPz5oMQc
x+k0JlkckpHkLhV6c6mpqeFzTIgNelvT5EQ7cyZ1Ln2jndri+dKaUzF6OsyX
Rr5RM6I8zI+7Z37NahyX4poB8uS+dAIPJR1DDBCXpO20dNfnJgcZE7R/tGqw
THdXEe/quYYTn3/8qpHltyHcW+KVjb3WQnGRIDlLgy1vhrCy1FoLpryHIa04
x67JdgGKjZc0x51yW1YyW0vW9j4/O8eeWOkhXtf34SaIzx424HTuUIPQnErV
rvhRJJ+4oaUJcQLPMm+zrGUPVQvnv+E80HG9NLtvJ8sthmgAORPjIOncURZK
35iSWFjJ0x4/PvhknBZATdR9FrHK7ZgBwT5biRjtnvi9XjmTccgD6iluphtp
sEnO8vboDMmojwqhe/tVNH/Q6xXrvlmfWiN5Ry8XJwEzIuKtjhmawtoqcEEx
fvNG58aanDYZzFZNkQq93MnREVofpHD8GnV1SPAcJ++tVdC+qPQrh5juWvtV
RG2mJQXUpExBXRfR5MzOgoo9EaFG4T5bw/m/WmkjNcQ+n91ald5H1ZM3gOL0
E9UVo0MqnpEJkaDnwaUdD+IaHlM4SDveUFjZgCgyN9fUPFoCT6QGvti4cWYP
Ak7dS3+8ymHNS6cHDfEVr8JVLr+AxhmgfFz3kSl7GCOc9mJN2X0v3UBk/eaj
ekT5y9u21AFn5HCr+IH5lyvTl6DdtlLzrv4c3wcyO+6xGec0EXf4hlcysk+L
r5Fkyz5PWCQt+9hL7cO9soCxOyQ9oBDwBhzNQ1NdvjKDG19b00I+iJW04HGL
v1BERvC+ZJXFULXPrbazK/loep8372ZkWLTuWi8ljC5sR2Xf7K5N8mAFTvkf
ctyivEda1RohbzlB0eBCuylyrokhr1j9wtODa59cQF7kJz1ioYCag/iKakQ3
GpmQN4hkUcFy0JTRm3jIpKwRvJO1DUe76YKi6XHB9rguVaEckQGbuX/mf6TA
bKKATnp1CmJreFL3xTMEYqvZUAJyhhcZnVE74PGvkLMm4tPdugibL5zpdzMm
IOKp0wMdF5ggqQm9wo5C6USmtSgCi2L5rtuAi2UnLWnECbZQKkufMjqhwgDx
gzkvj96MfQi4kKABCn/9/PnFTUFYwdHVlFjDdSuvJ9PRu2NF1wLhCl0jN5/+
Qtsr5XYD4hedBh0kD8lo3LOFElmU43QgmvdEqUFzWn0QmsTTGniHohFUT/oD
445bV43F0eMqx3IqnGh0sIIqQfTz2tqsyDRk0iV+zChl+Hcg0CH0lmTBMzvG
lz3cXKPZYW5lk9hUKTTFlnG4eKmGb27I6VIAC9aF9GGKOf90D2kfS4/YY2pQ
FiLcz6p/1UDQSSwPTEqs8Y2Y8pJxfty3UcY1fqAG994YOksC49MlCGGdFB7k
foW4Iihh2CEsevmt9SOxtoyp5lZ+kliPOkBvgXD8TyQy0ajEfsccctIB5HmO
K/k0VE5v8tUAOerPFs06i/4fWgjyy1rQ07fdml0zkF7aQ+imwB+tDtqebNN+
FY8UMbEeedpNUaCjIvWDtPDCkCup8mHJLqof4aiHp/Ewt7SpiPTqlrBLrlNX
cq9alxnr63EqH1hB/aNnLn2wg+QAro+P/6XW6zFAMsZpD0Hz7YXy+6UtXt4Y
JuwvkqECziL05cCJIwl7yHt81mWFiCeEl0Vjqm+zMbGppA+XOp/1y7VRM9Lj
vjf2EcCaVXkTBhQff5bPgHMnOZtR+OtGRn5IeDElEeu8ZlzkkQeS8c1Q/Ew7
isjduVIjuQxxNIXKpolOeSJVKTh3qaAA/Ymm4nGRAUDEeWF+Q9RUvvADEWxG
VCRfVqrmIgHJjrT70avTvk9AtE7/QuYck0mYnH/561l2LjhZsDwT9konDQeX
QHF4xoqNupB7yItqkX8Wak0HFNLkoGvBXs2+ZwGDIHf14SllSfXLwGUqwWs4
wls2jsSjBp6SkuWwwMzTJO5lHRFhzsfjRlhmAR+0g5xYb0Xbm1ml9B8L6lHe
ZWou277VUObRzqyL+Ktd5s13IMiBtB962TpERktiSlgKMYNdtKbhvuMRabDl
x7S93krXSgZKzBle7JFxU2IzGXVcQ7TX6ekMiEjYG45RQqL/s7On+72ONRPG
W09kNXGcLDAaovAMoOIxFKnaEVM0gAzqIGoKkWEmACpZTSZC2G2YSlnXP2wP
yTF7lh0lWO/WNag1vFASWW2pQEhkF8mWAco5iZwDqNlcrYcX5Hm3l1EyYfg3
2Za0N3IaYhCK6PiARcR3YL0Tdnd8d/cFd/zRBblettoCwethMJsR6Iv4gUUz
IrlshBY6AiN4kGTZ+aivybMZ1rhNEXwuJG7ro5DeQdYtuWbLGhPjbA2cH3Z7
Qk+h7K+B/d/gwOk/NtX08hOGjj2Q99UfVJz4RL/zJekv+UBUwXTmgM5YTeBh
QgLX7eoRZIihtKsN7qp8QIZNU3zX+GCf95Vy5wAXKQPbrpF5K+CJJA+GL0Hs
0p/h7hItGya3TFTId2DZTpDvODPAiMC+unb62v3v/S3T08JdEj/iEmMEO2us
UoEVZSPFcseBB3Fjqj+AwqKAgdDhYoApWWlyKPU2lV+DLMDh6bgmNIZrreo9
7bZ8sECGGNgNYYB4cUr63xjGR2Wz2LNVd8kO2uYasV0/UcXmbUl4uLi87lRU
T1xBJvmHaW4EECpv+2kMirBu+hm5n7QDaOtMTNX0TevT4gTZLZnTd9dl2Bgk
6ySkgeW3uMKbzJk/FzVnp7c/YdoWtvEko99JYr4GMuACN4fAYDaEUgHz6Cgd
hSA2h7aECllKCHkJk2aciULRL5bCdb+RkktDb3g2kvaqeG2ZUTnolprVvFju
awVqU5qsezwtwYfXynN8MMjjA3KUcvZKLNZRdNVLii+zgMEcg0nMPyy2HBSH
vuLKKdx985juvi00D7HeuZx/acn6Xu5PhM8Dggq+m9PUKPqFdIrynoXor1xq
yN2FMm1ZZQ2OyT8zih4FmNbhpRAHXRLTYx8NXUWiUFisurJq8IedPotwa3yJ
TLrIHYB6QgJxR/KQw6IhslGU4w1cCoecxJE+iaMkOqmIL5CPbbc8/z30klHe
QM9MuQmFyfRrctfTZ0HCMtBszOZ7Iv24UgM+kTIs6WcMrrCb5Akn2Vx88irw
uxubldfaLLHVqKANkUEI1ZOD+0MuznH5P39TwMbcki1dNQFDEwaRLmHEgK3r
omRnBoAiktDHmxbrQqzOjgxn1Z8vlcbahE7e/P7B3NdnguG66E+RdojlZ7a5
XXHq42UeQIZOz+dIn6FcaAC7IFK3xdXwfLMnqpLlTMH9DV3JjdqUypzGk7i4
hUaJazmyl2x3TPK/XAzjYytw/LXUC+zNhNjf1IbdsmoLooKYH5+fK1jf1ZVd
VEyf16ULm9HLpQVJPkM/iLZzYQmAeScQrUfz2qDEpri2Lx64lOuDD56b8ajd
TcjO6kNb0agEKQezpkBkCesGSjbc2u7HdNGIoNLRDeQpC2yZpLifEQSHCm9s
GX82KpY92RCvV+cUvNyYmxk7lhrO7REsZ98MmHWUJa54ICU8+BZdi/aR2EpJ
vm2vT7j1QiEzzBfsCIFoCKKYlmnqCDedzioSeSwGwkFkfH9mZ5z5/ec0Ppt2
+Gcx2z+xuiAKc0axHiw8tg8EDsiPRdTZ1ivhmhteF6mCD6JkknHeLcx243Dx
YPySBwT0XQqEvRmTuFAc5c80HMLJ/ptFlBDI1MkYOnWe2FsZKROWXpAUbKch
iogqQjR5CwvYBTYi3Cz67uTH84sC4ay2wxfZ+gC4wBPO9IhwCRJT6oYQ+sEj
s6p+gCs/OZW38mli8YZwvkIrEpwIl1MET74MXkgA6D12E+Bf+g6s0zpcTd0V
JTnOZlSNegsG7tvk8uTembV+kGMpqJssGTAssfCEWJiow8lmXlvaQKlQtjBF
dJILe/9YeSpnnp29WJw6SaEIAuejb9RytTw5eawX1SD+y1FkBXNdqj4rl1af
RzWZe/tABY5xfJAJhW2y7be+Zkrr+wghlQDpc5zPW3wZXV3ohFyqS5dawmrS
vdRXaUKoBkcH14ujPmyH1TT341PRrw8ddn47w6YB8lnNmwL0FYNHH7fKferz
O4mklAOO5ui9P4/b1N6aKfLFkh8gYjwlLRLrPfDnxaaVYqP0HTKeQLdN6/hj
kngjfjt0xJAIqdnoD/IFkwKJiPZqzjZbz9SQ+G69gqXaTk1+D5Yl2S4Um4Su
knbDchLI6FL22nZd6u6EIWBLvKeHsiGg/w6DETyU5srvb7coi+cZ7xA/P9/p
n+4ceFYGsvYT/er3THHnMTycBvlFsC0QKLZvx1cqf3FBjUJ2sW2OxF2n9tPv
pfvWYe5zv/V6bfJLW82EWzLCPJZ5B12vsj54Y1UhSkcDS9sYaS/Kl0OLxs2h
1SR1lRo25sEuirpUSrsTks+SDLUYHC2SLWbJQwq/C/p/MNN5ZTnPUyen8uUp
muPZZEJSFyHcgIaJJvIGOdV6AnoZIoSP3oRCisXjVHrR4rKUj4/WOcv2U2bP
Z01z9h1wEWST4zAMo4FALR/wO6o8Oz+7yg4NpbprlBFE5cXspB14McsF3DM7
lPKeGaAzJO+IvqgGUGwROaNrMERGIJS0mZ7NIS85k9sgH4SBJuHLeeVYhBci
QGBaq5jR90Do8vgh7H5bqRQrDTn1hwdMzPLwVpt9IYe7zTS1eV0kb9Jtnj1Y
8pcaPtGhcVbcYleeZ6vMZL3qHnPwYpI9n3VM5puQPWShi7XRJTGd07Op5Kim
62qzQe98XmX4OMeXAviFvLuNEXT2Cdkf5eDQk5/LDynkMnI+mi1qgivx6d4x
YmxuhjzNHuvj7o9mFSZXku/d/ysOzRP0TgumdT4wx0jSC3t1PjrZ3fjZN6NQ
ldFz6OOPp+CFx8oZwwthLNr+B3YWyIruNI2wp/gCMcjajheWIEiPHtCTDWn/
iZtxOzyuQmIaVCdYGjNN5X5Jl7j9jMFCuCl6w7K6fvWHeSc11mT3p+eiOi/F
gp7p+bF76dVHc7S8mfZHYU1/WIXcMrmMn01WRxIyTQkFQWo0pu9zaAVag9wC
xZ/VvQMz2qWXiLGfRLVnz0sQnLa5LJa3/YjEJa4WO1bKemca+F/vN4D+ZeWV
BHl9TqyAMj8qhBy2sHt3ARB2NFIpKhmALMP9R6L3JVJKThVrRHxuM7lUITfL
pU5TLDv1bC/lTTPqwIyv6Hrif+IhmmAVckBxAzPxfxL0ZM48EyWHD6qcSAk9
3dpjYNpPiuF+jLt1qLhaQHdqTJgMPfEcBRbEjdPVCK98z2HurbGg+sVvBqGg
9jccf1ix/+JFmaYg8PgVZ6hbCTTG9TfZZz5m4sNdO7qdzmJvWY3WnygN7fZo
SXa+k/YIrtfXRzNkDCdh2fUaWrTe0+ZOr56X9apVWddp2bWN7VLVa8+igiCL
y29rrx9Dd9n2XauU9fKT6jE+gxANtL9Orxo6td7sAKcnVBOXvXf4LUWFdE3M
wtu2IWME/5UoF9uHcerHZ6pDn2mO+7fOKkdA1Y8aKyCA/AMKj6gk5bSYT6dk
ScAgtn2tblWULiH/oTNQMpGLiQsfUiNik42/KgHhPQAAInX5zMUSvZGAu8Fj
OYL3bFzG80rVcwYMPiiVjAofm7ZAr/GS/gyxHRJ9IQXI/lqJImNAOhZx3yvS
uIQFkRqJbyiKEdbA6x0FLcz+JOuiwwstDaFI3cCO2yaMy18UspHA+6Cjo2hp
OPD1yzJJVfFItci1KblfpEFIh1g6Opbo2thY/RCN2i9f0THCDU0YJo4LCBn1
fw4qIZzNfutJQmW7bJ3i1+9umIjIuNjvD+jHUbI8JFSMiIHcqUjET6AX9wwt
o3+e4OE0o/YI3imbgmdDwtMNGgRhOdZdH5LgAPw7I8xDVoKrH/KzwfJ0jniV
pmV8gF09RcCQC6UEQnbb5UD5Z+1Zt+DFUJTBzWlbTHOF3T9fGSGKu8l07F2V
a6+ecYUI1u5odamQVNVMZ7qTXRzIVmRBpEBX/8cHFhQm+1081G5Nq7DA0g7K
tOCj1FFv4KRDz2FS5xzXLJzXFoAZ3Kl20PodvoyENXDZJ6rXL/nf13hXpMEV
DeKFo8IaEjeRbActIw3gpFyr0YyNIoOImswrT6lt4yCLffDc4l9Z4lVQU6iU
CfVJBbWC7Ie2xEcnYG1Nlxh7uh9Hnbl8D+IVcV+bE70xSxCNt3+zFWtis4S6
VeXFAvsutuONRqi2a2orDFTl4l/QnH1ehe2oulPnCdsSFD/KEKmMkZ1a3Z5w
kfzmigMZu27qiTkXzuO8mkzfq7isPxSJSW/3OYqm/HSDlC+2dzWH1F6Mf0wA
j8ri6RkjkUrW78ijgRcnnUIiTFjMe4IYEPLYcG0myaLA+4KTotJe5s5WWirL
ycU5gAL/x3btLo/uXjs2y39rjlKKlPtFHg47NtBjjAvLLrs9pY2LxvlvamCW
hBSm4ehqveggEHfpn5XQOQY1qELYlpdMseY2f2v+frzWdbmRdE32plXSJGGk
MbbA6mP+u3HCJgUmR75C3Ki4LZI0YpslnDyQwIk2LdLNzPvB6hKRC66NYi6N
rq/lu4s8Gs8+foAHeTb78AY5zbAPWHpWiPfklLFdZ3WTCYG+rMEhCzIGQ2Kx
nRglqmYeikY+vONoxRrwXvmDKaM7h1EKuDvYnHgw7/xrkRwXdO39A2thfcXr
b1wU9ilKLzyhEJh3EqBoUyVVXqwMO8KKVC2BGe37rCwDDJtMJPAA096GlQgX
XX+51MWMUElWL+vskdYkPyH5g/dM/Ms81OgzXvrLKS/RKFl9EtVci9W9gGcc
K4trvlwFxkV9jHrHIa1r/lCHU0CQqP/sSzfyLTZmeB97V8JnCw2EVeFLjfNI
7AQGfSIErnIFnGPOKIemoT0dIwz4ZNPGXHVj6AYhBoaPaW1/C8L8LceX0w1T
U89EzwYJn2PdW3++h1ObpkNYOOZq64kc8NjH1LK2aZI5QtxuSTLmuuSISAbM
W7AyDFOF09fbwaJf73o1d0RfQ5JcHY5C2YAUGI5kgJ2fJCXe7FMeQfPM1z8d
GAuM8C25/rYc1uz/7gWK4vqkAh8cn9reMIqrrHHH7i9hWFGYtMVZr/ewMlag
3MxNa9C7xMLnH9SL8IeifT8X7lGOL9jLj9uxcjwTjeIGHk7+BBIwjV/Q23sD
ZcU7cMNO8cRUFxKKfz8kUrf/5co/ZajZog34rtrAvxZ0Dvlp12nwAB5U+P/D
ynDA6OOkQVts4nz1uHjsXKHjPz2Bzy+xWWrxXypR6ALvAS6QqvlHvynq9Dnz
Vma9cR2XQkUDt7mNq8LBfVXUbRyyMdFl9ApV54BnxdgtID14EeBcFjV0IhJp
2z0MVUhLPmDjE81oYwHWpbD4ROo4FVHe3SDHpCLzyIY+FCnsive+YtV/ZnbK
wvvBMoJk0xiT3KzWTNQ0fi+fOy+rWL+ZmJ0RFD9yV0VcxEY3MKHjiz4SE+uF
HXQHYuqeLQ8h2/41+NU/qVOlnKZ7sN/SchsVFNG5dnVugaSeSJJcxEu7CTlA
f++NAv+uZWV/y75ajrvie5jVEVFc2ugQMMZGXT8G/Si6LrbmWp6MP0+NB8l/
hCGhAo+mclRTSbHc/jzKrabGzlKYiE6Hv17MGbo3rFyH7V7M+5lqwTeVLSth
6MqvNWRea6hJi0bzHZ4JlkSyQxc056qAN7suTc0WoZ5Z4vgu3u4aw6YQzM+a
WDcHtRn2y+lqbgiC/fMUGVaeJ3Z44D9QZ23RZdPzrzRkUBoBoxqtTlEEy6SY
U7zcgoZFQF3VCDw9jj/a0fDCM7ZoNQpxO4yRHoxvjj1mNOME1LTQF/uD6/d/
WSalNijW5JLYV4WWcqxkhh+VtbP3Ft+ElWVsnEdGMP5o3OZrVLdo0M2p0dnH
QdyI89ZtTSb02FlkZKThIgoFeNs4/PDwjbmZV5yNIXHguiArrq7nWS3im8UV
da8uimyjuXVf2XpHcMDCOve1XO4n3A/FRC0FOJgRrPcIEyqUanGIo1rBVMAw
Slj0Of4gixqQsBtq52dkXaSrtHkSjeCCrDEQiM0HwPJ+mgXkytvklnFQX0Gl
iKylD9aJoPzIw3LWhmSFWf8jGUu6JtCscd/+iHeX/F8auqj9Mzmsn98WsLo5
yOIu7uziV1/czFKACMpiKxTcRba8Z7hLkxpJOOr03L2P4Z2Z/2WDXFN3tWku
xcYS8FVk0j5xSdkKZVVxMQgc4CRyhT3EkX1wWhFqJ7gCAMGKSlyI+rOmyxHp
qLDjmdBDAuDyYzICVuvMN4LaPew9JWQR5ybWsnobh7wSiZkzD8+UkWkYV8QS
yZBnCfT6bcM/Z83jazhMSYiPg4BVfv5uB1nLvkQ5xoyULyBDne2dWRTFIO68
10PSqVKX3GUq8SW0kbyhWR0JXrEeJHzBZvNawfwpWwWKlsjV53fa+8yaz1n3
dONSDzezxRaFp01ToYLsSS64M4szfiGvhGdpag+RKhPlSEoDzk9jj99ILYXr
Aqb8e8zk4238JLTMJv8wPAK6p+2C8CwjwAi3omU5z/39fBp82dXhnt2OgoCo
cLRvI+yMgXyDp50rnpE60koyDW8rl/yEru0lB4t0cINsm/oCtMDWkbp25ChL
rfsImk1E/U4/SEV6mHG85doLpHLX/9j6rthWXryWhacOSOm3YGRFxyWijemb
Ql5TIU4e35N2f5MughKotbXCy0pDrUSyBz/8F7ztDW6eWCg9rK7uXKMNGp/5
NXxUrJgP/B/9eW74KP3V1RpPqcQ2b1w/5Lt2oWn5J79Dc1ddPcfEB7QVtzgl
oWCzwVua/PLJhYC+WL2to4Yx4qNbdsIeLN7gENWRQ+PnK8gnJnfpLyL+1Woc
3Vxtj1lmJ+CLGtI1N64x9rjr4WHhGLwLtVcSBAJ0qkOBcKybe3weaqDXTwfK
yVmf+qNDe4bJI7CqazGNHjkeENovdwsndXt36OX3BexX9wthn+2QITsh2+B7
/nzLUO87zZxyjJB762NqgRZUDonzplwVMUhIGIkDD1cvtysAK4JEpj6waGe1
uUBauvqRrB4pKrYdNp+es6Uz/byDpdwORpdIz6ZDZgIrXX+w1VJBAqwk2I8Z
GMRusXa+d5EA2o8rpdunJXJIfvUMGMMVP53gUbsN0zefrg3osoWPYXNfbadx
EII9kkKmLyy0Azhw+PGzBvef06YySi9hFU9WAK6UBwRPoqdq6JV/CmwsOtSD
4WWlMw0ZFhQ6JfAs0RSBedB/vTZs09+IQ8SekpO25DuXs0C6c3riRq4OnDBM
g0lxF92RrxUn3wlP4DXgB9vGGf0OcEevNdReCbNAlo+cDEhgkFEjJ6q80dcz
2bTgBKybkMijjgcLs/5jaDebWu+D22EiYHnr9cTV+86uZSCExBGZzmPV6v9m
ilUAa0g++cLB+VHxj54wGwgdpWiSeMuauyZJg4kLjAI1obA5wb0sz22wo+qC
kxSTvbAto5xbiAXa0+p12/C2twKdEUC0DCoEB4yOJp9dMZv/fz11cInjBuz9
gJquqocGoSCdz8HEcERN8LLwpW+cColOghbIlovxCesl2wzR7bA0tYJyVgPQ
IYpvOWoeo4OU4ScT86EhsEI/oXS+6w5YDd0SScx09rkbhD3PePsrVX0v6DP2
Qo9V1PG+cvjSq1jpodmlV000/DHRgaTB5P/moHFKw366CXB6RlEZr4pq37lN
i+Mphxpu0pEGQqYVlUYwGII3ZfYCdPD2ZZu7PM1SlGifYmabUPBwhHxxw45B
IO34gPX03v3quNiYry6WC4VERoTv6PnR37KjIXPz/Wj7NbXvx+pi53uhw16T
cdo/tiQe+3d2JEQIi6JgTcZHBOfuk1xuoSdertVXfrgGvJVe0EIfyvwz14vv
WiUpn+1QVjv7sQ7crNwgGiq42QEqtH7Wz/Rk6b87q8Q//t6JqWS/1vccFoXD
fT+dUXVhVBUj9VqFBWbhBfcLP0PRTa9GVbO84iTDJOE+8GBdRHf8F/EC1ZHr
Z6Kf3Zngtd40kujpj6PsuzGGHUQv05j6X31KdxoVas9L9nV2SX+8nKrT3SLT
Ne6jFrW/bFSIrkFrkkM1UrpsqGgzkUD3jkHYX/yms0Ejg78mNitwHQ1oZLn7
y31Zi0cq5064K4r6akwsX5W+DkOMSpqAh+5wCkNkWK35QA+7iC8DLDsMA6Rh
c+WMpqUfg13q1/HznenKGYFCs63XIB0Nr9agKAapYgKq6QRiNdO47anRZhv+
OOKFIW4RvxEnNMzMN+o46zXx19DdrpCQdHXeFyQojqVThcJZTolEatyvLdSU
JYIY0PC7jQx0bTvd9vMQLj3MFA34+El+dTN3HyeMQ0kOvHgDxFKzD7Fh95uB
nYozV/KCPRybpilj4mKJkJ1EyHDE4h7vzWXfGHcvZmvF1naBORU+UnY8OE1N
BVqCCCvhABHu9qrMJP1H+80oh+pjs9dyS/GAU+rizNgoXMG4Be4mp7BlRZhk
+kqk1rc9RQBVnIwV1t3xaY57shg6PTkuVgTklx5OqOtkPJHrtxneXqBW9hJ5
Ga4eY0MzaU5XHIFpK2vlrDxnprOnVltWTmnahFCxKD6UCNOWAXbAOFGqT9fi
jadMY0YiaIoCcMxFcGuj4abkpN6QhxwNgzcPPu1GvM32KDa2ZyjfXuupZFG/
FIS2QygHtj5kqvEU+5U/Wu+TbeOl46cO4Z50FsHjkyGCGYk+uoGrFLDXyC1r
LHB36LgqeOyki5So8CGf26mV9hTZlpNr96jvY9KR3LnnPTAMcZGZ3B38aeDO
gi3/T69W9KsoPiveyFbBkVx7MP2QV6QS/Vnw/ORDCavpP5tsJ3bAiJdHWT1Y
ewcsudh4DI8mdUWoT4NmbHAdLfJT08FPFLTTGiKkinOcGzPaEc0KoE6KsEge
hQ5s0za1piGJHSZ2L34W97aAwa56TILmGzwg5V39T2mzCueUBV+KpQsqsrZe
4iKHAUj1n86d466oOar+aBJa8aiB8GN9NqHS4sQqXIMhLkg63/LXxbqSxLJK
T9IIHBX+oD3IWzD8lFmbUTvrCaP8P7QeSGK50sRfahZ7C0rNRt+5e9wYRSOp
k1qopH0QhLwntZC5Z2/ITujko2fMiXoNsbmJnR+7DFu1V2x88zF/V0s1/Tj1
Vwqj8HRz6TDiLC/yJMzNVO3JtE+M7kNR/ZO/TdSHOYWhUvUWpxqArKpjF2nV
g4OpoSYk9eieeWpLyPpyk/0lemFbyn9SExdYiY/l5gqwRfv95Rk4oMSdoiSl
9clFMjMbJ+4mkM8O5vnKhaCRp1d3I2C4Q7cd2YTDAdeM0DQxdtY3K7Zv8ck7
am4u9WGZ96X1vTtPVMIlvygtl4Ol0N3hcdsMG1gcR6lzqrjZ+RBm6tmkJLGc
wp1nh+NzraU15wgfJpbrwq/fvxsfiWjWqADw6ZM0QpizFMKdCzyQlObGVl+M
614Lpbw5q9MGOlOM5iHqajdrcQF83X3aXW/trsWoJOh10EXAIOiqKVGwK/u9
7HqTz2+fqy0LFPijZKbPK1Q57MzH8ljXRIxooIw6YHexIiRTeLwqAbWaA5JC
ko/nnRd7EfIkaIuO2sQJfzn71XMEt7lM3BfqQ6XqFmvATTFGe+5RmZXGgz7H
53jRKk/a2DBy71CD8pWkJWNCLjRwWoND0174GZcXy9ulVakTaihE8nocA3bN
fYT/+vOWROqQReW2tL8zrVrIDRsFFv+9twPHpKhuDh9wHgrOEPk9gTE8q0P/
siLZauyWAoIR3oQxDC6JnTjObHuHFF81Q+horrAjEMg09HnTKJc1PlbPTR4S
MmHdVexbatVofIRl6ezfkqMyvAb7jum8HfMsw3pqrULq4To7kyajHtHLZS+p
9GvM2weow4+j/Hzzj2D01cmfjCx+kWk+rULV/Zw7TjK2td+BJsdOf/vWhZ6B
dBFvLZACS5V3/Mnhxal9FByrgEPW/QTh4kbrQDLwncGxXUiiCOu8f5nADUZC
aQoITCLc9Zl6V89vecb1uX6L0+bKjyIpx+96H+SwrJ5gLwJRhY1gMAtWcJub
iwuWu+wTxL3fXW3InPOEpyvsEN7sXUjN/0Nbj7IMZ0V2I/SjeJRFtr754HUK
qgw4J3swqFfWEZ9sk4XwfxdQ3+zZOX3woL7DhIx9Wfwuh5ATuN2hG0mlU1xi
seR7YpCeQ4+0ORMqKNUCXafifi41nm092ZSVSyg+ZlM/KAD38E07F/lxRq3M
kkDgqHVE+o6cvTa7inNcBN+tmbbvzKxrVV37JNqB8Z2BEIO+LQqVu+2VVzWL
aLtgne8CNNECbfBWMmRbceL1noO483j4vz18JI3mQShqDYY0js6yL14FqalZ
ZGA7hYJ3vN0ObdL0A7PQTaKCtp/m9BrOAloyRenIKjGcm4qi7JOeEMNn5wjj
Y6rFXbbgqp8fYvNmaG6dyblqtphYphQ7MkLTDZt7GFw96601UvuonG4grBrQ
nCdcVfh0/Sb7yMENv9vC3G7cXTOttqliqsOOX7wgJ32EN2FRI+5drhIu7ZLA
Ozls/u6ERb7MMI/GhujZ7JFWOeURhohnEwMeLedEjtF4x5gG6zhq+igKiMx3
8OUZAHJuxBKRKTTbOc5dRGNGmXsEwE4Jo/5wbztB958ljfOmt5PYEBrJRfIV
N2sVVGx9/XfPijievKWYDXGPS7FRAN+sWJyNf9DGxNk1NZlL7mQWrYZubNXe
a/nKYUuPHzB1GAhJ+Q05YnA6EO1vx7lGWUWbL5TCqLEp8uaEj9gCycqFobmD
mjBVFAHF37zGbrwpnnMCsWPpk9lYrqwEd7h09mLdinDG4iX1W0/vMZRxI+uR
ZKL3/7pKZoaxjlyOqVtQZwEd6cTpaUjpCekbUcYQeR8w5Uo2nad2OsIL+TAd
3S9p4eeov6Df/o0BJioRWchX64N3jDvM7gdDE9rV1cz6l2sBjx9IRcSqoO9z
9sZvsjHnrWkFMOqeXOmIiZhmqv5OoAqQ6BlQ+WZMOmh5TIPhmz5bKocvrUOH
NtO1UiCWec19N00Z0PMX2RiMxLvAfGyXcfnxr+gpCWet+sFGwNbUMsQgiioe
Wo6kozlQyL5wkSdbzhCJ2vL0k2qCdO7/5r6DeETihIKoxq4EgyFyd7WX3/ve
M2WgrXOSlvqdF+M1hbMnw/F8GzUSVGQhT2iLXPk3Y7JPtTcKW+fopTcxGmY6
GjFiPw6mZ06JiuMzEHvuzvxJWRkpQVIWLnwh3smx/tr2k7eyZeAPklcAREPC
WOhY7dly3A8PCov7q0pohC4On97MdwW9pPd18K8IVHbA0hq11OSa61GJ8Ue3
W12k5HHVGxUDiP76l2vnkKgf74IThjSwU87MUd5DEYUDA/9IVhXiV1xW1CAV
/CwN9IkGmZ+n498nG6C8hEscqHgPRS7tHXpXqDT+THJqVX5fZT1LzrR5F7x1
ay2G30rmHoGp5sKV4hm/sBiw3J4JQkzOckFkvGq+eCfWNyjSNSlR5A2xCRIG
rbHRqebEP2RZLSOwBsZWT6fd3TZLYaJaeuuykNLErm2NLVz/ry+iz4CpPIM/
UQSuq/Iz9DSOEQyAbZFye3x2wuVs7X/BlZl/qJcVABJzDY8QBT448t14G3yZ
HqvjixbmZlN+A5ZkArEA5yCVo+vpZZTKxFWNgMFXkC4N1ahgbnf2lxHsbvF7
XtRQ18d4mMLOIAW5BXPk7asAGHjQ+uY8H/Sl2UBYUGNv8phg1xuAzPcmAF6+
97T/GYC69+SRlm5cC4DjqJak/E1N2aSPpD7KC2UaNmg3ui8Pi6aEj6toJpHM
QCTWwbHUMiTpXvmyEx3e5KtMBMrqSzQpE4VlV27coVWQG6kLZTWqgeonhG+G
sD9AcyW9DIMWzvD9RZgkboZaKMgEZXNJLRKE2mlSODq8Rb0xP8yBwCMN79Qf
yCfHzCAtjNKtV4TOwBx0TT/04t0zhD0aBzeneJ4691fGfHjCVpIVdhCiewNi
j89mtOrRfWwDF6TD37bg62koS6A+cNdniZD9HmTrY3nk4rp8DxmUTz9GE7fk
w+Xb80sPI1+ieFbAkvtYHwksJT5xqpXwvou+o+UHkzBANBQAYnTk5KLYoRAZ
ZXZmFYDjcxL7ZewXQJL0sS8IvLVNE2Bv3rgCCeBwdRhXM5lnwlo88NDW0b7G
QNyb+9i+3WFD8VJJTTA9pVMzCoJgig5/vsqqrlk25+5QMN7UScmRf0qxQUz7
G6sipCxqS3j/RIgcXiVabgO8tqUL6wVtwsExeyz3wnO0fuveZMSEzito24h9
hyQ3LAYur1YGzHoV9t9Rmish8vUQ7vSPhs2g5PZl+YypWiQPqO0gCakZyaaw
XZ7K2Ph1jgaHgQKi33mmoC32K9X07yPUfY8VsfuynQsB7eruR+byeVbC4mMR
gcflD3X5dHnvgnwsLarbLdcNoS7plYUoEhlqQ2Ofp8o4itH5bncpp4+BTl2P
e/rg2/P+n1MXxyfSjw06zAJuiVaMyfuTHu+TqwDh4CRmxfs4sGwYNA9OVS6g
Kdj70DlMWZwX/y5nGGj9iXqSaN19hd5I2PsBWd87xk9pZGJr0EUo9vGKavTO
IygzqVbHN09mocz5Qms04KGHYAr17oSAn6fXdv9ojLeXkDHUEGFTCHEhjpvc
TyB2aMk1DnvtgtLPzlER+wXid+yQMBW27YrRiojyJXmNlB3JiXcbLx6CfsOY
J0M+ANnzROQMRp+5hcL+xEKRzorxDK+tmKFN7QbmOF+TkJVUtIL/bjZiV4WI
2RdwQMHM9ARTeCbx7KqU2OAZlnn6MZULVsHy9GYx6pB6xPlAAyVlCLbpNwQG
qZ/jSqWb7gLlCTAhLTiBJC1Y6xqtFR4NJdnqFS36z7Rgjq4n4mW4gVrLvbjG
TVwf+KW5MX+N1bbtKxb3oA10LYKvuKn3uHh+nFeVgGiRAfRf8YXXzGDzuJG0
JXYWB5cfOPSu/GHi/SDJzCm+i/rUjeLddF4qQyKGX3xq5wIfOfGSBBJbW6I+
8IBXz/bFnwMHCCT469MZmgHOyuwOXam7WUDT96Vbo8Vt9S/PfYLIy0Ymqjyr
sM97KeoURmV+R33fkAPbPR5NIM1WbbIFGF8aHWzdGo/9f9C8WsM2z9M4xr/K
HXVe65PlGZ9mQMfBH2duTGgAbegiCh8DtgWixsQ84M2lhaABxFmAKLcLs4rD
wCFZ5jXWGbSBsyOMG1uedP4HZX/wfMHZ3Au5ZcxFhR1bRuBBB7tQpjGOjL6h
vysbmYgL0UnGpzBbBDwykMGV2qnhqIscHLWxrz5bEBhJNs0xMGu6XDeDWUGH
j5+4sQqCzg+YbjioNO5KikrHnb5otX04Y7aT1q0hKtA1IsHWnAVNh+F395g5
qcv4b1ZGvGz50uQNj9CJm5PcVzIoKOaDkJ97p5KmDaWNI7z0oO5ju+ZD2vUi
x1Shpc6vOSNWuEQ7PRro2T/tPRQbaiEZ+RbeGTObSl8Ydm5wGbSYQMGqQlnd
A/YmJr/LViDu8qMDQ0oemmGIwohMJHcAX9krCu1ZBtnhITucAXQFKlkAgZjf
EkBcJDz2OSny9iqYoeR65q7UcwT/qMlGABcRoCIX97qN4g5C6t2tOD8h5OKQ
hMDICqqnXxHDDj0pDCttajs0Ypx18dxRqNsLpT9CyobgCN4n8QyDT0sXczEY
kDwb5kml30GDsLtFKIAN8xXkMoR0OK62QkjFsiSpVnK1fOSBWezO+y/V4R6T
G51k1F9iGCBaK/yvk0gVB/+sgS7R971wy2rDCJc8B46c3j4NHKHsj5ChVk0E
qXDtWlI8NOdxmDRYVAkRLEkTS2s6S5DJNf7aWy/nErIuyQA9qJPKhrpyVy73
bGsY1tATaAA7h3Y0++GFU08R7YShHegy20jM6rD+O8bUfAuZmW1p/47fi1ia
inlk7Xpt7a4FKI+U4NhOH6OPUIApH4rR2vbPo3zK3jlFQADyscvDMD1rrurW
5KCt8rYb6craZdVYlFCD+QtBMGUAR5j2kzjIKqNwYuPjsYMZmaJ3lzbTuloN
emXRwj1LDg1OB7PAmGMjZSW1UgSBKsSx5aVM2fnndJ9VwRkXUDQoqKscHl5n
RKo6mtYGKl2vJsm5Cczr2qw+F4eoKYP8Z6Y1hbq6GwaldrhrQeY98HuItvo+
mYT74SjdxFqOrKUnDPlQMWBwXKtbS3xlr7DVHkHfBgCIewC+ykhdDsUHmh51
zefIt2JynTLSEhdUM6imhZ6uPoYt6goSz4oCGlSPGwDR3MvpVtQZaKHLVF+D
DxcgfWf+tSxUZKdniTMzqzpKBTsvrDu8Cx3uP82ZRXZzOe2MYiol7Cgzv/ls
fk9sHScKp7pjR5ok6XACUm3qt9FXX3n2xGeuTdTvj81S1xyhAuev22G5Lf8b
hRSZdHZG+HoEE7+EJMJqvfuuf/oCm/r63qqJDmJw90nc6sv6gbqkstfbRpnl
7SqJJR0OvYYDRm7z7RVAHJAnjOl4n0Gca7KYVrpZYFrE9DeILE9Cb2QOcuKQ
2QDkIOgeSmDWDbV+6yrXX1/SNh85c+3WnEYgXT+dCHaq77P/CtWWvSswh1LD
aFm9Xjc1tsrfcJdnOqtOzVTXbEXFJ7vTvoRHnIKIHIUfdY2cF6O7Bth7N0bt
1jkTOVdaxFWJHVjTW9OMbVGsfEvTde7WfIKdBudKIGJTxRN4IHLBimp6akBz
iJkPNkz504Or2UbJ27FbikuYLbouE3TPMVJTzZPXKYuiMYcJQpaScvirjS8d
rQjguobaAmJFK7ddXdkUKy5iTClt9dzhvdIGcIYkW9k7wBr/hZ9HKOPpB2jD
cBGpPmhIvxFQxM5unv0roJAI42Oh27AZydS1dw6gTIsRCjOiE7Ovh1ojKDd+
QB48urYC/JtTjWhn9i2VpNCkZsZGEUzgYubKpsX4QyAwZgpAgBVZILCUkce0
dkmH2lG97OQe6fmMONSztDQ8XbjMmZ5Cs0RYN0K0V4GhX5ryqfwXRwHxrLZE
arBg1+bn4xERSfyiNB9QSI2c49GJf0Qh2M+gj5Ak7RwxgkZQR9shWOnRC+aJ
DyKcQC4pQa4vxxi92HJzqVrL0ZEFFnEXj1uCtZHx2vPEcN+PlJOeTKp0lcEn
N9N+G1VqOqLUZuPHMi9zSrOrddYHOJDtYQuDgVBGU4MK7F8D3ErE6xIR0jCN
+LLGQRCIXcLFNejoXXDY+cLPg5/Mwu4tvLbm0EIkRG2PvO4YN1znsU26S/g3
tse8HWih+u9kZkKkRoIVwyy+ybW2u03a9ELxKxVbsi8dbosV2VJL0tokF99M
DGm6dFTBYIlzy5eMcdx53kptA0CFVuJ9Shrh+tnRyCTxBe6j2TXVIi3x1C75
ligWq/B7TUwDas5vKMvsJ0eUhoXWGQyld3h1iCPKb1hsTuMY91EbYNNZEVmn
sfPACxxX31DziudRXvcHSnVEpmJHhiAkDJTJT/CHGeEPgV2DEyCCg5wyyVbE
9uEgGmtW5GietMXOKx0XU9ZF2Wf7UxF3zYDJRbPFC/IRz/yWgxgLHReRQo5x
UbQh2UspwyTrEjlzgMqOoAvJLr2wJ350tAJDqGsNibGygU7oyViW0lUPrcnF
stf+98rd3RWn2t60slPf9Jo0hvpSVA7dNgjffDaazF3Ps6cDRNfuY3rcWaoT
vtv1diERBGgWQvk4nPQqsPevP2KXhMUSFjoahkWygq29Bn3WYeZfiZHsNN6W
sIllXezsgkyE7yCjhoGXY57PKG7E9C9QzOOd96cgQjIK8ntoEBWmaBYf93TH
jZXNVgtjJ5URYBaKryF8cFzxHWhN45jkJddfWOR0480gpQ7smzGThfw03Hmr
ejuCelCVZzGfyIoFHORIcqldKuagqCtQ1sngPkH7CSlJtmgPsu5hkiFLu2ua
s0/bZTBJm7a5DecTyzZ36JBPajKUjPVe7Rx0hqiID9o3z5zadHE2JLGmOyvG
bazGJ7plzcEMDvOn2FwccArxK9qRBwkIdV4IuZVQKCiFgmxJB2c5BbZ0YXcu
FS7M2Tgk1ZVzRzHTXODQSpo9XVzXf8rTIBx8rtoN4yEBZbaBbXQk62iWzZz/
OvqEYS4nDydoF8Ek7YHpGRzeyyP1btG4qtmcmfz+lChpAjR4ykF8XATKb6f7
g1fb7vt1jL83xxYR6Hu/zPFuIS5SVT5JxvvPEIDk4XDq7uRW66DKhfNpTVkC
TFMAsxNnszhe+TvbJNVdHmoNAEtAufmbb+K4YliRyI5f7qOuynuQ3xjZjlMD
4++Nq0tn8VnbI8zC/WkOQl0KNuEOo5/QSLQmPQ8WlXXKTTP4T3Ty9DG6m/FY
KFsOcfCs13WwCXcAdATCjNpAbnWwUOfsm6h+o8CwUQrOEQC5cItUCYwIqiu4
mIGYADorEyLMvCBIw94cXnDMbwm+tQvjjCHwt4Dwmr3OCl6y7/xACOaCHLI8
NAVEqwR7FNjv3a2rsBxNLElapcxp+hUMpDCmBOIqZgg1Qkqh31OnU9LZnQ1v
xunG+naZ/jY4LecfZUDFAEzWHYCxV1kRLD5ZPBJQnkF5fkkr/teZiFNrBt9Z
HLcJYjy7uhHchKEp/Wbx3xLLoYxtk3+FckddGYK7/BmQaeZodaimHEnvkF7y
gMXHGdyYfDte9WhI1i9nULk8l56Ug/J2te5tbU/8kW+Jo8v6f5uOR5fKYOj1
imP0Fky2ZOzSUDrhM7VNLbJz634GI7AK4Yy4CT9BaKxEWj4krJdXLnz+WIwQ
PKKasOWWHOJIDBhuohou84f24kdQwK2D3Zi7vEWd67eG4YvixOC+j1bi/Trk
qGRUFMK8XyilqW7kjPuE09H4GLFK+0pyPHAxUhBSYUWIfAKCyqP68y/TWI3e
eSYUNvwzPSDyOc1ZKNIRaJu4kNJgvnOctONxpGnlh2m9gfZBaV85QUnP2w15
hAvDjBdnkthl8BKFzlT89fLOYYU9MUr9oE6aWttZARZMTb2gSes/qbuKQIPl
qCckYz9wJDoiuaYCL+rczhdEbAIqItm0dUbHcljfofMCZS9usk/EH390ovwR
tH31Thyppetge23okNRtQ+mnBE5lnxBa3HdSg2MTYsvkFzKkVlSIOF3pWvdk
EVzuaIqGWwE5IY0/Sz82bT1NaGTtGZYpuN/75834EI9u9vugukW8zeXeKgF5
eY7IP/G+ZV9cE4m0qCszsnccQV36D2G8upUohPWQ5CnYIvNkI+P6cdF+tAuu
8n7oUkUhhbbcD4tg/lK9ERJBpbHg04FemDavNw0ebl6K1ldAXRV5ULZ7C0KX
nqnugESGYVaHJ8YTxekI15snSNggq2YWjVlx1zkwjdJjwr0stMUbYd6ku6By
eNDjbpbilRkN6wf15uMc9OgpMdoRub1dZBCUCgL+zqhghPkj1NPtA8sXY72J
YwLzdeWiwIrgi+cYZx0B67APk8/Goj6yi9xdaJf5ZMSBd63JjR1WsbSkpx3s
5dDnRcuiueaIAE32JPCSL78tigV4FMvrK5rrDLLDECWFsxiUsV8x67q490p+
Ros0XTI5jx4xjb8C6TeT5qXi9SGGPchV1feK5c218O0MMDyxND0CmJ+5W4sY
si5kuMt2rS8oqOs3pzQqwnZmfEy/518IBaLbs/zGnACSUpgJOjzOdLk+JhWu
c2e6QLk8e1RSLY03dm/s9WyGoWwdx3Df0g7FS2gP7IWlZzb5hrAMUPm3yHVg
89UMAAgZkrpNxt2RkXSHFuUMo4VA8ec/wzzNJ1jy2PVDp+k3uuUvRkamgmj0
/dQ0pLABLVwUdCBc3NO2Fbbfgd6FOTz83Zgjm9SqrP1wwTkzjAYLpcfUQ0FB
t+K8JDFXw14ub6ylOv4RS8elSTSHoaBuUKLMuNYb0R6eROVYYtocrH7lX1B2
9uqsfo2ziIywQC7RZPKu713wDaF+GD9raRkMKeoT+nL7V6MpybUuVaKge5Lw
rYZTHHFWYETUKI/pTyuEoFNtSZDNLUyFnpOS3QkjvKGr8jGS0N+Pyw7okWjk
YkUcy1S4PuK/GTB07yDjsItnP1mzGsAIEM2mD/ZrOfFVRU4u3gEhz6Dnwvxn
9UUC0t9oypCGPFyPvgdYk6iD8EBB6/yY0X8Ymm+vKmK0RHzBIazBP0pBycm6
0z1r5TzvQiV3jqWTwnfuvsiaM/xJXAMK5PLXjGjQg9MIk6mN2jv/5aPejPYW
nHLq3aJVWE28wNOvE+eJHJJg5Fsil/PQ+e5qtp1X3ykJspfetZ0mckJ/kLe/
O0DR2ZlswRiU5rQeWlap7Igpt5+g170fg+XcbPzgTpd9KLF6/7TV2GY0BajQ
XtPUamKc8/Lg97IxkRoOLMk2y3VEDPNzX9wuaO7w4wzrAV9YyEDnqYivdNig
RZ3gKGiH29dRwEY3++Ec/ldngGslkvlUUaq7dOuVmmL9XFP5OVzWgwJP2CYh
LgO6cknSqo3wjvGSoozgHGd/VygIL/tkdjolR2T1U29c2vsd6uIhEDCf7dPx
fegw7XQcAqVVoCRaMt/9yoC3bMA3ObaXl/COLzG9NPwA/MPQSsz1NBxtxWhi
/YZCn+CYnnuk2Xi0ZpKljgHihKS8DkQCPGq0xaVwJ5JIVNM38c5DDkAF8cz6
aaqSp2o7h9kWQ1xUs3SAwpaxApQ2wnF6zZTQGtE0O4TfKfRIQg0d28zOKDFE
l3sLi11IGraZvMGWGWnuJVeNCuucDsvlkgCejpENbWJJqEWLi/7f6tdu4lvB
x10wRWpbaWNwhlimocQumZh7YCP3GaDyWrPrkfR2Sxst9XzQ8N7PX8DrFixw
yHc0REJ3x/OjaLLEJWAFrVHjJ1A0QzWtOzxDGwwZGfxEO7j8c6tKo695v9ke
Upkg+KxGy30JvxCJJVzree2tzeb0HNaSPJaM9fFEBWpouFoFDaNeFWavFajy
l+1dZuzdMWggbLDL5noozaUIQMKBE/84G1c4OwIFmB7XkCdhwBGarXwCKDcq
c9LLYaIPUdHsiVO0DLDoc1jaoP9c62KdNOU/KAxMcNAcDOhDOhOh7sgWvHJQ
PTlbyzNZ4w4FPiso3TZrwc5Dx7p7YEAZMkbl2SdWAv5eWQKXTcqG7RTX3Mi3
Q3ukh4ktZesVmc1PPQObUo1P6oFfJuga8OkRASGt11b0+N0VZLoxAw0v6r1S
T1C5Wh/a+KGGt8+nyk4hOHerxJNNfTNQ2a84FwqaJs07IXc51gUc5kuXGjUB
KCn8ZTk9oHUyyLkmAtLezfaXxdC379yw1+UjU4FPxpvvLhg1kn6VCYOhefTR
oDYVRdyApcZmLQLYaXxWdup+D0GBrBzFU1Iw5b3bmpfe05toWMGlhxC2Q0fe
9leCvTFF/MUnlD9Ijc6GFPgpW4mHam9AJIepZyaRfvcDItafSCqkheA/GPwG
KqzHJZ1IXmxSLq0/Vdh8JvlaTBaL74hdgbLg9ivQdkzThmeC3+lsGmHQRYoD
oPZW1BwbEPKgE/ffB6vuKhJ3pF/53GQ+J6IDPIWlqDkoHBgc0WxkfgFS6gyr
uDJY5dy9f2Z+bmfS4JiIYwrWQVWcou87CXZNRXFJWcax/IfBI+6nS3MgnRi0
k0X4/f0cTlQdBR+owblDLui2xpi5+bfIjPwUI+F2Ih77k8QazXQc0DYcrW9Y
x8yj33YhvWZWHDYQtO258aYjmaGMc17jRlub3sfSsTwVsNCfgBcIAeOkcnmT
w/3scrF6YzVg/4D8wWFeFimdNJmzhIaPf6/Vnep8wFVB9+2kCxdVjqin9Oyf
dhi+HM7c9NW9oxWNlyOZFUxCdkEgMM15kOWObTzn5NMvlrK8TNY3zHBmDS73
HZYW+VtRtzy8yOoDCngGq0zG2b8bOSbkmqPr+UQhMtB+QrqpQSRhyNuztT0o
HdlvQZjmMxBqD/u6PXeVF3KrXDw/9l+CKB0dzKCS0H9ZbKSik7fqNNmmy0rR
jmqSV1deJkgEqbk1qyswyK8riqzPYik3188eT1h6Vb1FnAgKh0yUcmNaTPed
nk1BXUFpeVoQNznlW4PDrpsMGq2Q77JuZLE2Gj7cqfCmLgnS9blhWIc8F8Bf
7jkP6RzGtSV8PdvVwory/O3yOrfvSPWAqdrXMJUg/lHNGgA8KbVarHmEPOYZ
KHnW/7+Ki7JBMOCxg8+tIwXIe2APK2CtiynSsMvgRQdGqZ4xazQhtCfQtcvI
7IuB2s242PXpy53+GQRawQVLaHDn62pGb1FI4Ik2ExcHPDmc/pUHb4vdsWmM
ptB8Yy8iy+Smesk0azX4W3aHrcip0lN2tQoRCHL8/PycIL9fMKTFGW3mQL9Q
1FbFfCUl4w86vDIgaqdfmzpcBBr053mMPCBXeHTZJO0KepY2xajilKsNtyKD
b9Gn7kGBviXfIIEql81bsd0m/WX0Iu8lnZZ0FIX51lB98FFmMhd/18gmTKiF
BkooxSdmbNoK3DKWA/oqpZUBBqVdhaqkRa9YlI8VNxeiXmgMPsCJyxw52tH0
BdukXlYOjxASdq83laRe0jEnx83AJO2Ma8GthlWvZtVVLzKgiMbITcc7L2j6
ZUVacjoNDId5Q04LDlWG2v5HdGiFdvGnydeU2D14H6L9HT8txmJr+ntPSn/U
+Sjh+hYULKOM1QtwRd+8tSmHziMkKYv54v5GB9ChkXK8fDBmMnpBYnlqUE90
77cwBiwQhYKPvHC+ra5+aY9YIX8KQ3Dzph+kWNrnf4lhiq6STK6rLKO4/haa
k2CEc/o6lC1CTVpP2MmEmPs0la8ldRPLVmb4cDMC9vePhg2ZPfMBgy5s+Exf
49WC8TOxnoxjWkK3JP5uVwsioecVIyvL1cmPPRwv8XIW9/XzUjpIf9MEPypA
Frnd5NqKsbZhzNrTMfQj19fbKMwOPUqe1xtNLIsJW1JBkA2TGf6HknZRT0rq
Y3MJHaS6Mmf+CxD8gxkrdBapffmHK6NTGL7kWsBYL7gaoeNTuJw/2n2lBlot
T+2gcpHBZoixDif5+iqJgK3svrUtq0PvDJM4ST8aTguHJmZxb2/VHfDcZBTW
GyR5Mz6CHHUo4MuesbtA4PYFWXUijk7shc7z6sbj7EXKNtPsItqS/0mIMTSc
DmDWHuGZBXh+aXFb8Uho1kLgwZJLYtKruQ9g6o2zXJ7XYXtsfFXSI76+ZCDS
Gw4SbsDZ+q4qfX8I91S7iEpdD9AY4kGM0yH59QR59PzhrCfTeL7prhJ8j4OR
PcsNLhGhJqgbyPxJB4cf0yB0nFnw0UBulHpmlxTtWFdqOs9RvPCMvwAyNkyF
9wv29w21vlyeb8dowMdB1Ps91lMYBc3/kiHm/JaB9Pck0rUQdAWMITx64hsr
rcfLsW8e6U9BWulp7ioGjmpzHfZx6sMVQDx9rmBfQaBnpK5NawfzQ/zWwln5
8aN/UFSjs5SlLlFl0NPdEHTGghf61V/hl2qxY+FErwAmatsPs2ID71U71C2G
oc/iD3izbpNEPfDVd2zP8OSPsO+gBNlaUZ8+EH7ZPWgkyIWo8eXEAblMfqs/
Qb0PvaWmcwf9PikcH3XBP6vIrWNq6zq7Y0k08zqTwdJB0qX0PWjYy9eGaGFM
VEGiRyeqGerMiWX1OtWF1KQu4WlDTDbv3xLGcoh0Cu13Bi8zztm2mJxIQR02
K1ROL7viGTk3cGHFO9tDkS1ko4V6hX6QlcfVvw/e2Q7Ca/hiuZp4wI0twZks
V3VplNLrXmvizrFbvGRzmAIUVjChGPe7RPR5DIHIPMbu+/yfH1ymbUKEY6nM
C3ceJxp7KgY5v4w5fZVhdoD0T+zJFUd4oV3QNFGFX1qfrolBF9z7AmBL/JT0
9pph1nhp1YB9ycrZ3XMzCP8cagCIWaQaKqlk+9XN0t1ClpZsme5MocanXdRM
WNL8z3ZIesWdBP7f7Ep2MOPfrdFnOYfhPspiYVTYzTYMD/YamE0aVJbWlMSQ
2MohU+28QujFgf3Lkw3qIlgndaXmztaAg3RzZUMt9cjIqvlssmu5Z2qYPQs4
05MqUjGWWUy73OzKG4ZDM8cC+MbsFOP2WgetiPnC1Un1hdYLb0IbyiAc3ygq
kbHjfvR63gPNfsUQMOwmguWMhC/a85Dz4H/mHBvc8Zpy+yre2iFxdstnMdFa
DNQGwp6INs1rA5Z/6HLSt9cv1zhaeJDbDtzSfQ8nAc9FmdcLcOIP2xudGU3w
UM2Wc68d9hC//LuFuEVMkQVeuFwEUFEqxcr1w6N9rGR9zE+XwbFKL2h5vor4
hK4f5kU2VBXKo1o13TOvlnM3z4KbUx7jvhix7lEZY7ihraaSZ4xqtNB4KN1V
gZuPvry0bhcJxX9uJEZlJMY52QRMnGm1XHlR6WQ6b2GF1mOFS7a3SoHj9Fws
0sQQfQ6E0UWZNhkw20cqU9+lDpgX96CRkXRZoJYeOMC4zkiozs7SAg5C37zx
w2g0lYa7v29hCICvRFyXXbOO6/bzQrxUo8IyNqh9/1CLI0vLCCPOQ/q0PP78
97mfGg3epBSbcLBgJ2pvMZxwQZbZ9Tu4oP6c3KzuOfkSKSXVk+U8lOdvhFcN
bfazYiNijU44bBV5fh+DOO5F/SkvJA0lTg478o4QWWe1i1uqoZlZ9zt4GLcd
lMDR5dDVGhTVLIWpYo/t22ZjEe4kCLoP9FzBH8yxrOzGMJv9zC73K10zuvf+
fupSW2SKrsGeuIpbE+3hy3+d7xEmMPv50oZk86IRV9TmbPGeqjgtkrgNlLu0
rAl3vMfj43Utc1fqvBrE1kNB4FNRrO5ZOSWVrfD/J0YFDhmhVMB7+4nRyzQm
+Xfm82ngddytgjY7SgiImxIpPARtm2hCB/rKN8wI7yYgglMGNIl4u0uYn9pV
F8/JBZE+JI8icL+3eJBdQnLs8ImJsTOXRbPv3gAHYcVFpFI9hworP1vZKQN6
HtUt+F7+hx1fuWRBA7SSP6Q3aPBatfsy74UOJPQsM1G9rDGWIHQl1ZRifbKv
mqLfy8S5z3KEwu297Jk5GiAPPr8Bl/TM4jiqxGZDNbFrVAvK2+hHZJR0km/1
BzeJ2illeTjp3+Qdto/0/7b2Kk7KHAkQHfCVQCa3YY5ymwv+lkHbxmxJzVwR
V1CVeZ2MvZYYTSCEdopMCI3gUDoyvcqKmFZXELVqMLnh+mfhMhczrAJoOjm0
KBhgnmXl4wbKXZUGAVPeIhbWdLHbvk9z73v3dblpLc27T1rl44KQJ6fUwbQz
ER6dOOygKztlhz9/XaloHLzqDO6iNdJSsrVnO04QI13M01Az8dfKUVQmVnCi
rUxIhb46EqC3RSGtS2NJ3FphSJQBi4yjZyBxDXAIlAO0uQ/ZyH2tmHFLRAir
NODF/Q/tmchiv65BGFo2orwv/kh4Qon96cmA7K76v6PrYtG5mDVZrtF3OVX9
2dj9Q/PixRyM7pdyscl2IsqUmidzyrL7GZ/m+BQYWXjuLVYSxWIJx9DFSBvh
6IXw6mE8I6zCr4+KY+mcrpl2hwUEFDR+Xx56skkVnl4KwHDMfg40hasEOmFR
06D0sBuh8CnspHxolm7TOW9pY98dZeOoM2pLgQDU7W7bIskSrq34ZsadghN3
gzzhBWlFN2C5TmTXS6E+Q6ajD4Un84NhBijP/saGWwgRuJahGSc0OHghPrvB
b0HTZSA3XASZ1pgL0GpUadL6H+O6ojt+wLSPvrgjOvjNdW7BEePF0woFoCQW
2ANmUFjGHaDrzwOzRUTqn6hHWVjtPBrsd79m95VqX914n/uxKeeQpw+VROWD
FsZ12G4k0UXLODMhZlpqPnDlG/IGJLOrsy05BMMEiuqT42k6SECdqDSrf2UH
UiWljkd68z8nLLOIyLUSHrVWV0B0mDAaz5r3uEQXTrIVuQ2DB7X61Su8JGM7
HGdWocr3PIJedrGV8tqVg77cOoKZL3LrZkOMgl2H7RkfJLbDkyoPAlQy+Ruo
+nGbNmx9NPRxnGWJTt6ZUouxIGdk5gRu2yp589Ov09HBtgSQyGPYn/LkZecZ
eKLWQNOKTLJz3kKk45lhPAz31P+1fMi/LSiLulsaswnn7ieQC8RhLH79AmCx
igIUaDVgYfMV1h+etKswRDFSG75M5WeOqMJ6L1ROybXIo96HX3QLdr78TArE
PVrtP+hg/dpvXsyozIjg1D8Zoun0hfaq3HQjie0c6lriYY0c10f6Vivgi0TI
eHfJjA2BIC/m6DxWWV41WPlZu9b5ag5ZubnfUTtx3/Q4Rr67Yy9/dcP6fDhU
3CsZHx0V+jui4qcCfBCs0iwm/SlynjfFVWZ+onWUdz5k1ZBkK24sMlLUCTQT
sJgjEiFZY2YNrIA634HWAZ0kyLVnIoIYPNdUopbF9IwilKhlqniWj1ZCDIo7
CCAAo6zlcmn/gCAHWtRZKmwblOVjh0HOvRWa7BhKKyHDScQXNpaJR3AjuBkn
P8m8JTHCovtzWqWwEOGMKU1SIlOeXu8Z2vToYW/aFkCd0rq4Lj61RVic6GW5
M5xiN+jl+dLP7aaIHs14tTOkngkIy1whnQNnMR3XCqCil8BIX0RrD3MYB/St
INgYvpP2gFRF1I1FKsQgIrcSEzySPUVbqluLspGI9LHDhLOpDyEiskEBDAXq
Gjpyd5JLdraKqTTxuZb7GkmcrKW4l+3z9egs8GQQzCCpcfWkA3ohGBsj4via
oWJ9yT9RnxgGNqUNRRvJVscSMipZBGoWzVEzaWkDIvVNgSIzz3q7EdgpBme3
12cRmZvdn7K5GG+E868QQMot/yjlWQ+eXO6gOWLzOm2eog8HSeU+mtDfskQ6
lSe+V1leIZsJimEldwoqh2wP6Q7AGohwot4has3Cn4aJOtRskD+aSo97PGUg
UFhTgfYsjnLyC9swcj4HUFv2r+TgNnYBKFM/JkBGcKiorvdRxqI79hS78DTu
MBkYIsoWXe3NAzQzdLu1lWyjXgoY2JHMLEhzG5LgBSXdtzw8FvBBldBN+mBy
dSnvbD2g5yegfwiP6IalquyNWmxYyEAYxSm9dztPUslbYhcttM2Wj47O18jn
58FKmMRF8tpzY77WdIkoQaHV/Hg5h8ah0PV4LxFDw2ulenbGNlg8tIVukadV
dk76cZ5fQkmMzQ+6KKvKTNc1DVNfAhGAm+ZoedTR4bFZOoFDgAQO2FlJbBzq
O9qrWp9ljQG/w9+uvV3x1lDRYSgSVW9mlUgMpL2v9kor7YeeL9DvwDEnZG7Q
xemIkSMD0fuezhItm+GlJHnWDF0cpHbqVdkJh52xZdRA+SpSs4QQOPX5GzoN
Fo7fuvMz0beU3IPwEG6EAcyc+gQgLWN0ulywShp1Qk+o3TSD9wBGzr5iHcXT
GSO0HAsaNjdatsF0q53a4LnworukqpTP+yLeDm9Q0rGxIW94GGl4VBPeovMp
HaueiOos46dZMVI+dDJYusKswNRQszn4IgeR87SCjCEPZ9cdzZuCf3rhODdf
Cwyg2dvs8yB/JWtcgL10dwgSv5HC7d6+8QGu8c+5y0ssykGAATwpGChFz86g
QEFRNGBESR9g4BEfkT14+pCQVay4FCn83rycdkX10+whKtzPII9bJkZjAm9W
xslSqK+vA9KnXc46y5V59MRu0XBhbdghW/XHwQUY/Nqn8D/y/zLdU3x/FRz4
MFTsuj289mAnyhYIe4Ocm4kIZPdGe4QQ6V7cdVXkjGyfE7bB5ZVg6HnJZVmz
pgAO7k3sf4nD0nBygFncXtgzShgoUy2AojgjnTFLa7UzjQjFOrMH+UeY4ji1
FIwT2z0tvemLHe/d8INM23IKpxFQi8ZrB++++FOHq5X4YhxNl+db5BFgx8H6
sofY3jbicPPZor11z5j07mg+9ldLiAAuNiCm0V2T4HNA0XlAN6L8yTdJChna
90dkOzQVjfNSrOYQFAsMTVG7UgU6de88BjENQjLFdtq2TqM2a3Jk5v62YLRD
vUsYuPlhZd1xPaIKMdiIZpb5imJEG9TrE9E2C6tZfNChE5G0HuF5XLnM6L2V
64AxK4JGtj2bgoTykhza6JbO6c2eczc0XwrknXGgmKxsTcmH+zFFj4igx/XR
oeBawOBvaF9TlzEPtNdMPlDNaxFtPlumwMywZ1zzUFR6cWKPLiMJjmIUOUH4
eZ84vln75iXa3IjyWs3vKDGnBmhv733GBKdVc7UWdJ9BsblntNBSLKDwNxRw
DeLAtwKxnVvVbuirAj0lSHdUgv50sjbQz7K+ZCh8em/hmKGHQ3W0fC8Me0vJ
yMQu6s2e4kLlA0MMexK6ySkqJBVkTe21EpuEIheNZRDMjcKGV/bJVgKEcHqO
pge4FNNT/gzIZLZuBbAhoXrRjYZDF5IUaEtxJlwZ+jDWa7EpD/31y5/zMyK2
RT04Q4/pf/7MU0rV6cA/JjlQ8d7eMJCpImV0FfqqeB5B78ylVs7ECbj8vfo6
Rqd9/BwafkhFZMGIKWme7OUt8MDaS+YwLe69MNEz02/or2Ne9xnYQVXUKlrp
5QqgWTZHBtTZaKRwLI+jDntLvwfSbDN4TrdceajEDVEcXOgXVGRM69ajQXvs
kTk0jOjtGCx21X8DLFw6RwiV3kl1yLRnov6HkMJHLyWWtL1EoKBFoJ532FRE
XFwLr0ITEe4lfKJQPcrqeCjYhkcvtAIy0Chy3eKh6fPS2bPpAYAzgybCjN01
Sot+LY/xbkvomjp5LfsBOfZRh/mFU3tQWTLvolCfURgn7+JjZPlpwRDLHWEp
K0T2fSaeUxf2D2yvUosqDxNFSH01/XpfJXE4i4iikSw30f5PlKJp8/7Mc4pH
/fxPZOxsrXND2Ur9M/Oc4cMsZEQT9nXT2MokntOU0Q71uEh2ufGrSGw+AiXI
6nIGEvAnQFUWrBf/vvGRgYUZZIZPI2qzlEcR5uFKcL7M0Id9i3a2YK78MGKs
plGqWuHaFK2m0DfIhtODuZAHbZx3x7K/mt34rNiuGAU9dgH2xp1Va9XJw6Vw
0YMZJF0vbyyLwWIRutMM73xcppfdwA1DkGZaJFv0guAftuKeE3G5YwbjXlxk
MgVPzcgIjbh6AX0CIBaExia1siMXIhyJvIIAErB8dBVhSNA1C/nDk7rhnoHz
bbKdfhoBuTCYqZZZRtIDlbvjck3uisyU9ZaSAXL5nKsAyIRrHaRCkko2s+n+
guW9EJEtXialc4/tgbCz0maUuaWRgCKb42iFk5mXLgRQSBk2+BaV5gqftKCp
iMlTKTyKg8ewQ9y7ZRCgApYjRiyUtuQHz6sFrfJU0VFgZhMllZsD6HmFOpdS
aaD6R5le/azM2OdCd6VnsD290K5G3KYNI8y8itVVARP0LW78xew+rH191M3q
Rzpa9WKduGMDnWmtyN6JqIHA+27i+KuZ2mw/Iafj0Eqfez1kOH4231gsNDB5
Q7cCN5+g+R7/a8+XcWEWt4wAG7DfkuzhkTSIurCINXAvp98fy6TjCb5V0ctz
lvHyBcqOqBxA3fTUtkjBc2KNN3XnAyR6yVy7KxyIApxXbtNF25dqs85g9JaH
n2sD2HnDgtXtXQV/e0ygj+oFu0y53VMTev5UX2qWwmRH1otlLELvqyW/W+Gm
Inb3xBANiYHhrMnqhyb2EnDztY9+M4cFkVIFDGxREAPFaKq8rnyh0h2e7zYr
1O5DKMAuNJGcsd+VgyvCbphgSuznFRmprAIgoO1s9J9+8oTULGCvvgQB4Tnu
r9IFyLnzRjoEG4yyzF4FkGYPF+aUOdhCi+7n1Ll+qFcU7cax1SBQVQl/AJ7x
C/wxRtzMZcadxKgMAD83i0RkltO/4lNwAsrJefuQyIrCiCV4y2wxVteNZ6+f
8gCaqmIHRs3+QEe34G7mcGMcMqIzaRzHGgHwv6Mv5Wb7b+SbXS/ystz2sR6w
mGs9DPp6A5GE0GhT78CfJatUsimQC6D+Xr2tcK1RP61MwmmOTk9miLAjqcm6
0HvO6R66KiwmIHX30NcM8IbqXslcrhwzI+pSaL5aKofuxeaEmyC69quv0o6o
ILClp/nazDPsJsFSyax2qZtNnUgU1Vt0SvkMQo0L9DeXYgAiKes/Gpign8gF
BydNKI1OQByKPUQ5yspeOZY6vjXEokiicMTsqJhMZMbxdBgYEkqFiY+PUX7q
VzeZMLuYWgR/2BeNY1dlleGhJLDbMdsWONC7Qxl/5FHfI2sc7iXY+emOb3oe
WQt+2uw9E9LZThfJzcv+YxzkfGQtujKNQR4wzdVF84yFEwxhZANBzVHKuO4+
vV1R0pxMWqJyUqXPq1N2OtLaPbywllyNYbBg+wzIISlyP9FiZ2H27aiHYPfB
bckttUZ+rrXArjjKySBxueo9fRFBFS+excTPD8mRRlLeqzO9MRjJ5b8n4kwk
4c6svxKOe1zhoQxxverfctLfdRfr7p6FJ43Fd/X6IFaPEo76WcgD1Vp//ot/
Ri+T3loWDlTvX17NDHxD75W+SzU73qPmc4EyWq5342s8+PBgyzmzDg9xsPs0
66qmg6s7glBrGiB/454DchY4wcw7IVR0X8TODmX63g6VEKGDkEVgWH7oQbDw
oubqm5QbxaAisY1uNcLvISHCMgOnxCvohOMduqJKD+6BVmQeUv6uYuriCIV1
mQ7nLusX/WIXgl0goRajs+f9WzZUMJx5gbRy4L8yfi8ZcjoyvZXdcc4oAYow
DdRkopS7U1vTkfxCe+jtQ5kZ/xPs/pHdEHmR71GLkREXSJSDHOUHjSFYw4xw
I1Dws/U6ViWf0UirB7MGJvxM2MhNKFn8GLiOqPF1eAFMxf++rHAhb4mLMIs/
wmKJDK8u3zMsKfFtfr+GMV1H+vpGjXGGJXZwo7OUggah+jNXkoz0nHwHsxlR
lUO1uezsmP3zBkgRLI+2FzTjHfHIZe9ahTWR4NVhYvA/n7PxsnyLRTFpif3M
EfolGJJDIfhprfg7deU9wn74WCNBDzXuI6UsBm2iMOsiO8am16Cb7AEMzw2i
m32GIKTQ8WumZ4tS8UVWpvhx4hk/3LCOGs+SZpnPdwDBqUKdTT2E3+jWX3pb
ns2gbUxfXWP+HN8+tP+sxWpkZfwnkjKh0Wma6dsvcwQ7TWC7ekcFNg8w66gE
0dvG0hoUJQffqigHm4xiGYLp9UYiiFpBcISq3wHLgsq3xZFpFvP+9l+zdXeP
oPHqbxf1yCIVJXMhCT3sp9qhCRiVJBiV+c792ZXWjAx5h4w6fvGdh2Llovdq
cgy1ndfRJvSKDNXmlF32uShg2BIKg+FoWcZ+9PXhiWpWsYc4RSAqYzMfjy06
y+xuB6jQNUGrVcRdpFGmjfO7UKr/oGeyq+OragGoPs5fMVCKX2fCPfJndE8Q
OKVgeEfsnYB8HhCgMmKac99ELyaIZ8LBw42HSNAJ5rEVD9vbwmtsryPFBFPM
un1aVselXdgNuUzNcphOtBNjvPxnarvavVRn2KeSMCSuBNj7LkENugnOy3Ck
OD0isDrg0EaPAAdKEgtJvr9N+udaz3YJ4s2yOlw4wRkk39QFB9COh/hi8B/r
Y1L/VlY00HirdUH5XGcCqAgYacalQ4Mp+ByEXoyEVazH+Y31bt2glSsDn1RR
E+852YeIgoOFTtDdTuq5LHbxaj3jiOcfwsw8k+U2RPGU4v+qTnzo7Sdc6JrV
iKBWagewBu6tPxxOXoe7yhKbVS0qgD8joRvR1PsH3AAa8eevv+J4hsoIF1NL
F2+iTEAq9LBGS3T3Lv3o8WUtk+NGjZthddUq9L3vxgbdT1frZxLlY1ZfKMnd
QlKt36o+/O1Z+tKr8s4XXEQTP6qdRli0RDu2yK153190lzk8wHh9OoUugLrc
/9C/vdy34/FYWnUGCC+5HaZ0PBQ197nf8/QPwMc97e9o5f5vfkrZi6GfbBTm
3czokdtUklCg2Q+i6D2eWG4b95YV2+Cfku7g5YFlQtUQ/ph0MX50ck8O89No
kLKA5X4iQaw15wVMIWcIgxkVHnA0GP60/StN5IzMJo4apKmTT+NvDXVxDbM9
ZeP+9OsctO4udlYNSgA1gFob2S2iRyS/L3dt2oa9OY0r40yfrisRCoreGpYU
iAQ4JTXJV7u4PPusC2K5beD/VGRFKR21Nqcw0tKxlOsR0gqgfSPsDc8S7o/I
VKLhvXHt/h5KWyW0xtBVBCOWzDEr94b1yjfBWr8X2h1NWsJUtKXnGXSCiZPr
8Og4M2yPRY+SRRZqsHWbJ21lK9T+Et1tebyKj42wWwiRVCRuOzkqdVWKKhcV
VGH59xgoDZK+sNI2WNpL0MjhJe60qP/TrzcvQ0k3BbVIhrOfJQ0OVcZ3S4ZP
jCiHR+9KIPvKH7KJK22r3YdJXzuR0eQgU8WEYvuDszvwZT9UvipVuyFOKikc
3O3chHtXepPk08fFaDQ44sjCPLQkIP51tB5uHi0rIh7PlGm+j2a9OY+ry1c7
OvAZjzCuTJ2JEPF8hLJuJlWzNuF/9HwZ9ORt0eLiT7e4LGuHRUwNyH3Q3fT8
jwn//wvNf68RpuAkxo6flr4wexFAGMvdX8mkcgvKIXl9u19m+52iPr/NAz4C
Eyj8TdM+A/goU988P7LWZj69EY0nkRrP+2/5NBsJQaraoIWS/b8jLpDf2O/R
fHYdL68OQZUOWpC/dEja1mdGrJQLpvdIVXsaTNqSyB1ST0PeVH52AoPb8ecC
wUJa4qGbcuFpKhIJ+ggxVMO89Rt5DXXruwaIorBc8CYNAxrNZB9nNWSxSr0B
EfEAEdXBfTaLh06E2lMj6HS7P+OL/qQ+N3uCeGAhRV0WcJt8J370Tr/VZ6sU
yLOssBzzG9V00ZWKszZ0b41BRTs5+arz1kMTEODG8GPbgqs7AAGb8z6q7P8f
iehtd7wpr6E1MkSsa1r9toRlVxFCcAr+ydRSS7anpyE4NoXW28r/WzOURcOc
FAt9LITEmcgygygyuLsu3xG5v/yd85G9WMr2O/bguXHSMWJZNMPsF2NYUEhZ
o0pgcZFyHyKr/ki8Mt+3xhqebksQ1CW7ztxFTo2O0c9Hdnk8eapF8EVpe0Aq
ktXq30GgiNuUIG1KpPjVEYpQpnzFoevMzIeb/Ms6lEWoyPQrRdA7DIJ/VRKN
e6sWQc5jMcCnjvo+F9gx0QW/IFRtvrtF+anR12bi9o8R9gqd3HZOF7u2GdzU
KasE5dftbw57e0nkinFofdAKMXO7WGsmMLKi092P509IM3PYjUzjKLwq1e4V
ZPsJmDYnPdkgNP9kfepmOWS3XW3u6ED69yEPct73qj2jGQH+PylSggVnY6EG
1Ic9KGmsr7tgMmhxBhuay3p4Mru4ixUBaJ8h80hNaRT0Cs+qfnVNRMFNqouP
TcvPqIpn8ziOXGAWefiUVHQfuI/YPPbmgJKE0XK1Sjob8pcPN9+fo27siKk1
flFu6/NnWL8j5zSY33JaSoo78exj81I+lNKDib4zzN47K0ky+umvUEsqOPMr
kOuCCm/IK65Sdr1qKr7w1hsbm7O7dSnoqvHEhNIY+lziTYj+nYnrt7IMPohM
NVmPN8PRzS9m/jd12rZM5cZnihqf5+cj7eps+2EeebIknjXXT7a2ZD84OV2u
LLnrXM+8ikdkvpgXEj+sncjEOE3YzUJwUjVH5Bkin53cA5+vmaQxTTrFl5Jl
byHkHHnbvkHF6jX1WzQ0Vrt0Q5dCHeWsTcmfK5l/xzbAVJgMUBk90rR2pL9Y
YcE7ZGoRdLlt3OYHaRaX8yxjlvtgmOIw5ClMyvRG+sd7Ul0jX3mJfI4Ng0OW
sCPi9Nzlep1uZcAb5jpPEMFk1zIq3yjb9dB7hpjPBcz+kDJuplxaNJLWjfA9
YjszcCNn11P4oJNGiLOcbECuJwapYsdx5kHXK9NXDeXThBB0/H0ls4DUte0g
iDpAfVSWt7IrJx0l8lC3vBAKG4hnenAMI9DILw46MEPpZsBofGt9Q/BcXxXO
rexcoWQLL6mrkvV4SjeRZUujxTiFxB0jZYIQVO61bg/x8Y4u4a9P3H/0f2NF
iX228eeILO9GSg9Jxu/Ja+2y0dP5L30YDlrbfcWRWi8qRbJZp4YbNb3cK2JE
wkb+6QAVg2zIya0D0dto8hZLMj4CxjsuOQwzK8XNIXX09iQQsPpUAidIvejH
2STQaolMM9cCE5WuGi2/Moxp76lPEbtKwBZ1GNGtKBGx/y4Hnb5GZzHWXSVq
7SMS2koy5g1BW2V+wSNrpaIJnXG++isjjqZWdO2XUyzuPeMA44cLWp53I2J+
1HA6DpOHd+0C+u6tWHKtKEUDteaevYBlJrJ+VPpOegUcZq6O/W0oDfJVdUqB
yNanFLQc+fylfAl3s5n74waAZ1VYL2RqlIpcvs6n1tdTP3bY/GpZNTcaiGuO
ZE3PEB+0XILLPFTd2VIWbXHu+0swAHUc96KcmWfN3nDPJECNsRxVpjJsGih2
PtANNpuV7vx1wspeNKDR98PjtCOf10+PbmCbMhBMJWcPnCUwZT0SOZCI3SSl
g0HxOgrFOn9WyVi8oKwfOn3dpO2veJ+TRn/2v474lNbshkIgKYLVR4YIgAue
PfXADMX4zN1VEEy2Tt5VetcyNOnkweTBI+zfTHPB0afNIqK+Zw3VvD5ZMOu6
I2LMb+pvr1dZnumadGoeMRnVIKcn9Q5LAzGe926nmjVPaOowNCDwquEsW5cY
ssecZSqM6bpz0TwZz0X1/dUQjHd7TkYWPrDJbzudOAM0goPoe3KLvN5njlZd
J2dlo/R0WOOr623vHOPKdHQXHOInU3l3UI89leLepcWMR9IjGDMSjizkangX
a5FFItd18ReEerY/8l+AF3DJpw+zqQcKcMENNbrXmg/oRlUzEPnyHYehXNVp
yRWIcismmZu1RnanMVmYibI2PNFAzFx6Ux7TTDMJv9f6NXU6igOqUHaQ4wvw
H0brV8eTQPbLlKnHANAB/4Wu0mZ8ifueInxp1JSO6mpVAF6EF3/IOd92lvrC
0Vy/9WbeJwXcax1phKOksJRDCKvONqyRkZumEKo7zPCQKOncj/xKeJFTSc7V
LeUKhCpr72JS5B+iI1yl72FGiwh1WvAQ5SISrbtmrTAqcBMvfwCOzb+H5AID
xhxgvkMHcEIbrDKJnfPKLUoMYaPuj0CVOqRnJtvTuIME6Czemqisf1CFKLGr
tm3xq0VmCzHOxC7sH3vYzh/YR3/b/7yNjN8h/3GNa5WpEcCDrAIIQkkED/F5
OJjl+NiGTNljaHWREGRS0NdvqU1hKslJ8PVd53ZEpVND/WfQJpI/LztEnqoz
ChTs/Xe56hn4q1v3qSxnl59myvT04zwVRTBCI4YgnqMjDXSgjCoRonc9bJ7G
OQKdUZpA+wTMoQQwi0IW8/dQZ58KyzzGL4rXDTm5I/7efKXDCA0bfQpbhhy0
EOu2/6CT2a0iGCkiCtDlE5ikzXLS6EqSR0yNn/n43GzsfEAG9CU+Judjcm0B
BX2CO/q4ODy9L5bBXHJWbryAvpUu4ALNbUhDvZ8yF3WdMMyXOIOdOoXNM4hz
uVq699autBb6tKi1uPLekbRrKm/OcQ8ZlzoOsaQe9X3BYSgy4jq+SQMG/9Hq
vWUkL5bF+JtfbVNCxs4bQtV9FUpR9SmD5xU2Bkye3WI4icFTJyHOn4ev0fPu
+Ya2rxa8YTa1YFE4vo+AzYgBMGXjYLXPs5Lyl88VSWL+2TMyjwP8wWGbgEqi
YHysW/suVEiYKcUuGo17OnKUdl0IDYSBPsVpgu3visvclymEq7HBHs1x2d7g
jpUKR0D2gGHWMHF/kPdomUHtvI6C5/0qIFu8u3FnXwrkQNoYP90d67vlGEq7
wb3ryvOG3e2Vmw2tov38Bua2UBMqBchFxrf7pKS7DVvFGXYH20PAoW9ORCDx
KtXIcM0E0Ue+yQzmAMLy8r6d/QJkGkwBvQ5rHdJmGqWexg1XKqdkYTeDyH9q
+LgByDg6OZSWe59TxED0PoEGX6yWmUOjRxLVZBmc3iG/xEHXkUkd2U1lkt4F
vt/HGOVCqnBQ//1hTPGJGVx4GBjo7xK9/rsi5qyF/G3QvFG7vJZ/9cjCjxcL
nVIxtmMWwhw8WLUsy/WqnjABK2dv1cNMVO4cRhb9DRWc+oGX8e7t2huacxrl
8TmMuxmLiQTBhvyy1pZvLVG7Yyev3BloPooeY2YqhcjagrJwYkp8NDPpH55j
Y3naawE9uxhrzYmbQsv/dV0OaDv+5ZkbLcl+/ei/twh3h4mXGaop3XTnztys
BazBHszWJQKCQ02Lc2Om6G1sm6ATFYyg04Lng7T7k+jTFYtp0G0G91xG4ja0
1PgH0spmLY3Bhg0YiBhzZQUJoBlTSpz1PjTcaH/sYkTg8d9AFiH1fTb8DGPL
TSvnq2OO3IiFDG+Twc7jn+m6VSEbz6xnuIgQyyCRct0Ed+jMvkW2EQtpAAKV
Zd3HYFjHeZTfrXAMikhKpy8M4EzdKkWFrQkyvJe6Tz3OQi/kX0pQltg3bxT6
UXXZkTkSD+8vd4XcI3SaEfJJe5QIcgDu4SPi1jAxH5gx264JulM8iOwmCZ/h
K5FEQcvZ0zy3MDPEbSrpq8mjImUWGLf+JGCs4vr0j8P8xQnfNPDhJaNeFP9h
haH08O/V2COzkUY/TUFCiSHCZXGLDs8j0l3nyCNDb3oZ/XvFt17YbxCHGwI+
tyENhOjOYYv02xdzFBe/NivOh9UpYmCoAoYcaLZhttILWt82kVK6Uyu5kXDo
cxElZf4bzVIDO16pubebYD9LGx5W2cd50rAVmO5Pdj4DnDzbZbJ/J0mRDiIE
KKhwV+l0dKGP4N9Dy/wPUPvXbtmNMbNEk9N2DGiOcqqtytD6hor8pMU/y59Y
K97UU1RzpaD4Pjouha/kbj2IpxOmTa+dPMFJ24EUFLlGRVPN9ZC0iMBuKxAH
bK+yTgEkBnvzoxO8l5ROR8VYtDUXrseEUEvvQ+jqHjQWdl6WvO5CkpDKRdia
BEeaJ12pk6hagmjXgupkflltfPq9n+G8sitDUmzrcwwIcoHN4yJIEiSOeqea
u52n5+Vs1iLf9nO/ELnjhVPXf4JMFhrX0aovcRIyMR+x1zMGEPLWEy00GZTE
xwKSJBVl7yjBr80GaUTco12Twccct1dWze5USMfVoFMwuRSfxS67gTyV7eGP
LuXIRsEHyX+kO/P5jqmnnsrzg6S/IC2Tn8qVFW/TbecYQksKPns0D0Ea13V6
q7AhMAP/VpEOa2HudN3cUGaZNF1itlSiRrXVgLv4GhKfJpjzUvS7RGkCxDqk
7bJeSlrKK3iXExQYK8hIk/LfioOxVZqhoGYPRCjxv7s8yoTTRF2qklyZ7PeP
TfIbU9nvnDGxV4taXtahdAQXGVMSbPvIgz2qKMlVRTHEsvgRqW0u6hYYc1ic
71sQO89HLeyVQfS9uOvP1koWIvALjRj+T5w0oWl4FeRlHbvqW/UJIiJvJT4x
DtXaU3lacd/6FbrwN3SJQ2PLHRRMx8MRqP3HQPV/bVEX8lwBNrtBbFCTz3Z/
Y7U/oUxdNKJA5MFYxzv5roUE0ICS2DFjSC4YUYumrWrcwKx0JBo5A/as2rwG
/yVjnOIjweZcYpqT3UXKkZmEw6mNvsSkEoMlncM2cyhThVmQCjx/dt3jJ83S
RBB0mej2MVnJ89R2YAkYe/JacuUQG7GMNW18FyHxkYRMHwXV5tRyl/KPJ/ty
ZovTBNsRSNKL86qvhOBV2vcYonfK6YrJN6YBPG9eX+QSqGxUm4tOQc+yiZfe
bAskoEASCH6+s8H7nxy4bhl0LJPfL8ebW+4VcSlS5thd/7vtroRobjulhSUl
7eBcDoxMbBH+XYcgNLQJWuJZ0QBGEjE1Vt5UMFPDaou3V9vdFLqpjS+flVks
ubE+lUn4ROeGrErVDj08HwwIA1QYxfVoahB/H/jK8XjXfxaGWlqSR6G5NDIg
vyWzQAMc9Kzz2IoOH3pi/y1/plcPerUw3Y0KhZD0NnjJYlLJfOk1F12RC4X0
tfUvzmsnCQzrEYcUkuhBm+NpA7KwCm5uPxFKxbZ0ky7+Iel/p90UHIaCZ7Um
coRcfo560/1ALQD5/DpL131N8OScOtS6U9C4gHEAMvUkOXikFM8lemeNgifC
Y7pT//3uOpEbQ0Xh9YEj4IVp2pJqPj6ZXNp6yhWZj45D9Tre6ANG1vcQg8IC
5tpdFyr8jhnz1mj2AEoacG0+iMe1OI7esMLsJd5scYVhST1M3YIGt4p3rn4d
ercUWIsVVyqQ5qcvsq9VGkWB1wvU1Cih1s2qH96bSUMwkyMPWz2TM7hikbjs
1lEJn7qzwnxooUG3I3X9LMazxVBtzfoPC31mjh3gDkH2Y2lVMV0Hwv8C0XoF
8Bzkt8hxiIpBa0stizJQBN0460yIpuxmPAfAzdQSTEUQDqy7+BZnUgSj0/rc
o4U1m/l+dfET1RHrj9y8Ns93DBG5HvVdFv0OT0TUCm5Ibafl+FHisD1oj2u/
IbnUgpkGOH7mLakARgjvu8ACMbdPYCLydA2zXpeDiLuLMWcHBGe9nhsy481E
ccuTfLnKVDq1MCapDbDIfnNc6vOibxtfiw0hdKUyiuqRdvy1B7W67e3T9vPM
muXIancapUYUB1l/T78G7I/bwVRktMLVDe61rKzvJbGXbvbb2l7c9HhR4imG
t8W5e4qMxtqAfLQYtfo7ihXOjdUGjf+ksA05ozfMLoKa5zJM6u551pdBtPx7
z2xkf6tU0M/ljTS3fdIfVH5laPT3hIy6fjVh6sXPnqYsnRshjPJ+Hua2u9xQ
ByCft/IOQlBKCLg9yYOXD+JGrjlISad1FNB8z65WMmgtpjF8I8l9FcZciUwg
VJG/BD3BcVv5++k5pj/PzZ/d3cnMjquAxDrTzJiwehVnT9lrQOKbykShMFO/
tXUOezfPBCny+qVeYjGBp6K1zj6NdAxJf5UiKwZ8JA4v5OgNRg9S/ouydNVV
lfeAJf5JzKREsZlCnUi5/Da5QqBtpMn5UiLE3GJ7KUPmpCO4tseHUKM5gFOV
WA472eIqxMkuId8doUR7BTgAdhG9h/inzsnJ83mFk5r7571JswKHvIuzj/Fd
CjRi6IhCQyuPjj1TfUTBnpAqwJBLRlCuvlSUMw7chkJjy+N+sO/PM0WKdnPE
nOu6awaQyaq0MxMP5PHVaUuulBldHUZa0P3myUYy74kyVqZNQZnzruln5YDN
HaeP7ArNbTKhqLuQ3he55/Uue4t+XKQwdNgzjbAn9R3WmZYxkm/rrbf803Tm
DrPuiDGu264SNJeoUg8YIy/z7YJfESVatglfwgCcLk3onC9YLLo7Wyci20xa
2Kfn65ZdTG3mw6wVGu5EijwhJCBaAm8Olv2hLhO0LgkxPLlW/QUedYVrSiaQ
VEMKyfes7rc3vJt7+qL8aAzSC8e14EdpqXkGsBLt1DNN34Blv8UHoy6OqQQc
2aRc4wiBNp9DedGKixPqeC0t6GxCrp2wRhIEdU+G2K5yr5ApCptmJ6Y5KJhf
04eMeyHtfxWrmKPxH7Ka+rLQTeGXO/r6QbutoUMziisCZ9dBrVDCtHZfPl3L
Uj5KKV8dbjGLr7hSMzMzRm+wuFDBB1F3w6TYixw2JADMjIVKeilY1xuYMe4B
k97lOmkojkkon8ZRT1kTObqiN6KAzuaVdYXVYzFepYt3zVBIxxl1fzwir99R
MU++URHdotTb4P3GhKl8CywQogBv0VbOIZV89UOJ0cswG7AjL4SbWvGjC0Ul
LBPfTizJJhDLwfeV6m20Qx4ZmqXBMb2YZ1NCTvSYCSaCD7rE8ExRRXcimQts
OMMLpcj0Sa+3APIIjnflUxnVajXSRo9LeQBvFFKi3VZNPsibsrVP0bDVTWkg
I7mITYbSC6OOd7W3GRZncANVIMyq2Z4+ouMyvPVrRaEK5hOtNY3WexLIuGxz
jCFKtlqR/eyzanLKHOBx8/h3mmwcnM6+enVYZlsu1Rd4pqV4gbEnBNFGOnWe
jwh52jcK1MG5LicAXUL+PC6N5WXpK13gmwONbFu1xAFKZQKtG+7xd9v86yqh
DeBKdYVBUtrROc75ksziQoGTN1qsnZanPbjQS7S95C23tZ3PaWcSRkv/X6sx
Ico+uizrHEaCRLxgu0TXgYKbtPJSHVZX3JEg1qE7Q6YrEkcprqJCVjAh0Vq9
bxuAie/6v6cnipENL/VQgOMLtBYcqb2Yg6CClO+nwJ1An7qTKZzwwwBBidue
MA6fN1hnh5Wd7+gOVghSab10HVy+qjJWlQknK8r03MtBdjZbW9kXcLQ0hJ/w
a+6g4unQFyzBEfZWfu8gCIzGZU+8sI2klt+nDVo7XH7Yqjbtz4IMjYI73LX8
m+X7UKylrJOi5U+sY8TPIGV4HozDyfaCYXJjWmsDoz72Sdo+FLT6R4IHd53F
ZdYbvcjPB164GXFlEHHhJi0/fG6RCUfrFSubpbIPSCgGqvuZGiJd6Pr+SI2/
yesovldOui/WP5awziynz5ZB4a2IPTTDzmuiKPA4dNKUv/h6CixzmFaF2ArD
no1S5T7aBvNXGYpYNSO0nO470U8XBZdGn/zhzdCrvm8ZBdOGM5F4m5JeyvUp
u/+UznZSdeY5+X3sauj26ApPY/MSWA1FvzDkgxqqjgiKWFjUqyUOjxmcOXbj
4oEK4dI8bq6qU5PXaPEmTy7bmm6T7bFoRJVJVnitXAemI2HfpBd+MxH2swSm
QqfTQ2NAhq0jQBFrAUEmFm8q0xkkg1zyPCCo5T4KzDvAZPxmsNeJwcOPNN3Z
IyGoH+C9xfRwsTlEdSQXsiri77wYtw9QBAIc+0tOHywYu+w/RxocYwG7+ZT1
iTiVV7M9k5dBWl1nUuAr26mUcJLVwHyCkNjU0E0Rcl1s18jJAz1/t1+xdZfG
7ECz98dGvJFprY1UPlNZZuyJVclLHfAqNJGnyPsxCb8rQywA7CGHMIs433ns
UdDMWUT+OpqmcXVuVR7z6oCMha/LfvF+rgaKg53I1n9Ek471KimMr+aCpJxR
tB8j+U9ZKxe2TNUeNJvRTDPlSXzi+PBkfZP0bgLrmGn4R3t0cQ6mSTmpH++G
WMVEMSPNr5PVabLd27EaHJJmMch7gyOVSgEkWWU52bw2lnQ1UOCGDPAhuI+d
jfABwI47UbTotkvMsQ0nlEFellHKj1pZEVD5wFYA803+ridoK4phGM5tw7GB
v5J5GK7rWyJ8CoZJcz1ZDMwPbYZX4RJ2Iv/qAyS/W6ToOKopzORJEuha0c4H
7XF+5q/VmENrFv/WBmMrgQhRc2TP7/3LdzvtcYFkO/Q5IpahpdexdS6tcXOI
AogmlyMNEpOTykU/TZ5gT+zJbTz3xLm53R+f6xGRh0CUNHOHyzNkHxaFfQDF
+XDRqrMDH0xe7ldq3YalcLNlTLMWkNITBkVjslUC87faCIRJBM1MSZYTg+yU
aLFiwLzcOMvJvk15PFi7AlmciyWQp8us3EhGAWw7+ECuMm/sFM1snAM0mmE/
olAM5wXe9LJiXj0hwSmkESdHp/MGZZ91uLSWzLkGapVtX5KtmQ+WuFDxT4JA
1xXkFn/T6LbePtk1PHPGrz0P0UWVH0sD9ORYlY5psESf7jGA+aTDBxIjISxy
j914bkRtKW5pYpCnjqljeSzd42xFQ6FvTTbQPv0wOpudh2lvrroUgKvlFbKV
HH+5e+1P2bwG5t5qzsOdBeb84td97XeyrYv8MmmY/w/mkFdZrqNrZcJ5LHsK
o+vdj14knTOPPtMODcwSsYjljLzsusIfpLcg0m1a/7EfPE1tQpPnlKQhK6l2
p9enX8hP2zrXb3rpEJeUWzsEuygksa56TdC8FwVXJXVXcBf4bih2hArShB0K
1bq8wZVcuklsiZ203C867YUBpqVQC6ZYsPDyi46uJ3CzTmxNidYKQGtTzNZ7
4zT1vHgafWEmQWJRoTWwsp3N3QiuMjSqpEyZL972DKP2zF3mCQg3Whtl46Nk
YEDrD6VVUPwdw+ihJhH2bdTRm129NBK7mGslCGoJt0QSmkzw/NGAFBJSKv/D
f0cEtgxV/bGd9OEm3SLZbC1tdFscFazRazo/P9hMVJZxb+k9fJmIdwXuhc2l
nP0aZPHmxEEseLpwspxcqcLeb6X9ugQA18AJa9GM+z7kRiJxsRan2nHU8Bfr
+MTUu1QHtJzQEAv3pArraIvbaFTFNlB8SizQjnez4Sd+SFn0+5KZtiOlx4LH
cJv1/s22US7/C+0EI5+Id9/rvcmi3FYQ3b4nEmOpWihHAN3PJD/Y4WP9UvVC
Dio7uJFCvMMqiv8jBF/+XIj375tpJnog+Fm3EpFTlBqDhkUhf02Ds7tE2L6A
xOD3oBMdP6/oAauyNqRIfroUcEhXurywY77WUP0v8ohbdZqlWknSAjjaPQIC
kgAS9c5R05rPa0kbe/RyRoDf9kMs8wEKaz42Kr3bY3w1Gm+37PjgwxIAF6rq
HefgAqfhHEChH5j1lJqmON5DM7ltYHPAWoFfVqCfO7X3SC53je8ZYztyP6q8
VWcu2Cs2oEjqeudst0wuiRC0Xq4DWLb6esF18kKJqR9RgJ9RuOnryWZkYxta
1Swvic50yLrgBJIYjMy2LJzW5y8C7ZTxuc+Z35252gkqvIb4+AzQYKeIAabk
91GSRxA8V5hKt48DC0+ehjWbwpFKo36wxNxbbtrWZfI74202OHG65BX0W/e8
i8RMXx4Z5tceGWVFWNRruGkqAt3DhA9YmJhIKPK8vQlJNwTRxGF3tAGHmeQ8
yaqYT1xN0bfprXdbMs85MUIX5rF9P4phhVrjqO+mYjTGen2Y3TLILxkWdBDn
uM0d5Gb7NfvQbp14WsNSwOtWT0wU1R4NXTg9hfDbqI1MP3ZuG1lkK5pZnD+b
n4GgmsKHWv7wNWdRzIsBoD7CuzStuu5+4sJOrnGFivqeveuk+6b/amZDG3Fi
DN3u36uY3qfLtP2Pa7WFqPm9N9x/OHB0QabQZb6NLNbQ8rWzcrBPvcHlgOoZ
FDCnG5zzmZawPu/x9No1hljmiS6pjjy0zdzsBB8NxCk3fyYN+aQ3pD61pT4F
YKQtCy7pEbxqC83L7iEivFxJV9kq2bsluIF/IsrN03qJQ387zqui4+3ja//a
ptfa9EiRImbMbauucbz/3MXvXIX8n6Tx4qaPW8cb+YYvfOd6qBzCmn2PDUD/
8XT9cVgnBIlzfpGxAPJZ2S1u9pfYl+uLRO7t+nnjeddRHUxj5cgnEbetP6ZM
vwhsT9lLuIfekGS1+MNHhjalKXjNPiryYew97RLKdPmKS0kkNemkezk1kK8X
TNIpp4MHqdqD0CSowdFdcrjFmEST+eo33l1Ce0wd0id5JHDyeIjC/85s5Cok
qCedoNe9EUs357GEtAn+u9JboMlrCin5HVMK8GyyBRUUA5XstIZ6EyF0d1M/
Rf8N1KTPmss7nhItxhFp+pFBqZYxYGl5eS/TEZfljv4waKmc/efwwP/1cUMv
rxGg/X8iYpNt1qNFnIgPlFPPV9CoTn2lS1z3pKrD7k9nDL1MJq3zmIqeNFJp
psgA6TVh+U/aZM3l/oFtpuQ/a/CqovQV8m/zOyoNfbUyIZvQVtxEkZ7DqXEr
cZbvG0IbQeO67HludgXaPQMjUhAGTgN35SgU5nrE5lpuz1fXeqxLOdOaKdSd
HgK7pF+GuZPPiieXDeK8omxUik+pQzmTksZihDxTzZP6UMsW0L4Ek204K2DG
EMEFZCy8zH4wBcr7rSGPneeqORay/D72qzYyr3DggCObXMILorxJ9oSm6kSS
XI5oXiN6AVh7+do+KZ8D2pJvF7I/36+P9tXmHhpC5J1t1AbLvDd/DkJNlFbx
w8pup9YXa5P9o/+QrkPccJ6hBfMHRs1LVrmsmqcDutjOcXJYF0r0odJmb7GB
TH0Q9JVXyltalxzze4s5VGpsSYgjuyHAM9tavPW0ot0zrCjrLa6B4W0z7D9u
GH516PeTLUlcxBcZUtwndwhEYN3zDYYjRxmh+GXZE5Cc4INqk9fFLjYoxWEA
i/MwWRYFsqTHAJjHdpIXjxZXUPHkK+XjeaqSZrfHlHPid9HQJpBtmBdA38NZ
vFxHSGPBG9eZOkyBHaLpd8nyZXFxp4wu6rQ/fIvY6WFTISLhbZRVmLPMk53E
e79BEjlJuFHwCujy4TkkNmnvT5wxC6uQqkIKFgAshk/YFtukQuTGSicQLQ6I
X1e3ER7QMk+ml1FwJxn+c2gb49Y2sJ2HywZUVqzIBd/fvJqbVgASNHnt5PBQ
2O0RAQhVga+lSJKT9p5YTMUVmbXde8ol+MOgTa6fZ2XPd62A4sA0ROTWRO1p
2KjbbNXMBYLvU1v/v+5Vfp0fh7CTcuUGCPdju7rVtvhuMC13ZwgD0llYLxga
LWwggAVVnV2jUdrHleif9GhbrnQ5kN8fe3ehCsc/G5dxNVut+1Rwz7qZkkz+
QXJlWfTcNbTn98NxGMsNPoJ82jR4HfNGxB2CqpLYUai3XUFZEaXBu5kn6z9c
ht2I5SRHA8wr+ypce7HiLZ9f5CUEYYDD0YR2F09XGDuhvWfTt370Ty0J83vl
OP361IXnuA9x1AUZ+A/yx4UUFSvqP5qVjE1BDUYHANhb4Gw7Gni2p0yjAhJ5
/00ijyJsixnLXcPkOwiL8AeaRKLIBBjtjZu2TGkBb7Sq0KKFFY5yM/S3KxlU
xhvyJ/G+A7t9UVID6v5mZtHy4PBwIIGOp20GM0ptegGa0OCQd0VoiX9ulpEG
aHXc6ywK8mkUJzjmlTvDpuT1X6yBEpqYjB9ceOyx6jVMu4qTp6QP0os2YK/m
Wu80DfwmvXzL9NCJD3pR8+FgrmBXHRyxxRAZvG59TCUvjffbRSshMap/bZaA
T6nrHYTESfH5uMaV6hyMrCwDjuWZ/2qUL3S7f9SswDoHrqmRLuzDX16IvSfA
ruBJAy3gbyUDaQjLttR6WOJzWT5cMDDIxXjmaAKsRier0FWFVLSQDCd8i8Z/
PCH4m+oqnzyEb7BUwO6/2skPV0Lbh1QjIIu1qVz2G7Tnt6wwvz6NYrat5nbh
bjQRyVtwS41R7eq0GB/kzDnilCCvwUEqWUIYzl5uqRTRrH2rw31/+SClAfXd
NO+fmHGv5Z/lbmVuL9Aweva+7rR5i9qS3dNjuoozuMafj8emf5mHk4usuj9l
a+Vq7yH5Lsi2hdpMMs/hfA+clIfstJK7v4Cf6qoxVywUfbZjBptouNeOb34E
65qqDEz8Scwfa92rPb/NhY6Hfrs2+VUqmZvlw7XMCSbNu2qjujHU1aen+fSs
Ai5677Se7fT3PqNrPmWpXCl9Q52PgG3g/0bliNFl/6HK8T0g6jjB8P4g3L+0
fKSZ6fm+qx0Tqajb7So7oXK9ur0euFB5ZVmcAPlbhmFznboH5fqE1OgLSggb
NSSPMvIix1KI5unjwFJJ1dTY7swu9atnDHvKB56GDX6uGMlwrnmQ1Gxen89l
H1/+DsJMPBOLo3gtQAEriDLRTAouBNx1BOUwJRN0pg+L+RiFpqw73ejjUyM0
8+Tr3aXiDVhtuDlb6FMtplzpYJ3XYnZWfOnXJ/cmpzxH+tkWfcguOHTtoAbW
wkZDC4vxs27IpHEBugR+z0IXv6kPwIY3zVJYP5zPdSiU+vzEvCCUrWZJukyZ
xBWkfalQwSs0dBZferd/tAXvcBsBjxeiA3FGyUvWbZU/M0pCWlO2QLj06Isz
asdrFRcTAY62TQ6kxtn7KNOmlJFIT2hVGJuBjaHifJjOp/PW9dIwQKsXu/RK
0vrJL1O7w1hfV9Qnwa8nKVPVnoInOhEz0VJo13fbyTKNloP3h0Tvps0KIwNu
1BPAcy/0sP03Q1g5uUOFH+tepDFbOlZ0yaVKGpTtyHQ2QNIEVB9UAQEFmxrY
1/bR2FXSq62m2J3MX9kpXn7eJoi0zkp3GQFJLxnP2l9NJqHIKSbSdKWXsohC
vZVYa4DHlCsCX/fqxFmv20+gQmBmNp9+ltDFEiznrN6khd1S9efTscSbxuAi
G1OhIMxF/NMVpYic7LtOpIMETwp+i6BUFJJTPz7eNvceoFYD6KpZfy9DKMtN
0eHxd+LxhtGPAItxpt3umg1Rxl2dj+Mkn4PZWTqGD/SqjHq+VAnv/6v5eObk
cX1LWL+0iOZbxveWQMxheoJdJbn+ZNXiSK82Ix/jpmd4EJ3xvUaUGcrZVSO4
ddh71+cKaWDTkYSiuJuq9m25rENRccYgMcgJoipbAbY76jZOGIMKZUq+L27W
AgrKQQaJ/yZuq63md3RRHt28b70N3A9YhR7Pxc1qRPqg9AuBq3Q00+jAA0Ve
uhoTEgexQXfcIZGbUsKHn6WUDo61wFQpGZ4pmRF5j8RAPf++IbKXpZ65cp/N
wDCFGoec4Hd2PPbtywoJ3wH1JRIKSLRr/Oene8hFW5heAzs0/Src/qgDdv94
wTpPPL0cJspkhMPQuzakGQV+PEYuys+EuoYi+sTZlrEyYrM2i2W+tWkBjr83
YskpzsZh6AI1SzkmQqsfwRfM7GGsqig5fCoqrXVlYHVw5GoYPL72XtMK9hjt
R5xqM2WovbXEl6RFT3sMtoBLz1vXVNqAATnvq3472fUCdgECoJYkYfB2dY+N
GSrF0ccJCG76bazrqfT4Kyt/WGp0+cbWGD4w9cifW5TNHHeQCSCu9mD5WkGG
1eXjXDohfwayCNqmnfvhKyrmq9yuhg6uePyC75NsCEBg8UFMfNiT2ngew4hK
difwUGyh5Miya2AZHHlYBtIo4rU24KclcBaPu3FZ3aLDqrQWNpFO+sF/R3g1
NPyCLKvZ1Y5MM3shpMttZUmChoqAcj2h8YsjfRCM3Nhct/5jjxvPA446KhLb
/s2/VuyeISHONyGe0JJ9a/Wz4ArvPvtUsvhFDdHWM7tCswNBQN1sspi8K23v
6XTTmm+sala0rFJsTgLqoIl3JfCXWEa0LsMY62ABxr3UfrqDSSjUBK42L0qA
mLgUD2RM8VF7BdA47oIqKGbgjRrg2BRxBOsEuZleP6l/95gR/K/V4gWjo+bu
lQFoGb+GJ65t1S0ZeFYgAODsOB+EhPevLALJ8uWzilnbOPf9iOta18s81+aZ
RqTOVANG28wWVkS4l5H2lr2XKZQsEuHMo5DKzBn7JAVOgD+tgifmn8InU6fh
NVOWNhuoW7KDSxwfE5MWaSDT5NIcOyza1oWRw6/NezV7TKetru9SiL0EtF+E
Bc7cQMAAOFJkue4klwYobR/v45qxiHHGLb9ZthKr9BtIkLvYBPAyIp9WrFCa
ZBe7QpOOIwyXIvSA7CXFM/VB6BpciHvOmPnYl8ToDDSeF7SA+JohpAlNNuv9
u7KK8HZPKnfw2n24wQHGpo5DkfqaYYZqoObWC4gdA2tA1lt/FL/ZUBcP73Uw
au1PhsjadHUswinvH8Ma4bCo5uoVSn8YP20SBrhUJNgAPjN1EKQbVCvW93o7
m8lXbM4rfLYOuY5YwOR4eYYOiJEMEnQnVdYLa2w0CHLn3P8+fD+bffHQLiiu
WKL3hx/zfOLcqm7WNnXyuIywf2Zxp08MEv0WPrV2pPUJqvxn6eXF5cmBHhDR
TwNQLkUwtJoeA3uLznj7XxxVKGyiOR0+gIZ+di341Pl9ZH2alpqj3DPe/KqC
bv03fwKtgeq+zeyPFi+2Vb1eQpVkXrlJsebXaztJDgql7T5ODVrbeWb1UJx5
kQ43r1m7KkOEfEa2d05yqPzbK9X3nHHkHsvL/StvFUlYe5b1VXR9hUButp8M
edEN00w+4tiqIaFDHcJypdioYSFP9OlOrMAy3VjenErJI+PlufzLCrEAGccj
npEngfH3D4ISrAklWsEa7LstvCg0PDshKvv5+taQwrIJolTZQM/fTLiNA7y1
CCGr4YlxNDV50bmXOpEY/9O30yGVuC9mCm9lb6dPa8nsOQZIOPNGfX0ikaa/
Q2tiWVfirraVtmu4HI/0KlSaQRURFgo9NfRFqrHodQWvD/Lty+DDUCewu9Sx
SWAHcSb8cUPfKwj3MpvjuP+DpJklm1atiqBMYPrEONVlI6lCrokQl9aqBcCz
oIZYH7nSlwlkNhkjXZZaRlDvI28sHo7CCoxvZmxxv0agTcqpZ4p6zE/tVx5d
fIuC/VRt3GhlDH6crikoh6xYn2LQddeP+NvWellL/GZhjA6rQTwBMz+UpYSa
0Xrvff/wHVDpqBc+jTU/gy9SI+i3jhG9Xe1hlvLx2GdphqRauYzLXF3/cetg
Yim/A2C3ubrs9wmK5HUz7aJe9Qb9K6G8w2TLgRoiXsNgAMaNeKi6vrFVmnBu
ZAqO5WJYY73vfpRGo2f5Ma0QD3BCIbN8bNm2MPlr/l60OjyxU1F88Zxcpn5C
D5iJd3roLbwJkH1E6RqeizTOC2ssjpyAVVT1YGtkypnlSxcqYLSCKmlrGOPP
HzmnTzKhPqrpnruOafdWrPhl3Fxl8PuJtkg8RVpKq8Q1FCnHE1bedecEqw+Q
tD9lnx03KkUEDpdcUjrSnhDic8iaL9zeJehXHcw1A4V2zsChs6hWfsNIbjTl
IQ4bfG6OT6/MZJuANdN1MXeUmb0gG427nDLFGBOaZtGZDEoZ43oJMKBJ2YZo
h6G85aqVqPSAAuf4lwRDKUgYTDebhL+1ktAjunPZbdRonDJboQKr11yRaEkn
oChrSufLPGpplIqJoU0jP2WdYU2/MJULb/J0x8e9rm5d8eh58GjcDQj9GZx8
JUxXn+PWlEJcDAM9cETGR3o0yKu2vfhcENaPdSx9u6O+YpJsb6DbGGfyK6FY
E8h5aVGc+AhjOCtwN0xluk6zEquphk9PNW18zRrzDteKYXxmTs8rEvL82zC+
XjH4snkaXCaRDTAAKRzAeyGRihdvrN5rcFyTjPh9LhU7T22Lu2HOeQsWbbE2
jkkme1f21mBF4nN63LcnZSqzUyzAbCOmXhtaRV2NRUwdS/tch1416vQ3ugXi
NmtH4099DkASkyvJMKDeZysqg6KGz77z01Wio93VM3M/EddIuI+jfr1IPIuE
aMZC9PbzprSn39apYoi3zOqUf+06C5NCDhuITFHbdNNoFDXKsI4fbbM+c+hW
ebjaCy+9NJuAbNoWCTkhGWMyFkKkHku2PTyZKazJ3QeN+CsPuV/42H9oPPb5
/2RewBixusPCBG39O/7/IyJE9cMLOAvYO5dfuBeHcbmpaWWfj8+YSA/kYM2i
O4Eeqoi8/ssuYmDCFLYlUaWVGWhCGNCM3duCJDA3UoZn+7asNGpMCsQAgGYe
nRgh2hbplbOq1t4XJlHNRItmHrarJ65reo1IIUUR2YnN9yQvGIOB+/7JCRMa
DPYNp6T9HYnV0RhK4ndcE9qqQfXKYVfnsuq3FYQZrnojhSmkabGaZPrK5U7a
W0fiKr9tGusCjpW2aCILBQ9TYRFZaDpRoaEVQyIJo4vUR+Ok8+4G0yOXv6AR
rx660Rtt5UBNyW27MX52ZrGDnp8L+TEhfZ15CslicANPe9kANDIRfJqnmCiy
q2ZWVU+l7jo+80hr5fWgdwJztkZN06YTB0CItdd9NLBIc9/A7QEGXXEx2reJ
BSGM1KR58Ng4uPyFuzvcZKT8CZKUg+2AkR8zWHhYquEgtdhie+6xcEdRJ150
D9tYBf6qeplL3nDvm/c/whjqf1B/QROFVsLuGMcu9L/+wmvxFKoDHyUmjrN0
/5616Lk5KRqwM8n57Juuw0HXYVZiXQ+XUYH93MMiQLaDs+O5huOesWKfcrfS
7TNPJlhNF7StZIYHbpNNq08fiMyWdC2LgeaGREk6kcPeY+n9DjjtJ63eFxsG
LOXMDf1SKPNhlTQhF+YHugGX9LuifCRjkJ07QuGJrTb/A2gSvtY6JtmESd0q
Wgm19PoZUZQHPS/7RoVrehyDkcOrqbEyVJnu4oYqLnwGSzibuLdAgFzf0mHE
quFDKHzHys/J01wGIU/8OVqlkt7+JTljvnYS1LxTEslRAxASHAlWfBLRaAA8
UzLzz8YtL7Iq0+/KrH7T1Lm/Pnsf+5XsyM/9l2EeEZXsrwFBfMPv2t7t3SG8
demtsZWjKbydaeLT7Hw/Fk2wpyET3iQcjNgNdRUI8zL7AvP1/8+8gDqO++sM
Vh7rakKI84Q16DWNfkFBAkwsiMW/Ruf7nuQLqIB+mlxf7Id23FWrV4AAoMlm
TmtTde/69i/mlL2dcl1taNpicBsLtJTlBCWrS6SruoihZHn9zv53Ul67jGBi
cH2gLGjCtGFA7lcxc8MFpKseYJjq1gziLfLbYE4QuLYkDkMQeEjGpmHK5xcj
zpiOLao4EUwvlJD0MlWE7HFf3ZjHtUJvqqEmev6bECXj7b08x945cjJs2E6R
oylnGMaI8amzPuusMTPYup41wyUdpnErGBhDgS4xFu7VkMG39y0thtGUbiT1
7bOM7NMf2L7IaISEE+aQyncIwze2jahoY5V5Phxu4+17Qj858rGPtUpAHVPb
l4tlZ6S7JnTIw7GWH1gFcwr/f2ZtXwoqlquLydAgDJT1/z8B3WUdsLvQT3+O
+HRx4Amd1bnkbfEvFNPDFHY7is4KkUoaQ4BPsTnq1wlMxhSyN0XwvYOBwtKs
AUhAneM8Ge/3SpOYfl2l7khz/pVHyU4m56lLdLVAavu0RNo6xOd3fe0d6jqD
7809g87Is+ZDSPdQpmW1YX3nCPi0yuS/hRBw5VK1KkgdNE1Y4YoBfrKzb643
/OjpgsqA+GSSzyp+cmamLeKdxUkqbusPwadLbTeQziCDRKoFRWzpW9NiVexV
drisC6mknG+nBlOhh7HfSLdsejz4nRSPmM39hFqKyB1wRZgRb4GIwVeI9xup
BUZLcnPHlcnjormy1nyxuHeh0Y4+TvL/8GO5cGNceaOZ+wiZKoEaBl2Nx5Y/
PcymuxX4Q3JxPDLwZdpDaeYGMtlFMRr0XfwNxcLmEBSvxuhaBDyc2Fw9nKd9
0N5hGhh5aemIpzXRh9ZgQo8x+GiypVwnmCOt2vcPFuEwCXmyj/yxKxKBWknD
IEW/nZn+Gukc8K6msW5YaUTOO2jJxMyHqvxjiJ/CTBc4LDbxCp4Z8+BELxvF
t97gqJdrEDBzHQCqmpTadlxTjZ8GGkH/tl/ZanzTVlZMC6L3FKbhMFEwTGw/
ZSA56+K8tEx9wDQxG8XVo7jh0yyclDpBSg+3DIGG6r1p1q/qAENyXSz+NBYG
8yazoU8SX7cNoiyye+4NqG9+hzgDrqF8/mzDhboDpIgiQrdCuGVyGoDWJKzX
Fy2t30WDuYtvpeCOiYs8QE1pX+YOhKlglVQ4tM5bk6v+d6s0LgAeY6YP2lbq
Lng0iTMyNyNa34O8WP9Bhm4pHQAEjCLC0oaxZVLFPbaIuJcqqsVKg+5ucqXv
+pePbwDG8OtljT+pYOeSx8fgxA1bwpR7jWdjSZgGBYECXsnkeT8WTJyFPdMu
0e2OtLkuPtHsaNbU1M/lXyi/wBxPirpf/QqSNgQrzrdwYd0lycC7JOofMepE
U72pxyJiXT0hLGMBFdbWVSyelPUtZSrCEfLsyxATp8QfPo1DvCA37s9wi0DH
48SUFTZH1yctfcE3RXnrITHvKW9hakN+3/Gi3upzZXv+HqxmBYawtJcFG8lK
Vwp9GjcSTIGD/+ZzdgcAE017k/pzoNpDYVFZZ2n53qKZ7DfGIPEZwhruVxNN
Hw/FW2kDQZgpeQNWhyZ//5m6/KcFk7fdslKpRwmRcfz6XM8bN39QefWuMnFI
CtYsnWYa64UVQBZNfrueXtDiUMo439e/n0ZkCHmKtSC4kTwgh6NKPlWX+T8d
DsTXKZ1URLTf0/q5WOWP7P9IvOYBQEBajtvMhE/198iVYQ0O76NjMBkJ1Q7l
J9AmG8ZfaD1qmD6EcqKRmZFs9TXxHP05iRluBmxUbknNgVbyLAqoc6gNHwdg
ubcWWRODPm5uwDbdHH+iWEL1xS8mbBc1p080cr2y+Vu11dZ4sWnjkfeFUcYy
9XH9Ehz1H1D3+tWiLlMBZvjaUOplLF03zXG54//JJ6NGVYPo5jgWnrY67ZDm
2meqEzqfwqY0p8qpN7Q3fRGRhDL/QYjWschfA7HgHo3T139uL8sBzR3BDjag
f4qCb9lB2lAlj5BLG+KQoFuZVYxKKAy1HmSZnNsmVs337dHiZN49K0f19q3p
neOhk/IxIyyimqZqzZtcTt9Ok9YVgqJijcocFw1sBYvWMUxf0z9l9lptQZ6+
BaRMF3VdcU0LsJ2rxMRKmZ4xdprBkt3+6IneAHrpXTmnrCm8n+A+FvLf5xRz
OFvINKnGtoixpyQJRqbQdRXXUDPbLLRvDhWQxnE6Ugs9wLqT9mNTPylIk1I/
Ox0NP/yyGkAIvq2uxR2uARyLtbf2iEsjJ/pbKHAWCkg3jd/9fzcr6On5yzmm
G+yaqjNeXivbfjA2LHE2n1Ur5ZR9sLcT+CNb9zWvcvZH02BOrzRXFTELD8hJ
3I6Y6XDG299Y3gE6fkaQ/aX5u5ZEQuHR8g/iIYYQ9hUHv1foIIWQOmiwg79p
onlRk+yCE40SoqfL4S/roiWPhAKahY4CVpV8wAa6WkpbYXi9vUkdoovq4c55
9Sm61zJhdUvKriW9LfuuiTORyFKRUsbydmBQoJ0lZG/xFqz3gGBsXvuKeAI3
IIpss7C9rrWQ8Wi6ml9kZHvS/14nPN+LD01TbI5vboR7OnSmij7FYm6LFggv
gB1OnzKWdbai4weyNYnraa9ZwMt97lLOmkVlO1avT9Y4S8Ho0tjheo8KkqVH
0c+gl4Kpb3Va3cV5vLhcjOtO5whE2IRKBD5VvRICU52EWk/AGcRXwJQB/2W1
ipxUiMFrutcbDZka91NNJhSM6mmXZLjgqJoluYOkIIlzl9yrfjnnS/Kb8xze
ejxE+mhaW7RwA5ygJdW9x6scR+xBLzGRGfJdWT6IEzChpn+qyShSfKPokGgb
E221STCy2nWo5FqFIkD0Q5QC+LKfP89fiw7Ft/aAUcmMZLDxGv6CjpHeMark
Gi9SLTOk+yPiCJ/JXCYWhndF4GNMvmAeej/vXsFmqTBOW9QWqwaEJGhozNtI
MENfwbBhqGLdZcB9+sYu3y6MxtJcBMmXpGErqvYJUGgF1FdO4uhCmQoo5VQN
XughbFFE8MRvygp4BwPOl5r/M7nI0FGSZSVcW7EQ0PKVyp+WiEqiEf+Or2ha
MLB7evo/urM+ugnBYiRFof6UavR2Bbb/R7T4iBYWfhNVoZBuM89+ptwewdCx
HFCtn7/fxUO8DcO9z/Np86ESizgeX1sEkB7S1zzV39oqcDylSoZGm1lEeSnT
MRQuaDAEnGhkGkhV+zHcSJzm5tE38hla+eshNj3s/zfB2H9Gy6QtUY9gSzG1
e2Na9L6U7uK0hBobKqT8eaaiAjjgXLN33ra57DfYjKVHnza7510nb4xdcGAW
00RSGcnHLwEPiEQuv4+T7L9k9l5W9Wp2lTtNki8iG0zF+O/B1FctZtwR08f6
JaIGYhztgX+xznhf8eDu8AJOffYFxgKPl8uFkA0cwIVEex30BXx1GzmzaKS4
R0ldtBZuBihDjsOCALXZ6p7CfKqWrDPLzq069ORundRngjIEItE6V5REC4hn
Dg5D9kG4gtlIn1qF5KYBZDszKYrT0MjnfWHKQcvHjIzNxoI/wEhbvqGoYhgR
mB+yleXxwOMDqyEEXErtu4DcHwou8DitmBAjKq7xE/ab6lstY8UU/eLljhmL
OjinCDl/m/1k4A5o3zBaToGORaE2kPgrcxIxyEmo4OWAOF1e4VQqwOVgTQaN
KBkxUgKAAJMmYQngkmJFMstn6QkkXpM9pFBfCE28HYXUmyEEwflnxAkqY/3y
6IwXvY9F3vmIBuA1GgHaHSQmvv3VTkBDkvlkSEe7m3b5UBtqVzfa6xmjW9OR
0iLNl5AOEBJ7n4WVaQpgA9hDg81PK+YGPQCFBRnWOpyA4jKyQzlaxlTxcwxp
rZ0HP9aC8Wi8AGv28Pc07+wfe1UYnbMMKcjrVSOdzv615koCK437Na+nj1yg
rAtKW8XhGt+xjgYJyojl1ThjPANER2MPyj0dqFjOZXFJemcG1zgVaWPxSJMh
A4MFyHVZebIBWrLFcMHtSOgxCgfJRO/DJEjZqIx7sDuQ9WZXbamdzAEkSAIA
4kf9cNVZA/a7T/Y26BLr0zHLMAkEuyTITUQJCJUVEF817Ii79ANcuJH07IBI
VbSFUhfzW60wTObw2WTFMRSgjsyj2hvKi/SPy6YhKnW3u9sp/hgFinugQ+95
YWPJ/8MZxgnWEi/pGxe92AxJ+A+jB60J8RdzUfHUvPUd/0XbThCL26nilmB8
Ix2kj707vYNa1/9djP0Bsji+zCbcioPhLHwvizPANmI1SKuHAJUnAM0i9ysK
JMNoqbRTIMqoDtCH9yPzLNo04MHMnpPbxLrBmmKowiR1EfrA7Ai2Gxp0+yzA
hsS9ly8Uduxk4llzu4e6Bxxhe2EzSzXKKPgCNagSZQCaMVM8Fqq+SOF2MnKl
5o5HkduwaRzrwnTm0D2df1LbdB6+2OsJPT968ctuVhUL3ui2SmHZzsKU4YwD
LdSyL/Jvmvg1i5KGZBWan3WKfcSxd5O69cVdpTJ/OA/vsccg5vabZG8J6C5b
B+S+ocQlOjdqIrSzTTdBf64ADqw03z03SMbmb7Gav2b0L5f9PpgCS5/JN41V
Um9Q0tKcLJoANLtuojlrWsByaaiq++bSQxvob6r4x30fysJXuAyg/HF15cve
zgsIAyux0rig5nup5TRqwAShhBgFkObBdROdGejZPnLG8Zz7XOR04+VLgeFb
34fWIL/QI/JGZ9PXcNL7qwvFbpfeGYe4B2w2s5EzW7iwTn44JCrrpc73jLop
JcJqUMMMG90T6NtJIubzywpDgnFWQcvybkGzRj7oHM8WIzczhFoU30nV0yHa
uH3fZjLzLGNituylbg47ajU8VwAU6BNhIXbsMEdGFPBuyGUadJANp1wDocvz
7odhc3K1sQW4pfGPV7AzwuVOrPDvKNvMXWOoHPl64gFRLsmNXlCtFXXjvgZV
etlVPxT3/civ1nyKpi9uLRQTUZUzGFQ1DVjpmjbCtWXF7QT5fhJODAsWlMMh
vJDuny/sGZ3APr3ndVZ7oH8+imApcmd1Li5IBWNIGzBM08Zi4mv9G9SURFOF
0bUcbw4hSSv/QUsC5X7EcvdE4ML0YLnvi5MIPVJ5ya+AanhWpOkm6CcNWmUF
kpMRbPmsOV/sIK76feCEtww0aNf8sPA9vPaaygjQwga+FVbPgeyIwKzZS29e
wnY6vanhnFJQsE924HosuU6XJGtKJ0ne2vdUHiqM90W+XowMKFjJLqqi/Z5r
V9Ub+H/CBckCVOrn/BY7GbzyKBZW2OTKHIafuN5p+1QfvddbXkBbSuNy63Nq
uZ0jlWT7hDfXVeEPFg0K6sXZbUACrmcZXIG917CkBaOXFQ1TMFENPhCMmPKs
sfSQHE04GekxC4L9t4ahRB98Tjx51l2d7rk2y0wLxDXtZc/FhKtJFqj1vcto
yGim42ZZ6JdBoshoLrMIbk7w4PWNLDY3u33KZqFtjRGojr/oNJ7BmqsVFXqB
CDnoB9MTTEGTqPrxfTvY+iX+lLFk5+UPGwBEg4Oxvgr1gBo7J5X4xjdjQ6PY
h0B6ihnDTVa0T/aVy7UgI97SgbkhlvPuVvCJWHmd/Lp2bKcqK9AC7dCK4fQU
vLc7kdWxCpXdB3dFp15q+8o+p8ZtkF+nFDt57kIhJXtYY8CN3GlIi4aRv3VP
Lg4pzxpLFE11t7DaaN4rTFpYJahlHdVUyXgazTy7TKxghvjciwgumugB0m+V
wbjntR2x7SUfKJJsRbxCqVTezE1gwwbsIVUEzHxYFAyFTYPrU8CLGBl+iLMg
TCKlYurkwssCkMVteNxZAxn56JDTxqXzPo1tLaYgJOEYKJncDrjX2l59152m
HIVLBcm0rTCoixaAJYvaYgZJxyiNhR+NOtGmu94eQ8QFxXG5teTp9zt2vxRQ
frDq68FlFT1VGsdXFANMeomoKAIgA1Pe5yp7YxZTDTDMZzw1DwKQdYAEV/Nx
hHAY6AEVAsrRjaelS9tVD9TeGL0pnN8XQbRH3RTK8fJhyJ5aYSzFBLR2Qc+W
HlkcZ7EIAQShd7tZ+gIixvKxVjd2Iqqk0IioEtFhuSUCMb/grhaMiCvRgzGz
ApvOid9i+YjFcxQm+mfaQrs/o2WGH6/w2ea+nIYwjPC44LyA4eCj/J0gQEu7
asXJSfieOMztfEgtUnvf8o4TEphqVub+06nhbrZjS1er3EoIrhiwSMUrzZV0
GH/B6EMRfoolTWopt65tyu62Ioc+e3QjPIWxX/u46BO+q5oMN2gc06UGGEvY
B/W6JKumSbJb6ea8HrVyxR2ZcE1M7NCe9iSbonTYq8Ma/j1YxB1Ulat4VWCV
sAy9bTa52R6qHDYgWZ68ryHmNspaI6T0xWGF+M07F+95jrn57LP0xJx14E8j
Rh8AEZ+meKnLuLMI4RLF15EpZI+aNbpNYu9R7eE1aIeCGjBXt1MSLRMOLEDf
Sw9y9uOP4DEiW4okAYUMkJN+CorWbBNdoDJ67RWR6BXbIS0yQhlZwEvdKe4N
wu0pcZddjTbFRuHXJ/Ms7/b4rP5ezTC6QZw/mqfvGlPGJKi3etFy5lEi5WUY
JLoMIYmy6nzMj1iKdr52E70D6LfPpAXEMd/3AfVHqSuvjXGdkNe/CIyzcB6a
r0YCHe/nrbMLzJgQgCli6h/9ajQhS5Yg8jRMhhbt7RYswonyHypRJk/VHlou
Eq6P8ZVWoAdPkGA6I5oU4YrTGmv1F5m/dxvwwzWcHCniDhwwHJrKHh8pe8OU
6NIOFWF/Sy+9c3poZxUTAmIcbIiZrRzNsTq6omv6q9C58KVobheWJcCzKbrV
WpLepawIHndVRB4ftkez8zWLUI43IXnCEL16z0Y53qlCGW2QEanrp2p8SU+0
ndy2f8Ej1R+UtuNiJJycjCB3CU18VpKkb/wmjQGaA+LR8wcL7wAKR9NVT7+O
g0K7f1y/E7jaVZbKstB8ur+04R1yB8vfSw1iAMTqdol979XkL5PPHpxonD/R
bkEl/TaQlkXLQopyWWXK9hz39XR6vfKKAdM8ST2uR/MabcD8yUUBFX3jQwf7
nO4EN/6tv9sV3jnjh8fojwXpjCYMLxiInvWVT2cWteg8OG4RwGdJj7d4gXtm
jMCi+uLFbO9lklpMcoFl0Y4lCQ23LoF7ZdNIBjGqs4ESL56rmxHYUSCK3WF0
MCQoHZezQIBMCuxXCGt68Tul4S5+GGFcPz0A0OSYkdwu5AwnzcZHhfXApDXH
TNJo7q/yXdzU3Ha3L1QTjP4o+w9bQ+IjQLi1s9jucEzoriyTmL8RIg1oyv2L
nV1jZBVt7CAqxiKwOnYa+LfPC+cZOIoj6dnA42/T64y0bLdAulATqdbtt6YY
fpueYxN7/S14ZJuIsxlx+Z1ROuDvDYUqmGcBwjbwD2i3dT/mOMqcUtK9u9Ge
dfK8vi7RV/VwAn+duAFm/APoRXklRkJORD5E+ck+DGnTAsEixwLE7GEgkC+D
1loTvgFyfbSA7vlW3eB5AAONNs37F9Lkpk2YY7uxlqhC/JGwGYYbeEc4xks4
VwaT7ON7Uw/enK+wuVHthahU5J2+J8EdS5FloB3F3mybNowibRJvfQhgK9tR
CiAlutBFu9hJk4X7MWPFFARFvCtkX+9jsRaaHhgGC/OjadSBGnOOJLPrEO5w
UQyRLcdyd7ZaS5SfK6z85oQyAIuIeZG9WEu4hrpn7oK+jkPvHGYiNDxUtZVn
uSf28I8ccmzdE8iiKkUhx2Y6z0A671GrViWHOlIJA5Bb2Qt+BmGsaFxNZ76/
JNMn1Ju+zf/A1+sE/KQj9Nnc04Hjjh5IiH9YcszKJNG7Qwt5dn0AsZHjcqtc
jSqMMpuLMAfMsFV2DoiiC2OzLBS+aBW3KkQG+gpyFa8WzrI0mVq8i3cObawt
hu8fo+6jg7a4VNepJnz+csBEusvSm7lLAns/+nd35s1k0+bWv8Hjz9SmdjX+
6m4hUpgafi0cWKIxdmMRbhy0Cwxl7v0DfVkJBt1I8WvR9aF404IS93afE18G
QchNaLER4irCB81ucAOvjCWhRwMt8411rOnLZAhfhWwtyMXlgGQX4zH9J/Mi
ahuMJ0W+u8IQ8vg+75cIs4GXQRAZw3hpewgKBvJbOeyXHA2qhtWjgqpDVOAy
y1GAUWHuQ41rkKa8f78no/ZB66kY/ypfxlo9K5eTNUHT0VatlZkSyvDk36F/
GWAUjrvM9cpHNyMpLrJWfbeJHOFiophQPSWoBQEQaNdw1ZKqZznqrDdujRqU
qOOEWJDSIsIiq6s3p+dPdRzDV05WIhEXwEpR7KGhk1ehB/wo0PSwlJSBM9pE
RBnTcOw65s+pzC6JGoaAkUpKbKfqDOoucn9viDlIPBnkq4VJEWi2gh9+lCoZ
yNuTiBTE38YkoX7hGgbf30hrxbPBbv7LqoZ9296uqiNwwee/uSRuaiCR839h
CbkPQ+bJkaFuL+fzAzEodhkNVPN+RHOHmQjl+Rh0gtU39snFXc0HHHnMI4jW
JL0g7B1bSXfahgjt3lqJV6bktBFluKZUaFU1dRIqmW8ru9me6h7ZZWlW27sS
kD/X8aIG0A8ktZV4y3ZjO0A8OfGYW1rTm3Hsf8/AozwzyL2n7E3CVKFMULuP
ImQjr1fXfmlIu/3cGI/bhLyHamhiC7kVh0j9B3HkntFYOlVfAcK7gt2UlNyr
YDpi6Zq9ebX0PC/3ECAEnJflWv25gb54eBSHZUeQo6fwt76O1jZ5Ll48nbHR
kOleTXjp/N0yKfoZ1LBkIx+X6aYgD9W9q/UxmUecS/pb+n2DrHqs3fE90QUy
SjdQ/GDefzLglLspQJHFUcm2Y7aHPRDIPqAGcThP1v0P6KS4FdxUxAFwsO51
IU50ckjG9GGIxv1uRma8mNlQYlpiFoKcqhb0v4kkMsZ0JLBr2UJnom1hPnxc
5RRZ9SCp6XvJOyrC3DOUKW14weGJjgVdCcrhAxk4VzcK83ZukjeFB49V7aG3
FY+BMLxwdZkXPoOhPdAvADgCJMcYEQm70iJG6GtHBqaTCTCw9Vn+M5bmLjeJ
0yikMsPw/pLk188vh66ejlW75tO8mTet0JPNqhO3O9VBaSHkXcOsWEJibeC7
xWnRGlPQahduVl2IRyaEqlLnxrfcCTnA6m2Pu2mJJEUlcohH0nMlA/tZfPGQ
OWI2+Eh7+8DT+LKlOD6xovBAgC/Fwa5/4YJTJrq2jns/+F4X9/gKq5Kv++NL
sOaq1bAUokkSBzzrl6aqyzAEFjtN1DZTcjP+PLMMcvO4dR8SEIfKOWIqMDZ1
nTeB2swrNtrI+SyP4C76jHFTCLD2vrZRoumJmWTNyIKbHNTQAl8coIcHCmNU
bw35LPl4C5vNYEQq+XfeLyKOR15DR9GxlabXu63HX8IeGHiQ+hHqyHZpMb0e
BMWlUdZNJy39vd7cnZLmA/J/5Ej8oifP74K6uigkKtre75kfUhBflu/HLvp3
R878h9W1oInQt7IzWBgdFD7BhHKZsEfDo9baaz2WZT+wOrAv6W7ZyISEep3x
aHzrJ3eZuH9x02CbPZgG8Ya4efq9wvNhs8tbrqsOqwb1NIWaeeLK1v9nTY/x
VVmL4+xAXdF961vVaDSKXhmaygGLZo8bqIEp19wB/WSI4unXV1pVTvFsVKsN
TfQbmwsMFy4KgKObqIogQM2eJq6Ysjxe6R3kEnmaw9NbfP7XolryIwvPNTpl
H+BXYWxHSlDnDRkzZjI74mk4gCrgBc8OBi7IRgnCgj8ScIYCnvIWevlQ5ONA
RNHPpIZFCySKHj4AIu353Fi5za/M1fdffTnTTB91uO1SyAbNU9En0c3rMcqr
xd5HG4KHQ6O/DdVtpQ2PUcUwdV4lussKxIe5+kd94edIgWSl8EmafScyWUaW
c+nG+RT1Qwg48GYDZwcSFMLLmoxDcXZsMRnulRUr+dn1Wpsdo3PmvvTDGgD3
Xqcqh+qkeydkcD4uVRXYF+yIB5VUexCdMpeScpIiH1KztDBMzF4ZiiJrQrn7
NvKSuX9Eglk/DssJ7pjq5tT9N++o/ajyGFTcT1ssbaB9eWbhCcy78LZ7rsuw
XptV6FyP+sdoOk/EEyGQldOskCoyVlwBHlge9owjW3VO+ZJBLdvjBLHbe/1M
6RMP6upP0Nf6K4M7TnoBG45xGlnRUW5oUOVpZJRK9Vk/qgiZnttmsXfKZrSB
equQRYhnxvrdnYoyZjbo5TOv6WZyUuzcclPJ4QbQtqEoDpWhuzR91VlDc5sY
0QxzHUCxXJYx7wTaYFu2cmeigBvnypqeITdVeXXk20mZVg1FDzW+IkvtnE5W
Sc5DDUNIYS5BemRLNZ11cG1ELfozl0SG+yvnnmOvigH9ROc+tWzmMrQGAIJT
JdoRXtM8oGjaVver8kzzJmw+J9wqUvJO4z/P/1N/hvfQBkUVf2MnMI6JghkW
IGmsyNwX47k4AaSte257VVtvpjJrZ9d7FuL5G672zMw9vBGJCPPmJIs+u+H9
u4QLhD7L6D/KcYYlx5Ka3Nzqsd3UYXP8EQJzK88ML4MGr8qkywQSFM4Sivkl
sVJgB0ExdCqHkl0BPhUpftGtTbiO/xSvZXJtH+ZpNjFYAadh6fI9XoAGcMZ0
lXIlzPfCF+o26xD/5PYBqlpqLkpF+nhSPETKY7UkCbh1AmUoShVsBZbeRIxw
N3IKFiIrG291W9VdHjOweSd/40mzohZ9c7piAywt8xFAJhGqg27p5IO0up2o
Z+DGmr5IC7C2zwUkrVhc2dClARlBx0mnmpbOonTCNGkjl8Q0gXvW1/o+/x5p
/ERvjVRQFhN7Woh/W7GwfO+DOvlV2chp6V1W9WOvW0gGAhlhDiS+ma2Vlor+
RRK5aBG8Nhk/HQ83jUEajgzd58Y+UbBSGDwy+MWTJa+HBx37WphHrnTQxU0b
A4YyZpcXEDdIVORNmWxIb83IGPjKKBumc16y8T28W3sIG6hNLTZznKkNTD9C
6J1gTwclZG2DGbOZAzeGx1aJD6SsjC6Wpgez2du9tdHrnIFIiKg0IkhHpJQx
Xx3aZAU5dcijuX89bQ9SXw2ue/heA6dS/lP98/5liM8dkMgFkpxxJsOf6YaI
pq/5Q7pEjNgYNHAgXwTnXxO8zOS/faheg2ib13LGVcPATZURXMGMHFkoISyV
tgjqvf948ZRHVjVNZ98KwBl8L62fPSk/bVLVVeSvamrMZSPRDDCQTo+osboX
lYnNPGQMeeA+BIFipUGO8W0xDajEUpsHICzk5Ib1U5B4GMEb1LCaVg+LJZEV
qOfTwgMkDN/D+VSyZ8i4VqRqeN7Wjk/+6+L56j66h1mc5PlwtX6t4KnABiAz
vXAHTzVrrdKh20MMfZj+yiujqtCC1Ngk5bGmACzQ8b5F54kKU1NWP2Lo8A2o
iWnz4p9ffxATxcSxorxCT7kN2TkP1SWBd49k+BeuRsr8TYivFGY2dHvg1+wB
xrUwrfgxIenKHzOuBO9/5dpnCvxaJnf4BuwTfyB+srRIx0gJx16n7tJjmQ9+
2jb1GXGi8lizEWArSTJpR0hBd0GvISIK6P2Q2doUutLfUSae9cquieZn9y3A
XitJjBnoTd37VCaJG/jN6WGi5vlfsYMmY8SYBCOA/ksCF7e8ujNlhldOBzmh
EDSNzEBiC5xPTLc6xEXY/iLsm4ufIJcOb4XogeZCWFWtsjyC/bOiiaFmK7aX
H2nxh37XcIohn+Zac8j9HeKLfSX55zuoy2N6e/Ty12NzOfj4PAcRnq+NGHZc
7rXjB4C3X7kU8NHtSlTbXGNDz3ZKcs4dy9/9aYBTZsYdGapwVt62ZU2wSZtd
f1HE82tog5+zorErR9QCK9ntoDK0Wh2/qlnnFLRrWZjiM+/TpGzqermKgPHh
uynJLBsgbaaX/thpJDDWZrkOGXCSkoPdQAZvBzmEpzTfurYLn5xvLaJev2Po
lRA9jhr7Tt9oqmsOyYWREZo8YjI0bkbbz8x1pNsHZy93pwYW0SXiunYRPWtY
q77tYshZbGIxxGtidUPty8K36SBm3PoqwUJvDc5VFot4qOOpC1puGoboqO26
qkQovY6HS1pR066H7403ZIh8IrUGFyPdySH5w9qJXeTt+D6UsrwV1z23Bj7K
ahvjsycBln6RivGaqN+eL5y/D0NgSdeJ1loDYu4kriINxvlBD2K37M1XmOQb
lc50A6LSfKyCMpd4BnmhfLgjcSxYPhMTU6WSpa+ID1bZdyiv3vLtJTdC0l0v
wTz6jdLRTdGv8WLKx0WyB5WfEQsvpSEcEl06iT64NRPyTsJYNneUVnrH0T9w
sLomso+6kgUj7KKvSAfvEx5Fxg0Dh5fh8po1xgbki7dFUBcp9ZXekI2Sv0R7
nmmhtf8VjVAnAs+X22WVJlag5Pw0V9YT4Bfo86rDwWaQmFqjvgz3sk40Gk31
Y0aELXujImTuTBesU8BGgVtLmJknOzx/s+hob09aVUmBRPoh8HvMsu7YyNA3
QrMOwcfi+Y4cKcG8krBry6OkW9bhNJsYzZBkxzwgZ/FJVJTIU0KSinWfOrE1
vm2E838HlOe+lhphLZ/4hYiWNJqWnIlP65TC0BeiGNcCQcQhbF/oZri8S/1r
oUX72Ntj1CVEEmChMOEz9sKFUV4KZR6m+rHIO1Q/SMy9xnyVtskRHn/M6waf
ADcLP2RnNi78q4C4kn/R9zWzzMdIqhMLtTSn6+XKkD9fvLDTzRuBJFJH4pyV
Snur+aIdWAH+iznvC3bxhxZBB2UetxBMVLqueKo8Ix4rG9LQa/OZ0VqSgCWg
drmtq+emHAwPP8qVTCIWwTMCcUfD9HLwxrmLC/yFgx+gR/Lwr/LnlfG77mz1
6VbcotqPRI6BSEoncgNSCoVZJ3JjOeffs4kRvvsYcBLoIR/vWjqDRltOoFvC
mQ2Swph+nNzVgRLd60oe8Xn0R7RIKFbua5nEfTztNyCC1s4JiJhDRFKV7VKy
40Re+hY4LI+aCS42bHJMBDBxjMPZ/D2xzEAM46DrSD5V6w3uVQRc9Ex1ALMp
acf2GYJssua3vHyNLMTQUYWPiJRPiYU0YNmRvr7ZuVpZBaPg1IqGXamUeHtq
kqBF8OvmuR4sAjcXcE3Krv+EnpKXxBj7pT2cyLrvlSfkOxLjdM9Rn/Y45ult
vvdjH3AB3/GwJYqNAqVViybeWuwwoF0h6zHPlDph75DkqXhRO9dKKs1YGn2X
aK7au/fQSfRkor6r8AvHbdyw8SRnIGBqVaM5ypqFT590Dwwf2g6q9xEPELTp
IG3PBDDjDUYBruEiVyvTA3FHCziSGURmm7zTRD+AVm9Q6CbUAt0i1T8dYag+
5dkA8VWWyyrh6KUg4eFZqyPjbbz6uZzUiNyUeos3jiFLcPJBRgeswOQwOrgH
T9mHjj9LSMs+LVoAt6KFzHB2h3prp6qaQ3qF9XOJYiwzXl6feRNv+35cIrso
r0zjfhbtbRUFDivZhkYGVG1vc94N1cLYIY978umo3elvQkzJO4VDLuybPPF1
nHDtDgUbWs0mzEOSg+v2z/I01fA5OkssDfhIJGIZ/tgMwkNvigs5zGcy42sw
iXycqwnfdeDDvx6yJ+M+mWesULA5snxZhVcYepVK4BaIHBPaZPJHKOqFJnap
4VQJXxbNBlHXndGXhELXsHMTUiFWlJmqdhavveku4xp9TsLu1ZOtWSeeqRaW
R+lSYOopGUz9k70orDJLVvsxQlObyKCS4TbAf/tv2opfVXxxIu4PekZidyIh
Eds4IjpEH3VpDLdXWg16ok5lPAuF6hE6G686HkowcaZK294AU7gfqRbba0mA
m7on4/XAaOfiUhlu/q47soE82D3iNQiC1b0uPD4aWuhAGPL4P16//qgM8dke
zEH88szt2uarfxWPVxNXpJftwSBO0FLVHsrJvS2RNl7BoVhesMpO5ds8vLGD
8urQqE5aKqLkqHxkDztRiQ6nhj2sPi6Z5tF49KEi07rCqm6SyKDmhFYIDj7r
uLxdzdpJJdiTX1ZhTYlKkrSFVKyjx3CzClkQK+AmxzK9CpUR7dZVLO4lI0Vl
xiApn5V+dyw9jMoNZahD8v49u9zZ43wK3WHEEGo3hnXTWkzEFwjbI+GrNwwV
+tt2b90s5aXaWWd8ZOD2/JJMX4PxeB0/w4T+z5GHGpF42BzxXidC0lTo+BH2
7efDR75XY5kh6EJcnZC7EPucg5nR0hnojZmk2tzKQeTOnW2mF2GqCZLs8nT4
v4TdM4l1cC2KBpJoU4eLez5gbuqcNWWmZGe2PYdYhxO7kkOOKE8rd9njEEl/
W5zUoXzVjgCF9NwD8NQnA9fIzB6iOnnEf0BxnWWOD68Apyq9Lr5/Cy2/Yk8P
h3ONOJ6BePcSZVG1FyAalWXcPl5LewDtR47Ny0gjWIJB0vpxs708/KDO+SvU
+qVTo6QWSeijQFQS5L6YwjcrZgXmmw0cxNul6l87BzP2mkkucXs0Z7lG1eiC
jlMxKbsqtygaUghZj+gncqZDp3vv9ROZUTXXvEIWOZ8349WQ/3IojkkYJBQa
xwRCGfFUaJ8DURHDcwRuaoRm5hLQyMAfAvNeRSoRlrf64PKLFtmVJwVXfkVs
DztTkFmhUEfvVM/o8N4JbrST8w/bUnJ8U6MZouRBBb7HCXY+UsRD65PoxjRd
9LB+s1HeK4LQ/D2y09q/cXxwGCaB/74pCa9N1MGIEnosZWFr2Pd0AkbQBr9y
pE6ZefPow773mRKAAbzvodc/9C34UJ4R5w8JRibm3TZ7Ky3AJe6rZ6BOdSzm
jlSaOctb6nz540s/TyjnJVCY9ytulKo6OHkB5JFF8sBm60dQdcEBDJCcFLK/
w+lhM258GGT8JLkNjc4uF9EXXQ+Q1XrEkOzeKF8q2g0sOiyxKUzf3E1ibwOO
2axKeoasdMGaxzcwjbT/ja40rVredB08MB5ZLbN0jLacgxyncsVLCXxHaU7U
k9p3iqDyue7kaSTn90exSA2a29vSMRugbk6sEUU9gqZZ0++KzZjVN9pmxqSQ
Z9/8O9tWiGM5CWVLCjgWM7rU48QHBfvqXOEk7MKSzgKJtUh6T5HMp2Z4RJV0
OL/9nB2KRWHc/eo4pWSnnLJbhjFDNB80kisQYcE8pWSumDugFxOL64ecYslu
HUdYN+3w4mLhjRj+JyXOCtCZG3zI1V+1Aq7Cbl/PickMvMpkTUm8yvLCWVP2
tcmDXaHLiMVZxYJB3/l8sLJFoIk8a9WIIVrmU7eR2LdM3J9+Zh1KUd0C/FVX
BqAB7sH61EtHkD5XeRuvCmCtwaiz0MKbxFCJqwLV8clSiWiUshKF/HgwQy5W
njHUgJ7MllhP4pqKLzEcfFW9tgDiVLCHMiSTopA+bxSaF13DxhoJ8ZvB78/+
nLHoZE4GRdAY7/WJrmjj+ai+3VfVSmxkddOrqogo2kuZWIX41pazQt6yGuDi
BiVNLFdoDoews6isK8wGHistS6q1ORwrEdRxnXBQLJ9rGh0/sdoxRHGzxubk
QXbp+/k152kHeNQ1NBHyzZ/BX5Z18EcIYx5OjY0oHnWIOlolbxHD3VXD5e7p
nQEdxQaPivTWhZO8CVBEhfMff++QrsQ38PYL1cgKVm13VLEv4ouT9peKHujR
cyNueS51obLPSEzSSnIgFCHrNh7nSuzsTTUcHUye3zVlIESqdZD56nSZ8tYs
TRUwkxgVOyCHEEk8XX0XRLXrzTcfAAdh9Mfzoz2qAomUTxx7gn+FG0v1bBDC
nXtc76h2RvkEpBkUDac8FDijUhfZrZm6ISbS6QRV7ylVaDjmS5QF+xnY4uqJ
MsbTPZUiBIZkAOtMFvT3jplyRHv+p0iKNL/pIe6HSQXqjbYLK9n2mrISdTdD
SK6PelgBgiTnEmEdbmuympG1FbFhCXx779+rFf+NKgmSbo7JylsAkNoiL/yu
3P9+JHxtwPRBNwXEskXSZqZPN6NDmrIHGC0Q2F21Y9+NuHhpOyz+LyBKEAsX
kMKLXJXq0+B7763SX6W7UyA5iwohCC434kOf2yT+4Em6GYxzX5e2aYZcoCgO
qzTAvqgj+HbYVM4gKGWgHv6UuW1hhpS2veRXJOHWTqkA9B1BqqJY0AOQJh5Y
ulj1BBj420/+uFsOIBtNKtlTk2MKd8Lb41vHAQbnfF2BMaEq6f+BPfSiso8S
evxnHIPh3ZNiFz5jlI45ZpmMSXhx0/6y+/FBL8XwF+xZE4hMZq+WwbCqfV6D
NBdsnGScEKKEhqqjs+nXrSrqALOvreTuwu4D1L7QwZD638a94Vh5q9BFDGON
3jGOKnMfCGqnzM6KT594fnsopg7QCVVK7QmCc6A47zTBEDM/5/vV1KfsKtuZ
hsASRHIxWDpccGhJIXURMyUmmCUcr0mSu1kxLvc4Lgc7DIWQ1ev/0YKQegYU
J0hkEtb6NX/syhmmeGde7Rk8M0fAhsRZ0gcbAAe3WiGTih0eRe04mpVYaDjs
brFAHLbR4Hs3sLkvWUAk3/fAeC3zOhsgFbcgu8DJqLNNkBVwAqWztU332N4v
y5fvC/J82ksDo7w+x/ga5WzlLz3UzzWu+uopDCSNixUawDs+R83oNLiRtL+E
Je0gZZ+sg4e7IBu+IcC/+vQwniTwUH+cTZ25I/Wrv5EPd2+QFA2vAB4XkMkS
vvsD3oKm+nYFgbk9vKVFuiuMTYiz6MfDgiqX/lcCt4EtOtz4Nz4Gvsqn0Y2o
89VnRw7eLCCsfQnZ0MmdyH8m4n/FAOHWLGMoiaC/a6nS5YvB+Tc/LuowjXcl
cVAbHQuYuXRVDeRShmPaRrx9EdllwvCDvLXnhC0ae5BvI7Ht2YjQhJ2BBVI3
IF2xW/tJKBVtIEe94pYAu7GBj7KcGLJBD0r9NxG3zAa0nfhv9ocodMUn2/9x
eOephf95u1e4EGQsqP1p0QtZeBsgX3xI5hoWNkSgHDqKhuw5AiwR4/g8LIZy
cFnPhfsMta6SkPqvA+XqPTXNbCg+sN0iOEsFfG2RVnxca6Wo5grK1G9c0jjY
oqXcSkqSnZeS6i/ORFmTyP3ddJZdsoLwMiA/ByNGwjxHHiLt9LmihU37jyRf
wqD58571R/V0C5OX8sGy5DPNUPtNFHjwG+IOOFAkZWPLpI9MdbDCQMv4uw3T
Vrhm+VK7O/oe6B2kUPrv8i/1MMG1SMg/3w+ET8NfoioIw5S1Kx51Cbe06FSb
YjIRDkHGrJoOCCmQDrXtStXvFt/a1nXjOt90/qw+Blnz9PndXK68X82vxd9P
AmuxBBVFpyBCv8Nsx5YpOL2AIgozU/ZUUlClErqHLIFlJmgbu51qzBjuHgHd
G8E9/nlbB/3WyQk0q5oJ3pliQ/jpejnuA6p9UzJP2Ge70Dk+MG89CDLCYB8A
Rv/YQSoOxvcaht1Bg2Nk/yRuXM1IgrkcXxqEyGXfb6ZkWTAj0mCPAvm4zfxz
jwrjM3i6gDGGmo24Ah7lJsTQcDrWEj3IB4b4tQEV+trkCRMDrwuirulah9ZU
yTCBhBUmuhes6zbR9LWHoNDa+hvdKMmNZvsxT2a9Luc3pslgW4OyBoJ6h+bb
pDuZR1IXvOVi/XsTvgJw+8X/sx+MhBPVFoyBhIj2cCJFbimEPj+p81ZI2Bnf
TiJalbfBt6n2rf774FoMWr5XwiKGAsfCKc7C38Z698brZXru/Jwcm5O+olXG
zV9St5AumaXZw2+lOwEELQyzN/HXAaHFnPjz809ZU2lZ/NLEWR3QWWGIk47Q
hbSW54ZzYZ5jxS1bR2hkGePRHsj/MQOOgLD9MN6NY9Kr5HRp5pIeryyuQqC/
pWu3+KRI3rO5LsJ70L2ATLeIArB5aP1sF36sUdXcaZttsO2J1pNFEO9hcPFd
bXmXZX4Y4T5Hf9vaNpHsLYMy6C8ojKkCNcLcrHA8RnAzG3eF7STG+++pDwrf
bvgqqxycSp65Fo3E03nCkBSZwVabN/4+43Om7VHdgyzbE5bzxFIpAdrqVg50
fqCu289Phy84PKdXzGrEwZuwQxrNlBJpsK50hugVL/ROHdi4iENlb+4hjUq6
XSVDdPYgjDHJkhzxa6CEH3N8HrXcWuJDvsKCVutlR0+FWTI+9qXk98cAn77n
r585Tp/hAmsYwzQyM+ntNtwEawWCfuLSmhuuyXYVacJbFBBDCocI8Q9CD8ki
nCTNiirumtwDUl/VLp3gDdmNGcKKqxC3UPdAR1zyHC9rc458fRuX5Ki001Eq
PlPOBb0aVeAK8c1+PCcCvu2mTJ9zi6ouIX0yB7xK4VFh2+5RS63aQA1NQu+t
QXQWG/yjnMD7diQv/F7dXnhFj8O0tTSP9fhu990clFbAiwSGL6HeeDhuXzJq
2PKqr4oYErcGgFllIW5HuzVVJkAmNjmjm0QKMF08yqU94Asit/AklJI8ZRgq
imr7P78HS8mSA6IBPs7YBsp0/NYFvBIzE25apNTSMJ6P57HncRZeRdmF3xjt
9OP8xmMqTq+n9+XA+/lu/G2baDRnVRMQX5WvY23jolJg4p/uYKGx7vg7aW5Q
pSfss4hzQ5LN9MWizshgcxeL7AJQb1QYUfmuzz053y1Hq1baciYoEw3RfvrH
gPCCZtCMy5BDjsM5a7gAQAt9Et7hYS3pbnPmaW1rylhbOLMHpGy4Bn4jJvNA
kMkd/sX5+iDmBX1cAfvZ7Os6kOyqmECkdrN8wNlvg6HCFBwfWbCZIRbzoJEj
rrI8iPAsG62yBjX5GUGQoE0uW3fJENGi9gkOTpNXMgCg0CoxO2jUIykj85jl
PDP4Z0L5nHCITWQ6JYTI6K4Zq76A63ed2PrvywJqi80tKWzA9LsI3wD/gndh
0un8M6OGAQfFTpyivDhR8fpElbaK7cjZDBMNOPpZGgKLST9mn+z0NY/JMoI6
mm3KQB4bZu3zstHdpY3CRshuQF3wUSrrPsnh/PuTTuA81qRCc5XIA6L4oZnm
qt2ttPWCodgEN0BC8HmYNq1ME3gJLs/XD5G426x2vXy5i1nZMbUMjkSZdNU1
AlH2WZKFgrsMsJbiQiScb/sdS2VKn/QQS+dEIWev5tsHzIqrDLQFhoKw7AQr
fGE/yZL8r9fUe7LIv12lyT737mt2fp49guGqu8eb/OazAZaz7ySze4xl43AK
g/PhVz8n2astx1BMrZANsvhV7owHkGiJSjx4LweB2u08+3dAJTj7/kDrjHBf
geMeg88AsZX0eu6WMzDnejHE3ZBNNb3Dug/8GGH3BX8dWpJTH/ThtvEzAh4+
X5QzPvFJn3juMueICmu/MARy1TMkOEnOyEfv8dar6UffPTsecvHQxSr0T9y3
YQE6aX00eAVEBJO3qPLacy/Zinw9BWzF2ZD3nLIjDdM6l4md1ToljrkKstJN
uAkpshK4UFCMEbc/3ItxFZQZb6U8zuzK8b0ggLWhM588PB1bHnBna9lY9FIt
yyDGhL9OsWkHGQsFdWUINhhPPzeGtmsQMS/Own4AAEIscokeXiH2VlbiPgTO
S0nopaxulA44lqePJRzRm+tq+FonEIvqQ56hn5Ji+oYPBaS3m+0RnICDCou3
h9FS1uZwomhfD5+ivSlgpGwhh3KD85jVVXyufvojZ+WXZsJOsc8AA+UyqcNx
b19YSlYwcRXm8LEz+QWSdlSJUqZUQJ5e9qwGqfIPeRwtVp9i9o6DB2sjHZLO
BqP2SN36qFgX061Ydm2368C3KT9mbQGTFbMRRUOzYv4nCG0erad0+rWoc4qA
+FfLxh2HycEhP+YwqyCEmm2sT9oCwk4S8g4smhEFTrAuil7BquMgTaPwyd8H
b85yb4IMRNvMQnIr0pZb1Qp+S2bgJ0X+bQ+coFlGx0mh2zfGztmhSlQPvV++
Gi37ZHK0yrZ3O/Yv/Kvggq8brV+NypNbpqNKcXbwS/pSo2fu5CKTUJ02sJvV
zxfjMARbHkeXe0ef0Hb0GN41p4J+YsNrQkpGi16mWQWvt9UE1TssIj/s6za6
yAe36o9h7uNObIg9i9LwlZqkSBccrkZPWLGLplKh5pwBc2Di3Qrqy/05JPkd
zF/ZRcCagGbvOQEZwYXm4RhcWWCz+gMpTkFfET4YDvzXLLBTaofLdt8pGVAl
k5ZkOFqugtufNH2L8BsUThvbPvwx2pHvmAfQQYfeaVmNwcqXS1Ixmqv+yyI2
gODdpav9xQc1H5dRSgsadtrZNZs/6/FJktyLQPci6WU52cPAKqy6yuY38tst
Wi97oonJM0LTDJPLFS7RsYb0eEE+V1829q3ZxyymMP/B4TtE630KXMeE3kPr
STpekySFHaXLz9wVW/ZK10eEBNzDPlhdFYXkcVIG65MEnV8zZEW3Pp/fUUp1
1Eh62potodhL64cPEv72gGa4+lqVdxOOXQoK6ydZvJvmJsSdOO4/caA8woL9
IVgxR5GGVpdpQg9JfIeiUMZJdpugogaUN1IB4YtkOLsjJFfyidRBiFO6+6EV
HxioJhbiclV/GOluL4HPmlHGM7ofI42/tgPIWRxPpV8HXNaA5G0fOJtk2QRn
FXPADZlJRNz2SSmYh6gqHFqR6HD+SlZbU04dyAMMv9EChL9SipMYkdEQpKs4
pvrNu7iWrOhMsk97V1PSP/1r0p50/YoNrb+FrbxHUtR8OaNR3x5ywfqd8DxY
zfFeVe6YBMz9RA8xUuDyARiWlFQIXMQYEiCQWdNw6Uhi1P4UM0HIkhI7g/I3
vVJXGU5FnbUmj38UAZconpjr+Q/+EXH/5DD/xGdYYqe9/IwdlE80CnNiIujQ
THxqAT/WUOi1J9BHtvtsuTg0Y5VYnO8LSHWs265paHs1jmZ6Gi4c4X+dx0C3
pXONnKOLXvqRjY30dnal56S1+hXQrWAPy1Ceez1xDhpT6EFlh17t5DdDlerU
Ig/cfx3w+JoJAQEzGUJ1X4iALA6c5c5tUTIPrFYnqVS5B8LUnlc7IRj1+azM
lWmi0YSp51qAXZioo8BANfM3EkFriyBdxzVYGhj77bupU08w2uZAYItoiqbI
XErP4ejvChg9TU88FTttpCoveEGnb4WZSCaF1G5STnp4C0jorfofXnkRQzAr
L5EWWSib3E4DajddoqKWqqQEKw1h9KQAMKzfmgk5ztxuDHnetKWK0SkhzdUh
Gqijy8BysUFnEGf8qdplBmqdOeuJwxpUuRwjUc4EqyfAtpPWguxaXnCxbLLT
c7LZfWqR3xHxVjlSoddYX9iB9cIAk09Z12fAa5uMzFwmGrO8dsistqb22Ax1
xmYnayr0J3FSb/WbwuXSn6e/qomCfJa1u+efnjyPZYXvBN4XM83QxuGzNBpB
NgXRCQi8B3TamsqWD3aISWEoldD5v6M99sun+E9/JUj8H7JuysmGj0oFJRLB
eE27/LV8tkIV3xIzQLdevDO7fB2wvBZX6kYMcz4LGd58I9vD28hhJaBiG0g8
2JIheOwUFMS10jVwAVbUQm1wfVSjL7qG9wgYrfnPzLYDDFE4U9CGNmAQyQ+E
tRndQvSGaJAPFU0oDAW/1gtpN1XzQPd2DLb29XAqeitVQQPftNFzd4fdZieg
KNs/dm5h5i/sV5onVdLITpJafNrVg7ZDtNTAu42QctDKiOA2kJQi+z9hqRzf
kC1JnoiMC0ID9fEi6RZEhsjHuES4cwO/vOl8QEIrxAJR9fZhxCj0fOOB0iei
3UCPJQxzJ7cLVYEMdhTRQmxMnVQ5gnN7h3m+O887xgPB7kDpp/Zc2hPyS0kG
Y/fm9TBpW1Sr5E45SjFqtRSqc2urtVn1Y/fzrhYH3qgFgbUHAFMB/HVPoJ0U
su1Oz+zrkkwf6Osi+aguk+JWMjJH7aWjbHjTbCzBJz8Gcsc5inuFtipj66vb
ixaBCFA8/QICHaEYlZHlvJRAPi+Iq9L0Fl+57HAUbL5G+oSskXisL39phG9c
Xan9LkfbweooRjdE2jdqC0ecZgHhXwHQWksekRJ8XCUwYwLUJhdHNofAg0VJ
zGxs7HopfBaIQAoP+d2F5B4EV1YIeuvY3CokGxPz2mpA3c7Haf+sfAeXGkdh
bgx80jJfAMRvWSgj+7x1D7+9iX8BL/le0AC2XhHSzYLG5ZAHvk2Dcxw882GV
HFi7X6jyOZGjqvnVFP+KyBzBOMB438jle36ohfA9JN59dzkS0R5krY9BNfCV
qZLEOVgdZkb7jk7OtIq4IRGbbZmLnJEES3ltI58qJNFUyVDoK7a+rwWhiagE
dWBBvWxNjJ6N0aU1hoQ1YWp86yU8KeZhxSuafaZGiGTAyLgpH7WdRchKIf76
xSVZgjfahKcWD82hgYZ2LqtExdaZ7YkCuQmrT9Al2rlWi4EJrGcm98LX/eji
7PdySEoQtF2NWRVjSUL5KARPP6iIaKXUQSTg999or5hYa7t9luxOcWiYo4B2
Wg4asNrpmxhNEyDRr52/mzFiXywJP1Tv1FLcpKBMN+v7YQJ03e/TGOZZOZAS
Kw8d9Rq7SxpNdittmwQvRBRu+TQOjOnX8XH1tV9Yk3KOuqGp5K5l+VmTcNxU
ohD9bNauKrVhFBwBJZCrBJahbipXA0KLJZmfzWzDI+c9eiXAeac6xgFzXmnp
Z30bHm0U7MMSaYr7fiQN5rtRkAFUTrF1E449wsl/OCYwY5C92qOBae5ZxdvB
Jy4KDgCjJ7AU6kf/X6bZjBNzQGDZ84IRmyzx04Md7TCtBkDiaPkgaIQHZtuX
PRFgoBCep0AiTf0OmFzrtwEvy0M27xiNlpnehAfNCbi7yKSVqB0CTj5e8ZwM
B7T0EYEQKw7ezC8sh/liuiuiyNasxQrYlNzrpR4jcNlx1lVjqesjvhdYaRg1
0YksyAY2AeKsZJF5fQnpOcUhntZAUs+pok8fiD3+bGHXETCA0AOSQQrJGoWq
KPwKj623KmSeQ1Yv9chDIkWDc0ZTmOFfS6/n+25upvA6DmWxFUS3Q/nI3a6c
+DmZzwWw/9Bv3AnxIXmLrPxAeastuCErdQYXMDzuCbssKdhwpEL3LZikeeKw
eY8MHBH15FMJi7TwYVZOinkgiizdM/URjkcAkTiK9sZISYUSYKLFmERpcLiN
1GaehPDcwwVXdZHnEk8+5nnI1Mkyfy7KvNPeDw6dosb3U5rEcrk1NX1v41Os
BMKKutD4YAib5cCbsEeAOeSfNOkhNAnxTZcWh7U/pF+IeZlyo0fo0rqQ/7Uv
iYzaF56qeTAweT+xhUb5Ai3FN7C+1pHPjEKNEodutcQ6ZSkOSzvOyHNk6iGa
i2lmxQUCNJupnpXN+rY07+M474TEcIOVt3htyy3jfDO17TbQZtiSIWk8WxS7
xIg9+jIOoIoCNAAMyxL5ByZN0xHn3FbTQ9vlj3KzPIBb7sbXjN1g6wWoHrJu
61aM+UqY4Kmk1sXl2THMNKyveY1ZuPk9rU7JctVvz5/oOQ5YEUVi3xHv2gmS
0rT6aVTnLqFbHa+prkI2FJLXIGl9AbzuOp+1d/4ARA6ZT9428Nsw6oZawmmd
Q43eg3MVxWoiQfAfcQz1/a/dfAgiCjKhoE/ANxB84Oi4G7fUzOD3kMk4lZpP
bevjjm5HyBJS9E7ILx8vJ20GivpDBrI0xHnvSajtmMfM06LuRICatoC5g4gn
EJqbJ4tSc+SDyE06XxZVf18M3pdvEUkZ8XktLBxBkUQDOcUPnYzLVyAeBtZb
6CFsQbBRG8wr9IMqdh410jUSsb4vQu+7v9NyN9PcOADU0s4yg5imNGEsAKhA
MHQSlX3SSh6HOuUlCiXsz3ur+Zy+N/uFkgbBprrQnvHED2hGIuu23DlIRI2h
+65XjR4mccZ87LXsa18j7OdpgJjKmLA+IZhtBQ2PcyOFt5FkCJehxDvn+ku0
2b0+rMld3KwpB8Nq6/w9n/LN/Bl8XOP5d8/fVRVRF+QWxOlpPssa0rjN11cX
SKvGBJvK3FzCowVI+1M/WLn+lYUA6AfPD3vzFYnw7SB9Saws+e0/mcUidfzw
zi4gYo6v6pB4cGq97RIHLm7XCPPuvA3sANdkUgpoJwcCUwY5r+LtsfHlyXxC
yLD25RdzFZfi/TlbG+IPJbdPfgFIV5nYJPLTLSORIXe2pgQxKAsTcaTW+xuf
WBAb+WmF9NuOxPeiG4U16m9dYev/PGse3r9W5QzOnOQHMaZ/Mem2qNyEaIVX
RWgGG28uY3OeGLmyNa1M023B36Btd6GAIRCPcKurQqMxLU3soyLuhi2w5n+k
UcBVLpUv9uk3SotPy/3ROCk5HVtLL89HxuZCkrcGm7D/8ft71d0JQzkz4bSK
w4DNaCBGemukOMTS+SnAjlbBL0ukknBVQpHXdEtiHCWeQ8CBSeXbNfPqLXKL
7J8DwuOK6cXWQy+KBJkq5KoRYTZHCwsbq9fXPpOMUf+g9aehil4KvFkQCnY/
TKYzsHhctTKj9bXiVeiqnuaFZe+r1djRj+XuklEpVNF4+LHAKKwUUnNoyyuc
07VDjnzBU29/9H77DmS6fMB+7HJJEMi1CQ+xxeeTJJ3ee1n7hEC4/F0k/Qfi
gJfdbmsHuIslYaJmJf/5E0nUD6Qf49Z6/RUcLI70TbdYNtfo/NFgSF9yhBP8
ghMb2gNY4x9+tViLj8p+IxuBLexx9Bvi6KI2MqlaorB3lveZswcZq81UFfCD
IIOKjKp8vE4AIHaZvxyQvgAmc+gxr/jPv74A2es8fSKKr0a5y+ijDSI3NPop
8ANg4ttzikkS5xT9Uor5UzwNmwbYtDiJIKofI2W/5stNB3ULaZ3dX0uDkD20
lkT1XkfKPYp2Xg1Obvd7L/nlM36qC4gbE10aTwvUe/Ktj8I4CW4oQQ3yHt9n
MyAzM+W1DX30FUSBfLTJS8t7YhiECxS/Y3l/AGj22rL6YfWEjguHoGzkrbnQ
3/98ptwpFnjT2ZOp/8ZI4zqcOOmZk0JBGTyafZLvkEe+jAQAWOeAe1RuYkcB
0V/ULOkzRW3+Or1plYamIF8iytXoxyC1tVBIbjBv1dDtoqU0/TLnJ/1984bO
ORwVe/d5Tkq4BNdZXEYlRkzJc6+fJUs37OEh1S4ltdBqCBUJC6KHngdqDzWY
lICpj+1lbPL8RFSZiJv0/KAudWjv3iPOG1ETyrgBQUNajdQsGV/ZvetWw8NF
eKQ5fcPlfaW0VpFZn/rHdZtxOIGf1/I088xI/SY6W4ZadL4rQh0tTS+CQtZI
V8XUJ0PrUfAvonux1tKx22vpzqz+gtaCVb0sZi7aQQ6SwixqUYGIKs28ijCc
dDgZEdVahG1G4Wv5UIZ37MhHLkt0hQIR3lYXBNtxsuNY1tzNkpUDZ3rA9JoH
Gkftj6uNlThwcvUW/6cGUi02Bj5dJ+17y+cl/nZscmX8aOGuD+vJlec0X5yK
V3sZer24CFCxOU0v9vUixVKfJh6hA6U2z4UrtqlPwGbjcJkP+k3fn2olro4z
lBNOHoOFCYFJzao6TR5SjYkhMzlnVsOkutgieQzURdVTVcVs7SXbYEvMDqrW
yKmyvB5r1weoHaIqv6FIyr98eNdBeWBQ4BOaxHmuQSmQrHD1V8usDZqgkkDH
2m1EsabeXrv0BL+TDowf0jgzOyFZblLrw5r85Z4LjgbxKw3UuMv0mK1UfRBW
WhWOM+vNfcXUyCHrCqAccZC14sU4NMvmc71UojjKCebeAZEvJfowpA2LBsJZ
yuXTvgOL4eEFFYbdL/lZR/XAc9Dk3/48kSKbzdWmZxaFL1U7chr4nb9iKHTW
Hq+dDLGa2hYyQ3vG0HWszyR832at8FCuUJp/R3zaSvUN7CiJd6MrMfVbmAqh
XKytl6dQwZXqkcVnTYJFfSFZVSCbMmCpmTlHefByDYgqSUcljNFXshNhGOAr
FhUmUb0eifPrTho/Hrh/Dr9nACvy6gdHfuYypc9GDhdzdf33MePwJnofJC5h
B74L9mc7A0mVLjtbzS8vFG1awzSDTsawmrYhJ2vkNgZlT6FHjSmvE/kR2XU6
zM8RAHfY7cVzEegxsGkLrqwcaVxshmk5ZumgFTHdrP5XnJnaUX8sIyO/RdpM
mp5OXGqMO3jalGU+mbdZ+cYsL2deuI+DaQfTuzev8lea5qL4d0qEvnRiG4Af
hwlQgYz0NGNcB2uULAtAWEnJ7qp5C5Qaokr1I0QXYxygaekWE8inWK235+Ys
MX+91VZVnjrbOdCExlJmcdVJSvlTAABNZZnw2CF70UefxA1zym6J54EeA2sP
BYvW79m8RTLHIVNTksmOZJh5/fFI8fITw11UobOwXUt8WxWEPYfmUxYnidNG
pykGYZkXjFl7Jf9AjQBuBRBxuFrUwFGij/0s31PrqwObqKL9mU4EzTHoETFp
K/TR8R6dzAfTJCTiFvq1wgoVnCxIjo+fUDbh9Xx/OvAXg8mI3I9UlAoefTJZ
rv1Cd8LNjQGuTEWYkQrkiFQLdljrTIWRrCJhs2DD+dg9ULig8xOvr1F0sBbq
fCNpzcvhyFx1fx+3tjhUeLsupcOuAge1XH9DUn5jDEcZA06XOMCYhxYghGbA
T/qaeGlOvWSpDLC3jWiKEDaJSYF+wOzmeoNq5LAyHZvzFFMbJccjqcui2xtI
R7GcUvHPCaf0Un3ePpoDhOQkH/1y19IT0b+EVp20PfEKsFbDnVz0HxHReSLn
svYmQp3Pa/P8dXaXl7bJz2ptGD3zcrLzHGwckhJ2Z0eceR+nbqwdvM1lzSBU
thdMYmSWHO1zksSU93n+LUI62mCXoSNv+31evCZo4N9rqh+JNRXyoz3Ygkq3
0HXx8AGmxReRrlKUR9V65tC3MTB+EbbJ+eENc+YmiSvJvZ8SWqDdHeaIeV19
ux+eopX6zW/KWbPFBD1qll1Qs5hVxcMX3jGhmVm8naJgsNhVEFkQTY8Px8db
ERzEDcIazoeeoMHGK8Em0soM/AsUbz+ltpYfBx5HSC3LeqWg78GJyEPOI/EW
+/xJPPo3hefkIwvNqSLmoQWpHlMmstqaSEhK7zXTd51zUB6wub2L7YHS/PzX
jvvGg3PJbW75j6bNqt+t0T3wU7eH6Z3k0w3tbEXzV7+iAC0dnpUe7EPt+KYh
alv9slolzyQ0j4AGyMAiOIIpF3ufIinynNVa7gs3U08WQ91Ri0uhQwhV4TGX
tysrS5xRrPIzw3ggCMR4YxaSStZoXXWnoXyDKMGpN1p0IWL7MNSs7K5r+q6j
3T7DlebxA0yooL1W7U1VELjxjm/MQYdGvPRRxWkdtn8KZfGEBYQoiSngNclC
5ljk3BLt9pYPEp9OktASjugOmywLugMTenC2+Hr8dyCaxs6lTd6mZNHX79K2
RxqaiZ90QtHnEnuvp00B7zjkQgvqxKxrEjketV3Ny5caGMgde4zARp20Qz5j
ltKcJXMX3snbw3LeV5A7TnZ9vE2wehiBpluxyW0htO4RO8+ejA8Eo7XH28Lu
9PxrlhJgrK8XumEa0/v5r+cQWnuI8L9lBl8iCRn3Vn6ilUTjKJyMohCLjZYv
siFk4mmZCBrLBqMI4vz9BT4RbD4queUR9ECe2JtUsx8sV0XUHGQWzrMGf/Y8
TKch8UUxue5kalY0J2LnMclQUeUjplWOx7OqUZFeiCswXL4lU+n/ydbeAl2y
ZkBffBSIbzOzmXFHCtxqd19Cg2fEO7FsS3WVjnvEhDxo7j5wmngdb/5pAKUO
HKyj+6SJyazncMgiTrX9j7suw0zZAo8mBJfiv4qTa+xS/1ciCOmmZRPhOM16
jYuKXP9Uq0vITN6JWhv4z+e1Lpv233Y5CK+LT+ExpYkRIYF1INZFMUVBefSf
5VEiaTbcMD5ETiVWTFd4kQNjNALvSZvV2+aYDn1TAHLEG4mOTM09l2q/Y0FL
ocQOQErxpL7/X7Td8cj9+woQWoJ8uv1oHMn+LvjRwX6GJiZo5Q5rkpVFKgE+
QqMM8Vfw0cawH6QVIQ8Rp2HtQX3pv9ARg10BXfWU+lWIz2lcvJDuBzdpl7a2
SzHtHhbxLTi6jFrvHsDYzJgBL59sF4RqPj64csTedEMXAvGlSoTjND0+dI1r
4bt+NGjAOL6uYFNrsoyGiYvPvxVT1uG+lkGxXf3+9WYu75iJAo0tvwpHu0K6
zXo6xfe8Kuewd0uBoIHZLtma4pR9ccTPPbhPUte+4g+WAhTMB3k8HZqea8nx
BxS0n6HLkrH5J9jNiSB4J7CrCGzB4RDZtshQAsEhj8cSUvfwzQCxV/Sk5DLJ
D1CW0t0L+6y5qgnesTOoOh1obvGKjcGamAIuPiR39OTidfXBR78gtw1t3qb7
Rr9jPD4JQVwN5qbkg67gTvPuNTOenzw729YDU1aF/bYoqO5/lboqMFqI2Xlo
NNBEnFkY7oDo6OnC9OkwSn7bMWElQDBaJ0GvwSxI7+TIKhv3sN7ecova7Kmg
Qyj2WzdFkcYu+e6QHjH+S21FOTToY9Pk8hxdb/T//Gz2WsQ5UcFd69csv9wq
ZgPB5Isa7FL8uLROpDVIVIwYmnBTppf0nGClqlvn80snSjnX19H7O0uQzsXm
jIW4dIjjxTKkdmH7fBKQo6Iqi17cGIlAbHpXLxfUKNRigru3jMIAl4dyquJB
VkBzxjFONLh2l3f8YTgJChpwbTrZMV6kxuFWwY9JEjiAPkcwPKDuKKi91M6d
MAahGSUW16dwjsIO4MQI3CBF+4A6d88Jwl0gdU9zT80IUjqWLR1fGJLDdOsy
Vh58BXmcBi11Gm7oO24oy0BAyn14YmJyvvfAHUTXTUMVopAHwq4NKisYZfs2
es4RQB5bkJ1nZmzgdTQfb/VZYlsZ8pmUt8yWSgGPh7386lbrHbSV/0toVEwt
cxbKn8vQHF4lnf5GhSuTrob0vuBsC44lW7JlHjGmcaMnxyyulpyBb3s+36O7
SzVZ7I8wLf/v0r3mhgpfAo5u6b8VyIAfTpregYWiC4MahIEtNONOjQhEF9SK
opS60YPXkGrvDZ3pumK6o2fZXGcx0MSiyHfy5797RPxClhFUtT2ZQgfYszdB
5hC46igwDBYn1PusFE8oTNL56YTJkCFI54RnLujTETDTAuhBn2FNjof9vgrT
Hh+e6YJHVFBi2y3w6tEdaPDnkehHlYe/l7epaoXGTXm4hu0iU4T5o2lJ5gld
wsf+7wK5ZTFRJE/WkSxbMqBIBv37zfSHMhQ+wI/dlFGocW3TGwtI1PZ/QDn/
tWbYvNEbaujX4fhxqtSA/rWL3yUumfs8/+CprIf4vH7drBJH9ucupu6Mo7vu
hzMmjAAF5MV40BUlht0KCYPLyugvE62w51ibeO87FXePracKh4g4rY+hoLAm
tb/mjAvHr8sgSd7iXb+SJWvGjCTbXx8Wlsnk/MxhTDO91tI/sH5oDZPDsDKM
nwRwaw76dY48DAyaqwn2LA7aAQVfaTkTAi6uvZjayVE3Oig3olJzvw4pY46G
VaNkBsA/RTzNeYIiSBDgNDMl9OE2T4P08Nsjkth9WZBCGh2f1Hjd26dTS0vS
BCz8tpuhAaQmXj9PxwHu08Qm6fCjNkuLe/1IPoVNvrw4rXSeKtgQLfuyBl49
9+j5oj1H/luELybXy4d2716TsNfBC7FHMFKHmiihuocjfG2x28uRigyDXaJj
KpwTZgscFCTla+3kgfLTuvkFArkzfwHS6SYM1b0xI/SpoAEk6GiOC3ACjDSP
hsusE5BjWBGQf5s3F5/idBl8hNVvea8eslNpt0AtHncgk/fCGt91OufFJZ4/
lbpyAnttWgVoCk7veaSOS7KzCEINJf+JddX4OHRzzmX2VolVsaiXpVw1fuKa
cv8fjW+dPONTnyg17qjHBYIzFdu6OtA8nTjVdX55sHTsu1gE0RFxwVA77Qo7
4UB3ceE7ur7gGhRdkcN3vEY7bp5W5KhIkr0GmqUA+i0ybpQ+IlWqy0eENaxp
6+PpEAQWw97QwneBBv8bTsP4MTLGPe67vA5cRg3pvjjAc2yqYBobeMsoQhrd
E+cARFPeR8FeyNga0WcY+UhJ3HVUxcNmL2+FozBXGHmS4wedRoa8jMqbnX3J
YDU0BSLr73Nw/1We75cuV4jilQD3/jsRsU16ajZE3NBdYAJpKoTrn3IjK+19
YFS0l0NfZv90tAKPL/WcrhT8bC1V8lZdy7Li+JDsuIACkqvWUHWvzpmsve8H
36JAYQEeGvBEM/KxpFvHA+HE4/Dy6kuBpkeaGwqNomwrjTwL5i71BsxawdVZ
lcTAG4BGQK9TJYbQt38KlFmLKjENjkiE4t1+JQhrdZSLGhnKN4VNPtOM3pVI
yKhuWzUX47kPWYpwznO5wEf99aLQcO5FC94FBtpSt2r54Koz2T0n8kCytaVJ
judGm+Sq2kX7r6qjSXxJ11LUXsejWhNCi+2ATzbwKlbdVpudSALkjL261TjY
+z19m+PSSR4XLnu2YpfBjfy9jtrPB2PL2UILpOrIhgQWvtGfSYBZh5EJLc48
s040xiFyLuA3rTiwLWyUBweSqHfUYiKO4a1PxFd8U/1mjdftnKs3OfwH/W2p
ov0KtcXtSXfQchdSpZsg4cMHwUpRszJ+FI5Ge/DRkgJj5b4+8/c8M3FJGuPO
koZr/DM6a0Jke7Amw545QN0Ap2/9ehkcFm/ePI2k5NbEJo+D9APjomDlwS1g
o8R18fn43AXPZXqsvlAKcqT0S4+QZtIsvWKTioKRewy8/qaZBhE6RZlQ3EOR
wt4MuIjqiL72MIGnl3f5fRgjxRPX35fiNe6cGtSObMBAnCvVyaqepA4EScNY
lmj6pk80kMEbDFQ4dIw1Tcr02jYu+HGid1iSvW4pc0Y/BvZHoO+NbtfVgsq6
I1K+GsDSz4j0v817EtCb2DupSgwoi94t3rqb+5O4/m/Y6AoG6tlgTRkw69Fm
jGgsS3cgfCtO2RCe+wUeCk1jr4sSA5ygAPmlZs/yCjDg6RA+wKtM5hWYbXY8
U2CZWcseX86cb7QJSDHntf8nino/tgFVYu6+NIDYFMud3CIbT/ORafJ9fgg+
+S4B8ue1k/Cwnb2Q1Qh+w+2Ul8zdSkaBhCxVlp9/HiGh4/8Fa/h0eLEr+R6s
0WD62rzo8Sgcit8c/mWxF+a2QSJKta0zH6pPSE6jvbupefLdZauiRmNQ1tL4
bIhmCLymm1z9ss2Uz3IJOEoPJLlhrUienKL5nc3C1/21HQ4FLNhjvCxHrohw
ut9GhtFl+8Y+fLc83EiIqdusP+zMMhXPGICdyw4iNYZGO+yYlvH7LbrLwz2g
2yV/i9E+1FUF2zWIEzJ5E4O5i13ps/bU25UieefFNvC/6TujekE2VeORIdPm
82Tk2yraVXbI+H4NVYe4nqkg4uSEjxC+EV3cX12+HIBT6m4mWz0KyBCcWCtm
LFFnL0A8fV9rw+le3mVmHKaP6/x5oHJfE4ty4FAafVVbK/Tl8G5PFPYhMU0w
MXaYi7+HDDtrV6hEO4c3sz6ctK0LVvVkBuqfF41olN83RZN45eqTCkGrniBJ
h9PxBTpKfHyvmVUE+ES2Ev5B7L9OrKIc9dyVyyumBbeAHX8ncJ1lPczFNy1M
ay+hS4/lrMsqs7GywWjP0fSJE9AUqBLReplJ2uZUZblPPRzx/gzbkXKpLdUX
0k7y2paFPANNf2UAm4xC7EA6zunJg970iiegvUnQVNzD3Q22O1EJpboj/6Yb
y7mqm6W5GIxDohpD/cU98O/SLhfD+dYpcV4OhiKg/mCaqnaP7sZo99+J1+I5
eXw9mLGla2UkIbUEnmT5t5KCeN0CEbYV/EJtIB2n+zSWUt992uqOwmz2xyaI
yvE7jJPyZl78oXqLpUV0cct+rIg1tIPfWM2uRhGrsqjwTCt+PmFQe259rlyU
f195atvf3/ep3i1vtshgJZ4bEqRcbDauPUOwEz27Z1CFzTEn+Y4+VAd7DWhe
O+v0fE2sqKJGCMwPpklKAcrWVFDhb6XozZdZWiWHegLiy5UiTiNQlE62BErp
TioPtprcSmhLJ5lsH12gqCZvDB07jqGzzP6EAJNNLT6JMKQQHSUcF2XtZpxI
4MMhxyxEoVcj8jgTzCjggycYp4dzEIB6AUb8ICETgxNN1q67UuUllJ54HKvR
xs5tjjtEQIasfi1OB/XQSCPl/o9gC7+524OUdf8pjRKYYQrHydhAYXnKNtwL
3jrrsv7w5pAqlrdFBVkpwLpgssvO8OBbzX91mrqRE3hCn8YUqCUnEDJXpJpz
PlnAQ7HVLfwgTv+uh2tH5WCs4OSITDgbdMkyUKeqrVOM+SD6YZYzHCY1wDQC
kDJan0cLVSFeJGNK2yd7vYvD3z534VL2zwBrVTvvR7msoeRZFR90KDM/mqpV
8J32pHlVrNy6tHLvXlkxwNpBNW6pDQj2+g3J6xVivXkx9M+r6XMHXPGowQUq
dJe5WqP1e+I0qhRssvyCctCDWQMtOBrhVqFB6babrQA8vxCMXDHh1NqTz7nG
FVZX1GldHdHIgDA4gls/XrkQeQomXWsZshmJD4id1wgEyGy1HBOw+GlBh1hJ
n1EZG0Qh9B2QC/1iGCBYgm1RbIIq3CeDEOuSaik3WEpzrI8xtXW5+ECrQqhQ
FmTfwYRPSogZAllTuGcy7KZ+zCjP41wshGoqN1tgW0ZzkkkygExSzCCPRg1e
eg9QOhlJk1EBGC4gQuJyIPbnu9euSKVgR3kq7PAuTrp4jFUpdbxJcfQp9aHr
6tCHJFyM+8uXMnA7mOmE3o2G4f6tND6/nHZefiEPtW5BfeqslzraNdSEU1Eq
D4Wp3+W/Y8zc94ZVk510eB5+d1Nn1uOWg8CH8ymV9F9qI8ZaqqDrALZlK/2P
sSjCtcutPjTSXnMK4YRzuv5kgn3boAKJNQvmw2RZQBGKPJ7LfrUTVIlyzISn
SqOTqArjE33++3n+s474tudJ01B2NApVFEhBrm+AVdhVj+RxDyDjAk9qS9R4
LyLKH+zqrfpmIAiS9pEvsw+hw03R+fEVuWSSql0zEidNrGVrQfOjio9B1/BH
TENTb/1XEQ5oKwBm/5G8cPNjziTmdpmiM4kE2m28Z86JeaQK6U5j8Y1ueeby
e35RA99Lb2hKC+RGyNlMEMC7tJS/BY/d85WDEjmlt/uGaPb6Wr/n24GijSkR
HWSDW1mdLojwGTsJ8RbuqdwkGjTWkgKtE7hHPeGQuefZG/ythw9J/mh2FKST
3NigXJ/9MR9Iih4+wFCVIVTyZXo1IY4FeHHdPiRuhjruzAdzluEu7/Ft1aoH
xm28CA07qFenkQkBvt9SKb/yz/Jffy3B2V1M5+p2LEQPHhcJ5jZPgZK7qJQg
Hjdmfrfh+Mb9rSVXbFyiJ3FtpC/oKN3iJhmWMRvZy8t6zPWpB7dUqS6D42ea
LIPC8oAXxO4LmWRIN2A4JkX7KKuTcQ+BX3wFvSvGVdSRz9hGfeUvdQtGsn7b
zUXwy3mD8/Bcb8lZmjmNpJW4ZX+xdW5zaN+9MbCIZcQN7fDRYwRIIECFtHN9
I8ZyaZbkZDVfdPue/qaiivgxvob0CsVXg7kvDidxFWyJ5igWFtxXORakCrPh
4+xsNJM1XYGn5Wz0RLigVrDpjFMhHy8SMDuKFWNnhZ0Fl9rWe/HFSKBDNMqa
iuPoC2w0nFD/WdD8JazXsZCOgun6B5B6pYU242Blx65pxHM45hIqJUQWfjrv
OOWZ8uZrdY2q4WBmD70LbcereMYmDDPd/vWpMP7A3cAQh4EIvXl1TpnK1b6k
g7PcT0l78dsG80p33nz1z9JBAQi4jTzZBqTu9NmnMwks81kmqq8iAHKuOrh+
+fpcPn+nyeF0FoPh31tdhGFtlGQsNEMOHLcHIKE/0w8m7No10tjCKnALtcxq
W4EqSZhT6pkrAq6uCiXTprx85SraOyLJnUk/0nEQ6dsJ5N6uEsHC173K9PxM
bvCnr3GCKv0KSCkslDDethBbaJIYtjwCH+9xz3o6dFYheQCT2xF9z07sMycu
vKRJd57hy9Hbb8RhgIRAkI5kdr/ISWbmDTkW+/hwuSZhxjtq+9NFeUK0nM2u
roh4EyqVxNbLSSaj99uc3ruOfXFrEVGXfhswXCk1xqS/KVMv669UROBulbxf
975pZ0Dj3Giz6c6IJA7ZnG4XGjq9v4jqovudGC+K5dasAOi7tL9DJ4TkNrYS
blzouKTaDTRGAg6cCy8u01yjCbDRHCKQ5qoPt8D7BvX+9BJqHcdg7ihZIsjG
yOvFqVRL6BqTvw5ZG/h79s+5vWVTkIemCK0i2vtT+zHukcLJOFwcln68vN+q
Kprf5iB43R7aUYNGZrNSCTzY7yQYAcLWCYqbk/7NJTN3dLPCrBuaWNYiwtjP
DlosfP0IIVBSzd0Flziz3Dstei//+xGCAtlPY7iM2lSLcscG6Sszk82Fbn34
Fwys8U2/lgqeqYPTtLPgTx5aElWwmj5IuhgqyMjfAraHyVEdjDTdqAf2jSBF
XT9PfgPHBP5O/1/avCVRqsqA0C2MQHDrps3OvL3aYbOhT56TnoLmzdTfKuNo
VEn3FBdDq28VqP+QZnY8S1L/aFVeJQpS9dJDtJLe561YBE5cfdGlFupWMnnm
QKt0GQdV4MF1JKKyCIphbS7V/YuNjSLiICmBs1sSmqZkWYdqnyL29EO2rTs5
TssRF4Qk6HeCv+qyQrGKohkneIXnXoUzYYNaKPCyA8DvvcrI46Y2iJWV4m6e
DFDSFPobVs+6UQsg6/Cdgb7I16ciGYA46gJOHBN2amL9Llr791UgeUCeLEjJ
P0ajLEuD6fB1Nz2F47IQXXzfinNzQDjpMJeNfX6NyBXY6lIkv40i68KYSxbz
hmg3c1S+qk79ENoBLHy/F8m8zM4iTKGSrHep+KLXLVZO0eL2qSMLfbmxnA24
WJgMsuExVfZ2UijwvV7TW8DCdxMxtvijiUQN5xboltT8bMbxe0g/toi+utEV
Ca8X6gwmFmMaQE/UvzI5X3KnZ+tmSogVPlbs2TwQkGcHytQ5l1sRsrRcAa1J
0dAjZp+grjH/OndxE1mzI+lQ4C8KLEcPORZyGZX7vyAaM2W5J4XD1nFhhVA4
P96iYJ/nsCco3bLLz8GuneZze9mytGiiOrorFVZCCk19klHmU3K9mOlKltz6
a793ZuW24DDIjdskcXJe3cOHPQC96oXlnOqlGFjwyfOproGq96gl6Y2AHHFX
okNkLj3f8NlNT0BB5b9iI/y5HFxyx7800sXUjGr3EvoFnPd0CI6BwRxPmYwL
uzm624h6QnG1qEedhakebLYPDJiB0NH45ixckS/7+heQegeShKQdTsm5HoIR
akBiiSx1Svamij1YfSA4NimvOpqVSiLySztA9cXkBzolv23gPfbkXwQGeh3B
xOfIZmULwGW0fuckXagpBhL4qK7hr5JjsUrLbvaVd1WJLDmSap6ytP8Ermb1
ZBEnIPs1fTsWaEcQdYzOmvBnOzNHhRIfdPDiVhB5rJn+VetNei8A9Jo3s2La
5kUBKhE/SSU3EhsucZwx1/ADZ0sXa/7vaFbEuBx8Nv0C+fo1nPmXQJR037DX
M5THOfmeXk4vkrzkN/gmdFWVNqvhzy8zZXCZNGOfZ+rgNCdfbE3dKYI9E/8U
mloKxySSTGEtYY39W5NvkoWpZ/PwHNi08hKUdUI7SrNHJgDvkEzSWChSAI1V
abgoEyjb1cSn/pmQTEk532Iw0xqxyWnkv40VPlHYBzx32qheQUZUVvWVXGX1
gtCEA3IzYm1wvnciIex/lQtn456atuzlO5NNl4ad/JjMY9/mkPpCifnI1ITy
yV558jBHs0VPmmw6RcpTs7Sp9CjfAl2TgAkr9JDIN3R8IO7zAXhY+QO6W7WX
ShbAqOsoi4Wbm9YbVoNEYqO1rcnn3y0CQ58zTILZ7x4bcj4JEH3UMdrlh8q/
D464RebZHYMm7lrgG4V7B4Ulb4QqC3iR/zeEMlByyuTy2mUbbT5SDC2ylMhy
KYYl01uLbP2WpwOPy8R3jTzsLrtm17/BYJbe3l7FSstmsmy6+HOdUxzKHBF4
ezqzDJWZutGiZDkyrn085GWSIdDtx8M7WWhbMVzwq7pxnW8+VKt0MTpJVuw6
gOXdVpZYztX6l8eA17PyplMQd7l7ryTsAxq8E3RGcnqax8L6N2f2z2SCJE1w
jG0ejzPmGGa1AeqQoCqJNrfNBWSdyJ0n9Ly64HYwSHhRmQOSpBty3LAi7/1V
nG3xfiI2v4c5lxLwS/Zc99DKDHJzxauTFxVJ2HLAvQOXC1BpofBVXW5i4TC7
BNlZ577cdx+vs0gYjxO4Qz587ye5KTHP6GTDYfPpAh2dVMdIKUNkrDftn9Jb
1TMteOVUV6D6WkVBJ/tLTjshEZtf1lxWkNhftjUy0JdI7G666WCgNHR178IY
75KaAljsLh9Lm1RJ0mNE4pOvg5cF68nFD2QG5jwoKayBJaioSRy16bbKrcA+
sP7xTfFi07zh61pHJftka4jWUrVzvleA1eMJ+ldZVIGOybboYeVng9RIueWY
nr9DyJYxNLiid8Dz9X16EMa7mgSbBHR2dAb3M/kHIrmLWKlQgiX86vAHUFaC
bQrctJN+PFR4WPdCz/NW1noBSuD+m7ASMUMYDNOgYvHks0Hh8tzt9PvIO09F
M8iZNF0dImqwlC4rofmOqhCQ+Zt/bdGgnpm71NEkfH5XJmbtUcE8MxPpp+vd
DAA/po84cSLmwxbGoHeTKtkQeC1GYHukf3uozX0mPSXWXlxCjXwrFXpMH/VQ
TY1HGIxtRF/wIOQ6QOEOayEJ9FcqcZGjjkASP7PRtzvJGrombafnPoiG+9N7
kNVyS+UESzMMEKPZbJnA42M6BbZVAqg10OdW/YnOWuelEu4OZc1uP2P3nIBO
Yex2fNvCqyT5aBlUqfTQ0szF7YuH3Pfx62PU7QP3npdf/MR5oDrm8d94EXFp
XjYcwM4iRdXzmS4+lvXh7WeQsym9eMD5m5kXO7/kA39JstAuRZT1oENhmM1K
P6CRpTCdrNWyZEt4+Hz0WV3W6rTVllsxUmWUcyY9pYWDMXktKQ+iwZ7n/Bbw
FGSXXl8FMS1NKxvs7Mc+CjRa/9P0k7ZYdtN1qt5eDx9TSdAOjQrxHyAjTSny
YFeEoVh1Pn0z89kEqTjdzwxHCEiHGhxxkPpc34ymUkiHgY1VzwXjjBy1mAiY
TlFqu4DV5OttTz+wS8tHe+V+JpNYMLD4oVfIZM2CFQGtoKw86m9Ix5zHckQC
gQ9BXIwHD1UqgsMjWrj5KE/FlMHj8MhQVaEcccuexudFPhi0wCAJiwo/JIW+
etbj9kzz/iERS/IOaubcOe7PMGaS5z6eh8WBBU/RZLZtx3Lp5vqOcalvRNk6
nLjJaLiD2W9p+SyjNQ9WfVS6YU1/ClCDSRvIVa2UHFM3+zapNlFhver/JVvi
PhGHrxXwxwWgiBSMqM+18HUUy7irNDh5TzOwUTvybEU5Bb4xrNJOvX71strt
sYP8V0e29dpPRVwbC2dZipHOxaNCQmzMP78BbhhuZKDOLiM9/sX7/YMEEHK5
EGZPgTbHs8myT/4+aGf8lDD3EY3xQ73KTeYdKMiGHUuEZ5MJMnM3MoIyQMyT
b4Jp08rBttY0CxZNuPKzlgI7U8/k0xeUuD4495PKI5X18KeeI+j8thGhekD0
z+CtvwOjTGe4b4BnVoy7SeGI52UTczwVA/4FUKMNK3qd1jAqTLon3B5zgmog
sgxNJrMe4byDeQyySKDqaYFwsg66H1FaZ18pmNtknVY62Kogl44xBSwXypzB
9ieOxmOgIPGZWqIm5P8kB4Loc4IPXFnhGT18XVNPh9mghDkLMa0nLkB+mbv+
6Yx5TTNjyAohHUhAmC/vZeAb7h861bxO/kQENSIgxQj20fYueaZdLZ+wLrSd
YWUYISGI1wyPO9XbvYY4pHScn8gVafgcbLNInrVzt97Glgd++iRLMgnB3UJI
ICXbAPpf0KLB4w5tgeY2UH5ZzIqbD6+J/10bD0RfoLN6yFiAIavxJnmfadNB
n8Mcyv5T4yZNwZolDFZ7zRzXKSkyyCfiE43a3UXgnlOpW6yxvEFFkPcE+KRQ
GHB5vIJA6ApoXDOqt8radmF6AdqOswIJElgaJRDsDke8ZE09MMuB27e8bQck
zRsdwYjMrGJhAp596kgWdf36ecreBMlqqR0g430la8JzaQiEKrZ5Y+xR5KOg
u8QOdVntASZx9R08o9iaTqDsw8E9Z6O4D1qD+bu1oeGkPCPBcJ1/yINMtNoU
WUmA2WPM0cLfLqi0czZSbLlDeeg7Ae798NrGMu+r2qbGYUqfzfLvFXFGYjJX
egAuA3xP/RHgPUaNtxSA0oIjYQC5swYkmZn73oBQfD9dqVD0Rj7ZXpVb169/
iTW3KvJxHqVHsQOiMRlvhbfbs2CUGD6xe2F7FXCHBJ2/RGgRs4q3018AW5OQ
gti1Mj17iCnS84aEw2XomTXX5IKFiZsfuPnppbmxTWy6OqSllDD6qgjx1or1
r99kAvjlFWRjVRlwvzQ/9AZqzlalyWUpmIs2Sh26PjvX/RXyPqxuUpW2UOqg
dFIx9RwZgu2rSbqRXWzYx4SkSjeLdBQ6ikMED2qYFYlaGUOWqB5AlmBg2FPE
HsIB3Zm2aAaIRDMfhb37K3tuUWaTuAdfWhYaVLqOnOkMlSgQk47XfHSeOBKW
PU9yTbe1s7+4pvD3IgUD1M3kQ6i0RdoLZPTZNKQL3nYN4XwIr2jbhgFr45P/
RfETJxQbJWDwLooM4FYIM+yHGx7daLiDqoEvctlJ5SG1roppHBTzdASITIJU
4cqpCAQwEpmKNAXQh5yt0brtOdFFaVdEY432bGE1d1H7Lae1bQBDEQZe7+VV
/1SuYJosszVOdbqTocm2OG5OfnNW7YGqtJfRbej60YLq+ADMLRxjrmwZlSRR
cXfbGTwzprIjLpaHO+2Od88W8e8JIyuWU6rfVbGb8l67Qv6MEdlYLh+jpeyl
czdX6QHElrTBYgbH7cUTcU4lKA64f1JugyqL8qNAYZwPyfqFyodHPp++feA4
/7dTq7TPKf/xFF6MpLKfUf7Yp1WCBhToxWTxO10gfm5vqCWRAxpvl+hTwAOi
shSxj1XWyYvnM1MajtmaaxRxkoY7QByUsqfOFtWvPwAlCjCjqftzueWnS2xP
PNvLZVXv75/b5tiMZHI8p9c238h7y+54Cot/v3VLVBkxgsUP7NzjUwspMs98
GuM0jm4Bn8qmqa7Xu/vR95CUXz6dB8zpeZZc5a3+NxM/cZxGJvtzaQwvNhyT
7Wbft6C1GX8ygCVsjiCJEZe2ejRAadxm/LIJAQvXSUE0Wz1nueY08ML3OjpH
mb5qSnCrM1wJzIF185KZovnxfNgZKKCpEEKimE1pC0aksS/wrnXFPdI1Meml
8FSmMtBwk3lH6w8MXpI6BINtCrOXfdkqTCxZOvbKJVNRbJc5UxAtl62O/fgn
meKsz7PDcyQzhtjA5BeKMSjjC+48u9KzLuM8Wbirx/unYKUypsJXMn0ES9WO
smsoUanI42FEqHICibN4+wP9BJcgJShtz626gAUOtIxq82akzRKoGAw7ztio
DnTAVq9Ul1D3NUqYjs9I1mPO5sLDVej5ujqvGpVUzXxBirQHH1NUruy6IDmZ
ZVek0QMghVdqF0fo0yqaSY4WfDXzGhgxd0z3Hm54Gtyv7dw4GGIFUHsqNXpy
cTLznZz1U+IUIHlcX2p90z+3wUMBPyeYXah3CNg0q2RRIpRgm/bpMq+pJPAi
+sXtvWpsYzZYwMr16KnNYun1CRH5mX0dF3CMCV+Va0qmWZ/R7fpcyVuv1oKv
eDI1f5NzR3NqmbDez+GNITadpHGY1qHdbOAzVfJFjIB/LEGDUwHPUjFKydBK
edi5ZXishzxPOMU1nKJGx+UWcSL1DsmboNTjGDtBAmizA1zpMlAB8Y17zhQ1
eSDxun8XZpy4C6O/NdCn2PGQisu7cXIL9UJYeIbYeMyfbt8g5s34BiOULTDL
GMNzuzSwdh4hGapmlI/Aa+lZQspVQeT4I1tzFElRhDRdynKycKReBJaUxmB8
aO/NfJWN5GZ4/PjyrBeW4JKgbLWzJtYxqZxIKS0M4rd9+hHJWNS/nwwDf9Mu
7ATObHbSYiTEYfdw0bHiIdsNQaKHgeEn3BznnLD06tUyV5FLAsuAnbyZ42y4
eQ7hUIZgub1qsvg3QJqNQ1NAe8rijbmRR6KMBu2210/M3Pwom0JlKjJuNYqv
bCN7GZbeNqoaLapqGVrQjX1+Ymks6xfpjPyoCIbEEOUeDvLcYW8faPxTJJAh
UZPrAEwYDILKKmJmFVQ6MVGzEFpwkVPQYr/Ide8DtwAGq+dct5RojfaKHMyh
rz754ivJf+xH0M7Bm1kHUKkDqDDhWSpxiAxpJwlRIU6lszP061lG5v7iZWVJ
goKCe5xmcEU0EegMlf5eaS8Djy5R4cVAqz02NTeXcO0GONmHXxITf7Xhk+kQ
H9lOC6kVHFBi9FA9dwlMJWeLfO9TVHdzRD1jLjTYvYehpZgTuSUpjvWLx1m1
NYE/P4AXu1yquqrLeMcPduQ1FJExYQItaJyEnFsQNA74BilR4K32s21zBHn4
adqjOMCorDMPBbjAzmHYzJDBCbLTSRhI3aN7zR606AW1FCIhk5nRhCb31wzP
zer2FG41+E69BsYkp6jEdqDE+uG20h624/Q1IDVrNeKGVLsa1fx1B/J5K6p3
0e9MJW5DTnjRtnR32llBlTAFqV97CKWIJ7hU7bVDgc2+NFQGNDTSetLe0kWi
fjfO8EgwRlhIA9QGomVrvQVBztFhr1FtmqiZKp+s7sc+PGM/E7NW15wTe0Fx
I7aU9Be9a7UPlLeKb5tY7KMU/HLu2vhurigAKYrUN6fIb5YYrh6WJ4uxOV0/
KkEXsmqOstl9qOd+93+ynPIf16ZgRWOLA23t12P8P9pQBgoGhFSCf8tBzGud
8Ca9H5s1OiZq99y5R33tFUcBe8lsLWQYGQKn2T78Ra18Ekiz6jcG1G7zzmZ7
vt+C9Hh6SxiOAGS1Ep5LgA2ISprk5Ji8H0e4FkfshskdhOixalcSkZHLmrp2
YVXu3P7LsfbCUELJ+CwKhYqV2k+h1OUp683ilEVcnLebWMnDTxdObjT4DaKb
to9TmaP79r7VRZIcuSchulmWEB06DQtk90jWfEoESXxmKb6yTokspvQq/XTw
uJ14hJlISTE0upQsGZY4KB0dOBzH938rjPlD98lmhoTDarYWlLO0F1pWzxVg
xbU8V9wPzkKBJhAGADjbbLM+1gLQMOCXnNzjnvpK83ygT09IJqpAFTwQrecH
Ihbbq8EVb26hteuhfr3lEY6sn8olOIeuBopD5WzSQgoM80/xyA55BvEyntZ1
lbw1QBHsDZoAFKA87ucgCF8E7nWNlEYAwUQDDcb2LZHX4qHpuFlCKhSa4MBO
1bB0TBxHmfGhPAaUrKvznPnPZyxMvWCR5uFr9osQ7Gz9r6kSyPXukHkC/rNV
1R4b2APi+krSHzr7seJ3oIOhYSxGd2o4cOWrCB53oIsp03T8F62V3gst2o+6
Pcl8KCVgChmRJPepNp+DBeZuM/RcVxOnzFdz4Mx/eFuHHqyaFV7WN6spuXS+
sErOuHYbPSUXrCumCRbikBs9vk4RrHRYqNWHT5a9smGtavHLgIzUFzPImedp
447u+T2Qe/amngnbUaf/Dx/eLomDkv3ZWqo+MMy8MmiVgnbe7mwDX6MMggNV
XimtVbN6lLIgznrLt0mn8RKEr/QeulTvjlw1TAbDElbiFIZb/ddeedsjCl05
vgwro9jqjd51ipcNJXP1hVLH++DDZdRI303vM9Yfjdz1kNc5BEncdAojiZX7
EhYvsvIoNp8LDJsscXLxnao5Jx9+nKfTyJwo47kR4KjQGlpusHNid9XoCsRf
wCm7eli+0SLOPtqLN/Br+r3TH/bC0aFWNtiKa6NCDMj2U5nIjo3VIfsnG0Ug
UTBWrBr0Sr7ySwP5u9qFLOCzUQJPrF22HWlnCsOnACmdRmiLr6Kpgheed56z
jJxSpjMhOxR9rdOlp4CZ0M/QyUa9Rvr4dh6lsu6gHqWtpYKOFqmKSSkrzEYj
d7PbWQ0D+3/nNt4kZbOFlsB/twok4tVr+kSzf7y4+mOfjD8WqfY+fq6Pgq7u
JsdgcB3gQLOf9kWHPWXhQ8BBvim3yCnuFogxdMZ/wsNcvJQsJ+BJiwY+oR/f
bnDhkzaAmFXY7y6sGwVqAguTZlmAZbtyVZKdngyx9oQZRQ/YMf8NPcBYUKfL
PZG+gATwq3tVZ8soddIV+ncUUfk0EqzP6td7IhGbOww3QesnZUWKsBUuZWv7
Nf2lR54A9PJ0ci1kQKmxlMigvKQepDWKKduBmAjCVGD1uuxxg8+zady0p2r9
/CYxTa/f5jpGgWs/drmr4M636mIM8JSGdgRzriBg2PC8Ic90TdE1EPOHbT7r
/yfvs7WEhwsKY3f6X8v/Dt04nBUGoJW6xpzTMdtLf/tER1vbVxFo4rka2b1o
3nmFYVE3iZe1JOdNI5J5YM0FwJmm9kJI8wATnR7lKl1Zq0IuULT6HBOpFBI/
LzXfXxNDw3uktOdpgun0GjUm+KJZ64WwNsTIdR5o83lsID/WDKvi5JsF5kK7
rp184odbSfYhyYi+Z6NxaiYtbl/zAsscRjhlY4/gg1zX8w+3R8P8HQ+GvZKM
er1oIombgFv93SteHp7zSoH6wG+OOue4RLAfhSFCQgkNPk7r18FWt22/4MGv
ka6OuaDuvAK2dKlM6MZIAnCRrRxRwB8qVhrgiX+/J7mp0S3NfmwQfR6J9v0n
R5CaMklf20Ez/CkoCq1blArrai7D8QjG3bNkufh3ZCmrCrRFae5eRfuSqilA
Mh94zy3PnRC+fCHX4/GFaHo6fLABiGwFBa0jJYIul95RDFgMgYNcK5DK9FYs
1qFoP4eF3ZAidAKdQ1aDTSwAE2Km7edQD9YomRzD2d4iHmY6qLtT+tLDACsn
VYRbURjLJUmzxBqPf+y+dYfFWiyk9niOMgFeRxjbgll6Dxt4ixdHQ8CeaNeL
HYAWv25OmapHZVbijg91RkaimMeMjsdAGWyNml3IJlJW5+ZNo+ekit7rBKOZ
y8f0l5zS7WPkegmyG9t44jTRAFVs1TgA/A1lpQ4uw7iVMIcaLT/WcQkTOr4k
P9MtKItUOQfPjFUwghWbR/2U/QP/lQa6ZVsfoRbAYWXKsmG91xptru2eTucp
5y6k+J42UkPI6IJinc+ccK6zpf99C/fqE+9Ai70I4IXBnDwUAUhFzUBuNJ+T
Bk5feu1ZWMdRIKn9kyjgBoz+TzZqRvIT4Viy0ENNOihW/IsBuSnW7ckgWcHs
dhnYEE9+miUWV2vJgIzQ+H1AOpWUGuVtRZXPdi//EZ67wdqI999LO8tkb0Nc
6VGIbRcCaM77EtCnbwBn0/g06hLW4TG59vVFjaP9j4oLZC3+WiqmnSR3mVLw
dWPfVbI2nVLSJ0P+cvaphFZjCIv2iNBOJwjOBgWE1OyBclHlx3n9gAJc3i2Z
VrAEgpqZGlFD5nXTmE5yYSoRctUB3mKFfqf/lfuwjZx6Hu6aoQt8skPQdw5L
n6rCCw6UzJFrb/V2S+KpasJvUdp+zq4dyr9dY1DDQQjHIIlU9jFHyfrGHcXY
hOctvN0FapKKbH9gJDw0IqW8eLXxgi2mA0arZbDtlK2qocLSFT3fFf74Tp8U
hiP+4EP3PuNN+2HJo12oT/uiR0eXq1e2/Zk0YRgYvzutTAtV+dKPD3RYtEbJ
SOAZ31/gDnfgMfZOOrluLrgiIggGNgF/KSMER4TDruIY/jS9m58LG0sOP0xz
XYBJKgeNVZBd/urVpNNYggmQo46d0saYwZu9XFL0Yd7R/fy6td9c82W9CWtt
MsGrQPiy9INPCs2rWVSJ5rlRBUfoJ4K3svVh6RMOBWPt9GfzEPKvpz6gfjCG
jBmQPoIAfO3CsvRmvCNFdwDxd+UEfu+mv9pytVekP50ZSI6v8aZYEa+rEsUx
YHt6jdG9jr5L/sZet0cKu8mqBe9RFBN3aVb6qWh2yOU8415+M1SRwaJ8SLZU
2ORl14iYxXr+Z2qwLZ/i/8NlTHiV4xCmMoXEwNYnSaJVkYN+BM9bq+10ltHr
U5bskJ0LlKicZpqfhsA3d82K8tSoarpFbvyCFwNYV38oK5d7B+mPEtSOwbyn
P2pIFF5i+yttlf5mpX/N2j1Jxo2O8wkWArOSSDupVE2aHF8DYt4g1/7Mk093
DCaK2mmbeONT2fbCk+QAfbTKXA05c3ucZQh7K5MGwyTmk1mD26mgdV9njez5
f3Esppw6AzzgGMPUmNpPAhX7zdXqo+eD89S1sCvzCEL+jaBMUhglAS7iahok
8s6PmH7q4Pjp7y2VZjUzhRcUIbNJpbLCxK3xpkTfb1PSy8jSSdgZkmdiyf2m
1McHuJm29JS+96XChbTiuYDAhTTRkR5mTfrdKgJpi3DxpT4GNDTTXDUGfP93
o458eUec9Fk7a71/lXR/OTJQ125kaWxzLbA9rWhO0cSTGhD5UK6UWPk/AGWH
14aFnZ9aNKH0zun5+AHdoBI3pxxgDeKfKLNLluiI4DMTRdRjcXILIMB4vEvS
lVThH2LUrRSbk5t1ixXgrJEjcN7wyI9jjSLuQ/sy5TzPFbyD7eziv3RLT5+R
bq3OaSAc/ERjTwZv0OL68beSVDrR1ROROjbxMr7cNwHJeMDMLIIyvla7gs9N
GtSWKGDPow2V8J8iJN4+N+sdmKymHKO06gxAKJuSjr5EJMRa/JNkENlGqzKm
//orW10Ghht8rX1db+9FkOP1rCkbR7spcvxnzQzblkQ0vL8YXD5DZWxEfaDC
wAZeO/daGG+svR/XE61rEMvxYwZ4jEGpwzcKkN7+kKBWdYrd5gDA/7uEesb7
+sHLHk8Te7hYWhHWJbIpvVZpWI02oitJBS1hg6CLsqnnzM2I5tJyJyD6McvM
TtNaDlSpCCeqRIFGSgkY90qQE5glC8D0EwTopxxdC4lW3inAaRkopFpR/SSQ
usV1IBLyI1Q/1Ws0jzu6tIdwnCjMAKQWKqv4GXKUE+OtXvykIzcdeh7S6rf0
SIoq0KiHka7Out0v1Do34n3O/b0G3pWmsCVTAJ9jAy64fcWw+cos3kjxZFp+
h3kRn3BYS/lmyhhbfkOocZskIXoyuPOk0Zns+vWf1TPavNpidcOLII5vnF1p
tnNhYYpoUaYQO9C1fUfHpPCJ8PVwql4Y5f6O2g0IVznes/U+lIViHlZKJapS
YJNcq+Avrkb0viw7TUmJ/7Iar2gFO+AyvcoyhCxiBTMUIftCzh1DA5Ydoo1M
jiKkB+eJRf3k/HEFFVolH8z3oHsIpvBtWNE0y3LIQR6nHvfB9m+ALK6as1m/
44mGYR67NxloRjW61BtUT+y9BlqP11BKcjR/3k5c2VIMVcMoWIoIC8HruefC
LazkCtCuoJV8Jdwv0QVZSpEdv9dLiOK1BUa8BhNqrtn2snS7gHcnbpSZMWkU
1BHpiq+25SrOWBfnFu6JIRGGAlgRjmL2vPy2b8tPDqGnCqb/Toe2G5wFDvfP
vLZFs45Wc+2t+ESu6+igbQm2iUQHWgfCt9J6WcoFtQAr+PhaQPoVAKkFwkP9
iM+Xo85SCzNnr9CWHz2ePMVVP7GYntkRoYL0h0NWMu4A1W+vWgY46fMoKsgw
3c5dIdb+6VVTYRj+m500xS/eH1J/vPsZYqABT0waD+14v+NcxmLCfPZvga/F
kTEtC8mgrNMwYvlIkwHJ/c4XCCTJpS04n2klq2A8HV0N3Ao/k6sJgSTE3dkJ
+UjyBBC++2bzlyta6W9SJc62eKEAzA3Yjnmc8/nV5nUALWSgNl3wqBlV2KNI
b2JPDLWRRKOxdlUXQm9pUHus2JYIdivwO6nhrvX+o6wy7F/eBoeSzSFZbxAC
GvRvmv6y1JDKkbUUZUDd+o++tf/o16/ppDQmzD0h/nCpgEW7pGwD4X2pHWPI
1Nu4Y1b62n0vFBQ69U7tWuAxrRcMDG0vdLeUv8L8N/nj7WUFcAJUWEMtNPKc
wTzbMBmoIMXcsncNVN+PEQ5+E3iy3yF5S+fITG/4u5AG9CSjFWGOO+m1Ikd1
6nwASz/Eb9clGGhWLZn29h1gwPsZjDLbx0JUQC7nXq4DewNAyH26t2UQWeFL
iQa2BIoZyJRutAoFFCS69fPoJVc7GWy4fj/I9hroIO2BFWgdEbOJ72AmjYGB
mOhaMde66REOQbOdrzJA73ucwUD1mcDe3Wk/1niFW6BWqFqSgY5RuKW02P1m
OWpYokJlXWo2qs314uaq1cy3RAdQiEJIo1m3KnvFBE8uVIMk6TphiHTeaolp
MARs3B0fPAQutN2GxVMKnPUXVQmP7wWFtotB620JwvKYmImpvm6w8vzuijpL
AxGtEHbZJomRsky+8xNuKhPckbioixhuBHMbWBM2Afm/j3Xs8OrI3blCkJfP
trg0UGDutI2rzC1p01X7qgsybx+4/Ld7eubqPRglHprWGQBuz9BkGjifwKTX
pNJEQzZ80K9EqJ2NzLYerFrnGJTEKEa7ucNNsSt+c+wza1eRpJRgc4UvCPUO
Gp7Ebvf20Q5Sp44h/vQiSYFVTHaI/CtC5Wz7Us51RnmWfp//CbAlocnWnU7F
APRa/KNUjJbKU7pd4o18Hnt1V3HkZZQFqxPNZ5JDitI9110HvUe64I/E6lhr
5sPe6jy/gbH2HPBClPylnDVZyJJTIgkx9XtsfwwJg/5GIwKizALWXbykTwPR
qx3wKk9VfDSx/2bJr8bZ/HIjl0VQFCX6Ku8cZESQF0aPZfaDDkFLj23f9pro
fNPTr7uXT66dRTV9ce851sU+ZkqIwRJu/ubn7gUibsiPLwJ+7K7RrOgQGlck
hbNWrWNCdczcPt6W/5ygcq1qabzDKwpRoTk30Fe2sxwnYL9jOngKAqNkbNGG
xZTadTR2WNDLe3JqALdKhJn3jzN4m+khJKSbmxWgjlfnl+epfV/B/cm+LII1
Ut8RgpSYC+FxA1Jt02tiCA2tMoav03dX/gaT+XdOZAGHMBUVoEansz4vv5zY
HYekyTlS4s/ne5v9cHIeItXIFR1gjNjuoSvNhfWy8fbQM7M4I5ctoECpSuwF
Y6c3MNuSgr3MUI0hDq5j6Qv46TiBcvi06n9DNER0OWvJQXFigHzIY7DcD/Kg
V8eV2JoaTHO77D9sn3CSt363E/202UQVsbqNZccAFLZEykyLwa/5clSstQNL
hFoNBIHxe06+c4T7IX0253NDX8FX/MAEwMKvi/3W5RhxGuUs0nOlVVO6aVPc
MSOVLCBcPC8CG1yoNawJSsJp0Y5hXWXNJTpwaVZPY13ogqGBL8GShoUYqI0U
P6JVGZ51sKlA+NcAgTKO/4t7DQDaISGmNpiNanKk+BSXhB/Excjg80RMdnED
cnZBKh98DurJoUPbO0Syx4oJBnsxyo2RRnch2dJwzhc70z1zMt1eah5PRA84
wSK80CXsFNJk7FnRJQ9sc+3PSO0g5e2b4ptXHZx3+KZfrj2X3k3l/Zmpq07R
AwSCaXPBrR6j3u+YpXtRQDMyzs9J1LrL7+wstiFs7Vjyb0UZVjcu+EEL2jPU
vsXN339Kmm8vpz3f76h8HZWZRnu6pWCIiirtt+hJVyTe6ZlSxDVJFAtA0wij
SpH7SKqyiqIzqS7zWKmaSfDdrYczKpEJJIdB7fBzfaN3C9fzYXUN9K3BLE1U
f0seYcJ/60Cl4O2qX1isj62f59WhK86qcDgUL76xNrqMj7sz1V5mRF9kpZLo
s8l1eGUYHvA2xYD7wa78G4d5UIBOosL0UqbGf3JQQhWMJvZ1xLFlFAx54ud7
LaPheMDBL8vcuq+8lkhdmgbLgvgNvV9NCNiUfNSoiQ8K7zap8OT8z0F7bsKL
NweQlzt1PTctHWd774+IoCJkPP4WT02c4Q+EKy9JU1lhzysmdXlo9YJJSntq
6cvlCw+SMMmDcL76IBWDTkixxEdrO2nq6bkMowxTszE9u8h+ozq8pZwBSFtE
jXwwoWypklJNJiR7FlHmS0+6F5J0B38opmodQcFihXUajHnziaic1zw9/7mc
bcvovrDMAtwdQi4lTEhjZjtdRCEDqdECQqRFG5gP+24Az4KfOUA73SJWOtvY
Mo0+dCCBPsELhDM3g1iEV4XA6mY1hzyt6pCZgQoFfw3nevHUkGdxdTXRpkM6
skANm7K8xXKFjv6QduxAvlqkVSFoNmh1fNxvg9yQX0MgUaCZy7UXoS9nLPMN
29Ws5HNuYTfS/I56pB+i8l6RM9zPAIqSHNJFzNsmuELNHFeA1tRLV+tHE45l
LQWFJLG8M2PWk1px7RBR6Y2+v6EVHHpCj3LoKOXGyAxXfzfEhkDn/zxMIqJG
6Lzs55p7HTir47FMg3XfUPCd00nR8E4uD2DrDeSxAqiGtqg/AHX6+aTtEpat
zAjVce/sFZRkoeaxLAbjZpMNFD9rVA50mR5ULXLPKx5vHwvMgCOphRcv+i41
aAJxLW+WoYKi2orJSkvP6p8WMoqpkccgi4k8OXpG6QJvwfyEMLujd9YWBlqF
YjB66AeFfjlasTn1t8mRLCq6f/tNCiN4fPMLzdZcYcLz0haayw6Ky5BdqMAZ
BkMYOWdqHuYRGfZQ2OIsbACHgkSjwlbHv6CLTde6+k+7hvMCfweUQkEEZTuy
Sem9ROzePdm95/pg5HsRBT8NpcP5fTqUQIAQn827myzeZW3Bu/yI8zPj2J/F
xYuW9qVbr8ny0xgtQD37KgYXsl1XQDB4VrNvn1IuBO+EcGSzh1/IhEidzyhh
VSaetEqv/edFiAGmiCBRhg19z07I7fRUIQDP/zcaRwOD0D0jo4nyQ49nF/Ir
1Afc6ADaKWXQMN5zzAypYTeDt8eK+jE5pQuKxpA2E/qXTGo9pioltKClitUk
jEMk2iF5vel4eiJazQ20S9kbK0IqjoiJJlkA/gQ22QGOSNAHlOADlCeFAEBH
JBf68kFKMJkOIuQl1ZAalcGWES0eAfhRWox1b1Ljbm+Unpai8B9U56jHjSbu
4SqrjPgiqHuiiXjf6ZQCH15nmXu3ZVfFMfA2HIH+kvsVyRX+sRA/krn8nygQ
40O7IFTGvxLZcopxJWlcX9ZuSZhl82QOLO8GaRQg43eS3VxSUyYMUULORvJN
RCiFGRR4nGK93Locl1Cbar3YYL+jUMw8rIjMFTKOhtUr6FFTzcukSGm4zMAq
MbTFUl16tOapi8uDVusMsBchXTlhOzqU8C1LZnoLrNRCUf2+WhSOB2F7yrxW
8iLCoh23DSsOE1gs57cLBYu1zS3K6Ohy/360nIE1ozUI0F779Z9m2pRJp1Hj
Y404ioB2Gy2Qq1Rd0T4azolTkA+T8AklObL4ekvoe4el+wfuvHP0GcQ1NQP/
tJiB6vyPKWfmgzJaERyC0AW14T/AVW+Xcrclc6FtLpIei2O8qKBSBqNoArEn
/G+DQnfI6iLcenpgQoFsd02bZnu4YKszRK84WiZudpgqYgEDlE5Ws3WVaY+Y
b4q3nfr++0KQhnf0WD8kNm2GkXqQhICoId2IER5YLUqypCIXTrLJoVH7RfVs
HwFZFcGxuIb16j1DK/rBgAYDIxMpsEnkhflsZvsKTeMGwAWfg4vqKWhDhpvC
jzTlKguLXwMbHg/slPCpCUM31MRVzoQyFKUBTCdZWAxESiQXUKSR3bZECv9V
WedTMt4+oqd2XwV9B6tz+upKxAODvTrsT7aai2ZfLtX4UZsiXO636qd+SkRS
NJzRRw+m3/MP/E88LPDpXx2YywBSl4AGIVEVnIVKuYD4lp4qF+1GadUZ/r0r
yLhP/4ZA5W0nvhm5Qgb1W/b2sCwnH79m48ZUf/nLF9YF13rq8jx4nmXaCu0n
901QqUUjCUNXX5MNoysfNPmvBURkDapDTQEGGpIgn7lUoijcCJXi7uLtFC1i
+CG4BKWua3BCYr0oOlHNNkhHpqXrI6dbCFIGPXTAKunQLv03KqWduRXxx1po
6jQtG5QYVVdGKWfWH7rTih/w6hJ6GjUGGATmaSeqt/PZlGNNof7A2kmAB2Yx
00fCt1Sbg52uRa0s+f5DsO1T0lMwYiyvdd9z+HnNs0ccOLyngmaI3rcTKwTR
RStRN//Cuk8oG012fLjCu+orYt5U5TVciXJEUEqK0emRpIsKn71H375VJWso
C075Gd2Mw5samK3esHlbSAK6Bwx9kaeasJXrSLqozv8ymzJwcaXtE7DqkbGd
usvWQ54uHD9SnKpllEv/L8PWyZItO7ZQkDkgUbIKUv5yvBcQBi7xnfQCEmHq
lJdBQvm78kmBKfb6SMKa2+n3t+JTQnwurcb54pZLjPHL1wqiA1ErtYKeIxSg
XRcmhUU2g3IjMxZZgq4iwuV5muNY98RRfrTwVKxJZ53+N8Qk/4G4N840JJ4k
9BTx4Nq49CVKRaaAMR0qN+OHQtxqMrhh+vmanXBLCuIl/ZzIifRzO2Mkm2EQ
eYw3DhqFuhaVcaHZanwldkqPUfagC9IGqKKMZ1wF99hN3Cki0ERJEiNrWZFh
N8sOu1k7qTDpnmmHyHoiBlJQYNCAtFVgKC+OKSrh2JrHkarmtq1tQQ1o9wpP
WlQiiwwyg/Txx51qzjbfaPsBThCel9p8tiWjaV/Yi8QgTt/p9srzckgjB7Dv
p26tFbQS7uCVT8OixpU2WRYU6MVIAjR5WLMkfr9/L56YeJlmvqasmIcZqK3c
xYK3rsWVCKQsVkGk3sxCopqWr4cYu9p/KSHoKdginqOqu2KIv6hvhqv5jXcF
JGcEF+ut/9OTgiOPCbr0hl6p7m++OyEuhZRo3RGs6cYh4N5Swhw1fLdnIDMI
TIzAS51i759lyqxm0XCta+GG1e+KyF1jh7sj5Vr1LJXUVb/3xEUyvKWWLFnW
LLyLHnhEmtZ0YNTUuKCnPB5Q+eRLuPhDMQM2kfFipgB+/FtnuHxlAKDy7zCh
JjcgpGgBOm8UZugVpIGBlNl3y7YZD9kc4aJWbL5KrR9evsuCuNHwGnU2Of8W
YNVl1F0G50Fzhg/xukNZ5wj7UjBVlZW9y00nUpOakllChvD1lnIKzSihs25N
sPquDJ2Vq1cvad0FnKUMtROHwppy/Jy/iHCHyBJD4zvTMGcz9x7yO6F9u/Wx
/QQtT0h1PXWjaZldclk8+Avb+3VrgQlDuRaAyyVTJBviePWczqcF2aW8yWFm
1W1r0o1AFyZ8GHXUsgn1yocF1m6MUg50z5fxVK9hTXcicrl1ZsDa558n7+1J
UPSGqyh45ZeuVmVvrXaVCiCB8k8GjknAOU3UbuJRW/dzdwQ0xAHlXZEGxWsT
CtyG4Lmw4OmVjWTnn1Y7OJRMprVwDVVCNUijfiY1Hj5PpOqtxNafW+FIPUsE
FnA3c26ELFDhALY9LNUFgaCtmladKTfyzQPPfF0a9gbSfCCZSaUPdAtu7qza
YiRMLF7VYAWRcAaoWqqfbqlUh9Z4W0Zo117PUIvAYzvL2pA3p3F7iTvlqRp+
p7VN+5/hgcFxtHT0MRmR8Y7vYyEuh1nIA4CFTjyzqIUYuSJHJSdXitHiApiX
XjfJjTH6JmtdpZ+sWGUoxwzRJ9z2W0y48a7W/wybyfvGy8d1woRXhF2C974h
jSRbSdSY+IxoRtgTeue1a+tBrjMu3l1XtYAyDi7CYOS6D2K7fIoDgnvO5ejZ
W3tsIJxYTRSI5+DH++Sxh62t/r+qjR3e5AkC6GVywDgl2Tm6inO5xyvavp3K
919geI/j2hU7Dzf6sP/CrAczn0SwxF/HYCe2Is/xZ8UuCpBtpgnC6kaBH793
YTGQEyW24UtS2XFSMP6y4bFGMSB/IPr9I6T5NH0/1/LUt1q2zxNmjsUBYgQ4
IBgpPB7blxFiBlUODlbi2KSH+OJurDeoAJTga8khzRY/MzKjT3DJF00mSEPm
5cmyTKfma8M85Uimv5DJfUw3g1rvj3t5v/wJHB75rImYGnw7DbDzngc4cd2Z
yl774oZDjFYCR3vrTvWIk8xoLjKNpJMOx1rbFofFaiE+jk2/j9NoGVBlz+XQ
b9TkrXYKFzbZFxQQusCi6pJ5FQYrZ7c/lj7pRCXAFLodpXNydlN1huo3KEwn
KPA9BTtYt6cH28P34PIy4AMGtgzwGtQcd38fRR760b2Uewx17XIgqgVM/sO9
cGhWldCC4XvDLTcSbQBgdt4+XONwKikV6VxeuvsJEKNaC1qWuSHe9isf/nv8
yCfRnJ12p8gDI23neH9yiOr//16NyVEPb7nK6r7CiUWteTvhod7p5TU8IqVp
ddzGTXwSHg5nKMM6J0r5L9Ydg4J1kHQE9+HL77hkND4ULJhBfTfi0eGej9xC
Cat1BuYIoAGfmB7lzYm2YhElmlWkWE5hFcwAzdgonH3Rq0xRrRBvsC3jWMGM
hppRB8+Cyox4qvGXKyu0++01w2V5toUyfBpYovQRfABFJKXheSfsRzujRP56
ly5fjCWwZDSiF9SF5hMzTlg8FZT8rWebhuGr3Zz3OgZx3XJuy4lifE7njIZO
mXaPMwGG5fwpxDN6Gknjfn05hrqSvxFBSDKPWsfrwWnWxQP/qvr2E+pv1yl1
iJB5y/MsmF3x/+OAanegS+UyTC7sqclMgSXdudenwyS1PLm98RN7C3g9NacX
Um1dPdp7gGWPd+KIuNTPtiE4AvolvfjVc6QA/RdsFkwk6sxuH/5kSnbf3JnU
wxzH2rkv3p2wLFXE5CZrCNsmhp06/hfmQVTJBJLgl4B0tLrxbeckEyY92kbR
w+dQEfRu5UyPt9CL7RCeMAFN0XNiOpEBli8RdLSsC6bESxZaamTiZiVlYZbs
7fewal0j+wTvx5VB/CFqkagR8iSIpEp8YdADX2P6M2yGkKx6k4IQb580W91U
REbVZynJOBtY4TG6sAXR+dFL/erMNZZweGMXhM/EYBxR3jEujKWBdLyAQmls
v2JBuF7RIIj/khrwfZu5rCuCnJqx/3dNhxTUx56AMsSKaNoCadZ7E+IEjQzy
HvfQ99Da3UOrh8C24jBkqJqukKuS8rgIodBjWrIwJ6MZQ/eps/oZkhqSmb5s
Tsz+cfyA0mVLqjtKM+CI6KBoHvP42OO2MJDWPLxNKP5wbnrJ83zrAzUa+Nv/
viuIjf6m9lo+SH2/mYUGnwPXR9DIPrrihFDT6E2z3EPLd17jrKHEqbt6jHMr
cuoLLBEyoIxXOXTyVmQrx5RKHBRMWM1XnsPGa2N0IpcNQsF3GhMZEBx+5xQ0
NCABA50f7h2mGTn7NJC3hSKgxzCxPhS4u8Lgmo8I/7Dk3/vkfaqz+a8kdbeu
on0YFVBvgA7+X6JMm6+pI/LqhlukFhA8w6POUK7lvEM4irP8o1KnT5wyX1fH
bjh9YQjL4cBYa8apmBfBb7mAfaU3+Uq3gZACxyFPAj+6RIrQDhTqxqmdYO8K
/AFMO3Tqp2weq6Gcr1fFZCvHql71GEKEPuqBUWhxuLLhExRD6W7pLL0iuCl2
CJ1H2wdVGqvBCxWF3IX9bWEb+uXud+rGNsX4sqK6oB0ac1EHaM58U2Ww/fII
rYr2vsF1x0zfRCS+5fJpmGxSZwC08QX8hBdw5htIqLQMhlBuW8UrTTi/kClq
HUfZ4cIk0hXoe9k6BsDvC+8ZpzC4NxJwrnJB5W19VvOflUzMtABrSp7H1T26
WP/fq4eRKiX0T/Ysc9cuFVvDywY9AAGfFkBx0od845Ixq4jkwWiZ17W71Sj+
O634dZT8ldIPfymCV9II7lOTtK7+7sL9V5KBZV5yR8MEKlPabe3Amnq/cPKZ
JCFr55+A3DrGvtmBNHv43vbGxC7v4rNP9JCg5aZWxZ37EmU8j3Lf721PeQuS
0cwFOlI3p6XnTXeMLgruL/lfreRYm4s60cB+xmHou9y4LQsio4ytrUGi6klB
vxk9aTF+9gXzzW9qaLam/zYd26B0qofagvkzT6wDWxOzdHr2KjhBXrXn6UF1
ULwyzvYS5K23kLaEAu0rY6LerJyMDlhhxNv3hDI/F80FTsacipkk7cS9q80F
X+0kqB6zuWhhIKs/BTTiRReWoai8ddQ2bnpR7YdTjxuXtnoIh1qEW7ogslM6
Q1fQRDgkqJu9D1LBQiTRYYRXssTUg1h6m4Cj/3Ss+hUbkgSfPT7oR92cOfN4
13Wtbi3KOOnLW3U/odOeetYVLQoJlDZFiW/dJHW3sr+tfBMOPxapgni5Senu
Kjo1n5P2hoXszEek0TZI2JVbQFE+pOnh20eXFVdDA9YwDmZODRQcg9aGXojq
O6FvalXG/CQ6s043w0rDmUKx7gK1Gl2SIO4tpgYRfXs66s5skpPnCHq5n6Y6
3ZvVxG+0Wai2vo4tsCaqKdgaWHl92diU/1Or9/OK50JcgnQbidhCB2JfnSOC
0QDbn94W5vQjJqWxl0nuCdyHFGgshxpU/FF4yhBDKhxjYYAo/fTLQNMWl+kd
VlmiTqjEz42bRkHGknTofZ5rjoDuahzW1nwqhKJV/sn0rrv7/oRKD8Piw6vf
pAoELcZN4OOMcgA4EsFnlfK1LZaX/xPTUlvhY8F2OVYxeCn3IayUB3815vwp
8t3ohDzJeoYjoCgUpv5KATa9984UoWnyHPfZ43cD8qmvyyjBYeBwIgKyz9yr
4TF/U3as61/kMT9wy8hyr7NqsbwC0tXE0xSDQKdT2D+j+ov0J1rMCibwnlDd
Pf1AhIA2erCw3vc9lroGBlpa4FDe11ZhOVlk741WJ0gft5PJc70hMji4z9a1
8EDieojwmHMMj3cfjs/5nWwkEy49kghsb+2jMsrcI5g+m1moCLgRpawbZWGZ
yT+dyiT3uTrP0XZcWBHKDA4QtEgnaDxd6jmzcP+Dy5FwdP+DVz4zmdWzM8hL
opJthnHoL6QI7qzoL2ZM/Ga+o8+nHaAd+3ThcIMymdpnxxqYqF12OmTz+b1e
qYmvzxt0+8cRrXhI2u5W/ripK3hE7BBl6anQk9ATzx4FBqPqF4mHga4mql+O
Hu0EqrUD6wgbpoyJ9MMeCdgUgkGrd8dvEeDVVZQAuKQaAgsOteLxjqyoXftG
aypnbvVX/Tl34avrGgSA9Ha6EpAnV+9PO6X2IuZ6M3gZJtBVW73F1oAlFfOK
06t+w3uSpXptFZRFotqKaX6D0qCy8gWOr0t9CO0AFSuvaZTqivbJ6+Ug04AO
7DOcveTLpcNfHppMf+kAvobW8i63B4cJV53gApslhgTcdLztUOu67C8fGefT
2YN0NFgpaYxIHUHfoj3F/hReB7+qn8bofMntU1Ru1UUMYql9B3hnuDKoNgor
e4SIp/UXYXOBRvYrFF57Mxfhi7H9EizWcI+sc9AQOqJv020m80U/CxRTClCw
UKXu1gkybpytRGaMloWdzS+H5+rpXq1OET0wqi8vTKzgGO/MWzto5Mr+BmoP
a/ONE6USpcxkGCvXNf08nNVbGUrBWxYfSi/0lv2W4kk1eiXSSHuiZJb3CHfM
iNEDgnBREpXGPvSp3S5xRKoE6VeWHQc1BYU6Uq9kAEvIwu8yZdFAaYvxJM59
WQh3s1gqT2lxlZCIB5t7H4b07Z3i+4gTQsNFAz6q9JGpwSExJdplCE1cjkqV
5XqKE4VhIYX/L3bIWdKdqv3YppH8kq5m5aquV1scJynLZXH3F7qRihGNR7xK
VGZA06ofT8ePDF90QO+4cR/MbXUuBcFsvTaMCILAET3Gd5TJH8snlRjvdOX4
7CSaaeyRkotRm1UMIaHmlIrW0FDo4RwF1MHzBP4/kjj3y5XQBedwqvvMFH8q
ToqeYzV+2oeWI2EzpRofMRaeo79nQ9lrBzIiw+Qok/JwEOFhUTZ1sqMqC7e5
sBG/r+roF5fVkonDT7GtjxMl7UXUdAnCqhtHfWqDgRfNdNd3UHjAcUvcx0g+
4Va015niNC+V2eY1/FwTrmyCnha9Mu2I7FFrJaNAjC5e1xXQYSkyEoZGUU+H
J1UbXANT5FN7ZbkEVuXhjrzqVm9mSMSOe+yG6k6sNbJgn5qA2FotMcev1Rxc
I7Xn8DSBM9UaKbYsbnFVgxkWhrFSUvvxxEGLf+hcICY/32hYp3750twpauw2
PFReGCXDm5DCIdrYUtz/7asMGngXzOb+COGkO+HG6PYSMoJkW35I2lxD16kV
mxmXpLuBisHcHG1y+mhxqSzcVzIe6Hk+BOchgZJbHBKHqbkBGOLP4gUgB06R
jmSKFADuS7d1VB/rLM7SpFAEZ0mzw9CahYw9bFwl7V+H0t1URrSMCB7iefPX
FC2aWdxH5mt2Csf+x2tvkFSnH8m9z6SrNpKU6QGSu+012IPwXvk+Tc9NPKAn
Sgzs+DdO2EG9Ad0kGPI/TZ+X5XtXU0PXntVoyp0bU5kTndaIfNAPf/73aQLd
nBJ9AnXJrG+wz0oMy7Ts38kVnzC1RAmfjWiQ6d+oJfVqPgT9P7QPaF0F9bPP
YIuBOuXCNGJMj6MlIw2KAwwV1w+ftXVqqjDuTGfvaHgIsuRT+DVHMnFKF6BC
dgchPE+/ANXK1JQAngFXSZUGyee0YftQeNF0emPNxGFiEiBu4KfO40QNg/iU
MFhEp1ZglC9mDmFk9ryt9/J8eNg3YkqfYSzZLbo/oLBZPu5bbn2NPhK8cWCl
oPpfKjIWBEfnatT1LUhv4Ydd71JZ2cFEZ/RBSVP9XIVPB9kvkZN4ToaljL2D
LP0mAZDSp30cCTFmaU7sW/SxY+x8eehVXHh+QKH/tn4rZg4S210qQOERpLt1
3vt/jkkdaE0hbCJ2ewihnna1P5Z/p8vi4+V+5+zAhBBXmX4OD5FNsIUdD6EP
YddDbUJ7x48CG/6L+dcK+tRoicwPHo1AJm35X6tW/oM6NOeLc4c14W0Y8Bgv
1T8QcrweRboHWPCpTnYuYB5bH+tUrfMHYh7MHe0FNZ9DgWjcLRglit6Uz0S5
KLSE/3o7QGMx9JcYq2chMYV3txTPJSmgysmAp0uBvHpShKfR9PiPdLWhDc1M
fZz7XyHPYKo7RVv4495OxzLwjkqgtAOO3RPJ3aa0n5VnzlNVLJCInvpqPjTv
I1vhWAGI/NbOG6BnZbLxX2KTi6mt0IdhojJufTXhapjpJkdETFwR5LtmszhQ
j+QV4JcLDTGlwJMpwngY9gTF8mpqxU/T8JEjn09X/J80tu1fky5ZzG5qzfCa
ZAR1bshTRUWfHooYzotGjIWuUxKjGiXIRcf+/3rwHBp2vl2+dgXAVbdHuWrO
2BE0+z6oN5cFOAwT0j3JcKPTmArmPw7p8oD/zOCydxfK+jWet/Aod7esXtvx
FW6+hKuQzcgkf/Y64E6pit8hkJBGPEIwexqq2gYxrl4QlEs8wI3/W2qD4Oa7
9cfRjejLDKPJORMD5ylzp4On75utybW7omp2uvHye12OOAT92h0yRp8OU+IQ
pvOA3uvHFEevaGZzw5YAtZAL+R3Y5E2hPIeTIAxaxbpYSwtEgG+7HyT1sHRu
JRmQUiIuSyWmrJfnTIdQN/TaDFE8qSZvdaimIRTaDFf+TUhDssC8kDiT/EBk
l1bs8kOryXfc17x6Tc9s1wV6OH2mMPcNFhtZc7zSiFSLCTwS5xwj0G9REhUo
G8hwNFnmu2Gy/AE5yGZiY4sVUnVGlaNkHHMlfxasoT+QvFXf52RuR2hwCve4
YfSkBVjyYe12R8812IABM4Nga4Fe5F3xAk96E+yY+8Nf+0BW12RONayMcNO+
c91J6FIlKDXpWgMC8agZW4j2Ph0dszFyoR/AlYNWPQ1aVQCO/EiqBnuXKgF0
lDA6AgXj2KOMmq7PE+vDiqVgdzx/wi7UY766oH0PZvBMr7GKcNCS5932pLum
L+IEozRJVgnjZVCGEsZeSzOpwAgvWOsMveaFnE2v+7BK6wXQHhioCP78SaGv
PYdsovSIOD7MqIt/0y+UnTratfaCfWjiYOfmoIyLf02xb7TUfVnplBJLgHB6
NBR54Cgly91adG9PR6Iq47qWl/13sdd3LxUa7wtU9NBW5OeaSyyW0cRmBWou
ZFZuWzt8Se0eqCcqz5WVB8RPGvrGiq3Qr8UsexC3Q07VnVQZOcaJh7C8B96W
TvGrh5F3SgVJuPlVGx1YbQfUDj9KBckeHEjkZYp8ApiOH+rCQsL3C00LAOwy
gAxsYawbq8Z4EPz9v/oxlo2GuBCDfUvQy87FZZ49WZd8QoNQvHPY0YCGmXv1
eTGF7iayzVomwC3QKarM15Zskla3XzSLwt4dPyzes2yTxzJhXl9ohs4dST1e
zr44dhEH64eiFnPlR1W+4ouBYsFC9USbJP7ahlPAXQ7JuoEg9GDWN1R98OlW
X4baykBlbzchacvWRIG/8YkY2KbDXjcdGRe6hNuTHxCyjdhzxr7XTTD/91YX
8mNHm5EhsOwg2K5JsemSsUama3glzFL+mmnCn5vj9Cc/uAqg8U6f+npZKVo+
0ReakWRAPpETlECDdGH75raVjQBe25SZeJqOPgz/QG9vS7WBk1vkO+Mo/ngS
A81tIyy95CSUYJKi79HXpmsJdUMMrCorlS1vfwu2lvW0FnxR8+OYW0GE2rIE
eF+vde+q06r5acMIIsQmWgc6StakzDkirwMegFtwAMVmZkIDetK4CeiA7w2H
0JIDrM0YkW9hZNSkSds05mpnVuMCsVIdPtdb/j9i+N6nroDvcfwu/NyI98w3
+DgRIZHNXs985/eEW0akzsr6D/VVW/an8Q22qzdj8TSzt5+IByd1bR4zdW+r
lyDcjb3oyqwoHsZtuvNShQD1MkZ4Zr7GlwU1BkSldmqCwo6/iKiut0IJ881g
sUCYl+2ACA2WHkyeH37wvkyrKYQrTgb7iOaSCwqazqFlUW9uILroFwJmLqDU
bCCrEh6iAJnR3saiLb8RWjbHrd51/pNpLInX6fDzF6eeBBtqK3NOiOZmFSMF
1SaB+Irf3PY5qws3PVKysJQekHigjTB91Wq0mYk7jC2x1nPm7U+TfBV3C8z6
FAfuyWqePB3ye3EGIze2FOJclzRHCNBXJnuYFHFYcFUdTeK0wX3UqLN4BeC2
crWqfMO4ghSAG196D2QfSW0JeFOSFZ5tr2Bw6OKOQwpUbZJglfUc+rxwEQzo
0hsDA8xJOAmTqetUE0smfR9UvGp3E1n+kRzCdUl0CgfDkPXVhJ1T0BsAIsY9
5gzxQW4Y4odFl1KWELyyzr6JZxAKozZJp4VUKeGVDnijhOGH+0X4Gq7/wJz0
DtO8tC/8psgMkr13pQnZLQUrXXU/uppHZY7utRWucvg6qCuTClikd8+jzEh7
OKUuc9I851rAdELj/C4wGd8MfUy9rm8D87TfDBWKxEFRzxWWh8YfV4rYvaa9
YeiEpTjJxovBLdgo5rieieVsSp8jY6V+X9ktphJvCDzxiGCekiAFZFOlnNg5
AiqZNkjRq1ADieLukMdcsCcf9+Osofmck94N2zIKTyyI4HgfWtFRWz5tzLXt
ix+3XlPOiQOrQ7QLkG5Ap1zkVRxQV+msDebkTGXKjXe2uuMMmOb7uxBOuCSR
bOAWiHjQbYMOPClu+MGjea4fjt2G7D9kJguyEcTW+yAylIxIoK6nUb4XB6Vw
52iAnxwlcFwVoeX1WNiZqX258zcQlz0kQCVJFsjErSQs3dGECd93Vo3nKLKh
RN0NrMTJGUsqLMIP78gF0K24zdhMSAKwLxYCeq+aqciqpGSFVI80TiecPvob
Hhqi4lyPeaRdXW4jgsi6Om90Rktgs79Dc5suaJVViPbB/kZYzN/R74nJbJu/
E1LBu3lW7vorlleIfTeMB1LNB1beEUgj0QbARs2STvyTbzMn/lYlMGsYXr70
e/y/VI5PH5U0KhAqWMt7d/1C3ieN6nnSAC2ftuJuyadZvQsZstZJP0hF4cIT
F+V8/lN7HKA9iRVIjOsOPj2ky6McX55vAOd6W3I6RxeJgVQsk/nPKdLexjkM
5GdwGsr2ti/SdhvMb0RpSZoTqATlDL+3vsRdpyQG6/XkhSi2ZIAC+6+ww5TV
2+wqJ7iUmgfEcHDBTRch50T1i/0AW85nIo3dBkb+ArPk55QqPxSu8Mv1sEOS
gnexMG7cMiJjd1qt1sCxqVbjxpvdVnGA6qEblkoo2SFttu2y3rYubD7aKOpX
8/+//etTn1F+hBVzJche8/mQF5G8JaEVMWhRxxrC/QohuyMGtgqdYS38+pyx
elPqs8w9UiSwlt2q74vpqB4nXxtoenv4v7xFKva4qMJtZ7Odm+rZK6bUxGI7
FJUYU8h+aEhODQjsD7XBVsRnHts+EcMdIMcqaql3nK146pxtsv+104eSq/pq
bGu+c8xACUnFDXc0qS1woBcce4UBGael+BB3wS/jjCZouNQkmZakvrxWSq1c
BTb1y5U7iT2WzLvyqWYnVHMw6Fd8T+0yS4Zn4FXcxlXtpQ4LsSrIBi0lDwnm
83bq8CG+/k7obVdBUZSfzNmEEhu4KHX9Jz28zlLfBkM0Ci6OL/7392/KU8RN
mFIGBl5fmwkv2SC6fw2LRRcjobNc8GBsVmUUAPz3x5Dw9iXl8uGfpVq8yMO9
bceYQ5byAPWlDa6XCl0hLj439qJYEyQfYms9bRc925qJWTXLAjmxKRSK4Tcz
XxtF3uNWzwfflgS+FzhOEp7vKxWE7R5jGNFyvFdbBMx9Dyk4NteT0eEpZzGS
VszVKOUeuLwdF18HZJRNlCnuu6j9JtmatPI5OJnl+f3mN2R8Uz+4UfoN5ldS
WDq8A+Kn/Yk0172EqQ1Kf1oNoVgMnTHAy43+X4+n99I7Eel2PDZqedtG4dHB
7n3IwQI/QEAGgBzuiVTW8RbA0iRxEZPkoEGbmE3VNQLxX3gEx4E6jSCkFk7i
fQW5YK6buQvH0FHeGbAbk9vW1lTL3PfS/v4IHY6ne9P2cJXUhNxzOuesDvEt
St0+gzWt8Q+JApY3+iT78RHtHyy+n/XoW59Vn6SSZOBT12WJp8G78eHF/g8k
FkFhDVPm0YzgUFkA5ZfbDIwCDVXC07Hyt3S/MAEOav48zoCi2CNnWrwb3BC8
bgaxW895sea+Zq2RPRSY0FV4yvJuWwEPwnlS21jcsPBblParL7TSsI0O7jTD
huSn9uxc1V44225irsg1iUy0SvY+gwHE+yoSveqNTL5lwtjY/ygcab3T7Xc5
oaLkHbJWlO9AWDh9pNMgayVlZvbEObGuCIw5QUBOF0HWd2ZqBWRz33SWPY20
lQPqTX7f8CAxdJdoZPDn4dIGOxYH05jBY55m01n+W7Cp938+pfZ2abQdM2BP
ZWIEh0zSHladYRx7HnlGAOlHpQ44ROYAjP8i2kujf1DnlJg/N5WdMETHJrG1
TA1qrRWy1hFSB/EqRLZlzEmczGm4jktUVIOqFN0yXGGDkB46fITeeMgo0sWm
N/HtvSv+GG0zLhEv1B7sxYKdVmKgRfnrg06+kQp6iWLwPQkDO7tQPxiAjJ3w
K+SVK07xyJgWVuHFcWoH6T2RPmCovFkbn+neEqttD5MLda12lojN6I3EWgx5
AEqwWZAIgkBijyS06vumfbhDUO2Mm4kGWZ/DpM0XN59TGle2BidGIJns047q
lX+halB2ETzc4grpS+t8I6QGQhIBvzoaf8ORXZ5ePaiaZHuXjJ7o8Tufw/sM
/aqbgO/Y5Mbr7vVbb6VjlBH5tdTLSQSGDbMqCX2uVNXPzov4RKBEPwRgWZmQ
JDnXjhuQhl3f+Np/9J/f4U6fOHcw6y08smnxfGlIE2lJF7WD+Tqe9NqsTtit
ajH1owse9pgnkJSRZeqBMwzJd/VV6U3QIo9/wfX7D6O+z9A3gnaNxSGBqzoX
ULa+L80TcP6H3tv6NkDTrBo52wXhW26GV6qHskbUL8ND7ptzbUaASzemWvY7
eTa8qIXbuSVBJ2JkTyOGVDMFhxi1Uer4PnKc95wO9vVEHIiAVBEaMmRmAu1m
e0Psj1IZ22uSyYMBuG2s0mZwkj+TrenpwV6ECXjhDqlu9etHtaVLnAQmcb/S
DeWnyqAnhL8GJ7ZawVw9boWN32FtodT7iCra/6nQ831U3fPbTWH98ZpBKbQ3
ZRhmCWvlWvl+rmUJoZofPeFkBIY1W/WSHhv3mlSjBBy+qAvdGSSp3tUmtWdf
sdomDNCeMRfLSwi7/2M1DrLBRe2fLjj5O16+bBJrgw6K2TSvddHdrMx10+At
Y21ReMXuhq7yLAfWixXC3LqVW9MAx+70XVdIi2TGpJ8r4JddXSiYgaj0qz5o
Flrn8PZTAEjQSlUV3LLS6ILplWYco5knZpWSB5ZjzMDMXXvTMshHe6RGfmj+
aH4oA9RZigZHVupkX6rJ4kqLS+nDxjzEKSF8CpvZY3FBFeKjY/BzAXadZ0R4
ByBGHSMkVPCDE3OjSsGlQ6AKPDJ8bG1NjBgWV4hyFvyCokhA/GI1vhHZS0Uw
mOYMH4Fveg2Py2ACTihhVVTOJDc874mO9XT7SnHZwjTtSwLqpHLv60nAe/pJ
lb7KL2XEMq93l63mWV5WVlx7Eb1lI+x+msMbLDKPI/B+MokqQUCMxFxQo10k
l+hDDmwRHzJw1EnWiNF+8PcNsFjjkyjBEZ6JiqRjFRZeHslqegNw9luBZirV
vUS/p6jNbAMsYpQrSnTBoLumZfO0AyaZINcnyfTXhPcRfTROrnb9Sgwq0Dol
lBS164mqrkHu8x8fKzYxySnMncEuDKqgBHFjjP2ARYl61Xa0PUXntQ8lhXae
0a3GBaRnjCac1ifRf/8/yuVTlLpgxxB4TpolRAzdQMbINKFUOgD/VLL0lixS
EnT145Hkjwo0jqWZ0mZ6kzroFRIMmGqJx2O8II8HIGCjy1c57Z7ElVOZvotd
elePqGmDiws7PxworvkOLqpZqeguqs/Ky00BAnStgj0dFYK/+k4R8JhHJeiC
0+v+Pe0fCIiY7VYSBqYbo+3MFfqPgmqyJWe8Ukzi2Gsfdve2I5SRSR8EL5Ge
7Zf2cNOObnOr8L7fxavtycF/gb2PLKIw+BJnuPaEah0SJ0HwgFx9evkPXcIo
h1Hz95rqqi96iXoJA9i9AFP3IzJkLlSNVXbNsUDmhbEtWNioIABujLC4cRgv
cxJhCPJKYIN+gkoKvNJ2kiadkNWUP7Wn2XVSfsI0VgRJBpBhkigycka6Kbcb
VXYJPE5+cPBUn0i4MpTs9S6QeR4WQdXoCsXyNtCbrEjO2HyXFPYIEnZlegky
sartgxSdOW5Rf6IYvTDaaxw0ApDAJfwFbXvdyTSSG0382Xi6t/xaaqIX8Amb
thSNUZyGZi8O6NP/U7TBrHUA7AnDjU2J2/jSDE2U6M86eawGS379Wm8op2fv
6KB+MqHmn36dE8qVuMsNMOr29pnp4qXGY0YXq+Bf734Ykq7Qk5nBbb2Ygd0v
febAWbzASL7CLXw9ff6xHCt3EzPMT4r0ifnk+pMFPrXTll2QtMMtNdfNdakp
L/qFMgBSD6Zh32BBh6S415La5zG0W8cjkdY/2DKx8Z+0Qg9XL3DPUeypkHPk
NZdObtQw52B5T/XdKNtHdda5LuNI5MYLdW6j1b/wljERwd7LFZHjnhkvYX+W
6cv9zyHg8LK90/lIwMC6REEhXgpy0Mhb81ZZNP8Twq1BC+HAY7GBRCVHOc0a
ZCBvmLj9PJ7Pa35/2oRSFxxTZ7vMSkk9FAGFhEDxBi2FXa+T8cUgDI+7q7sl
t4N10N6Q0o+Q4i3DJuDeVyihnPbPB5w8AJEIalAfhvxI3ee+x+hsYD60i2DD
u/Yd0/f4849kpas3b/83FvYMCR0JHaKLAAaMGZNp+uo2tRjYAw6DW01deOMY
TWiwOrSu99MgUWmtQafBDReisV4DlozXhvZjCCa+spnHUcmUTzExDHM/E0rJ
FLZmoSx7bHRhl8rDW1yRUsTM6yJdoJO3z1jMPRUJrxuqlnjGCNzEdq5SehVo
eoLTyFOPD69CQoYhZqfjFS0lxxobqgFBrLBnCyXBpraOMABx9NPupiRgL7Pj
9qPu6xK4WGot+t/l1DuF1BxdWE6RNHnyDiXzCtwPQrO17lVqELdVVc4/2/Nn
X5mJgHz2jsSphxkkOkVV8LDokSeYNQz2Ubu9kby9yPrO7IPSVnZR9057hBVv
EZEf/HpXhqf1tFq24UTadzxm7+e11ptfc8egd/irt+5i7EwwEN4lU2+rZp1l
awVQ1SHOCm/DETj58k4lk2Tl6ZtyDK0NnvNR62V8QGdAxDe7uQdXbjtjZsRH
Edu2fRQiNnlNQmoD+/HqqjP2sk/SBKmmito629jKXQK7dNOmGsEWNmMuFfTf
0PxlmuWAeoJNQGvX2X0KUa63AAhpdXoG18Ki4bza2W4Z6LMkgYIgiHCjerKw
sWwfSciaZQur1/6PU7ho5pDgWlS+h764+HovAQqfvs3ObVd38DkNFP1SL/kg
ZMKl8Ew2GjxN+igsXGm/54b8dDg1GOd6wgYwx8aY+xn0qrN5yKFdgQrC8ffl
cIk4r9iQfvMiZjHdZmcEqKvJjLI4L2BOrYd6xRrKAvIBUx2EB8KXjDjZ5cQx
p2WkWrYuWlU4Bj3sYkQ0ZkcU1S2FISzMJQKS73a7ssNiG9qajig7jMXtJn6g
Fq/wvPemDw54yzwBLhNP+icqo8O7etoVMpAaVwZRLHs4loipcUDvIW3WGxlY
qbbEiNhiNvV/bu4xTcn2A0B/VXOjCIzj0+f3gSTQkNhOFC8kIE+NI4QKprlr
qqL7yZUUMtJqToJkSSw9Vaxw1+JogZelMIqEqreOm6G5+bZX/jVDP4Bb5+u2
bodWZEAtgSpmPYg3g+H5eGMeWBIAyhu8isJQEV9EHcTFr2vlv1lEvFHq2OhJ
dPv5/IdF9C1IL/Oa+Xfh93ZQlIAivaV6tAk/eY55sudkIhGaRnmREMbQDJr0
NYssOj02nYtDDqgLHBkDTCp6X7vhaA0WmjWeOY4kV9Um46AlawY5LYNdszrZ
OHXILwTe6KKk0IeCwn7aKhLpYNU0GE9i6hBcH9rRbe382rQEXe9Z+MDxhKkr
pnur4MuVaDKq7oPMDGbh19ytjgPqiyacChGmpca3jTakgFNUlSqY2AXshd1R
UZDm7zK3EseKjVPFMct4OCF3ucZVy1WGfoHghNXBWdN0BUEUtYLmuN2a25hW
VJnlMmhDPUpnUQHU5ZsbQGhIfC83Ri2UsDCqkjhPZQVcMCKl+qLhkRVaHQ5/
op97h0u8WB4vaIOmAqibGUTlqTCG4t4mjZHE9m50OzJBhtdFPxJWiHx4v3gD
hGpb5DaC7jL7ljpahFspp3ShCPsW+0fuPaEA92o1vw3pE3/k52yRwr95TOtU
H1c96TsQrIGM2wjrPDkGJdgG2E4v70xkmTWOtCZS02AaNiSrtzC+DF6Jc7tP
lvYeLkYbv1aJtY2imjMrLcYLEq+dzoLY/o4ANsXze9S30Ks2jVxDMTqdeI7w
W2JItcDITSeTwRWAxNxbQIvtXURO8VmjyZOWnwyLMLJv/XNIIyT+mWvhSOD/
ba9Zqa1kIbr9LqHbhsPlogmIW8VR43CzD/MpDw+D0+mkxsR9+d2grmjkl3wE
fanqowRdkY6hRB3Yk0/IAUMZZXKsaYH5tJzJLVog8+b6qI/hb59xhH+1NYBQ
tbykCIwJ10FrBHAsTcHwVDBQ0O5xtUmFCUUeBEu4p3CrAJwMH1pqmhc3zhU4
fT9g3+oMsvArc+8PWwR/e512GI7qPMJvackeUAhiSO8rMxEN4Shuu+txZQwg
B5t/mdMxqdeqtrOwnp6aWpHTeAKPOp4IvrRf2ls1S3JDdbfrWhAUJBjfVER3
4W9ROBQ26kPnDo/14rsM8mFvfNHgFleht5q9rkGkIBLO2upfA1DH+k1LHf4R
ur8Et5C9Co/T/tbsnpLXhSHYFdgTql1t8AY3YDCNnk8azvIMvW/0faqtDXjX
w9wpyzWZm18EyB9sMPz8cnY9eXt9OkwkPoEIH9nUGdcXh4HuVNi3mYo8OzfV
M5WZeJcd/Yryi/QQ3K+lJnKbJS9KIYAGSBGjZevtnSGmAQ6sB123hwENNrPE
3Y9M/YchVsF5KO1QlJH3ybEiAdvyh7rHex7zClWnSiGa3UVDgt7QSYmRRYkT
sB969+8/XFgXkT+dahEz2Wdju7PXSt4PBmx6B2eUuWXXQWIarXMQAB+aOOWz
02UizJSwhe8IfBLoeBn++E9HKhY2sRyCxZN247jLABGFNXwDu72CQ64zrvaa
m8X6DJAqAAv/dzScm+YJzvmLuZBTE+lpizFdqZMmZz6Ia2bqTD3DSoJWlIdJ
KqyAlsIfFQ70eSMd+OZ8j9IzNTov65aHBogRy72NPuRkXHgkQsnWI7jzdVqE
+pDczWVnhMSeJ2rqc/Jg/wzT1C1jca3elZQh8FanQntO4M7StuQU9p4Ho8a7
47X4NWbUdvy7R4xUKTOlYX8sjDLTD06FG1VprvfwgD6kxWS0VyCigijpjZiG
FEKxTAP5eq8ENvrahY6mte9Hw9DT76hgcT1HnMIJTe8TEdW3+Xe1XHbkHtHg
jvCattfnrlMOgz03UntoFdkZeNaDig5+aXbxMDNqU6hjA7SLOIzU13V6Yrgw
84PfjCxaWEXo8QqOgw+TpcD5tudnqL4xENKWytk6uCCRCX5HfLWPdOhtA63f
fs7ywrcoB1HPcNYHX+KeOugFB5K2yRFTOsuoBAWHI/vquHsNAgcJoxtbUpi6
SyYB/GAQqDJMXi9aUZYCbtWaXjMt6/h5+EdJH5YT8IeQBkZpQMHDtTI796bY
d/8D6kEtdRdKxExsoX1Vus7hIaoqxCEtdYIQuGJTHPvzXk9kdrxssqVq64b4
K0tuCoweVGKUTaHm43r/TFj0yoIzccNNniXRpxXlf+FbyYwcJad3dkLEbL3H
DZ32sF+PM2xQeeJPXSyYIxwqWxvVRnxr2Deh2Lc94A9fwQfw9p+xM/Cd73fA
KIwt161jfo9S5G0L/kCgA/X+fRDPKpPl2CFuT3S5CAl4TMX5IINH9Jpz5ZYA
qH0BYXD0DyrcaOTasN9IqRFciRnWwaMTeLaoC8Bm2QThFnL1W+7QPR/NubJx
JMnd6Wo4y3TpYbbdHErE36TadQpVPLNLYkvsvEczqTqLyhFS2TNfMhg974hV
pv3VUeSNMAN1k2o1MpbHRTHI9BTFq7JtWEsxvedVGY3LYe3DUZuOmiYkuptF
dZiDR/PUkZtYI4p9eJgIsuSUmcr4Q5PNdmdMFsJgk45Whxkx6WqGfdvy6aQQ
7AyttC4tusXBW3mzwMuZ6ALNdwt7eQx42JegyOondoKKjN9pcZ/MShSmqDGZ
SAR+3RX0AdDi608MopuPhHY7NXpe3SH4Xwd3dxOCBiMF5Pw7/1VixXXvQbQe
61JQKEF+CVPO+s64/UQYOmxU8TcYPKBvQqFGIr+11cDET8FYdWqdehQHHUl5
XGSi8QQIY/01fD6I+e06ELJMXfMQep5+JodauaYLQVwZTdXcQoBXpFO04O7j
DRiIitax8R/4LAYMIfxWrJdgQnRnuTzE1fLwUgIuFA+Ccl5FH6QLTVHzOd0s
B9WE4azrFMq416XHu3VwZt/3YH8q+6J5SfHM2GkXwv5MGGYP6gfxYCG9KkRm
R1FdK/fKPBTFVaNH8NZcm7G8V947sRHPi+J/lkRrNXKZeWi2NVWq96Fmm9+5
zlpiAuRLBeZ4B2xUIdYHloIJvYh4djY29bS/CGBqMSRhR2DyJlVMJ7Hqknu4
a6tqEyIkG22rIP+4u3fLriLq56xKw3BaKoUOP5IS8zImylPVmNNezwRi7vJQ
19G06ERsvV2LFBx4xe+ph7oSvNtqS87nT72hA3JXrFaV75eazdLeK8aGYm5C
8njbbbpGVafNt4XI5SXkcfHnx/0hvDUGYGb01vEa+9S6saXeSTepG9HCF3jQ
lRZeffckwm2Wl85aXRRkqbO68kcw5oTY3nSdGVdYLh/92WcBqgv2VlZchZSR
PVMaob8CwG90Ny0fsWI3XuOgR7yTG9K8MvDOuo82U4Dq26/cG61ZmUpXk1CX
mfYai6I4+m65vc6R4NwAwPgXEU8WYjnSFx14qDLicBcpluE6tOWtmK2myRCi
T8k1/zf5h9DB+bsCWPQcdvLOxwoxRMvawhc62/n9nG2LfRhMqhwxeIMWHprn
AlKj4cafJTGapD3EaefhA95oetNpsBXe7RRBq+4+JWvZTe/Ct6FPgMXQpQSg
UKFVqtl8TpPlwa2tPTGAfSat9+e0HaC988D7Zt0A2PpFpXTxOmqIP9n1Gmxt
Tg7SMIFOEJg52UEhbHyWLliAXf5ALfl6HMBODmZYZVpuBuJoXJvj0sqI0cKU
dx/HfV+l2CevsZMoVkC4sfStQ0r70J0ng+hbnV4iM//ZgdVaYV1uT3z4p3mZ
A+GwPzILiNEJ3Xl/EOFRnGSWiflZ0pL7p2zkM9ZTlBjTCHAyRpR/eNGb97HY
z05WerhifQnSAUMZaxqHFbpY+c5x7P3u1dI8tShToXKmzlXcKTmMFEDuJVKR
s07SaxhW82iq4GdjwgaxFXMq1ddsgIwpk2plrkVwO4m5DHsT4szeU8EisjeG
lR59+9uPiEVPMZRr0RJch14KmKE9ZStqhCK9QxFwVWdVs9zXapPP+MQEqITm
w39naw0/xjeNfhg/UtHYG7GBPoWRGIWiGeiHSLbrEB/YNDgAl3a3QiAUVN2p
VX2Tcm/AzPJ0JuVtkTabXeycriaWuxGCm0zFWuyGaUtX0uRQn26bpFfjMS5w
Ne81fj3sjbtG0IuMiAD2gvMXHMVfQKmJEjVIly+YoQkRSAosXdOq+4CknOYm
2pCfq/HRpDPo/xrY652qiGlgvSfsMuvtFlK69HypBt9lwUY1MLhX5TKzAubu
CAFkFNjNRd31f7jqA9t9hQu/q+poJhiVJjOTEKqkCJOx1jcoP9L01p/HXWla
8a4uXWQl6jluS/Lhv9Hi/iPCp3PEUBoRGvkrsZiNeENM5t96iHfEfCQRWqJB
onp3zObF5EXzZPC3hTK8R6bcapyEqi3T4Z8uA2Dkq3CvBQcAMqlCaBIVcL+1
JKC0yid/hjMtpL5XOKVoS7SrbLIt9uG3pcRmrj9ERXsPVuwKkN3LFdWXfSHM
Ma0sWDRR3+ZFavj+LULV5pAuip4NkDuHbvDdSCkFG3sAAt248zcBFjuhxjTe
qAqvB9YjjcBVLKY0RK8aJh0bCySJN8Yb81zo5XW4FTXOI286Bk6jprHUlSXT
RPS4OOpoy9Eoau871YA7EivoA2UYtA0qXXAWbd7QtJv+4NjyjbQZKLibV5vw
gMoF2DwOmOQsopMIDiFSUMHXiIut44H9WLdGwjpIvadaLqAl4sbXtgSIlXvb
i3EppJL6z7p1EFCICQKciqtEER+/U7ZOF8j85S0JubLzwJO4vJVAk1Onbg/f
24VTrFUtUHt6ksbsn3qiFLBO+ZqUCzrabt23QvSZlEut8D+pnZUk0xSxStDx
7Zgi2WLKahbpp7MoC32vBjUfKxoGXzup01A5KriHzRc8IMKXaMwNSjEqmjPZ
86BJuUomfQlrQofxaYu4gKheAqbf6n0URGAhP/WVKq5zljtF1PSP/B4GgyNn
EERJOY4AIMeHpskkkTzdwJHkc58gfi1epi8oCBmfFkKuprJfkdPnjHNTJLJw
PNIFyzNeL+QWtxT0nbiwDFJ3HGnsI/0hA2311qMeJ0U9H79cstes+dRj/QEH
2+XmBcuInHTER8rznBfcZZLsHYwJsWpHS2R+SnVkEKqbjfM7KWrXFU8gtar4
PcPm+YP9JC8W1nRqqPDaaxpqFOkcXBAdeeQTtEdWf4ec2OQudqD15t67/ify
rDaCbaSO2zavvQMFKNWUB+TNCwSUxpyfOoRyH0uW8jfoz/thabTjHCtXIlD5
2KR6/49I2vKhQGQDos4mGalD5pGxIG5L9alnqCUnmsp/4wktQNMBz6BQMPDV
yL6WEKkFeGxUi14tJg8HCyw/W+SA8pgefZktESte4WHtx1dPjiOiK4xQ6fGu
wsb7SIojQr8/sRwaxwEHK3056TEkf6pFw2WyzIv8z59NKeiVzPDxB1SBO2GB
4DEUWJLLNQbVxq56+9wN6IWtl0zGYrZylCAy2ruL7JRMgLFNH6RictzR1dEA
zUq3YZDQYQbVTS/IgBTKtAqyQ0Gv1nwazWcm/nqDmn/dW+6mbmMIIcyjzyPP
dZvlc8/dD1j1Na8XpyPR/mqIe4VZfDMHu0VfFyY5jPhDu9O+r1VpnQL2s2CH
H7fx4rDMH7QthsyXvcdbFEf772Gegcfc2KaeJ0mQ2ogym42puF4yaez/BpE4
ToTViXcJZ2EcaXvIEJWhGuBPjpLbakLOXpLlirE39sSWg65yjI5HFTVm+yxJ
nS610eHNuB0PzVBe94K6TFROMOeK3XEmwSXxw5pNfUCaYymrVzr8udfPjS1K
FiZgqRQFSNMCwjwTCYl2Ns8gFet+krDjWeBf75fhUzETmE7pfUWpcdXJmKaa
640Od6+3ZgD+/DumAAsIEJCDEOo8dquhyJqRJ2PY/UOzPpy1ma9nJ5m2LgVu
M1567OO5rr+0JAuAZbBXi56NcqyyfpGg4UvAugjwCHcXA/a1CBV0jC7w7tGk
VGZCQOb1kFXHqk55y2/bFqaPn1HfUP3ZxsNpQJhvBMqdD2604Cj3nE8o1Eem
c/J/EoRZrvgMOS7JL56iTkH+U5JSglzal0LkkC8wWnTzV5HfPKsdgnDMNBaw
vV7F+qvEXFUva8oHRKIQMyLQZuCSt42HYzMSNE7Sp0+gNRdKRmtByvFS4fs1
Kxl6fqJvfBXUnlCGIEEc4ywWfpra4G3aFD4rRlFn9OPv6eyizpgPAwu1GEDI
rptn0Rjxafb4lRJ1MYDI5vCjJVOZdjAWAfXS83bTIPo/aci2FwNqfPYXEQw8
hYEiLDFN6XJEd9D3y3t71fXjX+xl6xLDrAiq7ZAcPQlhZxI//x5HDkR4r2aV
ca0Tw1RXVwLwempgnRmARwV1P7zRcdwNiC0zdjnfIUIShiOscu3uPRBSKNdS
9lz+LyslpqbSVajbxai+FYgGNirEdtmBTk4b44txradKgIbn8Pg+H2BwkKW9
36upRuP581yxSw7o5oLxP6g/aEM0yC8/hr4bNFeQvVU9F++w6MVoL5fKeUc4
kqv7lap0gsr7MEmbilyiBd1m1PIXoEEgHujCclB7qGl8LvD8GL4LWV7Z/5OX
3WjQktcv+PgNfPINPIMiAYm2goxxBG0NQYxKNhmIkxAEfX3vCv6EzCP8nCS5
dXQJ2wL1xfDRYxMFZJJwdzGmkKYzY1OoyWKGlrKjaS7YKzEHEzdWTLRnjYWO
CluPy74fSFmT8ZhK+J/NAQC+XsEtJ3pSUpuvXCQ1Da2/kSnXFZfcVBTjalM0
zdfXMJFE557hDIlYwCoV1/76UMbgokEmWcKH7gd8DD/aN0j5Pd5sGjoJ+wkP
FTcZ4tvJOxACYXVbfFZaO8dvcrREl7Z2hGgeJALqfrIMq2nN8sVjAlv7uD9P
2AKdCl6nfg73oCTNo7MiHw5XD/7VhCIST1vhm7Oh7kov+jhjQzyQBfNEjL3R
Eul26KsYy88J0LkxyG/jxxpRc/hD4O3kMsTngk/J2/jQF//XtEBY5v12IGHO
hEG7GDct7Ar4Z50dTT46CbqToXjxF5C/qiXnL/GEAIuWGtKM84YWC2E4fnzU
oRitELR4mDWtOiv9q3UHGISItBq1ILK6+zoEzaqlBm7+Ne4K4lYwvrdmik23
Z83zpqEPEXYA5fSpl/95Bd2YvVdXhDRdRUABai8+kGMgLrWru6XIwaKVL5P1
p2KKyGY3LGCvIBFe9BZ7GftvgOdB9q48skU87pHuB5xinAVDRmDAsUeKoz4p
Kgms/xCo+Kn6JJMg3J0yRg+D8yZo8OQ+tcV54o7PSCDm/n0kMzNr16SV2D0a
72kj6HrpMR0Ig3JSRNmdNDIx9xvnUIq9f8dJMcX9tHSXlyf/GLtr+FiGXHTN
YkHgb4T1YLuTpOE+xCWhNl/yiK96sIkwb9vv4IRFtv03O7aVXxbSbWoyxIBO
ZSF/V8S0Abm6uvyrwUZI8Q8KEqjASaeBUibe0leImzHchqs9FJYsv6yPnEa9
muQqkLIshq94kCnlR7rSqpWJBSAdqV0KLJrrrU9XtBenjmJ7y9LwvDnwHX4l
BV7OJOBc9LU+imsqJPxNYscuwmNpSSychu9WGuQKJ51/rSgFuJnetAoh9H4l
39WaoLWXfCuAEuOpYZMJOZNOfIet6CcYiGQm3av8JTWqaOg/MCrr5G2wIf57
HiEQAk3XsZDRP96Vyk9ESRL1VO/GQz8qmxy0Ffra+7dWpjI/Z0WjJIHyYdiX
f52lJJEhv2JTwN5dt5VDXg/N86MEMDBX3BbWoAWYWdk4k3vrrYs+d+RG+/vf
B1WkFO2FyzMNBxtoro4IlCrfC3HJ9DpsZ+6LfSZU8v3e5t813+IjL/gxlASv
4hBkTF/ClOi4PFEdQl5UcmMLS3f3UAE1s6EZhaw3jRoGLD1tgRdNojDtrH+Z
b+v+3sxR7J6go2eSwN552rTdANSt/UhCepoUXVCUTjHN6MqRcSbAohkRenA8
IU/dcyCUY0CIYqdxLln78Z3kecCk7LPyOn10OySSEQys4s04facK/Gw4SnDG
iIMt1pJPEIxIIeagedlnSow/uEWKXFOwol9JpP1J88WsXt+nNlN8sihDHxOt
VqfpZXMf398966q7qX1JSjo69m4F6K7ePMml3bm9E8CZaH4CM2vckafxkuBY
hwB7i0FDl8boR/bh1LKz2iJUyhfh40PZqmpWITPCQHJd2TiDGwj0GMYEjbXn
v8sAVlcUeTUMaXQ4Piv/q7jFlusplAI9Xp+QA/WGqLpi7ckC16RBSKNLtaRQ
3IgKcME0QRmxAavVTPayClxxpHAUoBqTXxyg0YeHT6cvYk7/uVr7qV+OgbKW
fxBn96E1kjsT4IZ1Kmkt0MxzXT39v2fe/uoJQnclF4Fu1fbTnnomRUz0Rwag
60XtOY4E9NKfZlcwVBx7mvcInFxvqfiG4fm3JSggzE2Jwk5K7p7l5B19HT2F
ebTLA0F3i2Z99iTEGoOaVeMQlnq8UJrUR7EbyfM2meCFcmhEJlwM0w0Wd9eA
iogHUsfgzC4dyYeEOFBFrHhFkW0GjQeRqXbwnh9zt8UGkLusQt9ccnfydLoO
e7Pfs8c3hBzjQxY8MXTzmTo8um/z8Z9JW8HufnQ4+TPzSsybsu/UrW9ZGUFc
V/zV2AZ+5Xnq2q9sJeIpsXGNxDldMnSz0PjGB3zhpkRUgLh2HZ30e+kjDCFv
xi3TG0KPL6rm/X9x11U5mY2Y+Wfzuy0Od82BpKC8Lv77qJ2fGLWeEsSLm3+q
pKktO7ISIcgxGMzERyDlx37SmOUHpI+vm9WagPX/DkiJtsziTNnF2SIY+fdF
G4kEJB8lupBQlBpuuVB9jnWTufkh6JW/W60BeK9GaIEJjXrdHeoLTh9U5kxP
rwFBWDLuaAtTXEpGYFqXzXE6VacOUf5X7uT8UzLQD0OJ1P0fHz2iUCa4OMq1
Ayv9vkXh+rWNVjLoLrW8swGWa2lHSIpHzMF1qHvxb/lc0Txq6yxskmphyfhR
NYHoy+Jn3mfZW7sJ9AEy29lOxJ6b8M9fupx+W/eGTFIlhQRK6TsuE/9nvSA7
bkWq3yMsnV24QvAB9GUlspvfclvVDMHTe48N4Zsu4KWOiJ8CI9KnVync8qKZ
no5K9uFEJjIa95Csa9K3wuoSX1QB+8vstzqX1E1+Jc5LUclLBY7sQ/cI+TRg
ZzUTFS/i2HGFhbZXUy94aGMO/cHq4INXOZstNLlGTvRArMI5es0D298zFHZC
AQMG/U6sVWjWmf4w3LSususTE1gUzU6f6ZZCHqMVu4TLWf17e9WZ42m2PonO
9XrKwqLDR9m6LHjeH0Da5r375R7Iy4urHRrl/1L8Nf37zHmXsdNg721k0Jnb
doP7INCvnuG5fe8TWBGSLI/+3XWsamFQJ6o2WLHCm7m2REgaa5ozcErC5vyB
M7sA0ubgZ97FAvTOIfdRYjE0ZZkR7zl1CxewlV94b6v78IrU37+MnEqW4TRm
hNw71F0XpGJ/9onGTQ40kS/c4OoBVaUuBFltRk+LSsnAqvHpAUfpLHLYFIpV
uzHhcZFsEaE08X0SjpPxy0WqT4f4Q8LdRwdaeG1r+1kRBve2ndo0fBuS4XfB
Y9VGKUWlvP8F7Fy+d+WjZLRQLZjG3qVTkCXV2dQtQzWUe2c83bvSoOSEYyxu
SWQm+QxgjHoEO8JG9dvnIEx3Dw3QNuG8fl0hVfmx7OoWcQODpGtb0VAf3XZe
P4NDhcTieCOx3ldcEPPLUCRvOnRK87cUqLBI84ONW/NE2l77bhXom4PIWGEv
VOjU3sbXyRTWz3QmimvqCHuwCZFhp8+FomNmaJ5G8Y0wm+JDKaqTJlbWiTWJ
hffx7Hl/oUmDKWXz86s+G77GbqYabWOgjK8ldvuM/kwGpFN/pQV08YdrbXj0
tsjCpQDFbKHtPG+KICgrm7yTKDGcTuR5tEfW2SfrNffVSE5BxehoDid3vcuH
4D6y8/R6voQVgTl6m1BjZD/55MWb+puj6CTbq9yd/5Dsmkq1Hta9SUundTHp
v95727oyDQWvZh/jndNhobMHDtklyh17RIqi7KDG2qGlIpi50UlOhvcyDkhk
uXtF1HcLBzv60dmvxoOhaPkk5xPU9a7FiJlqElyPFhgiQEj7ks8e7FmYsy1K
hN15Pi7fqw2sH6A811fsKmtLnZB9xs7342LHxPIFjAPGps+cxnaAgKF8E5AS
xBZuxJVPXfFa08jeuS7Lgj3i8+EC7C84wICaMzHhadYU5Ngznaph83jhdex5
KNTWvHu6TszeMZmVoJfUMX/A2EBgPwUAsOrTf6aS5TE3ov+AQjLFIWCmsbWf
EQF+GhQXl6bmw9QD7QI20lcBZFiLOpmFBvmSexboS/9i+YfAOeanu+s/AwrI
xYj14p0O9jBEr05fnmdjfftYN4sDdkTKD3OejlyAP4OcacB7yyk1dmtVzw2J
weEvo9TDj1UrbSnrpiwy3cNd9FkaGNEWb2QHE2KC+o30fGEaXlYkv+O5W+Ka
EawE6VCg6JLRI3O0dJCylk8EsVr929mkU2tqdhQrGOzg+LLrKXDikSVIOxeq
Pu/9qlc2QzAHUdN9HQNFVY9JNFt58I7CdG6qk/X+YRRzHWjkhuM7mQGH74B/
wV6g5/rb7EymO4DC6Ulu20MbOLongGVSDKroJMZN0GeqkFzNH246qE1aSu92
dKsRyycSypOyq8ho3p/reAodEwQB0W01LNCN47KGeuypWtVZdH/iicdwgkWn
Fqu/gjPyeM3PKvfXI4rS+XGYdjcSvDusDwoPCmjGX59trA5f3kBdyF2BPdmA
vGb1326lzpVVCiw+62xJfvPXJC9KT02VWTV3263f/qNHNTmG/YG6YEuXBQi9
ksgKmG2Q8xuzP2DKoXksDUuWOAR3Mwv1kY5NsBUgVQ4um1c1xD/99NDghpV+
1aIsh+EoDzrWjjJ+Eqfpl2lI4WQPZc3L9Rw0kkxhFySZkIHXgrn3Q4f6/6h8
M+LCJNzhM9QUCHrnZ/Mh9QZfdObGmZ4WmYxqfNk6y5M7mOASzGR+rI3QaUVJ
p6Rviga5mcQgWYXybbCbV6/btu28A4M87TZADmni5TpnP6pBQ3o5CwYIuKyT
Shxd+I5YKYIiLAvwdzTB78OdyErce4FWH8uXik74fajwe4wdBNIVtz8fli9b
g6p2cF97iyd/hOHhrjJwt1bQri0B2HxBCxCMI1/gv15/+eEqPbUT0ezlElYE
TKmljybH/79uGOwOTRJv4suM1clfX8QmCUDMv0L2F6zqZ6KA6xh4jy60YAso
xTjBHE+jAGNyW1e/daQom0640uns96kli9iYn0+p2wmbs0obvJFlY+ROtcuo
R8L95dbXR5xTRNJiT596iR7BqsNTWfpdIZG45EmNo5NCRsjrWsjPuK6QV7NL
8Hy5RSV1f2r10X9DtlyW1mDNnT/BpFR9Ienp2RltT7M/yuzRlx6XxpI2t3Qd
REa8rWiq/Yh6ejF+CqpLgnQJtsRir6sUNTUGqOo7CYg+SXSTGUXTT+xShwMD
K847RaAKZllFveTHUpLv6/uiagVImaMZjdSdGh4UpCtm2pB/PNRyh+fOqXE0
F7bwHF+GcXud5X0qq/qWciasaZ6bWNR4sQw5AsC2nQspvxMwC2K6pgHXrY5l
beaFp2haAFQ0+8Cvgsn3rStd1iAY1L3ENLVHPsIgysyJbdaweT/QOr5JPcQ7
SMUbXTejayb9r8hND8GxUoQzcIouEc60fk18FGQGjG0qF5mxTyXDJZlsGZmG
dldrtCWCHzqCkfqZlwd4AjIAhGs549R3PWo7W/JFzFCw8QqUhOMugvYUN8+v
9hvrF2pCWUYnLzDODZOLofkQMZcK6/2Rf+g6lSvMwCFfeXAkvxM9eZJ7hKb8
9xY3w1xxNvbBQmL8SeLy6czgRV6gHBPvphIK090YSEGT/s6LkYuowdC/MNZJ
+R1EfaaQo7IXshTW+ndyqpvRWCxrNbdqFp0AacYvyI5iuFza78BK6hkn+0ic
TOvWz05GSp1h84/7vKL3If+kKHY+yqEiKfwbNTzS5VRMCu9nyUQN/QoA5jRq
OswiSxFEWVJkAwNuyicy2ZqIkkZTZA2YAAn560lnJ10htA/FWUrre+HgDoT2
J9VuK7SNMlKDlwCoW8K7KXICzwXjTRmmYzYzylWaMTnZO8biOvNr6ayo7e1A
ZMjsTbDE4KLRvHgYzbIp2yGL3X9FUhNoMkJtS4B/ll/tO05cDphJbQrhAf1l
2aAy6J9w9dm69ihywGj74XRTxqyi/eZkreA0K1Wgz6NxF/R385r+gDXthmt1
4zMoKCAwgjEFNVC8HPiQCammxMyf3aDE9XC67/v/uqekM6/duDPpCNlV9dqB
xESTTcnZmZ1+WLNrOH7t/YEmkX4/2bAUjAv0Pgd3vyCXzSI00X1T/yVY2+to
kd0LAV3TI5ung48Uj+r7W9IZQF9dr0/ZTVqP1SMqP1SFjPHBTdiTUz7z8yAc
+vv1K1RWHgYJATpWRwgis1G1hP/jsODahhhjd/NoXzuRK0wFRa7XDt90s9bj
5QVhsG+4qHXHCsq2QhWWEUbVJJ31KWtPoXz4gr5wEjtMM6X3MAT1vtn3svEZ
skX21Cx2dPKMvhv8BFkCClKuupwW4n7QcUIFU2fG0l6CFN2bGiP+NbVPtBqm
ntRtOH1dTTn2yTL2jyJ+94IL4M1+RRgKRSKd66HkQhn0uSkCndjAlq3wna4f
XTP0qHH4iaC1BlMk+bcslRGhi1BGRsmtXoXCdD27G2kp7JXK35zye7kwESnN
THUssyi8+BE5w+WnzUATWR3XyfYhWq7z+bvOjpls4wRWWtZa6AO2e34Ut9wR
gyhyL5WHWEkQA68KdyNXJp4MV2qfiaBPOAvjSBc+6q0peNxMzfycXRdmilQA
g4fOK91pcEWQv2pWo/owysWl+sOGj2NYF1bhqOzb53t7Sgw/ZG95oF6QqCK/
ikY68QKPgYDOUUp9EnwAGdRl1R7+rcXDOKePh4kDb65utCf0Przq7y//lcu8
TjXuXD60EGQG2Kt03iOxXxfG1xUJ576nJaVzvPcrzGL8CTj+IMqfya6wTqBU
Y1Xsp5P4fvq+9MwfSZc4VTL8wMDtrukp5qTISwfkGAqRgauQwROfLcIYfn1N
qH8PAMWtapU7xvBI7qY75a0n8Ju3bLia7/NvUWigL0tsMAz65KTRRN9iGjQp
meT24yo8g3g9ENRweQCRaOyarXtoDtmrFIN45MJ8a0SIlnhHNpbbJh5r4/2G
uoOM2P6WUhd6I8U25nwyQtRi0UVC5i+K9MWpx4SYir7LF0GC2XjwHNTB+xdx
jc0uzrEcIF9YKkPOSUyOv3thg5IFQXDzrRIUzQ9WMJYy6epXiQIkKDD0AgDK
FwH2IFGnz8VcmRf3cR1BS+2+qrWMkiOeYtuw8uUauegEMQxnHxvqkJXz7jcC
Ko2rV3TsqhLnbw3IjM5lYzkduoLfKOgBfYNE9fNJ3cv04dzMGh07J4WrkTN3
773mop99SlQ9x5xyF5RQegaceHGYnxdD5DueVPZezbkMT7rw9PAS1Lf0re6z
CeglZcNnQoZPdKS2+G+6DYQ6GUMObSOqnIJZTTJRytndsMi8wK2JTMBfmNHi
9KYlqkLoH/6DTnZGAiY0AilRkk43JZJukoNJiEwzs5551u/fI2AoXPSzlgDu
Id15QLYC7rb9ZsWqSv/xDADx3nExGo3f74M/4JYCr+RNNJTdweh7jW1xchJO
A6+Rpl5wCUuiNZDsYQxFUPxypXE/kzBrqv3gI+dqbyvX7ni7UsSVPAG6jqyn
qtGdj2fGtwSVBHuSb1haxSgiWKzECU7NZ75S3iyghzlacb9ETAqM9m5Vp7Gs
tbtpec/lBAmNHUqDVA1azesqnC0X8KQRld4aCPWHJ0QZYE8H6b2Xe/QWjotm
iWdrcdUGoabZP+OQGHfmDrK2RYvvXm7iTDvM79nlidhNbGeuJ0h4pl5ZBWL/
+DKA32gdtquw+QvJmBEiXaFyaYM89a+TBE8rwY2x/zD4q+qfUeZVYsgsc2gE
/PbndQhCx7xNbZGwEktnc+/1sRsn5hVsIygQ43GSo5/pMvGqlQ0C88pwGQKF
4P/qIMS1PVQP1tQDXoO6uyof3eQG3SjkSg6PaJLEFRDI2nJmX+cG/C44k1EP
4WR1EWl3IC0Kjgk+EhPGRDsSzM3p3y2GB7NZcox3VldUFPVF2H9iGze7kO/C
a3pOFwpW5GxTpPmhdQMRay3+A3NBgjMoROXUIaVg4BCGKGJ3tDEGRku+p3Ge
SIExp1DVCkJryLTMI8kZFwTJZgg+udD/eP/szvIgUi3+nbFCg45OsH1MOmLo
cK7aMpldel7dArlP98dKSoVdlMHqa6IoMQz3Lk/vfEhgG6Nc1cKmC6huHAmn
SeFRYKkzoA9hDEceEwAfY3dJtGcRDNop45kWUh9OyCd5/2YghWlFb5WWDKmt
QnbJLz7V1QqJOFNsDbeRsRXJFpr32Gh3KuF4WR20oY2JCSHZN1Zj1HgZ52V4
6IoqLzXBZZLRz7pnTjnJvNSC/YBV2OiDzPu20/9kE2+vfeIGIcwSkE/lZXnm
N6CxbqWwournZgzCLt3AqkpFAaRzHjvlXTdMvwyNpM6LPtT662yl3UONDtfa
MLBJvlyD3RpmX5JdLUPBE3PI/U1LM/wP2IKzu26DuvzMTGRQvMLHz6HRp/od
CJJh4YHW3gd2mr8TnExNWkjZdKdsLObAH9Iy/YnNZ4Op3IwKkpK4lvvthBU7
buTXthBoSAgCZ7tT7IZBgfI2SJRJVTG7q4pO/rBcPik+mK2Ty+zt+cBgtuk3
QcW/IPTaoPmWxK97qsIfW0vsOil+S6TV42bAIkg7yOv3D4BCnpYs8W4Ko9ha
5Yjy7ET0ddFBFLS47Gt+z4D/iQ6zTFMD6PtHI+F4IKNIUGfjyB0SOugllr7Y
zQ3a4r5TnHcedAqhso4fDlYOst+TzpGm95M+AjX/lWG6bFGyQXJSl6fe4xlJ
9C4hDmdV1RUirPvy6cnVAOj/IogT0hqElc7VbGxOR6CQhp1A/H/E721nludL
xu+zEWmFdJhO45BzNbhDDRMEOCHHfX5cdglMOruUhbJVnNkXXqnf8bcXD5G2
fMjusrZP4SkMlfL6AzxH9ms3M94dNf+Y4q8eQaYw7SA481AH+a01uCe3Wh+M
6+Z2HxbinkYkyVFjtov8cmV8gIbW71AUGn0dwK0AqC6p2kNLZPYSxN48gkqi
3rao+y5BdPJ26l3A6z7UWuI8Em2MV1T/jOFYr7WJ4kqniFPr1i7WZSYJ4Ib4
EF8XbXFHN9EYkepHcliR4lfQsAQPu/M2zgU7OHkRAtTlAXAvIcor/yOxhcag
s/LM6hAv5geXfVKYt8CNnyOOdniy+ruAHo+WTH9KwOVUqMOqbHUOtdBDQK5E
x18hFbtvXxIei3fhUruaL+TI1u0WzjMmbHROnEU20WxqJ8InYRMk9ACsnQTK
m40cObHU9tuaGeOnlvOmtN2drQGdWdhi5AjYfvBmruaUQgA2mlr379VEvaNs
2mPlQt0pOXGy4siYoXxivgxx9aNbJxJ126EslP0ZqJ+uKe9ndgNaw4ovI20u
360SPOCNug1xovulumDAelkHoHehvFhpSWTZ59kpl1DUmA9ZBNeJM8Ym0Ka4
JcQ14lomBO9MiAc6dtD3n0ZhHia9i3ov1UzgWyJQ0M/ncEBHgB+Zw6L5fWL3
m2AgdIH6+VbmBgYLk+lyWESi85NIW532f+C4phoQ5qKY83fTHCrxexdC0wvC
N+kv/xCWnmZ89k491PpFdalvB7OWWFKNHTEAdwe/eUQshcCY0Ee8qbXwaK1+
e4r0fdxMsVPBjq2QjCoPmKUjIF36Vx0bNLtdZBaaArBR7fI3vpQPzUMBZf5p
PBePoPvFdtcnVcfZhYKa4QHK247p0DlRxGO7g/e5l1qdKTj2CaYjEY0i5iQx
wpGW+JTDohMYrag6tBU25XbGB3o7eDEhy6D/EMlCNXvs3++Uy0/RPbhySbyh
3vHDIbTzZi5/tkMSc6Jbf8g3jhyGxRyEcmYx/Q02+6DubDr78BEi1K6z9vQe
i3zQGdaoWk6VGFET3LEoEZnTVIJbL4hfB484biMG+GO2r+nPf71873Cg5cEe
4S4SLG9udDYVdl08fIIcqUjFoo6K+3uHyx7BNvK51V0iuhDlGHM0M3pmYU8d
1t7u0enHf9Zo4yWylxRtYfnFULRusG3vkTZsudhGzGkjPqC8GGlOgRMrQWwC
WsBZQ5L5xxg0ASapqD6n1vKFfxU5+wma69YRq/oP3iI+uouJcaBm5nLGitVd
iwMYRgFkbWxDYD5Dxxi/W4CyHZA+JlgUW9bym/vSkOBE5GPPj0Xu2XFjCvWp
OCenyvhA0ZZO9b5KxOglUv7cMLd2RiWF7r2gfNeDxN5Xk1H7uTy/pbzRe85r
k9z2xIUEIQF6K9rkUa2E3qVvU0WWrUE70nRo2u4nY5kh+59XWcAOx6xqA5SV
WDA2lCRYXWUXEzqQa/kZCLmKAs9Vyz3eVrmrMmkefncLA22NpGuJdaP+g/PP
Kv2+e8WKOss4cDTuUeE3DtUhATwLR8sgNiAdrAckJWyWzACVjncXfMRwR4oF
ox9sDI5v/2RxqNMUWzLDJihghIC8Fx83ghCc3rxOodw0mqInJAKLCNNwFdDX
j1jvWOhR6YDzMleN9jOiBO+FDYM4gKY//XsiT199BLXkl4X9XhIPGmIGfVze
Tc4lFSfKjNtU0tQdta8RwUjQ9hCNbhgFHA0Qc/EUR+AU3V8e4n27FOEnCML8
mT8ZVJaDRJAqHvdtwvvluUrrNyh3Ku2BBsfEj0vxZ7sss8sZjXE6q7AdPg/Z
2L+HW9suyxt22iGpmhmuNfRj8GGDkD2IkLjjzpXlNejAuSi7iR0BlDZFN2TM
oKIQ0CnlnecSjlPb2f7aASzgrzodQq0sLosNREj6jzbEcXZC04SHrLF9PU8U
x9Fev1xVpit2L/coUTZfkGJNVxpeyU8UUUa1OAWhG/ebvQ9a0CLYos8hAF7Z
pXmWbnOinT8qrtTQcOUtfOpl8sE+MgILa0eYRvPW6BGCZBy83sPInR0/BZzC
4wiNTzvatj987uY5GfckIssEiMCPBE7aNqao0OIHnSrF2nfcxA+tmJXdhe16
dPcmsXvL+iXhjpTjYG424lm3KRVQBbBVYasrOuRqFZRpayuhAxqQHmr8esR2
l40M4EE7/s1O2f8fPspL0o3meAsGeowum964pgnTUjxPEYqtz7PTYTqJ370L
LkDKxluARF9fnjV+eqFdAjVucpeYhLXbknFZazRuxnheCxSYq7W6pamJYsRc
5lp4GBdSWSb93cr0UxgsgrJkrIqqBJiuSBlUmIarI9TKj8MNOYfTdiSxvI3W
lmLKvb5Ugqb37ydWHadlduQiX14lhrROhJ/6U5891104+vLNCacaHBD+ifHQ
doomLYzjSXY7C+zHfBd9QdVsrx5jQB4SnM2mzMD2Ae06/kWtIL3PAsxRyHLn
lwuVBOm+SrH5Zr/6FzBkkmGBnM6P7Enqnasrnmv87hry5R1WT7NxDDpXqcZE
yx9EX+7rZgR0f98nch6ATW1LGeCjIWavUFWcqTmWhMH3lLfKBx8VVIvTcqqM
25fc5/I1JGyZsG9nbLjkY2/RWhLpfinAVzytg83InPDh5sw8NkRQc5Eum8o/
+/xl586V1Ei0naJOntRE2fItdeHxpfHf4w2tWmcxgHClug/B0MIwVzpSnFGw
Y3bFC5lq/LaSQwu7TkYcj5EzPp6XtpRICQFjGYLz2MqetdY3N0YTGhuaUnY9
lyDtKgWRiKsCrL71RQSJnPoFKCIAVDfEOlQrlIbpPLsgI87AO9bQj4GmsYEt
S+cyyGCwWp/7DDG8IyTpscTvhlF7P3zOU7NhgUrro47F4LG+YagMTK1O2sMr
UivtTf1dAItbCdD8TALibtb+GwjRs422lrfda5T3ShkW7pURJBaDfVa0egGQ
y1VsR+FiiqtS0eP742vWmyLbXWphvnJoOkKWm+jji9g8W8KVItm1hJtb2KXf
ek3AbVosbvFQ4lFvI1ZGYgkCcR5sjKPESGck2Z0I1E+UkwABl0tA/szUi7/v
ZWIDKO90cjIQ90sWr/HgBCrewz2YcAsIc1KKEaBPlndMjL/Q2k004yNzmy3F
mSpzJ2v5HQvJe5/ivgJsi/XXDkD19nMBmh8DgkCf8la/H80ryNCkOlzYXG0S
nH7/oGC/JoQkyNmENpjN/bKFQyKj7k6kbqi/GIizFHNxorxvLOqCysQN7DRm
8WCwl6kFBRiK+G/wYh28DfrTYfIZvzehubU33WXvU6gijqxvg+PZ7Z+6c/rG
UtgEZFJ9izoo63oTcZHdspvJuSglgglkA/cembhF1nWUYpFVfT+GX41eHOYa
M9zTDAir4xuT0zr6qYXMnmLLh96j9HctgdE4d+iiy2ltbBD1pGMsgli4ze2Z
qGyG/YHbz0oVVYJcOw5dmnM5CiP/8n5eesea3sT4EQBth6oKV3azihzkaAAW
9m8P+F4hod/Joz7FrrAhFzNp/1uGQFeRtU+B6vtpvlRLdZ4PeehAZbWmoC08
Foy28G5oW632wP//CSBUnL02+jkvbgdGmq21+Nd7OYnOiTrSgrM0Do+iKnig
U6snochtaa4Sx8VwxnAmasof70Z7mw0u7f2P0IhNaB7WAC6MZXklgQwJShw5
GK8Ogsbe/bmi1mLZj30CY6+U7DhG7Gbt5Vr8hQpag46v1Ar1GDdyox8BpCZ+
vzM7obZjILgOyO6OFVhyNbS/VXbStK8UxDag2yLu5tCx3F1eHE/pNyQqOOxg
rw3MRdw2WTrzaXpDskj0TJqrrBqbLiCjOIP9f2kk1paorexmEpECsI/Om1B8
Ci5rjxgEQWmmCF7kodMhKaQDZ0FMCLZDU49rivqiObvkNTprtJTuSFS6g92o
x0qmTH2GkfrqI/XSENf90khmsbHHgoijG8M2Cy/Jerf+6PPOLaPF/skYcifs
XZxYKia/aCh60iJL7x8EHtvHqJNtHV/EnJORB2b+tm0VDGcSd0pZaMyIwdum
uiSHhPI8Lo5jg7gi/bJsGxn9eeSlyYukkJGIuixGD6kbnzkU4RulQ6a+okwG
lBrI36X9R/iiCcwnlJmSxjRG0uf0omcFIMc6eCvho0qaQHtkuVtwvL4iXUK6
feOjk8NcVLBzmZd3jNNGbuHeLUZKPe3hdLb5j2jOeJ6CiH7jzDltRT+8sG75
JAvREHk94V+izkdVQE4QyZFehobblkLmoleWXmL9N5MSKgmsVN46lCCbSwXm
CnMoYL3WP6oNlW4uwp3g4s1q2KHA0/fNcp4wgTMw5m4w7IKhNa3u1yUYayN9
edtX5OWVxU9gJktLSyCNjJUVrhQ8ZpqvSFGBagNSP47Udz+cPVfT59UnBS+M
dxHTZgSToVi/LvK18CsVjA+1ZLnDeazuavHeFaa4AgFchq8GtYdOiCIYMt2M
31myNeYa89q3n9Gvy6+N915qQxPOaqnuDdiF9XgV5yTOfxuL6AjX2K4Ve1Ut
rXOzt+u+r7IWh7UJyYQXVbWUJ2g5Uybu8TApfxu1vKFw2PhmEPCNETz75pXG
icdKGHJW/UugN8MEiLbOXcl9mJ//qmfuymPC4uZFYHiQVe+8TsiumfuFsoHO
AMYxyUUcJRitle6414WJ5p7STHFFWeDdBoNnDR0m8UQYwUBD+WfWXXdDn5XH
rNoBDo2HWviLnCoJvuOlHQLHQPBe7CahutdCedRooITYtAQdgZAT/NNJtMuA
3mEjukEG4bmCQSkShp3wrA4EGyaQv36kMXsoyRGEvqYLhtN395OQQig98jU2
KmCPTU2O9c/buzDf2bSBjwtAATDL8pljKf5Opuk61mXFXKhqz7lDW4phrTCN
XsMuXoiE8LVOtF94+OEe3u4AlUVMhUclNJCHBpMla6/QjhE0hxJ/BOrsHwCy
B5+Fgb6UjCPV/839BqLxt1hMhJbVP5ws9ZmHXSPAJ1ZfTCV75sCooEtLQAWU
753/1aQyHYEKTn2aOKZoUDuSiXjsXKi4/h/mIke1ZKNXdklZU6XIV8SWHppW
3H5bigWLV6lx7Pt+RLWOQLnQ0Eunr9cPKJBKhU4ZYCQhU3PdfVJwhB0SV6XJ
iOIwO1aNRI+Q8BvgKTxgNOnagAM87ytEbeI/XHRuXZBMIru4GtSq2uT9VgBK
jVnBETBITUPSmpTQZ6PqsYF9mOoq0PVx3yzS6wSTC6Wpfm4M95I6tfbPgcAz
idALSYAfaIrCIrHw2oz3RonhDCUx/IZ0Vngmy8I0sWgmXFf4SeMJJZhPIxMB
imUh/6VJ+V14xmaBeBEM6W1dH7UvWxEUUox0Mg3sHzKbGY/FUi+eu8irZuNe
Eym02bqCrbbwOgqBwvOmlKQ7q50Q5ARGK5FaJzFlnjtokem2WLyM22r2zOTV
F+bfHimU07HRAp3xxloKoANWCRW2g64mkj4i1HlZsjYlRyiu3Kags50EZVPf
T71kVWHgTh28eLsE+cZCZWSTZMft7f3yS0KoqELIJVr23zgZe5H68FVNLWWk
3dHBd9G+wGPz70jkB+4UQeK7bil1lpBLQGQIJ8Kj5JXBc4KVpbZvRV1JBck3
isiF5EUuQ212ZkAKeoY+J9LLv3s/k27UIC43Ktr1kIJPVte5qr7dBj+iN5kO
UyVpPX05W3r6D4Q4AP60TsSwvSnoVADV4M/xeu2rjHWuYWCQdZJPkkeb2QYU
R8fmccsspT0uE3IVfQrzmWa3a1PtysnBmtSGaGfwl54/6pZz/1VnruOCpj/f
abIjRzkTa3KtuSGLP49VFeybngm49ynL5lGwLjSlDCV+willCf2qS9j/Qoag
B+7NS7Hzx2qGBbq47nx4lZYQK6PsT4afrLWh/6IfcI1BNNYisR/dalDIT27O
RAbFbYoXGR+ecJBlv3xpPHZ724K0zZ/VD+vBZcd+R5W9p+7VID2NAdG3BXOI
tCsSgvj9MDQTX+BzYXEDxTz4HGr42pQa2ke97vx1KdUqhFAjhLYgoULn0Cxy
19KWL1cS3ukqBVQnnijk1/dirwbxFJeZ/PuxsfuToYZYQ3qbUXRSLcDhvaO8
9REf9AyIfRAIX9alsIPTuG5LaTvv35ltU9SBmcWcdtzQOzwaf3UFdCodVuZR
86ESqI06bVDiazPm0lfZ+SvrcgEn6v/+NRZQ/TBVOaze8GalAlv2IkSidjjl
GogJEhg4uKY6FlJM2EQcW8piwtK/Wz4bVxnmQwt5IvrD6tjOpxA94yhMbH97
FMkgPHao6iQUD55J9U+QCFaW+XqhwzEDyZWRbVe7RbbR4LGGnWg8PR/JArQK
50e4uCYYnt9vlvCgH6SbW8BSAIgXkGYTFzTrRU2GiujCANYlG9ZnVtryo663
ByD1pNqjnztLNRazGdJRGnHB/kXdPNVKbTuok/NlIUtyp9Kr1atXLQLrJqMi
Z+jQNEvq8fJZPsKyODZxmGeMM4O7TcJttrmZW2ziBw46UbHRlzrz+rf/aJXY
VbJuDmlF0gB8dh6ZEnlQnbLE+2kgYxpyZ8OIW3H2QcbIcveRqKWXTZODUWwC
3h5FMtHoV6cjnzbz9luwsEhsMSJLBl8DRZEU8w5Lgu3SFq7Y/m9zYtEHlphX
PKAiScxHS9iiT2dxfzyE0opMvLrVGIZM+ACenDFcn2K3Vw5PKEjMkEmGdfDE
cr4Zys6JCUx3Pqnn9pUDLpW/TxsQLLFcB6eVbixpFjFy5KvMV+f3wb88oXBZ
lSQu+6BjDqcR6Yyd7xyJny3Bff9viDbVwslZC/I07wWRAyVbez6w1YjSP5KH
koHjJeXOdh9mxdcs5GdMl1ZlLzOqBh3sLDiBanrayAyfXdokYxqTJxPMGCW1
c/KOQIn0Al18/3RcHH6Wioj+Zk12j97SyckXA6oWL0gM46YCiZFitPoYfyDE
pAnK5272fgOX8ZiV0zuDLQtJQG4DCIjfYiqpky6M2yafk48rMq2EwwdnVTpW
tw1THtjabrOSdEz3fIqbARnA30dFcYL33TDx7auCRXTDLCawiAioCdmrIGQD
1j37y5ukjz32QE4jdLx8KwS0MQM5Q+fzEoY88oLLfKcQk2Hld3XKa6tfrCpu
cKoN+ov2AVvpxnqjoE/VjPzlBAKF+N/Ad3m5/vvOFQ4JlU6kZcoL0YXUs7V4
0nJoW7iTj5LXH1EPOLDx66NeQVuDQLrwrEm+2Rinmh23+ZnReKpKnx1TsTR8
1K8c8+zZQWHvx7D991ENVC0AUKBo0d3MtxCyPhPA/kenLSzzwqqgMy13WT4f
jim+8I8d0FVzHI7y2MVEuNear76F3uqv0dGEq8RFQUfuCgIgF196xGNLBv+2
HEFohzemQJTcK+R3L4wvEbD4vyd+bPQ9af2nBgC2aVK1OcUlyVj0TpOucCTn
no9Tow8Ag6cahunY4jty+yFXs+U5vkeqilZ1NDihEK1CrzzXigrqTn6qLGiG
CcjmT1TMeOIapGRhdZFPLPi808GbR+XcijD7M3yn268iX3in2bWOaikcPweE
VfNRbBNjefdcHESjEDnNZyFShryR87i8VucRrs/pDYKieGKga1qyIatBhTvQ
bFEuOADDVquMVEpp6LPZGockLz9helNEg1cvc4BGS9CPOfOfAYqVvC9q/Okq
Hk3p5Yz7o0PNmFv/DY2QrO6pA/ip4e4OCfZtjZ8M2opGWnCeaH49DnswirIP
W9jFt0u29qgMOxF43rzXz/CgpN/cGTasi8nuF+MMjpWnlHXVX7Fxp7B6/0V/
gnxCG1+8omyt1M9NeW9G6pjO69olb/7kW7hkLcSUMvOghSv0rwTug+jgA+Ll
bZ3kj9nd8oooxtV8H29GsZUAwE4W0Vq8Kf/5dqamgr1RIL/pn3Nwz72UO/VR
xUX1FIV6we50Uay53CmUe2HQp8U7Uly+2Taa35Jm6AV+46GU7tSP0+592kuo
azpgnPz3ZdGgYD50Q2vckg/Ukf2iS3NoEh4EVfEAw5IqkqYElE470+Q3A/2B
9qtFCojrCvzWKFINR+e2L4KT43xngjZnYniOXESC2zXlyQq3/IEAaz/FXWCl
ErDSO3Da4DHfVnYLE4TxpEy4dszS4FYxhx6trcNLHULNjxK1KyKM1VnefMvz
hPbLvqmmlodcxZhSmD33JK7rFSdeeaHXs59ZHHAK2YATjVGm+2CLIv9BWXKv
x3/SKYJJEdmWlRWAtC3liSyPA7Z6GSUSb5HEjNdROd9OANRhcr0KzkJA3qKv
PoDyiNE4Ilqc9x7S/Gy+E/TVKo9qw5I7qOp3K2s7lOYdnY6wfzfPo+Lv7P1C
cebO9zs6vDX83I/pOntfCUkna68O+MDRyH5WheYJFBxndApklRIA9qv/RmNZ
dcvGiePlG8eGMVBQ7Yo4AOaVNZhSJcC6ZLug3eHTt9vj8SZFKyZpwn9CMS/J
zioPU8fHbP5KydkEc/ba8FPiQdjF/js15VoQvkXVcgppqsjGdX5j1LEypmin
Kg/F3HQFabh7E5B0Ijl1rgGCn6rL0MXm1hMentSIggau1sBiunlXf57N21f5
bGTAWJv7VBYLaFC23LCXWabgneO+r2OIBZJuw2j9WNAtdqNEmrLVxy8MrJVu
Risc/G7zlzpPgpVLBpiWb1DjwhzcwQL2QJ/YBIfnOw7CJFvq48Lni1958KGW
WwIWwGfU5TJky1Sy+X6TrlTzy7+ZL+9daMQDKg/d7r2m4AU91PtQ1xdCD0Ae
aKOjUw8fZZSkb2PEi3YrvPczi/WScZcUciS5seOZEjzHfA+kThWFGCToNZSH
4h8/EP90xlv41TusWiS7MVYeOFIdrRIsOnZkKAmegc2ux4a/TukFbtvAdhXS
Yx2wKTF29dmY3Ej0DeGe9oSw6/Y2Nqm+4Nmz/eD16Qy6G21Gfk5C4y88ocbV
hx2QyuhESIGh2AS3E9HKugl2RY5Sd0pwwC8U+cN78AgWebWc1cxDsTogjMR3
dtCAoBeouv43lrxrnD4cHjefXYCkUAtVspYZK0ERykJPo/mI1jYzBpeQbL66
RMpt3C2mN62ZT8vZiJTkK+6jbgcui9XS639fsyrwiDTx5xXzM47se9tlMkkE
7Inl+Zhadtdfgl15dO4ulIdsoDbWQhzj+8+tE7sEPdhrxeg8gyvDVdOLTg8X
uDTIoXcBOT289Bh9/T1f31KHQgGZIkSbD+9Tpl1G+d9JkBMGPxi4KmeyHfDY
UiJph5I+5ShEHIhspABmXg4qTO+inkkqD/wFHmIeduRr9uOEV158/frb8Atz
MnRbOSHvGv8GkHH09aKpSQiXhp936e/4kCYeVghThlbk9+8fiIwbKmxD7eve
5EWlmWMAk4M38yUnf15ZeGQ7RtXzsbWf01ciqqTuQdJ0R13D2gxSepPtTda6
vSC/Uws+QXCKNVK6wN/Wa2zmb4QMHyV9L53zmGb+NfW/Cdq1QulFKi7Tn19Q
lU5AYTknaouRC34EX3uUhLZROBZfx9khXs4fbOl+7q/ikFmivWUVWQRcpYRc
Jd5bIWYOmtto/zCjzAqtksqfoDzM7q0u4ZFgXTvUXajTlQRmXXHazkLUJnV6
kQaZX/Usu/qXMXimoMHo5A85lT/SpKkWszGUu47snwXm5fJ6vAOnTvzhZ9+1
EpB0LFLEJRNZhOmOiWqsGphO4qBf02ApE1KYyMKvvbjTWuf80R63qhdr3i0G
U9IbtbeP9XUG74WEsW4MmEhpRuix1Q1flniVsDKPc+hcwzPJbSwrKGbKh42a
H1+R6uAiOBgzMFyNMwI5oB4cAm/X4UeaIYl1z8urp+5FClwpR/PFQRFTIFxD
KWeEWJioCEpxRcKHlJqZD91bKxMgkUh60aZu3cy05Wmp1HUyxJ7UYNwK13H3
wLIksNwqT3XKarxt0IJHRFAWbfd2grm8ZwGjxutWlVr+de/dIi54BNaiErYd
NXzyX5o5/P+/6f7+mg1O2ErgNO23wOtpVw8xD+1Y4YLQ7cS/Y3AryT35Lvni
1Jz6hEr6RpCKlF6toOgWdRpGBJBp5SGToE8LhF4hWplMSiF1mkkhxh8RHmCx
9qyJXsqhgu0YX4dTqGN7Ci1Tb4B0YsIflHC6tQcrg9oDVzLkm4DUs/IWMBou
w32Uhfae90uNws2wy17CK/h529HNmcirlxEY2KZvokgFc6mNSxmyxy9Bl5Qo
fALfdQ4Sp6m9z4hjtdF0xHi45RaMbMbQTntUciy+rOQR5+2umBPFNWHkpveQ
13w/VuA91NVSdUPCcw1bLPgbUCz+kyC0zTMtaDCOmkmnLt7K+EOt1nCXpQ9X
dZYSt4Ce9pw/PWKFUB4kpFiIp4IdZAEkPlE4PEyyhrxj2ZniQBYtWUi9C1PX
GFEJiQoGObB1H70D6U7gdYjj8E+zVfKO7507rrrTprR361/mE62JUsNEtE4G
sSvbawSGQPJxGsbvtGkZt3KZJksq8Vrh5Y7E8BAJjA2TkUHDDnT2Y/FowWxU
A90542rFmnfk23pDLQ2tAK2vbj/ABOB4nVfvjOldIMqyGvQxIHcRpsMW54bv
W3Fq1kgzQccEC853F9x4NLmsX19hTCxcSXV/5Z4nB3bFEEdwWP+GW6K7xduY
16e28RACNbqqSoohTrS5OUC99JYjYXoZTiRpNwFKalZ5TTzXIXz7j7maXufd
b595GGztPxlxEnHJKFa0q561SJ7dOMx1Qv9En5d/T/7clQ6DzKeyYDZZobPI
ClGpPHF+0bvQxeTio34XtSEh94tEMHcZftznrpW0Yew1t0+cUkeX3FHrZd2R
k/PCfZmTEFEcorHf/AZxXrkQzxUAuWGKRlFqfsH98Zc5mtKRgz0hXHvpAIhl
YaAfOIc1zwRR9ZbA9JADbotFCTTATuKUaBZpo4JVLz63hqgWbIE1Zqfjd6v3
REgQLwaGz4zBungTKYEsg02Ioyx0EUAOYwbMxawCrpPeUgot1aSNtU1b2VNN
g4vRY/Rr3fi9IFNf8TiScwJM803sAptNp/BvFIg1FlKnN8FClUD1ZDnIHu3p
Bc/Kd8oqEJfzVBwyENHWKg886kudBIszKV138Ry/x7WK6m8CqWuXXbbhv8pP
nwTkDm6CH4LSc2omMO6gBa530FrxobeSFovg3CUIpdHHc3tTUHJbY8zBdooo
Ld4Gp+wMhvfobfCfx2orOmUIPesEF4vspYkqaX2rPXFTHsWmBNsxuWHOkMzy
7GG3jMyidLbC8zawdAu53RUojhY1dliP9/KdAUTDx+sdYShjUsh+cAZ6LXNn
sb8jORxwf3LXDBXM8LPO7cFEosqqTSfLp2uPZfLsTx2DApfuZ9FOzd98Dw1q
aAoLjBd+mwSJ6nMFbEjxtP0JXe6TJQkBn+RaKtHbLD8GBBBH3b9kejL46M+W
DOgZMEuQZfuFIih+uSwOrN9XvVOQqlrKfzJouuS+pQwmmk5PbBTfB0xgMhJV
P0x8ww34FDYooQCZCAteGmz0b4Oh473Vk5zhL3f90kDJv8QrM4IiPj2IvuM0
+BiXMgbjrwJcdpu4K0VlfKiJKBD1qSg/E7kXbKRsa+RcfWl2GnIJnZp8EjEf
18PyBmEia0UgRDtVyWrgEgGvo3qlUrqUlf/7IDxFoz+OI35YeFB5KSZu/MTl
j/D9Jcs454GcwuIb/vDQCNFLydmxqplpOXB6gbVQm9yCAhuyKGBIO3hI+dR6
jOKDQ3gmUQG1v1R3xcA/dB5FlIsKSv+B5NjDnfKsC2n49enHUULI5xbbY++r
Xr8GbzrjPpGzTelyQnRDOdja5FS9M4SRsrWaYQRACdGMVujgSEEjp2SNkD3X
n/NRGe7yenYybx7Q1Y5eoX7EX2RN4zMsVbCY//pPRHZK3VP14r+3L5vvAEaK
T2x5W6l+9k5fodg0pTG+xBjGpggXZdMU/INVaururzBtBPIUhz0o7kbW4QII
HGk5i4itD7cuUCKhWpLutcagyQkB+l6ahQ0B1ZvlCuvipOPRj+Bq43Wihkib
4H1P2UXn6XrX5EZto7bbKdoscQkuqcqi0LZwgF1xzNQwVskdEB8soVfoOE6D
F7UUrGye1NnhvUKn3645fVGQf0xesHH9moXcrpprAzENOkg0VqZw+EjhbbhN
ZxmN8rB+pqKIaHeGppRWzbf7PEpwLrAmCwsKm5T+ZGxRyjRwnxqjvLiqu/r1
m3XLlyVBYPD8H0K6ft3u3sKQ0c0uhODBSA3lAUoiTR8BCPUd+zXvArn+Rom2
JkkV4vhuAvNVbNrNy99/+18AxN2RAzryr8L+M1yZja0iND05GaiSKF8/SGbs
b9k+V8HuKgJLZ9KafPXCupSQpG9dIcVQNylGzBufwc0aDFbo0ytyJK8CtIfQ
x4n5DvQJh5mZ+BPypXSsZeGZhfpRX+VdV2gfxkt13pE+racPBXTpvCf+ZbYH
b+Grhv7LKJ4P0fmchv2qkc2u6vd348SNo7/1tczaP1ZwHG+BDLeco5GnWMEP
GQW55YnPkaY651NqH3pQUuwQ7YoecOCDVrCeZ8sYFDyuGj1LA6Mxdkue1TxI
daEDwW7nr10iysKi+aa8Sc/0ZojrCP4MAy2D0TfBKQmNmRYxzOqjJyOPXutj
r6Jhwr/FW118O6Xt+xY+KoU/5dtr27DirYJpNigFQzmzoADADqUBiL47B3vU
jzijdY6Ot5/mHh+PpfGkjUXApVqCxAhe/qfuJXzjO41yXAV05vxJk2GfkrBB
iZpC/Sakn5XuHec2p2IqAxD0wStQV9jW4EMyoIyl3IF41yBSem61jXiAItVz
BUFJO8wHW2aLXeUjGyqjNkgYVjZbcHaCCYFU3zUfH4jmc5d+ia3VB7EiF1r0
91j41i3yHUErA27aKnn49kdPUQANRR9fbORTjbJS/UIu9Zf7BjhFk98fhPqG
Ui8ufUZuyGpVzY751O7AspY2rIf5P4mzGEggmpDtYyvF9unKSU2VULD1UNGJ
CUzfCqS4YZIQdY6ckwCcOPkJ4vihoxvUZIwX7haz2aG3Hfs49TZ5aq3NcQV/
UNGhDplLTdNr2c5FYFTnzsDu6Opr72BVbipItxcSzg7j+gZ2vWM+sHndZeML
YIcSAUrdoH5TUoTA6xVbfFqy7AhEDuYXDh2OMv7nJoGb5fNqvyi1s6VGC31k
+itxHvZ0ADZfrpaYfJQp6Sh+ZcMgEXWjxwkDDVLrrUxnTZWbMBVoLWPPioxY
lbwPyPC+kqYGwfOIy33KT6qpGErA1Jn58fJ/smMSEzVzIMSXAbIM4+DRfwjq
XZbRIV29Sv1CyS+my5YyKUXAaSYeZK/hE1KxQReZOTcqBTBp3DR+6G8+/XnH
9O4d0d/lFbpvGJnvM5kHeHrocY7YByRgFbdostyHw4c7BNncA153li/QPl5p
lyEIkTT1cGIm4H5BRvIgjGP1Ug8P8PMiNMnFDAvaD/sWR/zP4uFTksSIU+39
14YvuFAlKzh9PX3Sw1hAhvhQberlyITbcUisWG86k0+c7kKup6FElfcsRYQ5
ql6e5Sm5lWGoFDLiiGQDmL/MgTZklvbh2lhTlEGn6XnUKfm8n8ZRjxF2gGep
QRFGOPm4gOMUsC7JNNFHypHfD6XpGaBTR6fAzKIbiLSuEcsaV4empokePj7w
ea04j3p9XRX/5fDRglB6HbLNLLuUSsMI0ytTX0wHDmENWLw/kGpeFzvGTtoe
DxiEsHf1dEJdrcx9W52taIKoBBcQzZxa+K97zafZGSz4Pcc5K11Yga5sm5Df
gnfycvhNpAW0QgWN+MEoj26qU6aij0HDvJEEw4uw9Y5WCohLac3Yiu/SUjwK
+um2TBvd5UnGxcEObXwh6yGGgHn180lCj5tDHFpf7dU8FS74RK3s6VLhP1h3
bYq7rkbm0b9PyQ4WNHyTWSQF7im2gwRIT1Cdeoi+wc4zM6bsKLrghBjrurRT
v41h/TF+/bgVTUBqKDlEPOGypWFm3hOA6bbHqukwosnlSk6I1scPurw/AHMq
z5L4VOJ0VwQ5KoftxPziZjkxA0WDE95U/k814JTISyVmaQMSPj1CmvegjSXP
dp9c/+U9Thugtkwxh+Bk0lz8ZyLEFI/DhERkW0qHChYND9voEqqqrG6fSDsQ
si0UCOP5tPSUyPTbZgn+ZFD2CL2GJgHt6W/HLJRgd/oI9f5GbYdSFse7Ta5r
08hjgbMJ+//pRg4LmyHyZt00PO4XL0qb+oqTh3v8nVrAldkUvLxg2wyJKYbe
zuC4kvKG8CGy6aGxUX8Pmri4F6+WMLskksf4MF786h0qr1P5MoCWakH5iViA
DAwQCDGCLwKw4G9MFYtq6SzTZsi8DJr2ZGIJ3mDfIiA4rLY6r9vqvGg3rBfQ
qXEOfw3Vk4mn6VYeaNDKOJPhjwWoDAOEZLbH0K9VPj/a8COIfF3vhTbFlA60
uqdZ9OhDxwRhKrHjpLXuWDzTHJ/wStYNbm06IsiKIxchaHaunXgDnewp3l8V
/Ee0GG5ng2QMiEKELPPf3hZXfQ+H6nAtLllgM6Em1KMjNT20l9B5A/hxL3I3
Eo1l+HA4yVGzqgXoLgx+cTTa+HSUQDzhppWmWtAA95N5bXNwXp2wdqDfJsyW
U8wPIFVI28fBHiB86OQ48Fqq6oVKLWw2tcuBASYfJo44c85sZl2Bl6jHbG4Y
wedMU3dzmNv6zgQ9zLhoNoatojZorvj/r9ZzbqRCs2hwFq9Ozhr/H7sLmYYj
N4UxYfwBfu10j1rsAq324l8NxVo1fbpefZWW8v4Pw8U7QLVWccKvw7sTqYSu
IGJ7iutwj8wgcsFJhNSLAij/CJr0wqxrM6Rfw1L6Pgj/+tGGmshAYiW4/Peu
c2r0IPsz9tRB6Cv9dEy2r6TLFX93nk5R+Re4+vpU7uuI63Pv91i7EbtAltsS
jpJ8DpmUXYqgYVyGqA/XMWhk9KVjBF0rn1Y4moTOKYy9GxE3H8WHX2p1SAOM
MkCemwI7Jaj6WGTs/EBP/qrRYPXgx7lGr6lT6aGeVMLXEshxz0ByJW0LHPKQ
gLyJUH9Tzr5RjhoNmC1Issj8H6C2e3H3ijcXcJFeaN7mcv3+78g8FpJ8eC0b
ZwSHTHi7Cide6tlEf9BCNEX1FVvURIvZYYX1Qn95ow6pu6sZStSn3MWrj9NX
m2L72daXrc5QDjain0RiN9Uh4o/FtXQCIebJNpYbUn+kB8ZqjMovdZYdxMFV
8NWkZ5yqdSm+Ksg7xhp9Ylio2dLo+2nclUgy7sjY2lO8h8jWNc9fY0pfoDJI
zIt1IgUTpE9P/dERP7nlQXfRzchQl8Vg3aMUY4cEIlFIcTbluQSu645xvyAc
29V4ERTpGrIqGGW+cJ+447k7SaXgBcqUD7LOnu2gmMmMQcnugUdihhs+YY2N
lIoxVy1E9qM0dqoH95CDFEv5P9NRV9lNjdNfkoUBtx+M86Vb+6BlCPl1AmhL
MrJRVWes/lQ59RJilpLjWNSFErmOO6VPQWd3fE069ZmfiFSKJ8rOidA8qfWv
XDE0oWWlB84GK8AeavelYNv3Mfhhle0RktFC1dWT0Gtp+GY/QnvhfojTEcdn
V/GzLx7rYiebRV7D3eU8Hu+8uRhYNlWXbYB8Ly4cdFqUsu2sS5jYxSl9Hbh/
0HsR1DBl5He4zLALTTUnEJWCOxDtVHWuiwWz3ajc2NlD3oOAtgGNBDXhMOED
oMdb/cLFDtktrvhypceFFZmyaxGZdPo0RcjTvaGIeiiaCYVFS1Fy75e/a5Fv
EelxFG7AwaQXkaxmJ1x49TTR6S+DZUp5/3Hxtj0vXJASuqB/KXZhlWROs/Qi
AopSZXorRnMF7qAlMuscGebZIjEcjnL6QNsXQsdW+ESmQCLGiX+0TyDvhBgm
LigRU4uMRthfTnDWqrI3O7PI2+16EGA5rX2MzZba2ebMBHQ3IbwxFHSs7rR0
dXqtFUf5Q/mx3MvhnNrYfTxPGBnAmHZKhOCiLZt2J9AW4JsBLdl76vdxr13w
R8m+sQGOCf0CoKHC464BJEoqNIEuXhFm9I3kYZRuTyIy6u7IloCJ/MD/I6Ga
ndGIICbLNzeGAyLIOPJFmbNWSd1CPIDVlhAghxCLHglKCtyXuhxHk5aIrMIi
m2ZFzuA8+/M6EMa7yROEOPDTeaOvY4OMpvVNPC8P6mg6hWlsoWSbzWyhKgpP
KcsZrHIO370o9P+g2LfLrQYFNo3bLYX8ilqbJc1Lugos2KAs85mtfIXPEuFx
qz3Z+c0oXNI2orF4fPRHW+V/gYufCHmy79My0xDo0ZKLske91FC2dXJ7wRYM
4Zr5uEHhTzXG74Q2fhGkzH8wmkjN1V4+nQBEHj9xBcvmf9Q0XMuSRPbXygPX
o7j0kdNW4zE3SRN8HzeIRApMbvKqennyl1xjP8ZRwjlZIC5gSryTdbF377Fn
Gry8F1xAo1DSbKp9PpfC7X8UUpUM474BeKqWVC1nr3vzJuplDGa/h90/uHyx
/dtOw6fGxv6QOhuR8VWd3oBWZ7Cev3h290UhXLxD57gc7wGVpTB8RjYQvk5N
McVMOfCGpM4u+yUXDONHOgF3Yhne/b9tVUtGllFYzPqBRHB0nstGuP8ulXPT
GcTViw3xItvYDK/JQC0h2xVxpB26VH0/YhYGb+xItYm5TzTRymH2IqNDcFhJ
JhUx2AbR5p9kcmzLbPhhQ1sDz7QGp55SGz0ceBtsrYY4m7AMQ2vanyf5t45i
HjzKDDZKg1dmgICacCMywMYtWfobYsnCm+duXsLDQKE4nZZCChutXNnTUCyS
l3I6BTjfUTgLqXeysJ9mWu5iuWTsTrvIssQyOpstyABEotCV5bg3KIL8c7Jc
Fnp6UEbuo9sdjR/ZMTX6wX8EfNyGQlzXkFuJw7iz1yRM5ezqogcwlq1pPyW9
jClab3LZtNenFjCZXrZgY7kmre7GO+xQhKzpq3rXkIgo/BMur4mrWSNkR5Mh
DbpztR36U2B+y2VhaJHwiYWFe3QazC+ijotwAJVw4FVMpsYkH3zOEGQSr9n5
r1YyXXY5iO/+k1UA8YFLzMSBxeMEHaEnAVLzFOu3ZVQuN4Wc1J78Tgk49vs6
lowYdb+lLX7HFsW02c7697jQe8dBdrs3PpkJm43eWnL25liaPiRGQBpyjAMF
rxaycEvOC874AxpxqBEvuP/So1M0RyLTXbFXvjW22m19OOCmqwrHL8yT/aLG
RxaT0qvdW8Fm/MBxWLyA2p4ImcGc6MDIWqlYcIXfjfLZCQUdEqz4i8gHcjEG
bjPOLuk4xIIylBU4f8Lb2FkvAxxffOdoe3edj/BCmzNNUWetYFqrGHAd0d9x
FYH3UbEGy5zuGGS5oKY1Wy0o0rh1tIT8MUM2sJTm54AE0VzEvVGIUK44yWjR
L9FZbs9wdxRRTFEQITPRih7s7A1sVB1hp7huMh+ZGFlHNMTmxfC0mo4XSEJt
Kc+mT07J4ibi5wKd1/JvbSZVTy/N5warPORTYNA36FgnYKsgPtq95pbEbjW7
9wwvc74FlL8mUs5uGCQLXF9KeeErzLnPKjgr6QfV/Z6iaKCDPVzQXLG866XR
KKaa8E1/7W3H2uOUmJNjfosvhDFIoS6qBrTKL1+HA2HB9p/jmCHkPPB8ZZIi
p9+1YiShP+AOFLEQu9FmFPwVNBLtJ6fkj/rs7nI6ID9oWX8SY3+OwjY7wbYb
O+n4KurzlHsezfrAVQShf/1szdFfNKwsvT5aZBdQZENk77+QAQSyv4iF57dJ
ommqKGT3VWiqlqNkSEAdBMmKSCFUfPf7WdiSB5wNeTJGbYMTguo3mJh/ex7K
x5/RE/z32laB7t8CD5uBg6nwlyx72UHHp7C4A6NvY5SmxgZ/UQY5WnwIEYsA
a3LTENco5KfclCsgAMFfcJye/4eNPFij5VB8Oo16P5xfVzXuqSNqpdyOS++i
gLT4Vq8rKu8Gm2yV6Mc/UyTKVwsjSW/sMaVCLkWYdvFd9l7Lb5m1SVTofk1n
+DzRZRZ5L52jucM5MBlNMxbVeCv03cHdbT58jzmBmG18M7Buuvce9xt9qdOx
dnLbadA4Pyn4XFtUAxls/O190bRFVxvw+MWOYjOQu6FR5WThFz4viFh1Zp9P
ExVcOeFCyecrYnhCUZuDibXmKxguV8ocj9BaNvHk+xdf+B4swohSK60BPu9D
TZA19HeU5CbcSFxgYHADvyvFZABAINB/OvAD4HEeoZLc9rLT0BvJFoEBrz8U
AFeWdR+hzrVuB9VluBXSePOeko5B3rUKkj6p0JxaJikr/6ZeObkzQYmaUZUh
6vS6gGOw7rpnEjrfYgHBUXLWJcFVOfHAkq+LZG6EgGPeuUWBZPLeRuVZA2nV
AiIIRkY/KERVEE1/ZhJf6NBk9ZcnmaDjDibi5YUPtvVyJfeKWLX3vKns5jUL
nxn2t7OaZeTVEVJ4v6NcBImP06GxmlFooCbMqvvEwqh27mZ3731n7cYxnZ44
P9nR8+f4u/y+wcw5GRPzcGLz2pG9GNICwRK33IoaTr48QjSb30mM5FvgtmRT
8OuSW7ETkOqUGMLdyHmrfvialWgRvOnypoIFWo7o59Yhc8348d/qAWLPUQSv
QT6WEjTuYlaJNj0NT84tMsHpz+KywURIySTWnHfOnfogoU4F8Qx1vAsSw4Xc
paeZIxTLrqgUQGj4YMXE6Vm0l9eJ6tqLK6gwxgJqtkJP2spTTa0+U3K1W/qS
tX03bbtAJzPI+aP6lKTG1P6vtaNSF5I+sR2Kp+won4lQ/PzJT2xT0toZRRIa
adg7coSdkuTJ/cRdn2BwwbIsIP0v64Igf/GJg//Y5IAomJlHzT7A5XI3CuVM
pOgo/S3NDv+RpOYub+u4OD8xqNQUBR91FNvOwnLPbcx4q5y1qLjEWka+p5ew
9+uqzNu2ey3yPYlTVxnzMb1QNjnnuS6PhHU7zthFPJD/dPzD4+7XOpBJcIRW
zE7CgZDMtMpI0FLiP0esku9oAOX1Yp8FXS4zQOzpyTEmF+5RZedr6xfE6oUf
StLxq7e/um55m2/+mt+9fkznDlpn+EX1gD9CT8A0/7kLv8bMV0Pa0KZ0jsU5
PWmW/0cugPiRD+4FRhv1CGh8ghIpJUPpPyz1oxdt7P3o6idVs6CInvnRCOMl
6NoNyTTx8G/4wgVnqHE4yxN4S5CTYtEnygrhbXg22zKDLYlxvWD88bmSUQOn
uAtohepL0e328S2429O6uGKv84LsJMFMBqDzUIHRzHMRa5WEf8g+0eyIemv6
URLzX92a2qWJBSy73cSfdtLchPC+98PFgpv0TmbrAMnJGFalMWrzAtFcpJmw
F0rc/2aekjAs3IQfrk6K6UGQ/n2ALxabkrOxjxPXw6qUez4+xUlAf1IJ2pPw
+yboWZR1aErGroOxIi64CM81xuHG1rXvUWFba+z7Qk9PXEnzo2rAMKn30UoO
n4daN1K0DA/qelAN2Ir2cQfwqlXWN7yJvYQJXUaw48xwAQuw40+ahQpebAQY
X5qMhHfecDarJDW14TR+rU5+4QobkldY3dRo+3ivdy7lnrQpxH550v7H/uNk
Y5z+zol5yqx9ujD1bsdW4aPFSwltQwddhD5YImVmNRASBtAGiY0nIwJQo/62
uUTCzvjn7Zqfhiw//kXV45GEoxtigIZgXj5lVnBNDuOVrB5MslCj189m1tar
E0unE5oYec4qQ7EVS5nI/XpoUH3pbsCZdHgwqQXi5rDCwSE1nbgmN944Bh6J
yG06c6tdo3KjVlFcIBgjU/HkvB1i9zlV1+Xki4D6j7HuAZUd2BOPAgj2plz7
mqBcyvb8/whluSHzoQpetc6aLaTzMpj1YWjWAlZEoRnAMlVNW2SUe9LLcus6
EBWaG1X/t4yrD8uLVLlxl4NGJIva/SEMOBGEtrmGBOSIOq7JjI2S/OoeVsNf
jvepIygCYttoVgw0uoslPkx76jDV0U7IGtveWtIroRpyzwFvWm2iiQM7p3k0
6OeLTJUIM2mpHdzgb6UcCiM/9+dsPw4L/1zSx0uVwZ0fl3NTd52UrzzyoMoG
k3pnu5rSwXijC0uPK06Pw1KW7FnMCVB7FaCbywBKwzCKq5s/VGbR18KYFrzv
BGcyIRVY8OiNXBO44Z/Uan9Au+HvovqztlkuXHd8Cwhu7Hz4Qxw8tBQ2k0GI
TpGcLYO+XoJgqQqpnFvhwOhTLP6nJbGjm5xlU4UY+CC9bSv8llGT0Evt8VaU
VpbmuENCu5/bIuC6yz5CqmXooVAQUnSOAoajo/7dQtrLyKBwy9W+69fya8X6
Fciw+zA3fFuSAgzzCIIU0Yq7shfd1o4BYLptks7PRHZFueuL5Xv96XfhDYj3
ZNERbx5fSMfU+1lGGVKiPEL1yRfZDodyMts42MojO0tk+DCHf3gYxO3woY+6
b2YeLMk71eceCzikCRmjiaaqSYcFGiJyZOfFd6ds/jNIO/MSnHBEvZvWiW67
e2noF8UQ50/b4l8m5MRkSQisCLAUxXvx8vX31yXuPs2da7bqMIYY2wYYgh/E
IRg1pWnXux1oAfo9Ma5paH5PBwfL4psOt/3LtcIL9UbLvnhM0R80KqXpypDc
LUEVGJ+2NIFoS0cWHcJ+wvCpP+ibx3Gky9/kmpJTSZl7SqMvlmPNmfFqOAMY
YIn+ruczl2I8I+5mvFO4EZEl9Uc4lqcXOtsPslN92mSKzkU3txAi8MtO4w67
1h0GweuRlAd0rqz66ybThWZH4QtX723d8GiT6HL1xmeVNAfON2kcThBdFO1u
Q+XXfODtMKO0UTKFKnf8Pdillz1KZYBEVnSGr/1jKdoI0XoMOBZQi8iXD/OQ
TUwbuaKxDph46isGE6R6fUQH4b6QOGVBaxoJNJtm8ujlBOERb4cbEwpvCdAC
ASCiMJUjXGkoHLBVXHHEki3nxfYmB6Cd1bIdIUYVQAPZyLrouwUNU4+qV5LA
4YJZb13b434bmjGuXxLUHB5RFcHN5zz7DPrAlIP1rxnHyn/sCf1URRznn+aG
QZ4BGmFBKTii7jXR/HWiB5TWLg3ru+fIl6XQZhQ3KTytkAqjjlZPeqjFYUIZ
B1q1zl9h6cRfv/BDGkLIiua5hScROkz4PxwPtG6DV/bctyPSgUU0OysowAQw
rFhDdxF3CtpO26uWSrKShhmeX2lrkUh50iXfDhSdUJWe0WJtLxzMirVY0NLg
PWcLa4UY7CTi7l5YUeXXHEtxSRuOvHr6jsz4kEpscho9SKk+j3D0XEKolmpl
VoFC2KeX33mKOX3Pq70/LJANzXL1q/3C30X7IPsIAQFOI8LTkiBssYyZLDS5
iTpUe7X/zFyG4skSgQI4mgYET/d+LfPlwD7T+wOf+sa1Ep5GcWMn66ciEs4E
fcuJD6ZQeBsEnzQ7RVckV9wMEK5aLU8YmkIMsvi4giJIFKgpSYvtPYAcnsX0
52cyFP8CShvvi5QxkHHWw6crZxaM2hJ6+gJKgD4UTVuUXwmNSQKM4ePQ8j1K
kFeQU2syvJPVf/isYAj4lX+lzMbWh3HiKEJsmj3oVSljKvhNY8Lllkv20Xhh
GAy+c6XA11DF3yzAq4I+t3gzTzvQDGxS2jbbhzgmY44fMl+1PnN1cs5FPV/s
trl0RX7PK/yZHpE2QoSs1Eg/z6e8eZyD4FFLSIhGW+MJGoeDHhSqj37go00Y
n/GT+bSXjUCoYKRYdZKTpZFDSFpWuKd2mUp9+Sh8EsHLpSoJq5rQpd95xR6K
pKy1I4DqGWpKHuCvzlhJztlNXjdX8BDbz1M9Ow8hB0Ko49aDpVsMChXbCtwC
1IO8cIb7mW8l/CYIsp0tYfZj8ERLc08CZ6+Ja3eK41kdmwaBBwd+xbxjQddC
pfTOKR7ITpLEhADBkPPveGWkCKY1CR44chY6wpJEYbi26W/NWS0qej3Ux3Tg
IZEjqg4Bs1nBOsYCwG9VFTFa9kxMJsaqyPX+2m7LNFT37Cz5amZZ/Dpk/NvT
PDtzMekRIt+i4BeFOeiXPC9zeFLh7hIXDft+Hd6yKa+9fqZBvJxe6cRdab7P
MDX6cUxLrM4kopsdWsX8JAUvmSBgDbwgSJTKM6OsxPzrw+u1zwsEmKRHTfhc
SRDTI77TNL2H/PadQAIr1zK7WM2dUFOrypgB0e6YWZXsFSlyOWLboig9YH5J
UKJkIpOS7chBYx8lQGxbNxCcWP10RzZiLsaZIJJtB7HWhrIZP6Djp8TQBj2n
YxSB7eCvZf4UBrGa6nHBR9hlevgVCeL+Ec6dlMtFYxfy7T/M5cUXim6wSNV9
YQlst7/UJvfR7pySG39POiniy7zKf4DGdARNIR1lMOPB/FvzIF8nPbo/AUGA
8fLTpXxheZLkvFS0e+h97eVNpYPDrZRiXsI/DagTolGpQDhrB+4eXGhktlha
1OFNAJx05iDwEsWdKFnEmelhLdKjEtdd1gFr6AekbCciENH/C7aye4CvkYdJ
YaYu0G/CEAR97rQzQ5v4/2vPa9VDpOZ03zD1BHx07dDYFUnYobX9J3BDN+jZ
88sv0E7vUC1LJheUU0k6Q2w9TyEb6qgqzsSo9JTFLh3um+ZyBU8MLYc9kwGf
V4mSyeHygrw5lBOxzyvAlOsyOKjZnVQR+2E+bt8a5CWDeI1vAIpjoeH6yPiy
k4rEIkNT9n03nTJkb0GsADv0cz1XnakwP1uLmJzHV3a9twJ1O0+ZWSfamTEZ
Wzxa9PsHBNrAW+TBKOue+xVKkOJ9oQeb8eB90fJUVIX2MjpQhg3nqMCEI7tz
HWDaSYCN4F8OL6wtMcHLYCA2l1Y7zba4eUPsv2+5zr2UKIAXpKulCSOYUmM4
leXUttFxjcZq21L1DTZoT6Fr0lQa4Qigd1GC+g6TgbiABpxQtIeDJhdxX3t9
1/g5HOtYTFAF+dzQY1xD6CuedqGKbxzYs9RUzE9YuIaqE8FkfMhmnwkUZl3l
g4RVh4tAxHljV8AMj71UEMFIwlnYckuESknLgQyl4WVBzZjYa2qCYOCbJxeW
YktIMn/2fl9UBiJH89y0l0hqQwLJc/MMJkRflBd/LGdwgqL8NuGY1TGjNr4J
AySCxdXJqJq3ZlrKZnfxJSFVLOb3sXufwxM3K938mgeVRoRMco+Ti4ufvh3L
SAY5FoASPsBmuJEE3axfJ1Gqehh/1iWCkr+EZa2zxgLBZQjW8zYpiUCe5Z3l
i4vk1DZ78LV1yLZ69+tS1Y7GVZn2kEU5cq7J1MWrbLemLuEOlPxxGbpNsMBV
d/U737iMpT7eyy7YVmOrhxI8cXQFKKgDEHv7VkrKwweiCoBWBqSweJcxcyME
v5cqB1cRvLcZ278uPTaY+6SUbBnXLFN7AUXYvvWFf3HaTtveT84OnfErmTOI
15/ANM4OPFmSGtMyDZIpfE2taxrhKyL3t3wINoN011yF+xYt+xbm3ymH9d8e
qH5ii5BFq7jN4AejklQCQeooqyjiWkZY98rWc7G5r0rgeJ0UdEk5lMPlvGgB
dEnizqYc4+jv3kBuoSpeJ17VI9KDummlPyarj2TNhisb+RWRFQeHoKBgDRwR
3nMp4coF9CpbDc/mDdB8MLlezbAztpS3yZCI5VZlfRtY1e834A8q663HUKzd
wENr67Sbt13lUQ4UxxNfpqefd6PHplqsAAhnFp70BsAPCGKRhm79trXAepuK
O7J4l9GT8t/73GHRMr+e7tf6GbNIHP3/z1ULOs6ELO8FZgd3NO6O/G+j7Dwp
NRlucCq45Czw10jfy1ujcX430PU3+sDupyMKfPGO7Ig8EAH4hmtA8tLtEaZN
/oAkIPFhH3W2x4o2hN2Xix6H+KCoLGsWNhcJ+YZH5xYBvHJSAt3Mb2n1eNYg
R9WJWEYlwuP1HLx4b5LiraATdSqJabYsgckhjXaFX8Lu7s24IrMXOcuhmXM9
Xv6IDmFAhUFGhmJ1Owv1xjwFSsT7irVaaA/qDvaPvVjn4dCtbQ9NSTpoJ9R8
XbCcNF4oZwSRJ4Uccc+FT2Hk3kPojFqASuWjHZwnhYwVrGK7+qGP2GXmSqvf
k2S3lkxNXI2dGp9mzj3TdW66Yase9vLEG1XpbTn9/c4UaBYkiX9bubrA/Hit
cj0U7cQvr/UInb/LclPay13QBJERWCaE+GVLzVaYgr6A8I3jE5EOXg3hqCmZ
eDHgEYVnuYZlyka3lvn0AvxQBfjkwI3p+xvbkV66ew1HdeZFjK/TOdo89KmJ
Kf4XinW5X7avhz8+vGYjlNXzGxoc/oqdQ+9BW3aswAN6B3I2SvCsNbVgOkVS
iArC8AkGH6/lVSoPhpWdCQFI5kmTJ8Vwr4B2O9kENvZXeSxSXc7OfrpnznE6
FWeVgOmeEDHPSignMF7aAHHMCSsnBw2tU/cfSWLw/6tUeop9iXBdZNMT31KI
ihsUWaXER8++QWdjnd8+yM95MIEB46prAKYC5i2/P8jD1hoCxS6sFGPRhHDz
EZr9MLCp7L6waefVJn5Z9O6hYnmI0aS4kg2fd889/xBRUOD8bnD5MssCD1AU
Pe6/cCEJHKSyL5wYc1FlbGJrgXEiPr+1KVn0BgMtgaAgiF2GCcLEYF7TCbQT
rRqhsKxKVBGIk37LwfVUU98exvxq+f3Ps+FTsmvRUXX9Px2YxvBELFVx+IzK
BkajJxFvbfhHk/gNojeMVu7Jbty/eTstFP/rB6CAgMxPblNqD0gC4SiWMUzs
13EJCAbuRJOEsJPgCieIQek846Vbep4rWAWCx8GN7sq+SZl/tqjGv7dLuH9U
BTXcxD5oAI0p7Q+eNd+g5t6bLPd1v5+W9EXVkGpLC0m4VKYCAV0zlwcxc9Q9
L8Cifb/0eNyvGHmlYnnw4T90nddYI0yYnRcDc7jK2AyKUdQuky2w8WowFZOz
mDwgZT71C+C3P8x6lExvXBrZGQ0Vq4J1qixjVo2w9JuHSMeivdiO2AAOy36C
e8Hub4lG38bF4/YSMTs3M4eV/hKlcGE11D0pHFeyT0WefCP2PwTqAXv1RFcr
/kePP1d6bww/NbwlekrUMxWZXZ1tH9P37vSwQ8tz8nzD5ppcbiQhZnzHrcBA
wLjoCzcYJEzZ47hULJMK3ZYs1fYB1xf9fKRi4hZSrXCzSD9tnC2WXiNZGgY7
HwuPhB6u1yBgqqtWFOam++A7HJjDYBcxKihXLExrLnO7t8HLFBtvrYK5FjDh
vvUsofs1Mf3AHrxjXgj5wKGD4bQuKt+AjTn1bCcEDrwH8RdrnsXszUHxRMkI
y+Fsd2ZBQDUmVWb5IRgtsuoPKK5k+/XOgnhkYI3BFp9FXWBGIMHgcF4tvh/m
oAFIiSf+kpj2bGt1ZpE3esjmZlQzj4KfVoZ0ZuddFgfiQziU6fjeJBfMurZG
eQJYkqQR2OvmPyWH1moPm8F2X+eJuZ/sZWQEcBN+WuCoFfln0JRy6iVqWYpX
TTUfzM+4IdtQcAUxGsch1x7ENwLsvZLpzO/Ty+UC6O5dTeox7S5Psp7rpCoT
O1oIZP62nOV0CXxgta4sC7Om7xaftDZ9ivV/+76nbqlExRAOdwoOe37plmRU
RPaR7cJ20/XBQp0uqKFEwi+bk41rKbwUu4i8N1X9F0kJgZ128oiOJj3nc+9U
Cq6n1niX+M0AkhdQ5g0NdBPl3XsvEu6pzRe9WkgxlP/uN9fwFjRzL7+AZVSU
4EZ+dCiW+iJEEeJLzIg7IKI5jxuH3xjHp6ABj6n8nChmRrfzlGFT/j3XXBAh
Ssxd5YB9h0YYVaejzhSCQnsyM+Sk66+bDnC31Frnb2brvfEILEcoblmi9Wa3
3QQFoIfZqE6nEvcerCbxUadBmK1ZRktcx79EgM/cWmTcHrCOQjSOzka8nGRS
CSjvVF4pPdtKMU1Bo6E4OrduCuYkf3o3likB2iNNYdNyb1V4NScbfnnxo39/
c+eWmYKLrlZNFsasvSmhsEpkNaysK2lj17akIpdRQFY29Ndo5obpUhp0uTGY
9IkZUrCiWjqGMmd9vGqj8UV1vqUid8hA/kEmIHyslbE/P7AHCiGhr0mrA0Hn
ull1jQMYPRqNVm93AucdzQzp5g9i0nDZ2v0n/r/ImPvtG8ImdnfxAOFaXWbl
Q17XAe0hP4dw39I7rsuvMvmI05gBUHIATEOSxCBsE7qdv8wle3hWy8+YAjg3
UIwLv8S2voOwafFTAdC6/GtR3wK1uNxVA3RUR0v/CgrtmxDRCty940nmXOgX
OBUcOM64YUEe1HaCKRMSWpoPgqgLkwq/zcj+i4OBng8xvh1oF7+S55bEtBlK
f9PQiS+U8qe3sVOOUuLIBiC5nROnUlSgub9MjWsjgrkFhf1IsY5ZCbdkvxPJ
SiDt/+t2PXcFy7MojF4O9zyq/0lfUijZ/S6gWhiK6rjg3QFAydM/SAEn/OIJ
/ms/9BuRYibD+TqgZ5Uttj7U70Rs+RwQ94Q6hHz8tmH2BLm48FJMyyyQQg+H
vl5Q9SyakhkEGiwn/fm8bYssRbicIyr1qLT/S81+/QuJIgRUZB5vVTBO+DH3
qX8MUA0AXa/uxHp6GLrn8YvGYNdvH1xS2HAKcRwljHNfF+63te3UC+1Gatdc
YEzGoe4w+hyViuy1I7aBfFcaiKJ2SS/jT27Y4OYQv0PkM7TLo3y9/3g4Jshi
5oTKLbuG18H/osLC02T7NS+qqYv9hln8a0oChs94mSBn5nA+uYOYKO8qfah9
TRSO0Bu87b84jXEk7PeUkZCZV0ypp9SguzXYcaVgZyjxsnNHO8UdgtYYTZoA
X96wsDqzgL6qQ//rLt6lMshZU8BY6IESPVFBMJZP6kRjft49/SDbs8YPL7IW
FzPn7ggMqvz5kDC7twrUte73bvyB2gHYY6RflArBVV2riY2oExBwkseculx1
eZMIiw+SNB8FET6PjdkPaeg3vxkUcE1NVXulNtmF6+vzgvT0rKL2W2mDiF1n
r7dJ1DDgpdqqaatRxVgCdvxj+SIqQ9+laKKpU+Xen0YywgFSslBZLVq/GzwO
FKaOF+O+aqC606pmuvomSZRiTjX1fIIXXwlJe/kLl651LTBZKOYCWBwHXCtY
7gZ1jorQzqalN8lWuRLKuTrRkt7eKI3H/UnAgbTKc6GvqoX2Cz/DYohLlGBT
C/IS0PcKzaEk6JmLMXdB8TnI2SuX3ZeQXVYiDX8C12CF5IzHJUPrn7IIu9Wv
gvsaTmti4+yNMNLAid/PhtE3AX/K3so6eNkm6+PKUqik92RyIZew4D2j0V++
3bQCih8t+FJxrtJT0o5yHiI4lM7g30u1ScWOz+/D5rH2MItYcoaoqiGbZ8N9
gu5uFQ0aMJ9m9mnkUhDZkyg64gvGYOut6Xhk+CaP8OUIeLM6dsTWoU2U2AVK
PfnahDfFrXTKRmyKYj4/KpHu5tOq2mqnLd0lFeNFMag1C4kc62O77NH1V9+O
dkwGSFT+dqaboFqFDG0X2Ngm5sOwSfPOiucsf/ro42efx+KlgSJWujgBi6i9
waWdU3WXtDrE6h/Yg9t3KyLxATEiWouOk4VsqtxquZbM6SgE4mwe/xV45anI
rBFCs9ZpXRuwti34lQXqvUQ95gjGR1rvEpNyrdzytCARzhvhvT05jOrCUWT1
HJSJlwYZdZ439SdeAF2kr7UrikV32hqDHSoHCl7qihVztxtWt3l67MTwdy6J
A81Zx0GtBAJ1tIo27QCxmOGal/oeihEldPXrI1y90vRz9UWHf0+UAWjZZZ4Q
7ldaLtdVu1dicqtZXzSo/GBy+fe6+LE+lpsb+CNqYO0wgElwiI0zk0cjK2F+
UeLnOo3aj+OjQ15iyVvUlgNnEvqk4Fs9hn2bMeqXdBt+w3VXeWjQdOBLK+AQ
QU3RnKUtKNvwCn+dyj20pI7Dx2WVoRKAS0hQUck2yj1ennrBj/mwVAliruB9
nZ0oNuN6DGDm/2bQBtuEOV+hxAYcZBcosRXoDgsUPzjTABdVOl1wRDPIuR0q
pxmBUWUO453XfIYBnQ6sHEYoMib+DkKqO9p5GOB4DHbYN5NB/JiREtgBQEYA
FTXH2V5og++5qKQ4nm6feHIL6gk8lsEmKcF2ASxlWWBZa/XzTIlnaDllKyE7
KDa6BGnpmoefHVIOkN2eGp2N9HK/c3xKlvcNLwhYWHQt8iFSe/lZ8UT8N2eM
PGgXiIBAk24Pb6jz4BfS6Aj62ch6A/BrOY5JuTrMFFZQFKwifzXbFTpu55Mb
IuZGWaUdovcjJH2O/J+SIIwf96mvg3UA5IeOezQWMZMpMnII7zZ019EBtYYs
KdLY4nyx4AKGnCJgH1evrxNLSx9mXzwMqUMmP3L0udbMDhxq5K8NIttI+e/J
BLL1ijKT7RSOhcmfjA4hwu+3tXUV+76rpKuvxXze0LZMtudcJsEvzXw067Il
uXjYlRDT/9LzoC5uyMHsLTNuQZxlooUeBAvQnZvVzBTfAJDo2br5DsvZUpp3
fghVzw5n5WS/NjzzpJw83BW7vpgHsA+PJfP/fAy8X/T6YVJdRItUyIYbe+va
hzzhU9UwEqIQnNGFP4HLk/50ZUurDVSFcIuWjIwPVbUGukqk+YyzMzbLDBcC
vw0u4iZ0ZSDrqa+iJwJLCI2H5yn/JrdXK3RJcpWTvfXvf7RAwSExX3G5po6u
JO2VnVPpC3kwNEocNvDVSPshJVVnAEeLTzWtc3bVJtWF9KvrRwArGmfo9Tkc
IdKvc3i4ikNArr76gjEmddMPNh5hddNl3yRHOVKOBC1xLaUqDQt6TuYxEzDT
y0SBLfdXL2+DkQXJSePiARvtAg9Mp088IUWRLWmtoEC0n+l4ifGlXXX+KcIf
QX/bBnFa9Yo/8XGJ3wzJaBdYthqvXWhk6ro1caquGqERyZa78rTxGS1teKVs
kOYpNMwwFdoDXhuaSJU+FdEvLsJpAyq1JddPQzG4PhLG6rWFWhX4qPBv5fbG
16K7y2Me+01WL1D46egKl27e7WyqBo4S2WoMfxDxb5r5/GWWgVVogmewYk0U
iRc9UHl570AqNUmqaeUegzlS+Yco2CQKo1R0WUVPhkX7Hb683hlp5/BZZsU4
BtDVMeFGSZuC8zIPITakhSggE9bjj8GnPxndmN4g3yoNNz7+IoKW6lVblYNC
EZwZxegy2E88jLcDilo/vENpoRzB5/L1KuYBw22j07SsEBz6SsQGJFdPG0mi
oHCEc9sh8Z0sMoefum7w/HoBnkXPjAzerCH6EFWh6Z7xa5BsuGR18Z2/TYOl
dla8e6uch2CHTh8jdKNnTqu8Mi3Q/4rZaY7MjToXjazMyteC0TwOCPLIpmCU
WN59gdf2RDNTTJh7/n6j00N0izFiLveiSBfzKVuYG13Feh/PeZ5du2PkQK/f
eHq8VifAxfmBXfaXOp2cuUstj4P7FRVisCEAjgzmx4IgxfDe/XWqKkaNo9iv
qtRUCe6RSxRoa5PHPXXtbQZH/UirT90sfn/qJqsuOTI1peHzkRaCOYBUG+Sy
k6tECEspYsscBOikGW92T73/IrRW022rwrGsvUc/lXFJ8PoKPzZ54ggRKmFu
FR/3FrtckANNPRDlHQrWuan7c5c1Ug0hbLkmWOTgYO05fvGwhznmA4cV4wIt
iaYRJnXiD6MfXkX3vDg1+6xEFwFtxSpZHWls/objoX9fhfzagxwmb5WA/sPA
CoAVINSxIn0aGKcld7ZddscCBCT2Y9121BzjTEvCrVDmOtU77pPS0QrXnSkX
scT4KVwDCtiH/roXXMcirat/vuFsazemV+sdgk/7oO0iT9eJhMmfFFUwRvmW
ZHHazY9+TsfR6POnmIxpQmKNLyvpobtAGDASFGmMsnwJMrztUxxhtS8/nFa9
kWfA9ecsIP3/he/F5CX+eY3/ONZURCokrKt3Uin2cZwYvayeLXu/KEZ1xkWq
TBU4MxQqNOunw4PgZAs5TJoaZyxvWmE+QfI4Xyq1zEFf9OGDc4vy/gYHdCt4
aNEcIAL1qjEJYgLGOVYtu7eVuoGyR3uElbVUKoDInbapWG17SCyPzLblXhy4
oCkbA2UrBh69mdoBuOmnFSuvpt7ACcD8Vfts45dLt3rNhfgmiF5bSFzEygEv
ydNRM+6wvq0gQufaAj36ryida43ONjSQXV0wtJAryTsydBgVozhjKvaE0OCD
nmNeY3Y3lc1JvtDJStLsnWA8Hp2lEKBc6q2T8cHr5jUuGKvwCcv85DMFLl3E
KSbkKnJ5WTtGssNpHmUPpS6aGmFP6IDbGvW2pYtl2RmP7ilgU8tfftuyoBlw
pdZAJh/dxXXsw67/35iokPtTloTYyccKSG3GnQQsUUXuKInkw8GRZes8B8gV
eE6sbsaSHAI+kcjEJY+9Hpl1pbaVZRWpRjLiKYxnmmKv4/k6amloRePUfVzU
d3cw7OaYIuQSDa5OPzg9HTaL5SkcGayF0bsuWnVxTi6+DgES4k7PljWOGNjC
gK9i7jHhoUKmF+IqII/uVeAhrDb9JPo1gaPuX70ZaLBj9XiRoOrsBdcCaWHD
L9/Rzest1N1qG2nVk7yFdt+OCEdIWJhwOi/Hmc/E7GnXecsBH5K+YST9EaQk
7EpMMNJktIEytFQc+SdIc3FqwCvsUEzV8Pff48C8al6P9wELBFyPinfBQj2d
HwyEgdk8Z6Uy9BqND96T82FK4sMYVaECdGO7h36+RClb2fwPethk/w9kaSFz
CSQ9ysOCFT4U+Q5M3PgkBCvC7CzS/lP5XPx5yiG01dhIw4Kc912ZzlkQgVU6
Vxdlb5ybxkUfxNlNiVkkCIqIyLY133XEc2ZdRyWfUNjvSg000TuCjyDTTcqj
nL8a2UpS2zXwV1sQDn/1jawfrePWMOu6wK3cVSB8yeFgERT69CaZ/iQycy8X
7P3F0yH5PlQ+oJRof9ZyLPk0oKNOaIL6TiyIohkxS1pJWWzZFSLIAJZ9EJVY
N2S959pigt7MdI9dR6kKOH0DBI3L83F1UM6w9p2Dxqs2jNAW5ESotxt356Ec
VGKNiEHNxVbMm1GgPBJfDeFOS9Np3vn1u9T7Wn3z8eE4+9BBL7jHnXQv2eKq
z3bn0Dbo/P0fFfWWMZJzzxDLGqgkqTcjPMaWelrdgT1nUCWTixnCQ5L6FQRA
Fgax4+hZolQNIba80w970s4sAB5enrovG0nHSt2rQWrAHUw2xKTKezaz60fZ
OM0cV1xV1HwmHu71UR5rH3g95uXaIsfkc5G/F/ImgyTesbDNLlifTehpndxr
k64xelxzq2/Z3nBMK958/+tYehSQ+0kXEs66wpaggdy8BE5zbKSw6k4j2Jo0
V/G4qt07+9CaES6Cv5gIF7MdG9cnuGFUUfsnc1AbdcEajlrB953mvhI+NwEn
2juRao3j2xQQKCrEpPJEAtAfPrDAFHK8YJn/6+yZLGBXIEyJlQQcqucIPtVw
WVx7sdkkg3c7JqtES8JK4HtsF9Q+dVf7CjmRkyG1yVRXi8ab1Bmn2b4YwskV
Fc2ZNCyzTgpM2VvvXpDdR09DEZjivzM3vtnEbWgRC1IpnWvwVTRKtCP0nha9
S5EnExJ3Ux2XuV++kyYl2oH/FALqisB0d37QKwx06VDQjEQc2hdciCu197TE
gIOWc5HknLd/tSgVV/5//WO0/e0IdxMiKt5En/wqvWMRBNg6gFShQChFkRSC
57NrvrOAfXH6BocFxDxRK1+X2IUC6kJoilRvoNo1SchYx0oxxKXJCnsB9xE5
bC99lVbgD06MTOQAO5MvJrqV8SWrebEFYCq8nJwIV+1rXfYngXq4xFhHuswf
wcW7tcRpTeSR0YyzSMH4MIRbLUMN4Bh+5OjtsMjnrITMh6M8naBuDfvNsvuh
Fh7hdaaJv1zkAooW8Csl7eZiKM3q0eFen+emJPyK9+R8WDGQKNKh4KRRJ/xF
shqjbwGgQIDYlAL+Zu3jG5dIM+0zHPPY5J75S5T5WjAq5x+Ts+8Rf9hKepCt
Q2ypV9QNT3IT9Q94tNNQGZriyFtWD/RLtz+qq2qjvjWWnIx/dAPNpU8acYEB
XGWvFxjfAWmx1sdpK1edU8ezCZzP37TZtVYdFIqZAYgnia1q0cc35QM7qwSL
e0fIZPQaYmcTvMetg4Msgn9JLLoq0SeA/lae0Q4ijdADR4i1hKqbUrxSr/Xm
u4TpnJh6MyUfcOTLwRbkA6ky5rm/2bsKI1WpSwvz11WCCxqKWwUU26NjG+bb
EHFnrjLyTe3dXgeeI/McB6ba+c1xKzXzJ5dq3oLgGKPLUeCbIFn5P+XzIYqo
2fr7fHP4bUqzHN9NDsT0B9Th598uFvrXJ48/Jt7bK25qPaYyrqLjga1rZkyl
bt9qLlaxNCdCNe3vxqL+GVy4oN/KeL1lRNyDhksJ7HyU6Ime464hXJnf1bvw
ms+WCCz2GXRTv6QGoMhhzottEAtRtfFtT60OUPcCQ3Hs+BMHy5OWp0xD1lBo
KwvOeQGpJF/+N2bFmxTx7Hz606q37zLNLGgTNLzvT8hnEx//CIcddbAFU8hV
k1+S1R6FjOfY/sOn6DF3vQQZxrj2gpL4eO3g/dVLOoF7y7xz8rIjFyX1zc/c
Jx9J7CxyB9YkmCu5gYdhkY7edM/yYBp3j8WWvrsaXnwgA/T/lswYIqZcWwoZ
KxBstsz8vvo/G/0bw9gc4V5GKvEdICyiu+KnhLbkTx9YZhLEn07OcWJ9EkOu
EORcwLmggAbgEiq1clX6gcZDOSlYVpjP6ebuHhSE1KS9iHftZRZMWNzVKmgT
FTuFOYd7AJBrL/Eg43nJCftJm5TccCHQhopAmdICzmqH5JbrE0mp/QNc2o3y
pX7AtwGNsZq96qccEzbuQuJc6gr7nX25Vg9vVKLktyQz/qM17G2ChB6cR0n8
LeP7yqU/Bt/MMVj6VMl4Vli7aRy8/4z7Cs8yspkyrE1oKEG1GnCGH4CW3h1n
veImjkTV65l1GRdJpJy+7+Bgrniz77LpdMfZIwnt35oEfkb5/Cb3G+PFNvTy
+kLnGba+eQ2kVC5BVFRMTDBJnLQUDczj5BqS9TB9vEzZJ+gDy+BUBuo7/bQz
Fj2Et3/mOZIs02uTQ2rghGOiNhSWFsH7/Z+LxmwQvVWelHHZT9lZ8gDoKAXW
zF0ixSzmHcn+K7HBXMaXowlUamEh8AEITQ9hr0a9qlTeT35l/Bc6oJ9UMrPO
eY347xFZldWaNC3+RLGOaANgdimYAt1mbFOUjj8oQCnKiqzkhHzaOkr6FVpD
NOLuuwNRdyRDh8Mt3DXaFLxnzsib+15D/Wq7l5HAzsqjG83JRbJVQQMjoSFZ
tbG8QiWYmij/pyun9IJ/KIHlmD2oxgsOpL+7w3VVNmXIAdnyf0U3Fh2FMvvs
z52HiOap97RbGfT5s8Axzw1UGiwxPy3hkntTZRRkz5E6oHdEQXrx39EgUk2v
ZMuP1LT0SvywjZGaXNmGw6F9N7/nPPDXT5SWClnhrV7FUGErZoIUU+Cliz7k
p3xpH+PPvyZoI/AK5EXsqDac3nFTUkQzyzFWdXnp9CRB40QIcV6nZyd8ZnUd
pvovQaqNIBmmVCNY8tmxmzzoimQhw529DbjEA0SFak+3mMmi8ntqKATKzbwR
TuiHV4q8ln37I/OEpcs3PcnMVuo9F6C8w30rKQyhNA7ZsaMh3cZXkQ0YHtL8
t3OyUqXuxj4fPnfMc+7MDm5y7SzUqp9V1CPBFh2LZp3fDfytxvzm7HtcIpVr
pxSTFH7g1fnbp9svkJIC65e/gsNBesB1seD1Uvse556X4mxBWx4OAMxk0yNf
ZDu6GtJxs5gsD+tDgfCiil5l4HPoEydJgLjZGCUT3XIO48G9aSF/QR/AoQL9
G0RHH4SPUyS1JS83JnvRiJApushJOgeb8BMoxMh2tgW3cF/CJeYGl9bvB0qr
uHWb5YMIbDM4uVCuWsKs5Bz32epR1xBQtaz6jrRwA28oM6/Rvde44Q+BkcLK
nt9kwfQBNSv6H9Hq4F45GOqX6vGgw2wPyVncudBZMtA4r7MvuQo10joqSf2r
/34WL1XdQ6Syb0ZbDjdIQO0OEkP+o6XOL6onmmmkwvHsQdqXOqjwpPS53Xa1
5ptVmb1IP2zl2z0kN+2x2ilQudW7mXQmdt/FpwvyID4gxDwnPlj6aPbmKW1r
FhQaI2LbmCCnSX3IsY4HC/ouk9UaoHTBY9obghxoiOTcN8DcuKGGQ/sKGYi+
U0TgygbNFZuNB7wR+gy06GZzS1X9mn6riP3pw3me0U3iVA+jk7j10WHMhIIo
HXlL6qlXvZo+zScCM4RXimLDsykD5jR25t9QxO3+gmGHE8InfOmfLSLcCDUE
J60AIYX/xlEqb2PuzYF1nsww7lD7sTgHSffY0UhUYJLgTIStP0TAgQvlmaxe
aKVe1iT3OKYN0I+8focQk+deX/lxarKw2RrNwisTBoKSZHSPFhXz4F5oLZTN
DAX69vSf770uegZ9dSc29OGie4CJwqPUvWzXWnDs9+5YXBylt4ReT9NdRSen
EN5DQkucWiqkpQaMvyMlv+gGsc8gEOAAmOdsKLeyh5Z7Ojxl+wy2U/FBBy8v
Kl2jSgauItRuC4+XwjYY7Mz7RrKAdj1cY5DWLHNOWtggaotRyO0YXMVLfGW9
wGo6r8HbT/cUZycKhqQMwDQsVz58TJo8JdsnTvFRrpwQD0kiLUOxkbYK0U5c
cHM25v5tj0Q8JPnl2KXmT2g2g+YlhAw6CUIIRwYorK2V0e9tn6Jabbi9stEr
5nz0WY1htza4aww28v4qRl5rzwAFZNYRd59DjRZUkH6qp/YFn+2WlfldJJpD
Te5jtOUkgpHS+stYUhBFe+IFsBDrfAKQ2xJTSCwMY67j5nW1AO+MbNHOIEM0
faCnHxcNrEnd99NXrZa9AFqq0QZzYoUftC2rh5ZPd6sfRA6XjdMEs7Irz3x1
Wq/9jQU0lJhHB8xu9nEj8PJ8X6VmopcLt1xXeMtfHdNDm4SNWW76YSuoD2LJ
0rEKCUlhDpXHar0nbIYK+FCX2bQTfD4MNYiNqQhIoGk01TwYYnRlHsqXacqz
oGkvMb9jBfFayquBXPD+w+UQrqN8sY/iWXckjZX3m7xQF50tBEwQgKDL6tuM
3WLDdpP7V6BTKVsNz+QXSeq9wLsvfHU1xBnzXS3NTe1915zh7p2oIEjxOL/p
WK8gZd+hSGsH1z+fzd4A4ZQin1NRmBrAwrvJMjPCPs7XjQxxuiiP4GfgxCRT
I9v3Cs4d6hFoWzhhWdXa0eEIEYUIDZxqk1ck9SiZk73KiWMvJsR6wvHveVZH
ewPMYHENWb5vN+8GE2ff5eMVhx18p9IdJpv8SijV7cU1Ha5Ce+i6TZ2ws3a2
xia0Q5VTRgDGRDHYekdxky3nWBiHIodDZI70V31TOx4VD+OKQBfczebS/IVl
qRB7tKpNTjzxlaly87Msdi/cM7FH7mPxX18gZ9aGUvuP2kPDdEFXKF/7dDz3
hd5NaIQKpX7MXR0TqTJQ8hzhLCUt6+jUk84gz8U0AvEsgenKVFXBl71OXOn6
QDaXyPCiX1dbDl26rGMUz+OPDGfMS3mXEZbhpL5ubudOIfqh1GuOfHrxEZ6z
1behYLjTzLLtc0jPBmvxzUt1WAXhvc6mP86khMNqjpOs1CkTdToX7/PwYt9g
NexEnh9wM4ARGMstGLFcU6RURudUO9dAuUAZ7N4ecQGPCkGcU4GY8GTnY9Cr
/XufKFOwIPsVzTUGbrwDQTaAugDHfbIqxzF+/qw1w0kwJfmJ2xeQO6hVmYM5
+kHoeaYJ0DMITc6/FyHDPb7ztLRLOQYOgFCcdee+jplsVBeIlpRiOjZTZqtH
MWc/y95qrc/j9Mv+g0h6HW+WSSQZbE+MPQCyS5i2wvXcRlFnRGvOxOzUOAHA
XLMNlBzkux9CNGxk15bZAZ+5ZVXDzi65wmE8bSVX4gRI28AIbDhvvMeq8UE7
KHSvG1kSgmKlNG/oBgG3GfKU4sq1pUi+fBCOHIhTna69GcFAfPW8x9dhy0S8
FloZbiaEpSjvpx05C+02jvhsfs3h5MqSgzDn1bK1iqaLYxZsW9tihG27hWI7
sbMKUDZkremFeJ91QB65zB24cH8jhttTScJf/c4+unYDoNNY1BhXG7ZRB4eM
YLkefVBoMOfl6P8W4sLlFsfIVobuJi1TFWn6VCK02O76dBKgpB+GGxOJ6muO
4h9APBTgV4RaxRa/OGrQWRIhUL4WL0yjcuEtWILvjJiNyhfHPotncpR0mfKk
5ZlrhH3oRtMrgxP/r35Gd+9802ngVj38+8dJZBf0zZmWOo3VvZreayMPaQEB
M9S3WCcYMHF5TjclbttJOZv1E6AgUx/6s2h6aqgycuuigmK57v18Iyx/Apbk
vyw9ZSyRvZyTyFFVRrjlPMbZzliVkNRFfq3i8NosYMAXv27gVtQTW/9divv/
GGIUlxsAaNfBa6X/CHRpWc+ZgB9+gxoqsCDXaYwa/kOGTxIeI4VHW7MQ+aS1
55Z9DdG0410fDZDFYFnin2jF5jziwEE4iHMBwoKAxQnTC6VthuCWdB0+0sPO
Dc056+zAPmap19iQigPNPEag7+Sdn923TM4tLJyC5TJ77RRZe68hiGX5imtE
KTsu2hp7eocPbHjQ+YtR5Tven8GA9Na0WCihZ5q+NWza3VRsWTcWjyA2nN1D
U76BsDcVZMs82NBiQ5NesjfvIzZFAugDh5phzgRO0hq7V2QCBGK/57lWteJZ
j/mWZaAdMJa8L68aoi4pnKXIrxJHJGBCkpCuMCNmaCIlTw+z/YnaELHWR5Ov
Q8EBfdCNBYmh7RFEcq2i4+ix7W6MHq09919VFhsIDlU34IommymFzL5m6RNG
2uKZXL3iMxRaz2VQXEWy2bw0yTru0Y1ctQ+sEmh+0JK/WCrBtu7APUkXQ4wQ
YdjR6/hCZ0dYiAz/h1Ad63Q28Z9irCo2As8By4FOzfEMhGmneBcahpcF+EPX
gONrKG26uPI4bFMR7d5BObZp7Uu63AzI/XvR/t4rE0j3ngf0Nx0I0gBmY7CG
3k/KLsqS9+ekAgXYdXFQ8KqAvcd0+czNp7WGs8vmIOLFz3J88EkcSS4bBWl6
fQT/hqzabCzLE4DOxx41JFZt68GZuB3K+vVLuDwFlUHWsn0Y8MBH3HL/px/z
nqE2pFvtQLW4XWWiI1ple2F5ORXn4N90l1Iy2krjKffCioEsapfgplVqoTTC
M2PjmHXk4woXwGnakRfPgK4skDw4Tjeg0MLgm23VyJEiLNSW4DeWpwFxGXla
IBUO119zMGiLdOyDLG8+EXEgTJmRMSeNkFpxz38ha6HpJr3ZlybTHkvTyJwN
zFeNiPuuyyzxn5B2Vw/omobt77xQeI67U15IzEwUB7xgVWP4V0aORSNYkVPX
Ih66AhxcBzYU8D+pR+mnnTsMQdQFDp/knNOhtymCM6D3dJi7eKFDxecrOG15
AiXksLDopjZJyQFCNLUPbc5JTr44XeeqNXdNZhpsNmH9WNr/U7ccKf9c4g3H
dTj+UV4SeiXLBenyMrKHlkaFMncjWzcRnjFWIqnsSayprZE1fRIqIBUo/SHq
913xOOyC3Rj4zX+e2Hqkydf1hZpiSMsaDD+sqSQZjYdkvGTGyP6+1fXECzKw
e1svrsV5F+nk3X+9x3f6F5JRjOEZxXL9WCQY3yRUuRTaNTt3Wh11UBsuoy0S
WLHSeOSaRBJSEbDHddJIsTl21vVTBtmyrDt5C6nkw59AeMC8CIdREqP+hq01
H39MYIAA0iOLwTmEjXxOdh5qagbyD/lrqVTDplGUGvSVowxAHBQHzllKtKXs
5sojFgebEgTNOtLcCMdXRVMMS/A4nZ86fmLBJkTMHWLEPgOnem4kD9XTdbib
4oqHZJO+wn/M9Y0Vj8mlyRpJgS7DRnPBR0zmI73NPr5SgYH27/bmnUwsaCqC
nnHy16ci5x413kI/1Rcn6lPSFM8fBCIpv3ytRzbfkv+qbYYDkHQGmq8CsjbZ
Gw+J31MatC6Im5Hp0x4O7Mh6IJg+9rzuis/nRbx3naefgg/aJh6m0HCV/cb5
hpU7rcJD9jN3KM0QhoGobO0RRF0Zx/ekyi4I0xDmrYpo2mcudvZar8IzQ7b7
sAeMO/rOK69DOHiGvNuNcIoSU5YUz6tX/HwOTqX8xgbmTpbDwoqpoMYHBPkU
kFmCeXRiFRBB+n/Eb3Qnq+2W7Xrj75eGRvrkMp6zLQMP1ez0fyJHaUIhUjDU
uMldnQs/U2Q2Rp+b/Jd244mPTJEhPOPoS3pfXbtyhnz4TvPqqb5A9wHX4iTx
gvfItdPoigafOTvC7jJaaPwC9aBOb8TWLw6kL3BVQKUUQjAhLE7Clxbbd0gJ
XuJ49BelfBVMhvpNNiAPIJnUcysjI3OUHAEPfW5g0sjmtPERWMf6J+q/HLK/
bTzBeptXnXf22bxoS7UaA9Ry0CBRsGHqS12TjWHRWJ5DeBiXceTI0hx5gV1e
dPvumayV5sMbAQy9ZJW2FN1wYw/6KUTvDtC5EoXQvnrZP4dVBpSwo4fu/Gki
q7juYM7cwjvCIeX4Br1pq56r4xC4AxnyoVEs3YJsBJpx2dEqFJMwyPDxXCqC
ZqlRP/DX2VqtTKuEoAI1SusVqd4B3rUzMJqD3cbOvot0NQp1bwykcUbVyIIB
DW+7H7E1i4jRWdecWqh536EavKo7SHfr+YtTAMZBhu6LfKThIU6YxaCStw5B
it05zhh8EC/QLeN+s2zdcJV4ovo/1xqDsuCk7prgyGlZQXaWWZk8IfQuJNiA
9YBsU6Uc8i2F5uQRcRVLuCNP0zBSr/SDBe7PF0HnoZKIbCrd10ek/56dkxqM
h4kR18qdvnrdLoYHk+hDqfARDXBC9h22NkSDe1tjdYYlB0qTJPK0Z8C4dA/w
dTkZ4mrUIE28cawXg67Gvdg3wdBkEwBXRTRrwx4KB/R0Mu4Esjx4gIze+SW4
Col7nG+cB56PdLYAs7yvFcZNu5U6tyJHYLeHrxniaE60VI6cHLLeAWmhqWYO
PrY1yB2It5FC/5lj6fNG/UF9kG0FC2GOYFcgU5bd75ZJgA7NAMEqi7+yQc1K
Akx50RQagdOdrfFs+FvKGhPt11tjjl+LStneeq04+dIlvFcePDxPTp6b5lL2
XOyMvdHL+MsrQ34o27HCf/M66X6nByL/u2ePG17k3qz+tY7P/5AHaInQtw+U
WxIhSbww9dIZBtk3inZzlpImHGxZWbzgNwK9XCzCuUU1OLaiSyRXd8P3N9oE
e32YkktgJKF9AZC0iOT8gaAgBnT3TVBVK9v/dcNDB8ijQ3lO4Ht0bLphlU6Q
5l5GH3gibS7i/9cvQrcZn30V67jy9BhdznUCr2TPRViE56QZDyckFMl8vkga
P/VjiJI/ovvDM2ZVb2eNXEyhY563Gbfl9gZeXC4wzpqKf8r+ZdO5Y0oM6SC4
v+M1pKuPEWFKxYpv+XbCMrXqKv+wnk2cVWNg1t11AfJEpDrC7XmeYNA+ABrw
YSgTwdkjqn7Rtx+Y3H8ITMmUg7xzg7thqnLQHPUVxtgoIKHYLXsRwrBfE4F6
zyxEQ+0vvH5BIXirMzParQMMWWbNdxlkcgEXs+owfLixjba4zyzPLsBLHvXY
VlB6dZ28R9mMfR6qZ7EF4lEs66bFZ3V7mUoIz2ddhl2BvbtRg5i5hE4QQ66M
ZPK46DDaJKOYkoU3+YLKq3+wcnJm+vKlGBGzSR78bl7dfe8s0LTAFBmIF7h0
Y149c/XtmKiAQDbexiOstzFunL+3lnl8YxxFo5NlZ/4rderLUBCJvrsBFTUG
AaXS12TqHN4zDsN/KWYp0lA+/twZAH0003T7lGSZZRXmxgETzAFm/F+nZbNs
xFS3yft7W8GvvbdMIHfpNNtfLO8I2hfaRCCcihU2S/j00jLNtmO3f4KwpSKb
1gxCmJcj6keEACP2DxURA+j+HkU+qWTey4KyrxAAV1/JoevYYPyQIGocNMie
r3JYvv5mvkq54Fs90PkRI32tPkreFrDdK/Av3R5KovBpbVBHIFPfefdkIcyh
i9Y2/ZhBrKst1NZsPT1+QK1JVzTR1ZRb78P3GsKdhJFHaTRtxsavOMWHceMh
UsgD0xcEz1JD4gO/iEnPsVPdTJeWlSRcy83kmDl/XCn1c/TVxr3n7uZHrQue
fqdtmAt/XaaMwhuKkzEmnQY9oFlFJXTZVgPWB+36kaguT6T+sCVsjxniYpmq
MTdiKuwLFHjYbFyhUmjEFoQWT2dlYwT/NpBIRikksZaLysMJCPp4fSH8wvwC
LB5xO4acBuq75pMPYmzMiKjVHt8MC4jR00c2LISi08ILoreoXiitIksLAJAv
IA/90Tj66rv+7wbKoRstMeqY3ihOav9EXRl3iNO1QaoT8w33WARDAloKNR7I
jUXF/WwQi6EmmvABf+3RQ0pquCY5c/LQ6QN9KxMp3oj7NFwMsTv6daDg5/4s
d14IlM1K5EIBs6Tp352kii7ENsZDXzVEXE4Jr7sBu+zTsVcDN3Ceez7rlj1t
sJbebAqMOKixvc2f4EkQuWFmxZrkpi2xJsPJv0Mt/HHQhLcUYtK4bQiIu5dr
/lrg8CQDUlGz7yp5sviFIwrFw5hcwu0G5sCVCzkRnjauv9kIPW1vALca5Nr3
UcluBbpV8kkQgEjVTlS3rcQHjmAd9G4zmjQ4LemK2VixBo/mTDOQx3mBVy4B
A3gIHB1dNCg7Bvn5drdDTGDTQentAHPtNBR6JIc36SKMvNwDQ2sQX30QTY9y
Gx4DMRSax8loVdEkuLoy7TH0DdOloBBf+Io1R3iVaXPcYgUch6YEDd0rGdpi
AJjEoyxW1cXnClg4whT475V2DjEaAfTQMQvRCkEIu2+wE8G+iHLaVtK6Oykm
Sk9jNfrGWWuCN8zbuxsBjmLgLJ02eYkLcPqQaMkDe7Vt7BQ4lMYRdYYW7dMV
WYXuva2pvTDJyirWgtqr2CXZ

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Z1kxvUZ6A6pwKaxOdYs07NFMnLFQMgt2NVR5MKR5RKdJ8c9hslnSwQz63pqgbJulNL2IsMQbF1Uj0IhqVuqvHik8GKPJT0wra1hxuKAB80yrxPtVbyBlDdvuZxuBjXIgzc5B2XcslaeodZFtBeyMeUYfEN78Sx7u3lzsX2A4IXzLnEWV5U6gYlyO2tGw+1I67OKRfL/w6Pxg+cNr2D1Y/t3pkMof+6e8VFnEeyhkMURZZjmH8BLAFnfxiCuq/olqhk7DZL1R82RmEoXx+wbLSvpbfG2QL8eIpJRKtdLhMI+awtAMQlICoKv2h8eFH2hOLeZs4Ba40804bz4yLtmrVTp3GFid3pwjDV207PMVaZNJkNeuY/pJYW9E0eMbPA7pW31BCf5LihD7X88rnxqQHlVSdWYh3NUddyje5HVk0nH5pLayjRckeP+mvB4P/g+FitM4pKsXtCIE1/KiJVTqtwM5Iw9O4MRBl8mBzz8bKqS2a0/K1lQHDRQnRuvCAAGnJWEQsCPpIoN5c0oZpAwiZdbL52YSYTiVVqhihWczW6UhZuRZeMOxz9R+MJ9WgqN9G8ZBrCkw6D+QDPX4/9cn3u+y5UW2nIDEJffCBMpR/kuRRoJslwrZk5ZDEEmCfDKurHnPLZWN7/EKNRIgFauCRunvPPrtTlKZ9NwMxq3R2CR05sfVdUgaTW10ADc8U9iIllLO1mukI+s2BAfAObkTJYk4B2aiClczQ5i5AcdQODAnRQ8l9muDT0AQ8JIv0EWxdVNGNIh/VHC4Z+nblFo/rG0MV1XPawGUvgBVjKf9UFnc96hdPG9CIkAiQZwinkcujZqs4NNdG0Z1NyC3XOuWYO+gwaNIgE3WYo55d2HczMMpKAst0xwvFAMqJJtF1hL4sFtb85FdqA/RbrQkMUco1ar3tc/hdTt4SzMgtHo4GSo8zORO0yhr/SkgUH5VvSAJnz7g/fSlw2EhZbl45SxnHfxCCsBxBg1sWKrB6UTp2ZTZb3EfIuSXPav0q6TELFVn"
`endif