// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ya4+7Me9VUIgCCIO9UkhOxnzPAP2o5LlgDQ5aTqI4HMbKRy5+0cVLoaOSi9u
GAlzPgLuiYBmm2v4YGFnaJ5x7xvZPb41JwHg1hIvSr/lZMW+zy7GSNodtEyI
tUm7tP0SFihFDsaVnl+ROvk0Ji4vJpT+0/OtFRplCi5IZ41ugaxhBMaOJeQS
BoPEdRtUwUuDPQWQyKpF+3x15dAWPUulgAalHb4VhVxLEnfvuHhqU9NsQ2or
OBvF2/m4EJoiCUGit0LlvCekcF+01Qz5RMV82X7dqV0VzXYksGsPR5sOlxau
R+fWgcSvZXOBVrEkP125FRQSYL5VhSRLCglmK8VgVw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N7qo53YoiR7WEWxzrv341guwBJuW351SheZ6IOUukZCTW1Dw/FJrm/sAgOqU
o4IHlK5cp/d9SRVRn3gJBX+fjXpOF98hMnNybpWYOp80aHQUAfK2N3gBLZWQ
Jp1JZVUriQP5f0sNPU7PeS8crUiZjxIALMguCCoTNhK4NPW2lGgohFSlLx2q
Nsgnkx0E1iL/rbaEO1jxDk25Wh52wCB70J/XcD/kZ02HW+RTRBgMk8YgZthj
Q+qXHWGPW3fFrMZ59jj5jmKGtxkGoFFOb6cFVwc/t+YUN9o13YxKTV7+05PK
XmP2sGY4fSmojFDq31pwzZNu7Gipvn6sr3S18Ctuqg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nF+fEkCdMGt16BaVZAmMOlHlcszlyJvIMV6zZ6X2lIq4vx/2ZYn6P46oBxQ3
PEAOVPOXnW5tUFCnoQDhZ6nV8g2zwkRGg0ZHcSDeLdqlN0Kg2+83XyXKxsu3
s0vQj0Te3G11Yex+Vrc3JUflqnVZLG/MEuWwPflsQStyMazB2uHZ11br9t4q
fOzodl0VZ+5dIRyBsYcCWgHfowRSc2/nRVbWGgoKFhkt1+S+1LGDn3VrZ6v0
4Bq/SEhFrE1c96Kth09Tvdw6hQYRjug3QLJHvcpKowis98GFsCTCCRHFVakg
YGiaxh8jC/0U7ktZsJSaMf6dfhL4pPR/59cb6WYb/Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UzZi2WOowSw2rVcPq43G3JIsb8AQkXvtIy6VCIIfJY0ETMWtE2l7ihHgeC1H
mKe2FM+7x4afBMXNKkcSSq9WHZ7niWLq+T9BVi2oDCIhxEUeMbDXUKvbGlYT
w5nO1G6sNyyQ3f66gm1Hm0EGt+K601p291hJ4+ItdNC9RRRZk3DQZ3brUjub
4sEk1eYwiQgms9Ax568Lb2ctrV4xrt0dibVEbCfl2r6Ch8bMEQJ9y9aS+kut
HlVrrif5h1pbVfUJbopNOJ5RaXsG2q6V84NPnR4p0js+KrldIq7GQmniHRpm
z1/TPyA6Pfy3dT6NYWd3p5zFnnQKTNmD9J2ky7CKVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U1RIohIREkNrhR2jNVmLSuAsTezYfKfJe7nD2LCSgqbf2Pn6Gji+pOw6qjXV
Dn+3x5ViK4oTwlMzoKaAhJiGG2+iE/hk0+8JtCjBRcUWw5BuJhcUz27ZnZmc
822hCksovBgawL011hAelbLE1uQ0pJr/HRBCXsjP4jR+kO5Blt8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AE4dIxDS911N5G0c7bO19FbfhMlxpzatjReFnfeHCANnXNGuPhSzvUAVIO7x
KsqZ61s6VHDKVgSZg56SlJIVaKywSLBrQdtfKefVUulMxJPvm3sxF2SCkgDs
k3tT0ZkDKqNJq+ct6LjD/nO65sw3V0ARI8GOzntie6q1+rhLzUutaH3IiycD
MzeNmpDm4/SKFxPVoe7x3tNw8M/B3Hx7XrPX4rD2fy9TcKWKh80VEVzvduSv
B8vmRMwh2YOk+PsfdRztjyL49uCp3+W4qAG2PpH2ZbyWrI+oNu0OFMN9hJeZ
9rCQqkQHnqFJRepJYCX1wI8XpxiKDFfeOb4r72WUKj04cCQLKlUzcNIp+do7
DDQQdvY0CMmAPq+R9gC7689IcTi07qenWZrOvi/HdmhEMAML9toyVdpI4TsP
RowIQLxdxioqYspOsZ8Mg0clQeep4z4PntHY6T7fyZoI3THJT16Xz6dLpak7
JEv022762pNnBq690sYiY61qF/MMCGlI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FoKMUeZbscgYKXwEMASCa9UGzPmoILlDSPkeKERbI6DHn9LoeLaBYa1OG1Uc
v7SBsjsrGaFKcEpXynvnXYBUi3wvTqSV7+ebif2/Sn+MVSzn0G9qWB2KFN++
ZGW5Hi2ws9If67WzDBWKFLwkoBjZjOcqmVCaFqfwmyao2XJj2yA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
abMvlKOJh2OhtCml/q4rShGTC5Sf5YS0ittC3qw+RtuRVTbicWWbp85Urzlm
Dv5VkCO4TCIxKoVjEr1ZytzZfKw/aG4yd/W8FWSWCViFJ9Kn5RBlnRYA3qpG
Sd43vjNGpYMiSfUF8BYZoMhEq1f50XfD+DkC1BRnTNfInNgJfng=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10848)
`pragma protect data_block
5UNPmhgRGbTvxIR1KqGx19TGFQiJlJJ4sWqcTluK3VB+uRmQJsFFl704CYFy
txKzjwRTxMg1hQbDfIzFg1zzy34b3viy+DjY4Fkl7+DznU9yYJXYE2Y6NBBi
GaX6s0IsI9Eah2zziaoXgmh7g3nLEwOk5+bWZuhWBn9z3FS1jKSnr4JLOC2J
WPsmg1PSIcBOPgfR0HiG/CnQyogNNZP0rvsaTx9Jl2My8Of4Co0SCKuSZzJE
d1DJxBxQD6Dei8xbGV8KFzMOkzx5zQxdA3OxV+rNaxC+/xxvO+WiRdEiVYCw
i3XbYpGPj20Uj5VTFdrPHv8lf1ryBzgnIgpfgF3LERv6JVXMU7UX0On4Cg+4
0CU6nSAuszfCBziflIsPS9aWEEyzemujqjuIlxacf5xHrYRYvpRdVw8KsbWT
z3+/70ZhV0u+sGak0FbsdgZytJ4qn0llV1Z98pPCDjtXVL0fPl/nNQt2UfsU
lNM+m1RcQc381sB0y1GJhoJ3Di4bI+4L+vKyBYlNivgg9rpiHtxwzf+4qECW
lIAKoRrgv8+B2Yb018fpb2hzW9ULIndJsEzwmwo5/UJ/GwQzkkK5ZusiuVwf
czsfGCd1Am8kLD9RgtSTybH03R7P8kzXdvjyTy2a0CxtI51Xx9UZZ8SW09zt
Z2tgXx/EuKX/G78ImRcK78XKtrQ2YKge7f2kk+A8yB6ahpg37ScSFsKp3HFj
djXLKWfsQNzec7IGKAY7KQvQlFGZLxzIT5sdaK0K14EFRIow0qEv0wRWice2
nK2lbnbC3UaoEu7f+CiufjIshllLrHEjodWd9VOrgNrBn0hBLpcLfP/CREiY
qsTCM/1+mFhZqhb1cqEIjQ4XV4BS7KfqTmfdP5j2Rwtlvg34k+1BFvQ6hhlL
KxRq03/u0ig4VE0qxTbcGUNGoFv+1RuO3SfZigdtGwxmtg5IWPS0eyYzQ76p
5Mvq9IDf7E+Hs1tNddo3vT+ehKttXBjJwbVqu1sW99LwVloixctBcNV4dCzu
ix5BQSQy9uBzvn+ye/eS4pcLcW9aNIEiecuc3YUeYigKCotpH3PDnagDHDd+
CMjAcduretRMXs10kSr1OU1vFBOX2MZ+iue3B3LlD4t0Y/TiZTpYJNsmLSSq
kIgMdsOOr9p5yGG3iqdhMmx4zKTnIwuLo70FVp/gT33ct1u3Ikl19UTApgMp
eiZqbMaI0JEXsdWKwfvvZ8gO+j5tzjGHfEN8AtSwmLjY+f2C4FpXw6MxKBGm
r5hvAt9Q98WkyKvfGfPA0Ndlk9X++Re3t0XXH/kNTSSbB3XvgwGdsPrk1fhR
u42J2yL6nheGIq6x4L7Oc5JT/0e/5cF3Ofghc6lzTuPLBjvDUhGxI1M/XICo
5OKUVoUk1cH7sqn6T/YHv/wKjYZbmKD+83G6BSRvVcHWZAhgvcVOTi+FgFSC
y412Uen4EWHbOR1LiRAuEkxdhJ+bD0qjpjn/24D8CHhgrlk3GfICzDFMlrDS
aFto9W2yvljjupxwH0hWAtAQPWsG6M4jXcfEa5nx3nm1zVEIMEJYUXh9weQY
3AYmfBNBjNBEhv/AMCj07foKUD3fZNKt7o2qpWAILnIGhlVICxVnmQIq45C0
lmQqmExdWOLW9BPkMJ9NbDqp3Q+KwWWkQKhudeDcXT/8idIKnNy8A/zMUMBe
ABIgtkQJMMeK+hOmO5lYvmjWCxh+ZAliJmU0pGHB5vz1ZFa3l1g50pP+oYpC
Uz9YOMRFC9hX3jelygyg3RFshUTB57FgBNLuCjSp0V+PhksoY5O8z4isN9YR
YdjBPI1UsyDD/kQm1/74GGwWiD8hvFo0U+KF8oC1Q/5H0NrAS0pw3GUAXVha
iH/DvpjsF1a74dlzkGjmx7Jlv039BL6bTwZ3Dh6GMlD+5328cvo3ePuo1xDv
GEA96waXZAZuggM0ma53EzRdlTmpoBmEr1PXn5NNEUWgj9oPHuXO0OBO3BDc
QXFJHpvczjIqtJ5LFiTmA+OnmXvXMaCnowR41EON0Slq4utbeYFBIUX6vNoV
3RFfcZDyh6Eosr2EKA5ik+kncjZ7v6GgS4dWjwMDgrBTAJrYb5qnxrkCP3Xl
PsoreHRdoYztJEVxxlyHLmuIdjS/vKGpQ0wU7TZZx3Asz7JdAvrHE7os/rnc
QBupBghvaqo8zmuk6cXv05+vEpkGC3oV4RAze+og/KKgUH4y40G2YxAneZa2
Gu2pz78uC8j8Jv7ZZ7KNEAC17Kvd87ekBiCbuR8SSyVl9pryYbZ8IfWtg+yQ
PoxC1lAibsZQMCosN1ySAI0XV2162Z56gAiQiLFfobDP98pPM+sQQjDQKifM
QH8ZWKWkVTYHqEh9X3Ob6pRH1Cr1kddgPH2+0LJRCUldpqXh8Ju1gZ6DeJ7A
ENq4qLPHrw0kcNnj14nAEqIATANum9g5TkbeUDkQeGREJb76VIhsugEJqq96
nVOz7ZKfCZQk2YkzcteLeiU8kEN1K5a+PElzhPJ1xlqkjvJvTIw6sXN7d1qI
xq6yBNnOEGIlhjYcDtcDeApbTIC2gEkQwdvWx2tt0ATxZZQlc0c3pQjsFbry
1FowMs37OyrFzt5AUSEe1FUv+ejLKmFvO7L2Y7/uuV6LcjzYYNds7klJKioT
f9dH1czZLK8J/2euRa0PKtwwHnoQuE+Dxn74epnVrOA1m/8Hg/GkzU1mMMyI
Qm+PChj6iywAjS+gjvJNeKIyrDRbmq6ySL1PzKgKASaaJd+cUtshqqVuN0VE
741IC7TlpNeU3OqQZi7bDXvWNNTdJuAeZA/O9GQgR2dhEnDwtQeMwXVpD6JP
W4hbeP4Xn/Tj0g2gVotdWb8/zEv7XtHzfrM4mVKNxZxZW5KZCZZu2B8pePi2
eAUgJMfDWiownF3JwuSi6up1XyIM+9qTd/5UNTvZpIhRndd6xQX/s21eUWUN
J3CKIGDqBY/uWZ40GtReWRP4iwtky4OuvmbhVNhOT9wMtuaygMTFk0MV9oum
rLcoeNyM9giBfD/neecph0/J5loq96DijxwOrp8MyNdfFMNb3s0q7MFBtnrA
liwxOCg/ciRuUVywMtuAk7AU2WMrTwgB8J4FjAY4eKfCBe/Z0BO9whvx9ycj
fnD1N9do0asMMb1gaSv6Qs8/AoAjQCjefQXDcd1K0dqiOi1t5RopPqWCjzmV
xVWAMX8CoRSjwmEv1TiJy3YC/MaxP5kxHlJh3vGGOLCUNqjTcyWyJVWrTmTs
4f30a8qSpJBPp/XDqjpyA6Trza5//v60ITOzy7Jd6nD8/x5GeDnjg1iE/xOM
73lTQOd89Iv6KWXQd6PErWO4sTzGyimwp7wvvM/di7WYPRQzH+2kKPaoGMCA
4lNvTzLhtK+yxuN4UwZPU/zmh2yJfNImR7NyB8DVhN49HU+O0dNnrcM6k3Mo
qrkoq+NiD0lH3qpZkq9gdLPNcRKSBF5dq4tu10BCkSDFL5OdHG7WtSgKn03L
tMyzkbGooPXH16WJcRaMyE989KERg0tJSAFqtbg1XOW3cDLfnUur0hJ7+hSi
QAEADPfDkv7AjTsxmYkL7378K1nKF4Wrih8itgDUsFU9Y+I9r6ub2DOas+GP
pOak5JIVJXKPAVzo4b6jLbr5eLjm3w6vj8hHZ6/s4YMxjxIodjcivWiO9fpj
NUcFZf4Q63tpHHUEhNeZXO6zArXstSXtSR6rIdm8+/3y55ViHaUX8u6zZQFK
OW1bRFtYDUmNJkqwTEVzEn2jW54k6EJcrAfhZOyX1FF6XiQNdKqw8cqVGpD0
3agHP0Ux7DTyUEkAbT1VEcmwpYfuGujybng0kbZ8cCfIXURm0cAsm+VU3kv+
SbUDI2Lu4GLSPw+AnIiYMdpC+lPj9VZ5+vopDKWOh+3IvPKVhteTNFoFiejp
cPXyNc4mJH1+PQYsyBsjj1yyT3WACVsuRYkt4NuG/gYGkFI1sbGDMEUKvnIA
7kU7Fgi5U5WRxTDpnR75X8jwSuNFZ+RL/vap/XBQzC/fZDf3Ce1JpObla4sZ
fT7wWXlYOjumwvbew0fvX6aIiOLjLz4dAOFNmmGci3Ef2CEwSIOsNSJ2ohuF
WWCVXT7Up52gGG1g0bettkvDP5Z3RxWbe+eR0PZJosJDEEnN9AZrWUSD0KS2
37p4QRlSSe8WeNNvrg0zi2hG+QRrEJcMB3vhdpfS3rkUcKDOddhyxBFfuc+I
VqhUFKakr7w8KTssPsI77ZV5eJ5qHhwcXtHEikNqAEkQ+0O4oZQeBbARtM/h
p4fa9MrumyLE3KKIsXVA2Cq1wwd318eoX52cXctktxedRY2HWPxeD0NISlNl
X1aEFs/bpAHpKnrm5pzLtykdeJFyRE1tHmtGvW2kqMS7YRO6ZnLXbyz4ahqY
uI11rem899gXEfEnh6PMPocbZVYAJX8IX9KvLEHN0Lr15XA75oNDGleGODDx
rrQsmJ7MStYBskISNGlpIRtIN/Mr32ZcflwzexK/+l8RJ9QA0N06du5rLgRm
zh1+42lXj6bA9qOuUbvhJgZN4WGyjq2J5ntTUe26PsD9z5hGMN15H2GSvVLQ
82CSbW5LJ9B3RbSP7CW+y0D4+v1dfk8fhgAgSQcLF5PHIxAJxr5Ub8EvrHYG
/y3o830cvZypdBA2yvDiF9OtzSKuqm4LxfIm/5AuX9x21+75UUenHQarQdpU
ZQjtmotzjw+lIP8VlJK1zWZJhyk6LQ8v1W+wt4A/qRa7ULv1SfaSnBcRQBqb
AKFLYmuo955cJqmU/0dJfRd/Hp9EhUlsnjP57HMNkgjUjtaBhGQiN2zsZv72
X30mdZC+wv5Zwf5DQClA4jcIhBvCyXU1/Igo3AjbFUvXj0OqyHfIaWNfOYPV
46t9WUNJ71Zvsdk01OCYLToj/GleHhQvd6VU9jJYWfCp/uPOvQR9hjOlomSK
zwI1xisNggiD/aH77U4Use4XWfu2YNhVeKAxUUmf8OFOUPhqDdFvGUrsIXrM
+n19eQDNxGXLeufHaiWc1LSn8KuXfsOvchxH6IUwdPSNhOB4hTIuty3IOORw
OXAb3BA5Tl41zncznNrP+hnRvdJKYQEX71QZ3DAs02Ogf+dO2CnjmNOWwLyA
sovwdK7YS4n86+gMsnV1qFOZeCLvnaZHLxMSx6KmSGq5mj5/4jzYtUbez4Ai
YEJ9HHsaraeNRDqnCODfJ1ff9ZOQn4bDnWlgVQVk4oxw/h633s4qJeRUm+tp
HycRW7PNdZq2xw+wHDCQLqFTQPHTUWzvVdAxLsNzqEC8NPgx0wGRi3R6Jmoz
8/xSpwkVGLt5JJIaJvww9SVL2E6gaI2kZdKWs+ILtw7us1Lh9dBhEpqzF0gh
aRaifx7KHlqi1+MtVFarhpKkBO/bw8pV8YLfwd41eEf374n2Sw6vxtvnxv9z
rkv+jMFaE9hYAhBdQEEppHItqWZ8ePbRIR82/od+OoldNkbT9DJ53pCKApxR
ATrduc95wwvIQPxPwcuHxXldWzIZ/mFFRnyTxqfgxRJdXuzEcbVknrzDz3Qq
ZrHOX34sg1UYLsl0V00syJY1Fil7Vk25AapxoZTM14ejLHrmmd2GhxDs5tFe
+rx3weRyhpmSxIUYLTJol3/I/LBLJoQT7mb4Hb/oydX/uX02oYL1brkrtGJT
LzNZGqRue7ZTifDUfUncSCHfdpxDTw3PbxhnEvnmm9W+pMOQdQY196P+pwZF
OPW0eLaJyjUQn+IEIMusPmHG5Uw6qQ88g1QQiT11o1ld/mAitruZWrOGk5U4
v/zw5N0Zwf5AgNm0+Ph1Q37sMMaQYr9K7q1C1KOdZMxGX+fYXP5mtT0iLMfi
BVVQaNZ2usgqEp0Uw9c7xM2LwW03rM7YO0WiVVsfK7du0sdwMBo1W3+JTx4r
raBDBZhT9Ecfre5HjMxurr0N835HrakoYy+R00LLlDTE9pg/ejNnRHPy0C57
oCuLohrNteqHTPGrQWOAjeAN02qTDrukxUDLz+QVKYzc0Fjlws5R1qlPueTR
sXlMSJpsH+z5IPt1EHbcqaTPVjmjxj7T7/LEGbNb4Gmm4l2I5dydv1QS8Rmc
dG1qySP/iUlplHNnGBD1wuBmxe1mxL4ACEAICK5v8FqMCudWFJlAVojdXKfu
7hhyzCULY8mSwRGvyiWi/1BKkQyeUgrq+6k2RRODKSIHZzEyp0CRYT1glvOh
3rFQW8asv/2JTTtTy3Y7qlROqbD+87Dn36NO9ULZb9rUHXpRbY3Jz83dvjlG
WQENL6MP8C59+14aenpBLRCK95yqk9N0NlgCoZ3CFuCgfxLhe/bswLOscXMr
HZl8jI311om1ZkFH0OTGUyvXNAd79ioWuLAyJjZdVk/+ioYMnCpzJbZG19ot
H1XGCNdffcjekeKh7Ji0fjsN2UQscRXXagwh0VP751KtNw9gcBFVmYfB0fnR
J0ugBH19iKcAg2evZTwXC20FIqj51UoDk5Akc9pmqyfDHoYnh4e24tNR4zW9
eMTNWGW4ozqCzN650/xdTsh4yCGN6wxJhUJ3dIWRTTiX9MIqw90vwmla5Kwq
ay1w397Lzqr0iBIyHhVk5HsX+vpOI8qT3xv1uJxjotSHYt2CwjznSzC60k6t
CA0o5/tVLaWMhmvEOw1+z/QUId73qGLquHWPsQ2pM4h+MuLA3PSF80cdeEau
qwEbFqqO+pKzEOtZsL7khpO654KWBLlgD1ry+dIkjcdxAzkz3LyS1dWHxZLQ
HC8N8CwTB97egVc+1KzBtxtr4ySBT2uTzVGDoMKLaVCiiYYWaW9D/vqhaRT/
nE3cLG+IBgl5aNo4qkdmZZ15IReD5u8kQk8BxZZtUJMZVp3ko5q6vQvhYfRB
yl4IUA2FvW/yB830Fh+m2kCWdUzwWcKoiGsgSSd8ADgHM8glXm5Nm5QcxDjj
qcf1liyC+AZ8u5qjmCHHt5ThAoHSXf9hUnZUx9eiN569R25DHoymK78c2/BK
X4qDtDUd9KPQCLITldy7WaLMDUkxE+ObNJTM3YTLD2XoE41Cnz46mYUd305e
ZVlTfvOpnznE+Rq9hfTWI8lvK/LUwwms6+u09wPmhdh338GJYpcwGx4bjT6v
bUZsX9ZzjsYGq9+g7C4CooSBmdH/TsVeqXm8U8DBcz/qglqc1R3+q0S1Nqtq
GD2RQh8LofrWT2R+8MM4TfcpUbZ7SGXgEpKYEeWwfO62dzCUD7nJ+HcIFF6w
HPcGvmmNdfS1yCLLwT7jmU4gL6x3NH0edhcLPPE7va3EG48BMGhrCbjq0pUo
AVwUndKx7JWlLDQCvxtzxSjQi5XPz9E7as3oE0KJKonSOM7YV9jjt2bmqVsx
w1Y0mnvy0sY2lNkphSIeLuJzA1lA+a5vPQrf3jY7TnLZiLKQdLnCAn3PUHBX
H8OhaXg6Jtq+Nq88nzVDUS02WOxltbNS+mna9gZmvByQ3BmTpvdHM8jMb3KC
9dwQSkgdu3Tnfoauc2TOaQLK4+WU3gO3s9yOWnWjZcy5KPKcktlO4qvlO47S
2C+ub+VN8Cw1Yxb2R1LZX0JeOHkF/IQx0zl2mbtfy8CDM4w8x8lV3ByvD04a
EWAd8NfshywbnyRBQdZMdIwGOKNMdNHQd2K4mnZQagVTSo60WJVjg7pG+weJ
5a6JSDamOGiDc1n+oJuEXTF4Mj6dqFkB5bHz33UCQUugSbPZOH3wRZXKDoK3
sT+z4GYoforahn6jeNWiQxxR+HoW3zvQRt789XVdouNg2vjAj8C7I7LhzGet
VgwfREwm2XqcfQptnhWf17tbAc41SBBA6A4WeOmEGCu3PaodTJ1mkmcLJOUV
uxzUcJ0hfb9awz1lsvVPmSLLgH6Lq/WDDG2vGXRj/qvx/b924jBkyENLDRHb
brBEknjY7cI3gLRjC3c3tjiLU7fcmlFX9vZfERUd87rostWCGP+Sv+aLE5QJ
rBUtWCHMtpfnXm+QqaUDJanO74tdoLuwJS6m8TAjIB3lB3vVywXQFz2S+ZuG
5L3jSQF7p8rrUANiFUFYm2JagjguVTdYWXpS1XedAgsLEq2MWCg8AOaWHE3p
7oELE6fHlxYzft5fpqnYtMpzNAqgLJQ1e1V+Mf4Dg1+Ewbsg7rx7FTRjdJj7
FAoYs/Wa6WSV047wNBWZ+J7z+7gF3TKvDvru5RvC3JwhZ8Li65X2ZZQhWQhw
Uki+hhLJzrZBYgqH+Ax6T5GXZx73cGOQebybfDBMYbuE9Fbd9/1jztXXSr1N
yR5dphJL3ijGO/RqsHoMOLT15I1kmAHTLqby7ccUjkbd8XZHmAI8f/fRxowQ
kIupKnebEoSyvwOfv6zJIdSfe4UW+JSHlbymjxAPPqADaKVajBaj1/vpBMlr
K9lc8MyuEOxlLMPDlxNFOaZNwerwwKPhXVRIY1PslbIIZDo4xj08HoUEikGm
pImR8ooHUGXrCv1kIgDucm5Yddn/D5OQFieYcIxc5Dm6r6i2sdMKa75jxo1b
5bAVBkLjPNcQzBAN5Nnb9zLsndYeMVPvBGXuunY9vpLm2nPphO0iEkAYXsXB
liZD0MlpvUvzdcymwcEJ2ytP4K/tWHl2qzekUkvgzdDv4dZT06rXHENeoetZ
9NDXLpwIFfxXaQMkHSCGSU+pVip/xLfDPVZgTDKt5axY3YxiwLN9QVHM4AcR
iDqfrtrBekAKfj5VvA9dpBpVLV38MDmCK8deFkIRlNIdqZDMGtVOx8smaKY+
DMnzSFukjGJ+fnA2mUYgoQN5J4WYxdufShA+Wf1rYnZ51Be3oshJNKM2o6zZ
nqOGtruJBJMH1JIDd1OWkzF4QwYH8MHvZ075/EdTaib/4ZV9kwL944eNC4cG
ESZpq2MqTW/nBBdXlKHgKpm8C0JEuWb/X9bN5cl1/2kFeFOHkPrj07gjAGxH
LkRYJcHpqyN9vmFtQF2CVJID75vE3KmTggNMuKUHI3b/AS6vBc4y/AMR7NI0
8Bi3avX2DnJ0L6/csXsFlazGWZnjdI2uywQjpFfD78TxOgGwXlB1vWIBIsaj
9qigIzhZOasu97b7YAHUnwqAvrdkEeaBlJhj0sdZ7C1sN+vwIGE7Y3okpoCo
RHbSXQc17GLn3JrObuF1cCYqza2dTqePc3+0dapTddvXcYFgV/oIgr7g8KS7
6mpPTGZXxKp8T8Xa/c/OoyvWukhSB8gVRT4419N6v+gBS1RH5urwWuKK2HrT
9FZIZ+2Vsj7sb2wf+12lQhL7SP7bPo5ivhgiIba5m+URYMPast9qlZRUhf9T
0hEPQBraoCIGnZX35SFtLnwA2lzoO+MT8gquMCzo3iscosROBDkQZRmVhBez
jijEmKlyE+L2kFc3kXGNMCx+HqT2O1NL0TSqx05XpgUXyBNn5L6y/5gUChTq
6z78BivGKDa4WqtkH3h6JBPf9xNhfhD5k392Zsqx8sGSV5UhLrDx8DU3tdT4
zyjZCKlNnAYtyU+TsSWN8ogI2OyyOn8dC5kmAlYCzt0vO4Ab8bg5XNbv24es
ONHIMq0lNvWy2HTvr05pFX0GSi7U49crvJjXW2z/m/17l7j81Q1zQQoQF3Cq
Gl/YRSSIp5pdWeWFyreueROX6jKvUUiUu+6Hya+GTuZNeZfe9SqJz57PQEY9
IZJYMQY6AgOtyKsajbYEMVh+0tf4iNqXUNMB3L/GsHQLwb9OAdRcLD0pfL3h
WwA8AJyF2K4eiTMQhhSJuUXgEVy1pzHbqy5iAYuPHbaXFDX15/u11RYdGAAZ
C8qYrWylOHmqSqfwVoHTdT/1Hcdi53NB4LYuzAC0vGPC8TLNjuo1AiqFAYCi
byglHDrkYZir/KO0gCsjrdtUSEGtsZSmeXmRR2UwYXITza9LN6gYyEkvEt5h
yELD5lQXkTFOXTUBdfH7Eqsem9xl339y6b6ABP2yXRNYjDBggRqicfGzScx0
jcOgwlSj/bFmme6QKRkFQxqgkuaj6rOG5B+iRlO9yyo9AYNTQTJwicnLzeSx
tnKtzu6iveBNVepDtZ4ZHfi0G6wMBeb45EVe9nLNmazWC6sEmRpk8r6jCv9x
m+RRsWnZ/gs0Wh8v03KBDdUflYQNLMkNKvvwx/7STmEH+8G8S2eBbO8jFpdg
ih52OP/oXhwblj8N23EIj/WVLQcBr1SlzRxp8tXv/ibekuvX79DQP3Zn/qqO
Qx7MPZNhYzG8LxYydPtp0JfuRZkHNj6cqFwb7TOxSG7qoAfpdQ/geu/0Ak2d
j98ks6Lg+bi4Sjm/siosUcKwIAOF5NcPd+7Tajounjrr55/OIiTErX0raSfj
FfXcCmiV68UaaW9UiHEtJxPIEwRCDGc9JlxrWL6eUS79ac+k++XpY3wvnzOI
fKnhHkOUVWO3ubaj5izuvC56iiVTaDqgLVuWgzw9c6oplDYKvJJ3+rjbAbY+
J+kXsRFd9/wwxB1VomQluSbZgjsg1/mWQWrNjz7+v8Lt6eXXKy5novlrJX6M
73fWJYOAwMH8JmE5S7e17E0xGxTYXRrItpFCx1Jobm0O1wOlCJjDnQ+pHlFF
dM3b1M9iTVw/coP4zy9F7SC8+55OPtu85tOfcO9aPhr6Ce/MwgvnnzFUfY3d
/hNANHuGsD3nA1suY4lOKcFFsX+klarQ/9+/QAU7as4xNypI6Xyy/DkruzXC
kdd4WXt7AWKQZZgaVzP7RYleErBOxhVvR8ABa/PCxtxQYgMJggaskg7H1Y9O
ybZ7joPn8QEInMkA1ke7Jb2+Bqi0ZeMLhwX+0hFh0kwh5s+EZsPZZD0iU9l8
DH2MSSBddTxpZ2ig1NqfBESA5gbVhuLzkXsPULnSvftniJEI070g+8JkXCBI
WfqOFxpQzBMqw+r+IivWJFjCQ/VH+jpQ7O41Ke42lkrUNt9+LuoLIrMu+V0N
WHGqMUEt835OGBUEdzusTFC1qjEQfMsnEYhMIh89YrxY16g5k5vP8L5iJ3yE
hcQWVmvBplT9MIB1sis70A3xGCHYhJaVvKE5w9U7qajBEDeBh13AtayGGuRY
Q3Z6g4c++eeCmhf6XDvLf/MrE3a1uIutlcPpVp2ZPp+uf9tB9LUMdiPkgCT4
TaBrQg77kaZU2xbm9rZc+hpYdKJfENQ30vWq5DYcZl3OQHniN9c3/MUFw3SZ
okF3MlqqHUXAnUc1SW6rHmz+qRA5UzVv8X0xRVrXaCzWxHiEleWEibMJFcME
zSgDgOC6SnBatPSBXIyKqeGX5IkXBsuYwfzWjoPuGybNQZ3KpByjmXvUP8wv
thKtAUFkgoY1LkA324F4jXI7MUSSe6SVgM0upC8lOgouQkoggkSSF9Grnqrq
+GcKPhO5cGU+4cq2UkHMhdLMcN2TySDdY6qhKgMXw0XYZiwDqAHys7fgCzua
O9leRvmdXD5P2sBotDPahhu9zJ6CjWkMvSKzIRtzErlbiaIWukRRnhiZ8xXI
hdfyEWfaJefpJRprNoClFrlBrx4KU1QImSRdecfz8kzTLNpb52HZ50cwB9Fn
lkQAFgoZAwmblS/F4W0r8aiK5geAAmHfUPDYQByns1REU2JR/2yRXKvf8BMN
osGe7vwDDe324JMhHhMA9cFNFz9Zb+JFjnDTnAueTosqnuKcb0DeMQeZ05Aj
/ZSPRZ9DNmfDraC5xXYkF4AiZ3Q4HHRtJu8MlI/zWEa1ZwEcdbaMlpCtG3Cx
IXdZDDO3QBiGx5vznw5jzZA9BDf5meBxogapBf/k1AHnnU89m7OkL8VJiC7L
WA6YiDDrOjH3Sd7EnzT4iKgeevoCRRjf6uopXWX+/pTYYJ2RW0Q2lvOWp1Cx
Pj+znX9PG8EviFRUV0vRIxJ16gJBvYHzzQW+JXc/CNJG9UM3LT3w2NeX6/Dc
HmohxnIyMaXc0TANcYeCrVVQgY9QLw/UIYPFJinwtmqtPvw25fneQuyWn1Zv
artzbvf4N5XInbGkHAanBVTpB6c1Gq46ZAMn+eU2VucNJCAlS9+EYM9Djwgt
JsZi1Ja9mdQ+xSQm9woasVAeGqNOBa1B5gEKdLXNVjwrBYGQRKYVc836yiwU
vJzZYcXF9xhqLIx48L0e8EZ7+xg7lQwnBKXtFQ5fSaSO4loMXvLxAP5ZXs34
E+wiDZw9qrT790V6mW6IHiBSONq987A76rdQ4YT1yOWlrZent3XgPSw2QpTv
elb9+C2Eym3bZ1g9J9YYmAegwkvJlfKPIMhNrfP80H3ZZic33A5l69Wr5Yxy
1nncVZGNH9koTGRIN6q7vcv6Pp5ONRIOOsnK+Qi/6W9maMtPCMhT9WgBbOVU
P64ZIiTAs0GcU1ksD8oiV1JC8ZBKfOTqMJaSERyiU0azQJlW4LlH4enbp4Pe
IpXoay5sCoaFZIUBT0+GuYO3cywVe3Qqzjyw0tk0nU6BLmUwyswcbcC4inCG
WSpF6kuZdBd3Iv8py882yvmgLwvp5eF+UieFFPf5vISKQwjLA8x/rbU48MaE
2KemI918gu7r1DvbrK4bW0qIpwAJhHasm2kLoygccU6mYR5ckTLlb0MK3PE2
FDCdsHx//G7oZ/yGnyw4f1lBmxjojJCs+Wcmeq4789Tvu09dYBO0wOiQsa7E
zoZE7Ap3hqvonSChBDvcHm/VG5Agn+sFZy5Kp71zSelVz7U+8jE3YzF2nA8p
Nb8lAgqdemaBaTNjTMDp2pmS3a7KHFuPbVgNeoYpO8kq8rd+kt8J6xs42ZrK
+he4X1pXsow8xxOqZDZ//7ZOVZCyI5d8AZK034PYx9LX0GZ0cEAjUyxnIbaG
RMrHDvlndtCN5mxsFZin3ebCx4M3loNHpCN4bKn1PWP1i/M4SHDUyLfEdOcA
fxvEPhTmtR7zTN+8i6nZBKlv75GgL5x7pyP12WFp9u8BNuDdx/kdDAFtqrEn
g9LKh6X6HuEIjjnmdsXXerh2RpqTSHcz7h89g1k/EDNrF33ITzfVePelKK+k
HT/zyCvDasZV9kIr0o7GuzeBL50bdIrt48osZ4QqGcTrj4LLaP0W44StQ925
elk8nNUAP4eMpG85dONu/llT4ZwgRWJKYYd/u+3clwizz77Ls9beOEf1H/v0
kOPnfYw/JaRrphL0ykUwOC6nRjtlyhWwuzx9ve1vAKfWpU8cef+kq+7Exk8C
7cfEqGSQ3V4MDf9CMhqqWa8LzwJ2MdSjKuj/l6iSxbdXBCXPTxaC0mMUtJcB
+BC9JkxRafMlIxeSy9oRmbFhRBUZ/grPu4T5JpAPsDcv/GSHV35nQp0VlZ9w
42AHVGk+GegU3nFJOlpGf1KSUuVQrMyPbUoDNvvpnm3J6UgAdNXKtsE6B8mA
q1alDIBnGj8GmBq6qvyniOHtGEQtW6V8Woa/DK9yJXAp8XSETTOV1hojYlEk
unqYa3O+BzArnue2k5Ajht/GIMO7kzgb6mWyv2IGd0XkpMXN3RcFkbaPqDWF
ZphMCvXR9qgHpIoWAo0u5nxj1/MKpV82U+ZR7Ry4DvcuQQs9zB2VTsmaBBEb
eBxZGwfXotGCUTx8zcaqTHroSonAGXzMrhRrWQymT9uLzap1ULGEZF4gDtnB
ahP567mB6sOFy6sfjessRfs2jh1TXI+QoIqLtn0Xkf7bkYzmnTgFiRxtHtJs
hITgeYTnalsc/hX7BC1W//9xpbP04NLmtns3R3QYC2iIVtjlS9URO6i3fTpH
OI9ZmhG3NvV9rrlcdgE02TXFcC/nHsSOZcgD1LSpBthgQl/TKoFqnfCV4Mmb
p1y8dVUBO6g6YZUzGrxui+L7MkShb5ghGeLqvirYmaFiE+NuBxMVr6NMNuTs
AzQv9tsRXqi0zLl76O0FVe1L7GEnnK0RZ1eEQ3TI8mLfs7eki0Tfo4xsMFxV
XDEpmEC2SczyFAbXA4Zt2pKEnQd8JCM/5HNX0YsPq7DrL5ueUVzYmAE/IRHH
xvPS/XGCPuvZhMes7d0kJm59J0eWTYB/ZWqsFaw8f8Khww0vkqKOmiHPEzOp
YpbafQG3zX7h/bdwu6h4khVRtiv8pydlyCd84JBAARHr1Mf12npYSUZXvHkp
ML9+NnG2ESE8yJVROa+ozaXWPr21nAp+ptmQF9fY4dQtddVvxFcj5WvS6OdK
FbCv/Q+VhSEVZrdGtX8TWh6ucbOp8BbZmM1G1wgLMIYsOTL2m0QRY98LYr28
E41KshTp4C18kmuqa6zXSFnWo2fzEsUM1JG6zUd7wQw/8b0jDhvPj/wefRi+
x/IJ5fGZ6Sot2gOtGR72jd4JFCIXSlzDD3UiqhN48PWOzUCLm+fzqmBqkkE6
fE2H4T7mgwLLfg8hspHAI0RluTnInPcjguUODwVH1TosrgYYV9COtkIvPtsb
KnGW57e/BRg1Pbxo8A/7HUATFbxvMMWhwsX7DDrkQVHb4xs5QueBRgDT6CCc
xZPTLbTwciHLWTBdcoakvfuAG2PO7OR/77P1nQlp1f9F25Fgv0mrj6Efb2c5
iMYLAfmnKy5f49NtJ8gNKY6xWVC+oAMWK9w/TatVA6rL35I6rYtDOJz5rCQ/
seyI

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzcxyCWCyzznCnuSfBwpKrkg8TiSCoB5ytvmbwHay4aXhzYHFam/usaKtf+xqbx99NA9xasTv1eqcv9wCXUWFv5dY0S0AI/c0W1KwA+wwBwHmtu//N68GZ0jdAYn3Tndv3bLv9qOiGqvVaxMBYLN18jZfm/pIiwq3rCpfnhSyQWkE2AH+dn0FjvQzl6cPMmdVLpsjbnfY1rJBilQ/zyP+bbuzx4obs0lP40lzxRNFgrToPkhmhVBahhrchR9FMCM3rr3i37KmWcyaASM5lmL4XgdDbV0crz6udw+nrFowcWgOq72wuDX7jgAH1EzICkIqL4+Vbw975TxLPiaR7fEoM/a4IstuoRLdX5Oo5UcgoimH7w9WuNV5SX4flwmhAImL5ha1uyESp0qbVoshHW7A/Jr2BykTeBoI9EllJtTA+h0V7QnM64fGKZGJcE6HKw06i9Drh2BK6SV0HWOM6M/v+Nlo4rKH0TdjOSVQRkvIibOuDZKooChLJj9rixXNOVl83IK36J6hi3RQyk2jzGyEclW0hzY3KyzWwPZGw0XC0TRmd9h8Sjr7cH2REg9JGdsKKkgmjkhxE+hzOML+MdDaHt4Prslqs9Rbw8ZL1XKNGjGMXKLfyrE6sAbIJX0BX9d6ovLz1dDSXnUunbHYpWdQh2bAwfpx9wZHx6iUX/HmGtpXdRF26U+dAswePMmCjpyWT76HrLay3btYvMdVORizYCiJIu6YOhLuT/qAuC62z26TtMf5DQBpkRMi/kJXKVpufXvPe8vyyB++qysR/qRPUQG"
`endif