// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dOA6ddEOhRa6A69qA4nhCRgHqTYG1t0wIudRAETSLpqrsiZfh4nO9vtI6Rrl
MxhwBerTvb+iuOT/t5E1ypv4yo+RpzpEERaU+4V3EKLutktX5RbIkBmFgiDb
/Fo0TkbxRccm7KJhrGxSWLMxcYURk9wHrEMzlPdkO3hiRPDK0IF/1p84vVyd
gg4s9iOk9EyfsyKpoMDqqv3iC6xvIH7o7CNtKaPnofPy001b+YPK6Wxam3UT
vJE94BeUu1DQq7L0aLgNv5NyUja3gI2Wrv0y14qsojpinqmY2Em1mEhM5PY4
n4xNcRbFpi2G8WXyCcyf8p+i/D4HvXsQQ9Ez1T+JTQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QBnyKToz38dqDWtOO3ombrLYIPfPsQOjppaGiifX9OnRTV6u3zbuyg8v44wD
xU+iJr2494+YGoDp7N0Nqh/8QpoVZ2tIZGDQpMZglgpD4SmJfXzLFLDneGnT
g9fYI6dHW+EU1QyNO7GThNHdqOXe4k5tVgL8qt/IAMlcVRZI5DQQ811GVPj9
nNiQWd5Svs26dwTBnUiMQn6HYq0Efxf//19zqgW1gxuCX0R11FFMnxtz6RhZ
+AhDAfdE0o+zO9yJnBs0TGSw2mXxtZkUMSrIEpWfo2UxlAgmHmEB/hOXHTX9
xzR3NrsxA3/GqIYsxdvrXP/Dj+479bS9Tk00P34h7A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DP9DE5zkKqLkR9+KnzJceuCcDejVlC8MoU7JmSdbEaP/7qxbujmzT6hi3Ipc
LaqMahTcOflDEpg0XjFLWc26HcsYGT5b9DCABnRkdnhX+cSU3MxozuV+hAYO
owMScfmfb3mUuh4tHacQl1yNYDoRhmmMc2aNHmfumO6Yyfo4yOmcTs/FKelg
IMOfC6R2vGyMr2gCMUIIfCDGJDXgcbhRBqgY/hpTdFoUn5HSn8Vq10r2u2+m
mCvorNm+tJ0bf7oCkyjazCIOW9nc0lPv+DemV0HQw9GtfD1bFsxEwTuoeiW2
dsHfgUPDI/LSYMe7kHs24vGcmlOa0MUi6R6yDxQ3zg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NkfeMlu47LWaVJSjGfyWb+WRJcPhf+elA+Gy5gjl+bf0Q2j1Xy8jj3hZ0z4D
BxyPMBaWdbeVz5DQ5ooscKknLQ3Dv7vKAvVBfmVqdk2lSZvMkeJIdNHSY9Z7
GkjNufOj/XcU9q0PRxH3CHYvLTzTr9cJu3RnhXaMt4dcl5T/jcXQE+kaEtUU
w4BNYL/KigTU1XtD/9S/L8RXD9te6JqSipy06IE1QKGeBZwusc03MciwgKBk
K12uS9FHoeeDtjlVI9mWkQIxz0sb7mNW6XC8KLkZsu+0kZMXG05FRjmPARgc
TtIgDltcDAIhCN0vUN+vJDlHKTyaVb/faXCBwrp3Xg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FmdYNCXpxKCnmzYr8gy6OpHWacsUUsBZ2AL7ns5HOUp+OMAlCawue8Kml/2A
2YWkxgiVzn5QvpgoMEQL6UBl5CbHqmoXdJ04cHxOWSVqYy87TqPcQKnE5Ziv
FLI8nlIjtmO0d0sPkgVczOukKw8Mhd+fgP1BX9BiHcLCAfg5UQA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GXUSLwMpV7ZiBbHLMlOwrCAlfSBJDP/pbcjgSYlK0G1Wo7ITVHF46OfxoC6Q
UWuVeODKyA/rE6bkAsPrfFzdYclsKYEW4J0vPEVV9b6jRWDU8OVXeLeWh8Dx
IP/n3rGxk56VSf2MaVBxHTMZ/5euS7EmevV1C8s/1XiVweyR/YILmEAFqkeT
tWGmYZI5bKefuHWVGNA5SEg+Lph/l7ZA67fcrZhI01CFdXPKn86anOlql4JH
vjW6trJ9ibhvLC08i1UZsNAR0uoeHmzTEiEc6gVTTWGfCej3bnO7Um5buEQA
193/Sv8/xAugOzrRIO+sU6Y/gC61tcZcJTjFd9sC3x/vDABPs/ApWiOsTS+5
SH710Sd59Qu2lde/sgFNGTIeLaQmZJ6enXXNIeb93UcsxcH9N66A8ZaaiDgq
LP3t58CDikYPIN83eIyEQGsK8TApBXndkF5mXIAX0x1K9L19E6TjD174U/4k
tDO01ccS7WRh7UUBhAyKMjiv9yPd/Hdq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MwkszvJ3lRWFGWHembT9XWmAHF3cMP1Dn/17ywGjSZRxpAsnnGEx2Tu5vskJ
MilV7NLgR1wnEGlaLIX42n18ed+pkmQaQbXsRnT75KEV2V/dWd6Dl3WDk8/a
GcDoUWP10Kz/GvI00mTqlTMSX1V6qWKH+t4qgGl2/9HUnv5VxW4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
prnRxf5oVhSFEH0VxqCRzozy8xJ/JcdmFaG9kXdjTe/fkSRDn4IhShHqqvJB
cq6U6uVAZLvo+fe5p//wpokhcFbl/q5dF/i6YwHMyDUAlUHG9Fz7kbsp8Vj4
S9ZNo/BR6+M3hHTH7elNeDYfsv7KyPx41VRJ9Q7F9IlMa1mbGo8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 22160)
`pragma protect data_block
aHpawG25q5Qw35v1t+tbPUZKmTropKybyQtzjhs9+YOpnUlS3dktSycvy92r
FoBheXoqcjDmQ2skERotHgV8VdHia1vTdXxIft/tN85T/TZiRdR/3cW5jZ11
GwuDfLpPiR7+odSh7gm6XjWnQMyMOFqMTzhnFHg6/h7jyiCcfqY2g2AG60vX
N6PbNsK2O9KDrVkGNbvfuH5GZ6w0WNlYz1QgRm2uuhYUdnLlEoOdUAaQUziQ
IGxtMEpTlDMt0tpI8iK5UZ8r/AGZEFP7Q7IHW6+M2M5XtUnDXP/jo64BbG2i
x8KWQIGRp9VDOVAZjNZilmZYss12KVKXJRPPAdN0scp3zWvxkt2aFihXQ9dZ
FbdqfTCgVOA+jYYq4kgD2tkGDhafGoD2SINu5oF2ejynRQ750KQaSVhBQH4h
F/8E450YXUqsHLWhIZnQo4Q+7MZZ04eOxgCkBwekN7ezMHbIkySANndEnUOJ
3Q/O6LyLjesXWNvJFF+lrqzMOfxke4ILITD0HgRJBF4b9pxrRZSsX2HCZnz2
KY3CewXYb5mnC6kVINer6xnScHFKFPty8FGCOj3KOLvXQROeAT2kbrbM8JRs
B/R/qwoHOqVwdTRocfj5mPYLvPvX3JpyCilBW0tQoPVuzo0kvaodo6QZrJBz
NuZVmxpFgDxihRfZYwJ1+7WnCiEOYmbfhAkhEABRs7m+fg9LYzyn094vaeJX
wPOZ1nyMY/445X8s3msSfN/6JnTb0LiO6gi3ALODoVWcQtyfdGWFNBighEUz
Q1ZOpzjxyZ3ki6bIGSo9uVQj63a04wXm86hcDfW+LOVEXJk2QVoz5gy61op+
xFT37M8VhzrTfe8FIBlXcPCRjVRlp9fJYCvoZVud8q91Wv7uK807uVDhyVMD
hJPcGjRBw6X1o3kf8UxjQjWKAVkj8/oHCCWOxtj8PS3Wl8reaYqTltyN5K6F
d4SAfqar2Bsv1aX5QvMifvC+6TyazoHj4z9Tg/Touax+OIOaNICHQ79Meiql
xibHQrmAeRD9mF88yHmtQvFyzZkXM+5i9SJZMtFgQy834qpqeKLt8zsP1R6n
gUi93LoWBDpGKxclMrnQe0cN+N8QHjNkTqJ50zfqgoA8TcvbGoVvtrP9+TE2
ru0iH89BCxWoZG3KYGgGPMAe7xZMXS/ZE+r5vXwKYXRkxWFa8dqZmVU3OTTt
kxFpcl8owhGKnW6T35QBomAJmGXa3TNuL+uNwoijVwoXfqz4EEGSL38A+YP3
uBvf4OBi4HcS/P7//KL0bsw1XAyA89ZcznsMhq7ZF6X4pIFnyqkTQLxlWSP+
xVa8aNWw+fnRfcwhwk4pHTt6rDRJEBJ8/2Ju7fIVIpXPLTIoqjbU1xVzVliJ
aHsrCkuXhfFwRMPpYVmVmyWtUrI2F1q3fm7s92E/ioKlxOeibjw/lIid/OYg
R1+nB0dkDfpHX/F5M9ZI17j1q94nIRfnYWolqoBxyuc7Ml+dmRCtFjBVnFo2
WyE5bYKHIPIMMQZQ5NR4PgirTMi4wHw6RADxhu5PVVfjbMfTfA/i/fTnoZdZ
CJzK5eSZ229rW35cAZM4d0LTz1v5ycWddgjjAnEMzW6gkGWbkBe2Uog4Ll/F
2N8lHGovBXNOew9EVhhG2JsKipRBNeymttFa6X0Ik5JiXYjXRRI/xHIGsqch
CyL7akj6xCpC7WyIjDZatqDHbMUwnq8a+w2dseVuFgM9wEZsqa5fPLyVDnOy
Tr2IqcV2InUDB4P09vyidT1WcefiO4k4E6sZikeu39VxgWuHJ2khYfuXt8ok
dJrSEkx3wDqjmMUVPhjvHssTbbssVquRZseXlmkcto6452N1s29b9bf5rJIz
w4W046ZBTPpQFhg1dn7Ih05J94kMzTU2LU6VV+BG11QU41kWv2TGdAI03NQs
v27LecypNIfXlK9WcmWPl6XYUfvWXc7keayfnz8rHsaCwEiV21NSfcEygEyw
8DyZjypEbGFMJv4FFgJOBPTS96w/vBbv2sdQrVrHbYJUG/LZNbcfqr8KhcLr
upR095lwc44XW3t0RDsjPT6TW8Pq1MChIUt4JFAHpoGLEagdWaQoyHAAl8uV
t8mnm89yPxgfnoLLn2+w0UnKjZAbtJtA/fSE3/BwJMQVLhdDclv9vzsXMbo3
TfWK28IoGJ0A67vcve4HlYTFK3Qkc3h/GhQXXtC+kJ9rxktzOfNpJqLbladu
EzJBkAsdnYarqGHdGIbZGGROeJCaT61hveN2PmILH+ZxFXZvPxiWmZlmG3yr
4173Ud6uglL5zmyeWbwClqJdQSVGk4PitM6Lsz5HOFfg0z0diTfV2UtH0V04
yqgndDdEr7Wv6o9oDHzlEws9+A4PM8NOT90p1GHdnG6SO9r12MEzhU1e7n8W
CM+d9Ixcap0a4OMklS6SwG6tVzaUIlLUxpWOhIhDDNOduCtyMtuzc3K3VbNg
rDy3tLoKH2g96Gl843rvYdLsI/Jw1AjMA5D01j8m5h2lRea3MoNB6w1WM1TM
TrT7LlKrulLAa6E+txlXpGN3CQwTHKX6fNPcT4inRiYfqOVN3qEbhueSXUOW
cSDVJmnhXPEb3HlauEQoevsFjeUwR89VhhM1bkytaZdrlvo10jVI5ElPk/Mn
lEwZTWCVfJ6Delm9AhYGfduBxUxhTTaX/KxrNgWinxCGoJ2Zkeg1Z87VlN6w
Fs6paSsTLtIOknoIt1Zl/XtKExVNEh4tW3M4VUidpZ7BuzCGjojHB4EC0IaA
ADZRx6Hjb+P/lJTRlwA8EMTUrJABAJjJsJS8AjP9pkhyLaj2uvdbhCt6mCwn
fR1Eak2oN45V5cCQRSaNS0dU6uQFkPd6lvXragV+Eitiezs5PgDlAhkb+xiT
COpwHtSuQ4YRk1xeR3pi8e9ItbgYvJmNZmBZdKqhOKjPqZxpCDz3pjDYKhyd
XYPMNWxZKIadjuqLTeC8vFem3F+JEBA3o5remNKFCrXY+h83DufBVdgk2dnU
DxnxdJ0tSwUXFLwo6hkmYO3chMtVVtn4YF5km1vHrpcP4h2Ib8xXqxjWuMFm
ifvDAEiiTF7OOla583nVuvNtXh4rc9VJqeib4HERAKC/TlN7O9gm1/f+nM3g
VHPiBBlq5RA4APM/V1FKfjfx4N9G5z8PiOqbi4a7Vle9xaB+2lBtTsIx49uG
W7wzTyc3FL255OZzKXeS9vlZcxeVZUuD1QHLuDvq0BRUXGQ+X5gUxgP6WbXX
tZcXYMnKGdvNBrKqoivcOlfHiUCMYndcDEIq/pdfQZ/xjvfU1ejZW7vF4GJQ
/TpfKPh2SR/ftE/Cz2ArvS/3AaeEV2aX11JOnxI83YuUia7R5DnE4OBxqCo9
4NcJAT+VJUCCreQorpzejYwp4buf/bLtEY/ShFXElvs4WyOjESy4LbSOwxXs
3n5BCU9yc8nSd+5g7SOsv9tel/Bk09y3IU1C1pXlSn8lBWA0wu59zPuK5e0e
FZhxoWborXv0qy+fvW6DWMat6y+MNUfpsccFKHpod8lSAGaQrOEaqPLYd6WE
nFUA/fbl846hxpaHRe1jshkAxocD9hRFfNPeN5K7PWy06QYgiyPCFypnB1ed
ZjQD7akeKmcalH/I2+Xd3FDXeZxaqB789hCUSEJyyopRqkb2iRtjSzeHi5zj
S7mrn4+tXHHL6ZinSCsKM6eJmmOFxRsVT0m9FLkquUMZP+pnJnPY7ZK2rJbQ
L1qnEXKMn2X8hJM73E8gyq96HR6sQtQzoXtIFz7nqACCcJriwGp299M4xxYg
fKZuc/h7Qtt3mzkBxkti7msM8XAlqWP8cFlLkkk3wsoDFO7cyDjBSpl1a6HG
1dJbgNkME+hzdx9mRPTepu/QPmt4cCIF2Z7U+I+hWjpDbcCO8ZSF2h1r+ouu
tfGiCXJVpNkBIHKTzPeRPoYntAVUMwnc7bt1iR+dmwiLFDPdVFq8x8aM3DQU
dobe7stH8CJTW+Mmpd+a028bqntoOEhCTbgUXNTekK8LwWYWuycNAGaplhKP
UuR4Gmk/vn6E9DXL0s6avT7huB6XEQ7UGkWkzdvhNPqvNaWk3jBtPFpfnpCe
+4HsdbkwNjhitNb0SOFHs/FzbsGw6zz5KMCmpHebKP/hmuCPTuxK2X7iXu5G
jdg0AlOfh5VCp4SqFRXorko9Xyr1wd2LczW5AM2RS6gyYPIB/vl+NSjCSuZf
/faRp/shb8sVYgW4Mi9Y48HUoBSDlvaP8siTu8s9RLj09KL4E4U/04MldcKm
dTWN3cXRVQCNAqTjHmkT6G8GVqkHYD2D13lw8I0ThO4E/YuZ2CtZF8qQHobI
L0h75sH90Nf4ID4YWNgGlEsgz6DPp4nZIzs7bEBpn8B7uDf2VpO3Fof/xk6m
jV+Kga/j+dO2qI44p9g+V99qo8J07LleW25vEmfNs2THMXOLUXdBIOiXxo6s
mtPVn3r7EDeAB3uAzS5CMYs1czWKfHQseiGBKyMx1D4w+KOumESAlJCrQlaO
9/c6jllnGLNWQWu4cxl1TQtq49vba0uxfFIJdum6NvDvRFXtaAQzs2Q2t+Q7
GsfXW+8XTQBvoWs0+o10IAy03d5AGL1BAPjlsg6anZQ+tGdjN83UAy9eYt23
cpSejW5vPK37VwbjROrn8+tPv8xmKDdorlSxy41tCkBdmrJvIc6lDQW39jxr
5XFakyLudoNRWZfakmTJL0W7yZdKj1kYZlsT0v1qA6tw0fg8MrWpkiMVglAC
TxG6rfQfVE/FvkcbnLsSY+YBOr0y91kQN5iH7VFw30vFHwCvbKE+U8E4bgV1
Xcm8WNCPoWzTZPyEp0Br7iHaQbXFUS+Ng2f7oQvgfi49db752siymWwWiOoG
8qaHuOjBUxETE0UnHs5OBUOSN3nef4YQ5cGkrsTyMsLkOqZXNBK44pt5ukF+
9RgL9+f9JE1iDf7bPe2Z3XiVs/lnXBwd9c1gCFrs9VvttsBbGfYKdxdZlbPF
S1x76XYz1Q8R6gIeemy2/JFymJG1pyVlfyXHI9ROTRb1SWzk/lPXpYoCdspo
2xk3UpFWgS8Qls1pgEWSqWYBBOkW92qqW+WSTCusA0JPjMdOxhsiCuEvnd+5
IYnoQ1qIgR4khfQBxqkR9x+p/Z6czFaVT+khZBwj2ci42m+28c8sa8PylIzK
YMp92HcHd+ZwFcFIcErRlqwA6iJ7mal/VyfzzzVP0ThhLNJn/f3qEww5P3E2
4XTCeOJ2wWJ1z24V/38Zpvkzs8G9pc7yXL+3hWMrDNjO2CyZM4Rmfnad37Ji
0qPVtRE3dzPYBg5flOh7iYJ1NYhhh83UsEgAmiIaAFkvfZ5WSkdZ3tI895jN
HEbBXqBof1LuIJPL5WaaubuZG9so5LqbwmlB3WY/XGktlIblZMJEe96MjUkt
okM0mXouJcogBXpntQ5dVCoVPscZwHqH0mKw+ZEwEiv2g+8CF7sANzOTPk7a
7+RX1m9VAINHWl4LKg2/ptwefRtuyDGuCvQUe2abjAjpqKfKtAcNiLZPk/S/
OVI4SeTkI69sXa4I07NDclrHpfHEBTNgvm5EUYGb3bEw/mP8N5PRQyAE2maB
p6tCHtGzJFAKlqsa9dM8rqdJxTdCJGUQda6S9vDe1/GxYYeyQS1M3bKi8mNt
/24WzozOCEiGDO0I3ZMLiziiXhE9Ca+N+yq4GhZhviahVeoUMjcRbe2uRiwk
zpDKd8MgCdzqHO/nMR5M7qQjZLxsbMrVrasDYmd69bzMlKPdRzcQszTsHU0t
cL6RKApIqLSU2Wqppg1pT85nAOaM9QMEUPhay/1cxL3dFP3NGYLKqjJFUCzz
VlW7IXc3LTtX2T5M6AlhKZzTIEuVEa4Bm6TMWTk4QpuGknRxUXYrP315Aaq0
w2+kSpec4KrygThnAd6u0k8bTcsdAfTmDeugcgr7Y/zylWnpHUz/Wsok6ckF
vVeUboZ+7uqOk/M+HS3re1ZDoq5lzwFMB5F/C8wG7+8YUquGQ0nE9Bpwqq0o
fgJ20zpJqW55cimmd1e7Up6JnifdYUtOyInmgnRCK/6kPhvCWeHvFErX0US3
Iupx0sz9AjuINmYRFg5tfzrdMgLpTJ/r9SSTHNnMk8RpOK+jDRX0Qncm1mmK
Abp5xWHpt9CZYKjyma/GakU8ywr0IZckeJoPVJYZiOUhEIDtQSTuW4x5cZGk
E9ldcMu+NTsXgnoMpZSn4v+Qi22TJsqixL9wRPy2nG5re/NPCLpXs4t+KE99
SIAQFcu7f2tA2IEHC8HFLBPd67YVXec3ilEiGGNcsEL+ncHBiSO+RY25nnOS
jrSlDxqAkuRt2Lof0P41JaR4tzwnGsjqKb17q+tMrPJGxKTRkiGM9WWN6Q8a
7+FIpgNEW5jlUuWjtd50BQ8IjkJMV2SQyIR34QkEm2V2ANqI/ujUxBX9MDbi
c6lTSgL9PZ7kjpyW/iasoR8M6eP2UBmFeFT4c+5VKkNjlReHa64NP7a+5VkW
YK2cfYaUUcM5d+SO8lJ7FOqxGVcMvtgm7k8I0pZywIeONyt9v7+yy+I3cWU6
fyHlVK/da9EwflrNLUnRt2yzkeAaIvDxWwHTxYyo4krPzepJNrFsdihcX1cY
NGuguBAmJYTCbu28N8Bls9AYOvB8W8BJrmVdwWcF/ZnZfEodGH/gwFExZDp3
DmHew4LiZczWTovdKyfLA+tUPaF4NgCLbQQscmPfwHkzEASgYSTh37dQQ5w2
zh2bTyrvkAa/Fles4ig+16rmWYWm2s6twx+FjHWnTp7hUc6jfz8FcjUrmY0u
FMSGP862XDsWliNgHJFmkJaB5RzwxZrhR08lIsmNj8YsRmA1TGbCc1H/5FDY
4Xj4CkIF8dUH19PIq7phnP+X4lcHXoFCz6V9XCFEZSkeaPRKvzjXYAOhTJZ9
EHnWHMbAcPhJlRAqoe30UzJsiOeRKp+Zfr48Wqhub50qQ34RltU8Gq1TCXa5
ElgA/ep8pvT9VX5Sfnn4+VlT8g4EtSqRerng2ve3ANgTeZtyYgcU6fP1REs3
eWn9AD+P38JQQHQbWpaa8vOgMt3LrmDwqmysjGs2cHpBTEFYlkNigqfv6HgF
XNwlDdutPqLhN9sz2eAUzmmrqiWBBW4znJ6B9FCpKT8qqc+BRtE5xILVhtTU
loEb0f/Dvrn9fYhaY04uDSLpCa5bmSxymJZ63Bp5gt+AUv8mYq/5GMDnPDpf
D0AhzTHRVcTlwMDw5Mx0CwBFgy2SYyfMLFrztg4hKlxNEwshP8KVRyKpi2GA
MtftLXcjFzErKjjERC4YA15EV9Ane8nERnn0Jfs6GW2IZyvC5oW0DRlCnmjt
qv4WPF3SmHEsX8tif2s1PkEEBKCJFzhXaW33SUo5npsjUCnBoL5WhI9UgsE/
uJGexOmwshKUkkaVRjAC+B7nf0lFFjU1V1S7G5EvcNL8cbBlwOEIQehVYqL2
AWu1+1Ndo8VHDIKlEbwKrXNYt+JTezPGh0voONg7Crs3d6rmHzidV80UpzKp
q/VUcb+juirm/g1QFpYTfUA3h1HwV0HJWZT2eHngoWuntqUkzHaCObe52WJE
92Xa8VRaeYhsPki30Izgl4tCPRDuMNTCMz9kKE40GqRnBv/+ohdspTGcbRi1
H11FndK+XA4yuVlQ2ZjzNSa4AuuPTb3JHk47JZj59Ms0zwIETRIuDfKNYgye
xDOH133LOBOXFdN1/VOzlTY2iCphS1YbqyBEpscz18kQc2+Dy7m+x/xg/a74
n+0ubdCsXs88gYgO9BWR+9Rbo1dg2Y0WBOkzANthn46tZ43H2TTFXrBVQTQx
qpoaUTuP9fYdeuExeioPTuyyIANFma3fdHBlLO1f+igJbSh9mBihaWqbGnzu
XdgsOhNWbh6uNRRz4BDkmXVovcY8IUFeBjtcrGwoxpqXHhFryPX3tzlj/f/X
bP67cbv+5MdHmot+atrSrk4PbY2fxOPwqaqYttALHDmfg1vLoY/xzZo9EEKj
6X7lAiQ6m5Dm91zxvVFSIunkPa7imDDhC1qdhINnfW83vYYzO9efSt/gRZ/l
gNZPzlXxERQAaUwt9Qm+sFr8N8hAH18bfOLtvo58P57pkboQ7zarWUECR4s6
bR7hhWzCadvu+qE1Ey79etaHqxZk+wufwghjioN/B7bTxXZCz3Lz1Io+g3R0
EW4UIAjP5Hll48XJAqasv9Tm8PcuK0sbJKgU+xcI1/+kdPsH9Tmr7f6ZTFHq
6ogfZu76oYen0la+moGrRw7TMg6QyXjT9eyumxvkwEHULgUbNuwZ995WaiFu
f32tsUKY7I3sDRJQQr6f2elKbk6NyK53F3LhUbonfv7WibMEchK76racyEQ7
iWuCEPeTrGZheelVI7I2QsQtnUU7iOZoZ1lnCN6DEf51noZcUb5n/cbfEgZm
Jv6izE8fKxf8fevfLBKtjPuh/gmwmzuyugckXU1baec8B5vxTOINyZ4QrnK7
SvXpYfEf1UWH3BvX+aZ9S2ZtIWJS/RPboIfCLxoSQzxFUUURJH+uWAQQrIub
lzKZLM6wXC7dtXa/2de1lxe3berHakkQQf+6VFZ6uDQnOVdFxp6YxzOenGLu
yGD2PpOk3xF79QkUGvXtojS5nQdPM3+rFziTOFtSLh5rWrqmUa7+vvHEo4fY
vqSFc5SmPQBaipa0JeUhSqPw5pPKwx65KVfQMUNBWuNBPSGy3+S4TLpWkdkh
FkTjNL/BbGl2oWZFNSMWr9zpFU51HV5ATMdJKhz5EjypK0K+M/id7GXniZy5
o3EwEAXGGwwXgUk8EFnIXczk3mPINS5lh7cy6t5PUHjTaFsenRPd5pi9oUWy
b3im7Rqd3PScQrwUThp4J6Qfaaai6kCfh3i3qUIV7IOIxy6JAGrPXlCXCHRg
IlDDy61ihDtMmbg8213PoATN3aeVQo7XjuafuFYdzaDJmqz2AF89tlqioc5v
gqGOJgkEXulSqcTxaqN9gaBP2fjG2T25Ol69x6K9eC9pSntpcgRUyUKEJa7v
4izKIrNAXAi7vT61he+EN45XuMofNbHLyqq6HfH9aUniVsGTjx09ZVx9W3T0
NWpUYyG5PL9EIAk4t3uoTT4Ac8xRdEgCCvE8J/Uhcn3WcO8Krch0ZbZs9WSw
R90OanKsc/Ajr3CgafKnTck6/eooSoB0eGsiXj3YC+AYaBh4MAjj529qMNNa
azEsLwyvbxXOhIek+cxTFaULxpAKh1mqPSCfJIgDPA8AHXDeIU7VjhqN1bDc
OopGw3L/0ac4H1GG8qo3+6B5BN+dVaX2Pue07Dzr3h212DKXdp0J1AWYyUgD
4p+cVqu8uy0ww7bY4Vl+CjuSXgO2juq291mU1C7npQQoNLRNyqIYdV+3SI7l
lM+rFWNc5+6185ERhBH42fgTlPrLoAiJmmxyEqAOdPnrHf4z6LNvGugtLmmJ
0QjAlV/7CYTsxzzl3KYwzazAc3gR3jJcPeX+0iFqKOf5wzzicKVJoddLQ/tW
kaObksImOCpvZUKoKw9DTWvNVGeCOdVnaaWuKvkmS0rGDxpQKLG6AZ6xzA/N
hOl2IC/1F7FMoU0y6QiuHP48W50Dj0WoQJ8JIdBcZ9H8Cb44FlaB8/Sr9rSr
RGY8I1bnvvsrUmHitiPc4JCjV4mKRffyGX7Z6pobiHS+kTch30UK+Mz7/EHI
iPyBj9lYx5S28mzYK8OYRgN1bC4VCZsReyJVYFRLVsd9GKJ/Kv+w83DlQZqQ
tqh+BNTrlClDjlVToNTf7x2YaSs3wYgazNva5xoKC+SNUIyrQM5x1MEl2+yI
M18d069q82xjuHcReioZxiOlTUC3aiXGsmLhMbyuM3MNRMHs+pyPJ8E64m0s
tAfJJfK5A28I1UTC/8Hn+SvJLJmqJBAbqXq8Zs4apt93wfe1jvE2sp2OKr6r
I00KK0J/J4d9leRMkdsd8XTQ9EKbP8TpamoYBcXuZnNVizkpHfaZQndVs+so
6fjzJnAwhDprYq6eBxeZVU8ikMMEbSBomYYbJWyja1pRS3I3ZC7/Ydc4qvoV
8MNUtccnXDC4cs/VbWFqIcStwY4NFkBqi21DAa3g6ynC/jUFU3JPpgzvUzMZ
/R/Cvxg6H1i/5p3K/TtpSuvk5s8t2xw941bCPfeVAJHNEHfUx0eFBkaHVjan
cTau46QtbvK9/M7U5ViklTx4S8jcGInboqQt0Jq3NgMI3YUbCcJE0iHJ+/qP
XqnVzc+O/AH/2p4ZKyCXMLVcHKC2Ip+Mx0aUE1ZMP4w92u9eOihLxgJirTOh
HrwFU2IIKYXmPYrgxE4ixFzavyYiAH5sKxh1w0+nTy7FR3df5s+7mmNFDGjE
u5XpnCF83zJHUoQ1qWdV6pjqP+vF+nUFssKZp2QmA3/2a3QfOR6MpDVdoXtW
rdtzqi7wD67gJihJgTUyn6OMRmWkX+PU87Ft0POdbnx5PwBJE+AZ4tplOFKI
JuYLsbPiLIQpo6aBPIzvBFo01zRLCrhFodmrLU6OTz+Aerk4W0wM6dGu79Qo
zjYBeJMMhU+OHvBMl8hwB+RTgL5x6fhxzIYLA1FjJyxOo/lUNgF5cW7tTBm9
K3DoKtQT4T2CDdmzVU1tnS2N2+UJKcZQ35eHAP1/WwUiTFQXMQAbdGQ00dFC
csQ6AiAUQAKrksNmJ7jufuWkHoSAYT3lj7Eu8bMGK/IafE3mEP+xIJAkvn7I
GPBmIoeu27dmyznUTmfPIYqlK190mPPhyMzKARnetnBuBesjAG6UJwoxCbFK
njaylrh2WcmFP9xwCCdUaBdr4PtBNS8dpRmKYiupCrlnr01QRVbQUqO7q37I
h2JF3xDzfwpHd6W1m5QXsBIfRZ9nDvfnDb6JRjCfish81oMXlC0ROFR65Q0m
bPgxx6AlqzutRPiLqOCqF6hauvpPR37+4KFF1l/0mKSolmhb513yav3/8YQM
rvfqCP9wWiBYtGmxSx2tRh+AJZJZlSR+jBx936g+uLPtRYInoIg9O6rNLiK+
S3snk4bDA6e/QnV4P+jf4kIjn51/A0Bj/kUxzpyAUeYhzP4ryQ4hnGUUwp4Y
rEB8f3JoW/w9JzlHrJUd/y0FAOzdS+2J39qS0TA7jytaOiOFJIXNx/YWsXCE
fGbOGq2n73bZqsVDS1nyc4k/RuWVikxIFes8IJWYp8SIkPeUt6uAlu6FX0GK
3z4Qo84sC7UZOa95T4XCuYdOfSLs+Sah1FtBkqLhFq6b2n8+O+2j6PskBDM8
9jo6Fp2uL0kJKZ3qTWYBHXlwXATNqUIL7o7hx0HKsjfK3WpcL3S7ZekB5Pfa
T5odWmRVOj+k887ShrMuj3Wi/W12nFdzP8b4IqpbgcsvxwuC0yfP0qZtog62
vGqLIdNmMUsUBpuWzb/h/7W6GwVyBeU3WCV2YbyY0nmMxDh1/oXMYT3at1BX
QoBJqjK4gvTKCilFvUnBN9g14L+bFDItRH3ZQtV1qLEPM43wVM6Ehpbsk0rA
cVYSXlxCfbsFC5iTBMLv4qBHk9DDNk3fKghKWGyzthNVptQDL7CgyADCZbLd
Sy1VWl0Lhb1zQSIuVmBD/2hBdFpzX1yIVejVbldxV+sT5xzRjr6TnKFCYjej
+rL9jaRtYMaZAVcHNj+YArNiYFeWozjgU/kk3PWAJjAaWdtC94WTZ6+TExbd
2xkPjLt80jDjWvhJbTnZvjlUWBQls+84Dbd42fO/LGvkI/HyABd2A0fCxJgf
7F+dfEXQRlK+VP1LXcFGVvGvC0hH33kTF3J5kvlcOJ5A1B2HMMt5uPikdsJK
GloMy8Xh2A1Bf01Y9djpYrg0eMbW8I2lS4iWCGobUCGfQ7eaWdtNU6FMfeYN
tRDKsTdkTPjdK5sWxx/tev3JyiUtISF7RRUzRMajGFI9kBnbN6YTXMnxYw0R
XCXvzV90mFo0HYEaCCUiw0DwRZ8I7658aL8aO1r+naVf1R78tP6+5fkTm4p7
NtwYOpz7B76vp9wnxKd8/CDrRqbtRaXglGmv2G+CXPr0g+DGvMnLAfsfSCMT
Nq4ekZnshjkgCH/amNm7L+ZNh7HPhZ+61/kvHIfeAE+w9wuqOatZ5b4jFGGL
+b6zBcL5LJ+z0MKdj0N0sQ4p38aZaDTMggHufC9lQX2Z+JNhajkxnpNT3+UD
ZWZ3mED4EQa9U5rQ4/Ypq1A54uEhbtAsqlKUGbHf93J8HPuy+FXqqE/pERlW
uz2ewNueH68Kw0g1bNL+jThs/5J/picdtYUvynwdzWf5uzXd03jX2t17QsG+
seKU2WkRL+kRtvG696YJI9Xs8WUgXOnyDqr2zy0MSkYtn+7HR3wo5D2bvv6E
0FyNMHMLFFjNeL7A6rLd35Kt7ssi6f88ElF8axzFn3ITpo9PO9ARH9xpsbn8
93Bc6tVYgOX7xFR6WNQaL95yXqj0yZta9zUR1PZmOWHI6kCjGoj/UAOT3xZO
qVAPVEu6enaR82MKVbTam/Iix6s6dHnS8GswkzTZeDGhMuy36wMXAibiQy7L
4q233Cd8uAYv/BfzKleTwHLLYb+o2rRZoUxNRoNc3RgQ/3nq79Y8iSarjRHL
7Tn0g8eCowRFIukaLZqdGCQXRU2vcgL2DSvBpW5fDgpwU8t0sjOq+fyH9/M7
FY1Suo9+Vh7grozTU82RGW3BXH8pCExXLMi2GGQ7H2/vA7IWy6dmoqPCLC+m
xp7DpUlx8WkOVdJrEiNi5V48IothaweNR3YyH3HcETm0Rn6vNRZwNTVDhfR8
1WdiH9yInuEFgpRxWaf71FsxNuXs8wBp1WCdrrKQsQjboArUN2lQpTWMf2EQ
laPHCw7+a0C3H+64KxjC5PFO6M+hxbwF8RfOKnSb1VzeYK58rasFZsUtCbov
C9p0c+R5d/EiGTs5R1tHH7NWoKwkFgess2calUwE7CIpRI++bvFe+YvZ6L/O
2PMD7Y1YZs80AnuEsaNQl5OVpyaNaCReQV/xcdKHWzrNAIOJh9vL0Yka3gwh
grXLhChISk5UQk+Bg7oqeFnmIrvBIFgI0paTs21cIjWoHkIxwP96QlnoNERp
i42Q5g7J49RL6CwUEfGqr7xiE60bRjt5IXqyPuWgZ5SDmKzG6KSeFkK9pue2
aa8SojxqFOO+C6OyoRVswdl8bX6j98Hi0xwklOGvYs/0zKSdjPgfqL+dQ09v
/VyrGC1wrBaRdovbPq3VwnN8b/QfZbMTRsoPum9aLGm07fbaz65h8zK9aO5L
PxH0AcZp8NnWEvSidrnzr5g2/pm9y6dPOUFTDfOy6herxLLNmsOaPWufWVId
YIpe4gKqJL72ma0g+aPI4Srwu2DSSLkjLGO8kBTNp/wsi4iH7XGQrLQmyAF4
xLBLUqBapqRMbcdM06APCu1VU0MBA8NzB+gV4DituVR7R7LvBDQBeqhGbyWV
H1dO8R308UoWPKlkMoCvHhQ0v/pt04fZMEZJGEgx9zq+DhzEuw4OATtCiLJ+
aL4xr3uZNRqQAZYUGtVQCK8VoljNAmuw+Q80dbkH+tAaDKUyLro8mqsOvvfX
vRH824Y8XR2n2SugZjS+k+Tm0sTkZnqxMPI7+KVTGmf1IXlr9v4x31mNYZHV
fz0vmtGH8rB7IGrXOIAMM5KaKqzwiv3HIppa4E9o7vcEW2r5l+jAG5KRrGUb
5ffAWAxeMy+9rkZbPLhIEntKKlfUDENLRj8YOvqFBEpGR/57gwHYGHxF4Xee
OJJoJLmlooctizA5zErRHA3g3ifyrgqfH1xUBGNes7STGmamlFkoBkAcngos
YMovHI4PXIBXkX6Pd55YBlQJr5Iix0TnDvanwHxHdAWkWP38IvoIpeQ4036R
fX96WiH9SSFZqP48sY1UqAxfBb1tylzYkWmEq4Ig3jJR/Um4fCD9I9aXkCPj
o3YMGkIUSEd4JoqiA+V3i19QJpypD56LeKz+Ow7LB8g5RAUnQVojdeE+du0H
Y3u/wQYxMOSGWUtpfFQ5LyUlVBDwBkm+0tEQawrEqfBAeVSKnfTlNtzpwnhN
9n7X9uzeD8MUuvSbr1jp2E9I7SiMylzbv4++t1XbzFSlK1gxOTqY0MGKK2l/
8cgbF+82LLFr5G7o95A8gqILCOOU0hvqG2zsxCPAKt/51zqqhOoGWFiGyG5L
w3rVxljZW12fR16Q27pS34Nj46GHW1cXF5/lVknC6uDyAZfokdioZfQ2zyWw
Y1WPyYTKnF/w/jT6aQHKJGfIdAMAFs425qixIg+WCd2sWLv47zsI4uM4Da6w
DbC+ycs9eP6tPX2tq7C0QDiZCktybDL/61G4hZlbgjl7hNXbYHV+crWePPvT
cpmuVgO8dD7glGh2wif7awVi5DChUJpdWMGtGzxv2If6JKncscBOy4CZXmrW
hIfvi+WI9Q2s8zR5CfPD53VVYQNS2+H/Lb7hhLY38ueR2RPHXPeuPZ9XZCWI
g51ESx2dMpgrcU2rmG6lJ+Ed3OLOUh2ONCqn6gtXCyxH/qH50pJaL8Ya1uRD
rr+Y0Hg1K8Pv/4nK3ck2aLcJrIb0GWGKbozZokNGekaDRZIwsoq80N4XrkUJ
SSBhjZP2FVXWQhbsLemDkILEkCv3hY6/4PvqQCzN3fSHsj7uQLtQaqrACJY4
29XsfSQrz7vW7/86ndWlgCcVLemMp9HYpBs3ER4/Na9cGo86yxXG9GXG5OYl
wlND7qgeggzboB7O7w1zynigrHMm7tR2qpJHYwkoa/Ayu9P0RdhrjlLGsx97
R1IbYSxMY3MwyiRhiwXHz9mnhWjbxg+4y+0Mr0vaB8bnI8Anf17V4MVbyICU
xWGeb8XKw4NBSDCNSF7d27JaovzyEVUw5B+fhIdMpXvUg+GEEkXAfCg1Kiis
wWwLbXkNuMcHdatK5OhQMzWh7qKdyx71cu1Kcf7O8zHAYuwoQHvCqXpgk1a6
teEH0zfBQ2t94iBD7hDKflV6NXxXqUCb/lQ33JVYMSOqDgN4l0VbUCoQ4wgH
z7Ijb13aMS/DfyBmzDDhzV9DHWBl/p2vxgD3I9jowQH/oioH6USrIwwULnhR
wbfHcKyDCMPJJS3MU7YK+HGCvQ3BROJ/NbjSdRxQXRyoR6H22ECB4/dLUxl6
CKFz/xugwowg33tyTftyzt9nuaMEcE3aoQia3CBQH5+n9s++HsFSKZ5IZsZ7
KsMQBtD/QdCsjG8MRavZ1/7KVHQrP0d2Er9VvmxguH+C9KLTKeocHG+q7fVl
JA/zCaH1xIONyABLFKC/+C/moBn8u4SxD7yHYXyEgFmTl98FZZ7uIZsPkP4Q
EOWCuR23a07TVw1Cypb0VsqGfQaqfWq8+42ayrWcDujX6pmWvqgtgWJghFDY
MWWgpv+K10zY+WyzjTBQh3Q70nwtck4C+HDAG2ulFbGxXNPB4vsgsSWa6OmV
qqqNnSBW/mWSv+T5ceESrfsV6eVR8VO1pdcDorETCAPr0JfF/T4K5Z/KJmNY
540Cn5YmMXcnkaPMZNDX+FNukVcTIXEPU1FIZbh2AxN6gLeM8+vZT4gyPpZN
xRDWqaaEFrQuC/EWdVkZIghCqfXwb/r2ARPaHE70/6iTJSw2rAI/acsOuCYu
Ad96lUuBavbjskRMRkGbSsxMqrlyMKDVyfyukC889juJvuKIaYRY572N6aWJ
UN+Tqjt5S36yijHSeyGtdIdY6TOk6YXrHsFCmhM3q8qGUJTyhA15Juxv2e/6
yuVrQO9Q2nNkOHnAOju3Shxw8szec8oLyBoUYrMaUogeHUuvQ2PUYh5qVx6g
XhhhwGZ9W425UNjkCXd1lfOvduEVaHmzvQA+0GZSMbQuqS1mOZHWhDngioPq
Kno52E60kD8h1a+bv9YkD3kfuEghryZ5EET0SsR+ncTtYBLswtUzO4fmawqU
XQbJMkDkniOjjNwpwDAyDmSL4W7bp/VMj8cOE9Bqmxcxx3Mf2C5UyyT5wbN4
ESIs0HQYageAQvNc4r8pl0KGQzAH2n0+JcSD2K92775kpb4ptKMxbdwr+qSG
8zCaC4pMBJyhF+9Gsz3LhFIlUqf7gHnWkApgS+oDUkU47guvptBvfIUhrTl7
jVkp6foPsGa+SuovH+tZtnXNnDN75c+y1bGIkmcequFY2JfaH1ri9G+ypul6
akZgdtu/yZHS7rAlolWU9KNL0MsX6f9Ae7K3TiBbH+NH9wZYF4d4WZweFW1Y
H4vjAprON57j08rLYCH+3NHZRz/HDxPjdzB6v6k1AFFPeKSFFwp6KI6PTeUo
EOtpvRXofD/b/3hawgQryb7xmQO1P69hy9+nK9mXU/oVErU0goKGTT8IPQH7
VmdkgRED72vMR7Hb9jfI8VcCUc2wSP/z1SgDelizP432aSUpSm1GJYPkfwTr
wJOBEFBJKaOIJId6UvFldRd/e1FN7A7Aii2yxt7sxFW7gT9nSxMtPuxQZYPK
9P+sNEWsJBoXf7+RM2DCc2nTafIZLzB6rCmx5V+xa6nV8N8FVKQ9DEhPk8JG
m3EaTgtBo6nMEgrTKdubTBCwZF+IVyoz5IpTlwITOPkiFPZTKPS8QvQHg4XA
0jzGFCs5wYEQIkIsIFqYdV9tR3FtHQTfJSTYWqwLv3HNPZN2QvlGX9oZLShM
Zyg+gO5WxecvUsQEvXwClvBHGFWBjEElqb/xUIJmEDoilwvBdoIM4p+ASiC6
HExC3YPpbxr4fzVOXfS+dzfT9M8GcUuf0tw75g2AMwz7c9MdgvBz3VVLllW3
W7V7LKNq4GVZaX90ML1xhZt8+roK553Z9pBaFt9pqdmZftBqodv3fla3+/UB
VDhvn/Wl0E7nldjVJ9Uhsz7AF/dbejziXbImqgqIwvggXVqaCZNM/6biYu4z
QxCZ9Gv3PMyxh/9e6dzkQ3/N6hM730RB29psWECxBtQBzVpLAVhvHDzaYw4z
r6Uk/2066e2lljReWiOKlEIhhdVHoRflHYH92ZxLm4WMKaki94qj6D+43+mZ
3i/uEzuEXQIKPUben1vbagP7fc+1EzIzW9+GI2zloNUTGRt7rwEcWA3r7HlD
fjPMKngar2fXNPHzxfHbp1ahp/OHsGmBvp1ur8vJJ30CzcBm7EPmzRX+s9oM
QEeddSfMPZmFTEONyc/1FJwDcZjr2sZ786ZDAIuZKUJhwOlzoN6wAtThuKaR
hrc7Nb2ksQoGWTuchaHECfn6QocGs7D1+qE0VeMd4qrmy4tk/FZ0vJtk/U7D
5od9vkGa9fI8qHp2AvParTKDz4e3F8itATeTasfD6b/gm0GxpbYQRpBhctgP
sJ516XdN1a7kAIAs1Ca0rpk8IfmoLnnPgJqJAXB3kz7tYgGYBWBO9HFN8isZ
Kid2/OndTzzLx2j+otlmgyeCcNEg5uKfVviVjr33Q8f6pI6QnhO+ywTqzg+J
pBJCK38B/0ZzxWLAdqESuCeEF/Wiribp+7JFK6ZNQHPymwd7FbknXzDNYh+G
9IlJfZlg//Q7ZNpLK+jRNOs1ox/fXXxclUzuHsSeG5uS2a7fm/3CSV/nhP39
lKiaWUg1OjCHmta1gSHR862ahvPmZYpDuj90BAEHZYrcy0c0py6J3jExNdvy
j8mz6Elf6XxXHJ91DLkk+8GyjbEGFUmrg+WR9MBC/4YmdLzIe3Dt2nsdK1Tr
eQ9uKDMS9dL9+WJGST58PA9sWx5HaTXFL6xaokkNmGPttYcBXZESmCslyWJG
zRgzas3dlQKj1J7zOGKRCuSmOY2mtnJcl6CjcX88cQMsP2Mr0eMk9oDSbCUj
DpLwhPm2jLDAbMoTEsZPdatsOo14pSP9IyCJWuTdPZ/MvcQR9TaJFosdPWrJ
VDQbmrLp0fNVgFjoU3aHv0FyyRv01ajZSHI+wN3uz9huDaKtxggHFuLXHrsd
BaBHDDrFlXG4JiXcRa+Og1t6ZFafotoBnMOLJcYvnrF5qllm+8BxwnJd5Uc8
o2NbAfTrfJwR1kg2HMxikdPhSasj2Ck86vEaOPOLb+NQYNn03FgkLhGkDhJy
Y2pB/XC7dKBNWJnrRkXxJLBlap0V/MhbIchh4pFDHOuPUF++oewXwQTaXsZJ
Hf04YWI50/hU/ATIoVfOHG2cbvFRAAMinlalzUmk3H+wpPmzn/rGFse0MudJ
TTG+NSqbbdH3NxInI3NVt/3jJpkEZiW5jqbnsuZj8D6wlGiFFxQIt69eonb8
beQN0dpF/fQr0emfPpRkzLLMC9NOME8N04WxAKaWgysUjGQLMDZQetQXTIQb
gsfL6Y1hnn7uv+pdgtFXRuF/0tDibRDAfj8/o/rBtYdNCdCM2V90/1IswymJ
F60/Mpfq5fTouT5d1wHxlXgddjy0E3gO75LEPcw7kLztq6mnhX7CIT1WmPOl
Ca7qlSJ75jEr2gIlSj2mEEEXvximLY/AWegGsmp6csGXCPcTl7/6CaSFio0a
bpmI7S0GgckOfF7x09yepcE4E/+QtUdjt+XhB6JBVulaYrFHgJ3bq7ykMaWF
rdRHOHzSH3DZP7REvM8KUrEeH2QdxcY1hHvbsk0bXlalDqEaJbgma03ykL68
I9S/4UU4bVni/Cva7RFaC1zTnxOxmvZMoZ4WZ+scmU+vGHkzk5q/mCwr8ON6
I81bd9YVh1w9Lur59wuVFpcliNLKRtjB7+ciXVVMeT4Gd7WfgWS0Kf+yaKAw
uxDF0PhZIMHfQwcWzGZRLzRf0/Wbp8kfLdkJ7cFzUjMgGUCU9iw6F6gAlc0q
XyYmDbRjeVr/wcb1t26RjPmxTL1r2qyuWvskBYBgzYu3DaDFTLQUNVV/f/sp
YA9xpnK8sUwzWSei7GSg0kblK9tzqKyAxVS7ToZ+sS14xzucorL4k2ON9m8f
SwIKn4Qpc0J7Zr0VRZnaRxlRZh7ufEUQjDYW7ttP0U7gOtgTLIOAal5tPycW
DLNCbjtUB+X5m11XFX3pc2UrB74vcjk2LIUxTGHa8WQ2kzkeGYu3b8gFBHut
nDcCzG5fsSAx9EaCN4zbVTRMJNSGJVEEEGIU9s7HjFC4LWLeXAXdaQEkDWNM
0VO/RtgWmi7PwEDRNGW/rVEJVmNc0xIZt4LRyldlgXi9UyFIIzjEdq6Op5qU
3rnBZbysdPJzr4owIgD3Yt6h1awk+kRL1e9J4xaKfW4KNwJJx75MqwKTKCRc
glZ+1FVvzpYcnY8ibn8A7V5Ch+LTpjJQbqxeY05C/ugXrgk9boLzsfGDcpeC
pFqkp9nU3dkZpCK2JSCeHC8DzuCH/WLbPzCX35xYVSY34SXH5RH6iCpsuZZD
zMsJAaRk7apQbH/7Q36+0S5JURGO74yPjT6TdJtGTLK4rrJb0WaLUad9UFTm
fdt0b/TJx38HTEtqPy/rL8ExOHOg1udnkI76ehdbV2xMdZXmkPlJHdZUbrWP
QpH8dm5DEkq4Q1N94fC2k6e1M4gK2u7DY/ys0KZZuTUFFzBNiGvult+gyyJW
2NRAOce1swSPSJnvvahe/VqZkWjaEU9WLUAtuotmoTAWuchi6738zRTTt1gA
0kYQWdt4Lgj0FiAogoeBKdGX8mrWZujKCHuemCtRPQANEfyhF1UYBFueP/Tb
fonJiiFWTp4F6LS8X9fJyph+6wry/Hed91LfDOJ9zRkVmxEN3DRtC4n46ER7
J+Y/4YbPSdUvgcFKB6JpZjm8xjPN0X/ADcEwlcAfeIygGCAhS0gdeoxpgpsB
Sg9DnTtRqj0u/9D3J1i23fvW6KfJ3/bK3SXmcY8mVOLtECzpTCNC2T3JO4N3
kLTE0ymBdSH5rlb0cUgK7jOefvCt2jtUoPW8X+tWlBg6ympglH1xaTArOGt+
LRweY/VrMJtzi4+K6i1umSDXJNcN4kq3H9AHQ3mm1ZqUCk5WcO9VlvXcOtf1
0LjLSA6LctzBonEgCgeDt526t62mmA5SQfJ15qpfhM9jyf6hlxfeVNKyBIAS
iHP7z7ZdXG80QMW6hHcDQXPGQK7aJhhysmLqbqin7GBDcHrJYoRQCC24mNSx
4sC84JXjHZWmIQyZVddW+K7MdP8MekSwgxk5G6GZyb5Tl0iEXGgmq5wbR4uZ
+PiZuCWipxHv3YyOqG5zeAaqeChTdhhN/e5paDDbc2O03tpkxGxA3LjfBspN
rpeyjOIBmHbJWY1PWBfm8kgdsrGxM9ZFutEenKUJCBn0S25jW+cLPINhMZH0
L0nzjNId8Q2epYwmrEMHZOVOqnfKKZhXBsDk8dktvQ9e3rF6c+QBuUc5jF97
j3+JYxhxQ94v+iGjq5gVObNNDcxeHoQy0Mat60r32f9XLvPmWSKnI0aygmKW
sWF0MI/8yJFjq/O9P8C7AGx3gKc1ogS5qicu12AboUwOIJ5le3PJ+nh1whgY
Ag+UJ3aH8NI3JkyXJEFUW7sIqLn9qt8DuYY9ON1Mxo40TssLhjcT6fOmXIBR
aw/0/lonMV0z/l/C6NgjvOYmPmBKGfsrVtSvMDpZs+S8P1//gAV3sV5U3azg
4938FFqicWa8XMLymO7qygwMBDFQGX3Alc9sJU/OYBskeISxLXP6mOPvEr0y
09A9wK0qanw+x/L5cO6HoyeMBkMOfZByebiK9ae35CMBw+ITR2LctuSQzY5G
MeBfJTHo147rcEQ1gnVXpzdOgzoTtiJYqaUPhSDlrlMjsH9ILS8158cZYN2o
KImUbSlpH2b7eOmVD7+JdjolIknvQNaVALXuzr0xpfICQjnf0EIymg90gqrg
JBfMSRKW8BQXxcqwPnIJhyHzPUCcXrEx0EcpQH9DcKye5XImZosBNj94ynD+
2h7mrnu+RU3PVQnnKC/gaJQJYpyHKnkZw/9kjPsnUUVJa2TjVpkEqZQUjFQl
zQ49gkcxHQhyCnhBVvLH1zMTD1Apqh2gRr49BYadrOTwnksf8kaXYahD/AjR
F+tmOjx37QD8UwLd+ajvxEw+tZnvdQLn8Yex4H9NMpqg0xPtff1rgDKA/ugy
QY9LYAB3ovBa8kkE1fg5isYEQgIu65TWvwOUbL1KT2EEWzIXwtkWdviN5O4L
9zaL1iNgFBgMRyVfsLpEyBcSyC6/rsNrw6d4zCRhbzoy+NYGeKRP+UjLq7d/
Oh5Ph36LWB1LbJd5BwlHZnSD1gKJAcANrTboEa2KyV68aRdPBwMPIeL9IEQV
Qir5njvH2scsvafTF2xDZ03GWhc2OuaAZM3tC2aN7i0JiRQ1AkLv3sEjvk7z
IdAW8WSBfZrVpw+skmLEZALOhCI97ixvWjYTO7ecSBgtL8KcVvC4RdTvcHQY
kpc3Df2oWGkZ6bPl9OWOSjqrKI7s/5ekpV+JH3b6lvCYzxyBwHdzrCVrIgbE
dvROMOZMvSDxnWYeNNn/jdD84SR3Lwl9j5bwyqh1GVoWEf9UufXxZQL5zXwi
CL0eyrA6ghX78KiQSF3aywBcdgWpUatPd/ZuCtpVF8Cb3qqYTbZViqWrZraP
7PEbew6pHNbccL0HpX9sbdXl73Z+wbCBkGrR6+cGIRZ3X0QPy3D5t5wk08TC
TiD1hY8ufxkYf3UTkF7tnkNY6fcpR+NXeEmPv6yMXZbv23weXt27mKQvVpgF
M6okM3RHtJPHpfpCse81OtgImoVYJM+p2DZVUk/CXFnrRFEqspAvw3rfPotO
YiUUBW6+5ASjfbyps4NOjhdujjZdckyFfKlxuCntx20uZyaUYP3V1Ez4u6ep
mAPQHSc20R3/RvkCgJ5OFNBntD+nxvn879xJczFvufDQs8l4YOgfga+LzN2k
pDNrLdkvedUsp4qFFk9A59TGhSxgDPJSXR8mYdiIPIyDB1a9bTG3cqbuetxp
M8ZBgBlhFzA4sVpKKgCrBR/7bakqU4DrvxUUUHYLc554K+1fvL0zBhuQPkCn
Qap1QThGLoAtyMBMejrdJZv4LZhG1lySt9m9ctduP9Wy+sdZqrQv2Xxxflix
vLnex1D6xKc/Bdo7gmXLX1dveArX9MP5uS60PleZv7GqhJYIOzp224dsLcQi
z3SP0OkyuxaQEWA3oT2Cdl06GyIagTqwr6PRn3cF/oPnltyYymazfR2Lur/y
kQPXkYXNbe842NUCF0WhTzH/+qvGjGL8KHT7V7UrNIAv0hR37rxQGSBmqjPy
R5avgWoIGRn+oN7zshdhJSTs5kBDpeiAo4XUdU9QOjAyAa/cBuFJPp8Lcisp
DxOIB4VYC5OtNT6vd0GzaoJrXzWKlxvQDj3qSS2TDl9v4In8Lz9lkR6FuYBV
ZrGZgstDwRYeli4zSwhn64orZCMJB7QvTOkFodibAejNgIQtw3WFR6CIcegF
ce0SiQl0+5Djn9DINOvC0b6pZimvwV8tGn1S7ytFz8Wp4i1kguzdDTXSCAma
kJnro7LL9ahD5JEtE2iNiddzYn8DXZDKWVnaRiF9pyonxrFaCIVV3mkbyRcD
nVkb/4otOlyPPteVf341bD4Pde3MGf9GQoVUCo+nDrbwZcgB/BSfxcBHQmwU
ILOUHaRt/FimzWSDKPzdzw5w8V9viADv8aQj4hY/3iRQ2ILtEdIiVvUTVKnm
2NL1l3Fdysgaab6QWkbI2IerUauStPsJuvC01OgGV26fS7ul9/BzX26+WVop
ttfyCoFbTlwWhoxSiVePhcR4BPG/O30tJ+V0uUQSi5jWcMdOws3cx56Qw+5u
088xu7JKWWZi5BlyCbUWnysjCqA3bN9zBg/aXRZyRpcCgWPdomT/kQuwRkYz
9pXGyUf63z75ijeGoDVAGyJy1xZN4yTPIfUEmOvWi+RqcZz0pkYaG++ewRoD
A/YKGG7RNLQnj/4cVhwlyLGcZxXgo/yw4i+aKcdDjrLFrwxt9zjFvOcLcEd4
qXzkjH3s0oNW916JZzqvFUPuCYTUhkNNFc1Fdlbd4sRaI8BZBQpo2sB2Lh3D
xnvfgp773In6Z8zwSXmvjV0idzFiL4L8CmRmdnDWuWZaaI7GLmqRSbGYpiw7
Cc9ruNF1YlJfyZ9Z5qjbVOgyjn1U3MOc+jTXJab9V4xd1TcdWduQnpM/xGUe
HrCsiieYtDd+mw9JWXWR/IIyofn1AdxxNUxVGjlo2YsgHNJYAWR0w4WVso5p
jykFCVqC7VYbuYTitargPejMOs75JS6RzfxVUJvA2Z31nw1VZec5xdtRfux+
L+dyH/V7pYdjoy+f2DKGARi0jX4f9dwxn9IYYhu5RWKWlyV4QNlEH8H7O5vB
cysTlxBeBVKS5bcJLTqPVdpVQUObPO6Oy7czAMZdAKcKaxwGqlT1LDaqhCaP
r696iAMFQLfdkGvHz9dJ1RwIa4bf8T8Mdyb5G570EXLKQdaMbiXHww4XL3VO
J6GwH6piGF5tEkP2AW7ORGdnsrUepdL7p+e7kvcfBC2ImnJB+l/WUrfa+2wN
eY/GRpE3K3uvrP7jmMHKOKwW+NO2ElZUdPQT5xrLKQTq2LHbcnod0LRv/jXx
BxO00fKLY2XT+ofGHjRbRmz3Fc7B7a9HtIrDz4s6GVGcB2Nzkl5ZGeZeMwSL
oEtlYV2rnodqeP/BzqLx7le1OpfC1UXJLwLrTdsbvL+Uzj/dTtHFq+juic71
BhmZ/6DJuQQmrRf33dMvyvsTrgtXErl51RKWG8hhMPxDRe63qpYF3V6T4VEL
gwbo+8eHLonSkpH8gi0rTok17srwvECG3B7fkAYwYSELRFD2JtQKq+34nKat
5nWf8ljjjaGFw42NhcQbYTZJKKrgtJd6lm6MNmOq9pQx9dQnkOnpu41IuWu0
y0Gv+lS9cTz/uxdrza3TljoCNZ9Tx10vM0d4ohYxsFEhTafpq8oIF9MIrG7/
Ee/FUIszEdNHsEGxazr0IaSjtGXU2Dj7MtFx+C6xnPCOI+EW2pSp8CaPZ0vL
U9AKOM25YPkaFYc1F1rzLcldGXnv8gg1qW8y0f6weniKc7Has8YH+jVagwBE
qW4L0D1Sp+VkUAHgGd0OPhImPLAMbmIHfEOSBH3DQr3WgCgKiqGu4uQWFQ2k
O55WZ8DvEY6udMGdoPZhDFuHLRrkvQGWNU9WXkBtIVixXLDd8B5+mfgTSF6+
hZuN7uQ1wQxv0yR1wxm7dxIibocmB9keFPNnh9QWh7VubIRuffq2iRAIXfPh
E0KiYY9/0KNZSvGrmNYMVD0Co+gOsQBEBtgSJnEBv/QKiYfbKEGRvguhi+M3
jqDrZL7HndwAfrKhap5Q5DhsUScmS+v26rOPFMibn6gzMg5lSkr6kZij3VNi
LcTYWsHv4PKOgVlSn/Ipvj+/Vu8GE1vTJnkHRyfQfOtskDqmjoGDkQIh9dTD
wT6sl8JBqQac1VGD8suGTpftQV5ZHjcBr+xW+2nrh8zTBb2Kzs7/S1mtpsGj
VQY/MRv/AgfcIYeHIrK5do9XqLq3xX+A0qfcK4n4Cr+yBDvRj/2Rw/68+qiN
6XoQvnKDXsUo0LhiwWyLuJLgAIhgIZcYjeZmLKGVNvbhPMIhEkDdbn1fC/oo
wuwlhoF+d5LvFgoT17xPkrFP15oDNs3l0zUxHb6y6AwBL+p7YHwxcZYWQq6o
gUaIAOWpkWANb/x9tjlDWTf5MWVMM+X261hfDyJA5uoaFBLez7DcLb1cBzSJ
cjBIzj/cFswNw9efJc5ssuH7tp5wMp1jqtnl+qnkmRVAcPdw50jsZAulPLme
yD9NzeL2oC9IJ696y89eMw/W9vTP20Xe+0kcC2UTv+AMkEQjRpsiRmhCsUKJ
k/qYeDvGgvU7qPK0M6ku5Zm2pY5jhU6nq1At30C0q/ajfTUW7xvmJ3Ydre1L
UTCQiIit+u1Zr4qOrrH3SVSocfY2hitdrgcS2LFztJQT1/UHBEG64tziGzHi
OP/OIXFRCzycYd3RMZGYD7dtI7Jhq72EWC/lgvND/QM7v65mRQh2j27o64A5
JeSTQ9tAmXyIc12hOxRLuZk+BstAryciV240LjFw5rruY1C4Dq5OkyoywqSP
Y1yN7lPyWgHGccgmBkw2N/3F6xQ/01k6tDroy7cXjdg0vVkidUkmGe3mne0N
QosLaua0tu2XUxU6FU5mg1WQIgV2YdmZYan62iR05mGa9z5OYc5ld7tB+CTH
pSEVNv/a2qVeZDG+777VCMXdhkIdPIwSP6XQJyfsG8JBvrCB2yRk2TaMT/UC
CTs5mtObfk5D0bhGFbZwfV8j0w66laVjQ60uIlMqxVDuE/glPLSE7k/B2A/Z
FyjQhXwwdMm4IDMmjYJB2EbEt/z1hvcF7NRmRZuMjv1i2NvTai90CEg0hKi5
zGMd6Fy1to1VfpDmnkUhVnW2Z5MRMmi0Gy9OHYejP6grSz6DKLeChUjnZx/x
sr4GQFnGEQYq7jT7fkk4M0PApmPg17AccazYqg6GkqHw8yIUMb93mkg+T16Y
mRd0uqhe89IWw+14yJPv9ywK/Bs0L2Mf6eLZzaomq1rsMKhzthFpUxK8bIi8
iQOBYnIL1v4fxvj7oH/JMGYvxoTH1675DQrpaCEQD/waXr9vzuc05i/3qVfs
spEftK1FvaArrmvCLxFDNiRii58m8udRJKGdVdacvdmphnhdqy5d2T9czDGB
McIvhTTTb2+Mvp9A82vcixJdi7R75ND+OJMjn8JIARelq/oJE7rlE+EWXxMX
fHZnW7CCnmBQi5rXFt2zNxcuQs4Gtf+vCxUI104Yn6uwc9446vqstNQuSkho
3JKyl/XRhupahN7Tc0sOAnsc5gyPI5dYVE20L+nUPWi46dFq015EuWs//IJl
V7fZz+oM8XqTctJRoyKj9mW0skoWoh4cn64KsKpYVDALm0S1/x82FN81mYAR
ouWkE34xg5gzy16x2FYoIJrcl88Ru3/AJ4qzLVgvaF2Oq7OR5kctgZR90GFz
VJ+Zuo4v8vhdDcJRyVxP1YE8H17oJ8RDcMM2JGlcnLPp3QVyxEQa4+hvlJeG
uJmXs0MFKIDSNJWBZ8O0Ac+t6pF7KhwGPONX0uLSTLT2lvDUnbtRffikul13
FXzgXqoJr6fFm3+aP6RopVqMZY1Ap7JtYm/mqGWGKXumaBe7AA7w9Hq+f9Ru
WKVSnzjTVmkvQV0gj4Vp4AVEjmZG+/xsBTqJTcyHUpWyWPQ8kDbHZlOzTPAB
bZfjujdPE+1eIOViKJ7/JItQa4u8Twfvw4lrdztT3dG5Zf17cGtnBMlnp4ww
DIRlu/FGNcR7rNIgsPAXwTjYyuIGOUXPcHhQahTB3XL/kg4gTBl7YryQieO6
KeURI74UPhthtl0smbuStUkL7T2iZ6BHwI2d0y2NAWwjHLsWkyJMhwfz3xrM
PiUQ99us/JJMyOhzJoqUhLI4c70ajlVxuNK1HICmNTWdmIUIEPVf8EyanGUL
6y1E98vGLR8qfLkN3fCLwuvTKjuU1TQR41uFst2wy3CexmgZ6LTdUe+8WnCY
VtRdPcvgTIT4PN1MpT5ijzYK2vHcGO02l+d/zZAPHUPqRSgWa6UW/1twuZw2
ovX3y6flmFWFB2NX6uPNGNyhwxDuUHeIRcsGVtBrdiV0ANmhT3qKsW2bCihQ
V7ProMUox4se/LEgt1ArYVgxYDVXSu8S3p/MrzScpkdWb8J/GOlBO+2QpNU6
eCW3fsi1xBpSU55qK53TSLt66COlCAp8UliQot1faT25xR67JUK4uytw5vxa
6HUVToLr8RfqOCghxSFZJ2ib/HqwwvUos51v9MecXgsy1SXl94jTxeHovGYa
1mFh11f2+n7i7Ert9OoCGPkVj2ZZoCsg5avbVoIw2nN5IU9T0QuszPCoEsDp
Xzj1IBmYMK2SKM0ICilhBmLd9dhGSR7qjI4Fe5BxFCiPJcInjDcV//Nn7iOX
ULW+/RcjxGElSpCxkLvmDcm8a48PeuIPRpDKjgIeQp/q3Zug+x4jmjZyEPew
TRbvCrrUdwD/4ERWLtmSJGQpdknU0tGw9Jolk+Je4uAXBq94MNKEnji5iSxu
POXqJT75/bwhczzWSCMreTlg0S3zkcdUvEbWMGIR49+F2e3y+yWaWl6DPUi+
WqDXLmHR/f2OP8qbsCw/7h7sBqyXWthJvf915hyCSjE1E+MMRNfN4peoa4Of
c5uUFXN0Bgo3MUtjy/H/6w7FaS/F+v85ZyJBC5pSSmLuvQOVl+/H3nPJrCHE
CbrWKk4rBM4oM5PSMg17BXttu+ZQMkg6cr5a0dnGFoePkmG1i8I4vmTa5HzV
zs0j9bC7yqLU2/UGfgEB5yPkS9ToAh8FBTlutUeCbok5KSnfbXmntUtDfWTB
XrpT7MRiBsPBMSj844EuFFZFS9rzDO15wZlWZDeZBhM0UAA2lgSlmp3ao/pm
0kA6DgnU8iNjAhu/chKm/ipIoYXnmw4gOanbI3Ulbov+yzmn4O+CBnazz3Ol
6Ngazs3IdotAQ5YuSxpwTt1l0GpvDFzt35+Dci+aqyEzPyDYfb+jU4vGfCrF
CGp4WUl2vFaSJ8Sy/pBXj7D+VjRGVnJ/RV8hfCJn0eQUQa7gk0kEx8nol/RF
dp8x8yGJLzz8OpKCcU5m/aj0c/G9yhWvq5DthsABiNipYUDRcSF2Y/nBuUJ0
53UL2xQKxQExSw9NV80azM4fW3fFs3rTMFORN8rLZhCfJd/U5MQXIUTbE+Ol
mjXg5uzA3r48/SFCTpQYb8anMKxAfPOop/9BdYOqPONwK+tYVIo+9fnXWgyS
ZfIVTzvw+D2vGseTh2ffyULQvddOLMw38Rkb5MoQ73WSqlWngK91ueaTPuuW
0bAhfHwubAfiYp71/AAmTtyUtucwCvhgkuiT9qKoOO34I65SDAIhtIBM09v1
uZO6Fj1lNTCHqN/itdyRuXb+dMN42q2OSFKM1EDLpL23KzRGlIIEJ/lNhYoC
9ukJYpOw0USU4HNa3vlU0+g1uaZKl0ArfA0eifK7kG0Pmng60ltvHwu8H4Bn
6skzQDKpVB1q1UBJE6easC+z17uFsMYGbjpFtC4J7yqT95blkYp/0ylJA3gK
+ILcO18BxQ7+agX/xYjwJKtKREZXYvd7JLmGAkodrPNhNiVOxP4Ov7OIExsO
gVlWnSuzRl2sjykWVdwRYGweXEgvKxZeOcc0w/jsQG8n1efqbN1tP3E5d84/
sxRdT1O1Am1lISYKu19F5iZwFHRNoPLcye//PiwHQWwI/RMoDra+C+/76pCU
Cpe9G6mOY4AXpK1DQWWWiLg6HjdmFZVoMZo6nVZ6z0mVwEu2DKMVeclEYn2U
etIbA8MpwNjaef+xnH6EFnBx5u2GU4gdyAF4mZZz9EgsfUpYSft9Vw4aPyYL
u9jshqE+Xq1y2KJbK4MtVRSbjmmUM8CujWr5H47hDTcIDuaqf8wt3yKAJ/Lb
SdcW5ze0sSpApw5E4bA+ZQfzrhWq8DtQgV2JzxeLWkB3ET9obXCaZuKitQua
BZ9LP+yFLLVXPVZsuQzOuKOfZgfESNd+K0KzB/ky4l8NBb4+NyCbnh53DdNp
byC5uW0Y5A43ErCsJwN2GcVwCktkOzOTp9/lqXRDnIwqr25OFnI5MOJgW2jq
awH9MDPAs3b6Mjji+s6yvsxHyo3mk5IzfdSDwn2ISw0qkotU9d0WsPedqdF3
g+o4/1RrLgT7RHwo6ay91jhTGqpwzGzwZETz9Vqigj2BJll73hrS2YGHx29k
uo5bhTdHA24qWE4yt2FjognBuaqn2mFNCN2Y3UFBLanin/zVHZ9qevHK9nvK
vZE6OYhO0ajr9/vzBGe0JX/Ydt4RG+v3gPWn7QwPs3cwDxx2BWHCrz3Bcpsq
Km+kSnc6khAQ4yU+Nhxb5XUpOkdBZHvZebXSf2wVNaTpswOgEWQqivvBB4sw
4SIv88jgokI2u54OPi+3KsTOB2ufOXd+D3Cj0/WnSzIW5oWON1OF8KMoymoV
xKb+rAwrkYvWt0DyMoG0498RTJ+1n9aNTAIf84xuhhr16FJ2YWZxo5n7faCb
+BOmsv1fHSwHzhDC0fBRz0briu7r3NpRvgM1vy/lh3MJzG2hYYnpHovhTXMn
u6dVupule+jU/PrWytCuPqILcITaDVtLFYswPpCGYlI5AFCWWYNuLi9lhXeO
85FYg0fLmLowJho20XT9WO8N9vfFf4a29WROhuaIXwvg2t/72J1LtQo9sX5Q
GqEzJXD4wET3Ho1KbFXmPxKJtT8fWLXfvmeOrDPf5fKP33rVbP6ui7swR/H7
rsjO/s3zts+/s9zdjOU6oi2Wtd/CasBlLIqMhWYO3rgIR9cIJ4Jcu8kaztM7
QmPBoAj/r6J/fp6gNDnpYwYbAz2OzJzrsnGIqDzH790fV0H/NDkgckYF91iJ
yoCCGUgGGoQPPS2+B3mlL/YrVNZGbBvXDfhlGjHs2pbdjDlsGcpK/qt9H/3T
HgnlIcN5ayrv403Mk+wePdmRnVSoiabbpWK0/nqoqW9Zh+tiW1aZU4VVdW00
ro0Wsk7ni2x55vqOww+3lu34+uOmAZVRY06QIGnqGy8ns0+jXSZorpamSmVj
X7HMO8jlOCvME9qMqxernKmc92THK7rRBNttfPu0AbSje/wCEtbJNMfSGFeQ
Kqs5vXVjduuOndp0IA+CaL23Pnb8ISSTWdDP50J/nAxWJe5WsjX9UnGTGraX
NA7A2bPXGqD9Hlb7IT4YdYCZz0Xwvau3u15JqPVm5MO0YOyYYa9OFi8pNo6O
umDJvqQsd+mmBkbkqY8tpdJ0OUs=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzd8Cc31NFe3Q2KMSt+VOjtoln1vt/XQqnjpFxmVZqnRTwnIh6d/ZcB+qaFyogJ7UaLWi7GHCGEx3o5/T3dsJCIl7JXX1yxParsTCzxNj+28Fz6/m46nQYipcAQxutb2yMzuJcZXmqAQEaSsT5330BkmJQNhHd8BgvZt7B6tnR9erV3zHjlpKMXp8RbZw4NzFJ8bI6LVJ2wepFuFn9xTDH+RH1ntbtu/oP1GQ4ms3DGKPTvo4FaMYTnsODZXzEhM7LNLmzCxVW/fjteRnQqS9XtD9zL0u4tSuNwTneyO33bZ1WUz+6fKfqNcO/1iAOYNe45GTi8jRoybktYnj4MlKnzatU0XZWpyCdKLlKCzzh0V8IQkMiZZjSNMiwmruyjtrLmSXCYJ6F3rIe3YjcTL5C1OHJhdZGPYeWu+KOa2/VJ8Mtu1khS1PHuac7qgsTfFXua5mroHLSTzeBH/xVVlHU/BkSfR/QOrk828gcDxhOVmNX1Ya1fuhsomX2+vJVWytFxBMDlwt8bV3Cxsr7PgUumVyNhVkvt7u6p2vQavOFeE756TSMD6Q6WWllTjLHJy6r33bvqC0Y656jvubz2YUERdasckiB/QjyopFjMuBcLl54DRtKkRgVsnFmJyZ7m41Ol/5C1NRJp2jPhaVJxnEYMuANI3kn+jM/AmC47dJLdMNL4arHaqlB7g98Gde2LVlED09slDhVQGRCCRKvTiiIx+WinKSKivDUuJ/p0TXgqNfIfU5SIxX6EARZiATp86TTc1m8uYr4SSnzkerOfmazkn"
`endif