// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xjeXnTNjBNSO75b9EtuG66e6vdtDrGR6tmRPJbQWvpsKcV+FJHrwfrpeAfqq
wbZsh1zDRmMZSs2K0POawdFk2qjfhPa1fNwNfGtBqY6tfIkAaKXmxF5tpE80
cT1X2RFwmYzpvj5dCK4zN+79CLhZ+QINY0cwqIVmSErr73ekxyrZqKFb0rMp
ZMnxY0CEBrwhMKmtVHuVjwmgm7cvw/bfQJCFGn/4H9XcVfmZZy5iy+5O9Ve8
OHkYP8yFnt1J+MWijck3nlRS6qz4FBJ+Dflf+qgV/9AVEXUZuQ4WCYihKq9w
q7qiYzBX2UT0P5y3HAPPgpjPzMLWWDiosOSbePE3Tw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ml/LR/6KO5VR24ie71sk2LIl1r3qA02Jg4voZ4rEZfiMez2hlR39/skDiQgd
7jXAMDIzjCmqkj7yYYm9w+3QZ5jst9EOsCnfKNLb7N89k6urNpUFksI+1rWZ
1joUrrJ+Qh0wBe7pJlvJcPMW6QB2d2gA72/r0CJaJWPaVjctelc0aRAQ2n2H
ro3A6vtyXfCoKnt2Jhjbf0T8IeU2fmYVSUMXMNLe1dgpeElsWqlR0vw8M4rL
mu9EqBjsFtnPdCuWbJpgbszuA4oCha8bjGgZG4WpKmwg6tYFllA2Ar9RgXJ/
Bcd+pBt1CuebXjgRJW1di2PsmBURFlTq9J+gsjvbrQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WRguBCqKub/g4CZad3rYkusGk8Sjx/VvE7UbBbwy0rRQRwubMrRzgLygx+0o
Yc2xniVenIdmaskbvTw5ir0/+U0YwRY4k6oR+nE3qsPwditDTL8qrcFfSI/C
ZJwFbKLObcFB+hX/x0JqdcTdM698m4b1kOjbO2prDDE0oMZBD7nQHZpkKQVv
ym3oCqVz1WCb/gmMLjMHgrndLBV7HLqGYZMtam0qTSl67e2N3aSzXWr4z/EQ
9Y2lwCRdikMNvQscR0uBzLfeblDjyOI9TCHjYw9QbUFN/SjElM356d9zTnHh
j8ydv8P+1X1wCRJ6GGjHcUQB9K1UGyyykQxuE76JvQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I302U0pCX/1puVTGo1/FnjOXH5zpCNrPj6kC0NGY0SVjewI1YvThCmEpkydF
i/EIVGADbjvr/UZnzUKTB70C8vTjptxPbqe7yGr1y3IwT7PVmfYW30Hhhb2h
3NrvXrAyWe/cfTa+fXfCCtDO94oXIw7xWFUiDxbGgLfmSRBBZHZTX9N8p2yV
DU+DDJs8oOWRtiFSVrb+r8SHggJ9eeJuEUDcM//OkrotNwacYcZe24802QD2
NTkslBhh34/56xXIXeEE6oMF81Tr7P8fsUSa+jCspWKETlQHCz27tA9L5+XZ
k8A0LV5fnKJdE7TJ/DQNcd/Xkn629OELdTPj6zygWg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YBMI2Titbm/aaQ7wN2gDlYvULF407dMLDDj47wztZTOQy41h24f5OylshdeZ
wyJ301vLATLhqpU9+qmptnVXsggLBnolQaSOklwnvF7jmTCGqUEROaBzQXgv
vM3kEfGokVHiUO52nG4UK82YMArytQje2EjGbmci14+PBd4VcWg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wdVTXUm7Qj/cchF7KL3Kz6aF9Y3qXCjfoWGgaIfZEYEseoCPu3zo8U79Aip5
0fKRPirGI2OYYkOJkY95vOZK9k7cxzENRahUOp5NjywvbHAwyr59irEhBPQq
ppfjm2JcDC5uN9UiOAVq22EY6fPHnV+z6akP3qKBCa6OTSRw3yZaAwLCHHjy
2xfi9nMtvS+GQM2M3eJNiM1Ec/R9eRTKGz+LHNoQHMDQj8zbTubYMt52I8Di
NSGjoKgvrP4h1dJRtKSzp3qnmIFC0ZWrnV6Ss5Q8EssE/fbZ5KZBAtpoSkhf
6tu1IbgrYn9m7VhCyCkUblMV4M3ojf3EUkegvrN0JbXcr1H18LmNt5P6W00V
vbzamDDPOt7Lt3OGkUMGnLKAb49PE2QmaNwC7VHoUGdV1XYIl49fGmxCX433
hW3z5kuGyWf3SEPCku1HG6tdytxWcSRTkoaqsuTc0fhQwP//F9P3VZkut/hT
agjeTNVWThJ0J+NKS6XvpuLtnATS2pd7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VcPCH9MhnbUFxxnMc1OpmaYNqwnbuRG88TUTxyiuiPbmztY0DKsA3mRbtQVB
rXA0FUvGdxSAU+Lhk1RxjCsKGHLmbCzsxfA4Dwm+zPpDAuUzQXIX3xcu9v8D
YfTKi+Hk71yOVncBJ8hcSrUFUTZM8tEA2TuaHj3dECagGOJrk88=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dxqn3HHBpcoADhQmbreUBEKZ6x97JK7XSxLQatr+ZpuuB4iNNO0+78sOuWld
FUnHzTVQ4RULrcXZyafieIe3svi24qKbr1gapE3Q6cAzfzez+ZwG5D/z218F
tCMiFAIHkALxa6ZVlxgKObjJEdzBNu4HfT6POXzt/5C77rVOg1Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1520)
`pragma protect data_block
PB/8DxnPZ2Jtw6YIM5KjbcddYS4ikXltP3RJ6ZNT8cxCvjQuXyCdNAGmwAFB
8CgQ5RzY6zvC8HfqcpbIq54pkNTj0Wnuy64DAwdLCYsBIf8mkF6Iy8db/v5K
oJvJBGOm2YklcPuFV2/SkkYE6Cjf3pZelbuesiQwebGi10jJ4cn7STvBHdDp
Yxw3uq3rWWmF4ru5gulqSA9wKBlAwW4uIFcTlqojL9O2gzXt4plw7hnTZ1tQ
ytmTolD9VWKLXXz6ZqaxwyBUjgex7Dbq78IHkGyw5/3xC+KPq3j3LAPd0RmN
BL11EPft44W3QpQgByyuJXhEqKM22aqdJ6UGMiNUTBSq9qAmF2bJICXpVLIx
z7Ka93IFjJjEfFyPD+H2mY+3b7lHUboaryeZcKy5oplkGhzajV61pgYCQ3Dv
JVF1tIS2IJ0WOWJRZKfvPzX4JZke09uDUNc+14w+Z0enihiXzACE7LIjRP7K
b6rPaR7SxIOYEZ1+81FdiAeCIm9tlEUS15yRGas0f3Ptlx2brtvARVE/iiRy
AdQmszUp4CV3l0BI+qhrjUNTpKURU672nJxSZm3O3cQYykk6BkUg2iN2lU+K
jKxYy/PSRCT09DW8/1NtHAwDq3/SAItp2+AN56UA/PlIawQYOAUcs0+RCATx
dswr0xaviAO1jM0eIg3oSjDI9FUZwofSHJ4hQOrof5MnkUiJDLTfFTUWBUjb
2O7sx6UGlbmdYXq1HBK96V0Aqj38CKGLgYTrJLGZi1nQHrr2N57Xa8KwImRk
gmKDRN7LHyC9t+nL+4a6QIe5VWfPthtHk3dEv2ASrdZakgdl7pX2lionF1TN
R3CuoD/A6wMEZXRA1oTa8K/vw5OmOGR72HNSdAqr5SlqF7EOSp3gW396ZiDY
INt9TCGD7VhATlD2QLiSgToYY8iSLjF1+h+OUBtC3LEO+dBNfRHamLBmvvpc
kow4o/lyVbPJjgA+hltnpMvEBEyZeAeytEq0X8Rp48EiaomAJxkQ5UkQx9gW
dv2btYEvKv1AOgNU7TGck9ex/OKYSpJ/fDlLfEn09dXfIPUdqFvOAzPxIGDd
YWMR2CjNZci3VymapfAzHXdPE4OKvnfF6ruyXqC/NPe2rUq8LbwhEdIdUYkd
5zHtJGDvcS6Lw1OtCU/eavwwy7V/otgR8i5d54F8dT784hlVB49/apOSfxun
J1znkzLhHCg7hcBTArosrkTv02DfHg8ZHXxaPPZVtgJUW9nFF8eFwfbtrqpy
7oCg7ejLv4i1H+zkorbK4WVDVNtUGk6g2R0gfdYXyXAu3UdLSshFd8a1LPiS
YSaJa+miDPv7GVEMRQLUvwg+rG3IZdK1qXIh1zYO4/VzVwbVPjDEeT3sEsbg
V6a32+f5mzuSVg13snQv1wkGEr7MomQ5bVKh5NxrguMbwd4oTNO90oyg1/pj
ZYpmUYH+eNEFeGTOuF3f/OD0+0ESeKQ4KJQJjFH1FOj2I0jGBHmzk+lPVC/k
C02q8cwTbY1igBRbRLpkoWXC2Z69y/XDKsMX3Wmq010SHEcaEP6YqGlQlv91
UZC+tipHBZyuW0nxOWFi9THPCKVR2tirEN/Z5pJz9P4Utgy/4wA04kbGmS7S
KS1OlgLbnfdOyWZWIcJnYu43Gbox9J5CCrywyEAlabjT0kriSXatqeTRiVMd
PRbkRcBFQ6mpSJgPFJL3A11bezVAE8rF5iLlOBRKTL4RzUszxx25rykOYNYF
7VSZ26IpkP5oY6D01h7lvbxj+xVftAXgRLurSG63nNZubg5A8+NiB10yvm/T
Zl/Q86CAYUnPUL7rH0Dph8RNqhiL7LOec+eNyiyPKDsum13CmycqhH22qoUl
0Gka6SH4/LmE1Z3uUxEUnTQGb2O+rGSDJp1TijKqrYLO5KNlGIzd7dNjd908
OGnMpNAwJQEkyGya/xN1Mq8HsE0JmhZAFnkAvGuttdQbtui8Q94bpxoFy9et
vSVQFVBg36+D2haMfqC1hhahSfC2QZ/hGJrJJcBrt6WB38Y=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyLfAABc7w60o8fpl+oRYVrSKOjyrisN33nnvmyBFqEZzRT94X1KbtJxtcQiC9CU29AFpUE1mDEf0YWDuSiS3DQThASNBC+/Jw7wb4LoEiGLG/IREvJk+bisGNKX3UIOzyjMVEXis6nbmZGLNGLffkXzxPAI882sqdB19Jr1hyI2ngphWB5rWzGqziFVOtfkbr18GEB1aMT25GZHa36wrSkWrJ2nL8/y7N6/HuKe/4MzcrOkJcy7MxGveFzwevrOH0CrYN5Ai3dTAyQ1T1xnG2yO7d7IsY7jtUbrTRZ11dCDrBzmjnz/Y62qRAK2KQDEJa2tRm19JVoHRE2CCnw/rHkqxdOk91rKvwv//Zz/L9UnhP7cJkwEe++UKMrcr9cIo/LUFcOeCgEPxZ8o7WpZqZSaN/ouYHiUOgj2nNgVRTaPe9DprZEKnrPTKTKrcWmn0lkz8bOgjbdLUoDmZetWtn7cSkpA164yPOE7W6bMUbuvSa/AV2Vwc8TrAvzSCk6jX1RrTFEnmxFxxFjmgxOoGtlUa91j8JYwr0jXnfmBkY7OLpl2nF/ahaU/QKHh1THEfwiCguiOGlj76LLOfTPTVuSm/hmrR11KLAUQKMBTPfWZWuLiYBa4b1auJ0+cUZ+FPUhnKL4TfjcJBRyEjaEgs+901NrpcOx8QTYvigRBiHPe03SxtHUegatKtzEjaBarob10gvPbX8U8hbwEQQ5PDx+hR3bpaJc1rskVlyTZt8eYkPscz0H9Z/RUTD5IZikJdBhQ2CoMrlg7JrCM5Xb/MqNK"
`endif