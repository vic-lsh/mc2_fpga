// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Aa7jCUdPeHcyb2hgj2GdIvmSBMyRm9ROTc18C+iGgizmGYsxKotQu/VuEYh/
/FKvvk9CcT4jddAgao01OSUxHGV4Q8fBCSSmupoXIzQG9fg9vtjy8RmVtFP9
OUtw6ocuYyjhCSWFhXq/NDTUBFmhQtNhiXYK34OKENv/vxx+IW9zhK/Dkupb
Gz6bS3KRDlqucQiCCo2+g/k2lhZCX+evCuVpGekjB6VVFKUBDpZAyIL5rI1D
Si5nJk9uOXwDFX+vXJV1C0myy7bCqihgkzoLtHX25CjHquQGXT+ipoGDsvLG
XNuYLYk8HWOm8x05nLEdyFAWycDOIALc0qkZ9sQTbQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gWEd67FWYxt3okEUxKMpTPxb8lBNehg3k3fT5nWtYZqRhAPFNWN6Xxzm/Gi7
ZM5Rtdpy0WqBSv4+YA7Bpii8DE3lvUhVOQ+JJJXbOwMwxluVAVZlQ8B2DnKC
ROMSqWfm61ToRB3e7vebxkLH2UIjvxVioyDaBZqgIJjRqzwnPUh1LE7Sjzf5
nKPoNMknPqh+XIUk2SfV7QUm5dAhZrmDwRFvgKcXR1uklruXk1gg5yVrBUEw
S8FfczSfCdybRiN03lhm5hrhdPzRdC5PmOq1B3LOwLhJWnDuD6COC8OvqGi1
IWqde1QNgPtTn1Gtsr1l7aeRR7Fn05lHoozR/kfP2Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cw676iUr/FYKqz3MX6dNPufzT89ej+YoN1wEuEOJNGfS/MJJUUvLaS5x2G1j
HAAQI+ZNEExwNi+z7J72leB5XKfJdhUj6AobNiCZ/laZZrdDbvB1ZiQzGVp0
5unIiwe1IbvcNzRgdr4Sy/ZY21QtYnHbKuUI+1DtJRTov7lAiuL7U5utKjWK
aLp8lNGg8GshK4Wj2CRCSSf6amkOivUrriZ8K5fVQ9cKeG5QW6lFyq8dZbLd
PAUe/GBlQwl5L1NcSz2zxa+5R+GYmD3WZ5UoUKHNSB/XKc2oJOQxnnrfPLi7
Oe/+vmIqX6GqX5gUyX9czSzZzVURr6BbwQtnZUhhGw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S3Da2XeyzsKAawlD/lzo8KX/llOYf/VO05TDkVb4HcR60+7JGJ1dVqR9EuGp
GJ8cXlg0AuBwR8Bolm3dHW7dYTL8SqpCm/fSNZ5aH4pVc1/wikxHv2NQs810
LE4mmAW6qODxT56eMHt8Frl+QWx02hSmciPYyPSVqg1J+YlNNw9YyWhA37ZE
WfK36SNbee4sCMEQv9jxjyeSvbkl6PK/EbZ85xnqYG+NCZLXQWtwIW9NU194
WtcG6pllg/YDnlDWDqu3iPHYLi3k8nyPr1ImilbVWZF16CfD5orbC8XJMPPO
YjNnz9HWa6aYtPx7b/y6Fn1fJwt1P1qlYB+4Hgp5dw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RdCIjcRmWSrEO2vFYe/eHKX/t2ts16CR+w+vAirNN6ranFxwum1GcBOSrzOK
pSHwJIZU1TOs2uU5xmEHySbdOzqyiAOX3duBldsoU8axynuwmyv7P4oipOj1
6YZAtnVePB1Ehjy800aiE/2Y46QbhIXIA12HQbgh6XAUhqioPyM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KhfBMivC/sv/53xdxDIGwtnsfGiT3PBWlOxC02T8jPHY/EzhEcWSCCnMtHwg
Y8lpeQv7hJ64LmYddlsWvyR8jep4T5Pzba0LZs6lYnArQyyA1+zVClwPWYfY
h6WXBvy5V6mrpCYI317Eo06kU/Ad1EuieO83quu00rDKkXIHQUPcab/WMNFA
AWB0qgLNAKwByzisUImz3lyDPFFYT9J2AKlqc4wl+pRwvD7zqzbaTbcGwzGP
h18XXKkXmkyxcsVWMyir38Ns2ZZYwflTSmAgfyhlVj1fDOg7QTTmLIB82E/U
HwjhjqqDk/lnDv49BA+r02fIgSyIBSiDgsKzZzNGBs/4aMohVAc77jlAAF12
7OpSYVwkx2URrXAs+7vNg8m/yC2JEsuIKRNMmWaGl6Ms75JeMvoEC8X1c0N3
8IglO8BowK54zjr3Z2AB8N87SCYeWEQ6jZ6OcYkejSAtQpclyjuwtqcgPiwZ
BRyMSlp0FTKyWygcclsi6avGYdEHFgCL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DiNNX89RDINMoWNicwQ+qfKf2zLuuvcKFHPWZpWvCB5SfaOIIGbrYQEvjG4+
K7r/ozvKRJ2Jk6qMpUp+gQ6xDolt0YXuOEwhHch4raqdqTE7zq1J8EbgqHVk
9k/sKTxZPZG7ZUUAg8WpotEIfDLJ2F6ryGVpn0QIZsRrH0oMGh0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XSsf2UUb4t1hxUjt6EEz/LqrLAPdJLMoamJVSiePKkwd7ZumkYxuDtWe2o78
T+3Xjn4YfAiwwOVRIVZckbkoea+CrkDqIYXOO6idZzbzOR+ScDxE/GbzcDdI
Gr9QQBLSkBiQOAdot4+GEKqR+M4CHu+HPpQx+M4kiasLnqa4Fy8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 992)
`pragma protect data_block
VmdUA7U45DvEEje3CWN48EzOBSFgJ9Bq6idsujOYa0uksmPf3h3dqXW/WQfI
CveoX67cQ9qjgbhxlxRuzBskDixJt43T8JqhLJP6Qpxhkze2r98mng1JVINS
FgWtgHoZ/+mQ7IU3x0ZUkX6TBrVQM2m5yR4v7v8JlkBVXcguv6uef4EKc/Zy
ltCAq9ph0nfpEO82eluflLOe6G5+C4Clw4+vt7FL2RncNXgI67+fPG+PEK6h
s0UKv4JoNNiUjFKZpiR2rgQeymZWLSt2g/wdRApGxmmh6IHAMJwh1UNE5toJ
XZNAPoOGVJGMk3ZPG4A+edP72RcXgohnUIRMaQmC+dmHLCm88qGYMSqznHro
HSuta1qPz2fJxr57CWXW1Jzma0IeSCBV93/UcRT9v/E68Qir0vCAOgmhH8dr
FliVXunId+wQWHOEJ7b6eltdduNkT0njLWPd2ZxvC9KJinkUhMGE1QcSmS2F
S/cD2W8aqPNTr9ypA8xv3/FyTZQtQtvGhZdCz7t5BkqywkMO3ifee0jJX2bY
6qe/lQIN0mvGjEZTlGT3resJy77+BoXsgSSIEFhLZGRUmj707IklBCa4IjM/
4ccLWLGXWE/GDdI+qJYqjP5voT8rTrBZr4VHV/Vt/OfgYCzS5wyoKU831ZtU
nWnreQn/PhhXT0m8s4IFeYPgfhto68k5tjBYfUI8pveVKj0XaHlRMquHsAu3
qVRs+J//jAZy3Fj5bMq+HtR/sm/wTNun7pnqEJRpPfZQFCZGv0/HQoMfPqXH
EOcqtpM3Plqbv0zNPRl8V+uvxx4smWGqwBTj7aPMBW3xqVaDLCL1e496Jpy+
T9DphXwPh1HUSBz1NaqzrfMcZU4Xi0gL2bE10q2EZZUY/vOh+IJ5uN/6ORAD
NKyO5LQZTC6UgcLnoXrSSVrRnFcfa37LCD3xzKZwnhdqlMlGe4UOhIwAh+XM
tusw0gOCZA/KmDuprgI7Uu8Lzhgw5d2Nrdw2DDGK0hvaWb1ssnEW+JtxKpVL
+/zbG74Qx7OWwpqkhpHGDyhN8aGNnGBPHKmUnRnB/q/tHpoDbYtxLVEj/LIv
CVqfRDL8Obhr5FHMDJG+I+4ge/mfY/Yu31LlzfHqmlC41bkKFkAcc0+2o98P
5DXORuEBs7QKs1zkW97xQKPXRuCC6Isdw81ptukjqorUq66mt4QGlh/dpHhT
H46Up1I9z2OlNIqrM70wfRGAdlwoyfOJPY4rkg0/AgQT4zE9i4/0u5CP/Orm
Dl+pBWMUucbGRDFnMK8fyDICewPe8GovJecDr+D8sKzabmuylebZOIVcd/2g
1Kc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeZKgfROJigAR9FWat+EUUe8MONatM+NmoTJ/A8d2KANmb00DehBWAHUHqiDQvrimLou+meg/A4iqbJUOZ+ks718/eiIcyD9vBK89/2mUvklS2hSVYztcfUCe9HFx3iMAvbxmZpNzrscchqn2l8TMGGq0mdewog2uMiW+HA/EIGSo7HhWDWITnJN51TpAn15m2G7YIRmFYlmY0V0GkoxP4tLbncsaYNH7DzPOvRS3jxOC00tGBrLxiZk8lMDO1keXZVhjntwQVBQEogsXzvvBkakeUZlAXAZEzRYjj/YwG+6lM3/xF8GA8EVEwR2Yxc+gT5ZsmL4JS1rDeECMkAgpAlu+wKd0uaUMdYULt3j2ejhXj0Kooi9N628x0Zcc+jd3lkCk4fNpAXgHO0TYSS3HjbaZyUi1JmKcQQL+zu+vGdsnqWyMedTzVT8CvYG7Xv6XO7Wu7Rz6kDRBIBvrrZg3MVWOKdzM4Ucnt9N2As2F//p8msyHYo5N8fvrQdnZNesvVj3TK2gHpzqSnDaAib6M/9vTkoMhGvK0JVEbJ9StLVkM8YIHZtj7auA/CDga31TXhWMQdPDgT2L5hTdVpGr9aVjIL+8qJP/OaSZ+1M5FTKqtpX8yk5SiWUIQOOKWdoG+qeQdnRWqroO9WG6iaWq8cIz8a7TCKs3GG3QdoNaKenTnXvLPoldp02UHUgb4kEZiNjGWgNjJlltwOxQhBluBeQY00b5VVvaLSI8+Y/KaqjvzRGbaUoAFscw6KTOQst6DasjDvLdV4lHd3DDXW9sPt/"
`endif