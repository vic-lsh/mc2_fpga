// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QGfDsosfTiB17ugNuO4L8z7VX9e84cxtI+UPMBXoz/Bm/W+bDlnutSt5pUs+
enD1IqYu+HHXL9mxHaKzjgylXnpK6E5MTS65ecbvAOBKmbILDUr9R0UWKOVD
89D6E1CJUrNJwKEKR19mkJ21xVazM24kSJX8RFmWht2Cl9UgLACI6w11g4zC
an1dNSNoGYVRFUT1Q2sv0MSLOhMJAuhP1qBttBgU89zCGMQbWAlwojD6vZwl
yWbTTtHxEhM2b6T7xhDVpYcQEfatah86jdCiOFMAWyhM3Uvj/IEP53CkW5Gh
32a0xay+h0iYieiLtoGiPv2AM+QZZu2xi9mkbuDKwg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LNtW2J3tvY5BwayH7YggmmchRv+jHlnvbDzUmKFwdZFe+iSXUZyN+KByLu34
eQNRXpgvUAW72weuXPSqrymnMnER/Ty1xringn1Ol8NzG2nIwlNZ5+D6Mxzf
yXliCAou/wqPEdgGrBhdacjUzc5ZKMY8rewoid7UF6N/Dl1WMZ79xXEICnhk
a0rKVKKnaQMVxUSpqySVanRrB8niDoE/pxQ0flo8eKBjXYGOafRgC1Y50JCq
B6GGz6u5l5O3gW8oKkYQcdVEoanJyiz5qZACE82MDZjKdBoo0llJOkz2zjTY
iAhiAHCgJPi7cF0N4UVIDPZ+rlpP34LzI/HEXFwzIg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tKSSWS5ZYQWvWcH3VwXc4R08Pg36lD6aRECAgI/kqIdl+L+OIo7HsveOY6l0
Cw+6cSYenJc59cUUxUTSvq0jy4J6mmxp2AKJjcZJ3EBJOwF09BOsgN+Wa8pa
3HfS9b4n5FyCrHC+cKcqW99SGL7yp0t69gGEfZJu7Cc+HmYPQIjMtanjnWZf
DKO42w81hxutfqaAM+KExL2K9amu6nXgGF0/o0CgxEO7TR1V0PnbnXKZi83j
FwnYOKYi2bQDk8/tRi4rf5paZVomwBlc6Ifxv/8Th6l+/++NwXKzIKBqyzdU
vQEbOcPEMMFauCOfNvTYY9y9GmwCfXrFxZNJhkF6Ng==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
esZATPKlHEQsJZSZBdDVfW8uVV7DttixADIMFZ6gTJuDYP/p5l6EESEGO3Q/
HXiFirXmXPt9MtVyMpi+AjR6m+4gAY2HetqAmBz+2Ud2T+oV+RIbQgVbDNun
cbIwsn0R82NhcfbKUqpLRVUAcVix+6Xbhwtn17+temkiBx4bkWKCHxSN5FkB
g766YmsPnCMxIp9SWry9AQR9MxHQaN2BLTFOhH7E0FYa9VNAHRQ8wUi3f61y
3/kQMygTJD/sH2bC63jn+jeIU707q/3kvEr+j1kAffCDaIYIQebfMKvPrkYs
wr0cCmxgoCuDCQDUmmezAdqWCKv3P3wJqa01erjWXw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Jp01HLq60naFnH0OZcMe6PB4lMC/xjuNlUYEJjadmDwYgt7rNQ3f0K1VTykB
3nLJNpfTEEgXrNFrYrW1Za2Dj52aoonf0FrJr8fcX5ilmwrQi2kMkBrCPHNP
U3+//aDnOtkgYnST+nejtLe+xPZGdsBOrIax+TBRkD5KA3Qf6/k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gj4LqOoVoBAO48usFmYgmI8R1Rj9O+JDNXh4pURUwHAfpyQ0f6FkBmvjaIYh
IP57eCC4g0NHz5OsI7qQkWPrH/HWDVACZls9p175qv8KdoQoc1tsfKwNQPgz
aV71Jq04ArUpdxlSuGgG0fknuzPhH5oUvplklE11ewzalBXCB7umeCZeY/LC
5cpUFPoj3KYRAaOXKmp9ixHjta+HaSsmSf5B653b0SBH6DpIuhXDBcMDlVpU
WgLTjPTPXBYALKiCAPmR0YPCw7Oxno/BuK7FH03LY680jtgRdbmLghyDSMXE
5NIBDDa1qW7ry/g570lvuiX55sG9pQwIHwKtyQ6PwroRRCgvWT3mXbSrcfrU
7Kk8IBhrGT2j68j6cvhdVnvVPuZ7CSAM28zdW8s9dNez7O3qxUt3YgRY0pVy
NKY5LJkOnVOcJvvHjm/fCLLaSN4j6juPm6m7MVWbfzKL7oAyu0I1UlrGlPXB
og5W0CMMGrr/44lNqErOFCzBjsmj4YdO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YZa2eiN2fmYOdbPtDer8B/2esLKybHSEOPV3oGYiPqC3T6fzrRqoCyoKu7e3
wBxoHU4UhGVBgQBqHp/PkSacf89yUjldMkYMt9Z/aBuZlL5cyaK/D1afDPO9
Wie5xlZlkVV8jiLh6iCOyVvr81lheZxqCdEYn7RoU/lRuj8GOHQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GAUhzkI9A8unadNKW4umEMh/3rhxvrd2PcoaBmjX1tCoJe/eKppsHImxbvr+
hGps+jqESkfoFI9pez7vyKymO5+xxDtzlxt67X3JehTrSlglKkF4TOQHtLWo
oa8LXfWM5P147NV9Cz80CeLbxnaVnTopoBaebtTVFP1o5dexmbM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 976)
`pragma protect data_block
v6SKDGT8Jotc9W+6HX1+aq0OYlEyID4HyBg4XKFENDfX2gaSU9jMVTbOkwym
M9dH4zk65L3qFV0TpK5J9qQNqRyNdfMdQx1/C6k5OA1HZ9FvohznKhklLo4x
cX/ip7aJNQA5IvI748weQEaprmNca8HAMdGpc2zTW06AjTISznr73L0+7IGl
ExEUCN3HvxrxnwTCG2V0VP+/+AGXURDGcW4SWS3lCWd3Aa8eUjDCoiisJWDf
9Uc+2OeYjrh66c12raHaThrCpYwQr7zogvsBV86DqHIadwSVNYfw+Zd1IjBg
QkYei3Y/j35/q8Rf8qFH04BhgDFiSU2jA8gBObqLRwuCJoJpOLyF6jzK3AHM
e6XfEnwdg8Mpts6cOYRH+zVcodisNOi054+MSyQUjULgf0nOUlgauMtrmfr1
D1I0G/ICKjyyGNjdXqO7XIqz5kc39s9yyxLvDAKwwx05x4AozNelmBGxVFUT
qb9Qf3n86aExT186wxlwflD71R0nyAISY7ZR6xWt6ot3a4Kj6EzZg2rpaft7
N8ZkiTbrUz6YElDCj5rnzXHM1ckIcavR3NqMCBfBcNg2frGOVqBXf+GsxifG
OPH89swkAJ9kRemN4D/b4sZ/CuMKX47+KHuci1f0uNrHKRLq/QQrtVrtc/9X
9nt8OR7ni2qZD5FbjLic96W1ANw4Cknue1iqEuxib2rHtRY5WB1roDq8PQ+/
CJgTYIbKYbY+RxGhLv9LnNZtFrLv5RHEH5iH6bnoaozu2xrBQOwCVqIOBD7W
7vMs+nGckFiYpjNKRfLV0Bop7W01s0EpJb8mv7/mmaS+m8a3IGUmnpr4pkPB
P1crVszXbK4uzy+7qFQcBD/iqjqfPl20NowzAKVoPAIno7bCkAAmZPD4sb8D
5yixlfrabo4Antm17NPpnkipiUASOsO6xBN0ojAax+f4R5yfcGY13oZh9J+7
UeQ0tKWVO54gWKros6g5WiR3XKdVt54HxC7rxr/sL2juloJgALFX2Mb19b2o
p6Xp6ma34ZDYGrfkUTslCORpRtmQPT9Oo7h7xxKDfnmWnSeQ6biPYR1sbu37
LmW9GdjuGGti5vYCVsNBfgIBPX1mHKyKGWqwz9oNEjdjYWm5Iw8KpJPxHnZa
7rXvA1MxR63zg1Su7FkUa9AWTmMZriQf4pJeBTOl3q8HBzRMn+m2bq5Qa9lN
bEX42HwaARoYg0ciFw1FD2GNdVCBJlT7fn6sTI87OytKx7/zqosRqQbvloq6
rxgmzbngjm/pzPRtfKlK4Ho/d2QiY2a5WTKxD5ui6w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQowPTtK6eYzho42sWK+kkVzDRVO8983JByN1nK8qABiabXENt2Q834wcA3fqdrzLT8Xp9YPjOri08Z2FC8dLX2OPupTk3R3dcFPWQfEotamLdMRmzxExSMBQme6rNSB3J+YFIXkwITZuRvV0AYSin2mL7jGQ9oCJrC8DkCPyY1pr730sNGn/AWJWLXhDC7yTxHkXr6BRvU/mvUMDm5tCWUpa0Km8+iNyUNB2+qjmzPPQu1RIudo6mbC2UE8g5ilc5ta8CI4mQrNEfARmLN2EF7ISnyFDfElEK4lN6lkOmTUH/t9k4Cevsf5RS0GgqiB/at1C0dxFjGO6PjjFohvLMR4Up7VeZkS0RvdVvvl6E0CkyZiKhqEkk4SJSG2kHIGnz3AiB7Ju7W9TomBu851s9/EQWsK5BIwAp2f+StZbUwlK1B5DVUZy6TWyPQDPbaW2F96FfFI4AEDYu02MBeIKw1G6AlukosknAFQlHJmoD9jc/U01UQJvGX8TXrTXZoW/s41boVTZFDLPo8Yv3IZKZA4nyM1i50k9KeYMy3b7Mfswm63qgR3QtUivMYukpEXVv3BeoNgOB0pI5R7UqRf4M3uMcJZeFpwd9mJ6BFn1aFxOwvtY+hQtcx8AZaDg8wrv0HnEMrLs5cygyNe29zJ37dBLMLZmjhKAKzhulaKvnJ1QneQymZ0pjvtY2dvurTVN3FKRe3H7lrFBJBNrsnAQDtc/xFL5JC9ykVDAfeTsKTlZ9hHx1ekYz5F7+ffGcTWeJoMbRyOBbVBqKOEXZlAngiNA"
`endif