// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hZV7HWU7PBzJ06vyQxAAgg7KcMgHS2WuNbSEOQaXpD+tAxquOtvNpHagE5Eo
2P0DoNyzrcJefuDqJIPuaKDGpmY/54Xp2TSQHe9lENIQ33+p8wLZvNuHRawt
VG+kvSQbzOXQRax+NL6fqWMTYi4Cb/Exfv3eSs3iToBEAd4dQXs4PEYijI/6
XClKRHKqGKYCp4G5heVZlJMr9dSxZxO3ZhCYGzAi1SUD0lfHwmUnBy9BY/rS
b+6dM+Bw0Siq2afasJRkIhReLJaWHTH9jLRKZ8ZtpBjnNURx+iaru7LHVZF/
4A9bSeaVv/F4lKFs1N4QCJ5B4f3UEMVXIdB4ptC8Pw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P5rCdRa/dxtAIMd5BN8lx84iWRSQKmaUWJ352ovRdwPwnkqa9ogvH3hAmNNP
iyt888WwJ+eNFKDZv2Bfqbnd+31eg8zXHJowcnH173XdS7AYBfh9pq+flOK0
xRBdWn58EFGSiku98z6fsLHaWgYgeBrkFbYJKKIp3sFDhm1RAWxP0f2jH+8e
EusSJEHodjNDGj6KnItY/d8fc7VNwK5iTHup5Mpy8zXXmExk8+s4VjOMpId8
y5SiuMBn9m1Xp83WAbd9HqHmSkfRyzz3OhfDTIBmxsk9wSiFc+tYqNZBYASv
k63tBp7noSiQQhpkJ8XL5FhKafqoo+Yc1MmnKs/hwg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q0sj0KX8H6xgZZ3rikeJcN6nypUZBugEBnob3LMLUexe0U6wZ9uCpB2J9et1
EvFY+3APXgR41Dkg6iTY8Hzpn+lOuamoZ/A0b6QS3lPBmz3BWKqYQRKN8Hty
VqpjvwAfGRePFHBAmhZX+nq80UeGResIZtYMkmtFfj0j6J5YlmcYBQDBSHof
2HkKmBKm3OEdvh5WWH3kIi4yKWEATRFSiPAUrAqCn8vTpb+Q4zIEFNcMU1c1
ciWVDGFSQ2PTmXp9rFy8iuwDix2gnlfk0MbP0VLcdwIzbV9m7Aw8uc9uCLqw
GEBnvO9YxqiUPgN/5ud7l079xZMt/LWu0vI3a1RFzA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EjGRymZB+3tMu1VPsMsW89WMRFdfGDt2ssZJW5HA5p+7UIWQdH8zzcwqzIx/
tfNrw00OANQJS9phxtFDYFrxfaz43DuUAIieG+sQz+rZcIUifE0rqWvsnvho
URuvSFSaSzKrzTvPkuj7URZdNyNBFmuxuDDr4lvFRyqRApdYPrfMREqEsYUX
iOt/6uwmAbcZ1dlgNzKc3p9/r2NiQXDjdewlPkmpcsF3WFyhikFqlew/daqF
DuStXwIGPnpUN+pkxV39f6vIeJOALVqcaDh1S/o9BWwXMencD/9XU3V0E8mv
Si1lXSqFGYSS75inEySvB/Drmw2wl4oU0OuNzCgJAw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ixWnX+WijfaEfS0dqTX0/enGMQnERpZk4p1/XDjJ9tdWtzg3gVJ9qihbi4e2
B2oLOP+hM+YMgCfiRheDYn0wLwrbiklv1qBpjolyxzBJk2FXk01EFhzopQCV
7kztpJieW8qb8IAFm9/unqJWmIb7Gnb+imbWTI36mJFD9XHfFog=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
D5VvujtwtVLt3bRgDOu9wgwyodmzQ5TqZMg/+EoVRGlSSB5kByvhNJv7Nvpe
C6a/Hu/WEYqXBPEBIzEz1/lEAsP91CPIgZiZWmPjbtP/MNE250kzwG9OuqGW
y05R8/n+o1FwzsPpHXd/sgOSDQ205omQ+CQMqtNKUZ7AjOfICEXFcktSy93f
C1axq8Mx58VG/CvfyaYZOGbpuULiKm7j3jOn6HOz10uwUumRFKqbeemNKCQx
WqH2oD7E0pqbbX5oH2/7fHvxDgtpu6+GfUHC5/pgozzQ2T/i84ziRhZBzQ6i
0b6Gum5A5nUh5ub9UtJTZxuTh6Bdsjcvavy0By4+roIhJpRIoRDRU6cEjSho
brt7VFX4YY/jmR/z5adLMPJAvk9HMtgH/9ksqEfQB4oODVC4btvjf9W26uGr
9LXIOUaIKSxdG8eIKmZYUL2ThXIh73r040bRCwnH6KcYp53V0ujlwKYLU5ER
z98S/NzuO+zvDuOQ/6RM/2rJBjmE9Dja


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tDMO5387mDGy+8ZZUYkR0tuxwnqd+fIY1Jr6lnrWjYpRtFsZ2Ga6lmtJOl04
tdfKnrJRRf1+Oaqwdix6PTJkbPdbyXmf05crCsQ/HoL96f2dXK4WcLSDoa5V
/bWnTvPfCEWk7xA69Id4b8O94vM96FqtjOb14luExufraoHCXVw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KhaPwCA+KvU6YPPH+/pXgt0ihDcXVSe4FX6aFfEByhsZCYBcfNo0cGndO7pV
OiD+MLOZw/vPlB8So8FxTG0wg3ObCUWd9aacATw31FKmvBWY3mWqq+nxVuAC
ZF6CC0NyvGfHTHkKM+niYwOZcGFcxlU0MsTC6dRJcOCnGloBtqQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 25024)
`pragma protect data_block
B3ITr7AnfJUW9TFiUZfQhRn5QZZDZqPn7Oidxu4fdXOlPS2mi8ruLIp51TuZ
r1Vox5re/TM7+ynLgDJGXrdinfzRmdaBb3mx3cH3NlQ79HxGG0nDPqU8P0I0
bQ5VHsvY0xju6XfEZ6al5dKCEBXyXvQExjWWM/HHmcq39m+qofbLiME1KBrr
HiUtFMSBP3YbkXMit84f+Axeg20x2OHV5Rc+Kit/ajQ96eFARdScWDSEOG35
TW/IqYqTd0JjIBAIlI1CNVDmYNEIb8Mz4a3okryOmNB6D9MeV5sdXOtWQWsP
IVaYGuwU/M6Hcil0ulw9f7j+nqyZnnaKcm726Tx8NqpypwGe+aNMeeFBcqw/
8C7RWEKjYifekvdl6LHWVZ5wvPMn63kbJlf4bsedy4cROXjlig6lS/JITD88
HyD4q5qaol87m7NpcYTK2ruzZqFVai4m8APEfFKZcjFOgS71aDI81z/mPaAD
kTIRRyouTWJRCIkEjd0CIp3I+UzpGHA8wWWh1bvqYIDZ7EmFYEU/ETrFUkAX
p4hfy3P57LwOEBsI61jJRK9wFWjqJgf5wZ4IZWjNUm02ABG0itybtVVF9cvg
rjeBb+jaRMW1zeJ4g6WpBhFCPV2V1YXuGPifFEDGyb1NaLLZmtUB1E4tnen6
yNdk2uqvve+m32VdJQMXwLZ68X4lizVmw8WR/+Vt/Ed+Rqe1L8dGTiozS0u4
Aau/+d2j6j/trQvcG3PYIy2NgTwOxWTsHHW5yWqljX7AZXtiPBrDNZxzdnVq
PJ+LDszIHa3Dqdjh6+NQfpH5mYejMesFS4TEyYGJJSWR7IeNzGLSoCHcptVv
aBsnO9Sdxx3UbJl7gQJ+wmdB50WyjOHH5aS0PXXEAZ9njCbzNPmya4y/cz5N
XpJob7OVP7p85nCNCB9MFjsiS7vEJG3BprhMvMwdZIB89+pLQ0fDy5BscIlv
apLoBP14oiufvwX24Hoq8WhhKBu+EMpdKSnnI8kALcGmPCjDVF+VNLBpUj85
H6OsqcvlrBCZSs3XrYMsGc/4lEOe8jMOzs/+vpxl9PNoZSBI9OX5dZK5KWx7
8i/x8Iox91QgL3dz2yA/m6xt6hq3EPtgZmOB5iiPhGdcCU99ClLPogkIuGbr
v8ISzo2YXMkbGhdtR8qeAy+FitHFaT1qh0AqTEgGu5wOCJLN0wB8Y1V6j+ci
XgxoNf0IC5T+viztEkEjn3BQxNnyzvTiiI7lACzMTzJRKX2S7S2Bh2sAQZcZ
bABxLVeyH3dr0vQ05h/RL63BvvBc4rOUE2ifnjZN+x2D5pcDVHdmttBgf5Jc
t29IaiPW8MNvE+Pi28NWgASVeJD2spp13/hYJkStHtPMCeWHRvahyBV8irvg
iqmdhvZOVcoZxZWqtVVJS4cSyLlxH3nOpf/iPwpIdvLeyelVc66+HmfBaLxj
aMfubbJ13mHnOFi6V2Vtp6q5J4gW/uzR91L6Cov7kGGBP0zmGhQrV+a5wmZD
yxsOUNV5qQOJoi/xL+lOwo/VYwTcBIHwYsvFFcoERygL7e/zMQSEzbQvGoeW
b87+CgFQTaOWpaIOuhYJDbcTsgcBGP4Px1vaC/1njBayT4ZJDQOw2NFP0/b2
dUlLhlNLmb01AYoTjR4sBhDrgG3A4dIlxh8vZFiZhkNWblD24Jz1c1687AXw
YpsVWKHZn/fwwuI+Qn8//LhBUD+sxMi0+TCTnyyu0Cl7dEoTScehbL9fyylO
tOhCrgFj7TrZvDoHSqhz8T3iMrEidyfc/ygPMrBoa2JmHpPUZ35Gi42Jh8O2
t7L9ja9h20YNyYGjeuTFS0WhCEGGSPCFxFzvD7veXxWFoxuoh0FJ7393OizL
mku23xuSUc+5pIOwE8CBFrT0y5SAvMfBbk04xNxW8f7kxFJdn09Je6RysLhn
XfOb2BSskYhmhKpjilxTkTt179ies6SMIDSpL574Buo6WbIJS/AQpXPbiIB+
yfNWs1aKrR1CZFPz0S7Vaj5wfD5hjcgD1ko/YsK1ndFJbVFWJh+XLjmRfaaR
vB7N0sB2d7+sjrJ3X9ZhuKB9+BnYMbwJgOw2XmDGmaJ+MtSOFvoUkW7Bkh2k
Gq5CCk3ZkVSxBbLw6uADepQoYAOj1oI1DXQIc80fDuG0XVpknrxxllN2L78N
BJadt3xVDybO+wvlEyld/v/8vf2a3szc6E40HupZrl/BDNYj9qebd8+9K7H0
mgdIdgchvN9MfMmrrr4dOHWCQK5pP2HIe1LuRd0Uqm6cHgRtZCPJ1E8IGInL
4jxuRQEWa5z3Bi1NBiVUA47deRrAfzpcwpdAF4CrpM+5gGWDGZS2P7PjVZPC
Ww8RSsf6scKqadmDCrhqsZl9O/6TCYgEY4zm3Tp11Fh9DVB15CFPBUYisAjS
/6vBKim5Xe2cbL7rrg+ZUX1pEHqInvb7vt27vVpVltCXeaqkLE3jY3FJEkF8
y9MmQPgX6irV7beCtIuLJZXJhoG6NQ/qFL5W4WoXvGRiPZ91+IFLf4ybIEJd
85Zve3BfrmRMRu1YJfaSH0dc2cGYnEskf3FBSDSa4IU3zbwICyqpKPAFcoXU
G9GvD4SpcsrxPsrowHl83CgXwnS+ZEk9W7xGrBXfWHhBkulNEx7TEOQ37ERC
0blDd/C1eRGyUWNMTn91GUSh3Rt3fdFJtk1lan0l9EbJyCboTekOvX99SNUd
I9lOBpOR0c5ij5FCCjtRT+IR4+sVCZBXm6+ucq/hKPDvYXp/+KYkWhSS+P0i
QSBNitdEmG7O1BUByYwgab05QJ9pwPbDba8Bq0B/a9PSJLs06dFAyGlDyIPJ
7vyjX+RbC1VuCGJc/LoY4qVRfp3jy5qvsUh4BCei6j/luIl6kOcHHqmLyQW6
s6cmn6SrO8yN9yx66X+MSLHBhY7Lh83waTBtfor7SwOGW/+oaQuZD3kgbukl
1V0xZQhTW6bucPq30E3DckUpyoFlCDuZLQmnt+MaF2Vrnlns9WfBqtd30enJ
I6Fwe76iG8xBks3KfsrT7mcIZcuH8QtKhlhsbqpzI3v/g4LLI0i95yrbl9az
y0LzG4WZdAPoE/xcrOoluy78tqKyUKC+vYYJtIJr089lG7GKDMfl0MCDj8CV
dmF2MYkTrs6hWI2QaxzBDKNhad/a40WnT9sbH1+WAr7h+VwaPexlGTQ+ufqQ
2Op+Jvk5rIGkd+UJUMBFPctN2MLakidZA3Vez/uAMLl9NxfOXnVr9RzxYG32
rfhig262YUrAceWJL1VYVvt251JW1bFdgTHN00GExYvQQP8ePCBbvYVGpvFu
OWqUW5o6rL2mxZI1813S0TYlI6FkEAqveSg8/cS7Kn8kK/hwKLfFP/NxDTU3
U2bapx0haz6m5WEfAq1XhM4oqwhHCzYTFqS+dQcGTNjBJbWENFRKezQVslS5
LXsCi8SbbD06D58NLdoFaVSeNG128vAqFzCJco/c9GmGuFEogc4EK3v1B5vw
raok4TOJfTKs/WR4Z97NNn2GVX8dFa7H39JDCnwogpP90c6D8zbOINd0mIlc
FS/EUiUY4TeUdpTW6msS+81y0u7eeuRwZoA680sIYvc0CMj3eVgZdT+GOJwZ
M3Jrdja+q30d7VRQ8hdPPo7MoxLUqewNwTKI384TN+uxcI0WMiZHMsgFNIpL
nvfhzmLjxfjlyodPoOAYiAzjxnwwZ3jtrr48inoIRbKwTvfQRRGMcVG15Mw+
YkYuzTJgn6/8gxgmWE690JUwk3CcKkLLtCHPvEeuBBu96cjOr5m7Bwxw1qf1
wLdlPjXClst/CDtSn1Qzf6qv30SSWHABZn5n/WydAujDSXLTORYQ9ul2F9io
jbQbPGq71Nnpg+fF5FQhEcPAxr6Bmnd65Oj/JedCUEyjHPrx19i627hI4hgt
gGXbWfnz0veuKaaTEo2BQk7/aye16chbYlduxCgfpEuSoS/AY6Y7y8Z0yiuD
8J+M56SBAbfoIBY6qNuvbc4+2/1RKvpwSGrUaWkYhDoukGqx+jurOWTODnCf
jpJ11820OC0z55XTb0p760PykJQpDOG2TnB+GekwDCK2TL8RzNAb4d3uewXn
cfFVuj+esnZMjV5lNX8wI55z0DTepwXSJICDWX4oZYTTDCQBqc3MBlM/h4km
ifrXECoHHnPZBuPjT+IXdCEYyO3fP8EvK5ZojatxxOEMExTbGNBr5yYLH6iR
s+qn9WZNWheGSFDkP3ds/KfgNR/lR3/ODf5M8YAezQQ8yKPwayte9ODAsM28
Hhim2OEoxYwCPVCAmsG1rrBo/TAqmgH5TiX6OgUkOYocC6F8/i/UYhjwi8EG
VWw3MMD49kn6LsdcDxvx+nInfQ4DZU9gjW6Uxx6qWIaCocLmKzfmhwwU4gAn
SMABF+7UlGIzZYreY8SJg0lA30k/IIqJQMpeGzqn51jsHyzSaqFRwj4AIkei
5F2eP9sP45u9748g7Un750Sjw/1pPEJUh1brLvo17jQp8UClyKZyKju0gWeR
F73E9s/qoWPReBsw55HBbvWcUrukC6sCd3KgYW6CzMhLt9y7ApKEjPQNsfbS
og1foUmiUL4VmI+4PPwJQ8Gvn4nPIl0gU58JzsqYxdibXClgTgqRgYwP18GR
NRCFpKtl04YcULxZ5Xo61/HmM4CfF3wiZBpQ0SP2VhvxIja6aA1yWDLRicJj
CPIeFA+3HkM+hQoxFlfPxKKS5SSWpeFTL4ZZgBo9yRQUV9I7Xwo9IPUAxJRI
rtZN92rfwaCqdaZw8lzFC5I72vmcwYow6wmHOrftiKDpiOxZkubVwfQYteFN
0hxCAVomSwQZSXBSfiyypCkI6VMBeBLB5yeSgD+E0MdgYti4PvjkNS3eFRGZ
ccIrTLBwTwKzGHHcoPJCGGDxqWxdqctIQk68GHdTrBd6Be8H7m0f6Vzi9t2e
rMD00rkOao+WjbOF2M/andbHLwhyzK8m62bP5jBnUd07JiyW6UQr00+/EuW3
rW6lVSP7zo9HeCgBTmixjZAFHaMDUknHLZ87JiHAJDTRve6lfNn/YP9NOlSR
a0rn0trPY+ZqsVowJ/sqTU1byzBM61aZU+VakaTchPA+1wjWzxuH+nikxYHF
Jh6m0V0u41MvYTvzlHJedD1I1h4lU6DG9Oc4hZ5EiPtmdzh8JOtPEmWCWy8w
rJPZc4ZzfbVDIfBU4vTJXtCFJjF2TCZfUpj7wVaVhUi/5l62NYn/w0qKYXli
b6Yrw3ZPGLzRxciVPDVr8ENSGpCDn2wdtj/VFyagxUD9r96mccBDzuL6ITfY
fuO2bAwoa1D+yNmnMqkeYz6PYj4BdBAb87PwlJ32trSue/8+HwogMQ4DThAV
NY9HsxFy7mymX0X2+EVWm9/dg6lkNoj51Rp4T++BQ7sgzrB8IVLDxWuOpSjj
fNAYwFQNNrF2BtQwKlhCzWIkmGRZ+7DlW8ZiHq3p0mmsDS4Ct4GvQUxwe26L
1n0eITY0j/vG4ARf0p2AFePjZ0++8hZJpgtI6Pcf7DNfNBfIBBiujI3pfoWz
SmafVyizeVhBvP6O6SMXnVeTSmP4aUVXrOcNFO/iy4iTGtmseqF5wGOs4oJO
ziw5k09aYclOd8J5w9KpRZzjI0iCQ6X6HydxzpaAXFD0r/MnNsDu8ymlVc2X
axp9ksB4EUvAwqE6De1hzS3iPqg8pRklo3yQ9xI8AU3wckFvfAOaOmEspR1k
UafyNF5lkPnE74gq2OZ214Bqr7uuwCQQ7AqusgOh/cAtH7PzGWSYYD81AfTd
GwCEA2wTgbnK1Tw615W7k4Z7rERMwk88uOn9Rn0BCQbzl1HxEeDmoogPFkRI
Le2z+Wsoim0oYu5aZgLRZjCe74Ys+F7dA6iIZ33kmxVQJWxd5ErB1Lat2cNC
VJO6EMZxJa2f3e1ZZ8XFG06LVgZ9ty5sJA31Ffg9cbg5GpCQKeqF50F06y34
PfqEX5YIJPAnmJQ6uiYlwfa1jYnj67LSUD69HnUyBC8/VEemCBx0ZrL2s/ic
E/pfI5SR8FFAeAkSeB4sPXy/J9G8IcPrtbQ8L34xvdv5X8Apr074MjoJI54r
5XFpuyMpo817VUw+Rh9Ko71FQLZbMrf7ao23HdeupR43kWBJk8rE+rX6Ayo/
KSvn6wdas2DeJ31hKpNNM1X5j3+U4weMzyTBydVaWw+Qx2NBdnquHcBsGlFt
Lx1tMo+KINgCU9nqssnxS+pbMhpDIgslInRYAtHXqWbbYGpdqGqOv5kALdoI
J7y5X5WOSUAMBnLFQWQYtH/CKLzE6aP4d2Hrj51kchG55UHDCTwPD+tOqMN/
n5m34rmVvKYT51728S768Mi0yVbV8kcdHHvCgMF7jb0+3ZE8i5Wq0BzdZFoP
DyvyaNzgylXkRdcE8O/13dvODB60JsBPGozdmOBx0pkP+K1xY2QOZHfChoTk
wEIJRnb6SJH5VT3Ew0ThPZ4IgU9eR5cxTkWNUkypN7BLNxqX9zZ+P22n3ztQ
CTjk8Y4krk84Q9OrDAjR8o0lhQS+GfXAzgaTSZzE6kibnPgfXkmq0EK7BLCL
alFZ0YqMlktq7dVKVqDYxsnFSyW4BImDu5EytK62ZnPnr6+ZuboHDQHEPI4+
AdSFXH1eXlMsIHwNiBRgTHm/Ljk+1Gq/7IeYZYwzn4PEgmAhg1Vz1qPe8ngF
xnNgy6v1tz7Ut+ks31i36p/FUT1fBfoeDIfoCFnZuIaJCpU09c3PxdYF9QFO
27Ob5CXDXMDyf6C6C64ULlJ9YSh6BXARBrJAAcNkv/ZyTm2ku8VcFTCeVVEX
XGNc2VL/3PBo8r47bbQ5bIDs1qG7fUyKdylXapKYXFh8Ip/HtAzUmXc01/Cs
nQVsK0Tv3coMz4cb/9VBR8p4cEWayzzFt0WK4oTuwxniS4goauJ2cK4mCbs3
G0r0rKdBkJuSySq7g8wAg9Eo4IO9gYsCB7C/UZSDx8twt2QPbLHsTe12njkW
1BQ6NYri4GOFEig7n2cj26gp3tuOupczwPi+7mHou0bb6Phixef8fmXYFOj0
zWzZD8lNwFIOvpUgQVDMIanuOpUYWQAsmYH3E6/4v+RgyVULb7neogB4gej9
9xxEskh7nIbwd622JKFoUYT7LFyENNoO+N1YaEpERTtP2sUzpHNpIjO6hWZw
QBRQlDRR8jdtLra1RMGLssyj15GYqSaC8WSjtIoE46SrQJ3skLVtjaKHOVeh
iBBt7K6mcYdGDAuvgCSRyTKffv2hmQJMpGFqCBBm0xsshh2eqVfFVqvUps4g
JV9KZHMbRMZeSs25g9/38qkD9vRuGTlNcI/vm88QTOerCQbBvrxbcu1DKHJ9
khz6SHM5JxVzzbIM9QCqRXCARmtcS7vD0lSwWTW3ZsC5JUTZIiEdkrLQuDbI
jyDKk69zU9jFuzP593TRrPDgh6lrk21TY3GXz0dc0EWCdQBDa+Q+4kaN4/Qo
G96GtAoBwc2nUT+aEyGLGsvCVpOdqc3yjwbd9bVBrLNYqQqVZanr3qo1Q85D
SUXfKgRbKjStnDRC0M9hvUv7x2tbOoNEBXTh6P56u/TU9IgA7Rf5m8aqYVTb
do/fqGXTA1UTKUKKvWkgsy6W4bCRKxNt+w9+YAZzuNesAfICS1GJecX5ms97
PlLxSisOoq4sLmwOiQPJo2RaGkrM6HB+jcJgnD0itCMonNhC/K/MfFWHo4ey
pjF9j4WEtvVBJT1WSo3cW7FN1YXv11FeMHDJ2oJWmRoxKEnOWEWkIIVr5kfk
WZiOwizdDoO8GfBQgG9l5PTl7s8upo0ziQdftI2CkXQ9f/TPvVldZIvYp6Tv
hFo+enXG3mTctSGgeNbS3OdihQ/+1YE9pHAHOeuhHJTpmkBHH8mqcb5XTjMT
qsge11DFedbi70REBsoxLvzRoulvzQYHNUa+VCpZdur9+vt74BBIiV2rVYxD
k5XlZfKlFpNgvmJRTPiihW3yhGdUfl4uwKdCgt1aF0Zgqoqb7L3erDdzSGSE
y9me4tRe/hm2xr0snxGn4BhHIo8EgoADO6dzqda+kyQ3FZkN0Ph5/NqYerQf
zm+xyoHq3niJJMRRPxaczswB3Q+RyUAxmtqdX/yKi3naTPi1pDyeZ7V948eS
8hfFJSeSb+GRXpjGemBfgYssdQb9BmpzJBzTVx+eauiodHg4mVKeKOk+fMwI
Bf+pbyEKuedNBFHRM04/U8nHXw5Vf1VOduKY86oPQhQv5E91FOGsjM2tAwe2
eV4Qo9FEAy0GhF0SYPvGXeESe3as7tlZxidNRIg78WS03Rp0foVxTEgRqUFf
hp9xgCqy/1ZUgY69bsGib8Yaa7nz4TFr9aZdMALZ8chi5odEMGmLHGIdLwcn
qLBkW+k4nlrN6WWC1zMGXVpxSW+Ory4JoFDyiHBR6P3FyXXNv+5cRt2xy5VQ
WOl8KehMOV58NVz7gAJhc1dojxpk8Jon986XZPfyigANr2hTDiGTYXYnLPJQ
tsZUivFSHae/sp/K7RUBBAoeOenrFGzubdDMxMv6XfoyNvNL01SWBE508aeX
L5rY6S8aYo+BhQxTghwtQtPcKuT7Mck0vV6ZJ34XzWxq98eKz7Fftu7t8EM4
GyZFiOTAWcN9WzZG+r3c2MwJAFDHtEC///m4jVpnZMtRf0h5P0oI9qE2gaed
TWY3u7BpDFdgGImdNu4ffahtE+QTpRMbjGSq/aHU7xFCU0KgDfs/MeUGgqpR
vFw6gHH1Z6dw3PRlcCyKKv2+pWtYdXCQPqsKL/UnhyPUdod3kMdLiRY8BtkN
vxmg6xGgWXGNLVruYapKcMeAx/C76fDbyArPUH7mF+h7E9ksqTrVPoT2ClvC
A97h1aPLXHDtK1ejDN54LBOmap3JV+wqwszq/j7NZ1LS973XhtRqICS2jK4g
TmFX6T53+bZFiW7KtRIFIXpKlpa1n/EsMtdOqwkcX+Qz2agldgsnNFm3hMA3
2OXkCHq6LPQR/sluJjKIpxNjXTC+CiQw9MN1+Hn6xPJzrVs7BzLjWzpbWqEs
Rt8yzd9aTmCXrPZrlXf5i23V1swKt82M8neTpRzgslpqAbGV6qyCMu6pAUv9
p/+b0GjD1PLS8fBn+9U00QytuUQ8eqEMKzdggfOd5W322ls4KXatdehJYYMd
ufG30HFLqK2Qnpm82QCMd+lMdFY5inNiO/cSJqjwYuzropLIlpen4NWi1DLc
EoRHl40zvJxq+UCOOw620QcWiAVu/7HPG68rE3yW54JcDBKjw2vnNZtLhjHW
fV8iae5oFzvRrSqMa3mjXqoenlmhd0b/lS4ALVXlRnjCkQepa5mdnuKqvH98
jUQpjZt5YTVA9kO+ePq9fiuFcWZEPNUy05sUfWYtra+sEbvk2I2LSrzCeNuR
ygOJeCkBQDDDe9e2mt6a9+pdenZys+Zqb3uwV0WHLa7gpfBWtM4AHfCv0a0w
lLzjQYcPpgcp+XGl1vJ0xauLVgKkKqcV+xgOmmpEDorkyq0GLsw873iKZWvZ
YbkNNXApEQ4dHmMAC33F7oYKn4l2PlEL48yRKarVBM4U3BKcBgEfL3K2HB2g
7MXMXeDY1crI+814fA0uYKk8yemQCFm475xVl8GrewX/BUJxfyL+XTR6qdjA
IFEm00Q2zwBwgWs/Rci6He0tUcgLwTcuxzQJxcXqpp0v8XZ8CVK2t1axcd8G
g53u1HupFdMZmwfSYGelY8BQ0nPYRACQYJiXJ3nu/u2dajXmMVmwJO8YzRiy
OOCyg28akvkUHJcIy1NkU+I/XF0upYjksE5ulCDQqa3pyJv9APBxFE6s6f/5
h0fM9XQ3s3tYZaJauZRTJ7afw+rRJI7fEf9KrYbkdnpIqXGsMiW4I2V0Un13
7OsABgu0hXWzGE7w3wlsFarLTgIWsElgt03NWfPY9slbM3Ln9599IOe42w3j
gLsMVW4aQ6UbemO6HzQ8WO//gDQ9wJkiq0a48A18T0aCp9KyQscCW3npPbuF
2B1ucJ+varaqiIU94+bkmdzOszQyDt0LgvfmOhlcfLKk9KoWWiVEegEZD8ed
8PzMPFcFAAg77Q8/rrEtgstUyrnuOmWqiEpCZMow1dOBTUr8rsTjsIYqI9wL
SDaj6+6bwrgXwDsDQaP1niYHnbMFRctZZ/cpt8MMRPI5ry1FaE48Jv/RTuLU
NVArhvENdnV3LRz2t3/dcffoK2hH6nLjxVcHJ5ur3r24VXMQk2lenHUsXm33
br7PuHlI919xQYVD5Y7X533itW7yW7MhNcd0pGD/IaGoTmxicXUQcxePSdCl
MaxC0rV7EchY8bGxzL4w2fX9Ccb9NYWjqU5pAtxR3TcmQnrj3hdK8ooBYesg
TT1WaKP9yE0YnVjmWQv0tEyhu76pEPBJ8882OE65MLT/rCxSlUgcM23uFrPf
tJjl4mWBwZWvco1TQHvG+g+bnCp+tVaFhJDR/MOtSUda6jVF1DgDi6YMx+NX
G2GsQTL7auI90cnj5NFbhqzPS+gsRRasxDyDfJgyz7CaVrF0B+By77012HoA
gjVqMwTZ6/AfOp+uFPeu3yUA76vaDS3P+bXXzzYAyNtP17Hg22HeEZzDZLcO
/cjFcNEb3Hs37l+Gnsw1nMg5A2MeyJG+U0QtrEXd86X5wEbZbATeBbfoIQbU
zYnA6S49smbJh8HrNXX0TH4SBwqYb51zQEVbjyVdC8y+8/JVC+MsZw9OqqCA
vHCTGBXK1EbRpwXfbI3h75OsPjRLlrgyyJRSs4W+T7Cxp7iehi+UULBkqrsS
RDfAOZkPQ91DQbwUYsbm+3MNDZTP+2w0NGz0gGFayfs65rPt5200/GjocBDZ
UDaGh3EeC/CKjQbQx6lNvw4cY1UR//YKZceKAbhvkb8wNk7uXRS0jNdqIULF
1lKTuYUgCAfGSnCb/YDSrMSThiVZKr5hBwaRjYs5MEc1IDV7MunzWMazEAZM
7+pzN8D0gDx3madVJgKz4NDiHSOLeJ1mw6y1+9niJk/jfXJz/3A5NiTYejEf
+J/BpLoTH6es8Oz/T+sx3UQMvXU5o1RGTaAm18SyVHBL28NgTZjzF2BlV2sZ
Hrd2TJPXxPJCjFT96wJQ4dHEbRnG1DxznYOSxsMHveO/Hk6y/NWSM1meLIan
9UWP2Jb8Ymi+lbJD+8p98kPGYBV4YoTRjR2kh/oZnKBAdw7GW3szQ77vdeqM
uha8ZI4+W6eSLaQzA8yGrsZP+OCnsnT5JWN0uGUSJGyPZH3jN8NKhbgv86jA
gAVzcmCR7XWk4j/DWMietI/E21fs6zZr04r6iqO0TkeYwZGVOFEMVxcQrQGN
FrMuqI+OmCGveqpOMp9fdSNNRvBr8xuApbNfEQjJ2ABwYoMaAVoh8PhYfnjf
zNvdUt5Ca6JVZWxnMy4sOerw0jVGr4mCa7zUDkGgTPisavEg3IUmZfGqzU1U
LUVEEXaSQDcRvTZdAj2M1t1aBbijBcV9lQ/Mmszyycpv5Ne+OvZZGoAg2RqT
FYPmF5Dq4Tk6SXmAyPsOdkef4h1zSFM4Ml0DK0wX8XBW7gMYob21cu5sAsm6
QFo0c+Zxd8kuCt1BieFcC8M8q5HiWzHypL0vZ7vgWzyz2m2sM+ee6ma0QcWr
sARpdcsTnPAc9+pxI2IslCzL1YUMky40AzlvU2i3A4IuSRlhpXmB3YMhbw44
TfrIH6a31JZtHlkqNXPWw66FrLBZj/43SNj52Z/Rh1uuBIqKMJ46oaPY2tbj
GTFEBL65NqPcB9ubyUKte3uxLaOzE9RHyFYnShARBk/fyNeJXGLU3XCGIgVa
yJGHagzf7loW4l7j2ScewZX9Hy4wLBt3OwH4zYZtop+w1zOtyN7giNrxRkrv
uhv8WCiN/P1psVaq/G7TfFesPVJXxh994EOHguIeVpVDXqzRrPjeQO9OXeZL
Vht3dCDTOFFc1Jrxe8npzvfJxpWHpPLJpdpGaggvqiozgSl5eTyKwX9JBChG
fa6lbNfDH7BhA5sJIIbNhgB6Vv+0lUOwzQkH4d/YlYMep/w79JuA1yqEMjPW
KJ8O231NKEXwPUp4ZcOBrD3JT7qkxYf/NPQyHR2mAccS4dgNkkBDJcmBWWli
AxODN6WOX4TH5EXH/mQyEJehmP0B/rPmU2vjXG32hJ9zbPPYGiMng3iHQCO7
9x+/O6VLDnRlY7Whz4Az2Zf+w29L+inz1O9oTx8CEd/i/kyrymp2hoQ3PnqP
jP/G9ZlJx1ewEJ6KyLdQJqEFInSXWoJmuU7tslYgJ+34/OvZ/cmhqA4h0X4h
nFMBrGJE4VwujIXwwcRvPIcSOfirvD6ckNIW4GMC/oVzrw2NhqZfUMMb6X//
R7L02PfXrrktm4IHI1ipxtJ60wT1Vp9KniP1mp/yIYi9EInOwjX/gPqsPK7c
66vAar6PRx2wZvA40D76WxnWB3nsPP+UX7WIFcjSBYBpzX0Dp77XMszTQxql
eF8L/dvHHAVCINvavN1wpTwH0kR2GTRFa41JUsZWXGD7ewjTf4k7Nu/7fEPy
Qv84JwGzttjR2+QjRBK2lgWHK9N6h4yfTW+mjKZx/nMrS7j/ZxkPu58+EzfQ
2VUAbbZPEac/b1HtgXjh0+9oTyTNGL5doPCB8XcqfFrUqyMr1SoyTFwyiYUr
LpbTjUfYXHegy+iLi+nVTxabKRqEykKAp/vnkLzMsPxBL841pyMLjkt5P6ZF
TsXJMK5WnewIk7yx+TMSIiW9BM95kR6SCjpfsmw4lcd0SAskoopksxj3tOOG
6OWksdO09YVbPhh95vHpRZj5whEtJZIF41u94cJ2wOmEih88Zgjh/GmD+KgM
3BEmUkaARm85Kn3tKWAN6yF3r4XoV/VFOKqJEcz2eXbMnVKCirPN3+C4xEAf
6CzwraCIwxaK0wB8w00jj8GBPdnn4O7hUDz2qiW0naA34Iv5FyUr3QREgYN0
gOatLMjb2RYLs7okbxXkS0CESrp3FvMPtb76snm7XvMjaDuF4qaTyTo3yLWa
AoiS4MNvZz/YzGL/WoTgUyKRJ79EFO+zriS/Z5APad4ePjLF8wlayJYjq/Q5
dCra+Ca3OAsi0uQXuagA8HdwdMBLNdGvaTJ8i+ChGqJgQKj8s8CfN6MHIbQm
dy1nb2A0+D/Ot3uJvLIqDz9tOgNfNcsOfIxONBirp5EgqqBEErDDFvQOeq0V
v9f0JTxq9iY3suVnSKLhbtcbs9lb625OQkUgdngjRCYLIe9h08lzYLJHUBin
wgksI5/wisrxPuEfFlWz7bKqcY8VCOegbo17y2zBdV3Mnbbf9e86zqNVB+Z+
5SNjxkLrVTi/qX49WmxVbjbczm9XMaASKy0raxcauRp4Mus6MF6kdgF+JkWo
Mphl/VFUTYTyFWjL5qHWcd5mMPPzbLkOtOobgYyMkuOrz66F+XMa2MbgCkBB
lAiJYcsVmzlnVgVWagtgt7paXs/SBm7gFe4dk0uChzF6Vz+5mXokDUCYbJR9
Qm21c0Y3EDAQqQpJaN/o7vvbziMyUVXLLVKbVKGJdG5faa6COsf4RUh8x+Mh
C721zsJLbc99TVl4Zc68lSTFGy2V6ok8VhicUXRExiqJgC4OExi/VKF/+Ok1
Giy4IqT1FIOdAg4LsT4vlePsbwwv5Y/kjA4CvYRhw0tWdvJOSvOhWOe2ZG23
Li/B4SMUshnly7T8yW2iQjJigxiVhFFuTEiPn9/L1C8GiPg1xNqPdYe9Eo1b
nfvtH4j5SiiiA/JIuu2PHCqKh22pNFKhtubmmYZMd6KA1xJkLpulq5pS1R4z
MMrBnqq9H+SPjRCmEpmICFJVd8eTp1xnw9dgv0FkAn/pK6cvuWO8F++jUwxi
MUv5dNzmHfSPWLxTYIFmemxEkuw0tFB3geTr9dKHIg2Cd4zYR8k6/UIVB3no
4zkLsalF+m1oafOwKDcWZaqw+CzlK0uSjhvOa6yob+QrDMTlwn5stfsB9PN9
Poq0fsGu2ugn4DdOqvucG0s3j3C7b5ZzszhfyIxuhFi1X012yQsjfmwJptgR
+ZRjFDQ/3zibce8iB2r4fXrtd57uavs44iYzJMmuX+ztg+5mdtzUSMjt2QbO
8VJy1bpbDIaG5P75aRflSorI835GV/XtZEzeR2oP2Dcg1r5EYgwK6l90r/S2
3qEcZIhPkBzjRmH7k0cKbhlIBTEAGHFd3YnOoq5Tr5uyVnnHhdkqVmVFb/Lc
oEVhUlxrZpwatJIO0IEoiv+sVmlCgeigD9Wg3oNH23+uKkVy0/eTYY5kmwG8
aq0Yf8i9iURV9uvI2V79EGP5YMHip3BreTbIK2f97WUaoNXOq+Mnd3zil7k0
9/UuXTPTt6Tt6Xe4OKvMtQ6JxwyqPf8zDiH0WNYK06yse0gnQeUpmrH+VHtg
xAYc3KPWlnUp4u4PK8oWqQDEBIR0UziattNmhKDKB04XyoeCgeBHppLw1G22
rRVjtZF91itbQ16iHJns5lfiCa5EIMpCb4u/+5ztJN6WHVjlhIYeMhqvMneh
2YI56G7rFzrSspzkzr7NYbO7OgU2TGN4V6lDgmbrIKn6sdyFyIXEGkUWX7hD
Gx2Go/k7AZxsqnHEvYQve3rn1WKxNxfp4ic7KLrpY8NZ5kHWqTeEEd1AScpN
/BTePTet7/xCcbkQHyiWZFjBvAluZBPQkEIS6lRvUubxwcwthNbnqIiFbsmT
p6lAuqif/+RIqAcVC5HgAnCBmAARBDvhwiF1g17Z5xmyxoC+0xrKhPNWfY9a
5ek8o1dAOX3yqxSiclURBE/uTM89sp/lDq1Y7tsH+k+hTBb8+8dOl0pc7AA1
pWytVyQX3Fl7vOcD47ycLUztNTOFSrxWjHU7xgpp7mStAPSySvBeFn+vOAdN
rhHBF54alBQUz9YZHfsqkX7T6/zX2Oth/j2hFSsfhu1biHynWgcCVNbd5e/p
XV4Y/NleQEyn17anAKwAhzCA20qmmD8kpii2tyoFQT+C1Ku7MQUgtHxOELeh
ETxgjoAOKtt011qONVnZkUjG4XS3SG/QeoaLrB5mcUApCTiEzUTsG7wFqGpz
sv/QPMV0PDORuGROy0che+lt9Q2GAMumhAztjq80tG2nuh9XPBBlVSod/bw7
6CcdwjQIO1FE/34Jk2o06RqpMEdVb4LkUANZ1OCa/T1aYJJ3mySSzYZmgq9N
RQnfg1vcS7Uo1hTCJPtgMaghxxSGeYXBH48WOpMpaMQXt+zCA/zM5N64z/eD
SsUlF5niynJzmxP1C/AMvFHPGzOoTOv1jl5jKLyLysxsK26MOyRY3CEMc7DI
MbNIRD26wBlIJHUVYttSCsfKN1j2JtkFH9Ef6G+efyPZtiPO6DHZFQP0C4/h
jjslOwPntw8u/jqZucugm2US4fzOQPpBcLuSIjcbMXuS9CYhvDnWTs3K5mOW
1gwZ8t9k1K3xurwbA57Nj3L4q5OlbgPCI1gKjpK/85+B0JU5KAUx4aHkZqEh
bUomct9S5w0Y7PHCie8a/+Jxdst0tPy627dIZM03NfezB2bNAIhlkv27m11/
28MAN46b4QMOrQkoVyb6n1j5NnP4/Xo+oOFL5ZWlbZDYtT+bmAQ6JiljsVLh
aTi+5EsJ6dz8J0fNFr65pLvg5MKit0VjIS1ipuQvMD/Mz5RpWRbncExl4vlJ
RIck4RTBD3JUFbNfor9gXCIi4YcgyWT3dBVPw3ojonKrjVno+dkIXjwmxQpW
sVumO39bkOYERJlZdDwsncXACubo/6x2dab7btxR3BlAIFbTG3Ed4OQwMypz
RRM8lnxuEECmqgjntXJpM/NgMYSWOkIjSt3jI5IRnI2UX3lK1aAv2sNw5OKO
TaK80I7s/ecyICHng8jNPIvT7B1V8xyTtjRb6rDOo29Ha2OPWU7u+W+p4qi3
3E8Uifm+jBvnEt/uNG6Hq/REje5SRkSQ4T73xH7vHOtNQs7q9CMUpDhjDM/e
+VJ+S9YvyHHEkqjO6Twt0tj7HWDyfpcgFigdfBxknEIf5DgxQA5mZa7DV/RH
E1vsfOeBKBgPmvdTR/laM67LGH9XWnJoyPqF7wNTwZ2EmJ36jZE87Q9Vb82x
xJloDZveKcISNmuU6YAi6AlFyXRcuI/RP9KSGuoOHjYyUReM27VHaJ05o9nA
OjOR2WXIQomH0dDAQ+EQwrSZvCehgA8LD1kMU9d31g/vQN5hpAyWV4dUzkI4
h2wVb3eGh61ENEFBNUTNRUkAA9RYAv4+H3sRpe8jx7ew5zYOXi9A8vMLK8PF
0E1LNZsf0CnlW8IchyeScKPPwJomE+AaZ8erEZKcM4QnDY5TyRi3YY3CY3yw
focCygndQSpZc2scRolj5i1qJFHLA+n+KytD3Dsv0h3TYztRpqWN2nY4zTtz
Ivu59DLFtREShNkBccOOjK2afJ4q1gCQbG7s15kevOMHxlGqzZdUmAeP5dpa
/eA5C4nn4k1Y5hopmSywcN2tvpUwh4PK3PxSwkamtxP4fUnrj09NiQRB9O5B
PQkhfL6F9All5r01k/3QEzMcoxYD0URSqaQRLLVw5xMa+qAauu0VxAmUtDxg
1En35ZNHkJw+MyijWUwpqKBGoCNI6rMD/VFzsRhTGgkfzq0YOMhfsqahmrPe
7ScQn3VVRUoG7nCP315uf/aKNXr6pLy91fn29GoF8u7Gv7545ilyFOHLcLRc
d28sRg9F8Hqe7p/NerlxwFarVRKWEcpHGhbkpPDoX8xKlZteSE6Qs2+zdDZr
V1ifCigIdYLMmppdtgSNMTGvXkDXrMKwFLwJz3rRGqrcMBz/esbmzdVdbV+Q
ErvoEHglbQXidk+QhkQXdUJReFqoRxQDJ7Ag9co6A86Q2TX3ojzMPwfdRmzl
3TtvCwRGy145srlHYBH03OKx/q4ftm3r9+RwEPxbCNSemUm3IEJ1htaAwysn
RZTL6lK+11fmxLpArTxFjrGmBobTUj6SwtqbohWBoVD3Zz7nIze9rCZIgBf0
LmzapfjTbt5lY8Ue+rB7ONtgRWllnmgElk1rc6iqKe2QZ3S+XeRgbD/4gWTL
5Dnzq9SFLDqUIWRhvPy3N3CiKnbGAMcPXSIndQU7XocbEI8mllcBJn1Z6QoB
RHiXkxiTo4NhBr6rKOAeuoSA6Jd0C7GdchsOxcSFhAepxuXpzyUWyiw+Cb+u
/78dHDVVbSaxaoxXPSqFrTLHkHRqpmCDll9Q0vRXMZB9o6nHhpJbLZcH0unQ
lMZcYZ0ZRo7NO2ovzyJr7hg42d6cv7d7VQIxc1zbK/MTgPgKGNLa/CBZtL58
hdEo1M8KmNd8l09DoykXV47zQd1R2n5BM69vkmZptnyLovGy0BFZ1r6bLNSz
XlTv7RkpzIWgkxhg0Iir3ekJZ1ULjEmlxG0RUrKFWb7z9RP5n9wNsjhOVQnc
hLvAPOJpjv0qvk6X1IqUyxAPJdWro6HAOGNldXjnXPKFVtEOZJ6iCjH3OpIr
kSweclNZUHNu+7L0hPiJfak4mQ7pwhsGehQ6W3ZdTbNT+5H31lSEli/4yx6x
KwhY/ZEQ1ug/68ZVHQIeTs6BZnLOXSdqZsZGi7F3IhVzrnwFxb0N4pS8Pizg
HGwYdmR2jps8VrIhnv9HuVpK87qLkCIlnhAiHjP1XQujT3KosU61KianWoUM
y1Nd0qdP9cEVxVRnTyK9WjDqE3kfchdQuui2CeDrG9iSSZ6n04+hYR8gGjE3
bmADrhUVw8w+yS4N0QyegCVhPUFSW4PYZQfwRQS0A9eb5s3qEXZXEkLeWdAx
q50/81NJFeBqYxfJU/xbnrWYYD9CB9DQQdTaBCzuEbIKI0hWl2mNXyXBzZXP
0ZOmM/1JcYZR2C6oX043mmVKjm97Xir3Qb+zhsaayc4biLC1B6G6Zkmk5V27
VxPC4/ujSHLpYPS7zXFeIgoslmF/xdhdHzCrquSqkyf77d/28wdDNwliNxlj
pjFCrTwjTDDHRQlE9DQJ8Lsxe3supVTskoxCq6SiPZXg6e2EfAadHSbIU8yQ
LBai8dsCMpIdZNtgUB/Ho5Y5c4iyfeCtJtDCL4RD79d5o0qQQCJ8sh5kgzfL
g1UIuVsv/ImhpWBECanzKKUMSYM46ZM7r/81Ac935xeuitfMLrQmXhAN7Xrx
JzM8xZuun+tRt2UsM0pFlwAXd2VzJn+HGlIAMzqjGce23H58a78mLxaP63K8
jR0MKdHywJOpt8tS7n3fyUV6YRIl83UtUGMexZwgSkUQeY9wHN/FiTtcGFCi
D/83+aAup/Xqo9gbN9q+PlFI/6SIIqf2JpBWh9N+Y7gz8s3TyFJ+xT8djHQ+
RIAOP4aATy7ukmi7H1wHUEXd3LHVzbohAcVJn9jG2T/AFwbCIflzD0yOkCt5
ffVnZ0TSc9hHpO/wl9Ra6Mk1aX7aJe9u5fLP7xkroyjDmrY+H/0DjkI+IIvI
wIEwB4+PKUG7qt+sk40MrI24GsLZkZixn7QxaIIpo1iJCDAsu2bIxwGTRuOG
hcyqOmDK7qALToBPsB+1zV0B37kJYwIC8T5amfDnGhOpCLGjmcXMHPHy+CM6
v4Nbg5aodqacKlLI6Z/Ej5hS7CibdcrmOGWBsIcDMsbwSUDamw0LfB1q9Dpu
qO4K80lZHhkv/8d9gID2f0oJYDs+/1qmOXgmquDft9quy6txqZCKJnH01qAa
ssC8QqVfwGPrTQXrFQOR/CT/CmFwDVZFdn9NY9sp33VWU8YWFUxhIVL5gSl8
UulTmv+ubjZLTq+FBrJ1zyW5gZqmyy0EN9BPJMZSEnjGb2ASbI7mJPISce6C
jmiTFZj9jYCvhRVW0Dd1OT/gSzWxpuz8YmhAxT0Ci82xlZcnv8YjB3jTCN7X
XCF8Ls6W0tiK+UUPNiFZpug5KJ1bqHRuY+8BaQKBRORaX9Brs1sMDBrZc7lj
KMd4I1wKatKxBkWfQlLqKj5DkVkvdejyH9+lw2XDII78tPAWoSBRSw3PyAzw
ll7zv01olEP/OiiK3wIRrsTpIGutDv0QCaWVRFl5itFOSKINeEh5ONI7nsoU
G/gCQpqXhF81dfQcgr8YaDSZktUt0uoAmwr/Fm7lnSnfjmkGkj4e/lXHyeVp
V1vvlg7LR4a6KyNp0cTnl1X8BYFDSK1utaZb8IEAxwzdevK/YWkR3fgiFdYP
FZbA8lZyIJFTH5l/LXMfURG4KCgKlct4NOjJLb/mXLBTauccRkcgqGlIoHoc
lPm9OOBb/LfAWTGK/C+PQ13efcVfeaE0a1ZmdEIruZXrwLGOvTCvgSR+A1lA
gY4tdh4tkQlSeIXzrbJqyFSSfTIBTlSSy6vdwpdP3M8YX3In5hIFPkG3W12K
UOkleV/EDu4YwNJ6K49JbRoOXS+U7BTqg93c6h3/QLQyY2Jdiu6vHIwD+9V+
GtZeAZ0hGoqe1CvZ2YZr4zVbFv7SyJbG1Gl9m5we2HqmclWBu3XLY4ew0H+k
29rOngIv65duuOp4zc8M/g7Ux9o9gbj8Vo2JZbpcUBELZy0A4aB56FXMtS5I
iflIhfDpirQt0IDdmq/k9gEcXrlqosUIhgM3/6oOaD1R7tv6tie8B0bPbyu0
EyVT+5Tvr6+kRj4RVkBxPdHAY4HZNxwV58mfT3s+hJsy9/oF36J0JQRgyy0c
Fp4+RL040YvQGnXBHX9gwrWl55mcJ6WAYf0WEHTVC99MF5g04q3F85xjTqM8
fVgN1wYLNGiMrn7lT0qXvibUVRDY/8KO2RXNkyD3V9hqUbTpFZny+WRZsES7
51FCxsYtPEWl8JF64UJ6UhAbt855aB98/UrLeF4Fmx9hluM7Sv3VO/G6LF5k
7FFmTyHWEtqnS4Mxl1wOdwZdth0nCduwSjyqI7epdUM5S3mgm7EaL6TiEHsq
vwXJWZuidKlRRtZ+WywzmiV6AbefTElPjJn7kuRPqUlil8auyIFf3804oYhp
cRe5slMuhoNic0RkhBzrOwCxNueRdM98a9dvOGyXl+F4mOfu+33e6N2E9Ab6
MScOOp3FyIVvdXn0WRBwDQ81ItYg/zcE5Ce8/G/fatghZU2Pgb3IlMRvB6BX
5Xorf6tO4/hqDx8Xf49nFLK0qcabfUQkk20HXQuFzfAfIZt5kNyunJ/JSYty
WZbYbr8M7whIEOGygKROLbea/BOUIrHHuW9KH0Gr/+xQg+YQ3hZPjTlntX6y
5JiSnSYaoT2h5XfBQB3mwm6t9l4R9cOga/1bB4ZbO0V3cqUnjmD7Vd0vINsK
o3hZeY1S2pu1jSEiTj4+0JoZn16TTFuC9eThkw9gYhKTFguGkYUtiE1kyj0I
Og/i5555LfrkuuNdsnhgDaRVA6QkIoEeSYayGXRSfdaIs7WvZ+6W8Oo2Q+Mt
455aS+kRSnaz84/Q2mOmSqZQ7tUHZxqIHRVyfjnxh4DR1bDzgs1qtId/s/Ie
gEUru/9/JyDhv62Pg4/ZT4huZJ+aDtT7EJ2lcOcILpmcZy0JcNOwF4l9ZGVN
e2YNBEfBNN1iFSirdio99YeF0zs1nabfm8xCKFazQCR5V73QD5hLUYtnCSDw
OF/kbdyqndBmRZ8vo5vJlaIaM+D8uXzOCQRfPAxJIqAgExKm+30wEzANdQvf
8XHzAf2DBdUz1EQmluQmrw02FgKj3hqv85DPcdpqv40vkbyI6c/7aWoV7EBc
XQ5m7DrUzb/CcxtmpC0+dZ4dyGqtV9c+urNNWvO0Aa0QnDeF0/O/qG0ufL80
2Na0AqUhW1rOmkMNV094pOIi+WJTh5v08Jq1ONxVNq8k9v9+sq5p167EnlW9
rjjsUzRom0JDniYQJAjoCaKftjmrv6XApsAbkF97b+ulxUbGnrXE9h+VImGh
iIvnFfIQZcnCJFVt3UDPktyPLqMFXGtVUwtlhr1/jW1VMZgVUhJUTNnwnocE
P2V2/qz41+Y0PI14i7fF7wawNG9LECBoaQJvNHI7nEsJfkhI8amBZOIGc4E4
1Sh2qKgu/BPLITvX5UHXJxjSPFaz11xNU5hAnn/0axy8Sy4L+wwvpzEO6MyD
qaa209v7qAy7vZ6VVNyGUY/Di7PZ6qnrSiisEmHF7jFRoGwUrr6NixBNkic6
1ZOjWY/hzMOE3VFClTdsxXHb1p2EQNEzxaQVr2NG1RmbtEmaLm7/WwIHsAWK
A+wf2vPgGdd9Me+1BRkFxgGS0QgBmnzgzZUgrdcQatvcRoc2rFuqagmQBRqA
01FnZCdyaSoqXPir5z2r1n88oQyphxbcTdt0NufZxf82NAX+rWevtoLfsn/p
6DpBySwM8neGivxLowL2BMFp50aWcUb0GWVSHamTBFORH11n9Sn7Vkw22yYH
5HU3w4hQTOjx9jmmBE3l6oVULy5UTAgQHscB7mjngKEN+WgpYVxJdIGhU1N+
xlingGQv28WQowANeMlHmqGLhSyn6+CBwzQKl/zH5GmlR3aIvEhqWUpDyur5
DtQ8fZ3yon+i1DJzLbn0CdCcQmuM3MPsdkHgb7reHGiw0jjoUSzCST66e3H1
PpASjE2OV/UaZ7puqar33iR+AunmFRXUQsdRGX9MfmfIFnrjfiQ2KtshcNPD
7gfF15wAHT8BrDPSVBEbgbChAlPOv3rneO+dun3MhFIVrx6DwyE5scn14tCb
9hA62w9NHh965d/J04EUKV3O64pon5qgDjflWoDOKESWYmXsnxA5Ib/b8EDM
96nDzANJvh5Q5HEF4ZHSCt0sPLYUWnR3iuw1V+/N9DzI+jsVxrXs76kEgQpy
UFXcflglPYTydoluYPn8K1hrgmbG3hOQe6/1gWHLZebud6SvvWYvdu/2SUcR
XnXYboo+rzS0vwoZKFiexNY73U2XjwwYbJdECs13wErRVVgY8hzZ5LOR/ejg
7ngelkqBHCp5pVxFKahO3CA234IJBn9G2Md8Vrlf2JXhi0PLGCtD3kJgL7yx
x8/5TVmDEtAd7+rw8F7nyWkiCzxXq1/6juQmp1cO7oS0n0/Cbj+NDzDpzNmR
hNFhP+VEtN/wqKALtRbEpaisrbFh/hPayAe3ViDu4zN+kSnATXb/Aan3l7py
lC+5eWx7G0ctT0mb1nrr6K45DuOaoEdrSsCppbu1x60266C1jbJz70XkAH3f
ZkMvDc9fgaWDawsx3i1vKdQ1smLT4BMPJVuVMm4fpym/7umxYVj+kjbuRJmp
GZ+WBiOZd+B68cZbjogmnUcrjDhfqpBXbWgH1q8sBbTcDd/6fOCVs9QFGuFc
vBcoT03SoL5H9KKXbdDNPc18LsX1qOXMq5kvvNixA3RFHbWGuH+idOPXomiP
iDKwO5c3r0nKBebxtPqqWjQ5H+Q/48mcJdrfWiGLxNU1fKN5dNIFmYqy1bxY
bFwde/SxtqM95mHLoSHbYi6cwV2xfn7qTdnmiaZUXUrtzevohsIifFXnsP0Z
DIZc01TYE/0Aal7tSgtzLbAKrXLNSRzb7Wvb+qcbYuqlGv3+GDJgMXt8nHnm
p3sDNFXfRpjU0KM+1q1bqp+/FPiiwqJ7keSU41z3JlQSH+/MUKchuzpIdvsZ
ap58cApkcE3g8en92RNnQaZVW4gCr/tJgkNJdr5Kq7j3pbJmWEGeh5tNmlLj
EzsFOw1MHswvhz2KOok6GJEqFF9DZimRaIwod5QRrXkW0jqV6/rAuVL/dWLN
JM7/2PpTIUJ/c6PNBwZ38cdvNNpJW8k3veBliHbiuwe4cly5+MfbnVqLxaFT
Hsd2mjtBbHFOLAOFGsY6w8k4T45/+aYXXaUncl6hrtZgiwc05RPx3ld4SYwI
hemy77QN8ifgeBjJkDoDaD6cMtBKbm9QYtt44UToE+bzJ15MuxMJrUy3Di8m
Ggm4xl87gAuTKUtYrEFqbhyKUmMOzKVITPMUrZGNskf3h5CqrfPhRD1HfXW8
melNw7OA2xgZx5LCwJ/W4qhx0jjFy/enqKv4ktM2jRinmGZxmuY/qussaKYM
lRjm36vPYdbYFb8RXLIKP4p9msXSJZFpdKQac/pRTwpvVej3blt9H9lG0zy1
6ucFZPbrI/4jeUKXogpKdRJXQDsthpr6ZkHch6O1PljLOw4VaaMb860OAM9B
O6gToeJ2ik76rFd+rr6IVo7t7k3Nz4YSkarUlYq2r7GGtW0JajRHlkU71i1s
oxqc6Bb4mhhpcjE6ydWRjMqhp8a/lg7TVebbNsiglfCM6Fap04iQ0MTtyaHe
pz7zMhU//MANbJ/GVTvjxDNX8+nW1UxS/8e/W7ZxMPdmsUJwYaaTuuLl0eGq
EM5k4so8QA5PyqF0XYS2nKwCjEo4GPFt9qaQ1UbMqV4VOGJOPxka8fyBdBVW
8ug8bBAJLsP+3syJg7aU89/m3Hos6sXblV+yEeqTnC6S065KmR1QpUVobE7d
Jar3+zbgT1p6caoTKtfuR4WxKwuLfWgMertl5cckwQlxVAngDC9G8orLs7F7
0jd0FTub9MXfxxjXXtbEfjpVNVzqTEhpG/Z6g6bPNPLDNyhWRRbkgzptmf2B
YVb9flY+PyYvjNt2f1BVxPhqLQSuF5yjmysSEGx1SfF2GCYgk7J23g/QOhoO
fuIxMtGALSQznp5DmJbu+ag++7cG/fiNyNKYxQwpIbuFhFHMtG2tvEpzUcES
Em0Hacjk+iYi8ztnHwppVHnCC6d4LZOulTlgKLbu3QxeRC5fQ7bu8QcafTC0
/UI8U06/w1YOCj0+mx8IAPIrsPWKG+0aSb887e+1n4KqOOMm18rSS06lliv6
YOH3FLSWpQCugKUAxHur1byB1zNEcyBInK+4UTYe5AR90RnzLYum+UhZNM7p
j0HripDIYiLc11vE9H6eUClSdp1LNWflOUDEp0ljeYFt2OwuG97cv4iDnrZh
LLvX/UclX/gCZr7fdz4kKMJ9YBGn5wt/GPlgqfEiyU80hx0bUCvRrH96LDwh
FwCiPY5OLJfXBVjQZfYy6Zb/aUa56aQe9JlSltoOJbKK4ZqHHnEI1wh6VoyY
dBNO7hSv7zfOcFGSwHyp8riPysQo798Sj89khtAP/VHg1/B9rrt/LBU9lS8a
XQTAndtJFYYjUSTCJ0cbIKq14lSlXSWUVRPmGdfOMfnUC0MUBOs+9CRxNJNY
xkeqde7MiiYKuaKSj2pIKMbgK0zIED7QrxJBssOcBegZenfEbtpQQeAxU4Pf
zOFAe1EgktEGcu1b+yBW/NXMc1Sk/GIv1yjmdwaQpd5Pt+VQYMSl0ueNYFuJ
4ZKiWmn8P1ivQ69L6GKNcjPtm1/zP4721VHF5s8ARUwDiYl1fKDcvf4gBuXD
ULL1bG1pr2YEfRv3h/ypxdCfuq/VDXLrx1HIHr/kfwUf1Irj/xq3mF2G9mKa
t4Y5sFUHflj2KmYfx6iHuC3eGngXj8rkQnfdFNwWwGeAtVuXQyd805XvOTwU
dKlQ6UuFtFf2JMMIBASQioY4ui9dwzvnQnQwH+ZYiWB2XLWGOsVQaXji8FnC
d4ICMKAFPvugn/XsRX4MUCOeyUxg84M/ruvVxIb4p/TU4JeXrTPYFLfFXJ2Y
UST45o3bf2vkeB1bkXyed4LfXcZUtrmbZGOuK1OdBZ0qROKXrP/uyBMPe1HS
w5qHBy6sTIIHRimD9H9Ympgy101DnqqX2KsrBQRTClQFtwOO0q2lyEqYhRf+
gVY37Gf8pdUkO/2tzHBNoIN48IgDvvJ4IBql8w0GpQ31r5RwHSEdi4tmEPNF
VTUEkCJQGMJlPGBJpBnbVFNDdaxd/9RBw4wf/IJedyLgf3+ttSEIq+oN07Ys
wuo3YXFVH7fZdPP1v3v+ye1w2Jl5seJKJ3HkatExTMbnsmOepnRQRNMzCnF+
WiEP8j9mwFVg228nq/D4gdP0BXLkP5ZWMjaIm5Y27Sl4PTKMh9fXXdKBxF+r
zWjN5MW9M2Q/FPNHPEe2Xb4TcuQAkp6uAXWff23JKSkGk9wE+i9fGcSk1Hsh
MOx/KjzLykY9mp7XfH8AeTNuMzm4VND2bHL2L6ZvGpWNxsW5gw059NgP45Ia
D7Ft8Kpye3729AMYVEXt6DUtOCzZTgI4esMrBmd97b6GKY+jv3ynePtdbAKc
NatvMd8GHtywztpTfrNRr96JFPovSOzByJAFkoEVBg4LVX6uqh/B7KIYu7Mv
I1YWfDnkgifFdutAhfFIkyHP7MQtrKqfhC9AdZSAFRidyo9xG3rHZ9gQHYtc
cpCtFqm29zAkBH3XXhq4LrdmJDBF5cNieWpQgMWcN/uHEGLYKNsqIGNnWXoj
5qhuplgvvN9982+0T3cg86QbVo+bOTZCViDxLMxJFzuYuDEzB0153VcyzaNo
68tNFHsOnI3lVWXZnvuceAY0Qpk0DPiB61DqnEo9jQyP30C/ogxXn6NZHlau
RFqYu1rt8USATrp1ePG+9OxHpacRgRdaXlMtx5MeRBKleV1Mairqxi0Xcn8N
vBQ/ltPC5EvTBBwL3EKGjUOUINmeSGRUIzwZRNhdR2Gc9b9gkulgnwhaENs4
ieE9UrQ5Mq2y+THKMXhk9vMLuVZDFpWBSVGxE3AWhAXISzYAJlJRgA4ZbJwi
FA8YwvPfxJFUE6SpjIQxLxQ7LZiM0di3bhSTcKGDT+oHZXcrE1CcBC5fB2mo
nD9AQhu+PVlmmAzklXr3qcGUcW+c1xRzFES0gbPLW0iS7SSL2NuVdby5uQzx
FGa6pMBuNxQYvg5B0AYVVQdOFDIv22d6LCp+EchtSjou2bCJFSQmHKvZgrlv
6VRM3Gtmo2knOQ6S4kJbaHO8tWo6qgJMq35SISyFHgCEonAIfFQPEAz0IIG9
aW/qIxTXrVofj2G+z/qSSFLhYdK1qkmFGr7ektMJVOTT+yqTBsMKhsg/SI1U
OdS2E3ovcZFYjH3XjQ0w35dYBJs7F9p2ac1s8wZTtRsvtj2AZfwCY1NyqAWp
xKBQaLsD+B2/GTz1PqwNwtV/2f07ILSI4CoUNe3OHWgqeQ44OE4yB+SDn+va
QV4vF/gceQ/qkAA8+mAkTSxlvxabrjcEAJwdl5K3fQMxQYPspoYgBdDkqVj6
xcUVTlLugQXdy6bm0QmFoQHRGs8n2HpegntqQyY3O/X7LF+Iq0DYgsuc5K69
7XrO+VrzTnTiIk9kG0sklaVdlh/Drn9WLC/XQv2rctM+9DPxqj5bx5v6wbQ1
LU4fCf3V0KPlD3j/YK5EYI+Q3Ms39G06GHGclYbIY1iOlaXqXgA8Ha/sJaXw
EnOHIaCQpuCcSoBF72WRR8zkbUgMosHDVARgcIxpwwZXNhHM4wOBtYglOBUG
EyMDDQJ2J9O14upo1ezkTpOrePqZbLjNdwmMqrY9eECPgafOsq2Zhc6v43hJ
QA/MmPaXDw8FLlVgybTwCFhtSk3i8rbugNOtUOOlqB4XDLQVKMX5p+W+0Q1v
naCI/2ojy6D6XRcOkfY0ZgKCuaNta2+ra710GBPdHLm160LUbnhZA2UPMBBp
9xbkwAN64OSM2on5Hx6/YOgOv+7BkgSyVvkxztouBfdRmp2RsiNBT6yiZvmd
MOVna/KhYimrndA3w37Fu/xVHarL1tSQJVFg6jtL0zohPEaFXe31raxsPKAt
E9NkQrDS6TWK4axSyj3xTqZXHR2oTyCwyiFwmzWocbhhwVRRgyB6zI7ueoNn
UMXHKob9EWaQuVCQ39EBV9baGsnUFQoiXQuPewX3V6xYwj0lE+0PvRUWbGvc
heg9bDwCL7/JTj91uHowdpdJzIn6snRYvznyx+a40Zs7dOgThHnbEL8Y9UeI
BKt4xi64N6a03R7W5nQ94IXx40A3X6bGxcLPTCALNWuoYz3z+AX/Jz31KhLd
jvOrIJkBtW8HL/jsbqUzd1ivyMYCeo8pLDyOEj/cQIfxNO2rTjd4niUVWocd
3LIImHSTeFz2v23yMxQqkpFApYGzKp1DXydQdePH+Ij2CEtBLcX1vS9i1zl1
k9zIMjH317fzg74RhqArCEvyEWtjI2ePLpRGlDWafq1spDG/vPl5XRV8peeS
wTz0ggPWVgeEQTuR1lSJJ8nMue1cSED+lMjZPGGVfM5FtVlX5dZV9nRu4EVb
/KWeKXAS4NbAnGUZvmysvBxwHNIhebPjg0Brg1PZIwIg9T2W5JfZi8/MyyKO
vZXDZ2+5eOxSR5OdtW6DrM/ZKNEJUsj3142vBuSuWjDzmQRh7zwR+VND9p2s
uGr6YAki+Uxsqa2giwUu90hpYgb0KK8vEWqpaXX8z6s7rwOQDGT2vfEHu+DK
VC1E4MZteuV0EJnYZx5H2wqgKfMQfjEYo4rgn/FKKQIv8eh8LcZqM7TJuj9i
A0rUdoRTWQjaaJUWANsRVe4DYkKgdfCEeaoN31bNL3BNH2x0ZIs3Vjik8WDt
KRKFpAhtEX8phTQZhH0YTt9e1ZPmWh+5rRLb+9CWcNqoBaYO4Iw5OYTRPie7
DEFUAUSpMWye2N253KVbCFlMArVBOa40K1NgJPqyMIfk3pAYylaPODdAx/UO
ShP7Qjj8z08ZAMrBcHFcA8mZ6Nsy2rpSLYLfMsGA0WnnRKdTzpc1FrRUow44
BT1nBnSalz6GVCXsOcHYWoWCpOxEQtlyEZMkBeck+NW3t6ApttKxxEyZlxXh
N52KbNHWtQ/bwaCSjZFLhR6HbDvY3Gkr5VxXlGeYL3Ncr8rRhgr9NYHAxH/e
5Qq6ScECkskhqA7fc9DhMST6pAYJm2kzzdcKH8Smuzj3LmmnLF+W/YNlaZri
KObFWuneJZvDz7VLLB5YCFCsuzdUZuQsVD13kfKwJuiBOIhsuVyOPmKy6xua
D4nd3VVTJ/e5Yvre/XJC37WGlBirmqgWZ8GnxQdaguYXk1pbRZgbis632nRL
XKSSH+4+k6WaXYwUg/8UVgJPfahCqhC4iXuDloz0IQ+s1Vu6oXCJWT/ixh1D
ficFvcDMjMzcSvKfQx8rVUiEsxmVJ96e+9/XFn5nl9P9T3UI3GWJvMP9gVS9
zTOSZ5LQ6+0TelXjZY90vq90P7M3GUrMrnyKLNf2wGxfU3yuUr71jYNS3wEk
v8TMjOEaYGQU+x/oDqG7rrKldKMa3Kf94SnfzazSyNHj6N1bmz5ZGUw04fgC
9RtzMmhrxC9TXB0JYiNOf5YxyVK9ruoDx/OGn4aRCTfwhUgAlinQTeR9+hsw
neNnx7rC1tOYxmLnYEWkq7i+u5/EbQZmUE7roNMBR2cHPz17jRFIecitlupa
hfwKKAdvGkJJU2lvDlSm55igGw4V6PC0Jr8eehv/1cdG9zimHqC82jeSHfNf
847qtLbvXJVZbg8320+kz7K/aXv3ueyqkHiVjLxW29ect6xcJXnp0Y01cZEM
HkKcdhin1TUjZQXiCQrhSP1vpDEkRNGS61RTkKlqO6rDR58X+Ji25AcAtVhv
A8b4CJCsJqKW9q3M7Odz9hvsIMFB+iFhfQjykAfI9oyX/SSHCbM1jXmprJQ5
bfBXPXlOoq9taPOfzHrWl0I+qLeJLMGfCkIySp+thCDHOEA0m+YHcKia4k5M
LJrXv6eRDFi1HT4zy+miBXdskoFd81vNpZgYIjU4K0dG7CZt8frjOuA07Ikh
B+1ES5//AxLn8/9lNKGa3vN9nsuX/Ii4YvWL0LeDoYiIEnw8k+jsA2W12p9o
JGTjZsjMtnFzEtxs2slCzewm4O+36hM2dT9XPQ9dA9hzU9ndpqpUW89KXwN0
r9UKqWzhnyK5PTGbxv60lAiBpDGyr6vSFx2WEyEaSpyC2eZdFb45dD4cj3rt
OFPmuCnURYK+U5fcWZB7eC1rZQ41aNmpjoioQC+WufbkOhtIa6fWRgODNd4n
GYAFPubY1dNRXkaL/yurLKi6e0VIk8YKoVlDP4nf3fTfKJWrBxLtHX/Uj7/c
gXbORkHASTso1WdUnxLkaUFBkkGvkriNpICSsCXXdI5tFR5wzM6YEUjM/y3N
P9ZRz3wBtKoyb30zRLZV86IiLt90QUqflfhrxk+TvHnNURl2T0G2GQy99R7S
tT9NUZg/Q/mKq8/zzH2ztGJtHQqApGLiP8Oq2U2vMwWl53eJpIk6y7fOscLK
G7O9uL4sm3elw889DSGPH39OJUPVwM8poX7+8sys9q4a2lgZKTpVp6DWTur+
lu6IcZiN6Er8cYzH7bk0iEIjVhbQdr7Fjj4gLiBTp/K0JUMRepACbI+iPgvJ
Q+ntV7g2xcynMlVXrGFZdUcXb/9OMSFucDcTvWz2ZaJJbkWpOOABbyXdEjTI
u+70CnB51nNTiUXGDskdDFD6PkwTHsFSRJYHokbh99XdmgsloBDdyWsnEkAd
b7fGiSMQL0BYvMbQqLq6LTziUwIru+4JLhiTx9TO8HC59hS+oepDYfotONLb
ouy/eQHOiQ0U/+g85+jdubsJqeX/go0OCZ2nXsOGnPwB0zXU6JkIdgrtrc7A
GuTbP7ehMx8oFt07CX3spKdYVHIjh8B2h4Gh/cw61gkgRJWw2T1LPbU5pX6m
h0gpJtW86v7edmim9WQN6inV29DCFwJh3WSR5FT1wKVEdW2/4aw2YA7U56kX
fPCZ9MJAMkNuKhxpbswyvqmOUrDGn+WxhA+TwekRWhI15AfazvO1/gi/wTRl
jjRKpg9/3zls5ouJJSA7vQG6RVHczZ/M+SOngCuBRdGym6naM8AoEDWqUYbY
RiUs4/5GhN8lbXZ1Z/JpqRoN1RXyDaB4hU018UypkD/xTH0pBX8JA6CFJzjE
C02YeZcOCjiM3cPru1Aib9+t23qmd6dlunwzEACvzk4o6Bmw43RlGSvn6rOW
jbT6K/jtXqT71FHJUr4oNOEzulf+8tCF7UddKoCs4Umw5dokoMlYpcoTSmop
bEKMad725CXcUR9wEc8xGZmSXFSZsG65y/novmzjHNJpfjjJLe0Z9NJG9kh0
3SgZ5ORiTMMMzQKsvU2FMbcsDRSgRInJ2lTkwHaTbnlwlwDeJjp+V3gcZwRk
kMH76K4F90kxNe7MrCeGaM2eUk41gsIOWTgtHIjWWj6JaYCFoAh5WWmW1U0x
QYqGbo94t8iIiXFdhsHKU/MN3NySiMti7mGcjQjNCo7INxLdn1ISy5mit4Mm
r/bN3MP0b46HoxlpGplOYKuPVjho6BdtaZ+xfPv3R4Cq4McPFPYmnTMSspEr
FqQr1XQoDR/c4YGY7M1auyErWIh7XZg2WOQlIjUu3a16ZL9U2AqfbDcOzPol
DyAtb6TZ6i+eBmQB4JgGS1lHn3FbbNPeBvJKjx1ipbahvNCU6c75dqqBH3XJ
5knbUYC7CDfVV0JxKjQi34IuRO+0BBdyXK+F96/AgHybYg1iITgbvJ0ZrqEy
ZtRjvaRLyp/4sqw7hii0d65i7v4rlx/DsbdpJRAYb80aE+uJwibe7k1TFKCz
IO0j/X4ASDe71rJ7fvUG237hKY5UEcOLBkshKOxzyLRRmnZlpfwTedDR5kzU
oCmx0CHWNB5PtQgtkpM2FwNXKKiJCFlRBiCwiDON6H8CY8q0MZ0pFyEqpURH
BZUhw9CUPprqOyt32Dkddqp56lH38yvmlZaSy3GfAyzuo8TeeNWRs0P1TEX4
lKYk4lVF5PSkUrTdMK64cBOYzVyIpn5kYx+DoW5i71mak8twVHxav4DiH3q3
TY+Fyny5X2YycgctL6EohXVSckNhI1b8Bpq7jIjf6DPL2uV0wtv8mh9pyVI6
AJBKSdVeu0McJoZPeSX4HRwZxOcKDQCdsaxgXo1o9N+ZQXPvq0lqHJPpap1S
isQkvL623knKIGwl4EYpYGIoTF/v02NxqytXCh1E7rPPHiywFpQ6CZt7KacH
iM3De0bPRHjKgw2FLreZxVD1yXs5bRyio7BGZRyG1+dcM0DetRsjZW4wu/iL
8u8FxIo3jWGD5q7EvRQL7aQEMWXWeDHCWT/EDiXEHCdbZIpRq46rhX9EWCy/
deB9+xXy8GI3StuTLr7ix0YxzilvZDSEfzWRNEbK1ST7HyMnmBCqqPqwjGyn
yRBO28Zx+ft1BdWlIyPTd4KJXOSVnLS5rxqPXYQ2flP9k86O3gr1/ggSk//S
ZJhMmlCaouAUlg7JyAp1MJVtR941mp4iNLh9QczWJJ7JIwVDiQ52Fhvc4Ycr
u52cCjq5Q2LxIRHMSqkpAJhC6SWdGLWS2eKXOG2aScBo3emx9kak99NTaBmK
9fyZjO3p39DpXoi0XSSJSpkkZJjF5A9/lcltUeyCsyHxFHD3PvS/ZerVKduG
Dqjx6Pqn3Ldg7U6YRYS222DHzCqbpzLN/2XUVcxgUqID0N0ctHFcUf/Xy5Co
oTeZrxA2bl5Wz30m3scKDjMC6FPsigxp46/Uy8QHUMebeOnLyfB5o/UaJjh/
WOnHBBQ3kMBCQXMawDTXLmuanFC4GLv/gr+uFA0FMqpaybhmvWKRxyxR98n4
auK1pX+Ne9yrSmVMZbV/TQmKKvRwI2PZ/YuVBGM9RzLnOzW0f4pmM54AM/uM
E0uatZaF19GKuNS5blsaV6EOrRDLJ3E3bDGhBER0yVv9bpWt+UxKUumxFZDM
kolJ0FQoYYDN8pw1MKHKpPDotMLPA6BYfqgYt9nfdLJyHFeWb4P/JyJM1Prm
D+9cISQt/0Bvgz8er22hRvcSSvGVeFntMaMuX0W+Z3/6dgKPZch+I+2lfqae
YTQKlVduXPgjEElGq8IQQF5tkVpVFXVCLN0CGwtxqyNtuemNjH0TTCms3nmz
NC1/U0j8SlAtFB39hhea38bbNTQIvBBGZKvMVSBjU/fkLEke2rv+xfxsWq2O
PDmP0vCNL58iwknB1gEb43E0NLxVU9r7AYkiyDk2QmL/UKdQYCqx4wS9NwRY
lE/Ga0XqWeahDv/ATEBIzsij0ua/yD1NMsztM2bUGkd+0r++mQlDm9/4wdKm
H42lNswP+moBfApivnrrqRkZMIV4SRuN73RNDZ4EPeTq77MYsDseV0x+DTT8
xJmMCDQourfhprRLIlMjiLMWX406bqAIloCOQ3da6X0FtgLwlJ2xamFuh4yS
ImDkOZTd8pldHzA/Vi5TXczxSyrVPjd2c4M0RdA4P1oh6IFRFhvLfZsHmLjz
78xjv+QGbI04XlGemH/NPu7XxhLDfMTOHVq//lSbFyKTHZWGNsmPe4JOwFJy
F6mGRMYr6aZnzmZ2GuMxxI023GjJH2XcW/IjV4z44dSpnCRLjNnoBDFyaGQA
c5T4K7YJLmoMA666XQkiKVsBGqTTbD0HjlMVKaIAuVLW2/6NXkHfyOLF0DoO
oPR0rjU8oDZyBcX1qxnNThb5z1nosVTU1CD+k19es0upaDLZN4RHJCe2Fgsf
UGQcJGEmU2cANb2BZMm5+SG8+nQBKYmJKfSEu64HYfr7PBEYVuv48lRRyJLF
IpxR2WWtikoKSldVYwBsJpi2Sm/K/H0Ma4ajrKIlTpN0yVOFqQN/1R5znSmm
bcoXfO8BpBq/vchRgqZb64vlXA1tIE75R4HbYPe1quHWJdTgJzvK+6sy/EaR
aAB3qPfU8Z7qQmLmxRTIDpZAhN6HUSKDHB0vxuU3z5bLyPrmbWqvzNL6ek4z
l8YRwzIrL/is6//Dm2Rg2Z89Ek6idZRbyEfu6D+NSAJmDpLMbeGvnhBtZ+uK
FjqXsnQ5Yc7QuUupe/w8D8rEXguvxNJQ8MHmj1BEjIaLQdW701CtKxrP5Q6M
+p93iG2SXT0UY4cWYfMFt670A0503++5ZjNEUtjNLT20PUFk6H0LNciE2lPd
0XdqDBtvO/HVnAluKvqZLOplYawMnoI7N4kiOHlDzllEP/6alJG+4MuK0i9a
NYyq37+JxcjZS9NjLiDTTMuDQ0jMgwSqK4TC1Op1pGRL2K6FBXsxok9dlxqI
GWpiQb/FH8+4uOM8KmJg58oCYZSByrTCgCNYmfutZPVkpaoqKeM+/ojDDKyV
6rbhmXklcgS0F64mW+rJvu1Jq3UHVWvQS/bJ9+YgBypgW6H1h0uzaH+AGmgU
QjFMdIwRF+GC+Tut1ivK667L9zAf8WXEEcfwHAtzwmio08zJ81WAGxEQfyq7
bxZWfQqQLup2llRsoF3dgSaqHXnggD8jfe1sS+n3bTym18T6oM7N6qxzQ90m
o2N8RVEWwHYVrtDJFlGjMnsMLN7e2/GPQMYYIkUAhWYOZ9iZEs7PKCd70awS
stUL06AZhlYEuZP1IsGciyrUaTRatRzUCsmFU+9/Hcr9MsoAjuG/w9QevCE5
GzuQ4oI6rK9PCARK3rxhkNfNOEQD57U0mhmhnHAGHPSwP54Tn0mHF2ioC3qe
X7/1rUyL2zwdXezjNblkjaUzmdCG/zyobfF7Yu9MfMxEpn/IwF2FdR1PfIrg
RdHttkKVZhwWTRD3ZNC/rnlX/WiQF7vrLVawGeXbIwruhaL7mfOoFHcYvJ0m
ItyuDqhQ2rMLdZHBtoMi8/xp49mM7vgS8mQIojEgN6ozkJKwufdOjALIwakG
ho0WDA1hOBEi6jgWvDQmiagkAzv2GiDukrYiLpv/kVAFQ6zhbrUbOPNq/HS8
b6Wpeg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1IIuOF5jMNd5R6sZskpgPd4bGgwz4JRENi2BSRJSkX+osrh41KxwHwB6IMMBhIk9ECT4Nyff3viGFTrSj9s5u5uYynj2aggAyweQ4HU1q0uhHLVUNksVMwksBPd/dMfWUoEch00ljsWfXG2g/KjEhpQDfVapFz6lfwMW9xMSXGM+RIVdKXVWpU84T5+h1mEIHXH+bFDu+IQp3CHIzWH275CWnVuiE03Jivz7gygSdPXz097MjjR5mUtiYsQ0wd4S6OSOLevQEmPRr5wE9RtITtvi4v5tBKArjUy16v3lflzJlhXd//6/qqrhyPi/1LnHf/YHYM8lIxFwYPnMnAOsAPNpjiNfb4EAfZAM3+BOsu3mCOQaHqwDTg7oqy4X54MiBrDcPex6MfPQ+m2dcdHRWZhEjPp1iXYlhtjBKP5ciFeqozD+7x7j1rFnTodC45h4frI1msBp0/TLR7TNmiPadtgkX260zIhO6w2ndZSeoojQdUAarejv6GJSA6yfNzi02qpoHVTm2KlPIh+5Fn3fXFVru+Q/pa0SpRyJ5lMnVH6gSvVbOjW7cNwIRZBRqA5r/aY/W+i4DPnNaquLmzJKddVL8iZrzZgDzzPaMpr3ABXGUWyX8vqS/p0JDfLy8OStC1ArOPWa8DmOdO44FI7yQ4ld7sruQO1FP9GYNwcAF6zOmk78evRe6pW1nx5Dm4b/RJFfYnyplz86Gr1DkEDA1AkIeZTLf4BuQYNkfm9lZZQb4y/7VOkzQn3+rip/hsqCm5Ks5/KgHWmiKIGb1AvInAk"
`endif