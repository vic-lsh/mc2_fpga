// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jv9vOqT4rvjhgd7pt+C8hWOlSh3PpojN3CjBORrcDAxz5vRTV1J4kMxK0j7o
xwm2EJbvx60AlXL1GSWmPa8nCJcYRPKn93MEkgBvy8hGKm7GqX6jNpwr+690
LvXK7xc600lePhgk4iIdNl1MKHAbZqhfaD2u5pjbXVrNfUph96U2isKZwroo
hjU/wXjrClk6vy7r/uhmaFCVi1sunW2G7FxiAH5KCwa/t5+eJsnoe3IIemny
nxXR+uFrKE9BmVgvrYd4POaCDdw5tGNXQwHDvVtSkFVKZwm8NzQ1Ffm/qy9r
Qdf++NE8yPJQKA8Ng5ByWI6cjWbuH/iwtEDIJZ9qwQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oHjGZOq/NDYp7rh8X5L7/VLgs+YjFLamsHlbc0VyO6BjOUtzZnx0lLwnuKX0
Nqduaq6fTBnFyknaRUlTeE9em9QfDDKJZiQG6W0/AkExbNcFEliERjNnyrjf
v83OFZvVW1GwgY6d78nnB+JyOhuVK/kVr7be6AWZZoyaMrjXk/w76sZZwY9p
A0s7dis0yLVKJvjJ/n8KlP6X5jor+PRcQwH5Vg1/DRee0BTXLUiTeii5fi8r
/arKIMehFz1bCO0FYSB9AzeV5nHYOqTQHQb2f0lo5yMVF8cdfDxrnexo3snt
GfhUQZg8+IgUj65cri2yxLiEytpmlpKi4qavEv+Kkg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IFR4ScXqJxzso4qF8/hLryGgI6/IMxuf6ipSJt7aFXV3q9V9chREYszZt+sR
1BP7MSqsN3CRdO74eWjrl2LdPdYdYNkThWDnYRWxX62BQkZA9PfXM4TcWhC8
BncGhL++Ex6MfqNNwJsPujDen0HZXw2DeG5D+ChX+osZWNCarFCc9iBq2Vwd
7ro7sFmKBYPY60bP2VW5f/RnWW+/wyEZQpb2JEyzaa9R6aqMr+/OouewA7t4
ab3KMZpLdlY9I0npWP59EHbQ+s3T+nUL+Rej1NfwS7vAe2SG8vPYG4UL1yzk
76O2Joq8cW/QdD8H7aO8mbDO6UV/dwc9kkS8o+YhHQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Vd9OHbQ/S3WeSHnl8ViwltN1pyIy/cIO1r2Stb+aOmRSdTbBJhb4RifVH2eL
MgDEiDjzgNjib96aGEH/UU793OYbL2Ok5HXQ5yFlBWTdYnUMiZP+hPWZ+cTs
TbCYjSZ/boISIdk5icx6jFS+HUkpHgVXvRI63oGuE4zdSGwSKvPtzYwcdqTY
zioLcAD8T6FO7TOn0prR7y6UcBYqXFgqlY4QSmGNDSMcS7zC5NN91t7heH81
De62iiv4VAWsdCHkkvhFq9ZDBaC3ST1k6sSzCpADxDHgMvHwOzrPUwN7wlDX
k5Nzriprs3uMPXMyMUC0G9iiu/k/2mNUjRLjm0redA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eBwkzixkBfbCjikJRExK5oBFoKDvCy7iQuSU4jGIeUGJO/EJQjKwoIL+WNgE
XQF+n99kiCbYJ/SU2la4fPkswBcijNV+UykU2Bao/eJhsrhX0KKmtfIFE1io
U70VhSIMKQBuwtkKIat6UsOsleBCoS5PMd+uPbwR2bKgTXWtXy0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
l4C4T5p3niiLZkRWto6jE42AC5/AUqeqYS+eEa0EMDdlRUIqDmWPU6XrnJTn
8QffKZ8dPtmkvncRe1B8lKoQeRsnGI6n7jnRju+ZAA84xeAiU/SN5o5hcfwT
GgrsaMG5KMlsxzSyBVrEGqQBDquqmPWASiEhTv+P0w0sjS7mzRSt5NMxbMGm
C4D6N7r07U9/3PRLdj/zzvowU2aLfbUHzoSYfwrQ/YmLsU/qGVbA8NKmRp8/
tOFFIh4uuiFEJiYXQrIYp8eMeSxL276ZpalGy8QoT/uaoHSzAk4HTO5kgrNw
WsiTOGHMN1BpvUaRD5ftW+6luzEP48LvTF7cedTBTRc8ib26DSM84DMX1eXN
DOaA28F6EFV2OoqGW4HqkKy/ohn8TBE0+QYFH4jJIN5NUvhoNCITH9xvdSyh
6Y2eNH9b4l89feN0QBT2blR7/NQ60XTktwqQo9eMR59jM0o+EKWkanKuPkWi
pDpUMDSWdzJzyq5YOUPa47oVCHkkCUZn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mmqOAjHXR9yLfar7Qc9OTc5g+OMfGmAoDLWL3AUvLXWHEbwHZYzhfmctYlPi
LhnFYHoJ12qvgCiNzj5JlkUvCuVM2YjOGt8j0XyVm9/xlOfLibSnfN5VUokQ
uhxVSr6nbdLiKNlf36bL+Nm429cAjhRUPrq1b0x/mTedlmCNQQw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CqsI/g8ik/ZnDKxrtDGtqRsx9U/YZ9kPsd0LtggmwDzbqThg+Id/4bQzTf1N
UGW49IJKrAS/lp3UjKXjzL2MErHPHpVOBMggqVY4JWThJT3L+8dG4MHsS1LS
VUhQEhQHp3oqF5NI8coHQzrzHKyzXpvJM0+xVgmJJlEIy0KTeFw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 166432)
`pragma protect data_block
pnUmUX+sLpnUg9mtI2tz5AEt/zrzdt9nm3+Hqom9xABwtHxwbvjDX+X9xo/k
yrInmk7Wt6L5UVA8LKx3q8xXdzPxjEhWvMzgaU+GBAIsP5xgxexEnHZSSiFP
K5SIyf27p7mHQSYXfGGZoPjvF0cVU9Tu+mWc1PvHwKBaf21RxSDPVCLudw/r
fDttRm9rNquvUWQ0gBFm4IHtVCGitH/R9Qa1Ewi/7YM8IvXie1qEXrlgzMo2
JcK13WUkB9eiNXI4tHwovewcNRzmpAFa4pOKKxzbnhuSAeYKQCfYM5d9sOsp
w1Y8NN3v0hY9pzDuBFqq5gQZi6Vym1dD6MvGmCgA8k8hXbUzTXdZgz8yMWYl
pMSK2IKWhgMQ5pj789tTJg6d9f/uIziiV4/7hbgOgfIaXhTBKaoYbqf81nNd
aWV+VboMUJ/2gsdDnS9W47bBI50IKlA27V0Nm6AUnnTbVWEuds/8jIKN+w2A
9UpHpUJGIHQWYohtDpPwCHilQ7H3WPLVb/4JPHJygvBxxtnFGR47QKjFuTG8
kzMqaTUUq5NuTr0jA/L2rEc7emd3U+4eWedF19MqjQeaof8TDbkk/5Jdr16C
iRmjnI2FXyN5c3I60jzywsZ9pVToIMRLHra3oruS1Wb32PMQxKAXDxONF5Ah
jsLHD9MmmJh/D0E6P0cuJDPhAxa985+dG3UAMP1KSMkg/n8XpiJNVuEvtv6G
gjPiunfQmVwlofd9bGZoz0Rh7fken2TmFMaeevkVVZoAgGyO7uAzjWiHDQsx
7OoXVxP5cR7JFhtC/TPeo0Jxr3geDja7eM7wHbosDdKhGLkocHlL5aSYEN4W
95FcgLw/86AA48HEX5uOuhLEotobeWs+K5DGScuGErT5JGC8j7/7V1TGRMiH
T18jDWD5JBg7Np3MTZRBwTEFVMGsFrJd9VSQYtRpyaAam4oZGXsTOxVcNH1h
pA0d6kk4NkKt6uRSIm1zf+kqfMPj9VIaoJ3azNLZDU5cFTGoBG++vNmEW8yJ
4pXbM3Um/0WxTuY7ygvOZkUQkL89rXUb6VoDwdCKHEUDyAze5Q9hFnfng3FY
kBfzQzuF+Iaoe7AQrnZCi+4h9k2EvcC/avj7ac0N2wv66/0CmJykNM/KYPk5
UvHv5C4LB8E8Kw9U4nId5kcsTO5vcJuWqusx+ZUpUxMT0LkGo8d1nImJkcB4
6KOPG5CIFCgyKE/TS1ez7XieiyErTJiIvteB36tfX16T4F0IKl5WSW9SE7GZ
Sguv67Eaode7aiZWrgK2dqXwnwWuYdR+0RpSBc09VNk02SU1MLS7IdMYueyU
aB++/QZsX0YifDWIJf/9+7/B57l9hRLLy2X7UeEnL+rht8kVWfDgduTPglz9
diV5YOA4rkbPbc9euTv9wSnHVxU/ynx/H7P0YU0cjbC8yZzjApxFPoUc33Cf
uZPr9LnLCx3MIHNosT3OLYpOVVrDbSybCv4ucdF1XFCpyU6tdpxJ+N2Bbk9L
PWgW/uhq3paiWpbE3/xkRqU3H/lK3vb/671bt4o3yDerGh2sQJ/R4/2BaQjI
QHoEUUBU3oMpMU6y/XOshH3+o8jLSMo4xkjg6+nUoJRNBC2GZS/8q3vHfDzN
3WvleMrnUYJxycreIp1YTE1uglHADyqctoaUCzW6JMvMBCQ7KUdsZrk9D2bQ
9bplS8OroTFM5wUAPQ1cqMEA944zko45levFJqQ4iZ5fJPc8SjTuhYjgUn3G
9jOso8hw+9URsNcMOg48i4QlJmIOzYWcAyQ++7UPFkXsM0/AjTnC8kusUjtp
oE0GXm8cTqK3e+K6A7BcWv5s3qxFqLMXH/sBClOE2/2+O2fPtIKe8PoaPAKp
sTYDeW6nq0C+PVHqajRjiP6yahMJe2FgHQvhm+md8bwsKeShMtMgdLiU8fSm
sZgu27herNYt5zSoMx5a2O3I2DIQEOdUkDQZn7tI5f71L8A+XxkvgjzJyycO
HUjV6+OCB0eM/XRjTjWT9uAq54QpggKvh1ZAk4KL4ytQPPby1KtzH4XmonXV
2XT28PU4BxVh1SQWwVElOAYT4K6ma8Y2DdpoXJlvoGBnQnEP/WONrNGHp1Wx
sq+dLtn2Uv5Guy7Z80hk8wkfMaNZ2kV67ibLDkIORNkDgWGYVmK/fysZ1Owl
SP6R6lwlWq883KeuaAGT1FGqLBmjhxBKn0PsZKJpdpRS3Diz2y4LfHkN4592
CHUlNb9qfoB2dy12Em1vAUi/AVVlfC4RoVczD1snmh88l41p+JBlgIOgGF2i
UIC+0zfGZrNtVcZcqZnojq1pvBr3K58GL85AJdyPciwpt3GNzESNY1KI1sED
tLn0KlAw2FowO9hwL+o95SQssQ2W91o8uBGlJEZjHCpADXKf4qxfKX3wYGyU
6R5/NL1XHf9PlL0dBSbuSFAnCVeHNxdOZn6KUYrcuUi2G7aZmiSac2X8x6wx
WzMrNutGViI6N0DWqyUltFkhDPF3kJdDk476FrExwpHTiPcwwKmcdEiKxUlE
RR5gT8iBto0LpMt2bIoStQHBRJX1e/cER8Kg9V9O7hoJgEvsWg1hAUgpEmog
LpmyAcuB3y5PYgJUZkozpG+T49MfyUUF0Eczbkz24+oI9HLEfLjwh0F4pZ8T
smndWuZOhzDk/EYEZ/iJ/KG55u8bequWqAuhI9O1cSOUFLOgqVdkjJ7TyL/L
s+kqfqe9Ci29C0xHqvfdAHHtqj87Ba5jGgFxAbEOBM2Sn6qRgO6zodLF20Vu
3IPBv9hgYjL3HbHDppZzb8JdUBzXBDNmvbBqR0LKkmo8B+6xyxR+Gu3N3tmy
WcLPdmKcGv2uaWQ3n+W0paiqEtpy3RfjGEWBFJOMQIlnmWYJHVrBDrdSrhSs
nvlmupkLbjzbO9fovfKJzvVaWhVzfBD4n4wPSzFydwp2AcpXxqv/SE2tB0HJ
Kf3lJkTmLpql7WCIK8miG43ZDJyxu6hH8M35Eb0JqRgId5QYZkQJIGVx7O9d
Fa1v3wAxXQKPfAAaT+H7Roi8rwgoDrlN8nbKOv4hrXwLo/y4tO+6vV4pt34s
irOFdFm1dQwfJaJyOy63x9L9NvKM2ynrlGBOxsoppI7NOTF5H759UNRGSA2F
Sfm4uwCjo8FQqqMBk74pLC4xxzzWH5WKl2CAdiKIaFmqD2uKRcT6GLHNlk2Z
K3hjcW3kP9qk3wM+5XGk7US8kgxw0Fk3bO58sCRMlmyrksI9RjiuturgJ3eq
er+yHyOFIz3TF93DRNHEkUNjAcWDhuMYXiCU8PFQ1YbuaFELjkph5COAaWVc
UVL0ghaCyDPmy0A/UkzvSlh6J/8jw1drlzsQ6HDwwaHm9375MlljU5EOWhdS
ACOkZl6pq1IkJfQxNRhxHwNXmcaHgnrqhPBVl4fQmHdZ6f4XJczGm5Ed3Las
1LGJnLnn+ZIkgV3t8GeCa0Re7VRNeKC/FwG7cB0IWlXd39m7x6qiPdCwJWPj
0WnjX8FrYSuHdnQ6tdo+kQkIHCQ0fC3XbKwRztEzny9Xf89B5hwP+h0ppuq7
fMtwBXyoV/yIN29ygBp4ZiVa3zHWORzGSyBqf9x0myrJF68nbi5sY6fvVRvc
ANkzwSvXpW6i25feZKGs4/6PevjE6spatWim2Uq4GatdnYQcH/U3rvmY3WRg
HN1aUIqOdvFN/tCHwQM5DoUO43Ms3y1cVg76miTJ2830MWJ/7bzwoJ/4jnwn
8jCshMhp3x7L4+1MF4GZpd8nnX9uF+95uFjMAYpZPuqAj4ZlfS+oZNRKFuvp
ohenmO0cJc0GXCF/cO9lDY7HpJl7QMXNMtXj1sbTNoxK8d/skmOXhhXbj4fv
XHxsZrfyw3AAwURFx3IvqA9euSFLTG04sdSPqiSwtWTtFbkEHo74xpVjgzph
s/oQI8Aeo/j9gebXht+DI0Ok5E6EOD+/kfhi+qCdvSoirXgnzalJcYommMQn
Zya8tBXHeXBqbX6O82Oj/eW7wnvLP0LQzFDsDrlxgPyUJFrJEfyBN8x/cvtZ
4Klxsd45Kz9MF3P/jN1FrKzqzlG0ib/TV8MIUz8xWdritJyC0OezlTPvoSvy
zN3kWUyCxF53CP0hWp4Nuhv/Wc/C546qC/oKifX7mh61j9Vh/GpL39unI6Gl
B7E7urzNQXd6xvZjrytXdIx+asaKnInMJRm0kQFm0LzC1X4dw/ru636HPisc
DoBsKiTM+lGU8PzA0lQfjuVqFS6l7jMeZUiNtkH0mbTGw7uy1Is+Fbc61ASw
uqs8HRGNpEfHHpcmbqIyTq8wNwFKvKqempwdqLnhY9TqkHH/79CgYDDoPlaF
dqMgh3n3d1+p4NUg74wRwum5tbwynhxyVzlOZWVETJxYpc+kCfssJ14HAGD7
775Q9K3dJ5yhw72IcoTkTU4LPnH2Jox06v11ZCKWiX+Z5HSJPyTV6N6EGcyW
lqkCSGILy+x/n+hBvBtqy0DnMQ6uRTVtjeG/JynVxJEzu26Y15y+gGfgOqrK
3X/R/ZYnYcSbLT+2IDqoC+XQvi9tc/mp8sgZxjnO7cRuoklTVL79J6Vev/0Z
P/Vk6UhayNvU9eCbf77+6uSvaeWB5C/K9t1iQ7vaiLqdhF1b+LXMeCPQnZYp
VNfUr5dj8j2eBoCUBHUZMtR3/pZQkbrRJLpkJc7ulVJqRRz4H2DTowZBEci3
m5WbfSyTTl7o0M5D6cNNUu+xvNySzziYJBduOUjwBFvU2cqABMJOB+LTfb4e
lAr6WRxPo1ARTr+uiZZUNAf6WHiTdYL3ocw8Gxnm39dVgQfKMIo9XzcpgCK8
BARil4WxALco9b9d891M9lJ93Ogu7t6AGz3xI9pCOQ+jwaB4uWp0bmZUz0NK
65OEZKijKo3Qd4ZxzOL0bcWywINeYUsJsjtmtL8yv6YySzvCSzC50TVgs23A
RqxG4y/AeoLTNYwM0Yvsagjra0o0SVCkSdEWUeQBeSe+hEe0c2nyy7c5iVhY
SLfb1T0RW0hhjnbzs8X/Gs2zUmOc61DII0OS9TxlCZryD0TBB1gX6fxPf1Q3
8wEBlAQB85QwRgG4IFChvMsPzSZKq2JhObd7JyPbG6PyGu0swV8btKHSomfF
9ROTrJphPOmBJ/MTQ2Wzx2re+Qht/OAi3HDm8XurkEsq+9rpNfl39yLC3QT0
+x7/lpmWGee+DSROzNH3Ev/APBRc3rMS2tjAVcRhV8L7gHCIihuOQwiKgojZ
Kg3lU5SkljufrP3+v4ZX9W42BXdI5TPdA984xpnJk6lQumrIDmMjcCRkR8rY
uK7UJyTGmU2y3ozS50ZU4j1QZue1z+goL6+mLtwxIH3dupISQNCViKpV+jJ2
1sWUzy6uQaeuys5AFnzjNsw1f5uoSwk6SNrwcLvrUiNwpPegAVpdKFnWg3ll
e5r9s5UXUewscaB3lCMgAICO9knEH7SsW1AY+EaI61CKd6Gfb9Qpj41Fh/yi
PdGmvcH+YnkGRZ2/FLGbA/ddCG03fdzb8rWJ8KWh3GtgvmfCzwWvBc4yM+OR
hGkrJ0a3ZfDadr9uY+9InLkjyNH5eZAZYxsOgudoHq7WT+B78Bmf8PzwSiv/
P7mvMB7k+Jfg4xDJBZsJL+TvH70RNdlZmOBpts3aiC49BInu7HapXL5KM4Y7
Jgf83xB7upr5iSimGpWc2XuRbwaLmbyFdXrvoM0mBlW78vBG07C0VePCWKmM
UiF4ILV2vOm9ZRJrOzeUAlm4yXbWHCo+/rxmxBc8UNykwIOrQuqwOlH5Xbqj
Xc7gvV1HncIFNw9Xyj1U1PGYfV7wXc/XbGTJR+MRWbDM+Wu9ETF1M4LP0e16
S1tzr6Lj+DcGloEjPjRdOCa6e3cIVzlfuitslcTpspc16tziX+PbPk8zuNuK
Kgpjg9h6yuX18vpMitKzsudwh3Xx+7FxuG5iWehL3L9MPgYUPLGEc7njJM3v
K/bMigDqnif3IPei6mAvKzQyUsgRUqM1eVl8EPMxKfrVg2YXHelx64DSsW+H
P1kyq5m70ZJK/g+iSbw9rMqXwwCnjs7AHMqJfivYKADNmxBwpU2dkhvAh3/L
/esYZQStgsN2ca1pwSFrI7euRvJvcWojdq5UMOdSKq1KM79B5QenO0nstujj
vmcKKuhbTLJd4RaU4wk6lszCSXOVVIzoue0hQHjIqTaRqUBqs2YCBxNxG28Z
FNFL6+EGpZeCX3Il3r2gzTS3BgEGb9ZahwLhn2/wDW1y/9Jpx7ZR8v4aXSZ2
EQeEAPazW/5zjhxQNp9H9EzhmLXf/aM9jHlyYV/vouVEHrXQcm19ABPlUV05
56erT9+AAB/Wh3sgx6p9QoyPgH6xM6oH1tQwRyc/VAfFpwGphZR/kVEy9XP1
Mw5x6qCMutHewPD3OOB/iH2IwZjZ1OumNiKvE4G7eARFx8/meDDx9trP3EVy
/TTsNXsua92njpqgvyMNNF7xwGrXaWnOTy/gAGRETmtgDxC0OD+UlZO7YjWW
XyD04VbvM14O/ynL2wwijtbq+wAxF9nZhee8YBkiWOmd1UuTDRBC5/uQNJ5V
M0Wuo3FRe6x3NSP3bsUQIuwCh3cdaGvl+cHrpGjUYmAfT2QvJmctRCuVWmHK
gZA9x28S6qIiMEpkmKsqN3xUcf+e08Dov1C+WT8SCWeNuuoOlP7yrIKPQPBG
KozbdruME6IIbv2tgRmChaPjuxcIGRVZ1Eoylx0Ps/tYq9mxF1p7S1zkdERx
WEbMPxYg1QH9NblvFOZ3fo33mR6xoN5IrXgloCBAUSHpm4tl0ocXrDL3fbkO
U28b+88zsefPQz1jez2a1bnGgdXbeTexxoenaEgsxz9g0YujmxSI9lKk10h/
cVmsEPbONyyGGD4yo0JCPbc+YDSt0ikLE0LXH912pdVINYlub6GS/xkPY0lP
dtnzVP+0kdFyxhVmXxD0I+LDYieqNzQ4BjYb02LinWr5bUD8X4iCQBdfJG8X
04rqHvGOVWJGOrvveFW9VVvJzT+jrI1afwtbpW5R09TnFVq+zRTGjO05E/bt
K+NitqjoX6pO3fO6reeANsnTELHAqRqCd8ViOQG6TwSavAE8dwnYk1XIdiN/
+2fDVMn49TJv4Ncrb05j7gNhM8ghdbFsaAlIT2YDY4Yx0h18g5BtKhHLF8zK
56dVtcAfaea3bUKpZiqfwecgXyn1tX+/eLm9WtJRfaSUKqsV2GRUk2VRQAHp
HssKLDhfY4sIqKbPNRrDMA+ZXhGJFdp/Rfu/eNifaJCGB9boVGFu3Ft+eEpu
ErAV8SrdfG0swzr1qGPFDyvTUl2XQBnVVvjX4XsoIqv595oNS+qxouGyzS8T
ugstiE1E7PutpxoC32kEml+bg44rMET0bRHCCY89CyZWskvIF+Y/QO8mrrV4
lW/JrbquQvsbottWtekjJnO4oykJ9H4MBpSO27RbKeVC54Mh79RrWhplAML1
XQdwnYh7nDQ80xEVwtmSaz2B4grfL5jQX9eM2KMFq4bIZvoQ7cjYHo2WZz7J
7mUibElA5cGyXuYbJhN+JdE/RFaapcMTjJx8/BR3PkCfY+QR42NhkEclC5h4
evYqFuJ6vY28YsVbqjdlbPEMj3/CY4T32PR9QD6Uqo2zj5TvzN1Up1znOJyA
HDcWNqxpiI25eCEOpm7KeIa+WgKr5fcIVz5m2pTbt8txvpPOiH0vFX1mOoL6
bzldjUyb0UgQSCG+FmqWWVZ++Mb8sgBYmMxm2qAArtJfmYsCD7pFAWzDRnIP
gvYdUsRO7ONlB8PSNY+GR1v5aGe5Da5cYV0OrKQpoecJ50Hi6qE7UhdnX1PV
35U5zLHhMaXTqHMaMPrm6BLhc4yYVnYlF1ncOEtFuAS1WaYQimbflWv6QmkM
CDUg3wehfQg8zawDvOmJxnFhrBT1WhffpG4wKRID01jstqcpIZQwcos0sSMT
DZXt+ZjvWUYxfBo9BcAJLU6qbk6zNXjUDwzlp1OE4Od7zx/c1hpBTEeJ+Xla
LpBvdMJKWgoQrbDUrv3B6IQOfw3B6Jb73kHTskzLUumz5S5idEhDYA9o/0O9
UJCkdxnGqMdAIiCfNHNo5gC7JqCs/6xoHkCEjbMk8BV6fdn7ZCwo0sM8VQro
fbq4Vc5ukaCfBn4YpCpj0NwVq+ZDFxCQ9vtWEz+pBR7qXbN3PJsKBZ7Hpi9v
/n1EIH56Ibrp2lpvBb9HpHI+PihpjNdv0AL9J0LjGLgni1ntLaZDhUkX98n0
qZer1FqjvR8y2WsZcGuWQRw54a6MAqeczSQJKCZqX7f7iRpDzxYxWCzq9tGI
kyDOk8e7hpM+XY2HjGJVtT4xbisHhMA2y3IrcSq7hTJjQNpjAVIfmF280m19
Oe0WB6re6ARN4RePQz5J11tCmHgGzxtTAE39O3Zu85tvMppg8xuLew5AqTM1
fLa8V+spf400jzP115QvvUlOJ2uar8v15WyNjVrO/OnqAm+KXkEs/WqeKHk/
FJhjycSuDmN6Yr+HjOiNNtiw144pEKzF0SuMMTW71YQDfxgAoeyLWxQ0u15U
wbIsDfHbSK7KfvnyTAAbbJUuHACcympCwLDEYS1Cdi3GV4Nrfkm3NpqlyvKU
n3nmvZa7F6u+4T3RgpOwAk0huA9oRJXQjKQodNAdJBqVaYB9XE78PFv9jdFz
K/js/6mqbA1H6wzRXqr4q5W7O1EZgbgoD261KrIupsKG26sLXlE2vBpKvEj4
vl2+X8moqgyYy+fUdvQx+8WyR8tCq7CdgACZDO79WNkbNTb8KXnAFz2Csd3V
off2SP5YNFUKkcipJ4skdUo6HXpOlPRt2SUXxf/9suXBlLi7miguhQ0CWrHj
JQ+dwjAG2AzQqXnohWokg8qz148BJAdr3pr8BcBjgiDTK3eBp62ACMkGvgg7
PBUwQTPcylpge0CuzIdtEy3EE2D2dLJc0ZvDB8vPFSDYmGQem6WZyeD1AwMV
vYKRgloHQW9cEDghDdRsFBEKX/V65eua1q/sgnQwdZMUk3SaUIjflRyG4kt+
LdOuUc/xHEHMNNS0kSGuQeDDyHvF5Qo9QX/L29vGQiUrvyKpTzJ5pfgJ3sAn
4uUeICTWyguM5ruu2C3h2ACKYwKnTHCwy13O9LxkD220nv02Y1hgsCKvXFDD
6xSVe613IsOLodTQWadHLznZakxdXP6bN2GKdevefPcF8bsDhcnele8LtCds
T3KK6Kr790lbIpZxjU4Oxx5pkHYyxWOTtHr2EybVoqXdraiegcKoCBKEmeN1
oyVujvtSTygitwVw98x2Tmgl9LXaMa4dS72SQO9YkyrTzeBtUO58h6mU431F
IXQSIAFR5umVjTCip67HUhyDgrRelrjsm9/lZbUmatp7RvZYfP7IrhmZ7g80
34oNScqfQsFAKxoNWDprO4Jx8SUGo4mF9BDGmcfpx9wSfHz+2T0werT1GY3k
JQaMm9xdon1/7FeILrqwzkTTakvL4edsctasWKuaT+43vSiaEFcVnItXWE+w
gTnQ+gDkyuevE8GPwMoEA9+/fGZb+O/8Oo2PqT4gkoGNOEUHxgOEhRA+B2FA
+Gqb1BMb9Kh6GRcAucrNCklqwNP4a7+SZfkeyNT0bshMdpuAUssD8sKqZith
za02kbX5Wi20csp2e3Gf+ZtDtkOruRKRUIjthfyefyX/l2uBbG5WPv+dwGh9
anvRNYpW+1ON99zY3pIYfKqrlanfS5M59Xb9PrlDckGo89I9tWNsHHyHldy/
fOmVKY+dLnas14F8470SMxV2w3TWJ2D8fkdnxed91HLU6nfXneb5vShaRmtt
b1fcG2gMOmYJLcFODjtbNmxc3uFdYDo6kiSQ0u7Wd/zwUHUGVa0jZuNeBo/T
qZrBfiuO1arLRdPzJaRoNh/IUhprEUMJz7XMQ6rHfal1kUhS6BKTuggGTHvo
ggUTYH7kMssv4Gl+LWA6KjNMPYSTzl15OvSsgtBJM9C7p4RADODCDRMAChik
m0Nc4U0Hhp1x8v3zdIMiU0M+mR3IjUXl9F3+tVQQQa0wWlLPHz1HSTBunyih
SB5DbnnpJieU7rfS47AFXj0nx0x7bD/rjiEtMIL0Bbg7acUFs3zEg98bm39C
fPOxry8G/HhY8l7R66PPkC1u4ni7a/UjoAfMfjRP7zWXYBR5qgBSbikfhDK7
Gj2XJTp7XBBtczX+u/xgsjkvIf/Xzx5XO75wG56u02wqb5tbljj1aTpgBWG7
jW2D86Ro/8mHGR4nShgaAa18NkP+wcQiQlOc6oCLsCmvf1WEo0MB+hTOxE9d
wUR27K2JTlM76O3oiQomTVOAsHE6B+SFa0FVr7dpvtYCvvOfdUdc20MT0umu
aAfNwg3s+1mtPWiZuFsAeHtf39b/+QXgyvLl0NjAyBH/m9DrBdcplmhT+Qcl
DSKhM6znqZEW9RnFu16zbzH1VUB+mx2chEp15ngcri9VGzwBW2/cu86Q61Wf
QhFzfgAQir1yohQzNIz6v0UQ2V+Leenn6getHu3jMFgHqTh+8ouMbF6qKbDb
2L4C63eFc53bs9ID/EdozxzdUEwhRboKTVrzo59TE6y86P7w3Qud+4fJ3XXe
sWgJmKk7dMm4vqbc4GW+0o/RwGsvaymuTmLOoclHk1vuJYW3WjC82PEiTz9g
ctNzN/P7zrNAAkAN7M2xT/ufIx/GrvJR6d7cnUT2ZMoG1pDCMVS26XxRCYQf
JJd40YjnPZAaWFME1k0H0Co0ZSixZ+IUAxLg7GR39wUvzFMNUiDJBTb3jhNS
J+kY9AM4FDVKHyF4WhJPgjLmTDhnbG6s7HjgRNZj3yvR1ybG5ytAb4uh20fR
qqpCtw/Ez2opIF4f0tX7Z9GsJbNh2i1pB0WxaqS8RE7pKJSWyRwPQU1FZH4v
VeS5Ah7avJd/cBtop+ijI19YQ8NWb8FxV3X705kTWtYcNzDjVcSUTV3ybDJL
enN6yZpFM3FndEb/xUezInBsE1maFaJxbqxpff2wxzo6BFu3Tm7Qre6CODw9
EJf1+zjD5iWxeDaqAgbL9Qu9dZFmeVL25/bJD4mudk+zv7/fvgYQCl79qGQH
YnR+9ugrUJI4+aOrgIMa7u9hAHzzfrSwDNVqg1ay8p44HRtiQtTuOH8lTDac
yWIq7TBrHb+858gy18siJ+pcLkRTa5niW/K6NH4pS7aJGIhhLL34u6ZWWpjP
RMyp7S45U22Vpc6UqrCaTxevAhcHq/f/b+uhai5vsKaenztkdUCnhXZk+OcT
qYv6M90fl0KH5cEHW+TVlR8VVTksQprisaady5ULvYZVW7zNPUf/XEYmuvS/
fA8+kJfA4YBJa0l/e50XfuuBvR1QF8Hjjp+Rvq5CCaFJkQjIB4pN6tbFPovF
bi0iTa65S6YD2dIwCVOlWZwLKFp+dKsZVp/ufbCJM0VSgHkyaafk/WgfxcGf
51707/8s1GHPP1wvCuar2M+c9mMVs5uadiELn3T8P7SuCW5JglstISLnjX9b
/FRhbVdpDeSn0k6l+NsLizWFteKkocQXSQHNlXEkiumMUp3ycUNQY4jakQ0W
QZowQfsKvfJ4c5EuxNhf+OgUrq4tCclwZCP/9Fb4d+0yOBE0raHH6qqBJ0PW
rBMCX4HoiR937dMlhfhs7NLw6y3WibKHvhD+NPLk0dsWCL1/fMwGBDJIVas6
TqWPtP3FyOFzfAzi8AEb6wqU8dbwmhNTk7RDXpxY2/YXoRLHY+9mP21u1D8w
pJtE0O9Mc2gQDnWeKlTuuKKYoXRSvV2Px9Pv4h5LA9KHXrNFXrJYzg33Q1Ji
gmWTU9VuSldKhntI1mANsdoHF65JY4WjMJI8Pbl0i5F6Za4gMW/2Q0qBoFFn
4N+QXmBKB/diH/Uk6wjIhAV7P6W4LyYJ2rw9OXbGR0ZXhthe3QRh9YFEgwrB
MJbACK+p1yvqJ1PUBj/eWiBo6XoN06O6WW9fKmOPBCGET/3pddypKFuMplcS
rvg8jsm66PTawnuv9ukPGcUm6Axv47JTpnehe/LNc8Zb3hVRohHhXiTVG8fQ
RTXBdOp+N2QXyWV0Znsk67V5Wz/4CRUDNa/ImKL3SEjEH1cvzk98k/9yo7WA
S5pvuc6Su/qEqj28N9EkfGp2Td7BYlEamNEKhxTlh/b7VvF+W/AapW67TcC2
Q0P3XUOAnUXJoP2Rt8z0J7Ud8q/aRZH1fr+hKyz7BaQCoqvYeQdkCI8U+Kxh
s9FgchnyY2PRb9VTf31pFPyVkkCB5ySRomRVSz8ACrTGPkJ00JH+UnLjF2TD
uMRU6rbzUU8ykhA/w8zW3XJZxh13XbnfmtDRh2+hmcYtUN1pQl2i9Oex2NVZ
X4PMSP9Ca6KnNXrvP2uV9c5aAmjRBzD5ZVRhSP2qCGanHeA2EdbL1732l0Vq
0wkPMmKG3xjEGL6yUp3nQ1sRgIye4Q2SkNCwjEItCNzaJMzNiRt8QdlqJIsX
KYbyDAZ32wfDnnIUSoaJoUS8z+VMIQ+CXTcUo9KUX5lPnyNjLy5qlNujWjPx
fEgUDqwWs6vxg2N5UckvzbOek+ja51ZlllvnxeAHccmwoUdSR2LYpw3efp7j
wEhqg5bGHT09XujVYK7tqNT6/mmGJ/IGEA4O7wZqTpCUk6aXE7qg8dcjQr39
8Xzyq23kCLgblkVnrdtWmDZYYKJTHafjMPi3FkKvTYDOcGvKFtvGhkc54loX
DSrRfLubeLFvrOPJ3TINh0sBqzX3luThWsKXgUmdra4ksCe+EwG67cJIWvxz
lKYcgfe0vtv7lMd7Z9Igv77YEJUizh8KPtlmFGS7Z5RRxxJrcY0rt77C3nj6
04Uv6AVg7dpQ7fQasiYFOKepP0T44KxWeR2D+enbWyjVvgoVlpnDBP8SfTe0
ry7iRysoJ1uouDUtq6nm9O2Du8BqC2D25Jmiir4RlVMjx+T7JYtt9AdXhRBT
xGtCkT3cvww9tArlSmAfYvx47foAl6J6XbNYYTrnIDTAnlTkBbqtNyDSVF/A
H71CRPcaD9SzjGP6JthHHANBScL6VRxh/tqa8kySKCC594+joVhmMCxljKqR
x/No5HF8NhPUeBFOyJyq00QY8QlYVyE9Qk4SOkNXaJ2RcVX7uaizX4sgqU4J
eUT991OsMLskokoqtDA3YIUFBgebXn+///CEnJRZQR7y/RY+LNtQ6eY91goQ
54bB23s+czJK1Hmo4ECj3S0747pHrLkDQTlPUYvdRjAVRL0qkaMKwQfe8GGo
taP1TYj1khrupqiFXUTT5yLwgQAJ8Ucp45ixZHif162vL8O4HerJJ3BmwI2+
UCKEa8BUuuBa6nRmBxlaEXisVFxikAdRdCw5HcFI0P4+Xnc+wIftgoP+ACjr
S0JcA8i6zG9uRmMahgRPpzb3onBERirLN7lhkdr5Rn+G5lNLn84ErEH53G13
wM7JEovF1y9IrIfanR0NLj70PismJ03PExqGbj6Vm76BR40pKwVyIQaUZ6yP
EqhlXqkdekQRWjzc1GzLC1eW3SIpJORiNc5Ug8TylqnZsYvmAgmRkrCjk+KM
lh20xjx1c1IWqQUa7JfPEICrfWlzX+egCEKWFa2L0QDkdPEPVbLYl87RGFzA
qKvPqs1eFNu6/rauqJ6wnoiEb20Xvg26OI5uXhPBcwIfT7cdiMIL4n97cO0C
jEtCL5jPnutRqfRVJEyQdfUdiMBbgBuJAXWWM/O6AC7SUZ6LgvadBXM5WTfT
WsTf9EWFdClYny5C2eTSn3HAcbpqcVQ5wdtMHSjQ/mvvjX2RYOMUn5uUSppp
14piD9Z1gRdYOLmID0wJPHyz1F/T9QeGnhoJq6FQMd/HmKgerYE9cgVEAerT
OKr2ScxlabKNluoFYGwTKLVJyIUpksDawCPirY/yiZF77/u03vn5rR6SIREp
mTY9q+hOcQgJJIZSBOhAr/hMHVjDC2rrytcIwgdGRp3bofxZg5UO42kGJKHm
/XLsPf8FXsPe9ddd9N0oWGgxzSKzL3t29rrjnzMhc3fUdZgeOZlMJ3O16Yt4
BoQfFl/JIjSvtasUDP+At9Ll3oxvCassJcbPkNlOpDwg1w8ul2Tv5Oq9Lqor
SWSwQKYxR0W29YtNwXUV3VaAgJL0mroxcUalU7feP/VgkMwfEBBvhAX9AwzD
aHORvgSVrwPEami8hisv+S4wUPSfmwDy5AxUdMw4MfvXiRp/KMXCzFmHMu0u
0kyfUuYGuOY7PzGbZS90roXNf+YHB2JNuUUXppIu0xO55Fw0CoucU83yNXJ+
7JeM0R78pHP/Q4whRqM9bHPrk8i4Xkmbqn4uju+UTgxfGvcG3l/K8ksuGuDt
MHfNG4DBFUM0CquhlCRM+JjIfaGdjpfzxOOPftyY7n8ZyryEuWOiv1koplN7
355eCd3a1Go7a9rr1RrEkHjBxSYFX+rXQj7J1+WvvEj7vkIJq1lYy9WGw/Ut
HxmiKaD/jdlx5nPVpc+hVdc0VlEuBIBpyBIur7W10lUpG6/ZQd50sMKbnULR
mo7Dkwr4ZJGQfL75oQHT7WDhjlMAupoQJdM+SvF0mBaFANq49Sw8bBPe7j/r
6+1J5NofqrTzgm944p91DFsBx6ehmJ8VeRlq1ULddTWs0i9VwWIOERUBtXw6
TOROi0woOQtxp9BI2lOK0qzTvvnx6IOnm8TlQQs0QsnJ9a/iI4y02E9ctC0W
ATsKamwSsw/zytcELMeJqzLQhe5Pfm1nrJ8sTPFYglZ+dqup4vxr5t1D1VHf
/WHpuOagENYHIVgdJIzHOYzD2bzoTpSdyKjIOsy967AwnE2mqPV3jBU0EIMr
2osvXpwOIgOXJ61fSbJVuKT0fM/IGuiaA3XPDar7Kka8eYP6llLjabA55Cy/
1T+8xbjpViCIYAqgtOYz3Yk5gHNtxweO3GNpG0KAfUxcv96+P/f0ozPM7xvk
/oqBSsTVBxGy3YVwib3MV/ZyKbr0Kypcve7tEWafWK4dLvrwX/SZz6kUrNjJ
3HPM7GbewsUeUw6Linmr3wGlw7fbf9tckmZIaGpfvIYcnqF0cDox6midopyg
McN+hjIgwSK972f5C9ivm6BNv2LpgKctDy9D7Crww3IsfQxi2Ws9RLBoQ+45
VDm/cO2OpSNXwUEUfZXBn444tHmCMqKtXUAVEv1i3z5igD+hS9Jv86pVV3DF
6Bhlpv74qpRdJmjWRHG8njbouOWfs3isSeKXJKg0XJRVNfAFXWBg7uB/jej1
iJiBPESpvpN2ThH+8ocHXdS8Y/o2VO1YyW4t0MEYtbp/iG/gySptWL2/I70K
vG9m7VN1bo2i2/tsU+M7JD0Rje183ufBOB6Mv5T+/k6o8yq0vpLErzoPY3jA
at6f4hytAtbyS2zZF5ik2WGpsZXGKh5XKqtc8JKVRbZ3ZDCcdl32mvVDRkJ2
A/lX6i7d6xLsnY4qmy50HxEPV76ZZFBpzxBnpHCPvHWUTQEXnUnpRJIdC9ZA
CP2b8VJPtZ3EBq5yegU5CJ5nB2G1zwMDsfTaJ2rrCZvDgUORBBhB1NVmmcKc
eBsLwpfuNggHsSafA+zmcsl2ob/fcGX/HeV+HLTDz9UJUvYBsExkJ5r3PIgH
eWYhJ7LRgZvhTjHw+iMJ4uIkVf2Cp6VirvJQUC0J/D4HYZt2bJYN5pp4hOf0
QfgtyEVgopWZ0tI0KeV4g44M9a7NC5xuDDOShRkIRvCOrDH6MqA582zDoGWs
Zz6qSaqbEM28eN3mHAJaFjMPrpA6GRbDmT/K5Ux/iam+yS6wfu80l2f9lxb6
KlQIUE/PRXBWZeUXVyANQB3zjo5m+chICyHyqwQNLQi4d3PY5NxwtbHUuYMn
Tn+lirr0pBqxyzSS1JNbne6Uv3XcYqkzRXax8avg+jjPR4Eds253VkGMMLUC
u05Zd9Py/mbP+A5M0ToEPAmU9XRHPdQN/ofxQkOGHjM+rP9VMJJQbPPVMp4O
qtVXKMHCm9I2wdvRBA/e+Bg9XA9sTWxevYW+5rLYYhHuQWuPLubX7iKGK5Mf
r8AY43GQg1WmLhr3HSn3cTTSydBGMMzIvwG97Re8Iyu25IBMQm/VyBBRZbF4
0WxFF5qQZND3av7LmU1JcaTquv4fF04vknYkMOPeZepf7XBX7GGn5EdtWR4e
QWJvIyqiiEKynbpLHmZxXkev6LPDic+Nr8yogV3rnWal8XYEQU7jn6Q1E5bq
VMcHTJmWL0/m2U14DjqfWgpTGg9Zr/HR6I0bnVkdfexHIZYcukRmOwGsVMNE
KyRU1dYI52LnG05BKDVHkLIITl1MH8oZDV+4zSyYFnesCXZL2u62xywNvD3T
A0lh5W+d7EVbpfMf2QrCweNkjV4n7+suvmCETynjNzVZyNZOnsWceg/KzOac
xbIXe669rh23akD2VwWYWvEvUm1QO22gwnLYIgZYbgJMi5bGN6ypr409PA4D
TttliQrER2YYvLJXcUurTQZCmf9RvckbLieQK+XUf4zLHo+CbFZQf2nBRGWY
io/oolc2CKvoqgPpBIvMxhkI9oaPNNlMDgING+MZ2hiJ3gBWaOXGlXi+YAwl
tyGxJ6ANLBr5wXFnEQMrR3OVdNoP2RsNB6ictDKd382I12e72ka+z25P9t89
zv2YP+KhAG6WWPAyrDKI5OZ3x52OyaXA3WZzADNqaTOpHMcYbOrZVJFxJiiX
NTErIda66m3oA8kKjzwv2fj7Z8MJxPkYdV/29ggOMkF9cJ+yctvz2CNgOyGc
2CmGtzwP7Wy6WyUZG45qrzIMKMhln/yYDZX1Zd0H9srDIbV+FPHBh7M4SADe
LA/Ky7Fpc3pFO/mk/KlgRyYJPeE4wiWg3cOxBxN4Zzp0MeFljO+r3zeqFnDR
a5IO1Pofop7shHJO3ScsE10tukq7Sh5PtNXz/FzsY71p6hc5TV70ztwV3HHs
MfAahrU5C+XNetxUGOUy98igwLf+KvS2JYHIS6vYy0TMsR29UTVUrnYQN5U1
oHNYRy9t0d3jxeXwRyMv2yhzvsPLk84xlDz6fA6KSUK2rMI+xQX9WuSFTJIV
L3a2T7VNXpILWxFXZ5288ulwRMzfX6eOs6MhkR4LJgHkFCRXQ+AeOJYCkCt5
4/2HCr7Kj7KYexlopcfs2aQHRiuN61f3d1i/b4wsARch1cXR+X3l/zPx9ibT
CyqT4bmE7VHjt9Wch/vGHQ8m7q7J1powZ3EKt8VqKhpxlduxZIPe6eAij5//
M1asM0D3BTNJUw5EerUE1BqOjb5XoP2DBVXQ+H+cmhRUL4c61bWWMI3EXf1W
4g4hLqERWUNmtNACvKmewfIPABIGbsw+Ec9hOLLwtZs/canAnUcAY0wEnUc1
ZZ9w4VbZ/kDodLfk22C/gIDTNF6B6ClN5zm8Ko85Ul8o8y12CSvzrkZl395y
LSo/4qJfnSJXjTHAq/3txpmFrDLxYlgI8H7ZIwfUTfyQrc/Fx5jIgdegV4Lo
c94mh88enWNRlnn1EtvhCMZ9rIKMLrNO8otnI+K+G6YYWLxuMUaA4W1P2lA8
F15oMhMTpHjS+FHWsVO2n+w9eygJqp1oBL+qQlQCHwWKJbAJ/H4PAobuyIkm
UH5niLf4Pcpht9+YEivViPSo1pK7yFTaXmcToyHU/C0fiu/gmCAk9ZQKVjYX
WsAdKe4pN1g2B9gnPJ4sZ8/vejx2ejTb1nEfi/a4V9gFqvu+xlRcvWoDxpDK
rALAkwrUJa9OId7j0LdXZGiJlQWjeMz1z1NTa5PMRjw/q99IpKB6W0idobeX
xDDgdMeRuLMCsomoA3QznF6xEdXBDB/uptohUYjxs49rJFZeAvzqvOqJ1lnV
7LjD5Igpua4yxh5SdzjuALrV3De1GX+APSot4Hqd/PxomAuezYkbIqNfs5KL
SspBB4NsZ8lVN6OqbFqDuc23WSLwwiQrMS4L9DGZRwz/DPwUJjG+cDMyF5yA
MCXrHwUM3QBQ1ckDCCzW83cCmX/ts7r5Aaegm0PvCjki2xgS6qotG3rw6AEj
gaOMAYGMVWrQWeSLq6IeQRF+H4JBPMDQlinQSSc0HtpYgqy0NwUry9uoP30v
8vIQ7jlWUIbx4u/jnEzwfVgVBpXos7YfPQXhvdNxyTixbZdz5iQzgyecmdTT
VIx8PVETRfY+pb/in4zlT1jAZXGkDyxeHper6YAQsHz2xT5F8CwVLTJjlz+5
dNj5J6cplb1HkCTXYqVGHh7TVGUIhNbtTlTC8vf3t5qAh4WE5doXWuaael+H
SbSSPg20hyrnRkSgWYiWIFGwRSlwUN1ueOp5RJ/wLPWR/e7hYMqa9f+35ScZ
GT3WiQlkGuPAW/eDMYR9pxnmlOndG60KOvsUGGu6odrwEcfHcdtkVFVWENmR
X1+r3rHcLT1n3qD95SfNUnaQr2emgIAmcUroQ6W+uN/eBN6dame3Rb6m07C6
zbEUXUSb8WSutcuh2zcOxroTcC95iyfpv9zJeWC1l967vf9OgvFVFa5Krw5u
0kzThjeAKqZGjTURHyIu6+tX0n0l9XbZCtS0eJLr+bXuTd6gY/qZm7+38IMX
JCLcV/unWJYMd115eleToUySJbnEpeafieJeaygo0nu5RPW+gYYzsTupfQqG
GvEIYJatEotKXL3fTCBnT8PPks/LPQBNCS4Usef/LUfVLq3wt+2VqwqFKE0X
lBl03y8FS9V8njTg3zHrzgPT0krEKLdQHevp3LXdfNf1fSADmr7RG5bXrIni
MuNXXO1Wp+3l8rAmoHXRnVSxH+mXsDDxnIy43/Dbmxdg9sXUQV7pMYCG+3fN
vu7QFF7hr8eKhQgjmY9shUgbqb69s06k6kZTT+xk/honlMytCgIIiM2js+Qt
exM6kCeH5B8pfg7eMZDH+ZBYgbcKpKKcPH7Scw9IuPDjy6PInG9fDeZSfKq5
oCSe3seuvDhUuXnM1cYTi4OtzSryJBr/Rj+jICGGaaZ0DCh8f6ih1f8fTNdh
5EPChAmw26TTyATVV4PNR+DUPbC6peZzOO+zuG5cbXV2Nh2mJLyeF30wC/hv
chytAYQjxgfqYK/CikK2/UL3vBCa4NYcHpzy92+nKh4GF6rQcmKIIbkHwbRt
VbE5TMhy4anrA9sB7iAq134MjXp1L6RbJCEoiEuLRWDwr4y4CB+FLPf4ys+t
64I3Ob+ea39x1YaqPUjzdJEvc8jSdcXlPTzJ7dwaxkYBhCgSeohb0sBsHDVp
Kg4cdFkK7GEsrXPXWebwY5KkbZsTE9gk0vK5VXWZWQcIvt3lfLADR7WOZ/j3
7/OOB47BR0DqfypTpSpT3KD+Ww94IHpH6wFUQnKAYOJ36uNTAX3aP0UPJm+L
omcrg46EjqTwoaocX6L0J4piwDgfC6RA0IMQZlO3av3IB25JRqMyADyJ94nu
nWuXEbVOPi3OcdpCOzdQXCjEajIZbfhe/1BaqTC/fN7dgX4s2Ryjd/+gaZd0
7d4OQfFkTjdBpBUonJqTeGeIZBu4QnZM+UxX+6KQJy+jIcdhOD6IIrkQrTQj
EvB2QUfEBwnIn5woSjA8ksYlo3aBroEzKBCitBwqabAsGAsHNBM2iEV19FcJ
dW+b1yEmb3v6NS1cIZl6G/eXwtMuY7iwdv98zYqouguW08DJ0+6cnPjiUyA0
yffWJjaavoiYn6uzZ0iaaTf7N4PlkWx6wdPEgYXekxng2zrvq4Ye9x+Q9yYl
AAMt20wYlX0+WU4UfblLBsiTafnOZER+l4V6YlRfhY5CLl70NQmPEOK3wA+n
zj2sikXTSXglGqvAE0HXeej+rpXaalyffldwFtUh6satEUmRjvNynCujjiA7
wCBOUa65jz4zcW1V5yJZcftshV0zubw2lWRxa1sTGsBG/pEJ0+sBm+q/h6Qw
yDsd5YqaJ9wXGFVWreiKItLzQ/H43ov9S6P7unfDdD9CmRJWmyrxWmhJwK4e
w1u2cD/tN9WgX+3ySnp1zp1omcIuWNMHljDRqrchY8PgUmY6M9qE7qFJRIjG
qEin7ZegRP9xsqcor5cB1Dei4dWHWiBymBItAxuEoF8XNN1OUX+D87bx46OB
JgVngM79zP/fPLtGa+WEdNzNZa1S48DPQBWid5IbQUGFoLWpDazC5GdA+95J
fT7mFPTqyU+w5ke0cL9lsSC9P2Qky59Pv4O9wOEjwZTrrftQLGpyZXpB/wvJ
1vXTiYznIsWIQogwlNCaYYWtCih+aBFLvnTP0Ex4JTX9CBTTNyMH83ttcqdt
BtFNMHAOdD2Gez1sX85uNoBfKdjyKw+iUUA1/J0gqJ+7I8WUkC5BBpGiUeLj
LwG/4FdZjatO+z/CbtgUugpiimjWDV69kW1+FAcE9v+v3sbKhWmshKJxiMkm
slU/OB5J1v5CB/ZoQdSCJv5BKm6shXxg3FixkRaw+FTAzZ8HWNKUUMsEvIFJ
Lgkz+rVhRtl+dfX1qKkkOnQMPo4hRMN5sqlPMXRLr0HIIUf5mKKOIGVNOfLW
OK6PATB/7sszNi+6E2ycYZHMFOias1ynH5c89QvpiLpg8DGVvL7BlyS62iej
F17fGIkCZuXqDnGdkU6PXkqmN72Wc3m+gHsgLl4n5gOux6PnkazjEXLfH9Kl
SPXDRDbl7JcCUv2VtZo2isuKv7XIjBqCcGv/BxUniuFXGOgtgpsUUsAk63/1
KNj9DKvuGlkBV/TGm/uLziCUjqTshZrMMeyoyApmakdqusN8+OfuC4GHavyk
JYm0RRjVfc9qs2m89C3uQdzNIIFzURgCQBSOgqXvb25/d8MvxqSQRZrkZ3EZ
jHPXv6TPpBjn9T7qS7q7P+RbtMcp0uDeEd73yMxrlr8J4ek0oKr3PR/Yd2Ch
tcdhcfGST20DmowX5RWIHp0uikzQ0zKRQJeyGjn9RVlNYw05yWTJ76Eh2l4C
VZXb2ePcoFN24LjrtjKAyLLDZJjv5zHGwC3bVypS7J4Eu3vMYYPV89aYVAcy
DELOmf043wQcsHkzw0hoO66iwdXPm+/5FIlAzOIVoCUFTqDO4XPaulF6JxIK
9wNtfYSWNNjKhbkdXvZIeRypfalCDbERcME3GQyde9ujOoMBuEl39mNFqqfZ
Ic/Qu8A/EXy1ATBiktPrEk1q5GJH6aX9iU4AJo6lg6kfL6WpxKhN0WbHVcI5
ydV+pdxIAJPAwT2I3p788E+NHsoDna5qiLZhB4Sc9+Ho0jIUv/DudZN+MNiY
bVLH0sb0HvkLr6bcXBFs1BkkdQPhTrmo/7GnIexoaHOOrVGSUW4RH77cXj3n
dBNadIZEZb/U2BaokrDFP5i/rKdFGv+/S2rSC914Sdk3APVADikh54v0WwpZ
erXtdKFktHFrpyjwEj0cZb3ikoebfxK7OIPVeCpGmkCuxynfhwjD01l63jfq
GgsTZnSXIfo4NrDepULNsllSXnH8UFRr9ROs6ZDjPF4y6MQq/WL1Lg+vySX5
dNu2aCPOZMBteIrgL2F0MnMFoNr2sZwEnPZwiES40BDey1VUK948TEKgvg9v
7BX7LQ4OA9R9V6rE8XYfocCLm6t5YfmlRSs5/AewfIFrQwNXbePf7/2ax0ig
Sm6MJwCKsjwGD2VtlxzxPqg2oewAA86GFaRNvO3Ita5Fc1fGHf6nZCISNGpg
BuC64v0G8uxnzt2qJbTy42I2EK3KvboHe7aAUtIRkAyPGvlkwO4WnHMegGfH
HsGbKkvKajFWoWadGZTwgLTPcKzE2uJJcXZqO62ciAHajPmckNfpKBGBhF/c
BoC6Ma9M9BwJBFKN05dcJw7q12YMvAmk6vsq3SlWh4VvUIZFinlCKWDXD4yV
lnesCzUEJJ6NLHTTiz4QvqN9tAnK3v5U5TBiuICSA12yo8JGH0seMQL3F68W
O15/yAak3yscTozwlZ8O0DfIigQf+sTr8UBq+343SJXUhuJicvwr/QTS75eE
bj/DzgEdRtwkZqnyJIaaI9foMghK9fEwMGM3xH1Y3yMmg0xLMRe5n/QAnpcs
x4mTdQEITCb/HMk1jzf1IlqimSwxFwqO4OZkBnJlf/Q5ZWTvCNYLGQVWunY8
XYXpzSr/7yGOwYX48wgoiqd0hvUJ+prk8uo2pRLQMWlzI6D4o8ujORNa4HNH
tjZlbjWHdnj+p394FDtPIX/UtGLApnQIO0KgjD3HiuMrYWtfCh+JtC5aDWtZ
OF+Gaxk7Sv5meag7/chRhB+wJP8ux1TWMCgjm4L6nGPbM/euh+MIceIloN8S
ol5NkABvVGeiP0tkQflfXiyB4vGX15jFcrWE4nx/OgHJevjdiVVgMyVkhde3
t3LSSN5CzdxmsSJFqoO7OREq9iAUkSka6n5e+69kOFvznmoohvOOKI+PAqMN
ilrUvEl7ZFNZAhgclwDQRMbQ+ELlZb4WpKbiOnZJvJhnwiSGS+H2vC1nWn7f
RADbCfHD7n5GpFJADSqCJ8819KYFMMmFlSnOLUoJCoGtPJNc9ziuJTBp6WPh
ymQoTExWKYssutEqnWr0O241/OnNi7DSrsAYj894UtLLOicYhijL+XPXv/Tm
GYHEEJMC4h53dUWDeLKOLm12PP/LLQnrM87MfamY1mN5OpZVAj/faWyh96uf
vwC0ceWNmcszMD6GRyMW313GCGfUzeZ3ZZ2FMdcmYRE+F/hKheSBu76cx1Rx
i5z2A5kcRmaxFdwJJ1pRBYJgPwte4fAhDZ/+aVo4AMniKH9vi5zvVhDzVUVZ
AeJ8A+r7Zn2mGeXJZWTAU3pg8twipIxOUIgOlJGkD7e33Yptxr3ZWA76/nOS
Wk+jjeKVGXcKUtF/AQC7IrWGQl4yMntCWPwb4dDbp77muFcZH14vjJmL5UmC
LMze9EU68xB2mxvKcplM5mG7Mm8FDfVcs8TIgh67+1Lmz/uk6wMtWFhsWMVB
XT4o7Dm9k2j5BOFfKYQJs0C+UBeq/J4jk8aOxxg3IjWSQ5y5ohDl6bobKTe2
srrVCen5HhRWruaBc32vvTO3beq86a82bYSt8TcUnh07fJZD/qe2mdUkHqmJ
/glnmgWeLX4c6WiNbZ4MX1lMe5EDE+w6cWTzU4/ew1JRrVKgK/2durLOQPU6
KG+KGeekSlrpfxxc+DCrk1z8VFRrx2dUHE1kDgvfJAJLgR29eT/cC9V6mfbw
KQVbN3AuSRWSjf7Pel45uajPYbMBqfuVQG//tdgg21fPh6acviqWF5xrIYvI
TlFzR/gigd5rQb573Ah+SSnhofzzBm6dPEdKImvMCsr7va14xbI8ZTg3X/HF
dd5IMgiVxUNSzTWenJlhwmHXuw8epQrVajyASzPY3HP9ZZspCisxF7bvVO+g
14RAY+Lb7g8IMtSbDy+GGMlDa+M1TgKeNzEFONH+ggz/Wxvjig+/7YhwUJYy
DxOXZ2BLX6sPyDQcuTiS8yCSOZwbFXEzLad4dt0bDDhagqSxuUdDXGmmezYp
LkkOzhb8J/bV0cYztgU9yFm3BEkutNQ2bm3dbBmwtcbDdvfsIQLQlwKUP+0G
Y0SBnDVxf7h8T+BmV42za2krXHAX2ZWsw/YDUQ8LWak2GYtz7Dm66DKHQj9P
l2KJ3ShF+O24W4t7kBDC7KSBXIvEmNEnas+YQx3fqP6N7dGu3JvbXeBmdq9k
+W4foNyuxKx8On/6mjsfK3irkVwSKU8/jquriinYkteajgORpA6X3YWjiO+4
C1T9uAhTY1/nozBi2pKtsAHZ5OcFBrW+QLCNxtynCFjKW/Y0srSwIycg64+H
VBuGHvZhGAJWVJk5oWPRV3Vc24A8ogmcGg6t3hwdFK2YAlCXTjYoTm2Tnunt
a5ETba1AZRd51A2ObklVHX8Hpw4UsoZkIoef88L3Rl4VBoA+F24N4Vb1GouS
6LDfizg8P7x45knx8UJIYrXgNxab807rljhqTabo7bdAhAEtQtd2YaCaAVL6
EK+CljKFzBimC8boRQZj2UE6PCDD7KF/DOd47pb4w10xyVIjuoiI35k7ITx/
9frPtnu2arfwXU++lE2yjJTnG31ZK67pJUHmIMwcdR7rMh13ZMPduehRvTPi
NEkLDkTBYmivZTyUIepfMGju860b6sY+u3ID8rfAlfKapn0q3aTilQtPjHoB
OFtWjRbG1GXuPGrtzzNinex4shg3LNeKfn4cl3k9Fr647ioQN3NlGaIAvD3j
1YfDhYHHWwif4oDxz/+aX5ksY99DFuf+pJIySvRPcA3M08nKN9nT/zlluQlQ
5Xt1pRX91zQ6nEqh4rBEyvtqMEzOy23cADjcOICCsTuCYha9QuD9UK8hTrIv
+oxntaKl4HTlX7z69FPv+ZiR94ESumGfcNZZhDHY7+SopRMEXo3xAsoKCXp7
TdVUM7XI9eYWL5jxhOgJJmcoaCJaFApFg1s/2q1px6VD4whgM/g61ZbtMkIO
x6XO9c/8XFJx0RHI/I3Xvamjz8c4aTC0oaFgmhbULwA1+hp2Lnqmf8N7v4UQ
1DFVS1Hfb3IbmC5ZSvDWydZebcqy5r+FQ9Tliq69SpUNGj1X9NrdJdDwbX59
RSCWQVjewgB1kwHydveo6qBojKGN/PdktULxh5wrIRlo1/wt85OHflqK9+3O
Ucromkl2OqMc90YlBAq8DZ9zhzDSe/UzaeDHHASZGuxUzzG8xh88oQembe/J
kDwoZULbhQgsmpyDKCWDhyhfV0/MYjVCTdmGVUITMwY7E7oJHQp6h/OtvBoO
/YeLrB4PPe33XIdyanpS9MU1mqhHo0NehI5+P+o91KrtLGNEEXdCCalIGbhX
qekgWf0d3IBqljQj0ZARQTiv8oJe6rHL1VwtJzWcaS3Jx7a5AN3UsvgaKV5V
GMxihMYF3NJrAkfr0ir4yt7ZZjeEUG98Dc0G7oYHKF1U817vrfxcN9CEwV9j
h1BzfZFMJ3Wc2+RgvSHVUq194DIvu/Mc3cOu05Mc15XQfWmNXY0GEG8Lrtxs
nesDWzM9btVdTr4ZBvDy0azfd7e2M/g8Pd5EFvWwVeERvchoI6jZSyjicy1z
E+SYMHCl6FwA09f53d62VDNkzWenVpwRbIXzbCsGYUDb/9qSOkKQcua+W6tY
kQ9B5jPeMGxRznlI+4ZZY2iIEe/ntUaegbDiSJ5/o8NUtYGlzz3PZUB/+o51
7GFcvUluz1YlmnmYbKXQygLrqjqBx1hMdD+CYmnifE/eYar9ob9BfdmUee8J
eKTYTcTSBG5No63McaoAV4YZu4nArIC98MOa2FdvjO2ajKbHwiCKsrywbELe
NsbXVOj1y+8ZDx2sqoLkcWtNLwkVbKFdpVSqeUtvtKXkQU7s4r+R5izkTtUe
biQVA8rLNhcUG7ILBs6512HNhbYvi0A8nFaM9XniQ4Vn/7zhyhw4UminoOJi
x7NIqpybb1OGKQZBYy4E21YyrrXLjQ68IsSoPyhejrx2ItaLlrauhm4kVs8/
R4LxcAZzGzGXc9Nx4uvqUq0mA7pSLisiF/XXxxDr8Exq0Awgnj4g8DbhHnml
wdHexGa69j1VcUOhZCMAihHfxvrpsAbusfNU/69ZiG4IYIuA2oWtupvklchY
jeJA4CRkFQ2bDxqmLUgUb0+pVyQNHbt2bzZyRRyc6YwzOVH3Hz+ZVgaU19YS
0XK7okivKx228+BfwLHHuCt1co9VbuGmfplsSxlLS+4V1R3IZsx64ceBwpEA
9g+ZST0PTcFYEoIJWPPa6wPzLT+VoCXShEaOMqUxxZHCFugysPxbWLylDFZA
U2+eDwj9WxE2EvltPqM+O869NC/43zeNRz2sQq4sIZhqj7d93BezBQDWosgz
43kyB2wplj3x26zTsj1VEWuzRKIfj/pnv9AWUEYm0PhjIlo4B1qCEJMl6Cxm
ryvQmoiopgYP1CdhU2hFht0HaNs8oG2ckUr9d2hdvzjcaH3/X3ivUw9G6M16
/P41//pRtrkhg1HYFy6NByasJ0Q9tG99v5A+XT62gVM1FBfwxvIEucDar+66
w1hwy1FjlzWXBqvRFUOCUT/x03VeZreKN4mvFCCOOQ0eSEZgrv5jKSLeUCHb
zX0XjlHgY6cNtSvfJs8HkKKyQ+UMflJP+Io1EysY3XZmArDpASjCClOF4q9J
nSiosUXWb51Il2wKmbXHIUPn1mLfa5j/6soN6r1FKxqs2VTVTe+1Q0XBTyu1
uMzMh4Imc63Bd4oTAg6fJBPTCMPIw7nJy7mImMHSR8vIz8U4nFViq5HjUTkI
b2U5m6EZAyqShTE6tq8N8rKMW76UTYgcDvBdfJWssew5c2MKeNzIjcFE5u1W
xB2tSWigIlm/Yr9oDlAhfYuwWdjeXRERJui40UR06eOBQ44DUDoACBREUjHP
dEgFn31ATUEPGfIMAgRrGUWwQf6lmHH9GHOGO5F6PjAYjVtSnHIorXkzmGkb
GhOzLPbb3Tl2Ic+QCnhdF96XcXYU6KQfSONMEkkslxjBoz+ucFf7qvbkvkaF
bu9Ws1/eBf5ooxXz07C8cCnwqAR3QvnCnOaf9pj18471tuMW3b45F5+2T1q9
Ru6cFVElJSS8gjOdxJk2wTl5TxCLfw1jSjWKlGoOGksRHfMUWIHurkRTYMU4
oj7rE338ZXrTA/yDKMpn/tneM5kCX7I1mQpwLNGbNFkrLnL502AKWu75Qmnl
vHK9/SwXm+0Rm/M4oz09hxqg2DYvvD3F9oRmcZJ/5SIX/GAxatoUSAE5+Tms
5yIauPqM474BhXkzHGdy7QQF5HsrGaQpk5MtcO3z7TEtBF+C56+WU2H2Audn
6dT2miWDJVnQJ+OudPQhJayMDSewwZ/25sJD9wvrFtf1bgIfdI/UKUU4fske
rmE1fxrhZLXPYHA6cmjzExytmVafXj7gdoEKcxEO4n6w0NhjYDMBCIClixBd
tTerE/kN8SFEP4ecaFWWH6rKSbKCXIpHJ7xPHAmj30GMiMVVNzTxbQwtcUDc
xtgaIUaBuQYHbE0sk44wIDrWQ2pPBYOxD3i9whByk12BBmL2T/kjczVA1+Kj
tgSjdNfX68eDOxGoLKab2uDXS7wPO4JN/hTEGdlZ4kitpq+pxYFBILPXcuqx
XTXD2sYpdzHGBZ4iFnIF9MhFhGMvaHIUbKQZx88c75quQSyM/DRir+cqF7qr
pfo/KDcShe9yY6EKBN/bXUFwaM9KxZt2kI5WyIt0yaPD1szexm9S1yGo/yvh
sSIXamojF9jjtmUIwzxblGdMfL/CBXNHXkE8AnDH9kGfDhe6DH8LKc4HpKBo
cdMTxUAjvgUdhBR92wbHNto+/kTxQvEdG3LOYQtgVfIVIuaavosFDmrCed/r
fKWKdWjiY1Q0Tsun8VM1JOsuEOtZoXVG09dH7/Vexw4KmauRu96Lf5Niwiyr
oSKWF6bLh03llNMV9oVc2KP3D68w1HM9vuyW+Dvj9UhvHG2PSsMMsUvDXI7v
rYV4R96A0jxyqgeKZ7rmR+jtNg/rdsdeY/UnQtDqWSSgxa1iK54SZQEsmf5A
J+J3LOOabVPCigsIIAe/eok9bk1NA5xcJJ+L5lh+yk4/wPMRoie9R0tbD7E3
GjOSsTK/dmAOQybZVj1HySH5TDEW81XdBBPKjMz9B6RRUSB1Q5Fa6eMtcnWW
zwInCmPtPnV8KjmhETBbA/XdrpSebYTlYDZZUu0H/Fx5O0EZZ5hB0lxHyk9W
9jhiUAEDaYn3ftQx488wsd3ZeK5oKQnJQybOuga61xZEQdD7kRgoVMAgMHyC
ob7kJEhWNGQ6TGh9tweG0Rze2kPnkYgqCzbugeO50PfAu0YP77fBFPJfNMtR
f0aQzqyb6sNWPcxKgwCw27Ni9y57Yi2EDrNyGDMKUPNcW4OEz4/CokgVNCP3
7dlcORT7j2QiSHT3imtWRTFs4ZQFPsjJxfI+7FVl2ejRM/bAnvXYrFL9a6H7
YNYZPM+6PkoUiyOUgqYiXXpnSAXR+EwKxWqYjpo3O38pVG93gk87FRpTLwca
BFW5Urjkkc/fT+pn9XPOjzk5NgszeOgTH1d3/hDMV5+me77dhGZey5vaSUri
LCGdva52Uj9zKYT/8JgPfLN6xFopJaA+YLoGaULvlKzJ5l+ALpKqZON8tmDr
OtcyKA8qb23jA/nyoDTLn7FHy/RtQDh1bjKgLcyx+rko8d6+fT/qRjzFlKGN
586BAYodvmV/R9qQpujlb36+JjeHW8sITTNprN/nX2Nlvcef5Gpv+H9kctv/
6f2ZqWdxUxLvEHZHcvHhJvPhUc0ZX8BZvjYg0A5X/zopX5TvSOA/FudRp/qA
M5EaYyPNCrTVEF51Y6PW2vqVLbtn48m++k8uBEFzUtGatGwYVH4Bh95BpWUV
/e6XjnSSDj4D3zoRc7KXwU7qsSVJ7MvgNWf26GaQqaLs7+6s4ULxOKlscN7c
IKOPW/JuH5Id60jTzPLZ+uJhhkfKvfIslN4zjLk7Nr9j4M3X/Ypl+5dBLUgO
Y3BPvx4+XHIInc4kewp325V7fU355iKSo3fDexLNbzF4H/g4iga4BlUr+AZr
Sd8oHH6UcAGLvtKo+x+gYv54k8LqHLBBYcFxCbeAChD9CkvTntHEESXMWLzw
JbaMwWt5GeOZ5ByyjkDCRsc6FJ2W4uI9aSuMItxCk1xliTG/niJEiwPenhGZ
4PJXxoc/osP2BeLxKgrxqDLhhKDp9kCn+NnRebl8IpNoQTldVxAUCviVNNFv
xnmOFl2Q6Fln27SqGOqrxzo6/frWhxBSRxMtwoBBgWLKsFK1hJLvyiwaGIhN
q9SPhOWlgy9QBx/Un1Krp/LF5BTt/K6OF6KKd9EMmqVhGBWedKaYccy7lY3w
89vpalm61oeyeM///U9FCylrQq80q0nDHvWygNzx0Mexko94t5X6+09Wua0l
TIpRHwskAz8losXUPt9OzTN7OGI+fs9nma5V4HzkMvXK23FyGjh9I1/BZ5Av
E0V5/4NFzunTvLZD9dX9ESwelyNp3RBZZTsZlC7qlDw+LhH5wzHkFMQn9Hof
qHoy5FDTy4SlTmvCtUZdziRk4vGXguMfu+HHYuBk4TejisPsojrrje7tDEHi
cNeNozBfnYY1cHUsjceLXivZkMvajLuAK+q8RgoRBzTOqzQw0i4DhurprQq3
GuFVWeMc3k68z+9+YAz4Em2Ec4S7Cka6mbiTteNUN9jgVHE0GF0Ocn0Ib9qH
bc4wibyTupjrbEdX62qWfVnODgVt2U9VxoDhXw1HpF7NLNf3r/ynBEnzoFU5
zWrcVG2iUbeKfu9TWGqwXkoDETdDtQSXVeZCmPr/tJuRvobub5VEPCCTTjI4
eUDCjOQRdj3TmZ/Qw6/sIPahMEM8pmROAKP7bUybrEwoHwF5AvDmgu4t4qxw
IXpy1iyjPcdJA5MfgG9/1611RI3bWEEuRYlYGF3vtmXHJcaXObX1kynLgPI6
on8X6wvR5638MAoweCXR1YEMLZlLpyZEmqH75waQDaKGNpSshnAMg45Gh7sN
IRVXuidKh2cLkfjyH1VVCdwdKzFd0ogC2xXCx2WTQqYSBMhj/N3q56LaAydK
bpRsqWLkoqOhScO21f4rWoIgsDUJqV/iG6yyu42kuq+9PchRG/7Mk/UAyQUS
UDJcFgDQAoaFB7lxBhtQHuzb/OifDW1hx1UdpvyXjyzi1IppUUWZwycqxd2k
JF8gEEKVf/MuGTbMwvdICZR9VI0Wru+mC+FmEbocNygu//OWjvq6EIqMtKm9
zqeGxJk9p9Y9gCQMQ2FA+SD2by8ZUjspHWzaO1id6eUyfkwVtJzoOGvR6bgG
Bq2LTmYzfLSQ8dkK7/snsifG8le8Evrx95M0x3FNlhX/w8TpQxzdfea8iDbk
ixdAgCZnzZgoiHSIDC/ofsr7aWPAYs2ZaTljc8Og6qbBhDTShNYLPTt4pZS3
ZTXYs5HgjfLlw0163YHO74UvqQPSa6WtSJVkDUuv30CWtygtzXUUG+iWNnAp
6w0std8f4itvFCa2YHWQkf/VWXYmAmRIH61SyPBzfWcr5AcbcpAPl+8x7EKw
yb78Gz0tgWKs/DwjisCLqEhO6TVJlLMiwJksf0mhey/Ylv1wvvg3L9ckQLLh
P9PN8ysprkC7xzpNoSVO7tw3QRXC0/SKe5znqhvjT1iRSAxz2+znwBAruad1
DJNRAB+kEZ0rpX4OFJ1c0YJl4VnHAVx8Z2O6KbTaetMLYXsaK/YH8/CpubhK
j32RZV+Xgu7LlMRawYL6Zlf9gJtRnUa0JNvyZ9kNZ0/MDA6SoCqdqnHVeLnk
7JWRBE5D8s0XhUA/H1BkdvaAoewr0MV2RGpX5CNADDL0hKUAjddPZb7iDKjo
gv2ImP0fMWKhDYjkZss9S4wMGvrnMoEtk0m2cvs1l4e5QrBZxmgFK8hbkxE8
SSRs3EIfrF8Fov9POMQsfz0VITVCDUDPnC9KmcbF68MRLJJ/MErwVaig2tNj
OL71og5rjOkeEeexzLi1YkIXkDgD8SAAc/j1dNm7pnmD9jdr0d/d087CyJS6
olGES4n6x3jhGY3HPziH/g1HEGGqA/FOJKk5mjzcL4u2rt4YdVJ0/Ain64vy
BGBnApB5q68M6Z3L+0+JLInpZ55e5ECQg9/q0owIdTABSETqk1R9c9tpfoGI
4cG9bmlFDbuFlnneqgRMHYWoQikOvl0qCmCjrjVA8yHtzHbLKqRva1oSb6lv
OX5ZfIFax5QrDGyYnav224Zii2RrrjgRKzg8HvBrCxbuyuMDzpEnkwSqGZzY
+Ap5FqmEoyzuLmmvbdWsJ9ZbGOs03jsRw8akIybahWePohffVZokFdRI/NbP
rEoV2/gDzUEHh87Dh/nbSXzOJ2U0HUk4CXdswIokHO6Yeh2pHd3SNbsqQqEN
ahRTinSGOSXGh9POZ1kbWrSvxscNJuBcHc5zgGEbccKcm0XqZPqr7N5njCAU
3lh3B+ksbDeIJdTgGH5OJLCHkNnR+Fc1kJFYzRgoOGsQ9s64XjUdIOTilNQW
Hdkad9FcQ1KcKI6ljjhimRmH6lqHVEPRGmQjYIqi8pN6UafS/U24zrsNiM4u
6X4Gbmd7OVEY+zvAqI+A3yNVhBkl6RmYDESdIkv+bN3GqJjUOxU21/XHR0nq
AuGqW2l+HgKGsQwhXoIT2PnBgOXbPks275ss9fZVdAVLCQHWHsJZPljvHAV9
P4uoUOF1jqFq7trGByUzCmXuDwaHOsB+gA27Ufm0aJAuwqLfX0dV/YMiD/Qn
Tt/ERjjlzbxnjtuXzJxKUIy1rp348ugk2JmrrEHBrPK8gpIOcFcxKN26M5Ts
wSS40IiDSF+Z+UIKKL7yNtDwxyICV9tCPSLVL+/LkD+lLpVYZUw0dfA1OkIq
4VbYpqgGPN42/A405kM34uIcQ5dv0YezX1yaPHhNmIKwoC+8j+HrKyaVbzQf
bYmEL624qylYYwpOwPw0m4LHep2uR6rfn0KYaTQyvzMvVDxWjRNvjCVK78Jl
CeMwHA8BX+lZn0HJ2+lXZUq8s9v7uKaie0AWvImV36L65vVRqVvGUmvQ6ao/
TBsVpB3ipU2TJQevtiLrPO6Z88P0hHgWRj07lbWRVSl2ZszjyhKNq2UkQ5xq
vktAm62apBwQUaHab9LuuNYAm8vBbxpWyivCMekC/elM2F/8o7Es6qPP/Tb9
e0dmU4a+vybmTBPz62Yiok2HaA1S0YkmkjWcZ26PcCH4iz6LNJkmbJGZbwpV
WN6wXoMIuZEfMA2JJjc/Hyoxoz+g9hVuX8DdhJVYe095tpaWcdNwKbgwK2zU
HTduMHRu4I/ujchfq+xYDYeYx32TTbwZtUIvy6JMW816R0Uu6CRvn6X96Pa8
QQo13DK2IjSHq7DXbmdtBrgdX8IpkkuE9MBrU4dNx7tbca8rKTYSKL2RU2u+
HTH7Z4tUd7qKEz4kt6+WpRJ0RwZdGt2KN7sLoJJaTsLpO9YCFo4ZdD2Us8g9
sOKJmwPUuR+RQpYQhA23gxDUX2I0XPxI3zE17x+vqgzvtM7QvMPm5z+a9feA
sZdGovgTaJ+hi5+4/daMQIr4sr33x5gMmiiuRQNL55M5aSoZvRIDu+w2P1fu
+uz2vc1HZCuzDLTReJnzpxnpdZ5OWrIEayyfQvgxtoQXMZm6K0GY1TupPUe/
2jriM8kQ/lMJfLc7W7RonXbHV9fAH2O7E2ykWMB1mT7X0m730R/iacbC41SB
eBNfox82KfYy9KtBesT2yd7hUzMjJCej3ulgUsuuI87vEkTj/3DGA3Cdy8ky
xIFukGkbwKU5Gf7P19uKBOxjoxsfmA8YeeIJmMVUsMXPbTbjjLUCBXkzHVxU
xN/1VLdZ6+NwMpnzoTLbnEZh1tnPtbCFCNQ+PDpg4g2LiKBsYCBynnAymMH+
x5dWQoQnDrjJLokEMLCJMBosFLOihX+fCuRZMEhoPt/IF+wFQ99oOAmx5deD
PtUJz1S3EU25N9AyMKbKQhi6n/+Y8Z4u++piHozpqRJe1NK8AeyqDJ5MuTun
eGAA/4G4WPrABvRphFFg1TtrX/Dc4M4ad+NkdQ635JrpMB4iayLbJAhRc6Xy
F7su867DKR2hPleQkEZxFYarYo7HAIkRtc5ikapq2lbEpVIaMaUQXQXmNd7h
7TTwvWvCMiS3emwYIYRN8x0zcPA9u+7MZ8Bc2CD4nsXePtTOXK4J2t7BWKyf
OZxfleHcsk66ak+sldCmWgSRou9nkhJritCbHPjXDBil3/6HspsPQJraveQQ
5d2dyeyuCPUGiJWiLNyscSHq2pZvzKe5ZOTa1V3YnqZ3G+HJAPphOMwxa3Di
zzFPoDTB2HpWj8PE3B4vo08DDYS1HZgFkZG/nJKWqITgeskGrhgH0RJxvZl1
3enNhQCx0z5SXtJgo6gkJre91HvSD0TzsuA2hIlk4tX4u3hoO7k+sATmrYNc
Rnr4K9BIYt1Uvhpr0blKN4RXWJj4oGa+ao1kPkP0sWAkEim/lfBiUkLfzIxP
8aT7FDToI14FDfAersGTD6jqmoaWZWzc38f2wntE4wJWeix9y/0mVFoU2TUa
YAUeTh/1BFqtJeZLFCnjUfuIQlHTZ1PcHb3TPB2N68g/yZ/a4CUlT2hGJNdD
SO3vYJh3X/D5wAt1KUz3jnhgN8X67CQLc9kXKjlCOo3H+cOutnKc9NBLWDur
qAshHgY9jfrYnI1BB2cjz1fdXsigT2VmE5lJrW6u4YkYwaKuFs43RHmBASxp
8gxR/22YcWYl/lUTe0aAebA63NX4OwjoW/fJd+65MLduZ9z7DwH8cL8TLmd5
u31raYWp3d5i4ODDZxw+7BDaKMzH8Tdm3KbyCg8U1B9azCyYolzQr33QRSZB
CRui+A2At0yszb0dCh6Ryu0vn2NkZl1tBIveqNz6JAloAl10d2pbKYdSEmqX
drWO0DYJufi5bqV49wruNdi1ULGFqNo8q8P6NulSXAl0QewXj5it3y6ILz+M
0iBeLWZDTmHdzPJSFjtzc7bF5MjTdFKzlBRefT3UYTK1RwOEWA5rlEic+l9C
hQxOpRFQysR+VHWTboohmUmXpEhRrsu/dnOZrtLu5JFLxAJLeCeTa3KOZcG5
6OJPIO7dk9ZSqz2kbeicIZ8kFdxv5i0jslatXNTUFZdJSNQZBWhsCB/tZ+Eo
IeqK1OWyWG30t5Bafpl3jiQd3Y887mu/ru4p8460jIY3GER45AZxGjZ+XK1K
Nt1JKsJMGghlTcKfyQm21qXRa6Vuvy3/qbQJzKD+FTWf7PxfROJ0SrLGZoY+
SxWQc1AF8pW9IuXR9HuH1dX4obkQ5bjsgX74yCDBMFogZ2wrlvKoryNi2rlU
EsIYI6dnlwAPpEenCOqPMeXGbpguZccdNhZ51CXdBFYj89TAXJ/dnwOCdrL2
a4fy8oveF41Kck/YFBH6n2ow5jVb/2G1kMDVuWhu4f4ejv9SdO3gG/RPaHKE
WpTy7f++3SZPQ0vroSFeNR39PNZ6ZEMcyPTjxVChgUspLm9xF8diU4E0YPRp
8dxivONkISJMD6CHPz8I8QyjzjK9I9Z5yukmRNrUDNWhEIrCKQ4Y9kkeEB6C
RtQ5ZqO3jZg7pfahKxcPtpruyodTlPlC8VugALpVTisA/GRWcRW40m+CzoGp
iFod7p9HFzhtKyrmKhkza/Yzhp8rPGlibn2Da5gt0J2bOEDchoOPyDbhAHIV
RzXVBHnzNR46ofSHe/83hfLBMKHPVOnTqhfcl6rHiVp4BL6CwzsCwJikL1UN
97547lLm0zZw7YBcmvBFIFEhPkH7fIIom518LNP+FgQvhunp38W7iXThP5vV
5SXU4jR3+LpGCuemJBW+22do4MmDTWLwPZEVMRJExfyxvtH10/UvzgotTNsP
fpE58fJ7i/7VOlxcBCBuAshu6sFY2CZ0SITa/lZrTgFjFIZK0AAPuhYMlju3
HqE4p3vkdpMeB+uTPmBQza547iAWCdwTrR8N87zJGIygt+ABsef2a59filSM
kmNzk54A4D5wxKS3piKjUzYiJWmWRcRXgbyYVJiRWrLeH1Y6ChrXU1E/Y07O
Kl8bdDffgOiVXnHPib3225Y515stFR/9VNtWsVBCIEwnh1M7uFFnfnhq5ozC
DT8jA2utOt1JGvagW8q3FkO5cGLAyCsqJ45kWwIBBXm8W5T0b1yUOsVn0GLj
P7ojjQK3nOx9JEgJrz8KfcvY9yrzekd/xma2It823Jg8/JZr5iT5a1SkY5fv
ZyTOcdi5nB7j6aC8fX5mO3pu7+dWYmnmnPrknqEOsBUXvnoDYD8T1b9+edDQ
mhIX/Snf84cNsvfMii7PNbgLJmteoL+7GPOHPaVbVHbeLdhdjmCng8lpO4cq
67Dqxd4ZeX6hXl9W2wJCPsvUFDRlAgfQA5yqlWFq/ZLCOqsihKyvckU1PUBR
vOkKppgmQJoT160cngjB5Q4NvgrgX6QDRbR1e+ObT6fAooHp77B5BnI4Dmgm
YNGPXDdhOgUkRw+x0nW2DZB0sEUJhFePYbLpwWWT+5tgTP0cvOr5ATVlBjkr
CRL5BAz9k/qShKIxL3+KijgMmrKts1nuZPLcX9wbo9iBLWT2qUw+j41P0qnj
v6vXgIIhReSlfrkQyB158gtgblmy19cP+tWFcoyGhBSt/yvZU5Wx7Oxfn7rO
1VS6tYjzkVgyv61z99f51rVn66s+IcZMOVI5Rd3WVTr8BU41sisyUbISccUe
we6gRqbcE6KHU4JW7iDm2zUT9ud83EGxxFkShD4SF8ruO9U2BYlQcWt3NNnh
1OrD224urY3HJrtLhfUhAd6NAceqNdlvl4bBIUO2FQ9zQ6qQncSlWTwfq4Mf
C/f2DxATdTWtWoU19AjY3yL+xq5vdwG7DvUQOISF6e1D4ju8MmMkAeM5ezhu
6U8c5DMOY6ojyc1ZHr6fZu658O6nKvBK/jSxbCGqRyFgsWBXtGuChC9Xiwyj
oYWp6JjkiOWOL0/iusakuxUPD1oORQQPNGsxfrkip6Mgt7IeKAYjQ7yEskvz
/3zH5c1ubo5vI1epY58BoLKisvBvJGnuPkm78x/fuuFM5xS2pqb0iG3orTAM
39/YIYKeqjSZw7t69tMMm2bR/ycyjmVPwOVjQNj3DMUDYJ4DXD5vjQMbDylW
IdD2Pj0K4nM8E5HqaKlcQpt169zrzK2yii0Ya0ru7dEIjkz3Sa9jxJ+NU2R5
HKf6ZebEjvmZOmvGRvvE0pS55OMPId377t3ReSNZBDrK11BdGS0c5mpNB6+6
jzTdgYnmR9XZSLzsEeTSEOMXSl+Vf6vFHGmJ1xfl5YEkPpMaCje4zYTbbNAe
c+RMkBE2UQ9xRaCVnF+SfhtYsoF3q9TMJlfen3mXY3RVHXt510bNCRd0AskF
dcItA3IDnh5k81pXWZk639n9lbzV7udktDz2bhSMRyTRgMhm1Dhbi7mbZM96
XehqUlOer+C6YUcICN582+ddG6UHp8jVASBkKOoKy5o7M+E9C/SjeviEyOTQ
iWA5nBaXY/IGJZHWuuYGsjXGfkxmHi+JYA10tqc84vWawxtaVN+IoacGKAnU
+biz+ZjD2oTzldCQ13lMiCmlLLWyxYh1WY4rrS+tpfiwiFK4RvalMx2yWE65
GDDDwB1IEW01+Wohbk3XMo7bJk4Kbt5x2WTF8jMo2co/9ghWsHNZTblQqY31
XOdJSC9QdfePdEV6LJvK55ux6AnBfkAJY/pgArWd3t4BMS6vO/bdEVBVtT5n
FG7Y3DfpWYWaNW4Q3VaFpN6mWxqMhYS6FFVslm6ml2ILdsJvdUU562SaBEuM
hg48J/EOpqoFjTX1B70JJmhs3Hr+mfVSDHPLfD4n9NR6H/nosL3kZVoZSuoM
z12bboHaKdFBFt0OShZtcSkUtd8ouRw4hh8ixTgwlxMZ2eqy4H2AbbpaT9f+
FiW/cr4CKrNIxLu/bfYq+52LOYUSUDGj8M8z1E0M5e4bM1uMqiy7cpIgca2b
XGjKrBbmoKTWhzd4VuBNwGOpbQYVrzv5hdcNVQZU/wnqFjKOnLOV4Kbgnh65
ie7ICauxEa8JjXkprT8meGAtOyn/iMmqZDsn72OkZIaI0Af3EAOKNI8oCiYM
OtS/1eDX+9PhrOjrunVYt+XqLl6X9vTW/Y2ZRmoNrAZoi+8hhG058bFCQts2
4CIKoHRxTTULEp4iTNy3JW2MPpl7iRri2nUGRBFXdmNenpE1VfAPocU0JCiu
iO/KU8rsYkSDOlAfubqcQPSej1Qd237Q5DePvCVfsZjZrAAh9jYZIn4wV41A
KUWzq3ffG+ydVwIBlI3mgLESxywhohnaPPXh70oVBncKVq0h4okZy67cPPrY
u1TNAxlGsTiOYyk+8IzuDnJlGV2Tjc2GGG4mDkqPBFe1/e8GBK1n7Rt2r3/N
o3x40GRHs/KvDiya5zgiLmC1OWpNabcT2GyJvMPUqedLocaVQiMOmmf76Q2V
wSQ7S/4epCUW1SRfBEiEBrJG7oWuXWnCYFfYs/BxR4/jTllXXMLK2/A4RhS5
BLA6UJSIPCN5Vnu14rTDWcaBidfO7Co2gVPSapBJNzCNdPqiTVK5stkO8q6k
ZEAupVbK2Z/dV2s1UIxdSj+3qbXp7B5otCLBCbAx8XQO7u4tGlsXy93+ehz8
h2Tz26nvIzvD/fG0r02xYcqMeOK3wohYcVfsJWsL27GCsLbrskhSSbuAbPeH
ePTugnCG4+I9hOdtLNNYiDbglDd7HmmR6yTrA/RtcEKprSuJei1I+9K3vm6O
zkdGFGSoj6cBBzIBaAxeDVIWoybHPFeP8OHSb3TjfNkPyu3FQ6wHGBtcO5Lk
r2oXBT4mQ9g+jNS3YtE+0se/s3vPeHo47CzDdhpMgYTH8JkZvgZwNguRnbyj
cW9ViqLEvwzc0j/djWAuooUnPN/bIRhTBaau20sc77EBetXInvloUkCE93Z0
NBHaPd/4vUDu3vaX0nz0VB0mK1kPzWDFCopRTBLL8D0ABaVrDELPkD7t9aF2
dLonwZdwZm34YIaJLpqyuDK6mAbDPEultStUqrZrqL6Zba4W8F+1jQ+L/1uj
ONY+YIQh6e4uAUM/ygmJX1A6/TQ3jqwimrm0NKLMQjpcMdvX1lK79Sd8BXNf
M2Cp8tku+XTnVSek2s2b0bFpq7D1CUaeIowwElT52JyIZEidwWp56IW7Dx94
Ai02RLvirOi8gKXyvTqe01Zx/+pBGtewsclvVXlbUPzU+393++4BZO3IoPUN
ov6CHOJK38PduhFLIm4SFWKEa4fKdyBhhc5iPWfsQFx20qcw2jKtt5HIS9qX
iAziWw/LHw0PyL/ZLZuz/CrB5H8An/h5MN1KHGiUej4AmOGvZA0Lkc77hULM
QM81s51EetxNJbQeuR1W7wzGFoThjZ5IldRReqPz0tadSoUaDEBUZONfZREG
BPc+hhKlrKnuIncKjdYX3Ts5sf5fjavQUULk3SWAVxOrvm3kLfcCLyOgGsPf
3ASXuTHe9jPTkbPYBm/6l7rgm6TyLjecJhAb3QZkcecW94ViKeD/sVkTVzXs
AU+pJsURPMt9BOxkl/NMMn2nL80GuzJFYOW1EYBGxG6PRq46GS/CwUFhOd9q
zbDh0Jh19yJ3VV8LA/GvrSLE4Q804jeROD3VzGRZPoMvYRGqpeO42ldvq6eS
XNRccRuz5+hO0AoRyT0YOmemdRwhYyow9obrnCABuz6l04RgAVUayMweJYoU
JKwBWlOBtoCKm8/Ql12tOsWoaUCnILQhgWP4bJmWhw3HEq1ht8VLlSaL/cNU
OdbcOPi5AahicNkYb4BNnaLCD13vAXaR7yThfmMLtl6PVVyGes1zixrRxbcC
xauD3iMrXz4CwBQGp37onQJTOrFBfL0GULl19Biaa2QCHrhpy7K+fAq/lk0l
KnbsZpIyOXnEkQKj7f+gnPbUpCK0EUOrecq4rMvHYe0mSzZCrXypZJKybj1n
tWhIzblUDmkegSdQgbMdH1tu7OPZZhNxwn3xImbsKgIfr2kT6cnPXNuCdLc1
XpY8Lpprr9ehH+yMnpxga6N46RoVuhVncKGQkm60vBVlUtJ0qiRYRi2gkKxd
Oj5lFiIaPTwncSYnQcuPta28gqLFdS0pD0ZpBvW6QK/iwNCxu55sh8o/gESX
ju70F8Hs9cJkoaBnJS1JSduC/op7ga+cNY0tUzBOILVHye+rd8Wfuu7H+m7x
z5aKlKvotSeZsICjwQRbBKw5B1cldCqu7mnPSOMcmPn3MK0abwUHTRVuf4Ty
0xkRS8Gx09gvV9sQDca/y/yUDLEK5tmxIiyGpTJ8mA9rNvVqzNT/JJNVaPhs
P31xCfWxjVMqemiQ6YluXXpDnTTMl4puKTsbkJhbFqOwq5P5rT0aO4Xh+qzl
wZki69szLRsDiXZm7nIAd61OFnN/eS0jPKH/5ropKAErW8Z5IjHzINe00J68
G0LLFeMcycPCJN4016KDWMN7yMUMuEN9X13gVa+ggXPoQysxSK/Kz5Q7z+z8
Ti+p2qcV6dBZ0MnYqRBAujpyZ9SsUl9yinCGxjX2HmXBa3HcZxfM83AruEaO
neKL25fl/3tRnVW44h5usZWQ6ZWKO8qRAkxSzi2w13mzdPKXMltv7QNPcGEE
sahWSGluy8trdFJsjuPIPDh+vpgv6/NoIXxFfvlh6uAM6FXqSHelj361mwvt
xwNN9GUeUFKs2LkSY5P2RovKZwb2auPKC5jBcmcILeP300/x/8iy2t7vvflp
EL3ZYMNaehfz77nKPjeG6lyiXhfecsn7nfyRQSC8LfTTUERcLTx7T8FQTG6R
axXRZyG10MmqjA/NQCogci102I5z69jXLqUKsF3MFb1AjSO7poUpkBZlJGtx
Y2i+Ryl0G6uDvLFKbfbLsZBo0/lu1kb+MkVcyQBFWnRLe+IM1wC+FpSDVm2y
beOCCWqaHoOjkFa7DHKYLa4f7lmc4Ajo8f3WONIKWAGAPiG/YJ7suyUY01HX
l0gcrHY+wy25xO278+qkYrHszP5JynHLDVabdd0l1IoNL+lmp8C9ndPn7xDX
ws/1UvaefssvQheBtEY8hs0gxZniwuuRSD0rEbddMD0qvAVgGOMj34fbkonO
+9UhlYactYIFgiOVdXe5DkbHl5CqHhDa6BoGcLirIc2eLzf8n8J/9fdHtcZZ
yY6jjJY6AQCc5ZR25KwkRXsNAljpnufmq5dNgCEV10BAJ0HLHWeZDsDDFhyE
1HyWVlmvlIxMYR780F6CvgZ2Eynk7p31v9zH3hkIk8EdprR8HUn8OiEfiK0W
m0R6VxNx1WnXsoKal/1P69id/vciSJlywgE9L7c3Isp6mVvl4LQqL7Xlovd5
F+vAewdfx+JQezKZY4+T55BlbJY5TNyQf2srflVep1ocI+mELsuuhFJkhcsw
ozRH406Nm1CuHFqzr5+HJl1/tjANHsOAN0m+JkrdYHXQRLVLs8mPIDPvbnXR
GbXhlZGyUOwW8mogwj2gSM081oOa3sHomIuSPUgv2y37uM67tp6OBEEdccS0
EZ4pW8MrtLBI7/x84k3g6KC0bwvKrVUzQ5zG26wQW4Uo6HwowMjl1sVQlkoS
S5pwWYmOjITCKX/bmTOuwt+fpyKHVQoA70nOwTAttYf1T6YeRpfYAKLgpEOQ
OCxbJJxZX4H/Oz7xVACSN1Njrj5vvV2hr1n6gEtw6KAvnJr/yMpkQEW9YnZy
TFSl9JuI+TlTS9AC86vx9uuxsCoytCIG9zhpzs9TP9/qC6j2WFitWAgG61/o
74uotKScdEv2q/tEJ7ylZw2541RoEJj9YfPsZHKQ8nGu7zBZLT+hHOn+QZHo
6MkLGcH3Fwr4w1Pmk3zDB36IYhVorRgrupkPO9UWPaL1XZu5cswGIbRJJDuy
sWsnh7Antpu6EHcDHZrv1YyMcCnDlUgtLVo2F0xOtZo+QfGQ/xHQ7qW3r3ep
kjU1xwdhPUUBU7Wc0yrkgvTOjnBYAEtwujWELhVBMm9jddPZKbcXr+1N9iBY
1iYPAHsVfxxB2ZiowIyVMMODrzEhvddlHaLY9XqQGhJyJ0e+8gAdPZhWEO8R
OpbBfkOrzGN5lsW8VwvhE44LKCQ6gvgMrPkO4DMwsuZtbSIYWKSuT5dHlzI8
BF0r0QGFIcbcKVfO3jzYhkP8r9anK6QH23svixpZuwE/lh/1eQcfXNzUobNr
1WAC4m64dAW9p/xq2yi+0xHFtnPlVI7JaiAqjDNmnaw8L/T4OEZ3UulnHdQ7
D/NZU6pp1rJUI+/Pr34zIscr3lj2lAMMgZ3LXADzuE1AMd1QmIZwOHYyBdv3
4sacEkBmDgzNS+JzAt/TIzfmhvd50I7Dh4PrGkYO+u6YaJxiJ2me1BjTAS4p
otEJGFFUQzo0AiEWxiw3cGURqzBesATQSv4f08Scqd4naKQBJbE0XO0phDv4
izK89xuxoaiLA5OTnzoqihLebxm3auZsiFfBqPjB3xf6CQIIdxYQMQ9Ks5ow
C3MqSxLCByC7ur/l6XNDO3CDaJgE3tKZQYmtWxmY3yodzs6/B8b32j0xFflY
PKOS2X9KBSP/NYrNQ3iwEC/3kvMRWSRjYkC/riLt++A6W5twLzBoC84XiBls
RkqZARahw3sb87znPwPVoPiA9KVoHdh6aC2ZBIPhHmb2ey8mbTvdeEovFyDl
XsfSA6QowGW6TRXO+BGx8mwcsa4cCHsr/RsyhY1izuwZ+6No6f94gA0feQ1C
Qc+X9DwBpZ2pqNn/qd1QhB1Zk+NE+Que/XswLiy/ImN+76P3NSLK6FrivdYd
kbnSK43V8jKknqbnihldMIs4wXORjn148dxg2HjpedhNYETSGYysmcMk1ThR
euiVY8jUErTx+vksKk+nw3Ojwc5wjIJCo95lkkxZmcFfwMYbsh3cG/oKUW1P
0PpMvfvlCMUe4dPAliX/YDmFvemRBs2jxPNcjkcuR8AfbgNgDeuobW2ZTWla
XSGi/yCsfvN57KzcJ0aWhcRAc8Cqc7KTKwPpz5BxqIyfYmJtk55qYqTfPIMW
jkdwVXUuAHo6s4UZYzn+fRngfBVXRarDqNqC1roUsYk/Oa3qLVGgDCchlTXx
zq+T0YCaC+Hxj3R3AE4neAE7SSr7DZVYmfzmu9NviCLOUBzGzUiRZIGFMMKK
95pxLUGAxcQtHYVpaaRMpjDe0Jn61KKzHSmKRFWWX781Cw9Q7agK64cgPJLw
u5cZgawfu7B3O320s8cC3r9XhbcCRQ6uhxf64a2wLGkK4lfi5Fhh4yq9hlT5
UC7T/ja3FvQEZW1zFZA0/12fuzSpI/c4V2wbJp54YiZr5pO/QAOizPlqlk8T
pTomrTQK4fr5QaBqCrxqbHjUzKIvgyxeviQXq0ZxsLrYlrRSUDlDa0zh3nH4
jzBsb6mym+U8m/Jr/WN6qnd3CflKAzLSwKDyJnqu/9+Ytmrk3lIO1MqAoIiY
2/oE29IMkrsZ8xhBo+3g7CVG2CHmV9kO+oxUm7xUDCK49jOfelFV9tJsdRZn
JAmPB0b+16Ofzx2LhVzelBl+BxmFB4JsfklRpKLrEZIJenJs8C8lf3hqcpjj
DOlFnHnqiK1yewGQlZsLWME7risIfc+cIkmug+ejwPurWmRhX2ZUbPeXRL+p
/EXpSiB5b48yF6IYAOGxmaUK6Nq1LmeSPx/osnGOvySGuXR8tO7CHOcGE034
Cb1L9c3+nZNNlgERTOj60IZUBbWMwRrVYS8cAyc0ogsQDVWFcGFll42goWXZ
9H4mNT+T5qg9FEEKMhM0DEG9yW+KziuOBxd9rmV4V8DoBxKBoMj8SGMfT93D
1RUDOnmu06BklNJsDZfcM0w6Z7+nTltUjv8uvAVdCZJdFqoOc+JiqSMTczv9
EcfcqprivRKtYqOQv5yWprcW4NzNlHd+9t8oOYY4ckQHJkYx9aYD+d5lCDtm
tIZqdH9UZHWCJoV4qqVT2TP+vKNTo2Ep1SA5MhJoKbFNrqxIo8SjmMTUUfys
iF7d+C0RE8igLieJU4y4JDOgcvaemwz9JXFc5VSnyEqWqd/BRBdhqA0bk20i
D8Q838rsDFSRwsH9Zrb3Ua+dXp94QVTzqmJ+ubF491+SP6cPdpgMp68FeVcC
3RkNrxNkRQ09pstMPc314mZT+cPTtPJjG6q4NfOFxApc74DSR9Viq5XI0rMP
Gqs258Pk0AfNGmHHkYOieIYCWTJRyWx+Z7KNKyFlKq3Y9hRkNIZeWlYv3mVR
MimOrSqBo6PuKvQbAzpQVco673A+IYC11C/1yoOiLzgzwq1kiQkI/G519q48
wp4Mny9QUw1IMb+x2e9kSgs/DUc1RU8RceJQot2Xh1KsTq8Bf4LreE7IrJ8U
JDCbdONomM1DablO+DxLDNPBCziNZ/097rxpvjeWYO/P2UmM+OjvGHybti1g
ZD7MPXwmWt2aCDN0pXSbYg8TYMyzuSMqZkh1Osr1gPk8v7X6BuYEVM68+uDe
22KV4uPblvc/3jcrG/eROAXSiQBAZn0iP8Y1g1uGuINHFKYR1xsJ4RNpa9vK
MLo06Mfvuy5tI95Aygmh53J7aosE7s7mpxkpJevj/g+jkdL9em9AgE43PS3s
nLY9BKJWTvMJwF7EeHDP6UZ/EKaKcN8DJpnt8ZZi/C6zLPa+7ogcNyQV7LMB
sdnTn1dbNxv0pY74orncooNuGnZTyACEBA7MYy5Sp1d8rxsmVE+4PN1RThHb
YlnXbuFLy0I6sC80ziCp1az+M/tygUW5gI0PzVvvoP0h161EDvAYJ3iJusTC
YndJGHboE/A925UMZoyudt5EyFLiFrM/vos1opBmE0CHwe3qzAXS34SgqFix
zoRFlMLVzn+o8DSamZHLyxc6hO9+5kKjdN5Fcjl1EifcgoiznmdJo0hbCzph
JKJiM01m5a9R995ugSAJGNSlqcjZSaWe/XVIkbPld+7oCCxfVghvpNFO5EPX
WtxNJZUxHDEvKuRakdwU5s+cIGPMl6WxEDmKKKF4vKcyIq2QRUBEOSLItQGX
VBZyWlZhOlEbmu/MD0T1Od/m0oB0BjvhEL69U3Az9pP3o4naFqL/23tlfP+a
9xLAmbkGg35Ex+E2zNipB4Lp/9OzHUk54VhzDLHfZLdbmvbDadrvz4NriT0A
4V9O/ZMeqYNk29J+hCqNegvG5C93jYXKRmDO3kD76QC91cHiPS+2P6i0r1LW
WCTp62sWGcjXsmpHH3ZvngZSjbsuZbUMtFdBH40HxPnux1hvAce1YYb6Awko
bA+SPosMKkaL7EsYiLb3Y5KUt8gRvWGsRLvrhkqFA27dumU7DLq7jOR/HU5e
C8ExwsJAfWn2PYFFOPVxaty+OGDMxKxHTu7L/ieDCM6skKBtjvDPtlwfwMYh
RCb14MYRn6/9G0JBiSSrQqlBbE/ejox5w8cDDygWHU1kt+Pq/NDcDOmHYoq+
nGOPNkZM0sqKbgymXXKqHyppsKs+MslcWoTgjor7slwBSi1LBPwHGcOus5Mr
T5muUlDjkpdRhhizqtUf/xXl3rsUUenQOC3wrGw1Ax2msvWgPP7tavnn6akq
7f7dMCngLCM4IRj9d/rb3tXPrxPZcopz3Xmi7YYE6H6FC8MGNYxw0a9CJENf
dzdiSn1ir2f6Hi7Ai4SZHjsEe3X2WbDHfp/wqIR8ipFAYcrR6x+Fa+LYPMbf
o2PpNIXJV6aKdNfQTeSe61lxi+836YTC+/VnKf9uWCiwcpdsmVK8c0vpl0DD
h3BS4Qll5Q5Hu2efkIiGSnqkNj3e2WF70spfwcFeO/xsVCOaFTJmTMv5HvoG
ro74Leg/4rfHEbeGMP3sC6rLsFFtWwOHot8gg1y4HaJ5nCS2POMuJpLnJmDW
Cp+/mkWlK8W0B04LWAXwaBMD3nDQVqtDr7T0rhMPPSp0d7C0nDf9IqoLJVuK
TuQdhk6besO93q2Y0+zDSF1p5102J3k5z1lIpRojPYXXQ3bJLDuCaeCFRnp7
Psg6MJuisiHcYujmuhy0mUnODkaOnnopBCI8PxxTVnhUybU3KOWEvdkgYWSn
tj77C5F5R1+4SPZS04GIoUDZopPmi1iwfVjOfMvS02JbQFVo4b2G0ohbJP70
ZGjsi3vrc3+VyXVMaQk0JDeOViS5pjqNTIgCiIchmY+M/OyU4dlN/mSM4YEN
Olbvaokqf1R+WlH9ZC+PVu1KXb0dgOx5hY06uAGucLEHiZ16378RUjzKhs6l
H2AZkJk15zbrMZoZTkwEPmqzOJRmaI75E0M1wR+qK33gBPDX3KocbZRPHMZ+
x1q+MSntVqIUlrrtnXk7Ph6qokipXAqSZ7Gede4QCcJ/5cQ9ifw3N7A63YYq
Dp9K64KyLwCka89FLyQYfjSQibJssPFSNk/RLFa3/MsxNQDV7gt+gdkd6Xfq
PJsa/JPn/N1RRbCwDy4LBYmkW/9pC4fwxDAHetGWHRUG7om1nxBsOZniWRCR
w4PgYknxm8xEiBaCz01AC+TfTUXsuBRGsRBdrCNbYL8joqJ7OjjIcTTqEmLl
EFkLlSuOmFSMf2ANUCD1pGj5qqdgsE126XvS8Ym9hSYhf/r3SSnjmpkwPmcA
DwNztlbZTCwqfsquU8yjDsUgC4SMqcx8xJYLOT+Ir4TsctgshaGAzIGooEqC
pbJTdT5mvhWV1dgX8TRUA/+p0L1s8VgIHLP+q6QwzK3HgObTq7AhNgy8uoR+
1sMfZhPaSaYWyjuNSfjjg2exlwekQFhgq0aP/oiWEqgsygR4PSNyBK8/WCJz
9fQ3G77lhLOFmCKscXar6X6cbuGQ5Dq5hoYC/sMNmjwKfWWM+BCem35/w1KS
Qz5qhmDRf8VYMewAFO/zTWM4Cra7VVUTF7A8DKfNWzqBPdVlZBpR+QCdLCWg
baWBRTCMyUA6D20A3SzTzVRL3eC+cKcIKBKraikfcevql5DafAryHrlc8Mnr
aOxpXk4XWexyW24RNObO0dVz+tNx1PU3RVcalaGMmhZbuXkwlJmkBfI3E66h
2KMklo/RrM945RDoqpP9o45RzNOxMdPSlp1rzhRK+0tkNWTHuOVp6VQIGNyJ
4wpXIdHbJyqPvbDIW7bNRPvXjAVYVVEgdrk8bapcUh3mmY4BpXFIBtUw9crf
Gy9vWtr52HjmOY7xIbOtXu7glbJhf+2PJuiNoHg+wYaCvPi+jsoFZ0UECyjv
vz853w9QxDHEhWW3Z/xl46GYA5+mJuR4r3aXsi31UIMqYwP6WVD6WOoSLfZ/
myMwUumdy50QiEB7fceVAQDwSaFtjcb4NyWbDQQQ1bQMZJHriNjHZAMDxPjo
ka0QOmV0svHeELmG4UCIgyCwxtifvwrx2gsUCRGb6ZBVazIpCNdDcS2ciyg2
wBoq4wreTn5Bn2iDebznEJCwnxBqqlom311v/1wQE3kS2Mb7qQu5Zh7UD/sz
LOYGdY3/3gNhgICdJIlStvZlM4iR4PAoPSERd+Ksk7ghJHmfS5QsHQtU0lHG
wdNNFfcASQvskSwg4fzNbdRplHuxBO11PGu9oONd2kbYuILckeosf8a1TyPl
F8tNOrMQhWlJT3otIWZ8Mp7C2VBKIXcvR5u67YNKi2v5FIHU6rP5nAqtH0Vr
kPYOyb4Y64mQ+93m+6HzCXw8wXvOufNlt7yVhjoB/Yy1mTXdezV0gPHrN16/
XAWbADpQECg3RV+Fq9blrL4/kQE5A9kcyLVcdP6janoaCZ8wVSkguZbE3Erq
S8sypmJfn+x0pAk5CVYTI7m4IqFWZapSyzFXx7/gnjS9rbl5ndtcUkO8/c9v
J0t9xRsgSvFHxT6BCh/RP0O/0FtTZR840+vD0cdC5+jbpFGHQLeDON7bZZTD
VTJbuuSmLJvQAFLqV1YFN52CkcRaRa46e+Ctwi8r0C+zEjdvhWIxiGCH+dhd
b4R4feQcjIggBxj9LzU0SoHQR5Pp/e8NqfZcmp84fv1QdvL0PV5r+kMwPNOP
7REo3EsJghf83ilBIiPgP84uanmqla9xUrqSEq/tUD0J306QMBB5UpPZ4ruG
GgyzA5UzOGUmYtWNZrrO9xPOJFeAjFxukk7SlCXCddx7E2HgKqdoZ3qugDCX
P9AAw44Q5xlcCzMHXgaN+67EBXQ/Y+B3lczokMmffRcxl3dxhKNdL8Inm/sM
3AMKWB/Xf+5A+LDGEelpVuZ07jzxCp8pqujKzsrxaBWKcQtz/pTvJwk9mX21
VquOkXewbFZzLLYlP46axCwXslT1ccuAYFSNnci8W8+Sc/i/dmJNC7if+Xe5
EPaq+7EZaUQXKUI+m4X3dXCYykDSZBKINkJyMr+5A7sID/08owbkx8fi7biW
EtcC1eIHAmcRXmXu9jm/KJRd6BoPNCmFTWdltHf7ygpn+cdrjJiyJiz7CbLm
7EOn2jiJ4W4dojqlDKtYKS0TZMuva+dpOi/PU+ebzcrn7N4ZlIeI9qeEF+Bt
WkZHHyQPKBVRe7dlDZByTXlx0kyd0ZGQdh4uzLbiquYbPlJpdgYMgSJ3vxSb
ds/vu+vGyC/tnfb3+jT+Z4RnHSniEMFz7lDqvSrLhNZEiFkMBh4o17L7W/no
ifW+yIfqW5wFN3ekCFDAxveF10bVFUJ1u2Hl+7wy7gv9WOZXgBWK/pOEjIIR
dAfsTKCwGv65TgqcB0LK3CJnZNNpmTnNFmCjankhu4zb9HYU0ru3LeTGXWe0
Hn7rO7XdBwh8XzUa+t6ztsXWpiGBhQ8T41hBTYpfQiofc00qejFkwgVrw2p/
L1wIByB1NV/wb3IPKTWBTSqrl63oBaF+UM5NXFCZZXLW6hNHf+iDXFwZqBZU
71fvhhAy5MLOZnJTsHfejQ0HgjYkLmhlbNFaL2/gqsTgEtJ1YmCSpo4Vtpr/
68dUT9FGuOz9cQrqZKxpfLb8Rgq/JhZYt9DnhMLbiwlHnU7EGBwTT44tZu+Z
6bWQPNKWg5H7QkiZ3HAomLbZKJNBiEfabjOPJCbCQif83lW9OH75uAJHSUH+
xpaLVtYLkOXTwdCFdFy9xILoHXH7m9yzPMBnVnz8vvKAz21NCIN6xHwfWX3k
i7NnptjDa4RgRrdcfKjD6mFFrjqEGRYztl9k4hERAoLu4Kf+jqVG6M2CXEgu
JsDfNGKsoKy7W/j6eyiTJVr7dPorqdaRyIKY69y7BG9rAVaRPC78ybrKLwdk
PQpG1oAVJcUdLJt0vSnNrAgNOJIlbAE1WV/p3VevrJh5uYkFMLpLKIbND/8h
Mse5cN81t600fzFBhYa8PF8pUXcIUXjO99WhyrOblwjE87Bh9XbkxpGJQy/a
sRyleWjgM5QvNVnJyxIJ6NNwY6W4FrMJphCUdKY2ljez7YMJ0VWhgHuGvIf2
L6K1GPoVJO9QqG5566jXNdseLNBCr38QSkBKPsWWyNYSFBnPAMOuRj1w6dbx
D7ibDzT9X5t42M+wZZ7hxa9EB//HqRa89/XdV1dIlEQjtLOBSNtI1s2xgaLC
g/m0epOT96nfWABJbwLu0DVqPTrTRsmBI+6RhN/PTswRTLQLpbXjsiO11F/G
c3h9/TxoNgx0YdOuE+JzJsNIlXDrRsIQYfMlg5M7fSSqL1Jk/rtzFBrpzGNw
+jajTvrBtR4h/x1wjLamct7Dkbx5rBIoGmZTrE+JmWIUwaKTJ3vynY+ybrLw
VlAINO6QPC+jqh6+3SLzyzHbVNZNkgXSUbDJQ7sYlnNK7KH7K4asjKv/MdoS
y9ezUcWUgwVFjBhGs8/aHA5xH4d2OS6mtPr3IyvJsr8+HbvF+0hC26wX8mjl
RT2WNvZfXF1C4F0G4INKoWkHTyMDpocSaaXsenLQoDGuUg5wK5+O9oGSHgm0
dNmekrOg1P4T+HQ9CxOi4VuA+y21pi2evMJTcL1U8xWzQ/BxV5oNpznb1zfg
yEW4FY+9V3UA1YA/Wv1LmBKhPThE+T/jRxrwn8rPMAizHPkW9Uw9s8Qvkeye
MCKh37NmmmlUDuXbuZ73dFuuJDbBPQhwpvNkS5lSrpCspjglWM6gU/1+HyBD
chVbPZk2G16JbFBscO+amoNwh5V3nx7B4xF/FMj6jbjRPIgrCS1xB0b9xXYc
pTYP6GagvkF0sl2uMNUs8mp1rJ6vhn1zn9qxUZSmgwX8da50WtUx+b+z9va/
dRgPN/IV4LwpJteuvucZeAK6i1Dt1O1T1RuZd6Ga8cTW+UPlFjv4WPU0/nOr
VxjinvPuqaflFWltHsAjNmuKUhFfWeK1fnSmUF6lwp4giNJY2YjeefuWyw/j
DK/qfSGeHa273hqDCy9acWfExNrERAgpHe0BXYgKFcItV939KydtsvNuiCKK
kZjjyrFNfKi8H4p9OKWl7QK50nE5PL/y1OKn39eaQhBY/kNV8tn0r0H63nRU
EIZg5rC/5fvPN6IZcc6ISRg/qlQsuS0oYSEteOknZ03ea8ztzosP7eiomLNE
2ofzGJceAuiizJ/00qjbhuasnTz3w4LzMbrldQfq6eGWGUtocw84rE1Vc4fI
9Y+munw6fYSHhoT/BYDikkGDNy1EHU83srjeUubVcyUw4L9cwx0B14nqSOBT
qKAM+bjsCiAg8CcFZvPLkGpDsYRnA6oZRnCQsl8zQlYh+P12xPZU1ie15ZzV
XRykirbANDNZVZovKeE8EQ3fHyT+R2eeMe1DuQsg3pG0W5Zn+pIKDo4B3mi6
dKQCVMWE68NMIKkcYmg8x62D5yg4gFpnVLtxPEsXkKc651e5ac0DTnlIvKPG
ACN21Nd/YW1b2vDw9v0Bq9hLQwm0rnpuOhpGUraVPIn1YFeaC0/9yrTh2Vps
8+LHeh11ySTpHe30FNhvJzSjyYF5ngHpfR6I6mM4V9wQavcCaCW+qYGzyeVj
6hlR5bOIPv7WAxdHhLTOmbKP07BdAKkuHyACVbNVyDa6ZnW5tIZsuZdEij4u
pUURypMm7uoWKH56Y/ldXtDAzrbaR2OcxRF78/AExnWwZb3pITd3UVc4HbDz
HdCdUtMLav2xPSr//VHQxznmIGyZN0epbUm5YBVZF6oTCfa5aWtw/dTWHnuX
4NzImY59vMg6F5QlcMQxuzu+T49ERkjJGxkgFKZ2MWD4QyDGILyxjUE4ze5O
tInKUoUX685nb9iQQn9O1Nm3jlKPgKy9EjAcMTefLzlLRT57Wlo2npUgJTFw
gRny+TbcPHM1BmugLu16Nd6+0uizUwCq1R5ONqaKHPmt5hL9T/k8Z2pCoAW1
UUMFYHzEhuMFMYvjmnrVHz07HxdGyA456F1vHhESbyzluUs0gKrGNiqUnCvB
9ZNdGMbGVeDZsZtLsXVWBEohkrbq4krnsAoVpciK9WjTDmlZRTrItWdFqyOO
a9x6KPz4kePc94wuUYLMZpt5aEcwhPdIyRHR6mIAvsHkOSTcnm5BtVW+AmGq
q3BYRK4DWw85PFCFxBuxGhUd0A6HxvjXKNAa7nrKr+GtDFhI7R0DhDwp8uSy
UerQ3U1rQHvY+xHm0fsp2CJgTdtQu4ZvXeLrbJRsWTwwe2w/2zJQ92VTNCc4
V6S/VpqKJLivp5y9f2wkFj0pYlXKT6qX7NE4c2cQ5uM4FSNEd8cNEKRE+Eco
fe1SvKraLCiNQ8tzpIqgJQCfvRztkVQbB63hgYLYSJ/LcC9YhFpKbU6MmyH7
b1mpjjbHaeRBApDGLFoo1lelW5Jf54p8O2PFF72AM9JisOEwrykdo2L42UkS
3kSpTt5Y+urnRNv/U5uMwKLCgnSVf5wGVWTZEPDf+t9udIETbMzqqEtUSZjW
bNxOnDvo3A2yyElbFw0yyQi6VgAgBO+aDbjZM6SbiynxQBBWeUOpxa5oQTmR
OkiF8Sw6MCmU3TfqQjdHRxCLSRCkd6q71yYveQA/oLAPV5GdZDLqpKJyFx00
2uAuRzAle8bcAj2D8xDduEZ3z/J5gDUJjiWqRUwCf5+SxPws8gM63deoX9QP
fWRbzf7TdKckCkAF9/0k0iGM27qeNQD7FkzLV9t0q6nSwun1sWJ0LzsiCSbL
ylyWLWgohz4YPFoxFUD1Iz199O0PxLkHHSWQHvk/vST2FFl/Y1sbAexaYKvP
XRRHXJlGUpqo8/n2KCoM9KJqpcR6kRen/MzfqSZDawWGDXvWFURA2yXBQCrV
bv8wpdbK/wVGwf0Mf8rMjCn5d9lMaOWNN4h6IDIzz4G3kIeJClT0Xa3C9BiS
4iRDLkjMO5DCrKeBMEcocdVEToRbSatJnMMQ5SJ+KqfT+9nNR4eb6OjKiBMO
Mwb+3LGhtTCkA/ZPGtz/sJMv6O08csxGcywciSd2Bk/OcM8LL/PEj3kxD61V
k45R7+ssBnNRhAXSZraPFVODA+MJwJTgQ+UDVxEi2olfbIZjcBBywEN0nxvO
C6CVG9AD1lVnWy6hRxIWmkxnM/vuBuOahseW3DObx3prpNHDlle+43/kh58k
yOM290HqRXU4QbotXXPQNtGAnY05ccI4QtXrGo427Bh0oa0/55n/rgIZiGFb
KbIG/v3kGqstv7QjHz80FGXyUNajsnv0ExGqPnebUtB9y1qHY0fnPeXWmlEC
djY/89Ys4xOyE7uM6Ygq2fAxdYOGwDsAgh4PLu6PDPFcaWvWXqi0AnA1gvQl
sKKD1nBDILgZsuAh+d8ntdZdRq1ofKD0Aq0h1IlgLP7xlzHIUcu47htSmm+g
UDF1YbvFmdl92fVYf2WWS9OfxC8T5rYpZTd711glrrIYnPx0QIAXtBI2kX3r
XhpA/aivSV/+YaYoLqrDPBvxlLOcK2qdPTcflUM0NiWKOG+cA/L6iVoADJZx
DxTa9NsukE5yqeDfIXoKdm6Hw00+Jq6OM2S2CH482BBG02n8axZrb8j9Ys+J
pysKCgXQtX8wXYhiriB68SPzwaN78RprOCyrsNh8er+RkjG0E7Ja0uaj714N
JtH/MCzcoQ8juViWffUhoFsKaixm4WJ/8zQ30Q2LRwC2jtWFzCBABsiyEp8R
/niaJapkH8bcA+90UVpdETAqv//arlfPFBIy6mQHsNSNbpw9i62ZiDayIYeY
5WiZrrnBycNwzJ4xm9Q2LBKzhKukILYGH4tVKvQw37wSTLXaVTxhEeegmx32
gNXWq5Hq7Ft7rUwVyNdYiJwoPHlQ6m/lRqVl0Y+4EOj7XTGv+7T9YC56DkfJ
sAz3SfM3wKqHoQSd+0ZBhh1aFrlmGrFBTUcJgFsCvmOzv+2CFw2N1n0P1Lwc
QWodWnKvbnD/KGoYrRTNJFiEuSyd1eYUM7w1XWmmo6msWXiLn5uuM0RmPiOy
LvaCE4wSvs3D8OdO4RvBCmf14zAphMlC7nWzwvpHKPl5bMWDmugrjtw/rv2p
yqMMJaK0JQnO+5U1axJggsMeXADLRDggde5wJYUnCx/5wONtyHGFnJqH4jpW
WK1lYyOV6m16sYz0J0/5kZ2JU9eguI8lGFA5BNNO7BqZefrBzLe5/6Oav5cT
DeHFe85xC1hhn5h+nM3OwaItLN6VK+MowYo/AMtNqMpDaB95XJpjsSSpC1K4
f5aJCyxZO1cVOLyl7GNQ8XGLRb1o8DlgJ32BpErOJe5RIDuKy1MQzvZeoywE
6lhSClXbhATmJTVr8wOafcoHa+sDQNedWXbU2GDuulGRQx+PNwivgfXCMs0n
B4JdHWE7RzJZiT8EYye8b1hMYWFifWIKw4SB7k6InrRBF0fO8jqUU9mRK1d0
VQJ9zWxiN/vgyaRYOnvp5m5nSiB9DPh1GfgF88/+X1Xy2ZUCkUXUjWg6agcO
ZZu99J8O+tf3+4BVNfXIm2Cdslx+S0fRMdyTnfaMyQ67fWoVaif5F64j9IN5
LsmSghHBurxGjCSEpOQj3TB0msY3QjLrMBeffrvz0j/53Og8Z5z6DloYuzpS
MxpZ4d1TaTHv+Y4AQiSA35dHv1h6CDGwCvF3kBCwHW3WmZe3/NVlW8fcpt3v
LXIa/ME2d2fnecfci01dXkUVcJFanW9xXTkJ3zBiHDXaIHyTuc1jFR5Bc3LF
67NiYi7YdG130PAMmqtZyXDf8vDoejqlWUSb0gPRO5HKvWk0eph5oYV+rrCv
A9fbTxLc7oOvuN5UabtpA6X6HlJbC8ObQnNZWWgYDM2jj8b/01FoCOAm+5mR
YyV0k6mvLMZ1D0A+tJrbX88aaxhRW/nms22b4btnPdoYuwic4VSgT/CYRlMk
RvqGv/TguDubHpgmlB6NDxrl3+8+e5elMYzfufWw++1eyvzJ3x0j2jIJDSGM
Dz1YndTaxWvsAqyN1nWILgeMCWhQP+s9iky0Vgi2rH6oCNxJDS8y28HUVyH3
BDbmN/0CtRasnoKnQ3eMzGHVYwG6BEyue5rEIKYoMZLa8B5s4a5NqLlL8qdM
kPQU7ODLZEly9V8Kk3uPAo2OIroNmOO0otHnHRmc3qmIJzPKSeP5bhnKOOTC
ogThLbw/OEQrtojImJIgEhQyHgXRTyFS4KuUuwnY77QpSINuCy2D+EseyyGV
SYq7o2ijbqRWR2pEDOzzMfZ+oTxSnlfuaUlweaT2OaIU2KxS5r2azKy7QCPk
+mqy7MCffWnKqrIz/w41MkEiP8LdBhsl7/ld46G8VA5kTEZ4ncMmC0ADKsYe
VtmcK7RbN2+wZOzAGPONpRdTUOZva3c7LQLjzhiwa+U4TcCWSPfqcLzHVAN3
v9W+QNZIqRzYepXedI21CeElEyQpcL9DY3ISAPP7T45AAaDwzb07Kwtngz2r
eazbkoayTGdAH1iXZBKzyLyA0XQRM7XXctGz8vBWal7duaIHEWtwOSkrxdIm
ecnQH2y1gkU05tUIAsS26DtslHJpW612V2qIMh/tUVB7AqdNsR5pBFUoyKBt
bWJiowOQW9FUQ5xYEadfrlMB1IU9GBKqA4by/7WQSUrPQp523FiyvfWUyBZm
x9dZ5+KlgBn5+bnnnoH4RN5i+XJacOA3uWQCeaDY1zzH9g8VlTM/EYLTO9/5
tMmr3HNGQKadrZBSZz1zjaElkeZNHiwXqh2ATm/S1+jvlVNs/lFqHUZ6POgd
6ehg10+KSnRXgAopy9wP2QCWO+sFPLzx5pjkKCBhUxgrklREnmOgdxj14qta
Iy8cMlFIXosQaVLHseb0McXpwuZ0OYeOee+gPPdCa0iETyVtpaIJL/6AZ0Dv
8zC4hu3fw22zxajP728f/zd4fflbr2xInBUcHreWvh6ZdPdKx60CxoUTrVNq
qSYhJWR9HCJ8ektCqGuVC/QYwRQCVe/BJQLYtQKuquFP6Ggx94h1rmS/GSpB
IZuEV5cChlcXi7qQU0LD2zi1wvBdcE5R8uRXr1zI5V45KNiobKAv69R0S5Xe
8duKKmzZQ9+UPX5B70w6NNSmIfXnU1dpVe73BP43UiOGJYRSnx5EI+nZb2xu
hzZcVRBe2fo+2KvBk2CxCdjMHM52eIYGdBAEBcbnyD+ClmZMLcWeL9f0HdGB
gIgfRf4GWEotJ9rydlFvoYfe6SoK73mBhLN0fy/gjHEd8ZxwGe8vWNBmVPb9
vGuEkXLdpyL3GycCwc+/hfZvAaQ/kCTKxMDAO7oQ0L4BsQSk9KgGDFQYbnJO
zmw3QxrUBgwd/LsHloAcpH3vwaiogng1gnNHPfQbCS6eYlobaFExDplTRUGz
6erNPWsoHH/x8MSRyy7J9Cdy4LmJwBiVO34xsItBl9NVgPFSnxdaZDr4Y48k
ySZ3D9fUwC+DHEoq39Lmtoq6kx0P9pqB3EujVunlhyJoan7iWP4ksndlA6vj
VsJCfYuV06D6Bxr0A1/iKbFB1Y9R4Xvc1xRW3piKy18gwwIW9y5Kn634lBeL
XQq3+W27I57G0Lc7tXn7EhV4fmcG3XXXYwQxNCWdMwFNIV2fSQYognYj8X41
enYUV5ExmlCZr+4HpgMxLQQArGixbiEsZb3jCm2qQnGhCMr+QTvccTuegCl+
ibPJhp8IpxC75Rnrkfnqxa6FVYgBUILn5YXxgDlRd7nPAoyIPlywZz9/vgTQ
mUi/SY/JI+oTslp5pKwnI4Ov7TLUK5leoNzlC+B6C4Q3+3ts701guXALTNrG
IhacUMPPpEDVttonaJ2bEzKnBaPA4ZT1k3rEl0GAXTfITnXu4M+7bjKdrdL0
dVWwwgAEhQPhKWxce0pJcLKxv9IXl8vCQFOz6Opqxv+5kEv6iRdtdhG9OGgB
Txguo9ytuatoxQ98Kv9iCcMPgEof2q7PDU3ZbmUzpkhIjRryHco106T8JiFz
CyybgcimNpjMSyWbDwcACIPlVmF+Cse4qbhC8lbJ18s1hF/nNulbeEoC1+W1
UMAHo7Y6xrPZe0hQkfvWQB7yxHBsYDcJDeohvAZmcM5Lm7XsP58goVK+ijY9
gSVCfTRg8Ew2xiYYvMU+994YUajGgW7vr3pE2YOathoapGyByDP1YRxetsPa
hAJULLm3J9b8Yc2EDliVE/dGheHj3LaTg1b35pVGMZXoCaeBn8ncQawAfHwX
skKCld8Tq2Ls98qZp+AUIKDwFj5Fi2HzbQVvt5Ty1fao5PD1fPZl5UrO3h9M
5te2pfsQeAVBndQFFguXSbtiBXe5wRKJ5eL1qydhSqyjzWOaP7p32na8egfA
uE+dqFQds3soHdFIvifyvae7zBzyvD5PGX5WV2yDEG0Hbq0rY+/7gtYwB840
50xjbAeASA1dHfdfFngzrO+iMpyQnF2H4rIL4uMqajNoLRDHkRSauaC1SBb6
csbQgOt3RUnv0MA16qK/Kv1BR/ofyXIUbMDtlNKhWnwxOS3VXvNeaGs/i87q
QJguvRuVJKLt7jrjg23S3taxloviKFABAXP7BMwlvYfaFM+4mK8pdZ2iC0iq
NLdMs8En9vTEAhurh3vhM5O7PRNdZBAgw96eXsWgoFhidZ4aI4JEqTci12Ib
Ogyqr6PFeTVrtZizrN0D0cz9WecQvA6eRTMRk6EfrLDc5pSp7rhnUmXs8xjO
HOdl3p1cWQdVg0b0g68z2j8LPRqW5R7xjfsScjBJ/D+wk+pjmDzR2fXFD643
COVglojmSTxWLGdaC0NLpcHFceFBvRRk6RPtdrjEFA9gCi0awoxUFvkuwFGG
fr/SOz8xp0Gy661biczdYV9u1KtGckBJbEbYpRLbBdzOzpOndixdxDJDWSnB
LyMxJWXWFRFhGtxk2REac4Aqx06T4c1Whu8IL0vMNCr3klpzfe51KMExVdHj
dRhB8uvjGGwijkY4v184MieHBLJOLtZ7ilPSq+EP2BUnhzZMtIJhH3U/VS37
FNBOb1/X8Zft5pHFqrXRQgOaRS2p2TKGzyml6tQ+2WUTv5oNu0h7tk3JBHVI
2P3wG7malmEZoQDofCDCFsPslVZvR5JoDgDPyzLHLYD+9MgNusM7OHVe1h8w
z8dUsh7qAqEbV95sposmvEbPlhseS6tQmcaiCdje/5Og5yRwNr0f3JiBPlHT
IzncNwjasiUw9wNGm5T5DPpVZYaVOvZ+HWqpPVjHuXaUal6LJCceuMlTkhFP
3Q4sQqtwCL8gzYAp5u0Pbpo1S1zSt2/P/0DlElTH67U1kaxue8d4TjzdORz9
evZY44aU9pCPqeaeAG4X7MHkGMwrySUZTdxH6IW5O8omHBaclf03zYXtI9vr
QpQolebg60FzT6fSR4HxK1tE7/exkLwn7zZXAqfwYewf4f21S0F0SBpvgS3/
jXtug1uxSvkAqBU9nQgu0ZfnDORj1PhEBMbGpuOO54NYHn8346JLB+ekfG0J
POfv5502tjMOIK+k1qELYEyyrQ/ImXgSJk88s3fDrOXmT55+fGU5Pdzkkapg
xzPMOBhSuKfiiZovHvzzbnpA5jnxztlg9A25DRYlIaXvnDCxKs8/Jkhuy0ke
pnCRttjkMdyYWbJKMAMZ4gUtLb0a6jI4+Wl7UQPDOFVDBozly1sIjeVKA7oq
YNYEzOl2o+gCbYQwW4MpjWKeGBuGQCTtWDfOt1VsuQpr2nMdW3k+bLLXBt5F
kXtwVoYqv9AsQJEZEAvDq2AgCoi0QwMzykQIXxPQI7RoN8I4lgtayDSvdQYN
ti9FFzti4QawEm6UNETlciLGcCxdCEOH3fiz/TdrAcm22EiOBvTqUxxln68h
KTmXfJa8hEMwOKEl2N1bd2UPXfjvofWq5VJ2TlQ5a0X2hIH5sYOB2AIM15aB
NwuxzWQpqfUqe5KQegftRENyfMNfqCZSQVTFZORS5pZfHA3aA9vXFgPFWbk3
riIQmFgaBFKGTOZcRvb5uVkheKrOrcouEcaYPvKtwB1BXMQdgnAZxGTlwphx
2QbyJc6HgAmwx93dBz40JoGg0/DxAq7wxMShR84OuZaipvHclaGtq68Wu8LI
THwlEXV/pm9ulZGmvZmQ0EmdVzdu4auR3yfe8WUbmxV43UVepE4qnZmFbmAR
TPQQw5jWksNqMdHyv51x/wJsQILNqpTfMEVgzLBFn1/X5ve9auUGWiFI+uaz
i/sGyizcmaCJnjnzxTfchyPLnOsC58tCKkCnPi1LVrJbuT8qog2l4ipp2zvO
Yy/90pduS6qG3u3sxqTkAyWZp5QFtKTQ6R3HAakTNSVQajA+3QMIENt28ARl
gnLohxnLQ0EcqkC1Oy/Pvs2XlRl8C72nXLEvv1dlzUDfgJ9RSctLfnUXqLk5
doF4umzvvTgB9Muj89jS7AoiWu6Z3wuJ0+IeqBsqDmEBtSRT9z5Lm/8ZWiQ/
qB6Dp0FhmZqF9m9YT4/I3On2nwz+aeLvrPT3ywyioW0aM2rYnCoqB3lRl3jQ
TjNyt+s91CaKeWhQwIlqxdGhjRGoksWJZk1ufaJFu0RE7T6txL/t2ZcmUkux
u+Z6v6o/lBiAo+Cq2G4k/qsAYmlWooTJUgd2jOWomuDSv0vc9XuynaOUYVI3
V7COxHVzcLU76BRfX+GH+iIiHPmf2+of6TddhDg+HhgJkTCuQ7Zqd960lK1z
E+8jaQKirGV7w1djaugrgYAWN4o1cVtCUjZ3+oiHkfHOAPmlNtugPfbVgfpA
nrVSomBUESNBBSDMAuBU6Q0OvLr4FWCNcRrlXNsOZe7f5KEnMlfaYlvBGDEq
cts6AcdUx/jTVD9yke704vs/Dvi983uAds34s6cR1tG/lHHyxH3rfKINm5vs
igg3nQV5gwsJCbYkRY69JfbWU4DKpANzLiXjAz4Nok4CHiLH1klA1rtTw2gh
AEfDxors3wihgIzo9cKdcv77prJkS1LoHwTb/VlV5QeK26mEliCxbsVgY/3y
7RVcrSWktXHo+h5ZizkQwx1thE2rgzlx3SdEmZH9Vn9Yz2lu24ZDyV2Fe1k9
0xkWhVVwrVK06Dp33+Ar9ill6frFHdCBEpAFSylFrvi1fMxKom1FBD9jcje3
RYdrL+E+zzimCUk5giZZNnyl8pm99ZRIaXqq/OVg9YNInlNg05MKf4hbde+y
imjcD/WWQ2eUieH9MD5cx4DGuNndWPUm2SJ7+TyS+viMH9GRi13YH3ICOdrk
/2YXmK8VFzN6yMKx2OdLIvxANgVJiG8e/F4CkCHrpkBjqDzmOchB3Vrdc4Mm
bjfbCUU0TwOPTysp6Aujeau/3TAEoJh0DQ199fKILE1Zr2j/RK4zuQrGs6Zz
BFk4Y/dI4Y+AfgIBg1qBr+7HPQRmPXZ/Fj9y70Hw7uGsW3kRUKH4vipFrtQr
3IY9Jm0wEg7He5LBAlS52EnNVM/P41f2VQ6Ecs9nA2luemKiSPSIYIMFRWeD
lUSdwN4vf0Psgvkqh/I3MuoBUtKTS8UFRszDsch+R6tFEIudjZ6xILMWjmnx
r9Aym1JIzu7PniW7JwzITIhOSlKpNTF3L733Rj5l4RweQuIHpRSfEPN5Z1Ht
9wVOYvPiRbxR0GtFtM7fsLyD+M2vFhiuFkDeRu10AMlLm0Cn7+vVvLSgK064
5ANXHurTZba8FRTsvTGic6WwLkhTWkwF3LM7QfbZxCIqN203n4KfsUizS9rz
08b224pVBBEW+SAZnnk2lpC2hjoGk0T7g7ztYiYgBDLf1tg1FimW/G1W35uw
OuUVqCVjdCsi7yKgKZD1WiI3daliRwJ6ABP8POKaGs5AFfhrDUz3sTnZIKix
JeyWzQk+Wr4DS4wSLCkhx1jKgJdR1+x3af4GCeIEwHvM/uNZ0AqreCifrgm7
7of+Vacy3WtQqdfeEaOWYhiSaCw3ut3aP+fHfQhQk/Sm6Yk2Z1F16Y+4VVfh
nwI0dYJGxSEjcodS8flMq23456poSHSLMTwv7LMKQD0jIiTra5U7M7VrnJrV
F63RJlDSz5H/48FKb7YSxz36esyY8x1w4inWCFD2llnNLlFs+EbZKlptI5Fo
b91V8JJVapXuVkbQTGPs3NWumr9V3yc06DPSe/Te0Nz0Chm6ZGc+w02UDFj6
XHY/MeEQn2gNRXeFBZy0BHWFuFAs2DzcttmS5nCjhV/Rn1Twua0UMmyTsUlI
tJjtEIqnMZP40AsxUVmIsjsIQHI1mMbPSSfl0E36RMD9cp2rrKDCLAKYdC+Y
M0zxSskPsbfGNRizNcgxdxfXItG7wj83qg+uRTXZLXbTXeb72823bsMe22az
Z8Uo6DnnrE8AIfnicumPRjjsKflJi4Gix2PJIrsR7Ilrhnq2ZC/2D19p4TbI
S8fMtZRXr5wcevQuiIEpbOdiU0i9W2j2s6M/kiAjP0o2FjRD3MRXmOPQJ9JZ
Ro5g85YJ4JyWgcp73st3XG0Z4F6z1UWrM8ushF5T2lXrLSJS9kOFUV17rT16
A9xYSmdU7zygEdZ9l6TEhS/aMpZLv75YSkW8yAdGoO9DdZuWcQU7F+r94xYO
XWnpFSWJUnm3NYC03lXDU26u5Uzp7SgHzBwuC8DYHO0K9b4RimxPDNPMb9bU
cHCvmK4gLiBuLky6DCq8NfoL+tDhks6kSu9GUx85jnTEfTke2e2gBlprXeu1
4j6wNeXcrM1KvHOUo0ttG5APZ2rMkM9XCmVPCG4vr7zGPmGba4vMugV2iwME
i0U2JW29fn43V7OQhRNWN4XLCnXk3dslHs8chIeUWZFqc16yNZvzwDvkIvqG
9bqpPsHt+J5Cihj8OcUAEYhOmOXl43DK77woufkhaJ3lTIeuXfmx0afjjyZ+
BvXUbOtp74YEIAfu/KsIKaITxxluQu31OHTPsEmxTsWdu6s+FCoxcAzx30Ni
UFVgdxcg96mTYS/xEyfWzUkbNJ+a/D+wa5B1pkkyiX2JPieDnPeboiBIeMU/
Lck9YKV1uicYBPfI4ax+SOapQdu98gMvh4dIhCu1F3/qLugLTQ9F/HJGoA6T
AQ9EookkzErPaWwyAEGTKnUJyPtirQ+IweKU4O5D2hcWTzO6tdWidaF+TUgV
ICB8QTeljI3eOXD4MNDtGkIUI5LBNDhC9Xe3AH9c46SmNLauUcQlZh1J9Mjz
cf8X/D3Ofc4fxFbr7dKuJarBiDj8K70CoYtS0lxXSLYxHubqgMBLepVMIrCO
mhPw07voYPUVdWBPLNbXIpTF36NloDdk03m4AQAxKIfasUlrsS4oylMLRUsC
0u9qyoQKNNQHEWYWKVHPIG3SkJtKFgrio4zR8npYSx8/KywcJ5JfhAa5XxYb
LlzQfggLiTlEdI5attU9xCW96zK/sJmiAKXfKmjjy8/blt+ltS+6FmTx5n3T
innX6x9xj1ZBkO2uDTP2P8kJKE8Y13O6OXVZTSc9nVpiOG88urQw2lO30jHL
tBPfvKFHiVrK1MvXWXzTXhA+sh5H/D33PSyf8R+LN+O7lxXvh5KuzM90oXZu
2Rjab5RNfO10mgP8XooRYLPq6nOZZgZrNTlzK4S0IxjzLl5O2RpkVir0yOLL
QV6pAr7bJLUrMLzWfISeBOHGkbxE1lZP7BNZyH3zjKY89ZwhNp1yY8yt7gyh
Z3NxjKTqWOEkpWNbX+H9MdmGcxbfk5e6mQVhmTWbViTxIon+IsTVEyb0f/rh
qpD3nnsFepZzECvIatjqcfoAG32znL2ePZvlc6/lMHXHXUHZweUmdoBysV/T
UFCi77TwgY/putdjXHhOC2TrMYSkC5OGm2kLDkExEn9lC4/DiIg7MoudQv/S
urzpubABc1TOl+z5OfzroKi40qZCZaoJ5EU+bsn4WqQWdnYZqn+/Xr5xlmA9
65WLg0kXFuT82Hpz0M2gJga50Okey7qGPr3NGl5EExU+zBF51lRV1VQkOD07
o1G0gw9ShOZHa17bJ+xNaUAfl33nnGW35rLDBiIdIuxAHxAkHCIUNFMfTFRE
75EXDyxYHP+b9vo6XLMR/3JThkjP2s9mz7Pgog0YiIFyCAjdxzWrlvfefmEW
XppXknYOk79LHgV01t553TmNXLSnac2uK438zpjcEW1jQ+OlyX0qcqoz7eZb
tKAIB75fnKsmkxrSyqkhPEORTDKDQc2RicFYWvX+MsG6EHO6McqA1jXkOPG+
sXsc/bG2hYGXqP053ai5Q6KuQG31vCtnbWpOyeNuam29T9OgstJ6rX+YcveY
VRa6dEQkQX9jHmqfCx/xi2tcn5zdUKIp7X0+hFh6jBKnxhiCdBCJt/OAiLcJ
/LLLATmN1LxvtxDOuVua4b6cVTYOKa3hVdMQS6ekjzZ91KJ4vjW/2hr3eyHb
fxBa0eqRvVFINqiBkRFhqhmGS7CahU09IEplvIMKVoU1A+kgEZteaer/PKzx
W/0r6D66b6WDArwP3fMP0lBDM8D8D4aQb6C06KMMxDtaY1g8S71oNdEwTH+O
gFYU65zygGncZb/wp5IFD0L8UKLweJQIUWcx9U61bJQ1/waMoVsjYn74odWi
c6HDRPrRfOKop0MQ6al5GdbyMcwm3QgeGvyxSaBdy+lBgS4sc0lhY11yLAEL
8gocUV9CwZ6oG/nf87Vpu3NjsUFHIoR/Tw+L1QuN0taQ9fwAEiCSBBg3SdMT
wQUas2RfmYqZVZ3spVi/1jHpCZHsfbUfLLzmhAKafIa+NgiJ90Yi7jHEghYE
TiAHThREm4YCbtVk6PuQTrRkMWQAC98ENrq/dIgvwSwREPGbVXFAmdlsRF7l
vnwvWCXDn6TFCRyyGqQg7ULSCzEF4tp3l3ZW/Mi3evPRXB01IdB2PwlSYHHI
kR1gtW1ihtaN6UTlqr3UYdkhuaAQAkZTCNRR/TBt2PKgTrWdcKuxnHqW7b61
gdUlAWbqbRe8Lon7hBCpIljg09ttqddPSssh6ZfrZpKmDHMpEKNSgzpZ/ujV
Lxz2yN+eusCsSbMDXBn0ZtJw3JLgXDb1E4UB9XiSsd6P4ttCbwPAbUdv6/OY
+NN38j2U2rlRDoQlg+eUUzXYRiZOsIBWZrBDXg/3zwSN5AoyGeVdM3GExF1I
Xo9tFT5ILOhYtOVWuTNPaPluPpb0aSioykEMa47zgJp7ydsliwVvOUDyoaKr
YmiB4iKfyDWvI33z2Xm9C2wJ0eGnPmRdeO+hEhino9WdrqSJ6jdUccUu2zHF
E34RbmOX4YrNMuKYTg0OtXRb4rCrIQcrQ7sRpHp6qipM1sF3wRnH+MkXz4Tz
9mGgNMtHnmuFhjZzmDLrcMUIc+HMjDLjVGOY5fQE1JF1LN/ylMgCigRYfLBl
dTASY6WgqZmqVOioNdOGQB5p48dz9n9AvZ5fQFuSfkM9148N7WZ6c23oI0Px
2X4Ofs0p+rVeU3MFlAvniGnkVqbgTSCQmyFTi9uj2a4s4oU93D3UbvPsK56G
3ohYK2ydv6nguhPpC6peRgZL92S+SmNN5XBSKcQ4y0B5ll2Y9jn4mP/Op50i
4hzj+M8A4zoNXenl7Kdt2F1IcU7Fd2Rg8+EYXoQeXZLwNIPtR4XLTgsN61KW
Ws3DrDgStSTnk4bI5Ijr2xPD0U47p0Jm9ODbkhrcaTlL5gLX1SeZEUhiCxP7
XU141fk5iz/sxBLsxOziPuWQM0Ylc8GWOHQMKvPx7zoKM8DCmX9pDd2jCe+f
m9gsj4PKpbwLiw7N6c0Dae32d+WazxN8iu6Ua4pYohx72yaSJzXCBH5O5+ex
eqt4luyD3TYKgW8GcGRkbYhzNvuQ7r/Yetx91gi0Yw0RDIWizbXKOMuS5EY+
mpk6ENZepVh8Onhx4J5KGh2sRb4wL3XAN2dqoI8MptNtqrnDbZoq5t9pj8XC
hS12LesWfpjtRyOq4S2A7Zs8NCQWUphqTzCrZ1I8ic72LdshgMn2ZMEKiRdZ
a66E89KIv//3bwXPsiRh0iT/H04EDCpwKBDJ3tmXpA3+J9JELJo+DqlhX6Dz
uezLDYYjtaVMibe5irr0Z6PRQSGv/UWDENJNBscZO8gScSM/oeacWnKyj2EF
fkwB5FONcKa3IgEzCbVJ3xfvBTxmxKH7bscl56J+6sojp0LkSWwbiD3MA9at
UHeKTWqwiv/CIaVYAe3sX9V0AitjnPwBEmfyQ2wNd4rbuwGNrHR6veZ8twCI
ypGIcs/MDuUoyK0S+YlmqVWc1AEkKSd4P+zOPyixiSvROeyFxvUUWRZfnDl6
+uDjgHntk+AIy37lJF1g9+xVyJLS/5BmvvyY6/UgAlpO09HNF0Iw/OV5f+HJ
Nr5vH7RjI56W59bkB36h02LxNjA595bnC2Rk65XoCfjSCou4pLkaFkPIqNQ6
54fUeYZydOvXRnTYByhAJJG9wRpW4DO+PHAgKAbLtDVLFAqNbJ2WRR9k8IPP
abcao2eFBPGwqsTp0owfvBETEL2liFMTaaUNuwtllCCfZmFnXJcdbQbJUNzq
84TL1HqIcPfqE/3g95ZlGuxPTZTJbghHF/nVXpBgzmHDRTLq2dVUZhf77NcP
7zFbYwl6f8/PlWaWHYrK9PPfwBczaqShDCOgah76kNB1t2wB7VtyGWNPUkqF
Uq+vrabMk7TbOxuGD6emYKzyj/rEclIB4d5LdYaTKkSEgSsukejWpkYdw2H8
KmtqCr78VZyY9Uza8GvJEYtjlJ9/HLgxQPf5oyAGKuGW5AwXlc+/XpWN+A1g
YOWRCDgxHNWKnxPNXFY20AjE0lL3ITY07cX8IH4wScUgyCyIRpkWSfEEaaRi
+iXAio9bhSW+ktaViQFfFvidGOhddig2T9+8s+fQX8eY68m7RkhvbbAilrUk
vV4fz/+x5M29DLgqHTBBVE1Yj2KJTTqpfdu4HSpvliAoPIBQvWCo1KCjSrBv
sfPhd9CJ3OiTVArYAX+vgvPC0vDY8I2p3GZ3qas6tyEL7ygutkApC75f9yhs
dVmc4iQ2I/eBdXoY/XG5K/AYD4yaIR0TiABE8IqFGiKhkINNb6jvWHRkPFJG
bkXs3zkvxF3IEiraFF4e7EqDp94lpGlP6eDzHh3JtZpGvsYcSaYSc/5X0bMe
rimkYqQC1Gr+n2C0yHLb3kXghGiSuZWOV7hLlGXyJ7C6l6DnJg3tMi7FS7/Z
imEPQJlwBznBfKTPyfXFZCea6LCTjrj/UsuVWGUDDVuyn4bnVP0b/snN8yf7
6fH1aM4vRIf98CiKc866Tfc06ouTVszvp/xfRKTl1Cu1TIsqgClsWsk3Qlwe
YA2OJgzqAM2lDOCPR6gTbkuFztDadgLVZ7jN6IoOhhlaMAXg0RyFjUM4EgCz
QINl8JspuV67XNSyqYC7mGt70d+WhPxmnsoyL6MN3/UJ2v2v0Nr/eMyT1ZPh
tQZps3j2FKo7VSLQTKEtfG4aLoujUtH3XeLrsFLl9SYTR2BqWdG/A5xKJ7nl
eDiMG02Wp6gFZ+axTdKjE3D6UFuz0ipdqN5xk6kYlpT8SzEYOOFzbjIPnzdQ
e7b3AlGav32SCNg6rw/clktz5NrM1lVo7qh4QhCADy21PiwdTO0ftIE4ZU8c
REm34hB6odLUsuk/t3tl/pshOcMk1f82ni7GfmXQ4/CQ/C5A3z3HKHZTCvge
S25Mea+udsMQsxeIqruNmHDrgmZ/BUjsxHelvgFkxOBj9shZGlfW4+40qu6Z
HWap45RE3I0mx6VKSQVn/JShAUFlJe9E9JuruQyMFTRLVrsNaXz0bNPLnzSK
yTnZ4Jl/W3GkxF1+YhtVwZDbdlzeJ4eKDzZ/IL6YbuxYS7wyxSJBon+M2vlx
b2x3mjb1SjKUSyYKZu+kI/AtZ4Qr1Zb1M97dzmsbQYzelmn6L74z03gUFnjs
sqxRqqvUz6iYOrXVK+4178ITCB05Yis+O8GYsQeM4Dtxwx4oqM2gU+HgxlTM
xAe3X2crJNOuEUFoMp5NhXGEGp+Sn7UImDenRKoP7kjcZ4+sr1WoFjxsHw/2
DGvQa8rHTUO8wuGM663gKdrencfhZqrrhnDHWgt7/u7RrV47SYfupF/B7NmQ
PdhoaAc9JqxlgPUXb8UkZWFSgcTmZFRmuP63DcKPRgNdQSgbnZa+lf9L3Trq
tkyWkUBVYOJvhbbUenmoMkkbmedmMAkMcYMPRdN1Dc9ymZGg7pafmtY9S2pC
5nQtDpdRCpC8jCzmspaOHrjfKJxijJTqlce+sV93A5F3KDjcoPBiY6PvYqKJ
BFRyTvLx5WQM22JdCFxZqBwCIRHu0KyTt9IW4yyH64u1loQFCDc7vTLagBTK
2vUVAN7jss6iPV0fFnX03rOHHv9eZuRHgceINnE/2j6cBS2etKEBqP2r0QMw
B9F96uKrmJpEK/rkcnBXZX22/MyfrbWmIKY5jiPOHXaay6ao/sPfZHKQHPf/
qZmExDiuYUjkVCa7D3JuN5sG7B2xEYyv22Vp3ITCHQPp5KIRVnIGZqPh2uNG
HmaQjkFxwgmmY/8uOalDa25KN/aWJsH0DPnCsQOnRPFfNZ7yvl0PCNbRgrr5
CjBjvlYcX5OB/XLYQyJITdENd6T1Q8YMCH7gqmYBg2t9WLL6uPNR6BeGH1Fq
tY/XL6LJMmbmfKHRbcdBE6LsYKmSdI8CJnsvBR8PVQN6f1dDtkrXx5HGSWs9
8wGyccrjOZiFLtOpPRid509B2slv1gfujtFem0bOJ49ycBGWYv67/LelM1lU
b+AWxbKNFVRqZ7Kp87BSc9MesAhNtHONEusOOglmWZ5s8jsF6tClnXfo6rJO
3xJO+hyUWls559RHFhtBC1Ex+r7gKHB44gNKczI/8+KUd3C2cSihxZHthVgc
uWP6pfAjzwgxMVwDbkpHocYotExjKCHCFXRCGJWt/XQrXqGr0M4zUI0Oq1hy
nrZfWHFwm2PK6hPj/ZWfaNdjwJex6zs1gyqclAXMUR2jUQeXBFquvpQlB/HZ
TYxRCP5AvuUilr4udlL1qPt/0hf6hIj7VRlYrltVEKuN7TDNDzsVRGcGyIrL
gJUWA0m3OtNhIcVBFCOhrDA5Tb4xs5JCsafzNlkWfIMInLx8MADrm7Esv7Px
W4WQtMFVBU9USjO+SldR/2xph3Z/RF+USIGQtZBuTvDU3mNE4Bnl6+fxMLqJ
RXB+rb/LSUWhvny+kU9rw07v6Kj83P/vlzMdTju5Wq9x/JwewpvJcEVo6qfk
PEzHRX2Y+IM2NDyYuXPAVmlnibr4ivRrpd7hbsPkY4q6X+ZHD7IOHWT+UDiE
smAGwunDiWOFPfB9LomBmBhcZfMruubkd8gO4rKs2KZsgEelzodQ1HuictYc
Y3MOPAXVnbxGNG+mAYhzW4lLjFnxeKeGgMUaofayjWs29MqoIUQgA9hd+QkB
UskCY5hrNDc7sgmUciK+uv6Wa8aPsuRt6CbG5AR2jQM2/tbQugqJBBnVM/yN
QWk8h+EfmJSmNTDF3IrcM8YTyOr+cWPFoQGDdLwUBA8QcQ2hjaPVtNSlmyES
T7hW362feeeuZ6o9nmLZdclf8QSe2FT7o2RPwCS9UKjt8dWUUgRvJjxfLZjE
V6tVVcMYDcY3lT6c6ndAIpl5Erp7xuO6pHsYjMnkyDirrPozmnQNf2oYdljH
grkB48AJNl/45mquqAggIudzUdLron1soZNeKwfXb18jBdoz/At+1kMDFL7+
jc4jypUVWePOtM8MO8KIiG2B4l88cQEwwgONUozojCLEMcpxqEdrL8qhZP6u
fzM1B/IAY4GB5S2ZQlHJox0JCsyOiv5hLAe+tJaYS1JgNtdFKVMWPw7FRhJS
DLuNCww8UXYPcAGaT3XOWt1/7KOZomLuNqp01QIX/jaihMWFkCGe5ksw6XQC
i+w6ejIJ/Wm7XZTiccfCLJdyKXgCEtmr4rPPYpEuPDk9PtNyEzBkWegCZEE9
bAcvg7I5PbkucYhhjrfJslAT6cJE15K3G4dlOLt8MEXdPKFNLYi4vBKrgbXM
+lNK4pEXKMfPFYQ9JguErRopykd0/JfN00AfTXu+GiR85UqHF4LoD0mZwKi6
pZT1qiUNom4Zx77i0Z2TvSZHqk3fQL9rsLxG2RLnmZlNqw/NDat/Qe9geXrB
O1T7BdL9hMm1MARoF2J2DSW2Bpuwx3UBOS4S3Y8kHo78V42Xpe+2zbk7h6UH
HwhjdAtY2lz0ySj7xXd1lGKsnAWpdvnrfDIhs7/Y6y15A3TXgEg704WnZdyi
t2KNYomK5bU3FRNO+saYJkLDeQkD8H1qcli9MvXiS0Q0DxRMOvn9IjZd2qkG
GgYn5jQ8+R2zKrbFwFADhQ1PZC1mEwxfYmqFUeNN0XU1JkV9/9KhTjUHQGWh
9jqDVosVYZeC/kZKtOcmrPDSoPTj8xNIJnK0HbvbrC+payg+ZFMVhMiI7r5S
jXGGtwOxCfb8Uy+HyrM73CwSXGZEQ3kPt0FBgad8qCYoQctaFPDD8yLHjJbD
yCbh59y+EBBMTcc4wMJ7Q2w2Clvy5cMONdpryZ/OA3ACWOdMp2xxdWr7l9Oy
8juZtSkjeLA6XaG6JKg4dIJR15AqFF2A5QFGAdgVdG0fObKJnLWTrSyZ7nTS
PRxl1Hr5aKg9mYihPpQ2/1tDH1seUtcdUDFuttpI2CrnM09G2dSC9MAM2+xC
9pFcMPlc51YgrtME+X5+/UGhPYTv6Qc1G5aNwNJ2xNBUFicTvYCh0wSFGJ4u
IaRCCcDM8ZrbmQIDPbiV3lXrfDRMvY8kx5McGRSM7+CDW8H6LcRAaXe8TwU5
bRjcbUAyg9I5Q1tZ5A5p3B+qcgnimOwG2vxwgX/dJ+0K29Whe53Egyz4wtOu
Ec6KyrvOLGoFsANfN16C+DwGczx4ayXJDM4W/fPIE/HtbvfoI1MFIg5bbWkx
SBxvc5JpstYwVAbcr9OIKP+odOcmdzr4/O6rCuLEc9NUoikAy4ljPbx97Qif
xUmXSW7QrxRkDsNFdq0lcYpnUJstVWnfe59EByYd0k7xGY/N8SEqm0U1F5jU
gcOVz8xHbNbr78MoiGc3+QshXqVXiAXPXW6AZ0J4Dv6YADFJWBuW5kH4VnmG
JXktF7PTA5wy5HhFVJZvtXIH4Uthc4LcIkSrlC4YwRA80HUfrfK4YUCQnfMS
HTXNA3CPaFzuouDwGqy2yKyG/z8UOqOndhr2C0RiTdVUA5XtEGl4ZnEXEnU6
t2kCuImdOSI3WAT4ADK20AzwKILe/ncWng5Bu4Q4J9iyKaZqhUBJisgHBpwH
nPYCvfHATVZcKdgu5HHLpFGmKDsFjy0ZexTE6c5D9AZ71/sexIufO4WSTaXu
X+DF8tHs4IK1WjGtUMmhSCreLa1mM2LEUB4AayFmaKyRL6XH9xhMmEaWQRUs
GJXqBbSpNfD/zSHXl+JP9MsY22UEb8J400TdnvreBOAkZebngtBhOESL90Mo
tJfqwk9XVvabFZ4uVyRUh2H46pwMvbLjg44i+lqPJa1Kiuqlzvu89gqErQn1
BNxX/GP2QQ2ZYBMe0REK9v/UvYkt1K0ENRXN96n4QYPOvsAnJs8Ophtapmub
whY1wJzvlOhs73hxfTmaLeK1O5TvvmroLaU1UTaSn0pSXdE4s3z2mYLjK1nG
C133H8drOCgiXekxSIM4C/bDFkQoBCAehStnJ7zAUvY/0ug1t0zsSnnLZ6LH
X3XhwRhR+F+tZ+muwr1Jh8zmCyjVkoN9aiet1AjnMAm8Tb/mV+K1ral+16Hn
SlONwlSXCzkmDacOxXMfzLuD5EAh9HGnlx6Re8D2BzVWQxNOSmPPXjM5nWzF
mlMabkrwq7i8DD524HX1Hrkc+rDS45gWNmeVahke9eHgWot8BYPCfl/MIq8R
jjT2LLe+2yDcvceQcpDIA0ybaWVQJmGXXP4vkvi/wBrV3RIY2N8aGK1TGd66
sG4d0m3cUMdwmHtbvpjYxJWeTnT8R4zmkWvU3h5p2OOFeHxVa2D/7JGwF0HV
dlaMzbEXoi4bXUrYgutqBphPX7ExqCJXdWobTbCg38EliV92FLGq4T4i0MxW
i7KQm2Z9WdaIsYliDgZFZiasAtrz/gExEpP2Tk0Px+YsGXX6uqyoBvUgWBl5
h30r80isa05Meq1/oPerqU8EBDZwrwHHtx7r2I4nibA3aamXHPmU2YgvsLrC
5X+euJnrI2Utgypbim67LC8Vq0xMQ7VJP9CFk6DjhFqnv547EyXq3Qq2Vptj
OlR6TFs1xCFg1MxNYYmSgItmtLaeJRKE02Yf0ejsg++e8s2l3/j9KcAQP6Lq
FhPG0jYT6oQpEsOfdwUJlkuJADrC6pnYaUFYqsq/9KEuyrEMNYh2gkurrdgm
biOnw4/JwcYS0f6n9VFGYb+fNfK2oAY36SYAzeHBCSy+5JfyXYslF4QQgy5q
Pyc1zsmS2Thfh8vjC7gD9FlMxARKhpzlYskC+n7cy0K7w2jI7fhFHKdJh3C/
DmU8u0XJ+Rbml7ki/QO6Ochwbdo5jxaS2MvUPI9yJajAcLHZfLWhTcxVuRwn
5UJxqS2UvTEWLjveQ2owWZPPnQVVG3RC/Py9YRIGengqDxggp4V2/aMZbz3K
82pukw1nVWUL06zoBuG37tP9271cWdXJwVnSHH2qihMHQUqCTY+fzHraEZSD
K9u+kTzXxdvXfRgRVaLgSHG8eEPme+IYandNsaxKXcsRG8xzdIvI+ZtRy7iT
eLIREFSzBK+U9weQQIPAsngzZX6JQCrKVQ984UNQhbIMGyTGJoZEb/7gKs33
j1Xp4ZpHyQur1L+1UfNA8/GmGfYpIla3v3pwKa9kEM6zBnWE1a9ZHsy/eOxK
7DVADD9LyFnqE5liZoeJ6Y73sFnQHvZPe295S/BiBLhsRm05PdJEbA8UrU9Z
jcgdjqZmGd0qw69sY0CqLCU5Mcea4YcM/ylufNfbYHGzquxJqG9/xBC406Fb
H66rb54PTRqpiuNX5v6JhztMv61xGwedt410k583eIxmSVtp08oJRiSHwCRu
xxU/9UipTMeX8AjI7du/QDVRakV/zZoQ0lVb3faW9c2aWGIGJfLvCWBm51Ju
fCZJO+MfKLAMHTtB5FK2W+dtpLJmS1K2TBCB8YJmhXenB8TmnwmIOu/4h5GR
iYwgZMfXdjmI95R6Ytzg1qpjuZTBRkcagDuuZLEMF+LbantX06oMDOUfu7Ca
tPENnIvPcjvF/n2U49iTMkyh4/RqRhJjocELnsTtR6OWz7SpmcLQVvwuffvX
ckTZUC3AgqGguiSB1pN43XKzBAHb6dIcmikmGI08DGlKdgKlbMGQoo6Hi9L+
RSK2zqUYREoXuILUD7jPgidmQGa3xUUZGjCAeT7JxggzUZQUM93IRD9Wk5O6
gE3mV6+vKejng9k93kqPU84LGLjBRvA/qbnSx+KB4Uz7Jx0qWReKmFRhVcNu
HAqsYDxeagrT8vmkX3ZzQWgbuWM7W0vKw7R9TQA2NChhzejWare5XkhOKNjI
qCiGKEiXtuCzKtxUJvwImlq1jp+1LBJACHon+ZguQ1jMXAN+CzdXFD0a+7v7
3pQFCbf+5kba5TjTQBx1vrYz18wXzyQBTwN2SoUde5aPf4nf+NHvuVJsBhw0
Dp2qj+KThBfQcPAtGy4i//Gs5UnO7s6W3xFoQT8KXAKbYnF5M1jAtqGQCc70
g8UDzrhpkHXiCK7vbjjWOKtZxfiYV8ZHovTw29OQ2l7pCb7RwDb94nm+q4G6
bVMxl5gZUff0+lbU9kWE+jDTTTlyOkbQGnVNYCn+/gIF9A5StQ6aeXZhsgc0
z9VaMGhoYK8oBotjsGJaKAyH6SS4MDqa2sXICX9wIfmi2xiArUBbtBP4cfzH
1po4KwvN4qbEP5T71oar7rVbZuiANrGqknMvzJ5g5xbMvmTul4fIAmvPrqQq
cxxfEBCWIJuoKE+NWInQ/sB3MAbKTXtJRcJC6T+f2L+e/Oa4TGwTKcsLPyPT
c9IWZA9+hNB7x5khYHY5tkRxPnF21WyK0H6wSTBoepJ4OqfBgu8eb1Lb7For
C1ddglxz7WLpwQdpxYeVG6TgRC0Ydv2S1sSM6HF5WjZVAfsUk3zJw9wC2S9V
X53FqxUWXMq0NUSP4gpakrvSVKdahvxT9345+Kjtn4q3CI7FlAylBW/9pec1
CiS+gkb1B+BZrAQ4IVJMyFp+s2ROCW5Fc6t+RSGXzrm08iomd2loss2Jw94R
EZ9TT8BzOUoJxd9m9/BZrCZ2RapinDlsBaWaqDMZzbla3yvkduB5RxVkDRhj
B83OKMbWEKl195ivxFSe2mV67qrhQk6TFmm8q7WPGNeDmDRR9qRqDR/dTzYn
SVK9lF5wSXHQd15lx/iaRvlDJ/vq5426kNXMoF7Rq9zm6tlLZlDyg5S0cfQ9
MwdFklx+63AivSIcw0nPgI+0TJCMw+2k13nz6U6Yb+8J6ems02MQ/rqhX7hb
qgFxwRE6Y7hjyvFlH8xobyH+tff7YG0IKqgmUOiIZr7YqDHlXw8ApzTSF3SX
Akm4HxPNH0gs+IgoUVq3rqgPDhcYdYPEjjFbEQKMc5NLC5DuoYybfTX20gof
JVYm1tBtBNOOv9CI7I2zhCDEFqpnIK5FxIdMGr396dOlxEvZ0vSslHhx6JEs
QHSUcWVUpeXhcjz5EpvZBt38x+8XPQZG/RDYI4VA33/4PQNaeyO8bVdnx5ub
Gf4qHbzISBRhsBTWl4w6WTkNWTnTUowKyFO2ipuNV5aQPXQJ5XPyBQVAFSvL
NpeSWI62YCaNC4C3ImKXtZzyUlomdOcS0t9UBSpxTJOIVRrjjWZsg0MSN78i
eDYCjkKkB7nkUxlPl9mZS7OvMteq4wmhAnmpDgMxErDfDJTkggdInan1hAYQ
MT9cNq4W1hHUfH6O2MymxFDhwJkNNiqSl/1kAu3sQltihkJmofdwI9TmWi43
gzjRL8Nc1egEEhWoeXHkEHmUkbBLWA3fGuAau0kxwgXPwjKQFHdwpkWOnGtY
+WvVYpvz+u6Jnp+qZxgQtZntks6vIiYNVmgWj36cLZ7lwZQndMQ82DLsX2RT
aqc+izryDlcfeE3sIqZf4/EivIwTL1dQnHwqqToER1pMhSk1dWPVITdNuy4t
YGG5GfwGssTgcjkfaMF81q5GZSrKKz6XNOLdIv82lp4kHxuxOm54UHzmrKDo
Qdq3umHMbtFgEBqPnYFmN+kwHiKNuJuJ2IpD03VnIKqYsF/EHMLwfXgDkP5G
kSf7+6/vJg/KvlMcWOV88yISObLhoChR1xP/mwcZvmIbHXnMSGBJALkhCN+i
PDKnuTjAaoUHQ1BNVOlowaZxktm8Jx1Yx7+4RcMj3xp/c2fIEa9jkm8Vtnsv
fGK+P2KaHMQ5oDFAWhiJPh3ns6V9y+noa6uSTs83gmaZkr3VL91jeZFKelH7
Exi9qj79OdJYH5Cfmm7oT8tLMTP5FV70PgrKG3o8kAlanitHwPRi0UcfA8kn
JKaAyCWLYhSLeiUBKxfGXIu7TSH9iDVXaYOsbIda9rJrOPw4x5LGEkNR+7zE
NuASTDbAydN5nAolPoLvyTaqZO+GrUM9zo/8sWjGtJQX/15x9nvIZuI/I+/V
pS6IaeO2vho/XENcQdwlmRxOpI54OH//C9mAmDnq5W6bPxSUBDRXngc18wk+
HQhBXdniHg7Q3J5RZm8LaHC8zpcn91spRdO1/+uMbUQ3wiGaaqIG2lWMa+Px
fc1CWpQG8yxPsYPbd4yyqf8gCaxWVGplJTXuA12g5xhPMsmsDKQHGHHi6VBx
q64FWBuGFitOs7+c+H2LwMH5MQ1rg9jpwy4XUNRhZHdjtCrIMTPM2nBoms4C
yS8QQ9z5651dXY4r0TaQ5tb5GWLfhYBoSD8ap62pf2cClP1qF7WF5+K1KI69
XcYK+mQP9tdJthcwUsFhqahs8jkLtnyxdwuQOhfNMVwfyKc1+1sr3azhVP5O
Ocb3TXvkLhLX0z+a1afVsld+0jq3rrEPrkvo4NykXr2TdXJPf+JaU3NKk1pT
o2e4QmJexk00J2yxTRPPF0cUwPFl1pNjjXynHzwANFFxG4MmH3kRlGiBmOYp
N76GqmBxhXTlkRVnjyStIPfaQgwtzQVm7cQAQ5RB6DE0odqu4hpZGy+1stCk
4f9icutMPopYFYfqQP4vnaZZj4QswraSvfLTm+WjjZa7tIY/xODWPEl6ESHY
uhcyxyw6oZh1EWw1uyjgM6yPvZEnYynwn6I2uHV4pYVv0EEGzjMgwEj5rbqN
2qcozY79sOj7jVGEhxEmmpvNfVD9DH/C4gUknDv4b527Ov6cpwYI5uO0hv4J
UJdL4FPWICWyG3q/02aZAwXu6P3FXjdHGdFo0InD9TCe44IPAotyBufNpMfZ
KapjE2yqNtOnbwGJvU9LOk2uFLggZXLAUgdUjnghDApq7OGZKW+yYAGYu1x3
LuKrY1bBXcH9w4ykVfU7lZvSGHDMTRuG/JP3ekBUPQZuuQVOle33s3CHHL9x
JFNcQep8hfcfP9LO38zJ/hqpPuTn0uM7TLS9uZY/3Hj8QMuUPw8IisNK7eo+
6NkwmBuobD8nEvUa5Bk3zG/4enUiubul0Pfg9Pt69XUjPTyVHnbTpUV0+9+l
oolJJMUPK5ZRpwyUSzNCJOAywx2ObM1gmwS5FOqYP7TTlpcL3QDoJCNPoTXA
rTadMIurfzCUFnGjkyBYo/vvtA+QT5MwodOWGptAPAyyZW4Kv+uG9zWjf/Hm
r8nb+eT9O7M+gXOWLDg66chFPMJgBHavtX/QByD93UXvNhtNPNuTedoR8K7E
ahWcBkzxz7Aos7fbMK6z+GiJ3nm6LPdd3Y/Hp5MlPki0elHaVpKpN/TGlMbf
xl3Ov7Cktl/Do7Svm9LSgkU4Lnck4n+a/m4ExuO/8xxM/zrhTK61xTsRZXHr
G+ylL5o9pKGSSDj+ls59jWIBi6qH0vBkQCWJvFRq+O0gUli6W3KCnbJ0x1uI
7SZ9yXc1tr+UZ5jMx6umskQzYnA5mZIgHyYVEFAJDtQcyQza19F8lMp/h8R9
D5BrMpDZua4DeoY46/OC4ZIzSd0QEMoI+fuu/aLjG54gCv70WGb3KoZfJqf9
+g76qdGGSgdxtsW348Vd0OAucXjciml4aFxSmxWOILurD0uD3JUsPplA6k19
uG6dvCQgVszV/qlLxZ94ZiEVTT7S7oalTeQ5vrIT2Pr/XK/T8aEZ0OUYp3jJ
ulISrVQt8+O2LJEaL8Nvzs7fGmq2fdaPgXiSettQMQOeuHnRgzD58olGk8fj
5hAQhgxgvqutPo9j7GboblQtVfNrl/tDpXctXARMo40WiYPig/9ZZjsfcq4E
BrL0uLRk1XT0kiKFVp6HsED7bFwqcQBNG35WUdM11yEv7NkPFn7fmcIFHNih
s29K48CSvNWu6tvba1A4z7g7tjZ7ufCRr0CYLZM53huJZPzeng1E5+wjpZD7
40bcvSp70kqnNG6+UhwXHXTsKxYxHb0byRgaKzvXLTzcRQu7Sg1K9Sq/DFY1
mPdtP16Udwu0xTAWg41bPUtkpXV3FgIB0XEzQg0YkrytTI1MDJQgNM0OxnYm
QcgwRtuO53xCzjqrPwAU2fAgm4eSC62NxGoPbJq6F/DYJTFbsdtFdZp3Md0z
z4d61mwzgx3hgF+cQML3pXeolLSizdlEtyhVUlsq14++8RD/ls11f0x0b3A4
SzZbHAlnQO6+YOBOtPUiYgr/+q/UBHZ6xrKgxhMecaWDOKasHT1TlVZGYWMJ
sUBtBKKE51NkRE1BXxfUNRs3fKShXZ/ADpIAjFV+wdSJioJAUSaN5iHAbuWP
GYIFQVl4GfiDsm2TGejZt+73Fm3jcMhjNz8nWdSd0RLFtkgnrbKfvr7uegii
atdC+AImm5fFKIANCd01l/WNnlGsYGT19pqfuIVk0kfNj7Ek18Wdo3fpslB6
uN3IpFX4fX/cs2qKIxtryFnfqgs3lKXdFsxpEC6ohd0jalgFeDNpEwUeLBBZ
S48vWZWU9YuFEpPPEptGpu5V9u85itbHgPJdKROoKJnNla0SNfSkpGUyTzYo
TIEXtuTTKYN56kwt2iywrLJVEyc/zDC9YgFnN1vj32+iUYAe/FH7Qgi+WIIx
ikQaoJBW6zZ01iThvQcY5uRJjoRQdlVu0zeFnN9X7+prDkFeDY56pWtBuUTg
eXSS5um7lapSJi7U1Hb156t/weDFpedJF61yxI9l2e9Gl1XRVWI47rB+abBI
yfu4swteYjMV53clTm2SjL8MuPFJEVBeCLpEqtK2/yNqcvxNeJ0P6yQ2v3Ff
xgOJ/FpG1DRZGvnu73PB2blD6LVipyHOAS753Sfc3e7BNRvrL82nEHIT06kk
XAAyApemoup6w7hiiZ8dw0yGXzVw2JTlwhwKn4Snf65BhABJ94o/xppczyJ/
J+ksQ6WcCJsWoKB8+CeZebqRal9uC/2dAF34yVsAKNVyHS6jJMg73seTy5wx
uXVUl3nLIMn1qxJacXeqW3k5mDfWERamz0mN2hxBKzz1zwlrju5IrZfUw+0j
XUMXPsVP60QJrDXtgYW4Y9q25Qxm7mIMvqyT1+i6zKxdpYg1TcR4/lK/pYtz
jxkUo39nR9NlT7veEJ+DY3iJTqLjKaLwHP6+0GWUVRwYL9VeAA7Hg51QRL6O
Q8b4T3lnISTclAdQLaeuyRwr+xHvsyiw6nwitL5y7swKdh8rPuXloYsOUQ7g
GszNTQ9OfqnNOfcmalsCqDlst4QXlTANNaO+v0sAYuddyctWaVFRqQ1iaODy
84lzCMdULuJTNv/l56jxnixKbZ5rFtZtOJ6NL0eShTqLCMotB2w0HFuYkmS2
9Eq34htodqW5+E5hUJmUcO/f4NtFlMLobpf5DXPqoNVjtMmYVWRuVHZiWDq6
80E6jkWwKrHxLHkjIQgoRSB+ehZ0eWdyknLW0hk+cWabqJYx2tMyKJm+hBs9
10cUD9UOSGGIjzGJqAcBnPZqqtcjrEKioyONNsHjO0ifIzoWcRMz7710a9jX
huSrO20Y8nTvMBgsl4ye3mcHRZ/54Ya2gQoGR+az56ZPPw9mrcBPhKdn2XBn
ruG9X/VpTC1EBGOtfXfu6CCpDHPMWSL6diagFENYzvffcg6eSxjRzWNRTCwv
avnX+HuPoH7X5cPn+mnSCBOKVsZGwx8LwZMCsuu4zFFnbxTmJ0KVbQXDX9jK
Qb34HO9CVE7PxcOdyUy270ujGPoFLhWkJmSI8BRV5aSC8/UUkaF6m+cdsOV6
XM43BFhPzz2qG+1waCVG553HkftrRfLEGSGO34ShZC3CzVNUOm12sUKUZQms
dAjFAAW1TUb69dZDnfI5YrKekOSXBtFDb/4NSfoSyaKSlUxyULit+kbxft79
O36pb2YnnYuku52HAxfKS06RCNOZurSTlOdF0XyQ6gf+njllvoyR/ZuxgbCs
x8tXh+qOGDdl1AZXk3qtD4jJgX9Px9YnSBEKqUU+KEHNL5u2arpMMyOd7eAc
fuNfTnDhZF9HhsvXFJ2PKuMHap6JhehT2tyjds4aa4xQABS18rhcUl540FVK
PCD63m2IjbKtHTsYQobXDFqXtahjn9NpCOOwXlbv52qYf+d7Ns8vWbHh8kjS
lDKiapQD9aYbYmUpaLuGzOsdtZnYhRVBP2brw34P7AW62igj9PZJ5yj8M11p
yLFAREs7bORwgOn9eJeU/Dkegr66LrBADBWlnaimZzGCgH5yT0YCsjP4C23L
G4SlgN6UJdXfM0h1/k388E1Z3RP0AVx2kqt2agOD9uo/0WLiNxad8fLH4Zv1
Sw3Qa1n2GR6eiGW228S2uJIqmYFqJxvZwGOpiOi9h/XmRPL8svmPwL6wnUaJ
Fxl8GIoQbC5/6vPV6eA/MArm1T5ucKSIUbh1ajWL+7NEhC8CJht6k1IvUWE/
+6YqZ5QsqLfwEpfE4RiDObnFW8W3ZJ2dOwETn6XsrUciYNZhZf4nIJJP4LEl
0W3fUOIIdoKCi0SoPmhI20EoBCMW7DBKaAX5dgLMc6iO/FMtJ80eaUCUFzxc
xnJFO6iRXHyfzD9U1C0C4HAimizjowB8n3sjKFYAErdmFfy4DkjFGL9EFFvE
Xqgrmo9cKgKmX4sL4F26qlBFeZUeC+I0VVK+tFt9g9MGl6LzD0+MG8uvRRc0
n5ke5cUrtUGhHUI2XhJ2lnFb8OqiXNrN0dIgbRshsrYzLvn3OkSAZsIqPgZj
aySnXV+rhpXQscN6vXHftkLxMQiBePHiyAH+Y2y/qFBmV4PAOFjTVqjYw/8H
uPy70UIEXNsdknGrteCtOOasufOh7L+UeLbtzCl9U+XmEJFO9RegojKP+0j6
8nnpoJ1D1Eij4VfqQpQRHcVoJLyHuNI+PJEeiFjRzJTH9JdwhwUM33xQfHLE
Kl60QwQf8oj8qs9bJg36F8jULkUpwsau9l3Xh+T+tb1kQgrHg1SZDQwsS9Z/
NlOXjskmu9bukkzomqmG5laT/PqMa+EuUtI7Uz2x5eNUdC+LNL1fsDunJySB
W07Nb8WTxOr++wvd67UA9Y1xhSm29hP80iys+Wdcg5LJibxOBs9SeQ1Zi0kI
ucEj7K/nnjYN+Dc8vNIaDsFisTTFlIlYcr41kBUpjGF99A2bH3r/sLlVQKPW
g/Q3bWqbmTNvyoMnPP8suiRCsDjrhACBaFZWyaYEj/P3PR9HRuLxHhPGhnWT
0F0fAMVrHxqnxguSMHB/vSdw2TK1Pm/auKriVQv7iELYgLY+8kyJ8mJTJ92s
0663Av3It/9E8xw/RO00mgbpq7HGVWya+LAgAYsZ/QUagLCp4O9JSrpFLP+A
wuaCtgQ5LvjXXi9wZITLjtDgPZRR43LAYsWGEmAzof4BbC9fHJKLVRcQq9MX
G+zf3lk96r8os6dU5LvBT7Lo3U6rsFvkvfuAOZ4njeey7eqZ5BHyrdIXft6N
gOVgYBnzTOiEe5AwqDkjmyyE6Gtqbm0KLKrl3ngEku3mXBH4yjcOY5DBqjB3
zEonO0Eqo2MhmkxXyRmbKoGUXtx/ldwO3TkKSTjIM9EaHfz5GK4kYpXgP01W
+xzucB0MA/c525Y7n+Y7/zS9YTwlPSeSKcZ79yYVOkc1qSnSST/tTHRjJWfc
CSGEe7BPtDLQpV3hgNeQwWbkX38R0Kp1A9BJR9L/VYTWVMlUYO+z1h13FmUy
7KgY9WX3bQhfaZByoiVLtNx8KQ34WREZs7niONlJBDLODhkQeULARcf0uXrI
gIin14ulCyGpJU2Xkhk2NUo83BBWpmLNmyhd5cwZRIjBapVV37e5qAFijywo
FdV/yUtimGZX4JCA+2HYh9q3w9b1md+0375SZ7uNSGajEIYTZAIIIJkO3xup
n+fHsfoWEj4Tb6AMYoRab7UBRk3HvoLpMyl5ULUbMOapsao9VBnAwXRD17/s
JypS88mHnetcoMz4YBh0cUlJ5UNKuBqRCx0xqmbK8MOP/5XdbtbukH04TlDF
ouWrJpoVd0NHE507cc8k71V1Eh48BROack95NpuuxRgXIqKkCwbuCJTEEp3w
BbOQlxHUwPwiqMmzUYi32np5AXthPvJbB2+AuHw3sYmscBaQ+r2cDD43XcOT
fsEOme/GSBxlQVq9YdfRIga8PvFfAJFE73+LLT8S8GmO9li/WwgdAlN6QU12
CI0CHx4HhZ1I8NrZtliMIC0+q668A64O4ztvllfsHUjL5jXTyjFVig80o9ZD
oopyub04Nvh1i5M7NH73SWzI2eQaNhFkIQt5UY/iPVBD2PfmQg9r8kPXcSdI
W/KUSuIvs6UYdMRg9pEQOW6yDyauJTra2jJcp5V8PJxjSdQTU4igTG4i/igg
tgm7fkISy8ZR7+isI7IiSqZ2J0mcSYtPoLwB83BDPfCbgXLTQl5l23HtIpIs
Sq8j64wl5lVh/XXdfjfsiwtMhAJD/hQbaDaMI/sFawDBLEykAWBTRJI/RNpv
fVtZ31OL+miHT4sw4hqNCv1eJ4vDEIINq52wk48KBWepLhOZihKXqKcfOJqR
9DccBsgmnltHmhHw7R/H3NLVjt571legfyZClzhCo2Xfpm6c5TjLDOMb496Z
KT5wnUnZTuJZTM8+An7UXhB9R9WvyTz0ZvPH4qQlLEpckM2qrZLCOeUBHNua
vnbTc1w7XL76cEO8x34SU8nwnOSyFH321M32KvSZ5Gqdfv8SbTYwTHuz2oQc
iXPr8b2afUNZE5X3aoCoSH+1LwOukQWPEowcKJ9y95aEIaXscV+eUY6oj9yD
s6pVYA/yFB1r5Hs+xfoFUtNMbqRVeJE5iU7jqdMwvL4ImJhCWxNRs9nX/YBd
+/MV66G/wgFK4+8mfiW30FR+uIop+dHFx+D0/CUqcWmVefHylSUqfaY6zXgg
ilURc0U3H+xjkgMFSWyoSSsbhgO/SE4q5s7/A9U5jMdlscmGsF2fqQgnzP1A
CBVAL81fYl50qZuCMJnU5qU6OD8PSFwd/kR/SEbboEoPS6RKm3s/K1inzfu+
ekwatHBh4p4U7kogxy83J3HnCHWHr/lNyinM/bW87jISJGG4x9juXoxLfm0D
fCpcg8DLQef7p1aqULuzTsvm0hXXFjNCEoOT5phCSM/5RI0eP77zfo0KRq1X
HOwo8fnAYT8bpFU37lvBVcNTYT9n8UJM983b2Hewj2/VrupSP+cXkYh/Dy8N
qHbEF2RSNIDwR0hwont5r1lfgwGPVhSib28AANCEMwOzxRatpApLrmfiY30o
u3lTy94BTRgBUPDwLCeIyZlfhxevd3ElRQ3Q+gz6mzuY1vh/Tku6QXBZGdr3
Gcm5PzVaVP2Iz+/7MrxikFpOHgaMM5LH6HmPZ2Gqh1TDETDF7voLCPeCqQ+R
DkN/ssUSVVtpYfwJNJuV8Ub60QDQI2PeLirqwTe9oNtiLWhW8zRmCWtK3sV/
o9+0Igimc13nVA6h0aFq/EWPe6MPIPz9LYcZ9FVXnBcfrxer43pPTeJ1pseN
altSFx/cETaqUn+1hUwTN+wosTKgE2Uvsp/bm2o2rydrO5czs/oN0KGGQHyF
GnCK7ZDnp8C04GLtTpDh5it3UVNcZSjTL3d7CV9DhKJRMW62nyIH2EMoB8Up
1QyTcE+4BLAJGjrhJQwWhSLEj7TUR2zR7hw7DCw4QPk3pbwCoCenrXeXb+RF
WPIGVesgl9ia0x/mG4qhu8rD2py/EtycDDCv7Rxt6LdD3AwdFF1CPRak691G
QGYFbo3yckop85spvLMXLjBdq+C6dlJxWx1aRHG07cZtWTC0P6iPJYJnueOV
cb/76B4n7SjptVi2mvGFWb29n+tw6KtGHsvYI1KT3cpCP0qg4X6TfSDqu8fh
KnuI+xq+oKogDmayrRkzJ7wpxAymRw+3UDLjHxFrkA0wH8wSv2GRFiEo69It
1zmJJ2DojNmlMS7DMw+R/0z24gdis844QH1t3L5Ix1w4vBEK0cPJcBBm92lr
AZuWwz2z7eGtHkKaRSVv/ezerkmjVubzch1wPcZ0ymLmLJ0tuXgV6udC16Dz
Y1c/lpEcgttavs/sw6+tJnn0q5ytkdFfRgCTDtGjpauWfXGW2B4Ab9kt4JKv
IXVNvODnowd8bV+d9uOji80ohiRAat9tLzalA9DMjQ2TYuxAWGa+HTibQrn7
e8OGmwjPoHYwwCyeK6Z8CK/2C9H6natdCEFQGF4ZXQaBJ3zClUJq6BusLVvU
JhQPxxkPeLTVM6ky4hhXbDvdwlZgUTWObOVPjiRCTrSsaBEvNwOITyAbN4EX
Q0yz89yodRL46aMKIfZ3+qbqzDLsQc7V7CVn6hbw757JIJP6wIZ3SSWe3qwJ
FZoGHEtAwpiGxql3GD0vLNyrgU7VnT1k6o2zD1sZWlC9Heiiy/4E0hzmDngK
EwpxIgPBWXuIwmL65CdOtW3bTbfkJWTwJ03MILtAV3thhW4PaDZC8AQCIj6O
br+hhRLhAKXxI0uF2vqjcZhiKjUZXCCcgyNVQ6RnczHbO/lbrYUc3jpxt1Mz
AodsqolLLCJd0urce6OfbI7f+geU5QXiuGAZs1Q92xp5GuGSeME1sAmBiFgg
4gzCb0QWwo0pAAWsOJ8SUBVE7wnqmG6v6iWEPGtr3tZIDxKk/lwspfyEousf
nQnAkhEQulCqhK6K1Q7MazY6jiwWbisxSqmW1XZi+wYRva7rbd9j9Q+STNJ1
JStzmt5oZvzmaS51VJtPyK0wSf0hKxnRiZfM8WwAWJwjoRltXCZC5Nlv4oAD
VkKkuCnaNRQQP4MAUGBem4OuuZjc/VnC8NmA1YSf9fZMHo5CEZ8y8btIXi8x
Vf42MCoAujTxnJjRhYEocR/soU3NEzG4ZUXKfcdUgm/iVcnmhKUPfrxzhl8A
VnmtNl7QJK2kBFizFQ+VP4eLM/ghJU9rCG0bj5xDrECRGN/lOWNtOh0u3c0M
zUzxWtyD4MTdw9xQlyzZU/4FWHrh68vn027fTUz/qYoVnMdRhLQ8u59jQ3c5
0Zs47U89XcJ2/xpByz1FP7Utu5O6WSTOVUhSz4WNPZ5GqXHhJhzcFkvPKoFk
B+jrFJXZE2+N8ckrPNcZ3EbjkJGzoWVYZOoTklXZc8PwpsndgUlw1QOh3PCa
lRJ6D5JC29JbAP4bEMMM1DyJfObO6tvFCZNXvncKZi3gkY5eJutYTzA1N/Gz
STRNzoajD8GqCEeZg8gmssU9l4js7gUL/aAuNCBi8gEop/Hsreuu9sUSRDaQ
5KYnKGXBGwLWGNVD0ON6VB3oZqoDDU6m2A9IZ5YNTHmSQp4/Nwd1OcZXsBDy
/tFvHHbb3rXpdLngneuK3ylyIk/qQBqG3lRg1gAXKNY1JBcaAkiu9WPkMq1a
VYERmso+x/AGWAIWYwuUO//SmZmBhLeXXaBRFigdWCFBiAboEt/wVf043KfT
lyDRjouSY2s9E/81fiGrgDnBH/3j5yZx+QsAwhIoSReoBQynPcqwAHH1AtV9
cjRdLr23ZFdt5g1Q6tJB2XJAJ2PBA16AnRX2ge/vvVw0N63no0/FzNhCYlsG
DbVgDby9bqLNvme5UNdqX54NmN4z5h131xR2G68KhwnJ13MdDX1RSymQ2+aX
OA42ejje+ZoHqmaXgX7GVFEyz6xMfDy+tkh7TUYixS/PwGisZ8Y/pxu7519W
6LE0eHNHYjYGlNlYAK6XW+Wh3hM4eFfAhavpfVG7jNN79ySFsgb/LP8c16X4
LPZpqdjkFZGulcEF4YgJqIp/uNzr9rUg35P6Xf71F1oJI0QfyxL9SCzIK4TY
nrxe77iBhhmfaJGBe4F6YcDsdq4FzO8clWnPMwbFJjKwk2aWCtvAE4W13/lQ
k9t0CCg6eY2qNYeAn/FxSMclDqXZkDGbbjIwMJv4qoKe2xQGuvCVW9FDgO7P
4kotzYxIer51GiTsKiRZmTf1iRzwwGkjv1cKrBC3c8HP5p9ghA28em2jAw44
BAylBbdsxEZsoPajhbJIgMfUHDvPOM0sWJuxnu8j9309/cI7JoDM3RDR97Bh
3Mmap972Aq6gMJAI8JJDXwdHArfImJSu1O9xgFvUNEO4GPiSFRpK6t5K6bIk
LLZNiCrspN6j6Qkd7cDeLhAjnGlaKUCTt4AkFYpfJZg98VhCW6fnEVIPVYIb
Ia0jx7j0Qur0OIp3a/XVtr73IBtBBfRKwYsBR/T5iurtfx5zZDrxYu1Gvzh3
8QvdR57k0Fn8SdIf/2e9dBvM15Em9BL4OeHjkL7oxoW51FOVSP1rwdVVCf/j
TdO48dOj6ly2E06llhea+n4q2zXwGy+0Ohmc/370Jak3IJYYfHOp54hvYsyb
Us1feA5tDAYVXcKgKa2dG9WolsudGbSSCqC8Nsr+t4yEEC6KCP9f4aZ3mx+E
gWbfQnX8atjs0ct+WghRCkoEjmOJG4QKQgPunoRHeX/co7g1EfZNf+/H+8fe
8AijkkRKee5UrByXEfRpt6vYEkmlox+MX5nEAkxYPHQir0pr3Udo64qU8Xzy
2+nvRtopB/F2r18Qttq4ru+uU7zE5H0YCOfCu6xq/ZIPKuAo3qsyo6nuhzNG
7dxmMcBI5eLVHHO24a6oiCD4fgSz7KetRnPUQks4UoCT+Z1G+dze2ckYR/xl
rpujlAWxDojPPg/2cKhpWFUzLYHKnW2A7toisosQ8Xrg8zPg23fEThGXGXIE
i4cYaTWjOytP7p+5IQEcALADzeResYQHOHiCHHsgBugstSpvxgRKDux/Q9C+
YQgVQ9q9h69ZO3XdCbrlRh4p9DvHlf0kEnwSqnWaVz9NP5GyTNahMV11uBKA
wwqFtiLXoZqscG+wQSQ6W0qXIyW3MtLZEeunxsMopywOFgDh+9bcUduViBG3
bZYlNBb+XG2guRVA0z9i1tReyGwY4rsY/LNnkKELIyiKqHTorKRgQqP8piNr
FA3oPyP7vQCaDJbujXCaY1nXT3CudNsEWEpOzQq3sfNyP68SA/8efiqBj2+8
J7JH8G1sWBcnuOz9a92KWZ0mTVnOHMvFTnubg1/Agmk4jSwzVZA08DQw8VLj
NLsbYbpTSxBDaY0Dw1u+DC9og1VhJJx2QOJU191nE1Jbs7FQk8hWP0DiMV25
3go0o3F7bOISx2NAMYasGt97Yse1Ug6Kr/bC6olMtFleQMr1XE6ewJrxdq/A
49DcsdNMbYD1RrsNdJ1g5P87M3teDFa4Z0SAxn6BYqk56Taiztohvq6m4RvX
KVCAm3/pGl7QYxPdDRk1nRbM+G1VbkpSEAOuQLCEWaaK0aBgulNfrD+8mbGm
WXDqxqnRjLaZRYT8sVpUQU5AzH6wTcDcSK5hQcQuz3KngA/J58Qbz+ffSJUK
DEHaVqM219CxiwBB3Hm472d26R6lCLLxyZSLffcZJOfJoHcmw9VmByCgSJSO
Cz6FZpsllzsgo1w2kbA58EY8jtqjs/eDzTx03JcbYkreZG/Ke0imMNFtaacn
wXOgedkMYmaJgqPRLZLAY+MnzohYod0EpZGp6EMfrNsppQv+bpPNRQbSAwCr
d8EMo2GMHzbgY6X6KvdHquFe9oVKHn93KHEoPK+EkEbsrj71WSSJx9o/iu2n
OGUQByr441BCBuAD5PsHI2xPPbmolOEj8HEjEsk3+6S+rWixMa1TEL4dFeV4
dkUkHSDjk8y6oVPiqU0/1K0tm3ZEt9+sCnLjLmLID8WbEb9aaTXILrgiRwwT
pi0VI3cLVoEV1nuw9Onq0Z+OhCavRPWTgg7t21iDAwixuTBuMFi2fMHC23S8
tzMmYv9HagNkNcb+vRQxBNqdYV3Xo29ZWNpughl9/X1eApYOa5N8ohxnLxzK
55ww9BdrMgS2DeOyjjxDXaWZiQ/mYbAzyZQjcg9J+g7xmFYKI5j5U+XIuLhs
LdgOiBsljtHeElXjqeoHaFKLGAFTa8yG8J6NOeRN4bhlLp8ID9emUL6OEY9s
oCqdR4yNdjUC8krPzF+Eh2qM/zg7/RlrJ8w3lcXQgIlE7saSg+Be5oCTeBYR
Y0EQqJR8MYmVWTeRq9oaq2fiIuisX0CQbvWdUZpSWozXg/0bZ+9Xt4UvHsrJ
KJLcYpI8yD/MogbVDSawNJeWJ+rkH/Kpy+tXFlBg/I+J5sHQ/rZ+KZNfAIh7
E/qj8meKEyR+97q674cwJ1s5FmY3y+kL2oSebo3boLhPZ9frwwv3PLkeFws3
ObZV3Bkje92Khl2hOjPsg5Ip2x0xyxZRqVFAGV3CqyqaUfxJYvIYLmOZl2Fa
Cb5QsIh46xjZwQDX37q5IFGTx35aGLHD65libwHghT7F78gfp83pnwLBbKXZ
jXC2g9bJUZk84mphAsxNqxktackEQMXw64LkTElFQpQGAoQivb+44cvTiKqa
IxeM4bsDlWSeD/8gLddcFTMtue/upVeOmHFAgmtf8gCh73EoKhGnJUhSP9/g
dpqbk1TZES94zKOUHfqYaLH1iKSvZnmcOZ0nf6KVXM/FeVt7tbl/u1yGnGKf
/4fyFj7Y+5l3WzwGrWevrWBRF53AJb4czO0yGMpk5duL5qjsb039alt2NrFj
UAv0LVO68Zbpp5erTSiGv05DBNs02qw0j/y8dqdznhjEVaNZ9Xvzfyu7zOwv
TsiVVsMAaKsXNiedFItXRl8sXpHY9sxN/lj5zGtUaBBGmDnyzJ6biPjdBJMC
hlyFtatr7eF7H10kYL0BMUUmAPY4F4/17THoA6+q9Co5SG2stiRC9VTOZ4Bx
40EiCI0ZkDKyncnaEfwp1Ic/Y31mOIRpD9G6lrbttDWjrjWQVaVV3sHjfIPZ
e2JC7IyhLiQiCgWSGWEkbpOnkz/NFzHk60qAUJUC3mUebjVi8TOqwt6FLKTg
JZRy/+H8B9jWFzHlbIOqMydenWdLW5Il+zZIcf1pc8WzJ8wLJBHZWL8wS++i
zTP+XhTD50OEOo1xo0Ck2j1wpVbunxJe6QBaX97eqe3282OUxO0N9Q6Is2Xu
P44fJ1ShKPAvdxJT7c1uOZLMuwGmSKFToLbfGRWF/P1cc9Ee+uuTIuk3+vW+
BbMnnSniQ+knQ23aLeGbdOPr/43K2q76tVLpCxKtRtqV4uJFimYY4a/ees9m
gKT/X12IUHebgzOQuDuYeXGWjaVJEwqGhZCn+EqDenoS9e/QM+b9+RR2YXTD
rUBpyFl+uy/SKXGhOMggq7+MqVPMtEwhvf6a9yaqaomGsxjnM0bqO+9yFCpw
HaILCFfkBunp++U+9zOWehUsDGlXWk/s3xsh4Jak7SGOKvivVF9YBn+xSAFS
US9Vz3CsK1SsWuzMPKt3KRoix4WCEG5fck5R+Ij1EInd9TqWluFemHSBHva/
qaOq9ZgE0z+r+Dh0DVB6Zq5eJV++C7xNzkjeiqcjvxgXG1FDyeeVNNFPyxw3
OSLrVY92VUenmkDPi3aC8cZ/3H/nSxhZNipGsUXQY2MC6D03ei/mUni7rLTi
i/H2i+QiBcmsLbqCo68xMCPWVTa9y60O3dl3AHY+g9UisgHRfkPyr1K3FJ+J
Usg2oEpSr1xjBs4NAEu+PnCUVM9wy7sOSNKNJJGVsuiWqpnLATAfMAb/dLpV
lutrKGKQiJtdImoIWOZUf9TZNbc39PWuUi09XZA+LYnsJRBna64Pk/EobES1
rzuhsczu4QvI3i4m0T123UKC4w8hS33vaxzw9UDdhwCuagW595LZWX/uwJAC
elma98Sq6yFIqTMAQL5Q17RYyVw0ZL48QVDyLQsIoofXKXwgu4XdpNJsI21B
NWGoh5YUeF5pHWOrCF+P4/JE//J0UFoInARjm3gP3WNoSlZ/VC4lwn+1J716
plHEPYtVVbL+TcdyBYZbz8l3w67jzwAyi9NW6s8MeMnqoR7YqEU9XCcMwj6U
8HW+stvA39cnuSNzFeNdd6/8nE4y8GGG1kuC3V2CSn6SKxqseDMSdQrbn/cb
cAZj1niWMj+dq1qgcYneu11lvbB1cu9AGNUUofEtCpfQWJdxTtiDaTpFeaHV
7GkFR9XZcGcpxuUMW8TE8QAqY3Udde3yNvlF5KJ/jnjEDq6Nkdtz6GtCuaJ4
6rfaxrlGe3AiH3xfL+HKv9eocZJpJvHAVbc/fAqkpG5LiLrJfSerMBTLLPst
lqlI2r477eVdT0P9eHkDBr9tbEL0U1FIrB6B7mz7S48XGUw9frJNLAaz3uTW
7hxcwqeKGxH86kSU+GZAsCOisDwahNB4fj3PyeX3HzfSg7S5BnhOGqTDQCg9
FfFt+W94Iv6SOoOZajjQ4/OYdQ3y/nknvikOqo+qKKPDsKILO5/JIe0fCqjz
R17887PvYb3IbdPV2f7LgfluVsCfUlj7Kbi6doRRfDYYmN+95xtn7ifqUoLV
nykg4o6mcZzoaAqo9/Nu0DNVzz+5f2jdO0IClhuqNYX08nyQ7IRLCnAxqKUN
BUn3KoGQIHRDakLwX8FMM+HHyhY9J362Ar2JdkR/7f0rhPh1+tD75urt0Gj+
RNy4WrE+feccP0fwD5gjI5xjMxmQRvQwcxkqrkW+pH3fzzC9NrPmrxHK0NJ9
hCusKw+cIIu/dXw9aqH2OiUzpdG4AiDLpVwzIDZPZRiesX3bIgfM0Xv3XcAD
wvz93RL3QP0ktFzvnuVv3Uefw14CfBssbavLDLIK6KnV5rc+ggCLIIncu/LW
WeCHs4dYtSJEv9q3J1ROELDVHkBPUDwIqfoU9DfNQEUWCO/Ti9Fb1vQ1gLfH
qix0E4wP/JC869cNsGZCw2f4elYuoTELkfWgH5i3UzLJGs051Ag3C9LYEwvt
hFtVr3ovHzHj31cXz1BvsFFRWt0fHfozRcywlHsC3qj3J3O+8YUYSGfYN9x5
eGd7hKSGbC0J+ZyRAiACyd+h0BeN1DIKd9Zj3bYz94baFS16tSHp1jKx3vNU
mRGDLfxYNsuxqkOmoQfpQWAdoNr2gPAhZngsp61tWueD84jX/Tu9gzy4AEKm
v3j1brLs1VfS7o9qSDGXj2WWaklXODckGLbn4jzL4ox87m4soTNL83NVXHhA
LiwdKHYJYB/2UsNG0jOlHLOCRlH5rWOE+fbWgiMiQDXpgAUxSlKWCofjK/ny
VUPbaKhD8OxwpSZoABN5tJ/fO+TCylNqVzRz38+Z0QMuGtdZDJil/8iZXN6C
onoQEHqyDqtYWx7qu4NI6DClV+u5RbePV0R/ijNx8J7JITZqCfqhrJ1mbQ4/
JYaEFUMcvM9IysZKorPEZ8dCSoL8F7OG9I62utlPfB3y+bltdMR4Jjkdo4SE
f8DSzfIc12C0q8OushD3ZcvjRM5uCa2bRdisldmJcAkdTWgakzXiSEd8ZPse
0GulFG2CiUwQjxX/uZ7ptuMkgFLbiAWrL5LnaFbSngcUjNwp78ByOw8kNwJG
nOAnV+RIKrpi1hJ4mInNnRRJEYCRkVmz/IsUSTFcZ7+3MekqAfQXIP7ZVamQ
VUcLbTgGYmWnCPm/DnNrCfcYYUfRFNzG5qMCPvwRE4T/f6rMugyNqXHz97RH
HsTA7EDL5PY+KB6iEDTC5IvIckZvd7QOTB7AG6g5z5vSG+cHrAFjiJK1ypeI
KJuJvTX/p3WTkogSCYYXQ3BKQ2thiG++dq6qmAxvaIfftRIQ5rsMaDxb4gp/
eqBSTwiXuwQ0nWBt0C6JipSSMSa2ifStmqzbEvrbtfnjUeqg7U7ZlOQurtlX
zk0xScpVSGLkyBeZjNITxh6qKNLwVSQkcN8wovkdL5f5FxQDSOMS8SIs8MTG
4tsElL9XYvl3uXSBjwwVXAoIR5y7xLtNfK1nQoQSQnctoHBAT04Ah74NluKO
EW7WDYDJPJSSgGY3bR3fRGUPDWQBgTLnEra0+MbToCfBqg4xh7wivPx5SeC4
ttiKB//eyVr905IuWh3Ek9hQZx9FnVGulnALdo2nERSRm0O0KEeqA78oJdIZ
lkc8X8yaqsY//wpNQNFkyN5Wlo8IsNiIpIr+UdZlJZEqoIOmqWH/WjJCZs+5
tB1AikL1vSiDYrvs5XYrGywu87mETCq9VMkoxsW2hJ8ffZ6AlKFvI4voRIye
Z8y933MMnMUxJ00qyJe65gaoD5/+zhyrbacfzII8rYHa9fPkK65DdmSlQgtf
PKeLOSlwFGjHo9w4wMApl8cTRqdSXL0A1MchULpH3eDhDhaffi2GmKZyYjlM
z6SHgjbMq4goh9ef7AwMBB44tmux1dBjpiAP8JvNoR3jBEoJGJrPX5Ia/pDw
XuIvWT1vopATbQDNow8MITfeozZEwRYX96I86xJsPcvmDFSGbGxxu9DFQslb
RmRE2LIdd2ak7kAiJIi7jL21d4hWgT377xlXANrCDFkGGLdSRhH2aKVpbO2p
W4cL/M3/5r6sCwObyfvsajgynWuBBHKQXu4eVNfkjgOVzctbm9Jq7+3h+sHf
Sj3CTwxr1BWY1vDbYtybQR6l1sQyQfug1ghOZiAw0MaK71fbYsRtGSoW7cPn
F9GnwkMp1RAlyMy0EWDR83xXe36njc+DV6524e0KHE4ZKEXaBJn8vltk8fnd
Jh5fiqTPS8K5MySGrYq4JXea2kpt58a5/GNNRWttlzCuXv3MCGeGRkUEUDcz
HS1jhjPjxDEBK3bgPCGhTx81qmYvN5Hz3OQwr+g6a/blhmBvvaeWnkK1x2r9
Z+Icx0UZwQoI4SdyZ+loIyQtUJgyWX5vyvAQLqRnMfGrh6KSYUCaHNMR2pu7
WsB5gl9XqJmtD8V3Ks52Vqnunlw/DffDXYDIEDKtD/8yLwdyx1I5CUOeazW+
cu5h6jMtQiEDF6YUixX0Nvwv3V50BPluUHsrq+6iEQfRlWs3iI5gVWAvAhdl
YM5U2FR00tzDvjZcMSaAz2scychzSghDSet+qLPYEtPlcM2gFUGoRR1h69Li
5tD+CjD7GYq/Zk17Ud9mXSq8PyhsmplFyEmq/6gYNOG4m78nhoIlY45xp8W9
BW28fR5qapVXs6hvZMvwDgiFcUW8Iykw8M4W7/fNoOOxgGEkzG+wHWTIbXRx
lKXFohg9TxKeoMUr88UH+ipkjEBGzZVoiGqoBFYyjtKm1OJEyQWoK9dZzK3H
oKN8Y3Kd4q/DuN7bezX2cuNPXAROGSVBgw/nb79Vv8CwZ++59xT6h1ntGx77
QrmwAXy0i0XOzXIDiXxPyVFIb0+e0gbd52WzBWbOkP6I5nX1S1bdU3FlcXxj
e9CYPhR4OSvZMhZ3A+ztqT3J6bVE0oOzg3NMWrVojp9zmgVanUrhXf6vWacC
XyG6Gw89d9THjGI8cYuKz74hti0aluAjpRjxyZ/5NedDL0ZIoEaMOr/YSwAr
zbkEJRc42WW9J4z+sbaugRSARec+9svAb+4SVa/L/FumQOx/R0zlskiznzP0
5Doge7ThTOPjsnCpMwhO2pWJ4fZXm9xsCzYsP/pNHEv1jkhQ6D5BYI6PZQX9
yHjj8xGIrmrF/jADQyt3Lf+iAj7cMFlrnIS40OBEfn9JRLWm3WgYNwOe0x3Z
Wb9lyoxF5OKGA+rAQmokpK97tCreFmAmj6XVAAkpDKBM1cpHboKag0zYfLDR
gFwd32IWoT2pKsZJ480dzZpKDWc2nwRUP7PL5p/L8ScbCS/Hz50ssN7bistq
Y/w/Weu2qmjNg+wMguf2uZzHLwN3Rx1Jboz1HYR+a7XmZ3fWqsdeBMDDeS9q
OtHO5AfdG9yhlHV+zwhRBNodliAiIdTp4Pig2vDL3lsomQUNnxYYrpXwVaQ1
C5rx1/1uFMAekHPQe7sKhNkodIZi5OjhXAqPHK/SY//Da/1FagmcHxvZkbh2
6Wb3Ci3UFVhHrWSKl5Sb4xVgIK6Hqsyb/Ij1OLU3cDl+n5iR7G4GCJsOkhuc
pMiMQJoVjG1uCElIY7bQfoUAYTsO+YpZujW3dGRnp2c7rlcWzvu4zZKnm66Q
2STpdRavS8RmRvBfMvKGkbZPyZGB0wRj4tXb2+3lWyGivR6ehNZuOl1FsD/i
yKG4e5C5U5kU72T3sBG7iabhDVEbCiYsAI2nr1ajqPcL+dA7EpW1gfXMdEKD
HzdGM5vsTzWmRu4ocxB00w91v+zmCHlf0FnWI0+KPiCgsCto46g5tTdc5KpN
/25aXRbaYNfTCRbLztM2hMW0KShuTB23koL7UdyxpMy4WOYiXxxZS+CtJbjy
VycjZSJXDzIewqZ5r7fuAljrEcQLuyArfraM00HCUgaoV6LnIVaMKQCBBJbW
eIDfoYHh8CS/N+OtkrVUzbeFLUozPcVCGqxPk+uzrFbxCsBIB9yHQNKcoIN7
RfPxtulkxmkiOF2x60MWNl0biQWt4HdqypxF0R0GYX33pMIrPSypZ59Cr08v
knpRgElq85T0OBWgTtL6ukJ9WdsKLdss+qtT0cJ41G3cfojl+KSYBjpLz4nh
OcS7bYZ2CDJQwJt1Z0YCQo8pNiwmczjhC56KHrGSgsAL2Q4EwoSBKPyC78bc
UPqaYJTC5GSZ/kzJm9vdDriBBu6qCRnI7vhUcdRMEVcbAgmW6zzx6Kox6pxu
G0vdaupDCNO+eLfuHRtpCceMQMj7kQ+7v15i934+BxdcpAtbs1jc/gzIVocP
fpZYFf/uckfBN6biv8j01KfEouq02DE2Lx+yuaBdAzX1KLgQnAy13POnawzw
1G8Cv169LGpJ2K76ycHmOGE8FjfkaOrw/3r3tOr3TGeDLadqi5gSfvzYqsGq
Q7ECZFzysI3RSaaTVJzO5UPRbKE95t/v3llgASSQFBFL0ulFUGoKdqHxwqlO
yNhpb6CBNjv7my2+SH7h9AOhrm8iZSDDgy5aAQYpcA6m/6D0iZTAozXs4VK+
8IyptlOy2NbMWWMPBo95v9sY9VrIr0ZRfPy+siiSZbUWjgvZiQXDHKfkFdTL
zu6BLj5XPhfulTX0h2nrQOzxat4mDQ/VxSOw1ifwwUO7DJG3WnOgdgF2dwpU
cb2g8S47n0iLk3/hOOwwkUMONuySe3mnus7ZXBBkTXZ4FtTaLVZLUkrVsJUA
QZ+yp2aeaGIfkLJDtgNFoVGd/dNzOsp+AZJYcR22RiDb7RCQQMjsBYxODOoP
8zpgNLec6T5JoAW9bLyRmALmfKBK9H9x2PhY3e8U88K/2kQkxQroJM+c3aWm
fzflvyeqmwTazPWzoPH9bFtaDjul8VkCsFpHc1AmOHN5hZ6saXnXrpNuZBqN
KAoUSCxtHN2GrN05DIDkPBve4ptJS3C6bjntFSaDYynPaP7XslhSoNbCFrFa
UUsQHObnqMCeyo1yvgTMgUqxEv3MxDzPQJiQusY3pKODw8aMzwKGD9s73LQL
pSIM3u0u9wDiILZOtfWEGDWQn94pb08r1dszcMwIFKV1uG3b0ry4SPs+5Nhu
JpstYM2t+ORaitOP6DCJYka6lJii8/wwsK9WVjOfFguNJHdkW5+rcdRBuuS5
uijqdTdGy7S/PJTfb9O44MNreLZ6eVWC5EfzGKVtIPUgKv4ToCdAAZqNe4RU
gaPOT65S/Pcl+ibFa1sgPdYXxv/dbTAmEn9tdfRWxhrrbii93KcZprQ+XCE4
d2wcnaNN4m8jH13lKp9Nhbih8lUySYvyM+Fpy/qQm1+P138lbjVuCofs1rSg
NAcEvBKpSGRV2In8uRPw9ySxqAp9oD7mc9E5LYIB238f/izL8IbFW90/yxR6
zI5NpgMNltqOiRLJa1P+Gql+LMpjAu1Acpnfow9G/iFPFil+m7MecXIrmX1c
lcPpVRROdlOGj/Hf3CgW7JwKJht+SrEjZzdcMe3N2mtU71zYZlCnwkSUSiVE
14vYE1eKcLozZ/DgQwFXqxiQVYz0H3lYDaZvDxqgWFvUxyPWJgpIvml3knD8
IsPKNaP3JUTxLsw5xrKSsAc9ntlYO4Ags6WmUSXC3YKuV7CQx/bVpiZ83oZw
4DxvOIU8piZqpQjnRtgByKk4EcUL/ua3K/2qT83QAMQQBdjPFh01oy7pA3ZZ
mHhd6RZ1ayb708A1LLALyjLN0RhLLNHRFedNiQ0qW2W7jQesc5Sz6ZlBVrjd
9ZEhNN6Bbm4aaw/FTmo1OgvTogcEkY5tI43kRs2jnydd7Kkp3y/3EbWqMEqb
mxpBwyEOyKTRH4Av+T8RePdYPrP7HPhJe5VtZ6soRWf3fCHODJR3O3w6d6ww
zGSWItRvIREx1b2L0g33+AUDtVhPxtvKZbVLcO0EweaFDEisG3tNAKPOw9Sl
k/9uteVCdTzh6w4eE5MSHvBYkKL7yGY2EvzTIKbsYUhH2kcY9CJDQWnFAMTI
S+TZmDpSw3xR8e7Gsk6znU1izKDzZsTPkP/Sf96AI90e+Fp5rwEjn4itezH7
/5Oje5Db4y5UHmtS1xqW+vTZjZ6llMzoL13ln31xyUfm8DnD/dsZlr7VX9NH
Bl3HdaTiq+XK3MHg+00hCDEXRk3QG34LTGwT1YYKpy1vQXZlCEqbFMik3l88
K/vUFC5MRle48HFNHQNY+8lpOG0wQnjiFGGKZ/RwykwCUjAtYat8HDJ6SSFJ
uv2J8uCeHsrXSpkBafR80Nn35dCy5TENO1we1WDGCLJLmhzGEzxAY/I5F1KQ
6v6y7XHSFH9ef3CwyzeE4ageeclpxM5xwhPVLHi5FS2OxsUHT24nqHMC6tQL
j1STRrqbayNkljOSUGs7hcy/7bl/tcCyZ7tSBnBhkmGx41XEqgBY9BFbBfnR
7JkU2eh1X8LniWoK14Fw8d8wLr/yiW6vdYHQ2FWJuHeDjQIIUDpvzJnMPIvg
HoZvCA/vk02HHmjrfsoYW0GF2c9mDxtzfBRrKEQbzDxsjEW6x9ANIoAS7vGo
zx0LCqkOP/qWm6eSYlYJKR05YRTPlGNB9d5NaZbnBc1/D90s8t7oWFVmRzAj
T8vYcIreIBMoJ/LLC7Ehck2IQkZP4duoxYI370NhmHug+hb2tNuP3KpRfedT
roIw10+5gEJuwDebDTYxXp668XQsBA23XrPEfvU4OfM/8b5U1SOxQo58p1iw
PDkBX1TTcNpKnj+xFmlIzeAZRk4EcQGl+Vbmj9aj9GgTyGJsTNgVl/GItpaU
/v2zp2d4XMkDtpRxCDTQOwp8u7JH+DswK4vbGINmaXhGJuLFTSyfWAweLKPK
piCQdMA7TLNtHj7yjyOGmU3c6OgBJahlsnazSiq5SCETM71vd60//l63nS9S
ULCpYTDF+SET7FRyERn/3MIiUEpei3CO59hR6sJq9AAcx/vNhd9YXgb8tiQG
B1NlwPJOnM9w+GjMUolvXQ40FLc7flxhuesqLLD1YW0ha0dw0X/es3958vvj
6zKxTGLraPaY5r//ispeDxGKRNido70SwNwZRq3tROVDtkCbr9VLfXgL2bqW
2qWmWi0oKHTyoYIIbns03D/PcEMjeQFBiIfTI5dXIDPW91GZod/6u8YqnIqw
bbmvk7x+0XTOGkkarGPALEIrhVmJT8hVswvdx2unXH8qwZCQ5aNaeYUtTFde
txh8mHs7ssw3E/y2QRdMHqo00e2bis46sSud12vIFkC6N6e1Z2MpXSRWS0HE
0wBp1IDJ0T+O+RseDaDgVoWfRVd8PPd74Y3Z/7//7kIQIbOrEKYxTE9+8VNs
Imglmih8fRZkbaXmxXkmSE6APu1k8STwM0N0rNWuMMBccpEGxrpZM3u4Wk47
//zPvA7v8SomWfw+YQWlUoFAjCoowybLi55yxklOvmsjshPpUKKvK9blgMXE
zuVnvbQe51YENCznV7HbkxQ+yqDSP4kWdx27cHqO6+k3+AtiYvhjyVGK3ttd
xDr2yiwrSj/qgcg7vkWKNkSMJwA56ZIZ8E7hm0lW6KVPYhwSLbsPzozKYek6
FAcenHYQDxNbKK33UBgnmM0/FVv76obb+s3sCNNukOUw1W1HuN2kNOW/jccq
XxRLVKOXYzRonv2UO4NOimWB7YaT8tvXvqB2TgDF1qqnu5gmtB51WxqcD4Mu
vBiE2TH9YZ8SpmzMMVkizaAsGMh3LhlUdVO4jN3MKhkc8dTmg5SL5icG5tsG
IOwhjhtwIxKHae4hnf1Rz4l7+7OO1IIgu/d/C1OMi/Qj2YpthtOhWEsgkqJ2
pPDl60wIzop2kxbP98BMEqG4EM1IoYKxJE5d/bygJPSAI3PTFMdVWd9Nufc6
0MjMrYklei6Ztii/RnZ/urNlXl7yfGIJbKGeFvrFIDF/Rz1pNJgeawnNnRte
b1V16iDTCFd/1NsHpteA5C8Bt1SKB9/fT6oXmD3EmDoEpqgZAi1OGsq9StfQ
5xmzzSBjANNXkQKbJKNwJ6BHeknWjkfbCWI+zd50ssQloT+/1vJPbIS10bLV
80+9y3mGRxJtS0p1E408gzD4QiP/+Z5/nEVpWAI6UujgVpQjB6Xop6AqZtsZ
vdNvni4KgElwypE5NbAgepqwJZwZ3IJOXSfHNhVfyO2U/pdemrCqZUz+cG7e
802qyp7BAWQK3QbF8leotuAzYKMZS0LfclUwNP84Kagn/MenX358FUMlOkbk
M/MnZmMNVpMjqzEv3ofNmVgYibKI6n76Cd2JvOgS7v5K7O+NWbDpjUD35jwx
16eoobNOrF29TmrqOUPS2rqlsRoAZLdMvDUVyXbROeUFFrLEtUBenaiZgrL2
2rwZzlRdQ/7eS7lm3YNRoBII1HZMY8GJFL6D4sr4BpJiN4MTAvs+QVd1cu7I
mbliEIof6QOOO9B0SiypEFCPl//aCfVQe7hAgwk+xxn/V1zV3fqnSEL5Dvyl
d95ZcEG1HNOARN860ANw3DrTTRAP5yVESdVwOmm56tqJBjsrNXkyDrD55YTH
GstFqp+ZMhGOC0uqDnqMJydZYhtMusAajQb1jqmYxXXIPSHNunXkITSfVBJn
4EWKdC2Xv2GclREXuTYruzxSv9utjpMC5iXh83qPZ1il8LEAINby8usjb5td
59hqfWrMpeJXHAzOrI5bpvF0QuqzsVN/J/7gHitFuBXyFEPVHwWxr2wlbsqz
gulgEnf4F1W1XQtO6GwiBo72uuDa3aH1D5Fq0MgMtkDQYlkLfxW5bfATEnwY
mPfrZDi3Xyt9NY4xLOs7xZoQPksAhS7AZiG9cRvUeG4R14VtIHnDI23L/gUV
Dpp/RRVju4lApi/F8HJ1HO7H441lcFvIqPNYuvs9Z1qYifXXrj2Q3gsobhwO
ZPmJJROlxQXp+h4TZixobwOXya1mC1J+XVgsvSDRM6RWw7qloG5Zvotntp08
kf0en4Ls5HGaw8t8toWzfdRpVqAQZDgCU2pVSJUjV0ZyUdlTclvmHEHcNCWW
r3JrllV0TWO48fCjO6XqMajZt8o/kq67knwon4DUlrY3Cu+xc2F5UgfTXphN
Gg/LoZZytw1fMblVvaqoXvDcF++rEgP55mh0gvw+NP5Naj/5qqPfYcx0Niqi
U72jRnWAVvGAB/RKlhADfesN+z9UsZz91blLG3uQyJ6bB5uLabqY8jUbkFVu
JjDjj7hF8gh8KzkByYan/k52juo4TG+IFwHejqq8cVsQSOYjIT6rM+/B/4ps
L2sISoDc049ZiknvLq6CGRMXi2CgowpT8zNeftp3DOzOobutET2ChCGpg8PW
n6/pk3yJmwPNNzfddNVr+nskLfDbtUzbnaG5OXPJeBtYjsFdOwIiMoiNHT60
b4jbrsHsaSC1zgf2roVAPZhL2aF47uhwVsWbOpcS0Ld2fjDxfrINd0kqVuM9
Sx+BgQnzu6Nk+2bThdcz8Im029kYRX28Y68cYn7knUOp+icRsANLVeektJFL
zHS9m0HdjYABWQFAZ/H4KnaFRAsCo1TXZmACO4F1v7DOcxmbSuMwOaZt1asR
B1GWryvu1qpCVQzlP7+1zPAymi9mnhIGTY66e8Og9swDwd5h3h3OGrVaB1bv
zx1Way1Tfe/sPQkAcMoPY+Nu3/5JDgvlpwNZQM+AH6yOPceUJl58h3tGttrW
ySNGqQiAfhqaMBR4mvBduYFOOpHKf3iRyz+5nqAelrFFpjsA6tY+yrNOzSXh
ZaxL0SZ2l53CgD+L2cHcgFIjxw8TqpUTeWZdd4lRcQaget1Zl489gL3sesIm
RItq41igs0LKqAwGa2YNv2Qi/8L39uySm89iu+44cApRb9ndMaNm4So0wC3m
e0y7831rWeRw3QVlrIba45UjnuH3Uhd8jXwyv8klR4n3LSXwJlVU2bT7sg/W
lF9Hz43eLAxhh4Bb0Pz+ksCmJzbT6QU0JT9NrwEIBbl2HsXr2KLQF7Kcck5d
YeD17CuNUoLLUfXrnoAzI4tezvL7lrXMv/GQVd8wwvjk0tkwJOS818H53VCd
XISwftJyGTADoqxsND4G/SOb0G95uAfu8gmIrDdyz6t74hZr/VmcsDQMTFbn
iQCOco0tV3ULhdiOXObEzosViihDY07EEQVjcHaF0zhs9+nNXqwzAYMx5cNm
CT7wB09rFbbhAupRJ8e8ByI8T4Syg4rMlkoWDEf3Zh+Pz2ZlhoBr2ojdBhvL
Yb9n96Kt6jKgC62DHLxFae0JGOuNtNSCQ7XM8vVRcBkI7BO5hCucnHricWw5
j6TPZChiXFnR+9bFmej9TOiPd2QAW/MVzwt78eozjVgh4nALYRtPbetwIrJq
J5ogh6V3tZntmCUOa+dlV9UmXpUotRElOmDRNuemrCdG7U1nsgGlN9a78FCt
i4VGUXN68aE+iLvfkJfIPDXLo3UUjnkDtDh1QGcfnCY+goaJsg9qu0ZdV/ys
akg1OABfnlDeQkLcZlxbSg2P2mWH3Yc+InKGftxgXayvm/5yMTh5elLQKfhZ
Nluohcj0BR4tyQJ1DUSFZ5jlZINH4zjhEMvSuULFWCVKei6OpRozgEFM+23E
0t478NTOYJTe1qTy8/vRyy56GxuHBREHVp8w5BC4rXhyJQOnZrLOmNN8x2Hq
CVIVMSHRTirnZshQrTceKFIQblCBQpjQsehxZVq8L74MOA8zpzRsrJhrKL1N
BXmND0EnubBNupTjc4s6I13rtkmQ5YEXN6mgGZpIgIcvnS4RDtOdbC1BGSpf
s2kHANP7mTFUVLy2XyWENOSInbrI6sbRR+bGonuDN48BuMGWsBU7vmlLSMqx
UlKROm0TJXMrkP4b3et+aY+Nd0H/nDXHFSPFO/QQIIDv3N0nn15f4txgzkxK
3FtEdxvsmBlx+6MwNA/BJNjL9GJxlbRuEg+tXf5IcfGXF4bBcDTfLqZ1j5ot
6hh4h/+d01K/J4GCwxF/9Kv4S03RLTfF2iy7qUAA2PaRh2RwaGb8A2tSgt64
tej+dmX3h1ZMWPtpV4QnFt/ZW41Gqs30TSgn/Q/COzfQpGKPE/cRRooHkZjz
AdJ+S4GBMi1A7CYMqErcA/c6eH0OR3J3zeNc9slU8KuRB0djn6QtyT0nxZ70
d8vtLDyoMKWB5WFM14cLxlBao+b+xotyDSMXAhL/w+gfTUBKdX4nplcdjuWH
yU6y1XSiCjIz/EbE/9xui7YZ2yIZ2g+42q5YIXCEZzUpDzTj3e1sjUa+aham
yftnZn13jSBzSucexowyTan8AE7mAmum4ZPQsgdAjVYYa6kylaXy+sn8TRod
XNMvq7FVtE3YTqb978zafFsTPZ+ptiU3Gq0GJoPZIZ/XDyqTgHXudQhMsGy0
3HuBgBzLE8f//gUfrMfr8SsbqPRMmwz0ivCYS8PqnOuxcjKi+c+3t2PXp9TQ
CRkNVSqQitnL0bNoBostWfCeuydr0orMAjuCas9aXPd75QZhKpesIa5ev41c
/7JoCDFDcFyvrn2lQ7w0VSgjtDvaAku4eeJhfC+tLGpxo+fd6aClzCGC77Pd
QdTD7AwKXhIGMPMsOcVrWA/U9JWLm8ykNehen03kVrGcQPmy60tl5b7O0M8d
WuaaXN/JHEUQ0D5hcIIS7IHJ2Z4RDDvvbk+uBm3z9KKmdwASEdgrfsh3w+OY
kAE6pYjK2l7PE3iZGZ2bkwGeeb70tGLuhSwkm5nLJ97AMJj6cbtYx72iqYmq
cwfpPze8X1uJ8W/tR0sS9xtFA3tejc1diUQqivQdCliKH3JjJGDhqOEo+H+g
oJjz8s8kqIvhDDHW3h5T2YuH7PyRmZ8vc0yJ3ySn6EOApSBkPIG96dc5s1YD
xWrliRYZJWeRukO3rF9MywX4OnAovlHolytjLyBFh5hnw+zlYQv7pA/QVxJx
Fve9mHUAIuvvS6VkRlAvc0WVBkeaNbJHu2DrHYtfd/s9uYk8k3VT1tiLbnZf
pZYzvGmrKpAtbSE0EH3/2Uybdnkz0EE7lhZ0W4wOAqApq1orSr3veOfbRiAX
7vrGQAF4vvenpLtE+kFjh28JrDvrWv0cLPQLmF/BUhMH8WLFKNLn7ff2AWlq
JxfzpgodJiwpgHLtu/Vb5iAVl59FJmIJ7PWiIq71IGODKDC3jADPsa0eD4EB
FZVRMKSVXJHKbd/xFRH+ngwiad/uiArjHrQ1bpODHhsjlvFgPyLAyYsOFLZB
H1smFcJq1XHWAtrRM0snxXJAWp+yYA6i2yieXgGZgNazcb8NQD7g+C+JzYJs
wDeej0n+HcrZJPXOt/TZjt+R7+yZPbfJCrXWl4VOIO4QE7PMXWuXlXvCLv/6
39mtAB2ifxmiTbFXA28QPQW97d05y24lXtUb17E78fMrveiKZotclYdz0EvS
7gsaNAbVnQGNTYMpYwoTwIdBa/RyFm/8Q517DQkP8jaA7wlmkZeRbYXhEugX
fH2s4oI/OglkGOvfn7Ti5HuxlzzSJwpc+PiaSVvvJkwnNfpY3w7WZn6wJ6xb
SBSQw95Mo6+rL6SHZH4qaaeFVgb5Et2a//l5vQYXkLJb+YJGYJNx5G2tE8pZ
U/f+a4PkYVStrPotVHtJZmY4PVxa6oAztdJ8PIWNaxFaJEqt7FCRkYE/Bnfy
YslgykJM+GvKXt2pVbc6IycqJ8YejP8vNCM4FX1HGJ0c2G2wLxKYN0lliw8i
0BFMm7DXzNm9XmHXwYOrhAzCzN6kmlRPi4qL2OtiTUW5ilaCN4REzNHRgNDk
jVCsqcaR9EuNXbNTsE+sf0j8WmwsmQ9WV1fnZYEi4a+JGWJl+rNfECpWoWGK
yNgoT5d+GeGVP5KmNpPafhm15ASbGX6rXABlFwNWnrDrsu2c03KfNd7Hf7DD
wHD/mFMsBLWqzA4U8QYi/T79/jutFK0q3xtcaksPSMaJ35KtXIvfEgdeDgyL
h08bvzm/0p2WvVM4cVP5YWNywGQBZCr9Ks5jRnwrIrE3Uhr5Z1PaaMsynEQI
CvSbv5Chgcv+3gBv++r4gfFh1mla4FJsqyRco4XW5fTCqkSwzQKQ+h9VNEhA
P/5u34pwS1QDvkCVMl0W88T+N38T+K/b/VelTfH4xEeRlEuQHT0zxD7x1YAj
L2L4ry4p4eFIxe/CXf4769T+INDQzMmnFJdJ4m9KJU8nkID3ZAgXacDyyrF7
l/a7V27yXPNk2ua9WRTSJVUs/4A9sznPUbmn/gXVupxEsUwHsjV4QOtl8U3B
w7iCLA91BcWLwNwK3brWSuMHnKb+b2CENwrxLQyC8vNvnAgzVs8Z2XaF58Cz
g7o4PcFHH9DzdPK4i8/rqfkdhNeD4HLp95o22ItEmGA1lqfTsdi8XQ1XY6+5
pUSJyy923gCd6ViYPOlqjOgrLbf2j5EdSZinaRBdNbSr7/BmTUpMpHh9J6dT
03PfkJ9ka/02+QeZqOjStBzU8zVKRtbyzmRQBnam7UgTdSsnkkMxK98tN/1T
fTg73lM2a5xIirdzmnMzDcIchFSYjdoQZv0Oz/pgNZotfZNYEJ8Oo/pGsZVE
J9Z5e0bs+QrCLnSHzM9P91w6Y0mjZbVJpGnshG5vKQziWKa0+Y/mlkYFnPl+
8hm5v9le5X1L7gLEOVWqzR41I56FFqH1n0t+eMQSY1UZj4meCU/9u+s6ZKSm
ajqbW9Cn075ypmj3OdKEAN/x+p78mWjgZXMmLr+GjjWh2VGbW7Oss3/Dc15Q
zlJ+Cl9MgMVgzxbXerTXdvy2KLPVllzgr3Sr1yODX4kJnsKf44kfuEnbRWPm
+VKeUGbI0WGePa8CbHKSRXOarvxORq3Pphhw3dgluWmjx7ObpXZ6W583B9Cn
NTVqMVi4iJyLWAHeYUhd3tQ4/55mzNUS+otA2m9WVXvzcgjCs2KdLNwOxbW7
W9GjqFN7HWmdC4BoMPqgIHZtLkLUuHrndgUvfDX00qqan4SjY3kS8Y6gwcJF
Pm46UanpgNw1IUggytWGMsCyTKQrawm+cTH6d4LXc9fZZ3BA/Q1/1o4Az7Sy
ayAN6vuTXeTUPnLtcBWRdKbjRA35quqd0NCCfLgQvrBANNzWXC0dswZOsNI7
2lnyD4AxoNw2k01Yh2xWANcE2t56z+XtPhNHv3ADSjc17EmYMNJa5VLUOscl
B0GJhk2ar7OO69qLR/MMaymNjqyl1kHIrs6BTEFkIXhupXDehetTDvWAyHy+
PouaKV+xNe56zD37VsrpNJXBku+K/KoVM5ueSJLxQmA1tBYYK3g+Bd6gK7rk
7fXyYe1Bfj3tZjx+xJYzKI7Eq7cuThKfCAyUg4LIixiUZAmxIgcZfdotzgtz
HPoxqgGxUjcojJ2h+nvo1xCDeRh9iE4RLgO7+77suUA1ISOvXfyjxIg78f+9
aWRi/JIxVe0i2mHs1tnYI74XVjLLthYaIOAVHG6GaaLu2J7PucVQc2F08zRH
6hskM4cgwihxTYg6mDYp3QgJ9cJu8VGhL5eCiJyK/Lkd3rHg+7EE1go13WTI
x5vn9tXtEBp1kQNktHjm9H6TmeYBSs9my3mNDHqBzBeDUTLtaM1pQtWwTDqf
KZlSdzgThFX7cklatHGaXBgNWEBWynLduuf2s8cUxZ2URmqPP0La4QErxuiO
jrNa1XSsIdfxa7wTBuTGaRP+Dk2CD+CTwtcx6NZEIQA+h677YTalFCGS+TEt
l8YCGHnAzV7TYXsVQYgTIGxafh5b2WOwF0J2gZOsL3NtWpzxNIONxsQyLSHf
MbyBSHGAqvyHjv3XUD83objxdj8XJ7TDfYeAYxHaKDF6ttAWYUbs+PbId04r
KR+PU1eS2X/aXaBgzZoLoNVXwGw9Ife4+FTx9HxLu06ENPzE1i6k1L6MfMBc
2uN2+JxScFDlgFOjqO8M3EeF5VyYPTpmSZ6MLpSbxTQQdSt0VCUJtEb1PrqO
msotqMEDbgRRsSCnO6B/tnyMaxQavsd9LS/KofKk/gWUhqpxUgA29nPzb4Wj
28rLjKKQnopSlJpnykHUU/ySuxwIgJN5s3+5NGL59knpMFb7x1GY00+zJUik
5y1EaNRj3ZH9uCxEKO1bWEVBRAV6vU1xEa7WKYr4iM+CHz6cuIaj7tZuvRO/
NtTnCZlbVh5JURk8776ac2ARAgFGxesvVvcAVlrtakkaI9Kl6qXr6GJkLDRJ
FWjWbZ/mTWOJKlNruFOYPyuQ6rxbwdcbVbIQm0pcvVT+oBsZshaetA1cjO3p
XC+UagERB0bpZK5z393Waoga6rmgTas+hK0upaSipGPbLprDhcM004izTFO4
JgxKCnrgHrtCW26Olyqmq4xFUqVdqC3wyQtTaxJMEsstMknxTwxM7B2axsWB
SqhgUBi7fbnlHsVtZkZmoUpwtciWctHqjGHb1rGFv2BXfxZtYD4ewaK+hlQM
9x+qwvx1Yab0yr21hwTPrODWiBVXdN91hyHsYTgPIVo+erXxY0Hj+nmnwB7s
fX+nBc03KZLO+1z7D+Gq7FBcS48K8m19aW3y+PBzwRpQtCh0S5dy+Bwhigl2
XBAxaRspSq7dDfjEdmyIQnXQUmwDgK5WnGGbo8LZxupHJ5mIx3LPy4BESeR5
e/GrQmfTGkwrjitwCz+pw+Tcmn+F4iuPMnLtLN28gCP8wt1p0oGUryW8Ujf4
Swh8iX4bew0aaKKg7+Bxn3j1MIU544SxZeTYpX4Xi+ZCGA6iNKVyInjCXVI1
X3qXXWXfufAJpJWP8hK6TeXxSQVGOmJ2xMn3179MavU0iFj4JQs/hePSu0mD
5C3XiZn9I0GTUkeI9GC655QQT91ZJ5FZEd3Q1ceZYzq50MEtVbKYk7aGJ5x4
9PCPK7xOYfqG6A7oAp7gSpjDfA97KhijeyRTm+6Cd0R4f8iAbI/7QtgS1M/y
yX/FQzSc9thBKMQNDXiMjUigqcvjQ3tMIovug9KmStjbIp++So4SIOkpBCDr
4SUTfq0mL0QgxuzwGgTP7tEbHleM4X2XxUY0yvOdhGd3dBme7omO9xCJbuqf
JKSnKQ9xBv5jXOcHwe28KWR2s0nTbMmLvIjHYhhpSYiR3q41X2fZMC9v9YTZ
3WAZWXwlSOIy8dxJzrKrnkfLZ12ySaV32m3lipohy+jEgh+RGndY1nIPggAk
GGa0ipCjps0C3Cj5ZDSxvy/iAIKIqQKSMuwl69U2sNuGlmiN2hu+aKCwXxh2
piUpyi56tx8dyYUNARDm27cmagepXe2pqCF814U/B88p9L8zk9szXzT0EWgE
LUVLLMe1xzLs61SyATyJf3taCJ712hSdP00Uo9TyYZmcpeXm9pZ9kslVcf4V
9MpUwMCkaoSuwOg+XcAmfdI7JTvOozoaqPDfzQxdEqUIxz3VxLK5RlRkjDCW
fxubfi0NffEfQO25lnuGTUy7DkS6CRYZDK2sYUfMG8c8xyIxXE3ivc4phDok
uqeogOQUVYrh7P3YECM7XIWMtIfKmugMRB6wVq0JmE8z2/mub4/plewtZ5l+
+g3OmMVAU+fiR2Qs/so3HdlqRBGIfjIw3ll3KnoydX9/AzfHZK0gFu5fmxda
GS48Djz8PC50iL1yIqodkjJFRakS0RPrxz/Z7Cno767HS5KuvAoocshgZxIU
iAMl/ZqNnOtDp+0QnEco0akSgdIc5fAmzkpIE7msUZs3PW0ZbWf+59h2IUPf
my5zCiX3yvAZ6+si5WuzgNfcyfr6fRYiOdqz/LAjsWZqgt7jqUyY3BjlkhJ+
FJY/7E5QdizMmJ91vsXRqeDdzuUXWR17gk4UysDKsM8D3IylruOPaD9wQ9vr
us2CLRaVV2Alvl8HB/2m5jNBlPSRfvumLWb1al507JaGUjdu4W7DWgWn14u8
DWCz9GlhlRxyU2aSQm7ekSybggmYakT/OkRY8upamjzqqS1Dcz0vV5bHR5AW
jKdvhLy12B7kc5honESJykG/6ktG81E2T+NsKrGQ1PhfUf8gwNzmUbpYUM+J
eKax9UZKMt5PFKsQPB59QCssYTqd9KJvMbqqO+hw7G+ntzV1pk+izx0fxFl+
1BTVniP5t80eDwtWhJvfltW0IIcxP0PQpgF5wq5Hyz2kMoOgvYRVEoI25CAe
HHBRC+RAghROIh/WJZVrFaKmiZFN2OOSnfNBQPdu1pTisUjqTCEVql1JlMTJ
gZKr5a6zc1GWUNbGubwW3ArmvW4UaE1jr/Rerf2D9cyDpXdPteFs0ByIupDc
1xlYgekLpMEvALYICBxsXxwyvFJs2HAhvnNrRNqcgAKd+1VFJI0IK7pz8IbM
RhRzXecoKFKhylMp9MZj0ihOeK3g6GU942NiPGyThy9inRUvzes3ZdSsjmNu
3hmklURP/wZcaok+ngdxoikVTS+Q5rTQej4s4BAqJ2TUbnM96BDa1DkFLigl
nr8tmd1+ziAWiT5ET1WwoHTjqscJjUbIJvHWfAg6fogslsaCoRjy5me13s7P
VJRczhfjT3xYVuQxYEEG5wuJv/+jm71FJv/kGYYJak8fzktmghoLpgCL9lbu
StOLokvEg3W97SfKJK3pDI50+/3ubB55L6SYZtRXAAjGQBlN3FDwQOM6wvPM
n3coGgQdYwvoVxmzVU61mlTuGW/Nh/qZlampSrTtNH1quxt8pttmj7CMeJeG
KsCh+/fCo4MM0rVgdbKa8HAVVV4K2nsx8txA89UBnUFDFBAd+fNKmrHGZ+CF
ITfl5+UdvU13XQXE6anhaKWE+SH0nmVX/t3styh8A0xlR/xmEhMLfJ8NbXOj
D2+/RO04LtpVONSCJxewyyHtGUl30ObYNZ/d2wKGP67zM2+MAVx0jMjHDUAW
UhKAlGan3UvZV7/OhzI+rALYrn/RJ5YKnNyomSepb2lYXEqdHp2rYCaslGv4
J/MPewHzx/137nNS7pWX+US+NHMY1Mz9KjiEVOqHD7tyTBgELUCF5466o9VP
R1Nsw00VXqPelRfrTOPvLQLvlZmvhh3QkHMo6DnGRu3QKY6Z8sADSpj207AV
GstGbwHySSQiRGoBiM3yHzQWNgzC1kp5xslQzwyPQ/Mk8aP3Y0UYIJxnx7oh
AkfUise1QfyCYZkFpJahKYGO+weY0cgryDZaKLtPHEwe2Sf1oFcMF1VzXC8o
G99mBnOrKGd7Si5Tc0kilZSzSPZU5KXfQbaW2AaQFsYcIoy2PuFSCoHP3tny
ZR/QlqAqHPDcelVnuG3ISSPuX8N68XlG8n2fWSfzmzYR30zXfvHj9ggTMA/+
2SQdn2l/5GbDZdqDep8i72OtsmfIycAuPlAcJTACReTmafyuabkr8Js3lneN
Of/TYG/5BBPxS5Mh/z9+MJ+lEKKw5JflKz0aezVjcIIYyQZsdsXw3dm+RDyn
zfVzl7dkFoU1Eu3vVp2n2Di+0DytOW/zs1grfo1/JjC+DvKv/vHH0heEN0Cq
CMKusRAa08wphAzIVFwTH4Z/0yohXgdnBhGIj2Ww3ccoodt7dofVFCJwRgUT
UD/W5S8gjEUaYt9ypEqz7WIFxz9SmjgeF1D4a8WMkc2ppY0/Y34PaW7/dqqY
iJn9s8BfOHofixav/1/t/4gmgLsxpSylhjYWDgcCmbKnKsPU+FnW+d15fn5a
MN/WMA+xeEPIlsslLqIaE3fGiS305vYxJtuF0WSXxFHU5Nif8IS6nVVKzySG
IqjcF+IWvOb+Y9eLoBDvwWavOPc2fj0tyrCjhPXEpURGX18ViHpVvAZg5Ge6
xL3rLQ3PjPrXVxllRuHjQCOCFzHiCccKQ1qJF8q2FFsS5j4A0i6UNK+mVJYh
09zls2LdPY1t4k7FEyjhPmT1EluPBVuhVxaLOsd2BJzFGot1pUtkgJwEMVkp
vLBAGfsLEMvzJGfd8zrQki9Salj6qOL5oDbNyY+9VGjvGrMFz/VblTFGLTvz
v73ueWFfIG+WLgrQJQ5O39oRiZtz40kadYEaCQScEiDhhNpz0XQGZrlJq08P
+nJmCioKAXCBOEFsmbxT3JFnnhYsbWOSMzLcdEV31CdWiZ9cnFqRtdiqucbZ
XwEeQFrZwzjOjZHUVzJURxPm62j2yk+YpezFM/gxeDHuqp6kLVe0PbL3hWL7
01i297ZakqICgD7LF9XF2A7m4y4IB3IF83um6/uDGMouW+pRe5H7B4znApTT
TlDXdsetq0drqWoZy+b2SQeI3oWEOeBjd/3dpgCkNmyG/KlsvbQIzrgdtaBf
Id6WnSkEwD7SNxF9cAXuPyVWlyKP8rlh2gCe+gpZ0pJZ75adS1k9nZAi0C+i
K7Y83UAoU3d6n3XkkhQnYUcm7YmpEqg8dNvHNMVuY47cUEIBy7Bjj435HSmG
0lGHdm38JOSvhScWiU+RInBTCWkx1Bvnycsb8P04Y0DVXUs+Lequ+wmHNS8b
z4nMx0b5nw2RvS6eCS3wJKhb3g+Bfo6ltrZ4rQBqV3jnb7TznBvA5yYnmd3e
FSxulSmIffJ641g0dPafGS52VnxSDrZzexl2Gm864SlPGPzTVpAuY+duGk1B
CzgZrGjTdZ6+qd3fLC7F6HeXOxUspTJwa0/UjXdi7R0sB2WsT1TgQU9zHwu/
ym/5DCYFcVHBcWoUxVhAyd77k8Q5TuNvkcexBcE9U+fic27OfmufNSrPMZhb
FoPzr/IlVUpeis22MItHf0LbBMyvj1UiqLjZsZq+5xxdK+hNrv6LJiWmUxbQ
u81eKspLBUK0QHBGYVBx/IWDbdMLKZvYDt/trN7sY+mHCi1O5Ntc1Tejtjs9
S7CO6p/VcO0ZfXFT74zK9D+WPXs2Y8QypVGR88gr7F6oXssoAhIuTKqxymUd
GEGMxJvy/fT5htlGdxkcjunGmJcJWnS6tVbY3u/qFD0dZLVtRfrTv3VF7wPf
6VELSDzfv0HMJRQVCBLP4bFZiHaO/R2h+7psM2ILX+I2LCbC+6Lhjl2zgCtL
p9qSJoNw0LLFiehgRjohGtU0rVOKUSqlcOPRL76qX9D3opz1q4/Fhwt59Ewx
aY8Bxpo9U5bPZWgZg99guQoMrGBrOz/8eCgTPFRJJ7jg4WEApc9PqmoGmMB/
/btyEig2BLjE+fCeoGEO9JehHi2yg0+nu1Qlom61UTawAYPHeny6s5eoOi08
VKoe7smytHER1MnzXSdi6uOU1R853Tl4BupHJfUZfkuDMWtKl6N8kbm/Z00j
uRKHOZCt2Lwnnjg+ARsLDi8QubzeC8rfk7+Ut+9mF5PVrPDrBM/TFbR+02yG
qK6ht2vO23GrnM1CSj7klMI4+Iih7nYaGce6jGkNid8XT7FpanR1Cm6eQdVP
3a8Nowr6lIo/NC6HM7yva8H7d6SgdG18amiO4/jorV2g1JOeKwVh6GWftFAe
a1OCM2fI5JHy8vRX/l3bJRcdbYB7Sc4aUZlPpSPy+K3bD3tz/bGYbwYGXZgl
GaAzVfJLy/R3FNIuJPD57ecyGhwlgtjvatIdthLOaRJx0JTX7qk9Vzas5Voy
0oAOYwTrQOzl4j0p2fLMRMXWqHKpOuih3PmGxiJA3DEp0z29vRY+6X9psxv3
niuWDJAQcVbTKQYy2KS/DY9oJTQyBGWL9ZAIHVdsjpMOQa7BWlVLJQIJeOut
SKe8tmoVJ/bYMDY6PZV87EqxI9MTn2491sihZ/SmphQD2GFsTo6pKfNI31aI
CiklqH3zCKNLhPRR/kTayX5u620wgOesP1MF7jozXhgrZ2m0mKPFeC/B9wa7
aOSnGbMYuPXRfFviK5283epIHDKS5cGc95NX3tb3OPEFC94ASABhMruUA3U4
STuwr0zhFJauwP9KE6h2Pxs3e5cns32YlvwmbvBFoFWQYnjZOIXZOs/RymV0
95wU6ni23UDYhJs8fi+KevE1KctHpVFA7dQtDgM0IsMlA/9RfjvqO9FK5TvO
QObPipshIejQP/BFyrGgM8AK9NNu+gNUZrWgb1ugxz7CMt7ZuihcUie21yz9
+0GxERqZKi3pmR5UJ7lIUjVBmJ94m2L085aRu3GkvHiwyzOgx7J4D8mVfFyb
ltMZ0JkeY+0tivuEMITsu2TS0GJYfIZQyWKMp37R51X5t20IH2A3ZlHXnDWG
07622UYCUNhJR+puhGsynizUcLW8IjLs0/YyTl9cic5qX0OkhoF2ea+009rM
mo4J6zSfbACtT/08CpnjfwmdWjhbD4f9jlvXwDaj6vuX0DpdXyfyq7vdHpF0
0Yvt0Sx2q5E7LM+6WVdZb1hWwH5hErTNEFGAEDcp1reJY2ZryUAyucl7kKs0
A+6bAUenSRaIAqH5uaVhQ+U+zN1KObWWRLluB2KhvZVyOhORR94KZrnq1iEg
A0IoTYeq96ss8Mt+YHjsOo0SkHsCstO/bTihpbH48jF9ZltjWET21v9lTIaL
xcW9nV22cwY7XX/4cBdff7UTIr6Szai7E3cjgRv3uwsV+pCby4ttRn2tyS05
QrUf+aozoIw59if5pzZ9Tt3ZB627RAhTfbtFagW6HRA+aSIjg2Mi/poi1EjI
WNTpPOKvUdMHSkWdtxmRZKQJ3E9soPJ6lFnOYWhWluFQ0Gl6k4n6xpi8L7V3
jwzR9tZMRPuuWbmpKbQQKwvJth8MA6OXIPc27ZBX53gwOpxwZli4LwcrpY5p
fCI2p6Vi1jYiOM/IydK0VYxOW9Psa6R33UQNCqLl6hvsEavAhMXvj8VrTET3
31jpaKCgwDSZ1g1metNrzHle2SEXVSAqxO8Lv9lAMMxBJobAZ6N8adkJLBhi
MeOEKKnrvmCpmhtLFUPWQ42JZxcSptv7dmN8fLCvay0Xxajy5oD3VioMJ50p
dq+AYyaqePFNijJ1aih7mH5RJyPqDFz+L68tFnO9w4DRBW3G82HTu0icZ0oI
tOhwrevs5GTmvnkyHudDEc8dpbokQ4CBDmO+NMbHyp97bVBZpvNrzu/nyPRk
oWB19Yf54SK0afW431PFlFvP+c6i8RZqx4svY4K333sMnWanO5zlGedSGhSC
WjIULGbr95qZ21FzAsy+vYOD8fbCgOVvQkJK8u1LMYY4w9ZNhG8kLWLFWyVZ
ahSqZNkH7zkfaTMsnh5w9+WkgO/k/EtxntHTb7tW207OK6+rpU9xx1evTURy
Zf+MrfJlUrDVR3Na2hqIkez4yhw0H/qglffanC5L0dVPkqomMcSdSbsaezo0
SoJDk1Aj2XFBLtA03i22HLPs1RI5c+ntGFPqCTNeEv+9CHXpoa0gwcbGxlgl
Gs2AJEkw6KwOWyPX2TCV3OY0aL2w2ReDD+Io+Pew/P3RDcUWLNXX54x2wsvP
KZuR+UXOs9R8vVCGzNOwk4a0mtVXod8ueaiPlA2PJNkh8dbmL6PpGK5HeAet
m7UqwUi6c7fKO2IktPkGyOvUXZdk53uWW+vQCU+MYEeB6qnIr6iVUalo0+ju
rznKIMWVYyBAbda92jdzfoAmEuVK/84tnVJImhJv9tifsmYJ2d0Byvt9OisI
pKPokXtALfHZlCp8DXfhevY3YPcXtN6MZPKMb0emlO+YtL7ihCZa1Kpyg1op
URp0bMJoQc0mkKTziDGhLtL2dOTjJK5f13hIgwmZM4aWDjjVD0020D4/Th4H
SpQtAdxrEckYskwoIMMUtJpiNF6PW4Tg+V7Ih2Sqo3ksOgENEJuaQVi5jlgi
DC8YgPCVz9ZPlhLjidX/Yy9P9qPc4aXysnxNcrqgsVnqZYVIef+t1xrFosnl
N/hjA7dD0r10Z097HqWraRV3z3f++/nFj9KfIFNOHqrQdWvNNSbqRQGG5Htb
TajMljHK9Z+4DTmEC18/qf2BjdXafusRwvIWw2TQ/tzzjpN9XzcD71yzPo0u
HTAmpYG7BRroDX7achUmS4savGL50/skgr8lj2dDqDlRCN5A7c+EWMb3XTpm
mbf08PM8L7R9eh8mqBPflLxxX/TZNKcMV0ouDeWi1GS24v0BfFsA0zdhJykR
otxe56qu872IHLs2Mlki3wnvsZQFEDynarAX712IAg+4JxKnuwpUOZqiOoUY
9NYF1/9UtzNF9VhmpeCxmpUTL9m6wk2g35YjGqdN2W6deqtP0i+DyLb+MAJO
LRF6V4y6m1jOHNvR/wJg4v21qBaUxfO8OzIQ0zlq0mdu/L4UYnOSUU4vexWi
bud8OWwhjsKa+eiiky4nwyojnZ4+5ipi8qpmrYS4Q29SYcERHKMwLhwbZZft
fjYAW0+SdR+fp84b0ma9QopZlgKSzkdXUnPY5SxHQ3prU4Fz2nn1cpjh0ljM
ZoGawlK1dkkfBsqApI3iKphNuotAv0nXW7asa6ib0Jtd/O/CljpPXa34g4xr
Qbn32g/SNuKSWWBe905/KKurRD+rXrgEgH6GZvqTqDiYXxPqzTthFxE7URco
PrIu8tAiMLRwgLicIAYp4TxPyId4uqCzTGBzDl0uupSMuG+faGOrx6uiBsHu
OjGPF8FGHN5LykJWME13XK2Mpf37bFLQobdOzrDApMeONUh2Z/4L93BSfjFU
oo4wccVLKZQDrZ+YV5jQu1n6r2JQLgw5USyBHHb04HMTwaXmTumVzTP+uNns
nFrGvb76/F4pYNEe3VBRMmtQrXsaSIHEnuvtoiOnQX10TJZhws+1NSEiXwli
VDR/Ah3vEgm3RhwBLQjEvCzXZWE6KIfYjBQg7zdeOcIQsE3EOgls3nl5z1Ew
t9VQUCeeXLYiJjQ1160xduBjqSO78pwc9dLl5LmQMhWYtqDHExHYoPaCKRq/
eJmgkMNW+W1Yj97rXX+p6BpRS4pyIizrFmGUrRDrupngFUkhTxJSDlonMIP+
gf5HCXlgvG5fbIKBzpIXa+sJ/e/kxP3UdYS3TJ9+C4VLdF77Q82oSPtfkqG3
ZyCU3a1pmFcMKMgrckwq84yLuSrM/sIInuToaV9AwVG0nE4SIU+bE2nBK6B6
wlO1fboTHE7PmST537SC18hflgnUT1f57wPY3XcAryJaVgVrI1zEZr2BtNy6
IyK08PVSOhWEBJk0GWbD/pFNIZfOmVL+J8xv0OI5w2BuWRaDYQYYKwJR59db
MAMd6AbZA7djcjEQrLmEk7LSN90lgTHvezie4gg8x9nkOJ7TSZks9+rS70jo
EUysZpxQ8UlqhjKYFJp+J26HXh5UZcgZsQldjdJqKkkVExW8W5VBTyL3R/9i
mAJILrSWYpf66UX80TSv173AOxc5YTZlwfNvveOuki0y9OTp1+dXy36pyDks
6gMNtrBlNZk8QaiaxWkIu5lQ3FbzQweJxnIU926QpCMgwZ9z9N5i3tMpKOPA
98CEt76rj5k3PUy9fS+Xix3EKbEc3V5hNg84I+Abn88v1zFXKW2tt5fTBqW9
pDkIDZk+eSaujkcGWbi5FffdXY9pf+6vITAL1XPM3gDZyqX/OAC1rVHOSUli
P/RPwcl36w3H9VNSRlW9XhOzliHiC7tR8XucFTDFg2UqeZwVcmRW+2qe8hlz
nkCg2HHIhUU3WbTghIQL77g2GFYGWrrQfcq937Yszr/J/vWloMrJatKRs83I
EasZFnB333fQkphPzUkybE7uBIvDRWyTPNOFHf8JN2zgP9I7OVTW0Nyev+tf
BFcRvd8KVUdHSOnfQb4WKpRY05NzLPfFHvj1Xlla0SyoSWNHSuaFdn9PQGCB
mphFkitcccqGG3zX2PPNyJEJddMJQn/56aeQ9CZe4Cci03m808YZ4GmFdb7n
FMeDXJPNiAD6Ao1Bebf28TnjsGIni70sq2TY14QHCg7HT9sc1lLiIrzG5ows
AGeE/Nk7zIOfIJZKFfb0o4hpttlg5BVFzVUZfKm9TYG/jNWjoMdBKrCvvqwl
o3V1/DK261MWhXJVZbbygeEPogDuNgtcdLmsgss1d74Hv8uh1CEWRvIHTAoO
irFW0In9rms8TFP48ba6OCdrkqeANif0fyLrCooausyJyuuWwYnOnQFHNeHh
4oM5uDrgQWpxBDsHOEv4NGETYTB2MGa6eBPoggS4ITN1DTm/JUbp+P7ZdnVq
2FIHm8S8c6Nd7NkXDZSoVXxSLApwiYwt9uBIN/NA7j1bctijWNTtY6wHR54w
K+5uNR2wiMgKY9bmRR/mTwaNMFqfZEHe59ZOEAfOCRAVDeB+bj6fjVc5u49B
HY+mF8fdxCfU2uPf3qBYehzLJ4o2zhAxLjlBVwU7zvHk4NiSY7wN44Fgta5x
qL/Zy6UJ5NLISwxCoSaaRL3DveDOKUSvGZddT/picg7Qz5KOiDFwE1EWu1g8
5pl6bUzqrecdz8MxvUXJx3DlVqfT3MsgYx8VvrNVlH2gBq+fXjhH4WZ3YwfI
2ob6BraNqpNixQ6o6TQQXSBE7tEPKUXGnR+TPRqV8eOrOgRnddn4RNVIKkcZ
phpuc+8Ky/k+DmS+PMnJfwXf+z3qtWWOYykX6fk269jiaBodu57m+nSQvgSO
zgNv3windRIE9XE81voN0V8hPXyy3BlzvyYzfiLNUpsbfAN+YfGllG4B0VhL
5CNMf6Ev9cVteCE6pkHe/dNNF/8vTSPcWtmqRIS27s1exzUQDyq0QhQhoihg
0LVOoUvona5Ip1j4wEQ5S+nS0gm3uHfHZiMOpPyXb9kO7ruc0qdFprhlEgMq
/R8t/37WnKbJBpq+RwCecQ+IRorkwi7vONSrswlYm+vEJVQ+gI3+fkrgwKRF
65fZPFejfG5fVr+VIwSH7fmONDb9zfnXIwnQqVFnWng9kYZVD6CgqiekqQa6
QbavOIB+xUmdoNIfYckwYJG1YNVZuYWdT6byA8NFqp/7NsykXdZIPUR5/7b0
DuRHc+U0oGdfO8a2vLLV2cn634vEObgkiwV87dGeVSIo78KfjNoxlCUVsiVt
26Bt5QSY7qi9H134Tta0XZ6SzX6Hf6/UDH5R+lVnOwU00MB+aLlnX/4z0GVW
zqYGE0jj7ONMVDq3AVUVS6FWpGLOUqY5Qwp8+7xgQjFVmubzIx0VlCaGgKNx
FXo3n/YaDa2+n+f7VxHhJoc72AGZwY/pSA8/jRgiyO9lurFCzJCEVwfVkFmL
wwRzOJn0wBOriXPKMA+lWmnecp7LTvyNKdVdfJo6+CIMqe8mr2B6Y3HDNzI3
SJUbWzVzx0n/CCIYCmqAx0ZOLWnPS8ssDGa7dDgclg5RUUCDO09glnY9QPxb
MRkWYHte9P6w1eIBV2VSE69/dqJuhdD2L/mAuk+K83uqroC5Xx8wW6KaG+MR
Y9BhHaG2LC5Irn3nCdYDdrsq0qCJahKWOtIeA5/LqW/IoYebUHJzfOR+asNO
RDwFI83tf0WgaQkBe5WBi1gqYMVeFqs0LbOaQOqbVFZsG2PhksylBhn5GmTg
nWAm9TW7JzFQXvaaS+Ypw/CFLp47skMiLPztmziWRL0gqLXQjGBuQXJMztSR
+K5o2B/BD1T7w5Q0ChuGcQp/h8CgM/LrQrX6rtF86KotCiMW56NAniufPA3Q
fBuXnFpkwG/APG/cFw5dtdd0xss8Lb14WhLYlbTWbe8elfYd8t2UbDG0afX3
bzZWhpTw3062Spma2VHS60cVZO75xP/h9DD9X2MaAgfvyiXI4ovqmPBWrLzO
F4QP/aDK8YBrkT74ksf4fe/I8z9+zJmfei48VXKh5cfXTHRZAIvx45Bl0MEa
JJWu7VvFj4g605yxdQFUU2mj9K6fRcAwKbUt7GnutUo8ktfZktj0YIgx7+Ap
Yd3ZNHod0G2Y0v4nYQErZIWuNh3B08VKNAltnpfg6HvjW3U0veumC6ZWjSlP
8u9J9VriczyaGpCGAEVAw5qIcOsvWvUjUlJzhY3JbC2zihkuFDKpQe6WVVmE
3y8aiZJ/If+9LWx52W97XycXc9jMYgsApbQLZHkSsmWWV/de4jrRTqK1Liiu
/uF2Z2acPfpPu8NHKjhvSvVy6qKjgtrsUYKlNdJ+eEftXCvoINGxr6k3ORQ9
c/TMIlBX3xVNfeFTEiPZBtES1rohtIXITpDZhtDerZM8lxiIxNaduCZT5wO7
SMEps6/mcQqZ54LLdwkdOwLnGEC3qCZMyow/uvAtxwF4CgMm9M+XiYIpKjlJ
+WAn4zGKYjVNh/1OExT35/p5BD+aPb3POJNcdDF+IvSw803mqPViJ+DQseJz
rIvVU8gFxDZJl4otIufwEVx5ohyEaUPQsuUeVUJ1FyrpvI8yJ8gdxBMUIer1
Fe1bXsqRYrdQP3fG8He4As547SxHeGmCEY9IHO7EqFniVDN4m3xlZEbv9Vwe
OLp9u75UhWwD+5xMA4eyD05KF/Oq6GySWL6J2mq5VPd4A8iGPn1KRxT8ZAXe
S9gYZ3MdAsKNX0Azijxz8nRa+H/7ghE+BHWwuAv24Aj6jrUCh4W/naStSjDk
d0vjYtRolkj3awWPW1/qd/P1Vp/bTk8USZ9gMK4MEV0bbazVgc5cXXPh6Tcb
0NrH70YEFHggRk9qeCwA0vfoiTejAJQX2dg6ZdMyeVGFtzYil6VurzJJWy/P
t+SNzUKnZu8aEmzF2G6ureddPXpScyOWlWpBALYOTUlRQnRZn+LkxGN1wjZD
uzvpBtoJjAydwznY7UNkR68hTipSDeTJI1JyMOtx4ryFButL+ZIKIElUUZyQ
uQseluXG/i6Bzs/8hOWW7SAXJkfeUAT/24oPkZQPn3U27GZ+tCEHojBWrS0l
aATGXaP3rkSnvh2nMMzOutXAf+mQDvROr2tC9+4Z3hAKaVUNxIbsv3U8k64y
XrrDWOZvd4rubtM7GM1vvVhTK1faq8wZJp4St3Xxu0xv0Z1FG7flKlIJk00G
U5WSg9/bgmZljDkGPma4s3B7J5yEVzBYsn7niIAY7y6k9DCqniwiYBWj4p39
ZYhikTZwYJsglGENywzyU3HEbmWAXHXckUhvfr6RZJpMAeWXP2YCt/wtsteq
ZiM3+LYXfyzIToizmGRl4Fv2xU2ZQ8tenGCC93nQusOJhxUs9UrXjWDcr6Bt
bltAlinsowc2YQlBzQFo85EkxtXEQROGuV0l/y26h6bFMbNKBczNxFJ4hhcS
d1t0sRbSOQUNHx+yDmEaHlA40430iQjZXPDvXUEn4WVxaeYeHSbDyhdHfdfX
/eiPNPHoxqjl7ScdU5HajI+24duxdDkq829NRH7aslfep3doTixaf/2dzzjJ
A07et2PaQYC+ZtFP8q98hOPgzFe4cHzk+2KqCDyhVzOQJjw8sKBNajC6DrM4
wirnK30EHzXMtjWuvJUCUGREQ/qA66B2VTfgkBCTcOlSWtzgoHp02XcK1Ovi
AmjotYeY6Ta1m73qP+WwHIMdBEquNDkncbWn5ZhXEeXQFr0ugXEaqmHF6b25
HH1UR8TBDlV1onepQL6Lyjmb/wCnsjYuV6bp4BRowfX49J1IQ5En8a5xkjL3
UBPKc+GRn5PgJO9Wwd3K2YcK4rros0n03YPqRUvXcq+xWDkZt54oWDfEyqRM
yZjZn6GSEHVRMgMUenIH+NTCC7IMmG6vAOGDFST9kFFgNKWOE0H2CNQ8V+Pf
B7usMjpLU+R1bY7hLsslncDOLgJn0qaXuWHzdCWzHuiZYn90dz5CZaMlr7AW
XjMUD1g1vdyq8D1RF7lGqOk9QI7Xq7ywBMTH+68n9MNwdoX/7B6WV2qJvBkP
kdjzSynxU4yQJ6/J7crgidYZhRBAqVQbbmC6T2HQTDYNGk+D2uD5F3CkaU9V
ntZs7hQhxWaXYxl0mbCBoG7HA/ehWrkSE/7dWBrR3FwTlp0APlDHN9nMatKI
2vlqBEHrt47ngetj4idlhoIHs1B2QJPr8obqJUSvFxbkmjq5LVYvGmDetqWR
PvEcw52xUSJiE3rDolxskL6nz6spcWCwq0ZEtSU9mOCwNl33hWJW8uouZrEy
KCdwzgJmvrGzqLjPegJj2ITwtXqC9jbD/JCe5dYqxozyOeY4vML9ZugJvbWJ
13eTijKwEMhV6DqLGJlv8ZaJwsnKVGK6MaOKFuM4oB7Tx20qOWOXpMn+3z9k
g+bbkMXOhtr9yivgLIsvosoc4B2LRZtSFJhIfzTZCmVOoBT8FDO94PxQ8moy
qC9MVjvRNZieAKsFo6QVxsrqLg48SJOwV6VCRMOaXxA+CN3yS+fIj8KXylqk
Vqm6fxIo8YYQSa+/jKIuSHoHDBAb0AWBi/ODw/UrmRLufhdHt7gU4kCv96RB
vMdazf4YUR24wNwjGJWZ4wwYs5Ug1g9tM4HhXTQmhg9EzaUEVLnodomL4cmg
VSqZdQWx1dYbjOYIXb0LzWdwvoWrXgTIQqnuCInLNYBiK4XgjH+7Hzc+v6Gj
SWHmqyE56AnRcNG+rPJPAS3mMZVSW1O1yPCi3c6wdwYmqcAs+9uSUz4O3lQf
hRXD4vdlpTlsa/vNdsiZNEjibqQ4dA5qG5H6hSDHpdGT1Td3Y99STxz8ivIF
Xnq0R0wKibM/+FKqIajjkHlBmWUkRWSYPZjxJsZAPUXimx/smiI0WiwmjzMf
ugFx5/T4nOcCLgiu9oZr4Xuko/y3XttRV5GB12xX6Q/f4XM08FacsiKyPHam
5+J/RssaHSHVg6Q5KXstzQUzEMExuyDlaTgeuD4fIIit9PvqSewVepBURBqw
DaEhRkz2aHhv6kQJtYDbCucltOSC9/9cNAxrvYcK6JxSa/kzMplmRCJYNPH7
f+jwGj+4TmhfRtBMU8222k73fLND+lwGsGCMWENivewTLDPngK0lVaOYUbJ+
qBlC7u6pPA+ThJJtUXR6Nv0fjh5dndij2crP5iEJHs+JbgIcruf8M/ggMxOo
J4tEi+RYjjR+Mt3G0eho8qp8MQNEEEY1OWqMiNaHOIByMvMZ8yviSnZPCR9J
Fy1HSnTqI3UjR/Wb1VdV9ejGVBWJs9ELeh3CbhrU9JRjEQzNyz0E6Q8cPocu
Rxh9xYYA81FRD2EohSGqgDfAPsK4k/3IstlcZRh5/tXWo3TVbBuUAeLdJZvA
6YmzA9jw5kSnu6qdvd3hlg1EotpUw2oNG6Ip6V4blLbX+Y6onxZQZZQON7KX
u7IIU1CFNJ/ej+GOlrXTwI3MCn7WiBh4F+b1UOboevigcFYag7nTrga29CSa
jHNRb/52p3Jxm5Kj0nANb2msGnh/hjAU0AmxnvyKNvuu+QbK64Pa6xMg5pTW
zNmXWQgmkIIe4eJrwE/JPcveJ5y8cxAMrDf8ibHPuxxtqE1npf6L67tl1ZH6
yb+ygLQFm55lN4r57g+LgIbECz77wNmwSyM9hMlXvxPXrRRCaPzAJ+pt7UuJ
aA3iG0jzLJU3MARTzf/tlFHARoyAW5DYUS4CkacIny+TIg9wJmLDqk4JhAjD
1mZcEuDM1npoJbJKy00+z4C94jRRVv8Ikg/4FnOFRix05rO8DvtAR9RpYqBU
wbK+N2u2gvOWjxSAqkLP1R7LhfIXPn/Qfvrekv4/0PM4zJMLmABUGOKd7GmJ
3QrYJ+3DAel/YZ0XsXcMtOZ5HIJ0bh8NUpgEaZrAkQlduwdi6st8NYyI/juD
nhkprqM1UcVUptPiej9FLDgpBTvteDBiwBO32EhcREtvnVwSXxC6zrpBil56
vrYDtxgQ6k3XrRuxEvKu9Pd9H7eMg+neB9zCT5EJA3G5E5fgx4UiVijZP6QD
tsPUNB4QTDKJC6xaJ5UbkMy0ttFXiqAuaYcmicczbsu4aR78i2EBvn6g1O0F
QA+mbjLxAWWcQD7fzp4BFmuK0JmStgQkYl+EnX6wCN/IZdJsG39AqZhWg+SO
HIGQKvUUu1OI1Tyj7i08QB8IWZLubr54xlJLY/eTnQojRMqVENDGSisDl1aM
4KwKIGrsCAUXalCQMRN5cxsrn2P3OXzBeSoEqnRx2Xx61oZVEqwBOG3jyqLH
+b/g4fUBIzGB3CKNlaS7+yA1RpAPr3JE2nIfoIY8lCq5l77dxvGbF3qFl36E
oqsPphV/lRc3a85yb6zJGpWDvIwQrjqb7vlrHZiDv5dbxw17Dmh5/x9HvDsM
XDIbouhAwtFEGxlOiMmUajhYVindTV3Tt0Ug+xtm49mQzNuCosSW9JNW8VPW
szmEDnS8ivocLKdJn+2AMQeXg3lNNWsjRcfrBwEEQtxhRgeCwPF2LzfJO78B
FBnHFI6mJ5f0MDirSwzlg+XuLnOAWGxLBtf2lDrS/GDiICKdYsKVIxqoAmub
T2zFRY9Wxo8gw+aldQbZPZ5DNougT5RShCPJJnbH+EcAow1ciUY0zXxFW7A3
GLBc+YxizDeLYZ/7ImUeWRubFyaalL8SkZ8V600ELY2p8oCOuzT6TE2IAcr7
RNN03RJyUyCEzqyAScJlwSn751CdPbzzcmX+qiIQQI56YaT9BF83ORjPMYsR
Wog3rwbQ5YBqUraXoUuBwgj/ZAqkVVpG/IW5kM3OTLkgERJIJjCCzZm5ziZf
iNP7JGTyF69fjePRsk27s5Qjjp04AyUiPV4Tzn6Bhqb0iBEJXWnL7ShJqUau
x428rZRlAteAcoW12y4rK0Mzt+/VkR1QvFiQjlxFqwI/5a4j6mr0bDkcbz6s
zAAwNh+g4x5yhQwAcCFEsd1k+uzT5eHG+VKNay6QcMcWX/NOJBkm22k+Ek0p
iYtlKjNG6dxAHE4G0hkK/mv1Hyfc4BjXvdDIDurg0XJ7QnTszTNkOpb1/5mQ
UyZLBsKtnKh1JkIJ+6VwkvUWandFJyGMHOyPHOAhB55072DbW+bo4a5mfeFl
8e2MSLqJFoLB+sB9+Fbe8ZuVpHiMOjjHfoCArdU0/vo78XN0IxeKrCpMrgRd
y2I0N6z/UkY3F44CKHEDZ0b7aUaQ4S9NJtcBgJNe+R066OTqx1eoMJzAPJmW
tH0NbTsJXy8Cblfu4CdE2h6wadVIutrCqcZS7L4ApTlyRfoAC6fhH4K5EeRT
7g28CW41qFvfiDKXFrwP1Wt4SzZd5fJJKfh3wX2dSq2F9T1ZETZRoKxFljaP
pxBeVmR4nHoOzKgOeQNW0gkpLU+rx8RphZ3y/bYGn+0ck9rFIDT0FrnZOyDi
vhWmSbloamv2GiTGWmDxPG6jN2pfLbYPgX6FNvqAxtQEgG8xTKfJjM8D6Rbz
+pllS6NB64k9gCEEywf1UEPVguKGWr4s3tCC1gBS0NaHMym2R8+cjYelV4Dj
Mk/mIzlxmzBRk9pfaGSUZUkSc7ffYy1LHVKf19hv15nOIiisI7VsCdXtVLYm
1KaD+GudG6tT1NaBWiI6YL95dYiWMb4hhmkSGZwQiDNAw97YVIzPEsuqCo8X
BxhQgcfnW/oCa2lqRmIozhNilMNP9mjpu+t4T/MDpdcG/avGmJNcb/DHR6aq
g86RtEBmesgQokE7eRUq5+Qg3WnRxYoRERLIZqvdnLfjfoZbEPe3lbFEUHX+
r1rMHBYgwSZBIiFqfIgNyCk8aXh1AgXascukiFEcABx4+gawSlfeFJOVNF6m
PkpV2IbnRHp5E0crJGTjz6wDwP67B8IXYNF+dYim8MssRM8Jdu9Q4D/HeQCl
l/YRFjiIo8guJTAuwZTQMPDw4b1ojwW1PwzfLs7PAdE14r4v0AvNYKsNYWU6
jo/pp2N0uH4xL73kMDM+Hz905Gcn33O+vukHEuV0WN6YC3GY9Av3e+/zbRWt
LuI9nnsEJmyUW/SRvqMgg9hIOmieXjke3UVKemfyeZJQ6wlyXMcZP33MVQCX
blqLMdeUqwKySJGAqw9+yEl5MUvEf0lap3YjZWtz1frP9TxVsZsclNRX/BEu
LOl6ZR+kRWSdvQRShnMQPryjugPP7VnuONZofgCgYhO4gNQ1RFZMkMEQ5t/A
B1a8cHenyuyOZ9QXeE09bN8WYUH+bobAIPU/tUDN260zzXDI3GY69XoSSvjD
cxILae2gYRTXuSfJ6ssqQM+iuVZEXa4/kMti7D+h+ue33muSOqHv31QuJ3ko
skR0CJv/W8Y9pLZsNTk1nPorbf6hSXH8D9JwKfClJqL5vZxDok8UH4GbhYPh
FYQjxDmSB1inJRWRlhywxkbgHuKKlocdAsPMZRhN//ImWLi8rirsvEVk5Udr
tK6Yc7bseGvhVmeHloc9WOaAIi0mJmlVtg2Q3dDgxaSFKiCeBDt651fPyoVM
PUa+uMF1cKVDWO1mbPm/nYX7WZBy6sz1bGZu2PQvIh4ncNTBJh7yORA1mCx5
glucl+4kMszdO4anLhhtgHHW1RMTS7/OuptHgB4TaCK6e/2Pyd9mm4RG932Z
ryu/7c0rAsSpt4XE/PCSbyDXEp1tiaJY+3P7wDkH7MtmX0FjebFg4dG9R0GA
G8nZ7pAin2bXcxJns/yPMLc7N1weelOEqQ2WKjXqDXkabKkZVpZDBX4iwbeK
khrhVQ/A2wGUQjUy/ehRrK70tKZR1Xioy66QtkUFhpmh6pxdX4vl1gS/T4SG
invThDwsqWm6L3DRveYzwNeYugO8jz5EUl0bxxnJFN9na3Yhwub0pOmHoN9w
JBsWQmrRRJG6LIao4bpkT2zJsMPN8zjjxkztpv0VRcByX9p3fVxXiDVHXtK6
s3bwh6MHXWE7dUuSehlzwtgcBNUwh2o+k0rtW5wDYted4xP8pOfPIyG433c/
MUtPr0jJN7yS1sC39sg7/OIgcnhnE4g/at6qIwzYswAYNrnGhC76pixDDT0x
1BPDMr18cgzCCXlewKNfg4mkYytXBF+9udyEcRx4UFFcYoMziTtohOMoXNqT
QGSisHf+KysUYSEhSQr1/09Awzos1ZK5OWxOvCVfB9rCGLmJoUhOAre+8MOd
6xsekjmQFTgYV0Xya6EifeSbWITp3brR92Gm3R5hrmA4h95gFc0/R/ksuFzX
Pb4iHc/+rtnGNInK06j05I5Y2y4IobD8xv87/Zg4gYlJ2E/9LO2Tn+fCRM7U
/OUIFoCf0KqdQRII7wXpWtW1+HHjy+f6MqVmfO8iKtz0sn8Bz3LylVR76dAo
kbS6rZSz7vRCQ53sjpt9EyljwhoCMX0q+gp5Zdrb4oC2I8DDKIGeaHFCGQcT
F/bViCTo17IcEFFOYMM3Hr6V7swvbYkeZV3ZRYuteBbV7gkjqUQ6FZ5wg2dC
7SWftekQ3Y2S7LpwqiJNgVmrU5QlheyD7KUyCBtX6Ek+OqtyEfJUXv5+PUcB
sjlAgk2FrsO0hbghXFJzzBSFwA0+vw4EkTMQghpzqq4sj+xjC3u80IpcQuzl
KbkBdvb4PY2kiscmrKUJoMbYPgJxj9KevvS3x4Ws6GUznwrHwjUhbvEMT1dZ
pk/ZVOHP2hYZwQK3qhkQQaKfjDNi8rO7YNvB6Qfqe/InvtcsWlyDT2fnve0i
wmS+Zg6NGZ+8WZZf42rof3Aggz+6c+TELxL47lsqamfZ9QvgmLxpoVFgHeXw
p8riVlqjcFAFRjOl0Oj9K0KSqkMpUhLEURWwjCaOvA6aD2so9jSFjmd17I62
CMcvCEXR3lmeSD/EJYqRdqvAGYmmFVqlulRGyJL//ijaAcDHKBBuFRzKlI2I
JbLUGQmSkFnjHhWjYO7pq+iJ0YYZp2vh89y+SnquETf3E9FZckFOyjY9fgkw
vbBtfIGMWlsFup0ZQKFa1xJFfY28uuo1rSoH3dWn3MM5oXTlwuEgLRMJ6zGe
vaJRPmBm8Sqac6eOHvm8LDD7ZXOa+DhmqtTNtblsk6nkuZI9uTLaT6DKJdT7
ilrXq3Nck17VVlBu6o4Mk7MYy24MbyQZ25mT2KuU44B3ZlKQ6HBm5jlSG0Vu
ABmlARprmajBgHBq3PfQMdhO9xD6z6Lfgb1zvcdc9ermglqHSkj3CEBf3/Xv
8mGEGE/qMIy8xmXN/rZOKvk31pQjIpsQtw4fNWgL8CCbYmDkKAx7+8xjgwXn
oAX+8dBkWC3fi+9k5ocLyyWoSY3DuJT1yS+g5j4o6W4AR6Lc7H1WkcSpQ3wl
l2XYae6eHa+2VhcT54yycdUNmFVI7XcUTD56McF0qT4UIpKJrrVoK2i4DIAm
/n9WeVemSHtfjSIYmK+5x6c9aY5w6wzhNr07EVg5lmzcOHXiJRUmscvPy1Sk
rbw2OkcsMFEeAxUndpjyx1VR2Fuzz0YxxrHAscqY2u5cncbvT37cmeKIPf3q
mgQ4EnOA4HJC6q3FAjgpdcicK0ZSqR/oM0beySQAgHknvknKehiIoueScx0F
cvZYO2weLzPjx7Z0zL7tcbWRukqobmVjkarzGuaawDPas6jxFrTszsNZxTqZ
eK/scCLKVE60zsz+cMau+DBvJIjLwpXT5wZIlr8Y05AevzaBJVfRB8kjltWM
KW9wK9F/MM7mUQZmQXIjuET8sJ/ZcTKvUwafed1X8XlGAXd7vIZUjetfnNHG
sV/sfmzBF4wd7y6gLh1w0lW+BCh6gbyxz+uoU9FMCW6tqjTTxJyn1Xx0rhaO
T+m3k9Rtz8lTmxJmcG9i+UBxrYrnVGmOL1TXurQRb83POfXhi6Rqxr9c3PbX
qOFuZwphokt6ADVLtqH9Cl1d0Qzoft7Ll190gaUrsXw0DhsIQErl36lJJf3R
fikfndkTFwghIkR2cd2vHKtVJFpPvAVwoHJSsHT8rDvcQfJbPUQeitSXgj+k
PuHDxngnmxMXnTt76HEljeeNuG5tFQryqxm9yzz56PQu7LLDPvdUF/M15T8s
oqpZXepUECGyYGmNYndvai9g0CIJWfO2KQXHbC9+VL6h8sQu6rij2tB4Nu3V
Su0mQKpOAv61mBeVzsylWE/dG7w2cP3fqifsCSwqtSL7KMY2IXCA6onwMKY0
+Rsb1pDrcVQz6NiOHzDJwI7EnlNQL3SZZ0nKCzrZIn/Bbw/gNdRgSbTSTapl
D3vaEollwCnh0nHSBhFLDvoYVH1Z1l3lcUf1qU6N2RDZIC83j+Cm6B1ui6hm
LaLvutygIc+P11gXR1U5C03NBwjpVzYRRRc6ewqRr44y6oy/JAQyB3XTWukx
XZYTwmrBo1Ix6h4XBoF59zPIrsnbzkyfomblAGaIf7HodM7BxawCIlZjaCX0
8zBZmEEKs8o5tBkydOQCp19IQRvdkD9fOyOIbbhQOOiglz2Jjb8FvabTUd76
2mFb7dc5iGq2/jftEKwJejRtT3RjP2LPWKmEUo8Ji8n8zxMFJfy+hTvhbUqj
dbRhk/7ef9qpYXrXMHqueLHvLjtPnyt/gf+6M0yukv22KWtvMKQeaYOCtfdi
cXI1HT/c9Wr/xu4ysDcp4nRgYof8JFS2nJmKGnX/58kA1Ipdo1HNJabg+c9e
jb4eoZkPm2PHJ6zJHiWN8ws7KeN+bzkST6RcpsslFvR4Hv5hBF3kd6udjUSq
mJxl7Fygp0bQ7Y5uVFyJTXRX8Dh0w6bKp/m/pPL3nBqtPUFCHbqGR/k5I5pt
l/ra48XM8p0E3ToVI0R2HuUnd8zRGD2N8K6BgQtRmU2/Oby7bGFPJXsqxhSG
4JYTckma1+/POCdSowZPKXnYB/yPx0dtiWvUedXGc4p5IVOQDLW16SuwK1C5
p4YtRzWXgtF7FEBdEJxlOj+WetNtO7Ty8aptAJYg1JMl3umPUVTO89cOqryt
HhCSOEH6X3juaK0FHx5OMFnWQ+2h5UJ7Kg+FHHRmYu3cPwY7X0tdOxPJiDRT
i+WIkGG70nLzJk6ZRlNqLfnatj9u8DK6NxROO4/1u2ld28eFVrBDg8xioE5f
DLAGXv2ecyySIzRctTTxaLhUaGPmpl76PJ2x12jQVkNnyTdjPzeZfUGwpvo1
OPeahCB9umAZaHLSMJyWXmowoyqKt8kCM2Xt/j3sWdRm2LfbtpojQPQpaDEf
AYquH6PMsBhtp0NhtjcBFyRXPhciKQU7+15WEhKADWd8LeGR2XRbpsyzxGJv
hWHqs+saFluyCMOQJNirP+Ko7ETfp/OF/M4swLbMdr/SKmHCK15prbqeYIht
y71kwv+ilYFMRg0kqV/T1Nob7NHLh2/FQhPzm4v9lTuhkGmXdPS5o/Sv7U22
tVjnUNmzLX4QgXFy5pNTRcLOOkKIArAyFOsyC2eNAIKzJgNYvFjvqsoCYuEQ
yHI1B83bhJCghaWlNFkYUVSgvPmA06goIRe/P3tnOXfWbOuDejBgM/RiW5ot
FVIBaBOK/NHaJFT6r2YDgsUxA3xv9XIguYVKZxY71pcl14STTQwKX54ByUSc
dHPi4tNts3+FO0Yl0ZAebhGxsSNMEW5z2ciN7JzQknnjyNxXH4HEkIVtN9qq
fI+vH/tGqscKDjb5uK/CRjdfpmFFwYEPUDFz5192y0HOxeXDt1L3mLZaGTHC
AWBkCWf48KhjnRF5Jyc4gP2T/FqKMgVW1ufIyHVMDHIOvHECSpxdfky+/Xyf
97VEM0CO6GCY5J4XXyEhT7SEFHeQcEgLVh8w6rH4+8pozOa2amAi5QHJSPgQ
HJ7yvzUOu/F042D791XnUFBptT/10u7iv/4MfY75iL7F673wF/dyr2JQNGZU
q0aAEITb0zf/gTV5yKaBRqqpvB95mPx7jyvBAvZRhme4KHpwxAekrS9BNMaH
SKkz4vCcgfplFWFYEnMs/T5YO9ACBKMSS0Jl8hDEWc2lVgcCRtJcbPDFy8eg
BDnab3CLAKkLpO+u5xSVP/l9Eq1pZR4yPk8bh8kXmJBbfK1Z4IczFvPVCqEs
jGT0oapd9veybDCwhurPMSUXSkXPskdH/1tUQbmBz3fO9bHhEj0ZR7HWY02J
7YYM4R3j9RINAIyT2u8z5ccjPrQvOawWY5xqTcDXzuxwBsvV499xibrHeRqn
prktFtcqYAwG0QovxjVw8FSiMFqO2D/xvMPqvq1KalgN7FfohQ4xtobl8cWy
j+Htk/EGa7tNliPprLdHt5+4pv5Yd+pRm1p6VQSeuTwlVXmzgFsChEKRvtbi
AVQFRR6DyhkvlH4/hV5vjC95l5wYJOISrqCKPEhVic4Siy9OiFnii7rCWu2a
XNw+Gr6jnFZBftw2Ylvn0oX1P/9pF/PS+p8qdyQyArks77eWGlPGsi3m0n6U
JkxSz3IVfdYkhVoRoNjm+1+MfXV/FrnDlA7YnA1nWJJSrBZfbbITAC8mD2iG
lZSY7itMkkzrO2SOkyaqA56G9o8R5hjWPNr4V9ppijxJwGFst3dRFva5m64+
amORGkNhEL2BWM0tNkXw7jIBLeOQjPJxn5qRFB8pMmz2AjFyIkSY4q38+RST
F/NY53f0DejxJntuXXBY1RnrGf0vBWxUUfG5EGTNK+fF6dhJXgqBJFIpB3c7
bNTyI/ClPsToZyXvAkLqj0KJcEjpCQXJNfAlsPaPRKMv/emzmB1x9aMJ55Un
zAUJM88uTyooVW6GFxVI1tYRInm/1GOvffT/G/V6UV0fMNy4Ic/+v3WC3bbp
mbMfhnirdqSz0rO9Ikz+wBYGDVEaXEHI7xmo8O4+A1pRcl5L9ONKUKhoaIrz
npseJ3Vq0I7TyqfBJhAHaoJOaeaeixT0TOGOSDpi3f5XDee+l+xENxt8aP25
bMCZk21lAcZWe/3fvfhjizUDRa1z0AbERkf7GYOaYB/D70cmbx0iCC3qEPhL
4x+Iih+d44CfjQ/VOjfsUJrZ7AFb8XWRd1FBCR0jj5cvt+nLJN2x01lLnMGm
C4fdtbZnn9kEYUgWEO0X44qGo9F7i4wwHaAHtXqzBv025EE6C3dMpa9F/j1x
fGm//vUI9nS4k1M0TgJzAzU+5NX4NIgCussZ0sZEOunuFs2NP7RI7949mGrH
klVQjvZldg4YEGsEbHii8hA2eHVOWF9jgKlpxT/Hpk6hnzTzuxxsXlmrOrT5
NnRJYEnBxmY1AJGbm6prDCScXzrmeio1OksS+uN/85StBDAmLKYujRO2IOmH
Ue0j/PqCcLIABJmzBDTEWVeR3fxjgOX/1HgL8TMH+sRaYsU/sXwt87NDZzHm
7+nMPfOe8eSPvZxt2DdppME35N+WYrKvv6HDrZb/5k1RLfxT9JCKeCEUlKT9
oH7aTYl3Yz0cWg2w6XdVjm296ylOap3kKI44BvHfsDCAImVu0+hZ/WNTtx6E
hi/IExhe5sUkdOrSuM6/iqCD2n5QiTpwA7aoahjLMBRpnq/L4bbeiTMP0I5U
Ct7ZyaudzZRO2hOOrr0ITmHedhpJ0Kptgryw1SQg2ahO6tL7gptlUK4V5l1O
yDirl6JBqQUltGCOl/ub+jDV6SUmQ4H6N2SJ6P3mqqcasQN8E0FZ5VmOlAhx
354k4Q0YQV48nk48yZd7chpSGzRV8fiMFsOJQTrH9WO2bXc8Eg0oE0/4fddZ
MJJkkxBn+9Rrc/84+eIud/99lABnK6GkKQn8ubETcx0rvwAZ004KtyGf2Hn0
ro1pWSsnrdd/5/S+9Q/0yvfE8RD//H33zwtmYjJDl5csGSbuv9v7uYXKMzUF
1RD8QxHvcBm/O9uKTJyi+tPSZt9GxgJZAgJl2/GOTb0QU0cFm3UhbWhv0sFA
iBjTRzQbyKdsJr+VaZw7ZkcGvabEVZh1DpoR7kiOfwMKQ4v1MF2zv5xewJM2
e2omBq4tnD/rZ5OtpkF0rQFpRXk7sBKjkAGcND4IDHQWhBX/p2jwNl86ndJy
Be0s0ztZeV/HKCLwAEiHMDt5OMeUIIeu+vagfezvEvYCsTtrSQJ2iPTJXNsa
HxtYbhynnJgZiArJUW1J1O/eCMc0uNWxP3YfV8PtRnT671xb2Iav3uA2J1er
hjpr6AB/l+23ghdAcnvIfsEm7GVR92/8O3oisx0ZvMSJNgtLn9evltOxRdv5
bzyZ1G4VN6gJEa5ULVzfHa7B4SJO5UPIrQxSRRLOqECltYLmNX4rnhavHI6X
FQJGt2vXlK1RGSjFfXnqJ109COVKCwNGuBYlK+jyppJmAm3HJ1SMJwzwsp1T
/KE4NLx33YYjaNPQkMsCHQwlb6KRYYy1C6NGBD1kmNDOgMRiL3+ewCgKyXRN
eid2+kc+O9uBchklf6tMDlQDVrXrpX2aWV10C1lMEXpP45PYCm7h5ey7S2Ci
FpggGl6+8vO3syuiHd/ByHbEhiFprZrWyGbCdub/lT4tTIVzWbdvd7kVajA8
wwGMjIGhHgHvjY1O4EmI40yqFP9azVOprZ8zty+K9kHUwogLBBgxo38rGoWC
gmQnbBXNcepQJvfHUjLU5JGBL36R1lbsRnWvW5flhdniZA09jGQPax60j+Ys
x+XfMVtWR3IpELc6m8nROqzFpOYP6i7GSwgkmwTGGvFIpF1OCKOmA12xJW2J
yNAyfkN/7OlRaplpodv2XiPjWWCuOwv0VAbk/AaSDDDIp+sEZhkCWBuU1Lg+
MYbtPUZZGniZ4hVV/Kt76+zhSH8yfK6nqtZE07xBVbomUljVyx1umBMwFAvZ
CnveFJonUwVKBvjThxvfVT75UiqXiWCz56gYOAXmKc3BrFX7RQ04O0+oPg8+
MYcRZOaTcIOyf5/LA7W8arHL4jtaMo8w35QlOKmPFEhBXZ0VX/9C2AnLkD5I
76OUAHM8FRwm6ZxkbA976oTAefSmKtz+wcnmFiJVnyKPV/NtzEzKxDf4oi+P
rht8yMRNJb3cM+ccrBxbitumNL0iSUY/ssq5pzA1a2tlV4zh8dKSy0y/oOPa
o/POApUvvNtbHbnlObQPDQ0akNcFZhxZP1vn66Rfu9qwCA9IYftAs86xWg4J
Fp3syHZyiFGIhuSuJKG1GybwDNmLBAhHKhEz1K3xs4EF+Lrm8DMVIboMCTUJ
GUzN3ahZM8fiuE5o5sCZM/vLgp/lfBnmZvjv7SZVgwssLM6RER+UDBVajdhL
+1AbYjKwX8NuWgxhKbNuw4VWWegArGWmeD2Zreri/vpZnF3kD+qzv6j8WiEy
mX99LnLBRm+kuMa8/GUm5bJH4KnEHiP17Skwfk0Ak3LKrEL0Yj6veewjyQS4
Bkc1LKUNHR//Zzqn8A1RJrAWzgTwPPlzAT35WOlUDP4fTbr/ono3kHxIJzSE
Wrl1b5XX8cjH3KetAWFT/SbDezA5UvRzAyTaur77+swb2CIAtxbB4Miz1jRa
r8L0ZUDfDlt9SrWkTIuH107F+CzEzEvBy5H4isjvikwDZxhIJq1GK/RiugSW
5LHkjQ21Bphzu15nqGrvXwKt8iX465LnhluSU0BhE13YtwpmYaqIdIazytb+
lvz6HBQN7bDONTGWjJPILyNd+x2ovNkoQZqAZBYQjLYXGazHc3MBAhLSbtqL
WPeJHDdk36L2njywh4zyD2rS4/mNTyPmAOFxwXLWEqJv9Dnzd/0vsPWuoJMR
Huql6td7196iB4+yu5KbAgmK52y/buqhiUmyf4hwcwqpz52aDyYzYrACvgtT
/zZ3SI2ZOnBa48yQ5xrvLJD8v/n8raz+NL8VdG5QR95kygK/E8LI5+Myagcc
PT+srJB6dA40Wm2A5d/bErAnXPSTt3+MRXyixu0ICHhlqd4armJGKEzz7u2F
n6d8DCXd9RHpXnP8tF+aoif5++AkslnaVh/FDDCsc6/pYJhlhCErkWImJ0se
QV3Agz9sdR5mzgEaCGmNuCBxiGWsGRh0oF03/I841hseDjnIVS1wN55FtNMR
vBjY6Di50L30BMA7KvJaFuhJO1J7Wu2fWHyr8msVL624bTJQ3g1ilbg4oo5F
wqTFpAGIxqhCbjtfuYis4Jq4S2ugz7FxU14D99GE21boiXBSNvXe2rzNngRq
5dkmPRAmkeIN1Eu8dKoldJX+utuSEVLJrDsTvMarYbh5OzClyF7ixtvMnhW8
CXWLXHZwSfw1IVYg+3xjQL5VK3QAzOwi9Z+l0QxoC2K8loJx65+5WospjVt5
PwJr4dU903GYWvdhYOhbbHjFDfUhthxxyktFZKPSKVy+DlutU1de68RiF8jz
uLN0DmvnJzEdhTWglyc+7wdGrhrWujar42em+qa/LRIxdLLx6xr033OkY61J
J8hGaF8pLs+R2VTJYibe9Zb97l7BFOlk1MjoMaKoDVn9hOWALbIqnnklSfgM
630v/j5wq46+sC/J5QV0LyCqCnjshA4FNETh0YlN39Fm/SIVR1E/8Sa/u09P
glJDOltdbHtOKMs4aTAQgUXEaxLofwfx8jOaJPuNJxP5go4OPfepZ3vkDmoP
opAjg0F1cdKw87i06vsHA3UaULGnM9rrVCnYFvOp33Pt0pdTkqF89FHrCoc4
3ShmKrqkduPeACmZqE/go3BWg3OB/BSkenGpybS/anhoITeX2gGkCpOK9wxA
kY0aNDxyH0lnzwUwO9woahsD5np2JlwG7AexAajhbovfjOZAUg7l+Zkkr+n2
uGL/LXawZvsNJPX9ZT7LbUUGWTAFRNm88H891piRZk489QRlYsqLi3rpE5e7
bJAtgtpAHSp0hkegQ4UgTgly3p4bzXtVfkkTA/kZSh58z2evyrHpraBAN/9g
nDLwQeNuYNd4SkYK2gCrYgWNyXfPWQFWJWw4894veKckyiObPproCn7E+tzm
pS99sjoYjW7iOmwAyWom8jZH+O0SCwYQR7hYnN1Iyb5Ud60dW4DLowsEcnFP
95yqSnmvFJOhU6JJXzFzd4a+Q69taAkF34lL1nTvD/WKEXJpEcZ1u/CP7afK
cjGsPWVQtaNhWt/eqsgwFKplxAr+UVZZjyU63L5UQ7upjFWoPtVfZivRbMKC
wdzr1P9osi1AWG3O//ysZ4SZhuaygBYPAA+3a7+j3vJS1VwdkaAkkZfgCqrF
CNiBBvZQBAIo8UNyf8mg7jQEn0WtKYJrln4MizslD5SvCJGR3kN4GJmGrzGn
aXJYl39Ug+Bpj9Cj1BsqbnC1G86MTlagmClRxLpKqGsg190Ts3vencKIPV8h
Me3RGXFotQSsQkjx2u5SA8QU9j0XKhfqkAkBdaYFRo3hbIze4ifh7pG2aM6a
L5lw1a2INttZIz8m1G1njpG+kZ6T3VCJXpTebJSGs4syoN+PbJGTEi2MsaYi
N9eQGSFR+04ZVQJwdcfF8aQMHbvME+xvwd1BUYnssFhAAVFgAwbKmUT9n6CJ
9carqOhJrKIrLXn7/H8vOdJwCu4c3pjISZuL1N+WLRkkh4g5Jx8HPbJrVrZU
3+Aw63LSdeoW7YYd19m1OxhQ6tAiMMsroNWlz5Kcco1jtkAXq8vewwhgXBAQ
RnEKGRdD4Z/LcYuUK5FqmpS2XVxO54IE4Wtv8oj7ZXl0gV6yrkXaIt82KJCG
nEKD4/pZTndVK5px46CzEsc0iDgg5vtHjoknELBeKlOq7ywILyh/68LyPbbE
+7pCD75AhfzI0wtmZ7XwiwOw1s/AerCAUzw/LwPWPl+i47jdWp/dDstUSBC+
zMcI5mcXzkigF3+AKZSzJjguw8Vk9WhBpkYmFTmOGmmpydkfFQKu+GNzwjkl
c29Qqg3MCQj2hI2Mwx+E9mbK/xHfZmjI6ZA6yhIvUfu/ssg1eI7JxUgC12N3
zL4wEL1sqq9qsg6FKBqan4Q/0hz/CbZzAayqVSgkfGSGHkqQ4N/W7jl4uccg
sxtzSrw+FMH7zF+JxNGGde5ZsZNpEIQWffw48QA6DVnWZQeb9YTtWLUrKVN7
POVITWy3Ze7vfXGIYzllK6q4I267hmoAMsaim8BLghodmILgeIF/iCUtVfMG
yNW+PGFpcKRCq6qYMOkhbDXzi1vzNCR4Y5U3SFk/qk6iuL/AqQi092poNBod
WxzgF6e3A6KHMCpb3kmOGDKbX3B/opuTrORxWzyvNcEvMU9axBNfUZmi4+wl
VeUJJqOe3gEF3UmIgz1tq54sBmHS0L3/V7IRTMPB4fIA9ZOpMN1X8HQvYc0K
hHxPZVutBux9hYO9tglngQMccBnnGs251j4dxYPOmfOwlY3YqAzmi9Yhh+9X
Aqwav5HwyNJKRLyL5K0j3DFe0ZCshT9gRN59r4KZ1x8ANS830mgVEqrsz2Qu
4Q5XAbdZakidgfjH3ANJObPQSUOdS8jyaP3y0WubGB6EHc4ilQ1OSGtOcDT/
1eSK+v6L7q+3MQWnKXhACpq37b1UCq+Ig1gmW0jSGcUR2mlNipQD5UYuokIE
TDzIh7NNmgRLqNOzyBBR89URsg+7MPLomhOxITFcAHs3pmm6ztSooKDzWs31
2hm4xg90uH9QiR/NJ3dlvottLnpfkrDBKKqRj5EnRG8q/n1ZsE5q2Nj+psHt
k2sNcgRIqh3xxktiXv/H11TsX7jWMlxtPnyafkx/4OPHdBPuQf8GYIFgZ2fN
5dVg32hEtXXdVmeJUt7EcVuOVwkeaxyVPwYlHQ78YwQsx5+cmep6uZn63m7X
7A0T4MJ0AB5fZ3y2k3CNLdDQX1XTJqzu6nxpXbm+0+MbqwAbvxKjj+XfI7DH
Bx6umK0OeNyb8cukkrYsliXIYKaYWarDcM4hiD2nLx69dUFqb5J9hGMVPKuR
CeOnQgpSE3wLmtJVgeDxzQwwQaCBiegUVqedcmSGiv6K+SqkwIBy90f7GiB8
cZKLDyHVB2WAXhYMUAnJ3U9NDNZauppC3+qFDKFsyQWhCLgcezRqNrpPVJsv
aAVts2Rxj/MawsImRVvCFsVLTi40YSh76eBFRjtCvOWMfxUBwaMgJs2vievU
e3LpQNkx2TWdGsTbrCDSbwHvbRPzO7I82cEFjthtlAmGis11CSXru4nCFkDy
zCPWX7j0/fEDzyeg8Z1YTRulggtNB5xo+bzeEfDXHVOEwZ/kH44RiBY2PN7f
w8MLydY0SY184afXvjHLXPAud2mHBYENsznd0MozwXmdCictiOXgqkpBC8JW
PiwZClRv4Tc/dP6nypx7JcUbxT8DlCvTOoV/TcWg9fQRe2sacR61UrZ2+j+K
sNkpEyfZ3Nizdm3XVf5feGzQNWT8sjXF/yZrIGrJzTbv/lHTMSpc0apPcnaZ
sxeD8A3vW+Lxq2s8VEWgvVdnwymXsH0LDbXZuEAuSeUYPw6HOCa03NBGJIDM
Up1PUDaJhqV9IR2MSPM5mKWkesAKV0UKmxEcyKRwDE4sgH9u3kOuYv34COuW
Pf/G06gBxAXU3wORkJM6upt215AmdobIPgxvArFfHQycUHLRybq5e8PXBnrp
+p9hLetEjbZB2FDzP5iITKe7xW0Tglt+WYA5t+/cSZVI9uSp1eupAJm0pbMB
RfJGH5ZvoTgG8i5Oz2HtPGFp6MQzQS8gtDVEZGPqjpLaQMR+cryduIr1xQn0
qZbGcHn1OqZbdUidvLclkmxCqFURoor1keP6ATEzlNKQHXZOwt2shetSDCzm
9LGvj5MqaZbTbSmxGfhq4Vr9qox2Eri32C060JQ9dllbDssJTVftJAh2VOKZ
8IC1/JIQDcd+E6+uGs5uM2jdbdvqOTG7/TmPvsGSChVLFMxWgLtPgMDpjtfa
GxCjT/KAvfyVEk5JreyTLDA/lOXQtURdqnNrN7mLpFlImp5CvDVCet7RXa+u
fncgpCvv5e+sKHktpSkPlxhrcZdTjpWrLYYw0YC3nHmA/SJIDYE/4/eCP0MI
M5gLCiqabDeFkKwgB3s10GwHGdcAwi5ddbEHP+/U7vUldXUeTuBSokwKlyxP
LKQrTmBp1RcuYpNuOZI4+0Ly8+uaD19RUxN/ZBcGnmekEzt6kaIOuOg/JcNg
KrhIgT6Jqydf4VUjv34ekuEKZfH73glb5yaNgr1IiwxxPnxEqun5SzR/TUKN
JQlmnGCIsHLBFdr7/QHp0S4EYzTWiJbD0fHHdlM618STg8T0C3O6gDU5j0gW
YFzj9A7dSLmrVGv63eje9o+bGCKkIhcI1NpfybJyoLzW8B8cs3NTmq+TljVN
cM0ARUaB2Vz5Pby/Coe5EnKyYVhLcZYX6Qhjz3ZMROC4U1UoMUQlcXy2j9KK
X6DBvNJ6soWP9oDZASgejXrC3WP3m1gzNJ42NbBLkSooPvbsx0LlZtTcBGvx
RCDerkLhLqiI+7zHCMZaVTaKRjwqKVcXh+xEF6La2CtfOSCQJQzKTk5bdd/b
4rJEIt57oE84qxtIFx3efuhmuEPbR7ya1Co1o5eKHLKVXa6iKj6PkFFVMZIN
K8VLxdLGCKPymFPe56wIa4lxUKZ06FrmkGg1ZbqSip0sMh1m1IUDAsrUcZLx
U8a2iDOoj/vbH44BaJHwDXrRNQ064TXjZ4yx/lmbj7kKxiAxccp107Ze90rM
XQ0INPer4E0Xo6lu59KuhE8BruwgHHT/ELmqNUSZxzJivHR1exfQWCRzgW9D
NOfyg0MuM4jKPzJ2SQbHK+n32DMPZ6xmwKw3wbkmd6xGuNMIGPLKaaknWqVg
wK9nU1cNUblozI3juhcH8t+Te8BTgTIV0hQSRdwbH+tT6gr+BUn+hvL/bCYb
QsCXPCqeDD4RfQEmXWpU8h0elw6J//YG71e9YW980YAW5exy6PgohHTkTRvL
z/pdV5w+Jsbx5hUf4Ieb4TFJ4v8Vav8Tj96kDKKrGGwt0D0fMF4Mie2HY+Et
EGB5ZvSo6Y01lAz6zfd8u6KeMiYN2JJ+nDN+GfPpj821k9VWfvhEvld8QfRB
PyDOG8XuiTzQq+RL+c+/f8GqcZX7lJ1C5ElnwK+3EPVm8qxFFFV+uxC4M7Ab
g2VBlHAoa/1y5DKgGFmfmNJIzk6RhgyLgj42Hxf/WJJDgafnpLUSA7X2jhyA
CB7ld54o7uuzr1X1lUtx86HRr2eXjZLhBXe9noLGvUL5zouVFeWE2l4LBdo3
+oWMdS082jzzSpHeG+LZxcuNINo/3DFJQ30SpZ2NYZ0BEB/2n+R4x7PaG095
vL/hK8OFIZBxEzrWC8Tck4ZdLZNPSZYYgBLiUW7grJeaWIJhbTACXRY0LuW1
tArqdLytSt2seQCegkOmaCKCL7nap4ssjCfSdaXGq0bdz3vWNcG41xrXE0Fn
yMaYjEkB0cV4nOnn4qAVd/sIf7ip+++aQqZl6XBtg5fznibVixE6fNBEYXRp
NMBcUNs5B2WWyVNQCBWZFadcAtit/xBpp9xSS0kODUOMG6yjfYqcM7WF5YFg
VRlkpB/JV9OJY8/SBwfL7zx0qo0gzZrKMCXyMK6EiYXdnAqooxhmgbB+/6mY
FB66iCG6JsythRNdDz+FV7T+rWrlOrWn+mV5Zz+NWajHRzAJnSY2RoS+5aA/
+DWRt2t9KSLpEdgfgqeWGfi7/eeJNhp0HfZlUKgfqcgrx6CAm5XW1or/VFTd
VCXtQPcr5Wc7pJU8B3fffd3rMfGvIaF7gASBX4vU+fi0XfWRTSSvgaS+3mQE
ZGD3zu99wI1VhJU3HheFy3m6Da6/Im3ZdwpYJl1CcNwDbNudrm8+aNVZXu+N
k7TSiqT0jQUSXitj/OHUk1ZoDl4y2oO6jCnyrOHMPfSp385zkoWWrOQFe18D
gUKshIE9EDrLjofXBMxySSPtgkHncM8eBPIwCOX13FVZqWjoFIvgKY9WrShI
K2oseuM0BDowc49jLApKbxnZUjNXKT6ioSTK2Q6usDVRdyBn8Bj/9IfUsx1e
aXNtsDvXYW8cihyBpLp6TiRKwm6nmRZBrXO4h4RwzOnA3O8Wvz5wU3T+tuir
apJTnyQ2tHiUIwvidj3xTZAesUAJ5cRjvb4D6lE6+hCfyTx0GZPVht4L0Dk/
Y5B4ZxMYHD18G24PtP3zxfvizyv5XQB3V3Ga/6q7kG+N2Wt6Y/lv8/PjWh2C
bHRTrhnvDC4SmJ8qlp88CFkHHrX6DmJ30PXnBFrF8xx+Bok7GZMJf5IKBu0I
ytM5T8vJe8hOa95mHRx6gSMK9QAPr8DSndNt8StwnaZSKoFMmoh/rztmmB3g
A4gaAdEeE8OGaKqVBjtGxw6Ma8BnLmitrFEqyTBrbZpex//8KSOTe/50sJLc
9q3962TI8W4tBkdlqWOlkRwKaUthDDoEJeOPFf3U9TMLPxB/r3VTVsNwcBsk
lj475J3CTBdR4EQ1tC8taNErZIPdO34qFM3hYkIwiuQffHSYABR+Tk6JEN4f
2vkzqoGGbiVZRQ61ttnPJvozEDGdXuMoxVdJpFuP3d9cF2w6g44Y8F+LmtJN
aUqVCJvEAQbo3MQlk95EpmR4cw6tq7N84DwM8NJf4FYQKOGhuGT4cc1Qj4mZ
AtTTGMSMD19mwo7YXKLWkTTH8lKkc2342ffiBesmUuEGb4pUAfX7oAVwDs0c
CJhrujYNG9TVO+r9mmjBDo30vcYMjXsatrkDriOLxC8ogOLHMuC1vO8+wlTh
JWwIUqS40hSYkhx+mLjPUuLBc4kULAIbWdAfz2Xe48uPWdzGanQ3q8J8/4gr
encEkxqG7NJIr4NJD7I5oUfTd1FNGIvCKZg1YgqoDFsxYDN0Gif5btHoeHAr
r/aTghB8+2XDtG+Qsl1xlLoar7KL9KWmlxS2pun0dTlARhINhFSdWSnGKvTN
NkP13/YKaCu+asZyRHMPq1buTMB/n61ihjM3ct4a9NsCGl84xgK807BmKwcG
wAKfFQ3M15+vAIY9bcSZxEOEiG5t0OZrBAjXjpMKlLql9EkZsKd0lcqt0jqo
96ss8EZcbQI3EU+SN5a/IAaQ6/8VZ3djGRu1u5yLo4+q/AhB82v3Kg3GLdnf
s1A71Cw5tCg9ZUJPjdnLeBh5TkVd2om5qF+itOSAdFZpkIDL08VGChqooaa4
2BY0WYRdG1aW641UQU7+bFVrw+yHaE8oCjthDqeZVE66w0TOq6m3lP93uiq0
brMVkMAys5MzfLRtyryabusDVs3CtbYNOO2vUiCtS+gDR8xj6oDzsxuGrLKb
yq3dGJpdF64PS9DMmwKaAk+bJJgdF0te7F+9si0LkgBSgQnHvM1LNGqE/Nql
hVZhfwNNBYQlT0iHM9eYzi/X8rKoGVhpI/g/M3rh24TR2zp++XwtsQuy3ttT
LPJ8Uk+mN4uV+Wowf0wBa+/Xhm93P3fEjvuBkkV351jIb6FWFW8ZSVaor7Tn
cA6hhzEb2e8aKCVl+jHZxhpXxnbuQwmP7ffR8R+rzorjgCXIlzotA9Fz3Hzt
dwrI44N0UYKqfh3QCh1KElONSHGvO66CuN1uID+8GYKR7hUeiBJXCMkRCWrQ
0WkjODImlUlViApnnvZeMlfyDy4lzxCni2BA2m4JlAUcyCCJTPgQg6OOVeVG
ylfhMWSLonyc459x0R/rNgjP91UIbQMwjpD/wiJ5rJrrLYVKuRSZoFT00HFd
CC5OFsgcH4VupePThjbAqmUbGOxD4ypj5r+L/lScJ7f4VWjGx2v0HmK5Cdt0
bb1+bOvgfAd9A31AnGbeny4N7hFU6x5fy6QWHXeHgWZNOo1xBM8RTYxnDri7
sMJHNeoX9Kwu3e/1wRbzXBnVCqrllFU6H4n9Sbq9oht/feGJNxyISTJTzBqx
g8GHz7X1GFg+ZiZhT6O3hIfEwKkac2OriBiaYwYJYhnKy0TcoUw12tKZS/dx
u4DzJT8711NJ4tEnvxBUcVfogzrEB7GHHFsv3nSP66sbsB++7t7rwq1aUJwd
sqVKXh60lb0xGfgKT4pythM6dUcY6sZWe00vl4XYsDK1275aCQeciiyBellF
z2KxVAeskP4RY00Bbs16pxXjEWbwa7cRTZAO+r4LGBKCEsoAZEdFGU05rfx4
WNswj623OiMOdeeEEa9DXalTgJ9CxnvudlCtUmJGbMuut5y5cJyNUGcz8Ogx
+SyJoETeiZZtIwZWBTpyLTzTfo6uXhonx9x5vLhkSvWMDZG6YKA8yOt8YZyO
l/a9qunIDqdEPJW7z2lb2ZaW75ClyKxy7re/J5qbTV7h8cESK1nEPZ5wi7j2
SWBvrWdexhcvBjYCjVSYqX50hrQC2gq/dPEbqWRJf4hW7hoRsj/mpBDfw4B9
UvwJpNk4xl/AvmRKnZx+bTr8CRC95j+knRFzlkEAlAxaBCgOYx11biPAdIeC
+Vm9q+Yz2VEYpI/e7Xn5g7ffIaVNvdSK6d7MvD7w06Xj7LUEVfNbuKiauyVd
sgm64k5Hc+QFhAnGZvVZL9nigVRxyGvkEE8JGkaMNdbXfTX2mBTuOsfkh07B
eCexSzYdYkv0PuSWcRQ1vJOjGebMNNHsbZm2vS4hSaBOPascUAA9UORqoluR
TXjCM2HX/+2gRhQd9jhIm0xZB20oWRDjqCGDzhWqYymDOwccphveGcJQGQci
ea1IEIsVP5xpWPGhLQ2UdjO3AWwRRwhyeUWTN4QBav3DzicuycKh0UDlP3/j
DX05EkZ3KS9GMrxMzNfvZlBkZVIg3c6A3ifGmxMH4NJbq+J5HszoWmq5wswI
Uxxmx89sZTUPDnv+0Rp2BAAHJcCv1Y9Gy5lDe28tUrt/RjeRu8s8Y1ZMElL1
VR49TfdQn1bjFdf8S15E602mzLE6ORLJe8yuCF3UpijcI2ANkArXVLSTULbq
1szmbntcXG1uE/q+QRwq9hUt2k9nce3w9xEuLX0NcqYw+Cbqyi6dueNHVqns
UtSNjIHoWaoEKYD9q6FaH/wQXpTqEFWXJntBrCRGBbnhFow6xOKfPojhmJOj
PVjvo4CVx490uryqI/fVBhBHckMhtLLLnzMMETKN1izu1brMOQDTilXOD5+n
Ra/30/enrGnwYP5WY54t2G9aVKsIBIIRlXnXvIUoaGnF3C18scsH0vw9MeYP
imxWKxa5ISM20PM3oOh6PP5BLd0DCg/xncx6XRIhAuVbMqTvHBjLgl7zjoCz
IKYuUsaB88hWJW64FlUVEUBMJhAazn1eYt9Du0/qBriXdhXdXSEa5sDEfzKL
KVLx38e0dbuBewcyoQL6BMH4wtcFgzM0QQGqc7I7pDN76fz9H19MUNoeQCAw
m+YvhI0yC24nXnO/0Z5IMVbEPUnVYJCNeTyhGLInNwMPfZLxj6UwPDepU+mw
WQiDWfT/MpVS6TpUyGW1qKL8mRvASp8chQvf+FxIZaTadRAm6SCnhTSTOjJo
UDYDTK0lYt4pAOoda7Yre81dcDQAL5Yy1e9mpRfx2H/7PjjBI3Fc3HIW22nN
xaiuiSac46kq5hJsTQEE17dzbTwLbqk7EPHsUXJz/9s0JZbsS6TYIKf97FCE
mHf1yWt7rI9DmNR9/WXOcDktp7iw0GtXEW0AZu4FmLJD15GGpqeidZX98t12
T0uMDzICzyVY/b+wiREaaF/MMi++UuyrVo/PUP2RpvQHWnsH3GJdK68Dp8r9
qMdMfgRm/V+n5M5XUMsjxPfmwt3xYmTcz2NQmtEFmq7pSg+U3iTD2rF8KavP
AuVOsq4HeXrqBCxgYNBL2s6osk1s57wvRnJHwMsEAJ58/uvfnhZk+HYwWm+f
gNoeQAts0kKSVkfba5HxVTACs9yrivwFQwNT19QZvSI7uC9hA6UEens7QmhE
E++9b6V0VuvkZwrHMLoX4Vh86TCZBOPRSXxBBN+XVkUXq0a757xmRHf1u+bn
g3nXWHbqn8YfMEsFkZTijFGL3iiYnrPN8/o/1d3oJt9Y7E/P34Bgn8PMPqB7
VTwrDTGfjEtncr9hVE6yzC8uhf8teWuWolYfzM5UBnCG8k6ePTDSGhOfUep2
xzmx1lF8wde0qINLgd6M6n1B3PRY/ePj2Bo7OGl6H54Ic9tadnvLoSVMJItG
LblULS/aRs9PKXU26ETxsdHOBK9nhCtZgPOk5NWzFi+W9iyGsjepEBZj2btB
ycHqfLKy6IFlgLJQuK9WNzGMI5X7MJrl49sNGDNtsQD6Y4EtGNELqrdPJg4E
llKIMiZxBnPGEsNVX/tSfOQEWAVwz05Br8SfNSMiK4X+ycgbX0iqKoKo99FR
n+ZhxPP+2Y0FOXm1oBKOmg63SMKvDlFYID2aInlkwDRdF9mvSEKnNQ8AUwUB
1um83ALdtiLZAceFSQOp/XWj3XD1Nevgm8lwlAvdj6JtdiKilw0zAhKwsCsi
Uc9CIUvZ1CZ8mX22uk3i89Wi1KLJS1BPiKQDCU7jwiCIgNzAjAduQXdSO203
QxnU6WI61n7UlASPszOKpCUbjLw5H4OHfdc1jtXFOGttSOJffO7xBjnJ95ez
XpzL2IM6RT98Jy9c5Yhh+3irvTedRiL9khe2wsvF98AT/GyNMM0bw10Yqw8d
fVomKk7PbxrTfLjldsQkW1/VxYFSx+0BN7XsA8ELqW2zk+EjKNptzTnU3bN4
IfcH1wpPm2CSVArl/LFGjbHRgiV1pXyBytDPxLYAOE8d1+gv9QfrVfnT6dlH
Ou58yLx4dVVQ2W02WSOp3+bD+SpUpXer1Wqq0Ozx5c6p9+q8eYbcOBq6OwG7
gVkQKJYjENaODVLS1I7cXeLy2imHvgihmmCeFVTNy9iDoHJ2r4jTwxZGww0F
1rgvAW+TdgtRSwRA1jKbWaXRYTEnMGTIBdmUQcIsVHf6hP/I01bnKUvTzqYU
0671RuhM3nrq28QSsM5s0ZKm4Tj0wYBKUBVJ80u63Zxtt3xp93T6UscLKIv1
3896hfnqu1epec2UqCx/Bg8wexrOFTE30h8Dd6m46LawEM1xd0odAoKmwEfv
U7nE2v6D3RE9LHBwgB2FKpKRXxUBXqRQpFps36C7cuBKB4Fgpt7yCL1s+4//
+crY9MvKszO5RodD5ZKs9rg9ctrBbeHlOW/mF0+2Fmm5x0bl++VErhkFVNnK
EF6iMNZ7j14XtkTshrGCh6sEN1xjLn9pP4cDxB/dxCg6WIhyDvS2SaXP/BpC
1ViOaUB0wq7P2oKvC/8lXydfQtJ1F4UxCbybuIO0juzzXicqE8BWoQJeN5SS
pEwbvmos4tZL1Z5YgUk/tY4x2dU8bMfdRo0QOJfNJ7qSx06UkhWKY4i2W87Z
KBgka/iCC/WDbVx/bG4tBtaFuQs2DqxBYyp060ncoKjuSmxM/0DwfLIO5SkO
wwHhAqQla6NQxuqNwtB9z5t3n2MpRbMIkP33SqsnAZBuvmES3CTZpKD3TvCt
1BDjrkXrWc6dv93uFhFlEM0fr17rVh9UqxquJn/I+uVEE9uh7ij4BqEp3cnf
HEszteaW8JN4ehZQ4sdGuydsH6lFCKON+j4bWJ5rJ7/9Igyq8JgwBT5S81cC
+qNMX/Hmvjx/TxgA9IjEn31RVGF2luKuDhqQp7ued+dwKzcwJdWtBFlm8lin
NTnf0AhntOzKdEALCHBNJ5cJ0Eo0Em62th8ddXJ0hw4dleXQvhkLn2ycrbD4
fGF7dQg/zQp/8GpeU0WBGbIdRVFa47nmShmlYXiHZDaYWZ+GdXaQ52TkuuDR
iGU8L1mLp0RZyd/sXLNZDTwuWjzWUBeUfRB7X6MRR3knWMhYQ1azgqakoOUa
XtXZ952yz1QiWjZIILUcsNLE79WlNSVXVFJnfLR2Yeomd4aMg4Pl079R/rqx
WT/MZdKBD7uTeLrzHnEskmrAiGgvlmYlhl09uhuvm7I0UlRhQ5sJg1ndFb9O
giMgwR5NgnxvBKte2B5MjckgVXvklJooJPtO3jZTuiZpBsq1YgwZT0tJ7Y03
9IxI32BOo4RMvT0NQutqrT/6YkK6cRu17su63BySEQvAnTiLatNF/xr4IM1d
q3MVQRDwFKDNnXml1l2eBBWM7h9qwTaqGcyCsgloqaJwPWX/zuxzZSimxQyH
ZoV/LFbItTZNVvE4WubupSHnwTVK9LDiFNm35fDAJNTCBccrfovLgmQ75dvZ
b/sDpnovnNyURSO9nKoPgrCpCtF6ibWcT5lVUIQbLSoN5vz+Bi5vMfShvhDy
YY/QVP2w67Xh0/t2SyVSXThQ+Y7tcllb50W4FTGkymjU8VxWTCCVXgLp5sWh
YN4JhcvUraesLE4Q+qkju/aiMkEAisSqysXneSXSknbemuzuo7CHi9fUrkQE
ADF0/Ha/f9D4bXwcFl7oTDSseFNtWB3dg0euRdE85bxY0x9wi1TSwA9lyoMh
n/uwFzXCMJ1LuYcX4o9+oFYptzQNQ2TcSwrOaN3YV9s9S519I4i2Dg03DvnT
L2xIQ8z4vRnfwLduUPwq8GIdB3BtDn9SYDdSIhagKpRSo5AYZo3lzfzNI21P
U+ITFvQfZpNnOywmuGyeSw1mvhHW+/ExF/VNHKrdpZk+1KUno0PMCuclmdS/
61O8wYPT6az6mKvjYoAKsKPVSpCdpeOScdqvCB39oQqSqGBYHAPElw9yxLaQ
Rhtw095Kpv6Dr69eZlzrFzPDwQYUEk1TyIt59/DPXl4bVZB7p/W8b5rEYBYf
7XLyJp4JelwI3malvnrnLDXRq7cFScGNn2Xk/Nid5tnqHvcQsHMd0M37RHBw
1CVyTM4Z8p9pSVqgGzK5E/IeV6u2D3AS8cQinHIPUOnWtIUQWxtEyOoFStqZ
g/ssZij8D6Z6JoEG9ghSjwWS092dwiP8g05aqarPRpDMjE0jJQ3Uup2weyrd
squ7eOFrwFRkOdAJuBE9jLAfPGoJfLrk+4z+rwJGn4ahaVfUZqsVmLOtUxzw
/G6qgtVewlEdovfpB4azjTYsV9RvkspEuI6t1lzp1wtQ8GcMhSfnAdrUXp96
PhjnEqTrtPgiA5BTz7ETYcnrpcbrvEv7IONMV8lvuTdRg8pczkq0Gq4xNK3o
3YY8M/i/QZDHO7ID3obsd7sAX7ICSuoZ5rYycTMVI/VfGkjR5JN16EpN6TWe
qcyRneXF7GM25Fgpi0f0jx1+OtJULBPc16BEde9PetzYMlXmA62YZ5eoNrdV
CQlhysrAomKJfYnIXVUfUBDvCQyQIqfATWzCRGw8CT4QJPyDWdPwkwrxTcHj
ieodHCTWNZLJc5IcFtoJ8gj6JQjiVNMaZOq3BER1cGzGaw9m3SmMr8v6YY/F
UDqcMW06oZTl3iHZnD+FCp+OPwvm+7yftcMF5uIMrrIdcDD179FadyVcCMZa
wo4Ada1yhjEuoCEfPt/aKB2eN9OzBG/xyX3on0/mrkyq6XzQLIDZxgXwtSIB
ppV3AXxIYdYVV+weFSiZh7jNAhMCnNYdALZtp5X5RZjxufklvsZTbM8Bomhv
mWGZ0Onf94mNs2+g2wLzNXTVp+rA4y+/aQhGWvRy2Y2imnjgCPT/Q1pMEj7a
pG4roL6brvTegeIIcMdzIT5kmqwqhHoYgaBX9kMAvzH+HPQ0DOrEDqGpJ8GV
8PjsPG+0+qIHVCbuq1xsHkauKIHgK5OrrYiW7Sk75egzwFlhWQN0/pWozZHI
AjGi9Qnw1lMVZSltV690A6gOpjRMrVoaAHqSHciFg6XRj4PDn0Zmb46QSaGp
KHKN/VDmF52zQI0h444afXetm5/dFnMSIIx32VFZaU07M+pEsgM67UT+AMGA
J+OTUu/YJRiFbcGZo481ylmihwghhXQB8xPcVrRoYnUOr1+Uj6Fu0f/c8+JN
pJmaiOtmsFe4Nqb+6lLGCKuehaBtj2bZ3gsVPeagYxK8O/BB9z5PPyb2Zc2n
77uEf7vmbWQ14ryib/q6GGvEsYvQL4EyrlUOt1NkkXYdnWebzH02BGppuZSX
ugU1xbNYD4zE8fuLzauIO2Rt6uva/yVgnJ19iL3S2wd2Z9X0wvH6fq6nGHow
c3/R/fkB0bslB8VOANAKTGVvBYZMvIlO3tJbgTRY5EIJAscJfi5FS3lkE+ha
Vj3G07PkBXgO55P0ki0m4WrVdRc8HQVFg2Jlyv3aeKz1FtE11dgYFYkajBTn
KGQVEYDQh4NBnRjiIcFDsPb42wazAG72Pmyg86E3Vln6JVjaJxCwlwiDZ89n
ggDEhkM+UwZBOjEe/zd93CinC9odXvOr9inB9U6o5pJtX1z7CXwhrArMqZ05
G02xkJHVj4D8a0ctTfSL7nOZuhZYwuCkQl1AAbABiKRO9edJwsk7Tq3eDMM7
PIYnO3y6NlIOX03YrKu98ZmgaCGxN8qLm6xVOpfaiCC0vB9qHdxoY6YQkWqT
mLu5rNrnQc4rLw6YiL/PirDrgdU09Ok/1+Nlrh6WnUIxuvYSkFx2WAhRCEz2
btW55B0+pzoRmPFlxdQq/gIJwGiUa+6CH0/QUumQ8khNVAyLfY/UbNbivjtY
+qUkU7sd38rOOp9eu4RTpeThE8gxO00blDIhsdvnLfVyQpR3DfJcfltSVIqN
qtH8E1Li2dQkYK9MS6pYALctv9X6XTpmGLq1zl9nALxewf7d6gARm4eGScWt
xu1w03ln97hDCGcCfdvaaTKam/Xd/K0849+0QtWosqlMt83T3PwmVAja0PO3
phazaq/e8fp2s4tOkz5olzran4ooL2tTOWXJEzjNvwHhwZoX92b6Wh02BShP
Hd8Fp5XNJ/6kmsHUi3O0a+9kHQRPUi8Pzo4cBbPz5SWEhqJOMLZja9nteZv9
pXh/P13sa6iM8eMx20vHW+EeEoc3ZOOeLWfrYTG8xFj0razl+nzffS4z9wot
YKB72d158CXwkA7gaegKzqa5ZZwpyus/JfSXhZEZfthXyvsIbERmGnSNpK8/
DQVID41BRwVXYh0swG6piYSLr2dBhTi0uG6i1KitDvTWkTGlbMNCnxACecGp
M70aQ7NsVNiLalIM4DPaJKl6QHhNTPvzTjo5xaTKsmhoGde03+nl3l2uieHj
XQW//HMKw/Nr42jwvOOw/7MZY858r5YfarYbaXZNN/dAm2kRftrGTx6osfN+
pNf03xB3mMHEFhlglPY64rhgf2Cy+f7eMQp9qaAeeDDqzrqR8wUrUrEzjjcd
V6Dav1ETU+KzKuFjZOHVT/L31wl5RYq4nBydHnJyG1g8OsAaPSqiVi1pGHjM
CXSS7d47+GjA6y9l9OGhqA8SABzl5lRF4tjcZpwNbR4nXJgxejJ6Ti3jCkqL
4sjda216e+K5z0xXkYzqS+f+G4X4HOfdoQBuzGgZ5ZDRplHWmBgeKGQExWv6
Cq6qXOEjzZORKphQVuMEvKtO1l1x3p81WIyBk5b1VqVCLcuw0mdLQM+TWzyK
0Kt3BdlqhFQsbU3ab5OQVjMH5HHFOuIEcUBoxPqXUDGP0uk+zvJhVj5SVX6D
DgsYSkwqxyLp0r7zJ5cnu5YcijWNMlWGZ1tV+MeAniX6eGRFxpOFH5haUCHP
ppFqP0wDJF3Y0pTH3GADMOC0Rt85MzMasZ0+x/QyiMmQNK8luONsSaWtgrW5
twi6AR+ng7Gnxi8XZUfTxfB8HLjAujL7gcweJpIXwtLkwXDv2QqSPiMH4fQY
l6Jl3BXxDBUFWk/7u6E5d6xkjz7LLmjlKMwcd5mOgSqHNTGbIuheP/h5ehwp
ktROZuD/7ecEqMuzhsLRJ6IHwiiFnNWlC9jUeDdfztcjaXxnG6aUYcDk7X3W
pBW0+BuSxXpHvZiKQlRZyy0vUTEtOctdWWTaSinhI5v4qr0LE16q9m9F1TT0
LOWWD+I11AJqaFOw6lzBi6Uv3g7xVrnSnCqNWxiVxCM0YjMuwjFR4B0TLVrg
3haYdPSzqmdWIkxtu/t06CN/9JeUo6r+YxKuPG4QpX3cnFNoG2mbAHhf7GCE
T5IAunjZTVFAqOuSEK61JEcxYO9v3c2LwCnEAlmVjzf51b9ABnnlnAXHppOk
x2Qm4PSlv6dqoY0lpFKKvRzuG5Pi/y2ikTbqLDQBHk8783lI/sCrnICFobVX
u2q4dUGeqjxvkl+b1ZBXeloz5sglbe6pEEfkZb4pfIsgxdl2Vgh0wDINUwZr
HIMCscA2vdeXVU9NnJ6LAtL/P0+zWZdRsqfa3kEZCaf7iix31/eZ5Iay4myn
pUP6EKqGfDgcSnnKnTV0Kk64M8HDmj0RDf14/GhpACfk+6XAkxGoqozPdbg2
7QAkNyptEPIBXedJ1nV/48yJTRJzabL7ikyZfu4ScZnEacIsgGboSeWu3dcM
EBoJqRBy5kUiIdriDFD/UIpcNf/oYD2eMS40Zh41zNoJDDsRHQtz4sg+zYdN
E5mauUXw4PxAQjDfdUSRJ8cadi8Yjc1E+eMkuMw7qzid00lTVs4JHC7RsJ2M
UeEpWLNp5X9/PiHq/M1rGIqXkQO5/OszRx8tgTMBLiycwb6A1+j9DswmGQr2
eUBjvhWU/iBZIUkpCAua8TgIntMY3bbGugi3gFSSCTGWO5dSQYwO3kDBGLMN
RRAqWxsvNZ5DFx4SwwX3+Xd0ko4iekNsfLrxvJw3sD6371ltdHOPgxeJr7nM
FqBTfRWv8RwPNN40Qyjm7eG1mcHse1t3rWC63xntYVH0WfoDVPwLk2jBpnlm
/f4u3L9SfWlSQQ4G1AU6/dDWSIwmCTLdPzeABy23WF4ZQ3LJyvtMhBMtfiIF
5yLRH28//6eoj6jkGATGlvEeThcftkK1IrXizO5iDi+tFJxOJ+pHOTYRMfig
d8pWZt6hRTchjFLOz9uXcFFtv6OC1IoHEroK2c7j+CJBWXJU2bzrkokYZYIE
N5oLYpApSGAUOOaEJMnSQamCpy9PkBM4/L1XHq7qcUFcQf/avDP5hKOIecCp
ZsIQJMY83/wnk3/1U6ovPQtdjaLQ4EgvnVwSvz7bqO7zi9UX5PQoqhflszNX
ruqi2MG2IzzpoUIxHhqCLSVS+so32VRnSLqD/OHNm3Ytp4hBppHTzT6clGv+
f278TZc/FMVd+pY9+dje+9/JCIxd/82fBT8iqVX+QZBEyCA0kXr7emL4XG28
owVp8sg+He0InJ34Mh8Ln8uhgDuBvyu0qen41Eo8GeZA/xKnOVd5RQTV6Wox
Dcq8YH9sriliIX7/NWMSKGVoQNnd+UWhBs/z9ZJ6tjg1MaiKnF55kCf3fdvS
1/mkOAoOOMwqSwpZLcW37K0JpQGCuj7Kni/XDZJBcE/Eg6SGeNkGj55tXzPn
T3StGdByUsmVpqwD0qBJwC4NL2Bpy9BfxGNSi0quBY5KzmoEStJVGd4uYHOw
AyQyINTUhZe/qjhTXrdD82nMVYA10HQJQ1uoReZYfl7MZawQwMUhWtKKuUOX
MEKIt3q0gE1TADB2/uFs6BehMzKrgo6QHleEXODz23pgUxTW4wHWcISRgFK4
xP156HMxAcJ4EaFP8L1NYoG9xGMrfAW688zFNfvhzP5W30sXzZrmC7A28u/m
Ly8OByFNs2PMySnZub/VLqryCkdolYGwljkeuX5vZzmP2hPegRdBCu8VsChz
yw02zvme5CbdIVPL5gwACgQQWtmYRdAFIrHPeGtLjvs0j1wHewYvU9u0XxCD
GbPgz7CIpRzMTIeLDM8EMYLxz3JjYXUsLqw22NU7Vdu566ioPi+Xbpnck8Qe
Fdnno5yhDFQC+uNhN7x8MsUvY3BtiDKUsNLbwPnpOQRoBSIk+1h/s/1lxC+j
2QTrSmIgW9RQIN3FflIXRMTDJbzPX4a4ansk89Z3WlSDRY6IITTO+2KBByy4
AAA/yXwj8Ol81zM0Cx6CHeaZjnqDEMytZxl6To+xcWojCrKrzSCfWb4VWisj
RRIPSOC5/ZIrGrWgMsQXU/uYtLJnIRHsvCKp3E7+2nWCjmYXPyj5hUejYayC
tFQwk0Ni7uIVFuFA1DOQzcIgBdvQIOFcmDsgnu/vwLMsg+8GpVmYRWPGnHst
W4cEjvBsDwgKAsyAYjEXQZrmaVXokD1mYebBRMq+r6/QRegGSY/xXcin6HZS
3Rwb9UwHhP1a0NsxEy7hKO8/VaFkfsJcdnRUbHFcFWTzV12Fq1QJZKIet5Zj
6Un4jfR4sFngbvdALXNoHH/N+q5l8+255zpxnYEI3cr+EsBPQutLoC1mpe/D
V6ChCvEFHf2x5dtCQofc53F/ubO6ww4BeHLGVn9gt2TOduWh9/nHcJy5iAl8
fVQLigY7/MtoXoe1siPNFF9VJhJW1WTh4Tc+/Qnzn5miwN1lDfUm5Y3OjJIK
GvyJv6MFi+wq2J5eOQxwm0wemjwf143gcnjyGM7eKYZcFmQijof8Ib0pn287
PszAQn0wLRPCFDYch0fPDgJEFwZnN94sx4AtZTxv0crpqhD+jVBFaZJJ+MZ7
5XXuCbxSjHjyOWh2FbAfV6pqu6pXdZHXT1dGBD2+KPu8tcnO+41g63KArjXM
d5GsNYvcqT+4F5qJyG09RMLu7srYNxHed/U2Bq98oKxn+ddRlU1ql9kA+ShB
PoPYedo/KOCY1Emr3lTP2FdQBxWcmlvwmsiZ9kHtPe6cbNp6AZPyoI/dIFhq
nsCsV+rL9zffbYqhoqV5e6Koj9UDpwgmnXxU6o0ZR7BgZ3Ps5U6GyFv3OS6/
ZWR8QBheT4JKW6j4xCs4sdfqMLKkJmgnyjoPPTQA6JVyYCdW1mPU2b5esDhA
X4kvet3MkKv9+82UHysy/N/kWRWmkj4Br4itqCx69xPOr4WpiQZsa74/B+o2
OTZIuzar8VfXKHQURI0J16SRO2VLopNpRVS3D3c4gy18aMyBaTzI2ypDKAsc
AxpMr/fKKaEAJBHrSeF+vC1lSP8oLbC2XXCF47aTLiBRTO/D2HB9w0U5ir5n
uaiYFj2A5wPhbLYczn7r9wxMvyzmAweYs36lEk7NrG/8pwN79n8A/IZ6vXil
n66d8sQDgZK8ClmHlsJQHY4Wo3T+ZzCmZTutJ+Myc308ZuI49adm5iESyarP
GS2a5o6D5YkBL46eO2RyIVyo2MRsWrXBKda6+xuZJ2ihUAYVNbTkPVqibvZt
A4ZUDblCrLoUthfENzg4dQlfv43BcgKEgUVuYFRfAsINEZGohaPXPmYOEE38
smoOSqV2Qnc/2Bv2IWjusaeFxhAG2yn2gABry46hxe+tAzoaaLjM6ofuIhC8
vqv77zHX73DzGxUrGSh5DY64pITpd4mxt+Std5NWMdDpHnb3VMyuxm9tWr2B
3lgvcDfhtpTdu+h3/29vva/LFRjD/QHQR0gMevgrCSzrYikkuIAqCRw/T0/5
7TlohkEipZ7zdpEwbvfogJni+3GmEtVLT8apasqdy0Jr9s3FAbg53WICacFe
Yq/9shAe77WAjo9z1pVsDQJRcfMAS7eTSFkjdjvymUzoyqb77em7sYvWT1g6
fWjA49oEz4XQ2oE4n81tfhY6L0z4YjCr/rFZOiA9l4haNQngj2n8x0RAe7bX
csRmfOkFOMnQj1dyH4w1dEpXd5ilT91Hf/SY9dTMhfTHDMQTkQJIVaYEYa86
gpI9oWxkD8ZYaJOBqNe0CM4hGKWbgl9NSICz+aixgzCMIgcSTLwxvDj/EJo2
CcnAXNldJSvvV7NwqCQ2A5EswmAACeKED8nMYgz+bZUrfFmjzmg203PCymP5
32L32LfkTBcPw4fhAZHIoF5KFuBpMsizvlFJKYXEtsbBOMboWyZVAfZ+sAaV
F0V1q/ol0cJbh4gRD1eEFTio3+AvyYUcrY33pqmVeuEekVZujLm/1LE5Jg+n
5LTz7MjwrzJuelQFiPG/Ng5ntvrAAEyUII8bbNaPHneJ1F2Wwi+3u/rSSEFs
lg27x/CVgAarFOT6bWzzZMdlFKF90sqXxVsCTc1OSETR0yKjoZECAGDOBoNX
7hAb+25L2DO7kJnY6fv/fCNlvzvUGPXYCOqDiHtJscRjPQU2uGetCgnxJIax
srDVdvw5QSy7KrY8BVKW6uXpgOGREpleJKHosTupr6W5xxMgfyuFDUxuk31z
fijRoy33EPW+O0me7qWcvmv06Yqmcaqej8SbwFAxfCMIG3QGJuRxyeq1gBKW
SeyI5mx4YGcSqPzXO1R28HJfVHNlnEJFPjnwF6qFxrvs+7T5fJze7uxJG9n+
xej968DYvxsIoM5M6yAGyq/62TLDaVzoVpb/C9Gb5EcrCZ1kaau6nklkvr9x
I3Wq2nWgo6TH4V3rDo1qdaYU2odbeZEMkUEodYDrYEy/yMcHzU7rM7R1paVk
W6lj+phOZlLOTrFtfjGSIIunYjvwH4q9UeQHQ77KpgzpDXjFLBzcS9simlWH
8ezatyW62xndgYfjDJBrxaXTG9HDRhUsi3L4JkaKVnGYcgVV68uO/++i9ZdN
59oCrCAHECx5OAqra1GCK/WAIQJjdh+Rhm4ZtWBF1nK8Mo9CMFZXQHzxNRL6
xrszXtGvkycyp5m/nyoDi/SNhsq+LzzjkZTHlb50eXRJ0Be8wealH/3K6sF/
9KPnp6nfpn1lK1hZRequFIyFYwATK4yRZwiqO+otC4x6+AHArjAaJ48uiBcM
WHP6fkd9HOYXY1I7RLJ3TfZP/NxAFV6DlgwR09IWraR/0aziwPHXy++1ggEv
zzw633qeyC1ChH7z4MTCbiXTwVCYm7a7KnbhozIFEFmZ6GLO7Una530mcDSn
PQwlPq5AqkGDYkRVFTUGGf27wR3EUo6pyAhKV+0tcLhOfPMpdljZzgrI76uA
k+TgN26EluNp9cu2mdggWihwQld2aHTMZwGHqnU0cM2Uxersuw8KghpYDNZq
uc84gbN5vmWF2sjMXXsh3jXlFtBMvc0bPZby2d5B9Npj8z+2k8/uYAEjNrRr
R6NR8ZM5qy/ewCgTFrDiuFzMln49aeIr1Nqu6W5OEmizai9NqrnyFkyoGVdl
+fqBfu6GbSfDuJh+p1lk+9AAnxomY4s35GQCnCZ8nleAMO4IFg/dQy0JMIYl
9dtCnXMyCcAMTWtd5NcYmvk6qKcDbSUXxm2OTE+XESe1KNVNXfwr+CVBPZFW
KQRPpnPja1ivgYrER/4MS0yf+FproOdyh4+3mPmrXaYqOdD4SJXQ/G0pcli8
J1CtgrEWFw4ApCDP9XUpJtNG4qm/kI/Myu2Vwg4izunGwoNMbejMPca7SD8g
U48c4jixhfzAmnPR0TbcB691/1lDCyBJJAHlDd+sbNeNLCvLSLwvOfKZNLgN
QsyoQJ603gTarjK28jmNJg18EEBCZoq9cWUg8DcEPwZjBxJW9n/c+N4DI3rC
RsRnOkC3Dij4SfcE2rX5Ojy6TfRyqkUyD6+0CAzqLPnjOiCcPZur36t45i7X
j+J2cd13rFpKto8qV9HKXqGd2bs/NtwF2D6Lq/UU9BklMZV/Oao3TEcTJ9P+
cN3fQFUfMbIQ/aKWeUHSjP5ESKmEe+SpPVDeP0o2bQS1OOw2pOmyrThAiACA
j+K9FuvHLNgpKuyEA2dT1OYxIzWUPfcM7VjB9OSk+PhIrKIgzgzwZqaAB5Ez
oxzvgArW9mmwTxrkqKj2wZ1jmIZkxyzutgnPRuUiVoZoIpf5HE3WC9rsaZI/
gbUGWhJeoVSobosXa7BZ7lrYu1WQw+pQVJIJku/+Al7q1XWEmX1ovAC11n6W
PH25iazIobYRbZTH/XdpgZ3/MKA7L1zarm4RGROVzrOByce+lETKjz7bL0iE
IUIKabNuj+WRQvNQEkK7UNPbJKGhjOyEu2Scs7/1qk2noq+B1PnD6c7qjEYu
Z7khZUBBHl6qStCaxo+AZi96hOuciLARCygU+mH6VjLx/fDgIND5HMPon5Dv
Tpl6den3//q8wU2HksVaIiCn9Iji5ELX9StKmvdzh78L6wtL19Wb751p0Dm1
w2x6HtZZWGbAodvbh8g51QR3+Opky/u1tfufwihfJgoqYxyMsTKPpP1d6/xS
Cjsd7NELxeUsUmRc7B0k+xRWo90zzLWqZ2noT/MSgYQKX5QB8ckNqCD5b0+6
c+dyucv/OQS5+QpAWtfbUQQ6Ys47LB3MdA5LXHIOWKZwc4L3z9jEwLxlZlQC
nx5bmj0ilVKKCJaSTAdWs1z7ApVmbePD2+/1f8zQeywskWzHI8tk4/ze5kBH
b5JrgPKL3G2RAZAlisi+HuWzzr6XkrDsXfdjZlQ8KF7waiqR1hcphlOb+JzJ
0W9IyfAe37EQVBofHJH4i1e0JTza4VklfsjnlHkmBlHTptIJeECwehoegzHk
eoO/7Wo+vAGXUEICVqwHv/0By0zcicWFobq8yUngZEGAU1GGDVb4Vv2KMtRH
1/ER579ykFzORUAR3m/+6Ym6z4+w/TBVoXp1aeUt9Xw/bdT6qZ6s2/azXxQF
E677oJyXHUOtd6AfSEGnG/KRyR8KKUV5Km4sLU7dbLFTbjWeZU7fB0wG5D9C
iYEhSRI3/tRpSROmvsW/hpuIwpI5ETYyohFXkhwXZpYK8cUCPyzcn/sInLSK
W88rKlLfTVc8cvjw7ZUKH0H5jibEfcqCquddCH7Y1Y7UpVW9tzhfthoUIwGN
NsHR8a8S3EuOMj+3qjsawYyXJcGDyoNsUVXUyJQqVJdPn8W/osW1F0jLq1yZ
RPH3BLAlvIm305rVeDsOBpH2EcS3DbZkzl6XMJ+/77fkrmLyExfvRHYYTDcH
lbZy/JiQYmySKKieyiW/2uNd78QTA5L735CAAthQEhd9vjlmmqbu+FIgZ5CZ
unB0TrS9GgRbL2fYtMlJUSbqEX5B1+RYlSriAiyUHPnCPO7oFE6oSDAHaCJ0
H6Rz+HimZ1jGIIouYYcUBmtSo2870vesfYfkF/nXJAHgGyCXAnICySNiC60B
vED9vY6XDU05cNW3Ivy8cXPkRWzfWYge3fyupzj/VJayuXQYJjd26PnUdy5x
ciPPvimdxsuAb674qfZBV7XEBNdrwvA3kZV9OQz3+Klk7BTEAv12nEDZAYJm
LLFptJOEssc3UH0gGTQKirB93QB7aKlsh42k/Ky8pKpAuL64QH7TjefGY7aK
CnAnJpiaZLcKWs43NqJLfInvmlOW32OnNi2gFOhFHWO2lArqGPRUlQqSNG71
5hZ7erSR/wNasLJtwWiButi/x1CpbibM60fEUlT/1dNzVmDszDnaRBuFI8zr
fGka17O9WQLXBWNhVE80DY7RmiYyeg60eNMY+I0OKguvqCio0R4kInAwOTau
bvB+5DtiwuSNJUkYAJVAWaKuCmk6rq3bH/Ewlmk29IZUxGt5V5OBFAX8M4tG
vy/tXbaW5FsncmeQ8LXmq0gejPVWx4gF9b/RaJhQqokPXe6XKE9uOH+yFNbc
+ABaCgmboHjWj8YSzsnZNPEsCoiwFYkgTSW4cOAgg3DIXGLI2MvlWgOwzL9t
0Mt0nieT26vS4VfTThjwiJ0gDH7l0jnzvQIqb9w5vJnZN9GLOG6eM0Ppyf5Y
cYY3uA1mO0DVeko8mx7uGqmMLxQLrQzSu7jKjs5b0DzOK4zEtLMxM61DXRv+
WUN+lx585jKWaLbz2Dt+u74PnfFjylYHtWMMVRPfQ50FT6FNJfKJwO1JESRd
8CrJTowcg0VDbc4WJFJfMa/7Cw/v7OSAcHFBKf5iDEhg5TJcArzLiXIr3jDv
55PPdlwar9ijjvEzB+N8iIPjpzKFksu/H1tBgnRUFtmfSjs+Q+5UNqhVdWzc
WIyQ638UEgRQd9l3a+BtKFXMUshP+3ubK0PsNJIGTYFF26J4FY4wksm4Kpn+
AFhQJD8JznYlLbq6npRsFz8Rc3zJcQxoiLgFvyF7UQafKJLN+/3AXuzWehoL
l5XvvbwzhdxDBhCAVS+Ej/K4i/+pp9Mu8FvwvovdeOtfumgzVp0QmNBFKoEr
77qecZHN2ZXxJqEVihHYZldlKv0SoBebiXGp6Qj+ZTJz1xSBWMBX8A8Rp5rs
9x9OFeSjyksLioU3MG/UhJ5W06GPbWlzT000pjezQiopvyAx2bM+lOPd968F
arp98bTSaJEJe6ZgYV4ZMEaDJg7yUVtprcn/KwGl6+d1giHoX7en7dQwv66P
TdCUh17lrWT++ZJkPtxomFyQacQ7N2Gxm/mwjndPvytnrSSGQIb48nHAxYaC
Jc4y2UpBSOej3347Bug6Y1ZJKPZplDJ1OQPN3JFNJrBN/ZO/8jEyD8A8MJd9
boTgWl3/Hb4r4itg7VvJrfFKffp6/mZDS+7xogc6RCDRo3ISBv+Qg7gzLMEU
yAQfMro0VbuFwCC1XtbEH7y3pluiBUR3rQn6FDczoRkKKiiEhrdeoRJvNTb3
eu0X3tQtpK6apyE1OISIF7ZUh7aNTqvUsjHKM7Bt/dRN4WB5OppajuhXVGIh
8To5hWo2+qBXE3xIMirOa5PfpcGyB0nwtonOFjX03ZldNSLHExvON8M3Qugq
3nCN8ZpOTPlI7ppaI3GF8FCHuLGqJSMoo774KP8xiNPv3VSjAoEc49XYZBvM
MD9yhi3e0XFN86Qpy7ACsBMZq0aSl64Mh9noVjDZDavsH1unAA841cSzO8rJ
Yrbf69b6WNStFwnw2anRhIlIGLx5K5L0wap9hv56BTWTD3fDZdknwY7cAxld
1bYPuiIEWw5EKbb4QQjePwGOnbearTOghxOLZw2Pv1Oo3+m9PXzDyVyjQsYf
YrAhbZ1rVfWyXp3IMP2QAFWDZ+cW1Em6ZKhddYPZhB6dN1zEFvPUQfN59J+j
qzIQL27OQ7/22oZyijh/vzu89IlKqc/yxVCy/oNPJWq6u5VsAJVYP0MEBzRE
xemGTcjjNVqzextvSeEVyYGaTIkvTswLypfgCjqzsoRObqcDElaIF9J1Q41f
7/0Z10JjpbaoN0dYRCuM855yjeZmwuB72DHQf4ps9KzlT+yd010YaVTQO6ev
QF2tOWSNbrBF5stKtuR65w2bhKFaSd69nuwd7xw7tgb4PBSE3xl1kT0ihSHm
bN6yPI4ul83AjfRa6i0J0iTB8OAUksYgxftOkM/4cx6hnwcSyQ4d6MrvT5lZ
0BLsqKgk4K1rsbnHC1YAnVs+RfybR0cLgD4xOs4QqZSvu+8manmhAnVjlctL
92yK0SFvznzMLUY4VYJvnkW9t636cjx9MnST4JcX4jkYO7Uo6z5zJLunAoPM
uw1aMvv8yuiMVlzln8Oh4Msy3nqDwdGH/tNk2l1sgVfVWgsi2tPsQoj7F9J0
MaUMi/kNgnvvVm0xd9C4QQ4T4Kj0kLG0C5jDujhKgv+i5WB5Kc7p8GbMpKun
nvZpUYmg7Z8jl+kjeXFxRpRDZ0clWKsnX2DoInin1KhASIETKgmPBqD9kyJQ
K/HSXOTBP3NWu0mKY5FYMoIE7aIUiJK6pqd8Oa6YfjBDYv59nVSLU9vRVTYK
HNPF+2UYRmtp5qic6fh5UsHgqzTY6asuHZkivUA3U85+0GbIhLWClHWRR+s2
xama0YgkVATE1lYRqCaqpx2jzFW4x6p1Ukr3pkcZsUlY197olErNfwgJqHjW
goPG6QJHd0UA5XNDFOFxFCaykG/U2p12gJwhfWe8sEwUF+gtkZV/evSpIUua
WeaLAOy29DC6mbfNkYwmtU0mVJf/3RgBdHSDkQcma3H/5mS9YFTc+PqQjCkZ
LicXqasmDLn3fCqjpM/NTos8MqPHVv5iQMvTYnip5i2CnXaH9wGr3+tinhPa
HX92KvcGvCPUNgq49mJjtRC9Chc3auofiOIXOla+z56y85ghg7qCTvCZmntF
R+3uzVM1DOPtE0soGmQU6bgqXz/L73oD6eZp6rewDmMZFrfUg1EDumJHpqCn
FoHoy1TnGKUh4llt60wDdXA6SQ5Cg6tj67Hztt+lxR3x72wIrLTVEakcYpKC
/D2XTIyp/uNYRfW2eGLs+BxlpqQygLCeqZU37065+Ycmffl8wsxANfihUdJJ
o66N8RtUdTV3WrqVJQasgK8I3DwFMqLcQOv2EFA+owwsPuXUQkGMa2fUz8/B
OR2piwPg4j58pmjjExuMOOno9dCkTyl9n0FL7LqgcFbggoD5gTetEZInEoIz
eKDCjZ/DDi/g8qnmxHBS5Tz0K+65+FS9uBPW1oPyFGS2qhp54ivQavpVepVj
96eHResxaeIM6e3wgv14XOBjuwsp4Oya1ncTTsCc0ETEAhpQ3m/s4405c5zE
siNqeQidLuzMYY18M9akSJ7UdclbIrGoXyHFIhT1Ab9y/IL+YZ83gByKhPHC
+gTm9HB6rOOTXtOVOGzYDffPtn9i2AkZTeye97pSf8tr0jmIWYJqPYT4A1Jb
6Lhb6Zr7Pfk9fEWIw2W+eA6TrIkKKiO7BeB84nGDo1V+CxznnEOnXEhMTkAe
5bFgVnjXQW4FoTGyH6dsbnOJAfRHQwO4WO7lH+MRvRC/ApmnTV3VGFf7VEaS
B8B0ve/rZ+jWVKjwvOStt6jufGRBRJqxIar7OZBQdSMP+Ox7cfv+EmJ1nwvV
H/5VssT6q4S/U939+xjOsvoo4UjeAACOEGKflWf8k5LAjUI46bY3qIBwUxoq
rnAZBOVIrF+Xp89sTl9R5syvaep3pa9B3ErkTgD0F5tI+TSDO1iWPceZwiy7
2pWkyWrYxnxGMewZeuvsnwqnJYIqCJatPzUySBZOty9lHA+RTGb0bG2D30CZ
FAjwvUP+kxXodeO18PsyVHlEvTj4hIky6+Q54VvWlDvNGjuTFPpGb0XhGCzH
cJOTg0LXliJJOcQJEMJNOXvi+YlcoXMgXcg/NQk9sFulG5/uyLQPFh4IO8HM
c2EFfU2TziwYge81xspzyMIfD064szhQlrgKayT2bb76ViMX2WmTwMHHrdPb
RO2h5SgZE6yv4A/R/AJjOqY50czivfGa9agz1A7xVaSX2RLSbOhH0aHEEqaX
22Gp/rwVaRU13O8FMgpZOLTY80ttoEOenXgR4E2+aNrAC+RdodcWA6OGxtbr
BlBT5sDoZmxYVXyKrpgo/i5qCHY1kCTYXkPfh9m9S4kJQ6s2X1ssVZlPBCvy
C8zbbAc0FFV1G8/fTk8Cnf6LCo/6/5PCvluUb/y0wPq08FqxHWztlPF0gWSv
FowVyHo8/lw/bmq2s5nUSlvxYnELQkhNYw+K8wwqDbvp8UH5HLdkEW1RcmJf
pTpyfHFS8ZdfivQwjPlaOBP/scQXUz7rivAfNyZvqthMAeJbsHZxlDwCoxfI
zLQPXOwq6wtd3Ay63VjnrXlo4/8ewcYzYUXfVvEjcYG6hQ0TUjWS2AvdB0H4
CweSiUk4ZQagf9lJrcetyif3HhQQ6oxi+CHRF7T1SfFxTUQV54aOz9Pqna7F
WrxV3iRqA+m2sUdCyzrry8SHpk0XzGXl/eH+PjFRYFJ4+wepGVWPPDavug79
wLoTDYWUXAOzTdsIvFa5QmnjoDMPVXqImqIkn2cAs2XT2v8AfLtuwodAkrl+
KzjWJoza4OFjEaVrHheXrAq4N+tUWWd1J5nUvaGe5D2aTbFV4bXCWTU/SsKq
2Bs/9qGE5qjEXPPp/IPmmduHe3+Lp4MGgNa3EsY0XMXFO71ecMvraay2wWcl
IdlK/mmh6LmWEiAXrp5iFNvzGL/YU2rLF/m3SoMm4sK+u2NudExucMd7/K3M
bU6hchDi9QHFjRgCB3rcKm3v2MluhTlYr7XKv2N83143bhlCSw5GAnMUgUvi
4UmWbz+3Zf5RcGY+mFdPJzI1dSfPiBv0jzeo55/aNkqPs7ilJXRvV8he1eSk
cfvK70LgYUlEG1i0a933IojzyRqssfNXhW4S1OhdcDTS7rKOJo/Ad6+5Dz7U
VNCSIgA9ZZQInIGP0AWmko1g8OtV4XqypitJ07Dj1MBduCluz8sf00favdmS
SGvB6f3u6Li6VvfNSvKYVNFd8nu9VYiyN2bi/J90s27JXRATrjb6ZSt0ieR1
U0F4rPNOYG5MAkKbzDaDx5K2VjeKk/YV6OngCD0fug54xmISqeuzQfP5A0GU
xzCK0t/tVX2YFwnzQfbDI5mx+yxtNVsL5P6biPePCYy78IUvSRC7Zrt+Jilj
Y90PUEDakRhacQoFX2ZT7oGPW3xJ1xsvWXxz3TEIg6JIw/rgkry+rZRd1LNO
oWWpLiIdLTDPBQ1WO5ZlEvN7cnmeX/743/OMWgmmJPaiq2IoFKYS6g2KtNYW
wjDEsJUpmfAUhTTIav01MTiS+A6he17hMyZEcMyg6NYfMtcIcELxhdT+LqkC
JWSamenfM/CmQaYWTJBhBixpjvjBp6p1H/qe3wS8zOLsGaZSVd1EJ9yep/Gm
62ZtVKgS0WnovIRqkoqP8RpBVdmySaLLG/Eus7SbFXZJTr2rXrYmFGcNfgza
ZsR2kymdszd3xtvWKtoWDAUqbthS19F3K5gn/YbV7GikwBcUGPrWjCi5DTHF
mZmTE7qF/aivZtaCE40Rx76TVnSyvLONmgxD9eR2GKN1fAYrqa1PD1x9z+DM
8XCWZJPWJdoPutkPFrc0AB5MDUacLFrufw1MaeVxm8nnr8zkWf/7Yf/g01nP
JX6X+mxYYSvzQ7a5l9qh0C0i2iakCgJMhUoExaV+BBtk53qUtwgGC8PCyfxO
b9CIt04oYc8RElXY8v4rqCWARW0x4zTO7Bw0NEbhhycXXgf2CeaQneR2CHyT
z8ccqOWhORUIfljuM8vZ/OdA+6F7Nz2jFM6+vcAVLjJwfiAJfGv7kQH2Zwai
kGs28NQxvM3UPv9mSzqLI6rIRMCf5JVuYo4Ty8W1G3b4ME4hqSl/0/QOdGxi
dDzd1nblXVkUgUEoKe2grRRMJRFyVugrf1CgXAlh2D5262zvuxoMfshwEmry
N2aFwmLYDxlO069XOhrdi9nBPVN189jPTtaSvKPmX5iCp1vaROhTnQ01s9Hn
AQQ0YlRRCYGcCa+fYzv2alvR+SkHbAoKXygG/SUuwQOFb6aiZoHRTHtzBuGV
MteOAj9k5hsD13Ky+jahITIbXcsuvJz4iB5qG3Dvl9UjxtTlilTNFY8GEcza
+nwOuN05IKgSkip1IPbFfGkWp+dsBSyrXyS8kK2kblMm42g+hTIPGg0GSjjc
00GkisYC8LipNF8tRc7SEEWLi8Aat5D6rK4Ic5H7tYAbChKxEXZWAm0RydNd
jxdTgCRzFQhi3RRbQQWIjFveKHWMcV7dJcYb2/2LwvJE2ul3HQxHN4fC/LK8
Icj+ZhS52XaOtatSRxqqSUjTSf/kK5DYRPpyN5sS3pMLwZJx0nPNAHkFw69G
BsmYQgzAus6aH+TLsiMDFSHXvMpHEggwi1EdW5zqt5cwj9TMIoFDJWtHXrJi
gZ4/c4auQ2XVe6DP8Iw3/2gL2GwEJCLiA13yvcHtvVwY0j2/KThRXXIjQJp+
QJMUS6iguCCfNRnwfPki70h21ovxpx1nrGBbf5tREqC6hnZF67VQwGEPsPLk
hIngiGumdQ3M3SlD660GI78FBY6HXg2vjpSv+axgCBHGmDcnmGpvDD8Pnh4U
lCzVYAiuaH+GR3P79K/WRbAwToHj34tcx6F9DSVhjm1/TnGC5rvRProP6ppE
AS6/jgNKTwj4yZjpyz0DobHmHuPZodsGegCcG/8+zpQwUgBPOHAy1Oy4I3dr
O/YW8Bi6RWHsB7TNtO4FpdpWJt22zUNTPujI4VbB/Mx+WXtOtS3Fr0j06Owq
2/kSmNHuMNT0UnljmoteuhIpsaLyjQfBIWQ3R/yKrC5prIPTsEw+rQrdZKo6
PT3PkpRnGarF+pv4d//5LUU8Ebb6xp2lfXd8dd0sBtuCEnSKraFSAamQe8Nf
BR+F5/P5Ak+4kbfhRBM2zE5GITK/dvCyxY8e7T+Zhb1wSyioL6sQx3Z+wCyO
awDF/nOEJhxdhPHr8+kA5jpuiUIwQVP2fmlpM5AeHqIC5ZSJNB7Th7SP77si
j8twyCVrWO4Rlrez8ERtfzWv9zQigLLSv6ehaAxYnFMtC0KbbfkP5Ujrvzsz
sniEZTjSxX65kDPlVfJEEaUaEVRYs4PB1MJqntrsycfd8n9/mlycM+CeaRyp
INwZOWPnXZxZuufUsZJSkui69dW2Ff9JlcYHQg9Yx9VdRtzum+uHOyP/SWSz
HDI+om+icuUdkVSSeK54eEvQsTHGmwNUgFFlTJysP9ux99Y47h1qHQBgpudx
QZ1IkfC/jzsam2pHLitFsK4fbp6qlZ21FRE818zth/qCUTSdu2sWrzButn8W
bH3IQg5FQ4/DAghpBixfaYu+qStj8yFvpNxVTy65V7sl6c/PbUHOPIQ6/t/P
Su8uY1F4axuvmSukBtJmqFb9SmG9Bs4eFg+tFReAbRoLiVlCF5UnajchRVvx
+As5KBJxxcRvSgCWWeS6Zvz4xlOaYLNTHSpqdE+SPhixICRvWsgMsEB78pgC
VLZSwJhoRKAA+ui/Vy41ae0ZE9m4pUmfYvATOY4d1jVlBzR/oXz3Z9V4SOhT
jgapBl3EKkYD/WyyfzoYtNqgDMki6cEwYO/N55rugcBmst0WSBdMuPBIlUbU
9ObA7WzoPqshhvH8zEeqtO9CIEwtyCBaZQ0UXv/u9vvyq84Su0PSW94UwGaJ
/ft8pgbPMf1I8jC69ya1OvGGJCUnandU0Zyt4udaFFWYA8YmolD24xKECsBU
UZJ2anqAr6KMl7HJJ6In70IHErENxe088Z1DaZ5f2bKpns+2bl5XNiMNhgHC
dqRRh3jwcSpiudkOrbqQNA8a+xSFB42dcpSSTy7g9EGPUC7HfAQHiSChQF9o
PJta6Ea/eXRJmj4mNXUIXUXQ7K5FtnltZWZq/0bLkRWWQdTv5TduzmGsODai
eInMKrYVAzpZF1adrDs2TGIdMOQrjetIxAZPhCWr/fizZIdkVMGwWqDwL8ha
5wBAR/dx38dHzNPwm1574xkdNb5z/7z5heaD60c1bZXA1NmBn+kusBRAOiHt
v6GSXZeddwp4YFMXf3KPVVdmNhM9zqTE9w8jJNTzq9Ax8cbXYdItB9SlbWot
UCajljcO7R9pcXuETO3vlKA7rTLOeDYm7CoZu9WoiE5FRwpwJXvwBIGXYAfl
t1St8oiGN1mDh1ic00r1cAZE0NeuPMLnDVe7RRRphbO/qV0rm1aYBEQje50B
AP6MFI09babir1TgNemiqcMi27EkkeTX4Wb38v0nrB2zctoQYK86EW0TLhXJ
JD6L8+MK2AQCuTZcBvFEHsXHWItgYoxg0GKUQ9OiStyJOBgt/+lIbWuCVAiE
DN5inpyIVrzVd3LZXzWyhax+kRrQjnhngeoDXo/63XjLbKQqVmdD+hJjRHyf
3l7vOf8iwxzbcxrpNRaYyC8hguTRM4qeTuGaUOr8erpgsBdeajdrHSYsVTgL
oILFIA0qfRJ1HU8vteJtuS5lsRDDkREIHp90D0lzKnEzsJmSpXOwU4TMCU59
4MESCnKpMZXyHRR/pRdwtEEehXPKjMCbcvbYaKzMmTGo5BGAAdPvzmMEzIQR
sx8EzSCxC4aITCTbmk4hNNhh2piCqjZYKQv8v0hmNCU3WcoxbroycrAnL9/g
ZRmNc86C6ffUDWLYfzk15zGA5J+LzoyB/mZ5H+l+KO0qXNl/oTbOLwmirDuX
XYhi1sEu1fexyjVItVd9MFiZut3SGJZ40Fx6sHhhqwvcRv1fh5asdTA1tNsn
MIrsVOkUmaNwUup+HoZ57+sJCnjjsPq2wqiLNtR6g2JPpRSoVqZjVuhgVXG2
wSL3JNBkW3f/uuCVV3JGfYeQsltod2FxdP4gUdSy6X5CRX1vmUWOiEP2wVLS
EGQWaLwwn/DYK3CbmxPrQnEVkBES2+vdLKQlC9bfJ2eYary9txhWwTM7RKTd
fGp47/PorHHCA4B4VOesDZgYNmhmglPKZFkG/j1F7j+nuDmnkjOiOO9Rgspn
RTze6sb04JmmSPR/hjbYirSW0obJy+WQPJLx9wUrSQr1Ntf/OCx6XogWe9vV
SG8IzjyiTtFh0nclBrUkVPkYS21IXN2irE5t95bA5DJl9I6oNRptvSnk00tv
CztX6VZTUzvPzTYHD3iDbs8W2EUk1bXmJiJqTqrkLEEqE1TX5t+HaesddZeV
tWoPCpMfKX7AXYYtLC39dTH21DosRgbeJpPbziXA/iQLanlf0iSfMou0YzML
jL0BVoH5W5qvRA7J4FnQJzFpve5+xfwCWOmGU3u6Cr+totWPRmviHkrHFozB
bvFFfhEpG8x0jr522LWUttBC3lf2uSYcC7DN+abMniuMHBoHBZdADh0ZG1aY
rZKKV9dy+k4SBq484/f99qgCYfLTnn7eLLK0vS9rIwI1icOJdC6zOB9NVX/9
4bFD9OFP/6GHHfSshN0IBA4ivCwz6wmGnu78oeiImj9z7twmYieExTHa02lc
zWNypbnL62rmXWPxGyQxklwmVUPBV8hUFjQKr7VVfdaWK6q4VL71x2vermeA
YM6ZzXWWnZFt9gOcki3E82GldIbO3NAKGA2MuUOqt20SpjQnt0NtFsX94Uns
w1AugR9I5Zdn0tvKdxipbreOgT53pzFVpFJI6OFGECNcCdJHzLNgYIx341Nv
q8G7kSUzGaVW0pBLTMzmBAGpkDNNc4qJCgWewIW3GV0aec2BqXL8Gr/1o5K4
3jLfwvpfNGFI88AAWFwp4vQUJKG2tZ0sBAvvItjB0QeLh/NMX7/pzeeYrlkn
DcM3KvctIwDyVUj3Kwam+mwkzPWADuEGCA7SKVOgCnnPCMUK5mqfUGaqn0ME
OAV2u9iHJ/f2hS57XSaI+iQyJQnwtP5AWO47cdF3XplmWEZnzCcUrN5E5Y6J
NZx54eQqgh1xORZA7/ar+q6iVVAdkLkyDaRBrm2p/2dqUSNqHVdHyGPWSnYn
ds/67CeYPbjeNUktt2K7Y6teJbHBMzS2xOK+a+o3UuQZX9vPgG7JpczVuooP
LFclXQNgYhURL4K6c3ITZ53yt12LSqvHAPLkmsw7F6NZ25NrIoP8kTUFTSZG
xbjhGr+yfbxOTIv1PumiirXotIvklVWHBqi+bMWT8MjHKunuUfBo3tHOrVvX
tnx6hC5ex1THYpheoOGG2CJLmeNIx6iQjXW6V1oHh9fP2+AAzG/yOXUl/+26
NMLXNycCA9jJp97KNaWGMoaXbqpa7mIztiRePxo0URtLtNphulq+grppQkt0
OcdkBZ4coDhVy1bfUzK9PCL1VKocCoHLdKuLxqLwqlxGGLYx+AM2q4y6r/z6
/7CnuE/JyIAHAPSesRlF5eE49O00cr0AZNSeHUzfjScSRF8VkX7E1FmpalT9
Q0uMpHqWxhvAfZ95hMB1Q5nldh8hlXolKJhX9SQ9Hdwj14uGunP4/Gigz7jq
ou9nE7Bit+7FjOxm2HTm9E/GAmW0dpSMSVtGch4rLndzKe50sCBb95hLn98y
pne3WjmIU1Ah3yiZcH+83AvqQphW32McmX8+7XrYW306l2+pkMzSH1ZekojR
2egIDXO+e58sg15ZDbYWjI1XeFgHAWarnPbbzQKPPgwgoozBdCBo+2vveufv
9yg+PhJ668EbXxyssTilDyMvuOvHxwfeb+WAYCOUn7l7WyUUrz92NisVKZjv
BsX6+vSDVP8EwtgN3eaGOOZ2AGHnt6nPbtPoRt+Mm4eYBqZVge6Dv40IL3Wo
8O6j3YMigYEbO1F8c+tRoLF1YsduyznxIdfYmIKgh11BJuNHaevkn6kSY91Y
2ybvUHPBUdeW2vcjcX2AdVhIq6eeU/QTYvdHZuhPpNrj706qS9R1JABKrDgu
B6txSqcSbrPC8XuM9qIehI4QRjp9R7b2fj79Fp7v6CettCFRewS0ZWd0SE59
TIXQnsM4Y2/SBXFm5uhCGJ3G4mCSQdEhNLSobJIySmrIH643jLb+EJJfUsZn
Z2s8HkDUYu0M4SkW+rlhkawJDTZI4w1dv7EFdIm8IKGOholXbOeIWbEXHi4y
yjmPB3xfZpXa0lY7BdI603cMhJ4NcILyEIJ1UlDD3I3Bkwo9km+ziqZeTx9p
4uyqr/keATW6QjWRWaOZ9rgbc9/iE511isILKVLNij73sv3Mcm9Ryyb4bEcO
O+uQ7CjnP59Q0I82v8S7uoOosQNWQd0eHVegh7LIQoUr8kt0+vD8vBZchJTO
cJNlywkcRgURAlZLDHlUNK1YJxysgqCRN/X9KIH6yTYq7jHoa4rNNEwjesEd
ONKr+urefm50MBZ79AFo1S56pv2kH9fyXA3vBerUhiVeKVSLjLcd09K0Dj7F
J/VKYjda+8lJN0CmVqAq+Ai50bgXPEBTmRSlM5aOLq9ywBMl5xyaLFn6cZ44
0xxekNMEd3JrO8FYNTK6Wr87UpJLwpHPxNAiy5C/KJ9+KaFAJXPHjvvoXkCp
gZKLR+X5SbWxVZzLy+b23ap1jaNRCG03+8MjSi9T7zwca993sKTbPxqMuXkV
JRHA7YmCdTeWeJM4Negs8dtv/0ipo5rMed4rHCaZCkNLbMbf2NGd28IDqu/h
z8d9l11c6ja3aCiaEbwv444UCmFAyAUdtOPWCq2fynK1RppQJUhq3Wz3vBuV
fDIGiKbbJLxkTTwsG9Bppd4PbFGg57jaHqZnRDTCNxjO/46KJcQsFIUaejIV
4MmRbqfAs4cdVAO5sz4hUgqimhcQn0QfOwv8x7lUJtHF8cVGyGyrTriqANu5
I1Q/oI8AE+ATD/vD7IHsIH6sgFZWhwQysvRuymkftqwpvKvn5vqemh2J1aEo
PjaSSbrZE7DJWBxA3YFT1ojOAxlzd7eWtDsggp/RaAAroUr6W4HSj52HhtVr
p2qIA6AS/9VFk84wAMecwNljgFKoTLE6IDWtbwsmY0BsRsvUYpzrTY8nYLuO
vmvsXe34gY5lquBDbEY7G7sEjdrxc6tcqj2Fi529zS705LfOYVd318zaXAKR
HACIDkc98kNrFvRQXb9c3bryTguJ+s8yKN5aVkUzpQGZZ2OdVyxe8ev2AK+Z
3sgK0XgCgWHzDcKB2qUPG4dn8K/9yivon5XejMUVas3rEYmMCuWeuy/R9bRU
c1E4QmCthma74iN/AlJ//lKnIzfIZm/J+NAraD6IHYVbafo/JzA7dvLy38cG
38gk4x97pl7+VMfAodPdu75t73jgK6PGh2ZlgRDagJkVHrhGJb7FOwcUrvXT
JHJGkRxgDEi5q0R12ABFelcdHyFtTEjkmjOHPo/vNa/+yK2IZPiZcJ91TeuF
nu0b5GRs0i62i7ygQRQrep1H9IeVEnYIEW305ZHNOY3j/NfDe/OCVYTIsh5n
o1Xaugy8Op8JVnUIJIuONo7KiVF7vlQK8SQSEP1jbf9SZsr0poTRRwMI4AHp
SjBLaP2N1+89YRvJSwZQNnA4ZvcnmOgoxfa2cbOxlVASZ+XwN8WP2ch9r6X3
pCffoMceA2rji/HBQCPL+A/9vnr75N00H7E3fx0C3h1f5NwDquPGv3lU3zjA
jxUKj+0FSS/OfKvbISOCn7lPq7h65g4Qp+f9gqFfUdZaKG86nSxauqUtz+PN
+ANUYJRZED+c14mL0NpbSMkRTVowcZVyHnTgv+TuJKC7W44xaCVaI8yj7fvo
J9w/w+5KKnvxW7mTBzOUIuecHBwSaCBk/AgwvAZ796ohR9MLAoJ4dlf+uQZD
umwqk7FrXcObDawtzf7iIhuGQxCA8KwDfzk1xGgQaGYOXLMLtUSASZ4eVnKG
k/W7dool9+Xre42D2V4sY7qdxUmsGBoy9eVcr2oGItj0xl22fZjpTLLdDN48
V9GnvevzXEUZF8AGKFsWaEQG45TZyPSVF8ch6GZPhRcNbWRs4vs0/IIWjX00
tx3sMUO+bG33lwALbIEZj/6C0avtorlttQL1Jx62Fr9AghPXjIAhPSPqvtO+
upiSePryI8uKJ/npiu3PqEOEQdLjwgma0u1E1d2f0PAwnMFsC2YThAOiEgdt
3iDrZIQ3YFtBDRd+o8M4LVfhdHqTDGQuZSrt0YAK/nwuAR30ne0ttM08ZYU0
p82TiPDX5/8dpgWUSlH1EfgvOlwSlkjqN4E9AEDSyi5QeRMzJLt7UorYhive
sIikJ+Jrud7XT6Tx662PtRngDSE1dJwoaQBskkWDjN1SuoYKah8I5e0JHXq5
bNMzfUOPouUa/pjkjMfIsQIxTiQNuXQAtUXDKgy6KKL54apZIz+hjzKzAeir
jMme7IEKgdgzi0pDu3Hl7j3cbgpFgXPzgdXyNKq/QsmTENy/v+OWj02ri/wt
SqQCoB47ON5R2xVHoRuN1MS6hjBWMTPVQTE65WFMhXRjDZyWhdfblIotz7eS
JuMS2tprMj+nVHEmCMtWW62aisSbUco7VR30hd/eodE0s2GxGzq0QjKDF/DF
vZtTMVs0UoAI4lj2vLv4Fii1y0KPEEE7nztIRRO6/5C+1PzKfTAze+ziu2CS
a22GkFftX0aOgZTOF+6Xsc5xLFEeqbATMosdTqD0vXnXK3ojkTPB3UjmjNy+
KxmTymBD+REpkTZ3fuRZfRN12t+bD5AWBO4DeIKqXIGdDWXomwtzOb3a//XS
c1xmwUPI/etwu5JM7O7ddPvmNIOOCjdh+O/aTyjedRbdZg9eKGPxXilomsxv
PzaQo5xjB2Q3v4g4hcGN9oMv8bFmH3AWUNTxnK64b76k7WEqv/vNDasvFHRJ
CvxDTxV/AYI6F2NNN/YDPIi52gN9+/4AOUGnLXtfoUcfE5jRL1efWo0nNIDL
RPMpMd9zcpzteXtrudwNIzj5fNspEoAo6uU6Vk+Iyo89zwUp8Hs6NlrQNxvq
tPyX3oT8349NtacImorOwj1fDn3jy6LH5LXEgIwaUsX86/BxnjSIck9LQT6n
wBY+d130u28goDDnEP6yAVPCmOCT1SDFL/99LQVgDJCs/3Qq2lH5H5wPhDkX
YRXu7vlJ/FC/nFMoSk42IUUHTFcKk+Z0ehRJDy6I/qcJcjQqLODluM81mT1N
8H+Gvj8Mn5Kpxu8JZi0O2djVOzxHt0xyWn8M0qR5Y1J1o8m07I6CQfBCovbQ
VamY4ujF/+GRi64Y/uHAEPqrCjXPYk9KPyAccPiz1ZuojuibtVQH0rI0wP7o
DeJdCdWYGECuMei+ZT/PprHhOxj62KY8MpUYNH8ZDcBnelpuwI7EllKDPp4u
aod+X1I+EQlWu+09GuxiJKWckG3ZdOqHYOltmK4ff54R4Y2g3/oaPek1f5x7
TiD1s2Sqs8o4iQ4EPhjwMfy925Mk7tSEDcRVxh2h1kb6zQcu20j+oSy3LZge
Djp8HtKp7CENrboqS81yT8k+u03AT+6HVgHmLttF9fvqKBJuyLETslHtPUOt
DCRfyP/AFn9qm6lm7vgGBboaceWq8LouQcMRoj/rt4UlTFtaTXeM+2ZiqC8q
M7TVNGehreIbNEJsPYkEZ2zQo40uIIxuRYy3CSaHhIWDHDZaT1sITKF7HxT3
Cwe1yqx5h16SlhbAD35BNWwp31bVwmnUgyqPa+w0NXapybHMpAfl6VUQuYcV
Qb8wTSdUFleE4EW/sNE87y5a1cov8cAnseE+fO1bqJHCh25jxSihfXLacFVb
NuZyJQ4M3VdLcTiwh7ONNZj2XzDPfySAqCXEdlPDmz83unzEPX91AAcwvmtw
MTBxxw475ZyXum2OhCxI/+Gz5tfCNQktVLR7+d79gRgFUJst81CshSYblsIJ
A7v1lWw01wZdWl8/XN8H9g0p2r0qwO1NJPrlgdLPxcug4M8R819S3sAAgmQz
wjJkTa84A+tTDLwtU+P3p03X5nfJ1WSQhPh+AWMenoClriYVdf2XR3OYjBxH
8utPuShkCQAAhc3mEymFlr6xVGDfKwaIBtO5WheDaiMAOF7+ZPzR9dXADOAD
9Op+e35+KJDEgry5sEXsX27lYWOXWsL40O646bAjys9FpygoOvN3p8mMwVwa
xGns/r93CKQsfcf9ToaqSPhQ67HpbUByDIqBun4grwNraVk3qwng0vN9YTbi
qTuD6almLoPSyEHWb66OgMwLCfiQQifzwRtSZBNVlDpedCybxXKqB72R0eMN
/95LAya0HhBJhN9wJ/1wDzY0LmDTEkDxjT7ddaqGgfr66+2oaXctn54w0qpr
jqL87tdb2pQMbdW2VhIi5OeL8CRfQ6jvWofLr7VGynHA8DZ5939mLkF7z4WK
9ubEl4HlZZCNNKQCa2GujWrb8xH0uMxUFhif4SR/nzs0G4c5gXIg0Jaq69kK
9VFBagqb6yF4ri2SS54xmRo8zP56FlbqjqlPxMm+AHmJ+kvNphw1UlIRce7m
nba5rbzco1ixVVIMrr+PL9rqK/zVkfp1K2LB+WM0c8EahQZRd5egjWcddxwJ
xwoTRQDwowUkri6OdTvF1iV9q4qdZMvxyZV8MBTQn8NXKGYptOiY30PDWPKq
O5gnWDtlhMn/ZfFQOBkg4i3swwRkEGwJAvlHnv3kp0dSHrgCtFwRUPBCZb3s
F7eONabhBSs5scjvgYmIfGEI4/i+xz7KzcTTFU8/6S65cn1vjvuo1lY/DLzp
gfHY9NicX0CoBqTKGd8mviMM06IbfmvtIAiPSzdLpDKhGyMP6HCvfii0+X5L
QIzeCU9hs6wGicaP7FajXEttd/FQGshAG9Fs36J18pUO4xo1O8lT15lexl9+
5dXCd76MNKjXHUVuRya22n/cJrwVoEExp71kIuXbWrIfiHQhUxzS6nEcP8qd
kNj0GOUNAttCinYaywkolvwlq+UZyccUwLluaWfePu69kONOj4yoJAWchMrD
E17QbhGW0KUm9MRVokVhjadaRfN+an7/xQvFs/aH6IRkZ3XLjeiYO+JLQC2G
kpb+M7Olc+kR6VAJNFXZmuUJxJ52w6DbUmLtxwOtiwxfJodBxJTtsNhgr68+
euf1T/3RDwtiOAITlolhYKx84a443qvbz0SfH5+SpF2U0O3Gbp7A7bQnlyZK
tzVcb7HzLo8SJrGOjKsDG0ZUmP8Fgeoz4j1FRR9sTywySldv+hwwj+2CVLhB
U88Aggv/SZDAMbn3W7deE5W/A5xeHhFYADxmk85dGWLPIPNOuuHEnk0tbgAh
iJ0Wlcx08nbKDHj4gm15FaXX4JTUn+bwhaCiSnLSumVBfMajgOzwZgBvTB6J
XtT9S8KdAYYo0en4/5yZ2N2HeL6Ja1o2hRIm4/2fXR2nuASg3j6R4BUMBwCu
5p7zeKviLmU+uH2wMz37wbaBIk5Gave4mqFyZKrh52qsHNaN901YGk2I/i2h
khLVzJTCvJoyUGLnvz3LSQppBzqL/D74KZe5WoGMW1sZVrTe0YHXUs2uYp84
QIE56nD6CpkDezUEUfh/zTlpvkQBPgdmDUtYE6D7XvIVeDy/equP44PeSt4R
BNfqCO98XZCcFshxfgjzL3vUdMLpmRXK5vbJAhSuDmCV0ilyebjZrq6uC+Gg
g3IckPgkRY5k4u+++J0JQ2XzfKtuSS0JGo3Ydf4bjVue4q81YhrIH9OthmPC
a8VSmkiB+77bG34EA77oXD0BOdjUSECUa8r1EG7D9GvWt0jbfBVRG5OcZmLE
i6TFdsNGX9LE4S+vVQUCYNvdke6gJ6V7/8pBZNw8auF/jM7OpjaT1pVTPpAk
aI1FHtG25K8nY4CXw8dnAA02mhwGPxWvE4AWhrilYZbj20fhoVwYKGAfD0o3
gFpzpwadD5MPcAHawrpmHg/RKKUp+chZhI22A/xgeeVEjnCGGIkETntfUhKA
I3I8Q1DNOKBy0wtZNJ5LsxWRUYIfV8nEUQ2rG19APkfNXodCTVzcfGqCidKv
jODl1Br2dmZQAVziICYntEvz5ArXi3Wv53521MdgBwe9hpRxP0Vny8KyaEt1
l8YGGCUXNUqFrvLzkMho91NvDf5NLeBn4w2FldvJ1lTY4xeH1bTDCXZACEOX
9TXXE2vcAz3AP82q6GlBj/YJivJYXeUrcJeArxi5cbd0Oyoo4O0WC6Q8ZPM3
C21mYVsU5BbJZGB+WGMOFKechKsTV7BxXNrF0/oqsIs8uSmh7/Qu7QtpsoV+
/xy1kGqHvk3yUq1PgG3Sd79LdI/FkWblNPVeVl3ejJzPjbwCgXWHhw5dZIAz
Z2GUdR546FRfOiys5nLiVz+IBIv+n2+7zQEtAlxWjk5LZGdkWRU4knBEjiRT
Y636vRwQUrEk/Ge7qigFqgBS7JcbTdXR621vd5Y2EbD+yJpSFjpzKK1DJgvH
MAWIIWx6D7wUt2FgyzGtiOI0l06ZAy5ZGP0SL3yhk5A4X6wfqW3PFi5rDmTL
BEbH3riOafnoO1rVFg+orh7kdV3xRmdRrOU+vxu61udT46K9EKRf8ccecXVb
m+sNYcf6mj4JfNMaeldDJoz5ell96EMTXY6nNSbWiFXfRKJrwrh0SeMg2yyi
8gz4YaqP39GrvOCn8P6HNoCZeqtn+sOGPXD3NmISIMo+OgDnbqxC/zUDMxgA
yPRy2x4JP+QTzvA1iQ6zzwpsC4Oy0+sBr0JFB0/UHh2QEwEnHbPSBu5Hqvnp
sdmbnwxUqHT053htyjZvhb0wFftFiVA8n2El4VaJfNTaWgJfR7IirhkNz7Cp
OSrLyOtHRLVIMNgKcB4YFw42hoYrcDL4Zl6UgsFh4eO+LlSbVrzXvFiLHteH
9k+C4m6QlIHTKq/7Ex0kQQUMGz8v+HcBJQH+E45ccTLuJTEbvvO/1zWlZQdK
ueEZgLLb9vtbLpd8bBtGQU+DLOf7aQViiDdzfYxrG0qyQLOoMfzeNW8gIS6u
QvFjVDcHy9uq+WX+eeHBt/2mMvt9W/+s8wKQqP1eXksR5zqbcUSPqCikO2he
e5Hf3uU7B8MK0jtNuod3yi2mSwGtoa6+WaUNeq2+wynmjVsR2FKOJ/pzcibe
Si93RmsMKAgrJFadsMx91wumNLHlpeTVmexKg4cKVrI9Yd4DKdoqmEoSUDRp
8++4VWRb/s6xVyXrkpCDXFdyN+2qN3urgYusmqFXTyX5cjlBz6S3GEsWI0Pk
autReMsAhZoARqNNarQN//Vo+DaUrDLwdTOXS9FL0R6djV+NOku7JWADmiSc
CFL+QR5a8Vnles33WYG9mkgFng7uG1YaHLOCPeXqbQwltfKwxyD1CVLbdRGB
hBSs2yQgUBAf2g8hUgbED2qCHxK3UXWrLfHC10pqGKiNjC8SxaaEeMcZSg8w
TZCPEh0REyTG2g4dsNwTlpOIkvgkCRksJM7bqNgiKRY+LC/v87KeN5wnC6wV
RF7beiMTodCy2+zrTqg2mFMbwMFs+RySKmHjJDNbYyiw2dmqD6qo1NqTDgS8
iCO0aiNZoznFoRHHd68MGDIwgAlh7ULQYTWX6GDUAnTDP8akWUYGEGFmeE2i
knHya0moRVgVg217rR2P0JlXClE+fV3a/gJXdqN7w+6rUDpfeN5nE/lCQ4EQ
gj0NGSBynWIfcavcB4MQIcIaGxl+NBzvP+V68+JYGEyETc/CnSpPLaFNoWrQ
uaR3vmNQqW8w4RfiLUcTjIpLVA88ilbQDUdkOcXnPdeQMd7oMEbomtnTH8Wr
hI+tnAyAV4NhvplO1GifrG0Lr844AF1NYbw7nMHO0hluV/enXKMb2vh/FwhM
W6FG8B45ALd3VlGIZ7yd7MPF9+s/94LRBz7caIxhxpi8KUJNBpYKf/xHDgAj
BpfxIcgKZSziHe5NeKU/u7kiY/Mz7xDXouWpBHdcgRbtkcAcFh3YWBRsrt/A
VIiEisw0GiXverXltbYgwto8viAUW+KbbiZyspaTLquzEDuhX9oWVVeGhGpF
XhI4oNxnQrFeJBsLyFY8PIvp+JYBdue/sYh3kMCvHhiuG6pCt4L3nEqy6UW/
l/fe9dMv9zKjo4Hmc+4LpQbWY6rGmVAcGntYqOKEHOV/552eIdrARRP1XJff
x09c2thvRwAlWd+nYmtn2hnmowuF2ZqKcRDdCbDwI/3A4eQ5vpFS/IkT/Xba
6tZS3GjKKovvPR54zju6lHVbnrJWlnFtPOMnETnvdGjfbZYFTbUE7pr2XtaZ
0MiBKHtrls7LVyr7B/X6prXKlwP1LZD7ibBTU1bzYS5E8cuHEELlZFbQw5nt
xbitjinlZ3K4FbfU43NQjrmc9ECVytEqH4GIyw62edCwd/zdGfD5BGs02/L8
Cg6SNxpI+1XHdDsBZ4HNxAXQcFxJBPCrpmczdlod45Cbd8vSyYbLRAjYiTxe
9iEJrVeIdMsna9nSQ/C2YRdORR/p2S7qp8m15/nYOG0lisjAdL1z+i/+chE+
RS3QM4cDpYBXrFR5OgWXcNjzCAbC83qKcsaxP/jCJZnSg8nlCiB/0bWJpP4f
VqGbTCYQ6ghdR8ZjirbCEYZOewPS2SW6k/lmVY5F5dXdC/m8iO7cqoGNo72e
hKvub9NHMFqB2csZ8tSZMZzKLOvy79lLd4GtmLSy0M1upVoqKMEkBvg/p+JC
YgikmWWHWuD4mbJgJ5Vp4phr2qcrDdh1qIuoakpZZ6pkGiYJ2MbqFehrK/eX
5kV8Sll9dtJJ4ldh9HY+o41e/gOOic1NW6+JGCa5nE6l+BgVqPDGeGEEzCsp
r9Z46WdUMuJpOD4VD8jlBqknxRmhKkOxYSQDPvoAEZ3wvHb9Pajz4VgqzV+R
Xl+VNmj5HLP0sJxx3DIrUgkhzbf9mjL5eg3541Brk0l8uBNcxRdXPvFQ18gL
1slsjlyKBiY7mmejcunmcrPAPaaKlWmz/ZkoZpZ63b12YSyWwquYv9pUMu2d
eki2bDSlY4Gc2+ydaVAFjyo9stTHNhAeVSNGSrOmegrjZuUYCdHHVttl+Bke
Mezw2YSx+uBqHIi4lIAHNsmIZXhweChRQeWlq52VsGXitYSboyaw94og4VaK
Js4nmzmkXvD1wqUMUFRPmJefD2lrmfD18PPtB5/MyHgTb1+m8KorAV0emezg
RVwmlgumhgWBxu95WsLyyaxMw/duH9yiJGVSinZ2Zam5rk6W1c9yMV82eV6Y
DtIWT7pCvYU5+vSSnQrObrbyV7cv+Swk//LT+xyCq05wBRpeYkYMCuBDdoWH
0MMkYkeCOiDvFl4tYD6oN4XYd57wg8jAUZk06EynHo3jTuWRlwdduxpTgExh
Ia+6FU1RxxXVClDlbDa8gBZ9K1vrWqpc17E9hS5+8cvnAw0HtGAOUpqi00Yy
LFxtfy9o8fCu1zp0ox9f15NSK4zlnzE5/SvYHMUkmZc1vNOuscqZ0QJrzlBf
JKUAYEJYj+WhfoEoP2tU7aE+yi9tbiPBkLHqVSiSx2EUHwtl4XWCFAvCnPAL
nA3gNG9Z1e8ofVH9DwOKAbMzyoU6/8iQ9OjK98xGf+Y2y2LL9HD43ZVhkOeT
7mbZKfaPdbrQQZDYdPYC2CGzDbMZDdLsR6wKIFiNQXX/EROuMCKdBe4zmQl0
fOCszxqUtxZ+WpUxuaUfVLzAcUfzZwXrszMBHi2/BVyh97pCa2NbsC+orJCi
8vSI3FDYbR4rQKS77K0f5GcGdZbKZh61G8DpLVQ2ptS8umjF9tx6vnqiI9OX
JBm5BkzYY8lTbEZnPMEs3ikcEqqeaA2fWa7eW2DRRzOLpMUR76ixS3mkfyKR
dZICjnqUKDbqdsZGCJPY9ctxxC3iEMFPy59Y6mmudLZ8ajHs0O9t8/pE+pY0
eafdBouV8YDX9pdEfpWBMwGNW13BgfxZbc5MgbJet9exuuO2ecAyhsAQngBk
BCBtM4rq8jr4ktlYBYQKBCyuRRwi2yoMIfnKkTG6SxrkDxy89qAmTFUp9tlp
idprzu9sp8/jvM1ZSI5pZNUph6UD94Re0XQsWZ5ifGPfoqhCCvctZqKebfUk
gBzmRG7jGGndnYjWPPmNoqqy/rkDdyIvk3p+G1H7JJ6BLc8UYAPTnFbzsL5w
eLVgwRKBanrK40K/20KTcu0uEujNwNQz6o2FRmgxm7P6it5A5KaKx/fnnJrF
LNoMuS120u2yzDe2Wmm0xrJ+EvF9ZOWeEjp9PDibn+8SCbR5atSQ9HMN410y
25XTLDVvr30JMtu8e14NSSwOQWsFUsHfGijrQZZjoeqlhALfr0s73oj9NTMk
DcwKzsLHGFJhBWWYSOc2lQaUJdJPdncPJFHlJ0HBfAV5JxLbuNF3kgxJbnYc
0zdrq/zpbkE/BF7aAFVDX13JJl0xGjuFkZAFW5+JyGIvohejgn/UdboFr7Sc
p+YMl9Uwi+L//qZK20U+S5F1QDHuDy/RnFlo9tevxzFnj+N1kRRGBX84XzFQ
fR+Z/pTs4QYLqB96CkutfzKuv0qItIBnqY4UKZoHFbv90MBlfaymxaxucS15
o/jjR8zSlG6gMFokRkp2057bxdbI2MVAKnIklAf0TOuwKsknDyBOTN2aY+sC
zabdaGUzal8E9+EpvSAAf6s4MEBTCAm9JNtyKdMcqIB/HbLbSak6kVnhEaO0
mupGz5q3j8BTy2BAliuzC1S/yEzyX0zeXSzzjN15IkkdgLxG5tsx731B66/a
goDf/VkMlFKtc84EPX+e2aWbXccZqyem4sbqexsr8zTuHCA1dKQlqYa156jz
/WwQ470ybLbZNeU9ZUobwyDKRTFKjKkTXEryJ5XqPaVoUmsY5i5ZmqvaXTCX
4lbUg7/z06SdTnR9c7J5cznqDrcAbGfL3hUxeR1WvPH1KgDDCah3ui7j53Nc
xjdf3xzgrfUbODNpzhRSIt2z5ILACl6MgtmWo9mV5jBvuBepb90NcALKJFM8
oP9fEku60gsr05OjNztRUBUrzs5ruG3EHPONpPQNrdqbVVwoB2XGX4ccDWzk
PlG9ToTJIaLKjJXmQAEHdxT6BDa8g61uhvYwyLVib400caSjG1jRJrn239VR
N03rL6+EEOgF4fdwH8gzVn7Z+bxNVJ48NSB9bdli34r7DJ7Zu5PpaK04TlRY
8SdLdNcdm+b1ILhRCZ0pf0qo5PAPrXS+DNrPZOAFB5ytV3Pwx/eoCG1u3Fym
WXsFwBvwmgo7dqPKfCg+8fOluDFF6w/mzm+CUz8WirgEnDRBxnUTnIwPZ29O
nz7rQPvMNdYiHX+9thtLB0WBfIixlo5HbzqmuzQExMgTiSR5uejbyLqovtIE
N59KyQeFFFalZ2GtPnPl/xuRN77kYOD3nf7rPExcFaT2nQ3HSBaiURjeHpJq
g09TA6/VpuL/wyJxkM1ccEyz0THgFDoi9VTy/06+CcHv7Xb1RV4PLWWw4EGt
2iMV0zgzVzJs2Wv4wQhnpRcVzVNUzwNnieEBoD9jW/4k6YpZ6cDCAWZmtZU/
W0y4LoWIClps3qMi2SaMw1LbS34zOZZuFGEL+jIfVOD5VBBUwNZnGlDuW4X5
dOZACdj0wYua5VYbuk5bVgxcuNl+o+3lWQs2zyO1sF90ileZhEbq7+5kqo8R
hVnus4Peta70ZOYRhbP8mQC3gbBcJXmn0K1CJ5L6FEG4XJQPrw895OCAFevf
f3l3G1hnd4+Z1NUGE/BUt58+GYCGKpWB3taT3qit4KfaraJL69SIGrgi5Rse
hnvEvGuZJfAh7K2KnPpHRGQDThCGTr/5lSk3uYW9FsfxvuGwFci7sDBoSahD
lnvjzRUqc2VG/FDC2l2NSoladBNh/MGsfDhKokc4ksWKxOHXUTDjIAOSJ0o+
2/eN/AGS4T6kGsCegnM6UFqGd7hdE8NQ4yxa/EZhoopS9RovoMnCEj4AL+pn
dFFbeHTffZVqxUmUzqopoJJrmDxMXevp7/nMkx/+dPlMcQpQNmLdpw1YF291
6Ej7ckv4ZqEs0Ic63iq2BhGENKzSstLO+MyUESjVGsZPuVr6lYBXz/O0Idsj
B07GyBXFMaSPGrvGXHLEUIVzhFlf2Oh+QRaejKgNJ4vnE2YAEgKxczlS7T+u
D2l5NBbnoCZl4n2RB0VpLhs4ka0LN+4EOrdj1RifC7K/tMDcekgPcs+J6rHw
bWE4AC+xF4/mN5Ap9uvR+MCaSFzyLoHhFxLelQ6ZxaudldUy4ozfV+P6JAOy
NE7oelz4zewS22UCRUfWTiiuHtCAxIIjMlByfx7hi/DvWqbz/namWJfTzbxB
Yqw6XHHlwFIhmGgmpna0SIizqhoD7d4axjV8jWVk6sLa3QYfvKCHnRoAhlRN
f+E/7UQI2q4vK9ilKlP1Y1RvApRWip++FLEBU3kALrTM42bXlLfqA1brXlzD
04GqcIieGJnfS/Ned3ppYKYJnQ3L0eVo6zWYoDMHTZS3EF1w9NRrNuAF6e59
8xrb7BtB4+W+u9PmtwCo+oH9uv5CM6ySxNLycqXsJzRamsP9GinTnGFBQzgP
lhlhHxokUBMUj6kMCZ1clBUcsBexZ55qDv2uW6oU1LIG+dAfulQP2bsxiR5y
uwm79YbMPUEP7f+0K0LvMJnPHYi5X/LzPUSAaIZGiIbuIIWM1eL+2vh6H7u7
1tRwytpy/xVUOoR6zy/0PE1svA+t5Hj9eJsyCaMYxlqVzve1snJDFMrTry7U
R1UV/NOhEIgm7QkNzZUOnPkXAX0rZRTObMa8yln44aKr3Q+0XX1COc3Xangt
ej/hHBh7mHxCGg9he6rjC7dv73j/K7OwVtZfLILdONR/kKaKZpjV4uNr6zOt
OPBBbVtnPCgbFxRQLb8S7d9zr7eohKU177OW9bGkgc/NFu1ClZjyj3RKXbFY
JWOSdbaCMfpNbvPN5aQSCjIZhwbgx0Y74hkSqi1YfQUFPdzlXM0AHG66nAKw
C/CYjExydJ3bugYQI2aBj7PJlzZvuaAhoP8VE9nO0oqsB06AVu1twVe+riQO
xmV7Yq4BudbQd6+DGgkr2V7YFgYH6Gz7X9UVEjjyl+GMpo8S4FjNMB0XkZE2
kL8vsnPZctDqkTQAclEzNLkMCXH/cPiKk9tMi9v9N6x53aVlDdS0TiL7AHdI
4NSiz1w17MmN6tS8510BBqUJf3Ie/4t8Jnp1MCvIvv5BDEuHEajmqUlcKJ6N
RWzPdmU3+7G8gNkuSgUu4O7Y42O0KmbvpfCFJT26Z4BSo7A4d3esK12VcKI6
8WVAUWWG08wDQ02BTMOZLdDRpt6uRLVRWUqq/026N95hzkJYG7ArTyyy9BkU
zQGdfZCvkKlurn+EHHPaWPJp7/IrJYXiMgjTpFf4LvTwswJeJ3VqFYV20tdv
lRMbBQfa2GjZQX1N1xxl6+nmT0qKKtqwdGWCnPoIB+D75YGjpecSl3o5S/7b
xLpH9x3VyragsRQ8WGkCjwoBfFjhKD7V13WIB6ZDtRM2t0/WuuR/gamal+ia
3sT3Ks9JoG+LoPQfqlXk5wt+rZSzWOfDELVNkOzvg+97icRV5Q+qhT/vYdRg
3Fsm73IZU3e/dQz6HbshQXFI7gVMhL8U/3CMRZs71oqdJ+RTVQIXm+/z0w4c
hFRyZVdqhIDpeqFYHKsqjlratzViXebG6poMv6/EvOm1nksnJTykTwRI+/6S
4glB48OjEVijwwS3iqzsfbySH45fH1uhP44SD70CqYAWMzXVdnCFMEdxNTaX
n67RTGR5DzS2xagcunr7O8UstF3+g+DUjKQQUYZg+FQWFQL9FI7GSuS9Nzs4
NLT2EoIC6scVp49hdihpOu30PpMe8/+pkN2Um9JQCPp98Xsr2t7aAU3O6GGW
8lbtBLeU4G5xmUfzItVcR9Bb5stqwkFciaSfOfolDm+UScwGWMHJimEzd8ch
5jizLv1ucBBpqGwPno9mU5QklGjh3+dVQT65KSe84UsNBu6/Xt4Y5Tk40PLs
ysRmgRrpUlq2l8nVjJF4J+7bfYZbE5LdrFMeAtSgscXGDZnGgxsQdhBe6yBt
NmhWEMrNypV2LkuMYiR+mpcLrlUtnuZhZihQVhcajwnAhxIlMJGhdz99vWaj
mYVaQi0Y3pSBqM4Tl0Fuz+JKOHHNVXYjr4TkMxQMoq37IwxSfx3ilLCDWha+
H9XIo2nBM6jznGSd4AOuH5u03o7KmQJB6hZEwCaH9dLU42tkMfRte4jGp4uE
cv2bZXt2OfyL8DftcWyWEsjmWB53a6IwaJNKjbS9XxAwO9AreALu5xFfYGBA
3+fq+FYk8LvkQb/goNqIP56LCMnFBZFzwuz7J8pGG1miX2JTMq0mdKL+03OZ
wmt+5GqxouN/rWygVzzzteyKuuocr1VTxgoTFFXNt85VlQdGS7vBC28hLmce
XOrSRzMCjMfkR7ikHBT7HLWA3MUx33LHFLVhPJ1cKu/c39lx21fbTstX6VPQ
OKYGkcJxp/QdCGFjdrxMC4rxkNlsX1BUmdwZJnDElGwpbvjy86rvT7smR5Ku
sOgHqCS2ocZJoLMw+ImdlmRD6dL27ideVVl2/UMxtSdGiNUmAVpQ+sIoBfcW
4LVSm9e6kDHrgrEh+gpu6bQpqltZ/fMmGjNFyGzRD9FsdXE1bexvjR+7EjSj
Hn0YWBqKQirJ4JU38nhBBZFVXN+5iym2F76UCPsEO8kSP9DNks6hbCRR5E9F
8VLlG9oa2gIL2YSv7vfGx/Euuux08y9uGouqbgvzkClyQ/hCmI2rL5No9i6l
RQllPHi82zgFfSMM13a9JDYtIJ6oIyWKGbx9OUMgh0UalOinDD8CetUPPu7T
O65iYFJPgP0SE1WDSi3X8tfOKy6RxbnY+jHr8w3wBefjP5D0FFy2ASwubqn2
nDD+v3qbk73I/9gGDfJ9gIj4oOb9GeLJGdnNqRp7buVhns7U5WWQOXMemgYq
giA3FhM2P7YvEBshKZ2kfj4Igx9fY8RweLF654kkS8nJMHKTyJ35U854nMfc
/H6JYivvrJ4dwZoRlTkHf24JcPoft0ahmVoZlj4hWnThrRnZL/zZJrymk+rH
slicXfIKb7WNATjZxYMIw7lLMcx6c46K6bJI1YY7zbabOAcJHwp/OG50G96E
0EbwNfQWjaE6UIFpHYBkQlO+4rpuuOl9WcJpD1n/KgLVqtMzUEDtYlF66CHX
FDEh5D0bv6T6kku68YDpOfsacnCdYIv0cew2Aj9jLN4pEEdbAImyKU8E1xJG
jQV+hYUtpOWztPjXm83eRaK4aNrF6tuSttfkKEiakQ6iUAx59DQhgZn7MeWZ
E4jelvJIg3HcftPyi37fcOBHZyu9QQFrCFGUo/vMMYOqrQzM45oJF+Kql61F
74GMEzdSiDQtOZCfe7aWhbpv+s0DFycChq+RacepN14Op+Efv+ep5ew9jsOR
wtu/SQnJiWtX1EX2kgPh4pw+WvNrOslHlS0fWLIl4QOaPcF1jrpLp1L0a3z2
K6usGaYHbAP0uaZocVN4rW2pwPgKDxyvIRjI0pUPJQVD9S9aGGpL7iqzcKTj
4koHZ/YOJeQEfvwyP7+Ifi5nR70vCcezeqJKbNpcHNJ+OMA+4TjK7vGBwRTS
Ln73H4/WMrv2dkp7pdkGhbe6ZnirkDSbvs603lYpcYpEYJ+UbLyFen3SUFiN
rrpU71GOVt28p/fy0e5MG2pm4KXnkqYV85Hxgp4p+/3Qn+ItG7lueswinWpk
XQXhkugx9qTCVyc2V8Cv7Xo+GSJqLoTgNN87wF39RZ7AIjCcOY+hrOwnHYzY
gFORQHzsNdyIpwEi5iRqA2E9CwpSn7x24SYCNrkwrgpG3a+uiopBUAvG6Jdr
Pkf2H3bx8QIkgtm6BkR9oGBEBHQyZ0xu72YdGiGEkFBvlFk0s2fCWZdOXHsc
YbAM3iTJy4E8BN1TeWG08hT/nutr+FA9WPHxynaGP5y83ci1cXWHY3UjXTm1
TrLvM9xZx7c4ouxI/6AstqQipeYXFQjRL642w0MoD22OFQyjarw3mImo1q5T
w8jNlKQiLaUwjwLWByLf4pKWcSrwvsNjLOPR4oL0FO0HCoKwNaxI6oHCb3MS
qh7NIV5KfMikOqQbAKxwbfkDBxlrG0Jvb8z2ZcfzHdjAIq1OLHSx5uhJbPTw
dwJoeGyt8LWn2IYfKsVtwGxmEa3i8axFh/9NtnjfWxcZsXaHyFh0NF96aoeZ
MO7B61+huecS2cuw+qrdi7AkkxOdk4zx7PgDm1ayQadc5VEscFlZ9l9pg6gH
yaBIXpd7DGiJJ41IALcrj95JbS8b9fFJtYFAIQZ6A6bFN9s7JPm6cM3T44Jo
KwPcNMpuUgCA/GOVkvmGLrC4SUFyuXBSyhZNp2PTAUTAnlBrUpHKs3Ets/gL
G+QiHQ/Tc2H5FK5xWYSqGWqsZgdPDrZ+xx42R2he/E39nxBlQmZh6yOuciob
oJ/UQBICCUFjcS35+9w8vJwMTQhVJwYBJKCsa4ELMLEiIkh5x8J9fi/tnr29
80amYyE9HJGeM+9lcUOrTOQRNTKcOifIaDcbqV1OpTEFNGgOb98n+YmaxcYt
Xrq/HbPnwyKvq07U0cgCVKR09eVS1QBSbINeoWsPPs/R01OCwfCYf4yWaXuc
I7UWQRUF9hfZtFNnj+FGx/iCKgkXJ8xs1rSDlHC200eTWwKrGcfcWpeLsdH9
Ohj/ayZwNRA6I/JePrKeyTLVER/dcpi1mW4g6lpP9tLZgUX7xl3ZoLCEYvg5
oW+W3NwpqGkTAtTJZc1B9DbHMszfToPzlf5yTuGsouvcYJABAXZ8L0uOQ86c
N1xZARw7XT/f2mazpuXw/lfIMqSnhpHhQRopBzbk2ZEuF+d/4x5lvsyvbm1F
UKYFEV+zZ+wSRZMxuDaD6KjJAMObVvmhGOGysQftwo62951+k0NBAF9CdTDY
y9yCcwTNgqIrmhBCT63kulI+h9C4rlNxmzQaLH2EKqwmSRh2TC/gsmYJMyxo
zoIQIScAh1fIsz2siNbh5dM75jRUoLE0BgBUeR/xzL+VSkNQu8ECONBN8gdM
E8Ah5SDfB7oAfrKNizwEFJtNVATZGo0Aa4rVFj2kB1H0yU/+me5h32AMe77F
daLvXZQQvNgHoqm7+J+6ue1DgF+gQmIdbHKCauA64u4YOAMWOVbsmOqeh+mm
SCh0rqgKQidGIvKeIRV0ODxxxirbJU7H1RLEHFHoXKZLblQcntSrEP9ip1tC
g2fXgBNjJxyHszvDMWUfewgoxP4IV6sDnKke9UdaiRNA7NwaSS3hf99eGsDh
/Y/eIM5wrQ4BlzTFXHDgIGuc8DRDtMFvJEISj+GJVu2BwweAU8ondOOOYJLP
nfwuXfoI3VDP/h3YC58biNVixo1dfSEzPBt+gtnkWmQRLMtnaVQS03qimCrb
K118Ja8YjuMH8jMXKv3SckV1B6psR1LHMApBCINPu+W+8V/WGuEbD6d8F4oF
YXUxeA0JMuQPhD3N4GYEdeZR52f2unsUlMqGsZnAu0ExVS5X7TYUam2PGz8P
vNghIYStR2nO29d4AIOVYAkyFeIzpQjKbNrsW1jxxtSvMELnhLepHEIM0HJv
sKEGNzteKxgXw8AH+K8E6FhujOd95aGE0nwC2DsW77kadnYsD+S2R1lscIDZ
X53+/CT3HPN+thX1+DmOlqIfDkOXAKDp2zUWJugpxU8e2B4Aj8UOA1Pv3XQN
m7Ow8bI/GKX6z3KSSD3cxeorTjPyy1dysWrHvkWDeCekuQR8x41j1KaqC3fR
0C+vRhpKv32Qv/zPGkS/AefinBQMcxgeXGnN6CeOAgZkE5kQqzGNpjLkxMx8
h3+gr+mchEcj3Bu/iygWFdJkCKuinPA+ny1h1pGPcaMT046PQcB9geY7wskY
3gdY9C94SInCxenK631OM0wbyGkuGjSLD7pYrw2MBVzgGus/tPOryVCvZ5Lw
88iDGa49tis0WPapoHLTM2S2DiPQpM1c0UAz5BXKOyg0oZaz/CLuWkBAoq19
NjP6UUvnXeb2z6JZG0RH1AeT4S1CzJKCk9mtJ1i5AGFYETfXAjOTqxH/JEa7
w3miFtqm5yhiZpFPEscOcooSq4M63J5UcmTZ8UuhoVOUvSsDgPNWiQGhuM4e
Et9xrei1jx2D3DdUdvH5bZ/AQFYDcr/F6hxZvjauKXfbBINnS9/uat29eG9J
xy3dx0HnQ4VZZgd4a5X+oreuYnMyMY2PF/gVtgIWym5YPoC77TWl/T7iZw6r
uCOc3GzcsatDem/oUe4w/u5xCrlLxpk0vYh3d3cXgjuY0TEKdKlFi45GNJ3e
dXV4TekAaR1Am8y29JGrMgrbUI3VYv8VW+bDREugrfKiUV1tlXA/HO1fzlUg
fHa1QUYcD/vDTBTw4RdZviInsZBnowCXk+84ol6sk0TeOULAjqaahOLXVexj
9dscnAChfOluLXZnmSmBb+gjsZNQ6LtGp4HnJTiD29o4GM2sfU6UNm7Lr2O8
r0JGXWzwClD8RgjyPRrARI/ht44ZjsN08/nVhWILSf39z2n5EwAvsK/dCvvv
RbxIHe9NFZjxghlyc+c6uLkp4S7HpBvHv10QRMVPJu4aEgUTSo+23qfvZx2u
SH4T99dY39w1vnkG4dMS/pMk3o9uC2EWF+vPbg+iW96iMZ0kaA9u7UY2U7Fl
OR4/jHnMUup0BqeIIJbdfx4Tc6SH2QHiI6ipebbn9JfN1QW0RbwL/8Ho3gYG
M+zU0qQQ2pyXUVYjxxARbc8mBQchteHL4TcBWXnIBsZXPJzSjKrNtLcc9lb7
JTEL3I6aKMtJZg2cwu9nkmY43SRh9L8MWRvudL2O0w+7JiKMy3LnJOFZbMhV
uTzgYxKJU4pPO4jL+Fh6Cy6z+81l/SUqfmi2V34V6NXnd16OaolnXfAZhGLx
3/O4wD+cLz+v5/mz9tjsoYLTdb6elY9xqlOJkeOv3JB0s6gYsvlHCYp3WnMg
OYo8eDaqgrn1Lyxd+GUtvOENPXJPx85htLgON0GBHV37Bmme54Qv8RPlRLAa
AJw2n8exFdTSkOdLA0kGP8qAnsAuskyGibqPgJPaFL9+1E4nVcwK2QHdpXGY
1CbUCVQkQkdH2WkDkOgyQfsNlE9gz+LPPJG5meWa7weFCTr8zIvgbpsuzlv1
tApPUtAKRA9AymKUvfwH7VKzioy2R3N+4sBg8KttdNf71AyM/hfkivTI4FyA
3Df5LrE1mygmayZAl8aYvxBsgJLvAURtliEu9jBpVtU6wervA5Nx8zGa8xXe
heRbXlbBZK4PiYefG1KzEY9ouavm/uxUMNA8MwN8dGOvwXdw0ibx7zenVImu
19DLycO1n5BJyMCtpyzNCtb04r1vTz0Z5VnVFjHqUMBbNfgN76+jF1HeQwRH
uRTcxpj8nJeTZeDhU2pHy4mdvwbPpxpAauQQngtM983slfAmj4OhydfkJjUK
AB/c7FZf4qTe3UbXaJvngi+rgOubdCYqwsVyk7RwYdAMvrqkub5Opk78ZybS
ciu7aGfsrQ60OZN5oZTGWG1a5S/SJmqUmgwFnL68i2zq7ZtPcAYCG3u0DHtc
7CFyzJW758iy9Su0jZodR41tlRyEz81UVXDhzWNJ2pXghgqSEj2Pu6gFKa90
pmpu+gF7reqU23i3ChUj4XyUpSSw7UzFdwz443xRSC4xB2FMVSQaym4p7GQQ
uDjQqk9+KA+dZ2+ujDwcyO//Du0B9chE9dNgsc98WBCg/xYOrLK6cu3lsffl
9ZoiPD0/kT1JCAsbfoNbz2T/ZKkTuHav1KFa1tpddkkHLN0xPFyHBrvOL3CI
DA6FJLu3DtnGNLtl6SDXA89voKeJl02JJjnxbiRppzv3nyianJxilUL7/GI9
L5+z5LzoUETW+YOXvj3+RJEuyPZQR9/wsnRcgniJxi6EJFcPnNT0LW7fUHZM
vTrfiFUuAM32Xq1fdCiv6OMJZ0bSo+zrg5fpWvb8YEfHCVPdCsuYNUfGmoFQ
d7qrENdyoklEyau93Hky7zYhGzotEcTBtpdCk03cYCZgpptIC74Yclzlh4EH
Rs6EvCMjR67M5HSeaaGOckQdE1uJC1GOaZ7wmORWQY24xu/a3TI0sJ9/4m9W
kcc65fzb3UgbD9JvRcuPsGxG7K/HtXHmyj8Iu4EMhleJqcNARnmYoiFHxTDi
DMqQCdgOJVqYdOG7y+XQ+zbguaKs8HohEInCvrr0J/OE/UlxB9Onw7UhqTjJ
/eiioXe9JZgRT/r3zRkJrYYjvkmwpZsJQSSs2p14xwfCQ8fKJ+sHSCn315pC
J9wqQ4xRD/oG3LJjTgJsETb/gjD+ZpYB8Ab5udSq+t7XB9eQSW4su0ZRZSsV
l8u95bYfR8Zww8+jTvpKN09JMTQ/4bJQps91VJGOJXdrU6TY1ftroa3Y8Mdd
JaDUKywOn/hlmgIgKDGkJf80Gn04FLv6thP2UVaJDf/ugNgC/HTnuMam7Bv6
WJhU3XoMIoctv0eK8Xos0ByE+JXLLqW2nR2xNFRTyVUd6qTzI2vTgHax3Tzu
jQbOPbMsi3Xz/mzTNn+1ZTbjLbZCc+HzzHZlb1n9kKAU401zaUtszH9P0IXB
I3RWengPEKHVQKJRyknX443zsKnp6d3QubjoIDFhk7dz7ZAlifyYtSa55Tjq
Qm47jzPRl3Q/lz+PJiXYsfwZCH9vhHF52POM4iU6laH/VDxU/CT7TND1xq1F
FXpzKgqMfi10plIaidHL8LRK+9MlwSw2WIonpzjFFwZNE6hcZRKkqKLnUSKr
0nB/vlE24YtEsJuspQwZoqOlUZxylZZ7CpOgoMzdtZyR+/GLGnTaSzqZCiM+
Ca5HPiSzKB9YmTlOR94Na2zcVrP/IL/2ESvMiKjb5S2Mnuv5DzxNe/ZCvAnQ
C6AVHfqM/zXrZhZqBBM2+dG9iZWrzAElBI7LITnxYrnRmZKi0cXISaslB6XN
4q64kfAknoMBlV10AUH/ou6H4wbZLbhfZCSLklLTrpwDRJClVt5tvTOwTmi4
R4njiVNzSd5mb4Ra7y62m64CerBcTYGoO0bi3KjwZMfFaFQtVcD5gFezPE9M
tW2JDik6azzvoL46mFr3/ughZqNtaIcuWG8aO50swVlfxeYB1tO9npEcyvEp
vhtXelTMgXdiylz1kUGGCC4tgpAiyTV+09bHzHrRGRvw7oGa1YUoRRhq+fiC
T4iEMQX/atn3GeIIBA60VR2A8JTN5UftOGlkci1/Ta8uPlixq1YK3PpHRV4i
HRKXmmOf2eo/HzbOI2Z1o5hrQosTZohkoxoIEw7PODPBAak8UbTmcLXwZxXp
VOAcVQHyP8NuIVnTkK/BD+P8p1qeR+JL9F6byVLjt6KXcxRgaFHNXoGVP8b0
4GgfYzMF+o5cpZ2TYGg8ntnOOh45mMLbrA+c5kai5Bn4ISwLwPugVNkwq7QE
V8PbhmEJ0gK9Nf0pTk3M3ZAuKfSCl1lbzdu0CW0/4quuox8TEa180pHo3+Np
t17V8ITY67K1yk6lx9N10LIc8+fUafuQnOy7TzapkQEtzaEAD5uPr4TX8AfG
PRmwA4B/BwgpGbYbPwBuF10igZtpgXkxTsmJ/E9SeAhi1+J3byf0mU8b1jBc
WbMuXfunHatKA1RWDpYKlQB40rxAERXWV2/v69smnrW3au0ONamTHdW41/l1
fv0W56wXQpt53kQO7uKxSVd6tBPUv8v1NBPhBDmIIqnoiX4VTsduPo7tJbon
HYvyQgl0bxEtar2I3FlhseuTBDvj7wtFXiBTaj/4+MZIl2J9hIvN4+As+89S
WnbQXQRgP8fMn6SYcRhb+wfyPw5V1ApCIPrrCBDNGOI5wXQCYcVfNt6TpzJP
rk999/MDNMSzHJa2muslw7Nvr6RtlKiao2WEto9O2H0bk2F5dZN7nz0dzYXq
claaljPUBZsLQUVjp9CyVA4DkIA6E6oxWOR2HwfChSr/VhpRK8R5NvXXHrNV
90J90l4tFjttXYl/bhZn5l4DtnXaaih5ibBkzVCfYeS6l7siTG4UyQ8pCES+
WBhqVeldI/+ydl9KjE94n3N/8zpRYyMRDef90MrqOgchnd7NSle5APJp6bZM
ez8yiqMHTzugb8IkJS2w3XqpQoIKpCtwCy+6n0j4lSw2lRfTDpmDZc+XB1Lj
R0xp6XVsTZupStRZ2Pzew4xtJjV7CZzwTlOmc0uHYi1/9tE4hlIP3YSCJqhD
dHdS+sTFtjf5Uf0RGcjYKveNRD/kq9G1F5OjrrPGrsWZo0VnWX8qhgVCD6s6
xTqv1Y2NfVF5q0uUbtKqwVS9gfPamqimctpfYlOH8vgl5YINVLqE9dSyw05f
QPPLzojiKfcycphwEw3a1MapPkwRwIwcG4h8eqnlROtYkY9zUu7OqM90VhJ0
q2Kms9/IP6qp7Mi6+hpyZc+GTNDrn6oDCd3vTpkrKv/TDvGN2gnhGNyuw67T
dom0ufcVmYgm8vxoPV9k0gf35XsPM4FjbNSSuCKK4ZucfTdVIWxc50XrDI5l
NSrsg1A631l4SJpiGmuzp5hkhvjw5aJsNwl0rrF01E+iYQCXNL6x1+Xa/4Z1
1MTuDjN8Tz806OPpqnw2HzmLU6S8AfZW6WxKcDL84Nc9N0vwWF4hfKMvnPxb
tazsR1irJWvQyz3bzmtWyYq5Iuu78dNo14BEP8i8gPVhVoLz3LxjYHdmk0aA
mufpr12MMO3R9QRcjO5PovlU9X3JjeWrZKUIBEM8M7xo8w9OzNC/ysguHBSk
bb95zQsO6xHXroTbCLDvYl8mDVdANgVlXx7+eGDunAPjQqum1wheC4474quM
6B1syHhwjYoiw4zG7omFRgSzxdhOd2+NkyILrAPfeB1ADdbxio1SJ7dfi64F
jisZNENBsAwMcM77fLrUv4KvzyZF/ZxOrU7aSjcIaeaP9TKfP6mqPGluOlLL
jqKCTbUvBtS+Ob/fC/+0vgJexEMEDDNpZRYoQLiF8ifodqRlISXEJxXoY2QV
WjUIBw61F+/Nf7f/DoAXGAVW5Rqjs8L6UlwZxYjrt6h6XIzuosUObcXPHfQS
C9wA/yubEFFUFnm/Qt9febubHcOe+ImEV02d3qGVQUdyX1eF78cS9qa0cq/h
NlJ0o/XRZkXvFvHxK2H1pBjtmdvkDAtY/o91FsE40ozTfVRKdwXmjvg0MwLA
3GfMbXK0a8Bbafzpy7ZEBN47+YHP/PpNFfiYV6lj/RpdNO5Sm6SRQ7AiBy07
ark5P9aoiC0KgSCXi0DUBWJkh9jYV8sULpDom9Elm7Bs3tgFBVNmXnroMi8S
wC2ekV4fN0WRsfqX35lBLi2ftUdRdQ7kaEQSaVcmkr71ZtisK+eUy+tsjyVJ
b0THJrkwWBT/MB4Ato2ID5BfDIKaUMT6afpmAQ4YeXSX2FWtjJjMkrE5bbKA
2dPtRZtLQrfA3U0Id9X59q5yOkEwx4zb9ccj1WJTN77sfn/nLDk9HpBSKcAX
oLHdFASHtCpBYyLLnXbpnFAyK3Z/4Gqya7rnOO1rAI63D9ByEM9ycCa7OOHL
f7NqaFXXVFH/sp1D21b8g0mw6ABAMEvAX1Bdh64YxZjejDLN1y1J3Zj0SH2Y
/xQVc0prLO5ineM3iVzAD7/ULQmO9BZN5MxxXpsMAObiP+iifAVp6fE2sV5a
Tm62o7+jpPsEkk3OKrNAxITLpCgU3/tA6mcAawBq4vwakYN4sXKE53V7ZOTw
ErhXr8Nay0s1t5Q5ulLT8QGRIoaj6NiYKVlQy3PLLac64mTa0DA51ev0CN0c
hhmQfoLh4CuezH+FynwK8FqUxvWxs2drtwqrt5iUhX/DeRaFXABLzE0IzJ47
dch2sIOgvFtGqByk2P+duTFgEW+vbe65zXB52B/ARzKv6Cz32cvDh4LNQozq
plo/qZqdmKHFSHrDsyzVCbGxCDEIsRvjPNNovlsx8sfxGsiY/KFIyYy77B8E
XpVfLUPuASdgu8BmeJWdZhvdFVNt90NlJstXWdnAgSZ2loxG7GJJ0GYUWYIt
7ce3LZhiUKz9eCpwBXDwhOLjejLo7/Tfl6Vo+iuZ2aJLKQPmLABzypCyIXXI
1W8Bm+Rj0m7wl/vL1czqR90M/BnKdIzGo1GmnYfOzMT5Hq53atdM9t0wWeUK
/N5GPPsKjiMqHvnYVMmM6lIbuXQ+9DDk07B3h3H8tFu0TMOvNdRSlu2sANCO
racXeExrvrEL7/z718DNr73oWMitaQM/ouSvLx3hJeXdd4ooZWZzIRgt/Jgh
tlVfsPzaOvAPUHqA4iJJchBtJ7PhXCYcVaiBBMY1spd4JP/cJYnHP68mf/jA
lfVlCqZYItcjVYN4e909TtmeKcAcDlFNMHU16lKRliGPT8L7kkoJ+5AsUKIO
mZaYX69OEHyPxHk4QCNBF4MRlWD3tvP73wnT1vB7AcJpG4hESPfe0l2wivLZ
EsI9+uU5kQe7jXx6/hRei3sH9VlzMlOZfl3FCBNQXxTDsOfVD2NrjUMxzTK2
HC/SmrUhz31CzJdLSsLxkKNbOY0IbH8I2HO2VUWRH9R5qz/6jIOCOxAVR2By
VCEgGljchbr/TnI0W/znKdtzw60Van8e22FjmTNmZ2f4nOfmOz/yGmybc7tW
XpdMEmsUPfx8ItvC7aGu2OXlRIF6Vdm9/VUcqXYIOS5XZA/l2mYHmdQ5RmP5
OWzHTSRxuft6XaUq/kv1hNJrDtYwyzSyiaXw2Xll9AhK22agedgMTfJMrEbD
Dfr/BI6RmFQDCJnrNWHfpCqeneru4vtZNtUFEea0Zgi0W9X0IVdmavTLV1YI
nOwnNgbFxPsLIao+ad5Ss4SKf8cygsdiwyloArAb/drFQYHyfBjxspapHqbw
AnDCvOGPOO+abi3UHeqSFu/+LCiyUYNbBXE71qH7rdNKlZw7/bfMvZ8tg+0G
os74+rU6l+5V6CrJwYjS065FADNaHus2rYc2lNaDiwNhz/POZxE6rQO/tc7W
wLIgSthMuIDCHK3/IcLAiRQ4zSkWnphC2KVJ5+FQ4ZTsU5+RKxsDoIurRdVR
NRdAhtn0qHsfqq1Cc8OwPiS1P4W0HuTkKvpBMqm3KvIBAaysyiNBw8A9HwAq
WUw+HS5xAqVtzGVxj2nXRZ4dpn5yDHZQyowuohHjaKHRaVKWJLHIGPzWd0Ux
YY67tkrNd5gXuHVayvs+XMyLt3UK5hb4PHc4SoEEE/5IusPpwCNZFVMiCrXx
rImWm29iU2/kYap6JNOrqigWivxJERWlxH/Wj4oC0A7+CMoFhr0sLnAqeUBw
iBY0cP79Tastj/h6jiND/lnVAvwoN8ATZ796sqh8r2Q+bSV44V6egjp909uT
cFO9GIiEko7oAXBl/QeNOQwC9NDW1uF0E8RITuWFWMIBC7Tu9ly8jwoDJWdW
7o6KAFBaScdQhAr2X5LQmIm/VY1UXDa99hn4WQlhjA5ETC2KkNrG4gvBa6iT
txzNWKqvbPiTXf74yKfaOECJJN1jdyccBgrogod1VbjqiU/a2fJcHk62Jd/X
GN6kf4vI6a4NoPoi1ThD4xe9GmFjZH4BIjm+9it0hF4Jema1pR0qAuUzd4oi
O/CgxCB/HWjaRINw7wfdhVqKRagqNtzL2jNdJQFou40nd9An6zwHHibnfO/n
D6EHnP6wSbU7PjZHRT35YSWnv/T128iSQWCMFQAyE7BoibqH4oqGNOVUmsCv
bL2zeuy+HMGKhM0XmF1gztP7W4qIaB/dpUPOUnqG0tEB93N7dHeoTlrwOQZU
emRC4zF8r1wP6VEHjZewoA27FO9aykHShSPhQKSkAeEVNLrxAysjTiqfsTr9
th6j1wKxd8XYA9PxWnNUaACHIFy6Of2TByLJj0A3oiDaYrgN6tTRnBbPXpVX
vgcbx9r/hFxsnAp5da/QJVVbNAApmdSGBEFKqLQI5XK0NehuM8ExsCRUeG4p
/sBeMIt/uCKJoESIN9jdb8VHQih0zJGyQ8rWzv485dsjf+mz5G2yK12kRtgN
ObVBoxli+7ph1HuxUbiJ9ibtrPl3aFoApRmsHpVJ3Ierhq9+OlbbjPDRxCIo
Qx1RsQ0Owe0KXptrcST4swBo/hiTcDT4UtgqUBuge099hxRaxqgP9TTS6AZd
BRuiHjF0ZxzyWagTaGIaYaBo5NKFH8dTqIF4IXpS84FMzG6TLpDD2vA55AH+
sOJmdQIxa/h+UyDbXm3G03MQgwBJ4CU4Dby687/HHS9DHxlRL4of6xOSigYa
uiEIb408tvHYX693KyUCwzxq9KAIzKKZCvaVW228CieiTCfF1fXbVV91x7dk
iSNB0rOW13/MP/91vBi6sCVoSIRg1KziPeJBbi++LuCfVO6RXMZoldfxJ+1J
xOUKK405PObk9o8jdhKAK3nU5zFNfic4le6uZgKm+LGjSJ9A9/ssI6ZizvZp
qnsCMYj+aE26TaLKAQzAlAQOFCFwEsujOAVHLfOjWO+m3EoQ2Bdl6z3OuUgL
Py4/lakyMOcQr2ZSZ2gfHFYr82lhdANTFOA2S+ssR/zEFwPHHZ4lPmHzPxuH
Oy8qQCuJTRCXfzLIzzHy3RJTa+6N1iOGhWIqTA9MoOIAOASUuJD2Oa+2RntE
WHrW3giSkxUPy8YXDSSh1DEWO/nC5a4VurAVARO9VPnFho8N0SxOiKIFzoWO
+DnepCGSC3cV7vhaV9uJSeqdDwJxOl7/EKHkTq7sqbDmxbSuho8XX2lFzjMz
zP/xgNBRQUJzqq7982wBhI7r0Ap9TRA2mDPjhxA8HcBTan/A5sNmBLo6PtuS
X45tnZG5gwVVm2fn568nNUEhPKock03RS9mc+n97NBLEmaspF5vE9IfHdBnb
BgtCH8zBlQ9zjQc1H0KXMPbh1vCFfhp0GnYPr7grquc1sBMCRljoFTrRuPkG
aOP7aESXI6mGwu+E91YdWublFfE989bLLvW0EQnFs97vcc8D7f3PqcJphVeJ
1xDz1yArVEa4ObJFSxTiBmOzspInSBloJHO7ewZPuRk52C8Yg4/UimMKCkDw
wrTAXZKkq6CLnLq3cI6UXRBnjN+SqThYmWVDHtFWw0N0T6rlitpR4L61KbhS
SG4Efu/4wi/XNgVjB48nnnJy5DCuRZThJO0VMEa5/MU99xTebJM4rztbUlNQ
7sQpc8eYMndeb7YJi9oZ7UJP6dEsa3ufphp9POZAOgUDmweC0JA4FNj7OH7m
L33J7sOq1J19Tjb28S8JiZ9nQhDSwJNeV2Wj4u2o+nImjCBQCQ0tSP56TG5a
Ss4neSlILZMVTwKfv81FNfDRyWqtpP4A3CBhGc0isSmK+vgP93x6JqKLE2mo
4DHVjkQ+KDOV8AbXnvwNtjUeQLeDvGD73Az8NsNCAN54Li78iDUbUwkl6RM3
m+lisPprmd61r2fkA3/+cwtnb9ztG+uf0rqZwZDjRx5OR12OAnqtKez3HUOc
fSY7sqcMzRAywIMiu6+pE06nmn6o1OpbPomI1VXZhq9mjuthzWRw4SE/5IXg
mMeGZtuzmt0ACUNMmMorGhL0Cd4ecuLmmuM6WuLbKRD9Tc081kR7rVPA6/Kc
1ufehDzhEfvWMpT/Rb2pL3ZIG2a3Y36fipiGsyctyGmHMbSJXDDIjMR1S/fJ
awJOYyazYaNglCwgwzVOXcNC9clgsvzXmmzFYPjJuc7SUg7/PJVXs4pKpEMs
927iolDBDsXzlM0NngX2GRtzUIMbz8dqrHxRDWEzmRvO0QES5fiGo5+9rb/9
kCDHsayUg7VHygIWfdOM4QB/TTZeNKh29BcY2EUK8rBDmkq3OaO/y/2dz4cL
zw3hb+aMwbUbIPktPVZJRgEfuNrFXcwXC++x1qiyShFa6rsg0abBdOc5n4Hv
Er77WyUvyxZ5h7qDwdpHFxpNuebrbRo4lGb9Ct9FAjFK7cqz5RBW2baDpdin
gWLDOxgBbjSppw18hQMMkIIK7hJ+2J1dVYIva3I4BxAIR4p/WvqKs1m56zci
+j8gKPMSngC4VVV7lDbjMoNVs/k2YKMLX2A4ZPZ7anf9VgvTW6XS+K4r2rf/
MeHVirnae5FnAyGYIUWW0bQI3Xfcv9W9ZSN3EypgKF91qP6QF4HaXRAwJiXE
e4lqRRtfY4/a7D/+1XT/wqIMGgu/4m0kmed9subH3MwDQj2Pu6NoVuTtIcl/
aFe7W0hnqdWN0+Z8DVcFZOUPPibMl5cEHu8vhUljAliAYyHpnrkymjxadIRD
fnKMVCqPnDuklMHvQZJ2Ty0MpRFJYmSwvs5iaq3sZ5drMFQDpC1g5mwsjPBe
eQ+Be/ndKOXL09FuyFQpShyebYu22Z87bjyi609Uxo/PeeCUwCThQEJ35XSa
zMDAPD7bQFDiQLN5YNIS1cOuw7/Vrs84HZFItohJ2XqfGFRmx/3v4p+BCgjQ
tahfmff9uminPZzouvW8JIVxPPOrCKPemTgdDtcSIkOHdvNpguDoI6ZMaM/8
rlou4xdQy26rqi+4zSdzMt+P+uTES8x5acdDSSAeDJIetGL4amLvrYZ3+Cu7
hsL2yAfXH53HQW7od9lRHs5V4GVN03AsrJHLvlm9aYbzq9uza4t3I2biM2EM
qPMWBQhWCc9T+XkjM7s0XdJaJSekPuQow6DH1+laW+DSRRDlzasqsS2Fy7g4
P32pYKo3RtRfjPXzftzc3zojOjHJUdp6707HfnB36KgqZj5kQcck2hRu5QDJ
MwR05Qp2I33gVowpxocx/cwNJhi/50tgQBVa+uLgeljZrLH4SDZ7cNDthy4M
kqb/l3Y394spvvRTtjv9R7RVnx3IDr0laONE3v5NaYCiaCrid21B07N6wYF0
c/nvEJxuHh650REnNffrx7mfw6dxR+bYLZ0i451S8R93+cLGkRJmwSI8a6Rr
j8cke8r56jxk+RFQhudzabyDFEnfu+LVwFL/S3hFC1ahKTf1IO4UfwjYlhUD
TjW0XHKZAeqxhipbhycxUJFnPW3nPvkZFNbe1JvOhTho6eds4GoYS8IIEHEG
LR6E0ot/FWxOwtqFtW6A/4NlvVXWE20+8hYiaQsG1U4tV1lOsL/mU+5JDe4J
ReXJt3qXPpgF7ZGrz0CUPqbrgKc4oG18NEjnlEGQ1qp0ds+Bapl8YZNFWhMM
LO/P1fsOQZj52GKoRI1/Cjc3pf1jlFcCcn+OVNsRy+e8gn3MUdKbuoNlxedy
oFX4Bx+qD2A/+KGH7R+vsG5G8durZi7uviDPGkj5dbETEwBn58JsTfqHOECb
RjDg++SLDC3UBgxS7uxT0B3HGd2jieYg9nNRDUToy2GAV983XbLrk/XeMUV2
ssXdaT9uV6J2oISH60ps/tCKsTx4P2OxLBwDNLQR6dbDurETUgWIyl7f9Vfk
i3fCTz2dXI0cHr6TvxXQxNrSsmx7ryl7i02eyTJvef1y/Bp6hPhlLleqJ1Sb
CxWqCnk6mwgcaYnyjKsBkD/CU+9vHTQ7oa1hPL5HPddWQDvu9xg16j/gLngv
ohPU0Hk65L3LiBQtWs6C6eui8tdrr8N1OujFNssBOm7eVvLsC0c2FfK2RTC5
EfKrT6hk20rh0svEOMj5z631vdd9VfRrLOFjwemTyfNsMaas1NYSb7a7FlQv
D1D3skrQYmol3CJoj+bJ3418MC/u/04EODEa+rQilI30h5d8jEehkaU3nM9X
MOcJOg4mOGagmxv2UPHO4ENsSN/m//arbjTXSpmeplY+1h8Mu2v+6AlSbiLY
g2MoNfeslC7jlZT7kyFea3ToYGvWQvqcPi9p2Lb4BdLmUagLa36LaGhcKfoz
Ovwg6erAbJpWOQKK1SDbJxEWpMy8N5ERf4gqkS+9Nr8hHy4dhjVPMWebR1Jb
Ye+VrSLiM/JJ/PdzR4auEH8CbbGa3yz3M6UPDta/YJiGYb5kOIZ6iVqFdstG
gHrlpVcYwKj3MNAx3id3P5IJWvICJW2nkdFH4c3rwrvD4TqkwZLHpxb0KMwP
C7n16NGBMUP8EPz+jafzgw+u4ZwtAObbn3K5xVnfXeDiOwtLETQeyyTOMpE7
EqGfy6+Cw+oQ8bSc+9gdNARK0KlY5c6S0AUZpF9qhmDFOYsHBhlZyysl6xjn
X1TuOMm8JEaGkh2I6/8vcwrzykBOq+I4alk6aMcjp6iHAZGkTr1JCG788Akn
bFqitr8NbkmdwEDEQuS9sqgeK7oue9xFQ85nNg/rBFH5I9TH2kdr4BdCdj5K
6VZT+BREeZvBNXeC6P8KYnGhsh99U4quusOgYrleSoKVODmaf1atU/Qapskq
KQRXhQdVVpqPraxyswPfVK5CTY0mJ2PFe6gYonKU5unXPLDeJ4MUPp1DtuvN
IK6Njz5/ebWsQ5HNt/OdXg6yrb6ElVfZuIvcLp8+sAecRlujXw2XRWUuPvN3
ufT2rZjlzh2huXom0WMQRyEPKTscIfkW0xY7nkqrGXBGQ9v6Fo925DktfEba
/ZXgqCE7IcibvA0vbquzvTGxDIKU/AV+SpOCtsCJnXEFhw16n0tdsUOjcgCN
k3Z+5ZFDnCh11Dv1qqlVSl+t0vARb6U+fh4m5kIBAvctqDAcS+b31rrDJTm7
XhvQesSS2fhS4akqI/HpJt3u9UAZ7DeNuWMuM4DPm2i3/nb0qTqEiKMjm5qN
U2sj81Z7zIa1t92V6fcPeuQ0bJCuCKoWAWydoaK6PgJgSdD1vSbuQDENU7IA
0Rx3GXKi7B8ygSMvwDojzFjtFCjXwnpwTrXQNNclDCE4BrBMDShh4GZ29f/k
O9o+VaOtbTs4/QB0/DaxzLdn855cL5V64khJLYGbZSiQsIUAB6jrew06y0z6
l9bo/rC5zGf4PnrUQPHUxeTGu6yfbYnmKz59NDrG7doNu5ubo1xEe1+Dxzqc
gACx7IGxp+uJs2eJGvJmf3De5XJHPRskaQuJA3/nPlepDM277BDQ1t6P8R7q
f7q6dCEtqICtVKhkgM7pspg7Gd+X7VrXtNOdlggbnl9l9IrgTXFr21hDolgw
Cq82NNSvwWVDRE5sKEwJdKJuEEVs+HfmkBBhboXmLXJDQkBNGMTVY/Il1ai5
/lbRhv2i5dofMetFJt4ZdFEZYt/SM6SMVt+hikcmlS3/s86Ew+GWTtcVPneb
mrZRAHeldRV/94ohEAFQO5YkozA8RmN32sdXVM4iWwMFYOgpdUl/jnnhB4/E
wJfjhFAxMoMUg1ZrwnOZmBB7Saua5CUN/3ee7M0FzpZaJ5a9Fo0g4rdzDlW4
feDXAsjr5AYEXVr2s+rbPNjiVggCPmYp3HbKZeKsZ/7NxmQ71ZYi4ZNgICTb
o80sVksj3uzBtsnlPoDVMj9CuV0qS7x057Oe0icd2aDUtCmf00jipgACyLB8
SpR/tnS/wnXE8w4JjYw1HPkN9RoCccP9/oju/7bDihVfH/wFwQdHoSM3z565
umxN7zlRB1C7ckUz0Zxb5uIZsFEUUu2HMwQelhn4mHpVRC+x4LgYSGq2mJX8
vmhAQj1Zkxfi3oJrRvA2ITmmQic6yVUtCmOv2Ns86k3HVp86ldyuiAmVrsLW
5e+bvpXYOcxL1V1SxOdP1XtKycVfomkcLw15mxY/6rW9JTsevXSm9/e3gITS
uxMFyhrl09ytR9BqUfBmVN7BZ6YewKHJ21C0R6dIyJv6f+PDP2DNz2ZSGiDc
fmgHTXYfBaigB8bX4sI67G/clavNvIeeVj1jeaeexsT75E6Ieoi9AyZRWwaX
g4jkMq9HOyTV8wne7qzvOlJN+r1tWXDYDc4qk1oo0zFtcc0lxhUpuO2uDU4M
K+dqEfddQR1+sHzG4wCbReFYtrTvqfQDB9ea344JOZHchwLuc5+pnwRuEFnR
7wE1VHXOmoye8FL6z7VQ/0sjF0vWSDFOlYftdYGkgT1/ZYohNtjQMUc5pAk1
rZN/ekSZkr9yy3SJtLyV/ESbmPtToEzy1BhBCXPsOO417MJt4csOPWA+NcxT
ak442Uyc5nngNTmIRsBVRMFKJbA8eX9SB5lo506iQRTzRprDcVYbls8QUlfK
Aj2bG2Eir/TnQ6DnHmdl8cBQJPo7WhKYgvO179NiYGCy+0ZoYKSny4ELocgg
0T8VS4e7JXJRG0vaedxCby0Vm8HXaahMozF+/WOzbMG4LrIj3j2/9DCx4Kq2
HUP98Se1VOM9QSmiuNaEWgRbKv7sEWgPgCjKQFVvIGv8omQtPBJwrwpnMJtT
HXGi3xLrYoWXiXwr6PCg4Vrr8q/E/B3ppoDA7/EOpmobUST7B/tJ887Y5yfN
ZI5jdBxO1nQSjY48m4jjoLPnnO4z+pUMaFDhXViPWIrol074Nc5ICksxoyv+
LnO+MB2RRD1++ins5JbHMLi8UcQ1HbeoPCmDxgs8bNi9LsevyQ9NUDAI2ES/
fYaZ89sM0Moe1QF76zpNIadH5r37UUfb/By6yChuc1ZQfHJqLGKp/8jFeNY8
noo1kPFGkMo1nSH9udBXsBKmNo4gpeDT5NZ4et8ZrLIpyObKnFcwyZC7Cc6M
a1aUomH2nVJM8maDH16O3AIi+zRrcDgahtpUeocxQmuV44fIZKjraU74MgOW
AY97QpKXqJjBmgRiGJxcVJcANYLkXGZA9Rb7qFMzubWCpKCiH1ObOroFbJCe
JPO0GthYWL9PD33961Dr/vHTjnGyJeEzoXYUTS1wGGmsegxwX01AaOrKjSKV
ejL/iQ06HuXbfMN9dwfGMxAR9i1X8hGAqwmyiN58Zpq0XDM7MZl/q8IivP+o
DfyA6dD9lJmuGpqCUg6Lq0210/WnFM/dKZ2bcHRF6krMcljBWNJam54x3FrD
pcrJqZxN0pzZwZaMmqjZ/K7SJnstpW/unizGOanMv4z4Xhmk1pJlnvVuQxZ+
sOgYrLW2qHFr1prDhwCX8GoIAb/Y0zxgeYl1i33KA6WSON1bG468qzV+P0u5
bzgqy60AMM26OIjkBfU8tabJN3XCoxx4mTa+/2k0WUWX3NDWfrGCB/Wrfdjx
glJvu+sZkufNvMJZNh1LJ4Cp+rCjHyALxw2rHdu0vkenr4DCkJcuOWMA4uuS
0EuIKyfJkmolDy8kWGf3bl+sV3xINOwvLpJKyx/VWV212YiOYCY8W6DO4oED
Dwz55vqabg3+RLd7PyHDpndgCgCf8NQt8TqlZz2hqbPbnrlKNBCW+IdslCUt
g7EYt2mALXg23VldQIIZ2gAqJFk3hll9TMEuFvHMUz3Xkh/3PPqsajJBXh5z
ustfbig0FB7NUnw4NfQ0NRo3PA0dYBxGJ17YULKuWrcBZqFPdW45hxd2MFfD
HCN/3ANgRkAGNI323hfVM9w/RFGx1RsgnK9KIxQH9Xw8mInKiRI1Jd3IBqM9
295YaE3kzS8oLkR4OIldVAsC4miai/IXHRYHTvgZwV2pDwRuLF4jLBKjbI54
Yi+7QzHeF+B8WaC65Z3+E0r8MM+XGG+ymZfOZlnFkyEJ6zZNwykOEqgoM0Kq
6Oht5n9KekkXvpBrQJtM4BmnPvwwzgf89kf43KDl3DbHQDEzW22edGUVy32n
KOa4MQoou2EDB5Qu8194uJEc/BqrlsI1LmqKrzVRY019iyxtx7qCXQenfgkK
4xsZM3jG73ZbUmR1YgcpCL4LdsSVpCfdxOkntz4JHToxl79kAWi4PBMadxLL
ojHDZv7d8IoPnpSftC36mk4kj6WGGo0VQZ1Jb6WqrfVGZrboggcY2NGybhXj
A1Z9TVekjqdVDp5AlIl37OvG+GKB9nOaYYF4AfwQ6tZfBaovBPM/bs1wvIFx
w0ICs++wvhXXhcDyk1maTMABuUOkv0Okpx2M2X4pRoRi1XGhYOrmXsKEYrqj
Tvy6Jr6lGZ15HT+V3hLRGwRrV6bll+BfUcN0kWdmVwmKqiwJvU1p5reXisSX
m9pclCwpLqM3BpI+qI37dRkSny4EvAYcE2Jwk+OMwn/EJnTKyg0/1BWr2jLU
A7aTXLXQCPc8tZvyM2IT8y1KtEKLyu7PAi6XeKnU7KIhFQ1R64NMg25vhx80
CJnAGuMMXOd5NSRbbSGogLy9nlp6g45nL1Yx/CLtFsKoAPjcxVmpxU0x6OD7
kTDsCW7QxfsLf3EaAG0LMHi2w8HidENSfu7B3+PNSL3CgZOdt4ktYvKwx8iJ
nmI+VHondbdY3YXWrmxXMM/P2aTdDrbz9mNL6UAqKQHBCYrrCK+ptCFqH9Uj
cblQXuuDdUq+voikH/HK2+FesL3W1TdfI0lGZFlD6RKUgSnVDuK3a1Cc7TWn
WquSoO/dlYYqg6mBckUzt0zJ2rNyqiJ/jMFG4TmAJggVWvFIA5JuLz6U7uWu
Ov4CrKfDWBUFQHAhNie01vRDWg8g0hHPsossI9a+NQfxPthgkF7F1FHws0hM
OcX70535twqJuofrIqOft279hf1aGHPBNhbKC2pS85z5hEG9SvJTTqvSPyYF
Etbx4zSdEqSmz8ayQe2ERfbHf9psHnts7ubc7/H3RlKQfKzxHe05Bbnbd0EP
GvVQSHHTC+NzqpmE6OjZsvRryW9t/4bHDfoPCGijJqSwwWdunzzZ+n1Z1dKs
G7MnYdPM1bJp2FYtuxKEhDb3Y9nUd6j4MhreaxbMO3fFz3Sz4hFEwWRTjSF4
EiSMkMNmDvW8cXJ2EP6O3ykE/9GxNccuLkJn8zB3DBYQWT94y6Ei/YpAwsqN
V9+1xFK3mETlwkL26KZkWQJKV3AiMiZvObMR8uURlaZKk1YHtc4faD8TInAb
pqfjXKjlPGLUsS9h0tTrrPgXc88SjsTQIqtDq+MbdHOqTGupHX58NCFU8WoJ
ty/LdDenyS7ggz5tk2XvYlMGOssxG3vdaye1IOKB4CkUxcLpsFKG7VFkERDl
YGXJZXQW/yjPu3hb0VXe92xlP80yTH5YC/MowraobCAbDWpT9ZM4uXyZM/Da
XamZJYarykyOer4JQ23b1/MoDQzy7pkWBFPhEvVE3bAyV4ubkmlxrvqi4mYu
nV+gtMqqmXoEamvXYg5P7tBisrJ6TUdM+fchqn1gwkAP8vwQhXRRInZS4VlR
sKmCweFvwWvovWmmSAFEPetDqQxJYF9b9thRlG53gRkTF4r4b5Ad1ZgZJp6a
FRGeYOcl3T1zS1JF2rntKsGyF+xh/4Bq7pHttvf9g8bQ6xCt43p0GC4nR12H
tDO+4CqaTJ26ANWFPc5NfcPi5JQeYnpbweLEGLbzRL/iOtfNBhzoSZJwkElI
x2PboXDQ9xMphYktb9k0qMToqLkXSmMwPrqaDuJB00xd0VGBE0lVoGn4cYlw
qLvURhD5CE2B71wLvpt/eJyQbu6A7jeN8cqsI0u5mOuFl4ea/W8qCeD9NxHm
K4yZLudpuF7rYU9PMV5wIhMB7lUa2qNrgrYb11emUJD7ExuwRdmHkKoKcgcy
XbcTlN9v9a4y8M66CfeYdQDlQQpMJXsCNmErA0eGHSPWQOYVnKjYy+mW0Pb5
nCDm+gYhwt2crJWlVdVdSVyPiXTNBwkt8MvaI9wBK4L3D4P2y4dFk+v9YHgX
h8dJyyjZ3WrXZ47B+92sVhFa1/14Jqh+dnMNv4GLauu8O4BZTv8lJusesQCJ
TyS9K5mBHIQQpF/rWq3wtNDRnIcBnkkDXS9uarI+XwBQFH/Px0eaFqs7Xdcf
ojdKokNBAQ4JjjqVBI8ZoCbqb86Xex0Nv1UzcmWYMv3dBQfRPXZhhxLPipDf
zb17mCZqo5ZX+Ex/ZmbiJUaircTttJaI6thjJqyB7wi1O0IjOgaGtDqmNprN
ZFztO7Dg9gX2LVkrqtKNjtNcxRez3vO9CSAa0ulnNQM4FDDAjq0SPs9P8SRP
tX8wORLNekOGo/NWP6lle5T2FD4dG5nL9hNAKU5RLTzbBVBAZWZvqX3ZvfVj
uTWqrQJxL7SfcV2nUSiCI+oRrvmqsC9FdPIMiTg4/8qYfQZA/AWUI8Yi0Fu0
of51LkNqMqU+UdfaHYvRMGP2SlXB548JdaIxlVgtgp3f2JWDZKkWSGfDOyan
4XgskgBgGN/xLT4kJrGWwxH6e/jTvKBe7ZkXAIqtpX3TBuvy1G6y1dka+hUB
mdpDgIbTBWbqahA2n/JAkLM7J42snRO2BJHoU2tlowCsaBMCD/6PCNo6SzZU
abU69hzyNUjwmWobgCSHZQpXySMcAy6OxAL2WOStNWBVLisJaCQN1azf3cr1
rcgCUewKIAG3LdJ7LdrAExq0c/aNMBf2vjP0qV/HFtwbQ26i6OcfiTzH/AgP
tg8zYpWhnIxITneiFgsGWpSe/kZQr0A9F/+OkYaOl2b2ybfNOU8r/U4wplw/
Ho3KoKvJnKo+slh006loe7/yfWLsd5a8mvxen7aVTc4fo4twhfTQkqemjzLn
6jOMoSgumNd3FR5/9kHV2Ckm5XcCHwakpJ7c7vXkjoplggg5Vvn07JunnfoQ
pmYJQWI/PGwSyxjD/jCTkZo23YdEk+Q79cQByWvMlLZHIYzfmNgKfn3HyaX6
jLs9Ai9bO54axGPvFZJbSMhaasX6BZNFouh8i3Z6ZOw1BkF2khsgstStZ2DO
wIWS6ifmWKlWvdTTSC/DWrpxCrS/vlW6I+LhfTH+PUZZqMNCObLc0W+HwRGn
esbvmXzGgivdP9CTipmgLXxFGwtxTSlZ0s6TWW2L/JOUWp/zNCjUw4t6mi9F
ECbbdk4NZvJGyAVyueYjtcRoN1eT9X5uTJi9PWbFjpjhLHIBxt65ivfOn022
HMp4R/iZ0J954P5395sgn+H6Ri3GLL8Aqk8Mclt8e9lQ7PyOVNmXFpi8/LSf
qwRGdKYQx488cvkVpcZE4NSZ/zk3pxv8ZYq+EV4FSkajymJNfV4Hozd1N9A7
iC1pp8tnL8oGkI5Mg+4dVTyGq1n8nSHzGqgv6v2yr8S5A+Q1juhhEMM+t13I
XFk3/RiA0kkCXwaLvrxqJ36p+JjHRuh/MIgGpS/7N8qP8rCNFNu7b6couAwg
LSRRB7n7HZwDwScRSurF3ARC9fmQsv3CsOohIIhraaTw2F0AS3PqldCufxCc
MMW1Us3NReX1bSIJQn/2cP+DHdW5QYg8ZOx5uuhPqsS9FK++346Afa8vsM09
TOCHmHdvYPqAOj/18YZccn7mpCQWwI23DZBKvFvq3dntjZyJ5cEh11/ii56i
z3pzX/wOqawISXjyYMfuNnyFcXWGIQFXeZf3d8whEpT+L/eGRo+cV1SzMFCY
Ss1uj6HqGvpc5mnLFFiVfhHiSJoO6MfYaqjohjpLyLIraCpzhH5xriB0DRby
0LfbNX2uWV9ptyGP2cqVE+WfIH3pt/dEg6wqK/DFSFdVluTDoCSZCXt31TXd
Zi/tagD9EgmL6wH2T5wefrcvU+XHQe7Mn5lOeMqCD9RBPaqtoQ2ploKYLby9
2kdnZjNESYooqyU1uYBBuGB7XA/8pp4RsujZEZ4YG86lpw6RoAv3Fw8jHnSD
VGrqElt+EnUgK8UrWZQkp4f7eojO7jxF6wcoTREwNe0j/um/JcWtnjm68OhT
nelynWUTog1HjU9pETZfCzZ2KdUl1uJunLL4U92aZctysbUEzU4m8H2AZ/NR
nawaLC9bz9i4GdtwiT21OkBQWN0AkTUic6tPTNBNKdxNusGaej3hKx01rRqQ
i+viCZLYUt+G5x+vTjbfv2JlmKlw/FbMC/9VyMREjf3x1vV5Ib9hUBP9ojAb
z6no9Hv0OX3lI9lE3A5+Q7Yyo1dzTmFmyuPVyoJ7m1+00reCpBcyDECkV274
B1rPO/lGYHj+Hth/XJUn767+KkOt52SKlQ5Kod1AbqoHQiMQVMb4KhlGoyBT
GK3mxpoGIqhMcTvVQr1AZcxPC0HA+zbP7WuOB1QXG19Ds3wn35nakw2JduR/
YLAtEXjzR+nBOx+C1qdAB2g+fbzXu3BDZ6eZzOV5dBSnKJbozZSzMSAqVM5c
QsrARu/j2/rEUHB9W0lFJbFTz7Ak7fvspz0MDk8tS4mU9rLhPB6jlbR8V4yU
inF5EKTyzk47RZU8FwRrC7RnhYzLpmaw7ZmfYhl+sr3rqetlpHO3IdGNNAOy
cM2ZosioWK9SNiXbGV28XJhByq97aG6IP3hhSgZLtY2558IA6H10aEOsujOy
0Y8DGW9bRn5YjtNK3W71LMT8Ihy+VH+6reXHp/JdUCdxrWWhAk+xHiM0iEB9
ZcpH3IVVi3J6Kf2+i6h8DeleynDw3YdPuPHttkN1AMwhX1ikm/oSB8ZZbUmP
91ciM7mb/BdDIRo9Wdx5pePNrtle7BHtpcdm2DffaeoBUH0OB9BB9JkQRxa1
/Pcq/jHeoN4KkpbZlNV9ypteN7sB45nJo1BGcGqcGYh/VbDK+/nm8gUBxmx3
2chizgkKTgzJk3rgLlXC/TBt/mdLvxMYcZxkzQqpZao9YQOBwVJaXOUfMqYU
Dq5A6qIrdTWf0YEWO/mYqTpl4WlUVfpg2dZiT+eVtDj2tppOafEP5OTTd3ej
uWpre44qSn85zPtJTM/eR5XCyG2zM+ZnVwnJAB22aZv/NxSQKAF2n/TPv0QC
+bxspn1vKTL2ahIVISduxN6febCtGykbUhRgLj4kQn88KJ6KTQNBXDV05BHB
NPbK/f9zI42pQ9G0DVD6jJagnpnvcMb1+g1iisfuPDfYaJfrXl2Y4EbQD1Z2
OfAiKF358HZnSHNaC9gJCOS7jNNR6962UfCrMlTTFLeG3/euuo+Qr7bf0gnT
z1s3nxBMZ1355FH3NaZ2b1jiitbH8dunAQ25ND2MM22f1zs2HiBkzrxgs0U6
gF0gxQ8Xf228Xz9FcCSMNQp7Eov2qMYvRvi0eEe0iAHYBr5JX4xXO3NfdBtl
mLwAK4yFCfOho0/cydSQ2admfbLyzYc22Pd7kC5bFId+mqGMFgZbh7dpKOQ9
DwjWBJbUedBAOsNu5PM85CWGbX2zRV5kIx1BRkyaV+cNqv65bN0s+mQgjzQp
jWCDs0rLkP+XqTTy6jf8v/3ZkM00YufmAtFiDcn0aCs1iU3UFqj1hfjsell2
sz1IjlCyCkM/1LHoDeCsX0V7SZDSGXQIcoYJ8F7bFqOjCGlgTa/bg76U1COJ
VYNAVJXKLl2qIh5J0SWjVR8b7RfR8r9LEcXgQy2EP8XUGzkBHRPLz4ZUwrDF
BDpByaqijFGIOmtB8US6olcTsNM5Ey8XLMX+sCk4zvldoV09yEmZ8sKQADTi
V16SE6KhcVeAwAyQVO8rStrkr3UmchRzEFVVYvvX7AUXZnBN9RRJhE6+wEC0
55HrGM1BhdABBpPB1Lpps2vLeH4V3qCE7ILMU4jA11SPmxVVf2awralcTKan
JHeVKxebKLurjvh2ezCrQHZ+VCHAECE7fUXcefd4bP8FD9n8ZmtSwYXABD96
dsOcRivKJzhW3Wmtj3APD0U4FLqS3Fk7jrFXkn3I8sgzeH6BGG2qlv1HolF/
7z0mfbq65+3vyju8PNmpnYGbw9Or71TqKSzCdxN42hyynjxa8+5l2E0GloOP
1s23OuWLXdYGK4aPCrAGd2erWzP0k03lFOn6L43Fjs5dqljG5fwjkyoa1lVW
BoymPVA0ZO2eb4dIipoMwhP7St8K5lu85rauA7sRWhFxHeLbw+dHu7Re44ug
YdIaroG/RCpMnYXUoJ7GKpHVW6GvhwtvqPORn7MIcDREFh/XGcFpzrZdevel
uO0W+/xCZhWjuVqreBRFd78y8BIAZUb4tOB9MM1JQyjv05npVUbI/MqnV14Y
Jlt/lM+NY/ZSx1Ih9p0UKAOUKXN3v/2AJvrZwD6IFFYzTNCIvpQqpYzI96ms
jGyKeSA2bLKUUmCrVX6Os10AlbIihFBd9lw6U/Exz7Te7mvZOGwjx2bFPJUi
LTCs1WPHUMe7MOyEZLjSM8UtC3m0KgF6euBvNyvGzbQWAT7S1Tc8VGVJQ2t0
GVd1Of4EZKXfLaDBUrAMjFEFU47zowpBpDJl7Y8y80h0EniIiPXBc5VjSOLc
c0OMWTUlOnYIMUNPAlJATvt+RKwlWqsz+i69KlKMP8dTUdnUj/a5RhwD+HIV
7f34SKvuUYl5Pwh6IpXH/wK6K6MN+6rz/vxWtkkF2m0/ImgJruzQLZrqvKAX
uTQrAJgZqtRwLkkTN3DdMUc2rVDzv1j0AvnVXmethkjCag8UtiL9bBOrnpfe
Cy9xmHBvexF+x+OxKu9aavS3BmVoDV4x97E8ag4jCn7ZgrIstJ6OaKBLH+3P
x2fk1RsXWOj1biMl21REiaFEXxW3sMlLLWGlBCA01mR9E3rP1PRkT680Etfo
bvP5nrWaTCTskRRT7/fzTUoHSvPsx7GS4ng7Ft3btL9HE2QIq5kcaOTWZ0Qb
PVNdYtSv7lSq0J3xUsaaBIp9BWtkOMR4vVajFFH2hvRu0/f6e0+CP6rcrrQa
uXtKonTNbqqIz8SSpZ3NXZ4BmJj9GW3cToohvuDmUmIkL9lI4C1hTFeP98+C
FGAwGEa3ey6LvK5dyV3LBg1GGiGYjeMpyxC1/+y9mKKPGmFadwHQMANu0uO+
3rrENExq+96R/jcPCKjYX308qWrVdlFXgWoxpAK6yYrD+52YfTuEb8CRYLzA
RSM282neWnda/LghxSXbEWlaU8rejv42SAENpw5ZdZ/igL/Rtp+VrBE91gkj
plRJ/WqCP2HyW+7ZtSH4dp2oEdzfz6zYlbBLGmYmK2+LJhbXTxOYywmBNuFV
GY3TaLLBPf4+uQN0kgZT0KhDgAV+Wp5VfBEH8RQKbXRi8+ldrmRvP4Eg8sWZ
m778WrOPY62ZbVSkKOt1o6kIT/SXwavewXD7s+opk+atJ6xqIAhlWUZEspIP
25tADA/iIaC5rpUjNfkO+oa7I5KROGeXKIzOxFGcuzC2J1JgObkOFlL8Moqd
DgfDZ9cp/6Ixh9Qdb1zg3NPVDwvzLJqUOIF2qBwdmqCTFe8F30RxgqzLyDqN
P+ddnqRq29HYsI6eJSt0faVVFNj4W0MKSLAhA2X0aK5jHGMBGzWhLYb3Zugj
HVJStpnR0+beUSHSEieSQlv2gtMC48bDi46oZIBlFK9fmVwW+cC8qdw8+KjC
24iThia1K2rHFTiJR26AzI6t/rZPMcwK5uGL5ps9VpByetLEoF50G7Oi4AFK
3HZmpuchtwskeYBNJD66X0rPV+CM+n7x8IIanUbEs2Ma8Yip86OqY+KDNpbs
nQH1fbff9cAQmc/qdrEm4Au7GN5ALvmqhg/EyscFqTU41v5pjIkwWEsV9v1Z
qOxdePWShSYlYFHyOd5S7BrItwyg0PVLr+MJ04z3sNslMWOcmscqAmsf2nhK
CRq16nz9RD2WtiqgGHPNgdaxpFyvYsKym2Qbl7Z2wcmXDFRi4fDe8tciMDjB
0XqABXBMI4sVsjA3aZeFSPrT6e8JUKC6mhUYXV39TP95NsaHIyu/XQAwSwhY
Q1gphePgZxsVHPF5AtiHzqAxu9RtaTMn+YRE3tsKfqBQU4696/vT8SPtWXhE
52/QjAMy0hsW53QsY5eYsstVHWF+DDom67FdK/iG6C+hiKCBVhNGaaBe6xXp
hYZ6tM1gQmebHcrnoYVJYr3K6heelww4GOIdSILII+ttOQ5NwMBVPnDI9/i5
N3dJc7b4rVjHaO0ns+TuVpAeUQ4hPJAqUmhCFiKmCLSNDDlXJnjNV25zGYbV
OePR7Szd5RYaWf0/DoFl7p587BRWDgQcd9UzTKE95Qh/s1KYaRsBzKNiksm+
hwNyA65h7ZqfgQNoXMUhI5XnYgN/l6yO0EFGt43k6PXnCd0kzF4zouBZ55oo
Vqm61xBcHIL6hcvXh09V8uHyAIH2yvb5Pdy5onUJH9rNgWgzW3RhXX2P/Zmt
r2AugXV9NfYXhyz7q7kJhiU9cWxTbQEQA7BmzT4JoLj7cMup+J245gfcRMmg
KLBKTf6OHTVi0zXvmxXUJzn2VCajdrg/YOF1rJZMAWKNvpG0JdrUZJeWbH7D
3gVw4d6JTlQxIVpspWMgvtMWSQScJgPt2+5CN10gI5D5wU5xU/TEsyLhzIK7
tqlzBL6wM9MKiVe3cSQpz5svwcAXgdARI6UEL61uKxXGB0l0+EYpDeaZ73DG
WV9FvpNhqmEKSN4Y9kEbxYL112XTvtfHuEBYyefR51cysY4FJsyrqlRPd/8J
JgHsJyXs7USkyPQXwgswXDfHKHFQaRrZzdWw/uFyojqWEyWQZ7pzhT7AsRvv
5AG1WCr7UVxSxe3D6Qa+f3OXGA41N9B3WCkDVrcuaZORQJNdemySDkmUUyZB
7+AIrfLmfGoCc6dgaiJTn8hKSUfnEwIJUT1tRcA7FnJHLPbfLGU8sfkiUcPk
3trCh4Bey2Wo7frhtKvIeZnxqn+p2zBtza0rCdetopcj8rA/ZEoElo70IKSK
EJ3ELYRy1dtLTcw2kZQ9D11PY4SB8Q9Axt/tRLDk2Heec89WKnhs+WmxSR2C
VRMSKsDf18YRXa0ZBXvrnjDxAcM1MpY34fL1yKlw/5Ew/AEFlpG/494q9spN
6NxZO/D8psjr/joLJR62l/lW7o3e8zJmLAySUWeZ0LK5H3fz9YJH+qMFxKgG
0ytkjLCLlwmUJvj8qUlC24+okfgDuTJJFjXinxSQNRw5sbSrQ/azVWtLJ58F
sO8kjQWmB018AsYQeuhgN5xE2IlkwIXq+ivUa2gve5nzMD8ELnMWWXI83Sdz
2L+62sIC85T5huhxJ0CiUS04RQcfjKj+NiyN3WBJ9JXn1d9a1BvRSe05vT0h
hKH9EFwOiJ6X8vsgpsArqk0NbPRwS50LyBalYBfXw5/V/q1GAoEDDbCqOOBk
gQ/T/QPI+xwrROXR86jcPcaBY1AjGo9ZHcRpCTg/KNfpuOyiF0KyyEry7fRV
Cb/Z6UoaVNLc6LwIsE0VLgMxsEEESitzg7WkYUGcxFkrz4ROhOqW3NHvdMOs
TbIyvrU9Jj5jvXC+aGiUA5V4olfKPcZZzSRCtg9Bh1DbyVtmKbndHs+kXbFW
LcOqmHqmC9WVc6Teiij51S0dzdTXQ2tUeTTZEquYfe6vKoSp3mhqmWxjxLJn
+HhayEYZhsdm4KM5pbyAzxcL8Ehp9eMXQwScmhZg4JHXZPS7jxipm7ACFYQ/
HpbNXcw1++OGcBw+WZ65RMWCJnuCu6UvIpF5QBVuXp8pLqWxld02s+1vz/Nh
kUwbfaGypGGRNxNvwqnWKLO/0zKd3g8zsQfJEKio/g/XVWnsUi3uHhH35396
rcoCHMQBNM4KK4MGLAcpTCsSqiCkEpYbSwqAwPHLxQUFC/pfhs2JeT8SHzCJ
VS3XPZAbk8gcsDMm/aRPHUM1W2YBsmx+6Hvx1xUiODusL/Wsk7rvAlgdpKqK
QdI0DkTwCmPIaXSrxF/nd2n8CQ8lRhcGGN0pSEjjmyIqkh72BrJH98m05rw+
g6HxXbhQujdAcY+g9DO1hXUeuOUkvyR8kQKuawtn+2npqRGhAwlURkR8JXbG
TUAalE9z8Y1zWFjCCQNXVwAbEN14fW6p8cTugZMO9ixuZf6b0Zlu0KkW/0HC
7RK6ICIHkohRHh+51wl10QHOIp9CotpbhzVJPiNbTDW6jCk7B88/v5A+GRIf
2RLBifm0UHAV3P1R+gKDZXwxyaGgHeuJuNnABk+ufxlcamR1fbD3B15V0YbW
w9BgooeimpjOOoWSJrNM4Ujke778oYK1OwLidg/1bJr4QURdvKrdzLsXlm2P
J18BAKkS+W5qldMlGg24BpDACiej2LJueGIL+14hDYesybK+EeH2onkCnD7W
ijgX+sWIz1sLB3ib6hZhgx29QYtcDH0LF8qPUfbvDToti26VfF8CSY9vsYo7
SQns0wpU6nKSmSDC9o7HPk203KpUp6ZFkecyOaG2E1wbhMQDXT4+UgdDs9k8
+wXhn38O5MP/1Ffc4CCH/RZen3xwLEAmChoIzzNbeFHU5UdjFPI+7uXvx1AS
fFq8AJSp45wbla/cIwtAjyq7HjMmi+LvyNe9YfjcOTl3Rs1LqXrsy/BAoSEJ
euvjUts2zy2eOPCNkfS7vphyun7o1WMtA+jafwHP20Wpl7MC84zlzCGl49tm
4HAzPzea2kEC8lNZ63aHeoz5KlxAdsXOyxjiHrQ+uQ4H+12nnE/9/Sw/z7TS
Z8uPfarDqU0OSX0vocZq9WUA+Sw9cocFO79y7zwtNf4ZWKhyCZ+eiaARF77U
Iv9DWjHC8d9EU+DHqqHGH+PeVTp6gJeG/GfL2eQNU5v7Z+7kt0ogOSv4zk1s
XYdXgSAbsnR9bx27hg5KBoN0l1Iv6LifAU58wyPQuVEbx4zNeyuFvXmmjBcn
jJqSToIv2AeEKC0/YPrEj3L7F/srARAvhzhH+ubvhiWKEKdb0XgjER1K7327
7/342wuNmHvyvFylBlkpThP5F7txEdP/AmSyU82ntTEsSekbRqlqtipvBJ8x
Mj5y2DgwPG6cDfBMiQ5sS78g+3HWiDbj4Hck6Q6BAwtYuKKiJqnPQf0Jk7vp
KxoCeVKG5XocfoeJb+wiB+gT5NQuJup+sMtOGUjuKK6dsreHKypcDdXs6w03
WrI3mP8T7QkHXEDSx+5irsLAfBwhC5qw+GwyXhylDxWLwjdrMMHwZqhYqPyt
Gk9sm0MdeNiFIp9//AnQ1Fjb00tTX3up8Dw3QTBLlGZ1JB+sPpl+O6mh/CtH
H+Nd2Ozne/PNnnT6C0w0QumnM85hZIxQLQsKRrUTUqzsTwZ5MzwpMLEoo0H6
osWlooy/udRnECwq4A0ppH5DYiW1kmTyZPBCxctvMPu8geh5jbP34vj9Ibxi
K4uTbpuikp/gzEXsj0wAcAwLGRnb5irx/p3hyuKzIj102/Nq3YTJsMlI47qL
0/hgIRAc3p2CDHaFyc0WtISECjqhan/CnQcEq4wA6Fa+zstXelo/cDzvV1vE
dIta7XCNHQzKTzZ9t3lkheapdnvadd/woylse5gmtvzUYXOeoRgfujU0KcC+
9tSvZNkcHr7AMpLtntDdURVpHdn2woWQv6YvatroVHz/f/f0Ai09clhvspQJ
jSdf1IHeKLlLwQApkwdyiNtPTl4pbkbR7bgkTBUrjRKkZu8npfLufPmLI1wB
lbyKune0tejbO1a3M7h1a1BqPiD4TDq8oQzSG2Rp16JxP8h5wHDT2dBESfBK
nGmNMfYXxmQVETCAKw1FtkXQL9+VIUBBx9u+FuVUvjc58HVG0sKlCe1BZ6Lh
GT7uU8WtKuVLpTzKb69SSPuvDSN900kgE5tbFMg2g2X5rul3l2rZTska+l7D
5P6wBqmhmB843ykTVcEmGw1Pjbh6GQNCrTJog4ls4Ft+9v3b/NraoiH0yOK+
nNZXf6oWaswewOo8G7ZQ6lJrDrO3nLoym0PRLOIub0/V6o1Fa+h+xN9vRQL5
8/h+GBMoojoHrdfkxQTZxURB1hd2U5VQtLkVdCB7Wi/H8s4vWYrHBnRDYgP6
aDgu/kZvHp0j8iACiP/ff4IMCxzoxpfadurZU9SOJjPEHRqvyzJIZc0l/udO
6f0PR8ckWkCzcym2teRbAS9wDSJtUiM+9JiUUQLz+/beunGg7HeEVoT4+vY1
enbUI6ZLT1x58MLUtA/KhYWUtI8SJxeGpZpnumYmKWnQg+bVp9NXN28oZ6q5
mLSu0uwrJQhuqfuCe29Wm8Q/iew6DStmVHHmuI+yhGd2uZUO2nnD1D+u8TjZ
t2WEr3uurgdr/Wr0GrmbgkbtZSOW7SoS5Eg6YwTQ8CaCe62lGk5h5TAGWpvo
y29cyDvN8fh8EXVe1KsXCgMdm8ZLLb4cw41p3UevbFSEuk5pv07gZfl3iOJp
m3OtzBVOSliYHgPr/k+nASoWe/LPoK/i0RrwJEhJ5uF/uSLVBvH3Gb+FYszu
lRHsh8/QR0VmleH/mmwTUdUAbmWCv+gPngjs9ytZFY02aqxtdr42Oq/xcMTL
U4fmh8jUuSgFBwh3GQMbl5l6p/jkDJiG/lw8ORzb+epoRxhIt2gUUPJD3x82
oVf0cL6oPzQqpRFsEGwMZEEku1J21kOsPxAN7Bh8+FgsL3iAxHl1X6bkIWs8
C8Dk/V/NCV9iw8XpJoJVdELXfqCzhwhm1dPXEECPfR/PzUi7BzpDtQX73mVl
qA4cLDkj8hQpmd6eXDfkFpp8pfiM111LzxaLQ79lU5jUgFf+n6aVZeKUHHEr
bm4+qBkj0gXgrms2SPGMUUIzfdjf+hCpHY99ll6iCxEqtAL9DuYwufWgcyHW
g4cMbxCV0D4zYEN3+IdU+P/V9NFyCLikv01gl62t1A5V0CRwKq1+kXI7Klso
WkljRnrPRoOAmk0RmxShsljcGRY0go/BIKQA0VzHFPCnoWROqVq+ay5AmynY
OHQxGycC9lZwaD7qm+sPzNnc1aOtxwNurkssyElRDxZoqPogKuopa/281VUh
QSbIDMZbGk51CtqsfB38UhQsUoWc4XP5T9lSSqqeQxbC1/UIA3UBrITaeb/I
UgWK60cLwsoeEQhNDcdymNXCTh5G8dg+T5SF73kJNhapLNg8qiXRd4nUpOLO
oIeRVm4trejhL7KCKveUXd9PxzpFE1XkerfQU3Wbx98rwafoXntJ9dC/6du7
rg6wcBe6oe2jZnUqQKKmH8N2FBzdHF+4d6LHIc/46wYHfbesPpx87Bi3Yok/
eYTEyez+vqex+VcRkMA+8kGIwixZxnFCCkdNZRAUQ5DkwWmcZmphrk+Bw/om
7SOF/jHdkDWZA2fLEzmxFaDYBW3yJWm2LcTfa2D+iMSW9O/yZYyKaPwhxJ39
AHZnkWMhkazMygqj52oyl0XI3jrbBNOHkxdDNYleSYRkBCS3E3oXpn6zghtd
VXAGTvNRKkaRUMMTEhl2rPK4KUstMzZG46QdfKr/JTw4Zqo1WcoTMLjWXzTH
hFS/aoWvl1Ls6RJaHPDv7yfOjDzLo7KJHO4JWViDWWaB8aRn3rTB9hngw6Qo
wpUsCNeDMW6xKYKV4GALr/pfO8cGTJXJmIb0Y63/hlZKuktCuE249HPxWJcc
rmg0BP8oNK2TzYVlouSesNQKsv6vDUhJdkcYtKahBRaki22umUJZzd/Hf/GJ
farjLXnJI4ewNkJ0sbWeGmiqhZaYISP98vDD60cLA8oARhnb5pQdVs1twYnF
Iv1Isf3h0AW7NCWPFuA4AstTQjKHF9aHsKTM948T5VKhLYQQAFpNj6TS2JCi
3jfCps41J6qRKYbzKAaZ1Yatvfc+7nReRVXrG6QoiwlwdECdVRUeU8Zt5mR8
WiFDP3YCtVyjuisxeAqDM5oc/gMBGLgespz4YQmikqCFwI3rTn/Phsbd7Qr1
IpjRSIvhSTe0uj9tw0NWmSUov92rkFZGzT6cOKn05Ce6x2gMD3fwNMTyxEaa
zXhHIic1v6ImGF25Hh0WaIN0yDx4KRf3CtctYELePi/12S8R2tY0IuON6V60
ewfgOpFEjuAzR9tZNW1xykIiqX14jk9crspCJzU27QdcTnCALDLgFmyZH75+
M4gsKGndHW50ZvO6FKqg9GP0sv+/Pm91CINHmi3pC0fzHpwsWUIfwsiUDgur
qMoqX4b5ygHtrdsk245QdAItRZnKqQEvJZ3z5R7fyVYL97d6NlRAuA9R6O7O
qx+qzLSXgO1y6HRWB3uh4w2gFIGFuUUeG2/YcWbO1+rz7nJNZp5U70OE/pLH
NoPgsnkfOkBQSs1qQHB/0NVPtI2zX+gs5Y1v5hK0VQQ9cfBPoJ+/xoM8qSzw
Ydt+bt+c94UrTJaROQI4MCUN8FGpxPtvHkcIWlM1G6D21lXQAcuDQ20Deva6
E6Ozp/LsRvi+uUbovlQHX8jb2vkctfWovJn+k92tt4M1Up6isRmhArYRNVGu
BXteob0T5CA2OL+cWlPArIyqtFEUPOK7f+bZjW1vF1iKV71DqpUnsq3L9e2b
30aBCcyd6oDFxV2bL63dqCsMwg/bAiqcVLVAz/ZRo8cwO7u527szK6OymskQ
FK7e4/CUU4nl3HyvmMk1ngJsC2boLN1Ug7fbh9V8gWh4Z5kvhNLwk45gfK46
NwIiq2XdEwUhEiNC6Dmy54fLP0cq8PlxIds1fwpDzum9TUL5ZM4U07LDwF80
oVDgz1DuOeJ8vwC8L3JLxA2KQzSf8XiAJ1uLPDxKJcPH1k/LwWdjrXI4JSHR
ujWMlBE/9zNMQszdSl30BB2IhDn2ho+esPnLImo+Afm2BHwquIqXvF0iL5Co
zRMoGqno62VbTqItmRakgxKiIdWi1mEFuc3G8HoTqnpXrRdfqnQU8SGBItrp
hWsNJaDMOVueRgI6PWreDutWTDujBbM75e44mioyKLHgErSj/2THy3XJ4AoW
zUoyPYKJPoZh3t+yeO945eAg39BSFRxxyF+eJyTLFTQ0funNEkQb967aqN2B
6GND1nGYxNDqwcqsIjhg/rQyqcjrKZTSlmjSb0yjb2QljSKNnrBNxH9latXv
hrn1UBWv93Gd6I1yqPbohT2BhMMBBNBpNjDzm7FrnZradmV7gncOURI7b//G
+IZ477SX3kiS8A+2Dm9rPF6pCvTYhvERMnRFah8fLUF37kdQCEhqfbbgfUaF
W5zqsByxf3SKSe1srLhhxlVFdonjoU2RGLhrzzQmtl7QnFOA+14Xe+w71vDd
EJaA5l7kyDN7aOPF2EvUPgqt7yzfirVSwl5e0B72x0+FZEbTNOaVVM5aWuD7
yQStKDjZlvRsLiPDtxWyk7WRPyc2N2SsYjLxZALx9zH8GujEcN5Fe5Ygdpai
7Zl4EO2MJR0ZbS0r/bNf1vUyhwm2uCTLOZqcmC950LRbWfsCziOIn5i3cfLc
cghX5lU8Qk0omvkASPsq74jjf/J7XwOug/VsmwMXoKBhnZPtj+2E05bMdu0g
IfsU0vA0ymCkXOfLUM7yXJ7Uh4/jrrCvE3WBs2U3Y48Q9Lmm7HCn9TwaoG3T
Usj66mGUCyACDhkLeHKJI4WJHB29z036ov4ZIMO3HNonB/OwOVzf0SIihkfl
nyDfFbOWJkK4YkpQxqpD/HeeS0+1qkuXh0z7/Mo5N1oL9J+cFhk9zBefnS9X
UmMKBrAzuv3I3nbtv4lp/07qTqpXSARqWcHBt1QBSJXeBkDgZZTbJsd3QAd5
7ZRPvFfGC+hsbTDAo5tLXM5OsFKr50/Y980/fcfU9xN6eYGFcnZ9H6y8uMgi
GDvP2LGy8HWlE7NoBQ/xCaa47/31ArwjY1RF2lrnvSnTCj3ckf5w21Ho5nVZ
Yf4tF3iiXoE9awXNqeu5m4TJZVjePYikWVWMSSPBNbL4jFGQdHdnPyyF6idz
K225kr18Ku0Ssaq5YOn1vGZKfINZwLnjbOSD8luQq1ruJiQOvjeIIU7mra4U
vHDcHFSd1vWY4FJH3IQbllUPEmPxS0o3WYEH/hTs99TI+HqzEe9PodZbMQL+
vY2moCGfk/QCvTYZiIBisfnz8OLzUKKFSvnbLkXdS0aQAe+iDg7+M6MINnoq
ncYtMg6LTShBFJ+aclD+DsmDqbvG8P5BHhqM/oSJEmuV7uOgt3bqtDV8MZ4v
/DNHBREFX972fZ7tQuC8j5/XUqmqrr2ggycZpLXv1x50UxdhmPnaJDEiSYDY
pCXIsSth2CIFazSkJz2h2+voeqxI6JFRJC5Tc7djgfGugT7xS2JaNvxVBRKa
cr0CErIoXbesBn0pvQ8MkYOsZzlOVGIhE65LmnTuxY+E4V/ZwtXXfaEo4zON
O3UsgmXx4U6D8LJnLWBXKC/sRlsJ5evHCldQ2XzWg+Jx8D9xi1nmKp2pgvDc
mxWJEO0bcvQqXV+wVwGedNE8zkpYEGaHXpT60UO2F4HTHvmwfeSFze3Y9RY1
iPwRicN+mqbGEjtFuw3N+BBIkx5/rpQRG84FRLBkErHluh7r8OsJk4pq+p2o
z+u9cW5K4H6OIvenhpWDl1YCkil0t9qo49MOUiJwL9sWEE6OxT08bio11mU4
Tv69wupALXLOx3ip7MvJsTOGS0QYmqQ/vzhs4Z9LnRvGcRAyEOn0lwlX8jtl
i4nr+ozer/HdtnuABvJR4MwM1aRF/FSgQfbQuG/Ow9B5EIWJseN5zjNNVRjH
ejyBGKzTHxlFKU9+Y/2gYQY2rifwescfGLroKMx8pE2yIZ9oMGKpVCNARvU2
0A4LD+xs6pQ9bZRTG0DqCT6igRHTSPoOmXlg9q+GzTt9se9ru555xh6GCOmZ
ICTiAyqM+D6UVWshKHpSU9OFj/C2kRHke++eXPbdGCNiNbElgKFCn8shlWDO
Mo6Cq+V7/npXS8cHZ/MOpOzqSwf7qXLDMpsHolir9kjU87ExT88RL7+QAV9q
ChHrKkZFlP6lfq3g2TisTV1bGC9ZlN7z14FfihvWvnf+5gthzP5vL7whO0sg
dkNj1Kgh3l4yn3LIQa6rS3RfvH3CyxD5zV1a74+Kp/+1MDhAQVdZmqjbb3wU
Iejp0q0fKyWMlfKCEisCzW8eu3cZr53hEkMXFmgyWdZA8foMZq6TDvjtG2TP
dlNyI1YElWWxShuQhEChjoSDUNgM5U3E31VNulkR5BYq9AtNIwV3J2pXmDmJ
CIahaEWficMFhMAoK1sKm5X014EMfS8T86UOrRALNK2NviBhQqOljQUA28w1
TjgYAB5ED/BYTUR545A8Tm8jHvl5TRaYi4NlNy164Haw4w7wxx3LxvomW1wE
tOc8kLhm4pm1cDO6FroXZID1I3CNoTGTWqDGufx9E3x7EqZ9wH4baxulFQsF
b9kseBQw0ADbElGANuQqz91YtAmYw7DDr3iQ6ktfy0NOKpdt/Rp3okJOymJ/
HCtL8X4C6fhB/m7GQ3mf/OYLl5jjbb1Fgdg2zhrWBlW+AvMrZ0mZaC8+hzD7
UWACdSUopIV9Iu3I1ho1VnuTOLSEUHI6M35tWVQlTCeG4UlVz/t4mussxVBq
NOtuXKKIK3BiPOpnQcpVIx+7JBToZmdM+LljvA2X5YmaPNhpjMxVUDRl8KWE
JhwMqR8S3ARXYxhiyK7YuFtel4HOG6RZe1L8fFkG9kISXsejfNkHYaPwE9vx
2UoxHxwf+1OYGK+XW4bU+nXBGD/sPFq1KND+uajEdZ74YlhICpNHQZrSc0Sa
4gJFIdqCSsjO31UP6hyl83WEn/e9VQVeITS7Z12VGL7cVNBE3MKcGj53SqLU
zxRkzjRZ+HlTzjP0yfrqVKfg9LNFjW7qPmMKlR5zDnUjjJbuKmQDWc6fnC9b
l0w3br5Nriy2/MC3OilcRm8MpFVCnz4+tYlxGoyLMPMJXa4Oj6y47eKlIVdz
KYSCA7jjUWN9S5HoCf3+5/dXX9gHHbNtxwki0HRGU9OTyk6bDXG6kscdql16
9yngVQHt6/xQP2oZzWaX0aF7gQvEeH9iK5Xx0NVHhzni7JqYPWbnuEZI4KfV
YaVbH2tFD4FwM2GK4OddWCSe6NDgrE3lYiHIks28oPbkZBnKl1NkzZVG3EQp
77cJj3ljuSanKCHmJKPLscz4Pgjzk0ahAhieZ37dCFO7bTncMTgXUYZKlTBv
MxLtuG9gUBEDvdQcs04ezxcXkE6vFcU2uGdZbFjubEbe2q/sJJ58/dwcLvG+
S1BYQR2EKuqOtvsDu0RC3r+ZpEHMGe4fl3lS6EG76jcGwK/yrV1LKoOCFpef
RStdwPsPWDbkfLuKWKFNy4+9ISFawpqxaKpfaSZZe2HFezRqKZ5xglBZJWcy
l1ZV64wL9/J49yyV3y0vYXFN3mjiDW1VgyV8f06Sgm+aUxOe773Mu6papcAZ
IpLQjOQerwkYWh8mqT3DAB0C74YfPXRyDgAx/8geKALROsAYFdVZsELyLzOg
pHcKQkj6y0YwHEKfKGAjjuuIT1VMvXp+R8ZMnKLh9IsLnWWyypXAWpLSFcDt
zsKhFMyO83+2Uj0c83sPenrSxfKNFFXuUS9Bd3xilSqKVtsUY85e/wBqu3Ij
41dkunxLXO8sJm/Tmtf/+0AdiJ/QrqVvZjWZhOh4vWuk9CbZAWsxLtCRFiY5
vrGqLrUWB6HruKMvxqn4D4RXfQ7JpuYplCucY5a1V1yizAErhYxZ8zpRtYyZ
vN5HpoG1FtVeo2LtytcEQgLaj5S546qvhex9nfDEUhEfOQmN7e8W/pG+6i29
xf2mEi7KZ+BjC6B1EqgUbnvPMaUI+0xxaAeSAmKRyixhinHT+rKKbM20Qt5s
og3LsNUDSAfDwaXO82QqK48C4bCZYN5p+X+ZH+EiFc2jeY4N9Fr6NAywdzcp
AP+Wm/aUYH4SX6b5slOWfoNg6UG3M1RK6JUk94ea3W4PeaoGjXKhT5lKscoR
Z+s0vL+MjP3Vx92aVkYuzvQ7pVeyR+CBtP62kX1UMagdbD6gmaUIqI8Q+LSj
Dye/Hnxd2pHZ6pVUfU78q0zuU33VqKmkA4EPPRZKFmaysMvmeePr7rWXHFqT
ggJDeUIMz+1TpZG+UFLqfEpG2xGd/jIGxh9m+k0Y446muJtf1lYGjBMMfB/i
j0B79ECycBdOYrXNHzpSvGffaDaxBzWt/YnRoVfE+8y21/fyeIpq6TQcrTwK
Dk5jsHVQt6qCn3NxQGRtNeLyvZp9GA+P6+dAUff/3W16b01vxPkZGCqSrmdQ
kyuE32Cb5+0OnKJ0QAeP9WlEBBG3PpJoHDkVUDKmV5pIv1JBMZFhQaZVTJq1
Xv/ctu3gef21pgU87tWqXvbr2RxdKDmGSPDHqW3w7ZxEO3jJui+B3R3n6egj
eMlyLZUoiVlzHUDF9nw5S2Nu7C6mIVU0+P3+lpHEtJpwzIrOYOlenFFULI3S
PGPAL61H595fMuZXDSnySuDmJCz3bsyfPqRpb0sM3cA+crI1v7uLy9oT2ZDB
NaqXKh0ej2xS71Vmq3BrYy/cJwehUeJOcFfhprY2LcruINOUjPalBeGY5lHw
l2YwvsLL41jYlIJYBhV9muHnFHguw7TVFqDWPgfbnVFGdVNpEes4y/PK1SbU
CdznO+jj965pZWB9RdRR8s1ilForrWn/UzKE85UQh45ARbcbVFaf8ev/zU45
5ex9yWQ5foFN+kh0/yN6W4WXlKcMXdEDF5SfAiG9x/uBqdzJueVJuVOl/56e
81dJD6FFG3CvOpOi98xuz4arPW98I2DNoG62DZ6YcxxrTouDzZ+JRu4B5bhG
dpVCUCwaNd7SKTKztfJQjTUGJVHM0EhMxiMcqmDJvbAe3786/iXp6ssKxL6x
d72Lb/FU9lcmPCx5xQP8gJoZUzgQaq8LWZDTrdrnGrtLkg7VjN6tKgT4qatZ
Az4bhHTdjO9RJlFX4znws0dFm5gYB64KeKXsM+8TXRAznLaiTpzwExDKf6O8
q59HrXGrdNguljgyMh+sa/u4fdOOTQ2Dj0Uaa/pHk0FGv40r8GvUqam9opy8
Xic58n8KABbFiTNoPfYfE9YnWN73zEKlU1rMNMuKQbNODEQ5RLMk9sc1pLIs
pflikpKBbPjhA0aya56PkQsDJLKbOsqeewE+ZQiAO8vpqB05BevXrCEBBCwt
YoKi3dOlIM5+ne74iB589ffZENzyl/Q8LjNzmd1ro5Xi9Qo19Tg5Ee5oodlr
ktGlgftRNTEkukuzCm4CWXzq2R9/R+QtFfXtIPTGxAz7EckZZN+I5+EIn6iF
KWx9FqK7nQC105hh9VZjXLg2zpXAZAtP96yGKpe+Z262oLGk/FofUf9Ll6Tr
4fb5yHRQBsjqioZGVtrrKOz68OMFmnXFUUncxF4L40iytECCyShnnp0DCITS
01vhTeLtGJV6IkB/qObw9OverbOBNHKTrTkUKD7bS4LEexn0UzXLH0djgNUM
qF5Q+DxrBMjBcekReQERpYY69IuOngoTA1CtnyzfxvTrWrOW94ye7LsSDXj4
my4BrcyjA8J65d7yOHGD6iOsAE+qRQOAUCatrzknGI6tVLwksYW/MSliIUxm
FJRNsnSjGXqndiBlicqYcqaZdBYythetJHBD89k8buEYzdqhZQZKjQiIpkWG
R73ZqlDQXO63QGdCdtLcECgfAj1MrwZ3vvTL/qRF6oqfC3JheiDSOmDk1iQw
G+zXXLamhqcvmbER+dbh0SH5hWnbzrPhkdiJjjS+AAVBU+8zjMuX3zxnqreH
E52CfjUN8/uy6bcdrzmQb2NVg66lQB1inwBQuqX71allingDYMxBClduAgay
9I2kHqt2Rfbi9esJzemlJHAiIx0L2NVEYuPY3+8rTyyAByU8DpXnu8RzdHqx
MLoSkM2lcQ/HK47TFgDbOHZIFDqjuF6MniFUKZ30YkdlBLCC7YhF8P89UIRO
jRNmbhemJsfUKHMy8Pq2A77rM/RwboJImXG696f7AwrZOfHnMsul26rLWhAY
YehqHJYYovKaTnGdU1tM+GQhSnSAgMpp1ojfACRbBwrxz7I+Gmzu0Ir4tcRY
/UNQDnSx5lSBsjYG55T3e5Gf1S4SBbA/p877ui6SP/sxoULqlijOhO1rXJgN
SNzbd2ybK7c1dItYfvg4i5Z+OBEMG8rjt9RWJ+1ZkEYBMJGErp8hwFf1UCHP
T7OCsu9t5JmTmaYwyHWxA//QPNx3kRsnasT2pjZN/opCOChdW5gwe1gsXiix
SWBTaNCoiNQWqbdz3YJhcARM3VErdFbbJCv495dPjCSKNpCgC3wdp0SbClyk
+vl6/K6jqZ5HVZ296W4TPs9cEQigkN8O5q/SgFFm301fwH8wzwOeGWzcoM7f
meJwkuEUt0FIuzNvcjgguKHae2fg3qNXTferLS4ZJ9U2QQoyEEyy/RNGwe8Y
Fj1njHK3+VPAi1DMn4L02X7/MGulOq8i0lWFQsEofN1oL0KnvoThqY96nHWe
WrQe1AatIEi6UZFdY5sVG6ummc9hib8RE9TWza4adjjPA0WrG8Qd2srJieYk
wbusrWjKBZmyJPLUAKy7ZE+yrdbkhPcCSOYQjSYKsEQIOwmZBn5RzDO9/fSa
+4OCo5j/FInfkpWw8XMXunzUmE6NnRDibpHjVf1vU2w5xkdIVcXqMhQs4PG7
ck7fNBmorSJs/tduJS7axPhRL9kKK2E99BWvhGLl6XMtHI3tATM7gVFmiDpA
Lbq70lHXJTY3NKAzmObKn3phgOCdv5YQjLuzpDhUCS+PMoYZXnKWY32rKQkF
/tThi7QdLMPGc00fSSdxd8SgCCNpUnyi3DT+fDftg65cvIEOVt6BXEV6J7/c
82ChD7lVE4pxfbccTvrUPAzYT5DWf8Yagu0irvpGcVBmnK1N3RojeDSqQnrA
n081gAbSVouQhJcgNYFmRZ/0u3OHr2TbvoB17dS8SC8TLsdJB9ipuQH3RaPm
2Oaok/ozC2CJdHm1y7V+7zpizguH0UFdMO+TWl1j39RNqGDFpx3aeComQkl1
Wah2hawXnT3DtYIk1Do8IdiRvexG3xBOijFHoPCFwGnw65gLfSAeeAyDAlXy
o0KZRrys3lMMfUamAuGMcudLTK+eAUntko+gGaTzlUCGvnGhWqbo6KdxdLLi
Wn4q1Ngq00i2HGRjnnsOc4CUFUNVsrIF4IklMWKXE03DjJ0091nWG808KR2Q
TjLILhg8iWKjg2ixF6rSumvG2f3QSipeXDReOXNVqqMS2/It79kR1sKHZml/
jjE+pkjrGXH+8hyz8Lt/qohOFLSsgbL/cnBFgdPe9Sfwk6Lc4rkBy0Mt+mNO
eK7Hc8uL6AdruXEd2+2TGeTLsuvsqYowr3RfHqiuqwazgVvPFs5PlHB9bDmj
8d+LfRP92RZUpIv3U8NpkTQoUgtzt7IP5FH83FG/sUArW8T5gS//mSQ7AGYR
fhXTMIoUPhaGPQU5zgu6fszSw9zY7q9tgXcELunOXqn0EsEhbU9uW7n/J5tR
rxlw7UPJw0c+vhkwKupv5T6pweBnU87wJ9Oj0E566gzlwvLpix2PUd1ilZsX
KbIpMvbLjJvTH3Pyes4cK0fkfVRREDkc4NdW91wm6VMhiy5aaPT8yvVoQV65
2YxfD6A8gXdGm5HaInp7PbaNJfv0gV7mDbn/eOAphEmMciIntD3gpjTQSJ3c
e4pq6CSVarAB0l3DwQ832RF6dmRSgzY3T0J1C3VIIjYzCe8SlAV03DjXKXPH
ydx/tGpo7hcaQbt5xJZ1iSuAe95kKlUuRcGhr8t4JBVKWCkayTCTmERMMm6S
9YFXxtndpqGdQKgXu6i9XOqgSsTq8s3PVSM0aW+cztpiQZvHWsv3c11cMeHW
bB0TGwIR0vLQ6NaSefrSbIOhy5GXrfoud6N3r4OaLMNTGhnDHyIiWhmQk+iG
VSur7aDY8kTYDvAMA/MJniYFAkT0b0kdS7wbwoeuelE/o3/J+keXadTyCVct
VSz+sZLN6DWYCxBrM6l1+nBNWj/RCyFjm+Eh9hv9I8MA5JsuFAbJVBzkclhi
K2PeGzxWR9URmBm/PdRJpX3yAlzEIdr18TOkFIOQ//nMDqtW4mcjGsp34DQE
jNXf9qwI9lLN5aqL2JRZ5jPn65NmF7d3zhmZNLWzeP7Mrhk+Q3yRzcU+/4pf
bEDC0tJQv6RAHMaiFJxcjPqskYiYkGWme7QmxZSht4+riC2NcD/ja61WgOtx
nMtmQW9Uez3A6wXReo5WsMNKtOhoh0GWomqYfJl3DA0SGSyCGB5wrCqQ5Vx5
gLT2qCmQ64jAIgyjXIcZY49ksJGCxOaUGeejBZk87fJfwFSaFbgoS4PcB6sG
LN44x+zk8dPASWeUNQSSqS+PHfd37q+t+EFZCZUcYWbJyny4EZ7WdNZbHGtA
uGYh+SA45eP5CWvzmPi2gb+WpeZpqf8w/GNg73IF3eq2+bP1cI5gE23U8LAm
74/xDdCJFipHufeSpRffMdIM3cnpNZ9RoJPioXqTY+dtDutfjX2fBN0kmjjm
fT+nZ7XvgvTSdJM3bph/37DiKsJh1hZmSn/bzjzxTKAChRVFK1jQdDB9o2sa
WiVgIvse+fT7+f+tU86HR0ZsWEn94SQkz1O6U7+HvwPNrikFtP5PdjxlEGvr
ZBOyXqLUoVV1JxJadhGHdWo2rol5lG9oY4CJ1b12KOmMw9Yje2/Tm4KpKwbq
a53HtnMH8+srCe8uALPdtvzXTjbhuLDT9uGn2+Bytjtp56oGAEAgZwFS5yvD
ugxxb3ELlKXYEgNcYMt2+axlNWQBaBgrA6eOlCDUQsZoTpCl0cvGzHSYCg/T
SDHIqf59zsktDpjIixdF3Mf3f+M4L2NegzrA2vuQTxxOZDY3Yud8oM9hFdAg
RlTidV1WxhF+qyxrhrG2+cdTEm8Znga8XjpgfElhuvieT+pDgBs4tVU4Ibp6
+lH46M7RNb8eu+XYA+NU6+aP9i+yN/tRlMkZhBxgyV2TZZvio9w8E9zV50RC
PbxytHQhOfhQvg8i0rqOI5wvTCRG8CWdFekjpSxpTek4NTden19URS4duMg1
yCc0iOcb9qa1dnEDQQBRir8+Inb2f+s/ZGujxjBjFN6w/up0P/co8tzIwIOw
nOxx/cNbN6CrbVnJIdSJyCpsy/zfcbiB0C/dG+f5aS4iscs5iPmmc+vJzzIt
pnKNxpQYXb+8yX+SYkR9QUIEzEND44OCwHwntwiQ01mxIUlAA/+x8/8T0CeB
dfMJKCCRTP82ssRXNrQgZs3Pkfx/ClBx/zlRNBCQM3QmksJefYgXUugfxhHa
OersZ6al7zQtf8Exfa+cH34ZuO8k20zDhbAnL1Ab2aKIbnf8iL1nVpuvW2SL
38iGnp0uOe/ggh6VsMebFzCY7qT1jGT6XymsA9K5or7OxynAgq7OVBOTYFO8
xXb4UO6KXleOr8wFzjpbr0QwYuJ8pfYSHpamcQcqIIZiEOsZVdy3tcbV8OXy
EsOpIBb7uoR17jBKSSlrEp7fArW01d+leBFapBBFRmH7H+USLFiMTSquRNpF
ys0kRFJqJcK1uo8hdqSNykvJlDFXSvORRbQE9qjAGZ48582Vn98Qx9UDizT5
Hh5OAz/Arcqi/As1CW4HYJze71xowKayTBzzEWbAHHMVhnQUZwE4477jDfuN
ThrOmi/zAsqhdcDSJGaZSiKuQu03ODnY8fk/kUdb4KCTqjKQOBmiflS2q7ti
e/A+vAEHoH6oBqgACLbpsdrsd3+a6b4+uHf7kmq5URPkh2RnJKE29+ZPpM/e
uNs5of4JrajvfUXeaunFOnQwMIQbQPOFHQeJIyvKWTMai4ItcjLPpFwtQhxH
IuAaMfZJsi1FpOXRq31K1OVDVTPsn44i9u496rhTFPomFtCwqiKtR0+uY/fv
qSboLDm7Ze6VLcdA7pHAKVi6a45qJRhN3brtJXXy95UBIEyTL2eW7mwjpP6L
byE4+krROd1GSXD2l/nchrYh9NKnlOKUXznHhRtEfBb7ltRO+YCor2dJSfg/
GhC2zsdFAPAxtE3rNYWs63KiTFgTPEOw2lxoHGphFLgTUY8Sx/6p2nsNIDMN
KHRbxh5i0MJcyDi+TbL3gXhvI9njDwXxNqHMk3FuZFopSdbvX1Ug3FHuUHmY
Gm1Dv14fsuwv4K15L6/54ojb1mAh9t4JTOPJZ5hb8PFuPMPeU8eREN4Heaoi
hIGNqyEE44J1c6MeUWCm8u9BLVyo975A+N8z/aSJvnXQ/Q6Bn6Cli3wcAS0b
7XwKGUIWvoxo9OHagJDNKXnGI9Wmh1K3/36RDgkx88Yk3ra5req13SSvwBpe
n9HsBFTYnx9maJ21Z9FgpVGdcqsQaSId3b1UOq21FFvd/jy03wtauF82dX5g
wQrqcr7qs0Zf2pjPlcG80EFb9ntRTbrVgBjfC/ROJVFUol0sPW4ubf+15Xa6
Y3i0T2ZDU5L83u/zgqXGuKpGFDLiNuR2N1O/q/6lcChKwYTPlJz7TifUQyIK
AWpx+BBPUxvF8VKogiNd5Kc40FK9GtxozYf6MC+gJV7+HQdL2txqFuihFGmc
Jn+7WntpOfnZxuIp/2io4/5fjsfi8UFu95xBqWDcPz4VZCNVLbrkNH1k/e+w
eESi0ZtM9aaTmSpbucRj6NOa/yKEpxg41RRELF5nyjc3J5Ok6Q6AiIFGRpGY
4cNLXvg17lIaWAMRf3xDYjiz9oEhEJa/Znu8tlqzL2OiGD8uI7fBXqU09bUK
keS/948wGAhuM0OWyblWE/ghzanz+1+hOVGg9ydPDXKrXi53hE1hMFMlLNRh
cm74Lvunz1tD5lJK6zt/1GNrQSbDAc2mIdqACp6nVDuH2XqkSWr9ujnMPV80
YXfS2lSlO0Qz2rtLAfh9GU1+hpZWQRRsXszYQuFtYGRzeDJ8wawutP1uXvur
WSV4Qt5Ne6caYCLMiHm3M5kE9pzB3aD86FuD4vL7qQt9CSarr1FRIb4HZpjd
FZ732Mya0E9JbKaacImSvxIyuw9aU0VuRZ/V3d8HCveGwcfcMAghuak2pDW4
B04x4o5HeV4Fn7oSV8D4YvzqbgCFtLTMJIRwS4npKEN2rAg1h6rjYDoJzIVX
9yKey43M3OC0K6ng2gqq7HyRnpYC9vYLIhecVpPCRJadmtqfCEwInHlajOqo
P632x5pZFvrm0TeG6NE4tJB24NofT9ZGOsiLs7XYxl9BosLRbZ5QTEHINCiU
nTLAhX/6Tuk+bjEnT0dFT/k28P8V0ATOKwslX7Xd2eoBX6fp4VBAAX2ktjrJ
mnPivgwEJsoGOVO97dKMtVs/Y7FlVWR2ZpaUnJ4AVSmjdzx9q61uPlBXvOf1
gEEIVs+PGwlHQ3yTUid7+DqvEGT951CRW7VSHuwiH6h4g1nyCeLXw/JsmAxL
8Bwmp7GZD1EjOHXxEJFkagaorbTviVW7nU16n0lm2UvX+o7CwuyVo7HAJiqs
8P84TMlMB6zmqeWAO1mZhTbs6xFy/2HGGHx0upZJpRLDCi2jZ7aHQW+TBTJx
cpkqSk087ko6/aCsESsFJOcVO2kuioBUxXl4/uO8NUd9SA7z+QHMCVo50hKA
6Zom1qb0jAJGiisHuKU+7eB5JQAOTrFPHNz8JJMkAMtorxChDJx0s720UoKs
H5ojxd70MdV6LCk/VdFbs71mPntl4x34/x0aLTjO9saGZ3lgVlJVVyr0qNXa
g47WUhqtdVectmvrlaBIJTq6VB6mce9okPXFmd5xLMVqxvMTjHioupP7fd5l
XzqSxS/Tw0y4yQ6KEKdYxSQJcKzc9b62KKrY0SvbS9d/e79apL6uLRRUryUg
/M1NsvJ1nb+AJcdya3RyeMLhQVbD5egGXAtqFyknTA84Dlc4I7sVE7NLxxZ9
c2ExOpVfzVg++BdWGDnk98o46qiTqaM1GSquNGp3bTDxrSDQx4biAPWkeyHa
rYawyUgn4iWCVGvmOTaRkV1rii3gJnqVXH+7L26Ltd27UZzrPZmgYkabFXs4
j5wg1jOUqVt/8babsF3ic19yE4ddjpjFgelopnmZZhkfPRPTMsNoJzhLsadQ
AfVhsSqIi1cN/SqRNWpKjTDA+0YVlvWuoaiimlz+g+QhwYAjwnWd8e+xO+Gt
FB5xODeXlQ3G7wJ1Uxv8dvHqF4M7BIWg1TeQcudwNBg/zz+qcPaNwv8DmaFa
KlHoaCOxmtpBC2seX+RVaxpGShT6v1DdrnW20Bp67v8YeLKjaiaBRCvdeESy
ORYDUh38GOHv7AT+m3GNX0qXKhw/iZLy/dVm+j52FGTaxXPIv75PU1n5ge9i
6+TYjIMGX1PE9WYD2uFXd29zLIwLZy0yySoPjC1o1kMeB9x8vCi3XdZn8W40
7fU7XobkWaZuMXN8miKitC2j8TI3MIRjzJi0FmxDP7kChtXxbZMPuT0BucfW
WAQutuFhr71YFSFIW8veL90G/ocg9Bdws9ykDq1cM2G1M6aQPJkJz0P4d8dw
o+t9HH7bybw2MSFVBCMi2Uk5d++2S1NHuGsNI4/TwMyRaQ3SCp9zIrffqoZK
0hmTxF/zYkDETsoBWRubf3Lv9f7uNXdHezqesxKX7/+9k+tzEuiTkR3YBUwP
F9RnkhwP0NdUz+hXZM6FucoE5lyKbK1IL1tYnVb4sl6qrsbHpfSY7rUDW95d
4EpIfi1eOEw9Grlfk7y/sefRX2sMiVIOfb7RRgxZuTD+jDGoa8vfzp/522+v
3nCf75YPEo7NP78FjXQSUka4C4t+Qw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "hmRb1hCms2kg5lxwgzvVC1ojkYPyZtVhUZroYIGDp3nv41l/XQfn8gMXcNw31HDDWBFvru7tQ/av+VlNCOY8CAEc3dS4tSN1iCLWoSLzjcf1An3u0nZDKunxPUWY57wMTkfTn6dFEXYBYGQG/cgNqAwhgy/sA9kmZ+yrzAG/xfCgRlDUR3RpN+hQPPycj5HNM2pIgRPAeD/5T2qj/frBFu5c2+SfDL19Hg79cXZFl7VeOps0cLpeAUG14n9bup04lJNvUvDosxI+S5hm7k9jBU/Wx+dlV7hgTVPhI/GnhI0+yjq65OEbClAJl30sRmlDPgOGgToMfot02ZFGpKyPldO+4dHKtQle6N0NTVxZqyaz6svfejlrnguJIj6eXVjoFyKXsqXmLg9BiCQrQykdki8vvLupl6k8UtQePtCg0xL7INxlHaS8WE0sucNAORxEZopqbhAsycZx6sEYH3DwcBy9Nfhp6CCSHbO6bstJGo8M+ITaYjjH14X4J+tsl20aRLm/V13Brb0DHOeQhWHJ6FpV3XfCaaFu9H0BgSg0x9dIpHrbW+J3VvP+ev3A0FnCD+ARN/1mDWh+V6PTc2ePMbWGjbAWpUU3Hbn3AzM9+6LNBrfZAtUi2a/xZmhl/eZQAL90wmrvDvBRwaGwYYp8NTXBYkYFxu9jCxfBMpIs4iAwmvUXlz6FuQ3h/pT2QjSLiFN180dog9kqAIXAutw5WZUUQRfCEbshyIFGNR9F7I++/pWxG/1ASCLh25gLNDdQcPDHqiQvL0Qgq+MNvx7jsvSPS3rExUcD0Rq+fwzXJovNyRJQljnCXF+eYXbFacdlh1j4BCAwsQrqFqlcWewJ3S+CpU7eCVMxFfrgQledQg4Fl06m2B9JHDbjonpDdARhQzGB7LvLNgyILJz7zy5fxN6ywCm9s8G79B7SOBa3FTVFuxivmgP3yCTm0pqYMLuIhKdey8gYJ0/Ukbjb9AQ4wUB87OCNfRzsyiDnd+koU1/5ZV+rVW7jwlbhlWXM8UkP"
`endif