// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kMMoeFjrZFhT8uOktnDm/FOLRxvBpCwkJBdWJks+drPh/ph/xOEAZoqAkdxa
kVG1jVeE1qaOHYtfZIb8mjnMFihre59XCVgd2BZw0IMy3zpRDlsKzy5G/V2g
TGFIUgWs8eVDovJTqUX2YGqUGdoozuqufsmVRnLctflLjMX+LavjfF9qGA29
SoXUWrJoDrzd7lm8JQtxmSlEdlccFUcn/foEQIwyjnZp5GStVaGjMGI0XXwf
RpwAuSgq6vW6+2NCFOmTS185YXFW5swUBrkoVq76RfnH7LWZ8NK2XOgP6O1J
JocbVHfa4bPuOEplMAk2wDTO4f0ayYlyBqfkiNiwUg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qsUMH6ARTiQa2dBiH5aVPnNKr0OpVCAwIbnanVph1k1ED0INIoaQf5b8N2Nq
uFjXE2RjI6T7IyfaCide9JMde8RlthgBPE5O5CeP3FOOgYbNJ/m01iVtb6dm
a7E8Jmn1u7Q2UuxcCAREDjv/GO7rwx9QHyv8nofo66KYx17j7iKLqcZpS9Mq
9coFLX/zJN6WAEWdQEuVSi4dVjzav4Kt0j9vLiTo6EN3Aumjxxvqg5FJtQ4+
9eotgFyS/nFupCsEG6lwtODgc7ZNMyq6l2+14lYRLV+VXck7xoTPjAm9txzA
ob0r6brhi1vud9jwmVKMvYi0amFxqReNJPveuLZxHQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gJiaobeCzaZ1oQ/R+cvwSAsak3OzBeIYU3hVcanY9HdBcMVA9gwJmOwQtbx5
qqhvzVsg3ikJwk9/tR3EX5qtYBs4+jLshIrUdQBdcr5b/Vbb0jL1VRczX1im
vKHCKZVmXYCR+rP4PDZDneTpOt6p3lOvIImTXOasjJzo1m/m2YbxeHT271mx
7rOZerVk9bvO1rL2Oxjjh6kpbHNqQ12FubVkyKRDDjpIECviRCoXM3jj82Mh
IV7n5EMfBKre62Vm3VRQa80b+N4XdXPAKa5JaI0ON3jaSAsgWLU045v83/iX
QLFhXwhtHCeY648e6w3upfuhTzYymCTXHHJbJ0FJQQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MC2T1CBiGZsUwAp6UPxeDtFHBx9mfr0rGKIfPBscu0QMkM64QdgvVYV3gxVq
gmjNInh9vS6hk/6N6G+f6HIZWNSxTLcls2m2pvHVNlTSvGPmb+b3+VyDDTjI
rjKcdrWnbn7tq+9EZwr6o1b0PJ27JTYoHWf3dJ6NgM85JEgDxYPzOMiBYyyt
sZVb/DOsrXd3VfmQiUiODyjVbIObKs7JGHg8I9eboVdZqc3W7v/PDg37OCLN
AqhEelAvXrxQR/FkJYWZs0P2IoSBewQ1DTvMlZC+K96fLHuUI7ge1Tiz+O8a
5fhEIt84Lf50jQb+TZ7zObaNe+PP/jEtjyMUaCkNDA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ideT1eqezww2BYyKhawyvNHkJduSWvRqQBPKx8E07IJSKAEQ9tS7tT2+n/C6
vYzJ6/oNSSNXuWSgwessYSi2CjXoQRwg7zM9PCkcYU3aILSOYxxv8QX4MUDH
Unw/m1xN+Sut5RdRgy3/grA3nHNXlOhKmGT6eMB/uXqGtF6+oCs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QWywnXP8p8BMWVU9VX3o8msEo5vo6a9f5iTih1OCnQX+hfd/HjdROhNTuppO
emgHkhHgGcKoQO+zDmCJGXhcskuWrezOf+sdQ6n5UQk9IV9XwsaMIX956NUE
j8DC3SQC+OtQvnAixc5ZcH0escbLeNkv/NffLCkvOb8vQE96K00jd99C6MJz
V0wPYLqaByK7/gx5pWDn4O/FfWqf0Lj30PkxPzakBOXshs1mP4aRnfidmQyw
RO8IQx5DJOwaE2IJ8wNAkj28N2aDdF8OTCMHLzGgVgKayIYa7smequxJ7zxc
7FxLEmorL9UL3Id7Qul8V85qxeLsO3V5M4c5z4bHfQOYndu3vQ4YdhQJ8RVU
3CZRkyOU/NXRXgseJ3++CtRYdhaVKhstCNsiA92INSZJY+gYMTGEmgi8SiIg
ZutlQAtmLbMAVBnhV6MZWei8ASeixePojLpQogUPBbQ7hFqQ4iQdbAbwBsAb
92bhSs8pG8zwTmN5KfXO/8oQkr0CbnSL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ikIi1O/YRz68o2lA+P0lrYBRZz6w35W1vwdBTEuAwK7z+Mquew0cGNwYhCbt
hl4CYFqozalgguvqa8hkH2jeXuef2uzO46wDq48oIu6XWCVfH0eNcxCtY+3A
UDZ5kzqa33fJpCHq1pMUSLt3szOLi82PqV7Sa1w1jF4xbzCJb/4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
drclnDthfWLI7uawUAcP64JmqxTTVnM9fr09Fac3o4HsxQMWYGXIekxRz1Yt
6o75/TuD3zDCSgw8h/SyuF+jIBsgIP7UKxqRDiTIfLKIcOlRESXU5OWeUV53
/hmT/np7oR5/KOAaaYwmWspp2tW7We9SQQSuoFE9fxpxvGoznIs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 54384)
`pragma protect data_block
kmtntU5UIukwiZbsJmLy/mix0qwgNXdIG3Q8Xk5gNNCYcdvY0UHiJoYsIv5i
rIYFST+U+E8eQpulqfFLTtZ2476Siv1lObzJdgnI8maWaNXLql6U/G1qaAMj
yLmcmzOurivSJKVKhJzV5jUBiROxkVJldkkc8wgr7E1IymJcesQh5Nr6Jzor
vkBZ/8T+m4K6WRvN+RlGgWuvJEavWYySWk69GYfQvlr97IvLsZEDb9By74PZ
+u4Jw79fP4C+wFtaigy+QwmDwlaPx6yO52MjI1VXbsQR9DWNN1jcI0Rj8Sch
MJwwpQi3+14MZ1gKvJZwpZpBiTF0kZX0fkDY1Y26y9XbpiPNMm07xT8g3yCk
zHUyRMWvukWCu1w5fbvoYG37YxvjtTjRzaxxrt78azCXSqWgKRlI0GcKKtPY
Mvv80wJLdZByoWUKGCkggPk1w8SJP/Wf7y0hVUWPONJn9PZn7NJVW65Lde+k
t+KgWClYZmQcU0xbJqp2FPNh9xH0yuJ/tLAt2RbV21sEMyXIlnno9fFYg3H3
rZtPqE/gEDKoq9CsYQ7i0qyID6Tk5wdPlh/UIrRzzMxxLKsZOJFYzNN8Kxwq
yJwawMcyY5XmGxbJY7ONmVRqUqNg9Xr48yG6I/SxaRXs+BwdkV7BW03LVlrS
+0Gr+yHg+996/IsGULyjxKLFvC2Y4mPtWu8t9TZwQTsIZuz0dC3+aM17EEXp
XI/7TNOC8KK55KZ8PqEC3Vk+hVymsl1+GHOdHkPyhq8dq2LMQr78qcEP2ypt
mi+ZkDtiRZlwfThCQU9YI+tCyRC06OgdzxzQ2fg8nOjwaqUyyoIvEN0d6YDX
C4Hs3Vm4GBd2CkWLumq8qihHUz3XXUqdX9virs+bQsXE45NsciEM/EYIBuGx
hw+jytnaG8lTQO0LXw0j4K/yvf4piUeClrglRwlIRbyvbZ+3TZe1D5oeVer1
ooU/sHK+u32GyjK/Ivxti1PcFDiX995Y9S4xpphEvua0UxGaDAyxvkD7t/U6
CCoucSMSu6z6H2Tu/AkHws5H1D5at2fOBiLL0Wqt+GuL0JVJ3tuWppeFXuma
uGdUohjoQsNeUIdvgFgmubX0Bwi1X9QQfLz0sNmHkkRHmHmuaKH9TLG02KD7
RXapWOEeScUqDh1/vOv2fptn26BTDzlwPEF+zkr1nANizj6/r98zLmNU76tF
aGsrVAf1UfTQKB/uidsv5mV6poFAjplY9p5w4aHidVqZEf8ZDtuSJZxC5Nyz
/vYld3RS0GBfqH9Li3hG7sBmWncIrQIx0Ng8VZ2uBEnpCOwHnr6Lmya6whh4
uF8Ba4LrlA928q0nPpZbU26lMrZDuWpAnAl/nELaUT4e0+o/++96rPSDxOYL
zkWMrVMT8Hlbpj3jXU3SwDq2sK/v+ymQ1CUIjpekZ2hRXf2P040Zy8xlJ6T+
+7ylFeBAv1fiaubV37iN7N0NGrHn61a91TbnxB+GZDIWfDlyo59/IiznkAir
rbzjqv9w7FtcfUUKCJWpJSfGNKbwtQ/YqouhaaVAm8A3DxBGPiK40kbpSBoy
8oPhxKISJ5rOJIi/KanWTfvs3WUTJugatzQbT68oPdkB+hxVu4tKJ+mHgQGX
xoCKP8HbkajyI30KaklYAjBxkB9MK3CE+swAk3zd9n17AJhVku1TICqAAY1l
D+rD7aDGqiYI0Tqm712AbRx9GNEVycJiIUfZhXKBQCWDbNHfSPaxeGtsSbGI
8Z3D6RL7dib7bQR24ebUguZue/xVUPhDv8HHeiknb3VZy4s0CBJewJcBT0CJ
W2MuXH1+WpLS94vV9MvdKdtnbLbjIwfhGVayk2XdJBZ14KqXEui+LJGfAGGt
o79RtTIXkVtOqq3qAbXUq/433qARrurbV5ESsQRFHc1cKa2VETjmkfBAw03A
XV6LkPWMXFqkDv1uYUtk3KKp+4KQlRzzDHAhuYJArTXH8lrSCyOooI8dBgP9
ZuED8oqdBJ5YFEabaB7yF2NSmTe2jRv00GLDAQ0iDR9bIoF8wjtbqjRmZvZk
ZMiOQ7XcsGfbnQ8YlZ3zoTX5yCONC1EMxanemGiYholKbCkQBllMtA+PYWhS
tJOSwYJC6mT76iWCk9OqTl75EAWcqEK/1YbydrFJJhLFSd+rZ5ScrhcRkW5U
TnuTbuhImlqMlElzKE00B360Pw6kwDPilGCNGVYfTpFSrZj8Pd5YDIMxTaib
u4RsTqpgf3KMPTuiGRHgdvr2JnHGRR+N3L/Bn8IXKhbG+aMuwfCBpKJhtPOP
0x6kXMrHeszPAzyiaKRAqxI1nQ6DUSzL8JPz9j8J0tkLcDW20JRvyOYjqFy6
6sO3nxACbTJH2yr8HrdbtorOqIf/DPMS1Me7ikyKqR3XCRVUSpKPvJGDvN8X
DYRX4lIbIeKsadlOo0OKmtKRUMoqEWub3zwmAqFqeU0wkiuIZgjFboTtMWBw
Y72SZqEPej5/XcRltgWvNEQf6wnOXwIAlGSdHJPUa2PD9V74XPo8nk5itbfm
HY2mcNHkVERH4Q0+kcugEr95dS3p7QJfh/NG6Dk/txn0faU/3/V9HAelHMBg
fyDLTDwJH/FIQ8ntRBvehYMaCBeq0lnKu1Ql3RJzcdqiOuunqY0dO7VbEQv6
hzTcOuVqvSA8jh4efF+0e5xJBiRdv2P7Nb5aO/e8F95pxQ4v6G4oKwxRegSQ
/7Lv4kGdbiCsOUTf+O7RCpFyLj2yuVou8Ex5xJ/JE6jn1mLkvas0YSnmkrko
+n4hiZTfCFmcKllTxJKsSmEumMRUAP7sCbqagY1Tu+7Af8jntchd98HsUR73
Ndv+iatxEgBpQWsO+Tm2MVRiA24YPFb5uHA8liyDB6raC2zinIdsxYRkDv01
e5Ze4ij59RscgXzX8LDJCW0cAdK34XHZijMU0bu1ZGKkvRi8WumN66IqCajJ
Vfbhw/hREw6B8MPEThJ69iQWDqY79QgZl0vbEdpc0QBkgIprB0mZwGgAwLR6
BC+fFQpxDNtyqBeX8FlaXTrlD8nNCGUZEhPgAgEC4kEGbTXhOhtwQ1Xbaw2B
SugrQE77sYVQ1doHLpZRscxlmQnM4QH8n6PXMVxqUz/bBXbCltyPdVY54+Ue
05P5my6jxU/RFppl6N9VaTBw2dHfa60PZDEmeRVCx5X+dt+XHNnuAxNgYYNU
EDKnzGYr+PqTAiBZfwlc/zIFaVfrrPYAp2/jmCBN6N6H5uTq/AdCkR4x1OOM
1somZ0MNz2Lo3l1wb2wRHmhES7DcvL97qS9qzNg6JBl0H6Fe1ZRTrZwg8dSn
Xyh2gw+4iNhmqGnxgscz1IMQCoQku2+8Z9AR/r5MILaeuvykR4Ef6CXlvVsv
C5Fu0gQdOI0yY5DHdHyl+3XH+jj0sTAnXCqkXEe2FrC3Jyor1V96rXZkZQLl
1m7F40szWI6dVMTJxlRT2Z9dE2x3Qp3FxHvuOI2Hh1XQr2f0rVK/zHrYehZi
jrsfrOjKPgJH1NjkY/y6TrSIcKzj3/VcVe+Su4h+7rU5odXYPY+A6fgFON9/
SFG92u7+RFu4CvspABcq/nEGvup4OAWu9BERg9n8b4w5JwpHSedtTdjsFUT/
VwPnBxnudKqt5ZhwoZKEwpg1KWIQGRygiy8qceMLEZkD/CPcj7im3pavKD3i
EwZt1hmdNv7ttEpwOI8mEbfWNAN7LDjcRE+eys6vWAkUfuD2eK4vwMM72VdG
pmB/ckjojsDdBy8emtUX0/U3dDrth1Nd0aa7wGeBuwVstX1UeGSfa1trKZFX
/vEjiWdZzkIOSveIqdhaKc51kjlyqi9oolodvJnBJPY6jbdHVjbEa7pAu+6P
wgBi1SEC+xQ4OTVf8Lw0MMbNIiTn/eNndhViLluOfeJIbW4hipQ8tJYKV+vY
B4AIUpEAaXRRHauMLOvr9iQ7BXUU8PEx7eBtuyD6vDdmxxcdxXi5Emo6Vij0
qnSxTAmITYi6OuCUIpIbtWv1AnvIZQq595FeRV/MeS7JZZlUPIda847kG3BQ
XyoZ///EIOwf/L4g3+x+n60CTMqHDCUzmYfrdreG32jzGKOfWdfc+DO5zVPU
KWss4WiwLuEP5jARrZxbJkReEOdooV0nLg/twYi+hoY/MJ2ImaexLJ0w/3rb
mBgX2FYXVLNJM+QSu/LyabNtlp1rhP/sLU7vozsatqYI89llZ1nwQGfDXV24
9IiXFjWSdi4QDcb1rer3uJoNDOCKuq3OzJZ6kPKD/5qcjlZxkuXBmS33ZIkP
CoVyc+HHVPF92Pq9snKpSJ9Ot1U9r3PiF5nwBb0XoPsqWh6AOQghFSXcoqsR
HOYol9yEyXHmJgyGUnkIzRWIj7cIkBfxXhtFidQ/z+nfQBZhHpvPTIeGou5Y
blXieOx+vZo7jO0TIrRJvPFgy109GpbnL0h4WQtI8tp5TueUC/O+dcIrNSGc
z5UafFCRT6jvHHWNftEAQo92oKvU8zWS+9rdAKUYdJwm2WwM9TInk16OS84h
uhbp+J0fEurCNST3gjs55hJb//ixIf22P7a1jLjMc92+IhWUgfblxEfIHtUC
AESEgf8146AfSw+Ox/OM8JJ4UkDubcooMSYS9MVgMYGrdO4IpbXmHQ44n1f6
lBUjMpYxI06tgF8e45vgNDKEpc0GwY16qKJLlzVFe/NqccRoQwojAc4Q0vgJ
iwgF3yMVkEbqAVlXwGlTbe/+ggGN8le+0RH9E/eUxMdICt0QFLGK7k/BcHI1
OfSQ9GXpH1UPlO83SSRRwrtOG7mTWbNpjooHcYjb8hOksP2VgdwfdDh4A1uY
duddbW0trvKmiZ8r2A0BRnyhHMEuX6bSFhYzDSs/OqL3J3TkQCv+5VcfTFnQ
wcl5jR5Lp3i4zphWAcoHNI/w0oqniSAXVsYh8tj/aisKSYTiJtLdpYk6jMGF
WjedA+jls7wmI3FgkgQuBjckrybB6emzaWatSYoILMBxoxTqLK/AzBMJUJQl
pT7kNhFcS8/ULNqYumAerCnQIlua5Y7gAJ0CcZEhFyo7yhFyN7XrHAmzt1zz
LpjufoOvSG3bQHRMW8acTNcT7zi9HzJKBOGYnr4P1bEb7c1S8Oxjz8Y2L62I
r+o+rQN3muTpJVJOkHwSGQXl6uIODmGxWohop3Cr7cYiCVdzt7+XnohJJ5v3
Z8byO0mK8yHozdSih3pK8gJkTRV5iVbO99hTkaInjpU5oLTWmRMeNat8p3cF
rnSQaeVL4MwElgXB8W5AX5eZkILSfwTbLQf+Uksil5BL4htiU+Bhk2zI9k69
8rnTuqBByETb/xbWSGXLuNSm6V+UVRjnB2dm1g1boS5HAIQ93jYYZBuB0nry
Wov7EtJH4jBvFFJfgLvl9c3IdGG+2a1xE6fzzuHv+INx6nL4OTnlbWaCbQtn
E7XWw32wXPSueXjrOJBF8S6hIgc255+5rXx0eRS/hedoGnQqt1EH2MJT7EKQ
gHUcGfp+IWuIwVh3q2/u8EE++ibWDVKp8c/e1I3mEtDZi5Y36vHGDjX4kpJ5
K0+5DGvi7L3cw5Vea6PfKgzGn4WGiCAy8xTG3sar+vdObIwOPx+Peo38yNgb
2krWoMfur0PkIqshb8hNc7UU7ytt/clzXimCqkSwgWOOa9dNXs349KXSyf82
rPnE+nNE/A7lrZufKk4nLIMkEFPAx6T5Yuq6XZQDGD5OIctE2OYc0b6LTZah
spZIq4q65TmgvHMebctxpLy4jPdVC0EvvAiLg5Qd7+QxBu0hca3S2018paNQ
Pc+/93fZrHsQ6LAGRBywEsy7IXQodrQDgrq0QVnfVNTUd8VHLlyBsO3nm02z
evVJfLzg2N0X3R/xTIjMQpwMhz7korpMYcrofsYo3lpPf1E2rqlSXzauNFsm
9kfT9oxwWOR+x7CSDDgdFnVAH1k0ZttNZM+MIDrVugd6No2p2HF00rf41gc7
THnV5r4HZHJgpGWKfvb8vdt/pc9VyjalKjMeF5gzgKHzr+6NEAhplSQesoO/
2egvyyFyBkGIHTcHbxy65Tx0sw081/xYnb4y0MkpZvH4EKunGbwUvKlt9lcr
nivUuoKOb6ERvOzK00EBgXFa7AqDjuwA5cmWREjOmVenv8bLeYQd2jVQdv68
xcFmF3KFc8tQ5RjcMNCiwedlQRkSTv+ZYzhAvHuxKdcgvQqidrQR5L9OyEDU
ipMcLRjF8qs1D1hCpNpIu3/t6Sxhtp02/94FFbPTAtygsDLF2/5RsKucNucy
b9fNGFsPJFrbxVHm4xwZ8bsv0qwzCtNP8ZxmF6HcR7FV9IWxH8KLdKDM2wvJ
unl+QD3eucQRmZCQfoTDlJFEJncCK9Bi+Vo0UnGEyZqgGROGAHLaMlj2G+iV
oivfaZR06yeZqXZCv84vaWWlWP/kTAXjp9L/zddXg9VFKFH/6Xm2np3PxkH3
ilpwgTW6wkYeG8Elaf1xPONoFEuYCVmj/+Ti5JJlyOUf4KUviUkgwYDrSHKi
ZAH8TCFTptDg1L0ZXghuWZ90OClzFhC3rOYBRKOpCTSkKkhNoO5Oja52J1nI
BGvvA8IAATkK2CMkCWx01xVCpf32qhl3PdODsSBPt0LFzucSoSuFhn6mHB1W
2HvyW0mbBVM8oQtrBQTRYnkBfWPdhS+qiaHv3+0RPXpOGubZSUQeaINF7oa/
enjGzwxAMsktwK6oDe3DEYFhuSa/Kmij7mF+c2u1FJKJ/cIq7B0uz2UNC65t
39qS3D6+/oSv4SP/AJxc1NykWn4t23HU3Jc9FTagiAQE+xPlU0zlGlT9Qc+q
RvFW+lczmlCu0maq0kUnsi2GM+raS81HRJGx50R7NpsJpTJkB8nq7j/e/VvJ
7Z6wMgT41AZrIcaQGwzluJfkOcQeF9q6juvWB3T7dAfvR4dS0o4Iyy17emkR
SMwJsEc2ce1Wgovvb583rL9DuqaqHHUi7XWv8PxMYIVUG4thpF5dBPaUuSzH
lPrKCVTj9zvCSa0qdPowTb8JNtpnVd4AY1DZ1FEBopdeotdb7QicFwh5PFWY
PtyQmiUquWcxVxPnJgyf+U1Fp4b/HTYvl1ZQ1Z5If+qt7oHSqJCQYnnqf3kh
1VI/NzCmVggPmoRGhmEUeYuV58vJYbatIDG2Y9KtGDe5/KQUmRdKlsAbdKKm
+5HfWgi0/vdG+H4XgQK8ty2aYQLqRZHOEAzfy1qvN/JWHf0QfkLhpuBzvE4L
WCDP/Y3AuJKhBb4zLN2IlrnRJNHiosxSsItt6dW+jmbRONO+JRRUZS/5K4nD
8eRt6lCiHUioKbFgRzPt6Z3YUAxUjwXptMdi8PSQRAQxNj0qSA3iNo49+64C
5u+vLVvjjC/Y4SNhjh1oIyYaSTkVsdPa3EQBeNsVyyug5o+qfpRUj63k0JiK
gc6hhpkFQdC0ANLMLVTS0eOxVDqyGHSDAadyyYMovdkH5kKnZt1GdNQA/53t
ogybGLbprRgEW2bxsNQmdhv1IKgqTkCB/Dcdy0cCAIajtEYlKvTpdmX2Yu5q
LbgmboTyY2+/DxNckdFTwyiCrMSIpXNMT9ogqK1SpARwAemvoNnKGPAajnTb
7O4p5GiwfpUu0LhJcQGJbLzorhux4zSjX1QS6+YVN1oqx05lhlnrldXVlZ9U
3lEk6DGAy4QDyWOR051vy7dQk6DpZ4wDoHLezi+iPssCa5RMKdpYke3HdCMF
allOGCMQ00FaGZ2wR1w/ngeD5mHUf3G0YqVowIHPBt/S8hOoJmXCmnoKCbnx
mH70AhijQFwBa3k+rTHGb41mqNh5nk5pgLw4gvlTLTmm2i6i6b6Xt3zVdf+i
HOvMBrY/a63G8ZUYlJRENafSksxJDqTpvirLsTMu3njkfjIQL3FsHZ5D8Buo
8zhvX+MbHQhUedXznC4R5cVXxJsNoZdM0Btek1aB8NKcyPWTt3tfE5NxX0u9
+VD2c2bswdW6XdPRbXG6lY3/mrYTFxp/VAnbWs8yUyGCc6IjKF4xG+rTLcEp
WdesSqUb2EkXKdQegO2XeCZ+WhpngYtdaiJ1fcF02ofuQAoXrZOtg2Mc18Ke
ypAhP9yNLsSnqQ6iaW+V2e7mUXEoBzQfuRUTgnygWtxVTv1plN6HUeDsMPjy
9HTycAFzS5Wit8Km+LEMTm/zuFhFyqO7h7T1Wpii42KjoP4GVeV5iMr83E1+
IHxwIA7HqyB+2OKa811e+QRXJvIXZNPQ4msQD1elnvCs0U5IoFsbKQzw36Me
yOoxrsWmSi1luBFutcBZOdcaBPuHnjfFirKXdKWo4Z6vyUjrGe1BrJnPAQAD
ZzWP6/aidk26E9c1nQwP3gSMv90wyFAfiEQEoFDsaEuRznALPKzy+fSEcGWd
VORuROYq/SDGmcshJM2srmnConCE+FEDPC4kAzpnCMpGRQxq1dy0eCXfboTs
CRslEeNfkB41JvGxEVt0CiJxHsjObnCfptYnfa24tKoZO02bOK0y43t8F7nJ
6VFowx0YM4vPZZ/JNGDu/t13r0Q3s/6unTilm8B7RZ5cCu8m68rAG/RiJFv/
gD4MsPEHntSr71ySmA6mdNdTltllL6DQSQLk3c/qoiRWpHPFnWz7AgnhQY/E
/MdQ6agQ6vzUtpM2nbaVm8TvwQXNkRDzM7SXDHvpXvD8D71umPNbzX9BcfrT
ja3+/Z5N8uvU/X5bolOLck1DU5S+0N7zf04eLzSW122Laq5/p1BDHKoTnK8B
s+5pnhbPAdmI4W8VDN674OPxNDjbxDLrRrBFgSIt4e7N1IUtiBVxsf5BCqmM
u4XkpP2V03nOGcrZ6hjc1FxrLYJaz/KTwMa7haIL2+XevjOruh6ATBe5W5nd
lfgRldPlkwS+xBe/JsfW2rkjX1d7IyaIxt+ouvYHS2zGJS8zrG+h1UlHGFx+
mGfMNz1HFG2fhZvLmPzW5TSsn1e2DURpJnzYIvelXEijFIqTu29NgCJU0E/w
9w5RTfaQWd1RBvzG5dNEjq9YFAmZKMIY+L0LiWxAiDijrBosSNnbv+KFrp4M
ZwkAr+IAwIuIEay+Sh4JFy2ZgMUZrgg1hadlBT6BQP/ealjQUZSE/5HysoXO
YKvNBnoxkooTNsq7NEus0jl7F+qmVwkkYP4kGPjt5QtEzrFQgMqEmzMJ6S1R
ztUbxxujzMzCMImU9BFG18we3NFrJeZuRZEVfV8QgRYgfWwP2Q3f0o8/v3KK
wVrQpfEkFjOcEOQ6tRtqg60Srl5mKOav8ZyWiutI48+o1rAPl20c3HLW7x5p
Yftof0ifIHzjZpPQ5xl8xFmd0HnONhlDWvKC9DTmtWRwUO0Gz3WMT2qTgQwH
mM/FovzwyQl35hGTAvcshfxxzWGTObBcsTQgQwEBNyfY192r98UGsipOaRE1
AxebLvLKkWWgF2yi4ESVDddPP/9sY1r3z0fKvLT4Us0RNVFtK1VeOhZkIKmu
Ab28FVmAJbTcCI6MdJVAe+EbuZRYlN7hoyVtYFBifrSo9fGbJQn0mWfrOH/m
ONCxjolEiy+gTEpqTypqFj/fsPQzOFmmwRmBjoYx45rV7XhS/dNdg6fQT6x4
02KQROxVbALmkKs0yh/rdztz0LiCTgCZURrK9HbmIKJ19LFvw4WEDiDWBTqK
SKWZVhGkDxDGlqgmG8IeNcdhalqFyVncfJKgyLx2Tvx1BYzQsQ/axz6M18YO
ZGc5qDqNCqWnLqvPAe+9J2P6FXTA0WOaCxFbpgs1hcfpk2PE5eNWezwL8nPt
ip43fOUtABZpoQLWW15ywppZFkOrtKlj6Oe6K6sdqgv+YRmw1Z+kGlkI3npF
FheKqKck+llupot5fML6cOGl7swwOt1yliPoYPKqY1TRyctG7b7PsiZlB+rj
HE7Js+GrrY1QT3+4dN3NHaHmWUvOuApiL5hE7X/0AWapiRJUyYVefM6pHZyU
eXdx9ef7v7jidvlIIuxWTgCB8Zs7JhiuDQPcP1M+tlJroi3TDDg4EVB8f750
eC78LKd9S9eRQ1g4PZUUlZY7JDWU7o7rkmSsS3546w6nOeYUIYQz8jwIJliR
xhqtQB0qent3R1aNBmdsv05qXGOJR/vra5cdWenC5QjRfZLipWM/q8BpvAak
dVXUaP14+Vb9AM58OANq+5x0+O7UAkK+7FPbg7Qe0B0VJMPbU22RP1P/QpH5
RL4XALj0KyU7cZVdXf+tr4Cny1frTUukzuuziF/M2xZO0HunVAMwYtsAgPRV
8A+7/rKvDmgnMPP/lQGMGbTgx4oRfKRB0KWBujb/E7U5E3Gng0JGnOS6/qeN
b0OviD+jsNHgBAZs+/y1izd/lsrnanpm36TchiR2f4C3r8wxDE9ZR1eZql3v
ETha7+okXSfqDTct1RYoU4OewZYwD/ef5zeDURNjnNGtFBaCHXck89++Zt9V
7mmYIVzRCYvpcZYkh3WxqtrAcsOgOVY8te7wGOT1X9EMS5dx55boKZoGX3Br
6ZIBKN670k5avY53ozCP+3DRh2uz2EiFJF+p7shW0g+ypNvv+Wp5H+rB8y9U
W4WGV75gP6wtGoXSwe4BiWDHF9mSX3D5fowll4LRPNIWT2jSqsIpQnhPLUjr
qRmAEdoOkLWmnWzhcqQ93EsBbEY8JTinplfNMgkYsnZreI1z7R6sq57/UMHJ
vdESyakqBBHl/zLzTjTPKEVoJCD9WBLnPkTSR73uISyNfCT2byypDbUA87AM
7ULILBQMdEYRe13y6Sqa342qLKx0760H87SY43RIXofo/Z71kNAqo0AM7H4k
pMYwQfsMVPF3zAq7+HcNn0uY4xVBKYo9FnCiWXh/RdQ4VqlLD7xU+jdLorzC
QW1+7GGoAaHDQDiDJf1GBBgNw/N2sFolETS7XEySR34d8dR1i8Q/vZmhiLLR
an76aaR8yQma6StGbBsKakHK33/NUDipPV8DH/Bov0zJ145+SJBZzr5+/pTS
W/JayCBHIpGJOCfeCyLoYsiNUpgrYbXRUSG17Lg8XKUVFSSlAQfz6h5aLVft
6siOO6wVTz+qkODg8DbiJfGFMBDA/4L/oJhX2sNCL/nZaUkaXS2JHTs9OIWr
EGq8VF4+2cqCV+qgGDsCqhxLW0GfkMk291KfwDtLXUmG7kusBs+TCkLGS8vK
bBQL4uUeKoFd3JDQ/Gsd6OSL6KLe54rxaq8/glE9WcHYNm58WPIf5v0M/XmZ
fXVorqEFzWjeN8sEHUBW/wOOwaFPWFP9q8lB2hcC0yRgtcJYTKRacBsSgt7i
BGIyz9JIdKYQ8NtY8+1kbkUMupg1UV8nxn5Fis8vNfM3eYwIbmepvIh45Q/W
j9Jyazr0fxT+vaTOOmyu3qJxmlB5ZUnS38ySuUXlm3BKal4fGC2PAoLzEx/s
Ae8yXM18TrfGosPWMB+obp2NVOtTaXfOqN3yMxEfl9KO/w0Fvx18l9OrN6CI
qRRZowsp6h+thF5q6Yztpa+dfg9wxLvY3M1LiTnxac3AdZ6Jv1nOavGR42mj
p5Cb6dJpQYPI95k/5VW6+R0dCHeajrCpyYzbh2afKefJTfb9NR7sANJZljEr
htlOmWFtgxRYZE/AEGHFaOcipm/1+VxeMsyLffP30HmDlnh6xS7QchDpaPpH
jmhfWMdlwuMRa3z4MfXZgSL37+XiCDDCJS3qYG95a9TT2R6SHRC4kxiF34if
ey3pewHWIxuJlw7rox7uSD9ZBht2bqeD4Fcz1qrCSktBN3a87KI47W2p/n3K
F4koOgrPnhJy8OxMHZBSd6y/MmYQyQWFZoxJz3luEYUgmQcLI3hBLbPr20f9
PDJup0zI5XnBWYXv6gnfBPAl3o+U5m+lJ3dQGYf2A+O5FMStxsAwL0RNotvP
D7b4XJLe7GrqtCPaX/AGTMICqzj4z5HGbaychi1sxMV8C+xo1IbjLwnp/iTP
t7PyD2J/4kRFLjpIU9qp52vdmhHzNAela5JRjHdX9wGWn0zHoKotWdN64Rp7
H0ykp3BbcmnHaegAbGi0/PfuAjqztqPniyX2aZ0ulfDQZubn7RpqKF5LJajv
B6D5U6rDGBchg8+n4XwvYOfPIN0Hh4fe14Eoy9/zajcRFTr13+Es2LIwi4QI
2EPQBbstSb6l9+69wgcYHMo0ABJoFDpAbGH9j/BdoQVFQmKS/a6sTyHN5Hri
BXvIIVecculYHLf5qBt30bXbeZbBuTu6vVVmuPRxfBADkJKo4xg8xO47x+Gr
FmpqhIAJ4Ah0YkxwdtfpiC9LTZ54yMNmKXdNZ3qkPDfAng3wpP/gNm/RAa1W
cu1+GxwvQp0yydj/iojskh6rXNpjJwG0LCusW/e1RS6yVwh35rXSD6qwvAGb
QBA5ES4Gj8ulVmMV3KhGupQFC8oPbLYVT/vOjP78SydR/7vVsbA/RjDOiD6k
ESpVrJ70QQPP+lNHDXYh3pf3i2sJmU2DdfTMwZQx1VoqgDLejdZHBXsNK9+K
8azrIQwm04eBWznqZdJMKDdq6IJP16zUV3B0PoUtMH1TR70LTFoTV6zlvtew
vlD2gXhheb4FuEkXlD+EmNFm8wCEmVHBnQ5K5+UWrMhOsJqvT+28chaH3kpC
B+D+EoMiy0rT6eTSPpRI1Z1VXiJzpESATz5nGesbb02q07BTK6AL65WBxCn7
LfGeyEAkhQMsMKkOD2lFwaoW4ZnJYCBPjc/kDUfMPkmTIlyIurRSqVgFZLhu
4g+AEDwiUlYgPrkyB1hwIHPJWvhsGu2FzNFUcjDEZ9arRKNY+Ix4s5B77RVS
mepIcf/YyTBaGfu2S5Km5X6NbL5ks54T4SMklvGyAUUijXpuqB2rik45+LQ4
WyU/dF1HpX8/XE6hR9ZM/Y1CFPtHEaYF2S+wqSjY8Cf/BNrUcWCrnSTCH0gq
FKL+exJN2ROKqKsivQIFUnGs9qriV4FyU+EynDW3GBNDFr8A40i5Cc+SHcrR
mAqPylxmgH9+U32B75+oWnqgj685ZKDzi3ZJxl7dpe/IvDv6zA82jeKzwqIf
dWGcxr2uY3Fn3at3SIsqM+MCFqHFBxUEst5loTwy58sj3HQIHTpSOi51Rgq2
a9l/hHdDWx2nuqqw6IflcF+IK5P2XVMIMUk6EdvC7HCZ2IToiXZ5schXVVdZ
fsHbMlxFzgWNOhsDBRDVWSCI0YNbPKFNV3ZYp8wXrlbFyQ661uvY3C060ocY
+CEo85yD2W6+PJC1482cwK5T6WF8eULs1YJ++DCHvxG6aljldzml1HA+YsCb
IfGT7uSmSmyQ0uEOMaF9RL1jYj04gtKf7qbc4jXHoTWBNyteC3NXuCJn1FxA
8P+B/0a0Wp8zXNd/Sg3mUvAA42UL8f9ctSxGLgK8FYjCFeZvYcMHyj3RzEoK
bMUfb97LakLemhvejlwhPKihMltIrW708eNqkMOgWZF+IivA7Z0QGDTN6GQQ
ApavruhB7k2uCzc0n2qVRDPqsvFznnGqKXrzQ/LOUNUlF+DukvFR38noUXTw
71kFMfpmzWEY4AkMVkgicekhFBkKPeqr6SMl6KkD1NQdjOj+qRhbw/2PQ6Sa
lwpajGbdW+4vGYcO3JAT/GzVMZeJHLwKU/69NEl/dLqjiHlKcZTjpRGNEwAW
+7EIRn5ygNikQwIs9RCWuBQqABk5n1zF421Fn0fVMML1k23NWNQi8hBxJFHg
F3Ne3KJqi9kmp6Kuw7V2eWtMr4PMpWqL2+bQyxBzlqyRCR9YmCaD63suhXY2
pjbD0Kf/JfBjGYnjLFeyLnXDr3kRQn5aOMYbiwROpAsc1NLwEhCZrdTxMA7Z
ho7pqygKTQAw+++YSaSgeB0srotZVkcNEyFZXZuykJbhPXglSPHmSU6RrY6a
j/XA3aWfQ01qDnpaJ8RI5KMBr+/Sro+iBdwIs84QrtUBDB2x/bI71Jk56Czx
IfV9fjtti/WEbQ21NDBRamk71C/R6+Bp14a4wXOjDp94uIzSBOCTI0XUjUgN
fq/z/RUsjYk81FclOUQLW7y6oyhu9qw4ownCsLXPsEfHcQhqp6cAILYZKtlG
/eSx6VH3nXdTJmhpnp2gxhOse6rndKL0kWfzA5FNenjXEJXhWFvlKNeuNDcr
NnoP0Kh+z8bDyWGrQZ91dviJlCFC/MxLeWCprK42UOE8jpm8BDCKlGSqqlnE
kUczmqJPwJImoXnRSg+1bdN+J56WN5t1wZqOEBetLHWdny3q7uhOrfV77MHh
aNByoLHDMIDcAnzZ3Lq4Y8Mrp08iCPjymEm6kecmYMRU27Ix8fR9N1LP3G3v
Z/vAJUBmNI5BmrZgSmOaJq+CuNBZnAamUsuicjXz5nNV9SrD9naFEZ1RWXMp
IzTw0u1kVSJkVdKp9SLKOBDxGVybo34YMrKDUHxtNSdQjD7674Lu9VijBdyY
xVOJvASlOqi+ZexHWEw0KNq08btwy8Hh0SLKUd1AZhugo59mdwL1qnF+6odc
vpBDz9MsvjutmH3E6E3ZHw91ZMcvt1xgtVwPVWvlFUmLKj03u3nQcSUzzaRd
5Gvq5nJuLDa4sOiPjo02/3begNfYaNzXhfhXMpMDFP97CbY1yEiW9ndQrWPG
bKuxpCtc4DnihSROjYN3nxuXfsD/X/3Gj96+2lNU/geVK4QAqXn1msS5SIDG
6V06D3IqBaJEhwUJ2JgquogDnOm32NGmSf3S5GQlQQfD7N+QDCCm2j6P5EP8
xf0UTOgFfXnNs8mM2YFU8g76y11/bdITu2WEcHzHz4Ry7SbwRMRhCu6pvsUP
WQyyu7n6ExBSwWDaW/SWB8FOwvAbn6P0i1G7quelOuNOD+p8CNRxnpK9dmLS
r1VPxvl0ATT1uxX+Tc1UhLFynhOPfuiPL8FGbEIwynbg7OIZbrgK6MfMbQ8j
4ZtQZWveMUDuaDGoGCVbIOKjTgN2SDxcM77fXUwnKBCJ+dVWZxeH4SVYMXcr
9Z2pt8U7TzJe2iXiSVvKotDEqFhp4WXAOzNU/QezPHR9wE+SE6Kq0BQPrTTQ
pqfSba43c1GKPqe+H1WGo5l0m9LTs+1BXlgY5oxP9IJT3XKZ8nIZUyutWx0x
Q2YSFbEbJzjXp2QEdQ1rsCHEW5WxpNxEjpaDcGS115zJO1s5iQOMNKGlKGlA
sODyqQJqBcetI0fZMkASIVLQjpCwG77Yb0AjkJZky0r4/6T3ACdSveMqVead
PnvppiLlLanuUjK7x/NjnKUSKBLCOk+o7oiCRzaRosNzF+pk7CPqCm9wugyS
ZTj/7FBktAyAV7fMM8S7FFKvzfq6+gYKkKDPQfq5SjetnD7JAyBBlbKdUGm7
i++vFuHiL47UFYpbXrYXmrY/tXSaNSfo6XTJjUPVNdUNOjjOb2OYgxXwDKBA
AhSNfqV4gzRYLmQhJw2dYYUBCY3+tb+f8XffXRUiHiFD7JvoUJairG5JWOV1
fcECqMxPgZUCATTWjKw5InpLTXs0sryxFOeqsk3Oh23o3NZqucUhFjeerAZM
q58GKZMsAaK+cj9YT3xSNNtZl3mWmzmMVaJc1uSUT/DbMJM158gx6FO850y5
IfF8ld4VBcbfb2HAq/u6ZYyJLKyjh1g/t1upmtKVx4yIE46BIGhxLHNh46xR
Vt4Z43o1/CicIZFFxbt4HH7ocaXJ/qjqU8K//fInDT1ITWsNzkFCWZrSMOPK
DSGn2ZmPkFV2zJ+nx3Mvd4U4cPQOBgbH9rQ+LHdXs/uq2KSVEZ7AfMvvMf+s
pHGx3/AOtAScOiGqwbSylsR7H8G2CuRJHHoyEup8vygn0oL1x6xuQD9uo8kT
r3Y24sDqxYfHJd9R0ga6l0XZ1n8pswUWdpv7Zd5qOg14AERZOjaGMciBIOIs
CnYEiwbV07hb9sFZIyoEktVugj2P8WrYfdq54b/mWaEK3j9kGMlMHSKvEdDI
cAxnwxuDe6SA0YGr13DdwgreNDyk2JkeRlx45xDgRbtsiPdBhs+MI0QDlhKU
KolX1LDL9c8BnmFnfGugbZtXUUB0th/BmzHpFP85/2nf2Uhrz0Ogjcm+ZIav
1bMIhsbdx5m+oqZTKKE6IecG/NVG0NWTz8OQsaeDkSm3C7PsHxmFOFPbEq0J
GXd0ff66flrakOVZJf5soxCI4VqkQnKTOhbwOza3XRWc02z1uwra99bDvSr0
oKlnJ5pyEcR84rDjyvmQJk0zD8CV72CLRXnIFouSFnKoGIkAI32zRVJ8RyE9
xWQD19iInKhRzwraZVctbxTrzHLGNXW7yO2A1hDPyNUHgjnSNgHfDmiEW56w
f/4MKZFYPpL0NJE2Vh3U7W2WcEW0foZ+nnUE6PB3RWLW31kkK1nlxarsaVBU
NubCRLFnaFVQAs8L8lqbKv7JxHQhAOInI4g2dCcNzt5K27QFvin/Ofkh8XUm
sQvL8srw2wXGMOUF/pL3cwRBeGL81Z3biIas57qIQ7Xc4OVG2XaFPKjDw1tK
J1ku12Wzz5jG3K7ahF2p3PDhZYiFZ8lIwF1ncn3cbz9FgCid3TMl34fV2EvT
nz67SDPtwem5KGc3A5jCzZPZJUPIC2d1onyHZxvYwCNYTebn4jbCFkAQmD/T
63KVcPDlCAgxCzXeOWb0c3nXivu3uqYdSrqSfcPBtVkE8JXM8v8n7Y8d2k9L
rCUg6kHaXMrzVK+j/zpfLpD7MqqC0sfkjx1ZiBbAAiOyxoJh6TQ7PlUIPP4G
hIFsHeOiI6X9NpB7vTuth8bUEotJ2El/PYrD3ZKDpjKOt4njLsqayORYHpBZ
qHNcB3F79G+wQrTKjvUKXQp5C3JlbpyfFH3MhcCQ3o0PC7KOkVsooQ/KM9oG
tAsqZZWoDldlr4F5ZtCmsAxKcw/1rPZlcm+Z2fNcuR+DP0Rf2o7oN/S9yaJe
+occwPvDFeIcvEc/6tP5WDhmS7EEm4JvYQIr1elk5q4Sth0wtfwpdR5Mtv6F
TbhWEAekUGV0wzOJkFlD0pjK4XPHGUDMvlKefaeM3dJw8FnFvnB3+ZZS8dcP
8yvB3/HB+5gprXm5bnXb4jvJMawxgcQBW469YMKuimuGX6tsSDqbXBvcZ9q7
7nMRP3KMFVxt8bBZtwDEfGe1KMMFS3wzwJbDIBx63l/fGkHWh2qSmAF6NnUi
5nRJ3mfoEc0J1kK1YaHf0ba51SNObFLN8P1HfN/imVSP/xNgX3jWZSs73KTp
YO6JQcAV7rl8UOY8Yco8eFZQ0aCMxi8wbIcyynWLx1ZK6q/vZFkTrQ5+U7+L
og4XxLxcTCI/7fSBeN8jlOzL6crNndDFmjT4ru3JTdXfNWYWEaTlReKvmuHf
v+jUrU2mIdxjQaF6qaxAqTnJhjepNw9HghVyf1cA6k3+tIVgMSzrz3i2HGPW
FBbFRiMvSpVNN8bPd2ujICgzSPxVul+TNfEPoQowB82jRz+BaWq+PRIAPAXJ
vDMDmuWT6IBBwN3LcVOi+HfGwkGxs/S6hMJAAJztPz7o/LwfpjJcPBe9E3Wy
D/gUVX3vkYFm8e/14K4/U/L+hUIlDblTbV4bID89J3EqTNWGrzRCt8MtWfCG
oKS/GzAcIwY8Nx79iUluPQXTjqs4QngzfBEt4FW42uNshKlGdZ+kxJa9iEns
vdd7hT6ACmmDwWEhi8GR4YSlJf7sNWUqLcUBAUxekxzzF6yy4IE4wPXcPcfz
cuw2LrZKEWeUvQLxA0tJWufi1zSTeAlDu9VORzuS3ABpQOLy60js0rUfPk16
b6AW11VM0AXeCZZOmTAr8pWOP9tvetunIvPyY/Jv1zLfGWmyxddTZZCiRdDW
YTgS+O05mcP+V56gZGoVUjf8AlwkcD3OvzJP9u8P2G/nsXRta/akFMcjcfsD
qYLSVTRUmVrJJMFr4f0Q6FHFt60jmOOxZc84+/xirQedO/i1ebItSTI4K6kT
U3Nvn68LwFYNC7t21GSEGTpIAfzHZjqNC+3SmmJ63y6n2VeytI96O4m8vC96
n64QWFuwG35KCr1+eTASHmhp/+C+XNjxMna50Q2s8HhwH41r7c1IZA5CRmCw
mBbtZI9jnHkaaF1dMwOPn1fd0mXu6RJO9mU5rSZhXNXkUUBorRgdMTyu4QLU
YMt004YP8NW78ZB8U1lb1rkwwPwWM4lAvlr70eYxmd4lWXwlZxXy5J+BAo/A
PK0DBv/5oJBwqlly+XmejG8siOc6jOabKGK+akZ7k/AWo4u5APXMTnzKnTFA
oMBK3NwAd/+kzIwvNb17rfO3D6/8MyL6wg+jSQwVe0CiI/dYaP8PX0khVOIj
NB8Ms3UKYZiMxdGXBOXAR5+1QGN4vOxV5Qw5cq72VwULp+YI93RaPm3VvEmD
I5qOHjW+nm4rBxpSwDRSeTFluckcDHShzAuz7GUdaVVFlX9Ez5MR/mjGb0M+
o9Vd46xI9tuyhpMI5pVj3NnRiglRiPzy9ATyJd9sB2SFEQpkgmgA+Vfzl+kW
gHyQHl0HONZWnZHfmmE3iDAUy9XKCZCrgytfGX6/V2C2z5BrBdv3MRyxDtNI
kKZHxL53yIEiq8J1fFM4CDVEdIAcK4CxqyCfDu+AMvdUBBSryb3OHoO9C6Vc
RxTMtK16C7GVOKGayJ/a+B1i1zr+vmKtq4gaggTJpI651d6g5f0QxAZSu0uF
r+uOpCT72fYdkaf+uEimhhJbyy9R+AZrOK7kRTLc7rJeh5+AalihPfHjEqN0
GmWO6rtsGASJN+XNW5EfaC95qTndlrFtEw/t7z695D73A7doPvbwJs46WPzs
/UeRmTRBOwP1EiKPQc1MVV4NayDT8vMhRab/5zsv55NZPcvhne9RV9z3GGP9
qlElDZMqcbDVXhcH/u2awlppCwivGV54gMhJucHUsliWcdhar6EhZuAssVpQ
7nvtJ9fvjBHs4Ex8XltU/RZxQszb8c4UAJPV88w/toKuvG4ydSUFh4sZa8Ex
oNpF8QJhJyEGtXR5ecoeW5tSGwnjJPSUGFe748X2n+UA7Fj3RRQrN0h5ObOG
/l6xDy8oGSWuCsLATuztO/5nQj12i2QzNhvEpLifL5m2fEc1Ras4gMbtW6Xy
6FGUEsONYyu/QBQMW7dQ2tvhRpzSOl5ApCXcL5MTg3VHfpAankdn1wieTE+S
z+O20qeJphWdOhP4J5U4e5Hcpg4QHSrG4lfmKHnAJcpwpwyu/clB5nRDD2CG
SFVb2/ruwynwJzuCB4K6aZqtcaMKmQ8JgSUb9423XwrR+6bC2wydhJEzCDZX
IN3glyvmXQLXR/0/Et/Fi6bkj1NsQU7OBZUcBciv86IBcY1KYWLsOn3Z0Sc4
vV+ZVL1urS6r5dEE1wXlOVea6/WtpqTtY/ZOvKk9hoFgvkaPW/tq+yJeP5oC
W27MFFCwXbnNmhLsr06PC7x0sxHElDFlffHuNWXJJxa/wA6fVXp9/edslFT+
tZenWP2kp2qLD61p9gKdEp8QlZDGVxfCVsXjVWFzlZbGxdVxoOB8FaDx2fok
ee4YnG2DcCaivlzi+keLaq8g0+QwSthGJ37RKn4EYgI9XnLC5rDGnPTT0aZc
qjUbPNSsvkp6uFHhzAGTF/V/sZ5EFBDmVaF/r+Zek9Jq7FknyUKTCmRZ7VFN
iIOpbEo76tHIN+FFoLFH/zK/FOLVRC6lnryT0KBdPkDirIHltNiXc6+KzZr4
2/oZXDLcQo8wpOy0x1bKlR83P4YOizAYOaHhEKzt+Gxj7PKWhuORwhE7F5oi
En/xf0muG/Sm83oVplxnP8JSAT2aKQFGNERgwLR9Wsl4T1ztCGpPPR2mmHa0
2/ZRTSHNfRaiyWuGOjUqnSlZJoOBGGxENJsy25zOAQISbyFDYswhb8MYXMAq
6xHyptmem8aEUl5Z3CXoQkrjbC8bS34ozgktl/+xo50Y44OpPG8xyrGWwaCr
LGQN7Y0XeZ9qVGZmhdOrtkCWJnZXlsu55T3NMTxVf5dWC790UalznMgz0PhR
IS0f8s4kL5USAjq9GHhNyxT5uVwzITr2rjWPBHFpGnlHXp1AJKTYG9YZ+Xwc
NFGBkAo/AI9zGPOO3PhrRYufi7tMucW/xXKwqFvtRjS825z3IAHZUE1e487M
wRELg453zJ8CDuNaqo7oecKcpDl0CIePJkmXHx6a4D/HAAp2qk+FrSg1MNYG
j4alwRoCdkZn0MOKleHX5MoghUSBbgKN69OJ5LYFhOPOC0M637hvIbx5lpoZ
XmuerMfJ6Hs4ALuPK8mXKfPC77ig+GHlIPgmuYvhZrWfK1r+t0s/Gi3KajxH
Oof5jD4H/UuBfFeL6zGssAPlDxicDlVwWGeiZWRlcx3xvSOhPlWSAjvd/8Ls
vQB7yRnwGC06GhJsqc0xp4YIQtrDP6G1GMox+JOFv5wN9nEwr5yKzRVsCHSN
BYQXUmU/5TfwgpNdxi4wEaUIj+aQ4hdW+LMIVHKxTJz3wFptyE9kPTiws+xe
qT6sclM0hqK7NHsDavDseDvDjdz9M8sm37fJU6dC1BLxYj2B2+HOmqIdm/Uc
UvHgMzGjjR5RHwfs5qBDhk2JriItxFHE4OR4Tx4gBge3W/su2WtRHHXbVx2l
5Sn8avw9fbBvaNwVAgRFwj6YBdyCw0mY/eIEPzQq0fltFtkZdeNBlWZCr9M/
DjH4r7ktG/21w+zypOz1ZouEsnD03kdamiJWGHEspimch8VulaYFaUNwSrwV
QulxmkB8+9yAzxnj0V/PT6L6LTmvtHG4fvxiIFGCsnv9M9S3O9IwNgtBrml2
xQgidxYbMh/XbvHuhv9R67R1rDLaMOVh593LZPdv9bFZZDOAea9n3tsoVvbL
h5ix/3oKBatE0ielnAtONZIPnHJfc+lPog+BbvLSWPbJ92RGeHfOXY4agT3P
TTJ6rItW1Wngop+ekvEy7x0tIGIbXAdxsuT2AwzgoyibRQHxCkOI2VP3fFas
OHZc/1X5yXw5HAKftBtRIYilCmnSAxyZnZaHJatNTOvyTZFEl7F6Ck8sJHTG
ffSD3pGB9hDjt5NEdCydSe+DKNovP6XyG7g9bnZKHq3lq7gPeVHf0uBL8qMX
lXmI9lofn1Fmyui+NS3xHvhJwjd5Pa+MkxPdeKLsYq5CLZfV7UZpeRjoAGAV
DwupfvqshUnUyukNXtM5xAndxdtS5JYV41oxle7MJcP61UvofMvV51ZAaw9N
KuMZ1UIUfOsooTkCsa/30AfdkGQ6QPDjKgH7x4eP3++5W16hnaESbDThrfW+
aWCtnZQeicoSB3JOpNSlw5D2XnWpCRzYldk33tCFZ24nsKMusKCfKUJDvl05
YB7uo84eeBsZ1EYjjGGvkAnEMBGBN4nv9FwKSpf7VYtUAgF3KqFNMTldOn7q
xWS2xuDo8Tf044I5IqPV6eO5vtlAjeVOkRHA3lzKDA5D23pwN4Z0hgsP912L
rZ5nuiFR2DdF9AhfcOjUa6hBnqDG+I4D32pnc4fK5tMkOl4ZeBnovrxuAYVU
Gr0trClJSczgJiU6znv6DYl04IRWafkxI+F1lQLul5k5+FHeVVwNtzg2z6Pl
Q0GU7e14ZgXzM32bN8J3YdqoBMyN0+OeEUhIdjmCcoaA82WeWwUcmNHnSU50
SJnY6WHfO+gZ6g4I9ATAKcXl6GK8GVG5MD4aefWzTAYCeh50FepOxODBZfhb
SUj9GxjALG6l3RnLO+6ws02h7lykuxIACxe2D0GTr10tDjlGOqkZKCEuoRhM
nI+29dFq/03Xo+7Jv6Wox8YdqcBzgVPHsXhubxAu5USHoHwCaZpQ3DAq9OGl
fXPmWaY525LLynzbGZbJnm3ZXvAQfvSyRCoow3xSMH7HpSb8FtnA+jkcLzo6
sAXW6uqG+dTTwaorAvXOQq7ne/2LDzM+JC+DMREaxIbjkZQSWdTJp02Quo76
ClooTwmawOYkOoSQBISchRYRwauy/Vy/37AONJ1BCHL2OzOBS4gdFgUbj86C
bPkRANda84/INQGJnnYYvF4DfLmjVCRaE/Gzp8/PBqwLVLWc3H2aHXQJuz42
wNbfo4MLiXr6A0lSGQEnWdENnbhidjy5FRl05yxcD8eNEK1WFh8W+1kZA8j2
mhqjjxq6sb8WnrkMAacH27MApbN+oRI3KCC3yUccw2j75pbuXBit/3qBwYu/
R71dS9XZ8bTeTHKuTE9zcnk5442NjVMXiPM3gvzhjHj8ij86dZUpZCZWi9ir
XQdb54nfzkCpcVSeBqCnywe1ttb83GFJMcqdXKoB+phdE5xpbGIYcO6BMePR
wGJab5Ayko4V5gZdI1saTt6M5tde3ZlGLWNZzaQzeNeoYn7g24k7HwuMX62w
51t4h+Uzj+1cs0MnYysvnA44LQBUKJZDgxzPMxMOCXl1Aq7HzM0mzb/kJ10X
MFte1Co9Icuq0JBN3ygUeTw8DA6X6D0+inu20stkPqfBMxMhqWNXqIdlSPV/
Md1s5l72h0oMqV5393HLRJRz420cPw7a11wIvh+xOO33ut5B7NywE3B+kkH4
yvx7SVvsPw05Fzgaqh8M5NGTg5qRqiIb0g+yI7C7dPj1GB9KyAFC1cp7JJnU
s8hBFyZdJiaiG7/Nia+DgvDTTyKIZeJ9ShX4/l3rNEDNTMRtvT9xFyBpAM91
KNRIuwVKVv8NOGiTXUJ9lAWc4HXPzkiDEkQ4bmkS//GER6F3zoEjToLn8EVp
C88vjGWK7VRWvGBqGlIF3F2iLvn/Vcf8gr+lrIndIHAq/+rkuKIk4lBWPdSk
IMZziaigkqyWxI1kuumzwtbS/bjY0VeiKAAHtrrt7/EkN1POpQXBFehq3X17
+KKNlGRDt+HQs8qCqZjwMSl2LGm4AUP/kj43sdTvsyF5FkTHOq0+8DBGU5bP
h7meC3o06GKE37pmA9Nwi59BX6uHwtbySEJPGDGPJRJ7JkUJqaCjcm8Zjnwu
P1dEBk/pcgrcWl+hqclM8Kp25yKYDxoP/EtZaRDS4Sd4hUD7A3XtCwtLEq0k
GFFQNA8APnssCQBq9hawwzRT3kqB3NDOiTkQBaxvPVmkr6NbP8TXqrMI1NEs
ukd6j/RTuENS4B/GvRXbqgUSLltROPoARo96JjsjpJFGepPujBgGOe5h2V9D
ZHJ62PwBL+EHOE/WdmR0DaeqRiSl9EyMzz8jxG3Ee/iAinCe8GbzTeRR35d/
HVJdSYZDXH0geme/0DRGOFD4dJbaqeZMY5PUgrb+wH2onz2WCq4yj80wtOwj
9XP0wWUcUwqYOrBOBwks6+vi20Y6cFBfUFlmFo52qL2L9b2vsX+gq0kOZNrP
WmrLd0p4Ybf3Su3yBN9DV7IPAOyW75368bZsVBkjZUv2iIYfPFvUr832LkIA
aHIM/YDp6OuRfUbiBliB+hL9UnOgPCRN4/Mchs0TilWvXAODsylyhUfhksni
w0B/wPQpCWn8fb2H37kyG1tcZBKbyyKx+RxU5aYeM1PIdLqeYDXYBc8OI19V
5SpNM4DQ3aho81zXgR7ukkrGNkHo2ig2Nv5rukoKguC+1ZkqDUYoIW6Lo/3N
K6vxn00KDrfqcasEbd8Wg8ItvjWXgbkKiiIr6axry6KzFUD2NdRMV3bOhCJP
WY8P8/uA/cZpEBK8U1BUlO9So5eXjmhj5jxxzvcXTZAM6m9HU2wFsoopJqJ1
TOsYaWv8rT4kp2aerQRw8zJ23zwc2fcAWRuy74Kkul5OMxxo0OZnj/LYt8Ny
h39xxBbQ5EchhK5QRjBE8PlwcTaB+CYGjrvn+KLHwQdHX2p69sfZh/QiSnML
/GZleJ+3w7AeHyvMI3mVtM+wsAdkuBoIsnSLazIRYFsA/Blop7+LxlW2dkB3
v8nRmGD4vs1pZZVdbivljcxu44ry7qHABoTjg++xBfBNhWmxNYxs2V7bCws8
p0fVaibAwAf9aIhk6KgnO3DNkkHxoLRdrunQiGSenmVhSbuGldJX/pMEnTWM
WijNdf9bkwsv77ST2NIDUte0sGpFkajNKedx9OXqrfVwDfJTkE4zerqlVHjH
OOaDOpaqlKFa94/g0r00LcySXufbfOqxyMWaOFR+oHeuFuQek3pHpvqXfxpY
x6OyjFmFmO+ZjvuR42LYufxZS6w0VQSYEVjBu4DvyK23MdPUkXngfUrkFwYH
LZbKjNwUdenm4P1OXn9Var9GO1gyBD3eo56oPZYkTA6HNROwwL7tWNKOhsYr
HvZphUMpwarCKjhQkLTUyjdXd481fMjVxYbaetNMVwk1HyhHrOFGrikVbYIs
mdckkjVie/FpOBOmYggIfWIumnmP85G6mk/HfUrCcAbuoNLjk+cQI6N1+nw3
+zTJ52LX6W2PM7SlxpmHybfgADFz1ppW2tZOdVkKi+QPx+MEFPWDoUZVyN8L
71zg/ePqeZEGrhsbBUSD1OWYkvl+8/k317KFOEfT0jYIWvfv7O8Ze5NGn8QI
jqI79KO3VzejzVIyxKDRvoH2Z8asqslmDI46MuETOGflgJyJXGRV8mn2+CdC
awGoCcMS/ueoi7E6hiEe5CaiJmyeAUB2IATPXU8ogmiBKWes7Q7A/EFQ8s5h
T/27ntEgy6RCqHznvZ31zP1C231Blfy+j6vMdi5wN28+5ARybfe9TaIjYC9W
/3LHpKNA4G6XwVSZ/IpUEfKwWx3GwtQ+NWdwezq+j2X7J4oKPgxrAr1+5Mx5
1NNBEtF1AYPVKZO+iuh7btIyy0QGFPmbTX/v9M326/AOthH/fzVfxYA+5IAN
dl7a/tzgp/tErZg0YXoJ73L669p33VOJKcvuKaAZA+HNGocyPwUuc0cMpfge
gHoYRlFKkPhke2B4WmWCY7VcbXGY8mJDdXAAtgDbh6TcCSkhzR1ROsR6rC+4
+p6zOfZ1eX55JF9rwzm3zt8WVmdTUWrbM5PHCYiSqNN3prh2K+kCVGHTYbuU
ZdFcaRYrr7iLfEQD/FrQZQGGnTuc5yZCicrGRZBC9tXERD0y9qer3U+IiTYx
0X3kXdiYZeQafdwBBRfTp9ZXLuBTQ8G1rngMj8ajFnjtOjBtQqdNRg9HJylC
D/ygCiHJ8wJCgS3OG/MrZlZpQfyq9AeotrQSLrYbzDZDLijnp2bN+Mo2ijO9
1O2pvPAwzKLWe4f/uRzaaTtJLosrjvmNQJ++3DauTuXBU5VaP4FHvi7Rvk3G
iYa25QGf14s/8lBLp2/j2bnnTRvK/WHNEEcskrKct/DM4EknM5tlw33hvHde
+TZhiUw6l1RsleGoCO38YZpyxEB8P1NZSovOJVNyoBMuZHlq+ny5pTEd3h/y
PpMX3IM8mJsPc0jUYCsYsxPsVsaZ0Kj4p8RgnTXiAttS43JMc7rqY0u1FVhW
5+0dTkibqQl//q4R8oMvR2erEAZheiJFK0G2O9xdVLJVLO/WA9OR4zeCs3Q0
+LM+brIZju1jHLZeRBZAuSCxZs6/ez9jdFdiLfQLtZqqMHNh0AxRnOJh6d6X
eu1UqpoowZ+LMjMQ3Dq8tSH6SzyZpQOoVWk5Ib17o5upkByFOo9O5qJY5uOL
c0HDPsXWG1aRnxIjXcN7fFto8nRhV44Hv++HIkaZLh0JwketdrwgUMMIhtW2
iAaGHbGdeSA19XGPdabzD3oHd0efFTIbvsYpfgq0H197QkKNRgjm0+U71hA9
04XmarMpvbAReyW4IjTqOL5HctThKLv2Cfr/1AuDr5y6ObFWAxhiCIjHRbsZ
nrVATmChoBhob5xIwVBrgpXxKb1GvBVtPnocTnE3arIO1drdtBwjAkOaTq9r
S6OW4ySVgXS5ClxfJGB/vqrteXpvk4DbQQMdOEGfWsSqfL7cWAJi8BfWIyqa
WZ8IMJissgCt59rItZkutmbDNzpkrbBxxwYjXf6TrUT3gRxIRhkz0jvFUuI6
knYrzUIGs3sCnwCEB5G6BEcaJbP6VVp/+g09sGOAZM8vhMZzXKkPTqSbgOh1
73ZeAWDnqY4oY9d9SYJikjEyRczlZt0Rk+FmAgvKm1hzmJDqbVjabQwpWcUs
8CVD0BbhEL6P5fPSqntrKZ2pBcPNr/8uZqK9YdRcA2mNZtdXiGnZVx/A6d5t
aAPFJgqBGUS1s64JnKVGm93+L0/AQsdv97+SqvgYQQW176WL4p3+tpaDU/3X
KMjWo5F2uYadaQfRdJZk2HeaLrgSpTwAOc2r2lXl+1AWNsSAunUb2C2kXeia
7XM9ramDIAZYXeHszpVTdP9IENbmtWM/hhbuDq0rl3NDzU4vMeaSdVKon9/P
QhVSA/IgyQlM3vHdRpIBBpdHdHnZERdKQsDJ6iTWIzXhDA7wJdOyW8IMZ3fQ
BQksxJTcIRwHP8mVyVZgBoCtNyOLyshgcTH2wGfc7FpJjoXl1lY3ziCh9xPM
K3qx6pPUqsDkpFren2vo9ePI/wZb5iPH9pntYfl2V+JYOHhUxFYBuIBjzS4r
fl0BVJA5FH4IATbLZ9OYLarB6SAWUmnjJggbY+d3SqQHPoOQyceFKGBJQ6ZG
RBUKHeGK2n4vGpp4n01wpy1KHjjGuwRUGVfgKhpJv4i0Ki0A+G7CYrlYoBGJ
/r4Sy9eLPh+Vdjz3Z92Th/JJiCYnGd2iAMqmCVieHztkRaBpC3dpn2Am56uW
bmYVZsYuTLCnfiK8IgJ4K0baZNIDQVw0EewJNJF7f/P/Z90N/5IqLMq2238W
7UI058qY9hvsA5o93pN1uhFajBNbnbR46qY0RpgjBpamdb/k42nfpG8e744o
rBIfrYXJ9abQvGPkKUi49VAwYytZ8D0KYw1/ajgwdP6lR+4+h15sT7ovWcBm
caFvWTLLZGz1Qe28mHallpA0hcyQXpg99DrZxU0HMSvOtp/zfFS56yVd9C5z
/f5X++swilcN83C4fYjgjdoBiUvCZ48RtCI/Yq/79VyV+7/yAV9iPQ6UA1RV
k2rdjdlcWTZoPGWHzHO8zXTxkgLUDDuWTAgcwG6iEDA1U7Rp0x6lciTeMQof
3sA104LGVFqAkx2shOGyof3SFAfjEh8W5QRNkWM7aYsLSEuK1JlRdhapuWjz
w2fmqQ+ve4AcFWbbVR16AWW8Gi6+oMx8I+OE2ezmr4GqlJYs259Z0nnUnSvd
yYAgIssGamIcWsbdogpgOZ0CX5o7rxtwBhryqu7s6rQyg67Ze4pykHo+MJ7o
np32rmudySGAfz/GpAa7Mzu1lDJeK2ZnSCg8olk1wuX43E3oWfdYXBEqA42p
IyGyAxtf9BUMFKkAvnf9xip8cA3MIf6SONoMfyvFMuQlWxTwBpf/8mE4/WWo
Ls8n1fywXYkwIk9sBESwi8y8tLHjbbgD9nqMI3TKkYlG8udXMqV11Pk/6wnV
sGWBlSp+lngT+0iZKCasP8i2NujOPoRTHKyJFDlYmqS8GsbThXqAAmI0oG9W
xvJ9tymunoNkSeZLouZqpAuhYD4mxQRJPbB2RFa8JijWXmmaBZ0GENEqsFSB
yPe4NsQb20epb8rqoJIjKsBV5nFMMf47HfOxLt46eNrGJyxaGTeK+YHroV07
FV57rsERIhgnLStMYf16OzBo+X42buwcDjHzIZV4QrRa3VHSJu8/76V8nHcj
oo7j7wlf7t1Oedk3TEMO4sYoc9fCy5wEEDYLFB8nAmUgPoAlbbbOUaGQwEwF
o0Hf1tQO7MwSi8k6qaR1UCFJVPmuVT20LKEru9yKZqR++iZecypiRf8I6SNk
nU9qBaDiXN9WimZuQC+m1/+ZBi2RvYxmdCdPiMSj2g6j89b4Y/xWCWRY/ZCi
bJpo57mvAFSq0tF6lkCeWcVoWbwruWeuYsbweVCl2s83yiPM0UjZib94/1Lj
LjmrG8IlE+xqFRq2JnlID3Fw/dnzdYF61eUXIfmIijYQ6XQyN3xcUftgOMMK
eEOfOMMeQstwbxiYeAr/UrABmU84teFXvbQQkG6KKJrC+39dqx643gziu09u
t2+6RstHHwCIsiB+lMQQsZ20ovBqjD77VFgwerd4I+Mtj9qBGKL7vguKk1Wa
WqKKhL8ZyvkRaagIYH2Bykh6TuwOt9QXh+bl+grezq1Qou6z4lPNY0sveUGi
g/OanIpYf4XFtovS9NJbSkEJv4rcjCrmYFke3drFPWXeee5oWWOYZxF84k9/
wB4oqxXVjwvLYbPbjjlac2CRDECI7gGnigUc9qW0sIV3lZqBB7kqGIxCwIJF
Ax0T7chYhCVoSeonXwCHV4es8xMZq7iEF5omqGzXMgfYqP+dmy/7OFyFgYVs
U+nDuXm5Yr0YQSD6uRDyqOyPsCGO5cfV2/w/2mTCQz75NNnvjzwcQXqQD6Dh
Y6JSkU5EE73UbqfRqU2/+TMg/ach/Mj1A/uqky7KJbUtow0bIyLaaRl2B7fr
xZlArmC8589/4UQ6FNsAEK7ttGu7JdEl5ae/t7IxV95W8Dg4lpuYUFVdBuNX
2YXteeIC12tzDD34KOTA3D0dkSTbACCuDYg0ebugZ5V4T/X+EGqEoAByMEg9
lOEEzikV7Dd4xe7fjKIA7EFnoK19jwwJpSY6zxI0upB0vi+Tuo5s5n3ICEab
G4xlHb1GHgEtsl+Gj4QM0hiPax4MhqClbxBaktUUg/mZ/mrrzqvKTX3yj9aP
1iuSqpIAzBiYjomKfhLfXqXbe1Wwx9cFratEwPEZlCveRN7tS/OneUjNzNbB
1Lxx6FNiFxsIlHA8sQMg5ZgpPysH0L+kOdJ4WKp/N8snCxSHJQRboI+jFyCG
r3QWOUAxXHW+LAsmQXogyUCBF9HATpgYEH75ZOsByZfz1dFUPldb6NY6Doli
RDqaKXask1O7diZdqYy///N0y+9q2HYDLtS0rTKlnx0TQiYwIOQHS1cMNYKJ
XwbBjGocWZbRkm+9In9JV0aCU0rqwFl+MBcUvAZxSh0N11Anl1W9tFKv5dNW
A33GGGuLaIRtu2YxPppwE9HEgQgKFIKqu3yqTm9ieRmCEhwXMkjdFQHUa7cN
UKTe2S0Kx5qL/vCN5k+WBjMPsT6m0LHC2wCtc18qtU+0DopHW3vF6pCMfB2W
r0XVVJtQ5zdwcru1Xw1VFVxQ72B/IO7vdwWZtSoH6UDeznXGHuct0a/r0VWK
PAg1wOOdUg4+yBQ+KYYBQhU1H4bT5rLlaVe0O8FVHFRkoUiR+gvbvhzDuMIu
G5nKbELEZTC+rgTbAwXrOkGvBLvI86eou39r+c3F1QjCLadnbJjVofMKsxPu
WTOPnR3R0MeZ4mAFg6rpcfkItH6V+/n4gnfKXSSDdKt5Ze4UMcVTIz+F8oz1
MYFCWP+CjnGSkFAgT5qmYNvLSur87WjxVk/jBH/Ll372a9Gd+ROVa4xQ91N1
wn46+EhGa6CgYHexzvSP8NWYQ3Le8WNWVVnnsMskR3nTAfqJ34JkytiChDXn
xir/ccQthj7ZDgTULcjRI0/7jYJ7zksHjvx2ctYXiJ6FQSjf3XAYo/dRjhKn
soOyWrTvgmWbXoOvU9K5Zk1YpHcG8uf58gRPSgDb3Gs8/vAptw/Cge1Ai2iR
3YInpQdMIWWXqnpaUIMMUsKXw6M40z0k3UPi/Vjnnt/1LBxlndvkwOUoQYGA
seBJckep1WSDhm7G4KOrI1QOrWhvvzzDkq4sK0izTDhbd7iN6rpebJ0hRxFv
p8l094AoaY5/+qToJLwKTj886/csN7CFYFnzmsZZ6F/agyPmwnM5po23v4IM
yLWOPBkPI93hvWQKRhrS+80FW6nm43c0yP7/8gFzkmYjMyJaYhDJt6qx/FlF
jg1LPaC2sqauCMvC7tPQ4WcL5iSnnhjZkLPNCRUQokIPDuZKism/kTqIJYYd
JlB+hjERIuxPh1du4YAV7FXBvv3FW64gJk2vNuF9mDGgffGxrAjslFvSJdHv
gRkecUnOY+OWnnykM68uCovA35yFHZueOQdfrUwNeMp98lxC+ynTupy1cHyo
j8b8nFCs5Ltu2JY8fRhAPgRqMvVKv+zdhAKe60zyZMnzhNNu/CsR++aKa3uu
RuDGU2d8xCMgO50e3FxmbWNEsM9PIWMSuD3Y7uRk5izgmJeOmPy/fcDAjVAU
e0XfmExHwR2plXEAdOpaUqGvrWMjZrXkkO4NqAt1iCcyKB5t4Xx9IApzYESS
N1zso6AHUVibtd48jgm2fwsBFOQktfzA2ij7rxVQubbYdJPZw31h+sL4WDwg
03GEG+JNu5gkJWx8SlYbvu1G5uari1u5R2Nm+eN5ue3e0aDvjNV7v9PI61Ty
T00BTbvkezEe0spHJIRfdbmSviBS92UsPL5rTK0p9ofl4qQDjP29zKZtcAE/
lopZ0BLy2mpNDTGvGf2asUnPujZygTZw7PZKI28FA2FEQ9Xw9jy4pucqzFKx
bpwb74PfPVoIeKqj53P9u2cbzQl3TIgrjwzr6inr2PPrprOiwTbVgYb9MGo6
TB8rn7OlEJjbNUGRwhAjzL62n7Lf5qdHo23wGe95SxSXdCZUqG+TePVNiw6i
3+XyuZAFpT+jsKxGYXIixCMe7H8qoMdRY+aN3PefY0uXSuiRMVcSGCRm9UeW
wdfVi8T7KAaoIabQVvJ13nHH788v37Q6iZhbWI9ZtMz6uZCkJ9FPxov+IwSu
aHuXMyZ3dcpKS3LShZLlHzB/B0GO51GOoAJd3vdymRz16pG60Lksi7W1+n3Z
DnEVhwVpR6U5RZfXAepWl5YjAWjZ4jdaDahUlYfpwG6ouJ1xjnzwKChinyQS
2QGgOc2l4QLrUONOr58FRFEjTxyzG8keGZ4f8JzZdJ8z3Zn+xtl9DfTSigjV
ig88M9BuuU00mvDLDT2GEWoCNarQkRr2f76N6anPSws+Wz7dn5ZOkPZVVW+M
XsKHQxTkpohVByZQj0rzk5DNd2ExR21QJBCeqRlTaF4VnJ/afSWmKdjA+jRu
wvdpSkpucFSZ/N7zTQ/LqqPSGMgLhEiF+/lCOe9i0PkkyxRK8pgT6PwycxF/
KULQOPDsZHn3i8z9ZMbLULWlhjrLkRMofFhzeKbEibkFAaYdNAJ1tM8SuuFd
AlyJOc57lh/4mViZVwfufzYShzg7sUnxva6B8czW7xgicfGDyCZo1OfOvNJu
gooLkNtEnLN9fMZB7aTo2WlV/MXJ56iLRtcsbuEI1OjqfaK+oLXaE4hPaUjd
buSJMyDlVheafhtptx+xGgJffy/QTUj/Gl5ObWsCH/yP7Bdwcnr/u5FrJwBp
iuJy4oZJUkKGxKq5KDUvVTW5SrGEUdv0GxF40lc/TqxEuvxInXWaKB2IbEWd
c8R7zHHWNOU3uaNcZCDIgA/QUSPqqLvsi5Kpa/o8H9hCJS1c8GmcHxl+CiCG
8fDwKxbIG+80Ln0Y5ukrIMkt6METADY82cMIx3xm4wxCJP/1ETNkiCet08k2
zDqa486ZNk0+UKosFKnREIruhUT9Cm4kS+0MmFdX2O4DAkEcj6r2qAnhE+we
dXmCthCAooYpOu0G3omlG2HlxQJziJzgwKeRDzGZuY4UY+bRYHsY5jrjxTqg
kOcBv4IXuUJKfRGpRmPJ4X238wL74BvA2a0Em+HtIpA8iDxTzrgOnkkTX1Jq
fN9giX+Xe+9SXFFm2JH5U4AlrJsrCGAx4Xl31D2jGzrsBmAiE24PlRcYW9Vv
MFWpUWAMEwBRKJc53q6Uw2aIsUz38qudXr5v2uolBoYVmuc0dE7cSjxo48GG
RaGNMr23OrishNNoqGb5vn7SVxIexq8ua3qM0HCGTSGLeP3qM8zaLIdqdmYD
5lVdMAjEBr+8aBPJ0SFlbJ/WISx3nXLdryGq5sixJW+d+vAY4sphOWDAWdoM
4GRc9EX0tQTrJJ6I3IpHvO7ErXEypyUSzBYBXRd56MRUzKt++Vic01evYJo0
VEQc+Ba7W5D39uicZDJlp08o7mjiQOEYuwITFzsA+VuIDvzETsMDTkRcr1Aq
C2+6E/kJn5Oe1DjLwXPebdq0nxJbCJ/e4xMJOvfH9Jcr35AsKVX59CW/N784
ASk8Ds8ALCDhnVimxbuH0W2mhRbMNvD4rEq9JWo++zzNN2Oxkneg5wbuEO9m
DiKhoZ6pqTR4R88+SWCR82MLR32cQ1h27L0d7sBXyM7cqamxMeeRnJyia6IS
6zKPjJwWoCL6fWUVhncU99lHM5StIol+sAv1a/MAgbVCpsRmK0zVPtseX23r
arhZXRZR/dZxm6z01oNbSK2zTM9UgiFwsx2WfEvCr87XDEfR6LV2jP1jsQfy
urh734oahTaccmGUuPbp/0CNSz5p1UMkJoAJVZwbzcyaW3kLx0GXsgOyQCZo
BbS4kgGyhAyXdEFGvAAFoP0vBVMPmpBMuOYvrDmSulmNGLiF+9wHXgT5Dysb
l+T9FIR535P+nK517q+RQg++deUc5v8xf5G2je2B2LhhNCwwfOpY3c9BWAOa
1EsCFKzvkd28HD8Z9mmnOPnXbBpmBus2GNkQltdKcE6bqL0hBfdccw1afvi9
rGj58UpFhSTsx0ZfPl+Z7eLqJLKnl2/xsTr7EygVL6Q/DDRFHyWZ7pJRzU7m
py5E9ajlafxkej3W0o5eECrCoO2QvN+gpCxMPecu+8CkY79CiOLftMMlBpbp
XnkhkqWduL+HtsfClR05Z5I7KCVqXfbLv32tWAbSFKhnAczMORrfJe3USSKH
iNEIt4i6Dl9S5KB53issszgWdi7iMvzLL8gqobTIYdgTV08S0EssdRlpRITu
ZDNRgA2smedKCZcl58APT6fzE695aKh7QKEK8maMteuncvw6HrzU3+0UEJJk
uODmZiH+DRSX4ipwz9PF3m90hUEEh40ivLnxRrsuv8vxIVjy6tvgepoTDFTw
2DX6BNlhT0h1iPPbnqYMTq5l7XqZ+ZyVhAgaqUUyx/CX4BSiYfDT3TkKp886
ziPtGEtIQVkt7mUyhsUPhuY1gCRd9wEyDCqDrWLfwBmIwz5+N6cqh1Lelep+
9kYGXIwLFgsez0WbUBc0Vr5pxFWwQ5ZI0OoT0g1BCQdXC6DvCVHslA5PFFGc
OsPMwFUnrDYaktvh+jtmKOfqz6ooj2U1mF/JfkyKHtDQL429mvtU4BqYiKH+
n6gyaFOpKjYVl0aVesRn2i07xyJzxx9SUYVIq5tDlu0lX5ADSe/+9AXof2Jk
SckXEQ5tOyU0CEQAlulQhIVSrh+ccqbkQ52VAhA/CmSaDSqTHK6ChvDMvEJy
eI9lLiqzXsHnuAkTs2cTDnQw1sxoq9AkNq8UROJLokEEDVCn1f9sfS1HeQVI
Q/uMNivpOXV+SGaCv7AIVR/rG7neC/8KDspeBlwjq8t7keOT0W6KjiXKDOjZ
GhdoL4T8Z3c13ig629x6Yf6LDltRThgDJRk8afDyMBo+GXA10CgzUr/OP5sI
FQyVG5eekpxOIhijAvAhaKYaBazn0UM2Wku3BWsNbBHd+t/coK1qv8e10ur4
qsHgzmtBvveU1awpHxwrYVTz1tKk4+SXDIDf73a3N1ifRMdpeOtJKqg5BGP3
2RSwumRxtMiAAWgJKgWV/BQk+b7+LTjiERw+N8TWBTw+C0y/+iXtcdAOlSbu
0sakKAmQsAkrhuubeT6TDkPRNVw9UnG476NrXhNEZuKpqbEjg+V4U0CwdZfi
cOuzthuz8Wv78WjIIfT1phCGdlc5euURNjJT6Mf+ixeI159YytZ0qcqQ/70C
n1fYdaXDGYgYc9QhV9ecWkWk7h4tV9mkUUzii0R2893GIK94hzJ/JYz2Em4h
DuynXgEHmI28qZzH6OmDMok/I1vsCQXL9CKmbQjDO1gxDr9lkFGf54I/qish
OEylTk2fwQbMRVLkGe8w+NKJyBaldL2+UWZL/IwaW3EWNx4P10O+GPEBKkbw
+3CLwtzF5rXTb959xPCazaONpBENxvU+iGcSIHNsZiMUE2kiWFuk8X1yX9wa
brCapcMvgCNA9QTBXkIJNux69wGb3gEkN7jg/5pWp3dHmJvq2A4ZzNjem6ZT
m8zgKmsma3/uRsXVkHTFgzo+Y+0Pxg4hkinsKVMa6S4xpQG5gzZs7sZgup1j
8HpdS71tTIqdyyJL39+1wd3mrzqyG9AOBFAKC7FEDHSzb/GMrX5m6nsyfVWQ
dfg2hMGoJifRmwe+gnTm2yqh52yDtBB0dlg1crGlfFqPnf99lNbSZvHg0P3R
nqdTmbwVdtX43bVccsS5jJmS45vsFuJHFmxR4ojRd55topIDcM659gd9QR7p
74oJ9wPs8fmwZ+z7Y778O1L/O4Vhv/IdPICbku18xpVDByCuV83PTo0kduOp
qGw4J4aMMrmGzMPoPKZzMkKYqLRrTEU/htz19fBCZeFHlviRiLXXHFbscxiM
hHm6xovJ1sWA/xo6dCUN3npVO5rP4sDcuZ9d9ebltJe+y1Hw6JOP71Cp4YIS
6/zPKaHSgsRWQGPlalEdGBddJui2lY/bOhzfioLQ5Xk/7ibo0WnkIzGYmlLy
zVimeniI3pn55H1WEM/xQAMF4qk+Ri1ioyE3kuMTmipDct4A+Q0e1zYy/LGP
ylp87tQfvcCzlqDAepoA6r+olYNGR8AExMHRpSM3fBAK1HPLKLSqvDvNpQZT
qvNBBOK56X/xrlEdGQSRnNuQkfmXt7E6+K0c9n8jwoZ+wkMgBCpDZnK1B69o
eSf0ebJsjJ6BJpVQig+ilL4smV2KuxYvA78PGxTHNILyL5vK8qG2Y/5GWSQF
OTQxoliiCtjRpROV07VoCKHLCQVfrM4Ut4AP1/YcAa99ncjMf5wuWUUhwbX/
OrGyb+gRRUyI/xye9IoXCUj15qxgijNlBdYg5WuBa6HQRx+cbAkYkNb4Dry8
Xrfsq/mFijBj298DrN1KX6+uS60/zG/6MNC4ktfsuSRK+Z/l819VNy7vdiUZ
sn9rZ64FS7OciHRmkL9tYPKXkTcHGWJ1SfuzuE5BXKqyhp+GH/RsgKpQwE9Z
xbpD2vseDvAG2Ipjx6wg1A3xQFjGhsYXLmdw7RY4XjZXo+45vYEPd3xQBH6m
UZNIcF89G87E97o12w0tQyoGt1N+DXQ9rAuUn3COcV//5iEwR+C02U5vQ8Oz
njsPvl7FStjDRD5pYuJaEf7qj0i758LIBodZK/862EdjIUUbwgXbWZEjNy52
YK9ULHCutqOppNvKbqjDfPsnznbZ5f6fNghWv28j6JlT9qQJq3W9htj2Oj23
k2Zl6/YFv0V/raZdCWo30yUnzJAc8bhuEHu/fv/1drLF5NR+PHEaefLr0vB4
dF0ta2lbupu2F7G1BAeHMQuQDJ0Z1sviuBRrVKPh0R9fkCNy2tvId/jGkyoN
OVSLFemsWXXPyWn7oPneXLAtyglmHKXA5vOds8aczaTMDg44MukXwyOesjBI
JWxgFM/B73WCcqa9lcjej5a616gAmNY7ArCsmO2DTPvPjXbH2URKUB+I5D8F
rMipXrOqY2f5oeDA77XMrbiydnKHGT6uEzaDMHG3dGeernj6Lm3FP8m7ltvJ
9xoU1EPGnHKv0aj69HYOkhUeltsQGRK4lNUKW8WmYywCCNw5wB/Nua2FeD5t
QB6vId5fPLeHKZ3f61DY0BiBTgivkTMFhiwrdDG/5UlMJaG4SykLm4emxLW9
6fth2v83+yWQNjz34+AUCOitLqzASGk4K2HkD6l2QRkPZJENsDby20rHrhgi
FJBK0E9btzXvtIBCZkJAQ9bLjODA7foqMjW3P8lrf2+kHQxViX+rgZuMADO/
H6CbbWYkRw50HWCFimDl47vZdo8bL+ESXNDejD/8Qm0+S8RqqGVun5AxWPWm
DdjnoHkcLAH40DL1fygeOBI507stZXkv3BEpSVU5KnhdARIiUG0Kdm3TOI6k
977wlQSkSDp1xb+UbTgvEs/w1WVXLRisznTSkviYuqnUF2K5YAu38Ir99amk
zvbWA7KqHA1OsvhUpeiTDIIQSj4oTtfEwNoLV9vec2nTV+oI3hEwKuHSaKYH
tqJ3+zf2FqSGe/1CAJyjKzj6LY4jn4nK87J9T84uozCa8Nsaj6+F0zmwTDAk
Pdepm4rjts2RQ9ZI0JTXUCoyh0rS3DHutiVER5jGHjYs9PxzidgaaZJd1yme
fkj4IqWCS8BzUT2Dihh4BYYb6PRgSxl3eSraNI5Lyb6RNTyH2L9XifqyzPvR
Khus8MHIoBHcG1gtPNgM8MBbzopfaM43gK4J9+7UWM1Qi6Tx1umCbOfza6F6
4KJmNlXweoZxmIV4Ti/GfvSM2HgctLR2nijGXGyqooDdg2GRN3eOrBsNdo++
KMFGfOSUf17tR0JKJRHsHSFfavWNQ7EoHeJq+TVisMp7NK8BhEScD2o0stk8
S7ZkxpwHZHyF6CUyb2seJnFW5fl+kvperbmjUZes/cElNbLL3yGZ73WcPkCD
Otuw2HpUIQN6kagR5qA8qjK2O4vQvHJlVgjPPYCrjsxpg64vkKd5WIbyPCCF
t6s/ZaESlAhq1yE6pX0KTodWNd2mwdEsRbR36x1z6ZFvDaQCccB7m4H38BNj
cB1L6jpqjroHCa6HtfLaXhAmgeVLSAWiQtDQc+KIQ2SspB1W7A5PX/vNdiJh
tLF0sfZGnRxgDnAfJUwowZvqvLZq/x9kRQ2V0fx+I8xLUzAYWo6XGhatqcyj
Y6xv7BM5JoZ1vAELXiZlRRzwJkK/Ihdy0GHO8zrDFCfzXhSoKxP6x+hjFZv7
Rk4jfnJUwlQnX7sD2G1iV2y5ecaDQg4lWUz0ZdDxyNRLe/G4BDdQLvkyjSjI
xtqewYEo1+KZcqb2ovz9Z4+jeEgwz3jFKGeBBsQWw12Y1al+H6ePT3HcZB1x
M6wonVSxP7C8onUEeoLjfPobce1XItrWxUmqkgeemPi62RGJgJagpZqchIk6
XYiphhFxiKgHy2B9ZgHMSATT5JKeO8W4/9jC+kLu1WkYWEN6Rw7LiVGO6h0A
gA8HTD1D2X8O9a76r52V9MlAR1ROb7GgqTMlFXD5dEeUuGQABi/7zYxUBs4U
ETSVnrZaoEcubGDKPjCdx3jhvLLWG/D5wcpwTlMWlaQF8HmK7Yf+C9HMXTJe
tkqLO9DQm+dSISAMAW8W6rJqcu7YOxo2RxrvH1liI4FeDLhiu7XsQisyxrFb
CXmZ0i3ItqOM+UaG5CXkMykiR2AytXyu+Rt7di0Ko10ukP3//VQHN0TBORp9
6PZ5JK0PxbtQYQWxTODjv2NlVHeM/kGRXgp/IYA+FWrptlI7qJkzHMO0kTjP
mtmRgSjIFqV8HzhFSsyvYTb8isGtRs+KJzJDBLCSW++IwgF/9lgb6tUjPVJH
xBpsr0geCTo3iXd0hoxSj8ZsVraWoy4N8GcS/OHIiCq9W4pRmQ/cesWT8zoD
q52nd3ddj7Br7F2Eum6+dRGWmKyU9VdgIqlj66disYKo8tqySHMkXg+Km1Wr
yXiJgT1wCWNgEjCjNllhvQDQbznmQGDm7PEco7utxPerD2x7zVmOtYpRedeU
3rPye/Cluk5tCbxqvtzo7hmbDuCt6X09TvIfXLSl1qFiGiYOInaDD21aVYKF
hkSmgCZpIJDzL62hQu5Do1cslEEopRYUxVk1M/ZQoem0a3G6O+0620G7tUXz
sUMPOFHTAZgRmk6ijZ8S+aLRuIAZ31s69Zfd8y5Q7rHsXLrEDzBJcw/7mJMw
uHndBoI6YAxVnBqy+RSavPVpbxdmJjDWesVco1+BkE1SEGAmYpMnb7RhRBPC
Yeug4+8yYoBBVvzRdDmOdLpdoKV9GCeZ1lXzApe0cHUzLhoasTuA8KvF7Qmr
STNCob++Sa16YHaMgFRCzZFSILYqoKOC9964x1vPF4/k1LWNMXz/YDXSTdw/
So39OWTOP/3XNQeAZ+xkSfJU37GqccN4Bi576XK1N6G6NxcyVrTdwBU31oEu
6Tyur/IY+sfUEs2DfEsEygFI7RLjMRgGDCNqQHU95I9SVEE2gyEfScip7z57
U8yc6KSaOgAXqOt9aAIgAtGB1xfyjEDWOOkdKFgIMei4f6QmqPCjPqpZhxd4
VUt49Zp3U7KJgBmzuRz1+vxKhVqjV2LJLEsqJf3QXIms+ERbDh+RUmWT8sfJ
4y8GMMUf0j0x2nvA/F3YzRXjnKQK/hth6ZY3AEZDb8V0w4/IsoJF5F7RDCHY
QrU9+Xre+U94+InjhxvczR1IWwf7bgFT6gSPj2w2TvvKB4SIgcVQh9oLC3f2
A6vRPHL9OMWa5YHRH81y2nzJe/V+sizrBsu0/X1Pmo7DshuzZUB6kXdfDIAz
l29vtODzPy2aJ2nua1puuFXicUzaKcvjPC+0NkcnCjnMqdFF3VRLzKVYyZfv
EsrZvsMLdAvP9Ir4WLmunkBq7OkVFCr//lf5YEUm/nxiipAeOEdKZMYHH+1V
mPee63spqvVV45R0d5qpPfX8n0lZ8x/CJPuYLVY6z5QTDM+HcMREDFBzHgS+
PFsNy72lvxXpmbq5yYhL48l8A5cmEr2XFUDO3QfsJZOi/mr/vvbsfbdn2WRc
ZJDxoyc0pKS9oqRt5e19M/mzAcjP4gkTXwmgSkXAtiVIK3nDLwppQStjKYgc
rY4Z5/u/97K2jPeYvnq/1HFvLG5ZzrSj1ndv65Amu9MBI1DVZ7W5rlL7I7Dd
BMlbG7E/OmOmZBVUPD6pN+A6HHc6ROeEplqbkF884hsx2grt/92XsTLcHYbj
NEDwk6uD7uNYaJXerWxgqr8glzA/Xx4SHBRRkykYr8qJKSJEHt3NFz7C6zaB
W4MxOKL7qE/e0+X13GBHXiVlb3+VVWHERYhX4yjLetFUBwor+CFbAYLBqL/L
A13T7cbzTUr2WZ22UE9NYH5BCzyBItkyHuq6CGOPdDyjAiLLrbpKm0bJCsAM
Fmcdt3vcYV8Vc3XqD3QcJ69Mk1SLeAX/VT1zX8fBCoysIbyjcKgB27sEPuGb
OIyh1Mz2pkA3nq3wK1btpE/7V6O22KhtfOtnW0ZrHUShI7AK3rBa93KWetYd
h5aIIjsygL6CiYr3Nt+bYDyYvnZsVEeWCiMstABWoOWINDy2lYlj2UiGHM4O
b6dPahFrFPz2l64S0igjIOLbanNrv44NjksopcAerPCDg1m/gkKXEriQCZop
x39pAGjw2cpsc7x0Nitgczx8OpcCV08yc5fEJ0hlJ70t/aMI/FfNbOVygLgB
QLY7Vz1KV+ZC2TXJ7WItxskeUl6AnC59P/5xAQZOzF79liaFw8+MPPGbDqpU
nXqa5dKv4svp8CkDTCa2eLkwtpZUCBoWYB0H3IGEMSxWF90ea1UaUBGTPoin
wdFGdHS4F0WIs3K/UejdfvbRefac9m9pOmOe/Yb1K/lCmkTBAI5iBFUbaZIE
ecUUC0e0tiMKO6+IWsjNt/vN4Vyy1Xu3tTonJ2P0gHnljOoVCT6d9e+zfZb4
YMtVbAMmg5u+bUyhZHnWGqB4WOQ/kjjIzKJRK6d+mS3aJwCKSj4ncbnvLQdA
DdPSq3+cKZIR6q2bwdujXcyWwNSDzgfUNMtyrpCHtdJdlHTvwZGilqC2wBlQ
IrI4RBpu7okvsBeG9Tt0L/SpyKlomGAko+UWFKL/RYaN9shYRj+fXhQn9T0L
EJb9ZIC0OytPH7xx//XmL/Md3OcKA5qHFUEUo2/8PSnp/TgZ5fu8dWbtSKIJ
TWR3+c/KBGenjitJXagHQ/HXe9z13roCTQ3SrLZnFztjp/fYLGDwaX8gl/Be
VZ2Rvm8vN1b7Yv6UVqd/DjTXDIm4/v3kmUuEjkJoHQ5iCupxllQtbi/RXI6E
ZCiPfwdpXOHdPVlJhs63dMNlmVMduNHyJ74TmLnO9Ius6ZslulpVmusvmaWi
T9oz4ZgbSVg8KdhoAV8JBXKEa1LQJYmRF81/KFL6G1J7B1NA0MlxDlTfis6n
HOTHpj8RbqbDZ/YtuV1itJ3cOqAajFJHczb57mhLLxOXeSFomnuRgASq5PaT
U4+WJ7d9qJaZd9ob7Q8XCZfvLjk8eWKv0r4UzIoZLiDw1TyJ+aEC8aAs6j3j
wUwd6aXZatoE2M4f8p6qPHMhZIYJwXZyijNYYKgcPzj04y82yX2nPdsxvGyf
5o2tbCj06INtVQ34IUsq4DUbkA2hNBPe8pui2oPFjxW0WeMPUb2Nu5EyMJbA
4IRiJKOodTsKqc1+YmNbrvLiAsfGiO8HWf3+z30rUC/qS9IR8Sip4Dnt2pRp
Os06pWmWyFIy2MLobKMKhTEoE0VEAAeDY7BZL/TIYPorfrpF/tmGpMxNqnME
H3/adQVvcEJbjZbWigJAmB2Q/0coLh8WPLSTYwzZMh13PoJTiYmlcTAHdtnI
VvmfvSo/JVTWAwGUnJehitpO3+1T3/rj5fuw/LVgK/TMruHBIj+pjEG1b98Q
h06iry7pLmX0T/LpGiYoOC1M53iW5w0JfV+L2BpXUTE2FpVwuYThffmT4V9E
disQPNDNAc3rysPb6pqAE9u9nFTndP8+rTSsmLCiFlTKkLplzegK7YQeY4Lf
RJQL8J5W1jDDhIuHmZoVodz/i3eHnCySlzj+X2Cr++8r6UkOD3y9y4o1uEqF
qHfTQr8kQeYn4L0Kfp2L7JpmzaOzc9E2XFgul48ahaPPWK7dkyV9AeJvKjCd
Jr5dba1IM25Nwbstw8iINh3zypbVsVT9x8OHHphtOTzQeS5bl6sXWrUFkof8
XBpYdeq3sioNqY4JqflFUHPaUBqBZTEyGJWO35U2AHiTvDgqVSdjdaqLoOxP
ScCTWBxUS1y7YLYzpltp4sfJNLud9R+VA7u7Qs9YcJftLv532oKunyauLz0v
iMgdfkjYgPqL7ohCJKvOjaf1WIJA/NcYr7wc5gW3WCnzP7WxXeXdl/lKkR8a
K6KdD8+rMCMLcXCj1QkZb/KHirsEnbUDeWpoQb4ck8T9i651NYGa26HGTca5
svStI1OAmOTpPqkNBk76xVj4YKR0Q7ygnGOEqgA7vu4hHMrpMVobUBIB0+qt
o7LzbEsT7qfNs9msD2HBl5dqnJ+6V8yZ/2/TVd1oyvfATLuGJaUtbwFNkZ1C
rImndZx7i6wLhs6RKJbZYnfUd+liG2zhnrdiIO/ybuvMjjEPVS0beEFA8sRF
q1yRa3AeKf88GwetXeW93N02H2YvM87Rkk99OUfOkVB/gvpDPPBWQyKzFpBV
j/spxrKgB8u8mGhobo6Rs1CBW5Pdr5HnN78pAm0mrl2J0QnizevU3M+Qse8J
WLtR2PfKyieFV9o5a5z81QuYPnsQzITZuCDLqCwpLlYD+2+6itvVB4qJ5rej
kj4aP9X7J0VV1yMRJLBqmqjHcPQsvcggLHg5ckpuV3z1BkXXhtqaoiQWq4ub
raI0cHWsp1uhcndf9hEN8CsH7FycpPw0gOeNd4rfzvCWateadSxLIjKakBQJ
NYTzdNFOdHXg+EaC4IOnMHnIt01j714FtyhjEi1XidNFL1OTo8fP74ryJRbs
QfTh4+BgrQXKcHvGlCzBxCkSuBMZG/3sNKf15pIJAuPi8dGgCrJ7AR0e5N05
GoQKelVwyvf32i4wme+gXNZHmgjOIewekKQpuqroumoX3guCkZWsG+gEwnBa
a6lUzSNR8KPTBLUIdz8FZWPCBFQ0MU0VQxTUYI+vHM1Xo1f0MRjnfZQFr4Zo
yfb/WTm8PSv0KQEer02OxCPyjbjM/SU1euu53WLjjkp9tDf9NOu94voaZ6wP
6EYF2CCnX/9UBeqPjGAE6PGo/MsfO+8eQDHJNmgA71d4vVS4KBODBV+nLxah
YdMAsTsNGggKu1kmRgqnsvmsB8h2uWclW8wbIAHoQdmpdMqwB9rP4P04bM/K
J//eJaN4STrLKKK1ULJur8qMzQHm1LNZZcdfZsMYnDRupOqN6dbIHg3bw3YK
5HK+p7ijUhr/jyvlQ1eykxxUOtvljhJHlIn9K/wd8LYYPq43NLEwG44G8Bi4
b5eW4vxRyNI0ocubn9jTo9n+j5dN9icAnCmQwa/CqzQ/k5RZcakR/ncny8V9
ZgoR5vZ8+mMoXC7wY/+lz7hGdHTyLU1TwLB9CAsPdyCsGQ0uCgzVvgdW7Ic5
RdllErTEjN5lfiw13hwZAVmfT4TCm/m2DfVg2hsdzFSuMm+lFbH6wALSS+GR
UNNSTsSG07DxMNfadV0yTDXwxDKJ3eNu4FvMHrizyQmshsyPnCo+Lz/wvoA+
IsgJXLdTH/Ik19j+pHy1/KYqTzITMkJKFXMwiKcXRfJVpC6y9bQBU3sUPFan
JPCmPSFq0WDGBhyU1vdxCTEd0DKFeZkczTrnwV6Mq98NcirXui3HWmr0EeXA
tXzQduuteewcYAzJufne4Q/EcOU8dRXAPOrn8PuQ4DZrrUs6fOcvePmyOaOP
MMhGMJYO0kx4B5vPLGMRVf1WK1B7TekppTEXm2K+y9wwxbycM/WfhMLxthpN
uyVO1cmROBEBLsm/aB3CnjPcxmvwkDXzXrZGq2EUTZVPLM4MlY5T4Ffi9qOl
mlVS+JCUnliK2ZMsijZPpq7V6uVlgHqu6DLBOaXw9xsvzHRKGx4ukXBZIGUw
YBzyIcRhA9XWBOo2OuBEO8qEynMcUM9qIMUAWp/F1ynQkagVrYJj6V3jbqzq
AFGuD3R50AlhDY97YD8jzc3krWMDAdNeQgBpgf5GCjsOsBQX8rHPzixvjlYC
p/EcKetrjdRGHo5eTkjja8MeWZqHrzLfVUL4Ygmcj3xwOcuEhfaBHzvAJU4f
4iEJz2d0auoeAhrCe96NshoRiZUccljZl94xSWoBWOX1ccQZT5mBcbm5ccyA
AdXLAx9qY0uzAmlk6md99VUYgDFqPjeoxi2rmB+dXBbOcC2rU5T0qmrQIx8C
fN7jF5CMOYujk+Rj40jP00mDSlWQ5wadUYpx3P1nDTq1tzHAtQOnfEtlUTEB
ug5nzBj1eXtcGYgPmL+xguxSDUSyrymhSO1Ho+eI+c8/EEeOmZfLsw7CqjbI
vee4yf+CLbyEblmzFnZyh1tb/Kw5Ak6gQve6PIxikI2lxzeXjRrZE/CHoR1n
frxWQTQDltby5N5cgq5naPRDVSCQYZWBBV5hAC28BvLiKd+h5Y1DJ9+ub80/
LuPJ7btBbi9OFuONOk2sFoBXBjpkbmPOTepLej3eit9vEiSwZrMXoVHr5S1S
NZHmF9crp93qCblZSBPGeWR4gALF89gZvC5xJ8aGoFJCahsPZuAlO/wM1lZS
C5GxV5xYeZ8fT/Q3bktD3f9evnDuQ7tMEZKqd2oKxlBbl5e6Kk6hYvfjhP4L
fMYBbp00UbkMmnUelRvWcyIbZMiGjQt7+kQPGoFrEc1feJXukrSW7pyb6Mvn
OybGKijuNV/9CBd8Rt7vkG/GtzU53D5Iugp0/M4D83TOnSKk3E9kSlGY2Cfq
KZWzhEtTGfSnuyLUfR3RCKWCz1sJbpZYufTQ/wPQzuCz+hMK9Xvdgbvp0oAz
iCQ04636QlFkgmV4vsrDcYq2jDoLhKfw5/NEEO+06TZzSp74DTpYeolmDshm
MoxM86Z06F5mlqXT2fHSfnLMbSIrGJOV7qSDNmWMJTuA2Y4cUAd7AcfsvGi+
8iye278vSsZZUqeA6CCWusj+4IYNYnTqGCgGl42ZxdoRKHuf39Qrtd84weMw
olhvTXJH4XLPB3CQ+qAQ09VS4/q/5uJDdREhn300Ut6f2948YH9EWbn1VaIE
NllgkUVlKLs2uZxJcmkTVJO9O9KrkqUF6h2DerczRA68gLQpcEaQRtuejWOQ
4QK/wUOzUv3nGMhb8mEVVnMFBzcIzCwE4tXprnNZ9lZpWLeqMFAUIs6DOxeI
LnAbhTDCgGLidL3KXThSBBdo18EfHXXMFiPpF6Hqkdb8JvhIK4JIC+2Upt/A
9H6ptJlS5Ims/LcT3Pd+bGaS7vsLtNHJvyarsk9kKBsu6YZNCjEwLocOjsZ6
n19O3u96mmXEEt3b6x8v/fFo7VD4PRl7Xf/4K+RzYZjdDNtb9Lo8rUuZAEpG
Gvo+CN6LL6Peg1IHiaxyYOqDr0BPt80BKPfRW3QrCQfRRJw1Ldg+EspvR3yw
8UCdb3Bw9DWJZh64wMfwU5wItyIgS+u968Wk35L3iTWHL7H2fsaG7dLdspoZ
G+Mz8RqVvg39nd59eBBYZvWzTLMcADHeWi2PchuKRTD2vguy/qfXoGULh+vP
ABEV6VOPR2pwXJTlU2XjlU42ugbH/R7hPVUA19vbSu3lr1c6iM5VoHmZpxa+
LKQA9hsgr2XlL43ZTnW3bkmKbaIi8ytVLkCuDhYoc8ecXUltM772kn0CibBs
oRlhGegSp+GWui/tlQdG/Xc8nO1hQFTFr0a4+jucTUPZaIM/Y7JUNK1hBNmW
homAIV5saX8AabDDvVwS3Hd8BUEqxt8Rc9xa3kwOpt04VPfcLRCuhwqzWF4V
lRyOIemjw3grld0qXOxcKJUHHOFs/8kcmlPT0UNvY46ROrXERvD/vC730atu
APUSqiAecISJCV8P8185L3PmnrtfO0weuLfmU9WoTdPWgApuJs7U8vcGU9Mj
yvEvFQThJMx9I9tZklc3LRTgU9Wnt2P2hWGg8c4ZcKsBUk9PMpHGS+OMWZjn
YU0eC7UuI5CxbQAzha+crOl/taED9cm6K1OVMcXk9b6+xTY3rwx1Lcz1HoFe
8VZKJw3VDlrcgdoxedQ8Tw2MnuAwQXLYRV8WdXe+oRUBXjQh/Tpew0xyoVGn
BRwNe9IJbA3aghV0CFwUly6XUv7WwC7U+MQkgrJjOS+HzILhxjp4jmLQ78uq
MbKm6cfrzpcv3yWo7Vek9279/5aeldAVDDo6kdzpZJDE7k0DfJL83Q6kcZ64
DJRO6ojUDD6HRIqIE9mohonPTAIqFjqrwmLSgcMAXGHdBcHPbmXERWmDMs6d
MMn5dkT64DP1hZR6cLsEi8JVwGy1dgRWd+7PwgwoDC+Lgpvab/aWX1JTSpbj
HUEy1UgzmqXUW2Gd1ElYLOh20/AgKL6bznVq5w/Mu2YiOtmtS1STw0OVDln+
1pKxZKs3WYmSN/vFwsjJY1xOeA3LBzcKEkIqH11GDczyEQ4IPm6baJ+1C+sd
pAGkr+sjbXPS0nLlU4HnCl/Nea5ezFQ0fPmjREn66VGH8FksmQPBxNu88wPm
guH07zcY/ePmgfo17hL2w1p+vAfPKM4SSisdxQODQTrBya14iPLP/TbTMOap
RuigDoDyy9G+9yXgaETujYZm7yumqPeYCfu5Xq3XlBl6Vtp97vP8vgKA5nSL
ejfhQzYWxoJ4UJF5iQKOQKZYIs8+wEzeo8KepFV6OC5mK7cvj77hhCR3XFdU
1VUjqvl36YEFMzu3rVvbnRxZrq2VRPN1yl1EsqqKdGphh9l+QgRpJKM/bxkE
2LAFk0eNZAZnX6O+N0IMKG7LPhs/SJbCE6JqXEw++pUw4EGH5Mz6uCCgQlwC
48tJ/pHshRQXe1TvxaWd243nMl3NOxLIJSOE1VEBK+R0jpxjjkLaPTMKLrbY
kjzEhr/qLsaw0cOOOzqPaZfYp9qtQhNWkm7kDgFBzEUVZI+F/uxTxmih5uXv
5QSF4FtbeWmwLqsxsFMQmzTo0bPYpyPY8g3bDqFtyxM2E7nDulSUrBty3Gsg
mPuouZuEyY+R8Ua5ihol/nQOY3npw9zcpM2X4hZFr9bb7L4Qt1AMiFm+38Z+
0P5B1sq1vx55ZvA+1fg2ra+Nh9eVVODURZpOgWUvw+i1PsLwo94Jrma3lTXy
uKM1qEGILcVxQ26sLtPwaJW8yvnRwgEnpD7TPbigdEZfE14pgZebYFGfahdH
DY3ETc655pX/2kyOYS2OTDyI/+6YiRrVTZ6wZFS4dtXuF7KMbmotumDvfX9u
4FHp0vSuurM7lCdyIU3vEo09V/Yz6XGta3te1eWxGrJSYFgPYX7EbwH9lpWx
2t+jfxAaLOhWt3lruIFijwS2LJfPn/fbWacJL6/287DhxabvBk0ZjDzkMk6i
W9gsd/p9mpjXazTHWMyedUNgoYuhNuBm+VIMK33w9kUyXn1unE/0HiB8wXid
4LXacbvUI6WA+/AWQ2XvQR+pbO45mYRU8nKRx2d9oDG2uN8hLZRIexH1GJn1
7dB+mEmX2TfG55tn9oUcLulnOIL7FscurZGl1o+PafCIdPyavhTZw1jMg6Rt
TXlsTeAj4wbMMnNH81vHQd+yP6vPe1rhRQi65jnQx12jcW4UmFh76WCpro/p
hgT8wMzk1XFBOEzR8RZ/Zghj8IaBVi4rY8hFL31TKAJJ6CDLlqOCh4+uCvrG
JUTp/+VFRsWk9Sc2p1td/co/0wQvHSsa7Yme0709Ngo3XOSZw0pEWkFq+QSs
k92E80qvGAmGC3VFqqHxEpTozszWIO0LAGqZ3ZaPl1rmDzosXV57jf/V+DAd
aB+bY7PGo5qHhAT5Mt/RqSzxZAtMZTzGO2c2Lk+Ce9KsqydEwCCTGj/OWeMj
Tvg4cnA1PzZZI2iPPGkZCvSVkdudS6plECG3VlyhUmTC5eFEsIUJNfTgPj59
KI3jogETh8G8hEHkoiacCX0wsP0dK1cZ3KdTkT60mw62vptxD/g0O4tPykGG
td8f1rVuPP3qBazc4DdQK+NMpFV9WyCr9uVrlYCrUNuNvmahNX2VDYnzWUuH
30+WANQ/6Elb5SHYVE1NwnFB/n4jqzee+D34oM8x1tC+QtgVhxC05FyD8phb
/oXgMJf6mUWlXIUfRgBabYi/CV4IvEYPZMII5EV4aghtkY6hn2fOMKloXOGp
dV+dN4VEF7sjVFpGWM/pfZ+cRf35ttNv/ZV9LSIWrrNIYdJEtQ1vG553gwzw
W9345qG9FlrDlFo9JCQVl7ng+sb366xEfjA7VtiMCuxegJu1317h8n/4Db1s
JEnfMeVevTOYkoGO7ABTfr7Wt8/RZ5iL1AprrjfNrHMX9X3FTXsJ1pk/7v/G
fZoaZxTJQCYhp8wGQML7MagFOClFJ3g6vFag36lYN6Tx/mzk6AJkqeYErEi9
nNmt33xY6Nf9tPDvKrM3saE3jhgZBYWPCN7JbdmO/5b1osTNLiWdt5b2YI9J
2hmKV6bmS3TbJPJ0BiZihslZW5C+z68yZyrn2vJ8n5X7Vp7lD/EG7OyMypRF
2NB6Er3oY4CmTVCWF11EAOsIsAORTIZLj8SRMBlXss25Wjvi1boB1wewAKYE
jeir0gajxtkzWI06zwBR5JK7yn3/DK/UiCeFuLW4eHot33Znb1Za1RmJzzEF
UbHrkzyOMs4C+oN1650Eo/PefGliIduKkZyJ3Tdxi06AimMQcO/rQImprZJp
iQ6N0VMaKgXQBr/kUl7DUW4dWwRVF11IIrBjSX5hHhqZ26eJPkVL25XevQIC
CcrNeOfN8Y2psVoWU8ereYiAyjHdmDfL7vv5D6ICdLHNvRCFBOllMZyBIsGQ
PwUFBM3xsCE1J4bCrM27acy6sm9mprATR5ZN4TZC3+ZoCpClsWPGj1FssARi
w4ndbbgkw1wL0K+pO+KRagMFZMfiGSc0NMKVUPa28KrPxno/v/qKSkmmbBn2
BNuWVqNudMRiIGJmNylPipyBa1Oq7RsiIyhuxEx4XfPGbuiajcinfoOlZwWF
nOUE48t1hdA8QIQdXXX/VPfk3gtB1N+IrYo4hBicYXFnZnn68qJnohgxEkov
lMF1Xnzk81I0nVz9W/iIHOQdCcGDoZOncHc+kxxXVImbpaFRcBWczuB0Az38
6LWUsD9wkCUdUce15i6jJXUnfU7Z8MLREND8MBfWIMRlGLeTrcE2g3PtvzFX
khG55aEM4aaJwBUiqEYWYI6HsiHopP+m9r0gyqi8DYaE9jHA20kwIzzD/qD+
N+m1EtLGXEyiAdUCAmuf63uUgZxObcxwyzabYK+TIdBpEiZ9Jqm8dqicGvqH
bM/Ksu1HGmL67I9sdsAC37OUgqi+kw8VZbxvDSn/4A4z2bBWAjC20K1BXhGx
9tknE9ze3ta6fvHzQDIZ3awv2ZDU3hPu2WfC6F3Rgl0wWRBGdZGp90qlWpzW
t/7PWF7F/K0oNe566glZGVYpwh2JcPFxmQqmOPtauD7jHsfa4TvDr6OXyrxi
9VzQtvk4wKzYeNFUBuAtSJ96OXocIbzghnVzto+DTgRaUeNY7qO9Rf5POR/I
zYdAneAKjWTWhJ/r99swAlu2L9jMTjxfIN5Fs+8BT3wv5fgKVS0Wc2ifX2J8
9je89ZVqfXtNs+Juc9NMMi7uv7oxwXo/jUgGpRZwXgwftb0j/Y3ktDgLmdYS
wjJEgTpt6ot31JRrvOPCFq8sljY8/doclfTT0kq0WQiKVXlQ6HvnoTiYpHB2
qQi0m2CRt7pUjjdHo0MYc988BmniUK8RSD3u2GtYzxxOnNNfLCX7q9yiLMYd
pQkdv8+xjnFSx6KKnI/wR19uOtOwnZn3WfjZEVCrqdvvNRVlVk+UqEgRuPZ9
h+nEnkqRyBhMJpAqLTzXKZ40H4JhyxWNgGE6Xi9idasKabDBlmZHp+dYe6nb
Srbx9/xuuUwgjwoBU5MouzLD5YXUjPqGiIVVn5ixEEsmW48V10SEuyGbaKoj
xQvBIP8foAOYbDf5oryBOo+ddV34l0CeMwlz/b5oaKNUQszdXFDFBGBQbBgm
+fjCoadqC0XyQEwvgvPij0rK66Dmwab6FTCY4xmssQYkMoYHMyjntXjx/yuY
0y91av5jTuXB1y53LZQNguNmgMwjVav5yYOB/p9MNaD5uZ/wolBaww7ijodU
3wMwIxOaSik02XOWoTOsi68c7BUyrxEMtDxvyCZhZO0KHMtgIwO1S0Q0LbYL
W+KVXAUpMuZrDepSyRYFvuuyATD6V63ZFp0zOEHrNjCXJBBVpIIZJPniriGY
oopaVCqbLF1unvrh0JQyzUDpsbbH0jzBDMqBdnDsG+43wqWYdadRETRYk3ys
Hl03xK2l7LaPmR2s1SDerbLqmWjqM3I/2vZQj3nav73yWyECVJthOf1RqAho
tB4fRvYQ0WgqWH7M3Ej6ylNd6kEWIsbwb57+uD8TAR5V3jfYvP6tXLGUEsNA
hS61TH6NS6Q5VzafdruDW0MI7+Y7+Tj3kaxidQSZXe7uvPpmBgIY4SV/0h9I
sZ0EzXKO+Ohc8yn9pMhTelPTFSQVjm8St+h4EfXP8J+UXB11RfQhE6KV8jbQ
3Gl2n40A5hOo1VUlGg4vEHbjfeeXWWv7+ZxGmGYQ0FAFiV4GAHnrFtO7Ydx0
Evun2pgRF2legSQAuZxTrK5NffgUomYnBqjIKXnDFmFQK1y5gIEBTHbEW08H
QzaxPZcG8W1zRvJbhuo2S5jmrOR6REBZtxy7yI5YEMn254tnhlJxAkHP0FEX
Xjh/u7nST/Z2o+OibYbU1YHwFoflzelbt+ICu+avZrA2leKBRyzZIDKb6xEe
L/7Wxl0hpwvw8WW0NRaZtJSEp/te2q7DyEw6rdTCUzHp5YubdiEFUPkqdpYi
LXIhjMqkNzoAi7YlMwV6YG6p+gThlTCG7sfCP4ObGkkOp4TaA6Ln877qRThQ
nJ8xtB9s8Y08XCf1qXWc5O9j69lRbui4BFbjdm8jFjZ9xtjbg+tNjXA+vlMt
pev43ZEinxRnfNsVUrVqFNPNByEDB9DsVWB1jEar+/l7Ai+Ef0yPtFTxM1GR
9wuSlmITE8Q9Jwv09+LIZtGWg0kpEfWgcM7CxMaT1Ss99xqb+8X+FVJ1s12e
kWvskaTmSopBLoio80GVqX7tO6oarWfIysHBB3aqpHSRhaxGovzpJjvOwm7h
zv5aoUIBKQiKYpQXE3iBsGvBeYkiyt0jy9lFG0EPIkfFav3RwU0C/4J1toe6
R6j/UWkTH6rbQi+UrRYCLE4rMUHJP9/yxZZORVNmzCbyb5jB/sz1jAJia8x8
TtAyJ755PjRMfz/klvg2WvXPJfnt8wAhjTm3UBUiWwrcOpkEM1/6TscyYIeK
I+FrgvjzekPA4kjuJA9IJ8SsiZngt0bWIo842Xcb/t8x7DH0g6kgIi9waoq2
FI3HQSRCmSS82Sviwij1e/R4s/VRPIgxcRoRSqkxDFEbK2ijnw/LVuGUgBPQ
WxyzjewkkX3gFn8YQ93Qk4QZFr6UZvTQf5e3ueKBpH5j+/5BKxLnAjNXPZ7A
4bD4clTw2NfI/WkUph/Alz9FjbzHd5SI7xkft8jC7B4iS0saFNMZUmFWi8hB
va/u7j6/hTPvag8WxRUR+04bdqmGNafxDGQ5mMSKWAJUWeN7THPK5+tt/9mm
b8UVCMyNX7iJvxNHnOScbMbxEAekKx99Z4cPj8HIDeVlKOSQwT4BBu7qFL9v
jHWmoIVY/kKLMXXujUEwI7dDOIcdugYLXmVJ5mUoXl05XWsRLXjZRjxYM8WW
Fczkdv9O8ithyyq+VQdrLvBeeY8t6JyVn0SPFL/tH0eqfQIpAyHCYyH1WbsG
oGj7q4vK2lHf5L94eVXMiPnUSXcCkaOUbjo4NiiCCk+rSe3rTDbokCkrM5IL
WUJJW2iID6K6bqNko/VT+2efjvNXrb1Nuz3ZNNLbpqg1yz6z4ufW+Osrvqm3
pzquvY9LyXina0svaErmWpddGy37HRHrYhJteULEeZdhuP379RX5yctCNsLq
xAwILneGCFtrgwwXbrAJjvVvAW0a7wmmwx/IWJ2xNYG0e4woRwog1JXXV+Aa
uqXIvjKJEpOFumsl2UyxnRCCKi59Ytx7k+ufivdh1k5yWSLHYSHuHCDgeHBA
qf6cc4A8A197n6AtRuZZbf225cP0fjrmCxym2njokTsRPcNx8DYVyb8eBwpf
AfPkBbI7Xs3QsQjDFZoFAHEL5Ud5AzX6ggkKfQ2304uURV5NoGJdrrjVsO6v
PXO0EobPeTDt5k4Mjb8sP++Zt1i2nn2Jz3tvSJp7BaZivo2xzoEcAipvUxGh
U1HaZoZl5SCnYGpYpdFZ9O0Qto0pbnjOcHaTGRtNt02BeshkhygDluD1dD1J
IzweuxSRl62uZrYsi5TkD2jkUPc5LST4/lLu/OhyxktrcP7Fl8IhQTQpALu0
aW/QDER3oQ5+JYthCDW2DGTAK3p+KR9m+MW1S103t2HlSt7QVRkGcvWcSsR5
8wRNWgJNNFlAwjhKmABF2J5f4d6nIK3kJ5IZd4e8fUY3XFsVWCQtz2FHNPjF
muvo1ql/b/YRZwcr/2H9xCOvzKk2Y6P6QlzTHT4YwgCHH045ydi3feVbtjB3
BAn6Trhv39hIKQb1nYlYxA62R1B+TYcWd/6XeNQqnMAbrj/2CwpIhDDY9kY4
a9zMia3kT03KkQUTrtLAZv4nkNJ7i38EciFwhoTcbPKFA4KVCzpcQiTpElHq
9l1f/550Ayc4ymjrPRMbRWbJsgJOgBZGBV25QnfTUXH850YpMG8SRXe0MSvS
zDM9+KB+NSmnaZYj6qzcXLfrk8Y6fGrtJeFNtNAachYL9DR7VEpmumRwagn4
LdPhSpue0/w3AjCBy5xLB7AUByzi53MFqg+CWeJB72mtx/z/LFCIRa2/9FTP
jZvMM79RrIKFFc54+U8v4ir0d/5NxzXVTngMasU++kTjHXhEeZ+CdGCgrq3s
Fh6SiGvh08GsI0C4xIWNq7d7XHZjm7c97Nmk9Ii23eOaU2VBJYfZ7cCuo91C
06rspfrvSIfrSOmXGw3ygn2dIWIhotKmslYSxof/pCgJBD8EXQFapG3gwtH3
6jYK8+bWAjct+W/L0mLqRpv8V+bT1GY9h6UZ0baXvnVg3PC49JXr71KMSIhv
n6tHVT5Bu42+BZYJYUTY6jUSu+qGzayBufzvIyVaxabrbWlybg+3llMZdGis
4EwK2ywjitYavR3jTXTBvq2PC6vZ+9+rRAAJvaRo0f5aZYITDXL7wEPK1fKb
EXyU4c3ub9u+1L4Jd/c+I4zONcWrVOZh/vU4lgjBCajnkxvMFsN70IPVUMCW
PiaSOzZ1m0ort1TAOIcjTOAmCtycj9K0sKbYHE6jWLjB3tYmQd1GSV6rgqFJ
CYMhokI6ooFUQ36dObCSnBsMxqcRXPgC/fpSOpqETKkP8GDJ/3mTSmC504ih
kMHhpLZrkqNpV6WlGVlVT+l7yLj4xGWkA7nVbPXjRGU+WhXtbGT7m6xoHsZP
/TB0sN6yRPH+yn1ujSb8ngKT7THuL+uEvYP7TplOYgmTZxxkfHnmMC2+Koex
xc5HT/osbzHbwDu3aL3pzvkQ5oZG3bSte573IACw6KogjXxqLX1q/kwcSUi3
/PXdpf4egT8FS61YbepEMkPQBUVjyS8WgzFitLoM1yhiKjMLQhfkZgfJKQq4
yC6XoWnIdvNHxObCv4/qhzZJxzOvHSUXKqelc4LajABYtlpjlg+mHaJ6X8iL
bwM+6XWA2OwnduSwHkMficJo63hejOguqhH8Hndg1TU2XPx1TjMdJuxeB/BE
SHbj14mc3O/88h9HmVP3vMnXjygdNxRREFVBocZTQp24sH3bsCxzxzsSgEQX
CNOwxat8L1tQ2P3E7320CL2y6uBdolC+sR2EBbHldRPVjk++R6aWYSKVb/MV
90eErbYj6xiQxHZMnqW5SeRjB1szO0hGgNyTrz9ndpyTLS3lehdieuW8nrUk
2pZyESgyUX3qOSMmsBj9NCrcX/IPW7giiMxoHL0gN14AxrDIqaLW50eIz0Y3
6b2Ze+ZFXAU8gmmyujopbfv1B4TNeVeinDSAze2MID75pUKM5cW2q4rXSfS/
AsZ2lt1gF8ytjVzFJ/i1Yq8YYgrZq234Q9hy9dPf4f6ShV+m0U0jeIIdpxFh
rBdawoBKbdg0sACHCCW07AV1xKBk2H/FQ/35GM71fwmJS+SWM9Ab8r4uE9EK
YexfxwDuvwxWmRIRWJrycVCurZL8FYtTcrO+nomEyD6DvB2pI8K3yUWvbNZY
wzMz+Ex25nLQ/xqLfcIWJqvV2LOyWROsOgTAYkUcsR1+sRCDReTT3MogHKRU
anE3mawmAwN4E6kvRRPcBshYj5Nq0p3B6P37vnK1GiQfqrPs2WJgTCvKCi0N
bEOVzF88qjySZ5rA4sdyDYilr+PNWGWBF4e9/0rhmvxflNponBPqqCHXc2qD
YzHgL8zvtI3lugIQmjt+pu9kIPiGCQ6a5wuJW8cx1HbHaYhBLkpVICt6UC9x
TKGfLwNKoEMnIdwKlDX68dH6jhovy8fMAJ2hbdaCB5jE+dSPRSDKLrTJI3El
jw4h2KPBgZw6XlvCJmYEPHvHoZvRbI9+2uboqydw/Cw9//fqpz6wdeOAdsCw
0AHgfl/cEMuzd2M6dSNyz6A72oIUjcikbOI9qVVg50cth9hFk+ujcVqDA5an
q1+oRE0w4nQY73nIZ2v+ROEPCVBY2DPFvBnpHuU6EOCnLItoD6bSkDeIPzfy
n/kP8zOGXHGyK1mAaA7XRBeIv6a9QQ0BNJ/UutwDDq4Cc4gyotijPT4Ou0++
pEQK7JDWtMKtQaqOLDVPXdxoxi95kcqFGfr22RYooqxP+fqC5u7DypE+Aq0z
2xxaHSbMTeLVbkpG64d/MVRWcBITuqqHcJ9CGisoGnHvu59+6sL+RZpc6VSE
XcXmGYyJIuX/hpD9peRtEuXNd557jDC9H3PAijwXsXfECkCy3yPKL8SRue8J
fSfC9hcIbOqUmdr+tt/ewaWay0UFeh/JFVuJ+me263oZGJIcSvZ5wClkD+99
9UJgjdRfuiOL8ctrWY1wiieLQw+JufMhcFkkIaKH8ads0dvVXHo8aBznLmXM
ZXUZJYPuw8bHxnwayNnl+3ro4w4bxyI9iEFVgaVjnMhm6QMa8RZ/jMCDNvIr
G1TNB5Ntkq1qh4eUXf6zCtxLuaSJxOUDCIgBROzMWpHit/iwhQTigZ5jLnpM
YoY19u5wXX2umKsLUjOboku7tRxHmXYRj+4/j1VSP26IXpAM20ejVFROxttH
Wqgp1w3WISEf4Qnqypl5xkGgbfZA5yhNsxifINBYkYQol4Gof99/R5+AEpjx
fUrb0oySnYyrznc/k2XS+NF4k8ojB9nakeQvKF367M+mUd5rf/V1s9Nztx1N
s18SBQZIZPmjfiLZ2IjPrTlFlUIdJP7NJHzBt940KnG7Ajg3BWslK/IP8nhE
x9TUFsqB/559nMlcfIqENsWEzGO4i5Kx4pGG0GLz0DsCqgWzo+9oP0aGWRVQ
p4Gm6GzXa3LT8DtXWeOq7063O3t8X37jKSTVWLXEBOhHkGahoUa6Uh/S3LUs
fogi/edDOFq/xare4WD//Uy+6pJZI3ENLhyA5aXFvaLOXXjNmk+E6kfa5y4R
tEtra2SpoVnAO/w3m+YEGlUZaOAy3pA/u5iAE/Yd/hGXG0yU/gfDQ6hQ2yNX
1UJFjrpS4oBHOv1YVu/m7UfYAK2HovgJV74eL3lu29OUh0XQVT8ci4LkV6Kx
v/BcpRIGUXpFRneaQdSt+NZijYQ+GS1y7NW9xWiZhDbEpPaQ4ik0aO3rv0Lf
NNX+Ko4vEOX2SuaPnxBYWhGOZL8//JtfeRj+9Ha5G9YET24DGX0omy7MnELk
Z7JY3llIDE/z70wB15iKBIPNWNlyvo8UirQqMJjz9skp5V8+pqPVbghAASW7
32BwHrB2a4XaUGNxKD3REslcnUoWjwTvK2fWMfmuO4ze1VDlvGlyD4FcZJxZ
s/Gyh6PKvnNm9mj6ujxUQJfqVSAkmMOktS1xSVJjUdXz9IwfQQBShKKg4z6c
1bofhSjtd3lpbav2v7BF/emXro90wTJCTmr4cRNWNkREuUCIsWbrIZb5906g
kd7B5lDXv91XCHutVOifW7yB/3yN4rhM/0geqllOS4LsASfUKwvyuN/CbsHY
YwiC0zaWxbbU1lz/LkSuz/3RmjqQsbV440d+gKW6rjjM3lGwc7qUb0oKtGoI
umju5zZdjcusdXDi6SsnRPVIrzvKYm/ZZjxxwQSP4f41ZgSqE3zi38tmwI3X
S8aesQSCZ4xsPgTGueNtpUBsPCJaScKHNU5BRydpVeFwUT6HXms054P9C3oc
s0ibq9QWcq7Isdaoxs1dEqMCMchEkCixkHZq4RBjARQz61yN6o0xHk5BDqrD
ruSkWUHKlnJOY98PkUtz4BTdmm7u/4ewpkL8G6hXglXe42hFtgnGCGM63rbj
HtGcQBYhp1sNx5eBDJuuoZZ3egFQvaI0oxd7nylO+xHXSUHwlUUaX0E7rvG3
Efo+wVBFH7Pt4vmw6ebB+BvBfPe7prao/9ZsEV2Eya+2cqRNiSgulY75MZi0
De53flGk4Qp2OUbBtJSuuRtm+F0o1zDb098bY9ndKExcYHB7yvNqDUhfoPQm
7TNwTk0Qn4vFrP23COh06Qt3aWDNNKqe6aYJ0S7LI10ilTzzENk9kr554o8M
5JmtvGitjrvJViioaGjcbFW+zXP2yq56IIlH9eDSvFxYMdfsQwGGdNhiafhD
g0nj9MAECS8V4bomSxOs+RHvkopTb+LsYtXlUYXa47mOJdRAtBeT91c5KGr3
QMfCn8cA+sDm2lZudEcsWbAlSPv5fRa+mISTL0+s00a2e1hYoAHn93SOKb1A
o1gez1PXqUetStDY3FgpbQlHEeeVJRQY0I/bWY+UFH2l7h4C/SeBiH8oRwmW
3mKKSCAXw8XI1O/6/hkKsqOyQpKmZy/1Ci7ypYRwAx1Ep0AEyW4nWvBLYgMB
9TmDuq7jM/CbTpW9zFX91WhHnd/Gklx4WKUNUOIZl17lOnHqAxgCmku/Dt6A
SFKqnSrNrS43QH/d4Cn2PdkFkDaTan6PKbJatIrA4QOu6KhvDK3FHEr45cXI
nPLqxOYftLHT3HnuyOgCv5Cfwe5d6vOhnZ6hDk//aAQyKQdYugR+NnQRPWkE
yDRdMOZACE4izqH2KvGUJcQYMjYiT1o/3WOb1GAIcGfQTna/1edq3L8r0T6I
Fios5lOoM7WXxDjJ21E2CcpZILhFhcrJNbYjwaHCmaqMXex/WG5x1pQ+XB59
9eND0NAixxggK6yPd2/p2KOqlenFJh22Dq5b0nNUBF+PY8B8uhR9oZ9icrgG
HSci5yECwwTH86NJNL3EWnnzGyya4QypMGSxFz4rEm6a/Kh2DQHO6uVjuaiL
Xam+G4LRaALQOhT46nlnHq+SgGvZ/uqkSnoHUHDeVvMmVh1dBKriUImqA6PS
JYFqTv9IwTW2m/BU+yKrauiKVm2/UJmfeR65ZI+UYAOGJd2Bej/BV4sHoTe4
zM1g4RPFKQNjZIf/CqlzGsXpwUHpNsxW+Zwdmv2Etj4QpuZnKAf1F8C40lvx
hFA1KcaonwbGsKOubG3TsXqXshm6b947nbNNMqPL1LJZ+zYN6zYqKxnQa2Cu
f2HhemWgA+GF7+PaBYfGDNh7R0sXi5slSVirp0DUMqq8IaYx6emijYb2LKrY
zPDYSJWLO+tUNGqPIHYArN9H5TfcyLGsChouL+PJ5GXqniGj10f6mocawq/G
Dkd0VHoxtdzGyZVIDFwXBR7HcCkfsfTChzC26JOLPrbMNPLBncK8W2xqFMyu
0CGedySQ1PWH9Un353yQXgiNaEKfhffYI39eIzrx8b9Pr7t24EFBB1urvSQy
s+CSLRDYfu58Pir3DdFmv8hXczsB+f3TptOjcPjJ8elhKP14y+iFJYSSZvFA
1fMUgILSXz3kCYNN0SROW22OLtzKl/mLRSn6Lhs6dIyyAmFxXZEHhvtXF+P/
xLhNQGN6M7r/jcFQQxkbL1+xk9YuIoE9zvQ7ssk3/6+X1vUqE7n78hOeMwIv
PaVpuGuldz3hEMybuQ/6Jw5C73lVe2b79CLI8ZBosBCL0SJN3nkL2UXLuHTy
+cY0lRVSUs+QtOiEFhWL2Q7iKs0SwmO3IaeK7VaqcKNJA5mJKlEUSdtOxeV9
TjvqDj/ZiANesztqCMdETZULUTJmqJb7+bxsufBKNLr0RCieDcCvE2O+45g6
BGfep2F0MXzBmvptsZ7gWGUOKFvf/BvJGvnGTJgKIqlU2PCVuE+OVgYKurQB
rTSSiQn+ydxoeE9aiaOLrlxgaINwJR737mMnvWSB71S9iFr2zPMWLt6Pcssr
IX9kTO1KXGf9WiRkumcaYe/AIPTIo9D+CizjHsbD1VqLjBhjt2mnV85AJ98Y
pVA/NSjFd+GhYwy7V3itfNH9gU+H10iZ6Gc10gIIF5sNHEK3jOwXMIaRAj73
otm7oeOYhT0grQqIEJtMOqPwA299jmaCBkEzF63E7rnFMGuC+8qpslPDdB4Z
ptrEqivlBsth55X1ogFg7huKVz6HpdAdhGRSUWlsDmBSeiSTD4Ai6PaXDogw
d0At5pS+8jzHz0BtN+K6JDP+CUqOBJiDIQUE5oAlhxKifcCPcV46Fu9NsgDu
YJr2grYs27xIuH6YUo6/DyxUdCo3ekuoOzdHTIt43znNt/+bjLKFL3N0ZXuS
DqrqMs0v0uT7VjWOhWkNp4bdSIIg1aPb7fz7ZsG0owoloRsTtvKcMr6wTxeL
8ELoxUqGGCzO9GIy/frlHnFxAkKdR++bj0kUTLkmkhhf4qdzRKjOM6ukoxw/
O+SfHEylwbp7V0HOMSEUBt3E1MSJRwEMvFwh3YtCBPKrMrhTYOzgEb+jsxPF
W8bwnQfX5XxBFLAdyDMLdAPC10s+gvjxK0kFF+YhrLGYf4VmWM1WkamMPY80
FYvOqt+1woO5OEdehj5qyQ4Z98BNX+0G1V8nVGgfQ0JzvIZfvoqwUvWorAdy
2sYr8fkjtem7V6/oPD+ziyiRuuMxoaSBkGC6GVnNLtyHytjNBB7UkOYDDHbE
iuElLvPTP7lrLomiu0y3FSw5FTnOxJbf+cLaXF7rPaIZjQ3nvqJBcOubGFXJ
Fov/7rxxvkm6V345p0jHfxBJet5poH84IATh+7PzVs98nxrePCqhKbDR33fC
h9ugWlBjm135FsA66W/YTm1n2AGUPd19Yt4/Nf9bC6sCvc/Pz+PD7ON8wK7m
wB1Mj7TfIGtfXdG1Jow6Nvx2nMfbAPaCUYLM8epEF1heL15Nj4zxnzyeJugW
S+KxasHlRd4fkwQS/0/95tvpQN9ogKau2oblrLkZsbunbLeCgrKY6HgRnTnv
4EjQeOadxTPq50Gcs2lC0sazJ9FKCAcpzGtwkBT+Tz+W83Il2i1adYlwTlGW
Fa6aHDq9roddX5cgn0oarDO2eAqWQqQfcEo/bgPt0qBY1kpOMtRknLeRTJpu
CR1kPwgnNDwWVa4b1qv9oKzcimHVoAJuXmsGCZnC+5qXFMNzMlCyQXp80WX9
si363zjoqDc/DpgG50rWnSat5LMP0y1peeSk40v8LdJyrJ7CGzdFq5XH+0rx
TtmTvYp62LoZaNS+jzv7kXzojIHzfro0YOO2JSWueuA44FhWTiaagfqNdMib
nxke3PxnpRtfr354RjsTjWfnSiHF0gmGcsziUqbSCykWbecJB0LLP8SS/Xzw
jgSCDRKGzlB/bfSMHHitm8ERAGAkr8grPB6u4x7qE0oCFit/g2sD1a32YvKT
CoB+0mSzoq/wZgpPO+jHxnr3q2UTF6j4oJH1ML4OmnUuFQzgOgRUnFwHTKgG
93W15OvPMtwEDG3g/ib5/7yazAOGrZ6QhgPBV7mPCFGZj80K10eO4/aFloxu
Rsm5BIBxITpt4rOlD0iZKsxe2z2n77w5dQw6GuZyM8o/gK5r45dJVpixsPtm
wxvaeptVHoeiRF73lgjELH4Afe1s0HGZqbQO++lmKAewL7OBkf7awtcVN1b2
sWvEypACXO3iwlnscPhyd26KyqeuOYzRozI3VPG7hhcl42gdZkW4Jsov/WTr
meb0bhlvTIbrDVzhN9F+AA9NIo+xT3wwW8RxzW+xBUrPhzKimqeXpIdpR9+M
HSy0IDKdi/miFDJfccVu5ds2yFMGDQvGIih9O3K2I/FR2H1GzB0CwSqE/m60
3DeOjoM2klzDV9lfJ2HER3mWcot3cRWipHVeooo56A4aW1G5V2OOy69xUvk+
/0xUdqo/viU9pb83cMBIGpYnuzcT6rMJp1d+ytNJeuOWLOcsUeWRll/nFV94
1C2W6R8CQ8uLIeLS6KBdKeqzUexmLswoH2cIVBdRWxUUgpHbDjoPnxFzdHN/
ucZSM1t9HxPREjOxZFQWvMPgoZJLfnvlfURdo3NcRZChukEmTYtvHSDkU0Wy
H5WiTstgYs3IGTGapofDZrhotaPw72y3vN69In6nSA/clD4a7HKL3lgZP9vs
DoXvUiP/0dn9XK3raKZzx+bxdZ6RQC9DGwnPBOUSf81Zb9vOkeTxXuus4zNi
/JH/umCiluw4LhDq8T2VMUTJwcbl6E6o3I/RMBTCYLYTKphxZcH61h19YqwV
tU+6V3+Z9/WoDC0vO35gLrPkMOt6pHEFKRf1hh/hqD4wm23twL55hoBu6J1k
8fFHJFcknGIgjzoX0yoJLIcikoM+f1OFsEjZv6PPIsYupDU5d/noY7BrpoLs
ypXjpg7g9lu6BTZcyFu2WEkDp8528g2xeGJKn7kJUc2EeP38G2dEbYJpJegF
lZ++ZAYpgDZaLi+veu2BSnsXM75MaBpfDMRUhypUsoXgNGstjXC6kxtjTmEZ
fWRjr+lqBv1e7HMi5FiCFLgyKkdlffuSJigeHlsotDqiarfImfXcgbZcR7k6
esZpXUPg9CzfDvOS7Scl2GNk+FhVXWELDUcjVbOfTBgZHhhvVZZT2iauGKux
EGVlOXx55DoIxVXLx1mDlOYg70LgVVcFoO11g1KMWvyOUdEYa2Uoq6PLmeUa
IpCgNbMhj1ffcEbZ9UEFCCkee7jr4mdV1xad2Do+yugkZI8aKDeE+9cr5Wnh
T8eMcl1Ptn3KETU/HE8+aFmvTFUqE8e4NSCznECJYIQZuI/s/dS/B17pO2s4
YwGEu+wcPtHF7ZbOlawSdxdY/YX6T8LWJ9M8DqfC46WJMHOLKE9GPcIdoyWY
+RgT9yHx37ggXFY8gLozDsBD4T6wNnIQl1PLQZoYJ5KOEIqWvITkmCF/DE+F
6L74irrZbY2BloDc4gBfbKCApGE511LUYMWtDUiT93LT2V8BrtgQY/A2trez
e6Js7Ou/1QxEx7ia7sq7168+zBmgz47TZt/XN9GcAXyn5l1sHbDABrG+QgbJ
5TNtqLwDvAOE6w5JfG3US58STdEAwhbEs1T1VhEe2xkHjfyTIIjzO74rpYRv
8DWxBVDRMS9wHVJf+8BkRRo8mOy6y94qScG0NxzMq9uW6rs/N+fPK7c6Hw2A
Pk5z4TrGYRIU+GISXFSxBesHf7pnUyWQm0tuXQGVYPIMcSghbPKrNuLNvBwV
VwHEOF9kLKLoFY3jTgkCWdUawnEw3JBP0jyv80gICgrCb3X1ljynQJVx0sOM
I8zSMmlW6rgrEW2/lZKcua/xbJsTnyD+5z3JiNq6nQKkLGC84J10saJL39HP
yaIHHxpJe6nIgaZW+EmlT3Ds0rf5Fb8s8EUQjGNKxGnC1H1fav3RhtgmBSR5
ueEq/S/iLk8OE6L+68x2g7CofruCzOWybYYTB/Gt7pmnTTdGYkHICUMH3/fO
N2Pc/3ImhPTvYOOjeP1A/JWsnlUq+zbi1XXCBfyX4vG8f7XR/o7bgtFGnHkP
0sEP+D669iurHuxh9j/31YfJ9kRUH3RR0LK2tnAI13hbwB8ekIZohkOZ+KNE
bjBqszK+L/pi99V65IstxsQk1NvXm3C4FvJUgjs9fca+GaByuEkW2T56A7aQ
rqRlWoA8RD1Cir5m8DsXdE5s3eCR591GBm8NfzxQcjz6ci655VophPE0+TWy
UW4KmEgrdy2+gz/yUU2kgr9gz3yWZUQsHYZXYwrGKV0IAxLe3xvEBf6nD+J3
R6TzKLhxC336BlJJDt1BquNloZTZBB5EFxVsZXHAIycar+TT3mhn/LcoTDzI
K66t5x5b5fXcirzQPotlcSLUGKegpf7mUw3E5k/EQb5frdvdJDM6SMK8xm5R
vdMdbtrejZw634xeaCKWB8FskXluUP8bKnIGzAgSOO29dEWz66wJjjf9HBxW
6f9FJA9u//WafcUy1zev1AZHp808M+mKiYmh8BPNAgwNafnrokThz/BNZFhp
Y3zGdHYtEeRiaTzFXHz7zui8SFjTs3VgnDiOlgfnHzes1aiYVLB65nBfkoch
iOuBJnsDbJaRf0CZYl+6AtYhjm8pzQS+6utTzCM0kOokvTyDoDFV5l3y7AEF
CN6My55CAEXBl3lhA7J3YTKIyellnGUHl4yEFHsxuz/tSfG8tFDb8RG30b/o
JbiF1B+/3b1b/Hk+vlGYdM6GQM8hTmEUsGSZA0F/q8DsnFCysbDbsH+zjhHg
bsHnkJscbPYygpnMuds3y2rQgotny96Pelua7il8cZzXzwjUk9qNxhV23GEn
De4IWcrb8Plr/emVXEgEdb9MYYkB9Mt7LRBpM1qp52kFyUhj78whaVEogiLh
S9BAwuYepGWOmYhfCRivjhSncEN4WzLTEDhNsAY263AeQNtPv5Bdw5Y4/ubh
3Mz1OIE0YiUkg0xAp2619jQAAcY/P0hGTCgXgivPt16OYZT1hQxbTVId7iDi
o2nXS+PYD/HoWvXO7+2MImu7SdDYDJjzlXFrI9HPC91JJl61SeL14u03++ov
2PjEhGjV7Ewmkv9loi30YgOfNA1sMOhALFCO17ZqTFMeQ45fgitjZX6y9QM8
wheiKsI65vq8QLNE8Kg/ENcwjvjtw3kDO02f+1HTiifcsDEGU6+FUzEcWSvU
3xUKDdAewt7FGeKF5rRwf/vOGvisALsB/SOfsDs0IHVCdtF5IVwWVppCyBj6
bQ71yxefjfzaEbfMeRD/tJYe7eyZC0TWuAWRgdGnxJdnW39nRZzSb6Az4gRL
CXnXwe2ShFG/2+wBQJZMfiwSqb6l0ah3VAQ/LFlqA0keqochKLnKLAam+jcC
tE+18iQjczg4wTvSnUBAPnVQlm4pWO4OPMTvzO0dDrVfogJTtIhrRo3+4D06
+9+JQB/f80Ta9RiFWds/mRK+xnxYRYUgSfEqfJcWNhuF3ik8Vo7aNpMrnfBo
ivRko6FC5OJs60/oVECka8CYVmeF23ae5kiea2YYfbYPBklC+mAde2HqNUvU
eb7rAVStBZHJ0bLQCLCJlOaAObhoagtwFhd2xYlfrb5IU3UkXUJwFnAvqsE2
pTFWEaRi3lrhSY6J9WpvgtJv52kIjev8yYKHNC7I7+uDd/SIgnTjGYmUUa3D
8uClgCXHoy0h9oCiOtfaAOumyloCRVBfMduQOCQEtH2cMaJEselClRTr4EL5
ERL67u6y903d8FtYBUcRPYXUIpZb3mgpFqiEGry8ovSGSqSclLUjxDdJs71R
gU5XAQZxsKSj8/bjCGpK/PW4UXEFr4i3GZ95ckS1/dRABzHX7bDtiAQ7ZOib
eyv0ISVddrnNHFC+zt3Nb2YhxeJoYrjV0WhjzaWcUXiW9dnEELEkcxJoSV8m
g8UGiBJhpbdDLiePxf79VAWdJGbDIloH3BkQpXytenEcE/JI+gHs2jqQQpWK
+ffngcY4KxsXvTdrwfrMXwhYjMMBCz1IJ0+YgfS91aNGkar7/sICkWfTZ/91
tQ77f6c73WuDCQc2zNsBj9EMh1l6YUHPXQ+lrOWi1e/o5EqFW8zLfMoLGHQ2
ozeuypo58LZeYDJGPeBvWF3POH6KomnIuN47kvBqjJkyhEo2qm7jCITGEq2q
UOL//Um0cHFdFWsOrIu+fUG4I60ykSXzrgBje4OTB13aRI8wpLrCFmjfIEp/
NZA1xbicYX1wmgFdevsBB4nCft10SSvxZHdoBTmnDlsvxhItPMUM4ckRQruZ
v8WsNQOFV57dvu56Eju3zgKiR4tCWGXpxYv+2RSI9ZUf2Lji0tZDd5DXeDdZ
5hZZ69Mgbya/3r14FP2D2F2wYAC6KooXdgkicJ3KxqrcfYSJ49MxyLdOkLNG
IBFJv523c1OE3NiVDoqLc1phrmVJdrWWap3jzlzms6PNaVbYQGOwHm39IKdd
rySedUQ6wjO5DzzZhnZhTdaHiRsZf/dwx8IaUuRquEDfYKD0WJxMptqPGWw7
NneVuTH8qTgG8KUuN3nHDWhmoscTqG/p/KuwgEYGk98JTSubPHUnftEq70od
ETYvHuxzpLz5Yah+h2aX066xytbwhPEXvUEOsXeVijGhyTjixiYo6ZE2EYuy
ndqJ6zbuBsZg3CZojKEiKAORe6vUjFWnN7ALR6ud91ckUE2B1Jq1T7f7dx+Q
ThvWEXnEgjPoNUMMfCj5x5bBRYEP6c+uQKhbFXF3LOfz/X6b4S9X46/XlKqj
Hc83le0tYlnI783Q99XtRMSMMHQWHqFpqFaTxpx6zgs8SCN8oxZ1FEOmigeP
cJB7sjCL+g/m0yphuArrnH15IWMZdysVXgP25cIduYe9pssSoapOGSlX1aeF
zcS/rfMl276a23DW1Ro3sxIAX8ql4+M6QJUYvFr9tfSg5/2vC/fW0ryi4FHN
IZC49Z9XeuAvMUnRRYGNcyQ5q097wOiHvM+4hOwELLze27UpDeLE34OxmOTL
50bu49QU6ZZVXn1TRlGZinOzJmUzdKRCIndL52msipqHb9Qc1h5Ch/e0xrBa
n6NB184QITFIkrPk54Un/eASUlStsbdNdTpTdYELFLR63Xa9/pp58A4lOolS
+fOs4jSLNOr9PM/UXGQ/7ytEaLSWHpaAHyOdvCGtlFUt+Do72BJ2HsCUdhyo
CwVaIAcjmwMC7i0BlD8dyyXqg8N62ydZ0hoIYeRIUFgkP/oKmlC4rVrboVl5
xKggmZiOt+XncUpV2VJqgLGj1SPxRdof3KKAscQ8VladlaLEqOfck5OqY5ee
PZLilKNqnnt24fLLNSKuA4SmjjduR4yXiy6hmP7Cu/2i4ky6mokBi/aOYUIF
r//ZFpFNaPfl1rbCIuym5ERO1nIYCvLUI0hN3NTJSEzqYftQmaBsjfWuYdBK
JaycmQE6OkkYUhtOAv2MZqPhUZtyaJV+l7PvsWPaLOG193E3nzSlokCF6Oh+
xXtxmoVY28sqGPV8RQW28VYDv1UoMOLACbM+fBZQo4xpM0rQMuE2ZSre9kt5
nK0RtCIDSrMVhO62J4ZPgXLUYu1Hf7Yy3ZdWBj4sdt3eLKR0EvXvBe4f1ueF
Mlk4Y0SGGyTzjj2ErOL7RJ68r0KwOd5tCBb7grTs677gTWP3N6mdcSLa6hES
MM9HMaZL9T/DVgqmKrGMtUO6sGH8TFaYwZ/dlo2+Spv0iW/J/ABfoG1P7sQY
ai1XNvlgv/8N8CdHoGiGUdFMcXSoATrjnMb+69RBDoq67AqHLvdwuJTiot0i
KcICIqV+0WiDXjOMT/qCDGl+r/u8rtvCbZkKyTioqbT2kWgrH3ocdOE9KcSm
ElPAEdQ2Xl2Fmnm6SE3ImdiM1mV6I2WwjIL/Bu3roOc+U6OdHQGBaJSkcZY7
z0xHUmeeK6Jw5S1tBA6ZCzWffY1pRLFtEmyxtXeje5f9bWPKukc1FPm+52eT
OUaiVaycbg0FfoAJfqjV77/YGxaQhyPk67P8HSEqZLIPxsbVtloCqaqF7OZX
+dxndjAr3kRpjuQTAP7LNQ6/t5iuiAuZuwrkMjt42zj3WwMFbn1lfdDYS24Y
AF9Eu88KtnwmwMDrvu92BrZ+7LhAKo9yde4aSO407DHnqEfbCzwOhfCPLQIv
p+84H9olclWkesfvba82A5UBejz1TllolMEoXe9J36iS5tk4kFeNVdzv/EZG
NELpTZKMec75qJXXUGPcsQzuJ0IoyoRE7605LVpxkP485mw21tDwgypXSmab
QDn1Z7ROCjkrsdm90Z3eaCAow1iLCBbVPdj4o68DQGizad5JcUSSXtLepWKX
m2mh00Jum4EFm/9Imzl82q11IwwinpjCd1KPsiT5Vfcu5/zXV95xISjORdsy
i+HR8jJsy1n2inZAmiJRMK4fWQ2CekOgOfGvRJ6F85Dy00kEHvX/HDFWD3D+
h46iGH8LTkwqMc7vxFVTRPY/ANVh9tPelwZwt7yR488ORDExVPP+/7EmKpFM
rct98ecNmTp2mNP8Dc/TRl+zVKJmZuoy+Gxar7yhNxpLjZc13NyfpW+n4deG
okG0jK9SFKhSRxLU+m/YIx8d5Ao2WAJJul4tZS2u2fKilDH7FNyLFrQm8GEA
vFUe/l70KKdp/3A3oXsIfpRxtpbuXeKMdd1w1T7dmgo3gVvtjxrliffVsX6+
fke2yz74JEPUYZQJGdh09H5a2hbQPoxK+f70NBcTW0CmHtcMnB6zxzUpcN82
XSrKfpCo0gqY4aV1xNhgQVsdTl1rhwV/rRnt8xXdOJ2vmhOAJOIT9VUD/nKg
XwVj871l9V/y0E01FvRECtYbUsXZUzyXYVcWG6C02cwddNXqzI3xUqBdt/Mt
cw8cNk5rE7u6NYgAfZD4Pt2L2n/rjxqpwB3ciST0ABtvJsmGPKKiNry6Dptq
kpm74jB4EvkIoVCh2TMTrZ8r7TxBXzCqkkWudqdmUhtANJM1EjVlx8r25ML6
7ZSrlBR18IAvXbKantXZEsDa4qlrDUDiBppPvJgBW5eaairtkDSJC6r2SDSv
q5xyFKkJ2ul3F18N35Me3yQ+vJzKNb/LR5t/46L3WxHVw/Oio29b7gKtXVhf
nIGXMe7UsPAgrPvgeh04s4SRYbvcBwCPr9v/H5FG/ccbToipWdGcaYk53nup
wahnwv1m7SddS/X16FnoABy5rngiF2TCOJdmAwPK+ZgPtCXWXa+tqXpCu4Oy
q1chHHTfefVDBsLJph0HBOP5OUqkFtAuY6aMoChKJeMRzMWWYkHSVBaesY5v
8zsXdgcDn6pAkKQ9O8IyTux7gVRuoacXtiufhNEm1mW9aJh8wkem3Zeuih0A
UMYNfCRX0s5NnBFqxEvO2JPq9lsBWC92idjvDQRhHUfWR7WI+2HYU0rIZ2B2
/LfJVYNhJmramRGs/4ClqCkUkjpNisEj+gU3khELlW1AjWxv1Mk7wqDS/Yek
X7eMJDQR9LzbeydjdmWvEWjmMZFAuwDDaNlFTMpZZIh3EA4PAQ63Wd07aZnZ
nr2d4fQUjYloIbKpwqehPpGFBrY6DavfxE0Ts8B+B6vEO/iYId+bxIRQMuTP
8pmC2lCSIEJXgMyA3WpgiFcuLbsDQvIt6a+J2cftuwesl/R/2iryaJMIAFUq
vpQ/wHe4G7MO4chpO316ytdlLId66tOKgir60BwqcJV50VfJnzdMopgAoHWC
J48zIY9BkLtCUpY6QsQc6SQaVtrxUOsHGhndHBTdqQLlU2wps3eUj9Vrq+iN
4h+qyBij9LjsHjdMAadKNdS/kYfURB1B9qM0Yvl49ATk9WGW5gN0Ar8ERe2N
2AeRHpMGx5xZwbHQRwR87+yyCC8aEnz3hkF7CD19WHLbAPhrjTS0M9EM3Eu0
5uCLNq5WN5qeGWg0z6k50wn3CtStjbEbCD655rvusuBJFJWk0hdxuGf5riem
dav3ZtYJ6pasq/OEMrP2hpXNaFBr6+UiZKXgAHO/gFIodgbDPsK1HzATw0RV
30qw4eleDqpGECEmhob/jh+pa0YSGIwp5WjQPLldx2LzAjJ0srEFuTnHbdml
1S7qYOWmCUBRC0/osKORwE3Sy68iI88lKSZrCbC6tlrRM4Gc4tGxK6X4Y0Nj
qABnEnnX9HRJ/yVQdm0y55euV4eWg6fX3yodFOi1XodKpgVtqRrqURireATp
UyL1osr+ymxLLm47Fwftv0q86VlekNc+aZQliGKs0iB7KvbR/rWfZkH5xMEB
IIhzmIdhbh5aqFbzuIgWs5eknBHsl2WOv9B/0zRQDbEQ/fKytrqmMnbRU+vk
hlylgaeTrrCLRta4hUXnkmgKt16guXdBJcB3utnBmVqtn9phHO4MLR66MUPP
3DmOxqqPVR1g8KZDSbQW4v1CZAyy3+GWte09sFcPK1GUPWeob0DAW038xOyj
gjMefCFqcLQJRMCPvL93fzapJTomNS8gs3WX5twRanw78ZJJ0qi5gdXzD2B3
wCyc25aKFfQkvov6fBL3ka+ZjvfmT1hDuneJQcSXAnR2FJeifdxkAb1iRmzY
x52LXChBhrQRe3j0g2ka7ayoQZv/02q8GPCAqN3ySeEL2unvkYL4pH26s5sd
WUPuVOufH28b2kCq4gQ4o4SJVDl9c7Pb/TWstRW0dtlOrYY6ZfJauT/32abh
yP8880B6MXPE74JmP9XxiDSr1dAKMEUwHHMDA9gp11Eh4nzGSylUtP4BCaRu
pUzyoKHVLRoBysAs9/Ev+ioXWNZO4+VzUctAFws54CTjkdH9ERgt7j/mIdIc
dMriXtKRJdOcjPJn5TnglZQdPkNFRZIoEKCAPgrCKDXZsiYH9Kkosjz0avNd
HL6RJMRolrg49y5o4szJmucVJMF1/VDp4/1rRArRZsiB2MandxtxYAENtz3+
hDiq2AN7BbvwR7TEkh2TKll7mRFS5sjFMrbwFNYu0pgj9bYa720DwrFqgHt8
JSQLFRwGDmLZUbvjlJ35p6LTWn2EI7j3sD5wN1seh3nJ6NpLiSHycpDNw9Oc
676BSXI2fTwo4rFybevegkh2QY0sHzryoqJe2v3nf2tdDKuvQQ0ILaaehI8Q
sPaH/z3VOdxiSktFWeleJPz8Xlp/gC982Tlpxa7gnFPZMtEL05lAoMuJBssi
2RAr6vbGzGz86ngi0Ose/fsmciMZVop2vcg6e+6RnvhSBax1k4W+Z6ES6s8j
AhGYnRhHwpa/Z9eq5Zocj+wVfp1YgCClJlSBh4D25R46Z2cc8INoTIs4mbaq
zIQieV2sOT2XS6xGEXtPqFHrsOMJXY0dCITaPGR1yXBP+6ebsTEig30JYkpb
SwkBWpv3jSXcaS3fZ1L/efwPdIc9GZ6SBfh1ZOdtStciiFHxeLkV7CckTthq
qdqsCgkhEdd6nTcDXszmZp47FVinJfzKN7YieKIixQVfoYUlyyh1SrQ4zqh8
w+3pNFlZinIVR0mMi/klrj1V6VQvqpQEXJnbwgkDo0yY0HR7zfXYV3h2j4Z9
Vy/TewICxD9i/rPsW2u2PBfwmEQX7YoQwWfru4ZYRi/LE9wwq775nJbCz4iK
jA3RKsALqy3KdSsLp1IhZMvUAmXCNq4mBNRPUT4CJLn6Ma3FREHKpfGxe95t
oCl0ZBOkas3fdN6xI3UglMCfsUbSSvSy1Lqe6v497y8jPwQU/MOLcnoUKSSn
Lvg3hSL03NkVA56O9KIDdo0fujyDzc5CIrIbDgSEDLcdS+i8MweyPKUuUad8
wPdsC/UdSRcExunmPjXXl6Cw9vPwgKKByiDREYQPYktuAXQIIUQUI7k90foC
nyn0IxmNAnfNgczTnHb8ctXtMTv/1hoMKeooEkWLbSc/DE6L4chMG2UMgEeh
ywVR/50OTHyw2Vo7zeNu/QOxfbysVwxRkbdUhTPLSVBnpijMbz7eIFF3+OyE
N3Phi8IR52DUHIpopWrqDpoW4OKSjI8isd3Fbse+At1cgKIUSn+U+5uAIHn6
YNBecIMPy+QXQPdJG5R5h5V7kCBSxoBB5cGoNhbzl7afjCSv6uZYdfVe0W9E
WkbMPJZCSbs/jwcs1Pck5mXlyKbuZ0ubV8SifZe3UowK+Xa7MGiG0xFX1+rv
htMDYSoq9CKVtPioZFkvcl28v/PH81BuSgKpciTS46GjBkIRGkaKvTO1aREB
srNc8JKb0hxGM3nWhOrsS5nI7g7AnWoHRjjsF46Jdlve4X5KIQwVf8qkPssK
kUY9PNgbh7Wjj5TZZEK3SsTnAWmyeZDRnjphU3JLh+At1/ToQuIRxK8dh8iu
IqXRlzSoQmSQPzBVrSU4DoG61E89duL58f0eHlXUyPf5eg06jRRHaSJdNYee
cEM38YwMRCdwCu5/XwFrKAT7XX0T0XWHittcm5lJ5m6zyXXHevy7HUBAiQrC
fN1IYL2827x6UxHYvKMYt9ZwNAI3wJ4jxrX0mrNARYmC+0Yw2Jx8P2LHSHNE
QiNKGKHF7IVYdnEVKRo4PdAYuWcRzWp7Lslg8OpFh36axF5cAWwPVfNW9K7g
Zrxm1eM+HTvNSGcGiT98i3gh++atEewXLbX/ZWhxdi3OebymFZtOG1Ab2ziX
S104ekf+JcKyjZ7A4Ai+gTqwlAxDqu2Xtuum/qlO6Jin5svnR9r6bQPhF88s
HXWSwYGe41u0ZOECrVnSLrj29Tv1berTerFpLdgbpeVa6c07OSHnPCMdQyt5
F9QbRM3BDpOnl/yl6iVbSJN9ZyYCuO2MRrB7g7bzY0SACX+9upvngBayk7dk
5gvuWAqhaM2v+JR6zHKAtgVX25Gl0ZhivZoa/fX48cSWtoop3nI37MtgyOVr
P40lpi5stG8psbgh1A78v8SXSNoqKl00CREVtA0pi+lkLp4u04o7NWsZpbaK
UL8JDJahaxO7u/HpgnBKRv3xYJhdd25f2AxoQRHWYHMzfH8cPOh/pMHLToXU
A5rI65EYadhvtg6lm2KIrlin3KDYOZgHe6cXq4AYcZCdKOpb3btpwNip9kjX
v8Q9p37FdV1LXaKgsHB4Ho4NILVfkFYiG/z3qR03zuYNv1wTq8zeFrsQ60pu
OkiBxW7unTmBXjlRr+UvjSC73ctmxC/vJCbJ02hgBvWz6UE2t6ROdyney0d4
4hQdd5HuRIZZdpwycoodeKS96W8pIs1wZFJlJjVwHcY+fQ30s7W91xATJ3MN
WxSxKsaIsItZOxCGU60luXnV12RiX2m0EzTWLUHG+4pcYjTc2gazpGqe8gl5
NOk0I8A5U2JVEhz0DRLYa+MM5wXiWzUN130qZaDEmEqnKqR7zfO0kE2u5FWz
IZRspJabX1DLgd56HBsFLBWRWFrHu5sYhe9pFWSbckZg86G9j65QgOS1C36u
cH3VJYkmliE1m15433agyvCLIDp6mi0yGtfUfCWfi62f8JdYKxnPqIS5AI08
81LFQekqArHOl9nqVCpbZ/eSQVLCc/KuhYB8KT8CZUeN1mMjVu6XMQseMZWp
cDiXV2ypqt1jkIhI6MR7CAP0PtpX86EgW6Lv7FywKrZlyHoX8UXROR95R93/
bTvL9Avz90uw/Uwf9oTcBSyucjV1u3u0grUeRct7q8s/zp4kIzQuqszfkTL7
O9eejJHyodPUaMNcDmjNlEZDDscfRaAjb9afhCDelLBZFBPrdbtH3FyLP+Zq
zGPD5pehblkgUvjO9YZqEUNa49LsI0RLW+D3gSbAgFFIbMuhM9h80udSXZsw
rduQSZFBNlK2QB3roH2ZNx+CgkISjqun7NMs8tC1Q6fSzmvXV6NwYprS1ox/
TEjjk+zlzLp4k92D9iPywyBwXVmwyzEKDQgr8YWXZH0Svd1RiAb1FiI188/z
CjYTcXvZbDXbc7INI7IzDc7g6P32Fzh9lFpSzta1ocUk2bkxF5CbQ6NTwsyC
4NRzeHxAhPci3hfnPgWhqRR05hy8AErDelVHVw2amjDtcuB2UVOge+/5BfgB
LtK98MYR9jXKGdXAvBWNjX4ZpvVZPensutLj2ZEz18I0kZgMIViMFqgvwz0h
Wlb/VL/iW3HzC5JGA0n1hANwTNBoTJQKwJedsc0De21VwjpmhlZCCGak/QZv
UHG2bHlFyxHl0pBh/X49miZh829avxROVC1loy26Hq77lw2IOzvEEgiRPTE2
UxOBrdCUy+mIrOvOP4nU8EAQzH5tAEqnJGQjZBZRwmZ2Zbw6ihSEskYe88qC
gkOQpaZPtGTXn+0IoQPLomRbWwMsk6vf45vMujo8OMY1mHLUbqwYZCIcJsVz
pAMtQExouyizY1RusSp3X/66kVHBlKZ63pbb8eIXflItpjKJ+MePRtY9HQtg
l2lAQrPjjc9CnTJBsPKAB9XlBoR3W0e3oCbZfDZiUr5bj4gFktbtWHqxg3bJ
jE+QTM6QjMGhhjH+3ViqjU8E76Wvrptrs1858LfyYrUaHCUYUuHPgVw0VnED
tUrrgy3c8seEcUWf/PRM1bKpWhblKcaEICe05jFWy/uICgGNBeuqSfIT86uL
iWC9wwuQxYM+B2sc8kTfl/sY/zsCuFzYXdcJG9pl/eF1cBhET2J2JmhNa1xO
ASgwKL6gGM5c2SQSIg0lDzZJ+EBlLyhKmeIBTj3DUflXRE+wRQydUHoJTyh2
YANw1wJhhX8CmZNG2eWgDlEAHgRc8aVWtYQVL5rBED9UVT9CGWY8kRxTs1R2
j/468BiyKqSz5TtAN3Y467/CGCGwP97aS6Sh1UWUwXd8vz4YJANxUI0hK431
6sWnqCL/XnKMtF4CKSVhequh/8NA9817M60RWg2Ivo9CytktPKyHYk5MMeeG
Qog6WtlKQ38LszTwzQsPBeUaws6WUZyy2SFyWHEEEs+5ngQZOnmhPjohazWV
1mmVtUJ0M8qnGu/Pq8I2yXF6t5VFeDQWBo2e+5hklc/DdE5FsuvgWj6bxxeR
mMyGWBWf+3SRlBACO61Q7y3El3vSKXvkew+5hSyCI+ViIkzu9C9RS/Vm06Rz
pS4rNmzfNCeo5EeiosDHlGTb4gWiMyUtaE1gqFQ68S8SAtnuLmq/Ttmq/bA3
LpHf3a7GxcG/pMEdQ2jE9h1LEBXYuRvg4EzHjBcnlpYF8CrbKi9AD6Nrv/DR
rd2wigflDZpsLireQ07MfKg/zkLFby0bJkDtcAxPtxtVAoS0f1W1HkLfIgbm
JA+g54qrNQaIbnqCRk/YLM8IAzuNfqfJIv53P14fFBKf7mS5Gl1kH4vbXqcS
9MgwSoQxgHBMSTfZ/RNwcobpaMsfSPDJwgG9Aj0wZT3IElLph94j/1nmrD4D
iqPhzEVhndE82i05Fzf3qTLQxTlkpKfLz2PrYDlLrzGlZOW2wpYaQW5KfKXD
A2/2AeSNkLrbJM0VmgQ31dqdBlg4s77qfk1ObyGK/gQMIjJnB7TNWktR+HP7
R0V4L17HG7NJap/mYkzufQ79HrdDhdWwWZKAXgQdj77rAY1yDMgSi5xcDVdn
wgtYwAsLjzN/XCSeujCFKSEIAwStVpxCADxGpK4p13RViVh54MwSQKdk7Sfh
LElTCevo0XnORnTkTbLJ2Aoa9XprWS9DJyd+i7ZEhaXPdeRIyPJn8KRSXot3
ncTjTbxlPa7Y678Akt6PfF9rFrIDUB92MZHze3mSUiY+LYbHJ+O96Lpl/xUX
czAOoYsrCCYpzCkGWelDKje2Iy4xGdbhk8qfWR7rLQ+SOM+Nwm/qle8YTcL0
07dezqq6jItYhtpjgfucb5Ec2JgIN3CPJvrPzUkvIIY26NrnzONzGqzmJqHN
SWNHAO6XC1CcufxyKDqwkAvYdfwRd6fysLEtpCrclLeWxQ7hRMfdUdnPX4XK
4LXbfJKNTGy7hiQxLIM0F+sPF7uNmPwxZWKIi7zg7MsF12ixOGqd6Za+R09P
oYXcsYdn6n8E4e79vKXP6mQAu54ni2JQMYfOyApwYXSnOd+mKZhdtRaD+xb4
UKFbm2ssJq1oAYBoHl1R6ceW2opQ8VwyQCtbFvtegLUb+tvdLrpyn6k3FMqn
AJqrBtovqAGb1NIJ/P4lQ6vaCgqngtOT6HrnA8OqkCuU2CtMey1M0MXJNEZH
pGdc3oj9kmCtNnOYFGK2WfJ80OfB29fDyoPoonPXZEGlw0Yru7XwLa1JdUTw
c27R+StrYeFmFPMjz4/Kmrs6Y/7PxhicNwOnJKTUjdhbSLUPoO0N1GdaAHFg
PtXD9pk7a2h1F6pT1YEvN/ZYJOFUg0OBrsw6v0yxHHjV8Cq0xnPFHPpJYZEi
4JiXBwXQlHXtd5Cb/ZyIY7mBMkzQSMFY

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EpZq19609/fy1e7MVlZfOAYX6aD9IBLSRJcQR49zPM8Z2omTVP5jsamjTnKBEY9zkbANPqa7wX8Ost15/mkY/0kVTuUbJnvDWVgy3QDDc+QWepOkWOI1oL3y+XIkTcYDd9KbQQorn6UqJu8JwHdSRewnyeFryRNDicpkhYPO5r+gaizacR3+hUHLYrJ8oZzSsEC5X9rSt6r9rNp2tTRqSMBLJNXfeJLneKQoWUG7PYDgIageER6rC5YOAisOAY8RIZ0YKhoTCEcTCSZjWvjOPpuhu2cvyodAiYEUazFGOqUvozQfQZBMOHT63dEjVFsSbIqUfP4QRyX7uB7ovWqDqEPQPorOACjoUPvTNP08tEg8exOdF5/xl4Mcapcdpsa6/UGXTK9Jqd5yC6KdXcF9ZaXD090fChKlY6vhhvVRgX6jauQut0RsxxK2XJs3989ToVHbMStnIHQqaLjOThXaTMz80AsY8lzpRLCXmP+yOTAogZe9MpFvrma0nFmx81dZWrTrAAb+3Q33xf+Jvy7GTdYMw/qnwBJN8viRCPWDXcDVw2STfNODOfZDdUgM0FUtxa95huM1AKfQQAQT2dXuPjRPxvkvckqYWKdim8uk6iYxBFLgpCqUGB+t0Y9AP4sZml8Ec634tMFiAOEaLlIzovc7AWOZ7z7IupQWDqtZh+vJ/MyY8Oor0Bv9b5qdLMHukRqbc9JbSDN1J13Cs6SRvXC5aPYyH6FqSypO4USglXKMJtvV/F8lRPxl/2iDF6tau1/KQJt6rilswvCP7nH0gHf"
`endif