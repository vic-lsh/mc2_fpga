// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pYkeR+cDBAicTOI+TYYhnfmiJjhobNRXyRfHW+mnwp+UuvQI4vtKKx0i9tSK
PtsO/zaU8783TguZb/Poh62j9yk4iBqD+eQzRxBpabWCdAnRXtibvq5XXYnd
aLtIuZI9S7aqhiffj1OME3ehWb2Fw7EktKej4B4zltzoq7c4je49dxCIFRm6
eRjDzmbVaXyO5gHu54IC1QwPWqv9bgyTddCarjja8uavlMcDgp09WD6U9/gl
2S511Fsg1yli2Y2Oxgs/L52HQq44Su013bm+jjzugVgtbfq1m1GHTsEO8tQY
PP+CDLWo4Wg+54PbtWzUHxLwtIdRViJSKcVnamI/AQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I+2ZVln039VSOO1wKxveqLThWbm0Dgnfxv8X21tX17c+x+PP4PSokiogkkMH
wZSpo1FFzlG1KilAaHqO7QFcCFMSXd7LTX1BWLjyQQfDXdGg/SEDz8ck5BTv
YL2cW12KkcJBLG0UvMinl95pCMCTLZ+96BXjAM+abdixrH7dnydn30Dw0pkG
VLIAnp5jz11l0G7d744itrOs1jRnLYCvETa+d/sksmKYeEPUCu04wkWXjUjC
aW6JfzwgJC654SqwFDjDiW3FNR5/cEiOQEzSy5AZ3glOTdK/uY3MDZor+Mj5
Bz8SAMnmzhu4ydMvFWaiYI1IMbrGsZ4Ud9uBUb3hqg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iXDQBsNwhR7JurU4tunzvSKfDN/oof53aMULTV2OgCzKyMNZFmp2a44QsyLt
M7HGGeEwnUwLHBM8z4gEj8PAzb60xwRn0qUL7enRn2fsS1esVWzSTagwELby
WzOqV6pTdCGjcUzfrdJPVUJH+8dMsNQEsf3FFeoajqa+uRouj44S+bPWrFIV
t/KAu3WbFmP6LQegZZ7KCL23E8X6faKm0a+SDNccX9TWwDRHiZd3dOuedhcO
L3KTsr2UlkUQXd3uLjD3ORA2hZXrjpXEDZ3n5vVydIdDfN/2AcLqnUARti3a
P1isRHqBf3e1Xg6bPAuRWI5YH7/AIOS5kjLQmEqcxg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Awu5Z2QGsC+bI0vgHWirUoVvA8Lri2TM7o5SK9jy6dAVzorEjJxO0ms2ItV9
QVtt8Pmt52LIuq59JnTPP9eVsJNQaJZs9WaNL9z2pptH5GYkxtmfMq6Zkw8I
EE3izpbuJUudfyREt6Thz52ej0zAzGMp2W11MsFj+wHlEEVa8eDA+cckFLxf
F7mV+q8FCfIMwh4gcvAWpSqpOeGbwmFY6ZkE++6D9A74ECKoV6H0r0EVjq/J
3kZS2552Z3cxf/wPA9AR+Xqkn+Uec7xwwpPXdpYLnAqumEvfDPIhm+MMBu47
c/JDhf/60NBMIBJloHw4HctHqkkYpTGus9p+UvFF1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GE85fcqC13L9vpTeyVn9GNHztIU1yYEx03qv03PJXNISpJQ3IYGcd7KRVwUp
BG5Xw7/Y79QbWQQhEM/whfEjyNZVv3eid21xJVxGvQW6NUFjQjDCOIezfZfy
N9gOsndvdP0pfhlqSbkCyNyP2XxhrtS+2GbDZKToRSDS+bAlwWY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VwMLunvsHFnLb0mqctvFIadL6fPyakQtIcA8auPS2jje+y5Sa8OfWq/FVdJo
GEtJz50xEFw3Fga64s+EriELn5FTdIUNueR1YRwnPzfWxX1kB0LsAA0fKpHm
x3IGyAgS3Y7dOa5YP2jtKWlIwc1h8tYmADpvLgc1kBnqElyZ1Uijh5FDHVsn
Y1kOskzbdF+iJfGEB76D9kqF6aW6wHuEv3zjCB+ZSKj7mJ/D5g4rvbSk1cOA
p6l7vVUmx5dPTghtTKrmxH3CvmlLioVbPt22wBVpDMmZCLf6CRcp7ulmO5sh
xIytzvZzuDGe4PqpR3ius5CMMCftyzC5SV9bYmEbSONjGoOj03MPJORRLARg
h8ntXXtNW2JdK5UvcZ0r0eUUbn4cptx2XA8gGF1/BhUpqxibrOsnHq6serFF
t3+cf/Eg5BF90vPgmY2K3KJPH+PXzIjjCvSCx3UU4LJLBH2uYDc3Lr3V5ty6
4pl317fXhOxawFrY09uwfZau8EPOXSCq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Pq+Gp8pXKpl99SdDMoCLLcQwa35SLVhu2txCm7PISeJzPULw2tFDQBwm3Rn/
ZTRBDdjNYUYITDRnk8vHAJtTT+aL004kZ9T8lm4FU1qAhjddFnX7MG8dla91
9B+/RS6rfc7dbv7uZie3hspWscUUY3B8Kc1hn1FtMUk3v3RW5ck=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SSEZHPoZDC2tmjmywFjwhEdf3rzHrj/PcLD7FAzk1l9O/GkLeaMPGn7GuCQs
3Ys1LWvkjRZokz5YTbUm1w87J5jARQm3okxg/80YASw69K/hY5f88UMdAg9Z
XyXDb4xH6PWYCew5/OmJNP+EQDXBLNHTSvMkdc5nn1TEQdzmgxA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 72288)
`pragma protect data_block
gh0raStEMn9itsTz5zdLcwGdOzvy4Gtz9iy+uiB0FFQV+Z3C9jHBlUQhS9kD
G48oETsxG5ZYaZ5YMT1fWqRKC3SmiJfPuxBZircFo8jvw8ZZ3yPg3Hvdxm6y
3UaPGv0kIA9SAJQDB5StCTsm/rTHeUAtbYWtPU/8NRov/vy07zzr7eYxb+ZD
e5BMvwV9fktiQZFt2W/URWkXY9WKBFY13gflkE/sNGMlVqUdLDKcCNoB7bug
F20UQp2CJ/0MlLrCygsB6BrQZmvkrhtO+keFsXYMqFw/aloORXC6ABpAKadg
sCy/wDWbEnc0JRXOZ3TU71MUjPO4QGzQ+xA5H5fNcXBypXLYQyvFsJZgCwwt
V/Sfl49+wJOeTGjfdEZxBw3XrV3+AAbrA3lszL/nwc0G0OGpi0/sqmleaL4K
fcfAwfMr2pBLN39HLLjU7sWrOBDe/Gm/ZOkYIcQCie4aB93bTGxYLd0K/0IX
4j5ePEMvwZABpTJog8JCH0jQwOjehfaGhBX9VOj5/1xo0wVi7+ANkB+OuplL
WLnujHcENueaxpkQkLf0d1l0CsOW9N9/7i8MxCLd9mhYuD8KJT2dlSsNvVn4
gGjk0r6ukqvCZ7p0XHhuMnWVdqcCOVb8db2yKAb4Z8vIdfSojaoiL9CsSI09
dE9N/bjlvP3GDp4CAja6s4BFeoeNpmu9WFfFIMWrFzOSRKiHf2dHjhvKEmLr
6udSk0N/cugIZrkPgxGCB7+KZI0qXDb5olsDhHQCWOU6YzFdFHyvKguD5Gxb
fs7oIyUvLb0u1jnf2fpRg6IOKcOlxTA9YsloNlv8bHJHLlagW1cQC/qc59Iw
MMzRNXuayJbLIt8pTHH1E4BOo336w9QtPU53KlNMGbN2fVe1G1dggcnkBVtL
rC2JRQ3wrzG/AZ43kmFsnTQt1/bWtK/vfrgb/lpGMEHMqF3uL08DwtbTk40l
tjIPdrWyn6OZP/oTjRQtyOVdBPe8ickHiJ+4G33I7XydOipXXSOCGLo4OVl6
Pw6tSvYKsDXaZBduTem11VXxln/17RSyCs9DMmA6lflyiB5NoHWrWFZhcY1D
d06M/e4rboMjHSY7gXJHj3Vj2GGW+tB8cH/1k4vJDz6/jEPagwEZxEgX4km7
H6qrqsH4W3WgSWDi1ReKhIrnhCiklklXRPHkO3slU6oXZ3CTVPBMjRmGhMJO
ouQDyCV3LlQzyJgxTWH32jjQlyb7/SfK7PAF+LARjm70KWBIPnbRw4eakzXS
tx8wcHPHuHR3Yxupb23EMRRltwFQQBjj4FUDbEHi6yjDIMsV1x0bz7OXdAtB
B7y11yVbE76m1KPgraulhsOr0FjTHC95LoYQr/fCkPXQPHyeJfOH0DGKgErG
bMfIANSMYzyPkmESQBAIHsKAsP+s2M3C452iO73A7bIbhYaLLPB24wuStlAC
CF8PakfkVkuxRhpCAWPo9F3ug1knGTIG/Ie/uAXp0UatsCath7kFteOriW86
7WW9E05OVPeUQ1O16k/vAgPA3TGFE5HLpvw8ytHk3+i5Ka5GFioCwMrKvtXN
uu0CvLVXXaI0oEYSIeZDuVOO0cp/bDJQTIaLSYtnaeAooFxYASo/I2WeDH5D
Lp/9VsYWiVSzPtvJjgnkknE40f7Ub4SLGhOQ+rgyNscv3xINskIkwMCCw71I
Qu65bMUy2lJ94gW59EfESKW1MhTRbsw2/9UF0lOvWcVjFMXg11aAqYFLwIy+
wbFU6EPWazFsWTKhkfaXk311nfEd5qnN5oT6JbccWTH/paQ28TvOsVJEgb6/
NypV/b1plzM9AnTR/IVefP29KescPxRQKetn5mYNdG9acy0xHZAIDOtllHZg
FCQ1tcjqHoHhQEt+A38PDJSTmiSrknKG2QNn4b/C66di8lJIkvpgeS4htxhA
LdgxS/toqsD4zDJ0jhNoSHq1uHgHGrr3k7O5aCkDlhFwqkMiHxvW59XFcErt
lkDdEB7ldXfPJrRRzypE3Q6OZab/6sy78UzuMd+WCukWhg163drDSJM6T8Ny
vw8Z1AGubwMgQvm17vitOVTWYvfYJC+pQ8lULhTRnzQw36W+kR6BjtshRCNn
ywGf9S3jnzO8SO8Gkh2lXS1hcpkT9+75JbEU1Bt2Vt/Ptl6eHKhaa5i5XcAV
YdLvCTVs75YL+vZ0G6UPKKbamhUnXczoCrU1Vbr/sC3eiwCUxS+PJSMvbx8B
Itmla6V1u84MwnEX9nixMg2sKtilyUcLRORV1BwtwCJWm/Sz9nLyCuPG3dZ3
AlF+e3HvuxRlB9uEjp0A/gph9Bu5//qPdkIIFarkbmSAIxcpBUr7VwSFctEm
m4tJbblEoFF/HJU5Nf5dAJeqRqnPRjwlya2i371nj3YzdYWdufYp6oshn9+q
azbUW1DFMkTYfTU+9VG44ZaxScAAcqD2YjixlXnapRJ9GjAz0fRtgj5FeTjA
VEwj0NAilWON/sY19l2QAIiIsIGLNg81q/neq+V7I3WglOEfoG/Tk+JOB9nf
xMjLmqko5ZgR3gBVrCOYZ++85xxLxYm4xA0RWgJo2LFDmIb1JuIFjl98Hfn+
3YFnka2Yo+fEc/Q2US/fHdurvPPKhslxTIyo7EME5rtw334taqjaf15CdJ9s
bX3Mw78mDhe0xkq5fG8EKPu/EPZow6MDQOLhHmqxC2BnFDV32eUElrJvKxv4
qiWsHTg3XOrLazi/ga98kNYJunPWd80WDuV30eU6e7ZGNxZQX0BXnveVFHbH
wHtY8NE1SAQUA8RPhJzM8AxEZsrlF3oZUu+27NXOb21e0v38Um9UwVxmyUzY
cp4gQ2N8nJ13IogzsyNg6vKiU5VA8Iasw5KJPzHL4Zrv/UnnfVw/gQDxA/BP
q9bVnjfeCPhzWoXuy9R7wS6+NQm9a4D92j7f3Y8NVU95cvMbtGI8tqH0cDvi
g2zniSCemmc+wOIpC2k6GdA3+92fiI7tKHivZ3r2AclpTW0mMz4ljq6Jd7p6
anzqO9kYYoOyw/OfG4GK/p+NJ9neVACj3LmQlxIoYlQcA8HeMGSoGXVJ5nJt
XHvjOt19jHElZkftx2GGyxeGVtMHtrWyStV9v+GEHdpUeU6KAalpUv2z1ikj
vOGsllXC774ctiXkefJ0xzz56s6OdNlGU6ly5Mu/Xlm7hbFD2YXvkJzYuYXb
GA/HMRAXSvjEifha87wJqF0qfYk8woP8bPZhl4UrxJG7iZUO2xT7QFUVmvov
WwgeCrrTLPx9+us7S3q6BRYf0zJkGlqsqnWfXJyB1DoYVuXpNnxrCsQBzypz
3pyGold4tMl5jf0rbmkKLUFcbmUJP2i8jMtCT5Aper1zXshV5FoO48xJ6RTZ
A+za8SEGnbMllK6E9reR1SetfJ1LpmwQM6+mGrx+R/ab/tU3itgmBOqcJkPj
E8fcNmlmrsLHXRuM03BgT1M3glW6EdHh5tdiUR2DUhiFf8lhINqxQoc/LytQ
qiYoBBHkEdoHzjMBH/I/EqEKjm0RABJAepLsjcPJ/bomVw6NEH8UXYlPnY1K
DTMRDllqFpbFIi9qM9JEvPxAVgd/g283zJ4F74RoSSAk/VFgxgosWTv5Tfph
ecfqHepRfZ0bMamX01zSG9Iuv0yTIaVmn7b/7BCWEWsT5Ui9vDHXYDwpyj26
qyX7YnKXoSEPs7RqvCvEkxKROpIKQDkxHsEg8aHrC7M73zvHljlmd2PzRLNN
Q4ceRHI3DdRKGeON/LeJzfsgHq/99LxEpDWIw66SddTMw9iKBDIQK8dDdn1f
u45wuzvSCRnrx4Ic43AckqVJ4GkHW9VEu/mAGmEiroycX3om7HlpezbD1ij6
qh723s0gFLGAl/BVDc8Z8MeZ61+LT8G5Cjj3a23OTNfuT3LKkC9TQ1VdSw96
uwQTf2uVy1GrofYtHR95Wvqmc8yUKE8/F4IluOgZEPQIgZ3KYX4R864qz22X
Q7MDA6bjwY48SHK8bz1zBSxneXwZyM+WI4kAUiPo3oiKQ85acJWX96lG2YM8
AnxyGxR7w+Kw9NBF4R3iijmaoLdseAgy08h3dAuLfENUzn9+pUIcW+D33dGq
TU+dK3OEHWsqLY5W49mPmzktg0SubJcONK2ah8NnaAjGREcUpZqayHOjsxP3
j12kMzZ/535QuND4s1FLm3LwlVHxwaDsKabCAkZcTS87ayF7iQyUM7yWAp/X
qxFeyjeIubNUKjvnJCse9HJiAVuuF6s1t/G+8tNnpt35CHMhnlIlqB69Fb6Z
X9RUMs+QpeUgKT9fY4wsS1/jjOwZ/zyky9+TQWAYdSwpvyIk2gjcdDL9eCAt
e2tbupp7easEtAmemUdwnnVFuCvOqP4NRm+eCftLixr/d34Yi2XoFL/hOwlr
Qfsw68NkqeSmO7ecl87ZL+Lj5IBJlwBG8lDkBQ/Y/jK/L6XLakFHabgMjf8L
LSk/nKKAZUMji1oUS1xHtIvuClo2qotlo3XnI7qY3bUaPiPcqjP0hqlnNtJW
/G0O7s2lb+GXyDdY58D4gjoLIiDHLp32bKdCnPZNlf8gjUPBIZmjBZmP47XE
bbr35PUwt+nBY+hbKZzJs61NXo2hX05FXwR8ThqX+k381LX03aw3WJw3p0lP
PqQmpjZ6qAaytmDCCREf509A44nMsb3K8LBoNoCUqH+x5gPLBijrYSCqJ0mQ
dh2F1mFhV0TGH7iJ3/QmA4c7lY5zP/K+6uB3e4PXWNFAzrVFqdOUB/aRRkcU
TcsZq5OPU8hY5kFxw80FMdJj4K0mM3Wd7BvZZEOv1VpYQr8gCLW2b/EZl5/5
5FE9c1Djd+2ZZN06D5ubUd+62JTso8fO66Hr/KTKTiwGKKknECpIFufHMX7N
nWOw3hnoMacA9nGzCnhlTvzfTUktgLgYx0mOmFOZHcGUxXS7wycRlTJ6abXN
V2nyXcZouB5z1vGMTbLYMPKVzCfHa8QzkWj9pOFjXItvIILVJYiTYcG4B154
0T+EngH7KTqP58i+6gTSFaOb5spEwvnVdY7uJn44VbWNRBgBgLUxijS5415C
YuFOgbU8YtOZXMYCThmiqaxn6gVwOU72qZAp7S3O7r3xjam57dbahUeaIJlD
t2SwjHCXls2ikgPiq0hYOU0IQcPWVc/5bBb7U84L5fnv/Mi0zjEs5iPvIeV0
/KBUC/H0rx2RjJm6j4MvoN5JpufZp2adGhuWrj3HFyKC9rWyCXvJqthKI0G/
IpQB+w9C5MT34ACw9fiSosqPYdYMhzT1kP+KXpclxdbVRHuIQqplt0HMMR+c
6wdgHNM3kQz2VvOKTkhy5nST+5T9zf24iSzVwaV8iRmEV8/lxc4cpsVIeh8V
baDEqEdbXrBJSHLJLFfvsobHMMPkCsqv2+g9futOVijXhzpqolI49PLphzxR
pQFVFrcguS4B2FfYJcXHsIpedJ7xWO6NqU+LbtStjewERHLQHLKYRN8lHHVf
I6/N+5MU6VMzqiZWJn8oRzMllkRnvT3DLCgBYY2EOJYhiNq1ly14teukctts
zKXjLYtfh876ozieU+3BEc/qGANo6C84iIYJULUBVjPU1PlLCV4B2Td7RRno
hrYC3CKEnSfCosP70vtPU94TXgX24RLDfl/fC+eVJVuepxWPN6o0iMVjoGBO
IE2qv1FeMQEDq9g4L8lOAaBHWkurwvOAEhuEbLbd0DUH0SCxwEhZt29h+b5W
rl986BV1VpNvHmcEh6jK7egEiFWBhuZoMRISLQcAATsTubPPMBelX18ukhGv
9dHOs289H05YiW0DBpVEUi+3x1M8nQw+RkL5EJJOhfC88xszQBZCYUW4SD0q
rY+tlO5vvaWM5aEgemwm8K1xGPViIxlVw3GG5FZKW0XKDJee3Sv8xQ+taPxJ
sB0r0/evmy1eXqOh0OK9uv4c9bwqdvDfSCpWpKmEnNT233nZ8OHeD0myF5ci
PUiGxT18/O3CKNGntY86uBMGkUvAytHRlMP2aKTOQcyupq90hxDLzAnCbPtU
IbUc1xsOAIyEkqZtlEILXDpcI6emOLuO/uVfAAk2oBmsmCbK4FJXE8kWIVhI
350wk7EkgElGEEF2EWjXP9c1jNIesnue1EYwHW5kC+dbpunNV/TOJIoaTV59
YP1TgdBtu2mfoe3nyCvPMstl5enF5UDIJs+TjewQj8OxNdGKcC47xk1W7hPx
lIb7ak0BcRVhkxQ4GlmXDkCaYEaA7liVUzfxV9aw9HVQ/mu8veyi/72HntHJ
WEDOEciL4qfLaI+rGjmAp2iGx7V4vm5LgCXUrjz0s0Jrj0oPJfLeyxY9wSk7
WBh3PfydA4sghirUN66mzURnGsDBAsrW4pxMZubSMoSCz4PpaxgGHgLW96SR
7n2XIxGAz5SKXkGZHpnWPgS138X1SXmiXUvGze94Qq0tY5f8wMbwJJ7RSPaC
8jMsoyxzzzBJvd/mAeojTwv1Nm4ODgIiY5xp9oPYOPNnvm8jC98rTcPhRLft
HD2oFD+M0Ep8k4Cxzj6wQdhNs0ZzkRWMpvsu0LIBQ3cKGWmWZE49rkpHsJHd
xT/vBuordEkelS8uHJx7+WkM5HrXMcPIwyQBO2pBXbDb8U/PiVV/RmXDyJc4
xpzemvY3tjNu1p95IbcSllEpMAQg159n6WWzmsNDV1YkioOBR3pmnbBEP4FK
9ibMzuklbEVpkmeWDyGZm+uwMS8uZnwJ/9LFyJHZUV4pYmQot84VC+yluY4i
Deh6+bVVTHMrG5J7IYyMYt8pJnvj4kZAcBc265cxVHnyZQNy1a9UkRurapwq
p8l+MzWKhyc2HWFw+ziBgPJDdfwmyTC76pCTnhONKtLU8WA3ZHtM9ifawbRo
9ObHR1sFizyT7BgzpqRqLcUj8GE4EeOYStF26zRgXq5//n/du1BuO9qnOiKm
bRwLwUbwF58GP9FSBsk0dGXTUs6BtujmfIwd5fQ/XZmGVVOSJSHeYQ+HD/MR
2kKfUzUVADPbItwZJiZgRHPHMR7jzLj5aaKqvnbaPB3TO/nsta+1VGZ8Hefc
xKxK7uvkabRUP9oteOdLqg0FOWiqfyOWK4uUhXUinBqybSqQybaUCbuYDvWM
Kcvf5aaAyuOB1q31Bhueiv5eAtAMmbNTL6vuX69s6muHwP5IBI37fKSHfWIz
uFfUjlU+IfrLx1qEfzZ/8/NSpmUUe2IS6W5w/SZ+kqYkWtm9cFrEqR/V5Z96
3qoga3Ph1MQwq0wdxrGX32qipY/0qvJE5BwXkZ0Krg6PnZ99+mtXJ+bjtOvL
twXQYMI34iK08zjpogPpjQFO9k3FkvZBOh8OyNQtt3nP00b3Q4YBq9TkT9vS
bxjfq/+j16a+7vIZuiH0h0TjrLkhMdDycn1aNG8ka7+GYerBFhDk5ihlRbmM
HO2oj8rb5dd5Vrd+HMLFcfYph7z2sST3HXWXcMTRiKhv46iTcq6SOKTTQaOA
LrlGCf5L6Jnv7jQ/60zwlF9bVLSzx/C8dHFY1G6pM48E7WdnbnfzRyRtn37f
qASOKD86oKnfVjN9vbUBwMfsUwZNpogrbP0vIG+0hvh+7BtDNYn5TkhOYTsg
MVF2iJOaYzQ31jxbnFD6dbfyjxOzQC/nfrH2ZSDvOxtofaHanma/pI2X0Nl0
k9XDnUUY1EpexW78l8DlaqLMMRTUUcrh/ROSC9WO8gfUKVRuPN0qPRCBfSIS
FYttW0CJzLT0ijzSZMCK1m9gWNDyYTjuBb7b+flQtIufcwYgS3g20HiDMKwW
4fAwbZqo6tRwtheo1+0INsrw0Bm6B/EPrf/HfZOiqVoKUhho3ABHc//2HARg
oWyeqgwrSuBK4/cK45HUR5wl5nCwGVsFxXE7QkInIXM0AlgrHhZz0Te7izZL
pl9fdz9zmU/mDswsP44NaiA6TYu3dW4wtc5Fqp6p5bFU3KqcNibqLGs5m8sb
YIDgXJ5BcFMYEe5opeZzuIJ04e0ZeLVLIlxe2MNvl9ap8m6nYoYhDvrjlMWf
hK7GPs+Q4TpowbpsaTR1kJdJ0IhyUb4KFTKg5rvWGcz7jYTI63DfY5ecWnKX
XRWyb9HV9hWH1F6TFyUZjRb7aW+ZEVOstCaZscJjaFI6H1lvoL8llCxYLk9P
ooV58SuCMyfLivaPOu9W8gjrfg/Wa/u/3D2aKNEeFFPIk2XKlgZ4MmfIeHtz
ua6nkZpbcDUrQey0oF1jglOVs8Tzvup6qq2UD4HjajvLHUxJLf6H0ODy3CQo
inrnboJSDFXYP2ow+ge7ZkFUH7gmj++UymB0hUpr066aybjbg5ygoWFrWDEY
gspWQ2mePtHokpSjpcH4d8DAroMVw6+mBIU/wNOMXoNa2qA/tSXMlelnEaHs
h1a1uBOxCEI0qP/tn+ooAm6Ej4SKdzFo9OeeN6NSKDhw4B7aQDeltBhsiRpD
8zp/C1Unp+xe6qEdj4QOovvgkImxii7/y53CB6WXHPlsuH9hLYE5CLcojVeS
Viw2kaUgTCmhwuJ0tJAPi/1++ZNrMFl8nKWNv945UUGP5zU3UT9GxTQULhLw
RMqqc4+eY2Xl2YgYIL2w65K/YQ8WSOxlcdZ4xqaSQZgZGwysfAADXm2eCf+H
aemY1D4mCvzzwlqaGxsLIDE/Iim84T7DclFKBzjq6A2Tq+R9pD1EkxS+S7gx
43lr93hF6iXzW5R4MBkAKf8DqbxBJXtxqw/lsJmv5zFWNpzXN18oOSFhRNUf
xe163xPgHX5iq6n5NGHLCncDw3RyepAtv1M72G237pNhQ6nWnd+VMnoe6+eS
hk1BcBuwImH0MzV5B8SUjibb0sD/RrUOgp8HPwMV4O+5B0KqdMgBZQagBs+3
rjzR52Amtgv+1vrDPLb7lJqTRQdUFOf3HmiqLVRMZxxVfRkaT2tMS+9ZAxbl
5ujd03i3/MlBtmx4hwqxSvqZpCB+HCySsYjwmWZxVJ7aUIPUIX5R4tOG5Dqy
xVTjfLweMB2apimnR6e/mfttodkbfA3Q1MSTGCyJ6DeW7JMX8aj3Z5D7gE6/
Dak6A/ZEtRcgcehiBwH3uUjZJU1oYZ+ZhIwJZAckw3MIYWBcMTk2oyeW7k6S
TMCDKdXyHFZI4p2u+M6o6scIGxuQxHxfS4QoJKa6rKj9niBOWrBvAfTQfqWP
dRk6FIUwQndwf0XcfqGduC/AaXqkfIfMkjMjt+Mjc1ikShHFSGH1H7R5MTa3
uQnbjZJdLdbJfIROAbnLTxOxZhzdjgz3NfbbFr49W8Enzj9KLPjJOkq5fdOy
/Z6SWGTn+GBTVWChM92UMwrIAbi2IpzhUbY78rM5JLv7LAN8+5uyGhvqrulk
ZnkT7V+lpVWfi+0PX+CZe4opEg6YcXvpoo/fBrjvGS+9VV+sQ2DNAbQg2Fjg
TxFuD2VA1WYR05XKXAc+VkF1t8bLseycL0KwpeI1f7RNm95hFwsKTpCQDmAy
AXy1l/W1O9z7nDGeKAagcpMaW9ObBPR+iNVQnlOuVOOo/hDUk2vw7pamH5QS
ESrMP/EVS2XSvdW6uFpsXaUldB1sc9EyIiXJyZYusQ2M4SOWZOTyX3xcIy1D
XTnuAx3ekAFraCwVStotU/+IDmwzFom9EHNmG8wfW5OtSEdsFOJKJlVfgTCX
fjMCyq4MMOh5vpYGqMFyH8W9wEgadXvTU6G55HJAKmxlOlTfusJahrMyA8QP
E48fuRaUzmLRz3KprXl3G80OU+VmcrTGIDIhxsPCiAatfSejsScXFly6yrdZ
vJsi7N/J/ul+NpbOBuLTRAPp24I0SfWbzUANkJqM4hITvzExEfHv2Iudli9Y
q+8n4htZXw0HrY9VvikOy1GJ9L+xb1wIgb88k7DSs7Z1+PX9SVmaLnNr2nDN
POXIPG+ipo07LsxhyXLgBjIkrXCJ20AZOMUAl9hoeTqrm4cI4NhGbFCjsQBd
IX13KiFIqg/vdJ8ZEWpPoROjBqZmqf/fH+eksQwpVO4PcWriQ70TqMNbTVqJ
s2PfRFUu1Wx2bmv95Da7EGpPajot2hJIkHj1ehwNLbEK1uC1YhPIE2jj3F4m
eVgzSSJiKzxNUEm/PT7MdaE7ZSAWDijWz+QRucynxz48ldj6iNItR1P33+dh
Npx10vZUCMWKOPg3nqc33dMTu82dJF2c59oYr+D/tuEkiPr35k3n5IrBirrV
6H2XZq6KeCgu4aqIoO3/VNbyrhOMoiRMfg6QcXv1XtuyOSnfVbMiCflQF1WF
ew+8MlCEIrfzxAchEBMFZN+icOBjNuZqWI7qtD03bR1jgStxe2G1MKeeWi31
bv5XuSDrGXbtxIZPxZlwxqBYIVQVsyzTwIcc7f/Ee4IrSvy8DSGOek7J75Uh
65pfM8TZ4RFbNjppE1a+2ByuExoHocJLEvXBbjWutwWJ/UN5WiOWtv6YwfCo
S3uptX4naWFnlfz2jmU1fBNhS5htQqOmG8tJkSzCvMBSxT3elc0h8+Ccmt47
6RJbd1LSuHko0GjIjI4D0SSnWZkQfbzI1gQxuaZYREFJhyC7HLNWMUDFRWhx
Xc0uHH3QbJJ5qE8EAmqn46XHgZLvVVRX6wrXNct/mF/cd3oAA7+6SaefDZKB
H5YOXijoy3HSAxcIlh5C/Z0HJ9pK14eykH9aTpmYpaZ9Q+38h4gg75WfPWTb
iOliFB0s6cy374EBoS2cqck8+YiVPIknmJvh8fbReFUCf87YfE5CNTnZ968q
MLpDmHB1Je2XIQwxHm1wN24nUSWqEEUO+Bgcf63dEsDkCGI5Tl3b24mMLB71
dKjWyDZSk6/2rWKHoabNU6Ys7W4WgeNvH51PQybrHG+0rZhnFWWYVx3Lzw/n
XFpYfhXzbRnaWYL1UzpJO+wAdq0vj9c9h/zqbPHJm5kvHzxY37UMIVdUbe5j
ZUNjD7SGzfOkI6EuV1Wq9lmXFvK5ayGnkpCdyqU7nD73DRErCUIOOrNRij4X
TiUaALMoYGL0WDkKpKWnMeZega4/aOYpdIMjsmi/Geo/J/UFuHa4LTVeLEy8
+NGVqdAKf6aqHQYTRra1n5RRzTH1s5s2eqFlKR2lfN+afipo1mOQvQ1MCmzM
pZcoPY51TH0WN7YLCVhKNJk0uyHG0+de5LzBV5kOfIB8FGQ3Z67+IpqhYRTO
sJcXKEGWX4ucPa8h4FcHvZ4AA1j8GJGgbdBfMcQea+rRMpXSlkgMVDAT9Hku
6tuckUHPKEfP7YUfUT4Zf4uTZB3wyt1Q6WoeFHHGbt24sRaM+79KaPgQqjwt
Wtrz7+lRrws6woQYlyvGy4Y9qxjm/n0yAkJnrVzdIPOx/L49AmgEeHASZwfj
VWfsmGmNlOe3PYHomc+CShrMDApk+j8imfk2bGsI7xUUoQpGKIRL90uGVp6f
DgpnkIa4xbFeu7CA4RynmMxBZOGmEgiM8N+w+JAt69TlChkzJoJxGTVqPwUV
qiyshZkZkVWgMXPnWjO3pxTgHOpRTYpuXuC6qpEN2VPuWeiRtgiU5Zb2ZDa5
8xd6K7SQgGymQ0zHIGmJVQV0ef62Kjs69BZxx+ACr48XmoNozot7MKfUvBeh
piiCEiL6miZ1bo7sGxuciBLpfHR9nn5UzA5T7yI67XU3gVdqbWZkSwvYtQel
X/jJJOYzLZLy0+/2j4V7rBrQZath6dsNBkQxExkvczOjMcheZGPx881xGBf/
dYoS3oJmDrRg4eHySBi5do3mk2kNIfVufiCssXWE3+DspQPEPEI7AirG4P8y
dOaEQaei8t8WXf0BKM4lw/Q1jt2jY0KNnZ7FxYI1dHE6Hm7yeQlVzsq+FGRZ
ytqBauhwv0XlMv2NCoNpYaBCeXFFuFvdS0aPnqpRLbSqSS2HUc9/l3MywdK5
VYiL1RM2A2nLc1ShsBJeE99sKpZFY/yz2cHF5hH8bc8RNOjDZpfd3W9WJh4I
tR9O0pJKDiAy2e63QmVxR4jZ4QlTBP41VnFnyO4ft2bkkKejbGjdjrE1r0yz
lgLuM8pfYc234fcxdN9e/pWO5xCSBMAAZoEBXoWT9RWypiKZGsub4kpgg46y
fI/RP2s2bCIZ0zQVcp9aQROYGkQJAAeL2bU3mvJBR+avfwD6177GFoGgJjYH
nqhVizj7Q2CcCqfZdcx1wuYa/2gMB1VwxNplGpj+SvTqW6vz7Inm19N1P4Q7
Bwyx1QxB2pagO4+sSKnvakvwZ2SF7vzjLjW5zgixylz85FA1S4HML7pxms17
0k+8jm7+ODR0jU53XdP3U3aue450qPUajLLicAa2hw/0zieC809v1o4Q7195
HAZ6ReRZwLX21Uni4KYr2HwuYEoVZqKjMnjI480yTxGlGS149lnCCX+jxAkW
n36XPAq4coXp/yNt7uURzOVa81FyUzdmXDWqK2Qg1bvQoceAvOKtWZmF7DoV
HfCJW9bi4INw6N80kFqVww5bXxqbAem7xLH62AcRjtoMcQZkJsYR7kOXTYk1
RfNEk43llwNLqGSlX36RBUrEnHcPZLoIfUozJL2IGVTEjgwJ0KYjz9kiI1dX
2L0gzfKbUVGyZWrvoOJL9ob09JwM73xrpN0m9rBJuwdIg6GtuEStwgucJmwI
+JUhVtClG4ARWi5ypHFM6xIJfChr0V1cJxI6USHpYsjLatwqudpNJIN16nso
AsQSSvmquZ/fx2335y+KKoOoyvGRlCYXv9TnEPzdAO9rtcVvka/j9C/lHJ15
JJH2bj1UhrXWz68ZD1Bs2vIPjxRJ/qd/6gYaxbOTA8Pm78E0MZEtZk7pBWuc
uI+vydQZ6sp951EHa+w3fP03T6aMUT7EkDmPbUYHnE2cnjPazepmGfFvJSfx
5Vrv/PELohlb6hKh/u8PueCiUHp7NGadBFq/H690ZRUDDj5cTU5WFnNIB/m9
g3ds7Z6smn2Oxn55w1RN8OqzvgHeUW1eLTa7to6cEFbyzVAvmZ/Nbdo0oFgP
to4/phiqusDTppmbWOYmofA7XbK6tVCTjY74fJzvZEbsnJCUMpHgxLrTor/X
1YIO/PuEsDcv8DfYAv4ZAgFAouW17R1Z+e47EL76iKel2ipJ0RGXCdJul8t7
g4A0+cWMt0IwfUA23+Yw5017xHXSSKFjl+eQ/OOde/Mujy1nwuts2b3kingc
xGbhRF1OPsZEmp+F2EPKXiExApHfbzdlGrweEsxkCcNyfO3tLdqaCaa9YFyO
alLmOY4Ym6uwYPKTJMCTBvg3Xr8fQ2xbmzAXJ5gCe0c5YUYfjXrbbMlNz/sr
ygkoN48igYruEOLS/YwBeIn+zKOC0niF6jX1TQ4/EP0fqB9uZBxp/rDzS/xC
1fW0SwgN7fRmuwjkCBY3iHfSWLzYwmv8rK3iE4UnZU6bPY52Uq+RTNoXlTHF
58/A8Y6Zdleg5uQzzv9Dk//aTMGuxjN4Kbukccj9wl+uXAlN0BUPlISgspGS
lJ4aQBv/bOSi2kRtiPqwSVmkInfbbYcIHhlWuOnVBhOID5BlIOn28NbnTDox
nJcOid1mNeDJoftp1BkOsbXM96i9gOMSlsd1VKDZ1s9db2peo5n2226gjFtu
6XWO9KU7FozXsWs7fldBuexBaBk6E49Bd1JNcz7RBONrLC6ZhrUt/9EV8zIy
rTliK82UF0W9Zvi4B10hOzBif042egDhN7mci5J9Gw3RTxZBiINtFPo++N3C
gCld0Mr5I5ihEbDi+PDvNE5ROF/A+zbv2sU2J4I3aAP+yUcAZBbfYLMZURZh
H2paVJuu4fDlnKyYXiKWkixW4aTuHUqFun0Lha3BQy9YimvYMRn5UlUpSk8L
KM1aI4ozOD/wqECBbC6gDMOol5rNa3asImYt2YiyZ49VMFk15bsEGZ0ubQGx
yP0KO0/R0S9Dm1Vhz4ABwFAojHSFTUral0wM2QqkfPj0HbhYfdueuPsqVQh7
3r1QP4my4TiApVKYVzZRbLKxqtG3dvARFRA8yS3dKViNcdJa8h3QLCFUbs/v
KFTTCFc27h4j8HyHuKT6jWxTaCXRyhEr+mtzw0vajrwz1zijTo437dam0Ay4
isoYZ49NnGWQ/Z8jqeBzbahE6P0iwll4Rhy7ToWj6ZUm6CIddUEcq/tQbGMe
NMe1F/yweTjvPqqw95sG+THhC5gmYPd8qOzhbgIa9bNaNibiMuuE8HMuepPJ
lL5y2iKYxMkVQhYYU8HkCNbexfj3Fa4O2m+Oj/787bYf2VHC//X9hueE1/+7
FQBQKRXHn3tlr4HJ7mFVrDU+kD9W83v8a0pUNOWYYEAbnLwRzfUH/AonG8Qk
v1HAzXW5CSXi6DESPedyzuJwH+IfUM2MuVVbQScMiw0YMvL/f9Ww9KKFQn6q
qOkrAP3ZAIOjBzoM21xhmFavDgzxzVhNDljXymHlhS47jxRKdo6t0Rer2dfz
Aux7Tb02THpSTWAvA0WA8lAU9ODbWaXalgLGkCTykaJl+AgkiN58G8Yu636y
9b9hx4Ug8XgCBiSUiZMARyW4hFjjaKSMxyb8qnfAz1FPdj5ULaBbGeGxtkFz
tK3CD4tDKoBsmtEhG35vJGRd8WFwjU0LnYTBzUkcfZIidQlLw+pt8Z/j3bpJ
BQOOLPuD4pfwuYkEVlPrcUk949yuVr0Fe+2m2pV4EkZpUp/WRTJvXhLynhZg
HinIO+E3ADvW1hpu3ausaG+tfjNsB9JJMYoQkQDS/GwgO6mnIQpBbJ0h+K37
VR/mzGUwA/jsGYmIt6wEkNRuKHC9O+Ic2QYv9ZxzgcpSMNVRCbGq9WXDI+3i
aYfArRyQRmr85Ih0QWIQMWb2YJ+ShF/gcVFiFc732sJwxhktLQO6rUACA4tE
zP53i6UDX/zcv01SJys/ewr/udM2eEAjkAsibMgXYntZCmmz5smTkzKEg455
LFw0iGuCCDJeKwMV40uwfsQNXB9usgtrZDlAMcFL8B7kmn69yXYTramR1GfZ
Wby2WQbsu0gR9njT0LwSyo07AF95S8Kgy4nb3C4vuoR/cv04CqBFKU/J0QF5
7iOVnf3rQlN+mD/SaepHOJ9LesHYOXHJm/gMoBLG+eufiUJ6pqDfO/lekZu2
HgmVAU3Ayonx+GO/nWaTwXVstN5S3NWiCvnlXQw8+7iHKzwI5Gn3CgUOVLSW
cZjNKeEUQt66rTBrq+nj5hP6v3+Z/s6+AN2EntC4LxFVd4z7JbpClJEl34Oz
h3MoB2fkVmM3OtB1Np4iu/SCP9AJc2fEq0dSEaUJZ87apkTVYqijWQiBxpUj
Ol6C9+/GaK9WTDqlveaLmljy1mDjAcgEaB23At/N8F/6TPym+luACQfxEB0Q
7exqmAECRpbXhxUHxn/F0VSanxQVu6k+WReIKMIEBKg5TqGkOXEc6SHT0E9z
RDjBUID0Fwg7fcXCcWyS6G+wKKC1dXWPJpv9BSRLirloFEJGFUNOjqR4I5A+
oGiiHYH8AjuriMX7G/k9XS5eDZvFON4sk5PapsIw4K6yBDPk3AOLdDF2zvAX
Ou6zc2ZARuC2kF2PAJNmMnwBUHgXAZCsW/8K3Vd8TjrgmM5VX1DVXV/QMGCy
xhoANGATz981v6fWCixo71SW5YZVwCUvq9ZiDn1B6x50spg7OrsMA520PcMU
OWeEcHmecAFCvGE/ksc8FeShStcVcu5h9YwxaKX/x5iCNP2iAzx4EP3WC12z
d3UrizlzuRB+49cOlqTELHTiHzAj21vYVxCftMKAHvcgO3lcY6X7jWMZ+ZX7
U9xelMTBsnK+n9hkpGlrIKqSmvBYLEaUEzw6Yj8e805KcXVmQ/N6NGb97Ayr
AKSsbtf5OQM9RkqlWzpSPqLBB8Sr+T0talo5+9r5Jc36m7xfAfGMT+YDGpaj
W6HHGLWXdfbgNXHsCBV3IUAFd8HorBm5hfEaLYejhpBGMWQL4XW2a+bHa/Ik
Wx5FUjFubtNpjDYuJxK7vuR1ybKQNcruc7M6iQar//m7PxE/jlJhqtJeaxc8
o03L850yFmeXmMT0cyeOqgvpIMJJvNzsJpcmiJuORTkEIpV6af8Xolau1Ws0
MW1lHMePv6v5uvwn4Rk634lP4mVRn2mEdenKDPL5xUX4c3Aur9ci5nIXrQbO
o12m0wIUNdCATk8lyeHEbvI8JgyaKr2jJ6zLmyZlrnqfYL5Ei0000z9aHu67
d1GQdv293WbM0gEQyAcMquMG/niRKR+7UsBygoxsJrX15mxy+UITk5+wWE1E
Hf2k4/sgTMxcEVSbh6csDrMW2NKcWeXhhKR0nFv8zxOHyjm/RXLP25SIrNcL
4Ss/EkiLuptz6qsXQQcnfltz38tewkWGUzvm6EYYIHFELBxhbu9Oy5WLYmv6
PECDh/eejXIUxbUB/ZQQcWDk9wfUoEVqhVHyvIm+geCCQJuxMaEq1FuJBgU6
THQal1Wq9Lm9pG+gG1Lxf3zgErRdD0Pbw6Zd0QZ9rZ7wPPadlXaxtt0hQodU
leXiAXIvBB/v93m4XNQvR/TQlb/tMKw+xI84RGHi/aAMojBSq9WOcpAsft9E
Gp5IxM28Yj7tahTS0mQIKQm3gpyGJwabTBLZKeaGHf5FhNAwGqW9pzUxO/RI
M0YKiloZK/PjmwwKA9xhfOG4bMjP2/ZcKsqES1Uy6OsSw3/pUrm3DqK0uhxg
evySYhT/YMOM1GMSRZH8U9HQEPZh2502nwCOc8DlQHQHQeVrVop1V+EH41us
LskUOGItXQQvjHE6m4CQb5XHPeT8LxnE3bKNLf9659TT81f8cFXYbTdaLfU/
Y5e72pYpqFy+Jh6Ni2UV6C6WxpdQmC/Ax3DzV+BiQjYjYtN0J9gD2jAaZThi
FFgOqNlsB6Zd1fMJyASXs6Zblo0ES5wak9i+udiU92KC/N1EnnmrTgRZZGZk
OC48cFPqAeuWOD3bTa6dewYYruV/6Az2QnYtVWkPm39xjnEf13y53ujIMVWi
oPLWeLpCLW5poK8Y0/RHFcp1PDYCtogzZRZjN9G9BYw0AUdwdnXh7Uk4atDE
WDHj91Gv4TQGjUEONGKMZP+FJP16nrrgMwf0Z3RTZR3xmoq9LGcL46Q+n7+k
FayldFlJ181zljsaA2xVisYa7F6xT5Hnh3Q/ISHlATwxtfOIOVcIMLDhYLzl
8VAcPwrk2ipH0txovUj6FPMY1AkTJR28GSz1TIrVdg8z2BEKX9+BCWYnxar4
XVCVesjVLLIuiXPB8QTzrzVB/6o+6ChxUrQP+hndLRZfAavpetVPWVpfztwW
nY/m+owPD4uliXIboNvxnXDsV3yGLDxPIV1tyhlJcdeiawK4Krg75XiYAU46
K1fp2s/y+GlnuGUI8sywuuaMAuSbUtW4eZGF6+ghqDQz70N1Pb1JQtTsLtXv
JScO+tFZT61w2Tc/XGogSJNxjz2uG3dgBSI4Fg1RuSNwPKGj7+Y89C23tA7Y
gVQCQl8KRzkOzaFnu504OTqLoY+bVfgB9Gdp2Y1d+E0QXsfLyx5ueo6shjVk
cwGc3mZ1OxFCr0rWL9r8c7G67uvr322Sp69rS/aVvfHmLn8kW+8BslEQxTqU
jkP1VzeMwbKBEAkyLUMz/YqlS6XKY6MTbPl00OuZYOFCyFNJi07aeqrrivMx
y2Q/MYGkYyPSfBrHdxpQf60qcaUQozAQ9xS1Q9FWunOxjHv1KhgpFA8BdX8b
3aagdZhu+TFs7u9/foy/egnm/gSYLi4cpOkiGLuId36tnNKiczR1DwSIIAUX
qkYMotLxQHu4txAQBOFGMLVGGbY0tun5HKhmwpnCH4PRZE6G2oGNTkAU5G0R
HxTHmCSAdCeRfDj/tzWfOuxFmIUcLszftZTOEnNo9rjBF5LuKDtFs9pD/Ktb
lC6MwjI5hYwioO9IlIkfKHo0cy5V+7b/Afd6k5j3KKh9jLGFvcuSBGzuqRDo
u9LM14pK3vQzm6jyDRlvN3aAiyXoXF5y3rhzSkcre4QvZfHHyaUD9CrQknmD
GfFxg2HAHGm7dYw4PlokeqFGRYGSZPR0xLTiWeGEuQUA5wg+n+9N2GMH+6f0
BsywXHXyVymZhbislzQ2K8PSg8qWNjfPjkQQgndIKZdCMqCE5Qk8vSlJObj9
TMb2ciNn/Y+Nurny6FywkWkVxKoGIAAl1QPpAluAdFkLVwdQxzgpjTTJPB8y
nLOO5uvr1iRZM6GnZDBuiMr7C5D+KZ31n1h5ouvUNbj2gVDMqn/v2rUoKLdt
ixn95Paq9jRUdmoskd662O0lJ9Pn7BNAfIkblTf4geR8QNgPiouGQWelK5/W
uAhf747Ba1bh7C1FiDINl2Da3I4w5QtWQDE818NLCkYCrfCJJTNRDGKQkWHu
+FVHVDG2FLwkyBXjM573Og+eZURQ4xo7RrwbwSeHPh2Xy0NOQg/XuWb7KXcZ
rLnTElBfGUhokGX2+Pvquav3Mnaw07ABiplx3S+g3qaad2jBzJqIIG8PGMuB
eqh+3QVnnJjyunO4+rgw81gtCOx3CUZWYuX99gdyQEXQjRh6voVpXiasAp+8
g061wvy/BkxSd4semhV5iw5W3cYKPnMpLgWgHiZenppP8+zxdCXwLpkX80bd
1XRSHvKitX+VMoyJfbc6Q7HPSfocyYoORlo3XMzgJ7KIinZnhf08eEG3vwOA
xjdW5FfQrIdg/UtEP3c1lnorsp/axfZbS5XRs/3hzMg3mnWRbpDdeBL/QI8z
UCuI/MYl5IMIr9gUNy6lb4ZnAdQkN/FdLLszdbk+zGG+NURSJpLrWkjrB/L8
yKZ0t2zHcM0vfbJC7ar8KOiXYqvPgLQrGxZemAJ55fW1iFthAC1xA4iYtyce
OXzHVLDRizp8EeWIBuNb/KHaLLQRXRvS6on/WBbdSZ9h7eIYQLaSmqGOudGT
LBpWco/jzuECupf5j4GrO3lCu+9C1XMeD87Qrm/DZi/YetnGGaYhYRgvOUal
dVuOqVSV0t+LnOF2KsBEIgMOmeVDAwhiZAboPiUHNrwvFNTSeMsaUQIbXogN
fe5n7EWeR+jVUsHuTUCBzgl6MPttk0f64e994fwkMqadP1ba5tgaMs+nfzfS
ogzS/DhkkNfDqZDwhRGstHxz1pynUcWU2vhAaGIW2OF623ClvgYDYbrHigSn
YY4OolNL7Qck6Rqw3Ob6g3oT/CY1fRH1iRp9lNuRHSpPUuyuRfhodU2Gw5g/
iAUN5es5EbJvCFFNRg79Y1zdU5PV/DavRNKmuWqfRZdc82gHqHonwQyWW0vq
ESTH85fEz8L1v8idBqqhzkxcFpB1vE5Mcr3CKLkH0k7mGen3RNDZ2Fjvj1cS
M3ZsTvT+MVRv+HYaQOLsJ2bMlYDwwALCCFY7u35v+rv1mkkN1jtjwYBlppYH
DRF7Wp75h88LnSH419/hp54Ko9VuRl4lMuIls0ZU4A8AbGKMpKHruE3dban1
LdN1hRRwxDXXkPvo7eliYaFLnVHb8x7wC0Hgn9QP4USujNOsnw/JkK1st4zL
19AX5YZyPADW3xwpqUjZa+vn+EYSLJvq6UusnLVkMCemVu6XLlhp3ITnKpCO
bNFv0+B4rpzoXysy3nwjcHtJrcExMNEBzQKgMRk876S/vD6CNWYRp2KW7jji
MVn53qYNKVGyfHQswnMKL/gkqyaFJ9fRSDo1xzI4gY6o29xF4hM3ag3b9iUs
IQxv5hPxYQ1r4e3qRS7igvjjCT/N1RuTrfDiqTUd8Nq1aA4KRIYY5KZy5b+M
9Nqy69ga/7PfIEtz0JYXdL1jsbkKqIFhJN5RlT9rOKYNPqRrsxGYHCSRIX9b
L72P+ApXJ4JNS5tJoK2Fo+RFh9VyUC+qED2OFkdydCFrhHuqefPEgIbsjpHE
SaTrO3lJIO2TVWxsAQOWxI3sNdauVri2Ewhr0veHkUktkVD8g4Ha7ZTi9Sho
17Js+M6W3EZec25C/0DV7vsHk7XCuqLMIC9yiTgqZdE/iZ1jc9W6JjeFqFFj
0le/VoMpSMQhOhFzvRN7aLmlqI5v9OfwMyMAwcugbdyI3we623BlUjCVNrxZ
cxNCn/TIfkL5/It7Ev7g8fuJjWcQfefz+85/KxHtrtx5INHC+KVfsTvp2zKA
O1Z37genobIv2UG9AF5Y7ywB5i0POJtaFz4nUwUD3MAoj1KUmf7tSCEbNKgH
KoOZFVFyz06mNrBGa67NTP3qizI1NzGEmcBnppu1UnUKWgOAhC76H3N59Kcr
bnMmRFz47rz5jv0J38ODWlmtc0aIPkOd8qEKoKBdJxT4P5/K3o4opso4mfpy
KqnbsnIqK93xXNUf7ZBdlIRz/W+DLwgEvmOq5QsrkkgLfAYlXT/cb0z15LfD
qvqeUUvdsLNS6zaQ8OyRyS6cStTuN1PJE5MnpA9oxNFWWGo2J17yrwqmHiVP
9BdGXF0s8b3VFFzaRb5ofC5+N5TNint01NJknahwbQTthXX/g1amjsZaBbPm
hYXMmgGCivwFzwdtaOC51D5e2507VfsrI/gYmSjHzRBNv49AHg0JTemF1BNq
ukop/le+9YlzVlxI/TYTOiaRrSwWFI2pBuCNs+VgNlOgXqX2sp3yslyIqrpE
TMq78sQnvyVvC8F3S3PHACxZPLvs0Pch9hGAwMfl1pWhWwx5UvyybVoMI7uC
b9ocKBVM+PY8MFnM842S2rh20Q0sUdN8qrxwu+04a2RrKzfoif9D3SeoPtke
SJg3N8EEn10C7lPtJ6rd1eprD9Lpm96r3Dq2/1DJei9t+I8FqLLJRHoCuXNn
F1l0ynLabUNcyUnjDnR4zuXRRcSLunr8ATUlxplG1/QjgBZpum1p6OENb+96
AC1P2btjLjaSHroB1C5tcG/ZKkRDlKkD+Lh9RM98T1aOGnMvsJZEdp9GBsu2
D3frn6Y/ejZn6aX3rSxMwUYRcaI8MyhFtjjHKEuOymAdXFvsvJl5hm9uxbeb
/spKIW53E39sV4iKbxos/amob1phTzppp3vb3e0PWFrcPPXPKuz75apAkwTc
3V+s03TnvzcHqBl5eozZti2y2av9gu5nnEyOK7u1ELyfUxMN71o5QJn2A7C8
J5rZBSG9+7M48f31CldsqdTwWu8ZyRzQrY6lC4J4AcG9jIWYGQ1JtS1j50d2
03uSqV78UeJa44dk1ml8INuuCtXFEzBNvX87VAXMCPebIs1w14OpS97FXMWH
QxdkWLnd+53V8VjoB/zhUeA2CXb4fdM/OeQ31gZzcYs23S3iqw1gNxS3tKLx
XXW/sfukqPyAwbBQ2rwK4mCezicHUqmB+URm6rdFkD3HJhUdeeNH9MYqNUpk
wBlOEmBYgZYOVioqlrJEpAA0pDBVsaf973TjxZUWeq86zHaR/CocCaALzE02
sZkDdAMTTzi8uRff9IqeSqRMvG1KB6wZei5IFMMuM9zob+xbGbbDj0eVVlhM
5xz4bHzOfozzbCUYzIAbKcjqgY0oWnZaJV8cfqO/5gB726Jfl4LEU1/kzagv
CWNj5SUU122KTiauOL5PAz/6S/rIDeGd2LxEi34c1yOvEWV2ErGxAnNEC56m
UZ+PCUjERtYmDobmZrAmHo/5BcbnXLSaLhSXFvSYXPP6qCYFicDgw4N5bnCW
OQJKc6L9tXnSrzpsjDfHrnJGBiFR4yYKUi9mL/aqu3fMhlTdOg2z5KQWBW/N
tFjdJsNjEQOEwbmYWmA2FEP8tvAfWa119wBra0n9vp4LrljXYWCztWD4O2G4
jr9RtBNbnUorF2gF6+qEcrS/O4qolezagvopi820XJozVY68YKi6KlxneUXt
hznVO9TJfdJuGYlq4I3YXtTTpOqKPJn71/QfBSO/mwDcV9iAL9AG4f1byTUn
Q5K5dc5aUpvH1I15sLNM1RHVuSCnYkKnzYypsg+4BNe+MEPUNxo+OOK6Nm2x
spahIeux8k5o6CWVxwknFLxSlUSoIxGPvzzfwRdXQp+kvhLD9P2SzCXvw93W
x1TBcwBjqSfaMwqg2N958xCtaLP4Yrqp596VgfOQzPz6lDDMx5xVdXpqxFst
+5ceVxApQnBaXYxHAyhALMjJ8tZlmRgv7ui8nerCc5e665izWEBrxq0PRsPK
IPmv7v0c/Xh86PFoRcnfOyGZEVUAYyDnqTMuVT7F9HMhC5LWOJ9YeYVpTEAX
p/IpsrUgjX7GgjIEnh4BXnHXU2OxV6C/h5Y9Ilr0nyA+lE07ZhyNUeQ/ztWc
HBUIzBU4QiJ/vaC/86xa2EAZH89RweAmpA5o+wNrWp3caRC5MIJKb1zUJtg/
5AdAGQeIF1CEYYpkP5mCmGVgw4YzuOBiKKkPrjnPykUmZfAd074S8SaKylGb
41+SwtIJAhp//qhgq11+C77fcvJ01yWQ8PB7OpzQ/dOIcFmhMGSxS637YJ9k
kg0LfPsNhL+NiQkKxhUuG9dz1qwmVkYQXFZt+Baaymh0EEUfRpgi+Sa6SboT
aFjlUT4ZdIPXKq3B1Hocb/+sCkkH1UMtnMWv8Jvx3g5KwWGWdH4dECHvWkFq
6fYSfbVaZI1o74dVqJVBH61xvbT+BKHRKERGvBly6TcU3bV/9mwEkb8Uq2Yy
rmY3UaezYiDJbf7Ir4xRsp5fbyHUivztHmTCj23Pvq8BCSr8ozgnNYIM9oIK
YPlaBCqQ6e3PjdESXHV+/eVBXjQibK0wiNOf0B9GOMAXTOS9GU7r0ewSUT0/
HiWgUa09wF2IKQS7k/cSC8PodvyIf1uL6fkbIKsLPLYIuiEDi8tCbtxmiMBN
NQo9VUf3QMBCpNnwy8y7Ly6c+GnjyHVtz0iHOpMshwX/DzkiRyQMvnOCpG6w
jhHDDxekf5Q5m4Jr8YXzmUMwP3IKU8aKGHXtz1frEeK5ku9B5PbXEXNoZG9h
TAWACe2dBZXipVb54f6z4C719qKU9sZh+M4smftci367HA41Vmo1EvZs0Zug
jkBSDlNNPr9dtjndayANNLOy59L9ioAIHmjn/htgY7Mb5uCjuC+POwA8Kion
YSi7JZwa7T2qPb4mJoLaMhaTxMi0xRHk67kRT439kRaa2HYiCMrKp6d+glpd
pQoVmhgAUGwUfBYsOlDzFVpEvYL6o7fa102cXej8kD5dgAAneD/EXsCNZt7V
/bR2RtXrzrFUXJFohQlMaSpUMzSiCjjtT1euBlxNhQBsATv/W6ed6N6RMvH/
mek8lFCkOELgxf+5U5Pjd9Ywc3ngArk0zlRvPwS8eeNUPyIk64Gw/4EPJ8Ag
4evxgaIxX/3xCVWKlxQnSXnpO0dAQInpKUtos/RnZi/acPEBqA1Y9kvJFWrV
HB4Zr86xRTmSvuTmZ96y40OcXNGmKggARkFOlLIwpHn7XIOcwMAwRyaZNi0z
aNk2gwhxT+m7WeEeLby0EHFNpCMCv2n2QVHp5SXtRnnp4hyr85SURFrYJ3Ot
ioRM2wQsE5kXAO19SliGBlwW6cxKWiYxQpWMGgmG7R9DjHgIl+Kh6CGPfkys
iMDtws60eqT7goINgcXc2zBz0TNYFZSPfh7l8vUS61emW23WT63h5HaXbamH
NOklfeHmT/+Gps6dESrG9uJ/TeFPjdh5+bgvR+S1d+q7ZlMb3ICyKSq3RueX
sfE9tdnQNPNBgMdNQDV/9mOmw2EQlCnBaJrG+OpP0D+oGunVkIyc2apVFM1u
sGM8xZFZKXIoc8IM1KPHF7BfcxBaSiy90W7r6N84QJcG2AnJ58iW7N+CV2kL
++w0hxgRrpMy7LQvv/NcL4VhSRmLOB/NTMOwUDQmUOeecwXQ+KUWqHj3zJ3d
U8eRiTfxMDWPXU3ZqXxRHQ2Fvj7Y/5dzE/MpKP/3GRCW5NwlIwq7GSUSQk2V
nJxn3MHJGa72pNwEs4ecG0S3p84IpkqyPXtIj+GThuAAQ7FD6y8PEhy4y8wc
LZKyOyeIXofKdRHEWP9hNajWE94thsBMLNXn2UdAlW12kleUcXeI1MHr0ZeS
q/n1HoZWEUbkrHsy1EeT7W443quCpr28Vk2dmHVPceU6STdCkuYDm6kkv9vU
nBxs637HxD2Qknmqxrd30jzcuePsXGYsYghLanh2ylJAEQHJhaiYTSQu+zDy
bNkBpQo237RdpNaxZQ393IS+GHGNhNuc3Ayzegqn2CHa2ll8i+laxL+sFpax
lOMgFKs4xgk4PK5JtE+P3Ow/5ECDST+OwqClJUvO2ed+o2jGoz7yDLEAMAJl
TuZHI5rv1zxYSkaxFRWthOXJWy1Jyqh/b9LINw1dTkcLl2UEqxYvR0Q61ZFv
vU/I5q5aWqRTqWOcoqdbuQ2fLaxk2Mr5juFthQNBicXEUGmZM3qhSyT0ls/x
cQcw3Ef/ZAliwfK5hgigmdeB6Gkh7m6yA+qHwLDI/rFAFJUIrFdwACH+DT1d
aHhZeeHSguLM+gpy4ntWMCAPuUyI1FIczDmf/DiuwtbKOzUtvccaOYpSw1hI
LEcMw+c+QioZvVrwXzSsTpZe/401Iec8ClAd35els4wNQEYYfbCSrfusVuS7
5AzeitzRYw11iUri7p0m43xO7AUgmJQ7bOBfL8dFf0RkBRLA8fS9jlq6UM+V
Q598PcxDZrxlFmUVq8NakBw4PJVsqEnlfrprceuAS8V8S/RFj8VEwKN5lMzP
RJLfC4wRxZjWmA9OK2XinE4eClwP02f2xeLoIZpDfQRzfmx4Sj0SEuOLWkiQ
/E/AruW6XFApICCe3Kc3LG9dz4IdvbSy9T0YzxCmqKJ9mKkEKRO9TEh04ukm
yIVixxIqImyCaQLKOfHAFjHRkrv4QNaN0HPt2XDKIo16QVHuNi9bnY0MRy2/
yZ8zAGHr4Gk0MdY10DnrAvAtxFmE6DqLewlhwAXlfkp6grOuX9U+EepsDVml
+eJ3BeoOL6o6BdpN9JAvftcz5SHCpP+fG+17U2fIce4Dsrja1LYNguC4AMGL
R7tgzedL2jNNC4jxWrqXZ3OpNMzkPz3vAbl1MqY5ve1Sqrz8hKrlHKxFfrzx
StT0tvg496Vxw7NbtppGhQ4q8UgRI8n+FCMmQxWOMtd9DY5KRHIDBjkLjyH6
Jx4aCf4c44YNwy4OnvWoop2XEtQK7XRO5pd/EWVwyozq9B7NaSUehhGptDRf
I6gZoru6T64KYem10OpfQKT0f6TpMnSytZXxrPBLKpoyd/rnlVrkP2QsOnKv
CtNXSSiIo/IIxklzWSdZq5Sjwp5YNGvQKzYWCgfczeKPP3raBdmPLSMwDXFE
LAdUQQOHPO4aThjtCd3dppDmWH2X0MlieAPKXoOUKnFpQ8/ViMGT03NBXedD
yWoKlxGWIHXS3gSSwCrT0g6DmINi2yQimPUrb5zVK4EO9rDrAfvTffEtf9TI
jBIcn07nMAyYR5dK+uVBlfu7go2nM7BZm6fhSDlrBFUIn3Azot/f7EYSeAWp
C1uBBIZHEjDkGp45erM6kkbsi8kfRD8O8f3Hc0br4CyUWRzPVHVOsbHsoUIc
UVFzPAOAuP8bR26AdHqDV2tbpZj+b/dnQwDXAyt2yZJ3z6CHZzijYud6ALD2
kSfgl4yIQvklTIP5+hgtOA9jIyX3GIUtt26v/YCsLSc1F2Qy6MXCgBQiSKlH
AEQJSAvGyztxinpu2+UMDrpfIin0ugYTT8scmLlPR47KGMbKnudvYYVyUEFh
LDcDxWsp3ASShmTdWt1GDsXPzaYLVUnCqFOMaCnkToZMdb/lTWkvkBAzZoo1
GLXWyrZ6W+Or5FmQrnMh6i7bR9c6R4dfG9sCp1MaOVf1OnauQBsp5aTtkExE
CWfEeHNEqLPMxmoaF7JR4VpxsKNQ3U8vADSRTnAAqhFw64MS1dqlIIpjQwTs
SVe3r45DvUOWgfmmkgO7HjJQLzQSmIh5TxP+jXfnKyg8ytLgfqzgW9Dp1vDD
DyKUYk59nh1m946Wch8XkuLmm3uPhiS8vwiCJp4dpcpoCAgoY68WroMAr0Jy
fJQfPJg8xlN/K9gF+UNz8iAut9XR5TA15CAnVjcW5PkPAYVENS8rHd1LWnF0
8qWCw+73BprB2dDOA9Y+LnvFTd7xKc2dbb/NLPFSqrdBQRP0kYXsaiBRaOdR
fnuAjZo4u1KD09amL7y9mhOca5PwEo3COpXVLk0be4PNC5N3NqTnM9fuke2a
N9S/JlRSm0/nsZJCtou0oPgk8uYjD6vLqe5WBD791YxVw7avuq/ZfdPht+v7
3dQHoFmSLEufnzG+1P9PmU5t/El8k9UwRJ1yNu+5cfq/DMEvZ9zMVM/MJMwU
hkx9eZ8fEaIjySgDMExGvq2dmmwV8Psbb4Psz4BsznhygJQ7tvfImk8EwsQD
FW6z+Hvpq+Ib8yfBmUvDr4jT8zm2NcVvvqvSryoK4w8fNDxcIvODVL5C7rwX
fs+w1p8APgPXZJ0yM+sfW/J7zvTyLQw77eWfPWTctn8aM71nlzSGhzQ4W7hL
N3p9CPSodogUkQKHjudcZmZwQ1lBSfzIZuiLOWGQRl/pPr+aPFMCJSWIbdgc
Rp5UH7iPubPu0jbDToIuLHN+jBcyY07pCFYni0Bj1hfpPEw4gt6MH6fLLVAF
uEKP9+HCChxnsDeahhXJuyOiiINFi74yvyGESm3T6UZGhd80Hlc+ougs35Di
NcFnIM386YKeDJfDwE3aQtKWYJk9BhuKwJ/S/TqpsRAsVlt6SUoae3TOYSKm
a6gPhyLvNH7T/IrVm2Auw8nN5y0MhOuvK0+n0siHef45Tr95YvVlDP5E1d64
oO0bxAk+bNs6JGvvDgiBBl5jNQs60/A+ljpHcRq+DaBqfCiIklDIbEC/s1Bi
6Y/sHIDTmBneUcRukjwPtAPKMMD9WrciZlPlzl4lK5AY3qvXM5ooFG2fQybU
MIRZzdFwJ7Rj5JOBtKwurO9lGFArfHfRvByU59pyRpv+xC4V8OgYGpoBKFna
DPahnCeCnIuN2JHaDEX985gubozUpb0jJu1nP2+uihx8NsVr1aM9hXydsQ0C
Oxkn6MqwIfHhvz3za86jCH9sQaw4Vppz4PbHt3uGkxyvpv7XETdYFpHRYPGY
+AYpSQgLwbQ+9SF645U2NhPvt5IPp6rAJNR8lOt9ydc1ZNEgtRvQoQJoS7yd
8EAB5v3w7q+5CT5voRKev0aOUVOYgV5lE63mOZ8gpean+02xwwRF+3o3rnlj
sgUASd5BH4yDjczwjsb29Cu9hsXYyPQ+yaoHXzwj1RB7KZ4PrizF08W9UsUQ
sE7tOPQnlFMcvbXILpKV4RTKaGvuC5viGL77c1F5/CBMdXfCNxPCu2i8Y/vx
heoEfJAvEf+UgbAVfyuGcQu0QwuOzE/h0IuZyRk/Zp43NkOb7IelJqB2Nhh9
UlGPJ4t8vNvfCrwmSg5fgmliZlw40i9A9wPNXUVOSL6jWTvqKVCxfGOuj5Rm
klcfiTEAMIlNH0tLyrOhzsv38L7FUDYQBnOwoEc3q+WysMyAMsripOAGMOiy
K+thCMOBXm0MSWBITdfJttpyi4aaGRtvpPeg3V8rnXqy2Rq7HXzp7T0rSqdF
TPdpm/7qGYEXGT3XazbhUyOY7luP+g8lmkAC50954WeGnGNFUztDAnh4va3D
dFMr1vtKMddk002RKOrTzD8J9psuRwtr/fPWit6ZhIHuVkTOkV/r4Ghk3W6V
TkH0rrVHjRVM6tZJ87U7C3VooUU3NOillKOsD+RIxUlP9L1JhYGdv1SGPyPS
/cuMGkC69j5ItOL0mr2x/NOW8n6cs3zBmsiiehh6TQVT852aFWvY7d29aufL
offORSURV0hbZEc2zx53sLJ2pIrCI+DAIZTVpV1mWELdm2YWvFKllaK99dqV
rC7A6thAovA1KLiU8VmMvTpfnfka1HDr2NssrjTfryh6eWrXQ28IFD/Mz1j9
OoogUxsWZYgkBfvHHefRS193H1LXTYeYcLFrTuI5uQAnmzxs8XuH1cd9cNTs
ATnRIT+EswGaU6g/qwm/iFe+HA1O37K2DgaxssLH2QT5vd965NXsRECRq3hz
VGhfU/msR5sz9fy6qYx0SRYFy+6AXZ73wc/VOOor5GCZ66iNSNNLQzLPDDAc
SVTF5ygYy/F7OBKzMYZOqDZPODI18aZah9a8xxDOREYoQA+8WafKtzkkxWHQ
Dq3F5ymBTO5RWldkTKeQov0ZSWt4HGA5KtGS2nUszVnFNqp4N9KHRev9MDW1
pbjmDThCtu3+VSETbfBvESz7WLJcMVrZ1OPaHIbURcMswQgRg8CnJAzj23BZ
KpGE2xUncVFxzz+to8qbKg++NbeZ50eXLeqNbPeHJNXGnoP249Pn2wQkxD8Q
6R71IKI9Z7yk2EKRx4wn8ShzRlEqcPLM4kfdpJnz2CY6ZkRWWK7Q/6Fy7Vq4
vuMPCOcRZ9ZWbc7YAdlEeUTV89lNG9Xkoupoh8NJloO30PfFnlRyNnsagYjv
cCK21sAohHJ8w5XnpVKpDMPitBAL0k1Tv+LUpleJmp3ol1uoy9IX535zD/ZS
yxgE0avJPudeHMBkeMDxSewS03UcJzlIqArvFhF5QujDPdtjM16wD7Mnpj9M
0Q1MgH0f5PFVJm27tClC5iwI+1Hv8HSz/Y958T3P1Lgq2ohC7L8OjOZl8LYi
RvSGx73fIFq0O7Uuj5bRPcAOqK7cmN/Bh3x7TQzdw9RvBAha5qdF7wyrsjWi
phERGMZD4jB+hC1svQn9yxm4iR7nCBlxuJVjBe3BDFaBDeQa0NogIj5S/yRe
IvRclVdqsDvMYpjWYA/g88REIsXaIWJwrVXxFBtc/wQW/WOKED5ClMVJBDqr
fO8ZVmrx3wv+FYW+ffxvuITiFqb9ndWAHp4Atnma6TbeEY8TEY6cV7xLJgla
iGBVbnHp4wfPV6gFDKdklsN0yr6lijmzFAo3C8hYwtiG/OlxlqXvwd1f1vCJ
AmpElBao2SSlx1jK5uNKLu6aF/fo4qTJWWMHPRuQ3vzjSgWxpJttErwckHns
R00WC223bQQg9TzGUjr8MsGMI8QKxoOq99oOzgcqA2Z25lewYoWK27DfuI9d
WMq6wzrWg0HD1dHw5zujdJQrzvKzunAV3nUXfLgDNfjXOtItUbctApTio7gi
k0Nkm+mNHHtVO2u1N1u2hpY7LZsJW13golqWqPm4Z0EyGElN6A5nqIgcPcmB
Bx7qYcIAZAt35Br2ts0W9/d1peiDNg4O1egwlbdg9+ke0ymFM9Jjf3ogiR+9
oDDP5lVJ8oJUids2oMwGwk+UH+4LrJOGCvZkDD3skvSkL88PJfU9BU7sXCVt
VkEDzbU+g1BBKlLQumbhbhwHMVqG3xedrOyq+s6yNiAwK4Tf9Aq8GZMUqiwp
f9dRaow3atwq1Ex2Y5VTE3yUuHCDhZHS5Z9FkCRwmIQd3Gw/cvPOy6GkUlRl
FtEMDZ8tWJb9Ug8DZkn1AQ/pcsuAXqaIIDEL2WK9AKaHRl+FznX4rjkdkjIO
UPZdvcEyHJ7tOXqZtpJT4Kq4u5Nm5HoYOf8eZMGsUCxrUnLFwT9LZAVVhAXj
D44yYQnEZIyN0SQ42CaIJ/aXfh9h3Ghk5zEaRkSA1+RxpF9uqMUA07vQEHqb
xY+UzruIBAx3znMllmgUZU91vlI34Yhiz26yqB1KJDaVfjoplBdWSzhqYOlh
zQHPZHxpb8NIS8LPi4JbKlLEmw1EDEt1h4EPJLxJIuxC95oIv6b+vWIuyvj/
VLicin+Fgi8iyFDZbYEVm4oAIDpXJt6mZtHmlsNazK8cDZKsVwlyWiMOn2O/
ire1K2s15E0qmsTbEsro8/apz30e7uUd6hNnpqwpkgig3mLUIPEnP5hm6NZT
+Hn2aLIqhOHBtV3tQRSk/Lwfx+b8EXD9pRZXbFsYF9ItTE08ROaAAhz2nv40
gr8ZOquW444IUMpHP89JxM/vQ/OQL9xq4Co9vc+YoeclIoCJyIY4LDKJDnk8
mRrdBkFN8umBXpwtds2MkOBtrApAhLJRz9bC3+FVHtfD1QzcufuyfPYs7Mrv
fzeQ/GFSv6q7CJQnDd+xFS1M4UrJC+FxkVwlGkA6tOsPdTL6Z1+K17n2H5cI
09sz4hRxGHsd6K5Wvg2P/UYVpMCdbWKHeK6P7tTYFkVTyT4wqkGRzmroy+dD
VO6ZnPDqIca8CaFZ3NSHYznYdVqUhgmzapY/4AlV/0FCBWyyVsqboAG7VktZ
cJQs1PGo2DoTe7uihJZZLq5rr4nCG4u89Gw40Q5pL33m4wywym/XnDXErXab
wn98rj5cenvVc2WsuEANZ9PSYjJRfy9C5rLqsDy/+9euV1KdWg+JPJRq8yb/
k9rS8dHb3SyLerH4mj/qMbESMw7pg/suj8+4YEousjln4ytyxssYgell/Oyd
YXsLS8QEihbyrD0lp73wLlC9csN1NPsIlm/tp1AsE8ooX+FnSiBIr9udci5J
3y+TPER4KPe9VsKt8FqzptfmOqmeWxmZpPUMjco88Ql6Nm/uL5P8kXyMIryJ
HfAV74ZfGnyYc0RKITU8Dtp5dlhZryTUaXdGeXhlqnlx2THHMdbxLYQLv4GL
Tw3cURnIKg/AWPQdeDWX7sp2FBax+4lEll5NP8VodePVtZcXk33AnjmUW9is
A1vFAfXBOGw0A1KgXS7YUKz3chr0vCPaIUgswSlmLqEHc0ddoEzUigIDabc7
seHhSahCsa1vDTFANSDqY5N2a8TIK9t3UD9o+IYdwiTbP/b0LDbWTaRx8JKg
rB0uC5Mw7uQdtW6VlsoRK14pDGhOTj/EAsBpVoqjjPitV1d8zc/vUZfm/W9e
JSPSYSVF5Opf1a/D0GIuclbTxNyfCkAj9S2jAT0Qm8DxhIYRikdqXLg+WEz4
9SM4xNFaFrT3k++d9bh3g2RU/5PL+wZx62xlerBJHTqIsFqk+0cEvOlAVSj7
Hd4nJwRpfUu5j6fU6gmzqiRXyKoNkrzyH24U9ChvS3kNVw+8IWbbcRlHN3yj
EoNiAPOQC8mS0uEcmvmz6t5mpMXPcqPdpUbT1A04weJPIyvc7g6HyNQ/XjJ3
hJuG0S8EXwzkCwtBvxrDcnXLhwF/3R+bKPa4rIoRVbEt++UsgvgETCpGW01+
6RwYRNbPeftrgz/fUlXCevX3UPOwC0QNH/KhONUbjWfaeHBPe98L3CUEfDI4
Gc5NwLEuOmjeMLNgVb1nfJQEHqwHSbS2ZB8zLOvoPikdg8M2te13bkaHSB3H
eF70Q4VTXvRldnctViZPHzo74338G1P2gtdbxivI5m4wqZr2ipWI99g+nAcd
a1wn9Ny0dxcVtFv3ikYo2Rf4+zDkW8jIeiEnpI75qbzHoNn3yJj1nsQj0Vzx
7a1BAuV6smPVNeXroiZu8qxQYu+rFTc1QB7PjRGQDdhaYlAfhaOIH1+0V1eC
um/y9ghFzu1tolZH4UepoQdWNY1l5r6LN8YRYcBM/qZqcD/bqe2dmTGoyqXy
PfUZQcIvBD5fts/yWFyRJk1Dsx0X/PekoJM8Bloejym8hyWyWKGxly0PA4F2
EyG8IwkICzJS6vqFqDMcEPQVuhntcyna5R1p/g3xafzoQL0CJMPfI5bj71KM
UkA7ZCy8wZO+oiU5hXWLCHd8AZsQIgi0bOIX7HiSccLpPSUhoRV9CDqCifcx
Np4mIBicaPPgGh12QQM7su2fq/zsjX82xIwgd3n6eed3cKAR+RUI009lU6iQ
QUU0KvZkfYGM162YD64VD00xB1zFrMd39KWt9E0Pyvm/1k6AhrKfWN8+6PVt
venMKh/qjMYo2S4nwmTl3FXNF3FEOl1eCg1TuTJ8xsaTp8ry9P0gJYZWSmK9
XK73Nizz3ejzvaiXbGpuvxhYfCLaDd38GmUyGcBcCUYh8NsQbUmEmIkHQbY2
GWjG/bFucRhignIpt6Q1SHbh1GTcSckR+YkvZl69ypHYuqHqIEUy/Q2Utq19
XLtXkyw4zz18jizWqiTfQfF4Rmp3VJFSUx9xS1k8SiFV2YjZK+qmIiqebVTk
arC6ip7WoLxderjrkj7BKLcSkF+aK0KXRY0sIX5aSy6OfLqJ7ClG7aC57uSi
YFFUXIbIN2ISDHuAFdORPRuj2FDQd0oEKOELSsd83YOe9Qmpw4VWgkvxJuAa
YcDeKMRyb/EzrCwjmfTtVuxN31okq+FV2ynXkE+D+9Ng2XH09AKqYazpdcP8
opg6cE0ELAspv0mChmLzE75UZ+nDyjpf6PpwQMxA+y2zQiuIRztACH9QHT1D
OfxEaAcQ0zpEY2CKvFlMv+fQ4gmTlS67s3be4CxDQ+G1S1McDIRomBsNp3iG
FJRuzE7r0Pe9OrUcmKydLQK7jvaCuzmyeiHo++J1X3xyIcrtN6KBFtsCumcs
zfNz7YygOJ+bWeDZoAyuzbx5ywXJ3wF5gC/sPkCE68Ri6IBHZiVNXwCYzG/p
e+LdJvruxNTDm1ylQjs2gsolOMA63LTWLGt42VUdkSto4bIl049RoVqvqTGW
D7xNKL7uxFj3rM7bLBajW+2sso6SOFZ1TmNpT8eFCLPSgWiZLs/c9/FL1ZzD
KdvWWDkibujKf6JIcI4khoMu8FfCDEgnWNWmkOR639wNEAg6ZhIkiJiIRvHy
21he8EY01aPY93ZEMYWkur0NE6ksdD9X1lM0gscuW8Bn0AawQXR570nKL9Gy
c1jEDkqWExZ1LORGbDg2lJeP5aiKjtD3kutEdSRXCpQkq66GIk2D9BIOkMHr
71jQYGPpmlq6Ohs/S1c4eeYh0hVjkLvvm8qa/ofU9Fz3ztJDd7es8Us8V33I
snboWb0ETn51BUo4XJHXVQjYk1RZG/1bwMk9zZ2Mw0pC1x69OJFE2EGKD2Nq
+KS8Vb5eSjLzuL1ZTRBSV8KVh0N6QZMOm89xWvygUCxNu1+9kfIa70EDy6An
ulecGZa/I8JpEedJIWNLkpWPOEXiUxSA41VPe/9p+LzCxbtTs0w0TBraTAUF
zsTfbuaIrp670AjoK1JFlYhqpZ1lzEtsxzjZLIlc0BYtgQHdShL4VI27uy6l
TR39KkaOtlUD8zrcKDmyxVR0eeVI92C05OyZhaziE9fZ1cDsu5rQ+lYhP1nH
HlVK8UDKEg8nsq/oes/yUpJmDC9tbdWzCiLeZAdXWN6J/a6TqQCFVHGsROOx
n7TT2+Cln/AfMsAMe7KFYbIiBqand0MEDZqKonwBoRiW/2H5QppHQDgSy7Zs
OaJvTB9+xs/lybn/C7fc0Ybu9kKNwa64gZKyYKIvHZuiFrxXJZa9H4MoFa9W
/Wdu/bLSiKsIcbK/bk1gvCDCJASjlLvHWrBBJb/9SmlPprP8U8LgzLulPQMb
/XLvZkLjfMI394vdUAHkhfWMQVja9UtaSRurMhF4Ar7/tllPabEbBlQpdGHx
Vo65iNXwfdnIRm4BFoRhgfLD+aEq9dFkPPi4fCMzr0HsXyXkj8S4cHK+x4ec
vMhhfEYu90zk5wV/eiD0sP8c2EP7EHOxzF4cUWob230t0fYfEUP2rM4L6250
cwOmbm7mesqWfizPKlYNWdfPuwoMvM/hI38Rha8SAPgVTKzLfU3mKNEzUP5y
0M21MKtxtCB1H9mVwxQrdTSqoX6wgljjVKh73Rf411EoRGDneZNn1xJ73S1/
la6H9rl4EQvsDxwN0UhfVc9SkfATPfUoMuPCwSTPCgjtIazEBlz/GoVU/Gpb
t1ORKrIDMXjWsiIlad/E/xyG2XQNlpk7W2tlKE4hELnwLJrpZKlagCb2bPWV
5HF1WuK/B/4D+fyVoEI1MxfmSnqe46R5o+ngxKBjSD6vffD4MI1qe24EMtyf
yZ7JbIbmrj71r1pBhO7qOnD2BU9mqxkm0LlpAIrfWM6Nhng4On5YDBH/DIet
gc8MvFcIKP5fWmYswAXXkSX7qsZhY2HuzMF0eEgaH9Rt5UXkAuhtVoMUgeSF
0rYs72C3L78hUhKlPhxFwZqfvCXKvAMlF7X8bmRr9XgnyeYMqgduTW8WBga5
o+fMAStvjNlyrBGcLNWXiU0wcJmhiDUb8fZyNkl4O0PFcgOxvl7+Jf3mkCNS
hFiwq3XYlzSzZVsSoBhFsXfDtmQrcDHhvHGDp++rPiXuD5Xp1teal1nl0TMj
WdNC9r5jpf9jVx88IhNRXogHO92lZCexZXM2+gakx9/KgXEv6Z4WcPfMIbFI
BmROJ6lYoVCEEDOepXJcmRpo9X8TAGVMDXZFfVJUjIlQsJaaFy7sHdoebKoe
kEXXKiweD4MaE73lWvGr4b2Q6x7K6VRhKdCKOPhI22qzY1eHDGIlepaiNMgo
Y9p+Gyolcu16davY0qW/qA6iwYNyNPX0wdiiYABNtsqH0jd7FxCDIRxkhEOh
L5FP10jyj0+EZ6fHhapHv0zMRCC8nvMzYPBrsywzOgdE64V2CuTe8V8ZTD2L
jgKxlQ2vEPYtlTjNrcML7WqCqZ4clgFpGI+jhq7A6cS+0Kbh0VQT/A4+3hWr
cs7O6mbBakFQxUpJH4Rp+YfMBiE4ZQ+3ePVMRoQmT7MySeszWUnn/Tp/tVAr
C3wMcqwDKWpPTfoz3HRG0cMm+LJbiJmUDvv8e5Qs6+GUV1++E8/F1JS8JKAl
PXidxR4fG0hlkdDemsUSP+0uVy7fvWxTqi+v5ZJJPuh1SUvBUuzL/U8E8eAU
S+C+AmCDZ2nB5orAJsJDlg4007kWG7kVzbZCzArRgcBBNZbTbrRg6lBtCgAN
gJo0XxeHHAbOB/jf8y54gPp/SMezCKl734w4DRce5zVCbgqpP07tyTrkZb+i
kqZWyh+M8+VbWD7Lkw2UTG3SY/6UH8tHMx0+or0bqViGnQVg17fHuRaA4gSm
/m4UjqGMJ1rmMWYtnLjEAsWG2/+yQOG9UtzI9layjoHCsq1mt/QfTaxqVp9B
sjRDyXCjU2vvpZlMul7cBPEdwj+2GCys1T+jBujxjzQOrdGC/Z5sTD+xQtrD
1uFP8tieIkrYPQney6YrxyOHKKLwHI/2uwyZ0i/eq4CAfYkjY2ChWuwv308L
f0kA/HJ+BLkCLq+VjCO4wwVIGe8l9F07q4fs3Iy04+pEZ8qJur2robqzlItm
zgnhYk+zfhGpLUPYpDvhKuV7V/qs5Dlsr1fRHBFLCuPDkSqiz1HfcLQnOl0v
LrklRsokGGRbSKfLmEyBwlZvCEGzpt+md++cEvX23hNSHllir5siL/7aquS7
RwDmlTlJcp4UbOp6VQiCV9FMUM4AcpnHKEaRzf597xoLyDHMZW8We8chFRTn
8OMrthuB4NY6x+tZ8sLReXo2n3YxPOuzgj2q/NXH4gtc3+T/rLKzNqeX4FUq
cDUO1Gq3qSBMYvzG8UPMfRJHfAy5LEwVTDkUdJDQqgvTZGViJb7OD5HEKg9B
Km+ss5JGl18lUAUMlNoF4av8ZO9/gszZ3GOcRqUTsZUktH966mY0GMKB5leY
c5tvI5MNhfDZY5CDOfGIZHTeCLYmDOla7CG/y7UzCs1B81i5+MmrfSFkJdRI
HRu28tMwDMY8jDszTz/PKkEN7ImCrxA79fqeldiJqRCbO7JtRZui1MF2TVI9
WCOjgW+m35bVKTqFaKO9FlRqVO0YfcHzAZmeHwYB5rCxN8qVF9wbN2F4sbAv
LLfmajcvMF45kOd5ewo/+AIaVHWeRax7kPCQi8qOkipKrCBCHAedO7HapHIa
r7MwpDo9UHSx2Dzkn0hpDS1OGSuCW+a8GUHla1g6pkrXkbXkxIttlzNe5BwO
3iCmR6+Z68f+2zbwFuF6vQq5m2VZZTs4Ct0TuUxxuhxNDfLjxbumIlXb+Uyt
okWxeVWzaqFmdPwIQyjoH8j0c25boh5KVAY/0wxIOe9s1z/KoxC1+if7Og6k
XKEGLQ/IVvjvfVHRMj6ZsEOF4hCvN3U5TVSD0H5MCdhMLqT27VD47+raLYmS
U07BgNiLfMSLet0feusAwLFUCTdcK4rV9duyVfz9WGHVZtVFQIf9jCORuZQc
tjxYDPWFi1vfYWu0adkgi0VfpHvU0XJ3DaskBKOjh5kv2Ws8qbDBuXJ2eB0B
e1fUY64CG1ZTDhijLWze9koWaqC1ffQxyq2hs7UMKI+B6oMMhaVD1dYENbUM
pYL3p215Rxqb81ktbkH6mnC6tyk/Jt42afNUtQfM1BtG6GQZvpK9VGuGURJv
ykFfHNaOc+JixmdPYxvyIroSafUnSwrUF8Bv3mJiNQIaf5uhYBpvcX4slWTf
OWlV5yHylrxNo00tUuHDKs51cZiukqOrKawGvnTdJT17O9KZ5vZwJZI4pdAW
Y0Rz5FGZ77CAy3lxF5ThB2SY5JXciShuB38ykFye30oXMqkzCex1ZrLHfqKS
LYVenERKwkxSD4XmIcpfJgmQ+c5oPJnGMcDWo6ayRjTJrjAAWOX8uD09lY1Z
UFoLLIG/cwn8yC4NMRwsUQDwqBT/AgLghiMy5oHmI2xaATALmh6rNosbSKPJ
PSe7JYNr4CdspOkgAYpDnpioJ80f1ROO3p5OGDLUBbPUTdDZAW/8qQDIxPNZ
R0Fg6viPpQln8mqBi2Tro+P1TtivfZETUe8BknLWWGA7oFL0DgTxwjrex5GG
5dnHWMH44/TIBv9sxslAPO1O34ex55a4jwke9CHtFgPtkoR8F0INHL4ucIVL
Z/1opP9NPb4/tGBnJUZ4EzrifzKHeW3oiLWB4Mw6cbBSWrBzyeiBnlTi/7GV
ssobxbywPavMI2W5fShbSwYT6pBhza3gEFx6nQkAO651450+5BMSyb/CyP6S
x3zVEB46Fh3Ljbafn2q0kllMwDJgXncWxLtWStFxcH7Vww1piRGB059x9kID
NHOKncNovbLoW5ZM1fQNgACptQgFX/je5L5sGt0+pAYiEoqjdfxQL4oiDfmb
SiImc37LOnpQYvGQKoUR3lcneuc26z0OIDRsZms9FvYH+xcr8A328jqB0EBA
skHjelxzQN01y/hIpnJ9Mzv4SO5pmSAn035t0p1iYz5Qr7cijzq+l8+GLs4T
CEr0fK5DjYQGG59ssZH/qlwGvTlX4V16bFevliVHMQjZ3wO9ySnWQHs2/Bw7
ajVjnvU9+ohRSoMuS32osVV0l4myHoldqVCpHdt9E2FLUEdrRI4N7qs5GBAq
tjU7F/0MUHtc0na5xiolXWI5bQQQuqjNILg1rBLMEe7848KTLZFMlglgosmE
HHxu2xj8yuNRVqbbve83UTPlJ/RfaAW73CseRdPEkR+6VqRnAjEhFPDzjMui
KaDvAk8lzT6ZWVSC9rKKQ/jQDfZM0SoWszmroS372uNNb+RW6ruu+VhAB494
SzLgDJ1fXFkwWYns1XvZ9ANtrrkoEJDCGKKj5rgSOOOa4/HSbnMpoScRE1jp
QEsH16Q5lKkJ5jbkf6YhksXMG9KHLbiollcXhFW2IGJHu9/rgtsUM1W1NKX8
kNJ1qOn4p9S8H/GMOJxALAXD5B+eyqslB/LNT8NOm8tGOg3GuBMC8UCKVPg4
OqTFC2rvfBybciG3TWi4z8V7CMryRrGNMRkK+SFqRKQYVytMH2K6tBspqqdW
6fHkO9PWGIckJiN8TMIpRimPqCf2qL865m+9NlNToHNkSS9TJ4m5K8GikUxZ
/JF3xmSilUbP39gkNYEoA16CcHtSN3Xk/fduUK71ckxFiQe5kWS1VFlY4iAn
rNUZk/yBFOtMaed6Be9C8/KTNCjgjHEBEnvAYCQJ5g3I6Suc6JLekJaQ4RHj
ZsKVzYcW5G0u6VN0eDTuFqZ+/UBhYanXD0LrslZ9+sHv2ABOHlNAqWoGdnAf
YEf4MMqjuBI4R68xZoZZyf4IbTwKijh6St2ZGMYOCATXuEVG1zWQr45U6wHw
jTZipCILkcD69+X3ZLPukwlXodKPNJy1w4o13F2ipn5T80cqRYA5fvA/vL5l
0ydt1tIbSdOSVIpEXe5MZCWqA3t+4srbi5baGQregl4g4Tu9+1FlhMEANAo4
IyDSD4TyfOpQegpralrglc19s4bXKdYT/C8P5aN4LIKtRWQsDBs+9dxOsDAn
czD5/ILQwN/68kUiY1sNWKLW7mKm9et1opAYDHCq0aHL1SEYgSmkni0l0qLH
XPl9eqDQNYbzlhAiDrKJCCRyiv95mN+drQ/VgwZufKh+qULpZ+C/f5F5PCZA
e5qGomTi2aehqCwkvd/zbDeBCmmQGobXCpndQ3MslsYBsnLiX8z6qZdTwF1I
1li4H4Jei3lyPL1Uj/ZdT1fg/6DXoC2Xm6uYsm37f72M2fgmQLIxy/+chNEE
jZQjUexzmWTX84Mf//Bf4r045pDA+s7cvs/z+cNB4A8lbHqaJklAdZEGBOX5
NDNOiNYYrsv1hz/RG+WTClnG+0zlpQQJkjPHzHA407OSYzbn1SJm/DSWTe4X
m144Z2Wu/c8Nlzdv36nheUFvu04Dffzo4tR4TR4/4LMcgiaJlKObZuzsFLrP
e0mT38+UxOujD4rYWd7p0L2LqqyZy72Jkv24QPG2/HEkvjbadxqsmO4gNfDO
at7yR2dCgFUwvNze233lvbVNg0GND9ZYq44kan297d1KmXH2dQDTJP3F5OlJ
d2z95fl6yr15eRcotkxW1LzAto61P/AMBVekNAOmVnfF+5lK9VSqaT+kxrap
qkEAxoieHKjVG/50WMmA/483n3GUbimcn7/vR26ChIIsSwzdFTWUS0gJ5EpV
1tygN5+F2QRylc1679Ypb8jv4gjbTaQHmlaWsse1/b13+0E3P273vABz/7Jq
ziNyUPiP9pe4A2QmJOkyunU6d1E3nTCX+vvKyoBJigtEoDDh/FTN0oH9mYoc
XumgVYjdxkqj3dPM/tvO0+TqiBFEsbjhBqYf/4rj9MnQ3t0JWxzXTdA5OFrG
AJOh4s6nYJF3ppSo57ubEamdpc8zt60fIlPdKPncgzZPymXJ6xLVs5uqgZHp
n5Xm3EnxureAPgSF/CCPH4Jj/1pHBq8eEH9PlGAH1w2IBcHNH/qQYrH1dCyH
/fMosJMD6/rdVPTuodIFEOr7ixzoc3+SRevHxxeG7GPmNxrJh6xGcNEyMtJM
UtYwk8de+3Iq8tFcE26xwtEonaZkNx/WVQaM0tZP7VHLwLPmHjnYRx0KhJdH
jPQ9+E1aHXaKGt4RWF45fjQyHV/epUfKZhva3ZSNk+NAyP7jHRToJuFuGqOS
LSw5npBPoaIbgc+3SpdWEXwQx1/ZrU2aJZkaQDyFkPfzSjrUoyWbd+U0AX9H
OFgTX+9CAYzyUrpKSMfRWMtLbjn8+u2iDf8GfqT/oWM0p7BD9SXHO3brt/Q9
8Gun3gsyiHbSpfl+tG+3Ku1agdsHtIfbvnaK9fau1JGL29Utj86JH9iKkPxk
hfXfAt5742MzXacuGabCHb6Jwk5KQcQ2ZaKLQOJ25Kp8D8dWWAf3HZMnTxoR
ARLtuCVIEC93j0/qiJk3EwLS3b0YifoYesSBbVsFBbyASPmtD9mdKE9tfO4k
65vI3FGajook86+9I/KUa992VfGE/qXSYdWKFmH407V7UWn6cmbtKlYOje+7
DoHU3ICG34Er17EeA1jEsEgOIALmmVs19kk/yBu4yKKNIe8biKWPc8mFnRsR
2Sd2Wx++EZr1ZbTZhPHYqxTV4dD8+mviMbXyyGxaSPIERyNsIzCCmS30Q8E2
aVVr/bg6oJkv6aMGtdiX67bv5fTLTg8OCdRUMqe6iUh92wT6UW4kB8xCqdau
hdRySt6j0Z6Kgrf2WhyCRGhzgXNiSxIsz+smKLSJm5BxOzAPvCOFxgwXpXu5
Z5MBssk1YjfTGIfiTsUysOEaJZG16PtBM4Et8AUlkAox2oktqb84moksQHD4
EcS23h2z+KsZ35jWD/LEEmyprOinX7dl7b0JPGHRi6RdCfcr9Mg9VfHpa1qk
L2hw+8E4D2IZlWPHQbhstOPPM/kr9q3b0xekv/RVDpYMOYdnHWT+lqy0uwEX
MBCgL1Q5+NWzz+UsagHL5clOGZcz4SVzEbo+OrbZzGzQ6AYyKu9hUDR0paRY
bqsUE2X1xd5I7Ilf5bTn8lqy4ifWd0XUbCyMcDDBccuDqKEyO6WAGp9onoWm
776nFssM4teGjXZyXP6G+rpv4z+tJyxXUMKqJm96OLtvSGF/i/bR7Zql6zNo
eFWid/PAvOs1/o+JwX6rR0m/ojkc/h0whwettJVNNcN4KdovtU9SpSCghZuB
IuRa1DGLaZQepDiN3WpE3cL0kPWJ7riA4CRFKnXPOoDzZB9kjlVyRYexRVyL
9i3thgGspokIZi0shSyJC/7yrQUeVZa8SUIFd1DNUwwiRC+a/JKsQoxR2WsP
ObdavkfXfk40FoUelod/blm0z6YV0vYPtgmvIMkPnjzyvy2Zvfde/xdKdVD5
w9seBxqZ/ZLNwg7hVAu+mYYOadCgS3G4DJGveuUoPuFOnsGeqLqbffc53YvK
IkVeAYEt57smgyDAoSP2NSo3DyOoIAVTsysnrkatOGd+NxV13Px73QO2Uq0y
elzllQ926DTdT5NhtAadbH1UTJsMDmDD9swUl5gepyzZekR1jvuj6zeAxlJk
2JpjWrZD78IPA218KnntaTmzJdpykE3GS+cw9iDfxDImW5WMMzj6zzoJAWoF
780VtmGTi0LgiTGCnnoFLSAUoV1OUvu/4f7oIczSdOG8r6GvdE5hDuo2dNjQ
jTw4K6FsE6A64IxJWSwpWSvMMCmqx+0Q6MUsPD2wWAj23Doasi6DHWrQVZK3
r+F+qoHTti1jQpCbVfrbzBcecVlwbHUdvIZnI7Banj+3Y5809Uv6aNCNVft+
jWgUEdeyqARdhuWJbbhHPQ+8RISTaesZmuuoSqGUcPmNuIOl0Xp+vAqYPEnU
x6quZVcZBR+HNXSewECtVHLvplPaShP5djPRQ9nJrRreiWMyEh1YZuw7nrUv
QjWuGlkUuMPc2wbym3FldIwvkgzGDZZpaL8/en77urTHyYEW1KscJuYf0Jsy
ioDXS429ymItLQJ58awDx06xXceSWZCfZVDTczoar1+ibnRMy6xY5ZFRNQm3
dltDhNt9fs3xjw31zoPfIkFGuRtAxgGkPT1RcNaBbsTHsRzVxpKqIMAO0fWr
mKP8zyOA9lm4utWY1mPvAkcYC9oMzXWnf1izgqFjs/ohDZpOIOGMYwywRPEU
glOewXUJei/Bz1HnpGSxsrWSht13ThVXD0KlLP5uL6zUjxG7FlgCKFFfVFkQ
LjcHB6oljDj2696ZW77L8AlnwsK1NlYKG0hKTNoSRRzNzim+xwHK89nK7sjP
9wjvFs3l+Qa1K1kPeh5nwn8g1uINQ8thjnTdFO62+Kc9pUuNyeTeGAbnmbwz
8Vg6YB6Cem1T2zhMmPgLa2bp8WyaxMuiRTrNPOuPrtW3Gc7NZhwd/CXh6IRS
daB8cl3FbldKKTM8odlloaL87f1mmPCCTVpPgJSDAQSwCxlMdCr2u2FHN7qd
B3Je8gFuAeibm9RXw8LrPYUQVzPAYE77KOV+MawSmwrYgBQh1FVrbNW5nina
YKx6v57QCPu17Zm5XN/eDvCqHWhlXEnmTBqb0y6uBWspadEOfCzFrvB5sgxV
8OIR6ZgfeNfT1ppegeDCt4+TnBTl9TSCshpk5grh69CiT1o93brmvOCvR6A9
HJo4NhkFKVCdyRMaEegNq20hwQJ3+upMyiVthf8g+1lVcLQ3oiVE515DKYPV
5RyMPEpdDhqtBJC/Y9TWAHCRhR8nwFq8FwwD4wLkLO41zeXBfTsvyzJLoSIb
T33YEhwhfNaDCtcbz3unI2Atf0j4NK8BfAixQRKsbYstTJaFAGZbXb2t10rX
FzS/zouTUCQzilisS/Y29TsyUAo260ItHHaHq0XgpEBE4htYB8IBnCcULVna
sNE+tFqCcdYyAYlP2xzNR0HZdPVFO23RcThwDKtAlk6Y4Q/j24DGDhaPDZm6
80HAQGhc8ss4EeVLamOr5U51+jFH6pAZ47L9+peqwtVqog46yTsFbujws646
5D2WLJGMivfCc2dqk/DxRpnVx+r74cvBB8vwON0Hpy+9/E/EWMeKu/1g8uz2
K5tMOcBINlbkNO5cHy9JhlEhKEoNPjWrCTUVqOYba3JhXzdXteO7lLe969ss
FbpfnuUyhAx/tvAJOwnOul7kcCJMt/cWNatdBiUIsHL/hbYjSKRWKRAoq+U0
YrBHlR74gxkwV2Ow88Cf9xY0ADh8ewVwmj0M2GTJH5NbpxPhf9Vt/juHl++W
SWKiqrD4diwZqd9SbLm3JOcPWbJwQLlj0zVzzdq9eohrSWrEnc3vg1FW1l0b
tRs9QbpnCqiPF2JjB76JVw8Scqieu0Nq2EUSEVG8dGLBV2q6AOi0zkO0T8zX
Rr5X7TMJ6lNNPUkG6YFaAhzekKbU5BE4Uo6U35Zh4ur54IGJtqVTRdnPXIF3
qdo22MKVxoCywpbqj3VpPY/bEw9F2GN1mUreG18RRDhwOf94dytgR8NXh4nc
2FkazWS5xoPcYCpSjOGOfSQGKbB2+/ukAmkOZm5Pe0b3feR0g9P7MJnKNtS8
KGW9KNqLbOFeyid5kIVEAoD1HH5MhgZuyQkvci+lLCeeAzl5Edcko3tT0KFc
vMDzBqsJuRSnMf0Rdtblfr8eFUdZRKgAOdn4WBR97EXOfSlY3GDjMgpXuHSj
7UHMRBSAXWW6i2mbgngxJ4Lgk3v65DRmXqYFgbKyB/+svLzia787HzQMbBlx
/i6jVUGkNS4ffojGiGrTHt4z3QjGDCXs1/n+7iajpdR1BIboA0/io4hvS0WS
QWkNqhPo61WFk4zQPbG/wA4tFqStsiJ7xonPoS2JG80ClfIfdQyrQW/PUFc6
OL8OA3sxiDTJrAXONE8ZLX96Qid6roIN4J6brrDxwfYLjS3Q/esqBq8pAMQU
uHE615sRSXNzxJL5EA0DLfNmjFm+mEmxm8EYiNVXwZNfl0GT8itpxldulYpb
RjiVYGofj+q37Wtn1fz39e4Z7NB1HSzWh8RAH9AiuUvTInAqoy4AIvgeYJ5b
aNhhr6AX9MHxmaloZnazuwJR3besoOCTQELb08wHyvvCIjVPVSDjoDOYPoD6
RNbKX0Fq0Qd5rnKIlIdIxvqOyv8qhr7lSjszf5gF9aiUvoGCmFk4bJHwATw2
L2fpHJBbuiQKkYWJU5uJivI1k4okv5wYnDU/ytXvmNuFAQqKRjwjSrJaUOgM
M1vpUDMq3ojJ2gMya6dGa17xoERaqOv5uI0EpH+cWSdNDDt8bqK0jtAHDPFb
rEDkztSNgpbegISM2xVGDn5nK00jkYEm3ryAtVDsxOMFE1ffzv1/Y5qVBotJ
XqiT39/MWCdeB8533acZLVE0IeCqqn7kNgWo3M+8Yn+F8yegiwWbOgUEJULx
QUAkQS22w/mwfVCVVq3qHuabQ1VCTjKb0MKijSDi9LWIB8SPwGpw5+jvy2r4
7Kg0z6BwGMgFfuK5wL5+PntwFAfnghI+VjFwMhs+t2teZz/F3mY7Lq4Z6E/k
CWAdaHCoe3/wmSwzzFpimY4Lg4fFQU+PQuu49RKEZJkER/m43PgjVK4eNRDl
gSy7msAxCMSjl/cp1W6bysowHcsRv9v81wZUJLEKHbXluH1K+9v2cpIr3jIX
hdPuE9YwG27KorYTeNOn9/PNgN6mLhh/i/4eBXWrpfq6he81GLmR5RB3hXLG
WVoSI2KE9P+1Zl+PVkEgZcBsNg4csbH3tYHLXqeLZ2d1pg/5Y8NDSO/CU7qq
ZobsPFHzJg+ktJmhf/u43gfnUVImEWF/LdltzFpV9hamczXkuqg4+TXH9JpI
/uxQd0HmJiPDrlEBMTUNriaJ2z6l9ZqL4l8tK1/2y2whH/KZb4Tm5MpMnti8
xvhZnzuEPZdZ6DrRcMnq8A+fSRmdEY6r3WMnpVL98/VLNpHtQ56XHyUdXJs3
vkc/84rWYiVRFjJem5MG4bWFRtUZNqagBNU31cWe7qY86HMulzjfVTNYKxTp
KaAPE1DbTZFGq3IneoSJhdylCBsEGxJAf8uC74Vwc1OvtvUFUyt512JlCl1G
0GTjJ4c3ziDfmaEc9UiN2ju4ZaqN6OEuM1QZdObeaa2brZcJrlpPuM9p2cOl
lubpAgPSvn/Km822ta9a9oVnRUCQm1RcojnqezBD/sjQjpZ+WrXs7ZfeB6TP
+1gspvkRsNZgd7jGr8pXvevnmdLHyLW843TrYU7ZZRh/JttAxhwuAHnTG429
2XqD3BwS6uo7BSlG3IntEEfax8cR9+3J/9NPdS5cgjPSZpM2qMhT4bUXKqL8
R6udHXtX4nExhd9btCFA2ZWpZD4cGgV1dceu3N5cHmWzq/Kl2RXZUszh4YJs
v9K8xw8OOXnlUs5xskv6SIzapHdR3MTKNa4KbNjnAgEXGIRp6Ld7Xgmh9Bmh
EiIjSAzJ1zwrP7RWn6fOvKj08/gYQ09MYM44nYXnzsNUaqcdLynRz5zxBjeN
AOHbiEMuJP9KRdKTvh2mcDg+o211mjUvSGlOljrZQHP27n4lpeUt81/CB3nJ
0gdJ/Vq3n++KWLd4ZyT51RB6s+0P4V8aETQykNC5oFNtPEwvRRWjShnW5DLG
mwohmE+neO5KZpzXog/UOMEE2z4TiBUzOuwkzE57+NbEnWtdHG4eBAJUVkfT
vVewkRiyNr7lgHyTjWpekGxEQrOdd/FpQnHEhc++CoQcizNzooI8T6/ltqu/
S306pCxfIUiP8W4yScUM8pBZ7uzI15hcQ7rmn7s8AfpLw3SHw2Fq6CF4NqvY
vZV93lDxmL/Yhvi0Ys0JaIg0Q3Rh2rJwofQcT6oFbYeLTokX7axYopziPq4R
1Bs7pf091iFz4LDVZ6AA9eU891Ap7FUSxwjGs4uV0SNZNw9H3vhRNDAICdm4
1obfRsT8aF1wodqY5lw98isEpxtD/jthrGMENck3d8q2KhdWQ7eyrs8R/4Yy
Lk9Y0DPH2nE02zUSShgkUr72inE2kiR77i4s2j5VERRj/dK3ypxL+ymaukLr
gdH4n92LuvLdHfRz8O+HFxutFBrz+Vego4iw3cKH3iYUBGycZb1l/aXfRBHA
JY39zfqxHZoUFGwK4bY+TOz06LCidaUShgu5S/Nxz3eT5kKS1rrH7RpzhUF8
KSGBGLIG1PIm2Ylh237czqEPL/qKJIh0SAs4izik9LL5Y0xJVDJvKFg8TV39
m5tyeH+gHZGeBUxoL7emI9e5I0TIw/UToF0KGjf98h6hLtAk6l+UIxZ9xE9N
Oe4i1DE+p/QKaQEmZj5+5VtzhRztXEgGcZEglinGoLOqkYk0QKSm2AlbRh0r
QbDYqZg0UtsdDBdWTU41+MOhfl64jYFeuJrAzEoUwzKdBrUYf7Jgl2mlOVez
3Sivrq6nWbTEHWVqfMizFmsykv3OnoNAOy477ASGHonLM3j1q+RHandOLPgf
UagBRCb6igoIGv228tRQY67D01YPYCaxakwjMZzxlBEATBW3Nm2ng43FLknp
hWi/vil1ci6IHgyzurUZE6HfAZdUizyOuUVADeDETtU8pFVKGeDwR85CB6mD
CxBb+G3B7vVrxdOUz7VBcHQz4O32vVGbBCV0EMlIolyH3boBacZIpk3j9PZs
j/a4qjiYUeB1taF97Qjocv0Vw+VRK9Nr25gBrS5joU/yCsijT5NrUjdp+PKN
X6+Ks8ORpHTp+SlvTWDRISkXCX92Azt3CJalFJiVSR5jDOJhOweJNrsSK/+H
88jK8BjAC7SwINhf9qa8HZm4GiAWItqpV+/efVeXs4zThDSWYLiwTu3Ldw8W
gwN7xomposDV/tVVMDr7fSrTkJxVt+nrC20PzDtGMoU/KFIotc7qVAAd0kV8
AUPn1vgjw0dFHPFayXwmuw2xgMC/ngGlk96wJHE0HAooyHGoSXj/3umbB/OO
8FTVucjTGpJBRxW2P+Cn9ViumNd/G9VJv39MdbPSAgEujs6C8BU8EDErzcvz
dIlwr74R91066ibvu4T1b4vLsVyryU8jap5XziB+GbQ0M8DaRLueJv0xIJXe
joLcK3SppdV5cZ3nFdV9DGv+PRtp9FdpTDgK2fNTQfK+qpi8k/kiOV3r7RJ5
mBVUPiFil7lId08+e1meQB2OnQxYtYiUJXIhAkZkHRL/6LJPpO6jx0Ih+P8J
zoaCgS/p+YgkkqFeC4C1JHbAHGJ3BpBKngs2Q3lCzaCEIhIa2znbSnQ5pi/G
NvkwFMUdLZZMzF9EK1dpkvlXhKV0DYfEwSeZj/+YAAo/oi2BiYiTXLWn89ha
m5wJA0nU+nIbilZoJTwW1KlLGZbPlDMTiTAc6FuYupX96egsn3U2DNnGMQ8z
My1f0i56D+x/0yR4FYZRwnCdfqgUq4rJRlZwchsqau6kZX4DlxHNvW+F6N/w
8O+RL3N8VIcMFwPUUOZLmo/WiA5JRgoAb458TCDL6WkY5LBoIhs59SFYBUOa
oENPsp8DW1t4rqk8EswNEIdqAAM2XkYhf1yZ8ZmdJ2uociFSLtJaofh3qMrL
V34WAk45Tftvtv0Cl1Wpe7tguaMA84b1KKisBDblYHjNukfn9xJ9OUG+8ZQn
sUAEiQHHQzpB+L2kD59kQq3ou1QbQif95uXIR393Q5mOp8zGQrAs5Ee2pIPT
dNkOWS/tQUsFjAhr+/a3Pl9ud7APJpZZjUgOb8KICd7soyLwn+F3nlXIzJ1Q
RVuGWdn/ep7qTG8dZfJBFc5v+ebl8zs9N5mNr4uVUWAXkq1YCLP5b9gFzErg
urKcrA4jNJDygLhJGhZPJtn7V185XRUD2LvCSuOWQ74RgvKfxvNUKYROGeko
e55kWKI6GlNxkVy4+dwumpZtLfxtkJRoZdCIZVJs5T4zlVI1UpQ7ftFkWZk3
BBOd5FtQq4jOrC3S/DCti9CETWsyYR4dHS8HDGmS5NfurB5l2b26l7LLqldg
0siPwDvJhJALhXhptABFmliJF8mqRep71Yl0Wf1h0OQHctx2KvGNor7fd7g8
bDSF2grEIicF3YacfpCJz2BvBHF/lqmTYvUksUyRMKBuFESuchzAxq6NYNKf
MblUSKxBtoE3rEVC8HQSB7uIzk4TZRobQk2y+gfQcQydgT2JLr7uteHPkVwe
/Pu0m0W0q7HpSct4y4Tf7H+MFoRdnkQeBGFxTR//b0zbCUcuNP3OGsWaQZ0I
kQ8c40u2dukfrV6hDtoR2zK0LzzBSBePIf719RJ59mAjTnjKp0uSenLKkTog
1a3eTRFan5ZbJTyZT97MMjDTUtqZYxpSwMxz+H/+cWMXFbH8IZNnzL9jL9Lm
VJ6kskSdebC5QmA5+KlBAJVKIGSGf5XR747iCsUDUF4LreOvSLr1MyJKgxAu
eGY6czxPLx/TmIcRA2qsKS8oDUlWDPjA8dW7KPbA2Ov0rLJ1O3C8p1v8T8Bl
68zlpSUG5OAW8SGYvqX7v7ZA0gvlaEgUFXhpgUcLHoOzkvn4ApLVl6POsHsb
XLl/ZH2K27kmlqD87nRS44N+h3ETZYzCBjHa0uhy1OwKJFBPHz4/NTfwIGLH
0bu9e4mqcYNXbX1HAS7TbEU6/OUtODITo2MiqS9nIUYkkfMG+rVLlncGk7+6
Ac1LirZa6eMzOkjBLCzgsOgutQOsnSNQo1IGk8P0OTAwBCz/2/7X1vL931mP
1IW50GZhcWV9vL8dvQxiDctI40CVF8fGvxrWNUx7VZHxnRLd/Rzc34JjePYy
yxlbO/iq/Wz85aWjKZ6kjc9QGF7/0PA2SXYivUohL5ukxUPSGy0xGgp4NDdP
zUZQmN2JATgiXZFeS1BNZmzyXpsgh94jEZwYMIiTu2afcm84xw1cSQHTsVY0
5gHbNttntC0lZKKSfj5dOWCBnkuhp9ROltRaPX1JNiWLjFOB6bFh01Z4eT6G
eAwY3fMgem5vyO0n7yCgFNsKogJbREdJAPtf8MF2ubozZaEMgoSpNeeUgt2L
hr4AUb3dY91Ght+yzdUI8Ux4Td+JNg5bmdG26UEUh4fQT7gVHmjAvpiuDFIx
8lk/OmnzHj7RwWQTMZdBoETWJxKEtPSPSBBbj+VQkosZCWBt1GKp41u1n2S2
1XMmqjg4l+DBr8BZTWCO26KStLlrRb9TE7CxbWPigskUFMfPqeGthzkhHNUb
ZoWyrajdhSFZQNYxfnBDC1hvohGmx5jvoNSwtuczHheVeuJrfJ3xZ8DvbZRQ
HdTVocQp52ruf3VJgF3AfeBWQS8dKsWuowOSC1DlKpKcI6q4zJOeDblNJx5Y
xD0KHprP/mQ8Kss4sMCRfBJggGSd0XXPW85l5ioryNx3NPd9G1rq3N8U+e0n
UWUjyReCYozBPr++nPQO9W2mQfalnf0HuJUSBc9/TMrT4lKSIUM+uWV6y1Qn
poGgLABoRkwR21IKN3zJyqEotHzkwFb1+I/4Paf3sYly4+HQwVcKQ6fUmTT3
m3s1yj7Q26hqpm2dalTEoc1A3IS1U+8KSXmyUbwkPaFCUL5Xej3phzsY+kmK
wBHuS2ntUJ5duEYbQ/Tm+CRVF2kIrZcr/2Zv79R34eEqDAdOcm6XnFs9mOzf
Fdy1abTLTxnLRGwmeE7H7XU3oNegpOSgO+a/mf1HpfrtVhVeVn32Q6Jo2Jfk
E3RJckyMjHL/9ghT4TMCoSFFRfMHFMwd30rBAUdsLkKhKustrbJV+Bj3hgUM
dI9ZUQQK1hmVSsHPCQxgIeq1EXX+KrvhcEw1XEeuXl4xzAs9Z2L0oAEZAdAD
qZAXkSW5KZqIiLyJK7Q2VrNh47lbmJE/6QNa+LPBqM3ejpmBbR5Ni0wNCQ6n
fsC6dSojZb7QFuYsTQWDs4vC4xI3zUKvOTCPp9AeGmpcS2M+qc0iAH+ZwhAJ
uTpTPZPbQoipV7ywz/oi+DVuWcaM5/DRYpxAQgb9euVshIkknW4zOAdNqnqO
y6e90QbqCWZxFiZSk7eUh2arjl2WEsRIR9OpetHICtW36dOSLyrJTd/NTdLl
i7pyN33NHd6mKTYmFS01f14LouPM/YJiJVOurNimmX8MYlfTmmOLjo71k5EP
aUfLu1SYMbUASVgJH1Y8GGuAVajRNQR1R/xI0hyzZ926nWqwLAC0uCd/2VVp
GGFQd8+rHFbskUOLZ5WHlISL4rCf06+YwD8zCQXbPHTQoznzWa7uY1FCqsHG
I0M/ikyXgco+pwyJ2Sl377G16Somg5Uscn5jblGPkH+fLRHfMkW9m013OEkb
cprT3QUWtk+F8A9k1nfxEuu9qjoo/sI5wMNA9yBroTW/8yyBT/aRWwb8eJst
fs9wDj1R5Wjg/QdH0RKRIOIhL130kczUL7/WO3piwhDe8DJDzaclCMlBwviZ
lOWPk4awLvjCRh1czPiYHzHWVRKiYrozzquSfq6bW5/axgtu1u6GkntULAei
WfC8ui4H3T2R5It3nO/Mv8b5RiPCKIcVZHXZpKAAMM/RuyC3thh9gBtbwx7d
1gzHLqx30N0jrpsvoo7Rcw79GLfXGe9Be3njp336pdSO53JWxNYISShd3X/M
6hsFJHTHbR6B07EtDuNOffuF2YDQMpoMf79+cBsgJT8s4C6sU8ImZ7OVS853
36rmb5S1XFKKDZ8aX9blKG6TQLHfKEF4NCCSRxIDPWgz8WHw32j0Ze8HXHea
VQfQtmaDXT7FLasN08qOSTtKaC2qK9ahAsT0rM5vAPAy7+U7ZA1dRchSyANp
PM55mlPdmM8pBTW/Atkxqet5Z6NmZ5AClfVU/dCnN/1PCAPuyNh2eoNIi0bJ
kKCje650jF0lEjWMl+uS6UGc6r9Oyhwok/xZycsVXQIbII9MOrPz7uVckYGV
Jy1knehA83uP2da/C2pXBeVIIBoEqAtOVF1mcS+m03xf7QiS0BhtfUf3QbpB
msM7a0fB77Sd89m5KhcIWsW8g6ArgFTVx//X9pkwV7MtWLHhbUhmHvrVWn9Q
gGtE0S5SyQOMmeiRK67vekyxf2q71Jd3jAfU2gbe3QTs0CjD/cabsSLJKqBR
WHKVnH0ITSLEyP/SfAJwNrKeaOl4+g30pcY9trtTpmRjP+guZ7I/bMd2pGAG
Gbza8ZdJRirt3mfvecSDeGJ9iF44TQiRZa0ecqd4QDrsf2Q9f3/ZOJjVuSEg
Tew1IBSUqup0ADJ2MttyBI11qpXAjQUGSnQjsMkP/19hyGJuhY6zFCN4V1al
NoAh1RBDrnKZBeCwgyedtV51wut7PAhGBZkrpglQUrZR57L9rUa1WtJVoSeF
c59xENt/LEnavvg3UHmKw1Slex7BX8Dhad069/4X3SauYWG2sMaod0oGD1T4
Wr4wOiXItfOy0oDPpbGNXrKfFrJ9E9nfEzF2EVP8MPmM9Tma4e7GXDa45L03
+W+TE8IjvD1RHH93X9eWSmW4M5InLAQ2K/19zpnDt2S2Wmid1tO+WnYV7M/P
x8db5DF0T4sacWVhg3BXOy3nFhopg59e4Nepe66wrH8UHyMDX6+b+mpWjUPq
xh6303NQWYMjgH+G7TyorNIJ48Cztmp/akkoMZUlDwJyrCm8kUKGzgHHk+3q
NGShRjuOCwyR5kFGvsU3WM7vIpwwkSOSg98CR40XVInXMdCLJEtCIxcvJ1xO
rIUuM2yMJKmVdsBr/iAHxxPQT50zWYbZwTxA5K0Yt3MmYsFcYQAVTazXZJjo
vAu9xA7pfVSem0HVMCmD0rkFQ/ZrgB6GC99E6tCOjrhONkUc2r70yOLrdJLG
qpDneAA7NW/S9cegPlGpE1fhPrMtgjL7gvC7J6ijXVUcQAhW8N3KRuVNsVUe
cMcNlNhFPGCWldZ26mvaJa45/oqmeXes6yAz9oy8qkFzN6wXcNd6RlWNhlsx
G3puq6qITs/mZJfJ/rtSyIDzqdB+3g4dLyvO8dODN+ijyX88LoUbFPwqjrfy
vERpDI9FP9YabGunwHKNlTJ6mOHNReemGxiDK6iL7y3UyraamrewehC8f1Z0
HjccZFU5mAwqQaSqHCbP5AVnl2UWVgzEhqNSEGzx49R9Fhl8lIZtoBmBjpYF
VW4quFCztLAVW6S0POiZb67QLwquQLzpk3ONgmC4rXVR3jYs+h+bI1PhIsCf
uhndhxsbPz9TMhUqIdbUGqRNWcnKf7a73TXSnsFHvqQoEgkKcHO1MJJz5KpX
P3ip6uhgESMNLpGxXxF8up3UPk0aboXD5iaJ/G9/tShl4nBB9WQNp/atO43S
9eBoKsmPJfx80BsZotLTVfFWArMy/gyBayKe2F1B5lMOMriHdpOWrV7A0DPb
k7vHoYqGyWrESCQnn8fsg2pwdMmeDaH9OJZyj/P/4f06cA+TArRj9qYqkeNG
RCPTCCvZqoWtEmqm32MLuHenpIbUNZWHOAliJFB4ve0Qt0lslVqnWT+qvO/q
9gsmGSkaXznbtU+zaPDbuxbt2Ksicr9SUlomIFfcn+RGZAn339o/fMscpDm2
P18xpf8PMk16/OFr/8a2ShjeZTXRhxvT7hdid99F1twIdUJSV86YQacMyfUG
MUdCBG+PPMOXQ1Kk6MpavZqyMORlUkUrcL4CIR6JM3Ppskdtm6uBa4JmgTL3
Lvp64PgPe2MYFafq8gWFYvl55Guzq2vrrwVpPctUy1Ug910OarF8F6p4JMfA
OmZ/irGaeDng/dyffY8bBIWmyT/OANdSqyFR8Xf8BC2qQwA/xPBHfPS08HsL
xvKaoNsHOwAUjXyyY3CDVjpanVAs6/QofyivFT7FxQYgWjOtIX/tzY7H20CK
R5Tmz9LYZ5e2KkUbP2TVHwzpaJBJxvtIhyK39hdApObU7O10YqhKjEaRoEZq
OLVnh3UJEy/6VzwOn3g+Rc/j/EfcFKQzCFQWE+UDyb8aQzrWG3qaG2rXprZ8
5xfdPI/EgJZnPb1Nqs4Z4Z9PWN3vg4QmIr/sSZG5dJpI9r+cF5Lea2LG1z2S
WzFXFYSmQmCSNCRXzgh5g15tdmBLVQMBll8Ub0d/jqKZIEgGvhOjCD6QUM06
lN552K3JaT3Y7+oH1o7LyRavIpDyHYX4kS1++DTYDs4YS4nAJ50qGa2dT3i6
W+8pJjgYh3Hbo0RxtgE3/TS05KiSpjf9k+dIi4Gm5q134cjL+YG2P+kZZ8XM
X6x2uuTSc1kJskCiSPjgXlcVrdzX2KAk49Z/peqkDunkEXjHhEs/3125OeER
vrNEkJtxd83ZEY+OYpZ3kb9SLBsb8vhe2oRY+3Huerny7YFaATOykjIMHLqS
P0TcCPrin7LEBzNPJqkj+6rY5aEnpYH6vDIBhm/cmyfMf4kVkRitLrDrC/Ot
LCV9xrfAcZzH9uNVOuvCnilfsv+rPtM3H9OlGysKxLN3aAGwOOGFQS9CIeNT
bTZbx+FFM5X8KvuoAraYlSxqJDMJ6yM9V54jBR7BqEGn8sR/EWnsd2vk7W5m
1wonHu8LWg4tVUUuitj9G67ISiyqyBuOtCmeNt5FP963njFH9fPIvvhymbCr
KyAUlaxB0mwbzl79nu/oRJF+gv2Vepu7mzheO7qjjvmFt5n0zo61n1p98eP+
Dut1hXXD6WynLZH+9PJCbSZPTYqjFcIPm44niS7mbHeizxertEUy4BGWP9h4
Nw75Ib3RVbRfRIRTS++4mOU8eeSR8Wo7t1XyKDI4M04TQb5WCdQ0RzUljHML
0dBLm+4RlO801TjpUHPxRr2j7xnXHdZCsTUZrGfLNhUSJe3rnN8ToqmhofsI
DksXQ/+FAwAlSkZ29zC0taLeq3HPlw3dtQEuGll6tz19OE7a007imburL5ys
GBLTSzhDl6TA959aMaEx9kDgb4EGbxjjOGIr842/kb8/BYWEGUeVGSen7G7L
WzSqEJVGHuZQuLnwrkdYK3GYEFprg/CA6vzhpp/bXPxTBOjW7F4uuiMuJTEz
siVvi1JKTHOmZzAbZV575Kygo5ajSqFsFPKeog78dOxagBXILZVu12G+Q0Od
3Mfgy5NPZKgdW0KwPVQW1Q0eh9QprZsoTVsH3VOsqT9ZWY02AwbjSOrfbuxG
/pDTsG9Jx+ard/32TCee5HNJJA0M+rUKnTmYbJrEbf+l5MyfJIGE10c6PY1s
oNvVWV8yOhMEST2pSvG0XZzUt2/40FOFJND0oXD/VIhWrkXrCfBcvI5I7SGg
zM4YsjIrc1ykIKrt/Vv0nf606E61Oe5yHk3aoLDgN6mRIVGkoDflnS2ebHPU
NczTElTQfCGQX2SMLLI8m3hFg/MBi95jZZxJU+2IKL1hvhJtwXn6b8SQ1l9z
eOcbran43gDJrbv6UVdua4XCc3XDslmoNEN85gRmEcj6c15kAaSnLG6EycId
XqxPfrZ34JSKv5bGj1WcjR21oAQxLlIomTOcj5+IV3mv+zfV2dmzFKnqhZjv
5m1PnDwE2We5DYVxKEx6k2qHdQjzI4Jfz9mECdQI6mNcTXGCVYIFpBgFaei+
NCfJYaQKBagtsVQiDZZCE6xdkE4YJ0hbM2ex23GRd63/COBrejBZt2ZKMeQl
5QvKWhI+25Xfo5cNBtL6YRkhjhZY330KnzafVoY9mHMfBbx/E/gb3WO4VZCC
raSLtcEU6JFZn4EQIXhaa3bqJ8jPaDdYwtq4atb9gv9mWCrlyKxoueqVAgR3
jRW0wxiLzsFxuOmVVWxTie1H1p5XNPs96naKsCpUgNAesVh6tbOnYwzW1f6Z
bQpx69k5kbLZ7gahkJlr3+/Cv+NqiA4K6I7rTbpzZxOW4bwyKcdAlI4Yi6KQ
aRoBzCSyVOoU8bFW//KKT/0Fn0+pkLGvR4Lfo3KCzOYiA3ukxttHcTgCqhAm
IIDavZYHvjd9pfOEdLPcVWo1MyizkbO+BSH6pkToSNOsEC0jzivsG7eg3MOv
vckLz7TFOWSag9EiCYPOpych0Z02PkiU3IoGR1npJPeBXoHfA4sBtF2oQVTb
n1j7Vc/cITe17i3eBDGmq3bXOrCcH9qJYbgJoL3poa3JHWtWufq2wyyxLo7j
yxdLU8RlHtzE4lryHSW+ucw+TwnuT3pRbfnAlFoYiEfqkawLzfm0VMcn9rI7
6rTKcc7jVoNT3Y8oWxLMYCn1B+TcYpjYyCsOwovYpHFJvEYnM8L4GvBqTJP3
m9+MdMdSxBIk1CGauhAZrJQDC3FRxliVPbHbQDhD1tadXgldFVTAh8h9lPo+
9kPJ0MUfBU+14eEb0Wk5tawfhGA131Lml3yR4Q+LTWvtOy41wvVbuL7tDMHV
qjMyauqvdnTDGL2AWfvqvod2yu8QxaByGF4LZy48CjtcgOUR3NJkd+b7Wgcf
2hTn5f34QX3sdfkrtglLCTY8vvAMZ5pIqyWIOpjevd3H+IjS9BbU0kogJdGV
NhI1JL2nwQuO/kzBlqigjiVzcOZ2NSRNBlnukZtNHFQnpFZlgmzralR5qMvU
5bH8L3siKtcR98Fs2Q9EndY9p31U5tyn7zORo+bjaRhdG12YxGvYrh1PD2Vw
oE0z+6H83aOOzWqxB1x/X9VbFCmSzCCuf2+IGot/sCDs11/0ywJSyCYjjJ0z
Kr4HSS9ymRwcMqbNhGBhjtbr0TboP6wAte5xQ0dvdOOr15VgKIWBwWxcHKbZ
nTx7miLXJ7RFhunNeT1RkyxznNjROmVuvGbHZXj0yiDRpRQWcY5N8nb8wn7s
no3tCtkDWqB4AJYxrD4OvKzRzd3sBTdZRl3PLx/UvO31Mhjr/emIXCpPXf6r
en1NWdXw1MPmh1xDlFcSKx3Au5YlHdcDRvnzoKY7X7+M5PBqWJfsbc0D/zrj
iAzAL/CF0dVxZ9VtZ+Kew6YIW29Y0FUUO2TjIoIgZQyYTErzPXMdLgwUiEnr
733nIP5aZlNP1uDN0SDzDXXkQ/rJOAszcaTfNzjjrEo+8YGcVMhymKsg6sAL
ZZFbM89BTE3yEzLPxmG2IiFVVRugT8UFLVWHjLHLagoJtJoRM2FWeClePR9R
df66kGPqRPsI/8TWALAYEor+j57JVah3ubG/tCPDD0OwFS03k7rhxfgzHB25
gePH90t9jt/zDEo9qTfAF5dmb6llXa4vt77BOwnOfONk7MIW7qkqBo3g4JLL
42LEbBORzVahIqB0KFo0gxU32RRuqsb3C1ero7rs9SnGJFIjy1kuBJnJ6e4y
XXpkSFRH3yZaJ1asrHB3iZF+FRpBlqluSafXkv0gcHr1S5sRd1WjT7s21A/O
Hajd2b/pGT3cC+0bt9E7YRKTvkpw56SuRlFU/4JH4hRp7vIWZr1gO+kkoMTR
O8ow9L7SzJtfQJudaO9XELk+loVemn2j0+jt105wbZxNHjCLzRegL6V4oRUU
WQ8+nN3wEI8nRDwjXfos3JdvN4gqOOvWRUuRidzfIM3k+mnITRck63sfLKqc
rWWlBQ45V6hcdo4+GGIwfJip1wME1i1t8ZHG7Vt0XKvXZKhSZGzK4hs9oNhD
fAfNB42PCYcuXpFGiXk/j+xvGfqsOzYuE/i8tgMQoxBHRnvelS4MixHeXwmV
pcM7hf46Tnhq0gXc8lskNxzRwUyq8TTssF1MevKViL2WChe28Ie2HzYI4MfH
NBm8z8+MgIK4eGzrBzwxLIfVadOg8K2SlXAbfJqK1msEl1w8ddIywXYwqp41
JW92C5NSdF+ahIcD1sL1v70Pb8NaHWp91rVkOp5iWbTCnXHJbfmI6bJSXGKQ
CgfKtv5REcgxv5kofi1wjeLXitpXCZ2MtLwiGllwhljP/hgd3QiiXbjmLFcb
xmB0eyzOjg38h8XkB+7BKqRLwtWtF/0ggJkKyp7fbDPFGINB/lgX+vIaddCM
mEuBXxtA7CeMLfX0Mhvcvm1Iy0Yj99tWIqzjBt785FGMEngJ9JkS4iDMrRO+
+9vsdclfmBxtpgYlIHBstX5zAjBLNeMMzaQRxw80M4QmqmcTDzMWz2qSDANz
GzO9oiMktxfVvUM75QUf1LqnV8P/bcjsYFtoCbvNecKbSVLqz0wSTFXSeXE1
h6UyLLS2QUm9fvIQEuhGTYsqDPacMYVnajSLNN1drGRdIoCbqt7MBuF4sgiC
Mo6eoaZVh4096z4bo7xD+IGS/aPxwxHw1UDZ2XSAwaIlMl/qOCwpz8GTPuua
BDh/HDF8CHIJARSpfLF9OR3FCt7CatioIjXON/G/IQNM00fNB751NNq4wdD+
OkLa+yLulsu+t0sI4mtZsEUEbrKF+/FqkzgEmNGZxAxC4RKUn5FxmHAeEAy3
tVyHmgK2nSe1C5eM/SzTorgeep9mZ6GHneVAr3FPh3nj/LuODJgDs7eECVO+
zUbYfIIbZtZ9Ef31n2tdCAmfLPzIRj3bqyIO590pmBoaNGETTq28Zvfs4Tcm
X6FucG5DRPChoUl875MfhfmO8TftcYbadHhjDeKL3HHEYaDRjXkKQ/KCUn41
T/FB1TwvBSy/KcK8xD/FTdua+2CyE/WNzAqGeHKweBCcTbU1T5BrJPlacX+x
M//rgm35YQXcOGZz+jIWqj4B16CHxIv8z2CzHsD46ZumGgL8X+V2CaqRcrV1
SdD7FXBs7vtx5EEbBZDV83d9+OjLnX85K3pvZf4efwiljmpAlKRPS3k+2TDR
XWJIjOg+BeXn1qRxUL7dgGGnuFzvyC+DUan/7YUjW4RyuQFWPopCgWSTmV60
fpZbwUrQYLSuJbzH75Ek4C3EULstc2U6M4EeWH2bbJgM1shRhfwaURk1QZ8N
e39rg8yt415+kTjuL6J6f304mzB7abyEBraJmZeztyGI9j5EbjGlWHvWUGNf
GSEDkoUa93S64Y4p8qYAyQf4xjl8M9gT+bNRdwJOzVwG2hmp7WgzvhUiYaRW
BrKce6fREK0HmDyFGY4Hu6O7hk54dhHTiaV3sfIcr2G1yZQ6yhbBTKEyA31Q
wDrhitCbojd8EPF9PI27CEsXURnfVE84iHTgHBh3kAxvfMmRj09Na2HLxBsq
L5AZT7p0OPj/PuolQMIp4E4odU55i+aGjCQKS9l2rWWPu/ycth/Jg02t15ur
BsZM4EEw5FBUeMeYNtX5VdSWkIwvW7Kpg+sl51mVn1TbNPOlEXnRw9qKYJyf
TktUcpRe7dGIWPTh5C/H4KIkaOTU6H/WIMLK5kuIwR5RwdHDtqrxpjXZKi2f
hmEYAHOKgMGfoHu1JZKo8cBZ1NAJs0ZmO7Pg1R56m98I4inKKPb+N1mZt8nZ
oPpjlJTirAiurNwJ/ppdx4r/oaTqp7UyJ5gGIOHH8mWFiihD7PqBb05y+4pB
Q2so46VDoxV74gbhXKTNLknl+jf6JXUqt1+FK5pbs/OayDksDZ/oC/BPwOjU
J5doV3ef3D2pN3eYidY+tk39aTLQ2Uqt7l91h+Qus5/9bZCS+LQ/bawV8rW5
scm6UyNOEw1n2ivfVmsufrGfqUEQEA4IFr+lbkoOIRaZ9RPgVTmFzR0n3ImC
H9apFJ6aSJFX+yH9HoGJIIsLTGhEzBNOnQrSQzeue7zevAjfFwb/DAOABalO
HzC1P6qnfF1jclYVO7SkuikNTOOb3jP2h7Chcm1uHqX+guJpa7mexDecdRk9
eC/w8NC+I2sm82y0piamoJ6omCE2iyANUZlIbTy2u0shuuCMdxdfzpwIYq8N
IAPeEz4fVAsJGVd5UAuWmWQJfOR/xSvY0SdJCGi2oOmgIombsrFf/56mUHgY
+p3sbiifFUbEeV6fqUGu2SLl+2SKAdRHQpG8UFv/dSb+ue59bOYToK5fLgiM
1UFRFKBgbSeID1z5SZSzVW6z7iPMVVm1I706DACTkO4VRdgz/h5C8RDiSyQv
3Vz6csMVa9ncFKvmphnAXqsSeALsXCo3KVgzIctsSBiWCow/e+KQyCLLQS7X
VthScAf9iXi+jwM0OdmJajUalWyJUvdJ59eOw1Gl3DrcVpdd+OJoiL3R/q6C
Y+vU65tyZgRVNduDny34ZNZuF6UvEfVAfi01ti7I7veDQBtVCyb6iJEFt4QW
5O5eTqTOlMWKK60TUPuaG5bjNBP9UASp+V1mkyu5A1TmcHf0lMmGtUuKzX4g
l9TrSYAxC8Mb9bEgvkiGr2deE8Lf6U9V4z56nd06Eyj8BuIEZC0vQTVkOXap
KEotoO5fhlbD+G4chbnxPRzTGC9DaNnmgnPOpDD51IL9X1ieyUWX2kGNJU1/
UV/druoWcvOMi4uKDfb4Ysz7W1EvUiAyAEqSTScNjbx4jzwxn9MTmv2LMBVC
ibC0dT0mN+CnoJd0Z6MwPeN69xMP95wsjhswbSfUcy0WFTi59C5WRPKv0Lkk
zvT3whrlAxEMGyVoFkIlPtixE1rwmSkVCFL+A48oc2nYW5yr7CN/P+B7muAZ
+m7PxZ2CnNbsGskvveOJ6zvUSKSi3Gzklrcagp4uWOQFmCl3rreypICzDoLg
vb7QRsmvmlfdkEvHGrtVkwzbrwfD7hTz/k6DsPafv2q0sj8pBYHIKEC8srIh
Jgto2QhEsj1lY7EIrANFTqYMYbyD/4ln3Ha3yWSRSsxtEM7BhUjmPV82WRtv
EkR0WqheLgNKimrNAI2TNBNM5bdom1P8rfXqJEJOl7CGVa8nv5i7JZ93yl/f
D/jrQxkhjyhfzCi0gI9T+G7PdVBHAAhEc3dIu0VzA00KynM3xX2V27fu+PGw
5CsAwx/YrDWptEeztbWvv0t2p4RpPk9k+k2zuFprNpb3hT1tmFW/5C1++jrZ
q2u/HmPsS1I4sazO8Xrm2AQ3sMSkhjD6KKpE7g3J3a4mXK2uovpttOomQfbY
cVCb339EonfVk6INnfw1k2snldwqJTv42HQ32QSZt8cOjcW+GamnKkmXETo+
wW5rGQ5dBopzxBOz8uZqP+8pFssSlvo9ImKRtCsYjmjAVc9KFaZmArBoeiBS
PfTrV96mL4ha62Vq7vxomMRUeUxNHTe1VgCW5HNpUjI2zU0HiOE7VEdqFFaj
oa7et+9JlxyZ4hddT5iM0z4NK7jD/2FR0TaoV9c6b6zF7OmqW3EeTjFEoQY/
2k5ar0mudf2B/fFDo3O97ZVuucNu8hCG1EZWv1tKQG2I68rk3UmZDrpYlO3p
M9sLRQR3tFD8R006qpP5Y9AnQhjT76aAHLvk71cKOsIA77kKR7D9ZgVyWYWa
Q9YyWxZFWI5Wg6rNRadyGLEzU+jAurbaSPu4fYzHT6EWBubvUuMfxX2LM0NO
8P8IyjyIYPVw7uj4RXYYg1woZc/0Pmdc66dIY5dEQBXZSQcLB0c6Pym+Hw9q
whmpx9qx7ra7fKOgDNeCKAMnJW/rAO5Rnm7Q0eAY3N3gPZzpNOpkjze1p16o
vLlTgqApucLUfESCYVn0TUksk5CMiYHzEdC0MOpHZy6ObvM7kV1qTAZidDdd
rgfZ8V27C6fPlVFnsLq5INetDPpkPPPwnls9UqPz1vYAvPorIV0zJk5teGD7
3Qk2l+VvLmsbwDx73pJxWDw/LcHZ/fBKVzWpa785BoCgamdmYp47B1IKhhMl
4vQ3WxLBQgxDJ0bPOjvzIZfBTa6YUR9OMTVljMJVP1eLXZ73k2huyEOnQwuU
kkaCIYeYikHTOKLH1OtN1WAVFHuNxBNeMF4NkuTyE7JUJqFD3EgnLR+Nbp/n
L51WRHVQ2mfGMda5QmoqKRoJzcgv5FMTSMswE90rmrrEvahKnlvsjclZmHTK
P14pDia/nbBswoZfBTComsRkAAhrae5pyqx/8V78tdmJnvLU5D5+phsxv3Ay
kAKYuhQP3H0Jq4/UHxh2KjitMFoPoS1vja+Kc42Qnkleg6xXmLcEaKNVnlBR
ajvMxDMIDUxMF26T4Vz7dmTxT3nm3QCGm96X52Vqk9L18g0XedxKkWyqUT99
oujdNFakP6VfW/VozBBQ9vaIm4kxW8OoFbrOgVUXhoGH8LXv2WDOAZg6P2nk
Vx7FbYKRCSi2iPS+ZWfwjeq7obODbtkKFk3Bq+z8bHlB52gcTgv7YFyMApYP
GSvzTF81/mqJDDyTfuE8fGl6E+f4c5Yh4wB3sDSMhW6ieR3bwqRQGmGIzMPN
DbbyINDRkpyWEQ+fg1uJPAbbkoD7rhFo9WeDP3Cof6g2u9qJIf7R7A4SOJi2
c4PeclK12lHAPePq5oRq5G92JqGSlOpvTH7ZqxSlaf51DQqAjJV7hEu4H9Jv
+AxQ5X/nXWuXzePCtaqFdCyA0mWoL/+HCbtgQVElVmluDjFKc4lncQxdoM+g
231Q50wjsHIj70G03PqBG1ebcmmlkvZXPWxCft1zAxRKdXe9gOR1tlOKxjFw
QY7WyEDaPjOB2Xxgjd0vyFpKwmkO9qiSSvjUgI6p8EWVQLG8D1PfG68h6s9E
m+KXy3fFwTdmQPcKOuHsfHzfraACZdRhGGOI8wdl5+mpjRm/7lXJ+AL5cSC2
og/NMz1/DZfvZTTriBQlUWJesXPkq5dLAMV6/NVY+qu1KM0OO1lArMgKsycn
fpldjkt3itjHXjihdbjf9grnrduyEKod5CDXip9VDWxJPjC+uETlGPYQGDSg
wL3NHH2J3Rl0/+FdtJV5u71q6X4YrgXNXfyqOAbpJu8NYDACtpyuXn9NvexD
9797J/WeRzQspl9zB7SKc+lAQlXcqLWkad4QQOemdrQFTuhhB3rBw2FS1G4C
zk+ujQcTQyVwr73vWuhVEqpjjm4ER83GQG0guZj9Nb22LiOPcaJdc4whNzmT
ISY7mMqSQXQylPvXcpWaQpdWFh1HWJWf8C3t1yBYllhD/Hn3OxDXiTPO6nT4
F0vZSaWiq4Q5MIKEfQuvJa2B7dawbtgria+nZxmGZ9ZPg1kYr8v0qAg/B49t
0YEt3geYvlVOmcAbUDmPv98F4tYVRBiAuVct2fI3N3cmbsq+l2MFQv2NFTUH
AfaSN9iv7anUkmL+2Nr+viY52ZUK/uENzbWZVmEZF/+ZoNn8kTSH1VXNB79w
vDa5WrnGS5A5e6kFbYscWepgCLERWHKqWLgiX3ERfnt+eH3KgRzJWuyRoKVQ
jGXXX/t0JogVoVzKBtku9Xkzvxard4Ru7aRhoQgpC0Pf2CN5kfLedoLUzhLZ
Ovx3p3Jt/x3RHZghLRvGDSJ/YuyLyNsvsL3Ok0rgkQyxlI6Okk3e7kAFg/BQ
LdjO44DcaqQoD/or0i6gG30n/AIebdYNk/RCJIGkNW9lWhb7HmhCpMFSo8hY
yd+r31wB8o9ChK4+iv1ViVoZrmUIgZDEkc41l1SG/HY3MVNuSl6Wxon1AwCt
D5XLbSvLpeUo92pifBOwa3XmKTSA8unW7uCwbAIE8p2n5kMNGiCUiFdmOxLb
Mvyd3nL0e+FPBjqTZIHR7/BJSU3ycacHXpi72HF3kDd5hFIJA91bOaAfsj09
mskXyTlTRbWX26Yinqn6JDRgJ3Vn94mMOxuoFcCitGdbxdQ2xnZfubO0a2Ag
XC2rApuILJnwP6RcBYyv7MaTY6XmoIJR370JPuBEgaCboHNbDTJfMHfsrESQ
UKNicKYfhWNA4UzhPOxB8Xjt3FmR/N8OI+aRV0VlmSBRK3YdktCGv/Lqh0Af
jW+F/1RxAbv5Ptx/aQuhgLkFXPXBLyT+YFrv/NZN1HE+VFkCbzo8hObB4XFg
bo6YvsR4a4xJxnGz74RoJKjIIIoe34mj1esXYoD8bL8e/MZcsxPGqsiy5cPX
RAyWJOEOoiJW2TvHjea74qxclxiy2i8Dt77UoDwW1CQeQfkvwLNxS56I3inA
5O+xkUg2rjMs8V4XTl/a0rI0ZyzOUJrZqtLp0L6WCzvUbHU7j3wyYrI5VxRL
IimsT3msf9Tmv8ITIRgzRj+RhRToolrwMNEXXBNgGWWG00V08uY5uoI18l5A
U6ubYE0lncxzABVkiLSpbj0/qOZf3grQnaojMHm2gEf/23k/XX0eyt2JDBQi
E8Qu5iEKWOcUIDskfs6VmE6kPa0Dxr7UkawdA9QPj3GbAvjka3gV9BD8wOtC
+EZ8z8gRFY8AzmkZZv2KtfL2UT2xvMwV2Sax9GvCT4uSpnzVLcRWlLi36ATh
iuiH8JhPtwCou7jTi6TuuLmLBs/jpfNTqlp5s60uSLohJOP9JaxZs4Bjdwdv
LNhTLANVbMKngWbD44Eq+8dHgsa6EBkPnyis0Ajb2kfgFWhazes2/FBv8l1E
/SpghP57y2t808j7GTALYycTrQnp9Jsy+5PU5eQYH018BDIdPNQ+zUajvfeq
93K5vBnvliTZOECwaPRU5I8FiKUy6Gh2gJOC4q02Ep+KtlkWlWLAsnxb46Up
wHLd2WDA7kSK7icfjwWF1q/+8sX2eRtWc9n+V4DYWc6ZDi0PFU6TVBDLy5TH
nIux/+FBEaGfjCrRWq3vxU7YOHWGdvMhGrcGbDSxVYsuGZNMeURAlH0tv26J
eQqGyJ24AZmjGwkxpJtdcFaOIuYLlEn4nDrq710ktBTwjFizj0ea4lAdoSoL
qZ5WmeAcaEBjGMd2aPEP3arUpgfi3A1J4Gs9gTwhtpUT2bgqgYrZUzw9z6UV
C0XviW2NTiajTtqBQC4CHaKK9hrAUe5dLNDIBI2bZDkSMDpJJYiew/S2Mu4O
c1HTL/haDRiX7XnK7FBsWd3VC957YZb4Vq/Xxgh5+NVX9LLd2bmTATeOeiLn
WuxLFOvnKKGE4zKWOFrrpaaUr77GXI1eDvz9ZwQsUNw3VtRjNGrICtnW/KET
n9sd+dJNHzXsnzw33dQa1UQzWPI6D2fVb9sYoHT6wyRG0E373kUg6vtB6/nu
aBvjPOaSI+WUWVgPQ8EypKQNYmBDFKMAVdWCFQosYG7iPTyJwVmBktpaDjT+
vae5NYzUqtnUYznUU/OBQIaL0iYySHiVeVDrMe5y/8tsDKYpWoihfhQvl7Jo
LwqnSfpouBcyTD1TQUKYKIYC14knkei7rswyn5PTsJZWQm0nc03RllryztoE
VHURWayQP+uF2qiDJT83762t76YVgvGtRfUtRWtBwiRxpju61zQE3bL47o5j
hDyhjIzllCbrr5dDlq3Ugr2MmaMTuc/85m7K5p5cngrp6Rhm0ZRHoVVmpLit
NMq81zYdAwmuCjrctriJ9ZR9m4TT1UuFwB2xePkj/ZNTVlKgRb3SY7cl7p9O
vkNaTmf5zITHcnhmuL6v0XkD1WpoTQN3xX+sJi0MUQzEqrquRlb489fCOU8p
GCwfp4PldFk22Bhz/Frqj1O+5mjQpAOUqEj6FHI2HsGAglRSuEhrS7G5WjaE
BC+cokJphJhrkD+T2UhsQVORBp0GDu8PHhSstHysqTMOApirHwkTyMT8Xd8i
wyuKVwz8TWxK7eQbxourdYBt/jxOK7e5+nMHc1CMDZhmLPu6+4XgqPeccLe7
rIxuEPjPld2C7Q9ZYtffXGHHOloIBoeI1TrrM4u2svi45YwQPgokf/dJTbQF
vuyuhYg+0h1GNKAU0XhxYxr+xr6J9fnlrhBff+GyCQ/V43xF+c1pMfNWoGBI
q7m9xfDRAKx8wz/cewEppuIjVlqMH3wumH9mMYWZbNGtQr5Iz69nW9bVDiRI
mx+rlfcehLLb9uD7yIF+SOGBjQJzXSeZCWO5YKg4QNk9XPXMXJYrLCkFUYdE
AgTuGfh3x5bXSRJFyQ+dpCPrOhh4nVde38NVuD3B11IcfwLwDRZHcKUOtkth
8RNOXp/jeteMaCA764B2Z8Zv9C4W1NKEkwMI6UAR37w8GBOiRQSwsxMJp9kq
khgqdI/VkEow/bj3Q1mBbFtHCVfXrEmxuFZrrW8RiZLhIQj6w5UOyjo3HqQn
ulZkbELG44vyAE7pGG124hbVX4FXGJ7XyHp7AESpvpVem5B0n8qtfj5K2fkx
H7bW4lKcuznls0I2dkObY1UhYnSgWy1ALbr7jxRkhNRfMT9xvlhnxHX0rfBx
b+42694oF5kHjCTOx16+Hxxe5BAk2yiuqUYiGSWS13BfHaREdAPB+ak77KmF
Kd0nRoF1pa6rnXx7pBEmOP//YmqIkP7EL3Q1VJc7/x8oM4RGvDfeTUHTS6Ex
61bzziQ8HknVYjpwYrzRby2WRSQ3xe1p5zCfWLc3jIOpN3FjDZThIa3RTkKZ
QJqf1n8p6sqn0q4+VXEMs5CM8u94I7K98Zjf/8WdMzJssJhx6zhNTOAEjq58
TPIFScPGG4zV2Uy5H9hKCcMnxsqwL5yk+h21VmqnOCzfpKDuDeOS+OWE0Gzx
3QfZJFSbqzEyqa21v6COd8RogGNt5Z2XqdWac/Pbc+Hk8D3ZbqBAKCmyzGuL
lklzjvfHUmKPjkIEMaa5Ze7XBE6TzUl+7qyY6+sV1z6rKmOkSYHj6owYXiDR
/eyrhyJhllIJ8il7Q3zYFbJSbC3ej/AaudnlU91gX+Zld5UM3+UYSxfDDsyc
0Vch7eO5SRAXEunBxcSxziQGLWkjU3VVMXl8BYVaxk3GdC0nLqyAGCDiJz6j
xYU5F2D4aviFG568+i7Kbvid5Ojaiq/NJ8oslydmcAYE3OP1cosLxZjV0XYD
O7Vh17vf6Gf8AD9hyEySlXP5WxcroFwokuEvq+O3IwVztLwrbgoGj/jaFLcT
ZJawuvL2Nk5j93Ttp7oCK47zVpoVfONPwXg3x9jxMnvEnLCNP+lzvdypidij
BSnsY8a3HS9Mb1JJidRj16L5xqeKVq5STT2weyrSG8cH6v33iIGzkfO8ZNKV
Ds7epFMPmfeChw7iTRvDWaQpm6briS13bD3atKPb68CHeIWcmmfE2JG8Tl1l
Pz95EzrXdGyD0NA2qi2aQKquBLxkdI66LJMbhn/B7eTzleS88VmdB9yY4eBw
x6s23Q8JPN+kZXov6Z8cQMTSYIICFIUzr5N0NJz9w8s/8eqsJenwRra/mVh9
CEr3OpYeKcUW6KC0T1rSt6HcK02W6+zkCUOU1SFFmQdJ2RI8pAStU/9766kR
8TpZZXAR5n4UiUo510LNdXPDv2KnfudRHzC09SqXxpL0vqVj9tzUd2ouY6lo
iy8b5L6LemWE1zg6H6taXwbpl5bw+HRAjwTPohiYqCqx+tthhsNI21TTNmci
WX/kvvcK8VW8LWh2+Xqo8UcObM1/ZqRmdSu6CMRccxqldiHcP7xP/jAqLU6J
kQ4rjh3Qn3u5pT7o7W5kWoZ3/5Tih0QXZspe0JCP9LpwAfUipgff0CJ5q1hk
Ef5VVKcqRCM3X/crSvZdF3spFLCU+ysAbDjvhMvnlHIlia4GvK4rKZCcIVVb
GcZgqCQ9WzJmbHE0pZ056cfjZY1fU+pT69yA/fEaoi8mAZsItbCBm36lVoRJ
t+/uwJpO4QEJqnKaWUSU54P0X0K89EA43G6rO8wPvkNHaiJel7upuHwGRjU2
3XSBr50a06C1RkpmdsXWaOONBOViegal9Pa1XytZ/T2CUQqUfIAcwvMqvMae
U3aPyAPcJwAvoJFIkUuhX5MjTWFPRv1pNj6F1a06Pv3bCOtDj9SCA0WPfeBA
J9OHRUTnos78EcTU57IDB2TLD9TO6EvhAoljaiyrY/8aQiy0B1cccF2+kbDL
j1XmFKgAX8vV+50pTBT2h61By6Bl0FuwCMvGY05TlTR4Xw2FxU8FqzB8vf1a
rY0WWfIe85B04Bo2MwNvx9cJvYvF5r6mQKGHZciInL76+bHcDNgcAvt7hU8U
X/wIap9lA57qOl4/jXTuqIG3bhrR7eLIdkE6bhAmeMnJNLoIBjeVCfy5D54R
/xBf59YJu8fTvWqXh3yDVCu4kk5lbHpgIfGTyZ3rDVMPaHtFzf/shayBJ0Zm
ohFE+ZzZqi6D5L2csajKfKH5rjq7LRiLeAOVTr32pUVOAgBjSrH5pmXfVtD5
XpLgLQqrff5dcervlT0OkSyM3sZpRExqrMDZP5b54lWsFRfW9yit1mSYT5ig
G/TOBpsB6CPx8Gg9k9iKmGCEsDT8rg0CnfwirsxUkiy2fbxb2jFYXGz1EUah
wkmHUxptEojBAO7rgUYeXrbLovH2KNr+/2zPAgxHFZltgO9Q50sUHECRI/4Y
sImWEE91zjwlYXPdLf2b3rfkl69n0BUyEb3YFX+gO6eEDdpi+T4q0mXAqeJ8
IuTU7CAH9c4PGk+H5wUZucILKJzoa5JYaoOOWQC9Ohj6Dp2P9SsS+cRqLI7Y
rT9/B8JConJ41dFsSlGRSj5FrzfScNpUcoRmzdL5cxJ/4nA9vgUOjJFSDPjl
gRChQkGpKvYSXVjsJGpe3m41jFB6VUxqQIjXmQqkqDTcHCXXB18LDwVHlu9L
4wU6hKjNSqPDQ6ls1YkTGkvNMefGWWZDNF4Y+clFHOZtrugA+kjIrMHyNJe6
ygRIcrF1BcEwlz8M3YBqGN5LxoSIxCF1gBwt0fiVc+AwfCLVEeqjzxhpa2bR
flE8y+OdxEciLoHOOI9zm9Pls9bn6kvFneZEoUkMhDDQ4Mr2rXUt2X3SZmqm
B7gfnHaUQekRjjP9x/ef7YErWOEjof9rbFtVdbSYlAAtyzB4Wdk+cUBslJJU
FIqVrxbJpa7lWQg3B4ZqYraav4GhVhhUeA11E+ksWxvZDDfJrmQtkC5cDJVS
fvqQg8ro/GGnpWHIl/KDon3T0ftT5HamlCJ6FaMmW8hsMkX18y5Aqns7hLJv
pgyp5OphNnCN/G1QzIt9mw4MioLSFmoiipPi2sVzDOU2PNP1QUiwMRdMR+Dv
QIF/IVTv9BO7GJOSYL5hXuthrir3GaRpuidwUXfOiKccRjrJ5QIJihMJme1g
XMWuGvBIER/rq9C4bH+sdJpj7T2WKCEr3aCsV5dqoX3njx9UUJ4FC1Bk0t/v
3K9G0jw3DGaNVgcep1e8iLzf7Cu8CLSvKHRqqie9sJ/WBag5oIYT4thbrql5
AVGbvQgkCVsndUlIG4LLfParmxAmR7/uW70EGpNkhWwTHtMSMgYW2Z+hFHfW
yvxTFAAS5prKqvuuIIiqt+LDBuY8I+OkjznQ/CpAOYRQS5jbTJbXF1/V/uej
0EUpq/fOMu8R0mg55ZX3F/yxB/HPTojPu99RmoutB/hcVgU2ue7L2plOdnOO
2U9UkoBKTK83J/VcM1rxLaDjGeTVGnoAXsxzZJuXieOpXlh6w/ose9/JYWFf
MsU7ibhQ5aJciqH9gwx0gZOGF037XEHg8DjF83Znpz5CTBuv+6TTM8NZlbAr
pdiqEc6+8/kW+2DvVcicLT0vZVVslESlqhPJSKgiAJ0HTPplh/gEqi8dyco2
/QMPQ8bCsKSmWbL4ndeef8MxWSG+Bv+HU4LWDYdjqQkOaEGMQGEW0hNk1wIn
rArktS/yY4OJ45To6+lYX5J3EV3CA0/oqtSFmlSR1I8FSxMVAofgmN/bvtJq
QGBn6c9ljrk5AFzCiD4IA3pGIsZU0vhIejmLRMBwbh93crAEqaIJ+pyvzD4/
tTmNvxIULu97GmnxQUPj9eTu7SgoEHwuNyGM9W6ETiM3VK0x5ZRI2ZYVXJU/
KVufLaZtR91DOPFTibLYLEehLt3g43MdvOjYArIKGsj8YJvwtlfmAefaFhlF
XJZCpFnej3i3P31/UXonBLf4+1ATeCMaWsZFvF+snSWPmsUBEWl3wHn4TMMj
lsu3KtnOOa0ffjq9HT7BzSCz6Khn0VnewxCvmjcD2ywtkR7NL72zXqGCOfqg
876mvXp+/Dqb93vo5PDF4PczUQMm7ssbO2rMPlhw1hCodVawYBF4tyx/PN8r
omqbdLIzjcuelxpjtjdjzAWtZB5Ny/V5ufk9O3+alqg0VghIYIWxGMSPHNiK
OrFeBeXMeKFrjlUR5Vnwpsc5s/uO+jgmsEwrnFIgzaBKDicqvaKnXuokX+Pb
MfCuuuY4oJ4jJ53XcKLHhfbW1VRuNkgEyMwJqkFvArp9LNkBl3G59UwczJ9Q
jf0Q4YmcfRE9mTtkKbeyv884Ldq/EUBAZLs5rfvk64l6gMsT5rmEROqmzLcs
TFI73Ah/cj1RIgbqeBRTPFZrKVvZ+NCHVooGX6yxFjctrta/lCVXBiYuK10g
u+HW0YT521zXniui6wgJHiqCCdC6iFZbpIJEEWgPPXXohdcxu5c+kc2wMCZR
OayZdvKhdJLP96VINn6I4ClrpJbM7P9prnqWw2CthWeWxl+gDyfbn8cEe/0K
OtfW4ahdgjDHCHgwF6SaRvyArDASSCBNwCbIU1zpPms5uKxrgtv+RwdmwsMR
nXmaU1O0cP+a56jqIi8WOZejodXIA3zZwpK4xMtQAMORja8HyVtsutEMULS5
lZBatSZ61kH83O1x7n+gMW0UUmd8yVE3h0Jgn3lyAmmm1eaOmYNQnvqAlGYR
xsql4XyJ198t6vMdz9L3Ib3l+Dx9lCD+cUKfec4yCTa//QIrPYG4Md7qQxx2
8bHZuoXbVZCcjzpEBI2b76sg2YgTbaosODPf1yxJzBy7mPq3e5wSJiSYb27O
ntRkP+ezSQdCfgQfxq5wBHCZGpDaIrY98sSLZ0xyMe6SqNVihptA94zgVJLU
en3KA+elH33h7LjT65Zo2XeLtvAAuSAgjtfaAnqApgCL08PkImjJ1+IhuVl7
mzEWPhJ24hczRWivvgF3cB2fRoeKNE4X6M8LJbe0qUSfXovahZ0AAH5aT3XK
Ti3/PhYlVFnFjETHWxaiP+yLzf+5UPjbEjNfWtYED92VYh3OukJnFNnBri97
TY/QQuVKu+olLMxO/InKno0bKVpSBu9ejBKWlV8MB52MiVSrl6ezzhiMYQxB
qeTuStBqgFGIKH/qnx/M+jhl4kUch7Dp4ePjR1r4Pq4gPGAJT2xywPz9Pw/Z
JcCmO94kC6Ci5gJU2DiiqfAIGOG4C9FtnkF2YGmKW6wodWTfcTCBBBglDFy3
zNO5u5Mij1DWrx/A0eDslkkHT3s/7D3pVR2S6//msBzO9JJd4ZmNWyQzaq7x
SSPBYltSrXlFlpTuF87aShbRxGhC1g32VIigCGsKM1wsF9HQjGiuboydWfdT
OdjDrr5y8cjpBR7/2tti0ZJD8a4NOLaPSZVaoTMN5H0aZN5H6eQk9rf2Zq4t
+6Wl6Vs2x0EVSGEsSfuwyHH5lJFfY6HuXfTjwu4ou3Mi9c8w0fEykj2t7+lJ
Og1ZB7RmzbS3c0xARfcA5t+Jp+fB6JAbGGrnVENqb1MfsWYyfPZGF6Q5aoWp
KGldo3n3bJgJMR3vZMocpYMFXFjdRQrUrtqDdfrfjtrQlRzJSYoLjVI2pDE2
qrmDACOcpt1dZrYiK6LcX4RrD+HFcbnKp0JDdspjXwPVdHmEyLTRkmrHEBBk
e5Bjk81YULxRUhju2zPh11crfzBZL1fR7Xmir0CNHA9S7FzgxnxONqJpv2fr
J1gHlO6zHP6cWkfs6u12gr63zLhPFJV0IyNYNQamL0X55kE+s2JZyVSDEa7d
TspMiciISUENEpv1ar9UwMq75+cGr2LTA7RBD58ZmbgD5lAoHF1U9aoEzA+V
DZOeKR0hOIh8FqHZ0RmTuVs//j7WnxydjCxDj/+DSQYpspLkZ7XJSL4gtlzn
BZWL9+7S8YjfAgMsAIBWu2unPYXi6licUJu+k/8GgKnbRlFwufbUaCDf1mXD
9Pa3ziW32XplOhN36t75Vs0Ke3l/PlbVkJF+C8uwuNvTNjqKOT0dVg4fO/rw
MDLZ4fvU7W8iWDzG6QJe3QrYXj6Oie8o8yuYqi/91KE47eanpxoWEejNsV+7
uYDWK7daS0lABNyJfPRXcstZQZGDEyHAhwboqTZun/kLfwuTSqwcMVHSNnEY
mj+4sJ+SVxPH3WE0Q6FBfTBcNAqDomKc0jJ/aellMoEnPJoAJWKohaW9gYmd
X+Oqfp7ml7AsI5JXoHWILC+6BuNTnRK2VQ8r/RW7eYSJ3+vYm4UCe9jhB+HJ
Uiq1Dqn2mzNQXwX5PsIcXohZrl9nMuXHu6rJpex3vs9rwdLP4u5StEE75Ws/
bOq3GuZ4IP4Ehrgl8JcqunWDgnCQTOmQZMAUPHh/My+uIKKq9Dqu4Z90t3zW
p6P7UQXtIpCka7ZLKziuO8D4o2uinXz2QNZqSYUvc5QmCq+3fgC56hiWvK1m
Vw1j7h01XWO7QXZVqdsRlr8P39/EprnIk1SadEGfIJMTS1S9hRN7j1A35YxB
XqoFmvWCQECSQrCiLV/BGbwF0OgyQsdh+CMbIUCkKXb3Pz7PUEbAyYqH5nQj
hhLElu1b7lpyxmFmUY3Yl2QBRCH3JtUWBC04domkmUJPqXb2h1mopGDkOOfO
1eHvDuzZdeBi0hFDEHaLJmKuI+gUV25tNhQ+ZP3mzHdwsQMTpBUjVIInTX3H
r6IJ5XDzs5OSuAJvtkVZGrW05jHZasCXThkl4aXMpoyW2Cf3uNKNLvSiWAG+
3IiJ1IncZnatxDAsmMSG3S4x7z/HwCrEP/NspF57O2FMmmGy3uun1+hY0xgl
K0S/gRJsWGz5EK1wPAwYkRY+lCIzg5E1+If+AtOeHGOjgp8VimdCLZfJ5eLF
TGd5OwaoIYqpD7TlCt6B10Q3kcmThhwCnw67AN3gNsFYaUmVvUpH49kG0ePM
LdBAMxq2Q5gL1Sl4llEasVnF6qnaDhC3eIS/DWiodGHeCnJK7w1MSvVs2q8R
rH7mpu39Sg34zdcqV/yRxsaddn5TEFDnvhOqjS/4N3Aa2iWdnM75wWPKzmLo
g7RK00Li0NxgcfzmQ6W6p4ATaGs04eNaJrsIXA9RnRsse8N8cWc0Tiiq+C8K
aGQbpppxsM3+QMOsTlb2c5rMrQvf6AvDF2/atQWAsp7yWmBb480FfJNsisg9
XQIu9vlH3KlY+jZ0Wf5fly5Pp9tZG7Z4vmvXiteRViiQmkFRtx0jEbFAO/K4
TjneWLrq1IDRVQokTVMw5at6G6lWfQYoigMVMf7ek860Do5rcZo4jjL2PLce
fUAUyqkHBb9Li3aAzuQcZ/i2OvwQ4Pdzm9f+0VIQcAfNt4f27XNEG1K8fPFW
mflBLaz5dzPE21LTOQcP82fKyQ/k74eq/R79YM0u9YlDRpUb+/jjL8W9Juyq
kAgpC4ONucGePQWUBgi3wOQbjRI9ZnGddnMHCHAb2eWE+Vs148uQRCAvekRN
kXc3zRaVf2UikO7ultaEP5QMxmOh9cv0JFCSIJMx/FBcaoD4/qPBCEY1DJTg
9B8KyGn01UxxtGHFVtA59H0FaXhtIL6RiWuSlgLJhdK5DGb+91m68W+URb4Z
NR4uTd/WkmiSXeRPpwmsFkk2IVCKt4f9ONWSQGO17NVDWidl5FVhfFZvdAK7
cfQL0Ccm5qsJsqOaOI9F2J7jHHDyg6hDUKuVE21HRz9xd3x3VgLhe00C111U
I9W6lQUiPQAZ0yl5aKhNKLzPrWI7H20rsdKG4868evSwp6oiobd9bRZoAKjU
K47Cf9lcf/iFf4ZTzUfRmXKorOpHZzccpciGX9e9gnh8UPlYUulmq0UGPPUT
sISpBTu8B6Mg45bHj/+KlbVII2liXwuCbnQu1mFqJMzE6ZXAAWx7CnIaQbRT
vMGdr16nenlWBvvOCm2StsPWwuIUM1otBAlB6wLtUP7d1S1HfGV9p3f56gvi
E5meYOnsV/JiO4fJcdSNhzTYCZd8r8WfnVytAQkpKjVpk1KNVLSpiFiFY2sS
DX9dYArmIHAAV/whgq9fJLBrSudNwKX8pJaiyZP0182bnRpDNURrwJTy3fwn
HLmc71lboRHcCyJX03Ye6F9B/5S4UVUfBi9ReVU3oHpp4//Khzd9MBDbXkOI
Njwj9VtX/SLpYE5heRmAHcZz1+3YPNpsHsG8LL3kWRNOonqE8uuyWLzyLu/c
EjLfYlOdX10CSn8UP8tQMQlVmJKeVaIIoqU0Fid84lWE2ZyeBF68oQkyhlFf
q+shkRz7FIrfcf37iF4ufW+Q7Y49WcrwFWaUQHHet2pn/STIek2cIGA7xF0q
T0JV6W4jdnBlft/eN2+ZPei4vSMRApuwPWKv3LBECuI4qd6ds1eUGsVLEAV2
k/fNNxNyA7ufaZphvzuSYAuMyXhmbOXwtSRUThC98IjuSgJhNOwArIP2Sk91
1Ulc+vgJEd/YtNA1kuXkn3yVMqlQ4AyAjvWM7cCqIZR5T/kljnKLhZM9DE51
nCGHEGv9XLLVuohKhgEEjzq+25TOLYM/MmC4ZGmubh4SHBqahtkyM4Mqvu0M
LvC/XiByx/iTRxdLxkNoahoHOANxQ+QO7HwtACXSUO3MSt1jpdBmWbd2BSbj
vAQNSH3KdXQMqD/SRNiU5zl6vyuKEsaQEVebF9CEQso0mX0Er08lRGPUotyt
ksf95UFIRV6H6V27cnj5Tf4zKWgenB9FhP9kxRhtNxtfe3ghoVErfI0RshRJ
7l/WZ2FF80tZn/1RClkS7m3fSD8+Tvtu7B0DC66I1M/dOJD54P0gQM47rAeY
BK48abU/NcN9EJC/xRiQsr0YftD6EGE7SQyFxrzvNAfqB54Z7Z8b8jFXXVe+
H0xgS8LNez0zQdP4FpjERb6lZbGnvc9dXNpeezSHgpyoj7GMp7vNCKLYzFPK
UmVVhfaFKRXWSXbn8a6tkpbNI/b6sOQRixL8I3qcgNmH+oHWpFVTP1HnI3/E
gaYfV46NrP9E8JC9WSf+wlTl33PhzUP9hn0ujR4Gfd0hxcQ9iTAd1gy3Z+62
B9z3a1tB1g+y1BMr+UtP5Say+H/WmrL5jImcsRCrRZVCw8mrXRChmbWgE7Ta
8fxvDL5gO9H/NuO2FxVJ1t3lZ1LbK15USmVzpkn0l+TdTY63r4WnHMVuF7SD
T23fqToMwmJ9FH+MyeQSP2BgU2Y9+pQMmp4DpF71hQzytsLEq462VCtKSsbI
5tygOhtjc9X77s7elzmQSGufDvgv3R+cpJLwlxbsf9MkVo5mAFqD4vhsW+yL
GJgQwBfd5yq0l9aqN31m5XaSAJ6icZkRfxFCqIM/RjE/JrTXXLIAtKC6i7BT
2kWFQ9DHOS+W34rM9cdv3QtQNX7IfZIkkfMamygsDwbsU+BAguEnyvN2BYLa
pJGhLsvnQPhJtpnYjia9A30vMcK5bDWYN58XSGSP7gnghK0h3AgisNSkNGkh
2cUFwVYEJ0RiOEIuGjfCzn19Xih8o/ZXxqOXf+hD5C9g+3PHmBSJA8axbgn0
OMKT/km/bRxOHmy76YVe634v6hBsE2mh3EvPqA2XrppwslBiwPVDTtnAd1EA
MLsazj+8B9oshBaGygqhEQOkjrj040kZ/DwKKKYwhoniWI3tlbWJcLNm7lBO
fpFsFF9QuyzR5wZmdAeR00jmyxV9t+NRlEMhl1N50lPBfmT3RVCem6bfj0Sy
rdfdQf5j3RelQ9LskUwftWXyxM75BltwrLcIapRM1JGd3HcCjiKGD2ne8sxr
yptApOjAR4F2qp0GeIxmJjE6Yi371fGzPVAq0wojUjYCbMoz5DOz037t16lR
0B1qP6/t5r/rdIgn17NXfgyI1AMTYwmrFBO348Qw8PhJym4QO4rjOeuaRPpY
c09cA7HzCUzxhZjCybPHwXlwna1vA7y33d8o6DlOZSNfYIVICIUvZWNyZGrd
LCyGLWzpaWqP/L+7N6L9dB+LgxXlXf2cr7NB063BvS4z/e4zdRH2sStJBe1Y
irK6ut8tGtBMLEyx32abpqBJXa3xtdXC7DSm6LuIvvjTVyVNhwmogUaJUEl3
PFKULueiV7OoPx+LdQeb9s/8c3f6p7tRv+A+6ba7zgDXQ9waLWeJ7a2nzU25
Ihcp/oAtWI9rc3YL5sNbXa85GgbQwTG/ENohZ4fvPqA0dOLalPq0/Nukte6S
+NVna+HfUW3bRBZO5K5OIc3arbQk8Jqc4AyInL3SfmygMefafbEEaF826NZL
DgsYY3QeFPIJ4LajJ+Va+ZDmqQu2d7ieX89JRrcN7FFcYh+DBCSkan9Wl4Vo
GsX4k/D1HNmm14PVfycPKc6ZGEHzZSxEAHpnn4guJs/Xj39+QaEGcSQTmv6F
6JtBxc5aYTxHpm32mrPq8CIfRbgiyQBGcE+yaeNWZiZe4f8G9kLhrliY35NG
E3564hXX8JztIL9jlxJaGtCssKqKqOdo4YDisV/doxb35jHF2wRh4pOTFTk7
QkxkWnUFeLpAtHoEQL+h7rAnPnEMKpCDKNUppVWzf9vP4FY7+5sXwGQEvAdX
1k8eBVPOOUazIJP1dcm4XDkoEZ8RAPHjcY5mVj7YF6VJTSvlViv87oD6+G+b
MwEq8ex7eFag7aDfyk6KZQoFxNaSVtjgZTypQmtHAYt6Q1LGWCh1H6Qw/v+F
JnXZopZl1KDw7hHYUljHC5Izh5Bscdt9cYwVdkGnlI7Uk7qMUZvHjndGNQYp
3R2A2we2nklx2i5A+k4OOmE35v1578gnzmk+OJxAxy88gkfhjAm7SIGgsK3v
Fb6WioioC/5sk6nVmCM01ICqX8crKwftVV7drj+BYcQk9A7GiQ2Q8dRuWEcK
4/K40YGanPiNQeK9GgLjt3E1E5z4GcsL0/nAPB9Ci3SoGsoLQ9ki9Od3NZPC
+yZaQyKAL61tGeVGPDCiuz58jbVAK0VjCq1e8Gxaw/BvTcxobKd9AGJm989o
3JccYfWKzsCxOtQTrSXfQ6xlefk2g/mBy61p4Y0VgxT3SRvmGjgwDecKhcpb
ndLv6XOTUTdN2mAXyf8lMkruqFiB1rLti8hHu1tl8dbZbDJwpk4IkcuAIktJ
e9AsW3MX+1gvVUXP/3ELOst8sniENF2crq/jUVCaU18NcB8aFwPTIWO6jvms
tNIRNLCgnmNaGwsS0q6N0tej+1SzKBXUyx+boDYWKJnFjGO9ZwN7j2mHmcJc
VielWnHaPXg0lW0pL+eCVi+9ddjHFRdzpl6wl2kazqooqOu/60nLm9ZDJvcx
zYSuOVg2PZgD+NJnUuLdKrE7zCsLtGFFdlMZSmaA9KJo/7tUmPrNKj8zu/Jk
Nq0mqA0rN3WSZ53RVoeXrcwRYCWajqAttItVEabPtbxN46zC1RLV8cPFXfvk
E0iezhrtMZrtHbiWxrA/woCC0jvbBjBSQsOAg35PCycTm540HlAG+21wFPyy
KUvHccR4kqvKUGUGU12VSRV1dsnLxd/NZoNAgDB57ojfZe8WnY18rVqzHS++
tzlR5z6pHHd/bZ4cfrrtCza8LFJAVTeJuSyRoPWE4wJYgsL7yjX00QCYz3nH
TJblCdEb2UBPFiuwkQMWA5BniYtHHKIW9plU+usXGZ0PWCCtSc1EF1trCixD
IdXrAu772y3Pfd3D5XwZKIX2snL5qM1UB3JOO4+fXGNWwXlq7QzzIVWqokDp
LebkFaq8KxeH2Z8TrCgm+BUivPHUJy5IF561C+smm0/0v7GEwIwZ2mqic1sH
pX8IvvJixLJN611ReC2TEf6IxexwuV+sGvu11+4rcfboOsdG4hL9vBpZ9GOS
CPz1p2X3NlQbASacYIAcdyBtDhuGdmw7i8xbxO1OXloLqLvhabaZjfR/h+FB
FkhKlaE63Yzjx2Cj24eK/w59XJx/MPRPjm3HYVhaT+lU5o1E0JgvohBP8Lqa
SJ44dZU1EXiUolA/VhyzJ6gGFhL9LHMFsKtCvKbpe88un1P+pj6+Ezy0Rufv
vS2VZFc7fLzSnWyV4SsqA6y5/FsqmTHcBswp7hx7AlAVtBcZZ7mY6kI1huJH
PjUHSz0UJKjqY9Mt2x3zT2hMYMCCkkqo/butJ9Pvl3G8IuuCsl52drlj6Qbb
WRIV2o9ckrj6hPnexeUIobAJG6m7fQQBSkGxAeHB6OieB8RHzEIJgp+Br6Dw
2DGmvPOdRmuswscLm0sUPuDgrjADOPh/mYyb6t5QNylmkwHkjN+FTteBITHT
W744FDU7B9/OOcIsBGxbm3sky9qRd65SsYfC+hECP9gc91rB1H9k67sAKb9y
DAZXtooHUcxRKg5T0YmtOuVftkgNqhDGA9Ccjm0AGdhsk3KZ3xPdeC7Y2y/w
pK2w31mN3o2zZd1RsE1kQAjZKKfD6JB0druXndU6MsPYnYwKuEY+azaR94Dt
bqUcljyphhEjr7E16J8M95Zfc29KwyFfwLIV4EJ+P04hbwAbcE70mxmFIHJ3
IX6VTHxRG25fnGGqAGoQeCuDce1BRwXC9b4VoN+E1jrvb5yGClstaOEWDzcA
7Le2KhodTdKG446CM3WJQ8WL4Mp7Lc2DB1sQu7gQJtowcerqghgBRVF0jbBp
f6PNXG+8Js6CwoQOFz4gN9jBzWxpLz5mu4mjiZ+JdI1f6D/knH1N+nudOS3K
BApJInx2/NrZTkXlp2a0FtjnqkDG3cvk+flPaU3acuLOvBTvEgwS9rnusih7
O6xKwVczVbMcyVm1AVWYBF50jgLxegZfdVH5eVs6VBHOdmBMMSbsuzl8Kgr9
1HqwGklf7aCRA7QFx1PBpMRODh9xzGPuZaeygX5QGc8Y9Bp4vixNUTYM4fWC
KRlCQFweh0NPSzziimVxBhfQABS4zLOV+b81UcEkW8Nj+M652RJguAgKMLyV
uzxY7haNcuFIazT+qMyycH7ae2a5duCExlxEjy2Y+OHvjCPkurJg5gp+lw2t
FYjU5oBr5fm2FuAk/EmmMBsOkZEqPIoAgxZFb4oSQuoawb+IWlZ90rNKPyhT
Lsg0z+nsEvfEPomqJC1iS8gqoaT5k71GoKoe/a5+In+tHrLky7tEkiyiJSAi
a0yXuT+Tu16eNmL+NGb82/fZkrQch68Mk5p85hW796Ot5vz9a/BW2P0pGekS
Lhs2T+VAVifqgtvFG5V24yHKkMZIwI9e6B0DMu7RGiNEJUbD0J0bIrmG5RTi
CGQimcmjs5LvJP0rCZw+zwM1zg2YRjZ2HhexLwyD+9UufM1kgicFMDQ0MxF1
uRq636yeoyCvRY4d0xA0tZemtqsew34aRUaHrYU1WQu1a83vjUp73lmNj/ij
eWuiameajB9Li/iQM3ujoR4nmQZzGO+eizw7LdTI2UOxFp+MiNhxd5IK3Ch1
zPDRrSJDEOfToqv+bjTK0iHAvU5hlrob+1QTgMPbRZ1bP9lLtUPp6KA1Uy6M
hTRgMsnjm4NtVDsPHhsBR8dGbnbTr23nYqkb0Ky91nV5W/a4VtPDI1Jw746Y
StwgPCnqtYBhetg4d/HDF2hrGj435lL8Rv3wO5EPBgZxLaw/NuFHSWd7P0BI
H3LTCT3LuB64yIUHPk242IV46wAlWtiA/KwXZC2OF2Bt4204qhxYCwUB2o3D
OVxtrmtRt29H8h2lWxBbH18IwRx0/Gf1df6ZH8luGJydLcCPhoIOJTI+wUWD
2k/bhuiugF55jov/HL8FzxAyV1cKz+TCUIVwJvh1O/98Fh4WAibtYZCraoIH
OqqNBnkDPZ2rJsxKUuEtbCqBDczCrkJPqae53k6SZGfIBcsJSlwpwKCS3ePX
VeQYXHjlF0uoLZ00wAc8OjfQqYzJIZr/jTEtquCDHcLuxEljSVIoe4cotIwZ
V/NexvgCDeB4Q6To21SOLsVZiVO2r9Xp6ZbcGYnoDmos3EXh2j0NfQRLxdng
Fppo98qBhtpG6qOo1mPc1KYPsVFbqqS0V6BEpOTwE1jm7SzlqiGmCsegVl28
dipGqVtDWq2JEzhxl4rBUsQgQYbymvWKbxiIw9tHr+myoG/jko2kTWjk4ovi
Y00VCox+xYsx7VzosIf6QWUuSxRjGCr6l8/6xuSII/ST3ViCn+sYKygrB01A
d+gKFnHztIlGBLNhabxBMQvCY/cJ8WdZs9S/myGz/UHNvlZHEepEN20hfJuH
LrB6Bsh0ogiE57BPEEzslkdcHOzoqp8uu6Guslif0GGwP0x0PKmu766LJgMo
+fn0eEir5bVpMjm6ezucvGHHYPwzQmqYJnBIQ0zttjN9KmBw9qp7Jpp5+TuI
ktjWT3G46PjE8ol1+bsJREFij5jt5BRbR9y5AKo7+CgRcO2EyVc8cDJK1tSu
523kzIf1kFHQe0BFxJ3e2jko3l0qwR+R/Sm7lFatz6uxvu5bQiZDK5Dc3D8O
txQbFx2+MzYned1NpY8uqNehLpzcU7zSfX5/J1tek7FwP5aIjsB5MPzWPZIj
eKHXkxi0zia8Y2LT2VDyOE8SSt6wQ1LY6fqpMF3bdMo4B7olAnrvJ7r646bd
G57vHK2dgy9rv38foXJJSqAyIe4pohpEIGI+WPXYNELiDD4mc29VqQFxse8S
3YHSyFUc4jNJsetzJ1OtphR+zAfcpTT67pyBE6ofV/6/Wevd6N2zQa0mVaFO
0aZ2ZZo4k+0tzHGgew23a5lNcc/kLG+kw8pHZIyJdKIQwUWXdYGTIfJQJZ8a
EKkitWBYV2cROdZqGg1tSrvSycJKHWerTbttA1Y2Igdx8fWVbZUybZ63lbyT
EwufgiHNto3wJI2itpkZUM0xOJrx6grkcm1WvMIUSQnNQmUGZIwzmZ8frZk9
yKYZ+CgH/vYGyNhhz5uuH39QWH5mCjsxszTbxu6DiriHXUHUzbYOYlyQtWO9
Ukeq2PLx+rLn/MhwS7FD6SgBmGA/zSIourOG68S6kO5K2a7QRoR11TH8C8jX
UkaQHlbkh6kJLif+z8sjBTJRiFpA9PUdXSnDB/f4p8LVcXuPGxQjIaOUfRo/
BN9yXG63TFScEP36KrrI8lVNSy1Waiipu176aDlT1n7xhkaiMVtaYis74pv4
1KM1DWkiSZf0PZouFP5zlLGFog2RbKyT2gdMoPioJDbJ5tlbE0/I+kNL1w4p
jE27tMPV5A0Afd/XuboijMaa+j3izwUV/0zffXOD8UAcZVfrpCSrhKpjlkKQ
4HrJqB6jeESUDB2K7EMobKikuH0yfd/XdeuSGauItum2oFsL+gT63eXqaTRi
bNIBx5iXNfX09y1TiUMg3ylO0YPOpnuNDF4j0qaOpUjiIEhU9IXP0rBn+Azw
k1+HIDWFyWOWaIT4eFHrsvhEHN5wjJa9C4B5kVoB2vrG/KiaK0Wh3GaAOJgi
wSQ5gIRwpNrJnyYTf3bfR8TrbAzLN9KezGNJSMPlqzzKcAn3mHHdG9XJYiea
ZF5qys/ootc3VMZsQBWR1xP1Qc08VgAP4GkBAmThKmOHCCRuor95NIdG4fA3
78aaC2azNV1TikKyXECr3bSDDEKS2Jpf5Wj5K2UZHb+1zlX11jBLUMeTCDA0
m6yvODLpmAHPaad2oYIO46eQ9UMGbajrCSBCEyiQoOA8N5eJ/y1txq1T2kN5
FsMMP/cZ8/Yr/XA7H6HZf29mjwe22HlzNTU0vYiDKIT+Xi9+kMMC703Zur/V
yLZMfOMv6GyrXgLlkMp832MqsdpaIyE/091wJFLugtqwkveQ+Aig1oIW0+iC
XWFk72I8JZbxBI19FB5XKnx8S6KD3J4iizW2Blrv8E2eWwayVmZ8gHixjg8A
Huyo5wQwFkyt8R1hiEjlPK2Dd25HIkAIVuujpS+rTSxWj12b+FZ4aCAwLfKi
3RCDkyeMxsmMGNvyJIddIH1FnVXhyzMSnn1Em+LjTo+hz3uP41EAgcuxOA3B
bfn17YtKFshqDcdafTlA4Sz/r978xBsCX7n4opTiL/KF3xA0JNSWgc2mZBZ4
RlWoXzjKfOQ6UrNSkxrbla0f2znPTz5N7nKrHu25jbGY2x7Uufh/mUb7aHOO
xvsKn4iq2wP+Xt0pKf0sCgwyi8SSsx4hGhp+eEubNbsFe8GMIpXDWhxBOh9K
NEF+RyLlPPDu04doOo/MfEQqXuXMGubIkYZvFzs726ua3NFC6ukWuNKglHno
L/pe3OC7lJ8Fiq1/+LwjMRtq/5VTDVDDJqMMX4/s13Aa/Bo2JQ+YCVvdIDjT
lBQRCn9PxChlqXec+LHiB/FaU9ZaoersHr0JdeEi7UEkzdM81rZ1oOV3lHB+
ntol25eppEYOoMT3zo2TqSmNAVMF/tPgkygD+IhmoU6j5t9Wi2iQBnS38/+d
YmGRauGSW7dqlq3+CmtSdgBp+HlDaIXrWPBmCBg0gxFtMpRaSjc5Cqxt6W9R
VeSm5Q9El3L90qmd8WFHnhS+aAJkm3g7FDVoY85mDBYICyuisTKAAWePPEp2
74yxxogq8qqrowDowUZ2omWdBhNFmyb9F/LKvdPGZ4MAQqkQxvW70wR8Fbxe
M4n1BVylaIHQA03UKjFIdXv0w23zVh13nVubYBj4BX5fsXWwYGCq4Q/o70YJ
TUdVb0Bdlyd+eQ56hu1T5OSbVpdNV1fRz1gOSq06o8lAXw1auo8OnjdiLp6n
R5xY7k78yjftdHnc2I/CPrYqX5HC2Njr5AUJ3hqdosztbPhwDWb0Dmv0FiRh
YitfBFL4zA+IyDFJen70l8108SjrxlExuALLtpVK5qJHMODo2Jmjvm//nv9v
5bAXbPJczwhb/ok4jQJ+JfU6r4PpXGVSHxE+kDQOpOOxpsH15MbEKf8W3V2G
nbklWR2xROme7emtUkGoKTjCMVcOpFfYEzyNb6Siy20QrDoVHiO9h31vgHTL
n+u/Fiy7G9kIL7VFF4eYqLv8fSVOrd8eSod+CKaYvARLsRbfYfWMCn+pCdk+
6nbSsK5haNKiS1z7vgH1OqxGrV/QRpkBPWvCAwyQaYMPuGdyv2w2kM9wjbDr
jubgqnYe9OyZ3oIYRg1c/XZMZlqW/JMNCQdXwahxzLfpo8jbVFJzK9I4NcO/
J3W7glOplgOwLQzZVvx6g5XPE6iWDgI0Hmg9cjBQopINieOQL1/lmRaA73Nn
cAVt156VWLSCxKZYzW1afY0nFcXogkwOBWtiATChwLouBcYXXhdNtZSuPfjx
UbR8+G5JrcSyORRKJF3NOuDL4poT5zq/ncxVQjDX2sIObGbG3O1AEJRvzCiW
m2sQvJzZJIXvcIl0lPj+fsjT27nDeFegdpa2R9ni825jVHkvMNPVpIDo5w9W
/RigsvXYp571wqrfIN070wnEc9zdwKmNcVRcAzEgzx2OBSFrrhxu7qo4WLrA
TlCJwLUG4kvNe6gH7T8jl9itLDrkkZIbuVskVwaFX9QhaqFc40njLqh461Yy
pIMLaHoPENpzQlefuvG0vyneRgGyPoDEgX978pSwzJEVybcpQpSuKL+XmECm
mWfbad6DQd+Tdv9nqObdtGoB7UTl7ZdI6tR4Qxd0YJ7y6cEBXJEftCjsp+qL
D4NOJHa2GdfMPtsLulM3DCMDjRbaNpVBXwNFoXXqUDlkzFOiu/azLlaQ93DQ
qBSm6UvsXiw5cG9XayPziFqquwl/R9sIQ5MtOY1vXi4ShvnxmqoJ/KRQuWtG
HdmuSnBHcO8u0xAGaxrMhf5NZ3PSBBdGRaRmyeWuJ7CP/EKo98oClX6P/mch
oHbAX4m83guueB8Pvy6BBgY8TjuYfDLTrAYLEexNB/bOfmCoeYXQ3WHaDMNT
N73pM0sHTG5IC7G8Ev8IMv9EZBt0MSHCViXzj53LAsWbWnt/oCa5Z4jvttKs
csA3BDfka+taNYLAOX8kWDVD+R8UpGqP1LTrtVopSyARYtorDN+IgYvbPhHm
gzCIQOsbEfwIBXLHHazFrG1QcbsBC+XTw5//HLawImaXX6Gx91HKm7Vxe+IM
hHEYRMvdKUJucrKMapMOkwPT11QlUX91N4BUfcUI7G8/0zkF2R9T4f2rVGp5
eVt6jm7mPpHx8f48Q+AC4t+BIKJ0jH8OphsBJC5Km6beaqAeHd+uoEq8bGVj
ujTC2qUtL0Fd4FLXGpycniZKSz9oO1HCgYfbhMvpW4X0YAYfLDNRq9bdo51P
7xzqDH9q3QeibIQi8iTQ7YHOKF1Yhbkmm6sORp45iNOuRLMMMgx8DwJsO9Cj
3ZD8tjvg5Bx8ca+j1SbteDiLZ4/prxrE69+A339bIU3sc65UYDGV7JG/Gmln
GaYRIGfhKOQBKVEUduGnhvc2jOML01tcPWYajz0KKBVg/EiqB0BVVUREHKQQ
RF871WacJMAwqj2wmxO9PLO9N4FCjOKw5muvMuwol8DuLK2atIqs+9+XRYvC
eGUMC2ShMkHambgCR0iZ7YkitX3zxdwOrE2ZwH2PGNgD/21yooH+Rs/EwdA+
71gCIhvsijUPY0bHam2BhBU7SzVPd4db2/bfqCILtcnc1GkAOylbo6mvDlL1
74U9koKsqRiTtmSpdbfjJrQIQIvN3YL7HboSBBv12w9W4wap/t+gkWTMXmIA
YKRKQ2pg6CvkjHkZXYqtBHmolbuyAGMjN77HuwDHO1NQSvZUUN8O2uKEPIkN
PjwMMK7A8qnaLhI4PpAIoLuRq11Z+hXdt4Z9KiGyoVP8ZunigDkltOYUAsQB
aeMfrKH8R3q8qMBEIG5tasHiOaS3PWNQ7V6p3MNWQ5KRjQlLCArpHVBFwSWY
H7hK0lFWDnUMa/6EA3hqxQ+4ybDenl/9p69x8nNZyfM4Ot5xaju1bp0Q3CGN
/lqDaazd6uzo2i5KcS3KcIOlkFg/oyzKbyimWx+LvNj0tIjxwik0LwlSdKTl
MbYL+eeBp/hwtZdqywvzdig6+t3a0JAycEntPbXv5fy1IKOxL/VjW76MnYVZ
lUuknyEaX0/e9QtTj+tqdEa8bW/+l2uf8/RKmG98BpY63SscRgB+4F0G88nR
DwHYyIkN+MF2gg55wvsc/eViN2AupVIjAPPFFgpW0gJOJKtu9mlU4M++OyjN
NQ1dsbAPW0hGT2zdYIlJsS0GQkiWbzSbnZC7NmOIzvQNCK6fRl1e8XX7+cIP
Y1YunFUQQv27nlH8tBUxp7GE51A0TdDGJUXakYHwYzGqRobo6YaGRG/iVqvO
PGN8jf6jVjU/WMIv3qZcUSyaoS66QMFjdM6IS8TZ6MSegDp24A4K1Efh1exi
fcNCrQB6FBC3GeC7zigd8tjtGZ13u9VbsEURB4ugjlTm+DsArxhK2KRRMmqd
6qtI3y0XbTZRLRDe2e0+Wnedp+RN2IJ5VUiQFkSgZtqfEtLihm0oQaNcxW2h
sOpyhT7ES6W4hsmh5oGNvY58DtFTJ8QN57h9uN0CWMe3VLiMiRPxTQriYrbu
b3n0Pv+uM4PwtkbC3evs/zkhu1Uv3/i84yLcYBZ7NGwiIQ8sfigcGZCCUvEQ
PRArVSQmYYWNmjOELeqUBexRsRfQUn+vnMuuzKhictdrQ7BuPPudQYLAocI/
2LNuiiOl4tZAC/xs1yA2Fn33kkQq/cZ7trqPInLxTMjcG1/bpkXYVjGF5vmW
D1qqwOXUk8VRvbfRm5YrvNF/ScxZ/4TLrnQcgmdbvggK9TKabtWqssV6KT8e
fAtRG59VBGGJsb3s1SPtCw6xqPlSyW+g6gOE4mClyKrPgvUM3yeABLYvweH1
YpM5uo4QM/zJqMzs7IVj8NmLxJE6TsrB8dv+MRB9wOLoFuHa+4mUiicMK3e5
dyCiYyrHL17ik/jMfOB1MUVCGZZuCNxuGzy80ct1LPaAvcyTJeiRv7mNg5te
zHFB12Ih9VeqOD7rUyT0da+Gs05CyQs9YPs+Cfs+BsUsWNelXzR9ll9x5EVN
0Ld88hLsLb8DT64God+1tlvInt6LoObEsqyV2Op2qDL1f9GfVs8FYM0Dc51u
74KZYc52Pmu1p2E3gHPqHGAslhLcDUoypsG7qBntsIc6HMkKX4EdGzl7PyGr
TpNlnr90bRU/eho2RI+OAYfKmerFA3K6rvEFtZXW8WwWsAod9GxA32kKMzKc
pExedsKABvoH95xes57xcIkTSPxE8IanhFKOudhA59HR6yDacQ+LkHFdoBZJ
L6LZ0Ztylq8V2wM4uqpShWQt1NOpoz4jpLkRKdENpJiPAn0Qd1MS+BwepjgS
c4qesulTEiYI5jYRFj0EbbAtCNc34A3inA2W6NEvULJtJvO68LbCoOcoEi4V
9YFdL/5SZ+NPaeYtW9CA0uOJadU2MmP1gfEpyjWIubHAVV2nMdOerejfrye9
W+88ZH2FopQqlt6iwdi9ZSccSSzLgndoAp5ZltLTxGc9mb6NF/fzSD9fc7Wv
HI/Yo07W91eHIFjnKXe2e5SnnnVYI0bBKXZx2lnRmmqidiumyLNTNAotRNgP
1DSGIDtpHlnNNMd9rLFW0ctv2DAY/0VpPE82vIue7BHsaP/zouyIWv4Xec4q
W5hN1zXtP/XlW9GRiUWmgdF/roWSeaGmP2yBkHCNskmtM8XqaUDMeY3h2GTL
X593a4B8jb4f5H0oQF23KN7w2SKzOccb6+7xllw5WkYqISvpiGxOYMbQUAkR
UZntM0ZT/lOe8rhYVnnWN+CD9/8MV8k5yFtbWhtB8ZCgvq5FTJX4rwXf03g6
CigfjHxRPIcfVkihl92Sfv8Jx4uTfUW3OC0xy3IsmnvwK7kP843e67djJS23
32Nweuli+9V2XMEcbbBzTGnt4FINV7ElmEfoLpsIMI7a3zjKOcgcVxaqaPZ6
EMfcrMGaVaQqhCXZkAnlputMYbQfxvZZiWTORHEsRAeURMfXV1JcAkvLOj2c
i8dsaCW4yq+oaOthOG0xYiOIopibpLF6LFQSo1wm9FfX4WL2/Zw0SgsT9hNP
NU7atb0wywjOXA9TTd4c1SkBrvtwkBZ9psUMNfbxgxvGEAjIyrm0n10p1M1W
NYKZTWywpQkXZisYPr9+mNVYHr/tlc6pPFMGZ41esTlSF7ojxgs+9htp9zpb
KocGLOjjYnoqvu0CzRlwwCq8SfzgTkbUVt8Urr+LHx9Bn7Rxx3SB+FOXPH/B
BtB70e6eIISDbGLtR5k797Ho1JrO56yeMhtdLeZ5ez9mTDJoTsdMZjMk+bTg
xK0/59goyF+HweBv+9dsNnQ8CY8HZfRRQVUx5w0jgwTDqSCGowWfCqnAdLL5
mm6Hv8EXmiP4N6sgvjnf+HH76Q6ktzQGhr4dbUmUi7skrb/ePnF3EekIv+bl
kvxZs8b5L1Tk7hWMSdA6oE/Yayy7riIkfXppf5o1ppnWH+dKo6uDAuCNkWtx
Y9Te+YY+U7nHkVuoGAI6KVyTVCS48V5JXBaRjK8GVxM+fBxnCQxl0hSGCnu+
q934UlOEJ+88bHc7dRCxQULDiaoVl5SQNJpSmo1Gx/82uYm0JX/pqSZpBTtd
kQNwA0Js+eMZcQ+z919tMJHblR1BdnkyWdtPOEvYGftcYmVHRNsIh0DWXuam
517UBaVRd3ECV/zAB1sgrd4watHkM7ZXvSwtBE9UvJZaF5Qjn4fPmrzQlNfW
g+DWxTB3p2+psDE3tpZYA8QXqk+ogA8SJbttSj6n4GwxTyrBhc+jR0ZLY3tM
MsdX41v7RQt10Wf+UzF8og3swfKUIzbhwvb52yxTXlwXRH3Ae7HJMrFSNlZZ
lhXuair7E/r1JXcA27uy2nZmGXmrcCLk2/JYZiusiavfAncXBy/mkbPR8x8u
Kglc3SHUsE8rjcLzbqEapCQSvfRA+QMeTkf+6pv7jRr+DfyFRcP6HNysfnVr
hw4fwTU2y9o0P0QOMu/DZZXs4gVsukQZGwAGsughlkRPDtpvY0ptR/hfENfL
L2utj3xCD9+X4nHV/L15tO0hF5FMIJi9W3hDUJldKe2+djuz2P1ibHq6tPrX
nMZ9F0aK7k04YZOgTDNjCF2/EX/sDxu5MdWAmFkMAzJxabYpFHHZD97gMZAr
2JujYbiQB20UXMmI+eUJxEi3dX1ajHgPBRZz0a+p4zEjlaV+Ld+3pXRorSgS
Z1bCUI46H8z4u30DPtz/hpDMwuqIJVYS1JbZiX7pAwpzm997fH7jM4+2wJ1U
glkA4dVmvvYN28rHuN29QjBZmdtQ5O4Q8M6ha04MKghJkMmFCozgfxxH3o+q
1+pEZONlhpjZvKD3CvntyUH/U4EBEpRp/Vm1gLjdcABgYGhTcQx2PvLWD0Hk
H+JWCnkNXCuNSaA/o/YorHgIFqsu2EFgBQB5EiuMdPf0r+TtN5qNneYWhKPa
47/xVCsMXO2070MQe+3t+AUKPqKC8z+OOwOmBQ1WvVe7f3sM5LQf/xbWJFmb
qs/TFmwbzBi4K5MZjoDE/G1kyE3kSwVglESwxADRtGTzkJBYV0RaN6F+I46y
Q+DUvAEPXKnoicCcyiWcr8u2PEEkzH1Y1X0m9OsEqtjkY057RAauURxPUrLg
+eNK5O3Dj8lIRrS6xVfZwOWo82V4P6pn5Li+SA90pCslXcRA58b1/68sX+VD
zEg7WgZVEEv26ld1qw0Erz/ACi17ksokQlKSqmLaUL2fKH1pE0ua2GEyMYEB
ZMrlHq0nPNz2VUOAAzkR+//HF/9QI6r7hDGRJu/XSSfjZMoABsvejDNY1HcH
BAFxfRTpVJcLm41cx3691IxFjHyXKdcTeLABMvlcvnCQFKmnPa9SrMm7YcSm
Tx7JKnNttry+epkEIUg6vYxOLh7cX30exs53BkbnMF6IiBcvyUyp/x+lEB9f
Eni5EHugJZEpJiNmdzzwIIvRUsGzhzBxSkYkZ3qgyr9FeliJpwV4Dj77R7qP
exr8HFjIy/SSmeurWqtVJ7EZZl1jgW8OG5EyHZt/3BO75BBwgVecgQaB9feU
MzdYcWRMhDJrqp20/CvLAuDEgUjoRJGf7qVMyyHZs5u4tJ+pyBmTbgGW5U1a
NlvDCrJ7W9srW+ZbnOREpRUtuFAeMCoj+GLR9Ik+7xcW8fanbiN64QgU/3jK
3cPg84kd5oqU3ifJvY5fe5seVA4fNS+N8ow7b5+870RmB65juL6f1nhAu/na
d3j5NVCZdXSkfqkhia+0NcBOC/eBy5s9fDgUZHK99ktNOm4LwNqN6MmlqfM5
zv5pizoFIqEYRFhza4qipR5yS9nsYorOMNnZ2/s0c18GkqwP9OO3UC6hhJ/s
kjaj6DGY0F9CDZzYtMB/EvV2TmkqZsDvicJbszTaBeY6pbu5I8Nap6eGV9bz
hEOXIuf8rDl5ouqUZz7FE6UyA4mkdk5Hdtg85N+WYSzVe5FPzV7JfKbo3EcB
BenhI3aOCwlU2OujnlBRiR4LDB2l2SRhsehYkd2Sf3qBoFN4Cw4uy1jZzNPm
qUZkyAuuqsb64/fEAGtskI8O66M/R2Ft7+4DmIwKTjC0HEePckK785iMUCta
j0yejLDGib/37JBWXKlHa5j76RWmPyET+ZptXxGqsDH6VFB7j7bUeI4oek9Z
lphpt2aGzOGPS97TcGYVgCE78kBfUa3IUkQ1rR70t5ElAik8bjOX73DZGDMv
hcAmJIJbixlmfG9IgXCV9lZTFwk5qFzCoaJEN9Iacj2xk5ohUY2dj4DXHE8M
XA4mqrAjF6NNAL4tI86NfTStdQ7SbwoauWjF4hrhcNBuClVBAXoxibgEuSE/
k6LJZZrbNJmvZXNDs/QEuLyM1z7RxReShuzPntgMRCVA9RkmB/3VhNSv+EEQ
PS/+xWxEPMRRAxClnslSObS3l/5LyD8PbUMaHx5rjFWk/Dtbc6vulgzBjF1C
YjTuyfilTqZZcvjlQUr5lcuqljHy6YrSvXtpPWL+HxFNZjUCXNm3YkAUFIFO
kWadAD7CckZyRbAKYgi1iMtNs4lJt2hVvZVIdEOG/+JvEziGEqqHv93/K9ZJ
pcucQdgEhiZGcixBr4sIJ8OSyeuoLsZBhpJUrs5MReAx6clSj7p4s8NRk4zx
VaFAdwQOrLchTlNGYw3mqVeTIkVgrwscwpzXiJ1NuP3oTt1L28kd5W3lNlN3
/s+1kJ9O2szg0CZFGHK863+FI++Sc3dR+jDfVKQZGjeO2ajRI68XAEdF7Pjh
Vnyk/nXkfuJw0UmyDr+BEyGGF1gjlLpcXi+x3qEIsDURN9zmocMybU/9JJnE
ZjerT4kME8LpNxsvrjn5A+r1pLxoeiAGLZMjq06MvnoG3V0MkeOmIUY4QNZM
QWjnzv6kraM8A0c7WhHF7CSs/Ab5qpvANxqxufWZ/wnhhe7uHtGt+RF8zyl5
OUnPdtZ6x3F8B3PlWHcxvRpEgcudDmr7j3eETP9vLHIGd2e2/rh7BwO3n7P/
Xql7cYlkA/Zmt8+wO2ENGTBtMl0VhhRU4HxfrZWX1BKrWaM2kP0TFaQozWam
fD0GlEJb4HMp3ChMfvg15bIk6mWXWF0d3+6YsGFJbGbGLeMl2qakU/hlkjlj
aPFjaPKs9AN/IcB89mvKomjH9PwfWPpE4WoZqw7Uiqvtr8jpUnfDud9utToS
2PWbXd0CKvbtLFvJU5RuMyUTU1Qer17VcrlQVbNOFIYRGWz2OUz6d/59cx8b
ki8Am37s7cvyNU/xqXDoNcF6MENSg8OesX/yODUE+3ZCL1nyPiBRv1MNLbfz
vsFRUZIFP/eI0DO9nnBuXRK3JNIYcEZkESkftS+yDk5dNwUwN2P1EfqNoW6m
3tKoB0HdzZ7k1AfUGIewkQhIt8YLkUPVRBeHmg6M7bJlHmykStGU2KdFtSvN
m/Z2PmT4Z61TxYMi0VKbbsRKJo+4JAPHijNqfG8VJH9oG7uKreHIf13eu8/b
j1lE7J4gFcmqf8wTdvL2rYmszTDnb7owJHYcVYLHqPxuqSDFS92QU9bE8npp
s2ZucZaPwk7iHkxCf1/QUwQ/zxHBD49aWQf95H+QEKGBSwwpnUTa9mgY7WKn
jBGcR4PGqqZAm4pFQ9r8h30k53PRvclrQK3Rqf//bzn+K9ADGviIBRIQqm0y
XVVihmuK/FnU9o/AtUEluD3GEPztXvPO1+qwb67nORWXdJfWf0Jx5uJVfdCI
HskRI4jks62qjfjIvKM2asUWsrRsqeRRxLCIYEkglSQSSlklIms+qQa0ukp8
BCsKK12frrs7tkrVfej864FG5C0hZ8OuUMcAbScsMEkNcUAL25HEIE67RbNS
S6TrjnOb8ahDRjb+SEy5t2JU+Q1pG4mA8Y05K6TVgvmODSbEpq7gkSuoQsUm
HnEz+KFvq/wKZrhScPTFJwKdTLaugItiF3sX2utZvMucNaJNZLdfQHHPtrG1
iFOP3pkAysiu/vjheLoMNgVOqf9n/537bHqny79SQlc7DxZQpuYv4uTl9pX1
28gByDXmUWnl90yqT6HIkVnqei/TfeXFKjFU/xEZr9Ji/0Tcs2Cy3xg8+faj
Iup61on5KFP+bMi3Zc4a+66Lhqzgq0cnauwHJR++wzBXk/44P6ZhY2Ivtlht
Ms5iEB6uKZe4E9lOTHfWrAzk+5satHDuykohGMHZKYE7GUn5qVu1ptmPeQMX
6IVYYajmri2df7/ryeYtLOnAUMT5C9BaF9/gUprfcpII5Jmk5XSaU9iUY70L
w2NJIjunC72cOjGEk6noAm38HgwK0o2nAZmcnmbtdUsHyi0iwY6WPhcQmIKq
kUeDUoeuSLcJ+votk1SkCA0pHHe3vzWNVx3WzEM2acBAdZ5o68HiDIWkwImj
O8SIJytvh4levh+xJd02oc3yZHbLCWGXRqwNpMO9dgmKKQ0MtFAZFjXwIEMi
YkJBgVNHcStP5mKkEOUFBhECNY5j5lVAmiV/79NQ5uW6+4YhAg0Ho5Ms17Ui
Os8hq7HHg88ywEk3mxsWx41mYKlGIoQ27p+iocHoLWYxAnEm2VaDe1ezeHCJ
cdsmDhu0/1OgWxnz5dlu6NmPx0GjqSd4uCovgwstwLRiJCY2hhXYNkc8Nuw5
yFNdl4ACPclLVkrhEbhuAK0YxAEaKMMq03rS3bND8buolZW1jqpCH1UW+/i6
e0DsPibFAoIjmPPVNjoI0otscEayiBVkUXmst8ALAo+RkuW8zKAZR3QVUtAI
HUIROsHgMAOZ7/CD1sSa8PsMIDyopsG49+Y2RHjqOruwXIyUbgmfTE7qrmIq
vE5GCxNRtPrOG1u1hh8u35GL1DpCp4xa6t3g0IKzT9hPy7Q12JFGqcaSxOum
jss+eFs802r1znjB+fgyZ4l/XM+CcjAkFndyn+AIAtrGzZcg5mR1oMY9O2kq
i85+nK/8HAedcEv98iwJ4yzU3nFgcp8GAKzbNe3O6BLhw44VLHYIpE8KZIbK
L11CLgFGCyHCsL+XudAongro1WedN5eZDmikihe3XO2a87kgU/LDCnjRmPyK
rpezHQaUGU9AVk3hVk7YIcuca7nnpBEN4yVo+kbziGUloyZuiU8oIhQnG4L3
Afc18vWhMSdc4NJO3XgGR8GQASl3Ts7VpBFwpu9QFFWw+5ZQFVF+KQFNReTM
qrbrwQx/LU+abhKaGhA5HJgpKjaM0QE3urVk/haxZYn5wJ5Aiw+TjfDC+Lpd
pa6tJO9UD4vNpAg2uxlMU3jR5/qh5q1/QEtJJRiPP7x2/IFNP6y9wwtuAtUE
TH6YvpN8swnLbleOVwZP2QXMv63H202waXeR624Ee1n/C9pIFvIDGFCkvmvc
GU6bqPRlLfAaaKhUfTP0w+Cpdd8W4pd3WW8E2dI/YJ13CHhqHztCw9ynVe46
pTuJcSP0N4ZthM5JEr6O2DOWgFo/ySjPkqhtKRre+8DW9xgsv3gOgxJGsqtx
vfpVNXf/wSV3HXvwmIoB94IwCnJEBIlKQKak0ucKpF5Rqh4PyqNArt7u2Obe
hB8OyOL58oPwzA7bZlibaUYK9y34RdRUq/4/WxdAK2X53fEfPqps3rrx1vpt
jRnAtZgdtfzDToZZI01/adtUbjP+GYKRs6UN1b6tlwYTkwm1/fhIlqt0d7BF
CQLs2FvxlLZZZj02XjpGGi9jgIeSFPa8qMapr99xmcMoIDkO1hQxtU8Zbrzt
feaxBMxboXZ8jVHL2z1VsT6Aa5NxF01fjZU6CTcgaEKnXhrt4vYA9A7rXW8r
cJc/heNy9IOA0KWsG996kq5js5FEvfDfe+O2pnknZJYMCOJNS6I5Z457Wz3w
FXwobEEIGcZw2/dOb4bI++/2fm92pKttEJq8hXIWG0s4DWkdlXqYRS8l29zw
CclkiHar67IpqS+dObfxmovQOLvpLpAhx925UOVUo5hTdQrK3JcYc1SYT4t3
rxwcfy3KFjxJg9NJfGZBfC4yYnj7b5omlUI3mdYFyzyyRXfNyHAoFt69WyiU
1xvaN4jpGKsC7IZslOYW13BDkCsiq5wqPI1oXuCiNAMuJP/5w2FWVWMvIwaT
n9qPX0G9m9CifvhbYqBsKhWRdFc6e/ITH02j5lQ4qlvLSbhaYu3cZn/JaxmA
MJEaqFggxlzSY7/udn/PJz+QvnHTCGKB1cio4sgAYffIaCpdmeBvxWE3ZZhf
40cI30w1C6HDy9YVRwlIVeWURthdMWpi0OF7WnPNObvEmf7URpH3e3L/fgnk
QRNy47Je2NxTQO9a2a+LqUxxCjcUL+d+b6zYS5orV+pCBSBFcReAu++Gewf0
9MBt7tl5zaemdtIj9p65oRzXXueTinHEi507guNQntxv7IroCfUZT9t1H1nD
unOZ5HeBmW1nUahWbJYYURDJf6bkPpAloLfnQ4HhzHHQ+fbf7z2j5j2GnLSu
21atQsZPZNOcV4U/CX1PlhZL0dsScQ/1KltaaIpRJmj4pxF1kjlEZQ0zE4D8
qjR/BwayLll/XUgWo/fWXAoA/ji6Zkysn7rbeXUspe/G3ied9q55b4GmLzyi
G0fj/dLbFdagCZbgSxyvD0HCqJ2bGLLK7n49NzAhtLCfJAZbhlxCjsYueXw9
/dUXKF62z0UYe/RdpvUlh/8tRO7Fw0df4nmTu6BlcPfTZhgv6bAAV2c43bEv
ZDfOvNkcQgFDb80xaTy40WWtqvJi/86mSlYkiAnTubO0eSNiZI0RJtbLTYW3
Qn23j9nyaII4Oo88Cbey4xr0M5kma/YHxieuyGr447eWudtgWf8ZO2jaGQiU
wYn/wYJEvF5TWBZiupfNN/gaKWVNaLKI2c9ku4GVsNAyJqtUM0LQNkPru9aQ
bjke7fpteBlCVkm0hbZi8N5aJT4vZyB6MOdJMWcNdxZ65an+tUA7R+LejHmz
Rnzw/Q9ArbPV/7or9VYrtNtkhGNzwJrupTJCyUskLdMs3o5QTBvtSv/5k5dZ
XlDkxt1hOhflzUXLpSur3gMshxTCRpYdexkH9o4t6PQjwe7w2/l1HYaI83F8
XkcxeHcfOONbOeSfnWhLhEEEYgmqACMq4Mo7jlnfYZyEW2BLPhj2tA1f7CUJ
dgXoDibWkchV/2Pic4PdC/x1+CIW6CNUieydkWvujgFRA4cUJxQU4xGZZex/
DjPJhV0D1jpwiRinOQ7axIWyv+2wbsVgC7a/SzRRBOoJSYlFcYDm8g14nbhn
OYvfQACpU7Z2FD+D33eC1oAgRZGmovTB+opjwwECczaQtB7lGVNB5oiZGcmY
AWxqLv6fdnjkKcpD7UbDhpBNmJLbfwMl0jxIv0BH/ChWB4QqXRmYXAo+KsWf
SLGtZX8kHnqIni0UJSfLbYcyMgW9OiSmlkBKIHLpoIuiKmHJ6neVo9KgMSRS
QPJKp/vcGQF7wGhpVSas4UjEJZ57AVSuf2UHWQJG7e1L1cw3VSu38ksYrXZj
FkIqIZs6oruBCUCUSgh5rEAcGYT0UrssZ+qx79JRASLvpZO+LN4jBghPmYVU
jth1Mja/L1CO/x7dhYv5Ypwp4QuHlUmcriuobqjIwVHS9pIl0hF/G6xODTq2
2m16MX47Fl5iGHWE0ztzl5S9D+nYK/9g4t832MKUoGld4Ug7sXypa5HHH0C8
sdrvNFXT5dFQunWVQKtF8ZSSu6drLWFdvIaQ/BhPjr7juZXPt4qqn1gEhyto
TjMjtziKVYPjLo/odmONZ7OFbP/VO4dPkHsikvk0xBmumsEufNWVDUHzq48y
lRWITSWvn3+uELoKiHeD0JH5oHQWSdTsCqAPq9yKaBfqqaZI1Mu0wZ3WKfTy
pfG3MJRnoNny+cLCP3c1F6RopQNV62DUJYkNSaWrupPrZSuLB2Cxf6ZGWTCd
mzCrL3pJYtS20426ccnmDvE4Oc5lmAtRKZ8ADNGJ9NjzChJICubLmLG4Wn3J
/LAaIIWu7tAqPP2ZzRdljxHSNbgEy3XmkQZAFc5aYsslwHuqkS84Zu/g0Z6U
YuGMi49lX42/8/b/Wkalc7U2LlUDDTpKsEo9sfODsYvAqjE5jn4SZkuemyA4
gmSgQcEilmRFxLFVntq9pSUAWOflu7fPNWtpiRGT9i2Khb5doC6XoVscw5Bn
vqf7MfQlrHOejPIwAxhu560+z8pmDp+hm9Iw8RRVPWMK0FnQBM/SvvBshT02
0YuWmBFCqp/vBRxqQMFFa57WhRMO3913kpAvG1ShPY1dGPdgX5nlI6D2aeoI
NjWg3N/xlj6yTclI6TJBTxAnYpEG9+tviRpNKB47ynN4Nc/2D88OeBkMCMMW
JHW8HNp/jeGDgojI9n2YmEJ6tH33g8Pp8naAOEu+rYTXbv10HctLfnFEYodN
Vvdc8h3bWOP6vjaX/HB1Sk2q2tGx+87v/OuyW02LARmjDGdEgn5jCdu5+sHv
dV/X3UcibuSxlUXOOScXZNR8g83Qbjl0E0SnSP6FrU6Jr/6MJzEh1/5t4UMT
gcgNBoqrPVkAduKBu9ClH71WZuEt3x+MFr16jn1ROyGiIjl0GtVAsZN335ay
RTIRTYRvUbmoHziypxGF9wVZx37tnhDaxIt9qto2cOtwTmziN8QMNhh/EG8f
8J5Af5dEePZqqNIrt/MTgfhHHDRuaDPT7pjlMotGArS2h0GpRGg5F9Va+eZL
mSPOYuzl4nnAvPG4P2lK1JOuxs/KlgPCVbDnUAbOANUDLfPuC0+qS1Dtoghs
rGA266ubRkQ2Snybo4XKnEQA0C95I0JCJ60r/YETZTaYzaj6xYk2T6Loqj1S
4iaQLzi1dhnnQ0hoDfLwVBEtImH3a/MZmAJpVQfRkvvCGwwu+BmFLdds/Zs3
1ixTxn8eGU2hNdqDBCJHmdYmBtTBy5y0YxRNGixyd/g+Icf5BsRtFrlezySj
QI+FeJL6BbR+MPxGTWXjMERr02KptcfrXLLDj9c1hN+xDM1C7ejiofzgqhzW
hZ6+mIUhn9icYfyxb0qm2KYId1BhZbeBG4hpFw0mqHtk1JP0nGZmsSXf/XSb
j2/31cDg43eIBfxzdcmKbWvQ4DpRsSRuEmCB+NHoulnIieXz86lQs++5pNfS
gEpJyekwWZkwjGJv+vsGODB8TpbmCTn2IYrEg7/OGesuJNg4TVG/4Tl+/5TQ
Lx1FPInzIXA15BCzesoE2EztNhT0X456qx+2CVfDnA+W7ScD2A3s+dvtQGAm
F+z5C5eoIGa27uSX8/HUVQ0WRgvXqytFWtJdUI7zDYZRpzp5VNjJChrzRpK9
9nqTmVwK2qiOvgtmAziB2doSjQlmGL5e2DTJyl+935EtrpsFpKeH3FNJ36nN
xY/NikjDRIkj5OlT7sUTCYHAqVsMqZZA7fE5wi2Ex11/bxHozYrcNGUCknkS
B5Ib88P1Vq8P8+DngHjoeZOeFPXKO0YqIzkbHLVrcSYh9ZdrXKdE1qBcx+gc
o2s8/aLLlg0N+FB+OXA3bTH9n8t+b2Nb/MDR3clKfI1ROL/Fd/oYHtlDBzbQ
/Af6WyKi+b4GB/mTaKC/RrENVxC7hqDZBkLDKmiVqzYSysjOrT7pfAsGdx4D
qMacLOM/E1iP7vvj11+fHLfqaRReE+fzwc745ddfVnqyFpaejQl3fqM5f03T
VsQExQegosXTf4NIEWf0o5zT3UH1D5aeIT3hsYgjsgKGyQ4b97qsGf2SVV/B
ldWH08yawQY7Ih1mNiQkxQ2ObTLpFmSOaeplDuWX2JiNK0J6M9PwFg2BaCsL
llWPxuMYbbU8Iubt95tMJ2IZ1X/07dtXfEqIdj9dudrXCGExeqBX/Sr1ggYJ
s8sn2BX6RCT3fPZ9RYJ4SfKA63zBp+qHoxtz/8T0zgnlFkXfJU8BxNbOeMkd
xnLsXWFZVppmCSYyRTCMhYDbBPazrsLlztvbWwH4mFyoB2jsDTdlDQpNjD60
ewWfQ3dRjE4UstSaVsrDWtIfezNMU/4yEr3Vqg0mDIoWMZCgWvppOmUHsDKM
OHFJ8eSsyykkGz+Mv0LG7p83HNrREb3w0gYrni1r53LRKCl48bjyZsoADsIK
o56+ikkXzoNOiQ5/quXTkWQon017uzbNAcGv5I99X5088KdQqZIE1nIIMD+z
8qxTgNKhaDH4num/AeJlghtsvuwlgsYIqikN42MImXaSoAklcOmbkb5XucSH
+DoR53oRh2k7MzU2ydaCM6Uid3pECol9yOVA5RmwXsrz7ra4SptWWEFo5en7
M/g732k1sMHDqTT2ediI6tfaSTEimyDVUATS98lmy0YAUmaiNAbpndx9j4fq
y77SyzqJ5YQNcTpUtwZOxWNr75HMXk7/XdEk2tyDcnrQJqWRu6NdY9ePcA+S
WlT3SwMn4Wol0s32W7PzLLWrgqN0SH5G2gWG56y2bnswX4wXxzXLzwpum+kS
lOhUk0Pgd1fYWqm6y8pz2e+aZyTff0oG/D15utFWihA4NnnxHBQrxTQ7Jwx9
MnW+QDrRv3Q6NmbMOEKX+RyIWSq0SBOYRJciwkrbRgfYe98F8zz104/k5FiM
ry8RO5X+0q0YiYPenuBKizaN4NTebod9OvRkmcxAsPZTD0nZfDG9/OsOIgsP
kiZj8D4hu4ux8XLU2J2xUkIjV2eFLgotMP9q7hQ/zFh+Y4mPQ0DDqRe+JFiK
gNHPsl0qj0mFsvQsov+lZnoUCXEXszQ6TDi+NfdEbu+CkmSYH4hQpeCE+z6p
J0YEkselpAAdW5C6m2b+Pn6cfQ6A5KzwE5Xvs/AaFh03J39+yZrnxY/+dp2T
Te/BbvKVsdhhg3hpTOX7aRHzhxapQ9FqhrJ+9eiMop3mHx8uH9G9z24xBgih
Upux6XNQK/oam+7owlteiA1R1+DVNEo/5h0cxG9gdcWwtNoN2WANjCGNx6e7
61TIlBcN7FSYf6pvy3hMpQA0zFLBeqYOkotnQ6tPWOHL5SpmMc8Md+szxawm
B3EfS/0zQlOxjZENstDSkGb32BOKnYpl687ItFfChJX+uIAsJyOnNJdzQ8q0
CZECDD66xLd1N6fY1XaDnI1j63leP1Os5sr0kC6O2k30Ml0fvFaky5Dzk/tF
w6iIDZo8dR8qICXV8YhdKbUlWgD8GRi5tqVGkW3EX2WDBWR7PBR3bzzLzLRN
qwljETi2W0yBKNnE1yHPo0u7Ez6qKS+vyXJNshd+lLs23F1OpauZdKBwZVEZ
fQc0K7aj911G6CMz1L/6EdQduSZvcDEl0+ScRoyKGgYAgMed9PuGxz08mEhj
az/QdHjooH/a0Y8sw5YmrF7hfG/WcMaB2zdfxwl5MYGfg35dzvtaVUcfOLrZ
kWC3S1osEXbb5IpY6aHenMmkA2BxRHFn+/6qe0HyyHrmW3zByk7zWKhbpekI
jeQy8knC+sH7zFniLIiLsVz5RJM/6E3sO4fG6SI0DVRDbBsue8RDzbMRbKxo
Hz/v/s72U2lqjLsn170XI4jHqoJa9hNdBnudayb7O+lw5bBh5SKU9eq50jwQ
CIXRuFXAmUIpyV5OeOcbzTu0ZlIEW6yYRZO5fVBVifUGFjLBbyFWuP99UvTo
fHeCFi/oqSt8o5ip8dYsZGqOpPHhYsMt0aRzjGBYgEi1RmGmPOUcTdKR2gzh
/m42c0Tv/U7nFyDh5tdpgDqK5Ky93iYxABZ1MpT8ijiW6x8QQOpPtgoFldC4
tyoFjcd1eIgvp6Gi/qulOnKmFiGM4cvOsdEqThQRHH3C1mAhpUvJilfEFnKO
5rBKZCH7D/saV5x1eokumb7Pq5ONFzd79D14kMmLnisxkZ3PP2foZDeRiIp3
5kJOGqMlMnOPUyDkJHyVtSiLg1xHM6DznxhT9cO8K/qrNPOMf+CV0Cshek7E
tN5uBGl2murrkXXDGjk76x83jeWwN+PB6dR3UgmrTf9DAdmyCVOGidqRfZUy
4/2tuqNjiXkmKa2DYX/qKctU

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGMeg3deFl3f/A42YLjIoD0xDSIAMsdcfR4+Onp/TqrVIRMZka3FjRzQqBpDUP/0t+yh4lcSwnG+yRFYr1cE9oU4hmFpAdJkSvfdVgdy7Bj7ts36MfTQLNXv5YuT+rMYDet3uP14orEizbI8GC1KztLwK/+D0d3RYpNoGILarNUBePrKyOcAEn6s/Sbl+k5RPJlqKC1feV1fMNza+hwpFfwlnOmFQbzHdmoHzc9kjJcU4nARz9mIKp97dsjQcm1dkwv8siTjOCk7PE9B0/vz4Y1zb0dKQEIWtaxjgQ9mZbfPWo5Xrc6Iyl2Gc32xN/CPEfxQRbk8ZmUCurbkNsfa1CE/FOIci7J/3ZK9qwYmyzU/B98UFC3njEmel+Xgncj0HN9ZQcqkBDmPOzsi9iqVZcHlCq7r9ZvlfeZTfATrm1XATWbYPy2oEw471eQn2saK0VideTvvfdQ5gxAMBEkzN1sv8DdPo1npavR3LyIU7q27A/mJhwFztRJdmh9pRCOnBKdGcYM5l3+r6wazqhJlMIYBfqId61GQzTyBH+658kRfGt4jgtTdr6uiyVtD9GWDlhNU06HFf7IaiMr/LICTr0SC/R0W264K6TTxlHloW5XH149bG94f/55p1D3Crve+ZtH4paR8jJ++hKBpjPx4/VZ3U7uefV/RoQMNLIZlXuSJZv/tRSfc4JG+jUZGW+/jh3z2nZ+skO+qomZOuRIc3Fap4hZSOg6IQELDRvUU0wywmncoojOH6FBpBctiAmADAwFkOHER7vVo/hJ9WCrJcxRy"
`endif