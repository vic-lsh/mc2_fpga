// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K6ys3UiyzVMq77w7sj0+urekaLI8JdDKpteWPesap2ICbm+HHu29FSITyEUn
8DBcG1vnDBJ7tYHgIGIwcdzQGutwNq7bYtbNwamrm7kElgrPYU/Dccf4DtSp
WKDEs9Q8whHlcWiuDBE2SghB+dV1KCici3tsWCzLLzZWrWtETF+6CnufVB8y
sxD/afv4Yw0xpio0NEiAc7/qkoguakJvQXIH5Ghe0VYiB42fRw5J8t6fWzWG
O+e0c8nVyH1l6/BAkb5QyZ5A+UETqyx9DZE9z2ePAVpP3LKCpl2NA4ZRxRYo
3TYUg4Fke3YlaMtZe1JOec9NB1Iba1xOJr8El9gAcw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TiHR313Gmxa/6B6f1et0lG+EGwWsPjMY82LCnr4wSqXiEeuuVrDLdawznwib
/L+1I7sLiUIVl2Dj4UAoMTUelekpNMI/fDG0UVVVjwSvlc/BiqDmrvDQeKsS
q271pHv7xpfU9Jw1bN8gGwtKZnXg/y6i9AlnM0SVNrwJZCKwXEOFbUn7WZrX
dg8xOIsWJgG8sw6g18MZrA6Dnzy2kA+KFkJPbp6BPk1/oBLfLz3h+knNG2ZD
zWIDvu3W/2FBITYFE/0u79hddx3tusNOvA0K2eRmJ+HUzC1ZXiKb8hfFcocJ
RJGK0GzA/6ss3sepq+RyQTtsgI4+pUwwIaWtOgzGDg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vhQLj8z4BLwFjzj1lJ9WG5Rw/nBkV96CFwwKm4HwKDRkbVKVrfaupdI9ue0C
V9HQwUz2O7EymgOkIvhTQxzPaTtcsE3Dx8+/s2uFuwkn+BBYSapGR7nuM5tq
AhHaMbHs9Tv75uA99M80PNnrjgEEVtKwohCzP2cYkO7Zt7pg8QRA5r2UcnoT
5hAoufFf4G4UMye2P4+yGVi6lxw4UzDbIFe2LJ5Rnn6pzRIExdD8YTWRWZjX
w6UzVUuphFX//4vAJlq1q7RovGR1wkfiomeZlv8D8476+Js9Gd9Qpcz7YkKj
zX/TAobZGNVraGEEhqwO7L0bU094GI+IbAljPY7FVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gk10DMGbPM1S6cRGAl2lul2bT6lQtKbVcNk4pfrmkaOp2ZNHM2FkSIdOGlwu
lMgrIQPC712IHt/MAFLwaRllBLoLHsWS6QDllioKLzQUyCcB5slPW4nNBC8A
D6/Ojl9UBQKZIp3CDInemagE2r2yEQpBVUhFFe55R4zMZ9/+8JQVx9WGGFqN
Raesnzlv9d0vp7NhGp8tzGAO5xX9Sh+GDe+QpPsbqhtRaA6DY5O8VBbYNZBs
XmMZ4AkZgiTUTiZ93bgLKpU/7+GxOw/0brfq+mXFabLnmk/jqKapQ6Y99tXZ
FfnqnDPuZCtdYZfuPaImrndKsSf+BBWg/fsrZ/lFTA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L8uB23HTCHyv3NtrWMdX6Z6YJ47hX3NpV4oCGrPMiaBMCXgy2qbvmW5ZQLwT
ncs1EJqezBv4St/wDtiDBcaP21Mt76xHj8YrEciDsIf5kTmu2+Z1B+HLRUu9
fZguatIO67eLANG9WQ4Mz07/G0C1DDFDjGzQWgVwCb0vwr8Hn+I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sdFsRcXShiDX664cxKVzw/0EHxmGN3AXS5Zms4KVXFLAojTi5iZ02Rn9KLCy
TM+7/a6dsDcM9wRQAYJ0+obc9YTbi9Uwzs1ndUjHhviEpmYwEcO0VD4i1O+k
9XTBgXh7b7InbRjaz0qwBEzY+kzZNt8YBtxtRDL8HeYq/W9yKr2waDaM8/2r
Sn0v1hs1jm4LFy46BNr875imUCG/4Ke4jpR7mDmuEhgpqZ4Qu6xXqpGfBBVa
pS6Ks/nTuKF1OQHqnZVRg+ojLnXHO5Pyfo7jnA4tCzyZnx4eHvrIp4IfcDJq
iVWsZy/v/Yv8V8dT0EX0Fz8IFMdO9n6c87aiwCfQgy4BIDl2XPT4qswuz+x+
D7oVdbGqXoxJwvoGKoTX6RAXnXTRkCkS5ZK0S4j8hcSphI9gn/bgxqzl++FT
w4mzuhl/mT4smLueimOAsIsxo1xUlS/RLKHJEII/H3v3LhMIC4Dc+xAGwH3w
lkcwYXAvD53OFFEO3iWVaNeH800pg2Uq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SuwWbbrZg3OGXtUL1mNwlUt2SpjU/qIf18J+DCSk68miTECQDmo0nl4MIBBH
IALGfAueVy//7vnN9/2ZWspHjNltcqzFsGQrbE8Yc8Hq6QhxPKO4HH5CFCXf
u0LlWY5LQaa7JcUBFg+uyCGvMjWxJK4S0C/MAVqWoUiN+AGDumc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r4wISlEUn5m9vo181HAfT/fKfTfrq21vnOivui6kFWhJODnnySIrHkx3Ky9K
dHQGzGFUEEHu9RgXjLT5NmV54HNYQkR4IZ7hHvhdUlk45D0TOrTxduE9Swdz
Jyjv03HTX2T8RyNJ56NwvMUdxiFiazjR/SI7nqcAjLegueqrid8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23504)
`pragma protect data_block
nc7C/R/7MsZdoQaftrzKV1sGpUk3+zx1GGtearEP+cZhncGjrdlAQCPAWhLQ
lRfc5yZqARfjfkpLLxKBDuysBmcoV/I/MgbTkUJ+MakMBTLuWi6BReYbwFG2
X2goEV5Lcmngc96nUrkLhz7khIDmFaDnNcBaVl4En4rayv11gzutu3pA4wWg
+XH+GEpQfvL72CSoQqb8DWx/JKBsQj1mSAQ46pXd/t0KygLNtRSvytezrKdW
rwwIViM6SAI+XM/U6nWlk0QhwomH+M8YB+9y4mOIxrnk/qqVYRcMwpdID6LV
/RPLh4RBATpDUiqZqYJY0eUUZXPYlwLYUBH9RFjl8tlmDjDpjbjW69E+yOnK
yFT6n8vcM4CsdUcXnw3d015/lcPjk0lcuk6TSEXvtRV2l3f4VTLRLEHwDcZa
VdVQ7wHtEY6D98jwNFI6ePXPqNte4/gmn3XgIdi78v+qWlScEbEFQ1h50LV9
GBLQmPh2qxYJMGfIb2FIQowuk/GJM+rvHuC7HviJ5fvTu5Uto28XeLYY8dQ+
/xBX8sFZ1ANoqQmdoBZpkvD8IPrQ9i9YrQo8jcuhRXMNH6OiKjv+t/2zFIkG
0PS08mzI+UudMiio0IyoEfj95/s2riaIMPz7cSa4+DlGJ7TavasTDCw8sWcA
5g1JeW02r73o55tNNZu+XkFbF/303DKCsp6ZKA7W/LoQRS5jSPANMKPYgfXc
ucT2VcEf2IF+L/1AIR1TwL+E3EcgmpxyqU1YlcwH2jq19DgmdTpj5Y5pWULB
LzT36S9S4TFJCRXUh36OSxtvpKYzmFJOTz9YY+e7yKTzuuhBjEp6cNoJqcNq
EvyDKF7c5l5oIasIfYceTm6AvttuCzuMIpxmQO1jagK73f2B5NdsJ/ayzesW
iEttUW8Y1GirlhW5suN6CWLL9kA5004qe35XZ/IcOBvqkkoRiFXyq1X4M5K0
5iPWzv1VoxzGDFVvIzemnIlH354YSwl7BlaimLfFdJljLXXX1ksQpPoCYqUd
XzfCAFBI+IZnFL56xYKbLFvMNHqsLCo6B/c0LHvr9tE3Vr6g1Bd8DJP5vg9l
mpEOt4eUkPFwnbB6HxgfoOgLS/bl4/XRGLeqvEj1l/zctQKyyBsNLfIo7Ahs
IcYmfqjFD/A0CnIfDqs5401JbFHpiKTtZURyQLYyx/CcTpUynNGl2awxMoPZ
nEA7T9tPhu9Rfu1LSr134yFxrtJIi4jqe1x6n5Aeae+z8G2b2lvdpn+MeX88
TONfYa+i2nSfDmp1XY1UByzu+x4IaJ/22yeHqf14Gb6+2qP9pq8PtXnqdkfp
ONuCX2MNObSn7+zI2n6iD//w51H6pIwJbipiF+2CavkXwVhqezhMsIFkcI+o
qZwvYzu7dE6nGqn9/MvGefeZNj1Ii2xjjPpnGGWWUeIC+7Um950MKkjC528A
a01VKonQkIIbdzoLHVOPgJJdu/IbSLEUznnP6DUy8VSNJak0VZlYD8/zCVbB
nXzPw7FcU2iHY9btBSXIg/sn+9GQvAY5qAw/+rXSU6N62A1qT2+8RXUyGbGU
MXlKGmb/of81paMGmMFY9oHPDBrBNio5YJmPR4aeb/vga6ZU6FEfcdVyKxvN
EwW45AxwE433JYrmJ94SASiXKNwFnFJa41EAYwcfwLA3GqwWS7MbUBSHX7ac
AYTiuJ/l9QM+rDIYB5RcOh9ZwXKdja8iCFlxLIMu1dhVaJ10mhWWMgEj6JOY
gw/30x8q0Fq13UJFIyMIfNqetv8EyCAbOFM7iDcppkey50mQayBonAkKfSHa
QLx1aWtSoo6mZJDbAZAYyHkkf8WOZg+YljJ5g81ki9SfBxUfWaPajaTpQTzC
gVI9BpknAgqrMbq1+s3W1bZEy6+8aU9jShMSeao0efX6DljfBJPQE6alk0Oz
FD64E+Zpb1O8aX2g605b5dBiHGKXyhZHogjHY+LsJGNL7AfpVEnfeqRSeIN+
uuQK2uzWXlO11OM5BRnzU7xC/TsTTWTdw++wOZioJJ9Qg+1x6uoeycRcfwv0
lzwc8Su86rVqGtFWDFMcUppVYqy5OWb55h6ZO+KuvK9iWtK/Kqv0MjkAdE6p
MiMaSljkRvKBmSkC5rUUtUeQ4izwO9VoKE3G8qRYGms5w9l/0WWepr5EbC1Z
8bAVQcE/wWIGYSoWYkk0mhfjh/NDjB0nqtIDLVm24BLIgS2m+pZGiPvB/8JM
GbXg7YsvM2TbTdKEmOKeoYDozrsh/+jNrCK25nwAhsfp7oMjuqzBjBulmhTS
WKZ46ERZrpSuvhAB+ZvKru0MbouwgObW+ZthxAeM72vDrke/7Z3w/P17KA4Q
58TfH24TgsOadn03m0DMEp7mvw8YmxHzXWBy0O25TwbA3EPFSSIlr7PzDRib
8rhY/0wOzeYbTJ18lV7T3rtDXWA5Q3XitR41F8xUmEFgfQAY2tillrJOzFa5
beqzr/Q7qtOM41p4Oks6AtCgLKiJCC/qloYwLZ3u8nBvSsdWV71NrXOualnb
HuhV3NRc2lxGFq5ilK+giYleZR/oQ4DSj858VsqVBe86dJAsG2E1Z2YOXHpf
CwDwOmPM99TCYDXUU2DJzFEkqlhSWpV/zkkR0tUwyneGdjMdD/8NQXwRj8U9
AhzrKpB2/tweNpPOCL4Hm7KXPTOV+8N5qt0IdijA8/qdKfv0seGHz2VTjeib
Lypgrb6VzWOkYLJxiHXK6s4alWl9EZMao4R4iHDiwarg+xd7/oGcXsACHscr
KqNJo0TNOqKhNCDya1bO4UCGarYKn0vb8jH6clq+0JX9TNOuhUfUOCIsIiqR
e5y7yqD0rEcFVwb8clTaVTA569DVwczWQ1HCqCGMnYt6NNF42LbWBMdOerVY
qXAVLWdY8U9Uy20zPSzoUYz+Wgep1/pYd8HZOA47e1VOsX6Iod0t+RJrpPW4
68DVCaiPoQ1x+c6nAxqVqEM7ZHUsABFkjl9NJCm7UkvMFGMya0tbEo210Bby
53zcEnleSVQVT9uiWnw549dGLCmKJRzzCmLpaJdRWfJi9vBQJkwxVBXcwoGw
nneUu1j04b+16prtWJJ5EKmjp48Wh48/K0b/iHJxHk30kZ16JxfvK5a7r1Ee
VghjLhhisQLxXAs5N0BHIM3cxwVMkeaoLSg12OzRl8+KMZM8nPvR+/2b/Cmv
hUzfOJudTHrMSGgwJ4bs1X0zh6QRPBOVNXXk1A0jE4awkgKBxeKeeQeQyiIS
/WrGavspn/bW7qM2lGAEIUogcpfWl7wnF7h4KyDuax4q1HXHvclzPSwr5ick
yPjqRDSepkEx+IgQjpdEi0j+b+3NBXqLYUInPslzIKtSb5ly5SRn+Qsa7nGT
6GdvCYAG4no+mv91Cut73C57MoJdn+sJFtsJCkIadgA9cS8aj9O/eQIFAZIf
2+HSOrvnK3cjJqX2wlfOyDO6WrES+JSgSft1bR/RJ7heOxFqZNYWSD8/8i8R
03jBaQftOeUolB8nfkYl9yKMi6pxTd0JJQdMgMVuBtgcCokFIOLlozzXu/BZ
LncSbeGDkIs8qDAUrhDdVqbD9V+AGRR3kI5eiZ+yxtnokHk6iW73Eji4YWBr
OTGx+Y34MpGFc2oTr1wyicw5SQkd4SwO8GGYViOd8Le2WF+cdnygQilXgSt9
vCwvgxtKCiAZBmNcIsmRFflk+NDa/RRrBONs0ASNjQ9Cx3jnjEDkE//tS+CJ
+q5HFBse6uPmcNVBzxmFBAATWgM3H+MMq2xiQkk3gkmOAZqFe8lyNWrvtqq1
nhVPzpBubk9+B6Lxh/weoXtISwWNNFHNOBM/TFlSKB+4Wsy0LqP4otL4MLEH
OqBrkes+HSG02/JVQvnSr6P909Y0+XIioXok5zZD/UvfP3JscyOM3Hl2UMIr
ZVZuLtMAdX2DrXFX+OnKWweJjVmvwTB7SHgR98LuIHI7lJQzcsUwoyNY87lg
BwMHj7ZuWDniag9VYEN4/knbFeNk/wBthBcXoI9RN9UNB8MYTiCsjq6kON19
C2vRaObi/51cZvpRxDPer7ZWricwId/BdlnLqag6qk27nRpALqEQ0twcmc+z
4TX4egeX7U+S4hGnRz8JX7dKb+j25cQWxgKau+otozMrFsVYo2eKEHxR/VKl
DH2Nj3lAygx7NXHt3vxmkTqj48EZ/6/GW+hl2gZRgZlA2vUc4GDERKxLoXQl
JkgyyDPWnFw6NVKGWvV3Ht1Eexc2Gv//BA2XJ2aIRPIG94TYVfnY2FWlZQG/
tff0bNIDz4s6iI8M2V33INK4ujDFBkOmz/HO0LLjpMs04Sg5OIKy6LT44say
aAQqHIwu/qgZ2bcXrIhyMQ1t/rMY0GoZCDxJ5QfgsuEFDJOV+EK6mzLwAkfg
5aIhtXWX441G8LDte6bFuwvVpzIbslmGZgjCsDrCNOcgSnZTRXV/hIC+ue6v
8opsmhq7ZwVDCExcfJZ85bmC7UIQdCc3m8+1VESWUv3tBPOMy/t961nJR2yA
0gQg/JH6HbxIBXWEmhhL9jkpbYxATMqYhIoxDYmB6dJSt8BxqwxrM7/oEhJD
9Mh5lPzpDTYg4s9VsjA+TUC7szhGHDgzSTvuZ6UhP6ksJWlUt3LVbkUNzVHN
OwlS9AAWrmwNMXy6JPp9mg15mjIGPkwDRbpSy2I3ike4beNJIvz5l5Fj50rh
HOhIGx2RBYu88JxSmRKvKL7QP+0uaESoj/4+s///gKyn0J825jdak1D3W8Yl
dy1iB76K8FB19tswdap3ggI9gjMsRIZSCzCczsgFUw8Rn3CTUsJbbKMGlH96
oYAi5w6MX8FfK6v+L3VUhhyWRwAbuKUzcr8ItSVqAbKVKQYHCgsgeQyaiGgd
DxAIHhnVHl1+Nz2XQZGjZao8eZgdileNj3swDYkewGx/2x799BkJDcAXyT/i
O7pRHqIwAaHOTZc0MY+cxqpNPiCeWIv4wbFopVZ+gKRC/XJZG6pTJjfh+FdZ
w6DfR5/tEqGYjnu7rKzjseBWR5UnXs7XrFq6FFyp3buQe4DXlrCkdM6umBiG
JgluliAbqgm3QC+gjcfI4HTUwk84svp/5HCat/nLT+98mIA9HKTAV9u6BtYU
RWiU7oMuCUB6+OxWfAYlc+s6fjgLPbmZO9PiYpy6sxzSt9y3JKiRb2PmoNOC
AxS4DeVLDprPwSz2zfBsDquJuzpfcbBqcf/lC7f1/G7K/1Lzbusz/t2ixHAH
lfjCBsMNuV2pq2OvZSIXjebVkSHX8jXmrl8jnaRdz91yvDhfNh3iM6q3/d9G
JGF1C9snvKkeHPbxv7IPTBzWGlD9JHi0BsfqZ1NjQggTBDcUbkz9iu+p0BiQ
0ufaU0Kb8efT9JlaYyMUAwjAWWCmU3SwWSPEmhAdCRU9EYNY+Y89KEmJI95I
FXAaiZoQM7MJR1jwLgD47STKU3m88wUjtx6gEjSpAFm+/t5jUxT71YiQuueZ
MVzJtC06p34YH+NQc8+l6LPkSxnEK0ym3ofVqnqaYjRhA9RCAzv1Hc/ChoFX
YK3BOy4npg45IWBZk7rbU/gLF3en33sE6LpBLHbCdvUVMSZ7qNezLhfG0adK
VQ7xvvlaK7SPgiy7dWlDxBAB+1bMze51bTH5rMrhV+r2zGeScJCZ/8P1LKI+
GuGNzAbOYG0w1zpvEx73dAE7keAY/rT7a1A0llXw6vBTf7b4GTD7jijmMp6R
qMK3OxNLf8lVbL5h/vKafOSFhspzwDtMJxjzOl3QXts+3TRdmm6tHxkBnlU3
DoI5SmQwO9al39hlICFgOYR/qm4XxCvS+R8rvmlhPNHzhig9LIjsRZ72CDFa
zF08F6h4yBA66ZPXvVVksuyGDXLBbNWOJG6r1f3V0C9ZS3MY8u9sgiy2UKBh
orBhApxosDsAR9rYFcAYRTx8fdgjgCgs+FnWEoYBoUWgeGllwJFrGA6JlDp2
HMJcXa47Ez9bY46JBHRGvRmyIm4aPy6YYSqKnu3U7UiCaR2i4DRn37wZVSl9
opyjVGMqDxbT5eYdA1fZdCwWndZd/dNZuOsykoactsuyI2aC6jrkuqZG253x
AVLwuEsCY6a+HUR2oc2h8NvdHQ2SGb8ES/4dviHk4Ay4kmuhsypqgf2E6BsH
iPwZzylq4J+bq5SVZX2/ouDTZ0yFtz1YDJsj+VAFrPrWVAtgcDQ+YwrYDkpm
JspmgjssM2YtfyW5o2p00miQjpM9VWaUXo5HhTjC8i2ydufSarbpEawGEKjn
+JENxqcLCGIUd+WI+QYnB3TSM6kDUWVCS/FqATRlldrEMgtjwxM/Qm1LF2+o
MWQ/RzG8JKFqNlazhFmcWjeXGVHp6cVBY2BoXtBxUBA0vhE8Qiyh1nhji/2A
gMryiUIksqA2Pg6Kkq8igrJVv8dPsZ79OECOhVfuS0Ynm4J6J40VFwybMWMb
yA3zUIynC2mXpm42oEeY+5qM5q6Grrko8+Efsvt+zFzIk6Krp0BQcOpFGPGw
hcuKCodG9mt9/Q5k3vH1m68PkpCDA5GIT52QBec3pDFX4wiWn5pmriWQJl/6
PW+WK06Z0mQ7qMLJcW+m0Q06gl1Z6+1+Pog+wjzlrPZIF7bBpjyrQc1Itqte
faS71n01G8zonuhCcj6VY5RmaUsGl80THYRo/SPrwueErM837wO8MpGorzep
UXP/EL3PxY/ny1B3n19gY0JI9EjFz1EJdnfWRgSlKYxIcMzUoWwcZnZBwsAO
OMSOAOZUY348yi6dt+VE15q6T6QTvU0YhVqWREM72AWcH/1LZA9PGR2MYeXS
BSVyiKYFiQz8j6Y1OM9hwFyOiydyasviq9ODFP4wMPQji0GdKmlcA6L8dNNB
yKBLABvNaz5F2J8xiVpmbPKpM/jIPcPnQ8Jyd/oFCetmHgODEzjJ7TuvWtGk
O0irzSTsA6sEnJLV8MbCxj31PtuEpHclvlUaPn9gQP1wGgZuhe0quMHjGSO7
d34nFtLh+CPgulUw1Vb0Fu4Fw7SRiqvBj3DDC5J7UPEwkx7LviiTz5k4Vs6V
UOfJOGmOH7jKla5U3EPD2LdbfYuYItsUSZsEYWX3Vd740qtQiTJKUH1DyQJ1
31ZgGCFaBWl9ntS+VsRLcAF1esRbJCcYkxxpaZwCRNPHCy3C92h18NK3d1uV
ySsFDpybMUVcyBi8tYt6/W4ZsbMjgmWHwqtDiaeYhRm0pIiuZT7x2+jbtciJ
Mt9a6xZLaWhucaRyiQnmAgpzg7pCKQX+chcmoG2TGfybrepNnvaUtCOkMFb0
lVkrBNTsXbcUNO7LENbjWuXq1wP/b+q5L7ytDnD4HrjKyBiWShOpyM5iAiAw
romqGXX3/vDPbQ+uGbRrVwXdK4E8Hh+9JDLacdCHsqYRK+JqWPD3nhp5Nt8f
CKME3KDgx7AdxqOqZiBqmpzoGsfnoKvS/3jmhyaXhgRzSFEZDMBqblUYmOI4
CVehsloiagHx5ERBUHHXZ2DdmmimYTLrWHiZITp+c3j7dCOjpVv1+iJlnWCE
QOAbDUeQCKbLbro+OFXyBIXLBDanT+df12pfAhw6Xu+21qxuz49mAu0q4R/K
CF9MPLDraNgLPrvVkKJXmN9H+Erhft81GiJI1Y3mO+tX5KHVUavHypgX10YE
0xBqSW/4v/cDXcX/ODD5pjpSk743F3UARzXPHmxvWzTjRL1vVr08byyxTcvV
lpMXZyqKVup3mDQQ5ea5r3mD5WjFMqgFW8LgtTLjI1Ngly6r7j8I5b+X/Rp8
xGh96kVPiBNfoEP/NPCxl3DxgpDpIJBatoc0ycygUlRhfIVMJg6T7oateL5/
Mhv8P6zIpKkD4IhvVctATVlKRIQuHtqlqdi9PJWQcoqJbX98e15NU1Zi/iZb
4nxHoXgYutJ/QWEacPL9uFWDrPElG+jJI4RPXWFDEaMK7tc/ZIDFL7+REmLZ
KA2u4M3q81cIcfpXIEpsxKgVFpzxgmOH6woRfW3DdongLtB7xkjKuu9SLRXq
za8ON5jqcNtnQsGMlPBQ8nsg4B+ShOzC2YzKDnjxEAGfIm4w3IIsXnBaMdKd
HfzHRKAIVo7ITY2tvcYhps1C7gTqElRg5nVddW6Zpwxn2Nv0JaMY2bT4vFeC
jD+6Fvku0VXF5Muyq5zvRCHGFq0rfGY0/75Drk02xZkXtaj3VNuC97i8kfbi
tOLmkoceLuzx2iUWR3KwMwUVZq4qy0cfj/hZD6KPvwgLiq5lRWtcmxa7ypHn
/RFIlHctyEhi7igZFD/Ijxfu4sPKM73TpaGywYftW25pdlGCaMuVxv+RwQgG
p+s3hzmEeVJTkLE3x7HbYzMOL6xfBT+z3sgM3fKTjf229gR2AuzWfawU1HtV
I2RZo8zB4GReAlYogm/snG0XVZ1ActzD91UXjRTs+m4uDit796ocC6yTrCYP
mJVrRsVXzUZeuTawNl32eHf+CaNheqsd9weP5OV7/5JjQaEtCebYMT0tU9nQ
gA3lYwNT1IH+rs0piKeMHX/aqOryo5tBirLMs+UzGZdTqf4/mcg2Cb3nZNI5
KosDB3dPl/nkE0QKvv6yhwP4U2ONVZWuDnxrmJffrEp0oU3PirrhS6M9l1rI
lNqXw6oWdMEKJ+3eerv6XWU48MWtXGghYUmH7pCBcGn4ItuW6osEfR8VgYvt
DLF4NPKtK4DNz0mDPZeQ5HFj/T4hNnIoeuqEm5PTPleNoRaBpV/HBN4cAeMr
0raEdvj8ftaCzuxAHVhNSG86KWeYj+Pvv4xDaY46IislAtvNop41tZbFTnQQ
lmDtjwZzErH9QULHsJWVg0iVQcxZfUlOcbe2KqtHzo5useywdYGUQAUcZc1H
dQZ9zrX8wHKO2Mz4N/s2OAxmGAGQQPupZHU71/S6V+ngimCgmJgV+xZ/CkBw
aNY0UXtrkesVJYYF+7okiBoWY3qt5rcm+nwW2jaBdGQkWhvdFubkc1k2G6f8
kw59Cw+KCs9nL7BgN5WE+yFYdXbAZ8fIx5uJDvzNtgpiwgpWs3Q9jx7aBtSO
JIL8zHl51kvaWFVQ0StfHcPyZselw3Hq921a82xWmJj1cdK7IL7XbUz3FW0C
8vLU1vo2DFnzeADc/w20CXvFKs0evY1uHOAas2NnLpGwUwWac5I3zTgmVYbZ
TKp8yKW/S6XvEGKFoxZ33IyLfE8rABQY7oeffr0+cRjYb57uJHGXeRKPGWUK
c4Roa1S8lQ1gRB78T7Qn736ADaMnyExtMQq+HSClWnrFoDo+LPtHVcSZ9hVf
94jahXvsV0fzXzvsMLiACitF8J8WirQelZFPOqvZsiVPe3kGLSdeZbnsOtKj
G10kvTLIm+CG1t5mD4yHx6M1/81AvxEsEboQZ4UUfAe6IdNx+mbnIDX5Q0si
vkgATyoIxan5TQvzpgpICD40cLuOrqU2D7gTROYNIbbCzdM5x4bnSlb2i9eJ
oQUYIDTSKt8tq1+tW9yw2AvGZ5hin2CbZBXiCk/o8O/YHd8wAR3lUMKT0gVU
7/+xdju63+HtM+09cIoNIUr09o0q17Nzm0ydodlFwghwtBO7yRA6Wokh1X3Y
b4Ie6voZvu2uLtG1Wk+B7iheUQ0dqA/jdy35c6VlabKh9mmhkfK960eoQezB
XQ9cYI0f3azcAoJjQBWGtB1mNmyZ1SngTwSl2GzmacJ+FbxkfLCpTzATtuoJ
Fy9tvAPgnxjoLzwz8KKKG0tr+nw07JzHFJ5BuNGzBJXzkZn5bfhvgzZcCiYK
Kef0PoRxka+RWgJpnnS5CTmDJr5cljyLnSAd3c6MghuIWu6Ntfq3VtqDxRX6
dv90i3e1M+/r65uSXKFFy21AfgxuwYV1mNyYSSX5Der1SGKdJ2ddyFfdoExj
UDHhnqVfhNit4SopRkfyNjYhVN7URfojMToWGFlwduBjNbOrFKLWLJvQhBfA
v//Cwa9Lm0PcPM2l1rdpDILl4B09smGX9YIC+Un7HAs/w2Ot6qlzLtFf4nfo
RsJzoepjEdoT1Cgr3h33UsMQzBvvmQ1I8YGfEkYXuctuizz73q1dMiBKtPJp
kK+U4mPQUZicOkGugaqfCoZeqJti9iiOdzLnIpFXyWJrpARwF4m15gF0U6ok
KtoyGvdm/3c2CQEs+UOcNeSTXmSHve1ZuQ74Kp0GNRNuDPFFhsoDKd8hXfVp
dyuCYT6qMljbzsoFa7B5tVFfD1p0DQjDgD7fU7SRGdRIUJ+shA5gscaIKUFc
g2uFkturxlzq3uVz3tWYsdUX8+ekmK3w+wu6MVHjzhiATxN34L54erEV6ktr
ARqh1wTYfZMfEpU5dCZ0mHux15HZmuSbWqr3tSdjitoV8Ffkfd9QyE44nWw0
oxWX4l7OrcJSI+5sHPlOLjMMiyuqGHVWGQj4Y1CNxqZgM8XbvIxvuqIriRax
B8SVQ8p1M3iLlvNiEOyWmal3zl2Be+/5R7secOP2FL/O6y9STTC4XuFLqRKR
VFFN1gvJEx7aj60nZqBpfuOpX4hILOvnT/jueVCYMJg+OSSpbXpijRdxNGyw
lhQLOZuUA7OJSxNzXJyK9fQgrvlBm7F6jZLMp9ygDryznyefdUTm1kLDEury
Oefil4Sx7t/ge0smjXl1K7L+9QK6cIyNy6p4TmESgnAvP0GoxMKoP7AnS50q
Y0BCrudAD4l73eSYvlEgKOKPXPDRfViGO+8njFWAQqwOc0ZT5ogcKQEmRqUK
qiDvzJyuDKF2jRpG1xNJoPOkGvHhXvYQKke+QjzFDsk4ZQsayS3EpZYNmijt
aik0kvWCAkJeGRadAzfPsfQjHlWlgvSkQ7AujggV0Ws9IvlxYB3o0aZ1bykP
zTJ4vEPXcClza5k7eGvVJfWncmvwcNX7jRK4PM5hOKDQM8k0bSuD99COypQp
fbp1ZItSsqVFwJ4t73hzvll8hHJ707XXVIJeJMExGLyDZ6zTecyQEZ0N3DZS
Szcj82ncJSxK8let+LFVYBS1aB6ZsDIwz95Aq8d68TLr7BWGRhcjpfytC84o
xzWzm3qRXWho1wZKsbVNMV2o7m5OACGXM2EDfKR1UUhLdDOgSZmLk+0JzLem
BqXg7IIoyZjAqW4qiJVYj28cCgL1dzrMkJ970koHLHi1ngolka6EWk1NS8tO
CG0w8iWHXadMZAIRdYpF5+YxtxVu7IOHHk1J+UXRX8ooH9cjSdjbtpf6/6JB
X2n3Cw2nMkTVHNP/soclsQsG7QEl3qvzFKjfJd2fzhggAwI0wbsfG14nxkLj
gGwbOUN9BL2JxCkiEkPl1cfJRGp3c8bXq9iY/CZSXKKX/pcx8q73Fqi3zViF
sWcl+HmS4HM6ETssJiotMsOMLGqyNyDnMBZUr9PoTf6AMx7xRjOB/DL3KXLS
AltGjyiPwhfPuuuy1ISQ50tAk0PvHX3C8B5QhR035lghearp0Ks9q0dNQoRF
zO11lvEWBu+XhASPLoXXqymx5a4QBWj0J7XZjstomH9KZJZUvN+eLm5spfP/
WyJ/Stfy80+QDBJAS6FKxftFmETfuKiR11EOA+jY7Dgnj/0+kbTo3wlX3t6O
81glFfLKwXmglGUv8IFuveaK4kTU4UZykK3bnWgfPi0OhGyKW1qdp3T3zwbA
ggraJw8XTTmUmIzOLYu7ZWuDt9JSxA+gGZxsvIIEK3peBj4AbOxHc/IWjoua
qTFmFqjxokwO6xwx/3sJMsN6vcp6r6Ct4tgtQMzPr1yAmafSPhBO4TrvQB4Q
BMslsYXrxMUhI4/djcwkC5v0QfmNMRi5Tq+/HjTntfKrRz5Cab7NFoBvQyQM
AqWR61H5EGayFhv7t2t7Ducu+jeeX5Kr+8FSGpt146OBz63spkPtZ5HgjYbv
0TY6dqLg2sZjxSCe9G0nsU7neB3fW2DhT9SCm+4bH5pj3xjB8YjYAvWfgL4A
/zuLAMSK9rrNn5oBXmcHgXHrhnX3d+ndsbw1NvK2HqooQohOPADXEwoDQEVW
yAIanLc6Mw5S75q5VGumx11gP3FNsUz3iOfqpj9ub/2AMPO9QMDfJdsOT/YG
FTqdK2uq7bnx54CIBJl669TqrEwKwP1VYRHCJm6HBANbQNJFFEBgjFnnV8i8
6VZBw/T323efq5fyYtiCpXhu6UXc37NJGVQ9Rot5CYWRoPwxhq/1de1EesCq
RRCxBUE1dEHh7cYU7vaKErKihvPhPD1qV2R3JkpSMYbIPyy9197xowfjCStG
Ai+zdowUNb4meYg4sPo71EXoIpt5QSRAgQla5i4k0Q2pROjOABYzqZ6M7A9q
9juQpVyZR6zQ70E1W9+0GvUGBS8B4M39CGiqMDRzo+kwqVR7KzycrI6vBtCA
Fqp/OvZB7fKKmkSeuRqfOQmD/uzMS/gc33yGKTurEJpH+hkavEWGZrufAoxK
uJiSso5TJYcbRlCYdLj1VEcBrmXUwATKYh0V1iAHL8ICLeOCWOJNIgkvuOlW
lp0Llg786anP1umMC5SPHUC3+LyrHZPhIJ6Tp8s0Z0xYyIo0UtAIC4foCoBW
Er++OaZaX3EogYFmLhWbk37W4uQ6y/5Rw3FVaH+0DsC9vj0sQdYfaIJdoKJC
hKvREjVtb12zN3Pr6mkuqshXOJpjsorSuQxt76c3wZlzReVke4KILntIrwYU
eesMyorJf3gLv8Nkl+WYT60y9d0PAXt4uSgF+VZiOs9I754ih9FqH9JQcMIr
F0iw4xziELBKqFQ+erfdr1Y1nkq0JwBKvA15p0bw+c20zjrKC8Lgmsc2Xfnt
OdtNiLkUaYWr7ESDRfL8BJfB76cLxNFEWeq3DDK/F7uRRHQzFLqJDGLEY8mx
ia1CwwzWUVVyONa99RHTxX1/6JpM+ttB5wOsdo7QA17eGtXWSeXnMXRpWdOy
9W1b7MpPfWQWM8D1Ch8bPO5RPes70G3jklait6367RHW9ur2EWXvhoGyXdmJ
6tF81UQeE7A5m1TUfD7JEQdLK/XXAITZtY43n+lXMmBfZkHfOxC/SBETWscG
XgkdS2KIfJJM53JOWKUeKnYuOQeIejgQgYuasyTNEZm5jUdGBdaIAGY3ZBfR
UNBA6uJkoigFB7zjRq0mz8quEYEYVFXHy50SQUjmuhPiSnUg0LjxEoIkAHbJ
ABdN67nlranBZL8Ra1sDJ1aS+lnPjfjd92lcR+e2jRQwbplKjFFUa3G0LFre
Gv2HGJI2rVm1xmGvjlqlOZmzpaybCR+qsvg1BYYY64a25HRBcjeySWN8NT10
4KfEwp0fY+MzeZfP+iqwzerZoooPDpMR780OxCXyGS7bZNe+BSGZsGkQkiae
2s5gdj0yi5xnB4Do4PG+LKOOrmIHXfRzuN+UGJwlh59DnFP80b2D4eFcftxh
UN68QnAQRHrJS978QvaDevqZixmY+XbBZ2kX1ixW6dFSbMt65ttSgkrCzOqM
e/bQ8LYsVeO0YLYJMdgT6e4hQd+1j4lHznlRt240PTbsQqboj9vVWfbwtTEb
YrqJ+pRvwJ7zXSiEieXne1o0331qJzBJtHNfHmgpSeG4gDyFfAUQOxFD5+9w
IOTZEeEvusQYC6ravCE75RAGFNrsdd5AVD2gr2mZEwhico61sIUhcA7squed
F/gt2N3fDvFSUBHMFTwHCyTYGhItOl3ZGn1Ug/VDwhjK0xyesX5tPQ01e0Qs
EhBG5pk2YeovywuE12VNrH9il/whU6qUTmxb7yqMfXSzDrb9tYzobDeDGuar
QGZX9LOc3mLLwdIG10zn8KrKs3cxhFm2OfP7eOtkY9pqphtekfVQcH8WN2dl
N4fyVbS3prnUq7uzjU9u4fgNBHg7RJ+AZBNPDjgSnZXvMujB6T3fL2UEOUmJ
2aGzv8fJ4J3fzZ9JHV8JC/tLE9RfPw0m3CAuspfcaM7i8vYCSQS8IpbOZ4yt
0kJc89Jzex1qNbSicuTyG9vn6OO3BBlWZl7Wz8ohUkxnd041FCjWDdKP2/Ri
64hOgL/E7SfhabQcOPn1l0Bn4S4W3PJLLwq9qYbhk8saLoxBFdIZ8M9DQDtW
NMpuVDFfVnGk60XDdcA8ReZWt2wOP/dc//dtBr/9BLcgSQQ0JPyZyg8ZP033
DY9kJzoqduitVcwMYcljMnuevWUw47K9t3x4mpLHVn9wjmf7chpEX6wohJIW
82KYAxplQJzGOSjAvp1bfbs0c3BowVQqfEWnGoQPxQh82Ao4E761dpcOef+w
g0if6JLrr9PDMdkkK+9KEGsRbRfvbd4eSSqkg4t9/h1YGXIbWXpVwkoOyIO/
gzH2HAnP0HjBT0OoebIiIrTixRh8i+OPiFfaNz2jRzOXSolWeuIxmX5/tFXZ
BU4/u5hzwb2g2r3mZ/Tqt7IaKq5W22ePXl21jZ+iT96kB2YAM1iwK920aMxZ
rnyJo1RyKiKMcwx8cO2MTBdyPIsBjeHsHuouQN45zxMpUlUVCgHm5tUxB9T8
qj3GnPZ3+u1ARGMMhGhkiXWBVgAeWRMEqihK0jV1T43tVV+DQP3c5eVmOI1n
u0u9KNfr/ryoNDe9WsNQxZAGRWTbWn/zyY+Nfi5KvBDUAiJ2n+FdR0MCsQcD
7eLmk5nHP+VeQp/5CTcwyeHnj00hQZetzaWC+sXrl0ihT5lRysKr4GH6lp+h
dVqiRaWn0ZzD2F3Smeg8tmzf0mHBcvbRWgj9R+WJ6cB/thKJS9l2XT4k94f8
4zVKMV31qbcSpZ6nbu889AS23deaNOQwnXgjw8GMBQcYtR+z8c9qlqvWFkOX
2EgKYUKUv4aP7bT7nGKTG1AxuyK0Ey4QAV6q1n57gH9/pbUQ3E6ztHa/ydJx
VHt+4JIAcooOAzCcjIOjzQysl/ncA5gOPvLwvC3ZfRtPOiSafZBhneTTgChX
5csNz3um4lTvlZRRV/JEBSAL72JZrz6EQoGM6RLnHUMYHG2r0Ey9nM74U/Lz
pgJtIDTpnChFs2yiNBej15sEx0oX+/vrV3FdECrzU5eqTbiBDOgS+wNw/H3Y
hSExlyUmlxViIQUt1697j5zk5PptxRmM43jhi3M1zgtPNYcX/iO9oL6iRj1a
RAHgjoREKNkCOjtEBFIzz9/4s9kwZhBcZkFwlURa3VlAo8ujbExmchgies5j
7ccx3zN0vurrpC9+NdDPgE8m/i+2CG1jRoNTrjXl+HvHemgetAFG1Axw7oad
3RM34eCKlFfV5SFnOgfPLxngR4G8S4Sg0/IOk5OSnzTAr2PgTTwFVYKsfaRQ
vJ+4uiMKUgR4kpqym6oaVatmN6pzHEe1Cat3tfLQs8/i+jS7Wcvy80GGmuZN
XHOMuDzOkmBvWIkpwUYSCKDA/FGyz3jL6f/X2xXHt0kuBsd7I2bbT0WuMfEo
vR4echhWHmR7GucvyJjqoW341bSr09CaFZ1/qs5KC/Ck6RZHy3+rHr0YaVhh
IPwrsPWhLWWlTKjai/SJySNHAhYEqRkt//qVNiaeOZTWoq3Q2/IKaON699UP
0pdvc0WHD87+EmvjLNWmMIduvmBheb0+IXcjXF7LKvi5lK11ktsxRJes5EmJ
BjnGRNPq0hajW9xfStkENha/jW0SjXwG5TJ8zLN2Hcf0sLpNMgoehDyBCUaO
PJ6Xtpaiqamm++4CudOldbyunBlz5Fr4sD2BiIruroEK7sHauTebxC8SZQRV
j8itGCu6EvUGKb4uPpPQ5E1jqG8w0oL1IOQ6SOnjHw+d6nLtk+7z/yiZ+uEW
/1Xb1qS4JvYZKlX7GEApkBjIfuagV+w/4fBY9w4FsVvH2wsPKK+Yb2R7GjP9
qRLfl/qurF6elupbxGRs7ocW9Z2cpBjsqy4ivz6MaACut2wTjxNLU/t1qrGG
iany3b6R87+lnCMcnoZmHHZuELO+GyKMkhwPkAZ1DgzP2Oqw+7f97/i1UoxK
2+bFoIXSBHZxykTxuIQD49/SSNpIBsOYVRfG6J5V/IRNmogyETWgoE8gpUnQ
bVG+mZzZTHBRzQu6tmTFu2NSht/RVjLxx5Pgy2e3maDPVJ5YH8Ljc6KZ4akn
nSt/QGR6JZW68ebr/XzPfs2S54tGc1bRGds0FtNQX73zkZ5X5Hwbg3I9PD57
Vr5c9UED24TSXCWYEjF8qIbqWSjIziOE8ZjxdNofJf0MebmK5Z63kpwLgQQe
ucgd+QaOZJ/VulFrvfJ3QZa1rJFKb+TwNcX7S8iJjWHmqLL6AnQBBE4lUVLr
yzsJ7Z9F/6h5/GcvLJuO53Ir2Bo9ROggCGf/EuST15tN4YIjmlnvjlE7w69Q
8AcT/WXOCw94Bq/XR6nIxuFlxtstRhI7DDS32OI5IVw2ylogDeLcvBE+xQgA
nm+apBj7GtUks0NsMN0F/XY2wHC30ftxG5PBZLQwb0MU3LZ475a4JMln3mNQ
km/GX1e0L0TyThHLp99O076oxDcpIq/iwQrPNquqxoppcbx4GEUZUqeb0ZNA
x0DHhO7tU/674FyskTzKs9bGZHO2tqHmkBvL0DFD9jgb+MzyEDXd8wc5XRLv
Zj567GBSnZMQ7uvGn+33q/pqAAAE9sM+DVlXeI+6AN+LpoRMZG9sPegCRfI4
oWLH7SBAlroCMvT2ga+ZyfZ+ey763K+gjNb1Jk9VVKlUfhi8OwFfwsDHlT13
jhxAsh5GXwJl57/UfE1SJsaF1EOatsdMizEJoWELBfH/mYqnP929MYZZJIkb
oTzIEnlcnkSYFcrRhbf/IsPy/PGOW7y6DhZ375GXNU8XZrDl0jcJmDT5ZJJT
1uKfSZnbhQZAosHk3Ym01HQGczGPu8fQ/U/F/xHRGo31I7LrHs4bBMwSCUii
dzVQrZVFSEfDDSYRHBQOpMOaudvFAxYMrlHSAHwAEIaNXc7HQr7I2k05RxdE
RQTqJZPcwzcCcuyte3Z+D3mauTYW4Q7KiAeC9O2jYfRXOY6l7wD6bTH7s09W
Sirs1RRWUYWvE4+xYU6iywiFJVhozJaPGzBmtDM1wfEPKXIX+hlgOStj8hcJ
PLAA58QckWEueuWlGq5G7Kq3xu4uGK0++9EXiMUKr4vkDHttpzmPzikfzO74
7FI7hw4aevYD9uJhzMfdbxnhHr9T5ZfWaGviVHFwexgFH+hK1OCaFbk5jplB
gGD5yse8Y1mrTX+TZPn9mW9ldNo4MF8sUpw33+mqEsdvMldsffrjev1kgutD
gp7fSkbncplGvVlL5t8zJ8zbnuL8G/+mQMU7Rs8sclL3JjdVAhxKVlt3C6p/
nTAQFjHdYzxC5C3i6StebpeOQAw2Buvb71sTSkhFU51bNbYv86FJh9LNFB32
/b0T7CHkc0hWFJuRs0Bhpp9U4EXecEyRRuMZxAmgRZAHYdX2lNYDtgtFgW2t
T5psio06mGofRmRu/wvofGXGMSAbWjvkrxMRhN4wGs5osoabuxT8qPLYcRAD
WdTmdpaTIvnZSU5msf2QSHfYbjbTrbFcyVnLWDLHR4LBQ0Jv9zBxnfHZdfCk
ZLHmP9R+uDvwtj3U8Y/I93RXdpuD805z8aPLoz0r3W1c/IER7CA1WDsDSEJ4
nY0lV+30GaIBKZACPcd9R7yK3NcQ0quqVXltprdSN5VI1tFE2Q3cYvLve61y
u7ySYEYCyx0ckfdWl50Jn9TaeUxNzC1xz2Mxg80iqPUdHrDXcee19NlEYzVN
PIrl5FcJjVm7q+XfKJGswzbttYasVe2yWdiQFXFaiAOWkxY3loiUuKZgBMjH
4X3ziiewY33/eIFQT7krcTPVLhFzA+CAywDCsOBP/N/8NOcJgW6yYOSV+SFD
5cIVHxoc+d6cAEewxIXS/9Yt7YmGPIY3poAW34+YJVTthQDJBl/MxvDnvwzA
AW0SZA+dIq7AbOLQkVQtZ+XHFYuyc7O4wfAxU538q6MXrzJl8YZYTN/3Gwki
jFyd4zXTnR3Wgowxugm0IwzgrGgeQkVs30+7en++jFljWYbzWdrt+J0j5cgB
alZoXUtyfX0Y864pobquofJRqPg3mYiD/orAogOIR6J/fx9Fg8KAgx3shppw
hMO/IIh7jlOfbDAptGfvXJc4zv1mtqk27l3G2M7Zyj3FVlOLER10VDuJK7cq
x6pvDyiaCRoOLvuoTpiiE/z+mIcXnw7K6QzaxA/FglrRTMHe4EjKrQMRlysz
MOXvtSIIL6d8/N7AHA2rT6d8WN778RoxvDqdoaa+QdgthhtzrNC4RMR95eEO
A8C60bjY77615rHEZ52aKELQEuk8dpLm0z4pldLUdH8rxVEn/CtFME43O/b8
V8V09MhTzH8yVSiTUaTxkGGpm+h8Pmhun39b5plX9yj1ixTXKxJ5MS57szUw
8jRYdy+8bDMaq78LDSGCd1mHpW1+YwrYIpBnH8KBvcXnbNaFq5eFgpSf+/bw
Jn69oHYyP4YvVOhTn51olOhAlXPwNEqvooo7VSX0TRFh8RPThc/SRk8iowtu
aLzxvPTbCjSYfQeLiE0xatrNPb1QyAGk3/cj82tM4obVRKYxt5knscLPACjG
N+jcicolDpuYos5q69C98fX1i8so7DUfGJfz2ch+VMdmzFvdNhEQU4mAKS9o
WsX38FqJgqz5DRIhKnmBt4BiRxmgu5j+bo087hdwBpUzFvwU6xFVs8E4MUa0
r98zsQRJ4waTToZ4Eb+sYyK7EQOU5s+qpk1GFlw2Z22NefBHFUF//+y4R7gl
DnUQsy4GDagoYWbZQ/JDKn74EfiYFfRWzTO0rMxELbh6QfQKGhaRT12i3gzX
UcU/OM49Bl8mPvmc5d6yJgoB5VwbsmkCxINGYZuhMBhQ/GfM/VEcaDi+yFPR
HZkBehYGwUktccLp703gENzFw+2/25pNPLOj8sozDLgjz1b6/4pBX2x+deHv
NS6ndYu4BOjM+NLzJDNzceJRyKz2ig2+ec2rm8l1EOIynSxU/feWdx5RBh57
JKp/jqdJemG6EIEuKIHskkksFx0sz0saopXOYTP7BXFhYdAoEZgJ7/rCkv8u
3IZFyogohjHI+Qka77FagaUACuNQo+VffW661FCK9D6K1igGs9QMJw2Hoxuf
CovDSOmvT6hvZzUrNLlhuU/GS8vjzlde1zCoopNaS/FNK2wkkuLE2JDC751H
OcqL56vW965+7FeXcBSKaXcJm6NJMfqeRRq9Gk4DT4uS2xIoTTIDKsoYo9tB
LnWB1J20vGTdm9e2+tBHgTG/TDMxNB55j0iSy+TY/NmYyCBsm6OUE4cQsxwf
J8qHtnqWxrXok9y5uaXWsNQsRJSY7apFaBIG1ciGOgoDxtMh3Ewi1xdkiqgS
7Klvezqa4oU9oJyRQhEGyfOL75lden9YVr3o1XlLwsYI1skvZTenYg9E5eNB
CzNiA7RgomJcVjCRUa5h2l+/fFZYNTImKjHFZNWrqKQ3JNgaDjWvLRgN+mzB
swMqrI0UdM4iIgnsoALKgkEqqUG/UtAdcnk+m22xhGvGTsH38CLGtfi1S6ud
Zf/2xu6ULx32LK4JVL8cIucV8aIs0XHV2pJZICT1gdOwrAFwyEg9uJIKPGDf
HYP2mQT+/zeUHeyka79Vmclg8I6/tjjZ9Gj75bQhackMx84BHGWr8roPe0eA
ZPUSRkgl3Ee8py06eDjIsxH6xS42ucqhjPYrk9mzCowljpFsBK1EBAqtOIS1
gMvud173Jo5/cT9cR/8OyXthU3XTr0Z8rt1EFlrGuDlpYjDIGjgYgnv0HkyM
CBSjv1cL5ix0glGbzkeqKfRRINqrkOcXDsyJ6XGpGIM3lFtOhxUdsyDllhGA
hWphrIazScg6AWl8gmSJNzQrrfbiFGniqw9WtOY3F37lKAphuteJF962aHtW
HKH7L/HIvouxNlDrq+zClSjWBSsduznRUuAB92hTQ2C/e0ZGMc4l2nywZetj
F34CtLIoLMTXFExc5t0m6FfHEl2meDVw96K3Pqq4hUqFBf/v6K5oSf5t4M45
WInDnoL3jQwEiwvZLR7uHNGdgldvElFI4iqnUb1vB5wl9ZI3dIfoJ7BFRJ+3
KXjm4gN0NXzc0DqUvDVf26SgyY93o37ivpdw55m/egPtdDtqFiS6ikZKs/RX
l8IFHVKP7mLHlVuqQmANVw5IHXCw14X4vm7duP10hg92dzkYRSf5LPxLAmWB
zBQDQrlOaY1BjY1lm7bCduC4o9tho3eY+40ewQs9++QHVQ0B02/gbbApQTtE
1OANYIoXXoZMrJta0ALkwy10g70TibMUvrleJywRw/A7TdiM3AsMZt4VKm1J
UB5bWYIpn6CRiYJt1oQHvWBHdqeBTU/zUU11t04x8MjILOHIYsWqBFKSU4NS
3W0xy8bTeeoqS4+BuZpdNQjCz7zslYKBP1/sA53UL1igWGZ0jd2hLB+to7c5
iGV4BD9DHsSIAOX6h0TeIqusip6d61mTNeZW4qgMrz2pGRaAnWrCMZ6DPPWh
9qo/lPLGnpqlcHQ08dKdkOGfRQf2dh/dCwd5bn5C3PeHLHws1weSn+xuCEtk
sjO3dg2ZympJ76zY7zgmIMtt+EsukO+nNFTfiYdLnhlzuoU2yHKgdqhdGydN
qB++Z8CSGwn+tjWGeBtQ7O1I0A5COrr63WEIbDXxfagE0lVxzJmJTHmRCMpm
yCzEAuzW7D+KoSGacpB/Yy5V7nuPImtzUvPOojgAT+ROREOimULkBmy8jdyL
IcHc9HcAUPPK1YxvzMK8caRIXKOo17NIFVQwkW393bTDNFbyJ8dMBqFHtSep
mgwEb6R48ExoWdAUZyV17yEuJ1hvelgo7URCpz+DHz/VdDfKjNwXHiAWIgdw
vMcK2e/E08tKsXWCIRYu5KaK2Ikxd3Dcgq9nI7sgol1lJJl07Mjx4Y5VOokt
kKxK/PtUsQd4HS66vvfEX0RJnz43HwRueTIlT0D8frKOGGE3jbk7eM4eZuUS
KSa46GrzLSzmNV7/gT9AZXLegMSG7yPCXCgXXrOkC8OiTh4UIUy4TkKQKGe/
kXlxvBXZHGxlgx/v2R3xQs1sAWLGPJrIgskx76cOjqJ/Cw7Vz++Ft4jd1RO/
44s4Xf148Fq3aW4BGpsfnUEN0csWr5tYegiyl9PSpcv2XMnKaihFLtdXLSYE
fWZJBTrztrtSCoeb6qCesmBBfZIXVw3OZIUC69hofwFA4jaeSJEfxRJdP4BC
hmLcKOiLBcn7YnED1T2CrFDSOjpwT05BPtoF3/Kdp3S9hOb0HVugz0bBGTte
072YEoBjlnfZd4ZUQ88Uy6M9C5Vf9bVAKJP6t7OsaH9WJqV1aInJJ1Y416t5
2mXQmmmAAMlR8Tk4oMlVbbW0HU+V6nfQ3v4FHIFDbcsvBk3RVuIj6ixZhekW
aIp5Vqin8ilhoJsl9NJgZqtTBLJZSbI4LwrAYi/g1OswHUZitG2fuPqD/IhN
RMA4TgVXO2I0QymE5HM6d+cUekZbVBJbQ5X+sMlUhHr1tALuuNP32LijSuwv
8kWRpXtMSRidSnOjtIU3P1nuBHzIcpXCam0y3BrQGYzib3DZZLVBWHm4DO/Y
XeBwt0cnaRWuKfujbYSNdAlAaPR1K4a5KaEgl2EOO2wEQSn6bz7JjXhgLeF0
ai9wn+3I3bZ6UHcOHLR685/iuf40Prer6z9sqn5Jl6yMbC9kCEu3GYFR/WBM
A66q6TBXjYoWGgLFZzXoMftl14daC6E0zUSyl0IWFmMH91aHlRP4uym9Tr4Y
A+o6z76E2Y67X8hRP3xYOHkcPd9Iw16TaoOZ/TV87c9DQu1K03sMZxVlGoET
pCEW75dFT1rO7Xe3xMxMQdqRjNa8BWqbKbH74/xiX0BYPzv8W5XjKCspztpo
iuRNIBBsXn73YHb6T3iux7XPmr5pjE9aCTgWeDfz7sYOBr1GJ62g81o6Z4wu
Kg/DEng1QbLDKflFwdu5nxoXo/9rnmTthrTRNpDgirmvraePgwgaPh0vZjSt
m964FbUDQJx8pkz4FgcL3E/6XUux3K/q3gXiW9FR6qXkeJocyTzLRt+nO/Oa
GbhjKWkyIwdhRVGN/VPCZvgiBAfHlnvIs3LmXI9hRo6jdwk4RHI1tBui5g+S
qMcB+Kml01zuKTbZFmczk9jhEqlTCoxQrslV8F629RNqTDFlLPqVzAnyVTDj
ht0JIbHIC3BEZyrtEzQ328n2EJM30JyyTY1LMb6TdO+xbdEmqX6n0pvizeaI
gbQdqdh+eb69/h2caguH1QvxIbNSxfaXeGRAFaAKxKG2vA5vwxOugt0Vmavp
Z8EeH6tkuJ8xuR2glx8Ti1TKuEvjPU/Q78wlQEx1E12zaedVF+GYGTsMGs8d
IZGumPdVzFQuLn8nQg/vODAlP4T7SNNcWzC6VxDR4S+A50kwm/zqFIKaU/CM
StIlowTCAD3EP0OJrUe7vHmStnT0Ts6ivodq2tOfEAYW1gD8/iudYprzv2T+
PSbMHj1rDBDxdDcB7y9C/4Rg922Z27kye5baHtRc7muQ0l2vbmOdUt6hVKyC
1Y3dY264IlR43Ydpaa1OnM9K+DynizK3cBmsoCxgVqsi66imL9wVUQvzPLE4
1InfQCTDd8n92n/XQuqlkt66RCVZitG02AgIsOkmHh53SXsqbWmQxGpkHnB9
ZflFjol0ECjlcwsp+IN3RqHh543fd+xpqgrLWosQ7XfqsrQoS52peLc0VnBO
0+ZhDVGeIP5kLJp9mlkr0fTVas9Q4+iUbjWoIvwc/+snSyJeqM/nHxgfGQsB
nFZs865Tzuuy49l9fa6cf+W+cxvAVunO5Ye7bAe1LHGQ50TXEDYO5FaPdmxf
as7uSvhancVCGr1zrGjNm/T7Ti8MUaN9TQduQc/vc2dOrUvIXULlu+cwm8td
fPjmd5FtTgR37vbTsAf7Omc9sxTOTK8UYuA0JKxTxXIYeyRD41to/qRHP6Vx
mqOeMYO2XDi0pbFyP+iyHE/MbQszjAHThQoyepmIvjHeTsRID1JVgZWYr/Nh
vDsVQN9OBfFj4O84um49v/0bO6TdBJknJvNMNFWFEzr8z2d2dngPdrC9+Slq
vrbw3PuILELjhZcifjSe7mpgsgIk2k/eaJuiAG6J2ZE4YPicUpVKATtda7F0
E0K4vfPTlukD1oHTpfvEHS8/jcpLtzLngVeYunsjiKoVLZhtiwnmsG9+0cUO
197owKEWNpDvILWLZtOXDTKA1uG/4FPGSk7HMrliVToCcxdSGEtW6X36mzzj
DMoY1QwURbsVfqROxtsw4yeDqET7Z1SwwbpomnofUgbcixcTaUvN8qlZt7wJ
X0QsEobzbK+oIsbDtHXxApP0wUoE8kAd0aBkJaxbhDJoHNICoGOkEUIPM9Vx
rOjolXN2473sWVqsMYAOAQddh39XrKXjcEsu9+B4qm9A2HaFkvcnxqOv16Oq
cixdsQL+rVWpihlZAaeQkoE5wdu0wjgB/YuSQYaQMt9f/wEj+ukuGgOYDQjL
B0ZC3hzz7l7MW8YmBUjw8ZvwXaEdx16qOjOb1ypDKRna198brbb+Q3KvQLuv
w2+KMCyuhYWANOEOReKiouTnX7/Fkcn8nv4TpboJza7U4kHlulP9iSErBzhN
vaoG9Xs7gn8Z5J8t56UbALpEm6yeofS6sMokCwxb5c1pwSlGleAv3CGWXkCb
X4Jj7ljakgOdEqLnhUiL2OODv9TRtmoFk7d5xFvaK8aKx+Lbqr3BKBLTJrl9
90nFgb9H7XS+rjI/BtyZ2eioMEHnn2HEaMdAUACEgiz7c3umMg76d8M14PRF
HqD6oAUz9EMn13SOKhQkgxYeZo53Uo+dq9SJCX5Guf/vkujpnRwzonkNXnXY
D/MwvFsy/zlpt/0qe8wZMEBKq6GbzB0dv32IkzMVunS/e9zexTDntKkhOszP
GQWIH58x/HjPHVMdny7NDKrZm0Na4DpdeMR2t8dv2RsFi88v4vu/Ft3CsZGN
3OHtk+onLgfoLY8SLF5sA4EzfxJ4CjbwMmUjSUo2N7BN6FCq1U/C1P+iSCP1
+VImw59jgm9C/vsC92iKSTnNpNB9eRAcKGiNDb1oAxoo2r12Ve1uzaelSCzm
ltAXhkDLGp8EJcuF5BEy5zorwaKlOJWcuMFhJa0ZmI9gDrym8kJlBJDmC9v3
hoBXXJd6UVulAqdK6qyJHaBBjlRM+dVFG28eFnrizv2PFASwKwF8ETDCmpWE
13AKrYMqneiqfemp7040QCKbVH6yWbXMTsrBKSg9WXzrg6+0YpCfDycTg2FB
YSWlHhPcNf/VEu9b6OWNYnZNaEC/dWgH4b8DItTiIjgUhUCXFLyUZu2YB2ns
uVFLVKEELeWY3ZtAuAuG8Y/DipdWfLbMgJBTP2HRoxi0g0LTHk+aqxjNsUqJ
LjiNy6uZErRpRfCsZleIjgFKa5Mt5drsHMTb2egQFDgUGVf7MBTEMyeCjfPE
gbZZOuZxaY314X82SB9OO+1tBr6gzXDXJiipx4G0Z4AGzMpCCrcPDH1bKh/A
SE6b1CLr/Ys/7XOaNjB+SNAk1XUdpcQzASc4p1ANhOYVw1W6lsE3vlF+7lLP
wf7GcxgZjEVLWEniAjgRsrAXZIu7JASzvA7g5MkGHGnRAOV/0Wn7J6F+87gU
Np9YfsGT3JncwFkxpa4EkUmNYjBA7kcQRvlINDJ8MiGxYPJCoJ/cwdXf/cx8
zUA8gLAKdNKWteIu5NdceGBwGvzciCjraAsecEULqtDhQ8XUtNnF5ySq+HP/
i1gwGJPuz9Up6FN1zR4hNLR/58PWKMSdlKm5WAKB5NN+5WpXq2yZlNZCrhOE
OBhg5+U57/1AdAY+puCGbG3TIIPf3tB7jWyePRffgfpnW8ZtRlwdyEU15xUh
7CzYfU6JJwoSPMoxjo0pnqGMAbBiDc5issG8WHJI6QnZcv/PWxSLzkceoEdi
biGSJ+jhB1mjJSnqklb+9Pvz+ya5fxcXO6N4HRm8Q/yGkilO3dnzWW+y7QRj
fXA2FqtYW+HihVccS4HtdZXn7wKKEoF/SDyRLZ27L2IQjH/WGEM5mouvmoHG
Pm+WJGDRVFm+ntYMMZ6EU8NYv9+EXMcK2sUGFtqys0+g8G09CCTz3Z8vN5p+
4WVhL6PobJNI59HQdhF+DMwDL4GldJ7sliLUbfO9uUgASwOhv3M5Ssw2DMDw
Kc3KaNajblE6RClahf3UPzsP/TUPlf/5eAAY2ifBW5Bdmw4K+PZW5ZOCQt4P
kk9/++RqWCyljAl67oCYs+8ds6OyMuOjUS+TCpTL0E+lM4LA8esBHFnlOFNa
7VBGl0m2ja4z9ElIXhwxIbi1yxW+corWvBhumSTgXPbVI6FoFji+4Cuw9vii
KFUtfXb8et0oC5GnjaSY70aLvE1ZnrcdZLkzceOuIWYLot3EjfavIQeef182
vlCMnLupE2HebU8W3VOIKRWO66Rm6/B9sU9bgT1Q0l8d8W6NgQ2L/o+Gs1Rg
t/wWaZd9ldlXimGvihIqFJaWpsjXwN+Wyr0nXge7c52fCBuQPvxzLSoS0iWI
jtah5+Mi7KvSqpeoVJ6xTBq40f0VPkU25mcQt4by+J8DaOzrZ9JDpw3Ny/CO
Yj8q3g51Uvc2zoAneJow3tRyp15QsgLkfNyLSwcbXMLP06K0R0OGHyf7jpwU
xiO7+9hFvhOXEX0aayccRHJG5Eb/jBLIh0UJSq1RAqeTUX1x9eilAsdZsdhx
6udcFosi9yZ5UHLY33LxuhWvZ2EbPwDPNS+nkPlLHjMKjIRlbl1cV5SQvDMw
OeBIftxw6XlCkQ4Ic+fn/WzlBC6nEZbMKO+2tXxlGtY3j8XoMgW8Gg8fEPOd
ZNlS/cLHSmZXatcHdsfs+Ih0kFAPY8QJlwlHHBc+Cbm+PIxPzJ6JVV06pShX
uFrD/h0s7i9eCT5NIIeG5w1/2+tiYLIku/SLMYS7CWXCu1s9GXuxJ8pd15/y
SPWJVB6xG2bwV3NRZlqBLrnsxAtaXUWQvVLbPfjXZQDBt4NuwumFQacOQlfh
7Nz8wHLrCYikr4y4Tuo64KlkOcMxJby+OIFz0GYUjKFySh6beVxhtAuvCjpD
1CLrpZ304qeFh/d8KC67spoMItPPNeerEfxKWH5rAI7Bz79BdPVoWpdOczKj
H08uIQITNHdwFzHaJNyyGW5E1vtcCv+B4SF8HxFfgGCdi9MhsHB6qDkAl6Xs
7JRR3I9VR049oQTA/DO/QANHO7Y41BHdFBHnLmDkxTXcEKruoyUaNPQTmHkL
Iygq+5/EbsDpXDutP3AV1Z3uT3M4AJUo2FgcDmD3HCtPtiecnfmJiswo8z6p
6pjcF4LTD1hMW1UX1QQCY165nNVySSt9ezIwhSx1PrfrFXxlEMMBULwbi00e
Me8ZjgamUSeYCu4OvExiZRk8iPdfBrL2kTxxVO2WNOKLPsO2kEP2oFhrH/ua
tBV0ZjIc8xfha+FnmYr/viyxpVkFQrVgCpVdBVmDplFOoBEe7FqXFKFSItAx
KtOra5dPWlA4LonstzM31Ly5HBQLbMibKHOpOGMeCZK3M439HGSIATykXxPN
ZlS0w0sZt7fGGdMK6sL16EHD/pqIViXwurzrMdbny1eyUITZivnXa0XngPNS
Qws3j5OzpmmnnT9wYkOyA4G3IlJREHHRpHP8YDFstjQ4VepN0bps4BJw56im
W7bSCGnF1bsvTViU28Tg8Rq1OZ0ihMJEcuy6GIu4GO7lM5/JVx12GDOf3K5Q
Up7iDr9YcQf/gxZjErJnmM+DxQDIX/bjCapefBTwnP2b+UFKGf8HjB4EcBwR
seXtpGLv7B7q2q8LW74hNibF9aWBIwhVA5ZSjdjhTxP9y2E3olQGkxhka+2R
JBBvuvXKzaF6dCGurlvDNr+icq68VN62F6v3SRfE7pwdqYl7F7DcEghCQMDZ
4nsFMhijehCFjTHdJlY7Gj0IgTwiipbGlIJtfVKUD9AlSC+3neVmeqSyiEwV
EIomv4C1MEWOt9Z0bk+Usk38a/cOcCAcQbjW5evDEz8nGyyIhrdrd1qNq10B
zxpDlxqLpdP/abC6QPKx9aF0r9+EOCSv1HVV0A6Tbnb0vVUWEjDXKtso/mAw
ZSVEPEcTQh3fBoFkBALkag3W0X1I+sjqWz+9uX/kzLQ4lfdkrZDghAjQMnxk
KH3h6QvHEYSp1/+kQ+KFn3Ys9UgzQTYTTse/nIhZxOMv4wZXZcKcaOJs0Gmz
vbGvaxOTHQJ4L5wfo3NhilxJPkWsr8Ydsxt0P79y3j3y2AdXdPmt0YTLpcrd
6nSoWmjsjTTo/THVlduLhKD8rXhY0baoCJA1fZKsZ5r1EAqqo/ybi7Y0R1jG
nUpocbSnQJoM/NUWasOgDUzXyzFAnPD2TJtJ21SrDkdqhQNFA2bwjrGmeHob
Dm71CeoshC1Z7MYwZbvUdyTwx3u1cy2vSnlFCCtr/3kYzNEAxAAe47lb+tsV
HP1qHrIMWwYLd0OTzyF4upLvyTXJvEqD6QdPEE/9tc4gFkseixQY7urPif+h
3Qf3WK5eBZof0EJQXcX8H6KSnna6kmMFxglm/lJVyDFryAJ35kYNs+IfzRRU
QiuefvUuJ4UwujgO8nY9HGmMmWQozJ8wetmVe4PGiG/M2hbVRAJcw1hvJhVR
ekDfn/lnRzYK1UMhWjQDH4DBq4QXauIziQjaKVLpipWW7nUqGDrEiqCXJ7Nv
Tj3EyGE9yjw4iVhAXssDjbvdVCpiNOiDV6LbpfuICwPw15gs/hfOYLcPuVQ+
y2xJYO2eoK4tNL714osSy/nc1Eolpctn0V81hub+OwJO0F+1EhPpE4HSVrm0
LgaMKHT40N9DwJ7DwCJmoiqHPJPkkaVmh3f/sE5sTEyHRcpzEY5FKTsX2yHR
alkIsWAqdliI3jnVHOo5xSiHEhndvfQmHbMGAFXjlmO44DC/VD636V3WxWEc
CgQTDw19/xrm7Dx5cBOQNal/Vqw45YyAB+7wVhcUYhhUjlJ8RCFH1CGb0VAi
9/w0+1Z1610C1OfZP36UPvV89PMCpK8mCu+L5oW0vs4BUq0AjUBaT98swcPm
xg/8NP9JvlSEjSZkbFphCZQmowBZ2b05Z3SFUwxj/E03pC4iqgOxp+2L2InM
W7FEDdIm0iaY9C2MEasSslqDW6ue3FLFlgD88bDNVNjKQlxMF4PD5NyEQbeZ
Ah4PdVM/ZBUImkO8r5cw47Y5dxIxsccUqsA8ONOmpgNz9grm55L8mfYUdw/j
BBPBkA/NQ07BcYv7nAFOJpl5YAr2q6GrPawgxVCMH6V2pi4MDs1qRfH9c8tH
jph1SKhF3ee5ka+6+rHbYHcY8zCHKZC0Wx2SBBYCHmLE+R65hV6QYfaji7RC
sSs12Qeskh+x63dqUvKuQ/PmGggxPoGl9ft5lFt7cmK85dperTJ5e52HnmJA
1023FS7bMJY/GpCAyUhEuxnMRrTkQnS1XspYXJx+xKblrRfA8dj1Hcwa/X/e
490NjNPhtd14U770NADYNUYn9kDZ31kXxkjgDSZky8XUIqTVpk7GgL5B2jnn
ItkP2hJZ/lVq5+i+SIeBIhQgMTjbk5Ku3v7I3jByY8t90eEqZBG/dmwzkdcC
4EWT1vXHxF/7ErcWAgyYdC7bfPXRxxZOawr/7Sm/ixIutgVhTAnuQ3F9nsta
JmAGSuQCXZ5KpkJ9ZPlk60S/0TkC0xBa1nNG8EMRFGVcyh3ONFMiaRAJV5RX
vlvQw2CExl0vAl6NMp7Nnrjg1wy4jAEZaGbx8Fiy+jZG/+Y/YnUGuIaS8Ild
ncs3/IfPJQXg0nl6OgaOcCI2XRpGzUK+tOH4Fp6dicJzXl+ZxXDOfD+tU8EP
CdVnb733V5TSxY+4gHtjt7pLhqmfVVgHQUft5svrDBA4du/To5mfjL9A5pe6
8ce8FtT2PAcg6TY44bN3GLyHznXDrupOS6va4ewkFy6hs//PUvFfZJ8fkmKA
gsmAkUmV1/xSOY3R2PcKdgjKJ82c9Ml7ec0iK7S5uhD5jllEMdZcF9gYTr1y
Tly3Eoe7zR3c+Fjs5gIG/JIrHQ/BweUqUqI7mgQUSEO2SqVEVEO32re5GVUB
TguARGzbrQREyYntDaUJbHzA7M3c7DwwR71w9gMyGEkTf3DVjdNG2PmPI8c/
ZI7VqPMvj3QG+fI42/3++nopJ1WV/ThbG7jl1sV6MaUk6P1pnwr1xiU5haID
FP3iU6HdEHY5jD3K4bqmA52R+mnqqe1F8C5WMCIvTt9gUjtsaGWKL8S1QtlB
5WRGquCxWDzk12Ymqrd6OAmYveiwT0QE65pecnAl6H3KhSKtklWaduWttnsF
nuLwngVtPKjaYhozQQT57nokSYqpJXmOg9Ew8co1WztdHTp75jpy4uhl8fzG
9lXJASUA9zNikB/isnY4yIbpykqCtExLunf9DZAf6jdvYkCEjus0qxErivQ8
iW9wtRuf60r+pxYn/tMX2njSt0CgEVKUGfS/opKn5G9drQeDHSpp6wUPqc7v
ce45vGugiVM9QqrykMuKl+SfRociL8mrSjrOuJNLot1CnXATzLHN/qrKXzOu
fCzSvMBR9mMgKhRKBcJucFhXnZIe265JXicA6QxDnCXiestOrv0+5HmyKie/
VFsqKHPp7isb9NwNpXaXG3zg+iAecFVSr3qqkjxZ0A42+p6EPLqK96jN5NTy
CXRRIGrDthqGi/LHRAKRj9ZrVmqIzb66HUPEU7zGIE4CttRu/PTxALUYdSgh
VftpRtOWPY7cKaiMUzAK/lZ2txKQw22gVs+1yFJjZsKETL/JiDX9kW/ytQYJ
/EcNHizcAJm0nYCrRc9hZTexLTd7FArRUuN1bBbu1OndLqe/TgnyemO83dGM
KmwxEbvs6jB5ASqhTqXKo8C+P+yW0ilL+QNY5C/+JRWwOzji2ja8fyE927t4
8ZfreHtiJBMGejgAj+ieFPfRbz/3sxKZ1Hwru4ZU1wV6tpj6FJbBiz4FuMu0
uNvvUGfnMGefPkd0wpIaFc7gNljMhdCNwgdhim5wD/7/GSgwfXY4GGLac5ri
f6THR+2R5g04RK8GXuIfxhGWN6H8uwC51Y+TAaJ2F2fVvdvlx96rUync/brG
sHxL96TI3tVUxCEk7sAwoLNyGevpcH5zVx1jB/c+bbMWOay8baIRIikXMZNX
S997Lo3TP4JtV6EqJ4MkryfLDCn1lmkl86i7xz1yiEMJ5/Obn5Hq0gp6dZgX
E87MegjHU5VSDD8ogmhH2/BouhfwstfLnAV5KjWxXuVqX4x1O1LlgUt6ZcLj
0P+XUWdh+AuRX/FAxpxBdeI7TY7kmfgpSVqeMm9plJHoz5/WalMspfQRxVXp
PQBpQaXfnQLDlbiFVD+Rw9AyfYxo+kleqzug//ibqsNVNOHt3nLc+QtNfpBh
dUSkpi+GHaE4a9gDnCw/F/I5LYHE5mw8Xk2ShrL/GMAf3fa+kjK2Hx42sK2W
l4g5D60Q5W80nvvpTnIZqzE7/5kbmUkHqvgAqynP5XOfCG8x0pdCFNFDBYyv
5Kgt0nndz1dw4GA276cIr6IyRtRbvZqwfYirKe1dlwNJy3yyNoh0GmdxDuUT
isFH3rsK2tmovh2TMMaOdACdq1b5YXBL42m29gSISU2uwAvKoZhkGFECIQpB
5JEKW/LtKEg23vZ8SNAyiI3omlLbRaOLM+zwpjzwg2MQGU9U1ON3BScXEynJ
ke4HvjqjAgNxWGIKZT7D/d9dn3Xxh+cdiguxbVqAminag7JU42uzVOhuyW+K
J6Zceh6rt71bfs2isSs/G0MYoAUDnrrwtlHRWaVeWrmmrClMYG2rRs5tii1U
9+fjr9/9rlKzML077fnviCErayPKIiXb0UZ08hJ3aVrHPPf8jstcb54NZXzE
kRfcBray/EDAPOwEatJbvVMmQVpYdanI72i5o1f7Aj93z4r+IQemcdKQ0Mi5
YVFIdBlSWQ35aJE1UvMUtEeCKPenXpSat0NMeRpNJFcCw1z0Our+il9l8gbc
jsxZF6mIdStflfNzmm2g7sBB1OPqQWK51nL41SD5Uc0sFp1X8wLjs/Kaqfwa
cvwFGZWX82Wyf6qzHfVnueb5aBq4s3rkdZl7fc+3/upEpiBvJFh48V6kjjJ4
OSdkd9O0RWgZ8ZknNimtnS3dnsZavtFLMX9NdCuYhomWS1QQvID+Q63eJNoI
RpoiFOAaWznYpsAtYhX1HJoYkMMbTUOKTQcz8Id4Wh5ARNKuGhcdmwuyE70C
/vaWkoxW9S/6vpG1mtYSuV++VyJrO952xr7a4CEV6HznRz3Cc0glBy/nxU+m
99nch0iq/ORhYzH/0/SNx6kUd2zIYycQJV9SmVkyU6YJN07Ms8BX9kF0T0Xe
RNW9u6Hk46KV/AdiVEGTdnrJ3xSdsBDfckjRD8KCXgAa1373WQmn9Bxe5/Nd
hRLQCktteE39vPWPFB2yAO6f+o4YLe6zotrqYL5xE+/UMKhDBRnLntTg7XG5
whYEUDarb7KmGDlLJMc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EphYdS+yg1CQguGA8ovDPRwCmqV+s5h0d7IosY1c2kMZWB25r8WGjwq4Z3Xr3ko+iXaiTriUrB1Knd0RRkHnGaTGCRqIsnWS8WkNMbgKfh6rQxoH4j3g1Y/SgHzCPymzsX/zfM2eF3rA68zvKupbrnGyUYuuVPwSRhe1IqeaUtK2v7Oja3pSODeKSQeEUXIgBxtq3CnuxoS6FhaF5CDW0c35GU3GB/YS+Nw1geA7XAJHR9rA+sz5aVmLtSf58O3mxM61pz/pw/NCd9BnbakYEZ4wK5T7tNm7AQPKo9TRZ3QWRkxJXSHHKnb4MAQI2rCOTRSTWH2TPb9EkAHYtLpskGvAFRmDW5l+IeBH/uQRbXGwYEQDwuXipNfMc8jqz+u0bHVCLSx+5dIPzSTQ0rxntWaEDat7ubwM9Bu9eO7DH7NLJAsP10UOBSrBXHBa8ORr8I3Ul8Wv8xHJ76ZQDgX08hLSi3orkEhr4Sgx9XLlmuvYrMGkdg9nB16OffsrruQIMArk2jtqwpFQB4UqbmdNUPLB+iwkkhmF8NFJDTC9eZPDA5pdYlvObxzRwItQoYbtkX4It32YdrcoG8cFUAURI8TqxWDyS9T0htZx1gxhWlkXNUj7zDXV2z1qtRQo9odbZzG1TkgeXwZF41J5JualvLO7YlquPX87nqZSIN42UrzHmjDJZUvSmZQnudWKzWXdJOZV5OVC+W+GHki7z88okmzX+UdOTpHpJE4tjbJfHJTSw0U03G3NX1EX2RPb9LNDqh26txbmZQrryvRpRSOzg4K"
`endif