// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lE8JGPpEQAQS8jd0zfeM4UshrgpjGDv8r8kK7I8dyZr9mu+qCnm7BUtUhBiI
fmuU6UkcTW6EQAZeQCdSCH1+YrVpZ7kWlosfAxmD62kwfn90RrvT4PLuTHK8
tUsyF6GQnm+ERcnQ+Wzqyqgp2ckfhFqf8SBlDZGQuwlxTj5f2zWfnvPs0eMn
5YBb7No6hxDkob2Jr8W05Rk2MvWwcYsZwRnMFgSPBRYx1pmSU7ErpPSqKNH2
GrFnannVdwPfCpArAI2pLm6X57Zypn5B7myBH2yXYOtIeldsvHit25IkSsXQ
sNp2Jq/7Y96O7w1gkj3zGtfTQ9UG5qs1FbXamtWFjg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dxXFtjXNYdD/Elhbt91nVIXvUTS62PcKbZ2hcjgd94dx1JFG9TdzZbIoXbsy
MJM5DGWCkVdrN0mho0RB5DjZv36VF+izisOvwFXBp1AmeiuMTCKcJw4TgFcU
Jhk7o6LOB7rgKS1MywMrlK22GwiU6rC6L6jmopfZcbwoT8bXRCX5F7GTNCDL
u2dcfI7B6EKHbDzYQl22cyDVTXnjR300B0wa3O01m8PzTKpWczAAdXU/zXmC
QLSNr07XGrtm78TVcEX99hcIfxyT+bDVpwTA//0h+LkYV4lVlb4Ziq9gyz3M
dpPUd2ePSbgh+TxgTSws9YcIiuMN5JXHAd7OEvSTTg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y/HXXo6RUhrKvk/xdzxW7aR4lenxuvv3rubQ3WX50tUh7EXNiEI72lWsWR6N
azbZLWx86yNDpC4ZrFqDmHeIDxUMNElxxbML//2HsPObt62mOtN0o7F21eHw
Sd2JgAG3FxmKYrva6uHg+7HpVer6Q10pJGPeywKnXVdGueZX1IVatezpWmFv
D/ADX/TiDz1K3Ymv5KSaJcJzJAzzNwlhRAwjpU5SzeStb+5s5uW90/ZOj2w6
7fHXjldk/GzRVKcH3SBT5onLl9kx8o46Wc/ZOFpXOcJN2+KzwY2SeJTQ+iH+
QktOQqxXN0tPYSP77A4WvfuhNgwuf6bssy4EEN0F9w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I2pBbYzn5kXTrLxqvieLJvUiOmg+5IfhM9FDnBJDntI7GPunUtJbDkzGl7rO
1UAafChehzYdDR1jyfopTDhQRHxuU7EhDaSuO1YGyfu4F0LpomM7MzvSecVO
VVeKerNZ5LMHiYpGR31xsiLXA+q8Yg+qG8OiEePdbkYNHXjy5C2y7ObT1pDq
zz9IPgJv5k7ohp99I/+3QhgavLUHFxyRO/PBOgH7dFer7X5TTcrWtLum2P+b
7Ms6+9ynFgfTTyRQO5OHCexMjJNN2HyyFYuEauBubLtcXnUX47LzO9aZ9/cx
QgGkmhwVwvshWxG11VXjEj54Bddq/zZTfmZeaQiKPQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y9XSO5t9Rg6bfspsBf46haio1FRbgyB7T8I9o1+TTXt/AamaI16TcKwb+h/I
mbYJB+mR1p8wZdmA9DzSpMBTKXHN/s6jTFXWDswa3yOAgAds1/4xFVKtNEnV
eSDbnPQQN/mbvPww+FGuGzZP4hzfDInZcQaaK2VSZpTeT9ctPAQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tVlsFCwP7e6a5X9pwz63/MA1f4KmeGyejC2t8zSIQi9r9ZwwSSph8R69OHrU
kXmzUwRrYvRcNJ3PZvgClhBjwbqH8g0FdLMnGmc9q6ls+4/K4dSEUywSxTwu
KcJiZSiXV/udp6L8sYWsLYswgUwq3speHemTB/ounsbiNYIX0+GbhpuytJy1
l9bDfY7ELSCJJmabKbNdXa0nwq+YgtfixsUNuraODiq5tLv54l/QjYr3MK9z
3kVh+KkkKa2As2X45hd91AUi+ygE0oXD7Jwt0jZxB3kJeynthGe6x7xmVCZq
b+wHoBsu1vcg0GRJO1VcgM2Hyuf/VGpiV7yeTUMRsS7UJYVJl7XcQ2AFHIkp
dZZBdPm3KUxjbRS4c4qfOGFRqNMv/Ouhnx0WH47QftQPuyw18BYvNit05fDh
FPdCgKLegbrIfqGkfw2vmvWWW3WRkDxl4Ep/58v1TZVa55uJ/RCrKEQ295rF
1Xn5gkQj7dH8gcsboaxtzDCgM6MwmQKK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZpYjtuihs0JS/65j1GKvYKTCQtb6LszEq1cqBYvJRM5zlPMet3TyTYtl39qe
taypPUOrL/r7/UDxb3tTMEhcTqWCJTr5RJ/AJUv7NC2m0OpsDwmyB68mCbFn
9pZH3WOHqWEHjfwO6Br8cefpNWjg1hm/1n2Fj++h5M4jgKeOZw4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XMmgLbBxeP/lEMeCGStVnV0iZp684toYIgAJz+oI3ySDt65FvvD88PZ0jPuw
OkaJ1uDsIhfhwElW5CJuBGCAW1aIt2ftyg6e3Sl1IHMMkpax9v6HJ9n1umH+
9eo3eN7p9bC84/B4YFpj+PUsx0+eGcJorQ+iuEvuDNEQ16cx8tw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2064)
`pragma protect data_block
rxk79/ySfcQiwGGp1Q2fd6X7FJ90EGz/bZ/0tOyup/fJ2/N5vWgQvFxZAljN
jTRv/ST+i95m99B840m7f+jp/5hvNMnsCgkx1L9t8RK89TlOo5NfXHJQ5GcC
AAOtFIuKx/w7NKW9nSTXz4TvLkqDFR2ME1b6uGviA5UQUmS6XKrdqBzA48E3
oF73zaPPZHAQFau5ae3+TeXwdP9siBZupe48q0GBlWPxtFdZxAUl/suuHBkf
mo3J3ubLKhMwQAApJkb6CzUM1qUw0JIQJ3CxgjcJsa3zkrCu3k24eDSEdpB+
8QD73/jTANPmTXr1f0v2OYcr2ysQ//JlcRKDvCzCL+TaSjJ/PlXjiE/JxfNQ
3wn/pN5Z5zMNktxLgveIi4CSD0dPYBKijFlgq6nWF4xVNi9HEREM3oZNlFIP
02NIhkKZpAZUMGna5f9YM2TKFRrB8t0ETKmvU2hgte90b/Z0qF1oLTPA21DW
IB6KtHjXwyEkk5Es3FHTtxaDcWeI3Vpb54xsBFLPVQZ/JBjBh6cd5RnfPlBQ
4j7WEfbUFlQ51KVE7KqmEAo93rY5iys8xez8MPCundUVv/GDdCW0tNe4tWgF
2Y4jG4TRWB/SuuaMXN/Lmwn3fooxE43P2oVlqu0RFlSmjcHWwSVXeKSYpkng
KwSIFmWpXOfidCoxJ8QEXhlLVLoJqCrqJhEYD+LYkRxrFcC0iuNG5ZcHQw1F
WPqgB9DWnnMs26RmPYPDfXaYWgkWTvpu09xgI8KhT/qmJJ/fRygC5F3EuHN3
U1KrVNrenXf3OYeXYx+knDyvS/O89kydH9ucDk48TkXnCE4qRaBZ5DMvt6Qa
p7haaBfuy7r+jvsH0qZPQ2HswGsNHGAzFu6J83Ol1I0kpGWxUP8DUGT4vgCz
Fu/iOlithemgJEVhDcJ6dK4LH2wE3iZ4cfG/OLD2K56j9TO0+PGbdobc8PdS
gsFbmYebFyfjKMetnRABjA0aAf6PL+82a8P8fnbBDBU8GoNmdiH7iC4Abc5e
QmZNh5PSftd4pAdoV+nhgt1jfaduZO/KQTKelYjrkoHkb1vdwKM5EJRZFO1E
CY8zPAy6pXxSXE/DenpPIY4tqXdN3gx9ebYFYLKwnRxyaig+3uDlYS29/wAZ
VC+4zoWXkCy39XvswvIqupvrdJLwR+cA61lM1tlT1m73+ZogZGCZBTuWdeiT
eNqsBV2YcGw8GPkXep4bFsXTc5I7JfI4VN6C7e+GEF4/Fv22dV9OTHoa8kDK
SzRW6BAQSUQYg6kIxleZ4KBU9YDAhlPbJnSrYN+PGG+d4XRWP8ra2eK+opPu
MGEzB1DsVPlzk+iKE5ZIQRFXGQdHM4cXhMMzpQSgmVJZ9L9ZwpCcRlFXJ+fe
shptm+ncbSnnQBQF6Dg8fXwCqpfMhdZ/xI3ooOMFFk7LRlN3fvzIzxShrjl0
zvBWi2/yapkXTFgOYFsENABgcxrftiUlp7kvmXWeUU1Zh+XvO4E9+o3DaZDI
1MJdB/yvROVOD8DkZsJv8q+KHcADwwJHEXy50F5gQztJSNDQlyIz7nVyba2q
XfUf3XfDgy+V+11WL6COD0ROwEkJlIFHSygPg+6BYy07gbsQtqdCGO5+Fucz
zuOVPulcJGrR5BguWiMFEj3xKiPxROEv9cEUO5DHxHa7GREBwbwv/AaIh7tO
rTSEQ4j5teflW92Z3tHXk06ZgKvxMEasrkGx+PWuTmTdhWUSPBTkX5h04aQZ
vwIwPqQfyQRRZ/mNmyNbnWypq3sBakeBh70w8H4Gbps4Su/vxVKRT68l+sx8
WGB3sCQbnT9jCobwFYPx32yxZQ/RZmUagKH7FKH6vVXSWZMALroLiZdTYPLy
D60zGVCXN50RKK9krtDpV4k2c377jlfQjck+x3KhkH9VFwPfUphZviY1unIh
hzE4N2kBUPT4scOi1cow34yFXbDWVixLoNA1lq7FCo2Ma0XxDbPa1jkNA3dc
JpZXPrSJgJB9h0UfzvCloRMOOKRMPPPUVaK5uoTpxBOVeLO1PxYF/GmhDJwI
iM3t/S6DmYUC21u4WiTL+/wKy8dw0eqZMNiDgVw/tVCSzAOfVpUDu3Q5Td9M
EDeAMyFzn8d2kmnGFBocctNriOa4dcB3vYg7DrkZBWOVM/BsxfRpm3LhY4ya
8iXv9R6yyejTBymfcILe+07JDweb9fcHJeFpSx4RCx3TbKGI3RWHTqsMMG7I
LGTs7pHfRlv4ySWmSFp10sLkP0fCWldvZaQBwikfw0cG4M/cbSLfLOmy4VWB
zyewt9KiM5nXzNomXyuTFEZaoaDD5P8rvF81AT930WCvnFLIBCo/Jz3BRyfK
FZ7S2jcbSBP3qr94dg4IpqlwAGub47v8wfccL+xfXs3Rt2+4JEW+nnuL75nx
mal1GDdE4CGjkTDkbn9bh/Yz7gPw2ORMwwu6QcyUBUoE503mmbAOprX1OxTX
E0wuiQs3J2ynN3CyNveByIA5N6M0B6gPcMN06bm09WoHK3f2b/ZxVndzH6k0
TC6dWThHHl4NnMaCY5MLnMnqKn+iW7ZUPSv8vK10MlBMsHrFWXXkVcqjujlc
lY2HHSrGL6RQgcNtJ337ICFnOAJwbyrJbehspnBjtlxMFObFSi7yrYUB2p4e
Hm5Ma+1gIl0g07dH3s62Bd/yJGnA++2tesYKOUYCdhKPOyI2J0jy1zcaiyR5
nMKfaLGGjN2xqycZgp00hFtCEmgJtfYl7qE4BwT8T+K+on2HUzaw

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Jsn4SKOFgoLnMe4GQGdWoZEjCeUgE7/3f3CHVfgk8UVx+meo7VdKx+fcBeI43EQnZoDtxX++QGTjixTFHbR6NP+pc6Vy/lofc2nJvzUzAwNH+H/m2WkYi2NtZNc1ACAyFY/9ht+BLg90IWUNa5YYoveQl+IkrR5TwTKbVgEmCGzlNAZ1DUt3moso2QA8JyNwujGW5VgieRawANuz83vOpDnRhmCuyGiDG/QGaQPn6t0kM3MdDYa1Gz0W9N6T9kg2EtQpN7LEn/0Oxm9UuphhQmTNb441892jykb9Fz5cdxcSvbHCtfhDg/KuR611S9EbB7qJ+MVsUQOnWlVkzgit03UF+txJWnKZQxdO0Ng1jDj2elwZurg1P9SiBgNAoJWQslIAJwypZntA7r1vDYaR+mY66YmB02Dp4E1giKjv1xWaHnrH2zu67/HWZTi4qdUx3SSxWo2Y7dHzB46Pv/kgoEKe8cIE4lTLeOsM3Arf6Y/RS+SrMk2btomHYPnMgRyGhDdo/oUadaFH4S4AToQ3f555yxEiDNX+R2OCxeM/9qItQAaNOxAGD/SNV65PajXwLF/d7FpiY/IB/iP42fZUpZlX5bVAl6C7TCuYBAAJRi0y02/MzoqNpNzE+gLo87w86gEbKts0kRzc26PI4khzrlnINMJaZpSCFRRs4QOF7/InxsPOD7Dt0+Tw6QpghkWqDlWe5pCxJbzSmQQ6jHmSToY/HGqzM+4LJLhQfEFDHg2v8HKcJfh1TECPAybyZc2pz7hMm+utSbhbf3jjN/1L02"
`endif