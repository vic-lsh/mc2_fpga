// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YXGJwgxj3h3EeZkF04G1M6P76VcIPq20CSm5v+lrun2o4T3zEIob+wvDl43V
jWV4tKu4A89qafyrRAt9OqzBLaZJp/lJSZyIS/aKFRydBB1d19Y3GTdIFt4T
m5x2BzWMjIasQCg3gc3Az6YpzksJPjxZOOJGUFb7L4ndx7TJexGAycH+UEKx
EdDQIAGMTYA6dcrMznsP43zs8DunyYH5oglhhiOUhCpinxQ+iIlpn6s2oIkL
2FdP1rdaRoHP0wifFEE1dhTW3Wn1qaQoYhX6kJo6Me1HCXmlmUuBz8IDC2Lg
v29aJGlNmh7YEVxW+1ykG14GhGQdFAJl9WkwZJVm8A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iJNG3dP237H2mDVfDh5xwnb1AsTgJa/8jkd+E7SFuvh+OSvjNa4P20Z8F9PQ
UCvu7aZvt/xrAkpuEoFCUWAiOQxRYGXysnQfKLTCYyEpqX6Pb2jbFUp9rzHU
jOT/ReVllfjpWpt4JMu3T0L7rClcafIaxUpJr2vlpjIfM2z4F2nWuZ4IGK30
Yf7LkLRvbRYZZJqxFOXumk5UdHc7xEETKxU9zafUzHeEcbbqkNQZg9+342iQ
MVgyrUmzQ7xV/22sQZ7VVAJPw8XA7hl+VfuNKCG4umikqP6uUn4XITef9CBh
zcAZ3vFxEKk8SPyLdDaq1O3uhjdKc7sxsSMAAGgFlA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uUQotYt+Nh4+FGkZcIv0Js9mstAYmaDR7nvXqanNJR7XnrFFqbNq71EFftkd
ENhOvhJ9p4PpFjukF5oy7pGbx34zeDAXsTOy2YJFf3iKd7iGpSCLDN22VP7e
6k3MIA9FiKLn7MWZKb2ypKCP9DWCR/WC6X5hmD9+ACbInT4vc6+8rxwNRK9M
Ze9EVYApDvGoVFhycv/fgq0Ek47crQWF1QZo+Pa3RtSN3J855Jxzlo4ro3hb
nnbxMUVwZ/OVBTWYnkRurb4ZgWkMZiFGtRsyO9eeeE5JkFpizJczlUW9tg3p
7UZYfPi/M8voMgmEToZC8Wywq2ECrGRvqdW5pw7txw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ojn1/gj89qAVymPm8PhRfx2b3IiHBI8OVPbrGrHO1phofkQ1L6kMnVpjVxhL
O9wQq53qKnj74p7nhw7IQa/6TCeRgs9KgSksrWVgcGbpBeER5PfE0N40tozh
XzVDXK12E5V/CWmfm/s4jEHnW8FSSToqucZiYFlecxw7BFdLbRcmt0cDL73A
/PP4d+ekeMkyVEkBUj4NeuLsBrRXZE3om9d1Mi9MYbGQ15sICcKFsirCJccs
kURswmYQuSrzWoKtUSRD9LQJbekD1Kvju1NAvem1YLERQMhDhnL65MwNVFkd
H7x67z9plHJezFkR1I3qX404ASelTyiiZ4DydEP/Hg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OX7GrR1A8ro08WxKGmRtBdRvxXi727sYWALu/OW73faLookuuZFlNVkqYo6G
rW9D9w4PWy7Q4JHK4RsBIaCfrf+PdQ6Snsl6iw638XucUrA/tRPh/tHRcGOQ
EswLyEsKerFls69q2QdWvAKNXfA5TxR/z/+JOXgLlhXogHB2NM0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DA1eOxfTje97QodG1ONNNqC56mEucN6rAa9IFu6uvdCozGpvm+jMkhJ8FOFE
vX+qPjM9s1YXwHzmwIB7vrbXwzNDfao/Ynxevtox8XQitooMw7DrHEKWm2hh
tGLMhTFP0jkGfrrEXXFYYVUAyz2g/RTgZR5a4xzG6Omo1RkC4ZMHsE8/0EEp
mkBSudgtUbOmQxzWZHb1K/8pv/KlzhzdtRTEXSFrbm62QiMH+UJ5B9tPz+zp
d9USJuf/N6Tej7iXuRrG0yy1EUGQikZHx240lzCn5s/gzMvgS9mqtwhpoSEb
2Np77GgD9s146X41/vXoq7LnsqGF3y9AeUPTiZp1QSXvL0SrpPbY8LukjM6w
YaGRI3qUmNugu1LVfFb3JpZKQaZV6B/lIQEmu+UPazbliQJ7IYYSyZ+egFoq
thprIgEEVbnaLWaSy/scQdDbZVRz43Eu4jp/Amh49aHwrTGYYeZV+t5XtUlw
UHRQPVJ/+LTZrMD8b7VSGYrzUL9IJvg4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KGE3drPhJPI/UN5kJhxWcYzf4hK0X35v0WuUa4yaE8Ryjx5aXf1sXmvGw5cj
raDgTTuFRCr+E57Mj67ZFyQxAoieyeDzoo4H9ZoMHa4KhjCy8rrKYCXqaWns
YbxdRyQH6B+/3eTjzuqS62zhcnQr5v9z3XOBx46dOQ61XRWBD2I=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cPSd1yVhU5VfLQKoWkxidKOq/TjU9gI8jFpx71YTv8WQVAtOKzDbgjfTeMpq
xFz2xoMZnQwlwGGqiL9VATP5gy/YhsaMoiS34HOLzMbvhH0RdMN5Y/LvxBOh
8lOpph08jw/ae2gUKhL2R9vBn3a2fqsG+a+9ni0DKS7c+eIrlqw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8336)
`pragma protect data_block
TUXz43nfU5zuRTaef4KmbQNXjy/1RKy90evWMhaied4DE13c3d/HujbI6F1+
16MwEZPiP7bGRV6ugP4xbwvbraoryz2xYp2FyGjmf2Gu5VCrtr6hAanANdIM
OWVOFYCLcWxU0l3HYRT+WvXNP/ij8ry2FOl01OTrarJj05iPltB/AtmSPfTf
tmV0Ocrno2LRof6cEu2xvAOZLO0giCIKbYF7sZ69GhPZ2/TZa93RKpCdIKwd
zO5P6tt8IRLqFDxRSlFr5+FgkH2KvsHwrnBDhLhcPbjqe+xzlblk8/lkbWxr
PyiRjnD9u7+htkmAuQ1rOtS1xDmZbDd9PxFip99i/FZAd3IKE26cWABR8lej
3yg46arKGEWCA0sIi4zFgJAV1+SYhkYAbV/BOjldLzVT+UtCf1yP5Qt86dek
rjmPqhSBTA3amxEdFIG/w5THET4P9cJPWDm1OTF48vBC513O2elronlVEfSf
HjQKxBdVE3k4VxIVQzMR/TbRaTW+ulIs50VUZSZUsNurzhM7nhx9gzuSPhp+
uRAtPfj+zGWh3Nw3s1XtCmdl7FmT9cAnrb2iIjktIfBYjskGYU+Pr4keIfTu
E3gXOx2apARVC9ZQxXnOSovEjj3Ze/CydRAkg6LzNTJguSMcyU8lj+dxyZ2J
uXR30h/uLKLnoiw0FfnpGNXleTf9jihaUyuH6yCAcc4psuHEf2JTtR4mpYd6
RE0m5vLwMp2NSmTCtMAgQGmtDJRsua1EjTlnjPkKan26UtBY0/r/1GK+XabV
t/XYie//BkFqB9gXpuDpJeHOSM3Q9ZxP1wTMNivt4OgsjUT7c3ajPJIPPciS
q/kkel1SURghk+7NCD2MIEUMXC3kByn1mLWaaph9WVbG0SBAIaAR3nP72Nbq
gcQfJw+p3LDnNdQdUPWvEPBSO0yfFDn2Yn+bpi9hv/eHtaC8QAwxnx0Wn9Yu
sFOT0sTdNWJQYH9Jhvz+mNu0NdAQRIp5eIEpHOVQ8KummMQowyWVWroikZHA
t7ffU2JnT9NA4rTskrjfCb+/d/PUp96/bI5FwqUUbiWluR8hlWyUlbrOULxX
l1v78qMh/TOYdmm00kgLYuly7RAVpnvLOqdKC4AEYPXxpupS2ftVYwfMC513
o7raal7PptZDxArQ+qS+O0Ml143gjiYdafajdZtdAo5LWICRxcbSBrp8dt/X
2FzinuW0htltAU96Kpi9YNSWuPvDMyABY3hmHffXq4wxcUTU33DiyTowHDE9
3CClmox0b4M3tETOcloK4PjWGGO4pDYGBlMKLJnD3W6yQjTyElgP3u0xVVrj
XLxPkYlD5ULqHiHf409bB9cYJ8uu2D+zSRvYicVs46F1nXlaEJmb0rYoaOHa
4Y1C2Qi/39i7P6SzVkwn27eJFlaIfd5jf2o4tRNr0FOWNmOlrFAJLgpx0ZXu
bXpe/eP57bZw+RnKej5Cjugem3arOYC/PiKtqO6LbBlxvFdWCnIdjHTePdzW
w35s6HT3jiZeeOjqO337gvwmhSNsGCr5XFw3h0VZ8w3OAyhfSQuMAF0ldOpG
+vZFrQ/y/BqGDzLWkpAKOnjHFv0F59SpH2mof/lZxrWM59fEOaNNrUC0jMaX
MQqt+MkxwiSp/osh+K5LBMRJajXCPa1Mv6hADMFFMtKf2bSWXl/QfDWxXDMa
7CmAQMAmauzW1ygOt5UWpKRxfDcvGIYClDbi3bUDp2bywlCkgQCcIrSmLI8r
E9qGTN1WP1HqTzgXQyoI1hPWjgdRT4IAiVv5mcroSVNnQ7iblc/QWbuGoDhW
fm6OCji2303vSnwFCut9Pfp2gVPCwUiQWjGVw6RJghMAFb6msPOZy4MRL3EV
j+CKbX6J7/6bKrvlIbY7vpz2s6Z3APHZMY8+SrHjeJ78K0FL2L7ESj/Bg1N0
eAhO53/gVJ9NgwBavuIWm6eFrlLTOViULEuIjOewHvSQ+dXLVjs11FF9lgZx
VlsnqDKd+q5gGeZEz0cOKiN7TUmdbmCYTrng4tTuPojuI6RXgbgU+KE5qPA9
EPaO7QzNys4x8VJN/b4GdRYFwWRinxGdLeohyd0Ug/i5z/RD6iwC36OYbhtb
il9sZhgaT5SHH3hKEQ8g8zUY31cv4cIja1lZg9eDlsh+lkLKEaBII+K5qWY3
XTTEjTTqKkAIWvTTOIuAOaxXG0FDY7dpULGFkq/1oQILowW0YwjenOlWC9NC
175MapjNrYZrQFPEz187t7kqY2v84+zSPZ6JN+oRx9e8JpuYmfiE1oufLQfr
m2DxreEGaqYjAFi2QAup+p5bAZY0x3DWnAP3vVjxAHbqbCa+YEF8ZBOEPJTm
6ShKdo5+cICTvX8mXkBrQ6llmfQXZ7SEQJZQeSIhqK67mw4lsE8hVKIP4E1o
+UDBxa9UbGTVVzJHM/UUw0MJY9NDlPCieHTM2JKdoIj8Arpy/aZPl75ozC/y
FG43esRomZzqny2HBZaQuPjEnrdBM9Qg0xc57Rc8UIYeK9lCH9TtaQiX8GuK
4F40xAVxzcvPlgs1vNmGZTSrpZCagv6KT1XbQ1LJX/i0qr6JA4Lh1TXCGQWW
rUuUG8qbPuscFDQha+1JETm2mpg5w2l1sMfETGF9qBffoRMCelJPfQfJd5NH
z9XVRg78xc1oiH3PhsMs+wkYjQvLVebzWAi4sFM7j/vlrQqD1Qd9hh6kUrUk
BXrZGUyvKz1NXFg2igiM8MRspxQOaSiYSRLRXgUw6kPYELzWNSNNlqo2wwe5
5D13sU4VRtxsxdtaRxb+xtOPfonlraOhdYPipRSG1RjYB912m20nKeLXuOnX
NYrsQOwiYLZt3Jyo7lYQhS7OdZllleHw4+92NWPkFrPc+1nWrM7bAnapl9X5
yddD0qP5k40/Mhis3nIr7bLkkDU6WzMXN9muegFs85l1Z89Tedh6gW7AJZBG
UJwi/aIkOh8G30GV7dVYsOcsRy4ATFlk3NQzgoIsQhNmgE5GfIFuByUoE0b5
7IrcRwHWEU03qrP0PGtne8/bNDpHHLErSQYpiTfcpgOP4cHoTeXPmnmzKryI
hgwLQ4sCAVTra8D6HHh1LRSjp+qmok1D4k47ZzCawb+Ctws3G8NLGZWQ304Y
/nZN+aguo22F2BGjU04MtLXXB0fUycT5aLGgpvHf2BE4MevyZ6F24UNYjZgQ
qJjePZ9nlSfwKAdlBzQgWpTpQGDyEYO86GYbu1xKXmiUlehNtvJW1debQJi3
ED2sGq7WIkKcMIpAlpBXROQwrNqFFabY70TM5hLmUoCb1deqtYJuaoghmLgk
vvXJebJnpl/s2d0wFzYf6NoTRsNisPIxCF/xUjhUJn4FBRRZTtQB5FVMvH3j
QxefLYlF/djP3WA3mlXeHfaZ8GSmwcabjpgJGgCEPIDKme+7oPzbELQgVtl/
TEElDed+DWoFg66FiqwUzdQ/VY/QrtHXD/7ZONS0DUcMNBxV0sBUceZMHmih
w0sZK16tkPMApiTEE8zzTnTxCSpf3KGhw5ToOadWQ5a09fW5Fm5BTv8rPh60
2omdfahNlEkrTzwZewewqY0ZYsUsOR6WeQWowvLlf3b1tETwGR2zCBmxAH3H
bIkMmBsh+l4l0PV+j6p4qAG9obwAUQaoyITDvsG4K/ot4ppPtTZyxlDne4W5
B+90N92KqRgPtujcCJXApnW08oPfhOyqG+fqjCAvP20ledv0cB0RO+qqr7T9
N4/GCgKfA/6Bt30BpnMrFHCFk/Zwg+h/zvD3/sp9xhd8icST2Gbj3yBt15nm
mYqJLUv+yz5N9Lxl7uZqWY04grZpyQ0NIl58T9pBTG7VvCQnEPW8CMMNB2P8
pH/D9eS4sYLRuTJsdi1MLHBQsM4e96irCRLuUh1Sh5wIrD0aSucLh8hXrnOD
2nPQghSFY25pWMK1zMX0YSvlYjhTe1JNOy0yUg7sdDkUz0n3JFFq39SXeSO+
coooqjCiD2bfaleb6mS5lmrsAyvmEnjoSAE9dn/f6G6MPDUuQvt04b3SxtaA
RENAizTM2ORaCJhzNu1UTgxAxYHpk/x5Zg2I03p5oYVTiVVNeeg467Mdpn0t
8HFRNu2wzkP0u7t7LVT0n8cv3Z7M4ddaaB4KESUiq2ytfT45cgycTkgEyRT7
iHVfq9QtXJ8DOmUiqR4jfpmj8VtWboEcYxH3Og9n2sFXkUYfTZM6W4D8XGgB
Gh72XEOjTbtlRimIClZK7aiRegfX+VDl2BwP+jVwd+Fn5W773GqDVKbjThog
HKBDFShwYGa5SZqmHcvZY3KB3NLgMZ/JDoHDjhFqCr7zcKFVaK8Zc9a+kfEA
MRyKYOxxA5aLrD30mccUgyulTFsDvAs7ESMXP7aCCLqSEgUpi6eIquoWI36s
obLWQM5ic2vecBiY400x2nBQ6E2wFUfV3In3ejGjgFK2ohMLD3BXVpvgnfZW
/npgtHPy+xESTLpfosWzVtyC3Nj+ShgK8EpB4CYVBPULiVNEeMo/xvUsmY3C
Wos5I1u49z7ncEO9vuhALNGrzZ8gWu20H7RRw2hWdgcKZkBP/Y+lFvtTSVYh
nGixB5YZR6s+CcTvq/JV6nWLd+Abu612Hnm+tlckTevfAwt6qZg4u8ZlCt3g
jNzUiYBwsEeRAOkWSm9C4BSckzDteOrtA4qXEq34+aagX57AtyJDGiUj1hFn
ilnbJ1tmYYQuscGqII1vwNVbso8nrxizUs0Qyz0yEri2FTTh57QvJAlXICk7
VWXAMr8HmBnKruTInBzqZwe5kjw0XP1XROt7IR8+qkgvoT/s5OhWxoBr9z9N
5WtweKmIyP2cHWWyO9w1dKJYbNtwEHSwE659pmRZKI69GraT+hZmaAv9EcBx
wQCXChQK0qR/wYxWtYzI2Zk1YyOHlvzP7Bhgmf5ASL6gCGielOnzLhf0b4C0
Ild770geWwPya4hdOgg3cYL0Wtm77TI+OdxI4X7qg9WAgxDbHfsMEdznnOaj
6UsI6j5xRoS1BRn+X7DDsk3ZpdU54UM8+sCMm9LpZR0Qg5MsgGegCU8At3Cj
kUfyfE7nqa8nCfeb+gGwEpkQd8BTVIA3IAOe3/UkyX8b8ZVzZfQvGNUaKXca
iG9nBYe7n2oT+A9Z0BR8u53xnBRvwcfIAKz6ISkCAanceALolA0NSrY4VyOW
675kJ5DBSvr6PGE3z054fK37pypjAG7X0feU4kQtmEtNd5c7rrSVraVo3BtU
I1BSHk847Rr176u4p/hqevkcheUmnuRXmdNrsQnwtoE6fEMa2j1a9WEdXIuh
5FPTvsFJ3aKL7DLx4yeY2Mld9K+Ic9YnU42v7Eec9kjCc3a5mo/VTbazlalP
IkDaBDbphX/m3JDS/SxxccYZbqIovXN3wSMOQqc3fLwl0/RRDaTUXF/MWjzp
xYMfg0fCYS2baBayRbDDuwvYtSA5BL4de7O1s6dVutdy1NEo6bmqNAcFzCYs
GoK+9/jIuLA3oMaKTB6/3Gt79Q/L6FXK4UNKluqlDMfCvd1LT3L0j/3fPQZ4
7hlWlJ6cFaRki5m22mwBvfMHX0hsQowtYtnJF8Ra6fuyQYTIR0mBmpRWK/yO
XmQksO1MyTEdMGjf/f7McdRxo3lIh1MuVdKxOnK8QBbt4NeWkltO1oN3hrYE
otCjEfG34JMs3UYVQhBWraAJsde1g1CL4xosGrVE6mQmNp6fhg7ETh/l4LM9
z5+UZykDj+6UiwNUjkRBzLlFf/RblmG5cAeCZMtYCpgoqpo3sQBSxS0t3v1e
ZGOwqig0zJ0sV8K5PJRUKPPn+T+mwPLTsrVZfViJDaOJyUQ3K7uwCnOQK9Ci
Q72AZurw3vAGCKrKssg2baH9U0WKsADD6d0EeZU8C2JPXC6FIf+5XoWPZGyO
ka/e5I0Ap3nLZKvYzYPlNew8V0NkVgzf79+gg1AZQV9pU4OI6/OA03uXAXow
HDNMA4p0S4tQcNMljmMuGnkJzOUaT+c0ercoYX1ls3qAMsef2zfS/nrWDUo8
j40NeC3Lja3CsYm95ZvRC4WNVSqSwccsqCnoWUFsl8jSaNj9NG9qCf6/YF9D
tdlFrtCI0XJdeVsBoF52L41SVTIL6Y43LQbPdw/pyKPI8vX+gPFSZCS8CPuL
PTycKv6SfAi1elaCdQoNKqhwaDnFwasV8kql2eSWWAQ59R2LwqHvplH2PjPO
uwb5hgvxJPEzw9oIwx9yFPe/YoaelZAED2dnoMOe0ErcnieCloxtPO+8wd3x
nNu5mCJspQSsdi40/1OLUGaoDVy1CFiFc0jxRauAMoxgUjoQt7lExkvMbLfg
zNMIRqFGlsn9d0YM7C5uOEL+706PZRBAwkRs1y2dvj8UAAuRb7PtbDyal3ul
HnuZR6Zt/7zplwAYhI3H40QBcmtypR9lZ7w3/i67hzAsuIdueYddDbCDQMe0
ERBjo+tbCpv19B4APTd2+n5InBVenmeO7lhSaBz25M8VxkBithR3NeTyitRy
bpA9qPEmF9TLYUcVO/aAiF0skV821DCItJ81tfKKBmcSWOd9jxNFFXgEBxco
X+HhonphdI2p6C4zhPu3UvaQevq83gRlAo8QLy3AlrhpqWV8UtqKYQ8p0pRB
IfmxUusBBQvTNwuOvZtCiCSI/4YHVOI88f4GLtg4CRStHornuLmlqT0KgjVP
MQoFoU0vQJ3Mxty4DF3CFk5Gh0NvmNGzpnGVjmREh+p0ztuUV6nJehqFSaL2
A+gagzRiOvxFkKRE2m4h+pu8w4GLO29030hmoq+/SvWJ2bjGfyhoJ8jPXOsk
7w2D1Bndae7++S8woa2kdubtnBKh7xGZMBDomFVHNuqW0iY86+K5qaTIHIVS
EPXv8mHkqD0Y1WG6Vja0qfCNg7mzzY2G9zc5bjAIZj9L6M4EndOGmr4eTojl
6CL4JfELs2XeGo8v/Kyrsb9eLXZYnZUXPScbKBbBdjt/vNZ8ym+/nhmMQLM7
6XnpTVpR0YTbNQYCETLLxKSt8Opx/qMKSX2dnS1qy9rmeYglxiCN9NS4XEV/
O6INsrxjxa4aKCsH1YAIDkbQCL5QBtCMP0kAG0AMTFsC0KzDdgLQUlKopsox
cqHI4mvhbG9oQ1UymKKo67s1S6E25M1llqykD0jPrqVy/wNjA1whVCqcjcn1
AcQax+UKGuCTP5lPUQvaDQ6ZGgefDGvbBQOyq0e57GENByZlL8TugE2I5Nuu
Ps0x0dUH6C8aJE6Ch9YUyGvztGctv6zxUzuVtIfukbK3p7odD1B5q65EDAxX
VKW+8XIiXy627KxFHopr1Q3NMRQTHcI4M+wYUgw9HM6sW+BDWHGqwuyW8nHe
SZ/N/QD0bj0TJ/qNsF9W6k36UqfzpZFlN9fXwOS0pCo9kdbG2UkjDoSrpo6f
JRuC051CT5DFUNNpuTs5557AoTeJsV6hg8ghTaBv/ZIR+WyJkDVLFUrqdsWt
VKACJusZZBgaaAptYkoEHpDOPejABJZkiqdXSs8tQhKwnewBAriAjj1xfUnV
ystqPy26uPjedX6l27z+ZGyJmmRZ7jPb2aKHe5/wAOD4c4bge+3/bfJyDBRc
zimPCOwNCe+U4wRYflhTtbQDZ0Kwri2It0J7DxpfkW8q8TgMq7n84RqLGo5f
BiU4l3Fs5yX4yycY1Ch1fW4lXxdt4rHLdOA6A64Ecgey3247IUxuSYRFW2Rf
odQwN4kM9wOiNAjMoQJqvYRg64ub9eRbX0hFE0Bn9VxAKSN780xx5Cx8DTjz
F73y/mXRJUGwg5+LWobCZiTsgxzUEZDGRmabtubcjq0h5Lf6kn6Cq5Tjgoph
WN/rKtcsKTwZkIYzZPsEtcbOPUxdsehuD/D73E2jAOlBDGyYb4+0Y1TY5Kzd
jzX7a/5Y0Sc2EvG+QE2iYQSKSTxAqu+N00s1E175kWEF9+kkdf/HRZ7NRlEv
ESd2KDs3KTN4J3RCRlLC/IwBld9yHynghQrhkTblNCbrPCgRxQJAqzaXI/9W
jp23Mao2poQuv+1TZrbpFCfq15VNb4GWOeGoQCBq5gMDI6ZyrPAFk0CokMsO
tcuibYX7NuSzl5xlTh5UoJeu2A9g+gBRCH7DC1GI5yhnvBLomyUGTDrVrxrT
8clDRsnKdhlChRGkbjdwiY1NTcBT5fC/MKT5Z7GYUR4NL5jNh9IjNCZ31Nlz
rg1nQN9sxlDSYGCgZHtIJIpxdBzk4XaDp9Ml4CYg6+ZnYGpvv3CEOi+jRoMD
2sMpn9ipItD/lKG6Pf23lkOKQagMH38swYsyyPi/0XZdpJF1IdQOD6BY9ZN6
5fF5gsGXkp8UVa23wdeszuwiMpGYBFgjtss87yhSjwsfgqEZ3KV7PvGOJdwF
NeAo61++bxayl/XYfKJz5e+iObzzZsMGxn/i6orVijBQe+dkb4RJAKtW652w
6kNe4qJ4dyAukEuIvCaNDErh8ckRHO6KKYYOmAdOqfYV0rS9kp406VtzkTTq
kOODSlfvobWzPzNMvt7KGsJ15Q0m5G4gjmqS2NbHGQRHnBbopOJuLPU90IGy
b+z/3pPUiRu5kxh0SLB+ZAIQ1AGEdeIeHkCJm/hHJTeeNEGV3fRT1G7IA6VK
A8e4ootGk/QT/YPFw524EBCH1A3CzIJR/cY97Dyuso1wjzdu5U2RYb2COTVi
JuUJ+QnEue4REwGpxzSsQ6jW+MmodrMvCdeeiypw9g5r6vxVeARj77QnzVFr
c4dtr5JMrL+Ui/56/20VD4X7SXlA9hJL0k7qUGAcMj6utLwsZYgeEnTvUjOw
dT8A62kvK3YZs5Zw6SawqZEy8AO0TKjq3oExtFJURNF0AQVuCKkfWkqw3vjm
JXVMN0SmJN9BsuQdlmYea0iVFzpI9EqGUAaqYUs5xjtzUYbL3mjjUJAVzS8+
55uTZod9aKVLUSzhnaXYr+z9qcfFftXQUJgswvQQZr4Lz0KBCr6OtMSLb2X0
TRAyPy3Tx7H4TdXHIUUDUWcp6WZdgc5qC+PNV1r0YMLSkprEpXFP9nAuxDZn
VyjMjaK4Z7QqekOm8dZuUIfyMLkkVTGeWtwCjy89/V4h04iW7OjN+33A2nUh
DXiZQoFOSZ2yhmBz8xPkbBrGue9ZTylJe+vC0QEfK69H5Ud5gL2lMtKh8Qbz
PkCFKq7hC+E8EK7u1cDQveVwTPXaN088Gtq0JPL4eDSYvgRSNtKqBJlRQcMF
+3SJFZO9GVwIbUdbBxqE9Cl1WgWx9fI5uVA5NFvn2MOHKWS+txw3HDE4wMhW
NQyTqQC7SLcqekVaVFTpXVSiVq4xZTz57bPnng/Lyv3JH62EOL3DyFDUb+5/
UpOSCfjR0EKHQLUFoDsjqsUwuaUfmjew+UI7VWfdsIpKiUlsgjBbDjqKbCvu
MPjDesZdkq1pvTmvs+ynrouEvJZLIyi4EeHQnwNJzzdBRrvKJmY0B4Xk+D0t
ukTmU4hq6eP75WraOZgGCcC2HkawqI8koNfaQusz+bq4ui55D1RdOxoJWgG7
vc4fyytz76iNn/HANCU0CRSYedB9Z2TdgePuj+1k1FJZeKqWV+RTzsMnZHwN
TBar4jXqAeRBsUthJco/mEZmCoTmtzpnkIWPOqRqis5LgXvYhRF7mKoMfS3t
UZUYdzIDR6zP/+9tZ5B5xlSYGCKK6/2CTGM5QdYEm2Od/8JzYRbOrK22sxFH
zjJG0aoZc7b0Gmwf+TnVy8Lsd4QI4p4USFisAamMi9zYiWUgwPGpyjnTyrDG
BhFlJgGGkbH2r9ENVd5AD0SbQfoafwq12hHUJ+o/0J7EXScbIX/dfM1npP80
IoGhCFidb/xYlIWNf8YtRsabuQYe/VpmBvzzp5qX9gChOClg7llNU38zfjyS
W67KWKGG+VGEPifukt7dVVek9eVZviXjnaZ4r7EMR47gQF7imePbGHf/W+RW
nfFWE78BBLxfUNRET/vxIRLiJ8qH8ab8tXhJc9kAnyStz5iWxN4tA5kDpxVj
2KoiqCCOYd7q36r09NYCpw8DXWrdQpqnyYKjLEYVRjwecnf36Y64IcC89G+2
ET6qfe/7OKP9bDuvByH5qQA08x9aVEjuBQvNokoeQQvT4gP9Bt+Tn9qy7oYb
aK4X5r7NdRpBtlN19bydleQwVZwzyer1ZeAS08iQP6+DYX9YAU0RPW6gNZWt
fER1q3kTAa8EDmJPi5djBPoUc3Wo0eizmdHEaT1vI3ZQp7h3HjGVClCFuMbC
uP1gWHP04nx5pp6Ox/6s3eRZ4IyNtnz/E/urIlSAbOYo/OgQiq8G2A46pluS
X/zFTJbC0tFf+ArSJ9C5ZKN7tjMBLKVNONktXqiexou6eC3tChHYDz9/uIrE
Vx6PTW+awDB0V8FzKjDsjZv/2D2xJyVGl597j9ocxVFqtdBZFO08gFZ2lVHH
fIzl7dXX9xybsJMEJQ0y5dMCgTfCP6z5uxy36YLtlJKT3HMig8QFV9HdhgYY
xCf1U6JxFaqTON75zTNcJHbkwv8zhx3IJ10y/9ijzUBIa5vN02NKh67hi0SW
vt6DiASKyVKtdjyQRnv9xw7IxT6/UtvgqoP94OQ/ppu7+qDcE4STT6LCpLNp
CLNU4wv90iI1yYPSlLa4LgjqqtbaCcDqcq/q2+nMIol6kcCkwhV3xr5ni+z8
5s5Regb8S2eKr7ohsWRqDr8D3eOckrZ/aG4OIYllBDhpYdkOyvpw8DgbTN4d
P/Td4gpeAtmxCbHuI+NpbhChTbl4s/IKJ28OB/1zYEqdtJqvPWFcz1vpIxOz
h7XdISx0OApJop3BUEyzEGHWZxql3frgfVquITmJM6iXvVbDHQyHiFUKyYEQ
hw8le10F6Np9F+yqvjgMejDdf6nd5g4NOAVUzue1lU5Ur9UCf/fDdnEwRLrU
S41/4x1F8f/hqX9DEsMzJGRMzwl7ME4WAg6pV7JEns/pHcx0Y0mELEzNgHpS
LcRi4tDOTclIYtUUvgV5gWyU/gRpOVyi1sBSsRVBL1H8CP3h9ZFCK9OXB5tU
zCafI8mOYOxFd/gaIp0ZDH0Y4jSySGAJ2t/1R4i3rFxo5PWqDIvHuX1pUCbZ
LAh7LvNuH50yAmjKoHVB8YqJtOGvPVgGfBigE8DodYvTV6RDXj2FAmWZ71Ua
fRe/y1qRD+KhYYI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoxcmCvV2feNFzzH0lWMEwo5tPt70CYpWl7SE/lYLdu+ESHjgsLuBR5dSv1l/lWtOIWc+aCaekdHsTDUc5GBvtCsX1jQiBO02W3pb956fi+wZcKEs35wNt9bGkg2ot1NiOLxjjsqsO61vYvAERbF4ISAnGNzDHF40UMEiACTS3D0uT+YnwN8rOv7ioo0IICrAVwDqQTQepjiWBZbzinBzv9Gs0XQiIc+oPkP/q3538Bjf291l2XcVkSdmcY0GC+wPjlvAgpyuKxqvOTD4IjWxOjObT+7Xd4VvcqAGJ807YNLE7URZba30xsCEZZXure+MGMq0AQ67YrbznNkBCxQEQrdkVQMJ9o0PD0CsWputb7wmsRowX6RaUF7DUQoPFrxnQts4bP5yFu68gRFaneSxmTDWmZmzZ5if3TFoJX431Z1HHru2eDJjztUegx1F4vlcm1rDjTWXfJsUsm86WDc3oCqS7726lXjkenveU5eixZP8DW7hXkGWjypgnXzyLi7Ob8KatcrImVfgbs0hHhe67o9KdEt39mUi8E5fRkuDmcfBSmnyvuyEgSOBbmZOmEcK/iaNUQ7pK05DBwog8wV9uU6V0lxxXDhSBOg/we09BzNjXly5pTY9Kag96IW1CJrJGwTZpu1VXo9lsk6oW2A/8MM4voJbpIAMRkkYohkV3tVov1nh2cHer0CVvoBV14hnXrQ6HyQcyX5iF3GV77N+k9ipgu2s+X3kByx7RiPn7c4UhdXkLWCRDVQ3sQx6D3JeznjNiZYwCCm4WlYi0ETBsul"
`endif