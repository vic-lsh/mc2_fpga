// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aM5lrBtr6uDKLFcSlrJ7LB+7WtAhZH5O/gnytkIf2KKm9Wbn3aAT0WCA/j1z
v/xu239W+9MirwoXfpcXm8BNhr3M75rCvemQBG1J13TSTitTIOGxO96LXf5A
JRgkqfXPaCUq75Djzp/rB75iZCw8iUeYkJyAJX755GkkXf5T4WJ3D1vY9/O6
ckt4nWboaIT60IBZOOFXitfNUDvMhu2qOPUyLhFkW05UeBdKZ6+V+X/hoU/o
8nq+KSSSsfEM6xoy1y1oOj292DNNpoaA9m1F2azK1umJI7o/sp11LEUTEnO8
JcNc1n0+CarLUqj0xit92gQZ96YUAFHFYnmQ9mYFKA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
co7NXDVdtNAZUP0bpgXfmU1qyh8k5PAc3DlCv0j/FcYVhWiADanK04vB8WZI
/MH+m2HGwXrh8I+J5BbxOiqSnX4IZHjfR/vejwpu9GvE0hTR++7vbnZU4WO7
H+NyCJkZ1KDaz6PEad3mPOdPSFr5EWwmkE0ESUHE+FfzpM7TNkMsdMIEI/rL
YViESgNLro/XEjKyGupfqNKXUp38LasBnvn68QfjxzEHg2AaIJWY6e+22vqo
L0wWKfmJgyeZa+3hK2i7tytdDUcrrfhbP1X+Gp1fYcJU5gJM+x4YdLP8qrG8
1ZWXDh6TJ2hUbn0RnmW5ah30AkSS9PK6e3CiUUmtTw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aaenVfkDqcBa5u33OAwusp29fElLvIec0TaYhPYEWCnrcWRlak7cEGEFCsxw
9b0cTsc2E4SqIhZdn+/sIV+X5eL0Nez7hof1O51Wyz2DLV019TJ08sbSzvyO
90wwyrClaDxVP1g4FyX4+3lLRsSciCKAac4ECbnhZR8s1DDZ9/LZ/q5ihaAf
QIuodWqxa0e78EgbkbWcI+iSOU1Qm6BoC6FLZ3pYG2jVC/KYomN+jZoQMtGy
WNtH+785Tj0tl9IKn+0eSYO0Od2Z11fDqzPq0C68WkpM5CosjBcrabfL1dwe
SUYso0IISHG9rMoh/g3xlTA5Slr4GNufofEC9/AAuA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BhgDdEJ46qipNRtOGBuXK33kqEGIP0EKe9TtwcIV4tWy6X6x4q+ZM5z4DSGB
c52s58F5HqBpDHTsuibX3VKGVGCvyZI8shFAqDj0cKYNxL96R8Ykq2WGdfAE
ICwaefxMsrEdlLFa9klHTcSNlh0khQ0XdV2ma2sYliJDqRo9HvBKYStGPBuP
Aiy4iSLswr9Wl3cI7bmhOci+noM/XBn7YdkXNZc2vkTTdcej/zyT3r48gWrM
cU7xM79KQEAqBx9/hz5/tkKiw8/ZSttDq82FUuc6OtVgmeCx/RyTpQrFc0ON
bbBYFFQvnswXvfRVO+6G6J/BEpalLtnSx+7JQEdy5g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Vec6WapcUFVuw8+R2Bl+lZ+3RXdZNq3MzeOjRUcTKiqF7ZmLwV/2NjYpcqZp
0a12b+/bS8UAqBJJ97W7PhJ0cf+XPBfVmKj7jZO6Zh3msQjJs2WDayZaje2x
dzzLEpQmQrxnuguJ4t56HqX6EFkBXjz8N6JnzZCZhCI2xx7GZGY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dr4EhEizCowClz0w9TUgksjtyHQj0djRiglkoQJgpsUnUIncA/oT6Fxn67GM
MUQCZIvBggR4BP/V/ELPjEU3EyTyaRGFi/3O4ECJC7nEFhrpzZmtYysHpOQY
UnnDfBqE9ziJPM9QTxDRB6I+cE+st5MsOpDZptsWXT+rUYX56d9P0Z2giPME
PnFfsBpnGt9pyMOaPb8zzbMLPoAjY0iMcMuoq4LcAzOIMr0CY1J240plMKJl
SWjxVMDpGJ7NwlCBVat2TmRTmvVuDiRWOXRUsaj2OM2ypCmEmxUmL64+0Zgd
wwtDDhltEI6v7DQ4PKHRUAGAz/LYUTJISfaHX1YsX16avbMBpRdFJ73+Uyrb
76GhWEopjMjfAYq9+VVADAk3JVcMNvKDAYfYf4wxD2Cn6Qv8RkubGcTsPmvN
Q8DJzVVXGVSb8DhX7CPvcDSyYrSfjQ449ZmIL4w54PC1HQt9jEtnxsz1uYyM
GANI+VZAh8XQrtbLOuBtU7IKpeFswPv/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XMa1eY6akALQVqcaU2uGld5hmCX07/XCzIyYc4sQMF0uhqDFAKb9S7me8f4Q
yn9sILUQTJoBaaHbBvRDMWCYPAnGw6RYGByFYc1RH4IoO2gk+RLLK6W0Fume
CPiCeyU1yynJVd3BZNhuWeYaNsr0lt8ZUjMbf3d1QRtPtqZPS2Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oUVzdOHyMfieXmJOlgBUKiqFte44f3D5lC53xv4XK6zhaUHHDFTJNYCdRCYj
K5RvJnVQFbM24DJ8Va3E4qndO6PsHQURDkMc/XgNxzc+QK/8WY0XT+WfyNT4
ONCpxDx1T6d+NWD5w/rLNpMVJ1854wYx6hKBpHeMNMbI4SpsaxE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 29360)
`pragma protect data_block
RsfVPYq0i7CsZr0HkYBc+fNod1uZJoGTHuDxIUAhffUEIoS69Nz6n82ASybm
iuWcVplLBPp+z1WhW9gsI51U7rQTEKP23lbyN9nx+q/kwXAjqv3hQtqKrG8R
FKjUjv9w+vuY7KTKPUSjrfJ5qMAhQ8BzykCe0sR7Z4Yqc6mkS7f+wIXZ5X4y
Hjq/F8tR8qmGiSk1XJJOqG5izgQna2H7J7Do6pEh+egvrHdyvXoZUNNZwLf2
1oX3Ra9XztA7KyLwodBEjJUszKmpxl+oH7f3JaxL+CGdJ4nO5sKbZJeMIPrA
GkiD7kQwkIoq+rML70kF8mXmRN6uGf9NTK9y9vzw6ASpIdpqwmiOqX0LiwiQ
XwBsqUXIXKYMCZH5hl2rBJRSQz26qCzn594Lf/U0ixCz0eCYxFNihDz5oCXZ
2YFOu1tWwF1Ygja9tSGuUoORpmDPc8hUeIESmlEKTOW6iuFcAKbN3Szbfa2+
amWkiV26ybtvM8bU0h3sJe+37Q2qvFN1CtyQ/y7sgiQM5c4hkBGj5naaGv7i
Py6e14jlfkEjbQJpXp5zuHqOUPrijZFMkH9imK4feTvobstR0yg81LiHVHlM
mJ5XsnymU2NRucnMJzX4gpVhdNNwfLXQHIWG9uWDr70jJ59Ms7QkVfilNfN7
z4B8wdxb32VgdIIkJNNVpiUIF0/WRsgvXohEyV/+iDpJ4Kyxg2DSAW93m0BT
bRUA3KAw65s9YnYCrBp73HPcv8Kd9sZjT9SD2KGI2AMNYXoqcphmBjKgGPz/
uKyl7kV5eUHdptS+aND/GGkO/kMNhOiBwd51/dVfuGe64mo6572LVf6qVFNT
//XgBF52cLbYXyjtPGw3jEF3OrtKnRNzq+6Jre/PUA21NXqNlsGDZcnkXfm9
nx648E9kN8UWjGv+6Bb3Wn06+SJ62RPwdLYNfmWT3pk+VOTgytyP4ix2SpW+
A8OMWK1ssIC8RteGVxm3XS3/yr+xWfFOwxoWV3n3YL6r6ew72BNe3fGTZyX8
hIBvS0UEs4K5jlIUm0gTEvoL2wENHwu6gY2xhzMoKl6fFUc9sgcyj67wDQFQ
XqAEtOsC61VktEOeGxGbbNqRhiqV3P/47wBgdZY7kJXg33w7nEznya5LhDEx
NXNwd8yTMqfH3NJ4g1LXHXfEzi1Yn81/dqhL9/7HFXrQUF9LsiFwUkFWvags
q91J0TkqFl/OZWiWcT8j5TH+HVICL8rhSSVFGviNtBNfyQIpbK19TAR6cPTd
q4Vdu75VSjiZ/cGA31F8zVJlc+p2sp/fSwUUFi0X9VCqduxXatbLQAZw55Th
VFS7/H1iBtvTUuOc3oaYXDwAejJoSICQ1M41OHwAboMiQUzbpql45rHg/exw
zpjKsL9NgkSDcVRDlkRztmtW/BAQUmGWUq0XrxZSs6hJJh4cfNqul/V+GwL1
NZXSD/+ajEEpkrfkkCIzritqJVy5A6W+JivA8WsZYuWdI7txAubkyvaDPvf0
zbfiLEpZo2j4Qx84GZIQb+iXEzi9jsa87CCLQanzLbLSmT/MwoJAs9jLkdmM
x6hvcoGZIs3fM1lfkbwcZYllf3a7+xrTUfP8SryM0Qfs3HXYfE1VequJUnp6
tHlknqpvrrBsxrYtjxUClkogpyNOXyH+8V5QFTY6kXjrRJQVQ8EQlXg7lj+0
eIH79gNN8xX+++atvXCFVVfwnjtdjMsQ/yNxO0wbI9aP3cbJ6K/PFr+jDG8U
nqaRKDLtzSVJ2mjbuNbeP56KDj+LU30uD6+zkNRKYFbZH6pfY/Kq/shs7V3L
vxIkcfLVjmC++2pCmnWt/mTgvUaEomIwPpiAZsgFQeFk4GLaBqv3ESvpRFhm
MLYqfQNWvijfcBEHzpoQDmOrcOr7y6LpS+JBjXhlz+XPrRtd0mEH1LpWdCQ1
bASzzQvPmt03QArbsUhk5HlHtLIPQfzh8mKxoUqVg47WbvKHssktrHKuKyYn
OUWh54WmAeRNUBNXLrcnsaAF2Oc/vfUtcfJIb3ZQbHzvLGi1VcyOpBrTjSkG
CLBvtqVUs8km34Axa166Yzcx35A1ahhRFNENVzc/kvmlXIM6hvsNhxzXoa22
nq5QEGDUq0oqjYy9+hObBCDVlRFWVHUbDoaUSjDO8XxELytOo5QAzAosdNEA
st+o3QEqEX/bhlzhUScoqRuC3ODltVP6fl13KEXrESBDU+IU/QOTf4N4yZGD
x3xFO9udvcOZF0c5Yu5PLvOYzPD1hRX6XVteTaQ/D5a74jJBwA7P7Duht7AG
pgv+hg34wBCk0+xnKbsGJd0pVL7ZfFoi5elvmzpzEQNXIezb5gh8p7yoRWZu
jLwfyu/QIJJVeEaofRleud51uOh7Esp6l7Ccrr5e9W8q0sinytM1fbusqI92
NasV/EAAdivZFteyFd4a1IubRD+q72J500WGqRJUXUXfp11CKyZy2/Xw4EKS
fGq9JlP7PmRZ1Mv7LHEYJ1L4W8cmFDlt+kFmaSX+lrVZaTM1EmDL3CPprp/N
2icJSYdVYbE09VBM5q7kBJ0i0C//bWLFSiwFldnyiihCNMGDFWnS1fcGLqmz
DrY7s7nko3mXnp/wjaOLJyBjNQm77blBtZ59ILuTvpxevCG83c2i8Wdkzwg7
IrChN/i8XXMCKJOvthYtuYf9BbIHcANwduS4xci9DZ3bZnMw0hkOzHTKYeiB
vA1TjtlfotCd0KRGTBOAkCCYm2US5kx01goi8TsUw2z7hyW8H4AYDrTpnoiR
nAT0gl4IXdeaFHw7igN4FKhfdT/DpIFVsCVFmzIDaoNnuc4Kb6M/XAwgtimm
g+ffARrlBLxWqnEUmg3XvMIAHKIfdQeUQPxe8brirD9j6GHyhe6dNBrlxwS4
WRveihuh6MBd68Qo7QHT35rJ0L3zDIZANAn11slU7L3UNEGGqzu8RzG/vL0w
kaGm5lDRoccisufdePjTtlEjbOXLP8VJ347RJyrr0gcQmXcMF/r3NSe6V+Ui
sU5WAQr1fooLcpzxs/Y9SONU/ZtDfqIwhqHv/aglWE/n6LLXBFSKA5OlMJC5
WgCDAYKcvZmhe40O2bVJCc3O/YCeu2T1jtfx090CPD1mPZgT10S8NrmSz8OR
V1gWx0/Z2tbq+XbXMcEBgqneRA2vK6racVuraSdvBlEAlZwRfzZrCgzQ3GwI
usBXygtWMpqxH9846zSGL/W2xpuwSQUW8lirzo6DFyL02s4pedrkAsVChgW8
bJv16S7btjiCPee0j5Y4QhPVI563eN52e5plN9R+rEkxMFGqqQcsyNcXLnNR
ffNQZT9BM9K6aviQiDLbdWuqewpMJgZELCSh0fTFQ4/0cHvV5/xgz4wRs4wQ
ABbr0VQauHQUp83aOVmmchPzcIhIsmhxRDSiXA4im7veMWPi/Ai2uM/4bvyu
lgc3qcx4K6rpBfkccK0txpL+1rXWh0VpGdHFO4ITco5IvcW2YJW2ESFbWVPn
wcR7uxBgJs6hncVGjalusanAnqvwstej/yjyNsrwO1DrHJll9g0JwVmrVnNS
mk9g1mgQlI6ay1ZGrYyIDU8087fBdKN4PfZasFxDTzzNhsivMyqOmhygktSM
ZGmgubIHf28HVoXj05cQnVy5MNFO91O/qDzDf0ywU7V8WeH421qEiUWqiIzz
fHTmOUQkWArfC5LD87u9D31s1leBL1H9Koec4BtMdC/3oYEBCPe8sj3P8UdB
U3A4lBHxCCJUWb5LDJJsJyyzhOV9NQp1tKnWylwRcPbFO30Ws7gSH0sD+beZ
crcIJdgsTtlB5Ucz+iSKqubUNAAluRQfwBBG5r+N3YtaXlJltcOcm/ctkE4y
dP2kjJep8gWZwBzZtRLNhT++F+M84e/GdD2aCVgrvhPpxBDCC4cN3VEGovgO
b6IgMXJmSY8ACqFmMXyrDqdfPKwZNKe3m+eWDEvwVy7MgSLeL5bzNsZ1p7Mf
hmlnZcd8eyOnuRKtsFKBiD+PVCCqbwqhoxPfzXXnxc1Q8vuHoRl0G2cMNwCi
W2rYY1FoGtV9OEQkCDj2mo3sGbqm5x3olDeVBkRZXcPdhdSzAcnPXLEztvZS
Rvl5E1aKpH3HGWE4SWbFMKyaUrgMb42mCHy1+w1w8DbN+z+3QGhr6c8YEUhb
EnAH5VVyXuHBMthzn8eTOjMBbbOZQWTJNfhBHsnpHV9gEkMDeCEGqa0NnIPN
dS+prNmoe98ovm36KU6nSUNU2upPqEN5DP1QSYZUxTLPDXuF27fqVe4Zhhmw
TTPNVNDwxD7jWAWkMfQGOXwmsoO6qNM0g4WjB+9lbaVTUD1HJuyJY86M6evF
PAGXVi0AXS36kO5Kn+rk9DpMBYpG/VHtbRvX4N/rSR32F/2ZpMFt7F7baawO
OpH7gd9GNlBN+MtCXdOjgHseA0EsCmwrK4f9SFqc8rEfaLPciZaHwm8EUWP1
HVi6oF+gsaHG9hkpzmv5PHTE8+hL9kn4WkhYNEFYg96ZQEAZoOjDuT+wRKdB
9UXsVxNyl1bd+Ow2r6yEMIsJsTvOBl16WNcUxSgXsLUySZvW5AZ+bj2UQycD
BxCTCjTKpKZMHvHPNIY3H8L7OXD7XZydXHa1H0KRarqHjBKtnyP2YrL4QhRO
czwF1ZEuldfxgIyLzv6XFHdjlRxHdtpPYMdsNfEgas+DQg1YD/gpPwJvPCfg
Rm4kjT32CdPX9dlfMnLgF3FsLs95wEKt8l+FupPjGf48d3l4F99CMg/6JWmE
BqTOF3TOsvTogLFIkw+mdS2XneWQXboDwI8lDYVEAd2gbDinrY1dAODyocxB
/7sa4rKWGqrebDacq4t5V5dompVujTabeCd7DT4dJ8fUTcF7qgBVyoN87Kag
iXjrfkWI1LHU4Cs/UIePb/zyXzc1aSzDeA/Bk9tUHYBt0PnmbuR/WyE7ANRo
zhmUStGIn9J+phC6BU8yzPXebN1s9+9wwkn9HAwpTH36/pFDt6ACOr8ivzzw
PzL8Dm+eDjz4BmMsTBwuzgcXmty8WDruRcN/6VOagx7spNS5w4BZ6/D+nSIh
9Uv7mEteYfNbjDf8yd0xF98fdwcIewUynXiKr6BzQsQ/Nq3qrRZH6kS0/J1Z
Hpe9P7J51r0TYfllgdaXiKETxx/p9q+Y8uO3pgVU6ilgHMEmdyzQefNb1Do2
sjjDo9ggaNvUdP0XOAjq5vjs6gmgdx5h7YI6gI3AX+UVKRTwps0iVeUcCnej
+qclD7Q9qXKveUzaI2I4UMFXacxcf7xpIqh1g+Q1W89f0ONE0Ct7CI3uHxnR
0cx/5MvxzFBTUsz0i+X4GamEcwAFTVeFfl4cjV2MHwupNPOJWM+lkO4ra4Sb
qiImlyA5jIW5LG8zuqFyieNhU3VtWonw/rZz9TKUVWMcrKfDJMJ4FgW3uf1/
yk07P8mFzsyKvr7kgpJPl0pKmgtLVrsrPnS82ku+ls5Nj1s3zVX9yM8Os4KE
Nv/FGHFWrEc16Rm2BjqdBv35f3/HxSMaJOw3AVMOcocYXz9AnGagq3EmHaMy
c2SUc/Iz7UFAnjBw+Hch70di4ale2I3KTbK366+jpk6fib4bAlAjO4jqtbY4
odwL2btkdEt/GHqPxXFpIrmDJkLyPMCKUlnZE3/OA4X0bx8mBiPcFUH47iKR
fIjNOPN+LVvX36dcsihj5MEEJ/wJYa5mmCxMPbJR0gWYvppcwICxnV6IJPYN
R10qZAMdKJOHW3i4p2zyUZ7RSEVTQMLvEsg/L1/kuboJV40chh0TZNQz9vzI
zODlkYSXAB8aZS5n1vu+6cWMs6SNk6KwV7YxAJ8L9Yh2erfHkxWzL0eP7B5X
2ogJNap31s9dp3Yd90sTak89BG37700Z1vPF7iaOIsTFBgezbRWiZcyiGIIW
A3/MgfGzq8hDNTlrSk/VuMW3Yhn5m/uhRi3U8RQW2uddtX+tFlxhwnIE0fwg
jm+TBzO27ZP9Lr4PS8mFMQth1d7WxLhvsAyezQR/4xULF/lcXlzUew0InGaS
fMZIsgPP4SBP0eF8tM8pWuKbO3ehjMWUxM5QtPyo99WhW/bgJaPTUnfqFB5E
VRcs04ty6qBQRM1+uuuRfMLmjpSUq1K7gcH4iv/PtK8Pa4M6Vb03n2oNWoo/
XPa8dUZjNU1Wm7pLeh+FzuQp+XEaczcXLl65hDaIY3jfRVWJaUA2IA2UEzTt
8w/TIaFT6VVH2AVP01+Nh1iYbLZEjwSrGQt0LicwKAX5Ifx60Ug7aGVpxkJE
26UkIn67NMuKdIpygtiyCNwDoJslel5zFt9l4fZ22wp/G8MVBHVaf/k8bVSn
LXjxj37aMcbd+kzvEFfqtY3/A69pcEUq6E7Ob6Lkqp1lZgSld7GbbXW6AnvU
jdcOX9x8ySa+7KA9rNSYAeI6c/Yczg6IwBq3mXUcEOWdakHcMaB2A8/1Xl+o
y4VKB/Nk+fDLIvn/PQw8VDmQ3mgJbm4nYAT6/D5biESHLMmFJq1GPvXklviU
5Dzsi/bHz1GUn2PQg0ELytxOGRjkXTfXoPedKcDTs3YY1apI3YxpJ4R3xwI0
0aFXVG1evndQNMC9aulBAmjJczf8fHaRad6BvdT6HKAsw340xv0dW51VZ9oZ
EE/cSSolMxrnt+nB0ul/Uw7RApvacmkpxP0U0l5stRWmTQC0OVeIZYuUNg5w
TENGMTkSEYvAsQNUKdQmp7kiyv6YW/JFWO1pKiHW1DZ9RF7JuLMy60slfxbD
KVmVo8ABrgbXDuMjWDQKFu/cHwId5TZgINAzOAHZSQn939zBDtYvaMOLnWGH
gSTxNhdHDEnZAXuZJR1WRoF4uWrwvWesQtAMxE/Qzw/Weu8NZaTHIrLVDgWY
CPfSMYAe0NKH2+9UIP1ZrWo3jvCdLJMjZxpWf531h7cw6Ou+QKIkviJsfvhw
8Pz/QosdtmMYAzUOFd8ie75dYbVn1KQ4wcNodyBBHK74jLh/IfWpBVlziU+L
wZyROuraz4dpQ2kYaUXd2xTNTLVad9Yt2nu5hCuHg3Ceu+YY+PK3DBsWcktw
BNhqbAexq037TXjuC7/GtM0AmJRVBwauOT6HMvv40Jm76ufz7ztY8f2fi5b/
G1K8OsAeOKjHQTF9iVxnvS1l1dRO8X/Z2G32U/1RpoWv3MexX7K5FG7kIpC9
f+ZW5fepzwzxkOsgsp+nV7MyaP944C+uuwsFooFFNcVW2AnESBpdElwkP7NL
VQADkYf9GY3Mc4yPRW7xruYf+da2999a+/44oYwdnR1Rl4tXTcIjgrYZjCk6
x2aEOENElesAcUy70e5DzavX1fH/TsBZ6i3+9iITA8I7iXCvMRy7YZ5fY24J
VHdB5IAxm3D7YlZBOR8S2Risk6/jvRC96+qKhRr6smYYt2J00MSsCxwB+tdl
cq577e+V24TndIyUpLMYlyS0UcSRIBGXrOP/RSFcgW8JSGWh9lECYMAWQiKK
7T2ZEHchc3ldic0PBD0p1YNkQ08g5uoJvHswKKZ01PiXgQ6ODRm9xhczKtl0
Jeg8hahjobc9AuJ+b8G2PcUhSo1zNSqKYqJnduErB6sm8upSQaC1V8X7Z1Md
UxQr/FIPKBySUxilA8J9P/4a0LaflL9ZaU0shhru7EkgY1DmvZ1lov1nJin7
NaPbOTojp6tuGbHCcAqdjRnW55Q1ZX/iMlg4A4bewZpDc2AF/YlNJEW6ascp
pCMZkixaLBClcCGyzRBC/rt2wnT6qCz8f+PI42tYRYseNYdZUO/rOK2jGL4T
1mRU0sLpjO0BkwJ6pyv+amOeESsvVaYD/Y1DrJAYMg+OAvn7VYvOFgBuy2FS
J7r3Y+z4HBMugn8KYgLf6ToD+jaeltsehh4pCZ8y/1Iv4kvBckejNe3l9DN+
t57ZA4+d3bA5UjUDqoHWA8MmtbGGsf07FXXt8kSnR+4/iaorTjRUxiEsffqT
cT9mqQoWkEr3RLIg/XWDc4M9JEzusBH6MBkBDHkldT8b8S0nCC5u6NKObMOP
z+IRPVFo71sQpULjXyVjar0rq9wdh/3ij2aJMD4/nJQcITyPDGPpWnoS9Fts
pFO0hzUgJUEhsc2rLlKPIw7HqRSw9SthtYfTbBZcmAr8r8CjjHOjDeY9hzmS
L56DGxLrFFE/w7sSDXw1gup4B8YytfXqjU5XHLnmMXEzRMTvroLuszzzHQbu
waVTNo5KaQJfF4I7kTkLbZFEwENC18eXAyMZ9ljeahBX7qX2lXQIHTziHtXw
xHi1vzON7QDT5M/G3rTeVkuDgHgVKrJ4PK/tWJ3OjrKLSDUqBHDpxoDdRknJ
8Wvjik6dGOoUIHj6NKegUmlj3EpX6ziIjublnQI3Jcv1vAOFLAOpfqCH0VFk
tOzAR+BSDx+fm3nTaTgdG9Cm775Qb8Unaz1TZT0K1sKoJnb5ZcPV1FJaIM97
7nLnHC474p467rLOgg+zABgohW3Obp3GIkgmiOzitOHPPDioFX5OHZhnrJXK
m+1KL58rd60Mkvmuygx5X81x0uNCqbch3aseyUAgnUIOCCnPYVfkoLZvjDoZ
3oxFZqXdFgQiJzCpyxMNI70K+Gu8dr5iyVatkTzMc1lljA+BOmkMdKBZjl7G
bWUqTK6SPkgPPHOmodTSOaW3KhhBslH1+XtseCHP9CdV4vV8BY7RH985tEEH
qP2Z73pr7KxUQUGfROlcYC3SY34Kk447K4YqBoAuZgMApmaS8zDue4+hXlmv
sDLM0Ins/YfW3qeFyAskpaFfrD5PvR3d+AO0/No46qqyyFwxBH9pe/ROsJ2R
w6915AgjGbtDRNFKurDd7TuXH+CdoxKPdb90++zM0cBj4oe1c06GI8PUIp+O
12evgRbmlhd/SAuvkfD8pvW9G1S2V0ejiq44ZgKf9VRFwM+fLIvrt1K1+oFw
b2j/qR+KP205nnt0wPqfPB19XIH76I0he//bH4GAcrMvpBEpY4w0bCOViySw
6YpQEuCiKBYH+QD6o7iLSa2/voQNpE2Q/Vk/3FVmIjlnq0BLh0xCxjQ+kcLT
WYvTb8+PPd0Z9Vc9z2FG4d7zo0KI1sscXS3f5dz3UQkGiZuLU548AThxfI3y
ymBXItdC6FH6NLQjt6ifCcl/C2ClaJpPIHldmI56nlr+NsLmK0/UA8IrHHOL
Quitadt5rZ+wGNIm+/0cZ6DnVkHJZsLuPsRMM0MqaUifw46NvZ7cBytpDCoh
f3T56hnvSh/CV5wHZEuTiN7XK/6xaoDZMVxJEI6KmO0MtI/ri0GLTBIzZLI7
3sn/diL9uHJp1H/o2yFv3CEAAazcd1EOhi62a57vBMX1TOnukjR6gyZ+IWXR
mGDXzO7n06gwFvWwyrQ7gHNuJkea8fjwFv9jpJ+mkQrGfF6bYmExtm09maBR
NUMUXt+pSe9MmJBRKcpA0/idugy9bfAWriqLogTzGy7X4/m+cUb9XqpsBwf9
14fRtJCNF+CE+vxAj4tJjdoKs7Z3ipBwJ7VnqLIzn8tkSeCnmtwlIdN9iwPD
jBGH+ZNmsi/wlXw4iWur7f2mnxymEpkGCypvHX2WQj7DkPpQV44+Yo7OTVEi
B6DSP/NSon6CBhWxvjiPLaVP1U1xskbbvEKYTggNOxhnap64fnkbLt4Zov2r
lkjJJSeVQvc+KlwnK0oko8zPkc6YutQELItnePGVwKNz68OJs0oOe8Cj6x8e
Yb7ZygwuC9pqAGz5eBwuv8U/HHyiLy0Mmez5MFgdxxLb5E3hpRYh/qey18mr
XXn5Ki6G4/4C44JJS+IImphS2k2q1f/uHAWwYABpOTF7fugDj0SXOuuFlp96
nx/ns+4X6FNn96RV7SF9PoxG49GWJxnBL8HiJI5l9hyLp5Uuwu/C87h0t+J0
MOot/LPAijuED8hGUexYp/3Uy/CR6Y8nxgxjiaj9qYueY/+NGSNvfeuCnyY9
19JkwRfVRmKxBIjAb1FU1hUzM5BUjtyMdGRNpLr1DfsU0S/jGuZqVvr1OenL
Lw/DbtqwubLa+5l/eLuNnvnyVGitGWUsLT1YVwGZX4Do1sWHv/LIDiM2kQ1c
bjWAjFHgmr2jTUvp8lI4HGPKh/Mqmwikq+heE7of9rXt9GkHP+zplN2Opiyk
z/Bcrm+co6iWvP4heaiSKROelpsX49IGMtZOKSTmsuibAV5M9fL1XayPhXvA
bp08eBBEjW5UXWgGFTO+jcl1HS3283wAeicLx6TdtwINXSvxoFEDN5tkmodJ
5hDrbaQbBqnpUtaY1ebbEj6Z4NT6Oe2o4DHqog4Hip2Rw1daTYRJxSAx8pZ+
A1/FdidioEy9k4Ujai+Rsh4cB+IiCe2XzA4IVzlerKdoimTsFYmET37YyFER
RMQZb02o1hC5lcICE7/Gq7Q5nRhC9XMI4GUgqBwidCAHwQlP72wmjCLW3wTh
87lhN75sFvLwtnQ3HujZqWAWcs/+78DXXayjt3tBcPVYIwic3XfxZa0FqDs1
Kp6RJIiG+wwIK86uMvyliKLnYfJm10YvzSYWppKQ83CrMdIJrg9s0DaH00Qs
DzWIg2jfiTjDBu5ai50Y+K7yszFCaxBQp7yuGL3ztfw7MwNqa1YIvgMG6OvF
QCdTfRdWjyCAzENayvrxHrqrcfxTH/BL2izt1DFrHb61hl8Z3J9a0W8FaBh2
Hf0K4JYbIoddZfRzjawCGroi/zU3PMIW3G4A+DsgmSvk8lXEu/XQicNoQnvX
QrxT6SAkjf7BAF2jYyISe5HU2+Aqfwe+Vs7njQ6riIL4J2Qle6XrXU9r+Qbu
X7nJmQzEz0Xc+5PRMrRFbtGT9M95jM7Au3ZRr/J0HgZiKpRVzB7vNulGdmzu
xBCLVE2m5VcvDir+sqZqpEcZohQd31jKPFhbI3pEzHje3kVjzcGNpJxL/tqL
thWddLNy0wAJuSgaKuKM7p7f8nYq4dL7ynFRyr5x6hEESr/aRj9aaa0VFJOK
zXpfs4RfFpaxSBugNtIqmMvR4SzEA6a4hgFHCfIPzXRolu0mtnCBpGFbnKBQ
rziSrrMQrC9aBMdVC35en7INWzyOxEEuC53BL1+pA6SDUinFhZ1DsIyaW5iA
khp4iHNWCI1O+N1ZbvtwGhZyGn/ET07ik7KnrNVKUqN0dL21uYKPn9/xTVfU
OEkwQUWDyCxVmbNffBGnozbDvEHyH4/KZzgcLJB6d0wYceBNWZwMheRSAgS9
84uN+DdRqvsxUdEEdaLh8LC8S74FUhY3HwnvJG2hRv3mMiR0QVfx0sOOI60l
TQk4wmWjoxw/1Gu2sEt8HlyjCKBndHltrTuqimStnN3Y3HAjWYnxVUfWdG8T
GaRyeO/NzfZFKfBa9NjY+o1y/ywkGLoEEC81A5j8xoMIocewGfY75zdHxqEK
t9Fy+e1sPkhBlXs8nx0EzqtW+fYO3kh+f1Agz93mZcTtLvAymKAwCTD20lXv
Oz2uVx4+0PiSgMJF+Xe6hgirTrxmwb5wumov5fPfKCKX+0pbw9Z8B4glqA7V
ks6oL+n17As/F6j0YB2OvDiFz3AuF6uHnacMmZupJCsF4tchrgOSPNsK8WuD
0vaWGcebY+hzSBltJIpUg1317Gxu1ypyrQNBu6WLQf6ruD9S7/8rK/3xBhfZ
NwPSh2GHCKJSuTxpq61FTMKMnPmc1JAAh2rH8cpGpqfre1eXqViNFM7y9ZmE
kS8tFhajrCEJJybndNYCEHnruaU/2IKsAHLryXkUyZMG8ihUS9+mg42Uuo+Y
YX1hl1Yd4bryHpS6qEu80iJefZ1EReRArRqgSIP7VmxtboFlpXvlwzG+ngGa
YGgbI1lEcGQgz3i68OcptM9fLcSOYLQnRWf/a0jDoGAmaN2ioTbsN/iA9dS3
95rHKtvFM6iMSTyOKFSOrmIV5DJVG93pzPdlD7XeesAmtcn5ZpfQ4CALBR5j
SBq708U/UyS9XMjM4gkzvB8OBefAUE+gBPcfd2sAQ8n4U3fJZcsW6kGzJfsn
U92iDed+LAbj4h7QAbAYrDNPd8zJWNN0/fhq+knpNr2IjbzAZIJXiq9R6NqX
UXGCadxj86KjZYoYTjC90IlXD+B8LaJy7Xk74D9weBHjibxrMso+GDiUlFYm
NMmk884Gfm6kt3ywq/h2883hB7B08lc8mGIshhAGwte4tgEevxFSY+CMuFUe
MACG5f9VsMWRABEkd4t0OFlt5lWSEy3JlTiUXg1lpCO/kqkLpxaqC07rPdom
h5UPyYcd4Dcn9zcSzc4yb5Nzku77Ue88VbvUjvWCWwIg/ZjQLDIAwF5aPcoZ
QPh00bYW35xke5W8YCq25EfIpDQHDKvy6+8jgEMKaNU2QU4asM5g2XcS1V0T
FvfpyrnLl68Q5nURZK7SpT3Wh7h5cd4Llcf05aQEEJQxWd/qXsVWa9CLOLFp
hzfi1TXhVMDbFMjSEaxePct4BOlC52UlkGIn5U52JBBxBBVnqOcHh9ISbL7W
1OiYfsoA+BwxzSPXSIIdF7FG7c1CHj9Qh3Xr4lRo5hMWZKBiuOCXHg7iP2Ut
vRgyxvDdmjdqUVAl4BNR+ysXQPL+rYTq94/18dU7Mu2HDA6cgHy+//iIgEnr
WxJFlvhTDAcU2T3LFhQ6Qs3/NjTGHYSouXSRWR9ZGjsWWHNuytSunmXI7UJk
h+4lDjlktbv1vQhUHQ+2+p4RRknqzHVFVv2xVsSOygiR7+48AjYcLUIvs7Za
i+tF3w9M3sFxQ8ETgVg/54ccQeAMBovFfGpgbb7LjkMUj8TggzLFVZS+IDko
eHuryrYKG8bq/XkiXOE7vOjL5HUV1T1KfTnfHmvGiDpuhhl2YEzpnWKkXoYg
ILx6uQnnYVSjx+EC9LIk1Y4PtIqx7vW9U/lAz1dAO5d+igtQeoLPhLHCv7ih
5Z1ed3eicfN7xlpweysSnI0vpqT2mEJFxogeQGABTGObv2luOuNa0iHfJO4/
unrZaGeB8+9rarDRU7VPvBQqobOavag3Mv4Z2VB5EQ9L2bgvmV+0u73CU7TR
DavhxKMcfMrb1TCbnXxzC19ho2uet4/no1RGtmxfoK8GtOUON8xo39ty/iPX
KrCGwWpcfXXjtupd1cQAQv76qqoQiZA3IT/4wq5okaL8TRoN3km2HPIctWsk
FwbFiQ4NNyNC238VZsRS8g8pmMltfr6uu9IRs2muZWP6taRj1+Aqfddi35t5
q8qw1+MPjeqExr1ZqULRfKK/bKqayfJLWbieOisJJrUwzBbyFN2CJ09FtON1
CPxSRoiw6INqSmhqE4ycXcRRw4UKcbifAFFvAnZjxw4G71LHZ1GaNT0JYEd3
dwXMenbEd3aQiA0XDywhIO+pOsE1/glOofeTsN2kgrH+2MINvPv6NezS6GtT
Uoaz3tPn/eEB+X6awQ4zjec/KrQUu74Dgq1OQpoyVyvpU9HRBaphO4wfCClp
niwmU6bkLod7CKwP8JRH+d+eJbetXUkgJ7mgjmIIREwpSpdYfacgyLqmcJ6F
sCSoDrFfNJnpWxekHKF9tglag/u/7HwqIvBKaMxGi8BwJ7YPYL2oVRPy9ZJo
vfaGtNGyLtdkdCQJYeYKudJ1rBVVrHaI+oOQXgyOwf12Q+z/iCPjMrI4Vdli
/8Z68iZChgxLTNi7iAN+gx++ulBtggbvMXVbFGSg1R9I4UZ8dWNF61LlDafu
6+QofidvjwtiJmzsVNFLXSQX5BY4nnm9HZH9J0IDWGzRGdYbK4APx0IHLCEv
ojcn9pSQFurVWhb3lIU69O5aAwP4QsawE9ugYY1VLFdrpFte4DkIcIJlf588
wVvTwAhmZZdCRkkvGu01xlf8u/77Mdnx2YAn73jaZ1dfKBDjPRzRn53VuI95
woGmTpAi3b5I+JtObauVwBDlKt2/fc3tg9l2l4tqqdw5mXjSlnOVviIED9Tb
WKF4mUUXTTH7JePokQXoPKFZIe9d/Ndvd65+JsvLMQZrXVVrTVLf8nF2QFh/
fr2dxm9zr81hpw+cSsVRgmCEZowUPZXdGKQt2hB8ImcsViP7L4kukB3zez1Z
6gjrHNirpOZXXRO6wnkqbAHQ4eVVa5HI5ajTFbBdbco95SuhBS8fzUXpc7af
Ba+MWJ2cbhktuyTHHNgkg8Tfd/5nwbtOZb8s7Hmycwroyb6KhtK+waB5Jk7I
TxAFuJrSLxHhrRGEKiNwH8GkwQMX0oBmvKZiRw7ftK1xDO2RdfzTDmuc5F65
ZtlWzC8KFsrEum8x9sbOp0ssnUF42ynMqmrX7BFX4HS6nnuZlKSW3502DexC
JZbrbVs6B9jt/E9JVLOX7niZ3zxA7vN5Cjqygfs40pTf+2O0M8K0tXhAVHDd
/NVGIkt7AMVd/6UCv3HhYKIm/RwKYtv8Dvu8JNoqlE7l7oTezuZ8LlVqpyWu
kwGo9EbH7Lc0ZgbLkUS+5hM7XvCnNBg5IAmNKoMASwVGTOGY6iPYH7w5dAlx
M024Nu+KuuHAoFwmCbmXwnavd3+H/Uc3hnb2BaEkN3UvIgHEoeOWjASLz3X5
ih+TCWVPR0+/Fw7f5hHWLXN14z2u7sp+S3RiRRV0bry/0mhzAZpVGryaaCao
xkR4Pm4nRe4d+CbhQQfN4mDrh9AqKz9WxlEt2B+DHbJyacrrfawrL0H6kGa6
sJyTMh65hfyQWkaqsv3kKFqjWQw9zjGaA/iP2EMSYAhjEixsRb+89ISbgw35
clyLB04Xag03AIO58E7n1qB6l9WzsqK0kPNSP4kp/OrjWtR3vW3t+d4IiOz2
2pHlFRL+iJWI9Sl/O/2oH3R1ASAfLiFBaT27lP/jHXycGBoLqussdeMkXJia
ux7+ChoO6UYyNLKvgUueXZ54iNfsb3LvEHMJ+TAJU2QS2cNHnSBnhZwYZxg6
ejhNFM4qp1l0DBVGo2xlqwqwFLF8CpZgN3kdiEU0JZJe1Vj8w4p6c+10+9Jh
tDoQS0NBRNdHNSFcoRbc57bn3ClchuIFVWZuDmK1G1PcrwLnZ4qenYfjHHjh
VrmMVadaWFtssNSmDN9kD9PbtF6WLJFs/FzdRn7LbNwCIPkE3iXdOUxxnC69
2FMQL7u04BJTdAObFYdUesIoEuQpOccZ0w9rOkqL9IJF++gY1AsOqg0Dygtv
LnnOmxG02H2mMj3azU/6OkwRudifbKYNlBMe85JGKX+ULMnwHKycXHJUMSba
KkCCanXBBBcwJ2fKOKbwRd32RrFpEOxCyktK/WCj83Ll08ZOZeQiRECA7pMp
HQQQ4Bg3YemcJZVNLFs2bEafQZLEFhqmZC0KXjrG1Vunec4UsqJAJQOdCRNu
Hoddwm1mWEj6QDwQ+jzx7/W9bKNKVc2HenT4ZL0JdAeFnb92AG+ovBeWumIm
hGlOeIKwYF46HIywKJhmMxcyxOkOUwQf6LjfWW2C8LGFsmf8vhxTrfA7/olm
H1cBHG1xhgGyiiywqhOk70RaT/84C08G+jVuVQ648jBwLbuzf01xLFzEQ1/C
VfPxVXIJhnqI6QiXqF/VjI/JqYz3oV/djsgJG5xyYLbaDi0aOIDhI0lyyuqk
9rjMwrG/uqY+plAARO7zVz6IrVUBp6DGVYmxH+qqy73OjP2pCIOBfkhgljxG
Pxrir+oSJ9vwncsu2OYlViyUHild58m4DEzk5uMwVO/S19ehT3Q1JnzuSHHJ
VCWwXjxwtsKD4lYfdtpW68Ww1mrdLAvYi86Pa5NuQAx038lKSl07dAkfzaar
+0rH4KWNr8a3/q9v49tuErZ/lo9hnGQBOOFn1Fy5EOjXuxdllhfvt1G7Mi/F
3OiycSTwZ4IhxscJL8XZzkmCafM25FaIWWc/96OXHsEJIoENe6aqnDiobd3s
ttoYz/5T3iOHFCOSL/qhYHfdbVfTP3T1Z7a1DdVZV5epWZCesLXEVuexXGkj
AaaGj533+nvlANa3vLsZ0/J7hj2BWh/ogbssuBTex8sYi9cTvuCsmojNZqro
gjuLn/WiRSUc6wlM//kzu00Pce+a/UND5SorbEP+zsTbvem92b/jAnoLSER+
rXOo+1/M1aLDq1nXLdYyI2pSQo+s1t9qnbeQhyIDsPy0PGKBVhIHAxYN1VEq
dq9+dRbczrNSOTYx+bZycNDOLXUbsov3SfKJrQpXpGCWw3Tsm1eIqaiSBI/i
f0pWuwK3Puw6UlRxLykzjeu5BOQbhIqLFta8DRVAOeTiUDWTE1k0XCJ2iBFy
jKxzfuR0l84hHnCQ9KFF8lZxjFopjnMQq7tIAeBn8/6iLgP/fFxBAkG88Ivk
VpYeX5rQBmvSVBA5mLWfJarOpyiUFT3CPKpaOE31EB0OT3QjI3Vv1/pmFUk0
VgRhNBcEgll8kWZOmSXNoaLpinZzhzwUqsYgLY5quqZjaa6ZGGjvXat+6wZO
9DmIEIQ38f/sH8TRElrj6PGyzywPFEpqCaIT9sgVBGjXKXZAmTGO8jI5tVeT
38kKZlg2lv8w+Nf9igbZKUwqRSD/x4jVsDzfYNXjYCfHt3NrUyIYB2P9rQY0
3TZ1OH4TiM1YFD08dyM33DBP77syucV9q744JGRJOta4iQF0af7DeeSKgro/
ENbqCSQYz/PVs5rIP1CiZNQWI111YvwFK5YDVVVTo1XsgD5dZlgaSY11/1Iv
N/U4DLIvCNZQLDsQMt33GUffOSQxed6OtiVGx1Fhg1rBYyljqdwJVExwU3TS
ui7epEnVLs+7y0UVc6GeO3BZ1gc3SF8DG7TmG+vSXk1N6YfU2HmYZa5OqwO7
5mPRjMjlDUPDiPrQflOxezs4CJYQZC4acM8gDLWMzPc+pMLV1LRZQP+Pr5/x
jwC6HNlbbRyuRsfatWoUqcXgGCs6CgOATruutDaXeTuSSVJz9eTyh+oPPg3/
wmlAlPX9+u/qDpMscz5+YbhLNGCMrZMBTcIL8qYDYAOyXxj0RBNzRqGqCTmF
JBMnCWNx1KK17ybAXJO2WCJVaxMNJL7rncLz15k0Lmh1nouVLSFUmf7pUWWB
74uGURRFdMPYXCjpAY49EoZIcsuVSd5Yuf9KDLeqBGimov6nzzGPxTwj5hsG
LL9MM4RdsTf/e6ajkG8JuWH4TQRP7DMLFJChAPXoUSBTMVvCSuKxW6sYnoH1
Stw205jRgtWQ8v4GToo9+gx6OEsvJX56eO5pU5jz2A0GCVuuxuOScBB+gwL9
dNGs9zp++jPlwWrozwJgFxwF6mXSN1FFP7aeNAA3ry+KICmbsnnlV4qqHyQM
jUF4C9yw7AkCs7/V8o23NzyFDBLhb7R7K/PvJMWus8xcvdSE+f3DmPUkHyyw
V2krsJ6jo/WfYWiSloRcJruIkN9wDDEzzn9wZK3rnVO4TGcQTGw6bLVAx882
9u5EtRR+VaDr2nQbk9PyQ4Az3DRVH8TODgn71abmFp4yuzhwJk3oMqJ+69Xm
0SJiGKSW8e3Izyh5ATpYCkypeWX5T66iXVm/IuoIg6emANZP5ipKZRbC74TL
Mqhtkfi6M8xCO97Th2599FyMYkm1iQ2AkZmirLWsoVTm3NvCcdLReaqfljho
hLTcec1ZOf+vR+Bj3atmyx5mOIPWrDMoHITg6fbVYgZdSHW71qJbLuXZwmHT
fK2OR6m2zWm9M3/UtxvmU7DKuMnYklimeXlXI57Bhpm3lAK5v5XiaV3SCduD
KivysC9WpHmBinZHcWrwz9LuJaZUHG1zeY/TQBirQU+zWTBTQWIAZgzVp/ZK
pA8XUUIlq22rqrybNYXiYD6NaryE5pc0bzU7wuCRPO91R8CFWxtGTCFW67U1
cfqFlb1avS/GhYc6MDUE2lIWuNAVWoVWfr4d87In1IdiMjfqOqgRXDvdHpz4
OlF0Hpiw0aeGt0EHPB7eRTFGoeRr5n75hpQ01H4hQ+Pfje/v7/Pk223pmCBC
6biACDS6Qk3u/CCjBDtUxO3wmvF9ouuX7ZiodGg0CysqQ5vRojO/jF9gQFKG
1rdaGznXw7/WT2LovRf5WJNuCIKPMoMUkq+lJjwYlsMLYPgZ3XkCgUwg0s6v
uZCPHke7jswCkK8zeDuZup//YVR+g8batWXVQ2890XSCxuD1aa0ptO4Ivgsu
eBpvuvoJNUx6mWG9MDVo7p0VjT3zqqdIR2SikE92u23IImiNuJPI6O0UrNgt
8ngu1x8Yo6a+vZTG7M8aZcTUoxYxPJ0rdeDoLtQgbDoMkCeqSG1jG3Ea1Tj0
TcnIyz0TxsrIUNDkRc2qyH2fpa6QeErsGkyVY3MhzTw7VfIKrEDqRFCGA96e
Eiuju3Bs7P2FaoU6ByieBIfTryGiwTbwKD1WTXq+eUnhFQEnctEGikKKOpua
SJwosf6Fc+cs6v/CS1lAhTZcUrpx6rulNtor4HerP8kHRK9m7sDRVVmvm2ln
NxgkrcFWIAybHvSDnn8QShnKe6viYR5gnFz0NO/IxWNEQ3knTfdCjnzsDMgX
oBi5YCVCDHs04jIq8EX9h4NOpyF/n/3EYwlawa3sDeniEf3uVXpSa7HP60UL
g7ODtPDn70JB5ivKPf3eu1XrRNI3UsYyEucksFnbSLsouJEXNyn3d++lbfUp
o3pah1uvP3tbbQZTijxgRPRXWoTvGNcj26V6O2pQPOOJpynvZsKY1+fXi61I
7m3voTTp9Tv9QRAxOnKWerPIU7WsLPB1CiM2XTWoNU2mMsYV3xL4BTMNZeyU
m9trbKEVVWxZqqWCdr+O9PTn8Et1KiJMn3cSgnuiswRvKu9/WQYn7fqdYRuK
LwF9SpxPrZVvML5QImrTcTZiVRnbChI1nWt9H20/G08RwO+hi6TstHv/ZR/y
63ejdco+HeAGplhkr36AJW7RBP1R2lrYeSGJQ31f749OnJ9w/KXBdYsnUDje
ibQS4M5ic2TrF0BZa/DxNrpbpRVppBQMztJmbve7/T046NbkeOEpmrPuIKbB
qQDg8dReL5p3Trgi0AAAMwD+XsNOZLE553sZhRZyj3BUMt+EHwCHb9Be3rfe
Vd9bugA+katLv8kgXVyluK/I1cU5R+oUiHD4Ryz61knNKcW0RhUxc1gqoWVz
d3LXpPoJIXFE0bZSj+M/C5JS6Pn09kOSfOV9aMc2nrA8gYAl2Hbji+YJ1D/R
R/RuFX1mrARRSpBF+cPnl55qCflvmGRARJnlLcX8ph4cPzGtu9B+E5eU18Fc
Ahh+z4niH7G6C4yAobKb6EARHD6sOO2OpvJCTkxMtMTPOGI6yQcGTpcLou6N
2FLr7IFWpHp3BAxVMPLuqlKch/PiBnzzuz9cpXacDsOggTeaUZmjTbIh4uae
5kKvSb6ABkjyr4VNjXeXn3IYpIExrf3CAKQVDoSkcNXZjJoEGAdUKAZ2mO3y
zD0FwL20T5Kfa0wETi6X0fnYr6jikFvGIp7FmN2CKsEqWG1CybEYMNmh3Ufj
aVE3YlvQDpOlVmnF2qfp6CqzeFdohTdM1cASLYTQmswRrouBh9oEreduCbYn
q6xLKKLhEJWNc7P9KMidpfXKr8L4uY0JqsEFcSP8FOKt4Cw0v944KrgVTQDB
PRw2FIw55PdWg8TeOwPLw9SusvURcXHXbFK6KH6FpHKzzEXuJCk6/XGTth3F
SUmINwwq3QVSPwPOsHUvNMOFAYBAWJ2w8+/oiaVhkqYZCpSIh6HoKmpdiP4+
/XVLBT8KeI70OIQPhkDwvjOZ0jZLkplg2/xGFOpxsxEgB6pgt53DU76TmJeY
0i2X0WugJnRKR4uie18yA4I0EVrdCUA/u3hA6I7IzFYfEy61mNRKzbkt5GUT
0Xve3kLxJLnQJemW2hU0Qq6woNCVTN2nhp9K07Fu76fqmzzukPl+dmm4RMPK
PYuwSjIXRFb5myi1g1lsMcRB49M1/ZwhaDcfXBhLyfsVhKaf+zQ+aNEf800A
nrgTcRR/Mecv1Rl0Rff+Qb1CNs2AiHQWsCrQDCNBEiQAi+cA6woVVlaVcdXV
J3bmrJaSqrtRgk7n+4NGwa1Puqqjp8whL0OWYW8G5aDRB+csXLQUCtfOEBfg
zGbLkKhlrSupRM/XmPV7vca4FZF/weQQfJKYsDj8xspBbqYxGRUfVR3uZyTt
7J+RPAZXjBLYYe7r/pHq/i3tVF4AwqepjOVEmmw1Bm3ysumHgmwBtiud3owW
kDOXXcJq32QrTe3mLnlWpqhKsCzlJdPj+eslPJ8c8U/TJg36h+Nso0TtWawo
z/n9WXpKBuQ7scmeYol9KKG7NyXNY99awg46PUGnmK6MwnHf3gTpoS1+XzCG
vS1xxrDsLQFnoKKGgKE0uOSfRpeRe4gcYCfb/n+LgDRk+/rbo70I1uMm8BYU
+hQq9wNeYdO5PJ46wuCunoOuvWmpR3zvDdrV0za3g/7WLSSpRJKzlxS+8sRM
R8qQPafYnpPoR/c/QvzwHoq8musJDZP64f06ocPndpY652h06z4+WkHFgK33
uzwwb2mqPDfznfuhpzyhB8cMOk7CzXuuA54vjWtqbRVn6edcQkgrrWcMGpRu
j/fQVVWi5iCh9Ut6gsQGj8rLIrwxTjiNOr2KuPQHgdu5zRCTom2OMbuerQIM
LjzQILO3g6gAaYBzrfLQU4HS0gJrkn2rusZ9gMSJWO1PraFB5ZRDM13kmnIj
mBfp7aHsB8FzJJqVo/5FNHMTNzNO+5gtFWQcTrpmObsM8T2N5OVgf8ux99IE
IYkXc42AVaoQLLoNdZ9R8kZOsaNIStthcbGyyP87/yq1fqlDVz2Hr941RQqQ
5yxq7irhqrS4i12bxlvOLgJFO2kzyfUPdphBzQGHdQCADRgOU1dcIDlETi62
K8WXjX7hMnaUz6oIUpTYoKIdwIOkOiPmvjeLgY+b3+M5dC/1cWoAyd5VZX5e
k8gRWkvVi3uysSNMafpHmFBWxlR9+mT8KAHchKEye62x8qDnalldxsGt6aUB
ysZlKKZB9cpf3wAu/Pwg7a1wpxMFntc1EPzaa+xqolIYfzZU0wKasMEREDef
Bvm8SEe4Iw6GvMZGls0fyTDw7uHYkKmceJwXzCt5EMccLQObPfmw11l6ZxBz
weRZkNxy+z2FTYJFtkeu0F1WbTDBJrb0FmpL+h20TzCpIHKgOC5BfUuA47gJ
wJlAfHcEZugQ8lHe4+jLW9hjc2lu5w+3TGCr+6QVWPKfz44RtST51IL4PQdu
SmrODJ/D/R8QtOaqTLsqpwebnKeNTkPCYYvTc1PcFNibt6WKe1QvRQCLE5NN
7EuL592sOwxqj1FfcVoqUXVU1IxETpCk4TmuI9+blG91rQ/7R7YrsS2bRveQ
ye7lPECC+g/YVVkBUq/AZCG1JQimNfI6m6ndFSbbbTZp7wkMfSVyefy/WrnQ
CUQkVvCWgzgbJ0r1Y+kx1FHFEO8ZwM/tBdE7hmNORLDbdkTTGXvgC2g0lXoJ
e3hBfzdxv9hnKFlJpD3o0NP6JFZL3SWcLLMoagM2aWPHIKkEedsYUzs6l5L8
miWIlsGUrgUpoqDm5jWPOXo+nDpZIxeAzpWviGZr3tFv6RmaSQ6yob0WPwlQ
b5UQeGnj1JCDab6As2Sqz+jsAWuHeodzygWg9nP26sSskqel5ek4h5TzXPq3
xHXacXmENh05Xz/HCMlTxfj2ryHWciZNPlO8vm9bfq8ZVNIRSG9v7k62O/Vc
vqDMMvv9rRORfyq9uWUrIAPmuSZTyohN9OxBLWKCcT7NOt54ubMO6QISICWm
SNF74SaNcTX2cP8O+lXSws8ufkoE0OIjZ3tXAKhSm5r/iZJob/YRhmLvb9le
DRCkfB1lkGVGebtpMy7gCB6sOOclAkOKzEbZ2ertbo+gyf4vVIMcCh8JclBP
2ErX2xOsbMBhBRew1/sdfwXZyNCAyGSIRS3XXDj9dVRg/MMsLRTkndbMdeDR
q/HOU+YoOPkfU/dtKH9yDqfiV0w1MBF9TgPsx/3g+m5q8xlXxI4i3953W44e
4IuuNVfCyNwx2bNjlr3ZZZ5SeQPn/wW4Pc804AhRYnCSJW81mmsc5UmMVNG2
rqembKbTslIuHvRd2Dg/LKqhdeVDoH9J2r2oR9XxBYIFOR8nF7mRRhFeZrd4
bslFw++4cgMCg9r7KNxL8Yis7Y8b5l3fi7X4K2vrKphprFmWGT0pAirBujzM
BXjRJrHnLZAbImlvcllLHDMhyAsdpgkte3R5W5hkiQF0CPGWqzaJZCxqGdcT
hq91DKHwMSOY5FZRq5e9p3bivxOdE1wgrKzM2H3Hvz2O9JNxLcrDDP1ooOcF
ByBIPuZZ80tNhXaIwA2fACM6kpTCCjYqHk0x0S3H/1BSBx1Aa9WW9Z8b97OI
xL7gN4hQDDkfZzT4VqDSoKNJ7IAzKQft5XvP8EcgRooYAv3eLiG0LrcYXSlC
H+caATEKRHdbbEqXv+ngzClXMcqSWZ8/clTpb18wWLX6rsEUzw4MWC34QPH9
HE81jx8B0r8Ci27MpeYIPZ/tryQxpYcyhOKOdbwxL0xrSxHxPnip31dppWwj
HNHPcG+CCeh0PIvAN29B2Ea+RBv26qYZjDbu57Pzn5vLeiGxQ9fM+Hos0nnH
kCwDDpk8ahRZXNAyIxLssAtvikck8Kb6hL94PS/YMVBj0kEaZCksLvxh15+p
Xwd+MjsIJEMSHZsYWN3bXtECI96ykjPYNh9rB8EvsxYvhcrtMDiphf2qCnpA
0tLTqH2y+uLNLKtmVryoPr3Xa3lQQj01P33GW629LByOcRkOjpKhUCB5XVxR
8vo9OVg9nybeEu1zKvC1C1Tb3p4wPw5CLxfZ3Ueef80U4ZkgSsaaS7t67Q74
18n35g63eFGd+NogSgLJPVkWu3wvF8igKvJ0WAfdC7ljadi2IMitJWsK+B/A
NG3PviWwZbz40XcNm2VERcSga07HXuOFUT9Q0dEo6XEBZAbh9zLMzYr//aQJ
wIKNXLVXp2tQIT/pE4BPOumv15hDrIh4m7jgPyw7Oz8yCc1l5Sk+tDTGRnKJ
e+bZ8AMrh6S/2XfyKovkn338k8MgIodAKDMVicVon6TacuP5YClZ4xSXBNga
+UWzbK5vZuyGV8cXgjDAxR21QuqTR8e1KqeZvZhxkdQrPSFwZT4a3Bf3W1tO
VJIUH5VnkiqoEoz2hviC7b4Bz4415V2lKK2Y8HcEtfEl5HnAnCMXOC9a1+O2
nLSxnH55lXGjM0XrcEG498pCWqCkwwN+b4tQg5Qegl074PCnsmZkHuPjPCJo
CBwPvB8ZstOiQ7QHXWb82Nu7tNzX5tiEJ2cd+n+zJeay7tuOXCPFVoEAETas
75Oba1+2VuquLXD69zXzev1QJ1qXZ52S0Dtv/SaShupzjuTwznSKZ/vd6jeU
tiaw+4SFLM7/xX0MOHMSU1TJO6EsT/ZYSQdQPKUVHoU07wSVeVzPpPkE6HpP
TpNVpWstrTUx9Rcwyd64pIg+YsFCp38/b7T3BIkEGkRa4NBkOq4YnG8Qp2B4
QJb0oHlMg8yiqjuJc1z9mihKMiNXbZrVexAPL2rN9f5wcAgSec4H6XJB6F3t
WjgAU2ecC+liawCR4yB5U3Hm1Att8DuSi5GvmmS9QJen0XQB/Hmxt/CPzNV4
JngeaqrNHYI6tqF7BN97rzA6RIxFQhEFf3aTyRPenb0dCBDAjqdrOxLlkm1e
o52IhC4ax6eDGrS+RQ1WxugxtD32RGRyDIuNDtu61x2BBQJ6uUWu7H6T0Tnu
NLZpuy67JeJe0s4L4mxOoA4MprifNPqQKwbAJ6666osufymatOtS6uAlDFzg
14X6nDVmuaVpzfOcD5eeFeqvHZcJxibgkhlJO7h2ieTiGAiz/J3FMKP63SvE
ZTuhKT6b/HlrKwBZX0y6xY7N9rp+5YnpC3ZirGFxlQ4Ae5Uwzw1+pHwKRGb2
iG/m9wcq7dlRTK7syRxXbdGg1b45GL9vdPqjsY4NbyWL6jRGYPaTmag9T/65
VJj0JQpgsS74If/FvsioyuZD02NaaLok6sGyqu8SrAigp/Y6/s4IX17sQKJ+
8hn/FkbGKL5JE5cNTvUt/poDjF4+DnXK1jC695yD49hMKD6Ai5e5ATAudc24
A00171rGH//ojEwo8RSJjREnwubOoh6qNoYyPMqnPYHvo8eTw8ouXNtY0K8w
XsRIVrzo15qqtbvh5tKaxpqLHOx2KyHSCF2w1qjRQE9GbvTXE7LrCtjNBJrb
+OvZCLbfcKRWP5HpWBeOi5LurwUT6miid7V+Xk2j/qEEe///CC7bmVvA8SZx
yekxzJ0dklDih4Qd2Y7JNgXrDq1kU6TDCHYjrthbIJEXNNq83lynvLR0agOm
WNLDs9Ft5FApveD34bdbxoNFEnX3UQmUQYxpfsPMTfd9huw8ORpepayxpY7t
9l3GBNsG3c3qLe22yMVn7IYXD3T083ED2wJj53iYRs6rTUwQ8OHhIoD9lQtW
2SHIHRJ4P1rpwFPIgdkFTPCnnjr7AV585+uFH+m3mRcwnpX+3EDPZ6mi6t4B
aP72VYrXqfFERXukY0PQRd4JZUpharuHcNDt8syf98XvlWNiLAPyRH5KsfDd
H4vNRiJwbGUAUGkwVK7NabSEJl8WcJODuJckj2RKOGAm2SiVcumskg0havGc
eJ7Gl22pyIUMDOHG560lt1wayAfTnnocX4uR5MEjZQzzD9kpbwtUDMmDEcLv
cLXcXTQUJuuEB42S3r1Lrbj5hoLHZvlUCe6mkdZcrgJd322Z3s4hZgFKFVRz
C9rIiREevnD6yFjkU3DmqSh6wHYAityiTEBUsgy3ol5em9ZPVwc2X4plbhuj
cj1K14fbrF2UxaNdefMtKp0s3S9ikRyZqxmKJF5C94i55EwhvPKBdNPmkKaJ
XgbBdVvEv2g5wK7U41r1Vp8KDDROZJKNWQRoOleXZckXf4VndzlhDR/PPNdy
ZfzuPSGlkmwtHvJYdFLhovVhkGLWPxg9o5FMsrn/cc7G8QfKRHEOCIJp72rl
NVwc1+IrUN8//gpgSCfTi03ccdr8ht+MaQTCScjibjFMRlurWJZL1CjC3eCk
3MJHTTobYr6Y/cn2RugQ879Mn+q0h92S9ud0IHGutYL/oeNTSVWaUM0Efr9X
ovf+l8J1BgcJP1H6CKi+f4LzEyUDO37ToiVoMrzFJK1dFD8uTKeqR52M/3OU
Vbde+ZBCyKwrx439xlJzjttPi6qj14SuErIIGUahEZHW7e48zwn4/PE49Yhu
piyYG53rdkUK+t7E8uJAc2Ie0H43bE3lZyH4tB/iHqNIIB8JaMikD/1fdeIf
VD1KTaqVaUtjur+Q9dljEVoRn4oSuYVZiOVLMcWthXyHD+4EvDkvYEKG4Oti
1wx08DaLcKYHev7XC3N5iFY+qUyW0dPCxNSmxrmTVtMXB43KMCJ/esz3X6x/
0QJWJFRiXqtzbPw6qZGOk2NI30rYk3lXzgsGsnXsQrKONeCChJr2CDYamHMP
dm+jSgbgAZ8O3HYfLihMI5onqe6LnqvNLBc6+ofJNm1wVepDQueVng0CzTTM
WGm8p6/gs06VacaNMtnf5mh+wiIyZunEek+AIRTYCqnU3TG6XyrCjdDlHbLS
4isYQLGBD+okapcf4jxY97RArw/jRf0AI1XUFWeL2gBs4QAzmll/vaC87dRv
FGdJMgzFssUZ90ZKOCTR1oMR8mjleDrSL5irmqfpG9R4tG4fnsLCg/M/Yc3e
wJl4DhX8cjcZ7222K1teS+QeQmkue4LBRZHzp4mGe69QI50+jhEdc5JWPKb2
fRenTLaZkHLu0neNz7VtxJPzKWbItWmKEqoyiqP+5LW535JL+Izk7hYHo59H
QNkpeaMW7lbZI2uAyCT3Xj1Dmapgg5MJ8zdcXeqfBMKBY1gGAdwje0W2RyXD
JEPfsqXM/lZ/nuzvygAFTK3TsvzJMT5VIwJ5RkzmD8bYSyD/MY4ndaTriZpV
J6w320Nrf/PRSKOY51DXIHcKxRWy+4qQkkJq++LGhCt94DszKsGTKUxgq6Kt
ZGeM6JCVmxaze+xFANoQjPZ8UbUeK5dy7s+H/pOoF39IdLG7L3wnexB8H3U1
N99T1s6kOqv8RZm/G7F2Q/HENkDhJxgdkOv5bCHpXYVjYSMUTfnPn76IhQIr
CfAXWWx1/5OWxW/e0mvWfD1IrHM8YxTno5PW9ZUE9VuQ3ETCa2w08dH6Lo3D
WSVAYFFzOTYQ9y6I+bQ5ddnOHMUKoLgvOTF/5nSzJOHd2ZhuVtiTJx48JHNI
FBfV2MZB4DQmFbzRhG9HCYxrEBzlVvV889KvlVMT7FhTQIpHm2Op6eIx3T0V
5bFAeOYsxCeSogpVa9i/VsTnNK8LTlNKjga1+wms8Z/esnstL0gYSyEbfGov
gPUaddGX+QG67ogJgeW5K51rxzQdFPqCi1RnHtIIUnN2dTYFVM1KuG9iAp3L
FX7t2uR6k02dLaFnVzgFMGep9q3+40/In789ro7hvyys5VHWgc8qpLk/QAre
pFc1PnC+ItZ9GqVhNWtCvybQxnYYs+kosn+Vnv9dU90asPLOc4K0LSZxckwo
13mj9Kc5d2sjBr4eRX74etkjNaIzbYDpnk1o8ZhUEuxd7OoABnIxcUi16eSK
qTHeRWtjRQfB5j6D/J+lQ0l2h+lFUFE2rUEf6xcATHlc2/B0cbMdV4HemmEt
nCCLVRGcuSWJWkhKnUSLjnrbXeEfq3KQQ2tgPuYqpHdEenRb7K3BqvxjfXCa
6gFyRVzLizOgpxySTvUQLlcpuKRYvfucmmyH21vEPGnWYb7F4oKdmXOQhRla
S86jsV8AGi+Dq46304IFDxa76VfWEJ8nhQkNfhgnPveB6Y579fP5KLW2drxH
PqAy5h8JGSzG+qdf6xMZx7QZr6DvRk+/w7N/R7+jnSINb5RLIFf1r9FNxgrw
YPTaFJUGlInYwN6m3cb7Rfu07Xinbb0bWdkiYVzImiGtpffwONW3IIoV+6O7
6asaJaGRKgSLQIHMyRiFs81yMX1u5Gb8lJh2T6WOLEJWsPrpiC2OGtSIKnkI
3RrX6hh5br14jz+YhtEos7+JimtgGGOsb0BNWz7YmGaZFNUPJxeuKUmHn6+T
yahLrorDbahFAjsV92/DlCdVvNsw78p3b1CXR+4FQgMPntldyMZ4BWpvve9D
bxmqq+q/OWVL+I/MzvauPYgoTmEWNXRGcHXxsQT4frt5fRmjPc6Iy08iYLhY
hQLtL6ZwKcoZCWoKFahitnF87Wk54+yyrUevLCHO8oT8NrOxE+sK4HubmPSj
ZMotpsFVvLOV5tGwUYVarplNo1oRuqd6na9s3lHM9dg8ztqSLKYgTJX7XmrL
4JfhiqpB+iiJeZoNYJyCsNmW4gkynWNykFZK9MPFuPapiMPfArIQ6amZJClD
13tyaBT9RtQ3jWDgE8kyeaE1SLX9Xwi3YK8PSIw/38bJ/F81gtmbnaRfWys6
R6y/BQ0GRvimAvkF2hEaaPdZ0IK9Jz1JaqGjpIQYHaIS08H3LSmOlMcYmgOF
KOPQLe3EDvSSM7uCLOYZ9pLY8alzOkgPeKJXmPb0UFKqawo/9rBR79vrhXDh
BWwg0vVqBAI5tab1XFfmvaYMk4zhru3nxcvCOAl/+JCewo1NjbgJFfE+Z3EN
5nbX4xIpHIh2oK68pBr40MTzApG82PFRo07W0qThUodhBOr2n4hYivrG1FiN
IbVBU54hUgIYf/2ZYWe9HvKWvZ+og1bOebuX71k7h2bVHxyf7NvM+7GfytEn
MNXWMWH1Y81G6RuT3bl/DzKIJDWQw/Dihf2yN58wEzKr7Rhxe+0XfVAa4Hav
BFRKM0UgUNmIwI4MheknDE1Inm1CUE0bK3JKHADcVXL+5VcuJAsrMP/QDj+y
RFTM9p//ZEg0ArTrsu3Q3bH06F9AIVrqeyLiC//FyPu0ucIISSLHh8TGsWhA
MXVfCyZgUpUXbBR5rT8MhyFaBRrQXruA9jUTTGWZvXwd+d/O4EoHsyJywxM0
A6QwrGvwwe6ysalcfFuGoQBYUIi2WCX8Z7tayTuSqMsgdkWNWYQUG3GPLhsu
JKNHLtiyISyDu+bsMxJD6iRXQ/ncu+SiNQPo2fB+w6w035Lkyjk6R8BL+3zT
zXhDDYwx5kvnOSXTZGiqC8IaBjpG4CyowyytZox/b0y+zQ9Ci3m1ACs5BC3J
M1hWWU96ECiK0rkXDGd42NNLV+7bPke0eJD+h3wsEhSbElBx4DcUmtZtB1iZ
Cnw72QNUkUeH/He8ZLYvhtcvfFGmfP5CJ0cJj8j74QPNMrv+e3PvU6/Fd55q
tpF+zXjJNBbKqcDpRT3azmrDtp95xFi3K/Ccp/aFYdpGDh50RzqOg0vioepK
Offu2RNJZr4qjcOjDk+uif2JHXFgnUa2yO+Ng37J2nGoz/Qd7A4EafsvHYB9
weD+TkwY0vhTElgSVYSPLNWzNQjcgxQMMtrYyOWCocrghdSjrLhk2VmJZTKn
k7lYy/sWc9fOKrbPYqyiE1R5TE+T/i3DgKIyyGHj4GXInVKvIPr72bg9oEAm
TZb2dbX9yajvkK67SwUC582lXEKrdFaJbPP0gi+Tizz33sjHRctCqp9LqMLu
kNuJLQHKk3s2uYeCIHYt7i4VnRhXmAq1oaPXlSJTDdTCVELcFR9rGwTk20a1
fTt7JUDxaEjp6Htk1RNcUMa2SfRs3AyMiFyPhzGQDRLp32egjgxTiJjzHZhr
IIoZBfmyURof96eLjiv60HOOKBMpdNBGYhIY70d5Gm/DG/aNOpveqq3iCUBz
2mxdv6mt/xBXId4fW+7TMjzJSJc3VFEjmW23deaRRLMiHYx3LW3fD/oKX47y
uuPIJy6Wg/a7Y9hX8OzD+4WSJBAlSUqeQ8bO9BYkvNT07AFbu+Ib4Gmd72/u
L9wHjS3K+P5yuli8vz7D9wuB0cUF9DxSkVeRTgtqWBkmHvXl4D4nq+/QpZTx
AM4QibwusqLswKGw6aRqHUYNXhHGvpp943hyN6PgFXr6hq1JFM1r7NKa5dxi
yu0e7OnyScUgBCUP0tSBbUalfkxyzMhAKZm3tfDqo2WPepQG8cjbVGQjJSbM
gabHkWnowsUmU0kp9YAiJgpcdbNggiL+dHjdsAm/19box0cymeNC9T1a2vHz
JHtQl06YCW/7FnmcBj/SB0csorMJYmTTR/06zzxvFaBElFSssK60C7r/62Fo
eb/lDVL6zwS1zGm2IDOWYYJN7aq9gx41mV+xgDJBDjA1oWFYirdPrxcIwWzP
G7tmkTSVKgdp5FTuaQg9wcac9EUNYtlTgfOP0SYXwo1QWuJ570JZOgjXvKnE
Ws/xB6hfr9zFrhbVYUTmDU1HW6yVmh0B+heYJScePinS7WeTJyRgrkcHeOr8
uM+27HJG7vX+3V2z02zEYEKRUHB0Q3e+SX6r3CYMprD2Izi7jGJ2syOACYAc
ClRNR7Ons34TbAGMHpyweSYTsuj/ckP8g2qAjrsddCD590TMfC2iDaWQREmP
UYwz5vMEySKozciG5oXHdO7VmILZfyJ9EqQj7r6sjick6Dka/eRF8VluDz0S
+0RW8tGW6OF1Ran8m0nDkYC2KzsbhHP7tqJVVXuhRNbctNV/AqFN7LBX37l/
Uvtvcu/nNKwIXuzBRUJAf9oqUdhg+BxS6TxiF2QHZDPE4x97xTb7HgqUswFC
Gvrt5p4EBoGmsC7CxoWPs89DrXOYx8BQHjGuzzWtTlX4h40G2tqNM+M0Gg2F
o5Bdrns56cg3RRM3d/DmUZUs2GCrecs9gV8CGYD/VJ4idUM+u0/NXU44Hp5o
KdGKG+BRlSXrx+aXfUaKspO8a216oc5Iv0wyycXtQSWqeNTmak4ist7p5vMU
LuUjEQgjhIH5E0oSsJjt+GyjlkYxJBFaQgyztgHlnoFW86Q5nylDTToX1tS0
ArYOiSIAxjOiQWd3XNu3UrfNyZOuXjsK9SPT9eerZIBM/6b3CJWwtyiFOPHU
xL0aQ41/4WCQYknrqbgjYT923BuAATX2wMEhMaO+MAWJqaNUcqfX2WH632KT
+wMGLVIBGX1Q0Hq4iduy63uXJ8zcQjbXKzfgnI1gcHn5XsDlB0aqZX/ze1Ci
Ljtaju7dyYovG/7RAJWhw4+8p665aIncjaLMTkvOBH+wHXEGreaN3nSNVuND
B/yEhwgUkXA+Y0KJSuOgctsXQoNESwHXgqL6DJvgQdulGP6OuBUwzfjCNQ1I
oNbcTPPMMAmkMj/wFRxgiv5+NtESv/r1jsoGu0+6CcPKRnBUW8hrLkywROlQ
hZrJNAAklhwOtecV34SE78Mr5As1b4lI9qZuSHOGT3bBZ9cpdKQkfG6w6iT/
u7nNf3JOlkfCgIaNoNHr+aOAylXagLImhTaMeK31Pt/PoEUdxivlsu3g9zQB
0YM90yyyD0GZ0/wRUO1gZbwgA7mqiu9P9qJRieHslRksDnGHgHSohyxk7Q18
iP1BHbjFTV96vO8YFgEYromVMFkvbK+wzfE/bFC6h6m+ZjT/Ph3Wa8xFKDVc
yvBbJpwi5HbknNs+FQg7MF5BUMe+1Vdhs9fi74aUFDUKI7aCat8Ewh6qFq57
nyE5tWQGcbp7LF5uvZllNtXS9vC+NuWfczwZXhjYcWflumW+y876tszDUs6m
0bUfExaucrGWBwIsmVEPekQtn8clWZilD0+l42FGRQm0EiYFBvAs1ibBZCa1
oV/w0uGgDA/SCenhEmWuYs1PYfJGqSo039O1vnJiZk9mckudK1oiNYbBYBxi
DkXF5D6sPoNFL87Cj9ciAR8grfwJgB7wH2jIVXDHd9NbuWofr5NY48UmYa5i
jmqA7qzWi+3OVty6qFSJcc32aLYOAVNbstLcq8L8x94L7xGSyQJpvaoJ/XTZ
sKMwklaVrl6xFCHsZZW6gdFnILnpbbykmBUArKN+oQmEbg3/Oh3NJvsXf/de
nU2nGY1rvh5ilQAdKUtsvKHcja3/mOZxeNc9VWLuqg2N3Cz6A6TS/n0lr7jl
fGyte5lS44ZjC1769tgb99+zw+rMsiVwBRIouPYELEJBj645tV0msnlwJdXC
UNdMtzkgqDharCe+/NXl7xsfAyPkdBKrlADd4jIQVbw0c0B9EzckfKNGV/FT
IVVbR/DdKAiCkBu3NRvP7xBePHptn6SaJDbJtYcdC0gFNsyFF5jltOGgFGNe
EvtpZnqtt1k9/qyCk6SZQ4216GW5TQDqADfVB4jhtS/dUGQF+N7g3VKw/A6R
D7VGfMRcCOGyGH6JIS6fAZQV5MknjvD95yIKFErD6ITTnvRMKu1oTpnoCXHw
luajW0/o3QprK1mq6hynGuySzTUJLcFsrdo/vwaDawWpQ9is0ykW3n3D1wMK
gqPE96TAQrKMFtg029hwAHmR2f+Wfbu94tATu0ubddgzCbcfjraT6tCoSl9p
MCgdVoEI1CSsDJZV/frfk2nqVNwiP9eH/Dlaa7yhZZ4NNDD63mZYKDghFOKn
lBZENSLqMzDH8i6+PkIYOrsYLEiVCD3qaQgUC6QigHlRPBN0bBriXLPYsa3V
Urxy+SiZ33NaYzRlt8ik3YGPS07qQGLaWe+NKPt6td8qD+xfL7IfLxs4brId
1FmIp1GkMtHD7OPHdGZkD5Z/+fuyOgZaIjoqUqF6g0gqxpqPN73BCSKRZ4RH
kqj+7Gr16ppTscsYKv4T1BAM9OJ54SKavc8BJ7EeE/2iZ+4ChZcXGs5tpFxt
FaA7k3eIT/PhmCQsqlUbrWzC6/k7smx05wONUVGBMujTkglKqj2Pz7nmNG1J
k3aqT7leg/CUvYdzjsZmDumjbxViF5AVNIhfCAIuaYaJuIln6hkwVVMDwRfd
sXi7FpnnoF7JXg/B7YRs9gIB8Z55IFLCOZT1dz07IMfaLnW8XzYeNqe6+4mL
TpSR2lzqLvA/gsLfcfmJ88itiYTZuGJ6nvo7Blppi90PcxyVVxwcRlDc4lRH
CzyaxiU7Ch6E4/PKkt0AdQMQ5ARw0se2s/NrmWhYqMm0GD7yiZ+BGvP3q3iO
4zdRtUewBCqat2oMFVFVc2cl5H48TplTcng6nGOr9Vd90/ZF8yfbGQmc6zvA
Az++inU6/7Knqb2cFbMxKyqfKDL9iE9Zhb32H9oAWrM2LmwHw6w0y87WAZGk
hemzdZOS19HJV3nrDlyT7kSGRgy/xrWV37Giqb7dZroeJZ94MEpSd4BakJBN
9OJ8ts+iGKAIwWy8+P/01hOXNEWgKYyRzTbMj7SwMhbsdY9V4T/wPd0zypwD
EHGvBjMxuKPj1udlW3jv0PtsjyFIKLfg/ljnYBlYRGZOU9InosCEt4YQcKAL
UzIeAg0HDWojgzXfV/vkM3lOHZpfGvDRpTTww2oYXwGQYgAHM7S3Au4IvZZA
dewMrs7W59Plrx2Y4aytmsGJqaWSKzYldtHTeJwsF/LpbUsGl9TC7BQWx/sx
0loI3eL0FoDXRuvsnVo0DoedqMiWpQ3aq3dh+NbnHS/ImSj9AR6N+Ezc08wa
7BeDIJ1ivYw9JyaeiJVslRQvafbqFeAG+lb0BHKY6vRDMdJvkjWu2K2wrUAt
9Wr5KfK5wFKTa+/AYcGc7XHRIREMiEDYm7Jy2XYYfAB6YBBFSem5BCqCpAsS
XRQB0LIffPQxp3nKZ4577UOR7ugAjHZ8Vm33lveh8jLhdfPs8SGXSiLr/9YV
5kKWAbfhs+wzT7MHxCI9EZx1gSN9QBaGCfzXrZkP6YNcIoKEvitOx3TUHUJs
EKPhWwS2IVANECEFDBv3s3181FqdImsuosFe8R5Sk+LNIjTfv0FcWZ8lkxlg
CQBPisDzzoQf3VXj/lyAzGfUTEC9chtGnILv2bPGVN59PAEH4RDxqW2tB9kV
x4IpOQPSPU3g0eD5cq0fgn62iiIJ37UP4dwBrT4NS2FCL/acbKVjLYR08T7G
fuFRT0KDQwCQW3rscE7Aoc4gXB3uRZGIXTeG+YWlGiwO+LblUMYz4JxutcQ6
P4nOXJ8/dqnvtc87GJWqznPsQRHloP7uwa3ojOZFk3g+sFG2qLV08Gm/+aeO
cmgZuzJydr2VjB29lQhJD5ZRRnSihspM2oI2UWMYl8mRAvjdUl9aTL87oSRv
H4Lnq0vHUpLCpGdVgbTe2WAqN9o6SXc99dwVM+3rhBIHVN2M58IAAm9nrDOh
APZ/1KANYr5fZJh66REQOfYfuf3nBk2A1/tWUYqkkl9c1KHS23hQgE/bPR/e
llRMtXJZiXNUA3NoZiLH2YYCvOBsdLuXAGX5E4a3VbfJEG1UtpR9vxzePHTR
6joDGdf4osFw5euEHQpi3as+mXYFNhpyMWrTjanMq9gxHgYf67PzqOXUgAmg
G4wf+jMuAJXcbEG5hwoUZgDGM+QdWOwQfpJ2BMWqD/vb7X7OxAzqyixMcSKv
/fu/6jpHzKGx9g/iJUceQaf3T901yk3tGg/9EC+U6l/ca+wPufVOIYRIHLCN
68L5dG+KpnlUdz882hxAp/VDaS+9YP8FeYnjjv21wuUdgfHrHxVfMY/vfJKv
JOLvsflmNm6bj+VRVxjGytfq8z9IBR4kDCw55Y4jv2uRO5oAypxL9lGowZ9L
Nc0fL8epE/3mFYvcKhlcrFboj9JKIjWFyHV8t4hLX9etsK1nk7IItxVETpVt
gR9wR+Ar5xJP7cP3WRspxWGke6KImy//shuhegJE2kHYbRVIK1oahb6tPEQG
kx3WBlS0LS5MsJiecCCZTEiecJf7r3pzgmKKx91iSTNyw/8bgoExUjblKsdv
xMWkmLBxQ+Y8gidqFew7/fYTih1q2M4w2bgib3SzunhZ8N2ptzrSnTvzKPYI
JcoLB2IC7UsAz1gX0ZuaMAxzjtqI+b+LgqxdtGs2tCX8vgvHXXi+yyPE0L1a
zmNCDx81FrkNrbWRDFcWdnR5gisjhnMsQxOJxPpWIsSmVQW8O3rOHzr5XzVP
g9B9UYM1s68pPAQtdUbpWwAMyVVmiJynfxIRYuuLhIoRlZNLec6m3ccv9aQS
aAcsXe0mDkCWSupu1n8V/8KeqZ21R0PpGgDAazrOxe/xtfyIqDUdTp/KU84Y
h5HToJ4oVOoohQlgHQUYLp2j/jhvZKxi9yXOXrjUVYQLCoEm4ChQjX+IlTcr
lbr4f+ZbRxno2iu4ImJygSYqPrLuX/MyoX7KP7xtqoXU43sxPts+OUpS6UjD
C9x7lyDVmBJkfbndb5UJb4JC/Lv6lIeJMGOQiabJqHW32zqL25QWM7lsI9Ri
g45t0qhuZvOXOVsGlm4X3R8NyiK5idIxXRNg6ecZVudPXotl05uEbA8dIdEY
XK6BOJzz42JZvVJhjSF4dbuz5ieHd9bAXCHB0xYuY5I0rmJ0FzLLY2o3WEqc
MXxP1y5vZWSkINi7lynOjW+yPDSfH87K6x/LQKCCOD1u31gK0ZEXNtLHeZxh
EF4NCsy3QtMkCqIudjAzwMCVDzgoqYBEN015EbRkEN2/dRl+MgCY8dnx5+JI
yLwhvNfF5ja6tLyHir7sNJrLrt4fwRiIJIP/rBEkysxxcMRQCYaeRGNFitjH
ItJQ3GxXrZMTTl44SGUp12AzUvF+1JTBRqr42d3zNHjaoQ/RC/c281wGxef8
/aZTRPyL45q91gz619yC5I4MbGAxf55SnFIjqznNEMTrMpiFbrdonC13Ak2Q
qZLMHSTHCenWq52Z9MNDTcITki4NHiYPWcp4EgeAHpNX3WpG4GaN+GEZLe6x
8JGMt/lSprs1IRXQMUeOPdehOdqJm6gPWdIbGJ8gQ/fLofn0uATGUQgYyR/D
HcQkuGTCC6CW9UnRiRans0w8YsK9DdtCwm6xZzEGnzJF4wSwdKD9c7CBj1Kn
wia5BZB4Ilzsycou37lvASLQCVPAZn8rqNUIASX3KgR3iqf0qn4o+bGMrloI
51D2BEL0C6WEQrh4rAhCRthmwAWwsbikDtFCVnv1YQLYjhlYpsajUctJ+Zdv
NjwFEj+y1OG3+yEujZ2KpDaJECLSpj5BDV7XylE2kyUTc8O2Dh3DT/fdAxvm
hdUzoPhFfOBXD/Ioq0V9HHIXySag6k1TH/iR6PGYq0k2C45W90xeYxX4GQlx
DZP3f3afL8wypTUug+79sqANIThaHGbLH7geNwOU9JQgWUCOQH9xF/Bntbxf
rxsCAksX0rgUyoF2yfYtsVJx5R3t2v8F9tSd0saUsr4oU04HUfMW+AMYeW2b
YzNtt72lxsgEQT55taa1TpeKhMPhZI+p2Ky+dyuetIMv6zvv2E+XszeC0BQ3
+DiFiad7ZO91fea+KFB0RWVZTL6t5h1iK+fcEkDomcmGinrovt2cLWe8vp3u
+z52hjyTrEOfa4DuTYbHFTOL5Fb8wnjmd+ltFH4x5E5mLcw6DRyrQpkyA4LV
ZqZ3PkCvl34WRZmfBIQeOsGHuIZ9QH/vb9Pl6q35MHj8y9lBOZuuecBWXk/9
V/5YCBxkVKTIgPgDoCivClqsnWK4qwe/YdL7u3qg+ia+wK4ruB9obBJWLOfX
iRuOsCAg6N4rM8BWit0dpSd+X4KeY8ySA4R7cHnq4+oInlIq/yioJyJimj86
uJrdnkJIb4+P6wbFpcM84mFXn2/DaR3UJ3R0OUzSRk/noyasxw/8N2iKpOcJ
K5BuuiEbZW70HV14QEjqE6ee4e2Wcdgpxvx2L62GnQ/4i46JaagO/CSn4c8N
RROPpR0wxDah9V9p9OaZ1UeYSOZ5njhLyT86MtY7T1DcaA8XxAF1i1T1MqvF
tAoyXClQJ+sCOeT9h2EKhG7Q3OMXqR/R//c2DT7J7z/NyMfcymo8ojypfQr8
HrcTWltScDuEtV4y2E01HTl9zMgbT6LuSudHikoc6SVTp/HeSAiUIlmHdG3F
zuPdAvlLaGXxp5ul570ari7bsDbSle5kafkSI9FatMzadSE88H3EKojs5zQC
SvRYr02jT/szS2Yr81Cu38ydPqEmVzwqcUNZdqOgqC/WZa96/Ro7qiCg+nj8
SgC0ETbbwnEB0st077qgV3aRGXcViF5kSuUYj8LEZXXzoB5RGdEsjccY7T2c
xdYUWEGhOQvANY0RmuCSBTz8ZQM4MdLWOaptJKYxWCZECtv8Py8X35jEvQ7Q
2LrTtMCyO0sg5WEhr7jtodLo+FLozqfpTv7+eaBDaWndoeoDXITJ+MqLATWF
vZnGTEvYzbGW4+Yov5lxhLJ+nYvg6mL+fW4nhhLVIRtlTuToLnM23gKKhxvd
hQTL31+NaDt4EHIGApvEgP2VTRBDFg3tfFUWWG61I40fPDd1YpqYkhnL0HrG
xS23B6dmCrBRa0nE8vLT7vaX3X1vB6IXZyU1RsAfD4x67Aw6ZJHUAk1XbBGa
Jj1OPQmYky9uJPNEH3hbXx01vo7ATRFGbG+duoNf0l4ZRa7pbp8qL8LSufgW
pwEJvcLJLBpIanzHU/oIIToyw1sknj45rNvOgMktB+1jS9D9E6GePWsKwdCA
/9hUsEA/7YWa09+cWf/abcVXzrxQY2YZSEH4kilSk5JswbiSZ11/0SnhPRbg
JwbjQSftQ5KcwJxCzv9E7/JEDR59Nfx/oHplF9x4rO/pRqF0d30obChYy0jv
hMU/1cd081j4uM7idTOT5SSlkLhVUziOcto9KtMU5DyD4CoibEKChJZ/212M
zGRw17tlA3XraNTGtEcEviKRh6SxRG8of3/LRDLysoAHmy3xrc14/sIVrZ3k
RzSJoZLctXXt7smnktvN76JgV6lAm9neFU+bbHOAb/vf0QSu9CLnyhuAFxwY
Jx4h4u+2P8MyZCGZwwLDa6C63gAmb8lnLWwAQZJcMH5JAWhC4xRx54G3j7Rx
zgJkuC0yUmJ5TB1qkH07jOM/Wew5B0BiXrlBqnDd8K2KqtVWRNo9fTPeZXR3
ZfbTxff560cwnSe8fQOYCaLhzn/zW4WW8QTSH4/8dzpr2L12EWTO01igJtUR
3EIdxdGbd+bs05OdbkQguwXtzPguAC9qUdbGgY3IZx7ySDFc0IQXCKXC8z09
9XXKOX9yZNBNHlicsoKAVK0PYVAGJLtFhWppAIWFawF5wNq1XEBNy+fF14qr
kZyK8VkXxlyoazLVF8VpCSc4pEKUO5M/ECDKHmCE25t7h1yDKkBhzRlYYBM7
qDXHLVoR72+RIEKPGcdyjxkpIMCdbGP1MjuEIhmb2TFaJsIj0SFhb9AQzNTt
t8OXUUQRZdwntSFF3ta3gVFSmDYkXx3nGWv5pUrj2YHLonNzSs5cLsMHVRS/
2UCym9OGWEMczV+H3efO8fjdgbO6TcME7Wif1LqCPVlXmP0HGuw+kQzr8NUf
i6D+OUAwWFNG4rmCLW/CTJ+m4PoNcWcri1s3WooFDIrST6jkuVYKTvoBeDnB
pEX0C9+ibbhJiLJqZNJQufWyg2cPrg7adFhY8k64N+TufoaqmAh+GtpovRPH
zAYVTPdiIrP9QYA3Jm9WBAsD/YZzBeb5GTQqON/RN42WaNb/71fWVZ5t+gIU
aO8T1doMn/OUXDxGFaKL8bEaZSDZua5DMdP6+sLdvQl9y1Abbp4gyJ3Aggb+
OOHUWsLx7mCUhQApl0mTQ6QUBw22p+H4tV8fj7yZFT6meGVL+6i3+wl1Pqau
/VQUwnKX9QabfIm56rdXBkz7WHvb8YhOjyyHOsHnNrXscJDiJYNRYcpB24hO
jYkLLV3caI2mh/gzZfZCcOFj7fRergJtvFSjaCKp0eP6D6QSD1C7ZubueG9C
/BeoZbbwjOcivCIDwSxF9G4OogGipVWMn3IGihIUEWoGmQ3jpIlnljd5Xu4L
So9Kxwj6OfULQB3UrS90XDonD589GmqOuqBR+KPgp5l62HVDcd33bJJ+utBU
DrbiEu14e3k/nScLIfCMD6XIl2F5tOhAAJ0NQFApUtPuZabSmB6iDq2JzSlq
CuFJX9UY15QqcqOAiD9dIDGmBKwx+tr4u7toCKQ5jRtL6FL0eWZ+h7m655RK
Ep7sGoCud5QAgzwxvenRmrjpM80FljmNMmsvvkUPQLa5sWHf6mPjmXdbJsD2
p4oatSKeYUPxsN1qKcgWVAK+at2XdvnfQbiYYGSygLeH0a8lGv/Xe31WMDea
b52tdphpNVuN9ocwxCy+LNTkyUIQbGO8FNiKcHJWuYgKi22zwBlFhHaCUEuu
SmmTWB04h84o9bXSk367tMlafHEfutu1KHh4L9hsDixyMHpu42UzXsN6ksoK
xIzGMwmzC4FXnrv/D5CbnA3WAtl8ardNA6AkGkrmcYMtSZ7fuum1+BIFDmuE
jMWsBFYpehJ8FuZAgrRkDnF7RdXBxew67HmpCUB9Pazgp8ZI6kWeq31An9nZ
QgA+958LC6Cj2dnaZ8Lm6aXqz0Wh7x2s+t5VJ9KoXNoeW2Vwx4fBfK6Rw4U1
/VUKmqPG3x/ObJeFA9RBuXg6yFPViigsZZXgNpDnE+0I2cKpO/C0+IwFjSFe
mPyof3Ov/mqrE5u2HqdPVCXLRbWpIsLNsvqub3QyyUcE6Zn10uhgBgK399/8
CTdM87R06RO+d1aloOkEE2xu2Co73QTs0p4aHfPX1OnwWqFvcC1zgOxB3PbN
CI+PZ6xgEstMA5issnPejZgYjLjKh+6wgmS1vKXrCswYU9DhHXA6hmogUmPZ
IlfHGZ+E2/K8aG4K8Dyx3dzcMLZyH1nSWrOyLWLAv3PTQyzRvpUVsQ5SH491
vUoNrT5fle60BOhykXTWteF5GUcTx84C/EwXZpkrR7vZwEUmoEnGFsRpdXjr
4HYThExPzOp580bS1/GiLdMZanEQx2ZGQKZIqV9KXyHdK553RzOiIBFHN1ra
qZFdS1BEaQEj6lWasdhrB2YyZD6VySi/EPE6YhAdyMMOuK31X4Iy5nvupwRP
ogebHNKxZ1qy931EGOfecJjLAjhSuH+qa2O8bu53RzL2tylL9WqNHV214Kfp
/LHhuIkTwaKbNc1y+t08SQUB6BWIzr2punuejYC+Da4dVSR63KKJMac4ytIr
kKbZmGQjBx2ZvzPqPs9RTgGJX+CKENVHw5az/eAWnJoqJnRF7UXpIBsNf2pN
W3N18QHXCQJz0etfDoOcc6it/4VU1ke5ZxdE+q+BdaKX4X2tpgcXa+4k9ydP
gnkW3bZ04zTGa8Et1RYAuDf1VTXo1CUkO8FFlfaC4T/VyfSqU5H97es50zJp
KoVe9VfW+XYzPauOHHKBfK50ypTCQntjfs6vzXp8nBOCu0a948ssAwvcyUbF
F/HU9VwZITp5q+YC9jg9raEhIU8e5eKveFCWO7XYEu5bArbnwTAw0WW/I8Rh
mV6njC4reqjuizHKcfgfIGD5rLI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0whsQJT1ifPf5hLf8g46sL245gLYTLoHTb9aCBMfXQAUecIoWs1msS/bzpnEfFOFmxWSt9u8jdBZ7X17bjhEtREhkeMISGw+GWp2XjC9D/dFQdVAT1eOTouIxERbB2VY+LkxqunEOWCuV52LypvoyfvbK6cNI04izFkggs9/hKwl53TePZU9quSgoy9J/5youZ3HolgLCsws2a8ka2ucYWFJWwqy62Vlz6ZHa0i8gM5KvITD/epRvAnKC1Rd+AlCWwdPaEWo9GNSPmBA0AMt2apMAVwrci9imAvBZQv/2HZ3wHoE5etYts3CF88aWaDFKo9jH8RfjXF0C19b4E6dYutHbQLZnb90k+Kv8QpvaoXHds4QEake7gmmnPYXWv2+kPrB+0o0gu6KPlbQMubjQqJr1+rBRDWXCLoHCB9jM4oFmkCjveQhzzT8zsi4yw+L/M0RrANPaAFOUnfJFa/EllmszjhtJ2W+8yl0lS5XDVEZyLqhFAPZujQmLvCSC2iU5ys/+GHJQWxHm5l+NWsRMjft5jgiW3c9p1zRQVwzVhFI3p9uClpY0uSvR4NVXnf0pb8UUsvUgJB6SHTJOwzBzCP8U6dBXU4UxetwRUWcFZlL9MVIX1i6utpvTA3Y1zJAUwHKsg271pnYm8W57zQ+yLwpIVJmvso/mAZy40T5WbvjEI7HJ6hEB1VPH0AMzn31t2Q+fnY1nYiwha8ZBVLmrHDJwyb9dZiLKVzJe+DAsC/BPjfSfZwe71bv7YTFFrvjgKXKZmiO+Q/c3sgsggD165OV"
`endif