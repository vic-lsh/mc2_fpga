// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W7cD8DqzKRMTmW/VUzx7pS1dnv7KH/YOpvyfy9M5Da/qjd8IsQl54cqA7b/p
rOFpeoq1P91aGIXGkD6R8N/kCQQVzbF4Of6wUGRDaAgYvkilCbtwPjHNQe7M
meR3cvU7Yb0xBwQZQ56dhx/9myRJ16guWSMkxj7U6PcyFt7nPYRIn1Guvpgh
6XT5vQAlAp2bnosqq0REitEUfbrLW3nch5v5+h/IHbEYk0uy92rMs2oCnU/8
0OEU2WTy8sXqasT/Nd7tMylWjK1JVw2Yl3KrGPd2zDIld9WTqOZGztJUEIlC
16FnVmpT7aKGYSurN0A5gEenCAsSqy8nP/PYAJ/3Iw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LxdntBN3H9W8fT2L9pmxgTqRJ7PAFBcETmmV5p4M54XubyD2Wb7HRVlpVj4u
ZyETLlsFrFUkpLsTtUdKfI6+ePkir9qiLYvfHRGr5UxYnt9VEiRSjdxuGNKo
5162DVAJJH/KbbYeZy4hWeQdf/+z5vF1KdCZQgtAyY4tfw7VQsJ1QFZk6UNU
2dL27jjrMxJWfc1nMJ5YABPwuL3tv4Wu6zhng/bjP3fFkcZKX++pmiXsYE1H
JR5ZZSMcpsEl8suSDoMZZ8wNBQ2mQy07vyc3U/0OuDJdQAuEZByl2lK8c3i2
7zZkH7h1VhsxYh0qk/UN/NoQ0eziXyF8HTkiuhINyw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
r65nF76vC5+9lA7TbKjJu4u+Yx/S6qdD+uOSkHYoqDqlZii4Boy4cAgAY9+k
hIgULPap63mDS5gjU9HqWIUoe/gtjtvkuGaBLRTTiG/tr+YcaQmjDKu4uqof
b47VdgxwKY7VflP7AajlIGzAPx82EHL61jp4qCUzlaBk2oRb80Ek8jC2HbPh
Njab8fib3LaoP8XQ+3krBBKsS17CPrtzUz/7EJx27rQjlDzK9c5k4ZZzeAKU
HUBgBmCy7BxdkXY94Tkp2BNtY1MX8Jwnq9uN1w+meITEloMLmB6hv+HEigAX
uVtkbJSV21ilpKQGgPMZKN67TpES8H0rALYH2pwr/w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LSglp1UtkDoHt0zNbpnRNGHpeYDkVYjV00dvdb1S3R0OdXrE/SFTV4hV9bwz
EzkRTjnAqKbls5KH74qF37MhdhKkshUS84uNIUmM1aoVbkehdAmDbJ5mFcKh
Zx9a8wLA/fm0rpWBTogKDWSSopTUBqAGDLVSFjlrwYbePciv5VRxNfcl7KCW
EY56ptb6qQHpWFzhh3LmLdtYHabGWW5TUO8XYokvssUkA+uybpve5mRsT853
baMNoE1oAeh7EWiWhB5GAzGVoskTHNXeO46CkxFQRNmFcRjphErGdPpeT0ty
Ha6D7Ca5zxjLeYJhuKsQCGOPbbq5bHdD3l4ck+lWmA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tXXVTG5oKufOHpioeb/C2dDap71Pu7grsNs4PGhGtJsGSuIrmnVsqVlh7ECC
BFwo4bgRdIIVF4sZkVZHTT16ZR+dqNrGnJ2Ejsb8l80dQs04lMCM6oenwkWy
PlHs0RaZrKD/mr7yUC5W7cNzwbx9l4NqmTclOgEWZWiw0mc8Q28=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WUgFIsRmM16X/m6Eq+EIEuFYKrkE6HORZ77bNhFhupPCbSk6H5Jw00ghLj05
xfIAIqen2l0JEz1DqdzPu/9VXs6DKKW8HPgDYL/gy4U/XXBkKA0nL0GwXVqL
Owg1PC55n54dIUdNO81zqKIVlUS4hU3rBufDNGg15hOmPI98aREN9ZoHzmvW
HlvDYBJtC16I/a1Ts+rnUvwoINbc8j3gQ07nKtLkoYJpo3WkfEr9pKwDHKZh
1RPQqUV8xfUOqq89ZmTih4J71bJwjrt1zf6eTOR4+032tclSjUjOPJkVD1Al
9yszQ8Ie3t+/lt/mH5j+xgOtCimXhLbIoBrIGKVCx5VqoavqBkG8wLTd6zpF
AAZFX8jLNoy3w/0tAV4yYLP4+8kMB4uaMDOhalaMhAAjZVxilMNJhSAuBGKb
1YSJ67WdvBFbH7p1D5Ovyo11qGevNSAgRnjLHyHMjK+Noh6GZRoVzw28kJyp
Bovwni09ov6FTpY7QJqdASBBP8uiDHes


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VcM7izWvyq/RriLEa2LNP995qqZC898mnBWGZ9JetOokb+Mo9M/+ircWUZ4n
YFP6FMP4HC2hiRuDZyt/pwcXxX+8JMJ1THdN4gM59wy/XdlfdBB+lvtjvs3O
7zQQQ5ggfFWC/B6v+rgl4y0i/jRWqqjrli03OCv52kPpjadjCIA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EvtHNt+/pH4q5h7djvWOk2trKoIgPLjLskMrfoWAe1pcyEwb29ljDLbJu/0f
zsrUGKZ79hgVCSts9WAz4OHk4Lh+RA8u5CKD8FTudDlWMzDQi6Fy1DUpyHtZ
WMopV+Z/FnPXJqXT10g7o+XRJeG3J/1mbxz+tiDJ+t1eZ0KWphc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14960)
`pragma protect data_block
84ul/lx/GTJI55nZCXVjmrZgIN2AvCsFTwLc9RILYpoEvfZ62wcctT3jsgti
K24rgoj0gQyr5UtRAbmmvldppMoOGG6ThnOkKFgIH2OgC2ERmq3F1kmQORAj
RowCZ++5c7sjtHZdG3kaG4NkWX1IlhqHUdGBUbvUnZChiezF+vfnk/xfdbyh
F/yxrK/q4TCsrAxE/IcDlSkIkN1uF2iMlGEygKUpHrslDlNINGEpBSL8yIGX
hDJDpogHsu8MIsAgfMH4zEdZWu1VnOpMin0wyUdDT5xQ0VxltJR5tVkIM1Ay
5sPANKWLzBu9U63fyLYKEtrDyjKuR+TKJCGAVHN0beJ4dd8QB8iqmHMjqGIK
EjCv/dNAeuIM50v3gXTvuJNtFIOjIuiI/SV8nSIWwTZDUPnlEI8l7As8KWJS
ioZOG9iGjfUMKQnPFwDEXAO3II6YHxXyX4KnoCZD3CfUKhwp0VhMvGuvZSR5
6oYJdgfqt/o8AT03A6KrvBHqrgin3lnv01Wdt6smjrCbfQ4MU4R0wh3h43BC
TL5v28LSrVJJbyJe093J9b4PGD7QXZb0HXXJXm/o4xGFHTCjgm9TO1qQuvYy
JY7EPcy7Q797WrHRva8NW1UqKbbaHLaKY6kDjzhnP+E+iHCrtoT6itQeGN8T
lznyR4wwZ5ZHPlheyRnJXQjxFTZKSbojE2H3uid58hVbO8G6ci2swPq8VIgR
JMdwnsNANo6pY8NTKaEAx8hDIPV/3VK4Yh7EMbUZfr89LRh6VHL7d07frMnp
IOSk6SglXdPnXQEk0LMMci3+3foeHLzOVJBvPHiby1vUcBZtluaKYb55AnqE
eDdLa+7YG91YMs6iZkf0dspjKRLva1vyeuXdbVYEOr6zOUL+CdK4xeWGWWcO
jsuxoMHhvFdQOdu/PNls8jDaFq+/AKvqTGgu1O/YluaZaN7c4l6l0v2FNgRh
fd3Dsmx2jAF5TlFo8EwZUiMGQSTplhiRCZeN448AXxE4dBqF7snfQVtkj0aE
j1J1dTNoDTxTwGgcJL/jihj0Wzn0PeiRjB3yMiGeREg7/lvHkd3vc6UT34VF
YxW56rdQH0Qo/grnfzZQk8gmmdW9ipq8j/B7Rg2/8ioC+lvvoJ8s4L3i4nFf
HTSlP5K6iUNqvk1ySefZm6vOpEeLyCGT5dNaaSC3U1849rr7z66taZ7TMniJ
2BGEw6ExlzieSaBULh2xZd4uptFLNQtsT4rFqSspam+zELlERB3xzuKoNOdt
86jMxSlMcRlPQ33EpHdJ/+C9lnt5rdScDciyLFGoiJPvDmxRhr8a3rs46Au8
ErbemFeawmWG3qGYgGGa5pxXz5fLLQq6rIC104DadjDRyaHx6TANEGMvQTCZ
rfvGdhdnhZ/j4nWChtZ5DnyRWuNgkQ0vIQ1DoE2CbmGoT2eQRDInjz1cvOC0
nt7eXjEbG9uI0AEc2U8F7JyGz+L8UHLOnQuxyswXo4ZKCkOMhAIFzgS8wcIx
uBhRufartA8fdBpFXX9R2weJUrW9wj4qqZInH7t6iFBccVRPyYcq5LOb7Z49
tyNZ3vYMeiaNH70fY7RxVieLbWAW0wFxH4JTQCqC7VOalMrg/ryCjhOyphWP
vBjYou+fHit/HqgEBXvwDtKrPTnw/sEOiSpTqDZJoYTgIurf116lMhW5ZsjW
5597Wzisi7bJqtpqtZebm6dZsY5XzOhYmOyAtMu+LQS9VRjfgne3x6Quq0K5
uuBQtIMtEGO2AfC6tW8Se+lvsH2qgZGJDWN4opaA3I19plpZfC8KKyJBRBER
MvfEy3FunEm7IxMQyr1t6i9lJjSFEVOGJzD4lJcVmIlQ9zBoiKYhMG/K4jk9
aCrb83B4NFf3G2jd9Pxfd4J4vmQvBsIx5RcLIb77pkuSSviQzdGCJnW9e4F9
6xSqqJdyX0aTqBJD639aOuksyCQuL53JOlO1+M4MOigvEIeLljqo8bELJpTe
bm96olbC2nbuN0HbCD8EdNVsT7yE+S0FoXLCYeSl1dEAA0WxQr7T2WuxU3tn
yAVTQ2SiHDRjxnNOTR5oj+Yo5X0vZuQokgaOxM/nrPn5mPbcpleR7OE4vRoN
buUy9Otkc1RkqaJUu+yIJNQMizRuBmU1i8oMfg+TMNgW1PmHdBY5Wgojz3mj
GICFgdLKUYKm9VSkJ8bLgx9ASd2HGv/ZFkzRzOHNz/5Rgh2C55CVcFyPvb6+
R3yUTay3F8etvYIddiIPRAE287zO8gHa85GkuZNOqNRZbaX7T8VozwDuOyzb
CytG81GHd9xerTGO8p5uWDOQ1pEh/Or3FLRf92urYvNC0K3M9QO9fm65Sqz2
4eYIuiOjJkzHjuyVf2wPYwutM7XVN+uS/xfT28tKlCDuVYcvkhY+NFqwY31J
mUmkYISXhl59s6IaA7c4IfvxQj8bfva1bAIrxSgsl8fsNuiosRa2PGVppRtV
fkyDMFLc6tzR5Ur19cg3RwmbyWmh6w6cGQ/vNOSfQ9hdlzrP1QOpwjzqVsPA
wVmQb4DB0NWp/kWpwonxFs0sHvjHSomO3deBfo4V76ZL3gmFjvsJWJJgSPAf
30V93rl/el3XhvsMGX2tuxg1ROBgbYUNaHFXhmD6GPXa9d2e/O3gR64Y2kVB
+8WWft6dOvDxVW2oltekbvmIlHl4g+47dOhhi8cDGIWiP0JdeNQxY2Y8YkmV
ONhL+/7RDyP50r5tmStXECwyge/Atau5SgI6e5mIOqXz63r+Sbm2I5B/c3TY
zuGRUGaVcpmTVRIxMH0LRHD2GymW/96kWzoGrpfpzE9IdMu5fkcNy3mDUtKI
VxJZ7KOqBipAaZ4d4qsLtkRqCJwkA6E7EQwrwA5ubWkKI0irAfslMjFfmbIk
hcSR4Ga4fJ0cgbktUFROPrd+qIgNInHQqqxaMVY8u6eFAt2Ap63kYta0OVyu
EVmMUh+aNdg0khJ92U7Y8SdLfqPb45ui7anvYDpBhVQG5yaeHJdwZUFyeraT
zlyZkFoWopYi7C/JhZN07nCP3lRIZt+gRkgyMmn4hmOdyHS1wMsFL3FTNdJf
3vyTLceWDQgCiJlSFceI+p9dbFZUevJDEdr9QojiX4jXUQ4UDZvrpjB+4NxQ
CXzKd1l00ZNaieRjLIHfkK4UyLMJTWW16mGSuxK3JFWMLWNnBmeLu7N7VP9a
W8/EIP6AcYCfQZP93nIkXhbgByHGThrlcbg6PqB894S0ZUvLlkvrTeB2baGU
HK1mrBqk5aMyymcdv+Fn3xlMBUhVmnAF/h1cl5btXQMSFMRJuydz6jLuUD0a
LtqDry7rZ6uz7aofV3Vc1ZYkHCwzSUU0zL2yHS7HtUdygDmRnkMSpUpTrmQ2
MuQllUoE9u15SQHEY2fji/D4QIaFNAvkus5FhvS0cVuKglndL6Pyn4zb57OX
P9zYs2eVN9bnxISH0TAey7wLFPEbHDhTi4TZdZAp8GjULJQZdXhS3Cq/OBj3
Hox1POwexZENW5hnLjqrYaWBFYKzUYfKlzp+7eToS/ucAWlWdcB+07aBt6iw
vsBpyJAF7XDXJcO0frwaUU2pCsCX8K3iZXUzOqJFGSkwRclpPzcyMv6VRDi1
qhVc9lgr6/GtOVZt8uWj7cqPgJule9Fg2/TN0p0Esi/qZmm3ay+CsczWOXRM
/3LXYrq6BOds/VCDfkHcpFL+AQZ0z97hK711HGQtRdUbCSuzkRWSFD9hW+vg
0J5qaxJjnlJts6nfHa5k69j34t+aIZLDaRN/St35x++g775tiGAzAem6i2aY
CyJKmVy2C6gaj2uFbhpAFT1tPKWakEF7ytoDYEFHdrClwjuOUdlF79ImJwUg
8t06y0cL+A85cohqVsGy2LDMWpi1nSdrrQn6v45yfEv2Ng5iWqyaESeO/38a
FMu0mQp0ynMnbkeR5MrN5Pb2/a25SKrLYt5+OyCGE1ieAX4TsluNQ8vhnFCb
VbAyfrStSUBEwoK/1XuYuRu3weBsJMARR1Myg1oKFQYn05q4qlpXVTxHLcNU
zFUOK6/zUD4fOX12/cjYAQjgsI6mCeqmYWlmC0TopIC9+tM+l+3WFE2loXkV
I2quvpjUMLd8rdCrHkigarDdlNck8hpGTCR4/0rYK28Qd6hhv8lBpuU7Kw8n
sOTAWPaa/yCzXB1YDGBQlV9lCeEZUECWEmVqEvOgRTIg8bFNovRA06nASdXk
RIz3hKytzbxtcNrwJuCjTRgY9xB4zmB4mbQfs10dDo6U6/+j+cuLesz7INvk
iUtEIkTGFTRB1rn0K2KPnTwpMjMTLLTSxWBvB10mIKLnrvRIx0oivvDpO6av
Pp8QWidjfEL9n+oLrjvnsQLgd5qRVkEe/LA9HMIjn1ckkCjNjkdyo1Uw7G0Y
CLbFuS7BIDH9MusE4A4ZmB5855g43FZcoCMpiskG0JNfaF1E81XTLVv+AbpP
/NnVuzWI1nLloWr21qJVVazCflnPB1MQJZECMkTu1HR8U46LO9BC7hjBkSjg
qQRVKtssqHkyWNirHXfgOdFZF7GsQcQNnekFofqgHdv9Qd6g7CsATitP7YA2
HXkGfxugdWkxWKDgHDkFj1XwX2DAQVpdA9Qz3UD52o37tFsMe1+Tmb41M2DU
bPjc7mN0P0gZExvL/VhRISABNibAEhuN/nYOZyNdze3Z095Xncqh8Y1RR5HI
ucZOlgvI3ICvUUcNjx8VyCTJGlKtvephSnLO4aGLozadEDOobFaxwjBH6ymD
bAbVBK/iZ7OPAQlPXxDRUlQKNF/RwHHZVzAXBYO1EAgz+KDdICxs5fM482k5
+uiDIGTK7TgRkbE1wuClPwJbWAxJLISwRTRC0/bo4H1jzpK6cOevVlU0qhJc
BINRjSGH46ycluegfSsCAj1mvfVmBn4y8SdE5++iCWnzFLpWSsifesf8a6ec
9MBssAbLdERPTTz9w166CVIfpY22eGgjDWnbmpL89T4iqCpK9q0WAxDskJR1
6qGooW9tnNWk4ipNoMWi2fQzDWzZRvoB/08VXZsfOrAxSA2vR6VHDTzkK+iw
LvPoA6nIGRszu6ja1RsgO8i99dy1LpL2kLmUz9Y5UgYzpuZcvTULPpoz3Rid
oagQklBAGbVUJQpdnMvnVLvQc5LbHrFWzKHsusBtAVc8H2vobZd5JSKkZJ5H
0PYiq/KC3mRSvYiSpBXIUwQ+KNVOstspAGEhod4Go4o9jbTLqAftlyYTgao7
VsBVGgR3sf26HgQwbhylcfvV3Lc29ISNNMoDSATDatKO31M5rL+OOQ1S7xuv
IPMuWTp9iZUSNg/4coGHvdwfI812s50kHOReHC3w9J2h10kEPAFqpG5BmhU8
qVVDbJmg6gC/6zLzY8QbOtUED+i68MhTKyec3WkbqKNRTUNK/Y34DcP+7Xts
R9x/+E8lJEcxwTjkaQ/u8oqoO5SP0SvW+MMQYJTuci7OLaP+jIxHZSBA6Rik
kB+ouH1ExIeL1m+q4ME3siGMqZtx7rX/2eabWXvdj1OuzJpLD9SBgAFLQCMk
PlWoqy1RlGEQJ1UCvxcsn6MfwcwX1coR7owCYGem2x5NWpjXkTPvZDH+QK7l
jvkOAbC3GVTCDtP9kMo9vZVaMtLA8FThngOVQe+KF+fS385gj9I8taG3Cnl5
Gh/daQ45efU6vDZfR9KlPkwvQC1Hht9vRDI8ZHlY8SwZJ01289W6L3hAPVDZ
RIBRzJt16kWo6umVZCYm2Ojm69b042Fn/1RwWFxisR9v660fLFjLRW/jPAcv
5CGXU12VLWTNg0z00/usGXaIcJJqSFIWQwR1ExlObYrLALy4aAdhSruUoZVu
mLR0jYMD8tlsVa/P85SjGiBs7957n+PuiQb9l43bo9k2z9aIjLQ1RtgGY0tR
fMLd4VB1hxMuw97bEUfdIlifnImuqwJpePcKdchtuKPmfLz7bu2psM9D+zwF
Fy2P87Lvei4+Efsjg4da+ipG0Pvm3OqNv3g7Uqv0pbFcEJRv8BJM6UAfI0cM
XqYofZQt8CAxbjbAZrKWqc5E1apQe5D4TL/ynujgIbAtxfW9nvDKl0Wb1QMr
U8b9awFsHhpPNAh1OaJnoHPsjma36gR/5UpE62NmIjA11sS/fD4fNuOdpa3P
SV5Xq7Fgl4UhqDaUpnmhEJ/Gwj29h3bLYUIAhY6njI9fCIg7RAVPW/O3OLDo
841xK4lZaoLXIRF2j/ht7HMDfN87N7VlyjYJiBe8/IFR0HE118PIHSggWYYv
ikYvriLrVg4VyAymyZwMhTC5KxAxptpso3fROpqhNNotmDOkLPX4vbLXJtv8
ZQSMql/Fdhn70LeBqSVGNEdQv/sa+xAEf0DOwNoxj5vfzKwgsJkuglzACkJ3
Y+0rWMHDSb/iC4Is/EcPiZXNW0Tk21HPAMHbOovi9BfHKNbVGB0oPWyKGtmg
1NqkB9dmM1IGqlzoVHlj4I650L2cLZLJr87RT2Gq515V1c3ozWAHqFeXwBH2
LYpUoRvCSOIufpTUdwRqdJnOxD3a2ghPAOoYAIYrsMNn8QEPZa2jSWi63vLY
TWKdrgYhFafCVlKsTKEL+3b3RehUGimPIsMaWv33zBQ5hOlYUaiwRRKafZ06
DE2rcVACXD9gGPEZ2kUJshZCL/hk7t3cQ2NDBHWqVEcz6xhSW/YW72H8fk+7
6lHAodPNDEDeb9x9quCYI1o6Bp9om681NqYH48j2UGJTVpCxTYZo0lFE5/qL
c41CSFDzsZE4xHxPrXCrJa6eR08usO1iCX8iVov1ruUlhhETDYp6YcamY0Lv
1cVWs0roWOeFGPjCCGX/MLFeGTTBx7RLTZHYjk2+6xH09K3ddSVkASX/j2UF
j8+FaX4UlLBEBUTX0GMFDrswthvEoa0t4u4ZA7GiSHIdZu2wd1o4c/afs/8/
l+HjvbwExqBSLMpsUj9z42HK0ZJn33oM+q4U1uNPCD8K5BGTw47fM1cY5nmR
Q//m1V6/RCcMGxUG3TmKlsSRpTZeAtlSnZ99e7NvYbYoPBFEtarjQ4GwJIAe
DpnVsyhsu8J5DOZ3PtfIjT0iEgzBbcnRFNoGrQEJdYKp/SS37kWU0dqDOF7/
A6X8C0b7rT0l/XqARcVjA+BhRJ1I9b4vUn/By5cHBAWWNkF5ooWbVZ2OQw8U
Ll+0dkp/URGKDKpj5DwspMhIk808KvXsJTdG12Cj0Ui2ym83mBHCz3DCBfu4
eoV3xrLpl2V2FQmPeUpmhtzEEmoy7D8PBtGp3DtiqIz8IzqMuF+TyRCj89cA
plQoNizlxEWV3dQfgWlq7QPs1CYJPAUTS1LgJH3Ol2JI2H69n1fvrmnhNQtN
qhh7V23b4u2VWE0DDq/ydmNYT1Q/PPh7FMFqmF8D/fmjr1VFLjtQIx5k2jZU
zskQv4CfwYrjD/4fbFphf+73CH4QVrHjGewvub6o2dG7xNyElyurFgtkjOp8
afbzs8GClzDdRYQjHtC9XFfhAAgvVf6pfROVZLDrg3EXBkqI5YuvdQQ9MwMC
HaYLaGvjhxbR/Cjg+zdZeWB/sFH9pMjMi5phoI1KFTDvK0357Ont3+58rIao
bBcPDzXZeEhQJPYCB766yV4X3xqQ2M07YgrHcB+mK23lfyfZVdt859tqjGrw
mnN8LacWBTC47zY+Y/naYvnk4ZY5OZernyaPcVIG29RumdQtBAH1EuwtuPXV
3YyVVuD9AffiSRK8PtecoEw+vCxSTxl0vd1d3f4G/G2YqdtEQ3nF5icoP7hO
3Ua3detCVE4vr+N0kiNMv2rLhD8umkUIan5HvkAp4mOZKasBNDVZVsGPRqZB
zSaDfY+mM8WTd5twobm2vuUpsCc1EEmsjrHTOmpwE/aRgWr/5flIcRAWouTw
ZuR3/3b7m8G/26xfdtK5WusBSL9SN2FTRAoetblw6OEzPX+vWtrc62f51Dy1
UG8zo5sVyBVAWisiOW8fkx/X2+M+TVIrtN04yp8IcSS7K3PVvAuWYpACuXwH
V11/qS5QfM1S4Qvddf7XA2Qo20J19rdgCRLrbtg0omDGxEsd4V4vGV1hH26/
Usn1W8ld3sb5QpCyxkyHpwn/1lRVU5kcjInrnENIAntG+Gs9voMsYBbB65Z3
EzouNHjNHGs6bCNsiWrKPZy6zxbNmlrpHQCYe3QaAmn3E3JOjAobjuFZod1T
ZQXJEBmYVk3e0UpfHYYVfCBY66aD/QBPBBfEE5KWgOt78NCXrDVF7RTxO5jz
+8p1jMAAj82VxLJ7rpNYZHQQ9ERox50urmiRyrQd1fktwrnmHkF6DW0o+YNt
gW3c+9WXi7Uhhj1KM7ftQAbPPrcR7fO6j9WxB4prDG1lk/M7A9f9gynlsmal
qLC35FV4ajPFlNkCsgG/Joh8U6BuKojmGopm0ulq7gPUZw+kYOAD7RezkPUK
HUBe5WPW5tS1v1op3saaRv4lg7rgiEq7I5/UkZNCHHtolJ8OaidcMLBeIGIW
pM1VtzfJpS3LSDpIUdBdoc3rOW5nZ5Lpw0/FvxENgoGh1iLFn0m9ccpfiZA5
Rc2i9fMUmSRyiJre8X3QeblA01mszM6HVNAUZlK4JScuEl5GAmnYc3lyQwKK
zR0tXg7+C7K1re2G0ISzuga29vcOwIznR7FoOHDG5Bwta9CbN8ziNk0WJ+pD
BJjGbPyZPYAHMW+z+nQJqKk323060i/VYklMDov59hSEOTCfZ3T651lkU6Ko
N9MFDQ18ZrQUmgpCHYG3aPp6bQmdEpCeVaFQnDUDCRrFnDaIQ1eZ7CV4ym2M
IQeHEBh2gkZbbf7qTcFsh5C2kKLt1Pv/83EPToLRjRJH6cIm0RgTMTQu/T2E
0p+wpHf1KZUQtDwZ7ciFrvqVwDP6qAPhdIpZQ9GgH6+DO09JNESy9hPWv32k
ha9LU0nqEOOnW8x4w2SDh+mkOY9CY92UdtCFWp3oZsBjqO0oeljKQWDMeCYp
eai3UAHuVAJFnwzsnDWruBaZJgEXtKVWctxlsNPIRvjmoIzcFXANaxRfKLPC
SdpgIjlInLWMsNYBVV6nB9nXywwjxGN4SxUPNqCmreZ+mQCvxvglkytk5E4r
bcWTA1TBAwkrH+6TN4CVhxvrZGEQUgwIjE2taUR2TnLAWPAaWpmVB59mZmxk
MxEA1aH8JEfwX/idIpWzV+cLLWVHvRJhlBvNAKSR42N0avPuRgM9IYEfEpLk
tQg6mBTOgfnZyEyvM2svZMT094zJQXKCA9KbqJsEWjI7kcgYLVtiR92i8hfL
efm80UR8wgC0jKZIS1VIcoH759RqqAcFn4YAZH/iwzfGIhdtXN81bA2dmfmA
NKjkrzzQ9dJ2ZmGZPZy4L5AFbq4/JS9MutEEtU+SUrMKTuA/UjmPUDagLjtp
1XbQk9dhedMEoPVD8ccPmUObNVnf1ZE6Im4v1qGtQ1psXNp6lZ88my5rqu11
10tggxqtB7L/Pg5OYduEkHFpvn+SigVnbC5KhA9zjzTS++mTSeuFnCCS+XKd
QREigPU352RKYxMPrn2Tl5JOaoOonWG5PUhey49OvHmtmUAJqfTCJiIMSfKO
vLGNdEU2bJqS+l+8pPMByD6tAUqPegBlGfLskSj2B2BjUOSLqNoW3AyyuL7o
ZX+d5jzfIyff95EPbMm5oicBCMQHFc4r9ijbrBftqYFGAdAqnWnaJaOiOLVK
WzjTvX7PqTbgM/XbBXFGlo2t48H8Si8EAAHMClb3ZCPyYU+p47RmLnuWvufC
rh7w2nU9QsSwOOJF2RYbYas2JluMPW+QnCREXQ4Ppz8lcBxz/bcZoD+WXCkB
rGrZYReHuNYUp/ciU05JfVjn+zOt535LEH70VOfXwDUGG67UJ2eoWbpVV86u
AvjN+D7Eh2pU1iiwk0+JgdiStrG7AWzXAQh5U1jUH6egbF/K8O+1Uj4VxtSf
pSUsdoxuxKdQnTh/2navEZrXCV4m04J+PeyLMRCMhNhwGDB5dwFgrpS0KBqY
DrBJ1jVZQX5ze5TK7IOHY13VxSkHPDwaXBP0+klu1HqARqBRrvTN0PGaSR0c
Oe23EGjYb22K5+I2FP2mSyR+ECEjgI0owrnXMQNvp0zvo/CQwc75ioVUw3ll
KEabmnoBcby3bXbmnoLkcsR8EB8m8lxmb1/LCCoytjhqEcoBwnYCFpTIutO9
7gV+yFISPaDBsC3B0fl8ugXCQppFO4dYQbDgyYtsXrT11g3gU5t8CSErZhtw
s24UMMa0wb+fPWOFofLgbeEeauCrFnpiVd6FtmSGNyOUSnBxv4p9dXOf8cJ7
CmyfnC2eXv6HZJdos/1/HN9xMYbgtK4CrF5VOgJWSjBN9eXzdaPlxBhO7T1V
ZQYluNfgJ5UICXyVQiEMkxrFVMp1938lBFz2wJK7KDP2KK5ddUviqa6MGK2U
iuTIrG+BLPQX4gjIHyFa+sAkQmsWiAff96pF7K5vZddmFaSuoip0d5tSotT9
vP4u1UcAcvLk65dolt6a9EsGOHTbkVmT06gpguabNzEfiFV6pYLSaIEnKe7D
ozZz6JL0iAyjjUthZVefOtj66ZdU5TMsM44ifYXcUgALsYe9/ireZEVTLfUd
SMgnigX63Fb09xXD/jNvtzWR3KFf21R0i0H/ZKHYKCZdGZgcdrBzXXC04x+5
vE66PTM4cl+bqCXfZr20gBsE2F8y01LtyaYX6bDrchPFQTaErRVQXJQ281wr
/pgJFOdo6ehkvn2A/Ovq1a/oSRvfqCn0PWtw1gOO0ysCL1aBh8hYUXXBOURs
AeH0ttH72QJs91JlQAPb03WYN+1UjJjREOpgfb5ur5plY2hvWFOvC5kMwzZy
Q32iAH148xbFdCZdn/89gTlItE030eZdm1WnLD/fDG3fPLYzp1zRV8TykcG6
X8oD9Y47RbQgCO88pU+qOMqruRzclHOzhTP6u2nrGF+WzRk8hbUi9ISAlnfA
A4Lk710vrOBkhgwoqENiSKdmrS+zJVQLCSWP3ITs6cNL27/yTw1T7owqN1NN
a+J4OqerJZwhvu2rRqiKP9dqsJYzovcWga3+4Mh29ZWcbhwDvDuffJXZmJ5V
O/9/NWzyQUSDVjep/nJjU/+8UG+oLeStIm8Un40K4z3gDHPZEpz5YnNY7jsh
zfcrsyd0QJwcxVrr9WCHbHG/0kco9aw9PATvtFIQesF5FhFVdcJdE31yAkWY
YJ04TqklhbmgAl7SsUbTT7wVq9/J3vcvV7/ABQz1eu04Gv7/UIE9eEH14Tqi
RcumP218LkqSCQIbe30t2+tPw+o5cJWeyTn0noIBKKDb+BQ8xxld287Ha7JH
F9HRvlCqrELw/clYGrlzGk6PfJKdqhDMKIaDXixwJ3aosNabXR8HkeaITkR9
t11xUYPohtU0zOufXWwxlD6m1j8e1EE7ohw6ircisOcuN5hz1nHMzLuAhtCM
RJ1dKcK7IAWS7PC+9asJ5Zvi+f6pBVTVtgTj26yHEfHRg9soko7RGopgg9WU
v0YLRR5yCA88YZL8X+WdvdtRNQhs4+N7W8BtLAt/pajTJPa+XSvkTQE0hfda
55XQinerR7sylt1devtJLPbXbS7b1JrFfvvpVjiu/aY5w1VYDM7F4gmUcoE+
KTX8UkM7uFcc7188ia7Y96KKTOT/D3seRYR9iVhkQdWtjNeZU4IUkMFzccAJ
N2riBD11/zp2QpIDJrAYC208P5y5kf8830j3yzln7ASKc9gx/0f1Ks7ACqDV
iiE4dNdi/HocI/HDOF0Zw1Vx7LW5ZbzdCY8eKbYi5mo93d0nU5xoC6VZr78O
i2FoJ2EPtU2gXaTdVnjrZyo3E/WcRK9Z4FAZB5fbLfr6fPzRkDmvz5ROshhN
3dcYMDbiuCci6Qu2pGS8hPuuwnF2xCSq7NB11ENf5h3rDgCEfhNEz8a48NlJ
ugUhC4St1dREX6eEZrfXQRJXhhEOxT7YXCUgl3MkjiOEWYgaPoE+sGVt8/7n
6yoQyN+m4rVZa7iOa3LIhxkuKhBvVinZRQumG6Rk2IGGC+KaalQEx46epsfu
fmpsjQ20rwTtWS94iPPSZhn3e63BQsmSeYe5zLkKbQtYilXujz8YuqMYC0m5
xY6nh5RVeXkW/jSF5JREm+UuuwigRU8amo4FUjjZlKiGDce/dLpd86whUfkx
jUQnIOU4tvSzFVwpDn2LkSDFOPd4MhLBIc3MEkIl3yAhYTXPqMabXjg0QQFV
7/ji5STDTimq6JTahylfROTrvvKtmY04NuTpBhq5mzKXaJsdKBYrIjJLIqg8
u+uTQWPAKtHk47l0j2ETJ8E/SO59BCyPKia7nWV5s+FnZWjALJm43NVPfm8E
znO5KP06MyobOC15sD9MFHcH1w8VlgO10e7iiw4egORnJrLsQyMEaU0qnw3V
MLoGu125QnzobMh04ReY/uEjNzHPZYI9uL1MyuxYLZyK0XcZyONyT3ltvTp4
C+7vZpWVh9s1wuDSFdIwvbf6luGGB1Ywk46IQsnfoSz2FwvQA5BEJLoCaYFN
TJcb+sxtG9yjMJJ/hON2K68BGUsdBs3whHc6ibX/fEGZQzwSDfdAY+IpEBpu
i83E68nmtKhqQ7ewZzzjafpy3m7F7lc2aBCe8mzDY53yP2uWAVEOOdcO2lnL
r+H8izgKC+/RCcmyXOH3bYsgdie530+VwAwCehrXefgDKYEpnN6YTl94FFhn
+gIpU5S7BMANEuCFab60w8otu/M228vZpsnDlN3LtLk1TVHzF9fRJlST7tVg
ZOZGFTax3sy6YRMvoM53R+oFYB74c6jplqG+uhc3KqihyheQ2aJGifbXzc+0
eMW+gcGX09jQAXuvEcU3G6mJ2ZQxVbKUQ3gTOYVSjbugpCh3ezm9Z1q545CM
14D/x7roMg/hiStO79l8rT6vIkDSZkK4Atcg7Qr5FM/AbkILX1T2YFIi4Olk
b4Kuj7W+G7Gp4QlsQT5g7ADUIzJQwGlS2TZo+JJptxhvAGycDuLDyxZKmFRr
si5bmxcKR1aGrqnZd1QVtfvNWoCbD7X6sz+BrcjsE+2bxYcVqBg3Lswo0pqa
+JoPsS/v40KtADNwTUP7RPXZG2prMTIPAudAGIVJ4BMOdPRY55ILi1aTvYBc
SyyJLkIzV9mPjcjaxHIDkqwCn5aD6NiKj8TG9RgvzX2feWLS/IchU9qQqcj9
CIKYpeD6DatlHjf3Q0TdKA6BO/tjz0ETe8dnhMsWOqLyL2XrKBzugpWO72eM
k5kzmSfXEQHs6wccQL3S9IJlELqVWmLlE25pfuDLFKZWhxAvovDn0BPMC3mC
iTCCh+VOovpl23HKdv42pdF7NhZqHEwFSWUeSAKDB5+Apa8azLaswvj4jFnS
Kwzrl04kw2Ox8XFaBaUenoW2vSBncKp+/s7fpKX9k7mNJzAvphPOLGwX9x3E
AIkFXtWIIaiRD6Ws+/siQFpsY5Va9xrnbiPzP9fsgQTK3wr1iRyiHIMbkZbB
qGD7HqdWneHO0UcoTklmnsBb6emT1Xgd/lHAwgVnIiGdUo9A4g6ib+ZRSgb7
9yMO90tvgGnyDicRrL9VKqx9KoO/aT0w9lV0Z8Y1NDFG55yvjfYgrLhEev9+
T8R6lgJGElUxEUdIXTt4mZexdVKHR5wXfTc7J0AWyn1l0REOLGoxxME2Y5+V
wO11wolnehljg5e08iSkfyKZfhh+y8IHt75V3z+lFAsluIXdP9ziArzBAMvG
ApAB7GN7XNf5WCnsmcP734WYWWj6N9T6K6ujTlUuLyoFTmbcJQov+jJgfCYu
MiHfuoKp23uOLnVM/URo9Vxp9tHgJYeCGQler9orM+jgWSe7doiZ/kI2GFoY
JCld8A0N3+FwdRmELDb2J7sGbT0KvR6wQGWCh3RX7mwGCktI5O3spowuF0LF
6OlLpgFWcUxps+5JHyUppzYOfonWRsTj6wLJtWSGLDG3EiEg/BSTOvRA4iSb
7r+HFL870H2fLLZ6pOVHZpWVOgjOmS7OCZV7CMSEkcogE6brakr3VyVLSTs+
EAmDyY62IOOuAaHSNwZNu37ZjQ0mkXc74Pa+Ez80yIJffVOQ2Yazp3Gv7tZD
g4PvGD9L5s3jpw/ujbUIpCxuai4QoekH3mInmZGSZaU3hVtw1lQidBIRbz8O
xG+J41GkKOX0Vic4Vt5WJJWQkUieplS/5x6I74R5tYA9yqGsXvyIyUQ+MLFQ
hle8qoXbMVji27lxr5O/9YjSdbruHZFwvGgywFSZ1mDwdruApPtLAhwXxRyd
hy65tqYa33p5EtFtv5FN4c5yTNdz0u8AjvazixK7B/LrZ4yoiY9Zd8cYV06u
nxQ7+5r6RYL82spZ/HxfCtkxcSDIHb8yeGU4zlLGGkxVhq3VV4QCxzOAFbMQ
fpH5+uLTMUMmJgiI42s1Ks6huW2S1cT7jmo2UWNnnH/Fmwn1pP1dad9hoQxY
HQkv9SYwaTslyv3i4D8fVcqJRW8bmOSfUd9a8qTG4m8CqjJCWBxwzlfh4Hnd
4I5VjANMHA+wTQ1pPQjykovGRoYO6rMFaSYPSqtCcSVZBQ9LjTO/dwpEDrx+
uiOvN2bDx+JLMG4Oq4z0K7GKju/x2tyw0YkKVucD1WZwLfy7gElZJfGGFFbF
/02b7oMoujIk2USGVzirN36UzmVeYyBTkvOwRUtCNycOvQJzMfCRsI+PSQOT
V/xj8Lso3yZw5/W7dc39FEu4K3IoX8Mq2HTpWC+TUpC1hH/F6ei/pvD9xwOT
oZ/Zo7gxFLDPXSlUujBg7LuDZ5Qxab7IWDs8J464QWTwKQFoGywPRhYErzTu
FwwBnzzjL9qP9GEngyLRmYn0a3yXnAUetuNeUxAJmjjwWYrBxxQWSKgKH//D
31rwIPCqq6eOczXtXm4w4QG9eruiE9Es9mqHA0dIu7/s38Xsbv4TJnklqvpO
W0kSXS7x9HZ8638BOjHWYIT63Kj7oq4Nh2b8z+VnqDoRZKXpgH0SIZQSU265
e9mvSORDti+V8VUzCyhha1fMWxW/8H53Oq2JSssfLyntUlZM6WnLOgMk1c/b
CzcalCqLn9vo31F0JOxkcTmoGynVt+K4Rl7nnu7b4MoovuDfU2PuLPxCY9ZZ
Xe4VnpDrUwS+DjfG77L95GcrK5l/OYGzz3B2QDhwj19dVHkt4y1X65dcx3gh
XS7cjCK5oTPNdAOLz3L7pRlh7HTd+exVFZmmVebHBkbtm08UvMsvq4AR4yBV
1CmyjtX+2p660CykcxI7Lmz7l8cLoIS7lUrfnPux5oc1YC6aHbY89dQB0Rws
2XFVATZ01g/CSausBFn6ihxH2w6rFERm654MHIU0/5HARgTp3I/ROjgzKtT+
Zcv6VHWJiHeQ4kFEn5OchaMZxGpv8byd9qHH3KstSHk0600SaHod816f+pyG
eG7cDpLiCCYcfrvCNqt1gs1FA8E3unOGdbCUR0F8WINOWx0S3jr/o7tHu7iH
bXJ3hywe0u97Me6wZJNgzA759h7Wkl7gaNo6xRqiJ21D7dgKuttW025/peeK
KqKqkn5w+7Jwom4c8M4eSzuIRRri8PNtbYthssI3CiEHu83GHdgfMHDZPK93
17+/ChJydzf9ccDcZn2ZOF8hsLhgBzuJ1pN9Ww1npNmk99k3wMyU5hETGAmq
DLHIacw+Y+IhoJniwC9GyPNRXc+6gV0BQcW1KMVy5vgYycDTzXRMHkGf7T7E
w2CNJaCVPejzFXZBznxms0l8MuvgPD2DXp1kAWhgAvh1S1FkT10N2xwUT8+p
nHjIxdir6y+skq80Nq6NhhGpqvMgEjFU7U52aVZ4FkIyx08/74g6APxgCpfw
oeTdFdS7+mgmksfdjd/WlDwAhBzt+4dNK/AG9I5Y6swxcVRYSZO9h91DnGjl
LKPLPNvpksJWN2hO3D1RFCqSUTTYTuYxMpMfGFtoSqEW740662uN1xw83I1D
LMQyMrNiXuXUvFWoynXWJviVuXhNhzUE+ugrbDp3gorm+VX6wbWWpuHwv1sb
IaiP48+v7kCiG9QaWCk1BQ/ka16dMJN4ygj/IsQ9M6y1QxE8hXh9b3OT5Eia
mRmxlUMU0urxD7dX4Q9edBCRj92md7mQBs91UVmaOm640lyGVlyBWfmoVZtI
0t0UhKD7T8Il+XTXILvBN5z5QVrp36pwXAtSTY7v2GfgLt9dIfEmJvY3YAo0
oCi0+9+16pHKZ6NAMT3U8NEwZJdqC+4YhrCcVZj4PIvj7fgu9K/LqROTs8H6
6MVh87Mo1EoHexUOAtIvD3Ah2PYHmotwG8RrOcER+R2hYj+b8IClDCMo3jeP
jJuObQ96fSDcQOryEeIdR2ds3gUyNwHHP0jEcA2DGom58zIH6YSqC0UouVMk
q/2mU1o+zcYGZk1n9pFRZbcoDIfIoR8jbZhEym+Gb45lbPANpfdb0yX8w2zo
4Tu04WQX6PgodyILjHLJooMVKroUtb3tJbvw0cmecAjUhdVPWJpghrILqIYp
uUXiq7jDVHxK+DdEHJqN3Ch5AfeJJefHc+nK5R6uX1oCIYyvJlBkVw9GZqkg
xKJeycOlAtmjsiqJE0+foxILLgYeSU6/J+KJVWRc5rR9dRtCCInhdyp9VHwA
4PS2R197qPvNgiWWrOTNDy80DcuwdlJ2CDgSBaKuQ6jq2sHD5s0YI2S4emJn
zNF1C4xgSq2X3nMuJ9rIk+5x1d9WvS7WYUnSC+w2t3H66a7xOovAnO7QKODY
XwPccBY65UV+zKARuCLdf1oz244QIGbGGifGFZq9LFV0VmQLTFfdjxPPNXFr
I+uUI/NTlJJNvDdpEuZEoCQVz8Y2pp1ze4KSUBGaeKWvoRVnl/t2I7yi/1EY
mPItPwm+xbMu8nUXTFrklvQmTTu9HY2Ec3Q/tb4nsrgEVhFxwSW+La8f7owf
uNODWe3fxrOaz2oXYU4ZXXssWy5UG0EQqYQmnDJb3INvaukzjlCPoVQcyWUs
PyYBhhMq3XxyPRYr3DaD9DdHegXP0BMp79mYrJDqxOjV8CiAt0/drbtB4Mnj
RzzuOqCdntVfERu1CZi5ZBZgYyQNtc8JvR216/BLTxA/zEbPF2Es3JsAfZ23
ooC5yaiOWIopS6LzOij0nirzUNedwUCW7vNLgMRxhcA3MIvEtmYY6cXqMyxG
Ji2KfLdg5XXuePdKABK4XBJpQoDDpirXK6LiWwG5fSnS8Fe5dHL3mbCuzBrO
c244sOaq6YAMQ4NI5tSnvMWuxbWXQ9OhE/osP90Oy7q/WgPw9V6dE184zvQv
yX17jQSjzhJEf7Af3mj92OVozVI0z/P1juiRupiMlGYI4D6vFs71Ti1BSPSl
MwS4ojJgTaNLqBU+SFrh+mTwTAx4BW/RBeyOd+ux3yQNVFjSGxf3WmadNiJe
3Sg2B93k6Wdd/dVuShQZS2qejhkP6U9kU3zgnVKhYwNGux7F+t/uzARTKEQy
Hx0Ib5uM8C7vgDxAvMK1ily9uUuNDUfGEKWIYjAER7glr7p+7Ltn9EpBOCa1
W6Z/NyXaEfXz4g6pHwB8T4thgOzeLQkvJ40FAjGl/NZ91HsbmOZGihyuMxQ4
RJLuE0NouXAoU+o2icMFt0FUbODEVenHDoHzrfYnLtTFHP4jLzt1tAR1lfae
JSarBb9T3DjgPyJMcg90X50kmbgPHkdQab1AyP85sBTfChdaKDozik75d5hg
/t3so1rDVmlBkR7saiZAUhgkWyeAfnZNSbTL+fnqKwhXiDgL/Pnd9K70OD+S
R/T6mbixWQXtyDF1XePrF7nJf2+vfL59g3k/lsPz29LvVvqf05o8DpYT3+HB
HLIzQElsIeHtbV5yNxIucnmGiF2DXi3CHWcSaZGwa8Zr4gI8yxUS1Aaq39hD
eOz9EMmey/3U9osH94Ut23tmhWbI/nOKE0co/Qh1clVDlLdR7THzvidOyd4X
FO0Fmz4rvhkoXITz2sg8FoiE2oHVbWyyMwfKqI28sAJQjnrYwscRurOQKKIj
gIvd58jkQ5qxOIt5cvGMkXX2NRWQ57ijT3+s29hHRgY8OiGUZPvgVPqIKYo+
wmCgDZSRmAt4z5rxnPUWp78cIjR9GSCDhkVoSbI00Ys6lPsVxLdtRuadEyzT
wbhsRWRi1A32d8aAs1qNH4LG4XSm71LuVuWhKjv10R1TwcFo7wR95ntY8uIr
nbHKs8Xqvr+0f9pSWnwvH09rsQ14RrV1xColZIh7zkgGqD+gC96CGDaNphdu
IjCBt1QlQ9zoX8GBgNsl7PP9O6wWW154+i8GRitAEi6RxH2VYtg2e61EEMDX
hnbr6jx1vTq3VN6U4AL0tIf1pqvnUJR/OudCF8ICcG8Fvn88fRTh0H42D31X
Qi1rx/vmKmiaIJpLXmpgIOuVe3Z1tpZKsg6/SCCrZWzL6Pk6VY5VCr5Y/Ohh
gYWuvFEZnsHx+4WDZhSdvrVkvty8v3TJvZs9gMWPDv4PgPogHJyiyLRDwfLy
eXy5plRhaX0LYcIZZHkqsFTnQrgOQcmkzfWIpTVUq8x0cTFiBTPVqf7DfjxM
HJYikd+U+2jvsX91t9X1ksS5PRlA/KFxRtzVmn00xXTiK/I+5THqdYG835gn
mSLWZpKROcACzej+hFzXcAI6VtZLRB0wUtdrpEaO/c7uDxd7kF/1mr3rvTSQ
wavAzBsTuAa1T+I4y1Gvj66/UIBUzNVOSSoCLrZzQF+gt4z8Tq7w0gZB999o
kF1E44E5GK7prulQEi/6oApLxvlQeDJHBWNQ9MBsvPZdxSiJhuYK86S6oqoM
3pm31msNO5q/xt5pc9igwCUuCyOhJ4bfMo993lY+xuO6GrTE+TFaRWGxMWqI
8+Xy9jiIY0APiBRW9qfVQVNLDn8ueRH9UCUIs4r/ZYgu5ucmFAsGqFdqIFhc
B09vaEr9nxH+FHuHqgvQb8T07uf8IEvAiEYYOn5B6rnrFFpf82KJ7BOglzKf
39RfXRPaAVH+xqDybRF9czVMHYDXWlD3Gp2uuI4CFmmK/3IJNKv6MhW/0GSg
/wK6YxMu0bH136Tsv1dp0BjKGe2Qx6LyHH4pi8tDo+J13pk31u7RkQaMN7qb
xu6DyWalKC8SaN8XV6aXpqU1QHDSPrHdLP0jJjH/FsTWIvqFnTaDYWESoUTJ
Ty+gG8h44xGI+LL0ZHZysQ7BwUngNjPBlJtUDt6Xzvxv1e1kdv+lyjGN8GKP
8p8VL3NtaxdjHP6ivc9NkIdO/H/GD902CRcqnAUFQFQcEZQgjvpuFxibabWm
BdH0tOxK7V7PeXGlXe91NMKVrV3Ujklr+gvUla263oEVzrt9IeYzOWKeK39e
X5UoJxwtKnp5ePVoHFc0DJQdLMswm9KgUCLDXxE+PhF3fwBKgNleSu61gQ+z
CPm9RjP4wiq9mWLWHwAVb6KwRHDLMtnxXld54aBnyD0DEoW2YdVQGDBZ4NVJ
zyb7ILgawc/1QOJyiXBBRkKFO+WAfCApTSxbLVeGcb5NCJgWObfX9u6j1J/9
Mks4OSI+wI3s9nDF9zBYTfabECa+UGq4uot+bLmMoKFh3V6zox08sfYVxiHi
HdFjDpZWBeyrZL9s7pKY6n01+1Lq4wI5i53rS4RNE4tGs0yyRKWmUJo3HBdc
iZMUlt8hLEax5R1Rl3iWRUHngbTeYr2vvrmdGc3Mi2YzJbl1efi0mdo7W9qh
gwi6d0DgWbwJnSrUjehbI+Ax4tSzen3Prr47eNz+npzUo4NPV3YcvxCjMQtK
w3tfdVspUlhKUNd6qlPEMsKzf8eNgjr1bEAczmCHAgkmjlxFR2qz+6k+xC2M
q9XuPJ90JpyMLVauCR1x6Ypk1UZ4k1UZLlKbeGXR/BWbawXOrbBbtwOQDGxC
p8o/+QguaryByF0vSHgE5UXGUDEoDGREmZGtS+09kJreBftews0HpjQvoqLw
KLHxsTkPC2bNPyXQlccwRpaC78S66bjLm2pVagzF+0YqrBKDN1aPnJMz5DiT
HkoGaQ9fTnO83jCI0qqq5bnob+Q=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGOq8KwUedUxfK3/Ad2z7hVEmkEHyrpNnbOZWsqAjRjPUeVoNApd0wSGfH2q4W2THFzSHm45lyxRk5Brt1+U/nV3zYpXUkw5qjSqYg+JTQkkfLWievAUP/RKveQ1IcuEkxHJEXK6BmV7B1BKQjHjbFdCq2m2Wy3z8hklu1hqZ38tZpSDO4WyNBqbIa9vvpNY1iYkcxSp+e5tUwLl3mSuZhqQlcMOG01rt+ygYC1UL8RSFSGWLYfZQM/+EbyvRa0agx6eEBrzp8Emt9ONYTizzoavY8ARMoHc1KTEmhRVwDfCaZmhk7nKiZ457+TvxRIAsIa1/OC0Xx9OxCtPrnRuTCHyKhHZMwQOPaoYFulDqxeZSzwBG64lWyz6cYhX0SUHCU/GFZeTbAqMfzez1LRzWe7GE+/k3gGEhx9l31Z6DkemoADm9NBIaYtQZbf0NHdBCw+kGbL+QkWbBn7Xbja1yM0yEd2CNfXo4ms3Ntpk2e93U4JSJi6MVTzQq/elakJPLucvkWiL3hzjFsGRGhaxheyDiWo60vbTrx9yrteFgigKbmKgPsT3wRAEADiIiKUeVSO0c0UoV3uHUPmBfHGcfhcQQVLA9qe5TtdJsEgV2gO1Y4uYmQ4wPqn89g5lkwlCslCHApRBvpl8PKgLtwNNN22S6ogR4o7VrLHtOCX5LuEK+K4YEz7NcmXC2o6jmUkz7B8SVsGLYWGndSV+rnqFj5hrKowEeaPMFd3jKMx6ISTXUABQGIAqKXE/xvTOBtogqQQcWFgSX1Lz8fXjUPFfql47"
`endif