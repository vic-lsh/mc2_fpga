// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xQon9sbqpjXSbAeJaeFu0YV6A27haoNyQG0XMM4NVFb5m0ti5wDzV7tJPCgb
KI1waA7O5PlkvM/bmSTCLeUr7P9IBN6Hm49DBUDs1FBSw7gXEyvq/cTwHZK1
sFTZSYb0yZrMNY7faKXyAUorWIGz5kSTy2LWz4pMXKltNWpFZKh91/KMbIEf
66LjHWDBbHOxdO6WSD8VwBav99hLZshr5yaUX3CeBu+Llgr9ZGVgjUSsSTbh
Z0cINFBV0eZUhejygbI/lXBMVQKKIsRf00QfTAM5Sk4jHfs66JEBc2x/Pfdk
018222UnMFkyiKDH+j6s4qz8x2h0/b+Vr0cQ7f2+0Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VMB4XedDZNDhTWE+4XHlPDD1xPqRaZyHW7e0KxTpONBmGxjtlKmxYAlidUEl
6U9kwzp4kQe4pD6UqErQbXHpyyjY2wni6huAh9SW6R5VZ3A/x8tiV6/Cf+H8
rnIlZRGfcHCIQfEhqlBVUp6QCquoYdXAbTywFTDTLNJCsC/hT6pIicNwO5tK
lzm6sE53/6jvnIKrgYII/vI/oDd2MzlyQ4rj5cKuRBjkCnpyxHgwN9vpzfTg
L5274y5BKC6Q69p0/spJO24nUaEvXs771Rof7MLYnoLqsYqLm1rUEFCCZdj+
DS/nCVUwTmF45hVEiLbijNDvxvsKbjhCbpWkD8nLcg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NcHxM7TjXEn4fDwT4EE8j+k72AUPQWGo/cSMBh5cxaChN/vdUiWErjypNX6U
Q2CphHwmSiYK1O99TAuR/HevUTazdmbbYkeKHFcP+EmXboS3IGU/fQmWJ8+4
OH2tK2gSbAq4wYo1o4JjTMXta721eQrUu0YCQX8fdUIwjnRw2wy4tYATcpHm
rHkF1WD2U+knx5rYJ7I1EDg7h3ZVKb0ghEjpS45BNiIvVPekV7xYGev7OsnU
IvBZDccf+x/9oDsTjCNSUyJPxgH/puUGf7+BsRQuLQmfpV2wRWqUej+qU1zN
hLFp2IBdMMtCw47fpa1zIVWVsxYpXUtNwtUDz/v4MQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XF7Sf4xML0wKX0IV4NOytxEc41y7/53RavsGY3jjNEGJCuKwqprk5e8Zn/LS
mG67zZn48PedlGtAHJSADm+BbZ2uvAM2ZulsJlxjL1bdKBxdBw/cU/t7NuFw
Cdj/u36GB5qwCPUSegTsb8G9y78d3koQc1QykCjQ2X5e0Y1AnW92xMQO0jXj
eEaqaB3lmecI6Fv/MykiE/DRBZXEAiNrzj2kLJL8jCxGr11qWVSbgAZSJJv0
bZqp1VEGrK7jsH+nlYecZzDnywIcDpwSUt7zh8AYriu01td56d+49Yc2Jx4T
HthGl+iCQmVtiMo7zvuYOf8Rya8tkfQIOmEJj70J3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P19UTaIupVc195Z5vqo9zBpnPXbnKgZDJn99T6YuH9XLE9tjymAJgRdxsNeT
MEqM7q/OIrxuwtdZbxD7EaS6vjkoefe6VqMf6yHIINj4eW2HiPMJcRbCTdzG
JzgEF01ZkPhpaMTy5vpxruz+YnIk/G7hQtuioL4Y3mJFGjsPOLg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pCaiLfeHzWfhV6Om71lsQpHYcTzyORrI4Z+igH45WwAlLKsF1vPJwV47k/mw
syS2DKX0IGK2bctouWYa04Yrw6n+p+cfrSsEy3xgA99ALc902IG4Wt0FQDXd
CawslkwCO042tE4FS9eQ2dFjy38hnulxnd+afEyo+P/1o+DFc+wfLnwdP/0p
0lIzBw3D/QW3LPVK2ZV4cJY/hIOlogvZSfvOHxb1SlYLwY+DYozAatZ9lY8n
yb5gjJrEa1p754kVDVCpZO9ZhkK+Yn5lkgmLpjeGweSoanFV3oagz8KDMkwO
5tWV/p5ea8oazrny6mxx9OS8GcxBPMB4A11Q+AE5CneFJM6HIP9JrrJXol65
J2OAL7vRtPwm1hYwdWarLOb9G2WS02TvygQQ9wkXUF9BDoEG+3fHk0bWFN6+
wODWrdQEi7u/8l0aA/QmffB+2Kgd3RaJbcVwi4rHJdYGi02I3piqWnhtFVqP
jSLT5PWyhQTfkPrxmD/M5UpF0Q/N0qoL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r7XWUMGTjGAItbQURCU1/uh3ZI03mqtE4Q5TJhBIxFAPmfBgZbKikZCBdngX
kzyW2yMXPnUFJMyFvS6LkdPNgUC3gdcm4ZNxSAqKPsgFJHTlgKIT4FC4nt92
iqcyXICblExnU22YFPCXJN3MY3iY7K8Qf7Jr4jyJJ5H93aXOr5s=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hhYC6h6/Ms6vc/EUyqfN2pZRCkPnjquKdLoi1xUMGqq+2BnP13QWhltyRKdh
X9pMx/54hq+KCPCTvHsgWe6xEYzBKccPxyDEc9pc4fea8QTRF67yE4KfiyqR
+OYGaiaOwvyE74A8IE3kg0eucLv4rfY4SLcpYVuWAqYqczSt73A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28656)
`pragma protect data_block
fBixsOtGO3HNDf4Gw9klSeQUPyEgls3ZXtgpk+2zD50LWINUKGRRm4R29w5c
suafJlyd90pqyLKyaNWtdU+nqe+1xz+7xfgFvBUAUwdgvEzx98Pq3Ci1Dtvi
BoxnhDWYiRTlTBjiVsIjOME78w7CD/tYTkc8jRO5v29KilQiwtJIT9pRTLPB
wEVOPP7on9w7ZonJoccwGCCOXZV61QDba3SIZPGsPlnxkSr9WV7JqxyFQPZo
ZA+CgtANHHD/kBHo2e4Sk7g8RtMUP3m2FBlaC54fF2dhppbVJih/A77PvhFY
+fdojiWUrAXqKuolOFeqniIOoe1o0Zjwjl6b6aSFhInTWw1xZlBUGSkkgdiy
WkWUUPKenL+lTOlA2Xjfn4Ek0pl+yGu4q++ma0mGIfd+DBRG+1tfTBetUXZv
d2WY0XVdeohXM46jru2fF+dHpNrmK3p4w1inTvFpAzfY+js45AeZ4Emb6bGJ
Wfs83poqNMO/DNhnvqX5a1+a9gZVBPXKkUvnahh6hmZCsLf5vRE3Y/bi7KAL
mmGS2GsGAXP5CHFNN6qUuenwB0MDLd7HvW9uQ9YHglqQ22MCL/Vonz9oGnYq
nbWFB/y6OAvJQy+Rbq32To+PubieEx3miBatbwRVbSL6UW6sAQi/1P8cl3JC
ZI3zByyUYMWDMoxSHia9zcg1CK7rL6cnKYrjLutuKRHHrQ+S/tHZrx22AjRz
Co31EQDxTWU44Pfoh5Ndd7Z3Qy2BrxyZNRxOO7gEg3ZVegAS5e6+4T4QQNiR
q27Oy9s1c+B4OHG1nYFOmVjGunqllmYDcOaKS4jvKmZ4Mo+dGfyK0spobbbh
jGWag85S1O1tJyn7nXu8clVCyuzJaKG2AYBRTI6WN7kWWh3HRRZ+89f9p2Oj
pikwSedW6HKLFqSnjXe4YOtxy90nVnr979DeR0PFT8Z8RF6qqC8KEOF0XhGC
GD0odNxY40aYCoQeEUWbALJU2ZCxaQzOXEBI2XaC/cLCmJ50am3XvqqeAvbI
N95nKIX99SiyGIsJ6boMjsxK/H6itDp6n5EIV5/u+Rlrtwdc2ygEuJggVmvy
cipu4DegTj8mNXyKqe2usaPqWWMYuyRkQx6M8ZlRE/qalWOonP6tJbLETXlv
3ZWWsSRbmywRto6w3IXA6cAaODCzR6gc13lS/v0ouggepyQxS4luVftWfepx
t/Xe1lGKYfnkosvK+i6zGpesp1W34/8GDZ9ns6R3jfM6bNiOPboS+9I445H0
MS5ekz4a8AcuFNBRAvXIk/3YQwb8P/3WE/xnB9nyAjLpDgyVtzYa3a2WN7gB
7vhoTIJOcZ7tlSautGypulKMRkOAjtgOzHEYSevQr/3T/FDQdrvFipxi+XsX
kCksHJ/gfx3jnmacWadfZ1IEcEWQT1u+qsbCuR8haUmkuvlbzE6QAFG8eYRq
vrj5r0i6mleO5UdcH+zhIjOQoLOpZE2eqUHHp9bKxwQ5pCqVF6gVyROzYNJj
NSazmmJPvq2kYG6YrB52KWEMgGwrcCWkLcUllrYqZw7LhI9EA+L+MPPCy7VJ
cbu37otlOs+xJA3k5jlQ4J0DCr+ZVtfMglIPcMlk208f7j8G4fedKQFwq4XA
0mk0RwTJ7Zj17FwObH0OoldoH90vlUKwNU9MhheEPU9nQn0zoRY5dwlmDZbv
PLrVa6Bfx8V/jxF6xjvqbA4AS7JZHWDVCx03dVkCXseND9ZrpxX7AVkRrzpr
691GaTwTmNmqVkPFN487aoCcwsaj5AfaJwhN53K3xJdufs+sL0KmQcQIwHCx
3V4y1AzSP/zVQvL+rml3i4K4fmIRLSNX88mTFk6p85PoFxgqwTMkj3IOmuGo
eJ2iNDMRCXqyWEWbUoFqi6LgHtbqO5MuE5BSj7Viu14nRw7P26PIWNEsAeqa
vFs4cOcXFXVSwPDKYKbjfhwvSDZgoDXVmesaNGZKVErLCJ/J7vVYsu4QcSS3
aPg+hhz38eCOSzdDhcQQz50TiSRtbos4OisKtnnJf8OS1xSXkW7YM2HPd7fp
sN9Y+UJlLuG9Qy/lOVxIsZ6gHaUQxxTvmDE+lDL14zUfvKSrM9MQ63nco9QO
RWo3JVFHAEyaodSwKcRkMTT5jZR6g0cRXzj5GpQqR4+n3cMrihOEzsiiD1xs
Y8/nsCnmKY964mVnvmtVs/lI737O6oT3ZzGDqVLUHhe/hPIR6D17G38ZMvQW
980eHodNqF3oNqrztBfcqTD5sPf73qps35jm4hUEgwOMF8p6cyshuUl+0jDq
h7Z4RxGiE9EyWQUTqn0udRhowD8QKG0YnOlFf7rJKflXRhohkkqjsXAR+k+a
TV1j8akbEl9i36f8gGOaE/+iXHWiJ+GsHdwDusWkf+E54Uh0vL2aC8yD6PGA
RVOSgLXTeoFgH8enDAJUzJy5yhmG0teWPqnCnEXF6rnFoXoJfuyoPQNm4z81
j2vvZ0QwlmDu6BqqG4bEl6UyWYADYaqKoynxX5vf+YnokGWGQ89C6P+Kh5c2
imaIQKthNu3mPCmx6g1bPQ92ZH0WX51ebeWD/4Bcew2HoCgJXo8P3Nt/8IDw
0gAHpqfli5bs8saGkEly2JfEkEceRcZ53RTD7rc7jbRq0KiAzm+Vh3Cm2jvG
QmD4IG9CUzdgR9lOgAd4kxLRYRZrtCKzihGxZq9+wlMGn4R2D9D91USBRtCA
wQtFTd65lqy7TaGyM3Na10t429N0FU5xavpXQ+pTe6JjvUtcSR61UFzXT7Pe
9HfFhG9HmN6ah8reeJIcL/0TiWM+DYdeX+PWxPBKJc1XqM1UMAncL5L8zN7D
j9nO1Gw6VPhLuhwuTDW+T/Heb11kNMhjpD648ncsOSRewOcNDMNabPyUQ8mH
1PpAtMj2wG3+reT6emu1/UJ2CP4p2sQ3/G2mK4zwCucEf347NUEFw3FDUz7C
SW+HMcvvrL1nWZJJaAeu0cAwGjIx1thUKx2j2GUxsXbZSV5ly68n1/vwXEZ/
4Cb6WHVuRxxz0R3bUsbYNgjAmQVOU+feNItVAOhsf8Wxf/47m8NJjj4jFDDd
BIJWoGdjtK4ebgCYQslhwuVpbgVYyBA5WVlb5s4U1/fu29QbOagDJQT4BzV+
PppAVSxDkSNCQmjgVehom8lNAW9LkJU73Le3JcZtbGb6oaD5ukY1YMHwlZgA
KLEJxssSyEuNVCbP/HscjrrpC51rd6QrsO6KiLf5oyI4Kl5haXzzXX9n68WW
MvzjE27bst5KUcQfMJks9Y3UhGN2wJ3kzVgjeJ0efe3ptAfy973NWTdydSJ1
q5OIlY77MwlPhYtNTzHAjmPb5oZGPrbWRbzX/TjT1dzv7tlUL+NvdwJaOnRa
qlrH93sJMula3S73qkQfCtuPPq02jhVsLpThAig7zGfxsDuNdaxcY8wj+tcC
Omej38Z6TmbRhRmmgn1xmCyQZn6iqQQ4/RQTBT6gV0gUc29picqdwofOw96N
sSv80Tawci6sbWRUer9XZwfYdrnSXAPgDTGR2UX30SwzUOEAq2nrevUl+7EI
V5qKbU02w2i+PYn8FChWACoNrnu1Q7/Kn34N7o03+cIWNBXJyVMqVu+ehdgM
HBbx2z41XNWuQaPcxXpgKvBx3Dkawnnk5VnrNAH4eE8B7/zlsZ/sDj92/qOx
vOwZ2kOJ7503QhKaf0lRkmaNknU1JCK1/HgoBuAB0Lkj6GDQq8nW9cE44hJD
WFnzkt2q5+VQo7+rBrijDVPS3iPS4vrY1alc2YgbK2EPNWspfD0lK0zhTYsh
OCSPPD9rUga81qneEHvVudtdm2gM2Gag6nB7qvQ/lc4BtI1DAGSTk7zEyp53
JEoCrBTD03OqYa1GaC9uvSd+TKp8T2V30wVUb22+I4rpMPcYXU5mpMsMfbu5
ZCvaSpWrF1Mp6qyHtWEXp1HKU0/RHgy5c+rtXvwxBzcaXS10/8Bif0fnggJD
iSCsOIXEfDIlVm+MGPFQq8cEDHYE2+o4qxtn5WKySYA1WZTCdvgPvT2Ne+br
kXtQWjh3KpoivxEOZgU6QHhOPZIhPVTWKH3AC10I8BVOEtoU2GfQ02w8W4m7
eebCdzEBO1wrgmQVdzcrDw9GimyOKVO2YgPca8VUwjWZ1PvskYqNB0d90DEC
KHcl0AExeDP0TbqpouzYpBP2G9AAPXNQVPAGKzxvHm0AnCyg58EN+UGnm7VX
qmgNoDUY4h45Com900XHfX5A4cnQw2TA/M4Djx4v8+KzUSJZxnpTjslapZ18
V9LhkUJwCY7b6UZ/j273P4vTtNL+7trAgKx58bMUZUsE046F8MASk/QxwwVz
Bg+NQ1DZBkZeGL98joiu6GsXKXFyFx4RuGDDoLzEl6EyjbE5AwMBl+Rh9Cn8
rSYQXoSGFvTFPdw6RTWqmUxjLo7kEpqmk1Y8BnC25u01UKlUw04rfI4lpvKB
0BDgy9n1iFrQ76JOA6AdlK7sCo0xYuhSEXa+B772A/juefqBqAO11umo3m34
iDbnfP1PKn8GL9E1P88r91sj5TnoWLIftNGldo1glzL2IBM3pmbBD/bzlBJR
RpZ1MG8BcIGL1hv86ZXbQt3LUjubCU0H7Y1ziopeZfz5n5/QbpTW3GlT2Ak6
UWBtGNTE/JWMlt+hhGWgNHeGOpCGhLYKTBshXdN2visVnA3c+CtLSZM2GzzZ
SMV+qDE5wRidmTZ989nyCGYhtjh3Q8EU3a9ysIJ283JDgGcao6XTeu6+weCI
/s6i1u1dg+nyVy+TR3sH8rSADin5MSjmBc9QgDVrKEB/UTHlyH/1gJCE1Y9E
AEdQN9mZb/m3QVM5oUGwIjcwEy4LWjCdGgu7KguhbVhIMyR/vVkuZ/xo8LCQ
jJJeNTr90e+F8GFHUCilrbtuSnCfmWpLIUqRk8RZBIoFYcMj/xHuFSX/2Xnc
hRyFpnBKE/udRDgyJTjnk/ZOO/v3lbr250Y7sNDIcaLTXBt80Q/uweWXYr9d
Jp1zxsODkOi8w8OFM8m42f/X2WK43X3KvBzaOavDwkDWB6zOi6fTDvu2R5tb
Ipr9BTIr8gPvxAoglLzo79Iu4SG2LgQtUCm7OdNRgP1mFlrq4bdRj6RCm8Qd
iU1qp9NfZtZqj50Ew2HayBpXCn054SPSJIGMnUqH7MUXqM+hhV2tGPDz3ewc
LMKtKVA5fSWAb8u0a898sTkcCpWG4A2WQxpDrjfHpv+/pvE8KHz418CEM2Wn
FYqGMgPDMltw60Idl8F6ijQMxlKFfJc+9zniCgX2mE7HuHRTmhSsn9OCf9ok
j3bgRXVpPEMH7VhEMVis/CF/yYttYCGjZtsVVkCM+CaOSCWFTMLfnZxI6aXq
Oz4x50115FZ7RFnJ1oPu3cWqIUMcNThE382SMb68MO+idWSt/G4kWiIavQsJ
/gSJtC8CsOjuwt5d1QkhUS/HDe0d5g5ZkUb1zo/EA//bWvk0zpu+SHxYgOPu
ZszlbNYIDX+ExFYMtI/CU1iMhHWPKy/C5+wfgxSI61KBLebkTMF7rFZeDlA5
ZMVLuaao42S/yOn7+IOeEGpSBgipln86ai1Uqdowni16Bf/43/ZM1EZEgt/6
MtUpogh/eQrTP61I4lJH25VHDlEq+By810AuS9GWPyeUnhyiOpTt1g3ik8l4
yLBZOcWh6kSm4jv/3i5azcdvrrcbtLajXFZbvQxqayohl2kUpQ8sEThbPHl3
VkACmjZoLSpO8f3V/bApMXDbQsjp3JQak9Yvatbyiluni19sgIhnUmz3J07Y
o2Ig4lIcgxqwlUW86aG6pgkJ6p5USx+s1xf9bD78aKMFp/7Yc+wEb5+RRjT8
y+n2x2D6sCd9eTGlgpYL9zacxVIZoGAnNe/oiypXvEsAPIQEiBcDpfILS/Oo
qRz7OEZsFIzJSu1cOlnGhNz0pvDZYcdgGG/Ho5rySIlspnsyBnkAdzwQFKCD
tr94pSEGEGGwMoxex4NvnowupTf8ob3zXcDBiAaIEsHFEykAJmug4HM+PgUx
C4WfgQNN05eFAReh7x9FP+UszeMNBfVSmKF9exDMRT7NtQgatKkORn9sv7ie
rB5mbQTOqhZcyhkQAD1EJvf1g1WePa+Gyw92lnS8jRW9Vl6M0KSH61nES7R3
0BXUTaG9JTWxkmlJ3s1uelu9H/6Oa412nujJiyrNCmmrd3FqhN880ibxFa3N
RRtYlccVo+ISHDUyz6gkO2/nyhsRUX37FbctSLuAGQWQJOR8jU9DDo+LRmMA
eLFdR5ErLVSuo6QIMMcYz34V9HaxK8OOrp1wcC3ukuEFTdBqGo5SNW6eE0Tb
T4HpVBHspwoJbMY2AiGDvvnulk92mP5btPqE5FWOnbSo4HLsgaNCzEqqLXws
d9u++/OBGEWSXnWATfZELRODs6X2KU1HhoQqWtl0IY9R7dBHDLp/B+/R1WvI
DguF6n4tqSjXfOfw8e9zmBew0hGMgGVbYr7LhQ9Bd9T8+AgTatiY+y42OT5u
4dnLkhPdQKAipLVF1wu5GpNBHpUfXYZDDXdrgQJCDr6adkzkQEWFB8zIhd66
r+qLESJsrqjCxIG76+bZlUPtexoP4OR8dUVBsYvFrUbHx7De1W8mex7fmQii
+W6NVpZpnbt2PpHd3DM+/BQcnjHpjPvKt6PDVoM07fojceC3zysvQtWU3sSW
A3jV0Wdl5YhPSz+yAuBQtXPR6uSLObbOnnxnQU6wWy4GNGWmJtWrMQhH733D
sP+4clTbZYCsBqAWEop1d9141MVhavI4g92ENLNnvP6UCCoXt2mfTDX5q99X
Jhjb6c0leHlUsDytrIeGQTM87BAuJjbWlJRmY6EQlnQLz1FIfLwHU+vcTbp/
GuIxHlBmXkZyTfz/QYrVs3FrOpKE4IyKNYzNhRIuZY4CBBdxk20y9H5zgOhb
2OK3FoaC2SAennUxeuNENvarmKhOZmmyH+b9wMQctFJpIOyn81QhCiz6/cv9
dUJ5s2J44PfL4vw1x+99ekWNUY86w3OZypy0Yank0UoJM/pbMPN6dXhhHNvq
+WMXVCIRAsrWL8N0/Ljn/sP7tC2U02v9/5S+ZHD+E/mysHyZ5nKjFtLnCOJC
hknlw6vgtOMZwM7WySx8srOmSQqse54TAyRAJkfOR9SltOBsaWEADUVALgxQ
llQ+hmLBMOOoDkWi9rvNeYzO/BTpE6B/TgVrQthLl32H/XgNTAj3j+FIiu8Y
KVlBBGIcryRkcs6kFM45SgZoOpSLuJDJL6SikuK1mBUXQ6JXPRk6oGin404e
Bk8s8EEhFtaGVfsEAXFn0nARalOQ7wqnAPNvriFD/RG1IDR4oEPIr7hhTWOE
IdZmhID+Aa9OUA3iJTBA1GZAc4EbFBIkgr8Ilii8Z9KLS0+ke3sH9xRDX64l
kYOpOsn0xy21mw0dK1/XCk2OsekLvEc00oi6z5wOoa2OBba+y+PZzKPCwSn0
oqPHW2YZVriV2Vbuq8/cDF1TvBv2O/uyuYkwI9i+m/ra+OI+LIa77LL85BCL
Z+9fXxhM1Fcuk66wmTO91xcXGAJ9/XSaNjZi7HFXe8OlE6ERRUS2JGbd3kpc
KzuEb4yABemb9ZKoZlfKkJ4TYSb4Z+XhZQwlYPu002XlwyHmi1tpWO4vOeQd
BgYYeOWd1+LnXwPfAdpjzboUzuyUjX1mCpWI7B2BtGbH5KlKYCJBHWCTDdFG
jxPUWBLiKKuff6YI6f8boVrfULYFn59yFp8dDoHU5u2E2Sa66zLMV9nC6fhI
l4z2Gc7hWYPUPihlKO+2UUXGC2mv1QkmAkY6TTfhfdwf0KVS5TWfAC+uYnuW
Df18nbhV42O3eLe096I3Xfb4WB21L6TdJIXhrtQ1fqynEaKFuU0YGkCl+IHJ
GUQiGcAox8m9S6Z6txEYUreS0HGu1W92gCe59KXx17u33ueTThC/AnnxiAwd
odYF6RM8nSjbNhOYZ0+AA+ndJk445j6rL0XSs7K1fdfx5aZZR93Ie0uFuVw3
DolFdNn5tzClH1ZqtC4NdgJjWqREvz//2HjDVdYF2P/HgNuuJZKBtKjpeudO
lcm1+kqujVBxckjY0RwIov4U3IRskWxHegayQxbBMgYWvdkyMcpSZgoqiDZC
iKbQIjb+KazkBcn+zZCVtMtzP2s9jWg6pQhM97rdc2wNIZ/5npH18xiSIhyx
r23bkga6fd4IO/aInTe+EEMHDmy204TcVfmih5AvdrwfL1bginoo4jxY01YC
THKBaTYoYZ1c3kgZbH+1QhqEjtrEgHM880kBrHxDzVR+Bfv2qlB0UedO3VCv
mU/Y1B4Vnm97a+ymtHr7fAiABbm2ITDq5MrOYiUqii6F3CwwQJqhCx5eUbfC
8Mwk89+IrSwa+jvyRxmY2X3wBDFxr+F3FUraWIKvJMxIOtpId49UtqmgFkJr
yBB+mIjv9K8kqWVHn7wpupCRYgZGJquOyhOleg7FYI2NdyRYnEhS5ZKnO9Yd
lIDnvNqsNJFUbNxLOPawFXzBsVXuR02d5TlvI0t1t8MGF63uV9wt4S5KE388
ruoUtmGRMF4u8c8TGzjLPUNH5B+YSS0z0XZYV4tMODTfNAqSSLKS1F2puGxK
JibQo2OQwI1nJ6+nMrBS1rs6fv0PwU9b3UPjaoT9Ri3kdnTgZGAZcE+oAcBH
DDmaLcYHXwU/zeqBqIZpR/UMhEg0mdjmCrHZXi65yfYGshV/KKd1xomQaC6C
52VN9vGaakHrTDxEVKHb3w2SkhMgZss+woNf5DYAuozZgWOwjNme751GCL/8
9L8ba8YIdRUbV3oIzKrfaUk/BoZzw5RnNTc2ttAG6E6G+zYTKsy8Nny4yix9
0kK/N3LBH1Xujb/uRzjuU647SaqLFysLtetHA06aUzL1QdEFF6yAmLl/d35e
dEfCfdLYnkDbv+W1ICyUcdRB+xD66eETt0+lJnr13BJFXv2ttVMZOv7j9eBL
tlkTORrC05GGwbXVSIAMbm5Whkywm8/aXvzUt0bb0C2DLLQswNVm4lBYZCpT
v75q7vO42NWIQivUasrldNerfW5YuAGKh/YNWkWRpOFwJ0ZjFE1ORpY74no4
UklTeaJ/KJuIJe5XDchzrJBdW3AkHeFkhg77sml72vjZzNeJbIgtnX0QsGGf
7lUfM7Rw3MomzveuDdWm4stthUX/YuVv7IvcSB0xsvgVH2fj/Pa2EWRyySfN
7mxNAhh0Rvp2YuH2lGbAhm8lfGWNBmJ9C5L1pf/+KozAgW3IsVoI32ZNNJaH
qeedEd7aowerEweKhwFEx1YNpsuqlRS9hdBxsBffkV5w11szlfJJQj8+vIf3
bGPXYYnczsdPbmshw4ewDj1i9nJlVHtsfQ1/drORhyFne2NL+mT9nFAMAN+J
NjhpFF1C4Vf4w0qWpYSqBnu0oxrwRsIqyELPaiyksf3LD3EGjvxJIJwWFYVJ
Gb/O5cFgajTYeN51cXDnMZz3lQljhuS0TYibs4Zp3fDugAbeyBVfRuxdRueQ
w9PZRT+4bmcT/UG7kQ0x/DcHI1CA6AC3ny29EJzjOzP74MkKglEHBYMac6H9
gomSBVp2My1pDOxfcJh8bfvGgbRmiyL84ZY33a2QD9UVLTGV+AQ7EArXixCQ
1d5Tbiqfn+lDXgZdlojXES/a6k34gTJgHRIxw8NqPgDf299ckOLiTtvAeZ63
OTXhdT6jKLsOannGQaxCDsOQV7yeN3KS26geR2qb58uXqAZ/xZuFWj5Mk5j7
8oErLB9Ah6AdRPslGFjKHr+dfU4p1xLuk5qHmEmaIX70xtkz1PY1H4TAbtV+
9JHxwABCpLfmVlKfTKUPh717pefBoFJCArpojfgVUMeJvUVIggVVQY0m1OGH
gAlzJah3X7DeMw3zUTfCB7S2cYEQfCZqw+Rhf7SDLFeuOhK7BNyIdD0LPCzp
GyUr73TukvL1uqLJ+a1uTJexqG06tTdjzHk0VP3FvGRMr9ucMsyiC6KXOvCS
AyKjz4a1p6CInQt/gwAt0tVBr+q6jZvuIJJC/mZ/+PWzsbx2c8tt4osBj3pf
hfSbDoOVPsxp9YYQ4eSpNlbuL01a2Xd8Viazm7QlGTlnRJnGWLhHJVtqyjv/
gwaBXivJ5CBpdtYgkonaVYbYgUcQY/MfpPwcX1p955HCrCTd2TqYrHNe9FiG
LpTH7hEaGe+Ab3JI/YTw9w08c9jEIZNFxrPU4FWX/4c865pZmhiSJ6yY3jTW
AqzUeqBZ2/e/aTZwUY5Kk7xTwTZioz7cJSDqDq2s5HU/GY5aycc5EpLmPSEg
k3Dd927SdRt03Gwtgkvt54eIMA2gde+JYJSfB0P3YkLHF34qJI8/Zm+ibOjx
Q/t4rwbFZYEdbpTWS5+t5Q3qDk+NZQ38+W/qdqAL5g/ckJ9ELsP+QCk0abwj
XLme+SfDTAO96p70d/pJRzn8zsX3u/sc99ldL9MQ90zPqIwCWbUA+8jlgl6z
76+bD2V3GDFSyh/TPY8cVt33iu2HC0FGyim5PQqArfG5W0fze23sRLAps+AZ
lYV/PJiDKYiPas6YwpmPaUXHqdIZ4gl98ujzUR++zAUqypTGq4MVnzSq92pE
WyGhG/q6lj6FVXhsR0e+g6BLHsPq+RwPaEIl5y8Rd19tY0KM+n3c0GtnbezL
9kp+pISy2C67dDdSYKCoDnyJdFE7279j9Qf6UQalYoWsFLYRx/1Bqj+1B05v
ouQZRJZM1yLGkuTHfV04qigrLLhDhDxQV8lzPCzsSeeFcgWOu5uSKYrTKEoQ
2fyjAUzQXHYLhs4ULZc2ISDq+b5Ux6k6nSMX/yjjImMJrwEJXjuI4LCsXane
fZoHiapNPwcU8VCWa5m8dpYC0e8ggWAlMG4G84bOIJSn9zeMQ0k3aTvsup+8
et36IZOtMKsU00OYGAZZ18sO/TJtrUEDxZOTyvS8AWs3WcyENEGZgNX5dZFa
cUAJ3Jtyy5W4Dx6+1mX6O5NTqSTTk4eKb63DFPpN/fL63afRGLZWvRIXNdZ0
VVQ/53QXsb0RpnJ/qNx88pml1y3sJt+eRw3A7qTBBsovXmQISuF/w7eTxrVL
+Icjfu6nOyGjpD+IfRLPEj9VQcDwUkhLV4aWC1pV3Zgww5KWAGnQmJvfbk21
N+2Q1qTKo1HK+pAQ5tYzxQ033W36vQB54KAAcLPZEUYcnmKI1Ks5eFij74Uf
oeem/7H2YOZV0whnxahEAGkDcvlS8WZqzbqgw3dyJfhoFmw7gnwEIanAKJm1
c/tx6Ph0E87B4YGJlt6doyGtHwJk96gX3aurnXK1YD6YMyaikUck9Wp/x3zR
8bBjXiMb1r19ryE5izMJTrfX/hnT9jymNcTgCun3HxBmzpIEVqwerigxhiMJ
rf8DxzmP5yO4PmN9K/EvY/54AO8CfEAL4I1yOJatfFhoagQZ/KvishVKFG27
jfljqFXKQBbj8YkknN+dal+nQE7xedrg55/K8ij6Nlx6HQ3lHi3R8SME+Fwi
6BT1oLLsy4pxpzTtMMACXgcVFYORpEGzuWQsbAwyYBeeDPvcEUP4BSiq1864
dBW3CjVtkYKHEWd4IdafociOBrUIBlXsVoI6ArdVIghtUM/8OMch4s1p9HRn
yqiAxs5fdiF2hxtBn4B4zDIiSXhck9KJ/Kb6mEOW4/jqGQFOu0pJxm/FCN6P
is0E1maR1qSh3mB2tmAOfRjqj+YH1Z6u1S5l+NlkG1O7E+UtQzADl78igPmc
hEvGUh0760g32ifH1oG8f4h7G+5JUx0SMorHKFYOXQblI5viimRW4Z/Z1H3F
26r2LABnepzqaY0HYCOV8qn3sX998JwRKSjeltRMaVWBsySdEQBZnWc8BVnd
aESjqCBXz4CdB/cjab7Mceh8654qpWi+Xzn1m/X98V1cuCc+ijOg7fuBhdVR
lyGdkrmWGTio8IoRvmqIugG+RE5VcTU3uZj2Gy1a16HsWQgE06fZ8klkOEH/
0Dl0E79t1LfHhaye9r9adopm1quihfpPzOwGPFPNic5tndCj3Ujz/U7pIf7T
MdNqYVjr06Z1utq/EJ28S0H4BV/UTRvyzSXaoiy4j9JDtWpfMLeU5Geq78q7
QCHBER4rfS8+6HLuOq5kDrU/ZaNVn+YllgmM3PPNHSfm0U1vzGytWpU16UL3
wynrTHLkX1nWntcSz43cAIQzJ0X+Sa/GqGvBqaahAIGmZbyjFfCMRXPcqr0g
ZipOsF3jIGQ5xZrAW6rOHGL53+ywFhheEUjXLPzZH2GIUYRv/1a62RKS/0Lu
0w+JG5tBoeA72ThrHFLfs+HXPby9In9ofFIwYqpJkQiAqKYGUoRzNAA1PyOi
6thVFlKXQih9Gc24YFegRXe+3OJ0Io24EE5p4yxElCx2oAQuV5g4sostVy81
cJt1uH5vcIxA9b8VJXO0Wk3p7Wn3NMFmr8CBttoARllwvO8kQwi/68cJ4JcM
lPO7wkQXeqQWcXO8U71SN1/r+zHTsxyj4ijwiZfIziCnJyX6Ns61+R+Xbysw
T5ZKNcyahbgGoqhGmVsrJLFH9cBTtTvWLW8NBHiKXucyWoP6m3Z+ltOaoQ40
GhmMrdmiqYDWATV2/p2UIf14nVui7mJ/zpyO4xApLJJL7pP9KTabNH8chTbc
KyfGdpJ54u1yvYOz/gmLO1Cd/FStd+9Wt/pH33sqH4WPF8rKqUNM47gzFSm9
UV67+ds0qLEbiTmloLRU+3cJ+MH6zFPgLaxFfjIIbr80pIl/DpfpL9ClCSDY
vAxosQeXiVZPJJt7woNEIDy43f2jOGy4fwYGlmnEHMdUdyld26dYR9wqoUTM
6KsWG5LXrFV1hR610aQSR7Dlxbj7sR/w4TjJo+gkD0IaROraoy6/bscSdAtM
LxTs4wG5NuDAF2W8+5kQZ/qAaHVOoTvgTy97bsBa2hg3q4LAjf3A2s6fp6sL
9o12uyhcFeeNkSfQLFotMNAbKiu5OxzMAyK2n69+O0YfxOM7zfwQtPKpHqks
tAed3wT+YwA1VnXx4jwlaYxvWwxs76CaFGzHaaCZEI3oZckTF7j+k7blp2xF
YBq6EBfyzDn7wp+YoxRY9a2wZjliegRiO6SauK9FW1S6qL0FSB47a0opeFin
9Y7jBIy4OwYJogZAtfIPuTXwlzGuZNZYFQfAsZm6O1mE1JZltYuzXN2VUns2
rUGvmO7m6hR+Chr2YzYwe2Yn9mn6u7DoC0gqbgwHPdQ5Tx2oVykhYfS1LflR
chSvMtfUp9t28goqqre0sZZ9tYA1lgy0cI8ztTsGGJMGRDthPd/VoRuQd48G
bgUKoTPVnqWHybjkLRoEZ33RPr6TDWf1R5Os9mQjM21ZHXm1BEkGjzK3OAo6
vVE8O3UiVJzPy5tjdTeQeeXyFGaquI35rbyw5dbIu0PhDsLkhi8QLemRA8Ot
lAemnUDvo+oQGWkgtuxe6p+g00taNihMdWXrO5JP3WX23tCSSmxRL1jHEGeB
kwCLqGTOTrCU00ALrdTeyw0qatMwMps0URFDa28Z6mB8r1O0EarvuPbY744s
nHWAkJPsqUzDYR2W0fAR4feG4n0SHIQSZPBOniB8ttzkdEBr12XzBYvxFYaR
TdNcKqtbweBa+nNqj740qxY0BbZETiEPihKr8hDYZuFIsgNluOpG4wdh6rHD
zQftk4GEnWPRSJWyPATrgCVxTSGzJMhWhWSObHmY6H2k/qF1tWTCe9ofU6Ph
QVsUKbll+zpd+i8Tx06Kp8gLGx+Ztq3+cRlejmlyp2JG6qXV5Ks3QMENA3lM
qWuitOwVlSb9oR4fzbwIeaiYjMIZaL0JTRBQkzqFjIfLQ8rDI9HJrcRNY4ue
SDVBlNlEmbfqLKL53tv4AIIJxtcQZdI6Ml8GHgorqJaYhkx3Lkwz+4RPZwUx
eKxUndPgFLiFQZHEqj+GaRAqzu+P1rVAG2PF4BkDWILcWKUUrxdfaRQWsAkU
GjCQC9rkgo15fMzsn500pZ/7IvJETyqc/rVIZbGH1i4xahtvYLnwWvzmUZiT
K2xrUDQwAIvSqB7IBzSCrW1WkELXB1kg9MCunGj+e4svsxnXIMgQu4vEj19D
jJVM9T/NmITNbZ+o0x73uZHKx+QMzp5/J+LSXeGzcq2d3jP6Qh0eab/z1XUN
3dnMqHUtMBu9YpyiJBUQqH2VA+7TMYXTOeimLx1Y10LV7dKZ74Lfo0FIcMAG
XAblYtA0j9QR9MFVSeRZOSGHJ4+wcC2IzKiG7a5PQ26vywPNUDnFpio1VPQX
6ZaL6+t9KFkrvXXDXss2nYO6GxeH0UkYkd++2nCIDnifsRXKbFN7n1JXIzpg
HHraaD4g+3OefGoO8Jg+n4anl3kwbEhV0GupKtI8s3WjIJNHF9Bs641NEQLL
kbyt9mW80eMCgMiChgjOXbUSL/7vMImR8MlOwDbaQL2N/8N85VT8OTG8UYFL
1hwDf/Ja4A03PPs2EMUjDxIGkE74wPnpmGogJaI2T6HhKQYyz7rvAi3hGNbP
pbBWotJEEcyNiode1/dUL/D8449p0CyhLjbtWVe8C7CjuFL6On1NLSG2JDPr
k6RFCIa8MiT8ptDAkGu/m1rd5xlwVQYSam0gDkX/UN6A740Jw6aVb3x1Uz/V
LxPSFTrPLhGiDePIj5jOv5ZzNe5PuJXVvoE27XmIggxYKG2a9aXzoFFTcgVA
RE3A6OuD39g2rkTAQjioYQUMjRRseRBDylfeL0DpBbEANH/8Zue06oeeu134
iXgx2appd+lUp9fo2LO2u+Ipl6mesexS8x/WZ5oXWPiz0TQKqfxlbZWLqPjl
P4mUkVL5q7P6fOlP0kwPEo64e804JpaovMpudSsTdY4hrWZp0MuAMqs3+IVu
SblWv5mFGLVdR71kpoc/YSN9hG4sHtkxIR6fSq38CLpiHnGpMESl7BiixLYL
A4Z08CynQItrwSh0IkW8I/DhQR22E63dT7cgkLMNrf2DPSf3OIW8LfBiPBpu
IuAR915m+e+ZryQMZG7BwWMdr0sadpOQICTau05a6dvcnZGd6xcJoyu68glb
9hNxN7xFS4eVSQhBLtAr6GZ/cCZnUNMdXsBcZ381Xfug5al3K1GBjcVJwWN0
Hi4pNq+d7ZuENKuejujB9TZUeCffuvLJZPYv/t3YdBobiplCo02QRbWRa660
81eOMvsJhPRDcAJfDCkRG/uvIG/t7rmDaXcwjj5O9vVKmwVI8mfGndmMLQfV
Z2lFpINvwmHfoDwA2LUud9HhBiRaHGsfVjGaO1xcXfJGwBtw0savq8K9/qxm
2Z0XXMRvhKRWegcGUJ7Lib/1ZRTQrpk0VplY5p2GuwwtY84452bG9iKPyANd
d2bOkvXy6uyy8cAi6rsnm5oQPOF6VeKW6qunSh4IUZSTvkh0LzlT9hEH0TXN
BZva7uLBzYjPUasjJIk2S71hnyxJCSsFuNpw4VVFIggpA9vSnHRG6kHG28oi
a+4af3fZOIAlQO/vE7BlM0eHxlHFL6DZ00sWONcOWJq4i9bahHhMwtbvaznw
a1OQQ+1jPvtwajtPFyg5tPhva2sczQ8BeolLHqlLqvbQCCADRfCnoh0PxmOY
K+6nB9aGcmbqMpORG/KJlxeUHHwrKThEO/GjI04CtR4FcD5k1H8++/bDfEae
sWedcrZKKowPX/AeeYvaVKAKxr4HUcHU1iCvr+wPmMfc+k60hN0F/p8kUJ0T
eHxWexJd7nzAf+x0KXeBH2ptSXRoyxqnj9yNLyw5P8n4MTCUi1Rvwr0e4fH+
+3GmX264fxClUBmd1xsUxdqMfxXmyJ3GFvHgKcjAkM7k58/NCAZfThlEdFNz
Vmn7d0p8OhxAa1yoehtooo8vqis2CG/nV3P1bkZeVLP784U4ROcCSNn1lPqj
ILo8GtzoybU1/ADOB05BzEZpaBGd2/xS9dt6PwnWvUt1pmGrzr/1qQJAessk
+1SbLMkw9bgOY/V5+uNpktoGine7pfMeoE3s1hRTTBg5FVbhsXBTh3R3/8IU
KYNx+SDc21bdsQ31ogpnkrCc7Zn9r1wDTVettuo01KnMmMBvxuLmFlJtN7Z8
BqWecuapcL/5V5K9tlRpioyciT0syTe7WoidqX3RA1B8RefgjbMp2tHIIe8d
4x3EBtMmpB0abF5Zz2ZONJDpjxl31q0P1BFAO0TBUSwyKFiSMkYs5I+8XMju
2wBUCF6mqZvdIOniMH7f0XML5y5P0gRjeR/WiO4DkZZvavqsyIhgE5w3Ee3B
Mf8eXIkaaS8AMmj68gYe2hQN5FGX5E6pQfoIYWg9x/uNw55+mMKLfZ6EXgUR
Sv123KRsutElNLEzhuf8g+byJvUNnTgPhUk4t3Y9H0gFJXYkN6n4MAgyKkt0
BsL+kzSyRcMG9oPqMYUSnxux05ILCGkvzZfk9q7ZoGuZgxjsvbzs0++Jp3rX
fBqaw5dv0IFglnHuyeSCGz1/vG8hKfx84swwDGxf1yKPS1weOUWcCukWKgTp
kFqRgHIYUlbuvKchl7wY02K5OfN3nLKad+nNEfatas6xNZHAQUk5oAMV9T4m
FoEVPTMP0cHKkIcKeruJGkP8A/J1LKnU4rx9OApXtJ3qMYAmGdoUVEYMhL5X
b5SiuTXySGGFRfwBEnNjYvcdolHynX01dP6FOGhOI6RiR4+dpGO16eLhMC37
YUXl+dZ+cMDdY1I+3clO/N1pRLYA1gYw/jox62GAK+ZX6ul36zEo5FFam2a8
67bOFZBNITOzoLkZN8G0nvYKUnzF83uUtj6UYlQOIdmuJLTGLwTh3II0P/QD
jxOTihfCLWUgyApo/fQlhYDBLIPHeTXAfGtyAJ/HLhJPDtOG3dVcnFJER31M
g1XryXDLI1WvV2DxK0COid0l+rGjR5qL7BmQ5r3fB6fXLwdiI/WmJ14IwH/4
vOaR326XhPrkFA052T54MEd94fwM2FHCp+hOCw/djKEOsdRseiDrSctaIc4x
W2VSzGfsduuo2BGTnDNdHjttNXsBDA0wBY3ycyXqzZPlthYd4KiwCxuc6hHN
ABNWqzamlItHo1aAuifeIDTmFM0s1343H74ojbZBDbN7zxm+DtmlTSmAPI7q
7l8rdmrNajcKpU7Xt4XcKjWlqaAUPtRF9hBwMTp11BKO/VD6qpkGVWe0bIIv
nrpdbBEQZge+d7NO9ogInBS79xVDs83xBSBHQl/pwcuP5Grmnd1lgOJdAMmP
7DLQvvtRApYUO1XNS5NubSd7Us70oB3j5qJAyKKBv37dkxIobtvjkYU4k0U9
60At4om+mRB3VSp5OhIEvqCAGGFqgCaGXkVMD4Hh+SYvE+nNjEbDiHCt8Zbc
kcKI9Vt4AKCzNae7S0MHU7cfnOfcYYacAOxqMTJlyOe8Ix+WEq3rxRydl4EU
iSDna1+PIxTRuKS39KyhidthZgmv5b2rO86qtFMHdQCUo18oBJnxaduqcAts
mof8CuNrfkDOSRZapLuEYJ0V/qtFphJt47+89EZf0B+AqsEjdus3q5BNzlQj
/v2j8slaB2D8g43vYZStVya4cL5Rq4sL8A7HJAHhowOF1PsuhuAYwcYzz/Dt
P3SIZ4k6WkT60hCd5TL5Ng1bdhd3lfqKxfgvtsywNT38qkPTlcbiDwreslYT
gimbbA7EO5cEiZPwB6OlvlCbWlyfteOJN5JtbJ6SkB4jeVoMkbhtpH9lnHEa
i5jIWRmCHoTwN2xJp1qV2Oux3a6zZSUmCkN0zpXfNyfXtiyPhlHI6sIscTdP
KMJSEp3D36Mh2ID61SqKSz13bZr7UJqv+VLqEW9KN7vW5gln1vggesi5NHfy
16u722YFD87nLsoZP5tlrAhJLx3CspJYD1Xzt9jD/naG0R0hMrMZKcM8KATc
pb/RVi3uxQD9F79eetVYxAU/FldXTub2dr3gP5QG23nmOsYoG2l9AV3LNLMD
4yQHw/84XyvXOARcqlso7rdHNs7GbJRWzPOrP/hsnxmART4Mc2RpCMr1g5Yz
DH/KThSwCS4euBduYUhL28sQW7zcE0EvYZeOY5hnTOZm6JHk5t3gPOmO3j5J
PZ5oT2V+KE+bKFNcwohqNJASz6jIpCyXStkPiGZwl8DsgXW0pfIuu55KnHOf
lHGMYY5U2hiNratY/dNS/KoTkrv0U5c1dYB3CqBwHjwpQxx32B0gsV7U35jk
fN+NSvQqdVGnvGXxaAuJVL/pltH0SGk3gq18xxXjnmLO8kItNx0HZsx6whrl
JJkeDJuCIW4v4w/b4iFZhMP36MunsrXjYbSeJRRc3L2skiCfWy8k2gzPpKLe
wlvVNWQjbGtXvFVKwT0p/ongFkjJ2xN2lPzFQlkMILVqC+Qy5dIrzjuJbe15
E6JbKvvlh7sB4pkRexQ03eQq46XUTSsJ3wBY0iI4lOKv9EiAZQ0Mj4eNzXdH
JsjKuTHlg1lZLjdyCcZv6fcCM0w0OqLDN6Va1UpeBjKuT8wA9xnazXB0WgVO
5tY+3GvZCTmFgK2y6HrS8tc2T1JNCJlOoLs8+tWjOZi5ugA4dbPyCrvwUngl
L7HtpR8arr8/ufPJkaDtuAxtqoiZ8m5/frnxlLST7LDJSmSM1LZAG1uBFY2M
VxyBdAeTpgIAGvaqALfsp3IMWwTYEL7ZjBLJOJh3F+RvzVJOrhgOFYhFm+mf
SpTKduGty2YrSV4mPoPnwdjtFiHEFsMQlIeXxkrgDrebbBagmVnYFT9hdhUg
vccO3ScU7k4Gj72xQCNDlIh4i9WimQVTTqw3pQ2hmpnW7gyY7hXv4bsprcaK
e0SK3gKOFOgzhoEkE11Z7ip8Y6UXxQ0NcjXmaQybiVaCAYGW5kt9U/G18tnj
jXZeIh2CVHmCgesrDp3cXm0kTRqDiTG9EhP/P8r8hf78tNlONikj+jE1lkYe
oEmVG40cKdU2IY7LVthi8tD8eJUAW+8COOC6JWmTursxMnllwyC/5gEU9n6V
txkKudl/lFbTy39T4fbivcsfiqVE33RGtwHRgxkkMve4omN3ghjXLHtHV9Ai
tK4b2lzX/1h5FFxZr9kS5NDgSKykHWj5fObS2ICSqngUtytT2eE5oECoT5Sv
Xa3EAvfh0yw6jCiivgSP6xtGi+hlUglq+hGq1uRkxlR78wufrcIkHqRCOi2p
8RbTd+bgCLwQlF3zD5BUIEXyhse3wl9kP0xIUWksGdgElI3HEKouvBfhFgyJ
2H6Q3K7QltzaHE9cL3Qhtfgnlwil2vWPTfP+dp4I8sZRnINwLmEq/pjEsCO8
7cmOex56IX9qKllyXqIPeVNWbBrctG7W4Z/l8ZX/qTx2LTKjCFUZ+mOsly6E
vcKibh25gd9g36hKvQtbGDqHulWlT9ZYygx4Bhw1afuCizZg5z++RO+Em2kg
rLSE3nWICGT5+b4ZRuFxJMhi+5g+mp5Xedpn5+aMnIL3r6VMdPBmKcW/oyV4
TwDqnbGW9Fq2qPIijWVikxfeelm73qya4neGVcJ/HIrjxsQ0+382hGnDYpxu
bP3oCvsAiqGhW32WdKHaJ/vqPX5KvgR2sLt1Msmbv31aHa9jRGqF7qMWA043
decZNC7EpTzJRh4O6yxY92soi5OBpuzoDzijzxyrzKzkh8Cw20TIBB2ACo24
OyippwK5/zZPu4H1txkynZjbUz8OmheIuZf0wtz8zihEUQ+BX0nQrhK+iRVd
J0ctDSHmCv0H6PGjZ+9IBWQbeWNb5YlPG8S4cymsIPalBAGAFBVc0QzFXGF0
JQ3ih3bmAS0QOUzqD9ZbMVLsUMaokOyFEsM59G8vp2TGOTeTFTVB7eA+5nQg
+enF9XNavJ0UhsI0Reoh2gDeEHlqIct7H9CyGVmBMqcfGja5BcZmTtjk6Btl
cCz76MgJDnn8Nv/qn4liW2b5vofa5ze/QjUKTZ9jlxRSNFn4DMdrkZhS1jC5
vpXiPG2dA8nZDQGfhcx4vSM8uR6zInIkHEnvlyVD8qkmyQfbG/wLsosRzVDW
pujzoH9Kmi6yC718wmwS1bohM6bSaDuy28fCpWQeWeT90f/IlVoVYXChVs5j
XALD0BJQqbheJD5R9zYrK3I5lLq+375tZve62yyY3m678GIpQaLFgrhAeePd
jFOfDDz9UEjHC+uEiU6/30aLW2OLI2n7iAzBvrFP7NMlpXrlIonT3oD59RK5
x0b9H+zbq3vRw3TTKecUHdtu+JdFDdNRVoQ8WCagqGvapJ8XNZkTcz0EAKxE
kvAl0xCuJAcTbNGuqQHIMwdRbiPEF0LdHYc62M4+jtkY64mEeF+WMwSFB9uI
AX+GEbv/JHE3vDAJ7U+GCN7uUJyIL+aozQWFqBaUDaG6yFnqeWRPL9TXtBGO
/6fXb900UxCxM1au0W+MHmdr281OXWQaTGpjoBxxydBMoNQZzDUV5vS/0KAa
MEcMTdcPjp23waVcJpHtOOLzWzaX++gMSQn2Tj3YmnW92vVnXQOMtaEYwV/p
EIYOWniZmaHGrn8SINMwEtWjYIMEO6SDKIpcvkgEqtk6t3NOu1+ZknrvszEM
ZkYp2jhj7dYSEEu1krshcaLQABftUIRZyhgsX4UOxnbULMGX1RfrSHiw+1V3
35+hz2ovoFEcdaV8jpozf3g8oZ7JVhLyK3N6he8dxULhLkhWNBU+nS1Lep9S
Bd3fdi0XUoDd1AT36+5Hg4z29b4X1fFTnGle6hpF4Pi4lR+nGdFZOHQEdq2F
/XwXvkY6SdLssqhihC8ZtNaLBqtHyDTBWMtYYw8771k/w7jQk9LCtj1X2g1s
XVkmg+YbwVVS4SAt1Lh7jfHiNKF1vpFAfv8rQXmZ0+Hwlo1ZhjN5jyPqhOM5
VJ4OuSdWJZhdHodNKb5K+ZgQmRaopydkESBo9wPCsfR/2yjwUDq6op/DfLRb
iit71lWK5ZeotVTdnmGv9RnsGvL7oYUcdNIqmG6GfP0Eq/GkDy66HOkRKB0I
W0YayEiSlxK5bRv+jXamwh4mfTVZ8NaJZ0J98XE3R7NBl06K78CDV4j+EL3b
pwAfbYTVnEYXsZo91qh5giGyMGj+mUJSpkyQ6Oy9FZ4yEOolKbhixVx/h1Ka
rMbvWccRCm/CPEQ9ej1EkWrGT2OYHBGUXnRt+mpMcX6PQAi1VVoAfdTbNkqC
EhUe6bvTNUQ5M4JQXcVK6Rr1ZPXCIXyRXtCWXRjg8x7Zp3+da3Q2FHy9qdA3
XlpyY/BgiDz90oyoyrDX9yBQI8kpTQO2KWmuwKZ6LXWagcGe3SIRcRbEi9ES
mAop21rzyqbGIn/EGGN7NUqVvpRe0XOaqXfitLDaR7Lj8MoM+AfpFTqUihlB
cug9glSdyJKVcvoPRFzFUHsa4idFTvbyJMwOr1wWs/aH/Z3BnZ7I5JjfxEKP
L0S/AAVBJ0WnyXy4CNsupfgiRF3G4e7KBM7KQ7KixS+nbhk8PorM0F92EDon
F/z2b+FeI7Vjpg1fbB/CD1fWGjVgLi+uUyPRZ+qe85sxI1hsyVVWXf2GQNWE
6XTQL0VWx0nX8/Dzr9H5vb6LBZtLX9ko6APptAR7cPVCLuGFvt+INIZ+XI6L
5CRTgdGC0jpp5CyefQXP/udjpmgfUOjb0mPJpucMRkNS5WbQdW0T8pY9QQmW
EmTS/lP2zY/2fazHno2MbBY33m+sbhKA+9zQGJ6d4uPJYxCagOl3WR5B8leZ
Lxb+AOLHWC6YLtCvjhPaQHqerNYpgLXRTdLO/0vBNU6Q+btJU7xsHj76gllu
v70OuRBb4eXk4hdPHGVpjDg5uPvFyO+35KyXzORDUyjyG8uHs2avMZ7ABQNz
8n+dAfAdHm/C/Xe/GoSrnhBFoY9sgnZ8rvWMh2Zftl3C7vWYL+vyMvx+VfpS
jKwmLE2B95crPDaza+ofyIwQthxcqvZi5GxMAmx8BlzEXHNq3c7lQB2Qjb8A
HL+ERE2p3xZ/hbVEhXRu1RTqka/udz+GWz6QEYSfOvboT/EkfUOzR4OY9qaJ
mBXAVhuX1uGre8eOT5M6BrLfFo99oivPHzl6gEtYBK5TxKzzlOh2fLyBYuzr
TpbPM1NWKiL2fgSYN+1Xfl/z2Pf3s7NaxWcZiYooGdLxIJv6F0GBZlxfCvXm
J1Wneh6yHuzCOCxVgSHpnTBKoLYnBKuCJsBcwhOuHJFJ5jBQmU+7RUjUmHin
wjxonc2wUE+WIXClV00kIXbWxVZrichAAE4kOH6eWgW51avtDeMbqsLR3izi
whZamHXxKsMwwpnX3XvlAKJZB00R+c2PNd3GCk2qk51eWTGGsmVqdEQ0b/zf
9WgOcuKjgZ6Qe7QcxQfVo9DBY/NWEmd7yXQ6xrDytEL3ZikqgCgW5ItI+qpH
1KkUYyaHNk9geGj1jDunD+oqnsBhENUgLJ893YJbP4wMESHIZLCf2demb9B8
pCHdJEDmVqIynwg9O4hyfq2xsINyOcTYOwLeCjbwfHPy9fZaeNE8U1WAVBG4
OghpmNK99hTl4f6rJgZRRVcnGhHc9QDhlJUkhNL3ybVER0wM8etHZwFkOGoX
pMHA6N2QXBXtZJl0q8gQZdtiqDhfSXqwbcZHWRI/86fqH5ETwMshaNHbgDog
QB3wCXpBqBM7Y4qGfVjXulxUapKHdxGvPvG5FACWVkY68V2RqMiB2I45vHCX
4L3mKuVEo01osHm2JbxUKZVQWqHjDyRZRxtJaBmodtG940vLBXbvR/uTI+j8
kZ/U1QfTJwbNoKDWK5vxxpYF6s/RdwOWPoAv4UDxvInjHnNHOb9ZZehi/HAS
bQI5MPFLY3GPAxQf68jW1D1sBQoX2PV0brOLWYnTpMzBxC3VdsmT1otZxADB
kPqX1+r0+oSOeR2tSlex6bHH9FrU0ctLO7b723RlByPFSQqTJJf9qaTU25tF
78k8FUwg8BQc5gA+hpDLOpsptlMa+2WPwhM3en1mLQMzB1M/92sbpn4Y/iYv
4UBjEDQfqVUH0fhNvOrwAPNanHymGzdZSDmlevyKJF+pff70SXUtID7OnQDO
2ugjU64hVG+mBp51RQPk2Wr1DJBKckgoYnZZrq5s/CyoCwCsH2d38cs2meXe
rx09KCNErWN/h/uZKI2rcJtU3jwXXtZGrPiNuIgzNzaO5G7iEnMCvEgpFskD
MBoD8t9kXk6BYiFVE/pAlCdupxiqYEg6L42vXpztJ/a500I5KCgRiExI3fm6
qCcsjTmx6Nd7T6Lmc2gvMRy5ImpydftOQyyKp5IuI+eJ2NW36aC1AjKZXM6u
oWVAEN7jN8U/YJo1BtL38WQr7tWa6DRSxZCCx55GxmZJdcfY/EF8T7Jv4554
acEwm8sorm+Am4Jiszv0Kgh70eBAoge6oK/CVbuBn7GJoyg1tCf9I70HG4P5
V29nAo/Ip129yakqGYyswy5mhcel/iB/XDTNRDqNdAK3QIjtIXxVdNnKPwf3
gXJwVRFWlRO4v1rkWHSYq4l8zX4gZFJmPlVfx0+7XvPY+aT8BKody1vtJUbX
MwlT6A+m3WrXKn3KlUcHGGD5bNQQnqVoP6q/u1lFwiEer+41AgGmyI7ORjJL
0IdYKajujqlKKnM4vkeoymTOEMBwkfOda1dU7s47MQESzlrFjZLiNt9dyOOo
zJVD6riBmv3TlG24ooAX3QHqqHGQqR1x0ru4Kam7v2AX9y1lK+dtD1gTHSx1
vICqSlFpgKm9dwytdd6nYbte2VfWBSioTc981QM3cxMSqFLvULIa+iBSlNeQ
uK22aGIv+cjKWxXufXgV1BNC0nMR4sJ8WCzkSrraga21xQTr7lhteOwTB+YX
G++vRNUhclTrkN55m0mbZR2GPZlagqlYJZB83k0tR9oimphVB0POFAZp1XC1
nHUbv+pkh2Gekrqbntcuj7xXcy9AvncgPYNevlG/X571NxBjp4hcMrFsAKeB
F6IA/gpKIfVwndVlQifLQudHu97JqUExAuylBaajKNlxBw88ZZ4mRvH5G2Uf
GYhg93UxjD+SQI1tQdnmOi+shLpaYZGZj8zrvcLPkxm48wAbryrroaVMg9Vg
eY3AVZAZRUZ7ui5qg6cD34L4VCQs5/vQr81VRaquZZsEHWbMDGS1NEhkfZlB
aG/RTkgImzLBn1tCxoJMlog87DTkdYJBxtmSFrDVsCqJBA/nM+gDlMzxBKjy
QJNiJpYcIFVvecp+j8+gWbJlFvxj+mUYi5G7Mpd32GwMxMNnvHfpE03nwNkK
8H5GQoiE7sPxFVRCK7aou9d7kCRIv1AqPpFXbZQjRiXi5ymTbnAc3Gs1OU46
SGlx4j4M27+aopfvzT4mSNlpx6BLUf1PCK76Xa9kONRz3XFLc6b1FU5LVEw+
aH8xwt8WIEIOuT6kYowzz0+8B+jF+eBIT564wJ6MiFvV0DkWa9HYGvw64rDk
PkcgqpYaTn4Wi3XFvm/N2j7LFQDRDExBV4TUlAq57qba+kSeUw9EM/Vl/ARD
SzbzZlZN6YZJE0jDyJsD/aGWg9fRr190uteOrY3nTLSazXlD9K6IUrszu5ZL
lQNXWYN6LdBJZ1XqEqIJw/nSV++MQ5A9yj6vIVKDUnVRejaWCw5ZlpQJTxtc
3vLP735UiqUO9b8hexUzR17P4+KgeNy91hVLDdm7s3mKNDewGnMJ75Vtp0RQ
uKxUU4LePdu2Lfj0nY8Te6mU/VWFySIzWaFDJFTtWDQYHi1GXs02OoL7938b
Cup59BXh6OLrUbA7Rf26BrbqjLgU+jVXcNIJLqE+WWL4tdJTd79mlbyiMEBm
3P9D55avheIsvE+Tb0f0vczwjJQvHzwlJ5OQCgh7y8pMItjnVbgriUCRXYvp
IICEunsPiWN9CV3xVFMKU2mXYmUYq3XmnnElleSYPuB8nuBx0tuxLN3Fd1Ml
OI/i5Fdz4SoawZgYZ51I1184r0WYhRWRqt3fwMxV3OEiuV5ETHtBCn1GV36b
hQx3A30AyrjDKRZ1AJeA+Mj+qBrrnCM+1Qvdi/7dWJ2m8mfCNVOjKGOgwcW2
hM0U9n3KUkVqiaf98Wl45lvhBUv8s9IoPsKieLTn+FfYLS3zSoPJkSNtvCMY
X3hvyxoVHpv8j2ZSQNyjyBWvuu3M9AHS5CJMdT3P6KPC1zta2oRDKeq+cZtv
lRD7Xn4CRiBq7qj2EIMMNdG/yUW5MQLmpipiZE1Ns+Qt2YcyqfU5FyOV07vP
GaET+Rw/UjqPFPgL0lmfk11/5lHeQYfmfXvxKfaDSJbJnb9qrcgHSGmCzTef
dEUzuT6unRhAEtWmC4oGzpRAIU19P585CkcP9n7cnBofUT9W6NFp31bXe37v
qAOVcN5y74virGVXp5yVCTr4Yd115biO/fSdZL0nebvI63qmqrFVzwLphH7g
4SCzYZ1+xzw6gLwOoMOdJpNCnD+obXrpmqQIEZYuqyn8pZzaBdJe21Mcaz/6
GK3kOyxgIla5kp3G8DFk9M46FcnawbEGXb0DAw14ybVsLK1CakSs+5sRAskL
/iJFH+eNU/ku4huJupn7FSweM0KmFK4VwsAhE3VNTYoRHwe+kg+UXAa7mpJJ
6ILrVJFQ7IXgiYw7WDiTzNgHUXfJkCZEVZEEaA2UsYX0kA9UZEresmgousRL
O7Rlfkeh97i9tU+lPdqzo6bP8S9LnvUDFKDdQmwM66thcYRbA0pgPUvgdxBH
PyTD5XvoavqdsddW6Zy7km2MFQXlT7foEdmmux4NrHB5pLvmhl2RAF1VMGBW
vzLHoJWRohUH/+yHwbnXKecFpAIISVQoMfy9wl8wqxflNSkw0BchqSVfzTtE
EtJ5GJBVj91GIqymwIXOUSknU34VfCBtZ6gwAJ1pcRBs9sWGdI1zmuSH66CJ
YoOTny2qGb+t88pxuIkrnBH4uxO7OX+g4Aez6wb/djXMTKFIep0AJi+01MG/
Lw4Ot1qDd9ei4vUQKSStPjCrQhf+a88ke1oWo1g0JUj+69guNd7mR55oOZyD
eGgcKWeBvDR9BPdSkQlDzRKp0u6hDDoDCWcQDkWWS35uhuTmStQMvyeQUVJk
ycZQQRoq6rLHkEN9dZbziiu7A/kc2K+2ZBqoAdRsomopzJHlezPt4OKhd54q
M4HsA3HtoTOs9QFe5TzqO6QxFOl2Hd4jJMJKNh/vcA68G316V69hsyffTQmW
uYYs1tCV9BgBEMW6GjvcMijw86RXMgi0wtTo8ng1AxoFsHlzs/3iPGR249Tw
/WvrwmwNFN63qLw9JgmMygYLw/+crBxtfkhFGo1jBhPrzyRvSsr+J6N7qGmO
pdIdbXCwly+JmVooXU0E8Zw5tdQ35DZQQkCDnU+N/v+OjILEVzGpOd/oXWuC
wpBW0F9HaTvNyTQ6IREYamfu+jDH6W8LM5lP4pPVck3N3dW+iBzB2KE/ZgqI
djIRSPv7jgsyz8/+RvT8TuoU3H3EnNbGyVOMgFIDE2uuL9Wp1kj8MIo8sOUp
CAK1ZlJ7RDIfI63MqhApwvcbXbvvv5Q2R5vCCXjdZkAgZg4TYi92aNwmGi4r
3mS1G9JZVYrfdClsk4tvDGMWismMjInOTCnfgix7zUrJHeFXICqrxO+7PMnP
rPfMFEwYwX3E6nFEhiTdQ2Wx1PHDyO+4FByQt9AUtJtZHpxw9lgM2SXXk+nH
3cP2VV+rMcmHSyUXyy8jVRrGnOodP6zDyUomCMY9ekQbMdv4/hqipVIyzxq+
5iladN9W0bSlobD20rz2MFehASHDzanUja/OmtizUzA1jeZPfNkd50HxRPHb
f+Es4oo0Dz0IoqMejKrUneoEBcb+wsnLRnYyHthYgPy6IzS2oas3YR758IUq
ELubjeGCYCvPz9Nt/UYWghjmHTp0J70QZP+7CruLoLsrFDrA1bsbG4RfpAnL
vuYhFMRjHzWqBFMMt4GjrV2y93JfPk4qbTlwYZdTWitGjAxgpkvUHmJaji6u
hEJDjn9pzeSS8Ie1oI06BJZLRI88XIUdv7nILy7ttqZ869IlR3PCBIC64V5q
53nj5VySpRWUMMbbxwDm3/6EYDMX7qffmgvczcA0rGLUFNwHuwpfqc/0zaLL
ysQaZWFgpwGZc2kK7VFSLtpk9cX6kkV2RJNnw4BMNjf6kChDGSPk+Uaaik/c
JCQp6lSGDAWMfNnlGDMVUj+MWdsKtGADfmrwozW8BLWWt8V4t9y7GQRrFw/N
5ipESxPNihHWsjOGpldWl+99TyKkOmKe++XaOzTSBntqXpVj8bzWMFWMv2GG
lX7HDAiqWlsAe54I+l9sESKDQV0rMvo3dzc4dCPrLTWQ5XhMOc3vGo6UbJE1
Qfu2q9UFH+k/xFGJFH/iIlbpN0wzRxCLhERdilz0Ij6Pp29qxRj/QzNiTWwh
uWzatEd47mX/UwHdl0VJHKlwS6FspeDRJ7fFWfENzSzd5yFUMkS5VlGGDe5E
BEoqip0Y+KeMIvIasvL0HyNO7CH1q710FzlraP/9VEwdPEOrqoyqUNt5qID1
ZOvUfhBj8ZU31W6YrQ4Hfw/miDT32URCKbXgEqggaMscPA5/SRQ3hyCqbg1N
0DbHoLvq3mi0uzvLYEJrznZKAxak/bnWvXCc8cuTaXE/1+R558mE/+jsASJw
+RdhVQto8Z8lnSlLLWf3TeEMW3og1oPr6jvq+XVlMjMm0xliq4EaXx1v96/N
7tpxgVGfmKtShMCrCzTASKY1nM6BcGsXwrfmKgPNSpfXM5UZAT4WKgwsE7ay
X1NWP5ELBNwk5dkZj1JbftnDemDYm/4Q6J/5IbPSVP1eR9VEJbOrahyLlGMT
fycGmiINeGT2sdmHDLLAv0B/P96tkB0hgaJbdV0zyUm+KYju29e/OIUuC4PF
bR+iJ+4G24ecfZZdoA3BBKezJ/9ZwGnXvydsWU5OI3T+RnaTattrFcAA9aPW
qBn37ncvcR6fM5hRH/ziUsfIKvLe999gE832PK3dOVbIHi9mv9z+NBal6bOw
a+nJHMc3g8S3wF4wRN0VnLk5MjTeZqUIi119RhP27k8Sa4XbDd09bTd97aTq
3FH4xVjdTcAxV44CohvFrU0F8ZoYBvVqMFihFDknl8EeCy5/fAnH8eSkqYW6
ELFCAJThEshz9GZUbZceuUROfDUfdsZ9aFWJFeNiaqxwXu6CTqPvDjc3X80S
lv8qPmoMwXM/9j7jUxYF39e2AjP/AdbmCrTJcWF/1TgYau2wSuFPGfXBkn4P
8wtwxhZCUegkeP7o0OidWHkMV9T3xsjcg7MQzvbFVBZVq2xjgYnIL7vpAFsp
MDh522f5WPPlXBKOPfKHTIFrxid/ZWq2O1+RH5qfbeeOL+irZ2vxT2mpv9QF
J4dX28T/Dn3BXRZVxhq8KRC9pNcURaGwT4auGf2VzBTIuxX1qwj+IULMcqHX
n/LSos1nB12BQAAdDMwt7qq6nvcw6DKSttewauubmm9t742XI9/64kzcODjr
hmbde1XcqlIDFn6Il6EDkazsCe2kdH+WE/tGYxrrKBO3GAdxDAqmSQ0fpQAl
nEV6p9eWOeIXHqugCNmSrwAsv84kMoPpb60AOccOkSi1zpe1KS+5Fppxd+t5
qv64gEyhWVqSiLdX2iBt/wFA68+Tg9qGUyEnmT5nqfH8fAhP2U5zEGSyQGgT
I+epKcEErBaQ34MschtIm66NzM5OvbbN0HV6QxGCIR8I8tJDb2FD68reSxs0
sGd13tRe3bRmqH5u+f3CH0KubkH4imt69dOMRtBoL8kfr8y+G8lfsRTkQDCz
yr6X6G0ApXgUMQx0I3rQCqFkAwsvwc7rdhv7faC1dGzQFU0Oa4KPSZluIzi5
Qw8i+n8jRZePDrH8RL6p6ugLWtUwlYdsURyZ4U+kMyiFazMMyvT90v3qsrq1
LnNzWEoH4UKGAUoyLQsZf1NysE0VQFH0MXf7dvJZd6c/X3wCsIEqjkmy/0pw
6A0hNvfhsyJH79xAyqmP+TaIhAHdPolGUy7EEZREI0Pobvr9A4JkKvMuxdf5
C5Tzeh3EOjkUq7WZSIeHmhPeSF21CZz2hw8Fsjenm8ZrZrTVYPduF76JOa+3
wHdUb1EwuCaj2B3oga/jikLoEZDdomn+fbgTvbrn/NGcSd5LB4mRjCxxn7FB
gc/T6sEXSMeTHkTwL7X72MLotCzVSgjy/QWxyOjPdsQaHNn1nxhwoaY1vbQz
tFEj8EdQ3MDjXTsCdP9ryCWRpK0Sw29AJ+HakfFU4QIxmj7Inhl+CmMI7/BY
GoLxlwDLEEqwQVwfBFNgjqWkzbp7Y9bQf6e7UXP1C0NzlDZJhry8ssn3pw2L
rTJ0U0D8puuE7OYENvjOXyKMgyeigk5Rv1IOjrhsa/RuzyRcjO2zHnNTdmGO
saZUnhDVGj2/nMZGx6MvPuAc9OA7J80zCa11YTyLS/id1ArHokvyeI2th+Yg
rKnzDi6xNM7bOPUp7oi/9HsHrE4z+TyneWImP6/ZbtU6YWn9/Z0GhEVGO2lB
10WUQ2tTluQa1A5HzO5u41BXP9OgqeL+6KI1Xh+ubldr5vSXEvEWWLdyk3X0
6OmrMsZUO4Tow8zychGbq6RaZGmfgqHcThOQ+94kuIp5zKISB98JsWLd7Iow
LbTPsuYtYeIctJlzPnWvOG8eICicTCZK5BwWAf6hHnIAyxfB3d5eFC1KMolL
uXZEeC0V2ekzsZrTvbCx5jlcgt4xl3H/s5ArWDZLTT3MfoVdfEIh2sZWwtGa
SD0HV4FRz8z8MevIM58kGqbOfkMLzCQ3dk/j68p1f+tBinjRCC9QOLnNjKcq
GpIeAuWLguXz1gW2FwxtrNVLQG5es59p64Q/0hREalb/9LMEHWrkcGY1ZoM+
aN5k6Mu5k1Bd7ZYf9WvyjVD8CuU7RXxjImjADydu6JYl6xL0j/fOGRoS3spr
eRK8VTrB23adACfKBmoTxrqmgxk7kYP7U0GsHqHbA9F2Q1VuTHKihNNM0WKs
SYdthGyNseqj32dAdK/371rb9ieUD2BA48s4bGzYOMzaWq6cqOMCkPG3o3RV
atc94FttebFaXs+VdkUJ1d8rYwsqftQj9yLo2lvaKbAmKuMGjVDNRj6FkQRZ
K7rJgBFueLQfcsYZoNDw1piuWOfxuq8s6zaw/LMfxCVJsgHp/USgNhVzd+w3
DfJBLDPlLGYBBYzCDU7l3iIKmCx85MxcWP3Bh80Ie3yVzAdBd4PvQsrlRESj
IoIdWhFoGkjJVW297cS7cejWziIwKnSwCrIk373+DkBEV+a5D0/7JywOkGY5
COauhgEgbEx2U3mA5HKKXY+Lju1qqJ38j5EPMOpHciGG/FjMe6eudkwVpJ7f
35Br0sCNnnUWugoNrOyqYspvtmFXbB3yX/OqPuyi8Or0cm/vXICiWVOWGCuT
Xnih/Z2x2AjxtTFyMj0ugLRy6Awv7SzD5n2E3qHx9HXgflMiTQxvf3aNVrmN
dl+CrRkw9DjQGithvf11w9iXIg5OGoU+bbVXo0y9DLnfY8DS96PigcJcyQ4T
50eckQQDoNVCEXg4eo5s2f+DznC+pThO6BGymezDwHxaLlh6xihYu8NY/XWO
B3SOcCquMdbakix5QzQYZn/qpfn/kySYuD2Alx9MXyivDRdhPGk58Rshk9M/
RbHwcn1vctXTHC2mYfM/0k256TqfgWmjBETks5ytN/aFgblfiuEz6GZu+9AP
3cXGahprr9q4RBRwBqKKdki8VVHHM6uQWoFWae0x/uTGp80zKzvpoNuqp5g4
WaXYi9ChVewb3OB96puDgg9aAYms4rzBhYfXX9TBPCPc6XSRytljN3V3E6eD
idYvbsTdCzTDJCnQ5F1BuiKPB28/boAdy/ur7s/ja1+7pthO1bki5Q4+WiMf
iWU/eyGViwCzQ2NVvOs96AAj8w/u75d1aJ7bFk8HnBgmwXyjLz48EhsLcElO
C7I5SZkYRYzoGL6i9mKTeJu6eA9Zw7M7QeQ3c5OVUuBuTcziyTsrvH8puQ1N
Apif+2fK0D2laAHZ+qkNV2NNvSHGDUyQhWsD1/g4y4l8ged9/y+o1B/qLjQN
mtZUsn/dbvL27LZkOcgcZypqAEwHY4xEsNR3WifeZJv0hI/bSP6RaPn+x+Mp
3lIb9LnQ/VMr9WggU2OyCugBlHcbJkAwiM2D3z5fYhPtHlVxp7hiJH827oOw
bt1BAejmj/IPIoLjSstoDTf5iGCpVSTZ/mTl6QSODYGqaGOeKWowT7H1vADx
FN2rIqt4n8BXPA7uv2id5vqu0h1mbp8JPVTKUuTGzJ4ds3eks7LHnj/kQ4Um
nmWWjWYnxX7CTGfeMNz5+/A6eKQ2QEHwlQ+8gd5b5yFlvyDeZ61IpEMO9vRh
kqMouN+nMBO5AsM2XqiomuSdpxouKPPSPWinORDmVvSOsnJUI0i/61h1zkXE
nlGBxlJ062s2AW/v7hquuGGU6M5Dufq5mY5asYuD9VL9BGwPc2WDADb6dBzD
LdlyRMdtVezUPjTWBf8dkOSy20DzNGo32gPC38Bj8UREzZC9CslRNEfCMEDS
+lr+Uf0Eamx5VDTM2lKL5nT91b7uFcF5a0Z6ltLvDllsnfY3CLknQIQ0DX+w
6qfgjSBWRhuPRPGigKZO0WkmWU3Lbk+KmasbXfkL8pdxrtOeOICLB6SV1+ns
w3hsAm3Y+xeza0o+ZLVK4jhVyawm6RNyWPuKCvtByx6fOuAt5BcsvKIjM4cu
Psfmcl6/ka0q9lWoth84/6t9FlESvDCJmHPrDcYBRHF47zKe0zP/FfAD0HIz
fy8C3HOegPYleniq5iFp9ZinbaaZ1dhhrTTLcun6fTOyJov2+qh+v8LzWe3V
6r7vPUN5ZpimL60BX9yeR4949p2uL4V7331wffAWsld3cM/WUdo0PjiVHS+4
7E2tjblueE/z61CfxZUSJJ+MQErXHpso0If63g5DEVv628n3e/MhbS9qq/mR
+2oJri5pGbZo2cNCitVLa1b3VeQ90BmGTvOJaA1bqQvkx/qPIcG8udtbkUZt
Km7UV2rGJtPzSymfVJMsakB/TcvVgRWaplR0YnhCKHm7QKGIsBuj++iioAsz
zOYtaD4QOX+GuaCPwOyLUUIA/GYpSQPoRb7XK61MpXYfyDm2pGYv8QpM78d/
K8C6nLNvvECHbQx1qoquQjmcLB+rdYphemhD/wewYamMD6wTe0ocMBl8btWO
gJ0X9ysIJ9Wl8/SNfKFVj7RIRW18ROyeUaFG/n6MCWkC3itLTdX6nLvSMUdL
QLuMa+M6FSlSZXlPJe8MPEenTTDE2TnvB5uflZ9yXDQ6MfQWiABESdM1LWVc
tWtGAjb5oylU8LpLl4ksvlAEeU3hX909C9k1WUDgqtylMINGHLgPT/D1wUjB
XvkvVhyGDEddXeLHovW069qBYbRy4AWGJ7GOkguodStStsIR0tyiyQqnBu0J
c1AGLpyP+iRrJXkJAt5hwhitVbNUgGVAuLyv+HDhQ5mpobG+oATwbqFSZMHH
h/m2U4bzY9Xj1tA+on82XAsc0qnIUQ0Z4wu40TbLqzOUJfTpcbGxBQDK5rqr
mumtDLKf44RTJpiiV6pxav+lrAspS1AJBU7qY5aWX75lN1/s7V4h1LfnJqx5
+uNtk6/YeAItuaNdB0dmP7WgA+OOIzwR9ypXCg3mD+2+InatsXaDb42bqRnY
BY2Xz+TNyL2eRyJvKmdQLEBoNgV7FShmSxcFODklg+nh+MS0zfusiLI3dr79
DBGnPUOGYXgxhyJj4bSBWPV3L4KtJOInrG8xHmNnMb9yiVUq/v0q0l7PjmbN
7kp9m/gyPY+RrN0nAnsjZKqt9oqfTthhZYf1JNkvmDCHb7RR5DaSuTljIC1i
HES4T3MlordRIV6qiVg/rjPwbz817RY5a6vWzIbHJdJi5pOVswTAMJHwozvn
XSmurz1kYdVGJRyFp+gLlxmAf2x6zZjmk4V1LlcmbuORYQBNdgjcDzUCmTZ4
YWVUQ5eVUDpvCkSEf6RJmNoGUHAR8Bwv9Jl0FWeaMXXLxy5OtHnRO8emYq+L
WRXIy4dDInH+pt1aUfx0VvWv5m0w1eRXjnsvzJXCAN+T8CGAltlqcgKejb2a
Nfwl73ZQE/P/GX6rRDc0rvNFvdNCVja6AMIT0FspFhXrvAEMmvZVZblBAE+L
p0nqT9vfef0i/V/1mfaC5Ou0QvWL/MmDHn1NrJTQjsa6hIAdLb1nMk52nPeJ
RKsNtG/KGxwaiAZkQdVapoQ/Yc3HLdcGXE8FPoY/9JXz4qUOUFy2W/ZWjld6
iWHIUesWFQuw+KL1sVSzi7FtYoq0P2qI9DrgWdTZXdV0ygVFh8dY2u9lm1RK
PAF9/LRXQkxTVFGepeRVvA9gC4AucaSKxlkzP3In9Tf5Q5ZkzcuSSoQZ10am
N7Zqo3iNmAKIqZVIdystrtQE9VMEstl/1kAhYGt9fYfrRhrWMLsEeUQ2FX8c
zmKV5EzsweivQ+mnNU0wCuVUUTovPskfytaIcqgLh0RRk084HY/wjGKgsyt+
/dxyAfN2w9l7f+SwFtqfIX55vIssCa0t9Jksymh90tqkp8XQE7PZpaRb7Z7E
GPQ6JqkCQHI9YyO8Wq72XT/KeSqdMEdBE3+8EDdH9xXIcWOIXEr8i6GKbYz9
O8t12gfm6tSYxBa5Resi5hDQiIJHk4fA8wVSNf2p2i8QqBE8ovhQ9pXPurZp
+EhxAMTMZmRq8gzHzBeknpoZLQajwvLskSOSrlQHLqkfYG0fFsBGKlcyW9y+
YLsK7k5nD4o4FyLTaiSwnUlrVcY/D3SaLPTs3ESUmXcDpPKOX+JWIgvdfHgb
82M0J9o+H9vjNGrEWzs4V49OkkKR8kClrd32jeAOFY+JwzO+pwruGFQxTdEB
MUwp25h4knfrsKG92OFkHZLQ+JJ7k/n9WVzbXokrKeNGmJu5rcCKuDV5xTBD
rwnyXgt1BVwdqWHs6pq5r3+CLUQeZAU/fPoKlRxsDiik9A2/Ml5YbgUBIEiP
ApVae1znOR0nTukSV2jV5oipg4BrM5W+6aF0sY8FN8I1dYdvLnFCpqZ23old
rie4gAUPFCe2mx5rWxLOnUKm7e9UXmHCCTZ+DjsL6wGHJSiPFVkS7R4h2CQf
OWcvoVZrb/W/mdGbh/nrRXKENrSqsFP1KbS/BvQ5qQWblA34vJvHOQJvIkZN
t8n1jrqi4V7/ps7DrgHmX+CvRy3t8HLkbZBUs0Kenb4TRRmEAKXD/xg86eFa
zT+8cZQYk0FnOmTZLydg043WYYB07TM61+nXupVG2MEOB8XJ4+Az+9Ks1HkJ
q8pzTytseCNWt+baOutOmRQos/d221jtwgbGhKhmznQSjobms3zXHVMIdmKe
HNEWPALyBv5brtDEKwJPerDQM9xdvyRPQyhnR9qDYtsSC1koCdj0MF61LtBV
4TKZxgbW/e/0XYHzKrbP/SBZLCCfbI7Qj2TYw/2lJJBCT5GzHSYTcsUuURtz
WBXY8B8wCvZ0UbOv/fzuzumb64egRrpEQzQlrpcLLHGg0TF5AnXlPH4evDpi
52Od6sECig7hRsLXq7yN/FaLA4K7YOkpgDw2WD/GLmpmVW8oAPabifrzHO3F
HMTS0W2GZVLV+D5TUZLJIeV4AHNY5mgVqQSgyE2/UnG5N+EtvZJGz+4idZeS
lx9DDpIIdWS2CwAy47k38OLmCZkVGbWs79dJv1uUxcf4SG6JdiE43Y0Hr9B/
a3qENwIlIVtgOOH0HyA6MxMHCZ95fAKBwFt1fnlqKjuk7vytIzlnf1r2Bzh8
G61GR0AUNjY5FmUJ0ir1X9miBHhayalAf0d3Awxg0eqT9Ejct9uoanz/pgTF
L6OP+5qlQjdiU/58nhX2d8ea49wShStXE4ZHPUiC9FJkH4OlgInHmeJ7B/eY
SWrerUwUaINu8Ad0BaR0hSFw1sfQDCwYlMtfIB3ikqNjmOqZoHRW8Gg+8eQW
PrHEbofTJtakS1AU5T3NKXk7fty8HKPImlOP0fXAEtlRDXpiyC49pB7DjUAJ
29dnhWOofspXuUbbcu2qpDmnwHCDvbCOOMurNY5QEnBZmbXnPPPPwQdnC8GN
P+/W9iigAee3RvYdhk8oK2ZRGDQe7ZtR1h62B9EVhntEushWrJ9t+SYtu5p1
1IUWZ43SCtRXtiv8XtfMcZtkTMPzBicIEPqR5cL88RHD7j2qL+qEx0Xfiean
FxZfsWgiwCkEl8fvX4SQ+h39kLA724alhOBwBrXIpgDIWqF4lM8C7MEyHCkn
ZIGMD8eFeJaQsOxMCVD5gPtAS17yKzkxLnmY98ko5jy/CTDmZmrHeXAVa8lV
wGxEJoZxeTfKaVBFVVlUZCp50NqfDd2nn2j4QO3G03y07JhloSWIJg/njPFY
3U3Iiwfqg9xh+EdoVPEQh7IrCqN2lksczOufiVaVJ3v4a0lFKBkg5c5QKaoK
QPuHY2rSa8XLnqv9yX1FnrGewaUsxOnpQVaQnTfGh1gVkpx3uNej5BzSc573
AEEz4vrf9HDEw3jvrW7mV8d+/HGXvcw2c/j7TMtreFbmxdmvl7CAn8qVLp8X
WKOl42j4Jsg3VS8OWJHI+uKqKqzsQZF4JEYUXEEfIZ/L3b3B1HbX3hcWeuhf
vXr7EqJzZn0aqZOaP5CAf5tWMkFtuP6bxaVdzSvmuBM3Nm0GfcV9wDGB7oxz
hkMdrEzbb0BojwHPPEwNX+VgQ2xCvFNmDRPYtc9hQaq+ROjKsvPrtpJOB1sj
8YIEcnpGu2ZDQQS4PDhwPpJdgistIDfTHxio+9ndqJmyl4vBe5HjQf++LNZz
xyg7PCsSWpnXaB5OWkRX3gmNr9bDdpHIVOr8cTYVN5RRCqzetvg6SSuxcMH3
JUBrxRQKi5lmtwWvXzHNyg29kjK2YBTkvapCUlgDuRpuyHxZQX7pq1U2LvAH
8ny+JKAQopfp0JoasXPGpIAzXJ8CdOzEjIRpfAiffP5JNDyCml/oZXgm2/AU
PWBEHGLoSA0C9vHP3auSeArEHaX0ASD7aHeuR8qUPunqrzPgirE/Fm+NMlyL
TAwF43pO4eMg5sixEL/Htuu+xRqZXGYK7eTFaNi4FToKbAZ9xdWRObBLTNmy
moD04QebAdjyCXe/FogML9QJQJ6XU6OHffJtobjaUK9+oNfQzvoCNzicO2gE
E3D+1NtIQrKiVgvpvtkw9ppH9o8uZK5R1DzHY/8uDlEg1RUG8NqKX5+FC9JG
eb8eXNHd4Nm6Uor6PbJPOoW3BOYlxLt4xUPDmIAj03EUCuELMYrdHEiiElQw
2hh0XDCBIcuC31RabZuQ+Ik3yZpXW6t2eGu5z054VlfTUP8B3zRn+hnpCYmV
/514d8unmgkdLZG4WRichbQfCR0MBAiAzD3yJuSBKlNKNevOGzQQytLefJc+
R0nDWTzTCTpHuBBq2eNR71L8/K466CBg20UFLFdoll1CVjIKZF/41O1t+nrv
mC10iZIv4wVqmd4nT3KLODCl7XvLLqLM44wq0v5US23VYqmxrTDJ/y0Mhj/a
QYKzSRB7AZhDT9jdK7BVSjoYKF9es9NG6NgwdQ26oVO+Ur0i4JsVjRU4A/Cm
5D6dT1O5jQiHOIo0bb3ZUl/9W/BfRHKc1uhf1D2EFqnhosUHG2M1hpFMCy+g
dBm51bPpuHyuWffYodTUDFFewtDaH/jYrgZvg+BMnvSgp6gDAhE5RJMQkjvL
hxgNSc1VyQ8pIVKMkQ9pvqmHLFWNq6/Cb1QazyEdOJsa+0GT2tkECgZ8AvUa
tiDsR6cZJ1I3EL+oluZkWPAtfJ5ehhHIMauSptj3kvEOo37UDPbQN6DmVDBV
fdqIHKu8FSUt41S7sOCnCXLS5Y94YnQrrRZ1qYW20dlBk3Eru+PSiApwHumk
8CI0q8G5dhYbKPzTD+cgAEI02ge2mKGjVr0+fvZEzAkqXOCKlbMc525cxg2t
8CkqeTKE9/o+3Fxk0arulyurjdQ5FrNROmyD94LkQMICXFZaNXpDnJ1sDO77
z/eb70bzVPjljhEZilVEQNsqP5xQrcEkcZNS58EjOhKrW9tBTfZEecf8Hmtd
vjdbmuMes/06tMhN6+FD2nWQ7r8RS4ZAjGF9JoP5leldZpyKgql6XPHnaLQV
1l34AQp5mBJnopThOsNzJ4bUUPEMjJvZejbgEHyANrbE+MGN/QfU7II0eJny
YovtdSddYKgVChBF4y3p+hu9kVGYWMav6W0XOk5lkkZNNzxH6f9ZUmrxRwlc
OaIL8txoTqA8S10d6UK3mc/vVbjiH00EnEO6N4xBbBZwQYdZS6T7jOANECtM
mFHh3ai0k7tIy2hxf19ALjM5Ne/ZI7lUA5DhS4KNRBgsFGxzOtJGPA3wZwno
03haNHaiSNmdkLoVxBKpbKFqk6A4N8XXt3A7pb9bRjguwvGJ9AU0qGnW5SGx
Vej07d5Q1LRfflKWUy1SEyyKOb+dSlYqu2yfcc8ff6P3OrUnpF905NjakCDh
6g8JylWjYJnUQXAY+dVe9xz0Lj6g2nQp+Q6SWqw+mv0J9FRymIrQV/2hI4hl
40ghNgCminGBdZJo9HLUI1qahaglUxljJQFu4GkCCKmI12plFwxFUzcAocDt
Xf1xiLyAAcJDaJ0t/+XF0b76Qw3Tfef/BDIpGgDZJ6su/CR3Gk88JFZx2VPh
BcTOkqTYtlmfscuUdwdGFyTvt8jJhB8/gkMHI9PzYTFb2esImptdpCdnSF3n
DN5tLeit/TQRYsce0SE0itZrLvFs00yicZXdXXzwQqTOVQmv62DTQs09GKQF
Rll0+NX2zukClcyZpmtyHR6MEZwgECVLFt437slKGCdpxaIqwqWWMo2NNcU6
nAVNnBxcW7m3ymhBZOLTKXE+5Zh3Xfn7ONh//zxdq1Utnet48cEsdOLCw0xz
cJEvHba9yGjwx1kV33O+g33qrH50s2t4u7AYvPdQVtaTBqQwGSa08HHU1+GR
xovE9whDJ5lP4L++oUvQ2gclBYkee+WCCJJuW4er7igVow3J16Z0qPXAfuLh
TFqzDoHT4Qj0VxCylBs9uh5Gbuqrh6NBwPvu3llIjTtmsLsAUDT9X2y/TYcC
GLePGtwIOzf/J8BWG+9QIXX00uLXq4+GQB8+S/6laikKcHigDfVTnzFLtL0I
7eFdQVRAJyP7i2hIFd1OmXd0L7BnDSu4TiIZEoc6an/AzzlkDJrZchfUnjKM
o9E6Zcr2A5sdlYXhrROW+sbmg3nDGU2vnHhuMDZ/8nz1MZ1m5RBDs1q8EpHD
E2YcSZfGJPc/hYNMWORZ/910GrBXy2NwyvyhlOs3Jozne+V9wz2LFh0yaIvz
znx8zYY/aQWFZtylg4s6GFBsR7E3vT6YyM7dd/RptEBsBP1c

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzf6y4v5kzzfWKspg/4b+T9vDVsogoPfm77q6ffoDGVrsF6KF38sqxhla8GToaBxdpMGF3DJW99DDD3O8ik8MnTjaGuFMnaT2WMVamaGcNcOkHnGP5/Kl71Ps13PdBRGYK6mUm5cm74X5OzXM0n5Q8c0Y+OcAGfNZpG87d+UbjHLD3ddv4HntRG2P9Wv8MKA++J0fzQ3xh+WsKqNcq1MAVyQb9/VvyAdbMeyGsO7Q8AgGu1JH4/TNE6+aQW8jtjdyB3D6HWxoo6wHOy97S+PACcX0ViSgXGqSPUrj8opV1CnSINpUk6uJrOqEPIIJf4HZ9aXJ4kwErum+Q5ls7ZG0WUtE9G9UEaVKD3UjrC1Puw5XEL+RqAatDAMsyK4xAUR4Jr72AtgbqQ8Whsz1QjAajwcdppSPLTiB9vqdv6zkf3nSZ06lDSe/ooYAnTXcZxhY5SOZfbh4s0kwEwN2S6owpJp91bobKoLfpmX9xsci3Xyw7SldanXdgs1unh4TLpGtcxkOISMwgX0A2bG0OoH2zm/9eSDuX69bEIwsSW594DNVBinT9NQxROtwAlPHJjLLKsbPHkh2EMoDe4BoMnA6/zQ8ALeA2Y08V6ySaMcKCyM2FGxHdNRMEwf91ipQSfMrI9XmUJGRvmUvPAhhbWc9Gw4tavycsVGsapb6yh5iLOa/CjzO8kF2Ag1WHxVqB4iecX+CLABLOEksFQgu8dLgadOn1318wyjrVTJrSG88zETew5DMUHf1+f8Yw7HzVR1f5PEywAdEO7ohUR/8RubnZRi"
`endif