// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DZnKIJK8zmn5iaat0Cx2+OkEWimZFBRWNbyVzi5EjYIe3uR4FJ5I5A7YJw4U
zCvs6XdTbedO+VQKYElqFiQ+ebAlBgO67VZO+IyJEJvBe0HVRcae4OwBplyO
rAA4CZz607u2WJcbjSZ04OiI1leGuOwLmZyAbuztMHPXv9aq0fQEZm28Vl/a
S4W/wTTy4dqt6AMLf5jZL8YTZAagSoVsF+5KnVLYrD/aXifk+AyoRMgkieis
BTgdCiQFdkQrnRU8smAEnWlXYIcXMMzcWiLfAXcs+iiWBf/9HQA7hIXfrIHF
c/heIUEf6w+OBXCGKYGoelpotmtcQSYuYWMzQOMCHA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZSqx+TfJ2LhADjHJZuYbRpuQhxY0kf+jyxqjESjZmtQS1ZQP60PH6Scn2he2
LWYOaAKxlhUIegj9VkR/m1K3eroJdhTYBGF7LwOoYVc8Qu4vl+M1Xofpdwui
E5Q/9RFPOHPIYxw7WxTuCPCCynejVsd39NTOiVPlL/VsKgqU1wKCHVBiRPdX
y0e6+rJ08rNYwiMjfK7pcNL/cSIhAAq5HKqYWZb3/YCcsPZdk+yS5ut/2Nb3
lZtjdbBkf0NKD84lu7RXYaMo4xzwZdSSwQrs0ONrX2aD0H7N6+7sbstvrjfZ
ghuLsqbGol65GQY1XQ+T8KPC8TycpVaEssvOTNu1rA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QD/a5WY3peQSH4G1E7LedsfC1W7dGcRg8Hiclpik6NMxlhItAOg7Z1qAxASU
/4nnI/hEtcPWnq3Wmc4h6WFFokuoA7ADku5lMZz/gF8NmIzMy/CkERyxpyRn
IMDwUlWLeijJD/nHMDuGhbD+wZt9EEBF8vURUCIPYBq8wVpBRjNFvWWKNPIs
PY75KkkQgCc/pd7j7PQHgS7Z8v94LRQBLnCBE7HOK7UMnOEHyMxaEQMtVvcT
YVYEg6qiay+dA/E2UFbEggVVs99wa3tBnE8iRj4xBCZeIUoG3UxsPtyEPSd5
X52MMrN+7trhLu3O1BEAC9BNJHJRAJROwpLIhnu90w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CrRKlVL1fG44aTvNPOk1O5eUok75yNjUmQ3SLAU4bCjaJwkt5NASHW2njIGF
Bw6OnaikCal9wz2dsZOOSfZWiha7mCIl1+EuT8Ncx3OMQPLEmDc9qGoefZZC
0wFrHMnubbLiaF0gN2duyrmbaJpm8Ck9qVp9vVLMSv//ukSqr4C9QK08yaeV
avNRA9b6GCbPlOBJMuAXz8UUXNBVi7HN0lBqR/+xD58Q+/DGhvTQMWCEtqAK
tmS2n3KadXyIyS9jXXFUp1fnpAPC7ThYhpgKYuvPUUiukIISj2Ffd7pKSMlc
bbOoPH0/f6qmq1B0tgJPoWRA4IyBCDajHnV+xrOsoQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D3wqFSLWIJ39Zp2fiBnlc6VI2mkzKjmHXZyxzveciXvtTj7OyeN8H8uYGNPE
quHCkTw4qvaMsAwosn6Px9y2Z7En/7bJukqevU9j8MhDJqfm5UoZtnL4Pgkh
c80JzdReTm073DZNdbP4ZUpIYJ5yh8psSh/+LNA9OuSLenk+qgA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DsYYNU5ywUqorhVZA6mI3d4Fadvvm/V9z2DGuYIEu3E+UtGhbUGuUr2+7BgT
g0MpupSjwIBQunoyBXc8vfDoP4UAZ1ARbQXW8G0v9/Reoc82vK18z5gHe+Fh
xd7LTy6viIS+bYna/Qn/GA2jn0SFupqsOodeG13rIzvjcF+bm7klbY0hntLj
UMe7UQ1DllvPLCerSXQLbk93FMsr6ymx+cx4MnlYW+Z9EBIxBtLDxpMbZQkz
Ysy17GzQJmBMqUQgt91l8P6bIKPrW8UceTvnumjD97ltQSqNWmSu5sENocc3
ospNFpIWX1jVZTaRYxQCJqRr8Pc3ekoloxZadv8xNWEMWRkD3VE2MvicGN82
pIQHng9jrlHNgTX6Tl0hETDkn5FeELN/mmZ1mbVDc1QNWTFYwTDdcS6M327H
7zSoHI+0DVRRg15b2SkSpWY02nkjA+KjlZRDktAU2dQLNdn5RGSRyS69am59
sRbLjcxqJxfYVn4wxsUvLp8RrTg/TO88


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
liyoeVcMPGyX/mAP4oz1GvyGdzwZCzfrpq6UyN7VEeJj2BxuVxf/m0Jucbvl
jiHkGhZwZDjO5TOFnYiZ0zfaUqPCyf3MomvsPWTv3LgzfFAmzio5GEXHxrP3
IAjoGVgbLjQPAws4VJioEC+ObztTNgdh5zhOSZqx5nm94gIbuFc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cXg6YiK6ucpaVtvPfqnDezN7H4E7iV3YELezwQxxuBTa4PKoh3AiCs972Z4Y
YVWtDz9aptj3cR619mYphRaNeM1JB2bQ+cipR+QSMteb9pG+iUxWO9BfkLIr
R6rqMY8EIeLAfs31YhWso5kMLG0WjBjB1i4YRQHX7fvhfhmO/1E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 74416)
`pragma protect data_block
jRHCsyKJ532Nuiq4BASM96JtVNgtW/kK7wNbeZeU+mD9/vkcRqXgCnvOayYT
pAeueJ21c3G5w1XYpbKstqegNvdG06tD7y1gnhkkChuwBx+vK2p73zVSYIXW
HjggX2/bxgkMcB0m9D5qkWdCCs+S/08zZ4uPnFU49Zz0b/wu2uCHn992K5Ui
qXUoMH5rjV9UPc0Q4WZBe29HB/WMiaRjRmV3y3yHg0tp/Q3tUZ/67Ag+11P0
CRLKbmFxgbbdzKHAi0zPzpJJYADHytzkeYrdaSHRvSQ3bszZXSjKfSILUemg
yf5xCSqFYLZGEH9K+nTev5qnecmPI0eVmUtoZdZIGRq73QOOCr2LC8NlEHq8
C76UQqt+l3qmT7xREuS3UDk8JdbZ07FG4C+U2jGMbc0iG6L0FPU9qvhWyHv0
lSlYLH7jLLeLdQ09HRZLkSKbbC8dtP+MKeyQpR4G2DUcJBEDGAha6JmYIrfP
AyAne5Pe4+LlUmfZEo4Is0AHrOMlctyygZT5j7irrjFuDXQ9dwgl5p2mLFoq
/p0YFlNVgzqqcQOfVU8lgH8lEbtAUhYejptV+Mpm62V7mGC0XHXwA62HnhDu
bx2KxAjcgYuN72vXjU3Q9tv5dHX/ivEi3udYm06tdtp0hIdMYJ7AM1DE9epo
BFzCHBuDFmlM03mCo0GWtjeMhFT3lD1tkgK71TPSDOsqanNHpdiLF9NXxQM6
wN7b2tagact31rA2VyThj3Hf0y8vUNLFAHr03njzBX9RYq0Zn91BVZ1I3W+d
rHwONpRGlvwpjyYUWjwhe1/7tETTk4xjcFaDsXZ2KnBV4GwgSr1pNl8DGEhr
duaJ14i9PvrVE0KI2xMHTM3JILIw2eftpQ04RUs6drelwS7yLHT3oVhmbwkg
bV0cOnpx2M/NO96MFHz/Wx1jiruo/ZQgQGpxq4K0KZ2qmMPbfvUSGcZpeRxg
xv6IKrc8RUjYGP0CG3lrSn/y7iDLe/wregyZ0lksrvybw5m0XWFYStBjmWv2
iTPeS4RdCSvdwKGvs3h23gsWO3oUJ7B4OUvS28AL61CO8JHd9GSukfqws3xk
h6lW/W1lXG5h245rYDUMe/cgB5YpOehax0tP/KzMbqIF5IWvdrXoAONUC7PH
MvEvLzESRwqclV8mT6anAz90QRf2/ACW6H6N/PtQ37s4Czv8UdDwx+zaRxum
yIoeHoNwHjRY+ufCBv+DUqrdAYo4d1kaOl9u8ApoXuKuKipGFRQO0jInxrUt
E1JT/AnnoVxD83vnSFTB2nM4NWPJq91Wcz5j1pJLsitLUOmQHdOdYrMV018o
QynRgKq1xzInr4QFIZER0lnr6fEEzkqhMx9V/nR+Qx2doW6MP+QDYHjZ9Fkw
vR71wJiXe0I55bO/+KYyyASqiSZSQRFdr58coPvUYz86e/L4rGeA1h+Uy+Gm
t9PiyByz5iCWepOo22w79ifZStveYcs/O2bHlpuCClhbyG3R0WSZNr4u7/sb
2AH34T8dKU7aD8gyybH8Zrxzi2aBz77PlFkDrhYXtD4g+WoeXAXQqJgJ1JcZ
JSxniqLfvGUNy37ho8E+Aob+C9bSpjYqcf3TRwV6jzIT1Kkznt6lwujNWMnN
e2+OSr6o2ynl9WNrcE9CpySnCnbsJzLZpVhMHWJVv/sPS+sw7imJW1yCnadH
o+fp0dqUC9KebtrwIKbVugQI40EcRYYTUxogJujOp9YTi0MHFdxHzF9qJYVX
Ol4wl59FRsBpvdbAbvPA89pbSHaJqwntkbbCUNn0uw49aDbxEiTfSCjZKxkx
HlIWCtd4B3aLr7eyuzQyVYZjNiukOW8az05241fcBTfDecW5FNC1gQRJqK8W
nRMAP1UuLKTTghQWbM/Jb7qlDP9s6vNycgBqLCiQaEMhHHoa0aRv1Ipx2ptn
kKL/pWKf3cbvdlWVsA0hb0xVjBLCPXnUUlAe0xwiMwyjBVax26jbD3ZpimnL
RWi9LeDNCBN1Mk+S8kk/ywPxoYXr0f3qiwc+17Um1cMx+5SInRGrcsJgFFbK
SzaqW/RkDqdwUDrD/91LDwiqGa+iZlS+gvf7/Qlzm/rNzRg8czh/ac8mE+VP
3DHYT3P264UgLgG6iK6HS9C1/wwQwgpNQ5dn0WmD1ntLH+lENWEGRO3XPL6q
D27+ug1Gnv3dAbLZkfifHS4r6fMzeQXFRi4oe8xw+R4IH289OF4RzyVImgyG
S3FAdgnuOOpRmW/EQFZQIP4QRZitppa0BVkUsUlUR8otVPaq8rzlgcjXLsEh
ynGHe68lmk/MCbGqIS6iZNPxPAhZ0PU5fTQnxK1J7ElJ3RAf/8Az0zsow5Vp
R6zdA+qnegguIXpDKLKdtZfjhOkIB4Nt19L1GjBezjc1jL4mDUiqk6XqyUxy
DwJ7HAojuHEhF7hRxLYMO+zA5TTGM32PB2XaxvT2oEKvv+EAH956wLMxvETk
1wII/oDGWQG1qKIn3tCBjCaNC0D30UWn8kBnEzQvrFU2oaseZ6qUQgoCUiE6
a5vfPooapSENsCjqsWD31mhGtMn8imaHSoZ4pkm3VE9abitmdQCh0FtwIX73
cW6USQY/x9oUCuDpXY35DJEzIdi/VHO7cySTkpPtjzmyVuqlTX7PhtpKDx9K
YnR0MNMFakJKlRGoCfcf4IfIECr/tTXniC+itOcjqh84U6c5WWbQCVYYMHcq
N5IUjBxERWsU6zpikdHrSShwRuTJsly4IXP3A02qFkiIBcmG/1c6hNX7vLtK
2l17ojeRt8pJq5F9xa0yj4g/1PBzzbJ024+7O4feNpEUznWpXHy7jMf2wSNx
0SMvmvkqIEa8lSYKj6gM8g7GaWpWNl7KwlnJRVT3EhrPYWGrgfoF3s8B5+yV
tJwM0JFgx4llDLj8vPPzpB7wQU3MiItr6XdffviQtLaArC6ZY6wkYWC3PgaD
JRJfrB64mYrZC0VKOpPnaEFCRfF5DmhziNn2A6mV9aXsRJzYFGydl+EGZ0m3
6/uvXg84E17f5wyVxZp+P/e241JBx+ybr59VUJMNZhuCzqB3ddc38/r6QZA5
VvWBq+W7CKvAu0rfRaH1oukvILO9eNhLcHDZlQG1+X7WByvVcln2BIozoeHA
g5vzFx/sSQfDBFcmAxuOAts3Xw2TcenzP4r2ikEz9DrfdIZREz3SKzYuJWQS
vZ5tt9WltqjZhb3skXLm6lP6Dq/5IjBB+iImHcx2lpJkDEEMimly3Z8FNOLu
gBgIZcMMzGkG3OEXO1ltORsdolArNJHjM0qULmsXShhGPwGy9FwZoN4zv9qv
Qt8aFh3Sa9GyKDNnPt4QPLHwjjfJ74JG9R7rsECEWAT0DoYHZR2o+j/VFEN7
lgBfZPa5MONiAybJ2mHow8Yi68GTiNppTQZhdRF8dJ41zPUXKjdwlsnTLgsf
PjyOsHU0eRr/REOrx+v1o7GOaGJcaBdA4EMs+pPGuLpP2H1WoQZzsX9GM+Sj
+6b2Iq5WNb5pQji2gUL+jh+Jqlc26RACmgfnywiHcS0wV5AWIDFbnV2tHSzJ
A1fgA0ht1i1HDQHHsFzLWmQIM4Fk3GCtjOUSRBvIsZb96pDWb7JD4ZvAjxDA
4KTvhrXGoDjrczIq6P0Ev6Ajk+/piozbU5dr4uLDmFv2kXPVtktxHz7/Pheg
o2jdiTk7pRvBlfkzyNbAQ+YNQ4VBnxy9JucLc17idpTbu0ILTob8AI6ARzot
Z4SZgDgXoyCGabC2udjFFJ5qcoO83cu+e/kXueK/fdGtYMetVMOuSho73ruR
/lKE/+Bft1WuOJmbs8pbiBfMcg/B+fShDYIknomzM1RcIBiQ6GpbUhsB9nTh
4YCiEk4zAH/Pk3+YMskv20aK8EaSNfJNkci24pHOlCz2dTIpBLHEOLd4fZcT
LyLvYfu/yNZZi+K3Ihv9Pxlb7bZJK4yNloh7osZN1bUNEeHVK+BBuN+hE+Rm
+H+klcqMQqpFNw+NX7YIaZmD3Aiu7cQA/gCZhIUIXG4G0urTiVE3jesbPwVu
5fYnz9w5qcgrGAo2JYMDOjXCN+HjMxKl6uu+Mj+FsbaVUCO6667gacjDDt0A
pb+WH45Rs3QIKtesv2fF1Oxu/uDXvdXCneI1f2ZXyj9X4fHV1afnuW/Wlw2d
7lEoF5Vx+kOEpEw+eYD7ZFKg2ZQb7r3A60LUcRDGTONG50oKvwB5/x7GOVv1
OYSHn/dA/tzSI5VCL/HCgeumks/BOPMOcnMenyLy2onTsiPoX8mWpX6iko63
M0w0UZLMlUimeFq2fnae06RFLtdPdP22kE9K6hiwn3XmpaPMEc2kw877pFFS
0w2U3GI+qoTak3HvxGTdVRw2SMifvAvTF6qsqXVQ/nFJIoeMeGFcxS0f897S
qX2rkctuyq3D0aOvvmxrzh+xxKjWWg3ZRzfatCjQ3eR00vll/8z1/3WDAgGn
2ZVgd3PHO1J1yFbfNuiVf+0RNaaAFiLSJHobHYQSt408wpp8lsxVe9/2gf2k
ugBl90DfzazRwk+aWqgGvxOz/NYwlSlv+B3IOOBSvbxy0FYHmc4lhADPVLCK
aDKwWP5OODChpqxmWBrojL95d1omPEo+5bN6cbvcmlBtcrNc7wY0RBSFurbK
h0SH99dJssUZtTu8KoCQfYuORdZkygbqgGjwIJaqC3pNSf+GKH42CjZyQFOa
PP2THTq7ZfFzp2v2LG3NyJEXcydSKTiWsNOhmfTCYQIPMKBh8r5FqQ5I+9c+
zsuxe0h0RiWhccLy62njBZrY76QYlZ3va7oDV3yBQm3KW28Z0eB30mXVrORB
hoHx6sZyeoY5u4nXrh6maR+JLN7zVs7Z59l65qOYdxF/Ur9mV/4QBQoBtVsQ
6Em61Q1Ko8i9nHrN+hco1sPOT+G0Q00xF67B+PivwmXslY9jacwfgr+1XPvi
6wB9yM5hIlraD9mkgJKM0fM1zHJcCxaMlRAYD/PwAIquBHjNUa8VB/9K0LN3
ReogYUwF/J702A3BgB+3asCl8ufK0fPoGaLOPDu5lativOwbXNNBieZn/+BF
0YIowmeni3Jp2MSanp3uE/fBidB8PGO5D93QX/dYomGkMktlIjWHD+1Wr1OY
esqLTkpr+NM2ona592VXuEqfYYZ9i8GsY2m4TXd+cgfJD6hmYOtj+sOeBMXj
Iz5/19VnoLo5yVKAsX3uXGsOLfu4zF56SZ5yBg4HWkxiK0l1vdRjVLl0u+cO
Wi2dwQ3LOb2Q6GKGs+ubWZpgYMSUW596X93bH7QlgiaZPmG+PPZ4ygwAPkz+
L559d1QA7968CoFUCry5ybewoj7zLM99FtzcAnu4ab7CPBqXN2QEbNTJuJSe
zbr5Wg6NNjGnTY8sJs5PZ6DMr8Hu9920/6n1J4GZ4VoJXeDUgb+QTTERoHR5
VEkOzafKbP7/d85cI91UBj8XmwK2gtGRftyK0v5iq21mhQ+Jk6ZuSSUYR4r8
NaYaFI9SlfCcQDzQiYZ8Ov9j0iwlFDVCDSZ8JQgf8JemRmlWwdrtKWq4HwUn
OxnhXTDqY45N5R6h70CyVGr7AGkdlzhVk2HsChP2SbwPlv5WlPdFNF2qH5SQ
znWhG+2jR6G3JM1uYFO4cewbkXvvU7qGtJQQtTaBNiynPweq4GbBuCRODKDO
XOmS7Xk52AdihGBfrFsZj/rqbNuU2wpnw56NQsrbSt5em4yXgHDSArVHwRx/
T5bRj4+C9nyr94dckJxx5lKqW/AYp885IooKwDU9vT5QBLARYNEIDhTbAUqk
r+2Ioc4qBuCTKDM5G1KNotYCLrlwAiTgE6Ld3KDVqobvU2y7iiOqrZIx2Kd3
fw324FC/ruLvdQTp7W9lu6g/pKU97rXqrJZS5QmcTOgumtpoHlPJ0dmUVpF2
6Sl0OpAQaon5r+grUkMpv8iMunKvC3G3G2sGAE/HjZORMaEHvFHNWxFWJnty
wlhTMFCRihkRImjHS9zU2Oc/vQ71GfT3mU/dicSG9+sxNbqWdZyaAckSVEPe
njieCMGmh0sMMW1xMCumHwJolwOxVK8Kqq2iXu+5TFsJS3V3sL/SQE03j8O0
UqAQ9FJmAkcXc5GBn7s3DaNYLhs3qckxXqdscWXLnRbufLEOCqtA5mev9Vg/
bKrGd4lOUJFeUl7rFZ2Ji7GWVswhCWqzotENzugMbvE2xWw3Qd0Cf5TC8HsQ
xJ6kVc0JC+kVCkywfEaeJ4noMnKApV3ejwnDeppqxrEhA8RYxZI4KQV7y4+G
gdk8kkFQoYXGkOHkDZWO+MbUhyvbP1FnqiDNZC8BqD+Ij4hRA9mIIdj/al7F
APZp4cilN9aevCGExmK0RuAK7FYqYsSjrsL9g2jxa8YlipCLcd1br97CYMe9
C4AgvizZQPfIUH5zO0GIBN3tEd1t2PZgbsUlG+tU9ODciw2HfZ7RQzPNadyM
T98s3FlY+U72WOo4mjgM0OxsmErtD+PITTDS6WB5zzIm/TgwEqIggqL0wdYo
z+j5GRO6KNOAZ4mGSyAdpvhtmMd+OObm0oF+84YnGUb/Znw0yR0sYnTI/flF
byYL7blIIHWUWuZeqyMuvf9KHjjz5HufIEbDHSkgzth47bP5E+Tc5D8E7nCQ
Z5TbbXqMpuSG9ulXmtP+HE1N0M2TAYYKZh3OueVmtEXNGlaYFHLEO/vtQ75f
7SPSrnvvNod8jhbl1m44prqwRvK0F5+gEZzlfZcdcAXoosxgfvN0D8IEthx4
ysg2X9skg66w12lxN6P+L37AWTU6fhiMfK5eJCBGG8Y110ULuilql54KY+T6
riInOXXJWbzdbnvhCukeuB9dloyuy+0mtDm7kSw3QtNAUMlakoPId3qACEFH
Rk1EQUCP/j75NleGHVFxLJKeNXuuYhqiWjzadTif+WkKNkeLmX+j7uQBHM3E
1+kS7F+bbXipWgChA/bOLQVUXsnVptx2Hf/14RzQ+Dk4NNpsS+ZhPpQqlmtJ
DEHUPmDoLkwYwJ5dL+H3I2viIffMpxrp1c1kpj5IVyF/oBi8p1yV7FATkwen
u/AkMHbNRJQXaBWnmMolYlhWLZCqaBsRCRd3u6ITK++PxfX8SU2/bIjEm+VG
SCbznbXepGry/sdgiK7gjFjwmsTPScVFfEAdWbdVt34wC7hKlWFjWQx0Colu
NWi3wmu3eb8FvAvrx+XzyPjDMkZzcZhWbJUHclhFzW6+Ys68D6fs/qqbsZJS
6ti+C0+j4MAtZd8FmzREWIZUVEVsVDnxssE8CBeGTJSBRsicnma20G79giCo
LGPtbGRQ1m12bJhF2zTeXEf0sU8x1Pyjfm5o8/O6QVZSFv45PGE0BRSFl2a7
ossgvT6xuqAWOyWong5HpL+bANK2i1H4pamlILE8frYpPuFVi/nfCDgAmRVl
MnQeoBPcJWRb9/jCw+qYsSj+ooLxY6PSAgmkLSmoWfbS0rbSYwxPyAxi2x/9
wr02MyBfuTvFVI5DNHwim7lYk2tWOQ2vMfw/0kZNs9eEeMCWu2XGr5ha9ZEJ
+nN5eCvpw+vKDTjvc8vBUDXgUqobbuB4mPDzPDY8NKX3XlIVV9pFgjyALMvK
vd5v8f2iQVHnXYLb2VW4hniCnP+2ta1EPlLjOYpXYAZt2a7mQzDpgCGr25Yh
WKar14mB9tN9bHfKUYNNyEt3IoMK++FwYKX+UaoShms1f9NdSs1CAgBZZpTC
hU8p1qwIik/9c3E3yWBMadaENAJ5M78xl+08HODoZfdnLhK7gAAPQe5rAr+e
wmfDuos3LWPt8n2S4F3b8vPOs5KQDkrMuO2+LfWqOWFZX5TILsqLf9bVVlta
8fbIZr0iNmD1WZLviyPueHNQyaGrIepczgaNVz5zdwoscfY/r1OG4cs+u1MH
wuCm7XISjsZKUrlwx43LT+jPz+Fv+6z70Ew+nPGpLIgq5puO7R3oKUgb8f/7
6wpfXsmN/Og/IL4OkuS2rreIUkZTjFPq+AeCL8JRrBBkKkilMGcypVmlrd0l
NsAp0bIGYbcOeyOhjQ/qxoW+RDO9b4tHv7lUkamIZIctVNOk+kyneUEEWO7N
l7c3tLfRng88dw3iDdTaL42Pjr+ASVpZ+ouhWxwdc/A5P/cO5X0b+vCxEE2E
2L3bif5aIxb23ovKPmIk0Cu9mymWvJjho18sEK09dEWJU9aVJb9qiv/rL37e
U3otQCFF3NOF13q+/yYE4zTMz1vmccC9sXjbnD4q1J3Jz0l2kRuT6c2/o7b/
sJaB/2+5I6CB2bKp31JYLdZ2lX7BeAQ+0rGBtoUcz4aniVyJXSyNJYRpP2Eq
4Nxs/eeQQiACHINeIBgXUGkh9dbfxGBla/gSP4R2o6P9sCXBRfrn6Ct+KjI9
XBFch22Qyccefl/pKTh9P/s8wyjbL4xQt1Lvx5KpS4kD26Rh8ixDlb9mHo7L
qS6gV+ccvBrvs5tkbG2JvIvc0tzSTE5ZrvWs66e32/UGKsTZnumbzvtA8Gjd
5qsif094Q45dyFYhTxXtvY6wpBLwxHYAuc8e82LvQL2wqXSPthn2k2h9/FMF
vIbwD9XX8Fi9iOsj63rqWrPpaeK9SehBCtBZLAbYfuj9MdlFB+5i41FvYF/0
jxsSHeBgvzrynfgqZ0nfjP5meY/jxhpKvBDrsOq0JN+UTG2tqUIk1tgjHeDv
exzK0xu7OM02CrSCxcFa57Xpc0s/NFjaKs3W1twzfLGWRX6U4gmkuzA6yOTn
G0VIhP3sex3kxneL4DsS/dIqE4meD3mM2ZitsFiLJuXNLZl8YcZfHlWljhqd
oVvXwPwD+YnLzbm8OxGtWc14pM+/oAFPg+7wDC3pUuzbiNSFIlhi3te6gCSc
+XtTTUy8O+85YNLyYfO7kOM+I/Hku5QrCZCkElfRgKBaApyk568AZuLWhj4N
djPJkJNXYjB0yxkg9lQkZlH2qpC8XKAGotPXH8K+5vFJvbDIB0EddHlULjFY
eGlGGsnwYsJHSr4vfWOdJAzd8BbbQBik6hYUsBp0V1xY1igQnTCf4ShaMzI9
I1nY/nbxX0rSbmOAlVJ1XQoSu0n37DN9rgKi3RN0zvwT1TdJBxOqn574i+N+
79Uw6MvQQR8Hw10UfCCkWH8BdB49oaiIGSVtKtoAYBqVreOKxDoTS00fZA67
Rakcx2oiuX93wMq45wUTHGj8ts+D3FzTT+PYG17nL5rhyDR24xsTOLvQLGjA
2YTkY4Dj9lB/P1nIHPt5WB7TyQ/Pyo+tk3KGesNucZeY4+mjiMzMPkQv0YoN
S4S6tPjlj9002hT7w8D8KZ+2Dw14ZaYFI0ax7D/jVxfHM/M3uVDikTbieXA6
JGJGpeFbvSeXRfIDwZVnugB+scqOvfjXmhPV/iWuf7UtzooobiEgZfttlee8
Yh+hi6bPAcuMYhBzdSAEVz8kS8R22x6XdgxfMEalyjRPi1T5RX49tuGuIvw+
9G/DAwgiSap/jeCTD27TZzDCctGnn3l0Wt8BVShB+waMkFTAjoQmDXAU6V75
QL6IHRratYkpya0NqzVy6ghLzEmbF+DhfXHw8vMaIgyNp28dIohMt9YxVNDP
WQFvvfVs/pw7BhSjyW+SUguSKwXZ/T6cxBEZGCJFTrZ53FOs7Co4se/KTJNN
Bv9TQ741bEHeX7Elqaa9A3ETZxQLZOL3vREG6YpGPSqSxno0H13/23PEiFHB
iNoNhW+jw3FbtJPevB+8HIr70l2aJY99w2jRDs5GkDZG3ctPVawGhKbAec3c
cSo60Tm4sG6ap4TlQriKxZdVS891cYrxa3ujqEEmZSvc3NYUJTUd08yN+aX6
yZgzGV3l24RqzCuc9WtarYZpK92iyQe6FJH0XxBqwb5i9DBYrI05mZlPImKg
TY5jWu3C83rBv21QJee8KLJ2e/Lf2aifJef9BTKvzpOSo8T3jx+lrRABxnH4
lMItjtabgaB3+YDp2Wug+1A3lbjdxVFUlkP4oWoLwZmuM4mog73wgfrvLiug
t2+2DC6avtYeM5HGQPuJVs+YdSJEpdOUYBEH/9mCMc2j8ViQB5feq1igmaoS
8Giq055zN/oMCZvLg77XtQyP9MZS/WtJx0mOhMmck7oHy0KXW0OrchXczyD8
pwcUrc7yWcCDheL9cOfXJInonEK+35LLYV56VLQDa3deKjDiwNqLDsw2RxGG
tz8A1TO1amAp3yWvSWvuqOT6kbOextXyZqcjsOFmSsrPWaiVCeoYHDIJZhQF
eT3Qp/Kt1XIEiLVN7R9f8osUPXWTA5L/htQFHO3neQtxyN+EbrieZ0w2Ufnp
HnK2esGnqD5AVO0cCXKcAKrY5ebf0tfWCaiBfMlC9CrgBlFfDxnp20wB93iW
iehAoCyoZdlqfK26sPtLYe0XVLnEVR5EJjchwfZ4ENn1/MVDFYp3fpN8hHdZ
dc3Sd58FqZunDvFHjXGqg1V3Hk202D9JaPNpb/sjh/mdU9c84eLkrQ8G9j53
3Ju3bDAwg6GkRzjVg+UwFDXGw8Ld4Bd2cGgkWO8+0PiUr2Tz53Vi4oTa7G87
P+eUu4NdOZF87Jpg59b299IvU6WNYa0J+zEHJnbTl/32FmLVvvwX5P61YwMT
61JV1q2InZBDXYT6NtJQEyA9Leso0zu6jh+zwmU7Jxs2WUXtl7vbxMieEsrm
dB/fYul/1Z37/yrJ90GrWnDeFrNIKa1W3dAMqcJdwdirl/WDVHBmI2u4yoav
22OKRy4JbT+fVN2qUZ/W9AMDsFghfc/l4p6sRKZWixl3JjzOiGV1HwTQqXpc
DI87VLXLvCBe6wwIR6XcyTVPuKRp/1tot6Wt9n4jEAMy5YrZahYniglzSLkE
HZGW8pIu5pvrBEXy7BwIhJxz2GFz7npZCkNtOn2+o1uo/bV411s/y38dL0z+
nHpdcbNj9x9ZueQNfsh64zkNLwcr8LgMbtcZAzKoW+RuXv6iph6PVCCGIk3i
eIFYLniad0/uchU7fE0H/FcLJ5Prfveu3lN5IJfP1yhwBePkifzK0ZMae6Q3
JdwKbl7YxBQ4BSaF4rh9Gso/C0tgNIxAdivPXgEvDIFrx04krywqsd8VIF+4
49UBLLpSo/CjSl/ev+hmy+6zlxxxdf4KD7e/08A3rhJevKNzNxp1MbJcHz64
dVJaKybc15+k/fEfepXiWqExqqaRRlw5xpW5esuANjsy4HKIpOzg770UxE0f
2CO+gKic9WQbVyI7I4UFYVI9GjxeRHpG6rPY5/okxSlR1v5eTr9ghu/MRAG3
BiFnmXvsN5Zm3qA88tGgOjTsJZKYaCKtzpIdtSS03RLaJSru2fMd70Q5YDTd
rTYfQgg+6amcIzKLMtkuFxZUPB6ncutBbC+jcmDJitPcUdPj18zNrGhDpmcX
NQ/M719tsnBfyNac4JNcEaK4s6khM6hgeOOVBB9J4FTXyjPikwLtyjmoagXx
PXAyUglQkzyxf/babxn1/o9PGZmdJsp7YFIjWIm/9wlg8OByOpwi37LUmrTW
/wIq1vPLou4UGmAXepXASqAJcaDk4svGXeSK7eOfk32t0vk9G0zrzowvq1qw
/0HiFXzLEHQxKt6i6CVD0LJov49JP+e/cOAjx/gUw2CytIBjBzNiFiPB2bu1
kcKpOhYAfj554CdS6+fBP3t2lYI4/N6NFZEwtzl34aSurWVDKix7Y4IPWcub
nXt/kHLLM2dS3T+CZr8L2/66JuQsbxv1rRts5LYu3xBEW6iN0UMyCxKF04ye
2sYWTQ/+1tscEJ/3mv76xTu9nytsgO2p+DMzvt8yBLgI5x90WTpA76gLhS4A
evbm+OajCyGMWbMS1q35iXjBhAfKXJwT/NbeqLWoVeYyheNTKtlVcBkhH1iU
cJ/CRfKMbKDb4FOFlCtCJ5l4xHYbtjtOMfK4D/Nrwf5dgcau8jJ9x94Ml5H7
VfPw+VA580edQl81VOXFDO7Uny3CqjVQDkTJc3AiopvV/IlcQlAyqm4UbHpn
7Ce1BE70PWPFWFEVZ9F+ev/nbL/2z4DmWvQNCPn3Jw61dioSWNInqpQjmo1R
5T8RVlJffLq5FbIMKd5HKnqKDH6I/FRPc/0QDE+bQRzHaf518Jb6d/n5wTlj
mfWfOSSv3Aguzbw65Wr4k/sQEfPeA/F/VXGWvcYcoHFlV7Sz2HzWYhlZ9/nq
yfM4cJLA2kIXfMIzuocr2DtX+grlRLcxOWHK64OYlpKMgsefXqDl4WfpVpwd
5W8BHDAV2Itq4O2Y6N0idtSu0/AHXEVgUh53SfkjdWUxfIwF/LgROxd5yVGS
568v64S+i92bLXVnnKhDpQkFaXNARxVoE2H/ybpqQ6//F41UvKoH/9EQl1wN
PsUCQv1Fv4QNfdXUiSPD9hOrM7BVFyMEh/Y+rzNAxog1CknJZEw8JyWl6WJe
c1LQaVdDznWSv1ehDZp509KHLuf/FMGB0Mj8hAQc1SSdBBiH9ytUfpsPBmLO
r7P2/b74rBmMrUBdSd1B6jVac6ZgtqYiDmAW0rrNOkJAaph2QYU8y4DlCVL0
7HknRfV5d6PKqKhmAT/ZBgGVTn49agbLua0shA3rRCIEO67UtuJ3jOiTPDze
VAvCVPv8yUvMPwk1ohs/J4cskfd5cvGyIg8pp99VgZ813Xo6LT2lJx3WtxQE
vrUnZxumu8Eo/vVKsf+Tav4oREdPt/czVGYcMymq2YJDVrBXCCBP4OOSHhAy
JZCaD051jxrVnbyEaolcjerhDOQcVHnkqVXmHk2dbtB6lk/+BbHM8Lcdjq9P
YoB4JSS/OWtXxKXozwWNN8a4J58rSjxEv5eOI73e6Zepa+jRRvuyCjrg5iZA
6tHaX4++J0I41k2r5g/rmxs9uwjjBrDWsblFRAXx+34P833ZlZyaGgqycEvF
QLO3kJBj3mltzmEVufpSH82tyiHuBtM6W3V1FmlWE2eegLC7GCwohE9Yv2dA
tsg04zCg+vuzhW/uduEyG1kUNWG7t43pV16XEnk0wHrxSjio75ZDxfDEXVWE
t/2i7joA0UzL+XIgZl99PdpjBob0FrtHcbsba0HenGBI7v/CeRNMFZYMujQc
jbf0sZGBC4uN+UvTeKVbpMST3tkqondxumEp9WjPLv6ppZqgnFDM7sKC1wbq
rQ7oROZMDOdi1W0I3u0M4GU8JcC4bYFMI034wXbOSrpcL4+kIEE3rnN77Bu5
34vAPrChrG4CrTCoOpjShQc70GNCcKqs/mtnRxegEGSVZg1fZmrfUmBDKwhp
mC9yYyXDTghmBMEIsQAipjxObBt8yYZaVkFn1PcE0bcFJdpAj1siSuFGj50J
Gw+6BVjSBo3Hw+wesiE6+05yBxF2NvY4Si7zGCo3MIdBK8xWSkfHcImR4qPf
T4m78r1klNwBXWiKaV65ETznqOz82rEJj/t5eYiXjVahgwlASXVn32YyeZh1
yR8ZXxX2YqOLHBAAkv2WiCr5K4JvDsTSwYSSy5U+3FYjjaIW9BPXYCnSSRv6
zWVZTuulhB/2qHMh1JxaHlsOX9mkOAdH3hnLBHmfMWsjawRwWeh1CwnSK0Ja
lxtyV2V9KRVk0bllxIVLdhMMWhmp7OrTz6WlfCYVmt+Manxa8vLKBfaHd67I
+DiQdCKaP9wq0kqG7YeD+E30+MHz9OfqxPmPbhem94t+wSrMqsXy3/nHY0bv
g8IlxQ7ijBqrzo2zS84J5RMI5Zs4PtjXncSQ9iEcNvhMPmGsPzyOFbvk944x
ueq/xCcT+F82wssEB73J9zvGqJacMNSTgnhKPmFUKpV4Tg6p3MmocJLDId3B
s3i4uOmWKI7GH+5LHjKQyZ79XWplqW8pJOSi4c6FcMZgAeI4vV+XfnkXHbST
kCGM5ZG3Hc6fQWKo8YUC3fzsPRH37nDkLpSMheNLFEoJ4Nt0JvlE5RzHRCx8
duSFxXd8Fu2t5Mgy3AzRyTxqt7e+FgCz0bEkuaSp7bMYNYI0SGhHLAOrT4ob
DjOSnoLMqdkVvmBI2s8ZTydUdW5DOV5uVOtclWeHW2g26CgEA7wvfNKNhWa3
6j37nA601KTZtVl5z+b74w1CDsnHn7PzRWdGxe7YnWtFbeYFADRtoiSiBN2I
sjvbkMVc9iE1Ta9ay4MUOWv73i3ym7BQ4r6Fm2zrrJu5LkdGVqxhU9zcKKrl
C1zWn+ur+qmr2Hymw/3uF7aAJKBsdVxyXb3Fh4oFECt5AE7JqAqoBwW/eNfV
GncEfYNtxPm9AP9UGxOjzs1jWWEpWSKG+Z8zUFlmf3VtPGl+Ji/enA+GsKtV
3qscn0eEX/tbh4HOSLplLfHlPwNRL0pAUr1/5OXDkmsv4omCt3/OIxzLwJIJ
DPEqNG0D802NW4Pwxc79TAa7PkgbH9G+MMgE1m36kf28OOmFVg6vc8itXd9M
U4RWZhMbnXtlFo4vlNee5JczLgeuYGNdW/TuUR3hN3+VaLP40rGUKYcew+vf
TuS42tMpe3fJvRHSb8d+ZUGoPUph7y4uisdzdi1uugYCEcHhzwuwKh2Hi486
6TMBiqH6Sr452oH0tDShUEWE3WeMUBIDlU8NVK5S3p2LJ39mhEggDg0vVGD5
6USXbQp71nmfv5qLZghKMVKiXOw+9ssWh7V/NfxVeaqCEB67aRbyAJjCLOBV
gWU7K5tFIJ+DuQqfG7JMS1C1nT8SGTPiwWZZLu39I0x9Wfqog01uDCJyC6QC
y6NaoHunIiLWCi/mwjjVIrxDMMSN2xhJEL0fOU2T8sKxVoOLJMdPeDPUq033
e5rooru7aGPwFmbYiQSnBSxPm/dOowdNcjSOUJqpgOZKVazGdixbOnl7Ec2D
T2IwC9YOxCNZQdmEAPswH0a6PNqFNfjAIYO6yCxbUDG0aCnKwWr2h039aj6x
MnQv/YUCtdr6KA/cMHH3QFdUpx/GKFY5ca2qfErGjevky9B9AA5Xl8EtnxVc
y/5nNWRtbMsKGUbwznLfyoxCI1i3nkb5sw2QLDGOCMd6Z/1txBa0DoKZxfFY
p+CqrEEMyrLjeh4c7bKkaPpum77Ujm6oFSXlX1+5n+kc8HEyKs239+GAcGdu
mKfoPvYFNxo8XurEu2Y4QCJAUAN1rDss5PR95ojb2OxxeRZkbtKCq2cRk7jg
FL+4AHgK/xeUV++L15mjtR5v/xAf+yVOIXVnrcfCY8d3U6fT9eJxClv8rJGX
wuQA8vEc1TGWxSWVn7nnVvqAYSTF3M+f2GFgf+dBvOg9I4wxb+uC4jn7FGij
kFPKKXGvM2S5kRnxHemDjBnTEoueMALc3cfsYvKUvdHBn0CD/0VggQaWiOSF
kn2RSfA0gtCXEm/VC08IW/IL+xTiUXeJDMXEzR3osmG+bhvdxdZVqNIsEDZq
k3rA7/cKfqMXemmfsICjGmt/zCCnss63jSoXvKwA1+2Bh1Cuh/37NhslAymd
03jdHQqCPtTIdhsa6zENGLog2yMxlOxYAjhK4GNtlwgMULH/mxj0cc1yp4qY
Zs9fr9PGdA1tM3MGAQ+B1eJZOPCD92wdRlko1OWsL4xbSkzwfk4s/yMej6/k
kyf7709OeOLOhMxVL7QDJwYa9tDTH6aP/v/OUP+tzqzfTkdpzrGAsO17bTL/
l3ux4+5tnMRj8Fw5l5eYfON3/lL7f8haMn1NUKakdwojbmGq94v3G1YxacgG
pXjcqGHPAFYxiqfVN3puSKaLH9PUCRiBtvyBl5+ySFtSuwUH+xa2CJwRzIKN
F6XmFZGToDKUq+FNYxNeAF/plfQo5gxfMogcorYJdRbK9x0EQBXOiigGmZKi
9rk0o/GbLe6pssXHN1pG/JfKYJfUfjRRqfRi+u0w/xlQLHbq/qO6h5aQDZwH
5l+fW44nyq3WjBuXExh13S307NQb24pfm4RAy+AfaNFpVJWvIqYyWJ0KssbZ
+Y4ByvBBfJDrLgGK/kyFKzoHBbJgx8vpU2iEDU4TaS8+UWOTKBhd4VferSjX
JyQrVb0ahzlHN3JUNS0eLbXZxRcVt4K0lsmHuGTBZwcRSZVR2oqqdydFJZB5
PepioVxiCgJEbpDKOsrde8y9By8psimnzFI964gqGgPRVDEgKI5QSJMoe/0/
kzq+cMmUhIQ0psUJ2MC7KXXo3rzKCATd0olyTOywkVwVzjp/JpRuc6XAUsLC
QOFBI26X2pt4Kvz9Nk+CpdSKZ9dRsZsDlBxvlxWNsPm2akw7GAvNmGz4d8FJ
nlQgLWTQTSDYeL3/0VWjh54rldxiJ1ZOOYSSM4xC5ZeOUoZ9ewQY9U+l/CTX
HKYmHwOVbngc9Qlb90dfSt3oQm9FPZ6iX1e+QSRwCnkryyewE2hzY61RpIjG
PLsbYNLNLoQ1vKqhJCMuSbOaCreeA2qn5jLX118X/iH0E84t/srj0eQr1nM9
29KCXrQTl66lDT0Z6C3vlB+4ae+51/MKyIuM2oLqI22Z3DPBp2IZKrHm9Ctx
Dwv+1WGKoYDAM/UyjpE+q8vtCH+KNA5T1JccN4Hcfkg2Js6LMUtNMu3TK9rw
5CG2jtg7sgnauDk6MCflOrMKCBBZ704yw2PAwzlyX9Tl3QjywXYTFTXPRUhm
+AvvzYhrTayPvacHuvuG4qlMYccRows6Du9G2hhRjF9lCpRyYfVqXtSrw5ff
vGeVOVljq4+k8XmVRE8hahwsPR7bHb3o8gu8CgGy0ounuLbfPRewL+uow1vK
orsWShKg3dDOC+4DUgUV69uiD10Shv2NNLwmMRFNBBtx46rEYVJH9ml/l1KH
85SftCeN49VfBpkdzrZ/6H9+SQBL5STmY2UNI7fAOfZNj+PPaj+HX3hxq/Wx
9EJ7Ma/su2FSHnHNvdzIMJ1K4GQRXJneljbQihFuvPlIJq/D5ZSrG6uHaFW1
E8qkuAc++KNE8d/MbEYhJCxZ7hDKGQNDdl5FyBi2Jj5ScWnnCJfuXdXppK3o
PP6lCydaP0K8FN7vD1InYbUFUMUxoqA6ve7ZOeKOHfNbyQaaGQfuUGjimdag
1PoFO1z7Z8otiXADjDA1FWi4GV+F1Vs7BuG9hlnpPBNe0EA+hKS1B2SoEpY+
QzepO3atBClK1zJx3teAd+801IZ/74WnKN2sqV+LB2PkuuK8spVLf93SUwdI
YI/BBT9Rj7wQ/3ea/0i/FQcairS3jlUemNDk9cXe/z+sYLsjOcKtz9y1Fjrw
aNpLaOlRTycc2BMMcUfQmM4ioRMpPCTNf+aMGNtI+jjGyXJdvW0hP5XzQ8ZT
0nALHFj/ZUmo29go1gqR6YUj2TVdrOWsnYxtjqTcL2jKfcAKYWHowUnVuhtZ
ZUAdqswcJSprhbdYjtgEeRYQUctyJqPI6u48lrU7P65oMCyLCEzH4NmavvDP
6NZGNOD5Mrc1VzzVHoantZCo/4ydtSVOatOezsd2Miy1+wCaRyWqkuzEfkbL
lKiqHPfGulWFSlKeYMOTa5POoSb28z1FG5sPa1LYNNsepQ0C2t9zgQG6Aq0k
vz/dDsoHKy67ZaHzEqfQMadL9zxEBD+gUI0s7vyOTV3l9nADktuRT+p7lV2j
9WmWJNFmizbsZDxSWT7mtG6buW+qt8MBRisBSilgWAAH64uA5Ia3fGJHF/BC
gTXpiL7NPd4H2spmId0Zn/zTnTtDypGogMQOI9sxepPchAOjn8BCy/IxsTiv
fcA+Xzb7ghHv1qxHBnx5K0TYgoNGyg7o7SDngCxgPwD8tJKLYO0bO7PGA+FS
K2b9XcrXtBwfa2UvFgvkyFMHrMqchsb4yVRMnnY6H795m0sT8MLpAsqa3FXB
lZhQFv91brFLgl+SB43ehXk8A+DUuGH6OtrTOEqfuQt46EAf5PIl7jOlUlLd
15tc/ABBi9rjqd63gRjQYihoCxWlL6AMuXt5X6mG6ftrdETjJYSXVCze+oL/
GSRrRDG6rqaeY07j/BEp5zDSfdkzRQ8e9KCz3QU8WAex2FOCDokxkcZmrxSz
SIhMiac2fJHOZxMH/PjwkqYYRQABz6+CWCquf+nE1z/vpHq/kqTMnx62n+YG
w/7sNPAI2yN3mHgQ0Bt19EefbYbqzSOEeOD5neVecj6jHpGiZ+WXOiDNx3w4
i6JPolOHLrV5LUax30lMJ7ECVem57C1RIQN4RWB39pxhBUR1DRp/D53Du5eN
2tAmRg5nem0+ylgq0X11DW1OyckphZ8iGpSgChhLPZkE429medsEwMmV/rCC
bwtg7xoH4b2TL9nd1942xiCBoxzzumjcOKqRL82dhRVEUMhjIXZ7ht7jgy3p
01nLstZ0r92ztT0xQZkJ907Zpw4KLLt2iy21EMjKIeHbGr7/j1bqZB922rVf
MpVY6KbUDyd3MRWldgzzUdiMNuZsz3Al8M+CVdFJR8dMOx9OjMcmYY/ZcS6S
dr6oQ7jlxmvI/rBDFcIY6LlJE7huh4/xkBa7SwLa41qTrbTiafhTCEPE5KUS
egSLHlZLOa9N2qdN2VeguocRvWByhQG90QGgXRFQiVFVquTca88Z7L31aXUp
ZhPK2NEFOc1r0lt3RfsPk0T5ozs8wro8DkOC5yZoXmXE2thyLylrkESStvAg
8sFmgpNxpAQntfWDuKolMUKgb8qkFO9H91+ICB67243SJdDsWyAWJU5JWQmr
D02Ta4bS2xyp+8zckNq8PnpmIwp0po6k1dDRMw4OMVwu4TsKpGivjaNpMTBk
HWxnI5AjD/gm2jT+Mj3R4BZonOi0gz0sXTaK1Pr3Rfg8y0VPSvy4fbR2Hnv9
z+IlV4JgcfciOIlB3PtqtHBMXQNrvHQ4g7haYgYnrNoPlkg6e9HrufnvwK2T
JNODh8VqYHfa1X3FPW48pfC65qVcFY90Y8ELWqSmCpXged2ISnJADcLCiamd
NPA/3QPoORI1EYfNQfM9dUDf9pRi28CfxHLghzpSQvByR2ObTd1kWyrYa9pc
l8VNl8iYbVEq0aBqH7TBwZBcvBjTJhlGlwKXeVak9bFa4+YcbqrW9/M9sJKr
JlSlrIJnSTaFmrn8O9p8SBeR5q63uOYPpxd2b4lSjCG0eW7uVIUoJ6ZCF8RW
yEuJs4/jKlB/h1QYwAk2iCAcCJ1AAyv5h1bNfSCIusvfhE9RwUQPwRpD1/HK
b7XzEImYF6FZzPrFn1irEg8cyQ6t9cGDZ0XOsihB2Jf+cUmjlWwo7JEJ0v2t
H/tmiSv29bMnoHnU7M3YM2jfjj6lQbHTLdCjFLAHXBWQ7KddxT0QCKUWsoIf
dmoxHhsDIBU9DKSoRBLHfiG/HcaslxV+gNXBd9wgGSqCdzilGHlbedGg6EeR
+GYJ1lF8PrkK8APFTKqgjhh9M122ZkkItxvX2vgaOw3FdDRBw01lynKHWOuP
f53BKTvqxIrwdre23m1SP+7y4Xwjum8QrN+8x4bwjZ+S0j1uvcDne3YCLtDP
oc+5g5Jqq2BaiZvWtlPMz7RGOLrCX7EBe8+ibgdhGZEWPYjRodn31S8EIxC8
73loId0w8J/9JCK6BsQmzLl23xQqRcnv+umKIa2TG1uPUE6k2i+fgRjFlwIg
WQ1xnXti6QezAIcqbnh9iW+CDLojBb4XvxV7gH1doELnIn81S/RkQtieF8C9
eGoddyoM3w7VbFIgJOMwghRW42GBQzAzJ2SEBSQccqT1mP/JSdSwyGGHsANw
8N+T5l1aCPSpJnJaZDbG4EQmfv//+ACAtMH9vrgHxLeTAC+QLGrCrJAl7lNj
M5DRDaZ2mkqk4pCXMYejSYNclauX7SgtGpT3ixqKyq5meQIuth3D12kDAKyI
Dk10d3Jr4garolpoXn9eCgEMl9j7HqG7mE0Y1S+Tmuq4TAA0m2FjHaIfVId2
ETu82KVUe/P3RAYOBhLGBug93x0uZCTs2YReKcXYlcnQCrGrjr+W767bd0R9
zfx1Ih/hD7+QjsfD8oDfIWvX+UtNTHYruTf1HvbTld/hgMrCYgPifjsTJqOh
kOD/XJPbUEAMQG0IG4pFejrVx1Nwht4Tl7P/wsuQquQJNkD1GPsVpJWnlGMY
yZa9U3uPEpxMhVZY1X8Qi7QsyDU8sf3toQmlPnZeMfO/jMQL3rGx3ddEX7xS
8GE9cn83l6ff7pZUP3Rojdn3O98e2cdUMnx1MQU+DQFNZhtqPRkFHdFo2Q3Z
smi7WEeEh9BBVsb19pK+e9mTIpJZOnMTeNgitYFplmPIBZXidfgxqhETsC2C
Nt7pr4rgWj7AH2HJ/hEXNoQPLxirWJC5mlMjR7ru79K6LD607anOH7jVZ1em
0FUsjadW6qQonUBlOXz6w/8n+nw53yRHFgUAd6/9WnQOCJXnxdeG+5XcWKMO
AMqFcTUN82mt7faWXbI+/IUMqEOhasOq9kyZQ9EyyyaK7hjpSMLuixKUJKJS
XnmguXadvJIsY5qPzWrgw5eWmjzkPSQJ40QU1zp4q4U/XFNe4PVlm65egaXE
3pKvzAnNcYuTvgW7WYt/C8VkjXBQZfMX4VVJZkwOV/Erc4eFTH0JxC438QUO
cBrnYBWk679F9FswwvOPH0h6vrq5s+wAkzfDDTcJf9m9vaDQY++XQVpy2DSF
bWeSITuZl83M01ooV+l2bokYbWYx80tcoAf++P/mzoITPyQEiQ5jZC1FukCN
oJNbphs+aScF/d+tcdI2AVOIgSaMRw0jopmYMHuoxqPZIldqvmyl0FiEHgzP
YeY3GfQ20TeOJM0ghDSmwe4FwpPOjpADN2TVfTmbVSHuetqPfc01PN/9nj6N
FZLdPNfgcHZIDESdDC7EXRagJMqja33/62yQ6ag9qQUPeIASGmpy24EpIg11
jiZ3QMdmFEFyBx/+LZdGlI++cbcsyPBTSXp/AO9+RAWwM4Y1+/Nq1v36ZtFA
77F83CVRYnXC1fXRbi1t5P/cH8ommF6AOmVEWCzTmgPTS5zl9pSuXo0WR54R
5xeoLgGvessvtqKcV/ilt1kozLrldNbYqZdf2q0FPcQqW+PhYJZRQwYrR9Cp
4K+lmOBeOL/fDsTflY0x8ENeLFsztn7w7vme4lB5DrK5u/z4cjUy7HrqqR5l
W7C7q/7+zxf+usG8ZseD4jAT/KlAJMejPZMGHiwkg3gozECAdDyUC6sb7hnG
JRaW2IVKTYCeSA32EuHvhvGpiA8LTXrlwtRJl3B/iEjx0T+vIo1H2EOX+L9Y
T9QbqYDuAKQJz0y6kbKAIRqD/jNrApgVn/THCZ1mir783+q9kufimBYC63Tr
/xkIO5Mwt7NIhNdNfvJg+So4JW8jZzU/I8FM/xK2qK9pqUDwtYpKe6l0MJNY
K8jm9zmlzQIW7wV3oeYYgl3oOYenX3FqLHFOc1shKZkKe2ZU66drtV20z2Eh
F+2PFH736ws3No9/IoRAOdoqEZHnyED61fCVn/eDeQC4rtjMUKmUj3b+m6Lq
yaS1NLlsLyNCbLUTitNeydmp5d/FlV8D34JD7gNuMn83lxfVbBK0vAmWrZpY
sBqD/xAD11ORBw+DMTJ+3jbqQR7U5KIWPqqFchnJGtCe8IarGiCP7hLfd3uM
SIfEI+S9PeUV1Eugzy3dD/e0GlKg2W9xNAUB93++1fd2JrPWcTL1L008Pt2F
FcjRa3P/+/0tNSnNm7n2Ln21u1VGl/1HTxDUPwdLhijMn0b+qc2XaDY/5zKM
qgyGP1DzeravoZYi6AtgiF+N4PElIk/8nnoBUpq0mzBouOOkCMJHrHi6kOs3
VXZBuOXpw35Gl389MOItvWP++1PiKFeynQ1drXBko/I7AqDHGtlrBDfQSJzZ
6fH2AJXDoMSWNqX9g/lqcRFrLRUb6OEST5nZfyutFujKB5Q8X8G9MvMegThr
1gnR+9CcNWe9mvbqZ04Nw774n9c4ni5xYFIv3QYH7oIIQWclUy62KlAUR/j6
G/KsQAoWdFNo9dZMueKSAU9B5BMb7YaqId5gMjHveUe4Cc3VA/LX2cbKg5Om
eGhHC/FYUNmF5UJN9YebVkAYyt6ScWM9fiElaY9ZKPtUHlUS2t+JNMFv+RHg
Yauo6AzDVpYt57OmEUszzUF9isjJX9+NKic7JbbLqP7ina3liR2jkMYuwVif
mu4y4qEroiw8JWHEdgRItO7bDJXKwH0kn1Fd3zl/QM+Ej34YH1kvHbeVpt57
groGsgnvY4m57CfFgDOXzixNO87EG4wxzQ7FnFy4uQDeLjItD/Wffa55mO/v
UtwJuov69QWxTT9iXjWNSR/OlkZqS7oT+Ym32FyGsfA19tgfQxJYa2qmPqoN
Y4tA9EKYc3M/1pF2GYISoZ+YgTXhpkYJdjcGpNLUBw5+ZbMYY/NzZfSie6xl
j92JKED9XHYtxJwhVhDUGKe3XcoJAauVSd7doOuSNT6Mu/aRX8RwBoZAcJwd
Jk/oWa8YL4URriEfvsMRjrVGhEStIm4JX6H411prTn0KjOsB6MbWrAYpVUhf
rDgDRZ5ukob0WkwEODPyABU/pOQfCvXs0BH2N6qQ5mQkyl1nQTNYN2alzT1k
C/ohesgqhkufxzXOzIxtAVHVuKb0Vr9605vchDfbWROcRx1a08HHAmfTCWKi
46YxwDd2JsF+z3mXq35+KPCFIQH9AsgbIA843kHacWivtGa29SrmbeXuC+QJ
OFXFr1UPwVjiEYfs6q4Pttq49FJx0qiCvsM1hvl0Y2uvacT2vb6503l0wz75
128rM5fR/Fd8RQxEPuBbj8GaAS3P34AvQYDCKjpeyHePSWZw752+nkveFCfH
fkQivaehDK4AoQU18ZkQv9nDStdn27ewpgV0fc9nl5y/CEsXbkPnJY8Uypvf
csciQ3a/CYcXGlxkRAkXoTn3zsOo1ObNwqMNMd8qxAukBpCwj8GJzOIHkyUc
TOa4SFGokE3+Ts9z1Z7mF7/sNvPQ+K2Dp/gVwBUgWMo66gW5Qmmz9OmNVTyG
6j91/4+r+mPefZBn20wTyZh4mrCfkr1ftHv7GEW3j/uV01VY3CSpoR4N9jFs
gMKe0oX0uobOgOIey2lCd8FVDHW+MpvL+UYZ1Sw9xMAP1OLATtL0m+FQrJNJ
zR7VgrrKTG0oXn57L6UnlC8z8cq5oxTd8e1bimyTkwz8k6xbiwwdL3nJfNuR
mWcRc8KSt4Q0cIkc0XY9bbg/KMTcKNAxUddWsximH1TVykAlmOGWkE913SHc
B2jzIMLQkABfGMhwLnfFS5OrKqAe9n9rYG0f+fB2j/vxNAG0YladIgR3GdxN
iviwCABqTe8I9PYyVOixydK5il4pXHYKtf7QxpF6qz62D/aYQAbGZZfyInTH
k1Yt+hT+Qb3m7PFN2kUA9NHZi288cARzk7ZqvMl4tlIKC97vCC58DZJI3ysQ
8wtIUdAuHzfM2srkmACzBDeAoJOOS4z+PP1KqYkwDrBdJxOAId2RCS108ADX
tQC9t6/Ah725egjfsp8pBzs0iNcTdRIGDznjxrdZcE6XzU0J1zknJGtE6mBx
zcIm4I9S4Lpw+UlodgGv5oyqOmlFjlrTdJ0aOdwakWeNmTr+3lhWAxmcQojf
NJTbpdj5XgdZ40oNTksqBbVNoaSgBJkpy0Ck4C4loeiWqWz00kFdQKz0hX3N
/YFX2/BqdMPStdNUd7olR3dWROyN1TL4UfA4flJOXvAFlp+N7piDOjWltEUj
kHho7A40Cd1CyN1HENQB7c018YkjXpFao4SVPtD5CreVv2Z7lXNepyyksb9L
Rs9uGQJaDkd1nHFP/gSpZZR/L5o620aI/lzLeLXP/9u4flW2JJQSKgZFATFc
90Kq+ATtPHv4JTXPSwI5ZnqOOMTp0OVmLYr0+UToNWvJQAUkz7JMwlD2qYeL
fjR7G+RH3Jyl5kTueXuMoO1E3GFHKTD8dd4P4T7BSjCi2mu/pOBC1EzdY5Fm
O12NCOME7f+oZw/KQ7JoH4Yh503utWInqrAYJt8/a7teaUmZ2XobW8HyNvZX
gDD/pRk32fhJb0BYUVKmNQclUHVKLDnfji9nJDZqSGLvmBBn46c/dWwHKxMF
TEmv0LhBhXXDsU66MX7VFPHt4IAATPl2eh1p2A0M7O31ZKgIIAZ1X7hgdU+J
8xROrymtFZZ94oKK4a4HWN23AIyABsLS5cHAD34Iih9xxRwPhKFHVaCMPVew
Bgn8y3RbCpQjuz0WUznSR3tJ3BZCVSYd8yHBXthzcn0VUXk3pjKt2hcI7PUU
LbsJZn5ZsYm5Sp0FLZ5lxhq6Fx9Fgr7ZpdgyNZDq0ai4C6uL/HOHA3y0XrNH
Y1oiarWKiFGFYWJ0nHtKDIyCHn8Z9AFRCqMMueXv5N/NJstsxAvswth5miRg
O6ocGVR2D686OLFD7t4QM77mX9/KKUW1nU1YGLKpBn3TJ0z8T8dX6T32n99F
6cifJBw+kI4OdhdsHNPpK71qtqaSklCSL0gmnM/t1osZRGRlzjCaUvWD5BHM
4y+B6PTXVEhXg6hrqLPsMpaX0VdCsiq0mL5TFjwy5GGrVKSRx/FPicI9yUUU
vprpxseUyjvi5xcG+hpuygbArtOsUTOrXQCfb0WAwOBkX/hcOZlPaiSzuMEg
2sCK9s3FFOZCh0QQVvre64qDLoQCtIyXAy7kmjINqHyjdHENXcP7QMkmHyqU
Np3kPpZjftq+buLbXu0T5hIufvkB0Ze3fZEfcySXaHybHZXul5vEg3sAxOuI
NQrke2uNebrhqK9sYJABOp3EzmKVQzByGOODvWQqysY15od1iq7XKqBhfaNg
TAUbQIYdHFbCMEV4PlGo5gImRstQ1nYIEwy+FjSJQ3ZWXScGlY8ZMWTu1gZW
WcAw4aqKFSPF+5JBGWZDneUcRg/PfCu/Y287aLtrArlRYoxnJlvIzhcR5yeO
3tVTzVVKEJMhTwOC1nbUw24FCsFW2+tx4HuPKdPxlDCrYCSrS/SDmQWIFkLe
TX5/BukKpB69cP9OoqrWFv5iXqm3xwmVFE8dgGHtTJmXlTJSda2/wEQk5nIV
uiKuuOl+1sv5e+5GePWqmrOLWPF+SBGlrt3P1QOab0+RsNvtQcvhvG716HCw
UFlEpo/uWsPD49eH7XxtdY3C5bV9jcnkO2zN71Fjh9jQK3QV1e19+bVco04j
+wwtGs+ER6mknvJw7Hn0NjVLizYx3wFVhn7PjDtpNCosdTr4FyzvbNAc0Otj
qlz5J0vSeSMEreAGN9HYO6zbHsIsVLW2JphQPZxq6vnEe4PxZbvTIT9oEXXS
jWyIg4QHJHlEQMO6Ye7WC3XSoh7TvNbcgXuCDsEVkC/9Rjx36yQUDYLHDVLH
yT7yrZFg3GmtM4BprO0hagyvm/75iHlgXsiQqY+1uzeWF1bKm6yuHmB1n5YM
bYn93ZeMiR12fhLPDxXeCyHSCjOHCGXs3jQAZ2y5BdtoZlpl5XE8NwtTM7zJ
EGf7Ugnt6QAXSj7JVcLELBYKPT2eHqOqqYjC9tZdhl3lOVXXZpzbCvdrsf4j
3SMsOHnEhQxwYEcACgR4W48GnNUXatkqzMBFQ2y2CwKloHnD+RAj4JextIYt
iAgWO8pfKrQ2QXgRbBowbgIvt3RTJAbsTuo1jHIYVGNiJ02hzdHtn97bdCLQ
IkxBGu9S4l4nGHs1ELjgmHJDAefYQ5yF4qV8fyqMWipblY5OUwCmc2pERmR8
gu2nXXehQP+1Z8kCApGP1xSS4HufyZ4glOY4uTF7NVlqYgfK9we1EjS1FyW3
ljGYQ5khMcHfnoktU9Sirv5qkAUMksh/mFlCSLoJ6WTak61rj1LCi6kR13PU
mmyL5GXDr3QK0hfOeM+LdPOs3M0alXUxkKb3uemmhUrC82WUUQVEumSZrYT/
pnhcpFlMrGlRYCHSo+4aCdMnQbz3HLwSH/BVcpH72zKM1BFHWGQI84Rq6mMS
gaYCc4yn8GkNcZ6SRd82Ic49+Bw4G3O/+etfcDT3lyUciZXm9CaCnvvlpSlN
PTa6Owlz/01IHm6ogYeV5sJ5wJd7m/oE4ibdddNTR2pVaiOpmx3L+0l8vq0N
roQ1+CTpNf4/KgsdafVeMBc2WSASiWENC+nNk5NjY9o8tdnKcqwCT2tD/pdq
0cpjVbIGNvn1fqfji7Alqpzm0rFE6Au8owGZQThgI4wrp9K8kwCQGTOSLMeF
fbNFGE614jKjjQBD6+oCI/VyLK/RC13cm4maeedYVZmGlqUEMPtsOjrND6CE
lPQPOiIN2I1/PIep47VbZnRcP1Qn1N/gtm3E7x7U5Iab4mJ/1A2cmhaFUkb+
XIODfuv1zurIyLRKhcx50LInL0PM1DC6cJrsR5IyMSKNfeNMy580BRbz8dh1
/p3NHeWsw+hXhP459wxVsYjz11xcsPFXkrRUoA8Wr5zAeQUXDpgpKOxGgawK
1O9NrSQEHPhWUez0KTNm8xHze6vOQ7mDDbrkAujbBzfYupzRT+NhwUm0u65i
lEakRctz32lpSPGK0L469Dlotu8Rqi0lxJbzW/zbbEFsPLw537jpTCLJQ1wR
jEdPP0+yQpdHAxgSX97gUwWJFYvtfKSB6cQHu8sjuWFqXkFab+upIEiG1knD
apGtPI8eJvl5hQ5DEAsxIo1+eEaxxGwZEoZgr0XdowrPzB9BhMlw22XhjqbS
4P0qEG6KyuZKqZ3TOaGRSpj+2Etz3PYzRRSM/nkfTR5yh10OhfSOkFDKD6iA
BYlK0FWhB3/V8JM1uXbrD6xLxfX9uaXIskKFRb5YXULf5dqEDTnjjNWlBsub
iXIIgkuM8JMQY73FE3QB3NsR2fxHo/G45eYR0LMoUA0MWIUbfGeUoqySW3vB
r63LzqHfiAEEwXKZVVN3BhsEz3TE/m2zrLG6eUnYGQ73bhYperC9XwJ6BV5K
SUFGab8BcvsYlOo5BeigAGL5YCEik2XyIzFRL2InoKUrNHzr/H3p4szkhq41
1bfYdvc/8eKq5M6aomgerEDeambcRiMTZSF2dh9qL8+PAD1c2f6gzwDhK1WI
omtldL2ondTHwo4b6Xj6ERGtlFiNJwlAG7IyERhZIKJafCYKOtLjTBpxpiDq
IkwCLbX9tuMzx2dJ9zZPVCRtiIcV7n81xIZoSY2P/xoVbo4oiu6kwG/EicEe
IWHXUUbdEcgodluggFwntiDO3t4Wzc45bS7sJYkZbCQLyUDN3o2FvgffKcY+
Tx5U9EF03M9t/KZkZ/Z6Kgp7rYMeLyWU2G7Om0ZXQCD6ydAet30GtNOmRKcp
2f5VoLpO4UfVbQsJF4Z1RwuGNkTBfRK33z/h8zzVpKcD6ueJQYLHckO0fNA/
sAyc0Yubx0zZ5WeipDiurhdj5fnyzAr9m+x6uHm4xbcD+Cm1JZTloYUkBPvW
3jUQksxbEjv4K/NCkcDkCaAZe0whUdtbY+hGEk8Yh2CsjZmfpyTOle8VuhaN
TSWp2qGE2D/072n5O5nzKQhRBHyH2G/KcFWAmlASr+MOAdsGLtgvZeefiP6l
zfu8yVYbU+9GbQZT/pA0cPTMaCrfR/e8PxaiM7CtOcjIg16jvDgWcR6r0Of1
EIcuXy96wxG2mZ9yzD/nyLlrxjjuSELf3hUDf1jRnGLFQI7tlrxHI++Q1KED
U+Rg5pxeYzbusAnzhwneRKXCSkbDPXPjNApNh9BXot9usqi6nxkAygQb/3Wk
G+gc3glVJEF740dBpgX+vyopGwcvgy5L/ZP1D6deRzuWZ9jgW/gik5Prpqyy
J1Dwes/Lh6bFAvUSNlWlDQ3JNeCwbHOCu/8xCJaxgE7dDYxQkKw+JFlSyFVN
vz1p3fULMcjz+hES8Kh2o88wZlcxlcsjLxXnhXdeCIuCl2cb8kRrTDxTpmM+
tz3QfU2bSTWtPYonXPJQyivMiAS6fcIhzM8P8UNic0gytAoaxEMpeHDRCGyY
b3m01NrLkNEQefjJu2FfmuCv4SY/s7F8oaVSTv5RpauSEXd4S4sSMqrVwQeZ
MuQ/j/FVO71nNJoohmxikqfUsqXZYbOt33j+RIV+ZHKL/UE/lLNQkrxYhXg3
GTMGO6ogK9xErqOAX+wMVmbCtXhZTzW6HFqW8+6hIN76Pvzg0EH+jin/8tO3
qFYD25FAZfkB2hNRA6qoMFBJJ1ggQvPYzWFxa+ZQh7twuPa73juNAZ9j9llb
TpeZgrAqL4/I3K3SM0o04+qIN3tdxRLZqyS06R/fNiTgk09AUtapSBD78T8U
Z87zIYgdTHaX8sFIZyYDjyFcIxyzME15cOWIcx7SdC/XtZl4y4a/OOszWtWm
FpEYrF+Va9ZtpX5ruR/UfLALg6gbDfY/3p1L3d8ovI7QUjxYK1UVNtymaam3
wvVexp3UO35PYLR+e6Gaw7Rhz3MJPsDo1zJ2yoIkgzoHBTD21668Zu7HMWGI
pG00yIhh/qHhq1EcSIoRElhWhihsdX6clPiohnOzGMj666rpgkXYutQvIHU+
Y08jH5hgTvoCHVlylXDg+Ey3ceOXG/9U+m1nV9ozed8oFtlPYpCFQuzEsdem
9Ygv3aUHwLQcRvFF2n9EIMKWir2h4Kj6/EAGY1I0bKdAWWJyH3sFuqpGwW2K
LKqFa+NJ0ArP0JOnDPCNRN+HXVFi28whchAvqfvxD8lbCRpBpkJtAPod7ztp
/48m6wWD2ZaGr1xk9DT7o4LxLrDpKLWD6pXTiw9NQ93dD6c9/WzSio1U0JOt
xLyKfLDjmJ5bwIAfCx4ktBzjizPtUSmnXzKORdyDoGx0ZeJd4m/mbHpzAa/v
910Aj3cl8AUu32IuTc+NLYbS9zEzOjg78oNNYg2l0oqN1PRDM8JcMW6P+uz8
RCud2jweQNzEh/TA+aVESM8CNTZ5yQHuIvPXoSfEIBkWpP84zcvYidyd/nec
V56iO30JtqgWZGpgYwWpwXfd/VJmSmS0iFMPVos1NV6ZC31cvXo9GB6ilQDd
zMeSthkt6dHsDLUtpCyKBzFdcLnkFYEQtt5PsTccaCytGFinUA3/qavpyZRo
e0W1UXWG68lHQAl9khSdh2Fq0OwFGUkCzVGTzcwzq2V1zjxgZH8HsSoxZStm
h49kvMfT/+2SDBIQ02PjlKx2ze+XL8Gfw7rCqZ9t2qYl866YFW3mvwkP+JHz
x77EwRlTWdIwIk76sOTFEFIhleohzF4+x9n5X92PD6B6rukC+ZRGJqMOWg0F
iqJBPGUwMWTWbXpcbxFfTP3lFF9B+4q6TKtgq94aKRV9dhemnGSDAVTVRkyl
QK2JEyaqXQANpTbLLczUQReeRb871es53sCPGVYhEn3bxHdOEsUagFEndUm6
Dmep22iMv3xyXsaNxYlzj02CfGAnwFDAbvxlxtZLVU+clABTVji2HkKE/BOO
KJxpCVZIgItseOwwUGRrj8DvbYKH7+PkoAhca4WrrKUL1HdnYFgrZPd9Bg4I
DVPNWYVAi732HsbH10f2wtVIQExE0pMBbO7nSFwcmG2WtUvEY9b1hgGVvV0Z
gWOF0s/sJglh64EJLwPCoIMgY2nVqkRgSKpsWUR0ZN026blOM3T8Sd2zYTqw
eHjPj8hURyhS9P0zYZRBJE0UxGf4Sfr0In7e/WOQhUDOUv7mwb/xUJVf1QeU
xGBKelIEHhak4qUz5mmUOqdpXKBsyYM/mc0XbDIU28s1MKVXMZdgwZeZKwry
c6Rp3cn/CAmdMplJco3RKuvOZQr1LD0JplYW1oT/w6RLwEG0+Qt0aMJCgltJ
5fAtaeElFsm3cz2PZm3RSF5pDycThuOFHwqpAT34/dU0htbApDGGmI8FM1o3
sIacL/hbq5L3+ssMISz/AtbOIfDngysX4Til/FuR+YnMWQ+pqV4VZ92Ee473
UWRIuKIULyTrFOugtvMgVeNXkiIzRdW3yLdc2ZbYYYpUuwrakvZdkUkSi9aW
poZYjWlFk1HNiIrS4ryH/1ecY6/S4esl2HmDuFxyMtYZJYF9BhM+dm2O8Iba
wDrYw9JAfD8Cli3KHLwSCYp8vBwwnGVUcgD6RqROKSiac+j0Rc6/SnxXD+Ax
h9QrNBmznAAx60Ymam7y62P1pzQy8de4HYEwtz1nlenIx/bh+hVxNt2s5D7R
59TM26M5CCvFs5k6u7DLfQOGEwzg3jlZVoDKdX9KZECggWG4Sno5vQOXGA/i
eVZVIiccB+JYPiUyneldVpqD+Wbqmus86gj6PchtCAzh3yTDsel6IpeUuxs/
SgOWRhhc7kBeLVZTrkvh/G4z6o8J0KgTez/XNUecwTagFf5S1dDr63TGRFOg
2HdX9/p26ias2JH5GJCDf0QcKwEvagP+6zqPGWfrORIYT3TatSD9cvwifjbV
ws92bC42TYgEVeK/WWiD6YiQfJMf3o+HzjWvgU46tANhXSf1yexc8tOlEvbf
KB9ZvEp6CmC+do5tkUDW+oeYFWmlj0/zswgY8Xvs7XjLUZfJcBlsRxksaMW2
f47FxdLIfjKKjE+/jz4G9VjowWE7FYRJwixJoLA+RucFh064ZmhbKVQ/6Xz0
QwS0ZQ22f5WQY64joc96pwNP6tprVXpxTshyw1jPCij6rCkY027qFUr5V1gq
D7M9kjlNRKYlHtGcPRKx9EmDuoBTFx0lhYuQPIxEJYVJPuYnpQ/b9KB/Micd
hbSu3VeWvD9pq7AggQhehGFAy/Y1v5d0DDgEiqliulekAvbmdRcUG3/70qL9
Z1/kVuPKzHnDP1NgxLcsomq2urZeUL3Qnt1yJvoPQKp1GTTQeZZPk+nd/rwi
VZQap4gUj3ACEyZjNMC4QGtiMnvTaavVmCdXqw70pD1c/RkJqjI/XQ3+8gK/
xlLMD2WpUPHrf5whAQe7P0cBaSTrQsKn3IeArSBjaNKEp0wpHb/MrRfN6ZO1
uK87lNbUoGOhwTClLdGDiu7QKf+sIQb4WJHUWNhj9SetE4jTlzqw0gTZ7XEP
Fh0qsZOqm9TWJPq6HEmoEzvWOXTcO40KZ9IBa2ksc0GPm4W5aawZZqlxnpL0
XgvkKvwxgDc7+5BHlvd/RjPu5JAc86Q5HGl7uQgSDxfvR/jGsdvMtk5+sL1K
RDEo498kph3Qu8WOt/2Kt1H7z4N8HwVXvMMoFba4o1+f3ZRVk8RWUWO3V0eS
8x3AOHK/tbbYGFMe2+yG+sz1Sl6t2GPb37ZXmu7pTT0Vtvz65IQDJfrq7U4N
Gzy/Xy4ID0DJp96sA9gYGkGMw38gPGOc5K/K3tIW31VTgT/C1YHySL+m1Gkm
uSrFtK05qe3Kg35wsdZU9rAloPgBj0fMzFiC4QwpLWvgx1kCQDsoklXHUJGk
t2B1icAjTr1Fju/MwZ4TG3ocTIVV67er5lCr9DO6yIByKQqnSfnekL2ZgROY
Qrrlq9sx2MvOiDdsAm9anKEjvoZ2Xb8NJ62nfxDVRli4qWCtgXL31EZc80qk
HDWjk2JvmnEz1jZb4Zd4QvtfUmgvSQ9zrp+jGHppUjmDvMSh2B7E5xSOa1vr
c11aTR2gm8UgIa3CkFAmHJce3uZ/h5JqBdZmo5aHC8MG+PkRjz4QckVZ9DvO
yR9jDhXVJTRr40tCa9lGffSUjY2X87lJZ6NkI6jaAzwz81RHoB0xJbAReU/Y
bb6yM/9Dwjb1QYDwQ0bUPBMQV7XH2TjWXb4RKP1F9eN9w+cua7BcQOAcztZ8
ufTCxjiGlXl4Elc+1dkxxFHbBrzHZM+qiTNdMaq6ywjOnU9TkPv1Iw1IP8vd
Qf8oXScE9Jj+OlYKr2gYgefXup9kqY4sJd6qJtE/xuYYrUExyipZcS3ii5Dg
uzCQnQUGChz+wH0lRUDytb7baPSQGc6JQMnPCk8kYrqLdXTq/YM8eiSmjHSO
op95TZafxPNXcZXVZsd5l4NLZJDrC6P+VohN8IE+76d8LeDMq9U4IYdgphdi
7JK343DKvt/Tl0hvc91LVYI2yTZoxRQ08a5zkzjQ71c4KhtaeawezjIUZU5w
PoiAfGiZK0fEXbJg4OzBJrcZC+0BL22r94WwdUedDI4QqajuGUWG3C8YmyBM
FWpvSu3ozFtC6RgTvVvh/Xp802TfqlGVRTC8hKEeTtf8Y5A2FcFxB5Rn7fO3
8ZKDeu52LfJoOOw7Bc8aQjboNGWiYjuWlpaa1WmJ+enecQY+CL6y5wdN4eiI
V1lbIdUHAMLOUHsbCKIyzm5o84hDqnw0tU9OD6iuDHNgU2O+IHXsuOCdQcQv
tskZRNlHHWxT5ZGFIDRnyYQWJpuhH7oHMtUH2w3W4tKwGIg9pZJ1rOdNjcu/
hbAZM4Z4J/Mo98gYc/IW0+8scjRK4uEube6curnK/ScR7n/XfSgQMYzqIB2W
QINhfiEhKUYXx/U3CSvVWGTD0TzyjUpUzRdIKIDzB1Q5xQli+8JPVycnOS8V
SeSTMibGKvUKbCXvy67IsmDcf5CSpywtfcuV34Rxo7y3AHVYMMk5Ck2on2/f
31E93mIqdMBSZ4FOEs7Z1pUyQ+Qw413FQtU+Rb+JtiFuta3XUGC4UJlp4o5U
39PpMwzhEeBmWghQzvOzQRAvLMyKcBGGde8XI0r24a2/xw/GPg5eO0+4HUij
hxN6DZXm4ZvmEKtseMUapx7eZYSMpnuEyNHS4gClo6I+BI/8ZWyzqsi6/DJg
Z35xxbdQor6zD2YmoG/dmsIQwP3bm1Ti/RLijYQukBQyP5Vn/+1vkLTvR4mS
BuJ6tPjfihgQ8xj96Xg94yp2G71S3mvlgtNAsLHjyg+F0vvIPaxDS51c9WaQ
TDOkCsbQ0ROlRtIm5elTrn2sxrsV+El/AcSdZDdfMQyIPr6MWBgPw/DLmlnu
+q6nAjj3POei8cWEWpYlhHj08gfV3CkclprXdH11ls2odMuPVLtApBbxNirq
q3YjDFlCaK+dxCoucBla6ba/m2xQe6/BUJ0tPXxpPp1q5n0D3ZOXOC1hDfDM
c2GAsfj45Hcn5goETfkBGk0OSCQE4qzLAxVhcGSP1KcqkipOLIhRO07o6kIn
nkeSaw952kUf5utcGHL2TKz0Um2tLtOcFQJISgu6H5haKtXeXJBqIDDHUB+3
vsDqsF1Jkj87cFBWUc8hFFN/TCVKuvIRSVqV3w+hRwoRo3yM/7LKpkJnMbuC
uk/qwHMwqE/OU6rV51zYp5iM0iftn+VIjRl4KvdDAWRu7v3NXqYP6vVuSFfk
cXED0Wd+Ba/PH06b4DROZMabZRlaxajtT/ARzogB2sQlft30GFxa3xydeGra
vw/DJr0lTCcYTEDBXnqSRH/RvuNyLgDbQ9xUAJoWLrIeIFPoUhK8cpCEAiLq
3U0bipc1q+OmZd5l93ErkaOVxAqtbNDsTA6j3hcfILXrBOpF4Og10RRJbul7
fONgZbNlsUVOaK18WnKxiG8ZyejTZE1HS50Bx1acZXpdpz8h4Au7U9MfSh++
nz4j0oGRJ3QErSwbRNQ2sO4EKr1bf2umf28TRiLdoq8+UAQfovKEcHXvN0Yi
HuqiXPIgOWIws/rMHwEiz4Kp3EgQN1CcHYasqzhGy8EmK5yiEkB38irKYdJ6
r1GcC9EKXG2VXkIxyOAp0CZvxY090wPXVEB933E0MGSAYuVidDV3Kcsu+SfR
8+YrzTX/rAD6FwCi+HrO6rAce8z/0LXn2/Pk1GXILUE1u9441I634YDpm3Ql
IPuB+tjFYc/0WWQoBK1YBRzxjYu10a482z/IfiGKP01t95QMU+O0C93VXMZv
cHsJQUBOZNhxVpsg10v/AWJPVfySyFmuK386Of2BC4on6d8LB/i+C16OPKhJ
GHrCQr3XcFsI8jFOqmavsIS8c8dBQpuwXb3Vuxhb3MG7Ri4mA0rX1w9gYHlK
PPr1h+n+sqUyK/Yw2RUS1GwC6eLtQOtuwu20HHS5ZtsvSyv72OfR0Wq+D5NH
jf82ja/cGYjx5oWUfbYv/NqbF63twTdx3ylaOyZslK9glnw7ReyMab1TyiNU
QbvmZ31vKuGXD2zzjCLhD6mS9wPHAVrVbOQ7TIXJFETau/pe/gM/Xl2V66Lo
XcjZSwcnlxDtj+I6yJ0H5f4eB0i/6beGkimNlZqyQG0eZTmnaK0zmmE330HE
40ZuiEPYNVP4hdGTy8LIio4Sijv7RGMz6FdMR/N8fIGDhX3v3YZsKIq0hBqb
ClbGpuoj/seVZscTtzy6uv/rE9vN7UBw5LXFSj/eib79jHwA8zZbmxNmEOSz
0RJgi3XdvlfnhkHOD10tonJk++WucvXF1d82vTnc9ZJmcDQD6W3HzXNT9YS3
it00tIpTPTknW3nq0roozkGRtZ4STKGrmz9fhJpWjMnBNKdLhtauKt5l6beK
EdvsxiKlVBHf/f3UrkGEeWNzsOy6043HU1gvATMLlJbhy0lrh4AjUh3gzAZL
MmzM4KQpaidA8ylJbGFP4qs6dDzlDQQhFZ7ztcO7KBTkQY0mALqSu9HziYD9
itFGN3OI4+Jrp8WExsqluO0o3/dcHNooSRG6MJEXmYPlPEEa/s35nTviXvxG
n5DMPmdpxNeQ2OtVFaf8HoNkiXKpxXwoc48SblI2kwyEbkFpeIWicdqEgCu9
pMDMasf01VVWp1H8JnL2osE8nBYxOB5goxLGEwAeMRL9Mmu03sHnzIm427ep
FFcnt5YRbE1I9n7GMatHiJK13A/36iyO6Je9ievmh1s7VB589L01+u+8o4Qf
P3lnb8GsQw6wx/YDM6ElqZgNqCmqT6uDa8jAGj8OpIQnPcfwyEdWC/+io293
0baXyviwmC6uNlSzFGZYjseN4ruqZe+Nktbxno8y0JiYu7XRnUoO80xRfubb
8arx2Bx1jDydekb+CyZSO+xkcu+JZQkaX6WxAvc81+DJz/X7+Gy3lixfXQ9u
czeuSU0N+ymRMaaR4cyRfYQoR2T8Fbv7MR04nUXgYWZtYP5rYESDIYv60Kzf
b01S3UgBroYtAr/MYWHaerVEPgBAoGiOI6J2SGSIYLIABKtVaId4UB7RPI6S
bdPeGdrP4JMcQSQZVjrPxRkJ1C0FXlNTWCu1OBXBLU5tf497jsxLy7fUR3Ne
yvwKHvzyLaobpGUcocvnyDjvLqCGOq0Gt1Qx5H0LVa2wA3c7TXALP+SszKt5
2qC1seT/iyflaj8khaA0LtHBDSSn/DHhcgjT4bMh5NC5B6uxoEI7XFh+EJyk
zutPLBUWkjcPWWjjTJrFMM7amuxBt0Ym34JoEiRJZ3TPIqrrCK6oOCPThmII
VJMXgDOZpw4MHFAy/mFgMCLwUvnwfE/GQGvFlFnzH6jTmA5omdwvkdNjttH1
t/yKt+TSzTsCf7PMlgdxpGzvRMS49t6MgG6Z7GY5sxRH5Pui9DClwO66Sdwj
2lQskFnmpZZxgk6hdqRJcGt7Y2vMCJE9xcOcn5nmTXZccUdpl1rggnFYQTSx
wuAzsxvbjkyA8wu0P468POehAVt/dzM/c8SHhdSBnb5dZq7bhpC0Chq8ZMc5
BoSV5wxVXYGmv3Ivphn4rCAfTitDCSkqmgRR0t+oCQSbf+DPsittOV6CT/wg
Q5O3nT4Sk7SgSMeADKGaSbudQ2ZDSxq/GHTlA5hTdvIxv7YBmWQ8H4QLDlt6
AwkZz7ePL26E5aGfDgaE7h8bYToE05Je9C+tSN+0UR9Q5UHyxl7kngv+SD7+
x2ROPFoXsLg0kDlVA23v0f7omCorjk/CvMQygV9jmrUOzi+ayU58kMgxCaqr
/aWvvIEbrMKpob3ZJWc4tTCBaEL2rIxMvDlPh8NtdEcI4Vc6PsLPucSc/W4f
H+RyHouDY/vaZtBvs0L0uvTh4pPd8aJXJw9crvy2fbwJs70suTOU8lKgsgA3
9B/gG7VlwmuVUhm1zjN5yo45aFQOLp+nPYrQPmCs31ZQClGYU/T6kXjwgCnq
qyzf38nI8hxf9B+PCWRJ0yhrK5PXOQ4iMG4DXLdeFRIcdlYDo3Kj+YstZ7ah
uKTte4Wdu5rR+wqOb1ntjnVkRO8fvNUAvFL/UGb8yXa64LfB/zDAxOifz25X
fC6L5tNnExmPA5K8O/c0/1nLUhMNX6ymnwwiASIcQhy1j1CVKxsGDp4gVuMx
l2qiDFPK/21m+2GvAnlvbE4EcV5S0PCRaeV8wiw+fYRQzMMshmLtzAlbTVtd
E8hhyb3V2OiDBFdsBdsmsPcUVhwHuJb5zT48h9I024phaCU9oh5cX2dDk6iv
u4gxi76Tw7Ak5+B+Lmq51uT/cJHkC9H6dg3UlEnKhC8jRQsRUc+bSag0Q4YK
QWma5+fsnySIAnkWUsV+vz40O/csZK/g59xMpBW4HW0eYxpigWw2OD7fy/wu
J/IuPPL9O/QOnquUc1u0cKaPYjFiGnxdrf+JsTtWJBRd215VCWG1hbxHObMU
OaYDt0+405VkjHxzMD4rl4hAP+psFtCZiB0fTepOTzpXUtpKsE1AzTsKfDEh
/NV7WTc0HQxGyMZR9xmOBXFVLFq7X0RRlkH1b5/ILeMcs2OEHs4aZSDh6Ehr
phxvWXDxtip62LZzi7kP4p6V6Xb6xIk3zqWB5BV9anKfcsRfgjWCKCQ9+LoQ
HMXN3C0O2zo7R1/+YXquVZumlF0Kt7x/RbOkHCzd1BgabLzK5ovctv/BvQ3c
jIZpW0D4Ti8/FgTcC/BOuGlJ8f2k2QM32Au38Q9XjIjsnl1DEC3fYoYo31kH
7/8QdHxGJgz9kzZh7hrFPwhk4a/9Z/DhOSumgtXyXkc9kNg8q1WAMfruiUGg
HDFIWzmNvlBE27A8X7CO1LNNAcE9Dvo+fd9bibAbIhTg1pQtEEIl2ypiYzss
dzGdeME9qq+uzdBnLTpBV5ZVN6RRq/ew0Cj/b2N6MqYA0DU6UFqk6f12fGH7
QvRz0UyZ00xyG0W46ZJV48xhdSZyX7j2pIGtJwHqM+XFL45CBmiymsjLaH7G
5NmVrA62M2A2gOsPp3Iy3acWvbFPFQh27q83k/pxIiJAZ8C1bx2RG0R2XXlH
MQOtozTcyVPS+d9wT/nX8tZtYdSgoiwpIFixIsZVd5AZsZ0I8/8LqfDlarZg
aCyrggKTtd+3v3bKB+LoQcC8zfLL3RMs9dLzO96zyluVcEhPN/UMEy14OdVa
mgS9Yjm+IVhiDrU8w04FEWwxu7/KonJ5IBMLYo0/9DQPDqkisBiwTRZsZNVE
HoZqTSPTk1wCuyZ0MUoZ2NsL0iPJd+aAUUYmjtyjwRMx4iB8quisZqQeR46W
+VhamwkefVQykGUwN83WeBiKq+FIOqpxYPpFuT9MURFQ7trdc70I31pnbnko
e/UOYZ3m3z4njHRtsNTjPy91wIVhQlX1wiofi4J2oBObwrYHFi+FhTz7AZHT
C+TNZMw4QueHLUm2A2F8gn/qKigTQugGlJYfDH9ITDQnK3qeQIxlaHi90Mwy
BfF3LacpcXsakMpI1lWB92NF7RJkOViAqNzlCiW3kpxVvRsLqoa5XZaLb4ob
VJCL1MJvsfNANlsqdhntWWSvKzxIenG+L/WKe6B0eawLPmuaHNnuN8Mqs8+h
csqAQZXK0QeA39Z+nljD9kL8yIIvvMUqSPDoHS6sov31fPbt+pHQcMnSx8aa
4X/7QR1IlytWNzyk+D6B3UXWM3JO1s+1TTfa14WKCMlUiWoVH7f3xvsTzBEP
owXj/6wL5lx8GLsZxJgnmVL2/I+MaMbCFkgppz+H0f94lUld20p040ZpqyJf
nfGFjRN6ratRdTuUZvAN+u7VSLcrs/QY4fU4G2IKLeyJVvCsHNfn2F8nBaB7
calSVKuPFMxOol+CcJmq1ZGwlaa5+oFIcQssTAvtg3m2D6kNIuq2kbxcqNeU
sHg+zjDhBWdx5eTWVaJGeKzqRJ/HV0hkO8wT/jrsx1mHYFPyq+4mR1K2sY9T
pdQH1iEHsTz9YFPVVENYxXt9VZL7nRmpA2JxJU+2TyWHvFidK2eTy3b8MSmT
iWHu/EWP8w5SUoZfNCbjEX0SkI0IFzS3ZcT9YCrOCxCuA5tcjdFc4qU9aWpN
YeDOwXxReMEQCiWYfFEHJ1z/bB+rTKG9HE4jxfZ5kDSI3zntU7ZeDHL8pay/
HVpiQshs3I8RA/cza1/K/i/x2GNJTwKFfr2C1hQacdKpM5qKvulpVSEKt4nB
zoTb3tv257Edyp7crM2vXkaYmQlyZrAKlCHfZKWkDXGIiSbLfFLmkWyRjjXr
V6Hxrt95kCKpLT2cuVEuXUAi6jSObC8MEuXMDpuxHjJNpwiv9LtehfauS1cM
pjK2tbfHYyUmdta6rJeBEjRYapPWd5cGp387yj+oPQod6TlHE5eq9n4jBeM1
PUD9z5DYg49bFtgHjpL63Gyrdd3hzP45SWhB7MHIobkQ2NrjAOGvkkg6PrCr
1H1tQOIwTrXPQPQXys44bzG35rtUiAZRsWHuFwWtm8x6ix+SyGdvRBjcIuoD
3eyuANyLQgPRsp47PJWMVdP2thIGZ6M6t10Pc3qpIkGk+UZhitHn72nE9IK5
fTbCb3yYJdP5rYjj7H5p12OsZCR2w3CrniIX4YepP6dm4bsXZcBfCsFQnLx/
KUT4cEnUoR8RDgJGi37X+AIXoi2CygjEH00+ayMI7LQR2v5DQDV27ACRnVsm
t6EDvA5issi7dxxaLOZC4sWZttw6kholVMoXSuftF7m8SFpzAeFoOFDiE5B0
fjK8P6KiQStWCA6tAWJHaEZseQItjrda5NG8ZSAFf27iJ3XvE4rs4FVd0VkT
Wmz3vZlpjvO4xqDQNVsWQyb3xDzOD/8n9V5QFS21rpaUyJb6vLjmvzbuALrF
V2VeJ4dRY9p3bjrQzL+aSH59e/hDM3KB5cY1I9lDgRbi6sKFz9v4Xr3eLzlX
IVH385lU/0mu/6LXOWbl5xj6h6gV0sq/K4+BYe1gRSCUMMFtmhdHQJiTXjdk
i8KBWLI0XHPWQx0+wlpRwjxb/+7zuj/6cVbHKMyyiCj8S2SwF8Btfs01PM9z
k8hKrLnDwjRT5Y3sIf3D8CU5BEZpRn3tYqIBKMk4CHx526CtVG1uelh/3j/2
9/lKLDLd8N0FLRwyRRD87NQPjtQezB3BeuK7NnlSyp4a2mlnf0GNZykNJnoC
EToQtXDM9aluBXIFSDo1yHG3spaU4aZ+zDvWWL4HEKbDmmroLgjNvPLWmwcB
4tbTvrjhnWurevU7LYxh6qR7k8vR5f08BWlSZEY7HJ6AJyq3WvlMCaWgQmFv
JLo/AmihXZs8n0VXYpLRCtkAZWqsWbCY/CK/ELNAjVW8T92JAv+zJsGEp8xw
z2pn68oO6iJFhyLLuudMTaZoWcgll83sIXgVrY7J8+PlcSyUk59Y4LTZGYyf
IrjBmVftvbshSTj87Sb/XRnwyQ5czsKe5LSCvl0TqUe7xXeeJVTX4iKYsXdx
f9q81awBZjX150xwrKO2jHswbD003ILc4ykw7K2mWVTWm2NDbqmCajNg8l1i
kwzF3JWMT4uAGN/uUiGDQ/XP8BXMuUi53P4bOCcGH4JJWhmvvaYenZPVGbKA
kxVHuBkxQXf3QRf0Bj/bbjFTgwzLfjyoLXSNjW5NuL9TjzpCnrrWF+oufJJW
LBV8FNoUp8lDvWorjM8sONwG6lKpD25nurw0eeDsvr9Es3GI/1OhWnlqb9AS
jGtAfwK1nnXvr7Ys/GGpRVVhGXDPgaVJH1lSdtWhdeuuJAKgMoqjYuoqjTNv
rZr5yYwuhu/zNyVGFppRn0N9iWDHWnCbywbNjJrlqtLr7SvlK5pk5pKcjpfa
cQWd3oPqx96JjMhWDNqp49t2Od2xctVU+o2ztpQDD2pjzTW1aj/ARHh7dQAG
/WInQHlgktDYZSHgr9b0gaXDuwnj85b6j9/qKp06jaExLp5lUX9u8EiPOhOB
1Ky/U3SW+R6ld6McDRtVlv/RmbyQRYGCszmAaDqgQxD4+kBBxLDnomgnON9X
V3iM54bhs9ZcyR2z61HtV8uB2NJidZxTQWHh+fusLGYDttCVtjGbwh5mPY/2
qcEK0W+mBtHyuwkL4o/wngT/9B2eKDhJfseVzquD0IRHlJ5l0FZ+vi/4ine5
1KreDjamGAzsHBAskIi2i03vC3ORRtfYJqO2js5pdGnifTyC9kO4NxuaqTfz
fjF2H/ZMzC1QBdlTZE1GXBleCwhmkqPZBNACrdazcVmBtbWWivO3ihyuP9jb
XFwicfTvtUD/LRKSrwFhMm4o8K+aJXi1ChWfGEfrLhVYyhvPaML1+mCqI2EY
REhFMTcNvex6S+LLE0a0bdXk8LQk5jk2UCf7WBkbCtVWm5I4cMZS8BDgOBYg
/rv/HnSJtnQ3k1kD55lJZ7lH2TCgt6Gv44BISzAdNzzRAqdwIHTDcbgKSb16
3D/uDviXzcyt3UbAq9EUgwPLPJK6I3ccNwHVxWiYPrBwZTj+vKOLyeBgCY8P
dAq2wNj9cN0jdCnj1mRqkYLMLWecQWL52mai4bHdmbGo4Rit6vsMVHM5/VOT
UsGCZKDCxNguj6fAutqEaqmGem//0sv5UAbr8GfQ1jr0Pb+wtyA30eF4/s4B
q8qDV3IG76bYxXmXn5Wh1Mvd2zvv98DJXsvHuVGmZQCGJC2Jvj7KLlYLoIHZ
54vFx/N85zBxW+j7uvt0yNukwiNauQS137XSmbiTPkSqpGG8me16w9hKumDd
AN+e8RgiospETaJ5zWUkhv2WZeyy03WU22APzJsB1iHr8a8z6x2dyhzXVdGL
YvIrk7HWq47bHsR90DVIa1HtNUbySevaJuwGQl4spvmvBynVj8BYQxjGpHJf
zroA/7lXfR0DR7K9l5BS2BPRw6ftxtqaPJy746p3O8bghXR71sgxtOeCIDdW
DtcplN5KEkt+XkGU9CK8B86+NnZXyx3kego95Kgqw+UzKqQQp9Ys2mL1e+I9
MUOYmi13OS878bhay1ZhL5II4rWTzMjAUBbXwbKRLzkL8XtrhrwGxuOoqPNg
o3a//LZHaQHuLSmoji+w4cuxH5wBi++n75XIgeZSmuv8KYOKafFoelnRdURe
BUJZrFNIpIGGqFBQUyVCnOv+ETiFus4eECSMgEwSBhaTt1YaNwfe8yQLOmRn
90UjxYS9A9kk0JjHXWQf7hT8T/PSa1Z2WLQhgE6GNwQ6D+2COsRzrujVHh2G
+IrdZ0cFbg3Vm7KpGLGOAexbhfO5HhOU4+NX4bVcjnRA2be42cRvnk5iibCZ
MZU9aUTfB4v9e6MEpNFEigQir8PJddVAqfj4K2cetQxPkH+e0UOPUgIPdaxg
Qlxzi+KNJskIFu9O7XR3KnBNTxzNxHJcYSQIupgjp1GEBAhvRDHw9qRP/b3g
SlDw8Tl6pVrhYfZb08zAKMC7bCvucIPYtzx9Ma992L4FrJ0mjqOFHi+AVrY/
E/E1unJCErcU9ghML4X8+8C6SSy/dn3cM/hXYmsU/Xm3UeZBaRz9bJ/SXt9Y
DpAG/uzUNwKuZQHLRDJHtcXBq6VhurDwpja+mMbNFJYXoSGFy0i13k5bYwEM
g6XPUTOxfBMLkBkYBdmIw72G7MyCaR0Dlai/mHh/67KW3Eq/Ql9hu8Gq3/tu
NAte5/H8K/RWzH6zqST293CGuOCxcHh3mUDIEmAf59qQLKzunf9RVALMKJJS
ADRkIlG0t2dMfF9h9g64OtATDgeTh+4yMwxhWVqM3z6In6lwU1ddf/UqP8nW
T8qatLdGUcXCqcN3QTiUfftmRKpAq5cAqHvVxK+hfUKJyaRIkVeu+F1tC2cL
sYv3rBemJF7uQn6bO8OOhcjWcsBu79lrjmFnJvZlO7A06vhDcIH7/nb009nE
4zCOwybIitmqrxyhz2zGEnpwJe81JDqnSOBdrJdGnWShmUzZ6NdtD1t//aRE
r+XJ7DNy1CWHlQT8s2mNv36WccD//oGKgQh+GNdBINRJfGEReEbwRh9QJryb
aasSYNrYxNvoQe2capfq5y4Fr1IwYDCiG6SRq5vcRFsLt5sIyQNsZ49F60ta
25Oeddo/rpE//DccMXIg9SwS+KpanIQH9DLZTIFoILMTpXLCvoKwtZSodYfZ
oX64dZLeVjUMVMcVs0s2EPqCn4AfLA9Z8sSMMjNcImF92v0FQu6Rp1+ZJRtR
h5AYvyLeUjcUtsHs1K8JZYJkxvJnkgtDyorZlrEh8c6SyWM+YIMmdEQDd/zK
ObMpUKuU7XNIgYTFB94p7tYKlvbmGZGmz3s6KRloRKsKTkWN0hWxw6zjFAEk
lH0F6VXAa9bomZ+Mk35CSLuuTOYnzROKQglUkHo1b0ypR6DGJmFSJSbFwRxP
d6Bp6P+agNfP0PGgi1DUyfi6jwBYIvurRozU6AdIGatmIHGrI+S0O0HLENMH
U0S4R+hiNShX2tY9/ZpVY8CkHlVecSnxpxAj6kYWpZgDVLqyJFkwefcADmmI
WcUu9f1enH5a9Hhp9aU6/h+JdSB8uF2beuXKTLo11jmFPkKc5Uc6kmYlhZBj
wEl6R6JfSP9q6CUDg5DHYHUGunZeULwd77hVnK46wH77SiKWWah/0f7NLV5M
z9GdHaabYWQesVLUqcJhcGVyivUml8bw6SUgnftk1Ak7Jx0ciivcZldhlgXU
X56UYDHkY6qee6fKuP8z+xCb2Wk5fyWzz8elePofzySCUMs1cstJ7HSwLrE2
rFmDsg3Amuf0C1XE1oqBRQOWKcnbJw0qm553hcofsEKaNamb0+Jg77K1YWxp
m+x3ZwpHh8+NTlcSUKtqN+qRTkaqsumrheLxhXiaRz198Tho7RdS4d2KKArS
/tGlFBfyLa+lXur0RKi3i35rh20TjnTQVa9bIvpfArbHPzprFHRTVYLuSHIt
lHtI2DQpOLcLRaanNtltalzYROZtGsDmXZijm/Zbny/YsbT5O4xVh0bHiNNk
dFL0ZQ0sJGZvYZPXptrg1Lywqyz7tY60FVvUSo/WhDCPg5XvaZDrDOvy/mxH
7JWRVcTx1dwf3663cAhDo1JXhQWSLEDnZka3fbhyf42Lyvvo8jc70nQG32+Z
nSr71w9F/0tBfaUYMJSU2e42m4iAtZUN4kWq8DCgy01kmei+WBWcTdcpArK4
83p0NnerBLUKgqh8gZaTp4FEZJsdfhBN/klXBNI2Wgt0bBOuqA6SrlIfnI61
+DphJFvibSAMS7m18bxjVzwfNI6XyTriNBIN1w5lDLdFJQE8W2pKZBDuSrTD
Wx85ezsXj0M6/VNiabYpHTQQi3+FRbUleJzHB/7o6QkhsQFrg9Qv5HnuBpVW
LhmaFOwHp9g5uWK1M5TGTQTa/mY65jzv6xsoleqvPYUI/EqpqnKerXU2Yfmu
7xzNuKMYEzlKZ0lXjm1dZwClctXUe841+NbYGt8Te2TyHU+tmphjJYX3jwYk
bxw5NMa7x4HYlQJkaPLbAk45QRDyQt9UP9nuWxIQRN9/Y0ZE3n7p7GJqwNZn
26Dfw8jBw8TGYybAz7IphPZNlqZ9OHM6HTMgD6WzCtGuej0QueX03XZUOq9u
55O7vegLirT3vi38omxDd+f74xLXFx4oDwH5fVNq76YzB6jGZkDSwJzNcVUb
1fRVTaSF7ADXhszT123mT5gb3xNkrawJiJp9xd3TFnoxMSYAKp/H5mgTORUw
+j5Kd9JpASmotDTt1tma7QrR/E31NevQs69tQ1hTDTKESUUJVQ3bnKwcSAai
f4Gl1a0AZc4MlhDXLGxJ9qw/y/7iMVCOuFa2DrCHtTwPemP33j3QbJtaSZDS
QCVjeVipuAzbCIpMLkOYEco3VBrdXV4/lSPfCgy+9fEVfkcRZR+pEgrQpa9W
k7i57DMkyJnvBmVGgHvz4LDo+a3s98rVoyPneVcdtUFB0jJekrCWrho3+7ys
Z5pNFgEbf5Ub0Qql7sDdr35RGUugWXg1Tntqly0KbVrpY6fOuTtTEdCpxxIh
GN8WfhTu2bnpc6U3aTUoBdMW7TLwBf9m0BdGIJWQpaKxN67Aj+rK/XOi8t6C
EShFmb6KZJrrRlhDXExGK3BywBHkug8AXoTNfQ6K4WUOyl1Zg0V086w017Ee
HGetioEyz5/tAL0L/jMKLpP8uMyZbNSSKJbX9UCEy07jqVX+NOEycQ/FlQkH
BH86Vqd4p+kazrnPLFVQQOP3SR8b4cjEig4u1ZpMj/a0oL1HzPzu56imfIeD
5KtDrlDsV251LRQngkX1OwOMAJLhaK1spmFp4RmzvCy9UKY7B4hiuzTZLTxC
mgBM/BBaA4FPKXyCMjNO5hji+eBpSNbpEMAfCWxLzIkWLwI0A3VTQzNEqj6k
Ybaz9+N/wBC1tS9rCf4XFeqDmOSi3rL8XSY9GZYXfo65zUwSDWyqGKWQ+BJI
R08WMjQzaggQa8KWYq0I/0akFNtZ7HMEzTb7RWUBW42e/bdnt+Ex1KEqPedN
J4kkqw207PWdMpnuegfDlVjRzOXi5an4ygr+MyIWCOsfuKgOz1VnSGUvNDXw
6Ikd50yJ+UrVUuAQL9SqMO/Qk6wEnb3ka6Tt7xrqzL68BrUKU8Ts6saXf8Xe
XBFKFOPNsZVKRRw4oCIS5Ja53IgZWiM+XJGjsohUn2Jv6IibO7eHvT7i32Hj
odVDgVFviyeXK0EMiGp1uag+n2+hj+v4wOyksjemkqLenrYPdjJjpnfA+DjW
4lGb5EFItu18aCfrw1vucI3ZY9cPtVpZd+ZrZQ2is/OYkZRM8ao39qWGfaM2
TnklIA3cLfOPKZShGQfI1EUM5CgD5CrNlLOcJLf2MiFF5f172KSotspCWs4l
D4cNtgZL2Y+qwtqJ4lJPeA7B8wiUVQvXg7qvax89ohMCfIX4dQJddVF2QoC7
3GYrMnL6YBLle5RIgdF8Fxwfe84qs2nha+bkKBg+DHK1VJtDR8kiDFCEHCi0
hqZCzpfKPK+0grGaiya11BEg2Nw4r36Q9MjHZNwc1ubLuaT2yJJAH6Kdfo1/
XFzfRPVTiKQqBTXyuz4Kv8NdtCkC7ACNjD4P4OHYt2aNuQXNpLKe7f3ha4LT
xcNQrc14+8KbGXXsb5KEkOdCyod+oC2W/ULiYiNzPWLDpmStglu9eZKOsE9K
XFLtilKmJMbiVowFzss1mZI87jYa81jmuwT/KMgKahwuF53SbrV831vk+sck
NZr0SdBYaOzVwThE7XGE37uz182lZOh/BZJobUi1UPEFpMbS4cAfWZ/iO5Lx
28Cu9cugEwNoFgeSuW6I3Zm03yA4Emu9t7el9Vb0ndqBxZPje1UVtaGpqRZY
guAmpFFefoVTTFOjAn6L8jE73j1o0hgiULNforPBAOmLVgUWFZ6UZ7RtPDJv
ccLUBnQSS/laX9Mo/oAozswzRGwnGQGQaaolBRN1X1PvPIYO/3qimexdW0rb
a5aQI46VtJyH3sNMWoKBXTJIIhyGDK3BPd5naTsYV/azG+Vdwu53tjBmWDjv
40FC/WCmrGZafzfYweUoKXLEHhSaiilRf7RwDXLuqX9bLUSQZKsxPS8pTowy
K85HwvW02Lc15IMetXqCjNzq2gB/beXBuyq1+dsj93ECyDASiWnvO0XzBGba
Z3rV4os+gwklNOXmAwnr+dCeSWRUHetdnaxMbOXYoJs8h20UiNw98woFvH55
uwDFU7Z/5niPCvo+vtBxLNdmBgaRIIPbTuVPGwhaxp/qNKTd9yVnNhkgTzqi
EeV18TnYoDOJlqTCxmerUONEK8sfMkcBTG7kI2H70PGrrJX4sGueMkhfbYps
ToA9LY7GITU/FreJSaANTEkikSsB8kC853YMT9RKAOPBvxaKMn6a6nAmn+vE
+vZV5011wqb54su21tk5XTFDV7eX9Drp1+uYLq1IDmUXQ3seeiQ4/FgSAfKk
AQJP124kfQSICPgwwVakSZdLcLGm+OG3Ck9hZeKjtNL7P9IEEG6/1SPllVe9
uCS3269YQo3GSa+4kMIr0PxeAwAwm06WeZvqQRbMMDmFUS668zisqgvBUH7i
zrSOEbE0a0afZL03mzVQnZQg3iHnbPPFPt6L9+ibI3P7ph+/bPTc1v/k/3pl
tq88ZV3h8rZrqnhABAvX27DZyKAv7KxYshojWxAkC7MJl9FjI5Ufv1tqmDbN
Yk3dLfVJqDsYbjPMi5vmURras4m5jHmnrsda1czvovCnepd1BRy5prw42wES
WXwrWJ3eSxAVpaYqzDYW4/P0W3DU5sRQ+UfFnO6VlW+Hdqgsq9qVWGpH+mZR
SgcxxyYvONq0CF/MIwXNaXQj0iMo+asCLh5It78GLYTDvLePODOUUR47IPYP
liwXvB45qifpxvNDbiFjTUqQilUBvePVeYXFEZe1pzmAsQGAdkMmpTiClMLs
jscjgF5qbOqgvnL1Z8Pkp8FC2RH9ijFLwoIIO/RxIrgcd6rCKsRjNJYMhP/v
cAbk6dN33IWLYURTj4c0kW64X+mlth2OEgkWbQb4V0jCZAR27ju+b3CvbOiy
YR9mmRjdCyQF65l/BL9S2GY0oYlypmmV/cqhn5BRIiC+lsxzIyfF5NG7Lm0q
QNoN+2vXrgjZQLcSihGsOZSuL2qvEe3QEAwTd8jBqVgKbGq17N4PG+f0vX/m
pHtFYZE5dv1fwA+/KOuhJkSnKPoqnaKFLsOFlyMJRoL/E64qIC7JTt7ED7aX
p7gjEkXiVUFzjQCusCa3tM+de03FFWKQlglCYpdFjVH+v/R5LSmfKEw2VnY5
QsPTMOZSjVovZWydnPFqsfBS/040A5ptP/wvMySPc6rPq+qgsRvBlo04R9wB
AjDyCFZ2UURzMR3y1Vq8XHsYzuKMKPuNjirmKug5Eaenkb1BlErc5V24MYj2
J1pW6lRxdk/S9IYo+mfmbGGXV8kzrIejUoHHQA8xgbjmlA8jU/lhfieBQFT5
ha0LcsSDJ7NLJIWpqTIc8amNGetU8MhPdmvEJ+5oiD9U7tFS0K4XvmPtWpjK
NcIPVjrLlDmQb/MDj5AxlgDD+wtF2U3hA0KBVA4j+TCGuA+e16urBIDtHhiS
i4jcPdf24EiRnFOfpC4C+apoQUaZFxxWiYAz+xDbgRojNoik/Zo/khCXBjkr
hhUP/8JM40AneMSpqe6OI+8XcGAECh/10/z/6AyQbiR4g/+2kM3Jjt28vUHY
U0k4JKZ0ocx56y6sckT9gc0b/N+TCUYAkxxV93+i5r7SW4MY3HBn4LEu579C
OiNNNOpoy+FHAVpUEgmQY0vnpc/n9BiEE7XEqnxLzm6U+Os/Mq4GGDYS5Pnl
X26FbUCmGIGMUYxPUARyWvAoB3EZzLdK1BC4rHGpCpvy28MtMcbAt6HzdGvv
MHQTorZqzmbZV9iN4/LDZvfjEu+WU39Vu0/WLjhXtiEp4f9n+LXdTzd00DVY
v5boH95M17sPtKCjgoyMI9pEyU+HPw7TyAxvkjagvmLmZkBYmjvzDw4g8gn5
zuePS1z8Uv9lLAFznIO4fnLS1yOeayvwr/3JrMgtFFDruEWf/Zkqh756CII4
cI4xESbgtSnfSDFZwjZjJQymkNGva6/rgHC/Kno6XJtodzti/yAkAmEjY1qY
MTyDKvRuDzrMHSvB9o7LSZv3AnJvGiGedIaYrMRkwsXrhgA+VRuWb9XhhbhH
sQWoVgPPB5mkxIDcOWX0Lcw0kzBJhk37MY1hmLwEgc+oFpTjfmgZmh7bTt1r
r9L2AI6HgVZibQhVGS/OclOrkQhEfOBVKE46ySvHLm+i/g6mY+yqTQewJwHG
XFC30myMNWPZBkp+xop78/s+XWXtsmBt80CXT8zkuse3p5r37dJY8KTvMMAe
4Nef1vY5XiT98YJB8s9W5QwoPlVHHmbOhWuekajBNZoKmyGAt613HI8YgC7s
22zElE1NIbbyu7gbGinwMscRVpxFyK+uZKtJbaliaMgyeRdLAUlpkU6+sSIx
1dyIom0ErFz5uRuDW2bQK2ZrfBf/mSp4sYX2zwKnZ9YjVLciORLJ5ZohS1wO
NF1z1DFM2Wn7I2LNphEEVM3HaEX/0pu7aLLmqg7h0EAdeejF2ADn9jneK/Et
BHuV3ySwu111dF3JFSOgq+iPIC23zY3BmJ13ofIY31qHS859zOTAlzjcsF8R
pHRnv4iGbv4Z3sKpI8evxc5+CDdKwYmqUljpEoIaEzwLNzz++XChBDqMTkR1
QdTtM2hUTWTI59/ZpzrOhEYVyQURLmgrPEqrBp3F3R+oNZTiVuI45Esxy/rw
svl+GPXUTmlvrIleYDkPaR+SWJLj6TE5H/Y6So0NJso8VCKCcyaJJqdri0X+
+FLQy4oTLMhhmseuSYOABusL00cqKW/Bbe2Ml24jg27ENVBQTQqtu6ZurEPF
DJhnpYfUtRg41GZitIesPYrj1/9gb1fP+Ycq+C5nvtkkicRXDHFohqscikfA
H57QLPJNzlwWFWTplpaaPkeBMU4aDfNVZ1IIsPwwPEwI2ascRhwmRRAl/dge
YrdfmOkmnZNXRK0FNoMI+Ez92djxDuq5R/5IDGuLeGonOfPfTBk58XfTzaVl
omSwOJewScWT6mXvMsaZViOKHeVSbI4o0QF6RmrPjyxr7Tb8oafVJgpMuDq1
WUy5ZJEgsYpDfltekOw3YVDhUxievRYZ4LnLP/C8E6uLkYfxfw9xoumW5v24
dn72Nqt+QlF4sx8PshDJ3OqhUQdhpZDtKO4mF07RN4k7+Okk2/jF2BDb5DrH
g6BgcGHSxMeHzZXeznEK583KIMHHk1J8eeXRr8eGd3tUVNN1qL2nJx3A7j17
bq90FKe6opadNmNq13omcS1HUPqnhf2wHb5+6kFgiP7qq79UgsB8WV8aQzT+
9FjtghjCW+ZxQx9YOBIXM62CgdOqNvdrmOq/9GzrjbcK8EQlrYkZY/XpLjla
FEOXyJYEta3R2AkD+xE07TxAw62G7EdCLnK3D24/G4ff8+knTsPMDTqlpY80
s4KSd5sDQpPl9TQtJWaVM+/rWUyYTHEfBSAGrq/zCLPa7yDQ0jzN/XibVFsq
8mQH02j8+Rrcu8jMSCJHOyA1ypslZsuEL5mIpVnYWYpeFBu7/JT/9ea9aGos
QZtSrEWMS8WmlthsCJY5UccZ1OaEtO1xha0nLFCHx0hNr7xL+8Adka9+eIqk
pQb5N+hMjBMlyhIaxfnZpS3BufQ44VoFjYIos4RvSgyBLFVFIuSWRfHECP0d
1cf3+xGYRMefVAncKgQR4vNvv0/X58CpkDFGx22WHcKS1OBc2W1ZVAb2U6yL
sqXFHmrNdAsbWkUyZ/udHwAZu7aafEvBVn78SEcz4QckW20IsuckpIoPbxmV
mqd8CxOt4jnFDNpGhxeXACgOQ8LgnafZwQHK7bI42kb6LcaZFYFPs8ZeMwnJ
K4115AWmYdIdgwpWeyNlTXOFambz1ubrJn6ZNM6VVhXq/GurC6ebDzgq5ELs
h/XBLMxnGCmz2LVufs9EbZqHdQCOVf1y6yx2ghF4IbzFFQ2goVsH1Mw4Z3o/
5TSU/J+9IacTGg6dEM768RSs4nW/+OC5DuC1kfMuVl1BglWaql1ZJwP3gU4n
7h36hT21CCzAhCBku0r99MTBRG3uGDKzqU4nOlPsihizZs5aUP812hDHee4B
p1FVaukKspblPfCqaw+32LxMkgfngs6WlQVeyL8bL6QSDTz4WK0YMF57dRAC
Bxk4ZzbXlHCwTAREbTsx4jxZPW3hBM3sYBLDbxQXwiJZNgBCRS9B4ZoHw7C1
HuKB+cXsOBc/guEjcWjja6qnd6HYj1curKpN5CUb9nxYK3xFFFlVhZoi7gqy
nXcKTWDivBURKPNs2gUTQ4KNN0Nr6T6dY0ZfUDKuqHnNN8SjTpDrJpl3tFv7
sQxht4X+8D2sRGC29Duyp5TQ2xxmFGqpo57+ymK/yf5MNN7h9W2HvXEvJ/g9
zo/mHbHcW4tPtdKKibno++q8CTRYnoSzpHbzPwtDf5AhJhXNHLSSj+Rh2Crz
VD7wHKWoP4tkB6dkJzRcdFE7r0TODPl1iPg5ECrpxtSVlPLko+iVI/hLwWEK
11WSoHTX2R6pjnAOu78jaLESm6pXVpNnDKExMufh0GY6CPxCF4ZdaXLLqwla
qmtH3AWrDo8xGBEkBi9j8YQkNdBOVAWpWs8gU+Zz0b31qX9dVfojm+rfwZN+
Kl0nOnPxXEgXgPnrj00Fle5549slg9TvYeAmQU0NiFhQMFoJieJOc1lp8Pp0
DxpnmxyK+diQVUQ2cQjFYGHpAltV7pXK2XSobzEN+5ZoEmRDOuWlRK8ZnJZJ
qg0JV4/aE4+MHR0aVhxgqXf+6+Ok1hLDL065qYvTpjGUULx/6Zm8m/5iAfcP
jJfajfyYXjt8VbnZBS6FCp7rYVWpyNetQKaDV/WeGnn00zwwaQd96T7rqS+Z
t+ZnQOdmu4XmtQxyobf8gx7iQ4THnJ0AcHkxQ/k++JfMVyJsT+zAy7xcYzUp
ZGOrL4OdxJrQPVYBfYXBgCb9etdAM+RNztrMa4DjikNEd1fTQgh9Zdtb4TpA
TR6gsfSgpPwm0DTiWoM1da4Vb1e8Wcpx9ntv4wefmJ7lBI1p2sGXZ353oyja
NljAo5Dm4UmLnfezmz64D9ZmXh7nP5CoJaV4VS76mPUg/HmJZjMQXQU20KXW
++cS8fF5tqzM7iqbnvHkqkwONqGC65irS6HSHHvzPJJ7UlzeMnsaP/YiQs6i
WF0aFKHGmgfL6jwarcDkPy9+63J91cuVl082MachbFwud4ronrxcv2vMwA7k
Limzo5cuftkFiK3sfgi0ZCb/drc1C32D+AGBOaD2EJ7vfAiw0TP8lwWrjkE2
E96D42S4DB+dt+4S8xwNEs2tWLmav+iB6PcSUwy6jqCoTYO31ILu5VBq0YJq
kU1vY8yxLNCDCn6Erq6EDlDXar6lHDJF2+OacyBf0swdPworPxBVhO/EInWd
j9H2o5ZmaQsKMg0s1KHC2GZ52HxjFYvMvqFdxo2+jiblHwcDocm0Xt/J3tsd
OuOyP2HCqT8bqXYLyW/rPGFD7nK1S8C1fHAYXLPdsVNmgb+LSaDPIY8FTW+o
nLiuqUJG8HPJ+6YGilmcu1i7XhDYaQJn0DHL69f4LA+IFCFTm85Zxe/QWi9M
4PH6ug8m3D2nT4eFL04TnN8WZGtGwawWQxUp+uCRgUaSrV1insSNpTEdeFlY
XDUdy36l6OZ5VOmIqlquKzHZcne/PGa8JvWGd1w8tm6IiZiQxYRk5GZ1T6ZP
rmQdK+KTC4TKzAgqm/QJd5Z0u+sme6NZq/4yIRd/XrYSNOviwDKVeKGA4Y2f
SLMTNhYsQjTJHIMPquhtWtKz+zMXw10HQM+u8SQdAbe5jJLNOgTR81pj7pvY
skBeNdr7DTVTHzPKj7Ec8v6SzKLF/JOKIX+3ZMks1bvwyQF/JmhnBTe7jRM9
zVTaRpElRks7t1Cv+EWw2DrlZHBy0EXnmOGNRwKxFi5El9HOFkdAnYzRVVHi
oZxsx4Oe2/3eYWEg0cIaGrKIlvTBZwtRexxv6upJvn5BKhqAtNU77fCD5Nn7
GT2Tqyea6HZ/WmNnpXoAaR2m2WNrQ0gxafMPlk+6O+lURZuHuMNPdR9V0f7d
XhreSJi+ITYPXfQalQHNyqNJuQL6ObSOo1bWTOi1OKdKtnkMaMEAZunq0ZBZ
6xXrOk3poeKbkZHYbIDigqNnbA288ntMSe9ccfJ086dmPqewSR4d/t5ClXUn
6UkGimC2LSlX7cg+5u9puWTwvocEc0wMQsv+YjWYqyN8DVPr6bjmP854cNgG
F671xm3KZHuzGV8gl7Xb18ZH9nBOvQGh4Vh08S2g6WwdXjUcm/l8b6udS5QR
kTezV7f5VCql2ZWQ1fJU5ylXLb6f8YCth+nETUIC+GpXhAZeTW2LLLNWI4ft
ewd2yLMDxq6Ci2CyDzYTqRRiVB98GdY9LmeLg9U2wtu2CTBX/loW5EYD5sel
yK5JjERdLDpQsuLoyHcdXVdrZk8WX36sLRmXqywi/Fa1kKwhwl2gYSkAa3b7
pcWNPynEjcj9QaOjS3wyeacWfPOTtW4aEUVdHUGKTqJQK54GlgWtI0f2W9/B
GsqjukoHkpA4R+Fe2PLYYimr/nLhAkWUh30PRbMlUM1OG53B68N/2n+19paV
kSkXZMX6FTDRsSnn9NPOylhO1uUnpX8RMPCkIqbt0KEv/OSAEviRtKSNgqVm
c3Tu4zG51txrRB4tA+QU7iwDAKNfQQRe11QcmMfZ+dctlpkvBrWcshjvSNJE
zME2giAWdNa0X4mq9pe4K9mrD/oiQe590BEqL3Ja6RsfQ9UNVJjQ0/egAJyV
pwpEUJ70oGZJBkkzETbDhZIF3DIdjAbHBANRHqAwrNuvoC/nVPsZpoWSHdiq
KJ8gcD6awcYfV5fn9G6/JJU8eE67+8aIWU7jIIcWL+0M9RUCpSZZSsOsDKl4
/fZxPy5sMwqpQM9EvJFXqVrvefWe7qqUH3cw4a5b1jYcKGc2c1uyhNrNR3Yf
9Dt5zb8FxDCAzCagvoCEgfC9AZka5Y72R6plWDR6MmsjoKX81sSYrnNBPPf9
M5EfYSSEV5HkxWMLrzqRqpFcbeUeFfkpN4STvFuQ5NbHyzXAwsLp5BZe5VGW
iY0Pwe2XI2aT1MU9UylhVK3vsg92xPVrxtn4yAj7kQpuYeTgOVdhNdlgU2OT
t8+VL+rRJgR9QW6f5GzNFLJ7BEMtZ12tblxYBgDbC9mXlqeXQKvr3wE9sNYE
n31efgqPeKyf8IFCrTBEvf/iAsw5qJjzvWW1VEGg4w+kqZ1a6UM74ydGYq5h
LBUDTVpJxVrcdYuxjW8WKtgZJuc6ryReAXr1sbFi65wyg6aPT2v9iMJhgGtB
UFkPLn8C8VDNkE9Ts9lzHRXZbqhHJAiG9LKvzKt8pXBacOoqyC0rtLa5FVBc
vF0K7AB0kc+5B/kMPexxWwgFT6hwJAGSQy7hCnCu+jLTY7dkfv3/hTGhEx5L
V3aw+GkRZ7LvtZIWsfH16kDiEDRv36Nvc+CcgKouzSfxqRaNMhZWAcYyV85B
jEJsOvrcOiDoX12dBuxZ8G4xuC0gIzCXPgrf1qQXmlYaTcb0N+HYtupdCZ/B
/CL0TWyc6JO8/2pvwDcOzZxm1i+DGR9JOLeQudCAHFgl3kpQWd5ulVFKqd1P
Ll1L1K7ikCvQtHTBK3b+UnRjSILcPwmoCOfyQCiGunE0avteC/kA5yBV0oGM
PLwvq3yrui5yuQNjCr/kgb5CbBEohv4mIQ6wMLREMj/I5PKCEtxMp2YlqSAk
ZZLpVyx6MWIkErnyOfAh+grNPpKpsuU6VcWFCWvzpLtVEWqkRExzN2PPsnYu
6Hs8pongRViESj+AgRhF9xm0IBxOCQ0Mz19TRkWxiseOnvakBZw3q6jioJjK
7Sth3tlreUxNVYcYc9+nGBdnP+I/AZ4pcoc3u5KqLRPTjmEw8+cuQcNippfp
otACUOxnJ9ignZGicQuXzRSfP2RotguTzoVMbt8jrvqNtRZERuEZTK5+CHTb
IE55HU4RTpl9dHrQNmk2uxnCTsboNCWrEK4+Xkl0b6xd7NxbH2wOxilAbW6G
q9jDh/EMMVDru6QcC899/O6vmTYKA7aToqC2z77LGCAr5qMRSADrJw0OBLRQ
vdc79/PqkX6zVecAvooFyjN85FEOVotTWystWh6r9KNOAH5VW0CvoRRM5qPc
TawGonEJ7YBpyc6vLxEAaLIwM3axS2+HgL0gcuSEP61dmvqZPcU6Ek97iZ7C
8SxcqALN70BbOGY1xhm8b11vFYMqeTvCAai8r3ds/PIYLGqrHXaiqy5zH86c
exXNgfYVYA5Sa1ssmLTosDTQmyNF4kfDMbQhYZOP10lhKKKQWjYVGahUVYq/
AGzIX6HnNwioS/+jWiKNZ7S2pcb8uH2Xzw5S6DX1Ic7CgLcibcfjeQ0m1UbZ
pN9I5NUuK4libwStpnt38mh1y5xN4Rc3C46m+ZNmqOhaJBs7TOOXydnro8tb
BcjFuMoLMxY9p/YfaYvLG4WU5SwB001kpqT/i6RL1AwMxb3vB0Wvwwz4qB7X
oONiClcq60yG4dqo0rzSLV5HzsgPXv9+NBHEFGkr1FAdJQigdjka09YkZXAh
+8uGyHLfNDgIJybv0fKaPjgY7MHLedFclIYn0056a1Tpts0x19kYJt3iizK/
OSLIk540z7lYRM29ARprUiv4ayUih0Z4T6cSxDs3McvnMYqeCZfyXcpg0Iwv
0CAu3iyKL/LVUlWIcLqR/DVy2jWV9y1Ul2PoxR53GVlz8W3zjThijh87n2Jj
eXU1xlusThhPXrYPsIHYiR0NigMYSTwoI0Ac0Tox0P/360Tr+OKRM8tFUTLE
kSKrAsGMkDqqG4zsTnfeRTyRaopWPn+Dmn4HMfI4nemsN1u3VEntRH/csqUT
JNuabNhzri+myDcT323xzLmKpHbvFgC7zndSge9tZq99ipzqe8dZAlGr2hvG
7AsfbbHqb6iKftzCFusOp5Kkl2eRKC8YBgTL5MA7y0px9D94WHn7GclfBEXZ
TbDq5XNUaNyCluSDHvi/SARZbnei62MfNYXPykF8vGNFb/lDMQEnjDtAK1g5
Kf5RNy/rVRJaG3Dmz1RrojpDmUb22S8R+bWd92OUz2AcQKs/HPPxeQ8abTle
OB2laol2hnm0b2QrpKHkl+nza1vofKIJRNxmCZ/bRZ5RP0o8nOjWUVz7TMS0
1RWkSTAB5eVAXRaTjsIv/qEBZuQWx3NwFKyqCWnMTzzBE+9yHUgMY2dWOda5
j9SvstOVayUPTj6ObNXG6MO9/GF4WXqhgPGWprhXB7snyWLaZCb30NhXIKtC
Ln9X9ihztBbXTjtzgtrNeM44KEC7WfZdWklVQcYv1c2HTZOOoBkODFIfOZqM
YzKyLHvvsFC/1XCvM3/igkYsoikXTDSY9jDgacIS4tVqSjiA07E8P9lBLRh5
3kxCLxcpabL4Q4nv+pnD2DwHvPi8tqSUIk2PuNWKiky8LgFVaEqhu+2jsBDa
2DdRvuUK4oG6j1zxe9gRJGKjNSUpK31VnOEPQPU73OHJt0e/oIiLZMvrJcUV
9XpRVPr4kDi+MzHCxr9nNxfF0fgClSNiOuqWHBMHQztrMKYrc54hJiZYiuQg
31bOBVq1N4i+AXkuQnjeEztrv82umUAAX/irpsQNQbybwi5MS9AG6+wSll4k
JMKYP3vZMq/Zq1beV+nOhcPC1z49AovMJ0x9cbXNbdd0AHlqKZdVYxn+9ESq
F+H2IFhdkj11XqUH3hKtyplJwgTNjagjuPaLfKtk6Fj3e5c+0JoSxGf3tqA1
gUc8HT2Pgkp2ONjyi405pIyqJKbe3oWXqnQLDddtQPrHOx7D2X6EAeMcHBAe
KyuHEkR0tga33cFQsYZ9184CcLB2OgsN5d/yxyiscnhvYPXdCJV4W3V3zt5t
yx3yauRpIQ7+SnV8qnql6ATPnireO6xcyybZykxLnZwHkhSfbAR98Htxy/BF
4oJkM36vT2A2MN3q3OdrF6gGaq1EuMKDaLPMje1bigNm/7NrqtlGcgOhtW3L
1LEJxP1+LIgBBgLilI966NY06FKAQD5gIhcO+POoSSeFEUZ8wR1TFWJvC9AD
dnwW5eYTzfbjtHrKJuUhXM9AcHYLd4d/tOiBppxsqzBHQ5aSfGQ3zpHezIV1
S5fiPSjc46rSiQxerVqlsP/97j23G8mRjXrc/C0jvTQ4cJXjUkS39FVwN20j
9HOZJzBojo1JIIorsgszFOjyt06VEF9yBeg9MY2zRDr8go3rP8T47H/7x9eo
tZ9+24ffDBCPIDSHfWSCiSMBDbsLrdVGbjoeMF2w8oS8bspZVQFUtSUuqknc
oipMz0SJ4aNjT54hYVyntu+eHw+Zvx1ptdCWXTpM4Fhnroe4P/VXiLk6CxX/
OUJ+6GvH81JbV7ugkI3yFW3F+cHvDY6NW7iw0jFKIyBFz1cvdytcD25laQfJ
F7NaEbbvHimxi/WjWRj/3wtkYPB2qEG7vrjBS1C5HxcIJ/3xbR9VGy8qYuhp
Afglz8bX+9WGySlj5/zyAm7cwKipB6TZMzSa333KCNWHaFG3oStHsF8S+MiZ
sKzcKaqv0/5FfCyHHCykTwl/Migt6edjF87sTRc6pwFtskI5ODdNZ5ZW5Wq8
cywbmpV512/h2PFCu1DGd2m0s+AUi59MUOXFTRtW1qP4P9xJ/4AL8RGWzCOO
yHEu5gchC2SamedH+A8lTgpC2sEXuBE55nasl2urdoUgZWPlkAsA4Zs8RnCW
3C/glG13qf/MEzBAVF3ekaGmwn/kyOvSqaaLWpSQmeiWlRce20EydNfIymC0
TYBjdhU1iJz6DihIv84SpOPvZsKknkSg5RX7HYcdaIyKmG96cvlxp53IMEnM
OYb/YhZkCQb8FQNOapFx05rx5B6+KInnAIBmB03r4qgw/4YFIcS/epCIojw2
+r+ljHpX03MU64y49r2+OyknRiK35+fPRxfhki/wA8E188veJhFG9xNJdnLQ
VCIkKdn9Kzo8yjI0d4PpDtsfcvLZRs7qeNSKHd283GMcm3jiVcXUjiV/Uk+p
9wwchM7EasOgAOs8Tpm9UT4Ix26fSbuj1ziKWG0U0oBtTNwSyQfBmJMZGq9d
XUhOkSdtT8lUXWV+ojWxtp5oYqk0kDzFI6j7GYp/IFs0USnpwwYQljF1s1vV
W177+mw3Be/hLHWyjC5nQCF1lGwT81/Ae4TeCfpWzHKGRZ03YApYiYrt2K+z
exuDNDwArY14i7jIGvwbLfWwduaCGdTepbEPgmaG3rpnva3pXSbOv/byYLbu
DGeizyApjd9PPxQvQ9Ap3QxP3FY71CKbZfGymWu+SaXnqpCX9RLLO1y5hKnZ
aMWOCx9xMD7Gb3Kk/6PNTu7b0mYiXAxhgPE2LHgwaOxbpKPppee/MbnCMX0E
LYMVVjguTk6kZMY8YPg2sBZvBu46XBGIkVjG13tCdBejacIpjLcfT2j9etsj
x5m606mE7RrN5+LbfGoU6NTkedmb8ZCc0sJCAanUx+DfnIH6V0jekPjNkI8x
3hzHdN6uxDnzqGVdeQdFtDBzlE+m9t4GpJ+Sh90p36SniQ1MChDmhqAJyi+Y
Atbl4Y7NHsUXy6jh4Mwn/0QPl6us12gSNPJTj033A9PYQb/0dZu7IAHl3owR
t5BTvVfbZTVLbuJu3P47Zeub/pTyiGJhf/9TxCB4BR+klq4noXmhdApUt808
IJhzIdcESmFGUgJ4MPmhG/hjIPcDOO7QIW81tIWzldo5iJ3AOpWi2JcsXtOn
SCbOJqlLNFKENAsGDaqebzYChhtEm+VpNMSX+XE1DYDW1VtaseMtzWjEGrGL
1jU9GBcBN3WHTGWyhBOLyq3YH5Erjr+dKuor5D3j+qUXm1DEBX89JedV8Fwx
n6eT6dznTXkmyN9r57UFW9gEgtHn3yMixH1+RAoJOB7HpsEkBjC+jpL+GRXb
PZkXLmagX9ikTkVmRrjJLJ0TbKsNV0l5FWrKITbiIC7xe2DxiUe8JTjy4i6D
s5c5M3Upt4DzT9q24CpSdo0UOnT/eIxNFujqZlcYy/lLJTCeobL7+3sPPYb6
cjsOLGiuONSQMDNCay5NYBaHXHcBzpxuRHdN4x3sNS3fvFlA3dMfj8UfcSdH
eFqEMXT/Jx3ZF3ekIyVPUEivnUX0TwsDqW5jW3SLScEnJmevaDCXo0w5N9fq
9nXIdE8qFc70r5URfhuMrXIFhwFs5mf7TbxbfIvX+EJvFwJkkx1GhIQdgO15
iUlYz7GFsru7MpKrkoRs26RZ/cuXxHjP/W1uyUf4EX8Xtt62C1WDq9I08Q/6
BRy7mBVlJEToYA2UAN3diWJCYK56cTAYnY837/q1iVED1R2wL+wGUGsU5KTs
2TuooQEweTg4oPngGpbttqF/bNfhzAQY8tqQ2xlxgHkR1Wl8jLi5dwVbtFLY
NO1WEnWacDS5BgRm4PKNF8RC2Mm2IYA53V2YrP6ncLe6Z/XTx2+zwIBiJj49
8xllH4yD43Et1QlPvkcZz52YfQHpl6MIavnsjhd92CT1F75SDLdTLpPIW80P
znOMJw7QJm0wyrfOxcuzn/P6Bu1jS79KLuLyonFJsoetH4pKUPkU3NJCYUdr
gH0Uf/OjualHqbu7Q1gKM3WXRVpuZc0iroZa6AR3HiZu4kyGl7kQ0JusX5YY
AyakJMClzfELwvVYxz+baHGIIfHT7qzeqFeg24cN0EDk0keS6yjGgWkM8tnK
V8YdEUu2FLTPC1E1NwGFy+AYK+T7qsh0Br+baKze8e6T5FfZhTzf7uI5bl8Y
/nxPJDpzRCQw0sd34q9IdXoXS2qFPkCfXbz1LfYPwgIUGCkJxB9Ru4SsG7g0
K3qpbPHF0c/oRKV8BCF64lcy+AmPwO+S8lY0byspwhEM+fDFkECpwSj2KD7T
5FLu09Xax7fSTx2RFgBSjxZOkMYAM+Uv7X+q0Q0+l3KomhLjMfzftmWYXNpy
p4I0wQBC4r6gVhVwwMZdCLOUtnsvvvZE7TKf7Z0/TUQdU1xxnAQkSH5TUoDX
WwqkaBCvMKUVytIPoAKT9lBJpwnHrtHtgZA3PxszFv4yKimVZE5U1BHUhx7N
xnxosqL5xwyAu8QOH62Kw9pPM2rPn0feD2AUqxXLzIieIKh7Z6CFsttu8LM2
5u2ypYd0LMkWFAolTA6MsIVv6EW6oGvVjkWZTVyul7nELu5M0y8MvfNvvptW
juIBt4rOvE9DYyfoHzlxFQ6L/1QeEyjx/QUYQJp2hZc+4AVB/jwLiVDBoBIf
uODDtOtRufHzn0ZHIxfKi68+mf+zamq6WVTZwH8K0rxG/592587WPkQJvGIu
yBCiPCrzjXd5gq0sMzKB9r0FpoYL7fMhZM7E189f9Go7AG3fOXC4YVt60Fsp
fnc7t+dG8vGEEG74LZApQRbrIAv4JqgVq8yCZTVpvPgfQrKfCRy75DuYynhP
LE8IsXYO9svvHg0pJ43lGJovsh51ljZmlq+XkjFkUFnw4oN0oTfYUi5xtF6c
IuRJj3NS/Dh3Iy6JICSTxXmSCdt3wsDQH5BuaZWFm3P9i+BqyOXVJfr68J3a
7ghoDu8Nmj5oy2VNHeSCoZI6yhUBTEzBd3a8DREYvZd9oVzCbN065fdj6HZf
rWYwd87U4m7ktmguo3tTtgJnGBClo+oRG1+f45OGbio6lYlOZXgO/i4hO7nh
tP2bFMKCpafHBopqmRs1otNXIRGe3s3stbEmjW9fo10C6WSIYYH2hDnEcOmA
v1Py22yCmSrTUUfG43KtbCRFamJuYMrsnEkUPy5lnl41xL4YYUXgSg5FirGi
wH3JSPe6HNB8SNu0EoRYJzgvTq8FHjfR1p3TFVbDpZqgs2MoUAvD5rGMM5au
43GR4RO5hfFpxkrd4dz754iq+1gXjwM0LUizA/n2f5yDKNl+jAHDpjZ1xZOq
M6SEbRR7drDRldQ6Nlg+umBcAtVnzN2txKrqsGVNX1PLk/u3IdJv8aNtIH5P
ypCO86c/0ppQQWuiUVF0Xd041AdCTK5LcrASNlN3w5yUlQV/v05MGbDblf5V
fR+ec2gJ5XY7sUHXylsQNVIOM17clIOpKKZqYoTnw75Yhjkeo0mV3QUZYJpu
fDqd41NoRQ8LYc2ytRFRijju0vBkB6NZjfHgRk5voTwgSE0Vq2vvdx3UMFwv
Bi2QxQunFlfjbk3oO+jMOnDqdCBYIDfFQNRSeli6cyut4Z0wGX0tRdFRk1/o
+r4PJWo3cZGhRDhvVt4GCdogyN/WB03ChGbksLM/OCXuUxMFzw2uEhYQJYKa
mpjTknt9q9jJdtnM41WIL47Welj1X17o1dOMyN5Gaw5yvM1siRr3E+7S695u
qNUyDwZY1imJvIt6dN4aVlpHQsaWmKp/Ok+n79aO1ODjKGejv11wIrhhW3zU
ByLuYUv3IC5A31J/PN2LyHJMMmdooEAsMIWAoh7PeKfLFxZmAzkZa7ezmlxZ
iJm5VryBnOIvRyDs1qx3/VPXwGvo27QjYABCLow2yTyvvt5QhkJBjXRy/SjA
8EHTvjWMaadvjGzSRqpa8W87QXtn7J3wF6BQqeQcAUUfxRw/NrH+AtdbKqu/
hyPgwpZ6aFEzyFRQhBoP6NRPlAdJHRaCGY/avFvF+hsaI3HGMjhuUanjYUbV
qWrSYvftDV/1TUteVdbMJwCrhn8Tvcl4gijfYkH16bJmYWNycCXJRSLftiOu
hqPbBEawJstHAgsvqQgz+nIlA+a5EtXlJG6X4xYjYIhjXo0l0/UZQ1PLEDBn
XhclBpPRVg+0boo8LGoaH1/7CTvC4kKlQ1QNk0Vhd44bTf2wiX5T2p8vSL7g
AuK1UbFxBY5gdE+FdIeqgPb9h53RpEB3QGK8UqX+9R+n3/KPomc+m+Vv9Ucl
EMt0DH4gWrR8nwNh8Ijv5XhsnTsEm2R2qIBnRtkmWAtlXYQsyRAH0I2Oz8dS
zge0M7cMwQtrN6bWEtBIACO3I9RXNm8FcCQwEWmbli5knUm1lEgwwNnymGAi
0snwr+nL57iXfZ7PrAzlH8iFBpbdABfAFuPSy1bLv6PAf5RN3MPvNLCvfnv6
qBxQ0SI3XxKoBYZIWmWvFDB7gajN1RfP8E1peoZnQh+tbK61c4zflf4hd2Iq
uXOXpCfHX1o+moUdn/eZp8KTRfWNTMME+B6yXWntRiC+mTSsebe9EbcJt7TF
WF5FbxcHoIQaG5hQ2KQQqzwRJDHUasgJqyHUXq64pCtZ6MVTnDGqF9B6h4hP
y1YTyCAjPM2d3MZ7szz3IV1LdOYOOhvRrzMoBLWpM0JjwHTXSLF4BiKQDuFh
tnwZnR2RjTWiV9M2XLjPOIb3G5XXdsup7VxjxYkWSh4a3nxnNDnFmiNsCnhA
Kfjxmeuqb9KHw8QKnIHYa6vorwCC83BX9p3i7Lf3/X3warFTISDMOWh5bjZ9
rSKZMq/6ARRL8sgLSodzgkjXGY7vlx11B2akIPIxe7SeSWO3DArbgG+jg+Hi
qYYzl3mfCQd2ugzO1SfZfDMQCSYwfOeLoemQ+lp7GC7G1xYLyhmpAeheO7vJ
lbZc7J7BMJMkwu5jibt7zeGMKm12kqVBtoVy6YfYiRUbae8NzXZgp/cZcZNv
R59yImsJ+Ex36R3sNknmlYkma1KS9XwhFdBvyzVhmrJ7mIoNKc+Hnd0iEIAI
9DRSZVJwZl+QDmTjhPSZ2FsyEF0ismxPWpW+T4oHoJAB3iUshHHhBtUDcn7H
U+1DbnNvnLm7BuraXKuPBmecUyuUdipJcnVyBeWTMpiybl8vCO0sulUO8Rh0
TQKdZQXLHxUIPaOp28pv+mxR8f45AafswveiPjViOfB4zwDt97zZK+n00u1B
SCVZxb7zl1kClpCGB7jPd+tuRlgBZz8FMCN6GWXjH/3UOZGutE752G/Ih+cm
S2oLX7WZWBGJlOh/p1/h52blSN3wC6YuRncYG0nzPUvMfAxsxSR9dMtXYy4Y
AlyNmC8LnAf4mraRThJ0pQ1mGTcBU9ZgYIDGmk7IbDtJIkb8W8T/m7YAKGc1
xqKIGkUjrlGPdtv2Y1AUy3Ipui2Jy6XJxmyjOyiEFZK9MKe03tp7AesR2gEd
+BkGMQBTkAkxU/FK45Tv7pIgGeDptm+sMkW//lu1adixKkmT8/Hm3zYIs04F
kMcf8YUF6/EN9tMxac1uY5g1j/sc82qr44C3j47oJkK8ShqhNFemlMUJC5if
88RbrcxJycngMvQ5ESIz4jN2buc8I0vHxhrMkFDbtm0dyDYj3wy8OTvv6Fi6
zN26z31WAj/fiZfxM2rWdMfrjWWUTdPtbClJzqyF5TGeAZMvkwnbs6HZ3bPh
LUoaJcWRHtRt7YvqDSjMKgYtMtlMw3jEomCXPRxX/mIr+NcQMCV/yy5MY9D+
sQXoD19+n187FuVhmBtG6GPsKJh0PScCJJhZVl1i0JCDr0zEHSb7p68uHwhs
8TbB5lZF0Md9zrjkw2y+DT38ph+ov5fgOXbUEAdPk8V3olY9fcP5pZK+EI3N
FPe9nKSBpCeYmnFJq+4ZCg41UAWhNDxldzO4LDS0txdfSXcFbEjWXmClnaJf
T8L9HOsuTwWkPIoXfl1zMJ42hAbBzj2eRaVno0LZwPIW9OVg6e8jA6PJyPj5
nxs44N4D3GLR3RJo25tT92cE83LdjNuPNS5fduB8KfOZX58g/jb524ni1c0k
wQJhm/iAtZJwYC48QrrNWDFvlUnRurB3DeXM+I6LVqrtnN+ehtxRkXCGK2ZX
CAqluXxVyOYGyl8zntuO84w3tXT5mbY+ooxX2a+PzCp1ajs+Y7qgUlpvSMdF
ryYTYvE54380T2UhGTwOQyUDcSCmF49u8gS44MJl3VT5SZpWbRtxZJpyBPJ7
9C1WaAYKt+bPw1feJGZnGJPedPLJTTRrUWRzvaVl5f0bVws7VS9vahW164cD
0geM4YPxxDApbrazA1jsDZSDTJcDDdkZ7Dv52pqD6c7Hui967Y9phdAqygQm
HuAUWV2WD4kZbqPp4OgKaSt0+9eaabwvUfOiPWu9a0bzMhF4+DOtUU+X/5VV
kv2CfWdVetsxcjvBSIqtEFj5Gj8/qysIIeMRfpX9qhxhr2M4EBR4k+DwU0k/
cpfLWWWN/Vt6v+yFaMCq30UrlVTgI6VxK+OoKgh3DrmsD5KHaTHtm/qJtJ6U
5N9q95oN3FNlwZ+4uNIL++4QKnTXETx7t7NYHeaf3kOq/EPhEW1AtY6ExVJR
6cPp/Kj37A877VCg971tgXylzr5FO0kLZJ9uuPAhQc2J7eyLHsO7XYrSx3er
2fGgqqGDj6trdtIlLVUgyCR8uqVIQfHOgvKNl77Wd8zXa8w2ppals0hp1tdq
96uaTfM+ihbjonBNyitdD+O8wJEImoZ5BfWa2ji78ADToHLo9bbrPCh6MN/p
tCd6Wm83hV0fmzKKArIkjsdItl0mZ7JRlQedynykF1WtFbdJPu2MIh7xsSXk
mqU6rDmhx8SrVh50HH7GcQ1Vy5EEKTgGsaU/C4Fd+0NjdC9j7VuxLg00x4KM
jDVdUHQGFir0l28OLzntsjSim76SacYIo00Wf28140uzv9XHFYOnQbWXoV1C
FPJ+IK0rtFEf6uIB1fFwDtcG90iCasvfri/MnnlIIoik0rPdx+aLzZzR+WLP
YAzvjSMqrGgsX8vJIRfhDnjpz178CqkMFfqPGxMzJ2JRxeB85imaf+vSZs+q
F/zIhyccYtqOrVhDKTqXtRq4yiFPqq4yGXayVPfcwsNo7fUUFmas2wqmCOfz
cPD9dbK8gH4onwAov62bHuMn+tNeOwho318iYLZTg2CdhF9FYqygqbk6lXet
+m2h1/vsWE3A3Oh0N4A4V+A7RPs0emAv8OG5zzedDykZUA2zPH4IDzfZqgJd
6kDx2YoEeawatkOMeKRsaA16G05MHv7pY2duX4/bXO0qnuDY3ikSbPoGAq2v
6b4BNXzycHjvDKJcQJQLucXVZeSTB5CmU+faf+eDgU6jHFyCh3HscA6TMTV8
85Q1o+ZBnv0ga9u6DPYMWl/FfeO0bJqEIYq7GdsKslahacSCZisPKpbGov6z
VuCTm8BWBsoy6lBfhS1BC5q7DY6kshvePnaX6LL8q401imFyXdmzgXt3gYYI
/T5sarJDM2CeyCyxfCNJ4JKs9gPFHeLN8kMADaHrbrPQgd9q8JQA6RNGOILR
j9tXH29ldmLekZ82aPAofoQ0O5D/nfEkgYvHYkqOwOjBPWSDtiEjOmZNyxIa
uKAOmVBCgopjYVXFzLgg8CyzKkhYS141ABuHvDHnxD7Q2dLFhW/v2+PE0uy9
56nUdSBnZ80dPnA/qiC5TJeuMl/acPP6Z9QUFDwmwdUQTIQkR1vPQqr223+c
Vciuqm2HzQ/OZs/0GWsDbaUGb/UYD5dKm8OIO4sEZerK+aCdoeSUs3CQ8TKM
UPFNnZTdJ/IUi+clw8YSlbyPc2h79zMwgbeDDAP7kzxvsjsD1s23eTN8epfv
RiiuOwEKiG2G2c+ZDfQ2QJfoGyVET7FxqizgCm/y1f3/X+r1a9eeacQXHEf7
xotl+uexFsTg3rZ3XJjGtfdB/QlXWe/KQMP1oenEXALZwvBZUxi6AbNLdVhO
ZPzZr+FBp5plWmFXEEuJ4Ja8wbFzF7qY9zhVi6GAhLoaiEZWEIiMUYqKxBVl
0jmDoxO+aFTZ3M8P/NrlnhUgqRlMKDjMBae5g97c1xpbItfTsoEUeIau1t9d
gdJXrYtl/DNFPo3MNv7o3dP7agQsL5NUwPzkjSsngPdlZ1OxJVuXj1x9a0Bi
0e0Qf9icBE999SwxlD2xlyIvNvWfdbs0CuhtTFhpuogrrBwjgB9uLrQKg4Vl
92LbDcjhEY7F0G6GJhbQTUamRyWV5XuGIPQ+ZTV2PGveDXHtZx2Zlrpb6arZ
RX0XKDbKuIGRQxokN1K+uHN8JF+vfHVt4mDFQErevnL3Rx/V1RIK8iZrHOHr
03+hogcDr2SKWZ5JOCU7kp0WfHjwF/fzkGpudbrbEr2pt5AQy8PRtcC8m0LI
CnuY3ydiLiMfTvZAy1jSoKjGCvKg1qq3xUVVEHX9Ryr+XMVfQx0WTn6VlMl/
zdiFsrJ1ib82BC3lZit01I3msiJN1zxzuYgUrGiNnLSOCZG19g2VAwscrN6O
L3VOd3bXOlLamcNlmREWHMo6oYaCpCA7tDnCoJT3xVRF0iIRxbIu87871xRf
qJzRHwhAsBak9B9ezsT/oliN5rBPgCJ9tWBAe/iPimwMOaEKnzCmjRaqVQk0
7xMAk/egIOPFcw+tAswGzwzuQSkuOBGdqFQNae2bowe2aoatSStLJwXL+N6S
B8gp82s2bo+bJQZACqIXlY8AsSa+dLEZyFAx2QqxICYJ+K1Eq1w+7lQsjEfr
7J658wV7W4SvV6mKVh+0JoYMP8uUS72lwjOZsKLOVTiEI73Jf0sohM6R9LAM
+oXMccGko4ErrXRgdR21wJgRK0ql9CIa+lgalP7BdGO0G1VAKLiOY/5X9W5j
LZqff3RcP/HDZXhAhQqgLnwvWmIiGvgZX8vG4oTjYASjbaLFG+p3ouy3yK5c
E2npuxVR+XSG1fgCQfX1kLQMMjQh/imijCY4wx05cMHcYb3qaSxas+NoMQS4
NKFkNxBA5IC/c58NW8E53mYY2XRvKxVhapCqHYhrEte/TiZVDL52RmVxnqG8
LGEs/NiHT+DeZK5VLDqBev5L8BvmrB5WDSyJwPKDAtvxZzKEPpgXYV6l/Qmk
6/Y7M/NxIvFujtAMGYj4G0FTLyMtzOqt/NYm9n5T80fsY/tmQZYDMLLzuj17
Rhc/yVLLrWn4bTg/xn4Z82Cl5/UR5xl6DEuww6klQ3P+DCA7qHNUsuM9z+84
f93oCPZtuJP+5qHa6QbKI0Whhd4fQ0mk4oaAW7wOzQGOMcho13GXJKR7hzzp
OPeS5m/fGrXc1gtXl3rai4qx+vkEAsy95gHMYAmz3Awi5erSoGkFUrM65F1o
0i2boEBgj8Q2OeV1R+b7DKzL/WLu5rmwSdeK/uaNLpI9eXpVpgjB7n22sWOw
XUoOBwcQjn7DFLEq5n8b91cbyzKsRZ2eAI6ZFmLX9/5o/0ZqBZsSn2DkvEGN
ZXqQePP+M+qRLIxHx1kpbVuiVX+e7AeJiMZQOwcCHFgPrNVwZL71BDi3mkZe
bU8A8wa7ogI2upd1qilKri47uYOdbx2tqZ+THE7AyrFvhOQpqiHCEeR8GWYR
5X0dku3Os8b+zcJydVay0b9wDZP1A3d8CD2Tg7gwpg+0FP1DRDSf8f77N1Nw
RqQ1C+uzfu7tN/uc1EnGbgAqXoVCMoGkeEIsmxj2G7suR3Zbqo6nh4EWdf8C
y6yP7rIMWWJCx6kR7+0rkYwCoA5G5a7xyqeXjQG2AUTgtgoS5QjBqpsF2mm/
2KCVlVrKK8oc1ED6wB5h4gGVcWO84gZ4b4kaypJniZrg+fM7ocmSD8kG/tTQ
ymYZ602AjoobTV8j3Gt7v5TSW+67KqO4Z2G6xBEC2XN1y18H5LazY0xtcN5c
lIVvXDFxjneh4jyVyXcFaMfT3Fr4vxXqnErLaCKUqkYFq0l9QjUXAV1TaUJt
raqIBS9u3l6iw0CDOjNovPLDG5Fahjx+ptZ1Z15hTF84P0lL/w2QtFsmPfLT
/JTOdPKY+8DW3EM8g+tNu1GNc8DmC7qOu4fulw5wvxiXLyDF3dj9vGvhFSXB
kujc98KdnXsECYdGHGcVuoeHv4JYwZQyWP+lDCDn2ONWYO+EBsFy2yKREyTT
f59n2ZM/sVggonIoHeg7aPD4/NiBzNlHdfzDCKhVPHGQ5WSv229GtcSmQt6y
myCY5YCfZB0ZPF807zNB/0TFG7ye+o7QH7jPtWXIwjpqEL9eZxctCSoPcWqb
rUCPWRySofmucHZBLkAGWcatq493yYXdaxa6PsuE8uNtg+dzewHPkxRZ1CwE
GkkrM5Pp2I8+M4cA2Eubd73fe3HYiMTNL2TuTSozwYfC6sHoYKKeF7tPvSnw
oQ4PcmVY12AieurI4gMsOpcXfDI/dLnrf//g93hiiksNSh8WImCICludiSun
kqLb/EdrsZzItXiyJOR4EP8qawRv9+mdZeO9hVoW/BilNt75bidxSuuAU4ms
lZOosqUaTCYwp9CkZETOPuk27KgKw79mNWm2Im4np5ONpOotptnrPMXqy3nF
BVAdMz6nU8F1rx/ajIOX+yp1yD5hQPQ/1bIuXpRpEXWMcZddg37OYgWFhVph
iQ04npuNHaf5YHexDHC3CmW1QTgKAmhPLb0JlA76UUeWQHNbZ5hABiTxIYXp
VKsqiL+gIu+ESrm6pEDHcuY98Lr9SiWwVo5IneZEdbSblSVjOkgBoPpoNJcX
ecHIQ5cl33C6b3d2D/JWAeWbx6gaiYkL0Tj5OBsmrQ5HFXZG93/8boimSZC7
tm/incJ3Kbf2ykxy/9eg4BFB544MQujbXYh901MTugFOP518qY2XAAmAT361
k68XE8N3YrAB4SJX8aMy7cffvo18Fwa6i7rodKWcL7jcjhdZQFtVeHNFPy0A
krh8O63CT3IGsU4SIIznhzTsLqqYRRFkP8cwXmKTeZoupEG5BUXENV2jmIJL
b3dVD6gBbiaLETrrsSo4BGIMNahj1MrXapQxO7SFUjTsyNJcoTKaPfM8fTOS
ZXR9TC3c204Za5SdLAQePk57C25cHysW+XknUSbo0FWGI7vOZvH4s6yZfU9+
jpZDAewZ1DSKW9MdLvkhKJg/0aORG3GyiqIPpy5p06S5irMU3gQQzhcKytaM
CZw3PeFai4U+uix7jg4r+/Q24qzTR6IXefn/tVkf6femwlHU0QcVomGVThew
+6zDtP9c5rxU8Li8Q5gh4VxKHf6mLW0cLC51q9bNFKW9g+vOrfAR3s2Sbovy
nOdiNiCy9+wycLQwzTYIHwK2xsK56Er8X3AiE5yy322sAt5Jyl1cQG5RWBnq
7K0AfTtQ+oR84XLJxOMPfEJ62+/wJgJYzxVR4JiyLvEU1m1EqNNX7coS2qtH
A3iYauaRYpObu2oyhY2mgxGYROWHA+MKfM+cNkx0TOGcNFpQhV1+VFMaBEeO
w56ACjCmjqCBuxkUqVzwPUnsoJcbKGbElu4T0dLFnNRWaq/FOiMNpX+ukokD
duUNRhaxmINAOuOA+vqtisJfBxsJN4nW7K6kBFyn1ueYjnu2LMPCHlPLrwea
ahYxQF3roBg+YJXfR7aLWjEmfrcbn9tNVKUJWcaRNsubKybJfhy5lUze5L5K
SMsxPHlwysfiNzB25lP9ycyrgroOOr/rq/agqBi+3tYvf5lwUGI8itKCLl3W
XD5Rx8OTm+SnfxfmMDNSNlrqLIdfJyjw6bau6cXL8v1Wa0sJgZE4AsMCoaBv
kOS3OAnfxpJ+beVztE4vXeXaJt54jbQaxth24YFLO+yWlN48yDRS3pw3uvVi
atR2v5/Qer+REMfht2i6FqzLxBWyWfQx2A92cimW/nrSEs0emBo/RfI9vbIu
cHrWOcXLODVkZ+F4dez7sIKJm35cxh/wqDV5BRaHQvNpompbzp7sMToSSSEf
W7b+tn6AUC5AtYudzep2nyW4WxVLFw6N7atK8LFHhTSUdeehxpVpBkwxmUd1
Lr40QgqwXNsr+0DD7NY/6dCjXL9kln7TKq95aix8GEbYEf78v22WO0MHLprM
1sNSTgUKClEQLFCgAXIBiaZ3NKaS9Uii+kYpcTYGp58XE0q+THF/KPW0LFce
OWDf7GlvsouHevIC3BDMy7XyjcmDm5RiBh1PRo1Ld4V8OTX0R5n1H+2EDBVt
ZlKtfGEsiNnCIDoUwKK1Cjbej6UivWFrQVxq6SqTbnCAuMGw7uMRhBn5D9RS
gR2CsFrTzeBHVwv7fHWFlPqz+MecYJNThNwHX9oDNnlV7hW9GfCD6AkluWqg
yUO5loQf6gvySD9709Sn+ur/rDY05gfgZUs34OqQe2Fo4VWJCgtHDEYlHz8D
GLF07CJnPRmeR5hsqQBxfKZfsCUq/yf3QSqDvCri4DwNhptBA4TCDoCmq8fm
+Z6p37nWCKpR1Mu/Etajd6MvQdTX4/+VloVN2Cd8Z+D68vcY7HfxjlCBvZxb
vt09T4jvwaiKKUcwgrykgGk8ZQz+1n0v9XhpF465OHewCAfPVYEqr7K3+y9B
FwHmcK2AdXiB7Oz7UAcE9lMvlxy3WVro/KN1hpNp4hNNAlsl1TwXgAkfxb8S
fkSpWsTe/qa8DZs1gqoOYoOJKSAaOrCtT/MRvE7scCttOQ18lB64wuKAy+6m
ookb8cVlwd8oFsm75xy+HJ4ljYI2yH4jVSg2NYr6hJHdL/belW9DABexMFHU
/wh01INP1M1mN+0E+YbztNW9ZmoHiF0A4DV7ANSBiwaf+oqJNdaK+4v8SYI3
oc57yyaGZuVllXY3KUtGxf2Df3yhI/OKTGb5OWqNRNsRtDL4HvJ2y08/VSWE
/z7vxToTivEGFZ6LXpV+WpfHBks8/II65dyURufv0G8UPOuquTAS/1gmxgse
+OqvaZsXiZsKAbss6XEvmA+63m/2e4h3DeWXOjE8Yck/CQAKsjAXDm/gUwQJ
6unFWSpXbbX8DzgyFrqWeCb3VBj2+dbrpEM7lznknNN+lcy3VqLTvtoh/2Lj
dMlwn2+RppBYKmV0uoggNc6hjAlRSsqxApo55XCUAEl35w6ID0OB/h8+5inS
1KCnTFTE6B7H1n1trCHkz0a1r/0WbFEZu0L1YMulboE74AaDkWpZy3oZYrkV
VqakBELuhc/nnKhMnEbe0D4XJ8UG49lc2kwhFD09edP91WU3ZcWl2mMXpN2m
eXe0TTx1wt3Qa9F57mA8L7O2R03W4s30/mi3LH0e+9gJ6PV3hWlg/TuJsSxb
4zEJ5irUYmVamPSvdw0kJYhO22a2lQA0ILBrVpfYHEc8uDk2aDLAHIrYXLYe
864fv8ExDjZYsSXntcdDnlTbGZ0bjaTW6CzfaDoLrH9W282ZmR9KzAt9qErO
eqSaKoi8zB+S0frIcU9vUt2IR5/KpVeGkMK50862MXfB6MypGPIOuVEaniSH
wNMPQ2PC+n0ZRXAhBB+qFLhFh5TORnKGU0N3WBw9AUnLTYBUsdN5+LAQj1Yk
dutaUDHHcTHFQfqXDTBWARx1a+TqjWR1n03m47FRurKjvp9mwJBBOaUuBETQ
WYograzHs/iyxM5LvTgLO81i+uLwKbKmx3CaFG1OGKLz4voh87qhpXIJJ/dw
ELfUyJJ55C5M2OC4+U8Niy/6BJlBFOz4/GiaHfliklK21VEjabNDjEuRt83r
cTxU0/GxHegPC0iHdNzrZHbM1YE85qKqHBCucF8aMKr0m0RB4S+zpsJLMqic
UWnzJJ+C/cZ2tiMdMDRTVoI0snLpr3bh4Hemvb1MNbE1D8+h6DctbtczNk+U
BroMEMziSmPLiP4nIS4aFzgaUOxwV7lhZm9j0JuRLO/+uXvsOuuutzJXbQKl
JdgsWyhMmPJ+OCSyahVfor0u9DqTinUymIM1oOaACTRiZeZ4sHqPaHLECjU7
stkxIg1tsWIV6D0iLLs7fHpk9/kqhfTapwOLKdrefl3OZWSC1JnBwhmGcIbS
OKlmvPPc3cPyS0Y5/ewktL/W8QCEiY1Krrof2Zu+KoF06CvznKbinAMye6S9
lgYCl0bYdEsqOvn7Ju/i+3VzikVscrY9PX8AnxeNcedwDjnbT7YSE8y+PE+L
6YfnFyrtNF2lX3M8NM0q4NyIF9kEkKBVY0ybauqpw/iMbCsvL0jkSgyOLcHa
Pr7rcUwu6zgj2GzGKjpeb/Yf4SDh3Jw48qS5mbxVpoESknbFWHqeIswmTNbg
Yyop5k7rRj7UwSgaumT7BH1j7KeFW5iG/X/q1QIZh9j+KrnmIlNxva8GwFhi
YUcoDODlCON0rAmYl++7PuXTpMyp90HkcuagP+dkr21Prz/GS+pCcl+RwcyS
+koFuUlwRrSnN0PAt/h/Dy6Z2wfRGSl/xfQSKU28A/Bj3BOk/Maa9669p7Gw
9xysZW5KjEPUHrsKZN3W/b3f8PYyb0/DU2yR+LnnqQeGrqXMF544mmvwmpCR
y6wKY2oswEwbUzUakqazCAWPpQj8nmBwL8f21XYfkINp4kzoIzSXOa5qGiAe
ZtmQ2Gyjk6I02HyFIVpejl3SJJNeJNFjO+IbaBlRC5p7dClZdNvuYhASnAjd
XwuaSTQqj78QyFXWzS3p/FRuKOaTuVVIf7hE5VIE0hscL/dHdAcFaUgKJ8BM
HOmUR6ZcgsJ7CRkE/Gl1xBBn50bNAj0KTRlakgwl8XIOBpJ2Oc3+nf9U/jDN
2hBbIMQG5O4ueS/wAFUVLUDkJKtrIwePAj9oUhX+suU4AtbQCEYeMmzK+gxW
9tIMn6jDlJQ0rutP+P5syjJC+3Turc5VD5miT5IAMch3ZErHuO1HSDluhR+J
ct9iW223/l13KzwRxcseWOd+HxPujjfrmDgjj5TATlmaGdvQu43B5hzvsRhW
uzeo0MGtsi148bt88cAVo3qTvFrEKOH6dm5b/QbdNyeUt6hauGANNNfRlElA
3QFfYqYh1bAKn+iEo7jmH/kL5D1WQqyx4KwrZPzSEMrj4xV13KQojREag+DI
wbkg8Ak69YYF+Xr2TmAporBwaLuMmjLw1F3W6cgk+uM0EI9dIg2d9MUvebli
0FlW6EmqZFsnX2mLOH+Q7PpCz6AKdn8OLyQOMVaG6kQGq9E60vCB8gP0ktyZ
R49o9aLe2ZKAflYVSTBQRZGJKMVCoXihlffpVkmXMhdXbi7n4DtIu7Zo5T4L
Vp4ha+pk09ADVVNSyLfZRkK2qFfK1sXkODoA5633CmczDyWSMZm/YZLhn8Iv
qsYW6Gj/VxNM+5/yyp/MHU0AFu1WnZ5kJJNOFQCgQPa2/ox7T9Su+H9pu5m8
1GE07WoLW2ljaOZ+Z4KfRqdIhOrZg98v6eaaglvUXL6McBleczGRDk5M1zUk
TlyACG00z4g4zgGwiZB65rEo01HBa8OypCbglwlIvDUjWsy1kevmOUpSxo2b
pjACg4Y/539QZlCtowO+G3ghgJXy9VtcnBEkdn/S7EHF+C3XQ9yyNE9zJh6L
lz77Zx+LQJujcL+AlUNt5s897WshIKtUfgN4j4vPbk4s+Z9k2ZS91JMK1wlW
1vRUEs2ZRlT/S7pNccyWsHbq6b6dvXz3pL/Jq1FyqH21NV4TDTzQwNBG9Are
rAL3E4ojyW+HKASAXzhFzEfzU8Tb2RRFG8+hcXxpgIBxYsM3UKTfsZWZXf4d
wQPpmnPGmK7fbAljv8wIvDn1ODySzQC10wQ0XLaKluWk8lYQUmguHjpOSXlh
//v9yRlrDrmE5+JPH2zfX5jlXBUOuqWc+6aAXLkM0vsXuHZ3BAmQmSxZGu3E
ZH2z6u5vbvt/5IfXx8yOKUNgGMeO7HzilE1qi9cZyD6fQmRxpSmfwOVO9UBM
Idh4TTwg2xQDXYPvCuDcdCopfPO2Z5W/E3Ci+KydU3atjsV1Ya9E9AifLhIa
bpA+OhumMrOI3Um3M9WE52uCZY0DsqOl5PzMGoAjnCC+rMcMrbd9Y3STwj4v
R5cIuQIytsnZM5aU3DudCZueuJurIxHBMbg33kBEBiLc3Xfw9BoKqO0k0eRI
KWOVz+Zca7jyKooTqLdTQ6H8kVnlxuXgKBg4nPpMIC3nmwv/PYzSMjR65Qyc
ajz4bzSDA0Kwp7O9wwC28p8Mn5X6wVl1m1ZHjqT1iAoJx/zxfOdLiIRLa4bU
b1dwTVCyY3s2sacRWRGe4T7Ds9D2DiKxOAtxtKqqQRtTUY+bdscugs8n5poy
Yl0fY+Tw3RzRlMK/ZJiSBAzW1ESIng7yjUuKAjcuagPu97m58kuUJJOw0Ldm
AOaZm2733FOFCYxWJTL/XjopFjaIeWQGoUJqoBdoO0xpXJUoTv9vbAVhmmWX
Bgb46aVqsi8i+ugWoW0MrRDVKYdJ9bDhGVjMQaQ2d0cDZHHj/Wr64OxoKp91
xfGBpwxObY5ebWziJ0tW5OCbLhDg2Kk53PyRf+OH9iQqM/Rfde6rYLSkzq8i
Pkj9R02NvGDlSdwbtG0LZ8SUeQii4r4ZyOSuSIW4aZxpn00YZ518aJxdtzqV
ckp1tmVXHK2azIZF6OwfkPH6i6XoghqXyA3lKXg4/mnRig7CcTMawdjdpJpz
KkFZxt/kj57Bbr4+3H3AB/2IjOpTPoThLeigdLCgY9oEjWN6AaUH6punUOKM
tVIJAr0xua6tjPrME3/e4GBu/pmBRmGOiSHmRgwEhJq+YyBtHWlX51BJo1KV
QDYE/+OcCjMoRpwruNlRa4tskLVvcfjzq+5bKQSH1Sq1GqIPlkU2Mo3qQrY7
r+gOWrl2WS0y9k26gAiGV9JwIhnC+Lrafn9APxj2OnfqnMHGtq2MC33KbtIu
iQRjgbM2ulp2okaqeLelPzEZKYvBGNJF50xdjMjU+nvia3VgsOBTnAWQWtyM
ePEth0Pz+XFj7zB59Rir0ukoqb0jg2KA9vGmv0VS8dxyCDruk15YvVf2jRyF
W9wF0u3BE+iFH8hB3piO7JqCt2eaBIl5UYLHWzIC6L1NS1t9LZ1dkdJgZbyf
Wapyf4xeY+8OxwyPfRRsCWFc/YHRygklvZ/rEwHfkJFv5ORHhiWwm0ZthDxP
WjmMpx5Fa0eCeKGIwG3itz1D5TIugO5E/uruny5QdyKfETyTScgg6QU0iv2H
TJp4mlsK0UMc/2RjNnPZ43fSvruBpQyhbpb7IC99ciFF7kWF0fDy+k7UdCB0
kE33m2NL0GkNxhewyaRihV3O8ts1sG81vFds8IWEFJ+CJHTv6ERvFL6HO4I1
vcPtLHlJuW2KOOH4PX0PJAnCVojYL1KaG6bkFQOI+r7sxhlQNx2YHnsxOrXj
gKrEKT7mT7ef6ITsz1nnxD/5ECzTtbzp2AxyNGu4wz/dg01PPEEbF4VvY2i6
qPljYtAK55hqj+rlpoNGv5GVTNhsxiQJx9WodLjo/vPXLnzH4C4UmQRYQQRp
TPgCv3xXtiG+3RokeyJzJTA0LS/sve5U7+bhLc8et0ybjULWJYOpXfeGpNW/
B/zerBFsnjn81gwC7pnKpnL/oCqrhbv928Rh7BGOtGMZ+yE0LkETWYRVv5NH
l41O9X26A2B+xJFmvCZqBJHKyMIm3Y/weBXmYes3qM8Tu3JRaxoSdyZnVeLs
EwpIJ/ERyqDJpzmEjeSf/mUDiWtkZH4Bj2GfJ9ncqgS5yfIYMeWsrmz3BuPZ
SAGHXtHixNHqLnkdKZ9HXURc9PW/pG8G21BacT6kF3vc16zjmuGA1KpheNPV
OHYneDwZbUTor8U+XvTD+Hac6JockwqNjiZwnOKHxHReDFfo0n0nEgqNPD8J
NjXGh7i0jDeLycz50cj3R50FztlZ4RgctJcMbJUNSrfuBpOf7KTfUi4mWEy2
YnMK/qPsLFHML9mCxA+ZT5swpk/owgWf2oP4Wuv1eKg9wUfiwmNgH2nx3sS+
Ev7Nawis4In5VQb7QEvM9f05PAHpfGP9cbRbeN9X4yjqM08Lasgt+87ov6tI
GK+yeE8GAQISMHBxSueG3A19DlRFbVtPpuS0H/o5dIZGuxopH/JoBcLyxak7
T0o/EpQG4W3wgYlt4FpH4WobYT9jSDh5/bYdERZOlaKqLsYIyZaj+LIaM2if
lAf5xGtdk1ZyUaXf8XFa3Rhp/sap14IQ/GTJQ/6p2mZVkQxDu9CIygTTZwkN
DDdXSxsa5ecEaaj4OHRPRDriik5LU6Rz4RfgM7LFVSzwvh5DvyuB/ABYw9t0
mcLI1ltlTO68ed+h6Nn+BQclvhw0kZKFBd2vQQlSYcGgg5beUl23F/4RfBsL
R+G6x3+rnRQ9PgpMtsxocKpcHnCZ49No8DYhEfUu4D9BF9XLYzP8alVWB8Rt
Ek9SFhKxWHddQjQqGflExG7LDXx7WUKQU8vlE3NN+ohKvq4DRURb1ilXYIo0
ToEddR9JWpvhcmIyhT7DbMeZUzfLzOdB9xlO0NHtKyRho4ABLLPbXvYNX3/d
/FeuthLB72WrQ3Ne0t8VK0DWP5loelLT8ZTFRMfGGEaDzKzl/Qb+vHfUaS4t
5vDoo/kXd+jskfXiuUyqNAZb3a2zXhSEWy/ar0t+VYFzxjbfwwTPK9MLP1E9
5uBuq97+paV1ieYC4oi0MsgYmL5gIpkXI+mfJbPLhmePv3x0CKwfspk4G4qw
VDe1/Yg9UQ+sdwA/LHks0Xtw3SghzdnO3kAF2LVW+yTYrbH5iHTiUnDFTKGe
gZp7LLhIfceBLrM88eLP3BjXePb3479LV35dabORuAQp4brH9s0qzGs8rWxX
vvSxYDRqIf4xlK+wjIpr4zcfD5g9zogI1rINvKVksULMOHDO2FMa9fhNIcen
znwDquvmlB9VoBhtJ2yuTXjEl518eYfdL1sfIlFY4pv4bhyu+faYAbt3kSd6
/qx7T4nU+9c378RUg7OrwpHGTv3KiKNgm/47tli0QLBLq7UuJI2GUZ2PpUSC
BMWNRErRnzcThNjVwthxToDqQrRzo0U7tcHtXq/+w+uI6Hzq6IwvN6VkxGnB
JrXavz+qZDimpiobw9xCZIcDBcTnV4UDqjBv0G9lu3kBqUKGR6WKB7l/YclU
RWfyv09FjwQLBMXa2wjy6i+0hU0yzAIRut6T+dU1JN7c87uUf0Y+7glOd3U5
hkHRQRCirAH8yqz1Ab5QiKZAF/Vd7rYbboyXb+Swg89j1X+9rWUsrn7pcFzG
YITCu+EoGcRxGEGhoSkmwiJo9RZArNfLsixiqPTSWbu+gU3cSTrgb+uN12m+
KIKYRBGKsahU1g2SuPDAgZda3ILnTDfmStLrtjmoaewaRVjk8PtIwFgNLTPR
kqq4bMyqtM0WQgLQXA1AOHWgYHzMCW+eRjWEm8/TyRGJWKG69Bh32rwZs180
ajIGlvOdMkw1qsK5P9VjsI/8K+6I1sL+VP1qr/PHBwMOLA1opFdZahSv07rY
T6VAAxZGnfoRUsGKyw4eug0cUXqv+glyoGwOexotNSDHjMTxnTuUwNevNzJE
nSBesdsMPXlZyOOEVK/Bgm1x3cBFxOHxH3LCfBpKsfYhPU06iJ1a0xIZlmz6
tKhYEIog/PSg7qpW6l1I6i/RS3NA6AjfDwbB5aIXtko7l5ZQe3FgchTdoZLH
8BveOzRdF6QuILftuZ2E8jKR6C96zk0qiIjTMlbXejSoforYNo+PISpFaLtL
7t7DPBEi6nirHHO1Jsj3up2CF84iAZ5Q9rTvqxoBh/SXLnqR+RxV3egCk1m5
A3HosydrnVcL42EeUF57PSC5hyxRlNasmCDxeRmwFtRJu7smuIWlT+Z4ymM1
mwOrx1HJY9cI7nmazZ+RZ5PaJuiDDu1q6ebfMPuI6hECXghHy//SWrmF8Sw+
Lv4X3TKqstxbwB6G2wAvLv6lZwU/QPzIj15D8sp+3G5r6hS49pI2WUWDp71H
84Vff7V2NRNZUPpV5rZG6M8LN0L51xnxFD74O3Ie4Ldsx+KUhRdJd+vPoZ43
Ip3yOibTdLJLqxu6u7Je2omRfYkN+Qfdmd/9BM6xM623yGHEYR9Qw9+VdsmN
RCKK0Nz46x9yA1qBYmaUiyKVFZymWcKxlBXUzSvkW6xEYvTuftmV8kXDzY7t
zTyViaVCcWHXyY47RbuH45J7L+1oxAjJvpv5ePe20QNRQvf/YnCOZdHr9/yC
QLX7mztXnZ3bYRCeCB9uzhlSA6MF+x6ctGxPko0I8CrZ7oqgaIhFGfbItS/m
qFdHQ9IdypRO/awt5scblF1SOxyQ5X9NGhSAnpTyfcibgSWb9z/fA4T/lcrp
x8a9BQ07D2G2dhQChFEu1AancHKAiaN5a/gA3jZQJr1kUOJKcSVZN2yHDEN5
xqDGqwn6cTuLjrjhtwxe2A4wo4RX67NlYpYCHo7FdY4iX0pPRiLnWskFdv4y
lXvOgcNkQ2HPqUcFqcCZ0VjM/K7TzEHD5GTye47qvUGppyul2iJPdq8CO7sL
80nEomMBeDryuHQXi5DCfEUGgSZ+O5/oVHbPZ16n9QAd4kK++XFUGAhgBivf
HUFE2T1KI10sv1bvNH3GB1preaEpeddLJ40FoRsdrJm8EdCRWkRgEjYtZMEl
TRJNox2RcxjWnX+lvzgF6UAkMvL8XDhQkaD0wbxkdn7L4TQ5lo7NjCrkV6iK
CCHeJD1TPoIEa3PGduMrRhCSG2+ZEpv+uDogLhUCXUZHXD9JZ7FIRvES5Rgx
bFegBWsAhPfZcnbWD/aihs4fq6MgrL0ISqSTviYXn0m+7OKkzH1TaoiwVG8V
Y0JJQkmf+oqeiRYNlzc7rucjyeIMt7F9GKlQ9T3fZqKHDvRExiIUGSIk/WWR
j3VSuhf6enIs/h9FlmRZ0VL9pWtLQuwNMfNzwnK8FOGB9qcXBMUgHnftXbxp
GtPfblrY1oOhPHZ9nE7hFoiuw1rRjMoBRm/MghtHd+o31J42hXT2xDpzlzcE
9kjnXxjOJBeY3p/2B28NvN9C1eFbNtKz20UJv5GodhS8k8f2yhEJcC5K4bhN
me3ZYsL9P99Ta1+aKkydHIyZrlpuG7N9dH/4gl6mfUlxZvtwAKDEELHcalV/
AbSDCr8G1wItpr/pMahRyKN4K1CHKVsWxnEB7pJOKNHm+v6GbZ1SqGr/tFad
dafLOpaMepyoh5aXcqxKexBkq1xgGOgt6Cv4CSdrlHljqCdsLMCof9Do2zQR
ChdQLS2x95EoyXF+ADgkUC0Bb+7Wx0YqOorUBeI/V6CbGRHeS2kgD55mKcur
QqeNFzSZ3BRwWxtbv/LYVMas/NSJhRzdXEkwr54atK5R2pvfNu2SJwO19YEG
KPqCRot+FZlFQfxJ5FhZFbrLGeUfNFzsRqCFG+zmeD5cuWrZFJiVfkSea0kP
XRT4be3EaFTFzqEC1zGhAzSjnDCc4CF2PR7T9Zqy0xaloVig7SPuVqA8WgEC
lYI4CPAnKRBnvYElPVNsNEXpsbQVRTuTDZLRGRSraUZKgRPvfyeQAHxpkKSe
nMNS2UkdiwYybmjr9DVsumphYmH5KQ6ZmXdQNXrnRB3vjQsExGQYScvpr8qi
icdl3XoA+3THrD8hi2Luko15ThqQPz2OvhRgZ6lKcPubY1PeDoEcEXD3iQyr
mj22RhmXiDKMTVlNAQcCew11wpSNSC/mvJGykQTZItvNuWU+eX0Fb84xOYO0
85L/UAuDOqfXetA+xOAf0pMeckrMsBs1DORrXQTF6fzJqQl0kml+VIZqn3SU
BSi1Ol/d3/TQV0fkk5m8P0jqorbE7EaWS1s04hod2hUHoOq/3plk9Nfb7Oz/
cx9+G+KkEyey7iXNMFatende0Ua4wtt7FvuMSnnRNxvsaqqHvB5P5mYLkXSa
6RwfdyWif17WS9uP5elh8lvOMxKlijpfurEWtJ1Gh2wOgl6v/n+4e1y4ayb8
gVligZaw8IQjyYMq/pPNcOPL+luG7oxIJnKPodSuo2IhhfAhoUZOQwDzwHwR
JDay0DC4Olpq9EVg4U7KahtsfVkmHvKz3RiSGt3mTymx3t3s/Hb35OZV6Hka
GCpZ7K88LLp3sGkJ1/KzbbZJN0OW6cuHK5/dVtE7rOwSx0IQJx5L9paE1Wfa
CBlS/vsHjnhYdizHsXIEnXMCnV4pAl4pi7t0/9lTAQxuxNOckCL//pgxiZxV
2Mxke52JsCo7pKt4hvfElxQaO1q+UNs6DbrF5pjHmlxT13RS3/bm8BwRSLUr
ziNEw2C1Lk50bvB+PtneLOuR+X8dntibRkoXa249NiZofWGcm4XUXKx1VrEO
ESt4uzAj0daJ6flbiwfN4BgjYNr00i7E3gI1o51pvkY1/HynRcAXy5ws+7Wc
ymxCIKK41Pi+Dc8ukOJwky866uZxa59KeFgxobGMno5/fzuQD3Ir6U/1fq05
xnM562dJaaR+rPu7ISPLvAsnfPrjA6rMwRGuFNWWYj4rCqlai8eWxqqnsrV7
brp5xE520LQapdw9YO7a2bGnLI3a6zIoZvbdGHF83sLBWI6KXTTYVqPAr9ow
54Dqy8BDCBbriLS7iMgsxIsT0p77u3ubyO6Twd/rUWhiSfdYMC+PhzQkQlKG
L1BnJkmypDc6eha/YyFo2nsKb702zsY4sI5Xi6rgzaTDbFSGQ9S91sCOZ/p+
RlLXv0Ujr04kBx5cGYsfoHZaPR60kUhIXwQwEfI9lDLGflhqknNzUwBba/Ce
3VqrhRI7OaI/DaaTJqHMaF0VFlKXr+k+Jy4Q6GjUbh8w7qE74uV/Rasu7+fl
hhnKEVqjIU0wV+tJSCxmroiBQmkHA1aN3HkkM0OxgyUK29dgoMmO4Xggl3CY
TGkCKU4kr4mj+Z+kaAyW4e0YDRyVeKtHjD1GYQElhk43cZuXGiGWMy7NqjxV
FXX703e2SCCmupKCUnkEu/VZ8z1VHEFBzxZL9rL40GAWb2iLpS4TigzoAenX
PeaKT9M5dJEshZy6Z/uiEP+EM8FFknKC3x4TpQrwWQ6rrWzhln91TTCLDrCt
ha+w6OwvMvGS7WZikhDqkUtjfbXxfVKBrcM6XG0D1fZwbRFcU8iBahecvHdM
gqcAknhmhLEUbRnf4qZNIXa/n0K6cwqIWpePJ2FErqp1OMhJQ1n1kxtPrMfE
xXcQqgxROuRlZwTX/ltJd/ekycE9p6KDWUqxC/962Ae+2xOAx6pF/PqLS9ur
xtnHT+UuKg6kN6/YpyVlYWKz+j3Auvh/pPOMnWLZQ6TdjBQIHK03ttp0dN0l
51OWR1oF8yb8g3KDq1PcxK4X5P8N+jGoF2Uh6coYU3Uh2XUNYT9Uy2rv8lTD
c82szFFcKESyd4TZUYpN3sMs5ISJzmN50REcI3Dr/zQ5CXcgZ4N9vEHx0XJK
CweE8NG1103BA8Ao+mxj2h7ebEf9bRtTt3DTyW8Iq2J2uQDcRUF/37PBcu3u
E3UaXPTHwoEAniOyQ2+xC3LR/ec7+mzN5Kxgy/hjTRKwUIYNO9qj7BlBFJyk
yE0pIVghtdtf9s6qW+nmbCDAO/oxAzT46HVqI/i8zsc4c3d4Zw+QBRjI3PFu
A8frELD2wGDv/rVCIURif2zDaomKV2+t3r6zhXiVZO/zKKAs8PN3CAEzCvoI
4fju7Bla+9b4qAWfM2zHTk2KiIHkzP5L1TPT1/bCAjfa38wSrI0yAd1/PXv7
7phLB7QwhbHfWD8vHuI3V4AJ7Z3LB6YxAYZLvNkQyH1BiIpZcCLKrrSgC9xa
idPaM47hEMhJcoQf/18hm7ZTdsgj0GE9UTqNbK2+97c5CNr/Drkogkw4ALZo
NM2ahl8CEFrCoTHDIYhi5KWtqQuYkmpusbAIITseweXhdqSd8A952+Il3xp/
lp2acLmmYB4KCKPH25dcp0brh8CYI9ksnJxha1OK+COMJjQqmZt479onKxL7
8hTA7pETacBRDzlhujIOELo6Ws5wkMmSrcaADvWyL0SdL0mxxcwvAhCew4QV
r+Q0dcdveME+ypI7RwvBj8vQSw1xZpqnDzyu6y197rUH1jOSt+4CFJff0kSu
78cwPkpc2kOVFgM+X68jhyd0bV1pe/5psJws+Fz1tFuG9kElg81BKN234xZb
YtwiFcaG8Jb6oz5b04DtDS753tvcdjbC6uFX+SRd+xw1M2uxiHprOY0GBCBg
m0sQEQv6H8L2pq1Jn5puWYFnm3Wf+pT65/sWSoV3lcsB4dRfbJHgUcFwc5Cs
SiSKRscITH65Z1V4mmBu2Wllz5vELBSk24/VtIArstOwWA1ivm1JkoX57Nga
jm2dchvlTkBjvsVmVUgiO9Sqz8YP+DXh8rv5qZS1UH6dLOfgAWgmkR0R6rGc
Z6ygBEqF5xLqRMWcxS342YnmcB/EYKvCUIOAz5QWvv7FTWMjSmJqWD1o+fg0
Ohp955E4x8lANbwT6GP4kZHhFMc8HceROVEXZdWsozSKWllyIBLta9uZ+dIc
cnXM3nLakVF9h557OCTExDH+KeueglloO0LvIMDzAgX7uPop+NAJfELWkEhG
IjQqKqWkvfXuJJXX7KC2wMO4CJPg8OQuuPN/TsgSDsuvHN9SQ1Y2iP8WAJOU
Cexka9U1TO5OCSz8O+yVJiDv/XE0jA/eRzECX3Iz0Ws7QOJBP+SNCwO5yZhm
gXoUBW6GWf7r6jvn8DVxJ+XYhFKx56yYB54fAerwlCb6W+S5csNR0MtRMdU/
QiRiRdsgh3f8D26ai3t/JjbM+FGv1jKjPzQkv1/gomiVjLf5EsqmViX8tJfz
7b7vlYkL2gESf+U7U7KGqE75IrQ/duGuq1Ev/vZuZCxhpvxwxJvVtyDpqcgG
3DdW4Nlghc4902fDUhebPmpOm+ghhIaqPQELVKNUgsXxSO/1+Zvwus5Z29ni
UbSJloBLf0e4uJniXbjrCovwhLzohUHS/FQlhGhRQyElTQt4Sh+f6exKtawO
ds2msLUjhP2KbXElcXqUIdiC8tWh/QELwt8i0vqe1XlFfafw49ON+6tdbi1u
Y7cA6ORGAMf2x/IqyFrlT4aZCWg1j7atj4QHIzOMHGjEl0KKVs3w+VFrqNv3
oPBnBGzVMZ0eX13Ku3kQOp4pmGbobwHOT+6NCPiVeJP1S8MGnCTNZn1TX6jH
vZHcs+TeRTIxJcvWbA4aDqo6wGnkvVcZMQzymGEIetSsh4hvXm2kpG4a5bda
1bzjtRp/97BYVwJgChkNRCGvei/dogoYYXOVOgwmggyF9piL6mfz1m+yaRQx
SIR5rOZVJrBtLs/JdJ7dT/EVZtBv+Hpwi2+NOQrHXB4L6rs4PXn25d9n8I34
D2sYufqDJmWhntJBOWfoJba53Zw5wzq0wrbtwIy+qvqq41CV2aDWbRWxKmPn
pszXFoQ3eA3GAODton8lLEODUkxrR8ai4q2Guk+ZoUY58C6jlAKoSQTk4+ui
p3Pylh/DoTS9hNbWKxX6acN0nlBdPR0RzeP3/JiD/8h50/2Cb9aUAmeX6SpB
AXvLe6nBOJ+UcfgWVejRGKkUZz6w01EEkrTcXAFrJ10wxwhc46UZwgAf0nuq
ryB48RotEcJn24K9j4La+Ns0/XRdu9psVMgiTOIhL03Crf+RQLngEXkcqqDi
UtqxBGvUjXvSa8rZpYmVACojVbXVb3cSxddz6L8Oib772DSypiqOiUM5cY6C
t3vmlwRT/RMSUotvz7Wu8LoXB75+Npwc8Qx9MjQmsXUR5iL+DtXR1kzDBrDb
9aP+RpNRl04270rF1xYTaN5H3MlopI6M/BjwxgVgKFK6jzwgA9qSTs9tJIox
UEyIvIVD4XVpbhAwa7cnLqAYiG0XFe35xaSkycKB1BqK7Td+6TWB2q0iZR5T
+wt5b4reqayVGQcf2dEap/wXtv6cJpoHTPLa9TL283DYVluYEYFgp+oKGhNe
3dLBfZbwKmWWhhHtX28DwP9laqNt3cPffZpllcFD12u9J0f0+1H/Rv6JbQpK
vj3Uau0D7peyLOg8/OF72essK4bUBa9rNQbVrypSm8OKPfxovsVBniKPlnaI
qeLmXJYAbbeGd7L6qCTmjHHsVgCuOqqtIGCut/LuIaSLRqKAwvxak/CoY4pv
JgUqKHknU3NNxfV+MAE/2XlwJs2Mj0aStEF/omLAo752UE/PCNFCHcKNyrB6
R59fso051WqAvzUY2HuxtRS+zr6epUm3bR3Y0D3aL/HQhzbgPsKmTMt5rGlz
Ufnw1CleHTNJq2jMpq2nK+5E3tneM7RxjI4Qazk07ZNzObI1L9+BKNE2QkrN
4/HXia2rthx5sGSE1WX+i5ZHdFS8qFzz9dsWAn6lqRw2fYftIFx/VMvCgutp
8lW7DRrBbcHiRExtFdhUorYp9s7g0mwT1wWrG2Du0E+9UmpRPNSkU4WMNJOe
9Q0VRZxwS0Zr+T4VyqidB4NtXBamUs6mr2CTA0LktbqQaqy6Bck1HUYxFihx
XWkmbj0bUYEQqEkXc3fck9bo1O2846hzAKZKM1Y6Nf9FUcLHAIkVNzL7zeJn
k0lozIkW21HVRugxKCTcwaj1xg4fUqqdEBQIxRnRETFRpRfo5QeoH7n2ygel
TmQfRfasJUuQOqtCMVEP0lTikvATcV7Rc7oZd3x608433tEa3pUy+Ks5zPwW
7YIePfON1i5a80ZsXzdk2dUdeYbhs2W30ybV38CAPz5ANBafru9p4Aj+n/5X
kW8tlwED9wAldYnK/FOzHlZZs288s53vtvWOu6VooiV2Lo1tvPcTfqFQyTVT
fThdwG1NHg6H3Mta1BP41wWGYGOu+fKJpi4HEFwV3e2HJzLRYNcpMPJOejRL
cQBONCbdupXSOGnTcpNhwmCy49R0H1GTDco8Jq6rXQ8NH58uuTTnvxNRPKk8
pC6E0q58kS48zPSmOHhf9aO6UDxjvltH/RRaXjYo46P4c4NQVhjtCyYQs5G7
ZWUHR3z85cDL84hk8s8gMiKM7BHnNxYelx3zBd174f2M8438vXepGumwMIT1
AfCCQvs6PKXY0A4pFWvuRP9H3joZk1oyHobZuSOzpTpiw9/7fcVQGA0VKZW5
lfs+zpjosoeJMbY0Y7Vc+Dg5bfUwOoHUeHqIon9iCL7aMUJGT14bWOYfjvy+
wa3jyIVHHrHJnfYBQYN5Gu+P8Rm4ChceNnknHm5zr/J46+oqhOUMXa5ULXSE
O9A0CfjEmAhGLFMK1miekKtE/VjMXvnZ4967F4Aqq9ehKxGx8zCbq40QX4Nq
NapEMXLDY0m/OvgK29HmguIc3k9Q201ozxtefdCBHjgKcVynU0HytjtTUgn6
bpKKKxiVVHh7Fs9MJSCfWlneDT6JntCoG9ewZtjaOIJK8NCxDTPtH1/4nZ1E
qNET0OEJ8QBAfiwVRg9HWWWo2ucLOraDJpeuesZLsgRovMkLZj5wTZ5y6ErV
MqlnlzWfzCDTT5kFmmpw0GDe4/vu1k5Gfn2NMPuULrFx/2V0K0EFxgFiplwV
r9rdISJnFKftAV167exmxkZkf8Vr18aF3uWt9O/TZbV8TlgmMfwdpDHfKOJl
iYRg9r9RIj+0FePfZkCDFC80UnNn3DRSdP+V+HEzo/mU854LFGIUMvkc64zV
oeTIEvk/0/HSJ0rzRzWe79kaLk5uhZV5BBvbITSTIRXuMO+EqOa7lQl2dIyr
fprsojUMzB08s6n32s4WL5+yBIbWOTeV0HMmUkcxfRtda1cvT03SRmQULv1Z
/5064CRtXCAgd6Rspv7BKF2vwXXCVYbk4MnC7yY/s2BDEZnQvjoNzC3WVmCm
Uol3R6LUHjuTEig80cH2ZOORae+Dj+FmxLqU553mdh+nIeumRnFxyzVITI41
KYQWO0zICboXd01Pg2S+88gxxMzdK+N/6snH+5ohBuf835vRyvqZFFHjwwzy
bAbFJtnaUN9VvOqRJVwD4rxk20JHz73HPQmPVkVxOvZiWNCya2uiQE/FzYm+
oaJQcVVXdIQx1EpvG1WWiVcCxmDbEIyy2NHUZNUhRdVHy8rJ6Ap1qnyYPbcZ
0wVYKykyYCwSYDA0swG5zniHBFLMiztI673avEiWHr2vX8mJPBdHyNVj3O/b
KW6FF0AQehIEcXG4gqaQc4gq4yEwC3oLIjBt87SgAgthSib0+cxxx0v30nIn
JmSUn/h33TSa3/XOyiBBHt/4CvWhxLXdJ9bPVCGQQrr+ZFs+uyKvI9qL3tFs
VHYy3jOG2E9WjHstr5st0a9OFsJCBeRX3TnPVr0AsKK7tvkmY/hIZbIMyF/v
arXZ9DikFn37O5UVaGUihyNzyQfGXphwVWyuyuos/EEB0cKQDyvby+BW1KXA
vXNZS+oeLYppWg8wrHvuw+IBHU6El6WyQm+La2LSXHqda5WZQ28wciAUepzQ
1kcwJMFAc4GI2cGaS3dqSanv9xzYvfTsdCXPFcflcSBwjM7ztpiOdKGWdw/I
kJJZFrQJIh9JJag9A1r1K/QBaV3O3AkxYayWwB7O3qnsecRZx7ITZvgvwEtA
7t7lQUykuuDWZqHFcKR8MusTBTLd6cLECpD8iTMgugV7SCp8GKubHFF0JX3s
Ng5ElS9g8n83AwlCriyui0Tp2nJFVrbnda2mHUqOl5ayzmb8u3aoHBWM9ANC
FMBa3SWjs3A379YM0q5fUJ4hHpPRmlqk8yh3gfZY1jnsFJ1U/usSu4kVHFFH
XW+2zPloSWVjVWJPKKFSqHplEpGEEvRp4iQ9xyRlPvkz1aogOXiavH2WUhYp
golq19B5vuKb/XFthVqq0L3Z9YpfZETthmpQL81xoulQ18EmE8Iym8TuuT2o
Rncn4sBJ/854tsrWrLDlvquAM0/ygtOdLMTgOuoIT4mGoQhsEBqepcA3rYkx
qw4U4vP+P8huEnIqfkiurnWjmpllfimS5UUAwWkh9Nwh2fN9uxrpy8S+4BL/
M0Kj+xsIZ+YO5nQ+cmOeeWl4+k8SDOnX0t+bTY2SUztGV3C4SFOsEz06Spdf
82UHjBbP5AKzYWyOB+cmjyO2N7nSs6HMMr0mT5ZA5fMIx781iY+aPem7WDL+
aLAxpgWBMPq+QUqeqY43SiB7xHQftRGNtly+12b+Pj1PUBrx3SODInuRzP9g
JzI7oh0AfGo5AafdXjhIsr7JK3L6RLfB36HPdRElU+vFSKpv41u+k5Rlt3VH
ZceLKwqvYSoO5tcLA6t27T6UCm6lh4+o9aCtnez6gb5pgccLOAuULFz9mGfK
kH/zvGFXRa+V5e9zmk2k1GeV65TfD2Tn9YHt5eMqKWLfSJXUdf4MU+Zb0/Vz
+Nfgy1EF42oObNfUEisL1JT3hILOvEkPiSdM4sak1AQM5v9J61RBs+4l/+zV
JEAnFVXhrMMd15mSfkBCEpGtREAZZJCrrNNsjC+qD9D94W1N2++JZ7gMNpFG
yl2c6FJkmC2V0yFdIZvw7hbroDKnmFzvaSGYZIuKHfKtP8cBi0hwpsZPSRm8
bF9+AgP8lBmCAPkEpfveBEe51HJW7gy6NUSHahI9+UKKGpL9Pek0p4s3ur4d
famfqcWZx2+m3wozy59HZFeZoNVhw1up1PulSuC6TGPb8Xae7AI0VR6vmhlH
NAG+gSOlebjOY71XSrO/M/nJKbmQ+SVyR1fQ/fORDxpCLF0jdmw1eQlt8w8x
4G/ghluul4BOW/bT5AO8MwbUSDZamhzWMHo05VGpB4UiKVfb04niX20mYi6J
eFafPWbqBEZGBxgmbb5GxHehJuz+ftaXyLkbzkNYcKWYNc5rYyb5HZF7IUNo
KMeBRMuotIuSjfu5jIU1GYo6sRVq7op/Voh2TOu3kK0/c971wlh0X6jZGXN/
I3WgllYHN2k5lGZUiynzHc+BeM95o7pU5MJkbpaIOPFTWMGdPJ3uFoAHd2VK
jOTp0qCGdAd6ygcKatP0wRzB9QQNjwmdIMlofC8af/zhVG8nu8SGyCPSVIXW
95jRZ2LUGCP5/uNMoljUPyQFuG//TMvB6LoOdupWPjd9Y/dHsT6iEPP3xH/b
Kwz+n+SQzaNBjd+8j/IvBFIoaC6f6W9ZpQufOvS7qP2cOHPbN1JVa4gzjMpP
8R9dqZoXc856AGlfs8X3QKqWwCapLkDySaf6Fvm1n3bR9hbfu9ef0F5Fk7kT
nX6nOPJpC7IQ0jF+YZg2bGjgZ+ytNghrRLw/cNcXD/91O4TBFWVGtrmttUkK
VATP4eRtNA8FInG2ASgq06jsN3ZFeLTxk/pdiZwpjY8uAlOWVEG9Z2AEXbdg
oZhOmT43+nxgp2HUbkPYrJk1zy9AJQfkzvCDwfUyx3GrhMN1As5R+X7e9aLU
3pzi3PbUQD6FxSz1NoQ8m3AJSzeCkRvIDIIH2CKwsmPJ/Qm/I2vjJf35TJME
MZaWAyKVIfDg/wwysmm6ad4ahGml8GBwKdIUZfBRz1zpuygGbc2repOocrBi
DnaFYbBM160BxrTBihFx5UTCErxrUblpWfGaLtaq3f5rWAdxYws57vlI3966
VckcS0Bs2r2r6itWV1BIkx0t39yFUHvB06Zz9kCHh3vgFbgo+cS8f6Y6Fbl7
KLz5hQQ8uSBoG2rqxDq1wFiRMyL5315jXgkAuq5tP7Fn9UQfP9ChPurq+9vY
5shtkfONu9L93evqtiy+NxQ7RIiwBRSOmo6BfnEwv+XFJO+W/7W3EJi61KP3
KToVWWp1UiKqGAClHLvhz5yKbmOgo8X1ltyBq6/D6sCFn5a1pmVSB22Qax5I
Dv+qTBdKK/cOTFbkZSrFUFWsffz31t3rokH234dVGVtgA2b0M7ofvXdV+++9
u/rQjGxTtHOV+062XnXbRxOJ9bXAvn18xdfgaqnVIFGuJo73+6J2CR8lTa9O
/CnUoL7TQZD8YBWvN0yg5EeWm81AImMHh9LEKHDFIzRtEONrcVTLrdhZJ0o4
KJAyKNluZ8hSiMNqLdtV+MPE0xv1CyAjF6xdhAHkntiTLoFBkjh7M7/au5SB
SkNF5OZ9thZkzaor0A0QrV1GULu6PO98C4Fd/+uNVdZ4V4e8jy7Z66HZJaxw
ezGCL+RhX3l1PgfgXBhH2MXlBdibgOUV+YNkuSGXC6UcX7cqZ32yIxaP1S2b
Kodv58yodpLKxLGQl1VWX4Ts+d8SNmNnhLJh7uNPZjfcpv0t99DP0shVtB0d
RGDt224h2NTfqLQ3D+UbkIraCVt50AKAafupzzSW3melqd2IdLd6JkEOrpT5
FwkERQtJ7vE/2brMo1+2Z2lfyUFQpLX9VXbeYaTVz+jAdbs6w4snLaNqdTBj
DpVLTbJQ5ifVwpE3D/eDV4wEuWOpwK4qhOOGyc/GL96c8ESoE2iZv7nTd1aV
HzTN7MY90HbQUvpbd4JvTwlgNniJBLpPqaIM3DCJDeypHe0aYbNoz7GWOchg
AcovHZUNuNMZHNh2Ry1AdlvNxQ4Ev3ZLPRJjGY07j+53MjBewEFe9tsfbqGQ
fO5D4xwh/wstndJoO2AIM8bIFetYyavi5zS0Wy1L8uZhwzkzkgGC8Tt7keCf
UG7pxsyMOYcjMWvTpHByKb+bs4iDy8syZPKxT0bjEjWyn0L4KfSn1ft3wNc+
072nQ0GCG/lmXxQPRN8X8HmjysBhsNXljbTR3iZexEf/9HRrPaY4BhcoIvoP
weW0j70GlZ8kviZahnKo452tWf98ev6zwO6Y/Go+vKf0f8ei9x/mwzo36G6e
XFc75trPi7KirXVa3lKujZNou3A4zRNTuh/dhuoBr9VS5hX7kf7sflpZSRfs
ZKJBIUZGpJ8XEUiUL8k9rTFWy2yb6vB4Aw0Pa9k/fjFdWxqOY/2hsFdRZ8dY
lyhgy4r/Ya5ZwbE9QlLgLbji0t4ZxpPsMSWCjQQ3nrKwCHCx6P2mDALJv8Tz
5I6cy2S04yriqdZ2ZADM52m/5mJPyQExYXUa+l/IcntUskhTd50KSH1gi2uD
+WA9rT/GYdyFMDev7WsBgVZgbsJtGYP9Ku3Rs0i+JaaIYv1c/qdF5H6Ke+y5
qWlzR3R5vAiRF4MeKEvaxGloT7q3xtcQUEXRkGq2AbiPtIPLwLWZL18+jMWI
xNlRzi3BjqnncjAYmKxRJwgsZgm8DtBafaYLieJ/2wAJ9f3gBpRwON6CBioX
7vUBzISEmFB/q6kWR1ZFMzjzZ52gTizyj0jb4q4RHV7yKhXcn7X2Za8jHYCF
oMw+2YAf1UXaO204IA1jCT2+Wqzxn5K2mntbyylTTVGr95f08PLztO08LUZn
2dWVf2Q5x4PiYwvVSMODYgpGIuaTXfsUAWqwBP1KwX9ghb979ePhOvdNooFW
eSBl9BElwnyh18zWcvYBqiEv0erUgUn6rF3VJFDzwLiLNt0GEb6yg3yWHVX7
Fhasa9SZGczPqY17GnqKSZc6aKQwi1NeTo9nMTzyY+Y/I0T/AqrpkP4l6nK4
EFDIclyIFkGb/7G583BHPYo3m3WXbD+16b37P35VUrILr2w30HjJhALogAJE
xXouf8r8EFkTacqDbCVjrA38FEISBs0CAUs69sxP7ZVfNYMFiAaqE+15dY8c
wnB1JSj18H1/WcY05QzDCnpp97nceBH9cyulgcmptMFFkXqq1+8YoVfWcJY1
tj+wL34SaXLUegUc4uJQ8ragcoDmO1BsaD/P7MPS/ZshEJwz0tvngn8AGeuL
9Zj6RUKkTrAGH2LNJu7UavSi6Wl8rDQOJrIpiAq9Z6wJ+1wf9D4LOnteFqLJ
R7VjWQ9qso5Ovr3wfWH65pz6f0RDgIF9+HyJLoknivj1ZHaim+2gGP34N/dV
PNqQeTpM5PzgDoXfaYb/DRzll2aUPz6vsQ0enoWH2TkVeLTJFOOrklhaXSBO
K8Z6HZeVjWTGTuLlP7xWgVwNEfVoOr7TqqatXEkKpkIWyvsbtwW+aTt3UeYD
nUe4GWBu/99IhcJurc6+N7FzekJb0wXc2zqapW8T5bCtHnj+c1PYVSJliV/w
1OM5lTuCeCA5Mm71Oi1nma7/EMAYk9GCFKCbqtTmhMlH2vE/D8/6fIc4JmYI
Z6DrmNYHx2xCNy5r/i1fUHf9dZajX1XR4HJQcEpJf/yBiUjLAFJJXqRku5D1
aYxQ7Ha4B8cKkpvYJySIiNczG7re/CwtV9fCIQTgjZJeaohpGNlb376odFQu
dfpDJorAxW1R2IVcRm34ziZ+YAd8UNn2dDoOUYYNoySC+9wSCCI7duCGy1RT
5vAGNNaBmoQvxNHHNwPDTJte4VsYyei0fYkxSjT6QP1HjUtggDFoYdaUwNed
qBKaJqDPlQvM+WXX4gQu2sVK2/sXpkqg7a/s3hhs91qYRPk7IbxNb8zS/qtF
35BqOE3Jc8qE/xkTRHalixxapkysFNUr0STieJbpEfOPpvJ6n29SrkZk72H1
i/h8hRLjge411E2b1TsJwtZmOupsakNQIWvh8isbp1mUm3+ipO9G/MLPzsLh
eBiRuuq/CSQTwhQ5lB3MlID70CrqzgkDD5XGge8AjURGVMqN84CcB2WXSpii
ihskvWdAiiPaVdMudfYuyFZuz59C8h2KHREpGPll/gyiaP/soJL2W2Vmjqn8
kmwg7AYvaswUmTwlLawqBHsdLejIfS5lm5XUfDofy6aM/yusG9yihJLviG93
kZzs+vPY2JWCVnpJRQt72SwfHTV0jZQObWAWKY/WmAAknqSEn+/HCy0x0uRn
zXfQrWQIwjahbJfgJmwSovpW7znbY6jN1DEkGBAShmjvVh3K1xTQLgTgxyNY
ga2wJVefYIkNMSPjxyA9OiYrrSMRfmJPH/7uAFn43z4owyhgGC4bnFn1JtCz
WgyJUtJGUC8kvTFk37ioK03YHxquElFzpQRk8neWE4j2qSd2+icjDNHpVruj
tiH/L9RBkZ6rhP889oOJ9Xti6f4Z/kxs+x03fsPxzzho3IDcloel3mIVFCrU
VaBUFjQNJGgNP1t1YZFL8aA7LcvMN26W1Rpht4lFnriX/QL6SE0wWQW623Z+
dRhT1viSnXFq2I7WHi1riVnuw1OBcaI34xW3Wy1wBsuVKaDsDGBb/IR4SZAN
+GbgpyLxm8AW3ABrMgdtVm+HEGQjiVd1Tk+ZCft5SRm0jcidXKGiqeqcPOnx
dxnWjt8FZ3f7yh9BcLOHAnwkYpGGGXxICFAJbeXEf3bnCk8IFVqu/v92kjGx
TeIzOmfCZBYjzCZF0LukI6bF9Z56iRTuPpgCJIbdWNUXz4itzsSBFaQUaVvF
uEHQAEnwFc+fUYmid8+Re51qexiV1l36M4bWrhDpMbCRhTx5lwXIx/6c3LII
j5vBVCr5/8laRiHopsVZ1rZpyMqhO9FphKvZyE+E54Q3IBdCBJBNwkvGa7UC
plssamAh9Pk2o+92FHZxXK/m/Y9SEvCGPwjypWNM3RcEXCSTwleaXvGsMsRN
tgxARbGvE97IXWkhTe1M/H399/2JWintFzIXvYf4GZI/5jouM6fxuiLXTCt1
zfryRmds0TMGDEINmXiuj4lIQsRsLBL0bYMjLF2otZQtglUxCnMjMp/MI80Y
x/iuEks3SZ8CYGEguUARsHgVQmi/2s90SvsNUYdtaiwrZU3NyjckNz2B/16H
sHRV5GR7058REXG81BJIp1iUKASzbB8V/68kMtNcfhrxl/UuiWpWfmgNYXHX
/4LaJ4OcTZswBoEkfBpDWcQSEWRHQtFqU2UhewQxtOa07wWY3iE8wSysm19i
COcMOnaHbLFOYI7d8/zgpbrL7SVpqMT2EAX45YP1UX+IcNTTNy119xLdL2sJ
pdiI0Kmvyu7XQ9h9nMrQK6ohUp+ikdG7ST4A3Oqln6DPdKhDVGU7kp1gH92g
1VU3rj+11aMoH1U8OLp8XeuNylbTIkz2VmiLA+zygZmgp3XLiYi07JkN11+o
adkXk99fMi3THPwbed+81UZ+HSnRnN52PXqrfF6XIgvNlzSq4Z0HOYJt4wMp
RqSy58xozDUAqQJT6luAHJ8R7ryK89FUFAswJTowrxWuYjkJWTX6PIU0bPoC
Y8kyHiSPxIQHyReJJ7DZAfmS0CeBaD+sa8zw5Soq/6EG07gUXMgi5EwtRxak
M6dBf4f7o138NewVlDnEU7T/OW5FGPpNpP7+H5ulWLD891PIxtWxCxb5wmv8
FilK9vUJPwvi0Dyl20FulBaY90ZsDvEZKDA3mA1A836ioyXmsSzI9Y7J4MJv
H/HLh9yk+s4f+YCP6Ndhk5/QwfdzWRE4v/A4ymCiugU0CupVD4RLpjkbWDWJ
/VI+4xltdPvzNP/MRbDbTGYc1HnLJRIfAF43qB9RxXC+CDyGrEzxOqBikGsw
7fnhTUdmAdty7M41OhhboY3804dvPUinyPOE1euFs1M8QX6gLqccFPmmOGwq
rnV7WIfzrPDmlxBkljB8tWiMry1R0RMsoa8BR6QKMp3VfjESJGrOE2/1QbC8
ebp4ZEn3xGCLs5XB0uIYiSt8i/dc8+LeZqwhG2j5YutNC0klIEiW4z811K7w
OYG61mnM0tLW7KLjvpjsmgl5Ue5hUNXAKaKAGMoYw8tn3OVqd6tOc9ZvGuvz
PJyN/I8bCwZOpyENF0EnqjmDmFShI6IULWWJxJHzLoIHGDdl1VMfblRyaBdj
S7pXOzaLRbfXtFZQ9SAot7h+MPOcGQwwMsqHJd3Wt6vnJ43dDvUDvh8VFigB
5EohgkI9TZqu8wDcUfD+cXqLZa1gBgtR8FIlNAPuuG6eDa4CJeAtNecJfSv0
Kw4cvbOPoCCmAfzFLgH0jMEol2K8BBLoQfpcrYL2f2Gi3aFxzs/+yh6wB7j6
kfgCW0gHSNQrpJo1qyQT1ArErPyUOd3dPbTNZDIEAQbj5K65w8zY/6YWLqnm
26DNm3bEzcMH3sLUUt0sXar6FjcX2ndCWP4LWH9C+FTgD1W275dj7bVDLSei
ydTbVu+5feB8204h+4g9V++S9fyluNoew7P1VGJO24AVjSAbp0wSv+BdyNyq
sGCa9/iRRci1A77jTWJcf1mrW6fjCR4erVhuofwjmmra+hIZVXmvQEs28KuG
yieQiowo+TKTMBjl6BknMGlJfLYnKc8hGYGJYhDkdoOKuIG7/Jwjceh0nXag
lfwCDEwZEnoDYflVIkjhE8wSSxVZWzA2TLN3KdfNkPOnEYC1eAfWf4saiwnu
Zs28WO2KH76Spshr/xitQKh/b/v/V1/LpWCJQif2rN+XaNw4B/XPLmCQDicB
tXbYYF8gmy4Pi3wM3BIRvC76e633M3i2kKMKk00e9ysUWyaNRcrgWBxXUfE2
EP2jvMeg2bo6WhM6vldROlWEvJTwfz5QNZh0xc1OwTk04/oud8kAbUq/RHY0
zbnTWcZiX4epdvGi/UOe+DvLU7wJ5p9eLQxi2UwpgS2RqjeooQoYqZnS0ulG
OUn9opg1sWXtySSAAtqBkxbardUzBVyzUUFVQWhjrBa7Dsd/XTn3jqAct7Ek
r7Imr5BdAeMciBRG9W2RWpcJokeupOQ5l3JiqwqVwhuJCve7xjKM4HJWu8Kz
v93kXgcYYFB15TyXyps18eM/dzsJeaQ2i9kvR2d8ZG8lQU9XYEF08Uu1BL5J
arYv75ecwUaKctKReo3vFH3GPIsjfwdDUUy+faM2CmouQ/+Eibi/MLn3+xfW
4xMulzCvKc7+lYAz3v+hVvBRmoYeX80dl3kPP8a8hCXsAldPLnsQ58TWg7S+
VW0jH9ntnbaias0RjOPkCo3wBkJ/6QoQoKdaZIhzsvQWF1ifIR/fkqPLHQkp
tiszpldda7hXEbLjzzoWlMcK2pnq/3birFStR2pOQVbXXOas/hfE4CU48q+Y
IeF8ACiked/HjrZq3FgWUaDDQkV6HbcnmYlNwBlsmk0op7vHoxLUVIJCZb1H
qtlQoWhFfxhprfTwQxZUjK6OXmXbEicwlCWJU5eup0tfY29I5TdhYkA3ea/8
KiWunZWkqNzDx2P2kymQHiwa3x8BT0OE5dosU7qY8+ANvQrMzjJn6PEtYr44
ylW9HNqIsEYNVc7VnWJRb7UbC8/prRqbvwKsr2E6GhfEaZl53kEvnIyrZmm6
a+Nr53wvt7KxaXd+BFDKztMjtPKE77an6TYxvYpMW2FroPkjQzohvMhhHbaW
iq+zQ4FG6v+HutYpEYZSjMosFPoFVA7KhygQacuC+U9lSk3xHG9aP3kHCV0d
ag6aGMf34xu+GDLUNsKTqHIpzZibJPKyxAO1C3QIUcUlavgIOgKTB9gbD/b6
W0bh/ob6CUJ0qyxJLMLOy514BHrxuL+Oc4JSFUz3iklI7M6AH2/txZ0bAGUO
tu5GcUGHvtr1TSQuQLmRauwDNZiInjdDnx006ZGClpepdUI/AL6QR9IHv8Gw
SU7hI5kS/tu3rdTjCAR2v3rXtJwXdwRSAIUq8aGKazvt1UIdBPljTaTvoQT8
YmG7byW0IpbMBkg5OZznSC+5uic9NQSgRlxwQmo+T88yGWeTAHNdkwzxK0UV
n8GDfmtWqbvfiqud3fKrjAIYF5y0bRLf9kj7MwCb9gZFkOscWYQ5heeBBPAS
6AZ0VN7pMX1oJZvcUekGMXmm3q4kTsH7mU/vjm3fsfeueRI6hzRjODJtNP9s
0SxVhT2h5fNgvMquc9KohKi7XqVshdGJdDIqJMWTbP+LP1vp7ogv9Z1l3VOR
y0gXruZRERtduk+F0uwUOVl6IarA894oxycTuYMS/l/JxqidNJAIenmiUQ8J
H/gSvOe+2axSHrkrYYj9x3Dk94JoC8UUZzpN0UfJ3OJFtsg4el4h7YFVXG1R
NmdGdkanJxgIujOudZV9ZdBXK84SPg60GvXXFTGiWssgp5f/U/87D2mpQUVw
49+S7hegDoM8K+zZbkQUl3mSqi/gE3DnKhH3lVBu1VvBaqrDNr7xbMF2VqpU
rb9+eqAccD/lW76RXiOtoiifBxdwAwAwzEcoa2u4IqX7Eq0F3gYUzFCYNMGr
6LvnxJF3CQocepp+/IzMieOkcBOUvuAZH/mbYuc81l/5O1a0VodRL9OrtdrZ
04TBsd4VdyCU2yDAmk73yCf0tMK4nVArv2vPEJXFAibmCIMoHoEASjEK2qdQ
mXnkCjJczqxrvqyI6Qhur6GHUFlg30ExLZZxwlUXTriZd72DcAF4ivf0ouIh
Gx2n8YjF0HLh/T0LbfaLQ6vOKKAikUh189F7fLBHLU8M3FRhTs49Pfp81UKY
C/gSRQNO0fyZProHgylb7Fv1OqtwXYy8cj/38p1B4CPfzutz2V+PrdszYwcC
FIHy3Tw73lw7X8VDDmdL7oJIT0zUQCAtYQDIyhiGYluw+nvJxUDj9mGItY11
4o6pnL1DOIIozjN7ViyQ3c0+wqa7DgwmDsMj5UwdEwoQgluBL+aSOawUSCvm
Isgni9RsybxVOoVcRu9N6ou7q7JPxBfCkicmo5YXKKFa3vt6ha7HRx0ItX3t
WQXHzAK2QeUawdNWun62rPMM3yxhowp3rRIZCBzAEAlSWvdsgAUvzj4PCxwC
lqkMI/EgCeoecMupzk++KeRXgQAckEvoV0JirPcsWJHkNIV7nddqFcttxkHR
3Xh4/1xF8cmHgjB7ZcdPkSPGJ8iiTDx0f+eEJhbC9gjpXEYf8dFfgKnY7ZVs
V+VF3KaNl1dENLeEWYrETNgafENtqgg7jghs9BHqVcf5paLzRwSn2LZSxKG6
wIIJKA8h6xqtk3W9ND4d3ylAk7eKT6UITulrZGlurPs+OZt7Shx/4v03tV3N
iuTE1RFv5ASlA0DkbGz8+TtXNH5hMVSd3MrRjz71er+4YAt7m22c7X4P7O3c
jHe+0NfztP/YG5LR2F5mh9C3PjmIUvA0Y0CxkS14qjigChNqK45BGb2i8RDu
WpGhk4tbgWDM6ZFplcU85p2Td/YnBcVezTBYpENeQqGF6WcvSYMGnnFmAPgK
a1G9SZF1fXH+40s2ij65nKwv6XkBH44YZePYFOrkTacQlCA74Pw6DS+ch+AI
JVS66Uyu33+zyt/SxZL1McPgYavJv0BMJcoPRLRUO75YKc6LyWInL2zKBaY/
/B2kJ8QAyZAI9b9EyXEEF61m+CDCdwgZ5uQ/LKRojQxzRZZocnL508TVEm1g
6/ALai3T1hRCtxuScF8xr4DDUoerA9dwTgxeZi++5mOfedil+3/2T9qni608
VfgOjDh7NP/oVYJFgWYL4H7m57j4Up7FtFwD1GhXqTVH9YQfftXs9i3NwEV6
anD6yuQvqZUn1l/bHpW1NcByGrvqnSn6UXL0dXhU8ogA9I8JfbCXyWBMEm6O
YiGV+x7VadY0WFcboCKhfhY9Mg0IRTojKfuFxPm+bB0jRWXhQ5y5i2WKN18s
IXpknK13ALO0H7M7qobJcQp9Eccs+P4cOTyWzw4X8N7jUZV1CU+6wbjd/DSF
JqYfm/vpX4yZ00g8/WbsHq6Vozt0UisNQPHhmPPRvFxMblU5zY9ziQpUCzXa
FIVzXLgbJpq4AgLejtvXwpFqM9llMmGSctaxluB5B5XoOffx1mPA/Cl0WAUD
WqlvOj6cRQ01lTItv8nTYrxf615OQ6Y0eotL/BCLr4Fn2oASrW6fD9kTbGEP
mMOjuMMqR+tACidvq08XzVxgMXIc8o8xZhf7rqKN6Jf0M7eZyQWZ4B6tc1SR
ZxC0+vRgU7E50xl9gr37Ry7mxzKF1xNa0AtyAufEIHnJVZBR8BCp9RUJTYve
BmU67ZTxHcPDHkRwMeod4R6tov7ZQM2q2HFEbPSGlXNTEha5K/qOyxSdpN7o
10wDZOrUVGSKy2D5YVxzz4DVYJz3Ug5YSwPV7c5LjrsSNl6lOjhArmnTEaeb
pxhHaHDmaRUtYCUvScrZ030myiMdJpLkzYu+CFPqHDx7Cj2UbAlnq3PeG2Xo
pnEHeOLpBkDQ8WXDxqaJM32fLKn26u+79ZxBP/gZ/DnZAwbs8En9IqWOpSVT
ai+1SYdnd7xj+lco85ssXv+wtAXE5JSky4ZMg95lGOGmLM7WiOpxRhZyx67D
BpSsfbyuRWDjQpvF3Jj4/WLLWkPJJW2qSKMA2djyXzqTx4/jq223RpND/15G
OVK21zxi97HUQ5/O0vkBgpSoc/wSMv3gM0gKc6/6Ahb/9YYqcO8BXJcoqN+6
owjSQK/pVYSFY8g9j3k7arWCVHhE5ACELCrvswa9Pwsdt+GRkNjItYzKYq0y
typrqDgOWZJVVbBw8tO02RozzJHQUa3xqyTai5JPCA3ez0Bq6ikBhZLZ6lxd
oaF7tABbbVnlRUx9wJRfs7QCyclLGfZI0B47mxMU/QVwaef1W6XhoKkTP7mD
bHispdJeXr33l/bU9tSnEcGzaVuGot8T8u0MrXcrBm47ovOt/kJa7rwXtTix
N4CYfVp5XqodVOSni3QOw+AkiquA32EGwpKlSLE+BIPF7x4oYiKHCbC6vfQ6
ct/NkIugeJ1qHri/x7LXpZhtnio2QEudwbtIFGtwFghyq4Qb4FsIMYhncW/q
HajB4odDkDLV47jTV7SeGI1rfD5JekdErG4Yq4AoaVnUD2syP4nsxmeMrq+h
IxzKIKeHgczl1gX6LlkxXLdSC5R3ogcz93AeKKW7udXrkvypfV49MlOVliTE
luWtUSq2f+Jg+xGgkbQPw7TjEZfkJlQ8sOv1IYb/YQhfCJ2mSKBHAsV+ebv+
EXfU5b5QN8VOpIOWqJXVaw0oVb4gka+XPisIG9p6FI7Ip+3Xb6chNTjWe2Yo
r3+kGyaFsTcQpfgP2Mv3WBZ5tfjjhqkd+dyZSlyONiSM27P8T1aFM8Ehdhlt
JAHyzrqv4/+meM9dGyrWGxXN+cCfZjbg8ARSVPtgMySZ5ACM9Ppnem2xw2FX
g4bwPjWM3VPPTS6fUPLmJ/O6r1CsV4Y/1CuJKe09MzerRtW4PPMMM5diLYK0
4oeVR7j7kzMfmhOA29wCLwPAOoHg99+EVXaVZeKT4pNzPOfjyRbFiG58j0wC
lw32U2tlLwTSPVOOytt8VmlGvyOydd/KWW4+sxaUPLnt6spOH7wOR++H2p5y
zZ0iAYwnCa54oQDFZWBsdhngMj9ul5FzJOo6PTKLzvyBeoJ86MRRo7jNosmx
WKf5dbzmE320fHR35Pl8TPOhy9Y6ow5QzrNq2niJDL+AxrQuRRdpEgHLU+kE
lwxxpJJh08Ktx4h2NKY6A0O0Z40H7aJHygv9YjidgZqmvPATGGjYo5Sx6gPi
K+azwo02YQW45p7utBOwRMMTxreQ188uA4luX0cVipMygihzqWV0usanj2c0
KOGIPhQafNNmdrYq8A5mRJvqOvKeDCIJVsosAzi8AL+38SeGpKWB62p9GMfF
NfqfyqVhCjMXdS8pwGtKxkytjRxXIf2F+QfHAHehAMAVo36DwPJbJqj8gaA3
hg2AIzK53qJnAXZwTTQ1QRk0ZY5aPu6BS7P/FicgVw3GussSiZqPyq3g1+5R
8p5ZtYsE3ClZ635kObzIzxkKok37mOhJSRtjvJRZ04205qYkgUrowgw1Eymm
vZFeyztdWjryQzYwzTcp6ywRvao7+zsEshvFq0oVxjosjUn6nihpn6mcicbq
SJTPIzx5MdT1Q531Ws4tQ0vVBSrqce1Yxk1ITIGbYRA0fIzfcA7tCNM9evOr
m5sAxw/KcV3dbbLKLO5VysTC946nx86+O4cdmgnwAtjGKc6HYlVKfMxcRtOq
45oiFXGR9lVMIonFh2SupSTgFx4JwiVJ8qWwvx/g2cYxgDTI4s6I03wrBLPO
6iFphqZR6dP0/Ampl5BfeWDgnX1ESoHwr0fnT16fUZwouT5yw/94uD/oQY47
gZxYRH0beLjwGdJ6aleO/xKl34pORtdN0u+cEnkqJ1KNbJouYxOoyB8tw6+w
whVq1pKjAH2TTwZuWE3AXSo4XPrQEfary9uGUMzocmoFqR+BVnaYllSJNiVh
JJUPCqBysmaLsPv+Nsrz37McjcGdoDP1yzCIAJLYzvImiaP/V+qPFY44zvqn
LiuQwK6yFq3kqnqs6u8StlVcf0Kgr0U3KI43UlErZH9AWGQRevtiYbdzDB9d
tdrI7w1U4TTEjX6wCC/XlaMeQSsRqRJ5cODa2NvtjnBszv7vc3jMQIyp6a1l
tVN2b/3X6uViRUS6iiq1CuPLZdj+Yi9Uma4+aAS0FpygAdfV6ixZMtHDao+I
8lDmQ70sVJkouerpdVxojKvtauu+/HAXlycxj+gVAYtu1rC1gNcaolsYy6ax
Q48xBqnyx/DzQZVuEcEZD1PetFePjhtThDwXmQkx4qk/XlGyfT7yzmmwDLit
23xgYVurfeMKbQ7SaxtfhT9m4dt1ob/wUpyef1LJO/WYv2jEnlU2031ACvXg
krR1CkPn38AGdwlMdNBhUsViil2tttS82BRUgdlu0zoWjU3NTV73ueIQQhqA
f3+vR1nKO/P3qFf85R0XuMsRreMqKqIRTQBeuuHpcbdC2O2bXLor5UQmNvCx
hEs3A3TYxbwdOgDBqmOxsGGKL4/RfEwUno9mgOj6tnJpdcaq0dN6eX2KtXjy
Z8XKpML2k10TOMeb36k25Iuoh4Bk8vsQWxD3VHxLTgvTVBqR5M4gXjDgcqTl
Lk9WP94BI/f+R2wtCXNMu/LVIemuLrEXGUtQYPzaSq7l6h3AUfpt3dHdMJO5
nSVIEsuLJ7cSwC8oTjrfoSzkd7SaHNFFRFnUeIW1rgvOtyhynNTVWXdXWdFt
eYHldHyQBimc46Rt9Yg/sgIRE0rCch2cZC/L8e4HvFiOu7X4pu9WHe+wgXsF
tB1IGf5nrIuCFJg6Jlb6EvbvSwXRuXVbNkOq6sXQoGcpoUyOO6ixBpcHgnmB
73ZqL/lyIEK8mZgXL7PdBvKfzKHO4dClCjxld9RDtKPft7v+n0by1+O0IRip
dMlhNo8yTJw3oip4BAM+ys1nnNLQFu+jB/Ecgsgx9K333aN+kzS5Yx+wctag
rSENZzU3F6h7pskxlOFmSEoznFdeLvBrrnev2pm8R0SCTWBucySqEmPfxXRG
HdGC4Rm35I0p0JjTG637luWvbynj9yccP9sOUsIyo5eyjDsox673e2pRiD5v
hSqlkTJDPrlwyGWhGDoSIru3SXu/Ey6UXP7Z+G83WubHQgEnHcl7fWPCT6E5
chP2qfwP2hzkQnRBcOvHXfWd0GThC41uf1j3sAzUuCIe5gQHFJSCqlIqCJWh
bQSTjW+rFA6otGT4/pKCsDN8K2SQUdVeQzY0gzfeZk12NeTm+TQeTXWb2ykx
W94NQ6/F/vi8ks4i8dl8AVsh7MP61Dm7wVbWC470YSmMBk/07xJjGEU5dBlz
sjFcjWWobrtPpSAjGwUANmMPfumOSB22cehuXrJPfDGxgy8EMNPrIfCDQYWD
t2/6dacu5V/5iqG0mgiM0k4Ni9AWq7IKN8WArZDTywDL84xuqfVZcXpcMO7l
qdJdBYyKjgcARPW/irgt4NWWTN79RMPdhrBynxY91Ptq/aK4hInzdZwODDv+
TMlOh72mi0Yu3X/9ijp4x+1JS5BEGYhnFKwH48sf/A9juY02PZQoodhIRfgy
NlckOuc2T5S9E7l5l+O4acuzW5xdkr1Em9r3jx6Tjg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTr5OMr7OOn6p5oxcrBcHdh/FIQnx6W1VRP9lJyuVPzXBFH7YjzBRuzd8VpWeuF0ZzO8aT8GYhiua2U7m+gKqrhkqdwnt7oxkDLw2EbVLwvXwyqAqDvxbMRK/NG1dFYn+VUjiAvwn8L0Tb1anwyrrCCP3VTeEn3dYQPhM+hlHvrIMJjg4jhtFjOlh+RHPId6+AtohdE3KMNzLW/TRozh0bflBPMTysafaoqrxoHNApRELweBqOywehuDkKtryivM5Kh4kf7XMk18vbgkBuhwtaEaF7a3XObotO7h30W8RXWBJ8MHLdkWdG4p1QV6oia6pXhIYynl7SIuXJ8giLZUeqzlq3tA4vqUFf9obTHcZtJwmY/WgsnWqZc5w0aov/UFPpMB2Qt09zYxgeaGOvX7yhNUfrqZlhXgjaEDyjPoA9graJWd+Wym6EnHHHCvMF6VX5n60z7JQNk6KsER4bn0NvwD7wQwBjwMSWuToduKPce868a8bflZZXxZTNYHAt2Uy435UQLbW6kJVmj9qPxrsECXchOKKzsMoViO7WMmbaQNsKoCwQtOWVxK7pcmuAU2M/Q592Iyu4b57WbEaQUveABJCK202nqe3e1h6oPu2ABpdmEXJlVVMjx/DNAQIhQTjk6yWsVsDdgm6SuNwhhe3P/EnOX9slCwy+ouz/zkKmc86nmRi5fu1N3j4oI5nPb2ecVEHqBs869MuDf0BHpopFGcjWr8AFxhsSHd6EhW/ptWmdU0Tir1/nVHl5550UFdjgX0OEtyIqaOs3Y2znxUTbk"
`endif