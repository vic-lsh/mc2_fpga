// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k3rNekr0hsY4UMGz5F9f02jeD8+OyxX9n5z//ClYsr2FOgLkR5lOfX7fEJUj
ZrTpZb7D/qIzzbqYfaA1b2EkgJKduGykb0vBAAL99bJpBNqY4KldEbKDuuW6
u0uhCUWoO3APrt2EfG07OafT+2GZ7DR9F4tuiO8gqeek5PhNCAe5vwIWULg8
/EP2uMYj2s8sOzM+tK7PBjWpD8Z5TcSZGf1CIjNuJuvWt/w2Rn7fKcv5kttX
+b+BiV+cO/Ffi82b0Rpz3RS6lXEsRjXTjiznKygZ5XJEFy+a3MFTdtiPIpO5
49FD86mw77MI6n0SmRLQiyCcNc8PTIaMEVWGya9++w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fDxGBDF1iPjpyd0kh7cv7sLydatibLf03tUjsmjqp/aZaXRlmq6x3pcy9dNq
PQIs3whh0LImevedWO6Y6BAjLtHXbFZ903lHdF2dpu/o+2/w1su9BkxLz6w+
XXK+nIoWVqZBFdtwIhu7j7cK3vdjY03iEvujnF6FfLzO5kOFdPlR0xBdBu+r
qauF3jeEWr3nHUf41hGbBrMN6yYOoqB71CGj7K35GS//vf6SwTSRKWqY1Fec
jwiBWH7F48hyo7If68AW5JdAMvOxXr9iyZmlDBZnd4AFo3tNgQpQsvPl5/ax
K02M4NzHDyiQjLj81YwQA/v7XgkAxh6nlwnXV7jhAg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D0tT3hDqb61edx79szgdmZdyevUfYDRS92tROXqAR2dST2FLEB8fgbgvIwXx
om2clTdmpbkVypZ6o2tqnyVxo/SlvfREAXzwwTk03nOQcaaQoIpsZhcnN5Zi
HIlsGa3WGKNrqYV4HkrKVVyoDhc+yq+1H/aeaTGXR/QU00UPVVgQkFxt//uY
2Wnzfb8RoNAlhWQyXPXkFoz+TmafZwxTW6p+Va6p4WSCYXQwW0YzucVNeauU
K+TB5Lep2OyoJqaUxSyzBbH25302ePn7btLGh7MJ3ZWPim4ZVOUsK6USDgRI
VRYgdz1gDq7acCdkx+KQXhi2/c8XfkWerk1okvhBTA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
StibywwI2LEoBTVjgMSzrH3XXzfTVZP4DCP+jmoYzVh+rNLdPAR+kTYRHUrp
hz4S9IE1R1FfJNKMOO+2RpckWBuXkvTMH+ha2lyQOOIqy+8b3DD0dAXKI8QN
onsCIQ4mKS/uQmJDHxCL/ebD015V8iy25BHgHb7ulnaogCYGRTfF76lWx3Ig
jXPz74NdWpiBtmuNJwcyVs7sw1L8bamavT6ba/O3lfTpr/ds0ux3UOe4BonK
lfuwoWroTwxyftMcFxbbYknSMVe8T7GKFTXnh6GwtS0+NQNZpJuIDRcq7264
sdgx0hkssc10o4xyDfUmP5gwhaAU9fQyT7i340J2+Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z81SHyN0tsZKUfRTkPjSdILJW+Iz5Asf88uzSziLvsoZSXm5Bg+cF9fLN8Ne
XpeuaP9f+bRPzyKDF4R8+iHh27Lidqty2pwk/UofyS5ZxF3yNLEv9SGcG0C/
eKtCn4TuiAsPUEsejtlmXzqEKDu93Bo9YkVao1rN18ddmd32vOw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uyN8obdlBwa6lEyBG8z2cjMFuSsFJWe4fasiS80yu1H1AvorAY/9EYzfithU
HmhGXgfneo6rKQg7ClKVMGTr9YXnqbp3R/jHetuMvUK1t1JiArQWL3zaegLu
6IoJ1/mvD6nJUrIVAPXeG5NtvijzZYmFJMXIHsLouthFOT/CujV3lLs+WFBm
mJ21z+0m2GXYtpeU31UucwDtkGT1MgHLAPtWL4B++M8BSEp+bBkxxiHmpVt+
+DHIcxk5ti/PhMEEy+CiydgE8ctZzPQkH+wcdjdmK5VHWtbq+6jxiIuD66aV
WELMUZYzYGZe39cGgtiK0zTjEpHRpgmUeLTy4Y3vKvIYv73/lzaoSyUdgEY3
8ngb0aPlYZBaWfpwAYu7VBx1No5yfCRPLIlXNe+H2pHf+POQ17lKyQhPz47h
K7P6xTOtXTJOqrHfuXfmgnuNq5xPABecO785t5/qRO2iWWQ+xn92iKBuEDSN
D95JYB5iadaUX+tHjdjbMWb/xGSfrYHH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XVSGITEz2aKwfvpAMqRpLI89WIprP/OiTZNySuadsOOp9OmPXz6GBkg5xHen
F4So2FA8ai5OjsTAa0PqNxqnEIJj1HL9q6/uGqEqqinC+GeKwt/yvfAJy8Rt
xzGH34tgHw3gq1V7AeERxF6doHLsfiIknE4GYv4erJlL66s9slE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lf3vVksUU+EbZbQQrGd9nuNEWjQJbxyR4SR/21bBCoocndD8b/R1+RJY+8MD
q1TxENRlFV98/2F4qKuGUjn4RFUZHgFISxjsFTwvpWY71qaZFxUjZR+iaON0
eX9NFlxrWfNBKx2eWn71C/IRf3V5Bq+THFMRNqfaFxbHw14OITQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
avRhDZWILoWXmF9//RoC/rmSRnzhb3rcCP23JSBOrp5Sxm5MdY7VRbNv/NM3
dLw7FxME/jTAwZTOjPmMO/w+FTFzkwAGha0ReoikI3GJYEK6OSG0WDd7Bnia
qTlvIscinsoYAkgOFt2fq4tRDBQIAeWgLTAWbgK9Irbcet227INXzzO/dmu3
33GmB/9dK5SVQ6fRWuxrcBRENupdPS7SzhP0FuQjWpSdzn61s9xYUnxN6oxn
BzKa8N7h1qorQgrDrLpqz+PwFtxWMuEchZUNuFj3IcMFecMveCHLrJ1YLSCW
ndwzi2MMD8y2n7QYc1K8JRHzyHR+GRImAUtnDXp9SfmOIzSlaK2+i1Gsg/eg
s0d67d5dkMLJUl0wDKdbhMgMC4Gn8MESDlTe1TgS3qxcFqMwn4JuNGh64eIr
M8R3N2d7ho7pOzOAGTyCbtKyywD0WyBJAAvya5z14FO6ekSfhyk1fAWNsdyD
cc0bUq1i64/LO1ZjZK/Ws+VR8/8LvxLv9cDDD6bVdoKBXYNVSekFMnEfq6H/
9gfoaiba8clltUS7APmojrnItT7Fv10fd8sZx6sU6H9JoWVbcco+IepXQPbk
25qknK2jkKinv1dO+OpNQbueS9t6ylpeVqKhmfipHzyMdr/lMDJhzxBRuTLA
g0O1ArZGu9chTR7lBKg282JA8EH0YhSqt5pLmabkVtOp9XIrBCFJ0vVk2c1n
vLAZYI+FQKOEhHT4Uh8Ndi5fULej14SrHbOUnhShjjNx1UHd21WH8Ci+cw67
/MM+fQU4cdJz0JsCidBJuv6BMELC3L4ZbEmusWgxNA/FZU769fF/wdLdznPi
JIzkFOCQsg+Vj0nSI22GBtSo0oJZTgn6RjiKaTl1fpyI7bskqmp3IOOvwxBS
2kZtjxaVlSF/OIS+LS3t4AtMLQwju7xEhRDsNoek/gD4ciMO1ay+dYes0mAn
cpo9FJEhbYXwVDbsf4Psau3szSLfyp/TBbx/XAPKtjIKBumxJsg1R0C4sjiK
nq2CqZxC5SdUnqiyMkp3nvCINRnjev14uyUHur7h2elirv031IGybD0GzPyI
kxRU0aWo60XVEy7odJpQx21M4cIjk6E96N1aZ7GELe24h/E73/H2V9/3Ajaf
ju6chpcBYKCexA78DLdTievbp6XPt57WuhCukiK/JNyLWs9hut7odNbbGvMQ
CvLJi4ffm7be5lSe83wjm3LbM22HoEKGi+X8W9EAV1iTPj97MaMOrs2/YOGV
npFCfJJmJ4LHpk+Xst3dg8tFmo6lFeibnoUZXdmujsuID/W8zG7bitVunmxn
jLrTraJ1GQHpD5uyIjPBLtWCPhzizeRpxK93zjCOf7D079Y8wkdzrgXzIkI2
/F9v3LiUd9CVyFpPiTs+iUCzTg+sXq3LOBYMRuqAtlm6KYxZWUU4JlQbgHHJ
lji/L9bNCAmivDOaDQCj2yAeNDipdUQXLNQuYTEJtkpn8ZsL29WzpAGBNVYL
OCPFURm/d1T65slXa0jb2VN21OfANfrG1TPcH+/wWJNccXeojDZMmWeoe0l2
4NEkXI/fv8ZEiCLBTC/x5LAGaNrYDTtPU4/Bk/nL3u6wthgI3Ox2dHmDou+h
5bpyHrMk4N6e+VObb2AtHpwGXWSYkGJaEP/yqqKyH0BUWKPAjNaKD0RoU8y2
Y9OqwKa8Z9AAchbbndplbYj8WuWomCTsiE/9MB5zoW1pIXRD8/OmG8mD1TyY
3Yom5pkv83vXSAy2ESro3TNEa88H519dtUJC6zjkmE7uTCG8OsSpCDv/GtYw
yynkUOM+Mj4lD8A2ZlHw6ceuM2tCoq4U0LY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdzh1OuETy5nJGMdZz7y0OUQYvtkFkPrW0ywVAxF8hHFxUisWyxS+pAeQQdnooNillkcqVi9BJCRDhQzW9aHWQkw1cccNCRJsuLAX1/seAQdiVGSIU/tDXZrC7jJcwclew6Gfydz5eZ5rOzBPlvnxCctO+Uz8Ik5lYQ795Qj3Ar0XuGFum7rBnE4y21DdWHbcDQRCDLOqP7RnQOxmJsMRg21sFdAd45c0OKkwsay3xqn4n3WmQIUzPJXwbvtUb0D0I8zpbXCs6V5ztbwLRRJpxspMqgizB8/c/6FZAMIwgKkYnwICd2pubQNIOXpIk1Fp74HF+J2VOJgoA6rvNf05qSdHLWlOCQC48Bz94jcA3TSAO6Ffxvq2/breGZk7Mz0XrlRz6oTirmn9YVrxc7fOS14lftrZ/4migupxTZO4FemySNHeVrUBPqkd/qzN+6lgvVIqh2VouFGxMl0lU6QX/Bu23hcb0fOX0SjQAoxKkkvvFoVRIn4Q9ARXzvV3gwaZZqfygsm+U9W6Zy0Ohz1jsJnHMqFoI+Gihfdv6bIskhZ3U5AlyeaUIUPS+LYnqlxniG9XJRE4EPfs8nbb4lrE4ii0NKMyHasgOr2u9XQbslDwY3k+ERnc5U+WQZeG6sEPTjtNNZyTvf6LR4WlBKBRs59vh5rR3njCCT1wX/BrUy2syCW6tViEE9utkD3X/Pa7JZKhBUpAqi/jTfg0yqeeG9pNx9ZYmjzPm9Vq7nfvCqZuFK7sihVmKC8rSvm4CD20owO8NKC+FR2Zg6d+HqzsBu"
`endif