// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HBSzr4XB+/y4vVxWoRw68dzEUOBUANI2aOlRPhYxO8El36VOZvIByaZbZ13P
rPbLy4U4UvADvJHJ/fhlxp6BSpjaz3oSQNxqzDVLqJVARnMXB/yYYUKpregN
zZ8O0L4H8eKNKCSdys8SB5ZkJ3RlDaAVE1BZ+AYGkQaaQJ2F8DqxLte/DbPF
/maJijCB2aY6uCOSGb8C9fvhBtCwJKctLWHYXsYv0zZdS0rUNAOMCpjnPkqL
Pp46T2qUkCvpLSeV6KsZZav4QiGNvi85KSv0MlWIaQjKgdNbOfRDvf9WqZDQ
il5sUI6uz7Gp3wBeM7aDKpaskffXdTxPMaSAsrOubA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qzbmvCMDaGZEsgJwk62rAFe2d8tL8qsGpDUkDKFJgpwUori6VNQPcHcE/rrU
3pVj0yo9KP+N7810il7NXDqM0q9nz1HKsz85fzVrK4PLHh6vUFuk1XSo9RBy
kpQ/z2NFLbDJsNe9DilUo4l+siLqqnUSH4h3h2lDRmfgYo9UgaNGROfVwwFb
tqCH0mRC+aORs4yxyNbMA68+JiJIh0iIMMv4yI16Yi2r+n9bL5R+eMfRst8a
75f84ELiJ+yTohlijuQbkOqFP4ILcFliR7vHwBQEupMiS8Ab691r1kJJDglL
TZpBaiWctYezxM2tPxzHfuGej0MPFF2XTOqd2/MUCw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XSXLM7CVvLSxe0sBTXir8AZH7ZWQeicmpscltWLrt1RG/YohZx1fW2brwDW6
6iy1QrFJbr0jXhc6HxYhtOi6QddJV15uszZb7O4008UK5mamBGR6B2FMT/ah
gK5ufVBETu5HuoeV5b684sLDYZpktVsKQmmIKx4uFtZI0Vb2jY4+WiNxxxI9
juyKooK/3KH9CxEbYpvU169rWDUu0vPPdmFBKVvJgqltMUJNXzsfbsKb1LAT
cLRwe3t/6ew5+h9d/UzadniDBAcEjSIfa2221J1CgPG6IhTr4CCUDu18x96F
Sn0j+OWxZS1YfQKpcgoyY7RTPO/weV0EMvMrvbwT+w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Z3QUo04PjKNLTBC6ToHkmwJclalbuRoijW9/xuHbDRFHjXYAbrUUyQ6pdQAq
7s5ovGAna8Np+DzLhG7Y4HKSAkvzT9NZsuhdqnHUPgt+1byvFjOOsOMSYU5K
dBEPfza1xJxfildj51jwAy1WyokS6TSuopySryhk2A+M0n4rc67k0Alfgm4Z
NlyfDbnaPt147vxoNcJsyUS/NxBhXxVZg/NdIfVkMhvgq43T2RH92FzEl3vq
65QZmX3FI4rSpio5Yt3IdfUPxSFx4GAgLON4PkwdUIGpcMt3ILea+N6+Rw+7
Yvqxyjoxy19entl1gMnxgyliOSUS7PWbeZp7Wo1wag==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UCGHJqrJyeqSIOBLqlROfQbXnJ0k6iEF365rShgWKwUMkyo6BT/676XcUCQc
LTXOl2ultZ4aGzBPcHBb8FJTcRC0SCyCzYNj9GdaAOSMHwZrh6Mp+W/budyS
OBLDVjiMSLSmLlcDMYnNK3cK01OZ7Uu5zIroPMMTwP0wBcSM9cM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
K/iPu1l5vvMj/TsdhaLVcO7xxQtddSGPMUqyV7HXfKLG7zVtmdR3NNfkUXlO
gxIawlu6GzYmD1Aj0CxuYUtshbI8SW225QHHs0jXf0vl6bczIVBdnLNhmEMH
ryWq1CcdU9YQUKGOVMJWDB7Daj06bzBVxysOFxMLlFUGW8kh+bHONIkUxrCv
enYSLceTm4dIupecpUywZs6DIj6dIhfrysJmpl+8LiSsErZpaHE9xGXjQxPW
CNUS4+63QyIBWwccYr7gnkMdlo6DS0wumQSlSxRTOKDvnZDLFzl2uIJEMyhn
eZaVBurRRS5PaXt++v9xjF0cheaSh27Vi4ET6826Xe5PIhZqWUPWu+szJC4V
rrByX8/1UnbSD/OpWnpTU1KA9mv6R73u8sW5fhjnV5Vy7O+9jyfuRcMRPl1p
RJkPi0b3JKXozn45Y79ktw8Y0moNOykdxeiT9aatfhzBHMEwygT8E8n28l1S
TWvuDD/HUlOCSbFA7s6j7+CvRNVMXVZt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f/1wU8NzHJP8rt6wtfTJxkn5no/BdUExR2zEV99nWOPlizjaShp6xti+j2nc
ulUNqY2cOW3YucEjCfm/V9dtweRRoYgSkUFMmAffiC6JdqfR1vl6GllgFS3y
bE2y6Gs1LFPLPt/TiafSfCvUGTzNq+vKKYMHXMkMXGTZBDBwvvU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oXrRO6O33lMEOJzdFxLhpIfz4jzAlbu4PEB0sjsKPj9e2j5igWwTeXLhMHf1
cJTn09Ck2JyQUnRXrFdOylEvmyZksnxEQN69hEtFrJg2bwXcM6L8Sk2j7+BT
jfOUEAzehZ6sVzFBFxagLvp+TMhSqoSkU4j/pRt8eGDZjfvpScw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11008)
`pragma protect data_block
8ldBa3KN5fi9iPgQWf4rUopDZdv0H5DSO1d9X30aBcE+7JYNxkwvvW1WHXaD
CfnL5FFBytP0tZCjM6BEgM6Aer547hIOV1czru0twbELef9tByqxsfuy4wJz
lVTmWuv9McIDteikzCyiVL6vqClfmf1mm9dYlMT3+Aki1NWKIBinaJ9AHefP
fZZkxIfXwLuxwjPggBLNTLcefvmao8DD/rHU1M+V1nzefeJwdPsdwxndKo+W
4/L+mPJxiDpnvqV0Uy85bYSjFAqypqfNRKUynkNP2LVGcc7DpWf4TlQyb0QN
CZrfyk5JUd6pvmTvqiIp0KzN/bqYEq4CoYkM6X31a/JamHa37gnLx/AJF8ru
zgNv3Y1P2i0ZMEf9vF3DgtncCdBzkOkYGPUFWhXRNKyiU66vbWB66mTxci1k
bTn0D3GU0iG6WLVWqvYHVVKt5gvJBg87VBQtU0h+aI2TCaKRok8098ezhC3H
uBOixuUuuEPDc9tWlDRMtdbZsdC5RMC3R/FuKSPw007nLr2erjzgT7E1zjf6
8i90+8sptbl2eOGi3YLIw84LzeX7BW7xN27K4F1QcprmTEDXaZRdZMqaU+zb
3TTzCh396C+HSyxgGOSIMX4Purma8DQZNYN2FVEO2NeSUMsFugWyoGsMmHaO
scs5PHSKr/jGMgQwb8ovCJGhgzEpqqerrPwl8VgY2gD0hRBclY+Fx38N76AL
dcT5mlq3KENwbl92nP6BSa1oLq6IdM7jBraKnJIJtNG8y7k9XueFU4p32hh+
RHCzg81e7lwNMYZLgQMUCZP1TGNtuw7qHSnnNCaZXRFopa/HT9FwmReXXElx
JaZrR1lcUbmzgVEIAft+yPjAFK84wF3Y81EHo5rSp2SAXwXLrC32qR+XkPlH
E+KsPAhncmqNLcOLNoabHozGhz6ptwjq3OvsyHfzXyguf1Vflmo7Xr1sT7sM
6UbK7Nf3LsCb2exKijNWsPIKrXTugXUUfOzPZaCKUQjOSK26nxAjABkCmk1a
M1AbKMWkeF+1WmI/6vQQgnhpwpvGdU8aP3EU4FQBRTfNncs3ZwFxOOqaw4r3
EibLtxbygrcK5yz4jPXEq/CS9D1YaSprUz1Qxz/rT+sDhWC/iUoUZ0hdcmy3
i9R9/QWL5H5ZMMA8sL0iyEXIcJpXD2T+uGYrZG4Tlrqk/8yWxCsxmTQraNgv
e5qloHMgCpwNoheeCnoOu5ylfa6cZUfVhqIezlymoF8YEfvPGsOEfi81/dls
SDncFzZx2nukYTnSeF4fSoSYBGFm3zG0UsPlY7951MB0MjDWcK3aOkQBonCA
kkTySRS+so6rpgOrkyBHCkgqbFO3+AZdW1OJ0vU0FJcy7lKrTwTTg34J15zb
9cbHZSbEUreW1nhfMUtoFv7MNuHsqHdvTqk6Z1yHnVbx8b1b8waNV6DaXRDX
4M4JYMFRuJ67zNqOBgXKlLLUIaTB8ZbxKrBLNX/4NJvfEKpACHgbzvua3zSi
zgTkjdPQ2sOXuYkyW4U6axOpt5QWpjNPHftSVBcP4glTbvFePsm+yuIeJlVU
rCkuhYYvz2wWQfjE7Mf4vBbvKc2FcwGkrHARD4dsbcI97+eIgfz2Wpppl4zo
bb9hlgPsqDZy4LODku+3LKA9mWs63HXkzk3J6wnc/EhJ1xCAeo5PrbGQFjTS
H5y5wTO9xSI5g0zBZA4TbDApNnhsqKz3bG1dyPWDnwfih6meocp4kaHjRLg1
S1k3lGw9TO2eolSqle+VTLR+QhtkJabks29zCHDvWsvBDVtVJ+wengvC7qIe
+yjNYvlHqPXKMBAvmFILDNX5JDMrJEB2fM1YgkRjmgl/BOYlFGKdrbbx/Wp7
jTCFhLk0ttBar26NegefDGjUiMtGAwoL54OWAWAAgxK8znijIdTxAsRNcA8a
26WG0iMQJy2RmzEGsH/QMxkEfa+2VSEii+04QsfV6MDyz6TgCQUlo0bOVE29
MuMzXr38mebHNxKqbKYn/F1jLjHOQHIKQrdVvhXbTPGd5YVTrj7JX88HLJ0g
FZogkY1+IUTexe00sKo+cI416HXoSI6WLe23DUhDjrbjtQNhF7gsLPvcXDOR
w60w4JJynHlyG4CZK8cM0asFoHmgkMgqyb7Btb+qyt/aSA92ql03Q+2lVdhB
nhtCYlU79g01OH8n84YDugKgFohZSBj8R/O9ar/oFYv939XntFAuFlyqJ55Z
Uhab8Nhgl1cYtNx7XSrxW0P54JvPt2v4MAjWWpw35c01+nL/Ls3hNrTtzDNf
mXwSsMHkY5zk609dZG64B9XMP8O4a0vVAiC42INqPjV49Mi56gAUbR4+EPMr
rUcMiu7TQpf3OUphWi9wob+dkR5Vv7iEX9+wNGw1a6VGcQNrCjTS6culgwLe
qSLJV7oSKsUvsblBw+21uGXd5n17l1+ydg0xLONOlcnU97y5v51dtfnoA18A
FomwcXyy23bYTdrtIx2FuiVhFLL200DiB/FdFU8eO1PzZi7Az8nvIAA/TtBy
Jk6bcXE2Ch5oganrSZabKKd+gJBvlsY9w8XW6hdD9k3gYubFuO4XZd5sgob2
8JiFhlxHY9vnjTaSIz3q46V7/Oem/vjxUiLsV9L1eE/yqaoZR58vvMRHUbnk
O/8EUOqNLP5QV0S0OLBtV2HUS7meEZm2n89wCHo5kkWffjNrtGGBUtJjoFK4
5KEAm7aDUzRN/v7v0sHYyV+2TR5sMuPTchpy1+BLVr8sVBCTwGPxtgdLL0f8
IOEtIKya+cbGVqq0zte/EVBHcfD55itjb4DqrJyl3c0tIm+JRvkwdrl7ia22
E5oStTVbXpjH0IshWWGcAqYhw1yD2g5fPtD7W7QwAqkEy7UPtFaWmuYMPzTk
pZtS8iOuS5m5KGxhKRuIhbafzjCgkdvYVvHM5c/2wL0QzaaAZo86otRvRhey
+u/qQ7c409ukufwb2HPr/wpuLioknkCKbXacf1d+8vhA/qFjxBhPJ/Au5ivw
B5aZ8G1rnElEZ7kCbiELB1eKEDRkaGo99n85BgalOW99K/Fi9VbJ6LxkIh40
qU0I9KZlqdLBnNfYN/2uJJonHsHisx9jkPS9Is7QAp371uwW5ePjvvwfpO1g
LnNfqZYDt/2TsUKvJYz7SOitzXK5rZ9Wo7v+Qw8qip6oNKFURp8Oc4j5rolE
LzYj9M0HgBibrHY3erpmVyVkafhI/Jq+xg4ZSxz9WGGkeEmeBa704IGJNQk9
NEzN5QVm80p624r87eFjbvCEt8PUK6V1xp63D3IYXoB/QfTk1RsxQjNMU6FC
YiGaC0IiLCsbgqnjmmTsCZpdgvwpTmBq1xwX5YxDyXbdPsq8bWnpaS+s8fmn
VPFekw3D+E/X/gG0zOPJB4evb/NYnayRqgzW+REx9O3N7mYWXR5sjkzTAyoi
govUmzpX9MYaQ89OBU+6SiDELymi46LsBrQdYBxwIg6jSJIqygsxVME36EdG
QXn1a8xl20U8ftlS1n4VIDZfo4vYn01l6zaGCwzvyPS1qMBZrbkseX09TW/i
9+FIow0kL2TrwBJ1G5wq0urza4t8xqpK/KKyFM5s+ESRL+Fxgkk7nXIyrUC6
wVmIM21aImfG9IFS1MVVO77+fcvJTdyVDuo8tiVI502aSVBmzwXPpgdZessO
CVIzXjHPwtlAExYvFZFgXFx+EULjmAq9h3ZzpKWG6HL/qbkg8Vl6Fb0iunZv
zpjIfFy6/2AVPVODIvym6b4KnY2dcGYUFPxtvvutoMTQl4OqTh4SFIT1x7qy
j7xnuYY1Q/7EQ6SeoeZCbqjsTVMJN/GFSWDYaS+xm4lFAIdVF9YUBxAWS65d
l2zM3g693BUhdyGWw6u/2y4027hqbkCj80WEKOYoHSzjdOiCsUHLN36NvJFh
ZAg5/HGMXABYLy0CAzeyprUXTs+LLYWvDQhuIsAPKQDMAoFyYRz422QQRXOj
o7uTWHjeJfYfYmU+I8l+qQONSfRgapcE+eHbh8P9L0n9gyDAwCSDWiwV6ZDX
g62pdQA4ixR4k7jedlBZ+Br4DpLyw9CnHXnDCbvPsIV5KTf6exKG1xigQoyO
3QDWZksy2VoNjAomlSKVC172CG9qWosNEBHijvCnmZLspbdOPs84lAkVVZEk
4FgZJJltvHwz2ESkQjO4N0TQcRHhI0H8DRqDzmNoq9DfMuuKzBWPRtz7QS0c
nX3AShX/9ZhJGghQCSmxDE/G3m/tlsP8gp4DsP9zTnM2DN4tsZ6yrbn/Ms04
4vUecINltOHzw6OH6HxN264lPwiPjPwQB8UjauQ6wtRJAaLqFo81dI95wsiB
zwccERZ7vtHCdk6hUuc1QbuZXNlShZb7jRZ94+EzdmkQxxC3sqG7FF5tWUI/
hK6XXmqzDLyukl1VT9C2iPs1dh02zf7ewLknnJSRtDq45s1KrLZPr25jtw+5
7F5QjLvmYuC3yY+qptqyYVSt5qGsX0KPFVx9CyVc74NtZrqj4Rk5M1F/V+Cx
jU3Gf02PI593eRZqUImtovCMjqjWs7qNTYSHaPIIDAvRB9cxaaNt0IkVY9bU
s6YTaChSD1tb/TrBFAqxtCM860cYpJuJ02nArsEugHSBOe7bZBgnBSrO9m5p
kuXqP49poT9QgR+cxymxpTMWMNuEf9KBL7KvOXGVL+L59PS+jEhdxjNTUNpY
q64PWDTchyEQdywPhH5GYFRKh0CxleIfCXKiNWFPnLaZvRrE2o+IkQOHCf0e
0eRa+Xf1SFTO1BEKFV4c+LPstAuMTGsdBqXWPVtxrJC8rIXaEGrbnnwS9uOk
E9ibdaWFtHuZOP/91/8bIQaKhMAFpsHsdjQD4rDaynSx4Wp9dnVZfM7OnPG0
iB/ZE1gOnGmjYebi5yH9FXPPU2vcHbzNwDQGIPBmmNSR7JTSm30IrY0iyOI3
42arHT/yXBPRRvqCAK7j7Qxsj11xVNSJBqL8J4FWMI8gU0jqQ4bgbfcCKZNR
9nWrIkoqIaMxF2QXyQJXJeKxDrQI1AV4ayA6hCZS2CEG5Y1YaUcCnrC/pv14
qgJKC4lRN+1yXpagqejojI0GcsUctmF6QOzkZPdgI7+9jVx739dmUq0Xst7q
aNcklitja8u6fryIEgZB2wjsc1Ds7ILeIej1VUODM5VUz/YAou6tjPfBJ+vU
0G/7sbEDigWo6yvt/HO3cIMg2ETrhW6I8RmZ/f/CzCcMhnkKktrbUemSUgl3
zT487m9suwAklb42SeNR/d3fjb5UcJoEup6JlRjRsovVZrwlNl3kY7pjhHFS
8clmVUla7KTh1xD/o6ZMANu+ZqugdPgg5Uw7hvsC4ZmylThj28d1h46iwvxq
OUiBdaQyTB6qwfI1KCb9R/Chv9blLd80InAtdlFcTleqjSp1S9ou++O22PkX
gnl3ksqNEhrMN2xYVv+v2csBzoiMClYqpdopeCeZv0h4I5iVD9Z7QUCZkZsL
VMRY1hhSgLK2PniHufoUKimkBl+8B4vDdqN8lkMGwdZs6BznodCZHg6Ux5Dr
r5NBjRjCk3Nj+YKJNF8wKGtGfQChjoJ7Jg1TU7adNyS1iQJI4xRls2d5dgXn
WO9biu+tiJiJKP6pDG0hs55SYrdr3dBWOvzPX8sMFDqUtv+caCdOFXnW0hFc
DdUB+eW0bK6xokHBjrDulNKzCV2XeC7+me6gJS6vvm5IKeQEas1q5YInqtSU
NIJvKd7B9CA0ZjpUXy80ENYhMZCK5sXLu/AqacOdT19wwMWkXk3s1Bvr9xuj
3Ahg/5WeWy0zCdXuoXUa26pRdWP8iF1ZybT4NMh4Ib/lUNBebX3cVV+C4XRl
Clr5OCpTSvZJDZbZoN/Iq2fM2smowwaYj2w94p9dNo2pO3YB+bBS6QFxFWOT
QGreuVztZQZtO4TXf+clSzmxIWF9g0Gsfi5S3jz1oUsQHiVDc8sKSFLWkSKr
JEDFXxnzonuOmkjoepxtcaR8AG0Ibfp1D9HYVazYZQMzr4VZt5Hn9nfUh5pX
yyFuzaMj9oK9XnVaauCHqUvfot4XiEednlnHae1aVP6zvyOw67Mp8ZZJK09t
E6HHnHlY7l+tK5pes+dpdymNXA+VlSdf3I7TUoS9/DREVxS9O/vhJuXIiVLn
nAg5KDUw4sUfksmhJ1z4A82VdDO9TNAu/UaeENAJUyiNhuiw+kFGO8wljj06
9Rc8SyWItZjsuOjlfi8qg924sxAm+PnMDWCFZiK1yvKrNFaw40QOXQyQFdp9
Mr9Af+IhqnrcsSCWolalvi23dxbY/ec5RTV439AKb6f2D0qKAz5D9q6shKxV
o5Yk6/cV4iZe+qyXwJpHnT5DxgWUD0E6QKr8h7MhPy04DTFKH/8wKnhRhYkn
YdvlbLFjsKUw8ozwV1DGB7/6rThKgXX3FqIkqKso27zirk6vJQom9J0YUBC/
VgEyzSH951WOJmeNj/WmPWwrER5/sLitg7rFsxCi13AKq0PW+ici8HbKFwi0
0si+8vkqrs4+PBrZlFZOLZJQ4d4W1rqqPHZSv+jHeDQgrlFaeqKB12W71Pnh
GZ+PG6hDy94FaMGrV/mi0VEysZyYQR6ubxu+EEhKKrjWfWfZB3mPT9FqKnf/
Ig2Z3x/CNxgvwaXBXHyoTWRCvK/zhcJBPevXkjU04LKSPM+dYH0pstH8dkFK
mWk7yz1TgoomERMQ2Vbyngm5C0KO09PODXe72rTj8m6P/I3bVquBQ5btHQcM
migGAU1DLdskgG7uOeOXYTv+G9iOKC874gnIQRhTnt4A/U6Fu6dpbpZibvw2
wCNGtVyGT/c6PYTGCFeEe7gGsED7oo6O0p3q3zh8IXHaiTvnPDyFqcaJgjvT
rLfZctIEbwrHs3KbUx03fD9B8tJE9BR7npzZnt1VLFEZ3gpM22PJsHgq7vcx
RVeqkvVJL5JWbqDqsFvBHBrXYc0GMMlqAPnPfq00xwNNPdTMFoezYqSXnBbz
BWJW+hWyNiyJ9cQ5/VRhl484w0SpOqeYX4F71VVxZ3pZF/mD565PIRFGujsb
43DoEl8mL73wiq8jFYWoTLStnnIlseDq7F6bF3PXjQ+kEGmlNwGmmK9CqrjZ
gjA3zgnQrqhVKS3tAkJMr9FvZaezcNWlUF/Er1ilYZG9wQkSj+EcWigFDopa
H7s4tJV6Ze4CRyH7AVg8k7L3U8s55EuJngc3LHnomaMMFAThjHjg0i0dIPjv
uoZlw0joIwtcDo55P9bXSixE1WKWjZM9ztVQU0gV1uNPROIcKe5ie6/ym8du
/lh+Fub/OPkQjKKxNDuAzYmPUgkFYJn1ZuCeZjKYshn5DLhgALRQ9RlDcgjp
+8xRAEviv9UVPPZa2XD4BMA82y88pYx0EjUQjkef8XaNTW9Tgg5mCEbRAQjc
TobnqMAsFkARiCgCRKe+Eu3e3aPwulsTQIE6j4oHoVUIPsGQCdqVO/Wnig2y
IkuFGsy+NXFX1uxuadisQg7guXAP79oYrzK9/N+r/QJvfFjCO2pcBT/0b8Oh
WQP6ZV1OrIoguhqTFvRvqkEPJ0REB0rtp7leqj1YBME5VeAfgqsicQekdUDa
EnLD7BtF5yQ6roQlCsiAtwdIpDWXcs9C7SX0OW2KNz17Lwjrfnm6oHK/w9Pt
ngWLsKN/T1In7eFt9VfoHxpHjjx4FFD3jzetRyV+z84jRstGj+VJrs/ahkii
vOzYdsZ/mA+hw6DzO/xlM7+6ZB81KGqhm6JVFySzXD+bYqOt5v2tCd//GFPx
UMDPM/5fdSFQFiVtXsMjJQzsCuwNP/PYX1hReBgktdIfQ65WRE+xdA00GSAM
93Y3BNCj1XhibJvv628e/U5COyrplZAwiZNU9jgReAOAiIJ/rfZmuvjeLP7c
NVfTRXNxKD1snoLjXx+VRobboG3LqUhuE3HHE280N2IzAAeyIt5/cdqMZ4ZM
A3ZCqee772Ictm8PFb565sDRXeul1VIs+4j5zGirqdkiifIYFnREToc5coxr
Q7Yy9geF7flDdxYDg0KqzskVIC06C5S9DL7zqYd15VMtqmvTVoNZZnKJ5CtF
55sn/jObnxpRW3WIxT4hAvz+WA4KJS1PhTr6WiIUgODaPMWIh//nE3hdysIE
OC0+vHVSGSo0FOjdKDQ1kwCyUEM9mjibwsbf138cuNy97u8BehE0iYFztK3Q
yS9wFfVE0y8KvrxvGP7kgGqtTnb6sk+dHcqLfWIF0QlbAhGOQaWMZpNeHBtb
+YVhXcugIyY7hi87mpwD/Du3QauBxMCBFCfTUhRO7u1C6s7EmOihUNHEa3dJ
4h77UqOHxv8LNZhSMjon0kefsXB3xpPFF0tfH4hHXn8y6rzCTiZj89AvcFsp
cUAjqtWZNq/z92RbJROT0t7aGcgVKYBZyUcGqk1ta9AeMIZ1VxBU3quqzWC7
QvtjICwwRJEltzexkDnL3G09ndEHQW6U2hk/uTfAgSVG4l+i1RgGANjXXlpB
VYW312V+YGYibNHREV/ezS0cPhdc29uw6mr7WZ/62lFhuc+kTPbiabkClRBH
pWYxrXtoYukcJrdXRAdJvCP/G5POHyxEV9QrBsWY+j7fSyAdhRokFcGXvW7v
E+qXrMcQYr23iDiYl6iBc19Pd6b1fktIAoecAX8rPsr5RsIcPl8IUTVK6Uw9
uAUHVwEn03/9ZMN14wV4vUwexf22Kqh3z2vVNj3UbEe6cscADTQxXNZBeZmr
/lnC6U6lEYdJbNS6Y4xPOrjBaxmVOpCg1rB/el5wJP6sGAQyGKLlqij1bj8b
72B5JpBIQWjqv9d2pE5L6l79/Ht4RR18eJ0rzvp0fcWV35IfCNWYMufo/eSG
M6G0tNtsR0dpAquFH3NuPe96gnRcAgdKSg3fRN/r9a1/6gGVoKmBjSCm0zTK
1a97CzbhydR9u2GPPCrWcC2gfe7wZj67Ls24RWhVzN+GH/1xA0Wtk0N2a7uw
Jqm01hwNqV1FfJxLTZs8yvUNU2xQl4bqQCXcLEc9qXBMmCBUJGxACJnP/fYd
7C5koAD4vPmw2MnnyRVuJJMAsVcPJf3ovmMYjvWBTk7IyQGvlJcf6l1H05p9
Uv6q+MPDAI8DEqFAW0ajRH2oDmZ6WaQYeAb2P5R4rl9eTPM66KlICk04KNUY
AFDvdqA/WBAlPeICP9C0+ZyPG5v+KMUv5lQOLbSxmybfaGSoPQF0k0vFWrs0
psPqkG7h0HRyUIyC7TaoAld+jtFV3oFZLFL3E1glh0n9PJgnFNzVQzQg5mlJ
PZArAGLBEhaUKDRHF9FqKyw6PjeX1OXDjrNj9oM09epiEcYKrU9agYgkIw+F
xA4tSHBjZ8BJ759Oq0HHGCbIYPmcvmc1n6y5Pv236I582AuwxPPdinbmkvch
YJmwMPEO2tKd4bCmBNQl1E8mYDIfyCcKtEB9mjMkWRe1Yp+ATtx61MyC0RXh
WeUV5IK23M7UjqZ/yC+zgpQFC9g7YdNWm54akhAMCfgsv5faKWBb4GxfAIoa
Afn5/QakZenjcZCdhNo0Xl6XkcasU/tv+LKlSg6yzlPTfticFM2bh5/cQV+A
G5UBYK5FC+jSbQJDY2FIM/P5Ol2FDrlkkyRsRo+fSS/tA5hkI7sWVSSJof1e
FppTcH39VbBvhXtm/WkXRbrMaWAeSZbqmbvTeiVMqJxfELcSOpzVIowwXl2Q
EFQbsWiKp/3+VSPvKSlo4kFALV08Nvw6X2WvpWExM57E/gI0tg1bNEpJkuVR
LbAtS7Drc93vVZyBUL29uVXLfALdHXyl//0pwIMubjCkIEOm0MM5zoMz7BEu
8CcAgOIb7zm80g7K+s7tXV9MK+jpVP8ApUTmKO6HBTLUlz4lF9o9/IXlkaaP
U6jL4JK09rrmZb05UB8PD1oN9YSwnfMn/TDS2D5yfvN1qCSh5l+fdzJUwOEH
Rk4u8W0IkXFHgnvFYE9gHDpDoS2oC68gOd3v8qHJfjH3sp0t1Kua0qLGc0po
joXof4K44oZFfxh/kggLSD364pB/0rdDps43gxocPDTK9hcp08YkDlZz6iJt
CX//NO7wHeUM66PmAUKQHRFontM3gpuLlZIz6rRSpPima9WsA6quBc4J0nTs
ZVWFiL6volP0a2e9ig+QDL5p8nchTaam8DT8JEMou4tlYXM1WO0tYz8/dWiq
pgpCIVXZZFn0A5nqaSRIWGcCja3shuboqI+wWuQISqcKQfcLxc01xqCkhhGA
XU/ruqa0cqif8UM+iLDCjhCz0cD0FHTUgSk1r2XMoI4E12toCL3Eu6sm0VUv
3vy1eXFJLtPaE+sB8bUCnBciCDevjGOl66i/1ABjU17TODvSquey8dnEIUvZ
TAkchURA9Y9x47jlHw+clqBz3AtHzqo2/WUGSWxEHkmupd+MeMj6FvTSNGSn
df0cgsqemR/yypsk9LjXSh84FA+2ZaOPls2PKNvSnZuF3o0R9zxjKBHnxst0
JX8WOACnHmyErDvFj0WsTbA3S74KZ0J72nhGtFlsJxYikOQYI+e5eg6JsgUs
FCthjJhPtGECPOS+9+5V42Q/qZjemxDQTIrZaq2kE0SZSLMAf62inn+2JKnD
O6D7cTscqGCzy5fiNz63TnXi8nc6F5PnHR/Gr6SwNq/mypjRHs4I6w5xzoRs
1LRAdpXl/NsB8HlS0+rlhav+H37s7xxvdG8xqxr13ourHhuMir8TLaFjN06m
hZOWt2RpXky3oVDCYbA3ZuVGRpTLu5VYrBXWHExQhx6Ep81iwA/rGMwE/7by
8YEJ77tfMFQzTaiMSUGs5TjTWEOwWQSHWldwjjllJ/w//ZPO5zF65LpnXtqw
DC15l0lqaKU2IAZk7SO6Nwz7t6OWiPTDhPxM4mcX7eedNjOH1GJ2ZzNTZ4Ex
c6ye6qV5Atzfa7J1k836WWOIDdbbI0kKxMGrsD8GbySMYSR68DMPdavvSGsa
I32rt3OrAY7zgAtcG1tcydJDlGutunKzWvZaqlGWs4QiKlbZd2bWfuFhwY3z
K/2MD5iVP8bscDnx/7FM9LOrGwItu/ctaw0eDPt87Q1KztuHvn4/yHG7WxYI
9NPDu2TGxQirv+z3qhF5iPwOffhDy4Z45ocKNVHyQxB5DTwQLLihK6ojAsWO
wo2Tm3JvSCBXJIcGIPwtacol3loQ9wBhk1urZMOJa/eYgFk25JRqETK1hx3a
7bpOt3B7GXx0j4TGhP1Cqu/P3UjqeOVdveSghMPME1aB+203QY2iXRPYjBhG
YBIAQf0OwYncOq/XGjCaUp+G3ros3rOcLj2CUpBRGK3pfW3oLuyMXof8h+eG
rttTRSky/Dk7VwTAQ01dbWkdk5d7+S5jqVwcEvthWUE/e3Z66E28qsr956FW
ZJrRGAf0eJlfNYNhQYE7ClkOCBaDW0IquyjJrVwllQt05Gq6eQ0OhkF0W4e4
m064J2JjdcAf45g0A6elinKaLe2q8+jdFD+VOGq64bhI7LL0e/nZKHP7LmAr
GH/5LJXy2aQndYg6qBhCzliz9X2aiKyQpszugp93UzlDSQiP8FkVk/B/3O/C
hIV+NmPKuCB/B4xBu8kc20cUlX78wIW7/R8F+uABgIx3mOSMPCy/uRcMGHST
h9iGHZ5lcIKOG8y5Kd86YX2jVqv2XV53dHGuavEMupWkcrmMeKrsr6f0kfe3
7Z3YsBg8xJMog7YTL9mwLZLWCere//fO9RWcfXXa4DjG4gVfnB1KpUD1bLzI
uQO+BxzlhEuoBmh6FY7tGlaO3BDChdMb26Jet+179UK4dgAA9sQN+ABiRcs2
RGTMtJfCY/YLsDus23IXCZCbcpAoZMjuA0BSXFedWPjwLDc/MPHrAkHT6fRA
t/G6Me+tssZxePGPBqnj/B8hYCl5+y5v7EEjJDvbSWyyUG3yEjjuewv4XFEo
41IilAq+fvKwryY4GyxDWR1F+VYUiu66BmdBUU2HcEFJJSbMvI3Q/3HQ3xWi
l0nqTOpfOOKieiglTu/nd4ccMm75eZc+ll1u1MchDs8roOVOb+hKdX3wG7+Y
bRaXKd95SjK8ZmBg8pGR6h7Xholf2sYqjPSoPawZBYGpw9LZOrMpxaMc1I1R
AglhLhsZZSmMF/KJCv8779tn4u6Rl6YF7ON8mo04WbL8GFkI9ROc9BQwsKm/
p+t1MO6oWQrtPy8g/7i3omf6QNctscjKCBDc/TeNiJ6lMfZm19jev1VkakaX
n5CDgutqmiqzPRGGnGbKC2EvgsEUrKA5AY58wg9ekzrRU81qpnUn5aFxNevg
Ad1bdmsppLTRiH3e8RuvHMpg3fvOJaaVImVuauwCJxcuygsLtqf3+0SLpKKv
JnRmJbuKu/vC71lISObrMHKawyLAj3e5+kP8AO49PUaFk0Bohho0dMuCW9Io
NpHtnc8yGMzPJl7sqIaXz/xY80t+wg7g79CHO5+dkMh31B027KrNBuMcqREd
xUYt1KHVG05odmBTTidc9WJM0d5Qj5nO3orm/mQi1Wl9M5LtcQmjw1md/pGs
yW1skgcCUp7qOAKluMQcTd9UxyFta1GjuOjGcf6UXbJuOkMypPiKrSFNHszk
EsXucl4BNxh0kqMIR/VrT7bDBN7fVYF/29ou2FYxpDNASVvx1+ygTUduhZij
sG7sb52oQQ4X+7AFmEA04NSgawuN/tHzWOBV16PndKqruVHUcRVVXrTl+JYe
UYlKAEkHxWZ5lLfXJDQjJdsFOx2UDRKoceIss7mhvjKZZFTdtC68VRJMJoWg
UDumqfHaidtZyBA5Qob6nbWnQL1lPdXhBdW9yCwPsmJHk0jrVm1lSquLb77O
1HhsskXJJ9uHXvH19k33lVkvkFY1LD+KBbq8JqCUqZrNNEE2gs2pvrIvBK+2
ZDZSyRDyAyxnJu+kjWyczFecgf7L8zfVqPw3rZGqm7nQzUkcBRmfNz0Ltu7v
Be2imbBDQk0GMzYhtElqp5uuwy/mJlipT/AV7HF34U2I0LLq+6FuJsV/Uqu3
PXwjlg4JJDdoWJyLOyPkm3PqdkUM3kAyPG11wDwXQybU1KHEOdzL+GfobdvA
pBH2/eszgNp2w0EJTcNKAlSbDbNNawtfAtSMZSewz0D/hlOWOcn1m0HhX82r
HcOOp0+PbUYylvCRiA6QCviJ6pQKmlAa7RGIVXInZBBQmC70k/w/YMUAtXkV
1kKKejDTXCBrUrbFTy18pDz0ONPVbembK3xub724CJfl9cAdp0eJ7dOo1S5o
iWZiblm5gLsXF5vmTLOfApmXpoeC9fPG83MtU19W1lcUZIVWfRzO1HwAbxKl
SX4DQnYYqawcGDwvVqXJGZWiEpDkoDX4brumVvX/IgtHHUajt9G1kA5K47Tk
QmV6JxiF0EG8Hf6JCXq7TLE61ZUZwM8iSNWsFqSOZSjomHSjhi3Ecm7ESxLr
T913VZ/b/v7RJ6hMdHUgsnfAxUI1IHwJ+ECbv+xtHoptbPfqSJMOvEDFg/c0
z9DNpdUS4SoBB1t6CWE7P3/oABP8WY71+HnjbBUpvLm3B7+k6BPL1OhmdXW6
7C8V00IwJMBqb1B1Pxfg8UTgocMtNWSAFMfkFee3QyykMBfeqQNleXuE3BAV
B9vpy6WBNElbzgOa/oMS6wOqCErzxTwK1xXFqY7uP/AYcnTNCUxqVuBX/oLH
1x30RlP8zHCC2DMjtnsZvA+MMu7d8l8YCp/xZocZdlpUeLCQeCDzCR8t3fO4
G4X2HaGu/GS919LvD1sng4mCngOi7OVVlbDIlEc6fBY7altTneuM5S/jH9p8
W5Ql9g5vUbcLY7oFVWE+ZnoT359SNye7qzX5k9PaQlc5cNgNvddMoUFyyhmM
r1bCQTp12tneT6FC8GkRXkeFDnPapH8u/m40CnqkjYEcuMwPVIcr8Alc0zac
NTXowsEI09CDWSgscdR9uByaiU1pqUv5aimCZnYGVq8GcOyLFYApFv1rEZOD
DDNbUvuBS5LbD4YLeZ4aZKewGZ3KDuTV4QFfUHga66P5786l1rZ92ENzK8zp
aSJkdi8hdWapTkduIESC45acCwZPNM7ermDs4zy/SHScCkyRK+Rf6TojOeBo
nY1547/tZllURXnlwwmQp1tB6YfUAmyBpOS+MPUbZOwLbM9Wi+KST0hwWKn+
HK0tN4T6pQV91T9vQ4+xXlnNqn6D/pbszMfYnIKo+E682hvrGqzPpws1UKE4
uGoMjC/ZUrTSKZzkRKTr33nC9Ud4TwGlqX8L29SdPN9FWEmTJfxaEcyEvNWL
hmageRFPwDVfK7m+Wuv3V7NRdqGKL9grRpyU5Ysc9mcwb5m6FFFtyn1NY1j8
AI9SELSD37mhsTa9ALsRND0lZnqR+VMOVkO57VgZL2/ERpo8mHm20SsFAMOm
+/ZlUkLFIZpoRiurr7QoDCrApsoevdZ0B5kG4UOK4ETcIf0NGPjBNOeKCgEl
MWBd/tlMOXsN5jLeSlBVexlU0AUHbDwnmSnuCRi6NYoI1dV6GoB1+oiRn92P
VsEw3kaXCveTGGjCYB2NuTRgxO9IznsuCcVwV2jJmMLIWf4/DoEkvdSqckl0
sT+dUWw0IwTLQ0ylZnweIgwODugktT9hTBw18i/P+p4xLwS/D/+E7d9pZ8Mt
uh+nY0zVKvehlT8Ce83dJdZV7TV7+S/aVNuA0teH9KUzHDtqpHtj76ZVlpiX
OqeMw8tyMnB32W3IKPE1Fp6zhOB1pv5Lx3MtsA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyK4EWC1pi6D2Ax4o2qIJIFB89MY1kWXrs78tJ31oemPWFG8tuvCS/jHZmghM7iNzVtEWotFDMlLkX1Q3y5PGwlBRa77hUsdRT4oTX1ktxotOBpIIF8GM24bbmTaNaudYu/nZEHjfT+jb/9HKws1xV3+P+ccdWodv6AUZkOSw6FBAMw4qpBxF3XSL0XxDUKTS4bPDFlR9h+8Ed9nb/RB3GrnB0+akaGrW3sKV6OmQG5FmHLj+5Ejuu8OuaXZOiXW9tyDSJ00rXhUmrw2yaVJAIArEApFR9bg76+Zkk+C/RYPHkqkx8V0UmlzAx+xf0b6h39TSQkXFoIiutkkLjXiKXU9Hh0J4gjEntTv5sTnvCmfWrSRoxXnKjNiTOz5BaHnhQl8xzcXNgipGJ2uqalSwHyQbUIGEeyjLvI5dfQGGqwFRi8Bn3igbpRdfCSvoHCtKI8zxV1lWAzYc0Xf43itgDm1Uu665ScXxhEG1KyQW9yg1VztQfSQs2jnfEMCeXFA6dZK5LZHYAz9DoIZNqQSqy4xLpRSx9ACd1FlAmMMSQ1j71u9HobYzLXyWl/uChigPGB3JmI7YAAui0fiuDuhQv2mbhygvEQVjSguZXbqs2VhDOq7pEna59ECumB/h2eC/a3MBJNtnmzBJw7mf9c/mPu0Xy+i2xgiECegKubPrnqH7aUFihbIRdUb9k+vDMDwajkSgCJtIZIDhTwaKvyWmUV/aNoF/nGVLf/qAni29USGPjQplCJo+jSfAbO4qTpoFLTfWVdmwMS8w2AlkeEdYaNd"
`endif