// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vriZPnp+WBeADrc8sNMmPFe3nL6S44efO4rA9ygHe2d/lugli2srYN2S0e6b
Vh663IOkNZBaGlxZvuaYf7Z9aS0pPCJ6Bi0Y7d0E9bZyJffF+cch+trcpKj0
ORpIh6SMIg7bKuFRk1QKOu82b4yWFsbeNW4Xiz+WVLcm7iXMc6+So35hhFBt
lisBAKF5gpB0srQwh/Xlmx8I+TqTEGO1TFY5INjVI9P9fmP5BA+ouwUXCgIL
ux+5Rrt5CWZCe5wGiRg7m2rxFddeLW1VLu4yrYXMqxvvy78fy6dl7PoBsMJn
pgI1u/29SfqtSXerf5YfApa/9+J74AEJxbq9azrBBg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pJsqVpC5E5HEv/HKkAtog3V3XbVsHBLVYsEb8wKm8BVUTYq5MniGDcoDt/B8
27wLWLFGQ+zBv84+tmRnvsNNqLUxAukLt7ARSWUiaDp9o2uLbww3DXGi4OBw
W0OfZ+04tUhmBQbDgN8GN91vlSxKeBBDkbtBfptIbGj4qMXGjBo+K7beHcrX
Gfl1FnTX5vgIjSK741TnOONxVz4VkuvlEEbowdJKQFX4eVJ2V+fM933oTq91
G2Z9chnMPf875tzHnoYSOx8InyPwNIXUtlah/KLf0dbWUYRRyjrzkUfDQCf6
4TQIVlCiJwJuGrx9ESJ5ZDeA0GvKWgtwbFZs5Qh5ow==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DTcTekqbRdfj7hvS+BEzudgFEOSugiEgEryUZ9xz1OcFCm6jX9bAfi/lcd3h
69JFqnGenDsWV1WyKq5AyFQAhkBIPPgQO12MXFrxqqGHwNRpu4LoQiErQ6wS
kinxT6AYGXF63D/GbtsNEfJGjdU5xIn2oQpzhTwYx/E7NsHGVI58LqySYC00
wPcRIlUruEOslCjjXR6Rn2rlfXVDC5Rg5ut1xP7tHcIBmYT46DVajHAjpN04
oFqL/IZkV/XVH1wAYYfbEQ8a/PcQwG8Sonf7KS62ZLVNkJoOT4Ki+0Ny40kp
oJGYLixhi3xoCPEHIYH8A0EcnuZ/RZ4nHZb7YMIzUg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bQUtNU8C1YkstUYrZi+RL/HzoyGly/GBtn4p+l5WTgwyLDb7Fv/2gQPx06hv
gxkHKAWKM8w1KrOVV4RIF2V/KYiB5qVOEv3fCQmyfP/aFIEJM9jtWGiprbus
VA/RQ7z1U0LgCHL+vVQaP1rABBLSptXG3HpDB+7lJH9/exDAfinIDbVNfEit
ZGmodfiJprzNSyOh+ULOqf6A0ByiGTjkk9gm5vVttuzuoECi8xdJeew1xUsn
4Vuz7BV/Z3GoNUiiDK63EOck2O0OVyWaeMGPDHw0e6qcYhXXTpRTe65lZGZP
3dtHALPHmH2e9BSSZkVk7GcPaQEZk05af742xrlyMA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mIcMSH9pXXdAhmFSixHQRXfH7JegSYc8XGv2F9bqeB7rDJYaD8M6HI8cf6Vb
saXceuTsMGVdtIRyPI4CqhUykVGRIew9gp2cXsgS2wBgMchmE+L8foK/54OB
bHlRBwsrulvvcj2ojHkxQA+tLkkfvBxJOKwZ313EWoaI0M8XjOk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xqvVKmhR3aFifOYcbiObmQq38VF1sTni2O9BhfNt9JrmbO4xkKBKNaBDMATb
o72bAYiJdHYvcyf2Iv05ZupiTACUg/5m+6dbojIufzSR0+R6sSIC/BAR+1Mz
CLcclOI3GHNviO9uFZOiTMTXWud1Xe/Uz93fq9oSRw38mcTgSpZxwMXWZ2Iq
sNZQ1hSTgGhbSyZlpp3bSkQHkcXAyzj1hiHsbMJAqCzNI+9guNWrnquPFKD9
NWr0qZ2wdBRIPJRLKZsU2eC+tpD9fT4C4y2LTX8/F+62iQiAoVdnihNzRPU4
sblbHmugryr0//7MDO2lTvMJ9LpL4wJQA3xSjj8bODGL8Y4MuhFz0SWnHMrM
EB6vSCSKDllubLEezGUnBQUyxsMLaGL8sec5cCCGLNrADE3jvltUWK8gnzlg
pEbmevfLKkowzmBrjo5F0weXKdx8f2Uaq3y0OxoNlfX4nNNoqNKfRRTZ2zaO
axarJyGFbloR8AlWzdw+eVKwN4BLt8kV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fDF++HsbRA9KsFc0Otaf8BwJiDmMLkHR5jVx/m5ucYSA5FFJ3aZ/KXB+vnNt
Froce9HhthcJMvWz1Ik2BmCG02Vuq6ASXOtgKBZNHhICeW81p/8jREKiKTgb
B9+HUazbIQp2Zhfo66BmmRqqV3wQ5QypfSxoYm3f7y6oIGD+oS0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VxM35jif0ZKpIJre2LqJg0gSXbk5tw6NAMOGuobigZuwuE/VAQmqW/47xA5D
zLizcBT2km/PFVScfn0snxePGtF25J3IBBeZj5Ysir4HZ9j5rNW1O3F51Jyj
OD9+zCf1FTpGi2tlw2FZCH4E67cU0WV4o89k8s5ZXZlD9nbk/ys=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
vaj35FdDyshg4KSw4GrNNpTj7FEbeEfcDvcFP+pqgAhdlE+MRUdwmI0kV+q4
JHqvBvWWUBafaHoa1uR6j9xS+xp4YpRzH70q3CGEq66cmriSIIw9MN+5TsL9
3b26pl8RY4lcZu9vHowC49YH0dNTUZiF1w0efxcWO9XfhcvFIl8yq7MTxOHD
XmIn2UgnPmnCvEqKWiSVq8xuPgslOmDi4/W0XUO1jV7CCpOMv1FeOwQAJmKD
Y3Xbo2nd6+otlqu9fZhusITAWjWnh5XGYsaCItuDGdzCkDK4B6p/Dfr8WwUT
1EI1FS64pZUMX0syRxxbXf/MBDwg9ynlJSM4Ake4837s+nzGHfcorPLoRDVk
dFCkuurNrPa1sUP/JS2IxjAYRX5yCa4DnuWY0BpO6NmUn2eMmUbCmpc3Bsgx
L2axh59yj9Sv8QyXtXULSWbg7b5jBLj0dVCbzQjIb17CTkrUsnAzWhHbZ1ip
tYUaoYcMzPzRNExFwvbtvtDOVm2cr1QMEJhBARE8FRqxFChWl+6TyAkyL2Ue
XB5vkgrOsDpvxTuDxWtUUoDMT9ccMOJ0t5734CQN/HeJJEu3KieEZ1nIARGa
rk9ymxLl0ukOybJXlgtuIg4aYFp54c7wwSWOh4DrXfJFQSzpNAa1WVvBPx0a
gNeaQmiICVtxfTs1cbQ5HJPExOOGkb38CYPFzBy2NShtO3L/uQc3YgPotm/O
YL1jZJ5gvDyESsC4/pdbbJZk5W+jXLDEmhIx0qV0BFofFmynvrFl+bazAvrE
TZvr1VEhwdwbCppI77f7zDTT1F87W7RNT0DF4G0cVpq0aaGM1sKH6c/kVg1c
k8YS74OTAKSNLkYhAPlbKgjNtsuGmkIK5mrDirfd/bnBAKV4KiN6JBk+bNQR
bMK6MZDgL7HejEKB+4Y3ASAWpSLaLPZrNrPV64IoAS0kOybehgQ+FRHn87no
W5ysMarqeHL5BDqvBVmxBPpjybeQ5gh2c68rjsCD7hVz6Nkol+99lFXWDuvB
TY8wmfZfmD0WqAKuKLXbBWfgNS4iTcpE6zeH4ueHN2DAoCcspV8s4hsjpDBl
7JrBuSbMfKfWTOb2IObfBdEOPBPa99uGE/oV4nehs5IKCZszAEb5l/tSvljc
1A3jItcb3DXbLJMMszgSNqnhDgOuz3qXbU8IzNt/l4Cj8WYONcYlGqDAR94O
FtnUINMdQ2iaLgynBuHZT5Z8JVZk5zkK+Y7RI6u0iDShNT5VASQQeZSBdkx+
vL6lHPk4kdbTb4USrdLZGwzofEyRQ+OMBLwgdmvyDTICN+Zi8xMEs3tDeMmk
b/aCSPzH+8bgbckHMCnlYlIuhIVqpDrNRiRvmp9AsD+UhCjb3h8cwQcfbiQ/
J6WTLMrvTZ3EwHwq3RjbFfoq3A67t8KoskXbLHW0pEFLMv8WJGs9ltHeGaw+
HVkyeXCbmKQGb8F5YtEs6SSIZSE5d6gq+4Mak9qXu/6RU8OSPq4W94J70doq
pLwkI0Arw9zPFxY0W7/jWCOUtTiuLVw01DyImKTYH9ezoMAsLnPY7ihmAttG
7BtCY3CvKRdYJ/ZV4p6ZQBUJ0KNZmACub+k9JrKJWWLajCRh+ClCfO3K8HIj
FDiCRPuc2qMyWYuTIliH3ibHZRd/1Prh659TFn69pve2cn9DOosxdDPdSsrH
Ci6u+JDzEwX7dvRL+gRBxU+Mzss=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeg2exSGfSY/ilai23uepJ7JZ6IDx348VBvwZlDpdGj4AtOBZQJeUtVY2y5qFZzus6pTHuoSglppT/0DY++s9FqF7bvhvhHPSuWtLKbvZ0jYA1OSRsZI8bJuqwatJzqTSv0r8tWlUN0zAOk0PTM3GNgpnwFcp6B9A65fCiOJ4a0tAx+GV+0TTmb1WYQHiOWMFVtAgJjsZ0VqZzyT3B/gxuyOCdtQyqCO1sJ3gFMsTANAJibxV6+gu7ZAQY8oFjB5w9G7lHVnlW8uCmM2hxa9uvItTwOvVzuPx+ScjQ+GI09sJiW16era4hNl5QIebobJUAPbgoQH3LmUE9tefnVVg1EAE8vVlMB4n2+yIfOd6Sw42BtS9VDZAXBSbo48Srd74+Kzi7Fi8fAOFESaWwSl2eFcwXlUIJoiG4pkOfGC+loFAWfW+mLctAddQdZEdoncNBASDbylpULvBMzJq/Bt1cFWsJ5S9PGXvK4o2rgYgiCox01NqCml7Hc4ncIQwR9d2kiDMlToYVC9f4YIM2L+L0sA9uGL9QlnHemlxo5Spnw4bafJ1QLRh2Yi8iQc9OzyK2QvZmwV1si0ysU4JZ0+gzAjYipQWJGMObR5pG77Ugk4wlaCo8YG4VCFu/1mBdkomAaW2jo/aUlt21LAca79mwGftr+SfeIv6ahbkLvzB//chnxR8Mxer065haqK8fPyPp3rHAN67Udz13GHC1zgv6jm4dveHLpl0yPIq09eWV9vD5gFX4CgcDx14yxsOsOKYf+mh3LOssPkcsmyKBqgwET"
`endif