// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RvdgtqVVQgZRAdSTX7kZcZ6s5rowf/SmiII3xrB+avmuyIMD0ElBB+3ezJdC
zKzIBFmC8t4gQOpiwoo5gTs6eLZ5EfTQTneG0fjhsLty6haZnKecNNBOXiuW
AG7gmDMd5D1tWCgEgTfyf5fQZYzhQgjHEpYC5ukO5u1yRZWimeYKhrXsXg66
BvYNjWVl931SSdyhTt49Mrv50fM7NwXZsIzZIgUIzrnDTsBi5fnltBCeN/U/
L1NY/E+SAVAkDL5FSyJWQilffLX6OvbulmRwS6T06hvk9Um8U88poyJFPp4c
qCbc2ebeWawxnQVo5iqen6WNEallpAL126lvy2ZRKQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AQn9GPp2RinD2q57ntZ8mhYRFJIKPrcIu8bRbsJauO4lUykyx6/E9ZPShTIF
LsXb28VDpSo6UgBErCMaURWjn770NIBmFrBF0wRWFU1A/rt2MGDaRySFsTSM
SbelVINwM/MYPC2hzsOnA1OZSajLWh8G3NNnatadQ/sOp925SpCbOAkYiGP1
yy1g011DXHGOsvS8v+MuTh3JdQT+nxBFT0IMuFRKeVA+d7g++qMXbqRtBwF/
M7GnFTG8anffzsPMmrYi6uKEasxQ0nfH9riZGIQ0H4pIxlCSCSEKllFHXWL6
h7bhuEyDDzlvTUn9JInnIQmYYBQPTHgs6Tmw+ZMxkQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nIAKBvMfvTQYEtvoVmnSa98CW71wDeYDyZEk/U+nyM2Egt4WoI8XYEwdHi0g
xOL2CHvR75m1nLP/KpR0qruqomtySCUkTnPy/hLXjrwW7JvNVynH5bhIZ4Kr
ftmRPt3Xf0KyqNUVzI4g42SbyZhAvqm/gVhBBnM9+qytRj4RYKNSbI5FmrYn
FT9T/Vi4d6cQA04CFFlGT+IRKSie8gCFZGD6kalkFNEiHmnuKRVa2zSevDZD
SXHbeXpiYy4CD+rlHMThzVsVxq4F5egn18CRSDlGRJN+tn2Blb+q7xW7AhrZ
0tHB2CPTRHgOyf8NTNmfWC1j62Evk4dXSILL76ppxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kurvezpQMsX4ILtC2seuwtkh+WRCXiTydQHQJqIShcbZlKxfE0g5QFDLlgka
w+2FqaPjhQmZJsxldFsgbXuFWNlO6TJFx+3mTwc4Un4Zs2CEq2Pff0ijYVeJ
ffjPTt7sdIqiGI5liIjfwcqFHGBUsLWxFmM9jrXeoOzVtEReUT5VKysx1cj0
bS99bEICdn4nuaviUVQPcg8hBYeGvmMaakQKpmZYLMOiHUCTckHkY+mSpHli
zXbqWqlJOdmCz4/kLt0NREzg96gMZhhvO41Rlr9u7+74N4UQEU3QSiW8bWmt
0XWBuzLqaHKGTvOJ5DAAmEyTOi+9fIeeWad372YPfg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MY2gilJqxjehOhb9zrn4CmqfUF3Q661lfNX1c6HGcvelHj+wBs1CelMabSaM
Pti/xx4Vlrjh3bqVSLbO90z1TpCPkFWopRo0C4tjlTuPWoJqLM+o8gUOcXzo
2GePIxadUZYck6NdnYbVEqYVRQmesHa8C0R/NscNK8etVs3EF2Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GQwFG8W+Y/V8EGW1J94PoBVShCTN9vVY3BkEfhs3TzhHoLmDXM7bapAz/gEu
rcp0KDaP3Aq7wufQ14Hka6Tgf1kXft3uzoAtgsvd+hu6MjDlP6YjNDCIGZ05
6xYo++JSYgOQJDvc1RSYVUs3q0NKC6phxzqZmDgDb6WykOPfmzZMG691T8cS
8AJMIZGB7Bb2yL1MGG1kHP58eczBtOPnWy69PgDuOWFa7De5q4JzK5LHbC3l
1k+9bUhgT272UpXtzRAspIKMNRQxp4+Nc7rHefs7LNYab3wE8ZsXxI08P62V
fe3CF921rfMmOid1QDqvwggpxYLzORwlap+BLZEAK0+Nzl8lQwntK1RItlII
80tf+hQXFEF5bBD5o0HvirufQqvlvARJihdJtnsEbLXOqUOxVQ9Oz3fBDczi
l7xxqyu7yvQaHuhnCT+NHrSmHIALTta04OmZUSjsRTfOIyfazMhY9Z2YI1bB
KWE2tA6Z+61JN+xWPU7hPodRVsDrH69W


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BS4t3UycGXKQX67Ynx7i6O35Px1zWbpEoeTAYDeJ45GBpdbCdalnkA2lkWdt
kStCjIxlfAwJ32ki5SD2LQFdAeWKBBWTd3XpcNaymKrSFAB1RZ35ZYPp+yQq
wcXL2jtiN1XBSN8IYLfSilHyZPoIAAMxJ8in79qIsZcgKeYht7E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BIMh/j08tAD2Waae7v+TdDDEB/ikthb33CJYzsuVVjo1gM7Y11NYl8B1Pyrd
u2TOmg1O98QszoejUOsmdI2cRh8QlKjhkWduSr3uGSKfuNiz2lxlxKJIlDUx
0xIxUMQQkYAOVLxzn6GP7LHtCLU7m6BMZ3ddk52Eoi0dRlE2iDE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1824)
`pragma protect data_block
mvjxMm7kl7eG7oAQwH9jOl2pn27sSs0qDcRtKkWXuVUCQJ9H1HzO2eGp4J5T
ZCQ7ipJyXnuHv7fmKzl4xx+TuM5/CoJu68o44nOTJYqxX3Zek141k1hEQ9aw
SHjtQ1yDOcIEqmSwX3aDAHCAqk1YZ6jSl6tXdcjGf1I0hC2idNVtLRT3Lc1J
zwDVg1ryytxXEHVKDztjP0fodFbYkvZKKACTRiUjQ3L1LJx5ifqy7+O7K4QB
BHWlpoqFhaCTJ0yrjp35XTrC3DZ2wHgxx+rk082EQzyx8p1m7PaKoUm4BrnO
hbRrjkVModD47lKGO6IODA79DFo7k1VuCZdB6FO2hfdbT/QLDLkS9lw0biP3
9ublOpwjysUM09/vP+0IEUmmvQX0H/4wQvegPWQPbyLzdBQNQL50LwrUsP0I
1PqlECgDoRvJnO3qx06D24YdbIBuDtpM7ViyLcmyPVGVRGP/fOeu4tIVTazX
i9uLW1cUhBBJmRS5jRDRjnrkUACPpaGrH+y/igOyUCdviIK01O8P5lOcYw+l
v6jI29neWdHNEuW4nHlGU13Dk3aIUvOxMi6yENbiD4Gx62168BeKipMJd+95
6QN+GGLIIXNKg8TlVqqoOpos6xUj6QddtIgqusZv1tmDPmc/B0E65+4DBDL4
g9v72jJIGaII/TrXx49pcY3oII4z4Zyp4AxswkiKo0QnoYvsDzTJCbuqmk7A
J/qJYYbXOJxPaM3Fw4IFo9j84S5qwBqSUko/wdgAW2smUBaARfx2NEXWCnfG
H/ZSYC6gwjukZ2jE0aB2oTj586bStldy8/mEeqTIV900hKxXhRMyW4Hw/2LH
Qr15pVG6D1mvEyvUPPNzoBNBjofakHObwdjfKdg+GaDzZ0A+GlGTJPo9L9aV
w+yvm/RoSPjOIEgvhocWn7cTzNozqA0+MzHH674n8mGwQ9Al9fTosQ38D4df
L4MG6nK1RW57puri+LLPmYwk1/5fiQNxmrQ6ouFWHiIHw6wfF8SIWsj5k4iq
2LX5tu++fUst4r4258gkGjAzVQxTLAPHs5oQXiIgECwWPct5YQqwJDSxSV5s
0mR3/85hq1JGn0//+WQLkgk1t+38g6E7r5hiPYsRwPIKlmnnqsPfEttiRbvV
6p2+M7iCa45zR58ouaYWCOFBB6cob7QarOAlMC8hcqz8VhG+KKnBoN+8PYzy
jeegAoimbQqvOOhyJBmlpyXqy8OGHGhSLJ4ErxKB6iA8RVLsOdnYrdlofzds
MhlNizu1O2k1JjZWMuRWJgLd4FSRR7R4nn/K2Qp5n024mEBNLCiiFm/O8iKW
4h6EtjoomQ9v0DoqZ6HXTdk7Lc3v1Wb30+KLXbEuj9tACtrZokYN4qEOIS+R
XzsPhqFATAgU7Q24xLq9LgJIYzrROKioaDBogXqI3fvsPwA5KUWYjjV5fkLx
hJMfL4Tz573Ls7Fu93tHWXHBZbiYf0oCKHPIHFFkzhNpaL2WWWsm/nEIbkyo
oeW47LcA0KMWJyYa5pYJl3ZUic4OxIkpj+WTSgyq2ttyYf6556DI4QGz7YFB
JoteQ8C4No5/npOOSc5bzDzsb2V1FBBDP3oJ0NsnGovb10MFHmxy8UNlaOHu
9tclMv2QMmpX5sjFVJAlV4ydeM3ax5QBNNQHWio5RNK3mlaCrtvJDfn/65/J
65RAnZtSYwpKgSzm9+WE7WpthNJYnqoasQVkxpksst26lpBF1gNrZ387Am9E
2KHSXhuo4kk980hB0cWpt+NGgOUvA0ZpjIUxBmto+ztQ2K89a3uH5cDsnUxD
9E+ADCH/wugemQG6/zRWTCtU6SKl9JVJItvkITVvqyJCV3x1mnphf3icEMzl
5e1PDvCZVTnyv9CDvFacd1WFNagJbueN8YvN5tDalDVChvjLzyhRQA/Lvfkx
ZNhRjIZkVbwvyPOWMDk6zwRPE0c5tLJvRdwTUhkSpm4BHwU+qCHcfRX8Rn3/
q7VjTcXNULPv+1ayqIgaINauSziWRBNXvS5MfiEGqvviBok7+h6H2XSkcrbL
DUPnbNQVvQ7cOg/jysLQRzS+c3t6geWlWNF15RkQTsF7dsKxEccDl3Yyvg9h
cWbZ1/ofgDoRzxrvlUtYMdNjWAeBrq0o5RAJyCN83teLjaYjKVPicg9O0vAo
m9VTrhum/qLkJRZoQFNd+2eYiiOg1QsNII6D7lmrM2yk4DWZ2INSKZaZ+tro
hoACpib8hbtZpbjgmyZ4yFBDE29LnWU8oSVYkZR3XyxVSCwD+tJMp/U8BeB8
RZxra87uClU9wDZrbp0l2EU4xHn3Tpx3N/YE//u/MhYdiTIn0pLqTsn7/O5I
24DJOnY5XJcMYZbybN247qaEict0jb5y/NtM3OYzcbvoACkBYoz7P/flhRf+
TxDrV6FbJmXndt2O7SUsr/zTO6w3rfej

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyK5kLZwm2TJpjjgOMnvD1btoqqxCmfSJ7bQMDySnpbgLCKdPmxAkyQsGWK1XLAvJAX2h/U+jeVH5Z5kP1fRmSYKpaSMCSG22twLY7JEjNuFvnzj43REpAH41g6EbI+7duKjbnE7okm65KJPb6h8c91iBWsSJn62hb7XUZddX+T6CCXDBG0P4Y23cQ3CNPyvlzNwN7sGZFWtVK+tIwS0s7qFOaRRQfXxm29bcMeiq73mjoJYRgh4XCXFDthGROsvhcisnVmkM8becvpwZinWvuBDYZ929DnjOKXLlQL9e96mLbO6O5r/GdGlrqshrIUHmN0LBMUrtseQeJCaWeQH4GMtwLVcgUz+C0HCDZ52gQIc0LPItNAKfa/CCzHuSKRNnAFtFllfbUpf5AKjh3Zy/d8oMeWytTadBTPgZws1vWMcti/Kxbhc+UMOkeukq8omGMJBApPXQrcFNXjiSpCBujoAYcPvYB7oONhaSWnqbXcWYzmgDI8I55lkZpFABcW5CSu4BtZEJCCkIi9eNJCnUsX5e/ejYusw81C5bUvrbh6T03ugvyWEemNeUKF/m/f6IH5yqesq2Lt49dnzowAr9ihSdSaG5lR2Fm1pBLM8e5KuDTzkQEH9nbeq0249NMM8OrBVUsCo30f0sM+wTrloBitoGLnpv86WC4HFelzDspHsvfkQcvQporYHkEJuFClucuC6NjNTvHZmC8slqwqw+b6/nrF2cHPQ7D3doz3pfI/j8l634LzAO6okN7Mw1GKAwhF2MDtz0lPMigt0HA5PjbEJ"
`endif