// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X2eeWsXH3Kw/LPWA9T8qQ5FV+BLnSJ6gVk5eds5d/MFnGBRwkwqwLfoK8qby
yH6SJNUz71gioS3LIPDrBl2aIKMR8VZ+jJ3worpwvlkHYPLcnMQ9rASNRRSJ
dNtFEBWepjuqzI/rEct0VEAgHxCw5e80xZc69YmthrMiR0hyYjP0dZniVg25
riWUh9KhRsIL28HzAqCnexLQ9fmN2mwlIDGnnAQdqOMmU34zKVUjkG3hATCl
T+NZScdOcmX7cmfOGt7/iAsAGQe2b2yfVhU6Bj6w6TmqykXlecBV02ZnNsla
UIpyGejri1PgGqoUAIulj0T5lfcBFyO5PH+ClF1GcA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cADuGAC7jHS40Qzih6Ju42NpDxHCsbffGJQH5ShegEkbUAWdyYWf0hZ7mNZN
dnStw1PcGBVVcOq4LNmSVJcT3v1I6gXaeqeQ+0YakLU+FTT3osKZGv/bumSV
p6V1DnnYNz3jZouUXFn5ZzU6cbqBIsJn9K/Yyda5gBgdJoZjVfGbSqjoTTti
ma+9CvXJ9PaUtz14a+IDcEe90uX3OoyBmFxEl+ramFdlwBbxfAcDcDFXwEUI
xsq/hsxDmt/8zd5GuZ+7156wtsZGcIbm4bt5B6qcAioHuMYsbRefMUW2YCXh
Cb2UphGCyfFJ5AC3mWrBRH/1o+FFaIJ8p0JwlooBqA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q/mcLSp/WRaeRImhOiFeFoTmTYGUiu+Z5XtQwy/mPGTsxdqak8ymaSAWHecp
7oS0hATgv3NJ1NazTZ6BlSRFkzb5fV1aeUJfll7raSwAjYDKP3AaLzQNE/Mt
6knsr68guCrNd2h5vGpQfsPkeivP+ks1whZsRzcVVE6+QFDPXzpkgrwGInpG
bN4COde8whjQ0XvbinshTAz8GzzLOZMwKMqUSZgMvD9RIgZ8cmz5dnv8T062
y7nE/8spB3aK47pneLh4/vS2nPs7O3ab99JOCmKZ2o8bXOhr1m43kVqOxURm
OKMW94hs/sZgXGlRO4ViFusnSI/ld2XeWFMGG37CsQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nmsQXVRCtFhuXfU3gmwWoNr6Oh75ww2HFOQswc3XrGrVWdnPeLH7UXXw8mVf
sYKZfiGcc1wU6rorrbxLXZq3J7pSRx1Evt5EqsyvfVoZzSpLgN0YB5Y/yN43
wQFFEyZADOlsYE9kLjnd45uIuZs6pIlFpm0TGyHH7/u32iGa2g6Eo9FdEy66
t2hTBHMGrdV4RMd6UYE5X3Wrv2X6ZEBKxUKBWuV9Prp1XRm8T7CbyJDyYo2Y
AuXvNy6EioKfq90u+TTZ4IeYmMSdBIfWbyG2T2jzKnTDcDSYnItUHCYJwlfi
rOzRX5likTfqAcdZ5hGCTYVB45iAaV143hNZYKijZQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GfLcmQGf2RthVc32Gq0jkmKQgt4N7X8f5OcqZZGFJyEutbvjWg9TFYqRIPfL
77P9tsaFgTDrv8MRa3f1Jx9OKwwyDPAqbmA9R5oHd8TzEKV/PJ5jMiv74gVI
Dx6Cals7YPX4LQJ1MmeAIHpU+H5/u8kJbvIuhncJpINPF4Ve+sM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
StysLK17avqKtA13yQcq9qoaWSr+lApWMGSMHDCT1d/0E7hEmt94lk+wU2KF
s+9WfjWHM8tHnNPRTLFE5Pe0JmxuLarIeEqrjN+doojHw5bbx+pn4CI8jBDJ
8xyN1/SLYopuZvvCYUqV7FwC4MkeOm24DdSUM0s8zD+tJ1MXPO8kzzf4nFvo
JpkzgHePCs0aup2e+49+PpNFK2zY3Y57QvkQxK5uqHJ5PeL0CV48LNsll3vO
Fwo3KoUSavaVPjPdITnehPJG+Iy2bjcPWZ+Imlo58csFlr0UFHMl7eA8nfAf
Xwo8ug/fRTSt3MO8pFWzI6jL2bUSE63hHftnv+phKJmguQZK6jDlDV4nCZjm
zAXpKGcxSUbsjFUSCopkqexRLbz8w81TsvnkTrLvMbypsIUTYMlw1tW8Ue0p
hnNE7niQUVsxn7MkSTw2EJW3q0IwjjvLpvnHbIrOPKmnnjR6wsTVweJVEF/z
rI//uBd794FsSG+lfZ4Jlg+JG//YpKiw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mDteQVz3cYUWYkSK5L9uADc8vMEZprarUPeFFni4nard5YC1OfrSnSuOhe5t
vX54N6eqaNx34+VK/eawjkJUm6X5ldjCLAGJT47jbPDxyESzaQqOGxpcEPL3
jVJ3na5FaxX+XlMYvNinzk+oEWc9j89cWPpGdODJmUEM1jqfG/o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FPO9QVwKERPp5LK+0etJs1MxAFJzAhWWVUCt/hgSisN1vGOXzzRq/4Ti+8Sv
O30MMoaWng7nbXDt2fnoMdEMvdU7OpzOfKZzc0m8auXwr9EW9Y/RkgenFxoK
Y6EJECZ6OmYd6R+r6osxctoTYytXl1avh1nNAPncsFsCudTl1PA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3008)
`pragma protect data_block
b3hZJIhYrtJEOFGJamOY60R4QudaWO30HhO5xkgF4VYOSgOCdLCXtrVuo0TR
ukerqbQioqaeOs0b14cisWgaBRHRiWlATPzOQgyarRGK4Ul+2O1ruLdcRsJ1
zuAkfpAVfT9Es4R3CwhKDBDLdTsdmNiNPy4AaYU+ZfyfxoZ3kGpAiOf8Z1ML
qbDd0Yc8hGvggi167ETJp5hG/xn3awUd46YEhWfIDXVquv+OYJ/517LAaF55
nxtdy/7tr0W2G70DsyjE7Vj/JS//vBcwz7Z+33rqo9P/+khpVSEJachDNNVG
NZG+wWGNWjamRxEK0S6+XoB0kfd556NWKTq1XpcW6dR1dBkH2OH/foMgTjP5
Eb6n/GLf9/rH+ZMZf0NEMHDSKuIdUpVgiaqeCSkd1yjd8/pE/RgOeBqnZ7o5
/S8OMb0VWCXI2NdW7ZYkZv4L3+/KY66o0oSpGZSIgE3624468cxI1z8QKGkk
V8zjhc/4JClPWIE2UIEbPC09jLykVNdZncd0AmQqTGo1Tvm4EZ++zHGQpl8O
sWaYbVJjF49iQ5Rg/At8Ol7vzA4bMWAwlXV/WI8BlPEbv1s3TJ7fouFeZ6vy
d8Hp5BfJXJcQWh8FqLpg3AySsQqXWpkoC07l5db9+/a4wrBW3v+q9oHiNJ5k
d8gPnMQG62oir4FQwPEgbPE1APG0pjCisXjivQC5M8+YHiVnP4OQFCja7k8h
9ZE9ovu0XIAmGWnlXOf93IBEaNZYDWtsP26EmA/K6LzjLW+pB3y3HIR/g6ut
f3/SwdYspowo/kKLYR6lNuKFqxJe3JEBJq0DzXbyRqr68JSzNgV17Fb1s/VW
OL2IcULkfPF34Kvq8hSy4E1Zyt5tVZly7ZVwxsV78smdOWIkKPUcgGHVXCfx
XZlcs1UcpbPFggd44NnbKYYq+cpEMSFwol/ekehQGU7iMJWpjvgyVWILDwnZ
+S3964/xIieQlyoWVA+zj9PYIPhLZ2qmL521stfjkLgBysVALx8fTpFpepFs
si/dhC6Ef5q+QjBW/HOtp/iu4/aCCtTV2a2/X9uPD/Q/+CVm1a+G95Uw/KFI
w1K7/9Geyljup5b0Wqu9Z+dY4ec+83MDpBgft0s9ybkRAq+eKbKBuRhjUxgV
Zaie91Uk/jfAcr0Atmv+R/l21j/YMS5A5OWD+WD8cjX3PPCqg3BzXp//mGSh
1l8Rzl0ADjve5icnUKAyzrSL21af0OLhvYJweQ7+dwFESN1GKVlGhKK41EUL
Tf7MLcpihIBoMJ58mYDotKm+Xi49U2q6xA3Nl29W9j1a8F1xjOdFRQqTXAm3
F2M0KJtvIdRvE68QWcQTiioWMFiuEk9N7TlusIbfkJIiRjwTKHFzDA4VH45y
4KXzM9H1cnWN4gwj8sdhYi3SpYxX1LvqBIk/pEyL47q4g3HhqHHADzn6h5DY
pOEPDZ+LBeEU95HdbwOUcTSUV1mz86iimLZaUZ1S9U+DWNLDxkQGv8t8vxGL
5ADj2nNHwHcAEfX5vXhEAjHrz+BcRkL33Bpvpt7Z0oQygl3s8ZT7I1purfDF
awsIhKWnuHtm1dBvwxk+DXUwdXELmvyfmGvrF1UVkRKtD6Bx7dAiqkYXJP/Q
3o1VlwENx14lsMov7ticXNvDv9+ema2jsHZVql+rj7UfP0XaQQkbB8p+dql/
eW/LxfOtE9VWis9qgs4vrgH3i+PtwvCELIdjOCgFB/zb3iMvFCNjvKWp2uVT
SgqeXK5gKUJbSY4T7+CtnbJlQNN0dQyucBQhJ7rYaBnOZ0wXBAo83/gWx9tM
nvA7WlRQ8ySmN2GMwf36Vf1oFDMt4cdJF0VdclTnpSruAc8v8CdwTDBrEnEX
40gvPelK57MTDbHiwuRCJI+m95VFgGCJNJtHTmqKu5tZfXP3e8VaIoxtkV/b
M1tEaXAZuXMSKV+PEvWBV0yi818AXAsylCHEE6uRAGRKsYFyiIuCRFjbv7TW
RKe7faiKJnBLQDPEprkDivlyHbYyZaTWnuzrJi2OR0v463+Q4H632XLCztKb
NegJ2ElEWSsSHssbNNoZlk6PF0GlKQnyx4tGwWXjKFmfNcew3ljAPzXACUqi
HSVjDXkh1fhJLZ0Rj3F59aCKA7L3ltLO0I9TmYv3M4SQhe8WCmCA9Oo9MaYl
N1Qk995D5dp4tvpIP0Ganbmlsi95C8Vu7khIpJ3cycRwZFRMee2yYcGtND0F
pjsAzY0b+AFqDZmIXWGHHMxjZAJJg7CyIn1VwQA1uHEpshgCxMNJDK3IAPWI
tmHrto2jMWdu5huVZd1lbMI88PpPipxp6n0klWi8jhffgIgEod+Bzxq2OcmJ
inIF1r6WZpPFJBUqKXaU0EoHlwCLmsIWsOw5wiy/8SX4vOxbxp5JbY3QDu3K
ZzF24LC2Yn3nGnbUvp1uTGnYDXWZk8MzGMu3g4KGozr3AXxESu3Vl5RjEWE6
DynguIJsczfDuBflj177Ty9P8ZPyAciO+Ylad93Gb5ehByy8Cd/dPsPHImSZ
DIFeLzb/Ls8kiHvm2uvaGM0faTxTC14VmKRdBTZvQF6zJ+hPLyXGVgByKm7U
aTRj6fEm8DUYCjTh5mUVF6rRIQTj7IwKUCgRHvelLbqkCbcwyUEUW+cRb4fS
qG4Bv9yOG4KJJ00rmiydjDRg4yf4b2LDVttpiRcQPSq4GzPkHoxSaPBnuqaB
TUov5/D3fvFsmVTUKZC9kJP4auAV/5CaV6ZzxCN8yUHOqUPnlFdNTA1FPBVr
etFrr+T2yoIpmbUJcdvvHx32fH1PzeU1PwEgk6FyqHopuJm40F9KyV7B+6az
mO9q2YK5sTxTgL/kpq5i/V5IgjtEExOS7qlMyexDege4N9M0wt08eCY66Y4t
Ib0zojNMF3GWNj/qk32oNaKajdpb75JNaOBcMqGFT48FcpgSpolulHpc2j0G
V6zW+10TyhlMGWs3sb/oDxTDmBPcJGH3lXKatrLtysNWSu0wUMYJy/hspEHK
W22K7Uk47uBGCcaS2ICXPbNLUZixjpYdNuDywtaoJorX/Z0womQmdFBUDnxp
lYVE2spoKN1FT4mXObejB9KEP0Bfn7LuIblT0Xr8TWjEHpK4hKgA2rKgq5UP
iurAPOWYLW/kHdsfB4ZN5mrDOR8DrNh6+LdVd0JN74Ng1lF3GPgw170NQnwh
Gb7LSOmh8vEz0iNB3kc0/G9IMIHJPxNE6ehlbZhb3ktkVOvnF2tdEu7tvCgQ
vM9Ty1DPUvkOFaHOF6T45RJGGjnU+kASKbxt+Mm8ge9xhTmmH0xdfm4EO3XE
g5OiBdJLph87tID1Z5VothaCua5kQZubk+i+UYDO6p80eXIcY0PWAcFFVUTs
Gx+G59JEuRuOFvolRA7ncBOBGHITIMGRRoYXpEw+dG8NWF9WExYCMVHNLaWB
ZJZwwY6hr1XHlpF6mV5QUl808iWq+TatRg4FKuCOGq7GqLk9BobmrwchyZgT
AcFX/BsaySIC8NnJAF5X4A3Idx5HZlCTA+49Q2SpywbrnlXEDunJsdT8aLwO
fNRSg7sAbwWzj8lnbFv6Scjyr/3+XklrOUqUVMG2ZylLc8FbHAKhdFEpW5YG
5m98BZrAlbmCB7tJ9RVSwoASgepk3n+BFnmyZ5CadKdMF10FbZLU8rpFo6fJ
ldQhfjN9wLn2UzNeaYSuOAlFM9QdaRax7sIhPKNnHrwQU+PUuOrFnfYZ0o1o
kXBbKgJBMEbgormQfVb9D5IDwKFiAHS9+qtabp7pzDNwfP1/ZTf2flkxRvYt
6L9rRnAOT7apBN4nb+0SNuxADzTiXysW27H81jXIcUqGb2/qq94YSJA23iuz
cN0368rAXN3TpSLUp1JW+HpSMYkGh5lC/SyReqpEViuyiwEhofdjkXaaZoj2
WzK/9Y+YIbBaXi0FT1In4otCcxiholNyNhuLlepDP/FuvLnC2Y5hvx8VlyDi
yE6RDvGOEgjvJLbNRehREqyVPQUcUxU3/A58YWxeJA74WKV1EuY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyLamA/MstiUbdciFbKk+V9lOaHScn5Q58GgVSb9b7gUePul9VXoaFIbXqDgkCH74Gpq3lNscvgIp4nqH9NmZGYgS3skRUcqQ2hTKrM7s3dbAt5okVRHbOG8xUizRcPDtg0boke33LE0BL8fPPWZ59JaOeJnGKjX43faDaa+eHk8iYkgH6N1mmRUES9Cjp1Op4y9uPI52+VrMClAfKS/+HVLTD4YjF1vBnrLyY3yZ6X29p/m/vbYRrvyPt/plhAkn2excjo0jv0rTB2wcqjyXmvc4Lj31pLSp59vtGEyVU1WZEAqovuMICgrhxp+dlY4Fw19lM3D1JWYUC5MOGb3BhN0G5P8t5hPy803RhwWCgY+c+ysLsCfhazeTi0OG1SJ7YXrg224jlitoIcxMxRGJCH8eV3Ui2KNGGnqiPUBPyYMZ/2ABxat21apPYbwoZWGr+arfJF3BTQnB+s/DFEQJ4iqCYVMQ+pNvamzmmpFeqIT/IHqcoDPOvm1hEHfBtUSQT3DgV6t4kwWy3t31CKmA2wL2nqisqIo8OaUm6/9nHUuqz31p2go55WClbL1ozTdE8DA9Mjcs0kzV12tbM0uJnmFWYBvegE2KxI1VMhj6dKobBtxi4KyH05u+Mk/xXgL+lffy+LzkzIlM4X+M/L7lyGvuIsY3Ve2tAHsy3RAdDsYBK8ovuOlzMpnt+LpQ+6pqx7L8EUJEAtPA04N4s9k58ZNCa0NSUxEoo25I6VyFN1Nn/U7th/hfGaCcyuaI7B72tVjGijbHexwssTrVKdb0MRC"
`endif