// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EdjzHcaDwZPXgmebbXQmQwwhFGQRh7MZRnRoiUI8I6UhmINWO4vY6LpyIdJt
0cMLmcud6gdZOX67+eRI9XSUo5MK5FIKn6zCCfcDpXfk1ZWHJK5h1hSmKx3a
oLXfIq8FSWk72fuk0AB0+HHl7T7ZlNl0uxfuPNecnD7ysEV74UulxM4+b/kl
fO3mp0zKT+JQvAijwAKHIKwp0DEd/UWLlx95Snl7FrieF8VkE63dcafSpXjJ
ZljgTKTNmm45bkjuHCim6RjTNsHfEZddYJowelOQ0K8sq4o55FyIyLRmu7Kf
DfBf2Qa0nJLQP1CzjzHTVFhzh2PSnPnMxKVxlas1Cg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jeKZKTMIhJPZx9lJwacSng4BtNDs39qlY5YjLubDtwyuspVuxCTRQEGbgHhO
A6gf4RNr6eJyE/QHW8An73VYZbjapN20G1mxK9CDKcLnGYYqNVjKxW+nQZVF
VUKyiUFX+KoTKVLYAxy9PByjPE1+0GNqWY8ZqqKGauyVxmFOdkQFPeAwoPtG
NaFhEHQABLQERHHpRigJ8lxGFvxCLYtFimjfc1ZzcEtxdPBaH8sJ7/vno/Ws
zXBJqWVzXYWSFm/qFtqUSbArGKE+n+lvFetiif5bYjmsY4zNRsq+wIYj7Sr/
ziQuhZEw3LLAzFl09ya4S1NMExd2iEKPXI8AQapEiQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YAVeojCBQlLwlG/ODB80RwWGq5IovnCBaOoQU+xOH+n/okT0HLYOwVjnlzRE
XVToIcQCERm89319L7+NtkozaEkzpVnCMIHSTqT4VBLDsigWrDYmfIbVl+0r
nkCwnyNOFbJeg0Cl4ZJqeafaHKyaA3DUEdaC/88OQ3QRnufsH561bCQMgmtS
4Bgc0npMNGO2X2JMuLxECU3ak/xab+3Bq86pk//74Hq09evOlXMqe+yCwFPv
p4oyOoBwHI5XhtJXxjlOOkxNPFmy1alqFN55/UZajcpyDhuWuRvRJhBcg/As
tcZCuWOpCShc3LZGlqJ/H7+DpzJjk4tGoLiTevdURg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iG5G8d0G9Bbok8hFF0NEzgtm+Wy7CrZw1yUtMfVjop8lwECPWzf7uLjEszQv
VyhnbxZPI7xFTxIDAmWmfKNxk0SC3EDGUJMtFUP3CUicVIQ7rCLIeKcpcPlf
HMNkDJqpDaVM+5Do0z45lxhjvAj2DCBVJofV38obecG52gS5lqSzRBUCIYMn
n3GmUJkvfIfwjvKCgESqc4sHEBmvas3w01sTfnAOhqp19xi8d/YHw1rYroho
0oWz8xkRKRNogbFtGMQadWs0YX9Am/n6FKfDLL+D0klW9vRlPda/FXzPloQl
YdLu/8zfWu+apk25ZkD9aYdcq2HoSVxBRNqoj+RghA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aHBW4zH/kQd8CAuBk9sZG33eGhUS4ed7cNSSA3zboExTjNKlae0+4ZiLN+G9
0wrEFvB2B6cFOLdibGQSex/vKhLeURgYtQM66tPPFNrmOaQiPXvwmSN1Mt56
BA5rtOwtSovvHD7+7kgmAoXTsQ/ZKeUD8caQTmq2+Hq+1LqNl9Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uZJkNfr2XmW1zIwHIhpRS77JA+C/yZnKrNr56/Ofr6SrcoWnZoTPyC0h7/lR
dAagqpf5hTNy+64rlXGNsJTaamLy3B8LAoIua6jOeLVtT+UhKST6eVoYypjp
fPEI61c152P6fPQXBIH9tRCNoE3PXx4m8Cd1tBA6deV7N5gvLo83pUvlxtAu
g1QqB9YAqektFg2Zx4iUI5ZBxX/9HU4UTJV9gmkTB5/YmGlvQ64PNKfYAqXC
1eDOtCLvIDda4R7esxZ2ReAABrtCROSlIw1UX9lmVcfOPDYbJ2tLC5M6jlzh
5G8IFRibuy1opJawU48JtprW2cFQnNWl3ek3idQCzrYPc++ZPaU7UXFx4P9N
cna5qzN+2MXaJxeE2L2hptwYTrHdyPjwUPlmqi+mwChDZyHJJtBQelYwvhbS
yDecTkoI0UeyWlIkowi/mqnJoqnDnjS7shMasrZTMPuzg4xCA+uLnts7EJ/j
Rd7Si/cf8pKzvgx5js8MMQr/KUH1xqWD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
suqBgwuXyO5SC7/tR57+CzgKRO9PhrRciRSRCdV1DwiuoyjBwo9qeMajQHyO
87wLnltqtlWnrqjyKJkJ//UvWPmufHIwPZWRvxCNvR48YJoO3K7bX5EqRYjE
BhmcjI2bOirZSQ/E+zM+5CBFaeJ1/B7yBT6Gzak1VFbzaSbkGxE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TZSYeHsJklcucXRG87FEuH0bWf2RM7LrR06AUpHhIBmL4EWYiWSiwnZoq8H3
WcLy3rGYlZpNNFsPEhT1PV0Bvm+Ka13dltqxytVGT0tv+Kyk3twodx7iCEzo
hvdfgJU541gKEeI/nZ7skQk+20eA0qBRCVtpYVRxQJDYAhu6kNo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
jRz9pJq6T4LZJp0YKjRn/EG1F/o5h1QgbDNnZ9z8ds8TzTDuOwO1GxaRfafX
QrENx0moV4y9JaX355K65TxGiORjvyHp7hIgHr/yfWiGdVLVBk0iWjLUBGFm
lWoqKNgnDAyevXSx5+iW9+ghaHZ40UASSkdjicNyZD3mzG/zp4KSei4zNasB
n0JISws8m+punwYzyd4sDEpfBfvlaZihE6hJ04gATwf98s2XfRnVSZm9RAa8
E010DIZjAsXzX4Wm2UG5uGX3jWo4JThvhB49QXtKx2AogYPpGK6KZvP2Mfap
jomW4bn2REbgfC7mchwvTFMhz3l0NJEUMdInzyl/VuZTgGxfbRc8ZvZKBJE+
Ghy7oDQhM1i1l5DMwEI4XjooqomKcvoe7TY5X1ROWxP46WUkjPGia5/6fjC0
3RWmfeoaDLEFcRrXDvcl3cKXd/LcDA1q0I+wxE9PhVkvAqMUbykcMtzCMAKs
NLHNR6kIVPJNv4rgJM5cJTifi3K2HSiMIhdacQiXhHTkpJ8luq/z6ZpIs9Qb
jPqKPeO70JHT9oxlOwtgiNyxigD0sLmB4vBRVFd3K8ehWoK8shmelmlNLSAd
w0WXI/AEkdMcNXeo72+ujZsEY9XBDIWPibQd0D8Ent9ySSNGLd4aQ5ujRfyj
C6WWtbZwrLiVyYPuze1qgwwp5MHUbQywia7V+mNfFITsQtW0oZ7bSpYgjLZC
Bqd4ISUEis4iwh/IjLbZIDVikl/6JhVtb66i5vz9ORdyjmJaIK1tMEBcpt1O
jfMGzUG40RZ0J5gS6GfCl7XKRN59We0dWOJgTU40LNroaCY4NlEBV+L/Za+T
Po+9LGyy3ko1wVmHxLdZmBkbdQusvjaFQOgufuR/qCWSP0404IAze4mUdtki
C3V/8dPadK6qwrk7vgvgj2XT14T3JvVaqZLx6wqifBp7KAhsdg9VrhPeKnbT
5QLU7H/br2el/QkxXTD2awUXDPe7dAJT6skzANdJUewnkyR3OvzJUtevyzO4
1d6wWDUvv3pKmKn0CtarWAC/IvSFL7cZVLRIKzOp/PSqtQcjrYhQyqs+Pnki
DrNVOXqu/RdWctA8Qbc6bQSVoq/p3b604jhZfK3svc5pw6wcPmlpjQdThCey
5pW/hdBgQChWXBLITtxrIb6S+C/QXzHqkN14NI2tdQVhlOT8XTS6iKknaOxV
WIaB1WOgHz03nAFAXlm8wsSOgFo1lTs3SIcYDH3EoR7fpfPaCH40LevzvgEx
YaM0wJuZH3hxHK1F+rSEQTgZTxJJQ2KgtYpBLf81ZfUVsae3kXv33LHDhEZU
ErxDg2++8TWlbQyq+6SNyp2aiVMm9HSPjizqM2VAFZdtKTHn9b6evpjZOjQu
aMVJ7xc6WDHE3htHn8iJtlM1j4ISodkeiHiL0Mw07+nPdX1bsv4KOsq9m/pZ
0AkxRk99rX3GrRWVAu+ilfCCQzbl+q4TdCvaHOEzgQgbE38U679zS6LzOhMx
hZhNKYKiXl6WIdmHxa9k11UxWo4sVU9kxz7RVZu2v+ZT+EFU4m3XdW+MSRYL
SILl80lGNEXHGMBhBO8MWIoeyoJ8ceqfyQRKhYcL8HxeV4QxK0fKmSHWrmbZ
CNvgLurJhqao360Zg7ZbbrBXRbiTXa7NxXU6i9Lry0Vy1lhdeMZHPMtJCvPW
B351+f0hnZ+53xG9T8zOgdiNQQQ=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqetkdApfPNZzWsIoGG8CsJDYVj2ZxkrmwyqXYBpmmmNeDopHF5i0w3h2NRGqVH7gdYe/M5TIfDEeFFOTKpDKAPqgwbuuXlR7xPpBxvZaJTI8inGjE1qySMaPNMeGAxdTFrOZWOl4FSEVr8SwrhBEky8+hbbU0ZTigKQnpofsYNIdQpV4GyXdAXvjNZh6PvYCk6/UtKjvfEqJF7d+v0wsyflTRRajRMTcXzL6vt0vnSgWOvJXXXDd6ZAYgpSWQSXRor8EgIsnAgwHlKCcwAy6UkXg3X4P4Fs6xTsATd/xb+zcD2guWP7io4mwGf++TBR5VeLErhRXqEX6hwDoGmT9QUV6dbmBkI8mXHMj9ok09KtL43iDazhfzsghENAYI8mEfhaM1CCr2d/tnCZlisrprjG7sf6P3Gz7KBPFIAADZfBAUMTACeuhB7Y25KJkyE95NDkr873ecybBCrKkGJWRlMrY+tm/aIC+RxgUhW2QvQBPnYAJiUoRql1GAAdURc+o5V2nfapbL1HnQuTGJqsrrCnophZBQglundXM7Zyleql7r+MG/eGkejwnMymidlOyjdy5bSqMNULlCsAj6KVzkK9jQ6KVGPdKEh2kGdDjmp5rX90yE1ocww6zCT4KCuh5z+L0/AQxjx52mkOTY0NBoIxU61DPr7QCYX32GjjT3P3ykNZGLlGEue7RUBmHweI4Dr4dttpxJc7E7aR9+clBhoyVu4Y8v5kWj/XDv1wqwyAVUaki5622/O5XmKko4eS0YVJdGiFtnbPXxkyxkS5Biam"
`endif