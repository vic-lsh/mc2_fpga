// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hP2exfDz3Px2439zNMIIE/rYKmfwxTekftR0znuWs0Gd0JLigMg11sJgKw00
Pj8/mMv5wBhtapmSPVrYufGG17ZqoH+pUP2aoOARxNLXjmFuEy47CKY4i5Y8
rRSDx1tBgmAXbtzIdUF4BokynkIFGY/x8er/oWkwgOwkoIVyOsf+DCoZI581
ETW/W0k9H0CyrR4J6afABRZaxGredthAxZLxfk9AnUpUJRuPS1pcuTq4X+J9
HpNgZ/6Y+fhF8mxQNek4XEfFRIlvLqn7wVQhFRk43ToQ6UXZd+VZ5h7uoZMw
rFFOG4+swNaRf7qBE9aS3orAkU/16Y08kc7RGsi4JA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m9+D0irE5s8mN+SAo1wtrs4yuU+MTgzDhjCqvUST50c2JFqnn5UNFwTrYPME
le4pa6Npi0XWpa4GZ9TOdTtB9i0dB6CKUqFiJy3eYeljjrNZ1PQjLyYEk98m
IPgaQD6TgnaH9vaYIgnLgdrj+y64T3R2DMwZpaMDP8Z+TMrZsA5oDKnFpsZC
k8O7j4+DVnsi40E99cv0jmkNID9isbmTzCyyjVabJwABxTjl8Kstv9WlLyKW
ICEl9J++RdaIOK5Rt21vWe0pb4HzqYWCeimkVwGcvjID1ONiYa1Q/XZXBmos
QQ24sSAPjyZD7HUjsHKSoD8QTqP8VdaGHwOnxwfMtA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l8ThfE9DiDb8+3ooWcRFnwCQxlGPx12m9UIkh259P7ZG6KiLOLfEAspxmglu
D/jWQ4heKhcKr/xkksXiA8d2ytOXKMg3gBSYV0rn1goqxXMhF+YuiFo8sOKQ
SAEYsz9kfigIYG/WC6d7VJCF8nJ1jlq8ccBkEeSLNQxRMLonSng0WmNceneC
mA9kPXVXdueO/PRtdiHiiqsR+g+GaatebIOU8AfQj/UYq8FIWzTmS/Bd5M/u
DNKyHwL1nF/6KDxB8Rgem+hptxfq/IW85EDBukC1IztEwX3lRTphMSTgxlCb
/D4u9vl1Z+w2CUlV/UEscMo8NNjDRAcGCDqttg/YGA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UJelTVApGltOWskyDdRz5abxUfKMpR5FcfghXItayQ5JOZpLhgOGkPuvFMvP
lpXvNQ39Os+FVx7/TDNfuUmSEqV0tTvAZFs7bDEdUK/guf1jKmPooQMUXGAn
ZixdQjUrUKlkouRgbrlYahKHGnmQ8oyOBWmUpko23c2LaIrBNaoX/LGXkQCG
qc2p6EjGLu/zH2spHr2//gelXqhKj+/iszRSB10S8OlAkQjriicaMZHKzIwL
g7uc1T9FItq5mzGhw2lbvztAAu4Sx/QlmCJ212HISFeD4bohXjZ6+zKmKgWh
1dCRWkwJ0CtEeBYlyHQn5F4P84i1bWkhCJoXP5STxQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
galSGQZJmlMs4eF4vfnVU3nkoe9AsVbhHpdJfyfrFIyaaVdU5EUE6En4/RpM
5tHqRy4Ba2sbplzRw8UPvym6sG2talxtp3rZvi7BnASK0CnwQlYDJu/UKl1y
czYPq2J31Bey3aS9YY6adinn315Si95rYRNu//SGw6rvbSitjGw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VMOmlgRlXafBdg6iu8KSvW3sDdfQTRi0fiNLlTz/3OojyZ+0RxdMN2fBgSSZ
gceIm1UqFLVF8tJXR6AzDN36NavZWgLUucPsb7YaUEfe7Nh+QABTlZZBI0Fg
GbaDSnNKh9RuOCA6BTtb3ng9EPVE9zo22VM+riUvLXcJGOCvnQJ5dNTe5yWc
tNOT6cTa9Xs4wumKDFFttsFmPj3W8SVY7QclygYQ7MqPgKMK8r43lWs6STOL
+1M6081nREUn3QhrFSiK+xmX8LIipHXOocJ7jkvNJ2QqGEBcyZ2zRsr6i/CN
MSh7X7+QIZy5gehz1cFv1ymHqMk7hRd8Ii8FQ334ApEn+h4zA7xHfG9JciKZ
mLksYFnULbUo/6n3ErX12pgfz+3zccd0l2lAJTl/htQ1t68uN++HonOdriuO
eAv/vCk6R8XTmBKW75ie9QtgVqyZXDc+50oxVc+BZE7Ca127Gu8LbxdK6Ajt
upK8wcrrXjKVNdrdxJxOoPcA8X8JSLNv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d5dSGqjiY/YysQ/eC9YGiJpSesFDi/CZyqpHawKV8WV4Z7G4neA3q3Bh3xHZ
sJ/S2krXwsNly+d58CcieFxPDPofhbD6WOJKdh26cOY51w3zRYqCMLkuF8OW
DnBojdc9xcWTP7FBDTxEA83x1sjxk6pqqbd9hSiKaoXPOoPSVVs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Vzh/+v4lZbHDeSRbeo8Erex7kPPvGw68IEa9HCEJHDAFjmSKP3TnRX5W4xfI
VuscXCYMNMu3w5mC7IR/jd0D3xQirwpYOPzeO/j/nK4slTxSR20PMyMwKw0+
wTn5r74m+8P43Qs1byeHOIaBR1nMGqMu64eXbCeG8u2Tx8vmAYw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8880)
`pragma protect data_block
kog/7EpfOMGH00ujDMyvIAn3eZNC9nTPi7FtTpPGf/sdS8UYC48khoxYaA3d
xD2IqyppUfB8A4pd6BFEK412e27W6KlUDXimgdQLWGlwH42T/D/Hn3xt+4kg
eqcMaWB1YeDJ6tJ3+GgO3ZAxCXoxkjEPWt6mL0doZozKHS9VkfP2YxBfrFBd
zhdzHs8Xtd1By7LBLMttH1GFCsIXfm2fX2zCw98/O+jQ7uEOzyqn9UV3wy/m
SyqNW6sZE35I7nD4qKuWb6UPA2sPHETsQg8C00LY/aXRiT6UkHl7+2iitklA
VrVhHG61cIMW8Pc51bXbeB+Mkdg19qEAnTOAiMOOXdP/EH25JyOjQbYV2gj5
NONypuKiMkLZCE9S7IFk6sIvYhJxVpQ3fHyWfRcF111HHfsHQiGNMJhZuny0
laAz3AmNmUPodcMTseF0kIw1kR671DB772MLhyEy8YK5runZ3FqeVMtVbhzm
WKb8Y3c/7txo8rpehuHRslMCaQBs+cNBNJANMdVtMsJsEOt5e8we575eUP9j
DM0T4FwIENfa9MbpMrHfiJh7hb6+I3Zj1JrcGENu5OYbsTvQBk2cMkoWmv8t
aoCIfshc60FAtXu4qQTAh0Lyt9NS7dDI72+hgepbzs1WXRkTDhlIzQ6iK6Mo
3IobR7VV2lXbEEm0guukCOSdplJaGQUA9MSawd31v+hMKJ5GXU7IyElwJxqg
h14XuTxOZseDZUR/ZCoBKuDVwCkwOBZHpZEc3Wpa57i81LffZsFSr3iarqQA
SbjMR2YO9b1fGc/NH0h9M2pL/6JWRGnUC265YoyaiIqqCUGPA2WYftmAFa+u
Y6zipjzGO65w6E9TxoLxfZ45Fvx/fx2iSq3j2HztaP7mMxzypp6MHMlnL6tN
vusZRM007kdu4tC0Q1/ugVoNB3wEjhdyqQHRKM9E7lQbXzWruMA7mh8Ollm+
27VCSnXzQPgXA/l1onuXyhzWjHUBmoVfDdW5b7MYp6ngbQ9WqLgUIhEwmfNy
JUY9W7SN4tX5v/h1QSCS9mEB9yTonwmF9Xq/401GeDSoERoKCIx96aZA2pWL
q8dP/NOXX55WoPVaEW3N6fYj/q7F0S3C1U8mk4iaaXAACgmpHfToV20b7sqH
lni9X0ZV86RHKSwSheyCqkd73rvQ5dnkDBRySeT8rwLQ0P2MoQpuNuswtV9U
B2D0d4jjH47hwx7xRPNpUEozHt2QLadcaHc6nRWR9+lLq58avDTCrqkmAqea
xFPFgqYrjOox2VunUlEUMNgpQQOWxM4OGn4jDK4i0tWXeU+HPBsq60+kZxXI
nRF/ST3OA3G9yRjlnfmYiPGeaVYQAkBgVz4+314Dx6GjsQ2qOWwtmh/mkADQ
INqzQKlTSp73OGpDcxsmdGolZL439l3dXBmvOcUjq1TN6F/6HqKSY5Ou+hlu
r/XqpQ7fZf2YCzdtZHscxWwL5P/IYkSjIDe3wKPOtM0CbOQFMVjHgDJ5/sYH
jQbGAhmkmkMgrQpWIzrqGiNn6v+dAwpYbGz3gR6leCJmLhEX4J2NYOJeE1kd
46ooFQ4PqYfJ2GY9ui3RogRtGae36YXL7H9rC0FDPMqZX2LcJ2zFsNiKiB+b
xkZGkYljdBxVkJ/KqaNwfvwnxlUS/2eYY8MQUHjZQZvi9uaYQMMF2enM6giS
UOfQ+UZSdm8482xhjfeCf1vD3hV4FoKfypNMZrTP7CHErmMWIEqCIQixgXWu
2PHliVk+1LCLtOBe+WLU5jZDsB5YnmJ6ORchSDoDVbzvMgApri+6OJO0fN7S
Byn+XlRtQmvOmee+9yz6ZSGREo6UkQdA5BUYguFJbhQVIZKwVn39q0Mz5fY+
bFTJ4FmZ4e6YFqtdMA54aBTEo1+VVx2TjeygmeYCHW5OoZdQaYIFLi9OjfMJ
0uY1u4uCAp3b48MLw6PbhVDbB/U4DLXGNRl9Wc946RrBFEbHgwcqJ/MMicVK
CCQJkogF93gcVlRUP+Mnt4lW9IeMWZPkh6GROLTA4I5S2xx2WaycEL7+6S29
Q21YVXrgowVDdWUfCeZI3gEU4Q9+agZOGlzd1t2BDpNIk+NSx4nmm2O6cnp2
k5u2Xl/xXT9FlX7PvocwkyRG1YNbRnKrX1bsUElCyzbG3iHDjnxGhZSFtOE+
IAceI1bMKYjxBK38FVdl8r4SoxlDQwrr5GeSz079esAXjNGFk3hyIoQ/XpgG
PNfOphRncowASoRIlsYx+Wd/+0i7QN4dsGrNiDAxaClZQSQbzGmJ3DRLvqFm
dLsIZNcURCL/mREa7VAP0XHw1/MJicT0DYqT1vL72fOxLYuevcMdvXffNdkk
xa5o89t/2yytlfxOwJv8inK2I3Dep04h9HAr3HIZ33CsPRoPgO/0tAVLEqmU
ehVavA1cneE3AcbMB9RLQuDQ0Ym/GJPco+z5qTkIEZgBbEWmUCfkwFLyka15
2JKUQDsR/hzk5oOcox8sogp8HKsnG1a442bOqWPYR8ZSJZ0lGcXQwjf/L0eT
4HwhN4WfMwfmjTDRVkcvJfUmESGJA4JsZOXyRvw7No16m4+ARcvGXo9axLVI
grV/NBCAzSTalXjYqoekPTBnZ21x2ZUiSFksg3q212LHbOdil9Z73A7KW0G3
mpPj87BqANNTOJJ35+B8KtMZahPWhErY60obmGW0/U7w2lt/QWbCnqdlxJQO
EqfBQUJbwS3a0S1xOm1lfQkE4dTZADWGvMiMzsY/7WAP0X7uO9Jahe7MVANy
qkd6V+QyLtJq7KctU7KNPQ60ifPtI0cXe/DEsk1MH+O2EJgeEKQuUQC4iC0N
5XfmaJpnupCmA2ViAQfE9RyW2YAwZYzwRjBTQZ6zL9l0sGpQ/ff2RoMnxgL2
my394DEZKvhxLyJscCK/630LTOaGvf+2jjMsNmkFtcCenNqE7haI119RpoiG
XsYXeJk+iWm+VRKIHbQw/2/IJtMsH6APJYq0RqlzNjlSkJaXdp1LC6NhUz3m
SbxOOFbSOq5gM605XsqSq/TDRtrpMWL+C3sjlsby6quBUHGHG0sLWTE0qdkM
EI7C1o377RYNz8nBKnXPYP0Ap9rq4TWXgbmDh5sKc7DQOhBuiQd6tP+W3cMP
UbPSasOEMjebBWwlBby7eDhQIJzicSZ6XQMvRWiiZCz3emc53Ocl584zXso9
eDQ0r0ysSNUG2YDXspkRUTsIG70NBaezi3puWSt2wj6NWagsfpaW1i6QYooF
Xsi36UYIE0l6XTyZ58vXwLMwJ6Yla0jjnuyQ24uHpSbec0LIVXh5Rmn7fvIR
rC0Mk4RpuK9+O8M53wkVTsMRmvNRiFpujXcTTJceUDoddBsWWITI5zb4heXZ
lhKnrEYSvWOVH7isHS/D+rh141DxsTRTLCMo+1UYBlYa8XMdm3qvs6Ct5c11
4IDwyj+Regyqlpo+hKvKo+1PKVLHNAd8X0ZM6l6xJmiqJvvhxpMA+XCzWGKV
aGodh0y8CPYmMIP8Bnx6FF4EkPIA0Oh7/0977JTq1zgq6IbapHQSPe22awbH
NOwctIjsUIWF5syQTcUXxHSmxFUn5C3Qq0HspU+7eK6DZUb9L7ScGlMcDKsy
hM9NJizVQfIlqdUHhKAVpMCGTByw+sPHAQUQtk1N61YxJTghSa4nlfrSKs4d
g/70mAEbjOnzHs8Nj+cV0Nm/0QKsQtIpvNBdhMLvBvwTBI7hkJEcIGnUfKdm
/6lBJFFveeEfQ/gqP96XOmPFr9d4ekaeHSQWpIcb4LlYtI45fKN1IeGbsQNd
n7AkEFNJURYC6vNgkAYzmkt8OY5GrnZlrLh7wlu+ECkzNJYTD1rsfycYMBnF
3ZDpCKHfa0qJKmsQK2S1R4qitAipDaeY0T869ATC9U2VO4f0eo/4D3a/Qx7t
kMI3PybFb5iZlApj3lcuAuef26D4iwBUNxjSuf9VTFhOVzfT25cpDWjpPAuq
7aS3sP5TYdcoJtDuFQlavHwzSiWb46XiZQjZ0ee7/S6DO24geenytYAHb33R
r+vG4zUhx1UuvWJxH88zhHMW8Z0QHghagmVCLJaqAybp6raw+ax00P4YjKZU
xsniSdc1TmJF1Eaaqilaf1XiLuhJDwt86lozCIOK3L5YBJMv1xnD2JMNmm12
NaA2NPL1P+FH30YO9QeRX6drjO3CrVPTpocQBpPbiHytBgsB5ES0Ur2TH0+u
sZmVkpgGvIg53MptDpIsf1BO/zwQInfUhoXvq2Ox1g5Av3h4h/J1z8Q7iwwa
FcPLt+/9AloG5CWUWSe2BmN447X4/m6p8U4pPie75Y3mXwS0niSfrEngmGDB
UtEvt6xIqAwE9dCx/yIYi+iUvnIk9wi5W4NA9vSwqMu+he7WtDJ48QkWvPHK
JtYYLmD2yEG/n5CCDTy5VVYxAsnwsGqEnry66zzLJyc2q4lMb7Vag1+YYXbI
lCryLxeAd7qp0hhsVfadZAMitqjMo/UKhnNu1gRyylFnV21n1dNwrj4dswA7
EfD//NAAT3f9wBhd7sr03hZcx0zDbBTEIf+I8A1gvEOSYfyaiN55F/SmTllS
YjTHw2vWFm3mWa1OebII+d82lDhukjAtK8hQsX6xsECijFHODsbaV5VlkdU1
k5FQ86wPd3aucGJ/vqctWNcHhsjRmSO/eUqjVTO1SoHf3Pv6Vnwd8enbXUZw
dzbo47P8wPtfmWPmieGzFhMgb7NwFPJnUnDMFGaF0CmhXMLLEGri0DuPVqlK
wxU1s9aqipwEuX6XvZbSObz6UlAxIVQvwGXmOYGReLzEcxzJrdUyWQMQCjrb
UZWXE9rCgy5C5ZKP1VoeTH5BFvPD0Q9HuKOX8Xrq5WgbciwJuW9HnKrPChDJ
V3NpSMwiJgzj16NHSHovqSTGvnK+SSOJBFZ2pp6y7X4blUZmGJcQZkUdl2aw
sbbCMDO+ewgZVYihAseNqN/6yiNFij8ywOA7E7yHo0p8YEOuQtxKdX0yvCqe
6GIbpP6nvIobLrEOS4xRBUAl83fHcZNXvIbUld1COuvGRHgn8/XgqDmTksvg
hBeobPA2KXnHSqLYVgkLQoq1acTWKz755/mH1+tmCYQYfkAV3gTAyNxYUyOj
G+GKTXSlntzvdu63Xty+26p1gPFCxGcR1MLlw1URhaNAz2BIbgnhysUMn+0g
BBi3BgAiYaH29R+ar/oZKvzWjU4kz3Z7Q8kmoOfI45hrZslSZMqNUlHciH9T
Rr9oEieJTLb/Zp0iN0LCfLohZ8ArOu5Noxw2YqNIaBVK3poWlxtGPOkWM1P1
83mQpjI2NBXDXPBluHZcawR9hkr75U8rQFmVforEYCZUhXAKqtRwT7dixhyN
QpzvwfElNsGlV+w8diFhTr5KNJMkzZDv4pikphioOjD1gVUsZVjjxrO/b6JC
upTpUFwODJNiZJ4QPchUmrHIqmh860yXQ22HH+0r/wB9EvxYY1nT0EzDG/qs
D5TDxeLaJHe6SmNJYSxdkvc3B9yDKnof+bT2cQ0iyKPYg6CrXPns5UTBQuLx
yyMow3G7qWfO4KbP2Nl4VKYynl5OAFx0waHNhG+yjneQKe2chL1zIrlo9EuL
+lSMoFzz7mPZymO5IfZQmvR6aNoTnaMyBxr7HcKNnxxz/AZ5L/8fZQjXU1Ci
4X2IO9ErkKsSTZcU8o4Ep/u15KwE7TcnDF8KaRh5eB6AWaYUjmxcn+PeMR+G
Dwyj9l7HNNTMpU52G8sZfF0JqpDhDVLx0tShxa11sKa3IRoUvT3zQdJeKEY0
Y1YAfqgQO8bcfCKxcnirRm+MCnjJG5B5Cf9/aKFQ3WJ+MRUXjvzXLoxpRn8c
4lI07Cxs+XJBBJ+rnX67MnsWGx+d2PAcJgsf3GqqZ2Rhf6FkOekKDITWGoGr
a62FB2wqWTt1SIpPdi+dkLkcw+S2lm+8LGrNC2IP5G/3gpwxeS+YgrWytyn0
OHP5Fu2ikTu/ycKwM+LrRWrMz1B4YD2Sj72ZOdvse7ZXzplLEDXTHdgflQAA
/HIuR+753RVwsEhFu8874PupNrrxvDgXPeC/Um3+VL2Vp6o77Eao6t4mrrE2
CSMA/76vdLONS2ChCJ9eMZFLMuJhBMTy8FwPuJSV5LKWLah9ixL8MDZUYXxE
MnInl2UjOOQSfUK63duYlvz9ZM9MUADLRZHenlv001AdctEPjLr17BZUkQOW
dib2Dt0mO1iNBPyVMq6vdR7RBXPjHl65H2IpYZLpDgcqQ0YgxokXOxQ9lZYm
sCBO7FfkekvGCD/CPce6diRABdxeO6M2wtaS269J8lb1Xvzeu4YOmwnDSuXk
Eh52DUQ0i/K7lsD8fVPToljpx2VPO0qVX2qCjhG2KpcYOzFiSmtaMRXtJN+D
z+ShAXsr6vNo0qR4H+t6VFCepvLlhXEu1/N0iGF92Db+JKzDElVP9kkS6RzH
K/RSp2FZhyXLzDARrzIihy8xji2e2RtBpwDlL4IoF6/Hpm+vbJotS/qJSgW8
7fvp9xAMvvFgOSbh+EHcfpQxvc/KnW6PaJ6PPhmfVtalQvJwbuDTA5W/8D+B
RuQBS6aB7SZsjgwcFON02zop4qZdX3kVzGjdqbrp0Zs0sP9UXcuu5kdk9iOn
BAK+4tis385ZqyLvxKvK+Qy63XcLXxj8NUcD867X93l0G6+bJHyU1i5y/fSZ
TlYEnY2m4ImFWcxs9uf1sHa4vAtqHVZnrjbRE9+w1jv+hIzzFX5LBX3AYZYZ
SKr53lvKCgElLEVa9c9wQFNohbqiTTJqRBOkjcFj+4NwzdRYSOAkY+EWz4Mz
jXjMeWYZwvySoWd2KfyWs79zLQy4s5jZjhf1fOWlONc5YMl2m2pVXGyBs0r4
iegG1lL7kAt9mTo1y/29gT4eW3b+sgHdM4GjUYkGq95pt5nlbGbprk1VFYq1
ayI30L5V4T7JjH29yMSsxUT7mKjBGIjmCY3bA5na8SresJpsDVKY7cC2JTsJ
G6y4l6XPm9639uVrxqnKHCrutNO1nUV+tdFJpbNF43I3jH7lmoc+xCB7wqIE
v70EFe233vJzad3CPN3R3Kjbs+9hS6rSzA5tkFykyWnoGdBIUiWIb7iGXfGQ
maICwJHsmLgwCwDHmLv5fXWb2WmvXZZgHxBI/ZOhsmabBDgy5+wcF9k9YUz4
Yclzc3EqLWDhoIT6zNhup+rw7pI/2s+NlRo6I+sgs01tWe4aMRpWwfpfb6JE
vJak7ODx3M1VVw8umaDyNfqzEEhIhLU1pt1nssJxtaBkZ2L+fM2evDLJs3mu
ByudbyYQoz0U+prND2fGpdbwhbZi5OIi9Mbybkw6y/AvMm0V5rPoGgJYEzSs
hUrLKbmAQ9R52GxRONSauIQBiOmUWSZ7zR9BJUFtrNGYqZaeE2HFCG/MBZfI
PSCni9a2esJnT5Kdc0AWrUNoeXE+t6IRhcjyg4GXcPEjNar6RnvlB2zRZUjI
RJfMvcDdBqxX4Q43LJ/jJnsDu9j77w/hdzKK1O9EJFhhrT5mWPsJAZ7UoQWR
Dq4PBWiTT8F5pdL9IJOPCUXD4yZ1h9/UHZ55u62T1QX+5Nu2ti/gC2LzpUmU
pGhFrGRinmVlC4Se3v4vsgR4HX/Sb8eWFdKGJs9vScqluicWNAQpE707Fo2h
tSCubPj6B2QUwP+s2Ghsgb3z1EPPRI9BN1D3CGFu7T0+FvJoV0CLz6xMnffh
gqlbNZbcNRViVHswxDaYKRtNc/ZJ9DMfpxd7Bk3XkMp69xVzXN7jkmRQyWTP
+kFpdsZhjSHxY6KhJL6S8oOiAlkIuqJa1i6e0HEacVoiMPIQfXN5L2cjzu+x
eFU0mwtJY4kmQcMdOS2CCu0Y+ChhukYiQXFBEZqPYoAACe2IRGROyoq4Y2ES
YV7XVFBUactIUoq9/msEflg6DvsS+9XRmNsjLR5SeWPVNM6Ys1LHLGN5Ip12
A1DnxGva4x112n1L9yIYeFHV+HPxTGpSkPp0SE71tlN7EQumIHB2qxBL5UQJ
HD1jKebTjyjUkX/q7nDRKhxeyMX3Vxo5BrKNYE1bBw7DwJXJF31xF+QScnBt
/GTR7jhlWbABsxmiT1sXrQC1vMjVDdyvWrI9tuyz+YDnapaQlcZkAnwetb+i
SeFADUJ+DT8DxeE+Sm9x/Ia8KKnbRKfrpoqpwNYrURAi5KhZEO0PCCzoVLRb
lv3abEXZT7f6dsfDsQpfzvLi2F6YYZEClR6azhH8LWqRdO5jeYUwTch68YdY
aQawk1VE/JMB0dSavtwdAX7kXh5+LVc+3s66yIOUaJecvl9eSgdY0mjHz+4M
PLALxEym4/3l/Atz2QSynkvk0TjZR5WPJJWdQ7tnTlCtqAqW2QHcWFtn94KQ
f+FAWljl2rXLgWYOBF2fqKyDZlNxLu/xGD0Bzbp3motAV6fycvrKIKCJae+e
xg9LJMR6b6USIysN0ZUE7z1snOs7g79SrxfxSMaBeOjhSXfqaAeAJSGWGI83
W7ep5aAB3H4Ju3vJL6tjfOQt/0lyvNyLpG8NANGz8fASEmCpF2E8raY/z6/e
dgr9k1aU/XURv+/uHOU0i92jAFpqJVS24eUHUp9FsAEM0lyJb+3pdRrSW+qG
7zXaHnwTjXM1MNzecRW1Ip7faZpycVf3pQ8Kg4qtmty9Z3r0zUb8SOEvUuOH
zzRWYZnZXgHeZIG7plZeMRk8Y3W3HH5KtD4Ee48VPvlME9gX0ywF2vhdBCWA
1LZK6A+f4NqTipDLrRSrYxOHujn/f7FKxVjjfC8Ax98UiRkWwDMkISvvxvqT
kNEGcyFualKuXhnkuAuO5O0MIL+iXMzejPG8j00h1SHVM6thNIPYlJP37Z9u
yU2lZvfSUwfUvGfkiuTWS7j2VndSuJbigxL5a0O40VAQreupMhvWoLk/PhC3
PUuyOC2m08A+KWn2GTEnoYXgBxFFBvgxeKak1mS0vZRfuSLQiikiYmIc0ryf
n/uSQbi3yJPtt/hJISjBMBMT/03mjlFDqJF5sXCDx6FPyMHYazgIaZzZ40Hv
f9TYYVlLfQASBzhMGXXbNW09nFakeESl6nEqrdJDhoCKgATZpNBZScdKgils
tQVh8S2h2dq7I6hFk0d1X51Fy8DGf0ZnsHJAEh0MEpUkv/i7LvqtLtFsirxf
jKGdHIEODhCAuEXcWcXfolYGesjPzMJVeUhjRqWxqSso17dAQXiyFw4moJa4
04Gw3f86EIhsu4n/h+JLLBck3WYVu6pNazWmZXY2thoEWGI+MsoPUOZjxF+m
+3tREI9J9yTND/z2Oj1GeHDSmdf2IMz7Mjv2n+ba/c8gZKQVdKasZRzz7BWi
sZMRbnl26XVLx1JMgvA4EXCUnCG6gq+fo7Ird2nahySV8XA2yWqeAzJ3Zro7
u86hUQCdp+c9mpDPOkqjO1KFGUY7qSkfwDwwqcB99fQX9vCISg2pL0pBPEXD
EIeP58VK0cr2EtS+1oiOsKSy7ZearLsjpNoHGwYF3ubkmEYZwLpC6sViJP+B
HN1xc/Qn2v4YhielUC55TkNcUUB3NcKJnr3QFgn1vNbEiOr0ffTfANcxBMn3
pF+X4Byar9Hetzuz2bP/C9liGVcfUpilXxA2knEWhz7+SfEsAcWNq73arNV4
nblqwXAJaCO1GGMYIxhhRqljpnAd0mStQNdF/xVOsMDODNwu1GZuR53GKS18
xDzjO2zxlfhrISw9KHwT5lVSpHvWavlNyQfZyXyPlInrIkIsPMsU7xj7yMmc
xSpXOTQmmPSdHFpTfEAl5jJZHLUrghHZZB6MZEJpZF7RhUgtru+HBYgx7z4s
xdBw4mmUPJn4yzdao+eNGNxYJjAht2E1FH4iWv9LbaOA9dV++ASNXhMsaoYd
cXOoSoML53nJ1fUXWQ1zsM9zUfwl+yHFYHqx5CBzgVOceFny7YZ8tTqPk4S/
25risHdQPklJYVcNW7xKdZoZhtBab7NAnFmC+FoWcV6+e1SWUVZjw0pt4P9o
KW2kC1MeP4J5Y6EiZh/BLZ6kY2htW7P9nLWXOgC2Os/8stNVqArWIMN2O8Tn
ttFuLaAnLeJPfIUMf1IRJbL6acsc28/qg/GZIi9ImwslhE+2L9tz5h5gi+Me
C3QfEDJEeND6mmZU9JOL3m7WDfdqYpz18ZfFt3nt0Rh59X5eWK/+km+d22Ii
Ubolx6UgdEQv+SbvYnhrSmQ/F/4mEiuQUA+sfw2222G9WILksms2GGFpvEDo
kAa/vrwz+Yhr/GE19SDSAt8SmDSGB+iVrk3CgYCoY+gKjLtEQXB/ILuuw6QT
R4OzzNE8IAUAgw4ErmuVThaWf11vTHwKFWzBNEvSSyHHBP+7q2dPIpKeT861
H0xYoNYvOeeU1pJFfTEdbfGDrk2XBoG6whKyyd+fRA19HkuMISp3RyXiysJY
y/57tiecuzr3X9NHz6p9JQoMYQBRIX2Y/6oySEzP1lHTTaEntElmE/5+IXdf
rBkwS1xPDc6AIPeV/bdW6TjB25RusCbED6LCAMQW1+pVOhZPapo8uQ5agkr0
xrC5jCQ+ZjCocM2woVAsWn6C0028hL9BBfvt0eKecySKgTOwotequA/d93XD
w+m11BzIlHVUv9nkcEP1j61kNtXfqFOpm5A0bF1KNR+bb+QaPwNMUGQyNalt
/fwsu4m2DPTphyY4c55AStZyzaSPDENTwa9aqw60rHRFqxkVftat2fNJtI9g
GULKvtnu5cceraKIIWJZ1ukbG5l1urxCy/IF8PB6lJfOYKJd1/3uKhq1LOPI
ty42I2uD7kWGxAfvVxpVOpo3QBHsbmR+seAscbfiLw+4TXlwFABMIUCWoT8N
hxtwtb6bsh7iShIZVF5nSTNzP09h6TeFO/SAEsN8nn2W0HWlC7UMxHCHGWVX
A8XBI6aIYaoVCtKSImL7VkTeg4uc8pxE5Y5yCOLdjnoeR1c9u0xD8a03AZE/
kIGQnRZvwHG1RochNjxYaD/CCQ0cR8JIz8qCzhkeXPpytMxU/71J01lJI/V0
pvGVRATlSvCJ/CsEkfvzuslBogj5+vul2zEN8axMQuAFxHllaAfQth9ozaRM
zfQ9qA9craAjy7kWAwfV0McyFzlqf6rYBMn3I/v+5WLyzN4AF4wGf2xslad2
1gH7s3uzkH1WayJZR94FZVOdq4NW6zwevKZdRnormVbvRDX8r+6UBX2nJsn0
ezVDMNKNKp3ycKhp/dLQmNqIGC1JjAsmHrjRZfQ3/hkt/l5lf07zKysHP0tE
syQX421YfwFv/9qe50ESMyMR1EdGfauITddVssaSeSwV9HagcSEzenugl4SH
Y5puwWWWYsrGS5eWzUOaezGhF1X6JCmqHR6Grvb5qqDBNH/NQ4mbW4xCTaTW
7WAUCJ4S9q126i38jucNP1QamzhGjoR26O/bjcnrD/cmA5tp9MTY98BkMiD4
DgfnWkPLuaeh0UmmnF8nmwhE53NRPfVnkRmfLUQgAHOkevlLq0khI9ToQUIq
/CCcijLcN2nD5XpyJs646YNi8A05NJIaXFDdxi1jE+9JQGc49uxz8M4AIFNc
CcQm3xfJkseqRkUtHA+txOV6pX0iVy/3tnmeim97wWLRc8Z3H30guLmjs6QT
W/Jsal6EaEdHxhXOKvKp8w4PcOqxT4D7yyrlVqmtz7gdP8uCYu0jD5wQsaHD
0hrJjrGd2pgM+SJhNMo+gA+GJ0VD/pZsfttThoUY0eIKXfbSdHBiuGWSt60y
hOHjiwEOWq+Ur+7bCuMjY5gaBwFWDwPkyluVUVtwezo66HpfK9B3BUKDzSi+
m4/G/VDO5WeXsxwpuxqi2wkPJlxKkG92yJXMXmmA9/L30VxjBVj6WQS3OXtH
atQA7FTnmA2mjZ/THYxV

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EzCD6YcoVTu6hvlb5+rrI9ZnPkjWU8K0YCnIYRYiEL2ZtMFvMYDj6sBgzZCRzFdh/0oYbtZ+GHnaHxhnXEoFUXOMDY7kI8nGwgOdv9Hy6r5NEHa1Q3QzxTObWhp1oGX7zwz1liAnonxS5MJgXc3HhMocmBROrTED1pBa0gTNPlKrOuUwa+DXri0sk9ou5ynJzxY+FXikPGwLC1kyNDKoDtx4OX+mdDktOxpURMDjXOdMfWKJh9I5ZvU0LrMvPcuT8OWtCdQlXuwIK5FsKfG2uh8yL4i5H4ibIdkhr4FxSzrZgfmz8yoBxVgBFahuFLp/5LFhKE7QfjDspQ9Z9ofFUHcux9BRZRXAuUQqbSD7af4SFLHQQQMGNf9bMuL7Oj+Jm2OgrGAfuST2QLus3qvCiR37gFglw0SVTLz5qx9Q9QiERPxCoX4f7ucsRrZ/NF5jNZgtXjS37HwtqAtMiqgRlV8JOMYz1TY7eL0dSTTDc95dI2ktBRnfrq8VBKd97gpgA0NBbB4E5x6EHU7+/AawFDJMiq+hoiwF2PcEpbtb8zsQ59OxuORTstZNy+V4gm/MaDq1VUXZrdISUiJY4YpShutSAY+QZNNyoo+Fq9oYflG54T7riSAlGAjfkDva5EnkSTOnMHaSBB5qzCU+fYEfgngmPSvBzXm6GHQyU2TGYUS8e14IvOyKTURVN4o5gRa6XMXqE3IgcnTau1h21DHqaXXw0yBgNz53yC7CiDZGMyx0aD/R7edKm6hAICV6/TjhAcjjmIbiLaOGT4B6c1+P2T0"
`endif