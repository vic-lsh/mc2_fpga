// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NdA+4fpx6uZOL0ZtuNKcH3weVnr6xZu/S17acUf549gik4HZndP7XCceOB0v
yqUkVfGdT+ddpI5kND1t25IZfsdbI4Rtzsou/3rBEEKxy497xfhCKIVgwzmQ
ogQoj6tYa7y5LrxJWb0UOm7TPI4tZW9jDrxuC6jZ97KEC+rKXRPbKitDC/UP
Kl4g0e5YeDilLvbSJ0iSrJ4zsdvfPmxFO/fUv9kQLajpp0IsW16IeY3vrtbJ
0NtfWJnWE4GyoAUhfDnQMFmrteVvr8bkr6kSzWz8mW8AwmOdvi8MeRD2zQop
mn3n1VneACcwZBCoFaXs2LgmlxJ0fQCjrU0UY+8T8g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
htFKPyPMXpdXzZbEV0zwReMABlqLX85lOch4WHyeJV4l+pN13AQLwfRg/2Lt
aiwI5PN/PPkzninhaoV3rpHN+ojAGMkJ2klcuYWxEJUUEmxZs8BJWaYjlYGH
kT6uDXpAtNkZFN1zUYggWPsgFeWsyr2V0oEsx5Kx89xI4kItoKKEeaSGh/WV
07BfTF4/OiyDS0YC+Lvu3r7O3vVbhQlR1J7YiMeA1m/IRNH/oQgSg4Pv/C7T
NJEHfinlj3XgfI6rwol91sVseIxcx09rghhcbamk2P2E3lURoZ1RkwM23//J
6kmJ+9JWPQLNBVC42/HoM1wyMY0svaezf6P6lRGcmQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SlwRWonVOv1ayDLDUsHF1su23GTx+BtJxbvGDDu2MS/7O/9lhyHMferJcG4f
oh0k6q5cGXamTqKHYEPmlPS4EDUNWNZV3f671ETlil0rilSBZKvohSEVYVH5
VBm4Ft07JS13Ny/LmhvL44Ewzc0eA4MbD236QbfLo8dbJvFRbbaWhv3Us/H+
uoIXAcr5PPbwfOO9p8blx6pe8sG9/nNiPVhuDYh9/yd3cDh0LgjqHb0esgH7
Yj/1tue7YhnyJ6eAw1Ag+a0jlrjkUMTitCOU5Buo3Jdt8oExpA5OTiqMLhUd
hWYoRcrZeura3mDF/I8rIZGyByMsdWqXm/vpWGzzCw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
evgNPTuba7ugtQOGDIwj70SMKoRNwYKbqr4h8vGmNtBa9Cfcs4Z0JxNPQyQO
jkzeeue650JBFGazdcYVuQun/wZnENsRBUlzmf7PlLbmvOEJwHe4UUA5tU0v
i0T7LPNmQsJiHCPFJ4jAPQ8EAQFrSK56oNIA+ohri/m91dT8mRQ+m2L/sRJz
4D6bTmy+qupNL95yTYIqUck7Ynp8i2ooauTUfi+KjIU5d5fU137b4+S087Tc
02zdlOuUBYLVeIzspRfx49vxR7juvQX2RILW+KKvxMc0YAiVkspSROqLeN87
AItHrdqvX6GxNZoqrtY2gmuOEmpZfaeOqYgIzdBUSA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jFp3miHDH3x9o7F3JDe4edsWPd2uypn83uoB9o6Whs4Ezvy51+ZcVCLuUGWO
QPrRbC/FQCMIlKzgCGXF1YlVZn+dnGo1RauILkkZ826V01S+SB9paz8DvNhA
fCQj2sfKsyK4O3y0pLtc7Jaoje+NPfoDfzwPD0RXsAGAUMfalpE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VWcl+0JbUXnKCzvEufIcVK2DvtT8Dnsc3e0LwysAm/N3koQ8zZnOnV352QYP
4JXt6djN0SVfiK425uc+IZIl1IX6pxHPvEWfvyN+nVNGqIo/Ti1ngvJqbwsd
Jz3VuQoP8GGmW/v7lStlcQDmYjeqdjXXfxV9ziIS3RK6BuPHc8oWyDKzYGXa
F0JLAfmJHG54VLrFMXuTLUnqJg4hmqc1dCVsIDY1FfSPr7AmdH+tLE1GiDit
6ltYVCMnb4vybjmKtOHTwiO5CZhsWMnQDKk5XJIkVROfDgBOr8nFw4dF3yVH
tDzCVE/InBfItBKzoARnP2EjBgMtzr2yrv61xVgGx8LfuOxmeuITeJDfje0a
Ogpm4jO2RXAjF2E8ODt0HBF4Dk4/WBjbbzqmiuWyibg7+Y/OtjqRopm2VDb8
o7OY+2QmLXtkyIjvGJMJCK3KgylWI4BLItEw8acNBBHwm3Kk9byO7lajtIrP
KOwjbcxSo4pJymP2fdA3gB1udknb3f1b


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VOikOnGBZrUImdTTzkgl84ZbOqRFyUJfCCFL6zh1+7rsv1bjy1t4+bjyBp7l
d2gaWvhmzpDp2x8BdjH97kOv5O8BBU8yrfG/h7OyxebRohTGPgSgvvRXczI9
8WJkz+6NCNMsw6J5wfmROxueMFPP7HNRIBWfhVEPgLmuNZXcN5c=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SfNjIK20nxwuH5vwtVxofHGVAyIMYyYmaEmyDFeGL/DSHJSq/1un21CFoPID
blStoJLt8AHC884w6CYQcYYcBQA3AQXjTJ6GOf8NX2pKgpDPlMOYyfZXbmi6
Dd15FrOZcL1j/59y8VmdAt2qjpghJlBuh+0/3JXpJR8SCupcCFc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1344)
`pragma protect data_block
3Jw59kfOiWWrJ7R5yRINjE3PoHS39Bev9GgVRaU6siCI7t1h4riNv4mm2JfC
sSodiC7d1lxWx5hjq54pDL8rV34BIWJ3LJD1YSvtJD2G7DsmTaAKYIN8lHov
MZef1XLSXtw/xrTRbRSXFosVaFWqeAqHj5nTzGEHw460MqC5Yk/nVrMfMSeU
jeES+ZP9a/7hx5dtTkRr84lIWEn3J5fv+vSdz4Q/oinwZ/gGzvwkuWh9eXMz
5G/g8Jgjovl9Uz2qZAT3Oknds7pjfcqqnNZT5XB6zifkBUvnBRlF4xxjh4Uz
L++ge8njIlpPicbgm9fP5RwcdKEoKWZuEBul7cXnyx5uy7+ZF/M+45vQsTwM
04CG+wUjBa/2DPNiCD9/g8VKhF768F9pJEk8/jszydCOjzur3cyyq0NZwAjW
0l9fG5Jm4cDYPWd371CzJ8DX1cHB+oa8ynKssFuQoTve/hyaLC+QN3m+G6WR
8aGmmSTiw5IlaIa8ZKPzh/EGpKshG6JSTz2rk6pdrfmGl6XTgkBGuDd3/pjk
Gbmv/UFb5aZtelqC81Malyb2JvN+BgODGpypzXRdYRQ2BTp5Mn74RXuIvcxO
HuIDIWRrFI3bB5lZ+RxW7pPd8r6E9YFQELPV1xQSV+bP0xJElLm63kqyd3ox
XZBXMpS+VvSvh0elCqDje73nY7pc2fImW+xlNMTDf0HDQhe8mjsLhkugs3Ti
/643qdyEvswJfuE7s+NyCnZxPEK/NhSzJz9QTehkgx99fnP9lwq3i3ZB/WFI
mE0LeN0f7CFiIq1JhKp0jM/itGf5LHcfGcnfSc4peHwSr2AmadIsceFAlJSW
QlEn5f0SntEbrwh7BonnLQytGA7iZcoOs4kv6jSnC19hUNd3bwsbMO6gpmma
ELqlff48XSHDMWRtMSV3iZCFU4ixRQb/m8lSWxsbktm1B6LEwdao7Z5Soij6
cRRiKa2ddfzrEcwANhJgDALt67+buc8cvPFoxcNKCiyNAkH4htiHSyUmnzaM
sMT3m/6UyjY3Zdlu26vPiiwu3fw5wG03cog0TOI8kswpeo1Qx2gFFRCx+cjf
WhLy3fPGqG8l4OFSPMJOTHxK9gkG5JhKnut8oVS6uZJw7rL9yhFp4uBBvY58
l4XdIPMRRPxikrXiuey81M7/MSZbnmgE+wRFJnew7eyYPHVzE6YnnRudxMZ6
JrKxc1rcUrzXZpQWwD50TALY+v+lrws0E6U4VkMIJ45VQUZkfzw4Q59oOxVP
fJIMYCcvDIWRWlK4odKXa0BWGAbiZsyTvVQvh4aSmkt9dbdoL/de1sqKkkGQ
50letfHLzkwSivAKSdkooYoCMpONks6EKIzMuzdjeuXuPzrbyZsMgg8YD/BX
ykcyHzbYc3B0HlayB+3SQjcARxEbO+4RMSuzOH0OcsYye2IrcLqVB4SHZoz2
CIeO5GDysh9+EufyPBta8QX5lJVPa8Uvr4xegdfxY0jKjLTc9jtzi9OYxmb1
K12CHs2Do1zqYrE92pDmDPoXlA+4DWgjVH913jetibxcHdSTRNpxXqKepW0k
D3AXBhAFUSE2D6rVmY3x1Scc4eVhcFVGmmhagKvpbbY75aShtYjmXxOlBtYA
qedgEWgOpKx61Gv0KBSN8FRA2tV5nEhcb0Lg4N77vRzdvnpV0jUz3/f1hSdV
kpGmAST0mX8vGWtTDAvWFtw7UYcc8vp22QOkbkaYIvaSTiI824EKMSHZYcMa
L+YLC4JOZ7ULaJNgmIr/ZGy1Odho/vqvvkR4s6PwpgIK/ljLYBwJ

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQozcLl0ba8TpjT5MNKvR6Cc03vb9I1cM8DnXkjs2u1kELpqU0wgnFXG1onnMattf1on/WIwwYSzl1rbg3n5P+OQ8gBPlgvJQIeIueF3AWrRzeMpQXO5hBVX/hW2b4BOTRtXpT326ebxW1qSyKiAeuVKCjnMOrpa2NwklvwPiMnqOTecKlC4CsB4mehzR/C9KUWYwvNA+IU0iDvdfsDs7Q+C61mWcRt8CDxZqIBFf7iVVCQyvUbRlNZLYZM78YmfnUXPDXX2pSvbHg7eP5VLLaMtpC1UZ+2wMkGCFTcxDdpsiTeqwEC0r5LFFgVb/iIC8hX5UzLV2K46k6HzNOIiBfZg/ETb8WsdXMshx1kaI/0Qa98TPeTZr2Xaml9/GWky6mmMT4pOVY7p3ZgS1yzGV0iE+FwypyAIqDAttgmYiJco0obgxggNTL8INY29AeCCa9UV6WBDsgf35Wa2aMJ7L4x95oaXZUg8T0qrP/R3xvDL/R8+WVkPQKYhZevcgRREnqh5QEyOUSJxMyYX9YL2lyzExIBbHXwl2SsxsMw5oXaJdKm20Kb13YSa3btbC0+LBwAx7SPkVxtvjL9kA+0RXBmMmqSfpFPqGi0iZVIWqhj5RqZSOqsTUOOGW6Nrts0Ao8SRUIpwILFnwExm4RxjSEybFjCbpdF7JdPFQOMsjn/cY/mnagIO4BOJ9uDRcjIz5qz7Lhmh7/PrzDsYTaWnTuIwA5UoirjSK03OHfs9yaWH578RfEv34g/7ah0M5IoXFfd3CuIXynjohNcK6EGadtUjS"
`endif