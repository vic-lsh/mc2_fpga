// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
znYT1u1Ye9PJU8veXbE3i3ZI+qaD3DNtkhKsT5ZYFHupdngBOuZWAWDA8nzS
uwTFT7tBOTbC1EOPUHWueIxkK9Zdh3sCWGlIi+FbT1o/6Hb7rssOH35QoOJ2
kIa9rNs5OdRkRmpOlRcIRjOsvvsctFquRUqTMTKnIqW1PjNf4DguazRjhoiq
PwCWdwUdYzpnaCbqaOtH0DrAo0aTpHGu/cYPLZCGsQqR/xP4Y/P64Z7s5SQg
N/jFr4MPcpLM50tEcj0TBHQigRItYRT5gjjoUpwsPqoFSPZc2Wc6NIBLO48K
3EdBAQUE2tYbdl3rnk9YzW2WZV8ccTGXOG+Slnn+Zw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E4fimrJDFKjgwhGZsE/T2Ff+eIrLbQc9q3HUGE0y6rVTG9HZGIiKeySMKXpW
44r9s7l2GBtUT9UzHzwPGynwlX6xKr6VxKa6CdA1yirmc1NKMdJWmi0y2gxF
DalUbnIfODJAvJr6rqMR+sfYUZBu+zrlA1Kgl/F4twgxS14W9VXL/OKQbe4a
DlxbH+fyF4CAIwa+Atvdg2qs/PBha43RnduWOUsCCiKluETVnexiwLBv7n/1
O2oz6Dv1rFwJH5VtVHpkHXTw52zDSJ46V+LVI7Nr8FKC5vaaVybirz2oB9sV
hU0cos/Ynwwx+WPRYxKErPo2YQLbsfxttJHzX2SE3g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vSc4pxKiCK+rf9I4N0f5Jb/toCc+4q4z5Q51Fqo+f9kZpbpkeOTWt8BIx9zx
KzGNNjBzDj5skJO74WUuDBMsqyIcdvv1glq9iFqH4JiA1XMF/RTL7ZjjKBHQ
6CAbWNXNzVMsj/TVS/YsvOozkjsNz20I4G5in10FSJgNd54Me5NS1vU9OpRp
ep7ihe9CiZoW+FtzXm34Ub30jE5AnqiGzE4rlmPNC/JwJWblqokOxElgAXDq
EgaC/rAK56hPXb45X7nU4tz0kGxwUUnii0OXGkDjXnpC9FTipLzrW0nFc5mr
loRrvz+LXsrOM5AdKHT6fn9x+x7gFZ1amrCgGrKUxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oU06dNqXxXAvq3Dn1lFTbJJswBVwG8Gg9lue6i05ALpR2XiVTq8gN1k1C5P0
KnIea+D+tSuP7dPDA/RJzHI9fTultuKnY99WXF2tGTgsyw1n6oJeZ9EOlyiP
oM886A+K8qnzcFn9vE8rhTxc1EFi7ZFfJ/8DbB6H+XXdaQygme3zbEHM7N2G
vHHmxUy7ourjBTtuifMyc1kn5d+DRYwCNZllvdUtzCPCi/VgfRSW9ZMdbDLn
AJS1tWisrOJC2NsttiZqMpFV8c93lTQx0p7/gSuom3zS1qbtpzu6WxgtdWEp
sKmj/y/qDkFjE/hF1d5aljkHCwdwJFE1YC61LMQOVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JBqt/ply4NkelMq6xRVu0wRK5r2V8VysoIdf7ffMNXvlPUbUy6EiNwlTQKOi
qbR162qpdpnMa8bEGWQ9rWp2k+h7xSYKoGUW7cRWpiB6wsIeRoANTEX0YSeq
bz1ODBIn313HlIahuT+7mvmwTkRiqPgPfU0nzs6LsD0Rt8jkS1k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LtJLk/J4DZwFAh23qEPu7X5yRPdzuLuluGqHACgr5vUnlv7uROfjd/2Y8/za
W1Cnj5b03m4W3DYz+2JhmIaYtRWU0/w5ZBpbbqSzqhrnDyh2juVZxWKf4D5I
B5rJ9teAKTpZ9ou9foiJ26kYFFWlIyQnNaJnj3W0dntntGih9IbYj9vlcnlI
/7XtShR5IMf1iyksnZAjs37Exkdel/78k0zTz24sRz4fn34D1aPG+8JZoQ9d
pUa6Vug4UUpQM/FWg5YIUAGhoxfFXgKbJA0BSMtFSrutnDT6wXHUpMHh8FL6
M0IykpJQ44LA6P3llrN+A2TnMjIeKXgedjRxzqqq6/mrjheI7IIBOMQgfukz
qkqW8cFTe2Zz+tN3TpxzlUYDKqhv6gSNC8dYlrhdWeuKHPV/50moP69yI3Vc
pVrQp1II1RJV5X3WfkaEwoCHWVwnsmdAuug4bLzVdpJVIjgHa1DhBxjiGOoo
F/1u/6mikFAxLQveShtG/O60lPHtMgeT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XKoCpVzNcx9Jp48XfvSEe8MzpJzFq48o7SPqpvTfOiIB7BbWjI699qauB0Z9
0kDnfbbzXFUwCrimuTLyNz85IxxWnthiGFvhb9ZLvYj19aQXh9IQqtFTYtyi
a9l/GY04D5+kjyW/x4c+kMjif9FgM32TcFCO+h+kUgDU0y+mYIg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n5IqXYtpxjKNMIlOvghDRixnBh0U9zpmoLsbT/uK/VDxpHLLE3olA+xCsZdM
4m4rSXbmwc/cmlshABBCKh3uaqICtGBUtWVJDm1HDRW86l58cY5aqp+4SnZq
vvwYRiI1VC1pDSl5YiqRcCRkjCC0pP6E3MGS6ZA3a1cChqGVisE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8544)
`pragma protect data_block
Q4gvFH/1GMoOABJ5sLAjZFEgtxLPEZT/IIS7CuBO6sp7yNhgIrtti8iMPzFy
Zr0ilxWQOKCOjG29xROxPSyqq4GIXZKsVvMKCWQbnINpE51ZoHldhKGkHgRd
T5nKtWhMs12Q8uu6e33qA8xTB4A2sWO5PDDKOtaoxvYsb5HlCD6NoLjCKrip
hj61goQzj3TvP7EIIlbzk0RYfFTHGgODEVk+zfRUqeXD1NhI4i4lNdndatSg
9j93J1Cti3b4M6gpzy40PIb76hYtHRfSXV3pWNE+kN+cZD86rRfW7HGzMCHB
iwywWjZZBsVwPP5CjciaCL+mN45XhxfvIfAi/K1yPyfpvHgUUqw23auKw8Yr
x2Fw4EbRqLPY+U2uaotloxvBLvgdOFNLVwmnZkCNbtgvm4bAnXBF1J3t5CxE
c0WALtoN+p6Iljdh7nJJYuISIOzqc0my3h6f4fBTfT/N2NKo2zz2WUnhejzb
j9HSasyah73eL9HfesafoVWdtJKKCSZ/Wi2IjIiXVugG5qOWDxbK6zRh8X2/
X2Bpzp66Hp6SWKM9rY+jXYtThK28PR1Ee451rEUc8VZ4qZPh8Qv/+yMXtulC
B4j42ATqDBHGo/UaDtMOSvc1uQXWgYYJjqbtO1POJLFxtXuVqpVD+CL+x6lv
odPqUcDzStCu759zjb/Ug4L9b7QAq2drkr39iccb3N8OB946ybYtw88rFhwh
u/2+fkFkMxbFL3TEuqLjyqXsRPpHroNLvCj7r9DC/Ooi43PxFi6tWs0yskAn
djVxZiR/oSlM3Czbcv41kOL8O0ZYI2TMZUZfLWNQJXvYAp81pGOl21DpGjUU
sR26C4EmVZKguNADJcnUd0TXPEZgo2A/9CIl9RVGaXpC8FDdj7lN4h6Ofqbl
hCzbTuGOHzj5Sd0bpAtY8lefr3JXRmzUq60jKhA7jZ+yo8GQE2eJp9OinuQC
5nY1kvHOwLs8n1IXtTk0u4uMNKs5i4u39QoSSONEg2yWhGQvQzy/RuybEmvD
3fZbFZmNtAy7PcnfD9jDLj6XyCeTojstVoYNZc7U3nbPBqpwl9woopTYv0uz
a+gDARe/h6FY7jc2LxQWyFpEhriT38gjilL/k+jjjnISf9ov+RIksVbHBhC3
re/fLQe7cZx0L6fJ4D5D7WxnVhm2vAO7sAv94mTb+uDLcKUo1mTwC091wLPA
fuD2G1JN3vCjl1OtdM+DDIBXvPxiMiV0D2WWZ+YfVeJ/rVaLwfnX9lBGdrC/
4HTUqvy2DhCL5rMP0QW7Wzv149uzQYrQ4A2mLL0IbD/b3QLZ+uB3S/o4d/ed
Vx3+Csy+o/XozVFPoatvcD/oraU2OnOTAGigms3fDzYOkPswuyz5QQ7op2Vu
sjGy03jn8ISWtGzjaNQH8WX2qVWOlPcZiwZeXjFUdEzFBum+zBV7D2u34zMq
OeU9ixB8gudm3i0F3Qh1263Ecpxb5/esdddVk0+DPjd3zF7PqlYnmXDBPcFP
HI4vUEfVVLDvJP17WlSAiI+TZgNniGf/wJ+MCcrmoOgu0Vozkg3yOckJ5ukL
SEhRYyM6AbKYtJSNg2RpdPsK/6G+f79Cj7C86mDhWDRbNtQ2usHnTNfnqmQR
1fQFKUdlOp0Es/HeaHu4GMoYJiz/VGJONAs7weBz7W2kbwVgDFBis76Mz6cl
9LRyicENgSr5dvSTY00zyqKlCXOltvW4lxet8Z9czGPF/IVId0opKMHImzTy
C43fkxgB486flIZex+03EttLyzk8K9fJePMW8GHJY/toGDKPyCK3mLDmvUi+
G+TL9mW32ktHNKYqx0G8NRrRIzTggYzumSRiTkHMoRLOQpMCbQ6wSyxBVbrI
mSAlhaRVkDh7SDOR6b3M0xjS3lU966yGfXb+C6Myj2qxvqfbeydygBhUHmgg
AUAIW15x4W0JxiXCN6wIbQkXuD9aMVJhxuMUIY9QOizqZF/AR3a9QHmebbvZ
qx2F/+b9JSE6xnV5VOv7XbjHlWrLqtni/DcBrkOniHKgaC3mFyXBAduj2T/+
r6AgyqQPs4r/wEjpP2Q/X59BnkrZmcYKIp2DTzSJeaMruApCd5BE3P7CfgMU
BQYGT+DMXl2ZLumvef05WqmT6i0IVRM7flPNOgGtMApaNrL/cVm36sbefN/K
ri5YKo27eSQVdmRIszIG+SkAPW4polSeTw5miL3aw5u1GDwDpRAwBfwvdOOU
kdntULpEIz9QQW29xwO9OKgecHuRy6s6pi+po4wIb1CBwmrO+nginC7mNfeR
z+KKOFR5VlUDoHpd9Ucnh7rKm5bmqLni229Ed8EcDR0S11xvL3gGcbyB40ot
3hHGmXF4qroHlVe7aH/yG0OBoLnsMULCAf6sG/qYHedI7QDb46MPEY52JO+R
q9ntsm+J1eDd4jC6mQpl+jvKnVMAJ+NCwMEkOK31Wy+uwFkGKeBE/caruPLT
bH9fVeCosMbHU0XLLRzrKA5zFv6GIXWqoSR1ANbfWokgQs0R4ZbrejtiwHHs
IhPYVN+haBwWGCS3rt1Z760AoKDRbrgDHSuEZVA6YuUgHDJ5OxOreXptAKtG
3fJZTQEx4D1QMl9FQfYp3UL6mL9u+rI+zqlIjZzohAn5w6P1wxDG8ak45GDS
hf2+LG7PH/xhogU/XXh1MOXScLSvFYC09/V1o+gNCtBWFQO0z8v7w2lImgmk
6WJYCHSdGatrUfhetlBqHVBukInKoIDiJzU44TkVU4B3sFqISIFJUQhYkj0f
r7ltVDuk4kFprJbrg0iDf8uOjEU8BoW4onUmIGS14YqYucX763FirPVXeaHI
T9rmGzqo+SDG7dQruF4WatxAaEGtq259KxnAenTpMAARWv5JCRmKkY6EpFEs
RWotK7V8EGFoAQT9QTtOqVrJyHr9CdjeCn+PkM2BhYskT33LMfHfLk9XEdGo
P1Oot9IYyeqsX/uRtxbwnw5ZUQrzz7ZIdOPtD625AepTTBGF7ocXAO3CXJdf
ieucTHIYYYvEDChjaJF7JwJe4ix+Zn9bFM2IyC3TlgrAiCXPAbHUv1SVCfV1
RlKovXPqupE5Qi1BWWXh2vKko7RR6w5lgA+wFGlXz7DSMgoUcZNd/zlvnN+7
I/sRPCpoqnyKYlxmL/uZ0HoavYEm7asU10jzmQokFZAzP7lhkje1kZDcejKV
8hB46WpQ0jBGe/4Hx5x9jcRAbOhh+wfFusEGAGz58uh/f0foN5qUiFOyU1st
H2tmR+5rS6S6/fMYrhLLVBtEHUlM25ODKzCQ1JpDyMyYS9nA3X57QCwdMkNI
mOhOiDpm4Rf1mqjjM1hxGoQEU7lQ6Xg2Md/Ii6HNYyG0nD+ujGtG6/c6I5KB
7Tbq6b792TJkVkk85uCU67L4wzrOgmn65Hco2lAS2GVaQavlz07VRuk1qYCx
ykrXWNERPUcw7Sz8UfuJJuym8Kw3w1RgnmZER2JeNcUem+Mp189/420fvBgL
xBKwBs2sYFFcbTfBma5jC1iXU/YKvjPLpx0Nfq2ACYrlA2fFF+ATNR9cEBZ8
uw4izkW2npgX3GjDOYS9/jJ7KqgEGF13Y6bQi2NCqZrPRJK2TjOH3YVk6qx/
h5CC+YpU7V6SvAGXSPx8re9tLiH+vPsA7+2wjYF8RlBWLUOBEJjReVJVkwrs
yS7vKoXWZbDRjzPaOtyJ/lZbxCn4OmvPUEWLTwS6Uvt9jJOq3e7UmZm1SiVk
CErf4x/iuIANgKl6A7VOIyKU9T0gfRO0O73JrvGNSjhJnESJvigGeU7940lH
46KPtde1be2jxEQJdCnF/iA3MJmMbWIwJu3NVufwbZoca6PIjOthbLLfAh45
PkurGJXrzeRtSKJRKIn+V2psjx3fx9u5vCYUcT/mkQ/ozpNaAY8FG35wCStA
8xYxivCcYND/g7HgeCChuqKAonD+Lk+8UXmFtw1HfThndGeA8ZLNJ6XvLtNP
EygMYikELcpcre47KSzKTT1/g+EfTGhg4ih2HpOHYu57NwqIj3VqlGOD08Nv
y1qN9Wkazw0FmzAPv2Sr+6wRPSQLVe6I9ueUqOHYz65T0+Fdk5LzQcIv9lnM
4ZgskkY6T8rWhtpXOvtMfUNwAIkFXuYJAT/o7MhYo93w0wYCtGkVYS0qIkfM
FG7zxq4A5JvLFw96w/3klgUiCFxe6vj7zJcyJc8ZVnl8vMOQ6TOC/gJNut6E
7kroQDYcGn143vxIL2mAO5EcGTTi1DauSRSQ02w/SUPYcbXNzcBScFefr2o6
oMigwc+qtJTfMDI9UcJ5pTF5ZYE+D6Fb4vR0wtBsL/jJT4Vr4A7r1kxdidd7
X2iEmThGUD2Sh3vKU9cK7M3+NnO9jWxDp3UQoSQOLAZaBJwea20CYcTSP2EC
1sGBC3u9PAJrChpXkls/nmOqeJCDIxlqXUSVdYUepVJuBHHJkbrVA6WvBqWM
K5IRsOUdfoKE0134XokUC7S3BediFJjd7C0x8ISFlR7ugK1Iwn2zKuZXBwQl
XmkUn5y46IlTehxu/Ihiiq9BFl9RKNYHIdAAW+sTHQwdQ0oMVlA0Zvb/dpeE
9lyFM1jRC1XPCs6hSh9fdlsvIEgbRfrP02+Vn416clxKhojTdJanXQJIvOgQ
FcvE7rgphKixIvym53gsb01+DRV7KGreG8CnOyWX7kC3vU6pcMdJmfeN7dX4
d7nnybT0A15KoukgyJDvoQUpsESQ4oWqOPKj5E40QF7Cs2CAl2eZp57U6AfU
pc1NtAkWn7ApdFx4PQnkiqIaZ0aoKztgXkHswmTySAUbMNkHyADPitdB1/3C
FncP5/nS72eK66EU8nILii2wGjMQY/MbyHmyAzi4DdislLx3gik94Bjc2Vlc
hIzs0wgeBg/vkH4PLxm9nOrrTzzeSf5i6AhriW5hR4vcH0d0zX+VTkurBrLF
pGPK7sTJSIN8/uRk7fbs25hWztQ03vpetMbN9brxmDXkEDtz2jBrabRpxWXF
gessjRxpZToNaFrWXYlVzXLSPVkd+rdYOcm0/HznKEDbvyx3V0tn6vvgH7Da
sKD6k8bal0RSA1/aeIo0KDgVJjJ5J/+HTxy5wXqUiEMaSlXTEVffgzJvfHzX
IxAPInQq+o6iYaedq4q4UVN3JX7NPM/D3w0kVQ88x8SJJg3T3gxhp9YOTG4q
Tr1bag+6724LRkKs8i7ZfDxQdL/6F/g9V+7s2P1wosMx/N6CC+w2Ar9R8VLe
vyusItOqpgU5llH5rPsgUKccnVESJODyRK2DzkJyNPK2f9WGPy9fU0ln+xh3
7pljrajyHT/NHwfbRC1UwkwyHIS8xCp18nzkrM+Ok6tSk503Df4h+whm7juM
i//CC3raUfd+irDb7vvb/Q2H9hCaqOVHnBQuWFtP/mKK1qYZL7hH4/SgqYft
2EH/vXtiuWiad+q8Vp/0CA/W44fwPWydKFenAMZpCLRE6AFLRAg1Ia3GLsL7
LOlmKuYtCbOeA7IebnHNiTbcPdZpKDPoUOAkzNhtXoUdiSZHPEebZ64WvKHN
0iIFPngDk9WFVTI+h6VOkHFK7IqWgLdgz85tBD7y+oRrOW5oONnpWdGDjza8
rSNHgKI/EL/GA28K1JFuAGcFwxZ88V3qzRT23YOqjQqXvrkJzrKQPQ/htzH4
fofHrROn/X+EVpHrJvvQDP49bi8e39YpAC1jP3pWaH85KI35cP3Mm7/soIDH
k+jNfwFHjyzdnTJ+7zo+0jd3n8/tZmMSlk2Gc+qOBZlWX5HV0uEyRkuSQHZ5
a86m7OVI9jw4fB5OtirTloc1eVyeyZpudODMADx1yCmvRilbe+ViYcjiGwgx
iP1WStHao63yWv7p9EkfwgBLOSOwwvlSWhD+WsBexwyvGdx8Kh5ZKMzJkYAp
D91lGSLlSULuU+LQ4zKYawzMaPmVIi4xXIUY6gM6VtBKhJRLW61MAqnnsXjL
8WVdYOXRr+OueVZP8hjK1S7iFprvNNPHt5CJNei8UkadJxLs6fTD/vzA4qhs
0ImNX+A8EqpkhBxRRF4Tz8mcoFzB3EKyGIvIBtNwS9y3rgSTHdnt6XWoEAed
af3WMQS8NlnAjwoL/1c0NkqeoS2ZNxqJ7T/tDZF3fWd0zQzT7y5iQd503vhY
z0AzG83ryQbRdE2Ukb76iiGKwBVxQJmj8aq9qWNmXkBBk1WTHY/ZlBk2mo4J
yO+6Z65noc+531QUjMHI5L9bV+Rub+43oD3wcd8iRLYW1dSP/T2GxU3aARCv
0PVnyFnogN1yDY0VC/UFA12js9EbdEFxVjMExNdDcIQ/SJcgzjaBNAt4bvuE
VnCFHdY29QAzviqJdWXJN42NZfTbs0pjHYfFo/W/E/+J3uvN7hB42vWFkf2V
ad4XeRAS++Ovg0pwr6GvIyNu0wcRFQaMj0a03AhsBJexmtT7uupgTDejFKcr
fi9NBrNJcYnpC4RD1Qn8rMBogZMnokYql5UVL+PIai9hGGXui1Z7NDau4yDu
OE0PPmI7Qj58hRaAoi1+jgWUJl+vuVKW1krhEhjV36TZeYFm0qUzum5IzXHG
OsprCvxsT2Xebynd+mZM/ACcGQ4XNKF0ctnrXej/jQc9DQ0bCeF5nYSUjp6D
dpulGu7Ih+bOAs90BYqR3Ww8KoMmcS8hVeCqkjWbrdWGMCWt7mhQ7ksxICXD
34nQ/+TnudvtG3fHFQ4XSxEF8FL4b+tD5U0e4qetdTsN36cioceDHP/fJt3L
yxqDPaXBE3xhCnV4ziejiUUwrBv57SWb4nJyGx2kuMxwKSIQc7gXsqFmtz/a
2IlRYE1BY4KHlEkhCl4h+RIX/mfy1ZsCICMXESIn7xiJyxT+zy3aOPnhsPKd
rNY9X1u2HX9RoLyZ2QWg5AnXB+NrKVCN+GZeIRCcTokBlhOEqT+WcFovdNHo
15LVuq85C5qv5XZctfD9/92hZTRPJyQpklqDnvtq5sb+MufHFx5vXlqmZmah
EA3zDdPKBV3VvBg9NxKyTC+5tzwdJq41EZ2QZKxAjrLzMSR/M+txZOkaJ4O+
VFYqfI+kqqQalYO41e9KrNBy3S2OSs+MIuAP7h+WElCEg1aqL4DcnteZDkA1
KC2uE3kYfripYSZbf0EKPunq+Lt3xPK6npyKZKT/HK3zR2MnTwnWtw9RTZLT
36zMosl0qbQFoj+PTjD618cLThTx4BTOz0EElU2LerAcKxMEtAYc7RGpCANv
ElZRTwVorq5VPdDRan9zLm8jfZzGyMJgLKpXaswUS1MUjPgsI9fu0dHlMXlZ
EIVgVl/tXjDqX5yTPQ5cqriiIq2Q01eqLJ8BR1qEWU7z7ZSWQDvylMLUkomw
I0sWD7lb09+8xM8PfokQTY+MVZAFf8X4TYxU+WhzKQIk53CjUsg1d8QuRWog
S/4GP+4dbbOrj8jUzyhCL2vArW4Oi9QY6kYM5BIduLauHFFnZFgak9t6nJ0c
QtF3dn/9YqC0pqRX6bULMwoH1GOiG6IbRcIyIdoI6Em9HsNjEkzfdYFyaRT5
Chz7kT6A2nH5e98h4dAlwbSGz9fhqcr3UrXq0u2wXW0lW+Bg/QWUD+mP65gp
/rGeShcmayvbnkWpAWT8kXZF23a7UcI3RJsXjGUXxoUa1aD43eYHL+kVf5m/
4cb1TfqaQCIOnD3eLSw4FOTTwHt8BG7ymEM3i33UqjDb+z7/yBHuILW8sMbZ
cnMzrcnGtx/ZM44pWPz8fpKLA8FEHsemPn3E28gIlWfXi/B32bZXSbIE4Z83
LG0xzH4r6CQbMW8onoRwlv1wWKcSfqwaWUfs/ubFwbMGyahL9Oycyn3EY81h
vcV4hd5yJSFF8xJRB6RdZ9CNrT4Zx0c0ZG0cnK9BkNPNkZCdkzwsgIxhVVDx
L1OqD3EWL42uE7lqPrBJWvbbxL+cCbNQTbktwSolYLzDi3OIK42CfEsis5zh
1WsGxGxW//hCWVZvUqiHpRT6bAQDy6mPN7xDw+kexcrKIuNBm+s0s0Yuy649
m5VGs+JWVjba+0XJjFwZw5stcv5pcWFK9qt9sN3Wm0YDXhUyFEO/ST0DJYLC
xEY2YyJbDXEIIwQwgxnRXgn8YuJEje3ThFPbd9ohWH/hMF46fcMx6ShGPLt6
TcQblRHQEoBfSDIIljhzyDvTTaZZbokjm5jTrRgWMGIkzxMSB3C7kE57e0n7
BXGhQbmpnU1SJIhrfedAadJqv4K//SYBcFHdAyLNTWiy9k7uvULBIV+9r7d6
I6Smp+yDZk4lrIzNTLrEdyHnijdHEhatbCIljKxqIbymogJXMsCVb1hC8qxq
eDWWrTrhBT6QhrAmKr16s6Oo3RZgAT6V5bNKFO3/98HaOzziUAD/TnRwgFTq
Ut1llkVWczR5hXYElUkXA8zt3NiOLaag/aRwbHDoZRp+LYXa0GHqyxwJWXdV
7xQ7mLtSj3cBWWlq22THG7i8SmC7zWuuky1yGmOkAHD9u46Tn0waNdHuL5xf
zfyKpmpVR05QRHVFv1cPCwO+1cuqNP3QzVy3NPFAhjuK2raS7xExExKoEYgl
I8Mk0ZSKK1VXzAGgt8AbzEFQ1buU4p3rTfxBJ5RGs6Bk/4Nx63dc/R67DVa6
2ctntQ5uSLihl48bla20/k+84j66jiyeqRfE+i59ZWw9trhiBgCZgROLAnvJ
BIa2ggsEMXpUpANK4bzXBcG02ni1QlwBLrKwFsJdTl//U9u22yzX99Wve1OO
di3pMb5UtZY0QMa91pfi9CSQJ/8EZeK1lzY14h0RRCMLA+lp9DZ/KE6Mf9zm
YcvnXPh+2S/XY0yuOJyuSamwZ2IWpmaDQyUjXkqh/53dcn7HCDfnlVbo4ren
cBsylFVnW89JdBY8lGJeE48H+2/8mdA+L86hXq9lwgYDEcGvZsFmoYr7YGSO
UOnjJy2vKnoT057NT5g867KlC+PC5lD1LEhv68sr1MWhxIkAFEhPvdOnZ+NW
Dkzwc1yIQGWwYYPURPGUME+gOSC1fzponEFvUWL1HLz0KYdLr5H+MpPXYf8r
15hfzND0C6zGyb8afj5Vzqj0ZBi/Voq0YTEyXuUAjlEC06m0pct94tb1aXX5
WtRK81X/IpYYOL7qrIqOF2qVzpTr6r3D0N2AG4J4ZsoDEmjFrSeLbNYLRYbD
gTVQh9hSBKAz1xZh4QItRkZgTTkQzAl22Gc9r1X6p9cdKuH6pbD4SX96WTaS
t8U+xze9+Mm7EZqwplJZJUC1dMoqdj6IPOle+Iu8bXOLuSh2Oc6cQstWY5V4
LU1SUuhebjYZ3jxdOcf+DcnZadtjI/8siRUmNGLChhgLLoRWeRigtU1PEzZz
mI8sqHl9Fb5G7F0xU+f1nWKAaCfwZk0tYbWQYdHBmlznmgaOPZdpN5epvr7d
fXWqxU06LVSr1T5/7XsdCuxYuq8xIUMMG93OafxtvRMR7uc9Dt4pX6CMRR4S
M6sDkd0GQgu1OFBu2FjdCGkC1IAA+nxRki2rGSdmLr9DGO5utieX9w6gXs/m
+4guxUeoF927rm9zBnInP5X3YjSe7sBFXhz7DZ7pe+mQCxRilHIhh7CYrDu0
b6Ah/XJUpwO8MtTcUGpxmjtX8867c5AvTJusK6uY6c5dI0z8Xna8aApyXnd/
HuWGvz6JWaLnbubLR53fC7V+FXeMhe0Tgy5BcH3V3VyT9kDN+iosLAmcXfch
Y2zxXmufXW2RS8RddupCUxITitrGfW2av9seLW/nt4tfZ1WC4SMLQtpOGxxr
6CZhC3QcVqgJkwFaFJML/OA1EQd6xmlWxt3cWtuxHE5ZW2QbN1z5xEsEm4jG
BJukUrj61fZd4yo6dnkU0cNquh+p8QVaSnzCZWm0mR/P/b5P+k0XCUpKyKYZ
jNc9MHS6bbm4P3JlivvM12WcL49gtUi2Vs97D1knUzxT0STtHEXPdMZUqMh+
QXLanLszyTB10erFmXQHOFBxOlOTXrF8Wah5EJCr1/1pAFx92gPOQ99ck2Re
DttvWBp+5ugSzzWtnhTpDiDfq5RRKm/brdRVQJwn3QHLws5dJUgsPS07huZB
+H1MqOf7JoTjId6tyeZXYf6u5iUaT3t5ifnfbZT2vyE8Yi4AnoHnOBK2c0jE
9ij2vux/Nt+BY3DC9ME+5eLnOZ13HSXDTQ6mxP/wkWsn1TsSUC1U7dMx/eo/
xWJ/58tb4QYlTFQ7QZjySeucOqqQU+SS5IicVlyqBAQBp6ctl1+XQKjuKHD/
DAK9RgGiL6OxzzqvepL5m0NHgrTFQsf6KWSM08eBBBHvQYn5xdPTwSgqZprW
0zrv0o8WUg+bHPo6ipHpM8Zehp9diAopwZuSCtXHmCrOjxSLEXSPtPZzK9eU
zMVslg3DGTsN8KuJNiiXB8lsXzRQOcFW/YTIhI7Wsx9evCy0L2bqnsavAuWl
HMRvyMl8Q7oN6xNiG9uGLtC965WoGeNPKv/L/sHDIvb3mh7gkdfgeV05Oo5p
aCjjO8qEHVeyhHlvWeZV8krQB3YwaTq7E974mFo5DVWEoXIr6AEc8tnvAVyg
n+C+6KYrq6DulwWbr0Q6ibtQG59BwU3VXJHlLoSjHn+2JMwluwuW94P+b0+O
K/yuX1LLozeaiKV9C5x44CPFVsESbPoJctBg2NI9+SH7L8cRiuejtb5Rfn76
jN3JdIiBQRL8CWcxEUH5QF2Hw1oZ4MSCGEhmKesxVJ6wzTfvmvNiZQaomAqP
v+qyK9fXu7FYzbsGcjHyzOp8dvJkZ2k2xm87XVy9kczyIHPVlnPM9ra+9njf
moGoGWjcjHKKUKN5e7rOnp97v3AjOo4FhXovKExtVLSUKz3zkv41uwJpdYiA
8uje/3MyNBIdYbKKWqUgW7p3jfIF9s/G10BdPjg83/aV7+938iGxrdgC9ugl
aEpPeVAB7mjbVc+c6LiCOVNrSLVE1zK88vZX9nopsYim4GXofSOQx020kO+6
LoIhpdJ9mhUjP2PgmHq1WdePyqxYPf1+FhnLX4j1aFrDhYtLi99BqeDWmYhF
08FdH3mCSuh3q9sVk7xM1NRfxadt+tHMKQb81AidZdnYwQbv8Ts2conFRdsF
m21dgkMj1BQoiz8oC9g5fTMno5e0NqSplY4jS2CwQxRod8eGaEGqR+Y1vkPj
2+02+P+0eYpinF0LyTKSuFV/qC+IlnYeyvnUCFw1Xw+kTqfbtDTrGjCyTWjc
iNbjqAeS7RSXrlO4ns80Phm14xYLxPp266m+eoqGIZ5s1jO5M4WF0nSgacvg
UuesW+tYqBp8Y7yps9DijeLzdgHaCITXar2+kyDt79hTcfdH/98unOhkqjay
IIZPnTvpY0390KINEUUmmceOii5K/fcVFX1MNC7HnSWP5a88MrcUcnq3SuEg
Cw5JyIjHYU6pTmN2lYxJIR1h94Ulp1V2gIk/caKA0APAogSb80ck

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzcV8seFSeltoMJ5dzRdZCbab1goMSh7UO0v+go/0Kq6hGrxxFKHC5dRlVfwdB8IL4nRvbeBJ3ao+8f0eLzN9Gy4ZaG1Ji30sYLXnlPAHdWTojJVokjjrb+sJdTpORpL2ZYVQL8wbyi15ntEaJmlx5hn7bvBCoCaZYwkqJ+oA/rcdS8D0O3Ell6JMozrObH7uH8HI3ZdpA8QWfXkopbHp0btrq6/IRjPQuSK+j4p3dlbjOXN1T4nZClWSAFqSi/tNcJ/hW/UnMflw4fC1tFrT/M6K3FO/iQbSwO4QKLK8I4FJpV5KUEzhPOG1FyHB48NxxzLHTRQseBh5zi+X/zA+JeqKLVT/kJ07iKiCxwNE7CMVjOaxTy0TGh4JTF6lle7QwsIlqmEOFJh4bv36FC8Ok+NgI0LdEK8qa/ROl73lExYmL3wYVtIqYrxAakFHT/rgqn5tBNmuYrKpweiQGJBhHOtn2evkqjU/7XiLko6zgdTLl0D62G7hBDNXM3OY0naP8c1mfCQc/zV1qb5rj2YWwWnlkjhdbF80+4CldaLJCfEXH4D6P994oEJ13ZtbUFNuk/JUHRlqZWYv8FN9ICWKBR7Pgeo0sFUh2jKMq27Z8iypraM7YYYt75X0KpKDW0Y9DtpIJwc/ulLXrFjDtqUsvVKLHrPwqN//Sh6ShoKkmPsNnUz9iLfqf4HEM4k8/9tti3E7LrQ9PAw3Bf2V7J0BeXvcieMvOSmjWrjIpyunQs45cvIIyQ2EDOfDMQ1noxq/E4tZG6oMjeUzUmogU5f4ESh"
`endif