// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xEPtfu8AzgILJXiedXty07VX35ug/WFz6GPWbYfJ2o1UodOfy2kFesKCDrMV
7lV45Po/NQLPJyVwX8jDk1V8FRT/eR0uYFtVx61PRuzVhTINPxlM7s//Xqsh
aDG8Ca82HjTXEhjtYtSoraf9drTNVKrc6uUmmxmG1OMZpLuPNjOorGfiTJeu
VIE7gKVfk81RYyuf23JPccNqw+DmctKV4mozHkNdEUaYEJ7doGFKF6CdZfDW
QEFXpvXa9iHGev9Et66VZsl1E56pWfTvEgPEvGqmb4KhsQJkJWwaQk//ppsF
DNl3MB+0NtqVG0DuTTX+xdVeLFZRLxzRprPMGBYE7A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PwlzzNPGT4sBMarjHiwiZuRiWeR9ojxwol563DHA+cSKL29ZkIR8vWhXPF2s
iApggr7piT+38408xMVaYK5H06LUpNxLOoyyb8AY4w6FB78/0Fvxx3kRAYgl
ZH4qIECQEsrn2opJiau7pV8UV3xzFYDgl0FV//oqyRmnitdCgceXhDn5ngGb
DD8Rpc7MAXO843uCyPnrOE+1Hgjr0A2RW7kCpzASfOSMtOqOJ5ohJYESnKi+
rIqjCloCQewPYpIhU/zpzeZvDQbp6n+lCAwuIUWsHEE/lBGSriNDM6x62ygl
iDwuKc+HOafjX8VUl2bm9Ux1QSJXuCwk+ZnrfDsXNA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
twy+NlBGG/FZuYPa/8PCywtDs2eCBCwenWqjfU0Xrpd34Eh4ZqLVsRoA7q7m
9pNqHQEqnM4GJvXHnJ6e/TAGHfq9s7IYQm/IYXbrEk2auFz+3wgD7krSHMG1
fZ/1+a22zOyIs0NQ7nM9PX2wmxiaSnqL03CVFxO93p3z2mzQvK1gNxj051u/
vjp0HohrJySmTTJs92swKeCrJevMmFuljHbK5eALqT9e2mfkl97lKiPLPgYK
JDsWI2+6oYLcCJOk/cnsTZ32cyuhYJI0i6nFMjKYKYmcFF0w0PrtQr8eordJ
CP98B9mCUxIaPOrn4f2O5337O/zl9OIR8oH2gg634A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mBZxI1IrDSDIiiMDGLiGppSNr16HQfSeGoghmjJwq8wBkU2wDA3+Vow4Hlvh
iW7/1M3PRTWA1pQVr+yDVwkQ0pQCV7s7VfhRmE+HWmYqomvpePDFhcGg9kTw
MUg5H+LUK4J5GxSi87ORAcND+lp9DROkMVXQ4phexIPai+CjfOlWBpNKnjhI
ZqgNN2WHPoYf9CFlcZrfYEr4wxhd3hHGZlH7lI5I9H1Ae7PNOmRgEwPkkCTu
31kdMucm/80n8u5atpM+pbzxyZ0Eew8cDU5WSbJ8KTmMHtwzLlC0qjTAAYvF
SQARhjjM6SAeWsQ11qKicn0WGTnkTdQ3DRJqkIZWuA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NfF1TeDiWAqO1FpWynQVA4av8khFQ+6D9WGg01kGqo7xrtWCS6mU7H2a8KbH
xEGWQOurNxX08F30egdza3tDqAPl3I0kmC+kqK1NVSVt4FG8yCL5rsBvmfAN
Obpko09qLm/3LG4bLk5Gir4pJH0gxd82jDtltjz9RQzbTMI+FV0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sLzshxrqHwgRQxehef4zP+xKBOHmQ2CqoDE7Z2B0F2Lh28qRYiLCPHj/56Lc
iywEyVTusM62Nk/BdwUfZAm5SnIQFc+oYY4mIvJVmYTF9sTzOgVA0FVj97Lw
POcwHPWwpuoXobV4uWAp9uuK9R0Cup4CdKHlcuyiBRLF4CLwfNS7FAj6yomn
1Qp8O2PApI5erbeYGTGKc6cAENpTqi59hP3vaYjq1geZ3ovsW6HGtcWH6/1g
HSxNrK9Q3ZFDHi4eRWiDAuJTL/GVJ+Z3Mcb8mmjQJGhGdtgiAEpzqdXXIY2r
HR2Ip2Fa6TN0p0CnQN57YeCSt4A6cAiT6ZOzPs3zG8oHjabK8iWbqE/2bLFM
AuinaVSYsVYNnm9Y2mRUHPkOc3GpJ7yTNDh8CSE/UHmvFLsOzdZtLIQuDqUt
wifJzfsq4iqiWvH5/od2UZzE32LU3bGcXAnRonqRVR7HeCxuSbfr7oXBuFgU
+Ieliq4IxE7SZtOdUiS7hDSVqlYwDKRJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BtSgEbSqs14aqagYGvE+AbwvFe1mYXCnPbJCxFVDCWWiHd+gYR8rVEOoNKG0
vdQBWG9dBtNiokQoKbTP/XIJwTjalNrOhHymnVQqYDGOCYGA20JMz9F0xaDF
ueJcwo2vE8SdVCrQJkFUFi8Z93vFOIRg44dqDNoDIe3ph+T19Wc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e7JP6L8yVG9eKIQll3TrpQGFKXR6H3bFF4b+cI1XqYH40JUVTKy5icnyKZTP
C0ZJRJLJuCoRZ/mF8WE4AppTdkrSdxhOEQGLBfWJWbgj96qXxfG4gQ5GTYzS
AtMqmdLI3MFc/lsCr/+4hbS8RUvIMEUoEcikpDSTjHEeGzHU9zg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7040)
`pragma protect data_block
dsmizcC1EFAbId/IfGnt3ReAUhJG06r1ablaJS9wOE9WbhKOYHNhDX6Laqyp
hDMJX2FOYOuHLfxl3f43C8pxcB7MX7x1aIk8byit1IP4Z7TBHjA9s421kpD3
tAkODrbU52pB6B0hQZhC5bKHaLzGlW0eBWIBMJdi+Rb6MzPa5CsYdetvWNbJ
GzpkwZ18Aze3eX/Q6GDAKRhNjINR7ElNx2exFezjv4lbpREoLkT0XLG1O4Ye
4gYxvycKcsXIcnu9xuLJC45NZrRDxmWc0aBfzJiSMEGXvpvN6/ct5IYTXQYO
CGLo/5L4Jo8+AKEeSv0Znf9fUoNMYFZhbWFP3bRxWYdcEQdCjCuFVeEKGppR
iNAIp4+RPvNIjQHYdJmSkBA/rtfl2OAmZDk9zPQMyzqKj6BzkSPt3L0mPiy2
ww8MMYoz4NOEwoxM2kscq/w+mdAbY7/hxw7MDZbE8J1t1OaDMUGT42FHgeOj
lh0wGHWzWdOrHXwb5MUTHETr0E9oBkh18fL2s9tCjLCNCItS8nQ6xLP9l2qC
mb3xaWlKbEFzoUnLAcAJYL2IJlH/gGi9DiBUWwLxvhrnhP0AJ/u7iTSVv76X
ztYfoZOZKPbb+h9V30cmfwuduKhwEVzIKSPmMW20SL38fHS1y8oeyVSMTYNb
kQn641Me7fQIp62K7QcTfxx0s9/e3ByfNL8YH+b2deZi/tbPg0HN2ltYAuuT
iGWC4vgqHYhPTSK4Ls7U7j03nktZcvqVVaUUlRaQ10o2IQ3rKIX9w49nqGB0
7eKuGSiePvoaWqCHlP2e6FFGMj92yG5rV+VG0TEG5spnl4yWKy5lYPcPQJgR
QQL3np9v+1HXHhTb31H4is1VY6Ms3wYZ040BEuAFkV5hicloqf7G/fm4LjU3
rQWTXX2Xq5BUG2kVP0IRqx62zy35CVTkhAsqUriHK0Vzgtl8y6QdbfKvwlJx
xnoGNUKabPg5LCLdyE0ch0rLe2T5fqn8NLGuwFgclmDiREdtda0icnFEe+Ml
4lbAIIbYMVKJHzn6F1x5tyMavE+sJJH+Ak0l6pjtfT+4yk2pQgDlc/HNfCSF
0TneY4cOfAxSxgjI3Q3dQW7V/t1ZnXirJojtSP0vxiFHBeSO697+eaqUNBhZ
oeWENhNQXlAECNM2WqCj1vbpczidk1Qob5Wqo7Fjzf9k+XV8fazpTsnNZs4i
JdeZkh5g/Sg3x1NP89zTsY9nuDWh0wNdqtHQeRZy1w6SAMxAszTQqBR1cqAI
sKtpDVicaC4UvPYrddEViQ5oAtqCruFlZUSsbqjsx6GFR9Afq7XPD3L3BlBh
4ugkWmL9hoghT7kOviZQzLvoD4GmaW2cyyK0kVb1jLhG23zU0A3dUagkN/ph
gYIbGHlexLELj83DG6hBvwTPnLSly57yC3wYpiutJl56LUzAL3kuvZPmeEbs
S3RTdKRCmuZitYkwhx7ckm7xefyXxamTUF1Ta9Z4paENG7wnJ581HFn5tHWg
rcjF2VDaPpV32ShzChfrl1cK/7ToHVruIy3MeWH3zCPpPujDEKdeMmMIRDnh
5WY6LH3mJUAQzjc0oAoIgwRZ9FokupxKZNp1Kx10RYgLQKbdM+MCDtMdbUF9
qUTH6ruu6wdjnT9IgAyGwjFHQM7ChPqCXw4HSfJgmWIZ5OvXZKwHPzTauM27
EPhA3clx8EPASRhqvrHRNHpGVvHsQc2+l1JfkWBeMkMRiRYqJc5AUPw4mEbB
0aYWZqdSqZZM8ht5R6t/VNbRZxLFbNVSvvetaarJdWiynxiT5nxQlOHz3GbU
Gg+kzVVv1HTS9DwhYvhiimHfPSiPF286Lbqar6ttASqobYYl5qIQOQ4vukVh
ZDyCjxXKA7sAwLoBPYfcCtenDVCo6BOTNsvCWiWe1NgLJoOAy2TGbdXpYgsM
46o0bOuGxN+Vq0EVbcagrNu7XP53XM6WEFllTCxDToqpSvhSqwMjihrQzIYh
h6MKknZcgLXEQ7E6RJPKQRwmIJj9LhMyXgxphaYAxLv1lu8lVS73MklAXPar
IdgZqg7JjZvnpzpcsBEhbZTONl6G/a+lWum6HlmjYGQ6bTaXpBYDRKCndeGI
e6jdEjSLIj/EMN5Q/Oik8DcOjDC0NOcYuvkmAI/EK49PuWwPm0yj7fC2JAeI
rC7dao17EW4MrodpjB4RbRHq8kaElATTyAGFNruzIcGD7ajj/elt/wB1NZPO
YY6T25H9FwQrRS3Sjw33mrmyEO+mA8WqklI0d13Nb23Ita+R7AoVRsbNPMD/
UEy5Vr37k+OT8BBQU+aQ5XjQKoTvZ5u00tPgtOzZgGXjWYQPCF0vUkxm0i0m
GXFsiCJ6aNINmNWjXewQILduA7ZPaN/9oCGApV6sOmt88BVPnGKfz05p+wQl
zgprcW5mkfxGFtpME9KaBpZUVYyqqCzZm385IE1xgs7QQ4996aTKOSLJG5vc
P8DmDCiX4vRUCC51WYiwqGrhZBi2nYQYIAWutNiQFEItM/huHzkHsXRep7N1
q7cLo6fywM3jfZRo1rS0zeTtqQUbvs5wmwezdet5nu3lYI9tKDoIoZWrhnoT
cqiiGOPu082m2r8yzQgZpdNaCKGHmiWi/vVdy2gj4nBqQOA7P7DnAxLdJmrX
MDF/AopV+OcS4/4ZKIq8IEFJw17mF9EbpeKGElwxP7XCmDVxuBgBpZsT2pZo
rsUQvfjWhtUMZyby7bi6bbXdyblEInfw/u6sk1BWdl24hn2DFZDmMWp99TDu
+MUKdYBf+SQAvmru3IcUkplc8Lguz2WlCXkMdj2mr5d4H4Ss6WJAyAi1oahr
dmTeIxPvzM7Rit+le5QN1mMkGLI1Cqel/KtZWbQBAzJpfwx157VnejoXMI+/
IoIGv+9MRg6ZbVQHsJe1Z3Iq87GUmFn3IhlZmbLGlLI1zb3BCV2yhWL7RBCq
XzoVw9RYp7+Oe0RLYJS+u+XQjy/asQO7zlwmox8HFMBb2jcqqOC7ynrCljsd
WniWGFopDzQtNmZPBx6YCyVvWIjHiaWFtls2BNp9f8uBLVwCpPIBPBnL0eLn
PnqlsdSVEbhql33qTjpSFADfkguoWa0rPMem2EZHeQ3sUZdOgQc1t6VpdVHu
ndxUwpNW0ty293vwaO2GMaYZqik0rsfDHYqcITOb7ziCuBdYPkQ3EsIpmlac
HGjt94WK9EI/8BQ8uHhJLWL1jvBPi0HLJwKBqalvuv2BDFbD89/oTwBwqOCa
8Xkvu6MiUQXEDVPYOB6GqzhQuPaBpWhYRVIq0Es3qiX6voDJ/MAoB4ZJH4/D
+IOvO+ugHxQTiLspeHv8uSHxjy0Nn0RxSr87eI4SO/SLlWiEo214fZ3ZzGfX
hbVkAR3YMMjNvPhvie0SvCNHBoxiJK7K/LnvOOmlansACJKYw+Xl++6HS1oo
Q0yoW/+qgDeZ1szpD3UId6pfMqqjIiDWQeWsSij9SvBqOxdQ1jQ0O3vbdi6q
JQ3c/Ac3+1RfaoZpVCN0dUSKuG8sUNHxlCTXexCIu5uTGn6oQ45/lcsVQ9j9
ygjFukUc6zHwk4cHs9JwcdWfpUlwLQnsaQbAB0rnYF5e1Oj+9+OYWj8DN8S8
/h161CJy6XmLAbwz6IyLGTY2yB0hLMTxMwSnA849qZZcsQDvWVWodZYERKd7
ARt4k1zAmebh1lmj7ZQyKUIdTk3pqb6wIsHF3qTBrYpt4nAp2Xmiqc9vviF1
Wbc2/xeVzMYEbUERsVvi1mUYetj5glL8uk0RVDG2euQx63jeeL3hyg/1XxLF
fVg96G1VKcko36TUinePt3Tiu9NBgNOhmtcq31a3tdm3faTuMOhK0d+squMa
wdjckcC4Ba9rTfDwkfXbz7ZEQVcBegJ1JP1SoF1WMIZPQEP/PlzB8z9KrnMm
gSCVhfMSKE6Wm0+6L2JZM9ulOzdhYrmSl4O6AQxpax+FU0uk5I+yBYGH6iAR
dGO8n4biREx6FiB7jaeaQ0LOtPBCK4qqPOqXTixcqtbo8JFp2LGGy9EnXQvA
oRWzNmj9/gDLJEXwbxzcTyZTUBNCmcWgma6r4Qe7Id8mbKMgX7dzFC6Gc1iE
SAIOZ0QiswGEkzfennbbM1yelnMP4/29Uh3hDM5xw4wGiBGbsYudVxPnX1Uw
yFU8hqdtpPW0BBHeOQMsKdabA/3Tl1tQshMd+VVwMurmWafjdtXIXaclQXMT
lDYz7spdd1iQwoTTveZPSpWRXlwovXfz9uk++nj8fHi3+/3w0uS9dzio4khA
srQB9ACtiVgXANMYlsMzRvkF5S3xtoG7R+h49QTtkGP7RgcXr3UFbCHxBPtc
MnVnMjaSyb6cPe1tAk8KOtjKFa+GnSn3eQBoc3kWBva9qsC6yvl36+TNR4Dc
dLGOvDVtHSAQDXbHt/pUIdsu+Kq8Zu1n2azDtAW5P/SIm+Fd8XTRHtRgJ8n1
2T36xA73EtmHlrQ4A1lmuWFLitcTF4xYjULlmRJGZZ4FsXAcODvMPbLRvVhA
pNmCWiby3G2AzMvSdSEJu1GoVKNG51ohrQ1MIUcAsoCWn7IFANvwtD5P3xZ4
ISj/TgrRs5LpjwXoscgmb4hEWZBvIbfXfye0O1TZ516IhNjxVlsgU8DfO6PO
V3WdvhV6McTzcOZqX0sg7kUVSbWeDeL4O4m9mrnaH0e/5LkjHCAiCqHVh2fP
aT4AFZbKx1d+LN1/nnytQIgkYuCz5cj4H/pLf9ZME8tbCuQsf+0Kfwd73PAS
rK1XVnDYq7ShR62bxdsA9dr/dkJHsepsoU0GIwXZjfv5lkGXzE3Y/R10ngjg
A8pTXGrXuu8ppls78XkHjFszfll+oE12z1ob0/d9pHwnSCtQQXvj1TIn/BcJ
sXVFPOnZViP6TcxfWZK6JYsUXaV0WgNVLm81poBoXmM2uvft6LhSv0fUj3xF
65R1Fx8yGhxyMUZizSuDxtYGyaQRo2aO6TNaF/6QXisP839Ng9EIiS5Bk31o
R3OyIM9quXYQcTXCiM9JumSShGh88/F+jVGscQiiDuxVdHhYfB7DGgI7NWYU
daWOk0Txu1P2zsVqBYJuGhTI3vdkQHZE5AhGL8NDIQq3yUtJiC3FLPut6CED
eevvSWcXsSHvZah4lOPmPEkTjn9yZ7rFIjw/GEXRSdIerZNda+ZQJxSJgJGb
OEp4m1r3srDIsiK7w08UYRCWKnfH0dJD4hBmkKCN6643tUmMhEnkVnNcJ7yj
VoJ/qoq2fw4fgOs+x2zHD2ree+23TpV3npCWrPSI3QkNgtuNoUjzKpZEc8qE
e5ljEJZzx0Tf0VM+oAxkB6w6+uFUFGvLpDOLTMxNdsNGSp5qzUty7n7IMGyT
EKIb0jhmrTvKpq9gYBWr4ScMK/YBdUArt4F6/dDe7EEAPPlFOg5ZJCHtUIpT
/xx2ymqD1T/mr7HAx9GD6WwOn8nXrdTXLGAld1lrPwXGLXjcsPVDkk7+ZlYY
8msV8rujy078SjCVQ3aTx0+rphLMX7WSxCqx+8JJNIOhNH2CE4AZRy1OYcTZ
U+iEhvN8a6n4uP7Bn5Ye4doxrgX6MG9yHeKArps4tgnp0NKxWdY7KNZnAdW6
zxxRzX9BfHzIDkaiYhUScicNm7QqZRCLTgoHAuHtwarrTgqWpsrrGhk8EURI
kImquxqbTnHMsVRHmQXmn+FngBIOqydb9XYHStmDauk+8NDS4+D8RNy9kIx3
g7/FlWm7WOe6yXs/wOKlp1nLuJiDZ5zVTe6bT+lZup2HvD/kTyGGDq3AjFxy
k/KcUDOpzbWCMPTY3qdz7G898HMd6SrtQwbYvVr1LtW6BG+2otS+xftYpKpO
jxWsmM2kozBTSs0UUdZf0mQZW+JekRrb7LfSZEJ6m0NDdf5qsInJdN8m7Kj3
/IW8s4LBr8Y+J/pnGXvnd2evmsAMCQTEY+iac8XyYyTBIv0Pzi3GNnZcc8TQ
3hIh1yXBJ7EdYDVpZrIyiqV6Ced025eRjMnh8Az8+Rwg8F/mv7MwinD7HGET
qFvzbN+LDcgutMg3nbl8Ww92ZaNKqNYP942Dii0PUgCT4shngplMf+00shor
VEIegCHhJBRVns33kMuMcyG2yGsSjkTEmfC1mxW4T/eQPhxnEnEiCuscJCCz
j7FiqnLznGcBz3JFlKgjO1TPRSlGxA/s7yVIgQMcCsOr7mK9Eb3kOXdVBPTs
ltw1IrHZTo2DYqBygUDoTJiI0iH4qsZDW0juq4+Ya/IYOVG2MH6Pkbf/rXjO
araou4+Dd2oQB0/FhrPn+cOzYAkwvDTQjhk83f2C89A6wO9wd5orSOrZ6f4M
OVIsRISs4p/EDqiGPgseB67uBAdvSX8k3LoBzUjPYlY7wLMea0NEbGTu7ikW
ndGSci4qLbqVCTbtyMrywwme3+RBgKsC50LSqyrHIv3F3IWCc99XeMsXg+Z3
SuJH0hOSU2BMXW1uMAlKQ4gjqqMAzUJdtCmf8IBTTy++njNyHk60HbiMJ7R0
SD2Mc2df1p/cVFiI7FTGw2X26UeBmLoEc3RRurDFd2lDQjh7npJmavSPULnl
AgHHl4EJ5Fs/Z+MnKXvAAe1jDboWjTluBAQldYCwSxBNR/KRD7xoMnlSCJhx
DLWX4YOTTRWjsX9v9beL/WPEl/3pwtSRvTI1wX5CrBjhkRRknYOps6d6/4LX
iBwZQprCfCY7HpK9OI5ZyFPRYpIwiXpkR/dH4zQbVPlJwHLqgaeK3YnY2h1W
CLMTMqDpuvN5QeSDvVyb7DuUlBDCRctX7VvbTsGI2F/8N/03QsCVITA7gKVb
yOMIpJAzPWxYxcb/8FaUbcgifYSs9Vu+0yi0MWNfA9BTIhJpoFTiI2SmAHRI
4MgV4h5w8xRSb/pkGB1i7tv7wXURN9aM7JEFskvqGYNILxG1X3nsFgiCCM3k
Hqb/VVHixgEGeLUluE1afALSt4iXcLqzg8ezeKigtlVIJKCmVZNEcIH3UrpL
0kKdEqQa3Xg3TykoG3NbLj3L+uW4fRAZqPo5oLxel+CqVHV2gTC5uVbLXdEl
Cok8o2YndsiFAYlf7OuAsUmHMEqHVKAN1DSaoaVTRvPwINyHmxtDeEY/8w/M
Udnb2Iuk7Oea1LGwcPOX1RW8R0qiFbFL3G3doyLgXZRM4XZYZwixVWw826x3
ol2tg2jcEcoLaeT4QvL0KZI4KApKahVSHvFQPJZUyd4rym5yWzO1OYQWWt0X
6SAB2vvyH9iZ1DTfCEIO/h1Pc/vM9NFdUVQf92WNh9XVghbTDViwa8OkmPbZ
Hf4t/SVquPxBt4hJ+ZEDLQWGFpZ3HcN4PKB3y9xBcb2UIa4eefAWLEit/LEv
9uWJB1B9JshGhsSzy0JA+HfzTUaVFE6/wQ8JSz+TYJUrCnwI/UWr7hGFfXG2
Lo/kM/1VEU4Kg+dcZP5Qz3apO1++SYlq8gn8D4OmrEuP1UrIShE+zfl0w6xv
HTT63ORHXlWzUcoKeobKI+On0IkDvqQP8EUn+82OtfVAKMzMGHC8JGiKa7k0
7tReNHSOYdJdC3poNyQoUsJug8p0ioMFQWVYn/6n9FkYtVuV0i12PURPINln
miQTDnLcXwzTml6YT2/TQ2ZKn9ZGA9Dgyxz/TZcEUzNTEc0s+v1ksmtnd2ZO
Q0hwINTQNT6vf1H6KuJHK9uMhBVYDd9jGEcd2jYNG0iP76rArXSxBpgr+COD
tG9P6eeRTYQfD8u9HMfsR7EPW8tvcnzNkhl0Cae8cDgb6XZymNhFWxBs6/Oo
4Efsi95K71QJwxSQqzjXYq3pqnU5Gs2Fle9ozLPehV9kLVPjj0SQbWdOeAir
BiKSyuT3cNwQU08UF5xuvtzDlRHrT4w9OE55ZDpqYAVWmKHMd1X65XQqJsL+
vBrrZAZt6s7lvMAF55K35gM9kdr8XopYJvHVuxthroNnEn7RhmxSZNJ2bDgh
3CLxnXsZnzDvcQJxf7IGkL8bBAVvpUKxjbzxLqs54h9mpLwtiivP1qPr3NhG
a++j3BiRP7jVg6q6tOFiZPyfQW0X8CXOBmwUgEMHkZ7uC0HARn7yU3O8VDIi
BuSKTJ+sMgeBMzG9EpLggN0M57AWAxs/Xun1MqdwmIp9XvO7flq4AZtLjBCD
m6vWIbO7jqRgumiUOVXUuInK4lUnTVelFi6tWZO+2Plr7t8JrSsqkfKBW8bd
uuIkOOD6gaR0uKspRyhDIMDtFy27hQ7ZfEcBDSHPJN8vGGWMa6wLLBKZKVt7
AE6Twlxq4A2mwpW0ZcYi+lxyqQvo12l77mzAA+yuQUyRqb3XTwBgKm0p86uL
I16Vy2OB4NrgFUsykDEMb/bie6DKdA/kkpw4kg30MdHp2EUf3WwuMNp/xMpC
KZ2YBjSuSfD8vNK+gkV2xvLudh3V4Th7mjSlt0ugKWmqtms9G8TfO58qFr0w
IDgnxuVEqMbZzivAqNp3y4CrC6WBNRAEHktdbstE2pVQOxFmfgx7Q8oHY8pE
PiSMW6w4KHJspzzDzc5nvQW8m2bndI8xuvIO5KBZ8RC1UJiSRQnSXUPYV7WP
kuzlJ3Oi5C69ELp9mCM9wu/0bs/LgKdZ7EgfYn1tgniu88ZsMaMWScpGhxfr
/n5nvXxU3I3cZ8G2701vOpktnnd9iycU5SWzYQESB6DVWbsiBWbZYum23PX6
3LpGyxKatHVvUJSb09SpfxapZurwSdGElmzvXh13qcX1qJH+8OnVLG5+7/k+
DcFeOD7aZsgC5/Y2DD49dDCWYv8ZCJ3p0U5OgKQZZrL776OBVlEhCZE2HDuk
BXOn4JRZbnmOKwB62QMc1TCpCAtf7oamMHSawjDg8z3g5PaflW2cpcvaPoUn
ShsKUGmmNk9E3x2IYXB0nXBGuUuAL9YbiVLqnNKmk0Ni9/dgtrgqPdt1ncrc
i5XhhmPD0CGSLVAo0Y/Q8i9b5541/CMSGexOtIUB82bdSD4H73ZfjqUH9nYu
xC3akSWDGS3aS0I9+ny31p0cTWxr0O+Go+6k3FbHx2bfn6h74q+u5YpvLtW2
9dgl8Fqhkm4uuhMXAXuhL66Dn3bEhqaMj+Cxzp+zsV/OWSr4fXybiLlN0r0O
JaXaS3ANpkkuzYgJWf2zl7bmktZ/B1VWrA+2+TGckQPM6Dc3dUTu6Vm6ckza
Ll/7u76mGg8uk4T1evuCBhz0PBaUpNXO7SPTIyPYelTexjNw3RqmadpgOKzP
rBSv8eo1RFWi4sgeom/saZRB8hAri0u3s+kzqjaP4MP9yu/Nxtu5fY2nX5oI
QaDEGX35eXUEMH76p7T5h2W7BhgmbN7A7VF8qFBIu4tp2nCRQg7J1qmg/hHS
4sJVhDBuwhJ0pCMUo7WjGZMINRY+5Y7Hgp00czhrZ2DTUoDkithg5w8Ok0It
Jwt97SIIVF4t6NQt7yWdvPY8Kd0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzdw2HovOzdHtUadq7WAyzWAZyRMpEact6aUukDvnBkFZaj4Dudx8p9ZjfAbKpnQ4ZDLsu6GEygGQegk//ndTmcOauvu8P05nipI3T7U0YMUnKSorTdHi3OyCo0uA2cg+q8ZaJzK8dwN3g5Blr4jESBVFiRN/f1so40oJxZVxAUNkvxm/ssROh67aoP6aLQFL6kBZkyCdzG0UFpREepCjCdF79gnNIi14w5e4RrzgW33eJjTHVfjBtQCrK0nLVDNbDoXXhTcF7jPaoS7VC1B1Ru6EVBJbfYnHZ9Y9IoAmo0Cg6+J8DzCAiVlmdFD1WdRu0mvo4cf4nLxH5894IPF1SXJ43qy9A++kjRz6FbLZvDRVqfc9D3eBVY9iIMRUUWKdN361z3kd/6LN8X6wr52AywNyOST3GUs0gC94+PwjkYBFs5o7tYjIIJXuAiiB64Nr0DB2IhmhOMftpnBBIayKfxBaPP81fstQUPzHorU5n6G6QN798bFmMfqhJ0ORKg4PZaNQbXm+JetsdjRE0Qo7Apexs2By/vwJqlBCUBJDtw+dyJTfly9XImNw13B4vIcGyejN43ajv0OqsUp6glcYMKH50+bjiCb80x+JDYmSFrvPg4obg0IzTWV9msh6pIXsPYd3M7ef/ZJ0PjNLZ0TJvA7y1VaLcmZtv40DFT+DkmLHK43bqcjRdqBAKBbAgW5182uSAj7QCDsl946UqF+MtJi9wNXKnysw9L8y+YgDWhQEUJfgck8lskFh9+I2A9pO+Ujy14h7sNoc3Q+vc7JJnAj"
`endif