// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wxYBGMrBXdFfqlCv9VDJtU0KKlIA3RMIjdbKVjd4ikS0h9FKrzNqRijWtI4l
SbBlkWZe/5chavUUk8FqE7gCcXxjt84gdb6APTxHPU7Myo/LoEpbX/TnWnlx
UdtK7cRRke8yOn8lB4mZiVbtG8ZTbtCOKITvKJD0v6GwDYncxhnmXfj/eDML
687BFWikEn0ubaJdZXd0SwALTmJrPQ6jNDXlkMsV5oGQqYwqTfJ3EDJU5Myf
ZJSbJt5o9vqf0TUO3w7u2JTxP/CMuIyWC3j4qV/Aau/YEr6I77K3/5x4ReRx
Lv2XdOTXopWsOvrEqpgmBZ3L4ty47q5LH2S9JBzWKg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kSFcE7boqReoqlvujpphmtVxqOIFfzooDlk/JScMzcq1BNOEoUPcKRbvILjV
2a/XwUZ3CI2GmCFGhomlBZbinnWcVUimpERfPIFB7Mm4ZiMSP0SZ1VSvMOih
bUtUYVjGTr9qy6S5spNah/DRThbjQVzeOve+1XCRLRaVvNTfZJ76BHNTEk2H
FnrWfYBrAYqLBlE4ztO/s9kQBryH7nQumX4TM6ekcX18CZQouTHCbuUeC483
q3pqH0fWLqgT+OmgaQbZQEVcdqUlmEH2gBP0KIFe8yNYW9JqeNCjjkT7r70d
BrcBQDfq1Q6qQsEyO/iUgdSuUEWlu9rBopWhNldhXw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
et/Z8sioKDfKUCkVHALUW+Pb+saJ0vCB3GXcMtEvE4362IV/t0ZsX5pKo9QC
Bs+emQDNX9SkHW70JlmwNym8pZxfAjWWrdAwRgtI14tGqgTLRo2/tp2fAR/I
KK4/qtgaFVZfJMfKBgM17Q63+w8xWlcNWlFfHy/av1+p7HA0RuxEB35Q7Yet
io/azrW23PHvmjtGr0W4y0ko+w8ZaUQlz8lC4aC2Tb0+As8xc9quUy3GIY8X
MnFzrSmFmBaPdqviVft+jYF3iW8tLtXOGz5t0JIwPbykLKlduMzbxQCJjHMN
k0zNGfjsSBcYLMhVirI3jsM/I8c8W3DVKCz8L2aboQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PeOF0AtvN1wtK47808rfEOftrlb0+5o6aqRtWhCTP4PbzqupZTt7q89mYPiF
fX6vY8qiySo/EUDwp1qZLFc82ZArUzsfGspgvGiJHcrOpSRlYUapsJiuM41M
3ohoDo8LCmFSq0Wl5e3Ir+G4HULWJt8gOSfyv5WCLLULCfcwHqpTsZd6gB2Z
hF7tVIGXVu7cfhseMGK3cbPhPYBZYcUuAMnMu+ard1z4S4QwrtZSu3qnwNEJ
EBK6ZHPXnrTnBWwdWr5Bn+dQBhQvSKplCp7kG6J253FARnjaxoeC0L6+kN5H
hp7JEzn5q297zcGMVqe8wLNiLox3ufs+IJUMwCP8Jw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hOPZD9X6OX4h4+NOvhvdFCZs1B1drC2MpcRNAbs0P6YOEROlytI+e0d74ToM
ryoC47PnM52bbkUJjG34f8iyWkXz97w90AuZYNw7N3Gus6SB/duQ4dm3jRwy
uDtGNouRyBapb2XCSIstK1y0Fe7Ca2YbMktMQLzl2RlEf7IgWjE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cOGEZ1lwYaLFIWh2OB5Q1xiRbOXs2nFOr3p1ru8/oWDQJXmtraTfYM08T/zC
Oeret+HrFye9NgAwDN7zFWaPt5p7p+2Go1jLfTNzf3CGajNgPAZ7wHRNwPam
r1UCEUBtqk5JQiUyLZXJO+s6DLZn05wswdz1s7gPTOHKTywSJ+5jJZjLmk3O
mkfhY4udIov4Qo+JtEw7ux6r5i/jbieuSADa57o7ceNeC0M3uq7krpVOEM3C
d/R3wEVt5mqtDEMIEnd0bQ7qWr5NjgkBqngx4nCfCntril8aXyjxy+oUZSpA
yXYPRTwUfJXd35mprw+Vv5p4Qq0JLQpxZoj6pNTqivVUrCYwY2DQhRiaseE+
DKJgJLj0zlYD3mnceBS5kHxJFNhhUHJhCsXul0pNR0L2xm53DB4PNEwBxCLS
A0EB142DbSzLypsHiiLwjoHRBfKjI64wvCqM+W3+yU4Zb80FFO6pupnnHmA9
WlkdarEL1pCbT9BiN8/FEI8XDSvd2Ew7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VBWvYUyKWRRwhnkcV2FuiwHjq2Y7kLBBC6sa1A5tDVXFsgbCreGNaF5hcf4s
rPdqOSBKE5QZDAdGvtLAcA5kwc/OylgDkwLLIIjeYduLvgvHjhZY3aZRxWlI
DcAWRnYUA7P28yfcyMAnV5yrjkcrqPCIAMLf2FweUs10nghn49E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hvjhN0WZ8lAx7xmX1L69k//5K2NAEKd8N5c+Bo/plE8v5od78uNKkafWjEOg
VpGiCtoZcpDQViONfX+CJFyWUIec1Hv8tZYgqdUa54hc8b3H5pgahc3P2vh3
ZROSJpY7TxcPkpkW5xeIF6+UaRbEXfYt+LTeGKCD+YIb3p4MIZU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2576)
`pragma protect data_block
adJgpQaqj9LCluS0JjCjTtbXGTEda+TjAfY4HErEY25n9VBsCfabZzfbrMYA
WO9HD0kiIuvI4ipkR2LPMrdZm1V+bd5DEnk6USLj73GPWh7Ou+zaGGQaoBVS
LbflLfaf04VsCjRTvozIM1h8YDQbBUBs+1My2lYToylpApW0F44uHhZLwPKY
reOrPemEZ9ebAfpbiB8IXDaIj84c/H7VBsVzsrXQghcl0Y2wagr+97e8xBD8
JL0URPnbK1FkZdrOcz7cuN2BlMXxtw4whYsEg2sxGRKdMvDzuOiE1oI+Y9Fj
V1opt8ivQxDA7cwrNd0mOPyCP+U5IZauxQMniIiz66oYtxyqzGVfYWxoHTXT
Rfapa6JpM1LVtJgCWQYz8Onfj8wBUNHUngGXARQxLgtDDFgv5ICBnzVSpP6M
XrvmoNXj5o3BCh1iOwgOiHwWmUsEAF3Hqfk6do2cSjT5d+22FYbzodM0FEJv
SYRirov2vwHZyB3sIaPYFyI0rLlXuHBKWq252P5Ei6vo/iHQrJ0hTl50VEi4
jl5Z4A6hF/FVKorZMbrWgNr5GpdneLMLOJHnlysv/4CeburXnoHayVPTmZse
sS8OCTKeftgp0942lWKTnyuaEvfaw9Q5qiGTTNSXcBRSuRrsnfkNH7t4z+5r
hSQbHsRGKziBVbFO0TcDC2AkEKbW2W2TXFciqvVmyrrSwV5YPciiAcScMACk
UEnBefXW3ig6CXTTIxVZQrPjhribS+dZzlCQL1zzA9rKvcVgLbGZlKSMH9Y0
LtQc1a3Npg91BjISLb3Ih0mE57IrvduEJ6aKAVV9cq3bTNcic2M11BDN9MYG
SUmucxTed1ThM0+2xJUbhx2Cs0l7b5GuX1VlNCLOZw5D9iiMBTmYtc39znnL
YZNhWQu0dQx3obD1JLSXsqeMW58+oCFqzV1ru06E2uwi5DP/srzhCgpQqLd3
Kx+4uOio9GGP0WPU6Q8lfah7XAk4h394LS4DhQDVKXPu50B7wEet/JfD6L83
yZNzsKgemJ3lGS//WS3KaCc0LukgiWaybDHoFt/XMQtX/OXaNxsD4cqXWrQ4
e2U25ozAbIqN+ZY9Jr8M9sM59Z3uO43O5t4/yaaHkO7eyKum58EToT5z5g76
CSApgvUUVhOtSN0p9kimNhghD6PYVH9/nZpo8dF7y+25PCH3J2a+bBLH93EZ
rjlTyKQ3Lzx4O1ccwS10QvsHTPC4Qy0lasENzOuK+rcettas8/ELoRxw1Axx
MEfpfdmiCjBQe+lbWeA14XK24FTzt3v6Gh6l8jEjdXxSIwKqjFE6aqjEsPVw
G/gJ1rMu0rvCshSpNfY9DD1V9mncclzerw4oQqxBbK2BxxqQMFwICbj3pBC5
TQ7VIOFRASF8x0oJHm/FmMT8/TKOzL2iUWZbQtSQ04r8efqhmUAwwJc6FJMm
+7fPIcOeKRGQNFxSjePoc9FwrHS2w0+/1LfuXEd8w9LrduCrrec9f/yM6jSO
/FEsaWgsBAhcSXvhD8wH3jAPsuIIyUXXoX1LgFeuj6Mg+pRlbmA5BLuz8CNh
1nildUaiQNXSliSIo+cYQA12k974aA7mjjtKjMvasMlB33EWPopnqgco0URJ
GcfWh4DMixbB/3pteDOqAC8cEzh4tMhA0n2OzqbNccN20dw62f6A4dcx0NM1
uB+c2zpyM1/rb0Ffks0mrN7MwiS0yZNeOdO7iNfY9Y0ZEpmFcfQ+oIvr2Zo/
ip4Oad2N66PlWozh9lf2DuwcZJ7G7oy3tt5ytwYJWx2iKq+dRycUrxvqauFj
jySJaQuNDKg6aiIih0nhzqSqTEf2HFctOFrOVLJwapr5pebZTafR1pMVsdtN
gBVhL+psT/X8Tt4Mqzon3NkzPJdHUU1m6qDIvw4ujpmdb4zBW1EMNtvGnXRS
bNJR4xwq2ymqnWgborETEVxK6CRuoaDzZtYqjI/wWNkGzb9e3jefjVPAOrVE
/F/2MYhgChsjdJDUR3WBK6k7NLMV+5E6iZ7/Rw7y71IOsyOdsdy7Qe+E7/28
ssAeTtSv5DIeWAKJxqPNBHdWgtfb1wKBP4mRmkSfBKO5D01q9PY54KKYon72
Eav1WXUMqZXH2t/FX02kRSFPdI9DTQXdPbeN/NxWDzkfHxS+Ke633bklmaF+
BHoT6KmPqEeLrKvOioKxHg/oquBUBjp50KI7JouM1y2kCYtzJiWPTVKUVuIg
68V1nGENHKZtPI4+mQlvzNkVpmhoPE22eIcLlDS+PBe0FmAlS/ikpWnAfsiu
6NxUEycefpOXxxM2C62fqVJku1OFk6/F7e7NaAOfgWzV5R5fxVQjhCtPwLTz
AOjdLJYA7eI9vI9r8+Az7rdjz+O5Be+GhT7SoMgpuu1Z/1c4f8K/wwzMdlOW
eQeYQuTQMRF3NTB8jK9C/8HfKgMS2DO3P2x8hSc17ikLMGXrDyEtTnrQ386R
K3SPjFXCkuBJSe0BSHBy76mOOKuHSbzsJ26C2NXJ0ie7AGBMpd2jDc5IzYmK
I7yxsXp8VFmvzC+6iaJ5/RaVaMtIjlJ6Skw5iulMB6pnQ9OV2ZBkThbdrFFm
fkAMXb6Wf8J2SF2itvFHybESDyhFYEIICc2fhJgiFifXpwm1pctvOv6k5Zpd
JBrnzSrPhOuuzdqQpW+WP+KYBJPESQsbF/7Vh+vh7F5ntS4fwbH1QreWBkU2
7tHmLfy5/VDL4ZVZ+QyEpaX/L5f8fwII4Eewpq7kWWnzfcWvBsjiFjTpgt0D
rE/jBnDpJbmoK+uwwpV0U8OCGNVrGlYuNPbCO/qG8wK7TM3NyoVEJLKLR7yk
kATvmMv3OqDSIX1RX0MnLrLr5sqiJK6mRYQayIUEC7G6mfWt1o8HM1SDyThr
/Es8V5hZ7IXm6tahqMCdnZo30DeByXA6bkXesBD08+o+8j4qAvOtPTGQk6Or
WYZNWkYKf+W5OyBNmi/ndR5lsIRo2P6pBZEy4gl2wLta1c7sVbqIZaYcC22H
9ABVKfJyp8nt9PyiXF7oYkmx0hQq5wtyZMj3dnVj0E8yVA45RRAfDdRqYSm4
0qhRTMowaCNC5szi0GKvVqPEClCoVcouf8Jkap0NaTdInBn7HqN96xOc7jYK
x7Zrn0sxjp/oI2fc9xsr566/bjQ3bOMKUPSvBxQc7a/nniCnhKIgEO8ek17O
Dx3I23UYjVrP2YBpe4/YfCX1Fpgx40/+x1JeHOlCNVH5I4bdJ6yBSaTlGRIV
hrv7dkEA9NRtOMBqhu2Y5akqF1NmzMGW3FlsUGRCkj92Nb7aEkMw1vG+MRm8
XmX0YxOaq1fGKz1CZEotQ0RCMXGl44T/sgt0YlB/VFxbnTfQc5jZLLGPyEz8
NtqxWvfGSyVeLdD2X07lS4FVEoFeUbzOWn9dAhDduNAKer8QYGRj7KBIv5wO
rZ6Bz2vFbZP8Bjw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1J97/sKukCNVLV/hLPBEXkV/+2S8WM03QsmlIVq7LnsndCE/LbMp77D9Ho92lDqv2VKEG019Z9QZVoyKeeWJLaz1DfPw2oRkHAA+fFygsBm/POKJqZ4toB/KkH3byUPMH5NhywnkaOlGIoU1thYWJxlPR3/1HwxonViHNuuVUdYz1TcmghWw4KgwoRxo3MNQuL9uWWebxud0Epsq12GdDQITgX3CVG+meomu8VA+1TAQoFspI/fz2cFIoYMcxFJzd3HhcmmT1sVOZEhOPmHVfu8tfnB3iA32Lb5Tweq0jDl52gKn7BvY18qSr/X7xz5+pQMd/q1JQKH5rmYL1WujmX0Hr2G+U/xO+NIBeTdl4A8oFf0MBIKaWLL4y20NyFhwcdBpO9O/KnYARTFrZvShToDucTa5Uco2+2MmqKBnMtRaAZeaDXWMhLib8KWMhn32SjF/+ILDmhp+H907YljWkG2SAWLyHvFlBUjuaCBKvTEdmMACyNEWBjRCGdtNH3JQzlWdYgBKgYpzOK7PkxSZQBs3s4VCl+QQ4yVJ5S36MZP7EwX3xk/R0wHbq7sqs0fqCVmnqH5/uOMSznfftSShmXWgE5EQcVPlEBRh0uUmJnAm2uc0qjIeHKhFOjt1hG44+F2izVyrgHLE6XLpqtrCjmknpRqsuayuIZdepVjPLifVTInluXjC2kXWc3sbzDxpKgxUMDEIoE2tR2D5bZX/lakFwyRoYouFFEhyQFJH/W1UcPEVC/rnHIBrRBZrQaAZLYNtfJN+//3uJZXeebyoGyd"
`endif