// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DL5s9BWXrHKOUx1xADzt/fOfek6yIbg27auGvEEEfYL2iH23c9n7hrK5CbRc
N4vYC1UUS1Mla4ygSqHsFMs+s8B/OsFIYA+n4A7swqBsGan1n797WIKWH9PT
BRiDxFzgVjz87SGXoccggTIDWYDX3HyGhCFcNrpPLGqm1XFnGP7hHkfXWLfk
KmS7naNS6OOOHNLYvJdndtY7ZY9Qrw2gPMSIx4BpqHK5ToDoTqn3HwfZ4sKn
mEHcgz/pH25ImDExLVTVPSnTmHBCw4k4AW9s+AhHDb8hXKZkaXfSLY/lzQbc
5g7LzozdUgXpgoTC6u7jwUBouxqk8EQkRwjBPb6PtA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CJ5WYMcqOpW2UqS+HFXwVPKslOAQo6f+/AePSvvF0/ZSuRYehz/cjI3rwxaV
5K7RWzHHzACCFe/X1J+B5hWYwsNqn4N5prWLG3dhsaLQGvnO+vqbv8q4WFNW
Nt6AQ2EhVTRS+XzrbkY1M7fTckMUeHjxLVJQvr/nQ0NcoadDObqZcrdVXrJu
sf09RKRRcGi4W6/Gn/Vvo6ae2I46dgdNfT6w7L64VLYSt+oBwhjaFnAzC1y2
k6SRk6s5BWVG9zljgoe9xzyalJRzMRh96IqXps7w5u2E/E5mO86OHpk3Z8A/
h0xV8WjWKkWenEKBhQg0Qrtg2H1ueV+EayBfH9831Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
t93ORgv0rpheCd+7gNEpqpdWLox5XfBvZxgMr8evmfkdOuaqwPSmIfIORNRX
3bYkIhETHZcmJa2P7dsQ7X1FPQ/tMqISbreElxqWc+rJEZ6atM8omUSrIr29
D9cSisG/BWaJrvTMDNGsm/oTkbBDewSRUn86nABJCWFC04Hu8dMID7UDbCbS
nox1nzwj3pP6PISCZmS0ry6VbVqHN4bX05yCRM1emT9j25fvXOZnvRxQ+iU2
H0tMvXikkyGgpdA9ILx060i/RU9aBZXAoUDtku84yoGuFsRerATkYgwi/qVM
tSXWKgGU85IwNkZZ96dwqQv4nwF4g0xduaI+hVd5FA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rMj+7Vvh9H/vXiFbIVTICw8n/W78Ps6EikHXbMxhEut8Q4htmvUQeYEc/1w9
d1hIVRBFs+5fky2jgcfYfeMXUdS8uC4hE49RVW7WtWuDNcg/iP9kRQHZo5Kw
p5iQxuLGs9zo3hCSq2wNJO61CAcSb56ZERaC34418XA2BiBl7XQP+Dvd2/GQ
S2/tLYmfay1HaaS1EUtlfgtTMXGwAZG0uzLWo/y2Yx5O7bxDKUrkpk5ewRuf
ez/YrJCBDMo88qT1zkN748lMOHg23YzZCuR7qRYCUFcH7zjYNX2RixWLLFtx
YYq+Rf6TFCNojH46NaGiK8vNx739bEp4SE4IueTVug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SreMTjglz97GR8hiCj+wYQ7UAcgmKl644GwqNkhCAJMc7gIgAF0jj+DZyeK5
JEdzgQlo8Y7IuSMtuKS5bJK19j1JB9H/fJH4oVoLlOfzrutjG7gXGNlUjwyr
VbZ1CPl3bfRCo8VcDw3va08a9yyyOJTrJmvxlxR2MOnUVi/cnqY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WiVx7ikaycQ7yovcgN2momUHFjlH/aUJffgbVNKwSsnB/8vAxQhfxz7NldeA
DbNZjB4/0DhJgRNUfn8LNBynBrmg8VfaZ6kI2Vo8YQHLb2XlvHjukNuIdagL
uioGaiRY3m91EaXgrT6ZnG1zQ3LfWtYXrWPrcVwJpV7KI0NbWOb4GyF/TTHZ
aj+pQn6BqyoP0bR9yMrc+NY6zOzgb/hy2DPvuBoRyFufz/BeMbxaI/XtZFq7
gOE4TJ+us+uSPwK4lH1jrzKIcREIGiS0rRX5ykfMUTeTHAVEULlqOoXTvm1f
wcZQfnH/8iOD3taR2oZiRbGeGrFd8YvE9Jz/McgDsJHtq8OO6QBO70EiVd72
lAVCZZJjEfqsERVflJzyk7sqlR/PM9wIkcFIkX3+64q0op4TxHX57C69ksD6
UVuGu4gLlGsV9AhgPEAcxy+FY7r6r+oRLFxnkrVLqbM9zwLCzXM4TKu+zwuO
agiEzoHI1lgtgkszNEbR+biYNKh0Q0AX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Sw+/sUgpy0K/auTY2kWdfUcGDXuaRjatapwLu/yeUe6xc/a1dKOYztQN68W0
q18Jqa1str/8IlcrPm+iK5AVRf2BvLPBY1m0ErXer/p3an865Ir3qo3/Arc/
Sfebh7b8RLKPrDOkqQdfw3ERsGMotABPoNT6myBGeoEitm2ov7E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
US2BkXwc6rlJkMbK4nmCYVwaJ/uNri2dizDN6ikdPPZwtY8b/zaA6spdDgKG
2xTGTXuu8nOkQuZ3yTXFsctsoYwlm96mw0fpjqvAJSCxUbhUkPjcup0jfyWk
MWaoKiJEnDD/2qET2oahCY3hpLsj+bQy5sGdQRzWIOC5qjNczRw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
WOUB0yMV7oJmzzgZJ2FPZy3ybTs6CB66NBczoXG8K8d3GuBFwKTP5cpAArTf
DnXZI2p5/zJc+x0gaUp8jmmNaYoKOFVBbpfRKIcq3E4PQ8z80stgVkmUW4IB
M3SPLpf2hd0uvnHLzpgcAku+0ovCAGiTOACOP4CBMyVHOXrVhN/hAT9/ivYm
x0N628sjlXhnU/ylY5PCJr+I5EZXhEmRpQE3kkJaz32e3dxCAu1SPa8l1MTI
WRZwtKPeWTVoldLC2V/P9EC6jPAGTwq6fVyJX5lAgG8mrHI36w8m/DcfTROg
iORsSxQJXAdOv1pDScO+NbozMA9/toPSe0S+3C286zT6KR3OGKmwA0hEAIi7
dLzSLTt4noJ7r0Gy26WwuDL1lc5Lj0MLJMEgMy+Sgmc526EDxyRHJXtTVQkM
KzKh2g74iuK8U+XIOIQRAw8yZsdgelH241TQlhtkrJQe81sKZg/0Eja8kNLq
nthLfHgRQc6OEjaA9ByVPphw2MVxk3oX208MYDP8A3c1b9qrKPGpHfgKDMH2
AiUygQkZV0/ZWfgTNKRp9Gvm3p06+wcNgY2PFJRx0wqWoIIwC06uxzIjMH7Q
Gynm+Y/BHNbgsDpPpCWPQC9/Ox2Bc4hOKLuqxvjoj5p0cSy2UYw6NReSB1oO
4Gh0wr8WQHelaTNYWIyW0OYLD+AfpKxN9yDECC17jEOR9E6AbGeyvHKchFPu
EYPzHIJ5PS9oi91vCSgnwiHItbj+w2iwP1ZG6bi3bBRtN50Ai0x66KtVV4pL
7lPLiQ7hYGrkGQ7NdsEUji6OJ/cIpv1DpFx3kx2CgTXTkmhu/NOGN9TGbFHC
QXy30wYdsXnYH2r5OOBSpGSxJRqcW84aWritZVSAVL7HILuqwmKLL6vOZngu
mMhgynGrzLlJPG7DmUWaDbGIcBRy87Bqiibal0sUT/qqcPG4m0qsl7XQNxxm
J630a0pxu6ZCpm9RjLefocgHZQeH0qBBDYIMRUd0X4FdA8kTMlRz9l+1XbZO
yQA4co9IZZAH2KDz4uEbTmcclklrfbuC4joNaEdLny6G73mcRFS+w53nX7tU
hL3hpA1gEoT7XrhBR/ryNhiUjujxXgmI6MFK3V/CjlBGwvxK2ExFZdch2aU4
SSCD8msTp+4SQo5wt5dw4CbVDkZCyklxORTFPiIe/bj6JCNFPqRx6IiT6AGI
6A/n7foOAWr9/3uBZIQQA/CZ8OnnLm7HEB6tPOEwZwYeLv1B9+g3zuv+8tWO
HVlQK82I/IA11BuX4NnttVER5kG2spLCHIEOGik3NOejByYZYR0pT4kErRvi
c6iyyEqn55dbrzvikKlfm3yZDUTumTXmPdu2eeflN0xQYck5WD1qhdrYTRSL
P3Tn2hUzsmPfTus6+Mo3CvRi7aj56oeoIBK1RkSu/0iElpeTYALe0uSnOr4D
0k1/ny9DRTN2xH+IbUEygLHpKS+qh+o063oczrk1HHxlxiKNqLDzqK+ejPNe
J+i3iOowT7H4IyDQIwElNjvTqM1wMbB5Jk8UKB/kZaopXszZvUevst7lm/LW
LAAe0gjC4lGaOmhM2zHZf9QOUdCL9Gw87rmbaBsGITbHFB/m9k4Mx0u6Pwrj
IiMGYgqclONuzLqex9nptJ8+S1WGUIVOxlNgiZKTPO22ZBgLvvl+wuTHNzMA
g/iAf1eRYkSE7MvjdOHN+dy8CoTae0AA+n23A4rdT4M0+YKE3Rkhr5Tu6TyV
VYjGR22+IMlkXz9eQDP4CjFZgD0wMpZP/81Z48ExCGAnVUlTPRFwwvfl+HQr
C+Q9ppMff4baN4VINtnGOY+mEa3ShuAHP1X4T8Pgup02NA3aIBQsC3IwY68u
0vDdJIv/30ZpCYfSDbWqZDNGK7UQ8V/gxssKKDRrV5lJlW50fLZU/AMvw/23
Gm+CbqMQZXWNgkyvTFdOKz6S6NkS31jLTP23ZGtqKEGdfFQ4HAc6Q7eC7I1C
7TvSNkezEMC5ejH+KDROTg2bjjpoyXSe5zs9icpCW9cbu900VlcjoNdlU6xD
DouevQShtXU+0pu0h8ezzvX+yxZ3504GOsJ8wq1zGG4flSIX0ao+Q7TTAso3
j3A9VfjmsrVYvjOYKkeFdZtyEX6owv1cuQhSfoC9Qp0EJKUAH0vfcXQz+p1D
Su7bNgYiERaQiQL/yY8In2ct4y/e6q2BE8hZ766UO9guuzaW27fWcvPC7IrU
OIgtOe7JLWmJWenL1sy8qkpP2mi8ZChPhuEvC1dhVHfDT3beAhRjjFF3vulB
NNeRgtoaV4HUQmFMaeYnPAo8IgR93agCwIQikE9TOzzwuJ+jrzHOBNsxKKYU
VRhl1kBH5uUGzsNSYodEKk61nMb2UXOQVnApNIZMLnxNXfhsBMs0czp8K8f0
K8m1fYIeolJLcsD0WBTznsgmU4lbT+O+BbB/Uxd5dCVBJ3+EbmDSErCqYTHz
ouHSWYxJLVoBycNPdOXIYrhoHc7YiVvNOIS9JkJY3/FEKudzGPf+qde2Q5Js
XCOe0D+MG9Lv3URFxfCBMW0BBfQ6CCzHRt6Tsyuy7rDQK5+Qj969v5l1CqdQ
2QQ+/BU6UMDkz8qOlIgrfpX9Tqq814K/M3yk9nJ8sY5l4DG9IYg/fwKOJLiT
pBRbN84xAS5HWlzMijQd0ElU5dt76szek6usCmPUfeWPFt1sPVr9F+Pr0LJQ
j04Vrs0yK8UpPEvUUexyJbc3v2NQ2wV4BVHNHg81keSYNluZBMZZ2Q8g6Y/N
/tPEV4oLxWWfKBmSkq0AaRIkXH4M+/cQfZGYNkSy0s8XVdS5jlPYXR72kyAN
hLDa9n8cU31XgQxjsgP4M1kaSNbEWtjGSWBRAdAuOo6V28r4GEtzwAPY6EGJ
EJBvGDoRSyrx9HUCqNELaAhiAgjnKi9PfDGiR/6pHWBW5FPo7lzWVsKPhCgA
z2ZiFssRrYLs5uAfS4ypdVjmAD2abS/USY3YYNRTMUsRnGMzUrutnuHONQ4s
WcX1k0NrlKhchxiEiT+PIkUaAHLkjC9n0uWddPhZIxJxM4eNbbr4d8xcMRYv
T/UF4Wd8d056libyBqkLb1y0bnrK80s2ckqB3jLQdhqY65TEQbvIWNh1QV8x
HrtshE0ax1sER/3H5lE2pVW9Hsgp1HR0UvAQTIdTS2XZxkmIJ5QjuD2UbZkc
Rul5hIjwN/hB13X0UqHMu7yesuYnB4Y6qNetCZwjldj38LAtB5fm6b9/975z
iGJtrCimDcjW+q3lae9qURrsSok5ig1MzA2acHRz0pxcbjsAOZcrl05xfLg5
bVPxd/UZnY+1nvCsuzm667qk8URNvng+B6S/V5nFkTncZ98YO+FCAEU+qO5g
oy0CnMv/wG0nWtij6qOKVhk64+6gi27cjUSb8QmbvRvaAVRx/xkz9t9btP8X
/apbjfwi6iCicxwP6eabYT6eb4LWZXUuUI6viM5rI5xmuH+V6DpSRrF47LP0
1yPsChVvYcJGO/hpYSp8Bd8+Imo4XuwRW1OVdALK8rYYjGGJhSxAdy7WBlDk
MWl85Z8hDjJYE2Am3R4Vicr2I3qg1p7QflFFSI3yMhBAIduUgn4O8dQgDYGQ
H0KgkZrF5LkyhioCM8/00akmlgOrVV1klwSwzIUYlXjPT4lU0GpeVz3PdCVT
lG1MqNof0a0Gew3X+QVnfa0BJ9ut6JaiwH1bsfiFFPQ3Q5F9SPLCy56ltibU
YMbGSzJPUu9xeIHd9Lvo0sHzHkW17s56iNgJn0ufkyoh72Nh9SFumpdftqUo
ilRbTV80rzrL5EyviqIX5hmcowoYLZjCi7omqptrcMAjmat/kTHqtFgHMBDL
5fgxeC67g0jXq2HK/yU65EhVsz1SHXQ5jXCjAP5ZWKQK+ZZzJJtcp2aw/jqV
O9YGNB3JXiGmXzG9wUeybmkxgQQsR0t8C8nAE5wTg4jlqLIqj0XxP7LCrzES
ErSy3pYCZyUYLlYLhCwYFfwwrT+EtkhDHhDysbGoUXQ2mt/aPyyu/p4WNe46
T8mEcdd3FQw674DYlqar9CUGlQiYO/atlA1wZ0ZbSVZiEvOld+DP/shqu/9w
v0LTmfKQzvIGRle4gkBhIohtrWqNm9P4d9ScCSJaaFPdeYksEHqwQWcPloH+
CGu/JqBaGXX5BTPPZYhja1ePDQF0/VPjG1Z9FATslTT9RUhb0yPYhy/gHLcn
flVTmszuaqrMD5GlcJgM01HNYJlQ7PfGTlIMklaiW2gIdo9vm4NHpnQtj9ut
NdruOL0CZXv22sPCwU43E/psUDFjK1rL1TP/h89Brd6VXBC+mcvMmSXFVV0O
e10Yt10N2ngTtil7b+78mHxPqC+12mP4/4yOxgLxlcFh+fjzHfPSL0dKrFsU
lUhZy4yqNwqqGiDU8TA9a6PaHw1LCNkxLWOgSsk8tIsWQXt9/p9q6ygY/1fL
FifCwA64IZ+lGflQi8f6APsybXkFEuRgvZqJIV4b//ol76utX86lnrjRZ8MZ
rDDrqYL4AyxsRjasxURmYBVV2ftu7hQhAXEyFEcBRKS4q2RDnj9ZxSlYTa0U
KTymhM5dJTO33mOWdSTzbFLbafvI9vqWayKXdIbQNJ+3wIfwQELuo94JN+2Z
XEFKJkIk776ku91WTM0kfWRp++x5eGo20eewzJ97OegjatU2arAOx6ge34t/
AvZSYgbdrduXuOeXM84AqDmRjYhflcqK5GrkAZyk0kXmWvDGgjSe9Zl0d6oY
66DiosEdRvENvmz8tIBh2Cg213X6N+CKAs8XtoqH1YxgquDsVP+ThTW9xVZp
rjmp28mYa+TmqnCFp2jTrtXJZXaMPwHoWbglllPlIRCiUbheVTvRNo27jS//
C5mX2K45PK+3QPeIFvmF0r753s044JKblH3lIhz3VA5epyzkrseZpcaiuFFc
1b29W+Hs3L12AQdWTREWoeHB6vYwtkTJTKl0FNgS8nflC9SzKiGOeun9GC5i
vgROvB3VGHvfPKi2q4UUe6/WYr+sHltAjkeKG0aSqN2gdpmK35BIixDIm49y
/OIlGV28eqMB8C8dpBCC2cL4KEcZbB6NZRgjDvno+SZ3UAwPTPHXj68Yk9h2
jsmUTLrKSiibss7SY4nsuI3z+NiQ/zjFFm6LzC9eyjNS44ckDoct9WONTobT
RywSYMRSH2MyRJBL3ySHRdtWwK7p4L90gAq6oGkzTwELYCwfS2+er2WP15Gl
IaqhsNOVp+6SMz9PqUA/V9U9NDdKEZG/59bphpIMWjsEIUVn4DP5ut0sJB2p
RInNE2XoLrJ4Z6SwjUpYPxbSzCFwDbTf3nvBjP715SZUssXTp2sUOrwdqOFz
6PguVDZDSSjXFNRmJKyJzWh5nS7Zk+S0tH9Ek7URyFICqFZpGsA1kZJEVhts
0w4FdZ4dxIdJcRtLijjSI2GUzhTznG6NHBLTUQ0YPhjAI7IQG/2h8tv6EfCi
NJyTzs4mwqXfP+PMAqo3FSU0LJ0FVVq6I79uNHmMG6kcCKvRIhyXVD7BM2ip
oz1QKuhTvzr8TZRIRBUuYK5aG2ib3SaPC6Z+cSJPJw3bs4XmVJeOFxyFGBvg
YdlHMBtL4uU/85uPsJJv1Ab89F3AvLslzCRUHwM0N3SHIRGiyyKAZWDwHGiC
9nMrnieuQzOeUyY7KmvkewbGw01eq9aKQqvdJGkveHH3pROILqCH9J22+33j
3jEhlmq97VP+QZk9DSi5WodRASmj4Z2GukgGkJddNTZG8ZYYzd7nMtoznKzL
4N9kwDbWZ+FK4wTozeuuQ6+lILVNjq2sHQQgGN0H0ho15zQIRnsM2uKP7g8a
eYLuWrZuYCmKl7OYmG8A8S98Q71soQXK5O07C0YfaWIDnUJLl1KRNhIeK/pU
rKcM9ls+9oMu3j4SyX/9pprtm1UC2E5Z8BUvdLYJQKUNHTOXgWn29QDVa6k9
BZBPwGNrlcJoGS5XeeS15dInYSKvyeQf4/ylzD5B14o4bSvFm+53nl07qhLk
dbtFvFpleXzotf1YZQ37fnEq7T3GTnE5sUDQIbO61fE/MujLzSIVCvA7ZsEs
PuxkidGcbyBSVSMg1K5Vb7vSr5bWy6dumxVXEGBaXouoge91lIR9SMBtW9KP
gqzlOT/2sx/PIXVMrkUZhFZKtoovPHVhF5jyeyuTO32DD+jV3REAQFR3I93q
2jVNCiXmrTn7Xw5MBSS2hYtk6ZgPthm57NB6I9Oj4S09OXQhwGMtFpGGsR4U
gwkEc763a0NdkBtmlEJFMXwnkZLEbflAvrfwAFD9E2nD5FUGftiTSF6hqMgu
WT8RgHEGEQ8FH2CjeR4n1roVxTnCV3a8NhKgVq3/FZdm4JQV29f5em5e9Hkm
r+dA5OowOkfYfL9kEM+f47zzIO3AZnHTYoKZc12nrqQb0QYKetF+KlrGOIn/
Lh/5ZASMoiknIiVeI96AZ3ftFA5ZE2MDULJjMYoYhUrFLvbVkTvuqtAavVdp
Jqr3DE/f/4O+jp6mFR2JJaDB2sDPlGsJEj8vOst4xYdq6MVoBevxub4Sx/M3
6sHMCH//asSdO4oqW6hR8FpGI5ncpR64h/2wjgajsbz9xkOAPml9uaGRECSZ
ohbFrsJF0hjolLE220/PIxp9VWl6AqcT6y4FsxR+Izs5fqHNXcLl1ODA5wCU
vorNsf2acj32xZJjOpan42uKmL78rb5oqErMOyvJtOMPzEAO02CBJKggYSAP
ULe80nhNJemdUsLnjUa70dHBBZWwkcg63GkS8xV0q42ad2sYWiTAVpRatoAy
LCb3DtyV7eFCxgyOrRwdld7T8EdusZ2BXGgIvaFRvR5BKdJlI1+LcfmTqaG+
Fd9Z1ZRLcZiEWWWByzFP0JGGy5J8Ee2yFTWOZd3/V2bWMq0jr/z+KLcn+v0H
BeiqJk8VpkzG9wndngKePWH8SN0OZxY09MJVxrJnlNVNwx+k7KRgQGbyK3dy
uPY36GRzD5MhS23OgE+MhgM+BXNpm4KZe569ql8O5nfovwi2+kPS40pTuIO7
xAORlDH2GjJPYpINP4rtM4I9SY0z14+bBdyCRvot81+9n1EV5W118Mm6YBM+
iq87CZ4yAbx3GxMt3N6WUFTXQPWAZWdGCgrJy/yBKj1khqaovyJ6lxgcwsXe
o9+b+uFDJzQlNp+8tN/ZIiA+b6wFEMVxWwFYLJsSHUAzdOAmoeJyq1I9v43N
pwGq2x5D5e6TtXYMKTJuKPovkXGt4Y5FaTPDk8pQdbdFkPR1j7Re/u1nwYZn
TMCngCgnK/xQSwTMgEeb+EDOfboiPLQHYYO1ggcazM5qXpuRYQxa8C7xbU7/
FV14cQuWyIL/G30uHUublFEkDbKv1UDiBz9SJsnHLKKERVmmaBan7yPTiQyq
v0B2FUmJt6AqwxgdrK6dY9gZj4noWKrI5/wxa+LzuvlyurEa52yAXKtaXO98
1TkwOxKL6nVST7dm3TwfnWehR0fOcUHgSJleRHnbMMySe17sd46MLuC6SRH5
C90gR14IOZ/HJ4nOGoQvx6jUnP+LbLf+MdfpO7gla9Er6CKQ+XBt9re5erxu
vy/C/4YdcU3F8unIA5qNMnm7mJ2yci11lM1Sqo8uGhC/iLTnPhk5V9lN8Pd/
0++lblhmbAmQ5Mdg3bcbX3n5GH3esl0JbXajKwKXsKlq2zveTgslTS6/7ecw
VS8gsf8XqizA5u97xA6I8yBhAovRi9lX537JisdspCw2WLwfJY4QXT2MRuQp
1xcFnOk0+rrgq7FM8RPQI2iPyJAkQH75ilEyLWgegS8npYjkqW9+jHyGt4eu
NOOcYsqIOZVjiBbeDYmvgsfpgopzdke4xpKotT8d6+vxFegtdvpKnFtS3jhF
q6Ju0srQp3G57rp1zC/MstFNwpNGA3dS4jWRKEY4A6zvZVIiGG98DGuAG28/
83CaITm4QI6PC4+ZiEO7UxQVAEOSFk07esrXRCTXFNqnCPLYoECR+rF7jTpj
+rdfUtEW1yUp1tm4gp7DrH078ROcEkkKY/U4KiSnONUzLQyYZpVaqaW3z0qe
uDN5aZYcZTaCRhjjC0rpIbrh8eS54tum+n75FJTCBEJVXBgaboWZZd/4hqsn
LStBpKnoI8Hu5kKj7KxWwZtTT2I4REcHlimieby3A9sbv9T6zEgVO/+ciGs7
Jw+Rg67CZWK2J1830TnhxRn/KPKKFdVYIFC7R+Vn8aa/ygrlHUbQN80tXk68
8/46TNfW7trxnXwKGuztHNeetx0rR3uQL5aqP6vOQEfNR5/oLc7aY5bQ9Vrs
6/0wxVAhec+4CUd3SUb5dmRekggoGJnIAAFSx6FQ+Hwyp8Sw2mgSNCJRxbte
7+iqaF6Y/UliItAt8deEZ7CWDpScQaGq8OluXYNpdWphK19f2Z7C0WMxIPrM
dYT07oVR+jTVgFhVktwDR9n2ud/ldjitgiog1afLo/ZhsuDC5+4gOMTUjpzu
mETve5oUZW5F7lEP7OS8jMMnbIwi0CRAgHVZwr0EijeqxgLmsmKWAFoEGcI0
4QYYW+qy4AY4RyBnsJ9bZ6cj3h8fVar4UGMh9+5qsbTDQW+cNZGFrOeFf8s/
acZ+x/qk8GamCujMww6hf3k33G/ZTVK41IPOjgN2wELFYRCUVgSnu8A6xTA/
ZOtgOAEpcZvPP87AkMVJ1+gKHEy2aqLCPWHGjDRK680NQfJZwNsD02p53Q4K
roRIoUWh1KntmcsYG3crgpIgdyo2gcJNJngiw1WYuUeWIQ5u6Muu+TX7t8Nu
u86+Spnw8F8XCeZpRRFMlNPl4cjrjOoLALtRI26jAoI0ujtOQO3Dhti7h6fR
Hui6YQlJHpvPbJUwWmFyKWmGVJ+zu57VVHfhVbXu46fmp6fS2MnQtV7BbQSF
ZHJALE0K6lBWw5FeU4LgUeHbkG/hzgrJPKjYllOnndoe0bEQkg1Gj6pSLe6j
ILPQYas7XBH9gljtT92ZjaB5BGD1ZLAURyjEU6wlrD/auuYbnzGmOU9aBFdA
EhmoNcSBFU8Iw1ggq+ku6n1XJ80a1rsJ5Cwd7V2ByMqSbWB9U+DSJG+o4s9p
TRjtcmSdLy/qjBXnSDSjnL25kgRmqmdyV2BuHJSlfd8xK6c4IygIW+kACba/
elI/PtDsXRGYtT+PwjUnI7iwmhs6hWHbFkjJm6adnynYNMdnkxidRpqyzvLt
exGxBn1xK9b3qhlSlACiPKrAQomZ5uj0p5cpomGQKXDm23TQDeqz6+vmbnNb
bk7vLx5f/iob+9D2lkQ2WH/31HLNPCC0kaYENDcVb2qRxat73urH2R9v86ZC
xhs+zGprm+UPt+n+wI/NvXgNltAxBDD0cMezoTiX6xlWiG+iiM6/dOEtTCjs
PgXfXWUrSC4TnlOnKl/t9yLnJc0nHk4q31x/8w+oQYPVm6n1Ba7DPzRYOD0H
J8eptZ4cZWYsbgSiCzaFNdULXRhpzAnaSULGlHpSDs/7uz5RT2lxZvu6Iwco
XXZbkEXGtcBNSDb2n2w0S0W7LgFxUgb7k0MyrbbkB7VJnUfwLztobZR5/Num
6INtqecTX6P5ZhQosaYhtDlO7fstgvNlOBhRFQ0s24sYSMbzwrw+2tIcKsqr
o2ezlCqUiQgPdhfHqs6YlBHalWUGzVdM96uJLan35QO+6IEHbDA12A2qlV/6
+Zxl+mTngSGXb1PfndCIWJk0Il4S1eGffOh/SgazkcRzdjKEU7cWBatRgZ+Y
s8WT2TkzcQUYb1ljwRQxzAmUvgtpzg/kHAOjdkqVG/j38sWem/UeB//wg1vf
n96/idsbW8OaWAn1SAVMdyecEQsM43JNQHOQpG3OXG1JcrHjCw6K712ltrMJ
9FYaPwUxcfvYAjx3cxyx5a313co8UcaUOj3WeiLSn6sKu8q4I2BL+8M+62x1
PPeywMAhtwtwngKWSK2edouBl1m1cnStLQn+nhWa1JMqgI2O/aejwbpz39tw
v2FtWvU8lAxt4coAw2uqbCBvEJiaYXAQsZbJqRhsU3AtFPtFHpzNcSEmoeLP
LcWOxHYdo/EUOBbAsg+XZGnzXGf/pbAQKwnxCjSILPeWm4ULN0EI4RYHSzKH
d7h1AVGGwKvpSWxcXx10awEdj+Hj3qh/xnZlhNNedZvxphGkOaMy1ADcGGrB
qamH07bkUIowkvhPHqUYWPi8o0IaLcvSwbqtScQFJhkLxE1ovQQJh/y8dSTe
bkXwNIHDn7aAnTXHhLv63iWt1Cp866S0CnXXbtSJJUYJPELq4zvumJnAb6Wg
3zGRkn7R9GrWtc1FclJKNmfGzovh244icY4D5ge3LziwFu1pibfSoMk+nX/G
w0CE0XQwR4SlY7x1i+c1oiK5iDh0gWhzMBtXSMt5pQ28C45FMmILXJEabo21
X3LCYIS9SkC57xUBhmJgsPxJZR0IAYZrtp7HdycRUdHXLkQ5Tws41Pk3ziuP
9Mj8HOdNWi5e1wDfUkuLGwwadJoM/dKCSeI/QDOT+HuJICqDObNoU5LroJxp
wGXJ5cYgasjorTgVl/Apgn3Sf0dvjHBW/yCs6W1IKlCj615l3ssZ/RraAPNU
ZEwonKqctbJKg4JtGe7ZCJNLbLrSdSac1jztUBhVXssMgAbg1N82BVipW2Vb
8s8MX6YCHrISqtw54Jq4REdm8ObtRL3NzcEEPPdUn1m0kKY902l1S6HkOv2O
RUhAbevaiwk2gBvHuHzOGMacvXEthtS+sEXLwv19lqynSk8/Ll5jgEpnR/3o
3MabqQwCg9wXXsMqxLXR7ZVS7YBOJLkW0H7rKO3f2PpgoMub+in15jPmMwe2
9oqBAqf7huuW54oA7I/TQzEMemtrqKc7A3zDKefoOlNzBz/rn/5cE37i3zCm
lURWujF4AY8PY3lkTOMhELr2hJEDdTsH/O7q+srFvl46opDKvE2ojJ2da7bH
59HnvE0r0PsAoP1IV2adTReJiLMqiySuPw4fEEflf7d7PYuNlfzbx2cV1pet
ZRLByzbO7frS6JZe8cyumTgVbMpzSplA2AEv9RbTT1B/7d5ngN0g1/G5d5GK
ahZnHv5SZNSplU1MRMeQzE0JW8Hs8l1aXzPu2J+7KE1Yuy+JFeJovn2aQYHD
dovfaL/j56rIF9kkxAzAVlO2EPEx4rOqg+68haQguoJWJxJyupl0RdVcukgR
03hYa6AhGaH/c14JNgoIv4kjWMwnnGvh1hvzccMLZykCGs002idSYlPf5Mn+
Bv/1OMhXZZ8FWG5OUaDNrkEavMpCXHuAPF/j+nai7stpkXdYptq9kziNqQVb
y4UsHOUq/kYwsgMvhitQ/kJyw/odc3Q/TPxV4iRPoczJBxDb

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzeesWTUFe31H7O6Ut+AqPdRVA2XyFpxn/PFJHJJUtXG1urykEvZQR9tH6zBbaKMz06jPIieVZbiSmjSVDSvCTRbU/y203m4tXudzUpd1/YC10KXiY5RQWCZg4fF55wGUCfvNF8A72rYonZRNVOXYhG1gyWfSoUiYPo+dvrNww1gqO2B0NiU1u266wEUcQNgL+RGnUKaGHQEvzE0HSuRRvTSt04S6+PhNMN+pnzxxmHQYSHl+HIqbKwv7UE82fVAq/NS4gR2om5qtf3Fx8SowE678J3mT+ZJYUAkHmSJwy+dXp5VZ1EKexwKgIXAnugRIKbGz10EzQ+ldU3LqOxtd87G1+0dSjxnQibMHlRurTBSLPB6qQ4uq1pkS6kWfBY8YQi42SBmKlXaRSLj+eR3vPFpFrd2d1ksM30b6+skneDkk0j2VjBh6mkSlEb1rKDTOicRSPCYTf2FHRxYUWa9o90iaFqrqlSxX53y3DrNV1Oy5lsP8tIAWc3XvmqcNFytp5mSKTZJdMAz71/7chWOHWdwrBq7nZOSrLwAn9rAnBIdzGWcy2DG1mhHd4UKUx0/z/mXcdYiy6xMBbP5B7nF+FMmfi9jsS4PQehGkKDhuciCnm2Znymk3LKnfaBFdgwYeZ76tDsbT3yGh05iHdFKZ28MoaK8g6wAmSxAFXAqS1MWX8pgN9PEhHPIiPKqwfNiMkLNt/UAzovI1SyPdUMsEILjjmvJHAvMFHd1ExWnmTxh9gMvK84sqqJe+0t2ARdGTUbr78Kn9rtePJhVHdyMD/LF"
`endif