// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
loP39Qn85z7WpPgF9cLW+IvEt84BZQxfV8PnK/dGGOjzoSDkUCLVQi3zF1Uf
lu1K/KD0GCAqw8Y85Lq3S2+eb0YjRFIOKnIqShMGUfLVg/RJA/ZKN5QG5dY0
KSPSzakFBEqhdRq3fpN43bju1x0huuP73wN015gCQ9lVXP+RYiIZlvNQ425q
1FD+klgRhcB7sijJlIKzV7KLRfFuMkE4SmK54riEJvPo0302RBeOJcb8jbK7
Ki01YwMgcua/E3gGn7IT2VjEzD1S2BYAmviCvZkV5Ip0a6912BPjXp7fS39a
zR6prMokIcOyAttbyfn1v31VZ+R8Ow4pmg6gSwTjxg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bCseP9GNnP+yMB8M0usN/iNUmD9JmTrniVxLVdF7VkDzJgrVQEhrhiZfxJo/
d1tyaNDWEYlNzb0b1ddNZDTBURoHbeJ6Z2GFd9C5Id+1PNE/o/IJU/srXALx
bN0lGX16quRMExHDr6U/EjMkv0cbyHAEqUON/hRShQQw8maWLQJLDEEZ+ie8
fSYq1QXhwtHGHzNxHvKYCvI7Q0P12D7PpitCMUcZIMtjesR0uW6dxH8PTh9r
hVw1SsagrCavc9Zz/BT59V56jt3J1RG3jSJ4KJT0mNL3YWroDfX//qfBinIK
/LP4nqAJKK2kcrOckg6Zkez1w5DSL6LMdH0usVLeNw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gXrwZhjJJT2hz73+mM3wnIjTeU4Bb50gFp0PCZYlNoZ4l81rPkz8+YiC7Yv5
jQKRUiqVZ2kfAMmVGYyLQHsIhSDIMXpzeMdWXnexLc/a31diqCnsNAkryTSA
akhGzln2n0BNIuFbL41viFpI3EcJ2kVZ4dZqyfDrlfNMk7OeK1hl1C53jFIX
q6bru4iy84Z3jvu840IoyEKYt8/7jMS6t7JJfQU4HHf2eBXjR1WMlD/3HmfS
n3rvLNEVWI0clXX4OsFZoBp3A4nCeM1iibs+kHfVhADqr2/ZZ16BF0pCiVhl
kYpVeHWtUHT05YO+eCxygwyDqsR1zYoyyQLecT6BFg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HukVmaEA6wlWeAaPl3AcxdmuNzjNSchPOFvO/3GWv2wuFAC7lpufQtqKtB45
4B35/5valG+mOfbVTCAx+fXaoWWnKfKnb9nat9wDI4/FgX4scPqNb+az9b2s
/RLhR6KlCeCb2/S27DzANSofVDWIjASfYyHvFyWFlkMdq25jDGcLL+00sO1T
+NAQCJd0+ujPxNbwhU90+d17BdxOaxPHRvLU8UJVBMZscYyq1NQWlqOp2rjT
EaTeAkSmjPE5+3zqCL4cVcBl+wO0KEgUNvx/JINGYWiK7DC8HKqpLsubA+ow
YUxGVOjneEk2ur1/7FCHtvNrB8vk2vvXDB4L9V9uxg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SY5rZ0hvEum2ZyKe047zlH2vTak220migC1SFM3J8DyyuHHfmk8+4RnS0KQK
X9SlLVHfyaY5UASt+d5LqG+1pUaFw9f1/JlSFqhpxpqn+/zBhVaR7pBvk4RN
8VQWdjCrQLkPzX/KeNxxwssneK4lMvLMj2Xv2qjSWGldKbiCqjw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B8ykC5VxGxPsJXostssnuGt9rNy636QnrY0H+6hdqJrEO1dVwux7WAYlWuxW
51hlXKcJ87gLM62XWFHR+KY5tUvOATd+z1Xmb5YKZoFRefqgZvX6uvw2CD/g
m3yndJAZjT4RzyP4LJjP36QjqufETmMYqCcrx1DkOj+pH5gI9780W5b5u5ZI
sJqc1moMKVQp+DM3qdRMMQFPdKO4uQ82Hm/feGx9DMnqiS2zenHXLYYyESyb
BKNeHbNByjEzbihsoeZ+hRjAtmVMzcFYpAyxarfX6GGLlL7pepRA4HuV2lW5
EqtpjfPhH/3uNnZO0IawNqO8z9ZrVSs5tiUmbCnTE/be8U9syyP7kg1XY3Rs
HVu1PsOdl0NuMHeHh3IEt063r+fVW4McWlq0XmCR7AeiRZx7sNMjCbrUQvM9
f1zYAYbjZ1wEY+tHGw0BSzxlnmJZ/aVc3coRqJ5/JBH26/UwTGdsZO8sBnRW
N8ug2YxtN++e/ddrMqpy3KRjk3fRRI5t


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
k7nd+fsBbk59c5YJwrVbRWoGa5WEXTzRXX4TYdCnzFjQEedpi6CbXz3sVCmi
by2FnJPl/ig98eCX4WvVjI9WmzXGpegYQwqBmbabfRNnDGonJee+bZ2JHwSd
vu1DhwV7ue9+uoy0YvcGlCbe3qePMy7GMCXGQHlX0w0mNAim/h8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ja4DxzCtav/ieg0zSO1ONEWpf1N9hXHDb4GmqMB3qjWL0Pxk96nSZ9y3YblR
ddi8nyUhRNc8QEvQ7pxcTTR3O0mOB6VTYpL1TnGdj93rW7zTp9ipsEpNVknD
LIGATNwyd8/y2xbTAwZMq5QR2oqxUZ7o1oNYA1gKtNsHIUVziBE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7440)
`pragma protect data_block
4sYNi2iugPeuPw5aW2uq/MOimlGc4YDBhsalkRcwM5kGucN9TX7SPkel3hzR
CRtNWh/yruvDXz+MvKJiURm/zTBf8ikW3whuwDdGJNcD8BPWeUwHdYjUoQHC
v6aEPeQA5a69ZjJ/8/Wb1CFLUjroxoVqdLC9YoQjY52IIfQr13DlQ1xWNT5I
kIiv5WVWuVmBCAKkT1oqUw7kt661xL/8J0tAz4XHOgG8RT5quIAjSLb+gJjB
/MedAqj7cC9WTeCOk2wQPjMArBSxw5p87Q0NdnUPYuD43MUJAuOPfwk2WZm3
qEeN23NKy0v2Jka3a+Sa+XO9lUqwv6axomy7ETgjFe0GcxjdpiDY+44+KIny
4D7X1UGEgcQSgJBMlUBGQWSNZsVLASu6YfIa6GcTGxp97Wv0iz/3RP8zqs6w
oNls0/fc0lnq4TPeRziSJ2bHYJHlDhSdZDsUtrtJfZ2O2jx2ejme78e/R/FY
yqhvtPH8b67qfXk/17fkbKkcBFc6XNq90bUwCX6Pb2StrNPPEVKLKB4/mTbU
kpNUUcO+2iOc/MiSY0UBau5nLTATRLInnGaa8PmcHnX75XlgSX7n7e2ISKTd
7cNKOsfFh9hVpXgoEe8J+WCEUqrieIhybLO9wH69Dn7dxKdpXe0EvQkL6ymH
p+GGOwiPwvZiturr8625KcdIqjiOUEQe3ay45uJPEz7ngs1CTI9QkbfjoLPx
7LHY1nxFVKQ3IWa6Av9sGOpctaHVzdvhkBhdTHBYZPa2cqfvRZDFUR9H4ELY
0EyPykE2EgWSjiPrzUGhabiUKKOGrMG1V/Xlf/1VsVDPTCR0Wk1Yz1PSjDRj
Mts+FeVO82UveKlXweitlwalW1B2WnWPxB1LAm66IDdvARQsIAyZBgvnM+lX
HNvsixvQCpxpGY5yjS9jj8kE5rX6LnNviPfW9gFSE5jpEAQSl9h5agffHgRt
i4m+EADwe77zcWAF8x+mZry9r6Zgi8AFoM7kPdYMS/sHxSdrh6YPSrfL8iu7
1BvSVvbAO44bK4PvSaAY7pGOdPL0kVIr5GPCgvcblNMi8NA5g9CdS28w6q73
cz4Zn1Z+p59YxdLwFWTl8p4csqIrUoe8Ou6PnG4v/y0FQJx+Fb33QjAcr4RQ
jlamSJowH/POSZpN+y6Vx8hrVXp9U8dXGGePmfXid2u0V3wQWwuhbDrqggPS
oqPUiVaZF7Sfd13SrB5rgx8hhr7O+VGARX7pJ3tHhY8K6pZ9AzNn7n7RUnby
4OOufCGJ7fOGH9WJAhlLli8fPh2Q3eJISDN+RZpi/VxaWeF6tSUQdRvZL4LJ
+77f/ncAZI10g2DxSHwY9l2TG795ETIME3GUYgikIqRd4rV1AHoKOFZAHcgt
3SqOQUqVwB1wVmEYnJxfcoJExbLc1S1L9rvN0IEYUaCQpYlQ9AzGeXPOGTxJ
XD/yW2uqif+kzhkROxOXiqo4TbySrQbaxNl/0+KKtqO1EtHe8ruOzbWknXN8
hIR+HtRd1hCU2oycB1JLljE39P1+wr/Ln6+7SvrHm58UKXTQQCvztTnA+z9x
uy3sCyS2wdr7Km7qzvNCZ0ox8s03ED+iGxO0HfZgFLAiWCh6S5dxqzlRj7yC
BzQ2KEhg2PJp2ZMbIMEfMRE/gO+pV99G97fjrpqEbYZVf984kPtnLatZAZdt
gPl1YKGuiG5oY8KXRniumGg8MjZtcIRCPD2Dp4B3rKWtrSZxCggiUrKkm29c
KOmgJFZwvuFli0+GruxIlmMbAq6aLxXoYufBP9GdfGpMNnqopyPX6vctgRmm
O5pCXXSKft9F8xUgdwaHsYTzL4vIH7kmh5H3PBi0eVujHD5MIwRybVXuzbOE
AYgYt3v6sf/+sD0pIW9O+z88MOZeli+/Bb/0HdejwZNa6Kxn/yaZgd1ADyW1
05Nh/RE/K1FGoOnchCuc+5hAIi/c+e4E2tIlDBN7U9t0xWldBUymBFx61uQA
bxVrQwdzk6xvyW2qJXZDRaLFNYgPPf8ampGuImXyt7OLJB4toEAfuYa4yRY1
3aDI2xqsLvYk4jB6SG0sqGkXON15qTnBvXR2O//Ytegi0cPVLRD1RjPyHy3I
ADiAKMhJEGFUTsxDaSUDElFqKkBI9zm5gVgIEPwCEZWjpJrZ/d0SLNLsYu3E
wsldoizxdf5CGi3+NM9p48y6KepnixRhm+utAnmyhy+FFAm7VDv9MB1rui7A
WuWvhGIJ9UH5690V9L/VACvWEV417GwRuB0/WJOEByUu14B3SmdKbZPyjpYc
uYMrSfQx6KF5eaUuuDt81Vp0N2PJkdJlQ2nP3KSDnkQ/cxmIrrt7AZdDfHXK
Eug2tToWIPDqLHBEV3CbQW5ktaNZIcjRH8bxUaOrwbpoADQsMnYJXTE1F66F
XZ/f7dCRSFy1E0/vZblwuserh67TXRJou6ZJhqdSQ0XdqPDbvtp5WsJl9zPD
xgcXp4YdfnSDd+/Sch2TICTpRBzqnUPxUGQn5gdvOcjDrQ2XD7NbJbadC9hD
mCuZ8MWDv1AjZgdUwpTl0r8zqsltce97Dk3n3relqVxKTuHd+gxjbtccFycI
qn0t2EqLNuCKRJBRAjUr4RTQR++jHDZPxdyYYH3xvad1t2lWyBxP34h5oVp6
jzO3ohpnCnrUld2PyM3s7k+lPTtqpkVbKvzCLH6tSiycjJLicf0fPsF9qedq
hT5rvFPaJ5YvpG/ETlrimGLkcb04PXHKmrVt1Beg0aMy1HBlg5B/AZjUn2b0
PEDIyFE5Q5jnT2OWDSdGiylQMTE5wC9iqQ49KIjV0dF4QozmnAJDpSO7h0eN
HOAjspOMJcInoPN9vixjX6Dxgx16g9Vtmf9UIu8MwbnlJV+MXoCLGLyV20tS
4DSHaNtgtfhI3cIHHU1p2+whbadw5Q6zaHpPgzTsvE8vNVLKX+E5QIaq+gfy
vkaE3CeY1HndhG+ZF4lWeKut/DFIu1nLZNbQ5ZKa4OgD0VqM1/52nvC76UNQ
6l+l6DtdYo4HFeTS7O3tN9U2GJ58pX54TbHGgQgCTEbA/dgllWzUU8JmAs+6
qBdsNsOwKdmSBZ63mPc5wR2rMOSFHft/cp8SQODfPU7oJy57t0LsRJt3M+ru
0sVJJfil30Ac0gPThCkF25DJLaKqDOE6XNBoGEmU4QycbAY0Yv0akxx5WMoO
dndwTokOtf6kK9VHbrIKf74wSPp0NDqh3CxH91+GO2nnmLv8oMBMP0zGC7em
WdHzIhEP6ORcy+XQjl1pQWXYmSpZErGdsM+ul8vjJQ1hxnHnAkIojOvmW8/s
DLZ0Vl7JLzG3h3sBlhz4IsZJLKgLYQ3YlbXB53OD2Iyy3KHfl3Hu+r2UzTue
HKrc2i6hkoZ12wkyRVgm9dKbU+ARM8HqwuZLkhH6husua0NQ35uS/k+sDugx
x1m0ZnIulNz9r+kxCEJtOF3vWmdjHovOye7fhL8H2eKeDfkI6A5P9Afv8en4
tNdqkYI6xoQXOJMhyezT5lT1SFwgprRPGZkWf97+1wXXGdaA0tAqkWH7h1nH
5jD1icUTufZj0YjaA9ctvYivm7CTPxM4ND5CFXjAApR7hfSIYjsPYKQYe5x+
RoSic9l63FXAtveBbqXw9cUDRW24XQKWDgLszsrMWAfqR8z0F0sKyAza/dHD
D4aEx4ZK7aY44M8GN7LnhnSdo3PDD4ftxTlk6yqRK5CbBtDJoP0iYQ2K3UEO
+yiXT4C9DmjGtE5S3iUofR7EyoY+TYwdfGGYbkvsZZcksMNUm1aoN7aL3VjR
3w0CFeiVSX9F3uU7ONcZlIDaMqcdv9/Cq0mtFxdo5OK55kzdVeUpr2S2tq5r
uUYAyLde+nZdAcZ+oPfU+71G+SpCGZBW3sJSWtT+FhfjGgyzMoy6mUna7Rcd
pbR/D+gzh6IJVMbMvfhsDxu7wobSJun06mwYuQHYBP0OHS/57b8o5t/wlsSq
POrc5LDUtZyM7goPGeSpwzfNiHwqjHnSp/hZV+6KZT/m0rccEdCXTeHA2dBq
PfnFWgOqMgdACYGKJRue0PGTZOqV52/RXZE+lLje4C/xnWbmPOxygfmoqjrr
LOUDHYc22s/MCFXvyqn+IrjzErFNq3Jn9ZUfbYo3PqFZl4FuNlDFcUZeKjGc
X/ugArkXDUFL/QBH4lWZyEYxMk7ho1gcbxmKCC5juCwyqnEet6Wm1OJ9vEon
bUnDzXa/aZ75T/rOksFj3Tm8dfOnBDNhXCdXGtGieqXdK92+msAYSp6TBx7B
TzUPD/hGKBe6XScokwPyrUY1pqHBvNfIQQEPIylVdv55azPmPWvI3FDnHTUw
Bo9PuknXHs7vh+F2i8KvrO5gjmKFTp/f1RFC1RK8h9ROwaNPIh3N2qECHapb
6QxffqcLEJO/RDR+l2G2gpPTIE9BNWsVWpvxbsbeRIdogQsv/ryvDSZNd1gS
ykbVZWQ5xqzNXOL6a4IFo6Ye0zaGlL6U0i4OUWmtXHEfMWwoyKBcSwONP6sC
aSvP0DMfuPASRB+iNc9LrlIoonv16Ug1DiZZHaOTgLEhHEpLT9TpeKfOuCOY
y+kUesyUK2hFKbUIPngIRhHP/q2MOqgYzlATFjuB2yHHPgXW6QszmN2JN+9F
x25rvqdGW+oSZ5Zh7JKXvV4agQdzCUhpCLzu5kyor9OX3N62vIR+be/ZjWgj
YuZaWPEaoTwDOXX96lpd5mk40nUIIHdSBoGfE0l/WAdnRQl3yppcs1cKkGRj
8JDrmOW0AJt/Lw8M9uTBLlhcOweijAHoFQ03+qSem8xDblZpzjiFrMY1zbV8
8gXhDlPoRH3bv8iiguGoAyZ+K0junkM9NpR7r2hyd/Z8srpk0DFPIevU/y+2
XblS+KfEoQbpL0krEhPAlO/0tV/HW2xGK0XRjfnZvbsT1DgJlIHI85gSaX6b
4gBDR+H5NlARQC7tWPLPtUOUWk1VQEY+jf2381d+CqFEROh8XJExBalqNU4u
Y2/qPL/RIcyzTajCSVKnEdEXrNW0Czih/L+9BY6C9SorKhXJYDRtgWuFlQrd
pRIZ+CYHt1tLUiisJpNkWj7L/W9XuQmbIjt6ntGq1+Y/vY6J/UfTLfjEJKRs
2iRp6IMsNiB+d/BZfU4DDLOcbWgkGyT6qRm70fEAYZb/7oEziWPsCgFNix5T
8ZBwKq/cGRkIj3OQrkRA9GcadzgGc+ntg5DNYfsrKZNantwIaqHJv2Zkto54
y3Qc4HWOiJKXg9M74SHiNFz6ocqLgaCGDjPERws6d5F+DlXT5ou0lV1PQkYd
uH4jLlT3MkebuF/oJ0WKmbRZcUAdm6xVGO6nIblFk0VERwA9WQym3VmSScoT
tSsfTJymm6Zaf5qAswkGUJdwuXAzCmRP5OhieUO7+codwYDzjZWCximU1Hv2
ucHc3D6rum0lO7Ek8MZnoEfn/W+ZFWCu3n69WNfVsvC9ndWPwnJsrKfcMMJY
WQ2mw/Oo2FImVHfwlVLtGvwnUTPujMK2rxwf9Jd5F5NwrxOnIZQkzoFTdFoj
KGwabQsjTTV/jDjxkH34NLj6HrXk15ELcJD1k09GPw22KZ4n60Z9W4oSNYMF
0WUKHh0j7k2aMWMZHU+5/xwoQ74Kohl3CJUTUQcm93mPZCYMxjhvQiAVIrse
dChlh58Qx963LIeQMrNVecyMGTsRiWE/w70Mpt+mtz+sSHzjWTxN+M6y63UK
WlFW17lTyXQQrFkmTJcykBo3b3D+kzeHmod6AfbWVZU8E2ks5p0wcTTCXy+n
Cn5qNTAg6QRRbzFbasuvkipMpol12T3bRm0Dvz9gTXl6LflH5+NzBtU/3CK8
ndtqsKjBvdEeiFjo4hjri5syXpRYucdj1S6BRbqxIyjH1SRRsnYni71cBhfT
rHQf67xBMIVgyys6sKBWMaqs/W5Vw/dL7eNt2QksuM+hhMmHZ2acgzunFPPD
OmAqIbFuqUdbsx1/jgRAXPDZodiBNmttfYrqaK+fQ7+8Ko5GsADH1tq6PWj1
C4YG5rEXpzrHhsz8IVrQmcDvujpI2ltbdce34M7ZqgBt+pRALpybjOcoJYDN
Ty25amvNnJ2g/Mi369U9Mi/TTB28Bx/8XmoNG+jiT04hAG0nArS7JvKlh/5e
FRcIfgPiRyF+wUb+iR/b3SUnyvYDCGBIubMXBiK42QJelh4QKRvzZN9oYqDZ
IlXYWfJNPnUaQw6XsikvNxNhwBZeT9YcsRuNLNgBV481eUBTECSJQHvIz34b
d7W1HpMNRtCmforE3jcpaPS67q+QQdwjclBqLP8W5ybfHhpeYJ3wK9fbsdfN
V7csK1K97D0UnJiCKIKjeObfGdZglSyeQKToKFiNFLfAH3WpJDytRwJ0mzd8
JcOIBhuwdibKj9z52CXh4BUnFAJBus4ASAmfb5ID3MJLlZV80reBa2Z04ObI
ATJjdkF2GH5UaKfpqA8/MdEcz8SD5JoNDb6woiYox5AMGB1ybMEjKOtIsAiJ
F4dTyfrPSDoVPEtnS09cWJjRz2sWLIFs+o9N0U10zvkZeeZaI+4X7/joeCTA
vm2GEpPPm7rhQ7Rr746rnEir2pWbUQrlQuimqSByGiEKZvx6/oUmSqZiVHWV
3+ACWWY6EN1hDUQ1QUPP3uWueNWXOXTb5T2GH3rDhiGMHMK6GVAPxsuujr9J
EU3y8bSIxEWubnBgtSRRQi37IvdoArUlrVebjmUjdACrei/nTf87txlB9UUt
BvntWvnV9Nwx8mhBAbvu57vDiRNA7+ILetCKZCJb7nOjbL7fUh7AelUIUloe
cUtUx5IPTiHD6qAUVv0giApqNtGWFOog/8Ce9oxzpR0kyADdS7SVc/Zs8YQj
nwSoTwDkJAgSOJZF0ulwLHCe1c4LNoKEUqKuaGTsxfnZLH8fva/jGek0tcnA
6e1tKUiYij05lOvVGoYxmYpk50nY76tGH/Bm7tpFyZc3jlk2dVvEr3GndSwc
8843HzJAL/S+uFngTthMSC1dW04dkrF7TL4HYZ4FZlaTcRHhDx1zgAKEd5Fi
non/wI8hn56dR4Hl3CfmdL8I+ITWuqze54ld03tovRCpkaUNDjiYdiJtL0M4
k7MwC7TO9O1cyNjAfXyKX67X3bJzVSNA3pVttRU3dinvaiUA2VcWi30cAXRc
09R96AcfnUA3twOuiY3bO92iZK1AFH7MnAQe3hKkdz+juE+ti0iiFYgMT5kn
pE4YalvAkJAsdqRxyvWFweFa4jndVgH0zpuC5nwYHvmMxCV0Xl/B/0PllaP3
R5EjAKrG+R9AmE2eA53LHcmo7fDXoSp8ylefEgjGiEp658TzFBT87MKAleJ+
VAp77da+FxDZyC72k4MsnbTZJA6VRGTIgixPnSp6jsBO70qph5dKEOh23V/X
SXqjBYAUqbV9KxtNIks6/0P7XhH45gBD7zdFSegkqQsLlqjiaECHIwleByg+
0wIvkCHAnmjTbAceqLV8IzJXTZpNHhfoHiBqYLRzX86kCRMXIRehGh2qZ+7M
IcujJP7NLnHpS2xTntCni6oqWqn9Kc72hp1Xnf23jIIBBLBEk1DblR7u8f3a
w0eqe7658sUh+RjbKu38kZqpDQgRPw8aYdGv0jIghAvhK7PspnSEwdQSAWAJ
5bntYE3KOWQ18E2mk86tg5UhcAGuYv0cqEBdJNlR6n1+c637BcAaMmf0z21e
qOv9PXUwSICKXSYNXRdZUTbcUMdbh3WaXKP9i2P+ImPm91zIp33+hjYfv5pn
DF8nf+RT9EbacyBUCcSUzNyzTRdD+fDngGjt6ak2UnHduxUc2VKFgWVwcKcL
AjRz9rfYvxHNNe5//kScahKsNoYodniH8KI/3xzPS1VWgNXErYXi9J0rPasN
fQxR/cfSZoMwwghCMmpOi3O3K+vOX13dkxrxiex7hzrmAqEQJZnQ4o7DdkB9
nE6Dn6w/xEqecbnbKOV9ZArmsJdiXV1sb8yYiY54gAPujoQgk5uPDObrxdnL
rYKI5cbDH4/Ri4Osz7E2CAV9+v3I+F/GCqFQQzYMUCjPc0I4EprEm5WNf9o7
JMig8XPWOVpw2JTWLDk5p/DVJ9iPcKeNF1j7esj4qArvG15j6nYohoYUWOWu
Kx+CHRVoFztf8sWli3/XMOX4E5XVljJy6NZdUh7whUqXcH0+iE5Fjnh3m1HB
DWrWYMHnONeb2ojxxn63YldZ0z6mut+53LgJNh1xQHbJM68MaZlujjheD0R3
XjB7nkdOSuHyBrTB1XZYVx9Kh1jGeniV/s+MguhgpWtYlVO9f8spLuD1spic
l/le48nPgmeByR/ynsvkgx/3drwGTplMe+xutKyg4FQc3UlUXSGIcZP5AFL4
Mje36ZwvwtU5fCb/BqTW1+LHX5XkGupoLmyXLySDOJ1UO9dP01Ay8G7BvZIQ
1EzNj4J0z3C2f/csNEO4vj+vesb84csoMXPwViGoTdoocqeRB8Ka0NTIu43n
dL5ARg/nGsPN9qp3yDTpRdRyckDW+PYYgvnsDEYvwk8cXlzmR/umR1cYGXHH
nRuQG1e9g2h4g06VSJ+D+ahX8TvLI0ueCPxQJE/Xzx0t1FwoclDlQFJ8s9hk
wyjIcM/5N4FVHQAtuJ3iqk9WhRejOusaqnfhlMMhdAjvZD0uv2KkWlMTxHU6
JhzwO9sF1+dGGI39bpKm7CObKbgnr3Sm+ytG3QlU3z410ah8bzaxpu0JAzT0
pipRtcYhI/jAZsYIENr9wi3HToHUXpce9qwYLEtqveVMYbTBaOfQE53Yjxkb
d+Zd9j2JKVNNBcDco8HcOQtsFTC47ZdWEYm7tuJ30v3/IRBwJuQWQEGrCw6x
SRjslAqph8BRyRo5QjkF7VHb5ERCq1obPGH/HCT9W7lR6RRyCDsiBDw8UF9N
LMy1//sxaYAW7S2zDH7kQj3ShX3MltAr2qRu7WatnI3UYHsLCnEzEWwP9zXZ
D+PwLPMFnQ/JR1Y9mF4zTOpr2l0JpMQsNa+qydlQXczIb99ATougBJr01X5q
qRmg1zTYPH7oayOEDoMExkCox+Jv6OnbuBKo2DeHfpQSqpgQ9imguN9UwYUr
McP8AOEbCHVzfBG6rFlKiWQXhFr9LvLZ/vJ2dmYwOqiJ5L22OhA98whj+aTw
H8EcpWOPSg8q0cXn9Hhd2ewfhSlDSGUkQXQfHGS6dKm5nemEtU9UB0aFFiZf
xFHVhnRUI3ZS4H7D4wVyhQxXEa4nGbe6t0H/tnHgsRflbs682SzEyce4Yeou
havcLewl2dH3RXOFieka0leREnR95rbMutHC+BqZKxG9gzXhnlDpd/ivxL/Y
9H0I8MNlfIpW1YJopuaNWtjiGoc1BTxSLODZGBN8SG00cNiGvuytB2ggUiDG
QcSdMm+lQDKbGIGL/feE/2LBoTGMDGpsC+tINVBx7ujC3cBEzPrMaHSPoUAv
BWR5+OaALFbSUKfDuy71d3hT+EVYTeptez8N6vNWFe6PsVAyIK2qORJ6Q90K
S7qWCSvUQ1ZP6IJguO9IVlqf4nJ1mAfGpC8C4egPBZLphqcNwyhP5Y/But36
MHOZUayX1niQ5hfbh+YiMph4PbxjEcYENsl3hL/UbAeEWjjqhmDYCHhONRfo
3Dtbpp3XL0YYacVUgYK0XPBI0y2Hzt+jNPCI0f+DnA94TRefkzCx2qaLcvUc
vHO/PJ0muG0gVALTkGLUSm1O5pMFDwFPTAUyCT6+I+gv66JfqNu2lIBVQsZh
8ZIsy0TtzKsxQ/oeMlRNOQh/vYij8mfPzgCHUdIIbFmir28PH6V7SS3TM44+
GqRq2VNtixOT5aIMQ1gQ7rlcN0nUup9FQhTfZZRn/PyNxXZZDbzrbvvEZHtx
Xamkw3iUHE0T9FdkA/P4+pZ5b6+04i3nwG88jYzi7glSRHWG4+yG90EkdgM4
ZYGN5PdE3ZvhcogS7oWY

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "uNqNhMjjY6+eXlQ+OJq9yNnSIVY1D0OD5CiHuujhYhAJ62wFeOdKAsHRQJWRoCj81qiY4Mxu6yEVbCzi7Pkvgv0W9/ryomy6FFy80PVh++TR5YVo5zUdTBm3qpK1m0rz8mdzZk7sNdYsiG8eiuk8Aote2A/AXeCMC7FZSbma2MS5D5SHrya/QPc50zZtGF/n9J0iLP0rILV00ShPkZwO/1deotx3YPp72fa66Z+XTa+zh0akwsns//5GCa4woaY/3oh2CBRoV2qrXUn9AIjL8Tc5CJ3WJj185YiXxWE+vG2yYcn91WvwMppCJrpDppTdnR+TAjEpvqywZgm/2cQurCvl3+68UCBTforrsDUyySEptBRp08iojag8P33pEl5ZOOeyqUumJcsUc4DvmOUVYvBxPIiQBGl1b5gCf6Z1vtuzPnEFmPE67PzzsNZRNvMi9E+vhocZFaeWRZNk5eEDpKoeEAB40I+H5bUmbMKq11hcuwffMVYXR6Bd6+iPsTELKGJubUJf4OXkag5yrFVEbhZWnaUDnPKf05HuPcPKoMUoDgtGVGBuHnm7qJLP9N+BvXCmCZHYiZFEAARlDC48uD0jhGlWh7+Vv65JTK36J/SjJtoA+GciiE07Tm3Nt9YuN1c0sf3BQATSuksTvm7ZP4+qtscWo+QIf/jJ9lBQpIIgT1Zyf1Z2YSh++wd0Kh+V5T6std2vQS9rPoyM7eKQtdyRe0yRyKRfK7qYVxjz6SFmLNd5bT3qWdKw1KRKrlPfiWnABt09yhcGFhqu0wR8ff262/wdSDV/qw8XyrL1VxHOPPOQFkzyx7A6f0aW1tkd/9wqMDrwcuZhD3kOTu0J+bZ+FhbPrlqc504HVEFQjrthSeubus/jzvEDEVGcoxVcT7SqjGcNqTWl7MzNgsBumFLbGUmUOQakpI5P7YZ4D5wwNUpTBSDve3Rca/szNFgXAXO28PNUrF1HInFJEhZuA/Qyhg/bB0M5uGMbBTB7juezSbMYFx7kliJ1CpNKuuaL"
`endif