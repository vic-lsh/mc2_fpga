// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WYWiFwccbkmceem+tEH7jezKkZ4j0yWbDpbStY7/0HaBHiQm004lxCpovjKe
5/Hc6cBNW5zf47ZpuXoas/qEtbludN3reSgHQcX1VNe73qVtQ7iMgdnVPs6C
LOIeb8tKg5aFSc9Vf88/0uHSAXCDacTCq36e+k90EBC2lsysunAI3m+Wdsgd
5c7QLSrqK9B55Gj1pTt9UX0L9EFZMjWd3XyC/gfDqCefhH2UcIgoHQnkLlSB
j7JGR5TrAeMUVoECgtu00pz/V3Thx4sIE+CLFcPtxPsQrWxTwbBPpdJj1dHu
1NhKjvg3cUiXosWew2ORcVMNPNuW6Wyc/KpuAFKDYg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RkzINIl7rd/BgrPNfLYivJNPS1GWLEtNoTJEGHM2BLhlcZilZvz9c/Qb5s6s
sC7sYl1jC3cTKd0ePZr9yw2A45VluzGfJ4ZU1Pq8PRMhkDEaZ/qyQX89CUgM
DWXTMiWByuZuJCaeKtez+lYwz5rMP3qaXYjGgHjJvhq+mSULlcVHKqDPU5Wr
FCZZXaH/ljo1zk7NW4BQ71lnt41Qe7NZXmqkWtAF1KhDz47LODdW+5mjdh3O
PGXxM8uG9vJ/EJXjT17kPJhrxVoBnCTC1MSrZtVZJVeGRubyYiQJJuZ8dBnY
wEX2xA1ZHwCYVYdRIBaCbyXt1LF0lQiud6zed0Rdsw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VhETFfEOW5CF0Y0q8cwaCQdbf8PTtXWiU/Vn4KimOvEOKGgAc9SZMLDr4+UK
fmPnlntl1cyLAUrKP44NfKAwhxKMPCk96L7gKr74hNbkfa0HtesYK1BKO1W2
i1jn6066E6V6f7hYBjLn8o7I4mhnZqmr+pU8hY7a5MyONtaANXBO7ApH7dAd
TEwmR9L/MpueeXBfD1yOeGDvyd9ylSjyyjxPKzxbDovMlInZp39OmocA8AeS
BsWlUVisxKCHsjFZmtA1FDooi3igznDBb3N4moFvISnu72Jn1A5LAuRP2/rA
txa+U7JqyEr/EOOyPs4k2U8Kqi+mo+9OUNV5sTFgtQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kasWHbXOg03b4E8xJsubmdvLOdI5cWyY7qMKzWticIcnoNY+5DCbAY6I9UXl
gQiseYV8LbjYPigAn1X6K3c9w1jndXwjEvXQ2X+kgD3A2h7TQuk3u/dWq07t
RZY9FMDdF49Dbjw2XFgLmvEbhcHMC5ThUuddma3P/TgRRIfKzFP0ba2S+D9A
aZ1SOdx/GKcbJxRm7tfipDG4zVkihjOrR/Yflv1cB9gAEW2Aczf/yfUraeIF
YXCvI2OSha6YSwobctF8AVEChJYcbhaji/Qem5YTMYPuv5vjBwgTfXTFMN2h
XAQq9ETZhLdDQ3qZzVCsq3x9k4VGQQFkUED8RsUPFw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JuRLTZBtd9PWo7tVdtMhzPKRbR+8+/3rq6eBZ8RjQ32cpTFB61XVkBoS4tTl
gBcxJtqRATb+jDmQZwuCdy9gPAU40t2N52Bp4HS1KY4uyqkegUnTcHz801Q5
xgfPjQvMS6t03M8WFCc6eMX9CKRiXIA4UQSApUvAkMpa7tUEafo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ISlSapNGYOvKIZWNhVEluaKUvQzoz83ryuChUhjjx6gioQE8KpzR14ECn9Dy
HchWozA2DONZGFLE59e33cKZK23De6nSAACZXXwMec5h4ihVbECPmW+oVrzD
P60zejWMBti8DSaPpxa4t8oWxWN5/KIpbtSIil/JaXQBIS06qRzjrnQtoF7T
ihARTXzxyEkjHEhxqK5e+Rs7H0VkyDaMoMdxyso+0+VZ6zIHPySo2v6B8V1H
/rWYYKLN4V+JR8VZKiXXUIDKOEmsJyjDE9Ih85+4ibShSZzon6ZW+CSBm1Lw
L0+rUVbL/Kl1b0aURsZPLN+eKXlhI8RiXVN2YOj83RIGMxVt03Dl7qwmnpVk
31kGP40QzP5Rro6Q1r0b5ntAUqLFLMjlfoJITIhkuEqy1oZAweX4PFYubq3O
dKdriD6wycF9xwdPP0mQyyllm6xmNvYdnaie+WNNhWof6I8yWZoWd1lX3jK/
Szhd40Ig34brnwdZj31CVKiE6O3muZod


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oP+Oj3X0sgglTOWH35/z1YhauO8Sl5a4ZZnHDUb3T/5Pd8yzPsFGuUXU9Pd2
l7PPcflbungNFwdTaBRQ+q7YicQuOVjVJFEbXrpKvwDGswh55GDeaUOyvsXg
hyu1rT1z3Hm+UqyhaVruAWc0jzsWAYU49eHqQZVZPSgL3ezSVZ8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bKWcZaafA6f6OCmlUyfWSCXd/nqGyBaxHhL8AaXmGtEFSkCGDS4jMqd5G94X
O1euph7x88qBe7bboWa2XfcErIVvqwB5QCPoKn6YpAzshKX5BN2JiWYBw2wl
lyIp2EYLTvZQA+YLKy3jFVKoPx+HfUdFgbOa72hd0dPfGhllrew=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10656)
`pragma protect data_block
w+mV2GbJG/iQJTzSyWo2Cz3LieSGk/jyBvOJdiJTCr0UsauC1bisEeF8S+cE
7JU2zLV0e4OgmNu9Q7L60TgrwRZODmSVnK2FaTnDGlWJJhb8iUKeayPosBcD
2h3qcMgv9kVmeur4ZGAma5muvpvnunxo73w/uwjAiqQqtvVGuG99xVlAnNzU
Az9rI6Sfwq59NtvP/tzemXhA8trdH8tLrxdasGPsXLF/sbFLmcEMKSvSbsxa
TLf7Cj6rwoLaXCZrXCQZx8eQzaxks5a/OSD4zggoyE5s0vyjJ4DofN5wnqsG
1yXK3DTqFJbh3VsIkz07ZX9pucOGyUr4isUAdShSukIOGIA4kYWOMk1Wp8Le
RNmFT52Suz0k4tTO2/xanqstMDdcbYva6RZbMApa/proe7N8ID9WfUR2S72f
C8bTbJbqG5upVGSt3NvLeK2uOUFyvAVsNHpHCBacceKmPk++wcn371Qc58aH
0hepkuwgzn1iBsD+7HFLejczTSqELpmEg5WFzrYGNZoBC+nDnblAqUeL9vWY
sM5f6/LD2b5bFzwJsY7hM/T0s8G0nBnhEKcPMsvuD4q0zz6DaCZ6u9Dz6DCf
O8Bymu6YbVG6N1wZxj5S+5AgrlxhbGxYSIVqUeFN9OWFv67ubGPQ0tdn10vN
JhCFAnUiHhu94z/MNpeYYdsbqdIKrwAXgM8f+hjSB9bfyDX0DVJlCBN21j9h
2jGSaSuWGcJXtg0w8crmbLUtYe9rrRwFHc+KOGINF2ji+LrUBiJH84ONXlXW
e8hZHVojGQjmXmMMbUm2Qvo7vBTrhC18rXmweXXWQ/NS4a1nnBm7eSVInRyg
2engIU4hNMxLYkBhYkax1nHJN6Q/iIsnwKxJgLfrd85iuK59aBzjdBLCxXVU
SsveYraPZ5U7EcEl+qixW1U7x7ygUPag3S/zsl5RyiK/DuZK0kzbyaBSPiee
Xw0A5N6WtR2vJMmTc4Nn+FB20zRh7lt9bzOdwn8JJ+k9d5NMirQ/ZiM22Lgv
ToRMJhrTrm5s+/Y2lSJm+xUtTqoM9g3fKk46JobofcPKFuDPxlXcgc4M4DA5
IDWSmdT5p5pdo4AQ3G3sYapCtujQPSIo5bzpkABlVt9gCmgxAuuxLUhxqK8V
FrP6/iiKQ2Z7n3q9pQaBza1UCgPHfRfjHpQlok7lftc98cETntFEeDlG0CaX
hXONr5h6K1TXkV+/6rlKSdBYAywOvGkkkh/lBl6tzyyZESZYuL6TfuFrNqbz
d297hI2AQKUPx0Uwq2bdZgfhi1oLSbGxavlbH8OH3fPnLDtIlChBxq1U65Qe
jaxVZeyC/IdgU4ZY5uXQfCqi1DqqCsojdm54CPaj6J2sW8JlNWeZx0jkiuFb
bM3Sl1/4dnAgEPdYypW7CoNE8Z8kV1Ii0Pxf/tU+lXXMoWu+8DebhTAQse+E
VhS1VfqwaNojycCcTqA4uKakpPWY6rk1YG/LMIOFSJRTKr4EDlQt4fSvbmdU
WHgi3FpT2bDVJCuczXVgcSTHKW1InewbXcLzA5SQYQAEQ2v39Xj/CTZPh1Ho
YSQCaiGrSbQlgNaG6rmscU8RGGWjJKiBK0VWlGfL1EI/sovAVk5px2QqrNpS
hoF3NUrk2S/+0ArME/xWwS3uDwP1ETICz0g+GS6oBqOOzIYd65TGrVzPXMiI
O5Vu8TUq1Qulqu8Yxkr1gF8OydC/PijSHi8XuAlmIM5OeeZ1839CPlTK0fnH
gWuzQGZm1xUVLvwodKDnPCFFqscae8TTFHRV68aG4QrbO01Kc1UAMVKrKZVw
RMuMINmiBRSJ6MhRHE3YRx0Xui9HKYrfjIsdurvrY/3YO10hC4cuiOtHgG5i
q5juGf/yS4JYvAVkjmP5kFModSlt9BCpnX1jk88DuA34E1FUM2fPCC86qXoN
4Qk5dFWDtBE05fA1F1N5T+AcF89VLA06zrptTg8CU9ii3n+6dLBGRDVHI/lu
Wyi09rREavAXwtkkdw79QN4KP13n5Kh9J+AnqSXkGcZe/aBbBycqvyB19XOf
nBvRO5+MY3lQt0E8MuUv+QoaU1GSzZX63J6Y9Z8OYZyHH0vybN7Khukzd8un
0zCvk+UGplZBAj9+cC7CZBztRv2WfE28nv8CY4E3A1OBNS2F+yDG6nThHkju
4WWOVZBNmutqZCOteFswcky0q/XN2oJcjSstgjpj/gIowzz6X7/sFVSkJRTk
UBCUYsGPIkdNkT2+Ug4hjfXdOYFrk7+pOQR0HniCeJGE+Hx3xv+KzSwbOFXv
wxiat0UoU05pHlWKtc09Ocd8nrsFOpcWqaZo1OGzJpIUfzg88nhQx/LHWD52
74h+IS9+t8z6VjLMbBEIPi+2gcdYPACTIHn9rhp34S+gxH9INrkD5IfeL/+F
JRNyHWAz1d8GI6MsNPItAIYL7u2V7OK3qRbBWa7msq8hdNfwlSLpqpQb4elk
cHChm6/z+4eEw8nrOLd8J71TqH49rR+q9ykG7yO+D1v1XKI0K0YDdfdqqMVJ
zPRFOmeFfHKE4C8B4rBGGbcPxnpLHrzqPgpGzL6CgRMFaYUkmdxw+z47ulqd
N7dWmVZdkGPciaa2kJtURxF8x/f3CMNfZKNDtAanZYeVf0VppjURJCwXN3l7
yAotYei4dpwfgvWth0B/loEaRA//mvZkhBcTow8VG+09pjgE6CWUn0/civgO
f/qwlvSEzSzSbm1CBlT5P99vCP1vUMBmHr523vbsnN6kg54kesKE72vXWDtd
gYBKrCKpD1Yt4CdVsoQkyQNSXG/hcQY/s5B9GlNr5ufQ+Rcio0a3wDCDAD2W
KULr7sROZnPinIl7weiFd6VM5bEYKZ5hAkdQ94hOkxyXIbBKrwMvJPQn3SOr
X5bCDT6RzXxu7iMekLclaq61IVMv1TNN9kMI98hshgQjhARnXXp7u89suULJ
FE8xTiNSaN7+it6m9Hi/7wgcIj5Dh2D/Z89Rjc7MjymYdjyEenQpAgqFgH0C
kFnKVidzkRH8Hk8x8T0rv3eMbWS8OQOiSnv8X+7IYY+SWSVqGreeUB9u8fJJ
SjF4lHk9Ocr6Eq0oKGmiBKs/e9s5CBZE5UZKEi2xVs3Ws7paHrXpXWN4eTFK
cX+/qAWdJ2812K2ciwMYixtvV1Y6AA0Vtt+Q5sMsPEEegZzhobd3SKwM4hGt
ftmfOXDSF+Zu+nf813O7n44gYsr1ACQgmDPTzCu5ael3yDsg0FmmrArqCoMc
hy5UEVwogKEY3heXXcB7Rf7KP6ddQhjxH34fX1zEQcgyngALVgVKU0IZuFc4
mSaz1u2rQ35Xl+h/5K79efPFTUe3zL7Kenx/1xuHZfUydKWmjzzeAYrF/VE3
FCWk7njd7uNvcp4OKx33MllxV2FCk8bpyfiEK86/UdTuZtUkkhyYvycClfA3
E62ag88EFZ6neGAXbiQn8osY9mt24bB/tTFXr5cvd/305JMjczsJMKKK5s62
f6vKe5+INBikF1RPaUJBp4i0NnlCM7cT2lwU+9Btzmh6UKP3/R3x2iQiWngk
X/rE5vyUBX4OXqa+Zh31W84FNxo5/0p2JleF5LHZG2fuZAq+sEr4ReDb0tu/
bhYr0TLUv0X13TkJ8GQCOYsxkRD+DYG7gnp1zMjoC5TWJ/YSSAhP3lbVpJG6
3w1c1xLY0JM99koqSFYmWmMqiuHRUZp3QvEQQpQOaokJYZkAIhCG767VPmx3
QxrgZhVzUOdW7aheIiYY/7uVNkd/qJCcHshZ8o0fcr3c5KwAoFSHPA+rwRdz
S0aIUsdWlm96019h5x/3Oe85ZqoqrSgyxXdNMa18NXBeXfzkyNwoJPh9wXab
pwLktHFDmqEvPBs2ULIkNSt1tbBL7PRzDkXJRRkDoA7LpYVB6X94k8inbbh4
gGzpLHBCyFOeVYnJQbCydMXSgsz08y9unqQFpEZdt/roytH4WxJtqp1kbdBV
P7XIoo64QjKC6R5Dwg/GiQJul6CpJqGZAOu2HWqP85aMDM9i/kxwds+t4x3M
m51fBW4XtdGl4Zv4jxdD1vaRImIgkvE6YxweKxmGP6EVDtXRxWTzHYbEiGaj
x9hnm9ewxvTVmoKqPolMvvJsdg3f6p5oVyHq7Khf1dnt2VW1T1ACWaBhDNfh
EnFTHuRp8bsA5qdaJgPcFTljaKCTEioiHLak+w8o6n9NFUxDYAaz2uJHy/RQ
r4zGCls7U6sl1cgJSIq5bxnAHJgCif/axzgtea75njZwPLpFocjJLNSOLkh4
dy5tsQ0tUkn/xLgn23tOMhAmIhJqbbogcHkZOPKPZTiHa7P0e7kN1Eoz3fAO
6wz5zS36dgtskbgX6ExNMLYcB5pIPLkmebzXzdNDXpSzOHmzw7I7W08X4SrE
8dYMmMARhFQVxL/QRn80bfF+0koS3cca40RFgwZ1j8RYq4vJqirA4Qlpsjzf
nZ0q4FBXA0WZnMT8ceb2+Al6QZgUwL5mW9Qtfww/aZezEJTKDZ2VbTNT+9aH
TvFVL33YGQOEY2r5IkakQJPddqAaCJ2Mdv/Xeum+PA4uqv1t+b8UawJKOndp
rudccv9DXrT6Mn1ycSJ2Cv2oNR7nt7w0OoxwDCi25iVu2LqCQGapkZaOLj8b
Dkcb8j1EnegmVthpS0xE3t6VS9WpTfqLJdX3rsRw7LzQoY+ixXFjMbHfaqK/
Par1+7Htg5/sljJpcMdb41LuOiygwe+TcobKr2oZbWfaBqsJEGz/OjpMpScL
0bkSrGqYgwGkGicVGSadiLj+TiECsM5J+bwrGx0CXJPD0ey2pF/oHHtghi0S
vjwe6lTdd4XDq3Zpny4UUSkBqyzAsorN2ACOSVApgZuUsxVo/wr2fOhuNRsY
ujKRn6SgrOFZVvhJsoYLuFBJVWs6rUiGVlolusqUxRR7OtCn7SY1KHE6lArS
iPZ3YlCsYlbbgxmId+KbqYzhN/a8XufckafyJDPmfqS2x3mXzdJ8GhYVNyHz
P5d9h12FUimoK/R7/o6ZvK/NMW3wGpbrgcCsxdp5hVbkHl+tr0JM6sL+TIXw
KZ6mbrhE8G3TgJZPco6Q//3LdayIukNptPPBSFLlACm74IzBkmpQlyzVMW8t
ABWVMkCfyQlsQdDwa0IZLGn1jDYOcjYMAR71r7WIKP2bdgibCEbE/XL5311N
l4hl8CYbhz3LVSppzfzsYF1eYzS8gNDduXOIaDzqgWHrrLNjvGipEKunSXwx
mYcB9AbM2PzMfO6iRfkXyuJnwl5qzyevOHw3b/EN2WJfxUK2o+UAFtblLshb
b2k2NDCuI4wl3nFLcew5/MgXLR3TWQ8Uk8m17DlO6CIzHIR9OAkFPB9Q8HWu
etXV/DOo7+/hcoiQFoSaOCPzca0haw9fn6k1n+ti7z+kYR1QocCYW97B/Jpp
l39udCqxxWhSE1NyglmnbyzOsXqysaj8Rhv5Cfp8qVVgBF4LOLqIhHjHNmrn
cfywBSnrME/L4Ys/5IV00CikjymLcvzzaB92su841HEYpSF+OoCGgQIfRz4Z
Jw/dPOzNh/hBl2U5ovKTqRdCoP7btCpvMPr9mWcTW7HYPy/R7vChCLvBLusM
Y0n0hQc+m4murKnGHg48JhzkQFye7D7KwsV7ByNp7T4idZ5tcBalSz2jCb4/
VTJPWLlJqMplDf1Oxdia+o4dDmkX6goV8pgorfdlf0StKdSRjZHZAyUOYIAQ
qBWAg7Qths1X1smprdV6prIwbSXt9UWfI10xNuTIrCgBU4tvVyosq48cIY1L
QRJasVuZp0O0PtRzqg0RW/qMsgDi/0QmqNPppZeD2Wsz2RIW6zLAC0ibSMg8
cKh2GNjwdyzxcoMQAK7wqx1rC8RiOb42nWbrz5yYy1ssyAG45Z19qiFjLNMG
x/d/sQ2jbmYDJxP7CZsd2uWDstjzW0Y+MxB9Kpd52kAZFXrH60Ifs7I5XaGz
UAOoyBSyB9d7q3TV2bYei6tA6y+Pdzq1vfM+1oG5PE2wpPA8HEw3XooKCJ2D
oGFDVGx2bMFGPNpmVykesVVdIvDFehWOaEddYQ50dlkjWpbelhy/9zYKK7nN
YRkN8iy5Rn+633gFfYym9/2dJ1xrezw08zoUpgPqrAs7GegDmcyuR/vDUY5n
/ZUeQm5c95SiMUXHy0tXNdOk6QEIOXr1oWYwbU2WGg9n41F0GqipQO83oapT
j1lT2Bz6xbs+gX52skeRxUvqL1YJIQczuZ7PzqWrg1SVRmC5jKdf7OpQLWHw
t33IAgvfK8KN5BAfEFrhI6Qgm2GUDkVQHUF5taX4RCLGCU4el9//BKBTisAh
wqXbqKBXdJGfYWPC/fxQQaIVC+RshAimf9yBgUSICEuBuR5hktZpVS+ahyjO
LyqV2SX7+pXuj16h7iiTFJnwVJILkO/XuwADF2yipaKsdy7ZTTP8ver32dkM
e0d/RifXGWfPLOl1GClYtQily5chyRvxSeSr0VhdNk7yohnLwbciJtZIpcjl
aapouXZT7EzqjKSVvcLiV10D6kbnQAb0Vb0e2Od/69oReHykNEnJwC27/pYQ
mJK+KqnB+5Gz0rAW7+yy0Ef6Hzy4WdqYpjjylhapiTmhP2716CVDY6hkDuay
BoYOsfyonj5GZ/Pcaw8VIk/+qOPF+nApwxKpRX79BPp6ry65855XgAxnjR5w
UYI+NMrlzHHIPzp+vokOsFW4EWS3bXbSi2emP+/6TET1j3F/Bf+L6ten3w0X
p62d0n5EOWdgTsgQm+d8UMGQZ5ZDo151AUmRKDV9spv/7x11zDGaBF9X/3Yv
YmybtPbWx0Stc15kVOxNxBhCI/mNsgolxv46Ze+26/XIv0To/0sb/x6b1eOj
W0xYeaYprVkM2R4hRPDgGvluvvq7M1Dy3Y3r3s89QYXqz00OWSVQo2QyJzU6
HeZclYxjiXZWiBXYuOcjOBKCNnehLiQc5rWnBTunrDUCC5ssT8/SY7YIukkr
kjBXqTtGMDBA81p5Ha5pquMOrmrZacOMj8RTAFKh4BpqCgJtyDJOcFk9QUnx
JA6gx3M+y7yccLN012FbbnH/6Yljx4drK6nZrroXbqef80nijt4FVXc52BtZ
dMVKKD0D/IgJjtf9EZ9OK1408cLXPToOPWEwQ14gq+rVYo5zC6TI5XaURlj+
AeUHc6ieqWLXzcud2AhYjSHw2CxalwbcUbZSqVO4in+p5cjZTCqGHgoTKvsw
z0MRJWVhpUwlQsV3jpUFC4iXoTCy1FNHTenPqwKEKfKOZEVfe6OFL6QNzD3B
Zgwmc8mk03AYGr1kCU9Q01oSgKrwsJC234xYuGrDyrvicF1KxLLbMsRVOBfl
8Su3RadTd4ARh9DwRICdCfvDQzC1Q2ocKpt7UNKbV8HyTDydpVk2Z+XI4VKg
QW4IChEP+lkb4V2cw4iBxuYwdvVL4nkCHc+aw15En00hsS6DfdScOeXhOXc7
TksE9GI2Vf3pfZz/l4LaU73Br2bQfhi26xDYcQ4qNRH553G1migbOccTjxup
e9k+hEpVOgfq/NeI+dPdA6Ce2m3YIQYUWDjW9l+wLVK+YbFEpLH/MRDXlhXd
plHdmbw9ANMk1MoYzJNg2QNOg/yDxvazygjeYR7oOx1N8miStMUX3rYV4oiR
u7yxE1bzmc3tfycVn+qlst79iNZPgc3TDfRxoyRwoPTy5uBkgtbc069a6UPG
yYTdncNndKlvp3XfxZBxGT+trwHRqV00N1AVWMK+oZYNNCxiybt0dThQdMXM
FWANrf129lHnRvmlid3XUWnV15fanDWd/Y3ovR6i9k+LZiRCKTUVenfh5yvs
fCuxZPEYa/lsqp/K9xQH13HCv3oFXJR8MP3mHR6QyF5y3zQcNnQVgnCrJdbj
l3yyLWiRvLNbtFuZAZG1qUOKEjnJLf8aXh09G89wl5aFTLKj7japBH/vTR4U
4bUB+MXIEdZrATdnXBFze5YiT4V2Mk6hNFNWXnPgC+tI44gRS6S0tU3+lRez
EnJ5yl/tYlB3rrNVJ4wba1/ek6W3Ze757XLWuy5xxQ2p2u4LTnwUcBIm87pk
2TbwblvPasZ39uREQmlrLyjju+7WjnyVKrfd91FU8vlSuE/dw5qEW6U1HUxa
31N1ye4Rc9flwqseloPb9sdZ4gNg96sBIDR2Mcc3hvBkskKNB/6vAOFp2f7r
MCV6/250JBDUkRBORx4YEPBhPJ5ueOssOizyTyp8fxAYes3WdCxS73AJGmKE
Dgk2Uu877TNDTSGZ36C6D3w7b/v2OG4IVy7G/v3neG75SvKwjC5zhlDjxPkp
W0JyEwfKm/YIpNWXYVFMzcMU+z9XpGTO5dQx3k/AV3xYU0Ncut/YL0MOmsKl
S6BeFHY6762hMepybOIKggO0U39jPF+xAks+0lftNXgr7Ss/Bj04Vz0G5kwt
MKTdJtey0sv2EkBNfZ6D2nWKGR8tBRUQcg0xvU7aW++eoBfBQJ84ogbMIPvJ
b4qP5XO43spZFQdq0ZbDrXbsIx/JdlKNdHQeK35trOp0kKdohW3lpNE8zraM
MeizUsm5hRVye04kgh0YoKRHpKo807pXacPwb+ySxQXNumz2fQjiCpXrQ8sB
6XKRdc5vvb1f7f5Jk7oHunmRnpLbsSg7MN8nyAM/WiTo6roAEuKKTj0a3Yd+
aTaWNPWmPmG309Lk95im7+OIH+eSBmYZywACoytm7hoNXNmGaQ4kHqHbRc6f
a/6NRtaCuypn2Vs7UDY7t1X+J+KFGsVmnDdHkUFYPXB0lPF8upXYQeXTeO6s
3URKgmGFs1qMvxDMKB/bZHoot11hQeG4EVGRHkIlhbWqm+6TOnRR7jXfeeN1
GBcQqalFkpSGn3F5NmVyv+qwBmaEQDlEyIsPEiEEoXcPErnhczqpyWFZyCzi
GmP/kS5ekXhjm8pszKmKibMd2nswDJZdyvUigIBsx/zC9BYzkMhjIG+3deeN
+SAAOCBWMyOT1lVpwtmIssGbq4LYjZ4AW1eqe0XP2i8Dt0K6gIwgYxR/bxKw
SS1Danli2iEBidms5CNuIkY3HA85kcDqHHWxiaLmbR3GRHhUq6WPfgFHphVA
LvtmzMLNLFFpgtyTJVf/TOx+zXPDE5jHkMOw2hnDx4+1wMkn0pjnb0pz0Hjr
QzmVTXK9k4CrGMAQa2diZpvMItxd/avRvwWuCL0nz11JL9Jc4XfA9RAQTcs6
IOHH1cy7PAsG1aec5ofEVxkNM5IY6JfkLTGKFOQrw8OgZqMQJN3YJUxEjLgK
0YzKG1W3/ZPmgRlDXxA9dxYv3OoaaQGIavO8XcabkWpL51AsbeEe2TbNMYQf
qXf+yjYUtIaega56bY6+/Vqpx/lDeMAo3YCSBgs8xaV9q8C8JUHg5TNfEXsr
cMEHCkfKZCapc2qpQq7oNPPtRvQcJ/iwBco77h2PtxXDhS6Ht/tRn1bC+zKx
6KC5uSCeC0LfTSIuRsnBunxxjw8St1WogWOVslh+IUTGjigwQ/Ro99H4WFcQ
AQgAkQZdphKRvmr8ugCTDu2Pc4K5AE8trJ3CQQpq0krE1hC3nji05ayeOoLn
PjgXdajlLJQq5jtygbQUwHp7H2lBRRnm6biVDIRhrxDMQ6FeIpG24D8cyv7g
uCr8uloHqV0vYS0DmO7MbTHaQ6+x780s8eYp0Nwpol6HPUG4bq7jciMMHWqc
39osAVhcWyc0G0bDNVyFzM8v9ouAWXi3xAMg53nq/75h/Bss+MtHxjguf8BN
hS3GUxdrohI3OVj4IvJoADsV1kXyDkCif7uzVWezO4BDft0ljI5YstyH1POT
Rb20TZLfppTaMNO+x/qXFuSgcNFN1QOVnb7MOlvPmxDju+JxiUlQkq1BEb0Y
z0AxJgbAgKgOWdH4vMDGZVhKorZVraD00uANXOwvjioA3UAXSaQC+8WEWnF5
Iw2x8nLC+S0xZjsMKx71DmEOIen9rvTR3Gd6Sfzeb4o30HtIuk5f6N4X1Er/
GB/GSjBy03SkKQxzvqYMInKfL/f/sEw5/5+eFfnDTXFSqzFU/dDZ+sFts+Tr
dcKj5EDXYbwuJ6QPQ71MgkwlO0RCDVKluiN98wLF/a3H99jchTtKtNkaceg5
p4QbZVh6Mg+YSmL0OQoadZC5DysWK98NpZifGVeweAOHZMSPa8pGwM+kXHrW
dKICFM5hI+YgB9Pk6djhQwq1BC+B2zaNi7qUCRmv8ghUJqBAi/P0l03LzgWt
GN6gCqOYgzvof58izMV/3L2rI8TgPmWtppaVpQq3y7XNLNOFnPontyxFfzbh
AEq5jyg7US/X13P7VyVkmd4uxqTaFXLumO6N1Y1v5xZqSQvnXBNX+s/g/ki/
9hpchuN86z0BQEptv009PWhG6XxH7pjED/XO40mUjqYJdhWhNY33mZPytsTb
8u/bW0n2d+CI8TX5xY+SAHxOFHSlpJmudkqqAejXqj+/V9bfpDJeuuWiJ02Y
4IDoznDWLu7AH2Y6Q/LAFZxbjIPjYzdWJLuJcn+bQk1x2t0SjQNq+/hpjxkI
FSdsos6CiGo3ohF7LA6aUDdM1XwF+B4B2te8yAFP+9ei0ThcubmU8GMMO92Y
3Gr12/165LMPMla+8jfhHc8vXau79hz5D4kLZqqdVGVT6o7xo4Wa+rOrYtjY
yb+YGqEGGgRSNFnu24FADR8S7X5JK0YKWSZOgj/FuTUm624M4jNPH3n3b4FK
StUvRRt2trOJLtZkxEGnM+gdCuckfNDJerZJrofTImUS83vNXMaXr4uqak5F
PD+c1+f3zadPi7OPymHBLpDvpUhKwQDBdxW+IMfHotOTajGQ0ROaRfBD6Foj
nBukArfBWw7JcDv7maIaLyKVWR7YmePiKTWphYyMs6OAJZdo9Qpmf5HhdQ6j
jvLEfQ7dfAiD0NphL2n4SuRXIrgiJtWFo5/slKzKW+Q8ryxVNhnSHGvm/KWp
vWHPPAuEJP6p540iUtkhheoleiXRknsTvT0CvT0T9icstxS+XtmyeTXboUbo
rOYhbah33EVklhR4vG8REkHAfAO+nGtYwFRf8q9qZZYnvgGIYe7C20f5d1MT
iXY2s4JKdynP4SkCWj7QiwuZbt1+TjtBX0KkHQmrv+ZM50HZCcGt+y9Iz4rw
5lAC9/ygnDieugergteZVxHdKHM+1Tj+fvqWuUSlwTiy2yZtZzEs4NbMmTEk
XEum7xE0i/rVptAEg8ptn3zvl7rM0ETvp3C5RTNJNleZ5aDrqNpm2fOeQ0ag
vkQi6OgN5R3Qed4jgBrDInbNK94J3mFCK5Xp7eayoI3PxS+aoKrzSme5WOHL
qvaukWLXmKc3OgphAUBtLJnxGcVg+V+7g2rkrIhDnp0OjGGrqHzy9TclVJPL
kB98ikPnIrkLZ/lYbUOunotXcZNNRW9Xyrh2BTIyP4gbB3h1KI75JlwQ6LLU
PofzjN8ia82Oe28q2JT8ejkfU2aFusMxzPnN3nlJ94UeUXzDvbU/++MPxvul
Kbu4S+/A1z8nrSlW6wUeijRfFuGPPzjYp/yRcra6XYJ7n5NBxTQlb5f/Y8ac
y012Tu1hmzLo8tP4fZt8WlWX9vtDGSV20l4p0x+wFMqi2SeMOPOUvi4sC7+c
K1fImTmU/nAaQhrRLgE8wgpfWFFORG9yKa+1UzXCg1cc6Pmqz/DtQrL5rJH/
Q/WMfiQ6Y6wBzO9xTEs5O52NFN8UUabk5Bjk0ck2EDTBZLW9NaiZuvzfifwN
tGcnVEM2QCO//KYf1QL7338sp7cav9z1BM9SikHR4bCO/zoROiPvGgdpi6eL
QVegGsZfIO2vR+BvpeQLsbWxkNMM4Ev1iHUe3vG+BTplp5U5NApVzjKVpBmF
eYmiNvnF0HkZ0As3eqAcVuCWFlhxtf+rlwU4UGh0o9+VXGgpJ/G9rVB4XT9Y
LDX1+fMTFMzSAFSAJK1RY/SG6oPKLmSmIgIGrMPO+sd0hP6WnlccVzJ/T+NJ
rPBN6+SnNyzgc/oQYXXk/rtcKIDN8XJfm/xqEwOPX3lFzIdwfHcn09sKlvOb
L20SgOyKU4hgd8cd6SO2C+p3mhCU+H8zDGdrDjEd0ot166SsDmotmWEYjKjX
gYKK7/X3CsT8bmJeO7sfs/OEPEf0h7Gat4mNLVB9w/hQ7V7R0Fowfg8QfT/S
mt+GwEL/Hh5GJuxgBY7Kv2QsKzHvhZqgoJRyjPe3DFwsALrFwStktfFQcVg8
UFKw9L8ZEjefiei/sitKx4MJznYmfjoiiGPDlDVlm0jx/axoFvm6XZ30XKaJ
+bBK8N9Aatn6267jZaHGVr/IR5nBes3bmR627eH5QATHmt/4h4inhy8pF0tW
uAOhviVonKrvOqXN5vzhJrIMZL3L01zYoUv35OXdvtfEUxRQm2rKmv7+CAqL
Vlw5wEDTEOqjUnrDrNEPJovDN38Z6id+zPaOGyi7/us/lJEBxdckc3QvQlJv
SIUlTCnhJU/7B1sM7ghWtzOI1DKwNBLzRzKSAakGs5UQEMvse0mMkm5KVkKf
Ef7IEJh481mxDcItVAMwG5nT/p1o4AHA+/NOicur49WJhwcAc6u06tKMg3pi
EncPTx32xT8sa5hS4vOWk4OgPi2JI8oGB47DkM/rS7zzCq1GY5xRe0K41OTc
R2zZBNGEWHjfB1CMzEZmI+6jvvqQyByBVCdiPM5ZbCkR9c/sXD7jQ4OT7aWQ
24q6rc/V8DzjOaafReqnR+01AbZWwLjnlyM6KxT43d4KZVUh/lx16D5NecDi
HTTALybCI3QfxHgseU0yIg3Nj9WH1wOYDyFLHTMYHSMpSLPKL6erqnsUZAGl
A8xZaL4CKi45qK43gTWv6J7kZg1/kcZYD8JNAL97R5+VqDhOlXswh4aoRE1d
idPvKcGBAnDWH9aOgvGZ8dmzYEO8ivmhfVfssmQu9zGsNvZGYxwlV3bnu3YJ
21L6H3LmN+Vtt8IL3C/1LO0kSTmIiQdCrMQUinmOVDWDt8WupZw3Yf9t9X3+
ZuebfrMXwftyqSwaQxqK8gHcMw440vF2QKAcUlQhonc7qblvFDyBR3OJDBD4
codamzSd/LENcTkjHeAr0cIK6dE2X6U4M6wg0cuQ48LdkqhRQsAwN6qbaNlU
3DxkKds9DlazouZJGvdaxx0mNJq1x69QRd8+AdcA4lzoth1qjdhidO7Rs343
+dnpB/1wuWo7FDHvUtFMsWz+F2h4ZjTfZ35hfzStab+hSBhfdlvBJL7S8ZqN
Zdib6HQ8l1Hgcj5kTydI13DpX5FQxSQuv1GbDDPkKH6OJvccSs4IX5cdmjqT
pQD2jxKBuO7u7nZ2kpa7fEEgSFgZO6kcl4aMKSXgVd+8KyYilWNRLBPKFAZC
QVPZO2wo4vxTDgzxdmdW2tx17ttGcUqIjkP1ziXMhSRjGM/NUvwlyv1MZzr4
Z5V8uiNMf4F+jNA3VoJuPY8/PZmzcWWKho+G9Z6sTg+P0DCLJJkWbC7yR0gV
z/8bDtNqP2sNmzQLqAZWi+Xzxw1fnXoyte8e1ij0Dh6gLDOenUGoJ/OsJ3p2
MHlv/49REniXQUnDUJCszW6sIKGX0fnuEaVUiV/+Vx5wHjaj5y2mALUm4ItM
t1A0Lm1HGOkiDRQuYV/SgRNe7fB6I7R98ZArEnY1n8YWPfnS3cUfEfla0PIU
w0a1b83ls33Zb1tlhIZ4TCSO2yDoqSEoZt4ZYpSppMdTa8rDIFwW6LOAJroj
MWxfg5ZJm2J94QOkJwlM/MuZsoqPld4NKjjtzKH74cg+tmxIhpnkV/fI97Gl
hAkubcSJ0jaGnPb3VlRUrhOskZWNi+wCqywb0RNd01+b69GLzxRk86H2WD3h
LFJ7IL9Jix+IG64eYJLSh01Fj9yp9tvG0kng51oBYQ3OUnwC1SG1hlrcEl7S
547p10SwENVqd7dN3nmc0FBmSNCErQRC5QGKFpZ9wqZnGDPwosisiVfCCpvk
kb38HhBUt0muHY/+IU3IFqKFhWyEl+NwFIY9s9z/t4s2qDEFEoXdLImyZMYp
/PRfUKHYmdODvtl1oSS8AIWjFt+ldE1z88weUxMdtuly0OCR8P+qm2mysN5K
ILxisAh3tspMjCZEk1UJUvtM/dSDZORPNyNcI73zwVSzAuZio78FKJSEwslG
RaOlY0/bOUZYNdXAe2nzCFSqY6qCFcaQLJNDZhccxlDmB2P+wkIVLae8ALkw
xjCOIUOuLDJTVdDasi3fgxdHOmNDtV7Pnjxloh9bKh5BPero

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzcJzBWApgXuKCYB23x6xiXwqfVLEgko0/0GXABzRurcB/eJYn8GRigCOMpgR5jca+Nd5Qxk/E8cmm+TNnZpSwrMX8IvNbBBsNqUl7v8LuUt8B0N88a7oXVOLTSi5QC3R1bA0mo88ere6X4Kok7f60I6tkhP5aUurOkmkjXj22iWXeJ+sbu7dsAO/lokczA7QiR7QY8mNR+woiAeoihn+kVScVGoE3u6MfB6uZqaM1vZV0Z/3WXfw0x3GX4QZWOovrM+GjfxFOAYC1I7YOWCo2FWXR/JXQxOtS6PrcskOzyl67s+AMeNpO4oRZ2vOQ09dDAbnq7NqZsH+JaAdK8wbaVpMx7Tzp+1rGLkyxzLRhPtNmixSiY9bG1nNPQ4vOhgKdgyt4J1ei/dCDnBtbsZEm6OW6cRiRYCEue6rAtys9Tyyin2E2ai2AN9zEHt/YaQJbb782iQu56jccaNJx/uicUV3LlylLQ02PQYl6VhhJ77UulEAHMeFlXt5297D1ACjk6DHaIbIWuv5pxUqO68rAZXZVibNYHbzgDOtXA79wn7d30NSS93SvMGweOtatvrMzSv3HWL4UFL4DQFcDjSz5keinPp3zyhkUmGKd/K2g8tZPQs/iUx4pOK5Aln/UkxQ+UvDbY+36fIYhH4qTtibJYXDtClhRNu3bNKs58AUGgXL33YxTxpVHjvIVunrW3rbb6gL5n3FjiEL24oVOSuUFsznK5sE0CZldSF6lBp0ZBs+l2MwCKx9bTa1sIRm+vztv9BtK70JNtM3jvqIy4zIQiN"
`endif