// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UD7rHaW8sVg/P9UmAvogkCg71/LuNTLV+RoUpWVy6Sp/bxCAhl8xc7Ukyk9q
O2XDCtaUjMRePKRhtw1qzDwq9OTzMbvAsdGLT5u8OhXMBVYZbKmFPDYtC0Kb
ZmGoG0suNM6zMh552dmz4WJqu5Ap+56nXqOgRQrKyfXbExpbW8zE2BuA73ij
dWk2MDGsSRABeEB8sUBtSOq9tnwXHGDw8MX0Oq3qZqpAiQfqKPjF438O15PJ
PiWtE+sVGoQD9SdlT6ps6Z5OEml4cqOnOfoOnflkBzcyoynYp4cHBh3wK5a3
EQ2sP5roysf1fxuWZjGJx0MlL7hdrqjCpwaAnnn7kA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XP6a5tBgxgt9G8oqksypOPoIlDNHlkIop9G3qbsDRgK1m4csuybp3cAhch6q
oFAm4c8J+d45bO8YuyH61OVAdhfjV7futv1EWZ6vO18F0pgFiyxr0UZeR1Pj
RxFu8BuAeHlDXf1/I9WS2eFamYCqVdV81iqj2qin+der+nB8j8V4ueAOV745
REyqunC7pZdqN/owMKhvNOFYmAlpY3CJjCF4eiUSFlL5JJli8CtZp7MMSfj8
QymrPvKge3n3PlAJ1WsFjXhKQSISMqGkAdO69KG3IiRkdvAldSNDnIR4ALU2
UIm7oAv2kM0GJV26Yxt2iKePRYfA6j3qRT6U6WlIqg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h5pWf+zQYB6slnaXCj2Zq8j19tsyZf3PQhNEYMpr6r9B0YbCH63ZC59wjUij
hemL+4lQ1G2RUJpLkBArnuWa21EHKFHjjJhk/Ke/fKbBmAs8x9nhIXOJKJR8
i81LrPiNEcXP4ZrT7p1NrBrQ+L+VvC3Nwo/cphcDSNamFOoRorWVY/r4odzo
4Vgb36S6TlMjM6qwwuJOVRQo2B5QtU2HgaDJLVoTOwfzjDC3fUIKnNHD3ilz
lJ5Id2IqxPn2t5ANggjxmXMTL2RaReuW+JMopjlDlPVilsLTDVUR44ve8gcx
6tMcXPmawHeYCNFQIf8sqhGYQO6QcShKFHggC/jFvQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KcevPsD38JCYyTO7AFvB3r1XJnkD1M2IHyekHrGG4f2T8IUqUuQ3PVx0u3uq
+TOAIS1k4yDVOMl59r1feXUAi1h/EwL3+qXwx5Ph0gubfxU2Ci7RZ6YJsL7h
xsgEj9SQkZV+T8ybjVtvPYEjfzi7EjmWygqY1k64roc79kH7k42XcBtqNaJG
ihN1VTD57wdWhPvInyZo5bAqk250PaFQ5oq8+yEGfoTGIDIWx9yW/3AYUS3M
MTZuKVMOpGA+7uo3R1eGHx4eMog/PTbzssT9ymLFJhdynVJNNKQn0CkbT8UR
ftPvo7lMIixHA6brYgkO6Q4Vtify7tulffN3V+Jrhg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FeFPtma4O8IJ0X5jjfRRvoB8zOBR30u0eFrvUw2+Awb7+R5s+HQYk82oPasR
ltKp5lv+q/4btomw+CyEcoAPIjkzRM3nYNIE1iObzD2Pj7VL2LXRakMu33Sa
I0FBVMXzBbbpd7OE/TSYbWnHN2QnrV/ATXvHFsuymUyRQ98ybZE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
st0QPpWw7bgKGzCUPBUl7MAOyjRH7Rqtrqj38DZkXNoc3oq1RmIet4dCs4SI
oRIILOOS4xnKTzh8tPe/EaA1WajmduC3ALvKaQroKc7zqem1mtZE5MCMzUQk
5RK89UIIRNkgQ4dzSd4FgMJxS8mI2+UXbA2w4U7Kvef+coKIVfg6FTsHpHGB
UfdJu3NJI1c5h5TeCXmrA6L2U5iRQ84/qmzssQuY1FK+y7/BfqtyAtF9efb5
qogkxVb7T/xh5VWWZoTaSp0iJF4bSs8oGcw60EPW79CigOwoj3+bU1Q9lSHo
4ZajN8mUwxZ3d79Wt4oByHpN8MQEV4da8uJ2fJw5h3v7y3pPjfQ6Qs9NVCOq
EppsVibV2CKmjcotN0QrhOY5FPXiD22HQlsifin927dMKL4Q77+HFsskqpuA
pynujUp/k43F8dGvvFG+o9YwOBEaqQQWCVq0uq1yBlVu0kZOvMQ7hhexY/0s
m08C23aRIddC5JdzEmp2CUoPGzSId+wz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DGOnR6R/tGNXv6oVNPNaCfGZRrUVisP90E3baB7+FqXgK85TQQUAeWlBHo+7
QIZD7tnFfxT2cRzCBPiJ5aiPUmA4CCRqsQK+vAt8uaWVvuWoPdgKtvXipxDJ
eB95GDfXVkbVQzyL24T+CSha+N4MYBdavz6VBG8SYYmBk8VGvOw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IOVfl+BGpkK08ZugLrmzIv74lPAnwiqDRD0Tf+5b/VKE1HEalYu55gD10EMI
GmlsVC4m9uEQNDbno9u88M4HxdJGLA1lNi4esrL+PrrpuXKIZmxgcdrGgUqI
ED0BMBqaWL8Bt7hXGz37f+4N094sE3drTZFz5d1jXWxtcQr3Bkg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 56912)
`pragma protect data_block
JEdcfH7SwFN7lGX82JIWqYYsicFXu7xBUVAKOkDqKiWv7jgJN3sYVqxMfI54
5a3vyPh6P+vZwGCx4C4PHYHnwlLvOJsmajZFnTVBWNPGFF35JfUCvAkJLtDL
GtYEGJsIxGSB1sX/b90kCbd7dZ0eX9hFgU13trdA7/criE4whPB/GzcP8d8a
JZc6ZxjbFUC/qLG/bR7wz9/JXKzOZoun2q8w8wGQdWBc0zFrHvKqFHmHbxz+
dtXrmzFUafgNzwYC+LP812mKbUSDiLsMmNTe/sxTD/Vr0kU9O0ko5YeY6QqE
E3adMVK4wR15UO7M2ApowYF+AAVxy/8hbPIToCP8KrzvlSltHnByiKSatVKB
6+bEXUTTLDaa9FAxnS0kq5ZHslvxKKsLtlmVDlGv5cs3jza/nDJHp1FvEGyM
HPH0ELyNCeAKoqOIKCZ02a1EWKxo5+zFKQbMOFGr6paum4ocXsLuVvsjUNzU
96aq4CwVs3FdtmMcf2LRDfiFADUmkDqq3opycaXL5yr5fpyReeZF+wU3HMeb
Ln79T147CCV4btoiKJOhwJJKhiOuBlK0ldG7gOlaa/nNAniy7Cmn2lG9bli8
reOLFg5+/+xECJHGKpxh59eUfO9E+h9OCegQjTIy7NXo5kMWL53sQ4GVsXNS
fHGCYJ3/m2AM93GHvzq6awhjTvKvUzuP1ld6rsp0hc+W84iKxpsZa/4sKPLQ
3OL2OtN5ciHei3dGfPiBszq0RyD3+O7USqQIRWcLeiPMi0l1r7XAVIvHafzo
WB8tZZiauKFmBPc8vp2Df85LDXyXB8P3HJ8X+FYwhr3NKLOYlRIaddy8mNPG
4hdiUpdlNaSIaMszNLz8vTQOOaUmcNPHcICj/hXGInquO5NQ5E+3J+q7kq/F
L8VX/3mZGyKKGVirjKZSHbZlD39OSXvYIqSyLvcLLHbj4rTK76e+a50fKq4J
Ngq5KrR4YyR5k/ZDrIUbFvzcuD4PalYGr8p3jn9j36If1aeP5XW+7Wy3D8PD
oCBahZ4LRih8EfadsLGaJu2HVG4avl8nFA49JKQddZb2cnnupLZoEdDqk1G/
qi7hqUIEGiuSp2x6wBoG2Y477+aMqj+ERhnm1ChLB8wPjG4dO6vUJKPl2xoN
SArB74pQNfMBFFzK9MBr4gyhGJ35lyTUaijLVyJ7bbHEySWKhgN9a5bUio6Z
m3nvHAiPLPIfxPlJ+qFcMTPlFERXwIlitUv6dNpd2KrivepxDM/Mufv0GTNY
fjgnyy3fBP7ZFRMQmP7oGEOMfSj49iL89xzEXw4JxWsK2irMdcwag2J/582D
tl0C5kewJBw+R+/HAIy5ukHLbHEyNf3LC/VBYAGBapWlzfgUM+zBY9UYKgHq
mgtK5P8/V4Rq4s0SmV0fhUmFiyTsDteJ2ZEV8fGHdDQ5wMD16vgkVf/EGdJm
RUt63mivYfTIMuqhPHEaRoF6hrgBD5IN/39HgIaAKvhSUz8kIqKkoH33smZl
LhOTVag+kl0cpx5yyxnMoxXrRdtNg9SDHXqvoqPttq5Izm+88ncZR6PdNqaM
DzK5YTrzdLTr0hIKg7MjCFUrLfDE6j+BymDDTVdV6Rjsa3bCmvt0Jq7BNhxG
Fovfr0M9Q3x7N5O6CwTwuv0DNFud3a8EeUF8GOGyfAcORnGjXv2ode5scsrO
q/l5vOsKVpTq+tm+K3VLrw//TGlfzI8da7LUvdYQwF/sKFO/Ja9yIs9B+Bsx
qacLuyze1Zdx2hZCxFPL5mXHrmA/TPqW6KnqX8MJyH1A9OspaO3ncUCw6PaL
KiRb+/sQcznc+opxqe9eE1f7KACRwoT6G8jFnULqj17VP+1xuAEsSfRXyAv5
FWBmkWyG1YuRtEvmVoCBQpMIjyHkSKmzyAdaKy/POyQfLfMkoLaUeIRiz+Bw
TomhRIX6brXJT/wkZwVYNQ5T2lwlz2mZ3w+w7ViBWZ9lTqO771f4gzNjFT0V
EzVr1DetOTu9nzK9jVuwxZBNXQ9Wwsvnt/TLSqvjbah8DjnmQ0fyaJgWMlLJ
IxehG8X5CYlip9pJdhkggqdKM3JGFa1ZoQ3SESvzXpfk4p6YemHYYEDTQtZv
Q0KIpYjBE2JMcWLvDALrJCrQUE5rIOMxfumrCkyrmbC4jzcN1BXkVXpfqoqC
jgERC357XxNJen3QmshkP8fY1cv0hu5Urc8LaL37FGj7H7V+0jYL3j5WSc8t
n9BtRXAiPnSQzb6GJWdE3oRZY4fecrv2SPcRN6rdAmfCGUQxDs2bgD81zKbu
GPGp80YSsyVvsUZk+TOzryOGHiLZcvs9uq2w9cD1YYtgJ2/yz6+Mb9V3JFJg
xqfRTbNDDj4RnsmNah8EfS2vGbskR4C/xIJhFNrn/38PBuQTkCp1mJh7IEWH
eKFsZv1pw1lFMV3x0eMLv9UCKb6RKZYirewzeLyk28+nAahTqDiM7tmChRZh
NrQ2HJVx1ILonSuzVtI91nqOrJpEdnP1VFMsgoaERmZk/LavKBF9OihVu/ZK
jSSlVAodC0mMwgjWJ2jX4tMzUfmjpfzcO/NNe4CWBoBwj0VzwfR4ZExvvjOs
CI7zdhNbYlJkCRME09WtWl+YV/lNTcL7CfS521BPY+nL8go2lN2NDf1rtq8Z
/iUZPZwsdd1ns7CoAN0S88Dzv9BxDjV6SQmn6vVpD9VuRbncNXnepe+Vc9K6
3jWjfT/LAfL8be95Xh6LJVfZU71TD3BL9Kf19PDml0cq2QMo7mvSLsdvJgx8
IscSR7HPOzmZjMdXgjylyS75BABNLB5laxCxpo+ck4X0DDRsHLG5R1BggIAM
nfGxh38jjCPgeOxfHDuWhcfa/V44RfxRzh+MeSVVJxvfAPO6DW3uDcXBGkkj
pmPQiz0vgl0UEkLe667qBwOAdC4zzyr9bvyPPjg/LYRS6jwP3uuibNipE4CQ
P3eAtqIpGtpV8lw4ALjykKm1EHf5olWp2h4r/BtlaOrfMCb7vhJSizlumCZP
mrV1LjeVmydHeZgitCoafLYEK9vxGQiR25Bd+lGw//+rkz5ipWdZy2/KWZh0
cnc/Wa+8ccucalnYOm6td/8m/Mr63BuFhRan0r9SRIHOboJOxyDGBylTsmpE
cRyCOW8bipTbhX6PeIULBA+CZ5pb0zBCFkM6egqJw90M0pu+UwExwNz52bLe
EZehjCgpucCGVMwLSEdUJYlWhYW659/mHcCe+LyhVYhpz9C+Otr81nEglie8
ZHWuJClyTwDqDy0rYLiSyEBFJ3R+zku+qcUxTtX248iPSyoAeCTSx8G99TZs
xqHyVLc/LyRAkSnvAUDOC2LegU+V58t82Dcd0u0pjqO+sn7lkv5pJsymXGRt
7p2J9HzTuyC10b0VH2oLjYmOO0qEMbSabCBRrMqevLmQ3fu67/julSSLqJHP
vW3JjkM81rx48Eo+3JGmTC445lOi5TCJpI1LHaluVLpzu4DSecrcIF1M2y/g
fWoSNDRFMMsfZzvH4vD2MchZcuj2rKOUYHIG4At6LkRdTa0TTQ7EuLTExcrW
HWIzZCr9v0Ke+BwPbgZ+0HAxUXstsEIuwPM3IZUAA9XlWEYSEAYrd+iSh/yW
yjVY1bh/lEH9J3rN1Bf9p8EsesGOO0iGL3R1Tm8enA0jwjJJXYd++BoBaDtO
TnUjzjtqzDbYjDHAMg0BX4wqzzr1MAtHQio+eMPugfGEmcGDAKLhg20GOQJN
e2Goca6/ucgoH1ZrBbrxXCTaMeEoncrhIIhXUr/F/6lq+PoXRJrXEDBeP6Gr
pZlg29PaESFzY0fRmJ0RxI5mPY9FWzNb9SO/i9ppYQ3Vg45T7BBnY2m9wIwY
ggaokjU+kfkeDbR6mhNK+4IMIAO38NA3tQJlLf0Jzy3SKthrMPzObPe5GzPS
3/NIqVFSBXVDo1+nOfFHfSuZpQfRsOlTPeYpN+NHBgQAGJchUy51lupi4xf+
FeQFjAGRo2J5xOfAB/aONxB2Vd6G12VWBhZaiS+6rS6/XS/vSw0F9wGU16kC
/q0TnC2iHFdh+bcnBvzxSFziLS4BFO0bj6hHHLyXxQbtcOsM2zaNgbBZcDs/
Mys3dAanfwf4N7G0InyyCgyyDwkg7nKDCYVtsKlzzX25YnJqLbm6et3SOMCu
E5MgJsTMuY2FMFAnjPP+jBYOdv6QTrHj8AlJSy8k3GnvDR/rtn9XS80rO7y/
wBQYJVUTdcCAd7HGZmz4cRrGoDC0j/QsLtefpVRlnFolZ8dnVaE4pDeNKw2M
G2cktz0NqtMtQXiwhX/XKgarl9rB6ZtZV2HNcfDn3vziHU6JV94/AW8JPTbd
O4zpCa5+cpQIF/Ke3Aq9gw8ikE4YlKcDELpC0J8LiSUiD7o+mRRX0ahL/R1q
aBTN7eTViUo0lzYZ4kX9tMbjqH+ORMl4EvailK4NeSHqP5uxugkyEdBSZIJd
kG8c1mV7uAlo8yXubUpeU2kyeW6Idubm0h2IFYegPSJn/f/F6a6yPZ0uE2jN
HHHADt/znz2K6E3d3PAnu1aOptNFci276jRz60wp1HQ2fWtu8Wrd0ZUYOlKt
amd1XrZ48SGQJtwQfnLqCLj/9ZZepwjbs12Zjr9nkW6/VsDS041y+K0OVL4m
DYP4UAg/0PQvNxgGODpV0xyHJsfdtqWO3gbBEI49yTje2kIk8yqB/2lNgJ1t
UzbuzmMB1PYaNJfXRjhXarG0pjNELSubmUIDUeXAqHT+cPTYRKAeGM308x59
mDvphAJjIknWLYcF/jEiqlg6OPjSo2+vCHUVvzsiFMIXOuaD3puh1Ihn3rtZ
jGJfrutaIYmPfEvsHYawelv12vBSpfK0kzozfrVu86Uucx2+rnccUKH7kgFH
qWOlYewI34+0SWcksLKXAB9Cw8cSsGpX5bd/gPbHmN5CHeQu0rRWN5rm/N0X
tjQnVq1sktc7CK/wjd2gNLHYBGFr8X9f1q/IxmvuIYBT1QhV94Z7rQ3jRH9J
ciXFVHeTxHspOS5aWhX5vO2NHN1n6HpgkRRxEwM84NujiP0HbdnRSWVtpq47
Q/RR8GAK99ANlI5ZeiBT2/9LFTn/3jSe5vryLUHasL/++bFF8d5oeZMufp4Y
1UxLuRT249rBJd9ftreAmhZesi9cNNULKoo2HPhozm2IqnPQFcd75FWdnP5U
U2Wy8+5K/Li3+sJKwsmsSAKsjG6LNyZThGrs6yHOEm36X/lmupA1VgnqFnDU
eE5HeEgNDdbWyWj1vVyvdVAj3ctPNylDVqWKGF1LSBVc3YttD9AVRAmTGkVA
Uy7hK7CvdUs+osYoGD/lK119t8UThANQoeP1/2bQ7A6jf8VhWu8kEF5PepeG
Df4dQ5zsPGG5ox0ilcq9jaxH/gggFAEimo/fQqPAmTFaWaZHRjr0rlSqgRWw
pu69tfULF34fi62BD6dh9V+9RUp6/ar1vNr54ycEQx4dm81ZxttZGXc2B1M1
2X95oE+Wo402b6ByWqEOCSEqccP8tSyREtZ5PfCe2hTKt8HNZLPOGQyKgd5k
MyIXEFZyNA7vA9Yt4LnwXswSuepLjjrsxoe9A4dh8kOkVutVtSCDdXZFvzrE
bMqqYuf5Omfu1GGZ3OuPb7CkF/hIXPwg1YZuAd9z9wo2JndrJ/O+tkulYe8O
CycP4Pw7xgDBswoFjjewjRBH1vZkEKL36V8k7mJe/88j065trrIjMdWpTZWZ
92ONPQFhcYw8WQM3v3AdsjGELpUor9K/fpx5Mdw69LAD5UwnaV2fZmAf0Z9e
+EP8+9ThzdZyBlfgYo2PYwaOM2Ctdrlu2nLLo6rByNUttaVlqi1mfayDyHuu
/Ayh6oYT5XH3nkkm1/sTfCa92nAGWekVIpOwVyQoM5qch32hIYozPU2L1WRu
QmGhiAwqcdIKfkGB6ZLa4w4PX7EP/z6f9EHuwQYhIQjlT7V1lrPKGKdfSB71
lYWkmqyCBfYTeOERzR7+irZfMbXkFXpVNEOQg2gsxAiAISV1LXL3RbWiPnzT
rxAAfmu9HjMukHxLLoQHR4m369NbnCpyHVNinWzwc6JnXk1/q1MR5r7f9I9S
wUMjFE/wJDeWA6hHIfQ/f6sPNA249itlhBULUrSH5l7KsR4ECKmp+Uh8xOSo
XQWSCVwKBYl6nhgRvU+sIlM/Q4RMW68wLfnGPQAvKObwR71HaRiKCDwaVBao
4lX/3U+hdi3scd+xMubW0KKbh8m5OCvUl0X+jBWZRPPp58yZNLArBcWTgzh3
x7yXLBEQvdTXEJiX7bDI1+yfWSbqZSdCKDLgq6+PniP9+4L9G6OrL3dU8Xcd
DLmy6ndfRB22pjf23yywZ0LQPR46rs5RD33mFRtTqAPTYMKsgaW+BrC9frxn
LUrCJNOEucQKCEGelURekjj3RMtwe4k5dXQsvbQLM6nTHWetiIQTmd3aOyNm
NSr3r/g1l2cGf4wfljHhz495w07Tb/FXdGTxxhYz6cRP+AeNrj9EbF4gCrAj
txUddXvT+LeqbG+eEaUesVvYwu7EWXszUvXRuiZAq3qALExDwvLuRm4TFIFi
miY0iyAPtw4kGDeuW3AFvtMYi0wjDxOAOq3dCgvPl3OLT5FyFwgLob3QBlxn
ftr9e+WJgs3pt0FB7R+0YeWdDNA18CApB2ezJ1hR/8KL5/w8sSOIIaDR36Yq
FQ+of3QlT4uKlrhiZDhIHpmR6x9AFXech14osu8iQYDKYwoBNJEWlPCNxUfW
eiPuYf0W1KAWULCGFCplij/F3ln9SvxWkxaQuVWEaZ6zC2ZDByFA0F5pV5Cv
Seh08dwGoeyhPU8yDD3l4xVR3sEgvJgIHI/HEhsXHBdiZo1GDf/YG7ukRO31
CIjS7+DZ01vfOB/NueQLufCzuurZ6rK4hNoEfX5EMpK+/+v59p9Io77kIIuN
aJZ9zRTV1j+K7HZPUB4f+4i/KCI57q/KpZxv65aeuZdFLQTtXOhW26ryKO8Y
PfY7YBBgIRNZx64Ou62V/7/g/nlN4OxCIOFcnARIAwsGo1CQcWI6J3z1kpr1
vhfaMe1mgh57zTbvM8yFvQAZP1c4aK99oUhOkRGSbBeJnDvuRGwXZkRNMlMl
0Nc4uJ9oC+mT65XBjW9mUNWoKoYDNgtwDs5F77xTHtd9rvnPw8x7aeqEMvs0
nYD3fpw5IulLQjG5JN87lHgq/i/Hud/ercVHt/ZLGZ//dq+NffDoRw/V1kcy
xjNe6b81tMuqkvxQZXi7jNlA9EdJ8hFQ8rgiOGm38ARo7LURlnrcR5avsaaz
a+M4Xg3CAYt58pjwCNXUYnckRe/xczxqZO62l3W2bCkkacGBtyRtsxXG/toh
VctHuYnFT0iGf7Gs3mw78Ul43Otnj283q4bxpDbKM/G68mRWns5ioWFwMjud
5tuzfem/ydG/1fGUe0TPiR5nmgIfgK9yrL3KR3XEGWzvI/lC8Ko2iOVsx/xs
d4JonVsge8gbkjuy9ll/x4fbJun32FoRuyFJPk08SizWPJ5i5683qeLwKWsr
Pth+SD/bqTOLhq4zWv6Twsr3z3WIMWLDeEtY/Vu65BbEbHG2tQsBvoqTOLi6
4t0KePUeGv0UfzDUKl27K6y+8HvZgt7+J5vOWEV/uH3dgCaLiVAUhvFQaL/g
qgN7ak53QL/QPf9bvkL7/qw0mTK0FofDMfn8fDYW8lRCKIhyCUStx1yXVawR
ffxVB3oIoC5x2WzWSDabhP+hDOIdVF8dnu+2v/M70KPMj+rlne1DGGEuaHFg
Enh5NMxnYFwHIbEKacykgcbEp4o+Gm/fanuhPrHDHkuuRzW8zU8+GiVPggLh
gcog7NgYXRnxt0BJXBd7MtP9kTH8FOmuGKIlXDN2M3NVPMtMokYh+5QCSP2k
H5EmTC3NGuV49StCcL7iKuzzG8JxoPYMAaRGZOAfBvpv9L8Q0iSxgCoWyE2f
D0OoT6v0sQ6LKqcnwYep5cimBBly/nTSGRQ7L2rEHeyGEoHtMN44mhwJlvDA
e6HjFs2ci5TVUMl0pm6XTX3YbTjAjW5uP//3rRCsGla9p6NVfpPC1Bbtt3ve
s4UBpW1JWMP8sctcRPYzlYpT72elMbEaHVGmU3Qev8Kya7O7tLOqkpf78K3T
WDuPFLheIn9ksz51PsnQhahW6gF0v2nbEY3Svj+a4hfnu4XokY8/aslin8px
f4dTvS/n6vepArkSNcbYl6EARFrJiKj3Gqf557uj1zHYTOUudGefwGBUS+3a
CUQbvsymgFoIkfNNGi3PVBmObiauTOphWeQoOIOD6xFqz43VeQ8thhtPGsRp
/HJShXzkS8ZpXWJMZkzrUL7ZXgPR/9/5DGiCmF9ZLZwclNw39Cw9Kna0ZeKt
fx+I05opLRe0ZY2C1YQIKm5AcztKQas15G/b2E13J3XXXAY4+Md/+xhxaMhx
5Ov5HKe37TrjlK7GjyX98JaIyyppDZCyHBYRUu02O21Z78oPy4Frb2UXmzQc
4yXNK7QxWwSHeiS192ka3z7MlBizHigiirWnreVWjbXAdreAzzo4gUjE94MZ
wR683pmleQ8HSVjwMYXfemlhKML8a4ScmgLBbipEc1WYRGHOzKn5yDex5NA3
6VUOcaj2uWiTJRjBM9NL7nPolOrebr6cH3s88n7pyDPD8+xXpKrf5a4eONkl
fBT+B9wlKpiYdnmIxX5/wESrw7BBuVZEIqiFRv70re4oJmNtFOwMoOx/3Btc
qU42L/DusywvYY6qGjNh525/+euPMbVtiZ96CuZ8u6BmMX9CX6zEblxQ5Wty
CVsYW4ALkbKN1Q7Cdrf2A8V4IiYzDd0nVbgWmu0BDrIt+vt3rU8ezwiSd/GE
OoOeNtdoH+FoxpRpK2wUct60Z376zv3kYwNIa4Rmtwyll5E+fuZQZV8jW8ad
wp2JMfEl/Td2/CbwohT/hLePXL4b1aoUHDNmP0GMizdR4nlm4nJRDlmQUSuk
lcQaRPkj+PwhQbHwOnPS6S2NrHE82Ej6lmWz03hxS2yq95uZlCKNkWPf4NJV
p8/nhNkrw0yDa579evbaUN4mQUkjgdeIdsTQmKVcX0uSm0y3sx3RvCex5vlK
bEutcdyNJbaOZupqOtVe8qyd3LipLvEpocnirgzaxHiIsDJ2sXdcUaGqfJjJ
vWwl0t4zLIc5IbroSGILtF5VQdIDbIgpalNUEPrN3yfsbRIvs6bDvE8tfEq1
DB0qE9rnx2fa2SXFq3I/IX6g+5RhuaLIzpGPM1xCVXpzUdDZrOicU+hDQpi0
02PXpnlsZgN/5thHsh1wj6gsObE0PMSv7wEL1BdINDX4UDciyoYVVuXBOnY4
v1QqSR1llXSkPruKkQqSdjITaS8KpJ4MzPCBWHW/Qyttyi2qGzZ+DlfcelKH
2my3mCAVb25ucbfOhvAC5g5ZhjKvklc7DF0VfJ8ohMYgLGx392ZYqhLv+lET
nxQ/j1a5okx3uQq4rDffLkFwQOfh+/PWNHQ+7IWsRO9O8eWFJZFSxEoHIGLX
CoB9PfPkNRRbxGEd99ubpGoRawUiml7briKChQUEh+G14IiM9Ts+b8C8cli8
nh4OlP2bep8emdZe942vD1fVi+hMMiOc2VHGWPDvKSxaiKWvGmmPjKcYs/vs
7DK1nn2UCjbLhgZ2rrPfad1wWRSyXLsDsKz99m5lIAnRE8GoFkQS6dEv1crw
BT/P5A8A7edbJNK6kNZOci23L9kEPeqsqDpdYGnY6OjbGSH4ARchtwirurs3
u/ZlJnFFgcDWAvIVsnEhINSETnwHx6rnVRmhJX+rBF/AtePooby3HKiak/k0
C9Y1jQ+GbwnNSRx6ZKoE0SjXe5Nma4nFBNNGw7/SdpF/BsurY1u7721n0YGT
KzvPdbaWqcYsoHk8xuEB91/VwXzYpHmYruwZKRAm8pxE3i5vbkH1QcKWZZg/
t1jdfv1W6THZm6pcCLZYn90QYeBqKepTB6xmSSJD5ad+T7farZ00CZ3LBr/J
n8KjFBMtjtxC7xyrTMUCS2IAY8urJ80QsnVxhn5Tb8EeRC1UJkAbI51jVB3P
CITJge20EoqSCmMSEPicuOFT1/wa1qKBqj+kViw63PTUU81S3IPmHtvKVXnE
T8Jpbb9fsgIzNnXbA+lRHs0wtbP3TH0Bxw06rH9rj5bwfWYG2cUi6dvpTsnp
llJvY3YDAdacUEY9QHq4ObJEWXgK1bha7DT0EcSuqTgtVt3EORh40sIPvhSl
/YhsTPHpwYY7wmbjqWKqCtLfHs/ouCegvw/x+qcXfddLNRaY9mcEuiMwX6be
tEEPWISomfLTOAX8y7a2BT60TgcD9AN0nC/J8v9EZA0ExPYhORIeeomHsWNA
RS9OUdM6c53yV/tCg4xXYfDS8K0BxFE0xfmQTqeQYFgqqkVaxVifeM5LOx1c
4q+FfdPLBhn2nnDafc7jZlIjLpKOWAm98N5vVFJkALkYjoRC28GZkPJykbWB
AgG8BPpZu3ovMsFI8hQ9+SgjGQqnthUWZyJQI7UkRIIQzyIVxaB5mWw80FWp
kIcNBbgslhvxD6XArdVAv9y8G4ss2djbYFOPAk1/b5shdP++14DSRU6Z41HL
ICS1SDKgAk3prkAlBmzns2o4ME54MUwDOrg4kpa5m4NvZE+kQt+JIJitOVSJ
pWxDMjGelxMN01WegKwkG9gBV+hX+5fYS4DXybGUpRIpZhaIpj5XhqfILx5h
G4jRZy3PlpyUVneBAkh1bicL3uWX76FBwz8mvF12oO1CRfZ+AzMpy7ljXZ+P
2gdRhQH7RZcZYJn01+xxIhVqgT72AnRedM8BpkwH7MV5Ya62zNTMOzPv5g1+
FeOpMLhraWOhdnDaojPBUQPDaFcFpI5hm9pDWwrexkVMfg0GRFqSiCkomyfq
/pRnu68my17Wse28lkwg5CLTOSNwY+g6JsX0vdfAxOw8kFurRD6LipK3sgSM
ZKlQl6J4ywyeVFiE7BOB8rLV2uq3J1Mw5ONfN486RKVZ5sLaZSnwD5h7DmUP
tXM0do7hgDsqUHztjhfWtnQElpDCoVX5rUiJaUdgA9kkep95bJS/swkMu3Vo
wIJAsnfNXPkKkTFOLx++kM/gnlAlkutu30Q5zglYvw0T7W76VLgHAvJWfGl4
51pAbo5jAdkmkO0Dj+2fIrva/S7NCzCMWIOb+AdwUblmuPY5vo43/W0AGGVU
SsorF+NkT6qhrBGdh2v9iFC+HN39njRjee89RGbZjBjAAF9XpFyRldnvwzWi
MdWi41f5HPfLJ0URGyINitIhbBaFYfnxDJ8k41aK142hD9TPFGCvvgIAFKmj
XkjfnifD/LHVgbPSYga8uLhP8rf8d8RSby1vNOVbtGxwZn4cdMf3IGwODFFL
v1TiZJKaft6m6LrtzmRLf4C3R2kb+6ylHtHXA7QLai5FD1UwKtutKq4w08x+
JDx4pRlORcCwmX84RqjkkkX3cSa7mu9s4yWm8r9hIENzaAiHPUs+dIk1QC+I
7GiddcpSKJljLuMRZ6O2gixunEmibMrV/u8mXA+JbQE5rUxAh3RlQAjcNrUG
ih8zOt0I9I9xuruClNyJ81Bu80cMgdJUmmSrnNGDoKyD7hEgisE1dXXNgb+M
9gkhLsPerB9qJ2mkqGk7BIeKvGA/36XJeP5aBDRZL3lue4UzxVLKquSxM7xF
ZOzTu7UXFeyjlX0T30v3Ho0UgJg8VTLAn4nc+2riwnXBeFz+Rn4S0/zF0uxF
iKZe4QveBaB+uFAUn+pcIGx8nrHZckwPWgpN1osD7YBgm9QZCb6HoOB243Tt
OTTgvH+h2vvQ86RY+oXbB1b7Yvlg1g831b4fRI7tQbQ5h7SSskLqC/oSqNIS
RkNu6YiAXD1KFtQSfuIx9hVtVfl6kG0jVcLt80LIQyWvrkyT+0Ip0lM1sKNM
iaIvrIq+X37Zz53Gb8SEpzS8+lgm9je48VvWGGAKdxTScrtSLa9o8I0YZxGC
yIylowZLZrtV7nvSfa439RBTSfz7ncrTypcoqYXIJnRGUu7pMyiOdX5Ea1bB
NTmqmO7au9FPlDGOY+gGoc2Zq6Vj2bDUUlTT+d+4JWdZVELIlWVjPFSH3H5X
Cg7fsJ5NBDG6cYC8eymehHuJhjCNSWTxADBw2lWn9ZFvAvT6hry6iz5o0DgN
2Q6GxWpEUjdYJMbRq6gjchXjWLCChA1I9bhOlGUwhxokxhE/Wf3Ur4xQFEAl
6e8ipXhfeITuC+TN7m2MVyqfMyZO3d8DOYcIsVvTUgB4BjgNcb7/Pm7EFZNs
lgXaMwOBu9I5dL2Sikryrv2HRkwoaHl2arqoCFwN3ttKnI6ZrDB108jxvFFf
KaRkR9Br6y+9rJEhpQZ9OPokOQrpuawLp8EsoPiqQUjXGZfMN43fwX0Jl4xm
3YSc3+PT+ee2gD5kjHSEcWHMnaGr+7J/WiLdnEUoJT/b1iMyPItbkgGSDGm4
tHUj1kHM0jfjvteIYp75rlIb+5iSEuCOk+OTPdw/ZAAvH+3vzi7vjf48GX6R
s1Ea6k/kJzREY/eM21yxNKY5VfQ8VtaYaVcrsXIyGrIiZimO27B3XgeaUafS
FLKw9wea+5lKbhjSx0F+OdhooOrCMenFOXHHe4hral1Qmy36T8UhnxtfFKyF
GvEsAp6/ew6fiC790oQ/LnyDBdjNAtUYCrJmuxhwkG3JCLiJ+L3kaNVWRO0j
Bjbqxby+b6rhpE+V7aZ9Ju7wmkGwBFwTCLbnwHoSfDt8bE6OxYFtzqrmf6+A
8B8EyBEqVO2uDJNwlytCRIfgHJm9NP4Cii986rF+RlRUR6fpr5eeUAGfT6XO
k5PdbNEVw3/AzXtu3TxLPPbSv2YpXSizf9crwBQbBEjNQrV8WO/cnETpE1oO
Eh2N9mfyTsjsTkSLNgZmuCrn0bNjIZ/lFtTzrU10YgDh7VJ0oSycZS7DE4Ds
gORNqGijzddFlIZUF1zhMdD3kkb47/EV9JgglVr+hYjX9zG7MrQ5EWuU5ZGu
K3bQO3IxhpC39zdLiwWIuYGoin671zrEXgaLjMF/mbblJYKVE9rmC+wFsZBn
nQ1V/2KzltL+bXWdb7AklpokkVmGMWjKH2geL90kvYftIj7zfHvQl53gWmbI
AzWATVDHcXRfJxDtJwXGKWmZuzv3+Tf/tJw1vD9ZkAEcZEGwmgpCE4SesSnV
oCryKTaHrndmr1FL2E23DbOBqFe1Z0BNt6AtO01my3etNGo/+szHrI0+jApC
rlIYzzurj/qkNq6+Z8bYEEo2APbjYIzLca/BnBO7wm5An1TCkEnCqPfHHTha
K6w6+5xT7TKVmVulygrXNwSfnefMqlrL5e5SFMZ+j+9DtT8v03n6zgYb2n6P
TBThmgG8lQzj0h9upS6C/TgXL06amLrKyUQMo5o35jRCic5PSRa8ObOyJ+Vl
a1ypEjlu3chIEaUMsj7SyDEfd/3JBpzbEi+DMmLhNBaCavEVDvdpAZ80Ycad
km+Dq8MG6vLr47dbqjf4XrjFoFNTJqC9HvjgTqjkhK/ud4TFhFvaqNInRLqb
1LTyNYNgptgRp45lkoaGrOmrVZYMJ3OjrfocoNhNa8TOSja4Uk8h7aiP4KSv
Wen1tMOPfTF1HYa0WLtcdSNvtNRQEEyYn+Wy39DiBkW9N7NXFaYaLe+Iv+yR
iSF2rBn/Z5904oXLuX0DNHqcO8/AytTNsSNRcK774z8Yg/K0iwIRb/f1SnDn
DPiiIp+x3nrJLrBMTjpJ6g4aZGmY/xBhs2NMTpodVOSQ8F7iO+i8wftvsWWL
3GUUS7WHyvZ3LobBoOQM9hiK3ydwH+Pf8BxaEgQUwgO/26hNSBqwxcXIAjyn
duEMOfIKXjHiXTUWc8hNNbxdF38IRVH5PZZM1EYQGu31Inlc3gbzKJKGLc0u
DFYWbna7SkGBWBfx8EO5eIw+DpOpBb/tM1Q6O3QtflcLYr4Dxgm5QGks1cOJ
6FKDR4q6hbH2RJm5n95MDmI7XvGgxwkHK5GJiEWrpSnIr8lW9yrGbfiveJqG
nCk2r/dO5cqTsTxQLjckLIUHQlelRMk8jb2/h/79I9hGmZqWrjwaTfM95MJZ
nNotCwbZcyz5Hspz5ddFi0OQGC9JhGllIbW6NtDEgWMyNHuUyR3Xr6QtVmVw
kUdccN9YFm1dg/ozxZBa3IbvO/uca2SWFllN9L+I3Mrm0VjraOvrCwl+h7Y+
kEiID1cSitdUQlhVRBkzdvB1M8YbkEKfTSs6DvITM5RVHAukTn8VCTGzmUsk
h6xI9fA4mvbycSY3rHBIyCjY7vBGEk9q+BcgFEuqRliQfJozN64H4KErvT8c
voMZ7+HJKeKfECsV1CmR14oyQpt9CiVedBG1KFaxmzYZU4393ZPJd4+jMoRI
9EHhC059mJ2uRA5tEhYVyRI0An4hps5H5narHzVDf+iszPNmih9pbmnxxz2y
fca/BeJtk9L5dmShHmFjX2VhcscXLc8rmsWpNuhiGW3n3DhI2xwt8JbU87Hy
JmIOBKEnQrzpZDM8P5KVu308nTcYskoF8df+DbARhn5PIcoseA3KSi+Hc5pw
xVa7MdgBibbY9pt07f0mg3KFrIfa+1EnceMvSmR2HLQTU5qDN9GftujKdq+t
E93wY8aIm5d/zTNvF8QrROCcWOdzEa/wZoNP6acM2lVO6wUfgJRWQC7EnBLi
Xqz1i2ZNR+mSlnuEd2nIX0NOa1SwYjhh7X99FhHJFJHQZ16bCoe4j7dC731R
UrBOrlX49sieTXKR522GcNOVnZ2MbYKW7LLdQ4UZmAfSQQWFd1fBpRHFdRFe
NtDmZ4gzyUMwM4FJz1xTOyqz3yqwnijB1LjDK5TVYQ55P4lVjkb8sGz+PCGZ
jTibflrvn4gb1PIeMLtoPVXbohIzHmoXYLJ3ol3n9q3+e79jQI364EW9XTZw
erWdZ46SGaoxcxFRlfziZH0EopHnGKck6SFB0sETDXaZITy8fIGEm7L4SLpB
hIidjal7W7aStx8CC4+jaYB2Z8DnHNrn8PZc7APHq+AfUt+kTty1QdAPogmx
h7GHYTCUdkjRlZxjfPYpWROnJmuulU1wjpbwLaNK4Ozxq/+f9GrFXVqiH/Yf
fwRs7aHN7N5IpifoeYiKSW5xDnd7hgFECawGBD2+0Gi6C+t5WW2/xibNzQHt
3VTPecEM0Y8LFCb47MVD6ez45ffjXHkNE4JGH2bnfYxSdQUMhPe3HjkTF1HZ
fTUloCWCn+WBADHsklGVg51IbdgaF6zgk82wVZzdYzl4ye0l1YZOHKTB5a91
ZuIl9R3nqFee878yDeDtG0ezph2viiKF+HlGaELgqgE2Bp9CeoNVB8lLPJAO
lnvaMfJfpANElaSkdjZ8LCiQ6F6a6Hwj5s3e5OndS4jUlYGTEkOdT7yiUM19
NR2Car9phPoFjNkeZDq8jJ6tqaimnmWqX9CC/2n0ILJxJYQUKw3pq34bEpdL
+AIKIFfJttjq0Sgbzp6+ZUQo+HLY9+92arcnxkMwTFQ/Bl+lYEtuT5ynAyoc
1glBSIfGtwspg1T1OBlbfspNiQKiQXMo28t7s2+3/FZskxUShBqN2qWpL3iz
kXlo3srnVvA+tFHuFE39ZlZV0DBZotChSSLFadGiTxpGVoiDPC6Ru7dIPIKU
4atjhB9rul7Vp5lHzeOW+Os97YDEGsOM+2mA8WgIR6JIJ8TAP2RrX3dOtSpA
KG/J93pRSZFY0cn6BSqvUCCtVrqm/IEKgBf8Y3/qTUTJ8bYPzfUr07wv/eVL
wyVFCdHCItfXyiDzCk+jC3sgjBB/XnqoegNTCDaCCvMBla5x30OrB9eZx3DT
AjDuqwN6ynBWkdGVW+x7dzKeSk8cG0v5eYl960YR8KtI3w8mXJf5N4y4bhUU
ykfMx7YML57vwkibuMGVUVD6hEyRmTPeyYHHfUslO85T+T6SPYG5waIC3Nhm
6dCe+BTS3nZz0K/SIXKD7UveOrValwWWeVp9L3Z/8FJAxIdWDPjUXzJlz7l2
4zSYaMBTF9EY8XXyGX8aZC8cAfZG8fuv8U0mt+BvVog//K2UrBBScgK0WUbx
zp0sbtDnNvL4eMKTo8Ep5FTpvUDo4pJjzQBtE9d3cpQZZlkTbGle8maB8ZbK
5plerxgXUViQ/3pn6XswCWXIVBr1E2Rex6qo01wLXv81EwIiw6En+ATodpPr
01+72WEDIzlURo9WDattXCnepdYyp/rNDpPubSau4G7bBcUervFohaIi5bvL
Dc6OGGjRkyF6Xk8qt4+saP/0NwttLif+te1AVLJK3Jpi90OfX5OEwUMS/LFj
WH2k/xWUiuZkzeMsOSVE7Frpy7bRRSDAJySqvIPpYg5RaOrGbmd3HczlCOI4
RcH0YpGqjyQIReIFiENXXkUfO+2ht0uzNDIqHXY/yepCNKsGmaF6pjhghZEb
0IrTOYghHJz6AepRawXCy4xagzeSGFH4KK8Zz/vGhZBJQvFb0KIvHduxskxS
0qW/p6tLGAReKo2vAdwEvDx0hXqcNjdr4ls0+KycsFWgXt1zsQF9aT8Jv8Fz
A6SoOXZYHCTT+vbOPMLuIc1/q3tK71g4IE1uEhU5stYG83gG7aRvTTxvdWlu
WgZsHKlLW7rWKKH6dike4Uxo1b38HX6ZTvNxBaV4SCfpMmUzyBZ9vO1ZE8/o
Z4Xqq3dFfi+Yc7mKAM0krhUbzfTyCylttq3kTAvX9OTc+eEGKz16AqAOk0DX
wvuJ+zsOZFZ+CHKWz4RA1/3qep5MIIR1u+aKuZCASE3Xxb3ZxenDxO5bt4FQ
iRqqjW6cj2Tib2zz8Mevp5krGIp2CXJNLqVVNeWdU6wTjtVWWI4wrrbIxNp2
TEmCZ+Y/7hev/kphXpehm5oKUjG9u65pIDOO2Y2R1KmCA8KZMB3UsIQZwU4w
aaEnIxvcawtB7ENHu80DIWCkNYFZ2HdHwLvCiagaC150cJ2JVasuZPpsPDOw
a1Jpq8eS+SSHDIBpjz5LMMXkI2hNIc1TD3r5AcKHk5hzcKJd7P9+lV/14flm
jmXW319gsDAOVcKAY3N/KxWbkGaAIjqry7Jfv8ZIyw/b775qD1y0SEZ8zSD1
Ng+wkofZUI/Q1GdszGpce7ZZhxORRSZBabfULEp8tKz6iKMeOpPJHNoT1vMn
ybZIIdGyYj1PFs48MtndZo632rN6oO+hCy7EIWA3bWnr8pNUTyZL5N4Eia8N
0IOS3pMT+f2fSxD/x2toY9yrZF3vQWRFR3CUKgkMUT2w6FxOCdqOcom1JBOB
L+0FkQmGOrFSSh5J8EgwDL+48Z9GU8hJ5VsEpZuMIN+4m0IjHQ0Yt/0t8DdG
kkd0i8jrtNruG6qVlP1flRV+FgdaYqST8TnyxVo0xPHb9R+qTE0gfmKC2pTO
+uQfx67wOhgIGk5O2qErjfldyZk5fJxPMHjSqxBc/FNZIkbkiXKgQU5g+Y1y
9v6AqoyQ25AbxQHlAebWWqLMynVfC8GcgfKdr5OY5aiOx52A8ZA4oqy+8gIO
pNZ5P3Sg7f3VCm7ehI/kJVsIWK7P0qGQQBYUzgb7XjjzMQGmOFF+je1/lqA3
ruSHKAYT6BxCI3uNaODVjKQz8uAGSrzDRV3yq5IeR2Zjdn/NRXnx3DeXJx1U
Jx6dpI4mBHGzyVT/nhoHxdQeiK5a9FZsONiPnO/1ruCxxgskL8bVDS/JHzzd
84Ab6Yb1Ce91jXMMRmO2/TFQjnDJ0pAGC102YAXfjB4JTfCyxpyIKohSuBLB
++blNK06Ce+/KnPFse0npkQdAFKzX3a8tsMTYOiNEdzUYOrlwn8CsDxkJOms
yHBJ/5In+CgzO6lX0KyNdGyiXsueEJ4XzhOkLn9nNUDvEyoKAZPYvJKpgOcM
hmknAg6Jer9tdeUce3aWzqSpBPOGgteLJ+fz58mNdEKQKPa6MzUtiZPlZtCi
BJw9VygNkhQAPDaj//RYJ6h6HYZgE4drHVoh2i8gqgziFpfxEpf39AFMcY0p
M2rGdRgzN4eD/SAKucqe5RxzqfhsOQewT7G+Js1AIc83aXLVjXYyIZid3a0a
Jq0+c31NOcKw5dgQwYdSFzHQPC+NOmgkIrxnr6ZA/RQO7n70L8AjMAc7TzY3
MFUAe5fxGG5KB64kQK7/D/Nq2u2wnMNNIhtAv9swer7QJR55Avvm6ep7a5gN
Dciw5N4cznk0ADHAgiAhtBOINwh5AzEZmyspGThIgHAMe8x5xg7pwE0DFXPZ
phtSPl97kfkcmbdixxYqSQCW0dNF+3aAf7qcztCZKq/G8iGhMpqaGHftMXWG
XSj5GUzOM/LiJzrINJUO6Mupz06GFOOmeqhw1NJBuU36fsQpPrY7Cc4wunbT
L7LISZoal4mcv+9BRO9q9uXbo2ZiKzyx2aN6VEZewlqJekQAuHiV0STJnSkr
G6Iqz8ZcC+Njh+EbisSmjkTL1oKcbsj4jRTtpD9qCcJ8GN+36wldOOxcr3EG
NThcEdpsVZBvW9obRFKozTT0Run40vgm1tTHiLvPpEORtOs8MJdQgJ6292Z8
uJn3A2d0Zie+Tw0sxZhgqygK3TeX1SiaRGZxq5kpEO2vHMAhK0+0nOqLRo4R
B/uC9vrVwWiWHtZRuNoh19UkNdBG+DqgGm6LrXM4U7xJ1Or8ppZYtb22M7I4
m6W5dEMGsHldOZIfb/U2Zj88hGOPj8MRnelpNUEpcmRoMM7LFyekH+dzGC9p
eZrneYMNsCJEes1frK4JGTppx1eqIWye8qvWmOHGT20NbR5QM57qmkQ9QTWo
UoARVftoO9RoWY0MOaBuAnmubiGmxQwrU9scV19nC4RGqkNwS+9yVhVUu1n4
QPnWcjDFoHzbOjO2K6Pt9wKRufTpEPPfjoWNArlIzeKOEsdhdf0VQsoHL8Rr
ldOoBnujUuGyRlggEBdUmBz9GtadciWdINrOBnI/HXzpIhWrA2Z8WuSy/2Bo
r01IVU4/ms9+fPlJfSl2a3lIt2FHdRe55hE2gXBweUcbqtvDKDrSp3f9qo00
fgSBQpkyb8jOdxN8Eq6upoAe9/hSW/dfoU55vgqQT7D8zUazGrL1BH9S8gl8
pfPWDBGPKo0sXRnbBvQF8k0coGr5aA3EYEARZgTMsVw5bYf7CnQf6kx4zHJD
W9LltAHRt/JxYx/mxTrbgXbjtSnQhbbqTDr0Hfi3H3LIWD4vdJ/GL2Quoedx
n8t+IQa2wuR2rYSysU/X+dNgfJDUKapdHAGImAskqGlrjxDZlsUVRZlfPNFG
Ot8Tpli92hligrYVZSS43INv3OOKJioJVVhElb11VWIRgexcSp0sWLk8olpu
rgQYuLIUQZ7Pw3BV73WZ0A+bpN2v2/RMTYZ+eZclQb7liQKmlprHKajjb89S
sIeJin0+4Z+Opftv4pppHbvWgHsuNyVMNLBI/5ZqtQtwNKbhGuu42xD7P/qU
oaBSaG7mioE22lHyhxM0HPgrFOlKVQcNbhEYoufdjOFOdVyoNqD1Mjj6kGhP
3kNgmHwkOHj+RJEFGfx4pUmIlrtMAUo0BiIJcrV7nrFrSKMgaTtKIBPUYnZM
j9adYfEQ3T0KP8QNtjevDMjFHGuHVmSisx2ci1+FXQJgLHrt0iZVbSMZb1lq
Kh7xm30Wca3BURRQk4i3cp37tuYM7npkgzhoQxfh7OFDXWB5SSQAJ7sqO4dp
OuZ58VfCug6W9yCgv/ThVEwwxZKL7yH/mzbl5KIFI2l+NQfcPoMzxbyhvkj5
Au8AdQ8vlyfATAj6BjCfc0nQGm1NbS2l0tZUNdhZKT9XB32/sZWQrj1VmGq/
caUXBDLxAdtUXaygA+oIJOI0j4/nRpmhl0hJ1fmvk/4NEmqO9O3cgNI/cucH
915ZvMuuYZpCEyMdAh8m2VbNNr8KjZjWvRqRwqDfT7LItHF0X22gFDuu9j9w
rpygU8Z0FxaqbtYa/mGwGBza0SsfUi3jX3PRhBoS0WlRGDk+tTbRZ8/2yJxx
v2/BjMNxfHFBR/8Pi/F4STW+c/BEgvoepCwYRCcC0ovtJtrta1M7L9plrEf4
O6/a0taWkatjErL6HRDD5bSPUTlaxTFO+w9OFYqVCQXrce/yPttddarI1Ag8
Omar0jz7sRyg/ad+LGvHvVUwjT2gley13zelEDONFNWzYw8TmXBdhBI04yaj
S4DB3obufkOMwpz6qizjK5t9C+toLruJSm9tOU5yG4CBssb3L4jRijlQVksh
JAm2/WxBxedRPI5xuoP7eBf1KXWhlhH7T+25/BInpsNope8Zv/AFKChaczHS
nFZ/3FcB6mOOb7EtqP9pBPUXODE+rx/Lu+v19/YdMQYWcvU6K+j6PN1qcZQs
cFMWbmuBnBC6+1GNgg1LGpHcf6/kkLvk4GvU/qzntjtBq4zvTaL7AGkxZV/t
4YKFh2Y4/nRIzE7vr+u6/utSi3oe+qyCtcX7L8rEPGzTI/+5jkavo4nkE/24
iP4H1ZpGn+GlAidVQqIFOirM27LdCnbOrtTqW0MQOvlIJf//dO5wdo7Ysxlm
2t4flkijGCVX0yVZeyT430RGG61xt6MLpLcW3QgUJWXFBjDD86ai+pzDfnIZ
bMqMmFAzw90DtpWqVAxL85I9E41R4W+X2BvYj+Z29G00upAQBTvPopbCktww
lMfRL8dub7xOOZjfHFU0c7g5lV6g1Pq2I4bfi3+RstfhGD4bmQmfmjYLMk3H
4uGY1SYhngTnwDJJHIXmAv2nyMXC1AAi9SSRSwpjJic/VNKUjqDmkxB6jhFW
yJfbF1zgNe9ud9hhAfm+WKg69s+zfe++fUZoW637TZp5ctneIfwvGTLMmhhd
AtIhCHVin88Sfh3Gp0ErcL2om4CAMynMamOIqfjFNWFtR49yUPi4msjj+Dib
UAHnX2jNDybx+UV2535iGlckzUDKbMPh4jtLNJ37ddi4/+N/O3amatjfF/8h
vUE4H7ikoEZAvXnwzipAY+23uqsaOwgtuT55KEpoaPD6JfZXv2RudxHXvZOx
uf6ojkJUxGLSsc6ghquMu5m/oNTFCHH3fIEGUUwNAutr0vk2+mJt3M6i4r5t
erOmnHDUCMZxDorGU/ptqhHeIiKFYLHTyHKaFtjU7Q75k/tUQ+PcCCScaarD
ud0LBPIpJwaJ0+mq3gpk2x3PyRpDC57PKIZbbzdsjroxyBERMISbPz/4aoFq
bE44CdrRNafmYbcPB6AzC4NGOqNn9U9E1/46quAq8XN+RTCxVRY8DhbcomyE
k+TbkGGOj0OvshvvDbyploT55OTdpk3LB21g0RP64+hP2dzApYRCzRYCzL2P
XQQnfNAdMytD71csZteABlRr3WfNvmU8tCbUjeb3c8xThsDGBmGm4dcfleZX
MeUsPo5SWu15zZtMal5uMKjr72Au4seNgbJRBp7tYvLmcmy3hI0rg3ovVjEk
UqVMHb/u8DCHzW6zEXUMruovYs0IKLUelB3t1XtmrixZAP8nchWgOoRuc1UD
wl6IH1HD4lIYnYObLC8zG8ZXZXPfJY3DltNIU+Jqt/FXbA1YWt5jUKDqU+dN
h8ken0vL6X6ztpJw1cFpTDqRwJAuYq+S/oTMVf8ojkBcHB/tIsf535O+7BWm
m6sjgF/J2HCMnWT58aP4YqdtQvsq8uzktX4ZR3fCaO51luIa/Im+usgO1e1N
mZwfnbkArP3Y0iStZDktrlvzu/YGwe+umGJ6xrrKHHClBRXSqufcfORa/x1h
00nDx2/p30WhLSyqlY2FjoyWlSnVbCuO/rQBWRjsCxtnjC5CyqMdxWiFNGoa
Swqa8FtRZMJxKE3K9wj46rDBKb0SkMAZVnJMIF1Flyy1Sl20GkVg1MS1lPhL
EBjGb6Eqbhs0eQSMIU2mYk6qQfVZUkfZvK6en+TkpTu5+2ehL/YPzPGaZpo4
FyNQwEvmuWzo17f9soRI1FPDj22fNK7aQC/8e8Y9H+EcVE8z9J4cp7xI4tUO
4oxo5ySu2CS56uIh0Uf+KBiqTJrnMUdqI3FJv+dbzt6Hlrso/POVgK+P84PJ
QbxjZj/FvxSNrkoPcMj64vVSIcdTQE4cMmW7szTCAvRwW0zQAfW+nxPIC8Hh
NZskX/OFEfZbWQuuV0GaDe5UG2FdDFrTC7ALJqZ/P5jIf9vgQei0wuBcGGgh
Cpv1kcRJoAe6wlfYj0fpVHktfJqHBhmfwAIZCv/mulX/9GjkQp4dDYAsNFzi
cPPAY8Gt4cUCSOGFaWdv3mYvxHMYmxbLL6kzxtgP9Q8USbmD5Lz9We+aGz8x
NTH/C+YZmfrIynRUYZst1orqtC13CKGb4MU315iOEa38SLAl2Pw5yfNNmEij
/W3cWmkxg3LiQzInBzIfwFumBJsr6qRgrMXQkY6Y1fgyvT2kXCscqj7Of3Kz
jU0cEa4kG1dju4VE0XEizZi9XCtt3fuLVPrZ4UG6Q81ljoNaiESRpzb/19WF
kuoEHQmGM2xczvxlNYbGkinr9wQpFAOEZZTtmATuLVh8L/hH6zaH/azPMf/b
nqFoLu1ZinVtT1XhRmYG4Ge499/UjTrCXC/1hNcRrAi9VSl8nGPeLvG9vLo6
9E7Y/RaETg+Fkbyrsna3/0y/53YTFSF9ourFGFlEUPwi9rCKZV60X3TW1sdW
7GE++x7IEp5WrQ37t3p3z7BbisoxROcia1a9yOOM4wgImpSsGdZ8zxDjrEF3
xlR4vQRvql4J3IHI/dIgQUSRh7RH4x6TWnYLNzlqtLBpHMjSd8Ahux8hcZFy
x1vCqTbAyNq8UYtgGGJMoYzUH+RfGQWX7MNTUzITE9m+FcMa5QOuOPwYkrcv
GXiCIWA1x1OJpI+8NQvqEQ/+fymprguZm27Yc65e7BljnE/a1AMTB03kttyG
5nA6T23TLP5y6d+MMNcTtOf2Q1JjTbsMTHsEMdJuC9NcnH+SQ7KWW6ds/8GY
AlfEN2TBpsMZ7NHvh/glwXYUjYol/xKdt7e72IofRVpXiRV5EKKMr6W35KFA
a+Onoraw1AuYztbDcW/KKpMScOhSViIQsKWegOjmg3BxbI3Ik8CRBEW4iCfO
/GVR2ByApXJAZ46tb5t9rvY7JBtpmEMZHl+qNFZwdQzAdBpM14lRkxACjHLi
CEN5sjcaXZ26AKch9BLHsveUaaZabry2m3qg47she2Cm4Nb2qqoVUjCOP9B1
zXRqRB4x2K/wumifasQEXPBh3/sVR/h5Fc8fRtgHNovjBKdinbP7Gn3f1r/i
CoxhAa96b//LEZS7hbhTPM4MEGFF6MSBdYA1lR0bDikFEpLBtC+3gY1bQvo5
mf36EhIW9J9qatzF+kOBUus8rkvY4SoU42XvRBtIG86kLD6qqNCiRPRwLJBQ
+tzhYqy9PC+CPl0hwVHiivompP2heOpOf7R/aaaiREhuiQkHUcAkEKyWLydf
SilEUOaamlU/0iX2yKArFZMpjaSlyn/9Web4dm3mTOzjf6u3G121Ihr5mI4t
8DekNZE3w6EeARSJVWUbeAz0FwMmDpyrdbMWcYvo97beSlt1Waa/pTH2BIOa
rzhaqOlKxlxEehVLWqyKQHtu3R1nIyos6Aa7Wv6y9tdIIp+cNt8JkUmSYqfq
NRCqM9ZqpSxKuHcolv3JLZ82IJ8KIccKshD/Jm7YgxvTUMY6CW+D4eq5Te1R
BCDWLSXikUHYh7j5SkEIUsaYfiydPC7j4G0cvIrX1hnchYnS+1tC5EtoKXKD
7CAUDiV3if8Dx3NDlR3dAjWhvP8gHzjXx8aVN5ukWcHFEdGYKgfKQvmiFNE6
Xs00EELdnHgAya04PMV1gtPZ4DQGibotIUMp1W0YE1KN1kz7vkV8yxUBAoHx
FX0KLSsPvzyBXZBi+RhlZgapXJLV1exUfjLjsVKZK5TcQKDXDNGtWoMX1zCb
28z3hU1z9Y81yeV9+TnRedfrYRn5B9NzmyUH7HN5CxD2ZwMzYMqjPrEfqOjX
fkvbeDDdR7yw3yBkTOs1cDXHsDZrZbA4TqfM3GQLfn+wuNOYAtz9jBIaT9ae
YkKqbs9ieNvUxor/7QPvR3t1ZpUCyUTxTNrZRCCxyTy5l7SofYxy8sNhszYm
I5UooPYxZvBQCVPmBMvw0bSTtT34AecxL9R+rbg13S3F2jRBzWRhqiYCKKws
mdOhfoCoTLPrBh7sC62WsZccftLk8tPxH/y9g5PHNPv1VLVXbKuK5h9nESyI
Q8hAhXC4YXrH9tbvNKybRVo8N6qJy3Bwyd1p18eJuryaRyV10Rzsp4JuGBTc
6Zmax0giwFyB2hjVaOOx7257ff1VlhKnCpgLvg2nb6tV5LqpmO3nWuZJtHl3
ZspvBSVjI57CoWWKKYWi4+8MMOVQFyMK8VSMEM+wLZe6OrzWyibjVj0MBo2x
BSjikBoHnFT/mZx55pYY6HqcSExJCdAwyfKqSD0i2GTgEnLeKw3hmBkcwErT
Q9PFJYw3xbvcsJqqjT6mZu2eYRcIvg/xvgWMdDnfFDyT9URb2YlMML4yTweq
QecetmGiOH7/am6CtavpCH5jHvLCjjm/K/BxhKnPfP0myrk/vH9Y0ohIp/E4
PXQEyozW7yD6Zp4lqNkqct9YOnjJNENLdH3bwRN7tyvbStMzYwyq9Lk5zIFE
i2jA9U7aLwcQtLZRTvQNpgEqHy6P6MiuYqOAqm7oWP3jzAvnqNtFR/Gqg94W
VKhhpjA/QisYxFovm7sOEc44KUq+sLScVmxDYo1j4JvamIGRy6rcfYN+hhIL
h26fdjjVck5vjiAK2XXwpWDNs2lh+BU07pZlqqG8lp/HM10zsSKQgQNOInFq
QHho1154xFPbM7X/NSizjRg+Ail+zjnAvj4H94Ci1YSpfoRi9RNlDiRn3srT
AVhikmkoiCzY3wXHLGvelwx0PM/M8YZyVp/UF/3AFJp+YtBTxSlKORnvj+EB
hWhWgRdbhMBdf9JYzqIfU400c7iF9lU+mI4m1tfwoZeQHUD27yK9HniKotul
LJGl/PUteJVeL44F4/KogFIIS/ZPi4dpWJDrsCChdZNu8oQ4vmSLFPVryzkq
IOkAIT6DFHxGU51akMkeK1qaFnwbpVCHgeKgaQGLLP/KamOCPGU6EBtBzqgI
yz2cvpC9/ZrcCc8LjHrgUCgzea5e5I9UFOrynxHwDZPU+U6/m0xSqveMXYmQ
7+9sKtICFg8yJjz6T+pSGKNynDc2TpoO0ALyM9d7DBck/iT7l4qxX12h3CME
83rEnG+Jr8hjnekzrs1yqnz7xdyXQLHbxibiE4tyEhPRboirjjR+NZE4t1Jf
sL9qafdhjkuy9xTZm19GoKjwve/kqw1uKx/uB+b7LBChRobid3ac9uSm4KlI
wMcEvd0UOlqQKR/P3tvk5Gxz4EVsX8ynEp9SBpBmtor6PFkN5wBF5gBbSqoB
+z+Y2uvwfKPwlkgpIrR2beTHM4YeE8byew7gYueydVZb3g/BYVQR1lkfKay7
CJnUBf+P1OwxKtPHGI12Yd61ZO3ELqSRaDL1620MV9MmjAH4GWbkQbbcjI9k
AoHqy/gdylJJKE6nuPhCaNoWKrwuYFSUJtBG1OeETEfHwe1ah9+nYbsfzHYm
ChF4t3jpYsZIu36teikieoCPNrG+s55PBqyW7MQXyLmtfOnmOgiLBtbWSDML
ZKMrjCQVCEZ4gRGNIhOVhXEuwR+ZB+EGMAZv4hIcg699UaEaMDtm/+CAdghd
4F/c2/4XB/pJGrhBDXSh92mT7q1sCXswOwzVC4QJZ51oZiqytWXknXXJ24vm
6xippPDy0gv0pP8UlSfLa49jT0+NKCqrPBazImtPDPFwGTNmoDm/tKoqUiF2
ULPJOBkSmxoDwgcdWfzLbXRENVoWmWY25TPeI8+K1AFQAB3w0PAX/4nPGXgT
4tE4oNavkFPG3rfSJctFNONMdON5gIk3lg92O3sp4kngJAm0/9/jvMNOPtZD
u4BprmdvUtbTwCt+j/8bG1eLFrsfbqfShTRAx7gJFFUM6wGaAItheDouBW5s
U1P1F73o7xzZuuEZmnLFAlgxdhuTIFEf0YY/anX4/jmZQzkN2pj2K4W4qX5w
9tZC7ZzxP7IiHoq4pbQwgsLRjtVk0IIMxCVIlSqSvQLy41tgRVc043GWPewT
GSwrRj49IKOSYa5/xXHYPY6ytihWCle8oOhaKVCgnKFzQ8T6Pq5ety2ogJh8
k6WvY7zJcuOaTUFmsuWfiQWYdK6LKmy/wCNSmw64vKtAqmgB7si5hqX9xD7N
PAT5NnTIeII80Z5jwlLx1oAFYiRoeLg4+oUKDR4OqT3ArBVKggQIdGDTCkL9
Q0UOyb62KrYfDyGcQQgU69dy0N90jC9wbAe2+b1eNXvt0EAml8IhcWZezNMr
LPaeDe2+kResXeT3K1xpsXvN5T2Zp1c6M4K4DQs3ZHlNho5IKzUpZnENrS2Y
ZKK+qOopJj8GU3Iq6oMXxSgjmmH9KHH+pnA48idPrdJtl1Spxme3M2CNkQ7l
lTOH4gGzH4FqsBZIgDZUbwG+BnM2M8XXtkf+LAxdPbWGol2hwnEtOoUJO5QY
Swe5S4Kday8F/v+Hpest94jw+1GExuyNY7siPnlA6+LcH6Z13DiKOboKKPrc
sw9v/iwtazwF4KOV/Yi6olf6PkTTrqsDrPLtnCBmBdU2ioUkI/hZbo2Wbg/d
lDDK98Bk5B4lJ1KXXUhufwJIyBAODml7nAF7BFPcWQwh6qKXRTFJQMT1grSv
nf92ulo1WlSSXbVNUeKhlx5qZQ0/d7BRx7QAzVbtvF8/uDS0RUwNhjbHxn59
InLV/6OgkCQ0vm4m1qtpbCUKW3iKzxh3C6zc/etYyawtyMNDn+PB/CNRTxGi
I/gRKrzB30sbKj6yiSlc7ykS/iFZhe8uVPNoKVZBSKfw1Bu8wKGmaydUC6l6
cyoo1G1nwhNH513a+tOMyLBo1GVAlbBEv/H3YjXMZsROjAxnlBKdqh66UljW
1l4x28Jz8D7A9VQvofhXWnVX4ciuP0OUkSv5xSL74AUMqtf4np3f9+UzSL8s
dHbMv4GI0xQYWzoFdssIXU3UWb2y/XvFNhFcYChQiWZKHkXWhDnEJo/C6kmR
bxXE3hNECjpFA4OZuMQp4xWq5vdaM/+9DyqTyW/z0yzQiM820DlcN6CcG124
CzVM1Xwrcf0NY4grQqgNS1gJjDt2wcUI1GYSwksbS+3tmh+WiOR0GpeAu9uc
Kum2nsrwbI+RQ6+/U44eUIkMW6LiJG9oAR0q3jlbxwWPgFnkdTAGgRqcWKZK
yDeH7PiEYaRcGg8dnTYVJzBa52VdDSHU2ysGLINeKeOj92pRTjcK4mLq4NQI
i1SY6Q/2OuMrSWMXhR6Q3qzhOec0BFrwW+NVwALHDob+sReewfHxne+YJut7
4aFJAom32CUhAxnQHqaFuHJzF/kBuGajgHAJTYx4X/GRdhrrCBosbpEvYfMN
qw+m70bI2wc3XK3K8lqQj/qxZ9NOkTAJmazLaOQhQCASIPfP18LkvK4IB4d4
zH8UqzhXfDd8h/4VAIyuTKECS8fcbRksS7K9NuCCv7aCysUcTHZRfVv/3fMW
4dkZuvKidRQft+aOSdHKGkQI5Q6H8llYRuboR3OZhPZtBb8SawzYoNO5nxAN
qM/1jQZQmie4n+HyjdFZipcuuL3XJlow4djAII/VhsnAXI18ewKEJ+HobKa5
6D0mQQAA3voaLVbTn8kgkDh5bgT8PGGsqlL6Ipup9y4NBSmAJVF/9Ykif0U2
HSk8uX1ds5w5RAA5FbpdRicrn1TNRdZ5CPeMaXi1+x5lqOmvBSHmioobkFve
JZziysi+1jU0gwI9GhY3Ws1geUtAGAatF9mLB9dyw1IevufvmiBB5pV43Uzr
ahgzAvrjSthgss+R7nmHGF5zEFfSTbXR9hI63xqJ37MD7ZuhEtXKXNjAyDj6
TjnteyBeVXHlk2itgXUn/wg85DIChI0U54PdqSL8iLhzJVQwttDxJ8ME+V8D
nC9zrICBSzmLz6r8RI/bMgWp00H0PCiOWRr0Ps2HEGgmLx2BvWFUYABsAwbp
LcyRsIc4YuFN0WkzIejo7PySimXTr2GvlNgCHUUA6uz1Bd9PzAEOPcEWD6l2
935aDbtH2e1siTZx2QOBZZ7aBSr3w2Tx+CZwX7gaizXVn4RjB4fkTWPiRCPC
GJB6s12TbLqCPKAw6vviYx1RtcT+7dVAJQhhYCnR/+CwqFjlh3gogL8F4yLu
CmSRGYovv4orD9wfMuBC5C/qwIcZuUDwhcymczhSjfFAYr6HOnX8z1MX6wou
zcyJsn8V7YvFWpSrTp5pWS2tWkdSaGKBX6U3RlZASEWOId0SxeIYfXhk89v6
Z0WH5gUpHhpQ9AjAGBgIY8w4w6cyEa0WhvkyQI/+3ONPsTStaffebcZCP0kZ
JlCgDbSqnVyDKLyfH8EuZwc6m52KBgAOVcqpwRESuSC6C2cTSHuz+I+N6RWO
Y0Xd0CS6fDMV0XfbDVGIF5VJ6Pr9CW67Mzn4SAgC5ZIB60yhh6pvIb+nNJn6
LSYWaFcTnc7bYNUcvFNzYOHoWDEeYM4CwCIwC0gicE57yMdxzDviA4N8agGt
yTihI5/dONObKg7JF4+RX20ny5TZTtges5YbJVPXV8zpGfZCTuI5xIcZnpTV
r+rKCRo6n3qPj52nkj9CSVoAXK7NGtKt8h/OLKVbI2gFuMa+8e3MbqJl9H2/
HhSx1kLHDAlYYwiliX0CRFHCb4ul1vAZHxzIvV0vqYLRaRWayKHaoJioIyYt
kcCqOnu/4XM81hFsxWSiQ+WcJe3Qm6OmIIieF1+khSCli3wJ/0JNWdivMRGS
I6bSR8CRSVyROdF+TgtF9lTHyLGKzPyAGfEnibHfFGEZUitCEm7RZZ4QX9ON
bYH+ik3+jXbUAIWQNHckSqcYCUtHfxKXr/JpzUcfneIc9xc9RMK5M8xArewh
mfP+BYPqahEHZN7IyptdILDP0C7s5gQtkY7001C2boNdAiO9ngY2Pd5Ub/k4
r5bUTcogRe9AC0VfVp9CsfgCnMb1/XnrFQGmb5BRH5drj1gmqUba4H1lHeSA
Y3A8jlcd43m2xEYHcfc3B5Xi+ZPNB40zvi3O0fpaPws3hMyVsEDUEwZsgVed
rFkPrDrnCJwXAHlKBdB0Cxfq2SDqzdF6b+GYxu+XBe3d9BC1UJqA9wx8gSAx
g3eRqDigJB41SQvNyoTWfK8jkxA8c7Jkd2E3OA/SqA8DAds1KWQ+LAjqM0FR
RdU0ZubyMsTnKkUq4F2TvXh87sgnJtP2EA3s3tmm5SVCntOjM4RF2YCfa5a7
1MvKGlQCul3/6azKw1TuAXTItvBct8Nzka1BKQR2rSt0aCvNWfjrUKe/ZVdr
nVVrgaM0MbRsU7r8JmgJx76E82jdopa259h+g+qijCw3QS8d8SKEJh2JFI/Q
zlE6rH8BWkwYD9peKsCc9+gsQ11rfLaSDg50QN/Yg7/RxB+NeRywoQh2o0md
UDCU3qE+ZQj3HUkFg5GhaPVZkeA38AhAGImnVtVZe2nuQtN7oqMCQWK/Uo88
E/xeoqAix3AsExytc5bZhXs/lqsnW7b+lhya8ZYxPi9zfjdAzhFB7Izw5W89
67Z1fivESApvTWsxNDPuELZiSiV5nT1zVdbYmPeVnIcMV1zrgrMv6JlTWAz2
xw5Y+5cRR7AIT/DkCe044uDR8XkPNliUQrLYlJGXj/P7ZqIpd2pAzk0IPhiD
BATUOjSCEorRT5d5Mx1hXyInRrZPksr/fciDTEIixMBDnvPiDD1rpCbbIa46
Kmn/KCeO5yrVHZ8B7/M7MJ7LKn0GcfS+zv/wuu7Tmm0OES+tWRpf6z3CLz9p
2mFvuQVvMA/LE7IzW9eLrj/AOHp6ser3TrFNPnHAGFVFPK38bfj6h/wYeKgp
RjCRXm4DPt8inGD+NpaeesX+UJfwnTa2WPDUauvBTO8HS3fih1QKnYklAtiR
BsMV+/y1SLTSPdekEo6xroemtKpsIKEaAScbmYqhvcJpJ1C5pM5iSonejKuJ
76ibMqjGMVIEEYlunkbPheKsirKaJ9rGH2mGz8f8yp3DxuB1uZC+bQ5JB3cS
7TVysTFB2Jy0J01YrkFozUEJJujI8k9wboqqBWfCdxMwaWRtUykUF4jX3uj9
1fYMpkwQHozldFJzH+OWNGZ07wWjnBcngbOpWS9o9hcVtv/ZkZZiOoQxXMsT
77VZse88mhrh+uB84wwUF5BfQAPU1sfCdxx9k4aBC6v3fzXP/cUrb4PVOV07
U9+J2qiQ1vVdw7J5jpnl4Q0Xa2LJusDGJlh7o2ec68eMdIlds7s+r55qux88
zJhZsPw/SB5KM5RbY7Wnpn/MtQQWkTUy9wtiRusEFoMsuNV4JqqtayChMhSg
cSoSO4HrIrW0urUkkzR5dVtaHtMaXcMLo8eefCIAFf2fC0VW8c64jOqUZO55
6K2uPHIwsN4j2sCRjzWOvRxbYu/oNyg6Vi5T5p0FSiZ65+BW5nL5bdA92p6x
8DZvMpLsu4HCKTAbCZl9MVo2iBiRScQNzacR5DjKS1uyibKTgLfdI6BjG1V8
dyc9dViCZwyalob+ZZjrFLrIb7eGodpTkBFoyP1M7qmAGIqYgxszbYCrWKP2
FtxORGWq3oQmaB/4odqkDnSxBYX54XlI14Cn0RWdjpZw6qoRnKPIoLtcRtBS
3sxnfPlj4PObW5zwCefdETqAAnMnJ17lDkEdXNs8rKfA13422xAMorHOuHgi
sDnUf4V2BDcPVdCoUvx7EIDhabx7MSNcL3RpTrKqc0u1pMXJgQ7s9PgQsStZ
5LflfCReekkzGN7ncSJ4zMbnrXllgn434nCotXSdecpQwNkI18NDDu4YJUHD
1Jwsah5/DVWquWirrJKu8rgZ0JyBmvb7q0UntqCQt3i8GD1GxHsMLMF5IGI2
P+AnR1Qvk55rIQe6ZX0kjJL2XY6mgmoH4l32qfniGk7GCAbb3tBdSigprA0c
aAN6Qo2zDK7XWAFZkm0zfPQ3rvrnrWbljLQQkyJpimB6LddKkvbBl5GOswch
HtWCsS0xreqDHyiJETnUwdqUBH8iEZCZ3c42W26J7S3OcwXIEIe2AM0vEgnA
6UgT3wsg/rtHJGAqColPPYsR3sW/KIQgBcfCN+Z+ImRooZdfDjbVcjNb5Nok
3lIYjwPd1ntEtscL/7gGJUnsMukU/RR7FC7buwgtGs8qDAf06+ib5Erqpi6k
TRGBIuqiWXr8HbmmY7hY+cmew9B8PYP2+5R52kPsE5DTevoUza4TddO9tcGu
cRMhDcPvS5HqoYltP6rH2/4uZFuQnIlgfvttSnmSQwyh3vMi/euSPwS8kYBq
+coi1BrmH7KUEfVRiJc7yR+LOp+cE3tZFAEl/mh9AUzLPmL593wjJO3v88JX
Z/XuHF9cM0MlBJfgwxYGG/fJLK0K0WjcxRMc1qRYA/U6NggWsZAxWgRnv1FC
m63S6rVt493l1LHX0I2yxLvlqa09n1U0EC9zJIMVj05U4lw81BEyJX8aSkJ6
6F5VUWGcRILHFRF+R7XCYUUbmIriBePZ7llwW/m/1RIM7TBTnFftt5JOM+Af
PShJrrTgwQpR7LYgjbhPVBtRVsm6SWCpfT0vj+hgZ0fyhYD4iLbtY1k3l6I9
qNGxXvO3u92Id4yFxLxFc4osu9gxyn/gyLicQYulewFF5u224MmWGnd6rKeW
htyL0tupL3K22pgkgj2WBCTPq0mzWpFhG1dwOKQLiHIk+H6Bi90gZkjLPbdF
oMe2JPhw0VUgSKDna+6xIMqa0kpED/aUgov3kuLzYAliomzwnMmN0KSiMIPr
iy6z5ZsOTznz7FyXXpM6XgAcV4zze7sWSZPluN4YOfs9Jxg4DHs0o+WeGLjh
q/UvvsfyUy4IcLA7mHf2yookUZLLbTplg52QX+cXjqJhNhigDzCmj0Ie+xpy
iaPS/+Ak537r3DsuSZgTlGh8mHAXp8kcgSNjenHQC5VsoXqkWjPCKewzjSIX
tTaloiPDkPBizdeMpuaLjp7vJe+fM56X7MP4b5YMDDvgI/nopblgzFviIrAc
K/945DlVZSWRY/o46lZU8oBJQnXDnC8N40R1gVJUQqWbOiMkORVKarIuQtu6
HTI59ISGS36oLXgqmwatxoLHYi4tLRZT6Ah8eTL3LEb85H39+xMYJv73PEIu
KMwSIHu6BGalHKwomYX94ymnnOwf8T88T9VrFf7YDoX0zSt7jGE/OdmcBitb
+2JBqn5iMtwCydirKFi4oUr5PzYo7+tCFnoElUNAHwbfIt6+981HE7LDeuoE
Crrrx//TnjfAFvBE6vt9q3iccDtIewG6RhlBNJS7LKIUFKxMveyT+BAVHwdi
OwyqD9qYxtmUMyq4RGwk2glrAOSR1mxBfMEMo3ndG42OMg5sF77yq6wBjb7o
yXOeOPzLGpQHpxMCq18lhzKTUTITXFTXWcAq+eSgV0JW7PBNweR3DI603aNk
xiZymhxVeyX89EQ/MsFovjSnF6S7TWeqlR8N675G3xgoMRENYcrDWg+nwRXh
sRSkAA/4w4gcNlJYHgtxMMnuvbjctPdHZBxqfKqCjVlBvltOVKArlohAfA/Y
RG4O5SgfWx2gB6VQ7+4WlJlePW7nItUhpvc95MTm3R9BZmcE+TMGXUktSsL9
1/AOMMhLzHi4YEjLINU/lpp/BDowhjPNBSEBBPj2mLEYEP7UdV7ykQ7hG8Je
X1EA5EO/3XwsuQg+lkJS9Erg5rloYnlWnQbRtzWOxMzJGtX/+o4fsvFMJxq0
P598m/ZLC/9KBFT5VmcQGELQhd7A83NeJNB574XsVyh6aqm+KNxfLCzzjRbA
00wO53mbw4thuvzrYLVOd7dsLE6wyGKabVFpKRcyquxQQA8BJzXT5oHXkxNr
AykIwvg2KzEsfPamuBi3rGYnPau55HVbELs1f5Pv/WhKehlfhbnd03U53RvN
HQ9EIvHW5gqE7VzhMYHPPTjvXg6Bhjj29WJ8IqpX01oImBgU+KkUS41pu77B
PT6UwacpI4+eqXxY2U1hU3hJjPDqizgUhg46IrErohWuPNzf1Uc3+YW8rcRf
sNbwG5zKWaA0CaF9Pi3BjCpQWEQcVVkvNJSn/cik3LDbW6Km6JZD6pCI9GtX
d2nlzrL+jqi9VZUjyeEQZ2I3phwUZubAXsCwx+wcT2rPk1c9Cpt61IZAY2K7
OMDejds8V1cAUEna+CRgAciHorajqQjC7HzafDyZiY0eYFza6CG2t7f72lIl
ubqtsbb4TLK4+AgsRUHwEOZE7N4UPcBS2w0/z8Q4/gaCvHswY5N4HjhK86Nc
UIkqqZEjC9emD7r7RFvtk/7aErqmdOohCaO/eE4TCGz8LtMmxo6XWYvYbTjv
Sm6zEmAQXPdqjxAWGPnaCVMZ6Qg/hNFP+BwBKUXOhCJuwEWV5iEd8zMSE7OL
Igyr+h8foL3xQRz7RJd/4Deiu9q4YvlyWpZNUs/7FQ5zWayh0l8txvjfp5gy
XcBnYAKHWf14wVHOCv5h9gQypucsfPYvmTTGBTX+/p8UesEH7zXfyVDddGDw
0mYsLPzxGKi5G5skWji1F8BVh3v5ZqGKO9lqZY9C6E4kDycNMu+rPACxJpJ/
lfZ4bYQHX4a1HFRN+M3VAfcoEPyegYJNJpfJRRRk42+gUbPqW0kSZvv9/+5j
etOl02PGjNMKQvAiX25qFegKhZSow14g9q45r3QyAMNBQIgL/rkDxeLRWuKY
agEV62ygojqi6N3aefwthg9Xoo028tHiqz5OZ+wjadGt6zmgtdJGPVC8+Zp1
TS+2myqxcn2C8wGvnp1nCRpJ9qY+Opo0eJRx1uMggYo/EWSbnhlgFe0jX2GJ
SgsqP3Sdz1GSdVqPJAyJOLV1tm+YZEmQQ/XSOE7rETCNY3ISzRNPhul7VPkP
J6wthxwcC8HbysYSXSxnyVuEW02QLJkAiYi35j3B1Lsvet9SpXc93DdWJ3b5
cqsmlzvfeH7ZflLBtEkGmIhabFJms0mGwmA/fgv5s/Mblh9UaGmPO8Bts0F0
kVRYHF0vkg4Z+JsJRIaAWScmfWUdUAZO45diI44Xf9iLrsxd+Yk0yKRZ61hK
HCj+2Ho3E1DiyDjncq13X7MF+UAtt9HzM2t04TBdCNFhrGiTRM9HnRTD14X6
0YZaf+zmM8ohlsueBJELJXHOSZOLs2/ZqWqop7htFsbsH8T8/RubWrNG4wjQ
Je7BY/dh+y8u0i/vHeYUi/M5kmJdqP+Ewd805jJ0cFMxEJw3P5DPLAHqoLUi
vOJpwVyczJegF9Ov+I39ujxE/akilTkfODEjkSbGO/eQxFcEIwVZgf9V89++
lHvRQOYEyk9dhIIFEBVjZpIm2sMg2F5ER02xnK6jN2qZaF208roNOfFVN/YT
GEXf1i1331XPww62wGok1Y1WEU7cz4FMAu8noKOPQRXrJOFS0dyL5xPM/nH6
RlxupNM2tCCC2sXMaYC7G5ONb1/S6EG2Vp/2hRYfYm4Zv048KnBDFm6v3Ue8
zXyAH+6yf48hZgPl3OmZYXbX4uMdoMIk2Cr1lV6cOU2Ee5BqmhtOIR0SPlKJ
7ZlVAaT7wJAtCoxwin/WPgXIGznr3wVqo0ZiuD0FoAa/y7buLwgnaMFqNsOA
F7YP5UemhQACO3gTm1nhYVc30BxxlDDQEZ5ILzKn33AVbdrWHIaatHNUvYf4
bfeCx5x5xxnxwfLM71vZo58IXF2wGh3CR1bsLsLGpejQbJLCFWd9hRtMtOZX
JRQ+wDey/FGY9GI05JKmYPZL3ECv0LcIVqChDRNMhJSAZhZwkqKz5E9XMLIc
3k61UTbRbn6DQxc0Gz5GPGAcuNfEqxC7RasrrY371OWtK590jhV8afNtVAh9
akd8AOc/V0QiaXRK8zlIiecaluKzDxU2X2TM4HsMDfOtfDJlBxJGeJt/r34g
NjZVEySWs/5JRSLpUhwMLOOX1hpP0/uLqMjYAJRwRuGlS9mmWOCSJzzZ6GJ3
gFDuSSc4yVyxMDu9VpcoKkErNw1bWQLOKs2NDREA61YLwjj+FLvJO6V1Xsxl
CpGd68HSNTntfG78X+aFzfC/ZTPEw7eJOQrkHwfaUETvqz6R5XVCwvkSQyip
p59EKpJsc89wDsL3qyLFL8NDE2MzTQ4LN+nUSvPuvBgJPcSIOtdp+yhA2Pir
C9w6CMVq+tKMe1K42s1T8xqhSN0VK2h2fnOAL8a0gV3UHFQmi8bH3wmY93wk
63c427UP6YNXbxn43RiVHWHNlQXWew7fNQQh7I1Lgww0QucfKeXEshXBlp2A
YnF5FwV7uL5IW2vc+WgOPqnh+HQduQWaGrWNjSUrxRJD2U70GUaAaAMEXUIG
bot70AqEbOPiF3mzHJR2hwpxHdDNsjG7udwLpZNKaq277th+mfpb/wS8Sdwn
U4uvSllAXKD3h2odkDTApUdnXsPuIJk7mhVe2XysOk4DhbcAEPwiPny6xPXk
SWVu3+/aUpES6g0WCGIaQvJs6IgssZuHPHLHxmF5RCtfx++hJG0T3N/hg/AV
6Mv6C2xn1G9UsikBHqOpNpkl0DocUpz0mlS+13whuBjipJngrPXPMik9CgR9
gbGcHVtAfdbh6T0MdGbpIvVKk+5IlqWZrd3JatV2WSw0gjYlSfOybBcE7RJx
VYP2pPKqFoA0gG2pBrk3ZZZBxWKcukJ5HBZh6Z5l/u2dgrxUuHQzHcMCBjJa
aM7ZilMe2eTwxJn6FryqGE0pq+rOJu4O5qBLKjrg6XgFjco7VSKF8CcK7EhH
SA4jKUuas0RJG5l3u8asAXDMYRrnk1P68XxA1Mj8+vN7iV3Ef70XpDmB217Z
VQIxTvnruwYdfgJGSY4cTnMCYBCv4Yl8McoVI9cMTn3gYhULt9UVBRR95Kin
bysNvS2ZYRXPCoBzoqGWR9zjMEyKqbWCWE6W6GFQfZceoXI6okrtIiuZd0Hl
iX6JzHk7m8vDZawsFDwLfk4Lsk5WNlPJLzb6/nska+Zjdi3zpDqLp3F+x+Xi
qvin2Oyq10k3HpRxBgjbL9jcl7aI139bxBd45BKVxIhTPocTlLo2DwizY2Fg
ATRCara4k8E73+EeAyZGwpmUDjmhXxBklnX2/tKYuL6K+TsKmlr+gcwQLw0w
XjuLlxa1MnNhxAm8Q3RFFxymj/YPmBkGr0pVZtzjjBP+zcg3sfgwpF/dOU+5
3tEjaUwNNItVbgkopclD419A/t376vFGI/t1cnJ9ttgFTygu+QzQhH6+V+Il
XcR6dRjFSP1SP8f1uOiNEzwiaDGU7Jm4rL7rpRFaEozRpQhEQZWFdWeU1icj
moBHP2z8ATSRHQgX1GgblBf2HmqSsLCm7SsUG0P3cnX6KWAYta7bFI534/Ur
RNEJSPteqMwihUGMWsLZ5KGuJje1G7rfjPKEdsChA6nkChKmzM4Pi9Zgx75N
2EM/wwsSTxYkOdh78APhWeJ1csAcQAIIw8n3HU1bAX93vJfp8ZSqMfMv8GsM
VWkQY1DQCqnznLjWvqI8tz2LsEM+3C3NJisMLiNR+mUYdeUrGyDJf3uo+A8H
Wj+zR4JgrBDvUO+Xa8UreOck/x5bXtbDlfhg280CD8OK+7Sa4KvkeCGZACkg
Q7V5QqdIQEFb5H5sAz9Yyr58dTqT7nLNLhP4b+jE0BqZMPEx0Eo8Gu7SkUpi
1AHrcgmTWvymksVgsZUWWLy2G7eZOuZehZdz3v7UXoUCs8Q/h+PNtgA3Sb3C
4Ilok9+LtMtLM/pfe5cIB/qkuhS/+/O7XLC5cfCi2s8dBJ0XMLQa5yuDuMeI
c55HRgk5wdLpjRNhJaTNieB/ZikGtQK7Eld3Nym0vnYO0+9YJsSrqVPMaspZ
yh+oGWUhr6j1KkCSaJoF402wZJMe64vD0w1qJ/Sc/RqKq4H7BKRPMDDfmPZP
EWTVUrZVSw1TAd0opNxMZM+wzsIjQFKxqsG00Uel4XOlsCN1orT+19OVjuSZ
TZjGyneiQyX8wjxqDjpFf+T89C2h3gtk3XED/zI0jLfuq3VWt9HlbJTjCC4+
QoQFJ4pYQsNSNgGu05jFYSEVSD7a9oa+YndA0GM3umcH68RI7ti6jbVMjm9h
t4JZoqSY6bdhlYACCSea5jhG0hkffRJqSvLb0lp75POhaNeniB1zCqIdbt0L
3gIqi8VT94V1Qjv5LJSBku3p8zNT+Vgj1FvB19rEPdM/c6IEA/wjr07wn9YM
ozABflQXLTRjlxaKOVnvSM42EwcwdDbX96QJ3afR7JbSlwuivZTcCJ6LjRI+
770Mwh6FdCQpuR2fTdvCWJT4s0L3UF8sZMVkiTEcc9I2HR+2LzmCSrySelU5
qqFG+JHRCJgyhm2zIx2kQfXhNZMHr3LAyNY+Y4VZYzczCC8o76XSXFHhfSOw
P7dzNcqLqQFIdfD3ss9v0rDX+73uAJ54clhNBDiz+VYAXSGVuQlebskV1HTM
8xf0cnPF56ViS6KN6TEv6q4Lt13xno6E4yrQIHdCFhZq+mCYJgHsL+hWcXhO
cwmjsljDzBJz1yPxAoXV/YtGD4x7QsBL4RGbu7QXAWne7sjZZ+9e85Fw4s+P
gNYjarp7w6bVH97usPL+LNc/o8rEKV2VlUBDINscwj654JZ9JyJfPEwbcj0r
bdeuHagi+j50uJscSB9mGaLnti8vvirZF3xqmWddfyCZpRMaVMcGzdzh2zsj
sIW/7HnTKGCeSeuW3lM5feMmAypHEIPk90ge9wWZLxcMEze+GzxVgvc1Y37G
GpvLt3sk9ZwYSj93tDDNht5xTzYaDN65H923noXqAP87p1ylu0jQvLhEwTRk
zP3H2FrVDzrnpoQU2aYpK+lOWG/fcSwNtOB5Wmm4AF7hzftpk+67HPW4KZd/
87t9CcXpRj09j2Bk+TdiKBDPZSA8kqybvj4UTgM6VA7BiFMnhHHCOseM1fk1
FTcVf6HsgmKdKKHVU7AsynA8iArKu7xFfpPYg8Ai1ZgDDIl0NNNyPRYIVqh8
iNT3dXVXZ4+bJyOumL+5Jv0ZBO+uwfnfWw0g4GyD6oLSm1ikZNiOD1bH9YbO
zB3EigTpKQiDUB5F7jlwZhZFlPJru5tVP81gdebQ2nKJtKjfYblpCPTCrXOt
jlMi0sFdzKwZ/gpG3pOl+u0Wz4nvuD7SUKGRGDFfJdR5aoDxZTpZZN+sj7LC
uwMvBlSHENtJbeALLdB2SC1GgjVSJvHdWY5Hup+Dbe5+ToZ9an6dZ8ruIq/u
khoCzWgyY8/N5ODim4AmiVzfvl9zKrXYVDNQGptx0NpZvfiy/+xxvZ038g6W
cWl1OVeoqnY26j8nc46K43mQ4URZ+clknAfTLyLrWzQB/5F7W1EqRWVj5yXG
szP0XowSKHR4Q7O7U4tZxO+M1zO6kGVChmolgu4TFOhMwhlqa4zqhNoW/t9+
KxZhX7UG3e6eIGY+kH+WipPicrkDqz3uYd2bYAtXze45KChYDqr+SVL1OJDz
SVkVwW/IkGpvrh7QkS/Bt5e3VAFoAxSPqR8zwpM4B/zWbHvjUNtOTsNjqhpN
8jCJ9ddRv1AhJcvB3Gdd8ygrZcgQTHIUFe5CiLiRHsFnG4VQ9i257dc/vxk/
kPkT/I1VeKIUTRNVkpQW5h02oBxdRfX15fY2CBtqYfWBwp5p8IZmuIihwqQm
XT6CEDxdbeDCmmIO+SqL+yFnwflOE7L54aUHh2xIDDWh8mOaAM1E+16NkOWe
YWgr5vO5K1VTxC626Yis2XRLMi2B3LLgMdjCcMqS7KW8lAt59wtunukvsqtk
8aM0HPRVam0vqfoBMo8Z4l/+GZRNNSLmM6wLdkq8x7X+MsUmUeB92RXtDrsH
NIP0DAeyDvzN6HZBp/t76LLJFafvH2fkPITUVNHc51XRRb5Neocf6f8Ztn1Y
Zd029Dush469Tl6Pbg0v5L86IKlw8ya9CzweBV67Htv2NByiUWYY8cauIfv7
k3/Xmbk9+A2Lf4TtswW9Q5VSbb9y2/+MTHG/4SjoWzORcQ/nQftYBvABN35o
uzBCtkaSRCTreO49saq08vE375gESsGYzR8uhIB71Obzyq1IJgnEV0lID1Kx
ept9sva1XJLwsckIUKIu6xTU5me+3ja7Vu1G5jGVoMiOg0lZD6cLvl6ZP1RZ
xEJ46jqJX0UOjxhGttVvSyug1GyG23TUqPlmb88pJtg4OLuvvbb/hlyiyCOo
KkLV62zyrMbLojaslEL+bCCVzsXfYBqWocvXapMH9/A7siAmMQcrhcPPrdhZ
4zQULTdRR01OGXRjNVZ+18Za46hN9+JriZkGFAQDHnYxzXBr/9dkEfD/IiP6
AD77WvanTwD+xyJJCbKqpa3J4GzTR0dSN9h7itjs8VrIrowsnTMTo7bAXBYi
6R9xgAO3YJK3Ya++6CJhd5Lb2yDxYQTEt2p3wq64E+Blw7Lrcl37ycyMtBxX
rct9VVGA7/s8K5lBA/COq1mjx1ihLoOxskyZuuV7ZSZex+wrBtTOqpoicJxW
q5FDNIpNj5Jd3qLsVe1Kb5lGt3mLtArP3PtvSPw7QhND4ZxGe8ktOZgcekHJ
sRdt0Iq4aGI0Z2e0YEWrunaPa6lZsnHfWS3kjXj3F4bBeVnEiXU7uOw+b7p4
31hfdpHtZjf+4mCh4+FZapoKSSxQOpT9YaXnyx9KzSzqJOjt67JKRFbEg1yi
+Xn2/LmVhskKjQyHcwgMSBWMUgq3covM6Yt3pdeqmcTBbfnclgefWKZ+2QEA
YNfqrr+LdiUsFaycuEM6FOILQrHOs2D7UsKVbnf6R3fVC8eBmsSWWrQjen00
3/jnazLi3cdLJY1S69vKFlzWFNquHSJO35slZeczTLVWAgdVlqH0KqwZvqcD
9DqOxhUkunBaR9bGbsavTbqOGWQSgSzLB2J65SPsgQDgdarvvY60gbn6SMx5
n82mh8uWWbSxDUV4LEcrhYLVtFbZkU2DSGQt4TsKywMaMU/P0P9m2Qe/w7uh
nh/GzLyvacNSzSjAl31heQPm7QHsZFI3vYEHmm4Q2jolsEz/svOwhiq8PMi0
DmRodinynWGB13cH1Jif4Qr+e34obPpsDIyJvD2bpbH63WdmJHc1uXAg0UF6
yht9a7hl+QJcAmCajl14gzVlojT4GL/cWWD06JkqH6+tBqUkKZKdX7kL9RnC
LC3d+oa50Lq2PgMJYsf9Kn4OXa+j9sKb5CJX+j8t5JreOEpRic1I+/CiwIew
t7jFkvU6hDMHa3yIUcEJ52IHA6JRGwv0RznPQKfkfU1QqoVSTmLuhGbfYhsz
6UN18ShSQcNA/sERa8OmRHORY1OgDF5+XKAtEFKDV9mHsMKmNxyi5HXW55GX
JQH9cfayL77VFGKA8LvIL/I8YtX3J0MI0SW1gHmFvlbYNdUgK5q6PQVIWy1B
Q/5CSi4SEbox5QT/a5AtBajlm8tCN8cD8Yw97YFq9bjSTa1MYdgsSc2IWgGk
5PYY0XV15XTGreZpHWPThsKCbQrgAXYVdMBk1I/7CB2Lvp94k33w0uKUkhXc
i4tVDMyevi1Dx6XKDI2EASmMn2h5LDtF+FpRcVXXN3VKqexAEvev/cnxftNT
8CF39BkLyMRBAeu2Mgl216Aq2nBd7Tjxt1ptVJvfGlcSKM2iz5Q3VS6qBmjM
aKY7eFwVW/rxz6hVaLizn21dQzlKNirVVVcdbhrvpcYRIit/ZNK4r5k542r1
gS8gTUNBD3LgLdJhv4diOO1SPjRRYNX+dEZRdPL0veDoaxCOzl7hjjNc6pBO
Y1fqrxyaVPeYdoxS9IxpfRivve3HNdaboVeg8rFTphkvFlQiOVA+SeBvif4I
tHawlhkrKhX5LOQeNBXIeKPA4QCSS2ITScTxLpv/kglVI6+bB0BHc4UjMQNW
tWVjhgCyXw5wyxYZF+jK9i+ITvBEjZMOVMbbN4jQ9q2sR+zINspKoZicav79
MaXe7fTsz5Ni/jhaZcRHH7DeG+C+lS5sWyMRTzgsQ5TinY2OS+ZLtFq3Vrko
oBJzevP0OVG0CMhs1w2fiQxyC9nf8EuvYoAjr4Xi+GTl6AZBT9ry5idK5DOj
IfVRZHtV92E6ECJJUdKMOvLatSjtX+jn0pV/MHnr3rKXWWvbG/SMSkJ9lnoU
HfU6mKTpJEASXO2Slwai+cVx7AmQBnl5pc1A1veTS0oQTaY4C4jqWeofHS1Z
FlMNR7bjFOzSOkovspwDWzauzR9QsucH/MwSA0lzeGAttfmusmudYmsQ4AOH
V8x7kVpNtXytnDLxs/JZQ3O8zp78Bv0U+ZXZqJxPhxrQ2EnmnR5FkPNopTy4
dFWJ1nTaVqP7hJy1FAt1gq5nov0GWKYo6acrOxaaP1ol3kB274VuBH6Mq/l/
7r+2T07vxYl8LtK25tkL1yeFfpoYvwI4j4g8aB+Y04gLbbTEN9qkEDQhvvfA
gclE7th6CvwsAfIzHEmDpSWoMLRhEkmitazA0VepLPc6Q/CxygNlqHGtnfd7
f1ZDmEpKf77JNDy7ie2FY9DyqSvE9omAcs+8uY3PeIoddkMw1s3qkswyoKLf
lwQDs+P9cJvZMKAU8o5T9gziHl523++4BpTk5kLp9WnUgFj+k2bJDxlvGlKi
Q0lreAKMbj0maGW6AyrBC7kAQQlt8tIIqlkm8FLfvw9W3JSBKQs5bX/vYMN9
BgfC90RpC+qB9EfDlL4/OV1isiYMmfNjzwQFSBq1PsfaAHH6aNlJeDk0Sx14
vbdDUntJB+gxjO9D9MJ5fi2zInETxht6Ak8T8cvG4Rcl1LuZjbf02w0dUPoI
fnF6zw1FJi0GrYjxkTA2SzPAADrINJiBoRH7m5UOIJTMi8cUdMNzJ6K2mJGc
UoiWA2eq40k0YJ6a5Xx8j6W70jIr8eGoJvKvEh5IKfKnNwRC0koEuEpnX7z9
yWT6zdD2IBzb9MdKWg94rmVhrAWO7m/3yXvtZStPkz2WZG9LDNtWAxyT4Qrj
aqPyZBfY+InTe/aHbr48AkkPKV/l8yepIm29egZlo/aGT+F9ng8JN1AFaEox
KDFJt7DVqdyJTg3XZQolWlpgvpYWI01ybTzHIo4KBOsCBQbVzyQm0RLjfxJ2
kcdVfMhxkRNMvDaWnW4hU4/pRXYIuX89FDLaGaq7Fz6svReHPbHFO8O3ph+C
EYN02OfvxtpFRlPmsp+dhdFuUrggnLaHpNIwIfZcktC12fr6X/JWd9btCOiU
v0leux4+yxvA43FFl8jsQr/MHWpsa3yptmBkZTiZ/48TcOWD/O6H7yRBkW/k
GM9hJjVEt5S0IvX3cYKcPu4vjmAn3APJgBoeytKaDC8nXev1NLmuO5TYR+Z5
HtWCwRxE54B54Zv0hoY5Ilw2aXEO6kEVfuMVDfZQyG+9IxzzcLfu0DTZ2xNz
PgUBoY34W+NrDjds3usVDk0wSE08Do0AiMgdihnDq8+m+YxcOyPpVeRpRvwG
1GNuIxu8FgrwaNmJ23zTS5Q5wlfaf36Kz5a9auDP5lhyXTzdQkfd5KvFXIgu
MUOXjDWJwbeP69ARwkir2R6cHrGkfImjMyUqWD9FsVCWFRHp7cRU/R0BQaTx
5Gz8xt3VEB1/qLSdnOqcr7cnJub0HlW/t+ZUy5PQd6H5f0cg7Jof1oMC5AAo
IfwgV/o8wyFRDF5A/0qEDKGoG/i2A/3xFbHpw1UZ27NyNqghcWBiMgk0vmPO
SXRdACylmo9VRCpQiDY+O/o4dtjHmTXfL3XE8T71A7utoLs/CeiOTnKyAqTT
fLd/Fmnao+B5CboLoSSifAotIC3chypJwsgXk/U1FXZp5RUA0e9HuP5adW78
6Eku7Rcyu3iOUAcLIxTiLD5QGAq4UH457yhL+FaeE1H+xLvzuNJx02Ja/wEf
iHP6KYyHuBZIc45QZJU1HdTR4C5/JHHCm/RGesTHBcRCLfIUOKadt/B+Fg5J
YyglwsPWJ8vdbJ3803C9upLT+ElS/tHqrjjlel9VMsZzG3srdx0lW9af67bG
elmvn8+2KCfZ9GM/AALiLMb8M6ztqakD2Dx2rfi7s8ZYHv8tmWxd9AxBzM8u
p5forapFSvY5QuGwVklZCfRhBOsU3CgXX412ulPGAOpYlx6LsGOWScgbx1rF
rgF4+a6BBkLcYxbLK8uoG8GAKgivXDkjUbjO9p8X+1scXB1PH8HDAOeIhlpu
b0csMETWgUkO3SED16OBRITLLv+J18HImxhqUDowhMWMVDoHZX4xRzG/b5Ta
ZlRuu8H7KIQNUI21GinW2ShRXvTC5ye818FW+bRQmdMuAV3FuQGT3gaRXIcP
oqmpSzk6bdmFst5vG+KTSIGJdO8DfF6AkhYeDNVWc6k7P+CPktTYmLIVpoA2
vmOHB15Ab5rlKnpgDXGYFcv66XGZg580WJFcMl8OvFmhpDzTYefWAvblRDWu
V5h9zz1MQUJaPF7g+JbecA27pLNl4X0B0DJjK+8X6dTlpxId7Fl2uiVlj/eH
e0cs/46BmEabvmoS4AxZfl6wqO0qt8250HwC17sOSmo11ywrRMo/n8o3ShLM
nQAJ3tuDpk8aAPmR5urxNZz8vzecjEuQkXRXBUbu+KOwBnvBbd3QhnDT8kZR
t0K+73MvA+9u/OEYLrzKHfQYgK+5uzM+y22T0qqIEjkPFsOSPhwZya0n2aZd
u+wAivooQit4IxF0/3yFyalQuBkSL26PViIZAK8mRogpHWT2RqVDK9SYqyQg
mk38WsETz+9uC27O5V86D5b2u5U+KOoNEwEouHY0Wx9urau+1YcXV1vIhXCr
RV1cy7X7AIHw9P5HDQLGmmEikQuOq9jqfej+Rsffmm8mR5xuMpNQuDxiZVMb
O5AeO0EDyfABqUOa3F7iPE7QWJFrfVHCX2cm8ww19D29CAbEL3GeDHBCMKyb
Wc2sDeYt98UAEPmfutLnPbf2ayqX01vVCMM044j1Hel7bNsmbKVs5S9sbx+q
PGXYfY49wKcCdXPFHbKOwlXQIo5l/qqgG3w2VbuOWTei/cmAMGcYWs0xkSx0
T9tiZmhEVN66PM/zjFizmIZIm2W44wEkQe7Pu9tCbn1YY46lZzAWyWlKfRi3
kJcHYX9lcINKDG9wxsN0kgScmX15eaOO1wO/hyrIrmqkPNjO24wBNsMLiD/J
qvDOKcoNfQFBzeZRQ2s4PiepjxK5+ta+cl200iIdb6G6BR7iYso8ugVq+/lE
Ox6CKmdJ1K4dHm+pGrQ5ApLBOSacZiMP1sDhct7SZCh444GWoPJTKomS1KHR
2lsmVhjqPZnO0kBsU22tun0jVNmkkBIvJ68aKI10FO1boDhJA9F76CW2Gffd
mo3YTvrD5x9c1vWXN3asYvzvrVWLyRL2+D+m1avE9tUeVs0uULTS04yOEt7n
1XNl7ddVxO4H/jM+Eh/WmmBnb3beAiBGNap7bhQAC5777Yxqqn3roaJa19T9
xGwhFMz1Da5oGIVWT69jPJ6eLKo+4YNDPPJtpp21V/C5ZzjeSU1K9X+D1TK7
XlrzvobAcqd9yD5tZ1Zo9pMC8rCoyXBBIMW+vGAR+sxHz01VOPYqzuf49Nx/
x2dZVmw+y8nfQ5MKUncKDecdpP7f8fmEiZ0amBhmxxDaDUZ96C7UdNGeibdb
p31Wkc2QLnhteWTqog1ddCvwfbdAk5uKJNg/vU+G9F94MtugcgULWWRtoreu
QnznLEmDNxjz/2NuIFp25Rjaw7qZ2ne3oa8SjtrM10rZ5hRHf38j5Y2+83+0
IQofPx7iANPLLxcS5IZ8Mc/G1fYVmlVWHWvhUjeD+sKMy4oIVIL53ML0DhLH
aZhyPXNbXjidaBeN9pUfNnoEc4SHAXV1M+E3qg6TMcM2vJhogWXgRoO04Bcp
x2yzywZXlo9CWhQaNaTgm5NiZtnjVbwEhY7s/tPNJ+/EN9vzk4wbUw63IFjW
eZLRiviacumJewhjUWnU5iPMJxK27NSXTzwAQ0pKwQxgjdWOTVaDYTqet1m2
NVLxdmx5e97rl9r2uGpKf1Oab57VaDRLrDWqsXBUWBonLEW/ImrTm5nqNlMU
6HvtF3EbpnsZcwdoICAybxkiBuSG4mQaeKWlCzTlWg5GbDzw5YB37vYzbbbP
vGBaZJ0r1+1bydFvUMikX16SxsmYRsEneJQRoo4OBV8vXBi0fVAR+i5Yi33B
5Tr+Dz/HVMxr/lCcayShp9hOl37ntNw85ca5exYVjS7Fzk5kLsigQ1zxXPj2
v+FMUeLEQtHGtG+rUK+8fd7FkN8peo+suW2RYYFP6sDrdtVha3RbUyvbivCb
KR0x6VeLjxFMJdLYPqdv9Wr24RTeFcalhZcwYgTPloTt4jkU6P5mgSjpBtOf
ztFWZKfyJlbVGDTLLXQ/axLmQU95khvAHFpL1Cqmo06ePPCO9AtkGoRD5d8k
jADnUz5pyHJwzagRwnVVPLwwDg93kEgTo9YnpW09bNhVP2fKB9JwENFuA3MY
DzjtTs9XwMGfmcUWAgQR7Z1ZEjc3m728YvLMIV/wwRt2E8l2dZqhCY/F/DDS
JtzPl1tF6/IjzxEbnpNGP3mooloL4DNvL2wdTvyObsiCmb3XSm1m7jDVrZ9y
jb32SMGVpdZuCKnSRjLFBe4V8dvNstTDSAA8OjpwhR6EJ+b9YXrSfvRJWHbI
df1a67gBfLQ7JwfQ2Xta+p7hVDFIg1lpPOFoHOY82w8xs2EqB4LzyAkhh6u1
BDTMTg8OfgM9TKanxYDf66ke7cgKskQbNy30uI1O3AARcw12qtnuHbjFlV2t
qZQYoNCFmx8TxJlCX9dnB93QZ14brWf6thvbDAHSsSUqZMCwAXuXDTkPk8tu
PMjkcaZzFnOAsBD/dtYsK9kvqHr2N2GQizguxCJ8l6Re6/no8rZTADMINe2w
wKbop1IDODVAzDFyuB3S52/OQO84Qn3dDR080y43e82/buvuEly3lcAzKoLK
6f7cY7z4dfbearg/eHkyAHegRJRYIqs3Uy+Fd6G9OsGcMoqI5G8WxGjA/40C
/qA9woAbBijbfZMYRC15MKAg3J93FwRIqeBlSTzHr+LBhkzrjrmCp/PYUqHa
Zo8sQqU9BNnfl3eARAvNP13QDvkSsKF00idmKeK+T8SyvLm2Quvsfw+OwSp1
CBg4BIM7miwYfrAib8jPFZ7ORpgsm+k+xg8px3leQRSGn9P7KooPOzx8Td0Y
vl7d8Mf+UyKX0S9iUURmbr4nlNMyb8/y6LoT6MTJ2uH/4D/F6nJYrhjh38JG
P0rqq2lyTrs0Y3wmp0shd3lqRdOMr2ptlMMAq/SsBoBHJwAk7qLTLhxKQRKk
1g98NXL8w6/cP6zrZWPHphw+IbDMAYiDuufgaWPmnavFpgH9KtepJkukvGly
JNGZ4EkQbceJEMzkjfJCaPlPJ0G5gRicm9OzqWRwSkUAd/uSQrWcar5S6bug
exJ4oPc1D4lqoP0hzcwExCp1XZuCon/PLDmd+hgJtKNJVpFbmX6/DC+fp9nt
A12Q72uigscBv8a8+RzcW692/6VxZjydFfZQSA/G43KAZlozUUbMJeeVNVKn
jRgQ/+1Sz5hXYDVV+/k7HbAs+MJSh9fHhDIcIxDdRhsrYfgUjZPyZLPIDfuE
Ipx06Jd4q1jUdU2T/X8dem0YJthHIUfz9PQnghPN3FPfJIB9ZKWqrAzjXlMv
JBHpIrLn5TMITKxk7bRokldPxFYhnnr+nOPIzBRyD7AK3E8Ez9kSGQ5d2wlX
M5lIKojT+Vy50dyFxpR0KMnY8fNVzelvh0QID2nCtXxu2VJNm07O4RssaPY8
hOIYoOLeb7w5YMQK/ciVP8In/+AjuhLCbTE3l7gl/OvV99hoE/1rNsMFQ0Jz
d3YFbdTKZIu4UIgx1w9ZcNA7kG2iuOIItJ5imdj4KN14b61NVVyZmGdgFCqo
Ic30xN1WkWDWzCS1+V9tvR4PwOa/d6bYtvn2E7DBcL1v6eXitPBtnIZhtluf
hz/HJ+yWjckw2oiXaVBDaMCZWcs+KlLHzF7R9CF9wwI7HVE12d4UCuhV0q5R
nUJPNuNXeKX6aSeNVlw5fEdle4WoDbGClHP0MQQudDmxv/OSmodc9u7aTc7C
1ApZ8yAvSyE+zsYZdtiIypt/gMbLTP31c7w5i6d1RHd99F9gwrGs9yna4jvZ
sKSV0jrsHCnoioxETGLTFZs0v34B4j4c2uL6mOkfeZ+tM0i0SomsvaZrzXes
1uqfGEv2NdBAPoS0pahtbQlLbdbplYVs3Ce8I+0U7RNNUQ/q6VAxdL14pxv/
HMkGTyvc+Q4gXzGXPFthvF55ibqwFvPneYk01D94TA+vlwRn15gt4Xh1TcHX
fZ1/jh7EXhbUNraQEVk2IRcuTPg2GvPjwkwYdDePn2yP+tfCPfup+wdWyx9Y
TP74kFHZyTbOPRTg1WryLVyGW4M2/NcK/ltaZzyoawmuLSbHbZHq8zjB8En0
Wb3baK2qyL7bLTxk1zMV3ICL1J26qgI4wiiHdd9VuHlqnNQyMIvReS06ETLi
uCi/YrB/hNbta7hcHuzDYv0coi5nrNkGuyxF0/e28kBds53J+1epPMO0r6P8
D7CJG3i9A2S0OBtPeO5XsUv9QxBZC39N+C+4Rc2xi3zWMlNuJfqGnuZiOs9S
6qkmCMl5q2TIOcYTkQbAZB1s3QYvZ8N0YXDA6EpbucJdYsv3wiJ1DrO9xBTR
xBsCq2R3jNnrMmcI6BgKxEWOwSgrNu/ueHRyPJFMyzlyYI25QthAAeNigpL5
jchupyeG1EkykuQa7a+7u1jshvWe6Ov120qi6G8mxescoswDsmTscUcx6YVW
t2coiEF584I2S618hMW7o968emSyOU1g5DxizC0Z/LIWGnTdTXRDAsMRSkUN
mQi3V/WofBifomCbP4EbPgRaOCzXYB5eV8rM8i54kpxt5Qgd6C7JbVBawCmT
HNDU9TjLjEh0uZevVN/Ee84Ble4w3t8No4gnAj6mvQIA1OcTB5KS2/qQ/bvd
ZDvjILIoXKEnpg+eW48GutudhLRcnr3/T+6QFmmSyZYjcu4ICem3LWbbNOOr
l0oL2fa6GNNoZZfTR+ViXHm2mA/7Lis5FVjhaIT1KYxKumeRw81H6rQmBeWI
1/6Zf77kIRHaAKisc08AIxRWgaenT1eIjsCWlvjZWl0sEKZQgWCCe0eq5T8Q
JZ4bGGBJw7H7fWK80kdXlPtmklhiTzGwlKz+4aqtgGVWCz2M20KYO0Ju1dGI
c2kz6U6KZQWBfdpEYKw+6W51a0YeFCOLq7ftMoxYKdgO3EUMy0QN8DMaKezt
IegYtJN3tbPov1Xh70zk/L5QSBUFVQJcUPBO68svGCB5vVboTiipt0NXrJjN
yP/aX9xx+H/Bu2vJWod+8OEam/0xG0/8DBiRakdbvku9U2rAy2BT1O2ZLbvU
SaiIx/WQMlHM1pt4m7kUqBHifpAJ7A5EHCukNRQJaIOpQ0QFdTDYhKaafBgW
ggCuM3NS3VbVckDmckISRpawIZBpH1g5w3lLGFYkP40ej/YPBslTQs0I35Gg
xTn8PuXY5kp2mxkFsDIwP9mwTErEcntFCco7nKGRmq8SkpwdcUL0jV8EnSWI
8jPR1Ok9Gn9EvUvfsrp24d7MGPCy0pt4wefLjGM2T6h0m03ti77hnvyZc05j
88CSBNX11m2JBF/cDEe3FjVr7fIO8VLNrsQDIhpoD1aeA9S7n/QbYb6pmtUO
wfXe273VkirlLBfqI82QutV5ne6Lf3xCf2LDOOChvyMq61ND5XJTODflYAiP
EBHrNmB6JhNCcGkmTxw7x4GqvnawhTa5PvceXLytbbNxZIlSL+syyjK23+xg
VIRnuptz9AB2kzAcUJ8VGtwtmMDfn10Fv50J4JhaNJ0+kZfeW1XI/LuX3tGa
wgvTucuZ2tPkPYaaoy6XAVKbe0ZPHE/rvZ9NvwI6cuXd66phYHCg+PqSwubw
MZleHvK30yLd1JKoPtqYF/mpKILUFxJ6m0EM3nligLXEpAk7ypWpx9GOeFr+
otiiwC5xyffKKsGAWTpxGdIjwdXvL+lRUtlfvUlkOd4kBnwbRnbSbaQ2HWkJ
W4mlQzXJIZaoPY8US9StXjkYyXIRJJaszjdhwbdYdJCIE1gFF1KV1Y+hHl2q
yZmIDWs5lOTvIZSXDFqaIL654e60ueUMsABfV23BJdHQ/xMrtdu8proYyYfd
UxdhURG9AwNJ/qfy4keoPtWRxZau1MaWQGWa8Jo7wQvonGcJDet5rvDgoiiI
KCa7bA7dyhQwx9if46YvO+nHHb3Ft3hWvs/VJn6tnxk1+8TBlQ1TF6TgikTH
QgH741QrN6OwuYfg28pwCyc9oW0dl6xTdvn2YcEXXlrXa1SH/jZhSJupCVbr
36bZchCuJ1YIR2m+Bw0gN11T1ynGKEVD7bT5m9LynPe3ILORUYqV9n7dZsfT
GkbL+uOqt+o7+/clGoTxRWGx0Q7PRvJQy19Pf1MWir+ANPqFWlpnisNI0sTo
BJJAhRmeWIpC3NmU8o0Dud7QNAgn/B0I6WUae7RcXyNjVKLf1FU6c0ipWPG8
MnRxtFn2Z+GM5TGog46ykhlcv81jTxtvcNxItHlCGqKHf4F7PsuZ/D3UXQVR
soJM9KsT3LmyrO94KQ5EDRFdJZsUxsAO7OvfUWKfPV+GyYqK1cQIBKJ4Q+3X
tK4fyiXzK5V24Bnn2G0Y/AMB+ypWV8z/h4bClp/V0TXf6yJCBJA4KE6pER3D
KMxBXsnUrOoPP2Ljvu9QNRE7qLiyc3KuozsBkrAKLlj6nMv5rA1TqUZLPztS
grei2nKRCbt9AEzZljTN+tG70M+cmi37QC5dLAYccTAvWZr28b3cU5MTew1e
cZPtKK7nB9KzoO+WN9pUDkZeoS47zOxUumgJeUHqrXoHLWSTMZGe63yFhW70
P9N5HuOwx20jH0Nk2ZjUFyVPxWMBjV8HXS4yNEkd4D3jSDZcWXm2DyLENbRV
y9o9bwD5LscpFdWfK4o/hZAMuI6q2UaejXDE+CLJ/Kc+rJ65v1tTbNTUa3Pw
nUYyt+0y2Kw6I2vkhWOJJO+37oF6igNttPYQcLpdYBPoCGPrUGsqCvLsWuHV
L1ni2wygDW6d+qfpLUbbPITb6UUA9qxCffRF1Z8Jfp4PRYKc1HlwH5qe9n39
/8VwHtgUGEHnnu970nLkeRWigQFhX+GZRORPHfHKG/ydYN2jpdrXw+I+q5H3
a75wsjG3S9t3NANlMZ0FPLDcc8ctlBsD1f4mhdnWmeRC950A5qjbwulen9wn
ehTXwnu7hqDEksoRvj/M7WiFFfyb14yOiPp2wTOkLt0ZlepElAHtvS/TIjJy
FgWy1hRjx6bGUIvovukoIgeNBk/86mkalqXSbqli/w6gQibDXgSU9borpNgU
Pw0td17pRtfkOHnR6gcfkuCWlMJvUNI0WTQJ5sqa0tBf5hIm/+Ulhy5E/a02
pfxn362Jwu8+1qzncl85Q63JwthDb/Do7nkiS7Rw4IudpQtIRN6OjuSSMgbN
ilc1HcSlQQL55KCyWUZdzf+6iFOjWqrwAEa07NCjDffeO7yVynIBJD8mu9xp
4lRZgKxxvxBf/iI0VKFA398Zf1yEwfp5gmC18Og7ueMDmMTOQ4DGUrPMYgle
s9agFokDsxWO32oRFafYTcBKk2LVanb+quCL/CBLpOu/kebQ4cRaTXE0L5FO
YPDUYwURklphp+1qy5yLMAGz50CZ30hYoQw+3OBErYDyXED84y7z8xWsoc6y
OTizVrnNupTf+Bv+RgyeL6VcTAcgG9WrXBypsfFlrG0Y5pXt4saspPpK2PB7
lWrAyrN2/jBrSAXjxTFBsKjixFhOWnLeXPlw08IzJssE4UPdKJS8ky3z9aW7
Y/rb+x0vxQsOexzy7Gh1S6rmkEAUKLl9VfJVNwf0Xtx9CWSlMvudOgjK1EbI
rPfJEMq86oirruvrim1C0YVpBAl7pe+LAJHSup64+tqsHecmwIppDIg9/uBm
H6bdpt9jlCHNqXXdelUk4Ghgajwm5C5dEtDivOTQTec3CDC2XnVFKhtJWvda
xIkVDjG0AHrvDS31eQ0E7EsnHYb7/Dr7Ot6vZXabZxey5u/v79whuGauC3ta
beamGccQj0tsxyjZ+lnFx/zAx+QVfo/TjeU8p9o8dbKIdkSBsHiO50+xnRdS
cnuhcCf6YEymEQVF2fvVxbN8BAU9L8YIe9jCP5blnTRgblHJ3N/K0ELDs4Xq
DCfItNsqchnXZNl+Sgwoy6H9hJ09m6Y7ZtoAsXmaWER0vuOiN1/UasqQXf5/
6hvs5zhZsGYoNFrxTp/3L6RFljsHEiMGZ3KlSZsyyr/qf4AJJsehakQcTkKY
sDXwmWPwpPTrR477b56HJ1LUbfFcdkaRLVDVib++6DRI4RxMqZEqbhpWghHE
eHQVQECmhMdKtSJ6r94F812+JZW4N6nO0Ga8hRbyqFFiVENANt4Viap+985C
8sExJsKvggUAOrFbwHDnDiSxy82G8JVmamNM1DU1EjTSJ+0enVJj31R+K7Dg
E2NGuIpfiAJ94FN9kSQT/c3EFVKDCybFAMLBu2IVMmiBZJfh1tePdPTsrYpj
tqTFLsnqsfsk2W8oFQr+lJUxc6UoUyX0H7UUUyt6kyp+pcTvq+O0mbuaJ5zt
uLVgVk3K3tDdRSkP26MRktOo1T+/sa3VsoCa+BFJ4x3RBJgm3fB3ov/6VJvB
Ois5QN481oqnsgeO56+PeoekT2Ri8I++IbFp49hs4L/gUHOBo2h7ylXxsFoP
zFF0Sz13V6km5rCDy+3CmYPzBN8U3SGA/f0/zkS3SZoX0mxx+FC1H3+iY9ze
jiNKHZz6pmoBuptnf50B43KCyE+JLIgjmCoTsFtee/lxCpW6Pu2DrICUuPLr
A2HMZ8XSvjDsh0RGXMItgkv2oTy3yo6EVguLk4OIgWcaL3aRmsqVkReGYQry
+nEkWvStVZ1JmehN8OGWb1p/3Qe0Gw0fYSXacR4ZPPvG3AOqS2STDdavit7P
3StOnIjji3c938B98UF9+Hzy9fDnEHGMTyLmkWAX85fzMYaht8oUIccp3TYh
95jGWWReFePPde3HhtPbOiQWoOJ1m/U//2imzTwhQfQT1Q7TOOO5j2wq4+iZ
3s+cgEh5i9IVn7V0e37JgwCiueoILXKaxr/Ujf6YhVofoFQfrZx2IjBuUQBz
aD1fepMAkkCnhq12aAEP/PdDc2TAyvW8Gl7s4YEKKamvXExey3t/mCoNFqd0
1mfjy1YcO6W2FpR4cn8At/bptFGmO+mwQgb1bYs98+gjN0JBlX9jl9/az5/j
joBFpKU6ZF2J4czVn0OsVGKjZ8ZQ5QhZnoaH+CipugMxHQg3yILgoElQEopQ
pQ/mg86Z0SPtD1i3Rh6AMsaii4MhpSqB0h3VLYECn9Qr9oUFvNmp5Akh1EDT
kj5cCjA6Mx0PTPmYRJUjFZquxGEBmzFtUuLkkmCPY1whwJYbrnAtPFqi43EZ
NRMQe5CWuWs8413/DDDLWYp3nKfOqACDrws6ItnpXOTBlpKVISVUkLsK3M/J
gpS6n+sdLXum9pHRTWkwBSCsyK+nY0vxnIUetqaauDXGP4D5lv8LP9sOoE+J
09zdC30Cxt+2m8+ISTPyi+ok24JZBJro8yWDD/bPqSHsKgz+LOPktfgeQNKD
Z06mV3QnNjTYRFBWjsAJrPCnsuXF1P2bUW93S3da+OANP80THEjBN2hgsCqC
ZxQZLyDSP0rKm/8AMfsWJLTyPIBqGHRbr9t8W4YXq9Wwt957yqvSDdl8u+1a
bS0EsXDVy2jWsCsdSlKOKx0TdT/AkkI9yTOX5RkcK1c8lOyZ7SQlx02IpDcf
6OWnq/XQ30JiCXVOMNtu33tDQ+vTbqjubybXqcJf0BtPTMMuTBTr9NPthQqw
GxdT0rMD9IJ4NC0iJxVCzHBVrrO6DFUcZFEYPOBm1ZBUqAo3J7dHKn2lEhz4
wxGpJvx1elquvghlpm1dhKsOdUkyvgs2rWrTaMayEN+qhDjROkb2eZ6L7lb1
CBw0tC+nE6TpevxKoYO0/RfhJ+rKxwOz3BbAC1lP2UwK9FNYKUNtec+nRNsO
ZBvayH6S43UrcE/+1Qxc25q2fwenvI3NUsyY2/mexQmKMNTutrp7IGPkGNjP
ezaWoVJ63uRc4Mq+OmSt0ZU7NZyKWugPSY9sQYTCaHdZwdgQ/7SvXt89zTY+
B9vcVDpSMQwsO2NSU/xVYPXD+Jc8/NsYi9AnLdmS0KFFM8bEY2L/V4y5sPQO
vkXHUUrTnCHDCl+zKSVUG2Bw8azmysiG7LGnR2nghrT6Mt7H2aT9mdU5cUJg
B2RlmIBQ9rK2iB703bBF1oTEZqwYVolSRdpEjZGzIihFDl1kUzDCmHdpjjbH
g+G6AtvQUuaqtHtHmvNsh4+RjEOjKgRxuxw98kwn9sbnL8GbMbx1PyMkvexy
4+HVMHUSFi86DmIMng9S8R/UVXhJ91bKoEjHHVRfcRfD6i6Sd0E24LFsGaO1
IeTsX38G+pJE40WemTg5Gost4eltuPnl7c+PaUsg6XesR5Q3pnA3QjV2tWIV
rry+DiTtRF0HumQiQDkTJwM0FoXSRFb4q+z0gnNpK6sk/upLnyup52RHp3Ie
IPMEggXVWqVFDXePMIQdrN5TrdCFMt6Ty5xophT5RCfQsCEKbjoBuJlissqy
rKoMVJOpi1gmrBTMFBOiZjEcGM7xYKwvj/wfGUHvf7sMfyiHoBGr5x/cdSNc
HaE0L23KIMY68tXf1NDKEkXAfBzyY+LjOcrJqTl6e/7CXL9XcGUjTxCV5cem
u6ssbpJauLy2OkANVknNJ+rJygPPF1iLfUGJS+A1fikaXnfRQlQ3TTx58vWr
Ey2NtL2RDjBjNDf8zpu7bJDBMPattSuCUZu6iDoEIIjDPLqpJR5hjrk54aYK
uWYq/t6CW39/dO+csawIg3Tku4RGOvoNaCU2e9KB0glcPtRHKPaLSbvJXzx9
27UQKyZsWdhKNcT6+olDdU8S8tqJjWtvrel8Dgf95ETmVPsG3YO2oUnfPKmN
54rpui20ze0UlxgYsp1VF4kVUS3xDiGQXfvstPsOeYWMkadK5wPpXYFk3j3l
RkAv6DkB39LtwHCiv8nf9B2rDKGj+k/Xw3H1cCIIXpb/ea4pEUQOW1yr1WXM
AqGqmLeOBAUvYgYTbrTBKCeMrFL9Ct2nW+aUcHA7EDY1ZHs4oqOm9RSQLUyt
uCxHyD6QnAAEdayClUixKWM06Xwct24toCQyzSu6u2uO4Wj4j/u265yO1PG/
8vlemcX6LGKnDN55W1fW8RQtKzKJ6fKprUTdG5p77n73nt0iXWZnjKDuP/s4
PyeY7gOnfEtbM9BT/95rpS+NlrQ83LETRddtnO0hk57mddAYiUERZ8w7XcpY
meexqMagC1vu+ny050kmnDclEot84wAuXI3szOYJXqccU1hWIi2Zrgs1E+Al
FiCH9d2g5dWPrcDtgg/qVdh7q9/2yifDOnotRs30OAQwc+biYYccwTC6ZZk5
DEZdNWZEFsKLNWJzZeB04MqpKupJe6E9dJBlVdKBuySa9uOAITdHy8GM91wg
r7aiz+kgmnbO1cuOXgsIEIDWSnuGcukFh1wh2ueE7AXg337uUyuhXAkdShSD
7aais/Dtpk927TpcPI1v/NmO1Rhb6bHNqnbleCDYSHdKc7cGQm+f2R3Bz4Mb
ewA1zdjZXb4BPXhfI6+td6t1g+oYBbwIFCo4KgYw7cZDNIzLYpRYyyEZQlvh
nMkSpusY1lK10yaIG9rXqqNY+Jj9Yban5OwALQbj7/H1txjQ41XvWJ58/Epu
DjJBqXxNgeAILpNFDypIgT+Ra+bk3MChIRlRyBWjwLPG2Dqy2o584zKRtlBw
w0sESX6O26rKbSHkWLchUN+M7tKjfwRs4lCs3JlqtA6W0JgLVkPLbffjRbR7
SkU7lPg4I547g+MEu9CEKNYp0EZ/hZan5k9nWIn6WYxzSYDlKKSe/qAQ/pbq
7jLM88FSg8bjIf5fNvM6OyLVAac/j/fE8zDRf0jsTrCctGKSy2HgU5y0qdL8
7Rc2E9/z0JqDNTsUh1erD1FRUFJsCzrhUzVAUU4diRq/3eoo+wko43z+iyqy
WSjGZXX9syS4ZrMtRCvezbxxzR1INk5cGrL2+Jytr0x/RMCg40j1whIyI6oc
p4JMY/L84N70w4X2fHgn5ZZfyxUHfgnNsTVGWT7KHwxyql/xXa7Xd0tWYIFj
0pubpaVeNQNaDQR9gkq+nbczLFId6ROBapnwqyBsk4zFgByfrdkdcMVmQ/Yc
SU8xg9NaH+r1wYjtUwsF48ykzFhJLgPc4tKZEm+qxdtFT7uYnTQvyAxBPPM7
/Pm++ziWhVpuHdAn65qw2MkmOGh7JicLUdflw2ZtST7u/I3wE0d152Mv8sX7
ZDQQ1Xgh5jwY4AAXHc5t+zAglH9RQdkocY/+Ki8qfqju4jev4EbHNPeL/q6C
5uAzyzEA87TGI9HOLxHboNtnf7RTXLsJYFdlqG/p/h6192B4ob5QU4UEDqRv
TdnOdoleKryMRoVSmstH2kA+AbBrupceDHrKzVaH1Zj2rTPJa9OycdlVPYBX
BGxu+4qqyza0s1aLLvOpt/2FW+5S7fmzou17LcLhD3IE8ijmYoK1C3grsElc
Tp3cVT7rVHw0EUwkisL42xyk0J4cAYY7XXwtdLKegqhAEip02584uf9k6fHb
i+Ssl+70/uHy1ZgL+Vb/zMxxIvzSWLyAQtZIr6f2pP9QOqr/Rufo/3SOK6i8
vOoSjYzvOuuwRzT/V2BULQrvMz5f7umevvq5yZmmi85I5ozvbY7nMDUpMXtE
HOW+oWj1fj03x94IQCUzlBrDLYoWT95GJ3Xvwz1V2PfheIegbOgLL5cadjM7
miba6xDgvbgZm73Bs1CaOQ9+6/xpzBO33XfcvY0kY6IQR8+8U0FMhbbdLOg0
wawtIy/0IHANc7FV273jAwD11UZQO3xxOwPKAGN8M/USzDgVWqTgt/pGcS12
AIoxb/DOVd2f4dpNTc/kh9Um3r7VXlkZVdOgqIGzSQjtUJVqsqKIsfHNlkxK
kpD433CTw5jUkHUthEz+mpgMj79RrwPpXe7SsX2+GUMFJm02/wAoPSyNLVjL
YTSjgcKfjhu4cbD2i+6KvUUoSJF//GjQbfsue/e3kEBs8M7KKMcJsb0UtEYH
3sx5TrmT4S8ftEBpeD7hCjPeNPCYIH08XWYAObOgQL1Cf1f0ivxR3+I1lAa2
mNFR5rmco075dkKzCw4nja5PHMRvAl7/ruOxqpBvvUN9Yn2Xg6EqJphupoFE
576Py42qi1YKB5LyWUX7l1HDSSFHCUM+KRuDeCEajjWuoDVk6p82gnmZ7ytK
nnnT+rrBvtWYTsKBUYMuk55glpcGj5mYqa1TgF08KYLleTV9Bqsy+z4xwYf1
c3I4Nil5YwNSSpKrW4p0MonXc9JI0FRVcnQgEqzhUCRXxRXFrWzgAY3DuR9l
IOvEb8LMZYcsQjZkgbqmAQGsojobGQ0m2fiXrxVu6w+8ZbtcdFAlCymuo6Gv
r0x+MWQB+VQceqXwFRESokMY0+4hAMJELp6xgRLsA+xGxBYA3d87RbhYgkpZ
56COYT0ieuAYLhf4gBwQFL2n/HwPhIiMmUqyGbcCUvG9cs/mGvUanPnjagxT
OqgPLntk4qWV3FVc51fsTyErjgLKZXuIbZKCG5tNzDT3EbsqhfNnQxCNRLxv
mrAFn2rd3w5pfcoJTqXjh8FznoCKLT+BmlgR6eiP7Uf5NLw9LRzjwa8Exv8U
9Ivb/VdYqDGwpHSLeq09XIV5HUIO/D3ckwB6FL0aw+oMu5o8IhE6OK9q/S/m
SMhT1XDcGQuT4+1Qhy2qi5Z6lLH0JHGcrUFU2BtTGk2b84/f8j4jtaftpaxn
wfUvquapl13vBR6Ruq5EbOgB7fwmMS2/aAGTR+n+l3v6WnccO7JvodNdH0J7
MkPN4h4vCR8M1/tbMmRrkCl2xq1J9OGywcc8e28yJkT1Waod0TD1Uh6/eSvY
Kl8hq5mJ8NUyKtbGAqBF4Hf2b9cbg5qLU3ZzqpvPtEQkKKZtYEGRdoiTSpQE
hO9CbLd4GMAaIkiLZlZGw0HctBIj+3okN+mzW9J28sR5d2uUaFWY7+gXM30S
4dEJnewqgjLMyNsL45hkntMslNGvPf9YgrNXxScwsA0wJy/k1liYnbc3Y9Of
aArAI860FnoVLKX+o/FQqUy0GvPVnn3RvgTBzXW79u+wOfxzPQ0Y+sFo/WYj
dz6x4vpxmhehmujzzfasqvCQ858d03bDGo+tZi9y5QnuFM9BDugeILUQz3Iv
2+YgMvcvKo2v24dESK2JSIY15MmrWvxjPdseBSrVKizukvGKp/4rq7rnt8rt
4rMi+msP6JhqljH+/nkrZPxb9iw0D1wM/4/ozANcE7HxO++HAn9x0tXL8cAU
fUFa8nO+sQPcCmY5uU6NInnYvn/A0/jBUx863COdJtUpgDJAui5rxEwEvEkT
9uXcqENHFpgauJVXOO/XlkSAq822uA6gibE5y2KTsxH4XOmZPOoIWL1hpfvy
esKSkc1OHiPItLASkOqgeqsyDW6pOuZYbl1orsnfK87+lrL6KLz+rm+WJAWu
IarGpwks/dAvFaCOjzNt0QLtIs+1YWiVY52oyOr9L7uTbOLg1j+5/7dyftAH
OQy13iEGMdSMmIenAeTByg9F+8w/S/Ga9wyTKRgSQQIIluVnD6bW9h8eIN3Q
LPyEfAfmBPYHhT2MRIGj6wF+VCyxMcxg1EmW21N0tcnF+QEINSKBALdCIskf
oWxZzrFAYvUIxX6GbfIueIeA7IrLi47ta0SHQpvI54VQH8Xp03iB8Ma313VA
DJRCoUw2FSxiNFeIBaWzP/a1WJM7GIWcZQ0EFUpbhlG+k6MXpBLMOnuQqRnp
0AD+VGmhm6hFZ3BW6JC/YBVASPUuu3BLzjJsLMkbH0d4mTlu1JSNzUuLHJ9E
Rc+FbdliAtoFoNDOrx7XPwpTeGVZ8lPLaW3cHnzhc9rT8Q9pnUzBkfJyca/e
sY34HaFtgcv+Ta2Ux6xYgmcGIJSZX3s5xDnyu5T7/Zg7xTtRdqTCH1icwqCc
pj6BM3bKSRDPitoO9X54yT7smtOuYpSNHMgOU3Mqm9d1WWQS6lxSf7MrRSwg
8ekOFnTN5kOxGaALSTfBmy+8c3cLV9mV1YAsyk6vtPCjG7D4Aq7LNfPWyZuE
qPgzT6IRKu/WSBoTOyo9wDiLLVqFdQqELp5CHW0f1WjSLUV2Uy/sYbZxJnYV
A6J4Q12BUHNKyCoySjjqKUcIRIoGlSeRb3a8oURmj3Rpa32mpB2yerZ5WH9K
2DKvGKQg9+SL2V6h2mnxtySYkxhEFKd6Nq0AXGt1Wm6SWpIh1ukg74KBAEnv
Uke/pAG7Tv1jTA1kR6FOTvA2SN2KnasByEFRKLMzMI5dVlNpoHV8W96TjNOY
hfOyLUIEtufchJPe2XfJWCRJpZclsDuqo9rnXnNZSRq9U4EMaektoNjLptry
pHWFdP+OJN3P8HfMtcv3MUGuLGkHsFxOT3c/7600fCqwmCgoCCLwRyz3EEYj
WAIp9iTLRBIaHrL2YY0uAKQiXW9MmhJOA0rW2g/kAIo8Q6eJ59iyCvZ0jXAa
fqk0R+cOqT4g2xedKovHHkbm61xiN4HSuw4xbEuRqZWtQAWJuFLtVnzP2fEh
EVDDc88y+VOKC0DrLthZ5oMJUFM0NNcofKuBKoWumw0HWmEJWYfOW+6YCPbO
lJSoGf+NBzG0qhpL5ZywJUaRj+orS3xRANgtaeZOhKqSn2Qtca0GPkJaCVjW
SkVKAfNhGI7dh5wQvzf53+4XXUaKa2+4OxNkuVmeehRgj0xkQa1tFWyNwC2k
C5qnq3Z+kxAhzl8u7+3xP+dpimL5tjTYBclG9N3Y9lHD6BKi/L2EzDr/TQRc
Hmvnf4tipIA6/tgQaQN1O2n2GRFZjmXHd5higqJ+Thqb3Yx2q7UANP1jEnVZ
iFaUq3T1+eOSXAKm6w/W47iWCI1SlCdW+EviXSrJY3RzS+082GZCCJGE3KZ6
NtrOkrpp3V4k/O1IuvHOpZ6Cy/uPLV6xGN+FzRpP0Eyer55pH+xcNncSJHsJ
Uj0UwU4JEqh1POVfbraUwTrMMKDZSEkneTQQKOPKhSH2SpgbWaxsm80bUjQ+
FdLtA+ua0Wf3jNl0ZZETDO4Sjh3qVRbGehutJgRCn1QCpZzYqCvI8n7KDspu
8qXnZrtP6Ms0dXi7qRcvDXSXd4TPR5xqy0wj1vSGtDSWKECmNu3o5SmeESr9
l43kAiblKTRiWolFV4AqeLCjnkjtZnLliN3la1j4VQacU8jwGYQUnWx7G6Fe
lpgX8OoMr+L2UL3D8GM1AwXnZI5wlKHlIkC4GV2fs9SukwMZcIDPyCkbHBRj
UdAx+yRFBELe7I6A9p1B/+0Rx9y+cojPz4GnU134GoFIUWg0Zhz8YGB8JS37
+0pLRHHgm9I6Ai6iddurSMYQyffsihMfopKnc0zK8SFxwV2YAgIqnoN71FxH
9eaXqMSGsrb7momcHYMJLcVqJwt8he+axbhqWgn0vpgzt5+vpeCI4gAQE3+k
+paubO53RpCdCVj9d8GIQTNgfxRAgPJOqAAw+vsf2qwW4kNmkqS2yDvgfTb2
5ImphtQzq5Q0A0xRUscuKsO91aCC6Uw75/aNgUMbnlm3fXlFdTYsHUs49Gxj
DyTs8/JdwZXRdeUkN4Db2DrImrBoxlrnvDVMAGrghdy3neOIb2ZqB6SpML2u
JcOyZXN6YMAlzvn5WWR1zj2Y1YTdEmmNGM6gwjQ8aX4nIWFTwbsGK6Y4WIyf
KIkd8AfsEffuhWUQcOr2bMueaKE9lIdNDUsBIKJeLOF87zZhX+8tsuwdSMb5
cbWiYGV/RzsNAKifdrw4lz0x7ETgUmLfGPjKd31C1zTWzfSq1qq0DLse095M
XCmV7g36xN0fxxnw5eLPk0wQaNLcXThj5IC7jpTGDfKVuQIOlhuAb9KiFybB
U7TYYWNwU3t1HjHdQbZ9wUtgZNa/BRqtIoywkUZpJNBLjQhhdkZ5XZiuhsM+
skhyBM58UFXrw0PrnTVrvAmlxJQ8eAkewg+2s6X7QAAaAEM9r18Xgb0mza0I
yBXj7ASFyX330Lr83DWj0HXgAEGIycByunjCBcAHUtRUU39KFbfNS7yu9ujm
mCGBmZWjkRZrZc0ciuTIFX+3I9YavVIrroh2CVmSU8gGVFchjyC//pcJmpTt
vBooYbaK9FMQXaCmw/pxPftuJ35TozHYMcGPwX5fV+YOGPd3sHD1IiXNNS2t
Be+DyxOvggpvEekEZsZyQbBUGRYp9HX3esHVEK1K/iAb2u2li7fbLzcNfjED
FnzUxwCAXB638qlwmGEu8ScHbOZtd/68LVp75pRHGtBDnaJHX0gvkARJpyFi
jqziuy5Afx74lQMIZ+8R2xFnKIbshLDjyE1yuA18n4CBjeupx0Qs+OVN9O6V
853dFokCGAd6/mnqrtm6hGv+QSu1+FCvxrVlFo/3eQz+EGsoisiKvVKfazyp
fcvK1cBZpAT6wDG7CoDbHiYxHv6mSVO/0V/EL+WmiZs1UyAafPU+yAmA0w3s
EbzKMYE4Doq8EScnBITpzLX/PawwHxgJounSL8pOraZOgaUoAbE1ApBKANXT
l1uN5sMV1MWBaoke6k1SCgX0xyqd0Qp8cqWYtfd/oDtjqC+RF2cY/Gm4Oj52
vUf2GE0U+HxQYrgA7dMdg/91ltu9zeErye/LZSFWSFtqWp+eKsLDxkkKAo22
WcfR11lnSAUz9wOUdztfd9sd1RgkL9tPkdvLTA94ZnMFGqpghCBgXIrHN0W+
As9HS/PpirFApIQSnZCAb7+RK+3yVBMdppQ4Zk0yRJM0ms4EHffckoTe8QTg
6OZGsauOU0RZtOeg4azqSNQ/uZN6HHYx8ya3qFpu8rUgOizdtv39jdFgJZ27
Zwy3iA1PVgakMHydsSEtmC793iE/s2EckWrxlZ95pS+B0LcyEJxhCua9UKGP
UdKhG4uK/E5Epkc2gzk1e0lG2r+H/Y/vd7Snvm6OnWUFm1APWL22t77JpuTX
R8PTAB2QAVda9qFENCkqkZTPd35RjRiLBGex0p3jTHpo4KJuAbtPjzlre9/M
aplFDkpJmsdbY47ZjwuPK4RaCSZuId1EuX9tP7LjoqYwoXdY3IAjzCffn0B1
d6J7RAG/tcaw5DqUscKq/yG+GZ+EJLDxt1KeQXucLb9sta2jl6w1oUwXr8X7
/ivkigpWM91+L74HQPqosShlWC2kGvuvX1u85yuVD2GF1FaQZxd6wddGopDO
WkSVwpEWh86bv0U5RN56aXV0n95Bbv5tXtpHnH8GV50Vnn0MAygWC2lrUFBi
1p39Xz7ZvayTtLMS+Cai2ShFOgENCGlOOb6PeAu4lUKOR6W9Fwv/ooJ/QgYB
bTpQ811tq9WNiFiT9/09gj31MN1Ixk5tEv3mnK6RVxdW/UbCz1KnL/PgfFq4
H+oa1ojT2S9KUjoP4BYokRrfwFESU3Sx0TlaSTv1kYaMbJHL0PbpBknVwP3e
tqzQd2+OmI9Dbyx2Pxc8OYVRvBV76hkS2Fo3e4MQ1gQv7/zffrlhKXpsrGOB
qQXl5Oflufu/QfiCFl0iDYtTUwqKwumCNt5B0Y3WkRcGR5m+CVYsreL1jzyD
lGgx7WRMpwSO+AS8CoJL68gr7e4tJb/36khIFT4HHE/jAC+KyLYNqfoB/scZ
0QP8IqJFFqdtc+FvQn6D/6/CAWpTenYje5NDtWecW7HxWMG2TLFeoFGpk5BI
magBHIanHZuvG9br3aXRqCcnO58t5NvxSYCZb1jkkQWs6m7O6WHm+U+LYmVt
SRLKc24zpeZ4E9mWlYL+FMVemh/6n285RyBOa4bVYJuzoHHPdBVtIQueoHwM
d2YJU7zYkTxT0lozUOFwuQ7IDWBPzW+lhuUcQau7N5lNgL6AW8E/hiuGvddq
Ad9guYxEYsZhOasq0jf7nHGfubDubaVwMwV3BUAhSUR5RJMdEYRBupuBrPcj
lNnsT+qwmR2BZGIFJGCln4YmHWbmwmtaxphVfadcc/OyvcY3c8XV6iv3jmiv
5TJ63n4vNkSXIObsPVxpqz0+6eZ4r23WFLwDLrZGAXaJ/Kxqj2fOBs1rwGTo
JVk48/wp1Ezi+biAL2iYHPm4ZY98a9gCRoo6lLlCJRUxXZtCPfBjc9yxj+Z+
Cha8//R7cc7V22ZjdYecTT3CYJcRT47Sfbrj0CBJho6XTqkHILwy1pMUqWfL
tpmCJ/EsKMAWotmjqy63IuaOI05rARJPLsTH/Kg2KPbZg9IxPu/L7W9fns8G
K6bZD9YwLsygdZD6pAj8ALFYPTYT/71kPEEfhOz8h4Y+PVReULNvHFpkqm2I
ImYB8eSapKeGTOyHE1vRCQstNnEEGudlhjY8IxiDBJQHMWEUroACV8HlYe8N
/YBtRZqcg9zRPq6kxWhTBGhH1e2aaA25qyyPG3Dk+Laajhn3abN89IT4Hg/k
6ZjKjp5jk4xqte7w+JICnuHYxUyEzA3kGun+AATBJQRuU1+BMEyaQUq9KJ9u
JZDjdNKHtQ/x17AWUxzSnBsDElgqEL4MRDS5baS+peIrnNWpKxxpoW1ARzEB
h3hyrqxp9ZkY+CobMCrdyu0UZL3xiXhSfmCNelJzYfeeiSMHByKaWA8ik6rV
bX7rCdiU3tMC6VjlI1z6oyseaM2QUm280aaPy6Ca83jDyh2cDXnvTMskLwM4
QpbE90DCSi4b6qUZ3+Xq0fmXzkEl12dhJN6r+YphTRnHnnnCX9L7HwrGHgxM
Jyh/jcWpM7KZaTPOWczF5IwVETHbu1Ya2k5Ocz5psz6MPC+EWSmdNYeMBPp/
C4SNDv56cjTJ2wGzIsoimoMU6+IIXNf8I1MJTdTXUYHWId09q8QdG3+Gu3SJ
AQSzQuQ2fft9fmu7T9uGw2OFctX7C39iWM7g2pIexYPo6iMCSJUWFEL9cSXy
QU3oqm7tgNbYV3/fHexAJl9vcIAOeFpUiSyyLlpWCLdIp8vqgusBLi6ACPVf
iznhbNaObWU3VfzL2eQ5i/Y5pyDBZJpANQmtFVuMA8fF85DWm9EAXgDa7oQC
mGpKFQQHVzf/jefxu/3gFKqz1t44MihXGK2eCpdPiDvimV2MSuhbzkk8jFyx
GOpjTomU2uTsamU9D/vWwPRxCBWrQ+iry3Lr/kgflbzdR5vP94Yc5OdV+TYQ
oNdqIVQxImkHG2ZHswDb3yQh/O280TO9J+vv82TLWaPhL4lKYfG7SrLu2V6d
FR8gxusjWzsuyQULS3ohGtCZy0Z3O1QE3GcH1b0vj+mmpVbDtD+wOX5sX7RZ
ydld3rN89CeJZG2FWOG6xhG0YxbPzjaUKTWPIQFiNK0G1zEYsGOCqsOJDqIU
HWim2PR23zdygb+zrj6rcws0mXriXI1BGYDjHcaYOIKbFdHJW3QFMK7IBdkL
7fIbNYYnK6G0PB8m81Xb7au1emk0xwZHbTBt/NdEJ6+l3n3uwZ3kGSYHuiBw
X1JIpfZf1R3w+LHmCAxgTNv7Cg1kKUimmO+RygIFR/4JN7YkEF9cZIJFwVfl
54OpkKVQnO6oFOev3I86+od3c80Pu271orS3pY5jTj0BQZgHTbHRzuY49gtr
RXsJ+WAwnt3axpzFIgdJZtKlf9ktvqTusNVPiEX30ySbcLHF9OOwmeg6+n3+
X6U7YWVySPDhmh76sfQRLk0ibkBqQiXG0ZR3j7USi9bJ4pTdJ+k5KJ/MoNW7
x9Be22tF/ny5lAH9DSze3JhYhIDTU5/a/2hxtu8dawoHY772Pjlpl22ogtXJ
hy2r5+bxSD9e14o/JGQ3HWRmKLidGcefbxtz4CgScR5IiFQhv+6bMiZYzIbB
tRQkhoGvcrlyAgtUzmJravXEtl2mHa28racRW33BbwSjgkN9KEIVMtXuMYa6
MVjOgFdx2gKz9PK/rsfSKJ6tTTKwUJhZr3dNH3N3xmkcGV2CuYDZgqOT3Sp4
JlUiq3uKoi8z+L8wpefO09qp/JCW5E+M2ltRd938Y9rB1VfaIK3cVQOUhD64
JzixjhkkL8aGVJRKIsV10wazCm69PXi+N8lwu1tH3jloi0rN1vLHQHnm1IGn
1cqDXKyyNvddltsP/vqbk1iV3JyCD+E6c8DuCh4QilbroeGyCZUuHroik9/i
HrQQ2ZwnWRporv0tg+24EF646fNmPP2PR7b7UDnnoE8eqzoxFNPZuMNofbwX
/JDfmXkxwmNCwj3hQJ2Vho7gmEyZ5jaqW9j81C/P/aQAh9K0JOXmnQ/T5/50
8888BCwtfv8ZVaRU3j+pcrhJwnauCASjoSw65LiJiEIPr1pzNyJVQXkGt7L7
KXUTMFP7ICi6mIHJ0vH2a4XZPZ7grfyFFDv78X1EjWOqvxkfohRhmYW8MDEh
A0ishRnTFlbKHRzPut9SWi1ltDPL13/4lhJVUwgnUEU0Zu/xD66nugTdRGdy
a1m9PciNCFmxp2LeLNpA2gocWP0Y2UxDw/cy/X6TTNza3YBBbmUHvgcf1iQf
2kYHB0PhTRPnRqc/QyNQhNtIPZXj8pPWfiLKw4yPm7nxOh7zS+IsOxBISmmT
kuwA2/F9IyJjKTybETR3EDwu6fb4SoKKRXPhXMCVSNu7tQ+RSUH8wc/sgiro
Gge1uCDMjpzPlYc+gd3zVXqAJHlee0VyICnJepXvfDIvAJ+p4nYs4iww68B4
WDOi2rmFjddcANi8yvvKEQJytaKSJYvNjLEoqww8YdRuOiRfMBeUTyjlEYee
DomcjpYwcHdYVrM2BcMvzQ66hNfQu7y8nUaxpYcsq/NCvncYpgjzgRoVIcy5
TeN+aQboBtEKllj642jpHX5xycEZ2cWtKkcVi0x9rtsUNJmwzmX1S53BdYZ5
/95EETPHS/beck0iriqa0y7YtqIGHf7Fjc6ZWqv+ln6VZiUWARK7RyNkn4/b
uvA94HcDJ4ZjKypKwUaYZvVOSKM7B2VeQkupbJXgiyfMp7IlQQUoW5TUYIZB
pVDJHpTFaKI4slZ1tymovgnJkUFSUS99eqgO9WM1vp+nLfjr4DBmMjxEDal1
tUB8C/iI0JcOEFr3nVGA9oSHhU2K/LRlGjQDk+hpzh9nML3VOFy5EfFcHSVT
JvTTkFy808Nmdcu0px9e7QjnkyXXk+dbLTwHoXBuW+GXy9h602yANtmZsAf9
cmlM/t1Qq0Z37/TKuo0vUNL2XUasKjrw3MJDAtYLt/3WokPsClSrsGuXolVZ
bOVc64gi8JBUcvwvRsF1FGHEy9C0lv2GutSzvgWAsw+g8nRj0EQ1Quone6xg
+z+MUADq5hLwNmvqgQjp/5ge8sfEYFGZoMID4hKycdhM14Y47TelPYlOt4uG
VdgTY3oi9PZqrqJ2y4JGK+vfBsJq4lsuHV+NLnlT/+dn5vD8FUxTm4RnFpcQ
k55goc7CsuX9IVpEcZgsOJFynecc75R8aVe5jNdXpTcZkZkkaZXZP8f2bH/l
W8wOESUlnzkN6woTJeVGodWqvpshYQXQFhMjd9pGMIE7t4CNs6KSIjB5sOrg
h2d+R5q79Oo/NX7NycOeYub2PtH6RkgLfEqdHOZ+NXg1y7AcFORDCQ36EQpt
XRfnfEMvyTPRKHWqw9d9VZV11Tk0tr/t+Ff0f7uAzyR5FHE+ZLc/Y1lkC8Wb
1M7dYLIKhpAF6WFmQd9Ebnq6tsa6ANgGaQfjqDzf8NyGQE9FLaZkwdtEjLER
mom2qgLW7ZeOGE7OLRett72fL4al+UKfDq3N4YrZbQgPlY12V119vUPEnLQU
4FepR8Z+2BOBvBihZk5tdgxiW5TYGwlTSNCHxQc2DFOHYCWTGNuyXcmABtym
aUoNVrhmVRlqnHT9s9kUd26ra/ZBUIfk3dg/5emR51+/HADT3HYvd4pZY/RL
hnMVzTVvNRvIBC2Hoz3W7KmXuJK9/BNcGwshtDC+OziLTvH/lMm9rwluae14
HrCUrXNza1nkI63t7pkXdYnuovLXSqTwFwlGTIhIs6IhGMDvZv0FhVQoIs8L
VOp0EnsbZKa2wpYCeTS+yUHtVZrDeoZaPLMfWz+mOaT/1ZrofMzow33HTQFX
WF8dnNXh0Q9NOfkHj8biLLS6wIeRdP0itwGvHm7lmW8xGIiynMDWusoz4HYc
nXBzVFgvLyYOUphwkVE5OmmMVEVybjHxlT6/W+KeieRXOoXprHOKzHWOnyxG
TTJjAHGmmcJb8+VGQy6xKz/U/Tqt87pklxOUO66s1Ufl/4l1qswZ3Jc1Dx3h
BqlS21K2HV0ciab5b+Zij9W++dSH82KYP+YECa9AF1l7dCIHyg9KHNU54gDF
JLZJGnbGtDFeHnpHjHmWpWvfNv+fU9xQpLiQjIQindH20EdV3DKlOJptq9Ay
kC6RlFXHuDYfXcCLIpmRNLlqHHJfxUY/DD9RhBuxf7hqd5Ll4a716c2dj9gy
Plqac10SL9QfltXk3khF9fqLcHn+FMzVtwWwmifpl+/JU/IzW0uHq96AZPDE
8tBypPD9yYh76RT6mqf/xcv3aa3ZmppCf7KBX7f8wfamvXPlRIhLUXPx04i3
x0/ltxDqcEj3ARcnd7D8UIL41BF+vvEojl3df4WS8LO5TKAZOjoXUZr2fMUS
OHhUwbPGFNUT1Y2WtdKrf3qutqkouJm33OySB2Uca4aipgF4vYRwqMam/RqA
EnZxO6kK53/qDmv6Ckpk7zkNJ2+F/EYskZ/ybGD2J3MuAK0O5jBrGNcyl3i3
GxIy600JjYYNGR1ascLXDDGRapv2phEHIii93B48AXzNaiqo1rOsVcOz8gOW
GE9I8n+j6TJ0nlfDqUzcWCVY/Kzkn8ucIkKmZiqKxXAKOrkBCFHBcH/yN3bC
DC8Rt+7MIQv3hbtjfVlN9K9cclyYvtmJ6oJ3Q1dwHk7nOoATLgJit4WsLY2g
yBch91Z2IpTvGWfuBB7wIy6kyz8ayG2dnYRsV220lrF1/H5OQFVatpPf0lNu
6TdLVhaABOa/I23z4cBK/4LCl/aMy4agMAFzU3bWUdwk2gB/rF+c/3UV8s8X
HrjA8KxehvmG+r2RhjiuW1MQeRg1rhOsSeK93qT8RxaXAMzmJRuyhIv8Z32I
GwjuxRnKdGUUnWQmw896bvWWqHlNx8ducrIsfmSsUlh6mtz2IG3jIKlXEIlA
D/QjX3p0jP6XwHdVOHScliC4qdN9CgOBMUrMxy8TayU6BS+OAR8S4cHCPXsG
C1RPJnjpPI7N/D0FadflRUunflweH/+drgJKpm6RLwk/AkRC5b+Q+KmSW7Bh
pVwODMhauaD6Ddcy2qDW89xiRCRbvCNF5+1fv7sQtZ4PCjg3RAKGuPghPedw
9DyldpU2Sn4pJcBXcOFk4czECfLXAfEy51fV9WczPnBHBntNyvTmcnWe4M7f
UeJBj62UqDlof//JsWvjcIoVh2X3++XkacWsQC09fHL/dea7Dh1bM4ddnjCq
o9/BfIdQn5D2/mvsQtSb0++jqFzpF27VqUrLaoIjhV965EryhI8dm56ouzOA
hknvS0CFGa+4VKXScTIX+L7jRrIPVRHJnr/umJcl0ggzKKzI8QWbx821wu1k
bCKyy0PWlDH854gDEDVxGeTwHNFF8JGBPcBUoNLzca7v1aP4Ecim+jcYvZIf
0BtYObI/w4uyZ+nm2kgJBccamVGbtBV8clPQFNaymocdJGzpRF/BMtvJxo5H
9x+B1YU6Y7lrn+gUl1mI8gxoKglEETGZ7eLGWnLzq2FZT7qUtOe9eMBitEuo
AZ5o7yS3kmTNl/0P9pVQq1C8N0XlMMfL/CQzjm937Lx19oggmwUl9kg6qs7I
wJQpke8/HiAsYXUaMRUYCmVaw1knaWPJkY/pdJEH7l6fFyXcqSrQC3QfyTU0
39px6ntIRxjBEbVBJDK0f2YTEzbD4eFp6rE8OcEAm7qYXGgBH98PkioTlIWz
TebHZdH+nqxz9SBjU/u6z8EMj7NDDOxj6wW/CscDgCTp0BpbhxxrtT+zsYxd
KhszpoxcuU7xeLwVrCibjzg0t2nHxwz+twtBgR7Se4UumacZb4hzgwNswz3Z
kSQKmU6a/PzWjPbMu/YVaggb01QhoO2j/Cuo87fYlVp7KnaoBYQHzW/Sksgo
oaj0fXnEQVBwYQC+Zx27pDBDeO1acGo2XLBPiwz2Y1CyjP1y8eI9/Abx0A1w
JZp7K2/AJFxtQsn2creXzx62Hc4lsIhED8ew1brsf8Zrtmw6wQAYEnV0Nb83
k7I5l3bdlBm52vmEcVrGGIUzmptQv7GHP79aLh9ruEoucQcua5C1WSWfeR/o
YkyENLTdUlJJa9iAYKG1pOWwgBoqvNXLw+m7vxcmbrqim+E0++vaosIBw37g
HW+kl4bAi0NxnDRukOF+gvXPzFhfgu0vuqUY/wJ0uu5DDlFy5cjoUJYhK5wm
ZffztRnPa60tF0jtrKzXoF7Q13t5JbqeC8yPyyzcGjqKLhNdAM+/gXkDTAx1
7Ta76D80Dm7Dq0LcqYpFyv8Y31oXgEd6TJpFCf8tz6DJ7uxwcoom3bKQGKhN
xbxTCqAaxrxVmiJyskSCxyvv/AnsDCatlHMxtOj5KB/X5JXEawzQ1TNZ7HHY
V77k4jON3cyssDz/5+BReaFJMI/rSiCsQoNdPDjwglUeQI9P6T8f39/AQNNu
6InnEZmSq5sE1/71B4QnXUdvfxzayQNcUfAW2hvBDaC9J0vGEZw9688AU01S
EaM0TgUnI9pS8d63j735EuHioYAZ8qt2pLx61NY/SP3obeSDNneJ9R1i2rRV
b9Of5NOIbNJIZ64zELootpF7gtsCa/GNCmirciY/0yDAcFiZKEntkGbYR1y2
RkqMCdH2/HN6SmP2wUjuJc4KSo+7AqREXlcChwuVMz0b1hWca1g/JTPsQxDP
WuDJI7oj2kj2yYJG2J3U0SJ3Oxm0hasp0hj5Q29aHfVVAWHc2YC1AUso9IPj
oriph19ZnVPs1uqIKKIfSC+xUkprofMTvYw23e+TU3UdsOPTxWESoaWWZCmn
xySLcj8HAyiKI4QKFmLaWg7PpBWFZ4hsu9LrBM/y+0UUREsjDcnZuEKvr1gD
6xvpXSaZ2m0KvV8ehL0rbD0y0wxSYClm5BRBReuc9mXoPwOYHsRA6WVjgWl7
uUGRr6yyxmu2NUPqF4ck3rpUelcOooUUCqf7z1JdkALV35GCg/iCfMIgqJk1
/PPz7e6Cpw19K9gp1yJzrWMGJfoNvS0OK4MjYwBoCnI+QgNYlz9CqKbT7Vxk
F+wNeiO5AcV6O1ZPqJkmnlkpwG6kqQzZH1noSt07M+Kbz5QuIcpY5zoP3SM7
GC1GrEu5Aesm/sq0G64igFxGK0OJUZWiGoPmwuJKST3QVlnwWgsiDN7R7fMO
g5ZWH0Sc4hloRbNnTwufHRt/S+MsMk++ei8xcYJEqi4ivFTS9UOzM5pcSzpl
/yNHD46Ijd6SAp5D2aOz2DjqDKKgrN7k/5JHyYBI5X9IT/MG/rsQ0y4MgOYx
D94pYpI0xsSQFo7oB+4tOnJv/65+nVoxRiCmcVUFFT2L7pPpqIsC3Cl/K0g5
SQ0XHt6n+q3vE8jU/2TWwzzup2/q8QEiYi1CNynW6yUAvA01Z+R1NVPZQLxh
bYO5xQ1mvXtDyqwfhKxoZKsUEe8gwUAV4sGc9Uz+CIi19sonUei+1BqcnirV
o7Xu/SyC36lxit/XY5ztXzSXCTgaYJMr7fOq4SH8yuu8MCBvCeybNTwi/+6q
OXjAxzd+7PCcUAl/XY7SK9FZaEl9gLzqobiDmfXwAPPV+mh+oOMAJUnBdXLu
E7IHUEBaaxmbExmIQ1sa77Ni1x9GvAiCjSvj8u6uAsvYr/d9cjaJZEmGZW5r
pm/j1aJcyKni3/rIjDLwXXSPzPB3CgskQlfjV0QCH9faWT9F4/fSHuXrWngH
PZrXC0lBnHXwf8d2vmldK3PD6vQeKq8R6fWqKoHTE1ycf+IpJW4riiknMrdn
BTDYwVJ3GV2A8R+p5ezWqgWxgi+E+wD3mQyrWnCjmYFxzfqRR2OkucdSQ/9M
PunFGzV5g+mFULo1oOk+r2M80jZRBwVEN7ubDJJ8dpyas/BhuApzbOxM2fnz
TcdM0+ZPZIJpf9CPdZAa+XFBw6Erv9tpqXNLsJe30iPbJfDN3D7+PYDBXJB0
FMagz5tP5UiEd/HegMFot+OU1wTRX7TyrQm51O0FIYj8RU535Vl0MlW/a7KX
FLH6FoEhscveJ17VdjwkXP6C6dm+35soK/vQA4ZLvaHxSWrKY10AsA5CWtZS
yTXwwiYHFW6w3+RE53PxY9G1NyPjX7+fPvhZ45wqZS5afiNBUEEmAvx4VT2Y
0bBzgDRiWY/NK9lGc85s9frfBbFREcRRkE1pSwYLViKv1kozQo1bMEFbdAHD
Gen6SVnvjTt1SWpo3qUKCOgIzGux2POtbc6qBymP8dSIVt/bipKOkxKrNjkq
gIkXWI9SLLQcEe6XZK9MEdd04px8c8C77FGhzNmR1joE0fqYrAAchby/bygt
nHXnhWoGQUrhnObfq7TDgo0FLABWqt6WGk68ZvvCNdHn4TnbZ5i+QXSMvM4R
5ENhEKXDxQxFrSxO0N0xyPCnUSC/TsM5ag5vvdlJ0bvMRnG75npgvtXwqRhN
Vm3rFCG79K+ZsfAmgBSY3IbmF96+HA6Zm7lE9a2Ygtvyj5crMxMq/ZnM5vWD
Q5Ld7XLIpphD44fjnP/wAQddaBRUFnx5Pii4US41W5cR66GwoHHhWH9ojWFN
MJ81t7/SJpk5mygvedPhHApLvmMhwddbH0RaxJvXxKnLZlz9R4BThF8eM6RD
das26Vr31bqXDJCdLxZ3lb+jd191y7QWto69DI4aKf98YFmhHmt6bRMPmK/3
FQFjRz4HQk+1SyTBdi5djmKqmrGJG46OFkZfYaTzku8zfQDg/BOLMJbqSTmG
t+dP4KyEaym+3WTTSopcmdFs6onccvmdMCURwUMyXlzNAfLarvG/NUNmqTdt
nGiepikRMUiy1JlXCeqRiDMfgCJxgjetmwavpDeam8tDDbqlnP9sxOu/wlRz
TjmvMr9DtKNjndAKX4SNPKv0cVQmygZbFSIkps5ce1+yhOJTWRXDo5Te/37l
ljP36EV8bAyHbBra0wCt/IKtjm/ZTIbKLxy1DzXrD9UysM2O9yMcGOV0N+79
0wiToZ5sf4k6ZTZh//c9460v7F6hAXotlIhG/9K5lWzDcgV+M/wjxcn2yRso
9wHeDEvKvb7qfUq7h72lfH34Zqam4A1YAzAYM1wYQ4944xcaM5+ffh3HI6ex
A2KSAVHrLG55GCCvD3aEQrk5QooYcD3ZPt0As/31A3IKO/sBSZpmgakqI+NU
vlH6EXl7A5xY6feABR5s4H7p2saUnLKlBDO09snKS6CMV646dgqkEOufZ6wS
7AImfByuGeHSUH7ndNOeruzuHn70jwP1gi8zM9Qm6Q+vsihz1F4frOEnDTAm
pYISxTn8toKxlahrsRWSgLTOZ6kYyqpzbKj0PqkSYsza3MjXt1xFBNxX7w8g
O+xvjoPpCZ0sCoR9cH+hsVjIi8Rc5VR552/rT6urlTe3+tSMuHa9eZ301eco
j3lg3pMSJHQJ7Vv7X7aBLv7LQNQ2I1G11bDRIVJKs4YMk8r2CnW/Twn6Uc1M
5QBDtuVh2alNvAlQKk5XWYF8mOGA6Qzz4ydptgNnRS0v0gjI2wTYdjkdywgd
SPWaIyKTeheSIhrvcTEJk4z2CPhmnX8fM7BAD9GAMkvQaOoXg7QQUyDvjXSZ
BWscPoOzh7e0vlt4GJmYLh8RW6u80DNNuzwglxDjTraiwCyxmBba0JgZXQJb
pHnSyAx6vQjJCryUr0ZWlAn5VFjjkbhh74JeUYMgMXgwUIT8JzVhTGG+E2zs
Q98VP9GGm4kYjq+KpUGpLn4YazIvGucABxzQH/az03XzCLhtNC8c96nWfvv3
SrrMGXYhq0lI2F0nNBHetoXXSpYyt28fQKY2xLoyh2oRrXOHh0zdFBuAiC/u
FjdsuetLB8Jmo6EvhyL3ynp0S1/X78MmtQy3ilqmfh928o5kD4EFEannetnj
b0dLIhAP3OJz200UH4VKReWslW/Y+1eWdjxadFcF/SGYop2Tc6WBHzcrnujH
qOVT9cWeAo90ZDCbkGzUWyuUqNlNPJbMxKN2+S5oAIQ0Yf641KbVqJ2jCMq3
Hmm9hyNztzJW5n9SIniP7FY1WD5+AF7tjrLqhIg78yXxucWwqk2BeIo1wShB
6Ln9FU16mPGTTlZyv2Ob5wMgQuZDuBM3GD0WSGjXPNrk/Ob57QzLx0RsArpx
svgZLwdBgV2vvGUFxvRe5nKuLBG9AYDr0BD1+5zgxJAQCL/trP+a/HdZ6O//
9Oqq6wxouUPTdIvF90gGtK11rI4wfZlCWzOgMbPCj4wf78gqLOWc0coG2A1z
5UYkoj1ASlPWz9OWNBNSpFEhiSuPJu32eWqz/cLYHkMGHX3jRVqjsktrZ5dz
kVQrGev9/oyom+kkX/dmO6whZ3srq0Qmt2GLUnYHeM9hPFPISmncbEsWXhJE
uihwSaOERRnvB4IIjjogpl/mvbU0Hj+Wzp15DG28v0NppEKtHLiXG2W8TKja
YT/0OKghPXDOkjN5rmGgV19kTbwqsRwOWxcBoalKbu9nGxb8EpA5lTah8g58
zg8Z4A/mfMg7FxoTWSYxZ5HrVtEkGFrYDkotTj+kNP9F7BUc/hVsGCplVkwq
eLI21ucmH+Hzqe1AWplBrb2SI5R4d8bypr2XKV7dg0IVZ1b/Krr0wZvSN39c
z10fjyAj/LLnS9v/ahCl6ng5Rw/rz+gMODOa3CkcMd9KU0U6L0CooGf0sln5
CoTiQ/+SRlXnIqbbG327EL6sbdb1y5zj0HDIdob59o4E9nu5EpvQfKIBgonP
VVhi06XBb1HnHzue9Lp9kngqus5T1Jv/Q9HQkucjbe0AaB0WZcj3QRe2P1i2
puuoV94TgJi6KuuhqkYDOiNlSafi6NbatZe+gKhSZ2aPlVpW35rmskkeIYSk
8oETg8+CgKp3hciWD4wM57J4vH1N9NAn6PNeNzPhLsNraLpb4+S0irfMRjkS
dlSqlRA6vmYdgDhpeTjms7aeQu9xRJ9E0ZrhyX7gbXMRat+XkLMHZj2vATYM
GCDlVwJkEwJAH1obrtV/6owuBip71cZMgHj+HAY093t8vBdiv4nl+aQzKQk7
iXWkvzswDsKG4L4W0yURlKQH4nwcN7n0sDyLlt8X/UQjucf3Ei3hSEyiXlfC
gy5Rvebn7b+qEiLWOCRYKYALWTuOIApKeCh5ptPJfAY5x3Ncs1tyf0KtYZqe
MQfogMq8J7b0E3bh4cm8Q+ZJfXhUVXkU+L6WdkoU5pZPocgLI+MtGZMon79O
q2licpzG+lzk3UODWYl0BmlhAWyIxthP86zYvWUQI4RMsXiFy9Rww+Iv65rP
EdWZHRuApGqeqdbtJ1r+xRESmZkiEbDdG8fo4NtWsONK1LhozvCh+7OYeKF8
00zhXBis+c+BNQ9RGxVT+m4gHpGaWhdlpk+5Ip9GIQY75tzHc07XtEsbWVv4
Ti9P1/eZ0+IgRMyKKO+czN8tk0NxZlb65SFxZBrqd7jHejAh+KS6awLrLnqe
aP7gfjGHQWeb77jvCPTodF9JzGU+9H+isYiGADSK0zvs8nj4WIAwqCFZXBVH
6Nuip7AKadVQf/VZ/NDONOK9LHgCf/o1Ckqhe+d45q+w4dScNFwX48qu0MPa
tv9OFx+LZG/1no8pkELaaDbt0Wj9AJnqixYuVTU4oqfi7oLxM99qt9ixgZgg
hCni67ymjSiVyrbf0XBG6+SoTN/T5REazEGe6R5LsiqIEYI9AU4AE7MKpjPe
eKSuLk0KsaQfd7reBURQlNDawUu51ZFZHWGoh9UQyR3wuApfK4UghM4DgGtG
Lyw5I7WLymF497KrrUYBeEVUlsi8ymU/KbqHYUiDHEoNRIi6IGV/KOft+1RV
6z6rYSO80e4L1nZuMA3UJrWzZSTiz82d3BNIINhOMI75FpO5UMhkaVpZWjqC
IwBvMtFeApSPoozsteQx1YF3UPc2qdSSnlM6oauwNRSpNkRLJbGyLxOwUe1D
KZ3W/6Eaag+HGU/e7DZ66BFCN09IzW8JLnAdBqD01XLb01BuenWCKPIoB2Ed
h6m4SPTqhMubCdq0UofgZrGnt1MwoRMq7JCguN4+yEjaNpBvVjtDqjEes61g
r2vV8MPyxA04Sudlhjg+In8FW0xv85dV5RjgjtjLKvCZrVnS5uqaDqHeUzSe
XdxtlkgRYacdVq3ZTvyuieY1/9Pay5AeM1zgkdhki+T7v6gFuo2fDv2SPfT4
XtiY2kyPIeS8eOEGsMF50qoWBg+VH+prnUwvk78og2W6qiPLGpTLdIy7jgbC
2vS/E2JWVVn+LI9gpOGceOJvq4WYHjbADdqVa4/ww7CNnNxxBxEHIbstfk21
E0hhIWkkIV5toha0WH3ZGgPafktzjlOV4Lf6FREwH1JJVc6dRMJdtB6Bjdnz
SVZ0KhSPpKpWtimFgsqDu7mBtl8p/2LbrabGI31oTm80y4EYBBIo8r8s1In3
tX6O1X4EzLa35yyR0v46FcqdldXMsHoTBK/q6vPJYrNA6z0xn8Tl0nxxuWVZ
wg6OirW7vXBHJCBwj2ZKGAKgX4PiOD4DWlgEvYCtg5ObyvKt6Q+1Ui+gL9Sm
6dYckH8p3Wn4C5UZuuI9ot2IoC27rc6uVuvt1AGI0y37deh3ddna8GYYcWwQ
CJ9XpruFBkboEokxKHr4JIExH3g1aUb3xDbnDvjScK7XUbFog1gvmh/ZXh2D
nw+oeP7FjFL55ws6Ncywn9RH1ubHb1Skza3AORZFiFrwZ7GLQ6a2wE+BAgar
3aMgteHqulSeOCZqYhgbTQA32w6TrHc8ZL7HbS29J2FildVPthiRAsG4ebQR
H8LJdA9Zh6iiKQerxagjFMs8UVXYiYEQm1id57JFcM2gc/WhS8RaFf+QyTtw
l95c1M5Rsc5mV5KB29vJV0/cWSmHGT5C5+Tl5DGEFDp9mb6YtkaEDotBAwV6
32ul0hpywtjO8YXMH8DtnyrLXzcZCdNFVHaGhOo/PMzytZGEKgH+nPx3+jFi
/cG4KzeY/6YkN/8ux9/B89bXS5rOvh5tN9b0xrCxcds2vYjdlo2xyuGTgmJf
l8i25Pl5/yMnB61ofYItKsCECoFTLwU1jUdBDWb9LzwxpK/9dhIQow2Sfhzz
AO7Kq1H4bZp19c5lIkHCdcXublyzcuK5PgZQSEsb9CpkHxRJokKvs58H1hnZ
2MjApGuPGaJvXlSFuejwz84MtpTEDAWWohdyqJiwny+IeUFkLEtQARtu/Xue
NY8Vwq6doHcYbClmVaLviu/2F8yJTHO7GzyBe26GuZDqidNBZVbOGvNi6iTv
pqYz2H/FUX2HB9VwDRKAfmeCTb2M2BjDNKMZlYoJrQrU+506LWtqgUrCQKlh
wvjJ2wHCgvsN4JGlDLjCylNOY0zDv19dWgy/dw/0TM2tA6/pzPfZHlIUvSNU
MB8Hh4IFS3g/bn6h64ticZ6XLf4u9oJNB/GsCEzlTYfTb2S9x/D8qRZpVDxd
5N79VjGILV2bzFu4wQdnU4wf9L6RzinGs1BmgdteQgqUWxx1xBwpiOgSAZGD
SJ7cjf/V9UoLs/zN0mjXtobISZ/YY7UxKpsz77+mkhvziUsKqnOnFpj7zEAl
zNLmZMmGgeihhngf+HIhwixwuufllhKh18PKl/W16VRtispKl9c27KOqKstb
j0JAkzLfdoHaJFxtoY0sIZgTtgaJJ+6VN/zwMAdtbcGD29TVEpD9n1oa9D5p
r7zqwImQ2tQep8I3D78DZvdiHOIs/590HnuZQO2k+Gw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpeh8zprUeoIEkiUjxeksP9Rf1TRXq+o+bEXZN5rx9seqx7DzFdtnvl2LdRHtFTUXT94Y26D7957ZzYbxuH6thReHij/Cl+eYb0dcxJnPDY6uADpmqzP+2eeqWYwAXEAF1OJPpGw0l0Hwv3oayqMzqDVBUaFVxr8ImLTIn3Oplp2kOdCxUxOrjk1NllmfAf50UK2vUFbYnKpEZ5JbvuIvJgl36pEmoHYH+Pffm5Xkqd8uWPESjvszv6abgqINCq8kdoCQDWf57WO/Qo1QbKZQiQ8GY/E/VauaST2yjfZNbDoP5TnPPwp48LJv2bvBOrO/8ESFgzWJn94qIbwFWbJ6HIP/JBa7Un7RB9LAd88CyBkUXmbZJuHMo6t7B2Xzkkflduyc1bpWPhsMfcooE7788UEievemrLU6m/LKIdK1AukK6rj1xCQlamquIvpg0zXqtuPiICYiyTialWZ/89S6u+0qx33Uwy8sZfCiemfMB4M25pk+FHtlV+DcYLLW5+1VtmtRh8EOcVW2xX88hC54pkfSvgmo/NFBR6KM0e5bdGvvMrmsyDwLsPx8UAcvaF0NKODGxmTGfOmUhB2hvzWALt/zS2Na95mcbbX5shXmkyv4N6RUh/lviq32qxPtDDAebomoygqtdCDNKL/ZYtgfFjAuYw0jR0QrAgoP+t/t5RhYPo2NkaDZ4AzVDXPnrN9nBXEMB+jjLbpS+/YRNoz/qKwsatt6LZSEEdjDPq7RC3Uj5/e4UDF+6Lo3E48OtCahHUXqxk1oqPGWwU8QDhxbrPna"
`endif