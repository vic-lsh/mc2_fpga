// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CLGu1AHzg04KYF916rAetqUHH+8iTGwdAI+lmUkxMmQ2FOeTdVV4J8XQzJCp
KEkA2w3Z60B8lkMN+rI/u+fIoy75HnVl2kdWfFxS+gy3jVgVg9EdKtpjinUD
4bSXLyI/HiyQ5Zn/Bts4NhIMhMsGjSxxEqPfy5ToOiYN68Xuo1+V8FAwkgsv
ulaYOb7/eL5Mwgj/VLcg/dWYg78CkudaXn79eGM/DfCd5p1CsAyA6inaPWQw
heMcbcUosFffpCbUY5vlxVCQAY6/2jzrB7+tdHLbqjrxPi4AEm/R4w8tuoys
7OV4uXIH9O+2Tl9UlYn6EzUE9Iqm7wr/nHcWvPBHEQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fj4p4qqvHkZlt+DhgVcHxT3zkLDFh227TTLn13pnlf4n34A/OvJ27GlRgG4k
isJfvh0S3PZi2jAJLQiwdPxGEJS83dtqX5VnfmyUFzEw7YWn8+oYQBV62pdh
RH2rdhzvnYqDmjipx7BA4DXLmuZR2us89eY2U8ZfnxqH3CWaG4NPekraI1ai
CJ2y77PSw6d8UDju0v2WzyumT1nsTkK5TM3P+GWrSGSJruyNJVBNzP4KLZmF
82kNGGQD8sLBtD+/GiKMsLcI3+/qy8kTjsF7T/vq8vnPeEdALNPDJOu8juoD
CrZCDV0czsqTVai4vJ7IWwmD+Xv6ZeRm7zA5FplvjA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PVFjfLTsdLkie5DsE4XDgvcBAxm0r3k5fM6iO41UBXwSh4H2IGrznfJRkbVV
KxYg7Gth6AUlMYCQcU3MpDDNaAl62Pt1kL5z2QPviJB7f317BbIvdDOoy8LL
F4yf/61wZ9n9wjwr1UN0FTtQy7+ObD7stkTcz+x0RUmFp0WAPq8vs+N5DffK
aIcof6+b+2Fy2OsZoWeqjCqHcemUVr6Mb4h3MLwGYt1ENBvO5ebPVp9fkOCc
FNB4iYrreRV1BifuOr6lSphVrrl3mMRWaV9v/kMPqw/S0X2QeV9hrO+6JK9O
uYR+HVhZ78Tl8ukjueFhOuezQW/m6Chxk7BmOveI4w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eWBP9UpjUnAY+LLMmRsM0/frd4roaLdWFLoAxdcomSviXSWpsd2CUge/fB3O
3Hh2TtBTxqE4Av8Nip6oIStOXvcV5SMWBtpAZO+FQJ7HfW39vvpMkS292NSK
2mrV5+pC/wjdvCyn1rFTCHfpg7iBE6MNrV7eh+MtB6ua5PumoVfvJUHqPI51
QGLXWdCtt6U7UCgmhkIUVGpFKr/8gXxpFMA73CfRBUaHn3Q15tS1OUwq9G1P
/b3OAuEYW9+3/T5mhzpOolGPuPG4MyO8sw+bURvijKzD+w5Qts1sbEa6jlzK
e0yTbIVPDQRS4g0AASGGEmB2y82PJHhMLRMkA1pQzg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JL61wXneHkdq6p5e5PV8rKpFD17+5jZRaAVX06sLvKhUORwZ4Bq3cNdhIHOr
MbCFtIHS9EExh1BOh0J09AFsGyld5z2nkQMcBrTn7jJaodjlEIXNYaMrYmmy
0Ierx1IwOJJqV1mbzwXunJrL8LMHx6N9N4oG0iNbZRAUewv1zd4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Mk5//IB6LsMv3KRx9Li65AbMUxDhGH+s/jhp2CdQjAAWut4F0ZZJz0Y7mLH/
R+440bRZFJEqC6CZ08ma3oUhaHwzmDGb/KscHzdgvop+F9npn5BGgE7JHpE8
IfVkRDloj1j1/57X/OLNqYFDnp7Z9kGfQuHfiIfwzbBi3fY/KASRp3BZG8HR
eXWEDpEZkDd7pWYHSQZPKjhvsdLfHR1XbZkyC6FlEWV9sxVvwOSLnEHbVOFV
U3wU49fCvoAd4Tm+uNegeQsnDz9IYyhhX+ezMFlirOVtbtHK1l9VzTaKn0Vg
d7RWiUfC8vcMs7enqbBVQRijxwaOkoten/WMhGogIFBzjjQikqUV++FvBdsd
t6vr3t0Jn3doeWgZLYg2V3ACt7PxXQI3/ZwHhpVQ/bXYrG2TockdDSVgGcen
LZ/zzAa4lEohux8eriCEYnh7H/upmMze5TnpG/bAM8klHbjOV5vz4v2wBOoI
clJ/VLOQ4/rp2yECRTM/AboI/QLM40wy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OiXjp3r8xIMLXVuJ/nO7XGWg3SGAuD8JfQFK2DXr3yP/g+70n6TSbroiMfLE
Nd0Dnlk4sZneaYZlPfpzbGJR+9G2RQ/zoedDNIedzAnbnHQFPXEjx0HywGr0
foo4XDCmOw0ZFvUgrNgyWmO8HmhMxwB004YnCLsUd63ptQ1y66Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LDAby37qti60bt6UcGYePuKPqBLk+JTl5RiR+etQKYt6iff/4DFowBJ60V0S
dF0ddFViur37U6X4qT3tXN58FyLEKqubvScMm3HHCRhotEfk3frHOq1Ot3WE
C8lfwHCGHXmxYfJVF4UYbKSWejxlwILH8oAL/sPzzgaPgR/ezS4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3568)
`pragma protect data_block
HgJPqMm1GxMpZ5W3JmvrsIYDsRp8i9WQtsBO++bJ8lsHlH70cTYO+pGUFU6k
VtwwWit2o4g9HAxhqwoYY7iw92igJM6IZaTpGYJfeA5hFPK9KE7Ra7bAizKR
wW8n1WeSkwzu3Lo9wfspx37wfGY3+JfkpXez9MaiX1Y76gozaLQAMYf4e4v/
E1om7ch+H5jeXTVMZYtFtXBJufaCU040Z6s6/c5VglQVtyJ/9Wd0ecY5j9CB
srrgCLlUc0+dN45dAc6HLAoMLX9QeQIhn/yqG4dxip6wNWyHSZJFJPgc+gND
rlzCSQty9MTHgjgCqBZi/ka3D/nQR0226+yEc2n1NAJLuczlKp399IS6oPbx
12CgwJA7lUdyVwHIDpyNCVeguBIMGl9d1KqT8faTMqiH+rPN/kwlpNhSEDD0
g4qrh5fpridQMKOFj3fQlQql8lgWc/wFSu1Ligx7se04CTJJqhJ80UlBMwce
zCoIwOQMTiOna3qlLwGIDZK0HZ0EHoLviDCpPO97vmvGdEslcLu+YLWCME5h
ubL/J40DD4HHyVTumLDHiba+Z7fXmhLTKbXw2I+2L7rmf4KVbVBOX3p97F2v
D0KEbau0V4EL4UHkrw5yYGj8ckdJOVVWE33i/GWGab5JV0zKZXIlxa3N2LDa
rU4C+8K5ZIue0V++zbQooRYs4mg5xxI9zRXoL0XSRv3lFmkwtQLZpJd7RuVn
5GkShNeMzGVtBvqPNbYD8spScbRPfKBL7yy4RSGyfjddCYq6Wdqu0Q66bHJU
NNG6+UNkDbzZLkmPojpmcUD6I01+mCd2Q09Duk1nqWJQpJ9tjufYHh2INr66
bFhHMO6qwCcckFj5+pkAogmywBEioMhljctKeLuOFHQyaDSqG5q1wj60HBGk
KhelI+EaLzAwg1rifj72WxJ2MHYVlgb2/3l/VZ5VDwOMoVmihlWbHcXpE1a/
ZNw1IF21lgAoHLmx+4Y8+aiqrXHKub/Ol17AGKc3ehaktE44V8V4+lNQspIY
o7zaPVfWpCXd6GAfYvTUURWSbi9ngFTGk5CWWiD3kg4srom9gHeirpZnpPG7
77Wk+TUZZN5FpOkNZddVYnnmvTczsISQ+Ucft6E6YudKRdlrGgqVbDBy0FPD
ePhAo1EMIh1QLqI+OIQAg+a2bmA36yhnZi81UfYp2KDm4nmf+BBtbjkpsw3k
8iaAXKHTe1tysSGCK9Hp/6JL9/02ZDSg5oAGmb2khKLwgsDznofm0lSLq3fm
LtfyJtSN57oa6mEhIwfMB55z7+KkgBjyMMESvEHOT7P6yzTpLv9GXcntcHK1
NrsnctpuVXQ5fAlidYKJInoRpCd12x6EOcf0blzvCUKERbARCMu2iQn5H3bM
xVJqb5G/APYRdjcFG/UeCOG+nR+/Amwjx27A1EtHSDCELXwZXF77NAeklZcF
0sYVrxucat1urKd6s90J6M4+LB2HWM6o6kvjwTEW8ufswwmjedUsrbz+NLDn
Dyq63Ga/DKUXFkm5Afpj7Pany3nWhf9JKOaonridNHpM3VnacqWRW/SneiD+
+RVrUfXqHwMpW+pt5/Q+RPOitgmGxlo97LAq/1TPg5TmpEu6T9ohRnInFnQx
3voJdWKuGdvJv+nvS5jF3gorYjdfA8DpSmVTsM/L96Xxjdzz8YV8dOPOyILI
MxUvnJoBX5j+V0eN+JU//ApGjCKvAV3q9KqbzUysZA3gKbruJZHDVJcVAdT8
CLYGiituHeUFl2oDIC83abPmS4I8m3EPYkNLc0UD1PzQ18ogcuTYlv3yRWjG
MQ+906p1TqLBbRk6LVv0OqasZem9rRvUs7Zcj1ST94Exrt+ufA/ukuPw68eE
y7qOBD3VbwZmI1ZIGyztxNaEXpJs0iwucXRlZo/WXFSXUaI9InXz4UcgRNhX
vi/VV3JOph7+8DqssJoLhdFRDTDXaR+oGQ0DSIo3cHGRNGcDoF6n1VuG/fTr
Uxv2jYpV9F7OTKSegSW2tccXGwJWA//l1MJnAnfwxWDn4f2INc9wJW6AdedS
ddu6Mb3l+aXIUHGrafZ9xIoHRIoVM/01Mz5njMpUv7LeQjqoglWv+aAReUyT
dIx4kYYMrih1hfsF/9qxbYWX1dttZDOVEfTpcODtFMwP3tA3OAmvdhJPT2LR
idOCq8o3bqKgs3oaEn1r0bO7JDnkUzM/F2mPInxpitEdc/gZzpqvUxuijQgz
fHqr2XzuLxCaKvEAZ/iUTzcuN1VblbMLdX4i8+XHOPPVtSxPg6me6B/HLiMB
FIAePbZZcgEU9Nd1VoImZC4JlW1PDCLJZ8/MmxcdKste5q8TafYGDHcbyF+c
b7+p3NMRLmCpqyv4cr/Xs+6DUmSTKFKN3GsCLl9TuAbsEn2FpEswJGR/mzov
Sp5qvhz6jPU1KnRc6VKuFrJZXrcTXweDPvDNuVOWKvAZaxlUjD8+Whwqs5X9
l9uYtDJliZPKW2zGlWxZn68gz3dNEZ2R4yAzZ2ygTfOz1+YQ5o2RPlxQL+Qm
xdktvI+U+zemZbUPVUPMIAqd4+aiek+4JeXhI2/INk67C8rQAqw0q6Vh6xZZ
tSR7vvscPXJMqmBMepNOwNSleQlLKHCS7mUZ55DqfseOk2eARGXpoUEc8m66
LxnOt+mEr1meFk3ZKjAEyMYD3Jmsd0Qq2734smBqs/9luDdyJhQCLUWvnKMP
nFpf6Q4cIMWIiBRy9chHg2JlZwhzM5V9HXNBGvYEmwUkhyegaE3aUrKIqTDJ
a35LneJ1Y4dknzq89lHS8OtXAJciC/JLnRkP7BpdbD5mGPTuU8AH5y4++bAT
NV9Q4t7cPNjcQYtkLI17krqqHLPk2xMIvLErgGiU1xYFboWCQJmQv0WLt/P8
hSw4Dy1Qr35a/YkG3HhVmZppyn7qA3Ivo6/VBnezFx45vcJnRIIE4jHsxm1/
Wg955hkTrqPHoSQfvZLOLjkOh11FofBASEkBx8NU2NAm2WUUoZ46l+IXaNGT
uuN2yLD/MQrUuurxqEN03j41WvWT0vm7QGvECVcU0hBHYstil6ahF8Nzl+2W
mO9NBZ6n4KSjShb88Vntfr4eWXl4A/bBDSn2Y0QvnQzZ0s32zy2NP4BBJh3U
GhQC4+1DuYYoLWxedpTozngMbvraimkunARpqPbMY0QvalANaal6xflXFfYX
O74k5zJdV7SXXJFutYWHgcoHIr9Q8CFQFH0+OnDquHD4CD+4Q3OIIxAwV9H7
jUYd42syV3SnliKCef3Y0iuWXZTzFdp3dwlHnycNdDpmfFF4EpK7k3PEIMgg
ygK65vvr2EBimu27Vd+hMOZyXB5w8QjlVz/2t9SkMsRMaah92O/2W7R8ix1G
+njqxnmQqT1W9EaoK6gNMc3Fwl7ToDyHR7pYxCd0DPiXZy8btGUabqJtjzS7
S5BRlRoCa+Nm2je4SNIcxe9kQ4oesXlHm9ZsCOr0FjrwiGOe6Cjfghf8EIzW
wpDC7M1ihYM2QS8Jg1yoiuobThmgGNSCBtY++joIgTaIljRjCUZ7ch1VqO7+
gXs8kKEGnOZrHxDkk46QDTz0UPM2ml6LkIApQMq028vvHDJYJUl5XcAbWvMJ
/Em/alFmeBDRApNKD/WqhT5hQdmKiVSWRb8WS72eYs+DWIDJbHhHwdvuqljA
iZxuUTueLcA0LkkIxQTMBMYT+oFCYGgvyVgke3HNpWKzPJp4/ZwV6yejpx7O
ygmI5zjWq2YgY1ZkxLk8ds/w4fptXiSKyBzMvjwqLBEeejEWZAdSog2ywf2+
3dEmB1vzHbCJwznAaP7fMIyJ7FLe/7yTOzzijrm3/YcnRioU3BPTS/Bi+ULR
dyD8Dc2fDhbNQoL7RFN0jVLSFLjj4eA9yKjMTne3gJS/PPf8lrFrzWW7gKLL
aWB50Wp+wcAOqh82047O38p2si2TyggKb8GA6hrU/mkGDZ2YoAAUIbVRt5Ug
Zq66fhshwTvmEHLDNQS9oCgO9u1++FN6jSWfurRZ363Xp522C0D6Q06rLCMr
PJkry7QBgMuPEriw/cbAA2pAb8gZTsZXR8BvNye4qk8jLDD/bx95yzaX9sBG
hJVBSbk19P4/cLpIAvXr6HqhVbKAxGrOmgHYxhb5DAZLpSW9vIhpZBXB+wDI
qBL+O3A7Qc57EcAhv6WilMILP2cHEq76TCH9TEssYKtprgYrOIlee/mnRNcX
85+OBIOByVGdJv73EdH75d0A/nbDtFvmv3gCeuyuD/dM5jPET4m5EtHsHXqz
rgNeHRgnteL7Nwui3uepDeAcFykEuRlTF1sbihruqzdKid/O1YiG2j7JKlb7
Kd/2aZdW0E/nv9i92XBlJN9WRpFXxcJUoxNO/E4a/AsX9cfzl62HQ2RrAG0t
5sDZJu6wNugHdZl6zHN3fYtbVcUqqYezN8as3Zr3Jkd+ULgDM+0buZ6Kj0IA
w6hBwqAiB8TZowpdJcMDPKdToPHJHnSo/GbffiE9h2DWus5KTPUZBhNKPPXl
6XjH6J9nN7hPE0PlTl+FEKHi4l6R+dP+eRPfWd7hKSX0JGjS5t5GAYhV7OkV
nm04jcUIskJvGTDlgxPuMmE5M/qi1GCiQP+pKhch1hDt5IjbkBOzYCnlKVlW
XolL/+2l08pJxjoVcJNv8eGa40RZAmovZaJ/L6V3Al5XCFnd0uxndb6IbmNG
JxTO52fvRFn6SQJ/hfxHxILwqBNK8vqDaMcQcbc0PWW+4WzEXLhBMbw/PXax
e1FXhtcvbjCj3yr2kg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "221cqLfSQtZLwpVKjUxAj0azxWo9qWyTHel1yyBq9riDaTa7pjyEaEdGOLLz3wcrK5rHulca0g1g9Zlx/VJp3su79bVOdFJFOSZrof0/9wf6C4nAWrw+2PgJSzMMKpaFLO6gpDFruW5083aTh1M+Q5KnW16yLzHWGhpxtWHi5x5kzslfPRMwe4HyZUYh8/FwJanr1Um2jvkSaUjUKvojtHUTdbUpkWg93bqHvMIamsnZk3Y9g0YV+azZRNakOoKbSmrGAgDyEC5OMW/lUfOEVdI7GlIaomO2phjNVLJ7zmdXnDKPPFqJtj3wchI1p1Z4HHZ9/xBtTbfGXLs5rxKg2f5uStCxRtVh4sZxY0CTM/h2QPalPppMhZR3f0ZezRz0EJQwnsiDYf/8kDNDi4Va2scKC+RxmY9DXx0K3Oii9OoJ11M0pTF59gM2S6isa/skQi8aTjiaMWR4FTT0nztbEYIUdDOXut/rjWi76ip/9Bt8Ge3LsaKuQiuwawiIU2/wDfkKC92j0JeBKu9JmFpMwM52xrPTUr+HwV+Kmm/VUxvGty+PVvFW0MGubbgwGVyz3hNpqWAQSFtZFriOdU9rvmJROQwH6jHLXXjgVbBFu0N0owJs0FZGuPBE6qlgFwFOO0ndxP6vIj7DOfW0HyU+pYbl7LJs98Qjaxb+LHgxbTWHA56+cernXD1ulmeHojipGhSvWXyEp3efE0aAe1J47DQNzAfun5fHcsE72Hw2glpjGyImflBZCVTHtQ3Ruppzxh2LKGUESa7KTFwxngnUjAF8xkk8DKQNnWcGltZIedeekK0Y6t7dzuaOaXsZPKazl9pJsNXjuQHuXYmEPp17Scj77088/IMh3LilzRmUPG0J7d3HgIx9DdWhUzyfR7E7t8gWMP4Vj/Y+tttum+OQ1gV366K3DrI2KWU+oTeBUaXoiY88Ubt9MyD50YolNibfBFrip08larAGq2RZ33jvAmrdsuUWqJpGqJCCeLVnRTH6/n7vfFDc0kb2TJBZPNOv"
`endif