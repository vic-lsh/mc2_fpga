// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c21dru6DZRheRsa7OZirJeOYvE9jQIwx7qsgtqXUCzwBT3jn5mC2nzHgRe3M
N2yoUEgCQoDN7Z85OI4hnaAxav3IZjVzPENaxxAr6FPqODEOv49heg2EpDgA
CxIdi3Q593ZmY1Jb/Jz4iHSASOimQ0M1XOO91xb+fT23hvthXK+Ycz0oiGBK
ZIhBjg56Q4VbbM6LivvAWdPKfkkV7tCmu21mXSb0kRSbtpcehx6KvodyOU6U
9B094bTMXMcx3xyWhrQr8c7wZiI6ekl9xOJXl2IJZoz9N0GfmcPQfopUlM7w
KKYC8akky1nThbaCvotH6DIJGatJIsAeX4y7batnsg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
krdD69aXG09+CQ1DcWwXbUonhEfCJ1oEpHtcIQmop33DhXlqN0YjohWSfvg/
GvJip1m1X0z+G5TI7QWtwPvSozmK+r9nkU8Qlpwp45lvGJ7i8XHRyO4cLxDD
NX87A91KHHaEN9Kz6VNf51KlZCOsgVEzutdbn5/JvmT2+Q7mhSShcsbNDP46
7ZKa9/GerkG6aNm0rfBx2JCSovI+bpUfULFfgNAdO4/ZhBOKzHO04z/LE3JI
8zFMxo/tgrf0vNtQySuEaugzvo16F1I3gdyMChzLBM87ZioDje6g6aX6HNBd
Pv72IhJAKHrG8CpBd6kCRZIK/Hs/w5a3MGfwYVsa3g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZysvoB0C6O09xUcHwRxVHlsVtxVHwrn/jjPmJx/gkf9aXHawlt8/6ctBAVub
r4YOlUHdAUBZJMMVaxw8hXkvgxjRHh7bUKN5spj+evclEhf4p1uClH3SfyqY
qcDmFQ75nslahmrPGnEB9dAhebOYb02OeMrSzxn8jy3jzTE6GRst5UxI7/6G
eEllBsezBEoOScd9A1KO17+rX0EcmwE34IQx4CRnh7lgZULJvAcf4yCvP4DY
ddt50ONU20DJv5fELRvv3o7Uq6GFy0QzflSIgD0WB/Dx5oXQPYmjhTDPdr6S
etuiTu3k9/sFPrK3SZdxrgY7+nmu4Abxf85SWICc9g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q333uCfQzUuGMRUvJj0kTrWgd35DUc7DcdLLd3wEHEKfODZ+sSpb82I76AC9
68h4zpMxg7r/3tdb8ZR9LY8k6eDu1UsR2gI9ig6XLu+bsPt9EgFcQEw5jDjg
t86dkFlLAZFXGt98pJnE1wMEs7diJbUz/fz0ldtgErq0iw4qkQGU1wzSi4O6
kOKpcCycfwAamdNElxOHb2hx0H596bZmoEfmWB48niGM3aD/78TvSNc3zFBn
fGCsp0JkaVTllHIhRHGLNdwD8zCaVKf0ZY5IsKg9ssS2gbazM3DZfaXPgOrw
vidFrtp67YyAbL2sWKf+XUbyLC2sxg28e+Gz22jM3A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LsiB1jIWvzxcTjiftbjn4cb+dGbS9jxrBnDp9PPBHsQltEDr4dpIW7L7Byxa
EYvDPr49BS0lJQv9iqEIloeeUbkoB0AEHWJVb+ZtfmVg3ZgSesDj617hfPGX
wzzC1xda766G/xDNdL+3awpODH8X3EoW+F5HpKbxNpYng3ZRQXM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uACU6wOER047/cTWuJK8Qoka1MimBvX+r6YxtULDzFAlpnVXa9DxI+OFOkNK
H5bQpHpXOMlcfrc1NJh6QkcbE6dbfTqSuIqcetToJlbuk6gKwEnv4c0zCTpK
ykHeDMXtfTXlbtsGaSH0p+KtDL6fD7GOFjKkhq+XTJMp9Vmqufkis39ETzzW
bUpfA5KzPPnxfkigUd0UtFWt+JazkyychecAKOHpJ1rIZTVb0Zde++yDRkx9
pfqVlW8w1Qyw9WesGkNA00l2fUAFqQKCjslP/gauHHTm3nzIj8r+cLuvExsj
tL41qpCAXPSQF7znVl/5R+BLFwmwp73NEc8wCGbZsN5Yl+kSp2ZbWawG3Enh
e9s0brNDRLyVjGFVNrd+Whax0qAvjXFPt6VYYWGyRW6wB6SRSm9a9NAhpVln
WHpBZGOOd+QRjsn3JX8Gae+4ZLDKAfBeK22CmmBPJanCfwojB7YDF3/vL7jd
4KuiYr/lr3d5WTMRKiCFEwNU7WWs97id


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EZmHTSrL9Q9FqXx6NhHGbwfnwqWeNvx5zNWGmEtjiwPUakQ3KJl9HxaL0DGP
Yu0gEGpui8h1tBCo88intMLKDJxjVyzm0cC6YiKyO2erKrq2RkdSEKsqFxa9
QCyY6WM3rnnwiSoZX/An1EuPzZ0HJTip4azc5zvPwQ/6FmR4jPc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
unm0OOfz3tWZFiE9t0yTV/byTfVR4B0QoX4LYLw8+IVJhwgDJbcVf76rUS/r
2VQ8eKNN5dcKt5DkmKlM0AK2zSY/hG+U32QPcDQaBkRt8XQ15q+ozXNoXRyA
0LaS9JZc3ERBC7HEnHfKeYx7d5u7V31vQ6czueY4rqqMGL0zmj4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 151984)
`pragma protect data_block
isBusjFDsQSHD3i7L5lJL2OHN/Vhoc3R7gQofmqDf7KZun9zAdVZYQz6lrhJ
9myX8WkrSwGdPIEPZr7KvRTzhlcP8gpMqxl2AXqY3t13eGgI3lfxMlP79pHT
Bt5/+hSev/EbiGSsu+SWbKu+1iT0cIoiV7uYhgR/mS8LthErNWkSMzsQS7us
fCh3wF3GgtkcNsQUXA8P/H4BNO9YHjuXZe72PDbU2EGyS3Xi8VGSvOa6KX65
lSjRofwQWHaikiTfBBvPyiBU64p3An+JDWLBz3P+OTdIrHSoRQCaB44o8QS+
bVOezlVJsIWvI3F/yHXR+g0dYfrkIcYArvcFK5Nzbx7rLyi2OoPe75e22QTq
8sU8eNcyturt6b5qmGSa+BDUlJfbNYO0lHWkGQlueVkAiQmcE6PY0rgisWDh
Vic2NsTdDq5DCuIzhu1bO1CiGRfcQrHH8Pd1YSqYOztiv9XwbvRmBQtuiwx0
AinFltXDyGxdnU1ZiIPJp6+Lh+3oPJXZVLAzabmq4WmSFlhbYIfE4aRli7He
ZIZHmT0n1zJ3Z0DY9QltaMZvbUmkXYjR1mV0yrfa+KJx7IGz7IYhITNoJXyJ
R/cnShvbhNqJYCi1ZutfObeGtUyeilH9bxx2BCz8htS6fGPu2YxQo+UxmQZU
KVcL2cDHfV5hWWR1GLQl2TT1D0+fR1vAsjeFKUMcXCGjVwmGinudcvKtLm61
6eStNMfDiZpIAV5n163DOOopnwCKNH2caVDc10e1JrtZQpy0GoU9krNiIZBV
UOIyjyXHGRjWkNwVqT6h6qmIfZCuKq8xWkHifpim83BY/M2oCYwruYzUHS9m
mnXo0aQFfWynRviNq+1jjpl6l0R0/I3cAHaVOof9H+u3hx6poIGvao1slRE9
1s2vBJeKMus/Tt64e3/D03su23x/My45C3F+NihzOsWIzaAh0fXwYXNvB8B+
0Zx+w7FCsf6YjPJ9cuRCv5kW48Uv8pCOh/avUUs1UEKQmUYEy1oQnbQGtaDd
VE9iaY/iKad+PtxJC5cWOPlRKcoTA7u10GboFu75l6+o+/zN38gWL/upTFLB
aYWhCeBO0i47k3qMe8rtpa0XndhzqJVzLXo7zSoxrR3e6gVPfwYPpTnXnWQB
M4JBYSdqfmqqrk/q/8BB6zY/rmAlhJbVkzVYGdwOo2lcQoh5IXNdfvJVrVsZ
74d9Ul1PithZkOUIX/38OgwnUpjLnccSFhSpDzdGAMnVOtSRo4b6SWSP3Eu+
aaWyKaU5zpOrrcwwMJLLIkwDj1hXMMMZr+zjFiyixNjEzcEhIMKqz9lAKFV8
WGPRfVyxY4ldvSjCJvi5AdxR6V0XRcgD4E2wAih9Wqjd3x8DI/oO1Ji+qYdG
f3C+HUdeImc5ds4kwtEib0UzQleteMHM+sH7lOcJD2cR+CEt+PmD/nqxYd+p
iSUnMAR/1JOpNLDY10tgUDRnM+1FwDMXI2nEqjeU2aGmRvE3vlrKiUDTcgP+
Fp8j/DXFD2R+kCPDwUenP0viLL4FW827bv+ZxthhN+742QtK7NtEI/M3he4m
f/cm5djdiWr0y8SjHm5mvevNX9a7d8bdHyZyamtUIa4S2uKMHjTnCMxq1XpX
cqcoLtJ/wH2VpI7HgJl8BcC74w7EXV8cQ457MNpX6hv/nbADz6tY2knacY5m
Y2au8dQZesmITINIrHEA/z7vnBw3IQM7H+bNApq9jTf8fmUFFwm7mBkmrPYf
PGySl22QRi1Cv0cQrsGgw70lh4lEd1stfqojnNGGQpmlSDKiGcji/zLTlzDj
jc17xyx2RityR/ddcbIWojxU0wQM/DpnHv6jpLA/MJw9/nu3xcTLnC37IqGj
cutfH4L0ORuZNaE0RdfiTLAQ4YB44l9Es+mTLUekrzaxBqnQEhzoEVtEuT7q
2ourjirfyk7dCUmnzuRBI36/KX3pDjCjRyLVJeMjhZLBtDTVeL85QBBzhR7L
5HhhtCDeMxEHYHKE+q56TLh7QnItN0T8KcMqAaywrLi1TTKUC/dmxmNPmW1s
auZbcTY8BLk1wmQKwkfTLmItcDNmjfDNhBDFz2ikB45qtVL7skFkXNCRAzUc
g6+BltCm07NTRvvXGJPhsdDnSKanjDwTQBiMYFDY2T0iiSB4vFZRxVAQV1dd
q2A2hIodjMgg71SvURBkhYdNMfJ3oqdkJHP5rHqCWxph152oQlD/CViGu/Ir
InMKAjG56PJPHgWk+ukc79hQSsccoATxm7q6R+ZxAtSeKcaDY9LLTGL0CMxt
Rd2bBI31/Bdl4ZeGIkI7T1tuPmhNAlU/Y2DpcEruW053sVVZgpL5C39QB9c+
eg2b8E9Wh+Mh5WLXgg83GWA7NOePRHJPcxhC5Ki2PUSbQsjKl/NynzwUDAcl
0TGUFzt5x2W6J2IG25sQ13nRfbw8HnO0evjU1x+W1qdcaRCA7vyYaqgnlOpb
hN4sZ15qATiN6idXDQPCgRes8zG+1DD0aZUP57ZrtHXZXS36ylHaYHwsCfzY
OAjyElaAOoYLFfhQmz6AFy45C6XBUqY1JFvkeih/HVG0vAbcVgHRoe/HPOHS
nWU9EyvQ8ernRuOF0lL1evpu/PvFpBSXMO74VsEws8Hk8pr/f1E0IBbruYy/
Rh2ddqyCT0Ov1nMTjg6JobtnVGZvSjbPFsmFhelnChUCSdL89aCA0NN/zlWY
XcWGT3vCAHtYqXwA9BcpmTyTKwc1pFWxOAsRKN1Yk7+nLt6KLFziIyf1YYk8
Rak/2obqY1MIiFe+yVxY+d3sq2rXBhmLyO9VMiSODl3LhiO1DfmMz/eCiJus
VJBNtbST0m1vkJNWyTj709DWUXKAXoMqgo/3b8lewESEY6lqSexpX0GpbZ3T
1AHW+6VkZ4ntuCbCKOlFWspJ3utCujD9S2vwOUVVTVMQCvWxGrdISrRpAAkR
9son6bp0RlSrzSp44X/V+Kx2tsBLNSrQjfeHaqUqwA0B6OuPYU+MoVSwYnjh
6MG3+1NZ1uipYYbO9aMxK9asmEgsBPP0Pt2R9bxNW3S630JXVqYlwUst0F7R
wCYVp4K1zkCTCMf7gXmu3Z3yRDL3XI65Yw1VXNRdgPIKXAOq/oaTdnJfaFIN
hmu+hU+ViXpgAWANnz0++R5yecr0yTMQRXnBoKwtTp61jr1hJmMpyyh/fng4
11yKGZ93Vjp7hH1LyO63NZoqWUdCkOmajdvWBsHqtZBs4VhRQHyOmOxvPy9o
Smbj8oFLAmUXFUjKhSudVbmwMGKoOFuX4zVk8vceJ+Yn2jllVXlX8dzF+icj
ygEZxoM0AtbWufSjPjPUt0L1QbgBWPYRlusWvcVW40EQ/OsYc5YQTFVOMWz5
2+qEcGXHXjg8acQdbmvV5gBam17xGV29DMLe8CT1vyvx+gwIYvH3gnBSZLcz
zRt+ejqA0H3H8U/nT1gav9+5ponSroqMMZsVfG8CqmdWSUydmo9WvwRGcgD7
CJHESf5APQTFfSdIGu/ZWWphLT03YvNiK3l+jA8/PqO1Q0yIyFIMf7OWgEdw
aww7Qqc3MBcPAsTXAtlDF0tX2rdCNkScTDowi6sq+nIX8Ym0c7bF1rdiJEba
AJ9l6q+uvC918AmTSt1Sle7UKCroNKL7DV7gVpQxfsK2AYiVXTN6CgQby+vr
zFuB4IrhAkLXfa3V1w4BBtHPFoWrTGZ+M4gbivLHVPJ982pwn9+JRXEescWG
khSVAy14y7mERT65AOtWBPiv8vbDBwKB2TTIPoc8sJYGCQ1r2cV/iCQHzYwU
IWYDJqxCRPAi3pQRjk7+oymIHEv6ckEj6Fvmtr0G8vf1opeadaOQV17Rmk7E
/kjKYjVQKDPTRi7lqnR6HeU+spCAuVBR/bvZdUj9hdecdiReGHo9xf7QBEF/
Q+RVVtpOckhB2UFFqrSwnE+8df8AQSNcsKpzZt5Too4/ut6G928GuQIfh1St
m59/SHZPvNNVtGdJMXcUWz31J+7TlJuu9Q2N8oEkHw0Owad6K6pt0aX/Wby5
/rFGfDPcvOUoLlQR+cTovLWAAocszRNfIDPncFkqa1xgcMswAg9SHNVv87qK
lQYjiw86IJg4mLiGFTDArBqiwu/dq/yEkVjJ2bl603NfegyE+bh+cAa/A2+d
C7Icai1vPdfejXhBq3fE7nAYjzexQ2y+U9wu3lNxY3NE/fkZyR54kWFQ2HVm
BVM7tVWlY0BMWb2hmm/F9n3AnfcV4rbYxucyjCV47i59uO0LOIplW1lCwhaY
n1PJv44H75kVSqPZ9Ky+j0zJj13xKo19sMnhFF5Ge3wScYHZLmwhjMD/wu/D
PGPDqGEWPlX2McTJ8l99bfX0TCEQGu2M4+FRycf4LHjSd5rmIRN/UHkCNq11
bm8M2FVflZ4aRZRyIP6/9H1jz+t8N1zlu/NBLZzhWNdKy49RdaZTIHwSF75x
SEBr6A2PUg35tLuix4x6Q+sobOY6lrHnAqcTwI2IyvkpvLyV7tBfYhHkPLiZ
VyszAH5d4ZQJQ+xiCgEbB/APBZZFCoBtUUMut5lswX/u8oEsd5vCgX1H9eos
SwKOww/1Ru9TzmJgKZM8Xi7qwa3UQ6NspBvwkxoPn8TnB3ZA7xIZmZ8Y8GSz
g0fEXb9HlgRpeV+ZJQYWAlZ2M2HJFJwc65MWA0e+eQk79DiyXpdTOnGhW6bm
MskEMBcAU2QZjlPN55JrO8eyWOAwWPF1xxB6vFqWxeIpIOQ2CjPyLzEf7Tuo
bj6aymmg+IqU3FZkvNiO+2qnVz/c3BAc+qgJls2Ax8RVaEpYdfjY4TMJTizy
wCvFkj1wvBSI5B8fdIZ5YyunUGMs/6LVpJnRRV1Ky+dMorkykkQYHlAyXsJc
7fKd1vzJZgxuEFqL8AK05+ULNayMI+0J/SAnPoIHiVzyOGaoeCqfUf09i8Qa
s73mZTCtX9En73gBJdZMASYs34bkpyRR0LtUsWAql46nzdzGgG4VB33BhwZg
LVB9h+U04pMN1XI8RANWQEicVj5Ptj8kcsoZDATIiv8wAaccjdZ1f56zEyG0
Ce88+CAfDElhwidr3YZtARaL/gdrLR1t3bMcfoZz8CmZPlvjDOESvGY9sy0Q
JfplQM+/LD0vhBhjyu9UFds8Zm5iwbFhYCiValpZcXxn27bocnLINYjteuk0
KBOgUbII6T3PNKbWHGwuzBDMskaztwC7z1kfq9oab2aUyoXZaDhi9/+uwe+G
WS26saEhTYClV8W30ru49GzSDtOn4LFjf1JWdVuMRvSdm0toOX1jwuaTUpJ2
mQZMfrwwHQuqSscb3eh7dXYA8mV96Ot2TlKtqPQJWQLcSUUVf1ZFxR1/3F1L
g53THRu6JXesh2uKRn3PW5OwlKn8tedotwMoIyXOeYVCqBawPLIZlPPuupSh
EhmwfO1dlNlJsB0E8kG1Bq7b4MwtdyjU5Jzfu1Sfj61QjG0q3wqc3PYYXdEX
1VS4fkviMvy8L/NVBHrJmP9IdZND5WsIFaGj+4yYbbOHGpHiuG99vtTvXJTm
8mpSydwOL+8v8R1auFQ80dQ99Fd1gm5bRoVxNKObRFoxOHnxpCrfPqh4Vev4
S0ZfIbLPDlGtTQxyWAo7LEtTPByiFG7HCRQ80xyOohUctM+lRsv/GzIYRT8+
hRwYKqPMpdEUOhyxk+un5nyEs8OuMjUcZ+x3qyMuxm1eyTK8LYlaoV7BV6AL
uL4SDo/9u0AOlObgQ3kMfK0qfWGZNvi+Yv/hUYJ+GZasbMENU8CINov5m+ZZ
IJ6Ow6EbC1fhbHjuvTDVr1HjkwoLwczAxZcs9VyRsrmxNUM7gHQTgbfA1ipU
ng1Idky2DcqExkumm9+WxqPw6Bba0Dn4gzpz9FK5RSqOzlASOXp2c42dnKHR
MxL7rrOHbDq/gZEpEmCnr1q5fuAifztWm7zLE3V8WQzJVT54HUtdVseBp55s
lb+cf5XGgmr2bFAuOwzu95LZnd2AIEKtyP8auNH7KiGGFgC4AtwBcY1cQ0Wr
ISBkIs3boAKExJIdSNOuR3Xcuw43+mkIeNr+bgk4mFzBZY9P1o0iWJERgIKL
TQC8hNiJDzDikTrjpBGk52feBaRwkUHbtgEV52RdmtQTuZ7N88fjFLzjpacu
SKJ21tPFaF6TCmtaytZSc8KXRWOL2CN9gfIItF44gr1PcHJGQDZxyIrabS3G
2d/eFXwwXZp0XalSKHcOCLropLxdiuSZDAwVbIUsG5d18Jw2vplkpvOykl7H
ojhQ82a6LIIcGXrhytiANuFSiU1gDUnmXHXXQn2FB0J/FskaCw8O4hHI2KSG
K2oeyVxwrlyC0Naah+YAIePjv/iAyfcW8cIxwC08ItP9TPV4ZJuqsZYsTq3E
ReO2nfpjN9oLIvwT+OsPInKfmYhLYBkg1nTQfVCZ3ZWFrfopIbeDPU6SZso3
fu6LJW4c2/sgIzZnqT0hk1ezesKumO9ab8iPwPn+l8U9jDP0UwWeTuWi6DT/
ilLV3Ln5WzKCNZzKxGtT0KCTDm+KQYOC3GHCHGN0fhbG4r4bKuj9CYtRI7/C
trKiFuLKScrdETTIPwaE6287uqKFf5s88D2aos38C7T9N3HcHc6dpN4qmORf
2MUZxdZiH7lKiAIck/+mExWvxCC1ly4XXd+MWNXD3L2y2NAvqWY8QIEIRLaZ
5ju2U4MPfnHw6mHNqmF1ixjpskTInABp2wT3phCvi1Jr8w5AzCy2OwL0cgW+
VLYGgLAQwwJk4lmymp19Ha8tyTsF4PgxJ46SkBm3kEcMVxp2g+Jy5NdxsW6C
pTlmUieUcgQwwmNVSYkQX7Y75JRtj5ldnB8Y65SK14fnR5weK0elggGU3toX
8hcgY1jrrceX7CC+wwD17y8cfrxXRVjbw1oVQhU2ajsimdrtBO92yzshZ2Um
7HLSDipr9YuC5TreXEibouhn2l4MP+KvBwMVhrIVInVN/f/CwDUNrdMujeP6
TO2EUkL6p9Z5p8YQ/86gb3K17V1n158ObyGtz1FOcxo3Bs6dhy4Edxleti09
ckecnzgturNFq8DRQ/XNj1hdAp3900I0Yp4ReV8dLB3+dA7g/rOrEE+/+tL1
bfwOaXDLbAdiRiR3mV6Jr7RtarHk7AnHCyXbeSJt0c6QWEuIhxPwatJj6pf4
7aq58AaTgve7+DfmQH+r1iR7fvyVlKbJHNvihzhGf3YMgnbrIhRJtzWYAXbz
52AHRQetuuq/tglWv/bINHebIhnawopXa+qgDjguilofCnP1Gimd0ghu8wFR
3GZ75IlkOt3CzodMPB7J3ipJEHS3vahA2AV8H4OqNpq1quq2BVVA59yx+X8R
s6DNzzLgt0baxZiQrbTPrzDESBuftmbCPmNH111RoFVaxAnscF963Q8FTbza
zqsG9iWP+SxoyaVW6vINGUoBHqzG3JoigQd5k9NY9lb0IDVTn80m2hiixO1K
VZn4GFXP+zWkdKQDHLT+v31S4Gr2z5FZ9fupQZgMB3mW+br6I8BFCqPAC3TM
R+9HL4tSkYPWDm1xchLS7gChhZexkmowvzuyurbz1TY4KK/ZIU0xl6GFBkz7
Yihnai+mIDtOQhwS6vClmFrABYjbt9ocwaWlONCI13Pqx11jCx8TXsdVR4QA
FtTRKCeHOG5eEC7GUpSClM6dkcDTe1GVtImYgpjzHo5ydk6h+FEYKGcvkgpx
atdzrEuCPwrlJALXHbY1C6/J5q0Mw/rybZbAC8plguRZXRc4C+AtV2Wim/Iz
AFEAjl1KTTV7oSFas9DKr66nX6KaCtnDytaadeZnAdkmHfvvFufyBCwcz86c
DwS+n2wqfiJNlLOmrLfBcqLu4DEdJEK5dGt4r8rXkwd9W7o55vrW5rRSY5m/
UsIqJClAk+yX5bLdUYxKpMUxrEO0CEyQmQNvF17NPfJzccDHDE2QrKWfLsQ7
xZ+Xyyj6vSTSS06giCCetA/jqabrG7BLJCnpHehNmHKpGLZ5APkoeRJr1vsr
b9YK/RGQx1Qled1KSu8Ohzm4bNZvUog9Yo6YcXXSdHidZSC3vwpyUv3H1j5V
iJY13CvyOSBWZxlnTWv8/b1hcbFHkvS8UWGWC1l5sQSJYG69/lgEVtDMje4U
NVjAEvjGPJRbt72dKvGTfUA/zvFMCxBiUtJLaNrbhuMA0nQnMaikNDMi4YzI
DA8oispZJYSIt9RCZ8ZLXxqYM7pSDGQZkGf+KHFAii8DS0d5GzAFoiLWYhXo
+Thuf0kL2oOjL37omsZeAaE/gCjOznSeL1iwld5AVP/f5UjyQcsOHvwYRzKA
bn0vCRO3Ar/qmwz+ONowaf3T+kouX45QaoJsmdGy00BQFduU5Z1Q/tVGThW5
L3dI7mlnKA7Vi+xZfZEk3bxiOhP+L8eaZ9kR3ve5ZAKZEEKOEymK0VwPpMUy
vBRE2hznWkKZ/4O9GNXYDLYFcHFkhBkPw829TBwG2aSroFyEpB3dtbiQFPFJ
JD2KHERW1p1JtnkXVv3yRdiEHjcU1PJpr4BgEHVlasLsr2QI0aJdv0dNMlv/
xp/7k4qMh6WOBUb9zf12MsqtZgnpKF9eKXPEJs9Fp23Kxut0jTwDyuBZX5vQ
gJ331DTHXlAaa4UtI6+XqXf3JJMRBAWrydnXHU3pVhhYcOMDd0TYS37iZ9tD
mNTJW5/VT7uKMxhPB2oRq15wL0nIzMBtPF9zxp/p6h4DrzdOT969wGsdeveo
co8PxJkQfBuV8AO+3udi4P6fI8zpMc0xKmrXq2CRIYGWVgkqhVCMQ2Wnefi/
X2AEEdM+kTsV99/mnKJNPY7IpvL2Wqw2KltJi1/erG6DwWcxk5qRueSyuiI5
LMCp84M5xTce94CY6fOHLsMwN8NjwDHuZ9jWwOgHVz0SImMH1Q90rMejsWwh
Y+nyNNSWL8k31PKO6nigiBQqMuOrEiJWYo1iZ95FaALlaMnLWeI8vYuvYYtI
5NjdYCzd6H6u+laQZtNuMO1drVfZVsJoHd6BL4+LKX6/ZrptpKunRrWDUD43
R2+XlCwkkdM2LarPWzux4SVZwuHSpMzHVJrWkpW0inv/IB9TtF6xzsjC9FVT
1qd/7O4NthgSfTsmDdrkNxpiZ8IarrSV+ymb8gzIC/TzfTRUsR5uz/M15l3f
H+vhHX3kXlFB9S2QttZoK//AvIMrRQIPKg8GgRqhXbvEF2yb9Pn80JOpB5QB
dgwj1ostuAAkopa5O4XwPnQcwgMnF2n2krgkZR0VQf+R3jB7MqJUmc1Lm7s1
O+scxFYNXBgXLm/pZqUgp5RRzy88DvPQYDAz+JBamC26PHGwF3mNcsEtVhgN
cmbJW+MCfYysqnase1yWnpa8bqyw11NzBpicMeW7UsRISN8KmLpn6hUXUsa9
XtY/kR2187d+MVYZZt67k28or8O+UIqEANkeHwkt7jsnQT0QV4yAv9Zunv1d
Z5GE2CwVle/v6FT2zRBvqZyQdHEFxgR48siPnci/hvF9GVTqVNGMbpxnnuFw
5s4tUgRo4ye8w2GhGwtTorrMMnOsZolRZtdmNllUd304Vgab4ZRttQN5B/Lb
/M2cfCG2NCY1zoHcblkYvkCIYL9IXmG+2SGR4u2sZZ3y7PhCgejyyB3zjkFH
voyYNUaXSgyR2Ux6BJQx7jJSdKOtaCQgNFafUtVacILRsye21DS3wUNPG2yF
+8Tko/OQdoT3eFZclVhCVK5HwmpSnIi52AoC9Ho7T7ol2DqDQE+8RwedGlRU
w8ycZCQaTt5vufu5LF/g7wdUF1Am27VqWi790pP7WwjJlf18jTB5e1vApLin
hirz8b3d6dSiQNsLOnxZitFJgecmWEuf43RDwi9fR0ih6ZJ/K38HgKSKn8s3
zXrNF4o3xIeHXJihdcyQmdwyXvJzLmC98Mf0z2f03mkCk66PUFFhi2vbMT/z
qak7Q8koxJCtKKv1VaNCZHqlbQh5b2NPjrHa5Oc6twzeMQ1iLrkRiokg4fHu
/tZ7wx9Z7v4RVn/ITp1TvgPb6lUkiN/ItxHYjn7nT/IxkNRmOgyWcs9rIJ7N
xnVYngVjaR5jg/sBlUAg12gyX701EhNg9P/tTbkq+7/8ChnQjVRMlxvZgjTG
sOKuEaJh/aIX2+OD69h4CTn63X4BNn553IeKknKrG/ZRp1D1aozsntZ6IoJx
a820PqtpM5R9FJsM8G0GWZudtPI4ti8m2z6BJcq1RvdkXxYEOsbGzHgZqFQL
QvSn2/858JIFe/FdDPuFsbEl848pEMruK6dBjlZGFiuJPmxpxxayUDykATLY
n/ad/F1fa50rWfeuOOFrI6InhIusYhz/3/YM25XWi6nU9Bt/5SN4m382xjFn
3ruXN5MKjlnGHIQogKABJF4wp1y2lmBlCXKOx3/UrvlwD/T0jhuarH8ktL6o
L94zmULB7KY0Tezns+dpfDQvEG4LLsB7CHCJp6eKdqDiicdZ3QySo/kPQZxz
G2+B2Tozhvkz6C1zKItRLmjkshrWzQZM940TfLkU1mR+o/HChdGxdrFvwQPh
i9wWjrfmaerRo/Qf6G42SlV9Lyw8TGGu0zZA/GlLZX5YUW2ycCZBkjmaEVFE
itF1ppD0bHoaq9q31Z1E2rN+l3TvUywk0nGUGGjJqH6s97CDv1sNjGeF0z3s
cFI+HDOkCGm4ngGUX002nVbJFvR1jz2VHDWokUN9RtOG6YmZALT28zBaRnlP
lhdV0L6GLUGAUOQK58qEvdeyMWJdrYG7dFEuIcV2OszfsvjCD4nfjH8OsaY3
1Ji3egWv0i59ecDB3QOhICjWE4qsZQAt5oS165FgxImfcwlUNSSEnBtCR1Pr
ldHUODNYmKKFZWZcViEkhT5oKgVs0T8gFDhmdps2UaJYUhTKForOZz19k+Z+
O5hvvX7UUw4OqhQ+1d8huY32F98DEAPWMpKOQ8v23xDfb1rahT6O/f70rhGR
g+8YSwvG5REuNGYSe2oAxbRckpGip29APkCOV5LK8NRL5lVsoPpQEdWIgC08
p//mLUHL7Jr/OBOj1NJ8F6vRjHXhv9Mc1Rpz6JFimGfwehFQs9Wc17ysd/h2
etfUQUpQijFt5WbSY9JCwuOEf/ZpgPxUs/gr/vhJjsdYVElFyiWVWjoqyORZ
b7KYTP4UIb+4YGAcWHarH41BqXhcGr1d0xBE7Tw3hwIvziHx4T9iSSfDUw7K
mlOMWrKozipoEF90TKXaVK94iZBJrll9/YfdNvpMLr/16I6vI7D5J2QE/bbn
ekscbLhvUJ+v6sd0a+qjBKWLGRvVyuups48iI3yYfTsMSkFBsw77/DS1ZBrN
NbuX+EkfLOpKTZkNQzNbsp+JT8pWEhNNoOpiRAoGkxKSnOk7UmUToRE4ZeTr
Vozz5+nwZUnJAXWHx5e2LKAS4NhIUQ2uhhjaZ06PQ/a8BhQB0d6VvZtfYFqH
DjssO4Q3huUnxGFUL/c3qfTMPIQo/ofGHolFSzGhKoTfuUZlYkIXp7cvruzi
8oqbAHwlGTX9DR3IbqlunILlWZVFL4/6yY13rSbOKyFkAfm3BYtlPN2bt5mh
4jbMJn94CQ69DBycYABHd1K3UYg4llNiIWBu4wLodLDQ3r6Tbw/NTbr9DDnN
y5gODiLChgyZgH6il1dXBuj47UUj25G302yzyjOjT8gbr/V0Ds6gSIOtdcc/
qrScSNzaUaiKHg58S3r1BcUPP8L3rDG9kd2eNtOnPhLq2WVKQIIJo0OG81Xu
XNGVFRHmdPgEQ4jAFEPzEVDSVllwaOhwrOSo5ThmAPmvkWf+LrJjbvDGHIzU
c5OaLUdPOU9p+Ukx04HBDBZOREeT3qpC2bMbk5vP9pVGBzIP8HhuTSDPGiyt
rq/hwD/KBfnmJfWnuKbVdxXWvZVnPbgGLMGZbzS8ghh+OqaOW60+TcGhwmPd
d+EX4JRwaC/Dj4K2KX0CwwB/aOmFV7nDbTalQbSE69Ib7RcypJtgQ1Y+jPEa
3+4VPtVl5QTretPzntPUY82vTIaH79AB47k8Yx/q2ZK6k6Fl01esWl6PMCk4
vpW/dN8GUKeKTErQrMx/NE3tmjzoQqx0Z1RjAhBv8zMCxe/Uu7XVAwBuFUXn
Jko38TRf+GHr979xJGoGJQjf5F7zMHMG/+EqjtUdhF1Ax9uxIu8RuHafv+3R
Ytbkpf4SLJOVuyP4U5d+MHfqS+zF+UiChcUh6N8vHXqSP1rm5twlmCjcfb9T
+EhXBPScRtwUGBkdSxUtsXf7JQHDpexUUKkB4rWKGeyMPzzeVd+hVvYrjlGB
a8Q/jxfVZKI5TdBP6W/rHeNbSzqy2OjFIRdKljwObYomqBovMRVPOfmWO9bT
A8dFbazZL5WAkZf49X/bFONiQfvqW/PcwQVfnM/JVakf5aVa/bOilfCMQwK0
vsF01Scx23AIVtvvNsH9/TDq5b+PFabETjkirmLRyjON2Y/l+UpISk23ZWnd
zLA43zbSXtQQQWbWl2pVA6+5VbnVYKC01TglwHSYqJEOBUVlqZ2aWQP0I6ml
P7adddX615J2sGSE5z07lD3IUybXP0q5/z7tXJqYPdMK0AbJHUrDn4bVlA5c
hMOC0FZ8DIqTt3AbYfnW91yBvmPhvo0DjoBoQIoQ5nqaqVKWf2F54zH/S/yH
w42vOVoHm4bffNubqMLxj8DKPITPxfdP7PnzvkpfiPrOe7dkgsro2bEu4qIS
sFf4DKo5b55GUWvWtesLt5JpBbz+lKET6eQPThI8yT/9fN/6Eh0GhLn/0uNf
Z7nUcZqlC5RgnLxUtiGTBFcTB2srrSPXvcdr63Lq4ta2tJwo7mdTbXAXVhNV
8k2LhqMGsn/f0O+yISWdH4c/d0TDZfodoBzRdk/Pbi9uIeOizatNlivVq8kq
8fhVAk0tl9uqOnyahPyuM5/Dthf/coQY7mL6hsJ68VB7BqZFo0cKNxwV3jrA
erbBqHLbnZHlkmQVanZepKfwkN8AVGHa3JoP/7ja8g8cI4SW6rgN5N1fmVGZ
ceMzAHYfFPmQiPKvYvTEnjV+qSyggnRY4STOVvTsZeUBe7QZWZc/rDtko3f1
s6m/8Eb6s/fyggRVOxKJngeY3GpYxzBg60ZaUCG2bamSHdCColOdq9/6DOLQ
R9TS0ze8MJNDLJyR05J8kYD5X72mOBHeZ3lOeFxSHTYVEg5Yeif3VFa1JI12
sRntWcSiwFcXajokAtweLeGKGh1FGtkqdXmtCt5FUsW2ABf9AtMUh5dTx+3B
TFh2Zshiv1ynS1tXCV46PW2qx8MFE9U5MqdqAYejZ7bHYDExJ+Y8sAWo+3Hg
hK/qnS6W03utqENLY1jJzP9Ko1gNDdHA+DzBCafWFqYdiXxHT9TDONxcfaGE
flJkD8tKjQW5dNPsRbMIRquvG/Y5z5ZEgLWrGx6Up9/aPlINUgx1q6lf2OX/
kyE6mWPDJeNe2rvH0JicPC9afzlL5JNYF7bgCKoLS4FB4snS+nnfY4YFeVqx
PPdo5ln9Kt/RT55Xn4YHE81JmPy4W2pch7HoIYMxoeHhFIeODlQq4fBeRLnI
WknIbdsozo09foH+NVcQAHdDAxBJGLW+PEZNx73Oq04ROwhC+PZa9fQwPhvi
HDWxPOieSXypMMQetWB11P5k/SrsO9gE2ODwsmTzZ8uo+z+00Ml7/nD+S86o
JRMDpUFks5vxXXYFkM6jkfUa9/f4FyQmFo9Wn+i1JOq+Ko0Uqaoudeij3dRu
mE55JaMlIFPqh7m6A2WH+hOiYmSsakRdJMpDB4sxnvRv0KnZqs7yYrpb+N1z
7c4Y5mH6SrVKpnYRMGzp4yh2Fdfj9nGbhuGRWUkk050rv+eXhiaDbdjn8msH
BqFAV/N+ZTUttJSO7XC17Ox0td18e7OM+5yPc2GO7jDcjwWodoOgyA/PT8AP
yjTkgQi0qFxJzQAXu5ZLAqIiMR/y6eY4f4w/q+jj8NFA7VlPGpaerF/Z2n1Q
SDHgBFwoFYLu/9K2k+7/1eLTG8MfTrj507/xUjl9ZZND7a4nX3ye3aHnrKr+
oIM1CxMaAo2hSSFzFvRVzzzRvarjb688BDehiXgY2B3ZlZjtpXAHkc5PgUWa
krqUCuSxTz+/xnEhOo4MbE3LfEJZ1GqUG4BBjs3xE1o8TeyzizYhrs6uJrIm
swL8lDaEwruCHP4gMKZoCTxhMqoOQTCikT/XsTJklAlThuVoOkCKQr8uCmal
zPjUjTmJDDICr4U4zrpNM2yopuBRUXfoKgmwqarfeyvhSGALRiI5RXelgrk5
YXwLhPKwPI8Df+XUio+Al2lbQbdUNoJfWyAGY+ixegqB+/N/OhxnlTcm170S
7ezEjJpwAjkrj6hi32X8E+UyBRvE3av1/J2P1LrAs2P4oLlVb0ezropxzoVx
wt8Ap4Iv+920pY915DuOAxdZcFVFyF2rJVG+wpiUByvMOEr1mD8uXWO4uxtX
rA4quqWicTUEvbwIkxRPsAVlZQ8x3Gqv36U+aInb24Yk2P0awkW0iKy+EXFS
RVidDGNxkenpp61GRJo11zdQ2YPYgJ6E1Cqq1fuFFKyPDkSRn5hJ2EkPIDcQ
0bV1mfVWHrTxJJYAWfv0A8DFU8JafNX9Cvce9ilDM6/YwPaqB4/578RVD6KA
Yr3zHz7PMME+9JmF26OX2EpCuwWRHelr1idswR+KCNcVkrKUuzu74U/sfCmf
3Bg+/2fpaQd37CdeDaC7116INjtHT1AJ/wmN1bsYThGZ/XGn59M0PK9AApd6
L+6akFlh82YV8KhbayFDo/dlMW1Pc6r8ldlIz9yrwwKMGxK04KOhDcMWEVCn
LVY1GYqXnrUPWpUVXs1bYICYcJZ5zoeKobbGeL/NiPCZwDn5dJSotkOyX/k9
thA2nACFzk0+bolJAXQp9RZV3Z2eIbeRqrhxZaq0QiI9TxbGHm5q/9axE3Sd
7D1KWuWPJgGdWBzcp15T+UlLFgIQ0/qdtfY+fI/UVCLyGjG99kBGpRGLmPBh
VfaIBLQ+xk6iX09y/OBPjPrXvweAwHt/cEvppJiLF5jplA0lX0HQiPYxASEG
akJ3zFL+wKGm4/jys2T6ZYOI3ewa1n+uQ6E1lBDFyVWclx9uyjBFeKqNboxO
a05LOTnTyboKOnwN5C0mUQTyrEjvmJBP+NpwT30cXyRVyMUaPVK9FTlOS5m5
ZU8h+GaXq0LC6phYw+7UejDRd0cWcielXcRdtU4aTtzQ2dpjbXdKhJ2fqs8X
ulecQcnaFzdYnbUNUib7Cl//xvoYvmPDbSSUIQEZ57eeA5SVve5Pyc8PWLrZ
ZKf0WgECVOkkEHd48wcYykHyX18JaGcu1XKivRAVFoaX6e76tP0kZ2M5ZQ9E
wGjw69p22GVWXiY/haYwn3ix9UTJj60ooQXIgMLNrj4G9bXF4WUDE8QJRc8t
gd7o3ks4Ha0ci8N5N+aPy+hfUKwKET63qQ5QfFpLqTRmSpqorcxvdsTIAKab
7DSoLvHNUF+W3ohretyY6BG4iskE39kidS5IB6RakQnamlMSv8V6Oabo9N8m
ygtuO7Jz56iP+JYX9TQDzDbpXsIms8pJlGlvxgfQjqpE1sd+sQYVgW9SwDFZ
CS7fr0Xy9itMV7V5radW/Of0rRO7QSin8YF0FKERgc2JiShbkcj6SDs3BFwu
J45+WdJarX+OEabdaJJNHocINGz0wtyZEficJKFVqY9DxM19zmPBi8qCcZK1
VCBWrERAUoxtLldo0qHtruEjM0aPG8eE/oL2DFr6LiLeIOwuGQXxcrA2jWPT
sa5zNEnBfTsD5fScreEN3C7tcmUuw+ID3DbvoyrjUCAm/0uDhD/l9JQpRmu5
4mCuLFdLx8tT9Uwhu06wng6YABUtbo31MIJFWvXPSyBfchugE03l/WY2T/qf
y9nF0a3pjoggt4zStxk03Q1ES6JqexAe1z2RkN+DfOd4POnVR6Cli3OAe1RZ
kwZyWAC7Gp4ouSPnmdy2jF7JnQoyqVSEqquse6tb1Pe7WWCg54l4/X+1wGxj
3N1YtTnNkVkEDbOg14B++EweDAHKS75NMcnYA7pApDLb4MqQzSYwO/vEiUMY
xPpFNWtwGyGqgEakAW2k81wdShEyKxTjRVyKP6T+zF5LORQP3cEZCI96+AB/
mMWTSwsnQ1Hp9IcnEpDliZ6R1ToX8aK8NUhqxUCX7h6pfPyIBGSPayFuWC9I
kNqwfG0OF4V/KWXT5t10fhQ1fTrWah2uvGmzsRnNCNH18tEVV2sezu0KcrrF
0bw54B/YpZ/uxgI6NlDVPZ++ZI6y5B5GkrwuJGW/wMbkW/7bIRMq/cIMMmhW
lB9iHaB8WD/6D5+PpbWsXHfN8mvR+ma8eUGFC4CgCvyCaXWFjKIredLkykyg
WC2luoSyQvOZQYULOa1vpmJGRc9NIKfmq5VVgTO0aJKUWy4JYvnqaxKxrGMC
6D1QUanrnkdJuYK6+uNilk5GPdzO7gcEhxUvd5+79qoIEDx8YybO061PYxCc
okc3NwN5wEd8aIA+A8L29rRpHIaF98W+d4MxSuC1ZlAVrceNH+5tS1GTIhwm
RtjBsykQD1NUWEg5Nu9WMAPKYQK3ouv2R/4qWVESjLA+Wt/izq6PSjOlCp4O
ZQSS58fMG90sDCWHpKeNTwNQpTMeimzc1oMGzk4YACFUEuF6Ko6h+4Mx+Fp5
k0/ZDdM3S2o8GodSSbBkUNiWv/RUeU9Wqhf3PmPVJbsAYJbCcrVqWZ+nOngV
/NHmK7tm+ItUt6xm8VRaeoiLph8WT3O76sw9ZXaGDhTT5ATtatarwPXkylLQ
6ehONsEAuayCh/38raCJUaGc8Ue1MvCfGyBVMUI+pin/Ya22qJDYpzNJsDQY
a2UQtGDABpguHHdGn+W94FpWiJotDvXuJWIrS2Cfn/EuM85bAQju9hiAiBPT
a2VCj1cMDDz4z12ldFw3ekVogjVhimIwOH9mIIfzlmeomtJLCY7QDRXKrpL2
njPLfrC366ZXQf+ilAFxCKzmg7DOwHG0FEOqFJDT7mkrJ0jxrFQ7PHGK/KaS
ssgC3GIJzij2pkwD5WoDd9YiEuZ6KIzX0MDPNGf1dI75a4XKeu/+4l2ytACh
zgBjw+x5AHEg48tlOIFjlQ+XQVRnEHCMeQ4rghkwBF6A/Bm7+Zq628HzfVs8
EiN5IPeuTlZ0yPt1ZUlHDf3SXjYhk4RoTdVT9kGirJeVb2TUPOdvBtkRsl6S
PiEILU23uw1wtab1pUZzZGfCLOfeU6ElBJrtXbl4OKPHSYIvKpKKmZMgtX3W
TI35gQWsKgSec9QXviyy5b114RZT7+d8lffUaq/Pjl/W0bnAr4RBrtA0nDB4
m40M9AWzqkKLRbnb7tqxGJQ7jWsyXbxx4DQDhJmLOCS1Oew6jok8pHrO4mS/
Jpcih1no6GQDY2o0GE6Mg++WnbXCsTr2Ks72qiMYMxRdxdYAkEJ3bcPNvqbo
IpN7jPDhmce12Q98Y5f4/pLK4npc+xewvJWdNQbKpOC8lx/uzX4TA/Zkig8v
+nuG9KPUSSfik3iKK4l7NmEiHFEmM4+m4hMApVXcC80PjWHyy+yAnLPLecnI
d/IbaAgEKLXt8Y4/O9t24dLKrksgu/Aruiup6dFg3lrrACd6y6JHkJ0T/3A8
KVp2tvKtoyAV1WLaU91I/peiQp/pvAjHkMfzRSwP2D6Gm468vj4K3UgkIFD9
q2LHKpXLNIkxi03AAUO2Npe5OU7eRT/WBjqsPcLaJGmvNJaIal0Dbn061igj
GohVqb0RrDcjziJcNlVpw16pRDU/QogPRbLEAftL/UNhpkVzY/Qh25zI/nKv
3CiN7ns23z00OzYlEpUDG96gx6faILeAtqEEcgi3ZN2TY2z09o/r6tu8z321
7KfQKrwyJGKYJw6CbENeN/Oi1svYOkooe7dcWw82paT1OVb05KCt89OQRyaL
0XpeQqnwCcg/xiD5yK+3LJtIeqQ+wS4eFHoVE3Dfv/0+jeUYQnCq6klpjCM4
1ciAVwYL8lwZfqgatlMER2Y5vXxaa/iYwXs/aJWKJOuQInBwNYVWTihjIHLJ
2kCksD/axbiyfI7/1Q3HPNLpFEnvqn9QblXUUfqsVskB3jvPwRZbmV1gxd4v
9w8D6iYUDEmcAwV+zyCv0sBae4UslU047PWr+c/pUJbfO5rLuDoX3niFJZVI
+exFwighunKC++ayaZ08+4C5udoNWi1UbYabHzNSLSWJ+FlmiXJjYvHPbFsq
baIPG49Mw3iYiPwN8vr/MhEgARg/C4L9P6UdTJ3555ttw/6MzEF2vV2u3BRo
BCfuPzEk0L44YnB7b5hYHMyV2rCTQdapf1x1l8nR3+DE+EV1DHtItIAzF/qa
fU4KHbQc89Tf27aWHEN+v2vd7sKNQfZoC1Y0n4U9vMvm2hzUrh0mKZALz08N
opU6Rci8JGDLzmRIF4f4Ybl+GOgiVmAShTeL28kCf9I971aJwixGQhw9A0N3
b+7fVaIhmRq2OLtUW9ohqnpCwWFK/uKdpQNeLkIDqU0ONBBsGrhfYAWxAeVp
PYOyl4CO5Oz8QdyYCJ9bbWepMKFbhTDm0/cvsh8i2bMmQfm/5HIwwWt3uupm
uCUI9FulG9SkE6MCGy+1xb+RHn6si2wEknrzWgSqvjGkzRUBlUM+yrbxMWZv
r7MDPm/mjlLiMyyJogfYxW+uUcl4Bb0TT3dHSzF7OXu9AlVJk9iG5nj06TaN
n2TVdpQ7U/20AD+a2MnBRndaMEOQOKXzWzNlvGDqkFk/+Gi0mHQHg2eUo4f1
gIaP5H8U1wQFKpX4nt1DuujXSWBPAYMxWcdMYDJbv4Qda9KFmqVv72CLAeHr
3/jeu1/tz1VwPWLZ0MDGVk+ok0DcrPwsVvwNLPmqrLC6W81kTvJQOaMJkY61
8skG9xlJS/xNE+kL8XzIubHkZ4dCDz/OdKWJdFK0FZU3g4HUVzXobJEisx6o
Tfh3xrWT/IhTYI+0Tsb2IjmynBSsFsKoSy/ve1Co6H7aqrg9gWAeypr9ZG+g
0tFKjrdtrl3S+UGnf2QfcYupAq4Jo2LCaiGAk+8KHftPgW56SBzmSQsuGeBU
3KUOZLRiNeQPAn8Zu31DdhC8oGNGxaJT+TLnwOPZ2Kr9xqL0JTVHMHQEXmxA
bqUmTFHtMDq6ecR7aIhV06tj3LiwNXAp50ljkudUUHbwcPGAaHJQ7skh6ZQP
yWBn7OOUQqlDJL0pZCfkyP5xUHs5C0R8Kf5No1HIpwMLoYrpXEMsd8vGHPSf
NI9+Cx8nAoS2Ja+I8JFmkEzO471D9LC2PcHPLD4qFjLp2Nzxg1gc1Fokaqzb
2vckuU2Z5eDVqK+WLRKjeISsmip0TjuQvCM2vjsH02b0ry9lk7CR5DbeTFj5
eK9hPXsEToYsxJBewbNileCKz5VFj3hopwU216O3jfvBYAUY5F8uQNZwdzcA
4sYJ7J/NqlFFoVP1qxu15vg32gZ+cQQyUvE6Wbf4ZZvFK9DGDDflP2+VZWi6
9jzr4F3YXDUSkOLE/BgQpptku4g0Wd4ayEuv+eX+VRmsV89F3qr7zJc5IFRI
b0ArlF9Rsh1opK4OcTjURVS9nq/612rMpGMm9xWlLBNbS14Z5vVBN1jmJ40C
w5zwGyJxv1kU4qdbn0UbhKfOwnWyeqCPPTqV/69jYbQJJxIxubUn+JEjIEbl
KSe2BB5p0jA62iFQlDTSxe8Fuqs4qfw7V7Do6SZq9/pML4TKcEycYanj9egl
C9jxxGmjbeijWeatVEJLO+xowD4EVqP5wSnT3OZvNifc0/pbxpTAzZYYJAFZ
oJAmaD9UcHdeZcTySBg1dL9V09jbzGLbGbKB2q2hEIgYFxpqIiCUn4lByd8h
XGOf9KlNtT2Rbk6LOdzcqm7/eZH1MCk7nG2uh0V5cRlTq1ZYKwxdlSnNo0VG
Srkyg6aewJk6bHfKvO+lQBP7GpbSHEPZbJiD132M4cocwZDQqTLUULEBie63
CWaqDX0pjMuTxmz4UKLQrG2KRvhFSGQKGksxjA8eJOu3yXGDmPfcVSD+9f91
QEuNYIdXT94VBZk5KlSD4+JoAq/WbvuWr4Y4b6oQjvxJSbkF++SG/fbbb/R9
vBruCV82w9Q70y9TtsYaJwbAPi55K49tO0ufLXEsLkcxaatEvUF71rSx/6+g
3nSR80vsrn/Lizj+aW+egA7OibyJlfjGQN91LWBqAkbN28YA5R3dQxhNg2PH
WCcdiGii7uDfgmMqC0hvGBXwUYgBCfpbd4UEK4HBah1lpHJgVI3tpKr9cwpq
G6Hl18GD2r0JdsYa5X5kkj4tIE7Jx9qsESaYKAssR21V1hfkpPytU2mTOtfy
WXz2kZ9YNHbR8By30sh1IlTXN1SEkeCe1gKocig0KCilxHlEekfb2y5KY2ZT
HCNSOF51KTPTAkoA5R0w9cpIE+A1Bo2UHibakw25OC3RcZ/eqXJRU6OzkfH/
jFb8hwStpTdZbeAuEqui+3bbPeVsDik5i33DKXEC+Ld/wqOdTd/AsShxWjLA
9Byq4S2d4Jn65J3ucVSFzmq0BFXFaza4IxnTmVeEBXyzzbe1q+3HkbQ3jOJv
FBulLsD1aN2AMPS6gsu92kykHpnl3TDsoh0d3FpUVMqPupHi7Oz8sgM2DGEh
JiVzJuRuyOnPf2bBQZsMzXJLpt8oM73D/pYKxBMRSEE5Mo865+j8KgvkHzQ7
22fRrYJTtC9ZOpDAHdmfdFD7JY5wiFs8GVKZpYhGoTIIfLINRQEtCEV+HJQp
O17hd8wycQH9qdfrkPE5fF0pxn4kP5xrQN8NxOa9CgaUtuauBmiGlYEml8/7
tcw4slNYTre/evWtcg1gtjQ4vZAH/Y6bYtTfUhe0FM8iMNlYuqXrzMoUepps
+C673HbzV4cP7EiZ+rg6rp4usJ0xR9xBuQPNWbzpZSKOL/FqqFSXR/CRqUGA
RS1AEMJxsOWUJkLuZMz6hBFRofB9hci3U7yso8sxoyWVIliMpygNtXhubNu4
69nrDQfmp3PBK3Htv/8WpZwFu27Vg4dSwPQl8AMLaQF5EJwD4t2AB+rdPncf
LduDmfRz/VfNkmdV+NoaBp9wHBUN0QBuL5wRw+/XCEOUCWtBa2dTitUVvTy3
m5Erkgte8Q2USwxMEOLCpze3yq4WNoCUOnpCym492kqDD6RNB2T79e0pEMWS
9UUC6GuqXi0O9YtY3DqpDgw8sS4MMs6s8Ww7yFG8ujYdK9q8tlSPnZIZfR+/
ghFyuf8J2Fzjm/MXGqx+ACNku8c0EN5dMYmLj3CjBF+VwAIcbppRadyYdFmx
F56MW20oWI7LBcPwaItsi+u5F74bE2N1+xi193ODA0i69qA5fxF9Fc+EIXGx
/FPoQgwdmEkx0UzNv1DuHtVveuxR7aTAzDS1p+mqGspM5GabjNhPrzERleHG
B+ll3GX6sNH3Rdy5AivUdl/cs1jt7ocUSEKzlTB2sHuoV0IqJP6M/ADkpFVF
KblD+Dml1r9MMdSbR0CfYD4zSrjsbZEdBp7kEBDXksZx9vPwfmTPOBIagEUV
zMZW5kVoYv1NhCfQOJR9ttcqZyORsgeJ9WkqbvYTdJ8NuD6YpK0Q8j1odi/6
ERB9KlP2IUs3LoXwebUX33wPMKBdZCY4v2W/aVZ1VNsi+BPusfxB6FlE4Yw0
AE7fnr5dy2MJyFLHfMnbEho2e4AxwHVyISgdscaOa4tpj+9ZSXlPjM6ShmcL
cg8tP9N7uSeJJu2LMb2foKt5hT2PFxqZ73fkCL5nLE20FfaLQydNcLRzJQpt
dTleFO+qLHqkKL6xzNIrBCNQuT35wvwUA2Em0renAkPoHGHqWGU5ueAsMTzO
yMAfhji/CoxA5JGyM/wFEX6JSjI8nPsu8v5ll3ZdqUPFnl73eQ4vHa1xOKWu
6m7K6Yv4S+faMQff2cDkB6v3x+xSxNvlhi/6MGM4pYjjG6pgHqA6sb14OkfE
w9Hq5wO5pBApvyYQM7AAiBGWqgxRxf4EOMJI8Vd1bSioU6A/WTCF0qWtp7Oa
gAZIHpXAy1ETMeftHIiQKht26maxX0eOvKbwkxqSnlhAUBDphi6f5Ap5q9v3
Yt8uz8bogWL8ZQEyNUBS1DNNEMbW81mDGfDkwjHKonxFVUxg8/YXG4hwqkgd
7t2kICTKRMF1zikB5NlTmevQZxPVFPQi8cy/IJ+MwxjeGROwBFx0N+2QFYRR
HZrjcF2+Xpz8WbTYgXNYTrVl1iKYpc2Xz0Q8k0TcKuKLw9XR9yZmsyik2c0R
be7cUoz06q299yDm8csR0mUcbEp+XQIkHJSWsEX+QF2x3eS7GYGL4XDs7BPh
/35LOHlHTEMWlo8agJLnWoHYla7v6HkfthW7rF48NpUUlN4ESMi37r4HTn66
lw/T/w5RtUArJTbpHrPCyn+QMg6+UOGfyB/m0bjU8Wd+WNHyZ0zU2t0MuFNa
R+vV419hPX3+Ii30Wvi3RjUvqN/cmQ4sJER9RS/6ZbvAhdReLybT8IVSoGHB
DCl/OLyt/lv4fhs4CUeD/qEBRSgeSxfV1SVeg4ttrx5wuDaVHr59WNxP+jkg
obJuIs/5NpfDEZZJ5RqscIipTMb35g7i1eMLvnWK0BvzY3ZMN2YeoR4Va51S
GPnYGw5eUuU8fF6EvNWe1HfU+T4WxmRqXF/jK8Aoe1CiyzPs7E6E3mCVn+c6
SjahN1DKe5UAsA/ojVdM41W1hS4ezMP4B7PhCPMoE7U7IMJSpAyP+Ms4CurM
oZGUq7unEN35GR86TsUc98omwKcXDhtC4u8Z7Sv7lwU19vzraDaccqczcOZC
da+eeugqbt9NWsGTh0ns8/3Xi28tT0QpST3KO8LPbjxhT2W6O5rcM/WjBBy6
i5WvugGKx6l9cIVY67ruLc9Kbhk6ccdSoo4JG2FQGznY/iRIr9GyweoVdUmV
9k9+d7X1ktt6EpVG+sucf43knI96xJ6W/JdNZVYr+ZAhEPaP/7BXU/Zu6RQm
fMDqp+ut2JeEFVXwwKemc5zYVahPAXr7cvFQKUt5HocMT0tqGomT6/SqrnHr
NEb+hy1IZU1nskL6yopdUVSLGUOe+fSQQKvInsZRpsAqFp3fjATbUR8kJ2gG
f/lGXzQMdR8Abr9hiDRRX25XnLI85AdEo3vIZ5Bz1+/eeIM4bQtQgTXiAQ14
aHQYttEfMvlHSM5XbjhCm6eoVMETd/EsUg3oeN1S7IJ99KRVx7qxLB3L9hrR
0kZAmJwY9LnI13mqA543IaVV8ZtA5qxsqdXyMdrQ/p8VBHCtUg3nEZD0+BSy
waabQHH4OK/rkPZb6ZaT6CtnGZYOHcCYbGEvdOoLojR6D3NMZ0JnwztT7mDC
7TVC5brjjBFWOMSsUZZuvDt+Ll9P2EehhKakj6lYMyr/Tm1OI/R117+nAT22
Y8eGQBVTQeTR/EMtfp+nuTl9cos+wK7PMYAXMcJLfzujTlO4m87J8ikI5dFS
0254Xmbc0M3JocqZZyybfPcqSqsIyZqIYDZjk/4OIt3N9OOCE/uhimxfTMGx
j1rdny/DDwtaA/4tO4L7ctP67HJHvY0tvVyy7JooKgUXoabwJOye2DEulMPV
CpdeXUrJM4i30YXnq2vD5ej05U6nqLWGSdOT3cyOZ/AIbvSscAiLcRwE6FnT
T5XOxdaWVspxfMzEA+nxsL85DIuUMoupzQGYCo7vXpQ2K3h6bmFxmbeF4uHc
zKyMXYabJjrirZK3HBo2WXm3+pbsW0ZSG5WApQ01O7nPdDKybl0pSx/ZGPOU
tbulqiVL6x+M4tEtV633DIlDOqv/fEQfa8WWyg050PbH4idf7Ie5ROPcfnOY
GSx96TY7sQQxYQtcmcPOyKY4jcwVA1ye18wZKPdiXJ49Hza+VBahL/Q9BwY8
Amd96r7dI6knNnKe+JG/B96UCZj64cD1yloElLO4ZQ5vFh+WX4wyoukZgjNz
6Ijk7xfU+gH7uk9Jln1G8AUQVGtYRVNRo3YbARJee7JNENGJR+ePdLhZgssa
7+gICKLCWy/cT7vcNIfwkcmXOqY2YQUZup2FQFBT6CqZDSuHf/lCy4mTCU3O
eIlIEuZ1YrUiYGjHeDgnzpEkeNbdvf1BCd8c+V63ZVZlDL3y9mOAJbvhKomN
LjaTRtWG84OwWAPR3ZSEFD+hRo+JiXXC6fgO+zr3K3UMiocHdTGXvWhI8+ji
LxRWU/0GhA8nKdH/gG1U4RLqgg/OLM7Ohz5bCDUdnniAcWwZZ3lYbJDH6fQ3
Z63jtUQLa1JaD3qmGpfvQk2y6RSpDCkrF8Y1lIb2MH+ZbLbmeP/Y0bqHm3vt
2GWf80aE+VyaBYiAnZNsWmXGmTlX4zGtbNbqjXQJcsfSl6ZwNZHffLUTG5Kt
8mP4dPP32s+JYntDp5leXe3Dk2rkg50m3ol0HFSm5KuQR0k7yY8g8vrCDu7U
erSA5zhGv4MlAFFm94oj9g/wRyjCwAc5ibSxtF/mpcLCK9wdbi4ETAl4I+g0
/tvFwPG7C3363EDoQBfTveMnq91dl4IP7lTgloTUKoNCan6jOh16KXx5C2ye
/gBbggoncGZkDhHxVBhdKPF+93cxowKeeXNwyZ71WFvQs6owhg62+vj5AwB5
Rc5qVoyM1DWl8SqDDw+DfXEbMwVBN34uCiU+mUslJfCiWtOQJ0jptCyjxrEp
O32WGzmcjyM7L5wccWISGsjQmSCpIKVkgDHudTTgSQd1tji6fEPosx6LSXOY
anBB/6SEHOp4yJ26YC9e+Bxs/SczqhlCcn0gm2aQMEZ9DETxLz4cvkRPkfaj
jntxvJdo4jjTQukvV7MAYx3gnpwZsrxrq9IWAKJMXHGwWUuhN1dtcDbcHU7o
xoPZaWgAd9JpG5HjnhT5UX/MvvdeGwYHXKzE31rKafxJkwlOJcfrf5H3wtAe
o1ui/kVDRUODinsgT4ceGdyLTYWKyBviw2Bfp45xNBw46tlx3TwC6nMj6P/m
Rky95xSQ4tMBhjj+dG+csfSO9mKHVWo+L3H1iYJBp9pkTYVZO+/qDIQRqfEG
AVz6PmVxnkFUZ1GqDxAbgsc2EJnHDvePheClzHcaXrM6WmJls8bIkbZNJUQT
j+SgyfbViUnY+ufpRziZHPF6hmLkmUoifPncU7nD6kzxWKq8Wq7+Lw0Dh9RW
xo4NbsbtG63ZPhHdk+B0ZRqfZtlQ+OkqAFKRmy2st39FOU4e3Bk1Xda2iQ/0
wTKmDo42O6URZht7S1kFuqXErHLuQfBPS1ex14RqWdDuKG+g7yPTNtmVlkqj
up5N2hchQq8V+IESz7Rb+ZCrg7gm5nFLB6V/dRh7gI9qPpyzzpSLYSn9Go5p
x33i5OtaFmFazCSiMmy6QdxvhIxHPcFRzTCXO9jFTdYK0iX9Q9FLguwwxztk
NsrS+ngwsw6ZEKNVa5U5kLJZUuUHQuOJggwu5pFlHC7hs7qwPllZIUNpWyu4
rjDKr43vZXOkKlJjfUlC6lhIYEqDdBnCt5J7dAnL6EJpWFpd+i9/0TiN+LVb
FE79gYJ+fAoKUhyoYSV7NH2BEnuVhioOiLm6JqGVXvk5v2PikT1DmmNXVsBl
Hdl6LOf/AyHLe3DyW0fSd9gnXJd4bQn+Ig8kR7mO4QDOj+tNZe77jjCmfIHk
5YpFd5BkqkOXMBIDxGiPuXF+Z3EuiNp2h8eaGJyt1O26WdI40Z8SJ6USW+Fj
Iqf2eVOsf17x6oCrphB5h8Y1KDTrkdk/xiKQOkKZB3fwZ1VFaCP7D6CIo6vv
mo7VLLxTmdr9Wd4dY5QywOqcOOHkjclGnLnYpnepo4wAT/UOKehDD2fl2rVD
KzkX4NVxxTwZY/rpKz370V7yr38MD+RssvDOwRpzrf1gF80D8l8TsrZB1sPM
MHLMLYMYmJtVClxS/Cl0c7fQPJOu6Bmq1IcehFM7yQ6MOjPUMrsSTm28i8wo
91VKXZrjmP027Tef/iFRLrKefj6krLGB6jxsrDSA7PSWpCvSbH61hjEbqmKJ
9glMELQq69dbmX79aUc1IBulg1U/llo+ABzjyV0VM6nE2CmXWSP80/8IqZBA
ccVbngdEC0MYbaQoTqGaWafv5U8ZAKedKj7BwU9Yo/5UzdPY+ZJ8gunCfd9E
5IVm5jJEhm1XY2C7A7W/GMZVj9zrgKqjosyYMDgJewS/GuuaPW7nB1Yua5rF
3J+Ozt/dVr4xJ+ErqnSkY+tT/xOsDK/kV8NdtXZJ+zG1S++5EW2k0wsMCgOP
wMQ6jMh7UdiUztd/hN02ztabGr/Ezl0BROoqouXuMqryhNWcWPZaX6fd9lXe
u6haqZj4A4tEQvAuVmMfCQTSKPeMiCgS6Ew/c0l5NWagFa8WC1G1zpDb7+GJ
yOkzU+xg03+pF8hneNyE+6xBn2R5o3We8wgHw0Oiqow35SMyeY27Wj74bpLd
4y+msgTRiNgjZ8b4+gQ3rAsAFlns7xFuVN98SRk7xzp5xItsdJDj5280w0jK
1BSenablQ4yEXBW5LRrqFZQGenc7J0nVEs7n9S63ZpsJ2/9qRMU9NxiI/Viu
/fSwVtfZOP8x82VcsB+Bw7k8NpdbinccDsCuhyEs5ov6AU1yEn1J38awszkn
TXx86DcFL34BySaeF8E/uMAz9gbqc90jnnwaS8ezJTnqwTrwCG5ef6SGBezq
ntboKBrqdGWVNz/rDrNbLi90y1AhajGFWUp9SZtYxTpt4jteyKmKuNh1l/C8
KMQXfWjTMa86s0jCYvB00pKUHh1c13mOPjmlrmb2NhhrzRrQHaccu4kSXwdM
PjagoF+wIZlNEFHfriaJcrzyFH1nE1vcVTnKLrs6xI4Rhjz8IJwSUZvJ7MMg
7m3tYs5oLIMw4iVRFSDBuSsXUmrZvmTTzda263DVjRI8oewpVfYV+ZKbrP84
3w6cN3yykhPibPXf+dgdll2bnU6exIskghqMi3SlfRIrKImwzMAwjHgj28dF
0piyDvA73TUScLezlS6LkWCT0kq9oY296ZKa3BQLt4v7rE0qrgDQ9nyBZjaP
WdICX91xUuC1yOnjRt0Ojh3XJPOjFwocaabxJPlX3flsA8JTbpbZog9Omys0
AiV+AoVHN/7xrsnG00TI2u5cCgV5vtuk2lcjx/15fbgfQrLwGwdjqtiKeQO6
YZuSeY5938haNCdxIlnm/sSagsq2IspbyiQxP5tUVDr+e+XfyFHGtG29BoXJ
s3mBygqiZJTmlxRUqslKFASnPBk0BtAiOQdVrLbAqjLmFnLVubXze332b4iH
A2GoHrKXkxgI71T2jNXMy0VU6TgOZCkyQ3RhsrQDDtGryglhhdWldJJwm1O/
EsgqRGA1lKPcXuAavWH4WC+NmYulaecrTNJgJ2PO55XTPc2rYAj2TpVV5i9q
9CQ1eR4C3Q8RyvH3cAjsLSKmiWvU9ZrSftf8ZbOgzn350Trmy1wG/Gsd1bT8
toCVIQeTKMtJZ1uH1lO/EkjDEVSv/MlHDYxL5jcG03poxkRyHwGx2noH7Fny
+AZB3U8xpf4HK9v4yFJmSMSH1RsJQreQvoYnUBsS9mFVNEH9oCCIUiN8lb6C
VqFJzBOvTFQsjt9wYPks5SNaLxDtCgfa9UFTJbx1sTxdxzd5XVIEIMhAUDvr
RfpWR52oniflI0bJZ72D5DpxuHyQeUwJnsm6eLGx9NLC0REo9lVU641K7L87
cJjjxB+XMpBogI+xcQQsyw/pz3pkoLBxkE33o9tudDrtBDBvfGTXnAxrAb8F
ZWpO605nGPQS7CyUe5xqYjbXwuQt60/DSfw6wLrJQhT3zEVZ2mj6u8T2h2ai
lLeCvrXWLQnFutV3Qi9gSly7KKsB3as+PSNrI549hqGS8YQrjvzarHBPzdCb
JAyo1pNKC+7EoFbB9I9so5uefvI5287ywN8f3vnD9CnOTqA5OHQu/j1p//xv
l1wa2Wq+IOdI3r2u15NSXifb10W1dzUHMD/UiOTOnw0W9AMgSBhh3izK75+B
KFOZwBl5M5E58c3H34yGe1U+NMJaTxYxmUZ39rxATWA9hpaCEXZs1+/xVVS+
nlSPpniYxEo/3glyNOze7v6e/QIUj87aSOxacVBnc5AS2srgwlj9aHbYsGLc
D6GHPqauM5DrP8tPLN/C9AtNxchamcedUigjiDIZznzqBfTdD9afd8loz3U0
JI7MzeImvCz5qQNBY75JSeej32L+gYBVLRlwh1PKLOSz6nmGG9Um7Dsse0Zh
pTkaKqWiGTUEEskRtIQDJBP2PqWbOE2NzDJFG+zCURh5vHa4GAGUqP1t3AEg
trwPmElhpM22YUrRc3PUrPbs3ogjSMTZ52ah7Avx0YSOcoJZ2ytHOr3MgIO0
osAmry7FF+/UBSSwM1P5CElf0Qy7qjh4rJnVI6BMaefnDJw2uRv7SPEBB3RU
sgDNeEKfMHurk1Edb85nfTGDfHmifJsDerCndSxDLWeamy24tCcRQthBfgOG
+rGe5ZZVIhr1Q2iT44PAbBraFuw14lVH2RcC7/mJ4xGGIjxQXcSL9jSBxHdL
8oblVqrvux2oLOf4wpb4/s3LVHlRLUimk3X00TtHTqgra96tPQRS6SgGh8kN
nSja6Vum52nbzFO/fBNJ56I/pz6Qe6zMRvf6bisi2CpxMErh/QIuSrxgI5+x
9fMhihR0YexH2ApR73WTqCHV+InK9+YFIicn3VkQgiZHafzGYqqIvhmpBoCb
qFB8XaS+1BFy5dDh2Th4rWgyeHtocrTM5HtJFM4BV6TXMtF2dhbIvaBKlFkq
LqCloLN7Q/fahVrGE3FvJIzO01PCg87uKdOMiCus3Jw3Kn5JP1MwO0D8QuB+
kAEzZnKyOqlWV7GnWD9nXjLB6LG4wCAWF0C9EDjCPz9Eo1mam/rCeizmBRpr
QFZPHss/wn5Sjjbh+Qe+4OmI8SxvWqIz9+an+4zDyaPyFGATeW4XKPD6IgkN
ZTmNGfTH84o6tvfSCBGsMKTyVPm8OGlzousu1PKPPutFl6M7AVrk6OjqK44o
548U8NZaL3qBfJfKuvFsBTSJL1icZfJUbqsOcVuhSz/aQnS647JAx6huJtjE
1mAR9zppLManQqFC7eA3kveMahgkrY0mjhuynlCcPMHRnyG7tNypRUonP/6g
XIeV/ps6fsPbnjv4sCexRwmaJPe+BIJjuApbyPY0epEWsO1LdYPvQD2c/czT
b2Etc/Uen6wv2EhacoT3qzNXzMMkobgpQP6Xh1+zpE0ZfcEWpWSNTYX/s9y/
JQCUH6F6oakh5x0EFKkAZupcQVagzNKM5+cwzoATZDv+o8KnxlIlFwoir/Ro
xTfvDBZ8C4mN6Inx5bDfAtH4kmc+1pxvKykqo/PapakTuPcjWcoyXyiZboSo
C22qQNJFy85nUC86vkjgwkOMRLY5OIr7hjvVMeAkBOhqUNquGKtgddsYlVX4
xf3jfhiHW7MGTVZ7tWJHlyvQHxE9iEM3r46wCrrsXtIemYBZBQpFKIopBzDK
1H0lkA/U+U4PXMmzWh1RM33dIhpJ/MLS5JTD9QR947+uDj5dGZDHQ41zp79B
l61dOzK+SFU9leENjjCxjuexOnaaP3bugaw76CbAx/XbfLgt1O+hnhDnmf6F
CNKHBiWvQRn20kT0relOkHQpl1D7ie81PnxWg72pP3fqEn1bVYxlZLYmOhx8
8E7WCPTDoHFxoiNOc/JquovY23ZXSUgXWAUVppIwKSwujwh1d/cAAVNNIj61
Lq/xDk++xZosIaiGFPa1GoyrHTenTmAFXnJjc7qVo9dKILC2gMuLlfrEQoX0
f3zbU6qp3CF+8Z2M+WFy4O7IUWYqtBtsjYDouVd1tK/vgINGLV3ahZ5Gj0p+
xPOBusUldCKyVIC4zJsqRXD28PLIof6kiYFPHX7isnsoVhzJC+zIdRoP8e8b
x7LNGEedRgAFKng1idsTIs4LmngzAAywRe1eXPwgH8Zr0aK/9EerYuQVc6yO
zL2vhHMVAOGKDhYCbxhESLLsZRnEmkK1BzYA8KRkfcIawIE1Qj093MSCnmJH
bMaBSQfw8u/lkZSWPMyHbbo6zwHXDYVK2bartBJgPaMZYo7HmuDWMqAeZyOb
UXrradpQYwKJO6PPEVlHmT0rSrVwG7WSm115qNzz4uGcuCG+fqUYuf5klRD2
sytfLupOiZdDqwFaXsIizpphKvs7axyfJT/0FbUZtipllq6D+nLBtyUgQy7n
EpXLmsWbaCzYl971+H28KLm9Edh+eiLFE0JKeP8ZB3ciJLcYdf6hdIdObE+F
PfMboINGHIo3jYZ4EfVxp48xKr8Bo9LhJons6CimxVt25lUZ1W2CDsw23lTr
t8kBzdNZLCax91ouNUPerXleXB/84df7WME6d0hhHr4tD1Ir6znhFPOpZJsd
lomJRMI07nfADlyekwp+fuBTQr+idv2J+lDQJv4EDwteGwjxma9XsJ2HLDN5
wv2oLSLvY12LKImf47xSv4PC1x8V7BqRXTcItc6KRR7hdAXSZHd3ZLWvTrRi
HYvQFhIVOAyTjdXkbVBQiTXeWZQaRgeCJMQkCek3L2ZmBXqj7BMFU39sUJm6
pSybHFH8M9D8/gnxg9S1il442jlux8a3dTe+354WXaN8IoBXkwd1zy1Qa+Vc
EnQhl1WLiQIGAYN6I6B0f/N2Ei+XCtT/jCcFHplqAQChcWCrFgo2iqnbk4yt
7PWq62Ct4u0S8dGXO5oiZfdedBK+GEs9wEJTDOloKEMw4hwBXN+1lZ+qZzXv
d3uG5d0Trm/EYZta7NPK/Yta8No0nuNwfgDbtUQXQpRyqMoP4E88koVuX7tJ
qLU1AwwQxETYRAWkE9qtRifcIl9OO+EWdw/eWZTSYWL2gh/dUmGJWjwPwDdv
w2gqZeF8VvjTPdS5gVIe/dnrMN0dZpG1QxJDq1nrQHDVkgQ82QbMnACeys+H
tzUEpC910AvBohhrjj0jr3JiYIMsI/VtK6PNlCnfPQh33aPn/fGmx5MyO+XS
mqSom5qjJBGDr2mE+nloj9tnlFfZEm/fmKB5aTZ4iN/+iJ9cOrSQZTAeY9Lu
7NwtGpIc8x3bqFt3nkqc0bAe5PFtxq05Q4t9YcIiHg3t3jZUu84Zj/vudD01
5ljiNFVZtDfD6Rs6uqfU5wMgJD9yvWIr15s7z7nKG+OJXoXaHJ6YRNu6KWju
gdJhTAjZXzi0dDUIx2A1E0DsQDW68XKlJ8WJLoeyVyZvDG7kbZsC6pHWJ0Se
WBIg9Q/jpCEcJNKSmkqvHSV4qwF0+g+0S/9nu4lawCyLVHPeajL/f14RZjaM
qhWYe5DoQE037zyIMfvHXfeVjHwARKSPVrZv/6d5o3C5F4UfKcUMi+iQ6Bfh
HzMr7IW0/D1+3CMGCIxDhJWcDaEqAmvlfbRwFga3RkFanf0oWgxKLkfQJ8Qs
MrA7EWG+csD//7OsI20g524w7VDRmfEyxZBoi4WX0jx5BoobVi4S9inwcGI2
a6PNdBQlz4FDIgxGfgLI2BJ50525UIxyNCc/HdgmcLHErRxCJFZYPX0lvgoa
dq2GWzY7MN7Jax1sVvWUM4bVPuu8XeH9f81oRioVpCy1GEfJtdBiL/nKv1++
r76p4OcmDbiEeAIoXFbNSEieTI52iMjkcEM8rR054+rHi/pVMrA/EpqXs2Ix
6XmxcjNCQCQt9EKjVMZ3YjaBYP35fglWcEmdV+MJLDCZCF1ChrPSn3hA15wi
SKix8OVaTcpOHuYS0oyIxo90eanU7E8LD4CQY9o2pAkQQVSsPM5wb2fk3Mhh
CxM6mcfCUZ4oKdBM6+VRbBJKmByJWKPNUOCxJDOwFzcHaZE/DCIszyPwGNi3
mQ/qQdVvEz/gvEaXKLkkOt0cB2TLBBwJ4pylzmaZQ7d3g8FIDXXJW/WJVvxg
ROYdwCcqNk8DNwvMNfpNZLl2812gg0kc/XhM/cM3PRjy3T5MUOOYi3DsbHEb
ii9bsla8hUTwSK4TmgLu8qI48I8C3mUiy+KneQl7X/pBIMDw0qv2VNLqis3K
LPOdbQ2NWT9sz/HQRgxAnY69/ZxIHplEXizXInOEqJia3n9OGyTYXNRpDhg4
JWVY61bUxCVPxBd0DIUjfjp7OJhJAbRycodZG3kH5ZKd5UWLuCl7bym0SQgQ
gAlVSwdH5nybJ7UCihfYa/Z8zorWwvVGr/q4AJHrOJgxvm5ifbdEsuLNvOcy
ob3skHXujvDZPuhkhRQEdvuC9rNGBD0Xndh+yqxcwhAb9ukiv+fdos+tTs4n
1e6z+Sr3d9tccREZJ4P9RO6W936ubRoyvPgGalzKFKutakcAd6haGFS9wLf7
jdK6Y8ntrdBnNcKCahz/j/KL3+WjePBYjda87dEkBWzTdMVqPjMZqpVIn2ec
+7nrk2t9/ODNedBUFa13WTTj+k7RHrkZLKxiP/397txoJitvm22rGKbeAx/Z
kM46cKkjKI8NHqFtlce8JpMOHqy67keoXe8TNISIF88vA4OjWMbe1D8sx3ud
qe++6WIM052YpNJ+HPagaJB73qJXATDo+mdIh/gnKdpk4wCvsnjPqU/C99d6
H5F1GR//DKG+GulH9KKiUfX5/egGQwpMCApwcxzrB9NAnQJwIdvAs1zyXyKW
2wDJHTC4QbtDyx7dOkWqUqfwK30faVKfu2+9bbLI/p9c7/ABNTUl2aP5simu
MnaZ/dGFw5fNudw9TFhlTKMBBGxyxzRU6lYixTXJoRw3Cu+qf+g/RBeOXLe+
WbVAZdz/VBVuR9DeN4uWLr2gAtreamoFjmZdMs6ic1ZiAArWIPZR9l4a0rpg
ztnUJVnoDlwWMLF8vYVdGPybS3f1QDA02Spl5m4+g3i2Wsgg+f42PfIdj3mf
pJGRhNYZXXAFUWyrsmYpNDFq0yqpfhq+ZVRItYzBj3/DqacP3wVDQ0KLzYAT
chhskXAwBPwcvmCuIYFdnwibGzle/ieZ2ytuU1vga0i9QzLFHFE7stZSUchX
bt+QuBgRLA8rxDeTLEfTc6+dUWJkqAI815NRAcbEIphr1CFJroHZllxp1aKr
F1fJyHOI9DZh7gb4mrG400+Hn7z0GNC2OYMopZhoGopUk3erTq/j1OfB7sK+
v603xkG4jXplgnyLNFotUYG4ftCDGM/FQExqC5jzEBSpl7scsFbK25C06/Hz
mkfE0ZWZyENDvINwaIVudd/oPJ1/jWzUmHx+YtaSrvnF+mvlaCjMjD0Mm5yy
Ns7cIn6tVE1BTRb64YWcV2N1VkpqJXqeyzRAwycPMUwah/ebejpjR/mOtA+1
VyUjRAoJQZn0SnXg6jbnkFVQEm8i+DA+54hPXsCpQPKD3Dj16SKELGzKhwqc
B/yTwWXzY1Spmn9XmjB05N9guXHpnVjcyaIr61T1UtN4LhneNU1npPEeD48C
iuEerDr34YQY6bywbjFCepwqezzE2BFBoHhk8rexKAqVAxwgH7vjCbqD/GSa
cOKJC1vqrJC7eSJQ7eiFS6hbTlEd0d8n52v0YHDdi8cgm78ApVsiehth5+RR
EChfp9Bw6z9l25INw+8JIzdS4ucojnY7gMtZxpU1/BBIJ+ho6QmMZNdCgHTV
xcbloOwowm5Z0qNYtRk3Syn4Rtfzxmp9LzCpPj7brpaP9uLtlSQ5NHtLiHfM
7wsVP4Ag3qstd4CGtdKam+joC+Eu2TOndOZQC3Q4vcfQ07l7J07bAiyEax9h
4PHqL4Nq/GsxWS5aRg1dDF6w9Xt1kts7uMJkj1qKBGdDYEXI0CCKgaaCF2aF
yJwLeGkY2DrIGbV50aU+zTAdtD8K5m7hbkWxjzQ7c1rbBNYmClHCSN/1zd2I
cfmoK3Hjz/IKim438Sr8vPU0FKD5VFv5GSk+8TE4+fs8pfPkfACZFEKI3Lq+
0IQ7d4dkzqhaR9DtHPR7QockCHlZzXL/FigDEA0bxCEEh5AA+Z2brmrJw8U5
L38A3FACWMSsjT/wkaFhCL2XpM+ZNdDWPUzCL5AYwBtE9B4tw5nWLagArycP
2sKyqo8O4Z+OGJEnb+MmxSS7un/68aKQIOKopYxUAyodSIfwiTURHF3XKMzt
7Gndc68eN2G0UWmGR2Fb5P2/NLNSvMpHGHozrixsM4M+WEHV2GkZWngNJ1ib
If/CDpzpXEDyOW1lU7V1Bnzzf0Y2e2WoTASP/kQmqomORlQXHdgtygQTl6tj
j+SKYP49OeCIbhZqAu+LecssEobV9bJpZU5xz6iO6/XyN1qGunqeKo+HpdUS
pXXkwGfKfMaQ3FqlSVP1af8S/kRRQBOZlde5Qmq/qjox+zWlpH+mKX4+M2at
d92rPps09mQxq3/sM95MzdZXog93xzZm0r9ViD2yCc+ZVNsALLlvD+e+Rql9
OpNaHPEz+9xyQD663QSA/12Vj9i6oRIHjt2qtjyGLk8qIPW24v+j6MOmuSJe
MCpvnKScb67Aigcn8jci9ZPvauX9kXn082smrjl/viXFShplAdOwLTsCHwh9
Em3OO3X0eKC5/0QdGa1mqjZuRZUTEpuG7xyarEV+7XXlFdMJ4Vl1D0ptpO31
J0/3qUGxa2YMX6T04Ofbgw61ds7NS4K39KbyF5xFKalvqMBxa1vCxuaCx0ua
AR/prTKjZeft7VqzlT9SRS00CVcJfWOzD1gXYCB0pgukLNfamcbzlR1e0e3H
RgYFbCRkV1VY/Yp8pidLzvTiSiD9rxWH6SvffNlNuaRHsxRXsRt03vzfJe5E
quhPNTdRUTXcB4g7OAQJLDOtnNxv4CfeE22TUrei6/BUJyr4S9xet+lljtbR
DCZnCv/yHC2D6xeJjk5AwWzj8c/oahtcxuowxhuVtMKasssA7ztZiIHaJnEx
h63i8ErjkDcs9D6zj2SsTBL4ycEYZiQKrHR3TQDOtXO7UBTNln/rpztUhFtz
r7urSDPLRLGxe7FmKnjKxt2htwRMzdn0BdEvmC+LfDqJH+/QrKtbFN7TX0Ho
mq0Rj8lNzLpoWVRXkdEmT/QosreTghyU8trfy/S5khZZbHzRSTFlL8GYdvyJ
E64+YwjQl0oJyq4oA95mD4oCbDHjFPAwO0Rt/l9mw4BRkxnuQm9DRbtfMrSP
30vC8G5dqgSamK0AgNTjMImD0b28r/fPCP+2KwNMykXjKwiSHqyDzs3VnRtp
r26jxQZWsKc7vYOl0WcsFr7spmizt72i6HIXqBXwS/UQ67Ve2BRrz3axSFJq
HZijCnpNFg7K3jV5lfqUakkbOPaIeLSX/1jh2qgnR+rxhv2hYCknjOJkiXW1
yVxgKcrGW5up75ZwvDoBbgfaYSiamHxfu3GzbhKNq15w4Bd/fbH/A+b+yF87
2hInhRsAmZF9VnFoq6hle5UpeGh3wVwK/NnAyFkcsyolDx6v8pUlNT7Z79rv
FxpWOcNI5Bq3iG5IFZhFRVeIhWkSZ6GsTcl4TNjMq7ClNGZzBWzc0luI2MYT
IrA0rlBl8NNyyNEiLPRPA4WRWp4KppzL582HSty5b/CCKkO/Ve7P5Ywfhth+
v21fnWUek0Iqvnn2MW+FmiBkM3pn0OThDPtYjNLP4d8e3N20+Y6bOPMUxh7p
kY126uAeM77a+cwPP8KGymcdBpSRqsCgUjPb9M+XhJp8IQan1nNdg+2nVM55
b68hC7njiMeChJIBxDZqfnERtK3CCyFifdjpW3K54tspf3Vsvzf3yuU/uucQ
hZqVa4cSYZ5bjNDTmm3h6PEfPC/MWhrobVBBLN0vxAj7A5eT/ERU3iAEUtn9
Xf6iJ/uJgsJZRwr4bFw0Yb0zKVau5n6J6rj5myLUQmdp0Y8Hldo6sRxJJPj+
yyqo305ovkt7oJ5xHCKCmxnK5vZRwdR9QUiB3qwlGsRwW6Y1OYdX9DIF5CxV
H7XbEvtxL9irByCpCDPQjDNTA7z/EtnciVtDi6cFTqIxWRV8KSSmFLlRDnWi
S6vRP9PjlO7rTgzsl5iRJ9RtYugSmT7j9qkO0sYBGZKvBcq5N3kc7wmglUvk
vKPbYJbWCF7YGHF2B5lqUWrO2JzYVXZlXee3HC5ddvkSd7SMi0RUV4+65dF3
Aer7slUrtBZriJWeW0q060xN8iHA2qpfF0j9lMMHYuKZEzvbaj9PAMmAgRw3
rEHnnkZpVSMwzM+R4ScUO04qqOcxtpuHzDcdQ2Pi3WlW/2bU1GkvNbzvVkvz
4i/1oNQlbyXZv/rOInF2ppeJBfNDQ3KbbM9SpZeBvh4M24btIS4GG47TkhOY
jgdnokego9hg2xtLMIQgJC8KapP5ze4nyN5rkXMlFAnhVzTju9tfVoveM8lM
VClnIe8dYk7rVq2BEqJLRbnO3eVN+IOE+4P42fxsta8RpUd1qsiH8A5Dm+Vi
ZOFtLfn+xYUE0w5aNb7KwtIrFqYwoBAM24zTtpQnFAV5ReGichsw/xXqf9Qn
v+qgUdyFuhMHiz7GJkYyLmCwEKA4JbyfnFt1fHeIcssb1L+0nVzwK0/fVylz
hB2TpKtxxDF+SEXoQRcJADKcTHa/ia/FcDsuSsHR2pDR3au66++aYPzlS7/V
yPOf5IZfefqrefBCCrPh3mSYXifx/QiTPWXVb8MgEHEnCBdzcqo8WcAxUyfL
xEs+/6UNYb7GGlyDL1okImOtKmk/wbv/6g/LUkt519+cRC6jgsi6bmeIX5gV
DbnyfZ27LeCJr9MqIYrF6PfVt6psW+sJbMJd1dQID5EyX+A+KvxlX/9uftzA
QTG7hTreRfSUZtwI+es3woqjhHXukKZZfzBbOlWQGXvm3ZlTQXjk3e3UKrYN
71uz7eCEfIwx0H3cub23PEEYMYTUzDaD6+5QWB0sds6sh/ZRhEgzTptSvP+o
6OtCOLI2ibBiNk1T1WlBE7wd4udhcr67XvhAj9kNXs1PZPiV6elhtTNTsdiN
QouDDcPxFN/49FQI/qTZJjFYMeVrfz9vsLHZunKoUzI54ZkAcZE28Arc9UZY
ATQom2mq4U2x0uPQ0SEWJN99ukORPdLbUQ0tiAwFlQrmnPTSue6aV1iaIcuf
VrWN35MTh7p1CFrGK+dDW11XPUsIv9krkToMBx9RYER9K4CF+PBtAr3VVsnf
xE3jU0jcS+djoPb58gT9+p012ljrKThyOAvPUZLsHJ8iSf77YNKSK+5cF/gp
TBhRytbfwURx8dObm9MgGyFJUamb6umzH9mw/e5d0epOvXi8E7RfMFtorNfJ
VxKF8EJ+ij9MO3loE0qUp1XkkRgU4omAddpkaJZZH1qIOsKTHmRSWEYirgiw
9GPtfs9KGUyJy8GVlR39TwBxnAKx+8ms45KBMEHpCAFXydIWC4Pm1BCQliMe
8S54MA5BtL1AyF+vjfyJafW2ZTzVov2y1r66g8iBDKOV1pjxJnxd2Vklrarc
yGEzoT6aEjoOQ7r44GYd/xA+7y3p/LgaNtY4a0mOXyA+v0WMaTLsliDNgCHG
RL16QXMGhcodGICM3SAeiKiK77OgXvBO3ieukcgSc9ZrnQIm9wWultCcW2aJ
7hEfgzPA/Oro8J6TkHP9LfrFTwWNX8P1mQvRAhYcHmOOA51byiFm+0BAsKrw
Y4/M7pE7hjNrG1EuBw2wrP3L8XnTGShitH63M0Jmkcu0A+Xs7E8ydLmmyMc7
B/MXCn5jh05dRZzFm53eu5DQET92OyUII5B+VNaGs8AHobiIjPEIzoMb4jEq
UDZkdHPeMD2MtUsRmU8qRxgYSZ10lcsGkp5ubhDGNXQqI67IOoJjYr/WNC0q
PgaxrYobq5dD+RwG1eVTbgSFRj8M5lKuDRcf+XIt+ArDmEnzlQ5owJu4c0kC
BzNXdbqoQayCQ2YtChLJLaEsggoONfxVMQLzx0ZiYd0hL6v92jFC739G8r0l
ZJO3qJW0ZBRkbb5YJks5Qx49iNK8xlwxafZbXP4IkS6J+u4WMxbqGVKCafrD
qHfKJ3cbFzW7fWUGK+1Jx+gRB20MBph81nnfErGUlv9V66HIz0mIQb5mDdVu
pHqXvVS6g8NSqobCjcO4acmSh5N6IV706RbE3p98zbd1VAKvfBNNP53dEJfa
ks7ueaxTSUmh2mJxv868LNY/XLJpZ2Rpllq0h5bEOtSv4zPZVVfeEX6hRA6e
4hR/hXToD7FCjLD9/zECw2h45IsswQt9yRMZU3xGbgLh2suBIPcPyJD2nQL1
aD3IwGJgIQ2QnBdDo2PilFNJpgKrQsuxES+y9mnXDDasIqD/4dH9lH4tgDEl
9Z89gT/UnBkZtswL0E1ezPh8o5fSL3U8Otf58kmLsiMPZ0/yzvdpY8f/hDwQ
+5gwzb/Rrq0nxOXLV/Gc+MFjKqKArfxevvkjaLRj3kdRvRcYqvj9gs5ZOJqB
KZL/raAXLpp8u3HDm7wxxJsXgWJZ3kdgKewhwZGtFMmis4QVoN+OxqjCAFDP
DetM01gLzCch1/T0usohUas1THh7LCpz5GcoBw8hsSHp8ns6k4M/aA8yU6fu
j0D75V08mMRzWw6LHeRudFg4RiXCLAlBUf8MhxKwF+QF7irqMLh1K1mAQq8k
YsdJUDBXkO6M6NUnr1aty1Qt5wn7UipxrMi0x1ScDSYA3CKCejxMO3B6vA3T
IADz1w039xAXL+FQDR9aUQYGGfSIpiuysdpbZBRG7aU6/NdBwP7Tfm870M3n
tZTARZqSLxyBQEhhXNBqV7i0COZBUiVZsrpqIrI++fN+dJEi3RMJhif4erzu
vJiFXULe1BCj3X32hj6+QXIbfmQdkEEEHHhQJpYYLsLz3IDoROvRIufipJcr
z8m7Na+G+YhtEDyo45/in9VstXRTovTngWQ7JFH+OTPTljYDlkuMaY+bEhRz
xH4BCZpeaQdefWTPmhFZeYQ+KKgKYHh7rqJbplDknBzEXjQWE/glgumST8KF
7N0cQ+5b8rnjnn2XM1GtptfTxx0csMFEdWku4ZrmsO/lLQmhL6hXz7CDa1WA
aYT+s1ONZs+hM6/8UUVNd7wYxaFuEUrYEFtio7Lw4T0U3gDHvQBhgv5CZQeM
pE2MZKodP9j2LmAR7BpFNB+vHkp0tSPZb87kAmM0fYoaGz+tryvP3ncwFvuW
PwdZYT7zYjk2D4YxMoIydEnZK3gsHi/L7Z44jhXca692Ze0ldCPmSyXGb0Gr
A2VYSj4PrzGDBtNbY8A0pC7bbOUHl+PhZZhDRXb1C1cKJxGeEHW+h8CN+ZJk
mKyY64NmcMKlDnCiemrYFbN2F6sZp7cdrcpstzuBMKti0RW2/zLIBQerSqa7
MCdFlWZJtbp6/3f3J/qgZ+T8AanmOGcgpg6MOrWjiPPXEP3ZNwarMBMu0Yvg
eGkxW7QRU191CLSb+gAOZSlesHh4zy0ErBFsmFfL29IgUCBHXrnWrruzF1XI
weUknNJOl3j3dDik4WlkDlFDbcNePJyP/fr77aXMjlJIN+e8D/KwDbuoyo/e
jQX6gdq2kQdlzxQHm4sTSdESfs6xUXq7bZWMELuPGlS+sJAFMfuCy9ah34d8
3yh91YQ+kcYPG79+Gg6dmu0qBbIqdPl70j1FqW71fjuOboWgtb5jD3RV6BS7
Eo6wV/PdlUKoazapINraxfO9djOcxBPxeAAPTgIrF4GkUVXxURHU7JlFsAdu
Bk+/hBy37TLS6tm84mSXsOsObHgsQt82KAb2ZD+IWENFQSlKpWQnyS8WonW/
2YM4Hi3CYNXFwod1V2jBY3o1xICOHnwPALG5M8Y0rjr1z4riK6z8GKV0HnHf
YsKdt9wYw9KI24RaCT6cfaUBpeHqT7kxJR2e6wt2pOfwW642LYGcbDUSOM6+
tPbYTjSox5cAB/+zY1wwwMTFH2TwN1uaeQpu2ofpbcWqpbuk1ELB6M7uMoyY
YUj2iWzozxnX4UE9jX6U5rt5DTsXOi/g9wvJXzlIXDUWvk7wECqycXyGUnc5
rG6ER2xxy8+Jj2ZXfp9EszOanzomgwRpCiTBU6Rj88HIrEsuDpSnXH4sOu1s
WaeoIB022qNKevkkHMsfjLdCwcHBztmmoqBPaQ+TbcKJUsJ4vUe27NBBFNEf
bjGg9AsM7XCiecgn2N/BiR+zvq7Huku4Hayu41pyB0RC1PTiSMwY6GQtDvSW
FSRMzAotYYgmPFMv0l9IZRadSnWkk0kRz87yTcAvdf2FFjygUi+wy4GgxnzE
DudGnEqW+vqnF07EZhJZ0B8FGpVWLa0LWjcGq8+xNWGGcoR1P8RAVBvzDaXL
4FuwHtibHf1JJ2VxL8HyFJbe6ixdovtZdXbI3vhLw919aqDDfdr1Axc3cZX/
iHWLXOkAhSRy3/QBEhi+xN6ENCjiOXhWiZMrdc7yjfMP+ljsMvV4HPDou3yV
SMuUd75uOfp9CBVN8MaHa5M6CbB8/ioOA5g4SgTws2vUCL4GJxy2GYX9/jQj
W29kJKhC8XpPZK+keGi8VSF+c6kwGf0ewrA8t/cul3dUXI+2a1C/f5KmeRqg
fVVcYl0isaljoBfhsx1NCEM0Psil3pYRiyat/qxY+H/Lj+Sb2OYagFauiFj4
/GPyjIiJ9kGqjtfHNzDnTOy98OzQIumgcgYdA44ItrtgJU6Qr57S5doRto2J
+5ProswrIb5e6DyicRENWxve5kHzEO4Uk9k+Fkvjo5jgIgcz5cDjZJzGm3MJ
qQj0jczfb4FkNURBU0gJBwpVyOlTWfG5jXCGfnENqNNuoygv7rNgmFJ166mY
XR1M2NZX4ZAxTrK3snhDWE0Veq7kooVBHWVvB+hfSKbu6tjztDn3QiIAFGGU
ZqRwxSWWR7HmiibLzShN4wNWZIlc4mfeWVNMKvkqkzthzJJq2kcJ/zG0yvs+
u4TvWuwMPZqvABhrMXm2w+KSvmKzrgdcEg4wPtxiruqu9hKfyro22btyuQv9
scNXONzt+bex0UFdtUyTnmUtbKyBLTjfkAD118WOb9x3K2AHA54AgcosMVLH
eHY6F2pqcc0yo6jhNBGIvbSVl/RXfJEC5JBv5Q9aOXAuvcxONAPzsFPdOIao
wI/ghC83sVrkzRA7vlQYk85KQFTnuHij0ad6rUrYlLmdBlDGrAI2PXmYkf92
0jGRpPInE2+LvCM3b0FfyBiWF6ETk7vze0iZsk77ZKpaQplPSufFVpEv6vYS
qkNrANzMsYOcVDXKE1jOunTAcFzsOcXXLY07TxbeXhO04E+E38yNxdF241qo
3vaBYs9NOQsm885Ff/5wAcNbYD9gZAvddIim+hORyf0gtHKwahL/7yExkt9H
O33OC4APKbJoRe3EcARIbXk6hjhRnbf/rtIoGVRs6+vOpNkOF6GEh5EP1l0P
/dY2RDQXCL6NLiTzZqRxAXEyvOYtUAQH0TCUtQyUj3ORdS7Jjq1qtjhruETO
SQ1jencZlvAfgItvcKYqj3VaQAfGNTNsVfAD2QFc973TRESXFJWsEbfJza35
0C5GtXDyd6V3qsYjdk/itiiG1geSs1FNyWxmql/H8o19g/BXpSoDfKVp0w9r
Xw5zcBf5Vqw6eBBYK2loqQuFnp2O1p1H4YOyuFS8dJwawkGnP8cc/DQqg44n
ueY+2/8jbdySgnjqdVm9NSj5TpLiHaXNjWqihid2yLB7ZMJWf1ujlPH3h/Rh
Ms149Vukxi6efwJR3NLQMnaEZqOaUN89bH9+4OS4PNAz3z0v+QvetbGpadRz
hno2JfArQVzlfI3Ri/F3LyERjQvP8vkYwGUMwaABXtON5dw0U2f6oeSWXjzn
sQxaZbk+n+6Q+HgfeT+vePXjLJ/oEkUrYHW+nLlpxtIZOxuvdb6JH31ZNGCr
TeuFMEJC5zb6QeIoezSIVnxkeRWo8uyyPDKfH9GANPe94f1yHCGR72mc0S/g
MmsLBNJ8EEoCe7dkzHixYCMtT2sO7zPIGvIzE9t1/D9dIjQnpKeKhzYcHxYk
g4/OgjaxQDjXwMiCoJT9iX02owOcRnlYNAb6VbEK48Wosck5GMWIqzHtUe2M
qWyTRfG/UZdn/WdWdWFl5KFYMNNtPrOXnhWv0QuDaWNAeplFxlW19Lx8ZAUM
ECSh2GsNcrF1px3iYPVy3utFAGZlEk8P2toiQgW0WyL63D7oLr7852awcwCb
l6+mMcJ6WugBa4mVo7OK6ZstwBC/ZXc+htyJfi/4wq5estNRGt1Mko8We/hg
7UX3TBYwCAZopBlOQxe1NQi/k//pJ+beXdLvh2XHOP9XX3sQDIN/q9zFWxmW
LPVxNj+GzGi3t2y/A4620vfFvnsnxF7c/iuicjT9x6BLem6Y0z0cQv5NgKUI
8oZI3MTCA0X2FIcoi2i/hTcI1j74YIaOMfPlENrhJz3I+gyUsyi4ROSMhKZR
33VW37L790M+/sBl0AePmmREhywP5DlUvvLvV951kbRf9AOmTj4UbMe8v0ZG
DCEaoX73wowQ2tXiVqkdsEDv9usJ+iF7S2T39E87er+ZH1JtFTom5cGwOYeP
APchudzIgEndFElTf0+XOMsNcBiMSRDdCLkJPDgsqEPpwMRiddkn9XzL1iKc
Ix4cgZ4eB3YOiBsAvDIGyhx071i5KaqGQvamRPjRSZzHBBh0P7IyYw1krofb
tT6Zc/e4O7B2Bh7KSQD6VlH5Eyh97FV/xPR//tbOSD+mcc31dtMfJyEYraSH
QJ/vZhjYu+RXcKROrWYgvPyI0XePn95/oKl4ik75rMNMNEZvAo+dOCriLnDs
2eS7IX6hj4jTrlQ6r5OEaegzk1iod1Ir/HnyyX0QO1/JtcbOh0y6kP1twnt3
DQWLWTMuaYhJw77ACW3ZUMduR2vgrGYFYpEf9dMZ17PDZZi/sm0YvelKnmmY
u7V41R6qiDrCqK5IPNvANtQVz1NPuKpMY22j7ArXJVxYDvzGPpR6/b0hXB0G
jXq6Ui6SSMeVRg8x9/l1nJpYq9bLONgYe6CXARzZbS2gZTSeFT54IGWDGMI7
/VylDMxWN+R/MHYeH2yabkG7YCsYyvwd6XIKthH2zvzBFu3X7qjBbDxkXmF9
kQvjOmo0/ESCq04KQp4zN1xliiwk6eTk21POyL8F80XjCXOVvCha1YBU5/KZ
XP0Y0gQbixYPgHHPCmUCWZ9yjBLfwX9I9ZbonULdhkAbo+quvJc7Nq86fgKu
ZAE60Y62luA3dNVpro92QjK9ubmdRonYqVAhvVOTBlrNm9Jsfh0H2uJ23DU+
0Jv2/0xmT2x/xNMdOhtMgYYUE9MvkW7ZCkq9fOEFv5IA+68H6jQ4hisL5TIN
O8hbukLESjmuHI3qH6oV3sQNtCxfURB7MRqwRXr87sIgwoP2A80siLavjOcW
xwppUlk8Sh3n+5HBjDtApdUxZRSd6NW6DM6OKGdBI3wzqUjWnJE17IryTDdP
XBjf/BaeuxBcxfavZOZ1CKWRZVPlCIhdNZOxw77mIdnLgyfGGDZ5OO5ZbbS4
FV5aKJSOC6vYk3K3wNcqIDdHBKv8BZ+ofeDRVwqbcw7Lqvj4x7MuOs2DJ0Kh
jXy3XOqfiAIRFX87c2WtuLxzBeaIh0XL7IJO2YFXI6c1obRqCbOCFZGbsd3H
imsjlISqpNVMKjklKSxQ5l0I9e+S1ar8Bsci1e2jXz6RKbwi9sGkET1OvKpR
alHna+4LnECODoAckCyzzEDcuqg/oP3VXsJfQ7YrRbpfCmL0jAXMSOuwXS/B
VExABX/8e5yRsxbyeVKnameL1p0Dy0PqCSXXLSPTx4Co3vfackGrc3ru5mMN
0H7pIfOxqR0EQ2XXWRRTc9xJWIdTspb8I1SbdEsbMUjGfWDjVTMa1lcWRmDh
paZu8FaSoWS6e0iH7eTaTptlhGkfVQ/qSNV/iVEvPlp0nGLhgQEtRlVGfICA
K8QjX1a74gf11xlmWpVeo51bVOLyI5lqOZu+6glwwFFwV+CBmtGPoAQiZYUD
hoj+FJNh/xNvi6pHecYmJlsZhtQROSMWD79VxxzEJUJgYDmhvXEUYA1imwok
v3DaPkPhh55XF6LzkW+mF2+LGXCncikozNcHwLwoq/7hkGOdQ/jhr8kUo3Nm
dYqeIugjdAFZqFaXyvjL0GEOWXUDy1uOPiULl3AGz+0vgjHUoJz2upNR5lmg
6jg6MSH713hOhhDT+o4PxcRF91kjgwdSB93j8ebBj/9qBLwjkC0KBb0nKUoR
+BizVCM+JHGw1qmbmOElIYfJtCNirDo6GQgqqZ+6NclOeG6znAg8ysKstPpA
Z1gRLTJU2pHlw9/wLc5+trTDIR3gMwZ2MNUKPOdo/ZPDsZrd+IwCBS8wJL37
MxJYuoPzCf9fmesT557/MN6bT97aNtoxCT7xlI4FDefwX0a+62JVecbniMBF
vmOkRwEhrEGACEEEHOXQq1NkeAmcN4w+67tiqUqqMqIPsxULg/XbcOuPQk2N
33mJNep+vIOR60GQVrRJ6mYqSq+RHWtVSMrAJk7DIV/nRr6ql0p7gaOoLCrZ
S/y2tQgSyeGXwzw/A9LD65nd2C9H8bhgtlj+INnb/U6juWNSoGKTMjVPsa9m
511Rob+k2pvZOwnlbAP5JPcFx6dOO6Bj/2mGWCca9zSltwRRnOg+9gPbTrSL
B9gDixCWIpXP3A2D05+dA7Wo3Kwej0XOSeXM5aCok/UIvcnAacO6/Qq4MLVC
1Q0lsnK8zkwXMfa2h0Ob/foF5rtfemkjc38CFozjZb70fvTOKk0EPBBWf4FY
cqFZnCpiwbgO4Zq3nmQ1+/+Nh+Qn4eAOOeDYw0tkcXaVykzbTbFRfPsXB9rF
qn57a0ZSqf3V6Kcow3H3MnZNtyJoo2MkdJDAGKmBsEbVGldivfPuzm3dv+ml
wLPDPyDkJYqy3mof4/iLNuqLWra8gdlgur9iICGtpGJ0aJ04RzmMiab7jRc9
VzH0zOpfBrFfKpXUoxVRi9/PZ4O8xvuxvgPqRyZcqhMy2HjHQ1ZRsc2yVbi4
ZNxP46v3hGfROvOEbzRwZUWNH9gDvi7tg7loIFqHqRPCYPB6zkQn7l2iLOq9
oxNvpmL2MzBeFmCd9eXCtws8oCyPdp95O/U9fCuu3gsMeB1gWvf6/rksxSJ8
/vkR9n2H7EE2aomg4jRqKlh7s/fF+9XGbSWcoO0Gh1WMM9B6ZHNErLbvkufn
IpO+aVawVC34DJcOaS1NjyoBrwsHJSBjcqXX76jROnXyLrm9JSDtP+Cbe4rx
1OfVGhJ+rBpQPsaf6SbN+PjaUYK835ZSk7aTtUoQ2jYuO/V6MZXj7sfQpfXu
hNfBZJQ4ARz/uIi/IXDhLNPkc2F/2qH0NHJbR11ur+LZr2O5uGhEj/U9ddm1
ZQNE3xLvM4sqLFkkueBnDeiqXfrC0iRO3RArn8l2wi7w39AJuX2yWooLd1zj
jYT6rvVWTYZeihm8ndx2gu3SLCsvt/lIBh0SHsda6O/6M4dr4VwFyBfRyVbB
8vprQq+lVqRRagzYjVzLvyOmm0cm0tv7QUoZniLV/9kpffH+u1wwFECG+KCs
JH5bRJLYGQTCF42uJiWUUe7WeT41Npwy9KKczQf4pv4lsGsThZMDsAaFJdFS
Nkj5okG6h/6ThOBOLiMZlYf0N2yVhvuFxaE7ZA1fHXn10ZnMXbsNu3H3wxZ5
uoKTJ9xAh03K/TRojlazKPE/nStzsb7Y4gircRkB+WbwD6Xns1S2ih+rw9zM
WCRaZMbubzZysDfN7T5CjvvjXpqFCkKmvWwUjVU4hdoeNn2uuGgtAoSQQg8H
pRNiKMs12+AUqOpZ0SH+Wq4+YW6trlx/8hSoXU+0JPHuPJtT//eXFShooL6H
IV5miWlRSZScTYT8Q2atKAdEK1/sNsD6/hCHnILISuLWT+9w33QDiqHHB7je
Xar6YepvuY3PvtONfUoxqMUAmGFTd/GQc+Y1B9fcWJrou8EkbBvsYi6jky1h
+KJYN9Yadq9m6LQI0cC+S771JS2V0mQmTaMPbRnHaESPejMhlt8v60fslkUT
B7qyhQi+V5Yy1JY9zqHNqKEUl2eML+DX4GYpG+73e2A72aFS/uzzvLpgzNBj
pAykyjZZXX2wvd51jARRJEXzbfu9GZnVGRU/g1JEzOJlARGtXbeBnLO6LXKE
Qu86U3LmD//EjkR595sZBEuv4F5IaC2EjQPuyezNRWiY4oYiLcWUMmNPxccv
nGO5NWDxSOLI5xTtsmp2+Q+Zloiccu3RNUyx23WEe8iqrP094+Us1EpoU0IM
ocV4KaXw25wxl/W/yqMFKI7V0K5D24GywZAD8I2Vkntduj1vFfjHJP8LeOfN
OvGac/JK3yDrTDpeTJEFUdtiPkG7dAK+bfiwxXKBfv6fmkFmr71Yl28o+yY9
YaeA6y1IJRYsoefOiLQqUz6vpg3zJXS6gBYy+PBls4GVjKFCBn3VZujItHEo
hIfyRfFxkvFFZIfvwQM7JUdhXbe4dzc2f/IIbrYhKt7+lDoWIK01Kupj738O
eKRpPxb0/JfzkmpR6N1CVzyC0DDeiFJ44vXOtumWT2dTu/BUOABK3EF00Wxf
dP9+MV1/0nt1SEn95AJpZ8kpaItbMGzdwZOA+YZGsxsAfVD8yYSX8R8vQjN2
qDr3DJLCFYHqS5nP/aaM9KLZKnNv8A2+Xe2+4cmheNI2XK54CDkgdyrM3wIz
gE7sfPunh5gJBaUlew/PRa+UH0YHirbb7/BsBfizIGbZRr7eu4v85/9EiVJa
XHP6SUlWPH5zZLXXIidkstrrUClFnPLtaqzWd9N9cJucI63dk3Dt/afWi7tS
6sJ2nVkNTy3Fomx/2njZMWU08jryX6DzG2nYGCVaG5xq/ExSD0IjOE2xxoOl
UW5b611WPL4oVTurL88sx5DWZhphfoDpH197N1BuIR5xkuQ94jyTgE9t9ZRy
dy2p4KV985DxgUkysCNxs6YcaVX0D7zW1Q3FpuTB0N6qSjP8hoVDDAhYmmAa
dQGwTVtPJN3zjGL7rFUsczFherdKEOVWWBRdx1u3HxWDw3g9Vd3yH7iegDkY
lxlZWuyWmp+3M1TNQ8bAPUGNVWpjy0DNG/z7ogo01/86LQeXErxXuuSXMuh9
IpxQGAuFcv3SdM/yzaxBWOZ+VaEv454fznXh1R5nnifMt0n0K57Z0v765EJW
bGpkvAnzmrNseFjkq+xsf8pmL8GqPjat3dRor1fCOXMANnNZhyFRS+AaGemu
XCu1KyWJFFZjUYxRmpeo2HRAn3vyeE6Aq7HdfZFYq17JSSUXR786aGIdXAVo
NMgn/AtBVWreqAsnwAz/NIrIDMeVymYbFOY6TmZ3rPdv9z7n14w+1Zdy745O
s98LdZbe5qCLt2ufypBLLsghSJG6J11SI0XJ/SNhRJKHCO7DR4cY5eXFlnN8
pFOSU0e0o0iazKKuVmIxD9AKOOHA0+zqW6eJttKaGoa8x9sJfnYvUKIaMIba
Z+Ibi74KPx9RLQSt2AqsFsO/7jjNMVjheC9qSWB6J1FtG9hekW8jRkdOuEsz
LrG2bntUmUqvmnO5qe9NPIKlNxqbyTxWrrFo89XeQJaM9ueboQcs3vP5LZPv
oBtdbtjv6HMZKc/L1a1G75ii5eD8CW7b+nRDfqFF6SkYSpYOB3tsg2ypnlQF
u09DE+iUp8yKTWm+q3ZlugAHYevjs4rv8WsZ03XbuyowuNuXs5NErlr0vV1f
c/lB/ekFBO4In4ZRpt5sEFWY9iOjnm3lQXx0g8Fzx3Wi2cHQs/n2ALCL3MzU
eNObLzVHrucQnJVVYN8+rdOXfntKgxEAyPISRF2y0+BLU4RiVBSIjrvXgije
fdcLlLYcdqbdWaSli44eXFKq04o3PZAlOOY/QKGkBNFU7dLQa8Kx62dR9/Du
wcS7crRswSVPcZy94cY3cdc75P1ydyyY8LD7nRUYQKlBRndNto/Vz89xXBVB
9+08tSVJUVes2iFvxh3IH1IElE1yNhTacGPZQC+arHNZdaz1doI+SDTqJmjd
cfiMZGCtgPfst7EDA0/+jD7Dmkhc26A2pLb1CBLgIkZHFehatu6tDY+b1Xbu
XjSSSCblTSScc0k5Hzrqu3H70HpfUgY9xxcRUZje4E0kA9D9gN6M80ISmoNS
rsPi1pcVPhz4vlAlh0B6wnefNZUy7PxQq+pgjv7QyTtjGbk2PQhyEn/Fi+Ft
dptyPc8vLS3/10kyVaXVGTAUK6UQD1lGrdgfcEsRAdmle/g/QLOpQFv91Uwi
6sPJBcWIqD689vA67ejMIPcXqyRtzNZMR5fUR6onLHM/7aeOuO+Zff5w3S8L
c1lRP4HNqXWOlNKFgLsITdPwNy7dr23dd0AkbAhmT/5OA0lwgRZFefWwSBqN
huhXQcCzuPaZWQlC49GuDAe3yeMyoc/utQbuzWakLyJSq3dqAZC8iYDRfF0m
QP97fJbwx9xUZVNivb6bY/wVtMu7twT1SN0/tQ0chtonaIyy0OElA/4bXerJ
SgM3znb7oV1yYyL5cQtMIKx5ZFr8NNTZQAE4dg1FBrLvwQ46skfmtm+fMK7i
b6q2IbUOLA5EaUzDuOEfZr3XHSNyJf76PyUqt1vsqf7SJgmRHXkhmw0cdtNL
LvDgzBIK6JYePOYtieMQzvZmB2ocWXZ4xJStCDc8KRovizGXxeyOnh8Yw98/
zpbTDi6sx5+6+kzfDzK7j+3HuDP4MMz5WcYUTF6BSlr67s43w6B72RM3jUzH
m990js3iBm41hQtqy2gZfbxbq+Hroj0iVHa7h21gHpVnz9cXmFrCxQCaXkvH
/Br26qX3A7JPDp3xr/quOHKM9ZV5E2M7XGukCavo+BGomRyFphMximLQTqJ1
tlIDBAbydrozdoUVOsMLh+o74guViXnj6iECguSAa2bJE7gzCfqIygw3uVth
7YBEcM1Qq+bIvAbJ0jbmZGEtH1C9tedj3kqji5+tRZHbz6OHdyWhtW/vAesd
G6sKqhL4+//hbDo1d2OcPgODrwC+45tRFXEbrC5Clni1l7i2GwHMrpcymmGu
Su66zr7lIofAfuhNl1Z/nf7mQdFr6+Yk/A8ou0cQwY/qpOA2YHRg0xnJeqXF
mrwJkZSrKxXnTRMFsA1N0pIgbmc8pTomcY2rWUd7U9d4tLO4CMZ4agel9DlV
yra6vhV37Mqp1ICJfN/93WZfy6fu2KJYnyDl6PteMVhtEFLVApAHUd2GV4+N
iqQw/lL6Btf5LCOHTwd0RzMjZOD+XtV9KEm+HOccC0WRMkuVXDXpbr9SXakM
kSQVw7zZWYYPqB3fJjmZECMvkN+qAUAjS4GcVrIZ594iNvoanMJXduK7QRGr
j6mvM0ovSxbAZoAC0xxVRzZukl/ZX7lmqOC4hl44ezFIRLpMupVSoD4FkYFG
OrNKCRTxa94jB433sILwaEMoQmMPIYyrTrM2rZx+Z1tarjTXOv8oVEbSYkjB
R4OxalDuP+bVuH6exQ6Olf0sr+KYr7l3OFHDO74hEV43nCxbWCQVGVH4PsRT
/vf+vH0I5AeHCs0OI/rvoXX3qJmxypYrVBNLPY4ipSb3zKqc0dcBb6Y7EGFP
NGznJrZA7uSVT9LIM+TnYpifDT8cgRZE/sVdd3AN3u3SxKfQF+pyOEWFDv3H
ZVeJ9EWckVaSaDeCVuCsMGlE/ZafThIfBttb+SclRjnbDy37cZU1Blo6t8ZX
JnQbwaXPURi8Adj+N2EVYMcjYmkvGG7OgSHkDHqISQ1mEw3UgehM7E5ASVYk
IhUqQAfGom+3uTYG4xuNkeihHlJrkGvWjaEHdEYS89X4VaEBeYClPsPAZTgM
2NJOGCOb/vMwmetq/m8hx+MXp96y5JHM3NJ1ulA1/wyRd2fvSIRXCjGAW7Ny
N4+YLQH9eLtyN6bkgW+5oXb4g8raXFsQ3VoD+v5uy2vMNnyoCTn3yyvJZP/l
O6k2zMs7DB/JTBnGBiQDV1f5F22QdomHkawDOF3o4oFGNCLUmpyQDaXSK5Z0
X4ULqJahk6aRhrd1Brwix+xfVMH8IaRUOtLMtVH1YsXyuAAvTPli3d2GAYjn
a/mqHSAu5zwiw0OnXgEx3Ol1HIaXiPKGDK/V6l2t4doW2FWVrJKBO2I2cjrV
kQoJO8M1n+7UUhmNDgz4oD0v8B0LpRXfvqetoNSUmuTJaBY/bVEuQl+PUSHH
4LbgR6heoUqA6B8nNMeBVggakdA5gMz74pbIqTvk3W+dhyEk9/suOI50O4bH
PLTOgnUJOwzHlZmggTGPTXyZDXWtAMj6FarTj/TlyxRqY6pM+pJtZlrOUseL
hPeHlY9xqETpYBgWfXmo2GE9hvEmMQZUZPZu3G8a5KrDyN2Fzb1ugIj5KMoD
cxjpHvBUnbkv8mdAxFjscYTzshwXrXFQeucGW/3vfc5H4StETHuKHYmpsR57
XXA9O6Qy/VRgZtESTH+pf6Tex0IAqrOQk2shYhVgWMb7JhFDb7pLBAafW0bm
b+zqtar1FbC4MbRC1MZKUSHYShDvaL1Q+cmjuwrEHdCPR2qp8zsMPRgBb/tr
cwHEST4RDGRQZzJTTevkyTPSVIFjASxSbhr3oguvanSYETv4VS6jYBt/OeD0
NzR57Kpsf9KtilH8UXLyYBLA2zKmxmgAWqqcRItHYFtPisDfurM9uDbsuElQ
ItGs4TcX/cLBwQfmoNnjxZQd6krBQOFE+0BY9jTOkI5CO0E+SxVUwmSvAgZs
CgSQUaMbWlaWiJMiGjAXOsVdchzy06a5SobmRlXfdXJAG/eKFurs+dpzhAAe
wd9A86Z4NBj4quEda6AJkNyog4lFAn+Jx2Zz1E+qvOboUw4009OAF2zgGkVX
I6mjmKTqv3tt9vdtqKfKmQWZbh0AjG2zbfejFnhIchqPpDvfCFqdKq3x7FaE
fJqzvjb6s9z+IZ9+g3finiW50l+mh9YfP27vfcvUjTtcPJ+/BV3fbMnEUea4
xcWTQjnvTWO0cO6sMCF4PzK+9e0totfOqTfzkxKuuJaQ25MnkSwQL3YzBXI/
ze4q71aM/xPtdtGizhW5bnrkCGI4nOcPC/7U6el29d1QblmzNI76D3HfakYk
pFSGStZ+eCY3bpLgTRmH/vDq5+JS+FxA0TWvjpKKL+Izx8G08b7fn96uhqqP
5QI2EYXq0hsWKov7ML/TJk+XUHbFytB6wDHL51lM3uYEX2JGPe0mpE5mCxqX
89wy3IJmjgtxFK0coQHRfW5deciO40PhamdXt59Bc9q9IM8NYN9wv8hHQpzn
hm+5K3elfkahVWryY4WYHBcL8zOb8iS8WxoVKfp/6bMYqlFkVEp1U/hWqMKH
OQzpul964UrbMSnkobrBlON5X3chHvooFtgAENkdkKi2dlPsn/5+PdtxXCbB
RT9DebdVsgjm5tFdXCLvmfU2KgOR06sh1/ZUp9BCXiS2csEjzhbSC+g5A98D
ZfZJrPF8J6Awvey1cUD3u6OP7WfCAlyG5y/8TFxxRqHW1IgQU/K1nwQwrduy
Di3S5FQlC5gFyWkcOwkX7TyRRYCSc/algMof7edSXIoaogIffwAwCdVuCXlc
ewwrylC/xTTY1RPkE+eU806mAPLB3eMPT2vtcNtQyx4Z4jNuhWXnI1LzVGMQ
u7xqRTy+QggE76/6EVX1ir2NwrUVYr8/QVvtivAzk1eVn/1QRzaGdYS7XH+Y
9fPiqn0Wmb3fBsvnc6UJhDH0dvoIi+U6SmTqVdkzma9XtpylNkI2ZTJXUJWo
n91fPwJIWP71LPYnSXKrajGxe6SEiKRixxcW2cvr+2rURxiC7DamHxQc/wJG
Jb3c3wvF/thdEK2tSJUuyM0i6rX28RM77H8aC0P/F8go4DnhRMxD6zj3cRjt
5FjWFvSKMCCWredRehIcjJGG01RZ+INIHFNqQt4hSovYl3DhRGhTVDwYaV2v
P0I7/xojBUSLaMVG44l4nYnQz14zQ0ERyETI5eMrRsAJtui7/DERoQGpR4rY
Xw+2gLNp2a6j4PD/q7EnrgPFP1X0KwmkL9TJ1MfsAE78pRv6NQS15GTGNVxm
2OS7ygueLG7N9DMgGnZfbmk8ZDQv/PB/5u8bsyWNVSWboOwKc4KXgCGif34P
Irp5VewyYf4u/lvILqrrK7+pn+ojolCDmFkcL47uCZmuZGelmOJ8+jM9Yf0Q
UJW0IaQcukqYq3plOs27uYzq1t/2h0o3vGmDaFYOaL4VeJQXd3kLFnq8PFf0
r0azRHCidMXsC4Aa4BuMymx1AHT0yLZKUnTUttzJLdJgAPEroqL2UFv5odIf
gG9idTnEsHraNQOI1fpgRodhCLaQ46Jup0o77wmgVFmCImIEROGmqfeROy0o
KIYDkSeID6ArFDB/Fyzx80RGtSfs82MxGqt6k0FnIxk5PPhyEM7me+J2qbgx
ysaYTsgoLwC4DSv2pjUSN7+yIUn9kzVFO6+wkRLVwqSzR6RJLzH4YxPdz/Z8
IPtklDR9PUn+VneDXrRKdRGMUb+DMp1oobI9Zf0MIHwp+v5G5bhvlRI6Yj/L
vq0WkMhmNXg2TsgfrNQAaZnBYlm//Gi0GhFbpvkcfD0ky2YIbnk3q9VfdJpH
7uDGh90FUSgP8dfS2ZO4N+NBNKwjveJfhkul1/NDHpCxl38etAuF8LBcg8GJ
N0qVUIyK7BVZ1fhHmpmZe0WY3138IKsptC4/QgjwzkhBFsCktki2d0f4VWmB
negBRFHfHKHlny+F+kHk7bCjh4XzlU6JdrVbrqyfTKhqlnc666oafmWGRI3Q
yxIdNhN8RLc5Css0i5PgaWxWr34sNGv4LwRNn/AxjADP/gNir8hVmd67kfLL
LArbHZ+PYJKaFSwtxu1sToSlLp9Va4OJ5Y7LB8G+PISFjkcIebVM5HyrEwsS
1TQFrKuzBcYKkeXvxHSYuMWvc++GsH+Bk4CiOXGi0GZywn79e9mGGiBY+t3A
QdyNmGjYlBrHNXA9dt2y8zIpAd7ZHZBqjnLKRLHmBnBBL5OBipwtNMuH/dpt
zMFbrap20quHgtGDHdtk5S0zmGVkt09MoFmIhc1OP5wRb0vibdwFAZU2Tk3i
n5VtI+fXxyfcPtfsnyko8rxLs5TjrpZY0XXm69dVRL0Lt9BPXV/5RI5r7/Ec
xnf8es+QTkOXafBJ2LdFel+xFiOqOYdoBQDFZIB80WD4xtgTObOrA+4Z54Hn
6UQSpHjZ/DYOQHwUcvLpD98eHBE7nMEApqQaYs42rzmn7fh50Bph9FTY5ZTm
KiFDF30mOElvn19P1wbBOiBfDygnhDVmw67MmjZSEC3lPTS2lp2ioc6JAiYW
fK720j+c7m57IHstq1qA5PugTzbYhHLmbVbPUJn2dcmLjnvK3WpZTulw/xWO
j6RNoN2LQrFYnNAVk7+nANk7//tRJdHa5kg7lwaZ349+0j5lgVdGxB4oH7I9
QMF7ldaHmSReXvPuIuwB/SyAOHups4J2wmcyAc9B/aNnJlrYQtuES2qrw/RA
Ozm3Gu0VMcob0JeQGmC5Fd21EKlAEUjWWXGrwRJ3fHpMFqF2gbeJoh8rSRlP
LzxwQEIJoPqlapKRpoNHgBPknIA2VRrmNZf88DoVggs/WVVT1HjPwG6WzoSx
JOcTfherAouAOuQPSfU79zJB7mYMLj8haE1J46l05A8jMAFbf3hHhMAUmBKR
+AsBWGWQXjbKykjxlWcNIQLzV/Nuxs98VhQqLvBgqMqQ0gYLW5G98Si1gFJ/
qvrXVo8aNsD2znUY3dAPKOBRb7PtSM4YNwDJi9CNiUbGVX68gMxts7Bd0qoh
7pkwKXnkCQR3x+2i/1MlPY1QfyB4LpAnwMwF/tFcwQ/fAvETrOLoImgrLh2I
0/uqZYXcrmHO/9MNtSkaoFcjfoUQ0viDH5HTmPdFebiqoByQ8GKcNdOzT+l/
YzSTGT5j+CbGz65x/m2ah16Am9Q+yt5gTG2+pQ+V3U7YZAjvy9OM7y9qhZHT
9BFNWxDWyNYeQalrfZvLJTplLnukgLmHUKEQWgNw3V37SlmcQAnWfRej2aEI
l0JIs46L47GNfyceF8NmJh4IlcCYck3fT7VSLIQE7+v2MxmKU4CeTMMgj88Y
/AiL4cA07qxsdW444JSIE8z1n4MhSRdVPoZSxM1ellwVnujIXFZf2pkcv3Be
AGZmqzBeVshLGgzQc/DjkeA6SBktMfIXmZH/tEOaOBuh34x+hC6AjLV+aTDQ
/TCeYEWaJFpF39iLCi7NR/9DyFeDDCSAWH+GTOh4xpX6d9IFUX9fxNghWtC+
COU8TSoMLalyugmyfelaMhzixQFtwgCzPLqcTK6LwZA0A8gq4x+yuZGfe/+i
Z4hT5HV8ysctJBKYRe2zLURapisUxXV4TvopAOECutJwws0A0GsLuIa0hG9P
tM/YugXBSAflKx/Z6M5PG0QH9qDy7o2yb4QbKH7+KRcL4nECvjB4iX39SxaQ
TMjV99La4X3QzzvX642f9gMOy6i4XlDLfyvtjeLVM1YFrjO25TX+REzXDRv1
4YOZ5Dao6/IQQXxAuo0e0p+N+TFjoq8up0mHD3ZGkv8EDJaEFAS4CrczCKP8
I/sFNZLRcKc4eyuwjKyR3CtL47k5czfIxKwiI4uwyDlVuqNcFqmPKDJ94Wy7
b7nzPHdclbkLQXgUQMB3DaRjJM6Nz6rGqv01k56qfUiIq7s4Rj3lOE66tACl
DEn8RbhRlWpqTmO3gCLkWbUpu7sCfTtlL0/fPF6MLs0Rb3H2k+SxC4wk6Zsc
hEVTFGs8c8Mm5E4DHsiG6T1U2BXCcNHmQWo2P/3eUHza5oRZPeWTZ11Ud/iV
+VtQmy6wIGaJZ7CZH165pxgzdLYIDB5GGMKo12HYRj5F+J4r7vQ4WuMMGVW+
rQhp2OzXle2AaIxjbYxesmbbmLLbNXlKNaNn7T4QzJA/Y9AcigxgKz6iQl9w
ufrU5JytAknDyW+txn7Bt3cr6yUtIdCqhgcK+T444rSGkeHyGfjFZraa9yx8
CaATC02hWlpP0CWfOIaZH+fXI4EHkjxsvsRa0ptNTBzNrrArcMoYf3Oi0icP
B/ohozhu0/SMq0HPAbZ677DcFtQoxXO2G9vd5xgRHLuI+sDvl6QbYVCvDcia
MnP8N802Xny/KPxyKQ75ICXpXfTlWKXbqbZqNgFOI7Wtg6fiwRmbY/Xykndh
VwIQq7nWHKwBKPFCnZlvr1QqbE5L2dmdEiTAJptS+tDhKyt2SrH2vP6uyaCG
oqGjRVIHcuceHIobZGrehWbSW5Y5vxVSYibq6I2D4XKFDjeM8N1gVP303/Sv
DL9kt88qJ9Kweb6UTZ2BCuCJ4MCfT7JlIKfrrDe7ChRmRtaHML4rXJhqvy9m
G4Gt2CihBtFOnch5TvYgdfHw45cOsFfWkQh5k/LCHzeLTd+Tl7nHgsWedPmV
oA4/HLMIht2tABXWdtq+p71bfcj+dZOGBAEqMFBh7Zl5OFnrJZDP2uyjod9N
pVxklBqp8XddSOHdHN9XzI+R7hmUp9Rdi8vzTEkT3d+oYCkZfz4CUm+A/nt/
/8iByY2S5PaxgUYp4496HiLVDZ3c5gOtvdoCSLv5ouDTDAsywrELPxpuz2z6
UfzSRDC5bB6VOYLYn/U7R7f0ZwQhvGxhUThaAWv9JxmYX4m6rz25ZgaQZOLT
0LL5VuGhpq0gm4M8cdcX+pLa1H+NU5sAsyNWf3GeNzDrwK9Y9dAvBF+IupbY
4UNrlUiRwwGAhWUALy2QqylwEr8evia1N9yKdNNAow1t6U1AUeiXXDC3PR4Q
mJmrYHzrxAs2nby+tclPwcDzmZQ4dmOgiSn60OCtkeHYxJjdpDbF3oHA2sPq
tKcUeV2PPX5Bz/Axg4iQo2+cicSaVewjHI2jqgQzOZij1flWeXAF5ztG37As
iU15/u81SffV9F7VmpdLbTNE900P/2VvZJjn+hRBKtUPIJpuJKNtTE0Ixjxn
pNt0fOf/CNTbC92x4nyxdLK1Op6rg7DyYhtmAI3JgExFLD3vCPqM/dsE87Sq
4n+Ho+ZD7U62cdBDaXYtnwjO+UaF7UkSo//AICllM/Qkd7WeC5wGTtDgOpqJ
Rb7W0Ql9DHyavkVCqD2asVkP1GuaWb1H9BMzw5QzO83nxOqZFbUQPxM9MF7/
F9b8SYM/SKFHuODMHHBY9KqCpXizYlLl3Qi3WebYv2LPeMo8hQWv4RO/JB+v
HwSv0VGp9yDK5pB1ynM7YsttP43osAZ9qubKL+GDDfCvdg22rhjoNIJh2hrV
U0R8kMRDLGiqB9LA2hI0/t4rks+oAswFYidmWP4HXdFZObse8TnvpKggE2gx
h4a8Gqg7IN8blKGn6EUxg6A5Wk59MTumlOLecrCDm6J/5IwOc5258copKU9X
tzx50kK8N5DIQH0Er2Am3kPRSmfSyLAigwHNYFHhXfYCsDlCEKLNzfjVNgs0
ZvcZMt89yl4lveBiERozWU6QRy1hqvjTJKimkXx8rIumkU8KKRboPYrOuGMi
bL/8Oof1UxIn2t1k9scIirupLsfd7HrpgzdON2jY4TlFgq9xcRoFD0simCKe
EsuAJbDQE88LbkqEXoFTfnLYKiG4aYsqQHcRJGgMtokn76v/uieW6GV0k9pr
gtRaBZttccb+qDAQU0i+p3ZuktNALNDiaSPVQfQSid2MsrcBDBwxmt72hkgF
uXHOEOnnQuDmsqP+L0xuquNCX/2J+7B67oQPkl/SqwAvqPWh3gXZnfNUCdOr
m6FvCoV0Uch9rpeYCMZJgc2NWs+QNrnUjefvFyKP4J5f2hAWO70cetiZaZWQ
P1B63ng3pTbCwUlDSu87LLfOCZdWYeUcupfPQuXa0YfNnoS8B4ifkwWmfDsu
Xr56PpKfl3jQjRXT6wtfxBdrewierMbsOskMR+wGIAYg2n7ZBwEf1bRIBEdY
PFAPPTWwP/LgXqnxtFumgBcbCVEgVEzvwLph1j2JY8u4GYO6OuSoJmevfZJ8
MOVP8kuiBDB/DUgFAd8LGZlyouhGeF3f3SJfphHT8RIpEk73BG5pMSNYkrfl
mfIhDCaP2yrpRwuIcFjFp6y7ak1K/rhXZEOBANDojpJa+QI3tF98q53m1JMl
0LQmyREdiLwXgRQCotV+yGt1pokeH4afojhe+JYX+CruTnjufMLGDlbYKvC8
Hk4ZIihYxETejLCpl2BLHEdoBgwlb/YCf42uVmq1ln47HfKxylfXrgQ2FG3I
EUo4Ttd3dUlMJWegBavOe6fq4gCWf92uWHyP/sGmtkLEsfmTv2MAl+K0y5wd
MeA0+yNgDmPNq+xl7KQTbS6CQgj0yObpytSmoyZcYDRAvoz7/Q1srcJoC6gu
rsfzJw7qFgLBksWg5huZsFtfz6LKDGsMBwbtdUX4Dk6MX2fx4vWA4BlvPEGx
71SOWT967kWD1JNsoztvU3H5HErKsKBziraOyrmmiYJ9JO6U8gIUOqElbyHt
SW3jrGeA1GR3uOSc9nlwvwwKR5CDDlaxCaqCY2tfSlNPFyEGzReURrHAi9mx
XWiDRQcwu2ictGm7zeNTFVK9XgiAjbqm6iDEFcs1jFEsHsUItTQdLEP8kcg3
DFUMEiegWQOZyQDzVBRdeU+btpuO+PAaepSEOyyW2Sy5JrN80NJ4ELLajESV
tnM7duJsCnBP4+n/OtQ9EbAcebMBKolTBsbBWPYxR9rq2tX/DVflRA4JqEyw
TyBQf3bcWJOaD4Lg3Bwqnr7pkjDuHRBOlUANISiyzJ1nfgx6bfiUusbX2ysH
E4DiUzhTOMDL1UsUjubEu7RCWCiOGiKL+64o7Kpmi4+ANie9jJNkbYskMBtK
qUtvxYpuasRHgmnN33/gVD7RFLKmnRu6sIcOGPl7kdpVCC9DvCzXuD7vizX1
cn/ExeM9wtlFeqX3tg05pOkSxN7LvZU87D/av2IOnMisUaBn1rOEcDlLaOM7
lB95+N4/R+wKgu+sU4GKo9eg7b4JnsPAWVN+tDqxmr7bDUnUtPc1zPFbfHM4
Y/U1ypThOewB/otUUW3VBWlc+bgohwnTjHaIY57QUe0HnAOtQyLcI7MgcERi
mHAD7N3uXBlTFYfnIJN6mK7I3KzI+2DaK5PfWTSX+AP1OvkxBgMamiXFB6Qo
JstSnJ5R14qMcG/ehIuRFBBXVY+bYF/zRePzd2tqMlTHDp3KSyB03UJJUJHA
bNJxnJRuXzlPpNCA+BBnjNcLO4LJFJZCQkkcYCn5Oxrji+DJuJfM3c9nfja+
rqWMZIrjT8T0mQxICTUrXdNf0OWp95jKn2PPZ2OAG/i/2V6et2BXoVIBrfox
7TnzeP5gyB5z4/Bp5yRvvMj3mFB9r8pXn1sE+FjIGp7TLKHSadp/lPqZfgm8
n5nLVyYsjGPddC4bhP1vW/LzgDU3vgKyB5W0lvK86ss1TaYGvyZv8BCNRTEa
XxVbs4o5fAHqARvonkvqm485AE3Lva7VM9Ita1q6vZq3hExTJXl5RZBDt7T1
i5UBLa4EQxvTKD0fxJIXlV5lT+CTvFAyaJQHXfnUhYDivkxzv1u7Ila//R5i
OpZBmY7wqxauJ+ga5pVlCAlRuE4DVWgKVonJkGa6w27iIcap5acWtUlJkrnZ
vjrVtvtSxQCwwYWMl130LgT4vzE8oKUDAjp083ZFs/Wnmu0WL3Fhmg+xEW6W
dLZbOiYKjBq0JS0bgIxFOQcw6QTmGRTq3NMaKBRnPmzLYXcdbHd9u9NhUDaa
pXgKkUIP0LfKzQ6mOdE2t5sGaD9xwLqiwDcfYU3HEq2vCUmPh9j37e56+zoz
1j8qBkV+HcVZe7UKr43k7uVvRkebd8vDmqPtj9G19iQRz9JTzHwECwQi+JIP
B8YUJgLYf/8skY0rOfqVu9w9US2q7XoIxQs8RZBpss/wie7FdvDb/NHyi832
0yJ8KIX4As4HqA8ZCGNS76MJUYJK30aU3cHNfgUjQK8PxJiP8lIv+rqCuAGT
GNXXCyL3rki5AKgGBuwuHl2ugrtuQgZEhpxxk9h/bOC/SM3cs782nrV3E04H
sYjSNfu438pRxYDVw+/LC53Q7ZIZHYbF/1+UkpjoLobJ2JcBRDvypgv3N8AS
Lr2BC+sRda47qfIo5D/Z9k/+0ehD5ZUkoEQmopAa2LvkMNeMnqNFfZuwsEk1
jpuERIZaZfXWNBwn3qxZTb4cv1zQXdI5rqvzS3P27aHsrl7CiUlJutwVdTEM
bC9fDpxjJU/8WjzrnPqGSogza8JE3K9u+XyE3em/Zl0gXzN+jwOs7BcjFIze
c+zMc9JIBi+Lei/wO59DMuwdykZqq0T07MQQqx5/ARFQ3l8A58NogRoqhMiS
LBHTAE3Kp1PxsSjxG1AOztKc0OHyDklA77BaQ7XtF5EJ69UPJ7lB3/CdydMi
sYf51VD4lgp3GbmVAIrfXT+SIeCnebCSvFaiXbaKcww4Eb9THWWnu9hLFDj7
C7waiyHZqUp1PrRo2UN25uT5n6DoumKBgmJY3lyE2hSkr1x7+gVNkxqrVb8Y
PfG6ZN5Ksdikccrl3P3ZojLP8Erfnq1VgYEJPwGk3cUGCjVEJeojAJEl4lgv
3FMcFLKBSeV+6VDOiYiISPk0Cb7b3GtYe0im2IIqzhlJ5s0mVuSu4TNu2Adp
kLo0LiHSlSI9Tsm5pIQM3fEA0IPVIq8ocCw4plH2NkJtARaGvifevoB1xWDJ
1bp38y4Yy8jgSIO1Vjo3gaH7VSRuliNSZeDXdQXt+EhdAhtErTIwXR+CReFj
XTvD6iUlIz71yrKVRvIgDHkqthGkKdBf/yZLgoU6uKYy5haDXJkYecBRqSRD
LtNXv+yAe42DXZ+TbvGR+K6Dmg0BvEixjTCXj5Mmn2fyfLFHnJuFh2CT2MpL
E4sDrAWxjyTFslwQcvkjz/T7mwpu5r6dfwXwwhn0HO8cnDf/honsAiaPuF+C
VGw8o+h4TcBMez3Fc8tpqIHQL2iQ+7CiKkK1NIxTmIPPn24iLOuEFm2WX4Lf
F+jupPlorehNzCXvTxaHWu+NBMATxIWFavWjyCE64Kx3HuvYXeXq1eU3Tgca
4dcoi1xCOVaK5ZhOalUDQbjw6mhzN1IlGcafnuD9gPCSYdEMt3dyOcfx6htv
TT23RmvySSnCjvDEKbwrRf7bMfhsTocPgiTQ/133TYIpt4plMSj1VQewtp+t
SALhNSl7kvLe1kI8Yv1qM+1gBa6pt8ZbzPOQtPOmz1ziyQhHTFBPyolvsx1p
PBRXrOjQl9sUSFVS+TIbP4I7mbDSGRpXLk3Pnw0ZBATIoKHvay/stIv6edEl
CNW8Sk1Rb8s4myveY6AFETkIRHXKzdE0KU/AL52MZpCeDaKwICfdm/OPc5Wm
RyJTwEjXAWJ2tR3IrDFPGOXP2cKAqBWdAyuGcmdrX2FPDKT7SI+lGx5ypkf6
Pob3G84nZMqkh42DDMOUg/TIuW8HZL1gK3Y+oqATGgkih9GnGthHvU31zXPs
Ya1jzkzP+1bMxKqHLZxqb7lrKv06uyOeKZQkoA2D7qSPd/y5QJLvABOUUw9B
K2F/1waK4rxUviY7z8NjP+Yo5u1UN51E3DFOAGC0A6+DN0t1SjjUkA/7B8zm
GMoFiIdgzf9M3THJV/X/gYzrjYmuYgxHhKyP0Am5o6U+UIXM7kaqUweCHG7R
VvYzWG6XJYjGF53EKC0Ioj5oGXua5dJ7qqHcQU/Ar6o/3fTo5+Zj0ltKLH3l
9p1opOV/MRWZVqPpta26l+EZT8EEYbuTBBNjecFHZRIuXkqiiyuiOaxhJDyd
kmMuyMbIrA4hZ/MkiUu7Fy1EmuAIlP/GawXJxxc4Be3+2z77wlL5CKQkbafq
67j+ZwZ+HlhVpXdMUaO92FEWr2CzKldSA3krKPRjekvg59Ms6tkVIzICAKBo
AX3RPKg/+1E2PqbBZQNeV9PeV8url86aeCVEREtNGa7icHj71GhHt/hvpLWB
Lt2LLGtrBzxucW8MXCjvDHgMiig8vhaoYE9Ajfp3dFA2nvQY5LzgUs7IqLDx
VQnxLVx6cO6Ty1IDL9Nnom3S3jlrOcc3lLh5xiqoiig4LW49nfRcbcKawvya
x4yYZvwkhvq4offAKYZov+t4NZbdsK6CvfyxodrE7g3Lh6SQDAY8udvEw2nQ
4GooLDiAXmJ76eHM+knEGNCYmY2PyhWilpXXmCqtACXcLGMvXSJCT0ZSI7Tf
v+LuwHYA42SMhYSn8o+VgX0mChr+wqIS6JWJpWSe1mYIkKrvmcaSfHN8lqDh
MM6x7u37ZtT7MlaF3ZMcnOtB5AbvsyI4rKvS1pTQcAOofwaOKGYDcqa7UGMi
gYHdrbZy740HXVGKGtcexwDgIr2Md3/+ngFxXbvTZZJgCWSEcjxEdMM+99VS
DH4qHQBWRLbLTmwz5XW0QZ52l+a5bm+HskHeYEij0GNM2Loj/dJM3dMCT1JE
MkzPIzlHU44KTSLzssCvtEuxsxLwqVvJYjr6lWI9voBbJfxnavapWR4k3Q1m
ONhC3eQ4FVeTXC9wd86+VHs0ZSRZ82AU5B6ffiN4MWYHwWzwr4h4PzjpUdfQ
Zou7IP3gt4fCBNcudMVEaojT1tuHhf8IQ1WY3yi6eCOhBYTM5L8I5fdt0gxM
NWhSvqlFIE9fXWFUs1aBSpIJATVJXPCgKE9ft49EGxzKcWXh72NujJniFPn4
1upUe0z54sH332Zqt5c1yvTyAjZBCFxkF/DegglPzHf9Vdkuw6k53NKSnm7x
0Qh9s/0tf1coliPx6qsT2U8mpS3IpeEZvzvmxCEOHiaBZrYOYMwRSAxgWZhs
lsYjmlLdZtLrlvgkwBOI8nDRVZuLL0Jo0WnBtfWawGaf0BrlhuNjJ9vbF9rS
cK1A4M4ONylgVrIkIEYYrRn1YNy1pMVLVtY6RyVrEJRlA00do0oPNGXGL19X
0eJXRUIB5rwnxtRdB9zSBK0b1fBLUVcefkmN6+wAMHsVCzvrKdQbuzdORyar
UPeV33vZvfvYhSHe5+5WRbVhx+tmk3mD2RsNpYa/NKn9wzaMsY1Nk4Cf0iQt
4W2wUDeoentX0KnICYfBC0oSzKbiPIzc7PTI5EBnAZVPpW3U81UeIgzEmX8a
2RTDNZE+lQcxTGSMs2hBXIScb3/9AS9p6VoNUFLE45pgQH/d70eiDUO450cu
MA23GIgNOTYJb7/7o2R1Sdk73uIHdL22nMltwOmSJ8oMakqai5dLTnl1cX95
UCQaomvRTa1GX3i28LcaxZfzy+YLxW1mAFuKrkT2QmsS23ZZEQiCA/43mvX0
bKfcwoW73kFM7nUD/DzXMoE7JiVlOPJyi2RJe8oHGmC+dLAaX3KBfwa1XC2j
yoBXdkihyiklABgTKR6aPa5kpex7VpFuPnWiVKLCdO/jb3R9feGzFd3zeP/c
bRIeAdlI/djEr/QeBx9ClQab4eEpUI/wmt8+tKs9KAOTbKV/Fih3ZI+R38K/
hUo33N4N3BLkU0qoHFMIq7rykM/i2bvIbN2RGn0hpXFBD3cPXSpScRyF3CU+
nzXUyGH1kj1ZqDoua8AM7rDyffqwqME7ENt3hwZz8HfPTZBYUVdMPehlBIXp
cV8ikQCakHOTjtzMCac8cbExp1aC77t3CFLR04yy79inhqFsJAixBU3thH9h
ReOrvKwBeWSCdzaqdMy39oxS/qyYrInNf1uemKUjLFsRI5b2a2lmUvy84kQS
DyWYHo/aQMONgR4uu0qa0i8eH30o9ExatYJolLiu9QboSLB9sn6JxGZAZHoR
wI3JPcf+KahXQl9AnhBxhrWKgq5wvm3hLYwqLxUUvB8btGMmpQUpLsZcTr4m
nj1FzPhUxZSGOY8spddPKuSTDvzHSGiDRInT12Se+bexPJW/GUo/IG3+Q1Eh
JGRSpWGTxTudu82DWIfYxuLRYGAAe8d+GQFbu3RaljysfO2xBSTItKCGfpJ5
+VNGfnuO2qd7oGcjMjl60ZAqNUbsulTe7wAJNw6woSca+W0+gf2B/a7Qw6oM
EMFu7TF/TIdI57RtXXVDqxYZYtcsP9soj/BPa9Qrh1r9+ChXzcxbV9IY7uJ5
eYRf71Gjia4S0S12wLOW+Xg6NL5NEn0UfyQ15S6bqa0hes/dKXvLOJBzm/2X
ddDoIn1oOrxvL6WRUiM3bQ5HLR7HEknSQ+SFN0o2kJhRD0AsuI5fljAS6Gnq
1iUDFu/9IETIjKkOAl6MIp40GtNLoOjQ/SGFEjEMo7m6c4lW+G3RkINPehuH
gBhQ4eeZ0lTSC9VwVDE70qsaW9xHRGloCD1Sqy5QRmZ91NFQiZuyV7bcgvK5
NrgVNxQwz5v1LicfikJIiXnJpg2W6pgFDRw1Y4tHDkEqbmcTC2ID6CYS68pS
Hpjp+Wu1NLfwtec4Xwfiy9mZ8oqp/vCIZ2dQSK8+TOPQbDlsSFq6PMEjE7iz
he08KT5+fU4hNRLzkdAnGzxMZDMnJ/OU4YfHZP9srqn8Z4OOVQ8EB2psCoy9
Pg/IekDdlDttd93pFmNChC0Yc15kaMitDSCPGRN9tu1/uB/HmsMi/QU4xCDf
PpT/2hq/F1l3nJl3pAjS7B5Qk5o7zG+hIVGP9lV1dAyMP1GtK8Uy/7CQRLSP
iOEpQtMtFdyOsgqOyubTJzyP+KRqBPRwVQngob7AFQ/e3Og1ZFgYbb/jhb5E
jLxUNdaaW4k0xhgiTbOAlR1iUgOAn4cdkywn95j+WoZnQGg3dfChoIpZsGg9
X4rIVuCN5GMIBzgMBpMrSWveR2Q1nSKdkK1X1YqyM9ZHCzDvdB0rRKbEI6sG
AY/6MAr2Dxc6fIv+yht+/noW1SfeqXKgimfHQVUtxxkiNssxLGlYkvR+7zg/
rcBoXi3A/yZIVa5FZibJSiR5M2WvUWhFe+NreEWvRaevNcSbAR1tM9Dj48ZG
1USgtb5ChpHlorWm+i2XKMkoq5aqDKYj66pMbpc7gLD9wrVamfKKrdg0V1ND
SBgAz9XWrkhotzZQfV+kbd0OdeFpxQxMTz1C+Y6EFdpeowW3yTC5voo1dYXv
PotGKRiEfwis4BzXHdcY4R9y/cYBO4jNiUvTKBNcPQKh/I9zaG5DGm3FDFnD
B4aiVNa5FSygV0bzSgOZ3L+/5WYLbQSNHGMOM0jB6TRrqRQ0R/TzHdtwxcgp
d8he8bItVoWkMNiez4Nl/7FqTmqNspKe5tnVu5uvF46DG4KZczOGcE9djdel
qANMYVNRCX0EEELUqI8DDFR/cE9Atc1SsWLpL+wXaiRiQH+dodQSLY8ExFoA
g3GIcIVAVPDBNRNDEJwsuMHLGvDGsDApBdtdwKDggISgsr9cA30smLnDFLlt
e63P4LHqqujxmWtLqsWApiffi6ihrrayMRiP6PqZ2f2MNSJloBhyZg2ewFWE
RgmV0g6Cbj0EiA0WgnApHoXc2XkJcCaktzbWO2/55l06cqI5xZFbWbaDKwWm
VrxbUso4zSVfqBAhIN/MEL41ObRRsDt68GI8I8pKF6TSrt2xS8b4TVqoMmw7
hBpHLxMJ/M8A66N8Wkd7XKNrepUTGJuUwU8e5Q74Rk73Vy5HWaNpMCIPrKOT
yAAmJKCGGDP7r87H2Yx+qI/PXdJTRyZzGHow81tH6LL57YzbdkVSqspHLzl7
AEm5KONqx86DVhd2UJQVZxJcS5aQzxxlIB5RE14DE+y/59gVwr3UNkm/b7DP
KhkFScCz5Q+bJYSasGnDKcibxSII4MqlM/cxKPpmW+jHPTx28bb/zdejmJby
yMXlDDwrHEpXjo1uYscz00MAeIUeatOtbimnGQHGQviaDsBZ13qqZXsW0kZV
tD5L/mgC6PA1idfzvLKO1W+uMWLgcUVnuEiymGUNHGnqpWt0xYuE8rm6e2VY
DcYgQNnwnU1y+lbzieEW8piZ2Ln791qci/nOg7DDfoDvHjZwbX2mB2i9X50v
TOkruPxqaPYgnIIp4vZ33tWELJ7q1/q+Fj4WHhXYmokcHMaFI3ms6021/d16
jmQJHWWFblQ5cuOJeLRMmW48csjWZpK4fcmC7msA7U50GiNfY3D5v5Od0Vhg
SJgiS0n4Za5PlfQijc4U7z3W3hzxwgj3yF3auiRgVEFq3FCSrwBOwxDtLUva
aLkAoobj8zAbPUnrr8ql5jsIWC3qxIuxT9CT+WbNygrYNAf6wdWbA1aD5uo+
r6eMvNj/lDtldgkzk0QVQyXyjbPp7eaiEl8Qf7ZwFMV1rNtuv23OvNk1izH1
t2JkGfpq/kw6eV3BRyYfBw3zfUz1xu1XXD/EQwKxmIR82Db6UUk1wnDCbgqU
L6EcVMm48DSGG0v6aRonk6AfDVJgNefIEN6y4qGdgxiAaLfgyc4R5P5LDRN4
GqJR1NNq3P6l+v7z6T4RVTAJwXLx0QygIAgKb3Ro/gBa23AHOVeBpvv9ACSJ
XZ6cubBb4kBJDe9rx4t4cAlXhN59RxAxbkF+jHGwXFzSimhqWlwUF2RFyPvP
jSzJYssCIB7wY7VsDTcRnjLj/6K/rVOSbdqGoCmWmIpAyRxZ0MYuJJR54tFS
qOaOuGmO3FzmAGobuThNhsT9ZNLK3chdGrfKoyI/2TByJQWS75F7L/dmvZwU
kS8Pik7ABUisHG1WR2IJsAgafY3vQi+GNjfaCmPX5CCm3rXx9IIOFZoMFJzm
b0rP0GOOuDM2OGXHx5xC61WkLC0h3PP9p+PZ7jmca7bqsw9KAcDe08mFgxeP
j5Bn9Q+dXpnvbx90xmQ/aM5BdrJP8b+8fP/W8iZYdMu90Tt5Z5n2sDDXSzFP
y7ZCHxJrQi7dUpohQTXUeh4va5U/MAC5dk2pI7R/rLHsg7gUfZDK0vwNZD/n
q4sAp2iek7yYkF102IGg+B/OgpF6yB6liLSr9hjYUHs9YOow/agaMr9XGdr4
R+othxdRszpRqnsH6BFLiOxwoIsnl8Mzg2M4ceOuHUydgEeGHw2KLsfVnKZw
SO95khJ6Q66rb00myZkjQ4wGXpBOfPvx1egdszjuq07tUMhowYiay/CrLzhS
NCh8O3HzJIF7PuJhNJ8KTJVv/rJaa32X38HSWN7T/6DpDfib8bfi50rW5E+/
FX2lD3k0r4J6QuW80sDICBtcwQJRZk+V49BPTpl7gIgPvaRMRh05r7LYLdJW
ttKV4y6osiHYdvKoDJAym7Pj6tXgAIlWum6cRYSm5TRtFBPmYRC2EzMJozkb
TTJCzoRavSV9+et6lzbUUu/hfz9qJukTMNS7zGB0ky9o/Pa7fuvuTcJcSwCJ
dGYuc4fNJiluAxleKHxEPSZl4q053gRjGB0jgNIDm4GHITh1S4kF7F0ob8/p
ccNWDtzSzkuKFBmsVyESqVykkF3cq3NyMsIcl042MCYnToqiXMRrrhU48P+F
K0cW64fKRYzPd2v/oBTZvme2FN/qai9qOC5E3WDH3fin0oZ3JXwtS2unhtL5
lCRG2dMY+Lsxd1y18SBvbPAPglUwWFowshlG1mnwLoLcIKpMlNR+IH2DKJlC
3854eWyaX6KeWE2B8IAPlWpmiTcJb6W2AnvDqJF5yQi54ymmezfCZMoRsMX8
kaz2HeO5rvGgpJhmRpuhKVh3Bj7F9Etnf4ffIazzEAIE05sgbq9hLEgU2MS2
BEBkX+VscSLZ6g5dyYd/XWpO26lJcDk+Jwa6rL4mKFHxo0l31rzguZsUCTey
Oggu43bdePa4bo0wohkGlIuKX2AMVkCXL1W7e4dlcHwyQht+QRGB/jQQgOET
WvD1UpfpGB5qbb775g230dqhFQJPI/RA1fvn6HTraK/BIpiktIx/8OyR7vo2
8hXnJJTa5rnRExbptCQKqXuN4zcpE0FPgVEW/EjiuSGqfBainqQSjD7aY3eb
w4SLDNMs702pKZYtE+GQvb/nwhZEOE0CPzr7Us6clPbQlozrLvhLGxP1521Q
MfopCfiwdLEQIRibXXWafq7sp52AnmMC2BfnElY00UJAFxs00hIDOCAhIWxs
lNpw1fCieoF8RheD8l6cyPWRVrcKG50RuizyBlaXxoZ55o1c68yWhDuNu+gI
ELtNGrA7Ln8inNHXwGONNKgPu4uCv8eQsHwdXTMAZIAfSOFsFImQQU5OKJGu
tke4DgzQo6szWR+gj+U5TEr3W0aUq5QqW9s8BY3lSN0dcGqHFHATIHqszzO8
q7kIdp+ve+bk4rOkT3eDO+kc7lLKAu0BIcywfuBV8aURJ/C6y+vAI4K8UIoF
n31cT+r3Xk9RQqocJ7CAI28Rhfq4cr9Qx4fTtEoCJF2O+4GN0DrVyRquUHHr
MFvD/mA6neICWqp6srcwDtYNBBQHUkWTNkTnt7Z0+jPACx2LjZoBo78FDPe+
aWAJOjfdh0JOTM+mHyYpt3j1bZcBq7xAFNfIG7jF30Z3dR5pS47TOq74Sz3U
lnCqB/H1998zxTV4F85mxqKflwYfmIECHDpdY+Jhd1qjQ0ipky8TapHQomT7
EUq4pyi9vRI1lQvtV3THZwegokSfyB+Dlg1mSjYB5rtT0SDWUIs11EjbnZVO
XlL5tRRszTbcAUj7LHn+qVPHq3B/4aMGPi65xZDjePHtu5HGSVhBd0YLSDHr
tatr/wbHfJIn3XcYC1vWMtwprhLCl3cO+41+mszAsZrakrOYr9ngTfQSqUcl
V3vxUklLxN+MsSY0y9Cs2FvgrtfUXqxXYUM3nIhHSSN3I9QfCSTpA0w0RWlL
AmvkZa22WXYuC9a7PbYmetFbxubdYP07IGyz8G1yMFPl1yCklODVAB64nEUQ
+e4prKl7wivx8PyeW1QHWZVnTOiCokCJEPeY2gOk058WjYMiuS14rL5XOUc4
pCJZbm27ONHaOTRuSM8nOoQLmd/FKg5Q5iD4YhxQAt7xhHYVmjRxYGen2Nbz
OV6aZvFdCnSErvxMJQHJ/Qop8mpimJoxiudWSa6e6QRj4D0wip57onBlbn7F
12ITO7KVRrkgxoNi4xmqe/0p4X6ZFhItNje2gCGC5ocZLa0B9Xv33Otxl18p
vmrl0Qo/Pudi3+0mexKyejawZqOgLtT0LZZZnORqoQyX9tHbRmwozlzFWsxX
4ts0TuEM3VOk8S6EPJB2XHFhRdUkNTW6G0goQIh8gu0beFVVOMUy80wvQLua
WYYDjKcXJGg6DVrtV93WvGpamv0D8ldQbKDn6x/HvQPRtpli5CHGLQcmFRpg
1tPvuUOrU+OLwW8IwGlJWMZhDITkYpI8+7tKrLUVRqKO4dg8X6qrJwuVU26g
b7EQhs1uGnAdiwN6sxQJ9eWUSwjN3k4X4pYA+yd7g/GFCPfcD/A+I2a9qg96
9YrosXtDVjglCpcGRTQzMEJb6gkMfoZ3aC59nfHGsGG98lhU0Gng7BYf2fnZ
SlfeXDyH7OdPJcNyyydbMsu03aJCWxjzjZ9wV0OQBvDQRrPs4rbVaMeMEbmq
XToU+ZS5yqlK9B+NVK5eBSakP8TDjMBrIRiJmYr6LIODVffXrOwBz8h/Guiu
JucDVVgos4bsvdjsSIcyq/HE6/PNbwvl6nUrixdliHegXUjcn9rw6ftjszw9
A4nvJFC2kbL8LeYdaNy0RYpn4Asza3alBTWZthSoClcExvYbjRKnbuTwo8yn
DPpf1opyhYFkRrWKNOW4clI5pjwb6kVZWHp2FmB1UkvINSA9hb27CpTDtOuE
zxHyFEZ5rvIjWg5WFmf9adab7NzRSpCNqco9heHIQEVL97q9Tw2fl22TAqaT
RjNBv8vDYk7MpFDJgt2pxkLTttmXLpuWVNsg2FsL+n0ebaZjRH9STL8XqAPP
6WzbHSPld98rjVmM3wLNngWkjDpnpyvjrcm0uecHWV8mEZmX/nZAaNIFDN8V
uJ2TdWBqCd/vr15Xx0t+aUwoa1FfTp7cQPblpMOLJfXA271bLDKfrBx2eIV6
kXiN8dPxvq0SH1sDfJe/Fjc2Wom7X/DNtdinweVhzIQseQndTUdHXW+1DZsK
c9RQsg3J9ciQceiMdSuxQK891iDv2RG9H3jatnpeRbgb6yuQQwv72OByDEqI
4sfXD5WBqCNZAmvz/303rnvHu6uxeXCBbDhuLSPKZovSWBdqKRcikD+5d7K8
4wMG3b0RSfKg4z6RKTmGv9ZK1vAweU6o06bg1vEZ1Ne+Bxsb/vqO2tChhsas
LSnMGDdGPVxy0mJRcUDiSAyePzwuzJKUtXTHfMyQOmrLwdLA1yLLKs24UMQP
/g0Xmlg2Y2yX07ZG5a8HNtjX1ThDleCwh7STHpVt6XBA4PbYEEZlOb/OGZIa
xAhMz6oSGdIxSFVOmuYKZFPMR3d8C+eZrWW6rZaYupDHjcLFdtO6Og1yRTlL
2ILUOTv3qG572CDjKCaPq+Hhm/iX0FDvRFCdliavmaDBwLYyxCFaAqpieHZv
Xgf94LMa64/CYbysX6yOb3UjytfgglENgcGTPPbx+oqk5ahahSB13A71++N0
NRvJE3hXNHe8u8N9A16uwjo9dBT/R2dZ3FHFS2mJsseTvfDycKLBKLhd9Vsj
t/dUTbyLCHPZJX67W1DKfDm13gyDGR/OKPinii48PwTDzDAkfLsHxo9U9BrJ
kdbfpn3tUMGdIEhSHTeHdQuxzVNGqI+esatTMYd7hH7gn7Y+xR/JupuQp1Jx
/5JruLKGtT8rsQofytxXp2gUD65eI1jDrcAxjMSg5E52cn4zQ5W3E4XMaTci
ThIC0qLDHohPHcIxrYDatxTzTt74/WQoBIZkN+ET8nvXgi9Roitp/AX0Jtax
dgfdM4ef4ppNrQ8IsnLeAT/WO8560srjtFXHv8lbeCwm0GzmAGilMDYb/gKA
r7CMDiYGxkDDdv8PM2iOmGO7P+rbxDsnpnA/Q0Dl27VwnyaoPatZ5GoLBWEs
sqd8ZLYWh1LkuUJom0yOKa+AJnb7grnZVGwg3+jtx2650/yD/W6Hvyfa2UXk
8ScfCKP2ajH/gmkM6QBz3YrM7UEoSox/pyyBqLjpbQN9DK257y+YUGwBDC8w
ArYDkX2KbQ+VssLVom7kFmRwuNF+4D/o9i8mvpAWx0yotnpkKgfRe1K/G+EZ
b3A5wbbx3PiSdqO9iJ/4NNMmq9Qi31Ga5Co1QXZHs6a7RYYAWEiZKaw1yhG4
RPbDOPvns92DU7Zs1/oQYlmYV2MD/YLVKaZxgyyQSCw2kwWIys/MJdnImV/M
XLDX2tSNQYhDZGS81BMnfB5fzD2KYQezoTgXGaFM6IZWGfu9w2e7IV1CtS6J
OzKED78beK347KGjFX5NERnmtQF8fCen4orEsAH0wSxqzZ5YSbAiNlXXt/p7
vZ1QgVTqh1K14IVNMxWJvqDfmWl+F3cCeuoA09b1a8uNqjJZJ8uLY/2jfOZo
mXdTmdLrRnhR/5IMNlHel+2vqvOXAFvEsHBjMi3WybOYx+uLFC+QJGsQxKzE
ykw/MgmzvOmZxCY1Zln7V5KxGI//odFhITYZotipwltfU4UKnq/kDFFBVCOH
Ob5zgKDnwLvezBTfUxUU1lRrGVhtjkaDF/EoHBPFeFec5U5NR5xIRjXCFw2H
SkDunbvrrDwi6RZdOPBE7FdQ5mfjXIIjlTaJAGH7vhBoKJlzWlgyxh/RowM1
SRUsvhKvgIjn0mTQCAlBfUajQpEuJayTuvej3JTQWRdFHG4bRWzYzPoYuy8O
oCl9mcD7y6zOpQOkYoqYQ5T0Uo2cinKtT+D6ZabEV2frnw7J+O4XZ/CacT4u
uKOVPN5bD8EKosNtdLV7QxCb4oZjQ8jGVWX0qjEyOEu1wLlwqaSXP8aCnCvy
OVT5hFIDe2eCb44cEIHiaA6289vpRzNx9IyPRmYeFhftxvsItCr7WdHTPEvo
s9ESP1sSCqgxcrIqYx47ojG1A4g5pkw88MPn5pjZ04DtHi87q84jkd4Rqsy3
MLPk4UjgxmQz1g3LkUDZ1Mibcgj3fsZDiC1U1DmxYMpgfq+VoLYctYVwIy+c
x1GQOg0GH/Z1YSlFQ4bbSBQh4uScs2YvjfSl5DFisUUHGFiKLQkLCd/UVF/E
oV0bJZnnqKnUXGi4KyonUhhJIDmbIQ2K5NgdKaFHo4ZURtBFGij9ERPOdOdL
WXbmsRe7OGnWkbFhb9v7gbs7IORYGTK1fAvzdDbq7q7beim36q07uLAh39vX
N1XYTkUHf/5d5J7mXHdPPEyz4Wb3YC3lx/2p8Gro5+nLWmaU4YSEn/K4vYg0
a7uBQuttTzQ+LejrqQpO4KNeshg2Pi5Nr6juwK7avph6W/GOAsiuMutNqOM2
wladpaavGzWzOev4V9li+13DnzUzn0cBnPIPngfyaRqrx/gMbJoMwIxqxO5m
yjpwAq/81dGK4pDW0nMWAl4vFFB93Q8+7Fuhe6aJ76R+OWcSEn1eDb3PPYIz
+vcA5EAAE9s7hEjnwf6mprX1OzT+oVE9rJi4QCn5cKLT0CJEI+2JMjNphJ7c
oSi3jhMUL8+C9PLWZLFWsjV54ypaxWZCU71L6B6rNNv30I0wOrDpL76TULPv
H8aljlDy2NVT1cGC+kAnp2u4B3Xc/s4t0P0qVdAFlfsggVBwVvvF1c/4uBk6
l3mQwPviznx9OLSEEs8AJss+LdoYiVXbzb0aa/QTi91TgVnK7WXVU+eQgC+J
m8tFQtA6GNHigqVfxTT89dHlHhKSlbmEP3TbOtXKZQgoyw0/LrAvN7kaYNDn
atzEhBMiP8CxVLM8ZMGKg/vBudLBk6SAF3fMJJGftEjB7sf6v/qSpW33xQ08
hYgDjQlYWXvx8WCxYbdvIZPRwIZerMt+wp39hWj+6Np4tFdLqm+DJSmimzkW
SDma1tiW6iTczaqNQGcj1MxWbNeoOHVYVRyda8Wp4l7V0LwOv4UOtpLw1Fu7
deKpLJc0vBJP/rPXPwtxtFFzs98dOoJbrayFg4ez9PBmEECmehfxNIYYREno
qKJFbfPOZioFZlPGZKp28COrxL04/sNOpnNXLYiCzvhU+kUdYh3bx8D4jA04
5WQ9GhB1xBS0QrJ25N27yfwMUXmGle6Vb86L+PG8ecTbF414xgMF4F7Uq7hY
N+/jZa0RCWsZKYvWN+QcLpATZCyZgdQK4wKdU3u79SZ4ZgZFMKPLBJEnsD0U
hA9yoRu1KCvc/Qv8rh2AWubJEce6fTeHA3XuPDPnj0qwHDbazR5p8O2Eq7jm
CYrmOzZbTfayU3r+mcm43wL0XKvsgIlc+48ZbZDPBJHzXRjLY6vhbVf5F8QG
JkS7rEa9syB/H8N8ZMh10f09gNZFC6LkMkq2gdCWuEyVhczfCZcmP/wm/iah
g4KJl8YHhTKMnpJiu+0Zy9yaZ5TV9T1MkDRSrPcgNfkIfbrR+8abLWg3otTw
ur5aU7VD1KBd15tYAHWQYDBY2evclO9BuixuYOOWNuGLd/gudBAvHejMVq3l
so2QCz7Acf3n96BZ09uZH74aD5o6JIjoHGeMnLv1bzpRwQKoY2KMSQx3R6sq
O+f8R9R2O7vq4BYn4BpkfulTvJdcEcz6ds7hEI0hEO4kBmoMty2kQj5sXrry
+AsFl4mkbpKXRLpEYRKrH0kokPuOs24TALGHg25enqw2gtWESjiuPN9IVpC6
g4bB2XUqteGyqrnoX6RsEFULKmGsyN81AHnPlSTOUorfX3PaAIC1WSeAaMTV
/vgczxDSTRbVsYKBBb30O7Bfdlq56uB3LNQ3OOZSNoId6j7F7VFec3GarN8F
Vg6FUNezOseajqKpN2mm1/Bl3PLgVq7Z33yjQQpnyg52OWzd4/vwksK4P73T
hmmagB0US4eK9IXmCLRZxlpq/3gTZk878ve2dyx6dglyWW7AgpzEsNNEYGG/
gvobXiZ/CWlgUnClhb4UdFp1zsGcnvBve7xU3c1dfoRVkFlrihlpp2f6xHHN
O0tq66rZVpMayErVM4IV/a/bRD8s80ZvXUh7LlLTphsJgrX0v9BcLIA3oCGE
3XKPjtib4vCWbULPGe5rkkcK6EqYHV88wLXLqQ045yJTUpUJoOTnKTHQUE6/
ETFVV6amhi8SkaGh9Y/gyR5Clb9X9WQJ4KRMGTMXbJOblt/Kwgq4tztidkoo
BPtbR2GhVkZsRgcTHgFzTvimjrvbTic6rPkol1EMUfgvt8BIpG/kwzU6izEA
QNJRF87qJmGBhQV1z7WD3SzJV9GKy1XRYVfWUavlR7dDGwPuhvF8RswzQhl5
Wek/EibDQmba0MiRsbojD9KSOKeHTD5gk+ycvHSZIrLPjcbw5kwiVI8EDmVm
bI56ynYeDpHF/0qxmI88OMzRQaJiII+SGD8obUBImgTuMv/hC1s1r3Rw8rxk
LxfJ8Og2J9aarGLauD2XOwkGLwfTTw4SHcy5MNphYlLxjFOPAqJnUxbN1nvp
D3DMwzJH6XFfZcIqN1JH85LICgkeFbFFNNqlZDTeIJA87e7hzJJc6TGx5N+/
4QFawPa3QkbZIiHTBZRbGmbPfT0b7Nw197Ebj46o33DTUeobHJVrfRDSszgg
3epWU9M6TUfx5U5uuJvqt//wxyQeIsEys7PuQgVnOqGkz+QEdU5+yi9RNsK8
nxyVN+IkE/rAAF79B2WJT5FdwoNmc/q8uzx8h8JPZvOxHzi7QtRFVELv0cUc
JfZW20fb/r3h+2KA+DHlf6wPgSbuzRUllgtcFAdlNNaGaVwtXHnl53yDJ82Q
ZD7O4F8jFRH0cpnwlvDY60p20l/TkQBLhT/d6KXd4dmomgsVRSitf2yqyZop
3GdKiNIPMgae281NoYKmseOOFe4YGfKaYsHSCA1I4npAWTIDr4RWrpgCQBX4
C7hqFQ0HZBtwzzk/UpOZjFQRp2fZideqgJkMMfUcM+GmfifT4OySnfgfnsjZ
e4GnU0vUs91cFS4EkrOSCuR4qBxiJpNSKADAbB2qF1fKfsRj85TuYV6XO3+G
AKG1U+7LC0f4ZvMA745UFX/HI65e68Nu6X0NJ6OgXXt5Iic7gA7Zpj6yzUbA
guOwQrUEMnOCWufi+nJAujEkTpkrpq2vOOJBFurMuNjhim1ssHkz734DRj1b
Rj6Q3EAQ0JDohS1EOS78Pwd1bL0/Afzga0hyZ8qlnL6JhbxmuzmYT+H2NigB
C119pc0RggjN8ldscwK1qjRaM3utJlfbaBrIGFErV4tsKfYlHQrIFBj37Ruc
uBAjhPU3A8albWPczsU2+cAZPlD3A/MbHFH3vAdeMFNy6LpE068uewEPx6qu
K+58nP7K16THtnToFWNr9LKmEFo6IstDaRLMyj9nrpQ5UkLIPxoWt5185Ahm
9MymxFxFCYzszJox1PR0ZywyGOsCo2eV5E/OCu9RfCj1J4m+SP6nQx0GmX/3
n7Bmpj3wxWWwnMxne4+EPKGlIirqXWA8zdmnmmciHxy08rKfA/hoIqWPbNQs
QQu4/3OO0coBvM6J2vamtkpBYLPzMGrktFGMT+gTzD40xbneT9Xfo6Xr1Ujv
6Vbc5NIuOXhqiJ6gmimKYdr6vHdxfHqQNzEl86QOk+OeGP9tB7hgwN7Thph7
27WVbHg9E3BmT+61sXkDfD1q3u4kM9/OR2w8oODIESNJfhhWbqxKsH/MavPA
8zqdXQ/o2G/pV5jNhrjOIJv55jwcUlrsmTQxAFmK0K/a9RAMTpC3jbAK9DQh
Yu4VfrVxTyMsCOUdFvS7kzYG34T1DRvl/W0sMXciIJUZocx4tqrm9PHRo0uP
178s4OntY0Ql9a7NMOAgOxcwKb5dqLIpYvaDdyVj+7G4DYJwDT4ZY755SSbg
1juixdQcVj6Nd4Kh4U37WSFe4DjB9Dp1IpJnHFB1g4eQXw54GBbwLejPXhz6
W9Y5K0b9pXkB5lyIVKwhQo1+7zLdGWRwUX4VEGhAaoMYMnv5TsU4ZZwF69wH
K9lUDNgaUKQ6lN4qwLZUns2BqXUGkOAyo18uwguuN8D/PmV2QGqN2PkdEKLi
DWr7cgYyCtnaQBpi7OoyNCD4AZ1dHRse3cpa/cemc++ZI98+s7JlCfnUbm6P
7MQEleTk2kq5V+gblkaig5Wc3/XQ6KyUxj9bPYKNL4g/VR/LUvznfQl4Paum
jgbrqZZRa6ge27CF6vUP4AQHJMBDgg7CrmTQD8wZacsqrBmjEa/FzUseomU5
of5LUynn3iSngfGHrsV8W4YXSwILn9+VQAObHDilT61Gr3cJXvTJ6GGPvD9v
wCe57rt+Sd1s9i8JJlqshM6rrzWoxQTlhdRcyhx0BUmB0ErqvsqNXomHM6oo
OZY0XNGQtHB0XOOci2Od6ezU5Mayv6KRU3CVCwhojH4ZH1rgAJUBJ2DDbYHM
1pr0O/fgaEBJQgdEJitLCHdu5Rd7MEyN3tRSTLVQMpjG4hiAnma035TUO5LQ
6OtAIeyZAAxhZekXXpDmDginRNjYpzL8bqQR/IilPDIzjfO0GibiEPa2WSCM
i4YoJZ95lxy9utqzMJEDJ637GEt0zNJOU6MkHuEwFIHNngZsyE9peAMSoQkc
oxXSkv7owAaUUPRHdIqH2D48y9/lHPI1r/lq7oLZcvE/0WhAZDgUt2TLNHTE
9eJoslWEMkIA6MqkAiETtyxj866U7hfCn8BAR6Xnign0LkFHsVQKskwzukPY
q0P7tZ7jsuUO4973hI+mhzhMzrz9++3evrg59L6nSh3B26D/UosuOTKjyVXj
1kOcs9sxZhbM3Le9hxueIeDLmpOE55BC09Mc58quJJ5BGD3vyD0KbZkHNImq
iYe3rm64a8MNHzMtnWX9gsdxcj3q9x1kMdalZ8Puxs8NezRmHo4b8XVAUVxz
rRm1PWA0EGozrmCJS2TngJMfbp2cVh4wdHeKvfTqNn3GZ5SvV/wUsScNJml7
5h9rDpXbSPqBICWt8EX9XimXwkR6RMPIWVk7sQ9lKYOMXGKqw7aKCJGceK9f
NuUuBZ84U2QIJkE6zB+YXkN81c9AwVb6qv+CIqTjSipCeN93zBE6KGWIJsg2
QmaF6Os0oZCGaobtkAA2E0EQYX79vpXB806Al0z4FfpTAgWuT6Y6UTSpo/Nb
J5zRxEORcKSSfRRu6iwqPCwiLWa6B01Ah5Ql+cKwzmkLy2y4auAIBvrrrFyV
fX95835vxyXnxaWPnPTRdAxHKFXNaHcgcR/T1iWwgW81K57WpDZ/vczo6pnZ
ew/6mYAZ9r0Vt8O5pd68Un/3y9eooJw3KBuQijKIvS88l0ehKJ+5Yz4pVeyi
NZn3SW1xtc5WdNtCtfnwIl3chUh2B3wKmzfb+BfBSCKS0jdWYHQBJWG7ZhQC
NWe8ftmJ9MhPCWce+/nxFWPCjgX3K26ZwXsGSShFzBhncKeNoIdWcwqktE/v
tmFj4ZCCZo9UwnPCV1VvzT6R4nrwTWBL89kYoRhmPhbiKrXQgtz7HszUD+Xc
xuQ90dPakF/AbLSuWj5udrhLpvfgLYsAAPegFv29/tYdjuuzZ1r84qc/Yg0L
/krZUn4Nf+kFOaYwdwHIJWD1Z6JElwwUkr50NOOhjUNCWZFIpVLKV5vB/aHD
oM+sW+HXn5Aeh4knBcrsnoiAmZwvSVEbJrY9+j7bTuORRh2nPCGxpCDCC+//
Uxfm8nU8DC7ZC1h3UvYkYAEAzt3aKyTPnhk/vpz47DZQ31gu9NRD+PtZt3MI
oQnJCE14Y2+UCG1coSzh0QCCuouyzu80YXmdAgx5/pOn1Y26dYDFxS9sNy9T
PsezafIuOg/ZtXX62SZ6MZ+6Zxk70TS7GQWiq5sCPiGNSCT9rxVKjj03TfF6
Jv0UcSPamAOYMV5XwC76jpDpfr662SPaCA295rxFRWcn4/6fp+hhIwgh5Sdl
kd6kXcRFvppP82E6WIpji/zLqZAoQbj6q5OziYh/qM2bxwL26jNyqW3DuKHM
++Q2d2KthnhNxeP6/L8Oh10hkEBaUC2Pu2UsqWf45luO9OqnrJ5kUD9VXh8q
EpCtQK7FqQPIMQaxVjY+Mstdl4Do1fsZ0QXiDxYGDP7nnNCS6zh9h5SyDYqk
F5BKLfxDa+MTYcW9NZwIeyYeZ3VaNBAKS1JQ0fMGjVc/xG45kG0GmN3yaSR1
AMOh64oD+oVicFtOrrYL6lBYzWlBsNq+dvZJP35HUtcieyqSlJrdVUArBjpW
GB5YvUchJMbuL3L5nzwuPm/amXflinDdDXfi8HSoir/l9z6jgiITvlPy2/Xq
q1xU5ilAnIT+gziQZXpg1JVNJBKp1Lp70qDm40DlzcO8nvT/Dbi2GQvuTpeB
z03uXwGC1r5ZuAyaC+NCjc9gkZItrIG9y4OY74umRnyVTwyGefqOht+IaKk0
HdndDOh3sDNrw8RbB4jS+lfBhHEQiHZwyUp/3iewUIIdRXfqMndv5JTQUL5z
a/oiLiAscRnBzzWUYcWqgiRJ/GOnuNUmF1dIVQtwwCT61Gzahq55gNWxpnd6
YD5ocEr2sXmS682/HpAV/dlBz9tcT/0xCJAlHC1q+Dfr4UGKbuySw6wO77e+
ZPhZeyfw60jb+YPTwRfoCnr07iSJ7Sp+af6jyLV2627lbAI+7wz7IrspDag8
ERaImw7bOmsceycImhxS4WSjzpSR7ndyW3UVMfxq1h7rgjuvFuVpm087qGGu
fOjZHeQKsA4dpOwKyxpM+qy9yhgMAvoKbHOAkSXoEQLMnjvn+PPK6uMswkMK
Xg1wJbSJVbIz9DLUDSANfpWBJCpjZ8UQDI0VKeX4rQyJd8Im0PpDngxsy+iS
iq1jCLOB2nVZeo7rSXMOV2kFiiQYLelHP/M5GGQW2/KiwH0MKcNlBUOlDmlk
X/JBV8GbMDLxbEE08IdUgCWWcdqURgYd5yh6zIuo5d2VYpBI2okpMWpvse3/
QLQxOVj2qlSJYY6tUyCZwIqTWNBA7e0f9ky2WeSYnmD7fJPbDlam0LvhqUZX
eUgrFEu+jYTVDq3tuixNbO/CJY1nrB/WcR9trTDxBu/LHOxQycLP8SfVeiiR
qb0v2sqnt84a64UZIPzDJosD4yboBRfwvv410Fp139gNA4g10KwBgBcCn/p2
bjbMcwYcShYGgkJHElpfNCCHT0zNweWzbqxl6LGWxd6/OQqj8l/EU2IQd7aa
Dcu6xnhfJXCz5xVl7i1p1LVAh2fG92STBd0KMnUCZAZ4PMFs8WldFbnWKqGM
XTJxZI20CLsWTCseh32CiN5c/CeZJe0dh7g7ohg4fU25w2ZkvTnadnGg9CSe
0vqUi2567jDDJi1mOkpm61BaG/xuiPzBid22cZ+LOyqy2eoq6fClPhU5DFFQ
EkOk2X7S6TdO0ClBkm147ZkhSVg6dwIJ1VMTy5LkCPxgqF5I22S+3YiAsXWK
pVxSkd8loQUJvzkuFNM9SQmCh5peJ6woBEAR2x64xuhZxCVCH0rnEYvF2ybs
JWhgGGac9W2d5vaQbwif/pJvyrcQAbnfQx7jRMO2aLUQAaWGgzzT3RNnTX3L
HtuG9xO31HRWT5LM/j5orZgLDQ780hQRS3A20C3prJZUWTFxnR6R6TXerFfF
Uk8b6UTwNyaZtun7hBWPT8RdSWDVxo1PkuXzgBtx+IbbUN9HisVCwRT50Dsq
BEjUkuStGXvutfMZJBw2jVI0Lx9dWdjk2ZmqILesQIwX5tGq3kvFw2WQK24C
8JsVJZEIy33hLO5v/2cwUoqHYpFCFZad1mswr05pW1zqov8qPMKMKjq7tFRM
+MV8/I6DNxOBE6OByaUIdoe9W9JgwAk0xNQVg5tAYQ9lqYnYaCjURkBq3G4f
pgpzUP5e2C4QRRzjKkEkWznZuFxq/5wlI5SVYYb9DWLTwxrSMtCMZUHHfPTM
wVwH6a28hWXEOBxEzang/MlvXrN5eVKkqdp+jqxxLDog9kT7c0drMg82tZWG
KCXw2SMQ+cVLu32bA+6yBgNM3G8Ivndv01kYUY4a60u2GGQhOcYdH6gNVPpc
mtYkN7JzFTaL8V2Zur0ZdUFGJ7rriE/qdb+5e3zvavcDzorGjPYmDx/J6Fap
+/f7bF8Vm6TDWGW1PxrdCc6PAek2zme+rpXrSXSiLa2wJ3pTZ2Nvmv8ZODNE
4j3hWT7atJyqfv16gRl+CHXl1VGe8gMSCxvI3nRbRnzmCHsdyjafjYWkc3go
e1WPQFxoOEBg6aRENBcaV+YPwKlx2YuhsL4V1GanzxYOBhrmX81xY8G78OD8
XeBfwmMUzrtMzTCur5N/s9AGm1vdntDbynSO0RoMwILXJ7l8+qR2O48rM/D+
71uhwcJExIBXQ4L2IBJSdXC+sK0h0lC1mE3VKc6E/j9NalOwmv+KmB7jqIon
nET8xpGPO8XJwSLqLjOI2CeQuSpHNWBy3nkpPYv8qzvjYlyWfnQIdSgeqnDU
MI5PzV4MEcCUFSZhpouoVmBcOn4+vCYTQyRfmnSBbXvowRzVOBFkvzssEA7X
t3q+ur/C2RUtXxJT8EjVT0/XqFggLiJU4RNtGlxnmjwwS6SIL6zZ9rFI2Kmf
CmbIvblupnBbTw8PF5kAYvS4vVI1WHxfOw1RdLFPMEF4OlWpCy7IHgFuqf/G
kCQVg071JD7iFhGcIa0EYoCqeb6/kf1wYO/WbEOtmQNc+SSKVu4NqgHA+nTF
DbIWUFbGf63n9B8qDiddi6aNvve2xiyuy6pAjZw2I4pv9Irt7kNDgenjkIcD
EX8lWeHV46yHts7wBI1yWPZgJCO1/bo+iQi7UvC2WV0dEigjn/BLr/R+g/Me
pweoLobGqrT7wNG26Ivp3Vmgs37fpQPjAzedCz6LvZbkVTnDjlBYPhjNJW/6
kzXUpY0EAqTrPTTNKKfr9Re0NyK8Wjmc49FxaB0pcQGAxzOYIwNESegPOy1r
d8rGihsbgsqPGWfMGyHAs3dOhbouYrRUDBRulfkdwhF+MKuVyXB1ppIjr5TP
ardivr2FL67QbQN/HQJPM47wzwnTrPG90aUW449JYbdE4fDlfjypbIXK+CZX
BOJRpJLOhkv+khl4YZJjaJ3L8sVyUb3t3oZ3Z9cw2cHCkVxanauuHMX5mdAg
C8en+T5jq5eGZ8CL/i2ddhW7W40T9ePMUVt/nh5NC66KtrUNbkIHDUsfghs/
HBZM/fjMd6G5wtUCMOfucMrvMImpS7FSDHdFXSBqc/nhSlH4FERJZp5TEbtY
A13e6mwVV9LGEJB1NJJS3v5T9755sywP+XSETxxZk10I1bzyrtj6j0hKOTLO
i6xLXDoxMNt2cQTaKa4OR09QqCOLckn61OF5mqXWB2sqcedAiZRnfR5h2JwB
MXctmsEUQVjJ/5w4N6DF9+7e/OUPBA7onORMSsX9d5yewkE6yEhSZWTOV3su
P4Ey3yaITfz/ELNrQiJ51y175RhJ1CVP/I44He6XukvqE7wOsWEKvYmOg2O9
tmYrk3b3x0oPhFcCriF4hpKI6RjZ/3fWQaLjlMH4KAc8+lF5UIc+YVQEXKES
e44p+UazpcRQRVMHccsVIOloVtPInBdqUKuzvg6041caUqEEbm5dBL0mbxbw
Z4w6tTBirC8G6No702c0scfEu/UmRLgg1CZmh1oeVVCOrsyp41y1WOUeo5A2
xYt2TfJqP/1aJYXEEONnPu16ICJrmvQPqdDpxgVuI+dHzwx+BqnyVFSCbwoV
UjtmGReuhU/Tcb70++ZZAzUb2WBj6qHsdaZSE3AKaGxVXlu7MxGMl9pv1rDa
xM8D+ikQXrwom4Yglu/jz5qQUpqqqTgKH2cQ7V2Zn/xoZpVCkEIoSnPBRIHa
GWJmXl+YnxDbNMXn7C8sHsdz79tA/yDQcyNvtBN9Jeznk5l+VlQtukZPsALI
8IwEbnz5RbS0Yi8l0NfKZnUKowotY0kL65YJ3Qk6c9Ao3hsH0x2hhkCaVpqS
KhbtT64PBHXmKMFVG1f4CjEnMAL9S2Nuxx+yNlzgVQ1o3KDf7w+Y7vcKbALj
J74F7gBNG7M9FTNg3keUpTC4B4PqnPAySnNKimigJkVIafTMbYHZ0wYBWI/B
waGlLTvPjEPElbI7MhAGqi//T90pPJtH9mIux3n2xPGtlrHpyz1Acmp34FyM
rl6POp1a29YVnzPITtEeq0MGmssU1X/ptdbLrJ3+2NF2XiYNhRi9cZLDHQCM
KwVOyzul7ODxQVEpbay8KaP5cfHHkBaSJ/N64d7TZYCpU9AzK6BYyLgGtrns
ye2YGxQl6Z1jNUGSW/iah75coDV6D1GDU6dtcGDVZ0+NEyD7+Xer5vFuo7na
Fhfx3SheA1hBbF7YUBNjVmyRSbyjL6yn+ibWM7q+j67PxfbblOTXj2FAOhzu
Sn0S2gi9pdTBJ+xt1t2ZJ0zlklP/6ogSD49Q7yKpfVkGDEJltZyAD5YEumg4
Cd6lmITM1+gL1b/pgOZmnRRFCX6mzJMb5ESUmkgB00YE5EDpbvOgEk31lvN+
p12RsJUyc+qjuYklU58OCyzOaDrSbSSm4jP41an+EFpeh+nAqisOkkzU58pl
kVs+avNFCpCp41T4pdZgRNN9me/nLxXbFzsw1oxXoEX9o6DU9aI07wt83dA8
tVvdKjL1Ej82CKzsjvgmq3aRdRBsNUFGeEUqNqcotSMSFaDqpr8CP2jQrLnV
oX1yWX/rFl4Vwrz7qqEktbTyT17fOzT4+D5RTXOIgtEA6y81tgSy3SXwmXyT
Yie0h5s9a+HmRG3TKEwi59qePw1oTkYSrC/mIr6p0f2iLrahMHx7IKtaGlCp
1jSu+63CzJP4z76M+JucKEpSCmNUlsgbUJL3oSKzbeZkn9P7aiMzy/qhQYCy
B8ng8tPScNU0e7TZ8k72fcIqq4sC/qVOqw8Zt6J1lkhMFHraKX7GCS8DVD8G
tSP555AuBLlQRMp/hVA57I4dZ4S84XmldTGqqicP4qrSIjpiDaDRMknX5ry4
Arr2zFS6mtlfH5WMKSTaQSUgNUT5wZ/5e+udXJ9kp2+7RRdOVuQ/R+UOaUBl
C2+ipRgbiWiU/6xATSHPWulrbqd0PpJZMF2xJO1UOxmGLweD1s/xtAbO8/aS
8yXfZifVTxCUG3xq8Kf82S4l2Ww1GxsFHtyblci9joJYjk/hL8LtbUZmOykG
QhDGgFEaxNH/th580ohggEZXEvi4eTFVMuR0Bn8emxAxXSKo8ALsf9SE8Nw1
v7cPsKr8VRyIhJ8/C0Gui9+HlfQAHOJt1MDzCYgqC3kYEhDs3oErnGGL0z3v
zEeED7EbJsRraIL39SdBVpjjl91XNd9ATEESL2RSL1RzosmH/BaASOfvVCSm
xej+vwF6cqiGUQSSs5Ctad/qNH0/shHLzeuUDn7vd60+lYnJrPg9HO+00EYT
5QCZUVbycJ1Ue0VliiahZ4SLJKzfHeZK9w975VDYfyTwWhIEt5xZsQSgyw3b
kPPxtVIJ+PJnSeaVuFYLDoDSbfojR5wz8zcXdsDV8Ts3LblAvwM+ag/aiVMI
ehiNedA9jloSZ8giTPraXLUSTFB7/rsPXb6IV1vNtQHL/7pKPXeca0FJPLZA
FvvaqTAboLYeGZpdpel2E6vTZ7LJTsbuyH+fPovkS52Od1spQNLm2t5epL1y
EoYCG7WNKVrC9OB9fIMEPavBzWYKnJeDY4o8eWFzf8W+iMsfN23J8WIXlFlC
jzmYZZUqWLW7VgI3KEzsivfok/HSahrPWeqeBSVEnWT5SAzFbBS5rngGszrR
a8HpTHWFiPZFzgEerMleyh601MWt8MYrTO86NCQ3GsgwOJD7CbDuyjcupREE
MPdn6B+KRCJ7/Jwx30gHbxDQNuKK5tTrwN9r7DfM+AAKHQWS1H0mA5HLeq22
nMqFUlFBUeZIZ9kWp2Dqs0j9kvHUzVhSnWWkwY/7Z8mzVy0rnhoGAyRjv7b0
a//11xkYY/HZD3otfpvx8BoKgJN8TZy1PasSVKln7XS6blusk9dzO2L96NCy
VbziDxfULkFTsD9KKFkaG80GIaVh8Xyuteo5zvEYPN4yJPpNgjNUxKtfZiDH
BQQtQKDc/8/mKmVtTztYavTxrYsHtNbWmzyFI5kuWqi/+F6U8ycK2YqJwpr2
YSu333kV8R0fl0vD/ghmqPUL4/vBxXvn4lCnpc6lederbHPd+PK8OZmzmLRG
yf/714R3TkPQ5VPrmXAUjrkM1tN9q0RPGqc1hCNM421CFOl+Dhwuru/Tl6ZU
1DmP8ksUlVk5qji35kYdKFf5otOtgB1MJX8udx6jSZogxOEUxrgtTifoUZnZ
0yN/MjMqt6r+RdVYdsxDFABSlc4w91vrsV+jC2VSkHrD+VmyTxM6bM1XFMR3
/slzE+jDm2rQkbB8sZ9khCZONiaWebwhyUl8Wn7dRkXazXrsjA4dVYABfMu+
AuXX8swrOwggZVwheOeW3E6QoQ4ZXy3DmvMvkuokSukRZmawSkQ3q7ShiGZ6
Xosnq2CMqOUZ6FDttVTVdCDWFj/cBjGp4/TX26suYUHjjAd7L+B4R2FCgamx
hDjiJDhPd2sX2bm+eyNHdqUDpu+32Dycrg1/XoJUN1QjQB8RIwD7aSM5I2iE
KLeWCfgeRil452zQPZoS08jlJ4te0oJjGuiUgJ8IgMMH9Ff3/aHaGoqzTz0g
T7T97hsCKs9zrMuGoHCC3TS7x4cwY+CCYaBU9++fUb9+rn2v9hfxsyWS+Fii
Wdcb8VijPcZMUZw4HbyC2aCRiJnXr6FK8IL6a3LZG4tfiUKYa3Qove3iZjoW
c8+1w9XE0GYTHg+UoD+y47n4O3jM9fXiD4xGwyni+P5ycYhDhTtwPAcrxa3V
vLljKS72I55gBIO/po8AUMa/4nfWOtCfqxa5DCsNQFg8jdmJerHumblSI+00
+LOP2YBDcTESRlcQ2Tt3BZJaI/M8k6T94DFb+1cHxpFov00qEa67eYZvBJ0C
lqkiMgwh4CS/G5hptwMJ7EAKA/8ozFVTzzPFcdSwehADZzG4xc9V7Mx50BGR
Pa6RS7L0/p2hvAIJsGrgbEoAHZSMlf4JDjd3FGMf4i9oWLNfVDmgwDIc2ZxL
54rpRrSz3xO/wNSncIjV70JW2UfPc4ONzF63Oll1yUd/SG0nFfDyZe0Q4T9d
Meen0AleKoudPZbD/8uxA5y+eKWntxINbrNa6qw/UvJgSBOlaUY7NXzelBRT
OrBv5/NjlbYcG+SZYHaIAeBo0eewco5n/8XI8J3AXMKUx4+uHraXyPnwhp5t
gBqddMD9CKW+nxQO455SuzdkGp1jy9382bmzZp2yTCx5/OX0wmarE0Aifn5m
D4CdIA3U1c1knRPhyJfsY9mV8e02knA7jV2vR+zH26vHkYn8bnwtP4zaIhWd
IbX5zPuUFR+vqRjc7AbHOa0YmIsDan6sAqJ+BQbSX0B2BAEpceQPqkAbrNLD
gJUBADkKTviHUwgT0MPcw/wyAxSJRBBtSCDndGngPrSo6qDuVqX8qsjYQiIf
ln4Ss+ThOSh7d1nXAEnJTIEqfoudaY++btTxKuMExniE/EYd/SawGFoomCVL
Aa/MWLkAoQ9y7kmmIwLYdHx3RCUPHfm9zsZxir06e7ceX803Nq0MNQdXo5OL
ws/rtzZTVU1B70DTX6bbQpdPncNlEIae8vQR0tiCoAjy0f+BJyqGkV0r2+S1
L6ojs4cb0yDwwH9wX8+kKMOY3GPgfNR/MCv66KxtXIidpsxbsHRMRAj6nBiN
fsyksiZsRm5LBq7nAgArhvU366UnzTFiC43tP814mmFE3KwDCX/wPvEM8K+u
W1LyjSRxdfWXMApEDNX0a8vwv6Q51mZ2Rs2rJnaF0C/QnvEt268rDH1Y5Lg4
ICHlH+1rbbOb0R23fj7p92aHepWovxUlLwFCF/K4GFUYFFRtDLMEScseIC//
QJtOHz6ubBWvhCLkewjplHeHHCW3VVNzSGZaGHMD3J/Fj4/7Jjx8lgNrH4Ho
8coxPk8quE6Jam0VlCWU7UP6tq1Kv32U+uo1xgHuBtmS815uWwbMyzts+Dbf
gODmqOfhod5swOQcc2wbOloiFMtg/l3hHgk9dba4+oysnIrXsm7rjfYm/WhL
A4oSxpwpIyP52MTF/OIfKif25vrIAiBKzqko8MzODslpuCGZkh8ur89aJyBl
FC6q61G7pQUQMWuKvIE6Pef8E4wR/cxWDxcs+t4Jjga0282A+itzI7m04dZB
RLFNpsazGhiRproekvMByhkWMD9BLTAFl2atWTvMUez5a8W/Z1UMV2YBnjx7
UZ9WXeNF8uNnFBEySTJnBRWCduOoJ0kXlBrInDixhtLbI9K8O9gcM68qdNlH
/UjYpHiVbwCV2JzGmgP1vekr+jZ3rL/I14yN8mBVjOvZZVIapVDlIMuotyem
yjbXkGcUpLeFwC1qAt6HpMPyOwAiEHIfPTemfbS9r1EvirrqLSpUY4XMVBS0
qHXC4fP7Lw84yr22UFRGNgXkJJx8j0rRLDgSAFjrIqWlcVBMMjHSG10Wf/J/
/qWCEa4jDZBROl4lEv/52fFkkEPaXgApWcF6t22MJiSw9kE8Ksz3caLFqI7o
AQj19F+yw25eoPgnyz0FT5nZFacE+WORRH9XCazdi9LDtk0470GdiRmGn8Jw
wF0P5KCTpJBcGeAOWmybblt2xK3qfWfD/H/81sqqjd9GFYTqpLkoLIhN7I4L
ptwWBQ3FTyfeWRdLVO8mp2wrSSJ6cH4SX6CMspefz+TJKs6wxKYFz/OzZiyq
RR2tw5ulRTDDcg8VFmQnYFGc90kNd7rjKtZBwe3p4+8PoTSfrxd4+J75Sq0+
2BcGqDRH8YRbgRRT0IPUA+JFFijROoffErrcMpLu/Mf4kA9UH/p7TYMCSepN
FZW7/NcSJ09nA3D3PUm+MV2qKQ9ikhYAM+mpXQLHuQpX0Rl0/631guOBg48x
eIpzP3eivDwuRp4bJn0/PdlSjkC9Z0wfNNy3Dk0zpsFHBKJ+ARz/B1kfgXhx
4ELjQz9qXR9imK0A1q2PQXZSTVj9//mrLgQlbbcTHeTACKANZUhE3j1+FX5x
edQ3oUXznraYoiDS45p/6nt4RntLDOgNw8R51RsTegbf32HJKfftw9GjQ+ji
+Hdksqyayuza/dzdY/hqYRZfCI2ZYkBYgkbIcc0JeddT2sau5EytQ7S7fnxY
7vFuDsFWNdYglqxHDLIE6G80CqM6HDJUkC7bEmsfIQCg3JK0xeZLd9Z12mqg
UkaJ07wGHwwhEVaLmoSMqNDG3JETYZu/gA6q/jiF+z44omNoNBLVBFUrs7Dw
Tk647Yn5SBQhr00dXqROkjnveSfmEwYCAQpPw5b3EOoVf09fFCglGGUZWkyX
ONzDFoFTsaE+g+MyFw/Fpq0DiYc+VDbJImoC61Py8Qu1Ws43ZSm6Qjir0Gv9
bn/sZ/0feb2Mjxn3Sj3zb7lbhW54yDt0kNklzHY5JMR32AJvGi9C20JtjKa0
B2r0WtTIlJ8cKgUZW+x+4XJQSIsvRbxooyGCpYxpHGHU8q85ZjFRq2zSDchf
fr7NExSm+7W6GTiXRs72KnBtgITg/Ki8C2rxckvZPc4akHsh2CgTwT1YO9lP
gFgQCW1ZXGxPIEbCCFN/OCjjhMjABgqcUhCD51nAhv4Xu/y8W7nPM73lUnq1
49WZsdeKED50LFa5JBk5rczsrezXEdIvwSFcwjz5qUSwQSzHsHMoa5KipbwP
0xs9hZIvwe4L3VBG7l0wODBFrWbyeZ4bE7AZvNYvplQzJS2tkXorODRleuB1
wTIOjXZPNeUxibNHouKWunbkHDwlwccJpl1e4JaCpK7L0zzfpFHVXqz8cn5V
ysMw5OP4R5JrtgrpXAGMbiBoOhCzdkumhbcIikUvSqV7Cnne+vgAXvGBIc9/
3ffa650lhvc2sGi2N7evKew5tXGDVrWClizuJW/79HFEaFteDnb/q2hmWi33
9YbdyM8LqSSvIGpgOF0vEnLvHJHWBB6HU9OVBspfUg1D7EcS6qBf9z1+QDO8
h29nr0AMFqWR1rMAfxMBC5b6a5yLQb/S8uowhIq7qSTrTUmf5qGLB+9pyqLf
eTCXWxGqMbgFvILUMCe7mn4Mk56fPgXLiyJu7c612qxiRiA696ft49rO6SKV
4rWH+tVl+0eDCUO/itBaPPON6QzgO6GXTs9KLzWNIp0uEvxO1+AGjWD9tTzE
fO5L/48zVVz5/fdT8p7rCZSBAfnj869rZZwK8iEReBigWh7NRGeV0aOry4MT
w+tDkmgQLN/1s4C8vMoxs7X2rCmFIlr/RiP6BDW0RExQbW+CgAb6pLp1dMEE
6ouvBuAB8Vf28jFhpcoNTzUkaRJGAYV4mZ09nojaNc9gRclgALSkkYrPbR96
dZszaETBo33qeiovqOfcnrB8GHxXeci3g19OOYeNSVj3gfV4ODyLLjShno/e
ImmDQr4T9y5TAwKytMSOdgmd7fLcHQEV0f6fDSR4lobYr+zk620nIhmCDBRC
4QTKEm88KfSLepj1xN592QebhC6WMkdO2kHccx/K5YhC/ug/sXL9BjaSHTAf
BELPm9Nz6ZqCIl7WYg9gkxnJ4XN+MWdNdweOLMGdVVe4UWzPhhH+Q5/3TFXk
2hpiZWDGbp+pHh3wsj4qratRU9NPk9OicyPx3m83exzZr9E6g83WRzM2QyGd
Z7CoFuZSXac70NH1e4UzcxszoLEkhmnZ0sJ0r+iqhAXUDL3ntjNn0yFTxPp6
tr8bsTTISVW31dJM2bUsNaB+kFhNSGjUgf+h0x8bWj0PU2IeuBV57zt6Ktoh
NCUEIrIeRGFowC7VIlSTNbqwXV+An8Rxmwk04UX9eWHmXJl4hUPvJ+EdO2gQ
aSa4DnisIR/u7TcE9sieBdbZlU01oLAAuKDTvrd6zPYsPmotjVqQzHeItLOX
e6iID6ZCk2V7jIFYqD/P/YOf3QePjh3wh+FJDLD8UXtc6S+PH4DlEBdCJEaC
1CUWXmvAzqxe325RlvZgwjnpJylQJD8JsfP0f1FmMO5xFwNwLGk4FCo2fdV/
tBdYR/PTqazmhe98R/9NmHeAuDU4OAG7yUk88B1Clsh2cjjB2+4/zs5JkdeR
tEHRuSFUqGVw9KnOs40UUmZQXNIEZLgP+/uSIrUwFR+4T6zWepSxYiLNQ9DD
5hpFdnpsJbX9F9rZ7HpzsLRduMc0M/XqahI0crg9OmDLdUkSKsxCzNnh4/6f
ragFBgyNUjirmCvx7vOcfGfmg9p5/NJndsDZJcfLCvuoUJM9V0Gtt8fmlaIY
bR/dKdSYg05YI8fuH41SYTZ01TDbhHU1rIfHUAKX97j79Zq36AAhVwa7L9R3
dvn6OjBVOpKZDJ1asdHElVmi4RbVFpZ2HgHWTtSrzyEF3pjedEwZVA77VkHv
kosGpdhuXhKoBgsQB/Uh4bzZ4IOAPX9U8PBgxZ1ZzLZpDCGrKXE2OCdn5sjL
vOTwcuPxZhdSYYM0YTM1YalDJ1XwV94CMAQ8pXvQysDEzoUWgal1ruHzs4Qt
q67Z34/rjf6LHxdqZUn/iYFEUyBk7aBibXgJGa4dS4fcx4KiwPB4TNIL4rPE
SjA9O+EL0JqKAQtunTy+ILzo1DI/QYbXD5Zy2r0slkDk0SobVtTGaETYAORq
zsN/E4e9ffLEZVuzK5iD+OGWA7H/5o6tiAFoQjDFhj6TKsCKRfE7v513Xrrc
rXcpPvaD9J8JmkjTdv0SknFAj22JjH0ucKJw0+7s9227iMZ0XIxRduQGYRZ9
+SgrWTje9Aa3B9c/qcHfUNns6TLUJVHz7MB6eFk7APNyISszOAtdbKn7ZLkO
zLZQ1kwhUzKEygdH6NKwSENE6aG3NnZK4YvW9ai8eYe2RPAfYGkbXjRKYGQA
BFIDhCZa9Kv7rU4xsXjHOHGUAQkylqTDX9YOjKaT8zCIyW2IZsdBF7DEofq6
RShAPWddUAlxVzF7fvH4WYGFEpHree/sJfamgb3T7BmkCjuLMaBApzogw75y
JaLqEcfkhiPG9LwFAxOy1fYinAcy5DK0vv6FHK95CP8lVWmv0BIZvxA7ERRT
+8Hc+AVkLiqV3LCyCoQykkwPGxyQl9T6yRfDFEoLM2TWBmqvwDMW32i3QL9R
idBWoHJiseJXe8jAcKoNKH31ZXmC3rlafwrvwBcuuulVa/CTJtQnYPeWPJuh
DOroat7cju41r6aLUfIUcqJOpB03ibxoENDrFYbNSkTpPuyIdCjSeYwSAr4M
BZONz6uXYt0tiGw+uWnSEK2igKg7mXlmyEADzoCE8DSP3BXrqdq3RObrFG91
NrHXS1k/UCSAk7nyvVhDVsLX4k9JxQN395GpBQm0FXA9mSQjyjtOY3Svos6+
xvczRFAbo1xqV4C+jUsdYQzJindzR4hrujWCE75M7tdn0HYYzEdVzQCSO+Hr
8+Q1xxbuMI5zH2qddAo1RKGXzQn7fx5EJNrjN1G91aKWezrvFHCSpOL8B8cq
CtvKIBUrKQ5IuURGisd22TQSMs33tX6zWWACpwZloylsN+1QAbvRwae1qf9T
yQJD+03o7dEXR8X7wJ0XFEbKqJHHvVWErC/dxMoekc8q40aWS7fWpVQunCF3
BkxDyfdMje05jYYkLQLLy+s+ExXrdwnkvN6bagzv8vpij9AsJBEUqj7j+KKu
g/2uvV7HDOsBXL0yR4dPH+bs121eLc+LYSeDaVFYoYux4Mol3JtQRib4zVCd
ctcgRRyUYW71IBU00YjkzYJDKsumxknuopxqpK2/3moOsoTmBw1x74H9F22n
R75FDRXA6Lt9/wGCPugDZw/04ZTwIxiRfDMvkcssQ8IP09tY8GhiKU+1IJUR
RdoU0RQ4TYtDBLO3AaDe+PMjvpOTlwU55EqsSxkDZ8w3KvRStgZCMCUF+WUf
t1id49/44gZkqHd+5mt3K7HKsuU+gD6DYp0zYUV3trGGlf9yiaENu9Iqcv8U
o2cY6SgE37qeSxLKQO/hS4G66d+6uz0dZg2xzNtvSdmoucbe9sGuCwXv+HdZ
3hmDmwDAEBHCsD/28uQm4v5OvmYxKoLXlW3zN6b/1DnPWNrJQifDr+MnXE0J
OQkiYR5HF4XErCMwBN0+crgWhRnlIkkwleeq82LqC2AEhCXEVsRJozrxI8bG
NWatXCoVhUzMJGVZjEHHMK3mU1S6xqc62zeO1rA6hpsv2S9AERJbGMbZiukX
/QT7CGKNvt++hAnwX3BIJGiEySbfygQISsvyimaWp3vhhAKSYNZZjChiZhM2
zswi1GZhjZZpz5JLN06TWm837pkjkUtCB5mSIjCcwdSbuCOBkfloiha+j9Zw
1o2lWaZ/c0m76VRVZPeaAfzv04a5EgB2AORsjdKplvdp83yhAJZ5mERa1anz
BAwMDyIDcuWPCj8bkGBEfTe5ieaxKTB/PJmOruaP4eL1IHGGznGB7+59PkMp
F3sdoW/cgzVb/iQrm5UG+ddo/J0mR087bqX9tNBL5rhqb4RO72jaHbnsJIPC
SgB31wnX+3nOSfE4NVJY9Q0bIFT9/sdYLLlP1HSFOwQTppKoJcTEtV3UAqsI
okKbs/t9ZsIs4EcHUIw4XoZgNfQQTX2dUlX4X5ZA+9YLApud421PDV4mYEc/
s74lVzRVFycDiE8HHXR7qzmus0JK6DPGtY7kyqbY4GDStvpASZY+kxA6sji9
eSgneAp7b/bdjB8x2Nx848KAFPoTlS4pr9Bjuh4eyEmJyg+/LJo8txOgu7xU
QccH+BfN0ROe6NXbcmYg4VrL/lD7y+6isbozsIE9gidvnw/km78qqzg6MUgP
3j7/ps302ewlPEuvmmGEQG/r3cGzQ2BnOdhSqvRcSDMyzEHZvQmy0vSACAWR
l3zQuxu9dLroocvu1IXOeNTmTGNZiDkZrts7g7qacd2TtJ+Cmhr3ylhEgnOh
58OyfO6DeyKze5VcuCT7WlZGmWZZGSuS9+HWdOApKli0lkvHQpMr4TG+kx6K
dozpNZDFOVuhmZkMESA2ceyeiB1rvBaVXRYxLoVa5NP7bt9/z7Aj7eS1kVTT
lrG3cKuRsLfqcKqMpVmsBS3g1vRZSs7ahSolP1/RAnmcpU74XfR6tnlmuHuZ
JOUf5aWWQ2DSQEP6O/qK9Dehg1kKeskgRUHq6104lZtiE9PxMlsy2GodmZMU
zDX+1LbA532TsiNTcWMYj7geYbpH81uUz/BQAxCiqM58aEwXycsf1iW3o7gE
6lEv5uKEGCRSuB6bOtX41inVroSwWLf4v27eMc+R9HgbqxtGVe3MZuFLVhas
CjrBNAlPCu6BIxqNQMWkP3SyIHs1vCrlX3JhC9jIdb8cDHno/tAbD0RHWSRU
fnc/CJ5/jjFMGLyrZmmxiwKcV9LXFAd5dqQVcxC6RoNGE+UA/HUwk6Enw3M4
IRJRvO0F3PoyeOlqcyQstvhp2yPaL1FSF/kvYBR6BdGJynsG5Jkd6A2pWQ76
e1t9TU3DwBPPLksVSMaOyQu0GFSPXsQltuHm452TT0o6bsZAW6Igy9LdQQ42
Ir8KM9UjATWt3Gr2p6Yp6XrVXMzcRF7hDmSG92QFThCVsiVL2rMzMSGNx7yK
Xlve9koHrlzfUwDCN5delAqS1qNDA81zOt3h3RBbDMuamvDP0hskAcMiybW4
q/oo8S2gk7xug4OBqTBQs5XsOCHGikHLZ7DJKwlrlgBKnOgzQfYNn2CroA8b
Wp9CGqv9RsDmn++lkU3ahlJyprhuO/C9WD7shfb5ZqUa2gMlMUgQ252c0//u
UHf7CulZG1Ubl59MFOjuKXfwGUXYhkdKd8qqG7krevxZTiZI90u+ilZCSEPf
NWCy/0boq1LU4hH7FlHqC2qyLKr3JeC0v25aF2FR8QuNiVWmIICKsJcWS4jT
Rceeey4JHoRrHOqsKdgQywmLqTFomEnkHKCqdlsrr0WEGeaAZFZopeSqD4Cm
mfZ6s4VrY+caRv/heHDxQNXmVcFLe2CAd7da6xQwAqRfkdMyVYThrbJtpuOp
RmakoNa0cazAkUJ3pZO9aUYx4NHue73x+j3EjhyXoCAB3IjqAwVNTZ5i5Cx4
BOVlU8lCC3Pufvv7CX0AxpbYGtlHfphCYfq7C4j1Tbf8+vZJVvGBmUKEbI5o
sHEbrvQ0GdMTkFOB3Yq6XvKqfyCs6lzeVaHhlJIUM6BSIvcEcK4MOfnrQMxM
3aAOl5Zg/vBzTitkY16s7xcJ/EpShbAPZAxOIxq0aPOi3UkgxBBgwTYpG+ak
+ZJZxcEEKWbTqji1u9Aw9gFNe+XwMmgpzU685jtjmrFkXcm+egAuyCAw2kne
OUO4BD8YIX5UKq1tdrUiWPITsSV1lQLMKILMYERwJW5BvQm3gONkoKFC6L2w
K/1RllWgS4Ick5VxjRIHGfBYj5RgSNlPDpl70Z2W4nlLM8r/EhRBftDltVlb
y2j3WvahObqYxIXWHF49XY4FB8vZ4bd+Hs4AoNpQKSwQ+8JNwJ+aqTDJZa5S
Kte4yPWYEtE+p7g21QNUe8Uacjm0qtC4/mzcE4r4fneJpYzBld4vMOuSsUsB
Sg8T2L+C0Fb9815g8xVf0u6AcZGBaRa1rgQcKQGofjO0wj1ynnHlgE8w+M2U
XGps2P6bMdpnvuuKBuycR9yYBIF+XXCzgj7cswUnYFqK9BwERynjpnf9JYa/
GcednwqlcH2vWSTo9S04vhOJmfNfTYG0VIhK1KrWd8YbCkCkByH16ZizjCeg
ggHb63aLp90Js2AgShk6T0Zg7BOXGVm8M+bG1l6bszQCKd4nfAqb6W6jxoaX
Jgs72aSj+FnKGrL9U6TouJ+QSRUNt8vLPB5399HyQW7gYu0j9JT0R+aBI/3n
JlPrfTIG9bZ/IIB2XpcqlwIICdyWjfRg6l0mlQXc8ouC/g64BPUbL437Y9fk
7loyHViRogNOL5+r0IHV039nnuwCqPSZiI+zWF4HGfzkOQ7BekUIsGUw+3aA
BlatvAiBFzouG/qvD+1sc8/BPHjxgQTKAJtiXXP6FMBkcQ2OiQi8h775ek+E
TlQ6TJzU8pgvNQKlqNjWWEjvOVfkRNUnUN3XoOh6I13sOSt7573sptUY3fjG
+pmk3WUdU57EIEpGcvMEDSpwiHPh44XsKIrbsNllJy+6WNzMV+R2G/u67C7b
StaVv/HEIjCRqamZlI2xUPbbBxNVk6+E6gcB+sroRdLmy/+bPpfIkRY0Frwf
IUIIRvgZv/6zY5FZsUAEG3fow4vRpYrz1vv0/MebVMCXMK0QMEYihopMl3pO
wlMoBwR3ZrS2l/+SaLEL78HjbG8lo477zSg+DhNcU2pGf06ligouM1hEwjhP
I0TiwOZUQHgLAwPRs6RhnGvwGdqWAEpsTFuVnJbuwfS/2xVe4hIG2JV6mJeu
SUTzZbkgq06W2++3RoY7W+bg8Ma6y91rS0ZZnbSSpUwDrq9ve2RHTl5sy31/
TZDGSZkfJWIHxH0RYdgAcaBtGbvQRW3VrZxgsuOQYgGHcRH1SZ6elB5ukEmW
/A5OcRWSlDDlbEyaT3i/WccBVHpo6oupE2MkCOeoBpDedQCQP9IXkeAK0OBd
O+3xtSetx+8qfImtN10jlH3Bx3Olf7GxwkTUZ7evoWOzZOmzeropU4K8ChAz
Ku9Oba3cdGypTYND2Esm6r3h0NtFaLWJXHJRj5R77syodUrMBYIT1/M6+KLa
RH1rkbB+3UD+N+m0w9gdG6a9maf4v50gEMejy77h5D+2Ih1ti+Yem0Ll5Ys7
WYNVCRHuc2IqE8QTSkzUOxOB27IVcNIW867jNby5WJAz35C0UZTg3j5RWNuz
GOEpMx1E7FZwv4JbG37jcZjP9vElD8/+CJBktyYSaDnkvLoYqFvS1aArKdtP
XcbG09YT6r6yH8WcQojhzpbWc7IhLOqawD9OTq08LSbirCALOqfnOOH4lgK6
wotxIQ3L0SMCudl8ZztnBUBmJBiXNHH+A6qADAIgpKDQNzpBu52VZMYuaNJQ
6c5h6du9xBOUckJYAmu4SGD0+9FrF5oqkYY29sNhINVPSmokyfONfT8y5JKL
1G52k00zvp0lEWoYKAN5qOxGuvDzRPKKu4LaBegKBj7XYAUW0vK78umbCTGZ
SiqDTJSVZp8S1QNnG/zGicygRNzfHDj+yHYOhVxCFvQyA/Q5owXWWVbFVh4T
fGC4qNCbeSkCweVW8aEZDCl2Ge873UY68ghENNLDyYQrhjUedIEUqs+fwc8k
tiqaZzDB3WV3xDE81102HkXRpWCty0XE5va0GF7Zg5tuptKx+DBRlrOsTcpg
cnx71K7c/fxQyfTECSK0+t8BlECXqEbxVQ2SvaCqGMBCu+0wz2vDJ2xdtXPc
va+eaWeXVOnoeHJNgzhCGqEgRmp8SG8GjnP7HDa0SkmzjpOJUxgWU0qqmbBV
X4h/P4qXdTeneE+69c4hvW+zfdRy4HbvGCHkNbGl3IxgfI640mO5dP/jgY9U
/9jnkBIzLmstybJSWnRmTPpk888ctwUHO3O3b9pagZ8MjCjWLdjPr44Pkt9c
0B3rpI2AQ/9FXq/0yGiHQ3qyJZMlpMXZwbi6uHRjjvMw5VwRYAcz3ffvtIwz
gIfERmXp0c0+IFfEw6U/vMzPbzuVCJYe4FNTVF1+U25TT2y5/43T/B1bbv9v
L3lK8u/OKn32C/yVLMS1ufDDJG7tFWClJK4AfLs1ggwnuJh1U/GjciSOgSxl
8YM65C4FpaB0SxqOI017tGFWeCpr5lrpV/db4pP7ZHF7aZzs4wy0xTn8Rd7Z
yW0VMa5kkkceAuYG2pBnEKEMSU6fEm0byR56Yomb03U4XW3hEbJJxOGXyLLR
obQiyrRvQ/w+VMGdivzguzPOJ6HdQO+nQcge6BQ5Fw/cgfZb3FpncfC+brgn
k0z93ugPKRXEoubSQuS3f8BJRFHfKfrm+6hvCKsSfycCQaZBzCDdNGYzd78x
kWmIN9n+nlzUIH9D0vMtPva226CoQi4i4YLKsppnUI2ODkIV8+1BPoaD92im
WY+AYT5emKBQAfEKLhegZR8lIej7soerOoK2fPAx0vxPigT0U8JkeFzFLnAE
41UybvHAAnGufpF/BSCRR7l8RlZNMXeqnjW2ob6zbW506LdAe3jSUnYs8ty8
5pXww4ajd2wH+8xEKkC9MRMd9a+Ug5fI7SfmS3j36jMpIBlQrrfwsfzT5Q3R
9IyriEZmRMJQo0/HfpO8mBTPVw5+/CaZe8DtHm2R+mP4KTYZm0Fk3BPnqbcr
0ZV3j3p7QPKrJCRV2UIfiUB95+UIk3tSZCbUy8i3BrVmhtI1+DDs22hN20QY
G8nz4KgjBZ8iFE3/+arCB+CzHX49HVp+04vd4XwNsM4uu04DKDbOIGAjW4kG
ykiKawuHaTczWa+Tv0chFgDeguPMU5YU5N3X+/mj70pE0WbM08gktDTLgFGn
vQBpJwvL/Nlfw9PYTzcp0jbkvnfPP8LdYA24cPrnf56QiZUJ2/eji8P3eDem
IELBohXzGIznyZ31zfqhXuGAEtkeGmFYv3s+StQrtVRXlS2Y123rcrWyI/1K
xj4mtJEbKmTvKS9jaYzxGjRlPZzrcvE9kY+eB6LswFnHcSboRjfB+NRfDFS/
Uar1fS+rkuu/CYX37fogite4e7+w6xUeMaxNW5AQIoUHQh58SSPctJx0vQsx
sRTjKyxP9NvLSPJpQqwINu9jI57+4xx1GreYr4r/3ndjzN5mwoXYnUBQYIv8
gF/WvaJOOvC28wYMH3O0YsRgJIW81efQxgDfHUBnvSf8fIyy/9uDQF+AnTX2
E5O3Zx3R//ISrCXBpLFOS2JfOAuysG31knDBGL91oibeAYjCdytRpCWJ3aIw
QTWUaCJbqEauIdtwnKIxn1mH+rsdDS40XJBV9qDPB2IlJHiPxPCo010lztjq
aR/PB8QnbJpvHs3sFndx1PSqdDogI2l9asoRXP2wGZYi1HDD+i0ZlYJ9HbuU
xzQQ6MKHk7Ro7XckBKRXf9e6qQ01FGD1w73aZ6u0nYMev+MSJ8Uxsgq+kz97
IdPn0+tLytIaM5tAfRFJIiZvEIGs8M7Q5zxeESTk3s+SxJk/eL0/2EEK9Zrz
wbNfKZLMxGrOpL5Urim3f+sjWh1gThN9EEBwzA9OWP/SgdjuRVxHYMXsIrgh
Ce669g7NALCn/svcXYP0TgYUhk6MyiFuczoIE8/R1iPu29kPqYsFX3qfZXGN
2Qi3QrGiOk5B94/ffLOSEbmA5DmSzEjEmCBheosW1iFRAp6GNICR7udxLWVm
gESMfg/Cz1QJTdCU2RQpnAv7W7BeCljeAF2iyaA2iC9uUMj+gOpKhqB8JoC0
9nYO1q02OBZ5urer2iHXNXQhyVm9lsXFtCkT4UOJD80lmi3FHnQoZzj2XarP
vQwKFZIf1ysLocnumjgafeI6dPOP3khtFrvoA+whDKGQxXxewdFzohR+HBTd
9lwylseACxgTzgXnU/CCD6gmmbrqV6Ku4svpJYt0OZgEd11D7xsg+Dnskzyh
TIXflVH0eMeOD4KSUuc7dM8jKwHTDN975zXTA6BirynMzmhZvBb8zLxkAK2a
RdO28e20NSJHOjm2MzlbTSeIOCbxWBUQSW8tepznSL9zvs6QAnEUJfPfQxDi
han0niBtzSeF6D47yoCjElZbgZJ8GkMUjfLpIGbcL4IIRmsBG8Vzasseqoc+
mfyu/PZyY2RbUICP1X+UEPPVLhErzcAowbpyhCach5LlImTgoiV7lJWPzLIZ
YVw9dXexqlBjNQWtAPR142PZf1v93Tq4PRt/YpNS52ziZLU43+wWZHtqwUlB
52Sy421bKUS38SyLd90nRds71MLE7j8qlZZ/d/Dr5HOWCmSFQqfEZn5hdQn2
6gHaaqqjKwBbkX98jPZ2brYfqymv5aEjsC63pzeJQTXWg+7lpkbILgaLnttb
Y8veWhLseDZlgr+lbiF/Ar/K5Z/YGrZLg+fFhsz9YYFExdBo7annHGm9EXfO
/CnGKl4q88UEJ3+jXMgKlliiO34lIt7zO23LITcXHy1euJ+pEbl7VFKweR6H
CZgcSc2B7ExsP3HIbczdM17Bg0hbuIcbwVr91q4pxOUiCQTVH8vYyiWeh89/
ASS0gW184nOII/xMf1UKsOY4S/UhLqFdmV8kZY9V+L1GEz0DY99REHLQXx2a
xSupGUKgJW3VT14M82XjLNSwwYHOe4KzqeXLa7wYDLfmg3I9zB3zsVK6CmvC
rqXtLMrFX3XEYq7hmoYJCyjyFi5xOA/WoailugY6mCvuAspT8kYooNzmq/qc
F/xAaF0HUtLzni+GbOdP7E2XmDwXYYrDO0Ic+L0I1Vp0xAftHXFpGCsOYeEs
QUnfGckyRrirotglgL9Ltz4H+l0hCjY+vkngBOLCS7m9H2I551aMw9f4Fjly
mT8OvPwNd/j0ngBGypIQsAcZQ8flexjzQPUM5YHys4Byn+9K7n9nlMlQnYaN
tFuLnujxkLIMeCCo3H5qnmkFmH02TyOWRscGxoAELkMbi9Nu2NEtXmEKk2Pd
OF4r86uIgcFA9mZ2ZLLva/q6ugxDIFQ1lR5WxOPjA9hsQXY9CWNH8wx+NZtY
JbB2PmEDnRepCmRS/gbpZWMXEPumWzql92ZQrpc3DoSHjyW7Nchb7cXZpFI2
7N+VlrfBvsDRRQjc1KXFa73A5GL5mUVZo0SQzGWU6PEb5hbeMMuWQ640cbYb
mCxUVyK2tAHHW9f+t5nBYteHub6f3huO/JyxX59b9tI9r11uUGxhiaUByuzM
tV1/m0upslqeqWuCWBMIiW+4hIp2XqnVbUsqfv3zxx0gCISfUH2tgTydk0Qm
W/GKLvCB4NZgX7KLkchiP8TiM6mYhOcddCBZlBVDc01bl6KAMwd/Hfu2JovE
0eTav9BaCp5poqypNHiLfyL0yVpm/U+LsYUTvkuttQCLP3rJaSc16He3J9YQ
Etm/+5CAE6kPr8GfMXzIOWUvtdPKd5iH6kplECqnF0MAcK8EEtaIp7TmiG8U
UVs0lhMC0uFyl/DXhgML81G1Zg4EGgBB75U7f7YCg1a8f52STaDzjSmGNGcq
Eh+3/Cqnj43gvpkC3ErfhJXEUs8+vCB2t4/zh9Pt9nbtV9jA+25vwLF4iCn7
8iUxwBC+izDIPlbgNmhs2aLeFdQHW5pdaTwiU9D85rShEHq1f3V8Aur7fkBV
NQpyw875/euPIEZDarZGZMi/qKzEEWbZ+6lPxINJ0Dpt1WJSpN1bx6B9pSD6
0NWzKgsADJHHO3fZOP5gl1VrDEN7XJCPAkOQ73sJOg6mpNzertyC6ctQQRGA
W43G1E2TGjdPw+inPFybLx3eOMqeVEMWhvnKN26yY3KYz7OnA52gGcTrpNXH
8DIUhAE3NTtg+uKrrgZJWtMSPB90dCpLrQHVxMIpLTFtD/lSjCshmOXvqscH
Zl6NoTyvwkufEvcJpqQs8ETqCEqNs+gWiaaQSW2AyQcqDp5WEKUH7NHkJNoW
/OY9RjTPZVUbXHxnRlJF3fnzuao387V3EDvSyA3DDyRMyr7Luc90n/1neceH
89J7fNJsrahujMASa3T9vBSCyF95Qcj/vUU3Z2zAtAHZ4dHNkjijsn2s4wZ8
UH7FXcFMX6/RxBrB8DJK8uIppBVWH51LnVW2Nf3pzHCckWo0eHKKkZc/Hdl1
teFDoamd1XoqlN73j1TIgbvH9gGsQfPukEzLZAFdKfM/wrVzSscXdctOx5JC
ldwXw+vPo0rOFbPyQyn4stf5kryRRPLDigaxov9K3VuSaz+HdFPG2DKxyHPr
jO/uCf/NkxDjE/g8tEQ7QrPIA5JGWaqOS8g7JGNePBRSBmMVprXUYlzVC92W
jIULGdoJGf5bKaZ5WxCymQhmG9BXuJcRSuv2cFTiBVS7E/1JRYHQaNAakAop
6ONHM6AKOEYk6sZxuABeyp/EI5ewvrL2VzepHU0UrgCpEutW21HAAC3UfSVA
p4zAlRAM02ZNFyZjO7boVavQEH2DFpN0B4+wL5P5XcgOvmSZ4PXMVGBhcSCW
9Hv5NaQLeKqPJ4nlcOgbgsxsuiOVWv1EhEbmRebopc+tdZYbIIA4k6i88GS1
ecLoyMai4rywC2jQyqHOSoPc4TcADaVTjTbJYaFtFnHJoo4ygqpqUyfyPAr7
7gNyqve+BqekG6XUgfNZytTdqeMhqPLAPP/QPgKUxYV/nhS10AW2m1W3sSOR
XlbC7CPNbKSza8yrJE60at1mDpHNHBL528/muaDz77VhX4INajLCbrhJhgMY
0Xq1OSB7JQuzoPsnRTJhOQebig6CSx0KHL7hOA07cRZlGEFwZI5n2X6ZJ79P
gLg4iVlPKLJ2ACm/qumpMJKKEZBtwjO3Qj5En9E+Dgtyh7Wp+YuwMHign7AT
UhLOiGJrXr4Ew6ETHmHwsoxvcI9pahdeUNFV0igIziUaJ/umu4y9ra2TTXSt
uoxDPUMzV8G+3DIGkTax+IBgdvCvW3W/rQEgEHYpgDSFAGlDeSfB4/YDpMWP
p2AgT+MT/v+LKp2PGvd5Pe0CruelzngDX/Vdte4HVV8X3uXMwL91ClMpHj0n
8WcR+DKc387LEqFX1wwGkil2iAKCLJjq+SAfIk2cbPfuvRcBsdZbLFXZOY1Z
ykpcWGIaqHvLT2oQGD89afIZb/qFFEbF8DJOnY0hWPYAwcXF3ckFksPknPpj
c3x8SYkU/xrMByYw1OFvHXk+TL0Lz4ygtz8R11j8tN/g6FRDKhT7auKmIMFD
4b8K2jtx5IvqWFX/86VQ75rrxpRewz6elRF+egfAZWUMlTbsylQthZPwhujM
4amDkU4Ne7VixTiNx+Z/nuwKVhXgHcZUwO0kUB0cx0BxJLtzYM38J20rJt0N
4HG/DZrL2B9GQFwvntRPkMn8HqeEnlhSqSvXd3jJb7YEns119/AL3NW3jcOI
bJBGuPTawNQd0sfbbfKyuxfe6M2WMbQnwj3w5hEKVWz6MMkIHXExuOndj7iO
U2InHbti5NeWv39n8henTHszs54F8KoCesaFkzSoIznJUxgEn3DjWIr59qWp
EyjZ3fYMPq4kK2p/uvil1kji5VXcqkjW7hZCe4Jm1K7VhpzdnRZkzzRh7YWc
6CYj6JDFWwj59iechk2zOltpwf1XIo4gDIfzY5/zxwHL0SAwHWusAEmpRbA6
S3l+A/Z4gIaxheobnZje+2NFL1b/UQrXMRhaHcHk+brUpqhBADe87VtabONB
5q+QMa2sH8GdKK4w/4q271avbKprY6uXglYpne30lYh7+ylgjjxq/MjCwGeZ
AHSWkZZ2Nvku58KttA8QqYdDx+8Paj1VcVOpjN2ROG6iZGCxCjz/8MTR5nKQ
dJ9r3RP0xGav99Xj2yRfo4u3XE2UITJIvJW+uTaw1KzMlXo+zHEtNgz9k+24
ohcXY4YEJnjIfXWlFWGKwKLaZwViWQZoCJh/lbif8gNYTC7b5o+JZ/AK9dfL
CfkaVpiF7Aquw6SWzhilppV1/86LOb8j4wCRQufM7yE4vp0OyqBE3vsgQA7g
kQid2p3Xi6DHIUXK7zRpshghXRZ4e4SxfogJIxDd9j0VCYlTu1eOTbOdhUdn
Z2bkUkQQ7SwIVQwQl6Y9kRVahrnzCUoln2ZrI5JRWBuh+gCPHTEHh8d98GrX
ra/6iWUjXRlq3cKPzLJBzxSOx016URjv/AiE4IgPg1ndXKe2bN04vkhVhjAe
bF16hESV1UgGer8Cv5hkvCZvHlwXwZHs18Ufv/rzSR4RhvJd2VNLvTMxV7pz
o4j41c4jh/lAkecsN1al49rqAKy/Hxi5Bp6773z+IkhPT4AEwjgP/f9Iz4W0
enohcrXt2Ozr2hj0C46XQXa4w6OvfCE3UZft4znQyRqV8tSPQLAOpWZLLqU0
Z/nKb7RzwLKC+iJnGglzTJLL9Q6tP49fmwe3J2aEyCNdfLbCjpHYCzEZLdCo
tqE3WHvCUPqivUn04JvRbTcFCQfij+2/+LmTjb5sd0smLmD8NyKAptl2STP5
ZCmizb0twHz75sfLrnw0aFK8zfiXut0lrWe06NL2XImPlrwyjtQwA1IxYBgK
AVQ0CpnjWUBs/6qQKXQ0as+ZnvFmeji5/t9aXZA+FzY+WWeTGXjKS01oznR7
mCJqVcdOkOT07nJ6cvpyZGGURzXOp1dm9sc5cjVy1ixLOIB4ZI4jGuyOsFbi
rmyCdwvorIMghlkmISxSitVChcCKNrynu0gCrFJcfTHx6oK3o2A1lalARtDk
DmqS+smlxZiJrqtTLM3Z2jSLQ8T2EuZJh47Rvj43948jQ580pGu1fY9QmBeh
Vdur8kfz+X/Xjd0K4jgavGe80MWmlfAOT8euP3caMAUmGLwwPWCmxnSRrgPD
9mEEBZWNKH2LqDI1OaZE74mnxi1buuf8RXloCXbUQ75XisLr1+TQ+T7hKri0
pUNQ8falsG3rKdScx/m/aV6KQuDpBAXYrsNjPG4SQNRJ671fO6+Q4GGpqRDn
Q4TW89sB7Nbec9U33c9Y+GvaoB1j6aOeHuxJHI61nkx0vgXoYA6v0QkyGBjN
H2wyz4ZUMltQINIdWComWjdqKvoOwdsK+4ZaucuLbfClcVSuNCwaKIQGpjYc
Qvv01FoU7Rtj5Mg1hawFMGghpvROpDUVh2MReztdSdTPk/sAg6/TTwFLZ2m8
rc9NsT3qBTCGJSExinMpSw/5jIGeYrR8lfEJgsBfaNlvltWHHH79bhv1Syc/
BNZeBeR/3+6t6CZpi/8AC98x/Rjo/StvQ5ZxueRWffOxB4mVDkZSAPG07t+o
MBBs6cTF6H6QTEHrbRDZuUtVm/25oH1xLESaqJJLtQn71bQ5YXTgEOxo3+s5
HxiKPxdrHh+Y1G6Hwr5jvTUr7OWCr/MbO/vluJBNSFWY1MQPZJdbwQ77Z6F9
H54xZKkoL3dVmXy+wPI7g5wnoR437Vr00vPHmDdDN+z4vb2T80BbhikismAL
G0Qwqyep3PYfcGzN6Wfkp9lZdpcZ21w27cpt7EO4RIeELYC40m4ff+qZyHj1
BRvL0GkeSbzzXM6OIeDculpmzdORRlRTvKja6/t86bwS8jgyfNaEBNhzqgsZ
1zg1X6q6lKlzbSRGqnXATCb+FNOOfU7UpPD76MRZbm788vFNQeuV2qXaWLaE
MVmC7qOi+k95tlzm0cLZxLXS89KZLDToN6tJDy77PGF7tgFthIYd8xfC8G4C
0y53Dt+gAO3/mw54HNCsD3VK9HmNGAcKB6bQeBbpyxQbZYNeQCTyB0QG+WrJ
u1FEad/LKS0PWC1xYkroWI94vbBcED2AXALk5kITEeK4VNT4tvjVqMsg9cdv
BfJxQsByZrNrmpsTItnrCxSfLhWl3te8T0USe1zYiBKRRIJFPMC+FhF/9CB4
qT6dqbtSuIKXplsPpQxrz8OJmFrTFY6IW2qQGOfYgxrQsD3P2g1KjIYSVd7D
qSjcY6MrM0DOzpaxs/3vdBvioAfM5s49VqapYEK4p13mmobAI1hvGL2Ydwkc
vXYP8JayqsHkICBRdFU8I2bZ7+w8sIqwaB/duK+QZTIVCa4B/GMafE5cYUB6
ldw7E4TFDU6L66dTuunqfcZbLvZbwVcYEKEwlOGxuGv3r3F+OINVR3YeztqZ
AVA3cwekuE7E4Msmc41+MiLZqqbLZiuF7YcgbtlATKm1Mk476iio0b5Bul5S
H5LzlGgb7WPoq4XgEt+jSd/BOPnGY5erIOTv+aUrdkRPhoahZ/QxqQa4xGWD
yHC6Y6exyflND5u8CW+tMr5e9dN676NLf0xeap9aXUDlgMfDncFxcZ57vcUY
CrlNfNprths/ZHFUrwzJaloTja0E9Zp+Qz0nrj+cI+BE5MLO5XkAP4RjVpSL
G0PoaNpbRJYdG24YaQQZpKhfh2RxpoDsKr+MLY3EJk3VokwjxietqoZ8hLbv
dVhfbVNJgBiljlo1xgtgIcGgAAxID4445GxiBqlDoApLvZBKM6lrIKEOagPx
q5wwBjKUl6AqMtiBEm2MtefWAPc30PFO0fz7j/+MZd5WUsi8TEEKWxomHxya
eVpYGjoBajpKARxHKyjg7vpF4nieHDVdXTAe/GbWC0kuURye3E1cMUberyAL
X3w2XLBCXle0v/Cy8sTB2/MQZD7OsqgzcZtgn96sORwAbeHMQFRPo30bF51X
J18T2p72j7Xobm1HydRPAKT7zPbLaPztAmDAFRXX7iHOs1sNDGCdMWqn1jMd
9WqPMG8HM0Gu3mWLE0q/ow01sA+Ta+Nr8JjDBl64yCIQvVtHKq9xsthyLHFh
7AE8MalxRH11E4259Zrqify/bQ2C74O5DY3f0GHFulNbi0iQW0+tWTQn+Zgh
JK02PfbK3+k3ukYeggWhbtg1aumXOwjVyQEuRUeTat/yCYxk8LZsb7txuFdD
3C4mqNJCvRlTWkVt6Yfq3tGRRDsBrlz9v7W2AgOyQDNc6GhVI66AuxwjF0U5
Y6U4EOHFrCeZFCboBPOE4HEPjil7Mi5MKJmiIbjXVC0HfPpZW8vDPVCuyVwA
3z1SiIIucvZqq9buhxMrDqVKn8MJWuB3RlctXCS4nIqEAzyVKKJRUxNRpcnr
Yw8L78xDKOjENP5Jj3NtXfE3TTe8E7SV5iKvQZd/BhUu/yduMaaFsw3r28TB
NVqCJnZlqhQ6zSjblweCxoBWis5cmcySkUxpLNVhVm7/dAX+9TNO0P8NuAhA
MTJR8B3gIV/YOg49IqA8vmdY6NtAfdcrm9pSjJcyXOSdDBbbzTAiBNU8ZrSJ
eeHpDiEzTSfO+fNBHubMqYNbO7wJb96AI6tpjKWzCFWursn3C0hfnv3GOufs
ZYVVeUdfqXl2CYYaTEDAXY5hYMu/wGq/M74gZ11eFHicB66MsgBRiv5aK2EO
mUHAYrMDS0kpxyu0GiO4N+ATLZ1mXp3fFu51jr4SiT3lsBu7DvWd2I2L7VGP
gHWteZwR4gJtWifjxqxtdBWzFUN8wLK0XjKo+TBOvOMBcudjXBWbT8dIJDDv
Mqa6l53xKy1ybcn+87fSBodi6PJxoYxPM/pguRUoSIoAn+5CZk2hInvSA5FA
P34NjfKiW4wwQGskzV438M/ShTiVYeFEZbgIv2tB5V0oLhi8RKPXXIcFGI0P
/BWYIFSvW6N3tmQU2TBju5j4ywVnbXhju7ZjnQV1Ds4SWPUPYeY6YFO3bPea
/k6YULVrpme3txpSnruUsvO9r/rIu2aNsm6q93qvO5q/FDOHlDQiDVwacvR+
zWe5ghkruhrNOtrY6dqlaN+ox2RoS4LD+vPDNVCzYK9mh+LyYaP3McTgIkHo
7RgZA3iJJR3oC9TLDnpSoPo64hl5P3t0xnrOlzT9+7QvGwvVSh6x7jnoRAyj
8rI8BlP/HSMu6lD7CrwGjcnRi07UhtkNDtP3UAIBeycRQuRmruAeVEplZYDd
QFGH9c/LVulISMzipXO6Ma0L9CVuF9fH2XCuOTdrqt8vjSeN69Jq7ZKFCPPV
bPby+FVUMOudsSHalK7ulCAMzeYkOFjP9gOIG/A6Hu693RCG/g6loIGgV5re
InYM+MzlKEPsMRyLqO+lf6H+hZOCtIquedXsJOBRDPUweduhvrhw2dR5BkSd
bMAlCiVY363q0d78Sz167ZK+BcWbUycFkbi2m+dBsTfWli7Tlz8+jgH7IAtw
8oih+j58rctgDUnlSrd74Mvip+URCMQUwRuKoiAFZKSB/0O8ZuipT8z3jWUv
HmVYggS7OpgKUnx86NvNkw7fqiUEqdnAxeZEarjF54PGAmZV4oq6pJsLQZSM
ZYiBHcqFr4M4bmHoQV3MbPG3x7dZzq8v+5XDAuDRRxm2qBipZ8NXnvWHkUA1
BS4xrHD3u+OUjf38vH5qKx5P3MgR3zowibkg9XebuyuxTkb4ul9AP/FiJi43
HpHkLmfew6kSyE+Qf83xDFpKHTJPV9Pk5xtQFvdvtdaF20UYVL3K+QAmNQYl
Td2NkzdpJJattJw2QhNc0sp09IhsY//LSEX3vEg2AGDc1bp3VQ1X0g6AyAxn
C6ssC5VtmU1gZ77lBHYsLU7cPugx62bmSqr+RDX2U4cRqc6+VeZ2DgLRItse
YlJNhwxWlwLnNNxQLzLJg9mkgOXy61vHsslbMhaEdafeQL7ZGp0W6qVXFsb4
NoiuTmiJTvZS/FgAx7ZjXVU9YA1uXrOLooljsjjO86ZYvYZTDxAntyr3BnDo
phl38JtnKphPC57i5Ou9RPpvn+2a0E9aEgESPUPNaCPC4h+fVOf+3XB6Ykn0
jc8ISrsNaRScltIq7ifLZxnmCgDT03eVykrP/QT9DPQvOEnoBaU+RzI33y1s
AwlYdCjjVoRI8lbgdyIzxOL7cNOpjHhWPoFHm9W/VhS95sOjtqREJLhxWJfD
E/FxrfE60qFVxdQn2CQtbx2ADLB9194Rn+oRMSjsmEZCC6hqwCGhITMbwkfx
YoE7mjQb4S9OzSyG1cjPla2AFc6qUPRqXuW+PMRq6dBz6HYxj6HsME/fXxpa
HBIvsez4xL/HJJmlVB0QuJfeYJ6KSUa2le4P64tlGsn6jpN3jE2/+3bGE9Z5
BnZGHqcIWRBxyX5zd/H7hCdcoQGiF7EuRI29vzWy0yFEG8r67h44WYEcPvTz
lOQCU85AZj5R1CyGGu6/Lw6y+qnvGlfn2X/XhrOWF8NQWPlBYKsA4y/fW9/n
c7iaqDC6lWbJTY34TwaiZaYoBEF0YIlVfWb19hguFyOwkB+IFLK8hnfU0zpF
YfjGMPfGV0g6v4ywcDQfLVdL3hL5Jbyctvy6GHmQL0Vc0nHU+5KaEeQNUXGU
7hloR2xr5k1eCLxM0W/BIBR5jI+bnM/qAjFbZYJYiMPns/eOl9PPkd2BDEIB
okqiV+P3V6pO3ZVlNHRmKa5+pfxe73NQU9Srd2TowrkQonzkXH6H5qkh1cG4
rKY4RMphtcootWP6nJox+xvyeOsJHpi+zJgoKcYXF3cxW3mJxRSmi3aZBEsr
A6prRRVbFzrl/q8sg8u469E4bryMVv8XFe8NWcxox14RLb0sXuLNnU/HUTRG
yz5J/cIQynJ31Y6EMEDdE3jpMaYk51c889c3yFgwPGZkWZir5HPPBfY8pmO4
T+0UlqJ8ymxLXs4RFTmcyUFKRiMJ7SLwKAtakErpoY8cb9EPJmDE5zTD0tkd
BJsCcTlBaiST3xo/1mAYppzRwACDh9LIDjlSY/mamnmSoX3NRzzh4oa4BN9t
Yq2DqEnUR47q1Aq9o0N0fIa4dtC1y2HYmRb7RKpmDNIo5g8ZTTjzLadLfVFX
oeprRrZVTsne5DYvPWwnnDqybG5DsglQxAxqARLwickfLbV+6i8RcaQRIOti
9zTx+RgEAHxtETTSIp9zMH1mvOEi3j9ulQXKwA1MqdpLBhgIn6Z0hrPbbigH
EJzcQfZ5/B7L17+MpiUL8hFym0j2A8TnebDpBKU6ClkSdL1/jZXDKd0Dkdmk
IoLqifIpJ5YxDz0FAIc7ofL8DYKYlDgjX6LSS5F383ES9N4jEWL5Dn4G3uSf
MJHOZI/qA8PAdN6oev+oySM6fJMIP8aahSK3AIOL0H0AupwPJfnyFWRF3SM3
zwhbFOVS45npkroOHMpddM7cOe3qdiXeISyuaMMHS3nLYF2od+DAeINq17Xf
/2GqBFkbnl+fZ2Ca/GzvbH2LxdBrzf8Pzy9aSNd+rUjmrTRMco0NMesU83au
7/sUbCHbXS6T6mdb1FZVN/tfaiLzp9arbeuBYMp8H8gfiQGKAqJuc5ScIufA
/WLsg9ud4+jEoVQk/cVSFRD9WFo0g9TLeLUswQOORO/cFfhNbG09E+bTD5as
xxGjk1/emf7FXxz1TOzBlRRr8zTo2uTHHeCeqykELZzppYG9DnBSqKGevv7e
Bsl2h6Yau4DGPSN7T1GiQDUpZA4ETAddEBsmLYv8XpgES1+LWQiPoIxV6pOk
3O6zssDkQyydMaCJdmCIh3WbpdKq6zqbHlLBfijfHwcs9s7wIvYdddKP5Sjp
DsnZRKKLpdjFFyGFH52SBDZCE6vsAtDLXws8GcUKHqP4McYWx2ub2hkNhIzR
UtXiy10Zga+acwVoEMD8Ndc66UH1Jm+SNNmV9t3BqigG0+SewotElaawIb8J
tJRxLsKnf4NAAUVL+zk1coxKq9WMTjQRLM/GLADc7fLV1mI3Yrchhw++9MCL
s7EJAPqt+CBnQr5NNFbUTUC95icVihZhopnXocg033Z8LfIoGAtKznb816mq
mQu3tvkZeIxoS8SNal4oeVOfRYNOlR4EB5V6cJ8XLxGUH6AKnWQhLHz1xyrt
khstWW9Gzai6tev8WQkDCtjNlIR/cJGbj+XFzUjLuzktbTWD6rryh5dzp29A
hxsTB3R5EWniOhUrW1Qr5M500Lg2Ku0SIKR+GMAnnKvku750XT40wmwLnOAJ
iz+S8Kwb/DPxx8aCbhMQkzA0gYCcQVLK+MaY98T8AKy0+8BKS6epdxMFvIIH
zYewm97q/uHYRHnLGIgk6YSB8qqbAZGstlIPkgXHq/jedrIR5HHk/FPKYs13
WzZzxP3D8DFknP/upt9mSedE26Ow6R1wUIgEayK7CL7Tf1OAOOh4oJl3pcjV
ohQSGK1oepQOgf+S8syTvT99J5zWOBAaRgebIRxgqAAa4MkCVAnR5LKtEofy
8Zdsxtb0GkQ+ovLCRlHmiiSlXTZHEArkrfbm17wQ0pry9BmlifIBGNLJzI2O
CBmadg0pne7Y11kfqCDVnJTA696YMCX6GJObFt8rVVZQ6c9+49TB5OsBjpRU
DNWBRAGUi1F4wHVT6XEujGfxc6v9GgGfzfK6gmqVjgCcXdcRL/wi5itbjqLf
DsqZi43dhgKc02M4xbcpqHgEcvHs2PuEp4yC28Wjr41n2//1rOsFAK5okJp5
0T6mpcL7URfuvUnBTz3T99a7DLuNGPhD5ABorN4HX9Fo6X2MVtKRkwR0zW/2
cyHjyCE9TTeXobmTVFYzgVZ1RVfFqW4uDeAgVZI0Ak40w+EZbhRJ9pNRZbv8
MJCYnYYOn8nbZjDXI4XCGRlM7tZPS35UjKEek2q0bdlUSG4xZXvh34rOwNir
bxrPvHvGTtNSKpbosJluLjQ+oI+29s+N7wS9APQ1hTB2t2O7QBLeIotTVvuf
2MWOCsCBCnACzL3zCk4JWHRPdsAkqmVjwN8X7Tai2+BzCKdk/EXb026PULVm
rYt5T6AJCrI8V3yFMQZxFBstw7VpghptHuuVaYeZ3Nbj8EIZ6IHiux68wsih
rmIynPO+BQGQYEKQZUpgnV1xkPqhePGE1KRorfovIeSUeQYuOM9Hyf4LWnfT
3AMGZC5qZm7GvKByiQWBWLCzxoEA3CmQf0BXaXnxGfK8txOj6Tj6QGGYYvNr
uOPZc0y6VCWwpEY2ykovZdDhdxmjoFi0wDKkktcFDMp3T31KSaBjLjRbmlL6
Rbv+bZHN2e8En0B59sl4EEMEJqRk925eT/KTQc4Ex8WbzoefrIIqRi1Kbq0Z
tdzMhXssUfZXJjbdyi/Zswh6HWxjPI3HKjYag3AVewlDOWiEPW1TUmGf4/w+
DENcrZFqVRa82T3Oa+SJhhi+WUJotI6CCzeL7e/OfEyrNKjpefkNEKUoPHcy
YoY7mF6KlaOLFmd9616jYXGP6qc7ypw+tweQ2zd1nbMnbjrPuX6mK2epQfDi
U159/pa50yfvAAtWJ6Or6U4eqXHyAcEDqIvj2SP0vhoNF6VUeWrBcVq1Hqky
cyJ3a37dRH2T5RnOLCg9VWKkTk8KJFtXhAMVDtE/kzcLVX+aS5GWpTOj7/fT
LpTzOsk2TVfzgDUfdZcoDxkhloidbbpI6uNUbmePPOnHCwr5WdXWXhlEXuSg
TQyqSlR3JgrkHm49N1zecyDqPnMgBbZ07ooOSRtDy5gYvzt+aA6nfAB+/n5F
XVufCoBs5YiUsFleHcplLIFQymX38phllIG52cbwgmszRTQ/bz/aUJD+C6cp
GA/ta3MQl8AtaU6gzblAwXgjmZMU11KZ/Rcr7NYQWGrbAEcjSxQDboD9F2Ar
YJDqy5ZI+Hiwm3v2z3GRHpIGA0emCbfK8us6kgr7j/TzlwdM9dcr+dDpnr9t
46y/c4AusIFoJCdoyb0VKzEO9ba4xNapl65jIB+sCxYPCXCP2kTi9DmPvz57
Xoar1kO44K67enO7eQV7/D4clFn74UL1SLYJFK6Nj6N1JdQBhlgnDufj14V5
+MiIiltRUgg6ea1MsZhjDEphDIQnOUAqKhC0jWTVvcgK2o5+RfZAqfAF9XP7
ZISKvihcgvs9LdgfZKXyiLeaAtOwYnZ/rG/GKaq3aN58EhXcFHdV3a4bUNnj
hf5UVI4KJhuorthTCgutkzipnnb5VgItzZug/iG35UteCz4ioZDxAVpovYnF
X6LXIMM1SxweCmBOtcgUsna3TomQGjh4CWS+wlBCGmSBPBWCZwtXzcBtPDyj
7jSbg99/Mt4ZZ1kpUHn1+o8mGcKCsZzhQuMX2dwc1CzRjrRN61DekgBunMq/
dkFEjRpq6yiYQP6Gxve1STu2nGo4WsAXY2ToEQg8W0jAtlOdlgSipFZ/ycB3
Iks7HuNTqVnM5I+lqwAk6DMZxdBwYg8ZhMMdGv/hsKBLT6iMebdJ+oiiOE2H
af8A5svt21IZhrefy3JE6EYbwERqzfDVMx5Uw//Ku5HoPTFtNEzQkAh2olR0
XKMIWYYPuDqUA5xvTcm9RWNpRrK/zOiultHjoDzfjIuyNB6zsPRFTtoIKSvk
sHjmV5pKW++aSNRSeb4XE6XUjhxnbNQM47ZXdvkack5XRvNfT5UubSBbwtCr
maS29MK26hIaKUufcL5aEjmUpk4kDd99XSmIy6kfd01xmib9mK7OuKNL6cGu
bEJUXp9NUd81qSTBM2bU0NTU6S9gkfjG2h5+DJmYiw3py3YY/q4cEE59vQPR
q4Pk1K3ukTLcsSDHKOOUsr8bHwjcuJCyBQ9R4EjBl+5Nr/jcVFl4IlMJSph5
kqgwhGviRRyCXcz5btl9OvTEiKSUa3kR1M+h7KtF/q2j3PocxjjKgLPKBHQz
WJgu0QiHlB6N6Yu2Us4XPgy6PAooLg1CNcMOodNy5AG8wk4EL+9UpzlbkbJ7
ISXl762DKgViB1vPGXXaxpCvQBijDrJMiaOmV634KytP+LAVdcdzYrLYncb6
Nj5ByS1Nm+nXkkXoCHXlCiODt4+j/eyrs355tqtX/fBnR0Xa5N00i92Z4us4
+2ndMA6eSxFgzSrC1CtYds5oOQe1HZIYSv7NhLtmWd8lm3yX4ROYp0Hv/cgB
tdKxJdnbqTnNRGw7t1O+MS2t12sWcOcFnVFkDZk8c8ktz9nSgwVYaMAnd44a
tJUiGSRwO4Oog3yK0H8SnpFTNs02KYkjSbEuep925auOXEP2BQJjajuquqJR
w4+N8EGuH89MuLe6frq0yRIPZtQH77JDxW/yjAQNvWoJqb1hprT8SW1AZnea
PsHWDVlBE17PI3XiloFlmhBylAfqL4ubYVm00XHlfWihrsOjfPLGK78TdFp7
8ATnrpVQHjJ0gyHdVF+vGDLmPGACHerMkoI9yhz8B3vTc4+MLx1DTmNDCmY3
r7jbivadzDL9J/kQn0DgYgikUlJMEMNYHaAZPye3SbqRIGZezeHQVFIR3nq5
YjZp31TpIFbaqec+7/nBe9Od6ZjlG5DBOSACkCMtVI4jwdNyCkTiuf87E/2+
M3yLBDdNH8T4nJTAkJAjy7a/7wiqfR4wD+QSLAXP1baeT5vLwRSfgdy4DIIq
xS13WIHcqZWhUYrkA8e4PA/8cheR6TmF4xpSL7xd4E6kV9ZiN4JjB+AjDXzh
u6NE3KO+WSzXdlkzC4dtYV4/EdeIYlRn+H9KMECVfVoH9v6S2U4Gqj4pzBTm
2W5A2cmJ1Y43FN6jWSCl4MBFF0hVZxG9Rxv8D3QkwYO6UM5kqZqInzM5k9YK
XJhh406+qJgJdRd3g7TCYULUpM29WQt+c0gNFtQlxy1TC8ZWjOFq3VG5jKdd
KvebotxOWHyIeB5juJ68EI/SjX8YS+4xtawJchs9Crtv/SPouBqIWXzDDHqX
rpVvzmTIEt7YuGTkh/Uts4uj2tNCxyz5LbzJXN19h18cEedTWWuWQX52T3So
RG2Nzq2VUtvfWDpn/CTX11fWZOc7U9PYhUMKRGu1RSgIIsHs4iN+TnQCm+YP
5HAj1H2Ysf7eTaMncQUJK5wqPCmLVFiVDy7Gpu57qkv1zlTGg56W14OLy7OT
BvCvg3sV5F4lIW2V5baHV1CWF36Le6wo6DameQE1WnbJb530VVAVNBsXjJye
buFC/wp+0xzsaS4+Pl+OVNUwgJdhUjIksvQv6H5eR5a0iRK7ZZEKFR843d/i
Hgrx8WBrvfM4q2CqCcQiRn5OizPdkhb5g4b19+K1HBXtwGiqOXX7Mz6jy/7B
nXCowUwhx6e5H2EM4b7t0FCg34XO7XakRfqq/NbTJqCz5NCkbrlL/UjK/4H2
hO9ZvABkQJZK/CPBJqoMSp1w8MEx20pwMHjFYcMq95hAVxTncae8maCDHI/D
vnmeo9OOTggyxoI0ic0eoy21OVTRl3unytSYkxSixpQebvj66LT6j7/q0LgR
uk6LoMRWB1qooWY6Y7mPKeSKCLyf0PKG8cKXugS0n5hmy3MkSD5AbobYvywZ
LMMWXCYMU8wauOJMydF2gaUAyDaDaB9EISviak3Oqh+Qdy3wDt8RE7nRAwwi
DusDeipsazPaQC9A085uFdoerk4mZzi+SXbTfGxa7uOBbDX1f1jcti4BAo0B
CoLOMEtOJD4Hot4EYV3Cv4AG7UN9iaSrKe/XN71RmKupBhnQryud6uLSUQAL
lLJjXhikr7CXwP09MSLvsu6HhPo5WxRw/S3ehhZ9R8GO78KXWioI5qRkyb4T
BQPmStGMAERCGyXc/RFm82VsdomMWmVkvOXnlDR5dZEph+XcFO+NJoeiWuw3
w/lGxwFTI4pafBaLHNFU0Fqau1YvzHbtOxVaEGfOjmRaKkOsfiyEI2FCsiCh
te97sylnOykGHiYXsaSAG9UiAht40VSxBwCyJoYss/rskhUcDfNDicWMVJGO
SD6r+XOTGz07c79SYF5h9AUAEp5+YzhfPZ3jx00mtFfMBLLjwtlX4ciFNtO8
q7ItUWoQ9RTdSY4dnRmrx29tYQcZ4OVAGS7ovNpqIWEoafWYEcRzPBPYnKjJ
O+Q4Ap6L0PSrGrllDPfDRQpwTOI0ipedNptGdbQ4johD6oUk6dUiHk3sasyg
eAr8799u7PwhtBzplM4SQzGaS8NTZvXpKXtUGoQyix9XJdmvU7GkwAbDgUww
fHNWeX8r5aP6xMkUaB5KZ+VfXupYhe4WW2oJSwDC1ob21SnKrYfhEKaWPjTd
iV5i22nOFW+nI/Ka5CF0Zp399MXchjh249tyuqzXq9fDGDPjQ+303t3ZynlT
fWJhnO9NpFzOk9Kw1KpgwpjgDnMeNWogHD4VFF9E8328QJ9xI5NDCsDcAXFD
mVw3x47F6lKftKuPNTA6C7/HCqFxiga4I9CZRcZ+63y8Nl4FgUDrqKOXdLUx
FkqGvgbSx3+0qsTLKIAR1+Xxi/jejAwkXJfZyPwuL4GsHwx2/wUVGfxd6mIN
5shyje3XCjE8XRduYdDDWj9M1LItfVKWa6v8BxbKBQn+skD/5vhlbZ/C45mE
wnRX+ilDtRzvDLqmtcgC7hp9XVIpElHkVtoWxPedy/FLzh0MjIBw7DDEDIts
0+8Kl27u63cE72CHxU9UsU7jpYn2fUShGkoXBbeekIz2LRbiyr+M70sshx8N
he7r+OGcpt7Crgo6C2b3W0ALJb4JORQb03mnAiY5g4q39A7NYOntoKQkx+Dm
6YkhQFoFIAfB5rZ6H3DvauVDgmhLjAOm9r9SxcCkY8a//pZQycH2FPs+FS3o
fAsICHV7PPMopb6IJz+0r1r1wy4u9ENVpbyAzWq2KwMOiut8ykuRUjBbHoIF
4wENyvL//HDHaNJZ6Hak2ZQ75f6sclQPANawnsGAdpCf/b6FSU+w9WPtskT6
4Ez868Iyzyf9rHA8VfXr+pbT/ZTYhVTLfmArpD4mwKpxP6bInPRfcop/UpVQ
SRhCh+2Y0KhL2h/q2G82229X3tcUW+SyFvygDexoXi8KpYSFAapvkVprwWTE
f3aYMbL5CMEbyfGntZBcJUlnmg9+CQHdKnwX1IBuhOL6YVcsbkPn6Lbw9BoH
3RbhCO1bLV+zvW/UOMGckA3FbhfTPpqk5IsYTCqw/owqgDrqprTtzCP549o2
2q/UCoV5YnptpJAN6cnTB6GEgVfm/VZXunGr2JhGnUHO/snJjOiMs5gXxJbh
S80kkB0PTVm63bNR4DnvzTan2j3Wh585+YahZS8gbog/80nw8lQq0nNalskN
5t1k+UAlAYqlNWI0ofivPV+fbBdh09Z4pRslxmy9P8X+NICMjfMpMqiXraZF
K3nNAGS7DlXE4pC6D8F8ZI2lc5rfQsTZgAsTE5qSZ19LnzFoLUyomxBglf3q
WtXM3Zh3oUyWdX6M4rvI89qcJvY4JLNDVOIda8AASWBNGMiBsmCaQDIj0hJR
T0nLuK6hZpRAu2bjKxwKW7+MakF+xDr5drWiQ6TL75vyfhGCgKhc/cowUlrX
YLqY1jqiBheca2W/dj4+yGJk+mcuyXQ6b4kflDmTRMeWAmm1ncR03Jxd8hgN
WoorEwO2cQHMsSJvI57LMnLPDCRgOd/aNThqbJmIyasTMjyuDCJEivU8tv82
HcCGB/IdreoIybXu2cx5aAGbE83OdP6ZOdCkSvtxZasxYsbDEQS/Cw1B+Bcn
0EL2UdN5AK+HI/mcXI4zztrgOJVpUmmdeaaSwwFPxpuGP1ImYCuNx39eTftF
9FzkdGYnq6Y6l+zz6hic7hrqVaWft5Tjp/2YDfTapuekfHw2U4sC+/i7etSh
hRjlOhgNEMY8zGrVD0Hg39X1F2VBwPn3Y8avcNiZ9d1PqDro6fCGyyLpryF0
DP7XBbaAhzPiWQ5ly2CasgdTnVLtaHt7xCOodmkLXnE2amEWUM5FpQWgihwa
xltEpTEONub7tEuXsmDRGERNjeTzvnlxi2aIJbSMPcDfCjXaNYaid+TD3XKP
67Gq93Almyl5zvSB7HLmXQZ9Bx43Wa9KM4p453GMsqJQU0faS0aGGczPSx2m
gK/oZ7O9ZMnKQnuRxkalsoJB9O1SkZBaAfBx1JtDaTIjgNzAEbfRlMwqRcei
R/z14LDHUWoI3+EHOHxXwq2yKPOkrmpFeKi8t5xmgF1BNqTAGAxRLmMGNBik
9do/c5HxHJMUyefWc/BRnjkwEP4G7NRu7Tvegggvwmkma/6cg2ivrUxRkKfS
fpRA2P7c/icCVYXjNId+TA85PO2UNpeyK9PWSM+5Czy7ju7qPzfrg3VhWXkm
Aubn676LQd1qKEG35Y8+4GxuiK+EfkcBeeaK+toZgnRJF0vhtC5wlyPxqsh7
9b3OV5G0nFgy+SZUTdkjX+8JITIE9Bo0BrMBbO4wim94OkPiGXvhIWb+8SL7
BGzZaEMHPgnTj4aStUkdF2GfksWZcFGhtFjh/3KvcLBVtCM4S18M3ofH0m7l
5gxuYqJZkJn8N1k1caYB8hB0tH9UQ602RERKom+vOsI+K64cl0Z+bOBqEKhr
BiO0eazRH532TbRL1K8XD2fAmib2MCxd8dKbaJgg/eSNIk9iwvg9DXG/P5KS
TkYf4VSZmPOVe4KIjdVt0X6NAwOZLzpMDCXEgQZm++NJ4uFQKlwsZvPqwenA
AmnzpC2NghNM7gH7siUkUnRQibVo7dKF8VgkirbWPTgilvraLvud/jQrljL8
XSwmM0qX+D1kO2xl45aEGC3IKzaLhSFg7ZjBZU7xcCHGttCWh17ag+Ahtpiu
fO6v7cYSsY9wf7a37nb5fJB4AmGbb6fRPXLJQmFBzq36eXfoM8i5Pn1akz1d
ewaosVDeGGP2BzX/3swV1T6WLxlIPyeWR1cq2lF7Hlc60e7lWLhJSHpH+/A7
JUG8qXBMUHgyFcs9zDcXLNZxA4ZLsqXVypdJqiaom9ujlf+fkfsyKB0FND2j
lkT+3e+6giSXtLDO/NNLEJPO9NNl48BOIU4jJNNu8L/k7aSI6i+vor9YCKXP
Q0XRO2mz1fIWsboKHxBg3kHbRv9tqaCIce/SMqCgheod8FtkQhQtqKpK/gDb
r/NwKBTxzpUUG+4WGRaBlSj/3WyYrmoaFbn0xbixGPrP2f0zSAc5ZYfG3LYC
4j9OSRVLPxOlngQ00SvNtcG3I2LrNWMMpuvnswnV/WCSjkAa0LRUYy9GTZsJ
InCbwMjeuwjRWaZXEorFZITsVPMPwvphmaHBMjS4x43i3UcT0/DzT9TR4Ogd
5AZInLDJuT9AoJm8p0Ywj+9IFgfP0koL1M020Tp4+kVwVK3pJ7y0UjsTFygf
Mk3o724tERWooNYJXIcwIh5zv9IDcCT4GfENcQe30tEkSi+gzyAERv4C9hAz
acCx7RGZMMoh5HYxRDrQLCGQP2ML7xhA4Xom3yiXAqVJCjZolpJdyGv/mfqN
NWi2Mn+r9732wVEPJdvFYLLQfQkudzqiglChoMe2xO0aPq54dI82hu8BLWb/
IQNyA9G0/LjzfaIFQeDV1txvHqPgB+hOQObiTCxlqSYkG9lWwHN8QmQuxi62
o4YTGkXyOl6GyRa/wDrZnSQCcPCHu8TOnGlgOtCMEwEvqD6DUVro0MvwwwUc
l9ickJ5JW2cY5ZA614bX5FpIhRnhd9S+DgZAsR6cvWykglNAMu5NwDydYnDr
uF+wreTnH+esfnuSWEcRjqbSx5rfuk51uVyRrxuB63BD9xtnvySGphMVYY4H
apjhm7rX+9DplffD4wG7WCxnJEBrSortJCcYa5b/gDXoJzIim0eUA2m8EVBg
SuX3TsE0v6hTARqwcBdV0/hUfuZwHwENDbqAGLLsfVA65Na9AnbzAihG9KL3
QKqaT4f/5+ce0pKUY9/iJZOGcp471k1yOO6VJb9T7xVgGWS20CVcy0nzmNHM
OOPRR638bOvWQ/CTMb864mDB8XgRfW3dGk6KYC17HTdtL26T159xziNQuBeB
etSQ1uKFThx8SQuDwwIH6fQMdlQIrS43i+xRqwM5GNSGg2Q9gOrNwmq8Rq26
ehywxOuFgbAO2eowViR4OyuT7SdTu7ltZFf9TTsUeXLR9TIDZvmWRg9aNA8i
vcMWRa+6XQJ99770P5fQciMk6j6nr04oywi3Rk5dWyDvh9RqBlfuNbRYPb0/
F2/uNrVHiKQTjMOZCUIsVG6dNyFR7sz9LyK7RZB0Khlq5yzPj7hUVhj/ILMp
VFE/cuOqIg7XUF59a8Ua+zw9CTK4o9RDr0GlY1n0ny1hfsEYtB+xAlzPJ/cV
xJjTVruhenh5YKTnVs1PfHGhTJkCgTkl1OMeNM91kGNGMqq6H+QrDRadiJBB
TYQw2OWfwi5pRnqo2ZB8BByUm36+RJQipExsbjnxHm3Ul+mIvkbhhJ/0FgOe
jY70y2ergWfu0jPZef2+R7J/J3EoTpTM6eiVNT/kUxEOhsO21KRicp7nGbIu
XYN/0eUkjXX4dDHOwIKDZXLJGUJuyzfE0rG766ydn6zR58Qm/PFcHiMgI9xe
l+YHYU5xgle4Z3jzujpO2FIqvCOhILtpjwKhyvUNfbaNbFqvJ3CBYXBBhnSD
YLZBXUgBBS6+VBCDumyVXqlXPfButnLZ4il5YX++u4UCE0NbxmdDn4q1TDOT
fNv4fEMxasUvirTQaeIwt7VzqtRX91tizhWSyQPRnqGpWCrhuRC/cnovqdL8
eREtDrHwcMX6ns7bbXV/bhg0p2UTiEpIrHsqnKZcBp9NJ8KJpSnfhGB5M2G1
uA6NBpxZBaIpYZuE+oQSbVt1wfOaIEj5gArqxh4VOPza3REWGyNOkL8sGtu4
cXJUjP08H3/MxsdapUnKUTSUCgRsaUYMNAUPeQfsGmcvPbAkYvzZpFIoruI6
d7EuE1X+KZJwPeGcub0+5r5g0wWLMJEfxBN3OMBP0wK7KRdLIZay7z5Fms1E
gYTQJgn73pLbBc7G+K9RsdSSdyKcTrS8q6LvSmHa92qPvoMypusEWSsUsH8f
83MM+yeoQr6TORwIQWJLPCI1GrL+qfOI1YQtRmd1haXcgKG08J92MzY2LzfG
Gq8gPCnQmjU4IsE+zc6AmJY4vRJEWxPOuoNNxDdgKCZ842AzSQKX87LfxW/c
1NraqZeFjeggZIvP3TnJco97rC9NbWBM9l+8zZtNXSuCTJM54m21VznyE3Gt
KEKxgbtI5cS7lR2iT40FS/n0+uCe4YXOIZOI1io1HNuHlqmg3T6g7B3covET
4BAps92KRA4sV0n6shz6MPmVRnfs1rtjzAbn4NGv9S4MikYlq6/naOh6fdMu
JaXLN2ARGDDa/zSRb5/lMX/L4039x50gPI5+Vh75KNSkyK521xdUXagK4rAK
HEXRR6o+5vmtO1RPCCXCEHZgA8KIMYdq3Q9lxdpjZ/lP0brb7WUl+qJscho6
WPIIdkHXZ+XD6L/dpqDmNhwy1fgaOYeir+wmxEEvkK04dk9j5A7dPRSKY+9H
J2dH5Lgt11r2Gl6kndy1bFNfciqiDtdHOylSHCK6B4RhRF6pPDza72npTJCr
tQ6UjYCa9WQr1ER4g4bw2X08bUkJx1zysLjV3Jb2aqYGY7/JTDci06dlzqPT
6ACdWoGeLQkViriB4nelNS8adaWqDlpM1PlKKAaA59JHJyEjoGWUcBcip0hD
pM9dDPamos9RBqr7n6uNvpgBFa2JyRo+sm9EFGw9LdsZqZuQVogxH3cugBbH
u6rKQpDm49SlzdXixTKA3bQbK4rBgh69NhL9yExOxyjM8SG7b142TYC+BUSb
bzZiCEM6ds8Q0m8dYwPH2KTXDofyG+EBt7ry1htY9VM2h8gtqbcRlVX/7fUU
hmBdmsbqzlzvSaFYl8FBiPhbnCJz2a3OJ16dAJKvbEmwn0Mmx0clAKVvqdQb
5pDoc0NS63KbH9frz29Ok6GjEBhh8LR+CQgM7XFL/HPM5XgDRBd0cwn/yK4q
FYieO6meXVjUTCtsKesf2Uw1/tuUBQSvdE1XKOdfKpswKURcxmANqySOWHHK
qY6puUkbyufq8q0/Sgpg9Ah39pEzskEQFP4aQyVauX/rOW7ZaMCaaF7H0V/B
FxZ6z06yUblQk/RFi+iT5yIvDxHL+qFSX/Ju/gq7kgTzMK1+PBiVMg7Z3aos
CnAa2HZqgjWpgxtk9eH8VpciAblfrl1GuIiD7LsvAz4A0ipGhBTKU0oCT99g
l6j37/QIGY1xkrKl3X/7qxAnSjuqHIXDn2OdegbNGCJnixIBqKsIQvdVdsbX
pyKvSrxWmNTHRHUXoaOfoQZhmJriMWiTY87Hy3W8yQwgxuuEvl/uOQt8cNOW
36TMO0BvVqHHb8XXhIWZPT1OmitY3J1Tq1a8sfcyhvf8Pmjm/oZoYgpFQbDu
gfowOtA50KoeZgP+aHJfr16ABvROACjLswtzAg8mNw4YO2W0lRJrPF16ofHB
5hIcLbVzniCgLWxZX2U2uQO6yuKkczXtoTup/KzlMNZCky5et/RsZeS5VSfy
8pgM1r3knOrWsJcbSeOVur+jCPt5+6JAQvLI1xbyABH8H7x1ZVqjh6oH5NST
bhy0mbxItdYEXnYPgnwnuqWcuAOacMYxsPbfLjv8qF13wSvySvf63vJ3GiyP
cOKUzdm9/lWWDude8CDxJwoQfanrt4JowTrGb6z9JzXzEMUokbjNA6gfIwiv
LnOMqliaaZPw2kttfuyTNhMNZ28k8A8oDeqDN7fNjBwubh/fHS3bFmxu2NVt
tqjwE5PeK4q1on/WxfHYcS83ntA/UBVwUvkI8Gmu6M8tv76PpdhCf1mi9rlj
EfFbaYeW2DanDJxPpdENGypPx1UkX4ascNQu8M/u0/8gBHLzWbrYX9kC7ysM
ODXwt3tDZne/v6bnV3Aq4KaDH6wILDuOsYCDxj3hAbbOFbgk7Z6B+Ww21j8n
8RNJPKXC54P/ZEML1g6ZpDweNILE7z1VH9aCgD7JJwljjpN9g4DgWkeOiPaA
3zHTgQFp7cTcs25gYkKXWyc0q3iZ6Xk50OpqAZXVZ1Kqo6rD7jOvMohQFFeZ
HjgQg+yg61A4XbXeojyOY6hPeLpK+XWbHY6UVaTA5w8RFXp7GZgdA0zvN2wn
ZvZgbr5aUN5qe/t4ShVmrrVf1QbxnsCxXz/njqwe+H+T+JWoojxi+8fY0+qT
i9k0DHYdr+C0/jcJu+fX2WcDtHtVpGXEy2rjJR0sR8vcRuscSjGFWuWQb5nW
pMCIV2d3RaKOidUmSIob175y+OOSA2GEF4wELLkjz4tn06JZRkxDc50bw8gM
IOezG37YU4LtFySTisiTSInXkpcfykgT47fD5op81sVIV8yN4+F9BkmV7ipI
PYi3L5Vn6j8wk5crvDG+CMNHN25Ya2DycYCVE7VlhnKE1msfsNvTEoolA/hy
7qLappu1dDf0rBsSojgPyX5a1zsWnhsFwIhIYz+D3M5JWuSbm/uRkPahUDOI
m7T77zeUMirySrdEBi6q+s+C9Cv5tnnSSQAljuJcRK6k5v4Br+zZdyLx2yfD
PkDUR5N5NqFkncz6+Kp0YbdwJq6N/BRnOUfJ7/OIEBBmIOZF9eoi1/cl9Qbi
ULWRLG2jGJ/fcLM8FEeJJUTHUbBBVJ6xa/koKSAT+LuoUlGSBF4DH//ltmRo
vXYkYLMedgqpoYSKs2bm/Az5EwRPXNdwNdRwpYD8c0/SXPPdCXkRWxawXTfb
tOYL4ewjv7bYtyciN13vZ3NkYNoFO9WX9UIwqU0TrYeCcSqRDTi2los3qHyy
TW4K/2nYZYeEEam9vJTNbpsvHzRjVuJTgdQPqaB+PjAFWcIOw7A1s6apItOB
UkWt2YAalO8fdSxCHmViirHLtnK/VuN37Jyt8XhQHEhsb0FU/DntEmnZMTdQ
OPgivlROebtqZQgel+opQeUgtdaQTHZEpSX9TUSJqSY5/LHvO2DnrnGWNw6I
uJS+3tSeSx2Pvqq8IVtKQRnoTWuNLo6/MfKRoyHimr1nF29IzmfihrvbHMgs
rOIigKozTaLLqvix9dqQIUTI0k0pBon69EMDCIx+yFnM1pHzpdPwLS8mn2oA
Cs7mkPftOCrfvzEPNdHh7tCMpJHQWhVZvNM7rUrUQl9fwWs/IMLkXeeT4gXT
L+8lcYKWdJL5FBfAevQSODoPOtyVKKy8kTl7k50FCY9y+jKtv6dy8QrszLuW
XH0A6k8DHRtd+8NzDx/fYrJkuQ6GAPoKxrpiWJbq4woik/wNSr3MG6qfzPX6
44W09VSUQht/DJ5Rtj43ePt6yWazkDpbCQyoPas8vq74Lx38tnPD0F4h6nbe
pVXIO/2A95Vw8eM+reSyCI1jHnVwzNe4had1L0MLnzCYTGdQSl6GL2ODWvr8
dfF9SM8FCkh860hmVEAIAx/gatWqf7imdmH3RpbV2fRqpO+ih2AD7EFbl300
KO/dgCwWWFGydFo0LmMxuhdkmMe3N2Mc/X2I4ITzhRRN0FiUaZKiFN/A5e/6
nlJYaCzzVR0No9L9izMUxJfxaO71zMMNKhwNCamqzw3lhNqv1W/Aat0aTlZV
UgvTjCuaZnDUXH/bjuiSALQDN6FvCtZaKe8SRtN0VvYjmVGXJRiPwa+KKhpz
778LIzuo/NO6vMiMJJmFCIjDIW8gXB6e2SkJ0arMcbRb+FJsKnLtHAWdTzrk
qc/SBpNW4g6l7J94KIFBFSM0xoRfgc2En8gF05NNSJCZDKz8CEaQU8z+aA++
RYGjn1Hi25OHld8eoYRdOS52fWi38TI/2PxHMnkaaB24BeHf7LssVo68gDSX
12SjxmMYQYe2YFNWmqxhJqbuH5TzZDdbgfv83w6qLfCSOrjyXpCwwkq7Jrdw
pgMtygafvP58Ybo4/x2vyeN/RXGKC1Tw4Zq6IviKrIX3dns8jEtnkzb1C+25
YmbW/+Uv2iUjFpgc5apUSzWknai7DA4n01b7BS8LzYw8Nucn5SeHU0ql7rF9
5125A15IfnxgCcK89e5EAZGbSVvn8JfJbSHTgofRqgpeuAo1ZDOyPjp2L55j
IqBonxgnlr1M9bM+y2MP2lpCYxFpoJj9oksORsAGeQVfa4oVigdXmZ/cpySD
JfT38rtk1RnI+JEKQvEd3V3R7MMZ0vfZAFcbNg8WwugnH+PjOg+uypqjYdRi
Gm/1AfWB8fDVTYUFmk1oSSEh6qfSz8HwxIbPpyngCcFEAoqfDrn4PzoIQMsW
nJJFijqiMV3ukYzQFBnhKLJYwfZbEPLLk9gv8V9f9FLz8o58bEa7OD73iuhe
ldmnHC7xg3UWp3aWoy+7lVuWOdoE9Akxsdn1u6Yhsp04WZAGkB8OQMN+yeyC
WgEBMm2q77T4OLDIEMFEEKKsQDPQctzgcuffJbMD4bcWBrj9+iRC7rFnpdwS
oxXBssFhyYZxYg9X6SLAFeA35HhgODevwDZ22PVfJAnZp9qIxYaYp9rTVzHL
DaYeGgszGHaWOvJasHR7E6/mq3RrFbo8jEivxXY2dVqZ4YfiYn/PkadtFw1M
FtnPCRw1PP5rmqGj0B+mXGFy+f5iJLEbzvPAGUGy48XZ4DHiLD8eimFgPtZ1
9iCRt5U9aCY6QQ7ElKQ9jOe825Go41Iy6rG2nfTUweCp3kWsTPj/7kAKsCgq
4lOfrxykoiKKdNrVY0qZcm+Vb3zdIu/gIEQb8fyfDbragh0ZHEPoFOasR3Y6
nnOMotRciWzkRxstsJrTd6YHxXHP5VTEkHbG8e29ejPMkPVlvxRWSP/rZnKV
tCe12O874TIeKt614mweOT0vpJfcIJYOS+HfoFiUt3GltiC6la0pYm8pT68f
llnmMvzsHI4IEnj2kD+0n26/p9aqEWbKoHc6kdjlFElqi3/B5brcr8ahBBeK
4l8tG6lWMeZvQPV2QL75bfPecTHnFkm8sygpyggoOYonnOjNhxovIFsk9D+E
kAox9vKGA9vDI94LrqWY6/nZrdiDojIAY+csTIri/ohWmjqzvEIIuNvwNmWz
GAFAhrna72Iy6J90EaoeIvZu4ZOLcJhLYJVP2E9X7m56P/u2nUC8z8ODlP72
z36spJ3tEeM1AlWma8Xt6Nw9rsWe1U66oVxxw0OAHWfFlQ88UJO2OWu78d1F
SsF6PoBKbTAt+p9RQHlsZXfJaRC4v48pY2WxzGJRxKMAZHT5Tp6p9i7+TuRC
JDmqQFkdFYA4pDV6pn2bd757G60eBruMFkcOrcgcEnzo/KJwC5ShfC6qaN53
T6+et+vO5YTIPtN+XlVvjq82jqe/zfTWNnpd8Va2X06qYEVJgx8aL5YORQ0k
pWR24FIF5ZfDp+G5wyFk1gzkbnIhRilXj+tTPoHO6jRuZsGbeTPbXlPXqcux
Ee0Hku6n4jcCIamiPnAwjIcPjvWATykrazJ/baNk6J05erwltZsYzzFXmOnx
ua1bHzEk/Wqxv6F0/2RNdwphFS23j1G81bGWvJDZsBD5i7z9g4NU+gZNftVM
ZIoiEeArMJ+Z98AWh8ohOZIDsio4jLse5MR7vGONqYRwX8g3nAt1lOlzihh3
wC+yrJ8i+p7Lj+7SuiHgTRiE87SiaJwF7psaegjXFtrmHpwXJzQEYoLAxjF6
8fOfihXsfbn9tPeeoVxfVgG4J+07+tzryuk5VG+9adjhj3jEVrQU1IWPGUaq
FObaBkyRvbJZj7uuwnbQ46PVdKiHvl/7ZKUNlPs0jvUX/RtIDNEL5QmjdR3A
9YBk+FNODzlHX38i9sG9WdRCss5DEt5O3CH8+8R6hCcJtco8RQKeG9s+1EFc
iY6p4uPifYBYeXfKoCQQDSEWvlgL4w4ebTDCJmrSObD+b7XuWXf2hUU8F+mj
hXmiVDZvibjHiBxhmJarXlymGDIwMs8zt4W4uwZf7MQSkxHtU9y2cJdGZLEf
qsXYdGTgeHn9vF94eRSy45F+kdMLWc/JNxMTSealCYbgfXQNgnDoALgZUcAj
KC0iKwcSJfmx7+CYFFKGWAD7Ti7e+eGO7PaFWZOrGLfu1Mnu2H8R2r4icgTC
q1IsdCboenFkyhqsK8wC1CbD1C3iZcvx2FwrGLihVRdVf9vEK/QTCM87jmCV
SYjWHSoYCX2BeOU1cAmmyh+S1dvlSOYpDTRhfCibmZfPyLLHi3qVhovD/Bbc
b1JTkqqz+vC+33fjBLjNrOJ2sDDYZLZnxq/g5nqWOHOTIhsj0eZhbmP1Fi7t
Iw5EuuFc0NPTQ4WVcjb4Um8cmELwhrFV/ECpSv9pORKv9T/+MbIRP12Dhmhe
azcp8ABmmEpZ1DrKe+PosLyNlgy+YZTwbcbntHdI7GOp6uKiPLpaEYPJ3fPT
9wet+8Npm5pbqhSwyRMmwwwsfEvwjGSXqLaGuvir529Ai3OShPleb3OiPESX
WpbTFfz6TMecnZ41W/fBRnu8wxCDaJqlJsyONcIiwu1CTxcGyVb5RJplN60B
fyHBTQGzAU9O8za1zRJlPYTI37NukmG4xg1xATlg8V7tUWyVNphjnT9xgvgv
jR7/daW/NvIoIiO9ewkcVTsKhc3xAaSt2nYguYqgQ33HV5C8psdBJrFjoOHE
NJ7E5Z0lofMpGFYOcnHjYd3/8BiFwWeDo2amtbD9gH90JeCddqq+vx0wz6sN
PtURYmKgRG4JQGh9/BxB36eQifNuFGZ1Hn3rwuL5fFdOhi2ttASzedXKyTbM
HweQSZwLCOJ0p+JfoDtrwhjcSBLTHxK6UhhzIV/tFmSe5HXS3exngqZTPiB1
lFprGcYIbyD+Z0ENwiUeCkxUgiUlUhgn+5o5qJub305aCFgdjLlCgxrUWmep
AeL7PMLV2HjonIlO7NdHRDSkJt5IYUuCRESDbjmWO5V3zz2slvu5WRn9kOT2
6nWgOT4kzTbAU5JA4FhDpd9DvNKVLXFPs+/fZ/ijFqXinjWh81w7c7RNRr1J
BssoQoKM++IEBAyJpGIQDB25jgdohFZ139mnBtlB+3cGCXQqQL8RcPcoGkSf
47KCFXLwWuHBtUAG9/BURs52i1fh8RgLKON2kezs/0TqziVHyNZgPTB04CVz
F9dq03G6MBAEP1x5trfbRHiFVbwDopyEfDkDpTLTYQc53H+AQT1VaR53lT2c
9T8NwS7ffZug9uKt8fi0ugqTtxY7dk8fc4eMfIBM5HpsyoVSLCPLWhLdMTne
r2FepV6m/DopYVRgBUMf8VMD+jvUF+fgVXJ+WRbN5iJxQi0cr+cVYbIV7gMw
5m3NytDhd/VSVqrvBZAGCDwSvjn2ch5RZMUA6Ick55cfVXSyEwo+MmrNjENm
FNJG7CYk2L3ZpQukCJQXQcozJbCSCL3ixFCUfGohBUx5OyxgqiYg57IOoKRY
SKxsTPZiRf5+g8uAMUmi0e+W4KZv8xPmdikzX+DfXImS7q5O41UyB9jAUnrV
wg9JZBzOTgcgchJcZR9DOsH22gVGOTI255nRlTIhxAUfvOyJ9nhdZ0JU7q1I
ZV/jBXRjsFPquELJEADOBFx5XQZABQJy0v5mrBKtanYfj6c3u4kLq/llBuY0
CYB3KSzjIrtrMlLcmULk1bzQOflRilk1MLgIqKrftdNiAHpPM4lNJNBWxyW+
78Ay78eEjlIGFVbMIL+5xomjLdlWao+3FXcjrMx/Me85pNp6p9VXlunNXU+a
lvcszVt7TMqTE5q6HzkhxKx57/eMlIpGl56Ky+3Fk/Nfa2kmWc9jVWBGDCBm
K+ibtlziLmvKW8MH9kqV28WFb2ftu3kQMXF7udZyRzNb7x5SXjuh7p73V0Nn
hX+boX6yBGkYw5KvMFqG+yT1elOZJkssQzZBl5WIE4JQaXBF8EfK+zGgifF5
a2yjC05ZcRdrK5Yyq2o1AVJ18ZiCesTi3k4zHOeuTSpRVhQJhaNklhzqhrnR
OFjzsOiLzJTrAdimiBzZTpe8VeTXoKhd1iltHb1GUBov8ul5rU4jV/AH0akA
LYRdIHovueAvmTxsSyxqnx/JtJMoQDUobp9ul/Ta2peJshQxxRqqZFcYgdFK
H9bqkrEY7CawC6JembYi4ffe9dX1YneRkK7ygACA5yeizY6UHW36M6lEhUaS
X2W36zJif3LcQh4GUS1yNdp4J1DRqBQ2TFe51h4SApC3iPU/n+X681XDPsom
gmMGNfLJUZuByuAlrgX8xOsC3881XJXGHLVBIFquflYzP1kFZhGjKZTKjwF/
UYMcJuZkYV+rFCL1aGab+lfiPXKue9QIdjQDKcGn8a7nS2ABnugjoF/j2kGZ
XSUkaOxzOqWQrSQnztvB7JzkAG/Y+cpw4SPJPhgbra5F+Oc1nNZgpgQ0V8YZ
Jr/KVQXssm0UqAO1U/HEdZZC6ts4OmbH/Fm00puWTh+K85JPXfk0bFYR9KvZ
vg80zU2TsmvV62vl0APk1EzDfLeJL3Quqm5HGKoUFCR+1AbJ2KSj0MtMOUWs
WDtAcJJgDgI+mlHHaOt5C+vx6Vp8/DwpjTGy0U1jOHHo34KYcTT75YhTpei4
4PsNgZn/1IbPctEu8g9C8WJGTAbtY1ubt5S+/8NAERubUXXGZS/wf3Zj5pOT
NdX9G8Ud/WwiJF++rXkKOEoZH3E33XyBaBNaCss7Bazu2mvPZ+JjnVRLN6AP
RKT6lkuApMSWY2hFey/ehDJpiwYfmElQOa55REnu1d5d8QFMumyCPPocmwzV
QlHmw+XRl+uSD5BAVsfhgQ7O0BkpYWcX9As0sXKrGcmtpNra50yuE06QZHP9
5s9UQmNRnFzDDbjLIu2kud42nWRUS/iRr9UvSdmPeHhlIITtq2IMLBOnXh8Z
y+GG9uIZvpiVD0s3uJE0PKKnbp545MNB/SnhrLdBd21+wykKra1eIinCqNsy
E+o30gmChXpKnIxLt6KHgTzZLkzRNjX2l54Wka1WIZXvjhdD7BybOP1yE06h
UAtfPhh3Uz6wztfg7vqs70epz9G77HsHaVPfDMu7mBvaqNmDH4ftFI8hzJY5
dx8vhGVU2ghg4viAjuuB/zKLgcjpCnLxSPcb+bFcWm/VziW9PUlja7n+u+Au
HncgW9YgFLBuynR4qHjlhFeVsxTGIShjWOrsqabXrktNegWp6LhRBjetNAtw
HaXufOXthDKR86AWfs1QbSMQsq5IC+XYE3OneVP+mli4mntX2nVANdjTNFEr
WPsv5IDrvkAFW1420fdGvjw81Bu6WMeInp0nLZhnrxKtwkk0uTe6uH0rRh58
dkF5IVO+4AYJMA0GDIHl/d8VDcAADxDNF+86eaPBIlaEnQkgb1Ydb++KkD2i
2uyMq1+HyK53ykJbVrmKQJYBgzCfCo26nyn3E0d1aa0AC0F4r5cBmyYDGs3Q
HI/ePSx9eX1lLTotXphAdazxC1IW9/N8+TPYWD4lRSF/NvRMCSZe+bHLbTTs
8oCGUYZvyobqVk80VyL2yDZQicsLu1yvAwqyhvFDCR+nIx8h/W/7sAhmb3wU
jjpgZoGiYywO5+3W9rcX/2gOEGX7NdE/l7DSX+YFPy34LWY0KX6uqgwU6aM9
b/678YOKD3BxtP1/TQWms9H0HnpjCvMMLhUTsz5+ZA/3V3cwhRN4ggtEzIaR
qK92qEwnwXN2qiSCMoXjiqEwC0bX2CwT6A5O2bhK8wxMXwBPlCzdyLqfYodt
GOcesFPQMAJp4gzF1wQ0mhYGnXCNMHBla6rW9+VW5ondzlvNmD3rVsbmCj6O
l6hQ+mikMxp4d6ytPGWkefUWhrulwBeNhppT8zNKbAA5FOFC93y5en004U95
TUcCMZRax2lsc7+2sMOSICAHC4Y6to+njuE/XVaNJwQPeSOh2lRHEQ1fwWd/
sy1GG73o48Kb0YUrrywDjXyE8h6rLWV4+stjiG72KNdxQeOH2Dy/vU8t62AB
MdQ4NHesT0aI6FFPrglPNKuTsk/ha4X/8Uiy1ONTDt7Y4Jvd5h4QEihb/u9V
FJOkSlJnFyRabKjR0nrgj+eSndohbSLNE3B9K2BFLA7RmJQIXnTm2k5szGJl
/Mf7sxveECyjscg8j7m/MV6qn27T1Pr/tcC/bGRONvqTDNi8l6LWmulBbyP5
lp8QWIuHPnpmCswV03PUxCnggekbbD6fcEYURdyJwhXKQ81DPgdnKPwCRQ1s
WaBe13Wg9cn3KXSJBrqszOHaWjy7a7dC2rNFc9XLrc9nFNhoRu4ME/981DH1
N7x9hlJhfkF11PDEpYcDAqgb56sVxQs8g9gd1EzWEyRJq60y0q8aML6rZh7F
MlyaRTfFJHKM96ic0W0mtZoCnicIvty0IOuaQPwXM4SMqx2Fk/a0yOmYXlif
oK0V3cMW36EHBEtC27daXwIaxuN7CtzpKhlSGBBrG/6EJUOGnc9cpB3EvIU3
8OFPYfTYSkIuBuoSRM7Ve+8HnHJRDNC2TBPpiu9zu7URBtz9lwvx/VPoF9FY
uhNLCAgm05Qx4g9PXyFzEH3J/gWkr+l4x4XbfzpRQuDE+sIkHDJrxKtA9AHF
0k2MDs3lBM8dh/tDNiMcN3yT2oULPu2F7nJ2eclCZpLPvQwa2NyH/FI5clsR
mvlUxq+KT8ARQojotlgaic0jvTIq0TiCvWtOIvk1RsNxZ50rv12Syt0OJuPO
zWNLCMy9YuBMpX7VEmcUekDJEzJmmoZP2bmtwvYJcZoZMLvckHgEDuA5B4Kh
GqoRarbo2/eNS1OYz1IbGFVIsf+j/jF3WnohVCIfFqAmvKc+1C1Y0am9vJ5Q
BM3mTbIsqTUvYcopAT/PhvRKTJiSJKQsX24QfQL6fb9nfH/PXHQJc1KjgZyl
wrhau8clBGdtmull4IvOQfHOulYX9YQVFIwidz83i+6LAnWIf+YDYIt3xHBL
34Pknggnu/EGgT60ZV6hpuOJzkO+WrDmAhru9YU4lj6iL9ca6wOQA1PngBxe
QFfUT90B8vdgeITrQY03kw/wHDZauasMZMQ702rXeW7u6zlTAdN56zthGHxo
oRSKIshkBmXzRYaN8aJFZbBjlikvDDblFMoGPRoaXYHH6iw8FDviRQOtzqLw
uUdQIvwMsHZfG4e7rdnGxAUMxRUHBFgnrJN11ZryApELIxex+2+5xXFwy63K
/pDqTqxKIyhLaNTOmg1Ma6TJRvRyq89WzkkF2OKxQfaxRVd6IJwcOmRoKv/h
zza2mnGqoinc/vEnoF26HDHMWDOuktokleApJJ7GVej+4REokxXxBKMSqecK
3BcbQQ1SlcSI9JpPFLuYypbB/R3+GibeiAEJIobM2H6LE1v/gvvanXB4RtyQ
uyxFjbnIlDJQliHtAl0uT/ZXNPapjNUWM3ruTk5kivjkoT9qaQ9xWpQb7xZA
QqPNfyCWN299QA4j/CyS0tkUEN26RRi48ihh0MvidxViBy6oLlPPD8jKsMfi
RwxAyYShHlu9MSmUoba6T2AIa4I9Gn9dMEaG/IdVsMbO6YG3MmtPkMvndUbb
hT6IdqMjOUaosQEnR7gZybOOOh2IcRMdlRhOeyFweyu3THSmnpkGxHWCaut0
d4kriucyIgdBwFRtJ0t/wWBTrHKe7U4cFKRUswh+V0u23FQbLHj/19K/LWWD
YSk6RZCtakD2ww1AsgwI+8ATET1c8ZDDQdWonejdoPkd3lPB8RtAdoE1fQ+N
n4URDq8dGTBR/TscBKTBrCRNnGBzg15GVKZG/59Sqo6omgG3E5tTHyoghv69
qIufqJJax0nGa0vuIViEif6E9XPdlM7d5L4nefw8HBFBsWazd1o5VchfC4LZ
yOzWQp3rhNSXKhY0x6QIE6rgHa8l+O2m1Ef2iVWSeE3LrJrpqFbKHrN2b445
dlbj6kc2evNNeaGmGT0LsYwPqqJr53u7Jxk1XBSylZRfh4nffTx8dGFiUV3u
HOowlWaaq4+OQMWrJNZe1oPQzCFZc2J1zlXK4QqFysoIGrCz/7YgvOBkgbVf
mURYPUtsjfKZFyO7w3WOsmuhH+NTkGKIGNyvMVLKiwIaP9/oUd1in+K7VYeE
FHBQxIVeTzYhICR4KMf6lcGljNS/opjzAGhMzzuVGgpGc6qFMVC75JM9QBDr
GC15AYHhertCXs5ykDgrUYStczcdW+SkDxBEdQJSyL1cBf/TdfhUYMyDGeUd
smtYW1TZhvrg4WykjpJ3DsWkY5eQ9ZgfU9iwhXvrOQodL/HGar50uWZua/ho
30ylCpQhvYY13jMS2XIPeRslt2Hm9+BGzAY03sZMVi/Uf0OP/G/N0VYjVSIM
tOQXORUYdCvoydfEyD9RZvU+bY/PMM4q+yJn7aJ2B+KyR/iCYF7i/9aQ7Beh
JDjMUoPkWl/90IpFArqBT2yrNXtDA/81vrhoaI1SBejUKHeJlcuir9s0ZcVX
TH4eHyxheFEf5xUldmlZJ3ayv13Q1x/RjpbZjW8bYOFrnFlWeZZvpiw8Lr2/
P/moQzzxVCj5LuZATHYyg0a78lK6JyYJdK1E+4D3smrtN+kqOe4SJg0qXEbc
h1hVCJEMzVzYxcjHexQZlNLvEbp2DMTPJMzQxMHBsU7k2XivKfZW0xu4uBaI
ycOtj7vlPC3H27BBHI8FQoZT9+7bd7f/SqTKPRZBBkt87F9+ITBlKTmqZyeG
QQFRwykNXCoQc8Z+3TgX62A/8rLGQonOMBYKmxQXsGaq8BnznCASdjwtVcUt
V0qVgqo1WlgkoPbiTLftpC0C2Lq6FqPsfWT4EMh05RVH8bmiaV+FVb7+UgVS
4LVvUktkUsn8RRv/JpODH+7a9VCMdJzxy+dnSgYiTcyUFivp/YffTbMU5G5Z
y5EJlOaXfD8y5zWAS18TkTpK+i6jA47QEaIsoJCyvq3v6cX0DZuEnCi29pos
L5GcknktJbL64iomoeR/kJLuwLXrl1awIhilHLRAOfca03Fh20OjB4BWlbj6
UKa1WHIrvtUiIZrV9u7dHXVYGS3prCs4vyIK4CfRBh9E9yrYA1rqoUjyJ/jz
/Y5AAMg2VjQ3+V/zi5/T3ziM9rNe7+q+EVSd6hunHHJ2Nk3jqHkZ4D1lrV9F
VuwZWKdcwC18iizTjFiRYwT0r4Agf8haIQFJINH9fv2+RViQ7H2msWbuF14n
/aH/ixE9sd2Jbc4o9mQ3C8jqQppzy0wmvCp1YXEfVCX2jH5PUYTRZhB3bCtl
kqgziZz8jJDN51cbjBtCFnd8xqJ3K/aM+ULupcswBPSSowqCosAIufAEUzFx
6O+aaSidGdxY3xcH2FSpwJTvCf+qMh79wsmkNPPPs/N6IwyhUo+SjIROy7Mm
OL0HcJMt2nPSuLiIz3nCGAEqB0PVsvF3n07lBGRNjua21ZRH/7xEpDrhomPa
k6o7aIrrdAB1/dVJ/qzCctWR/O2e0KHo0i7Q7ei+olVjjEilghS5rjaI4DBP
CuwgQe/aLoYTXs8BqQoU8tLoH5U48qFhWUgOwHtsxl7LhqZwHr6SAxWON2F/
tskayyTM4VkscZrvR1uZQPRxAqL1+UnQvVNSDHL2pc4pc6yZijAas7dTBFS5
H0YmtJkDg1ze0L7oM9ZSCUNBrGfFaTe9KUsEaAmnpseLEX36YyLlxCmYMS5R
A20ibLDnUwbmis79zzvf6qQKqaY3scwrtpzb+7kCt9UlL5RgiNFsmNJdX1eg
nUFuTQfSyUY4Sf4YBHe7zW7P7Jx5J7TXMTw9AltMDEIbug8oZr1Kklp4RqCE
RkaiXxV2SXAQfZ/qpkcSayaxHrJ0I5bEBlOrCkCYlM5beNfxbWoOnzKiu8Wo
AXOM4nN57vpYLGJHC7WgB6vKcksmpTuC9qiTqMC1p3ameMP6C21wNjt7Pt5h
zSFHfcQ5gROVXsd9K3scpiIZ31mr6odTZpywUH6rufC4Zb1uUQlzJF3n2GP3
oPVPZCCuJoaLY0k2TPHsPc9QoV0mB6UTYGHX2Wt8GK5aDnu9ELWVyVHjrkQS
zvRPEosRXyOuyxGd2uMCDdV+8gtR8MsQhaqrbOVn0HHDp73LjACyBqpjOkWJ
0KOPZ6StCBe88baYuMoHB/e30FxHniAeyg8viKs9PfZ1umjLELx+qFIRkyuZ
vwUid0z1R5wsI+FcSrcdQhIUmxoWTwuFAdeNapIYa9FrlkcpZLVy5dZAtnNM
GH4zaXc4qATRmf6Q7nhs7mpXfxvhoNCxvGlo2Xzz8DdJ1nXmL/DSnbe6A/F/
Np7uttokHS8lEtdMzvpbeMwgKQsmtnEIi7ljg1aRKd25FmCZkNwSzT3OkD+S
L0vmRYn4o142iCXnsFANzyTam66XrzN0jXFRtC3bGkBZrw0BWrK1lzhZsmK2
LzkP8m0CUvXyx28+P3t9f79YMV4KLxCMN6KeSwHLkffQuxE1HPP5bMrG/Mlr
1C9SnqrHPoNS6K7kFBqxUvY6ks7p6bfKYjl8MA3eW/fXFQ6t1ma1X82+bTt3
eGWLLHzfw89+vRw1lF3xNzLyAGXtJzMiEd9yeAnJ+DoVThnIgVdEXwdzoMuI
cqmomVpi80M9qBTObeV5MUrrm0lgEsR6BhJUYKJVFTGTjVssjK3maSjob6Qc
Di5R9ueiZbnv6YT+h2IM0Lj7jVIi4JuwqcEtfvSBWc9QuCNmaniLd8QWbPMg
uBYyDfH/gd9SIk1u+dVr8xJG+wWtYOcdXLMU3kG2jxvZnAGBZHezEtnW5IAS
whbFM5lDviPG/k/MD6HGwy+uODj1vkyrxsM1hZdiSvRBJ+bGbCyGJp7tsZ8C
XVFELIRfDkJPuMZViBjNiTbH9CCWTrEv1v1/ycdCsbSYnVASdGtmKK+m5Uij
XDj7pvI+hOZfOsWILGPdkzcgFakTxK4AsiA6x7sjUWIpN6x0wvQHFOMvc42o
Kppdh45r8rrnkK97hhu2ny93PTFwchW93G8m6+y7Mw7UTognaUqi9jqEB+UK
Ud2wSxAKAAej4RsuG34nVQ6ZSjmETyNZJS7Is0j7IvOc9zuaJ7yf0TwjqA7c
xhL5LybinJtNVqbSeYStT2vlyYnnN3xiuHlwXimIv6Inqb03JWPoXONBjjBE
j25j8Px5AAzbfNJcWgMGim1/mo8Cb1tf3UyFaRb0TSVxfQuOr+emGDUTYDXO
Y8VTO0moER09pmMAmM6IDv+dBCgqJgP/RUzvBKE/dIwnaVpItKoKxhNXDXxn
3m69sg9f0nnQ4pkmk4vDEtpLDNYd39Hkov+9ovaUl9iS/Fv1JrnrxkCXtQXK
Jy1H1rwPoVF+TgVrcOzAt6C+gt3meohCWB+RLfVXTrDoD2+sewCXdv0nef91
gL90T4K9O1QRbLX+BqxlLQ8/E/gXahZTS0x1K+86AX8PLLokbpTyQ1P6NEES
TgutCYMKrjm+S+uvVPriNtTZp2cdFqDE8l+lAJcpPOQHO0ICqp1cpolQkztD
FlEh/+Y1zBRQJHDAsjTkR6FhZ6Ez87Cbju5tG3gZy/ghb1RldaE/gn3JDgQ+
08HaUkUIcXGpYcLCfx5S9NrvJcP2N1GNeiUZwgVScd8SUgygN2jIirGTHdY9
1eHwBDIC8eBqa0HAtc8YqpbhN+0v/sziXBDJGyrZjLIsBp4V5/8MKBJI2EMD
v3KSlTs+d+tYFYlKAF0JQ7wyBxa/YPxuJBVeo9zsctL79T1fiNYmsbcwVvpA
9g4uEIAf3PvvHy76DUXbb/X+jEIrEFXorGXViF7QgOszT4YvXL6060pe7EL/
U6aotDJWnj0dy4w3yOKHPRb8XT0CZmj4BWqDr3l1hlGCzNZgzEabROh4Y+bj
U+ZCjXGLUSEZ65yJ8lCam4SxvV5DeouifaOXCrUmCM40msddiu7fuSakkERO
fSjRspV/7x8qzZZbCMRu1VK9mv6pEL7buh+/EDiJp/oYuu9q1jTFrxgqMBEG
g61Rf+925G2x1pexh7v9daMSgu0IVWevGfOnEKR0fvU89PQ15h2B2cBstPgD
JRoBNo7CRjWSZXTVKn2YdM3jyFeUqxsn+DaVBfl4I0uDg+FUgjvWX63nzfvL
XCQBLg9lW7onU5eEh/ZEzS84kp/+7JhjdCHh5nCthKTB3CVjpjzUJZQnwXaI
ErS9qe9rkc33mTdkFD+i92YYaY9ILtg2T2pkVxVAaM7cZ2m2yzd0mrznzIBx
1+X9e70H/C/rMxqaRXQQUNRPIp3LEErNqQUzopVke1LUvaZ33H4Q1KC7BVyM
Q0QS8w8Um+kEbD3NJXMMo8SynI+rJKpw4an/m/reLgCeFmlsfO4F1lveDaHb
+2sqyVPhTKe8JmGCLD3yCEEPIxOjLEy0khupuQ3kSMXjguS9hIwhUkpzn/jV
0Vtrs5IqjrjUzqkm8svUqOJ5INZoMZ9IEC3gIIDiOllm37mh5LNQz38oAFBV
IAAiit78p7Qme8B6gHUdW2xdPDW4FKVTZfwAxXLK61MaJpSGrwH0a7SG/LHo
ETF6IaiH8oJAb5Jw8LvbbL99OROPe1b08i1HB8QyWn6E9hXAeg+q4/mVGKwf
PU+2Ts/J/CTQp0+7GaRiBgD4i5dAd4dl//lL/GHUHmOYQEYfS/MTVEPdPFTs
M/LgEKscgPm+p+9YSMpXJ4t25FsCQ1bbQ6mQcU2CqfVEvVztjhbGjV12dz5L
YomHm6d+sXJ0YItFqUhr+qj+QsL7FkbCM7KJDZiZlLEVLo0zV+7ubDrWaIG4
qJ+5c6vPlXNMtCG6f6xtwg9Cd4xYlA6FnxQi7fJeW7634BHuwcpjlMcSeu3b
TPARWt80mmk7cHlJ0Nr/IGFvifqRomAKDttyY5hDzULv4CjWLrsRe2jYNjZx
g/aFxao+s8MNA3iOPhrzpACX5UDvKMYymLldbxk3h7vhED9LJGB9OzF2K/ox
7UtM2kvf+OVGO8EacoGJwnD84pFX6q351/1mEIFsKBNIxeeE4pUZggZLM2Yo
S+fyYxE2q4DkE4xV/QNdyh7GMmzE4gq07SX14iZxQeZoBgVkRAHbz1nEsAzT
U9dZpVde5Eyza30IrPuf17BwaDOrmIXzAYnDzaOOa0YcaAc1buVEVYNQksOU
nTbBkzklM0MvYS9aIB1hQESWBSKlKez2NcJ9BpXEmB0gjNILv1jPdPPdxac1
4rCAMPqKlVEqWMl7LtXL8GOy5lzJAfNKaBIuM6QahbUKvDg53hjOEbKrtj29
0besH6oRM9TzBk45zt+NL4vbfMLe3s+nADFeFylvU9ET02/BB81KGzkuWizt
XHg4v/gjODXvOrP4qAHW+oYCP1v9uOckU9dmcrvM5YV+fBKqiH1twGKAg1Im
VvMykGwFRIv+UlZvn/E5kaxUHFGobb4le9GiJvUtRUZC5j7A7kGAK/8U1gyc
wxAyWQOnRKm5Yp/7K8+HnCKV7y9TXmr8h6tCL4zewMsIOTv/CkpKYGymU8eW
zs/Vjzk9vu3kthc87Gjg0zgqklbRNrtLi0OgliF2DNhoGOqjc0VgjpfCZY5u
RTkmqADSAYmuiYlH6I8TSdya3uKqoed8JTxx4L+MIbRUxKKJSw1SQxMQTy56
hWDHj985i3P89u/r1MTrX8ny5YzU6VK3SXFTFmgzd+mczTtqZ9ivJV40jIpa
elO0K8mWUZn8PxH5FfK5pxxYMTdNK251gMXUm0OtkDyCqJN+d0zh/xGbsr0s
YUTsPKSGmt2/5iTY0X2mhioIzz/h8Dw9HIVcK0lIkCOaX/tlKMt7XpqBO5PT
Ygh5I28reOIdMi/UxN5cA0r4eqP4xkZ5184OKmIZD/mwEXZyQEBMYZhgwKVI
Kz/1rNUHaASZ1GNxIHnvTEQrYKMSGNowkjZbiUOI2MZEToEmYv+ydUu8Sv/T
2CihOjqdisyRre+lfLhVgcSwsY2hw+6aXOPnVVe5pu5/mD7/LXcurmCSeQ2U
i73FZM60ETsMZuLlJf7Rm22qGZn9hk9AXnm6XSfDb2WrOTENj7NCog3wU6PY
cz0lLGNhUjdJ4jaAqx7gYg/9/7jfujxZcKrLOetJw83y4mgvMatVapG+7Erc
hl75YlSTjXAeljleXpDZe2RyX8KXCvnNLL/jiCijRyY9GDTPCiIGsecuOjqJ
lCs/5RF0tMD/ydIo5S10wHs2WfCVJAVscAfLLHo5CO+m/s3cHUnf8HCQoPtO
HDBqYLu9wMpbSbZ4yhghNOYJVVdEwOlZM7oRgOGdfOGflueLMEmDBgzpsla4
7Txk2x9qvN9brW0kuxX1WHJNbj9XmtMBl8VDkRNaMfzwxXTjRyk+NWfxJ+a4
7W3Is2PSvk68AgHPjAgAwKhrGpc5d0WQv3D046ZrwWs3z84vVcqKJkhZ5GQM
zs7/Z96qtbrLlNXS6b0Yer7FRI9ihbxbnVW9US8Y4U/8ktI0mkJVQGBQ7y1z
YK9uOyXQEIPaS3InqHYOHs/S07oU6/YZY7TQBFdaggi9CuWIhegHYpLQP4KH
7XanzCfN4n8QN281G1IdrqA24CJVx08gYGf5/dCUxK/7k/5ywA/S0pxzMDYH
B1eUJeISOWzYl9+UIheyFuHNo3mGNcDivH5bhCsyMlhz9fgbX/M7Dl7bxcmT
bfpBx4dB5TvnDgDLgqBh9SBIuB0Lu1/K7U1PF/mHDxHcAyAAIy7Jc3lpXfM8
c7rGzQ+yE6exqL3LpV9hTZCIRT0QLpMiKtgS4b3aLTBQoeMhTfgeqL3gEt5I
1P4MY/rFLKTGRuPWPmUh5WGaW07J95SRTX6ABk48g4QkzMzmTwY0V872iNcF
8rRXwvoRw7s60AeRV418TTj/4ySdXYXthNB+DFyjS1jZIowLViki23xgXMLc
WogWA33rgjcA2+5j6TOa6pWbBZZZUsrj/u8eRBLbZ9C5THxcJNLy8CGUEjzl
N611OtvJNljlBEe5w1WGvK6F3H1omasJDyPD+uyZm2/5O742OmjtopJ0Hmb6
QUJCdlooGmV3jwKZSf4gy4Ouqmblg1lEkLzVH7bMspg1OyAGKHCyiHLtTJU1
pMVoxq+CRTASVKN7niHhvqEoVr+cQ2z79ri2FOcuREGKtts/VVD+A+dcVvGG
nyDb0KbLtGJbWDmH1NiPHfrBASBsmqpjwmZfu2yImnY1mURpjnjOUIYmgeWT
Cd9bXznCiHUWbavBZ+KAYCkO4M4aQ0ntAnHBMryCBF4vEU8+mzHxxs1aAO+B
yOvuCOXNnwbVXzp4r5cHK5pbVjPFZo4wCHJ5qH4xvyzvmWYR/h8MtRLYHv8f
rS0DnZv0HsqQNd561CnTrxqD/VrW7uMak9eRLstb1dkPMRJ8o6H6oOn+74TZ
m0rDf9072PeYfq8CuxXMVKitQLNtblexlhSmTPoPl0KEAhbCVsRotDCCefxJ
1yBCn34RWRxr5kACGebnLjR+hPj5vRJBempFh4SPR/9wj3aMmxeTBvxLLd9d
L3ZWjivrBQJQ1XqAUdfgdGsV515PySy32eFD0ZEiijYbT2AFxIZID2JwIhVH
6PJRxgy+pA6LL8tgz4ynhZNiqCTx9oXY6C2/q6wZAr+EsGKrzez5I56fSMBU
wBP7/A5SWXfazcLBQsc8ktZPd6UTaC6m/g3dVhotC7O7WO/Tly/yCpzcIidL
HNogBye5/5V7O1Opm78MMbv9QPTi6gedeqY3z3ltO3i3vVUgPhd2+WQm5lPz
MitxWWK3Wv/XCzt2Qop+kxnWPxpCeU72gxxGHnTaqg2ndF43SmBvDiOrJPPV
07r6yPK0Q71IlzMXY9fHFt0Rmd0lY4dtlHTE4A9/wTFwNBQ0ozKfTwFLeYGl
zjLufadCIbqSH0MrjOIBEm99zsvvVhiF/dmALH3L3673pdUbbmC00W05pWS7
VSxKAnWkUV69TBjzBbVO95jxln9uRbhTiios6HTsY2FB2CLLDVsyDYZHOCmh
Yn8oqoO/OSOVbC9SC+rk2OMZ4EmQqm7SMycDMUB9wcgSZARfJw5rZz44k6qw
cMgfgU/Gd6hfXyCDOKEWtE5WPVUBCYs4lGOPMS3IgmGKWX0C6H5VH9AA5KCt
i3u6M4IA/ZyT0vI8KEFnDuCjdJvE9zTyCHw0U6RtrZbDQKjYGAeXvBH8ZBd7
jQCsCYFpUbQVq4WUdq3izc5+S1Ya/nhYQyLQrjXJ6XkUZ5AUT9swpZ/miD9v
+823p4PvPg7jCuyZZphqZoQ0saePd3aKg9fq2zHrnxCz7/qTpBRIofIgbyZO
mPV72CaAsaf70wNUMuPFrpGZV8pIz4ZGq0j1woHPE3twtndM7jHhsH161afD
RW32BN2Zvty6tOQjnpNeUYtPI8k8rT3XqPicps0+iDR+Ppwyrq68MiwU/fTL
ZD0t8acH2X8eoaTIwZvpLSSEnglLakDSPMpEvMRFls549TnDGpPIwRJZff+r
9FAuSv01hYlR3ovkJ1K/7NNLKkliZWxvLjwwBDVPioaSp88hJil4HBVJOHYD
GqWUehCSSNONkwfSApwRsM1SP1KnKzIzOU47sSiflvq1kr+Cq1rX8hwFd91z
S66K80qoEfsJ9Nbv6kKp4yRqfMjzX7WnMU/2VbgFEzqxczq7nO7qPVYmIkxw
09j2n4TCJJNt8mt1WxHQAIbqK8GtnBWYxlPzbNf4n9ogUDRm9FCLdK6gkr65
lQu9jdaZXltRSv4D2En1g/sBJ8i2TI2cT2RtWjI0/gqUO2/AEkrDGRytYkX+
xQi+xs7R9TRSIQ6q3pst4QlzwY/ztoWZTo3fVKE+3iLK5i08WtZ4Weho9ezB
9vroiZ0vgpsIuVkk45irwRhrgHKuG2HkNjQEcBX9xT+7cYwh1ZxqS3qO2FoT
0+A4ysu97LqZnJiIcVlrDWWaLmStbRA1tNPN4iFbGMyxOs5dtw1uzYUSLZ45
xJ24h6qe7lVqU8ZxaZN/qg/9hFls9eBl4VS5FWOEN9BEsgWHQLjvuHKwDNdi
clURBqYVVCKaJ2GOmY1yr2hkWcQYwuc1kvsZ16UfIKPGA2CSbMiUkVvepN6c
4d7y2YCLAAILONBbW9Efq/Olbqvhv/TEsffdCFwJtp4wAlz56oOaT0Qiax2r
IRqo7BXjloPH1S0O7GjhlpgCujsbhD+ptdg/DHk1onBpS6qXC8tED4D/GBBF
fnaJTXTlzK+qc5WzPASqpWWfSGLlsf9sFSDPymYJIiQxpNicnnbAKY2M0Dq2
vffnk+QorBYQrnq1ILG3kQBc+FTBPFpRDytkYfM4AkbuMEQhyaa1+sPbqCNz
9dISTy7PYNgmF3yji1eJTf9nyYuM8GNRF+FDE4t3h5Fme5vpCteaFGmvKf3B
vNLa2KBfZv5f1rdUw+CzKlk8SKXpxINgodO1Rej7jvcTQLx+R4nANr7hKOef
GJMBsaoE+W+j/9CBL8A9dN/GG+8GggzFEfnX4B3gNO65m5nDbofA5LxLcjgS
ZG9/jWe7S5pddcP+LxuRzYnuWPSHD9lVmwQuerIbPFH0+qT/XltRy676QXfp
JJkAHSrdCUeEZAdYAK8a6cJDwc85NE0cVwywGMggNUbQ8vNVJoHeshJFMEES
luaVJsimPdBk3rMl+jzzD4qtEbVtvyViA1XccKoPxpFy2xf2zB/OTpMAxDjP
hOAMlJC9jWAFtMqkqLhiNF6ZUq4qS79+uRB6AflPiQZ8RYpxZH7irbAWkSVS
k1uROsi2pnY78SVTSgNGZG2JWAgT/E75heVU3lL14puXAJYJ6nuv0AN5HVPm
tb/4qatF9Ijc/mehciuIzc1mSJW+DJrKXfgWdqn1n6Ewhdcw6hRL6S1G7xd6
CdlbyPFIKagUlXOm7VE8f1MaVlttvLeLsNA5XQvh14xDDfbbbKHK7et/CMbj
ZfGqHBw7iW9cHCrdH0pJk+L7yEyDGSulzOFWVjafmgDOfOBP3uvlmk6Z30ao
8gTxOdys2p142aGysR/8g6/eEoW9hrt1fCOPAcSBxAd6dDuvRVrOkmroP+ch
+kkkVy606I9rQuBeo+/0UVeK4y1kH4L/EnNqz5llfaxfR2SgSuignYt7zPqM
JmZkCACv5T6cov73d16k/OmUKfGS4Siz5324Jg2ZqnMSTZAED8N50wIP/Czs
IyNJI79jON0wMr2zumBPD/w3iWOIGNQ6VdeKxDymeNWldvoFIgKUtsMxggCK
97vn+4I2PnUDfQ5R6h6q8UpOYpwroe7G9DjVq5XIhcJu7RAYDCiWfY5Vtbdq
L6ei2Wq8wfLN7SPLI7q1/axzHdQBYAWbpFa7649DTEGsdfpQ2ftw3e9ewge2
QMGhni+Wvk/Rzo8m+0F2Ob0kFHOMj50OJWP8nMnCi6jKM6aSYfYT5zVWPnLz
pnlzfMQ302G05yZ/Kk4Po8Z4eLeXBKeC4Pry8xEKgjU+zMFlPfSzowCwcOqM
PcfCJSVPntbjQg7B2/BxyqQmx+MHOsFF4ScDWWKfCAnjXcfX0a59QlBfZMFz
8g0y8oVJpznfXdbg6awLaP0VENgGMHiecRqfNJtOwbAdeGY82xWLvbv2ljyM
KKaHJ+oOw5y7Ym8VyAwFUkwqUkNhtb1rqrCQhuTPjAgu2Cr8Xg6/+xu212pT
YqZUpJ0IPJgAbxLgTHGuPeSvmcLBywiKxsKBDNsfaGe5RuacpKsA2O2sNwwa
r4DyDyfG8v6sf+95P5ZZ0kdetxqdnSiGbszR43GOCAAu3WYqI5Gos6FTZbE2
l1RdOxZMWHiv+auXxeCT3dYFMUsNxOqBiaqPu7uWxIVxPWdNyfBoCeTkFPzg
yeA3/0TmkMxhBiMzW4QBvU7xpbsQ/pHfCq6wEXTE2cN02q4XpGIcFLxenAYP
MXhXc/l3/Js4w0zHrzpQHWaO020ey9nIRwrQTuLzq0CKCPC5emW9n2r7i1SJ
VcksGY9PH6O3LE5K8+j80uSNMrYD+KSGhbO1bMaUxrwxTLKnLjxklFG2Nv5V
ztQkNrkwyTGQQIigmnt1+F2kRyhhtNdWsEIkcehRzwDDTzSzrijebqnKMASO
pTDxS/8JEhUD7QVjGQvoxix5Ktq2gUcl3Nrz9fZAsBmDDHeClgHHaf/eAYsG
c5cA3IvyFeY6agc3Vk2lzb7+7rKA5tZUdIxFdWtUTB/IRW30CuHssbFeL6PO
wHqVkGv9ud8TXVa+id367CDApM6uP183blNzVc6Q5q5tEGT69ev2Cynw9OM3
IqkIyK1tmXfb8aL7clM2ildUWkiIfHVO5VP0wkVyn5GL722IhX05qCxpGxAH
t86T76MVmA63/VNL4kSOzKbwIr2jSwWYE3niKYmxcyLAlTKBXqbRNjwh0Pfd
ZCZeuHKNryvkZTHkzIUGRfa7ULtQZudhLcB+/sbRyvAi/CHNAIXcJStaSYgT
h1MiuCqOZ40na/dWY30aKAWQ/+smCoBDjqDWwPyylENaIHMM/ds5ZR+5aA0F
yl9zs1gKRpnspRQFyfyLFIUYKt2C9KWdUmhGilU+fMYVMgTIyq60n3Hd8EpU
KWJuDu6Glljb/CPDyAQ/HWznUzo6eX2mEdTfxMBRip+CoPNm5P0c/4QCAt1C
gpo2pDGe6j4cF8Vru+1i+pNw0GilW9ZzwLVvwSdhOzNGkQDv8SU5b+uIJR30
1sS5uD7z5AH9iEVEIRE2FYcIBf3hf3pG2MNeEPBpH6cVDBzpralcUdJdBYTT
87IfhNE5DSeY9c867BBIa2FsH/UVx8UuR3XJRLygJB5EUFzovcrxnx4Mmgpq
QYaIUMNzi2CdYoROm3BUf3qiFH0eo8Es0cKiXgezNNqDx5VaX7k6g58p1UPg
cClSfiKv1bLk+KTOdVmiJBH4Fpw+mmudSvT6ZQZjKzhCpz+6lxxjq7F1ATK5
66q9UH80taCCcSr5wgQySP835MlknwnGDKw6uLUlWNM5CYuVK4ld9yL05gi9
VXlWQBTUt3QZwMtIJXkWek1K03vumaTf1/KQLVH5RPPgr0mER3UoHii+idGt
agvcl8nCC0k0DOaa13U17gGNrkBXlYkSC8lluiRllTmwv4OuhLwChnRtsLd5
0isq7XZnXei4pfVUYZnGlFMIkJEDNLRhn0V8alu6dyqNMYx/lLZV19r/60tG
lstfEKpO8KJj7eFtaqB741iZHF+bZRGLoVMbEX0hg/EiVE3ZfmF36s7ovwjm
yt2fiftApSjSjsW4BdsMANAHJqRZ9HqEQWfkaNsGQnlxDeKBOXITNTwgsz/i
EK8gmKbsPS73JPADhebAFI/IrfMG2oLBobTW81QB/uCH0/QeElEjz2C/eC4L
eKvrRU4aPbYElPROBsR5slUIZihJD/j/u9YluKGlvU/Oz8ic+Phd08UZWVTb
Pq+oNzDlqXLyXT/itSMpy7aDrf4odoAWZqSETSpoV+X/YWknaX2i2/7eJ/Bw
HUCTIh1t0p2+6GKp0Mh7pamIFUSO1gXva33NXEobb0wVjKg5eVFRrkB11R1W
q+eWceZ5SJq7EumatQq+e7pERt7kckhbvsm+4iMTSYIlW9cUbsqccSe7MVV0
toLEvvp7s+G5oUOfYHXZijZqRvXozMet9R4wOZza+FkWofeisILDl7LMTqgs
z6+PjO6XVmxgxK26T6laZos6s6KGndVXPRAT/GiP55y3QDDeuV8dbOYklA8H
SICBsd29oUjioVZLmp0Eb1+ah4FFcLtaWPLUQOJXMTm9nEBbnYbkkzcVkjGV
FLzGZ8WEzgh+wiXxvPjxtNVqBSXOa06kygHe6C/stK+3Xl1RdN6naL13bwKi
ofiVnq1zcY6p3kJ5ppApWyozqqbBNmlTDii1B+vJC6sUzNkIik+5tM37OVgm
JyrIliGjwq6It3ySyDum6bcTAPlwWdW0YJ1Z7YNMd0qB3MMYfILWoTarihpK
2xJC3qIcnFu1QlMtqKRLnV/rCLrMbnEQVPkKiU1O3sSMzHCeWcjhjMwvEscd
7ly2ASRi4N8e5KfWo4ZlsE6qc8Cka6dc2AXuz/CqkeOqHNkL7XHm9KDJ7SUL
vdggXKCmmH+M1KDbN9tGJESL2sc6vj9RU0u/t2/GolZYsIqntDD5d7wYUxjl
Dln0nb15AwARWGksNoPgGVo84VfIvoGyPTsEdZhPKCJE6ZRD6qpYNBBblnui
33F1iqhiVT0iZZ9b8oECaUQ6l7NmRjfA2mUdxQyJL2UG4avVtMYusf7FfeZJ
DIHJ+RaOSUSI0PzIZ/jroHl8AbITxqs4d1mcoXgBBj9SzYsSoqtel2P+p9Dz
ncmQ14GtF6pb2ltqThuVo+OuBfBC55LlzkX99aaGJRwoVoebpAfJl9/Lmxem
e20AzrnylZlJiBTLJ0Of/rrdOuXb0yG5JKruMvShGi4cvB8CBcv5PIL8S3LN
yZT3jF3JmOQGVdLJJnTnvNBruEDN4eiykRkXfxPL16Wp4iLLH3OUIGWHf64t
8vnH/nYyxH5F+O9CmzVYEO7vHSA6t/3EMs4wsf2RQFACRLu91Py+2sEWReFj
zp2Dd8PUtfjBUgRXcnzfzW7C8RoR8GfFCC/CSIECouWezsCSX/aSONJbm67D
o4XJ3SkZhr5Ex8XSOu0P2cG7Hd2CPTdFUQzxVhg3t7Q9mi9Lu4nNrnWC44XZ
nXNNLUIa1NUo4Pjnvhp9DWpQDcvml1l8jBtEsmPOU0lLuQ3UmWYl+GryozPB
lllu0NHKzB3mSDdoaENlg6ifVm1zL0bSXCwT4BpNmGJXXw7IQnGpjsd7cHx9
9dkUVM89nkybp0bz8lXViv/Aoch1RlcSOoBvkVCM2X5teATvAyiWMmu6R6xR
JBBukRHL9eB1FCHv+W8f3kUop1/8PKIIyzkAMj42k62vinMiWJ1aUKj+QyeU
1yBWHWQ6XVxvcnsfD5v1+HZddgag8pePYIHQ9KR8zobYMASvZ7uC0AviAwXA
5qa2ViiVcztq6Cbuha8jqgZ7oUA5b4EM8Zgffhbuk5W7/boiid5FOCuJjgEm
hMIaK66kZ9Oml/I0TjAnO8lj80U69BYl8nnnsB/GLo2VUbj7tAuUPDtt2adI
h55nRTgyDOPO15S53V6kBfNnqauiXZxzLp+wX4FKeWCJ7eBMm7NM9Dd9S+65
gBVEFVVtO0+U3vZb+gmjQ9q8d8Q5Tz5XWbegsE+g7m4a/RTz/iUUVye/mkeJ
U54ua+H64IVVK/++GmnlgMX79gXV6kUkeDiHcmslZp60KYq+c73RrTwTVsKX
q7pU/BIQGoi3UyMZsq+/YVEwj5UhidaWyv5lSjqfqBgH2AHMpVnV4j15Qxru
ngHel/Y+sgosNfe9VDUCftPUbEKELA6JfQpf7xGjx3zf4umi1ot+rDwsSqiA
/2TqkgGe8fwWWvddGZPIZpkwS3wK1wV89lLdJ6dVoNICrL9hUUDyzTKTMq/b
8Ok/IeHGWAqRf3g/NaygVZSCEbvpqUH95nBwJ99OPuW0V+z6lRq5PnkztxAL
rjhuaNmV0qNa2lX1jy5Qt7rtLnvzkz9rmgixKjIZi5wye332thDALCWHFtGH
awdLNbAHEoH7D4oz1X1hGok8iSkk/Thqko5zck4jlqlu71Z+LaXtVgsYIyAy
wdtxa8LWViOOC4Uc/fUSwmNVRSsG2C2AZ9epgevWPTn1SzZ2V3n0Drqn/3NR
kLZUOCFcr/iXn0Z0BxZ0V+AEB3WG6aK87zj9cmw0p1KLS6m1wNFzYpD4zncc
Ys7kI8PZ6Bj6KZ/3Hak99mGuZkjYY87SUoaWrg+S1wNZoBefc/L90csjkTlP
ATvV/+Pc2v85yZ3KRmRquYqRAaAfavR0eZnyJ0JuB6cYWAJiNRgE78wsak3v
HLe1I0nhm7VmkhzMrFe/gG9kABWpZ1NPDl9fAwfGmXRmsG9Y995xo8o4Kcwk
GviFnPmvjJFk2XFCj5atw4eI/pOGYU6hKFOtny1OZME2fctaMvsQ4bxpDx6O
IG0keW5lOksiJevKc2cDBgvxEq/3EiSSIrUF9ZUBwrnXOhOC1tv7Xp/Zh3SG
apukeHmhBQnBD+vNcbtJ7C2ZHt3nXf+mmViOUYAnC/eAGoIV7nslIICh5JTP
rS4YPViui/fMHmiR142xCvO8cgtgn1UIdx++Fj7mvDM0XnOaHMAzRlUM5399
aThdqCeIFt/9DQFyIYvC7cGRrjukXard5vjnqVe0mpi1QjGf4jiPnEQt7UR7
eO7pPblFgQKzL1mR3HtkhBcLa9cxHvMdpBGF+vWZdYcnKj3ICJkMZKULiXaw
949BkDRBaava1Qwip/eHQlgWjgzaHTO2CAhXH/SJ7ZhpBeZ+Mgnj+iXO7de7
8ahCFl9oY3rWxospxucSsHxwNq+q/4CFGTS78mc4trYGedMTHmisqSeXGegR
aYTcK/XM71ildYU9LG0Y1dIv22QHWv8tRbztH3dPd135CWnkTKFnTy5BqIFC
KxlQRubZ59ttKvDog+l1Obagm5t5hAnQscqHbsT9Iv2QyGjN0qTeFzQz6yye
uurlDqWDDj+l1sKWk4EA5rYMgEcnEBdgmmEBvv2l6whtsZo0m3w+mcyakIyj
a5I1fGgcvmU6K5bqDRy++Fh3u3laogehyC35FOpFiRH6pNNd7fjpOgt+A4uD
WUJSnt5jFSFQgPFYP6uYpDGpmWWdTuLap8oMCt0zuX1J1LBU9rhgGD0YqQLx
2PyBd+DZJRyF1vkqZp8YhtwTZujzE9pyR/aM89yTURnsfHDYTG+gBgPf5DpO
LvrcI71MQhZaeUSOrxdUQdQmGGgNlWvNfXgw2IdBJgYU/5rCPc2hgZYLxGcX
d1FshubgkBt1xFg0Ar9B+iMVmcYmYLHvTndUFKDkly1rgGZg1tkzIY/nmFQo
YITbX83H0f7JmKjfRSsrikwAieGea+QRXlMdrQ8KAl46CEjFkWoyeORx0w5s
KK/zPXGrPh5b8ZrWjBYzKdi0JqMeuLiqgDHpADeftyi0ZnXE12djjJaW0g9y
BhCLwY+e8Tk8UDK/I/pcZ6RIjnjetHWdC9wrcSSC78Z3lOlzRuyeyIqXyQxt
owy4ezirqS6KRtrjpqyzbtNu2VjAEyANW40kMBZbwJ98R6prt2x8o+96SCi/
0/U4zo+mVW77jUd4id9WhrPZw5JLzUOQI8Lb3KaVbl8TNfPhvWVj6aCyB8Az
6n5p4bLdSfOtwLvfeTvfBOiJMDLTSDns0MKtOzH+ULGVBhZXNRTkRxl42lgk
9sqV56SWQM6Cd9fuF4OaVekelQRTdrSjbL2DwuqEAZONqN6w1XYBPhPbwSQt
bQU8AdtZIx0F2aD/QoYzSPzAJBcfci7mkSbyJq1nmMQzRqj7g7gVSNh9+zck
EmFE8lErqHTQnCwn8s6AxN/2KFDKtBtisQxrHmIbq8SmcWiV3PMVLg7AKDMi
7gk06IvoWz3++VAclFYx1ZlRIkBEp7ytdkuI3DJcpz/48K6o8UDgR56Ty+fk
NIPDYrHB+yjIW1TQwfsQ+6Qn60Atz8u+2S2UKmjhNlphqGxKXA4esC+/6hCO
TZvNHrUtpTfnDgZh5eXZ6bYsQd4IR6BGnsDKQHWq2onNwSw9Dg9zZZJ1asaX
R6HBPIGFCz3vcysOE1w92KKgGKIAdE038aXhXF7FU283yg3DsH70BBbC3fhj
FjJ0fGz2yw/OXdavWvtwTaZYEUseDvvvWfSDFybMX8yLNwtQkkU/Huvl9eU6
kgIeRLZS0gaHg6yUEFmMEFGunT3iLnc18x9AHlvRoHeIe269TGlHVn54lZ25
nc6NiNLVuL+aNMINYUZ5aX6JDMWoNcocCJdU/Pc6E1eBqRvT3SKeoXPJXfm/
xprEN5uFdjPv7dcoHCtpOiCWXDRBwsA5dNOVIMxign1sUExnugjMrdIiHV9g
aUPMnKqZ6feitT/aNC6GdE2tfDfuS+c1BQzlrGOX7yifIAs9UNrQD7tD/we6
UkjpyypZ0F27Qu5tUIoj07wfwpYXxRFAGjz3V6Fz+wbKCi8AntqCnouR+cTR
HMh1gEKXOXzpSxJ9iacwNxBIdi5sq0r3kKRc1Fe5EWMdcb3zqNpOCZ1lEWY0
6hcjtcEhzUBTcJ8ZLHCMQ3BKu86KUZO8nRg1fn9Qv4X10aKRpRGebWnnIyv3
jirRGFMD+YZOnRFepd4LpvX4DBAjsNANcxX3zwbujm5mo/K/zYavwH6vEc0J
AffJHk8KOb+p+LhsdPjePYG+eI/QjOQWNXUhrNE2TjGE0TSf6X0tm0g1Jcto
+CPMTRgJgkpe+RMhFwvQbrhTVHjIVxGTPf45svuTBloMtSGa0XOv6llFBEsn
WwlI3+sxnF+CfvvXI1zFfNqV26WP0GIq2rMZdoYN69WRs7GNAVaBZLcN1tJJ
BsdjLij7LZbAj4W0ovAhKR4f4JZOucPyQ1FjLMNtQ+GyZBTwCA0evoN3eYtW
/57nS3olJUanZkCoRxJscxJQ4aBOk3nOj9as7zh4LgWLWwna2xUwHlPdT4qp
SFHfIhng7+HgCejVL3kyac+KgFGLdc6YbC1aprDv10v6xo/jSMjB6J8GH/v/
GdxqrHCfs0fF6UvVL3IuZMwPfQ13ZqQ+94+LRwKjkp+ssqjkK4RFl21mQFdr
i/bkKYyGwkygQmJ9r1th+PX1qL8OWy0s37Q+Fnl42ThsAM7If7lESPYfuZVx
jo/OmrZi9VqujPJul+4D266BRcGbck/nCpvR5zlsBitoCNwUS3xnheMuRT/Q
ht299XwqCwi2kOTba89nBl7/aFdsMsbH0IUvojjuavDUoliZFK8aoOMX/HXA
NIuQwvLyaqjV9aOz6hXVHh+rVqqvysMFYnBQcC8/bK6XA68kTsyNVqclFuqd
r/e29jTwU34QrT1/CwAQIIoEziyplc8t5Op3JQn1psLVMjXObDLHOJw1FZ2P
BHn8xpCfkOVLFNt/4M5RNAPHheQh3cTCILz9yHlKLQA1bF7Au4z4BFhIllK1
dPq3NiWyFWOMUfL11u1VrzvQyBt0DomFtClxb47WaW5KWr6Tlw0BGJ2EzK0i
5lnbnCPKElxaKXRZJd1Gr7DbL1EO8r6rVqtCOA/1l0JHTSVNYDoBPwDuOfpW
jW5u+QnQvXGQYvwMd1MDHLrIZ2S1zdYZJDeBwPKATkrZGUIAajKfzVLaV1qg
5LQSK3ofaXLulzPIc9SuELF2fH4Xox+q30pORdKd8Foj76i7675LbocWWurI
T+MYMR5qaw4ThyYfVKX+4oTL9znbq3Bb6FKoimrtUQNvA5ZryvFtfGSnHCyW
eQv/uIa0jpsDCNDqEjEBgLDdyi8GeeF8cHBCrYZV8gR9fa8E7oHt1j1LxefX
zSZK2bEP16428RFFTa10nHpDhhy6YztyLz+p3GS82t/UkFOx0fRMKj6wAn1G
fh72Z6K0LNVJPnQL8eH3GccaS/fnDONqu+c6vwyoyqn1NOnCIU6+K2kUFlb/
NK/rgz7om6eqV2G2LEAZ/iltSWKJIjQf1bVCs243r3neyTFPDMuDxcQfFim3
A32niuCR8wMosq84IAY39zK8x4IKT6/FG2DUAotIOau2Kka7u6OU76F/hHRr
tfeVbqwQ4/018u809ZN0+MBBx4KN6cTHLa2KKtZrPm012erLyEvyFFxPn2UM
GL1+ElHUlxjXLbjLwya/PYOeShsVj67u59Eur2seY7XOc/Ih0/Zu2gF3k3jr
EuKCtH3bpRysThwW065DY/j4KSJ3x0Hh+x6UoNWDaiPVZCKIPQWqEXG9LZlA
NlabuEWGgFGOhbga+cP9b+kXUKrSl0WqQl7FvkN1sM2tAJand7k4Jp/EIIqs
8E9qK0UAnx+XTBa1uAJj31uPXyQuYqiEtm8W+fR/kgbmu9aYuqA24gqFmJ4o
XHe0iWn+cU93PKFY5c4i4NIumkAssM9zVwpQKdEqp2bGx1fDZV6j961/LBBa
rVg+4wGJuGcpNsUkJG0aR4voJCwgOsa7xtMascVGmhrs8+wZREOaFd2DP0IZ
IZdjmL2dQroXN8CuQ+jmviiwlpgjUqGmRJNIekWXIWCq5xaDh4RO8n8v4vh1
7o8p/qDfBCqYdwy4ZytZco0VLDUggVJFgayeih7jhR/J88W3L1bPGEvFWhbU
I/qafp6pFUUUhNmPV2SstN+qXM0JvHn0cap4TEYeWFu9y70L7Hpmd1m5+eBp
fXf1TNjFpc1rmCt7ZrHSqgeZSzCjv0kq4z3xY9mnJnHNUipdCCy4yk7qkJ0u
Xd2KdcJ9z/BI3bzVJI83Pnqzkcrt7QWWSnNhhJnzq68xgikE2HwHUvu12FW1
zqiP4MT5njMWdjkMpzKY6Se32425c2+lcYyTY5Wgn4A7cnK85aTwt+Ptmuz+
B75TvwefmLVqOT5I2L0gtlQnHHPU7SbvC7Oyr7sIdWDMDukQoys5T3sLRYv2
1hD5d9Wb3Uv84XvQ0TOgBjEbogQFaaconbWvzdSzK7/chudJTDJ+r1j7sGSA
fhOgYFytk8WEj3w9CniFvGpbVaBJ49GP/PhjNpYnlVspx6spzZIEQwHgIVjY
ezFxbUD/kOjn9Novl4kv7WZeTLmM1U61rGwp5U9ybVXkKcMRG8lWTCDKSDNP
2ffzZEpuS8xGjLPVSU0RD6en+8xsjZWh12kLBaBjhpMzN3xOD2h87D5WIj1t
PO6j3aWD8DCaBu7FnBqWMx/cp8Jh3h2DgX6nUKZk0mJcfzyxTwLNSMZq5783
1UQnHZ2e3pB/U/GOuJ76AJf8n4CTVAUr0yumrgTZW2+ouGIzAaw7BRxjjnux
8OvRpmiVY/VrW47Z6AmnTzIWsOE6lNeJ3Pi7dyNi8k5MN4Oy6g24zpEKfe/L
nKiU1HqnZIPj0at9deEsK32g4KM7Vk0cyEBAgSTddOZD35k5k7AGXOGqbvgr
w5vo1ArlYgn/s+SidefzN++XkVDBUaMGg25eZPIPXyrWB/rn7nI4N8lBUSWO
5fw6cG/yqkVqCHC8ehWpIPi8catuci9S9soh0kABpMEFMA9jYbnJO2AfpWzE
fk+KVAmcCIlu2SoFEmYBIrCgmnHw24GCdyOs0yQjx2IAnfxjnucyEJ9zjm+r
zJEMdPUVVwk+5q10ZsUhP7iE1r8xbpzlPbeRVvSwocI8LNAYN16OGGxMM8ga
1E8WF9uGRsNjV2kHTwkf0hWoxBNTnY7ZJLq0RZ9Pgy+2L+xzyp0cY1pbUvPg
rSoo2l++4UcSTr79VKwClyyDO5dHz8MdFHXsMTaXwPWg8IPdL0q2CWi8Rlsr
6eZGutxH+vO1kIEfKOqlSaVrne+XhFRYmgl7Xw7c4m49IW4Nc2/K/Jvzigib
0UfhkqSwXAyvhpMsSZAL+b/kvJMacy57F2WOZkXcBVm66xuRP98Y3lqf4pD6
L3LKtd5JTAUT7wKpYlS7ssy6B9vukcTZ3Y6XRbn3OvH/QyGnrSFRJ6vQ4+xp
dJKPpPId//uwjve46Azlk0CbT6gR1OevSjQF9mocW3JYa9ouhWbCNYW4fMcT
Z9BuukdTRuAxkQk7adGLj5O17Sa9bWqQ1n5DIucRg/w8dK/3DAWD3ye+x7Bt
v6XEQLJH8E5QJ8lI23507PQl509Wt0jns0mn3YH6Hg2Erbpy+FrW6mzC6sqs
8eFHv33eFSOn9XCzjV08DueNiDDDfsh2B689cZ+AsNplQg+nuh52YSH61akj
5q7v1QtRHaAaby/r57LOLeE5exYRLiVloTywd1i9G+R19t6zi54pPeG05k/9
CE9GJchnpWtUDfJo1uhV6amvLRZmhH5sdbjaGROaW487codSA7f14A+RwQwY
5qdlYCDI3aAvi6/U7HafgHzkyA2hdmnBLNhvVHW2J8lg1V24V+1dwlbN/zvR
30q07wD+E5pN5nDc1y/YDbOdZoRU2g37g/+GGcPdXCPqtFBnmP3qfi0AVMi3
xLHbiHg458gNkl8dsSqJUpCvhbnemKCKfw3b+ukkz4Ua/6ih8/ouc7HXkhxS
pO0/zmEr5fXOfxf0H5Ct3XuqXTg/+hecpk/QHuE0ADlybO4ukycbbNMkGV6x
gD3nJ8mDCh5YPQnPPJ7Pg1qTlKvCrW1nknn38dhZtYHIL2lsZVW6QXeuyar+
zOYlXf5mG6L3nUWjcQCK4CZdi4kfwC55zx66ldARse80fkN154sMqR6ORbsH
9twAUlspQW32uDBbK9CZg6oUpSUPZYqkCjth5QfJvT5DQf2hANCye9Wpe6rz
6lidAOAG/VfDgEIuAA01FZjvY9j415fhcHY7VrP3zQRJ9RJnGvF78ipkHbSa
lP0gMADtsqtCPGhrTG2u/u44jswniKh/EMZdorPmT8T4Jjg4e4OssU+PY/5u
pYR9G2v9orprSOF3nDvAs54Q9d+0NtBQz4MCv/tUKCyF1MTJsx5oiuAf08Wi
PJ5xO8yAKI0jpeBBK/xpvBHtSrbWddMWql+8q/8kuWCLui0poE9QAHLoanz/
IZ4TnsBDgEC8OcmKE/cFx1KoBhUMYc1JWcqFDkGO/pjJKyUREYtcy6U7Tn6+
ah8QiBoWAelcJvaFwP6J/acsk7iOkUBL6MGJ2MkbaVme1j1dCLC+uvxF/0KH
AmmoeCM0LX8w8vxm3PliSODBpILNulH22/5yyUiOlYamJ47XNxZSTFm9dHj5
xswE771LIlsCnMkb0/d8DaNdhx3JxTyjDpcq56YkpW2nE5Xkp7NRHn+Sdn28
gSw+Aetjdlld80IBiIW4CtCrc4I5sIcK5ltAegzHkgXemQg2Sq3gC3Y2m4Q1
17LfeJFjG8g7tUzh9ulMzK7pVkxd+MB3ANJme/UA1x+IV480kY8ucz2x+uil
CJRBCDaw6ZwgJGETMdFID6Xz0KVLFUbT1syFyKcIIyLpXZd0Vh96mT9o3GJt
84Wg088B9DDqRpRt3TbUGQFYivSKiUMA3VIOJ/LQO387eXBDdtq0JGEZqvFv
2g7pWsdt22wo2lGQSHjR0OGbRB54Qml2qLbcSX91VAnt+Hu/ytQ/PL3qiuxS
4D6H/In2VolHMtP9Gq1dYYwlm822MxNF7WuHkd18CGIlR2DCWDNfP2bc6pn8
qEa4LNCRNc3J16unaTCwi94ealdvhCgnWtQ4z/2LFyCGbJy+sEWLIct3A/P+
6Kgr5o9vq4mYfiLaKDtRlKf+SA5fi+bm2wMIzCWehoUYjKujgkRwCQGoKnvp
swucZ81L4abxo5TVRDjmqBfysk/9ljIiHEux8DwKaimUZoU4PfcfLVnsyhID
k7HyDKhNAyac7Y9kwH0DhQoWyrko78k44ZlO5YTSM2AOj4/Zi8MOERX/1Ixj
4tqK91qd0JhOrMgmqlt/NgmoEM/Pnd9BQQTxK+wZ0XeClT34J6vPiY1amMqR
UY33TRUvNNoBT9HYCrKB/R5TBLtsKZnmWVwxidZujh0HGX1SJqVcxqW3823D
+7zlYPruo1GXoGDrl9Ix8CIXgnwoYCedFyGGztPZlZrogHgPdfYs9EV4YFBg
Dk6RfapWytHYZaveo1EZ1jJuB6gfv068JDpLokgn1ZF2YRaZgYwDdGdz3DVA
mC9GLteanhC/a6exprYvL8byrV636KiXAcdYrU0u/h2QxRRnek+NttHTfUqp
Civ83F8KLFHHMTY5+jHW0PfA3vL0hZsrIoaV4h3E/kur2SYAbB8C9v89GYxQ
lbMdrxpFXeRysAwicoiFZ5Kn+j5bjjz3k82WFhcTvx8tEn20ETjk+6zCtOlk
QaoNiST8QODkdOvOW2gvcilXy4ODfCATZX+JhrCKzo1Zxd2xPUwhzFINx1ut
ONp/iYz5NTfCb+3j6xbNZJC8A7rC6lv0ANTV+cpGSqRAFnBqjEQljMlTg4RJ
PYJa2bgyw6PM2RJ+0Wn9x/6ntnhgFGtSgRgEFFTgWhOQL0Qr35Do62qm4Q65
5Po29W+6ShGf4+KbCwV8r+gd5uHQiPSltKoHv/d+t1B8/A4Fhj/svoCG8kMg
drv9CmmnCAMD1Uh9cX3tlHvz+7VfCvJSakLvA00BhZOvkzv3wl0AKBugGIcA
vvDBz2t5c4BzMxF4AcfljRLhRejbeOfhPOF/w8VoEKnFr68Uwgzcq0vg29jr
/8N5u/3NdQEoxzFBn9rVSUF3pa8FuvX+kqtOvgkHLPT10jWmaaoBPAxNEK0k
Pe9zoMumYUK+T+sU2CRLzywMKdcu2IitMdP63NNiwnLy8k8gugEICxYuKdMP
XhvQnZBNK6ZnNCmCWdHN06IUIzcHyFeyO377RMAL141F9Nt8w7Bn6C2Owc87
re2vLiaRVsr/2H2WnEFo5f08VWTpDuwDg5nXfPAH0shCRWXr14VMiFMmow5T
9UDT7isN2aDVPhp7WUZtDz31bHJLdU/NfYmDEjyDex0e5Bd20TPqtcjfLEt6
2bvs4oNXlPjyVFvsiSZrRDMl3RbJ86w+i/NeJmqvjzCXcaMi70jifGiWzO97
9oDuvlP0xXJml2I+ngBfyGmX1RNfU6AwLqeJRDkEj4W1gNStFDkzZpuRPMeZ
qYsplb6sWMZNlBKF3sLGzxkhn2fsNHVAMhvlfYay+fq0Wjdi+X9gGbBd7HA6
UPBJkuW15gGmi1Hbcw9lUwSTY+OeM/Ar7udEvTi4OSfBu8mRqN7EI9z93dhx
x8fPGEEFOiEoeJB+CEAF/HjlG2wz6VDFBpAslLWWCnu46YghFGKAMqZ4+5FQ
/5WhBHDSpwL8qZfXHAfMm/kv0nA/uktXRVPwXtJ3+s1QbWWLCLwRWj87SPS2
0wCHo3fzb6yCUb/JW+G/tb4w4fLEzDkuqjuQrnhNlJURV5eSTY8tmVu+Cok7
N5LMk4k701OpY91pC8oLalGUY4Dibr/o61GiBdrTWEvUU0/O+4I9IduXLWg2
Uup/Xtw/45P+6n7UF2mTQsiPmslejG8B/dtQKUCc8zVPcH2oipvSY1OUf/qA
EM+vyll5k8sPsM6I9Mw6Yz6Ixdya5HSz1dwikV996M7aFbWsJ5UKyhRcOrta
5B2GROUDmPy9QCT8W1fctGNZGbH5cT/pkEL0PJWgtgQN7/ZBXdDWxuf36g95
pKoztu9citKXJ4RNjn2BVNVotCH+o5wKHSxHP/OtcnVXBdK/C0sGNj+mhjqj
3KK5oX59STXdhBF92dgRjRZ2wQHDnaQ1jHkuz4AZxZqh7TnL5CvyL1fC1uaG
bgfy9i3w7P/zvef1Ml1g6Cfu3yeQSoZ8dZjA+ksDKQdmjyVHMuwfjZZecg+i
wB/cofJX/SyYUCrBPljpf1BEzQ3RSfBcGG5VwHm5lvNsCQN9RQ+dSxA/uhs7
FNJ9aYlfvOLEYLmZMfO8DN4y8hV01kggTcxH0N4CuvySbCFfX1LEJyKpwcEm
/NuDPtm4mlR8GZW0f9I8mbiE5IgWw7Hhj2wYfq+w3QosDKGC6i+O+iSaW/ik
6ytx+K7gLGZSiri0YDeqexkyWRqh2KRBY0MBPqClwoydZ1zqlfv453xm9lHv
bCm/unAtfpFSa1hQlSn1dvVfmRVLTmr7uSTLar/RlSk2aO4vCrieQjMC8d3A
FscPkxInyO7Sxgh0QHj+EnUNMWYJgvQAUknGSvhDceLuJLZqXUGEWKSmLaw8
w2WRNdgW4bcWspOcJmHtl2pyZctXt2RJXWHBPQhq1cYZJbEVpX+jZeq+kaRD
DPQVP1q2fHYS9YJt5A+qYlGXbYqru0Hj32NCrb28tfZi4M+GqAxDJjOG+Rct
5O44e7uVz4gAkpdWqXRjR1o3a43VWWbLlfDKK8QCBHTnkWR8hVZF3hvuHgEq
yU1Rs57KWuBHTAKhCdkb+NYUJK3F4WbqvWOOPqD1pXvcHBEIQ9NxC2i8TbH1
2rUl+4ygnJh86xFnsGaCiSnPj2AsqrzJYFf5NcB2R1B3cfyw0xpRMTbxUFpj
CE07aTYjl6U3WAdkBPHINkmSWqo3TyvD1nkoAfKcd4Ep0pF4UaNxI7oet9PR
NQeW0H0g4WrV9JqFXlo546Xfy5HiD0PMQ6WYkO9w/qFcdq3uLJe2INtlQly+
sfjm47yDxTMBZrx6ZabkmSwr07093rXvhZKTq6+LjYVbisGqY72mVuRA0x0W
FJ3H2dTirduy4h81nE2o73bSa3juDB9f0IqBchiBDb/VgZXDTlUhnVJTderH
AxUR4MjSgpuXtXUjAQWFXDhF6iYMPoqXNLMTpMFvk0dC81SxlbQuP+kxUWzR
c01MlWJbgM8kADI4cQaDYfDrLoDVgy60tc1GL7stpRszuNCRTvq31q2VaU9u
Gv+xwLtaUWubF/oGkxtkH8irW/8IsDlse60jXQzo//sgWc1JQwGT+p5R5EWo
DM/XP5pbF53KfeTBCQDBx7tF69VrssJKt1IWtbM1X77TiNpO8BqYBiAXeC4a
9NUkfMEhca5Qm1GJgF3pSb8aQu11JC8bqcssGCqZP4n9+wEa/OVXq578GD7b
HknlEVizxygOkoNzCiQmqQPqChFnKDJfZ/3o0Q0Q1ufT+jF6+TxavqB9tZhj
K5EVDkpu6pP8KiiiA/y8iQqn4HhKvrMHglyRpiKwF40tUt0Z1aH0TFYF/hJ9
l1cM8CetwCMtpCITq29CzpXJMg67cm7qkm/Tlb4g9gS/Ps4PDEH3vjFDgh1D
Es5I/7IfZUjnAO+IFxgDQ+9WfZECpPoXXIGe0dx/VwaaMp4FPHU+ESF/DEDU
68J3Jgx0M8iOISNe+75E+u/g1enoHRHhlGoxXNahzUPCbE2UnIFDEX2SsPoe
RQLaa4IsDeIGIaRDAlnpyQLCiyQVj5eERC5fNTkrpkixyDUocPh4V5MF5KCt
wCf3BlYA5SmZc2rk9kdS0XyTHWwiWZSr9AfFd+K3YvAHERp5bMdrDUYS8n32
hsqdgdE/Wqt8iev//nNkSVBvUUyP5YegXpYhofrRslbNAeOP5a0kXaGu+LjJ
mjQlsBKSvhSPrJr1JCh+xn/t5TNkqnqYAx1igznI6XLBniai/2qFXNSAFTLM
jD77vv/R/JwksTwOCaGH2Y1A2G3HyK/eZBiRrwofXxvW+8SWVAxiVoeQv9Pm
SFPuU6gu+qgvBgl0enN651U9hcukeI0YMfLGs6J86sC/pcc8HvQQCGHwh8tl
wBUmizGHV5kAVKYmK94/batlAVFDmYyy/DaCftgzRenMYP++sbpCKsUUovu7
pmWF084IrZPVHxzKrRcdAB2o1KIcEwVwoSyxNZlqmck4FC9eYe+OWxTWBYRY
ROJLGNet2o+WMbMSvwQpIwQuhEIXC+akqRv029KKLU6I/+F4UDM1O17RHdyh
O5rQ9eWXd0iv5vY3vIkzBHSy5cUrHMdeS0J80kqfcNkoq/Mg5rqtiyvi14Ex
XwhF9ZxDslyLmNTaTVx1kQAEWjtHi6MYx9SVt8CGlBpSSgy37nBVyN0KI9vc
kiNXKiGMqUpkonBQnjC7A4GZU4JpQk0fAG5xKYpRQcAKYld61Yqpt2iAJhOQ
AzfLePtBnD+RTuEAYMFf3hOsL5oQLkjspC0FIlnuTnRGyi4FSLlpAbWIFfCL
5Py8Mc22c+lUq94hO58X8LqPDY5HjdR4MsAPqusropLbExKEnKDku98zFyJ9
Kw80OK1vgn3wpV/BWgarVkXJVBKC7qmguVJXaIBXX6H4F6qsR9fr4piNYgtH
DlCdWu2sS7v9qwAzTOaAimG7uoRqTT0ggFVbIXU1WBbH1jJnfACLeGXftVxN
DJ5fs98Yt/AgmCgCyN5u/knC/d9Cgl5FPka4gGQ5y9UCd+xgbg7dYLgvBZgM
17h3XcNmJDMdPyiA8HF73DJ5ckgZ/4yreBE6MGTGjDhe1DVVb2aHUNwaBlkh
750Pw/9DO34p74z/8lTnSyf7u2Dh8gl7/ChA10IPlEnhPTbBnQjYHJ2uJvCn
X887YC1qIkszSsu6pLI+N1sO7dVEpxp6Lq3aVS8GI6MjnnjulnYGK93QTAu8
FHcgdJ3upBIo5uwelQQnrahpIMM6euGQsBXmAxyEfdgYUE3VWO13rRbTeaD/
SSHZyfhcWZTsTNIB4+ED4FCe2psBk1uTbXkeYQfXUo+jtCyAMimc7OtCn+hx
1prW87UQ6vj6Rra2K9KUGg+RxWW/8vP/DQj/tHl0gErjwL1pwrf1FlMAnKot
J3ZTPnZ74ERdJCzmN4wjlU8be0e/gzFIDNGtwlwiCscHuKGGPSSPNVyTHcX4
DqdpOL2Y6iJb7cVucYnNzEesjKIy/pHh2XHdrQfCP4AaUPYQYxzM7zR6e46l
CN/IowTjduMGrx1xeawgR303WK4R8u3NJkBd/zHSnaVI2+hf4kEHGWYhju3f
ATKCBiWqbC+rXE8HeJMU8SlHp780TEGZOSOV2L08xC25IPcw0dyX+eHk8Kz3
NoFUq3+6tSGZ6y99bUXuR03L7okUHjcvE/Am3U2YCoxvAC2pTcoVQ92XSaPH
5GZQLFL40mBMFw8AXU52IqjJDTo0Czj4JekfJk/0iQvXoxMq1ParzbTzcWMW
Z5P80GcV/AMfbKZhN3oxqSuRAfQLDSt9k/LyrpgQMA6Lxdg3aB5xdHbnGrhc
tFr0IdUDLlT53nYXGv5pUxXNwUCIwTOuMf0Jzte6V+R6XVPFSq1NDRJY3aCm
1jIctdsh5qWeOgnk2b8BcW8DJVh9+Vcc9gMP/0YkCNqBRhy5h4r/+syUpcLt
03iibE+NkI++c08O0c+5X85cjmqw9ZLTvfqFX2jZxUQwgGOG/NQNrbF9gYo4
Cd2FtkdqdUBdFZNGTg9lBWsy99aHrqOjp1EZlZzY4mrmSmQWr8ouVUuzT6y3
7eK43P3n0pCi7SfyhHTxZjgELlc9Tmc0J6Y4ImiafZG8FR1ono20nbZzsDtI
d2PlKgawIF2xSdBFIGFEUCmuTz7Nseod5qYvfXRVjL+U0uYdS8nn+QLGBalo
H4hcSOIQC1MKOhdZpeCxta03zg2RJAm49nQLuQeC4bAaBRVOkSA/BmWjuOzj
o3WWWd7oxo6g1MZbiXzjYZgJ1REkZ7Bh1XgRR8igY1h6jymRVDqruKZETBxH
rO8daVilBj4tsOqXshAZnegAB6ohjX8v1gNJyER5l6vyvljLRRftiPAXVhja
FoAY0lXHcee6SrW3uKY7zluRpAN0FXBV0Rydqdf1WvCPkeqwoKhGeis2T50e
FoiNiEYkuGvLCPa9CTXvNOEnuDQoje72sGYhQ+k1eYgaKy037JnCMlgNtAkx
MnlRanwPLslSwJGtOYUoxmbn/nThjec0lZ8fwT1TZek9VdqJ51ug4OVV34i0
Q+aMCYuhOygTHuMq+RPdXx/fduS20QjSs7AbYQ/ldkt16+rI4ftQG64DPb4p
JzwPDOsYVantu8Tob0U6A/fo4LqBUVGkW12cj/Eo2U0cc96JeqGBCmFeomkC
MbA1/a4bYPNEPSD2/X/CQlf02Qxc9eyNalf8iZL3LB9vc8WVuORKz3b7jRJG
zIBAvnX0RAq1aXc6qfrRWz/W0LZNQWoaaVD8iIPboGjFHZlRqqLI0gAW3JNp
fMqP4PPKCb6GG+z+d94N/PEapf0vJlFNwhzjtjAj0Nam4l4rMi+K3lDvgIgE
f70T1k09QX4pBcoodWWcEJPvVBsv7DaqIG5pgDYhsDHl7aCAJvPrvRVYZKNG
Kchsj7bLoe1Xzkanlim9HrOk5WyUjATlb13ABI1Ufsbt9mB5R+6Tfd5VvXrW
zH1XpotKQVR6PmkrP4WoR/nmywNImy0o8ZuFEhj3LraFZlgoMwSRpGWoHUj4
HIMB7vVkcAnFEjiHPwKm5Kd49Wk+26OajYqgQG0eMr98ei0v/oBkIs/AGwdn
uoKQ/kIM5RGSlgULlvM4AJprueas97WWZFuhgOJwHPAlOzWGCZyXiPO6bwDL
ZLQk3k+MS09w/B4XIIPhKdffj1EFkS5K6AQruqc5w1kV35vF8bvQJrxv9Ryk
aMIoPlJpeoyC25YWwYcA7WayJKq0szeole0Pm8TaWp/98WUd4egZf/Ur6udf
+tAZ80TMk9ALbJDm692Ila3+lO8L3njQehpBr/918KWPV1+Pq0Ws7UxCH5FX
X8c97k2MAn5Oz8Ll1a29hpq7e3K55dXNUfXy2sbH4q2XR0FNNss1QUCOocgY
iCLjUdXo4P9RZu2STs3a0xO7ExvexrFi95xCXLPqPefIvAO+3evEZ3xg6wJt
HD55SraKy2XvKWn3IqhQnYeW/p60VEpPYK6tgIoGIFc4Lo9yWRoN+wqzZrj5
Sn/ou+Aq4hMcjflPLccV4gaJDL8rEKdnjIp6T6VGGg9nKrs32aHfkDN2uFqJ
VZTYnJatlRfErG02xxks/+J/rFyugpMfOBykj4FsRem2A4EYZFi6962koiXW
uMOPqRVEc4AwHp3X/8ZrDBgbkwChM939A/O/vFjxNXbZKnz3os30d/q8D3+d
415qKvo/nnrLW7IK8p3gCuT2CT2yVhJReeKZ9URZLfsZY33tdULjPLq5Ra1X
JSRjyPFSzHgQM/Hvetqfo+U6GR9J1Z8g5hgAzyzlGd18dWfQ1cXKsJVijasm
gjV3nXZN/aBPzO4AeV8nBlDrFtx8sMHSfGDOmLnx37Qf8v3hu6pVd0Kpyrf9
wzk6vUdrKjJqFEC5JijEkemErC+TBh+8lKgqvb0oI1D7CzTQkaYIz5RBmi54
sA54Mv6Q+G2rQ45Wu3rqmWO1v2BPCIXopoJG8QyT4ScPVCX/F+vo2gjIEsZ1
6kC0pHpLF72hAAqgbNgoK1rmABBYcGKzlbWX+apM0cD8StDZMz0/NS1Mzqrb
1PQPWIaDyazOJN3NoNZuQ42Rskk5N5a4jQOOL+zEv+IcSw/TSpIIesHZeMcd
xgoWTABnLKp2Qj+LjUeD9CLR0C2/KoafEC5vAGY9UoSPfAZXIJJXCVrKjOFc
t9NECjk2dZg9lemo3/lUZQDW9Mxx+LvY4x2EvYaFUFxkRNc9Sy4IXLbMv6aQ
jvB+Aro4ixoCcYFW6VENHdyRvsmPa5qThyIhGln6aUhBxJRC6xeCG1rEVIWj
HFtwV998A6gflTC7QJoU7RbdPJc463aMxH0uUjwwEJNWbm8qqGnIvj4sxwqc
aWVM0H/5KHgp8NrzlnZKjB1W8tkrxL1dHToxisbsvnbyshnbw0FcIoB/h2fD
7g85SQEOU3MZeJYU+bf8OSdT735RrshLd8Aanuq3PG63bnVUN1+LzwcQ7CXl
PCjSZ7JTrjjanGsbJIR8ZGcufFnI7gSXKTjtg2cmdiy/vBdxthjq7uBGLqyP
lrNeyFzoYg53EUGBtvqcHdm9Fof16hUWeJwMBYXND7EgJEHwA43MpHbxsZDk
HIX9DIVaM83JKiE77nXH9flInlZIcEP5DLUTwxdnl1yz/Xbs4hBiH2zZ8xBZ
5gum4Tc6eZPsAk0axsko8J7I8snJWqv1M2W39NRrgUCNNiTRpkrpPAhPCCDJ
EaJDgI21vUNENdiWdLhz4btt+3i+LcN6np8yv5osJuU76exf/2NKiU6id1sL
GMpnwjGCgohngGEM3MkUfyNuAs+DVIY+CNcGbLgnAiMx5UVK/wdSvaNw/7WP
yMh9yXWGjlrb6ENQQcsZPRJJEP0nvQ4jBaKfHuPeTnecMokyWlG+GSp0U060
7oUWQz3CfL0VD52o2BPHEVkEG26GzJXPelAGQ4dVC0dNz0qdkBmK52saFmi6
eZvoG+qoGXhdVVuFOO6TatZm5I/eM0fNgM9+Djxlor5EnuEQWjjHVX6rcl/2
z9qN5SFivHOKlgZGeu3kI4NxHCYdkYkq1A2ob7jrSuFztJ3D6ndId6HoK76Q
8b6byHc707JedYdzaKpgGey9VP2ft234V2JRYwfjEtQxQ9GWgt9uJ9k5lPNL
5moHgqtHlBs20bL/M8CquANpj7dG8tFWTSyB+WdZlJ4ekpxfQZ8yiD1zSjet
pKkwt0TwZNxr8bChg2Bk4MzOG/Imvwn+hksbe0NM0Y5wqIJhKRp+qez/DWZe
z8nP6e/atkumRVV8h7vhVJhS3MfqSUr2QBzcuVPkoGUjmaNWoGSGVyZheylT
Eh0j7AQ9GwKimhXOPVBWOpllRCS5HOANGbZXPv7CwB3nKbb5XKhu3bHMFeEF
OMw6I1Nehgd9Ib6AhDLQcAZqpCXSXCtUrYcN/QYpfvrojT6TDnMRnn/EDyWW
01nkYdovLFx3WIqferlcKFXlfZ+QbZAvcFaCV8zuHWm3Up/Ab5gOcsPnGt6K
nAorDjkH9Gd7xvuCLqF+1fbABbh0Kv/mpIFQQGn273DIX3VygHQPwp0Giu3c
sU43QpLul7qZ2jxDxRu4w8wuuU+51/HSDMAlEto3+LTN/+MSHOdYXWwHxw17
yhgUutJf6o4bI3tVWrdEFGqZq9AUxGXHC6g+zFBGcZUfgiPxHgU/7D270JzG
5j32LGbRnhvu5YQ5nIL1f8E7h5cKAwBXL+TG6NPNlfvS2MLjZ7mUdiRmHUSa
UFyNNVdZUBm16vYVTcXpIj/c9+MQpSkteqqiI33lMjxWIpCFwMs5MZyNorrb
+Ak7WCHicXZmfGpv3spLI9xnwMLNwEzEVexUbR9lLyOojwHgjZoaNw+qrRwM
JyczuYkIPu3Voz0fGuPreQNmp7gQA7pThtnv+KgLActW7y4oqWYj7QqE6a8c
YcIsrQ7YW3ajaW+hOVqhI8XY9qU8SyQTaOPyT/WleCW4D3YFESV7aE2CTUYY
SsxBQoGYSI2rlbcSWoBhKuXuDtWxmZLCZ3TFzRjSJJ5wkRkiLmXNmnLTuDAh
QEGnSUixE8nuddnh6b+bgpSijaIbhheBYvviF5oYPI60zm/hZOPn7DcQUMMN
KhBtf4tFyYBKU2gV4CY0HbIrtvXt3mlWkhy0MK8+5egFSS62SFoxs6E/P6Oq
58sibSTQMPulx47UdJwOvvvj1aNWDuImfG5FRfGn1q2SSd469ysRhqceLpxW
R4oSEz826bDXWiwmCZu765NbJwxEX/59og6UiIHqgXXsE5q/m/vtguuYaIMi
71/lQolOC8KE4iwxclgHc6Uora8QiOGqwbTLx5yrEBjm7h0Y47kmqIXcP7Ym
jBUHpc3heLTBez2ZvMxE3BQ5sS0PUI81O4kNCcbsL+RgITrA14ssCa+97/WS
8tdU9tYQNIUwCcvdt8gQaNJ1pFfT2FGJ9c7cGKUt8XzUKytYKC6xgkVeNl1c
pgi6UYHjzgbvxdNtQY2VTOgA2lGxD+6utB0yJ65t6S3V8kdEFLxj2gY9Ue/3
/mvC2YKE61hWVITu9y3/HjWCCWL7Sm8s1IMLetP+nsfcJ1MpRZqf+NVJwxLY
C6BAM/vzGGPceOTYaouRC59aDpnOlb3mqMnLTlE9IFAkh8eQI26nWfrkVfhb
e00SRT1oBMWdLp1RAXE25LdKM8L77M2fdYpt42ZFnbxmXvfYPE6sHPUtvXE5
9UZm/g3RfiCep52MDBIF40sOo8hXxDScKInwH9L+ETKIL5Y3b2Za6S+Qkicl
XiuJqEBzE5rEcPTY2qMOFMfSZFn0clsspWs0eDnx9z4shv2sA1s4f28kyo7D
pq3/zA4tJPoNQRWhB87tyQ5yRIeJoHpgiQKaJ6d18obNVlesGcaoRj4LMYjO
4P5W5AR56UR/1jm8TFz0r6repf2PCCs6Q6putzvxgw0WICPj/8sB5H6ugVA1
rml9mxwLKcpcR4y5ZyRuKlWM0O8xfBucVRv+l3yiImnLY/EGKMwEYMCX50e4
y/uKDRTIcfFy0Q4wyPFMm2grESWYnpfGARMm4kcfJirybuKJG6FuoXsE5Is1
C6UK3fObjKVxqKmcrr8VTVQjtCNTPoa/ffvdyFD2HoHyqzco6QZTEne/2oyi
I8R7jEuD2MY3JFBJrXHrILOwJDEI2wwY+YH7uoejGmx/oHAJftTk21m5fHJV
go/62ia9QlGMASS/evW8bvBJB26MdoogC5zfuL3NV5LR/UE2A2nj81CnBqOI
xn3JLExVLlmY4UejgvxD5BUjK9aOXoj3YMVppOfhglbX4AjWhgh+vuUCmBsR
0XwQoE2YQkukeK9Df5Sr2j7Z3JS2NEIycMfKYag9yktyaszPjOvycjPpUNLU
82yRkUtLrUQ91FbP7KmAGQpvPM3q7S0UYa3ivVxiypKUBUXASwR2RWZnAEzl
OZn43A4UXHBBNJTtlGEvkrJneAtNRro/ii2BJWJKm0+uIdH5jat6Wb8d4oZv
7REzGYSUZK4PO5C+GQ8ABOlaLZMjLSQ81y6nfsxE3hN8AEngftBNz52D5VuP
ZslSzmBOC43upf6+S0Nx/p+CeeK4hb+TBWMHTeaAouvhUcZy+9QiUJiCljtE
pAbrZYrZ0adfSoZ5Q2GiIdyLRHjCkro4ClCdtC2+Rpd7kBUhuqv8jK7zBZU3
wu9fwKxvaojf/FhkvXiPEwv8gjTkLIgrT/yejfrXpw+Yqovp3a2YzQkTjxw9
T4DIIyzF88SwJvaO2UbR1RKQVY4fS7gQr4Tr/q6Ti7YV+yvYkXVBz5NCRupd
qkHbgt0JwSLZJ8EecjYuF//1Akw9X+/36DhC3wiBoYIqhIN9XfQ3n8NP7A9D
OAydjhT+o4jGlnrlKmMcdxvKeCq/eN8OJSK+lRpjQlxRIbw9aeCUDYCGFdu4
i2da0NlViyLaSc9nTCl0tOTit2GsqwiyClsJxhdeE3Omcm+3+XbkDzsmaaEz
FzBZkQ0/wZVHyhQFkMwrbn2QUikrdRarJkda5CYUdcj+P6KpNx62TIwNcG7j
yzgZwbga8iFNb3/z6c1TVgw0j0ifrO95SDjpSnC18aSlfQBgtOcKpczEtVcQ
SVe5QwxCYEwbSPO/nki7xS5lHAHZbptUIpH1yKzpVHHqkvq4j+3ReVUc90KO
KMkue8rCZ34XfRDDAiBETEAfPSMDRHWECtJsoXyypBqRfNq54Fu1Amv2gCxW
fA92Yo1BXzpSDjjhH7J8KLZqgbfYZzcy222ii95l35KErpmQfkT0sZK70EIm
s93PlxOxPxthKo1JTTQBJPEOai1gEaEovAzyD1FUqEDzVTDHASlUhYjxVJEJ
rKM6xwkTTLJsgLzISrtWTc2gK4WsX3lPR227H8OJvhFvB0wJVD0GjHuS5TWu
MJYeC+RhZttHMeXqT/n9Bz23iY7vwp4BaZYw4lE0m3ipD3FWLEsf/SvB7lkY
+aS26QTrbD9pcnVsNq+BoJSc3PO9TulNOb/xbJC4VUMQEyX2otDkulRL+Z8P
YJPEJwEMZ3E04cC9wXXG/UzPwP5m3THL2rUBTeM1I2qtkWDXIEerpc2uyYiw
uYfIeeWJLBnsTwg9uqhzladeDKCu5koWqMK6wVk70136M1omev7gCS73AGyM
tuFCWLXEH5q/dYOB7Dag+zU38nwljGXuPydZQMvKpV4UWvyIDZJqD+KY7uaL
D3XLg/x7NPkWoPlPTx6IdKYMceULi/W3WxvNSN+1V9En/XSF4NXyKGmNVhOj
R8p/Fc8YXQhMqiOOZiZSnIpDRBt+UfVFJ6S7IdboqmqPY52ZIwsyOFxY43wJ
5mBWvHqLz3CMx6M1r56lakDetso6dtiiLgNrSsCLRqN7GSylKAcLdxn1XGQ6
bipvUhudS8emqEevu2UU2TCd7/eadiJjuNXX5oRLIJKY+gOucVu8GccnfSk/
MYNB1GcXAivi9BXCWh87mgN4sgj8C9qSaAL+tkxOHnZA+DUXZu6yv2ym0y1b
LYCTiXSR652OslK/tnv42Z68mUR/AyMb/BdaYJMxVFSQu0lxLjnaJUxyfi/s
knxBA8FwZVngw3nERxitCcuudRoga8810WwJfSSWiaYEmmct9fFzipp+9Y0c
GcpfUwZ553UZG4WTaKaEbjRJvhLYvFliRecUznyc7cj/d86fA7ZoNLHtLOsY
SLI6jEq+jJs11wPLUYeuBlveeZTD3K2PpOvse52SooJv9AlX2voXgYH6EEo/
aBMz16Fh09nvAlSnaYB6n8/wQi0UaJDvux+rBYAmtMw0JoLTQfuuK7qItlND
PJbEiXzCNDwKTEFv01JB48xIwEQbMctE5jD8PtnGHOZDQ5sT0H8wdIyP8Ggj
ZxFbxVFpSFrakTvgWJOCOdpnwYTkX7p11JHco1MdZHygFW/55A86F5CCW8Ml
RV6NIB2L2FE5oijPKfdG7nX4fChg8+9PO6IO8hIO4eeIrT3/uiWm9Q5L9zBc
TFe2z4PzCy+HaiUIw7nlIF2xXIdPAK7Ne5T8z+o3+5eOZcaY12stybKc+fve
I0orKpo83WlkufYSqnopuv/eu9jF82cZT1Joo/nApMJL1gaObhDc1KC4ESgh
y7XtNBDzVY8uvy4YaAV8GsEuSpFDXdQ7sKEwYV1a2KsPGkZGP4rfvzRdEPyi
sXU6IFtzfJnRNzSgUF4jiQYVSyb54oazfyB/GEg43XPTjpaRtwvIgFL+HiRA
oWPznUSW1sX9EWr9108EnAnOGKeMotJSUM71GMFUlm6rnTDW6ccgw/z4ns34
YKbIxJYd6qGCnKlpeYiVHS+rRA3fUtfSbDXuiAp9DxbJHJCmQRcF7OTsudKS
wbFkhXqP1L8FgCMT34WiEBBr/sPvWCwBdqmPbpeXEHI30Ixk4/cEVeHICCEn
jEwYBUhrLzoXXpKmwkOgpQulIOT+/Q/85gmxIVtMrHP84/+HNUnj/OrSBrGE
mnTy/9V6U35aeicS7ih4avXDnI8tarANlN049ReCnES+phw0J1IWlpBu80wW
mqpm2jdSRivKCasyP2LuAVOPs2j825OjlY0fLtrT+ChC87x8qqN/ZDUfzBqh
lqT8lAYXUofc/SOjvy1zR9EpK9cLccFqKOAJciuJe6x4RwSmwZRE6hzWNATG
ZZXnkhT+S6dMVLDeB/BGwoBrvPre+4ioT1/FcId5YM5ExofXFIZjFDGLAi22
DH7OPVtpZ7oG10K6gEfEWYEcsHyFFiJUDXqHLNL84pCnkcpY68+Ti74tgAPi
q8w2AWOQe5fbqhh5rvv3E48PuO63zYrP7WKf1coMQXgHm+bdmVM4hb+RoiJc
8ZmrwAxbEA2m0zgynDGH+vB10A/+AWqGCGeYocVFbsSd7fquStnQn+aph+pP
6WaRsk/FvFhzQB0CoW+LUawgzx3HvfVVATTEu/WhcLkYxYwLT0jPmSzIz7JC
kFUkpiq1BWBvDlzDKPLfj/EpLvoK7/usnALbhLku+yPPznOsrQ/5zdZT0bMo
MqQ6OB/FOG4pclPdZSEQAd5wq5x7bNZWidXLFBZo6pbC/dcoKMvULgaB9et0
wf9Aqm96CVILJkcnGzKwaFF3x3RkQXroGHSU6qLarqulMbXvG75o571P+L03
U19W209SIMSvHJEHjF8j8uJ7BNSzBN5pmn4QiMdMuKNFfM4DL/L7xJtXfU7t
gOyw3umdb1kSkLaKsoi47XJ0jmM/eiVLmpD+gojWnIUjPkmW6CZsK8SmepAR
pbm1jL8MNJrzlWPd+PmXY19k4IZ9XKUx2+RLfEyPJeSmcxTFhTIgmD8dA4Du
PZl8O/YeSuEUyiHyyb7i6NAhgPStQpzwgDeBdeiNZuIPnxPVNGOGFouGqEkQ
0VwmFiLqwqacjTjkYdNEFVaUZVXZu/meMzaqJF/UZU87UIrbYzuQiU1eIEwm
SuYTr4aCPUAppMFw6vCS/udUm1MjouhneuDeJv2ERqd/wIJLG1FWYaD0AilS
xVauEBWsZnmYJ4QHgbCevLnqyt5mCRqWxCEOljntlNlIwIqLQGk5qyd4id2s
JFt/AjK0BePcN1ph46e1Tn0raEuegUep/mWodOBbN0tP1/NBAw1/vIl5HAQ8
24iSXDtDqZ3qNKXQ+lglqQvAAvsasw/PE1Cv40k0vgXpzB4y2Zd/ZwGbuQIQ
5MN369EDgRrkAkSkfY291kqm2KXZZ8TpF7woNjKfzFUIwi3qPFOkjOTC7HZZ
2gxauNKSUhD56w8zudPp5A0d6We7qC3EYpaY2SXdCb4DUnqdeL86TZtxo3jI
ocKEgTzyHL5LAi9mzy6QwLg1D8vVMRzyMaxTYSez8Sr/vgDb6ahKi316E6Ie
ZtMzddc74mApApdi2OBBWcp0Qas8G9jOcV2+7YmmezwE97870/hN6n/9vhkx
5ZrxDjtVvq++AChWsKWVlTkysUiAMJm9SljNOwLhK0l6vS2k7IeLwabQv3S3
+z6+YuuwJcpvELJiNPFJSJJxUcEqJ+vXlwmKTAtXOLRdT1hDfPQdLF5y6bAn
We5XJhsRTu+g4zaafg9lgtWKlwIij8dsytDi38NX+yZpQWt15QxnP6kNJ+HH
UOrBEIwnZ48yBRl7TSobXpqCt4qv+ZTnQ7nAoB3HdSU+0ysCTKULzsUCJEpK
WvS0ULyXK21j7OO0RbhLgjAZVyFEsM06Y3S4rLgcCYg4Jz8nLkNLAzYUVfBZ
XmC+Gryfppg2T/3mgDlmPG77Dl9iV/k0qF/bA0OtoggjOqEBXZ+3nNf36SEQ
u+Bm3/L9QZnUXiS/wfqV9KUKQ3BEYdKkIN52NaIQP4pV4yJsARgp36hbrOXm
9NiXS+cxmJdnIjbgOadZNoXfAjj9oFsGkCOATp0wQk/DHJBpfHB5s2oACXMS
79Zw1FQFPXNkfYWInAMGth0tzdpTgv0+r/uJdhBOrnHXclp1mjNPFfZfGdVJ
uUv690ZSPg6YsgnOk/Vpj/OBIdprUIUrSPlWbS2TuugJhZ3eLaBs9kljO6VW
aS3BaY4GXc7KIKSqX88m8PiAfIuIhiga+rRYOhXAwOkHWoF5TKJRMZgkCPQm
/9biY3YkW1IHFg9Ggy7rdtcXfBS/U28FZN0gYniMNA4B3fnTN8NqY8j9+KLK
nOs/p/xpZ/6yqAbpOMgSc9lazHgmuRhoVkgNKufq8nsUG4EAFMWZF8yxlHxR
ULdXDUU8ofCvQr1vJiGvkMBD+OMXJEmItpIHLsAO5KEo3egT8y9qoHNZ30n7
5mvuVB38zIJ0v6EqGHZpD6jUa+hCyNe41Z5sXFBeFcdnE1nyDRIrYbtBMJSd
AhH1Tz5/K9tHZMCqZOBbl+mbrnbvIFvnvme83Y5705Bz/jzjdrjfAU0WZ6l9
ELa5XsWRrkUIfu+cqKMEdGNcPFK8D3AXMZdWjyK3Err7W1M0W9fJjZhViZSh
6yWO7yIIIzGCtKnHvxJ6c1zZomctroPA26gafqX5V+VXixdpkQuR4hS/2ZAr
9eQZXoHMfhjFw3E2j/pAlOxdfLFQQnS/BPH+mb0MCBa44a0rYKVIZYUSkJti
2Vhi3u0l0lpAEen/higSZ5OdhBsecYkI7RNx3dCABEwoOLcA1eaEP1oGCZaH
MwujYU5RS4ZU1T+9m6tIrtpAr/Lp/oHwWqr5k+TCBIUwKNte+77z3NrwIReW
gwyjtyqbYTy/f7qr4eB3xc4PvYusGdK+5y3/CedYj1E0ZJM3VFkYKjbyuse2
RF5osLKL/5FL8+o+AjIWGSbLPdryPnrO1kjdXqQZI+I67WOrRCvPDez6Zq+2
xqa29PpoZtPf63pS4DXEvOAaEeoNLnPWv04BI4fAMtoLik2myTfA2AYi2yUv
JC+E2hORGbOLILA1FN+Qyy/3+kz8w0fFeZEiFCpzi1eH3vS8kMvbyXbnzU+u
pS0RsTHFqb3j+Hbvl4HFMRbw3SG00rJDaZOP3Zcpjj/TFuGbFfSOaD5hbGen
fc0bmER2NgF6QzRicz2teHFEXGRR3Yu6+mo3BuRLP/MmZlesESyT4aR1Rzw4
n+rkdNluR9PPH86iYgFTVNB9pwyS3Fix6ShqC8sUvzq3mmWVqt1HZDnTmcs1
m5HAgzlx4GactsIOZbjKghN6Gzu3TYoFD/uladDoRbyFIPuaXJ7Jsgh0VEr8
t+P9MypCXCObB3pxAa1jymc+91eqtRw/qxLvi8oukkN8LEu+hZJToUR34b+Y
LGQe12bNABRhrJxl54Gm+cHfuxHExJ15epWBx27mtSQmwGyJtl5kXxqeshOj
o9OPxmkb5mL4RSbYK4/V9Lc61yV4qvjZBqOVkr1EiuJy71HxQhrdVJuiinTg
xddv/mtUn9vv7FR0rySo6JTVJe7lyFbXxI8Cr/xXkOLT1MOK9QICQwhmCSAk
dFLwrEhkjRpBb8Py6Rc64naqbpEjFrhS8xn+2ReVw6uKsMAH/zDF4YqLQXBw
2JYd7qouZAyz5jM0gYG7GdR6p1RJc9D4NLWoBhJlAJBe86i2hsQZz1g943Hw
deJ76UkCzszV2g2iuuR0fMKDh4V0BxrD8l8c+gbECM/jOrYZ6nDxDdhxdZlG
Zfkq0YEt5VcsjIGURoVSCRktEMD5wCe9DKe7eh6xVf2iWAdg3z9cIt0oXL18
6cyd1ryVdMsVYOQuOhSk8J9Ymm68o34oi/G8czZ0um0sA4QzOOvhNdE4oXNO
wpvKqOYADfNpD4ZRczdGLlrv6Wx1FqqSFb8hLuZAmXR2eFihFbNKNG8L3Iu1
3DupzZpkEcO5wKJi3gHGfmZinAX+zjIG/opZCLndNyj5RuQ1Z+YLe+7sQg1p
QrlRah5jQRb0shEiiDeK1mwrg/ElCmceTBbttlF8M50L+eO0QT8lo1J8Egvb
5jCvqzJ74d0+SsuK0Wwx3yNt/jOwem9mVu1ws4Si8vX4jCwKqdBGRn4bLs7x
RmI5tnY8aUbulekwrfNn3AghnFMXTMSz9qcokF+iq6FRko2oF59JXar9WzZQ
Fet9EkpWKhM3HtMi1SkbW/MAPiJf5T97d+pukTXJWws83ltRrb2luY7Vt1gz
qkf9LBeLFh8YaWWCcLPT/c9Xr7qXEeSrPFiOB2VUs+KC6If9Phl8jhVgmHm+
C3ljFE7brezkhTxUfy/LS57+jhC0NTid7kx9QxqdQws8KDzrr95ARZQweLoP
EMiNjb+J08+1Y62oP9MFDoDCc5L93UBAFe3V22Qso+YZhzmcLdSHPfeGGI4N
tVVqBIKdaB2zQn4VIu1FZt9und/wZ//izasxsVzg+3pEj6kBS08Z/JAsP4FC
eTojHKpWdQlw9+YppyzJB4QlhLdKOZ+cunNlhxIuIaHyqiR+Kodi1Ub75jZY
m3IBR9c7I+LvrgklQO1DCR9rCqzlXGQBX/mBZgl+ENzTOyI6nZl1fG/Ag1ib
j2+KWrSaWQEjbStxxC3znOYep0KPFc4/bB2S+1l8gXAmrLuhD30l5zd4bml2
WUTw9uIMOIqVtVxjIWi6FL6wxCdwxa+Ib4przLWoqRp3kLhfVTnGJWdWWbGx
nQnmsTHY01ShL3N+dovNT8bOc/C4UROR/dBsec02gw1q8oNOEVsvT4waDtMC
68ROTUIABi4ZwZ2/8B612xwnadCVNJPNTe7R+U4TDEF5TZf7eW+JFB4p/cV4
GSZuQHCJ67y+cB9XcadmETFgVQd3ZgV8O09BlkKJiBBFlx9JFXzGsF/agFvS
f3UKDqbZF52H4hNCAMhJgunV5bg4CdBeN+9uSUpuKa812FGDm185hZTOU8XK
zTEp3USQRYLEvfnoUFbQtUzT9ARjXK3PyvmnPQ4zilxlPbeWIzQ8cMKctqMY
ZJ3f5DSEFquQx7f0noYafR6o1TPS+eiIvziI7Uqs4kbpgrhcONRBNHlgtHPh
uieo06Lt14uC92T8mK9ecKy4cf63z/kED//Dh4DlXGUe2fWNXVRg3jQhNA6N
UGzF45H1MsXypxDk7NxdysXLNKyN2IsO54d0PsLRhm9vQpdRsxUP+GgND5j4
g54EzAVJJtR4iUzr8Eztv9n9k/NXJOzP2IneO3YeEkRoHlvpXzLDtYXdmzIo
SKMyOsis8Cr8rrcEu7Gj+kFD1UkoYm3v6K0wUAuDJ3GWg9/xqGGoYSF11AAV
vWdIgRwK5vq+6GYPKtMLZ8jXe8LjWqkOOvPF4ihiKjCFw5PJIdK055yb/Tlh
vGuxRb7oE7TZODxxfO5aKIV1SdD1Le6P3TZ6J2ZDcBKPpF/1+cuoN81Xcq5l
mXNdiZgkneXQgcorAXuZObd5ApHLxF9GGK9E8RvMn4AuB+lOGgMlYI7l7ab7
tZvk3r0vOYma4DzN+elcBXaAI0Oj7OUxWzNKKX9Hm9GNqWcgHKwRoUIZTIh4
i+XZVjLdnEmXIGZix1ZNztcODr+ATy9+/8du5GDFh3ruwOM/fM9rzCSrFGju
d5KRLUZVemE+syRjh72Dn/7kGGyPj4VN0nB/78eJyHENAz+hdCW93RTJlIZB
pEJXWcEDHI3eu14OJ13CGUVjwh8ljXMuinnpFyn38TGVu9ruknX3zl1V7lLg
XEjoohw4TtDhpZQE19ljaqrsMa3PJVLpVLGv6q7EXmTlsCjTEsgF7dKwIFZg
e0aLnU6WbfLKxLA84knRaR34BfSBL0NFgKg/GudB3nLZntah91AWuuabLj4F
BcSugzR36t30iD7KRydxp4rGYeSdWM0dO08wk0dPcDjLWNLh5o9IquGdXTD3
GP6ZRhbSNLlBh3T+qr7qEMTEXlKAUppU1NahPpqmmFDMMUzbBBgT7x7ueofS
dQDlo1HdKCQqAl4ZXXxGsg4/PZ2mKzZ7nvfqYbXS/VkLyLOKmzOXgAmAbKph
lasE6Ng9el8M4GdQ7C3caIRZG7v0VhFKBg6ndyzjDwY7Q1oFFfpF7d2/PdpW
ANkcYypxGDnlZPigt0WctFBLq3M51dJke/wLxh9eVb81oSfNv1mqxItOfph7
1CpQ7aQ1VjcTou5oN7n/hU6noegvO2sk25BNrGURCK35ZqoasLWSSs+BqTOC
Exhb2D5oqjgpVYt66sKACM1T4WA6p5h0VH7n8MAv/eWte3AahPXFm2dDd9vo
J5qXD84StKaW+XRFIT3WbUX2ikMuaTixpNNfetVimUeaua1qn+1lVeQ/ueZa
sbt+sNF8Y5q7ZmNEHbeBg1FPSjYKPixBQ3xFlzIjBu7+qoGlb5Tyv+BEhPgj
6eXVwXZuyLO/yp4xeJi4m2VK7W6n4Sz2wbhbIYclAW/RCd61USGr9NaMGMAN
b726us8OdLNwGXVqSy4KtnSlKnThfoUXPXk9JoDu6Gm5qi4es1KGBs/Nz2Lz
X9ijzEdsnlHpQh8hbLzLSZfYtrGERhZeIdqnzsJQAkQLOVk0TqzPFWpWQ2zT
xzGv2Lbx6M1wmtfENy7RdG+diV4GZjgD1zHLmAjHrzKvozFB5WZX/rOHuumQ
O6j3WUhiF56RIiJcjgxcMTIHzN4r49IXaajou29jxNDVFQDa8C0E3yiCUC+h
vHAvcQmViRo8kYUw6TTUXMh2ox4HlcmAMjxGKcUO7GpRC2Vpuxo0Guzpxlfs
jOWglEMfb3u5txuLqrLRTF2fYaniTNqLDccjkLM3vSok/vB2J3fvqtZBb398
j6MHZEeM7HxW4tTX8jQxI1C1kPlHwbJ2kG+4CEgo8adbMphRuhrrLEReMHSZ
AdEW/tdHCo/w5hoSCoxrNq7J02N7ASeym4O9c57xCFZ8q4e3CwHnmG6Z0EPg
tVElOzCuI8B+3G2iEhkDwMaHowZEiYz3HaWfYbPShCLZ9c9r0MWB7gCyXSaq
ECtPSfixXp5EkvYbsIGgsEyDIvr7ayZqo3pyIRThwDdFSlxRFR/milXPwDXo
Ppwi9OCRCITbLHwR5bS/otoV9Yjhp3mnNXH+gJGZQyymaU8dYFTxgPfJdYfi
Krptt4nDB1SQorRpSYo0UKjHUUJvYYtBW4RgpL+duPW00oxfuuXgrftJAZib
VBpMiEmQ8Nvod5ZmLrWG017KxDK+V03W4issLpUhmDqKle6kKikF4+0tM9PS
VBGHzJqiMQv8SxiGOAJjzSL0OitdIkIjwGAB+0kMxYzDC35ZvvczYEQ4cZ7I
bBMN75Vlfzh9XkC0q91lUZytAcPMzfGMmVVS/1sZhrgXM6sikJimJOwzfplg
JyYi3RoUL9DOJ33nNxua3sa8Y2BnjOdM8s4QfxbCa1fXcB3eDYri1SfnLPGs
IDzwC80msvUdUr+7pbqy0dUg04KMjDMWRtjXzh29ifMbBWC7uMnWl/U3X8IX
jjPFyW7t4aJ71q+2F/2GIFXLwlg2wwI615IPH7HXP+GjOmGMY93jsPcAU138
vwCMBVUBva60MqOnavSbWm6qombdDqG78ryPcXlu5ajOUUNKXGGXa9iQk+6D
W1j6nsNmb1XcaFFqoWgplafdVojER66V/A2i+aTtOvBbT1CBHO4kfSemAfp7
0MWNS/73OLs6wg4bV+NJOIOIEGWu18TTZmHZZHVxY1GZp3XuUEnjK8jh3x4A
SCptac6mcJ2HlXrm6dCbVvobsv8DHqfJoBvr9tyqDqq1FPvlezITZkeCmqaR
nBft5wSighUHs97W027FCx76b7MlkAIJUmKI9owXJyJ5N1au8sunxWPgA6n+
Spr9PwEDfNr9uNTcO2/cC98h4O7fwBEaD8zoHnQfqZETtfMA2b9Fbo8oYDGk
Y79lvowIjxcYaUjUxZrPiCaStM7e8IP1mLpZNlATlYT8WutyGYpdimCsVCFb
/gSGCrCCWw5f5Avom/YRIR6B/+BouWv5egY3ld3A/GJXdLc6CB5DTQrFNtY7
7wgg/gOH3nNZK2iwsOhQK7iqV/h0DjFfCKj0ZZr5apiGrTKiRs7eAAe1Tufm
9WeyZoovq2U732v/eU0qM5hocfJnD26RP0ZKJW3McmmgBHPy0e6pSKSiyce8
ZVvWy3dN6Lng+QuzdXhD+Hdy9eLU9LUDakI5rCFtDVYXCDqyCN8a3H0wLobD
60NiR7pR8vDGZRKdoR57sK1RoXrvPq7Bqiz3BHYdZkqcL9dO+YiZhyxmOAVZ
ofN/RA33J3mIhOlLXydT1wAKrPa8T5DQHNQC9vTYlySKV7ttrxKFsRg//6Ms
I6io15j2GdPkQQcA8JnQZVT2yq3M7SDGAcekLYucWO0GfM1/mUk+M4JMxXB0
Qb3hLkRafZLMAJfmn0xOAvyJn4XTKHRyYoHvUC5YD5dPO0FOZcDtRksmk7Va
i2A7Nd5heEsavkY8UuA5qD3+kMWu9sB7wtoq4KYBaEcfz1uIZOhX+XbuEYrO
ndqLW3lCq04f50zeZtgKK/aY8Kr70hUpAadi8QBC5FSmJluzCGU95TXjNK7b
DIhavmR997Wr4noU7vU6FNszR1Ho86gI78V7MrM9EJTaTk1QWcx0TFF4dh0Q
iJ5Y4DPnlmNgK8wMrWgVr2XsduH3YaGtBYPLN0ETavDyDIhVuyEVPnczcdrX
XgvSQQB724o3vveksL40lavaS9yT/Cs4+h4c9lFPx3tlfk2YsidB5h7C26Tc
dMpsj/5Mj86V/9wKqgrWMOpPTmrvA99fOuz2Em7SJzp5y87/Ri9ZBjePL+uX
PvtiOgswOvCiqAsNE7ts+O1mAzvQQ5iAM/XtlI0YyKtaaKFdj+SUMQPlIcoU
RVhm6D+Dalz639d3KHFC/0luOxc2Ii3wiimY8YNBOnGOK1Sfy9KcMm5RRVwm
hc8vZmPMQCFcPy+jPGKAYqgDDQUoYfF7Tx90TcS0L3xy2rMy0vopCzrzJWse
1W1zhSHEUx2peCGEYz87QqBX1A2ENhldlifwz3KYaShBqK9tvSA/GalFxIdt
KfNjyAZsO22jytWjWyyofWf21zN8XaD7Yo5OFso0xxeiPkmfkaVRvbZOCZO6
/kLDk2+wI4ykwmekIe+3BuO4mHtw1CVI8jH6QzJSNEgh1kXBq/trQ8gJS8HJ
hyWbpKVa/kiNv/UR9y1AEUrzbpt+ZngWzhU4IiS1EHC8cy1L+nUpk2inHqIo
2iW/AcoWb55ldHWMuht70NytZ7hFMmHYCTMjUCASbFV+XWf+l9ZOGczoacK3
9oxiSqpnGKg5XP/L4WR22S5S5iSW02eQI7FH8sVjnXWh5QdpyT3KPktc4ir+
JRZ39UAh0o1OqGWu2MmAZLzGcQYEfCTKBQZe3T1MSp6U5ucbdDhBf88/hOnA
SAgjHbQVmYFndPUpBPT77X6UFCzzN1Sz8rUAQcutYEuCRk6jVRwbn80CK77r
OiEk6dgVs6kX/1NBbPpQqYD715R0ha6sNzU1a7Yn6rjRmm7N/z2FWbvI3yw2
C7KF2Bu9yi6aTHkH8d4HihV8Xu7qHrNLiGBM5UfeNrz22/MmRJImkHNVms6P
GyT/yJ/E4KQQwg7aS5x5wayQOrDV/yeWTN5LSYf9i2TGqt0PCmxW7q/7ptXH
PVLZG1/o6ZUyuMyCqX+pZi5Ny0ySC0y24nIyTxMSqVZVNo+7PMPXSDR1Pirz
BX9NtKB1+qwoae4CbgtHWBqKbAe/GjSyt1Wu9k2sj078zfNfzL5Gj2xVlgf/
ElI37w45OmIiOCbtVe6Fo3zUkpCTbpNRri+tAoPNeb/rMwZAZrBe+yOP9HgE
auLUlF8+KabCYkGrUJ+MmvxxmBU/whH5ivbyj6vs//FM7VF1/QuOzWQdN0F1
9zvayrEWfrdRiofOrpRMb+1WclB4jWLU66vCzhQzGr20jru9R5F7Q+xlQlfu
G0XdZZT03JAHILCq+NRei/1FOnjXNNGEfGYXKyzBqB9OmUBsQnzIxQnkPztj
clMR9sD1yu7BG1yIzVucCQDe9T3D5o2BGjg7zzAnpWN78jhPRuQuURllSubQ
ToYTiLZjwxL0T0jO7cBLnb1DSY5wpIZpHB30spAz1/mxYxmQHrY54MryUoge
XxDUlINMUvupx9I3pa7j9BCf3YZPGiTKIZtCFJvT8uE7BRGnWC4KZiidK16o
7Iy6XGe5HLrd1yLLSP7aC+ZoG15F2dWaqtFloQ+I18qZQcl4GzdtkkvnoKlQ
HGoorp9pF6eg9CwRTAaPt4gT/DNLMRc2277eUMr/OGLSsN/mbCY50l8vTAJg
G/BLhnECcdHvGoo1hG32FdjDWyjI4Es2fp9kz3cWCOBRJ7KU06M7QgQXPAzs
GneyI8vYESvhCwnYiiphsfFWMr4oT459fOHg8phmCw/wP6AkmDQoNuZpDnsi
C8W3r3UmrWeGBWC7Zqq1QuHZF59VnjzJgao3wrgNpkdNup9HTWDPHPrZXr99
1zGKuS6ecpiOCG99IEoDfVzrBA9rZdgpKQ1BM1ddtd2Wybf67eNliNq2L4Ho
aiSmKgokct0css43lUMoxK33G9NDlnViJd3NQhY7hSwGeNTzgI5QZz2HVbUF
B42sLzDtNJx8FX9qnpnVME5L98pOCunJr32nN3DyC6Wy2iRnDL4JJ/JDPlYG
eV0KtrvVTivx3JINHhgR3hEzac7D5jIa6VLJsY4YgdD3NzZfVu0SkPrSDu43
pE++CB8Flm5JiWj/Uf2xwKTFO69dJAnOjsdhzw10QPeGUJ7S3BH2Prka2q5P
IHMZOtRsKpcMpTsa8rdn1YAD2T4gvHIJ1roSF3AvZ9cwbfc15Yn/jSWaBrHo
oDJWY5Orx7HAURTHT2kXoBhREkZrW1PpXCsY934wypkZCdYy8Fmjy8Qh8v5w
Cl1F+WSevx9IQfrvojFpDVu0uAuFsJz/tmTZx+bL/ISBLgsqpzj+oyVr6xY8
jaNXmKhDbb6iII3QeI5BvU8834QfqdFw7+0H23sFpQeCjftCRKstp3rfmy6K
OLKZNXDhkQ9lQ+OYSOxj0lidNVtBYqTzVCujpW0PwTAQk3nvNrX4UbZKQeUU
Qr18+wjjNGtGfpI9oTAckdBdbsYxT9prSFV+QcEXUjBpSzWeiZ6OvcnHRgFd
L1R9i34eqtHwlfZ3+YrecjfPO06+X+AYaOL6KpwJvRlMNhplbRGV630WpKWP
+mU3kTchp/JuStk7zAp5o9pGxJV/GlKTuA5TSyqyePDzgv/lmVUfYpN51m2N
MpzYupwrYVCb8BlwAw1vCyb9yRu0fIvNKFRlbTeVHC4Uw2+pi9wTn7BYIION
VjiD3GZqqvKOTsPpbA9o5w5QokSJ8fMQMCKo6JUzNlhmNu1A18mDRMyEqnNl
WbKaKHrasrtxJ6b8nhFz2NY8EeDkbre06b/D9Kj5tl+fjxyj0OfxoQ+6I/5W
5DZknpFfLmaT2DcEdmT5mdKeFVEKr3A0BuB8WSKtNVdrU6muRJHwx2D/X287
n9SpHsD+p4wriC4fkwL+kTpS+z3Rqi8Iv/siGiiMCh+Ps8O0TaPg9VdufDqt
4k/KzwJMCJ7MRioPYoIzK3MCbAhE5D33NvMZG6/29EUKY2K6r2vmhOYiNjbw
d3GFqtdB3tYE9ge9VDBihXje8J038+LP+T9R16R9Z6Hm8bgZHNkgH8jArbV9
93F3A/A+ICUEfCH/zz0RZDlbmqnaTuYkMupeBQVEJOd426glR7+1JY6zGMDC
US2eN21L+N2PrVnKk0sF3dqnoWNQ4fCY44aY5CUU4braIkaFAM2+8iRWEqSp
MixqivaH9kYkvmwYck1ANfw/vlEL4AVtUK4riihJcu4H8Pt7wLhtVxGQojko
M9tTi5PJhjjLg8b+IrsbZQvli9s00gcOuZHT8vMdFYCF4leY7b3vt0KtU1P7
VL1IH2XB7NmtgHPG2ZGS6pIDb9n/Wf21mrjYnYgCi+WWevPOzZgFsXb4SSdH
TrOUnwNa21/414eFQZc5ccAzEyaErqPGfDo7/ZWtUzqQf7RtgVl2EK1W5bxJ
7GgdgM/MoS/uNJbB4Q1Ve2+A2ZFM3sUlYM2DLYbI4Ky6UnAn0kKJ65gpNGDh
r8wdxCAEoQdsMI89wEQJqoSGKMxDh3s7OnMLhliWoJOtoYgv+MLYPQtVmNtI
fyQJAsmFEj4F7LsbNaMDf/ENwyybVYG52n/jW/nU5kJYm5VHBs6abTMzH4G0
r+HLhnZTfZiwGi1NMFjavOuG7uZen5I14AGxIt+kChtweSmy1b2THsRWuQ1D
CTSPxuAIoG6rXjSTR7UZFG8g/iQRfYfMbXhxGrrXPFQMYaxACU61HmrSJdCi
1fBiea6daXDswsDC0a1DxZVN3GvKAGZct++sOkBzU7xdgPYbx+UQFUG9HkJs
SqPquhfGD0aUnr/joWwwwKdJCDluiPI1CGOkkYHfLUU0gaAFaD0/3kzDJpVl
Lvnh9EtvhcDadh/KCE5Hj4o1dvt5ZKeut7MkWbPX/a5vNmJUXwnpguhalpT+
Yh43dr7BdckgRsNv2CEucWgOwyZNiFAZTzNrPrZsLwWzY+RsbLN1j/cqNyEa
/yKCEWKFK4HFPHpbfqtE+ZRNgL/UsVcN9qUK4DJOT2cTnhoLdCnYwVXHvbi7
P1VL+/eB8USUJB7T5INvSZcBQOR8E6dzKEbwewkFwfyLJPeYhFh3sU2ZTgqH
sABJpeLEaGkjM5u/8EI5wBqKdxbc8nJFVNhLZ+iNVGXSQUMmOimgMSrQRf2r
JXh1EOrAglxRSnEEcZIWs6AUMODO2xfSXqe6cJZziEoxBaP4+O90o5K/tw0+
/ZxOY09jlV2XB0XbXJyMQfyF49c5EGh/TnNba3/XbWgTgrCKu4SGOwbf/DBs
V6XEJxddmggFEKcwU0ZCR1spFHWQltorQyLZiymO8GGueyrgP9R1eW04CLVw
u87vQAPdE7XpsZDY1VHRhCwIy0F+r1PEJnauAS0sS3Gsvx/zavs3cymhAjyA
bN6Z7neEwj3DlxNnPtdoKfvpyeJMN+uPLwUBaQJVW17pm7tpP/pAAYNdSklq
tIpTYisYcgx83kkUYvhaJlWYe2pVZP7DqfMIP++AuJhejU44H47/R9MZsa95
drjEC0ieXioooDtVxVjcPY4gkga3ke6JyO67Qq7ai4RPYe1hVILHCajpVGIb
O82s+nph7GeMbK4GSm8ZjFurB3jJV15lQh3FEbCyLqmABTkrjZUbN71lUVi2
hRF94yJLFnM0QZaXtD319FeVQaTUKNQoXszvPX7pQhBf6U3ZF3Nu2xBXIiIp
YhrSAJhkBeWjpkoGvF3HZRnkvZqokN1+wXGpDbNy3wMWOnYS0evqdwClfd/N
xwcTr8uGiKPqEoRCBCAfOFuOWTOgFDwEc8QCHLKP57WrCssMNY1J/UAI0lxf
mYUuqafvBp/CRqyc7XGfKS6Z3bUItj0UQ3WCwF4a1pgIbnMaBi7MOtRkHPl5
wlwZYuEuCUH3gTlGNq1WFPmQTkiImX0qbej0vIWXJtn84SOhtcISTeXISVMQ
SPZihh//ld0RHqcOt4ojPYXoKz8YMZdins+JoDpT+pLr8fMC3H3koc0FradC
fdItPcmA32Eq4o7cLY7tK4JNWSXdaGMq0A3K/fOpnphqqfxg4jsjRGQItW6P
xR3sUgJMWscCU7n3eYRLMOHz2gzq7xmuesgn0IH8L/4+sm+Ugn2/TkNjcWU7
Oc0+UU3NBnwtBKCcPmRSya40+zBOTtlVuA3pF7Rzani8GDjfCB8i87zKsBL8
61BVN4Ef1QQtb8GXaROVnk1HTcInVlAJTD2+vbwsjdRC3EveHAIoON1oEvyQ
N+c3+g8rqzvkbDAVFv6MD0q8dWK/0751KJnB4v2IQYXugTgluTE+POR0cKqG
bj/qRUlzkQ10mYYGQ30i4+GvGd1J+mqodwemMp2B3mRcguVX+tUUqIRINXhO
pshq8U1kQwyhcng/cJ1D9TV3pi10ocWbW8e0IhQ25+aLUg/PG1lp2Zs8s+Pa
lH3cVeoZSTdDu8NshPAT3ERdxm3B0rS48yWsMgvYF0VS7v8uZ9P8gfby7Ns9
/tQg4DSJoaC9aoif241Pgx0BAqBs+7BT9MrK0DtkUHBzGiTNBN3XzWT48Dfy
vL3kYmZoXH8vqREyS9ttWOsowB8e1Le32HXhCx18++F2MDwNYdRaNjyV9iRq
wSmNGMZe8DtISNsN1czQ4Gv7MYo+zZbEJFAq1FWmk23sxi404M5rriyFNswb
T+qhjQc/qHQRP+HZVn/QzUFsIgQyPhz13Q0fQcjX8MXSA4sG/Pi8B2TGy9TQ
YL9gP0131mBqtPCvVosfeWmvLO2cY6iuh/p+bvW3yN1LXXCbN/6Nq1HrJ7pX
sKEtw3RBeSaSWw6X/TLnAUYTWXD5mpLYL5tJ6RJD9D5qWhBoeskUSnrrvAGg
ndu8rmjI9vLEuqCBDQIrVEGycfOgL9GM3dyUO+4C/Cqoh13z3nTo/2z0dAaF
LndR3xLaijR00MxkjVLseE8Cj4LOQgPhAAMj6MkEEhy83IzJkkHoUcB+D3TO
OmulRh0z2dMD++HFDFji/jJmj8f3cM0h7iE+UxlldnU+BXb6rdgd8vexnTxu
VOKL/M6GiHNJR+vqTWI6NLKMdCDplTukHjhtkTQOULhusGDpKH6NUPpSpQ6Q
84EL9U+5dhrQUWKPfheqAxLUN2rEf18BAw+YCbcodgVdM83hs5moUx+J+1SC
t2+2tdGg7SzhmKGIjfPu35ihL69kH/rkR2YKAtS8qwsa0658jK7ZAgFxguQv
Xl1YF2JfCWXhvJttrGXSDW9SKZ0pOt7FqgYpQOsbb94Dva6gDCP4F1mjhNWG
eDfiRcA9icz5LlVcS717CAuBZ1RPkhZ3efYSzP0m6ndE6LbovRSncPamrgI3
3/iyAPeX3MKRXUY8LwUm595nJXgtBfat8K5DZPcWPbrkdGcA6C9n3wzdtXR4
uu5LljrGqTAGhJQlWXzwalVs0b9w6invtpFPU/kbY1QDyskA9nMP0225jJmK
jP+fe//Zt1Dy8BPWvIwOUOj8N4Nw3AYwV+HFxySow/gCiMlJKiwKFCtQTTR+
Fv3C3mIMzLDZ3EEnByH8Er7JeEmqMOgWY7ivU3ejnlOF99cTTCWmLZNscVBH
f0uBp6D7Syz0PqxMFyCeY/Ch/x7QFy49g5H4kiJmfG/w2nN+jsQWhTa057WR
0Tz4CvRuirIDppUZyAa3zDUuOSyKcSrU5XQH3OBYYKmgOIduoJ9XucqMdf25
hysdViV5gYyT+zq2TDRF5dWBMoEWEDSnnYaFbFb5H0/nBMnDJlIRkTks6zHC
9tJmyKlXhkSWn5LFvsbXedyG8EVFxSkQL/ax4ARnNG+xJMt7YiYrOQppGLjY
aUCWmilZMS2CUv1tL6TrGx7T//wDIk39ZREmrhbcEl2RJoL9mIuFeYlRDHH3
8pIOBUpctp8BcnSjgJmdcMpVDuiyhoCkEzohGx0k8xRFYzStuo0Cm0e8+GTB
xfIxGipKsw2vnHetOK4uzsPdBagJgsQBD19vNUKPkQMsoutLthYsx5OIRcSP
IsWY6QLZBFCaptQq4esP9fyM7wdi4h5rapSCTuKW7x8SIJvTxC1iN02XXgoO
bA/gYV7dFWMphA7Up7KqvFo8PxbjYlQUGJchKttlMG74oeyLS85rkeTFHYjL
JfqSPxLH+sDXbb2v+E7YDPI6dQ9f480Lkwh9KzqT3893DHKlrLB+Oqwae7dz
k7graXUn31YUwpB7ZGbyjLjI5CLIw98hvkkTLyt300wYNbrifbPu/zTGUN6i
PcyDlCVNZg/ecGzCKgbVgXXuN+NQtKDy1Wk7QKZW22RRqdM7kHcdVPkQA6uh
/ytCkRRvmCE96soi9wnAwGvN7wzC1z85D9a+UwwuFOgNEdLE7HJLEsZ83P0b
9UeFrF5kvKG966Y5W2TOf9sinHLhK8fB99JAhRS/XLFkAQQvP+0m8A1DzEpe
snWLLmRL8JPFoTEaUIABlSnkScJwRsYM9vGDiRyC5kmmaSo1KFx5dijL2jpF
OPv7PEcjEFaAPLw7RMR3QmxStFn+GFCRg11KyN92oSolQvaQ8gDoLjbYpiXn
XCHwAOyoOgTqmWpqq4yU5eKi2v74ulTfdhuApC5hgMPcC7ij/Sxo1vP2/HKq
nfrc90xVTpFZlOwOK00r0yiBMM3yIdMvtUJWP73i2o8HMKHXo/sOIQSPCHOb
whfz5YDkHKb2q+b2rWE2auKN80Pi8A9OvnKmg3QYwBsgIg1RkU4bVYd3tbus
0hPx2NJjICWMOJ9rS7bapZrfLkl12DiRumakNmoq/Sad4ZTms9DWOP4rkRSL
l7w3Tg/9GFGaUHpNZ+EJh05+YBcfGuRlCfTsDxk9m9/8Zl5L/jaIFMhsxAIL
Iv/1VDqvFM54BkHXyCHgRBXyJnWNT5BdBFNzYFtJObn/91ukopHjq1cca+UZ
QvEM8Z2RYrcZ1JEifrTDIFtsUt2KqW1FvlVfAqiEwUxfTRxRCAbboIU0Wi/w
KmqKTk2zIIQ4Am26CWElIPWt49Mv3QcRMTbwBkLyuK0x4/lJKnXI5SxGj+jm
i1QyYVjwjeRcuuXpGz9yceWAqy+6glKQluQYxD8Og6ILCGginA0Mavriqk8Q
GFCpgijcvFducO8WvFoAzRLn/wZu0xxcp1BFGy4QJqoTbZS8IUOuUtOJyM+9
mUcT1dChakhTlMsqEs9LO40aWjSe3Zo9iloGEvNxcB6aNSY7leK0G1getsX1
VN6e29aKwZtVezRngYL12rs45nJMfy1HDMtH15/inbhQMqtbiiYGOL6JpEiT
iNvE7lq2+uiDdudsXPV80oWVKUZkHHA5zdgmJg4g29qimqJlo22mniHQogMm
lQa853vSJYjA55Cqw/EEhs1YzSGdAJwRyNhUgQWEPlYidgt6hwvglNjN1G4o
yM1mDOKaUDe48JLlE4N1/MYlXhthd+Tvx1SBDr9/MZ29vrwsD0IZGzrkJ09q
BsrfIYplhKftZFp3iASOZKbXfSl7+kVvBvrf0JkWHmB2MmYGV2PskEro6qSf
yxUReVjeDO5ge82OUNruV6r3AKoXIu/w4Skc/27J60KO9FZa067QvfuOXUeJ
z7Dje0OoaUzxgZwC3JlESdYbvWJDiVXb4RpqYbMNzesGB6+LXd3rRT60czw7
YFytMFxTKuFktVEdHYqdgCRA6Q71s+aCn0H+LJhc52OAwYiYMGLh/ah8fCDk
ur4ELqu0jE2cOTC2QD9aPMrODhZQ1R3LXMY0vC2B+EWQpDo8NXZM5o7+k8Ex
tjVGPVGhtqqWTvXCUwh+nUpQzPBrrees8QBYvPMgho+1WOhc1XjfYwT7aKnu
g4MyDhHf4ObA6nwb/tU/sveVZEF8F5QcHYMusP2mw75kCI6Ea7g5UTc1i4QU
rCAkejdRcmznpjy3sRSq/fG+8Uq8UkVi2qAoOnJCssiQ5I1kwRiVSfEofMt0
KofnG5aTrDTzX2BzHh7ahpcMsGe12OEoqrpASFY24iHrTlGYh+shf+6NVBkB
XIV9dl+oIg/dLOE1+1BNaNlkhQk+jvxddN51dgeJkCUUlzbNespNnBpJb7rs
/mj4BPEWaoquCAb5EkA1XyNLsnwRF8rXUZR/D+a554hOTPqSH/+jkqb4FxBU
mQN9DZGc0X1KUNkBUYOwBHHP9gnE3mmduyzpPQMJPIOWGbZLEgM1gmYpYI0U
Dg4VXEU5b4ey+1FzTyAQUlD26haBVA22p0Q4l9Zo01s0apY8mVs9xqxJ79ZY
XXjQG/ZJcsYg0mZBAGYdYE6EADyeQhq/3n4lJlEDreM1RPsSlb1WXemUYREp
jGIfT/I2SIMjXeFLsVYseHbBk/tGTvn/tyCOL3szlPAS4EgJn6AzIy9Exyiz
bAhNRgDAVt8puEwkJeKUk67k+iHjb6xPnhm7Us8ax/WtGWcKTfQp/1n/LW3W
OIa50T1eqKAfZbJmqnX3Q1+7RXaKlDK6RDgcHp669ASfH+TFuD5p2UY1ZyIy
Z/8a2GSCi74fDPysFOMI1ffUrEPSJcbJGx02nQPxpLigzox1s2faChPVxvlt
W2s8T3Dhppa/Kd8aoI6VoOYH7BW0aKpIoxhRjg+Wj/5PLQwe9iKmIIPvQ6I9
KBsT1WJEUefL4zcKqS2fH5IlEIoB0uxaAdy5pxPpX/iTnX2OpnqSkZ3yM3Yw
9hkesKrfenRCZW1KGCdBo8gvo9Cxj3Z8p/N18gcqDR7XkVySMibnHLnF348i
v9XK9aGMMM16+eF5WuclkNsWsT3PlCgfJXfByqI4eFNZyNMWpRMm9mQoC1v7
gYOu6UJ05Wm59TAWiGz8EG9qDNSIDkR1YtrVYrwVuXo7CJPSgcRYBjxv3e/c
ucE/nLm3TpbqAgiokPEy8HHfDXu/FkozXdEVSlx8R+ZQ18On8F9Zu92B/Lc/
L3EDBmBUNmCgs32LOerDggIqx9U/AvOt08mo1AN3y2SnsoGISV7dG/Q+lvA7
o71wMHCD0xzdl14gAvAnSsdLMic1cVTn+nxgQhvn5CRd9FVU/DsdB9V30FXp
172VHrW0O4IowePEaZ4aSQsxvQBqCNRVAdfo7yNaH0WWAm4tjHInfR4lo5DW
EQ445LukB1+z1DXFYsVosgMOxkHiQZyG3gd6ys+uGYbdUWBLS1Sjdsyeebke
KZ9ZIDfYDlvfS1GzW4BdXQGBgjqmkG02b1BWiqWc5ULMQOlBtb0CHCQoMDt3
zYMbZDNjMODSfu5pGjBvV6GFT/4y8PauxczMlNJDgtA9tg4hWfIKjf7TzqXe
72hyEwsunQIbtbzKZFCHF1slIgLlNB6nZk6PPx3kynccUiw1aTozibWiV4sT
Q3lV1f2rdCFBfIHxbYQBYfWfnjdR0780heTlZ2YSrgfHFxYqPG3rPCZYwrw7
wUuFCjarzMZDlmk9lg3QAIWkutBPU9FSMaG6Tav3H4HPC8istFvyzrnTHn51
fhy/jtom1AMfj2Wf5wPkfMdHk0gaKdWtxMPkl/pOAR12tD7WoW3g/E7jRLHY
wjlGuDpSKwhNz7aZN/IXkOVLNE8KdbIDX1LkmvBe3zM8U+Z5CdPipjYzrj3L
wbDrDyY489vxQckTZQhVyMLLyyOrzsxqghZZHzCRpcEurx1UlQ9VnW4e1B++
M4DK/U6sLbvJp5sImM5tzzWDYSNrtuQMN1c8JjLwKom5CNI341p1vd62kSic
BhdK5A9juI+OalGS6yjatfS4zSHTlGKW/9rf1w6tzIbiqN7Aa5TcHwC4Ojaj
51vNAl5JauxVlbnv0adaiWdGqFvYooUCsHjxuK1YpTmtrJ5lUU416bCZcNSu
pmaKDver7Vwg129B1y3XAMAu1qrab8natTX1cKV0hZNbgtH/n9UpgBbu5B1b
xuqexYtRdTgCu+g9VZdXSR30CKKpJUVOUhYHo6FwT/IqgXLbpMd22xqDMdbr
I3aHI/jMuCsVN3avfi+clIza/t8KqHTF2FnI7v9kQCsyjDczmCXjx/6w2mT4
0M2OBw0PK2LSpycsoiZTV1U6ZZ7LvJNpUOnXeRDtk4KXJS8hUefR+7KCjkQs
V2Qvv6lilfWvZBbOtw/kQbZFu4lNqO58cmhu3akVZ7Ak75xgEKARFN+L8qEz
8oXAkx59jx8ZibOHXcMxMziPKZWsAO5mVczgwLtd3UjqC+z3It+VZu+ErDIz
y0ok1AbdHRifqD6xNE5yAzU+YqlI4kRzDaMgUARi1VlZqwxUYLC52bN35IZC
i2j5BtHh0AxMIR7UP1bTJFE6xFcaxbWX/xPh7NVVjjVILIyIDpaTv47HzqS0
uxPt6Sl8d4jPofXtlQ34bmhsHejbtTCxoBKJykhiLujQfozYuZSYCP7f4c9g
mtcs6WQ23io1jL2kxQ8TGVSvrmkPsI1mOLJ4EvLSd3jV5rtxWeMo4jygd3fi
N+xHRNg1HwYFO7h6ka/4F7R1qjPpe07XVQpxRzmlkULe9Y7o3cXJSCAgzgJw
/jUsKVcsD/q4zVXRrKcTOekauSZ1zjwt8hj5FEi3LMcMhbhx7Hv4faVfr60p
wrPrkH/ORBi3B2zMmNqLE111+2r85aGJ1uC0hlogvzQsv0lTSALUFha/SsAj
F6R+1jQsjU/M599QjpND/wIMrSfUlwuSOACZcQG7F9vE+KPvXuGGEDrpJBhg
iyrzrmtuBfwyxbKjML3Ha54Olxa1Fgj8dWL8fNIdpTsViEcswnQiHXS6Eq/3
EyQRXSjUmnj2/NOeJMpjOlNLU0O6OqzxKYxVASF4lQwzkdXN1uR4rwVAmEOT
V7wEWX/yTIQchLb72+9wG/nmRnJr+Re47tplc2ngR5M/HCx7f3ThuI2Zy4Ny
uR11jwyTSd6mDQAdwfej+LpWRAHjYPAfhdh7vhpucdeRTygURQsc94UT6M96
+XIhaYQ/gE8lzdF/9uZ6BostZPKXdRukppUctF0XjTBK517cVEvrbrNzWevg
rBRXT0VHNNLQSxHii5KNiGYyeBCURaGrpM3xYKL7LzxkfCUCnOuTDB9I55wy
iAaH1VrHhajrS/jyIIO55Rqecd9+ocxEL/V6ovKtjHnnuQMKjbQabDsUtmDd
kxlwrTTDb0rSiHlIqbNhelByPLaOnhapZrFTBNWYcUdR1Tfwm8dfjdWZd1jr
ir+9cA6d+/X3Z7hKfFB2f+F+ZCfKW5e5X8Sn6eDT3PrlHur+HJjmfnBDXnbv
RhXpI55tqXTIGaPUq8qAwl1YxR2S6tamFBtgwEpwqujwvyqhmMIlEj73secI
KuZiSJQG7if9BW2OwW+G1jhYqd67L6VouE5TqRrPqNBPHdRmdVenDAItUrqj
DBxi5O7GhvOhHfLNyqRBJvKhW01ZrgFAfvIOHdEpzg9gfOfS+0G5SkCfwvTp
7GiTfVAu/gS1inNTe0Zc0TXOMQjz/cHX7iBx8ETNJ2XDAJunWXuqQx9xG/kM
1phCbQamXk9iy28N873v/itWyvIx23Aqz6nA1nZY9L9ZOwb+A5io3jXruJGT
ccZtNy+CErZ/tENjZPXRMp6gNCGPf+1iDX/339tjFEOOCNZoxotLSqlkz6g1
7+vmcWsUH2DU3ncOb75FAlTPvhXKqahzT6NxJztkSvNWQsLOc6S2r2VABQGX
mrmX0z3qtfSG6BQUfD0uWNMi0YWB8jioEuYhNIyb7x1TqghCuBoVlSXa/CKJ
Dd6eUVLF2adeMW3DIh/snvngAtbTzpDXVZYgGVtWCpOrz0OgYMdBGxTt/eZv
IeoF15o8BMAoAT8nuFOyVZejJWsj1Vzcu0QWP6q9Fj/B9eSbTD9xxpgP5KoR
n9mgPETjvNdb4rNZXlCd7oNb6OYFNyunZmB7PC3OjhHhZO6k/uDGgi1dwWC9
n7WfjMQVZ+93wKgsG5KBO+B/TLXqolN5/pnvJR3ZKd1O2feQGOLhuJHKTAhe
oDTUOroPQiFHgkQoWxrrd33zx6kMmli9iaMzyqc5H3Q6P1vnlgv8q5AYPrRD
WisxXaTtHPYhsRBVDxKICvj4NpjLcaRD2zO8LqDlHeXSmbttePKTtJkcSEdB
xLxlaThGmTQsc5Z8yzFPInc0OH+bqHP5hx38uM9a9tPFOLYP4HyqA547R6cr
KH/FAeJd0b3qh4f8bJio1aVV6PRrjtIxVqfNJbSUpro1RSl+la/Luji9VNPo
of6mX63/RAV2Yp4AXFQ7ImW5FFihKs3jn8LDZk2lvYOXpAluR3y/iMKCY93m
5i79ckj5w9BIwdTICpUuJOcA3JtlloKePedbOAS6q6UAOIw/3yQ5ZZoyFUc1
M0UVrXwQZM9vsrX6W2lKIu8GpBM97NefrBSPdwrdZLcNuA1IGyqQn4YeZLDw
yoDAWuuDf4Fbs7ilz/mSv1LW9Z8MZZ0mJIslwDBwFWh29BIVLLOh3DzfMwy+
KHZA2PuiDv1oO0DJ5R+bbdUgNJBQguUakcQsMqfdaZmXkxK2/osKqACCAIuy
uAqx6kBzOcqWlUMHJlgGwWrWjNkH/WK8H+cXKT5aPzVD+1ouRWlHwtG7BcRd
prFCI/GpNhn+1r+00MQaSeq3g3KRkOvW1dXxxJKULRPXptb5oZzFqRxaEWUs
8wiDehwE2yTUe8Y14DH98VvdHX8kCgzJ3AL+/u1Qs4CDu2tdxXrxMn2fJCya
1BjHVTEiFshYfMdG7uE5sf7Li9nC1yExOhXNfIhKszZFIphPuD67QQh4CNsR
w+pC3t/7ZFSuOUorGLBkdw/ZaA07z0S/OhRo4rHAEOMnxWxq671VnUFuiJLK
mnG3qLy+P1L8u7OojC08wuNCa8780e5L2P1zDpJ4xfn68wyzzo6FgnW+h3Hd
ocp2eIss2Kr3IAq1Hx/20OzB2CjJIAkMQ8V2hX9oj9EpOnINvKwK98riBBLh
4Qfzi1J34rzwXA61HozfIWrkyPTwpBqMYLcC64vf/SmufX+QHnaKV9FCy/rK
Omp31TZ/wZ0z3te4yLVWe4tXxWu2a08XiY/cPLj5dB3wCLy+Lrur8l3MU3kt
6S1TYTL73gi9fcEi7RDzcdf5bRSjF9z7E9cJAXiAbm25AISZZE5lfTzT2B6q
7ypww950/g04xaVkOyAuZzANichg+HSdu9jSlWcKc2rd4Q2quoQNKaWmzZHH
1vZwajEaAFxg77srKbfr41Opb5x4Vfr8QOYpkX68TMoI1BQJUoJZ5fHGlsqc
ISqWNURLPxYH0ee+aXwYJkqdNp+pAdaeiEyFYHd2zUXPgvlNNfbYu0cVX4Km
QbBidPil/ZA6/OF8Dk4thEijUzUZmS84/CYk7hGK6Xb2HyikzDDZOWNQpiH/
0arW0ad/Dl5pvMm4IsKn8+y8XFiQ+9p2DlFIZYMWfo7RxkZd4YS/WzjUGoN1
TyyIfou1/MNXdnXzujykFdcWgo5+WR57L7AOabXJ5qo5/HCNGHziZQkMaqkI
8Cisze0+wDpA1Z/lc4tH+OKACNWBl2w3ncXumIXLQZfbsen2SrSNq7TV3VuO
3603ha7pFfOrPdDuuoVvXSjeKIe4phJ7vm3FZcbWy5NnptBE9+nEwt+qBAOe
dUEhIW7+zg+8ZSb17akwvIKJSVkY+KgOySZrHLXDQ84Ub7fw+eBML6cNlTjE
gFekKUYSQwbINRyPyZttOd+DlFt+WvZI5IGJv0VQN16cH2FgpKOqUTq9DlF4
WiBaeAnl0WxHsyDoDQdUnMFIIlPZxRvpItIqb4QTcjwwdv6cM6nLzwu0jIdw
StYMisTAD0ezaj4c3Pt72pbdpGB9KnDBqaU0rfCwCwH+MTbn8/2EIwGqYg/L
2lHgBFv968kOpzUbZGCoKxwsLHu2a2s8KUtrkN/ohRgQpN16ZiCYKgLiA+ER
8RSWZvnuKDx8igG3ZKoDXViqJdMPU5+yYdVpVTvMrcJBXOaao71KWg+UY3TF
vhSs7tycId62T+KJmbUryhWx522E1DhJFTtmcJRDvSn0KK+Oa1h96gX2qeHe
spWtKGgC0fGfQ2zCha2aReI2UYVbc4FZET2zSDGmJfnEKiLXIkY7qFwknqvA
qRxCDy7DxmXXFQYlPNMRiLEccFfxLE3I0IzHdyI2SbZNzKxuUQVSfVynzhBc
sy6lA8/z4HOy1H/cOL1ldmZ55Oq23we87snqTlj+78UDR6d2na2v3vNTI4hp
F6Ei1gwSdpXBgqLsfrPv7H2DqqHVIZjUL+kXtej7LeeeE5dPLtRb9twzPH/8
sMWMZ11CUDu8oYrTwPC4mPXOkU42RDHmmdzI2JRAivJfaRgnGbwEvTMi+EiW
apP3zcPDnL5lhjSGaYlv9ls822nw1XCN423HQgq3HO/1HVsen2dZ7v80JOBn
PpGYoyOu1iBBasygc3DvId9CB7lV8qZDkmTC2Xt0v+JhRqGRixJbOBaQ6cX2
LXqERpe3rT8gHPCfqeLGaNTTjKIEGzWIgY105l/AGMTdASqL8D/MH3TYGyQ3
oe4Yu3/aR1PcEWY4JdLcx9S0tXUDO/E86+XGbIELC4aqwvKs1w2vQVcxpbf3
n+GmnR3f/MFUALroG+CODl4yKZfROFoDt0zesOHsGVW7o316myNkkU4UkHly
M/ZJgBtHLPVDNjT+pDVfqQZLBEzb6JHe/gdEyjIPP6irHaXHT9AEdOB0tLkC
WPU5CwMuhp/wXYVAyGvYYo2T5fz+6ZzutnTobspLS/Gq88cfDfijg53lQBA1
Qyr75MI3VJyI3h6hOnqQEk6tR13vPJJcrtAukpq/jMyWSNIR/pHkJaoOO8MW
oDDZaeH2jQhEp2ujSs/v3eSAjZ5B3FwP+O6mxjn/ALh19L3Wo67bxcQSupM/
Kjmtl0bNihUMd0ce64IBKvDXa1QQQqPqxc8IbzSN3edTIZQKCzynJ/lM/x7s
iwaHBaVb46U0NLvkXDFavTdvRG9o4XJNaJgKW2PeEbZjXfMdFchFjxztIZJR
ydNhJt8Im9nSoQYjmM4ktBdy6gRehl96l5tHUo9imaUCEvY7zmZYsq3SDn2w
BuJdnq6guPLwdxytI1JBidEb7OBwWpLBh4IbbHSlDmPxBF0UjnPWuJsCq/hK
yJ2yyVdFoAdexcR/in0FIrSE8Dne157lC7N3a5QEdwWxFz22l7KYuyvHuDyk
73xfpMDE+TGRD4TnddZ55ZOOgrG1735Y17WpWg7RXOSh4iW1e4375/Vja7Ar
omyxrq8/e4Ri7nc0Bh0lRvcXZ5JE7jDsC9/L5eG1OY+pF6DMPXnnyxspytbm
8cyIX4G08HJB0Iyh90LMyAWdrF92BvKTsozeh+1Klputi+EGh99r8mQ4URCu
5Rq3upLy9iZ86qSx6xcOg29ANohPhdc2J4vZNKKtr7Oe1e/M1a3EuiogKmFB
ptxaOFX/1B+1iry3+I4TJ2rDQA/hMnfdkgDV2TluewtbHlEiBtBPaZG09fST
dvtKRexlZ7LPrUL0jmpDhcCCY+jwWymBpAb5XZmrXRuoOylJPxYrht2Xl3OD
WwEPlraTqiUIT0JvW1hlhlmqlIiSxsBYakRLJ+iYphravJFUKwBfgQxzHWaf
SgGPxslNSLC+BZlqyOrRCu2Cp5uilJrDicIi3lo0b6PaNa1N/RTmjjmPN1cb
X1QwQ1SwtOddSp6giV7ibKGs2/IISXGlgsG7pkvtwXEUFHuFgUbLwks1oKMW
YHx3pxCLSXjUxrIeWJWRJgR/AZjrJJgnL3s7GTCe1mT0w2H3he3vxrM+ob4s
PWBDNgV2dBINiBXq99PJBwZIzzxSRqPiBXZjn7p/wcqz75uewo6ZDxFm5ip+
+GNZ607KuTMmJ63iAYkLuFDYqnea3dEqThoBXKd3IT30rQ6RSN5/1R2GEzle
K3D8cQczPWQhzCN7QA0S9DYTa614yPtvJQwYxEoMhtrW18KMtsVH49epo1oV
99m3EALmwk7h+DaFn9Ofemt1C3cM0pQkeIfpxbFxR6nMujC0Kx221WsLUT93
ICUXlIDHGtRVc24F/1dOuO3AYgmQIoKQBe3bVeMdu7BS9FSyAFGGW51GB8BO
Gy4UW9CbGC9jcfCRMqTi1Ell40GpzqoaSCAiIzUXMSfcq7lnIWb3FD1BPzMi
jz5hcqA7PPBCwStqH7S+HMK4R3g4ZAS0iwSEShAVyH+C3puFpRg60XOF9+he
fefwAQZ+6QrM7y2bIOkRXTeUVtrE0E86wefLTwFc9FcanWM3tuDVzmV/FvSk
T5BqpGXhbDfcgJTtP32aCBhfxGmt7XooEn7LIPx8QJ6b6FfpjF78WBtf0XQG
qJmnZuIQfu6cO0jetEafH2Pq4CL5CI7lwA334SnZkv7S6J3+SEdSMUtwxH+G
RyYXg1fBfIX4jAqn/Xk0Et1dBTd9H/T42GyQkBvRuPHZypfWCN4yNi4QRmNE
H5nAaCd2Ig0h5HjnPkTfbj5PvXLZrnoD7xX3uO5EQljwl26wcpddI9Xsc162
GN7VRywVCjkaQUDllDL3jEJnKsTFxhaqMf0Pp7R6StIjq0u0SEa9+otATbEP
1xRjMicM1Yek+Mc0e/vFMfTCg2DYy8HHgx4DIdkt8BcuNMYUkti52Dc9lAFu
TAtaPUmQdDhRh7bafbVFI2+mJ9trEliET8Dvuyl8ckssYAINBQOS4Pp1q6m2
hIIgVDRz/4D1pSfBELHbc003VIkUEpx4DIw3o4TrLlTFERSZBv4dgHUs0R4k
uxD1pFzYvC9vDK7KZgGaiNqYMTOFsir3XMGTuMR7dlY2O2p4LbY1pSh6+331
PgYO9DNBLEJDXLn3DU1fvEs8OBAuYlSn8LwPRZrnholbGs69JVK9lILXM3+w
jVlm+1BWkS37m0Xh80MxXCojKkOIaqaJvLLdHr2GorWkk3oQSqps2DZFGZa2
3qgN0lsRylTl2Hkj4fmBFkGWzD3m5KOmsaZq0bqRU1seBC/oQN2EHDbXPW3K
VB3uNXN7gY4WRCUGTOEd0GvhoToRbBXhG7pitMdSD7KFWhjeK4BIvCcaeQNk
YngmbYalE9fJZr81JLbVLt+CyimrEhFWrAO0Y08k8biqr55xEXZSyQQJiaMa
vFNBZA3f868MuSXRUW+pWkhlk8D2ysfPNXDQN2BLMLEBHcMywYXA4YRWkFIY
gp1Ykl1S0FCuglnQFtF59dFaNOpl9k7AUZk4WaF1StanVFLoxr9OkvERsR/n
Knc0qtA/mySVo2WOPgtdaYBKRhsKbsvEHUtZbftkzGYvXHq5oDxD/sy/+QG7
oaZ3M0x3Xn4wg3bsoFavTaxRs63JvWcggeKv7xYbjd4M2wnvwKrpd51i8A2O
R3iT/1knaydvaTJxwgTD6K4et1ItgZPpidRuKfZyN4gpz22WNd9mlYVeZior
D+uWqE/414FtvdPKB6+EviuB6Lf6lt48XfV5/wEzz/JaiRkrxDy8lHRpLkzl
pu2FAomRLh/9i8GmaP1ipICLkZ5g8rU5YPTKjRAp2FmnBonmLqkzgkw1sfJP
qhYa4hLVJnrNjAdAnEx/JASU/2vCeU7LOy8bVq++Iq2fQy4IAg3jwzjX0xdM
8/Zt/qi+cZaoFyMvkHrMj/7IFdfQBbVT1DabUVnekidnFVLfs5zduxoVAe+e
70X6iC+i31vTRx/ZPO2UA5eIAPceC+KiEJ1UCezVn5EUw9ZpoXtZrlHnmtt8
avJT/8vJ5TkevuiLyFlD6kxmZyFz00wRpYeFp5IkqXCa6aEXOUhuPXvtifd5
JiLKatkHrw6a043MZtYIVw6gVeUD62O4a8jHrlwpuYjDNv+WvZxaBkks53u/
4be4S1jaUg0OmYjod+YaWNRn8YlPq0ENQ6M8lswgtOeYzU98Xjoq2Eipjeaz
qjXpSaPDI9sUl4wfNTdRyLZ4MyI0uS3TtOpiUB2RwVA5cRxqjNBLoSI0DdoH
T1kAZQvEmcFJQIwlRoZCxhCsE3gvyvekJ0PL2B8lWdGNukFXXmo2ZY32wImG
6DW6NmxYNDHfaZwTlrYTHJX2hNyLqbn8FFLKv1LPgphPR/E/xlnRDjbYdzIY
Sab642+atBuVWa90IobH5HtCIJUL0bABmBLA4p9Nq9M6aW0eEmlLa7zzULEZ
QuRrhIucnuFHlIdulrdg6NNkHyXp/6g2HMVMK2Ex3nP7LT3d2Z4Rsn4NYm8D
oCwVX0GLUInIvbymZbAYTXMVUsUw8MkgTDWjfDchwt6mhaClqc0cXtYrodTM
AfevcUgPnqqF8s4NnRxNNSk37Ss+QgCRN/3s+qmUNndeO1ucvA8wsRZMnZzO
EarC3fVzQx3wCqMZ4dp2ExXkhB4PrWO+EMgHwp3OanOpij1/cGH0guC41pce
OEGHZD3ZbAb92KTqIateH2HLUCVigs6uAiPiB2EAQIMde7hg8e63Q8XUiHAy
tmDNL6M+OqstKZw0onHeLWJdfQf2M3SOSWGshDJkLKq3iDQamV0ZgRZQH/4P
MI5tGTKPLqdpOG8O0c+2MO9wtU24JN9zU3RKbz+RbZERsBqQR9TT22dF6bsl
7ZsHTvXRZFnbfZObXrI4QwGaO+RsinRN2O0DVt+mW9ljT7i186xlE2QBHz0B
qxC7a/pw6BaFrzeT+aHv5eQ2q54Fpx/cFXDDcvi/AcRY0rNOixzjxwg2I99y
yWJks8LJP98uM4XOY5EgiWRKIYBYZCMgig+eT5VEc40F8dkP+uErwiOnYXpq
02lSVkjj45dt7qkj9N6GU8+rfKpAyEYli2++7Q1AMYm1G7gjntLy55MPQb4p
66UNxKRsDzyNEyq+gyQBGiKSjADgTHcGhrwJwmK9VvyeN+ptyIgPpLGEA6wx
OFZSFbNQd+4I7Ee2U6ZmBA/33FBVzY44m5BzjLXfpyNxEGQjFbpo9lZsiwP3
BZpjBhaUrc5PU0QTKaRTlaSGo1tqrSBSJEULvUXdu1H3VoXkiPKFXQg/fwDI
fm0oc9P6whB2+b87W4ycgqKZWiP/XeY2J6kXeFLHJgNzGOn7fFcNtgzr85Xe
EmSTO1Ma5G4pDLAFfj8TE//dkM6DRtTOQR3nfGBCFetq6GxzKukui7DoNV5P
fSSCZO+Q6B8OLGeCNg/iTyHz3426uVEcgMet04OsLv+Ge/AEh0nrgJ32j04F
lnvzFIH7EtXz7WsqYH1dkwDO2aRIX/aSTRTTxZO8N6Fbpr8SiHzKdVSyQc7k
xekqIbamKMv9YijEQiYn1vc68ryR1nPK77CFJXrnDwDCWr/0qX8f0KCl0jbT
YcxPr8sXkQ/ZrdPpt03BuBf4AD0CzDVELJ4o+27FJ5veBWPfO/3uFvzZLQ4p
Qeu1QRRgebMcBeq8EMUgKHBuDLJrrd32h8/9bYGgujWs4FuEf+x/2W//inLP
mYKZzRsEvWrxwVYaOX9uPEKohGwQhoNV+GqcUWGOfvhUWIT1tyoJbciupxtc
I+mgnS1JHlWRE2dJGzvEwtFpR6s0Dlnt/i6JwWL68KA0NLC3vJLje6GRwe+a
OC+/24qnobauknbHu3Rtph2ykpJoPWKCuxr8xBd2q/jfzOYxgp3n6gHOo2Kr
s7kBYpneRjH6DMkXvf34arhxc9ffwYjOi9nvilOmZ8C4JLB0nxTYxrwu4AEY
N8bCr958cTTBlkdmvDFKpKBV2HgxvFHPzs/TRHu8iZAu+dl4b6YudLz6BEiW
6PeAOuHPSBnX18nMyqwXVgB8tDuiOdvGQtDX0TpJLkh/c9mNxB0LKoyUj260
Q0KMbMOHv00lewAjM+TgKPF7Zqae/Jhc18NqrExW2n8jXxdCy7cibioxeEyU
SB8baZoQS2QgbvTHrxPs0YGuw6iRn9v+6T9uC1mamiGybxozFUUrVJJoRr77
vo+Pk0tuV6CJOIHR42NOANUKh0J+iiCBaUb+d6j/vd8xasl7b2CtX2iuOYj9
Ar6jB0z0TGWAhYXHeeR5My+HrjzpcHLXOLWEL64k4Je0MqLt7JSx2fp/oejf
s/6pxz8NYpklqi8z1iDnipwDTVVb69cESuBukf75oJifhyRjOx1zSaVPwRtm
GObGfeUEnLJ1ZVE/1huqeLwKQM3EbQlnqVff1Zh6GaWXEjio6+LHwBOBXDCC
GGkJviPjfmcT87Xz+CSsJjIudhN4yHlxjs0lpgwKguuroZHj97qcZv5dUjsv
CafpfstvOK5PcEUkfgY4O3lBGezXpQycf65LcFbcQcqi60uFmwrphO6kw5a/
ruSUN1VYjSbwNLoylEm+6KSChH5SFwQyw8vNXfy0XNcaArcuNe5qXj9xpYD0
NKvs/z5Jlg6zf2fr1MtVu9lIE5OlrmKeqb+AALaLQp8NKxFvaLTC0+ZkLR8P
MZjc0pJaZz3p/qywdU26cJCSDu3IvAgAT4O919JkAotEmQ2ujjuTRasz2xO+
SZHsGTa51yC4+9wqr+sR1fwF+bX5x0nggYeLsaGgU5XcHHuJc3qodTkdtldV
SNiNIvaiJwW+1ief7RzeC66lyRtRZbQbqTCcvp/PpNuDWfSog1JEuiq6yVMP
8B9TIJnVJMDE3vbpAGoy6/iNlgFz+HgIc537dOE99qutP4uKVYmfHZCUOXMZ
inOBPV3Bq6qNULENj8TEo2+BVdSYojnC4qV97iIkLYlrHGCYJINKlw/qhyNY
FRzK1OMziXHHs9sut97VtvWOsW5csN/Ajd2tt0MiYEIsO+gdvU1MO2ThTSC6
YSHnOrZ2A58lM3Q6e/ejDXi1PbIWjibXZ3cAZosKEa9h5bduwghEc9LyW9wb
WheE7YIYKRDsCZwNlcZAbLDKQXxiT/w3uCBwulV0xkRd6eecBA/znoDxRLE8
rdv94cThs0c518fM8XNIrsNfOIqDS9MElAfWniKYhAgAlF+5SBIuaCD6UBPH
T8RPvmnqBpaLb2R9QvdbxHNK80w6UuvaDk/aid6cETDVlIqUcRf9oKgeBI9Z
Cbn51AkFPpkvGom6wRfz/7Gh2X/oag3DTs8UnZIqEh/m8PNY4fy27OvqYonR
q4sZKlkWg74791rAiOh1pOOxqdULNJvaN5wO60/Co7Nnp/daXl1r0nunfB+X
Td6cnrPfn9L4wsidivkjAiOjeE7Wa84agJ95Jd4qR3DCGiIZ754/znfUmBhh
EHAoGmiJj0dOJ7iuWFItBqCypDDxRddsGqt5I3Ui63vO6+gk7MFpm7A+zh2C
NzWur0xXwGZTbzbrWbB0DlAVWSlgnsuOrNebttsHuOhvSvgZ4mc1ysZA/M48
W3N6z4dRficjQ1qvp2eMZY8n9MurCA41JTs7Q+ugmBICfqwUPXoUnsnTxwg2
KQloA1JCemn5urIdlyUNWhFD5wSGgD6618NUlIR+yEkIPM3LXGXzF0cd5oZQ
YdyXFh8mxMgwd/a/cCbD09axf9DDQ3zICbC/stUVqNhXcg/ZFalMmH5zEgI4
9K/9e/hdjYZlMjiZJjnfLiZX1UhzW7tMVfjGxSd4/stA8khq9KEtrE0h/B8S
F4UWJRT73DmiqBLN/RZ6HYuypt4k6QU1fL7RfLQBfD/fuZBkS6878oE2AgSZ
KIKecI55+NRBKybbABDYpOpZtbWK8TWF0v0l1ZCC3VOuYeqLsXYy6ohTQsGu
LwIcm3vMJkrvVTDO7TJsABKQeoXJ5ctu1nkwgrGjeAMhos+jU9uDkVESP4KO
8t6CEFR+57GUHgtVv6wb2yhNHW/eQTHxM17kNKztL2TpYHKPK/4ivQn8rlEx
H9mRGoc4W099xpmlWvT4uok4stqUhgExyRshp0ch5Pbsc4EOE8af/HsBrM/m
HBL+rs6H9ritFEvgPG+NEn7uxalrYWKuwCSg45HWnPr4tgNQ+1qAsoDdXC1Y
xgF7tuAY12daS63Insa/EgA40SprtwYn4C0IQ8JqTUC7RHa3F4aB+YCGX9bN
jU3DNBoQDgh/h5oblR7pEtruS2mC9z/kG0AdHLXu8g8SY/DwFN2TkNyUTJRU
qlA1BWQ/uWfMc83kNJLwL1AnttnhATtfmk0cyVVF5yaaLYAlAiZqSYqOEraS
yrUj0nLurNjM8MbfV0JCMX5gDNqV+jbIbjx4z+wiaNjBhKV4iXhPJfEsKWIk
fMfF7eo2ZS4itlceBPc2qF7zXJh3RPUjWZrYrI5/YGgLPtpoIG9vEsIf+i2Q
YZAjev9LXLW7tq+iS0RhdKYqgpsnmzTCU3JZednCELbQvLfn/S9PrprVSMbi
TTyEQ917rNNgRSb6XR+myZPKG5cdZNU/5UF144CizOw1MlyTi/p8CyCg7RH0
rnjT/s6W6VTwBAwNLm7Z/7yFVBuzRvbMk31V8fre993UwUZZZNqjRL31cilb
9jKPe8fMfpKEi2aFpwxFFFLKK5H2ChfCZe4PgXpxHsn/FO7PUQJycr9Eof3R
FiarBRSdaQqS8zP53cEHlNIa9wnPm9bBSFweFrPAph9vNGlaGmhPNKplS5U7
BjlR6kCsmb6lzRbPKXch2r3YxLTyQe9P0LwxiCkj9KGOEZJedRZVyp1MH3B8
uOCuUdQsfqgU7EZ+XSg/AmVxBDIa5nEQ2oSmj296/sIE/XQHEMgtQTcCme/P
17L0ofUpwV/053S6vh+NMck8C7lOu58Yz2MO2lONyMNJAc2xYg5CmkNMFV9v
mpbAT3XRCJnEdbnBVQ+rt3psRd9ZTuA0AXrT4z60x+Jz/Iq+texdhsxtUKYD
z6MjcE2ZmuTTjWM26oaH9HW3j5YbG1Z1BOFQKwnt+SLeRiiFhL5JRZJqnp/H
ezsaW6J8YGZ7OlXthNxPHMME+tp5GsuGIMvCT+whRTmFhzsgVZ2/qr0xrHfc
Ji9Ei+i/7brfnzkn5uKoWXMa7+sj86pMDc3r/Phb/kMh4in8GqfzbSDYO4UY
EVms3TCJVauatoyZtP+7VCkHN1RgiYIyttYza86opFCea85MPjUwsNPqvEQf
x6St/U0fowOJ8EdPYMxZR4p4+UdKl8EeJA1diGcZ8v3FroV4cmf/wZ7hM/Pr
zT1k99F0rKrrHqhtaGqoG5EnQCsfOz6A/o8PJqDoQeiz6xb3bcr6WzqpK1/L
vlcLEa4tywq+iPTAMUO2eOKw9bPAJvC7zDZZt5yhJhAPPWJNdkU+sFoaU7y2
4rNkNnydNwq8WwRDWrwepmW5bqCyGOkmKac/RW2nONjMkAgIz4bruraQKmjM
QMPvC4F7tbyPv09rYvXui/nq2Ci7Sv2wJe1R4MSKGxj30LqqgEt2Kwk+bIgY
wJZew6ihPEo9r8Jv57L1HuuOJXVNAbTZ/Ltf1FMwjOzMR6IdHaTpFezUgTZb
JrZPgnauh5VIa/E2+KBHUSofxpa8kw2sVsn7Vd0Csc/F2frsZDe8YV/1DLOZ
fzpgs5XD4RBNeth9LqWW54PC51HSNff+iLZBXfmjV2faMyE+5j7CPHTdqMCu
C761oqa+BmrO8RA3zpLRbb4kV0RiFdyYeq0p6yCPft3e6dvcpyMKD9ZVDdrt
EgNA84JIbyg/u7o4GsI30LiF85Qroh8mA/IgfFN51VNVMjE4oqTK+F7sgMYa
PQ+5ZATaZe6P+C4ns7WMQ7ayQryE2A0Qk9DyJ8LaakIZ2NfkRw8R0ofsmtEv
WpJnDoG4iMJ+ULoZjFdNNV2wr4nRGyQP80nvQ82us7J+a3RlrdUGFVV3MHGL
uzwXNHRveI2Yf41hc1IQiUJQdow/X5VkbXx+4kCmcU5dg6JHAb13S3lwP/Bc
98EdB6OG05VAVGB9zFlvG7knNeVKugvPhDokkRUQQe/tPk7Yaq1/w9sQxcFt
Cbdjm03JJ+iYrqB75CF6+6RiK6PGioIauvaMvIHXDGgKuaEuo7WwWVQ0OmnW
Ny+mFtrfyGsyvw4wANvvztqOTCgiJ9GjC7THPL/ptm9GBDAT4ogL0qTk1iAd
K6Wz5o1Y0745sasH5S38kjeFvNLfCW1Y5rTTP6iUgRQqiMTs55fUj5ZWPNRz
NvS2WOvZ7FkvowTyEJAiJ+z8tzwxc7bt9WrmpyR/Q/ziHe/mkGAYW7uiC/uS
IH8nUhjfH0q11+k0n9EOSjJwYZpzQHKLxZ1sG0KrYDWkHDsYifqV+fKyjhH0
HgCl41bmyzzXKAoOOR9yQOPb2Br4ZGkzPC5FVVPwpYkTE15/OJgmajBcyowd
8BhLhkyV84iR52fN2Lgpl3MuE9pPQFtX7R9SQwMd1Xm2lMAxwPlZzGMjm/wX
XvxE0ADLkKsQWPAZ+8mxGsUHer44TwqbMMzM+2Cl2G7/MV8SIb/1IE5paw7A
Ulafak0Xjfwv0coN14oETHBjbs7gdIHrGKYiArSvfi6IFezncyb0Z739tHKR
vgkTCG0nN/priwWTP3S8u0Laenht1IeRlWgmj7Eqp8NxAmluKZZ9YLZKsFnw
pYtbX2+rlP3gpNxwamX5SkzltUI9FXU/OeOrUGimLrtNHdkh7xrT+xF8CYEv
oYlyGbNrSjbbmT0DkKXSIRcu9/3VPCpxqWm6TCbUax8Rtd53+TtwRShXFCfs
x2ASWbDZqmIYzzdY3vQVOv/4x9lB/QThWJKkJqZwcWygKFz/9B1OKMO3u7LB
meUawg387PxHK/LEIGaNYJAdvT5fgnjNAGE7AZcXWf1DO9w6IfDGYAT8xAZs
VvhaOS4YKWVyLfMK05EqPvvbzLYnVMZLJndJAdrxc68KAqjLa1RZ5f5rQ2E8
j8b18nRdnBwzk+Ue6c0JlG7OCVccP4AoRJqTumwuZO8AzDsXy6mhZysOWd73
aA6tqmSvTP1YOf5yGTdjvlC4qGNFjzQ6MgQm1Krs3iRvCNmh/2qjw9qgJrlX
eb3leOO8q1TKahXVvB+nTI6kj4oeya6EE2IQWcodX79go1UYz6qOpvXmZo4N
lDlxVsPAx79rH/hDBSecxmbBLDf7PkTaNY3VPLRa/RF1HKMdwTmVn++Cvils
MsG2a78aOxZTqSbOY/JW7k0Hth8TzB8y5wvXKnIdDMLL4hbljynG9eOsPgjd
0LTuyCF1U+02+TnjA24XQLBW4XUsFuqqPR7+3y8T6WoqoF7L2CeaSek1xHSB
GXSU7BcfVqvIh8k3dUtpmOXFMIAg+25b4mI6C30HYv38nnZvFkQAEporyDZN
Z0ThLPIcNENlU8HQGwOC02OeLgvvrzmIhRxeCevtTj/g5pSKUJtL7vv6L9/c
iVXzycrLH3XzmJbSCUC4pv+zDLLydkDxvmHfcJIg0meSsuGXw9Lu+E2Iwkb0
Fq1KVE3CFI6faaXy6P8iA7bb//BPJbCInkVVyACh/rtquOkFgNtn5ZGocqHA
+sHET0m0VVgYpjVeDhT52PJaz/ORzLuAoPOulegkUAsy6as3UZrEonSYj2mM
6jR2Okw/Egp8PclUKJSbU/h3LDhIGlzAatfxhVOqin1BZMHpRKrk5EDxg3b6
7Rm8ncC3DaEoIADJsB5nN5CKz6aKoFy8na3tuIYPenTVI0pIRhdZbIbTt+jX
elrUOx5WdLzKymZb/l+ICklfqCcby8ZuUNFvFXmjBcMU1fBePZ2wUDUk44Nf
E6SFXT4rRKrD/RCNop7wjV6ZrW5GRJKxaCTJQGjL29FliLVEvOZVBstOD1ir
DSNJCm6ZbMN9/5tEa7/jQF0+m9+y+8GpWIGqB61PbZjw8ECajWWJAC8U4+FO
wLXy6O/2cwJcgzkWt0vHr0FzxYtLeI+NdrQH7RXMYxc//9mzOjJqXy9lTtMs
111uL/R154MGECHSokvaut16ak/ZvEd73K1eFPvusbg/RxD/2hnp+tZccCpK
ZzRW6FUNTHcePQwuZbVY6hJNs78AA5mOfu5dySXlg0dHMdpDd/gsRvqHPhCZ
nyJ6IfsstxZsO/tXJ+dqHkeESjGYmMQEBtxNTawQaPf/0eKERaKvs8JDtn2T
Q/WD+JiC4KTnvHYLRhiMMZD7LiPPnTdCeiRvB47aNT+iDgkT1BQv6jOAda7p
NxcPInUXdYCk71/Uuat59WBZcF/2tfNXeY6ER9asWzObByXp840XZoUPpx2j
kFKR++NxkVTkURnVFXKuzWys3+mCzWBkfiEfwVlufZX3PUriKbMCufiUS4DT
8LqRyi9IyCXvXlIJSgxZam1QQVMtPlE4VgtJ7Id+6e9P16lBSywwkcagomuC
QNfoWi1UgtUVUQez0gtUtncdDgueqk2j95xdHSqkgEXw1pNH6/EWkxgsrfqB
YgPMbxC3yIpSni9giApnj5V7zF44uYy+rs5NV97cZKtyDHWqwLIqV9LB2Ut0
UPSWSvu0mPeDT5JUpfhh0/RoWFeye02KWPx4JysFLrNuKryxkj0dKXRyVY2V
hhvsZzEJkPqTQC9S2/LN92Gx5cCeTR0/VqXzmg3sJ6tiFx5a8T93VeCMVh9E
pj3NdAvivE0sOzQA6odktWCAtr6caaXbdDxKxC3YQzBPHE+ggptHQo5hKXSl
OxwIegwqT3WQS0ZEKqBP+ye6LFkqY8B0anEzpUltM5SB0wxIwbfGj2HEZmoo
bbSzv8t7BL12PIfmJn4tFnCfPvZ1rsV0bNEOIw3lbisdYN9nJKeEGJrgffPN
jFImbmt8XDsU2Pw/oDw/yKxj7S8NJW8iLyxcOctk4gc/W4DwKVSBLsZGYLOj
qkNuDUNT1009dqJL0XszsC1/Vhn82+BUwL3DyTERm8RsT52QisHk+Ql7rz+X
7INiMKwGckW0Yxw/SdqeGkG0jZYPR68/b/xzP4tAIQ85NUmKKN3d9jhvrg+6
RymRWjy6TfEe2+Bhgd0KHxuF6OwtwadVSZGfe/rQgz7d7gdPsweChn1P2VP1
T331DZWaR2cPJTcAZ4s1zbHxiBwnu/bETrOvSKg8w+/OV4r6VI3dHowivA2O
enMrHFLjKhlf7gveTVYoAFRY8KhuuVHyi/1AGnFW4ZukngWJmDBcmvPx6ODY
9x6rKrTPr+ym7e7DgFypzNI1kNz6A7sRYkbQwIVYHE75gxjx6pFn3mw3pZYB
43hMcfFU9VLA4IxDgAAaG19BirJcPRgo3FRxAGVmFdrD0AvyfZXbsuBRrtCZ
/2dqCtHMruYKIBxtwStAnTNw4PnKcFm+nH6XkspR6yhLA7k3zQnSZ01UdNei
Itput0wOf0WmkjwVbtfxqItFPP7bnM/gd2Iho1dw8IySvy6BC9e2ma6hBGD1
XnTvBTGLJr9idu7l/jdmYBrUuLUQPWgNGDHj/cEOVxD/PZI4jPdpzzkmbR0C
aQXKLpWSkZy4vQ4RhmvbmlgL2KB5P6VFbrD5bRVXnZ/8AFzHqevdnpj0LuFW
cyXLVh9wglpUWqD2/mHd4a8+PrHbR207zq20Rshm8xsmsdY2NBDtUdciMxmz
FMT/t37n+UIcM/IhN4M+XOaz6RGU2dFgriI3496iRINAyQK6n0wijN17GnDT
R5CaNT0A2i9VwwG2wwMhwfFLsq7r4/xp0KyzqWkamP39C8gKd+aPHKjIfMHt
mfVZd5oWvZxLOM1rsODlPS4Pena55zz+pZJ7vPOnM4IgJ8bi122aqS9ACVbo
zcgi+OQBYSjGBHwZIVtUhDry1D2hr7HV2GKA5ugIO1zqiTXOG/JDGt9DJAz/
bLx2DuOsTRdq/lo+mIg/r+ae+K/77Ofx6kvN+aPTDHY1BPt2ZnwNcpMbIq0G
O7ih6uqXyTDOTTr/nUtnTapHpeolCOnbcfkAz+CXPs8k3o/xv+/6XI4q/5Tr
uYY8tv644oDurSeH0eqKw/0OhZmX9tzQ+0TLkyqqdyXBwFbXQGE9A2+OxZjs
Wc06K66HDoPQBFYK1nYm7dQ7XPVV5USkVN0HDpUt32jNBvcMj2JcF104non6
70JrcdYRqB+NF3bwujFZkoigkFVFXHxbvhtiQuki5iiMv/N4/9QR7p8yuciK
RcCrDZvBg1IPu1zXcKtQGYwxsGXZ9djs6PVjvrQqV2G4v7A7SCC0E20Q9Lx+
I40Xi0Up1lfoYPJv7hQh5ADmhjMpEeF2I07caZjtF4Guxo9xzPKjX9OIui+G
jwj1IeycPoZZTC6yWfmvSBhZpSzeXl6XfS20B5yFilHXlS2Lmxm7Gj92H7iR
KN00rqE2PTVmtRvx/jCFBE9LPnx7ZtKIJqW5nCfLyZYQDYGlECCh+2XDyUhl
l3V4SQ/D88NFs/AakJQXohzYpcQni0rPadWm6XK2CMaplclVY4tXNyikqa2z
pDturgA+wRmvw1flQnj1hvKrhcHdIXD6OnvLtMtbRhujxl+xkx1RlH26gg5s
fKfcRpMeJ0OOUkksMaRwXryvQxnHh7W9kKfAtzMOSPY6zX6eXFD9optHRxfX
15Fn7OCzXEnfnfEH4GZgmsYWTe+DNZUHKLxsDMsev+NKpimkDQ1B7VYTQdJv
wylEkm9VXZ2l/s1ijSfSso9r9kkw4e0oG9E3pZ4+umUiftfzc4oHB9IwBrYE
6TA/7mwI5j5W8Tcik7yYuA9aC4JhCAQVSBPSBPtH2gr4F8+hCIW2odZh5joI
Z+cIvlS9Q9TUOObQpbySB5zqh8IsSB3lWGx+diEReC+bsNNKpHFxnxmAw4B0
MN+skVuTAnrb4XhMTBOW7wcc2FXmgu6ab0y+yd74FjpzeSEOOYGN6pm5rA9m
h8wR5AXVY/BAZVAo/aqDsJH+SV77e2K+XlmgDWW3whCJJfb+Ohz7M6YFwTNk
TslFKfCrjfxsNQhe1q97f0gAcgfAyJThGb4xYjYcLjmvLUUyyrnqo4D3vGkN
E8dpPV/C8dqnPAML+ZIxdgnkMXX/aOrXXmTLP6PbvuJIYQP9JGlCAwNhfmKc
m0td6Nn/Q/ZjO0psZhvL7s+cRCLYXXZH2QKHdFF9DdC02mbGfAp+egoJ3k8s
Q1vMAntrreiQTDYP+Wd28GKJ/PmwWIEq0I5bRXzt86CKDCoWaV/Z9kZg1ccA
+rxgWTqI9sidHdK0rBROabT4w44H7Xnzcnk58XurtdTajNmIimXkco/WYWZq
k777lsILt5y9rtrMf+4wfZ87LMgL9f1yO3icbdlN5DKWPvoix5wok29kG690
4vUB57hppd6My/gR8PQxIKPzsDij2FKSOdIInF6h21yWhzidzOX4qohCKka4
LwkebDbV/DTFnjjVWj+BGDn7sKeLy8xn6kOJ6lSURIO+yBO9C6GU2UVcgUeO
fP27+8Wo+J3EMeGeiW6coBEdnhiQ7WPznvDTj/f+QAS13mSOR9hPSyQoQHIu
kj34/tObs1VBXxGRnxo7Ayo3fUGeBug0mIHgqb+Hlq5OJsli3IpyQQFaawnY
XP47QYAmg3eDS+/RuQtxkJasDvsssjGOiapAJTM2NGRg1jeComEmhHSCTR36
+fpahAzfpfxKC77HRSoaUW5bZ+US7h69FAxGQvpm0tQinbyACyYHJ9wdDtEQ
h4P/E9SR25tuMB64hMooYli9KQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "hmRb1hCms2kg5lxwgzvVC1ojkYPyZtVhUZroYIGDp3nv41l/XQfn8gMXcNw31HDDWBFvru7tQ/av+VlNCOY8CAEc3dS4tSN1iCLWoSLzjcf1An3u0nZDKunxPUWY57wMTkfTn6dFEXYBYGQG/cgNqAwhgy/sA9kmZ+yrzAG/xfCgRlDUR3RpN+hQPPycj5HNM2pIgRPAeD/5T2qj/frBFu5c2+SfDL19Hg79cXZFl7V5LRe8OQxEGYeA82EYwmGGH2LsxT3k6GBKluFv/tWB8+DXjYSYIjHAYxVhKHZ5dRa2Q0kxC/+oQ65N0o1UOAHLvAnmpTXJDDGVDJTEtlRNkkfSbqFOERFqr0O5YYo8EJ4AHT3M73izQVa3xqsdvzJmHa4AbFaA81cSJIoQoX/aOMmTylbJup47LS/hfC2GyAuHUH6RdT/FrcqHRwr3Cxc4JjC7ZeBcc6GcK4mXa8hOklIzLr1C2OCjCJLRKG22cTMnGIG/WoCPoAALqvPyrJdWLmT+kf4MmVjQh9Ez4Ao16qsoN9EZY+ymj6DlxZIljTRoqrzyFYiPgJbCjuUwloQlZrw+aqWS6FOXezfm1bZjdRZm9r4ak733YIaz+RURFjVeGy3wEw1Lz7u6DzbGwlwIay2z34KHKdO4VWaWvuuKM78/QYADdXBhfU7VRhiccKI4CvqhauyG/KvS9qqtXjdPjKcwgekj6q+VvlM0vwqoXKMK9vGqvdWaGMFiNzihLnw5/XzApp2WV+54eOUTSXmmFCS4/rOSC0AtwvwJTFRgPMiGyMiAlu4oX2lNbYz7PvBCcjuPZrRhMXMueTsiB0uc2flerbjhRKN5fm9NHOuiYlAY1gplKixhu9EQYIgQYAVd7hy/ARSS67kGgzjOcBkudVl9UdQFkv628oy1M+CdtyoYj7yikzY86mN4zNSFhThl+19ihTKcPgAoWBOigyUPvh23zREMx7a5FjiLXuxPpPftHZYgw7Si9gtm28r/4NNPIn57rGkYMVz/rmREuJOq"
`endif