// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xHW6lhB8jSocx3l7SDPM+exGLQ9ZUDyGteCcQALWR12yAq3zP1NlE2BU4dTk
yFucaoxQPXduKGpS9aAkghLqdjNSNu9MjwatAbitWCGJFAER1qrzwZ7zB5Ld
L2e//aFduR12OqogcXfGfnJxBzzmPZ7B4/Lu6gVsRP6mmp1+jhXkKRSxxrUy
7YX0iSkCC7DjKzT7hYUkJtNX5w8Rzh9htEXbpfPJawfmgcbjgu0bP040t/uf
fefj/9URhVSMao/8pJszydBUwupersy24pJhIWVCbQ+BbCoIM8NttePSELi6
vErn0578CzrR2DSV2+1aVCFhqHbcsLadV00S6ley9g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mmOk+s98j4zClUr7O2TIZSkXzGIZ05BS7S98Xjasy1VfZmVkQh4CCtVkzOoF
VvL6cCefzkU25uC9OOnAj8Gd9d+a/1OmWWj44ToZp2/ts9Geb6YEFLCw/jOg
Fez8WfICpD7HeT0Qwqh/LqnqbRuA5K5zKjxPFRiIujcSTnZM2Axodq+7tC01
HT+QXKotd4PhZdVMkenWC9H7o0X4LwCo0LJ7dQTywBbQ1fva5J1JRlEz7+VF
1qLvtLKeoUhum8roLWguFzG2+2SYK3njCpLTim/vvDHtWa6pd2/y7AVsR5YN
kAm5072pkRsFD+5Sjj6TtW0P9rU1de//Bdn+bBhhVQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BQlaUMi9Cfl157NRrVx5v0nwR7Kwnis/9iefrS58VnpSuXYOnLA95MjtKhgk
gZ8u6/SJnpUOt6i+uvjCJxJnC8DUqF3rdWc259nvokAGW2D6SfSoU/Gwyqdg
rtSFw2oQ09ukxWG7EpJS51fDRP4Bl2W4UlhGiSTJAKXNmTVOhM0SrqlXXMyy
79JjDic7D6O5JKaQbnXNI36VftufhDgPTQdwhDglK3irB7QWpPOM7MUv0fB9
s6YowwGwNkDw3/Y3vPLZoia/Q48Y3n5fV2aODtR5h2EHTqVNU0DqwFojpCKi
zAy2q69xgVKOxGlr+nwQSKUbLrFnqvBzP07x2YyPDw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YAfvquRMJdHbgW6GJYa3XvVNLGCBRCc0Ok3i+Cx9nwXT4KhvgHJdScui5jgj
1EWUaey1ybxmFeFb0NNY8o9CPdw8TTJgQtUxzCk4hdNcjwSdsrk5UHZQKGcB
QG/AREq8jiJ3A6znr3or7A/bF8+SjfWlI6XeUhy+wBvceqYCVxybnsLVcoJB
jn/yfV81prQisDFTmtrLsew8/pi5b7Hb+N8y17F0K+jM2PeIs1WjBaVQ34I9
DVQd3MXhj62dn5ufxdAg/Ow8EHxiwTHlMChwMPSDFJenDzJbL9I0kS62tgvi
JTIBV/Vqd2dp90q3hyfsyHCXBC7LKkOGL9CNn6Kc4A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CnKmChogYZHbqMVpwbFaZdksBOqyptuxyQp4nAmAyKLcdXanNRtAVfd9Fg3U
NvGaPva6yamnWeGP+AyP8MsyomMz3xUyhLs4RzehIw7Jma8GkUTTzRuoOcbd
zlyeSbXpXkxNOVALD6xYfdXiIiVzmrq4HaiFMv7+8snlatare60=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
I7zqePRQrNmRwybBfmjjMRuXoCdkmxxAdn4OisNKNWT/zINXmKUEINTY5nAN
0u9xAfruj3UTjjchqgiopiZC5/ZHgsAe+mrRCB+Huqk6eKY0i9G7uJbieP0p
pX2juTWhUlTHha6dKkldOKJkmu2j4ac0SYB6gXctg1Lhz3TjlRzQijwwZJHs
AD20108NfpokwZdGBqiTNyhAfdBAq+KWZDryralUNHJzwKXPmLB1mqa26PQT
KavKYXDdLzuFv8QXjzCqViBBj8XgMIbehP3q1R28VY81s2N2jGPdPp2e/NQQ
kVqi4A23ydAns0VP7X7x/FdNMDR1VQMU4mYFHA+sAbKkg6U0a/zsiHusfqzI
i1Npw1lG2jbmmaAIYUlTsbXxM+Xfp3y/ydo6hzjvyHqxpX68H9OVsBNQBmix
RdN0nIsIu71LqaTTDiDY9iVSxQTZSDkX4aCfrAFwK2bJfQV41HmohyGt50y2
Sk/42dq9XMNKoxGf5CGeelJQiIy5CaJv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
abZOn71I/pp4GQo5HNKlP0mNLQx5VZFqh18HU0tZ4z3Ro0Hg9xAGxhjhQITT
/LTMjbw1AqJhY1G8sgoPfKBpqWCCh/40VvrEmCnT1NTwOoVThdmbNyvCwli1
q/V0eEbN4mlRWETsGKa4ak/A8XCwvJgTnULQyErd91nfh2G3D5E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Dx5NXpAikZJR8JJS9+4GQvJR8QnOj6xdH3uwj5xDtwWeuFezJYXgKPw8IWIl
ZeHM/7GFmZnkp0/Dd7s0yYzAtdJMRWMgO8MqxCvYqN5v6W3uMkYlZUEyNUNO
VUmqMKPM0WDJ52MZJOCwYDxtUjRjH+zTtTKA9lzEVFgLPZvIE68=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8272)
`pragma protect data_block
VPJprUQCy/wiM8FVBZVNV1PrQ5OxtiEsUs+ftadx0gwCf50WMMaZw7ya3ddT
Dm1GxjRKqPb+wO6qDOqkPNBrAeiAbKzTqTV8hfVUuIrz6dHyi/Rj3rbQ5ET2
NScs3BahXZf8NebWULf9S2R87YJaTybDNfLC4ZQWbcTvjY9wlki3sZfpKNZ5
zA+GIuhE1alJ69VCOIWKxP3aIlSt3n0ZVlesqVxBDtC/paav+ObO1FoFYenU
1aBnXLgx+QRcfp/3cXJ3vR7phcQSEMOBAqvDXjXvUV980EkCCePb+6pbx5Ne
Xtn0uj8/K5nDVPqQRKKPZxavXE/2ZJ0huMk7PWMaG67c+IeJGcrPtXQt4Nm5
r/ZR/+F86D2l02Iy50tKPush48ghtjjWxb6jqYYs/KeoNiSbuWM7w981R/uh
z3bt3l11mN3tObjoYE2mDu7gInq6EZ7vndgj4FggRizZvt/hNGl8bhG1lG39
RF12YFUP38aOzcEOsR7ExDmffQrTli/dxLm1ri3k9ma0vGlFBZMUx9aCywSk
20fy02mun4Tju9iRgboHXyPtX5+ytIYkuE1Zyvu8Sl+gf4/+Npstg0f5RKaj
IwWJ9n7r7pEpdn+9AGAB9E7cBawMLMESHX5/6/9NEke6eJEt9yfk6VbETauu
Vk/EbxN7TVbYui53svLHKk3Y351pln6jpTVcq4xxbhwRus140tcvxtlNME0E
2dWmCOdXnpR+NJiM6jlUYTnXAjoBnoAnK8y1Fl7dciYVa22AHZoyVcXCdlHP
CdK+GX6Q5lwIp6l/FkX86nXaqdGepRN0PP6V29huafJj9ugWS9So1j8qYyhV
W8smc1xRw/hyOCwecEoRxWZJWVyAuAadVo20RHwHyef+oztKp+/egabZ4jSY
CIQIH6kIkIoHTeKlsp/Z3TmZ/ya9YWD++4cR86iFkAOZ524sxxsDOnvBxmJY
XCxAh1zPIGtgVg7y0p4c/cZhmu/o3r02QEvKponWzhZCDrfjBQQlEpsJliGH
bLrs7ROEWZouKUy2+DPMdSnkP7+W5VbVpeYFtz5CR685DeVgDEIxLxvRJQB6
PQd0r8a5C3IQl8+m/lVSfjSsydwcV1nHOVJ5en1Lh+Oeg9KUafbHZecO5g/U
+WTs8LqZwQX83Ll4oo7KGJhwQLYMdeJFVEw/i21V4k18CSEODAGzg8/QOMUj
bS3c7C/mDla4/UtjMQSv2WpaGknBfda0WnyQCEDAiwnC8lmEIWxSl0DbJ74Y
ei0zU5/ts7QPQP4ydxeN5EbRVZYcBL2cXfRNSW9YZ7oGq/qhqk7O2FvFiVDt
pC5Xq4kUlkVdV5XsSs/2aZlKszsijlSud2oWTOADSap8CRh85M0aThSjGVsM
ldnCxf1hn2l/zCaT8CnSXRvOSyQA5fBFaXw1FvtnpWclzr5tmRxTeehYv7OU
Tj95oxF2DimJ5NVaFbIXwP1Stvh2gfhtKUOYmlNUkNEXzrXyBfy/sxaErq69
0Z+OJgKpJqkKyN9PE1hdfbT7DoYUV7wlnKK6gsB8uM3PS9GqG5X5LsmakFEI
BPj2V4/06hRz5W881g4rD+fsAbbvYtEOPA/qmoDOeJ5HTTDURWu1EbTct11i
1lx8g/UjFshARq93V7+PpilHQZ/Ru+W+Qe4VcBu9BQoYv8KYXwP/uzQ11HO3
e5M/nbGitTQCLmFNnYrVP33XT+LUmzP7ESL30w7HyMpRuexM5t9qjLacZAom
B3CQu/GPGi5ZFR+JIGxJ69WD62kWKu7CdM1ubiaZrriY4+APyENwv/iC9tMW
9qEQQVMRjzzw5ezoKUoKV+IMS26vnllpPiyCDfobKnD4GWfGiaGvWT405C7G
ZcG2jM5NpXKyHoCnp1mNK/2s+7T4Um75/61Md5xz0TZ9z8mkS28SwvigQu87
5ZeK4N7VajLA273KJVjH3UVExH/TLcjnDoRFlsb7fc2YHxxKCoGGbfl0leO3
T0haWzk9wURxaRbF2lzHJKY8zbwMSlq2n3UPa93hpYKbR8VcJybfr8L63UnT
1wEEqHRDoO+kgngrHyFCZIHU4P4zvXUQ3SThHuxTOyXF4TauwHvTtf9BjKBS
YPOLNpeOsATBchB5dsWVqkJkFvxcKTQNzxjKrX9qAngb8ND7Kr1QCJoN87qG
1jCfzg9RlTQxaPe3QNE7C4sCG5wo70hTtgdxskAmzoHEQdsAvHPkxIVJb1YB
hBKZqTbCQyPfp2xzXwxhxcPeFjSqJyS0M9XcLHN7/eVjG1a0y4ZglS43q+uY
QeYJFx+nscOvCD8GmJKZgp/sCrOmgjlVqacuRmrKHqywHTrpz+iniaZMcpuC
ZNbHv3t8NJ/uCMdHsRV3pTtBMsSagCoalnOMCSbogseANSMndwtNfLONCBOi
0fzfdvxWa8EMC7kRmuQU4q9zycHU/XqibSIp5WuP+IHal1GoVzEnaT1hhJQX
jUI4qwpXUViv47T/oSV6P4q38DGwfF1lHjnKo8nT/rnY5gtjkyiqx7OCdiBA
tzb+Y8ns3eWsMH6wKNxAy6fkpZYfv3N7Ta2/swSxQ1IBHe4bbHvG1OC5COwm
afUh2xQA96IbwpeTfLmjqk/W5HQiyaBkRavThOmpvNtN9rKJd4zk3w8YxGyQ
wBlfBPh4lyr+SfEx1lP2mqJf8qKQrCjwLp1gIiBymG0iVesFt/OcrVbb06t2
JM4jYLzfkwyKA80j5mOxgM74k+Vk3SMjt7wAoPilREw0p33w2Efj+lxyAKSd
wuv0YCbNqLkofhH7PIW0ql45k85Bn3BUyQESbyvInXeSwc16M+BU3fQBEZnB
ahtYkOi4AWh4b5MLZASlSwr578MJNt5TuP502Wu2t+l80cUf2gOc2jIt/MHn
Oka54JF12cwGVLt3wJF6AibYlQNaWOCBwE5yh0nDJHEjMXsaIv5TrA7MmxsJ
JG5BZa5pJOesLXxBvKxnByTXA9n1TUrpF/kVKyTI267M5KKYntYHnfJsUpxl
0DOxrcVS8TgiugyE7h2V14dlCDNKbCLuhlNCLe6dtuf4oRZFrKWC2pN36aL7
TVOjJFscglcEGEGxxgHLoX35Z3l2HvzQih9wp/n4V7Eii8cA8A24UcoZl+b+
JqpxWA1XT3iuNK7TXSDiT2dYUJGeG9AxbS/G0ot9ZY0a28aGzQIZrcK2LPa9
RX/Q9SUqXUTZs9DTrfa+RUELFBzMyNv8QiwJhNgoq7bjnoNUIqM88wBUdz98
mTqnwoSb2GNCnst7fvzQFeXuR+Fe3uN1XhuW2UZZXXprNMBRqdx7WVmBICJr
qbJqeKE5DBEDP9KZk2wrfZ9t/K+5ohNEUZrHtBwyFbw/qWI93ph3Z8K0kzLO
W4kbpZ+uRIk67WwoH75al6y2Km7ho6kjGQCGga5LM2fkSdLaGW9kkooobhMe
+ilXtEJ+STPyVyGLjyPSUyoozOHIPatODTWTvlaaFo6K1NuxMIc4atHvJ+R6
AH9L2dxj68ADognu9rajkM4QN/sTUM6zkRblU+bYu17FWcv0MsWUdFmQHgbq
Xabl1SWL7iXsXG+sxPltKprsVWRS3G2LW7UOaKyGyDXLZE05EeKtEaGABdGj
CBKAzX6khDZUfhal6a/c6oK43ozlAS5KOcVKkv0SeWSPDsyvsgS8IK0WTeMD
ggx5Sgkpcma4yEwfhAJ+qtEJE+hdTS2PSWRQgt87fdQGLEV4moTaE5srfKKA
KBI9KRlAnkuQ/YtasY+k4up5Duo4mW1e9vmXKPf8XubL3+60+cNPRg+pohIh
2op3xm0RcZaJcGC2M9vP4tRulTh+ZBn3g7UFFoZSxrU4XNwpR+nI85SfMEUn
C8rGebtrlxRqLSbdEbqaRYRMCoNe50aPqvuD8pQAiOHLCbXch5PiC8hcy2EI
diif8VnicyshQ/zrkRWcxS35T62ltB5QXak01knJnhS2z3equTFuDTZJ4FbT
zTZ6Sgx/yqlnF5hAvZUvi4m7d8N648jU1PO8udzBmAfVdyqaPWBDHV92Ccj6
J4seprTMOQO1Eu0WJaUKDvY6Zi7ROo9aFJFPC2a326cBRBnLdCL1/WEHYIuj
y7JoXCT9JtwFE5aRkzKapi3SLYnWIFiJNZMnkre6DxQbGb9Naa4GG5INJP3G
1MCMOemtwtXGy5fRtSPb50t3sBpyxgSA2Aty6+pBaz1Mxxa5MprZvgIZFyVu
ucu5vl6ei+Zqxux/ovxZgUOLFyIqiXHmfzCMgUgoa2X03G5jyquJgqI1KTU8
1TvcWP4rivv5HVKEfPb01gNCVZrRS2PXwsnd0koxhD8zANpqLbk36TNUKDhM
YscsummUGs9lH6cM4C5prkSF+/gqr6dDk4+u3/6Kh6K6OlNp1djcwTifjPOG
pW0wmq3Vzy7inyOWSIcPkhJTO4F2pRKgWtufbWhCCKPX0NPwJ6sMQVHyd3JN
tPW6VEq3CFVDXDxh01mdVmUtgTcbVrQUc2ljCHfGbvDm3cR3bgCjm1nPyveC
PU96ZGI522L2yVz6dQdbzxeQktfn4xA+FvUVEYWYR8t2Uj9GQCho28vkYBwH
JAwAp4lUVu+5j1gL8LCnhFyRGFVeWVQ+aAgaw0WvlryBpZH1FGl/LRTnhUPp
PyHoFyzqPm/aC3eZWrVaUh3OKGJtzVoroojLhnTjHkcKP72Hoq5X71BlTEen
TqopxsVagDPEzohz11kqPyCChq+EeSxoFmv9eKriF8e+r3jr8RjlVhgp6Dom
Hu46Mhyr/vTAYK+Ou3v0eWrhFsO1FzO9AjpdidHUCkNz8oPtGkkGERT9I4DP
zX3h3aaI8ioPEZh2vlhFg4ViEfyFBZGJlZR8xdDtosxNI8lY3cm+97TC6BVb
8XItQ3ZF+/mjoj3OPM/loTBqABOdGQSv3ehBDvMAfRLhbemeY8WmIoPHRz+r
rnwKfN3t3Ob0hY65mKX+oVfcr3/bWTcpy0wj2W/b7roge5R3nV7v5KjegoyP
uklUqQA/isSfygQepm4Lr/i9zhvgsRyImDo4EHR2kWKu9C5rQtuYuTK2BGz2
QnExVjsONtJnnkRKLatTKQwTRyefoi8IF7oaBulT55nDZ32HA6a7Tfpn124f
8HQVglZ/eXfKdxVHYxSiCUXX/QN5He5oz2MF2gvJxph9wnRd9FbZ7C3hv9Le
qqixXbQtO+NTrb4wLaMof5X/E6jN315fMwfw8yWeN0NUe+2N51/3/zSU5i7W
SzEIKWbu1LXBRegP9lglFPrZNA9tMyxJguO9GV6JZDyMBJ7k+hWK9IDGS6nH
hw/llpfl7ot2RFMkgLsM24pc8s9miyPnLp28OtOh1vWuuKJbfrH+zcCKgtJL
rbEw7VRDvEqT32i4KyDrm6+yvvPPG01flseRwt5CkYk9XqQYsfZ1lM35WySw
Qj9VgCHgWtiVebuD4ENhmQ2/M6baZRDsMRA4Hp9uXsy8Uf6hgW2czowMnH3N
YGataSH9FY9fitdl3NuueifvDJfYsf7FHOJPDIVsIUCLxiN+ptIh80VduJaa
yugehM+xDrKD+yVno4vRm5cdF0wnPdVW5nkTb5VMA30Qi91Twd0oM35/CqDn
TYs82AYEF/xR0Hze+bG38bgCuGe5CiLA4XRG2GUVZRfNKbSctCrosz88t+yz
3hp4BwK0StZeq1lPgXHyDa6ABC/DBLJhMi+YwftdmPVkyAt4/nruZvLMrsEb
0fzUuCHybL7BYI5VYfjRCE8XlXC2U5I/KDnlG9c2CHcvPz7XHEDfX6HepgXz
BoOFra/1b9h0QPAN99/f9HsklUO07I5Ll+O104rtmzZOAdsvP0t9xEw96Ykt
OmWTuX7xCUXlXNdgF3rViuw73hJJoTKDN+/555XynLNNtrOlMzR5lPzVsCpM
Oei9TjDDhAN13eXspSao2JCkHaCUGYvN1WBv0AfE9Pg/wiX5ClzVH71ggdU6
/pbefdtjFiHArzbD8SRZQlBah/1Gj3nFXAsXKNZI7OAN4VqOWKmWmr/S4897
zs/mjInV4EbSLWCbJajCJ6ehg29SIcl1yRQeHOh7NKLoRI0pOiHpFhGuDaHF
f0DhaZUcZBGnj5NI1Ulwmk65Pk2xXetnBir3l88xZNJSpZysbo/Ri/N+bv9x
Mqjjb4auXK5YspHx3p0Arv9h8oucw6K21wRtWybBK+9ABohgsVvn+h5IhRob
KxucG4TZm6EDkjQM164DadlAZL2MsRQrJ2nbdNBCYJSfeSEFj3GneDN5kGno
2W55IbOxcsK6djH+EElCCoBFyeFvNic7OanZ9Qv5DAxasDeVt2brxIYyvJDM
FmXzEaH/1tBKie1qka2ZtdL+wvEUvc9JIiOxFJNr8JUeBAm//Wvx/4EULTWx
9vk5X4F7xVzexiG62qULc/htC+RPUAgaFy9xyKtFLRaLUwuhu83KktMARv0l
5FoUhTlej8hX+zc7EXZgQDe7y1ygp2gXCdCgLNwzke0CmB9RyWNOyeAaeas5
lcacBQXxvcs1uJ5Pr68AHDJcsdDfjcNsiVy02PqPnRmBkNvLuQUtHYF9GdSo
UUeVwNBPUemtI83iUhzyErF5aXJARRiXxUNCrf1cZ9GWijec56/v7E4zWqWL
CNEMGC68RGu17LaIBpoSA1c/44raiVtg4iNc6oYcRDW158K4CQbG4f5CXRwt
RzYEkqNsRp4L13gjkd/ZgQ+C5vGyvOdQbH2WO9dgKutAnKdt9HsNVmUCViU+
YxIgD+AeC74LSneVHM3FQdjznKpg7m5oPMWjbUsKhuieRLFXYelnxD64syKh
P0mQbZ3yZIkwuIvTjqh8drNP0EjjKTT+0uqu1Zb8cIdyg5OyPIuPfHXooGJ9
adF9s/AIacj4p2iNaLPag/my2fxg+TxE+D0SMoCZICa1V9BNWlVF3TS+9OZi
Z/e3qqvGiP6A85xw+/4ve74LOKnlp3an/RpTZVH8ODY2TKKsIAa6DmzqI0r+
H2oBze/rlB0M0XKXkHPqx7EzqdwnGMEmpIfIsG264YbxKl8crkGbt4i3cB6j
dOcY7gbfbuCvrgVS7JsKxDl56utbGIJXhwWnWCJn7bjFza6N6z1Un/XAxPPC
dgT0XvlYI4nbKG4eJaAphH0E/ZlJROY3ugxK6SrdebCaYT7zq/X6XPiQ8xPs
C5a/+QbIzbmnwF/x259qNMViBeStqHFFHHYHyrw8ueu+3WHCj+Yb36cGhii6
kroEorLOkkEcuSl7A0a8BGkJJR8tVTwzg6+Dd5Yg20523f++q3iWisi2Aoe1
xvaMPGwucESGP6Ya9bMeNQmneRGAdorkI1UYR6YwALm8Z5hHM93+Ogd33CJb
NB05Y2U23Iu41ikgU9rCgoECQgjZsj+wA7eun4q5TetZmltaJNT0J5lkaF0/
yt49U08omEegrx/XvJlVjoeKXG3AfHgNDx5FJWHIu9MavrffdG/ge0Q0Hk4Y
d2nfyun+4XcUGeNjCGBgYdIljUqNz5U2G1kZ6tFMqU8tFurUKPgYteFuxnLE
Q4GgkZ6tox7yiUkMDW3PJDzlULoX92BGH+d2dkzi0BSJX0HEg4lkp0DxdAHO
ReUZwNqvJ65jjFzwJR2zf+0wzgGp6fL9nRk0AUXtLSZJw40FMv6qMMFSvXc9
lRzVrHkOljNthEVfUgv2d+6aYiBvaL198DXQcTQ/NvG9Qr6DTQH62Sptz9tT
e7QJ8pJYEzP4fYBqMr9VLUDTblbU5rbz7sNgtN1UwQ60nEo6XthiDRs8jA4m
WlwOBnz142p/BJo6TB9VXGWuVxT5yaM2pABZxrOwjTIaHcHjGowwbHOGxSUE
uHjIGvSlLq2J3tjnaBu4azuTDqqXqkJ85wFy0R5oB6/WWom/c4+kyJim7tFY
WecK/xTbnA4iD/AWQhtOacVkX9jwDB89xEVya9SZBLnnf+G8Mu+PolYemu/U
r5KobatPlOHf+dfOb/q1v3c8xfPeXwvgI4cAIfcikh4ByOEXqhyu1mgZ797B
6HTdj/rqFFd04PPNiiRITmoH+AaFe8SI3v1PKwF6BW3bumyW2Isoj+ftoPb2
srM+k55BKs5MQJ6jJJirfQhkqARRixVtL4bBQ0r26qR8tc0YYl1p8H39laJT
9T8IRqHHEK7o+OZkc4W5AAqzpULItsxw44pBsNzQugvpmmhdRpYAurQI86ru
WvT4PYd/ezRCWnYEjbjn3ZsAAuzOFU/uJY4ReYwFidi7TczMuc7YMH2HRkmX
i+JalYWGLKq6MwO2A/cEJF+rKm2TqFNq+6Oxx+ncPvhNVY00FPzkTAgPz5r9
xyD3JhHhJfqZhzUrGzsruxWNTlX5QZoB+G2H+Yaw1nRau+1+gtPBtUy0H0yB
DSdCiVQ6qt4Vu0Q2C4QB9VjdeikawWqgyx2GkYwG0EWoKEqbvaU9Aots09Ke
YXjjEbZCKq1KYdDssHHLX+NAPgJAh46R9keK3u2LCvxK6KEVme9sRlInBIp3
NTbr00Uo2mE3bR6Bnt0zsTVAHKUQQVt7UBZaZl8T0uRW0E1KVsjKHPpx5NYL
ZZbcwkvhlyKAf3nujXDmDMCUWa4o5O/24/I7hASOMDBWIHvtAwCh7cL39CtB
85JM4T6LKBlVQWeBrrRF9oFpi63XRdGk2qBpHrC7QVnkL/JFb44rejrYsZ3W
mzhJintbeFm3kfdHw8fJjPBgQhb4EDTYkf7+Rfktrdj3nI3mwi5LCY5tH8xt
ZWvkunWH3l3iWpRezTYpC5Y0cyYQsOcT70Ymtu/8IoMS1L4ZIF7qIHP3sb9S
vd7z4TZKM7pr1c5gVCyheC258ogBejOHKf20ewvT8Jhw3A5Yr1dSmohlcfni
zLDLfD/+02GUT1sIbb4VKywsbzZNpm7V0bt5tE8NzAqiB7dh/cLgwpP1IHsR
7p61vd/Lx+0C5yZ2KN0ryMsh3biH9yBDwGbohvYg5DypI9YVQb2Du+PHb2oc
Bj9aV0a2Wemq93ELP8NvI1khfrTNdgL0jOWdubMfgEmQRXa+Gd6a7uPQXNku
HcRPdu2Fc2EyHrhcNrR1N9NQTxzHXu1jyxkJ0CwyCh9CObdDp6g4J64aoOeI
0tAHi3AM5v2qpKUUV6jNIFByFi8qDUDra69G/HI6t/vW6Z+CiCGrBSzcEdM+
gX+zbq/cftWX1KSqIfeYUey5tdV5MDYb4H5IYn8uRLn2PZwntkEBcCje2Bgc
PPoAOS0P0UVDzIZrN/s3uvumVuvtToXgyBBRX8NqIxu8wZI8FYlIyHh0iZR6
5WwUaTF3YIPxfrPhn7bw1OWQgJhYhRn1sgIZopNx7y7la3fGkFIsAaGRjiyG
si+QRLL3Y8NGoqSacPYlBLPhKsIwdEQbjRXW9dFleQOxInhdRhtZsOOrtBnh
kyHMi1xj/cHUy3seydQD/fTDxQFI0O3+rxzYxKqgGX2xJYbrf4+5yfwNF95z
PSiqyHBMUjVVnynVnhVa3WcBHjH9MLN+cw6ly97cpRhXZ3OuzM8LZB91jWHv
9W5z7EBi75baebSFnu6107ypFbGw4ow1gqtjNVEFIAewm6b9G7mnwX+hx9S6
S9udBHzdmE+ll8wuAuRzjLk2aUd+fqhA0NWx8+ZMLYeL6jXrKrBALN0BSBw+
GO0gH/R2fNxAn3OSkDbPSl+f4EVCB4dc7+F/k1MCO09f630jmfOfwUhbjGXL
Sl5FH1tHetwz0jqKyoYXdSmOAX20jKy2snV1e4QzrPgZ7u+t5Tt68MPz8l/2
qDKv6lV3Q0dj4qXLbZKdwIhJLdeE23OZlV5uDvcxSCGRFCOzZavg4IBPT6Yy
27m+6Tt8Tt8Drn6veu+/rxSOSCRw1dqQn9/2sKCK8CdzgceQAkH1V++wvTs8
poKB9MQ+Jj7va5E5qJV0qdyrVRlXE/QUuMxxAaTiv4AKv1z5Z3indMcKYqqG
Irigq6t6GTOF35xqZf6CY7ZsVyoYHntT6y2PhZ93z7MyevcaLfA+8mmUKcsP
YYKI8M/ghmCX76bTDYqXdkJlNZHOzjr3G7EoI+UL0V+hYbr1pNNjHWX6rvXm
ZSkAtTat6bGmfegVJ5LLwrdpP1/r+dVd1yT4v9dEdCljcCdMn84sytoT96l5
OOlbwAqUUTbGMC4ctoOSVmk+xSpdR6wcn0lxQXPSiy0XGGVt9UGQbc/SLLTV
akKanW2daSFUCrwzVsNue2cvoXCz54Qtf17Ujk0StA+84RW9CNVTB5A8dvdP
PY4+cHq/0eWTi8UzKbURgRKpLz6xVrC4b66WzC9RJ3wRWr+JyuN7cNtxVk94
qBZVkkUO4B7ICmBsMCFp385bzz/Nh10rNKdJLMKMkDV+QioSMHKFG4RpQakD
f0FebQR9W9nNOIKccrPx7O13BSTtfvaPGK/LMFBNrckJn3kge4t4yYgUYfVX
UA3YO7mpqOUIT525Ul39Z5rheUEOKFkJrQqMJjv01abSgW9InBrvaXlNCbdP
tENchMFceD8M8TVYTfJK7LaUb9mGikLW7mX+JfwPiG1Jwk9xQh6oBoVspyb4
SNzLTsIR++RWVOAyVTMpf7ztOSr5mJ8KGkNGKFZkJduQblrPauWCCcYnQZnN
x2BC2klnm5C00eBjTaSEhAHhFpOPGpzDmrc9Qwb5VImsMBCB4U+Iyuhy9Pw7
QcO/DC9GvduQAwUQzyfMcgSFbcqbbnhqR3xFX+UoikC1U3AdfaK5+ALOovm6
Q+HjsjAzPhe2dT89kG9A3ItkReyT+ghP7aXgqh2lEdMsoLxiHag51NNFIr1a
26zzOvphODMN3qIxHCy0KqUyq1vkE/TsKoVJ9uiPQf2yxMTI52e3PyBF/rOt
O/3k5p1feEXtgPghYwJ5389OMbmPfftmMzbL7Kskz0uPd7aR1NFxpYCl8g1I
VpyjY30Ry3SeEjCOM0JP4YZ6oGe5QpWLddFZ5qo9zkfaam11TfFTEdXv6Cta
hYpL2ucdbB3v7u5luxYMwRKtHGYxUSvo+0rvAeTiwRJPV3n75JHon2YuUenn
EptX9UUw+ITPayf83wurkOiyeVLlv/QdncXtr5LwGICaWsZi0w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGPWWPwC5++HygFGnRKRpLGL5thpM+U13sxAPd8CcD+HojU9kx1FKLV3suwbhdLF+q/F9gx62FG1m0pyiBqNHvvZgjW7Fz2ilexXlDhb6IN4q9aJenfdQdXDw+odyv10JcLo9X2/b/vnWxD9QctPNgdcQS6uhzCVwzqJYJ/0pC1NQKgGWiZt5w9mKYYxJc2/0bTt1EUnpq12lyifrODdXolOIBAiU7DSMYatTSVsHNFsVYIDCb+Qzyq1nIfV6FoNTrxZeGhnkPzcRW+CzhMbz0mIWQETUhgireEn61XXD76JH58VPZH+8dtp8XaEIhzpboMzQyZ881Ds7YFCcev8f7I+JP7a3UAEy5H3yfzg2LattBsWDpoDoZ92EnFYo9qNy+/Fuh4m88sCSDvXhtudm9BTWMTyVR3/2qfEc18wMYI6sa5yBaRZ/6hT3r0rtbRstbcbJbwXw6F8bSM2DI5Ej4rIERdvdMfXV+07rr46OxQmnUtkt1mswC2CfwdksvWeixuxcTZDsifH5vYDmUXC1HBCwzYV6EU3/FvMk7tQxSvGqfFmzRqXbSy4LzSxJWfa1It76BOgECyc6bk2rAb6o+FqhdgbcSnAC1Ck85U/LSNNpe8reM5ik2cLqo6+ZKjc1FIOirKsItxFEVFzJtsA5jftEwBEoRkOH8svvN06mw0gnTjBFqe80jiDlyidBijnsQpQBjOtEBDxeuPmGCCswOfPMlOWTA7I9R3McNMimrsuFjQU+lspfzTmYiAQPhGiTanr00WlSVkNeaU0p2ShdCAJ"
`endif