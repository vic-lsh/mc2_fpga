// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BzfkDLHnE+CYcvLQjpChPK+jaELKYV2+QBrzJcrnqFhmWtKr+ds73YjZDdDS
xfjVa/7+NMGer1P2ppWk51k1sf32y/tVdoSD3N2K6QpNWYaukwkhRZwhxQOG
G8iyjw4a/Qow81DKxJ7JRA8AO0mQtGukxEADWbZamRSMQHIHnaVFeJgJTG5l
GyCK2yMFsVYazMgE0rHvjfBNJlAMAwav1LbvO0Xqk4khwcUFfL2AUC0CRZxE
L6kMQnvVSolXk5bCGb5olXh/jwXRt9WT6amHD7ov/71fF4DLt+GZ3NUhW8wD
WC+YgtKDIUA/vR+UCfVOvaHYOhM4D1kPEKgCQVM89Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DhvMzwaVh/gdp1+FyNGQzTAYZ9jZ+fJ+WKhEoQmw8/3gMP/m4zvjU+erb5SG
aFNKUR0gxa2RLQJazPIHtYAn39DO2NycXhkyVfgWyM8BNFDiF+1zJYb1tOPG
313ziGzY7N0PdLzJG07CFOePyAys9vjg/xBDNb5nZVehA+RI6VtSjkMokFT6
bI3WBh90Z1Adctck8rmM0EI59QwlEH+6XqXhC4DXnLxTsuzyinRLs9CSQShg
MM2xMcVB3fjWNbb7SGV+m8++Zdgk9G1ouSyG9u2bOxBeglpp/QETrOZIiZbr
MQ7o2Ky4k1UJX3GSccUn74+vhnlycoz8d1gnKUDTlg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HFXVO+nYFQ0NOwuHY1qi/2Fdj7TnO5u/Z4irv0SEWDdtCpkTfJxV5Rrbvxkb
/9cy2mn95Zwrh61+atcwxMFGWFLmxmaDNOKzvzuHnN/ciAlNXCJ0X8CaUcbZ
MG6iZZSIZDvzBVSuXMhTWVSwiKs2h1TQAe6XJbwkIgEbST9j1JjBD5Vox5qZ
FOVNdwDbyIzVvr04iYj3sAUfaQDklRX+amwtL5Ol3JcD32TecWOWImE0FaU1
bUaDds+tApwNI60+MnMbuBmS6DMuKzoD+FhHLOlLS9Yl1AGTdX52bvQTGZw0
K6AcwoKN2rLzFpWWWHq4KcFmEg483aQobGdJMCsD7g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JtCjtOCoeBHwaE9TFTWlBLU7I3JFp0V0XsF9EyMZi5apgRcnlk9ZqM+fHclV
2KYdOuwkrZWuaLfkNV/xMWp6yf+EzxX0acgQUWnr08db5ADUgRaaz/8bE3Re
i5uSZKJDLLogkZ9cLJUMBPB6lpawYkUXBycniLvcxwWL9akU+EnH5Hbhw9Ua
MZlXfRBD5VbL4kNyVTOUYZCvmgLKUPB5EUDCFNoT1Hz8z8JhrRycFx3Gpu5L
sx51Jskk6ltDJ2JF2RCCD4xAJkec38GJbzdDBHXiWWN42J+pK3UAZtCbvSYc
VHuty3qH6d5rgnTxBpdrZbONXhO2pP7IHpAfeQZL7g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kAQihz4ZZKbM1GA4F3FxnYNm2G/a0dlDO5H8lRuZotqA7Po02tPY27omJpn7
nbzLfkBeIt+hvEfJTMHqqcjU4cqkxDY0buoProZJLOdQkiHRj8KaAcVsyuSZ
sFHrJDg8Fppd99BLzqIn44dwOyre/gKI3B2ckTjcc3tIjmU/+Ec=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jeZ8KPgxuCFbtr5NuXUcloP2To5Ai68uWz6aeVS8+wgYeHh/XR3WtSX2wJBf
9dNZ8Oc7cqAv3LYlHF4itjB63+u70FlJ0M+WwbCYROBshv5+Mbyi5KeYoI+Z
wuwpPpHJUFlYx8bCh6Ud1Rcljn5TubWZfea+nftVU9MNFcHd8TXyPHPVPq3L
3LPtpnt22zCCWbFtoWnnBHglEF0ozFMjgzL0WzOk+gRQJIn6pJD5OZYPoD7B
hZiVm8BzKbpSOQtX1FQcF1qBo1qgZs9yar+xX2Z2nPscQ/R5AHprJpH5prwK
K2RZ8z336kvq0Su7zAahXOBXXNGbjfNCYptBFASwT/Y3hvO5VjHxQ/0O+nku
rTaIcDxaCzuqeA/JLRefpOcsY2QFuoyEzF5HrospD4Ks1HxXIFKppqDrgqsV
Bock41OkaMlN4+VnDn+tEJ+89Z3zFi1B2uWrodR1sTJZQzKK7rg8SMvljywG
luC3KquGRsVrlXf8ZnQcxWquOnTp232b


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GK2yCgtgA5zVih7UseuZoRKy/WgAk6QTwo1IUuJavZ+CNpX2A+zy2V3hlJxC
GeLpWjGwrHwKolLFongd3FipSKT16oKfSF2bExiDgldteSxGNn9CTLtUB/XD
P7HY8zskFNhW8bTmWqKZ4FCOGv0Fb9Yj/mEaM4DsBD7WtIvIr1s=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kydaqbKq0u251h9yE3ie8/mSMd67pZjDDw8AiK6GKid7AbcfqHdCn16N67/V
Ue3zGEXvS3IxslXIRnwEA5ygYaDhyG5+4mWNrp/uOH3h6kfAUNXV/G7GMCG8
G8XVt5G5j+xhNzR87Hvum7mCh0e2hyVlBCwBKUGq/Q1l/7Toqeg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31120)
`pragma protect data_block
VbBWc7DWhcdL1p4iyAvy5kW5qoQb8G/PIiCZxaLj49FAS71dAwOPmw4lKOgf
82vDGHMXORavnEBw8ilGKfXPqmPVQKav3v+ahig43lZDiz3GzBXEw/PcT8rF
K4kHcqhldnQgUT0mhgo7+6pWhIy/pJaABqljtYew1hAEy8SmaQQI6PBX0RId
ZpxbqUy7zUC/n1oNLhYH0zPwavQ2rScpYWyuZVvrlcWhYxMjPjiKBUSmGQfY
Usg/XWKDMlHe58CJeyODYFJaAptY22mNoohH7o4G9M3Y4xDjszfkCn6qSdvB
rS7wKPEB9dJsQjQiWBC9eWB/KyCfcYTaSz7Qr23BFcppJcb8A3DKD6rxhWDD
ZW7Z6WHj/oLQLPdpZV5coft9u2rCqKAE2AINVV4Q8TUlQQ4q0rLlaJPOL+iK
QEcOUtnS66CiudFdjhgssghmHDf02OJYtrdWJJBEax/DpxKF6LOIN5myhK2O
7I0TEE8dAFO8iY5ri5x8Hn+EFRTcGBO+Bo6JiNX1ap0lu7EYyesf2fzhPbkW
Dwaq9ZpEmH80hkijElLhqW5NgfUytW6aUPZCSEkTmwkzZojU711wfk21dWX2
5U+8rGESxEN4sQ6+NRG5VDj2OoKvZwZCT4rNP1Qjge3rY50ZkK+zCiGNXiXE
a/YkWdVM53JaRSInJVDcT/HgvejIDo/tJVMSYiSbdgQdDZtNzGJirRMASe6n
JoDCWWowZzs7uGJe5TjuZyVk6lwEDkwE3pXiGU0xEFMjE4o1kPbQF0CZJRk7
WzgcF9m2IU5rFiA+CMCGeP6VzXVyH3JdJd5ijfOW9vNnMjjUzd1HL+RTmxKA
ThjmmGTF0ZrnWIYB620+gpQpMpFI4QE2VpAo1BPs+E4mPcHrP+4bCpVLtL0i
RbhkCqR022nAAm5QcAnV34Lrzla5mnGKq4myBX4IzFKIzRLsvjEmOYMze6cA
u2CSFu6LOvgJeF6ZMBFpdT//HKk4nTDmcD1RbnAaAy5DbKHXyR7P9wdME6jE
KO3AHu95FEqhYXhNvRaOaJnJhZqwJ3Lp7lbjOHKRAdEmnlwmuiF5qQSOxKw2
fcYAKLoCmIRSmY6bhpK9zglUP+c5JykAwnahNV8dq3pwcFJk1HoRJgd6COyj
kTXenMoZGerBVzec1AOhXF+03w9SkC/grzPhA2jD5TFwk5wTQrdMvTCjdHHG
W/+sdV/Xn11eLuJeG7ZTITM7QWIxXUF3T0JYK67de3iRuAcIaB9ZwXVqsEhc
2M/sWqraX8EF00b1Q2Ao9vE7w9LbOo2/AU94zDEGir0no3HcHKeWC5puZYeS
uayc1xXWIqoeaxd1yAPUqmHNExvrQrQBD7qNuDNUPfV8unZhlh3Xa8kXt8Po
LriZXQr54IAP+XAzEbStTMPwq9T+4i/TF3jeImQPYCToR056RO05EMEHYpdE
UVqWjeykMT/qB4bIlioC57iwwAW7c2xcQIuJ7bJjG+2l0kdaY14v+XuhsJRH
yMGLI1Lzf2ldTUr3gN8l4MlC5tQazIxXQfKxveyH3Z8hoEWEpHTr8e6pSV5S
I/dd9GQvAv+9uoLkcF54+6Aet3KhyxmkVy4R8u/CeSX3l60q1r9M2eOf4eeG
MLwM3JPpkFw0KR8aQg7JGS8oFavECImhygG0p8y1XxCjLh4109m2HMKSg+/I
0iNTfZdS4XFKBClBwyWyvjHCLqiftIMCjv7+H3MwmBYpSoMq+GbNKHBVCKTG
9rxiUF1hCk9CS7UKKEmgCNqyNTfz/z9jfjZa2nOm3TCl3JXr61eQ8ydKVfC9
5H2NCnjjK9x7KQhQYW74Y6z8uud6+33n+txmNx5AdwgF1aDS5tgQgIBnGJ0c
EV+sMJVGnpXt6flyrbtfrPymqlDpafeWdmtlErG570tpRBeMkUbs8CSRZlZ1
oTYqKbuCKF+veKvv2AoVQplHp99XGgK4THElPtq+cHSij+wt6SeCWS/CAVI4
b+mFXVlSNqQbfERW1uCstNg6IFDheLmPNz44PkL+xdEJ8S0Egkc73UBp9caH
RAqH6S49gLxyinpyn2WhPcacM19bjbiIdovnHn7d3Z8CR3l6zca17Hv/AyoK
14av6mYx6QCFyBpH+iS9428+E2sj0rL+jjOtNq2ew3hMyi8ZEuY8UJtud5qt
ww0JRZMJth20UQwbLym2l1Le+EAzCCN2kaWcKvZoHXEJi6Vu+hNWkQFq27Ls
8GeGxctctrXZNwTt13ReWbimYEndCIl1DpNoB5I7nMlpKNZfqRFwGvubNHBB
Tr+xlNk4bXTNAQZQ6dxCIpwV09aAvNTVStYz6fhmx1TRS9Ipe4+B7YN/I25v
XvIsfbDpp7pBE2M8ld7t5Xy9LD8yUNPiJrBIHZjo7Jodatv4RTxuyhOZSRLC
T+9Aeh0iRLRw3sSasVOyXpCdP776yiHw5FlmMDN9XWu4lKpmUElYIUe/rmpc
OiJe2rh6x1E4tYFA1Vmdt+l2iOwQGr8tDFAsJ4m9GA1GuwAYlHaqU4+4kNcZ
azE6AqsGvqXQ9SYe1A5VtvgNHZ2uWRIt0dFa6scDLdyQxVwdLGBUUpu/bEVS
YSKSQAMj1g/CeKzcABfQ33jKlbJhHqD0vTwKGCwwCNXgUe+rpJhH2I5xx/f2
4Ts1g3ynaLgt5B/iyZInsKdkjwYh8butf61ZervOZRmbdPDAAZivz8++474F
AprwlsjbjHWxrvppyLHjW5gqAaUbXbO614tc2AkRfNLU9wAl2C+3otz9RjD+
lbmoltRvGCd68X/eUscDRoGbmlD1BIemvqeKWgZuJfZBGtmfowlj7Vi34I7P
pcMiV7dN1N4b2YekbF9yYpTCxXxW47meeBf0ZWbA2Z9t2yXfOMENW54GIpeo
5THkboUxv7yJF48nwAFdEohu2s6khT8UkiracAdpQQW6JKRa14UoCgCNSU0G
bYPgfHQE3meKhlINGrtPtF5FvhA+VsMhNKlFEFhvwV4sMTLsZI7tif/Z6qCX
MgxyEnBy101YVgtJPeaksgTtG3SuY9xCyNtbDa0IrHZwQpyg0ERR/ExC6Bvn
ksa8ZXkvp65eMjbrATyfkcoiwTM6oybOU0WbX5h8nqgbdtBjq2ZsdkHW9q1v
l5YWuO3Dgxc0lo/t958gL//veWpir6+kwwbVQuNPIK4LJpuSnB1UaRfeO1M6
vlPOPkfQT0VkHnoJ4DF8xvKCK2IEhCV5KldaqLdgP417XuDoHq6Z5gqmrnoF
ebL6N0WNcxr1TcBGPIO8B3PSWyoTPI2i780unzVnXL49cKAlUI7OT/sIAydv
TuigNlJzl11nqgsfJgpggFXkVWAfjfVqA1xBm7UrWK5Az8Amu7SxDoM8yPJd
xHptC9SD0VBrmVBGRGd15KXDUQH63+R7HiTbk/Cfm3IJHWDgrLcV88c2go6h
VnF4HVU3e56LnVFHefcNZd92CEWSAHTLkM0KSVjB5bp0RhTDJpaf6pbf5uyR
JAOXCy5DzexgzbpLwsQoJLvoXlkptHQpvJcYf43a7o3OPpxFrkWPFDFHHDM3
q8UGwOJxKIg9a9dUVogqNGUaoszqpBj1GKrLmKaIZQJ4tdYPCk6WwE9siEN3
YIiDLCBRkF7+A10vUuyQFrJxpOg49TqnvNNogS4e3ULbrWkya4HsCuyi/KZq
gD26SVRx0Ht8PR4prx3u4/BCBDFgAPTvciQMn+roK1ef+5sM9jFFTD8Ixwlw
ndF/m265+M7p6gkyMTbWetJ45Vkg5zGxwrkRo4S++I2pdrLtp/ngqTT7Dy7U
cNGZX33HRVOzzahjImzUGzdIsTgGF8EWZc2CB2XzqoUXJIJ9YcrT++tofVon
BexkeKILhWx2XBYA67WDh5qMvmqzILJhmplUVG2oQ6YYF90xp+B7Cv7egEJf
PzlTFuA6wGuuMLtWIhtf0vqOToZKNxP1FNSUMGfZFolpzU7jkoZCWDm0MumY
3n0b2DWoDrEe4UaTuwV7u803uE8d9oMv1T7vO4SLtsR5ZcxDSGqG/Dgp7pGt
Y/HnLEjLLNG0mMm97a1nZi3ZRkgwK0Ogr2NK4ckMj8FBgmbVMbHgmg7/k7EO
CYf61ZfEpA/twWByW8KnZ6/c1b0m/kslS5m64GGvMfvpZYDUKy7e46ih8l1F
JFAA8r64m09VM87RwbQweTOUheo+oHApbGWKcynWYmZyLKEDggsRxNrtBDzm
Cz1OPOQphyh6kLzbp5usDCs8MQ2z/E6PTbLoR8Wkpi15/tsvjmMv+n0691S4
+VmsfTUYRZNvaZOOd2aB+xwdySjFg9z8FbwTOipGdZnwTLjlrYgeqNDyQjNf
zKvui0kN8hsjsZ1Ydta9Zy62krpKSzWDZnMj81eLuDwcpB/ppJmprk7J8WoU
yNw6DuQLaWSkVk4zCQM7o7GRwotAV9eDDpkOKmNPu2kkyfc2goQpTQyHCwet
Fhosa8DDz2qZefQAOE/YMEbQvfZzeod/KI9xa7OZUrRBb1OKOe11cjfmBYFT
Q5mPYDOUVH95R2l8AB26XinZ5BQggQMLFZ4dZTNA30RDhBjrfqRzs9MA84so
aktWTa9YdIQ2SEqV1mV16SGLUteP+4euGk//+2YIHQE/3jIWMUROLqqxMn8V
5XQpsJDD1nB8UwEMjs2H+cdEb4UzKuUuOEng7ZQ4yLFxWf7343gglCpnt8a5
nWVvHWSfPVqkex+ALyXccOFmQ2szRVNNdeidQd1b7+yJkUfh1G8rjFWluYmc
yIJdCEfz31uX+Xc+zV1GStUaoitHsQCseFmvknwvR+7DTK4n6p7I9PJpJkJi
ikzq6c66m97pSb5pBwmIHw4duXDmm0p9fmduxzgJhio8+0yKkKSZM9wGVPJU
C5ADtZUUObTu01EtM91jDkR9Gg6pZ5XmCShg7Ep2Cmmt9Hdwvc2OxjPIlazP
Zbz/Gq0lbpJEIGWum4h2r2VIMA6p/3lH4VULooVr6PZ8X8fadZbbc7r21jUi
ymVlfv0UchOtLSeT1Xo5DA12Wb7HBslnjXry+NBTPo1EfAkTiZIK3ZpczolZ
oX2JJKboqZ2v+VNzdhlBZFZX/sOg8p6/cvwah7yr1ri2OBq1FmE0SuOmkJjN
/Z7hjlxbRpaaCyquHFeUWH64y1eSAe7aH8/svkkxUUzyIubiCBtjfbmHnV5P
FYz8WvHpgdBhozoRNocHJjga8hAVO0XITsylvIaBNha8q/dFIr+ya3lmF9Um
Xi9Ib1rdi7QM7O2HmZSLsBKA1f/fXzpFGOpb8F/2OwOKnTCn+QoVhrYLIAXa
nHvMfHGJM/ZWHuMRnKraFgYcUhj16DMEyKER3v8g6ng+64MseKhkjBbokBjl
lWSwJQNd8C8WIvqcyOmnImHLeHsQT/iDE4/hF9+IsuJBvW1ND+5RqMbcpTVk
95oRD8hEvvXE9Yayt/hKzLcOqiUi38gpFV5yE6cWD73wlz5AY6NmbTg6/jjm
BIGqGx3+wwaSkmDKF5CG4yR+c8kKRnXj2QIH9+7II60xD0S73ASZT6kwFHzz
6OyNRk5hdJfSXlWRz9bwXUodUsylu0Vp9uxCb32bdrzQYV0AjPMitkmAv0jv
VoO+FakTuNXVfIqPAJzBpvpfYFTroNU3kk4yvjPExFxpl8JMVOcqWkPo+Hm9
V6dn6A8eKl9MyY1BgLu0PtJXlNqftRxod7n2CuO+Y44hN0hjQER7HyVc455u
sRRwTzF1ZLMjK46wsrv8QaLsQAf/Y6MCT8pZ9w6v4i+/EmlFDJi7xoDtmbyC
BsBoHxEyb1zxVWkHcivBw7BKvASADDKm6VlYHBZPlXKJvjRnqE3zPKJsCTc8
4nr7XWAMM9z7su/V03eUAYOaFghMOEonAZPXJQC5ksx15RXSkCl2BONINoM1
G+rsiEdCxRTVi0alsV0YCsGz0af/hpfv3iUvYhicm8VRt3c4s67G5Xor8VBg
D9dBVN612gHJfzsWOqsQ/Or0bX/IRwx9AUK8YDBeSTKuMdQZOZA1FUR74JV5
opDd50QS3tR2w7POAtecJsOxtkbzyJ53mHHA2qkXnGn8CP1vjiMTRdEMoqvp
TYfvJX+FuwwmrP0XAoZJZd6tLwYltp3j7xIs9YyK46iG8jO5uoBnRRJmCo5/
PaQaOmBeDaUVtPzvBWCbn5avBVTT8KRz9dYVsJLCZsf7pZVFAwauf461fc0F
FqnD4vugvUAHuXUUworPhtlSiIW2KZrAJc7qZeBEEZDGidrIH1EioRUFofpP
Hn9sS142pyb3nsQkGUgIZkGNFAG2vdT8ulsccjrl67/25ziqYdot2+a8wmek
3WakJ3SqQpPI0w6xZONdGKYehBlonJTjCKgOoazDBPsTW/SNXHmxTncT9AlA
FLlkW11SDYJQ7dEXvWMkPi/kTRHJk4wJkke8yoWMlgPsXcCU3S1/TlUpy6vv
zsPR6O6YrrnZ8fHTmTeQ4CUZc/6rq8UkaCMf+vKNE/JDrf+TSssQj2LlM3ZJ
uHdJUG+owANnm+dktT4BQzUsib8nUeV41qun9tfdKn+ZH4apWZmiTf62F677
7wO9tLwuuZYog4idd2wCfDgNkKvHqyqKVrFRMeLgFHLwq8nCYuPGbuzf/P1K
4dmJChrBIP/+c5aIrF+wl99IsKl3pjGcvQdbMKwmonQ/QGc0tJNK8JWOm+SW
AuojH7VFJrufiY59geybVlF7bt0nZxERO0v7SKtJAwN3fkUdw1FrP9qZPbuZ
7e+0KB3/L1VliQ+fUWYttVTJEtEW6d45zTzTY+QqUqXOq1MhHzwoM5/JEAEv
Bv0rxOVtJEcsvAMLfTpDQLaEKyQsLZBF95w7CRltYvtfzqwyyhCMxLWGcCCm
I4uRtqeNGIEtiaFx8he9H02syPqx2pYYu9mnDqoTKwq4PSYqnz+zbMshPDvQ
bWbOIRls6k5TyfGp5iC2agH1aWfJWvGfGdaGTpxBpxbf7ty4za/QWUMB3bQu
h3AEsWOZwq8ws/t1xcPjHWY34iyYTPLEUVvR/MUQ8BkhHoTuLrLTDzh7IdK8
3XxVVtjHFUKoerLsTvxNcBb6gQP8tpvJRek/ZIfILLH4jLMGJ3KJN+DTb79t
ektRfKU9d+FeVMEuNpqT60mlVcT36rxk0QgqlxpesUcTXhmiJl30U6NhnhxM
WsYfejDTvjS/h8aJQV/UTHQhsNOIhTi6jbw2489YBUSVgZe/1x+5XjNmVY7B
UIHpPHeI/88fWCLr0Oj7KeRAKTzQVpw/3FIr6BrQOYfi+Spncy6/03/f43B+
zkFIGPLSWgi6xp56rEcjwqKEDY0eXOmu5ZyAKHWez+4uhV8A29lv2dqiubhB
Ibc5WP9pGwg68FWFdvlhfW4+Il3OgV2kRW96d5YrGmu6OmA31BBHIhGbPB0g
U5bRqyOaGjaJH6XlYIKgo8OVhYJaVB4v4+F3uZ1iWZjBxTaCAJTsLXKCI9Sx
r1VrJ3Y2j7+ec33z7D/RMvTkWCY10yWdXJIQz17ihjJIUSTIHS5z7EgQzoyK
KMYDC2JOBzFJHKhVhb6Rdk6sqyaT2JF/IL8xNBXBcnDx4QPSJjd6ckkNpOBv
uPYXp3mQRbE0lnpdX0HxwAZTnHNENatF/pC/twhB75s2LXmyPRdyx6yEFxkC
oF19K6jF1OAVzOuKcsG+W0ZCRomJZW49swZcUkTqUHWYFUkMyRxZ3Bu7sd2n
jnomZJ0b3tKC2CR4cBfHWiqeRTiEM0ZSlAJZRrDaOXqxzaDSr2oByOkz7eJM
kTa3DrwirqZm48X7/cB/DJ4YYLomBLydD0/7iG7zuyPrvfdgVVJa+qr/9pZ7
EOkMshdin2AULEpFxj1iW+YzZT+MxrdIvcQcAsdNhJ4zk/vQpfkKt2d8w+B9
gJzO0bMESMYj2VlCIvOUyGsdtUaHj+r2tC5r25plz/I7UmBPvF1ql6hgkQ6B
+Edai1MBXud6SedwQmFBX11XMVfM+/rjs5db+1doClQk2TkSnwuETYPljAfD
lyeMm0yW6m+zwp5EQHla4Q8TSJ4GlNAs0ug5xfA6X025jW8D3YDsv6m8Cnpr
9rtkxLK6X4kdWcT7mYQWoG5xUy8p6EiUcIQTLJOlAL/eqHLqKYtW1WZppQqN
8opLEnFa5ZJj7RPg52U2lXpo0TmJJ+WE+4+2MnlrjVKMifl/H/p7BhxPwquK
w3OBd5rQVj9Z0jEGPxxygWkZCPS9/TwnuvivApiQSSmE8BjMFZpUSJhBHPv6
Ebt62qc8iDRbO+fDAIiohTW4tAcjp90bCTvxwqY9tH5vecxDf2Zn2663wHz5
W1l2wfWNJ0UNBbGbzQLvlz9UYmS+KKaVwwHDbmHhjly3dFpEzfabcKcvoYr2
sAzQuC2HjvG4jp4+gsUtt4gs5X4qD4OdV8XAfwcQsYOQizcY7csB0YfYyiRJ
i/tbLlvefgXBTeOFDk/REnptud3xIS5XwcgLmNXPPl9V1mKT5zYz7zxd8996
c4gffbtCJ28/zUTQ07CKSkbULI5RNKnnUSJiybX+uE1Q8hixjd32TYl90D0V
jgJeSaezUrC3bU1veFguWuJyfKrt8E+9keoZnutEuGsA/R5us+6b8WJQUbnA
xriWLp8FuGehvOPkcXf0jykofCk6lqwlw02OtrrLtCtR6/jpa6Lfg/OkXGmD
AVusRmJuejOAc0CQ/IS1PTprNnlmlUeNrkWZzEXT0ZzEUZvxxqoQc2r+105W
Xbn5rHSvGsVcgG10IHYog4/WIA7nGZ33fLkap8y37ETFvRpwSGQPU3fvRggg
go4ALPz+/huw81t1ZlU6qrL3YRJdwBStLrxsKmNiinT6Igw4Tq4BRLAsKlt4
ljeE33cNxfMc0EPHZcpB5uDYA+2aQmbFwPrmrel9hkDTrPHCh6YlXt78dEfN
rujVMSUJAh7qCHx0hXlN6y0bS+7ZXjlCWmcL8lI25TyuIjUb1x/o3MPn2v4G
oWszuHmOr160HWFliI6YTquUyMtarMb4BaADwFCQabYj7dKevdYCdmRBdmYB
iqKEVs+gAt9sB4iyrzGtErsyBkxq7R+Kc8OeTIrr3ocj9ag2lXIA0zF9hlbX
qtlpQOpeisN/6SC3goImBTPA2WLjAH0v7aObPVI/EzebRoccFwhHZnBTuv08
ncp4zrmpvceHAgBlscWeF9WTMfsfi9Upka6WdlibXpGDTNZyhKpBzbzCpCC3
mRXqvn4JnWHjut35dM/KaMlvyHhzEh+yOCyLkW5FA7s4uSGRMYUUC36VsAXD
Qoah2mcdY1tGs+N0/Dx9f/En8QJVI2LWT24TEGphuDh0h5vlnnYjBZ4f+VE2
Cx6m5s1a4RpRg4fdX1NM5Sejn/AYcdwz/CUYqfSXa0MshCWICtcXVfnB1yM5
/59yfhcIZy5XSVKXUuPp6cWkamnkqaH7pIC0cNQZyzLQnONTbBDyQvcSWwVy
8D8Jt7qdltzreg68CPOmLXPfPcpC1B4gsdpA8Ya7MorzFpK6d6loUgkG9hOf
pH04F+U7c+azjqBJaSlp/Wn+SqoNmp+OrZXp6J8PD5GMnakA3vr5OuaD3vdG
Gv7DNWYElw9nRdrub1SSy1MJFnxJF8zaLP5kR1vqsJqJSo2UjP9fTgss9DbB
c3hIwyRO5ntd4LDPNMwDy/iXRq6k5h2a786x/Af7/X0G7TbZAbLBHaLw/Vrx
2pKGayOEPskwegL+sMO3TTlX9AjDJRogq+e6nu7nR32hcqZgF1TfDkUDAStw
jRYqcApszo+AUaQSGH1xKFqOTuGUYA+3CtN65I2T0GmmKZnhrDA766gYiMcV
Po9jEXd9EHwiFNarO22n9H1H3+mn7WNz9/BqntNfZCGOuArFCAr2R2WeKdrC
d4NBgEgcnwL2sZ7e1opTCP5UELrTydkSv7Sqg3FB4TFUXqvPG1uHS/B5vLiK
+GnkHbbMm9nok4o20a7iqGTND9lZKa/5fDxPAWLY6CYpnE8yRWo4QVreixL/
Fy/z/QltHd328Snio3DB/f/GW0xeSKfdoTksq1FLr3nyWtNHcQ7SfT372ekO
KCp12S+8zSF+PR0n1FyTsYTWop2adqDtIhuZw2p7kfxiaN2L3fMRVWcs14EH
b0SNR2PVtF/GCrfjU16VrbXG562SHjKO6bx3KK0bN6fvIC5N40j2j1WR5u8p
xSKc4nJawQkdasDSUMcfWJw68xUI9kkOK1zBPqz9wzGqHpb01gBZjrH4CjiL
1ynS9C4Ff6I21ehjKtG4H+7xQDyyIeVy7JEawR3Bz6DUtb7SwbTe7PtS1dEI
/Buq320s3zuQT2Gt49mMw1v3cnfZG5A8Cpl0aSbCzwzroXieAsPQUfbO7N0E
0XxwH7LsYM4bQiMAUbJQzjq1raXnbCuuqSIZdotWa/Y42+fQZy77gTzrpQKC
u9TiTxs8ZpIeo0yc2Ny4SD3UkpqykDvc6xdIst38kEzlVmh9ECQ9L8D8xg3j
vtS1BF1joAVJkciPKHAl5iZOby9QSvb+yc3BqGHeYPNcs4tUNN8JzS+qkxdQ
hkcrnDpbIVDSyRu+20LObycDpPbTWrOGlfmSlMia1QW+1NDd/T6r8QaVEWgj
H7AsJK4plu86xsGTOYMkiFGtcGMw25jTdrfzGm4UftFAzFjpOe4NB1LYDMip
XW1asOw/DPkhLh/vLjTzHjunHyP//XVRMLyLk9WCk9o8DKOefrW8MY0pYQ/L
54NTwMNCk6c8bs0RsT2ze461pBuF+4ic18RlfaqcWQnrut3NtPcLJyq7avpr
F4CRP6QcCYH+1lAojdOyEe9/ksn+kGhZGtMABAcOHQph8wgQktXFhbjxEDh1
pu90hHvaI0Nmozesu4cbxkmj3533CLfFcuRaccZRu3PJ+Rk1yGu4ed9i8PWK
S2kZB2BhSbwNkenPXe7DfrAZyjc49ZKwPwx1kuu6o+LGHJ0LAym0KES86Vcn
oW1A1a9jXN38C4awpLFQBwX+WE590j6N6p5iOpeGEMrYuWTxjYfyNOaDnFlQ
ViBBNvpdXxIk74xqg15d2ShDb9d5PEwp3/Xqg6p4lDN7TPqU9DBCrdW+d4lq
HHDrKfb12Sa/v0qI3dVJzGOuAxaqLm1ferUmhF0teLwNzWbjCjZ8JKnXdFGJ
zYe9yzEs9QGGeD8ayj7jSjWeKpmaSMTLMiKB7iyNcXtk7RkD0bXeK/Jl/naL
bF274zA6XaaYGDvVZRFgkBsr4jC1oZvu1LBJVobWaPTiSqhMjx+ZA8dAFJOA
Z5RCspOYCykDnxsiRdjK1JrDyM2Vsfex/sQmQ1ZPPzMk5JWabWghP/GHOTrg
viKi61ZqAwrC5hzzlVGngzCyE8CrPHssyE75HHF+SzZ9ihviao5j6LSqYy4S
ropnCybDMTYnSMl/wsv1EUdDjfMOYUBXlbvFO1etZAY+V90NGypUj9XHBsZ4
U3qwertV+K5+/ZfOQjgIUO4NQ572qRt+gKhfayNIE63B6x3Vy6fBWE2lGKTN
8Uh3gKZzgOJ0iDK4ohVNDEz5aM0D+xjafvPuewvaznlQqANzyjGOrkfNuCvO
GsLaDo4HDd9ap0G6h831VWp2+9Iaj3M9TI7nGcLNv7JMbzvEHis8cTapie0a
WDUk9rf+MVYCLioZT+EHz6AOgdlt+6nM67vAm+GSaos1B0OILJMg0koip1s6
YNtNwb3QKXAfgqCOAl6DbYnn6VjBC26pLNEqeaNdjcRfHKO8BfiplbbRvNnh
wvxZA9Q/191iWInv//5h0Z30uzfd0+Ue+kc+uKxtmh4cPlrqWsrdCH0llyTO
0sxcfEVYMt7fgHuFnH/9s8gEPXUPmjdipFnsKJ1sUpcDVU0r2tTrkPoy8lTt
UZ/0tm+Tg2irWe9PAXAUD+NLzDo/evIJ/dZd1Ux94rvbBhFHD08aL8TmsJU1
ut3Gx84Smn7Wg0a4YJsnlBpK/20eG34+tfV5OAhXmuyVgWezVzH88lnrdTOP
B/1cB+8h8Aar7xNUg3Xki3BnWuYBYFriGM8/tN3bqLo8t3aJBGdzkz+a0nwR
WGYtHF8+raBkPXdo987oSbmqEvukKQRC0KIl8xP6dtq9etnzuEkChs+p2O7h
aHnpOF8G9PX7365nxbzqnqxhxtCt/devResyz44nDXdnB4V8VTafRQkY4fKH
zAXm7YqH9p5sapRMCbk0Hhi9l9ATL29B3UxA6VUPUEVOxiFGj1OZmyZsvS+P
wyxlOl/ioiLFheGCG0RcDKZu/DicqSksJsqghDnpqXFAtXeD48Lcle0nWdCn
rSaVHAkiS5QqSjlP+XGCqz532DVk8bh0su+VAG0XOmGZaAUFlgUu8Gz85a8T
lo0AjHyuixVMEeA74feLg3xVcyXeyHweAY6JTOnDxnZoSUd7/GL7zuA6gVnV
Fi2vnMXLOQYwZNhiDcvJtHwcZPOysg+VZHaPH5cwPNuV/ByuOGzG1FgAX652
2Ldlse0VpMBxEQrvaGnlnU8z/uZAa+tGmBvX1CbgvksWCFnbXVZ6bxkYPBtD
pwHRgCVR26IseCxHBN/joW7JydZZLHk30597nKLMxfYS+19oPSjrAS74UaH/
y2Rl+PdQeDYH32p8/UsG3Na6WUsGhfazASKKSRVg/Llq+PmaZAn8MymTroLG
CcsEggeA5FfEWwX7R7L5dAcHdpSB/gSNDj1uXL2VD67SLNyX5MU3xwRkt7Uu
OTqta8sVVrsxPoODIl1axG5pxLG6FmAK8HYo642sioOo8AimpVlrgFui4vQd
PQetUXLGQgCJXBhKxOJlW1ykKhNDw7RtWFvCdxHpvLWMe5JS08LaNX8dnjZx
I3YLUQydKIC9H//o+MNSRXQy2zu1c2IFKXxPaup+BWqAeaPSOyMtoynkZ3hd
QLDQLkgTI4D5NuOOMn2FPppDO4BDSwKm8+K8nE/8ifvbLGiR3Wvy11GYVZFP
SwNBkAVoX+ZRKW2hWzExels4RSXvdh+VA5GlpAo3PfnVObQdRc3rLmnOEWqD
eg35b2oCFk4rjArTMgG8U1ohBGqj8m102vgxqGBhNDpUePXGRcbCkRGBFymD
HZy3kPFWC8e6eEwC5HpZ5pdNDkjYrBF1jh7uDcnVuUuA6j+0+VPa9j11w4Bm
3YyayMRXQjNnoRwWVn0D+aL0+xMjdq1JscxkcPDTDoHIoMVWDRfLJTl/ravD
0XIulhTWaL91zxxskHDQSiHyqvVshdYFEGDqYjKTFLlw8ExnpSi5BwG1M44y
YNKGAQl1vEOunWCIAiUSrTxXqUKCAk9AMSjNRug4SWwjvHS/0Lv8ny1Fhdg+
5WceTVM41S4mdUf4ckhKaswB0dqvbes111eeGNHQclBz1ykgR8aYGIkQjZyh
4GIDjz1NPtm/X1ENAduClKnLUJXiSJtQKjy8hKzgXDO/whu5xhynqVOmceO7
LaqzGTy523Bw0bkgu+YPzN6XDd6HzX4zrSs70pRsRXIqoxqvInO9aUq+SBkE
IM2ot1unaCutfmxZ8To6sMoSFGAh9dkof5+PLOC+/6AnptaWrHhSbKxBwrxg
JP7H6Co5ZvMXsEnyO3vrMLDDeo+3fvVhQdJjkA3GjwWhna85r81ayF+CUprm
wupHyN6Rgp+4/8WbHxCwYNAjIAcXfQT+K/W4VDfTscswTRO/Teon++D+93Pl
MeyckaLFIAfPlEZOi5aAnAf+MbqISFhC6TVNSv4ZD3HfbZaV9mys6eFOeSoF
+kouqevjTfK57G5VUCKR28WvHnFJL7FxHjDhIRPxPhvYBhuAQt1v8u3w5C9z
TAwUUZIkJLH6/X4MjgOw+GxVenguXIepUoKmoKtMFfdr+bjB1dqOFCgatkXz
rqIJp6Wv/WXzMJz//hpgcyTkEDAs+Jm+ZSTPXd1E/3mueJ3StdNLTqArzjSB
AAuaNMSnfhcCRSf0pGf1i3fuaiKkb8Kc6aHt6/6FztaQ8rgsteEqnnRthgkq
uaWjHssV4jqBy76Zi6NXpnkAqNPUiHusly/JaImCWRycQAbKUGiDnC2jjuZn
i5ZjhG0F4sw/feoY1QXsoDew1VMkWwMWZCerbxWabDIGCPfsGP5crZsyrWKU
S6ILAW2l4hmzLmLeLhtlkviSFd32ZOU8mS34YVnZq0rxhiO/0qUJB6HDT0X8
KadY61zFxIrFCuUKXzUPL9bV4L3YWIcOAiyeDjbipdul5e3NzURk5XH+VoX2
vFPQUmdVCAfc8DhIDs3vnXAT9iEGecX0u/+FO0xjA6hXauLrQ1M+p3mEZ2tE
U5Icv6LbdW/gu2gZOq0wMmBV5QfJOBW4J6QqFIBs/SoFYVu/ZvPyd9kW3Jqd
V25GSWcNcVqcmo6hGJB3CVQsyZE5D/xtCbXxCfzU4Tdr4V+hZUXRhy/Chb2F
680hpA8FimZWt+PAgacHkxey/5hWhWVu8djJsZOSCuIesrWzwEvfsCsqDlao
rqurEzjF/SQrxhMgnW8Jd6fda9mHhIrniRsNwX1sPjA+/iKY4kpXoeDKmuKO
L3umhG/EiW+OrS0jUlxhMwcW30iwvo5AiIixl/tpx+t1+RS1cflC/bxSs3Av
ptrB2/WSizdWepvNYw6by4h+1Cvy9XeyzAx5C0s7x/iMEme481Z4mcBOARgP
w3KrrwaVLMHeK9FQeDYbKO7h0MZei3aqeiERpF3XA8byXs6dGiJe/txeRj+y
8yaT3reWL5Aa7sfipAlBzXbcN/DTLOvlNAb1etRCzlmzc5frWloGnohaOZ+8
tIaASiC/HRq0LLDHRCVs0IEr3Bf8nzL35+I8QuRIMC+bBAS8Lqnsf9jnRW77
mqvyFlluvL6rPa+8Z3+xC8KVhCRGenmrpsP15zuChQ/Cjez8K5soPpyjOQ1C
VWcED0s8JxfvUxbsj6xeYcaJJQST38YbmAQqPmnC52ZKIyFSueT17VWIgVhe
a3AQmMYd+a3VGI3X/f4ogf1h502/AWDfHmyMDT65BJfS4BjgrQL7COfP7Wj6
mAm/1LMQbBZpodvpkLleVPUfrqMFMDKelblIBUJAnRE/GTM+HAFOE5Sl6l/t
dibVlb9zkeMCkvOfFYwPtxsE8IX1JDSzVqh4LGPK3RZb9fAIiIuz/ZrqFe0J
49yYjWaZpfc1HuC+FeseroQ/8kCzFxjdsnxPuMljbIg8UYC223RMAV0fE4jR
UHyuaVUwsVrCnxd5KjnQzMMslm5U9ewHAY7n7JA2yge5wM/RXSKRIOw07PKj
57PhrmemyzR9IuYSIDCFpcsCiZrQtIYLZAZnmWzAnLT8poeq03hltDY1lX91
wyvMhO8fcygacwOgyRiafs3cEB6dLq1nFRmxnvRKoZ+oH6BZgs5q30sRBGVD
TvA5Borw53IrtyYnRu949PzMoc1Uvbww3qT4/8pSwgLphv1lXBDnObqT9iqC
VvJcNKc8GmLtEdDAEiDXpWVRZRWsvvDUePYiwU4YmrE8h4BdkOS37+hObJIM
40WV0GT+L4YlYC3zRrw8F5FdsW0cgLSq55ScM8S0L3R32UWYPvNeXxL7w/zw
sewGYHqx4lOedOk+NXMlKkwdmtD5zhtF3KOfWBc6UYA49csKKd8OH1vPuKcS
/GXVs86vwMdTwY896oGotb0UWzZbBRReOgdF3mCmwaiQMe2a2UYkWLz4iw8b
9VLAhcBRygne7M2SgjBSm0KMEiXSyH57WJ3avTIf6sp3LpDoYDo80esqevht
N7Jvlc8vjzfvUzk54WYvAUAL1/c0y6/2pDUaFitI260SJ+tQ1RINpAtX6IEm
fQtZJyKyftMWN6HfddDQPoeHTjXsYOloumuznHpRvQ92TtA3FUhfLSQBdgsa
UMocm76LepZdvBzFz7s0dh9seFLtMU9h5baZ6YU4jXCJNYAOO6VspkuLouLg
Znu3z1aDr/aAe1QyXBk71uMMk6So5tNAPvr3xPxgy+54WzBn60rhC9Wu21xu
/lytJJLN6QQ+EdBhD3vhDBGPNfiAltMdBLyX/gNJ9wAiqj5Zg+1nCXIS/PLX
NR9cpUUfpe3rr8n7cRecDRWjYrKhA6eHwZ7rTnziQGqfnHZBRYn9Fik6C7cI
y5zXzjg14/EvhBtk2XeHkEMSZ0FPVwAMwbBknvDKLAJPsRGjwVWI7AU2Pldp
12sH2//6DVt6FO9c5izJEMyoMqwjB4rxZEglbccXBed3XqnlCVUhuK1zpHWy
2EutVWnmaa3BpZJWluDxArqLXcM9JrlI8J0IEG4jfBVtpegDQj7/tiJs77gY
smvMec8feEB0KxRjGD0YXy2utNA3nA6VAMf7kL/qhyGT6g0ZBcU4OtFfuMl4
NG6CghdjeYRmDrQ0oGvZjuh+n3g9KRyse1EheydzxPZcS5TvBm0/PU2n7huO
bXqffIWdaaXSN3VDn9q53v0GtA3ApHodcq6IDbFkXwdL2LUSfXKK0CTJRSc+
dseuiuQ367ebJoka/eBtNuSUNW8y19j+4+nTMxiy+1E4suIJPz2ZldF73VaM
VfMrdSFPwfGOlM3ZIYz51n0o0sAaFufhLZJs+nESV7DAWhgMuTr0wvXWp/kt
/gCFe7i7CmckcuIhw4ZBj8iPWemlZ6WqjO91ULAe7g7Ke1VCDlNhbJ+Srm0g
5bQG6P8mIyKi7Wvo59OluSbCRS0yjq1ZSNqdxW4guHzzEmgmowKXhHQ6IqI5
dWslBC5YIilkAvy2k+xunVaL1ESkyRPKuaOkLv8zFf5fZXrqzV5e53LaKhnR
MrE5xSsw7XN5x9z+hevt4kCYUujqbJ5iVgSA0WfTkUnYX2yVovsXQCg5uONu
H8EZ8kOrZACnqT3CkwBdjqoJvoRNPly94WemPy5qganiPBxvF1EjPlm1i/CS
/P32crp9lXBqoPfIj4Gj2GghJFX5VGWVU/6y48tW2b9eXP8LAGcRX8ul5nJq
UVnsZQeMYiJzc2KvSGr0wsjwKO7MEbn60/y7YgUYJLV1s3piarYD80CXg2xN
CHefAqu8yAOfYt74REgLRgirws2zQRYPPsYEvCjZNWumlwOEu9RilltcEpSA
L6DHiZX6Rw+LrF9SJTVfiQB3dpZwuJ6zQSHb28kINNZ+L2M7cOUse3r8sxAi
zqTnqM5kKeQmFUJdS9Pup5E7jpvF4vmdYb+XHk0RBMHiLbrLrCQNny4E59pL
yehfJvrYTXDH74c1YMBpABFHPnBA0qTgM3lgu/JbKWXOZCBD6RrSgvb5LMTx
X8K1cziuJ5U+Dw1MQRa5rvIVWqWB9eVcAkB8dnLuKfCqKLdE7cAbmbrfpaDZ
pVvPz/OqNO4YRV3vWxbSKCjqTBj+Wzsv136dIzTtuzBClXsN4yxs7APxfJMn
mNHUdgjAk5H6e4JPfkGaTth3wuarKoZGoGneKVq2EFc3ptDdrA5OcPtweGY7
fqmrhjNZRZO/rkAg0GFTuZ9bTRs4TN97/cByeXg6QCZVdPXOfgZxoSZRa4Fa
YdyDVwZoc6uo5ZVdDGaUN5k/9aBclQhHpPJORyUD97O6ZswRxr7QCPL1KQC5
moC8+lZCXKw5RPc60JEEuniZ1sto6qIlDZwYS9K9m6VwaE877wuUllJT82FP
uZLwy327LNidjEhHSO5SfHtM4MJhrMUSjqse4k1cqRThZDEk7W48CjY4FEsc
duJ1YTgThmOBPUBivFaPX/xoLctiQxpcgyLHIpxLTMu8ebCQCszOi9H/A/o7
iiXdLNiljXxuIlA4+vAxalBF5axClCTiKzJ4Rhl0DEOJhkjyKXMVoGTnu/9M
ufhc+XdVhlDTuOeP1wakKmHMKHjC2fag7dDfaaMAL5edImgfhSmVVgac/y37
iVFgW789A/LpcKtDRMscQ9SfNC1p3iBwvEg9q2p7Hv5iDm6nQ6aLevRmOF0c
wC+yVdkODdZ5cwK0F779pyeToDbzFmcsZgOZJME0a31X1jMkHGWXH0VKOX+6
OMKOVr5KF5kV+jXsaZFEJeB086hW/aLtJ3TGFgR9aqAmRFpjN1zt/Qjz4mb9
JN221Uywyv5Cc5r8YZjtFjSi7jLBM4mHGlnhs58stgJBoXq3wCjQPYp+hVTM
cAAeeQV/8yETjlbDYRIdy8m/5I/pJGC0M8VaZknoHK4Wf6tDVTbcgwfYzlbV
IeVoqV4e5xK8/bp+s9iojax11W9Re5QLQiVZNZQZjQAb0Je1IZtajAxYrecl
O7WHRyDL5h/w2w7wvm8TAw8m9XdLKzlXiX0A9L0EkzthnEuZA8OGWjAQRqg+
qxrWTnKqvKN3AHht+HZNsPWJ0FexVnIqCGfNDq7WehG4k1zr0/T3fjsEWO0V
XBVht+Pcdc6dyt2U5paRP2KBx+q1guJj5GYCMc+xzUHDF+68dBI8iz84/EoR
IKzm8LN33iI6c1XuK2FCPTMsQIgMSxIBKU0/XXBLXvZwUoagyGeUvzVNnidF
n6mF0Bt9MihqVxmyFkb0DiTR2l8xAmb9Mq+GFd1OBstvrmKvkHPsM1mT/Tot
/7TyJ3pwcbgpYwkP8IAV+LcHw3KORSnAFhnOr8CHpxcZTsi1j2P258RGWFAI
GISBI8ObIuPUKXhrZyGgXYd/elpPg3BhPwQfTEk4Ym7eLZ4pAbfXlSRzS16+
u4kSjQk8TUONBmDT7evI/WfuzX+9unoiR8he365wgU6oSfZDKmg+kRAPdWlx
3E+HFFYxz+gcGjYeYjHI/BwmuXoNZ3r3iJ4eWaeZfrgL52Py/bhq3jbbaW0w
DNJpAWg8RFzVa50bwU/T3pvwf80huSkOpLKAw+MSNWNBqxUBGrEe1fQM2GFn
h+SzSC2CzejqZiEwQkwsi2e2NGYgW3uM8nGd/bSTmjZ/gDktYEhcMLTeFeS5
SFY6LrEUxH1eXTkHVYd62Nj0MN201w+198p4qPg4dcg9bEINTUVuaOIfplIS
TrwXV9emXXDUwnn8C7jhQoT7Honn+Ex6Kw2DztQw1jYo3A0EVYHAHNthEURZ
6ihk3gV1LNUbLZ5yaWdfPZSrWteF/fxv9cvmcvnoyIeTPfGk08bqpnGVHKkN
znoGMHNRDQOi/dHTkzSf03GCtj0D56d/JwEx38DsNemcKhdouGY2DrJ5ZvJQ
vN0vR/i/tP9nmhYmHwywZKrajF8PvaFDttVqUX53JUqq8D9/q6lVsjSVbeHY
AhqeKBdwBR2IJFn49Nbb/Yp5ZcJderfFGVxp/j3Uxono463LGPMDUTUBMfvQ
x+CtpJZnpqBt/czRL+pafEYn+IUSTSKRxdgIlJrN3lBBfUI42KoPRzlK5YO9
3U2d3KybHm+P50mpq3eOqKoxQDXDZqEbSi91MhV1Y0EJLa0Z31PLMJjSjSzy
tI8ddomE756V3dgvzpPN15NuNyIvH9J/LiOFdKHM0rqeAHJxcuspO4+x9Pq3
+FKySQm9GK9wJBHl9aZT7uzJ0EFEbk5W4wB1XFqXnN1YxswW97DwW2B+pLLI
DIwIx85FH/tmbp46aMIC9XpDUF2ujmLUj0Vk+UDTIv5S0cslznuAEAyxjAZO
d/kqqaLDsPwSdU/APj0eWZse8DTGFLnkSQxoChw7bbDnTqx9XnuVmJ0YlNWX
lsc0jIpqbKYougvNlxgc0HrqHSJt5+buG33nYL0A9hFVJKoOeDErlssfrTsZ
7G/Atee41o5ws5gUMv4nWCKzx0ES6ivX1pfkeNujSOMgpHzqEZ6u0CtE+N+8
d5GReDr+uWYcnVQApCRcMm9F4D44KMGhrebtcMSJxkbRoJdHYntHQ7s/DteU
gF4rii0FagXxG8JGbI8xWv74LoEteJAmmiEZkzDRxUBBESTmYeeRZf7JJvCJ
0y3afdgNZBpX7qP0clK4C4vXFBTu/48uXaTxJk8yRJFJmJ70YrvNqfWGbcu2
mfiAgUR3gbbia+tyWcaCJh4Ug5+rj8e6XhM6wXLr14WQ3hzDer3VpkaxZR0C
s8NF/cvHUOPPmuWq4k+bKIY4/m3tmGGBp04z9dStkHA8fXS3MMmtYTwdyNpy
TBPnRha64+KWb9PvVgxcdjFWSxZYw7j4y1QrqDoEBp2qKL9enyLM/0XkBnWb
CEq41qofzbKcSjz8dX9bqEUcD+WmMY4UCXTijbmueWBc0WKR6VNnuubeyWAi
f9gkyE4SddNx3M+NzjYyMIZq2Ha329YSiVzi7t4y/RVJKck4RaSC0UkTWjS5
9+YFpDr5SnlBdOPxr8VutCcgxzdoREL/Obmw7m8St/HHixdMc/iXISoxHNlm
w2Laadm6REik52FMCO+mco/edjJ55FDWb9PXY2m48nd2ZsCNOkObzpVvYfhA
CmpbNUa5MR6hEh22zT5CywsPfTSBN9UH30TgjA+dPNFBAcD0PLR01d4eD/Kd
SxrSMFE3Qn7/xajpEuTNWBYrGFqnHBWG7GfAh9cedQJh47yzANMlNwFVQzHe
ju1iw4Lp555SNG+c5cYos96rBrK5RbEdUln9cSoRp57R5990eJmtU8jwwGs2
HoQ1oKImLaBMNXMxh7rsRSOaUwcdyCZeQl4RvblwjxAPhmhOa5CMnHhUBtwB
zc4bkAwxFsHkLYuUIHVigC0JaihLFSZQ9UXvqQdjYV1Ef8p4dZ9idHwZJxYQ
ecmol9qpwPuplGWJiWYzly4It2qpK4/DzE+n6iCtBZlfpvzPFFyt2qve4824
Ig16uMvYmuJPCPGhUopNaHnPuWrAgatNU3yqHqc+Mz/UVF1ReCCyRu8fv6om
9lErr9TY0Lxkk/hGEA5AIxgoBrCiV68YClZxP9a18FuxhJkNCq1g+T8aN9kQ
gS892Gg43HdVXg5GJ1fer3HvSmbbkvay5Pvfv9qxFwDEbU4aysUQrH09mL3B
N9V/Nc9iVM73bB1YPhnTRPI3k5P7tPRrUSMKsTsM1qWBdLAJqoyfbQvwS++v
nEQDCvCsFm/U0txbEr4/xF+su0iQi2ZYgbizahNY8Wc3i/6oUN4eRw6RJDw3
0H/PiqPRoSAdkQnNSPHx5y5zlwFsnx2YQXf1hXlmH1DTKx40TMySbQ3DtPdU
R1+JlRC0hZsbyJ8iRpygqmG0w1mWwh97xzb3zSJcHOSUQ2HRsOTM+9rOlkj7
LwwjnX5qbSUzB2SX3NJd2KG1eQUuf2QjIsPF3+aVTcjzQhZ3OvQmG7g5bZKO
LjTA7j+pWBKyFo70nS9uNBNpSX2G2DKZ94JIaTZ+3TbzR6SKufsAE7ZnItNi
W01EbDudid6LszwfsZIuF1S8FYfJBXVt1/mvrcj55nDu6D6sko53N3pIXaHr
xa5xaqllhF1dxUjtWaoJjT7WBFcAAJyUtsehF4R8Ny5maNa3jtEQi9b3H7Xj
XozwQudji2y5MQMiXyWREpDNTnfcLe+NuWpRHmE9C2XQK4ikdgyyrJCqp51v
BYu1ZFFaTJ/E0RspmulPYlJVSJMbiIFEC2X97IY6vWSxSnEoqhhP6VIHDRzI
98Pv2/5DQZeUz6hs9qj9yuMk1mD8bZkbNFkU1EeocDFLYRwlPny7xsfX9k5X
bknBf9zxcapXTPgMBRDZQED/Rasy42RWDLudIRHHFhlZiielBlG4I9bR8fqo
UdWOxNnSmNB+l9SX9ulx8X+XkYdY6UHczN3nHNai0o7Z+wwKLQADjSscOG9K
tB+ShkleB+ovx+/ruX0wRKSZ/+AtsGnvPQMWwz8fqZb1tps0bBV6uClBOdVZ
6A2AMNXr+fcPkvYSMJS9iFZxUQyLGCfHmM1LFn42w9NaYfP3gwbFgmdttTcD
Svtplm7XPY+8PNSXxXS5uHy7SSEQIvAVGJiOZvtpGZEGVoHZ6jydvTkIkuF3
YKUr8XpywF8IgtTKCSHdrECX9UWD5ACC7ijXoOTxfne/VuQXGDQvUANR/8pO
DSrZvCN14JgsCmU3nwriL3CVCwmh4BqAqIVdeKYU/rza8u8dXMGWfsUSOuXD
H5z6yz/8SNQzynkEj9Z+OLZ1jRNRrGBegi632SUEXKcLYPGvESz89CEV+pLz
tmkmWVMAxu2KOHN7CEZ6RlLtQ8s7yqshYH0q1O0zIyz4Mkqc/zBfzQyrDADm
qXiXjVkxDDeBuJv1pnwTjrNEbFqjW7jAsFYoW6llLw6AIlYn/Nt2ZqRRn5sx
xX/oqpdu1kfRdqx/E757jXd0AU97wrCmo7P7aSkwnJUzqyRj2vPHog3UPD/x
OF9yEqXPTvknZu2/oKgQGL+kkkCNq4Qu0M3Rm5A6ZEW/AdZ4We3ZdMh5MloJ
dninjnL+m6gEOTTNcRqNhDa397O03mk30hSO9X6FYx+kU6qKUpmkeM6YH6kh
4FBcDSeUMz1Cy4A4x8z4dZCpq8O5z7OhX2WiaqkBZppfd8telVI4erDLm21M
L4cmE9WQUymAQwGB4W2684BxoU9YIHHHODgfXh58YUyJD32i/+t7cyi+wVXL
N1Q4jJ0H7z8s54OmI8x8BIhXA+iSXFp1TvgITmTkSaoZoymunFLCedPiSY8f
kMbrdFCwOaGGEOgWW4A74TmSWZxDmz/6K4VSLmt/c5bFxAsEx92tD9fM9pFs
85h1afgvdxzYRx2HdEejdm6rJA0+YGwAvjtm/FjP2kHup72W/5Y/lF+QqRn0
U259uW7ftn5r91SXGhwJ9zuMKrlvvV2yBAFdwfkCdSzK5igGoMzkxeKK4b6B
N4n6lEn54xmRNwZHHidMqVeUdIGA+LPzoiQDBwCOvb0n6pS+3OqyckEwGMy1
DZtfvBqGrYDyOMbuMfvOffSBhwM9T0ViCJqby0x2ThD+vPhiIR8ViWyx8OX2
j/OjTBKfPFw58LSsDejIcw/S8bjX7903YYIQK2tt5zPf+UQrFeQC0mYeyFDT
0ivZZIpBGITKRBd7mH5r406mrtbMgKvTigiZ5kR9j3dUdlOBum00UGk67tHc
DDE+Azom/4EIVV9BeeKiNt1J2Xdh14ipVm7wtKJ5RUVae/6YbAyVG0YIDxT6
BUDZz0MV3sp5Jm43VJ78Q7SY/nKC/T1ui8UGULz4Z8zMRBySU0oM1Zzu4rmc
RRBnWq8FwLu2RpvoPt9jJ16ckrtSQmKQzQIW31n/sBMhr5MDEnEASuzYfqeK
AIs2vzYUfA+7Bsz4gAviRk2bOluBJN5cd8+VwDN6TegC4aTIdZl/dEP2qUbK
I1vT7hySGSbYkzTuULZXYjt/TxqoquNtvjfC0eO/MHKcGhTq/5H2oyzz/4WR
tSXx1SqybqQNpR75vZGvq1KLZHq7KiZXnhhV8F08eemq/71A9T4wTKbsk593
k2WDh0+y3HCdMkRhjG4zbkhkFvxYdsZSNko0dTtC8LqPoymsR1qYNR+qowBE
pjC+4rkRhxcWk2leCYwASedtPqipueX+ZlkJJomgNMuX/IGXnYkPVH3VuCbc
HMlNTxIQ8carFiza8TmJPs24p5CjhEkYywnjf7uyPYmfVEhXGnTfHmdQACdr
8HgvV3zhe03cDExbE8vJjeldBjP49aoZIS4z1hZ3AFlOhz7vq8/bnC1pNqXu
rny9xkV9Durf7ZwT7pr9u2aeFYUZc31+6YQoQMaB2E3/lq6M5EZnxLR3leQk
zBVzsiyS6aqgHiGaffODs5tZAbEbbVjVcWrB9JJylOFftdGEj2uBkVRByis2
HA679Yl52B/3UfsHQMb6WTN7N1oHUWDtiDwYhrZJ0a0mcMyzM/eMvIuRfYM5
VbeybbRCSbli4GfJDfxRp2pfE1sMLVnHAaDRKzEoGlLKh6X8+iiapmlykgQd
oUUC8E9dLXm4yWitCD6gsricTop/pp7hNu/EJ5UuntAAKPSn0bIC/icxizM3
S5wsJCIvQim5gHhUs8SflAs2a/1Vlhr+sXhcTgBe93PI81ow9BsXm/l+OD/S
MRo4agdO8osBgUHDgAXTuDPHqObMqvrDRW8b1ZrQFm9DnXfQmMTGFjZ6ZP/Z
hkTYta0eJ1sujNto3zEASqcj6S9vR+ttDuLRds4jOirPZPw2izbfQzW9iTyN
SaMCzoZdB3RcfD73L17WQ87pyk71lAEU0XNtRJdk14AykTEOzkzcip7xSTfU
ZTAj4j7xWpZ9SEqixjFSwGAhf2Psu2YTTzVSzVG1qCXE4rYJRNb0OdjGMeWO
SLFpY80xWVseqhnCHS56SwIoKQjtwtQ/HVYS5+mzyqWYdAl0Q3hqJ8QBR3Xg
BX43mNcHYp6h1YhOjDbSp2ty9nrTQE14lnQA25k4+Tj6/oKQk/HR0y/cqixh
DJHcF/IApMJwy0RLYe4J4OVXeKy2Ve/7/KoNpmScm7xdMVoc7hOxzVnrKVpi
iyJTtP7mkyb5cP2tO+R/kLg2B36Qp7aZZWCwLLdk4JW+BMNlNDpZAzoRMAiz
JV0k2imJf548/tWbjMtYuNfdFeQr/wjqvludU3zLPpADgRcF3HgufsTJHi8F
OuBTl2BQ7AssUVEXtvntrF4DmDZ5me7NUhB7br8W0wOox3rfsMchNis41JSO
Nt/TPs7344LJCcuLqlz3tweuFMGlWkNOXgjLn0GYfRPl5gtC+uq8bDyH6zRi
fcrXa2oejjfGZNXBYQ/gcjX0Au6mFjEd7YsBuUFbMSgaKwqoyKAuOUc9vS6G
n0EzlqU4Wj/g2QxccUdYXRPXnOTLlhwnXuO2XFiUlSQXVJFQ2ZLjRrRI8Np3
CnQ8nEIRv+9eiKXkEnynLQ3tB+yeqHirzo3QlZ0pDQmc6UmlS7cUx+3JyGxu
kFKn6SfhEMiprmVX919qQ+d5oFLPn/kx9fs7Dof1LnzihS55PA3MQvWduM31
2yqjmcNIDABsklDuIbqM6jMHFwbS1CcUnDNSKpgik3Agpr65w8qkiExpdu5k
KIUQuYa2ksbFK/ZGeX6zFkjxydDuFMPrEPWcfIaoSZddRW7nV9ik988DC381
D1hRyspzqkm+bI7yL+32LZOo8Aekbfpy74K0/YnMD/5xHz2VsEgrrwZZZ5UW
go4NDHC3VsIhrb7EHrf/XPOZLKdbJQPlAZHhGKDGdsXHwUGpu7CHKR5WBKZM
CPaums72+oE6uze3+KpaFgnXXGvFoEXY5UI1/6odDrCKmSwoveL4u7QFLsvB
uHQRtKHWA/xaC0z00m1N/va6rw+gYNL7Zai5yO6Pb7tZ7aBJFzMgrNhnoZJY
0l6PO6sj7XwUmvDNQvKajGdJDsFTYxyx51DMM+s+P+bU9YhA4+u2AI74Bs/D
g4nwdj90H83U/gECe3PufEFsDwij+5rF17asLfmID8Ur3LuWCkd6En5vDhe3
tHmYDTCFf7edTcCWaboM/bTI2ZJ2flnk8pHprdfopii/z6WGQbimpaFgA+xh
GrJh4U7+AQnPZdlid6PPGuO2nIxTbaU05HELI2yUY/br1j4ZqkG0tByZKZIe
bFib+Kkhgv5WM3y62Ty2+bLtj4ADZzMPJRcVrIeUTWQu3tZ9L31rsaUTfCQ8
X5Gd4tmJntYRbyq3YNwjJ5wvj72QutP4V6E7qw5b76k7wVebm4T9xcmK3idC
FfH72mJ4dSdco8+G5MYtRJyvmnLqrky6kQzAI51tVw+zmWm6yIrBuEW4i8u1
KYoQ9b880Mwu/buaXFvC9t5t+CRiNnGmRJSwiHyamC2HzZDdiZ8Lmr1/xyo8
XdDK8aXH2hJTpQB3kaR7U7InnH1vSLQB2wIdVAVdkF/Xu/EdzXs7JEhOt6Xc
HAF6j1UptJSVb76cM53AiVTEf0RVu8JX2HLwdbIUrnCEhGgkJYVpFiNJoaVG
3fETy7y/msauxN8VXQkYx3se+inUE0miEpGu6LCsq3zNvkgV3NDlAykRa29/
Ywg51Gdz3yo7cr/Jv+qB7WuW7gdU8ZB7gy+s9qGmpan7T+IBJ2oewBAfZOh5
FGmbnJZDx5a/eAPwAKzGy/1KlNhxYO8bduItZjyi/g18gwqBAM5LyfdaNrZR
WY+2hI6lqUH2yIaLzyBE2amfbx3en51FbWSVcAaoBpw/TxXorwAipVlfYV7S
/mE4saLq7IMCHog6NOAgeNOAneG9znjwtkGIEOfbleCouhQFRuctdlDJUBpP
8azh1MlxyGrTaXJuq3yJajT/9RRMMKs9pyyrqFwjQ64c1snJft/Eoe+b2Lxj
q7SRFZQANzzPGWu3g2Vs/2vqB4RtVzGFdBXLBFN1C8QcOAX2mdw+7MKm7/Fg
lUBFqlD1UvYC70XB++UtTkDrJOKrq3C6kjZEa2BnF3aS1vkiuo9iPNqXC4xg
DpLL8/h3Ip1f1w6HuU8Ph3XpXHWz7wreIGv5J+r2xvJMYT86B2C1iPzNI8sv
Gx4AkCSMgnBhCzZahs1R4xf8OuCqP/aND8N5H9Pr6n6/KycWWi/f9VPjT24S
xi5c9iGrUqu+sf2dbYgOCv5HQ3OFPWUZ/+Ys/DNLOUrTVWThKjGEjNUDW3LW
swUJo7RLcJ9h5v+7vGLyd+4Al73EKWi/X0boznsszR0t+G22+sMZblPxA2+u
CnbdiCPXJsoLLc8nwPvCjdMvKypKW8opFFZT+0O2T33IfHuYhRGOn1EOCKBC
ACm597dc5GttuwhUaXLbrQQcz1t2jzbzxgScAYmZBd1aQO4vmuojqiFaamYJ
6aExZsXdyCuIDMVd4lDVFU+pF3BgkotrBihfkMYK6eeFPW2h7eEqtzpfpGHW
saVDP7cjtc8DaDfKh0bp9rhxNXh3vM8VTDcj1sQCinJk8kBSIMeyAvmDt0wp
C/znguy9kTynBrIj269PQr4FAjSZgtqAgWPD573F+VMgN+F23N9P1NK6ungr
+dsAMsq5GIdOo/qhg7/+DJo3Ghw7dBD5LfYLbHG47kKPCPIQyKhD8/dIHLCt
QEVbYf0OlsKAaPvwFenT8FtDMvMUbDvVTHrVzx26Hj/I+yZZ0FYe67kUl6We
YZOarOS6vWwivBXSBsLCMr3UBo7OXeuFr2BpPRiv0YQpMpIfWqkE7/A9lKZk
JoW47S63CbyFnyR2nna8I32HKtkidxAn2S41q9xgzEJZ/kkjQUWUrvTyRg+V
37CnzSrgw7uBeXwfLvV1NhGDvvLBVHAQbfX+ZQ8GWKYZ3BTyJB39fh5ZmPOO
FcX6V7BWoYDk+bSFRMHCgU8trXNVgljvjFCckoC3z7NRuQZuPbxp/kI4qmaZ
ixUhi6sBiupsBtGPh4SSPshAZlXSGE6hCfm5Sye3TXC+vy+0jcW7CbbXKI4O
5H3AP0PvnCs7n0v3y37cL5oxRxS4Je6n8uo+tDH55nNfqZRBtZeEoa2Ld7FK
jaP7G/wasqAQffsyw7li9fRqbi7c9pfSFUkAp50cPNbguFodTEF2yVJq9zOX
moPc71fcEwGRD4dnCWDzm5Z7OIhpGhhW4aEjCAcMotUZfoBtLuIcFgXtBdEo
xQwXg2kUDlIC7McQAaEL2uAH9LGXdwI7U+79lYHYzHRz4tLJg2rir+EXHNlp
8Qf6+k3liz0zquyVKMiDLPg2a1kTIYFD5xSKK6n4rYseVcc+oYWw/Ho5REwC
nzE/ku+5J9Mti3wyTp2H9MwCoYGvJmduOTjNfLbD+zcX+12r1PlU1g6fx6Z0
MOCXh+riyZDwKNEE57rmyRyNxzW+GIN3u6L6rv1IbuBsbf5l1g6gR1BPTJ6j
M2awRItwlM9p8F5YokftuVGcRR90qm7hGGRa0R1Qee3PX/tufADNQnz4JNLg
cxfUTHZU7oU+nRhwG2+KZqHOsWMrohRXlKO5Pv34Qo+eK4kkAGtSddFiYdIO
zAymCBpYUKLHrqpooO9vREVqkYG6E35+Twe8TW3BZ+gSwMcvJe14Han9OUHM
XKntarn2wzWlcCsJ4L9tmB8uBd5Ybd0+BThc9xwoxQ1Sr18QQYSmfOymu85B
gxknNQH9uM0qPUc6ZhA5jbgm/OSv/uVPKu3JHf1zHZdGpMtbQC+KpYixKV4g
9k///q4MZdP9QSQ/HpWKcDgvt5Kpkc7dogujWy1/FcIuWWo9baffvoPBZIsV
zvFKiGo+0JLIWHTPmIMDf9wvrSncVp+rtmTjshqY3TQYBG1M5eIRAbIH7W99
5O0gPfP3dy1F6/m+B77r9YAoqTrZXw9kEZ1enyeroosjbRZ3dTUlqUbu9UfD
qY7/0T28WwwivwJmhtPdizReYA7LL8YNayFX3r1e6zwcABUuNRxpkuG+CzFu
VYXR+twNPmcUK3uERbX9vRCp7MMgJ7b5QVxHqfOSQBgdrhaaJWZLBeMUyseq
fqI8TjNU9SOyqPW+CTacWdn2yIbZVQcZ/iywNTj04bFyVwqxveSmTk5VaZHi
dSP4f/v5ar3H7q6cn8Fq4lAO1DTEtZVTW1f2Lv8uzvnKPt4GEJAPoBmEmdHo
nvXdLr6jUTeqSQmPKNGxQrwwpjsCkmq5QKAambOld31pRtiN82QYr/+tdVJy
iD+Ls0vYBNGVeEUtPXvzfb5vQJkL3ZdrYXmvnrjth+Icm4ErMaAZcMwto/Mx
OHipjSAcuRBBN46+ozCUPbuH/353DghDuyr+gPS/6KX1PWImJRlqFiLyctyC
RyHYbbmWi9WOojzBpmOv6QeB/hxVz5CpaMTxJ0j2MRVH3qYbk1YGTXKgfZNa
s3Fc3gc2ZmGWoSS6/if32W+kF0cGvS4qtZUzXKtpyNsBnj0UG7CHu9IpiNRv
ARXP75nQDWUCsgikfirKG3VmtPihDvpCyFgPmWMxpBlEfOG7lKOVq7gfIazW
9t6s0k4GFYIoAHxnYqvkcMGPYmNwuWT0zC168CLDKd+Acw6hOfXIwxkzSHVC
jiRwCO0yDeSjOXt0gLaKBkxPIJ/ry1xjiMbjKEfwFxPinQ1XIzO/Oj4bxaiI
bcVELAOTUB55TtuHIwWYL1IfISvz6vdrO4bWmevYj3e3ltxlMo3pEWZ3/NIv
Wk1zavAWLI9bAlTLj+HoMv4J4QchTDo4DnWyH4vZojCBRGn20gZiA4IJWBzJ
av9q1uPvE+LjGxfcvlXY1AH0ywIe+ZI834uCPbLoyJVnfbpH5BrtTrXT31QL
5iH9UA+FMyXpUBNSjs1M95L2YS0QZptLqhoThGRaKvxGXcJWCfMeDOGbNPS6
LatMx+QKS4IB7fIK69x/omVQugtA1m1DxKZ4pR76KZ36TWNakxbQ65MhZPGJ
7OeaUAwjScL6wtds2IGmcdhxxCF1LWDU8f+1c+8DonEa5MvRZqazHva7fVno
qyECMraGRH352ljqQJzmgd3Xa3ospam/y8ETMsr4VWbwyk5wTyJsYIizsW79
L6EF1uR3yRucizDyiNu1Sqes6V18IOAaI1xTevFvTM5YYcg0ZJBKphOzTzpd
c0DyoHG9AnXUrjS0TwI/1qo1naTwHL5pHBfIXeZY0khaY70skT0+NbfwgPzO
ohFa+JpXkF3yR+GQIyFn3uA7tQZBgyDSUOtER2l+tdvbSWh6tVmURdCn50v1
+Bc1TnHWgRq83XKkqfjXXRXXRq26+TdZOr0rs05CA23KMIVbLTujqMAtQu65
f14EMuegx24sMhC0g6x1JMHN14a5MQo5bSBhqhmWUwuWou89bxbkG6qjbbnd
Wud6eEcjPvePCqGEcmi4Kr6c9nKz8xj2a47AX3WdXLsxm8qKJ5xb/tfsF4W8
VdB5QjaIjvxRQJQ0yk5eFvCX7Wxza7KdI3PLRCgjkcxQJnVAPuwmECMJ5vqn
rYPMhzFwuq7TC3n+frd0rcfabuufusy004t9mLoJC8Gz8JsXDB8tuCrnRXif
cV02wVSFTMcYqZkWIHc5+r9SXzC0c3xs8bwNNA865QWNIPrNoavw6Vk7WgG4
wqf+F89OaUfVwKdH4mArzbOCO1oNGQ//IBbpeUqu8xTv7isJ0HyiJqNZB/Yb
2VpVZjRSHchWrSfzG/ffqMsVJUnRRAnwSALZd4ha1jiMamZ7d3p/t4hsk+um
keHOJ98hnsjHquEyOdqsNTzUdLGodIzZSt5dR+9Ta0BAVzLM4Z7EboR/cygG
z5Oe/zllszRL+JOWERdJnQWXZd4yNG85/ozd9JtL1Cnefhs5ngdIEALY5Ggb
0G2kzVhJSW0Y9PI5MFdPq2D/KBVyrwMqpOc+EZ5xqElYSJcM5Ml7ADSdysun
iNchBpnOeiUaHGDuKNXtn8CrLpo+3nj8oBEDqUXbGarpQua2UO7nY+OU0/g6
VPSPJMj932gTQPv1YYaHBR2ZKXP+Sx9GcGowqGKZbJALc417qih3T4b/jVsH
UTCKS86z+eTfQMGX1yVANoR/YphgqD9+HgDKXPl9OHraYj1xHxXaT4Q2zzjD
TiZoKFqY/H0mz3f19noe7hCWwXeWhEw40C5GxRptSdb6NBElqRvhlBb4M4Qw
YKXpeuWBdT7qSZV++1ovAxtByI/fxRCbaIzF3CDkoG7M6hJWWFyGIVTKirAz
XbYAgKGUTTSttKFIzu3qBYqLIXfMBm10P3eT467O7JIgpnqOV+5Xe+Y2DSAM
Q/hyESMYzFzmOMriPNy++Ctu4fD7Xyo4Ij9QQgG90OK96FtN1UAz4wWfPDn2
NEptN2mwDhQ+bNbRZWGtsPJpKGSWlV7+lJBAkrOhV7cVn7/kc/QuSRW02j0q
GUTLBJH3In7srpZiQmz18noYB926dq8c3IQaNBWehc/U01QjCVT6MPNtFHtw
Zv658lNNRJnNTyfVxViIn1OGW3Q96UEAYr0JFg9/mattpoABfxGrxnopnK/g
cMmQXielLHAAYqAslRDvqzkz62O14XUGNX1p3cf1okWKOrOY2hTo1sq8reVK
ZrfXpA9sC84vZ5DOSjwe4gR3dm1df4hulO8DGxi4p6s3YO6PVa03NPmK7lOI
vM8YGIoJURdDOT8X03CshZ/0fP7KpWJQXCI04ODwDnVZ9nimd8ocJYAwkWiq
GGpIS0cYxI3LCevxQ6bJOuE7+5TeWyiUkDzVlsHCDeo+U75vhJ0oJ6aBDbgV
MLpqzglXVpFTUL/HaVn2kW/gY6P9rsEQBzUQosy2y6sEhm09C0IMRxDQB2Cc
6x0vojTOJYSjvB2OCI+dInphgdPeszNq8kud2hXxiTGdTVv3ZK3LYMRenboX
/5+ADxUCUcBaIBLykmPBtGUcygdcSckcMoiD9Lvu9ZttwybG5etk0PcZOLzo
+/JrwIOKp3hJS7pr3j5c+E7dmf9Is5WpapN2LIED7N8YqqGrf3p4vR5t5AuV
BFk7cCrydw1czQGvxTi7W9BGLdi2fGVm/zlCrxPv8rjAZqPJg2amYIA46ST7
UE2ughoN+13fFFebGIJF4E0uH7DCaxaa/RWQPmdtnvHTDiE8nx3TAVaJZ3ah
WWVz6hW9V2YEAkCULVpobkDOGMrK+9dXkPlz7K+U7s58eSDTZqu/GI1rgYqt
cy3+lyHTZW8pH3OU9/yoYNkMkJSPqQfyVsFNutrJMsGrjnJ1LqxiNloVNxZ+
curEyqxw+SpHm6+APxTdJBrvsnQjOMGcGGa5XmuivrchJJByQZGVDMYBxbJX
F7NhTOn9X9Z0oj81C7jKOz/10ASbOU0mAQo4fVTLzP9W8SP5ZYu9EkoPvg/8
YR2yHUX/kUoVJrDcWYKWJ5FO2L6fGGi+24LGJXpo0Ei3+VhUylhzRd1zi7it
7Bjq9TFYmJQWTbU69KZDbcdpKNtm6BGK2pgB9XajKCUhIAL9FrMVUm3NaOgo
aA4VWiSGEJoKGCKmFBexusOxMNLPbmr4Q8W3sPINCyQU78+PskI2O9WAh3Ha
vdAjvwOYXToanIQUN+McduJhoDXuE5L1paxxAdlW1JnSaFWxKjq/zcugXMrM
YSEfNGzBHOFi1ySXTlJb/QGQVH4Zxa6fAcRr6q58SK1KjqRulQrZklQ3Dpzr
PA3HN17XJDg3iUN+Nnw1/IAB6wT1K9TZtC/loJ6s2+tkhM1r/KIcXTXZf906
uPGOjVA6rRovCGpobHkLk61qp+RP3sTGhm2ZRFoll8d7qqdm/Dsir8PLqZZ0
wpe30LcHOoAoy9AnT3QKL9Crj46ouFc47EvzbJkddDM2CoYtOriLvseX7hPJ
cGCFmzhvCa53uW8Fym5pyonHNqD8p8QLx75dOVzrchPPHXaCZlNt3kvz90Gh
AGMbbws15qxLu7lYMD/tKUAZuoLE6U1iiH8JB7fiMy42H/4ogkHJW+lgVQ7y
Xf31RK/f7mdYTDPn0/nib0C69EcAhRXNqxFXQklPqozGsLwT7JFkzUyt9+5Y
iudF51a2yiW20g5PzgqyH0gj3Zy/XzQWeUCpjSeYn3oVF20jGk+hJYIBlj7W
2VAf+WTryawUpXPmvoeUVozce4mtzywOWKvat0h34FRgpqGWcsMxM6yJphzK
l3k7C5N1SM7L0wIwUyOII9W/n2RQYmcNovTysj1OPPv+6I4tfXDyEYqTg6/p
SoeWAJs/9MTJgh2Cgr8C6j6J0Zh4FFWoJAj+5+bK9Y7rckg+AF6eSRQ0dTxY
pMEr8NE0AS/p9MR0HQDZ7+madAYFQ2sTOYOoME3OQufbRbHASPWw/S+lsWlJ
i4k7W+Xxx1Dz36OTs5VgjL0SpgqkwNbj9MfKoQBYPGzCjFZq6A+IH6nyfyDp
7N3p77d/4zwZc4dVCJwFTSzVu/2db0KBG+X+Id2nzR6ROfDg///XIiaI/kQU
2aiKsmEgSf4/8VUjlz8x3JFQgqw7h7F0ENtI945f5WziPc+tidTSPF6tZe9Z
fIoKYIZDrq+cTx2IEz9xMopdOwULIGcgDNTJpxCh/NKWaLjrCImDeRYGU7gf
Dv3VDeTBAcIE2fJgDLaZF9AwzB3u6kz6kt+h44G0PXat7Mg1ZIbiGp0JlcvB
agm83oYhtYLVH6i7f05yofQ4JLW1x0orvNAHS2YeDFnmSM7hWSCXrdpK8sE2
m5vcH11nZHEe9qA1nHA+7SuMcxswhWsr+wJ72/5Zc0xUrNr/4qMckWRKQ94Z
0LIvn7/HtD5rYgb/H7P0iF+N0dNoUhp3DwzSlGFPp64HvY7Qc1fYWNNfj7f+
pLimGxmDUUOH8bJ1gNiEdDX9uEaqweTBqLV51fAk/ijjZHh5Wm0JLfYu+kTl
vBaI4qa55xcHc0bN3YkHIHCWb3iuCqXPOdEvAbr6IK2VphBjIPrTiUNeoqEU
6ohu8OVKmfn4EiZUrnpoyzathEGOb437I7eFSJIZI3MlDBdRWTO1Lr1CM7xW
aNiJbc3kAAgIX4vGr+7L5UdjP0P0iaX8IQL/xa5020pR7FMF8Lf1Yx09fO/K
2sdye6FID8kBoiEwdFpLPpdRait1ghuZmtIN/jdAlyd7QPWt2qX/kGaOuTCc
eMtpUlLf5dU0p79fALsAHRjSfmP4ieJScKolRSuD0N5CVrnWpG1rW0Ky+L+R
L9TZ0M7j1eKqq8YWOhPdvgUr2RC8HTFgfywA1mSYYCVfyEbtdkn6OVV/5EId
A9+73Bi6tIHwWcxyHgJcsdD9mmbIIqVL/tmhi8bb89nmnLOvIhMqNOD2t5nE
spspxpNYc6H/pASPzhXLMNwJLPJzz4yir449ebtwtqOGltD1lS69DjscVotV
fqWfE/REm7394hURPVzkj4+fgckWibwv92ozhtoZYIRUnZ5rsnqxb7sD7MwZ
W6KxKzBWPcw+anWxu5/3p6YYCSl1XCGFuq1YbaVg+Rkyg1XkNPkHgrFFkWCG
vC/CwmZIehuocby234p2GMvlsdOgAsI//HFpyRxq63Nly+Hu7USiU7/zWJVT
8WriDabQ3+KBXIctGSKZFwayaFWD5LOgNJn0+rZGV3js7YoWMKATYpp26UN/
VHNrAdIPv5YzSOvWYeKZ8jUisLc7c1MfiD+EtJ0CrHUg1n2aE7DIE4FaB6Bp
dDf0YsblfBXC5+D2IPAuGhOdicZikfUeJVggry9eA3qwifs3TrL9i0O1bdzt
n0l13dHMZs+o7Lu1HubG6nsNnTlvR5Q0/w1zggA5ZOk04Jk8Z1C3B6sZaYwf
4uokOKGJvyas/NT5IK0icPZj8BQa1zoeN9ZFTqiXxzF+FEJ89fvRpq4ZBEBq
gQcQZhQhBRWH0mAuwEFqk8I4kmb/3HTI6UzIvoWZu3n4YOqdQ6LNwuLLHGK4
sKVJMPamfD/wAvHnQTW5uV8xQJvNiudGWEWGyGt1AjH8oX/edlQqlRAAaS8Z
ag5quY8I1bNGmDpk11yDzdqUCeI/EYP3nN8fTkUsDVGTxxAJmRp2/glSVPrO
EM5an4KCXh3UJQ4gVk7kVv8tcTwwELSC8lXdQAVSX4eYFSW/L4oXqzJFSJ1M
04QZerwJ1BNM41vvL7NJ8ZMcwO+DfaNI3S3wIGZPhrXb9w8pEtA+jZxemM1A
YA93cBUsxn01nW0GrX1LvRvaVtpceQsxnP8c0ZTcsFxxzlfOntcog0EA1Sdk
lXRGe/QXiv7zPsgWcfeEhTPhRl8cs/NJ1r4OVSpwH9XJmmpZQ8bmxLd11JVZ
pllxtmlS1+Bd6ljA692gpuRLjdAp01k0UZPgzFRcrVQ7zKcIOMYsHCyoUISp
/t4thaaqg1nD1U2YVX2BrGdtOZudy3lRiSY5uwnnMkSOfned5Zz5L/Zbykf0
t6NzeTI2eFOHQgvGWHosD6gSdF7ogjAeLrKJaII4cmddbLMf2LrnLoGD72fL
CWMDXeNhJN4fUi9T1+gQDW9wpF2IuSE76NNT+EKwDxTn9LbiCwipghhcxoM6
kdXm9reDGYLT+JDNcHlNID4T/GWKssR7QzRw8CxStxWifWf8oAKkQhgtk+Tc
n/aSgw7TU2I53FnGx5Wqk7afpqeUhJttoJqBSlZHwGLjXWctAPPdmkKk/mm+
NSQhmJXoYTEnLEXOIl8mWogtXYnmWV6PHg42YNKJKBhA2AGrYVZdLJ+01V+X
z0BLlQizu4ASSf/USKa6q87crmqPyLJmJcSwa9yov5VMJJBFmIBt/m0JblSM
JIXl/PSglvObnxaZO3oNuUSNYsX9ZMTBTeccOZ3hRn7uJ+uk2HTk5S9uCt8A
PUQWbsDhd9AnLR3nlfpv3Sr9sK9rOvTk7ju79NFYFcJxqm+ZxzA0Pq2j7gce
cD0J+6D0PLyAzULMulG6jkJcuY7fFVZnX/5CDZcpswt7Wx6fFkJRPtNlMIoZ
xGT/1gHZhN0znXjrlx6boL285H7jytPMZw7woWYCDNIvSuUFxJT702f4HUS0
DaHDWZeJVG8L79+d5Rd6zeeKptS0OwYnlOSEbI+KcNcMwTkByrZ62SnDmNCQ
BMBoK5qvubemHponQjBHqpZ0mGug0fBM/JdaEDvYxuAgTrk9t/drw9TgWBSv
vCBuD32qwTlf7VuwM16oJbaqqbj8drfQSwIN+pSkpsoBr+Kdv07sW49hGiIs
9RIEAfnDygEPX4s20zFJAgHLDZ0bGhP7ILV/Ek9niCY/DYQVW8F3q+y8yfC5
nQTEhH3yqh2DS/93aZt180GasAcAAv3+TY1mupnenJ2774pvg1XMU9VXqKlc
iCY4aEsR6jF0eT1vdf9UAZUvci6AkJV2h15RnC8rpGF3RJrkRF6QU1GXR3wt
wNk63S75oJQzo97SQ1CBafbwUeQIKxxe4fnVb/FaIl91Fzu1vWciwAd7U962
Q6vwT7OqXOzvWaE2VLKNBLa1bQRuPmthGF6sZfNODqr3F/0aXiz0V+u1mG9i
vzojeDMPglqfi0IavPJGaU8Nw9biYLTmRvFax+S8Fg5FhL4SqiPyOa8+FkR8
vHugVcRjWZgvdtVEeAyXL+24lmOo+kI9EZoiKdMy2dV4Iffi6tSweRkgWmR+
qn5CkoArC6Ysi3CgiiuFx3Rml72OuSXrqp94eEbnzHKP8M9Jxt5IBaaGcwY9
87cxiSeCFiOswHTeDSoq/yOCKHxWXlZ2YknKCH9EqGXFKrbRKRnrWVERacNb
8oE/V+SVm4uEK3DJFc9MAhKVDbfOHrYU90jzkWmeOwSFgV3gtFfuOzWhUYPl
WueK/ie8U7k0FVLB3MT8x4omaSU8UGysaw2+2h7GHUCz1Cw7jDynFFuklaem
ys+5YnUbtx/bg7ZzxDQWNFOjl2L64gvaATLeaA1oAGYlUGXn2Q5/9vkPl43L
xNdn6yTjtW3PL5RFWpsC1xGLwTum7uUb1vs/03BRMXCCBMQzkQUkhyTXIWfh
dl3wz1wF7Dr+2Xac0E68t21aMyOK4ROFYQd+h91GZm0NQHjO+3U5YNGVeGfq
WfYU2GLwCifv4cHj5dEFJS6Dfnf36Epbpq2hN7xV5ADmiaZQ3T61YRZwTFGL
SoOLCTAh6DpxfY6KPYFfSdu9RWN4ZM35EI5u5B7331sNYo1Oxcu0l3GEqesb
H+2j+3gmidanYTiNU0rJHx6MIqT4UwzOnT8dHVkHM4d19RWYGJcsLHNF6kAT
kzdI37XEGsiSYrSj5u3VfxJaVj8+BKI5Q71hlm0K2xK46J7kZkr9WFlwiR/k
gztg6kksG5CXzfN/00tj807k9llN4dBNz22knQBE+T3tlTCG8lu914lkPisF
gtQAWnT+UWKfILvRrs8wTWp/FWTpJjvxaM+Yv2vUOhFopsWyOdSxjeXOYupZ
wozEqIpcIjqH6ZohRbKG9R5fO9706o0+VH8Vi/2gDHAPt6fHfhyHblacI5mH
oqCkqGgCW8Y3MXvochvhO034rl3Au3a5qB5npklCZpPIDYIClqDMf0EehUgp
2ECRb50AqLzD7tzTWzLtKFGduvw8Ly77Z62pi8MxRj6eidSvh5MhQX8XyQFH
OGUNIlrXFqG8LG73wovXm6y6hd0czGF8LoLjNAh5bSUHDAPM1N76opezF14Y
NQe1AmyqpxTNyjKspTEfRD8XLxEPUiKDOUbCR5UzGvxMsvpl6zZ5QIO7+/k7
gOVT2w4feSutpLCdv0yn1ZEFNhnWxzMEWdYjRXUiah04La+5GBEvWaU05/8U
Gc7+tffhsp7Q72QTzsTBzcsa3gWbpJqGc+NcEFpKs8Y9vnLtsSGIdtx/md49
dvCCUlV1OZXblt004leAk0C2CfBCqIxOP0gdxbMAQBHiJrtJ6vFDsBXMfG82
ulgV4AqK3c4YMziDgkR0jANDNrPpnv02WuvjDUWfwIurr3GL6ObcwliLxVer
N10yxLE0ixUB01dLnsaoaPLi0MFaq/DQ6lcZCdPL/nmQYralAHNlcNqTAB6J
fPtY6+ek8QPJC8QXe2riXZFjN8YbpjIO7PFmJnmBbRqtT9XLGIo9jzL8YuaR
yXMStIVCvQaTp4oUKPRnaoAehhO1EBjg5r9CzPr590tX7aq8ov4Or2NJ3qJz
VU9TJokY4fiS/tmxsUzeODXTrHn9xSQsrZkPHM8wwKKxsUfDuqZ2MNHwNfHh
VWSelOKHaU7Wo3WXd//v4jSe0L0qaVSemuV9GZRBWIlhVVzPPWSHCPgURJEB
0t5J1p9iSkgmn6sBjd+lodDAMvlMgoExGNZRdcMu4XpTk0o/nhH1uBHBA0EQ
E7aPxYU7fiRzmpw8QKVWOU58H0TbCV/Gs4lwwuV4Un+V8nHgQYgtgKDw6g+D
82n6NDQct2TrNd0D/3FzA0KqzvpIuoWI87KNguaxZYVSo/RwIVVG6Y1MyB09
R/tUSzya0D9SZ/c607iPFIb4PgboAtPPeg7+HyUOxUhg50upKOc5Jg99VPK7
cYN9CHPJaz62EOMNgWLTd1L5O+eFtte2fQ3cAJNfCDkES8Jb+k/yILR+1Re9
p8RnmO5zOJ4rXEQlYp82GVNxN0k5xyojhHNBHgfgpyaHJ+ZZ+P2yzm2bcT0b
z/hJB6qzp5QwmPfVjD35OwEPX1Fq0hd9r3Vw2e5PsL4mkulSjfaWsmUB/M94
4Q4jZRSB7kWhuz/tqnyNrBtc11lCAM+JzfXTcxrqlKXoxdLrnHu2hksYOgSD
9UaiidJDqd9OqoYxuwZWZPzK3rkpwugUqhVD6G9d2qDO36oUqI/OU4Wz6n6b
hiW8OBa7GW0/e5TLwEWbQ5FbuXRpmqBdcoGsNoNwsiAyeOLj5SvgI28NPxKY
OeQFGYey5enIeU3wV7ksV4+yMZSZF/94l+iVvQsU+7isHKk6ywGT+aYl/wWE
SRCCFJxULZTX2YuOtdQToHOIeDQ6fOep9iWFw5+HaDW16iKJTs8+Ff4es0f8
ZMbZFG206EQkA3UzB2vJGBura8Iy3JNxvwt+q0wjEhmMEf/QXIP0Iqvo8nYT
k3jEgAykmB3L8RYlR4LXywE2ojCxzHfG81LgcGIUx7zQ32GOhwTd0SOu8dNs
PX3ERfrEnMRFt4krYXff+D9zUPS7sqU7qgPDgiiRDAxocXGVoAo4OK2jOZ0R
3kWG54fPEqKEUMlRv24+JWfNspf+XluK6+IQWbKfnOCXJig2TWMDy8RpcPnv
MbSx+X9WRnQhUB+bKw6jnkOjfvz7inkg6GT8winl1T/lgSkG7rIv1EOZTgHk
y6TsWxXtCfgGBFbOaif9xskTLecE3zXw1qZ5xJOHC/WbAWkPhVfpTEpNm5uA
Ofix7MEHd2uJ/hXlFHq8Tmc5/VxOMFbFX7vZ/ZLHxPj9viWBUYTYUAqH5Bsk
tU5Y4J+kjGTMOFb5C3imTLuwJx5c3RBKhBQ2lQEetvhzzAvh2yiMn/2BfiVc
kd/JfiPNPxJ4mBLGhyloKTRRsb/roEe/Nymzjrgnget0TjHu3jG0wFczIISY
Jmir33TvFR5DNHaB/Oib/Xpvng6rhrwT0Z3HxRPSY/V5Ye2G/jEjkg4Mq5cB
Ic/1dCFdS6GeGWDQJ9gL6F3bGzxSLHdwTBV4lRsjLD84idr8FobbgQ9L7FRf
5lldLQYCQuirKFq3xFwQ0xPgCgCaGgAI6IyT3enNSb8oNBUo8ymf+w5DjYIZ
z+oz7aDM3n+RrxNxyBSOGikSTq+h7X4jEWNVmBx3XYeL3cIFIpqqb1aKTjMQ
0+eQyOpgjBIsc24nleq3ZWfJYSK5BeZ+HgnEW1n9cZr2FRSOjHqjBJVQ0+IQ
DkjNNlEZU/ECKkeFWztN2Ge6r7Rjw3OURvXzw1UrMhd1MkVl4K1RHMrfOh5Z
LY8sg5HO61BbxFLN/ZkE1cJiBLEg/AQahdPfMeNIQ+wbb4Kn6JHrzaeecyYm
BOuwEJ8BWpXKPpRumgEA1ZDAmBUiIfzB6iy7Dtz/03XWjBejMeyJAmcti1sR
aQMADeaOKnMT4LLUa744qfF/AEBe4OJJbvB42pugZXHWzIt4qMNvq/u6hEz7
iMLMUCUyPRIy8lW/LR4/J2ZdrKoAyrdU/ujQOYbaZIinixXzD3noFeknh3vm
myBZaLGJcwhPhcI43MDF3ATQ9p+e1oqknFbdRDp+3aw2DoY5H+irLUNGTSfw
aEAAvhKsNG+e+uHD95sUuZHaJqcdugOYkxuVF/bqZk66weDOL5OtAp3etNRi
vgwURbBeO+V7Lj5pFoBh3UvkXkZefCbwppB7/ZGf5egDiKhAC9fOihsw6LY+
7bpXfSrdcyxvx+DKscmdSwnEyss02kUxSl82RVo8wod6C7ynDluhcXhUnduY
Zv1P95u1p/5FIhykeI1XS3YJ6NgRn6xQpAnLDIHBIDgSWFvDiHngisnQikZy
8eIgZl8DAq3zFAARjPzIMd8jSmwF7ltyCjW2RGl3z3K/ck6bz6dN4EVeCgtG
WyhEj10kK4vEHIrB5Nc/emhjR3BX+RYW119wg7wX9WhOq8IvCqlE7Pm6ZpUA
jNIwoia2by39bMLa/yJExuVS1Dn5w54Vt9dyoBp0Zek2UQAQFVwSu70qnu93
Wca2A3Zf/EzwbndM79sKZUaI1ldq1LgYhwp/zR+UW+X2Kw4zlHX87FR494sW
LLEPNDIeXFC23lZMwGGeX9kvEhK3UdobBHMhzTfrD2qaOF8X3aPvdGHVfo3W
p+KJBKdkM5/v7uXVYetZPqoyc60Gagy4bz9XjtTBFFyWC/wLY0IoP1/0RH11
53xepfIqE49FSbnqvr4zDX+AW7ENByobCZAGUF/DASGd2DiVgzzEM2HrFTm3
RWZVpxiUrIN/JAoGNRiAiNKXPiBILLYzHP30rdRFbuW2SyOwXu8NBS2v/GLL
Hrpr72CModq4z+bOAuFn0zKM5fYZiLKzca2t1K5qLs7PsgLWkDT806ilMUbG
corefocOrjNRTuqSm5UE2TKlQwXdY2mOIYHx9FkWpD0PkeI0LGbETNdn78+v
11z3I1/0XvpCuuVjFrgOMfcjSTuaiqUmIczsf6DdIma3WJlZ1LPqr46Wvhb6
F18SMs/UaXxchMnfNx2FpA97h62D4q2iQFed2X6YZjPuF1tSwjX0Ay7HAOnE
HQNn2MxIwQ2jfrcf93BxhJYQairCje+/9I6XExMGLKot99hC7csCdXLyBIKl
OKv75Uk9Z8kslQJXVUE7YzB9e++D1TzlW961k58JPRdLpyGXB/Q8bATxq0lQ
3EcRgh/ZHJcJSQA8BZLRKnH4QnE05cJLzrLOAeevMrWLNzEFrqDxdlm+24yo
nLSSWVGRbkqUyiEmueQe9eBKJBLTWbennBwQHHqvTgtTCh2PcxqSOBEwfh0U
SD5xtaQWCUKNn17tMM+/d6MaprXd9rcMRrdOoHjMLxOrNws2oF8Vsb2l8XPY
vHhZX9H6KY4oSyEzwkeQAW88wVu3Dynk/tM5iv9nWJh0SjzjVPU0GtvJtKDq
LnXEsufkHPvo0el42IjaHmcPFFwqSbOgefIpQVGWY2Rd3oGFiTgoa9hC/T0B
+n1gcnxPsbVX7cQE2DVq7PPNybGS5wToIPLSNuzRUFfC1h4oLjbo9F7m+g82
l9BVcPUeVLhziVDLWnyfOEJUD9Hn4mHGKLNnpSf526Qe4R20nztwG/9Lklsm
F9q2nDH53rMGOw3L7X3KvWqfqIGgs4+kY0dTqU7ddI7ELyfLSIdhiziVo4In
5fdJqk8ZzDxzrYCYz/6nAHRyfiJ/gU1DRHpA5apMnJeOlCfkqrSyWjooZQx6
Jd26vyVg5U+o4xsz9jqkFxT9oD3xyU6pFtrjR0ekNvHEkbAh4DPMgykxfy1i
pmB9aYuZ2cZP1kHWjIp3uHfJbzx6wT2fqSdcQfpmohBDcVTyMNun6Z8GMi5j
myQeDwkj4jvtlScXiZtr7GKKH5nO3V+jumxqIRPbagB8PnCvL/gAVEAeTKwf
lD9+4P1cJIRzRgbr9UMiuXWx1NnuO3RFieS0MvdLwfKo4+5bMHLohOjvQIbC
f/gojApUUnd+ntJezwbJf143l+OuUdbRVmj8pu++o3s9KcLsoYh87UJYrzvQ
sKk3/qL9n8oY07WUyn2x22uCdWnqRrDIz+9G6Eyoh5k8h2I/tPFXb4LFGIvZ
YLIAlF9+J2V1aKy5OhOsU43zvbkyFy9JhuhIKAhL8B6l7iAaHAAJ9tLJPRDg
iMKDj7bU+S+rzY31HUBB5taTZ8lhf7gO/FdK9KxinNmbgdYQhCAYDEaBYfOf
fW2zn7JmKcJ8eRH23pjR9zRfd+5HfyMzs01ZVLSfk2fmrX/kOBsZPMWesZVj
3lO5wz0EtympPX3mWyH1z6Zouk1CXZSAn4Xtm23Ndo0EN6HqnA2+TM2G/FXf
GIsBHLZNO7nn3Dyt+285D1zHaxgT37itnUdliiCjMMhqgZMRW18u39DKH51e
AxRlh7+Wx8usu2nJdNZGNSGUtd8cAFmk3zBEhwgE6uNpmvnGpfYb7QxmgIlN
gzcdtc1wZKcrl6YTH+lV77Pi1XDbuAQ/Tg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EoXTw+RTC7EFZqFep+IDS5L5wlQVfGgL1dEb3AMs5NqU4W+V00A8Wdsq3E6xsiFUR5FnEaDb1EK1C/KBUkdq7rYJ11OgH5o9CIemw5P+fQMYvhLRe2HqY8FldaTfeHN9VDLVTQg4rPeeYpb1dBSlnxnj8B/Eu3rZhjod5gbGTtWeTG8vhVM536+FozyGpZInesYkENUGAB2DFcDcvKzsNZ6GvhmkeBEAdMojhWAzxKP2K5fp+QDNpkK/7xN6a89+mOmetY4Eb9V0BXG9ghrYYkO4tLYFiymloo0uCne6EF3FJbV+ZicAcGcjRRu/gc9A4rbtxB9OkY70GxIWt5MRbx0C/zvpZM2+DMDRYrVULMkFTSPCMpnndMM2eYfUlyQ4aC7nwsIFLLXI/7AAmYxzSS/iMse/6NFAEeBlgyEShb4yp59g9J7/BOlLKpBByOy1P6OV4Gy8v2WQa/HScuT4PYi//7pudoEuK83IyP4WJC8VX1fEBbT93br52TToXiA83cZfi/0hPOQuOp+0DfOfbus4RJFGc5hhGGIl0J101NW3vfED9Dd0IFAgVnDBHiqydf6CbdVQqg06ao7VG9W7d2tgBOM3/Pfo5CBkUjtQ6Ea7pKzaRK9cHft8Sw1NNzf7wJvYrULtG4sPwJYoBruyKUytCEpbS/ZNYmBnQ0OmpN3Ou4OV1sH3B+TkYhg0YauD+/lTqFvc1wQnTW9nXBdP+V13lH6DepWqLFZFvidel2oprTRrA2U0PTS194cjc//QY5grnzxboaJcLYhZBTQUPNd"
`endif