// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wlsqJZ8S3SJ/L71dltdnYcTotpVbC2WNDIsCrHKRcWKkMNPCL0txRSED+2EJ
IWgYvj1HxMIAONbT20vUh51IZdDhEDX4xQzdq6S7O+JkiWyuBG9B1JyKOiUE
5KNB8Bn+64EyRJxWvDbjnPqD2x1iuAn7/HBwoLFVlI7jIB4dZxL4iht0AKCf
0pmmY+oVLNYFCy44JxqYdNG6BOTatX7C+x5A69ja7RgqwD1RSToTrvw4Tbwc
ABMg0EpsPDHxRM2kjCv5wf9okTRx1SE/pUS8ZVb5LQSthoJ18IvWRR4v/KYx
dnkoo3/Fwh5W/EBfZ70AIk8uWHuC+LBliK74YU8Sgw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mI4zSYDJXlW2xeEOLPae26TyRjn8w2uBKnbG5EIhXQQZjmPumpgOd2kvSsz2
hV8y+IkePtyjyd3bt9B3dGhDM6Cc2AU3u1poQ9TR6VS73QgGNpyEIkIYup/q
ELCFjFdLYEVGzz7iENpj/ZYjM8n6umSoHfl7qh/7XyAAygup7nISh5ZchZKj
DdR5PIwmb6S2XiYohuZyvTXofW/N2URFwV7a/DAJb9o5z107Cer2NcYodd+Y
GATnEaN/PAdk1MJ02tghQcClQLwaWN+xKXNKOt/norRWWykg/QckQbBneK96
sqOgCszZhFbYzan6sQ4SmAnQ81jMB6TIzaxQx5fVTQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FE0Lq6Fz/0JrQUpJQjeaectFRpmxzKaFJS2NsXnIjFxlo6TGCU7lBP1oo2Sa
WjR/q7LqzP9J6npSW6ZtIjkz/TAt2fLx9kdjeGp5Mq5N4HakGSJFdRWcIHID
YGzq8vhCHBBSwwBlTH0Yc2nVwPH+LJQSOSyTH9C6/gFMMQdOYJje9RY3KGwi
/k11z/kPQET2uC1TMuJ7Erds92DVWAUlBSIRgBoKIkBGunxa2MaJqkekDsJa
Dp4I4nip8Pm2iwHWNZOvH5MyOAeHn4H0+kIscbNvXTcGGdN+GYR6TI9yoned
BVHYsl0hQZE9vzJMvPMKyvf1VAiOPdL88GkYa9URWA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WTUwUD2/NJhNvFMLBzciR6Fy7mbF/nDC9pr28GNIXnNscud5jDsjiX5jbrwU
CvUebBgF0CTmY/dZbMRWFVPVEdetuI0Z7v24TQ0+VreTc+AC8MZh8+Q6JiyK
0168c+y1QnZmq5OuhUQR01o0bl5uLprDAH0NCqMuumumP2Rgc7vWb4PneRiU
5wILhmX433ytOWJ4tlQUwE+kTkHJVzJX/tFBFhsWl0JZfwFEsTlWWpLJhJEu
xNfJ7E3Nsyeq5KteCzT7j0kkNfvMvwt/zlRcLSK58JRkOdpF8ygds50qax+9
k/eTQkqWdk/I/iCe+yWZUmjhRdhf+hHeXr69+7Pnbw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T92yqTGGTiJCmiKYCNPVVIsvmEuRXikN1/FtjwP0RSDs2cDMzxv0j7JzlPOL
qEsaZ97vRExIrZQXOwyEwUwqCj4CaUE24o99jJl4ZVCmzomRtPLU5EZQeXYF
joBxW17DaEeB8nven0pqjGv61ShCGi18Fp4QHAIP0JFAL8I6WCA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sMi8kkPnsGItkiDRKZfZhuJUUpNU8+kuNkVYU4iRxofO7NRyAuMhSroSeznp
XckEIYuEzPk+yJyJalJDaYMIvJd9AY4U9VPog9qzNW8vbREKaBqiOdYQ064f
js8NoAc94soKdLDAX8/xkPXwf7P3uR97vtNT4LZhy30k3YdrjLSOkNyiyzbN
hp69d1sud+v+EJA9l7JVIGNt/d+mZiKujV7y47NG6HZk0qQscLbInxy9/ck1
QuGWCeKZYOYR1S7OU/+4re7dkmw60ddtYpwq5h3icz3T+nYbjzzIkFTs9P1D
O0cM6IjKaeXNr0ULmeQ175YBPt4KBVaLH2nFbBWP6Ns2MST7uQrQP1+8af0H
auxj6/XRN1RR7CWy3yskn5iaC4dXE5gTKMq+N8RmvU8hmVEaO48nn5axOhXP
+ighGUv0O2T0GlYqDP//8+NZdSlCuEEeY1uAfN+6g20iHytqyeyKglhIwCR3
u53mFkk1iQPxfhSAbWDj91vsXxG0XgFv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f4+7KcMr4Pl4zFDpdBZ3T3PUf2t2GfiIbf3E9bjuo7fATZCBm/CeDSPqHmgu
pj9HCKBF4MfL7lKNPVaBna8rm5YYjbaVjDkcxm7Jq8yy5m4S83TaXgIrgCpq
i+ZbYojcdvUQVakWBNpm5Y3yDEJusuZKpo+ups685tsXJNA8Hys=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qOp5fwly+UEQfWHdEKudbc+h2u6zC2iXSZ1p01bUb8DWLxEPV4Q7vrauqlox
vYyTpxastkvbdw8/WUxCTj0BVBjF7Nm5JvdMVWI3t/lbwru1jIfIIy5caLRc
4p0+aqIRKK6N1vBBVcitd6IuHTXRfI9hUqDVE3bfhdCNhGPS5Kw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 76624)
`pragma protect data_block
pzlQi+3jD2YXVGkkrMqavY9baPwkKe+Nda2TXdYp/CYsj0VF1DpJPEcFxj4n
gKbe9eCnIQqUqWE91ieVM0ACf502dkAXgtvn0omffhLf7fVatY89KJ2SQTJ3
Xy8qOtHPmeWjzOOr+Wx1eOzqnIzn5Ll9i82GWDN1gG7kR3QWYnvILgao1U/O
q/0snJJaDgNjxSYueTol6nVdEK3Gm3b8eTjl57ijcNX9YzsWx8ZfPeN4lX4V
04T2zbq+C7jnvwHUuc/7IVnDgGLEjCMhlbi6+eV+5qTPF6eZDOZQNU7S606k
lq4zOL4fLnyol0SU6LtHNTAIvcpdA/oFaxwjr3NZesstguVXF2sXRVeTzUig
6JmJ0nUHHhPBTvN0QTCmFd0DZV/UtcK0yQuiL/lWCdGX5gLxJfwJTe1xlA6H
kThShNzZpBxlzm/9vMusYK4sfCFwCa548Dfq96A8A4/FW76YF40GkvHJRVKb
iePPG2oodDts5k36bKGJCeq+nmyslerxmc54uLporpjRZdy5K/djFxO8Fbbg
efv1VkWrMo/7tYJw7Xk+N46fAfamNGtyr55vMFs5OjYpsuyHOhXP/g93kqfS
tffiTcWY/q1bQIa+edmLKW45TDNAtPRQBsrph92jLlnwLD1goHvJ0P1tWfWI
wwp21LGapB8bTipmJKNs1Oo+EEF056AwgiBnHjH4lXLZC8OTr5b1bNsC21Ox
97vFu6ta/E6/6AW7JGOZ6MNU8nkdowbKwH7j4ucJb4zyi2KZvNT3Z20qCwfX
F5X1heqO5pai/O09GlluSCFLBDNvrw+9bWgYEzH46Au3Hwvnif+A3AhX4VdP
aoI0w3ekRAfrg7+WUO3kR2gaGwAgploA6RY/er3sNA8Y9ZcNIcl16DQGhuQy
m6Bl+CYTbmDAHdh2VSHqw3z7wamkaQRSex4zJ6gWqVTU/GYeAy6Dk98Gqxcy
xnTfSkkoapsNOm87NliPAuQ/68fCOxWaIRCCm62SI5WG60JCT2pOAcuqoCAR
dZM8nXS9e/g5mwy8SKt2A8X93TBjTTcx1ggga70ty2Ucamb1/J0R+eP3D+SQ
JrVV9DfhU6IYDQJ5apkK/6RUDlmEt8h99qtaVu1UTT1dPWyhKGcp/bp/Ko3a
TlKeSCuYy1gIDRDPtWwbgMSHq+YFztEKJoTOPvAAyBWfnrrAFGgrFii6SG2G
GJ6TMzOkbQlBEuqluCrgwRzuox96682vYh9PPETAxZPvAIWGqO2/j1zL05iQ
Ypi1MMU5MKtnDTsmBzgyktjQQtOepm61bDipZXw2uisaBiofp3wKKT2NO5G2
zKgLPYuAjE+heVbR2VoQZxcLg8YNzq1Fscbldh0WQJX9/fdYOZxAGaPpB3Jl
HwhI8L0bZgKARJkzYE9pcJZ/oegsHLgqp2/aAwJR/E3+c5Mdpzq0NbngyhM5
84pm9ELCRpkVa72+WlY1AF1xjA66q3AFzl/M+m25o5t43JT4HWHZIEy9yERw
gTHPReLLZWOArQl6TP7skUO9oDtcaJaKyF+omTvIdm1axF0HebJm5xFeLf9G
5jeSQhrpox32/3eXHJa6pOXAY7MVV1H0a/yZAu8BcgM8VNs6I/brCrwx1biw
MUttVxbJzWPCPVbkUhm/GuSo/go2bY7zFxp0xBC0zvSi9pijJZwsBMb971uA
trdf0bJxc9eItVFY9sgGWgRSosLzHXldPx5iqxjsxs1BwYNLRHXpdZMuTr8Y
D6soGLldGntyXcvFqsRXUy33J7Elvqtqkf7YhIGSaHQQQRU3eOmV2MLIfcC/
o5baMt1Ms1VcY7O3xkYNVX5LquGx5u5G3g2EYESDTS5bIx7Zl5ZaQsFl4ywQ
FqfjFZktbPZ89KYyRkYRmV+6IolowBSeAzWZnVqe+PXAltD0Sd7Btr7j5wPF
R9ePhLVFbVMZMpvLD5rrTwUs49uNxzpPZsfYhqV2/cntKaCRybS4V8ZWhwpt
gA0hYjiTRRTuY56cwY023VXvKmc5KOaP5aYYp2KRTNc5jFsh9gK/271RYTbZ
Bm412GoB1RUNyHXoTQaxr92tST9O2rSJxF+Tf4A5RZWvS98+XOw6sd8QZnKK
Gl6fvU8woOC1AXSZ0em7wKCehtvKXgUPWVlykqrICJH2LjaFbFUtTY7ijVFR
mHFhwuavwErwezOrl1fLKxUbkHhpDDdQj5mqxxOeqmM+M1Z/DylrRI2oFf23
Ju5cAxtaojY+wMVP2NXUk2kSMOzL4ZGjNd7SrVki+QYU4bn4ms3uQCoqxLCX
KM5O09Ks+MhvDpTH9Hvc8+KSzPmrYSglDAEVqSdFEcVQxBSJwR/AWVDAra5M
mQRs+BKB+9gRyPeg30ASRAvJdYxFmiIxsnt+IzwyZ922kPWTF5mwk/DB5fnC
Gy3/20+/XtegodKNR9hKlS2tnXAyjwvpOTqacn/A/aSiWD9lH6uSx9U85T+3
FU+yY1kbNhbFKWUFSoWz5ubshzX3azAt/gG6WLMP6RS9wua0n2hwPKiW59r0
H7V/ewxKiTFVikC2/MWCmsm8fukHwizJ651jrtz4ZEcV0OAnJnJbTgjhUTjO
KY2sc/ZEyIK193/9j8D5R0K/kmHK89RKacYYbUsq0Bwj6ncpM5wiMe8mabxw
I+KmU9WarVN6JswDJJdnKqy5UqkbnQiQPe1Nqr1YevYMdUy15iJU53QKwC1l
fHur/v0tuWQW6xvIPET4dFckFEX/XN5bOHIBFbMDR59CcQohhKleZYeFhgI0
X9bKG3mRNLVMjBfrMLdyb2sZvwh2dOpSZNHVsSrQ2Hsxs9NQRqjqw/nT4s05
NjWARJ8AwGELHFpG1PGrySBZr8Hwh3bzdijfui+5+9C6QxYwFVwOaoH2SFOf
zTlI6GGi6iTvGk3b6zHPdOXhQvrzR1/kQXrFCgEdoVC8zqJQwZUqpVyd3IBY
Xh9wi6O75SNw9b3VXdzxSxa2Vm2bkcpEuf7B2Hunq5VNO4EUq6NXjt+s0txL
YWkls/aJ/9TRhP/TgJNTRM2kdAIz1Ie6if7A6ewBqxP/VHbrUErbWMDIpSjS
Lqo7XBqAynrWedvqBKZTlPF+JRpXTIicImrXTpF6uTH03XjiYMn4U15hTz/Q
AY/H4LqSvCoLgDScoRKy1/EnP/RD+UKE3FVs42WZk2Y+1VRcSRH/WRz+lmeA
DisBhwYcSMKbebVZg9sKlT2Wzv/NScW3Bo+M4UwQesBvzl3fMH/UG6tF0KED
5vkpQKUnmtF99dvm34cC7cnolg02Kch+6ANRYfGJBlokoDwSSBqqAEgR/HL5
68dXaObNPQGJxrrCbel08n/SMF7rLErVtdenZY9XQGK6PKgCE/0t4hd/SlYS
TDrIyhG3r4ijH+iAF0VhZvcjaQxgqjQlRgriz2lX6RCKaRojypA15WL31xtO
ZmmaVUOQObqv7V61ZxhidNKHl21cwEHka5Vfi0D+J+C8QTKxgJOlz3Idr9AW
fpy517FeCyEy9vDVHbK3JJjJ4IC76PHB+KY14FDRELVKXZbGN7ckU7Zluz0q
rG40PtSt0LWSzujuwm7xbUj0rSeQ0CC2don7QGwa7217Pipa0GeULCXoLokP
Ws7L5BoJgdzKRMBRnjN58CoVtJ78NriYRnJKy/5WlNhDNrPKp09Q6lUoISgE
WG+54mneMeDA1y7dgd4/SQrYBDa+9OdW/X3e4czVCO8Zf53xcSpy/9GcM9JN
d5rENdUu/4qhkpMVFtvpE/nYz9iECqBEMs1pUxVmBDo9Nzyq/nh9LrT38tnf
y0gNyY2VP4xb2Kk69MrF5aN23C8dsvVOnAs460ceM8U/4Ya86DjbRbGX/KeQ
ayVknM6ceyVOrANbLGvsG/j4fz4Qt0R+8l9di0w59CjFHZ+oJzTwPBmOFA/1
lhLIc0WIvtcyKAEtqyifykmJXFS57hWUa8Ty+kGZjThXSAoFnEYtNJdG4JzG
HLpR7udJKfj03PhndTuWMuk7vHVAO3YlkSew/IIwmdXx0UaXIhKDz8p6v6/r
Ok1O10ifRF8Emwj5ib8EensMoPGzg9YnM4wmpvyKuENL1tjzUy2J9+vbIymf
3QEf3WEB3p2PmjRd9BnpNzMO90YR7k3oJtKhHg4dvhf1aB/gaQ2CskEO8CYV
o+XFbYPTRyOkwVx2xTrjEh1B7MNdSKbHEROPD+ghfBYgbX2G+o9sQzqhp619
Xpp5gw8EQxWQCnXnJO+eGGzdEIefadHrUcTXGgtBv8NEWZtB3pMwdidU+yAH
kO549/CioIWkQRYkzZsew+A33gsa416n++oE9ZrJEnW6lihQ2AX6+KIgC5tV
iS8CAyjHt+PltQpPx1ig+hK9toA/3qDn+MU7AdRXVcSfwTFFfMIMp1Hn748c
EWRwPCee5PLZcposuHbOCb3IOe7JKjc0hWD5UYpjVTnFngK2qnvjpq4/1zJy
KbHGBSaBjY9dWrDhoaEAd4aaFHZ9m9HRG3TqDN4tcAMkF5oUb5ZyPVpKFL0N
yiO/2w3ZBIYFTKuHuj3AmrnvxoSx9t3uuIWZRRzHDSuXlhxzArE8U513x/Bc
8ByvMtevapFgf4UH8knj/iGqBInMAPHWYtE8XWWsq+rPyIiGaw9yoiBhXF2n
RWKJy4iZJVRvlZJnBh0pNjEwjIhiiu3sLIDTlfIk7FmHN/WoC+v5tNDp+Pu9
n3OjFJ8lmug7+8zwIsiWpcigt5w+IXAzlLvTDvHneReQHKudnRXZhyW8j8o0
gT8eQdb9+8+AwJJwhanPyb8fQ/j6wqBR7XvWP1+ye12t8ib/DOA49GMrW7tH
k+bdHcLluRrKknhzyfxH/YPpCqwcnmCbf04zxcSgKD14CftAH/DgkGQVHPq+
m0jm5vaZcpN+sws1V2uguuRRXNdsCm8ZJXw2O1uuOme7dWc15WcyyeQinNSV
7jUOFddJenbBy6PAomb7U3zdDPG2m97a8nZzrvYs1fNYTMujdYZ+Qzhlfy/R
sg+WNNb1WHv3QJ7NqVO1lsiUQ6RFVpHyUTRr6t2BPEo8GYpo9qEJ40eH0uZ3
EgCTe8Kx/Q+ah+26/pTFudEiRmG5d/XEmVN2Ff8UlVmMAHxkEY0ATxaAmu59
gP0xRuq7rDGM0g0sg34mLiDOVB8sDu/QA+zMRkELHKcb5Mxn5YfNagoPXj9N
/AiFs9qbr3Gh7ltmptdSqIKMXmc9qgNh2RyYTJf9zTUF1FOxF38tmc0R702R
6JbG43EadJ9S57hJLQ3AXTIkBqS8qP4dgbs6ZSQsOEuIRhh0Oc/Heg2Di0Tq
ipChEZEBfxquxvBX0Mqy82DTEIjcWwsEEyAuSibS7Dx978i0FoBJVPjAlfK2
MAdhvnW4hEnSdOT/N+XNpJZ/ojGo+ADBk/lM/V9OtMXUEq2xodqTwyDnsZNy
dC8lumE5tVlLYq44xfhYZIjcN6p+UGfUT6fWBgRtM8Mn3LJuUaZJAIc7M+DM
E5vQlX2+dRixpNhPPvo+A6KdeLVxkOUEDzRJ2aQ3hf505WLIkQ6lfJo3PbZk
KBCib9zE9XzT9Vhr+kT3kEtYzECCwr9Xd5jPTOo+ha+8trdcz0TeUymRJTxO
mz0XuDsznWOVz18Na8UOdeZy61/iUlVqWiFfi/drGVwWcx9NGzWgpVvF5kfj
1+Mm0Vk7726262xd041aaLNR5j+z4NGxmbQhFd/3yUzJBDVXs9xrSHhxzb7t
Lk4VbWSLoZE6OgQCkXrslDpNzm5eSpzcQ/8xWsvlxKES7XYEm4yKYXDpXoqQ
ilJyPytSLqrPn9zz+LwCJbc0Jgjb5CR32jsAIAUQq9buO17UAVTk6ZNqrHNr
AcblVmATJwsi5Fl9dnArjwC7vhoAl8/K5+GKi+U+QPoYG9KU3mDazYwYpU/0
D4QWC2w/ZexA4H0mmlhn+w8aNeirSUTjlgkxQ+Vvg6UvpYv/REu84UgjJt+d
S0i2UaEtTCxTLJocpBdwCgmbpdVq4chyJKPE7p+9xuGd/+3RvP/vveM7tm2f
TK5fh4i6dMNbRDWntym7pDg0bWH1u/YX/E2OD3jI78XwWWV4QEvuE44JCHGH
Wg94GTX3g57HW6hnnFBTLXffOl5nerjB/q3kYcbuT/UhuSWC+WwfqknzH9xE
TAZL8readMJEX8R+XlWjOBY5UFKV6TNWOeiwxB20ovlrdRRmI4lL1AixmeS3
faOwtdmBlZpsrvu8cKJCDE8KniI22RXUBjG9h4uQIYxP5ZXwTvpEeQIy2TGO
EiPw4oVLAL/CfxPQzzmww+RM2r7Ji8+fS+WspRt3hVaaDCdCLhSKMWkPo+Y0
ACBfU59O3VL7qj5JASSZEH24+FgcZBMpKD4cMjlNTdjqlRhIE5CVs4TG85ux
XUm1h2QBMC48loWouA5ijtVneR15J7693+EPt00hfdCYmuQ2WsybWXNfrRkS
/zmdQd8TmEvmTayRpb5A4zBBW+Qrqh0V/efl6y5sABJG4ZQm4sjfG7YyP8Qx
qABG9cvAXUhuGW+WX9cxAPCCzPPCfEl4gXetsrQmCrAVNIlscVf4QftzLCH4
/viG26+YG25XAuSi3+RSzhXLATlkJ8Hj93Xm+3y+Kn55kVGpz1mQEdDkedny
qKBXvb5wW0aL7hrVX5S3n6Ec6FYj7NzIe7DvuQwNIH1K/lyzmT9gBJXD4Yuu
xI50A4KkK80ao7Ygxi3Ax5rew9rjdvMwvXQhCi70fNgsEFFdq/Ciyxg/InqQ
HOzQkcGUQRlXC0fMn0xnSlEcrKVr1uhAxKFWBdTvxGQY3mQ/ugckvgNPj8Js
QrsndxqlDfqZvyqfrNGhmWDxMdvUYwcXk4iXqsoQNA8dabwKhqme+7prdxBw
B5Z5e471vTXAwCEhbGWQX5/mwjFURRue5NNzliygoUvmeU+OfrSH5fqC9uaX
+RbOD9BckYx8Sh37IBZACWZzgdvRIh3T1iHsN1rgq6CkyhoHEjJcVyt+5Zh5
ba5AM+f16qai4R3PMRCTppDHDINwuP/Qfe8IFPDdwTEqd/8CxTJkn+nfoTOi
+pbYQk21Ky+51p8A7L3j9btgxBQR/2mMNIxxBChxMA9WKw647l2suOTHbsYZ
vCmf47Jv24XLFkw/3A9mJfvGYtXuAtuH64K9MKDeTkZnieV03yC6QStcJ2TE
2Ani+rsZXVfilz/fmAM1F/RgcPwgMgDRkTlUDEOuM9fHW/msNQBUTnPYUMUQ
hkfWIlEeywyrx6ca3ZsrvcbuY+8RnOP9DBRcpWZ3dHFHKlCfhjjlmVpIMPzA
PTCwZi0f+FctNIrJMAfyabT4YXeX4gOCqEc/Q0kgjnOlH2eMXAdGxfbbDiKj
6BD4Sz2XFjJkJ83gZzW/+Sdmj1kpqwYWhcEIJcIx71ySfR/gUrn9BWjdqjAs
YMA653ruSBAVpiTKjd0cZWh4sWHEU/A9Yz2DzIYy9B5APDTHK5lITyztQARi
vKlNJKzzSlEZykv5zPecwSPpXblwriFnnzjRst84pvkr5Gg/Ezegdj36j4Hk
tag9RJSXlWzHZaUCF1VlnFoKx72MP3YIhYh9PzNHu0WwE9pVcevt1Cz01gMA
tnHD1AeRAY57CHa6sPjucY3kO3rkMW8X7qEV2cRKs5FbhGNiqYCGFWah7Gkk
olJY5J1c2GNWe0RtbXzON9vcytbYMx0psDtgJhhzY2DCJpnYnKuj6LX+mQra
tVepOJCkHbLBh4Sf8ypBeMCon019HNeqnCMW/SuFemgPNHd3kUUfYL/Z9FGA
/mqCx7N4FtCt8zIpx36WL2FC43txZncKM2/iGkcYpruLUEzfdrtBPYIw+BAV
y0xWxET8clI2YYK6FmrVCavShf3h0OlCbnfqCOThumiZRmYEKeitdr/EAqnW
VxB/FWCtcizZgZ/JVo8kaV8ndDRFBfPN5NlwXKzPj1kMOs+Re6ReJx2Dz11d
ipQVXPaUXNp5ygexMYMdqSrVLMBe6K5Xq7DVsmQxB/fgwYu8IhUH2iAuMa7k
nvoTOTWOvimU+CWWQw+Jd6LaHhkd7fzBbFngb7+sYytF9oSb46bH4Z7h+J4X
FsIg3ukBRlsQrfxEvnKvyXN2pi8KGeKaDzH8bUFF4OrBFyNdqInciVtCSxE0
eVFfiog9XHWQRTNB5cCCtJGpUBq63wo/sqyNYL+8G0fZblnprQSzGPks5vN3
TOrO5nnVSLJMfzvumC67HN+ywH+2fx33Fcgwld5NWStOSub4idzTw2vCesGD
00swsd0lKsfnPnH9SxTVN11o5H8TolL3AKonqNZYZYaeoGLZ3ukhdgbBMJMX
chdGGNmHhSCIAdDgfr3mriMDFYEnKBRSeOZSq9xrGFnEBRvfZpDh2LZb+qaI
eAqi2qBOR6uMOS5m5q34Cdirm+Q9SHS0fqhzhqN59UD9Z0f38u/asQreDt7x
wkQFVAZPDPRhaod8WUuluv8iHoaAYFv7h3qee1tJMaEaICVjAhmcjSR1kfIm
I+hyNh4ZS2l55PeMr1ZdgMu1erFaLJ6+8LJ75UlTIapnhceyizl/4ZgmoVCF
UD1HXuowkF99bGNhJex2IK+QE4NK9VNO9YrB0ezEi6sE3GPVLXzy6BZeDayI
k9Qo3xrUmVktK+X/mfiIcZG1sWkA+bNnKFLk9gPBniZOvTe4Xs7DmPJV5UJ8
Un/4wONtpjVk/r5XbJKVxPrE/369cu2EPPd4CYi+1pW31KU4EY0HhR9XHPdW
4ej+eMaKYYtl6dFNVMF/EYDcZO4dJxNyfCwJ9PYLxzVms80YFJO2zAVpWrg7
sin9ZvFKIwCcyUH3iVRsPfssWGEi6HecusILERi7n4ttZPYRQri9pu/hmBP3
iKFVlj353RfJEpi8d6+snBdzkB20xU0IoKfRnklr+d9Y8UwOBg7RWw/c4Aje
5GWlbtTIcdt5b9AC4K4Da5DLCrlis6Ld9/GkxodWtPMGWkqyVcTxBTDopptQ
+RGbs5A4HRwYuZDQl7+HVahIPPjKGTtZwA4ESGGXCsTT6J0Nd0F8hNa1fsjG
NGwXgv6Pl1Q5O48FSXUI/W6lDNYNFnmDpFWXJWLQHib3JB49YzsPYeF/W67J
zW5fJO55EoJVEtRfrZmRZzXBFlDYEtsotZYBNcoE5r0H+gcMfZ4OyjaFFwWM
1bo37BTQo34/dLWYPSS2+kSl/8Pj6+MJAOEM5U0qZ4BLING8Dr2iKMjxjbux
iFyEAk1psEQtIiKlpKCEQSSIgKVEBBOm+Vqt7EojqGsqReDD8iPKLoi5uEmE
X2vQuxAdqVnZYt5YBai/DSnU6ubmLlSQvZD4kfQIuh+6Oh9f/qhQHkKJBh7X
27UwdQ+ervio7qsGCzARuRt5xY39ar992aqoF9PUuDpOrBUD2d4GUb6jePYa
668IPKysfZRQL9ONMVO3hmKHW+7OHaqN45WBeMHZvCtOLOuLFWYjGJiFuOAB
ktG59fkVb/djJee4vafFocXfIv9YUX8oauwkLyNVgJUI3LHhowumJKsWM5f/
rvrroVy/WKoteCSwu9jDV8HSLoyHSpiWFQ39EUX8yT5IBbzV2yluuEqq1ZtB
zzG7tgc2Ceod+RozMx7kAhnsfogbZ5lBH411T55iQT+v0/tbrL7J9/yOdl6u
iTgvMiRFZToIQUCCEfK8oEZ8V6TkWCQLMygCKVwjzp2MDKSkHpPoGTtl8Qfm
2SzjrLrLNFi+HNluRAEAMYWGzw5IAaLV3bfFxadE4VE774z7sud2avJDNWXT
JWEY6t2JTaXgF+l6p/PXWu4mPAgWxrXA/xlE3rE7JHAME8dAjqlEt14VOIu0
yQqXxXay4r5vthQqe7z7+Dl5aLmqjQGQ9JCYGYYBcgE49w0q+86eYjEehNnN
En72sTifxsguXaWVTL2Lt5+ZkC7BvWwRsDfpjWyYkYVu/kLDmVDbKnzLMAb7
jjvDyd3kKgFecYv9GxtkhnT80Eqj5MMyIQwnbUYPapYTJpRswRrBwNnR4i9G
g38P9Nz2l0/+5YfLw3gYu/8na3tXKx9alMwYoOlLzxee7fV1LJ8g261mVmvV
DuxgdfOUDbI1gK0WUo7k5m1GIm2NxAZ13qFSlE3dMYHnZxJF+l56r/BpdYFh
nR9eyuHawhh6dSvlAstr9A+4MWqCxwbexsldATb3nu0n3nv6OKye+/shApgv
zdOEjU3SbrN38x7/cjmO/VHGbA6zmUiXUqFtNbpSGOCBR2Gcovnu0eZScvtV
hduL+O9IUQmGINW6dCb7QUfCoEp4eTtPoF6+3ff9mTxrYqzsQsLMQ/014yL5
ZK1+WX3FDmRhcTEYe/7AqWkrBxFGwRuUM0QjtsmjZJ6Y5WNze8D/g9t3ofW6
NG0xdXY514nKh4GRPgkQgNg6wuQ++5dZZOa9NZMbsmZa2As+dwCts8x8Vmg5
Nrms7sL0ZAaYwhtjbHzJkd/15D5msY/71fvq7buyYdIgQayuJJiet2M9WqoP
WDmxOx8gZRBdrJ1Nf6GcfXW66CfLWocRLdzDCqdnteoH2xX5UJc3xkzP6h+8
PZMrY4pcQxgeBqavlZz456m7v733zv9DBwOuz5B0qBL2xEiqTfwDmjGuBFbq
vB+Soigg4kiyHjdh/M5JMxYaywqdiSdbSNXdFrd8oRoYhicRsu1t9sPhEIDp
KS7JnVXYTJKWhdVLaGMr+rGXPGL8f9XhX0W7OYWyOvF7aqzzIGifSSXZXPAP
f5oyT1exdtjTMq8u77AJbqQglGn7tHHaoHWIwW7RF/X1BoP600LUtiH4UQKB
rAbr/OVq5LVGY9l/fFaKfSQsUCWaoQwBWo9X+gqxAQGJkeK5dipGTbPxEIvY
K5b1iLtvfzsVIPA6mphafJDpc2wrSsQ3qyhtBnlCgLUPPL5EYG5y3bTN8ZE8
zLyOF8zB7+6k/PCqnONhu4yvTvAf3Ox3XoyZjWTTwr+//7CkmPqjS2G/3+Q/
WqNpdkuORbxrBhFyOJiKmMk8C1a+aJ2BRP8Xx9KtbvISS5X0W2HJkS/npGt5
a7y296+gB9Y3oZLr5IzukEmqmLu6wdoSaesgKmZiInpzhrevrZ2YHcv6VPEk
wWrPXpYluBFWu0zclYI8o7whAQIH4XzOid7iZO3rKgR34rrBeFRigERbPZdL
HWONQ8PbvsEkpHVq95sdPWnRd9x/aPu05Kw5sBB62gh0+UIVHtDXwOkzWK2C
nBo+w0MtvNvpun+pgVW2KYg3TsLOo9Mr3WGkq7Rj+tBF6eI2pPmq32/bJj+E
aQrlElXqqWeJ6/EpFfNje+MYqoLaTlOWdg8ZM+gBOlJb6Zu4uV3ZtzDysl+t
jF5uuc6RPMcaA5cFazjVYd7dwLWOk019phPxsQby+jbLr0zK8jAScz5qTusd
kjU9kv3VENutRrzUn4VxvtZxrg81s7II0Q4BqWRCKjM59Plj5g05sKyCV6U9
Ok+KQCBLjYsLLcYcAZbeRuoAu+QevX35szoAh1WvPsBsge1zf8mfGPHadOIz
HPfkXXKMDHLkkm3EBD2ztaxuNnkOsTj3h2nAAK2vIWJzO+ldrVpqkQGBmJ7p
CQLvXpqu3nNGjkUomPDQNH/YYWKPRjoVptBrkpxv6RTYg62AtmOuNokwc1j0
VLO/tsnBpugduPjnsT1WxgNknKediOkSL18hqeJ5HVcp/mlQ6NAs90NfhN53
tAWgktdJa+7n1RMZpR1OS34iuNyv0jfLdpJOszkP9QL3RpKglrI69LHNnVz3
NlRsT6bZPzGWhHIk0LScmdpaaTM2+5RUgsIjOdarKYv3OuOMsZMcET41DWRU
LHR7tDmDrFnNaT7taXnAXsoCToZNGWrk3wK/gWzC3HKxcid3NzEvkXBTmauu
Syx7B+xFy+sTBjooSxZs9l9LwbsL6ORhkR9jU0rGnauNcCyLEfjmFj+sFpT4
LnbEJUK9+GAL03wQbhJe/cKn48mARHleIG1CR55lrNkSSnC30F61H4iWGXRQ
uTJDuQSk76YQKltkwn89A1yOLmEiQoMrigaMpZwIQYAQJUU4jUiKU1KyVT2s
AE9h7Mu848dqwB9FqM8V5LghJAgwx7y8RbsgenZgR0eQjLhuQ46Mt9ruqW9q
cN1l/X/vkEl05gjXzwW4f5i/bwUBnViL5WXtcysgztZcVeOLOdp4f0vRIGAY
PYlPXpr7nUEoefR27RujD1G52mv3vSLEKSvh2CJ8ocCFuRgNVh2FO1sXYRMk
RjCfrq1J43NQkzk5sBs5bDLimMS7PhdrxSoCIrzMB//siCgcXaxeNp4CepI7
/1M9YSGzOyelgM7rgfkeqqAeDUuzEGc0lBG6iIjEDVDYH7eFhGeADT4psjWI
GM/bynHLtmKettTykI+Cm1GvpgATKw7+0F/us2bwOxNQNB0684a2SDqVxUx7
to6I4G2V0OmAGF1Ymze/D2qaWtcv+Hen7155j8FDvizDeksDaBZcy98mZb2H
VlmS7W9Z61dEdbXnuir21iU2CNBLMd594O9i3E7UmsfMxTsatA4KVZdKVywm
yfcRSWbBmg3V1rGHAm7Gf+T7OlzvucOCjPj3QF2x6J+8CUgMvZa35taEVfNd
qGSoO7uqvrGXrSH2pk15Zgt7eM5jbmhCU4ROEn8VfpJcH2NLEH5yInTONWqN
Phn2c/z/05CDS2LQoZNPUf2Ou2jaFaokbA4hZUqNFyj6p9zZtNHfP2o+FpZ/
vUdMNOC5CJVD6bZxrweDEY4w5Y+vDKU0eT+0ha7JPIJs/7CiHY1kYhHMCGuG
WVcL3Whv/gaN3lKvLgDe8SMIdHjJfd8dQ1prKaHGs1a4VzQVc9nBhRsg0PNP
iApvUDbSrEebpNlo0aJdw8kOvpq6br1cgADQwU51PbuBJ0fPkQ5H9e3+u7Sp
mREUxuU9anaLaoRMP4Mv8mGkOi43cx8MmbnWHBGGZ7GsQvGKgf/KOm4b116h
I+N0s6Ix3psGppNe/eBvRsk0Yg2XmRydGqQoLhZeiMU01hitFNUJsSpWyDkJ
EytSeMIA4/39JH2tvP+FXuTHvMwu3d1zht98kLBPjnBF5OR2ohuxg0FnEJVP
M2Ac9s72nzv/eYR3oj7oFGcOkNt8O2ApkORBnTG0aYTZ9BZnOZMhCtkoprbJ
vbeR1lLrkwn0SZtEKw6eAnqUkwApb9Lhf8eZiEBvBykfX11E1aqhDZVclCQS
plE7O0EDd0mUveRb02C7+RsuginiuB1pYiV4j6ZIvB5ys6Nvj3HYEI86tSZF
SB8Vv2l0Q35dMBb8NtAdOEuLXjY2CrNENebBHDZq8z4b7m7Q8MKiBIBnTWfq
bT09eMc4KQ8PbKd8EanlofnWpjms5lWAGSavQvSlcBNoJysXVjVwijFy5ewr
9s8uup7npLfi51O0l1jvDj0jPPVDUkt1GYOiQn1a8+uLy2JSUclWEKhJ/4DL
mpRXHJMWahlQOpucWonVudpXTlrQ2qofVF8YdcWTtXykrHAWYxV7nNoa9zXI
fZRxLXSgzWFPV2+uITlixDFZPRROOOTOWRJsZOdezPrBjXFuO/4w7TuKqVaR
T/U2rST3qKYU9Bka/p3r3/dndA/mkuupMAhAL7To/nMKAH0HqTlEWgh5OGL8
GtOzsxelwIBpFtX3tObP6csHWR6WT9+Few7o7FtpyS7fXNU1YnL0hksCQjby
frv5TTII/2zEKFwpKvSzqloHw6POz1T3Q//V8nWVtH7qSgAgQJyL54HEZwvs
SvZtxdrhuyFMiz6GTLznMUgFt+sRwhYnR6eMRZLxRbBzUxO9e3YYi3Z4JqJv
Fdmw2Z+Dcd5SK6ekD7WKGIvRQwV3wU5GjDlzuYoXKhNKosJDHV/MYXKj2bb8
62ZFSCMd79DefSfvIefkKCxhNxV/zotgQKOeq64qXpfV1SczRRP2R6hL0ROV
WkNkI6OtgYGSdq39kOPX2SIm9bdsB3JytHRaPjRkZamDISGffntnLhJNd65z
GaTH/JQHvTPiMKCInMsBlh3cYQOclIKX29LkzrBOdarkCfXfnYeeRosFa35D
QHcOGcRrzr6SVhSobTk/KsgErTtS9a31roi3Bj7PDd5ahXGLB7ubHFnGs2fJ
UfY0anhSE9BpTWBbOnz1zDGyAKycOsxFNFjmeqJWYXBX0fi4IhyFLQgfoU9I
HsNHHdWMGQ0Nl/xgV1+UUEc4B+7BXXX6LKuhfIFpgOgXXRFuf2lMygITjiVy
TvmW5Iyav/XUf9/bLI6ZfVSMIF7qwUzI/IeQ9kY+tnwR/fMFranIzLhtDDns
Gf0VHWanRvKqiYm+8RLOEh8Qgf3Y2jlkxNve1q/PslJqNCHiHWs580LTNIta
0AUB+Ky/x0h8pAwtfP6yw2fxR8Yy+xWFeppRDvrsj/PI5X194Xzk6VPgXxQX
1WI/RR5NFz9i5HG5BKH5uDFlD/QosrKMq7ej3fd2xs98WUYp0ZRuX+KbnNk6
ERboYbqUAUTpPtTzB0CSU8BCtf7P6ijhhEh9Y+KKKDN8fULbvHF1uzbuDfBj
30ZEPHK9aDbjXawefT1hcLN1vo07gaQuWvx6NMt1AmtNX2JwHVSYsRwK+zkv
AYx5C9ljYA2vpFeIgv5bvQdh4pMCl1mAPThlKUBRZLhcyx7/CHq82Z8BqoMO
06Y4/i1gR22Y3IkjRqBktD+oXKPw0FnakW6M/GB5/hoMO0IzoMN//30qnQkG
hI2RQ4SprO6QM2AvCYZHSzOqFZG4cZEfieR3id2ZLxklnhXbdO+1BUsMp8y1
VCuZk11mXvhm3urzFEwH4NGWAlF0qINM2gdU54ku0W9xXbe1Xg6TsUPxkV7p
k7lJx1nEElq8o8BfTj0u1exnThVHt2gKYTLC206buT/5UIfASihZoTMpYmDV
l1ohSuXA+HWcRANB1OuegzgBA1BvmaZOpqhSZtIkmNvv7iNhaKLZNq0jZCnZ
AAprCHij63atzzPL1/N4py1KAjkr1Vl8YXCZlMv9oufQW2IWxAyIYdEhMEa0
oWQ0Rcc483JqCjuZEhv3WKpjKEFoH2AI1qG7UWvkCYC5M6mGpUwgcqf8ju0N
VG4bU1mvLJqYAZnMvuzZUUREKIfjJb8HhiQhEuPN1Ca2PuKDQNliM31QTmrZ
iQMsJdtVBSmTzmR9Uci+4xIO0KaNti8X2uJKhEDjFPRfNIIL7M27AUgKUtdV
d2MgG4nRHL64W89YJaqAhItzcEOZmRrCBS7jB+XoA86t/BtoMCajGgxKw5+M
ss6jjRC1ECgbeHmpK23JmYVt/A6O/7zKL1WEaYV3BOPn6V3Z/SeU/qjPO73y
LyzNVe7v+G/7yXdxzm8Jpn8e+ZI1t4cwcLNr8QVsqZCVu6ch1a0MDZpBDBeH
tQYGTKaJRL3JdY2vaudKgdp42GX2uyEM0bqK8vAlezcm+wGlz0aF0BcYdaFF
xHgVAJZQwxraW/DEEP7QSxi2MTMIUc/b6ZXccC2yHtZHGjLxcAPZ3qb6LNVP
XZYFGr0riNZUYL93tnN/4QC2QxcRnj2sWBENZ2mIBrGoRRN7FJacnmEUK5RE
R2RtujIlJ3Jzv4XtFAyUXTpgjdLSnZgEcqLSTeGFfewTLkI5e/pU/PbDUpPu
0MFdmGyK6jdvuXwEBPn8izizsxauGo5tvA5nTIYI9599QvgL61B/NwqM32pa
EsxJ++3Z3kS407Jw7/ydtGd4k5yuvGGEXG0FdYlxuVTYuyDsit2EQjBp9zHn
wKTR0VoP683/r/0aOQTy+f85a2fOMD30prPolIFpH4Iz3PQsl1y3RfRzlzGY
zXRgBhPXI54o6aGtAKCuCGesnsKsu6pd0fTEMynOxHX4jJ0Vw1eufwpw2ZV5
Ri94WtvZyrqSCoboc1Rrvx8w7ZYmr4npU0xuNLncAOHJJRSLV6XZ5ThB9FRX
UW4AJx9CMQfGd0SRn3HS83MVqyV/5G+2BaOkos6E9L35MzWqb5+bwsdm7F8t
7MWBD7MC4pfTvo/1XGM3ZZaskCPdE6SzN+lfQbm5fsoyQ/mmR2RR4ccNcQeM
8AaYRmApYhQYVcOq60P9HZs7fBmq3avedAF4Y3OvXYS6NCRTgPv0AlueFYVi
B7+3psJ6+LhMy1sPSpsvuS71BA6nXBKx3BBTBgPwzeJSMl5FUstD7T+aBw0D
l4fsN2GxQIFPevQWaif9OdtF2gYIQvtf3+HeMdmduQ/EXLSi7/vvSbK6FPJ8
bZFGB53Efr3e/RwYcBJQ8uHj8u3IMy4twfGBX6nwwW59aV9oc5EJ8zv2hbgL
7X8fr0tAgorYp2sWQ20NYwe7cQR/31PDbwGJXAlnWdoL+0eImVmeJQarbMa1
WM2TXO8OHalN9R+bgwpKDNNsg1BTBhO4nmNkPXLjcUTwMpOaJhWqt95bsQpR
c1X3VkfoEohG85sDxyPQpfxtZlQLzrjt7jeiOf21x71t3xrqEstu7fpP/jyk
mxXSAqjVknMJ6yp8Hey9o51H8qmY6fJtmjjOlAd/Rav32Rw6pxh2r3i+bYen
bhaCf1UMSHNItUR5PQwnZ0RPCOnvGBHGoPvoDionfOwoCoXw7NiMRXimQAX0
yIbOUE8iUv5EGqDMTMi8stkK6Rfj9ZEDptzpJlpmJLC/yeorNa4V+SaUX+ZO
Rrc5kF31/z8weBVc/hG+4tLwkakI5GHzF28dRsVDpf32ryWyhw0uV+HFSbqU
2PGaZDtnsbzqoszVJf0cGBPr7m8JzyyoSf7+iFshjr/lqeBwI8UHN063FRma
z5/QfaTVRT3OOenm5gpn8A3+XRcNFnhZiI54bA+XsmnQ6E0cTtlK76i2rgWr
vbrvGTluGYiNkXL/b+P5W2zDrAcIbmSVlK4CJ5P/zeXnTHKm7Vsdwk7oiY2f
KlJ/2spicT1tJSmXyZUkJ0qZ2gRB62Poy5vXY9rwG3Lnv67HK+oKJ745Qv7O
A0Vx3xO4JtBEx98eeAmrEmAPXfaoaL9Q4Mrr5lx5kwbyltEMyp1M/s1abtrf
RJmdsFWmdCIGF4B79pT05K4pVKUPe5+3w6Yv0/F4sZtRAJILqFd4bzqyVs0Z
0GWCtNjztyHIS4YrJbzVQZSkrzQOTlLi+FTaYhelG4SpIjIWdU9/OlIlMMyX
V2qRcOKO+o3N/RC3tMCEwa+an34G+yh+t9NQScQv85UlX/93LE8toXBuGhHu
dMttTKXprQS5m3iMJYKTK+OYtBcSUIEGC2sBrYYvoAtzxXoeznU+6L1sFaAa
KXGMWbn0Yf9w3UoLhwCVNG8bW/FbhYZxnNTvR10eaxEFJAK9NsehQ+GjtEQ0
TLefGXSn3VSsBYeIIAfRV7dHpdVVwsI6bxG0tYLjULPlkZDZndt7zmHjBODy
f/uGLMgcn3q7wmbGnA812X5nyif8hjLTILHpvwEpK7mOYLzNV/PrTAZBoYSM
j4jdu16n4ItwD8VAC0jeQ/Ek/lPCacFE3Dmvhgpi+On/Z600NhrpAT2y9mP2
Od0vmtb3VnwVVTI5JhLTVdnntSZabC6gtfbdqVnPQBFsZvxLZDl/WQEhdNvK
Fmx2ig3JNzqm7iJm3z2pn0hfOBTZSqb391a8kUeVtrG8aCterW8B13isqGRv
rvKyHdaxdgIJwwP7/qDf+2pwWitsbIDmx5Rn0HMVEHno2ja880Rn+vqMpKR5
FtRRSnbPguMR7m+egCxLOSG7n9DxQ5T45s5ULWD+aYuHaTSFEbQUey5fkT6U
IhM6hbmAIzSYKz/DH7cKD9Q/FKEQkd9HC1mrrzJWdAP2LTkIc2Y2NzGti3E4
Y9hRZbMPBAZl1V5aaT1XjSxl2Ei+V5njmTXps4Qr3YGoLPeJ7Li2rCU4/qaA
ck/NoTdMMuSiEXQukQ13uwLp6+Et56aNZYSPzpVeTTKfd0SY+Ig7cai3qLAD
8lkvI6pJ0x/q4orUMRMn0U33ptYD4Ap4CABLjyz+woc+xn8vfiOR0gU/XpTg
wnfiHUW8Eec+2+uXTF+Gx8eDt3PLsm8/sVZ0XBcrYVwZBG6DIiX97u9nXx1f
CpRYoZfbFtQrAHuo+7z9znarzGVMdY7pcRJmsCOLeuXJb+eEnzDeZhr8h1wP
TtMYhVNUv0KTQRywHQRRlazgtIPOJjhGorHqs3M9lZeZYjIMKXxFA/84ouiV
7NfUNS+QWSnDMDuJ+WjttI/Hkgar8WEdG0aGMnrEPJtaK4lmWP1qDaNOt2XD
+rh45lBU/hR5g6QoUjEtViOs2MHNrAsxKRA+dNOgI5bSk71xS6CWmVF4MOzU
aGdPqcdZCh2YFHZvvXzOhGx0s9v4qLxrh83EhYIQb0K1zTezl+yhCQdHSKVJ
10qNc9XIYKTuBEXuKUnN+AL7u5Ub3EJpgc2JZBchbmNNQV3iOMGYSfwTNoF4
SNq5TwTN/m8jy+NU+41SwoNUfIWbNHWBMqUIXu5xe4JIry3cKEkWv261olNm
RtQTNyNd9pxrQDuT6I40LkPIF4uOFnd99UA9NuPJ5kcR7vppHhVCDi3U9jGR
Hy5DMVo77oV4ReDmUyPJgRLAo9rwyGhdX4KkvHoyjP15+XoTAngvY6dWMTKO
o7NMT2fRAdPtBDt0FudLLCtf3IhQCnkkV3Eznlr/papSgPfQzN/iv9kg+V5B
ka3wl5eFfX0MQSQvE4ZX1zQSzIOMGlpfph+Yzgp5fThYc0BZX4xCqrsSjVbV
fx7qlRAbfZ3LaEJzmvNhuXjDFPcAZQgL0LJN/++TikuH0T+cSaT0hxp+gK2u
gX1p3ugziCwylN/yypSld2psOrp7EW9wIdA14eLdH7x2mz2ZS1ik3ZKUbq1n
SJHAAzY7Bsp6HIcIEnZtX75/vBryYBJsZ7z/2621PXDGpHlVAbK9jfjNfJXV
US4lb56KdLQa+icAMH7ZcnOx965s/iGJG17pQrmnSYy26SvzN5CMGXvPTMSB
/0pA2sE2WV5elo5yIPFXE1m9uJvrGD7z2dMwQTP0xt39fz7bnOc9VyvO1I4K
WJO+K2JCSi/dKeNo48BJ299M8OyyrrtTt6vdZvPrCD98nM/31SJQlyJhX8BO
aoOtbRCWclhoMQvSV31VUX67Vo19ChrWPMVGZHQbjpdKppjdhzB9j+2mkwQ4
Z+flEEi0NtoBazH/d9o8Qe4TkD+CFwIYUNt6abwHRCcMRELKx+aVgDpkdsHZ
tF3mox05BrEaZSb2txeBeO9rZXDPiMtfyRPphdizCR35uRggzT+jb/yjdJzp
7pfu080JbGWo+pk2ZSPKIQ+E0eIQiAzWYoVWN9y+r+QQ6KSvCCeYDEDPQwaN
GdCQLPkcM68z/lZfykk8CR7+U1RvY5msUtukN0AinSWF8X5LI3UjMMfKqlpG
3443AmT4j4q+cnwNtYuCz1z0F8hKUJcSMnqcCKEJsFTYzME9tskw3WGFXGB7
yXm9HOfNm0nq7BxtDbI58/sp7h+vVcZDKy0Imn37O4h0PhIAlRPj3cw1lq1B
/wNrEewbqOfkI8xgfiZTZvfSo/gqUhbF+QAJjp81Xcr6/eSbXOdkIPWkiQ88
qSiefc7UM9mATSLkh34ryvp1FLEyaTfc7SJ+gVjSAhgmeBZVQP50CFC/mFid
yMPdU6oZHc+Bs8rkFtFNj3aUwQuhgS7JyMW6tFY+XaZbGH/BALB6RZNBg+fQ
paPQMC7eZ04ERvsZfdRA84sD4vYUrSBjnALoICFK2GPaSzDC1Xrdq2shFBc3
xm6fvLn7b+zke34zNFwCBb55M6U1XXLUepzXpb5W5VhWnPNuw09+RUbTRmkp
6YEcVHUduZPs9VHJ0SGJ42nXsclCKnvNafPB2tvJs+zTqnFN3FXOFrhGnTcj
32d9SF3mpYbvR6t5ygHyByu3cyKwGKxPnELuaojUUm8Tk7xBuch3DsD8lhRb
8d7+0nprY/RG6u85zmNLUq9o+neXAvdOP/jT0qviZD2o8EmpswkIfjkCptmI
VMhgBOyfb01t8J0Zy1YI15xdexnl6DSKVTNY3bmjSap3O4dQmEvgZAu+z/NN
cES1WrGHYXCNxTdHgGeLNN0qyGyaNN4Hz9mfbCUv3zL+7lS/Jg3L/hVUkEjt
LA4l0TOub5pVYwrUtoj8gbMp2DcjiGuyfKJcl5sf41sk3SCvUDaCdzgcDn97
RkopfD/zZ0wnYOyFT9sCTLqyN//5mincK6+t315yjZEejQ8T7aU7Hxmkz08d
WDHiK8Fubx+MGWPSww+vNOSiFNs/tGPMTLdY8Tnfxoqt2NQUH0sWuvLuaEi1
hgSGeKluX9Vb1MtGmWkKv/z2xQmQStjuuqeXQexibKLcLEie07PhQhZ2Fa6G
BJzmcCJigw3b55O6K5DJlAXqqQehssjSbrYuzq5NOp1GiA4+wq+EXLoBZnMy
vfh3tMN27mQufgkAn5i7oWMYGeT2wStaJ/VX7oouoeHHmUMJ3Dfthskaa4cC
qd08DUM9CYUO7KWcYCpC3paQHZjWF3AMH17hOn61LqnfcuG8nuhdKxkzBxTM
aYOP5wUpLUsASYyOCGoj8gypdzJf+kSTrBY+fnDHGTSz+Rc8vOtrxDMu+Tin
0oSMA1coix6gXz9FEfT4uBVnVI558j9kBVJKaP/rDyPBbAfDVv0a4lGGdovO
os/7h8fZGSGva6evos2HWRt7JkfrN28OR79gn8ky+PUCiV7RX0MOvirP+wCN
wkdVzfc/pI2zs+2rZz/b8lbQSBU5neRRkbdvTZ41R/7FrIcfMf0wZaOpzlpV
/Zo80r/46I1FKdrxEGgRW5zdBTieYRDpMfwyWgzAvcFUd1HVdoKclNAikVgx
YW6opbSm4Rr/yj3WFS5bLwUc35hgjRsL0o4ikQLgMzb1uBA86ynQu41rLgXW
VxVPb97qmjz4qqSSySz6otW161Q8OGtB4hX8r756lZSFbXWf9u9zePM27fSt
z09vjiayqgpG/DNzbaTXnC2kGFTnmp5z/Vd11z0t2Rt4KLGEADfCGD0XasKi
iVKAMJycmRwnbwiACbRvJn7bUr3y2KPDQn/l+upoTPkAv4ULlFaiBZ7GZMo2
nF3JH3nPZfcZLvo8LUaoZkRXcU5bpj6pF2TnII5eWVeYWWSIBh4RXVCi5c8O
lQLy9cj0A7T6YJeSYjjszp9XwEPzSdALYlsYqcHIPUGn7X2ryV78IFflCYQk
WSbpod6zdYOv3JOKLq2TGKLOYsFWFYzokPMcZ4mjwmhcjhpQ2O0G2i+ZEvzC
kSzaubLMsK6SS+i2ZhyHt4qqzUCvcAdIK9utXVwEDuM3BDg8dmlC8Ny84Eys
frmb1M5awLUIxPCoZep1XsDsHEuej9PMnBK3JlJN3kKvx5E7cIppy7leYNs8
IQUQQVqoH1dBeEuvzNhwa+s2jLxA912dMf07/9a7m1iCG6L5P1yyyIHn7qrC
h9T8YmNtEOljt0uhe7nshUaJhvljfOC02wjHpfrlIBjAScBhOEfzJDenkCV3
zqRWPZflU8DNi3TN2mo84w8EyGbg92h86RLvTwmHeqLjSdUNYydR6x/fV3ep
vLE7b5FRHZQNHpoYDOOKI340O8wmq8GDmYvOYKrC0s8og7B5tyaiCKMAUR1Y
XDlhLRI37xqalDk8kl8t0g3yPooc4ncDSH360lVePoRzOI8qpEpgq3WiPaIu
p6Zh8fzYx8Qb9NpmDVbTOnZ1lP8puHJdFfefw6eurvdMn36lJ291GQ8YvTDJ
OsuJF0ySJ9WCCy2gWyMClB2gJS1KkHLtBUSAUr3+mdU6BsamJ49hBKKKtK3X
JOydjJwgFqL2y1SeP6TowR8bJVj5lPxwUIil4ZF8erZMYwahrxvICXZHPRgd
KimBBDc6tzMJ44TBtmnNCFlauIi+z2AtMtafY56ar4Qc1gN3T77YHADDWvIi
8OvCunm44tKsernRr9OG6GiMpmD/rcs4vPILmcIONeqPkrHbmdFMNUgGFbEw
xmsVOLzMWo2m/OpAkhKgj0Kd4lYv0hLdqvmGhQCB9nJ2OzsPD9BxjwwI5g72
zNGLzca9YTgHGDrTrqcuYXguMjMFroktIovBfFqBo7xzZvrpxS5etPA/pwNr
3WmMmW35sFNojqbzytt0BMeAbKoM5N09mRjhNOASqTtCa2ZuLPqpYtwkxnSb
jEqqHgCERUhn5IDyeTdfVjejD259gv0Mp4d2kixOeYGmK76cgvUrfNGoVA1b
IXko+Dh8phpWFy4dJ5Q3LTgV/SvDDkYTGVzDB/HFpgsDScHb7aXMhTZYZ8iM
QG/XzPlGpSsL90iyqaJrjW+PCNxm914st3oxmaBWRh58j+kqqulazlcS/Lcz
dD1wPNPSkos71p5y4sY+fVhjNfm8umQ6E8hRRopfsqG3bLitzRXAUtX95vCl
tUtrPDJRaywgj/KdfVAhDWg14YeKlEpvaPW+3alHQ4wEE3A7JTPuAlTPBP1+
6sCbauAjaAUoSOW3hp6C9qn4AdOci7oS0oaX2C1gVFRMF49ZJWbFa3JP2HiN
Wf8sIr492VjF5brmafdjVExsafRzaULqdBqyxYQ1fUDLDS93VhFU/EKQsS26
gGGq+Hart9r+qpjzoOF4F3zZBnqejQ5VMjSMFMaQc4V7/1tg/7ZBKqADcwZy
HWiWk3f67Wy26mHxdavI8Nf7VroNvVoVQLnu2Simj1LUVQa72PWKgZYh7ynA
Mc+bPDFZgtAs0bSGYjP2hK4OIx2DgoWaIFRs1WfMrDEH2v7xxOBjX0Zxx1kf
bc75nug6+hlqSirsw4husquxRDIOmYlIsX5hg4SYaXll6EomM7jRRyt8TzWv
eg9/CDpCb8Q4EryD5OjmWqWQL+vP4rmAuNbkvbw+TAs8k0fscPlMf0IltRd3
k2O8B8m+Mw3DdDDmg+cPuX8Ynt4ngkdiDhM2PAMMzE+xnQmHFhXJHuaonPQq
AJqD5m1PPqnaUjaX0X5zSIQYH/M+BwbAwGeBP1pWlTyYpeslzg8lCmkBgaIE
h7g7z48jnh6YyGJ0zK4iXGT52JtuZd4+VDWpjnAdLpaTAp6IjJyTNvlioLlK
gyUY0Cj7eq7lws323WG7kiK4JhF+Lyy52+gMW56oO8yDxiet5kxfLz5yV1+2
+1DoYJUP3gz3CtKmJ1qiz2nDYz/TIXd2b5A3vNaeqvVCFOYyMuUqw29tlwU+
LpR3ietxIwC8BDo9D17pWgrYUmLOM9q85GlNBtXlfBDVDYBKzWbujjteSeaf
I0vo36PJdW0yF3ALZDh3fk6OTsW2o6/UlGtedkCFRa017q16C9h/4yBs0t01
hKH042nfy+hGmaCoTIE15ApFD9zE0wOZgROzXvizoSlkEfMYyiGp2rO9Tl5g
7drf5PF9/Pgax5sPaG92ltL2LqQCefHJMsuCalKwcOrx/kocQAUJyDsJAU2k
sC6WBW6bS47o22T3XkqoGfl0FhXTm9PwpR4hU/gvwEWrg8cpcU4/S6Jf095M
/ix7Ox+mrI9SA5TBxhsMWKuWh1bPmJb4E1+PnbHeemZ5I3GF0Uz+SnKoqcRZ
wcetlaJcf3DW1YA6HExlmgS+KTm8boKqcC030LPw0RxuqPAd0DyY/KQotJl2
X9Ud6ZLH72kwvn8T+UxxpBwhobYrD6lCvF6QT7n9czfN1HSePh0yf51ZOso0
FI1bVBDAnVTWVFDfOyyKubXm6EZz9BBnPyu+HhtEszhQ4G94qFRLiycGlgWK
EtLdvcAzErvT/om/n5b50rzzu2N4PsgCzo96quK3DHeBnCbS8N0iTfoULu8U
TyAVt1zEl5Kz/zQsuAO7Y5L57zCsjcf5cDFSCIPsEk+WZWkdyYGJ0wmSr3AO
swOa7QfBlnblivm+bN1D6YbhtFFm6xpPcE2mQweEE9PWvhY1ykMjlqZIrzz/
Xl8gU4F3I5dUIOHww3y73wfbjeFvPpnAMvTTqZ+VJdUIXu6t16qmo9yE+uw0
w0CmPAD4WZ5qEhlxoGQnTpoiQB1Xp8kBf6w1k8V9qhXoQPvdF8IicvYArP6f
KY0ATQSJCcetuBSzhamK6s9M7T6T82NctJwo3vspPokZdhD0uyVfP8V0ROaJ
ZQbSX3Vg181qUN6hYxSZ7gDk0zN7RscylbsE9kJwyDvijR9/j6zkPz3PNKUn
jCBtt0rSeZSPN4y/4fTJfmLwmeJFCyu6/FUBOvgLDhqKv0PwDB+oRx/avvwj
VEyvAqMHAPip3gF9oEoaWgEiKLabAsSOT8kbltL2s11eRE1aZBMwaomIiXJH
Fy/KvT8Hh97INm13QEffjiGd5SN1J+flFyTJbLLmxDjeFb8+s5skZRMqPBdI
IXh4+d/JGJR5HlhUCgJK4TpHfwHhTQMJUc0fuEnEsCPln3+sd7uLcpW5K8Jm
hnTylbfiqQZtRGZ+8mltYTa6SAk7kfG+lokr2VCOnqPP4DMZa3Uj0ITeCi2h
La7OgDH352jN59vkUMaNlyDpMPdg+rF0RZ8nq+tFrhLU5R2gMfP0OTT8/P39
xWQH+2xiEd2p3j+v7r8fu1g+b7ZXRmxDH+7C+oC2WLdLfl7dv0ScyY5fd7uG
h8xyo84pTxaPACdmgVQGjSf9hq9HVvbqJhVYkfiA8adCujcinHq9bQq1/9aR
g3mbCPaqqCeeOiEVRxH4YpL/iOa91W/fKuGq/ullRhHWNK+yL+sZs5QC3Xvf
o7YCk/uUByTnnjskLglv79JJ0PsJXvLDb38Vx7ys7lHSgCfOcMHVVO5VTzHY
nUYvuwWoRnsEKd3Oh2isith3ypN74OWc0aE0QSqXz3dMpKGdBZGqDv9SV8le
IrCkn/fsFD9NF77jH1eDQeMuG3FzsX1pYyNWeXmgmkckdrLvczsFz6nHeUz0
FoYGpXLHbHGEWhrgFv9HiVicCgjem9bpijYoAdbkpdx8jDItdLCyHhRXn9Ju
OsklOqhtkX4MCGq6nbzAAl1G8Fgvi1x92ftKaK86J8LqEt4NdZ2T9tWjbkif
ilVnaC37j91qXIEEEfbUi9oYJW31+O9hUswsD6+2k8Wd79EUuDKO4VCIWn2h
c7I3q/L9/oSdiojL8XS+dbEUgWO+W2yzHKhOw47mFjrkwOgyMu+eXMH+h/74
/KoKqm4d+Zd4qo6yk4NAZKwY/Bq+x+sxJgHYmNK2X3T6RNEJVL7u6XTGWMIG
iEEah0iwZaTXJfo86Dbit2jBMcuDnZ0o5ddRYLm/4PCuh/xMirGI7SOZxn/f
m7N58SJOTBKuCkaF8wdX/MLgPMzah9jTBBEQ4tiE+olKKUU/NzF+IJr88b8A
FsIyZoIhEYz2SSJsk1CW2+btyMEcjB07Nqr3je6gTXIxl6CQxi52KPnx6vgl
+fwl1DeKlgNu+9Bn2pgs4qLOYEtXTF9ch3MSg4tgAl+kfrFGNvwry92z1UJD
dHcEhi+w0Epry8+Oz4YTlgNDeAelxZEtV1l3cura9g382i/RZsdxd2SPhi0Z
1atDb9nxZ8x27aegUVmBswq8x+ysfqfoIIc9z/9lZ/cF/QP6rsoerXkhZ1nT
E/bJX2g1Fookks/raK4aWMMIp/4Pek64fnxVMr5Yb6e2fO9+p+9L3nNJdAuQ
x2dbIn5tIujEjRsSBH95Q8W/Twlg1hk5BNQPRucAJaPppFIBQJly+dq5xDws
bPRZ9ZEokDL8JZUAhnQ5Ook2FcYIKxt7jaNAW8/U0AUGf0fzyIR5aaUvZS+f
unYdkdOu5yKDciBe6xV5TeOoFYfFi6kd0RZCmsAIrtdec7XuyOQyCbedO86Q
a5tdjXqiqFQKlOTvYZxF8hcRpPXotqUH0yGIxRSuTdiNvh6UXtv1q81IE0tY
EicmbnmhvApUUfe7hgZvDRXsU8JAPWAPl1c2JjHmlZaiIgFH52E0My4Makm4
xRLY4k53OALwwxPBf5Mh02Xza5AV/YgDoRplu/foVfzeJyAYaHg1wjKPafnl
znuHkZbymvvGQk/XDbJ6pQTLsSk4UecDxOCTsfX4tfQG0KRUk/66LlOLYSYO
YZ5IeA3Pdskx47l58wpQp9ZWgn1vOOTJBSzsVQ132Oxf02h3P0J7S1G8koCW
BcduSA71srcyge7qp2BqG3WDBwyV+oPD9qW8KzxU2Anl53XXEbLsP9kAzYW6
nbsMa9W1d5+5PahPuxuUGsltjOOoLNuXHPHJu1YpMbacbytip3aq9WxG2jSj
CnqsIBIkHZqQMElAkbemLU/fyHWJdhT6E+l9fpVjcdEoSFLTxHnu5Tuk/qIx
qnYxMyCMrEBy0/dWHcieM79kqyVLc3kz2ZYWIJnbJkSg371DhnQtUVJtb5Bi
rwRiPHZVJfzK7hdo44CMUR/WIjAJodZ7RYL10dfhTSxLBGWGO9MEmQ228CPt
7BqXI6t6IIEMZwBPEG0GEeD2oUTifytjhwt6qglTMmZvXgvz4hveyRfQdasI
CTpH4ujCkBpnvNTOZZlEk3l4sSg1QqmI8JQIyJ/xBm5PtX6CWL3SI2gzh9E4
H3/6JP/4tJv6BlzsH8x1CtYLw6zf0weTAn0GMlK9nw1Wi88R3eXwTIfwNvO7
06vU4x8++wE+I4KE8REiRR1hzhUtkAnnr5tbavDAKZeVO367cd5mQA/YA+H3
POoJKQDr59RheXtTBn8XRd9kICYMIOTAINuDfVYgHuAfhbAyt4+Fa7YWjCEc
Ze68XlsqsRXlzO3GpCUlOGzFoybEksLHAykZ5fksmj1CiV66Qn+2mc7BRby/
0hdRy0qqE1wCyFdZJJkAA57df4M9JWm+F0I7fIOux74Ks/TwArnd4i8YZTMG
hhVCYDmzv6jdrjKsvdvLa0zuAbZDSbe2y1GVu2CGYtS+isqSQF8Of7IRJIyl
SXg/+XpER56XvyIKLhSikQjw8KHcXKDTYxW2KAL/0L02KMcwsW6e0c1/zSdG
SMYtI09JVCWxB3Sx6SB46SCdy98awfgcX1HWtzcvD5ycKzhUrvxloWHuaUx1
+FBiGaGqQ8/E/qjtUXQk7b9cwyt3i0QXXHR6DG/4mnbtWSwJE6aOlWYTHvS1
3N1f5pA42FM3cwx/ZQ3zFpr9FJuHpBtIEQOrwqne3frtdQAE0Hj+CAEt8jDb
jmDxJM4/p7OSg/893UAjL4YHTWiGP7dNSJhkHb9hV0l0RAAU8zFOmD8oetXk
zJjoVj/EvQ+M5VG76CvXBF4r6k72ea7EnMVP4XgtV2ydMNtt8NhqT3PUz1JP
5sdv0Ky7wLAM1W8P98AOECUrmq+3Hvj6VwcLFq4Av6bwqj919rRzHli++RkQ
g9gSPowE/SVihbs9L0yIG097Jde6JECYKCC0EHs5wAFwEx2c1YN4YWCjWwUP
LHTjtApaCq5NwLN7Jr0U8ID8zALtt48yUS1B0YE+rVmlzvEg3/jm1F+fdxDL
IVDgIdcU5E1SviqjFNqqt331ieZLutRZgZok5TA3PUyAP2A5ybXUsXNvZH0g
qgql177dAW+amann07N5JuSWdIrk31kgpvqX4HzP4dNmKR87U5pTsNlOyVPU
NPykzwCugKFU9WYKp9IyEM8zPVzoByXWrBuJx13MXPtMs0mPrCdAiqEJJdom
YDMYv3UV89OKiK/zTnDdcP8L9jVBVev8nqq2hRamStHmwyyu9en9a9D6NLBe
MlWnwmW5oi2tO1vHIfRNLZyDzHh/EK0OT5AqP7kDDrENciDAIEBxTQFunGib
dwzNtl0EJ8yOnjLKpu1p4a8gbzyT9M68MHCR9dX0T7DGTicLTVRqGjLwLoNA
CdQIEvkVy8aBdGoiIfmlXjbs0MNgKjJDeJjbHvDmxo4SUrYF0ac6pBhfsCjg
f8/WJkdArsQuay+PVfFJYB2QnVGnnqZDzgS5cLoWytcIVnIVbMFCB55Db90p
Y1YyIi4XZqbQOp+33smciTq9rwHrGvYlvhfVW6Jr2/CtWtAmQlLr0RRRcJv2
xNahS4+mY6KihzEWBh5sC+XNd6QpW7S2HE1HHksSoKq9qfcxrjC6AOpDS0VY
PBrWonkfLRZ3vCrRDhYALO37XrvrFt9y+f1vH7QuwBwXkcxoVpWwTV5kloQ3
BmKLE7qNMxtRUWfxfSzHR6n8SQPzTdmdZAvpZ2gYsNWoUvdsbZhd2TVhop5e
DMi7px1ziV/IqZdSJ8xi4YJ7xUReLKqGCmhzChUKvJlgwmnOCFdlk4Kr1BXJ
MUL6XZVMGm49zG8O1uTIP8BWgXHiigGIddftQLFAWfnROREjrAXLelLaSFbN
hZXmgoRUaFYAvYQ+s6KpeoOZ9g7L9bIShF/C8GVw68ABPtYTNcLy7R8wXUtl
gmMJzKezRyHZlY/uqafBbqXBSnfulzvA8yqKAg8+kz9qZC419wLeSzQSkBmB
64C8qWyzTpmpaAEKId9LTFfNZs57GvJ01aDE4L/wYFXaRwlQdjZCdmhwELtZ
fLY+nGYuCuNpu1MWIwwoBW0RCjnLH4cNCINWTV/C/Ex6h4RQoTSQmQbyYvMG
4pngLlN6RyacBHpC0/tdsOh+8d6sdDLJh03/Nf2Ur3iBtgMInhss5iJBH/KO
8jaLjf6PUWZOfOmG6aE0k1DytrxvjpHHdArZozLAMSiPu1uV6zzhDMYcwmy1
BxlqfTuFQP54aacU6k0ID4CNDXtT6G8gaOgbQ56vu90rHC3i1ueDsnO6NPBQ
hXxW0gtuFtQLpRdYYelqzbPkqxwSfFSZiF1jFYQRPTw5t7IjsujOT8zxCDjL
mEsUbcT8XX1dAzQmFaq31dlKUkHY/1vvCsKTQ46DCVTLySbuCAfFRsnV+tc+
YgySwaXBHySBUJwtp39ifQ5SVqLueG1jWdr7GidiWulc1rlPvVbEIOS3W4kM
k1urSq2/Bs4Q3Z7Lm1d+yo0SeudYPtx44vqXUssY1yaxMV4OFbe6xSaxyoeP
rsQc6bbv5AhpEtHIxiN7fH8M9kEHiCWFtQQ5JXhgmbTEUvstbaadU8d1P7K1
YhMnrFWivhuCw6Ock1A4ZDgO0kuWIhTusbw+u0/EzShWjQoqAUAjAVrxFNbK
PNoeDK981xNRrxiJoZjH+2IRhcV8AACFdHVFm5WZdwdFbi/sfiuU1vHQAFOk
bQ0QGRRefnqZf10DVtXVnaibFCzy6Mey6f6GVwqw68o8jEtgbW2AxDA6dpwH
o4ZrxOsVQwN9cnsZENh2YMFCLVkQHS44NeI49M0umTku8ehhkAV5J51yDZnU
ptLRHL9M0dV18BqVHHu9xklpQt1FcpaKI9Q+1yEP87Cf8bqXVOsK72AKv+Se
E9aswa0B4QYc/9DbXdmrT0VILpv9Acqa1y7dt/dCF7DvUSkPSurbb7rfAslt
9M5cGhkhx1PYrm+RTmxk91RO5BF8JjX4bWa5NkoxNKqWG8k/QOibMDoAo+mq
o9JoNTP82J3gRBnkkHFnXUtn3K4JDHjvQwXMOIln5t+08heT2F64n9/QvS8r
IvPk/LBYYNHy7/nXZAYlr47Jzt79gAnDKjJkUr0SJ7N+aN0FGFA7KXDdEZza
VnRKR5bNQcYT4QLrESQdL28hIEPu1z4Mi6gKlOeTKGx/5K+RXVwnZcdpmpxg
8LosbLhx6Jg0/y/zdOIkJv8AKEUddo9QKL+iQ6UmiMqU+AaVgyZ5agS6JG7U
a6qau+IasmBDl/2J/IGgQNkCGx8xPgjf48toOfrJCLZmnTabnmNijqmsxFdS
5o7QOu79NBZMuFpPJOQ/YMlAnWawrLqRzEoUdoW5M9u40vFqoGwaPSg0Z2CI
5rpXljh/aO3LmKkpdaxF0b/HLYvvyuLxtotSb4x52skyUmU8H3j81lVgjUvM
UsU/Ba4eRbvglbiLSR2ueOMzUGUfa8MfaBsQAfC7JFDL81I79/1UOkLXG0bC
Q4npbo57MWY4PEHE0zvkWTRi+zFs98MiMPqe2+MwxctT8MeGLvA3DTa0poFg
URL35iyZiO92LbRglMRvhjmmDtDR3XKfiKAwLD0pKCmuEgny9U9fG1CTBElP
fJ4gpjTqLsdIMm/e+p1iNLuaVkfhjighW/PenWY8oNrXSaYnMkSOCE2jjD2O
4KDydNk4vsW4qLEgwvTIC6TFQKU6K8LuGGn8r6QgSqxY2Z+q0eFLUheaofKT
fF2F8x2GZ3mB22WpJyQ/6sN8ZQqBOYVU26dpuNcSKAITM17po/ZybQ+JYz9X
bV8zyrFdZig/4wptDBGWTRaMxlsUrxv3FT57cQ6QOFU9wAUxHUebF4Y9ywdr
/YLKADy7CpH0lzdcPS1pKpAgwMFWmXDQcSXRLk15FHFIaQwHC6tLb1S3u/H0
WFlU1WH8TBImfIOjDwmdP5EldmveENUTbqe57Cyh0oR922g9NGA/U/siT4SH
/L0LHP5zxyJjcYOilHdyZVPQJdvyXij4+lHatIRME5Hrre26MJCpDrTh+Tdb
QizyLbPrvbFBc0nbgzhep6iCQf0VH/WhCKls9ZIYgLmyzJdSfng6gYCgIsM2
KGsSTjE8yD92uarDVc1GU6peoH86BAMblQWmaXgEfZ6w5C5wrPpGEg9fmxkK
zXHJlCoHnrvClKcj0MSMmii6roamd4u6OnyBqS2mH0vDtv766Zpq50hAxPLW
9BHRM23GG9uKp5eyZA2cSbBDpctP1fSOhd00TCO6Edo976Cj5yhKImBrFo7e
phf3+okakZTFr6hPee7IuErJ4GxTz9FVwDx/n9ONqQXTujpvQY+xq63UBQIg
u5tzl26aedWVPcy7DmVrRB+yO7E+wf31bieByGXLhpirr3JrrxwgD1iaMuSt
tOHFplk10yb+RrBMkojucfht/Ns8ylnzCI+C1DVb7vSg9HzFUc/DLy1GjIvi
VHIVLPiCJqxh0jEiaUCG0dqk2Qv2t9z06ZmFTPRZITKwuM0AY+KWpxtxnIjY
opdOnjeyRSfHYzDIEuuwUlBoJ+gMM1Y4C73lxCkNwqLnkFeEcRUJP6SgMym+
LlBASiTtRe5c3iIA5IwhoxpALR7uhhY7JFhYSzvpogyID2rWGuWkpXAsQJQG
mEl5kITd7E7n7PAwZe0nVlyYefErRVFmetqZD/TchKemcITiuj07wbEiM5my
8BL7ZzQkZDHJTr+mhjLSzyH9Of+9xVdS4rt+gEZ4JUqRE0dVfNoV3EpuEDhv
jGf1XXR5H3XTNUntBaMfuJ/YKeDFvJMEYIZftZBzn4xE7xGcIayJAT08wVPK
SNHwyjc/RF63ERz3lOg51iY4qKDnHtggdWk9cmDkaiq5XJizRzQV95EffaeM
zwQRhCRLJ1lffqWHpNSKUOqYl1WIC/QXaIcfk60NohxIm5/DIWBG+KfYNbU0
gJgN5E4nO7aLrKhtNJHOPoKf9ogXs+sZnSy0eokJDgH0XyeAOj5Un7ld6+I9
JArpoHmPv+/bakhbrI4QsM040YQ4RaL+Auvkxou5Cqj0dTw1zbNUdv+WfvzD
NVJF7uP0VlNM98Htikxq8MLaJyo95tNp+QaLx6Fz6vefdWv0C6qgQmtU+xLd
fLimZTL0r2zd0dgsZgKX4D/xGB9g+DbzXVuCBPjt0xj6yOxG7SXSU5lvaI7f
e4DayEj4XxTETRmM9wKiDrxTT0j5JGHpwQqPcOK3gzZCvRkMR4cptjgoM/f4
br9yzXJ1jb4lv+zY7uhW3bfVQ78lY+2YTETz27a/n99rl2oleVDPUXEPZ6OQ
INQ51d06GMFUTt1m4yNDG69xUx/EAYQyvTRJkB0iK6YXvhTQreFAEoJGE0Pf
QBjL3kSKD66wI+KLsjIXaUaEixEx5oviAKP32xfuJIs4c2IYReUSJ5iTxmC5
fCwn7pwNv2kry5Dkvzzuex/KExY2vVHaKuE8wq45+qUcHs1Nym48ejkN5cEd
2nCYteR0b3YqSMCJBqCyTRitlA0uQeafp88f6BJB0o3mJTMQYy1Ar84dUOU6
LHap3STI7NOf5VQypJdZenOHcEnCpdRUqVV6imE0YyvClIcSwnjSh1QYV28m
DoCGNdW+nkBSfHRlDpoowcCun2Qru4jQRKnnRLqv+LKg1TyFFSeqKGAmZSRO
IJKcvKO3Gg4DaOdgqGaYaosbCbVtfmlt1Du0VqVk2QXtG7lGM/og+RzV3bzq
s4i5xFwTbXGCo5XFEZo7S3cIniID/cTRfv8/b6SsyriX2C2Wp71LZA2wcwFq
kaHeCEDRzEdOtWAMhvN1Sp0ubPfcYUDgtegqwaAwdMKbpwY2f88kq2fhnCCs
KQSCknY4vO26Wh4GPbbgrWBY6SQnSroBph6v86HjtKIA8qoH4XRshDf/Frk6
e0N36BKHEGOoVbqiG2sv8CF+Mu9IA0O5yUB2NjDkiKtgtu4o6HRJc/3FgLao
mdDX4Y892XIG51FQQ3dlAuck1KN19H7pFpDVZvnn/iIkPRuGDLM1mW8raN4e
Di0z+sAFAshzvqaT3xT16Av3LuG9wWZCfD94PrNXFLFKls4Rz1VAHnIwfpPk
v2q35E4fV/2I+f7ZQNrf49kSY1zyg5oTyOxmiaAe9Bk2TbeZ93Bg/FWEcuZr
Jlij6ZIeVwUubVun1/DlrGl8GPs+iS1exAO0scdthFlioZSkSN9z96ka7PRy
HnEIJACChqmQhUrRp0GQpqbSvWlj4hdSEffFlyc1tpLXErxDyhKk2bwZOIa/
n4CGYwWI2Ytc27O3PiEAGcAlvCr86ZMJFLIeNQJgvxq3odz8dgulOB1VZKGz
b7tIP39ENUc0oXO2vwUZxGzJ9gahvOaBX2u/oASDkGFFQDwE6aICilyJGpIj
cnZgEc6RmZK3eRd5eeZplaRA9SVXw8QqEuxSVj04bsFYUc0db+qElxK/vkjV
YKCq/W5xlNcyoOwy3q34b0DUPuaodEzt83Zlb1HZ2NZC4dS5datMyBw7s5A3
daDBP16VSvH0+QaIMCpn6tFhJz/VGHxZ7zCOEsRWV21mj+KKJpKGMIB45WPz
XvrF7ihd7w0C3leHmutwpt1LQ1Ht01gn3DNgqfarLT94IjpYPo64+Phj2gV6
McZe5RFNKFDyJOZyLgZYIafzlYBGc46IWzDKUYJoqZBxX23hwat9F/DJDStP
K6xheHHtT7k+syk568jPAle5Ah789fs1sSndcgs+Au24bxTpb02trnWLajIL
43YYS/ofdDZANQEDzrlchyc/gr1Dt4fV2ME4VoqAHXtipP2cbkisktekoLAP
ZU6P8tbFaGLfhW/WeANTMc/ahK4BwsM3fBR/Tfy64KTJNmrjvY4arBnjBqT9
RWvHfBbf9F/gIJEkI0o8m9G5DmeJt5ZjkEFrpvajQJbsHiLsRLOKmAgwkdtu
PEnOhqjv+2ywkn8Be+3UU3OolGXMuIum5l4A8589UG0GwYzP9M1/muQJOW49
6dQ1Zaix4lDaRmptQYqp4kNm9nQUySTu1wbpUZUdBVtpC4xuMt4EYzJHDzR5
pVDOgblMwZvX4R81c4SUCKi7HU0ZqXN/kRMSPlR+9b5Pcu1R4TZRi9sHSbBx
Npa064zl7QXqkj5xkYe1EHo01L6zN8A/PRE63c9noHnr9CJJcRBgdZtoRu6D
4fJseBblQhsM81IX4LSrRXTAxlbXE/rWGYE3RVuOT2OJNHg9/HDzgu4/VgfJ
OIYhFuNwsWAgsJyWam/yy4okmnjauAm+LK/qEO2dnUZrqAbVneBF2gQb49+5
grLup1ENUKRMDZZG4L799qGKIZSriFISUjFVP80ARhxKv760oRMRjSgE05/z
pBawdFBKyj0D1QLAwO8rcLayB/SKkTE+jw+pQ5s+N5fJOTl4p+5oy4v+C26J
qDzswOmxNtdxIZun+Iz3DLNfARHO1nb92dtSuFZzldx50wp7BPrii1XCL5Zo
MWjo9xgaUPJCJ6bmSfKedIYVynLK+BpeWt9PuEuPEWSK1v+fMe+hicRiCpET
03J8oAlt2ktng9E57K3XngMEid0f5BuEFaB372dCKjNRVmx4W0GJguibQyUO
ZCbiy7L6qk/IbsLVPZiCT6GL8nYn/XQi9j5JDnPGIgSXoz3FD76UoYTP11ev
BJizgqL3yQmsHUrKmO9NQ0qdZSU2pnr038eUqlp6mLfryUd60VaLKwwEwhU6
oUoqtjPYl/gt2HYLb8KdHNp6jcrCvZ+itQn6bRdIPrtFFdLnSmqC4KfixqRu
rDsH4kAmcGC2jqUmXDAJTZeZ8pU2HkQjkMzCPpT8KAocrTmsqEuJwMLbBLIe
N91/3Dj8nsnKiXQ/1gYzShXmwQqsosnE6soo3UESYobty8a/q7dKbux40n/V
xZlAVjFL8yw7pnrOePxXm/FfHCWL1y+qITMWlcfLQYPcMhLSaSvvlZNGeFEy
amY+CD7vRBK6JZQu3473mKUpEbbPhjmIbyZJfLzFMFdM3g+gd26iIrpvZzbg
okybKUZ1ROc2NtthTwSAPTHhGuoiPtSPELOyLU5N7Jk8Ixo2soENaZ7/VCDv
pDx+Fl494ufzQRtIaJQ0XvIm8PtALwUEAkp8sIPadegST5vsB5tf9EpfNLR4
0cr9ycKPBDXnaR6Owzfna3GVedLN2IQ20oI4IEsIjeSc6UyuazliTRkASYHU
HVMvIEsuz4t8JK75sMiSlRb9Necgf/oYMRsoryyN8mE3FEAycoFCQGbLEeEh
Rovc9TM+Gf5XyttvyJpDHX8tE/o6lLOd7WKuc/TaF5QG9/cLD81E9gAIyLWX
NBTg0gU52h7fFC2J9/K+BFLB4+TQrIHd3o7qpEMbaL83JeWz+uojUJRWKD9Y
bEorZ+RVQSk6gpNUEU8rAmDBzziLp1g+AM8JaVKd1wIfeizlEwQkXN5BXkoH
ylWibsiEtVMwSinRfg5JmBPHj7Z5qBm5TjJZhIkozapJHbT2KsMjLsTM3ev3
bJ6IClZRqsF317JM6cH317t5ennhW6DOvVmnp5eTj8ksWqS45Pr29erg81yZ
Goqr/8TVH4sQUZ9Qp0UOcpHWCxXIlcAF+0I2kKGKiUnntUtuyGMU7Os7t6OE
C5AQMMrJRE+vGyiWnLjrZ1N38aMGg2LgOOrC8hV7t7uH6vI4c+AmofVWo+zt
c6mk6ccXCreBfJQJzkZ4+4kkUTpbpjdwTW0n8E5ntj+hOi/A8Zz/9TbOTL/E
cqt3UYX6ySW630qUUJsIgH8mS0fRynztjjgge/RPjFVr46I8Q3O/amws7Qv/
LG60SVYHiV0pWxrLNbEhFnJ92wyDHgsHiS+ftUA16TcCsv0pWC+R9kpNiEc0
O+Srll0eqIZNkKu0/uDigtvV1hsY9BmKNrXAr3FcL9/INw3I5QPDJgoFf8DH
kMpGkaMeelgrK2BB0Fq8ZqwvcA4fzsbh117aze5q74yKuqJiO3/IcRmq/GsK
+sEKmbpwR/ePGk/dIXCwB35L7PfDJIi4q8/uLTnUj4czd/6cUGfMtbx1/Xvd
zG9Xsa03Be0kRSd3GyffTLLb4i56g4LnBv3SwAPMl8Mvi3wndz8gHlaFG7mJ
i5fhiOijZuP/5YNghSHFkluNYteWdapxUkFWQMg9vOkkTsmduyMuUKVKbXm7
D/ZfxHqkRYQcawOj7KE/posrV5ykWiDu9wMxx4qrrhajl7w7gupYInMn/6ru
9D8pGzQfSoNWlXNsPfLEqPg1hyr8F3Apt2nviEoKgmnQ5QPRcqj8hEJlCsNx
Ipz2Fi8mJFpgX0143uso1syIZcA+bMZC2Vt/HXzo3M+zsScbgytthYc5q1Hk
3iWXLbdaxUA1aP1p9DwMdxxz2xXakXTqNZ8RHNKQf9QLv5Hd4dV0hW627ITF
OjVhx2bqU3USdMt4kIqvlF6EHrQaKGzxbNCLEbw4+osFV3PtdONn+5RRX4vH
3MxaZJkVkZ0a41MSlAirxo26N4q2xP69ZeoVKaIYRZba0W88vJhBHYt02ut6
q0RWmS39DufYGa88Lzfd6FI2xrj3FUPC0nZwA89VFMXblFET4fJmmlbY2D7j
owDBPKi4OIh9PBbB/qIKKzvbrmVGdyvJwTPMe8PFj7BPfNUhP7MeWt9lDgre
MIgY+O7tyuNx0zL5ucF9CmRB1mLaTMXUuOYWfw3sFxCXLUypglixh/nXx/g+
iHaa+TKyo9s+7KVI5/F1nCF3itpxuZkywu490Lg97WIuzFxfSYd/ZjQ6BSin
UKUPRm6PwvEDux2fboGupDKUXtrJ5g4rInL6zqg/n+bNm9D2PVw8lwvyWOzK
dnyHzsnuAd0sHyVkjpT/jKY8eOgbMQX0avmvs+jN+tLNX4Ja9NsYqU8cFiyu
M3/4H4BDtgQRZd1y902xl2t7jwlImfWz4lGFeK5lSojIZGzk0b9B1XugzWoG
sx96zWa3sAcetZKjxEqeEVvykihMwuKBu7TYkBTH/FrbnGqoWFwlPIwogLL7
W+M6lEfJC/Vp8T+5EFQmOE+8FbPrFSxEeiplYkO2Iw22fMoQVPeYqqPhhco6
gQAGYkBQGpg/EdrIWTOK4NyTVebA2nFEDrl1u8RULboDgiSOpOzG+dW5Lihl
wZ1qUXEQ2oXDMi1b4URcWjt6GW4hOYG4TwM2woN/pN+LTaUf6cvcfFUXxth1
LtpcZAHkrcPvSxHUZstQgUtoS5QEbZlpohK6PUs/8g69+kSCUgZSu78pVt8C
kI8Gky9Q9Z/xAE5Nz6zoyucH25X+UvT7byuYia/IAUm9H9pQZi0FxOFq05k9
7w66hogTN2+ylOPD4+Y7mcLRB0h6+QsBtbjsBw8Q+e/atYnaD2qK5cH5jraq
HHjAK6vWh5GXyNeW2DC0b5ShuhpCd2GFEtHOMMf63kEbrkoeIg2lavgaT2aD
KBFxBQouYgQl9kEcxvXsYyLneR++f/P7amSegdzbc6ZizE0OAVtDBYF7500A
/rTV9a9lc2pB+O9UZLBlphOSQbd4jdXnoGwRwCxvTQm7hcIWuKKHA9021e2/
Bwcs47QKpE9Q2GNcKY3MK092x/9moTlPjaBcawEsL+AnutcNKHaoYdswJkWR
jXB+qrXJKp4FqiHipWAfI6+Yp+8frbYKvExXsjOgBkkCmgYAnZfvtVcimp5C
edSR1ane72NcZ2wF3lzNgiYc8LkJXK9geRAx2Rsh1bpfhR2mHhCPKG/jWfne
UyS4Z9cg7NGZhshqkzV/AwTQfS3mZmpV1f1R5k3jDuWhDfmjN3RV8PAPGijK
SJ1lHMHfuyZwHKAdfaeOQi7rVZGxwIGJm+hRLYDWhLn4mrCXHVOvrfBHuxWG
1iaJZF4W14nbjxqfa+dn0HoTlEqNmm2etMKxsJfYLW9/wMb2cbAFZaf/VNFV
a9CRtP5m84TRUVVnjMkM6in50GLHw2c3p4XfdXXWmajlNuqvIiWWI9tr3t1b
vnbxWgu0Y+5ojRX+vQ49UU4b79v/m+D2c/UMfzFoW9J266fIgKs0Qsx1l3Tf
o1r9Yy3iaB04K5tu3OuXlDpPaTI6y7MYJZYSMV2Fj4VqYc5KJA5LenexUHt8
tWB6CkuHXnZ5JvBBSfB3IJrtl7kp620XQyxVicu9CbEp1t9/rGOLtKVLiiRr
LRgB3BI0oT+p7jwmqPduIEMfka3FMzOfMQx1p8SxHLcRV9VRG8XEPglW+urv
ytwnmemZd4VtWCjXELEtWMWRIrwkL9SYLPl9mFdiyxJSgnVg1IubYPvYD5Ol
YldOb1XD/6Sef3Y3a89OO4sOs96BZb0EXaWq7kO/h5Mhefvz0bSUNJVSFuKH
qTFta57Ngfv8rtVTfffmwqruynNn/2UABJbsD2OaR80oAC4MtkhQBt17VtU1
vs+H1PAr3tNwxEjKWbNBPke8Hw2HHh/kD25hd0AymuYtOb37AJXUsM1U8ric
gFImtBVD0LrGgEph2KaYbTeNtRtrrAeB8i0md0kCTtcmtTrQ8LHMfN86emYb
oio7GsuVDf9hO0GFxjOvuomGTqd8zAII3cskKdHIkfU+dWyH9B9JCVtCeyS7
W0HJ7ef8IN2rkNYBcOgSwuv5qd9v9lDhkSlKGwJbEuRW9mCRSiIrXBmGHzcg
GlwOLkXPmbTnpaINTL6wDQtctEp39pfzi01d3evM95Hw5jGajehgkuax9+Sp
Y3Ir+0XmC9IMcFOc0/EZRd5KpKFuCHNwqGFhy2Scdh0De1t4fmNAVrPzC1Bc
Uv1ZBUtAuQHoyx+Ssx+lhVTmvuKO6982GnyVe/wWf4KBSo/9jDBtQ2EmkuZn
8Vek+jbjjacnbKujyW8tp6zM//xohzhp3yN+YSZvpfa4YVTAygg7jEZH2gKq
pvXU4wtUpF7R6D7EsK3irZGTh7W8NgtbChnqfSMNXroUJ3YueNgFoGx/zIXr
5XuWRBiqWSjJmQbUwducuVEqRdPgaeSDdTVts3usyb9dY0xGsKZ+sZyOUzEI
PFKLjsXjqi52a5HjQdv99rIvYtsvCzkabfswNCu5bJhnD7MuFjcrule44iut
vYoz55hcAx6WLThsQDciUGMzLAoxMb8lP1WCdepxG6Grz7sQIesCIsat6NU5
nbRjp6F7YBRNPu7i7Xs64egoCiBO20DBBOQ+kQngd4qE8aCsJqvZ3AJIJQz8
hztHNNRDRJtEozb7CH0mcGUa9s47bXYcha37XUsadCUBM5hNEuyeYq/tC9jL
hn+c0Q3ATLjnYR93L0L+gMH8uADQL1pCpBWSFA/5pHRP7Tgdq57eNkElkNjk
9qnUDHKYm3EFf/k6gfauAqbZTAtBlLm3hi3d7/rU8zci1oi5vDjNQhfdXTzr
8YN0S6aGqVcerNjp2I2gdHSAAWEU055XCFHX0ujvnLgMSSBkZwd1Wcc1BAZQ
r+n8XFpZuUOsqJ7y894zrke3PPWXVAggy5+uhMpfsQhWtpKPURmKlp/ryTb6
oSZGdiQMC1KwyxGlQJlZQZ5S29oIWDsIxQvPjZm1mrV9C1eYV1s6flJbcXBC
YDIuVcGaCzIHayqHb2gsI9ZrFylno5FAVSndqCVeAYEeyb/B5mxeqEQ+QgVm
HO5tMQbnd3D/saSSdngQRPPDpLhl4eUBFSlvaZ6GN5768bfIxzf8ciPgs6kU
KDPy2tg1MujOM2IQodk/gnXGRC23U9a6gVpUjVrJccE9kjQQ/gENqVpUanPV
pYbgSwkv7AYhLg0+w7FG1ianmiJyyPuPz+6P+PdlsXp56b7tGYx6VkpquXVL
B95qdPosm+R1hrQBc/CqFYlmRy9FIJntTj+DzCuX5+djZHXHmdPVvzOiAmJ3
1lDdvBam/mY9dVgbG9qudEqWjNP5XXJVk/n/yxZUEhNUynx9pXMerB9tbmVL
c25/uliUnypAW4Iujj3XEweeU0euUieHGAoIteKzJHmSVabGixibRfC/JmLx
9x/seZohDhP1u/M2i+edfr25u1VZVh/EJVaHew2+srZ2deITYyYAoy/1qOXb
AhCrO3LlC4N0R84k3RBYDqYh47FzWqXZSIKGVb7CVz+14IVkhS5UD8opHK0t
Ijs5VWfY57Q8gHJU42Xy0sCbGqNV68ieTzZ6jamSwo2UjDk/bp5wQfKHAanx
HVK0U1nVUsy6nMCR4RfBW3FiibLR5HrGslqn/r+s/SI6CP5USsy1KZP3hs/c
ryxyhu0r1wGf570jZSFtEcomf3pQmWRbudYyQpQB4iumbNMuQETKqfLkAKOL
/hugyK+PtK9by7JFR0Jnfz6DQ9f5pbe0jwZAYYaRkdnELFDg6wd6rM3vR6jL
1bWC/o3Vztg5yVSwxi/+eVc+/Uh01geOBRPTvON3cATdCLWHK6QuHKmrLzM0
snhAB7CqXCUisuaGlRJF+zUXYWio+5AbyWobBx06adtzMVUANAcRcooYORJo
gLFZpH9DQ2U1Ix/l/2AZGd6dMKs4vWuaY3EV52NRQy8ipvTM6R7RgcUoIgzi
3tolAoc5Kmv59yJjtrtFwfthokkiSKT8rkjGbEO0HsUMbj44aSEPLMcnJBu8
FQIIMsf+dQY9+IVEgReLAE03PFeW4BwH0Wrm3Dk1WBIl6wA9hNrRo23z5eZW
DuobgOlO/QlSF9T7d+uCEGYQVyaj0ylokt/rQ6+7ecIATaYWmSab/85t09cr
iCRHhK7e2gd+BzgEEt8SQkD5FaoAlll6nga9IQZeU5pzMa2np+cMA//Ywl0H
acfB49bZY823z1w3A8cXCTNFvOQq1g3AYS55DYSYyxAE+haPrBqj65P3uBYj
TLa7YLJdqihx2h8fI2k1oIUQuSIwtnJxcitbGhWM+2FoR12XEV2xQqBTyoZt
wxDrZ1QBajhPPofrTvjDTlnMBTKSh1BJrScc5OM3utFupY/SftvdJTg0l+VS
7dexSchSO6rNfxpkPG0ZnXtKRLIlLmU/NlyHKFV1W5Sx7SZkvOHzThmq940Z
iOIsYdb/vmQ8qyniYYdGSi/NuuV2pocDQRvguKfSGGaiFQxsOz5laFAxYk+U
X10Icg/yrelLYQzlz9ZJHuZ6q7Ourv6I4q65zackWy++ied4awd1k2Kmqm+2
aHWaoe+jHyab7HS6nLKYsKIzMR1r4/pqG3GemzzqnLHUJ0dLk7xiWvLPdn4H
fBU1ekrspGzmjbkuCkd08Z0NbkoauUs6w1KesLoLcIDD2RYn/moLKNqglkDl
d7t9dP/IJahUvYrHVMRa0Cs2XECa+9pfAbWBoa0qkGHl3iIaFQTUMt8ImsZL
RTiMBDd1ZcdgAfcG8NgNYUHkl8FeW65ZvokcFuhYeWzzr+miFxOipRRdj6v0
i8pE1Z/uljQGcnlq5tq8pv7EYm2Befc/YxWlOHHi3yM8MupO2xKHSpE+z+rj
rXz6B44w3VzViVh6skrpTFCfOPKSUsOqRyP3hUgfIwcXxZrPT7FBN/vw9uwo
60Z9B4ravzfgBRzL+rcshoSRSEB1OweyAtaJMlgVM4gnyTR1/at1MRTpOo2f
Jynb0T8hFU6ys1/sY4CKnFw1HTGkZqeC/3ICGlBPO17OeSyOzhyXMUBla+L8
WXokzpocX6e8p2GjmgNilesgk/ygR2fHYXYk+hsh3PUk0O0lwLSQ3YNrMfkg
H0CVBO9oC1VQfV8rS4OWUd58AuxfqShZR5Gcj3xSgystAq1YMayybbb5Vv8Y
fPbKzXZW/PvpoH6qSCs3zJb9zUzTWzppjBsZHlxcMkoQKZVnP1ObBV36GJmC
/VulmZ7I8SE0kle2u3+m6W9t1kIRradW0K23LemYuaWVeJPz/6b6mUoSZJSN
gEnyZlUNku1GAOuYlPzdb/Rm2GWazmNlxAfCy0XLD4RTrxgqKemmAVbwMdON
a4cHHDDazmkFrwcDogD3Dl6lBQFaS6oJqDCuPsr0Ee1ORAGnSUD4wsNbe+vs
Okmw3we5eNeGMNcHpWw4nq6XJi2JMAQ0ftnYbit+tRQv7grDMsuMHiLIq+Jn
7tn5tu9dFd/fHpKwUhXGqlup83OGkl1obSXZC1COyZxrNgRj1SFxsl8pqmAa
Qas16kYFLy3uiuQcgqEHDpng4IGH0Vs+S8KWR6FzwzulReJ/1DvzKmPtTXKQ
IWHkxLdhTdhwO7sn+zIr4umpK2PNiWZTYDOLgzEaWuz/Omk8XNpBf7zzhu2Q
p5qi+DfpbCT+OyRw+xW6OmPaSA/7vq/KoBwQ/n++B7ej7RkLjMu8UF+6/RgH
LEcKB+WcwXOFzfqS3aNr0vuQ3Wq40d2nC2wNiAWW2yywogtXe1/3Xy2fKWzf
sE4D46COD0TbpbWSuZ309VudUhOAGXJxCFVbzYy65oe5Hn4yQRKeEOzRbFK3
OILShoxrTPGYrOEU0ofoiiFrXiHlxePZlvNSnCFCTr8ZBHQxno+MhidGF4NJ
0Z2GgdSD0a+80dcuOCzOvYNgRLkpGtv/wRdQSPCyO9yFNb7EW3bmwqDFSP2X
CYHv29Mbbqvy9GRAGHPDNjkralA8x7ifmyswaBGGfcmUYFyON90LE+zsHKQG
YtABMwboSuYAFEAPK/VFdTK0sIkzFVG4nf2MldRyNukbdsNxyI2S2HVgUtYF
sbxjlTqMn5cy0DdMdYhwTk91x44FBetPP1JpMBtO4e/lQyi8IE6qtvVZ8R8d
cLob8ERkAKg5yssoOkfEfOAuUo0dPFAHGNR9N4+2eR9tfNEayvYtVvo+OR/b
YkpBEKFKJinAzvBzSrgPiVa2BcnO1SkmGV/au6toSxZruAGt8OcaH0SEgWeU
jaJ1gsD/h6wj5+Sx19DtyFREutVCx/NlBYt30L09ZIhAN+RACAk662w22Gzi
J3pKMywEA7CIoO6vag4LmZYAuHbYE5FOZeo5AgE+K2TNaubUUoJGwEUAtvI7
sAbd71bnJ1GpOLWEqIwM4/kReyrjRri2u6pa5vfI9dR5qA7sxBLH3XNXfnUZ
ktjLwErPvMs6zasPRL6+Y6MmKUjOQqFbRhyCy6nuja2WBicDY6mZthXE1bfg
XpWyPQDi3dnz69lQCMkC4CJ73TPOyj2YKYI3+IAMZoV8wFXPW03iO21mSNhl
Gietja2YVEp/4cHt1I2aMw7cxxsDwezrH1ILQYFai6NY1K/SPcHqJLyfFEhi
QbOxzDXw1oMme85ZbhZc5gVVquubN14zfwt5iSEZBLRupLvKsZlpBMm7EZQE
V3C9m11NSR93Do1l1YSeFsiKWtQykbsb4bnfkKhRaKLBhueVTuJAX+0yNPy4
IgwMT6B79DeG5Ralu9ZX53qVOg7tVwhM1Aiw63YZxRH1/d60qNNKEbjQylBs
2Vpulq9poiRb72I1vfIeLaFHjR6qu1wGNnFBtv1vBRPhjFeEJZeIyhT1ir5p
8CaUJsPQ3MqeAnaiZcsxhnbEWcbZTnDAZt/RqdzLe9or39UNg73DCh/UO3HZ
7qwlxlrRFiyEFpaeMtUwJeeDDdhZkQDiZAI22n29VvBDjfyYWYJAj4MYtk2q
6A2PgDQ9yKPlubd37bXMwwO0TAoC0XILmu9n+/0fwizx22hrqP8Xc9lt2wiB
5GLIqdkbGyCHdbnXghqZaKcfA33PdacV0wzuz/36ERV1w9wtL0ge50zJCLNp
gAmEtXnoQTCrnhjAVWHrG5m/c//H4qKAbP6N/GQ/DqubiiCNaRCPDYlfethm
kxPFOOGkXdUotyRHpmT+Rm0N1/jcFWv+kZNFMR4UODbm9poEy3F0FRN3Iy5Z
wgPGQJm6OBcJeLmVBgoggGdI3RGCXQgwZ2Bouz5YfYb3/9DkCbAL0twAQeqx
AjoQt06U0DupLzM9VGfvzu37eIw7M4J+Dt2e0Pgaf7azdvZm9gm0NaIFnt5u
MA5tnbUDzSq4HY46Zsi8i8lhJtp01nGKdCP252PtNjD+z3MT5NqiM/MtLJZp
9j8ugxgsTFHzaUQ0pp/6QUdkZbNBwBUDILSewsZI9JLQ/grwbGIbkNYSH2lp
gv468D15sWQwUuz0xyoqlhKvNj79kb+c1H5Z7P9R2czoV1uu6hxlCl8t62K9
sgCA2iZAW3IyBRMFcYc8ghw29N9cCO1u52ZiP5WhhlHnaarpVpBLTRvAbSTA
dVKOnwPPiCPBHDGqXcnggVbfJTnbaU1khp0PgEI6YPzjUdCiP3yM/m7mHc6T
9QZqJq4eOijgzpV6cp0YdZ95juHMKadZ7QPYSFgL7owccFOc06jHmBfuXg5r
YqYzTwf1AwnHVgsJnbEsZn9+v7RnrzMsHnPjXkE5g9sMKif7JNLOuDOsDeFF
/tEuZZADmlTf7JDPEr031tgXLG/EFjz+iYebbNf7McMsrTojh1F4aWot5jdA
Z2xYIXa99v/Jqi8wXHgg9Rn0c1ZmONcWXx8PIaV/pnmnqHaHDoPXttp6MDSG
jqbqdM4R+ngLe+a4rR/x6RxYLpTT7i5CEVUjg/iyHgTJ4IOW7w89fcpT5N6Y
fXqXofnBc3ekhmBJVdgKvc53BXBKe1AEDW+HVo+yKRUBDpD7SOIX1PbC9kyg
12E7be/YMqXYZwL6mdhgr6/Lf2CoGtbcdJQ6o1tdKanPnNTGevhb6gYzGZxr
QX0Hw3B+rUO97u9rxzOCt8J1b+tPNY43L2UcbKmY5avUN1buuGGmcPBOI9rL
+wgS/xghCQmWsViTIMS/rAzprOfOQzydY4NLveIuVA1V373D9kLjAxFWOqdS
g8hDmmQRzypgB0DzPw9Rn8DkxDkDK4SnCr7GLNPIu/TrvnICH2fT8ZtUmEeV
TM4tQFygDKTdPDh4sK8LJUNhdEO3U3dWkcBfOsqaFwNNq77aqoWm+inkhBQj
+CgHS3wspVMW3aBlpTmBcwTLt40awFOe585ctlaL95MgdE7/HTLbqpbJXP4J
y7RhCTUzrbHWZIBcXgGiaOQO+CahHh/LfD7IWbvPJxDuCA5VZkBaJQFtPuSt
4hNY+RglDf40+/VM7wArgc5ZuqHBB9Bf2XzfEArhltGUuWmtnHqdeAskcRB2
GIVEKO4qE/2GFuxEUpH4u7U24QohZ/dLlLfkWIvmSsol53Pv032ubP5yEydf
SWN+y3zqg1LFOdtgTt3/L6X/AJoQCWBJpSRcKiMCh1dY722hMSXahklnKV1m
8O5bq32OM+INc/rZuZ2tX7ub0+cQ5UhF4PNPkGVvAE2QeS7re7XZtU06n2He
7ux+XYhfP/sMkVGBrMvuZQQVqNavlAIqBQYqPPK93rOJwpX0qLCZDo+F6WV3
gPrE7YxLGZgm83hXMtBMNSCRVKc8AQj56L2YDypv5EpJKoFTk5mxTcDsxpaK
zXqtn7DdjJJCH3ccxS4yns6A+E1vgaMLqZnciCdJBWmr7SMQS98OcrK27eEJ
+r2eXAgthYgA/+L2sJZvFwqz79xMD91BhpoRn02Uz8/x1o6gZQIp/rMnLDXT
7Md2JzSK5P2mOVCrK5xNMbu62F+Y34wb3juh50HdhqmYbKgHBNGLKuR0f2F1
NcpCjDtsSbXGwZEEIt8e2U2AxDrcykwaUcLaw4x6VvCJZzXTaIAoInMwFxVB
yxYhAgvanrL+OavSMcCPaZi/OtE4W7uLflafIjfg8VBkwC8ne6/ebufXGmmL
pkm6NFfXpZwb0B6v1uIef1E0Y99fHdHwpIsPoEFecXucD260R/X8fTH9BVKm
xT6G8Ht+nupZBsbAP7onsxnvqw0ZL0p/hqKRhGDEgynV5zEOFZLC3Xr2y1oU
VSV8sjDUx5BFPgv1oorhRl6NbxA925vlnFsWdF8VPpzb/+gXGxcMre6vBufp
Z+AjDStd4TPD4m3Judy+B1luz/v2qRYDfRyDaoUFs6kzTA3DDEDKJJezEvWs
WJzgLbAZaym+yG08kUoAKYsrK7ADn5pKWCBI00dJZv3KSTXoaOUW7xgNQ1dz
EWFL/hgVxhjXWOwJ3Imqa4U5ryLCW9t2G6pYW+FS5HKgeBGNzfqHnU92Rmhl
7tBCJOLs1YadOBLLirCEz6P/HolM4rQFWkko1HszU5hnXpXzK3WFU31mT+ns
SXwCpmWX9O49atDKne7WJ6l+d+MkNqQ5MhXRcCE00GHXHGqBCdPxBHsV6sqZ
sVl9rhhSrCMp6+/etVAdR+vHCsNIB/kT+33LiPA9pm1x4Mz22EVDe0bNMUA3
5dLUXjmL6iKXR2Q8C21ySBSm/stbfKHJm6IslE+3rUhk36zArtW0lLWpBGgL
VEM+/QaGsIcV7feHSaVKHFDGNYpdMmys5kKwmMUm39R+KXlZzXZC+3Dp1X9/
z+bfgGL0ShK0BS7QMw14AbDmFpynvS9wwHzeJ6c3S165olStojB/lAx/jEcu
TgcomLRHSwiGUpfAwxSh8z4/3rbaW+upt4CLlC63KRDqdEtV5FajeZ7NDl1j
di0tFToardf3wiZC84oGTEhfLVFW1BqxO0wOgqRN9xRHSwKbrKnGl2Mtkv0M
cAlZSTgv1jq67sTRsQ4NK62xwr2PvB5jYeVnpswpcAMzE7TqZl1C7JH9Oxbs
NzWWp7dQcxCrVAML0KAfUP2FUQepeyCvvZf6UVuHREtoRtntz18tPXveGIe5
yBEdtfmnrNa0GkHf6fKIWnYOLvqJLAfhfeBLU3WfBi5LyAW03+gEmY3AKBcL
qhO1/jvGSrxmrfrc9f2fuoBe20Hmc/eBx7eksly21bv0vGlmmmRf1NC1Bz07
3WGFXmkykSoE146JaBhDx/vn9jEXC9G1NiLtQ8r/Qkjaa4bTffyJxDDMnNMB
q8coJ0AUN6PTGRAmObvY4agUMB+5fHaV+c1cYcfPNspXIc3KQFH0t7WveTfh
hwHKZgC/hJsbk9LO/uh58vVKZAQc9qlgZXB4r74QLaYZLHviidviU/Pi8S6V
XKbd+ZD1qEVUnicUyYrEqjCX6FQG0yrghYSq7r3UyYzXqy/Msq3RAQK8DCwC
ABVr4DlAz/hPB45Eog33g7SfCATdIDqaMObzjVP69ct5rv4rBbZ+sRHYwphx
buKuMyRLx04/ot/YXCOyk3gN34FAaLRXTS9MF0Uhpwp72X5UILY02GaD8Z6H
bC5YfiWWFzx328+EE4odK7QYDCIzEapvFHERmajAixS3QCkBln3P1pxPCEaR
VIiXfqxVR+BFhuT+rsFxCpEvciv4TG6CsOwbaxVq9Ql0P8Jkois2GUlMq9ON
YFw3zmLl1S/7Xypq0EIRQVPpmpbGXj7gu+MpkzURC2OwUxfGw7OOMiBONBE3
f8TJD8i5L3zsmpq4igtDjlNqO0fjx6GYxomfZ4pW2bgx6t2xU/515zvgvOv3
EB/PrZK9cf41Cj5fPM4ah/f1z3OBPUTGCN4vD/IpXTfp6gZ7ftJnN0NuhYOm
OS+cMJlOlIt7s/lJXykB+g57pF0lp/Swk7v2GjgieoGIBnmJWUX6pBQxSbYu
qNc4Wh4Z24hvmFacyWnf5BpZbaTKqQfUfBAGK/ubq2s9cQGoqx5s7D2iy5ZY
k7d60F7nEAuzqcg7LLwtmpPn7UuJ4iP6HiuqOW5qt8DNF4hU1ZqMGrRoQehp
yNCzICjd8exXDyQM3EYch9b2MlUydvr8JDh3MHF4DHjPUaZfdj7zwjLrYuAL
Gz2lUheu2H11WCAJijsYSHgFoXD7nTCiu6PMwa2g+gzTPbjRRCXTOg2AETZz
Sfzhk+jo3q0jB7jXPGL750A8vOlbJK+RcPgkVgd6VoywVkmASFjqV4wFuuWR
NcaF61VLl5vsUohqtb7OqY6uTozDcfFpdhhoQWBVRO0e9iX5cNRyWlQWJ/GD
YQcXUzV9ARAJRUW7DVPxR3dg+9j79LxoXUz6zpjeHX6UeZ95IcZjLYkiBIk2
+qIHtKLYMvuz3q83XcvmyMLPk0ajBtRanbfLY4PndD7npH9l63feetiwyDaA
3Yrn2cBjBu3D4FfLn5mS2cKmqWom8eDVSeo+uGZd4C3fzLmfENmnettoxrbk
iaJEFb53v4FT7uV3Cv3yGm5rCEnI7j2u02+iEJsTlnzQXQTX9JXXqxkDO/Hq
c5idz81+gPlM5iR/eNyK1uMCTxammuV2nyZh8GDW+CTZPxo976hiGYSSGgfv
kXao6nw4VmHMUIoWFOdUgWEyxW8dWnDW1OhMt0eMvdkm0VAKhyw+5KxBW3SB
jKMPKxhLk1s5pTEkC7YfJzW/DJy0GKyTcDdmdHvHarnbo3w+p5YudpUb9eKd
dxy+kNuhvdsbdkhUWc2A3TgrggAEgKWj6cc+q5bdRm1hr0cy2soE3s6oAnET
MD4GrARWHn5nQgET+6elsjS41ebCx0plr/zAS/mYRe9TkJAm5ua1hjkGXcIj
Bm2vUTWgMY/kYjbXQEjnrHn5SpdZqr0DZtxRzBOAUzjhMjNZg1UsHXqVPbDE
/jQYiCszmoMEvT8yvcPhk2o68FObOgRCq3r2CPw/JeAXHHJL75+OMLIfruZu
fslcY+gIul9irozr4VNwtLFLQrYs945KHsNf8NzTvkdVy9QZG0rHVtJhGTgx
GHHzjquqL8Ep1J4POW3EtQs4xvkJB9ha3u2CwdHcUn80o+4rOVrvzzEciGhR
vYMTzNWJWkrAcuSCmiH0Jqs3pCIqPZ/1J770EjNSDcNNyJ91LtWZv48AXg+g
fckQSR/hhR8U60asgWaYleWt8qzxhIyS31xoaylCb0VljITEZwQuEHWHUIRJ
WmxmT4t9vdsi+9yDYmAnuWz0wLNeMNdD+XejTISLcKGPO2RiRlDKoXY485R6
L95jW/ABgBYcAtHUlP6KN0rSejXDkzTzZSpPPVVNtQq5khhcPon+GEOZ7fNR
6oJmkBhUBvcBkp0CbTf7+Y2UCTLtqm2y89sEFLPMXRrlUKyR4x73xE8ovDlt
CwVjk5eJycxlStFobSQYJpayoc+UHc0GRSI6QIfdyBmpzqiecMJg/tTtf5Fl
hN9UYCdP285NJy61gpW0VzKi0vdNt4FhdSvfWvXrfRw6RNOFVVCwBLLpdW+n
G792h1pc0uZBuMSpCfJ9vfgZubqpeLaHWft7GTYVk4bGHBzkkdAC93JIQVlK
5ZmKhJyOFKnoKxJnbzcc8qZk/05ACB+5yNXtkGuFj1IRCRhnoa388cW1An44
NILFunEW6Qu11nJPw2Ql2enRqRqEulzWD6wnayHvn6SoHssRXtNydCwmL9gu
SgK/V4ayVps9lw1M3gnWeOKQUp67uafYQ1I0lRA5IEknbYcEIv3QF+By+1MT
N2Befg8QWfg4CjnQnCticUu1ADg2whW6/zC8XzFUitck9O4qyoegTKj6BeNa
+/PPe85V7xWFqtnwh0x5BwlxSphELu1a7yRrqHy/+AXJGEov7Zc90MZeCjfZ
cMkmGfps66wP0mr7mFL6PtRG41BLwxYF0BCXoPbgMZVcdJNJ2sJ2AmaBVjKa
NR0kLYf8OulZA/PXY0KsryCiK1fXJwZzWvQylIOP3mJgsUFBvoIZHB/ojKgY
dV9xc6mOShAXjrtwFKjG3r38fQ4WHCzsB1WImmiJ4pBum6dUJ0rEmHzfuD89
NEnBQFnrRaygeC0RpaMpCXqW62acyUIDxuzjfzithWsKDxjnBhR1bZjBNevt
L9Ul0IYe/No5G79xHPp5EqKFxG1p271u3T0YHJHQB5LuyHT0QbodjFDnMf3H
lkvIb7E9dG/E0D8eq2RWnKFYoA6vv6RZOBkRKi7KyGqjE8yIQANym2O2TdZz
H9CIpY7Fbt6wYF8RXR5opxp0JVoryHlBrgd2c0TTyXk1peM0hMVcvzmFcw2E
NGVMsJcVdQ2hzA5Vjx1mrVwyblMOHSk1zMEmpumRym6/qcfR7hxRC2SfL0hV
7DZOSAVwrvjw8SM1gFgKruMLYAkAT66RPTqlQszZ3ftCuQ0sXZKkBaL2HCe7
xmeA7o0hGTMxhKKmZsU3lDxIKLjEe3O9gNzDfTnTV01nCszCjp6nd5XDbKQH
9S9repsf12ah37sgKKDgP4XHE9zMbDWSOK2EuBwQgVOfV5FOc/y5WYnAq4JI
xV5+NHTlg7NPyaG0Djk7REmK2eMiQwaEtX3SUoiEkhD06Jg+o4xPj4ZVygf4
k6kxMs6T4+ZlXfowpiuUeiWah7zRET+1lO4amgjlE2/yymK79VeMirdoT8pN
FSHTCFVRMWFee+URUTTjz1YJOW3R5k1cHflCqCBtmVt3h/ROqrjSRRSv8YP7
/9CYV3aOoFfsMQd7t3g5+AW56NzojS7vxLRXsOt4lRRUO3vXkVb7RHuRThmq
8yI8jd8mcYUQ99fnVfLmBXuKhI4FSgYodcTTHEUDYqX4kfEtbCzI5qNZdi1x
X4nNnJlctR75ZI5ZyuRFL6iK7VGpJZZHdYUTT044mMRKCYI6yyzNCsLtqNd4
xOdSHqWJOZOOUgg0ZU+REV3TUr5iefWBNK491U5PyD/cZyeFz4eK3wOEKaio
xF0VAa4rePBvVrBfskFszMDZMHSFFOHYkN8yRmJ6U7gXnxtqWR5027MEPDyp
AxotZm9VYGG2JVyDEjgdYQOpdX7GNw57ePrt0LU1rJK/2JWwjSARfeRyKq+n
0vHUOjYR6PI76+oTbzP7GfTkdU9CxFkTwG4f2hpyIDRKU7mtqgG/SVmNMv99
Xnwi5IhMc/lH8pswUZ6TkXhY3cExwmJGYn9vwhIBK0bgIqCVcGcFIKlmPCEe
D0N2cN/O4MCbb08tTltSh2VFHVmQZ8gIHnjZqTF8cf7En8ENlgYanOszfVHT
R04X14TdbvZJqGAzxqhlcM8g9qaDozxa7mwERq3rS9Pjzx5raGVHZIGE+/l2
nq9CUqY9/PELs6IcTzmJ6lTxfty1qlSTxoAEmOq/5tLf8kCb8pO5PdWu1J6x
NIvsQjPVWZ7GJ1nDN/y8gwwhKBiMDArPoRw+VR7pPhEC3DlJQ1WEiwBwBvfV
U5dUrAeesjrFR+lZ6RBMwBOkpQLXIQ0nG9JygUtK0R9DOCme6RqK1F9ZU92D
mdgY2zBfU78A2TuTtR/5FF1nUaPuYAxzZuwtQw7bbCxo0OyqF7P6iWuRtcCK
9YJRnnnVxdCIgWWldaYm7ImZER/ilnXaTDba9sUJuSNJUQ8WYtJZJ1TB4qhN
xdjkz7B999LKp+0zPwTIVTJHgD5iMU8TUS+PRW+uqJ/MhzFsonQ+oUVGk/ek
gaw0/8Z/U3uV+O/6lfDC0M090Ze5I5tBy3XCNDFUBWnxydTNgS+MUwAzye8a
XUC8TDCyqzqyL4WWUMfMWEYH8ojGy77hhKcSBjX73ZdV5prc3fW+YbLzrD77
asgFewiVn5UrlFlQoYg1TfNgkL9F6tv8oG9sxdbGSkGCsa/q7Ni+qj/ANTW2
DgvRb9G8YJ2T6mbV+tSnjGX8YZhEQIk7/7ubrxPW1j9/3vHoFwtgirX4kCYm
rML/D2HJySf5kE6VElaAPOQOIi3VbWIpnd/onB2sYCVYJF6Np7bFDK7sDKY0
sxK/UBsLPHQXjYf4R/+/mfc2FjTvdCHkl4tJZz5YF+PNOFHtW9D/R1l2LuD6
VOqfQtAxdsHa4FiweMrR4dRdLqgdhXB5tVpX6hGbCM3UQwNKk+dHAxOwEWfR
/9gb7pdKSmVFNsqKipNSXbZIDf2pZhyeDbQOj5Mi5ONy1AST3c6FEDZolaOu
DzNNWwaTtbZSt2ULXV839eFvaRRSESYcu7oDL22YwJQSB4YX880Dnyt6elTl
TK+JXNCwNlUYYMAKkQJNliZBjlpOqM4f3f93IbfF659gCEX2ynfkFObm1ygs
i/xeGqnq5ICkIaLRwJzMKgCz1W5wVOQGtyPJF6ubGSGuGLukOvvTI127fVdP
F8FpQxBDh5oWIYdHgPrn8qMD62CashPRM7QbPfXWsPb1otTOg4V+K96M+zrH
Paqq59jhkDDRN5USkKamXUgeljL8iZQwMD8Rod6sIiQGn2hKHjQnNvp++yek
wLauumcYutc3kUJxHDoy5ItzO8aN0jGlSP0ob414FpsFDicliOAcJ8VDh2oj
OJ2LleQSgeZ8qco3ZyRc6FSecgVik28hW0d9yGWddeHDyhEe3vVs4FGN4ALL
F2kRaTOEEWBjwccvBRaI1y1CNxBy6tehJbEfOrlisneQAn6aN2oEmv+gWsCQ
x/HVdEGtDztCnGI+F2sHecVndcUf9dW3kpv1hEi2Hl6LuIEAKO92OllpFxg+
W0QVR6ncGIhSEDrNEG9p3oQOxsnFs7CFIbaWcsoY6bPpA3g0YwW7OV5vhYOB
gTjzgzRHoovt3rEPuwiEaxpYTlVQJ2Lo8egjk5JzZuY4VeH79oZsZ0+46jzk
lXu9sxDTUvKwouhR1e8E3cZKkpRlfj2pTzc++ljLQ+Ps4jJPCLMuodRERyNQ
LAQMy2AgEebuO28u3F1h7+YUGQiZuOeN0aS7NwtfQnP+/pQHZmN4bWsu4nKa
a0Mj5r/1UqYD/wofrJprHnWDXfIRUQMmdt63BgBdAd7nF6OdiQEXZ3WpGA2X
dkHYJCdP7h+5JC0E3gd3mRTC89FDcgiqiwFqqR9ROR0e7mxdgNXzBm++mToF
Gu8002ZK/Xp9jYT37XqxvxJ1NK49k2ea/x0NjCkyyiHUkvP0FueeJwiIszVc
PpZJh4CdGW1W74fHcHY0DVLn9SelFJrH9nZYSFGGYQ39hYvu4wnQ3fGRAqeK
TVUbjU5dVgWMNtaxPQZckwKOA7agGSOkxBPcISTIuag7Yr5DerfPuzs8uP/9
ppl8UCe9vkRGqx7st+ZH32BWMEmpgqaYQjz0m9y8m3kzFCL/wZIbvqd9P2ok
6Tkz3OLwWniaMA/rtjIcMyeckMEkpZQ5v9rVpYzGaUmhgSht0F3w4oQq9A6j
S3yHCrgpq9M0Ll+vopYafr+JUiIeq9uwwQLmj9Y3Pj6gjIGf/4jzwIsBhuk0
H2blsRNGsl29RLmj+rQEbpTGgqf2phLbmf9OvIAgPvgBzVXU8Fc4ygByssGB
asPNfD3dduhkZS9FkmN5FjZffwej5EBvkjX84vEbOGV0fO4vQcHHgC75UyOZ
DX3zLzYPVk7ykhK/hzUlMTCys+63NuBLXF/rlBY5ouo+FXkpu4u+4zcP7pxT
B9duRHB/HY/+aFiuyH2Uo4h5WuKl4kx/qKhU3mTkHhdZ8T5yWFc10vCmbYuK
EY/uKrkmTBMRDJYABOnyyTfnJa49u3Es1vxWyINJTviux2aewEaC6rOQWZDn
li++GKXNZjOv6LXdDkt8ZOXVW1s7HSMUffrjZpvqefESnvdnGp95SxSIQuTx
iLoSZM1C5rlsqSERg+nKyRbYkDg/r+SqjkY2pSExxE+nhLTssaDhZAevS1zj
YCD5Ft1GMmJmy1mo/OLWeE9b/069+pgCyQsrpjiwCDtC8oUoo1PSTUJ7EA6g
tkTI78pYQJZqaySaLh1lkYO8EGK3p/VPfm0E3t7T9TEbdMqHDEzJXD7KJLmJ
LEet/+YRKg1jIH2cFErs9KkdJNoCYjx3M5Sbn1QEPKMP+RbQ4roLO1P2Ng0n
51r4Z2KUyhsrJXWsWZvO22Z9+1u+RHdeTJzwEKVGXJVjjdoF52Abf9H+MPd9
vawnhWiaufzmoy4DFo0IWtA+4YG72pMuHfM7o9RtiCJWawfys4Da5EA4bqRb
QAtjsPkYbVuk+viwa3lFONqRjR4naJAG/mIy46KuBXUKle1XG2H1Lr8ER7VE
wMscU1hHrMu+jr8Zbi6Gkuw88GAmgyVE+Qr++aUsWUlfy1nKMJhrO8Eo7zEz
IzUlY1BgT6r15SoMQUONQzvFUj24WLT3EZQsoE5GK5PXNbMIhysv1H9nIslx
QZLeSoxkrt2CcWZfwi7+/1AZBPTHGSfBOVWRbGqf71UohwhUHtW12VSevNOD
X5SGKwyLcFYR9MmFFlWRn2WEfoFx6hJ1amUGo3OoW0m3RQMBW2ifT7x85g8Z
OowC9MtBMsHOzMJz86a+e4Eo7mFs+J0ToEEbUS/IRuoSN/b0WRhy5r+UqNKc
eilFGpJ7yNyvbRrUsKlaq6wm4vGRIfxghCyqJuIzIbjK71YzBOULu5+KY9bv
Q1Ryrj93hBHcRjUyht8vozsJvTpm7Y2m6/WGWWxeK7ZMsK1XrDid5XHpG7DF
f6N3u31iEDGjZciZXLtbSuQCFhi+LqXO+qBHJtTb9oin3UIlmi9J4N4h6Etq
SFCe2pTjQncxrFIxK0IcZOCbCrZmIY9BDuW/KaJ2svqjH4a9Lc2xrkZ1giXT
4/4W2hgKuEo1dvFZnFFdnLbRCCxv/TCM4hsr5vAN2rjk5GX8AJ3gWWuM9u2L
kdq5Efgi0MGtHozoxOpSKBQDDDbP7A0+kg93Be0zyATT3g51zWCl+QPFGR7H
jGYdjkUGH1Mnvsag5ZizHQwe4GNpFWp6n1qB2LTMuI+ylUgQFgi74E50AeMr
Mu2M//hWz61bjteYTLU5XibNuDChBaAFN2H12T01QUhaIkJvMiOtIXnpt0sM
i3k5EfItwD9/g2devH3ZgvkVAh1EewhdeSRSEh1i0XZXMog2yMRZmE8RNGPw
vzOOd5JV1jR3cM2/kU10EdVs2YHqRMlfuUw9stZm2b15LJPD9QRgl/lU+Hdv
NW9E8ym6WN9d/zrdzReZGC8fKHFPcN+EfOFg4pRpYCFfXEMUbAUFp1Vw/CKu
c7xTzoNuNZ5N/1LfbwLKaPq6h/hz1LZxSHjOcSjQPApYO/3N8h8Y0KNzyAyQ
j4MIn9J2lW90BoiAj2wg3GLpoBZ5tkkRWu/tTd/LYdOeQ0uQLbrWr0yK9P4y
JeS/jg2RqThM4i16mVNWnJ8VF4o7tJ7KarsGxBdWlxkIKLtPBW/3A0kpTZP+
K6AtFDWUKM0Uk9frUxiKuqnQQs8ieuXB5g7OM1eSCPMQZQlur5gF94PjCt2+
FcJAX3AKe3Jn2Q29Pj3CyVToqFP2OscPIgMhqXJJZnBU/u5mdELyldR+n0Ye
PxykZIM60P/Lr6XInwD0lYjbJKkTJCK+/0FoNC7MixI9Wu9mpByPAvyUT+V7
JCIPz4fRZbU8ynAjSn70EM9wg84TarHQDb66iFa35j/5D6x9splg3939Z3sq
hCd7Al3lWOluerqfnw7XeyQGa6xi9yFFETzMa4moWUA739LZ1bvah8tLC+5w
QymQrRJA5YtCDDp4stxwWbGlIZz5FWXu4peCpm/o61Mv3vVPHl+vlzwZvEIA
XT9i/+hBDYGi7j/d2dpSh0zJRCTUBMdx9MjApZ5uqkM72kcjmBTNQJEBAb3C
cVkmM5YpojKvZ/EM/CVX1xuWRH1UTRkRzbcPxZRJlIX43dxbhfUAcqkk5pws
E/WdsUCh59O40QqEE8/bzR3+hphVtL9d4W/hQoS0xSC9aW5oiD+ZhwphxxLs
xsvLGOQvWlvqmyGv6dzNhazdx+nObksK1kGq1VH9S2HebtANwBG1IOYVYrAl
nsIR6pYti9E88vN9IMjvNAdIhQut1QS/if8QHak9vhuG+f1D295+lX2F5RZz
7WGIYLiYj9v3o4AHHRDxt5zOV/8awPV8v87oPvVR4kUk1yiepBH8yMrUWmsK
IQoyHvURKinFhy2sV0uVDLeilwslDMmEH4mOBW63Ftwh0osQjZH0gwb19d1y
kOHvBAnm5zPx/OiXtsqj0Te8sxp7nDg/ttQz6TLqoqsleOwNB3n/R79WDxJC
mtnkvRs4aQbt2GPjLC16jOQAvM2rILna1skFZCPVowDIGRjL1doU3DsTADiU
rcerDpA4ZFLjKb+G/v37tyCDzkpvXA7hHq33Xp5M/Dx5Ulmu5xfqutE3DnJA
ysGiSUF1ixgvE46DyMIewIJt0s1J9EfdU+viifme0y2etF2AY2Ex1EJtbXen
SWmPApw63R3HVi1mLOmoHJc/IHQ7y/U+sAu/N0Rx6/qHU+HPSpU7vHzTTMEu
HML+hclHx1VnZZzq2A6ywBJnceWmkQbOE2w2Hnf1tpC51I/9ZAD3teUlnCuS
GCsz8AJJXPRPcoPu/qjYoFhZHuzBkGASf7AHWeOjuVKm4oWaW2Mymj/oj9fq
kIxxiu63s1Uc+dGW1BYyF6fxEwt0DsPa2L4x2MTHaNHLRI+ftZFq5bXL2xOU
aLgn/W29RtSyMZDfUwVzQIdotvH7VFPoViWP5XQo97SM2IGxWXjHBbhiuHPv
yekwiTcBwRug1VkMl93aXdBCPGCgg2ACS3LZ/NETbJ2x9wHJbXHwQjn/A3uw
u4HVFk9GE/ILz6TJL7SdefNUg7J52lnITuxWODGJ//8in/2fN8xgirbluWGM
tgEAmYFQJduHqiUxZw4NvWz3dV+ZPNqGwaz+pu8eXMOW7OiiSpKxjX865H9k
bay8WBt9YIh4KZR8ovpB4Nv3dZgtYlBLvpc09Re3OsjVo8kmiL4B8FMtwCp8
futytZWFbP08tktlLibtNMDgJ0kbqmqNMMprpDCorjxofMCXkH9Z1w+YNIog
wsZqIghiBsMtmgWZYQqChC+eKN9+l1tedfeYyhCv8rcLL7ITx9sB7MZZNyod
3RSjKPm5srImZOXf0M2H9rk00ZiS81ndeg9TOrjEaVVoKKnF0Jh2f+LqkAaq
FicB9QAp8ek+YTsXchT+uNUJSl66x40Y39E9hO/jij5TIMdkKssmPmBgOESM
Lh2giH3JcnE9Ye9yzZM0X7yqKP1BeiKXhA5++NLCbyGQ51+N/pQ0zVq27Kmk
y1DEpV4Boyd9nP34Pvj7kVBLSy3Wm20dqQp6pPH53pRmgOZiry7AhBNFHZxT
2s2HmT32wZhdXKH7xtQzZH3+PruULX+ENm4FIKUMheSbJyQC7dydVsnfMT5e
s1QhkJp87ioFW0DFyH0W0fBKwB5pb5V3srOU2/+Uk4sJsboxGPO0hvp8uRCD
krrJjICyedThK+Zq5kADzAHD+U1iZJUpJlCpJHoq+mnOksc3w5TftfcUvIkb
zBQpzTxEKXk0AlSF7uIWXGSxpjwHyD/VGq609ZXmrhIfHwpFlBb2mDOVjEA1
Yok0aE9GIXgiLlH2J7EI9Ljm26NwY5o6ArIcAlESnmDfKtLX8chbUNeEgVTu
X8aRyL2r4WGkVCQY/jDDhV5V4yFTXKZG7Ky4KPTRLjDXfdK4aSwALbORjQkk
FUlZ9249TVSghTH4AuSFeF1nL6yO4pwv6tXalttB8XYyVAsRjz/ziSWw+zCG
obTOTA7cTkQGHC1/Qz4FLQGyo63WGmk3+acEyeqpgTH6dhUv1Z9JoRfxUHmV
R4X1E+tos+32mhhpjoHfu55hIMF5xiYXWv4/zvyBLQWicSQg5seQf3725Bjh
7kJwFYXayy9zdYRtnliMTl7/J1hKqB/hX5MrnpZ9rygsNofIH42kcBdqA9lt
EooRN5+uBX92q2pElnPCnh2XMDH2j8pVQzXNmAqvFXWrFPmJKQjNssBa9t3b
jse4zsO8dMMknNva0YIjpDgfcRk0byGNUgYDIMZ2eNy/0lf1CjlyArRmMats
3HadspSwmDmh37XpTBEIcEj4wYanMatNgj65rMO9ZAY7W1Vkzg9gKfcJU0XM
O1f8NkFuOiUEAyBR9VSzw9PsoAdaJYmxee/t6IZKiQck8tmeg0/gA9F451V4
OBfXhXjeHIbvVHIu+jnq/NmUkAjMuTRPcnPAT1UIihSyJU2yoO5vP/4hKeub
OkAdsb64z6LkJFPAE0pyf9/z/zzfwjDnFZX9ibC5EjK1JRhDUVgCcO9ssgyr
RUN5C0Mp91vRtLZ/0W8WYF1mMgG9I3vslbaLqvu7FNGSRwnVea+lR4KB5zxP
EcujuOuVLN64QJ2k/1fedvOJDI3p0gJ/6Zdl3/D4MJYY1B6Q+kODG8XixKr/
Ogykv8FbnyLZmG2VbvA2mXv/ntOq3nRu00ETNXZ0WA8s5d2vNthxii4S9hSA
LSE/WYyxzzGORjK0I6n8/TGENaQuApIHG4ct+feCjRDtsXKXTJPZ6jVs/x6F
N6yGr7WEy96mV9UI4G1xFKmXln7jNopwJMVGvu88nwKTfwzfyhkdxQj0x8l9
ZqPC9m0bLr0vZxXnPbDdadYEOinHkVmS+5poZUpcjlLY6oeKTfWdoNRrt/Dl
xTeeC2iqpO1zjtGjs7A4eXgRrj4QLo4iJnJ0Z6qbPASogoE1L/Zo9OhLILoV
QA9ZweXWIRAi+I4NrZFjdlF+qeH7lRzqYPQ7zjl+4qd+d4RvktpGQ1oGnMMd
BwhXspjVVhQ9HNwd5nFbdODrAbYwQIWbuLpbMHRDxcZ/m8Qi0IU491Bs6N3r
+bWu/xJeUWu8Pwpd+8I01775+zo/5PnaYPWnz2CbW0IOiJinDOOYKEIu+IIV
CQqGDuLFbXZnmQkcZXv+X4P6dzxlwByY02KfABJR2cqgssLaQhfiedNOQ7iZ
SD3PFYFw0PkP29IPA/rtdlKO3RXKKDNinDOvqTrRSs3Xnly5rO9AC9AY48LZ
OddJoZ59LPk+qhw1Q6Ct/ukFTZXHkfqIXfBYXjAeJ5MEzqLa5IY8DWnmVcOH
rFEeLtZs5/dnp2AAEyd65iOI7UX9vw78XswrZ/1LLdGFFCJTvbpAeQnryW9f
pZ6zwQ9z2+5mSePn6dL5wLaU9aqF1FddE5ZZjM6/P2DsZ7PkoLHlH1VEdWBM
S0hYeqPQ6pMdbO65e1TuHYPFLp9bqNqZq3ILho+Vxbt5exRPDpB1pVm7eEqn
hqbMTRvRoKdHwDyS6n5FJ5rT2hXawl9wk5eyFG9+70kO2fXfZCHJgFYPVAqJ
dA6thqxOj3gZ5k+3TI7vJXhJZ0ecvxnIaC+YlRATP1+RUhfV6fjlk7IFIcHu
D645uSF/oURD9Ba2Jnkq78Ote4BVGIjE9YdBZ7vr6OBeaz6YU5C4OZK0VslI
elJkyiw4ZbnNIcZrqQOpFH77QMb1KI/x8B7ZQBWznzF7UmylIvWQLp6ehjxx
s+fi3x8d6Sc/TP65YIs6FtuYv+FHeTVHQup5PYNft9zt/5YRgR/cPgOqyseC
vqpENeEMposUcokvu3GjDzXrh5iu2ajrONpT7tTyrqK11xyptLK/7CZ6ZjSD
t9HgGIQeMTsTOOHstsLjXX+PZrIU9aETyOOfLke3PuaTU3RwFD2HrnJJOQjC
IwfIuims81pZoKVKrGMtLJdPyQV1jAfXEot9KGs4FiX8UqU/Ea88PbUumxsc
GCqATVcOHbcXhrR4E3Dmaf1XocGg+bCWNPR7vn/YuYxqwG3b8b30+3uYQwqh
g2HYMkSD8cKO0pCUAiokS4MAivxBLLV6Jw91kzCaGiWsS/YPXOmrd6CmWWJK
/tlQ2O3tyns+p309dBVIa1MaY0WMuv4brIfysb0SDHpyhpMsIgBnfXEfLYSh
sdl0Yq4Zl9Z1IkWbfpdoRTAijxp93a24Zf+hGPLV54Ptn3EKOtq2yTIjB0jj
bSPnAnjZ+vRDXFsEpC/nPvRllb9Eq9pDdcyCV9yfMsUqfsFRQDKSN4QENBQF
aXJkUb845xB3AJwue+cn/azx5A8KTzKw8/8EUOdoux5HXb1OXVPU6EjdfL17
DO3g/EEhzdZlRoIltZgRGZyAJB442Q61s5Y4Qjd7sqRX9euTROETWHwBBq+i
EC6SyqCXuevyBrSC9XxnxmfyKV5i5qiQOaRiXRMERAKnKPpLO3qiMW8ritCl
aiVCA1D8V1M1BLa12aUlUfr2Q6Ab1ee2Bkvf3HoPesZJBTe2kfggUlFcxTWA
yERxbbbdvtJO0i8+ogxeMTBHa8utLpbuNViXt5gE+6ouoZDcrD8Aif61wqoi
uuY71zoiCy0ANKYT7198qVFIHyD/YNZ8iuedythYLcrW4rmTtoiEdgkt2qW+
LXnsOFLItJSU2czL6rxBlqilYwgYYTOD2Pan9PPKDyb4tTBf6jfXjBHKWiYk
NpC5+xH7HmIYQwM6AKCOq4uWA8NrqRoYG3PRh0sOM1Xb02HCqYn6bcKS73pM
YS/MP7Vr9l3+nx+IJCEHHp5zTz6KAurh3DGLnJmX8gnY7t7zi1SkdOWTWtqL
lWYUaVVVeZiszH4B20OgmWhkSLB8dKqDS0QIeOWsVSv+eU9SOtzkZjS5mGXa
avr7uPm9mRQ1Fp+uet6SJIXyWrjKEN53C7JxKURdQ0NLKHa33pgpkxt2gU55
houy3a52a2vgvBIVGeMfCRgYlGivdyFinBYIAOQu5CnZJ5lh3O7bvqXwOdku
ResEK3cSlqWyZH3kVUo8+p6zjAPRW0jirVaRMrTC7/DEys96rinzCz/MSIFg
SQyuZFP1GzKZLrI6+uwQBDESGB0V44SyDdkSKvMD3bwYgmuxAA3qBJ4OReZv
bInDgcxcKi5v9qCWoLRE63gOGxGT3wZpgCGKyeO38wfnUUsyWcvXi4uTlXBC
omhZA+FnWQ7X22QdWkDvEkvAEShCFWzU8Rp98HO0rrlMtqxAWTUiAZGx0UGu
wgRGnP8/2qISuHuRH6/NbvxW2w/NClAAaeg3XaptF2nvsh0ufFVvKQpT5A+o
gH9fvz8Pv+83CinH9rFqWD0c9BYfoe33+w3WqOcTwnyZPZHOp/NULqwJx99X
lXTlLiAsAIDwYWgbYAyJvvTnhLGmE2N0RiydiMaOyEbtJy/6dWNDMKcHGB8V
YzW5z3Ozq/UAKtE/6xrVQ8EYLSAbjtXeSdadOM3f/TSvD1sHbAqTIuH9tivR
+vqdecKGXRNv2vRp+8AOc059Q7cmgWKDE1gksSimRSEflkHsPjZbd74bDTWS
Jd0vB7u+leUnKXGQa7zWDs0spr7boXcINXn7ZUa8izOpSvm6JHOWlJkE/Mhx
tMccxsvEwM7NiIwbmdNIlVyBQRk0PzVdrjtCcID5YCxcj/AHEtpd3kKgQS/k
vEn5wXPu4YkzgZM5el36Do9d+JU0yrhZYLp0OFSAwmDmy48QKgNPBfnoltAd
5bTdkRKMZn3UCzEH6K6z8+CXz/z0XovFww6M/QK+AO92lXLbKsiHZOpQp1pN
6rSj0Mszm/hsUqS4WKu8Ly9J1JIoqADpEqA90kvcmZ0fmd6bXWe9wHRueINf
9JUFpDjVg5ow4byWa95BTPozFwm5zf5JwVKZHtk1Kjpx+D2BJrkBsOjXszjY
chsm1w1WimjmY5jJivdQ0oPDcISgY4aiU5OKtaTFxXor1Cpgk3XXgWczFYLU
3ZN+jthiFkb8tEHf4T8Y8nT2HHO4wSds1xo1ut4DVKqk7aMhtKYJKALgrcam
rMyBjcloJkG4geHGINw0O49RTNEfI1g2wy3v9rllns5mYamabX1M8tqnvx20
6Ck5pBEpM51LVu+TtnshEGVn0X/YoljGyQkN3IzYEYxS6IIUdoKa1Buz/XJJ
/CmMjkMCB3VdUDl39RAFrmQaXF9/v48XLcoRZikqjbNucjsxmnvoZEffdn/F
Kuid5NquUe+ftK+mf3xjo/6RZKllmteYg4B/yfTEJIcHDLKnDkVmTqnj3sxq
JNyZcpWwDC/Nfw2o7skMLGhmtApvceABaDaG5A6Om87vYO1/QTyGUj0z7PYf
YDOhJI/NPG47+vYQDT4YHZkJMKSoNuiT0DYyDXOknEqPu0vrbxZgCIFh0lZ7
7LC/1QNO+yEvzdBmoyvCH2uM+ljLBPn1vzxDNjQtS27eUVtH3e7Lo1KyqfNb
NBNRVzBS8CwRWZcpMwLYFUJn7GuNbWcYpLTlu2fPEqzqpvvCNN+j8KwStdfj
iSgSvucC2BhRbNiiEzceOowc51ryyfRMsorNZk90nqJMm420jbVQG4jLX6Jn
6JOKb7XT8B4AqCozSrpjY2T9mv0fxVA+VFRvheg8OMwxJKQ3NckptTXToc3D
vnc9WiuMLu329PwVRjUjWNa+rXq5Z1bEzsJyDKEtY5flYKccvrmSaAEylsf9
AhJN1nPh6i8du6ZM0xIghNzXpcapgw++8zZ7/LjI11XzL71oTPHAsPP9C7cQ
kEqlg6kILb2akzrtz9TF8cJ4EaacCAprnX1Z28fQw9mOhaoc8/x05gUIfFWg
n2GnM//qh4nqpEWw1pd/Ebwk5+WuhO/vyJFbHj7oeBgeNEXeTWFmvVNeqbCT
KqWuPjWy4TSr/ULzeJME2E1jYjL30Gc3jGiUSyg7574W+WwzHMuCmZDjxkHR
ngAd9gSh5mmWY8eHdPjWAr0pBgzpRDlQ6wpPj2QKTOF5FGTkVy9i82f8NfvM
2U9ZA0lJSL7RwtTet1rsEOsRuk+AJSmwvFuK4VMJLiNlbppQi/3eMPRKJumT
t7YAkFvBx/gXKCMMtiqfxq4rPrP/KfO63qfFY9MNHeTDtFs1prKEH6VCkMgS
wEGcbM8I1VfxYPuSBsgWv6uwIvovc633leLdYVMQyuIh5rkkTHrgyDklnXme
fZ+YJsQaki1wJync2a8Xt16Skxi7cHFkYHSEnU6lBJp1W1LoVFhGLppqjLnd
FLtNiCM4D/Mrbxbj9QVRfoGhkighirp1jkdCm1tdjB3yVEdREPd42uWPBuc7
XTwFm+Cj0/fsYTR9lrmPYPBBpgZs2A+WWFJFyQ9hgRHOn8XKbaUt3OHGqiot
zzgH9dkHYGyurioM2et9bMazAvTM2L8TvF1sx1t6cDVpN66LAXZmSLyQZ7V4
FXD2YReaUmAVv+v+AZmZZhyUUPXe67adaIarmdJXFa7gwFQTW5Czp2rSUPI9
9InHSJOafnT2HeVM8HuI1y9thnD4+I0DUouINtyMsQEDLftTH+w/IV9DUItE
7EsRDp5HyEqdAHFNwWEa4aMbApTINkWeRAHctYWNb3QS3QPo7E0AQz0DhFlJ
K7043Z0uvWKQjNnB8sGVEnPKUeY3HDKNif9TtYEbQ6Ji9FqHEOT6pUT7YpkC
8UYwTw/Pc/uT87+jyp8WbEK3nFaZ33FoZyCgOzUYH1vrtBChQajr4SlZuIKb
jLlSB/4UBWDeeXMWP027Dv3bYbKn3GpQdVJYQj7YmpTSmfgBJTyoEAQRE/dn
c4YhbQbGlyxRmqwBC8jIpczcz0qFdjmdllKtcFEB//g5d6myQPYEA+53YzQs
1iA4k3ljehYPMJEhfl3j1T3yzL82uw0mzNiXErkIj+EGC/XjF7CuBYF/Nj+M
Ikyi+nHks8d+ZWgT8djJeewzegVAUv6z9DSlyzYA9mex+gTvghlakV4TDz9C
9AixbpnxuVcObkc05sidm50X7gSKbDvJb3xqajiIwuzXP2MXNYrt62xxJ2Oy
JcxHa5JOHk1Ig8deoSZdP+Ugk4dGZpD9X+OzWM3t5t7USAXiMEyl6u6Rf68u
mdUACKtX6QxQFzgcS93Zc3KDNOYU1OzYDN9uABx4HcjzEpKOXTjHfYbwgOcT
E+RoX6J7KRXU3Dsd25QagfvSX84/XyxCp64QPhtqN14A/GbWHkLo0SGIDr8V
zBqkpW7utgRl/SPJ/0RQSexNunoXHLLkQAEHHmB1Nq6uf6bh1grB+Wq+R401
CMbpCtFaA+5oWHVtAP2Y4rQwRgVyhgyiEPOXDTTUvFB757zB6Or9UpFmKMxH
eCJ1JJZA1BJ7PES0ZVg2HvD2rcxhWaZeP2qbNoF4g03FoZK6qAnuCp7vouYc
vjD0p1IfqGCs99qdlnewukdfxkYhblt7tMyf3dqfhZ+YmM4UWHByKrl32ErJ
6AwplsQFL4xOZ1PZ/VM7DJB2eWo1mdrEiVra/0kvWIeb7bgSEoTsZHv9ExJE
yJ8pILZecjhQFxR6fWw2X5Q1hT0BvRdBo7uUFWElcexe/D5qXRyC/Wr0Is9C
WXGxH7B8OMzo/AlJwHclSLVDSAIag4OnHcJzuzBxVC65BRpwYiXKIxTSPvbE
9hPu2A/MUIgl9nSBP0T37uWMgzqZpNpHpo/EH0qUhO9mW098i79O3NzHm7R6
d19I/8tkGD5rf+KIN4zgSxq5bKNg5blpFWJWBXOkkSJVuCVBSecNJue52Qvo
zJqZR5nb7EZk6h3foL+G0Xp0oiz1Sb56JN+FMsZgdkgqgbBFQCPs2Kd8qx4W
rIlvkML/f+IkHbjTCfkcWBouF0DEZ4k4bVwFwagnC+U3ec5ZVxKlDVUKluUk
31uwlxsSbTRN0bY8DcJ73IMzllvy9uKUaKyR2RHUbeaFmfSdEAyyJFCbuY2y
HoEqFauQuY+OSeViNXO+JpJJaImd5GiDHwcbbFqf58Pc8itzOnUbnqKKRk8e
kyyV/lAdgPKc7hUekdZWoo0DaAZ7ViEkeOgUhS9I+nBUgOOQdLqyU6++4Sv3
tV7lejE1c0CoIdXLUPbO5ox0Ad0DTlwDEzATV57QQ7MpqgcHh13oBTmJIJ1V
DopRNVdfbg70M3WFW9+MlAPrU7v9RtQsnOJ2AeNppVDbNGtbmLfFLRJTKWbT
IfOc7u8NjJoGjF+ktb2mKr4TniT4CvrwW5F8114rjfnftmtnlCLlwILIzzKl
fIa9ho5fuFGDXTkXByVilFj+HPG9ARchGIkRhdp3Hk6BG/u+Cuwo3/egUCJH
LLLdPJ+0Q0BontZ1+25162QEgV6vrEIQtofcDXaKiI+zQc/RqQLT8JsUWHZK
OvepsHCgauenWC/VspGKvwbbPyAUitGMZxGBdgh5wxljxO+JElyAP9PmTq9b
3W+asnYBEkfM78J7+hhEimsvn21OQgPze7XZx4h7xEN+tWlyv6PXIkEDH5eG
vFlGolsj9i/6fw4NSYqHIuIjYBOV8jps3FgMqtAUezcSJgUZkS7fVqOUaxW1
cpAIRpAoireVEOgRrJUTMHIGkBJe1x/ffY/fht08oRi0lD8gCfn+dO/e+WXP
8T150ldkQKbieixnaVf1r3HAj8KfPzZ95Fdt1KIiIrIqaX/SpFuHYv/p7+/V
BvxOZSuDsQYpLq4Crwhjux9YyGuqmjOkg8ztdI4/pLbe0CMiAHMQ3YVbV/aF
NaZNXtC/Mqb0UQYHR4xOpHm1NGh3xpkP1N/RQveT1HdWvW0/NYilmWw0VWZs
So3Th4qW9WjZzhGYbxv/VoDMdZ9c5ZmCuFLTSwJFMdle6+DXuwl8VAcpD267
A4reHmxdn/8hAvpJ9sYp2kXeZRe0HSgdFWWgCfm+QVxB5I4Ju/DtSJgi/cVD
z96X2EXep3/qNrcGW2cl8+hlymmAXbIWwzYqJxf/SDi4cyHArWbR0FyQ4Xl+
3RfHeO/7ehGV+6t6W3mbxGrxgVkgkTx15P729F3Mosao/yoG/Qa00A6bpoJc
WE3nj1zoS3Mg+RJm83D3o0hj4eJCjYQyzs4BUndTb9k6onbdEYqjo3/EY2zU
gwJG+rkvDq/YVxMP/d1mvw8TiFN1KfrvDl6cbeQR0GvgUWvyRQYVYuGUTE//
rau8Il5AV6ztJ1Zt9RxKt0XSiOMRNQVwZp8Lgnb0AX8ODKTzy1IsAGBePjey
eCAgBQKv1GwiQUahUSKVcoCluumB1ACBb533FDOJUrVpGUZkAPqtrqJjBbMr
mOYB9fRZiTPhJKXu+Lq9l6kmvoURW2i0H0gK0AtvRl522tJE/FJxFZDQrz/g
Fiei9Q0gr5JDnLIwKFLpY3xVT0FoaDku6ISDhzCAMpBhpks7abwyXx4VbCk0
A1y8J3Ca6RICYVCLABgwBrKO6t3/8qZKE2kKQuYvLd+QnJPqiehpFXiqIOAi
omUUYRI6HWboKlLYIRbOYiqnrdX3SoW350LRw+gLcdTUHu8FKQGVA232KkFe
+Ol/jhQELod7R22qD3qm36ZWYC0ChrVvBD6rHRQYxC+Dg63Hf88tnuTMnayK
Udgbq3HSrzKL9FCDI5ehCM3g/CRW5SPKZlSWWsmU41K3EWH9I5eTnQOt0XM5
GT/JMDN0Prv9Nheh3zVFCof3DK6EF3Csq4blg6lPqr6FN3CkozSUvB/hrz8W
8J9LZJZCwGo0vr7ISeUe5+VDAb1JMfid8Rvc5rNnCYEVGLfXaLYQVTMyfyRH
68TH2aXCDcMVBaF/5MnMz2jJGlVF7G2kw+svSCqLvoWOSUtG31CuZvtyjWYm
sw6NmzN7ovd2QK1K6BZ9ot1gCb+xLLmpJiTqbWsfUpM06rdLdIrF/JgUBhUS
uiV79CTz5QqcifsEJwcZ2b1zJ2QMrVme9BHyHcC8HOwuK/NDi+4bYII9pt/r
ZOAUan2Scr0lzhc3yPVyn9cBiprLguHcJKst0ujubYRdwYh/OTZxXHLjD5lF
+plbXAeyTNKJrQcIM2or+xnRHhLAT92EzSB2SZZ7qWZmJzax6UWQEfczqHaD
YwcpY7ECGAA0zTD5uAhBxzd6a+9cKXvIG6F0RVAfO/RCj+/1fncoGD0dgs4D
5UW3WfLtfBp3dnoVzJzIHjoeKkjt1q00LPaeFPE7vY4ExFOPQiQgjRLzoSKJ
BqqDxrDi+uGks0LgxF+V6zU6dt/dqlIA8WrQNJgYfCez4D0G9+2D6EODqs5K
gsC7Iqj7F6AYsUoAJjbGlDzLsVMG0VtE6k2exOQRgzFe1vdqohqfg5c2dwaj
f0zwy/PX1gP+We90r9RT4zP2FS/AA/CaNZwPg/J0YRtrNvEYi1VJ9BaLAjn2
jgDUVUrj/x+Y6jCh1Ptdsi8ILirh2DlSrum29RZaXRGNTKrvb+tNK1JeS3Pr
IWTurlsnD5jPo8D3DTr52t80P9psvlLkf2MMvFsiNeh4GTjHUlqVBmjkUCKy
8kVP2JNFwwEiO1GRq3ftYkVtR21RLlPJqfOXHXA3014KG5acDIDZ8cfyTSop
NO/SPN/rjHiBpo/RTsM9cuKZdOOB2sLGX8SBaMLQriQRJVReh3ZXTfgc01bJ
5zO4oDdWGiwxjMYYUKh7NoPwLWn/wz4bc5rJGFXOFpR6m/WYzqw0Y1iCZY5V
S7z359a7mUTdkMF7jYGFyeQqGQKOr0gKMl8rTAu/J2k6HQUghVe/Tsj93XqK
7n/mN9VI7YVXEp6/ovibm7jubfmmnNJUoziMEp69gKa6WsOYqpP1uxe65Xxy
wGhOcnVQ02y+UmYBv26wcPMgSK7BurPEEI85R98oWGEshGbzqJw3w73L/ojA
MZr3Aghvq92N/5mp9vWHVKXXcm6GmOgbJCCvQ/B00cuUFDt1MF55+SzH2hpN
jtUosqA0lKupsWct8GlNaUFrc8OcyXYT4J6QWDUX1U9RnLQRIRWlzCGsIeFs
WkxKClIuCabnzxwjTVRUadrnyQdkxAUqgZb8tbHN/SGAl2T/dNY0VwnuL1Gr
tA76PUSSrbyl+kz1XMu/UGHQAnGDbjZBN4suBLF8aj4UZhyM9Tk31cM7RVq0
/HFuKHmqKVSrS7rig0jQWYMRw0OZPZWKk4MsPr67tUyBobxL4TEvSf2e95O7
bNQRqIzYRyChOT/KKBdpx293EaxskUrXo99eC+ovQTnmIGwESJ6mIce6K5bb
F1NDNBuYv0pWKHRyq5s8ZizX9XS15rpKnWWK0n/XiePT//gnBT9ygUOQR2c+
wepT/BpLrZcJ9L1qNi0G/hGm83ryavlGr5X+6k1lpGbwjQ0xImOjWao3DS1W
2BYVrYvGHk7yM1qcunlXPtiIi9ZdLJSIMOuWLfLWjXeio02HVNW8Iy3KJGgB
Un43mmR3Qxm36ZP8V6krSoT4wuodOdYe8sOaRCfmQQ4cRZGJORmDa2a+Kw+s
GxyBiSwrI6zMZ8RXWmOwlGA8eMgSX8pDZaz+DApjc5Lso/NmKkC2RGrtVOcA
XdpTLu26UUn/GFmiPWRcf2TRDlUJFK/XapJeDlWUlvq6FBIcb8MxkHbADQP0
AvfV0wyITEjnDMv8HSsbmbk1/yWs7i6uih+ePTTye3lw11YvX9HQRvJV0ITi
XA5XeisPIiAZVVrXkB1DMWsEdLOZkbZw0PLHzG8FSeqBeahT5P0hNGG6QSxQ
/KKpBUJdJKRjenxcg+SIskSbe/ry2gcqJ3cZXekYHrPrNeByw07eHxvV80Dv
zvz8xxj0ljX7hnkgSVesJSsb2hmRi7v6Pdhb8ZvmTFgweo2qAkKjlQjL1p+Q
U9aXzyH6PfO0oNs0mK36X0bEje55QyQhUJ1YYkao6d1G9D3ijiarFlRPKIp9
Ly1qsCXnmiMN/3W36wfVb+FdI1Ae1Q/suvoGTNxATuKbfKjKpoypK/h3YhHj
1RYmmdAlNHkxH5T9pHMGI/kRs1nw8o6FBeF/1JknDHEgMjqATKFCPCljApnd
ySesK+g+cJ1qpHEpVPGoITYamQGhlm26EVEaMnxwd5S3naTjZoi0AKA2hw04
OVC/QLWu1EN4hjGWihs1MBXLu15CvngHxeRMRsaoVXjqOSr0hZwLpmGN03+x
yXs5gLvtPZe1sWE2ALszdXQUZDAZMw+4DO9FEAcH35+y98f7G6KkSzf6XnkN
zYIqhfx+h8tTm3UH6rMk/n6cWLrIjX+HU3Z521VbKA+p46i6Gm8Ux0JGsRSO
SzsTFiRD/Unzbfw+5mbw1vK+D1JZbzKxUDvKNOaLWnF70GdzD+isb82SsVEk
HJPdAZyztZxs1CQGA2JtMKkPGhky1qZoKj4HeCoqYcPHIYTAc9lyiicWTz/N
eYK5IhUmpTvNWC7fBeB17W/yVazsem2eOcOYxQJKfKNJ9lB+UcZuszCPsjK1
zzDd8vsVZxiGMkzRELdUe1BPmVkw7F4fW9d5LnQf3oHQKWonCB77mldQaEtY
3+6YlZreVG/T/t/3ynBioBu498mGmA9FbQrewelMVQH45HfTFhBj8p8eZDv1
RU8XceDbX/tEH5fK+YVVjVdwkenhhdMWaJIfKBYFPPew2poCi52j4hOMmDfB
p362T0Z2NytASR8XlGfyF3po3uoS94ZyU2rPL3Y1S1mMI7j9begACutXx+Cs
tJNHjPAZ0Fwuvi77VXhrdzrpoFRXqArSJAnxKO6BwRMrHX0SLdF78dtuum0U
oxUdH6L/AbQ4G9pcOlTciEpPIyL8mlw3mWUTKP3LzLAhLoxkAWSxqEqqkiaP
vM9XGsDp2PrIxsUtA5VRt/vNII84nDHPx+PrnsURdeiS4jbtXjvcZFgYiK2n
GG/S61RkJFbixCwA+gC4l/7HZcoGsfKodd0LToaVsaq8bQGdgI96BmTXQKkq
ImdDTt32lQodxc18gr+lWjCRYhrDL4K4hAGFUdmC8s4vCu2NB9/RcTz7mmHN
Qx74tN/wCKpy2CgN7/Gb2iDB1EQjdbSWPhZnRi5MOAkI4OQyl93Vf53fFThw
Pw/Qq2DBK++ktz3MzaFENQYLGNUdt44qPFEUMSIjdZ4M0gaVRyv3Tj1nn6eY
zQNmiEWPiXMWcZeWQRuGB/Gq+DVm3ywHLkWcSzZlPxyLcFKNx6heoUp7XoI+
AkRqjSCBxQUe+l7Q3qQab1m72VaTx0nCZwvHM4gqXnXGAOKVVQewaGYBg8oS
FCgSLrUDg23QYo3Me0a7CaLeGH5WzwD3weX+VOt3Fh9tgZPI9Cb9yXhQF0Xm
2CXYmGTE8JW+1DQGFNjdZGhy4v1BMBzAPQ8lc5UVcgOGRqZGjRVRXMUe/sFJ
NazbLokbOM+d6vFVQROTj4CVZzBsqIYD4uUBItKPeRht+iTlAoh3kfL0yPOt
9r0maStTzpC9sJ+M0b2ksZ3VdQvSC9sEIMrUgBDk8XqwBIJ2QyiVJXcz7Us2
Zu22LymvOxqMy0EB2hH1qbrriheeLU0YKwKTcoidIKk/hkg3SMRHndHPvVD8
CagtjTuVyKs/xp6O6kDoOTlQS/V5nTCSi8NDEQG36IpNFIEUiG8zKltov0bw
RSI31ypfwx1ojR7jaRIwbQGLF5qH+SI30aJqqbVeGZaoLJYFRoQkkq8Ww7DO
CvpTqFaJZBissJcS2PBYwO0MB4UiSx+lkvCXv38CHetdMTVIppOeyB6+uYUQ
02FSVhAmt3wFrIi7ZEH5uqltU3bO4Nq97PtCJGSzJnW4yZid0I5oXr+0epxA
8o2EoZMm/D8lbU4EmfLDkIJgX7UrSCTQE4h3SkwsNCleV9vLBorBDn2A5OVj
WGWfnUeehhUvS9zuOUGgLBVmUZPGDYarzfngAVwWhW10AAygnfTdHcm/ZLBq
XpS+OuPIk5DABTv1qoCf42Uhw0EUwRBbL42jRqaFYVbXWFOUAY/uh/nX955R
nJ5DYketag7GDpv7LLC/8T0gKByJSe3O/ReDIj4FG/ypokOk2ISM2pPfMJkp
CnSRdq1ml/zMBwgp8xVlB2+O8mzecEPRbJ24FfqRlfk8BRshLAzzqbLCzfB7
Kuh0gZFfiTrlR/OPR6CFh0IZdqF1vNS3Cdoc6reQRUFFp7nI3TZWczDPenmM
loxSE6TWcnfMWvPGXlRiMJmvJoc6D23SvkjHfOutuAxabJYcMBlY3srdXsUP
Fw0NyF4ZbjEz8P/tikbh+WZ1Gje1rZJL/ROBDCDkU2Khgggj1kCpebxSVXTV
OoIkN9ckcPSyXUgekoWMRZ6Z2Y+8RBTDidqjANUTZFmkx0MiUpDqrz8PZmhN
/zHdyEN728I+KMrJFowG40pgC7mQ1Gu9FKuS5F7NyR9+ODjcTlRkueMItKBZ
p6w571H3WCxtfj6bJYR8iepIRFpZAcMi8u9amkeQaQ8uOZ1yf6Vb/6Go0FiF
YZBYX+VyhAMLb0Axw6iYP5XywFLT4bQ5vv4mvKVmh02l2feJljKO1OXMyNgE
HU/4pWqvoBKzDsxCpmWn3kDP8oJMb84iWIsACRUTgva2AgWhs+UJ1izfynZK
ji4ABcgQFkHL/89fSGQV/G00sEOGP2iTjKBYStoyWgT8Y71DXNfoGgFazp71
0L3PHhEXh8HG5NlWI2Ptl7wkDBHIQ3YGOH+USUafFNf4z8jYJhaIHewysNzh
Bl1ik/RkOe/v+A0ky46NZZehpOoeYmIlHsLBL8Yccfo4QP8KII+ilVIURij2
9VW5CvlT8E7U66/d9/B7tI9rotYM+1/uKdqoWPSPfkKtrM9j8F6+rwkRFZiZ
+SbFVT6WtmGyO51Ccx1HpkU5K4uCT2Xd2HMeOkoXU+qmgCm4EIqP2519+God
svjByV4YhecB8lvWkABs4h7HoL8faKbOYI+COzVsJbULthC7u0T1lixMMc98
g6c8kCr86nHXTmdnT3F/CuTrRQNQgwWIUIcFF+VxzSCkzuCY15M3D6AtmgKX
vJTf6sT9xgrLiLp8O7NGR9QCzRDOJBeT4H56mXskdh+/VHaFOnB3dOjA97UQ
Dq3rF9VVd4ze3a67o1OdxW6HVRsJbrnC9eGyIl7Aw5ylkBAS5K+yMg7TfCJ4
o4AE2DvzrzwLgghHbflJ8MMN/eDBmkrSxy7TyhmkiL1ZJKu+Ys9REkLiHgAr
59cDG/mwbGtzA6xlA0+DjR8RHNVBxGc2H700G8ti1+ax8VPp0uMHzG3sAF0N
6bZwf2GIDcHU45N3lcf6E5vyOHxNHX392tIJZI26PjeCVN45SgyDdQmpSUKx
fyXPg+PrXoEaMfcjo6mStmeT6LOEDJm1JmGoBMAkM4QvmHM8aH4PlEBVRob4
QxGCYKhPpfpsVUOqkTwN1Lmfy2qwZjqt9iFcaBlve9sIY/vtaFweVDR3zjBO
VMxTp9QEoOUmEUnxHLCs/6ItjuymTHoJhgaEvLQSwcCy/EKA9d+dE05EZlcb
n1xngwORtrBio1mrWKr/CYN5U1sO5jryKOyzvuFJY+YFaN4dp+nq+d6Kx2o4
3IxA3xfh2+8KLDf/jv7u8gMEfVI/UfrwS08UIOy7inBTZwkTKFXptp2/m7/F
pjMQFz7yYbOrBkgF2KetVxvTX7A6xi/B1DSUQb3/z5o2gJhFfPoqhBXW+QkJ
kgHAf8hDRwjFcYiK6frz2NOFgCeYLD/xzntOZ7jcZI2a4gq4xJifHDygu0lW
Yh7lE2kp55Jdp97PHE83dcC22TqqxlyUY9uXvHQCN4bewpsp+d2t/lmYrWhe
YHiJrKj3rT3KmrJShgP3a6viAQMwmIjM1MjPxQ2EFVBfoHioKVSM4/RykhqF
aMfPdPWJjXSHSQwO5Pmlixeh4FKZ5xaQyD2Z8c5ZuIh7OWSa61xbabiasuke
FKKN+S46sPFVWsawXgwyHq9jF1A27atHGRczYJNPQ0IrcAC8ctV5ahPe4YAJ
SH7aIFBOFJ6vftggCZXXnxf3EbIAVaXizESicMVPX5PIL3e7qgAPthRWYtpp
JZwKHZvuXdS0u1QepnMes2+nGd5Jpb/359hKWBYxqaRPlQxu/qWdSb3Suoco
5Libw3vYPmekQ+KXvXOY1zLv3VC+i/LliU9Tn7WBTMobcihcQhTS4+G1FlU5
ByNGUzjvKskK4ueQequAw89Jt3QIUWgTqT1l8J/xfPmqCwwdQo5c2ATZXJGn
94DZNgYs9sEUsIO5neZfYxQ1sf/pwmw2g/NMmHETOUo4VF3k/gQKPD8Q4DKd
BdrPAu3+5QwlhuE4lA3LG6/kEf2qIysSJNA8n4D7fgG5oNyvcARzcSkQV/A9
JgSK7ID/dmwzheIxrKCcOx1NmEOcH6/9Rl1tYAN/I8BrVolCkW8WwbFx5uqe
GySc0BAy/rrQPPA1yzkzPDqPKt1YdpPcEWlOAHC0IbiOSiBZfdicsiLG5rny
BODmGbjcsaEtuMNcV6zAhOQJb/e7+PQpZRqo8mHUHzJhulZmPuGz50RBVFV7
Q45tAh9I3jEy7WUijaBlGYB9RRX++p/AWsr8Hbo6edgVqj1QmDcC1A9h7CAW
erumZKKXfew3zhtfOXb0X6F50aE90A6v9T/UwZC04Mj0JQx6esEGYmH3G6s5
Jhb8z0grKhNClYmOoAJnlJpZdqRWEad8WikdaVsYNfuZJpyheQiFuS6WVK2B
6/lyD9pxkez+IBmdAhBWpFV6StIVLnJo8Ibj8/AzLh8SstD+pmsqF+9uG9uF
EXtkoxft75uJm3esdKTC/VSGrI3jpejOPx4nRfSycaajgakgORUEmbrsA9bV
3w3Y6sF8v3xCuug0l4O09P93x/5JHNCZY+n+wgQ5/Hx52s6G+LpB0Hi7w3QD
tbiYAJYK8HOW3bz9W8Gk53CxPD3iZ1SnacpBJ03nuL/e+03wr3s7mWZezE1G
fXum5bmqv3wJ2cdh8evwCEj+GGB953DW/7rx/fk2SWkDpmt5/RdYoHHPe0iv
uq5MxDlYugHwcl2bhNONa2T0xGjTmMf0qD0Jue0FMw2nmAbmmU4hvnouhZ7x
NSC9Svqb/HzGsjfQ7cqRw0WkyO1XnCU7h0Xv2OgSelrdVm34b8C6jjpCxWW2
TKcktfcQ2CpHPb3ygsnD2mJZYjyC9BQOzEwtyNyTYiC4nZTrSvbsSy7k/O2w
H2xRV8OqrkaYFkDn+K7ulm+G52dV6FN+2KLUp8rQGgjvRqSDqCpZzRVKLTSJ
1E0as+LLPs7KHif+ZW8FhinmB1rlq7BnACJkASWpqgUhq942MqizZrD/BUcE
lN+3WBYeTAW/PFvgAKMZqf9zSe6bXTXz6zapdziooOALLDctf65P+l10SRiz
o+nGLsD+dsXeEnJDEC4lDP5t25uklQc5Lea5ZpEHxR2AEGtgxd+lyfutGqPV
tkxSQYiE02Yh/9neArL9CeGPf9eR88IDS+THbvc2nB+HxUgajgfs10insZFa
kzwjVqFLX3QGI5cwrIQ2SzoiFEaZboIE3aCtDdjf7hkNJjbkkBOHK5hIaTKT
mMQFV2EG/y/kcCkvXLoGVYr8WJQZYIHtp7RM57he4nOsPFUL5jXmGWIAfGx4
TewBNmu7kdKbH4o2QgVf9ry6jSfkm4Vca1iiZVSApyrKMybexU1SKaBOI7pa
HjtFMgd1kpnV5uit9FX4TBrh47530yDSdCHuUR1VuXv0FgCN7Y+uaJHvtgUo
D8eOdi5P/IslHhBkZ5VqtfDzpwBMFmb/qX6Fi+B3WVjaNv+3elqii2uPwlb9
0Aj5cw3woo2RC2eDz7X22WToUqeBRtphqVktzdgWZYT6c1HvlHW6yJjsjmQb
GriRUDoNkFHWsFrULnJbkl6JkajDR/GZil/WH9II2bEw7yBJdLQNYgnpcdF3
Q1QFebh8/j//bNqz2DRqrc3dCiZvLzE9RmfsQlVZtHxPsCCkHrjUjW9zb43+
JyfO8SHFRIfGVOnksOIdmQjaAnmXyA1o4dYk5bALsyyviXfZBCaNnh0/Ri8d
ryn7Jaj3M4qo0F3JTJ5R2eW1yJGGfEMf0jTKoSYlV7HwX3RR5Xacm1lBWRvZ
5a3f275ijbOlav8dMHKOPxEUQ2R3GGizADFXcta8KxeDE4XNei4pdDwnaGxi
srVk/qEdlbjU6Lp8I6ieVFW1g3S2CwvgiFaIp016eRFNwjdGswVgLUZWdhRf
G3RmHFOXFzk7jJOeiqrvlDeCd+OzZ7K/DydMYgAUNb883fz4S/B8fRLziHJK
l+E86okGSprMWYkr/zK4/Bv8hS9ulUEPCbqjtnBCO8NVsB4NGE7KPo8rb9uQ
sb3c35M2U2dQuD0Pc9rMuLL0f4IEKc/2FY0EJl46DkKXsKkL2oE/iERdfCVN
hG90zSsihEOIVgYvPFXI8fLfm/W0zlZaQpDiXQrJSbsqmog1FlzeQuCa6mmN
GE3LGSBGOYmiPWn16SXM0IFquQXtg69QHaTfHarFRkWTEnseiFZljhktX+dH
1EzlDI4Mj9+cjL06HGAxO7H6TAqYk2iJv3hyWJsvEkSr3CWM+VCyuN5LaqCp
Bhzrp3LIJy+3E6Zo08pJRu1aUGpa2xmSbnLyWP4PUa7dACy6aPN/mZwFWNXG
KIOJG9tS9JfNLsVwbnef+2goIJ88tT6wUHVlATQ3ri+irwxWlxtmyusLqbgp
f+6qC68UlBeaOwdm5qQAYzvnGQ6Vpul89BqmtBeF59XciIKH6H2HJ6nKaQ1l
8ffnZ3XAN/jnBCs617T1KZlJ1kdtbw8Yvftnv3bdwmtwGGdbck9C4UhdEpUT
nedwq/1i1KrQmjDD3vybXKh13xiXh0nQPBZ8cU+zfOGrph2yp1HGllrfpQSb
1K40G6cmJuWi6YFNxxxbAhjt4uxUGHGwLMi+LeAlCKFbRvcSoGpZWcFtmnMd
7AbnVVZy3GiIErNSlvonj5LvT5GC9HRNUTc9l0ryw7t4+UTL4Bv8czhZMSgn
1CWc4HifWkGENAxKC7+gsvxSyO3eZ0dxNHMEVCLzcdnKUmn9JYxyL88aoF5Y
nqdQK+0UODglG+PxfJXmv8CNgkvDHmqyRmZtUrCwqXKJPCE3p/yfYpQNfUMt
ewWR1sBM1vJTuPmsxr1JL+sEcpSjybq7JSnGnsnLGyLWmGlupdnXAR++vODs
CVz4z3l6eJVLN3nnEtJtkRYG83Do8vl4M544CdigpEjhtccxMHtKqn5Pufa8
h3folbymadD1AeekWZS+jUNHqxS8e319Jx+LUJ+NzWgnZnltmX5GlGnPgWet
JN+a1s1ZB/K/hEgxNbwQaw3t2rKllSJc1QlGfLZB4lyXcgPPDQIAKQLL2du5
kNV452yO1aS4csJK/lBNV3EkQlilJXMhQ1WkfHRoWZA2QBSpe3/N/PhFpAbB
phtcThkvYu7kgjZMQvmemVYYFQDvef4RkvjrvJlZMbp5ivy4p3RXKZ9C2c4v
yQX6bJ2wDeD57WOkOZuNSGZhlTHa5EGvh/9QkX5nrGmXA1kvZ+TSVzdNbl3m
HEQrkcW6LAUZ9DZuaqIucOn/6C+KpIfF7C1wwefVeGMw/ZCJprrolrE0Zla1
/PuYOX8JxoxqIF4xbd+TTEOp5SWC+MjSnmO8KjEBvBiJW4BbnmZ+quuuZSs1
VDz4GogzyALasiPl01KLUKHA0Rx/7JdQ0ZnUZyonFsJTJKRHVGQ3rNL0pqgv
T6FaJBP6eQfqkutfa5aUxiapRQZhaKJJB0StGwAFspxr595MEbtuRv+xLhvr
liGswLRGWdoDuQ5Pgb82QPzhZMWs7nABX5EyDZ9NZSmdhRWGC45RID1G5db1
B8FNGzyIoUrTCEf0xguKxxz+zhCJIEQHQtE6KdxMtE4UISZazOEGGkVezF0O
DiOwHE5ZiGYM1qg52WBl915tB0JWrNTtpKhsXHrtRtWnU/rwm5rDYOxk6N2l
MDCIBocD32C9ynpxFcnXTjkVr/ORrFvL8I8FBxj4COZSQHuwVc4F4gdI4OiL
Qer74cJpHpcRgSaavfPkMytrjNRCkKHsIjtLK05MbxJcpHYpZmPnSgiJ+v2G
ulupN+Hn505sGUw6w80QaJYkTRQZDaA7tW5yYBy840sw4uFweLIvKVSnsbSc
Hv0T6K2pPMRLyftqpdAPKvt5xf+cVwkXiYrL617OOW9Vo2N1LVrWifzAVCY4
sLMzgpHIdPcvS72X5V+FPFShaKMr7VtZZbjF2A2ehwQZCjROQG28Wzc9958M
BrtRmXl+UwWs55z1z8chEECLXSLgvnpmAIgMuJ7GH3H/q+W0vCr9Uyo3k7Ps
EO3SnJXpd0HBnVGXRIxpl+ugJREHL5+X/rpJa7f2O7LegtkwbUhb5E6nSitI
auvvKBbGJCsOIAkv4K7BVzQBIkMiYfULca5q7+6JVBfWJZoGFB7o1QehiwJd
1zpjzu7zTjszeaF45lzoafCpzR9ZamvqLMyMCEX6Obg7clVZrXvQbyiR2LOP
bbNSdLPYUsxUd8x/whZsMGjseyUIWWJO7iKBVxUn7tuirFX1AmxWNiTP1qeV
wmQGHFTEh1jU2J9RQ+fPu+nr7W+c+E7Xcsi3sGURrU0EGG1f0qy/ZOTyhmjP
2LCNXJMJr63NZ6zGty3JWQ7KkCJG+5uEoH3G6oIbL42/ckj8zJfQhqb/XxQj
MK5xm86Bj6Tl2uCTTrQgaZbtYL3MHhXLuVIhWoG5R7znLrdP33SNFDBAEmyg
tmzaOPFbdSjDNhRFYWfZZoOJsGSqwFzVQODY1L1HSo/f2VDvY6PmgyuNf+PD
lHxoeJMgE9+68n3FViSMq3gh2ATh0zQhKrlXYMIA5M7/f6/4xYEoZRwSTf/U
6a+26KuRPyCjgWKsIF/kC75LZp4WgqHOONLV+hHUzUkER51y3x0ttJEQ5rhd
OoSVL6CzErjTttcrBbl1mI8rHyGivrefywhhrNE+ZkL9MhYBJw2SJZZFy+Ev
b0DSaL07ZgC6PThDrL7/m2oMnhLNB1815H7XeTvWzZtvNzDnGWWGHAMTsKl/
JGW5/aQH4u82gnhJRFal9ye4I4C9cQ0Ap3S9FnEWoYDVSE3sK2XvSdDA8ViN
579W2gHl8gy30lKMunlFdGo894/dNMYVesUL1YPWQZzHgkCbYecYcnwuZ6YB
S1D3lHQWpKIiRX164DE8ryuZ0FbeyehelVtG8kRWSsFlXPqAMLzKhsaz46Pc
r0yp4m5ef+ABs7eLt2lUjIEnFzTQo9YApGv2mWZgp5cXLrSKKS9XOt3aTR6x
Q1nMBjNzBFYdHZdRaWkvsA+mHdJ1q1lOnupEEwOtKLeBXJu9eMQpBEHH3ibi
47zAsNDkH0wD0LBNz0Z5j4tqwB7Wn3juMheyN/eSGj9h5AxRg2klw75Nk9hc
dMqeky1PEJr4cPcDM8YiLbuCIh939YMOhFCXCK/NU7Thda31sLP1my+CqVq1
RqFT33pRIGiNRY1iJ1fsGs2QJG+nIc9CYBfVgUB3X9FcZI3Bw+3LleuHOXHo
94+3qQIqb+Z9vEVkxkC/2f05jdXvx0iWotAsYgGCPYzHf3XGPtiwslHKit8H
SNFzwQLOUvrTsKLkzxHhVxxqVKRYs3qVt6wENpD2mboJ09nSImYOR/K0rghA
NFaCwm47Zva3X+hIATIfI3nGV8FxA1kYwNXVaxotE7c/NSPdWDsPPpxFj2mk
g1k2flBoJGPPGFoBpNT1QF+xiFqUrj8PEMTmlQbMltNhIkctM6CF4PPtto82
xcC4B6QM1m9BBRxfkAA3U05eK0BD/cQ0Hz+2IZD/LD7AA0SPJebsHYpUo1N+
NhXjVosHCtHm8FxJ/DM9sTMHauCTbhQsTy9ivAhRSmtaGHiHFkLeFn2kq35S
Ld6btKC1Vr3Kr+pVwNqy1FuRgs8gVBMR2QM0bZBJ62l9n9shkmPhJ9v3TZDT
SJYceLc339CqXK8PAOSpRiNWUZsAytVLAjiWx+bDotnqM+AxQyaWNgp8ht5w
HDeBAuVQhLkrNcKhNaUeKVFLU5FMbq6XKzh/zE5ENa82drOm7wv/2rTEka+O
8+LXMLSIpFcvItypHQLzwW+9fVtqgrw/aL1DQ9OM86c53xBatNqCErlu9aeI
gHRnGYV4aDvjlFbRmtLE4ft6Oj/5hRu5Xo+c/MexiREjgO546HjcgEOPEkJ2
50V9EinLFwxtAHFIPDlXSvs7nHOm9V0YJ/eMlLV94/1drKxdmSSV9oNQhjYL
dFTJi8jxLJjIvMrpXFYoRPU2nU9DsPU1t60o3JgIdZCCG36WXULrUxgKd5pd
AZKxx/ASWLKqWiZKYCQ5oC2u/CBh74lIwzalGfHy/WeG2CJ46mz83N84Dddf
wZyry7woJUz9D5iaWQyoiSE34DlVPYqGFiSV80YKoxHPemynqgu4xrYmWA48
xviq+FL+wZpq5AtobDqDyl5aqqiy+ElkPw8bcHm7YRBhlTAiNKY0MAX7iTRN
Atz+CI8v26nUmjQIav010kkG6G6bVXDud+pRNQmB5+DtGJKAvdyDEvSwNs3s
V0rVWIxnYCAw0JHVHX12VeT30BR+Z4Lkb+C56Zq6yuhfkK7ELqOXiEh/2Ruk
ddKlraGgHcmOiBMNTBPwiHsIs4ghqk1g+zl6QmFjx0TVT3uhvgmxBPcI7wFZ
N1YwBbDD5rMq5fMUCODnpl9RZ/NhzFta5caWHeGT0ULtbgM0OYWMw/kCWheD
iU56RNwJu7JuxPQsJsrL3bBFd8oxqWttW+oefro2MrzvL8gjvLg0FQNYA05t
5kPI25u7ERBHnXM7YS1cuarIva5HVdRuvaD7bdR6Q2rrsd+/zmn5vvVlSEUQ
RuJyWr/zu1jiGWoIh6v2Y6zXBaTbDJdnwJxIz9i1TDSalMIOf0l/AR4hdM6K
YZegAu0a0lX3d7SQOsbgXDxOs+Bo6yxYj6l+TKWD0MNjE341cTplLGC97H+T
TQpd6hWzK2u9H+/dO/gIJtMLLJpnTZlsOSdTdoTcmbA+AHBZsPMsIMilaMsT
7YQKzxj866im9SD4CJBwaeGeUGgXqnLWRtHBOnAGSAGBQ4f3LgF2OMzGdcXg
EZwjuID8Ch1cHYaS5j0y+03h0W9kFEl0rxmeeeabko6XEjrbMyFRCanQ3hqd
aleYnlyYRO4/O0k0uyIdZ1oXNLDT+pWfgmV4ZBfL2puYsaflcC2qtOg82I5d
IHvh2cvDUwn418XiACnm+D+qyWu4iASY5UYR73NOOpnMpGdTSVmQg9TAS6RC
J4jA12mtaUSsZMtbh+jzXFV+Dl33ERWlxp0ctsMX9zev/xL2Z7SI4d3Vpvja
d8hFHWKso8nhqKuZWACGAvGfMEUtSBefhhaCZq0/spu3WR5hMJFwMS1wDXQt
vAzhneF4OXqrbSQ/6vIBlxEqpS+hy8nCuKnfFB1PBiRVYXpEAqTWl6YTA69A
snDRCIf3Fm+ex4t8vh9tvS9hQxiz/9wMebLT8SJhuWwoiu1ih8uhxfu5encn
X26XMMo5k4FTBkjtM3xYJZgdT8i9Hu5cA8twYOO2iQbfZbl0XxPEfofwpMAp
w6BePt7gzUvANchBTIKP25D/b1u5j5JGd/nlj8O+OpzL/W55XAxGTQ5VAXuA
+eEppoatL89KSR4HHpZnEvW+Z6ugwOSG4zBnlAe754usRtsnl4GY0Zpb23aK
xNKZrg9mNUZqpnS2LssDXY4lVs4KQZEcDTmaeZpJekUduZdRgB3fSW0J6TRo
U+R1A9U5Bu7wiGmQ5sP+ia0izKZopHuJgIqNW94qv0LKiPy516ewO+hG0VZJ
ZNCkivim1xN55JTmxbb6blmlDYH/cbOXud0CpaZUVtZLQ4T1WqYSNrMHr1BX
nqKT6gIycpwiH3wYtybGutK/BLsxUcxrNtXCjnckk17GrW5lU1ftBDCEMHkW
NrLdTaN2VUz4y7txnbXFhscQJcmeXXKKdGxRhSDlcRqoBSCgyh5GvIY0x63k
F/ssTuQjr7f6K0HhHCQgqtDzZOkOcmDKZCu7YWZnLUwlS01j/BqcXaRH7Phn
zcum9KpC1sxKhW/Nrb/FUG/m4iaANBu8+us5XvT8R/EHybRsmBViyknE1RzM
IEDOjO2/P3v2xHADLJVLU+znJjSG7zLNaAS8+qmCDgT74pDJb1GETBb/wBLh
OJNbmCQUelTgIj9CKoJKylDVMtoFwy+ykhaH6IR0IPBPrExxM+gZwARIn5Qm
t1GY1LCLa2fHUsVhIhici/QP8Zn8qqDLG76a3btHEqZZ/ZpFsvKh1eeHJ7+n
EjXScw74PJXXOOUYJRFLzjZFxOTVTbe+OGwmmfakzirn0WnK33ZqXL/t9XLC
PapN4y0m9/O420ETIFpf42Zy0P0d510HXd4PGXgEp+9xw2M7fGwvUBvR3lQ3
mYV7dN3jd6reONOdlW8IYry/BwnojrTGhYV5F14gfZcCjYmzWxtZg4F6w3CS
vpXyv1pP1q4PtUXXGdCOHx8z/iw3WXno9GZAhg27ZA7/9n8rG82uAR5zA4CT
YY5zcVptmw6F8bL7iNs2FkIg9gYWa5YcLcvSS3wDsuFD9j9mvZibBALHpvqu
I91UvN93A3lpX+M2HwzSXYhYq8N46G5+ovMCTCN7N0xm+eslcoyI902S/5G6
QhMJ83AVVThd/yFfnd8jySF6OxLJrVHNFjCnnYjBUoxBl5vTw5CR8hfowgq2
zapWm3eZES92DRO3TftOSs+b+nOQeYcIQmIlefn0Q1md7djda9Q5mxdDWj9X
BWwuggh69bfe55M3vkIDbcM0F0e+XaAktKRjjbj3YXLfMA2pUIO9rpgxlroz
in6mrLhIyL1GnldrN+MJbNaC505OcrMNa3iZhFFT3d600PdtcB4+6B8ssBN5
a/CsZ2q4V4ylcxKCcF4AUndxpq6SNcNw7QeLolu7BNbiJslDEJzk2X1fauot
I6cVr3XBNIRj/DYXxDW6RBhNNpYxGMW4Goblf/HzdYwAEdUiB/QPX0yBvKKe
hth8ij6AJZ1LuFMMamv7RUkw2dp0TNzqjEdSSPOW9MDF+1McZxoHKZLn0jRQ
sdvQSssQV6GpzUchURF+jBFqWoXw0bX6M9BNUp5+/+YERCRH8+JfAhk1ulx9
Oa7n2Fg6PKyd6r52wWyncgEb9qsVG62prKVWg5M01DNeh0mQH/9yRgZKjfoC
F9Tbpy7YImLqvXz8Q5olCfYQqATVXEhfsIVRu2yAoBqnPYJIE/NO2lFWk5Qh
cq37o3bBUGK0V5bH0tCR7AkH5JnAZj5Fmicxh/iLkTjRzTa3hvuq6lnZ2p4N
GODDleyBsAGnlUeQ1o6OiWpz6ALQpu45BLz6sBNkmrIu4cSdg8zolsCxG4/P
jY31TTNJWREQZaUFSc9U0k2p6JGDqox/byVJBgkmqgdHC2TN880h93j+lEAy
5njCwGwdLYZCSKvXb5y79uwI9uU+SlLqybUe2aNmMl8SRwbiWKww7U49SpC4
o8yfA5P42V9ubssIv6ZYdV5uWhqiNun+agCKU1+VaLIwa0o6xGKOZpKPo0Me
aFc0Df4h4ycHGPgShUH0gfqgFDDJ8hGUBbQ2mXu6sZ9NpI7tPrwP0VkbQF3K
ODAtCPxgI6dTo+DzF2vAQGw+a3swsRaF7g8fd6bIvpjIJrMDl2MGiPF6pAxV
kiZJ8CPfBPn9/z/GW/k+R4PPFTRTnRKP6vX9hYeksquRnc5f+xYnhijFnR3O
HRKOqLJ/hbCIeIujGWJ5ezqdnrfvX6GQpLL/3OldX2CRwwPbvx+/y/1sG32V
cTs5SxMD1FyJBY4cPaMV910F6RmRe0P+H+1OylegFqYQ8UEc3UgpJD4gLRuf
mWBfWRfid+kvIgbB3XLufXsdkuqwNEYxcTWZaLE17ndfaHwzspSzyLPU+Fp8
msneiFUCmGehHAt8ED54OPx5c1UkLAF/34bR72VBQ0LwADQpVqaidTDucEGX
HsJVfdYLaR38P+21wCJBBghYk8rpTtMhtSIUJdhq0ZD2vCJfO2hFSe3yc/Lb
qJgoFC3ZAch8Vxjrjy8SkUMxaoGocYHR7ITVv2gs1fhDJ9cqsINJGUEpTOtU
QXNw5JWQ+SYAVYr8FDmvvW6PatlyV2kq4oropZ0BqKxO65PMv7bsbD6Xo3V6
RBpb8Fg9t2y2Yh41Z+j1dm33M5sjJ3XCslV2TYCACYcezPIpKzR+ltpokQLT
R79t0mttHzPVue4fHecI+If3yu3K9KXMfXNFujhZSyJGLZxm5MqTlYnJX288
k6pTKhQ9pxuHxvFYlTUuIXfyimd1P8L5HlrE0CZcWWY46aLcDme0xowArZx4
1K8QGgsi/lX7cOVojuWwK2Hmd6Y/1X0dlFwYfRKi/mCKL9JhDod59OBGe8re
K7TNvwtL8b50j+MZAD2Yor0BlxT25zQw5ZPeYFHlzBb2BGYbTvSHsW2n/AR8
fqQNkTJtzYOroPx8HIE/eYovPKNkhNBy/4is/6kCzjQCj4oekbUTavNOrMTO
btpexHZoDwHVonTUlREbkufi513X9KVMmA4Pr9rWRJtHU3FfAjWA5vFpbJU5
V0UHofIIGIct7Jr6qyw0cn9sz+pOgvgoOUF84A6+YjxrHmN0c1FDSYUn7PCl
QChVq6FQqoti/HizX6BXVYQBnHgBbQ4nqdDc1/l83OFfZSJJEKLhXUHUsH72
HDmq1stsGj0Eu9LyxWnGMkiVzRPnwH2B0TdCq6L/C8cjyb3pK6ol7uK72mUF
kCI2Jk91sxmIMjSREnFeKFmamM9goD6DGraBeKWzdaG2USpYIxuQfxGKF5YU
UKOejfziilGU2lxkpx/iCqbN2h5yzM3fNEEMjBidzz96VIvNQqeLoinNoD5O
ugIbZZjtn8BRzy15lR00tRkEmu5cmYwpU0oc2Iurr9t/DTKfbd1TZUXV9Nf+
2ieZa0TsYcm0StBhjPg/fgH6AJwCe8vH49tlO0KNo5ph4EF4x3O3UeAmLSxY
j6WUDvdLkpXV8kgrZAJ6mwQwI7IQt4obbb78RyY7HxXRMQ8JiBmM+c+exD3Y
/+ZwgrKYJ3YbS+OLvQkzLLfk9xfQO3CAXHU2cvlysoZ28Cnl3wrjRGC5KjB6
H3pn/RoMeMSd+WcP//trq9qJUL/rc0+BTlVw6LiTrePLs6jHTMxRQ1y/U2Hi
8EdnOUxc6wXe1/FmFBquX6EVnRWH9uWXQHuwvBBGHA4rGtYmpkPTNpEHNnQO
lY+FNP13lm+e+gGXbIlRAdJs5oATV+zKvpTSJ/x/RY17l08Iy+RNNyrUkeuK
shYS0751MyJDpoQRe0wUXYEdEV7oIpFxIabsMEX7CyCh54amr4eXdKOMC7Nh
ZNAP5gsc/ox5HtX6jeMvMGb6+dZzQxSUEzX3PbQ0KkjtkTC5WQeQdeR8JPYN
+4UBOFUDcal04NaohYGh6IRwLFDEHj5BlxeKwycr2dK0+vpxn1OBEcKzh4go
nPBsueoAHhQrTAdhd4InEAhnWNpc3oaSXJl1YwMI7LIK1sht4eMxKA4wbjdl
rHWtLUcagPvOnGRHXT/dvx0DmqZWFvaM+PB3XvyVxbWSoWVLzfSXlklloTTQ
fBtAOgFvphC7nAtuhoyIO0sU3Qe0nO6FgTMQ9hVGQTSsRKnPwhG8PPHiUw7d
Yzcl0MAvXOuXctRWsuEPl0TfZeycbgDwd+zKVlAaAHwfBI7v/5BGLvoL5nDC
lPmn5BaI9FXj+nOhhtx2y61RfVeg6Fdt5raCXUAawO7ABnfNwIwnO8ty/rMd
C5zOoNFi3St/GBh7irgWX8QnTgxK0oZXGBngNgdylAcC9dq99X5DHANJZ0x9
jOg+FA4p56enbxhVwPWA/LIXN92pOKHTXymSNPZQhXyorWqdqT703AZqSJAo
zt2ndYNFFNIiHV+jCPKGvsIJps3KHjNARpDar+tunMdSMSNSjGGut9l2u6Ks
lAxuZoEkzMfAVqP/mXAPCLuA3Rc3iJB8417ip2MtHN8+VDwnuZg8L4MVzCCo
puKlggUhGSqAlOthttazj1XJegF3+YF3JXJlghjQ8XJeNMFc0cMx2YFYSsK/
Z4jYOSLIxBpeySbOn6/Qb43HBwCs9G46OuNdxDC9gB+dHyR7NZYA4BD8JKGt
6qxpuJHzKj8rT1uFjFOCz3y8XJ/zO4BH5X+JMmDj7wdPdDa/4+JwrsurXFan
kUYDFZfDyXzbM6U07IXHOkVcBzDrfRJXjt3Rjh4iJ08XbpyiP0frQ4r9ZGez
5+itVrEvvPYNyKBwHJoxr9WpS3TPYEmFaiH9eOhWFma//c0Z3buil2l54nTq
4M45xkreu5iK7kChG+7oxIYP9lsmw/ARveYt/BPMxfxNCSYpdmozXQx1/Tw2
8D2wuxTS9ZyL/suEnBbiyU6bViWXpOj4tNMtG5r51E47v/ZX7scQMm+8y9Sr
N4khjBJ6h/X347ulXtq4lZQ9gq3SPIor1wfu14AZoWrKb65/9FLvas0dOHy1
GUgdjglMckxvsc5UrYLndwwMW7wBq3+vQigXTt9eF+1J8JEDy/a+c3ChhtW6
EEUC+C3yXtfpWqbAe3O54tsFenb9l0nHm5fYyknO4970AH34EWQmGZ4sCfeG
PAltaonB8w1R4g+7uZ26bp/NpPnDacqRn3lywHZpKqiFR3+K6WuTA+yozAEH
kyu68J26FW0Vo7rOF+5DOCVNhIsdxc4kEyAfKpmOXEijpcjJnTX/QqrGxyFj
Jf2L5IJDwWv9KdHmye69ttOOUSpT0IqlW+fELDyHJo42IgNnW75mQ6eV47I0
SOHORx/fKr8h2qtEOwMuGzC9NoCEfu9r4lT955gqQF8vKTB+37BInkoup2vK
V3XYvx7T1xrJPs0XWd9c51P4CvQ89TNp97iMYHUTJ+gYN1FYsvyvz/ipgiZG
suXhewsAuz9UFVLxhn8YmmQvGUshacza/0Qp2fJ615trauulBj8eVmt2T3uH
HyqWB+mdnZ6ejRxeQBAxp9cZhV8QMKByjdqNqe1fyfh/btnPg/3XZkDMTntQ
fzRSjPbP7UZsnwxq+slQUZ9ONCKsx2b2oZ9vzb2v24zhD3KQfuHHB1GsfEoj
KgoSuK5fHVS4NuNmr22E8BIX4qduO84/v58mYwIMq/yyh22xbx9woo0NEL0K
HAg2hDmLBJi4R8M178h9RdduuZY5PzxiN9iymqYLAzQvW/chsmFXReFhTUuv
UmtVsJHgb8+WnEVMyEN/Oo/xMb8vhzOw8LFh4IuKOmhQnX+DQWZ48WpzmERB
Hx7S5+ZWrQeAjEMyvjb0TnDrYBPH2eZwMnnL6jYD5mRcXae8CIKWyRjkGJv6
9DTyijNbA9K42tUd4A9N3bozFZkwaENLA+YwTnH49vbI+lLNVPGBrLpnuxxb
f4uirXXKEY47AeNJCKDsPqv5TOUhr63th7C3lAQlkUj9PkztG8oaNWa/inhE
vIIxkpwJSgjSWHTrWLjTys2c53vhNBXXtpwBQAKB1V2JxDdOmHMuZoybdZ6v
LLDg2Dmz0z2qu55jf5pav1vWBk1GilSIyCv6xNm3+5kaO/ZtgrfMmvJgfC7I
uArfMr2zCsBSd5zOZU6nJPuT8DU3Bd9Fqn2qd1/SWllZ9LjUbzAuL1QXp3RU
+rsKnghpLr7dvXUHAbe0/t8adI011fnjIsHZCaG2bpmz6j3njDvHnZ1Yalbe
B2IFqasFZ2VR1eHG/3jxSOFJwD4PLBw6gCfMr7cai2+v+8ThdDHkU69mA4JT
3/zN66QRowhRdeJxHa7xvUTWJi1tDgQXUq83GIL3fWNSskaa5QL6agPoUq4T
u5Rydw/t3eB3saW+kUaL0YaXVAfd11SAfckUDZg30foNHuwaPVyDdIZNzqLh
WZrq+Qz4FMd9GNx+CZfYHHEB/LEdfQ38t0+oHH/ED1VC8z5d/oO7w9z85ToX
y8AYBMM6OCKsAPFg1nGz3Ga0CygRFNyufpz/AFvxyVennpLJbVPw/AyZfHwj
d9BNxXBl64FviyEJ+P6CuUwrS+18P+fBhXkuUh/GmbD5xzKTp+4yBkjQKO9K
L7eXBEUO5yI0nzHbEFpMt3I7Ut4mhwiWra62vC0neHaKB8RT7jr4mk+CU3+4
Sft1PEhqYmC331DvQ5P76JFQw9mHl75XSu5txBbsG0HfwFIQFLKu+FxcIjhB
QMAkZrlX7BtIX84fkH5yEfWluvJ45BIEBFjjialtXOeY6KYU/PRwo05mV0Pl
syM+phu1gcyULV+BAHyAkUsRYvmlRfUNUgOQMdkAM1TMhTZG1Qf49z3A2Pyu
YDc2jJtQlCbmHwYUqQrXQjkcAiurAD473SK5zJQP9nq6INy6UjEypliXLiun
+9JWrMbWIUQjtsfkniMI4ZguZDjzhthUUZmdm0dKxYmTN9cqOzPrd38AFdV1
qyFeg5Ib2hP9M4O3cVM5wLZuv6EbN7GHUCg+eZ/eUoBcT8ix7Jrb+2hKkk63
dTmGt3jiM2KnhURHE++N37bvda/r1zGRWBM6ZH05aK6Yp332p0hUosK2PS8J
teknYyOTK75RkbqynOr3ud0BnPvwL1DpD7y6vvb59/WIq/GH21axS50YidfE
Twb6Ub9MGOHwSgddzw3tZ76s7ZEul2V8vjtq+Cz9X0iGku2b48+LgK8U+HE0
2NdPBSGP2rICXH7qZvm2nnhYmrmC3QWZvBSfFnVTUUFfQC+WX5gPO7OrPp6g
qLbnnNbD3aIwQwIDqT9zLRT47X+NbZIJGr6xtbRylBdYtKemmEfvANBENfaU
YAF11MnM2NENNF0IAQf1nEHkhPemA4j4sbL62OhXxiPdaMVTfF/L5OQMKc50
abr47Txke0bLClvttjfSBRU8W1pKVCNqFDm9j5hlZ9urwT5QRYPuKCaL5wg0
H0Hqqrt8b5zQ0dJq2qI2ibTcA30E/A51BxvsQSyj6zKDI4B7Z49aPuPYyLCd
VPFrlb7j52gBYcav++dcUIo3LJmNjjjwDidrIWQ82flmOus9zcU8NEdCj9pj
sxlRxfRo66fOsyad1BRldlOSYDGQuMYF3Jh8yhNix8PxJNVAgWNd3jITjsWh
MtRiJVf8koetb3CTXrJyx554zW01SKwKJVhS5e7Mo/DZK84OSLOFA8jlr9vb
KdojgXN/pR84ART7q3LK7kud6Z/bPaIEmnOEPdJmpqsU8LfRnbnggt8xJfqA
j5MHOBG5FYTKftHnCNidlO8ik7qhvE4sseZmvRCrD5+QZFO0NFvV1mbEc1RZ
tKgJBxMlPzA4CvyJBhBH6DDLrSdF+ScmhSWURjIUYi0KLC/u8c4vSmyEsK/I
QNgIbImxQ7Yff1gf+4teMR1YsMbvwbv6IXYxFVNXNhW3U5JiTKv8pPvi/weO
UH6ZOyP0EXnRMTQzhnc/fDs4171+Pqfq1GSV903j3XgBRAp4dhDDCGbBTqVh
1ywvdjiM0QmloHpNUM+WKwyokPVPxdcQPMqcdV2/uFnbu8cx5RgjbruR0y2H
Wm+Y03irYOgrMizRK4jL6JficOAp4N7H5G0F0vL9InAT4ef+WALheLDD+eRU
2E87PNxdarsoZ659MUOi+K477LiSgMLr2PvwyVZuwtNVI7n3OsZzGU36jtpM
qJd4+PwrVUMvw20sdvCDCnzLXKR9JDddhJfNUxkP9r5/8UT5YJdTrJ5JIweU
S8hL3UnRY8EkZe+cAXUJjSzGcgrtvJ6VZM/N9gnloA2d/gt6E5RYbDYfWhjl
tap83E9md34D+HVyH9IctcvZExlXtUbP9UJC/Qxk1cR07lqwdHth4RsLUr7q
MxNHNCwl0A3ZY1stcSDsiQF2cD7XF0tdbjWQ0NrrRjTjwPiwgFSKUEDwG6ds
bpiR4Ts1E0ZDLFvkpyV2GXn9RJt/wZW3E+jq6JzFaqh5BMkc5yl20DGFGYK6
L4n5fgnG4yfvSUI6f7HzSOI3lKo6h9WU2aEU13gfcZtdvv3aL+RdNUOJllQU
0SM0O0A+vMDdkHh8o0rx9lBeePkpQjmA1pl8AApD0PwWBpN49eq4pwd4JfpY
02AIzOt+NfiqmnXpL/A8FgpZRRsCQ3SotxPCI45aVqrrhhi190DjZ9X6FTVM
GacDTQGR5y/lJlWCd4gqQY2CjLPKhTvCSb97zRppzVbR2fV4IEGLNfPmhyqc
FVhwawK07wR3j2oiACRMjix2TDsWRoKgN0ujzeSrgJPSXYYxjwWv+Mw+EKiz
VmEgpf7h1+InQ9vjxJDaPCIfle7EqhCHwn51KKViOyWjiG8Qy0LPskjAq5Us
Pp13QcO9AX5K2HPywbnBqeYIp5aLlRaujaG+UIOldfqrfNPyEqFdJUBomnYx
G4xLzwqT6PFwQNqJc0IMdmjT96gxxD5gH2Og7OilzIQgUZ0DOSU8EfOWllBp
DVDTzHxSGxaFvUQ2ISG6ajp/SRaeLfbeERZsaNyzX8Uy7Dr4TVtwsmnJPHDN
bqfasGfis9aKVuBK9qi2R0o2TPTUzUpq9Ns3+Fuee8cs2n4nN02KVscfXcHS
J+LAGTcIaTahrUW3BMtbgZkzg13QVjmeWgIQmeVneMq6uutYALhiM6cQk8jK
TR5zxjxLTpCV3ozGAXayXHyKOqNn6KgK7wwrgGJDdscLq4Tp9I5rLA5RYzip
JV0e58gJSo0W1q4V8BJb0CSyg78t256PMCEVKRbICeY5FGLlwnxF35G0Yi8H
meTzlgkFtKwJ2Ov8RVXH5W4o41j8ZqAjaklECORcwarkhDo9pTiMBJyp3Umf
tDUPhGt0rFbtkwfR33/EGgb5F+z7OoapSkCPQCKky1ShcZwkWRQgnopifuL8
96hd/d90FqcNqP69H6cSStlVNs9Z5q4s1q8O6aEcAn4X7dEXvUVkKp1Ywx9f
MLNviH8zLq1IdGxLC4JPA0QvD7XlaexxacaGE4EFa7x/9YuDDAkWpz9sN/pi
1vIFQiw2vrC3qukg8RJVFptLxw4yrej37sRSxEeGsbKwdXSLaTrQ5D523wJ1
SfstpWCK9qGDNdTNbnoabw3LYD2IJ4cq+vkX+/1mMi0DlOZGGRFFNVjORH6e
7xKIh6a4VCpeJ/tmFPYoWL1NXFSH6PnIH7E9hMvymbmh0Qp27g6dHOmBXq7m
WNF0VutlMZo4bx8NKHjfuJM2xSK50XVbem+/AT7tLgdaTmujIU7wWDUAo3Do
kwflZiZcjPYgQfNzyHx7Xg6qJxc6TVsiyjIB2oFSSHF0tBqzyVrd4w0AW+FI
AMsEBobm96NMO0BpNBZqNFHAns1DHLEUFlUBWUaoUjLnSAi5LXIlvuWyn/Ef
0HTuaUVS4m0uZMqcrjBIDF80nGhWMtPiXW0GbZj/By2QcJxRijwOlsTvmDFY
gS6Ys5mrqm5ZwZbClKQq2V4rE5cEcm/bQ+cgSxuTFFokoQOWtsA7j2A8yPDZ
LEVwNKpulVXWVg+M9iIW5VySZ3scBN0F+Jy7h1W/eXZdX9hUoYrTSpXonlch
jfsLFPQT+6iWHiZmRUO4pEbQZ9Dwn7ieP9iCqK+MzrUTF6fd4wZ39WZRNM+8
PgdUMF+a7wQKiMPNypBnEIciIAhIOWS9BsG/Jym89oFzCGMvcaWoI+YTV+vm
4S4Pr70PcGYUMaR6wT4PSfWljBywB4tM4P+pfl7rL2dnDcLmkkoOxExRbdCt
rIdCxG9J7p2fVR1xoN6zpnSXE07f5dVKvutN/K8Di6CtA94Jo0AQd5M4Cd6I
BhlQEMAmHWYkDkWydUMl6hz7clteBReUJmPq6MJBoIEiL0AENx1lL5X1IXl+
UaH+aheev1qin9pfwG6+PxlFQbb/wf8FQT3lRfV/56O/aAJLLs59O272eDMr
X4EOiDZmuOHZ3r+6U0jjkIY+JgW2BNplvJArxtnDsFa2bp910abYiG4frVQF
yhBc6zg7FGJD4XX++O5md7B2JDThOF7C3g6F8eGoWVq7m2XMD/bbIR5Kf+Ce
2jXf09rINImuDgJ8P48CJN34eB18wQe8rs0WPMokV0ZLpeTtSP4RNYeRlzwj
ro5qjQNiwoqpq+UobwaNWed88Z2QO4SYZpTdENV29nIe0xdG6yUKNaXeqzkS
0Ce5QqnzDhS73Rke5CVBUqOEqeG/vGgWqR0DC0w4nx17rLL2cM8SvCLNdWU/
QDwCCTOgembKz7ToqyVyasSGMUz3SnEhAUY42RlgHreoKSI3L5FVMTPEWr9I
bgIEEh207dLfzkCS5MOlRrXm9LzetEsG5+2837XHgIRvsWdktGcSp0wGI/eQ
yavrF0pDSbOj7gqJXquhC1/CsnjxE7fGqNgqKlwh1BwStaDNNlKs+oeoqrXf
Oa/WzSbRCKUg2yb+r9usnVrXokQ3soyC5Bs+JE0M23QQCBSsqiXv23swZxRf
vwEv9HIJE/2KH9aIwoiiGMxfLxD6lGfM0J+Ft/YE7m/Y+upsGU7GRpGAAJdd
Pe2C0iDoic8QvXAqtdJ0b8SOQVd4ZANqQT20pWHRC6lV9uwelVmLZrIByYh0
9n/Cuge1OSK9wcNCmo7wJQPYmuNOns64htVX1hffI63tYxaL5SmiMQtQplqQ
0coA/fhJw5mgX0GSFJw6LlSfNUQUdpUFup6Zq1cLWZnZPuaroRQFqjXxSqkV
5vglkk2yMIOrzAdsCGXextW40cb56GmhOTT4/F4EIbR1kkCG5YGPk1Iayoez
dOuw/tuc6pVwImpNV7kI3w7clMpX9VCw0kGqqOU9bG42jnzPND14gM/rTEhE
dSi2bIV/0HN3jyUewYzMYnmvYsL4LV1kTmHe7R7z+HJhFRoTZnvbXS/TGXhj
eN4GmZI8d3IBITlmtJzs74V1+erVZcqTRdpNHxbWxDxleRDdSCRNJHJaSoTK
sFcQuzU588uQ+oxoqN5zP1+VPpQqERz5T1Vsy1BLuRIdpPwslPJJejm9r5Yg
JTMLWv/AWiuQYmzJxEy984Og3q3XKU6ImNzcLGmX28CjY9i9S6x/kBDGdUZT
P5ZehDnteK3RiBVJKTOlSKg4TdXqPsnjWewv/8qyYiXbrs1DWMap+2cmj1cg
YLl07kaAHe+bB1smanz8Z//dsSJzr6rrwap+rma+K6/nRCJmSi7BN/H8umCj
mlCH20k4ZJVW3WELIgRGSPJakCCONy50ebYLOEIFg5FW3YJ7kPoyF0Zg5Wlq
Z3DR769t2o2TNmJ026gan16jP4jyz5h/4ZDSXKLW9qsFej5vZAXQdUbN41nB
XB5UwnZAD5umfhwPexMQRsgM+roVWza7pMTlH+thA6cuZB59J7A5nFySVwuW
cEQ4NBHuuYoTh7GbEMFCFUoZiwaTB/pk7/hUMXI6Jx9YaBSjqLZvDtzPJ2w8
1lny39zeSkNS2/lJNrkaXYJjwIAlEr5/Yk9glrG7+n3cSYT0JnN7djjTAelK
6mqgFq/3Py3Hf76Qj+ZyOTaUMDAPncIy5qO2g1ef79GMDWiPbYQLchgo7QCb
1Vd0C4PepOZk3D/xiT1CKv3aDHSz5nMfAoS94hYqxur387YqUFOFDC6uyeSp
CxtILwGtR1xPH1Nos8d0D6g5+2vzIU6UAqTw+7W4hJ2ooksiGtQVCZZZkXH1
EqvgZSBseevl1/gAQ8XlZbdqDFpfFjfujd4Y+UXjf0k5Sfz3BHeVgFhIW2Hx
2u//GG+Nlu2Zjza0aq+oy8O9glH9NFWj91pXJ3EzhZr7qwua6opOAkqa8LFy
7Oc1y/oM/Ai7wkGyk+O9DwIt3BVvF1pVRDXQ/amDTJgwcnhtSWBn6JCpiT6w
zPqiNXSccxlB08b+APQe/VDV8qJodU3v8wu0CptkJOJZfumP3oSfqGEfCdDU
qEyj0pPqdjDQy/9ZfOgvadus58jwwQY133fR7IdZGfxqf9HEDjQU6p13H8kn
T9mIDtidJrww0GW/0h5MT8KPPpNsdTRxrQb654g0XU0M06YYHypGEj9OwMIw
UTIWGbFjSQhx/CfDITFJG8GRboT2jPmz1BqqvDj4eQcVXE7LRwct3I/z7fF6
PVNW0HQU5oYmZFyC4kizq++2+XaJfVLw3li+p1nk24D4Ci5ykBfZSSkyvLGY
JF1sp5i884okOdx+s3YmXTVwf1A21PdGjCgHRQXFakG2tJiffaOJD2PduQC2
w6N0x8OFG2v9I9IUD+yPk5+6iu2ZWW6oq272wZomVL2LJuqW//bLh66Xadnb
aA0y3OH1UbqwS0aIKu5wO6PW4/x4VtB0UdZbyuVRzxzxqh90a7ztcdsTBVPY
LsAqmK3RDsNz1GEkPAEhh13zSDrN8SIFBERIgwbhmQq0+VjX+MVWlRC7jK+3
+uvyJuJTITtDe6uBPeUfKSOPkxqUCKOCChoOdP5PAbOIlfN0RJFU+E8jQywv
DEsrW+vzMJ3yYU2M+JlitXoCUhh9zHikEqGh1AL+p0PIkmzjeUqoZyWXLuBg
IDXkecJ3D9biZ86N+7VsJjRL3ArHDcOFH4SjHbdKjZsNq7HGNDgDJm3Z0rpt
DbU5MgildYltELdQ8UcDSnV+fFvDfFXuYNWY3L4jlfLR+At0bjEzbxnNqAEE
7hwchndmZDR2IX5c9zn6HpYKZ3YW5kI10YlSac26wk4hGeRqZQ6kjmqN+mt+
ADypJIMPHSuRkCXXhTzdWJgM8delNQewR8WTcOEY8cpE0md5iJ7BsCWYRWNP
ditB8PJ1mourWvjpBZB//Eu3++lk2F3Fkz3PgqtMU8vwvT5F9PBDAF9mjZ2/
btUneKcFOc2KhlaGiVlbvlzkWV63l/8EBw40tLhKlgxJTK3uAQx/2aV+YkSo
q4ZCCKZCOIoeAzRH4q/YEGeHPk2X9Bz3gBfmYA+mipzKnyBi5Y/O1jnxPVNL
bUBwjWcHX4AEVEwcBYj5M0uyyHc2M1O++WSXUx7THE44JEhOrr3GCslHCRDk
O+WIi7Xgu44Jq6H7jvewKUh3hcTTIZ865Ya7kc+yollrXIpeMhYhF1d2PQIY
bWR+viuSbuhekWDGCD4jCg2V6koMf3wKT18DM9P7hg4wAYeeMlQupUa76Jqa
LItAG5OGA/S6rrkJZmTlDLYWr64sKR4GWnmPPN7fjw9TJFBjcAw0QWo2WSjI
5Khb/0mG9Jo3iFkytyFtyTZbfG5ulGCyCkVylCwzH3aDA9ZFT66stXVQzcr2
V/2SKXOYxw7IN03Ls6rcVKRB8/diHHLU1smNBvlUtJjk179sBGsHNqNb9yXB
OH+/fBkTANybxgXTx6lp7VI60n12sz2PBTxXieArgSF+ENjjZYEIvU4+J6IL
ybN1bjJfFyIdPYc3roKqrBrwACOKRXzlQOT4KxLY/242oOuooigW9WqjEa2A
KOvqFCgh9gs9QFihxhqHfbIbww96L+B3fPsj9fSW4cpwP2UjnlDKHcjmwDg0
DG66lRkj7aNRJOLIysnC1RxmzlNgOuDAJrTdBCwy+wI0NZqm4SX3XdKEFCAh
k0f2NQYQan5fWcpLvxRQRctU2KjRFAfReq+zHUOHcPS1nZq+d/VG/hMTGoBT
Zt6uy00zcuXNWJ1UgFk10UDO1lA8a/xoBf5dm1IogVSAG1uIfEt9b8CNH6a3
jxjiB1jab8on1DIYls1+jrrXxILksJmH+Qvy+pVKZGMkDKn9FRipryJvY50I
LbpKIhz+wXcMJotd2tZvOGNAog8Wx2iZmjEwfqTh9ai9Ly8cHW14mxJmJdaf
kaRoQKIq5R0DMW9zKljhMLoQhCaoYWwlVH3WjXbQ5DkWLG+3OAEnOJpLXt4j
uwhrxt89CEoiveMRZiiPtzSyvHN1r6OcaxRenlSaXGSOkNBTM0N+eMAXUylv
CdsRiEss17PfezXHObWM+UsJNcs/iYayKRAPIsHrG4sXhFQqbyVcw1CuTvOw
kHcMoaykdSu3UHUhMbEYm/TcnOoG3cl0OA4Kho4FxajxhT+DFfHNpn/LyEot
NDqtvSwseb3+2+YQegWrNuacS/QSeGUjIlablPMiFVy8IGyHJbfgEedixMDb
tzPlQjk9waJ5ICCsueGx2ZCDZdxRrRlDhgzEbwj7yS80kqTU2gwGCmcF2ZHo
FuqvsZQw+6ykG7SAam3rjW1KWhs7qCt+C6CLO6rCPsBmrt4L6Q5mXCZT0cE1
4ieRahfFB2DqD50pa5ZQ4rsQy4W5PyiCa6I5HmCXOjr+vIlDj60vkQb59dco
wbIhwqvmFvoLZDYCyGXZQGE8cz0AFfBfEns7t3FG9SLUJqQ0/fgJlSXUZ8BS
EgNwlkEKR2jLGgQj/gVd3LIc5Y5QXTTsx7JG0Lsm771EhV1PFDn96dBq7IAM
gajhIRhkJLs7MRL2vZ3xEnnkewsVNPKl1Z2ElSRlZ5ht/WaEyJJ9V41GiPre
e4Z3ZYjDN9nQfc+18FyCqqU1W0OuznTEoue4Fc5GEmpgwUdZKImwvSbJSunG
tTBCn7sNjSQ+ukA6Us7oXkzByl+jQS5mM22WtTOM0nPLHhlOBMS742HSATdb
fz2mG4adqtNXJKEfrJieFT22Bn4pecbytBzm+AbQc47/xQK/QRC8EbtwXw3J
pOsRhcVeT1Jx0wQAaS2PVNqmA9/eI+Gk9iXfgUUB48iZHHEDplDJugJSh0U2
BAHsoJSgTq/gfqk1WWc0vrQOPVoHT/z63/pvUf5ekcnGjVlKXy1k4RJP6c3G
kOF9WPHmu3KVmDV/Iqtk6pkt1MT3jCCG8ZgxXo5BBrOk7TPotmRJz8AHkvSl
bxBlwocd3AMc6HwMv/NjXHf5VIT9feNl3TcZVzQzaEpOQLhtbxgy6QxQ8DeT
CoRsn9AFic6kLy6fd0b/l5OKZ3AZnpjbPmPUHYiYvXuicJVTDCVqD9Fy/F0J
3dzt4gWSarcnhzAGb6lwNzCET/My6Yk95OMoKBS4QMkXu17eROGK4k5qTWAo
vk3d3FMw7DkBSKlONP5qAmxJqRm13vMnD5rEBfM9Chbd2xMEShBTCcSb6/So
L33NWpPQOInl7speU2X/abPPeq/bQzGsIrIOeZjBz2f3o29ihY4siwr/mOjf
1SWyNNWOba/AmeU6wsfNZZ2bHOLwCZATY+Ky4F9ETJlbynsL+SkrmCJV3Jbu
ziroEHKvFwkKgYhVaSXAXQeW7DKm3ZdCfd5GK1FWw0JUnjW1bZfTuenQcTnk
BAc36XFKE0GL9Xo5O1ZtivgrrK/KKk2UsiaDWrkDdu2YnXJfZh1i50AmvzBe
3JbenLOy1mpoAKraHF3XrkDaiE341atBMZezxamHCophtskNoQEUjXIyP92p
zmbJ6Pl3Z0YSD/QbPwkiw6StCS247UohDsIHZSOGaqpbmwvmtKIZJR6k5MAg
sYtMCxcpEn50B0E8gXdl2jelGHJNDwOmYGoG6ZIxVjbIumQucH0LaW0cFEGd
4BnlX/drjyopzRQAhoRNLRGhxcDX+2pLEIqo7uXK3htz4W1VGPb0N8rXbNTe
/ekNt3C0vVRm/7rPQRuxdnFywMXJBkP4wMAo3ikWmr9qiTuAuhkNSFVwgHc9
A+Ye2WrBl3aCoyioBt5GjItCwxKNqga61p4X01gQ+jvgtEMFE4sMFL9eBqzA
kOX+2pMVjNaEEGGJfI3+pBBJOdBoKVrYZNicy0xvv8FD8ziXFGyc1luhe1RD
2RgwjrccWa0lzw3qEXKKL7yBQ0lynpY4EMj3k7V4B6qB+GRAxVh4HbVOdZmJ
WqzjxaZaC+c0yLUDIyUwkNdEJkb6J6Pb9y3DHeW5QvtkZYxySCoBQzUys+7E
4eERS16kyvGNP+EsYzurcAy2GqvWWughgvpKdblL1T1oqH+49Fnoq2F1b15G
C3d03t+PoyuJQeFpb3GVPnRMOBuefbZ4MCFSXvqGRzfks1DrFdnnl2SQmt9k
j6iaCyvdu3oHiyuKK6FTHMaOL2vAh7cPAcV7JCwZcobMOGiKpM+kmf2CGL+v
UaxXtYIAvSSPGOiueJTjtd8Mx2yq5JZpYHC2XdGHV7IsR6iEIg1SPG5NR+DK
GboS4+lWJePh3xwSqVsdM6kpjyIs+s1MQ+g1+z26QrnKvkRkM4qmufchBbmw
IA9OmU3mPuYs0WYP8r+3EP4PnqQvGLXVviGefe2DUPhbl6n+t1jyYuRnKQgZ
DTarPNF+vqQ0/olRbhPd3A98YwCI7Hyl7mmtxq98USutf5DN8wErowshwAzL
qhocE3+HbWLIr4KUy4q6G56cEhAshOLM0iIpmb42Y1CjO4nuomPlxSvlASfq
UCdVc182/RzHVttA5dAmo4ZGcnEyzUIcog/R9uMJ6ehTXOYt5doG2JDRRUCY
p6K14d5+dAz1LsQEHnaeibfL4Z1vD6ARRor1bb1JL5KocFjrsZgqvBkPq2ys
Kdc+/4k3Lb/9YTavurhhoZMRVZQGb5kxM9gz6sq3BtDrwEGXuQvGpm3T2L/o
RZ+btoqFalUESgcZL3lyRgSxgKIThTXUTBUfgnf3UTnCVighj2G2yGQth1ps
fInJG5FlOCvk9IDxV+0hmOkcnm94YsdvrtJi2v4C+duzDm6M71EUm8Dee2ci
/55lHdxBQes/sCvQPGOfo7Mblbx0/MkuGk+ZElKVzGvfZ6qoIN81SQAhUJDa
PyxtNKW4CwV5lhJUtLWRd8AB9Wz4Una/QF1bfNeOhfazZDObLT86I+bhWjjq
Cc97QqKjDV2dBkl1zZykhNPQHnfJprTJJ6AGLiKcSgKBBpOM0wE7a4Alku8E
1WjcBJKwIKgPpcKzTYVHXZgkcNKcKRLlkdeAD52gQaoEhOsyE9hnoy2Gm8AO
6JMqN4b2LuMpnFzh4XRpPM7jxv00Y7q0HJuwVkcfHVUyA0nb0jyzrMhknUkH
M0i/oE8NJCFOylc2vEDsIdlDT3x7swoUTeKMI4FYcddqibjj+utc4YsBaZGi
CyPsdmlaT4YPSRXzdVL4VLDZr+QHTp2oO5lLnx+Xr3OJAgoGaWtkEg2Ll7sq
ykruxB83HoFHrVmtixtz7Oj5oIA8LDw73HumzzhlLJtclIT0gbk9aJjU5jLM
yIA+sf8vhCyK1z4u5b6NIhbqVGJz2opduBjzL44uEqAvzVffW4R8QMkqYMbf
OhRCw8v0b4EWZ0KQvczh7l4BqyVWGyjVeD5y1CZl8Jwz4cehhDaeAL8g8Fl3
crzUF2mpDnS0UTWU5SIwFdGmhYVv+6LxM80srLy2PimZ8W1jKhq8dZCgRQ6D
4rNZQOsD7MpchiCNM6QhqQc7SoNqSruqdWr7enAQCKz9tsp+HyVqK8/XDID2
sheddAkx0CpL5yEC1z+AumtWRaZeDKsK7YKN+MJORukiTI0Q9rkpKYodZvyV
8r0DI8Mpojls4NoyQQsTL7+mDyc1tgv+D3pfCCavZXHCegqg/oXIU8IjwQaP
R56SXUKDIae4m86Cequ2adSq0fpLgPeUTCtRjhWHJ33AIXmaYDHqNq1/w9M/
umx0do5dSDZynKePco0NJET78wyu9P6be7GKVjNEBG6Jv/1uUARJ+SpHoPHu
1bl+mz5w8Mh8H7yujbwiavPTkofN1gpAZ6M7c/171uSBRFnTx2SIy8XGBpyp
0b3+W4xb1d7pY6Ckj08K5QZpxoLeRkjJk02ayzA7Ugc6CRB9w3//BRvsy2ns
3bSi0tmNy6zNIcWBVhGv+Rxpqjq3Ee9/GeYQEBDv6Qg9gpmR5/S/LGQYuVhr
9z22xkZJ9ERC7pMJ2vuq3YSTOpfUb4TVNFAcTgeyA3uj8/7vu3N4sJbCavdK
WVzqlm9H90CyIN4EbH+lLiBsndKk94+lDpoWSt4F2q9RXHrDCouwc7xfQzva
7ONR0eKxFji2PnQC6i12jYUUnpS0f6ldzy/mjeCxB2EwupZHlpiYRMG9CNxM
/s4QopP6dDgY/KLf+xeCsVJEu6swKby6ZMDDM6tu7Yj9bUtLZYDrk+67QZXe
VA92G2HpJ/FzXZ8OPwUXQGMJ/kE2d4SmY4DCNKq8Z+HrvCfVeX0aC8f/L63R
2+k15mmgd6Ofkycf8bkM5XouBnl+85+QbVmr0SLmM3LdvUm/O3etGgjjowWz
4Wb2zkqD6lFOUSDxo79SGsVvQwDmZsqyLebDFDAVIP/iA48fig/QZF4BFU0H
uh4CQfjvFeAtKrPtWL6DOC+ZXAM4SmTfHoGLWUFxT85TYdIFksAIRMTw4CKI
CnGjkjIB42TB7TPDDdJhnZTi+Hxz0wHDsfHsAYBn4jLzKGhCkhlO68jfscUy
a15JufeDKoUe1XapaQSrHBjd+ZIjaKn2zaFgroEvmaIAvwW9/rjWMRjxISKA
sOWxyfxknn9nssi0zpyu7PCO/0D2N0VsKz76u+6NQk9g6oqYvl43bigJJ1z5
iEk1jpx1bCiV+tgOvSAGxfNlgILBZZOwDMcS40NAzUV7K7vEPHIkagSaz5yi
iyEA805RVukNkV0HMFj01GFh6iVZXebNLQXNoL7eaNbsW0h9MwrSaag4ylcA
/tHVPIXJNtZwvlsFNbWgghJ6wzyXtIKJL7b120xDX/JVm4OX3XEfc5P2K18c
HityoHWNUHGxXjVXEl9ApSnAcWg6B/IaGj5UQxwVXdqHczgWQls0qwwHe1/0
cR3JMbDhv7gv+c/bunWpWw7ZW338VQJjIqYwW7Yyyp+I8WvMpLjZtN2XOAfU
w8bHMnmXLJ5bxHm0Hq2cFHXj4OZlnkyJDAPCX4wG1mMVsiSKtVesq+kL25tg
757TjVDc6yRA9mBxwMONlu5INgO4yNbHwSGRyAk0R/9Z+B3Zei2NAX5XUu9Z
u688vG2r5db3zo6I2BHvBEmfAVjG6xtFQLnf4zstxjoqaF4I/kTeOEnRDOLP
jvdNcOa5Y8jDQiZDUt9ZhuYI8u2MMvg9hnh33injZOE6pAoKE1jBClrx/2It
/C6VcRKXd05zNIsoILrqpbzx89KYp/GTsrxqnNNpjufVd9TKCopgp9YYjn3j
/0rguRrvzqy2jTJ0mPAfBg9a0+Wzos//S9/m95jb/l6NcNctFk1qz0BAFbVh
YYViPrh7Eq0Y3qn5o5voGA7kBJuc2nZHPBiZKYCyyQeZJfvb5i3hK+6Bh6Mq
bRK4PxNTEUxtm1yJkC4MRhzFT1OTVDF7Ba0PJxYhG2+6hjci5bbqHN8Q+M8H
smKyYofMiybgYeJZFQ3c2Ix/MTnhVgqMpk7gFLkecKse3lnDtz0ufCkcoc2d
jVQDxDqjZi4TyH7JVc+v54f6XUpbUu/dAU71zrgH7TlRuqy1Uj3gpeh5pW82
JGgyDs2vqAhOUh2oawW3Pdf6klFj9QQUazxYFkKILUdssvJTr4Z7oBj1f4H7
sWzHBPV1tHpbdZzj5HpGQKpsOttZs8YUhjLsk9z+1sY1Bh56oEfcdauokvIE
Wy54xt+9+ogeMu9tVF95MUkNnQY5Z+xSClOA+1L/Tbg/Aknj4+Nxyy612D93
RZydzY7ireTeZWtT8s1lSpUc+Cm5zCxGJAqfEFzgrzneuc3RsZlcBl/xKRVq
D9jv6QXZN9YxrRk0fi+cqiwlk0I9cTJdiSaehuGDIBrYmAPrLgOn02+AFexX
vWbEEPHqBq9omQqVjbdJgWTlp6jLGZXD+BO6c1fvuVjR5I6roatEEsl3PZUZ
6shsuWhdt5GH2Hv874vDkEiZdUROzY9xdyzp3ZhhN5BpN3vYo5CtCcNWO9jd
vF29yhf5IB01xYQqWzVj5COAXg02lOMkxViAWZ5D2Ww5uoFg9Xox5bm2NLV4
PsJmE1cs3O+wjeIU3ou7wwKcQ33kI3n8HOvqsI/N30a4N2DzRaADZ7Pan8bA
TAAQog+4b85YeMTab320H8H9IHFbtsUmWsvd9Hsbpnix98lBjSuDbUX0hWOC
o+GwkUFD54mPeqesPp/Y1ko+P4aSn8GHxFdfmGGrRNSUHCt4tkkj1iW6CPRa
Vt8eCtUwEqpKka9xljQsNGsk293aiyoRjDv+h36wHcFn5qrPrRzWCazz17jz
l7BWFga+sX1Q1U0fBkqOioFiWjprRvMs5fFkDjKkZ4H22OL/0rTLS3szmvsJ
9fcb0/v92xr/VehB+lnpMuWWGs7uJYUNF/KneMUMBScJQrt4v01zOdS0qn/6
X644uflxuQNAuMxnmf+87OnzPw+Sb2hL9MgE76Nf1ZR5FLpSBFFMnpghohMT
AU84pUa8TP0+dcZNBmnc5pA0hrjINSErUsns+Weu3BDBeXc+TZIZTPF4yfIm
jNq9dPwCuySOpiP/e6KilMes2OCIwDIw9pW7CtJgpgPIc+n6vkfnpUgC7+zj
3fuT6xafbHrovRCEGYZ2BtsW1k9d0qE1JX7bFp9d477LltgQDkVs22AAEWZL
owVEWX/bhLiW+XqCifLJ5beQjCFQjXuHMWFHT6CGcgo+sbQhVufvFtCkMaM9
/dqTVUyFwYKSdCPyxxdVT+KnafkUkq8AA/LUeLjyTznLTgpiJJ98RxseW/ir
/wdREiD2gjFu6A8ERkx2WA2pzlB8UsZ9JqcKfKdKuOrMu+PgZgKvJziCYxqD
fAAGf0ipG7fOfPva4WPyaeimBy5J05P+HbT6iAcz/J9mN+WIIFh/RB/KWfpP
LH1L9f/QRa/pswWs+b8MoEZcH9gQyH6N4STBFEJuNKFtdcyCEG8G5qcx37Au
Lh0KGBq2o6Br9/ji5fx/5V44M7PbEa4p/K1co3pONlOFl2a/xhcuY9xjER7L
Isa/lg2q9UGCdln4sZs7fwf1Rna4TQNMG+uhU6KGoXUrN0qaFKZ/bJeZAw8/
zeFlxuliYrukHD8xJiaDR89Njm+YDeYEQiC/HK8gHg6FBwFnlTps5TJkaiim
BFFIsEFKl+Q65i4c83xsSdOFgvcteTWlMqer892GDrdoks/M2ZN2uUiTcVgX
y1Rygu3V9lSf8wBEz6yjLIglXWzKwOliRtx6h0RgxpqZ4bnff5IyFNeSfAUO
TBsk0SJmmpP72o4aPkw2ODilyK+peiBOe233E64X7igXrAqPF9jQw77gPnQ6
box9XUlODo+LdUQ2J/PxWEtR0wDLqTRVdgrVYYq/NfOdWZipf8QuEEOfl4UT
vMMs9e7WVjJw6ZR6B8J9jZgA/XvzD7ERDVJhSByMJBw06KqDheXkFHZAsOTj
KGaxs5p9TbGg8uptPo8CVHUrPooC5yX/Kagvc7Iu99rIcx0vOBVC+n176AqS
TGyqPxc2yPpVBrLMW8xnpjg4cI2zdLRmD4ZrUwMIvC/Sbik9k+A7Yy1L4EOs
IyQdImAUsi+luGQH2k5/6OkVgz3RlAQe2Ked86NUWhuNQ1JJ4JHjJ8lRFPtF
JAsWHAgtsePKM2K7Xgq6iQZSzMdmVrWHgnvulrpjqyXZFAB3xKenVyYfHRAe
VYxCse5hR2g0Yc5tF8lvC9LiGRP663t0M2EynkMAtXYW39XooiRH7GnJzZZZ
isOAWZajOMn5gy19cyITN8jm2qZM9u9ashMB6SvTLqHsEymhYpQRTqgk12vA
7jdv2xHKDU39zvr3cCOWbGpSqvaE5C99lU6E6edTsKow269wfryL7ihAzpV+
HiL6W3+mr9MlWw1OpgqTxW8oZuDubpQb7ktOsR1h3CKEG5OmaYa7dulhnz+y
J7kU4SS/c3v4m+SFIHoEFp7wbiEVMTZ+V9AwkhY4pehEKc6bfkdU3bP7tSKc
MuP6e+yfwdTVrwNcT/hafKwnKE4/lPdQ05Tm5IV1Kz4GBfdTujDAf/ZsBjfm
05aJ0q7zOeWAWQN9zelYFbq5fiDeIh5WRmC+U3zF1CRX8r+0YXVjvyCJjsGr
GFHL3WP53Usx0rfAr0bEqXYnGSQeeu7C0ur4XAJARhzGO4zi4USr6gdCBris
jBqLYerNGOKhtxLcP3LguceineM03Zgjjh7sZu9v1cp+DAcO2Xs1mzCRJHhs
2q4GfBvnXyBxg0smkAponBN3a+/n9/+ndagrLIOl8JVVZuKoLXnqloZRO+SA
TEg3BSk45vSRU4hoeR3hT7S0aa9x1fUblj/666BV7VTxd2brwuRAD3b5Kqa8
pWipWbmoMMnfRmDCjx3vm4YKrKuL6A3gXXeIhVN2tybOxLY9+21/HMaOjwrA
mVejbDA5sHN/0rQyR/Ip0oioOCXj79igavcLR1BD6Da3hVcPbyIWD/YCRAjd
eIId7MrCiAfzhbYZh65Gz1g1Fo81XHmq+n7/Vh+Ww2QLyEs8y2nYwx1BE+dU
2+imE3OVWnNKRCgr2nW67jaPixPcIm8veE2zSD112tadfEluNReAoRBwu9Lb
hnr/06YT50W7bcDqH91r/25uYYCKBUtgrdSOkZzzRRkEXjdwrnhTpqVODIxQ
Q+KbCu6E5Q0jjN9iIaSzkcUKvPWu9kw79LEsZqx+tKzfiPwqhklJFZ07fXsM
nelM9O/r+qh0hJpI9DUkMYJm8C6X+5OfrmRROE4RtyoJSXWyHlBjm5zKtyns
jpi+F8W8t60ntuons5JFMmZciFPgmnUTIjuiJjvDEfOnot+Xq8z2D4fbERKn
pHcJKGHseAZYpDCfKIOfxirDn0ShskfFauIgO6g2qaLVmYemV8yNOH5MTk81
nhTpsvO3wZn1qk/y4za0bLiH2nJUlz5rFiH6kFwihKvpVEDlAPg9RcnJ+beC
a+MyktITUnwKnYoHT5B4q5RXTlMfHWwefMagS0ZBpAFvtoXP5Y1dnKyL8u8J
1TVZ0hopxGlkqVxNvvskglzZxmObduqIVj/518D60+vvOG4ApdR86h6ubsaR
ZXV/3zaowBdmOII3N2txD2CHUV2qEKyU4+AlmEk8NBXEi49+NS/bvOkNorh+
RE94GcvawhO8Ap8z6sRTRDe4+wE2frlG4OakXy90MuReoTuQGa4i+ZfVHNQy
ee4iOdNH00qBwtbeKnbIpx8BW0XHR0piyy3V0GWiQ6zxvmcbfKzX3Rr4wuQi
0x3QXVmYRa9w5iP8WpyrxV8q2uPaQW90ogH6N0PUhBCkD2luiLFBhN+r5z5t
oDUXFfHpbr+1vklWo4y2lt+KofxELkYh9bNvZnaoup5Z/TuEbZatteVZ2Eu4
3EaIRqE1iOvygtETsixma7zfyDTpHGJjOK7f7KdSHWrNjEkQpEHlXna92om6
ZLtSCDLYaO+l19qgy9hpOQsS8tY0bCZIflUVNGcLH+NIVg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Lz9FErDuMmu8jWDQsLyQXT6r8FZwsWk2Fd/mAmgIcurvlcGvG569DcCCmdb+Qj6wo3bQuZETQ7W61v4I8F7ezmCfqaK7MziJXUUuMTN30O8LxQQL0RNe52X/4lHITMYdachhIMsfAPKfwN8z/8XVRhPuVXVIUAC2Kn13l2rtU4gsjJdk2HYZxVnw+7pDy2iS3Ko+n9+e0WszdbNmqkFe5oRk4SrA3W57cW19i0Lu5fVb4za5F+zioeyHB5hhq+w3KTjPDrxSDHphYIf8+g9OdF/ndYACSRO0FEubvRTU/NZlxjY6qVC+X2PnloDz2FkN8YzzHBzkQBgqa3W3PeK65Rl3OXsueWzVRJfJv9kSs0uhyjTbnw0e4cFgqR+wcwVQwBb4Pn9YtUffFpfYF6ALwLF4H4WLe9xBvIx6Him1PKbeeW+kIQ7xfBL6Dj16EKCnvp24ki6N/NmiLLE+wGvpBybA83oypR6aTsn/H6ezVyWywOTbNgc3CP2iJGailHHfAqi7NR46RSg8MfnB2XIkCCEKrNEw8Y+9HDJ9cRGta1bhHUjXPTosSWS+P73qiQ9vNlCA+y70RQnVtYF8bXCyMfcgh9vqXFv3+z7tgw0AdZF4jLE35W2Ws1p5csZBQevcyeGtoaEjGUntgDzxGL/3fx80hI4AnhTpVT24kOftWYcWWZFvC846UyJbeeQCDeu08HocNeeBQM1VJhAi9/+2C5zvuHT56JxzDSex7cOBUXqfmYtikwQ1j9wzfmqjFddDDEiW8pX5tmw+bXihVxB68P"
`endif