// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SYzAB8D7q0LIeHciMnJuKmL0GaC5fZXGwvUnMrt93GZAYFDVvZ47fZQOSlQN
wzrNV2Rwp2dFxLsoknjJ7JjwFkDX/I2FpzfziAr393x5sbBL/7NpVsq8XpC7
7Top5KVkf0UcMUtGgGWGLgjymlIHZy8K5SA0AYpFw4YSIYgiS6TNUX9MdiU7
52154Kd2iD9qN6Ual1IgcO9gokPjv3f4viVjemPcz5fNX02KsNv6W2sMYrxk
SusVtcuLSKJHCusqUGHJq4yfUFtYyn5bG72Y83X0wb2HhbIxux6g/lKAv2Yx
WJKUyMDrXoQnP/VkUyWIUcah1Zmflzc/34rnWJZlYg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kj+FEaV+aAf6ZGiApdZ3g7/q082rZ5dFgpZifOmoxseKfPuZesE1nBlDxQ5m
LWkR6ZOb51743hQNjXMuznSwA8Pe5AxQf2wKtLpqW8ZlAZjKjKow1SYbCojp
IcAOGp4WoK8na3ZQGqNzpvCSijaiS2tz9Ln19UEDLysYwZF/A9CpDu1hr5i4
ju/xEI3qUDO7xp6CoAhUZbe9PX73OEbW4E4FZRolayp/kROSWYCzmRoK7XsT
zu7nZFcB1Acr8Q8tsbldskNjKlHt5RHWvJ+GOw7PtanIPDhVAjvVV6lhPD6v
oUFI6jfpIcXNcFK6YcL1i8yROWkFSI7qWE9qQFdAng==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HJQkMq9JFn4CFzd7IWwCUrDP3qrLYH8lBo57D6eDh6Qw4OUnf7mN5yPizZLv
iKwpShpoZC67W+rnjqRffi6iYKuFnPAbBsGR2vFXAHLkQLRJM7XMHWqv8MBF
CXcvrSHu3ZOhgH0Ld9rdTMcy64NeDwGkEXKrVBmu7PVgpG5Z/3l9lo7Hf4YM
3kxrlqjFINWDt2agzpmetsIClNVVn67g2wsnylvsJ9rvkdUWx6CVAML6nCPQ
VpNa4fYbuHFctwfK+XnDfr748/jd4EQBi46RdzY0AvMNeTd180C5PQPnTdCs
K+wteEnLPIPkepAfnlySaOsFq3YZt3TKjDt8Tan1GA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WBITPKBdzfovmIBGtxiZDpCOHMVracbjP/BkL1jmoFB6Njk0+GephDZKUU7T
z/cLzsqGX/xYEQDiUVEaGDSeUjx7wbpRuFG4Bl0jbX6voU/VGtWeo6Hec6R0
yUbpev58jCFoQ9wspCRz9Nhg3QNJvsNprAul9E1IEo6PCpB4OQ+jcqEMgmg4
GZP+2tj+PXtCt8Hsf0p3Crj3xTbAjKyleT7gtRCp5cjndeamJJ+Pk+3h2Zor
5xwxTZJPDjG7z7otrLcus3Zbs1F7ZhKswbpcCf9hwi2ldldNlSiiZ9d4UJ5V
prSUlity34w1ODz0n4fsyVGl8RSchLehmAfNVIy5vQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CjFlnSfCwUIHcl69SC6r1tgDNaxl00MaoJybiGNCVHk188m5A5VjqsJRlous
KXnsQxDvRx3R3bI13fJglyjkjRttz9OaCTbR+55fZwzKvmnlrIabeZ/wxmJh
k4BVpclPu9tJiAQf4dnwdzPEcDpuxkxe5F/Y1ry8EI8tdzyOKPU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kchHs3UdLYwCa3V83o3lm9g5DDvO2ux4eIltCCwoVq+cmReFpMh4qaogg1oK
0IIPt/NM/gtOcOWcDeD/gfjvjKtPSZYakMO4Fyese0j7bZ4IWhwDwSHpizJP
ky6z8uDeJ3Q3/yj47cXIjETAXhetiK6xIDFHzGvPWM3ty7hvNU4xww0Ly5qW
+zx9fFS7ppUHYtdVKMei/oohOGuE0jaDvSR+TahUx4FrdDH4jPV/Y4wyPFjn
EGUNpLJz97BSpS6NaC9hHHba4DuNmJWG5a3lFGi7jJ9k+KBoLjK18pUY5Cyo
0FGa74AnOslxtJrTcIZY/VixQSajYS3/O/m8wpIg9vAEZlPOQUVm/mdjJG9R
kpKX24oxjy8a5l8xB4p7vYpGN3qwzWQNRZ8HE/nlOXLQ9Zoaj4F1oTO49TuU
kAtoXpOC7MjqYh/2L44bYDdotatLnAgEf0BjWpdhCfi4X62FRJaG2q93LC0A
IATJA6t0Q0VKCAAcx57KPdWF/VGW/kte


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D8t4pRfaKn69LGwqiOAVp+adZnqfbx2qMEYYJlU1GLOsJQh2L3kxQgV4vQE3
BxkDuS2pvzjN2QJN/eOiprjK0yZSRmGOk6+4Zzdu2ncayqlKW1qqr+7cIPor
S0HBPMJTHdIYCVe1pRxnVWcGDNQocbhr7N3SxaEs3Oj9vR1LN0s=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XDxkeeE3oCAjA24YEEN1Ic6i17Fiha2/LPqwQlDgXOgzgpQbRtudkxzT0WMs
sHa/VD5y0L7nHs7WYSiTQgKyu1wDNsXaUE8BPc5TwijrmGpy54WmZOXG/XFS
J3VP1K9gcQgGOCsf2IjtLpyDYig0uWUJ8mrUlQ2bjVra74esvaI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 120464)
`pragma protect data_block
hqpceYEIW8LujoItwZ95qEDXNWEvv6kHX62iSvs9b6o5lteWpqUW0MUMm1Oj
BwV0+6IS4d/3TO+4OQBl2iKtddXF+8V0Z+OOnxzBG4759dx8VOMRG8yf05jm
Zy9XNmrLoGqFy4htwYO6ybLz2fdzjtbT0ltr3EIwTS31CjJWeu0l6x26qW7w
SbFNRQdQ9UJ1ofT3FW1dd8RP6gYO7ruXq+jkZCdNjUX34NnjMFP8wXe6uqY2
58rzaql+I5uGQQeN2QGTpGxWdGskbwtR9mFK6nzaebk/mRWSlr/rbUDyDWIy
RNqxD84bAuQVtiPfSDkP4GeDUVHru9XcD+W93o6oPwTg1enZmhT/jElzdVep
bq3cjliMAMxmRQOOgvV2amh+cAkoNqQ7Jb9EoS1IwqN+lRrWufmpZbOnOTbi
aP6PJLe3VQMX6Jl18tADUYVtMX/tellEirS2oe+gkwfyYV70qOzryEAeDac6
BiuoJ+sVxhOl8+tA5HPwEk4IXkhrzeCUjTOmQXsNg47MmJ97uTsBVEkG041V
21ryJWHDDiH6Gs16dGyQ5mgeIDwBVDHtNT12dWrnmxecAZwrVWIoe3r6pEnv
nkdh+9+146Q8FWNwCssfA6bgze5zr9V8PPmAJc0qi/aWkDlfcuFxn1GRZnEw
Z4uoBB/+mKfkNmOfjxXPSwLleq5SHHRBX3XJ1rKVspEoXQrbmaSLJB6hOxLT
JW4GJ9+4iQJmHfIIF3fii95inehH61xHTTqHLrpTQ0feDDyRL8HLb3RMD0tF
X6I65hFmnKvbFuuOVgt/0tecMRu7NydJokMjpG5gkG/FQI9yq9Z/lNsP/XU9
Pj/DaNet/0puydBksxidso1QkvzHokB1g5gQAfjvOcy2aBDEeK8U/0oIbO0y
lsxMK63+ajua/fCs82Ww/ulV0zPk3YAvVKxAHZwTHghj0IlJhDlnofIKLN9L
D20Q/+uaQ9hdzUPnmgsvwoEqmYSpZ/ZzzcG0m7ToPXBTmagdHw/tuQVc6Q21
pDy2j6XdxrErD6e2q6IlGs+3zh0lbRdKjRSPq4G/C33lmROpG/00qUvBuHM1
HKGK1+HvJ92+3lC8s1A9acUJXiGqAGy9EmVXDX0TKGQgTJDaZXXTAFIvtrCh
IuNU2H1mKfGCy3lPqWtLwwlupI7gFnB02jL6CDGDt3mBgaEmXHE+V0l0wAXU
epqX/q65vNOqNKm78BB9YL72cxodXQM9qe1lBlefvtgkUhU4F8Nm1WWfWef/
PO6rVpUaDpZj0SU5XdOogcWb5f+Rw70Wsan+Gn6S6Lygy4SmWpNd1MeSS251
kP+QRP1+JTgD+fX8kE4J+ZRFZ5fiWvaACurYCiY8MThKTfmy97BF8y2am/tt
dYe6C5fn0OZmoAyVVh1oM2UjpVtWTojBSlWJ/QNyc8a/jo5+ARckd+trHEki
lcGvIF09TVvj/Xwz+Jbbwbv8hWDagJEpsII2p8XUzWr3cMHPyhIY2gRErgqL
3bhba4kFREzAg7LnCU/776PbMoInAf+ZwTE9F7/AlcerX5NYq03UB4xxVrry
zpaQ210y8MRPj4jSRhuV3XuZXF9izHPFV1gWJ9n99QixQG3hWX2DHJPwucmv
ZyAGy7cqWjm2N79mGZxN1M5VWfQyP4DQDcxbotNWDDn+iVexXNqDUCZqT6vv
fozRyCAPh40Xj11p7GfwAbRW64jPAsg4QD6R5p/iBOKpPdINcMutAiA4IDpK
7NfooMOu5RddO7h8gPhTu7euzjeEN8rd8v+YWMUxJc/Nj7FIDNqlYspGzqbX
Ucip6ZHPFaFzikdU3mDpZVbYAFuvv+PzmL8Z23v9dhHHXRJAovxEGy+sxP3C
lcSlntveZ717ui0F41iFSeUXc5rAE9Vs1/ZM1Zv3prciNTDv0uNx9b1efIqQ
z+XVr+PFNGFf7ZS5+ibK0GdiilXWvolvFhQ9b5GwHT/qE9zE+/b6eJcTp+n1
KOmXPxTLOQ42RO2oFh8PLzgA1YvLZiFIfL7Tg5lB3lLp9ojRUjgn5GqafsZy
u0tU3s7IEr0YzeIXTd5vU6w2kPDz85xiGOdPmYXNCm630SnXHsFNHZ3/fV9p
UWBltBRh7M9ZF3SlSUAiMbHAm2q4IqbKC3mAjoOboKgUg34oswJM5BGd1Ji7
PpN2jCGF2sDdElKlk6HBRgmx4NBOi8wXtYayvwvIGI4c/q1BhX1GHSmXOmo6
1C+jc/mIK7X7cCBWsUwwPlOMNwwOalV78LHF7KpfOW6spTdiWqKIFEnxCwFO
P/9ssMINE9dpj/lAXrUCVpveF1bWjDnjl7jgU3koeWoeHyq2GwS4+cOALc1W
+pL1mK8NQOI3iia0IodeIWhxZVdOBVQqfUVXgic6ODYQv5sMZfqp6mloj7wb
82kSQMGHb73UKZyCYWP3M66s23APUxAlUevORw64FqRUFPpak4CR0ot0VSrv
o5PKMfOvvawX3VlAXX7vk+EUPglh5Jjy5LpQL8LyLNkJdx9eQNH5bjpInaZW
urFt6uEZ2q3dlqqoBoGe9gf70zrYudoSG/601UCd9LkmV4yUp8/DNbEbvozj
qMyAM7cw+Pl6TPLnOiB7Q5e8CRAhi+bzB4hagNwJH3P603HnEzD0fS89ixpt
4Oie9jwv1HzinCB6aB3gVyOemEphNvA86i3uaL5iYx0SzixA1enDCA67VjZf
st1COZ8FmaPKN+mngtiowfijftAzFF4sCufh+hKNrFG2kEvttebb4BpmUsvE
nNM54Fu/nFwJo3fVk8NChoq7AV3NlPEMah/aIbAJwDKsQ5jp5IvlEXskSqBu
vC06usRQKZX9aUdkQmS2/QPCZPgf9SANGtVr/Hw4rPYZtz5yIApJuFdFBBi+
nMIHZuEBUdoJPUD6V+eeCBuiTcpj/3wGW+gAEF8NWVzvPOas3dMO/Q9B/lAy
RuapjXjL76lNg09oh0DUy2anV08uupAECfj43gOUU1iD19hDxPOoLNzXtgoK
Tyq3DsoHVTDmV1KKKUso6blnyZsB513dt/DZfPiXNuVknmigxJGNxXZtKrhX
lLcfXHgFFemBWzlGB+IKhz2eUsZyzt74KKfVMqNgwddrFoQYZ7po5UQAbhAc
90hjNj9k3/TbOuu1l9PTB8IDHC8i2LAXlS7D1bcpwCqzhNN9srNVTZ3EZ1bf
sjK3znSrlQDPXhTSsp7Ok5pMc/lh+mXbuJjp69MYuhH/ifjphQ/47Qr8hwj8
dnI5n3cGpH2Av3uZRaN+VbVHpZHaeqv4R7YKDcBAkm3G9Q2Gy3cfk90U5Z3O
DLa2TLwwWcJHK3jdOvOMx9Mr1k6xT5iatXQortY8NrMllfmE96+1urffABRO
mmq1pxXV/coKCYnUd3fyfJceSgK9CqEzVg9UebCQ9IwYy8IjsfxcQKoX52Sk
X75ZP+7pFDVw8RNR2TDRUyDbovnNQ43SD73O2oGf6DJf4CYhVnFm0KCK4BHx
y5WzSLmcc7n/XCInaaLtnawxSQ0pnRfzUOkoyQboJBGSO9jB73mHuu3bdKP+
rPWyltgyZ+P7u//2Y2QTfODtJUHmPHu7vAfHNnqTPCJcVyGOX7pU8jij1kWK
YaSrpE+PSi4kUfsTQmkwLV4cWN3N5P96f/+V/bnRL+cq36rcNWgNRzxj8LI0
q7I8cv39Y5lnAg3iev99pl9Azn2KKUTcyuJ+Gr+vYAzxU0J3zPuSIBT+8Mps
pFMXh1oB4j6qMV6WpTJD7tIoJxbAndqE5dc9kHgmhOzfxd5Bu3HSH44PZOJ/
8o/NqXT54KCyBFI6b8T3bo/2ZiQsepltpOuGmOxkqJoOanCDHIduRm7rqfm8
S8qnCR/VqxWIaiYGPdslrhOwtXEqv6O9iZARLwy4YAQDYUgXnzy0QndPyty2
EvcH3aHJIwKLqXPUggO9BwcILkvlJiQdb857Lk+lhwHt6W0A5/c5bL1volmJ
NT/bwGDc1a7paxikMedhgnqqV26e0nIPvZ7zW7hER2p64Kl6ylMWcCW9ewUJ
Pukv+N64FBbzG7LlVmvVarWoQSQDMjex7UcRmgSH13E03Ekp9HglHLPLX3cB
Jn4uZRtB2gc2OXdClv1uh/9nH6ahj9LhFUKap44DuQzt9owN+C16lPxs3dtj
Alv5p3mImFPEtj5tPd/5iZcjIsslwAeOowanYhNlNFyJIvBG+s05530WH1iO
1MPmCVNBZDOegh6QMNHqEqSWydR1XtsKw/0LyiuhCBVK6fpOWtA7492CXS16
PiTr+MUWd1BZW2t6RPMFc3JJqMcAozg/Uh8VNd8Ny4ys+xVrGaEk6xVtkMLh
Le6wPm7JsyWfdztBVunEOw8Ed8fV10TyURrk6qdTqDjGz+IJ4tzPZ8zlKD7G
LKaZctM1Yh666R94u14KNZUDEDOzhCdvPDwi6x/wxnO9yvLSiMYXLEcNz4UF
rByaOgV+iLvnnCYuY/2EMc97d8A5jbDDfZwRrhs3Ru1WOSqbOg/p1RwRH8aj
I9r1RmbUCUHFPiuWborjTvZEVoPXsumFeiJ5yGGiBftXKUw4cK+haHkiGzR9
DQ4PO4og2hfz6oUXrZUJIdBJt0Qi2MsrbWSIEO31ttTSkckgY5ub/3y+VwFS
1Di5eHuEs5aUBO7ayN+9An3E5r/tGK4SzGJJlZ8auw1POt3M1PdtNgTkRm9j
+uYxb7lAqAcBK3JGnDOL49Km3kXK4vkfTo9CaBd30YdkcL5Ib8qZoSCc/grk
ek+Ea5iuQNIi2MO9UxJjLOExU+iyAj6iXjdtvS2qo5MtcgWWhVl6QBKv0aCS
JtzEZJsck1u7YeCSyhpx48fkMkzHrnLWr0aCH2/9ePs5sDvXcQe8AmmByURo
H1dp/QLcZpBChGAxmv15+l4SBNZka1otSqoaX6qHcPi+jfOMy3UyiiEunv41
o/or9y7Sw9J1hzF9CuO1WPK9OlAtRozvRnKsn37Cg56tB+MAOkjjLB/BHaX4
xd9MhmjlEAaaWZDW/o8ENQ6OSk29TA2MwlhyLhBZsGBy1F33C2MivzF6t/mC
Ug17fwEoOGNJ0KicZ5vf+8cXk8M1dygYR6fJOtqsWIRMqOhwZjyPSU9C8nhk
CcdrKbsvIY8B5CWVv8ntm4m2wS2F/Sn6SQbGZP7bypkIt28/Q6I7e0KpECUA
COgSsgjTAVL5XRMhE+DFkeFezjtKg71EatGAivlEM1hvWhtCQgd0tLzWmF6m
b9SgYzFMB5JZ/KtwXaOhf37T9xU6pegel0ITEV4myglggpr8SlIjg0pOA10k
5Sz/EbXvoF9xPs2ifftrF1PJbue+0HHK8WwTCMcCRS49v5TfJswHmtD2TLWL
Z4moJMgMemE+MPCQRae0khvBgHjVT4CvR4AgWQw/kZ5PRwW7bbnqbSBj3/7X
8WyDkOlcPqj042OtTXH70nDYoo9hJGpPLaYvw9ocHhxpg9u0KSOhk3iZIa3W
e4BOP+fBKByEtUqtp1SYdykiUthRpNbj1NBOT3vie2nOePwKXjKI+29GSyXi
of+B2tt+qdPMJbAlzbS3W+ExWgBJYMj663gbn9ar1tGygBVaSSn5Z3K5lXv7
gDaaNR7ogEZzVzUVB5V1Ax0LplvSlcgPD44tsmMHuaR1Ye2vP00y6lGHo4UH
mxtdxlD6JXtfxCLUv5AWIhfsnMFQpkClwI+XCdsdfU8jTDR/GqHZQBrb34Oy
m6TWPol0z1P+kQ5x8llKpMYmCIQU1QPQ4ffevkffXyWpLJ20ilm7iaHN8WmV
+eh0qtZz5RiAq/yZynRprb8WfmZFWiIL5UmfYmxC/DtGiBlKDOOE/plTUXLg
Z1wV6E3S3DOzSpFz4r9d8ZwMBLXxwF1ZQyxJ4KiGZZ8vcX7fKH8q0UpjLW5R
TsdK7chp5F0dXKwxXFYT2tq+vT30BltRc34W10U8qdm9pChInj1fGIUVYe51
PLGQLZcMdMsE82MrNjuFlqWiRKLGKjNOo7eOVL0yuDXiBLIGJQEBsfDtZZqw
tHVYm3hBSLLsq2qAw3yd7mpyxaIbKueqTp3q5E1BinD4ij56bitRDA69stjr
FxcuiVpgjSOVHpNAKCCrhmP4nEvr1gYkP7Mqw6fNKR5z+sZC9gSGR4RCIWws
gOYO8Euv+vzEsSOu/4owHhuXHAT8hIwAgubR8iexG3n1FGiLjgiKMxnE1gcm
DyPUuxF8mhUtR4IfUmzYODuaPY3G1Ri/Pwt4uerWnFtnh5vs6uyiaUG5nnrd
VzPFakJjQJ52v4PQY5MmxY2aj6pFlFmct5L9R2TkM85tGMChqCp11+D+/UEK
Ky5Gd7i50teXxDNdROk1PGkVPvJQ3AVi3hPjZd3g3vKOke3Ke3svPu6UTih1
jif5Xzwxk4fAAGT+ZshJFNkIo8sh81a4Cv+C+SRUK0o85Hc2uv8tPVKirZKm
IRHa4Eum8XWyzJQwLvUTGtOOP08Wl+dhdF2YMTdDVW9Ea6iwRUzjFT+JIPRR
vp9mpGcuGxO84PM+tp+hzfbShq+T92MI0Bs4ebZ6IvJcgP2ySX3i6Y5b4hBz
3uSd2x+oNPT0Emx8g5VIEgpv/MA5/5L4CI4eSqomvi3l+Nqtsa3h0qYAKhER
XMeRIjXZPpyKQUM+wBl3G8CwRnfqkpxbuBb4SwP530DySOmFJLC1oo8j9Ktd
q6NIVnUICHyp8HjExu1I6HFE2fSYo1V+iJgtD7s3RvNDshdHursAWNlTCHtW
iQ9cA78avbmlkpwGLjZyo7FAbTalnpOwmtEqO7qjTdPKnPWrYjo2MhjJmu9T
SSE0O/kow60Hc8N0OlBPNNiEZJlSAvYilF0YMcH9kw1TyikAE+r5ldkA0R0c
ksFL0cQCCLu/n8wRuKHXUFl0AH0+QZczaoQr9VSSdvwpmZlKpozwtNCHZTw4
mAlyzP0g9QdMVFqn3OqLhSMTOqdEDKDTYtdKfhVZR6/iq7sO0kXZwApDU/Pf
KfJ8eq8jiAaarXxd876ReCRrDEmuoO/3hyS4eQDtRQ0Z4tOGckQH2p+rCSlQ
tOiU4l/ZvBtbpFCVYEn0jtOYMySjr+zI0TtHmGbyP+/4UUVI6iHdSFUieyTc
OEvGI2WnmOrQma0VsGHFR+FxAtOLjsZka3AC9Y9EqweKZSL3BG6+17jbX/qG
NNDHnw3IyFaYZVW6TqSR7WH2SOm0dvAUozQ+VdH1M6J5uewzKtY6cXpbdIj0
IHc7JvDMxqHZogYdn1GGdT5Y/v0bcjfFJyJo162q4YafKpNj0SD8Vgvn1fnZ
2Ql8FvleGb5qsHSi57ybpgv1V+vUFYZUy3Co800c9zaM60igtHOK4WNvZcTY
xuT2D0+zCKKjSqitaabkurXSxZ9bfLBq+9yW5sngjc8/L51Aafibfe/yR1vR
as/EWFF6dp8qktlte24Ew6KIsiOAsq1W3KUOM6+SMCvHctfZISwKPj9s4DSz
xOWjnPBOtpAicO2Bjy0nOOO7NmHXDono0O/M80QKnxEv5qd4QgSDENTWBAxl
RibomFzFB2XKWWKPx3hUwt1kRUi3UwVfCI5z9eSML2zcgIeJ3Q2YsNM2uOJA
AGCm3NSFL1dLNa650d3bEqfoh8TdypSJ+qSU2K1/oUiPH586SqZLAFIY0hxO
Y/2w5gATP59Mb8FwKDD3dpue+sDt7M5qG6w+iVO/ds0clNRsLm1CpYAFFFDi
a5VPX9ddnDvRYYPI2BdEH+8g93+sI3Bckvz9AuPNE4WqLTjPmZAhqZLnSKCF
d3GJ4UWmqWeGrVxipqwSGmF0N8/R84WIxshiXQGshnnkq/IKEUCE5PFUeSka
HzaRych4KW+zVaGYMaEAxODuXWOWU19LOTWjJfUVymj/RqWxa7nn6KssfDpO
UQ7nSfhbHAxa14HJLmLp7d0ARXGcbVgXGUmyQpn+HTaCOd9ZyB2q4jBqtAIt
rD5MJLvB1mA+Xa1HYXAaJFluAOXBoGxN3usAL0eco3noZtLelAi+PshqVN5d
OFUUihbkVLc5kwn+GmZXsYdvie2lOvDRhmmXW1RW+DkCUtEWZ0ealxMfO9Ti
lbysY5HugVrxd5bYsy++lmYCpXTlzYmHGTJOeqYqXcx8xB3IprxQVPhSctx4
juhvGGCULvGuW7r5EfX0QnfRauvJHdicwm02VovTvX+4LA6y70j3dhogT2vK
4E1riMunWn1XLGzSoDOzt8mWNtMKN169jQPIkr7So7lnQsLisb5HOciNHBrV
5DGBAqnyxdD3bK2JMrTV7UZKvw4YD1RrzwupILJTd9JA30TvjXUcTPASe9UU
GUeJoOpvfS9DcCfTi4BZ7K7oyPikMQRGxg7O5cZMsq66lmgQ8oyst7OUzWZx
thBEc13lYWxBWK15GsjjpKa+F7jnGg7yn57vhZ3Gz3j/wIr8Dh6eBi3EGikS
fUp3R/5mRDWV/B+NAkuqFVaJbztC0pXoYay5l/7T8PEJvzgwUjl3dk/FNKja
mi/W4Q9MdoW9t4hEnYSsApLYboj+IEGyx3QLq5uAyIkkX6KBg4vxHwoBuFVx
ot0xdbFhTN6m4LJZIDQOFfZDsxgmC6Cx2Nyui83/XfKoVkIJqUwOvfKf6an4
BWOGv2tAmYr0tZ/EY1IwU+gVmgTf5hHoyDGzOjCLiBiLVVFYnTDXp/LIqhA+
XSOeG7yWKZMbhpdtJYW3/6JeJkF+cu+VkrHvzFCe5nBmgW7BgbTNt36l3B1X
f8kp85ZbXFuXwDxDpl0vslmzd068JuKl6qt+D+z6XM0MJi6h1FTa8DYQn2dy
gwEejqbM7ObeixuqvamEPMfskbFnRVemR3P/ruyZCtCL5d8jmSU84WYeejMo
9D5SxDWX7v2WECFpVvrjyb4z33qhQo6TKgW1r+nt56OCWpTYGCzq+nVMKoV0
g0VCKT5apjzBlxuwHJaJynzRN1TpKjIwkNZ8vP2IBZNwmTPLxcq0jb2DeKS7
7ko/iRt1F8hikMy1coZ62E/DCeyE3L+p4qeXRP5pjI0cSPeRdFt0L9FRSk5L
DgCpLIzotHb+1jYDvuWMwHrTmKXXAbmuDAIxKBqUnvRoEDbwgfwANblXz5IH
dZ+AurSzhzTjX4V2/fDzV14/azTkL+PJTJIJ8rQO+D0CJ6imuDKakPUkqB2H
ENumsPaWg5r3aUnH2OB9xeJoOmd1MK7TMBryOOeNuT7rrmW5SPeBRUw3Infg
BEfnSfSvpupw5TIBtzmCT69HPlFHja3DZUCyFVAtv44DR/eyBEmTU26RMXDE
VLwWjdrjGtysN9y7ptpYwcPvxwYuWnUZgFXrfiSD6NsmbGtpcQ5hJoGkubEz
ZxZswKV96Z0gdwtk0lpO2cMaeIc8F0/AUMWPhfDrMhmfMlLyr66DuWCaiOAq
yDFIXxF//yEVDzGYFVbO7+DR9oqEDVMgZDKFFhfxINwV6r3wjiVG5n+xcL2E
SEkC/6oY2xUFgCkvI/EaxPipPw/P9TJyl3cAuOfY2TH87V7gRAKb6NuHteTH
Am6qRts1OPAzQvwDFqfer/r+aWylRCvpvAh9pOMGXp0AdLeuoQfDV5ymMUod
SGoKayIZhTfHYvX6onvOl277XuTN8iMytXNKuHqfD5Vm21CyhMTy/EBQmi/9
5tGyPfd/3JwABYh0jn6b4PNGM9gMZZ978bh+Cz3gFLIO9M1MOkWsg4c//ryJ
FXpDyXGPXJUcIvGLzA4Jwmo0TXrLoSI4U6FZejs0rKtcin5FvZA37jbJnEfP
JAiE0JX8dWVMZYSrLnNmgjp2bblDf7nmYikO15JTZWdcZx8TUmCE+U38sD2X
HnIT7sbBSIxayIHgkIes1GOqICgtYRNkG9Lz6DVsIpLx9ARvaFxn3DoBgnRc
HWnv15Ze4euxvXhjQQZ1V7KEYDKSpkphAWWU/BYIzwGYWG9YlHXNJ/T3vRw2
+Wg9/jkEmii8mn87C1xqQpEPb7gF0G3/XRFPw/YZ/Mi3PJUFtYt8G5iiPlYO
AnHmw1uRYpoFxWv0n6NSmBJwomdZqdFqsSz2lOTaxNX68LDkdrw+Sc+uDau3
L/S39XduiPSwKAaAdhhHJX6S09T7anjcLPnoPFcR3enslMO7cdLA/pfWaUAd
IK8nBBFjUxjanc4LEfAnkjCan2zZUt8opzCXq9rYsQs+iUWu55GWMism5GXM
ZT9CYK3Ae8It58usnOuBrVeiVp9xwTwW00EVUyHOcbZxJA4VZDxSy6vPdyQ3
bagxr83/bXN48QYhXHNQsQrQmQxC9FedhJXnz4Gx6mPqmip4WGkOCxOOdqrH
KMHaoiR9mStp/8Ho4uJKBUNptOUsFCoXkLz/rF1CPMZk1ge0YjnN2VcqIwRo
cJfnZ80U92QKCyLS6R7VgUdq3rb46tbU3kbDMT1H5T/pKmmfZM8e28M11AmY
C30CAdMSUdgdugUoPGjVHc5swSX7qnwC3b4Kx/7/VmChfkxiw0FYSVWBCBkf
Or816bA8bxhyAKvtihLDXTpBnZAWKWifs1gtwEYESrkY+MmqKt5t0hxgeDm6
dEBSnq+rn7Ji61vx7NrJHBfDzQHNRjEL01iEb6CRqEbYmhIFGSzgYdd/mplJ
nr+Lc6D0Jk8tnldKaekOOOs4HHhasm3cESo2Nwsf9VoG/gZzUZLlp1JCNXmD
gnfagJirXKEjTsP6/YMW9KpSAzpE5cyhCQ34okYuG971XfFzSgJ1cvAbb5vH
YVX3mOnf7bIKZ5n8vmYvoEqP7QPpYKwnsjgQ2yjralGiL7BYXn+u5gEq3//6
6qT7Uko63YCZxUvHBi/q75v+2TWfF4fKomdGMnwUv4AEQN3QcFFk97fTZ+ph
ksbCRaSb06EvS3vj3KwnL3CX9QAPukTNF0JPUhO4Z47O6XRVjlCCbSfhFxTJ
VkiY7kye11/jRrZfAlp7a7kd48+A/q6vj9qfnDTxYCpv4LEPlPZFQuSs3LgK
y2QGNcfzFtDA2bThorFNv+3BIbhu8mscdnQu4h8CuTZH2XGdusocOC6nOjXo
MJ8goSfr6U6IGlqdeUBcSvo3ytGMYacj8aVsNF9bF5xHp/noPXBT/HN2MB6S
0KaFkltklZ6h/K+gFbQTLSrfemQYYfsqjy4kKdDufs8Vqv5vKHni7WKGQ5t9
qY6RlnwUwPvk2N7KsPdq04Jse8MWGkRfv+nqOUR7ULkrjgm23m7wDbvWixAs
/YVBUd9erzsQ64oc8JGOe0ku3ZiwKRghaP4Ynn72kNl1ze7Uuuvh3VgyOMRG
L96YZONwCZMid2dTRChJHT7Nf+3bKZZba0ktku/IyXL56oL7KMnFTsM+MgzZ
3kmKz5sVECMzhMHUHdyo7RGd7D6cH7iDxB4JWwlZ1vYJnxZjLq+Y2WlrSRdJ
BVznuO+64eqOxPLQQksUsKayqjQRl1Y7dPIkUqzSjIvY79BPKkZ1g98PD08p
RfTbzyDPhENPfqtU7+gfUiAKSh1XYCpxJwDdXPsDchqQ65PB/5A4jK71ah9h
+1RM8Dr5Rc65+zVMhR63JC9fcDUTkQMfocoLYJ5OUPi9CemVpzU7L3lvJNsP
bisCdDOPlX/RysG1p+C27V94dLO6/nzNjMQlyEm/y6e9J7xlBOwokMKQIzId
VQc+E3mOorFqJR1K9pZeshOALSS7gCEoqrjT6XPGaOMuLXTBsdWfhK/NpFxU
cc2kkiQwAesgDO0XDN6jd4odZIeHZRW/rgxDYdx4KmGbcxiLyepif5eWLF8v
xziK+G2JGf2/ZsyImdRiIhPdcv3E/kU/FBWlr6iSYgWIEWRSkJwttHgIBcWH
uyfGAoNmZSrbGb7GSelmPPpGHXAaf3bhF7lFP9hp2EovbBNdPLnqgeDaJAyn
OG0ZmysT8b1Pc1T9ftO3+Ba44oalcc1N13PQ/umyasZySozqi8+s5HVOFquC
oP4Hvix/gdBlH8tTEjjAg5uY/yivbRb2ch75yFJAiOez+brFx7bmqA7ds1og
opLBTOX19Xm6LP3J3xSdrNu88FKgbkaS0ffMf7BpVwnN391JdBEh6sfK5bNr
cfjQdfc7ukBuJ1trCSS4QgVTJ89+CWeVjBngXu3TK9D/KzOCW00RWlpIoOoq
76m5j6fUuQ6c/Vbq9Os42ZkLcDjlcCSPvb9gV5CcRrFC+5dz271np3CJmf69
BvrwXaPy0L/PX/vmXy96tBSBcrcDr6h2oNU4ck8nebp1vfJJ3si18uulSreX
UPPEsBr2ZZdTVsx+8lzd6X/05b5S8OQuqGvLpUgZr7k6EJHk7gdw/8M5y9YP
6+SAInbhSI3iQPYzhogpjmqBCsTxtqThsxmhX5jF4TWMyyJZ7XhakQSxQ4ft
aNnZIrrwFYnXJoEWJk8nUm8LChN+ANVVMYfU4eNhK9nU2d6hyivQn5my2nJD
um4IeDWMS6ywPwllfnKNhWTRjkmRk82/gbRz/G/BeIivl5dh0yHCtp141+7I
GwvCzzK9jiS1Zaw55xU651O07712XTdfPYQ4OB+iH0O/GrCUd5uXziiSTrxR
d/k7+vIreU1bdl1Vy82XDy7Z7N+roDq5MAFV7sm7wuxcBdJtdreTFffwJrbc
NHgtx7/dDMSjYUr2gISVrGJejUxOjU3rRnK4TdgIdbYb3ioOxAGkV+mTqKyG
M7UkSkAIXWkNMJ1QZ1tgXL1gniz+lC0/BdNumRVYzbqxAQqUuuAM9QEzAg0m
+07x9g/JGdzI/N/dbS1UoxBKFgcHVGVzVqYNaH2YnCfwjwmx92wCNopqqEo+
ZHvfl1GltEUNlHwR+eIUE18aqpGv5uVzje6R4QVhfFCQUDLxjfbB0OhkyOhq
fHH2sgokmhpllOVJhsaPw+yvdS7TievCqgm4jHi9CY88rP/Iy6MljpQjabKu
rLuCUfCWfuxO97f1fWdx5s5MymfeNnj/DyCBN/6/4h8ImJMA9z1q44st9qA+
P6eankRcF7KFwI06XwOmQtsfsV/wB+MMTgRSlkAeB8IWTz/wGSGtgVgyIvLh
5w3TJ66R5CiUwxbcbGnJ1PcAXcAnbU+PXSWIoXtu/lOsHsF3c5l4EWuXZv4n
YUd2HTps10xv83ayjMN7SOtC2UiCIbtivO/QeGt+4ZdA2uLyWQdvB+3080PC
fKrXxm66KVgCUjEJr1HlRmoPynx1J1Apymo7bcaiFcNYuGTgihAlWncfbYKg
i6SbxyYYrFOQ+MmUius2meJCKJyeSzU9PjKYnk6H9qVvyhdOwC2GG0vy4gtc
KPN70RNaj73S10iTnrq99Wz3ySrozutDz5vKRJ7492L+h4yfV3ORpbSm7stE
J5XS8kM/tcWbMavfy5AKO5mMxLAVb3UYS2mzTgtmisO0JbsZ6NiS2HHt0ywn
4fHhoIzIym2Gjf5rS0bZg4nYgrxcLPWxw3FZqBCeT1BkJZjAwMdGZqQqsHnp
1nCIW2y0ZrglUIb5kVawW78Zhe6VpTn0PmY1zYbcgvImIRFZsz+UuHrunnTM
irD1REgLzxiHztWn5dEuV3iVeOJ6l1yFRm20aWTfGa44RhXdiUf3XhZYTU/G
J5yqUVCbciyMsBU0IU2LhmfyrG2T/giM2SHFjpdBOnRUcYGx7oIZ/coiZmcu
CG7OVeOr4S2QrjCCkCP2aLOdeuW27Cw2KHW/Cpj8HwcxeIWw/GMhuVTYumtY
4fJ45dD4VZP2LgovUyZWGK5g4mPhCfo3OxFwnQWIfu7CKdQ/+lLxoKfat1w2
bMSF9Bm3JpiFsJ8o/QHlAxaFvKlJgMwc/LTLtUo9TmBZmfAW019W0/YSq3xU
4Jmguot+BmlpTuwCis3ppMDTbg0+/74vyrIMYZoUK9yMeABZv8FXvgtqpYJm
JeynawPQI8aolJnno4yjfuwQexOije6TePNLo9StSg/v1F+OtrAFwK3LfAJU
MBKI0WnJdCOA+92Ty/mqg91nkQX01wzBSpGUR0QL5jp3E6LEKs7TCY/WHssG
9ZwSSy2820PU8KaWHVPPvjMib5GBkrQw3DQZxtPG+mcf9grCZY+AI+0dfD+G
6a0/v9TMFqLmKuMDl5WtGwvJSR8FjllJF6X45llOy/MiH67zsExQhCy/Qfye
Dd1lE1caOjkivKHChK0NEYjZBJB0izCIeNTfyeHq6EC0cedTjJ+MI+uFJs9L
sApsrFaYKEigkOcPC5+XqXmOMY3lKP27UwlIl2b8KYex27l1HfjIPOZRKzH+
Ry9Uh9deaLGrTE+ou4ekHzqKyBTOMtF6s3ow7KLYrToXTk1AawUzzvSeOh8i
cOC76xPIJ3Pw5ia4+6ppgMqqFBAb6M67i+LniA+IELuIm043qBM4kOuobPpu
3ZctQucgcjFMq/6PZUtc2giA773ggFOzWeeaZsm5Sw3ZHBpgFv++29lseZff
roxdlTo+C+rcgONaOaJb/aEeluS+8xmJCpWw/gpLQFHOht5ifQFteB7zXc31
yqC+B840nt/1hNiXBx6JDA75rAwqV8VOVib4w4BqVYcPjUkCE6MEb9IfRakT
xjfc1YZI8chSml2fob+tNNteptqSZzZtU4PMBtYcriBQwbv8QGIuJUEyHiOU
vdcrGf2myAllA9RdIxyuEpeTlRdyYKTIPdG8bPz5h0avNu99ZTykE5H1xqxk
mcd6y45QdcN2mT/i7tjAeDhZFMogbn3bf0I7D7O6Cm3qqf8cFv0NcuYFEcSh
5j8A8E3v3F/U6oQjBkX3aMXxiZx0PaLuxI5lySkgehF3BylVlQppd8LYLerS
6ogdubp+KNilF3MO1xfbVIz2CGhG9RPZjLw1aZdK04xCPlbRcdcZUWAWx9dI
qiHnTifEw9Wkb+KQOJSSDcELbVHpsYgUKIyVzN9dUPpSMMiU3yBLhC98+j03
xiRVzIK8FmNLefXu0nxrrtSxm+bf2oHD5F2cL7Ly6i2y2tes5QrI0uOF5Nvg
Z7lkClBxJ+DpPbmp2KQ4gir2uCWG8YxTnX3rifh0QyN+kCZfKGdFov/yC5EN
BKhPQRo11bg2og++wFiWrnsNAOERk0keJdXdWwhFRkYkp6CGgio/xOIW4FUs
WrP2Vhg1y/HZOVxT5AnV11MITiwgrg9q6UI5YuD9qGVh0Kcui95seySKmc6E
0yMaCcCxCce82ogjJ7njIxd0hyIX9BlITl02nY/O26ObT5SbvLgh/XuK/Zcb
QTmztgAaADuoTce9lWt2bGHOqqyaluAsc09puHfgQIt45jYE3wKUBQLsyhYt
zklYowehT8qMV4thT1J4E8T8maOiGrkbBLbxLj6rMg2gTxTM5LHxBR4nur3c
nMMB0zCUtkqHmROshZqjR+J4WMcOKP3jkcOR7UenNWDN+C5g1peZJ9kFenG7
hS8LGvttR3cMlYsjAFyZI9ESylllCtuW5kO0ETwEQEQoQE2iDV6C0PmZ0sUH
pVbIGdnJAwMlCB2szVo3FRADfhRDpxUJz55b5X8oAXA4gGO8jdVSMC39h69k
NKBnXBpWIJKVsuNI2L+Kz2ClXfskx9UE8y0IUfxiSCdibv7XGltEDBKYni2S
KaqgrW5ib3bHlPH5bYPuLY6YiWT5dX5vaNJWfCyireDA6zW15ktJcqQHnvWu
NuS7Q3AKljc/P5D4DHhxhp2VVUAXpXAFeyPSuvK6hPY6HEf6w9xNInLhrUok
k99Ua7Gv0wNEI4viG3Cx5k96W83v67y3kBNhGj/0W8SOYW2sCMKnc420ThNP
I8+50MbZKKnrPLZF8VcHfYifzJXrtNmaqMrBo94LauPKR+L+m9FWuHmqRw4M
gHc4G1sC1FiymkJKYbkevUxaYFJXyopUVPBBbBdpUfDzNmKKhqu7dQjpL7iK
lO1+jFDH7IuLNOC2UMWATrSIQsVoYfGGU3jC0uU22XP8vBzr973zTUzRkCM+
auwqhqpU3PgEdIcYj39MWIRel/Rnk3TT5toJfkASQGH8Eg2l1Sr1dq4o6n26
qE7Yg0a2ZPA+zUViC25B31Ihsuo9CIlBtvYVC92ANrx7757r3Dr47lQ0+Lo3
RijOYpmYGmdbENSCsl/Ppo++V3KoF0dz6jEwSToFPBWvweK8+l5lmRE3oUKV
6ntf3PuHCT7Lijq/l44/n3nlMb6gwG9NE74v8wAe+5gov7HlR27nyP/QSEmA
hxKxicUnLdeYaVP99ruNFpdwFP0zMxcJMfKet6RpvjZV+JmdgLdZkqslFhlV
2j6FcGNlSGjXPRm//WZMB0FgInugLZ2On9ACoxs+WhdQUFRcRDVfqpQiP8UF
zH1/PIKIO+w2BdoIyuojTsDkR8xR0iorxeJYyrQAtN0SGNLFC1afz16S1AVW
GApX1ytA6QlPQEM6lpkdmWzwQ+Ak9U9ax42RjVAWz6tBj5Kx17/Xa/ACdOSf
zcDn58/jGucw187Yb/PQUULNZZx4dtBA6Aqo2QnjAzicKd4KOBvnt/tH+VmW
vNruGiNuaI58dse7PExfQxJqYv1Z//TVeYmRqjQIEd5a3g40LW81U0Ns1cYF
jmaG+PeZWYY03DZX3bsWh1//lopPOFzTpbZLWmkr5b5OtuyL/Wo36n6uf+fZ
yYp4RQiLzmIXaDSp3ls/5UI6CnJKPACdvXh4rvUb3Haj3VqYHbYEcJQpSpC/
X9X0eV9Z8ZkasEgBtqpW4GDmvFW/KI4lIS8GTkD1vQ1XUmww941+d69G8ugr
pgZBiwbw4bqPs7cDq5ExcdgzS57xhBZMvimNMf20Sf/K7h6kFqNX8Q7g0EMk
H5q7+9BgBf7rGhkT0kbxPZEVMygHVJpgqQ2cGLq54vS5nIksYBzOcsTh8HTy
iyse/LybLRFvsYUVqWVANJtnSnqR11BdtQSShipzwPU7bqg6QMDrQ0W4ghfM
IN2kQk8EOVRbdhZlS0v0hjHvO/lycgHl8dBN12syqzR+MF6iHtfG5fpiafRa
x3kKTbJAnMjQ09a2TE48Cyo2plTwQAEPCexxyCH6kxpamHPEPngk2ZCuaH/L
ETpHk2yL43Xx6yf4nHxk9ohitiS5pZ8Y9B0Ui3b2N/1lWJDUcsRUSjP7pV9w
mIQLRUbmtl27tWu/exTC/mAqioS+FQCLDnjGB0nXRi58W99OpNSlzrxHqwEH
sttkRdRl7A+SQpM2Pig9EINTCoVGk7IDKP5sxgoug9EFpsVgp1N3hF2eA07Z
AxgQfDSBq8+LzWVaXo2foU2zq0axCOU4lubChU5KdwRo9fpiK1NVKHOeuTIa
rVTPwcO3OpaFmqzo7ZcSr3H906pbDjka9aZcmF2YtrSrDI6dt0ZEo0MSAhHw
btV8SBebTcK0mUxlUWNOn/3nvwIaXPS8jK5Hjyn+DtBMJ+/Gkl4iJyZDcjGq
EEm6MKiixtUUTj8Lz9vbrRGBE/8++BBaTb+ZjhQ4bN1sGlNTpxB/8944cxEQ
HEJXP58oQsRpn/mOXTXfhkccoczxRFMEbYQ+g+emXbqJ1gdGnwgR8VChRNuY
bVg4YKd2I1Yw/yteU2UYZyy2KdzSxEdT9WHnUZ3a69hLuPXq03CxLmyyGpuU
4ToF3QVPDsfZ3p3k4hZYIhc1QEZLv8VsWn4vyWahp6nITDnAnPN2mZrglq0X
3g/FRAOwFiUWZ1tlj8NEOjDsFT1TG7nP/ohj+AUnxTBAPhfUigKsKHXil698
9yGpCn1mueVvWg3I7ahl2rLxErmWsZuhV1wfTl54CMWQF5wKnWls3ggCWELp
Ha8niuAuNfcvjucwcSubuDsFm36rxpMBQWx3zyf79HM+dLlz7oIh91XH5KB1
6mX24L4pr5Ma8Vz1xUp/jCavrAQoxyoOT8xzkMxT0BUt4M7/6ho7AzCbtwn9
JSxP1pbDa6xt8QYCOuNU3O8zMWbJgzNKTmBMPlhvKD1t14BX2XLLGcyrA05d
ynENdZ08YZHfKKrYgx/coduX3Y7NHKu9VjM8d6skWs5K9KmgMb/PBkfCtCA/
AIqDDXVXkP7lFQkXTCXGyS4Nlt2XZn1bcI+vT0eJxQpVuf5leugctMWDX2Od
61PJ3LL3p3aUNK8EXPFH/ScwO1YLVWDxH/1IPZHbu6VeG7harl+Pj31GblqQ
F8hnxEHS9fEiOLPoG4CAbCgPyY7MZ8t7yBN4NyfPa8Q6uOtUcV0A1etgfoG2
/qDRb+B3ssxYR02oC9Z8JefCnLA8ngE0e1zfjOr6LHZ5M3bKuN2vWA2dkHWR
ERU1XWA9ahfIWPqb2nvAmna0+KPmUBJTJ37aX5KCVcDXyHt+JC6TpctnwEvK
vtdE8glkHiC0uP2XjtJkX28AY3vum+cmOl5tXS+uv+BLI4bG2onYDbYBSfnI
gy6QwakwGN56X+9rhnIKNy2sMC6y9AlWtp5FSuLAJIoaBLrLD4LbbZEhj4rE
mtWC0XADweNi+PGVB2LgZw17639kIR0JjWuIPXSdoSKvMI4BtiVuUSpFTU1Y
1MCj2VWRqIbXn1UP6AFUZajDj9sEkMqH7k8JTEXkM1+EKLjS497I8NdEzUzQ
M49rNjN8jdt3/3piM/eQ3K6Ull3dNRlpe7Y7CpCU9cWZYZxtr+TbSEBIqbn1
BP+0tsIeCS4IFlO+VKxtQpIlUkQgnvo93Fnb7XSU8OLoSz9M2929JmhA2Qhm
YWXbTP8lt/5pVpQHJMImXT6VMIxR2TJVVFVcUVd6zwVJZ8MYokm3X7xijQTX
jXN7IuSUZtx4LY9nmWcx6u/s88C0yjxiwviTWaoYv5DI0yB5jJJ8WkRjKgsa
MPwqiAqRc/YyOgml+E2spak3Dx1q3y8a8jpmausJ+IRaHvpXvN6JTBIkYPMG
/abugE4bQYIFzbNeWpj6qs1gdIeyiFV3poQJ6KUVoZ0BYITbL5xJVXwjl9iO
yangOSWwoeW4RGQeoRXZO29kz9qaM2rxN2awc0cZZNDfp+V5kuOrURyPaM6j
uHFH2kG/EVwUPyvvOsdPSnTbPJkGc58tI8+JQevLu8N/Wm7qBrbMsyrfV2rp
vhN7vUhaLDpKBrLTEMEgwUGu5KQjaldBveFNFamTc7EbSkPII9799JZVQvTb
UrAavNp2miBCmpDy8V1VoIOoxDEZiUA9NASgvPrzND/tMH96W1vPzzrG+yHW
ORTiVs98grADgYw4W6k2ICHkQxLsGkjFZGf623jRGyOErtNwV1TkThwSj7Cu
496xPvekBYhylkwa+pM9DgYPaP0vrAqZft5jalXt+GZqmex89rcNn04qzF1i
raCT2YqRC+WPLM8wNxaRMXmwNOTUU32UHLAM+Z3/pXFwsspbKekExE+hGpVm
jeBalFYj2K8g3rsxcfYamONEGOZOsbAOVPm7DEJrsZzfRUwqsPZrZYhfQSwJ
mJnie56xWyV9JGzigzWFC9BFROPbkvGv07W6qC99F3YLcoyoN4MVBWrg0nd8
uUUWyIcEZdGj1/6lgUXty3/AAnHcvVF0agIEp+kuTCJybq7wcvVkuigRzo5q
ZsEOme0wvmEtuBYyW9dUtNPucOC4H/1+FnSoIdpMT272OrWDo8LBjQsveynA
40TyJkOa8M2pO4Qh1rG6AKa/zRHAcg80kQl/urhGMyhcwsYHYOMjpOrSdPJU
3ovnPjDc5M/JNWLLfusnmcL5+RiWegjj6TOzI4SCGMLSXHXDuJe/FsOHnQOC
DUXgmjNTfAQSl2nw+3ABmL4cZGL8X9OslKYcLBtaecZl36rr0IN7BX3zDs8N
dPm53rVo1N4YX2W3extzABVrqYO5pOC5ipHO6bPEzAGlkDjAdNOQ4C+2/HeO
tql7a1jfSYe+97rV/6zJn4NIvmf6OsAZl6CEf3nLRYwBDSyuX7Xrp0XMDyhs
huJspoGu2poLym0Vo0cwY3P92bSbK6n0gzGsDrkXRmEtpDkW5HPSbKkMmmY0
Z04oJrj9hEV/yFR/e4vJISQ6baZc1cq8K23UqkPPiPwxa5SXI0lzmGcX+ymy
VnQ+E63bLT8q+zvPQw55kHUv/xEVqocXBH+sXOPXD0zB5efBjHPwhN5H27aI
AUaNJBnZDF9/5WodOqEm5LZg0flRCd20LbPgB+yd1HzQIFmYKRAaMwWNt+7R
B6W5t9uuoyw3oQ8oYhoX6srVVsBeInlk5AGYw/DMCqSUWbgw4ZNI983pyqPo
WdQsjyehKb8aD/kdCAD1dP6lcXqCsN2IZIHb4V5hNcqm70S6AOyxVoRptzey
rtDvxCmCmhnRO8Ccn5IjregAGmWMN7oyrE7h/nbawbw5VCFjxNC9bizavHeX
tLrg1k7TmwYcZS4i2nFot+r3U9MnifnMoJiguDMnF975mFdk5HqwVQCEvXS7
93h2Q3o6ROx3BLhrvQ6rVlryvfCglllUEJYggjlcLzZALN1OG8dKR+TTLvm4
c5/JWoPTAGY1r6h98KFLKlsW/GZvaok+YP4tnN3ZFrhIXDQ2fb9xJF/z9CLx
p0vGtQaySB4J2rtX/Rg8FW47UAUUkrGjpQ6H+8X1vngqSQyAaqwTQKikE9Vm
eDuA281G4M2dIfPBPfZryfXq/GlyFy9zyxmlYEyxblUnq2gb6+w4q0tV8MIY
bf3VLMX3zLd+AfrZmCMxVNS3I84rYjboUtEshpw+e9cGyUU/IZGc3D3p43uk
J6sY6uSe4RFK47I+Gl6DzJUcDZmOe0rwfSVgp/+xvaYmzJCck8e1a9lbnybX
b27yyQkWSZFw1yJUin+VlEpyGVIaKk8Cpe0UhzxEEQslqdIboROu3/UI8EKD
+aYZWxK7dITzFMVBOeXK8SzuNzRBArReCaqTb4+Nq6SkzIaJF+LE/5VAiCl4
z2Tz8Bv3z9/Ts2VQZOHNAAyv+cDXGBhKzoe32KbRKYx+DnXJNvHlDxBObVL0
WzQobrE+xzn/KpvgoqSx9mjISf2tDUFxbpPnps/3PFtCfhvCuQ2sePM0sVgp
ffC9f7NOFWkn9PL/+hZyCOyiT8xT3nE/Y7HljX9j+TAu+YNUWQl09vWnQ20i
bI0uy9YLk5ZkBq7bMV9gP58bjnbd/dEVlLru42c+do9Q+NvGP4unOsesJFgi
1F6NFhUaVsiF1mS+SbqsZWsmW+nLSiZr9/VYMspgW+CGUzCjkLhz9BnKYxQN
jobPhIuZ+79AoUhoSCmhMyF2ksEX+op3a3dw/hZ1Nqb8LhJDsi9IKpvn+SIB
ssfLikZOxgb4y1yQcCbvKQ7q2Zdo4YZG98ipFDim21E/eKIjHPs5UXtJxiht
7p/vnk8qJyW5evknbYwJ3Bn17Za13CnTzY4YPzBCz80MGpGdtwbOSsoCI2/R
dI7koXQkGyVJegY8+LgehwvRKb8Az9POKVGrCZ052swTNCqLMfeO4aLO5la0
2r+oZtPev1KJ86qaUkgQliHLJ5RJLkV+RZ4dr4wq7ICUwl1iJ3RbTFIMZOOp
5/nuLZnTT2Ph1hqsbqZPvZnmBY51aC4kBhvbOUSN/rhbhpz84SMFO3eCYjea
bwWDChrjdNnJN4zPW3LT/9CZvDTgej3ntlVV/b6yzdhJ3Nxh7rD8rH2029kN
9yPlQlqMM2JFtTTg+i4KYfPVYJObsjhk/DuRI7uih43PgS6klXy9812QcHni
tkMycIJ9zknGnzApP81PdRabHlAPrJ3QFY1s+mxlF4cThkMLwPSB1LzthCFM
NkEu3/60F1ZxVyBh9tV6vlniZihO4097ZkCvjp2fBJFMRCRk/XOO/S7jRFgO
V6SrKfnyYxGJeykbTaWcT0Fmaqst0hlS1YyIkeVXll2uh73oBlad4ECV/Kqf
kxHzZThtE8VZEi2hJfxTnpkueOCyd6NIBu159UKlUSXuhojSenuj0Z3vNuDe
olw6Xd/mR2lHKb7JX26pq8cG6Y+LpbOZXVXyY2frHgmmH1C6Mr5FKN1Bgt1u
iPopIzEocEZWSjKv1US2f3aE8gV22p8AQxDhquOudIhvfylQSzHdZTRop9/V
tFD5yZEOViqmm+a6LV+zDdokKUVnZNDTtwt7zlMqanP9JMpgpzpup4MXsudJ
Pm1IuHnvp7Tqa2W5mrEU8ZRA+tAtZ52SiepCxYxILaQlNhUb1qxgCrKByEAX
j9Z/Pam8gs4YyUKwM+nxDFLShWnhLKMJrfauX3U93IL7uuOxmKvekc90vvfh
h3DYsLoVnwLT3s+Z7sstcTHWExDypb6/EBNOzkl5EFzU7PsiRLWcjn5ZSu5O
BgGqxoMezef7qVSLrq9pqPT/7nIdOC4FRWfEk0ra1KAh+LpfRYreaLc7DPNO
ZWwnzZIQxF6IgaPPHRYyOvI+yoPxWcizjP2Bp0ZD/hBWigumG2k5B4zTr135
21/yHZACx1wGfwO3lCrAQXT8K9g41Vssk4+7GCmwjLKY9/Nav5qV1ekf2wqt
3ygcZ4759hdaK1kEwQMlWYcQPvcAm0rFcnsZAf/dTcdgAYyolCmuiq2Q+FoJ
rSR0I04K9wBR66zn6RcrysBQR5OYb3laEY8V+fl8ac35gcSou2Osmovlj00Y
m1eP5rJWsdd+YbqrQKBu4oJw/rTotVuWTaq/h5p8dk4dpBcSZkafbtWYgJ0p
MHYlzrHC4zi+fmBvFQPt8AiIeXR+UD36PRyVBcTDrcKHnO6nlcMdI9A+ALLp
bhAVDz7xNww9cd7VB0Cqm6+7/q/1YbQi7uzdnpeRuVT8GdUg7syO4PgNwu0g
/nfhNcQeZOfyyFToWc4nMJnPc+OE3Lr7hePYGNi7sFRhl4qHM652vt5taMgO
KoPko1ffDFTquTuoexb8xd8S/JMD/gUImFtNK6eLp8wPFnjwzrmamD/76k3u
9pIeCoBl0LJ+eQ6zX4LUG7oXbw30ZABrFyowz58O9XcabkDzcTe1qwoJRrOT
cZbxdi+/PiQu4jDY4h30cZA5JB67YnT3Y8jSQ4t8ME64H9YS9FFaIb0j5ffX
CE5le5jAzOxyamjQj7ixPHEOHEjqUv6b3zgCFYddLDLt+T+/PGW6T4Q+b6ZW
sns8+A2mz8FiGVhVFMaBbmCSwj8pWkb0vkE6ArtoaegWkKDeOvomGKqHOvnJ
3wL+9corBlUcyUg20fc9vmbsAGthsWQI1mtR4pJfuWmji3bsXz+b/wdl+JYX
ziOSSpaNd+5qNYn6vgQnynLENEJdL4XuB8nzIo9NmG/ecmbCkGfBNVe51wK/
I/b1VBoit+60SdRV5wyS3E+b2cjiqBMDN4G2pdG6NCWGhDbj6qblJwILaMKq
AKwOd3Ma1jTd0JnNcmlNlltv22f2lHa0tyU4SdtFJoz/+oFWuf/VdZ062+/a
mIacJ2D34Q5XV5zZeLmbSSS7SudN9/cyuUAebRkzZ5tU01TSxroQU+fhhebk
rH0S87735yp5C2CQWtKHzaC7JkOR02SvPubWTa7lcc/jTQ6bMb+SEDQnkR/8
PYdkMHMZeSu6UodZu1PGIAMlA9IMcLBAzVXZtb0CEW+gw9Q7Rn4FCD1aGp7+
Xo8HSRgUVEpRHCl2ODGvznAT3lnHr18tv57LNs7tdk8b93YphqxYbYmpnehs
p4qSaPKEzBDY78hoXNEDh9rlRSJ+crQxGOswjQ904/3G5+YuxVJZxvEWXZU9
VfT2CVt9fHOnxk2PUNb0qzWC+saJ7VGtet8ynjcg8cteFzqCpfyRVwMEPlNO
HAN1PM7yqb5lf7wDUECs6am8pVYeKXD0R2G0KGirobd9mlY+THPNiSmyW4TH
0OIxyXjykAaqBwzymLnVHUJHyWiryBn2MfSNWbkJiN60jDweKBm21XR4ZfYk
AyeA1wEmpblOe/7b4Z9WuAeG5F6OeUEgYze8wp6n25YOoLthPGqoM1LuPx89
3lc3xvv09mEt+cjVlqKVmUTt76Ffjn/yRSafN0gzKdyrgZCZ1+WSE1rtJcoU
H8J+M2z8gAZMEqWem9pvJldYj4IPZnmlKKH5sPfHkBPZYnuDfJU2xnmNmaVE
0P53OxmpYJuHcmfLYY8V6kdmBoGw6DWfXE8Nc9kmeySwAk0xFsfKWtDjIaKs
QLfLokunSMghfqu2ZvdEBXY8rpO4Imm53DcdGva1pzVRYC/U3lxq8a077CGe
2jcYiZr/URYLuOTcwv+jk2tG8eSMzdRDFJRhnIaz4cUSe+V4GQf54YOrLDh5
pMndheCM9J2EHMC8HtZPqtnl82HVTF6fVzP1vNuZNn0Hj9Z2pLaTJBMEg2z4
LzrSJy9S7K19pMMmIRkXiEyMytBf5Y38gPtl3T6etQ//eKhp7Ajx8lSG8LC/
74Li0dVN6UopNlF7TkKf5X5hkTXbwlPh02aSydIWXSJWQidfA3kWRcQIZ3P+
31T+MHHWHGZbHCP/GDBgJRAC1GOt7Ym3v6+qbYbRq7pZTTlcY+U3B3IKfsEG
+2BUZaOqbtAtrkKb3bUtohoOZnd8fzDlL3jLWpeMBeuNDGjLscqPkiaslOlB
CIIlwq7/ECFpFLv0sFKyi4oXbeQrf/J2itHYc9pSvU6/QhzqANaj9TBz0dJl
y0jmfQS19Sy0Y+H2TO+JSIN4MG9scqP+hZqbWAaSLmP3Zq3oYpPWpQoG2HxC
4mrCYsush6aAfS4omgSQpOBCgAhr/9mO4fddatzLda4MzEbRP4WJyMzDPeZW
5eJTCEJXEqhxGi2YYG+RJ+ViGRtfiKJSrReKYKyl0kBt2wuvTKI1h7a7f3qw
JztDf7o91Z4aFkYvcLzGcnJ0p1TObT4AZ+bLUlXZpYtRCaCStBNFLdIbNIvG
eXMYD4qz4gZmBFwRVAyvkqDnx18UxjZZ9sDMS+td4skeQMiBKaxSavuGGxuy
NgOOqfbXzmCNNQLp2jmZG9YGErfmTchxqjZNxYAMtlNcr0VzbVqhdPrRcTJm
2WLZyUU6D8n0TB05b/aOJCtwi7vROIZwYoCk4LhvPE8H/QAPmA51r4mv9zR0
4+3wHlcb3rFqxYMcjZRG8gSdCi759Fp7z88PkEq8BnVrP8iTPf8qlKuVIA87
tUPkH1Fprij3KuheGfTdPP9RROWX1x7rd0A1h+XsCTfAfM0WO0pFvKs/s2HB
yz8YG0sngaImtFYVvILjDVxpzMD7BvhBUcHnhzWhCLCMby7izG26tf2h67uX
HhWVXPShjXuHMrDHdBT1Ki312Mfz6R1GGi916HYunA8gwo31TrFVjiqIHH2S
A138ltfM1VBjLCbPRi5+H6UDlayC8Ye7N7Z/IElAtvSiymNsLP7glt7vo/Wb
jAA1O7NgCsTMDduZeaXvo3K9pbE+OI9T5El2NJq6+XoZZc6Z56pdW1UYbR5b
b34E+/adcgf60w7XcilUL4h/mNtUX5gv2lGSSA2Fe6v6veb95NgdTRU7BaJ7
Gm9/aZio+FuXsfVCTqA36yIXYuUUnExGb0EyBQ+A+aXcafcEcW30rw1wXlbA
Ygw0vanYVwBiX//tsPasfeHmScoVL1lGRfopjdbANG5l2BFoAIj9OUz4894H
PrFhEg59sLwRg+/wI3UB6vZwHqOrkDPNW6P3iId/9dcXtJUSQu6aRO/uX3Jm
5sKA76gRx4KpqDKZJivAhffhjdqVAhqfc1X0Q/9m/w2pCCI7UkQrmB0p8WiX
trI75ZJv1zXhSo1hq1RXSU2Wagvap0ijMJQsuffRYoJymER1xetv8ZR39O1t
zSoXHfVamgrlK5x8x/hY5BVUNcqrs7LRaMZcpj0wLVX5IY4nQHKxKYu/vv3m
lxsBJaIjxdS8D3d9KmZ/rrvsjXnbkvqBnUbCcEpZipxGm+fGnYwPw2k+s06m
QdWYVj9DqOXEJkMPlKYdq2VUaKqWcasrc/W0PFGzwiKjbSC9hKhrIaX8nOkL
9XZbMyyfRibugaMxu93s+Y9XvLFOPhUbZFL5uUNgzdyufH7UopQlYeZ/w7Mq
/bjqAfa4fNKuU3hYOFXwvZcrU3j5XN4o1wgz12o66c30+M/uqcU8zxkJ4g0d
JEZjOdsR70LJIPryXyOMm3FHPxZKXK3wEI00NTFkw+opQRFU+Ws+LTTIzafv
2muJiyDJ7nkMiPvmqyXrmKoiJf6bQOXqoC3jXxPUX3tR32fXW8cSQA8N8p/r
uGghREX8OVcQBPuye2TmNlZ2sJ4MS7I2+Sw6wOTXz7+RJ2IQnl3BnWz62ba6
A76dYAesYWi/YaMw6n1WThQo1DxIJZa8/MSzUvFCDPGqGZK1DGUIQUWUJSu7
GF02lt0jGE6OMVPwP41WlNrIh54eoAByPpf9KluH+SzjLhea2oH12mxSSfQt
Cad6KpMaUU6ebBvxw5t4XxcxiKRht2BaIz3AhC4xT0foOe219DH62N+7EgK/
SNln03g/j5cuxWo8EyDLW31oq7Q/23zh8ZuOADuN1Raz6THuSayn7ipq+O/V
ggUlETMhS/FwA2IkB9O8tMQhVnPsntnBvPAK1DkZHcrgshCpHOw2/Yewmi2K
hwmP9CXigBp/27XjtY4FdeXTnRqVsy12IyAqQppmeBDY1s0uPFDrGHUWY5FX
6NRRUGEtFdspc8CgqmIXEaelWROEUEwIf78tDKDrb7mgENdNJ0MRV22VB94w
drtcjRNAjxh8+PHX/RH6op9g74jiR5/22bmcQVvfrfJfl+Tusvmk1DnOzbVI
jVtQBOUyuFZlOBUaQdSkO67F43CF2950fZqtG0E9IOPjzUWWh2MtQ037/pp3
XtCAtw5aMRyvc+p7loZBKmCPtBpIpG7BTZNrSvzsJ22JjGy5E9NQonruG5lV
AIQT/Oe5oXMR9IfjpeVPPYNidd3VHmwzg5olGBegjmZTPs3+sKEtbf+VC6IS
1cB/esqO75jZCqR/qqkiS5MRKsb6mam/AAdFd+LLKTF+oYihdU8UitWgYpum
hqGKPdt8aSWIUfpxzeozrriXwNetM8pBnUPlVDj1/1b7iH57akyvIeUmptUI
0HVl5gUvsMtjOvfhCtm6AIoa23VWytUtfEFyN9KG8xfLZwiGMCMibeyRYf2Z
zXFs14Tbc5tbcD25eeAf0VnejqSvJdDrAbFa3Y+z+qbv0Ksj7ixzl8XkieU8
kK8HTNYbZUyIOrprMYsMjiDY/dMEdC9vaDJGO9jOhJo1PcaPt/2Hj/s5YAfK
mU2QH/3mh2yb1ivNStAdkVI3EmAmTSXqmHosFm2GS9qwiZp9sS/LWYE3jok5
ATAcWRwfz8Zt+39kH7wOYDmiE3d15iaKaBe+wQHI6mkCUq7PRVc0ZcYKiYqM
GWC5VMCUqioTHd+lTeV2lkFbmg8/lTSWemIWlCIXQIYI8UTrMIG8oTd7LXcQ
6z3kJzFe6lEL4sqCnvIYpYWSVcDI5jSTFn1kMOX8lNSbCEJZgFdjOtCtGNGo
/6nJDVqL9xl3Uk98t2tasi2E4Nqy8AZTFTZe4XbnMpsTZM+OEvaA7VX1g9nx
6vQ2DU2vL/bdocrb+SX2KAChQP1XGeaFSwyhovT/u8VGUnVkg7Z4ZigMJTO+
ljtFEkyI2PyjyacB1EzUz3p+jng1bgIPkKawD70u3UnEmMx29/16fq3gnhCJ
Rf+hSoGpsZxu0W9/NiffIVIxK15t/G+tul13lk+XGIYm+clQXclpTzNgjy1l
hMI+ItmZmpvlPnExVta9Xx/wYe3dSvKIUfkNpwvnps9dzQ8acB5Fm+kN+v2K
DhUz5bioNwEsu57LKRpl5zNn0zw4UN5PhZEhIBeDfEi6Bk7f4za15XohNGFI
9fJBSbW89b6ArjT1iiCqrkDQmSD61RsiyunX4S69MsrprHSA2oD4Bp5o7bGw
JEv9xjUOh9VlEiLCB9jMpnd7S56y8+kKlZK5t3ROgb/JcW19poJy4Oq4P8/u
MRNan3SBRCSbHRcO2h+l99Rtj7YQvET6MPn5szDal4cV30L1fnoNyXI6r4nU
ftY0IMJCEgFNRo6Gcd7kXPtfyVZV71WleMHZ63oZwZaEZYDjpxQFCja/GAsp
RmkhJT1S5bSZ2/6nZ6i+p3ln4MXeVqq62PWM7aqB//S4pfmWPjHuzgrgGr+z
Iu9nDiQ762MA/XdHpy96qqF300uS/qFXg/BOksr0ci0Sr8KkCsyhaDft2RJG
gF2BSy78yiD/LFEtVjM4ns1y3mHLuikLUeHvgD+sho8CHnaoxxEuUs5rg92B
+tbwx803cNG6PR/fX5zn44zIdlR9KsdERctOZ2wN85YhC9TSHiSRRGpwAl8u
wtJuF5MJ75cJzPpCmo3NUZ1G+bqO+sPueXlbRBx9IdbASmKmUGHwuu9keLaJ
5b2BmI/bM+rhgQXjd4jN0o3QhU9ej6P2DsiVxgCu2/fJEFUkDlIa78eLWwJZ
tL4oAd5n+jLCHiXtKZPXYa27g0cswXQ07z4zn1qamhsFx/QyFRMnT8FbPUNs
BBVle8SPxc6HvxSqpRY4WM6twzBH/MIkMt0fxI2V4m7QKoO9+CKe41G/VW4c
7RK2nieOQq9r5TQBIeAzEPxXvLKT+TcdgvAKNGk2Yb3ZvrO0khJLYdotr1gk
F/MJJKx7JKQMcKEawqAhn16gP0iEjA6Ey7/FfdHwUDZ26ohizG87Pp6+Latj
Tj5BXqjrAoz1ZkV68SwVlnifYoQqqQIDfuj4KBk7eY46NZI0l2Bqp7p8wzqs
Ns44f6NtM1O35f1iKfGx0U9mlayTT5pbaIAVacOa6y/rbDRgQ+86RoFv4wOJ
7Zr6QIgVb56n0mGYjzbcuRuPjbHkM1fTf8fQ+7y4nmc5voXenQhQdJPZBMDO
YDeDPcoR/9V50NR7LcERJYKPRHoT5Qxu4LBCgTQgDGfpgR+ob4YFZk40cwZq
60O/CK7UiB+O6n9GCChfhGyrKfC/Du9uZfpZuhsWVXcfGICbOGHQTLO6C5Lz
naxLe8TWZrMiOi7TfLnBVZzeiGxPrnuTMC0XHgIeDvZ3mBPgfAhlyWxzgYWf
iWUBpKa+8MgKNBYIiztozR94iUaWlUEIoOvfQ0JgsBiyZ95wOW+DhKomHBlc
vEF08wxEVEjvumRJFpUs3bzhI+yoJGW/slZbOVcY1xhZGeC/LDU6he+V55Ob
vK9/oMYzv3c7LaVPawHhph9w9MNmuNq1ETbqzasKyH6RNKBK0WZvU30zYmDQ
CSn+8h6YHoj5pcpzf4zOXPWdw7z4XnFGo7og2U0+gTFdHSAlt8LLvto2qSdb
u5ne179K7sKd3Wi+X/2OWzAtP+tk1az+un6BkBXvMfmJ+eU1mFLv3xN1ZOyV
4rycKR6uq64RZ4tq6odx1R4/cPRPT2J6aLPnGPXZ92uF2gWBeFpAqTk71ipP
Qtb+FXm3SavRgQbHCY8OTqftDs7f7Zc/ahSBr44m4SbYOpmotNJAS72vlQrn
e8IBB+mUvDCib02N8dUfQPSQJh83iBjHEQD2yomcHzF8dzGXjnV6S37Jf9wM
MoXieAMyP/agJoMlT+EnYkfla5Fc9yS456yj1NPX+OLZEqQ6jfluQnIjShL4
YFYVIdDlhoP9jRiJCymyrd+Lb/C++L95XoC02w2+jbQnD6VdtIfd+1asbH0u
qYBHBqXA98vtjCCm68oNlQSk2NTpP0ZJCKV5tLnOc/+UQh0qP7QB6FjK/gcd
NskpgHo51w67zPcSQhwra6odD/iwDZPKL3myLV8YkYJ2s2Oe0SmVXEvXT0Xl
XO2faENYZVa2ka+si5YddP7fOv/FhL4vgf6zBJXdzM2xRokIObGGTwtVgHmJ
Ral0SY6KE0c/+lk7AWGJGNUm4zY5nGyCc7xr3+lKXPjDgHZoJQuXJG47hZOD
727JDSNkci1Gsa3F57xJU+JJ3Hgtd8yJdCR9/0F8uGpuDtW+VhfFWVlRkD2f
kzWdlDjz5OAdxErIW6mf2KpSpZdz+85fsZGOcJ6jyBWyuo0+7UOcmZeELhNJ
kca7N/kKU/KsFNo9dHDNrcfakAUWM+qIjyOrywpzUngB0AcxsoKDUUjZ9B8i
HxImt8aC/1f3xEfn/y7bizIgv7wDVM6tNIIpPr/H0CpC9kpfd/Xz/PV2lRsb
pNrU1kKHQ3UVoVgVS14Znle1dltp1AKL1mdwgJgULnmN0lyU0pDEt6h820OJ
0jyKO8i3srBesY5QRy3ase+usFgAsGxVuCmVT1AN8FedcsoE/7aEm27JL+hx
9A4tUR15olkoszIG3scCE1f/kIy0pcgbHy8q6aQiuacv64JFFebdiQ+XYnaE
8SSk+ZZ006qxrZaTTinaBxGVJB+XvuEE9CVaU5zz060x+CN/p/pUsyU7sdLd
UauZ3Uw4+8SPSAs79AqD8YAsQvH77ICsdJk2KthlrEbMQaH0gtOydUOl/k6X
WuH8aCTYGHwNV0cVJ9Sx5geAxo4xhfYxQ+1ELk3J2pwnCbrSRsX8h8rjnaLy
X8K22sZS8IXxIhJ+zjPf1FRoicIxPNLMjJK07i5VPwakk8HHj9KsVEGb7KU7
GSmv6v7hA9j9djcnBFHIfrcLAd7x58T1KeysvzPOp+Y+glTC913totjTAQtu
EoTBfqz2dHQPIwc3Sa5VOvjB2RYEYMsK+W9Fg3hLwutYwlYsaxe1p3X/iOP8
O9OmWCv62NFL8yhPmIU/aDo+dYSVPHeBpBS1Wl9j8aJpK2TRRsQDEIv3S7zj
SQXAbJCmUfcN2uwIgkAcGTRfURxm3IqxDxkDEEHhmUgK+chARQ2pcMq481tJ
170jyR7ghyqWOi2EUY9aJBEh5Cv6Z5SR9VDyRc1wdqxHDbJr49Ec7S+eIJV2
sfgo9yJ8lkR5HhGPp44QB16tGbSMJZgr+TuwpOZNqnOtxqy5V9yRKE7TunV7
UdOBZnzgp7V+jHWdDVKn5kpaWTeISx64LGFr3jDbn5sdqOHM0kaTESAEbY1U
xJa+JvC5NhqYHn5Xzm9lWimPxdxclBvRNFW/9Fg70cca+FY7jxSLJcGEmOMr
9ZgqPq0jt+ZZR3mlZJTuabclXhbLw4tTJ12CMO6th29y6K/Lzu1Qga2GOC9O
zr12JFKn0fJTggTFwqiO1sHl6miWLla7RF/sMxcZ/FP9KVG9vBxgYx/napBN
qbZYE+liyx4j1guPTxnIn6EwvA00aRi0OkFOc4MlcNtYGhhRbrYj9yzuFBr5
1aHhByjN38y9G26V3thuU6Jrd0GgELeGxsFps4T9Tyf++D7xWZ8fUQa/yJUl
ZPs21jmJ59+qAPYd9VCuOFy4bcJVAoK02ED/vdogbeBmGSERqdCvNaZI9L/U
n2eAW5NGRhUP6lTc7eEYNJaJ2kSDnKzdGcFN/QT0WcVXdcdDdtt+TtQs032m
R8Y54JxOjL1q+gv+SVKYQjxh76QzaU+z3Z/ECtJYolSk8jLNTN13YQcFpinJ
GRbV6a0blrQpm86yDXBjnEXXJ5I5tFl7sPoWIJAq73NTLHY+GjfrxmAqswYt
j2QpJDCgJjLahrapvfQzmOnRvjlWyFO53V9TP7qycXLvMVuV5GpZ7R6AnONJ
2bohAS/oJGedlBBLvSv+DCZAPm5LSHR02XKjwVeyfdPPhrtz/eyFr5nIIwEr
JrtybfyNYsiUcE2rYr5iphma1YbUT5k/412GUSlEcpN0d+oEJyYr2iYz7lD+
EJime/YDBjU7PNcVGKJy8Kdje3JUBtzX+/1HBdLRBeJa2HSzeWTX8HsHVlF5
wY3s7Yku/EqH6WEYjnKjAdFXuNrHlvg6kVVMBRI3UDlMlJ9DRkU5qhhNkyOe
Uc6Nh3DbxE9kdmQj+Wt2UBQmT/qYGnCiA0V1rcuHnQ4eIPnodSVARj/m76fy
gPHluf3/xlrpW2JBSxt0me/O1adrUrYwz5tT/8cgOorTZf3cJC1Zm+tKk2Aw
UzwMk2uMttjpcKVeqUGAByMM24jFAVDFthIshi3DgI7GMJ0pashJmwAFyt+s
1YCH+9jGzkYJEjTEjEm2UXUFyEVprk0q614VDnkTzuSzaYZIjGzn7fRvXLaW
sDdLwuXDwjNpTWziLLVeToQW5CtdmhrbaxW/Zz9JW1oaRgHKvwCsWmffZkj0
x6qSl/vWzTO04YBOt56TTpO8qNvkA0ZaD5ib1itaBLNC9QKeoARRWcGls/cK
DUr474KLwQXcqNdRHPpxkLYqwhTE3dNFUkkV2eNd9WhcrrX0G0EZIhYGhzMw
FYL9pZje4M0L8MS5vdkHv1AaraZpVM2sf0hN6g0NrLoJyWiE7IxCK7rM+yE3
lOBBwhynpCt5jaZI1cw6v566t6v6NaT/8RjtG0zDiDU5H3fhCCSTJ53dEB5M
Hra+G6Hzus7Ba0GzAjxkgtZfsiOt8i3WND1cztSri14dTiqgDxtom5qeanit
rlV7tc12+ntE8FEJP/dctV68KFl4/baFckOeK+5HoI8kHAtBbwsuk37DFsj7
Ma97g3EEjfhYn/lSBP2UR/vcSXnEhq6GmSJlV30vDC7LX5ewdRos0JpdZbIN
wNNgXEL9n/HOzwOFNR62uK7ekiCag58LGREjt1/xGm+EPARRUl4ikB/uP7Qi
jpU4P+OtmgrlxGA31tBrr9+bzmAScmkC5khRpANfh/2clQLNyAzxMd2s+esn
HIMiZVZXHDmDq/KsUrIcWXNAUIAA9H2dJgqtrZOACyVxdgLYjsTJh8K9hQ/B
NyuceZsZftDLzIgkxOZgv8zMd0iVTvUuxa5fnXElJ3eE83KShABDfDT0wppA
ZBUfmNDChP1VxJfYjCcOzib983+XqcQGjrOcCrGw0pSljQQ6h++N72MfqZvQ
C9Qq6X4u2LhqNXWcLDrgKszJnIodD6895xV2aj6lrNnCGZpmH5tsS5WczvLh
K/+6UHmZngLSfZBWVDpNky/mjoKkLyDswmeS8bsQ90P5pxtXsFC3zPOdKqUB
0KGTxtfGopUXr9rYVO08QA7RBj5wGVlo27BbvAWcH7Q8fSV0jvFGPbUeOdj3
blsUSgVpI45RJx/uYl+vEs+iFHJbLVDIlfWLYbBIoWYNVCexuFHvSwdkh6us
w8qw3Eb8PpPU5GdRCzpBWrPJE+bgU3kD+dvs/W6e09aMNNyQG9Xc1AeRU6me
TBRAI320JNJ6SLrgAyVpzhDYQNyh83RUtVgAIyIpoNGalDnnJfYHPIbFjYap
N9iG0waZk17aOvRc51wEO/qWjJpe3hdvwmDND+7V2legGrz91TjupqWi0aHU
eI/4QOdykkDVLF/m7HQiKLqa2Gw5VFfe6RD+6gv/UICoBkIctFYOguVgPh18
k99BGXeLW11gPlj/2ABCdHXsmIKtIxjf4pxw6ty3EakAGnHqTSu5w73G0iHH
iKpmuCNrrdSrDzGaQP4H/cWirN38A2mFv89FCOfmdodZfuPlOXnbBkhaz1ph
hulWOmLA6lLf6XDOfTGX1TJMQIjMe6okakZ2cYDUybQRCidNlGkYLI4edrlT
9eBelQQNkQKc/Xb9uWLptZpghwj1l/mgLxW3agW9yR1JFvhM/dSnpY8WZlwC
nwIf1LU0XWTRMD24T5AN53eQqMA9KnOJtSkqSO4hPq+OpG8hzLmlhOdCJbgE
oVUtwpATmYYHUQDDykNzEPWWOc0jiIqEK4oIsaw+qNqAcq8R4PumIt98Sw8P
vpfZXTyEYDykIx4EG7/CSWPFgs2b5fvA+gUloObKvfZiIPQjTgGEjzC/2l3P
3vFqhxiXQcn/tzV/cTvlztdSqopN5Wq1p4Ar1UrNKXcaOmmNRCqb7hfJA3Qe
4PHaDFYGLzUDn1HCSiooco/OZAc2Rxhv1l02SqRitIw+RE10FkROIGYfjMy5
Vvym6dM+EuKDiKHud5HgQLf9BhgqH5tXYMADIC2LHPtju+h94aOr66Y2/au6
7+6XTlIYjRLxFGP1kZ5Sgb5Pl2eGdLz1Csb8jrKEWiXh2N+C3w3NaodBOjOZ
T5HO14ZQ4+S8AaRiuwL8eDMUpQmvv1P2RzowkyTqHr74rXb65OEM76UitRBz
8bIC+hRDdC4tYUFVxLd3xegGyrCURIX6wVv6JLLcxk0E8clOpiboySqcADHr
OMLmunWLtTWpvgSstTMGEsnekSGkiJ/GDwi+Lp8rVb2iyy7WSou+JzxkT3Ua
mCHp18mQRVwMHlpeKdWS+xJv3DHkMMZaqp0tODymoeJy41dG8LKWGEBgRNJ5
k0OOsBDmos9Goz89upP4nIRTT0epIpkJZsuJpIC/lRdOSaz6yYVfhS/3Iinv
CtsW0sUtEcEVJF2Qz429ABtpJ2uP+BSQj8PfdpcFetn7IJbTDJMxpY0Us4ys
RdZSi/pbL/N4L7MHdEEVg2vTOlbAx/u34K/gBEyGKGqEQDtG1PDixzd2hhxq
PwtHQ4AsVYysIRPFebOBuCp7ITJYksCJLQAsiil38W2Dp1FXZProZjd1doiV
NdothiEViud2a/Bt6+kw7EqEUoYcsZElYnr+URqGyMjNtSqYUjsMn5mG0Pqq
FizV6zUFPCSAOx3HCPRmjkxqNfd80fN0CM/89supe9aYGSMsfF8rnKshTTAd
2yKvWL06sFhl3Tfsmv7NwRwyA2PqC9GtTY1tBIcU/FX9eHuK4BWEIILzvIh7
vE27LWr8N+3SnHIlbaaEJoiZuJgsSL+O73gpNqjX40zCXiHYUaD51IceHyA9
PKSVUMgxBcGrb5QBg+iOb2PdwfcpbcofU0eSXQWJN+frjquYzDcV+5zsmbES
UvCJynO/ZBcsVnWjUbd+5AYldb4cgLFyupaQkoGSDVXwhRLaaHjhod6ngxC2
s1VV56rgfwznbUHZwpyiSN+rOnjfPMVZqbXBEvWlzs1qnIQHkJ5GN7+WQMR0
E+TjAZvQxNtXl5hY4CZjbl+MVeLcr0aJnz8LpEiIInucu0F78eAq0EuBGxV5
kt5Gu6OIjwI2bTzVj3E5Y+UoD3Q64H4e5tNBtBd2Iu4f3Iunc3oFSPqH+AWH
3MwX+oK/Ymj4uer63ZH03KlwZeFC7khliw6uG/vkXz27DC74bguXXoqp1BDG
gA0xeP4oi7ZqAGcrPqXNScYud7931o/rQa377YIOq6Aspi0LZob6b8D5Fs1E
05wkCbdbJHJSbpgA2lZiibjkyisSEaemmIRTzhrvOYkaeo26IJT+MksAC5xo
OJ82cFvVJMy8JX6LRASj1+LYJ4azcd/wOi6HlqgzUN5LA9k75QABKB6yMWGe
X6G+ltHheL37hmH0mjVOYQ+hh5q+CZKXdYlEmo5X251ktcscmoRASzkPA6nF
NcEEx11ol9yXQvORFgHv24aquE3mxeqFr+lcpVY2Ai4RiraWnSLJa1tUwGEj
BDchnUVwMiqKPG2qgXIAUfqXZDowv1G5aWdEr/W8dgyTiAFU6PpZodcYRoj5
cOmx4s2u/PR7qCgOC95U4wt2HLePtUac9Dg6GofmqYZifhu2HFYKm8BbUgLN
4174bnjFLOjhP9tnZCNX11A/VgdADG0Ghj9OFEdMtzUcShP9FR5ehy0jg9Td
LueXlE5A3sw70K/aQBR8wx9ip4/39s1BysykbvUsyX5MUt35pZd97VZ/zzHU
hKAMuJ4adGbA6QAUFq3Lys2xrUfwJxPYfegtDXNiOTsnwx9J/DklhXWA8hu7
ccHxnbwLcJTtvTsSYANLg+KpBW9qj+APFN2xpOEWOBAbZD0nLqFYpJp7K9Kq
LQIWvwpHFRLGNXX16oxAZ2CVTYbjqyBLutoDBmYPEbhwjAUiVg902slXScWe
tPoY5yWtBuEWKCVYDEotJsKT81GM3+WqKcVte0W21vuD2DQ/TTlR5stn1Ih/
ncRw46Cn3lhcOmYflTNsbYb/yhQvHJEAXjoySekW9h09KfM6hM8K5WDNNqQq
1g6jeHtmB3oitkrw7DCtssUxODwKVd1ahmnqqsIqU1UY8RNX19zMz2v9d7KG
XIJCq7bappgtQ9mnN53+X0a0xB8FHRrQHqr7UcaLGFe/UgDLk0Idu3jXO2YL
lvheaPuYMr3wpFV12tPn2iv6mmvQyq2qlsXofGYU6hWVOPUrqH+W/lZLy10s
cej4G482oVC94UIbUsluhKT4AO83cLT30uw/zozJHfHbiB1DQI1DxXW69TDj
sjKwVxsfFu1z8EZY6HQJgVL8snt6nRkmgaKQa+O528GK4Hxj2YGjx98kxzZR
5ZbeFi6skqabVtbgwYi5Ad20UHkx/QjHdUoSkQs/YKOTKIgQA4VvstawyvAm
UobnZxcnYGkmorZCiy4qkyfX3duyFZ4uqZkqJwdamdtJI2isyyECnjQEjaFb
rXkUOd+ZJ/KbZcFUl1zDyMN32ZxXj3/9BHEYTFTIzdaoPnc60av9iG8ftMUg
Zp6Exk9RdMLzCXBhGRF4pcT5b1Z3bolRZO2TKCRcs6yAkHvps1rQ6s5KoE5J
84/fvURgWL6lhPlM9Qr1rH7c6wDb+f7OljVokL0vQVJ7sJRC8c0hrKwu9Hmi
V7GBipx/uHsRPIZX63vlcethgBPz0kr4Gs0ht0lgz6/bW4aSiFm6PMLB56wl
cMywND3YhhBOm2dt12dpclvuId7ApU43gle9vfmgDsmjlSwtGyJmrGKfrsr3
8lZmlzI8WJ5F5ze4PYaP5qCwWWinE2BkYqPbf3Gmz2fU9yZ9IS7Nb1wnuh4x
6SrvzceAxXLzrPP/dGV7AZ8ChguEbRWiPgxiVHlJ3av5fcTfPX8ghKvrcu3r
Fjcfpki3WW/IFaFNqCVM81jNrCg+6MO6ltI0VBw0EbbSdQzFA9YkpfZ3G6YP
j723Dukr2cu3cGamg7Uj9ol3pzyiAPheFvGSXWmKW2gkucujj9XICeuYPjp3
D8PBvzkIj3l6uI1oKwtD5TSda1GVd+vhVAYPZXIBRzOH3pikL/ZKnPFfMrWk
NlYTc6u6WwfS2teSgZ0crlRsJygpDrjCT57bNak1wmeIHTHflUErJT0iia/e
jY3Rv42WEGTO+HxsjHCIxkpHOsKG4hW5igakBRcxjlpT8YSGnWdQkqCrKbBY
zVTioGudHZCZJjNJ12hPxWVE38qKnLq+DC9V/bjz5Ykijwml6eRb5o8NqGxb
LtTJeLKyUQzJf0UrHp+Qh18FalPufRzaIZN1PzfsMTgF/41/R/eBjUmDfyZK
ytaphGMWMmjI216URtboBWTA2NCLuH4NdVLZBIUeQ65oyAVhbA9CiPl4N90n
QI7tqmAA98aVOdI4wKbV+6HbCsSl5DWOLtppd/g1VpYhbXjI8e/i8igHNeQe
ICNcEcU0x8syglbHZzBuDHR891Co0Eqnvq2YipfFfWO5qNIlX0cQE/UbyZ7I
Rccjk8pe66SsC9PPpXzHFr32fN0otEdfSTDv4/kSfCkuhpG6GTFSmXL7/uvD
UjpatpwWXs+d3mrD30t2sqGxQTto592b/Uq5v8OXFhuenmKfLpTSyi4KxVGq
HiCzvAjBbOtFR5IJ1qWm8aNy2gZDs5T94Qcn4chg5cyYmiee9dnEOUO3Li0t
kWbOoDU5lX+1PpeT9uG2mJm5cg/v/YlqDk0phIgR8EDET9Ilw7Iq+RTmGc+U
w8uQC74beNzsW5BcR5gvj29U8/uEIP0ps8D4jMWbx/rvLV4tjt7cQKEL8SUT
oPXT0lQLBet3Pd7oVRW9hldbzhW/C9Uq7GoWqZR1dijLeqoLcy/Sy4vypCx8
Tdg5MOnQQ1sf2eDH9LaBwl64oEg7O/RrxdmBtahwErB1/WGFJNsbHoVJJJY3
BVqZu0C6Orf+8BXivwlFr/QwJfErQnVWeU7MvJmN/cSaVk3/iiuZ/rvOR6+O
UXa3LPmDpSmy1z08csKpJkVWwehX5h+oEnGqUpbsAJe4oSFhM9OUrcF0UZIs
J/0cJOJJ0fOh1p48p3sThTOcqU5kkrMahlZDc60dyWQgLswYSJp84XWSDsue
7iW+qroH7AutRC4RVQM6Bc6dHRs+U3xL35BToZcTVpKwEeu/lRVGDMHU9Ein
qOVyIuTzFmRIkFG/mu6MqWnYoUfcnQiyCAsJFVwBZFpGsL0lUmumOexkRphc
LFHS7PTfP9WDneV3n8aGbyfMITgwl7ltIiM7yA4nirZakofpprMTl7o/HYB5
ci04QXvTRusNrzUi0TBJPtb315dnkqmfLbkU7ppBvN1H0kl9UODi2Y8FGeTy
1lMbzAhRV0LvWO0ujssuvTFwBuM9BvyYhyaZWI2tFaxKEPQkq6BqkBlZlCh8
fbZQcOb5QIu+HHGlOIbTyRIVjlngmj4opJeqI63kkF7M1XTJYHKf2JTtV47D
800GgY5gHP4UtyNTsSsro4FwjlNdK1+Ti9IaqyHY5HbJHbfp4xDD2fdKXqFJ
yjoi/g48ohnlQIvYfXoOtGdBRWrKqwjqO+LCRvw5V7uwz4nXliHoLSMOCqBc
lUUTsvX2QxR8OBeE3oi8l1S+KnITx0z+N9We3vqn9DNGnnOvjT0mQj53jFDW
ZIQfAw3oe/uDTQ/NCIKdAYdXOtwsVJypns01I2IdZCghiKg3UtuAWos2YPzu
ANI++gDTqmrJx7krxcU17MK3O9NM4zMBzJPwxw5gjXvSi7m6oIf2zHiKtW9Z
DDCPz2h5lTheLsllDsD3W7Mq1oRIjEk+eaUo4caCByBSLKQth0DWZ8RWuWPx
RzYcT13BQcfUH7lY3BTTS4t8qMieJd0alrftX30uMFZnblFfLrTRF/ez8AI5
pH4xO/Ps8KXwxdkyEjftUPBfpOL2fAhqc8+PJlPOcZ1DCbeqjFvac9Q0A8UX
GFbLW9xs5ArNHRHmCmiGkT10z5cooYR9NkZdSiijbfjMzYRBV3SqDyr99/br
cxdK3isZNNXINM4OqV/7kiGYdYSIwOKWxm4UnYK6AC3A/7UKEwpSwNQWk2d8
E5bDQJ+ci5uqHar0I7cY0+Qxge1k2DuNXQBLl1W6mfA7WNTus4KXTbro2fLe
yjy4iBWX4AGXVwv37ikMfH4WItxbEaSkNdV1BUfuFCWRADbRyzPcdaov4uUN
wPZxXO0mKlxtgsWDRdq4RoQ1k8qlwCSJblVinG4NAwDT+6ddPMunnh6i8jzo
Moq6ec3wWs5DeyjtDsjNgi2Zsi8I+CCmO02a2OMS969JmA8u2QhmMmnhT9ub
zy2WHuRFmwvFcg41KalbP25aiKq9CMLz6dj4IVKKVctKd+DPvYBn/iV2hCxe
9ANAXydZ5EDfxzA7p/kTh/PnNItCwWLBDgQuzAPG9MjPC4aEmuViCWbRUD9S
/VryoU/hQzhxxVXZw18a0L6cKBiWeQfJpcF1F6LDH2LyB4LgXU8+KO6WABy8
LyIkF6kDY4raS7eh6PC286/bXDFF28FIw6pG2UIlYZnVnXItTvA0WabR0pUA
ir7HLZFhaAsYCtnS0Ezx8jN+MdkFo+P4UFxla2Y9IkzUrCMWEV4KTFANdn97
nvReSfcppdg7NZxj6819J+1oVSEFyT/dprwBmpYg3uagi6mp4c6/C0MN0XGY
5PYX6l3DCnuvl5N3pcmMQQiAhdKP1/XzsXcnTnhEs78rjtdftgqlQ3+QFENZ
WELd1Xb9hAP0GsCkhF3e5EsGJrnKFZDUSOZxH2tUWstQBJbdPaxI6tTIH8hK
mw/yfJd2U5Hv+9XlgW8EQMSHAe2rEIPRSQRWw5k2VN+CgjaAI+P+rB1kTFg9
2YMRUodmTMUqmwW+UW+wOSHE+/FXhkPrLsln9Po/ZBeFwlNZKglEWmkyRnmE
P8ifbxODPh/WSpwih1jvRhK7u0nLAGMeJpOtunOpTrVGqSckP6Wyx5F5PEDg
RWn3Gf/tNJaAFFgKUx+Zn9HhExWu/7VP6SrGfmH8N/Nsk/rJwx17lPfYqdqS
Fxouql6ZutWfNfKKKpwNbHDKrUdH5Hbq6Sgk6DcZIei88UHyxhJHUTqo324q
FkGBHbmwJgET7t4/+tTayCefqWiaay5HGL0TQmCwoKn1KoyvopxRB987msyj
BvRmZUav7OuQrfkkNqRh4UmjIhbCKE+mVyHIYJ98i8DzZLpEzDD5HHT/E30z
+Oq/Pz6sR/zHL34g3BtTiGWifWvqoVXG/9B5lGfkQgNsDKgWYDrzoYfVCjb/
biPOuHwl530wm1jN49kP8KmPjzwNNA0pr4Jb1b8WBEzgNxFead0v2LXKH5fZ
wR36apTHZ93iIGCb9Kl9yNT5mjO3vr0jVUJvvMRPdDXBUO30Ii6mnrTAzYxm
OtW0JreFfro5YeYX3gLN86v3UG/ioGFY4v+5y6yOqj1A6RJxrD1d2oyS9KjZ
8i/8+EB1Q8elPebkpyKaitM8ySzkbff7nCMMwy16eWVM8kX1JoJRa9mBofJi
3rsviZ9riYpHQoZFfFWoKspYPXIbqv14Wb0kWiu2iF0TeXC176EL/4zy/6vc
qnmpdwZOx1AfVfEwMfA5FH/fzicHe9hsec9FPwmF325ouS2/3Q2Un6Sj8KOa
571NcHvcDLrt4RKWcgQbq82I1wbngf4Sps398J6/0n1Bsf4it0d0OqDh8Lwo
68uWJMYW/XHgIacvploemaNg+XDOcMgqJXDgEbyk3/jkf264WclT20SKJHUJ
LNB0r7B/TSHtri7csvaJhsUo/9HqnZ/k8om3GJ0ZqtlXnlBLo8ojB86EDTWX
UwshzlMTyhoToHzGGygPyFvAkhTA/07zo5GK168AcW3UtccNKilGia3uvcAh
seRXVjqGWePUj4wu6RHHYhwGFL3kMCvHaStLjCWjVq20L+nKS8Ih2e+g4d5A
JdSFwJA8gNNCdByO1mQ7P9/xniTXN5SljzY6zroUkrzoX+2VsujMdEGpRbq6
1kmnpfxqE2/B6sNvTQshGDBYPtHUAAQafw/e+ngOEpcekpqdZxE3fE5TZRn1
Tqxa/T9li3LR08JVUj0xcZWZTRMF9JnxqqUIoEjen6opccERsVJ47H/97xyk
IbeJeZiBnR2jQYPgacCKCeGkRHRUqLXRaCyART4M9/MpTAztL8l4De+TPKqA
lyeSz5uejzQHIozRj2SWh7oDsna6HBWiyrY6fv74N91NdsYumTPYh75WcsgG
8vKLTpIhLzw3lbzQAgLo12zwfLCCiU2YN/QTCuFoDT7CyHcAQLcdNd+tGAzx
SI2VZpO9xCef9pF1BW47+b8wQzFSD/Qm3Ej8cmptrBU/9dwVy9fEUtHeFrUq
ufNI9+mRYjH+ZF8sccMwyiBBcs4GrlS2e7oAoZgYkLsvDgqZT5nuVePrcAzu
ib9I1vUvKRiTy9HwxEKA4b/hOYKlkKNXZ0inAo5Y3KSxFzoPm9EQzq5jh+31
ZqnOLdurPrw40ZTKWu9BjPj4fDYitubFdJU0sHS8oAqjoKQz9MxE6m+wBjAF
mXEbQ309r0WeYXe2m1kQ6dhmTNWWAj8sp/loXz3lRoPVGSrfszlzYYDhDN/M
DMQyR3nAaGEdJs7jWdAADkqq1OZAZ2yIkNk/302j+L2DChYGro1zMH1SffmY
CiDCwJw1yEV1fVibqSw/URdoAdM9dqqA1wgIT1j4wZ0Y69WfFFwUTZEPGcrA
2uRkt0vb3HM4+DnWVTBZdNuIpCuolY7I9xLpg/ji4AezG+8CufO9MKp7Zf+C
23y1P5TyX1i2PtdZTQPEGTH+w21Ar6lP+ACA8KmpMGTEFyeh20YDX9JX9LaO
h4wOJ99bwLfLGLiZ2os0ogLkTBGAnnmgXIW0Ei6toeY9Zjlf2XUkW1sLMbdL
39/ehO9cO8ZQO+L8JtmJlG0JqL+IZcaWYfctKYoFZqv6r+3tNljlPs62f15w
a+0aZpcAawcFM23FLQS9qJin2nb4wvb0bPNlovZ3Z9q4/WzFeXue+jC+9i88
0lSRjomHCw98YXcjw+dY+IwW4s09QdvLY48E+PIkk8YcL/ASc261WT6ueY4R
LBC9B4fz09TunTVF7Dqci9V/f//q9rA/Tc1RsD1wVV4LBeDfGvW+beh2oNKR
zZTTbJV9t1xlHbMyaAWQQXUc+/zqN7NxsxKKafwBn+brGjDFseoKZcXpOBQO
b6NlmmFuk0RynyZMFLys3QH6/lOPSjdyoH3AkHLwnSbWLwrLVclloyLPv2Gk
hLItMC4sftWmaBqiFLmV4nsidtyRc55YYYtlx9AdoQnj3mtr4n4O0jzGFQNA
KuwIyP+v31LYzCdjoZ254p1EnSHFl4ahmn0k6VYg26JUL+HosSiRebatjMxu
DG21qNgo4h5KRZNEq1W1FDRNKdSQuI5kvDlbVT2yRZRvgv7nasVgSOoLRQZE
alVFpMEDNJiBcgvMPUhLjGGQl9GXxCulSECTy3va3TP9wO1oZk5DdWKP8NKB
yFhNk8m1rc1Rgqlb943FfiFzqWPrFXR0dklTNrrsCRyTwX+v+y11/kUfLy9/
LCIZv8MM4UCitDvLBW8gesZcSHWpO17fKkkEMK2mGCTls35GX/nbgUpXpVr2
jn66flOLxGMMKGV4/oZ03PjlaFojIrBoXPa8xvBeAAEB9Ezt71M9VWpdw0Ku
H9Hco5LYZhMK5c9iXFbI4q5HmJ6h3kPl/gJfiv3c5Avrc8jeoDgz4jfggES8
Al0P0uh99Z2A20VYw32Ig4XlWFdPtDppUBAHINAlGuiPWB4I8L0kN1r2gyJZ
YPw//u2vTlJjW9cpIRCT5Yn4Ske1XgubhuIBJUL9z3/RUZXj6bR0bSHAbhTA
7bEMWIpjdz1acIPV22P5gjW2SfPtZn0wADPg4jQiymal6qlIBhXy8JrcsMpd
/wRA+r8QPIzIUgKjAPB20AE2K9lNC+gvC3E6y7FiOU8VMASDtD90rdiWcbL/
6X+VMXkeDDKbl2ecpt5rNEKDRsr6t/UAD4GYjra79275Rr5DkhCk9p3GTKvH
9m2oSWuS6nQZRvK7xt5nnkM2YyQVlr0g/dh2DUiXKsZQLxjlj02P462npdiP
Pk3sTv7TC+I9Y+PV4B2ArdLMfiRPyd17kMeuuH9+TDPFhnYymsfFVKzfXsvz
ZFaH6e3GWJUkys+I9LPi5ezrwKhn55eFdDlVKVr4Hn3ZNcfR2rKAvj4OXslq
YxCFAbcJ1K4AXRpR434mlMfdjzFbIMB2G4zgA8xHinde/Fa+ybpGRCR7cSXY
7Vrv95wREKkm/LLHMKlt3AD0HoHUJ03p/iIOHHVsJlD0iJnEaW+wdD7FNla5
Y/UbZw055cr0h2BU47Ja300HgyEEQdP92op0CztZYsnSs5Ptq0z9QYzCifz4
+dIixAg2lWTQ0DwnfaRMnAlb82y/fZZrejPSBl8JigBedjKXxaIsX1VFcsPD
Ry5q6cglYtLoHiEgm56dScC5hnURzOyWu5Vy9mydg+6SU/xduy3KykklcEaj
ro1FD53NaFuVaLPreOl6Mxip1Megbb2MwDVIoitQ6HbwuTAtKXg81SZCTIbb
8IZA3pa0eKoJu2poUwFQ/uvxhe92zrLmS0LqMkKvjWG1RTS2jm7hh4mbiaFk
uUKp8IpbQGaWlfRC8WVHiGi8NMAo+swIe3m/VUHg85Mr+vQc6GuwhZ88dijt
oVHMUeRZVunl1E7KDig8f2wfefphMai0f8v+EdJvkJK8AMfKZXE47PTcfptx
eLjAjdLVRIE5MdZSDEu1mNbR+nglCIoviHUMTs7xIr79p2LqBSdmMtcn0hvL
7/KvXkdgVm6RIunI7j7LGqrpEy3o1kcsGyOWAtV4uf7wVYVPOb4Ua4ot/iMg
WZN+O5Odt9cMyvdnbLO9E/6pRTmE0ycGNgj8anXdQjBzbD6lBlb03utvtcGH
n2tRgAn3Dx6EiMp4+p11Z1gCj0eGdUanwvNrrBX95+UBKL61JGoZbE2m4E5s
Eo9zhbjYYcOpW5uQvVKdxCX5P785oE+MMeIY3OwfOlwWOtcGsXiPvryJHxQY
7gminjM0VKt2+AVxzYGKnESAWal5mZl3v+HFPGYOesmk2E7c2MEtiruoqwjs
VArMnVnaBDRzjN4Ub2kiQZX/bgfjKOMTr7V/YrOWZvA3BIP33eIapqeXZuhx
KZUEDa5rnV2ZG1CHmlxw1TZb13IGXXWFJjueSiX0G/zDjxoL8q4g/brUN2dt
8Mg0eWqfbKDemzhPnu32FU0oekX8E5h0aIIr6+maIxqfEYR9ikW7Fm6PWKHS
ZDsdRehYD9BC99zMNapBY5BSSMZKK+jod2bRhhx3wRUuQLHNtP5Wskj9x4LM
hL3GLaZNM1oq3fMmPiikpyAPN396pV0C3aKUkyG79QcFHkV1ls+QJm//AbD1
WQTNBvlANJE+kt9/M+giUgaamd86mL9XEXca9dBtfVZqSeBN+PANogkbRSuP
rID8i03ERxmMsANQhwsfaf8rWz50b3ASy9l3gW+eJ3N0FF6AhC/Q94zXJ+3H
GKiOV8/UCi2/2TyuVFvo4/IuH5z90Jp03ARaUQYwCKKVQrsKurZXt6gZTdaz
Now91TtaCE8SacZG1sQf8IAVNgZlx+xB63/cCrBBKEDWJRH0O8TROcKziCPq
95u0vZEGKqMTMmMKan8PjhLMUC1r+DSBBvvuBclqeekHshSMO/UubUurA9Q/
tg+mHjEc080htNBuqFH03UEQeL+SFVcXtMNHMTxHKaxEnyPRFvIMD2ROWFMO
Yf43L30cB7vggKLloU1I/9qmas1TJhhIMt58OpcHXnYgJLYCxzU7hqE0RFDC
2REXywNUchUuGalb780f74Gq9RmdAqtCppt3+CVpzLW+tpM9KuGYCX40MT68
qUEVDqZAvfr7T80z7HdekHpVLpZJCZtcVnRX9rnzc4/e3eP3M5tRXYGrIsJK
Qcbs7v98juP8FQ6FQ202H3rFvhNY0bhOttuv2pSqix/uMZTW0t5KKB+MIenL
KRACqhVW1lCcNbWpuaj9/zLa0ZJsABoxdrQBoBj8cdRL82hwcXUj4RSySf2w
RYBysKLr3yRWVVyuXJGHVuM2xVpTOUVL7JZyaRWgfE9NcmPn8n1NQTUgVDQp
b6FSWXn/+U+IJSxZkloI2FXB6Xzrg/OOHQclGNbSezOnnhSpVuHpnMEozhIF
+Cuk23MLV00eCnNjQ4tNVF3uHIp2XrmPABjsqEDC+PvAYSXQOMNberaNYQh/
3JDPZi/ZxX6WYxLRlPZgzxCXwFEV20t2lL1lH+M1FD77z0yJqxzt8hREA7LV
6mhg9GnJrgeOIX3Dtes50dqZgnO3XyVOJMnnxFsxrF9ej9FQQ4JL/vW0Nyqw
Y1nzRiJnP8zOtztibN4ESJy/VV0b1td5EfxPpBQ70CYpUyb1jDAboxopFe24
P6SiQExXfvHNedIsd+Y5vtb6GjBMpwWaEJk7A8EuPGRP1/vPDffI6O9ai86K
J4HLwcL5p9EckZu1zNeQfumDmjsprEGeqezLuNFcDgRUHNfE8gOyPsx4zcTk
AffACatnLIdUndUEdFBB1sKc4cPpVN3y3XYI9rI6X0uAJpcG1m7utO78rsgo
wQQox3Cku3yZUB+fUMvb80jqtP9GKNv725uDU8/AuhLP70jnxoLWkbo5FT8r
IQTo6bkU2+728qESgr8Z1Mczj4bUQZuMljyvvGhH+zG39mNwZYkmGIzPCMA1
cYRTeTtMps9BtEIP5zXv/wT4mfxjvsk5FTMx0hmjLjOOfLoAMP5IA0XFkXJP
kHDFJagsOj13Cn+1kvj6ZX8dVOABbQ7Itb4lxJtJgsuqP8EOR1EpCcystueZ
CTzNZABl4kdZTNKUOn3tTe/doJr11r+7eoS3DdFck5WxW6Ojf9VDYQtNfm8E
yf5g5f7+7eQfx1pi3jNdNMuwHBUvVGL6X/ZljQoGJSl0maOMq1njxb8/LjUD
RuYHwasC5TEYQT6gMjttaXjSPGOz5+ESB9NGgfvbXKhtQsHuISmtNQOIS/WZ
G4l7p9M1niPDXx2shFdFi9fvFCgEzjTW9oSAyrdiIQ+WzG/3NiXhBd7b5Eb1
2Wlxz35DKeTI3t4Z0zFfIb8SCrZQzAf9nR7cn4OWelFe2MHNmdRMdYGzz+Em
8Sm3k/B4iOy5lfq6XcPlDmULkyv51N/PePPORDrfHsU9WU5mjlq83uDpsiqH
6H/RyY7twGzCvQ28hpas3042sSkE7J1wOQhWOQPRPSYhxuyAtsnquiQXuY+B
T5muyyIN1gWW1z6r9wRElK2fXkiTPr0A0YA0Dd3kQO9uKttK0ZolQQZIIYoj
gPjoum+qV2iFgJwR7ecPlbmKWS36hit9lX5EZL0Fz6SqiRj5Bmk3QUv/RU+7
4CE1kFJkUostoWoF1HJ7hH/g6MRqCOh3CvSlyohitVHozw5QpaJBhciSHIqd
W6Jtnl+4lksFEIgi5EsMHIzI/elyqrr5+8V4oXq8bzBaHKdtYgiTwzmQCEC2
BNU4BJUsh+hO5tNdlRjJ6PT8TCxlQtyo4hIbe7c3asYonfknQeZhRU7xW3Hd
y+FQkV377hEDEV4kDIESXJlOca0lDzMeuExrbpeWExC3c42brot+eiUI2VmM
k1ngBk/137rFOC+MZJ2+PuV4s63Rqk4YyDmgZCDBnbziRFWoVdTddp/b7W6O
zZ0QHP7dVFVw8gKIo7P+niVTNqFOw5DBkLXkLO2FPOpc3iiAncQ4gd2elimR
cy3p99utResxGxk8mUacSMjRjG56WwPKN0YSVZpjyHlK2+1wExQgtwrCY5i4
tYfRbkxj9g0PO4nwDrq01k0y4PI5U265IhQ0aUdfC28NUMdrer7WHeWiBqih
+//i17qo+Hvd62YaEpeB9MkUM6KabfhD2AN3AR2ix8VGk1N+MswNrZIqmGN3
XtETbfd7VToh/wqNQp4kIJ8DleJS/VEJpoQ589q6cA/FzmV7NIqGdlDCZc1p
K5Ww4j8xJymY1jhJDMa0WrnzcmzAAhzmigUGaVqhRvrvtWu/tD0mCUIkME/M
x9/JmdkBUctDw8lRtc91ds4Vqi7B7evg3IdobUIBpBne8XaZ4K3XGmPmilCC
E0glHbqNd9sGrXDEG843G3idJ+FuG/u+ctwm3T/0NfPelRpoZvjLiDT1gXzF
rhx0rABbUzsi2IQbYj0XLuwerv4zKHMBeMV4RcpYx+8pLGqas9KjnyQuhrF8
+YBicWZz2/6KASMvFALtbRFEJJdiYCXniwqRVjBYyaLENIRUJpkpAZq6Ce5I
1wsNDsO0hH304TWoCTE5FGSwcvxBtIGe/d4g3M1M7fre8MUEmqdPRiyhG/dO
53xnC/TGSnD4DaaWtaQm81uKDweDF9pOSa4I5b+39xTgwdnZcMFmOEV5uP3A
Qda/+51DgXwaFYAKq1JjkjGI6LLtmW1EeU4lYrXtJ1VR2sBIjhJXBGFQZ1XM
0cBlH/7Dvq4QvamuBXzLeEUMWUHa1/BEUn97REUww4iQ/eJ/kSTBlO1eihAX
laFpU8UyX37DpliOkC2ZKBqMr3g6A0czFYSm6gg1nY/c0LYeCcXfCJfZwPXu
xMUgerwZEU0HpgQ4xxSXHclis+lFZ99FhOhiC2WuVoovBoLBWDWGlMiiHo3b
URhdFi7M/s9diyccn0BF7cwVBw3Dw+nf7oghI9YZyQ+0/U0VHmrLCxStoVo6
SwshUYihm4q8mDYcQzfpqH7A+6yvndoucnPCRrUyEPZOqJnuAhQn2Wuryp3m
Txe0RlUGk2er4Iw79KHx0AE1a8PUkQyWNnr4tVM02BKH4HHAzYtn8h+kZgQ5
oxlOKcp292QI8tJDxAdTz0zzolP93jmElb/Lca3ACk4c47yzRkoNmvEWmTOk
7ujXwTFTvvSFeK0/BLkN0vWFEFGN/pi3PTkP6BP0bQ6NaEBmfaR3srbKh1eq
+TZUGCaS5VHPAf1tVy0iUGi4VDhQpiQ1ZrZEqZd6N90WVDgiC2vBhYyrTxsZ
8Gm9cCV38gXpEHJY8oxVuWjzFfg+146wybhu9kVeNn7TODF08C6oBEX/HwvM
wruD651N3xG6Ky2J2k9yldOPgkowxJd5R4xGghQibtlvMlmazXBlio5T2xeg
zkD55/KOOsqVww6wh1zfHzkToa8o7h3GHGYUijQm7RuJ7yQk7XNrF7y+qOua
Nz4FC37mYdWlEflgHJ43ClyAr9cP6xCv0pUKxbwNEFAWvD4c3ydrQSzQAR2Y
61jI6T7Hmd2Bx6O9TxFucgvdd0zbigXkMpuF4wDiXDs0ovFrapWU/9FY612+
G1gAjR+yIfsMh2doZgIWIIXz73SCVyk9aqklH3CAnXmMPwxGBwygg+f+pA6L
TloSp3GApeysWBwe3IL9igEUZj9rG21pz8sLmmyx00QdqAxTXwmdwLRZYtGD
XEmeQdVWzkReVjgAdGLS1QnFNtd6mbdNF+d9guY7iQwO8Mv66UYUzDbcN1Rp
+04DcCDpXdsSGzcfedht19E5b8c59hIsdYNu1bXnVvoJvyhJWxt2l8241Mhx
/lUUXNgYNK4ZhY6uV5qD9qgEPZoYA+XvmdqEwov1wcS4RBA6mIfrMvbux2vu
vtoXt4tVIlsHT7jRL/Iqi5KfVr9FGFZwLleb29WVX0oO1r/QcVuQx1c0tFZ0
+1wxcZHJdU8PWk+V/LbaXQVtAf0lo0mcQnqkdmV6/f60rC6gf4f57L1o97Zg
ndGLNsTAb8h8h+aNs4dJBP6Fu/GslnDZ9G58GNSnMtTDHDQzL4y4ap8xmtOS
gq6KwmNTxowQB1T4klbL9wLBM4bTW4/ag/yICpqhkBSVftH/rGAGWUZzJM6e
WKWTEHo8W2O7Z0Ls3GXTfTpGvwpwU8hPcIWyPtg+Jw5Udr3jp5XuJ+Cse/5e
hArtGKDiyAWzC1uyn2B9vdKOcBxlMCBdWNR/YgkDwcHDZSSmqTXCUx/wkAw2
bD78pf9gh5U8B2ip/x6K3kZnhKL+5LCws/NZnAm5oQUTyhCjbgIRlOJ3BV1E
o3Crz9HsvJHHlB1CnLw1HrgFyvjCpA/1YXTovZLzzbxopCGjjBjz7PkMOlIM
ETchgtqC32wkz0vLaG4QdQbrLmd4A6si4j/NZyZQf9Xn6MFbryiSWU3UOtXO
ccmeQ4Qq2okgRxnOt4OGvEYI4N5Ziy1gPmef/NNyUPZ9DMwnALjEUrhZ/oUC
u6UsvppBlY3OlnSh2iBXdYy5gPYSm2GISRl39M08QThEZ3bH1OWAM7BEauVw
Hykv4Sv8d7XqpK+4KRWiff6DZVAXXWo6weUSGoytjJtq7ZX0dmwa2Kk+8h3x
qrazT7TBHNnLFFuFGiwvv4zj8MWI1RR7L0upv7f2OkRsqkYlLuDtYP1h6WHN
dcuyPXuM/0+TFep+nCmfdwSulg9EWsOtX5EIlCYwAAVz3WS+FItec7s2TT33
m3VsD9LXQc0pdGflJ86JS6DiOWRYOGVQ/0QgsWjuerIpbmyestL0nHZiW0WH
RmNVr7ZmAvtaGmkBCxRjf643p56va9tm6eqaO79XXfecTK7itfTaLyNGJ57f
wsmnsiX+qRMg0hxUj67UC+Clwlru1zWrW4IIWyW+6EuMJHtjQxD6Zmh10rcG
XjKyfnKUWEpbx/BQCvVLH5aXOjouVDpY6ayYBidj7e9lLNg9xU1orCkYWCsG
URZJ5HP7hKDjbLQnszqZekTEewMnXoXdsNBpRLyvE9yn2TZWQCiXHczcE9Px
iJHKvgdHjFM5gqKIQHWtqab0rX2jnVASHuzj+LgIHz4DZo1PqDeGsd5ntNyu
SOYgxleRsLgP2bO+Ulf60yi+ZbT7MPC8OlKFKp/mOg6ZhCjCFyFMK8kB+b4f
n8n5DED+Pu2w3NHYkW1Kvw18jOMHrI+DJfDiAK5jRzjvyjDeOiNy5FRHxww/
5dsZn8AQN4ZeQn1Mb6FLR7BZMcQvzXVB9MInO2MQcyJg4I0jtCIEVJhxVyip
zj3bqpJo2dYTeWh8bpsfTWwPq4mCl60A4LNClfmGPqvkqTBPVpKYm9cFawgo
f1cSpc4llZ7xCIT8BfE/rwj1azv7O4W58q4Frvj/DiBhFx2n/dIHyf/mQI7g
D01mnpfXa1fz2aDsARaHcS5eqr7S5dOBWfpPAlcSHi2A1EFtVo1P1M38r88v
KdQgChI+IyPCFDZ2eNHyqTiZlxSDc9pnoO42W/UfZmKl8EiGiJsxCVY/PQcT
DbYE9Fw0Dc/RWnVwC4SGV+O81AQ+xXir2331kfJkvS4cyyP0qSO+bs4TtOoi
FOOgEVgFC/4reutUsCKdlPtE2CpoqXqjqauFvcNyWXs/Sn7P0JrgPKAlrI1k
uSS2pkNcklBJd+829YW1bF7Ok+Ba4vWRbD3FAwFWhJln3KEztqhQhhPxJiFg
M/WblA0y9kfftOXsx2JfuG6fMuJaNwxDWlN80N0Z1FPH0x3eZHL1pV7f7USX
T5gBpCd5yPQ/cWlA+qPnMo3sp5t/3zmofHXIYRAWlr3HbGll/313O9TVtGft
/xN8XYPrqjMGM/26Lp/eDUJeOUkzQz9JC9TqZcV9+beuy61+7Y3LI9jjn28y
7yd1ZjeoMXkAKk+YOE4xmPj/iVjrGFHrqgJAgM7UlNs7P7GX7p0bkAeg5qkx
PM4xgqo1AjcTGyk7SZ2DdablheTc65yB2JA/FCh6zBlUNd93+CbYZnywK/oM
GmkeO4dDutnIbZrI7y4KNhvqdQ5fxyO/CGlBc+Wn9e97BPZPtcVb/+0qQQ2f
r2IYhLvSdkh0BWLqGL9XTRMJz90THju2zbz19fN3Nn7wd9d/zPsrvSKV+Epp
mIaWWUk+BEGqzBfzM6ny+GT/1dVfEleahD1myHTxulE1XuduFkRzeC3yBfZO
vCdkgb0huq4F7S5tOECH3giB86KVBMDbkZtLrss6EUG+/E4leYwjjzQCewg8
MNaIdOBibHFuc4hjXP+getAeStL9NpZc42slz23tgeKhEOpaHl7a+4vIjkYz
XSMdFdBQF9j5MLt3n5GAoiXBe6nqLox7lN+m3CTKSyeHR6UqZ0bD8f6XdbIS
Dl8Iedu7ApTQwdU64iEQdCcdNM50QkLEK/m0FUw8hS8Sq/y2tlECB0Fb20QG
7hwHS/gTtijspT0d9Xq7U4/f5GZYX3iNlgoe00nbgmhwuwe3TnTIxu0MvWo5
MziAS7PDabCoeqL9VhnFTd7c4rQOtCT65e2vV+6cHuzOfRWjQ5Kip9o1vi0t
xHsxlknZIUcPE7o+1V7jh0/XriBvzOX9e8EGRZ2s1+Bz+IfX6yWkEeiakpVh
2ia2yMcVoeNuxjDWv/oh55G79eDuMEnQjL5PqXsqPABGDyuC75CuTAOc0jao
VzSIW0cWDqzM2JOIRDFEj0cuGYvL9PmCGxJNl5WP9G5x+J5zPOR+XdrPFBUL
nbG2cc2PzPP8Kb25jqYadlbR66HicabNo7sEa03PwFXk6nozx9gjGmf5JBaF
JJjqFDHjZEirnPbgtzvRs6zCu4aEw3k+zYDPeIFDjb9NwGdY5AzzCFUqznJ5
wZAOU5YspY9S+gWy9wMeyrb9ERgbPx1j35aitF7yW7TBBD6Y5xaoqEwguS4F
e2QjFc9y3IKRtTBfMFt7dYxDtS2cnzCx652Rz817FxKSRuw+UAZ9UTxBbT+9
aO+BfsXj3IsmpxuCdlLadYFCHsY+ZqATkTlkW/Pkc+EbygSuMOZcKO/fWX6C
PbeVD10TQzD3kf8AjKut/PpnC3nrNKlJMqYyHJvIHANsyXCnLqWrKQ005kse
UcdwOZoggoVPyATLcc5UTqAOEDohYKBACMHeRkggw3RNVvGHigePmGe9RqSg
TQpxU0mJCfdTYwZALkYW7CdgWLsCYeK8Yq+mtMnMEwy1r0ScYa4CMIbQ99Tw
UUDTUYY3bGteNUb+pqoa+HyHI47vFl1JIPScL98dI95RRV9sN2HDLTnr/cjn
PWTB+UnacEmwLWxQQ+D8+7uMIShwxWWzLnj9uL2naDeVvfbz+VA+xONvUCjF
cH9/StZsOuty4SKKBydP8ak+MgkKEdu7nXs982w98Qmy6YOX+vur218xdQHr
pr7ZTV120290T3GofAEdYmXuFLOicfZFn6Zs1CcyWfJL0Oi91/P5ZIcRWPIs
oSy9WJSVze+zQE0AOw1uTtX/2Ga9a0UhhZV89UkAV5kLeIY9Vqn6W9YAu8eI
w6FsfXFeCUUtyKH96YhnPoN7NjKojSlpKK84P/lTojKa1CdclvYasfat0ZjK
Air7QRBu/3PL7+Lm+Ot5zGNxoXnistmkl6NsB82FNDW9ADJUWOMgStHfdbTs
7hWY1nt7DTt+6z9CBcKSg/kDk0NsMx05q8cPWdQ+hJxDC31ZIEG6H7R1HZl3
BKjruZyPWN9a9rF3sLneWJ+A5Me5k0X8gL6dD9nDFDlNyVQMptnfb4mXpGh5
sC+pmROA++RY/b2FQgGjRWGESFIpxSuC5n0k5OpswVIJb+UYMyOpJigd5npt
kRupQErD9/m+R2NmMwKirDLb0b5n2PhFF+tMO9HzVMwxk2Yi/MbloCFTUHeW
3o80LmH4mtL8LjrKp1Mno4TulgamPf0k3Vl+5Eh5FtJmgrtY6yL1jbpSQrvy
4JnboqPTmWLR91TVBCfsq0rR+XS3HsBzmaw0BtW0FkA62n3OH4DYyLZI/6yz
oVBCDaCtmexNOfcxpDs+Sth+gJIaRE8/XOk+V7vc7jL2CWtVIbJcJ1W0zgQx
p8ZsnxcKt2JL4uIOyUmYAgDv+a5feuEiRzjGotoM8xilZl4ek3mmsflL1BAP
/jLVhjxjtOtpFxcA1S4GURGGxXCNJ1sp7pB6YWfs7AQhv6+6RpJjwINz/wxx
F08n1GDk6UQpSpEQXkHNys7KPMfZpBYw5ipcKosn+Tb84N3fWrX8kQr1gtvv
LMmi9agJV1Ldh/peW8diSvk0YzlqQejupAstsqvi3dmV2gPkiQMrN0mQEi3W
m/4yD7esYtxdHraFKiJ3s5SbF6vlSLZgyl8WqQiYzVReUeoPI+jbsaCbcYq3
qj3F7WCf/Nl4Di2N69eIbRo+vaxDui75iy2qrj2ZzTXp6vgrJLn0IVp0JARF
bp85YIkwY2jcN3o4iHl4rH5CUMahdGv7dZJEkQXx0C5YIfwiregWG6KFwIN5
t8OVey89obBYcWZc+N1WCc87dVyucEzA33DlvBJqghFCAkuIPHaXIDuEssec
5JLJEsmprJ6LS1BdfbpL3QlrrNi7KerpGUVTz4K/H6XC3bO0ezUidAgQVLeS
VyC/KZie5YudXFwGnAc3Vqdk2vTZX0rnnlKnkWu05m09iXMZjEhOzraegdVD
grEyqP51zwXICOg2m80oRPZTAAuTVePw+gs4x+9eOTm+ifHyFUB56elxa9LO
IlSO6ivE1/xVhh0PJCUh6G9F52o239S5I9i8fKHSoOjWv8HjuwPVffNwPG4N
KZcX2nzjdhoujP55a7Jz7H8RSfb4LHTAA3FcolF1bb5yQcju+NaQYecfdaf1
Wrp5vSi7/3wmmwO47dousEYD9dpLR1yM7qGS8xXWWdPnazv7sKLC1TtcK+gc
5M3DwOsVV70KDMHWbaU7O9xBEDdigaiC+r0SLO+WKeGUyJnDw/JTUCzdM4/i
MpCK9IE3ezAbz3lydAS8K7d8FEeOsjOoc7KVvUUde9b0QCbdWv9WqkqUZX9N
Zr6QQu7bo57Ns2kA3OfKd112Y9fRjK6gtZfLNzWK+eKbK1cCQ0USSwm3ACPn
4XWi7pvoo8keTCAwIdXnxRp6F9DEIjwcgseE+hKHtKK0/DUICeSnl4hM4VfS
vFWuAsIMkUtDDr5/1tYq7s1d0KmR+9WvXNPMaUaALLfa8KGtGy8AYyo7Aa3Q
KNatih34cNWM1mONL3h6+E0MjFBrKoEqpFgrCIaTUpCXsqTdbb5dRajva24P
8IGse9ZLAA1p+EELXqhz/FZUUULILLwnym02wqBjXap9dUmJjsQXyaa/76HU
NIzrwD/104MVjF/odPm8+Q+dTDmWL54ZENGDOZSU+k2vQEw/9RFQb6EKcuOr
8kHtkhq2v8TbIPdum+bqQwwNHpnx0wgSNAk161ca20Nc4YFNkF7iy28JgrBW
gkCWsQzsF7o9SDUm7FfV9pSaSrImT6131DwOOPL5bCIUDqPRyZLSbrGpHsiE
meAWnbQAh3lA/KJxc+Og/B/1SNRURfZCN7xeR3LKjTVOI1aTN0srodsm3y66
qyqcRl5FvaSje+qYcbgkzXj1bWJxPYYYmlP9YKHKKxeAWBYTec5dijKrrWJy
76exO7o5l37Q9/Xy9pa00qDMp0hqyMPAnvlmeNtygaVGfczXbkJNVjZTQCY8
+DLXXtTs8NvT3UEL6ew57SlAYO+gjRbG6mm9UrUkB/PLUbn3KClDqpk8n/4h
W/iKlBdgn/MTYOPXHn7rglzDf6logsuuHE0p9sCgtK2gFAF6kyjCdOA3Gr1u
q2A2ls0+IlYuPRFmsQBPO5hSNttmVSDQBwbpH5suIZSehLwF/JxT3caMr9be
u4sT3n9UxWHV+Piv6UDYQAc79LCvIR7yRPc57JbaIfOYIWtr+nR34nmF7QN/
SYw3pDw9XJDjrzyOHeYd2icKlUf/ZkGn6wjME1WG40vYNmm3PhKUuAGkmzon
cDbQu27fQIjyuK6/NFIoxT70q46R7w5x0+6LKpePkJe5B+C2CGqzFr5YqNAV
dANke67g6gxwK+sDYNrMYs4N/QABUYa+0vt6leJFY4qTm1yic8op1VbhnXlw
4tuV+y/ypbKZg4jQTFpVww8TeuE40k4cRLLSiDavMerMM4Kyb7OI6bHeLXrX
HXyAo8hPL5XsHbtHM7o3z3XOzwFnAQccY5F9lMi2Hl4U6z0YHfQz5QKEV8Pr
vRQMtL4eprDG2hVEZkyQZLARwi9O/w/b9ckRB3d8BgWzHorlZ1lg8SBRwm/7
ocEKPElO28Q9+xwk+8pCGoR9wbpbShWlM8DlCV7vJ2qCXjZWq7NoR3l0HEQ9
U3hbifdPEotyinERQWPxceqGZJsAKghnhoZLwtqvbOpNDsIQ0XIi42Bcgr+a
0PEV7C/D4iu/IHfIAYYSvQ/r5rz73i+SrLY9y6WepvNgaDveKSh6JGRmGooe
LdFzPZPV6fcLujuhlS/VRcBpEorfKhVrRmlqsdbVfpKJ9Pj9kIYAoTKqtiLJ
PtgMLKnr8F2tkk90BuDQfrN6UEwJSaPFnX0Wnbbtc7ZlOxtJbOGTl7u3UcGD
U8yuL/RHZ2YzjgcDnYqMnXN7JFae5Iyt1Y4vvuHQrgROJvNZLWLvBqeAUvwP
XdvXRdAejcuUNx/aR5za5vdAzPau14yntnCg74o1BFGZ96OqARoDHYa9GAsW
8oCEiqKD9/nhXhOm8+vGnUNb6X76deJdMjqWj3lvsA6Glmb06LadipoQDStq
s8sL4+uSMS8+I/WIZyvkACmhGFkZ2wcGtfEfuWPTPxRjdzW9O9ph19fu/Vdg
COqoW0SYqSTS2U46ZoXLu0szUpgyiKCOi1dQeHU8pK80TmCBVAbBiFDiMJAP
hP5FXpmGitUDZGlm9qRnZ/PwrnULvfRhNtHte0KdbCgm3YofvHdww6xY4bri
JWlW5Us9utcasoqJM+WKLmmghJlXGr7YmTEnuCHFDZO5/Uqepu8EFBe0kdd+
dBdKz5FJuPvkAiVGfWBKoRRZCYllPKqYfiMabUBMK+XyHKybU5TPutBsLUiT
3kbIbYROJMHUtlilZ612InTbLr/FbvFas8ST6U+0DHDXrl+drkpNGhnsk7YF
DpZEuTJfSp9eCoGmmq0Ris4nXUPdUD8FpWcTORrf29sZw49zTg+8vAgH+m1r
AYM01Y4P9ghDMs2TUskGbWoeMPYrXJCCpnbuIipePMedcH0+jksnZGXzKSF9
kF2f3ePHmFt0vaFdKU0/5VYco40kMfxd5i3lS1BFqmP75Zc2PW0Z8kHjqS7W
KdxKpalJ4CadUGly44Y3ZSk50DbOHiDccG9mEBM7z6zdF93ETBnvf62GAmKQ
3fTDmLNIyDOK8lmdhL2dHZw0xsBmgNcPlPsB8Lt2wSxuQxqrBXwKiX0+Uy6Y
gRuIui79rZpRWqiewRekO1p6epuEFukd4CBQr4n12yU9DQVfsIP4VjNC9WMN
Qlq0bhmhwvmhFuokX2Njvg1wAtpW9EDJ4dLwj5KUBWhjV6SqBe5G5fMvMkvq
zZLo6DYW06TrdK9uRxh0HQpN+KgFDJiLB0I2REvvUIfnT6n+9tXpDUZtE2HC
VAZhlObC0uDEBTeFKh/8XnSnmV4s+LAso8tKVe6qLmoU6BNkY+wiVR+apAB+
EC/wGkH9ojPomhKqVL0e/h4n2OkiWYMwqkHPnnCEmCYIUZ9sHnKVEwp8fZsI
mcYsDWnai0kCICvTDrI7NlY6qDjksi/NXI/MQLKr3uhP52S4A33HgzZISFvA
Bhiu/UxsafHKbsD3Sr/Mstf1DiaN5FSkDE7+DA9vz+g0rdvtcEEZhrE0K85S
M4uQkpwyT5T1ULsAAiSnUITeC2NyPTLPW0RQ1a/W//Rc0HHvVVAouMS9HbGK
GMbquv5/rEGmfFfa2Ozrs2FfQwtsV/5X3oDsHoQIIb4VYmScJ3OTeMXb6qa2
hhVTFj+5lgSnuvT55h/jxz5zsDKz0Jr45pyfX0iL1YSwFl8JepbX/dHUZyrQ
U3KZu3OScMMhF0XRMtWFp/JRQXk8V9WOWSM1odaZfNQxSW5c+O1ewUqUMw7b
yPfulKpww4ZD8YuDfTv5Xj3G7SMDX6yxoqVf8ZtWh5YRI7Q5CPtg+mLQ+kjG
mP1aM2TO4pHLOGj4pqssaWVw/MoMfC5nXF2CuVY05Qxt6vChiPe1u4f+tcY2
0FKCVo37Lq0qdsSEKi/QRVEyhKhSfQHJSsxtQVqpNHBVCFrG/cCRHWMogdOg
PLeOXB8+mwzF3+7aloYClzE4IDha4R+JqvVGAspFJhVKZRcIASYDs5PpEWa8
Tn/AzJrEQRCgHYNon86gHSQ6Uope6Ai+lQXjwv61QAefVO0axLoxAozoinIa
3HROgQVdFpkgmKKs4I2u2ZQmuiHGkQ6T0kbeI8zVNiYr+omiHJ2BzA5TpXbj
gSZNtEMPXHM7sGqHeWBovJVOgHcoGfQvqKO7np1QixOGkAEUh3dEv1pcb4hb
n5kJR4Sz20TKqZsg3r1jEZw5LkvAV20KQksckUwnw5P1VkKIt3mExxdXZP8Y
pr8DZLDCbBJFgpkEnnsmXtsnZazMb5PPhM/qotl4o3Q2ClwGZuisO/9JmuN5
H9a8Rut6R+NOfIMzZMkKWZ3fdwwfbdTfcj1zzWy3R9y+2camzQmYT1twBZcU
fdl5Vs/eDiKVLeleqz43PQlf6PHEdcj21Xq5MbaJDWM0jsywau38+eDgghDG
7k3QnUcniZLqupKPR048PHFrR2/915zSNk5pPGA8/EmfsHNDmVqQTsvpqwBL
M7w8fiy1BfFjAp0uAP3owcizBP4vo+eSmmY+8trz97TDZZyIvP/wwzIYKk8R
ZJ/MUIiZwQb+2qTcBpnXFPO8bykfjc4aVkFXRF8nqkU19BVAFnrHf/nYxX9I
lWp56xOH+FT9A3UK+YAB+ziBShLKZ8Y7aHg2m7PPuhtv404zEHb2B6CukH8n
nEFeeC3EWsx4fNEnqdHcfDDIpl0fJNN0f4tSGkxYgwCHnlHaCLhAZrhKwZTt
BOIeKYYgoA6kJpcQv3SEbx/Ks9LFKQCMqSga6Z0vOnXZSmCIVtXz6FIZJdIb
JC2e5tDhFDO4Jk4lOW9eAL54AHVgMJKpMO0SKW4fdU+EfYKLVpMkCoXDNIDD
552yMVcqmqTLWJh4g4pgJwUIS5N/92PQb40uD6S8hEAaWxw87HIkY3pdXtF7
1yd/JtxBVpANQjVcge3zho0hD8h6TUeaIIU+VGoprny0gC5cfa+4VgedauZJ
c65iF/MEvRBgiymSCuXk4pUjNyLGvicTAd+RP1v7jMs0813sr6ebWeEhT41T
BJXm2hdDNY9WabnjXbIV1k0KZoQsUaUa+k569D54DbkYbAnqiKNMTXB/wCIl
SyuLazwavEdyb+mPyGVd5u1lsRtqv+AcLCMH0nVP3y4sFBKSGC03BMp6ZwTB
V8RI4vxoK8ftbVPFLRzRnUTVM4Z2ca+XULU6mIhu5lO+kKclghUdRuW6oKgb
QB1ymui4V1KacNVBow1U9hJJEewetJkvW7DoDa9bZLuvmpmRpaf1Ni6jbKsa
2f3aGT1a8dy1TSsaem96ZgUrjkiLeMnPadAa3pHKbq0AesRee+IpNMWCECZ+
HviFnQi8YxGo8NTdDLYLUNarqrBdP1WlvptMYkzcLhsIAr7Wg3ocEVzOXi4s
DMXwLjwsfHhn6P1+UJoKZCk6VrMfwihZ905jMbuVO+OnEtoIgMxbjk2o/soK
rEPVfJzsjrl065x5ZsCMjcw6bWN5EtBfMKw83a09FgB++f5H4OY7zaRlb+v+
MBB+zSMKYrI7Y7/hXEnbywoPxZaZL8kb5u7SzMFXRETpcUKDTw7h9D6dvYf8
RlcsD3ZQ8j3qLQ8C56APPGLMunvfELIxCI8fcQDIcDM3KFLMAGXVBuZqoGPP
l4F1WCloVoxqaQj0QvADj2d9kV2DPntSWNp7M9b5TZ1AN1hnzQM3IuQ4EYaH
DtgVDV96mw2pkHe/dmHQSbdU5AxXmbUDHZz266SPRjh+Y4KoYjto1WjWPuML
L9zw2kmxkTCHGlRcLCGvfdAICwjXF4AnCenZbVFMwNSHa24LHj1DBznijlDr
QYWVWLKrit16y3cHkl4HJPsKwtXJPwbpRuBCR3jZ0AZ+gKFT/OeeGtSH2l84
5WAiHXkm6IyrE/fcJDgZoAX1ipkSczCVMbs79NYi+TFSoo4D4fEjI6Pes19C
R62EFbkl6v67YM8nSuzmH+50Gp0JJPaJsMiNWUPrYFjbJJUItxcnqASbVFgb
9A6IDvUb1qW/URRo8zYQxMrEGR+zKAF5kFXkKGUKuQoMq0VQsJE+i2Ec+/aE
Cm4/gsrZE04pOupJIIo6KPiWWi4PFmRvWNj2jDtqy4MUlfIEEE0GYrKKD53F
wEWhp4jhiInySIa009gI2vugk+/QsHZzoPzgjcz4Ar9BkYe6svfTut15ldLM
RMresiYca7HwRSWVu7xBQmM6Xt1OoD+4VTrRXObtcn9GsrLu46n1nlIe90VM
y91QwPMN30wlhG66FtnZ97VjULrWqSLenxraqadPx19W3lYp/bmq4ZTV3iFU
0ahYVgDs3uEK4RuPi7X/conpzajvnW75cwF2bdybNpwZZS0nBOAZt5Zok1+M
ZLexZILN1ueXBoM5/mBrthNNI9WDonYeuYlFnafbdnodma1m4x9p/RKi/PCR
ZvW07gnVhF4GoVG0RkP4PQKX7PBWLXq3gulJIWYxvFCOhaxO+f2KtKTH0fGr
QG3xE4eYDiT66nECNThyIb9WgJzhLPYuyVChLqONekgHWdeioiAwoeOstKW6
4ZEX21qOCbBvfZrBQhE0taLJPNan/J57nXqxIztLN8cs7wVSTwFju3LmGqcm
3TtqVeEim0H/fyWejMlWAwI8XSHw8gicC5iXjsQzM7ddZ540P55DLLe5metj
A19vl7vDALnLm2OoA2oPVfboq7JY6CUhoH7x8rKH7nMFiA82usFGqrJ7U8lW
HwGpnl0flfBNaI8Wt3z1+rSVdcSz/XvPM2vSmcxNSYzy+z4rNH8wRaY370DI
eKqYBJcS/984J/n9bX+feJOBPdL7WZ/G0dlXP4zWzMoB6+jLdd+ZPRJSMr4G
zHfBDJLqUMu2drbltCIUgfmTfB2TKaL+0340+YCKgQRPvJPQ0dI2UinkHFQe
Hoc97HZ31W3NTgPbNvo4tiybtrpNVGlWSkjkXGZcQfB/I9+hnfI91JFXMkJH
DwdCfyiC0ZcNY1t2HyqUoym6SCEWyCrDVYQX6bEmrshP+ZXNwzcLsiba2b2s
sw54uQQOMoGTCg0Z0g7hBYXFz5GXCauGe0aPou0WUyBx3Li6S5JxyptxKafl
uNwtBJTMZEJyQw2nflAy3nK3YQOD4ppHt8VatQv2NN6SRfYflcT2MP7RZ8Qb
zBeZxVRogEjKBmg5Tj5n+nAUcKJVbJxnz0/5P8mKb4jk3QvlqdFOm2mgJz9t
LlSIb30a1mOrwRlF2eeGeQ3xqRYXyZBgtShWwnh8R45ShE/Q9sRCLB65R+Se
Ogoapgw8PYEpRocyZ8eklwAE7PIxIMO43EB/nFknJZOuDdtKjjtxPUa+uUJ6
/iHtpLO9h4eZo1Yp1jLzOLrUd0k172ze0ciLWeTvZoSnePIzepcGne+i1TPF
BqaXWcj7oC5ljnoROWasSR/kWgzeQraPWf30r6S/Kmeeyu38FHffld0E/L8R
BbiRrUXaQkxQXqNCn13Gooxwj7SY5wMBtTFGlXAdLEgOQQJtfnV0WPjvTI80
556E3lyrPn9WaIMBtRKMP9UXQFKoLEOtcZ/CfQDLIAuvk+19VPg+3Fw+cT6N
LSeiFY0nVsL0S4qmKRcCDxooNvnvNfCT5dSdFJ5gYThLPnxNTyeVuM0PMtxS
deEPvJV1+6QxHRQEnXQQXW7nQDYgZDREWQlm5CuJ3fYwkTxdFOAEfDTt44UB
11g58+b4vlDU1Cn1NhKlY5nxDKK+RhNC83RRP8QoFaV+x89V4xmLnG/LP3Qx
tP40+6wuvYIWQ8fK2os5+YUEf3EnRnbVkUslBFe1wWeqVytOi2lgZi6CJrIT
DO9w1/WS2dZ/+858rZZuE0h59eb1tBw6pxIofgclZ1dmm8cY+7mUQ1az8Hw/
Ne5f49uZxM8huPjWKh782qWpf4vDHn94VazGofnV+ULNaKviEctmBM6OGmzB
gW6YbX83ssw7RmNv2/kMqVZk/oJ70KD7L9Hh0B+WdgM+L2QSUrcXGM5/CoM2
fjAxNa5B4S2cXBKzjLA/l37dY3cORvJo9/DbUfyFMmo2nMhgimqz6V4N2fOX
CoJszFsRpGh+tvU9hMwN6nCHe0n7irBbiQD4YNWkBXWZsA5W552wQ6XyK4gN
B9iFJNS9oRKL+qAH+rAad1EbcBFEG13gHvEbXl7P+Tw+kUlkthexgXWkJpEK
Kz+rQRMFKmC4mu4sLouDdUq5Mslv4FoWEGmfkjchK1pqg8zjzZuDs2BcCh7V
TlfzNSt1LV1c/RuHOwuw6QJ9pZ4BClHG3+eGePYkKXEVWtT6e0VAYbOxIaMK
HAYo7ejR3ZS+CJX5atU3L+iYFp2g57Lzskq0MQtogi5HhgWkqe/x/cp1z+H0
CrqUgksDduPmZ05DWSt5HH4iq/kWiomxkogzcDVjYqgfBP7wqUFH08lQcAPD
BOSRk3VjTFI45zMbUWNA0iOyMQ/4t082pKQ6YHd9LcjLDTbFYmknminzb8+k
qmUusYqhV5ab6F1NsBo0EazIY46vsGlZKSKMXJUzCtb6dnDZlBS289T9Oig6
TsM8YFYyuQ5a5CrQ9e6ycpSgxx4HMQyiGIOnsNJnr/nFQ4pLTEK5VIw1dr1K
QRrBcf9y1H5gGDV/CyLRsVAnc/+n0DKqPCmq2TUo5DlB7bfyev03YwcAwynW
CKIrnL9VMfUUNste/UQZreqkz/YldLdelvA8l/lqkiYv62Y8wFdSHBGcp7th
Z6vMMNJn5BwfNuUtXV2QMx4Je/bJuZxYViEUTYnHywNz148u786+290hSrbd
RxDhZleDjG3yvKaLsAsZ2KzDFIr+Oi53F07eiE2Xez1iIvw564ojTmvCL9cv
WcTOXoqvEeL4SxY51uvaPb2GJSEgi2B7+hNGAaJeU4N8OjUPdsHsp6pMwoM2
Fkkr5w9ejiyc4TyMeGXb5M/KtsX+Zd2b0q4Xz0gkL1tTrRuvPmQPUY2D0S4i
fvXc6E+gzjG1zmsrNkewPNKGK1sLPvi7HM/RS/EZMRN32J5gWNqdC9JHQTEE
IhlEsDfdAsyDawYtDwccyUVngQD6gB+Wev4TjwO8kp/kFzTsWrMwjdbez8O7
kwmIGh1Fb/iz87YWrlpaR1E4QNjxIijMB55sjkrMMC5nnURyLg2VzQt+19dZ
XZGxGE+GrHhDhS4Swt8kWSRjMzDMcXHbaFhDL8WpuXnnjCpma5X8OsJ63SjD
SoixlvA3nhuT5rvG1Oz4hZ2cYdDy/7oTViMeHPbJbC3X/7dE9784cn4Yy3vB
MPN8flymBwkPxCm+ZaeNrer0XbhU7SLVk1jtTPxvIc0a8tFgY9bTbKPVNiRY
/ock38XK8d1aq1hFD0BsFMPXk9oF20dQcapbk4iHpQoiRUz/YmP7I82+4EYE
9/6KO3H90iDvO8hsuwx6DwfeMQJr+YMBEvGlyjevfWr0RUHZFeradnU2e0dF
DFAdIVZ+k2SyFedxY82GCBZFO8yPdbKdZegPglsH5kOH/NwGwvSSOjl7kgDX
QDuX5CTVxYBAAtSELyjnTlCl8+ByxdYUWnXiqdvWYi4ZsTx0hSdJY+eRngD8
k13Hwrb05wiMjGUBk7SXFt5KQKNsr9DMdYzHufxoj9XmxGbxWluTkxmX3nT2
Xa2wnZYvZ0sxKc1FcsHROs9g3w0jCMBS8ttY2naoPAWtsy8ZXP5SvMohyUBB
dkW9HK1ASsRcjYBrkhyH6DjhQnMr+DQiEvnkqP98Hv1gXyPpcVtu4ghNG0UA
CmdNz9ULQ1XCvXfYsofxS7gDSzdUxZSQaRP1b7UfOqKq/D/13O9tfLro7xP3
V74qWfoyIBAWD5dwerl9aNF5lN4UNgL5YBDyUZkX8k5pltEl7z4SbOKf2k77
uHTeV+aPLC/IEVlyhDet5DFN8s5t94iH2dfaT1a7jaqh7iI0bXoFIuWXBuSx
6Yir36Xsb85SPoQ3BO/zLMYBDzKLw6pX53DQrC7oELZmssQTS/FfzdOl06AO
lmX2PfMDF/PgQLOQ6XFGAElZy8FZmpv3TovsXpAf50MAeZPd9a9qTTR2kKhx
bz9Tfcm9G8re9qY+FzTebgp4a89HkPwthIoaPkcFBW5qZvzD2cMZ6CGVdhNc
OBh4OIacU7hfzIOGB8KlXg8QcnabB7CM7Blq8hyIA5TA5v5CW1OX6UmcIrxU
Uc8jgtwoFb5nbtoMl+Vx/3svBgjJl0R8mcM7DsXudy6ii5OuBnwhWm9lku+S
YESUHmtGn+wgiSgaPlKHEIZrGDb295NMwEBBPhV7AyWQl9VxFDAA/25EAEkr
t00LzfafRQ2/hJ8YQBEmQ7NDjrP/7y++oXOKGImwLP7Nd9MQ5HwmfTc1Ob2v
qnD5ucSEjTb4kAcY6AnnGNjbl0XmZBgGRKgb/7O6hPvf646X0zMnFjxPcIcw
Gew9wpyAjfh3OO/L10DnIft5D0BRHSms1NOXXLGZ+0JlAcmR/yy9uIyfTBSE
7PZzQazgPop27l0/c+oLvss27rtCxVmrSVsAmydugyOnIaT5SpMZzPuDQFsX
KzgyuOxwX/+RcZlhKAx1zCQZ/LzYLvuLC8krkVxXhJNCuczXCDPNuFvVMuax
EARhpGbK/XxxZtRnU23mxuhNT8cai96DuXIo4nHu2rfSs3J7jgEf8DzTUYXB
U3lelb0HJZtVXyyXoO2JXIQlnUSMwOTpT0Kw3qizv883Ya9Xchrz8CjjfdiU
hHNWLewfzcSA0gcKWS4LMHdqtbFPsRD3nppQf4O8Id0eYGpNgQ8PEXTh1jwZ
4kM5ZcxuzgpZHwyifax3X+CWFLcEy2TulEDeiYSxlGfOwcjdiWpmFFU7zfLZ
SoOtifzmnBwRoqe9J48Y9ihr46XVGUdHrWjBbQUwQ+hZzsbxWA23Va64btAh
wfvO9JxCdyYDtbZUKBINjZv5Z2jx4uvxV3XzTmYNj8JtJ7qd9AfaL8enx87+
aQKh5xRndm30bOcYcqDIyCVEJHH42odOJ6DxEt9asf5WP6bzHUZRc3Z/lcVM
YOvmrz0IysSoOQpajky8WSy6lPvPyE/w7lG5bduB6l+IvdJWWSxgG+aNwWGN
u6vcD0A5L2nfncPQkmVMOtW28GxY4AKtcH/FFMi4ctU335AsLreo2nzhCSNy
4zcI6x9yApH9vWA0yxdSU7GUAxhOrrI1ekNzA+DS2pXJwTflH+HlihTdxEFt
NZUjuA/5MNwamI3EzJEMI42YSK8tpw/B69O/jXZci6tSNZ6AlLWA5sSmCX8L
VTgeljzAEda6TECENcCOhxSh/pVr2fFsn9V7hPuDgF+JfymmR5ueMKWi4o7F
GcTiAbn29V9YSj+xciztzvRrvuKbwuoSJlSgIOV814YYVaPgodsePFS7PahB
wknUSUYxoMCdcUwrclhuwxiBBo+nPrkXG/hjgj826y2Ij9YSrpNruRtYuWL+
QV+069sCZ2wtX+WhOrMHqyTdxHzim4fept8jDHoVnHXdpC+HJrCoVOlNtQ0x
H6xykh29DJ3WJmdoWgr6aDZcGC/CLP/SBugcLKfWvZuZGRUzeNSlAFmCP5JI
d53Xztn4rJbPXiYmIiKw5bqxUsm620SUPcWOhrBVLO1R143J1Q3qw4X4SokT
OgTfBXiuUxnx3JlU/HuI38QEbR+MsoQvJ8o2RFRLzOgAkMNS5J7MqZ/5Zyoa
QQSKmceW1g9lqOcbzbSTZPn+3pO3ZzfddWCeWi2I/TZ9fU9/kNI7j8fArOqJ
Z13uqjNnr/zW6rbu5HcIGKAiFcypWSUxqBl3/PNrtS4cf9G2hB7GHC3T1RyS
Ooy2on23ArPqCCTo1VTip3/ko/f+eBzCEKt+MKjfZHbdD9qUMPHYZ0HJBRxV
RfIlhhdr7Gfn2YQ+d9P///cIMr0ABGypwS1IVruHz2uJmZS6ye4nc7fNgtIw
e2rvYy/unlO9Pkg8t5H3GA3zljeKVUqfg8EjtOPAS5Wm/uLYmntkCj1AZfcz
P55sDS3Sx8apSYbouJmgzlXCyvSnLrERgnsYofT6mD1y/WXjxgOl+oiCfSf3
6XEyzhWjbRDP2/Xtna1HgCUEMzMqCIbAzIHql+V/IougT2D8CJnVZmfjaKkY
4F4hX1z52TF7AQyLYQwIftBw/gUv4qus6OMk8X08EZL/C2fDDdb8WPfFlZBX
YT6gVhlWSI9STuUnqFCzIfLV8vo++lBFk0xE2/khYGhmztjJ4bX0+EdH9Omb
S9bOS7fE4kOC3RPmYMlgUyXTr6WjsYKsxCHpJrTIQ+raM5KrlT4MySRbdHto
5wS2tB9xgaqPJxDOYNEJKlF6W9nPyEUR7GdLnnBSlRp9jYGGt/9OHtDK1XWs
TBkeNNZwCGGyBB7iwlpIwsx2jogocdlmSRxTkLpb6IL4VI+HQa5jgvAoJGrI
V9RZabLb06pb2CWU6QMRiPkRFEpYcFW2C3XHXkcNU31HVHlRFKRyUF2qPumA
TCZXipcTYVlAuQLlgT/Hx+QpSTQj+4nQA07BUfL8JIiEPSOvNm7PIOlQGman
4g4BipC42LuWvFR5j1WfsP7BcjkoOfLruVdhyjP6pgvfp49fHP6shynVQW+A
rrmEKFHO3DhsfuZgfmUdXmo7EBrOhJr6k2B9cBefOwPJlY+IPtSloVPlnuTA
O21QTIYvDvgjEGwvd1v6Aka9exwOeqPWAyZNHxs7UoCYxrnis1lITixQSwNu
HO1ko95P5UgGdOo6N2qQXUXVdsDEj6hQVVqoHWwdFZflMvbQOsIDQtdbYWUQ
U6s7X6aeaPJ81+Ii5gFSkNs4MMXhmWYvBQpeVyRR5EO021hfZtieYUqSPNWp
S72gwFtiGBvDClz4eieiLHD+lL//tnctsGM4GD9u5O7TYSH3Ll3Y3Zw1rPi6
EHvYzXSQYtSDc7kM//vhPYTG/CIPl1jDIu4XRWoDKNJ0cwMc1XXVEAsFwOof
IHkoGjpYFAMlALO0UfxOEaB1guZnKxSCn08bS4FR4Y+Q+G9JjNiKMGt5iXiM
y0rNKUDF77Qi0DdJ5iU2VsUBlawQWvBy4IogBEPM1qdOVgK5K18XZjQrno/f
Tx59icyIyRsn0b9vljyShQe9eQZIx4iud0woH/rkqAoi9mNA6k2bQh0wIEty
8hlDYsdmSJdh4zuAZMC5n0QrP/1PTVWI27GLsPQ5mcby+g6O7thSPTk3o3gT
0mljTRSuiWmAQE3TP6uc5OCx9s7nh/Am/XZ/kNGVl+SQFLopJM4aqkKkiFXy
TF65hLxm0ennjeTYYpFGv9sRzlN5F3cPOsxswvaUDxa/yzAhmNX0jwQXaqyv
R+S4h14YysOibnRjnZzvgpHf9OeQozQK54bHFdFpB2zE8nHdkC+DkIIBVlBo
TjU20ddUjtlCKiIArVicWJIG4JlsDoaRH9i1cnIsMAWm4eudNAAuxcWDsLls
SqD3UOGaLipq8JbT2e92BXRiBBZB5hRh6QMr1xsLtzjOByr2mz48dC9rTLAV
S+1qQ4xAG+oUPy43EYTQgpNtswRG+HgUJcilAaXe8fdpBystUCloVUHIKnE3
qXu52/6ZbASKuTKwohn2SCY7cTvTcuq4YrHlmdHERkGZ7PtUSk7kv2V681PJ
vgdhy3YPvilbJFBB3bkFPcs2iGFnf41pV8k/zKQC8E0w4SIjHLDrHo24dmuj
hV4DoPo1oUeE2FaDwMX/6sgWXbCBLH2XmoWjZc/5J5WJz3OEG7If+Pft9Kdq
2FlR4T1Y00Vebd5ITWdQz3M/XMPkb95P+l6jQVH0K1POibMvaj/lFwIJBvVs
oW/RCy5zZhwpzA7/sGu+kKfE8kuS5ecQNW5P1bzzRcvT0/JbI9DEJe8ZZ1+Q
jbLuxw5WxuiClAF8w3OFtWUSu1S2dNTpuqDt407fDSXoy5SaIB0sg/AlGx6n
uBRGN8XxmTo+pfp/eVxPMgJPKXuYCLmVpLfEovn5PCwq1FPxdJqO5ElT9Kif
iknCs7SI6QtDc0qAZMR+cgfAd1+LvCJQj8hPvdA4eLvZtA0gC0g3TKv+G19+
T2Hb+FXm5lNw99kxZ5DXonjs5WAQPlZAaM/sc5ooYJgU2IiiWaJ0lvgasJw0
flumChKyTLFbCj70fFxrbu4gOiENUtBnEiRjefRVLDeDxPr6xhyM+0XFmO9C
oDV+VIjjQTzSCGobsZvPsRuuKEcrfuwKAsh0UwKbf1WFB541Km30OIeTEWur
/m7dE6ykmogN1hEbOBn27rOaN4YbqLio9rb6+Wz1eBHm4zWTNzANvNhsh0df
mNX9csc8pCASg4EDsVpBoqCzpxDTc8RG6SVSGtbWX9Km5i2g2GlNhpTvVmMP
QLT0XptPE+Lwm61tgeyJIZgk3YV1sMLIuSzdwZKjBaDkp27+liA+a+3TPfqc
Ud/xa/uqFxna/y4Fc4DLlzuYHu1HU6TnJdQo+5zm6gf9nu2oBW08FgjcphGY
mZmtqeSy2Knp6tfiiwlrxnK9+l97A+SvQvVOb+WKfOoOSvoee4KyL5dQO2CL
8TGEfpCyU9vw4fkF2A2AMEIwoTAgnVW9j9bDQedexdNtMCX78WmZVACXPsRL
lI0abfZsm3fnbJepNUNGWrScZFlJW93cHlh8O+jyxE9eGIWqEIRffvZW5wxY
EILx2FrYCVOHmAUW7fJCTlb79GtmOjqHT5UOU++y9WEHSfkVUwCeLdWWQibw
oxYEdQ4CHZHyJhjb0XEE1z/SRI6eoBNMstv8UT1M4p1OdcV8Yjo6mSE1O0P9
DgeSczpZ/8S4pKPVsdDB8Ts3kc9rSDZExzT1mEJ6OddJ92jvKzS000GrqxL1
kLhrn3pIoweME6PvD+WnW3uiA4cx9l4vIZZvF3mRpPwvogPuI1K4cmTIOJ+K
DrSGvjliFgUlVJMp5hFQMtw3W63pHn6XM6ks1FQETBF9Hqr4fw1fOmcQ33xh
AYglMkPv5LFcwne0gWH0PgCl5G7o9gqyoWIMPE3QqYd6t6w8sNjZTK6IZiSk
unuMsa9c0AkTNAYPMtJYWVZiPrmYV0BRnksdnR95lZ8loFWi/ykTsWdoCDx0
MrK9P8JGfg0KEL90fklSzEyl+JMnbWDHjh6E+qTKgcODdmFH3eoNXtsU7EDJ
L3Q/fe0XKyZKKCS+mnVlMtA0yjxGGcar5zL+4RNxMIQowmWmgnxcsqOlv9Fy
ZbZLInPmIeaNI0PThCxCJV5mD6CHyTOtuiqXCbc/cCZGGVX34UDCuo6gq/ua
P+l9i9yDIofBTyoNskYS0Mk8HSpd6vU/fanw7qvhT738hid2fmjR720e3B9w
jJUoKKrL/xj6X2JT1FwNeDfKk8qDyi45FN+ceHJ2WW7OkjPMBRSSPn2p15Gl
kTYbkCVtYbMhr4gXyGibfE3oXT4pY5IE2HX8HHI7VQsvsEdBjywz1uouQ3IW
+jSQyVsTdawCjJAjckXpN2KghaQ5FmboG/kmIAnAl2OJFZCxbgZSXkMnteNz
aXJiovUxLw4pC6zM2zSUbo3wiEXnc17Ll8SlX4Sc288tzGUpQd4aSGjaKtgG
lIhrwtD9nce5gcbC29718M/W7dYU4qbA9hTXq5ecB7PauJjVayLGleyTkn+8
GXt+Os2elFF5sqPI6tZVfYH52lYOZ69yat1g4P3pvG+KEG7B0vJqgOCqLTeE
AMxd0OkQp7J43AGKJKdXvWAJnJGfNGyxYDXyQ3BGt4NslpUzgKGoSLpR+bgG
IfbmFDfdnjU5rozq7DhswqzLTSCgBukUjP6ljOU5hrykbwphJBsbPnWTyOh4
VrWHUsfQWYs9D5Z4Tspnamqe9SflNyJLtkojgv2FxJuj2F7BkVhU6xXVpYRv
LdVefBFwDB/CWyBSDtjYtHRX7SyBfr9k/XXuoWyUJ7i/y4y0kaNvDVmgRhVL
RPK+l7NagiVbXulI5DAXE26KCM4UeE42rxXuGwDCvmcFnyRjXtnX+QaAgvfS
KdnkeBEJedJe/hN/UcCxTYKWYWsqBWzBIRPtVF3yJXArqO6OBJvLZXKDaCpR
V0iB2ehKqMO3mWUzLIUTYh2yL3Oo4R71nnzkShHzV5dFBXztOVpBbobLmER5
eL99LKSxQvaHDN0SRWthMRIp8fRKzPGmusVNzS9z20L9MKMrcNhFNlcF5F7b
MTR/cdyMbaw0K5eN8jH+6Y+HKIT8ViDsnI4QwDpETUBlya/8bnWrwpdlQBtH
zmRRbydWYTUZzglHoFk8nF+zfe0FEEnsgbURWvlavcUJk6A2vWDzy1zPBf9K
jM+2f/fPgyc6H5lRB6F48qKPE9+HlnjJisRg2T4JV2o6VpxsxD4W+Hp3Uhao
8fq1sF3P3JYgvQh5Vk8gUwggzyJtHdNzwDp34XZsCXkZkUrjAu7Qa3PeWidb
6Qxjau1SdeMN7NwfrZ2gSrgye1DxPh/nhvauoIxDTafge8fo8x/Xbt9gUM5D
sFFsd0T7A8Bsc6JarAymGF0nK+eKOMTkDpq8fDvCAjdPN7ZC1GcJAvNuTIEL
/PoazdqWmQLMoLiiazVKz6YtLyUBk7IMao0kZhaS/tjjitfV/+pKZlR9nZfO
waPGeYKEuj3/9ruKBYcUJDG3vPSvNv1dl0OWuSglOdULhdWTtxQSOm9hmRHO
nhTWL2y65UeD9JqjjQwvk80D2DtzxJWzjpQNB8yXrnPWr1rrx0Qxa6ieU8DY
QkW/rZGLFNv4viBUcYIDvRkIpE4YGCGFtcP777UupLtDiAOI+Wdf7u/ST+eL
mDvWvkjON7klxD62FfjyV12zI59wmx4KZ+qmv9tMwv8CDAV/PHWKSnzy7kQu
f2pjX5NPgfE6tfa74wE5LuaLggX0f7HnCWJy1Bvglg9B/RgD74xA6BvEJ4uc
JQepL5aBKkx12nKPyISYy7F4X87omdBModeDdFJ6neVuWulvM2g30Lx8slD9
mfQBSDxKrvOLSwlmVpjMG4QHDB9xC9WMB93hudpGWomB3J1P8mIppiBJcr/h
xKTmqfoAVwRlNj37jwlxiX1bUuMQnNsu7WfUYlGI7HOpyMvkdf4X8ubMnuiZ
0q+OxaqURQPkmKhqaUjSVBD/X2IMcoIcs085E7XjnCK2oTKSxipnbugdkoCj
rRD8Id9pI6zIHoG3wrwlgFlg9jT8wG9jhIQ0uDf/kEjQgvT/SrxDgr1q7xum
QRXOfZt6GUHvURcs/UwluY6RAn5VsCAGnOdxAgCunAQPxktFI4h7w+CjBS+w
qd1+AjHvJFDazfO87SqV2bK0mWc0tsJQz1kILXFdllVt5xNSfrkVMg0I3f+K
5oKbtCyMSRT+haAOimeRL0afY2xEGysAG23dTrmwek7IvfjqL5eKDYedYMHA
xM/uldEC189g2BJpyZSAhiv1tl9d64K1yXtof4EoL/vb2tAXiLJBOQSkoTn8
cW5CC3V8W91r5SS/okMY0O+uYj4DFTdZjSt8raypBjX6hNEfTjk2mK1O9c6z
c7crQZb6pM4mu6UDbQr0lh6aHBAThzbe/lSjSnb/66DF1m4ZbksiFboe/Hcy
pHK/QuLxdsqmsh67U+wP0GtCDKRoYR/DJtx4WiUtCMuuQ4J86UULJ7lr1TYk
qLv+8RjhVwEYMfbE2nKCoxV6tkwwC0FFL8YvQK3eRx73aXEO/uHPKOn1h8Op
4F3/fDdfY/Mi5h126NFMVsuVkMZIapmHm4NDq5G9H+13aUyON2+1KEw4i/BH
biqyLFURatR0IVTLynR7C/+p4XaAPGAxPqyNQY2z7pevFfwHGkT7lXjsHT/H
dIq4/DAoEXV4hbkZwYcneNKP2VZwJedif7g2OJBNiR9T05w4GNu6dtK70RVx
65Qc4ObconJOysT9NXpnkgd9wLvAb/Zj7XwB1YRnX++x3o4ygTzqxHgTCJkH
/MHBMAxhwO7+oy0Vgt+y9AG4u3XB+iTXPnCpK7/sxuWbde51fQJb9TjUVNti
TjWmAu1s8FGWKSitrta+a7UC5PXpOZNYP7xDHpvAGsiJV/cX73aqK4UooPuu
FWludxHDyXzuL7aNMlnrhES/NR7p6EWI9VPhQEhpdclwikOpIuUrbAwGg1Hq
Q7CMjyPg1vZnq5oCRFvDAzahB6DV2dnjblmHCeAAmgHDsJHBzH2c+NqRw5Fo
UrVRvREPBYZjEYgBKsPcry9QMH0TgOHJzwr7UsnDjYs/+hBHQcOMQFFBOvsr
CHk5tdt9XvSriEZkA9AkUtW85mmmLJEZ/y08y6knqzr008PHquErDlGXCYkw
2oJ/K/Dnum2OaiFkndO8BBydlnuSa4P8LsylZO6ABuMAjVFUTO04M0doqz9Y
Oa6zi+Rpe1iiFwG0bZgBe10YUekj+OcDX/6xy2A9GzrdL8d/brKW4Iwc9CBI
eJaFMas9o3tDKIG3ZPqvmV2BZI2Tt6cKj9CoKP5nAWcVwI14X5gQjAge4M8K
joqpiYq1d1yIexl6C9ycaRDpYcuv63QnkWOrb4ELlkSadKjZoaPwzu/a48u0
j6yqhb6VAXp4ikBUN3TvDOaQ9St9Ct0ud04D3qNssPrLuRXWmQdK0MWXPLny
LeHY+lV+785Mh9XFR85NAstRvz1fshNorcIxKRPfpEztC5C93TeUYKlvpBUg
FgKx2WOsBwOqFDn/N3iJ9/E8TLrTA00CunIuPLh9bywqM7NRoA4I6MvzQL2u
YcsRI9Ydo+kC1Xoe66VA96OGg8Zd9h0UFZ5HS/u3Add5t823OXe4by7GkaLQ
uk8oHyDOQgNNnhvOu/tkd8QHp+Tg7rggUUUATncql+2kdfcTIIpSz4ixv+a8
WJaH7aI/ISIY9aLpF+sIFiVK2WDGCaGoAfPw3pOFZpWLr5bTMUU9rLm9K91V
/5Td3CpEr7c0nWYYpX5A99O75p8fQ/VllcL5hhsunouGZNJo2DNpMOCWMLrp
j7GLlXq3lLEpUco8rlh00BQ3coMc+9abGYjoUwRqqjEt1wL7IpkyChCJBSb6
RMH+RJRBbrKEJkn0sV15rRGiHI9KKiWqklxpikuVDNbXeINHhEjLt1hu6HNx
H6B2CY0pbb3m2TabCs+LGmt18aOH2JotWNftqc7S+ePoIunQOJwM0OOlvnEq
72z53Y0oUeZOqvPDGLbViemWGm1huWaCelsbhGMgttwPqHJFa3wCawCsOXtn
1YotmJ3phKAjqAeEmQwKDxbekfIJSfmoYuD/jMWTKPpdop00Lc5qpV7250j+
VrusHcZuYAIsNobh02Uq6cQ4vcFz8pJPW/XQaZyctD5k+pE7LhynLakWtZYL
QuAIrMegFQR3IwCyV1BGELmPd3cGRWd4GA8rJIUh9PeFPOTPH1FMAW4hDyEB
nrImzzM+Mrdr5DZMDvNG66SYzyDeVkeUXClgZrCAXdRNJg79WD+1qrJ4jbsG
u4C7kFeLXv/kCNBrSAG+xjvXjXFYxvZItXg2EjPl21ffpqw9yb/tPtu5DjtG
OPyhUrGcUqjrpJwuzCWHBA84yc+EOva7eVma5JqOgIMm7qWeS18Tus13leo3
z6aAUAdrQaVGaqg7rjo8HOmFLflQXasD2B7TWlR4+F/pTIWYU4briDHr34WR
CrlluoN1xEhFNyLaqXKmds3OKL1uftIwKZinvMZIKBMzZBIq+nTln8yY960H
5wcwSJ8LMF5yDT0Of70Wg5UQmiyHXSJ8yTDZeewvOH3J0qKk13AFFoGZiP+b
OujU+ZepbyVoTeOO1uIrwpjxX5q+Qh5/iq4a98rlfpf6ywjTduu1a7tFU/OZ
EVXyCi/IWqvRfvn//KMDx8HiGWIrnp1D5LUACvwa1m6i6Uvvcfj5blI/2hWp
0BOjgHXai3a6s8P3eTCA2E0Sl7SjQaDvIv9Q95ZLw36k8uNs5Wn2x9OUR0LH
yVDQeoLMr1MfVPghDICk5stgj074ZYFYIIDMbgBU0sIvA2dH2edLD6YhwLUK
qxhJBXauR+h2cSYvj2+2WinHIwTsLVFPu6EfZPxs8j23Zr2DuJ2Xm1e8okno
QAocbfF7e96Do4lNknol5ymRyPCPaVVZMN5phQuARPWC89zZVaMqE9z+DJoo
Wc//kWyDiB9ifTJ+trBrVbZqBBwzIqy8K2ppVCmvXCkw74jtZ+syKTnD8zM3
Ne8WLw5GGPBoYOtAO7PqYCRAlDXgrdva5zLJ8KQMWssjvuid4QOL9xh/IiD9
zUmP7J7qfJG9rUZ6FlmFv9JCYjKf99m6gOI0uK+1zspzidxdaziDaXEvAPW4
igxJqC6CAPLiy8VklT5n1r85uiwJ4XroPUMl3NKX1XQq0mMgYg/e4sessbYS
yt+5neuT+mqmWAvHyQvOF+tq4WRDeUojCZaa2CWpMz/QG0jLUPiPprbv42W1
nLsZneDzk0o+17Pw5myvNV5eXn/yfsVH/iB7joxxH/TZW2WO93osqt3Mw5+2
N9dmqLaCAoz19llh29HVE5DgucebzLpZqAiiRSVBFnh9Gia2BCc9WfLHQ2cD
Oe633W11wK4NgsCvSv1voNNxxK0dSnXp4LsQ+sbegQrNZMsF3n4RBDRMQGun
WPYx9jAOUiCbxTAmphqV6eUeiFB+hUP4xLqeRUlZiT6+lt38tU9pDa16ehKq
qwfal9mAL3JoAoJX3aUZlFPsDOfsfvlJmnnjhAiJ9sd+QgESOhyDNExuCHzo
DpdEyQktYjK2YIP0ZQ1jigKn+ZP30KTgKPfjcupKUXEiinmwxbnlO5HCQKeI
AlrF9kLH23TtBed48OmAbj1nvXZzro+GCzCGVv1RvZbwRNenJQHi4tYMJRDz
bBYfDgz/SGwVbsP2ERWcplgE7Wq/sgV+eXgN8UQiyf+IXvYBJPa5b440qeuH
GsXHAjJhQTojSpKT5Jtv5UZSjySL8jMR9KU9iO82zIkQzYi+agkYo+8pr4jH
NEBcMOkqGSU9GloE4JFLH3VOBpQZeF5BvRDHOoXJEVFdYHzmdMZpQbKLLH0S
qkpROAiL79MTrgqZWSNAuMQ269St6PsAAwpm7CMOynk/SDHA7rPM1AVXKCE2
p/YQnbk5RKL6jD3Q4x0Kr+F54GqMmB91RV+84CAKz+gOb1LE7dkh1d7XVBMS
E2jr4HqSDZpKXg4QcadVSnODjLmVuAxzAtRWbg5GhrON8R8MAB27+x0gxi1T
eaPMdUGvBeWXpjuRekuuuK3l2R05Yd8e8giMEwIWv3/DCf+4reeSaGAsoGw0
MacH8DAl7xcsl4++4QRdXUFkF/fcfltMl2bFUw3HORftdTrBGOV+BrKsoH9A
/ys9tX6o7zcGu6SCUhqiTAsA+TpyGYu4gx7/LHQuQWTgeuehm5Av4zn5kxnK
hqMTjh5+foQxoqwTI9mhSvTPw5Ijgmz2vG4pzCFoCujGbDyRqO2bEN+7l2qc
0n/ueTH1/upOr2xUtZc7YT/xDo069qQswsR5DDiKhA79U4UVegpgAGvoMtjz
7l14BYvVrUcmfSV9OcNRMYlonVOscDKJS/0cjupdFwnElGs6AZDlsLiXpUCr
+Oofu5kHn3vu67/Dx6KmtxZDlI/YSw9ALdKRtd6d24vc4jStHRNekaKjFz8G
wn/0gVUes5G9ZuADxikPMKCVZlfJom4MzbJe5bBvtEq9M4CeKbxoKVLWhOLT
+Vu9OqoBNabQh6wKVcxkDqnSZW3Wrr0DZT7+uKmm2QLnPNGoBB7P2nCtZPce
VmEm8A64yL2Ei3o5V61QPDet/hbKIOiBlLjxNac9q3eTdui8AWKkblg6wXXO
E+QBLIOdAmoZ0ShG8Tunf6KFqJ3Sg0rNo4rYxQZy9VPM9yX0yo689SgSmgK5
CJoRD3p508ZDUCsZyR7va7pl6aTpqv/gVhq9q9tAYRLSg+e0aftbh+InHGaT
adBV4t6+1Q2s5Xz66AVfDWxH951pkEkmXSghacOQG5al9fCsLAddcTvd674j
MAWF7IzMxw8ykOS/NJegT5oAcr8quLwzb3hmp3D0RJVSLecrnzP7snknMZQ5
Z/NaTnAF1/0ETvw/1G5r7oGKDzt1R7rPAkISP5nXQBSbn1Sum4JOST8q/c5Q
vebwB1Gp2dh2oUdKKQKwE4ScYuEKqRT2O9WWctLjw9aWAjw+r7JI7TdNNvfd
RXxhXGIb1oV45gCJYbETTZdgrP84hIcRmi9cU/IN3vMdwffMycDWTCiLGDEO
VE0TsdUoWdes7k6AH0dh98GQQ9TAui7+NFDQQGe6qjoxBUMDns+JkU3MSPAJ
TKh2FS+Jdg5oPkL7hasuepmREXO3hATc49NYs+CN4QG2BSTfoWHaH67t6PgM
uVKTVK464p7eV1uLqpJ1S31NyPJk/4/DUu+tBLBw4NMaeMHkx8Pwzj9OUDE2
/ncix4b1Rug5RIZXVmQ1XZ5cjXNWhfU11zOVE45oSXKh/NjVWyrVV2APMjP8
4cL9LlU0lnSUoriWOQLaBheAE9oggaEIwUcp5+tuYQYk4AxTbqfjjOksaIk/
dVU0AJuzPuySg9qFC3clUOR5Obn9RVvQDMLgKWWRn+rE7DvQ/0WJ8ZM5zXi5
W0bEYKXQI254tddQFJaZ2SVynmId6Jjbhn/VQy9wnhMfq/jZS6kNBiR5VHm0
SL+XPbVmRVVtM08sNns0KXOYR+H4O+qRkiQXeNNyacRaMKu6VyS/vBA/ILJZ
20sVaVfRpjv2ZTzIey7Amu1xrdWVMQnlCtCfGKlOt59dXz1rfieBoZ2bAyBn
oFAFjgslKz4Mi1YXob0ZivHsb7VE3ZleZWCT9ztehDSsDss2FIs8boORX+Q9
0vYZmJEXK4H2p75kQslWljJHV4stBifF2egvbFaxZHBfPcOK5lPBQKhz01UF
POWcyEOtqwfli0cLTiibyd3bqkuIlIyyt6I9g6CH8UylzrVSzA+ODIGW77Fn
nNIQhyi5GCTvAJTBzQv4aUIEx7DxvhVUav4hM5wJMPwziRCSNgUf1K0vQQpA
bE7hMv8A+DOs8Fl8R9oeF8oA8cosO4O1Fka9fVB8mIu0S0IJ24xMLXxQ0buc
aufAJikB10czPfq9tPVPR7EAKsboKBGWYxeEHPKK1gAhS1T3X5626UWmbHvb
6y1NkE+nsHnjhE/nVj8tsOeEwfHMfmBu8Gmu9nPqeQhs8Xp3SRdlsDOwOP6K
jxwmd4J64EDj1Avni8GK8VNgg4MaI3LWVlM5EHt3exIlUfgmKDo0Y/itkbdb
MYHyzhQVPdxqPslMvHJTbmBXWgiSHbW0QVZBCFg/DIylX0VJ/NK8McpMARsL
r8K1w243eheBz0vGX3ORIRgMfodmO9bAR/DeQBtp+SZ5mTAk7zuYHGVlotUu
G8hMHc/1+YpjU3bTlCwO0/GrcUJNWs8pDPpFsg24aVb1QB5c8UJVYiMyBhLQ
09onVUTKrIKTkQ048CT71O/ifvXKDVbBADJkZ67RP9el2Al7met9FCdo7ZHb
wM0L/9R8LP+9FEs4UGX+7hAkudw9iBRCLAn1QL5f7fW0yfTeqKr9mrJMTD2y
Ed4NxfQ+onhGMzBR4kfTJKZlu0NxGmYRD9VcSk0d7B6QJ5HwgJbUtM8EJrCv
wLlqIxXaBUToiXQlgeWTKV/zJSFsBCRHkQZ+unvy7LXKHjdYL4aa4lMwcv38
CgAJigCFEfrDXQW2jkDKpjTTkJPOYilWU/Hz5obwxPa1R5yZg7FbrSwG86Nq
NDllibr6/K9v3CpWVT0Oa3av2niAIeQL6fbkE216LzUbp/mnzGqGaPq6+xNu
BObNeiQn03YLTA3qxE1xFm6+Ls2wFncJnfD12Dsa08wK+leRfBy20fXfCvAF
eHVoA2vnPfXLFgaWSfM2tmNN4YapVHerQLGT+jZx3D8uLTb8UDar1YKx/SGg
od4Y6OQaQW/lUO+q67LBNZU3uLPYwk+Bxrmajm1EvMBBB6HWppRPNG56RWUn
xC2nzjvFIgH5wUqT/vYU/6A3CDU3dGwru+yWMhi35NkzRtoO+rAXjWudZeRr
J9NayxfBEWen9broZEVeuULRjGMP5hSdB/NjJaMALpskXIeHSUyFanpj1+/w
tzgBcQhUCb4blSqSfJ06Ohy48sEJs/eE3Uche9P/hsQjGq9Od69Ppv4bI06i
XdwDH6S2NS9MyNrB3vtkUFYHJt64zOmWsU6MkJMhmIsdZrHqB61vCNPbl0T3
O3fNRs5tO4UDOvLibLj6qgRpdu2oAyHfdOnIPEGogdgUKRz4G7sLWVEkUo4L
YfIM9gz2P479Luu/EE7JYZdmVsy/Ca48Aw3IRZBkoUebswvxug6Yg5cQ1CPG
1Tb2VVX6wTwQqKagNtrIf6NBHNkgO6zlYKIrR2xPoRpgiHgdmXh9WZhM1pek
+sx+f+3Flk/o+fAKoJCRTu8QF+cXYCuRE0cfXVt9YYSE2000y72tWkbJpqDm
obYT60CzVxPuTXeOvsGGEPAr1//gZ1XWhjTVZGKwdpWkfAbQkyfb4KeYIHvs
pCgUU7C+S9cVVlwDr1RDZsEiLW/WCkI0yCm+Tz1zu3WV69UIppGC4N+aqshU
1bUe6Lw8Q9FhX85NVAfs7Iuh43nyE2MqlvGiGAMmJGhMuEF6ouxjcFLbXG80
9Bnj4uGzL2SKyrPj+jSmlAiduNpt1/kLNoqeSBTie5YF8UDe2i1+3QMTpVUm
0QXAsLywk6CNBv6KcZ33IfQ+n4ZQAvgVZsxh1mG/ZSU3HnMlobnX6rMYZsjY
maS0mUewrD4bzsURhZRFE2wDkLcvA8h6pTa8q3yZQWv48UkBLBqm3ICc9I4B
7/2IhZzaXp1H1I3Wsbbzeuc+nFIhVDDNUxScLesBczR5A6phE05pCGLy8Ocu
lQRidpUQ36kq6rjhiNCXalgvUFMDWUn94y3Hxo0c6JMf8NDcEKqHaq/Vs6MR
khOb9q/W7q0iZwKoDtMeLbu4cv8UchG3VLEbdVkndu8sJ5z/9GfolJk8+unQ
hNfDInba5RC9q2URjgXvqosMTZ1SFearmUFBNPqQArU6902dPh8mXBnXBrUh
6NrMX/bCqGTJf+4ZJkYDUJ1sCe5/6DSSWS5JGk4q2F/8/5Bs9DnF/P10HNdf
wQBquor9lWKP4Cn34GZuxQ+0gCzANZEiL3AjZp3f01GX0rxKpC+9iaV2Hd+L
lBzAdtpuBEMSSIFoAam74DL0WQks9QFb/4+T6jQ5N3GV56ctdRRTp/LDEzxg
c9LYR8uEzJR0GSbbxtoomdgqhLtjgky/DLh421hz7zHK06jH1TJL67EZ+oH1
cBNUPfLdXaizld82Dlmylc+KE4+F0KhjkcqaD8bK6B9in/Y9NpY9bC8QWCAl
vAuh9o47jMl8+WGQY22YGrJx53OZeekDlCRE2oru35BnyjQI+zPwVGcu2ahz
HM3HYPVSv/aniKrU18kOPfXDeFJKdATOr/m5/dohpP1/4vfVZNqmFaahtAkP
/IK5cbgRbOX+Ai/DBTcjHgZjdMXI74Nh5fkwjTJN4fGBeUaUi2wIiSWY/qI5
LWKur0EOjO+SIf5s+V9zA1VlkE6mHGnTnSXk1RhslL+3pmkJ1ORZeA83edM9
kkmX52IK4g1Q1BjgZIsQOo+x+jZ/JKDL2JqNR/+7PQTjU14SPYyEth6Bdjbo
ub5S/jO5nyAyfRnusFW4k0vMb6ihLiwrQg8yTYofp2RNuwsksWGzaU5n4Tk7
dOA2XDSLKA+KhAiiXYZynT0bNQXjQ6ptFjxicGXuCmS1yS8zoVcctcPFiwdF
z9sr/+GFt9qYjXIct+60cm31x5comDTDNztiU3UbVImeIMWS4T6/RkD5zQMQ
c0jKrdEwbNUPhcSu2UXp+jn/qcGITgcwfvYSahvMXATAMWBtSwAjC99N84JV
2Uu5GBZ8OfLqgegtA0o6qQBgxo4Wo3u7vz/HkVlY0q8ThpL7BMthGo7Hb5xX
jQb0C9Eieur4zmvQneKgw7Sdrr/+vj3DlltiBeFnB13WMiYR6hVqKI0kunLQ
9GrecZHRGe7w+rzog0O4ZiKsnM7SU2WrU+iGy7uGrMrgYgAPTq2NcmHX+POt
Wu30onHmK8c7yVpjZxQNR+fphs1wUg1KWO0Eqh8NnazZgSGAnQehNthLteQK
fjH9oIexx2XTLZGWe47H+HT4Q+AiiIIzm9ocxFVYOPnGxgqCRCQJx4lzaSln
n4DNL/Q9ukKVfZOUxOF4Z6H3lcEHjuN+busOhabObyh2c1dwl0EsA0dvu818
y6i0mloXqkYqLxGHAmJgWa7dw/XUNIVtEmHmEzXaT2cH9xdcygk0z97S54ut
idyW9mu21jqU/wkEfqHbiGB6spZKMk5EdCY3Bl+8PEqRReVsYZN8V5pGThE4
nY4TrCemXH2r7avrd8EwwDVkpcioQkdlpUKmJmqFhu3vNmr4MaS0a/OvN9qr
ckyt4mjAtpUrhcOhhfssYorDndhDhmFd1BZu6XNG8ATNPDzFwidme68skTdT
aEE/+xFEAg19GxTLSmZ1FQSPDnNixAITrFcXMD3PtWBOLP6ASge1kvS4yMKP
avJYKzwHfiZf6zm9wmJF1os/NfOSpmBrsaR8I5dGsUqS054I+HNEMS2hQ56z
898xh5NVPkk226s/h8B5WDojecT3xDm6WL3g09I9ejoqw9rg+nvDTat/mKlf
D/FBWy5ifnZbevKF3SURZ7XKd20Upvqdc+sOQIK8zi82/t3SUbbKSjL6RjRJ
uDlVYKOc+ncH26wKEbmV4kkQMKZm4X7S/YQMTToPF4BGGa4rOj0NwzA/WT8j
8q0EK1Dkuw5m4p7m8nlAojn0aYXBxSgfysi5YZmC6Xe2CsqXN5i2Jgsia580
ISEcC1q9pBNzGfjFr0DpbppyiwPr5q6pqnayZnBUAu9yVnmBxZZIDox+H7As
e1Hpd425xY0CuAVF5dBaI1T0PNlIPHzklEvYAymgDO3nGCF7QItYa3/GofAe
db2b4VlAE9135UEZBOUekOCJAzTIwULFo/C/1gq60c4SIMDwq1M1W4UjrERP
ieQ7gMyZbHHEdw3VemeoKiZ7ee0ONG+Z98bi253A50VcIazxpt1SdofRcZFy
imib4Yx8/kGPGQERMccZdSXgtXKMor+omVVbS5wq4iqDY6Gx3HEms3qP2veH
vwN7jDbaP7TscCZ/wJkEutWBpykSq7VBj0JLLl2tggHnsbLTFmG2XIP3N+MZ
9fN2LJCA3F3wDvWb5o+kjYPVSE+fPSyrMSwy5idKRUHItVHgynvAiC13ToO+
PIldWIYWYQKBElhah4KnZdnBiiMFPDyHvjRFy8f8lXcyaOF50CkMOmdZjT/P
8SBZs9EkOsHd6txaaFkCObpJ8Sc3S32vpG3KdSuZ+t3/DHzq4BMZZD5EmG2r
Tkje1QC8CkZlx+eF7IxyDqPdzabXaJ7zwRDdktFDSqWQpMjOlZwxsUUdTS6Q
lFfss/N2+cBFbpnPVTwsWv5e7hxXY3uvHth7SpJc84qry9CZsBzgKmcEzz7P
sV+HBsE4VW4XmBYdWD8tWzIdhKCVkj4YqqJ5I1YzHuWVK9kPrLccJ1BvmZHC
vu1ZFpcpNXTlFf+Sb3RhgnY+l2KAeatUIwMod0rv4ZWr5Q4Bs7FqoOp1M6rZ
R4HJcexUrR9s7QwUnk3Y1hAzwxJXtv3jxPTUAn/RnsRKJhQ1AjNtKhflwp7U
23W1MTn9t19yCx5Wm77khxVZKVccihpzRl3bZ0qegOV9q3LGHP4IKFQPk7vu
lUOYwAA3pNqR50ZuM6qbPOmcWGTpwrgmPBVCxNCA3pz1n3WP7M9FTML/jTSi
PSperdUVyb9eQ7z1PzywBt89rJCtemFTVnOEsjDRcTnY6QoSsaAfGL3w/x6H
SOk5cKGDGusjjMiy1hXGWQM6zEx8k8tWZzBIruwFWRZml//2dugRWgA4UUXk
GNeYktgBHjvUMOaqMkZC9MNjarlsMmEY8wxpZtsEFfj6+Rj2Kz8n9TTj/JcY
4BWvXREYTig5pXQOhl+YvSe0H4U+if1wRikhAGaK1AUU9DqVXDCNb2NYtW5K
e/nh19oEqklSNr3ph9hxJf/Rt+4tMrbQil5YX6uTHGFgnMhz3z0jZI93glmi
0p3oMuf2cs2INnAwZcZCgFCrpbHzaT1ByNEkjkU4bxz8ekX/W/R7XXmN+6Rt
pUpx2+nsIGKixGVKwBQxmRmU8XUunDAFydV2G0bj43BsTZTp1IUnzQJEQ8K6
RYRZQBV3R2KvnYXQ1Bc+3y9ZxueN+1x7joeHvHxGphWP6d45MrNvpPYvq9mK
G6m/8fBBBcSLVp36RUgVRzSWWdglE4x4r3D4HL+IlzHM+AGvSuJNlGAShV6y
KO1AT7MXzMEu+BoVNBIEP7btbkYMDVgIhM6TgjQO9++YyGVqFlt2downpx34
KbV5pPGdR0n7PdcA8azgJE2ChYpq4+gn3In5HObWOC6jEDAkuB3dgeU9naJf
Mx9/TyEpsCaHT+fIgCHfl/dyhS9jmpLJ9mZBzSM0WrzQ07ZDpbXFrW8sDQpP
gYOvtcRuub6D7iDeoOUNE3Ro9vmQ7ttJJAhM0ujxpmCupthpddisMY+zEp6p
RdFtf2CxHpGqGjKKnm3+M69yDkJEgyXV9lD9z2KUaOSK34ZAS7C7zVkzyPnT
ji8B2zjEY10+ZL7UGc8TyC33HhUzj0YrVxsEluOXbHVUb9ezcR1bqT8lgVqq
amWllC3Borj85HeWQXvRpha9UIn+dh0FE051TIqfRYUBFtjAPPmDTsrOre/r
K7ZFhgmLuCT8R1sjHjxJGc59hqUfYJrJp9pYqgP1JztpeQc3aaNwBDXirYt8
0VWKDMksCOl9lFl/6mOB4qJr7NkaFzQnEuw8tBMi+0LdlPwOXn5hklc6MYs1
fy5wOk9/p4yaMzlXiYnvAStsQBiqdxYC4YFjX2sPOtdGojlFBefz4MCSHUp3
hjZv8TAoiN33kAM629izq4ar2G1fmNrVmp38Ijhl2W0XKXfy/vcZbe7Df0RG
ZnxLCqGQ5J1MubZMogq12wa2vCKBFyp/RsXY4anVMuKoNZ7roFInAsGTsCai
k9T3OHzFL/Slv4g22kUPoXjNqsr8RBViaeCJPp751bKi2H35N4PT/Di1j9IV
Rgbo93zx+FBWWJEz9syNeRRPuuU6tSak8zL6O/VQ49E1qEiBpEbaVLaxS/f8
FuDvwrXwk5upPg3JsIm0zMTJckQOWm/+jiEbQumFP3FIsOONM6tE5jNsNS1s
xf7m7WVaCGJ4kSCeo8BTcAoP4pBG2rMaP9wcu1QaMNTxcHQLNLl2M9szi1hS
O2hs5VdtC2fRx7+v9xFcpNLu6E+u1GGmfrNz1EhOLa06oR3PPUl9BaBStA0E
gF3qDGEMD2d6PxgZpK7sCx6zxT45V6PElJzhQGsrUvSTAyqAOgF6dDuj8DRe
t1eziW9VDe40os2vxcrm5zuYBPzr6HB/OMt9nVTDsLQSFzRTg4TB3VLnch8F
YxGpBLRZ01lISWq3SJfrb2RZCRVopk9MQQRH+Cp6OWBPhYOmtHjpoIgZsbVF
RfMl41PJUKb3JrCDUDhx7C/PQpcRK6e+WwysZPqKUK9GRtEaRMDeWuzGNJbG
GY3GXS1izrLQ0DcZwfC7fIdBR+1M28ipfbh4xjs3Oaiotcd9OJTQ6RpQ2hNT
GrLOD0XmcMoRJwEY6jYYWs8CKUVBoJxFZBe8Ps7/DSab+mnU/ZEuGaL4esuq
l9BUNi1brEwnH/vT+O2rAtRwkWv2MLRsWqSmRwQb/TnRuPYsQg/MJAFCHKBw
yb4u0exea3WhGXUZFdJbB6TwQLmq+3k8iVMkYR8zSWSB738/q5L0cJm0eBIW
zlO8wtzFMnioOxEB9jTLQ+wy4JUwGw8WRRaUba9d31iPGjqjEMLiNP+Ch32h
9cG2xmJFk6XvJoJz4IcYaLHDHfAXspOJ2RmhblVMwF6ER9/7T+Dr3HUa3KnZ
hbHTKK+5RDyH98asFO8QbZtlKcHh/5Ximk8eFJIEOYj94cOQKuTvEaEOh/qz
7N66f0VzwMZ126k6Nj7/QMsiioa5jZvRrMMxCGK8WaDrcsmF+relSsgIVOZD
N+aAEldzzl7G5jbf1lqyRFgU8OJkckPGm9l21RkFqNrvUMG+p6eZrTnJoxsW
O/AiddaiM+xAPeUari2d6wLQhOnMPVGUN2b3c6q+o+pgNZHFg7124raiMYlK
9aQOzJl+YbTylyI0ng3SYfb4vlxqErNpjumYIvjXs2Bqe+e9VYNDRImTjYRz
R21GJUxDXyLels/5imHW9hsOYKDGZIhpkJiVVsqHCwo5A3K6dt5/fGN7qHqE
/bAgUOUKJunsOEQ/iwb3QWNezvpjTSdI+oNq2m+WPPo8RTDSxCZ7Hsjnx38o
YD0HMeDsyErO/e5+/R1W0F90MfXzKVKLF5fQTgfOt2hwlo/IgOBVi3P8Gimc
1SiW6ROK697h3UV8aJ4jzd1qKyLAHnqMQnQfQ52aQdBpfpKOXnpmpkq4UucI
GKbVjBv/lO0LzSExN4KL0ZiUyoakGkC7bkKgxUYhuGCDqhAUfHNOAOta6Ijk
8EmBjQZw4XDDkA2Ux5pZ7hTDqlTKFTR/zn/KliK9wlD/7byZwDrme7EP7GPT
REk2g7DNL96PjII8ZuzJGMX9XPWcNXz5vGiJvw8wVQBeJpjJ3cJy8mcYd287
6VVyBhcBmySd9NGzPet38x5KvD4zbunoCSVmn3CDQnF+fV+c8hvafxaxHIDA
0MV4KdMc56Zwke/UaC+FUa2FeQR0IWW1+dwO1b9CmLnBTDreViX8KNJ6Svkm
VlTSRrwe/vhNkLsPoums2UDPoEnPXd9eFzUvVHfM6clBgYjDeqZMLYvu2T8U
QhzDYT3EqytCTu+XK/1ZGhir95mkPOG+PLqBn2JrX/9eEwChboPSnQwLgPro
JbDU+PbT5OkmUFZI0ZKd+4SWFmNipgwJs5ROl0laucS9maodIwWeYDeCE2Lg
ikaveoaga8ohACghIpxsYxqUDqNGB5+PgZtkJi7OhiuaFWGpwUtZPnN9RWTc
YQL7ZIgWjh/31e4zll9GEAFH8nN0Gm50d/kj0ihe1ElTzvnLEKUn2nILXLUi
xjmQaJOZaCozZegVH0YYdjCbKvfH0NWK/CPjZHnCw4WreXT1tGu9P2E00bTU
YzxhManYb+G7lhWd7i97DoNcLsgsIWJUHuqCYyjM7qNBO/ysYlRzhEm2Vrbs
XzrG/U347hboQkb8wdci7HXu8KzXrOgzQW/oWgydUgFhgxmIYRHvGbgzdEI3
pda0JZmdHW/uTt1XrX6pMGuJXKfxXc0zEjFmRJVtvSUg3e4nUeR4Bjc/TzDK
hpudLXS7oCdMclIYqkabFo/fJ5eDIz/sNC+8R7tejGNppVad+Q7jw8urwPVg
7NhuFY/c7Ij5HjeOm6aK3QoduCVcoz1Mp1s66SCVQQWhjBFYzxfYynUFbQTj
Hc+T7nghbxDu7aM7E0NL45y8j9Zx81QtPkg+YBPq2e9isMO71FA8r9GnZxKy
6GEs/CY4bYkPw037e3wAN4pnu4gYXFnfuLARTocZip7EVsmuJQrR4NOXtdjM
UkUMJOp5Lehxo9OW3TTDddCenMEMrL+JtC0XmHDGKJMS4zFaTtbNZc+5H5hj
tKvBuGuTV/ttuoP4T1vKi4OcLMYdebpe6JDTS17Z9ZWJ7EjOXuEYnVev5QnP
00+Vf4kPqZnK5+ly4V0YfhBbIzomoq4dSBZLwsNmkgu9YxmuPTDhIao1At1q
CPtEdDW4CJ/kCNOOene1+sN7WHeX0+IcBhGSbQP+7TAN8iIrh9viGu0/JouL
BKXV5gN4yX5AOPLL6cJMBhcH35PRGXs+eQBO6ROgNQh4taDiE4fCrgyixuay
25IVfqcykVsUikg8SGwJ/sja6tuZtQ0TN1Wgaoh0Jdqi3iHowsavoTSrWnAa
zw84mVS4//S2LpDL3HA3ofTTNH9+fpLcHiMXyyuid6vnfzowe9i7RIR/eWaj
7H/OOG/uzWuWdVfcpwkAshuqj8dsKwzJPHWNKwUYajrAJVmq2BXIBtrd7KX7
naggdo+dtvIWmynsfjG4+DdIsI/mQ5JnR2NNEK7pICfi0CMfUYVy0nQf6d/b
bFpfPKtNdG9Fi+dcpbNrbxuqftrK2zFHAdv+iNLUnBOQcLQE5p5ofSdllFPL
EIUccwLIIkYfFKknQledt24SPjlXR6NZz7my5MXpmMMqBOEPy8viWYZBQwTf
9YSSZT52WCCHqnw2fjSimTWXcts1lMNgmRAkAcaV9/AUBv+C2keOv2ghcANq
yh33HdbE7lrJodbpyF/oBVm8ojd3b88PEQWMGdr260qOCiJ2mx2spfUQjXml
cw1ixcF4Xa4YyE2codMR0vOkTaVGA70WjkvlbuwiqGkvP7d4Aa84FRH3dtLi
5bYXFv4HidkQI8TzfuGn2gWAAzmFFUMCCnzR0s2+QNNySNXed1eegYi8/jo3
3BQ8aYAuuPR9t0mvIiH0QTrTTRSP7/jTpKP6wPR/cgI0BEq3htclzEvGGS4V
m+9I/+Uam6K1ID1m0boxJ5dxVZommcOpJLKnFOEgRnYqjlDRmhb5RaoDnSBj
ohJFyPXpRthP7NZ9gqoKxiBCBrmXVcrio9vGPK58C3vGHY5xAYfPyk8CbYI0
uOCPLlNWZmCQBDhM/SZqOsbFT/0ijI6oriZtrfLivR2DJ7GZb9Iwn0yHB/41
0a+Lg7avPPEFQ5jXsJSuGnQj7bdJejaKl+PW40bIAZNbechEk6yuggdCPghL
WsbQUgVsG1po7XJSYIKa52zo5Yn7bHc/srqAX6r79sqizJRh8Oht3JyfnPhk
3rbmgKnE6mDAn0SztP11eaETE9AvnQ7e6yrOnncWpts7Dp5wQUuSm7iDfI4D
QzUqI8/dCXIQSitGuFcDTNY5UMvtn4nauxsL/SbsuxoRKlnQOTePkkGuEL6C
aFA4xnV0+AMETheS+I5WDRp7v0drO8hNLqimBzhy359+Z2EGjj8wSpQFr7zd
Zd9/BTal+vVXNoYXNmBqwEv1Ax6r2484T0cOcHI22hOg4MgDUFHgiDpnscWy
T5xdAe8wOEki1pgG6wS8050O2OLbUYpmueU0t024+wfZWfSCwy/d404kT6SR
JYj1bviclFiAls6Ha+iRoYwIoEMREX4GDwIjHHdb9VPiR1Ir1R89Yv7ro04P
mPolJuZVo8171+/cZpDLXF2ggKPicAXDENoUhmMZKpNoYgm7knF5VKKhKyPB
Vt77e4nmhnIWJVE2P3vgAJjrs8aKwaXMDamCMMzjvbfDMusPzg+8ms/osW3H
4cF0BNO9NMhG2Y7GC3liIhY7HXo+4RfI9kgQjNeL1fDvljj9WGmq6vuqOE78
hJGc+n3ijmtx3D4sEnR50bcFo/ni8aGT73hzdpmIRc0hi+4aEkyCDSgH4+TW
728kKdTXBgFiPg3gU2cnQVjIhCXDMOlPEBMqQkilDhBX847uira1X8lzBACi
SKzFHDszQQ+btqXTiPJmifRXmeD+RakHPuVgsikTBWCyFeEHv36fzovs01GI
itjjlYlx25xCzvd0RE9cjnEJDtCZU+Xg9YNRhLpI8lN9P4VGkaIpcrNPaGYh
9ufSLxm3/N4wsh7hNSyNwfjxN7pMruVYqZQyhY7EcJJazmWHfnQduLdtsygp
htD4aB47Zj2W/sRl8MKcisSsItH1tmwCUPi7zCH+5bnk/AWYyNMTdd0BGdE7
fctPsUJGI+fFwFQ3ZpW8BmuK9SjbFgiAPYr9CqBGkSrTenmSQMA52IWklNJx
jVVlzY4aOVcbG/DI1AhhPelt5TGa+4/PNEcDc7OKHqyPRpXDvobN7jpepEQD
pNB2fQQqSnh3AmbjVoQC6Fkb4VEeF5NRxSO1QHs6FmA0d2K3Rs0abn9AjTBZ
c5XNC820OUxWtQQ81lj2PddnoBJuiqEydPtGB3F+GjI0La8RgK73rBZbPBFE
lFAeXqyDittDNUIHChv7JkOpwqayAO5SH2O5iSTFhh5uEC8PD8adjqlhpTpm
pWsPcDBQNmnmVFcufMEORBPvFfZyXi8gQ5x3vbv1wLaeLdvG4BEoJSBuoTeq
PXZls2qG4zLxpUNeb5QabPivxbqAQy0hGn1Amwk0UI07cwDU2AJjI4rOl/Ud
f7yjlCy4GM+Jo21TeB3IKAf0TvEyvG+tP1vmbXmO40DzliVKPToLHtohKnpd
oWp/RV6LiT3Ael1RlRB53D+eV8iPQRKK3pWzo2RCtjQR0JZiOP39qtBFxxqT
1WG/a71z7UaJ4gXZ3pP2FEDclnXMzcwMKPuuY4cM1HxWGFITh1ocjHM7PsJG
cYL9dC/ZLcUbVkRJ2iNJoW6yGhXHkk0d3+9W+TXPRpwkHuoDd5u2Lco52rZQ
QZ96mWQwqNLEm07RD58DrST1gFImt//iYKbmMD3aDRxUYFkv+EA2w7rjAVrv
lTwFyOTp4kavR9SYTFiSZBBzD2cxk8NFf4STfgaFQ2Z1WgwuZQuOXMagdHCn
KJTjBcYgP2wiE0LK+Y1jqNY9dcIGY+kiVX66YyBgkxZxOhRLXLSi/rDJNy2w
sy8f/o2iohRL4kg8WRzK/u87adbx6Gh7k3AscaOkqVlF64HsLxncDfFbMf5l
PuBYL34K9P6OP+bO083Mh0JowiPYLie9JhMMV7J2TpdODq6Xou3XZkaYDolK
gfQ4J4B8D+WaWxwP9+v1lbg7KCJHUnDEzdSREpatAPU6TgO8HtLeG3mFsnR+
rBsbDj+H0O/bLMrjUdFOYvrj0J2luSqccSFwk1uSts25mW5q+uZCpfh1STyK
EWqwsFRPMHcMI0XixG+BNc9u2gN2bcQyr6B5PU98cMDz/yr6TtweKVxQ2MKz
KMgMxzlal2Q2OYZ1jRB/uipqcy+5ELB/yXYP+YOObha7BWQ0yvlkLHhpyOFA
I7WkKaEH0b0lPhhjUODPiKRPliGLSQTiGCpnXfoNPFsyG4fpmK4LFj8DGnJz
ckwkxbX4B+gy7vRPrXS9K+kOS22DYxaCtyC065NZbDymK+Mqs2gGfHFNnB0W
j8n9XqAQGDS7row6DIS2UTwuav1KBZtTj5IgTjyic/0TE/fxmwDZ7MmQpswC
K1C+V/+hRu2Vq+ZDOKtgDfgzSCWG7i9aKbF9UYjO11mxw9byQ4osMLjsLb4Z
MzkH4uJZEXSZG7Ow6FTtfsmzIS8r9+v2/KrOrS/tQX9LR/Ju3uStPGNFSchQ
5krtME+ooJos4gB8oL9PkCv+qXN5rUGxrpYKvZGRj7+LMe50GlUEtCVI7J8C
OoNDH/iwABqxCGkbxCDa5dqlcQmYyT3izSouESl/baVNNIyeX4SD90+vkr02
emKLMLM3n4VujEuOTe5jeAVxzU8q9boixIGAJoETWB8tZCWZ6RlS5YZMI+6a
5Xvf+2wrj5E1lrcTei8Zbq3Wq8uimUiqs9pGuCt5hTP/zv3RKCXtJYhC5yvP
PVYXf1w6puOjwWkh9o7jrtZACj9My/Qy6/tQ8QceorFMdD6ENkZzSvdXrGdY
FxuVHOgtcJz091fo7wmYyNcIYV9coheH0gjXO2cruEMgn/tRa5+8oZT/rttG
9U0gR2M+BDOMhk9ITxMDkb3ON1ZAwzIfmNj5UN4HIMT/JMmwwMcDeECeRmmN
Ehp4rHkKCRNitj4bMMqj7ZwdzrmR+cs+kMDBSMbWEzDWVTwnk8OG1O35AOh7
lS1V4tiSMpjbZupsGLQzuN4Lr0lnCSQYD3YTLfPh+4usqlIS6WnHXOk26XAR
3crwdFQXvgjkqndDBzLvJ63XKZpUaqxCc+ffjgd723LwHEURnHBrVik5ocvZ
BOr1OlKlWIMraKKcTvXePCjuY1XIa3sIDYdFLlqw7Pt4yzjiIIft21a9GMK/
U1zJ2Z1la4zonVXVWN5Tbd4zTdeReYtz6FD4d4AZXdLXt0ipzPMI157Pg6eR
Tb/pn0623smarFLttF0GwzVlx3+VWTHHrZxvL9AmHSGTXcDiF/E/l5CTq2r1
VB3aFz0isLbaRztP2qeUg73WDMh/1S/2EqdhA4D5YjWY/k7M4c1Ayi06K9dz
l3ZsuQUCcKBIry5tC08goq/ickR4btdKhTVL/g8tLcbN2njVBV1+DgjfbZvL
c/C/D7kZdjxr8gmxK0Xut00ifAK4eNdyEL2a52qdrVnhDc1QRHCC5l1beds9
Nnjrnbyh9OzF01y5LAf5oHMAE7N2wrbm33+XnTC4iYzSK4YVJG/TvsVnhDIY
dVsa9wGVIWDm9nqB6uJRXZKf0fXf8MRCM6a/RrJU5pqEbJWhv/nMz+kkvZPY
wNDxfhiFHCHG4eWTh4MJsfF52rGnvFZPsD9QxdonZFjB5bvLaPyWGmE44vg7
tVPnf0YEsSKyEqlfwe+cxvO69T/20KGbZRqC1/u29jKXDORixiKsb7j+Rjhq
2J/zL8hb0/34zWOYiLce/3mMoBL2+995jDzrFc3ypSpnU2gwPw6N13cIEHkk
OF1NPfmGNh7jHMx35k8pGRjw4OYhgVICFsgBbQ7HRQl8S+bjs0A4hLzqo5JY
VKSmPx7GF/HY4ZFac8ET57ReJz6pL2yaEEV/qvXCq96jdXDkDRUzMm6vwoCP
lBi0rolNRpCFKqcJo368h4a9HGGIROrErz0e+XiKD2cUwiB1m7zd6UeQoN8/
zgVhgtBxXanuzdoDHZBzwNq0O7K4lALNpg0tdHfTRsTCvonLEKOfi1f26fB9
X/lEboodE1GKPX4Eh4HDaEWiXgB3FUjrpXoxaM1CrjDqUHoyyeon5IYnmOxK
XcEvQo97trzMAoBofXDPvqB+UA0GIan/OSQlPD0lvrIKijHIksnho+nH1sq9
ton+1EECEl6W/KUqyFH/Ywb0DMym3BFj8vBYnI9iE9GfAbi0RA/V1DcvDcXX
lAnAKpjh89qXcbr7GOKmUBOjnAzYZ7RxBT38Rk0g6jks4aSmA/nvIOKsPI/i
l9lzSzJNv1YnQ8bIjxQmV4XyMx/iR5JW77jPRFxmsPRfUO4JuzLFmkEbGXC1
pNmK7seWQ3s9+/gqOfa8Ut/iO3AdRRAO2tORyTMhLEXo8RcuiphS214TRBXa
tycjqdgHedL5vW362vlodu89HUSqNADMG6mE/O62rPEB/RyMk45ueKQcy5Wk
LqM8WHbxFY+vWmqrBcJE3YYozkJcbM12xDevIJHk5Bk0/FnpiLfNQlx3uGuY
rGJ/0GDwNngv9sz16jwOCs6YbYVp0rhLnQntmI/Kp/Gf4HzTI0wLQUAHOAzX
bXQKsnk6k2hvLa86udDumuHM5+FqxhMG6uvMzzrs/BdyjCKFuYiVMV5G/h0J
Kz4U2trWyisK/jcrLwrBAYybUR3Dm9iV1uID8/uS2QFTPUGYGBfQk3uavMnO
2ACXAZmBT+qvDj2laQu+NgtYT/vmpoXluJrOa5HogoS8oycMQyBAPy2mBN0B
HyyjUc5xyzjvdzdydGsmVAEB4JaH7EeBG7vi7Q5t6EIz21MsrxiXIcCkjmIW
B528iUVWkFGZBfQpCvKRaOnGz/Szt5OwuC1QX68vGTMtgjmNq8t/mzaXGwoa
FMc1RjbDMjs8HZoom80Ds5lzWI2OLVg6plOpBjXo4sQjIOw7P2Zm1/yFAGQe
/CnHeDdSKyf+DYqo4WszldHiGdoZsQGHRJ19eC5BMeXpI5IWxQLd9nDN7NOy
5RCzV0dtOH9z9ziKWQXCCjQYDR0cS3YrHmXqDqD0pIoDSkQuZ7i/9a8v0hp8
9C8xyRZXvWi3oVz0ay/FrrzbjxWrEmn6jpB+9Nq+FU0dR27lhPR3EBJSASt0
5HnW7LSQD2wVr0S4FMrrCUen7vaXQoLNBUkII/xlJjFZfqpDBu7+LwY0IppR
oVFWTuD4ySvdGZaYE2sI7hFakS4RUgRckoWFuVkwWFLjXw6qX8mPnVfw0ASj
qU7lxPyWOHoquUeu23fmDDH6WIpHJ4PyqfORt2ShrQuVVXJW2bzgMlfzCJ/V
wif/2BCg3czQ8mPL3dIvh8v/A4KmEJnZVYZPif2ObF09v2aglpev1qT1oTFj
A8bVJGgc6h3bYU9S/oe81c2Zb1bDQRYGMzMatusymBjXv5x1m3NnjrCxmHOa
dfAD+T1QFa4+JEb1CCQjc2UgYUgM4bAaqojClDkdaOvOGcmSZVSV2/s8LKz4
vnmDgZ/ykTaQJInwl9jHmz11AMtX8R0VdVWq3+gvi3PodSAMrTMbdj+1vUvU
E5TO5LLkcrxmNT8jOl+dZTmk8p4byw/8KFzrk854I5b8ROUJofFeYX8Ha+MR
xez81DWN9FFSf+NYKe3LCN93TLUv8GqEI2fESGiLr8x6/Hqn59R2ugCkrZdY
hZIiuk4jVUZfz/Njy9IStg0B+AXXrsmdrHbhYodCLEKmUwwaLxHuAB5YH+2T
woPF1nCrzn4wD2pEOGmEvThrBxtMQWcAY+6qWnaMeV0Q3drzmlyMw+b3EY8c
tXkyjyhmu3qt1pSNqG5SS4djI7lZl7np1RwdCaU/B1NfkX0ak2qNs4aFNYaf
MEQ7h710EFZ+MsrR4I7JH/F/fAzi+qZVlK01OBTjaIo9DdzLH7Igt3C/P0UZ
ViXX7a0BDuYgotC77lK3+OC6L1goti/lBvYSIoQ9yyECmMmHXLV8bRY6yFX0
eLNasWWOqNIhGP4UUPXfckjfvMbRGjSCnutY+JJVfoozKq5HNZl9Oi264k8W
dytBXHjbzNWllji3m98/00SEp8oI7pnp0oWyp3B3fhuuIWqt2OmYoGLBuejm
IvVwtewYNHOKp0iQv+smxMlwAHO+5qj+sHv862Ok3idepph+qgrzxyUJhrcz
Rf9fYKsKxE9kAHEW9F8XY/KocoWwodrSdqcBxzb8k0wILt81Q6c0Euk9XgCV
SPfdP40ivZBwHZZV6iWIAnS2HZcWw63vrcgBQiJXwSR6ZivvOA2E7VXsq6tS
87FeKZYS8fTldQJOb48cbPQ9lx3WneC9f472VXB+Sh1qpSmscT6mM6lPFcKk
wWpMYw3x0/NF7xqVu+sSLk2TSuwfZB9fDebaYefSuA/6UjVx/0Rfotxj2M6q
NQgXiKWlIOMJhljTCW4qEKHuUuZYzlriC4fd+CvYhHyJoLnRxJP6C9+GeqVi
lypYqFrSOFy0/biYWBNCtDYkF5I5WR90Y9ftUGXuIsb3wgSFSEiyievfK9Oh
JtS41bX3OkdEGQtcax/Nvuz1uzppizoJYAyUCPERo+Ci/ERllyhcFIolREkL
U61zz6DSJqmc0OIy81Frc7gby76/ftwka7t8eyYiMcXJ4k1BYzxGX3TzjiBY
AXTKh/EE6p3+JQCox+lFchwvNvGD7owlyABey22w7spbWNFKj+KC2AfE6InU
ei9XOvVKA8NlSCwUyNTsfc5yNssMGBnF5W9x2C0H2Jda4GE/5LNb6hg0y37r
o6Az+9c1vopd8PXTFgtrc4Emot4A+YzAaXy6Mug3uDKt0zs5mY+ggLyufhQJ
86oIsYf8dS/qorVl0ZXlLZtgMOPvppZco/KNqox6jXTnB4d76SlsFrmfNSCI
MvpN9rO1LqrA4d5MysLBjmQx6bBuVv9RxKzTWeomDRQbMy6ao5N5MC0ozGJZ
fVN9hyYocMZxc314v3as0E6eamHR9mDGotZgUOYOqn9EH9hLxnoVGVLY5svd
fikAZVQz1p+kN3+8uJLj7bWM562VtUpBhQMh/21xOLrT1fs0LwA7c19pwNgd
y2hnL0KkAlgOeIbUZUpqGoUJyoSnQBR9hyOjNPTpWn8F9/Ni62JP7x485l2f
7rlcsc9ch3eBa+nMLV/SGv9fAW+wgMP8u8FWX5VTOisuJjACWPJgM2ulx8p5
OzE/T48NjvwbSwThsYo1COa6qRrPzL6HUd7hw+N2Cub22jG/h7+fErjGS78D
IkGVmEzS7Z6RIChWzMowFQh5KvTS0wxvG9HFwizV+FidgicKvUd8HrlELSgc
QGEREuE8hIfHPISrYSEB47D97J5r0M49bZBdYSezPZaMZHJJIP9NcXtCPz1n
RVV1pYXZK0vVBQbwOklui0mJ2aPAFK+Mi7cdpKNejMSebg0MAlikq9X+aJx9
JXc+tEjb2wuZiEnnl9oL4uStov4b+I57yeo2CyYmXlu6bZxl02xxDF5vZQO7
T9nJw/myNH4AjKY1PNBNxySRR9DTEloJZNn2UF0G+AEYCBtgcfl40yw9W231
XrGNAPI6jpxTT3TfJNJssKaIBBusLJGx0t8RfjKM3Pc9gyqUvCA68M50pi6s
aK0pHP9dxr4wEJ/bpCFxAcoAPCIQHeCjno+m6Z/GAlgvwVC5qEAskoD3MjGf
mHEXNeYMyr/B+e82dNvDMe8S3gISSNkNJqjhA43z7qlP7lwG2BAv/pf9zN7M
Cy4X47fKKLjNl/1la/Y7lUwxeR6qeeXR0clvelp9obpyDD3MWX41R1JzpPNa
5FSjoGQf52X9bp2Y+yKlnu+n7QP/Y74uPymP2puLJfIUd1YdN5UiNzvE9TKQ
uFEOn9fkom/HMI3LIL806/Ug7pcrEr3AdspnqwwJIsuOTD4YvPZwhRCiRW6V
dPe7qE9/4Cv4ZgfBN/c4cbNUKZIMsZcBisrTSAhNnE/cCTV3NRe6z/EbT6sO
0UfSX1brQ/sAmhIJ2tOArvioUMHIKLMlWyJasdJRgHS+pmfKW0NMrqEJkgmZ
3jksyS8BKtJ2XBV8OrMwPJOzdl0p+1Ka3XOy/wRIzLqbVvyvmG344AmILBAf
0VKI0OfETzum5tCKUIsAMbXW71XnywRvXaPKXXiyKhjpKuSFWbc5ISPas/kz
SqpS4WcA9sawRj9s9YQ0AYaDkRCH8+N73ymPjjGk4cSk2FF9AFsvJ2FTiRkt
Wrw42VUGuuix5/ow4K7ppf5OYhpGH6FriKexHfL5UBLWzCQL5c9ceBHAACv1
Qc+Kz+CG99uKudflMc1kKblTj0CDDqd3Z5hRb3MuwGTAmLm6LtAk/WCCHiYG
j+o/16XmIpWT4O6zpr/eKcu/KIFwMs5GJhv3tZzVToi73e0awJxF7gecC7/O
2FZJa/4MRZeP5GPzuT2vkRAmg0twTwZFVBUzj447BOSdCWuzAxAIZ4t+unb9
KD0v+IDZLZ2e/xAF7j5ZTsiNq7+1zF7wWMOcboSIIKH5QCqNERDvWNQE0m1D
9V7K9Ockw6V8AAgOvIXVM15omuaR13ARhfHC31M3ymRQitcZ8F3KGjn7+pbY
qrKd/AAlIVDwObQwWpS/cPSZXNcXBjNeuxPfSxdZpgSP3T1PMAFBBxXJbrCS
HRa3gPVFrt/yVrScM1GU2xJSI13K7yGFeO3eHMSvHrHgstSae3T9TR2iYOJG
/9dJPxF4oKP63f7lZO5OlAMRITDmmLvm4HOK2VgYa02jMILDa2TJZ4WX1SMy
3lefgJ3/AOqaYE7/GYKlKA3UVtuKZX3tN8WJVqlP8vhCvZ5uyqMeuZlJsgRP
ntg0KC2LKTaarF5cUhvP76G2DOiCLPfo2sbjQaPQzmsngjQRrfa5vYTmakgF
a1liqaG9r0R41WsOBuv2HE2nxddBO5HG9cMmgllwisrZBLwmoxjnVgRyVY+i
e6a2VDmKUC1Kp+OH9jXl8G+pyTo4UwnROVn5n9RPBcCQL4o4HUYGfNV6v0LJ
RDh3D7nc8xzzFJZ4FZib3XQ3b+TodaURvsl8CIjktq7Q3ST26D1rYq7VAMLm
Tz5eIgQGbVbI+mAnA2QfEQU598PgjoeQRS/dgDU5mIcPSSyaM3t8mSYRCHv/
vkZR7WG/uMHHVYRhkNST0BXSvziIAO9bkk2m4DWb9Y5UZkOgYInP7xEMs0BO
SRbPfvzrF4Yl0HnEDO3paKBtx28B3HlLQvkPFx0bqhjU1yU9mdL5MRZ7WLPc
h/Gd4TQVELy2FUSI7TrEeaCPvoxOlFQU/7doNx9Rv8+uaCWrbnBnaBh0VNIm
zkigVWDNk06VMEKJK2VzsqKsYGPUjXPk5VVVDi3xCVkmsS7gfKCqiNmP/NzB
BH8ujNphmg6Upim+wfiv2IWO/NJkU7ruvAlVGGIpvQ5lLoihB7L7mq86uHUY
md5hfiOuuYYvklcEpQ6gikRf5B9Jn2AKJ07jGXDAjlB+aF9eCLxWRr60YdO0
bOOwl9ujtlv8dyNAe/3nHqx3/FzyUhnfsmjiHJP+u/nqj123Noqu71w0AE96
c3zeejUKH9qqoV+39syal5ZqttVv5rSD4iTYgMITcuW+I/AvCkzV9KzBSc6R
NLyFPENlY00qmoyRbduEwMJ2YJtdJnGymylNB2SEtUFkL/0/IZnJ7YpSbXXF
jsV6NnmPXgeCG5279GeMR3OkrEFEm0hNd11vs0gDQwTmP8ZNN8F68kwFWTiK
wW3v4GZlrm4H/jgbJmPoA6BF/tU0BLf0jOSKwxzyY6rbhkx/OWoHecssbqFl
ZYlDVRlIMPwtBeE8WVAat0vrTt6H3/9CamQhViozDYN35Af641ukHShnbs3B
ZEJWnPwXNU21rqrSaYLU4DawOYfYLOy4ppefvL/tOx4iz3S3G/+8QCI2HfbE
5C/UUYvciNwjwnNIJtgNo+E1z0H3zk9AtenZFVpb34JOi2nFDY3B7P5gPs1L
xQbNaYItw+NiUyx4aSzmvyjJc4k5nP+8aH1ShyqygjdAl+DKrUvu4M3wRCko
RvEv5SR+HQEeCo/fWuMGbsYLvLZ9rr9j9OjwlCXoLQdD+1//UUlwaygvhsN7
/m7yWQrRmkDBSBs8NLXv+1rCgLTCaQ9qjOLOb3d8l+W+kweomyHHyGPM2Nlj
rtL1Dct27ysj63W7bhJxx+L0+uLmZ9wkYqkq7z3bsTKQNtY/NApmbHp0KK91
1lT7ZaO9GHrQMYyTfHI6/HDZI/t+zRTJcxi1n+1ul6r+1oMPmPRCN+4nPxhh
FX440khKajkJhasEVlWkgOQcuYlCWeE1+Ve6TuBhe90vTukUJG9ZFe994esi
lxs+4ZI+B8DIpiEYV+vB6b7A/sfSnQAv6iGpGtmZJZv0ljmdok9GvlB9RybI
XsqqTKLhr2yTpBfizFfK8rBKe7fKY0/37zG0dsebI3BUFo4wcewnrSk7DO6b
Qjt0YQoA18MtjB4t0LKegO9a89DEcojFa9JVxy66aZsxKpvX/zJ69IwKiNhz
JK9EchO8pOv+R55i3X4jfSLWYd8r12gsq1LfAm+GEhGrIs9S1X+qEQ8v/E/7
Dc+AStz4KvR27QLZKsc3sTt8dTLmSmBKdc4oUg2biKS+XGGYdwaX0PnssNYE
DmDnyAN2O9pqT4zBSrZFJ4GBBNZDTj2II941zavOaovDdW+zAXLbTtjt09kX
tx22Jh60QD4dl16ysmAAcZJBla1q8SPfYngfHN+x/Jx5oCoYw0TqDYDDMJRK
nG3vTayzGnr6O4YoHyEykirKWkGXJOGHHZJ14UR4Q4zqfJu/yuDHhrlEjxM2
M0b2v9IiuP8TGL2CE0DNeoNPlLmLV/rMmkEcKloO9eCHPrm9bhscJYtsdKye
Ak9GsV6jpyK35GXG1VH0yyag7rv8tiwbJdrf8SC9cm6JX/BpPMPHqtfAY333
FAduHFWBV8NDcLQet53mN2TIxcQ7JRDYd7lfPpbwC67zg2McK08b9qSPG2eB
gPHBuxcM5S1YztsdRL+BBgS9gt0yFVRSSwTRcvgvFCksADye3fzvPrHNTFH4
HLl+t4aNE3MMTwPM9GUEnWSGJ2OwsvF1PYD2gLQOUpy7Se55RIaDDpVaFoRC
+qOlt+k2o1mp2zxE4jiTr5V6NtLrgw+L/UyVIgmvEUyYnD70ntFET/9phFio
xv7b4mpLwgmeMnYfVuS62/bLpKq0upxq2FVz4Gm/wp2z4xo6Z5uBBUqKyhM+
2oqtm91bffQ+XF77G9ISdq1T7LCHvOU+WXWpVkJYwGfJbIdmCgxMHO+l1IaB
y3NIdTAlXKzfgvQLC2w062eIY+N8P18NTEc2wB5l1agIN+qmjej2LjzXTet1
4b95eY0qmtK5LFYvT9B3K2VNc9zkv/s/M9Jd7q6U0tIuEBCL+rxg5RIuc9f7
jlcHazzBaHYNwsv5s0J5kr7p71fIJS3IeFUayAywNO6/zWAWHgi7Kb3ftn6p
ePWor8qfGoty5hEv9IFmBbuNS8NNl3QmJzHfMtp4ztCtKIzp+pItbjBeHg3J
4KHjNpICnAhr7VWeg4eXrgkRxDdPgyyCXvaMlkX6hfyOsHXrU1XmrevY9Fbc
whhnCi0oIW0QGpaxU53yAcnPNeuzMKiN12s89QIf9gI3rPWnO2d/8TsVBHIk
Iu4Zx7BRL86q9IR22kVvGsneeqxAakBsm3wSfpryaQTPUmX+Od4dY5RjvGj3
5VXsAZLaIsvMsv67L/34LymQguCfjyeBR+bC2dt9YYqQsGckXA/WM7N8IDjL
IfRg2DmOkkPtW82zMhkNIX7HE6Lm5CXV8ACvYYaejX1EoLdXHdjKfR6Ci05o
P1QU0PP9ZIfBUUK7p6J4L65aXkYpLf56kx+xAUkz0SCYsJWlcMRw2KNyayif
ywCTEA0XjJko7WP9ZroVmMNvk9FK2THxWSc0TIOBh/WTi+Q43gqJK22HyrJI
2K4WAZiWc+kALgtVRNQGIPd1idJE23b8Y9QHn5cxT4qSRkDzqTUoPwj3Tg5N
IsFZAYbEoUz9VkXtKZXKIeu7Gdk5gkipSu6qaBwvYnlAb0JOLg14FsU1GhWq
J2S5W4UN0tzIuz+JiuOREp9TTXcYmlY1+NM3MpHnefL4rDPzXm/7hNBEPXS2
jrHcUJBDPvO/OXixxOehD+R9Pxr/ZJOLPh+ob1VwyLh68r6gywq7Ig47GvI+
xEnO2BT0ttkt95urPOmWuYvPKKIQgjZ5NlcZzyN6noNda4JOQ9sZcdnOsdfn
55viM50AKfl4TH4wlhCLQTpRyGcKXHm0RW72DTli0nXwWNVA92SrDDaWxV+7
jYqVUoS0TbNk7pEAfFmSIQRFhaQboxnght6FzMVB5AD+ZEqmvCJ/quhyTo9d
D4keiWjMm4ycMf2DvANRcCSCa0ZEbb7RO9PKELWa3L/SHeUfQsaO5VBhwiWj
g3Wwa8hF55yc9rlpER0blFidF2qG0ceB3CCM1ep07HzHM6sQrdwUYbhT351b
/Va76PU5DoBwjWGXxY0aTq8RSUDY2i91R4y9Hc8ZbFYHTdO6cNfMu4YOeqrm
t0NUsOxqifAv6lcbfDDQ12LIoVDxTF7V9Jff27pLAKU96cCrxXhqe++0Fopu
9Y8LbXnvtTaYXjicsCmntPYw9RZlDVlUJTLpnotjgoFTZClB73FMVpf0IMYW
UbfbE3pB8UJb+8BD5sHk4fEYLKh0/eur4BNfHRz+uZx1mrNJ7+wTeUjvJN4R
SwYdpfdeMbtNSK5LQyNl8B2MdJfWFEBtbbnC/miJvV+ZIFZYJ0stSg/asbYC
8lwG7bP9dASqMMotvtxNTXbFZmaFwhJblFt7B2yUpgu9wHDmefvUdOi2RVOO
cVysZPQKhA3fb1wSylTVekXfbpf7wfhrg21DKnNZnwvMiZDSs4+hwWFjIho/
RC856wb5OiYxuqkiWL94+ZBDf1WDs+A7v0oJxHcAP6dCHK0wE1I0fONXdcfR
M/wDYsqJDN9jnKNVWekFl50HdmWQiaQcWKk5E7BSo/Si7fObF521BEFSvlMp
Pe157LULF6n5pZ3RS78advdrV9gGoAQdgfQ9fFrOq+vIjHLS5jhehoz+zXBI
7gCjTBJ2YSOAWzr+cmxrneBYg5J6WktirGpEGUyG8yPyu9YUAuHHSAGIfvTV
RSgq9kUvmeB3w6zbffdXkqrZSeBs9aO6TmpaYbinMLfO+F40mUlHcQagcMF2
0cGho7ivBUQKsFKpMd59J1gPfg8CigIGNef+kn4c88jUh3knT/RP850X2H19
xsaQJUnU4TPcSVRx7v10P/AmeHpk5sOmFF54gBONFwHyxjwqyAnuBeRyJH2N
3VaqUsDSDCJUnhSBGbTjoVuU8OmZ/QqpXn1XpxZPKtQU0G73Z720JOUEXsHv
tZyAoMA6PoCZvNwulNlFGMEVwI/ksWIlwhNGw5RIfUZbNL0Ge4MNL3rEqyMM
pwroj/CG0kSUa6zuVjYSrsTUikdvCsGiQamTOm5t3tKwnJ6P2JzsHndP6pbB
tXbRLc7AI2T3XfGCcc9P1popyJm+yrsDCw4EHhX+yi1E+tn5ahTrwVAxM3p3
jzhVaBLi2BXcTKh1k2A9iBLrcs9+axNB6AkkbQUfOqKTOYNwM920Uho20jeg
l9ed6pLw2ZTSegjYjkD253KONzK+kkbyMiZ/WYguWVo3ygpmhOly+36cO21t
34KDel8gmEA9FII7kYAFy80zcF5x6m7TtQ+z5lxBhFysY8xSxccVzUMBSywn
4RLZUBa+SYIdgiygfq172pMdSRP+nmEsQB4JDA/mPuX1d0C5tbE4+gLEje2D
xVakFJON6FfELz0mmZYJgP4uKXuJEJ+6CIJWFkSkxARsjAdQ8YNSaFOM9/KI
O1XlgejgdDXuKhoo9GIBKFHfPpK7TOLurRimn6cDitUrPqjJLYEfoYLkw9LA
+N9r9U5ZlRXD/kuWGvkXrwtNN5guv/iiyKpyliMZAj5zWbnuJHxc9Wdb0j42
QvRIwLra4SHUV497/x9fAHXold1btKj2N3uqbw9RkbI7+DRdtIEdfo54MpKm
PCSoRkqL2+4XYwZ4/w2IHTcuTh7mNAbwkA4tLAxTM+RdyuxWiseZYf7TNvaV
eGsstXFofI4fhTc6aSb8o14nh1C23YZmnYg9IqCBKeA7p8glShFJ7FWsGHqP
EwVl5VZNBT2jWHm9mKmux6c2+Te2nO5eW6ck0d8M1fX9n1IisL35ZS3xi7b0
3fZ23JIVILuMR1DNp/97efiSc01HJm3dMaiB8AehU/kUGyMEQk2/IMCem5/f
0VOXRIksAKmw/z72Qhfr7gb9HohPUM1C7ELVAPZDx2bUfCadhqhNcIzxk891
V+fM6bsM0FMawOs9wVoRySfbgTDNHdScwv7aCyejPjN1YQio7b1SrhyMtO/I
82HkMh0Laf5c3UAv/ogVlhf/f67nsjuI0WkXaDgU3ZRF0oPTNYGXbqoCu4r0
N9o0yzi6blnF2DJV/3d2uuNeJ8wO/YaPmNsDcOgpATIakDgHifT0HYPx0ee1
BXfL+VfAAM179lIJWW1M45CgZNSaWPRcB17t2c0MOlkK7eR9fwsbCoPs7dDp
zGZRnas5AEnPbbFSY2XAxbA5QpUnAhyIjj15hUH0zl9AofOLo29znqK7BSU2
LQ68Ba9v0lmy/yuZJxVPyOMzfUXjCPuTwKcyGPrO0axJfBMJn0WRXbd+X6gB
VuSWnyQNJhoJv6P5APumw2qIIdI2kmUFI35dz7jS9RCLeaWLiR4+SAIG4K5v
tOF4kBF2jbWWyZzIM3wDP4TZW68MWdYNRg7TnVfIS/BaN94OTFXUqU0Kfpse
jhFnaHvMOIZ7lVjMLfnNJcqyHh4kdsF6wY2h3v+/JakamKuFaxED39hCaUX+
SmKnNcJT5t92xNSk2Z8YBu6FiocnXBWV9fLRzSeGiIgLncfXvN5oelYttEHx
aLq6KRuvxVF8EQM6XE8lQt2WBxObiRGsztAupZP1pPxwbcl6lEjeP+/6me9k
VpYdby4TBoRm3CDlnZk0y93NCLjn3AT4GtNx/6ilOsXplsaLkudu5YKR/vd/
BvVvFe6TPlagG/kODDXcAbtkkNttcoEU4eTP4cAvsieHWaLQmX/dcaoynysa
uwrDHavFd/eq4o++LikyEOvH0hkN39e/4ADj5ktCJGXhmruSA+u4E1jgR1QN
oGYPuqIii9lzgcVY3Yh3x+j/uODnMmaBnuuwCQX6b4rmWxeSvlpLSJT9y9N+
0NuBGnW39UUSQzIQ8Ta0oH46djYZgAgBFhMSWSuqmPS2w7yUCp/YQE24e+pW
LrF7HdhkWRXqu358wG2K2ConSFor/xcLSu2cbisKQXEyPGiDIPR6t0Amx9Vw
bhUbB+28h7RH7ABi9/4m3U6Vn3/TX/LaH982BsMOfqmEgQHNMfc7347q0saS
FbMC0D4rK6rQU/2PDidNAIuH0NjGwsepjq4kL9ovzSZ3rNG2dzeoVRP+AEXI
snz5GMPgSapsv52vBX+76gtR+uVnO1CAAKhG9EK9g13owsuo5xEGxVZkbe4B
keX95ILaj5FKrBu1jQEP/MLNivNxCBUUqWtmJNlyR43A4/BncbOl3OvgAlNg
enUYCO3ag5quoyxVsj6aVbk6aXVg/3gGRRbI8rnAy+edJQXCPCdBfERdGJKR
AD0VFfwuWobUUF5JIr0YvhBE9Me7YlqrDs9Q6ztziJoXEyaLRK66CulyI8+B
SSVXtBXru5lNsYHRBjOW/ZajL5yrs1mbv7VMM8KzzbZFvASi6gncAB+SZhgZ
zjD0I7G491n45UBg8kxT3/MLCfX3oQ0C+fMRqo5Hy3ciZe8dX/tlibBMvGGp
b8Yky6Yrg3upsgH8fhIfD104p4hJWX3MAGFUhJwjOjI8pvcfzPoW/pQ7l3Ry
OWifjbfyh2id3IN1Qk5aqPp7goinwbf9Uy3H8EXunZhyWd5181Ckwsqgtid3
2u75bf0B/dvkhLpUyoaOduBQYLBOzEPubXmVuGzzb+/NwqATaIiJE2tkG086
0VoUoYo5Q1yaXJlPVOO3G+LM2a/Yo02U+ENOfXC9w/35xljZtyo6mnIiiQAv
RpkoObhzOCJDvshi1j9lvX+OEUj8oeji9PdbS40D1BWGfX9GvDsfiFb7CVoh
iK5FOm/fH4WLcf5pMSMa2FP5GoMVf56o4oIIZ+5tUroZAAMCwRGjSTO9TGtF
/eUA7rv7LidB5P3u9jUcCs8qHg5rfJ0Z6O7Ot+8leZZKFF0Ae1oHXlrHSGyq
ac5Cpkr/j+SKBei3P6VFUil3YqntZWakMDccxWnK8o0pZSClvp5J+2IDPiMt
LBDNPanekcDVQMFX/mqwIkRCh/cfYcPa1ioyCKmW2/cK/IPIymhyijmMUG4v
stoH2RNT0Mol7+PlDBb2MHODUab9qT9ZWHs8PNgSg5lb+Q1tlRIClaRhtjC7
jnxJUCqnuCxhb3cUBaqXA9txo/QvvBWrFPjN5jI0hh71Xtwe2pX52z4udoWd
1+OC0BmIICKA78w7ULRFSEa4hgF3YkPuGunfYFd8fLNEkskWLW2tvIJ2BrBU
97Quhf8X1ny9OwjhoF/HAyEe5pDbpY8dg4mtYUcUswxxY4y7xJxZCCsM5Txa
zHMQQiQnFjlT+BcsVhOpevNTwjOJUaK6Zsde8Dp/bsgo/muZGHvzb2z+FTLM
w2ErXZ3rveSFzPEgfLNDf2iF5yLlwbOKiLw4WPiiTkWtct99Ysc5zaoLi2zh
UpdZx89gSvsVXbdfNRDGS/DlwI4cua4zGcp0KEkXUdf6NYk3ez2Hunl/0JiN
P9z3GMytC3lLYvwDkH1FyaElW8yBgjZFX87cmiJ/8HU4SmH+1uXVcJBSwm7L
FBkeiGp5PCHU7IdZjeqrv1F6d+4g07fLnhA8IaC+HPmb5atCNAjeJj439LKP
ozxJ9PrtWXQdCSs/A7c/hQ0GhL/anlKybmMSesNG6u4MONnelobWcuW6mYFv
Lh7cdPJN7MevMKvs3LujPng6bwozH8gryLLwUaiqIsIuz9P+ipYgr0pq2rn3
FU1Tlbv3LUILqrb1Y8IEIowEqklLM8SuT9eI2fJ4QFFXq43c5qp8abZG4Fzz
OiOGTwJwHxCJ3hwyQLuVhqE96ho++lfRgod+DOhytquYuwoAp7h8hvGognkM
h/71mpcElfOgXhxGJPMxNf+zkbpjm+PbHQWnQ7RWBeWebQEfnbc4FDOsnfSY
SNlKCvM3Zp9mXyFHvcw5b+EtvidmwK9KOuI/JeCJacUc4INbo5ku+TusuLCd
D4Ylef7v+J5Yt1EBQiVkgnYiGUO+fAbFgXTBbDNSOwhqpNwDi3plWo6ALXLA
vk+T9oEXQ0LWJLorFti+pylVwYGFQTqE+fifp9/jigNNW14iO2ZcATO1qM2D
EBjDwGbuYEKibuY5t4goxIcReaMVVmPz35F3YBXFoBBdJXv7vwnHdXVXKgqk
94TpsS448Dd/b67Px68lHVXLaRcaA3vTDsp6+kIb+qzSHBVTRLrZQH49jnmZ
PF2dFUPVvnSx+NdgL0lq9AoyzW/8RWz+pVP+bc08HeNpCs1RxIVJ6w4EUNlp
/+OU2/gQYwrM9xDe+8L0unKTPf+iS3NzZQqiXzUid6ffzRAiUI97UT2dW90W
2ALX+ZQb3tsEUePddLZ/VaRYOm8u+r+odKrsdcWUh2vRoZ1ShtlBohY5Xi6O
bZDwQ3Xl/vhW/kMAdkNtSjQSB47Y1zstqtJQmrLX62WQ6XFWLqCjaTodn9GV
p1GhVA1zwS3Y29ntJ2TSR+hpIOfV8SGzaHunQhfGx3oNSDtgQc9xa+Sn6l3Z
cWxi6sMZ9M3tfD/DlFfSqV5TXVuDRc12KZi09jwrFNhh/00vGZEiGWuYCbAD
EaLbyyCWMwOoNlNoK/HbLHBznyaZDoNH1lFNqGSDk4RL3aCkU1ELOeNIAnmN
HknIb2acqC6/A22l27X655LFYA5pnCoMVemQgptPr3b0emNTDXoEWw5DuLQ+
1hed09hMsFX8ZZg05Ml88T39HqR/SSmT5FR0ee5U5x+GxDqmaQHPvti/31JX
zDV59aQ7PtumwDDD6wX4ZkakKGSinJutfZgvZ161+ttOVmbII3LhnNirEBT1
UckvlEGFU+LHcP5JujJC3B3DHkjvNuO87zgp8vyzxqPP2FZC1GYWRfUNpokJ
8WgveyIEUzYz7TYwqupbqioxxzJUi2+uWDfIyf7nS24Y3D0SXyeeMsiheRKW
aH+MCl5SNJlYoHaPzA2CHMDIkgowYRJPiebMMNLTIvXy/EBlF8XapW9yhkE9
ePrIYPI5/bixabQfj/nZftLiNvB2yAe1Phg7+d6T0yZZyM6DQBOtpSSR09X3
IW6leYqnLJs5CfxtQlGFpQjbUbUlj3bYc7oQDTbGgua91Ygiqoqb/BHtmzY3
VwhxSo5oxAVJFCdqmvW0tYtRSYx4ljiO/RDTGSMfBDzdVjQQomVdqlan1hWL
gJd0EaDj9OCHVVfAcApvz6rHS9k5oORSeWyqgatQyyUImwMB8nSd4xCS/Ktq
CzjoxyDX+myCuo8gSvCNq3ZnGAe8uWZiv8TTxwWRmM2tHwGBLHOkltJis928
T0khqeG47pkQWBPJGNBZ1mApA1yJQ7lz1xIzT+747crx4cj1IsnoPqG9IaG5
EwfjM//AcI6QRwHHEOzP8rPJ8medPWoMNMt7VqCryjpU+whNXa4FhComU1zD
HCtytERtzoQVksWtfr0nXoEcGQfDXUodDh6j3shyQn1C5eK2Mrzmfil3acfU
aT7GLi7WjBhbIZQIb8wWC1qjhFQaz4eSUOBfGVUcxDr8AJmwocirU5lv2yl6
OOHCRyzwNISReajA4l37USRPUSnx5KhA9I2VGq1eWzN1NU98ug6LGct28Cfb
ExsMtRBRlM3oXSgOQutQkZ2MyPR2iieJBhAOdjycMzt2YKqTyxccNz3Em4AM
pw33ZVs7y08r19io3HeIj0ELdbEZPztxhSiDeIGCgaCqag2Aol18bdg93/qj
MsH3O7dfUqYK7oHh1pSheG0Ej9E0Wf8JbBnRBqoqeKa7DfLJmNfv8RxkS4x6
Q2rO5bZ1TAULztlz3TjIzPZJc1xzPpj5dbT6GegrkWMBTZPI/CTmmJpiMM8a
tNR1QP5EH7JAIUJ7rUO21JsLCnlW1dR3jJrzrVzBhVSj0TEfKU2uyGWv/vt5
+bnWxoIC1SUPPjKXLOm1hyXBvRRbHOARJCehSBTjAjs8sP12Yru4wJJ3yJnm
nHeXYBbsK6DEBShCxD05JRe2043MkrTc25DOycKffjV81WKvntfGKaykmwOf
8FRkYfWTw+dDZJYwUOizvsItskcjPYasK9U+y29bKKd47Z6O/yJeHIeN/kIE
CS5JA7fcBB6Jc+uAL64JfcEouKKPO/lNQ5yn150CZW5SZjZ9NEKz2qE7L+Po
C4htxWqdW+Hq357dggh6HSXNKvpNqsjz4qB8aaxuBufBjPRrmlgKbMNpc0Ru
6Qyosb7GtHhnBRggyz/9XtHXhz48xdtbaH0U1n8j1pHMTU0yjQyYUQ7Ru9h8
weQTYycMlrsYvV3geAARlIcD4u7QR0m/7cPJGHv6o6BDAMrCTmUfIoTVKyHa
uhH8sSnOAiOXnXOxiJIrh5LOM4NgWfG/r4KcFNKIXjpFKQEXFy06rvUEiDeH
Xlli7sTiX/LSZuKvcXSp7wgxx4OWHSZvSW4USLsuo2sdKphN+OWWX+lYKB0i
EOgVhxXKBNcCQNOv9XYIIqfN2PFTj+hCeDlYWpui8XkNSvaJw3PmcGeeQoO3
MenoJd8TryrjEpBh1NOD8Z7qGlZte3AuqPo9gXneArVkMhaWhrgk/NmzRhkO
yZOdi2P6fDwcVJpmZaURrIui921qyA3P/SIP4z37BY8MUIMb5kOj9VIb7+KP
xQDV55IGcLQdV2A4G6fnPCJsOC6QGqMp1+ZKOP6t07r/KF6pYVggGKTgx462
c60n0Fq392FiqIgY0YM9Y8tY6EJkI1F+Dsb/fe6q/83zBiz8pUSBLzm4+n00
drpCFpI9CW08DkutFtjhIMCQgtC8hoX/J99522SQtMnnm932gcL1e2/qXP5Q
VXt+aXuo5icw3IIlzB/s5U558JYia1bFWAcHrLRWEFJT+FJCFrGIRtmL6xH9
9DK1wCf7BXsrdDbIDuKGvTv7hMCaniDGh7KabaLeEA1F9lMmkWEPSj7ut2ZD
8EPRe0ownyzKN6NF07JVzKj52XhsP8STbpwdr96JlpQGRz8UBtS1yv8jU4u0
cXzR33Wkq8wTFj3nxfe9cAvgKWlA/jSdqU7VE0vix0SRGRAhGeLoCn8a3foA
drTQLgsO96n83VVIoBnlhpMoswQF/ATh/BS518YHjO01EdN4TfHEytkqQ6vL
9aH7OVl7FkPUhb7dR2cl2+zbwT+mST87JNUFaTCwyV8xxgN0c0sPf0j0qTUp
rmjcAGA+DDhDI+HvE3DGCSe1xQX6ENAApC0hGj4pIi5eqi4NaVmeAMv54uoD
lZ3bruqfTUFbBbKFOoAwU+fUSXcsglXB4m6/20MYuAzYpjoTIQV2OaQ047fJ
vbidOajU/FLMGcGWyVWneuWbxV6/nzzHX6S3m5UgdT3HqS/5XrjGdcib3vMA
4TrU2ghXRkWai6DBjb6cZ44k8ivAAU6/EPna6F3TxeCP9+6VopHBfzrQq91Z
32AhZDOSEOhVhynYo/msQAYvcIbjNux1JMRo/2e7Jr1hPxa0KlZlq+47hZ92
471lgyrOUqtKVYv9N5tvnxztvJkb9pkMjTtynWE0QRO815k0CxMh/RQKM4EV
JlhqUdaf1IoMJ2rsxHRUE3TunaBn6G+mL1WpD8nwAT8T9o+oWUu4JfPFOyem
z93k74qo8ZFq/tfV9S+noic9qc3Ulad4OZh33gRrH9ig/aoi7j1zYILsSI4Q
ViPOHot6XQNqErq1GDNjYHVuf8GY3mGS6HMejstQ3cn3YknQLwASSrEhWoRv
Rb5StcGkuw7c2jwjFf+9TzzDiP2+oDyrQpdibqzzbpqrWCTm0gZsceh+y3z+
GWR91Rvy2YaULC0oZzxQjCSFrNiX09uIw3/ZrWvoF2yQNySHZYEqpmhieMoh
MRi118CzZ7ENcoOy5dOORSARLEztUZRJDhrMmIKd2qoiGX7kJOvQZjqXF0i2
Acm9G9nFXq51OxJGj5MuzsQe9IIxoYXFTs5WWr0jsVp4rHYbZGWKgqUfBwcN
PXMo5cr22nzmPYoCzSoL/tT8Jlr7PZuJ+q0V1UEJG2G0nysnNTNbSz1aKCkg
247WpdvD562fOBGV2UNPAlwKT3RPyslfHfnFs94BL42uyWmo9QgUyRAd4Co1
sbSOYtyEZtaKxQR6WElXqbirUmNLsxLkNuSWebgP06jLIPxdelxox2TlLebD
5gtQYIOt5sT2P88oId4W8KKqq+/zMT7Dra8Ws9axw6R8l4CY0/Q1NtfJVuDN
LUkn0bKZlGnk+GiLXhvjFtu9dmf77YztmYwmOGmeG6MHC1v6PL6Ryr+mqZyv
yKiNEDwz/GtA4Ps/ra5KRm7mMZcQC0yKIgszsBDSK7P0uKMb0+4WQ5rKoedt
g3Y76RMrcR3zYf9F6uxvHPFpTUS7t50cjljaQwfaOYGX7ILNdRbKKFLUNn5o
NZHIdvP/oBx0FdOdFSqeecFCi8GWnZ9mbbAYe9ZPCBXeFGbsUfm9lH+Rs8Qg
Pel59xIXbq8QEq3jc9Nsy66nUEwVe1JKa8E0S6OeZygy9o5ejawAKhR8L4Q2
40Le+SEfWh0yBLlCEzu9xbkhROX+S2NC5V5EQK9CXiUjC+TBPNLSnjoUOik6
R/QmtP04/2Fy08i5D3KKR10THAAtgJbHT7Y0yi0/LtxV7TbjhcVkGNR2QsFo
HIAse6YB1H84lFzdoMlWEQ9Yp/GHOyJBx7UR+mXrgEftGFv9tmJ9SPRBp8Oq
jYKYXNRzmqBQCEHt8KNy6Vt/UwAR6D7jGmG4/buNltW3a1+FwRgClkZNS+9r
eEurm5K1onwrdvCJBDY4F/Rr7vElNpbj+pDl5cLeWkAcFX4FYs3xCH3a7yac
Rz9iaqNwwTbUdCtOp0GrAsLRwWb8CPcCXq82aDK3v+2BL6OkWfTZIotgHdOT
Vc8OsEusQg1MHh0fqutLXMXF+T1pXS0HzGsEHw4RB9G86acNP9JUiV6xW7fL
m+xXvlT8AzR5l2WqxW+Oh/iLZ1zHz8ocvE+6gx3Dm3XA6Fhe6PIjZlr/D7G5
+xRAymkK8VT/v+HmoPFpePGAg67GAX57QiM6rinINg3DiSafXmY2QWyvurHT
4Ycf51BZO+2Ky9TDiU/xmdv6DpFkxYr03Xfqg6Cjvo4EU1ePecuc/XezEzTL
QsZECB3WgpHNzSA/IEWMpUYLm2Cz2vq4k+XHyfsnnWFrWsuipD0ltyGZOMQr
bOaLkPvkBJa+QKMn5Gdq89NW2sawrnWpRG3HvmKiCIFxW+QuTnysvdBEzl2M
J/4nsCuX7wQdkUK3W5dJa+4rQvR6kDDUXTdbPXFAPW1wZBrCTJUtVb46onOa
C7K49Lm/qquRoQN7Lj7GFpMHtAOrUvuE4apVgYSulTNxpkRC5XhJA87ZmFaK
MTtXVDOIOwtGO2YDfBYkDQGUxAB7s4qcZaqOKThEBrXJggjBX+4nFcln64fa
8vCvWK0NdwiJ/hk09LEvbjBI+cJAdTQtfTS5MPXZYLFJyqSs4wf3ygwX7uKI
GgbYAEQWkdLkCCsth9a9LyJJiL17zEu+aeJcBZCkPJjxMA112G6wQJmofhDV
DhzvPMPYghoj6ml2d32pslF1g2mgcjmU0Gii+64I5Yz8eDSiHVM4hTL+gNIk
HJ/exzqMa9vlXPIQ2PQTzdeIEImBLBC6OgxV0PWi+SM+E20mR8/HG4rRuTKH
wqrqrK1jfUzNeiCljw7UHIHoef+XzKsqGo4qD6lJbzNttBvMv9U181Tlmz7Q
OqRrvpKaQor+ortlPJtKcZ9F95x2PKoPQ+3Uutt3p6WEjQwfu2OPN3UXzzfR
0tufHvyNAVCMcw9kQP+V2iXKSEXYK/ODRNUtRo/vOxnaJu5v21zB86RH1MBp
C13n4EXQyBgmIGSZ51x3rTKbmBRicJbC9wVar8hJQDDKO+/6T9RXKM3x8rXu
5YYNxBApejRaTVxNYDvLH5opfHyohmSUKziHoL3a87cABAs4466Eh3zNesy3
4xwVU61XyoE/W/47L3IXFQPKMnrDsjoLSrATaIBt2vCLWQSC58/PDW+Mkfs2
Wy0xQc5RNI1PM2SlEXX/MdxliCc/O+24hRAvgT630hdNDd1sw/tqaY28y44y
m9/e32V9RJujIAN1fyGva0Ll0eJ+ZvYKs1p0eFMda/TOzWhGpNMnMs2Dxy7K
kiBf2xIa5j+Oeoy/8+tL+RP2ysKxDJdWAPjRaSB+bu2yyqULe6bceD2r8Fmv
0oz0bLvb9hRqlaI6cgCL2r8BZloOWmRaERIkzNm0O3Fb2D+gqWqEUpUXdqws
KMD9cIsM1OwXPhQog7AQiFZE6eh8mGBT/TzU+wx6rtv+h1mH/XBqAIrBo2Qn
uJoopkPptsJg05hKlDy2KCf8jP/Tu3TppNQRrNIndZj5ugwxxtGBSsTSeiBP
QDiiMdxbKNAu/iyUqvkdAAM56ADP/gyx8yC2Foi1eNxLMUrMemuMhylhASr9
tncnS2MxKvLP6lKnXE3I4zeMzMRYvdVGY6ajy8uHtagGK+55mwvF5llA0ujo
mGfMeroVrvDfh9VC3GfLxNen+8la3wTFuvBXD2Z8kwVTf9ZsUC8KXMUwvWGu
y9L740pj6G6eRfSwyl8XYfOSvmSG0CH4+CHUQBx3msygS2odlrV7qWseTwJW
WrQfeHtDGDFU35SP0/ed0K1Y8M5lqyEsFrRSYUIaHOCB77NLhVuIKgSEEx2X
O0ZqEtxxHEpKsegtqz2PT9+hnEB8S9pe4Ji6ef0AtSotYHHkZIGEAFhva4rr
EfJihnwIrnNSguqa5NGSVOWMppDF/qFVCvGtc2sbEtnhEMqJT5kVnWNAUcQK
NNwaJAcAzzRw7aODQD8GomQFx7z7SJ7MjNXpYFp++Rc0uRnNM+QlqoQMxGMB
35KHIfIoSWjtzxmx2IjSUqbl0PvpwKutsOI98NLySRE+9YSPoMiQ5KPaszYw
Le7UNWt2UotMWd5HL/SyohD0DMdXi4QRHP0OmO2CLHmvrk0q5SXgtYfZmk8f
JEVkV/TacnnwwzXHLtLm9SQAyk2wTAb7klqTpQ6ghDpLz7/0sAlPG5BTExMW
MoFLn0r35bdOzaQnZf6BaCldrknBYLPhcad1IEJbfplEoR3q6Dnp0YQ0IE7x
Mba2YOmKgdMLfKWQ3wEuPjI3HI4e/XaDhVWzkIGWBpuS75Hh+j03nJbWFJc6
QhmuZ2yC4QaMjfY7PL+w/CJ6ELvAZy4ScUE/1qmKwUnI23bRtyOXS5vqBhsp
1TwuqzyG0moI5/YM7ZWoPFxf5gRMqOW3kVN7unHPjr2ITjJQ/1ZnP29QNOIk
WZc8dAVB/d9lLzk4P0+8UgaZd6kOHjw4neoVR3eZf2hmEcFIShgdi7qBt2km
ZgJMkTz6dp8TIESU9JMl6QFoH5/owtRgmZwFYP1hLdZeU2FnvMf6AHXtDgcL
E2Gmz8GKS6gZTaPH1UFg53/4lRn8LQg5rEmr4KFuNbsK3fnMOAY94BZoPJPF
GJLVgVY+GPlnJ0FPM4QNWfuWD/nbEPdT/ua1utDmstdSWs5eKOE+tZaicEBE
sEkMHAmvyIDGBonqaGh0cYWpdR0C6yhlNGlev+prL64lkan8EOqgkqg5ppGq
1S2xAqi8vM7KbaK/9ezteNpvBd+WPhogRyruC0qAYcRisfm32Yca6bPAgiGD
bfaUBD8lmciLGaEaazCiI7hJU6+tyrnbJgzbgMZZrdMSg9OVqyMujokI8DxR
l4/6OdKpLqIxEUb68INqkuu9hWozafiq2XshvBiWseLXHRje+p8gw6OwkiWg
8NUFqN4oSeWuCQs0T/Dldx4ks57gqf6ciM6aaSawaoRwpGOBCplCLoWWU4o9
OGOjI6VmCsk/B2qAAhGpXbErBjOA0RikSKR/kTaQKkZfjHQPe/XF7JxnICfn
PGD15fDA8R/DBfC+KUR78Pa8E/J3DKvgN3v/oSkhp2pRz8FqUSgG32Fpf7ln
p+uIz3ELAhh3gu+FJIoXMoO7nmLjTo30/KTndjPnahhf0Rn2AF1pf7vJTqfS
EKPzfErrlu3pqp/RzYG6RIfvE24Wrm7iY7B1R1pvAJc4KGWv9m9QCgRV3xJK
l6MBbAYv2kd9VRlk0UcfzphHNCtUkqyJyKI+qjuYkDuJlLKkNlR3NMBnnsSW
iVaidIXDgX19DJZTiLj3P8lEDLz6ncqSLE43jmXu7ts9SWktFJPJFvvscaPu
M6FbIYsLNIWVZMzQH0MSNN1qYHs6Unbg3BmEfSkLQ7o+BV9xiKyYpNE5QYh8
8BNLdPM6wmNzqgUOdsFk3M2ljrEzqnUc8HUHjlrY1GcSqYh2DvMOihulEEp3
ovGOsn2ou8bT35YWLTiBXtUAiXlukC64ajcFQpk0NTrIqoRoFZJMj47p24Yl
X2h0Z1rqV+03N9Iinvv7W9fOdj/uAKls29b5IPZxY7sN7ktWEONJvNEjm1aR
ekm/boHP1oOpFLd6rQ08rHXTfE9GGMP0lKz0D5/Toc1YNywlHg+BtwHBKvQh
7JeRQVlbkvTc+7MDRn326JqG/rkrvPgRMEWuVYMkhQ3qlit862vFPO6pMmoO
fcS6OhUtCuWtl7uMEligYAcG2eB2DMF4L8et1eitQHaNnRagRCJsUnif2Xdx
IAezSpYCxGWSYQyv10ylt5+OXDRt8b+7YLTWuKSutydSqZooCfchRinJpBUT
MzkaNYW+mUTrifM2vMgUyhAQNbAYB70RtOPeWL+E8Jznq+zHQ7xMCE2RwqHA
Yi9fI05R5QF/m3rJP/ruHV2VyD51lyXjBdEw/YJDI7XiTXnN/snah1/7t2nU
jJAHpAPv2wEzDTmkjViBlT5eQ6EKJBumWpVYZStSNMJF1CAbJpU2w8+SEvA2
r+OtAYYvZBhLbH8epY/1HlFDBOn/4MvgeaahZpUDdYBC7uU/QPqcu6CtEU98
q92nGhpikZl0sxQYmL2E7xJFxp1E0ylxSEt4IM0SEb0qJHa6KWq2HAh36Nky
jVxm9qCEEcKRXDhphd1V482AlbofeBhFqt2FpXhCiQp2dL+hPCoX+E5W+C9i
maTrYIpY3qyuQQQSeuUT0SmsZHyNltUh+osy0/r1vdWw77frlQO5q4T7EFW8
njLKiaH0/NW8EKeScoMsWzbUe482Dgzt/wqXnyazFMGaHphWqdy3t9oMLYPa
c7uBM152WNJQjjkdQuJvVy7++pItXtp9OtXVffbrVshU8aI8n8Ug90sFxesx
3Nu7WSSoPZDBbYQYWGbf9w4urX81qvqKU8ZPXE5scIPCYFILqMR+z626SppY
ISY0Z3Ol4DdfMHXk9cDwgGCI/iEt089/P6PC1NaCn1cIxWrqaBlqzbZeF9oG
fsKc9PbLgModV+hXcvr6EhizNkr1UoO9jB+zum2MiIKCbFMsynSWusil7RHD
2z0BX8hwYcwjz4m7GaW3DCAj+5rxjf/1Q9u3XevOMP931Ose7UKA17W7mFUP
Z9c+1n99FjxIcqftCpXMNWj4uZ6GJ7EPdH7I06Qv/CaQyzzxKz5NwZ26f5Cd
CGs72ZbfL3Rpaw5zUOiMR/Yla7s1mae0cMF43dLQsdIUW1r9eejQ1mvYnnI0
xrEjRdvkzVHLUcR3Eu+IhtQgEfrump7MkPdwx7xl/a80aNeN2lDzl7bMRZtU
xWjO4QbFI3dAkiJqYDIRizY49/2zyDI/z/9Ehwffsyfy/L7O9dvpfJK2YwPj
4FilYqEd3Q4RgvGCmBduJ/gyaX4cPA+ohI7qO4AD+KFbDZIJnOa8VAmMJESn
VIMfVU0Azz2utAMbfHsr8eL7yyBLZB64KTwka/GZFQte8N85ANQGEWGZj1za
0ABFFFKxSZwmC4OcFiJY1mE31ASVBdiuu4F7UmOWeawY7ggFQcDy43i4znNn
2fRanxXL6riwxm2sW6R7qR4aYr8ng5oxRmpl6kUUm2Je2FGwP7OMaOUhJmIH
7vfYd1QFFZpU9Ph7Q41qu1X+5uTAB+GzjHJcUC7sEYQPg9L/F7mI+8s2uQ+2
ILr2B68A6iKVFnp0Wb82Zj69Uq3UkbDnunmAKBkZZaXi2WzzvUI3MOmtCT+6
PZDSkL9bxt5JeehQZg8PBsPK6Q+uVlsZAXo7xHCoeAzOuxg/3lh4PDmX9D0W
6fwJYBBTh2lkrD+AHAWJuQtRqts5zTL4AKPtkEfNpXZNil+5I8+q9MbwlpqQ
OqKhXXeXk2F0/t95VKVfWH7E3WK6CQdyMIwi9X73/YNwsqeB5qVZCJQxTINZ
O59mEQ2xSEJriZMn23+CznVW4l/yUMyVXHLGtCCRKtvXdRh2C7P22c7RYhRd
ZJ5LBhnaTqha/Cu/ULa4uXA3M5xtK96hB+uah09ewhBRlVsr9giLxPuww2QM
Ez6Y01x8Z9w35qAnTiD4xZIMboO9WlbLpFFN4ievDBfL8NsjTEsJws6kTMpi
cZybwOJgRGsSqWr1CSHs1DsZwaCwdwZiq111DL3PlERGmQ1qZZZL2dEsSelW
IsUWUEcdGdPvppAJxnFKyniQ2OI5bN9lnd8yBtYZc4gLw0X0CCr0RnkCiU6D
/E6OBDXaiYnGe3Se6AyrnNgpWu1RiCvRpVEuPrdZSZLUgQ/PyL9hXIYg1SGV
bBmB/H7SFHYL/p+ExohMRruq4+92MTVPqAZpAzPWOHuA8AGORIYkTkX/kw3A
HLFohS8JWWD9Rk1oGsIJTsdmBhbeto8lBYOt0JtQ7fhROz4oWIXoq4PcJkQC
T3it4o+eLdtDSyKcMkp7G2zhZCOOZinMin3KKs/XxF/7PjhuTGuybjDfbLhu
hCEZBdGYqy6qeRIpuwkLLWNYgyzF3sY7zYaHi6i1dNk+r2nXYSi6umbG+zou
4YlRRWg4Y5okb/RYLTBcwq2vBEKadsng58EYgSlvP2N3qi9R1kDB/mbW2NBw
hoX3XJIaqepe0vcPI1mHvnbPt1W//W7pfwLlM+6R+6w7vM9E/uYYlvSZXaMl
PR+E0urt12AJgHvXU7i0RnV+2x/ZM4Jw/uaSuenC6vwTEkDJER2aImfgCvoG
tE8Y/fxNNTLnLFvhYFN8KrjtPK4mLucEC569AdGIrNrqSGQrdxyxGHEpnLmv
lgFfQMAilUXCNigKSCfa5oQ2rM4k1CZpf6PvnI4qO3XD2B2C+BP8F1QIX37f
MoU1esZAN2wCq37aZOFc/95znyXOqmU4XSXndCbML8uPTwTjXlwuC2WBz2Ie
P3AFuiKuWlS2qJW3mRgZzjYBIuTGeUDFm8WO6EO3p/Z4Vcp0PJY7Otn2Oj4O
Au35M9ly3unxDVMlOZmY4QzoOyByobjF2zjiM1pqm/C9VczbYKphh41LCrqs
lGFPArzB1G37/J0FtDyat8neMpgT2hpwU5ffkWdzriL1CTRfYh/RsVwgtl72
xYXlzn/zPWDmafhGxbacFjW+cxjzQBVS8U+E4MeoMT0mJ4eJXp2hcsyCdmMV
Q35U/iaTDXhmyh7oUkTvQe7vMVPq4jLEvEoKB6bPURQGz42R8PVJ6BvXt5x4
9MLDnp2MmqFi91P5gAKVDcjWGYFKlQMRZ3xzsa98n40BwGaQVYOSPcBOqY1T
HToWhWWCnl3PCnK2ig38AbalxWKOIrvqLHtSLB/0it0JXxu0gmBqwC71FIw1
jQ8fWNRi76hZ316Gxgb0S5SYsWiAZUqAMbuT0izyyurZjhzcU101FqeIfmcN
Xb3nRWtwSYi67qpxVxdg7uVAA1V2ZKVlMqKeuJ1ywul6r0Cwos9GxhyvfmNr
OMAAWJ+xJKEgT+ZXf8qJak/XFLhVQ8l47h264BoWr64eP3pYLdh5IxhUUAtF
C/eeyDsuopppG2H/PKUH+/gMFbRQlLwRkZd2voOcJUEnZzHTi4i0MYkHYzvA
XqdN5joWH1Pnfb/9bhyqthT5jSr1f3v9Ezlu/9iygrBDqI4XMj7AcsAaBabu
G6/OHwnAy1xQJN7EFduc7AXwzjYezEQGwIVB9ZAV5mlKroahScz6/5NasijE
IfHwDETs8u43kzKA4BJ6tKZOFwCOVgtiODd9Q7OEq0QbOvqTPLDoxdsrbas3
CYaHNE4ohNkepjSwlzYzZAPqPFAImEHf9KlAVBYb0VqZ3o15ptPc9E+e8az8
BXW72oVBO0jnmBtaQRDokU7o0FkiOM/UQgFGyoXNv3d8zKfnWDgd4jslcWKc
+c2bYj2AH1g5xvT0jTkBJFsgjgAmVF6kBQgOISoNE3YqqxH+TsUCbzxkUSSk
reLX0FgS9hmyM+DgPdu8lrc/xHbwjxzX8PKC4eoD5MeRVSzmOiuPGr8gtjDy
Nsgm1d2Izv1+Q8YSTnJ2gxxSTximSR+kWFRaHrZj3nMIXH5y9f19kNvUTnln
8zk9DQksYpGQRtIGcK75amRtZ3ubNGR66+yz1W4oaKlImw5Y/68y66oixvCo
K14VZewYzqOai5b+Q1nnnN1bj0IyJRgOFmrVah/vLN/1Do+O6Q1mHpAD6M7k
oNaLMteU83ZsDpagHsDhQNGKc5nkUIdciMf2+uR0F28l5Q8efCie0KY6ihH8
sWKDJ6eQQovNjSBYfyotIO3jPRk2587gEvKCKvCb40ToK2rk6c7J35bFdT6N
dq0Dtmt60VUb4h2pj9J26tKwILI4VZrs7TJaeLMOWyrZfZKj1ncpaM6coMDt
8nN1dqARwWeaDdhzsGv0VL0vyYFsgfb2agzH2EeOtpWtfwcpw3eIs3y+Na69
h+D9qwuoIssxqaQ2Nsr3nn/FdPSMlRBCMZR04THNyLQE0MLP4EU5tKzQNIPY
ceTWWW+pkxbp472uoLoSOzL7vSCntB1EQyW4IGxzhNekws/GUF9/X13ZpyoZ
h3LK8nAHoKFmO57og2W7w1/F5pW2A+uqNsxZS2IR0v1ReZOsaG44NeToLc7r
p5lzjMrA5iSqXs1Ta5Pt5S29zQa0jzpBQeERcsAGO9Yy9jNgdwmG3eNKYu4s
QZ1pA+G/wsn/geKcNJtVpWjSm5N/uMnNRtYel4DvpqpQKesI/B9VaGOJ5shX
GXnv5LcUgy0pK/WgRjAjuX3ajjvRjO0ZXPAmep0/OrIgx/OJ09v5AuVRwOhk
/5QiuB9xsPJd30L+H9oRJXVvmhuvxuIneDIydCwQamAJfVM2b/4eKEk/OeBY
dbs7dkGM/J6hKWSoPxNaJ/HeqfG0H+BtQ2UvBh8I0G1aINcM8LsQeLE3qotA
MP8EYRtRg5jwD9YeK2Qupe6Y7Pn/PbNQCN1qC08MhJfHWMxC8bC88hb9tzKU
7qw7tM2qRO1CDUTkyxsfaXJFSHH102axQ7VR/exReai+fwK0dC04MBnSnL/A
fpuvepwWla2o4TFmwXgigD5nm5SWsvzl3ykEJ/jbjz6jMgdaPISSFfN8k/Si
RAbIGRuQxR3u4QQqed+01oSe8JizJ5tcHbHSHYo7hgOnMEMVcyFLiiMubxKq
NDVdzSS0qpuMuXaIIyiSJEZUjEIwsx7HbL4xJhMQFq4wLIg9wj/nd0qvhAdZ
PLWmm2+lmCeN/c0/IFPXt3CRwNcbO7LeXlaNCvRQh20Y36IDGnqLtPgaLMko
l4MGRvT2gQKQMynG7EgHoMDxz4Il9zmnpqJ4fUqDig6R/IyWCLW9LJhJbU9M
DcItN9xvQ5OtqoKlFOxXLRcbjELbNREY9MWtPN1NBYUnWA8slgk+tiqvPr9L
1CVUjQP6cirIGvjbc2LcZNsmtaZmEUaXOLNI8NwWawt8p3HNQe1Sd8Con2fT
7N3FIoy+m+SK6lIbEtK4lCwPCap2Bxz9TDSAi9V9bEE8s4WX+COE04VVF4c1
2VWrZdrVDCpiMQx+oKFxji7xYJ32E/VMENJZ1HA4A8nApIWJzHhIZfCTHCwA
mzdWJhQXHvc7wESz/kUjRavgR9X9vKvcCAekEN4hoA4lPhWry92VHsitRUil
C+MrOVLISdCkez2GN/z7jej4OLERujvrM3M7aNiqnkal2yH0t/0GQrk/ZWCk
omcuPAXI862fqBorlAhMp6nFkXcazu3050I2VJw2nHQKS7EC4Jz0+L5h84/L
5JMoLnXBz6e4zTVRQ1ruNRTzhGFSHsLq+pvUZN69u2o4W4inNTQo60OehpeK
YZrjfzc38EO+1JgcazN7mAnRYbviU/oRXTrpL5BJn7eRzjcSuBXqiD77crbX
DH+f8wWllcu56thmtBkiAB/5VRAw7mTuO5SkkxRSjbnaU+gI/x8/jn3zjCVP
sXX9FfUNSTUsNCQIkD9tvQz3r3Y6QfeSQAx4kFlcbf5VER4IgoapTSEd/KWe
adZ5No04IKxB40N3gsuxWFztB++wa7EPIb5sS08CWMBYBpl6Xxz5IGArkTUp
nJNioTuOUFcVK+sESKLrmDMBTNL5zD83+hjqM3GmJevEjPUnT9IMbgLqVnjN
25asTrw0sPjlpOY9IRcd9Wk7Cidyf5zeQ4uJ3TCxs3SMBdR/N9Qp6Uifa2ju
P2r8KK9FHRHkFNIkHtyG0bj4O2KjykxoxXHColTnl1+iI6epUixdnHC+fv8b
dSeGgptPqpa3r//oWShxizYkg92C1HeNaobwpUDN0ONYcbhMPW9dOLeXWwKY
PyqpmONhpMVnPDdWKlQNcEeKyMQPtU4Rte2Sk2tmbew5FXvzYdmPBxOuMW4V
vOO0N96ndtuPsEwcwAZ4WBnF6OOnXciXtplZ0gHHV8hQ3LEuQYom8WPMSV6z
FzK4i00vFIs1GQ7yFswbS7+BLb93AB8i7Uvis6S/Dd4IZKZHXNRzNJj+XB/F
KNsJsxPfk1R9+cN56pYUI1PLtv1h05dV7hv7Ce1PB+o4dlm/OBY/+j/vQn6r
iIYWZJxoY5PDphzrzJDcqNMuRnHOTkPTDp3WmMjuA/XQRFd517TK8KzGwAXw
nM/ROygwgpxzlYqsZGqZ4BhVEmzF2cnta2m4uzuGy03ROCeogzvmWQH/TVmg
72e5WQISxw2JMebbuitVA3XxIyFTuZshqNgoiSCHE+XsHKHMu9jOf4ll1Ju5
usZj7XVH0fKGYZ5NvvRwKoGH7ZWHTTLslSBHt7KABZnIrxxW+ohbNx+/ZvEH
9IrFdlsP28r+ZbD0vzcO8A/xaN7Kyyh1yWaQm1EuSIWgP1MNru5TX7Q7PJmg
XG4EPq2N48QwZiHaFRVeDmA/Pqj1Ao7fHDvG4Zvsf/+M9vFPqDv+MOAUcmCI
eE2sDZ6v+Wwr1GtUKlEeWKsfh+UTiMtmd4iF1hu5LeuUyGNuB1JFrleR5ZvQ
pL0fzUB/tZKWY3e9C+aBnRNhVmm7MubB/IFDUf2dQMX92SPghSP1sculx6Wg
v5h4/kLiJtDNiEQSwtYTCwAR5TGIJs9k5GIA8/uHLaUlfztRUaogvFAAETeR
c9e6Z/yZuaLr3GfW1zP1Cs8xWmL0+soUvRzTnm7v6Nqn3fS0y1tM2g/h3dBm
26xv6XPxTjPoje1vrv4qz9tlxr6QgNoEMDwV0Pxii0TTz9eTDWu7xD78iv2d
M2FmU8Ssxh6CvznPBTXM7nbZ8XtsZabOWsLloUnQIHdBwlsHiU5mTEKUIXHx
cj0D5+QZI/J9jktc3heyomYtNYWC0FBpO1XOo20tj00gpoC0Q4oQcA5GET1U
asEXCPmn8FUsBJCzd47oJNZgF46+xMb/H5lMPrZSneY9m6ZMSQBCLQhZ991p
I5jFZN8B+oIAiDaErU1fHOMJhvKwxbjjdnsl/Z9AwdmdzrYRwYgE6kUHXUDl
n/ybOcDT3dDdV0ronLFFl5st/E91+SyDcPnmm6KWiWxD1Z9OXiudDcuKv4Is
/v7q23jUSnMGd31h+imSlSUn5e9o1787wYYrBQZl/d5S4D7HypZtA2usa+PZ
fQfzhXgk3seX6eFzZhYAfXYrvaLNk6PscHXqHoTZ83E3cHMuyEzJBaweNguo
foYp9cmHC38+0S2MWmaZbYaPeTF/SoWcg6yI7eCVlvzzxUdTe8iZhgNxiAgN
4m6DHqRAlFRwreBbsjHUC9glhsRZoiAWDDpNvdkHrqi8dpiNAvHi+qtFvT5Y
LvzGVE6xm+boFopfZ8IL6PC5IIVCiA9N9AYkHiczEBUkeXN6PLZFew9k9oAt
Wr9yHxgHDvVHnz2KXAlZIyeqVA92s0sPgfD2lyi2ldljPCXFrQn/VNQO/YMC
YN+at5LKER4NwKpy4P1ECYQQ9yle0Q8LYqwhiOXARtsdzi4RekFL4ZWwezmT
mca/uCgek7wQIakRW+dJYYHWUAr5zrlXv5kgv+1Lq38x488Puf9wbjOOYumc
XjDm0066yXJl+uTRvQkk7/OyPXe4CGPs5HA6lyLNek92zDu2KnvKk96ygTEE
tvgGu78ry2/wDVY44DIgRqPtvsFaRGHql8A17CaRcRzzRZT42bYzRi003Yhr
B+3yKWMU4X6YlLD9vOhwe9sBH8nNJc5VReXpAF3Jvyilsxd7DOWDh9jRRaI3
+0jKme+zc2wkOgVqy23gOEuQ+3YiCxL+ymBGqFUU0eaE+nWDp5U15hFZDJh1
plqJgWEusAmxSNyH9s9PV+ZrviU2Tlb+ToW9nKvzGmjOlpo5VGdsJKWG+oFm
J4d805SboDkBlLTR+fyuORLcaVgUkagjttTnZuyEnnm6encThar3JCOYl2VU
YZz/Bakq7NP5zbp4PUQ/sx6fWv0hmJQJXKGTqbqQryC8CMJJvSVqwqid8O5n
SRAGsokAAv4g+qx/UYYeVsJ9d7uCSQsvvr1RZ8UAxAQIkfhuFjEMnPEEN2bb
JmmPMSN6aalkVE7uuZ7/g8fegU8zyHZ3lhcw/Z8z826AhNhTwc6jjvgfO2C7
p7HBzaPXWrVzRk/2J2n6cUX5DaEGcJZzrQb0Y50dfzUwf6KouZ0v32vJ9o3f
wH+ZmQBa57Gz3bXTDxERi44e8Q9T/1/d+W/IXJgJjyEG9U8xPyIN3Ar1qTmc
bHJpARChzu/qdyPc279nIQAzpftjlCfx7VMekHGp+Pv1INtM9LtTe57n9UBJ
MziS4wH0fBs/hBUOrVITH2AkSifIAjXLP/qG8rG6DGEdM8Gt+7sP4SKypekm
fz/0eUzaq5L+tBn5jP6Y8A+CqNWiFu6ElgZgDT4Joqy+HX2KAePom8mu4le6
kVyNRgDikF3PTwwe2pgCVEnVffjLgIWST+YCi9hTyw10acpmcvG5he+bHekC
+R4FuW2RuAHHLNMnlKhffwqwGorl9FCT17PTCDg396pWMNVnLgRJ8tJvf813
HA2daPP/6DtiuuTlBskS+MLY18IWBqRIOvLaYXprYZ1qp18ZD/2D/0ngGr8n
9nWWzap9e6Poo+a5UnD06YO3tyXYgBL0VmzdrT2lARaxrZvFTm+w7kY/9BW/
KMQiPsR0C/5KFfUu/DsNNaG5Ywz4bLtE0+8mxCxDeAJx+xRqLyscEolP5nMs
V73asdLhdWXjOYhJbG3GuObr4Qw+CZ/byFGzZr1ehpL89Wz9E/lsszAwMvu1
D8Pvr34WDgIdVvT/RgCeVpb69R8/pk/malV36OLHFHbgha/WvQ2mkTXyrOpS
dU5jPaKjIxE/JKltEFpVdcEom48x/l8I/vkXB9A8CmloU9kAIzAN2YR/c96Y
KQt6l2Tgxjci9YcdVuTxfUMqrJatbfx+FJIfm4VfVqUthPnByOPGH6qhatu7
5nUP0aVTDQiPb9nM34PRKmjsHVDQgkg10Ehnm14uELOgg28pBNE0ybv58Kip
Y/bZTZroANQN/EpomB8kkaa7nlXJODcgJzLgIr/D2AFv7Cfj7HO08xEq6prl
OqlCp6xeEJAhhU4yNEP04JcZ/1IWOcdVxJobYnIulQ/ERlxtlHnTn/ZgH9ex
e+19gsA9UFzY5VsVzMmfaAmT0g19gXa+/kqTv3voZ1nDvAGmY0SF2MYpcHuq
yH5VfuNr7dNrveDv4DyZFQKiRBoUIYeyitBs452LvOxAkxcR9ON6X4wHRZwR
oiytUxNG+hgmzieG80cN43CsdVXsATAB0bKtUhM488Lg57JXgjd4xuSwK1sW
7xdwTCt1w2kdpkiUt3dRcri2JThEGDRxN8yWUtisKGNtViXIJKx0QZimugOf
0RI888R1J9CSrqUVnMdHx4wDijMxT500HqscxGZofsHJcDTUjdx1pLkBr9XA
Ixsokk6PnmwMBOJ9ya/K0eGWtX2/9hFdaVEzzLNv584Vnu9C3HQATrV+Yb1Y
dxjNrdskwUeQsBjHT2a/1TJbOU9zVudu0b6Pl+Z92/CnrwJn46TyO/8JoTr/
hY5+40WmDsvGRH5D94MTxpY3C61ZBp7VwEYBOgzitlqPix44JVjT9le0TdhI
GGnE1eoRN4O28GoWV5onk/LIrAovcY6IvER78KhWnoD7oqkd9emlz/sF46Pw
Fgs+iBIKn5jhyC38ofJTFq7R5oS9mP5mFKTy1dTwcnMpUNNFbwXNVLvBe9Bq
Hp1wT8pBKVlcjZ4xnqg7vTol/cGi/TplM2kEh+zOVsbHExuvmgk5woFvNNE3
NQ+mtK1JmsGQdBGl576rwc8OB1d9of3f/Ug5v2YbB+Q9s9MVXw8UJuFGS4xg
8SjD6BXbV/gI9at5z4dgB3gemzQXcbqGWbeblwcsljhTRBGfl+d9U6ejCo2+
FJ9afmS95VFwSeETJPgTFGQAnt/G9X1fRIfo1SKHyp3Lak1Z26BGvKlDPoID
bub+p0GZMFOuo4VSiz/7oYpdMM8c825gcnW6JdmGXm2FcsWl76eYRZGeJtsL
UTPGGY/kAZMxlf2hb6aq1NP+674mpn4sA6J2CUlmJkHZg9wRTd4y02sB9h3Y
4WjH2ROMslZepd482YBq/6eDi/nnK+feR2Ru/54aRe5zO0xwejLUmst0e646
664JC7FvSbY9fv/wF+KynXUkzLD1x5G9X32aG5mwbu0k1lzJCJTjrNZbv6rs
KrPiHhBiuAMB1Koe3mXks6IidhCHWWDQcglqSEBwtEyWkcdq672GzXZe0i8Z
YvSyxlhwHJyRpkE0cY+OugNmQIEVM5ROCc9K1E612S1hjoryM1VBPTf9voYe
hlpBjcmPKbp16wpHgHHyF/qoVAK54HlxdTuaxulmQ3cxb3J0krPNJ90I12b7
q7spefvemUwo2NeqaoPkMNcAzCv0qDu15M0U4JqVGFcHzi14vkJOSunHSZHT
ZYCIFvUZ3cQfnglf/JHmWdXhwmg4IjLV0+LJv1240aZblgp3O7DGYD/emM3+
MEbnyC9IFuBo4cVPHS14gzk1EtHV3TFfK5m93WEHphfSGBhj54xb1nVWzaP3
c+RgqTPUnF97ZmZaYgYRrZeGdcudCupkh0wyevI0FtbLMHV1/FuFwexhnuBX
OLtQIWzInJJMPtwGRkwkd2cryJ7PlSAmcJle1s/eWeJPilE+r68Z0Jy7Qf0u
t0F1dmmz78ofKqlNNdDSZu+1HRqLoYSpmCzbkdeGKcqsPFQKYkrfDOX8GYe+
InFEOMXQVOuz8zI93wb9zoyQlf9Z/QXG61dVA2WtKDWMro/aWhRct3lkPjtd
33LWPnHEhuZkl2quy97pMAX9pb2i8jxjJZd/ML3KqcXDiqC+QN0jTRo/sQqq
veTGfBtAIrMj7Jbm5NjTZgw0JCmaqsnE4uUpyNFt97g8ikYKkWOvUX2aX+vL
vcGeslsmlDomvG76cLSN1xy06aPvKJBpzsz5mEseQSNZgkgNt6KcC8byWu5w
7aX2sfq98UNC/IjYPcl70u8enhfiVHAKofl+01dssxh+GcYp3z02p0+Fl3Qr
VV96a409TBezq/fbOYxsnxDH0aNI7HnvH6G9f29ei8YnUP4VSMU+jES6tGIs
uPrn5/ugAzY8MW16hQod7K510Slb1bnnQcrkC0pI/a/b1VwFoGHxtcQlTxz3
xZCfHaiPkQDbzRM1F5qvZ5OxiChPcJvh+hl6TYdwKu8vrch/mfHt1s2woD0+
HyPFsmrzTulRRCJxPswFUuLXbmvQkV1FTEhJCzCEu7b7iTCXWaRwa8K8MAa6
TOGnWWMgGEPnEV6RMEofdFXg89fEMUaHLxCC6pXuFUENvs+pdIepDJn4DpNT
+ueyXCHuyuSJOmddr3FhcxVda9EIJzI90PPJ5vbtiJOFiUD361yF+trppUxK
LMwGqVs2BMQThEDBbOW1BD4NGEKNSHwp2xwvFkEydiOyzsi37cPY1qlJ1+gU
F8LyYZfxCSu2qfIvx04Jqf67Xso25hBCQIRX3ZEbCbZxlnNYzjDj5mJnt1Lp
OxqKamrc7V5P0hGsyR4PY4OQL34i+xv8m+pIr0vv4F8PjM/S4DRpzxTxdnkK
/Ltcc10nyPp9gBbLFcox77TdM3UCwF7JQ3BgZQF2srm6chBg5BKS8/Un8BTd
STpTspcQRzpdDpQ9DG60RwOh19z1D38RCTw3ZQfZBpR2wW/DlyWwxjbl2vlL
wEn1FVNzIpciom93BspulyD2cnCgSmt34DDDggi55GXWpMAQm/9GHkFGX8I/
oNd4sCwLb7HE1Hz95D1mYk0MkEm8XcpC2gvdr6yT4Fev4pO7YSWcT2EFLcsy
Gd5zHX3dvrecJZaOiaMmogY7s3WkmW9KwT8eyn/+WQkFNLro7C7NAmAId+EP
tBwfhyWpyICzM4fSVslifdbaVsgTxuHCUH2BMFyB4cBMdVT9g7BYrWLxWYfr
XXpqBNL7XIhNz3z4/YvUheWN51RJTYdPIbUsrDzg+pf9GPzOGImVsGak9Fx4
h9cNWHX4AmHQ6piBX4PBNqUyShyNXrkwI3QhCg4Ue/guPufKVzHlRb7EAazq
bPybN4WrmHOy1EnmgaI0f6IOlU99Rmg5XowEJqNN1obKSkPSshnFI//kWX//
Xyk/kzf+9HaEydoRDeqJI66zNXos2dKlrFqNFy9b7FAa6x4O88y6jIZoYGQ5
wvYUrhNoFfl/7UhU/iggX1O5JWy+rx5iGV2mHKjVr7BOAKovvF3MWng864TQ
7VNxXlfxQ9oFn4Jlf2SkBiomnVI7JrU3HU/LagEpwDU8Dnzdu5sFYQ1N8p0h
v7NI9pWQK76uI4GqGvyEKkvJ17BhZIhdymUe2uczo1oNEgAzYOglRJqS4kvR
OfPka3+Vy7MM9CtDHcEMSSCW2tE3NL1PQ27JN5cVtdmuw1XLWNWd5yxlIUD3
6NAkAtrbTEN1Ac6nz21a5KNcua6HK/s9A2UtANKEiGsf0ijhBdhnJXxRF45z
2gjjHQJjflzXxKNGeN3ANehTdNnERmXv/+mGJjuDCgvUK8dj7hMh4rTuZQ+0
GUxpkiVGcEugMLo6ImatUf0mNz6D25g9yBB10bIgWMk9TBl7ghiCDh+ClexN
Zd9vcUaQY13gTzY3tpiEa86IiLXXu0puWb8SQEG7KQLNIVjGAiFW2Ob2aNUI
NjI4fB6BDvnZYjk6gDOS0FE7ehvBAuCv74+kL9p4sssCLi90vzt5bryUPPl8
4eYzckwaaO9V0CHdXB6P3jruVjAsPQaq64GBzX3iTAh1VpAtWbeA6ON1jTdr
qKXVSV7gaAoosRJD8ZDmEKtXf9SuGE08xtZq265oZBDUzL1DPFFi7xQg0uuK
D260i3IKhiJDyPTMaZDK7ovfqmEUWWjvOop75ZCkbbC2pfIc3vHlMaFWzGvi
kVKARM3wtbbBdoz6f9UjFLvOjByAHsxP4NT+8CkMbASUn/6MWBCXckYxqOmB
Vl4cfmhb7lm3GpFSfVpoQEBIpY8y/TxcEtGwL1Rn7uFY/NXGyNeTtavw4pvI
4B328Nwjvlwv3bN9fBPOkZ6x3E/V5vB0m7F1CVqWIr1nPTdE6ZHyFQukh2gx
RCoOKxE7DdQZM/4jWJpxDMTK9qK12WfZQEurgH1nK7tTYcYQkHsFOpy7Leid
EApNlwLRm2rkdHMZYWxeQPktnfXncxyLFgMxd+d5Z5E2td+p0LA/WgwxVX1u
azKu72tfpC3bK+kGHwtu+ZzIG9+Q1+K4yq/7ix0tL1b/aLtlvXaYS67ASX2F
8uwCY1PgI4rQvTycfpW5bGKkGWJnYL9UGsoFEaR5/4Zme0oBDPCSdiuXb/kb
lRsVBiYYitS91dUBJfXtz6xndzcNDPD8eTQG+1M+cek2SkJcF/MWgpv39B8E
Wu/yLKYRJJGRtRi1DXQRqU39Y24HZ+6fbyf2DcZe0TAauanlLakwRtWbs+ar
IbK/lEoZhdUrtWGXCaHhzITtG12fd8khDegFGYkVRPRMF9gDeu7VH6dqd84w
yLymvtBpnfxt+xqBD6VXlWe7Hzj40JY+GnLqujxAy43QvjeANiIR3S/YtShi
mWqmjdyoRAWcYCZ3BArJW38vb+4fHbdGpGVwfHFNOGrTbUlpEEBKNB9gaMhd
bHlIXRd9IdV8uQmhhTe47A/cefs/SXkalxR6gor1NyE4IE42drHnggQ8MJ+i
CU62bRZ44mcxcdZBNF0k4Rggq02Ev4/5g6DbTXf1jHoRvwwrw16i/8I8ut4d
M1qNhSLhBMrUIbvxtZRpGauv4cDTfO3tAwcyeFqDJ0QJ9NtDwnMHJgtqn5Ak
P5d3NqCWcKcu6w4N51Glvn11hEwmzIP16KqVJHjXfGKBDlX6zEuzQklLiOAK
rXkfwreKk3dcki13frWWJm2lG+ZK1TwxtLKsaAZUsaDgQkKt+m21eHl0hCR+
Z5eyHVkTdG1v5YAhfeYmP2QuIWhWlvvKOVlQuCeVvzTxk6Hslf8/GPsdL2SL
70LNoGBErhqSvcL/DlYcINygH3XmFjPXjbcpyMXAotoh7hwfYH+WVxT9TyDy
he/bNsTWmVPe/7iD/r+pH4lNmMil6r1Z2hP2nWzqu/qLii2JarLn2s0dW+Sd
Zksepy8ayL73pocX/AENtT7AOGYMP7TDTOsD4mPOHvcst4yjFvjS7WzLC/vF
qawQ1/lM8mvuraMTCc916NgvCho6GJ8DywTypcKDDpfLUIPtXFrpP/kxQexl
iOj2scQqxBc/IHjlrcwibpMN7jM1YvuvF6Pmoh7tkggscTw7Rqd0IesAcgP3
L6PRBXzkxa46MvKgDTYX/a1VXczQ73Rlb/b3pr55grOd4lvI/oWD2aVm5uGZ
Oj7VKP4Bq0R9IvtND6vPJQHkY4lT46WvCTcCnJpKhZGSO3i4nm5OQLzzQJ2i
InDMlCCmesTi/t8iF131i2DmCmZinRssGDJD9x6O0O8nFiiLWtmgCkgEHn5M
OU5RXuqGoI+6hPIfD2JXi7QI/C1+oZtQEukz+vuTMyPJv/jrrixAG3laA/00
wjSLFQiGbB4zNJsJ+ONZaLhaMmko5GMnYbxImbpRGy5VCouVoi6K/AB5zdwD
V4gqmub4PqbDF4Re+T+IWOZmYcsuqp3dRDb4sCjC9eiL7MNg30c9w4KyilVQ
gBRV5XQ7O1P6sskuV0zgpVjsic/GtmnZY2XVMnW6vZBJ0VaG6Kao3Ak/fHI4
hFDnuV5LQCvdAIZ5MY4h0AdOq3kKodTtfygbcJNirdsp9l0yJOC6RS2koj+L
wLmmcEe2YrDez3Lw/fEGeoBdNnM8IRzxR4ANMRoHEEDsuWxwKsqOrCetEh6d
D1ErkJoawT4NDCByCkZglLtYGQAnOV1GQz9HVw522zJ+S8zrmiYuhEk9A/Pm
YZg1IZ6q/JjrsAyhM2ydvU7mKPC7cRiuHH59YnQK72vSUncqNfg29Qr1GOsV
BCVJuhk7ea16Ag9BzKl3yvP1sy901d5ArU2BimN5dP2/EcUfIIkUKBskx6M/
x6nF7T1hGrBBZRCR04xtEorfBozsywxti/l+1gh7QQPXRduVDEZn9V6S0rMQ
70ORMBUR/8tz2PrnB4fMp2u3OeP8h6MsB2903/u3IQohKNNKHshUhGBDIDm8
THjW3ATQ5H4DT4c0QhARTA31uvnMAvHtmHkczweu3Oi0OqnEflXDs8xk0qE5
jd4+WQKX63ivtTORDg3Vcmu08sq3ZkIx2yPTGQm6eqYDuzWJL/2JP15Vq3tj
2MD+7KNAbmuEfvKnkJ5LABsu3pwYiE9da+90QhcyQWeUslOaLXe5H3mRcDrl
l5ZUm5Ctq7BfcyNS3LPEPqdcPIEhDjsNgTt6OvWgOh/JZl3bsA6sYSxUl4ja
7SdIjpB0nm9aX5KQCTs9e+R/UwuVNoYHkqt9mFkcMEEkHY/SXAm6K+B0/s7z
NMr+NBqfb2q0ZQfBbH+2bOmDr74wfAo2Ydvtu0HgTSX1NPj2orT6QE/j11TN
uPKDgFCcvXMLby5EUAY0M5bFW908AIGYWUI4xRj0uwldUZlT96VDPYDb+V/+
NKADpmehplDdFpNZ7XqNoLRbUqJuEenS6CHCuKR8BOQZ2g9pzJ2ZzyzuONcO
HuWBoDjIBXNN8cnQv4rg47L8hyQDHz/Kqs+h7eXVUglHjbSdh6BhiIwQ+5XO
/RS1fRPDibwODHEEkPmTD1zVo3rJsd+fk2BPZh/norkBe1bYloYekTNZJU3j
/cmxkoOMUta0IFu4tMf8hgA5Gn8EYQWJDhL9wdkEk0Z1sm/YExpSNQ2DBN5p
30O93CYY+oGZgCUpfSeXQzXDEkCgtKNobC/lcSd1hvlcVqV48NuWj77QeOaI
CzlG53SwwSPgEaZ9B/UyfqTt2v1bFpCmfqr7fMiKsh9jkf0JW++AhvGGnAum
SKVMAx/WbxfQwe3PFtk4AOuYW6byqNRe1XTHf3avGZ/B68jJuzPgYBCmoY4v
Q797W3A76R679WixvqxDu/K1s4bxQiOGBZ+uDUenshvWgO1Fozz/+q21Tgxr
2XTltMw3yykDLOacPwjbxIUQ4+ixSllr3haquA4rtRWEhQTtWKDJpVXdkDg2
Y4TbA8wLs+AS2HJRtYxvyf+of2qaluOlqjIZ43DgDlUeA9lt3N7S6xIlmq23
FkNyC+0X1fD0nS45GWTk1KFxWgPrIW/cCEifzXL+zPRjnugednS4Q/hFysOh
N9jx5LkzlPDs3J7BvYu7BK5T/nXgaIoSDmd4FPd0zZZ5zwfCOifOfguunnzW
rolWCTVm2WdYArr1GA0NtMisIYy3G1PFuLCseerfM5HiwLpWAkbRzc5fusB7
H57qCv1/0Dmch1PAdsLj5FlhicEqnKiWLRtMQ/V1e0cZ3NWIubMItx3YfOZ2
EMDS2XFiEDCQaD9PYtEdoECo4ZBrrRCjuTWWEqK1J4uoGSP5008i6YNbDyrK
S8J6h1mQXCjRF1p9Trd4pPcmBUIwLVI/1iesAiDiFhtd/86QLl0sqGvK7Bs/
xHL0qf/2rDMk86Q+mnc5eeuGstEzNXU9bxssQIGd0DIi+6zV31gjqM7/jZco
sfC8BTyq5mzrMYu5V3YJy5T+oRXb4Gk2zxDdddWCWmm99HoD9PSEZnm1FCWm
w83mGgC0YahobTTiKCQq775sSTKC5j/2PO/nybS7nEjDuZC90RA0+fB9pqae
WEaD1CbUwOglH63YBAlttyXVTsgyN0xi/M1ETk4pNFDi1wo7/axUKOBl3tft
meRxR6q8CD3bj1+Z5SynRApxi/tN7wIk1mRJVVg6X0CStiRP0sMEaPqUqWeO
2YwWtbXIUYSQv0Fl1GjBIZnD6uYsmBlsdx85rHr8YYWf6ryEeli0w6ZgRIar
IT98GWK9V2e1/9JqQXK+s8sO+oZXrIRsETn11qdWOlx6Wao3E1Lemagfa6nQ
x9SIf9AjkY06DISKCPyMIX3PdhgQsWxVWSv2ihyPXPZEjRyk5VHjBSi8wL67
sa/5HY9PBeWmISZlDiqon5JtQ/fu7zRd0hnlLAteoM00kr7cAMuUXIcq7jD2
Z3/bK9/21/DQ3uP7hLoNEg6DSbplr2L2kPLYqdbJjJGwZsipSPE0ipyNxjHa
gUwszBV7COUSyEKh8ToSL4qKxR2KD6zlIT/FstkZCs1IKd7Eku0awyN9oZNM
sy/cBC5roMypS2GwRKWr3+7nCk5mtvLL0CHfNYXDTlf5OSHaSIYDz7ncCe2a
XsX2niXzb1WgHE6t0X8ui59P7P1502avZQr17WFAVOjRDyA9J4UpjXqvoTVZ
2hy9yOjrMYi22eLs21s0ndbmFOmTC0UPlc+3IeOqo/OJvxFGPQdQaiQMrIX1
CRCOVGRWVgjvGZsxrZZxGFhKqbi5bcjnRz97oiaWYdU1acVjOt+fAPuYk6iV
t9yxUopiazm2zLWA5AUk/d825XnmNd4Uq4XmIfC8SPuAzE6+GfIGzsA4lU6w
er+buyi5ub6i7mw51/K5xLXhqe3MZgy2Oi7HY8tFp/YcE4d+cf3bsa5FXrov
Y1VcCuVT5QOZpzZsgO7/U43oCubbZfCYPlXRBhGf7xbuoN08WEgo1BnAYRYt
060Ju3RAbti/2+q9tUWshyp7PY0MEtpOtLwJsQ3L+qzjrs9fEsIQq0d/OIZc
ZlORKZe0w7FyzeDcuq2qk60oB+VYME3GEnIPSnadBbfeYKY9qmhnzs6TYVkM
/7O7igGqwaMmkXtFM1M2Cbx/qXoCLWp5qoBIIp2juSXsk+K9T68Jeaed72Bb
ISswY7CJyGkN6xzREjwhdScR+DcmNZDNlkp9TM2m/SuK6DBLolMwIaBQM7rQ
BVdmdNmWrbMYdMcZABwWQUUBrdPwfmt8hS15piI81tQGn4XHyaUpuNgfR2tK
dO67tavRjWLk7gyt83GcbjcrG84rGYiYUPsajAzlSLVpun+SnbmRtkjODeU1
yMCKJ2MjqxzKOMrV2d9crGoAyQIeSZbJLySc5t/tM4afFw46bpjOU5l3Qd0F
FjumKaHrltBox1LC2R4dgCoGGcUyVwNbfRQgmcv69HTPgQnPHYP03GMa4b3j
0Lg+SXvqmFIKlVqTUGnX4KXzGeDz0dwIJCAb6MqcNWXWLgQXZmn+3Z55yNT4
kp0ZHPA3LAzXxY++Ws1acErXnbesf4uKlqgAjCP88pNoEoKFnJYVPOtaM8w1
YBHopf8u8sJcEMCRPxSnOLH3gR795B0zeuY079PIa+VNtrlU5KdEKuiYuCkb
sZ+3OBprKTTogpJsiTk4Xb4uc4YGiFVxTO9x3Uv9Ekw1QV9sddQcjny6gqqc
jyTdJkRrjucei3yoOiB2abvNytXuNfdL9daHMIe+ONqxEMailLz1iHmYO7Sn
IsQ2pL5crH/9Z6SNAKcwtqewHJYhqrtBIcJ9GxXTf81SYb3k2Pvbm3xa6XUD
WhZcQDQrSCk7wEVFyTsu5ntwMfQO24zpYVsjuQvvOA1MpxFD2q0QXy8j24UR
RmZUeGn78Vt65GHzLx2y9xWIizhmyDx6DqLHI7zLaroimeIaEKzDwmLxYYDd
/HFgHTW8yPLj2MVY0pHPIlhJJQ6P0GF18tko2pSVEHYIliHl6RjgtGknPCi/
VVQD8WmH8T5VkWykErYgokhTyna2a3Yxu4dQ84OWf4BRKRFp0YDkgssc5pZ6
U5KWpQMxDaZE+zuh+raOiagB8fnvzH6yK/Plp4h+OrsUMNCccm3AgK5KDZSl
ZaiDBwRTbQFg1y8M3UmyMuFeeQQ4/QStH8Wss5/pNmuw3q82quQnqGM5Iag7
NrnvTHp6d3gBPnP5LGgrKzK2AcYoNPqH2/daA0FZsvEqUp3eiy/dSKp1f5w7
3V/oVNlW+I5+8VhZb6Ed/t9TPhfVurZrMTXPJetBcocMdZPcDenfs5HkId6/
anZFqU3lTrd24vny2bfjI8aveuNtQnW0e86kM1ZXNl+TFRi3Xz25nfDrTJXv
1aHs2Jw4U51jNbanFsKcKvceMs0TGYnQd0D67EED7mc9j3DoeFbltj8Ac3Rh
BtA8wt9LVzprGYtl2jzSKgwY/yBaklXKijmL3WdqmpdUhmfLU+HsGWPmxKvv
LAtx/6Wl119c/CsvSFklWZlicTVxA0NcoJNwBaR4uU+UTl+bJZlZGbBqZpI1
WXD4b64QDqjOGTlE/O2JgH8RpLDXCEm5F0qXVDMk2wbJQ0kU26XOxeM5Jcxa
purM8ps7utfMNp6QCIYyvZjkMwcAA4/QyXdUsjfBeSGh//GMo5oCj5ufd/KI
zvFSlmyJ8fME5VREwQN9301yPlAPUOZuNK2DuKc73cahKy+7MNtXsOG98PFO
/BFQUMb0rXQN3YIe1aYulhhfCwsyBaM2nIR8GnwNueP1WTEIHYNB4ZLmRZbL
7pZY8rJlltQeMT7sVwO29U6zjLsK8OGsjaxUBDAz+S4wH7wxqd7YRf6PAu6S
//LQ1Olo3duhKBuHyzTBGbtZme5Ur+QIhsx61ZKGUkCLlg6FYJ4c45riebrr
OVu37FnBw8yN1uQOIvw/zFXEtS0R7kO3FNl4WrJjV4My96Y7K+kwu+Teblb2
rRWSW23WR6w6v9GGh8aKtQKjv5j+aGM9cIEqqfLT/zdt9hhiVu1qcOjiU/FI
2+mxhFiBKIks7SYmZ0LxOwc/O+SrL0eXYJWOsyusD68QkWov91vv0yi9Kdxu
Hf2t7Hmp0ooIM4goYPD+at+Mt3ZnaZjW8aPCUKC1qO2TwmerORQy4iJtL5ra
HR5KFmIUmoTQ3EZLFueKWM7tDPlinJ4pa4gwhQbmgZgESLv2yDOhhXn8ja+o
UJWL4YopOMLWovAMOIy3G3pSFUD1QzXm56uDzgwTV4AORT5siJRTWZEqhIEf
VbNWpT7QWTO6dPw5uANhH70vFRPT+noon2dKdyeKqkOn7frhJPdBHN8vWoGP
FveZzMzkvWEDRDibx1Ofxn7vUmzz7GDEoWFQhMjcud0ycbJ5dP2yfr0ao3xT
2po0twiXXsOVSI7kygjejro9+YQxXl0T+4cJ5Wl+dR33EE4yCB1gvKvwiwpr
l5Mq6womshZ27RlL4pGJF5gVDHzomScCWoRteSaWDe8MgtXIJWeC9FS2IDE1
UwsD4OSjuy9XJaZ/zsH3Yc5mKF8Bh3YZ4GOF9ElCpSk9PHXXLRTN0klyqGW+
sHfmZq5z6DtPj+jO3MZ6CkYRf9hUXOMHoguS98eUwjIHa18Wy1rplPrKOzYb
fj5IYD4b9prVgB2afdrHAvdH8Qf8bFSV9o8/y77AAviCgDqUnEbbV4GQiO95
MdooNX5pS6+UgYqWX/be6Dv5PNrr91b5B332LmKvaZzBrydY+4h3/MsMgKaW
wT5d1nb4sWdmHDgyNXZ90BTDhOg9UxqGLxC0rqM/sw8ZhTYsX/h7zzbAt2MN
0OJbpFTJVXIJLrttLYtBzNG1wnX3AUN4wOZewXjVkkT7ceniTAP8wTBC1mJR
PxAKLhJWbA36k50CkehhZgOofR9UQLz143TV7gAx+e2VPwXl+LefD57Pv1Nq
rcEiQEg9micFiGlVR5S1Q1yFPSOzRQMLuLzUQhDkbS7EcEpodZtOTqthUtEB
ms/J0qvKEOyDS0io22e1sL2/pmKl+5UwXLLhyIlvBP+w44JRo14VCAVWAEwp
FblFNS6S+CKKhAVnumDE2nuuqR+3CdDEWjHDIh/KWNoHKY2DVBpKJAk6eqrY
5QG0tu9aPNbHa4OKbwGgLymm89027K5EIzfZD5jb/pHx7GgOTNJf/H2xtk0Y
4i9MxZNTOFg45PpeVr6D1/Rv5Er3maoUA2rZboNrsm4UyUQemhpHl+cNxMJA
n72NZenigEWUhsKf1m8fSNtIEHaLvPVwL9VIDzzJ780CJUAdzs2LKE2XL4QO
VccKbbBYF1J7vw3mBq6IB5RIUH1wv2hOS9D6lziwUCRfbqOc+rgzq0CAEJsY
7Y2oeHEgiVKwn7sY0zLSSD1s7wqxfEsQH5ho/gJ/vjYGjTWpv0SED4CngPnM
OGuzManhdQN4u5d6LcxrO7o1ygIxetZ7h39tJDNnYVpGCkBV8x8X7EoIRw52
/seKhG0bvnzpXv8zW88JoCKc+8Tjwe4u/PgoyJ0cUgvIJC6koMu9s7LhpQXk
lEQioAdyFXjk0/LRT6jvscHKpzECOTMO59GH3Hmdku9wfDZsexiodLflMs6j
HClcp1jB1Qe4PdDYwd8K1O7b3m50YQ3gLvquTnIDv4g8osSew+nC9s4B9fIu
OdJou8lXUQ8SVy4mePfI2GzjsATGamxZGd8Sg548i0IST1W6Wv0iCon4XFeh
9eTX7b/iJTi/TZdFvXXzxn8Y6l3jOcBfqsES2v1/MEdrj9Cuq2ZLavFdAS7b
CQT2C4i4vPXQbCFiKPp8MaOvMglgKtdMfu3XSEl6Wffy88gZWMPC3q7p5Vvn
NJXVNfk+Az5A8tmCh/TrEM40HYxZI+kkJfMfN5vlRZJ/VOUwqCGSUtkCz/o+
JgDAgpou/Nl68sEJkCEDKeSYvyY5zHsB0pCG0DE0QcUu975aO1eTiTNhYH+p
T9L2qs9p5QtkpBdM7lHVDhb+oO48UBxDMSkDDyvMGs7HABiInpJDPX6Ctpc8
Tl6u7/oOHc4wOcjfnU1JdiDr033aFRXxuj3pXtvyo0Di3H6kj+ZPb5jsVq7+
iqdVVz9p/8oPwMuUFzN4Zp19gsPeH6v91grNt5ZLSVLrTbZJc6fLBUNNijnZ
QxpCd3vhDu8cYorNvf/cPKIuxsTXOsLshuGi5gpiCGN54W06kkvTr9ZmHfes
dULBeDXyzneKpU/PvKbPOChdjoRo/EOXuJ0Pifoz5M8wcReGEycLQifEBCNo
yJ9sxtcoEs55ccRFlIUmOtOyxegkIU6pNnHkeg//mYUUZcOPToIP/xPiyVKa
/w9WSaIMw5oTyXVppmre76iAIwS65NHxQeu59QzRBVKUr82RoAPBksMMUU2e
P754833vwxvnR3E/Oj01/usnKcBfmWGGxtuVMNH9RU7LRbMziHEjL6wfjr/n
lMWHEdKAXS58zhjI/MBD2a+rzAD8tImen8CB0cXRRaCo4U8S/hEp3zNJ1W1S
+4h33bo/RDIMnkjyoUgzawMBfPiz4YziQ0rV6HWQacHTSgZsE1x4XagZZWV0
KGE4ykLI0SJAGdSABBSpl99xYnLH89yGQdwX9aA8zaPHhO7HsrI2ew9VcAcB
wPLQSgrxus7E4FMN+T0KJDnjDd9XVqYAyCduu4C0kWd8l5BxoNA4EoE68F+9
0WwxidCL/8EgGjxZm7xVYE7Dl+3K90Qavtrg8hSklrDLWubeyNz7oqcQ0zPP
JzFUTkKL7TVIAXLBWCIuFBrJkWREx+CmZfBZhSvbmw1p5UJjLJq1CXl9NKEN
/QM/PFXP3v4d/GenznmlSYQivvLjNMy6m4zeTdqQ5tQoFm9GqBTfgQ0b/LVB
Yk2BgBCqCgaobsoY7rf/csTn5giXVWEkb7e1s7wql0gHMWMFI1qjiAudQxZj
ZyAdXgTyp/yf/Hu0ceMeIwWxJEvUPn97HZsS4b0q4SuUCIcR9pcunZV3TdP6
uHNRqXozp6caaTdQZl5Q328EJP3qfgy9IZjt4gb9ptYdMSTFkRIx5RKGo2Q3
Tp/DgxGrkyoL82iiB5TPEZXJPm3L9ywmuhzst2TeGuSgrUh/TBHv/VD+86yt
wBdNgdPiGJARF5lBkIskwgPNP/c3m7WRWUGTsoewYrHK+9jlaXcj9SfB6R2+
JpYn7NyjMH8JY6x6dC8vrc/CYMIlyqG6MrC6+j774qRg5T5bgg3ZZWyIYveN
19FFY2E+2JowWRQKC2atQ2jgR/t9uN+USgVf7kuaI0Vg161lnRIt/F5ip4Qw
IS89pUPPUU1kMa1xMpohOtbh6Sg58soaumpHOSgbJLgLj1EP+grOq6kBw/W7
ist4SXNeGHdR1meZYcEnot5WClrYJOSIAguhxhUJp4wMCxHvP+8yVi2CfuKi
KLnDnv3DXLLR5wxn6mh7+sz6HLf1jit0SNygFfpmm5rcfHFQDW/9d6aKnc8h
jBt7lecQC4EGN5pHEfzesITtkj3+kvdtuI6vtq7KAPAhhItAe4X9HHVRtzJY
Y8dFuQkWvh0Prx+y98JMat6nCI8VYwvYa4/BFQ57gDFI2/pjIujUuxJqZp9K
3VJhYz2r1BXrK7WEJcf7Nt0lsDhCj8QAAQUtvW1Dir/fS8qi+9PC6XZsck3t
LbGSMWnhIH0b4tmrY/l1pY26lF010xWMAfOlU9AwIfG2yk5j00t/dyTvMwrQ
nTfcYhOQRAnRgCRbcydKbcXml71bvWkj05PO+igY4sBEw9YtEo6NTkHs/3eI
aWjUiLOYjKinWxiZIxSHeL598NbIzfKe8cXfF9rX/LsQpDPb9QypfEe/Jdii
2smB63pQ9s10tJwGvOvUYGuop7e5Jj4B/c7lW0I9juGjdN8LuNmgrcMuh5um
CvM5gcettN+Dcf+u+Fzpdy7DmHDC/4npoVZrrMlsJsqcttoRd52PBlvhHwPr
MH8yt1DF28U3953jmyiKq3TIpj9LdHN14MmZ3dclXNsv544QqMRbMFG4TjCK
fHSEAT6lp6J4R0doqvhJNskXyK9Hx+FFKMtQIycv/8DtdGHEuhMu7+U0SaiR
oDpTa3MN9naf8qg+X9BHxKJPLkLusyNRR1EYgZZN/PId/PoPZta/5zTlEbSV
VkH4z+ESwSPvZrnHcNcoa865CquimaDn3wvy1nhlBCe9fU6iiVbvzebym2Ov
YPPHCk7MwoYlGlLUI0Il8szxiLlpAmnMT8f3GJD7QR61xElDGe7GvahUdXjk
k9MCJfeIp4WCnb3nm5gaMqFk9yXXsIkg6G928xc3D83532CvCBFXaLWifJ4Q
YLQpw124YrmYTkzd8SjIJNBbMzGbtSmXPIRWH6evmR9oXg37OjgQ3Ythhqm5
rBFIucGY1yojMWzsLiXgWZ2xd+Ae+r4CwgKcoknvP05NUANS/pS11uyp7JTy
0aq/Uab3pnWIGTEYJOCAAZ/NqLLxMWV/BWx+Rjb6EfTWDfSWuxLn3jhDj7Fz
HYlZ7nGifM8IuDTPtv+UGQ9kKHr5XOSc6AhEFi+htxAdRNqDFDHtHwjMyY6t
e6KChZq5ifZjszjja68I1Kjn7dKl4sHTfL/SaMqR0sPpMUCS0XHtgLgjXzPQ
kPOgVeRaofrrS06N2TX7HAajwtW+foYTswdjMiTXrjg6cHWgOhvz1xBlSfKO
LYWsKNGIX3SCeEsd6Cbp5fOOePOV5lXq4biwsRlIExrqOty+LtmLvr6KlR1x
grZvKZMmThYJMH+Nj8t8pA0hLQH8ZmsZOz1BlTfsE6sgGqdstqTxY8YdHrua
DBuP8/7vcMu6wtN6nKOfqqw8BhMhrOJjf3KpBDF5mx4QdhbfjvBJ2yf/t0JH
NjTFAE7f2aKNSN9mGW3wbyQTtoz+1Eu3BgAU6EOM9amTf0vO53ZKTUon0mm8
x9RNflyZrovs8abZEwVBUaCcAEGwtfvjrk1Ty9SK1MKAKauWcKyqKshxmfyK
FRL5CqZTOjajLBE9Zn3wqowEUH73FFOOKLRi/yGNJN8K30eNORuwYh5xUB0p
4/GkkNHceIfStPfQND0EZsW2njveRqDbab/wChN2NdKQzXMv1/XizXlOCL9r
El0rbbTmw+cZL2rFdejQSQlWhsapJaW2cDKbq53wIG1XjK+owZcA/nPITUy5
EtItgVkJpPg2euwRb0UZE1Ig+RkDSnVlyiKNqDni9GlHqjcE506k+5rYardy
soJjJtakdwUjbN110nuwYM9h9KJFye+7rPR7hEiMwlu6zqolKFM8X3brP5af
ZSev9nth08sWdJ256K9Ml6yyB3d5IRB1h3EgAstOQNxOZ7HK8kHNFCm3sN7P
Zv3PgtbmJVPGEVSG9uvAHdVfLVCgp/7MBUjEYAJMtiEEqdfccyq29nTCL58J
M4wvoJBCVU6asDZURujZqpsNcm5VyWnd00PdHzcHZVKWHJkWnn9MiKYznfxC
AGByr8lf8FYGx7sGmXZN9gOndwKvXsx6W/wrviUIYNRwT4FO/TKksvkTsB62
VsdQZEOFZMSz+4pomS+5KJoM5kDpIc/fiunWzBqO8bWcDyqCIfCr9dX2alCO
3kMtWKNccQLDxytBqVANTwKTjGS1NgJQt1THAdar2dv1RsfoGPtQjpFxUbxX
izVhvoJooPCEF0FesHUfIpWnw0XkJ7iJFpP6R7EJE2ENxhQholRP0pd6RweM
vku3N6jOpMWQ5REr1H95ETaJJQdM50MFhl7ULBGohpwD0RP+IMa6kYq+qJNa
uXxlW0UZg1FQ/dKno9Yak1B1yZzxOQ6uzLN+x2N+0C4npjW+nxkaZKY29IxG
ZEA1pLFRbxIh0iModuByb20/gjGbDX9Y8f0P006wv/ey9sfV2pJdhFh2AiiS
01DA3cOADyILFPSQhoEcZmqap63RFENnWNzW8s3xPpCNi9QuwyfOgScwT5C4
QBCEJtz/GcWn0YAWLo3Cl3DHzhbiPquz59rGFX2hpx9i+xv1xot7+x2cruab
1dmg4di5RtgljhaVeEGsM+9oQRnEUMSOudklMWRnoRgg/47qOxiCYDeT5J2g
Vpw8xLKcLUcU1CMe5E67fDMjpsZJQ9/D/hx1LRpLi+OWPR/zCH5lfLYxtqpS
qZlxFvkpA1px1xmo9EEIBMFg5/zrwX5SsIgdpDcWUs5s0kVgAIGXrx5ioKQl
tCWjGbpP4aS7U/BKloRaOxvoAQ3SVIzgLKdSdNwyxib7l+GTbDXeoW3SYznn
HtgXEAKc5T7xlyjNWgy+TmTRoAdbzwIrU6IGXJpvlMSHCiqQO/aBucx8EAWY
3V1PWTxgqeoJ5VBav5og35oUD3Er55h5XlbraEW2soaflwGKUiS/Llyq1SJL
BWFajU6Y94tK1TRocMLEWn7dwkrhL6GRKg7zPigwQWwyHuIpxONnwPOWjHuk
zhgzRe4c5U7BGwxbQG5X4MveQRrPua4kJ2CMJ/MqtG5BPkXkVyOvRhiEm1vw
EOSOEg77xl4zzXJw9gsT+p71CujrhI9WElJ2sAM3/zTWpoqoPqWbe0JI8rn6
K4CtOSxSBjWFKUJXiBqryO3czh+WOKb24Ib+zobHKcGGzYtuZHBKXM2Rjlua
D35lQDa/16Z1TgmNblLFIEBYcaHSq5C+tiEYGc0Qe5Wjv0OHZqmgVTLj0v8g
v67nGK7HGIDsRzObAtE3O4ZbxdgMlQqjTc5/ggopXJTpIEGG9oOGSoQGkMB2
ISY2fD9LcqRYtYs8YtRJsFiDFX45TACuuqyc/i9zlAZZL958Y4fGw4FGQgdb
4BUKkdK2XYdXtdVzPD0hpfB0yU5nml18JRlJZNiN8k4IBWE5Cz5YWJgz+q7A
4RhWcITPdLFePaNWyfCKhRb7ZhPltjO4PtFejrBjMqdzc7DZIvrf/qRAdwLo
Px/IckN+7wTLoILucnBvAZqRrIIX2oV9LNPZxKh/x/9K27z9dG1J/1WxBGSp
+4VTHwcYO8c3Uoo3gu4LeaF7E3Fsg6t9qDP4n/0GpfC5D4hhMNgSp9BCADVX
VdWRBN53JyeEJw0YkEmiGDDR70IL2NaHZrF72o1YuND4ou5cxSKoxiCw/O+M
hy8aqLAJRI6ytQI8YXTWw+hpp1pioxleAcwH1e+WeyOBb94RgybbYRdGnDa1
rCorWv6d1FaWOWkI29AHucQa5Rnin0azUnx1SAP7zUhTubsSFv4196tAlx4o
/P5q9XvDHax3i018Z/o65EE30bwe/THOtKZvvnDyh7qLXoPSIE2HwgkJ6Mr3
T3VAXtAfoyjYSfRdKocacsujfH2LUwJfB0hND8pWSEJJhoXJM0xuMyWBj2XR
K+1adl+TTH5eKAX5OdgE3lrfy8xQGorrDfPpJXIPfwpbD3AuNPJxh/cX7qaW
lDh351wyr5YsvK+MZWBJZRrZT+8QPVvyFk5+1ywXPtRiPGrsJiMp+B+Vsz5N
qkgz1a3/KaaTQDQ8eV6+LKWm2zBlPpsbqoRWQlnlKLK064pi1O1I7RTBtNBI
Nt2/hYxHQRxQ6I7PoKu5awQKxij1FAM1UvFNOehsKpBXUd14nLrK0tBn/wRZ
nAMtA1TLTuA/G5RBebXLARpZHw/M1W5r74ZghMkO+//cdW5RbBpqNJElSLhC
T3vGH7SkrZESL28v8GxVAi96oQlxqtsmkVw/LAvGIno+fpeMtT++TLpUPFqz
bWseW3uevnohCqp9Ye8oVokPrcb+tZK2YBXbgfK/z1f3loxEkPvibvlgysXb
4duSKgVxi60SzKOT3qNG0KQlEJDtX0vOQtRLeIH8aWcOJU4rYXG3duqd/9KW
hiET200kpxuZsWt5l9VV93o2FRxtuIn3JKqAMagOAsOFV/3p8DUpeDaLNCI0
S4sDBDKvlEi901CC8QUyTeg5RJYfnd9BQM9LU07unXVwFUaJrdK65wnZdAIQ
HnFKQK3DQm28XyYJTt8yPcH9dog1agWpf+Y6HcBe2H1XyVub32AL+Q4veLle
0cQyQPjtjfW75rReI1uUmMFrtcyJTGQzcbWOGBFB8qmR4caU9cNv8AZWFrnj
77VQKlhl0AYeBSmkdWXM1yMKDfI02u/102llGQsDFCtfDVEEGVeLPXuir5o7
AauNcdJwsIGbrt4Q7zRCJyrpeVm4rGJaBfCTWNTgkpvHMsZ5HkVKZBaR4LqI
XxjqP18Ub62zsQlGH6yYGmV1/LQy9+ENPSKSfS6RXYaD3e16wgf2FY5HV6AR
xkJ6yVyXDsXH6GhuZ9PCp2P+Y7gFOkmSJ4XYv4s1vGqlNAMuH6w6RhCiGxHJ
jpqFvxKgODF+ovTIszqPZkDlYryJVaU1FD6oKFsCtMW4DG4iRoCot9JzfMTA
JHk67TfGw5+wiqgLaDShlnuuJ6UTaudsAsdQpnRUBc3hUaZAXufWwYZO0TLZ
WICUFM1pKTTMlZLUTlhHtu33na3vjgz0K0HLOtLG2jsPm4cjflgxzHQ82YQ0
czHmS5HS/6OPizblCaZPk7yXbNHLDvmgLH5jCU+lLimmgcSb4LLkrLeUPCaQ
8CwsQ2zgLBUZLXUgAPjQztYw4NyYRGyc2SGgqXT8h6VPMCCLQXwcO/t70S2G
tRxLv/p7ltlmdW23Xs18ksBoQSff2ZhME24x/PPNdIEu7A1wsDmCoDZADzQ0
SRed8n3iovHDnQKvNIMS5sjFyu1Ed8BnXZeLqS2fSwrE0AXCSOQcc1G2qYjG
gM5QbfKnU/nANso31iEsYhUt26jN21HQFP0VQ1ILtzsIPR85BAno0t0pcnxP
VAVgErHCgtvBH+yUz6v7nwgmtofsLhdL4WNuQvQVZtdSQjhyDXfuMyOctLPZ
3FShDJGebagOiDUKUkUwBmWBrbUzV9h/pGbJZ9u/KzYfIYTfUtr67DcMHlkm
tCLNKslNYXFc742vodD1MRPwrjtLFSdyag5GH2hOaIi8B20hKYcr5FvagNAq
yKK7fOCLFiN4KPfpd8F0c+AvjZh6Whue+vn907dtGJowIlJtFL25WjGhuyOs
GH5yMHZDUGxNbvHYnqAQjyExF/ks67Xk90cR5e1CUM+eZYesgSYmPFPfgcy1
jZtQo4Of9LOv4HT+40/0OmAgb4IZ2thgqVXrPzPtZE9FpPEuhu9E9qm/jVwR
5rSwEYjuey/5ye1qhKWAFNFq66n0Vq55nXlETmdBuoU50vn0zXnfjXXCcHeo
kGEO8EHQ/ehocK+YkLkxcjlej6hyLzQsKyPrOdf+yq+nZUJ5u+aFbiPRTx+S
gS5Wpk6jw9bM4ta5IhU6FmS2PpVY//uNdDaix/hwu0t3Zd42H9llL0pc4u+m
4n7BJ9JeuAOIb545Mr9J4Jw0CXzkv2ZzgGrzZfmF8LBnYPup8J41pL3jflQQ
WhMX2vpGZTkQffULRNQHf/dKHVLK9OpOy8xPhknFV14t9yCiiQ5zxQhv0RPt
Vw9OTswCiFC9HFLTL3nyXbUer7oIV/mJSLGns5OqomgczAh8WVbbVeumv2Wi
ZyMXa+ZCyz0OlGVxxAaJmOsFW1QOYGBNAUf1200Xdfm/Kv+XYbgat7SD+p35
I2YJsAV7INFhvKy4Vbt7Rm//o6YyCU7Fz1cVwAV8hynsF4n5vRAGlKNTikwu
8R5ClMShjxnbqEA+1yClRYgbmRftw2doqx9B3yoUGgqkH8/bGLKV5a/Fg6wQ
LrRK91LRbbzQnBtxRkrK9wylarHMs+YFuwoPPqTXkMj5dqvoXfShsT+Hd6kK
K60UK5+qTOOD4NTDLbPzdtMwnQ74/2slakK4b4Ui90PMQNY6amrBiw9s02NA
51FxEZb/DXAb+MUpmyOepDr63DX2gyEe+D0DA5Zo4vgzz0Nqqv4mdnXKgjUM
icdssi9MROan7ALYvWeHN1zMTbcOFJNuy0JXFrOvRFKRwU2PpWqrpv08Jqzk
cYeIqwRsXJv8ICZo9PvrxEkpTJb0h4qwrQHzYJBfYOsg8f0rA/CihJtfDYTP
Rz8cnjKelDHML0v9sEwH0W2ihA3yC4hX0d842c58gz3qjrofQ5RtfrDYyDYj
j9eWEjJsNSDxYEllqUHnmCbB0ovuv4+shH7FplyESAclahrteO7b5MRq5FRW
YtPY/AOMJdq3pU961xKUx27wuxe2hV4NDbZsFQMKt0C3Wo6W5eOSvIomJ62P
B1Www/rCFoiOiRuMIKTHDroQy7M67If+NEcsQJeyuD8Gy7mgwEMC5onK4Lqm
nr3giVCDl6tZZfHsxQBCQdkPoRjhdXC/J2MHoQI2tZRH2hc6jlHMGs/HCHgG
ZUET5f4uLrXGh1UoTSYoyK8WIAK47w9dQ6WxSPre0B1nj2L/8w5RGNQyUfQP
MPqs4a/Wm9lRTh3erF4G3aYQpGRAB3G5V8sdxCAU5qOc6s64mEhfEtLyoaNr
Hvgl7AMXS9xc7nIZxGJAUckQN8EyWFYt3Kmlg9OM/ROwfzRumxFjcwedp9Py
eFNVfrO6TVvV3B+pehC/J3Uq5wK0FphgPdOab0TX3gccW/qE18/VWMVo6jHU
fdRNfJZyTr01BcV/+nTBrxWz6VLBQEJn8XJ5IyhIZpVn0m3++L84TodhlyZc
zjdYyL5jFqPonFRRu9NZjJyT54Dpxu2symwNCt/UukWb1UXcPcSEZLZi6Tzd
RfxHrTp74V5KS3sqV9skqK7lcW8ioN/pFdqfcCJWq6OMyJxTOKcmqpsJhMHr
+ryJOLkYlQRqdbeZWKRW77LETSSVHkcNe5sfPaifNfOLj3PBtVAJrQvDGHFU
R+dFi7Inj4kx2fjKv5MWPXa6gUEg45khKbgGHCra0vtHg+iefVXwAA1bcyRh
aXP3Es7NJ0pcM6IR02ywREJkq0d3qp1AmkFiPy+6oqFz47rNRNFljccP5KYd
jH/q+lfWRiJgzufB5V9jGpMV9d0GMw9hcoY4iV5FGegz5xBtqxsQ4+RmkE5R
PJgtrmZdWHJZk2+SLxMf3jsMML0Ruu1PgHKixZ+aDZEFlxwYyjWf1VWiT0LR
YjrKnwXZ//86IVqDrp4yPLkSPeMsGgS2I3ZChRyNLS3q5F7ad/2L5aAqmr33
sI9tfefLDkKTwDhswth4DW4/TKVW2zFJQe3aQ+KNeVHJSbZAuWs+r8gKgbCq
yyd8dy13y+NhyNMM+mGqT1UC2VsZ/r367J2hoWfqFk7Ug5ffw9++UD7bkzZM
dfQbMk13UoaOS99UA+xzZDScXgn6xSjZVNxQwkC3Ngm23Vftd7tTmxUaBCON
Jei/sGqBov0/+HUzIls1dtfhcLPbEYLSx1THUXe0LiHTq4VZBQlpp0/FCnZv
ubLvwQa6c3kDJif4tC4uUV8a/lkb1ug7RFLMF3rDDpQZbocK9GGI00X+eiiu
nHwEOUWfcAZt5YWek+1xBqsuHD3WDSRZiHcSHiJWmTNPS+UJVfOwLm2P8cfs
VGBTRwao3f3pxe/8ecWUCm/65La2fi+jKBR+oHQpMMDRnobCYBlVGocOTi3e
uom43ocrI/LYcBTBCNT5EpDDi1Jqvn4JekbkJYcD1W5hP5jXxxY2IEU2ob3W
8fhqsxMmznWfSdLN4nAu7vnFUuse6Nq65r3f0aEcDUzV0fIV7I4MdpClU9Cb
dNSdusvEzP7y+GV0i89JC+GcoHnn3lyjh2muUM7z8R6fsjvl4fLsoMGP8w7f
p+JBFxMZiBx/VbOxaB3Ie/+FoBTg0Q1UPouSSzg/MkHQH3Bw/UesZ3MrYkBo
LROToczLiYXtbER9f9enY7Ym9ZnNc9w1zW3+B5MSdsDmeFCaCmLYpHDNHBar
PmeA44DsFyQZvgsEwB4nOS0t48VNTIvFiQhie3lgf30666wF30vhL7Ql6He0
ZSy2QxNddTrydL33oyOXdTcOioNSEZG0O9OkUA5Q9dukXNF4JltcvO79HRZx
nfPXPcSq7QIgcTZsQC46ikNH7x+wVT0SABq60kQacPgqpfkTsBnU0aQRmBDC
YGzJRrrdzMq5Gad7XbH3ZWaGp0zpPc1hJoiEK17GKbhmsRrVexXpj9wxiq3J
dFlfzw4ost1QLmGQAEx9tDCJyBHJCG3E7xZ8W534tkioHQ4LKm1ESUPyQyIS
ZOxw6PZQ9qAxjpLodlg3cpDoen++1/x5nHMpB1VMJDld/nHH38x9bIcrp+xP
ZcrL3UoR/gqWQ63TpYzRpX3NILsziQluQiSJ9IliMPIJ8/mc+tg7EDK+aiT+
0PEDRgVozhV668vAXmy7ypoDEQPseO7YifNGXFRPlEhs3BIJy1JG//3ClCvM
26F7Rhzu340ZzU5v7p4KV0aixV+R3IEQBFabgOJDWpdvWINN+2j9EuIyvepK
SaWxvtEuJ7jZBaoMTZvaouiFED8fZW53OQBqebv0KMqDFHOD5b8ejBxZhja+
lx1Le5IItRm/YUajGSAqP2Z+5iRsGwdvwSkf8gI81n4LoKZUVeYD18LwOuEd
pf3TH7KuKCiKA3RJgwNcd2AwBlmfIwfUI7ZWfbRcnU0AgRu1AYH4505R+n36
cOYWteYagWYEdBQVPJeKFLvhrT95136mRnqA1j91tPG7hmujnHQOpy5YXQ8a
UBjqYLRevTUmcFIHlGtotgiNgUMVwUdxk1rOgpYm0OO+dtEV2hbnPsdDg8BD
7yIOJ9eQNCuFgpAntkCtD0T1Zm1Y+I+d1nOKHjGs70i5Rwot4L1q/ByKMAJg
d3+85/E6xgGzIcpcs+QNSyhsVTOWPthG1634JJ1RgI4oUyhX/oAnrBRumqR2
BjnXlHoS3xPVE12LwvfTYWXnNGhdL1OX3XM+F8cWEnDwGO2WLaVssBkkxYNN
PKEP64OnQpMulkHP/13xDOCFf+u9Eq71GkNLZBkzKVs7UU2K2XrOQSsxFMCi
n0jyJ/dhqI4+3w+z0ZgycgbTzfysW94RiQ0rTdHAewl7Pg7356wrDfzg+/js
U53c+BfeDuRo4+hfc4Xk4FvO/zkY3caEhZ/4FKuL/wbHrflxv8imqP9pPSl5
3qLChSEGv6HhtB3D+8PPiPYkRBxYDMkZYNmwsiG/3euQbb9pMNCwxkbwUOrv
DUbabhh6qCNCVS9FmFRVbBnnHbT61gbMw3fERTYYRxpwY/zcUUD+4kLgsbNN
Lqljvz+0NKztg+mfuWYUYTSeAYY3Wx9N/U4V9IeoAf+Pz4X77Y4zFodLYCws
hSgKRf7EyeWJ5YbGrampvtsC+F8eS/GcCcPZZ7MTD14r9ZPR/C/PF1WrVozz
h3JF1rcnHqJBUMqjUDQL9/FhvvsLDbQLJsAMw5C3Q9K72OHknObVWT4mZtBX
ugRNzQgzWLfoVbgT4++9TOi2RkIxYrBNECv8sKAkC9FOFhtIL3CIcnAE0Ahs
OcpSLLXioMoCmLT+7KQ4F77wiiRygmI/9qukJwqI5ETP2vPL5taTsSMeorpc
awng9F2SVYxcSAFmvzGDahVChBpxRL2OzdWi/byB18Z6Uq1TpRgwB43ShPk1
nqlRMYs2OSaHWVy+Q64FHcIzHz+eFfCTeDxqwEGcRIuCLLecUy8DcZBjdHs1
yY6OcaQ7R4bMtqgeoOkUkfYY1O9oq0FZp9zuVKJ0zkx9JoYAhDz4dvRWTipv
v+OOxhT3VJZiCgXBnTGtRXn1211g1a2/BfEe7yJnhubw3hTThFZSdK9S+DkC
tIc2UokymPaooRowtmNIejMYJa2lquM2eqWGO0JsKGI6RGJDkF+6dWyMq6Pi
nSrhsPFLKa+J/oHYNuPhWw12n/vclXZw7xSVwRy/QWBhVJnkj9xvDxYi7V4x
9l/YnJru2l8nUQtlpSn15CByTNLNeV3AR888U2cx0hZ5EhAN6LvTm2MMD1b1
Pzrow6eN4bvZdu0xUkGFtgjVi3m4YD6cNeTQ0w6QXjmAzrAycfCVnjMN1jEW
VA9blDrmJRMiemmcvmybH9CvePAwFIXkJCy5jxavMrBtK5r6j70GwBAnfg0t
0UTX1CW4T0sy3gcpxI+MndwFAg+iKPv5ph2jBoVCeiNASgelmdDRt7LLGPCn
xlXa7fQwJR2Mi9VQYr7pqQ7sooTrCV4oRetyMAEus1drdeWKNfCaNeNIERnL
WWCWfjXrQhMT9zKR5QG+ym79wsCYBUY6qqAoljJdk2CHM29pNoInQ2HgnGLa
Kyxkr4nMRmhuq+u97g+1pPPSNWdeWm7FTpvWVZA5/WoGITSv8fCIax3/XXrU
bIor/3N4mq4W3be45z/Ca2wKQIK3MkqDsoWPfFXDBBaBTXLixtuGP2hdl16E
oLdJZrccJtI2hxa5fDW/VLlLGNvTpk8Lb8N5IHyOPniwvJy8VhY9q4psU2PO
Tw+BOzT+Pa2DdGeFYc+sXLa8SkCduZX07TDs7Dua8jlWtij1XgMe2MC27g7u
dozx00MAsc6TYn5+FJcsISFzORfG/3WpWOXKfpCT3Zmx7W8aD47BhLjm+n/f
TlHpLjyidvQvohLIZbdoo05sKpcLOvtfqkUUTqZMUYOlw9GNbmriyYsc55f2
C7Y9kJrAnevNLbq4X/pgBIi+FGfnS5fQXggP5WzKDkj9m636Z5m/F/ZQ+9L0
BLkguKO1RfSd0IkEqGzaKrHCr6699pP4OMtbgmu0JdmWELCInT6nfhw7DDfp
VgQK5Jdz05unFN+PnOAG6fPMGGCuWnNRGYQ7ncFsNP4fVNZS8Z/fKRgNcKm7
ADAzE5aTdOrvMahIHcfzETlBuYaz/bP/uIjmXVLXkd7a5cbbxKyu/dAyICjP
FNttX7rdQ/6ubG9kWlls9eMv9jhjz3Iah/9IpYQsZfRw5a1WmzM3JG+r0lyM
AUANynELzvD+Z6MpasPVAyYbIPvhm6ylkTuMFin2DTGtDPAsfqiiJ3zTqI6w
SvIJGijfg0AV9ti2pYr9AdZ5zmmE6i270PIm2fzd4JIUuHkO/ObxE/80GIbo
6qk1FN2cafoONAMTGle5zxf+ABJU0y6iXCPG7wVCl55J8oragee5HNOW59XV
3N45oZ3Rs7jkZTAUrz6gQzMGRrxAT+1aEUq8jrUFe0hI2evGq7AWeMjpxQ7N
zf6+EuzTGkBuLolj/xrxRlXc7aAMdK9hK2M1wtvZ0vFcr4DIapC8mpFPaGd9
PMbGt1rLaVt8WAz0A/cDbSXMTixOni3Q/0eGHH84Ydyoqr1ZFSbK1D5RVVs9
m/jreB8ildR9ogW0pa+Z4UEmRqzA7cGs8Y+BR+BKL4Cle6P/lVQOY8D3K65p
eO0X4OUe4JWQ3aUAa7B9jhV19Oyxg44UdhDrBkuImvc9LR+cfJLebFvjumNl
vaKYHSAEZelmSNdpy8T9UmBh8f1rid3v/y8tD9B6OkMMdZONXYQ8gDeuzE+g
t+EuSyCWtPtmS0auzR/gxCeYua+KPeSdijHtZxVD9QAiKnToWqPfWdX4EzBU
6P3/P3uzzDWV0FqYRf0dUyIHoL4eRWRxt0TqcbqfEQLHjgPGL+Q+XTQZmYEG
UfN3gqH2CDs15gv77JgpvKwC/73HFb1xk6H2ubTMmwaJmlrqxk9UXin5LPmV
erJi1NGcw05+SyYavEIkIbiYR1mKaovfQclBTTJq9TMy6wb5zIe7KAp08mjl
uXB8IDivY9kav3hidRp8B40zA7lRk8PYZZpsJECWyr1ESE7oPMhbKcaD6MSh
sFKMjkvHaKexqmUR/2FaH/8BtupMnPqgS+ImPHKB3xvOkpD/uvzRJSs9NIBE
wp8lkUHbI/K89wD0BPfUzMF8W4By9To9rCgGATHNuQKsvTwiewCPesEcgN52
7uy7caLVeeX5+SAaM4OVT0sbPliIHPY540IHExYU4B/A2fSUVpjrqQdV1Zok
6XHXzJvsbqEEWHjzCAIkj1p/1xP3Yy4CkIimorH/ydIaa+dMABcqIuP0nWnd
Q4/wyzOsv09QsdQ+lSNNWx0/z+YdTwxELdWRr/T0tYHsAHfFvRmesbjmBLkG
3U5uxPenCd+SczKPD2RWZK6dA/ud67fk9Jtl8JLu1s6UNh867DKh6J+D0Y5y
kvmOk467RsJ5GLRqt2qtnD6Mj3JDmgtXYh2zMCE7ItbfPLjTtJIxkEz+NEQF
QB8VWBbSrCXN/7YFJV8f1eP9EXVtENaFB3ALRcomYRF6Ef3NvFT2Ffuv599h
daUQcrWTC5QZ9XhhMe7hxEpnfwNddReEAqARrlXrQFc3G3S7twBEN+UiXpf6
RMo1nSKk/Ng3PkK9BjsXaOFvIrp/5Xxf2Gf784hL5bspkRGOVQuzYLfS3pFF
egu6S91sMNf+H+k0eu7olXrEaqorFNJZwwF9GfcoeyKpw69hdvYjjBR3qHbX
4OrfV91WWCGkEDdIxdzP1FgXGG6B/QBq6KKtveurQ4gUBOqtzhBNLKT54wsf
yLyI0DPNy/WMit8smSTlhcELVQ2WD3/SQmwc1ZFaQzko/skXCAZVHl0i0XnW
O446XEWldQxaN2HSPLgldoGpOrvU91ig/31ctHNv+e21Fqi364hDYIP+qpXc
go38Fo2+FYuX5QSAAR8g0A25DGnhY3oOIPZ8j3cjLJR3YhO5rVfzYnYcQ/Qa
mvfuN/FL7HYmiiLehhTnUkP5xsggOI+xAXT9kZna+g5Sm25b8FEKd9Es3Pyk
NXzhXLQQNQMIwFDc3/jWDTCYKrPQreE5GcM/JgI1e4/j2tJgjkNaVejCmkTo
Dx+4WSX5COHZEx+Cn3WSUYtdGWgRr791XH1+Ok+y+N/Lyi3fJoVTS1G3kUVh
rHP4D8QX2gi0uknTJ1uyAasoJq2qqmZCvwXokCmrnRSF98Br1353NLPEMBQb
Hy6SaFkHPMOpr8h7MNHjP7giCVcLurGpL091IXq9J3TmG/+JdvemXEA1XvYx
dyhKQo+8/mooNse42ap+RSRh+0yYqjHHa3v/8IbytIz4JezolZrJXYebZ8+W
FdCP6tKmMT/Ju5BnhxCR4u98BfP3s29Ev3Oc9FuI+9hiZIkeaQg6RaKMYp1t
emDm6y7YTSfQ4visqkbQZKKGUJjCh4xPlcfmMTXWpotF8NO41MTfz2JBanHO
raC3Cde2CVNbcn9mZlzvr2dvNGRY9M7SnXLCDK2CsLSqSJ9Hr4KIkyjZRjdS
SBxzuPueMUzu6GARW6mR0HehE8MuL+pHrJOOw3LFgUSsLMWeeIu9vsvgvqBi
+9bZmUFVVMF2pdJFcEgBK0G10uKQsR8NGtsDmJDCTgVgywKfY99bu8fNkQIe
dI/bBaiXD12u3YROfjo8pyx/LM8MnoXn7Sx5PJKrWNxUoVeTmFSmvfzE5gm8
SoIZC2xc6+70MnLe6F3kzdC3zsAREFG6hJXLlwFMPBNYG+53+i0fdrEuSMLY
VsiQCQSzPmrfbZLbLDgqd8ecPZwXoNRoH6vdR+PMpOLWFcG7ze/A9+1r89G5
WxTQ05cbCN4wRCy+/5vOmn3M1mc1M8imNShwD4+IWYE42kQxCVJG+XkC+1HY
KDPXeczCqRydpt5pYqGpJrl8ONhPsecjCmDFU3BWi/W7eaE0KI+5GEswDS7R
jV8kTxwH3xJnEZJBQ3NCogjaed76JD6r6NizBeoglUkItfkWwKw77D6P7P+1
Q2DKgUMeyXh7nuwTcHvTV5e3gMA+0Ay64OHrF52TEieg1u38FB0PdT75cxrb
Da5w/FmGGn+PHNck8KFedUREw97xF9y1Bu3vsv0zr0IRKmwzX5ZvQxHmhixO
c6H/QxZksEcfzg5AZU/xkUJl/D7ECV4ttS/jxDpYQx4Ezmjl6JzTWfsgpyoI
7MKPhyd9gd8Rb+g7jHeYt+6norn2LXyUCLUflXwBCwg/gZ1Rvk70jvUV7Q+I
ZxbQr/+eoQt7vif3lbxESOzdlfluD8fW76t7LvuSbtUvcjlP2+gFcq/X1iO5
Fu/AS6u+Q0+0K3qYfpNcd3r4aAxfctAGKgmo2WzyVUVW+v4SHIvQiy7tKHaN
DKqQzFGCjSJbk8Gl3SE/Lrk51gdfxF1ADd3GZWd97ztlfN2TOEDXh1ZQwcNF
oPMVuRkiLFR9hZDXfGCHtvu8OpW0LcNtHrSBZzHJUmO1NBoeYFaQHM55fYCe
jrt8xteoR+FHoR5eB0gziRmgfOYhrfInJrpFvG15zY4K7SS6sFMkIzrkFAN5
WUPy5sNNoynw6ZuAUEOFWMnVGwqTADKsU0tqrUTj/mQaWWLoFmld9rl26pOM
I6mQKaGxk7hlSo1wEWmnvz39n1jyv16ir8LaPaF64hMbd1spUNgXmBC4nCTT
wCODLULpJzWrvEi492geSaQi8IADau9rrdAbD9Ip/8tATZ91RUZ3lwq6YJXH
2xMNzuyU6rOuYyrYUcZdO8p+68Q1asfLnlhCH+HAnc7hkW+XPmrF9UdoG4Aq
J6tDuV3cm/d2tEOf6ZEuG1Xv+0PLWVYnTJqfhtSxL4uveRwyNRKaUXO3yzKx
5e/wTvhasuDbjD0bIdRhXf0XkZdZxsrminSWn5dijBtMVcIBwCqtrUs4pov2
S/i0UXoJry+y232FJf2EUmofB5yqXBkWDfzjGXoXhb91vVmmJlzsPBhIE4VU
CqRXshOFHN/bUCOQ/MYJx9R9SVNk4n0GNDgulqdxu2ELFtONDFnztvi8VXH8
Hm5tFC5iG3TEydPSUVN+5+2ap+iv13oI8JqaJ5wMDV9YP55CLmkZqUgdecpb
2atiNcgSkzd2uT38s+iXbdZOffwdSVCkRmIE5RbLC4BgntWJqqLm2PNN+HIM
xjKPQx1iHo97M+86dQlE1hzkS3Ka3nMiwQCpS0f/wRfTUHTml6/CTnz5XcHK
fymWjyZWqjfHiY/yINf1vtRpUyh+DtwGMrY4t26uJ0SbntRCjYpHheZyNOPB
0BkOTrfgjmJhcVy7pXHeCaushO8jmjDpVqvmeUtTS1TxKpaBtfd5UQR+wfvW
78OQfnqrDrynhlZ9S8Z5EOES5L82D8Ad18WqwheJ04OE7Ojh+C5GUiLkWKUu
FJHDGonKanVNm7qlEamX2TeYNwsJo2z2faDR2vmCvD+1GJdrKfzwCuuP5IMb
qPlq3u3oPQKffD8k6dCRIIgg4RRxasBWhNpqNzE7A1pKbqVRCuf7xJtIeIHg
vrbs89KjvLwAm+4oEfpeE4dIJtXMJ/YUtmDcNhEJI/swLle7Q8fCWkPiYIUq
RwizNZ00/ZrXtp08ykiuH+EVSZUemoeGDjjEGI+urEYGdkkzjmlP4FVPKNOR
meON7Xo3koYngsIa0kw2eSIKBE8McgzYZyw8NSROxHXOPPAiSqyqnlD8crwa
2TQG5ECIS0Yymqz2QCvg/4+0NZB+sYISr1vBezpRls6+IRulE8dDle+YB3mo
d6gQSeNL4Uy90AZ613gbwS0OMpy756KnqGIaG/EunKbMbEuBnMGPcSO6VN3U
eYxq8T5qCMJyW4PspWZGdDGaYG0Nu7+MZyF/RYfZ+hFkg+FP3oylB79QSrFJ
+NWvmiA6gLppuAwgLibCZ5yyJ0Xuk1BrunPm6ZI8SCLnDIqDzQmJ4tMbIjzP
7YW3CV+cAmAt4qCxCjjmdtKiJ0X+j0o2npnSwbnseGvBZewJsJOEGjLJ16TN
Vb3tCMGI1SEv/6fadY13FHRFRmXfb7g06qQ8IHakI4WtxCKav4Y/TxnrR6KU
jiL1EF7f6Pi3hLVfOTiClmBOzPCuOc0kPJm1ZkUTZh9yNxxj7e9dfcj1jDEy
l49Ie0Ov7oT5B7cCG03eM/p02hmm+QT3YZeBv5NvJIRDM66/weJ9dtp4vtio
C72hCkAcLcdzbsvZJNZGn7nF7qqy+i2QEQth188StLd5dEV8XZB2AsMDQ1By
hbapDqZhwurPeJxR5iu8/Zn6IaBbZe8mtO7p/L7MkdBm4+7BlO95YWGG/qDx
4elk4jYoVeD74qG6NF/EDWtpahRHZCkncJ5Sv0x43PSdIREdXsLwtYrwemTr
5635L/xw6QUl2o2m6yYwGGlFkHVz8EEHgzsmxStRjY9XFdFk1WF1j9ZrH4ad
0D9i6KaS2GvsksUcwuJ9azz0yNsDhySu894NONqKHMzKz3bdTOq9QQ2ge6Fw
Z8YnXR6BZqQz7sOH3MLW/ggIgaqlVe/TCNmNiOnNJNMikNg3097jQsPzSUWl
n+hqj76jR/Zl6FW++TgN7C8d7kf/ykk/ZBEw76ZEBTSMJnmdSz7fAtCm41o9
5N6efTEKPklrPWRNFrM9wDkK8+c6WL9yS4eLZVb/Abt7IPXCNiiD/ZJdK+TY
cl7TjyoNfnBqagYuLrdfLCCBHGHsx7zh/PZt+HIZKd9ovXnD4a8Rq2yVtlD+
X5fFcjDO7eeIvbsjKQ4h/l3LIgVbrKN2s3gMfuy2CtNShDD5in/KOym6piso
EzSdb5ZLwxeJqSssDEXgEse1zijPYwh5AO7MEaikj9JrTq7Xresnmyw6DT9v
c1wXtPlWEKVHtuw8wbN701mgu2qbq33y1Ik9nbvxrvrBLJ8/+FGgJ6tmlz60
SxR0+DC3uGNx4yaqKzYacxQP+jkuIDviQeJtg1MrTW6PY/jadycC21QxBMxk
FINVTI3GCOZG6gXFFI5YO1P0c0nQWDGhZSoxlbfrgzg272NxdwW+/7ysyk1B
TXgwOIBJLxQ0hHTYedUYL8Uh7ZQpPlmUxsQyFPM+yqxgq0XY95VGLTX4xjV7
ACS+CMy4iK+a1cwLIRvG4EdOTdJdgfhgIVHYfYUccT4djV4CjFGLeIedNwJf
w8CETWAzfS6dfSi97NfOP67gMFlRh+yGo6k2FKTkeIQhy9KtHcbLBj6bqT3H
86yJJn6RKa3a2UODMtc/MMz+kgwqj6+IPu8CFLXcNObGgtEr3irxixI/iAnl
Zra6QcV2MdOLwZV54F+o+GJKY3IhOe/lnJH6orcBjEXSwZeBRnlNofoziftY
wEOJoOdYvbBhPXj+WFnymtr+cWUTtqhAXK3aoGy73OhJyNCydWvwQyEasBhS
/OgUuJNcaVX87nvuT6+MUmBL6YatmtULr2ClAhHGNkSSyczpmO7iSuWKYz9y
m6/HC14cEa5wREmI0vxXuAjlHXeRb2ZAXC0hV79RhFo4Du+ggtX6dSwqlLE3
gj0ztH8ij00/ybnLVqQteN5lQyJhz34bbV7NP3eItOlhgaCr6lthEsJ7Uxp1
hUi68FbeDlFrpZcX93bGqZym28HFvJDrqQEhH2hcwLK3pdeW9NFgpP2QvkyK
LHBKvvPobYB032hxNls91l6ovQza8lEk55ArCp7ip6sfeF74k1iUd7jRMQT7
v2869yAbwI6R6tQBiwF6efHoCAmr6eqpO4NHmcXKdu0FfXzky+Fe2M5GzZ8U
Ww67DDfVkv2NX97i63zlSigKTD7+7l1PoxtEoLy6JdbFn1zPowKu7KVC953e
hwXOXujjdVuRANkgefiY+jXa6kcSEoJ1GIV6KGwUfnh9HJ/ZcAf8+q8KtaYs
Y72hG2nfr/gmWq3SJK96wXJWxoIFbkKfZ9DhbSjMeSEmPil3xDxk0FBehxaT
HQVuP9lA/Cm/NRLOrDASZz8XfngeSB3kOdLlP5fJCODlnpTwnIzXf3BmmnK1
Hi4nPtz3kbAmD4m9UXFIc8zOA8fG2A63VAGw+LXaDYJVeCKtkoHQdfb7pfri
VROTud9cOpavbDVTqbONp9xD/MQkaW4SR5wm/4mmGnb36PmLLUnMIOFRW4+1
6dlhJMJ8Na18w/oDbqDOeGURguDr5GVSHtx4BXnTx4/SqKyH48EELvHtJCiS
IYkEUkK71sXZH2X4As90KUUmt6t2Gi070Y72ovA3tGEaFoH/4xpnfhD4tnUX
F8vamitqVSqb8GRDPSnRl8tub9PfhGN+ZNh4qbiubzqAKTz9nB+lE6IY5V30
BunOL9Fd7acTiMHHKXcSMpIxNuh/nX38p7m15eS0FuMBa1aTEJmcpxifDzbj
iQa5ZKW8PPUJv8ofu2O+5K/TllWjCtryOfyJL+eVnZlt1/CmoQ26OWN7w/G+
XCswERVxVD0pr75o8UmWkVnOYFotOxJQtKIrLVBDPHqegUt/XDp52SK0TcjP
HZwWyHXiKqYpegMbXLn9ryG9H3fLBRI6vxc2qlRq6dQSur5XrxBB9PcvM/YG
XRcN+r5Bx5j8fi+Rrh9qVR3saBrr1hJocffIVJQWF6qtZGpLpMFMal2UfZws
Yc1MT6eH/DAfgcR6oseqWUt+IJWAuszSVWkDFkXYXd/p+RjlOTyNw7SoGeyU
HQnk8wML74lwxYhfoFu6A+DDtnLPs/qWh4x0EA5vMk+ayT0OtwpVkutf4ukF
ZZMVGgTA/eeDwjenMh9ByNZoUnObcJ11cnE5uKUdJjuWOv6HihIoZiRT5lIn
Vqp9PIM/aJdIJ0N531qq3VToZOq4dL4JA4j41sx8imp6rBRWiAb9i5Ci22id
ZtgfME3wxGoutKzoymZ8TWMIVxeLY8oQxF/kHaasoJi59DDa/ogd56PzMWYI
IKMC3yMLt/UC1PLTggtoa+bj3fqlzzn/e+aecIpr41UfKpdkVLwSm97PD9VE
Kv/b0XmH7GyONIZdSXMSUmDqbZk1RiWTM/hyd1qBgYijRKkAnpEQzJIpY6qv
/yGxeP8aKa0nScvHS3xCh26D3sVm+kKZsgN1DrW2W3Ic/fAtXIaHXwmEa0jI
F8fJOPYBfPP0d2B+cmZ6v2laAjHyowRKiuEmg8oEL7jt1tci38nRgd1eO02z
hjRfN84ANxVDxqhJcdrU9NWfJp/pCORTnzhX1vw1c/dfKH2piLFF518Zmt2c
NemOjuzIEDPeMu1/YwSrvb4iGRX8/62OD04dTRe2e54uv7AWKL0RRiMqkKmb
wUjH7AyH5spXuFOSqtIdM2ogb3zl/MTRdnU5m3Qj6Oc61VZBNJZ7Jtuvw40A
Sdo08xUxmQNy1pPJ53zUr0Px8adiBuaq4OLTKSJcBXqDvD3g+uOon33ihDn0
nJrFWuuvZvvlS7u8d1BPnU6LxQt/LfpbeMlSjqZ/lXNBELpuncVPTenscLrT
7zGG8R1IzXTSOSMUfTNAMs6GSg66kXfsoxfIRQTG3sVjikwt63DNWPK0QG+u
KwMWgPFBlReUekJK3xLll18aiK81shrqon3Xq8O/0yVg5ZKzbCJuMs+e4irV
iTaknau1oLYLA5de45edTwwDmdCvpKUDaZgxdqRZWRTiSXZafAFXysLXJuLk
Ai9Qx5KmqoAfGorRQNmRBi3RDHiBSu1ZJ3588sOQ6EuUuwXjRVFhD9El9Hqd
i4iM2lx+eGmLCrlRdhDsXYZjKp7U2M6csvnBEJXdqH6ZdUAUAx+wwamT3YAn
ldko6+Mi/+iTvV3rBJ+IFEkjVUhbZ6f/WcDG7x7IHXPdY5H84StrwbSV1DtO
w44otMBLI6t1UL5SqY0sovQwAg6G4DCm1ALRyxq6skpAlOtR2F06qKYq8NXw
05AE2qCEw0V0zTQJXHrbw9Y/x1wCh+qGGmaEO2luXMfjDs8ZMD3tXQ+iMvxG
zw/qFNoh2bGQTXM1GV9ycWgbbDWAhAp7E0Q5rI94pxMqUS7rGI0h2PdG6tMp
8bS7Wat0+S63cnVcQz27hFWtCuKRpuZeDsvYHgifB2z8LWrvz4Tk7l3rPD+c
qTiLHsEs/Thr5SyOH4rdpRUYg7YQDxNSo1nfz0kbaS+Y3dCMGaMp4qS5CEzr
bIRLA9YbnEsXXpVWDc3QoqezBYHrqYWVvyxzi65osyMfi9NqEx9nVvCVPqg/
O+X1DCeIArzmSuHyRiHUWVA/8LDFOZRNlPtfXkHdvZ6uyQWNVq8HImxUs0MP
FBuzfQ/hnfNowN6ltSz2SQLPhMTVsTdYIM+C1lFtZEvo3JjoM1Tq9HBDeOg0
LewIPkMfehyuxFhDlgYqP6pB56x7ls49sY75lSJJlMLdQZqXQ8uHQPBU3cA9
4OMuOmDdKK08apZLPhkJi9ULe8OGngJoeDLEv9htXwfWJ+Psb3OrhsNb75uP
jYRR4+Nk7ysbxEw6isc3+zj2iqRAOmFUNlbBQt6coiUamEwpS/EL9unEPdOV
MRjw9+H2E1bLKaG7TWwme6NqQz6JwD+oAjHkM6QbpTDIMMGycmj5XVo5VZXB
pD8UpPJXKtgQSqPc4nm5vdiasSUeXZWMGLDvVjlBtGG/C5Y7J4GvRBzXoz4I
oYnhi739qlzZmxsHmIotSMWcS3gEW4DPKbWs7VT2iOJd3LIc0hwcEdjU7ae2
GbQukl0QLKT3pSSzbN6Y8ag76+aSMLbMm7UYcrA2AnGMzfkcwBj/1O4Oe4xU
b5e4XuBsJN2FN9UxqeEsQ7uDb88Jw5ws58mjGENHkueKr+tXlYTndgDxJBxs
3g7Wu/XqsZIkCXly8UMLBNW6eRYksGqzfQtJYkMjZzpO8G7aW9ftM1ieQYhh
nrZvwoBtBdDnJnfh8dm0+2h33tFxJfI0X4dBx2KjiVHi/DZrTO8T1DBDV02q
DETAhDaAx/vtD/fcjdCw2OxqzRa1ck7iSP7wft61kQ/J9EKrKEyvxyAiYnQ7
Bxwjswrq/Rpn/Tff6/DTblm60T2U+CYxqm/U3mkIv/M64B0FygXJoGvYLF70
9uWWL5qlaaXBta0z92zmWNGJSsWIG5U4WyMZ3TVA/BNSSiQoIzRbMYSw4AYe
ykes2skkz5rD9p4/v9agZarROalWrbAEBKLbsscmDJS9unsuUiVyB2iRRKNh
qwCPTf5yMEiHdGJje5FxEs+FtAVxoXkW5U8qOBqi+3WnBjZtbCGjAqf07ezz
aLYIRIWpCgfuIRXzcHlfAzsT54TN2FbsGeGz4qkf/HSzGpcCnuJk/86hzU6P
PyPSJvnc7qksfcu/QAukp4zk58lIyP+wh+COtSFcZRgmKKaF1wxQAvV6s6kK
XlccinDp6H9/0qOTOG44WJa4Lu0IJlhPYahx1i1VV/WgGxtcQtFTkY88xt2e
LlcQZxMFQBNxQZChv+XzLTs9JBoVzDLIUVbudmRnhftv0oiyoqs3o37Q6rqQ
0Vnf/OeYgjL9q/zAYznRqkcFSEMPrTIYXOruTUG7mgMWdsfU3LbDOLYgo/a8
JrGcxguCBdN2ZB3lULqJ6RjzBRIiSRwxj1CqoGS7zJT/8ZFt5ZPkRYnYB+9Z
dLC1ZdUm0wVuXMmjl6XJgHIVtqJAuVSHiXLJrIUlcAaae3BeB0SFHf124QpD
YxzAPqaeWUGRlBKvVwYfzehEiBU6Joo9gDj4880xG3eoxDx1J577eLyI+r6h
8I93M+mMGOLCa74ZNspoOyQ05WIEbrOVk7S3TUQuydDlGSaFM4XCaXUCKV5f
CIDkcKSCUu52YrmxqeiQ6rvjx2ERtYDF00axfi9z4d3/sbmVC5wtPI074pKy
CID5rJnQDiq/EUwZ7+uF2ZoAs/S5wmCnDVt0WTNqufuwN51adGGA2uBGU28Q
PRDkI99nAH2EQtS36TVGGud5s9miab9TJrXDDBpdCrv1VR/S4ycDzaChHwqv
Qdwtnv05vkCMg0f+FUBK6botUpJ7UXa6NpCt2J3+cj2cYqbCs7I+2QCKiH05
BsI6lnYrvWv0dEEpKHbg3ytRwTfOiNfjpSfHLo06ecP3uVZqADWpuL4aN0Mp
kh9ChcmI+M9Grm8tHg3NWK3+UAn+ypnCvQGdWRwhzKuHQfJBGAS+KqZnpmL6
C7J3qQfa+T9mx7s7+thHXV5yfE9Q08HLBH92Olc1hrGQkFu4KUmE5ifhx/Nt
rFilsU0g9Xf+nlBPXubVa02pqR6ItokQga2QW+b2QTphaeDfd76gCNjt5B1J
WGNf66qTqUU6hIWADwfiH6yRsD+ncmF7WXZQADoQxjoA6CGRkPb0AoqpRCEn
OPjydSk7wArsRmrmcrbQQRffeOiiurUENtzrKExNleB6CmuoC/sIHf6gaZ5K
VCKDnBIyHkFcEvJg/z4fg6ENENfu65AjVHujx2zGibHWQla1jW4RuMJE7Pim
aiREwSnFU3w2II7I7cKXOv+ZNPW4zMNpEJN9Drdwo2HmNb+eI3MKFipbhiDE
WHhlfWVaAT+bs6qZzU1flsnNigUYh98kZcqnA/kjswP8wlT7Roeix4GKx3K/
gIfUhbZy+fHZXdrTHKdiqxF7+2QeuYEd+xPOZFuNjSs3WAx+BVb0QIT+imxG
kYfeMOX6Wpi/T0XtG9ILK1lm0KXQX5MIHw/Yq94Y9EIocdV0k7BFO8J2P1y1
DhNDVuGhAQrEq557ngWyEuryG5Ls5JlRUTQax96IrdhWwHIo4AvIpRifVnBT
EIlJoghzLs4k55QHJlIeBLrdjm+LwV04eL5vpKfW+SdbMs6SRVAFV4Jo6LTE
0figLVXhSqOhRZg+66slMiHz1gP6AnVSWTvrPrXDrnrwo0OGjdqk7sWRDyw0
2jYvkV7AB4uLfeCFpoQLz4HVrgs9AfM6oIedFJTM9puOdyUxJJnD/pqPK/c4
x4m/oaOBoC7NPlfGLxXLcUDAQ56oHaivCKA795FJGV5VOqN0iz099yROs+P/
piONkoQq3CtC89NtdQk9ZAXO1vjmhAkK9m9VWA3XS46ekmzCm+kb+hXfCw4F
CPltfVpHeyi6UC9OSqMG/06QweWUJtPSLyHLY8xF6NqD/n6sx5w8wSfLPqmJ
bELFcw33S2qyMaw01hY39V/6XioAU6Mi9YfbQ+xpsTqnnx7ANY5fhXE05n+i
k637fXjZj+Vhps02Hjc4tb3ybzwJxHnHtYPMv7WwUfZsBZ7gJ0Vipr5o3UYn
Knq/oOb2V1zaRGg+M/+DBp+hm1vKpWV74uKVhjiiql2KS8xysMS9HJDRsmk+
S1ICNOZd7JmP1oJx4ZFTU0L/JTLam5i7eZKXQHuB/wFXnImykfkbYfIFJqN6
/f73ucyfMnMcLA76wkBaVae6X+hA294edMBq+Ixcaw7vNdGOaMoKO3/GaMhy
WwEU2VB7KzRNYDMMUs6WPXLNaYH1S8YAMkI/2ihVPshzVk+fNHcnhsav9inW
YUhDkZYd/b4yBMuDgFKnEYRkgWnQTY9SdiLc7VlhG9UTzhwIpASGr8yfiqZ7
Dr78DK+gvUZdj2pZfhskRntybGtAwBbgRRZavHrlxoO1NLAQBSPcZoFj/+7r
92kTC5vu+3E57Fplm66rc/BHgsd7ljqsT9B+p0uFBpZjmebTy+oMgozfiXls
iZzvv6BH5HEtZnPnhC1/yC0+CgN5auTYy9QT3gTexaIWFZhFDX97P4pEX7Kf
v0g2AsgMpqPzVBsq6v4oUCdhHdIKWARObzjj14DmuyJv//mgnTpP+tH/9/zF
3nR2QRz7uy7vgQSt2d3obDvIrD6co5OotwmxbbgbbjY4wxOe2Jh0iSDl9oEs
ce/pF4c2iuMGQrxyunBDUgdv/j+MK4EcFgY22xKHPLqJhBOADGZ9XL9zWdQH
XsopY/7O6R8WFfJu8pqZJL8f6PEl+WuJCEGk6yZItSVYlA78KRXr4ef/5RPn
jCpEy0+mJHmxCwOBObb3DS9OD7iQInpZvE4z3UoPa59WTsBwC4RA8EsQMIyw
+QseIbMDAmMRS1EbxbimMvnJjw2BO2c4IeUQMq5gZgFHX+LChPC3VYnHJwTb
+kSyAh1yLdWW/VPq5esoce3FQYgAEGdM4qGKtdCJmzwGPfYSsowB57VXqJPE
2YtxgHOu0W1DR2nYhMhH67UNiQh38P5sKlq9CW98VaPfXjCahdjSxnXcv57p
JcayJ6BVIOPwzYHSL4iHAVOS3daORHRYvNLPpQMMM7W9xx84F//rfdGTiJBQ
ZLmSa6GOxKiNObD0aoZRf+qpx4ndLIZ7eu41f5Feof/v3r79nDAEh8DsDsHY
ZvyniYVG06jlIZ2QVKZmxK2dwHP/LGOWcnVyZ+pLaNwhH4J0x6WTBfH4SCvy
JYyF44OE0w0EMqW0iWvjIot44cSHj1Lf/MTmwQr8FQa+tpIK/0Bf93doNRB5
woYgjDwVp5/qn1rSFZaYQcDOBFPq8xSn8Ss/7hH7G+ae82F3XgMfPIzIWWTr
aaO2PlR7tRZLsADH+ZdSyRhscUT6ligHJQEUDr0OP4boGAt1xf5zlrjZD/6G
Rd7blxfwRt3BUEHrEk+Hu8lbYA1C3qdoOaKV+iRG0o3pQMB7duQ2vSOJceBK
7HFEfPVCueuf3utQwQojlP8TUsHWGgHhw+4JozP3scjkh7ktA7e2pQETMazX
fc7aKZRrjtCGEDAi/sBZha5tT5U7jda3iqS7gJ4sLjGWcX0fVbhvv1BYXBGk
1qX0UKTbMf55MlUWRJR7BMc5XYUcuE9WFICSoBljsYs9+ZUhPdqD0lYm33gM
ymfZis+I8CHzuuUi5OoVU/wJ9yQ9Jd4q0Q4CxwGlw2jm+IDfxKBVPxPRm2Mr
t9QrTnfDlwcUZ3ZaPxY/p6GbFMxAc9DXpQ89mRfd+kq+iMiSJyxqItTiW7P8
FVk6lQS9JpPNuE2x5Yx3qht3lE2nGaMPX+DmPbmp+vA2JXZOrGtFc/3WM49u
A1EYmqBEefqpZ2OiwCo/rY9VNLfiTMzdAkyBV1B3t5NbXc+IjpcloWX2tE5Y
7zX2gPF1lpMeTuMiv7//pGtB0AnEu54W23S1uD9DzXol9XSf4XNr72Jev2U5
gOAzQihTuhWJJMQTUogfXUIduUOWgbs42hUqayDAIonsVPjqbfRVrpBeCGIb
m8xkDssyO9GIac2U2RdHsLc2h6yylJtO1rh5DuV3HpOeglDVSKwakowaJUq5
yjFtq0r7T4HyhjB8pHuxIOVPgDiXTBi75GxjIgD+WJA+nMsVikcftViRl+Co
i4Ih+HJkMhCYgQVBTb1nJr9flkRetouzhT8Wb+3bsrHv4EiT143GvkpLndI0
QAWPbv9d25k772sqkFGzqJkYOjiklLcl4iVHvIWaDcvKMt1c3agye3LUkOv/
eM5KPxH9wvykGJ8Zomxi8TOwkbnDGZ5+Cil9O83VbinmYBh3oMCuEumjz0Za
VaX3tLtQMbK7ehcxdwJK/7RYg43c6uxOYyMlGeCShLavpVoqP9oxuiGV66BJ
MnY2M69IgF4+DQZ1egO0b8j9gJVpkiHLAOfAyOcArOdLlCWJseAdXNVjNHZJ
sRWLHGMcwSwK891XQ0fMLMp2Zaxk1xE/lTJp4K6QdZt/51zfdD8Md2Qvx/Jy
tInC7r/zqm4iz1klyu7kx+C+Na9CyQCLT+0+9TNkgOQEQUtyNDdW+FKt3x3Y
yDvZgcU1LyP33ICvonMG01+O+79HdG/YQH/Q9TlcgOk4JK+EqL/q9rP3tuKo
RfjOF/KEVptfba3nWvy6pJn7vA8m4VVTm10zYvf14ZWzpvZKpJV932OxMo8m
rzVAEDrLiEpvXxTMIb8WMREFUH/lKHWSEe3YjlCmFcbDnhwB+UyTvydpZZhb
q7DLaQNCYCkVnBIRX2dJ0Bk74WDWvUggacCeJmN6rT38DxqerAlFG2lX1xze
gNOEgukNboLUjK3SowNTFtpYbQAEX/FnQJj9PxJhuRwhi2ab2UiyD7iiHlmf
FpSvRBajEab+e+AjNECvbig4Gjn0huJIzDoj+v8K177PjQ7rMlf606og/Z/O
gZh6uFdkxJbKAVszhp2FYOU7QmjsHGHj0C/XhT7bPi1+ZskcYJAs0L/Q5l0/
IP97WQE+Usq/yZJkGGcGnypgRPrAtMjomAJzEqn0rOF5h5Xmic7exbsUP/Z4
NMOmXEDQTgmqLSG7413mvRCzqlNChL7G/VtmC/Vp4BS6zEtnbRt6JRCpG2x8
04ruPNXgNnVQjTDZc2iImpERhXGFfzHssH16KOqC6KeCPnIp53J8r4JdLa91
0LACA2oi0EZ5N6g69wyY0JmAn+RTjPs9KL4hWInHWihFB3bAtePAkPXevszS
4ehSIPRlGQa8MFZr8+7/aqun1GNozC95uSG6U8WtSTVWawGPuOS5ziBuuedx
Kn5F5BbTVb//vwy+IGtG3X34ePwJgtxLlZ7DwTp8CMYlWUmNLBWtGzZiN7T4
bq/iculPBvQ3bIhESpCzKnDiWCNm9G//PRXxnlKYIde4Ii7m7eVD87riIflO
k2sjieoq2e3Ic1MWEbplxYJ6R3RIMPk7+bExQPUxgSgdW9w2KisVSR+lBmER
skDCq+jIwGiaEC6lxwqbgwNRNjrtutqbh8DeY1rFYAlTYoFonkWa9OS+CMcj
B2x8R41aSjaIkJqer0fw5ZE9vcJi57xR55bwgelUdtt+4f8k6CO5zIf8b8Y=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyIJCa7N3rfN55dwQXtMv6FbZBeccUsakqQvB8rgpHmeonjw/OYhvxtCDEqAfu1hxKzxLrRmJd2GK8TR2nvnjHuHDJ04ryg6BbtkChDvYxgps0o+j7q4/NdzbYw54B3/+D755TEaY9mmM/B7y2wQnQV7dr86xPsH/DKSDzU4dlXBRKT/bWs8jJZrxHS9gLutZEUx+9gSGoyp4k5mFek5qCL+Lo9c6TKeyVQwVp/TCymEWJhA6/WSI9cggRgye2prcRzJff3Vv4TvWRnuGbsVRuMJFXOTo+VNL+Ksfi9Z6sc6PwV7vvSPGXtMqFnAIxcEwDlCATWrCD0Xc7LheUJVO/swlPxlDxJZb8JRxSJPfHOwoajp/BjV3WkiKWxhkbbd+yWP83J9y1EatLMq12v2Q4j+niOaRmQ24XfJeoCQKYcZmFlRL8Bqv16Q+Lfx59vxFctR5queKmPjp8YGMn42jC9dxREyLgRDTeRJwpaJdOR0bavIX5TNBfT7/hE3ynqfEFEWD9Fq+GWvA2HZ0WIGBy7UHaaRRiJp17xrjNC2ZVqS9VQSHD6a1V2lsVtkEcAL2U+R465r/dKz9LxbEv5ww9UbGEAa3e58dBkZEzFavsgH9P71jEZgYAT4Y3GRNV9AYb1p6zQqQS9S7K6kg4InEvN5qRjm7dr/bELTEaLd3S8bzZLSi5ffuXX48Fesw1nScu5HTpqtVL6a8PV7PUv28btjH/DrosxHa76J9W/K0fRfeVPrNfYGGUudZwqeHRGbgDRk0IqY5vXNVOLtZzeup6pp"
`endif