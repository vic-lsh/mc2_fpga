// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Wsl1QsQUjGQHvVtYoCUFHvgE1viNvoRM9PZQeG84+3le5KzYiB0ShIP2CKR3
Y8FQtvIQoMwmSo4Aq3ll33uz9HWQQBgSpAhUv3dMbXKhEFLCLkpBtVg1+D+L
PNT0MOf/h8qwQAAzlhk2W5kq2ajH82rqgSYW3hPKQICvCErNb9owzZvOzY2G
XajIn7W0TFMJVhWSSMhSrkwRaO9EoPWQIffzlqDjrRdIUg1f7jIWFr2o0DOG
6I6Qf0OLu02fwC2WFrb+po75MDP9nqJDgnw3WUxMG/7u0ravIl7P7hvEkJrc
N29f/mYa1pb0ueoPKK+8J02zwTFCxLBDrTa/4BDUuA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DpSdoz6sooy3P2OjwShlvZScrSaTbNgKqzrX/64FQ8vReuLu+Y0Re6aAFUGf
1MK1eLQjlscgYn+bog6Zgtiap9uHQuhdKUfT/kREuavBQ/w8wexLUNtX6sas
fN9XAmIDfJM1bcGQ0d7a/8ZXy3NynQWDLwXhsZ6Es7wpkHolgmwS05o8Przw
r92uR6BPt3LnJXWfyhPLmIe8r6ZxLBwEmv5ySwzdwu1EwAfTZ0aIg6M7IRyF
08421u26+ZzR1TKHYab9NJ4Ug7ydK5g/RdUvK0jHW99HjYZuWIyNtfjNM4DT
t2DkO5fhATuvrZNBcbp8PQdByuj8c8nBahTaHt/SLg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MsT5/uSMOagYssl9tFpqI3l+UlGXCMiX1PCmB2c87fPsbCuaBJTMkVOkvrGy
FC7ZSx8y1RLLntWAAjSDzPxhYDvEyXqW0OLqEsreJ6mK75a7cT1rJNkyMIjx
REFBsAV/u2+ZebmiMVISeB2C7O81/Q3SwDlh0ez1rWKfXLvwmI1ol6iqxl2E
A5Y/pqmMFmj1/IvtqWu9iLj2FlrmYCah5CnwNpd4DHKge7ipHgazjOsToqmL
vl490fuIS/AJ8OA4Jdr0Ogh48ZybWOM+YTlVIfQNEjWkjQfb4//b9r08dOYB
uK8xEFKuRsSfD435DKeux373na+eLyh58IJB2W+InQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S8h92m9MtMNF/3IYFD2mUD8S5iSNa9ZIwKpEgLbekR6aVSnctHHNFZHXc5WB
t3aCWRlVvYcNoGBkfn/4Wr7JGFZ16mTEOZ9bvDsOfPfy80tsezdDgXfgrjhG
qONdVE0R9WJWi4Vb6XeJFN8PEJYrilyeu/i9ugUrW7skAJCoVdy6FbMhdcyf
rWx1TBbe/Ymy3TdrgK/TULgMQDbgiR6XLO/t5HX0MJr/pV+6hZt4CxGJ8uA5
73HqyDZQY628yg2fm8nyfThD3qQIAtda2cyDjqqk5wGNFevOOboE3w8D0gOQ
DZnVIRFdI7IZCOVBNz3O3HIHl0aNp2d4gcsSKKhpxQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C3XtNwFyZUa9gesFuhcgimIy8skLZXHeUFnhM65QshRkXHHdmOZXX3iv6d6T
lqqiLBoSJ6MMy7qBEqHSlkd5PNl410+BqVcYzc7uFpzknBbw3BIvzKZvQhlX
WUkt9Uj3n8IdkeUT/W9zdJEjinFzn+fizAxSL9F3czIWWCOqtYY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DuWKaYTYU/gCMI0NkhuAzFtNxEL+nfrvX4b8ssaYXuNIxJE/oQTrHUD5wDhM
QEXQMuEJiUGeQDWmt4HU9AGnMSBLEFAReSLD/3kYs27KiPVLjsbhUUbLhslQ
87SAwvQIxw+plJxEOCZpM66dmis8DOSDSpiUBonhN4dHbQALQyCbr9zCoG/o
mWIslzDAP28q94i2+9Pkm18DuQAhZyGfLfTGmNIn57vDgutx3MCm97nXeBMY
WtVezOVvz7a4CCFt0TVRL7zDKUmANrGUTvAv4x1UYwAY2ELVyJm4CvMdH3Eu
c9UvJWNdboXQJnl9avkmW3vhhRV0Z9GBG3jTpj4yI3DiMRv9zHrkS4axBSdS
m6KUWaNJ6PU/PCOXV1Hb7FGVj2pDWF72vPxzBvowXlPifVz2z+NXwuCSFzvl
IDYSpBLmb+iJjOgc4PxeH5y+WyyDxG53S/AmiVen73R+8zfrXe14o4318NLq
I2aaKKAYGZd9gIaPIV24+ldA7Enf2V0T


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lNEcsCMri4q3MQAgbcAEfW+GJ+qDYA9KqNGUmUDee7x2478WOLttWkMdou1l
uhVY3YRvc8R4QDfPhcRxMgJ3ml18S/FDyEf3il42oYd++45aIVeKjsUoFm/c
8iVuTO4/K3F52XcgYH/D6TamviX9zu/mxavI+JHutjqeABSJIDg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rgWD1ymcunEkA5eJmnS+egZgGRdRAupfPZs3EpeXW2hwpiI2C94X1FNakyvJ
y+hkedCERvGVQmjiznt5tv3+l59PRadM7lgsAu5jy5FagM48FyTNnf228ir0
Z265HSH3fGGlqMc8TX5xfyZv3200NlqTJlrby5UFNXhl63remD8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14400)
`pragma protect data_block
7pNG425ASK5s/g0/x4PKRzoOXjWsupO3PV50n86FuSDkp7ryEZMY30zlXtqk
Fc8NepqDyNlQBNCpzxlDIeyHTKK77Q3MyFdwGXroViIJr4oEPKQGP4Vc/W79
YGPETIzpOCPcqtVRAQiNczDb92+lIsRDmhtVCAOyCvu1MyvPX2q2PrKUwjvH
oDkHI5ni0M8N3+wez1yxjSPlr4EMHmyBqixiGxtk0yDYobYcGfkNflz+Y2IB
I7btbPc6viELPmPWFYKZtpMRcZ+VY4vBlwym4SddNxwrcLYTh3/AK8Gmffvp
A78p0WVEFIHsgRsTD94Dq6w+yvd4LoFsu45WJXs+C1qJtRY7G48Udm/T74GN
URg/EgtyoS18bsnP+yZc0TTAX7BI0e1Ih8m/0tzdcBqCV4L+NYU0sCE1HCXQ
5noj+OJRb9x8WjZd70sIGY3NHsjGT2jWMrCqccOtqUPUKnNXKLnvURvKRzAh
Jpo/iMMg57WcbdIh8eWeK+UWNlM4t0Q1UpMS+Z3mMDqceZUdOZuTdK0YyZHH
PlNmmjIo3S3eji7/4LQSUbNp54ZyrDhBdBOr8UI/+lVJqxzkxQucepNTkYS5
/8AIOckmWJLJNWCiinUi2XKN5O7wUlM/gUsfuFV80Q+ZPz1z7kLX3+zTR46n
m6y2PS1g6l29H0RO47ioFpWBo5MWE54/b8xzc+jUdplXr0qos4+r86euxqQ+
JyPp3zi7zGMLToqVGOEWFjaw6JlYarfv6SprtXIy6hkYlLYDBwC5Vkkg86BG
IDKU5/HEgFfPCDu2lm6pvUpS0yFRkAe3A9rHbd6LFiMobnKqryjg1VW39BMZ
5ayIi1o2ndlMHzpK/bPEQ1Gk9N6ufUWSWI4Am75Kn+cxgev2fNkmf2ZL4slN
4jD8h9kAzQ6kfRJn/JRdKuKzAh/w2lwquzjh3L9srcupdaXfQd7h5TWfjwB2
+4kcWK1pxK3EE5fx7Ww9XiFy9T78PsoTyIhqyg8CFJPAoI0gDFAKjwjwn41T
+m6WAKQJQKY/p41ZjjR3+fwuImx1KBOorvV4t9O6t3M65lapkKLW9KZ2legi
N1sKozV+GHz/P23uUGjTWc/pFNwrbaDpHZobdy0RowzxJmf6U0Ssgz/SlIPG
gQdeDJQQhCkNA4e6rvTtp7yGMc+KStk7Ti+2k145uJfkSBGVdeBoc2n7h7SD
HURX38ke4j4X6TcWlSwaMsvtK0oUvUFyT49kMsRYyVhZ90HvoyI+PpM3KgX7
Kt0v33f4KIEZ/RQi9VbpcPibbb2b3YAIngSMLgmDhp8pjO0uduwH+9d1geM8
eLnHpK0E/QmbbpSCBVWV8QHVxQuuFUDsYZWHTLIkzwWed4sMOhmc/0YHNRss
4QEowsESCQiDUmF5wwHirj0tryehF7tc5eJbzwEpSXEio7enpOSD56kfeNKs
cj3qVyOuHWbL+1PQgkfFxEglAGzWR/rXYbpYfeQEZzguX7ZGJpW5x0lD/JIs
HJ+ktcuNnEd6MCYwNgwJib0oRmBW9q2xQwTwnsD2i3Po9SGrniATNXuF/PJ5
sljoJqTdIYfvTNlldiWv6sysENiYoNgmjknp0YH3GGzSMtnD4XMxzhsAe6Vl
HYDELSBRuuKPgjB6kCZfPPDvmvVnuJIvT1/8MgS/FCRexEt6Ah5eejEoqzFD
P+fiLhU+5NNk+hVdekUO5HMHRA0MJOTM1IPK6S1Pe5iVDyWAxCJ3puMKqH2z
t54G8dwem9OIXtTw52EveSRaJ/VfLnKWseAOVo1K//kpMYcJ0Al0jWrHVTGg
7Lz+aTYHc404YBpKGMbRKgYWDH9worXMJlJj3KY7NR3opRDsgHw9kPv5QMp+
zEDv2NeEHPIMyyoaMgCp280IhJ6GNiiXkESQ2v7uUjHBc8tmLwLtdnyx4Ked
7Zh6VttNXQ4aamMaC1d+OGOu6uXuHDip+2oeTdmppIRWpQPq/RL8KrCJ1r3A
p7bLqzj/XKn2KPyOguA7GKvp8CIy49adX9ole4/AhbZpH8fvURzkirgzZRrn
aF/JpHZKurFn4XN4mIQiOIEUhb7rWS98nooZSHwkZqH1L7m2fCXVigmNTl7N
mGpsMLLMLY29Kg0d3VLrfHxf66KnGfV9PixfeKKYt4DzV1sM+4C96BZO4Bt5
i3//a4zy2UdydgdPYraCPMizK36K0ObFWkpdMa8RftPa3zJpIRzqpPwcGfaK
0fmOsZWbtSQPLJNS+yvCLXS8FxtMsGJig3BKxAgKiziMSy89bMcuWXdd0f0y
JzxzNo6Dmw2h2IEbDU6k8yK0DFdXXkP7EkxTABYN8BvJF3GWce3zR5XCQ4Lc
jKlx5A7U52lqnVYQF6nyiifkV7Kh7Cj9KOApvJ1a25ABpLwqj3zbTEblO7wr
Kf05zc4nXC9B2SJNTZ2TCxrIU6qFPj/Hq1g0L3MtXMgCukV04XryOgRFR8Ph
mzVIEpkYKwX8XMjONNs7Im1SyM2ve69AlU5aT78RdUzioFg2NHQxU1dmxOD4
95bySxpqpffPqIfDXhrc984Zf3vu99APdPtHytLzxsZriD0EOtoD6TrTV3Dc
wtnKxezOGrkd+EQJQTMG7/B+sWHXyns5zYpBVQkirAPpdVNqH6zEviViC4J1
RhmIbbOPAPmxp57Cp0Q2BmoIFJRTcp3ViM46AC9YLxcj7gG5BPAyGCaaxpn/
gIJZDNjo8/zu73zJDM4up6iobjaWDOoP0laNcxReHZico3LmKZf/1wC3wj92
AjdFaJW4kMc4AsF26I73e2XyriCg8eG27I0ImD6/MqDQSR1hnitlW1cFCLbV
gMcmzgqFHHWZNW7EqmbPluhkYf6BGki1rjJegDY5IuSXzbI+xlLd2Q0N/LUf
+cHPM4aXhBWRbsDoUhLXtTlJIW8+GJWjePhi4fboKgSwn4/jCMt3BhjV/8Vq
olTD2XgtDhPpfyeCeK/vaC/NY4rPy5fPEXK49iFMThlfsUYm99yWiYMN9W5T
lonhC0fgRZyVD1jIRSodFKkkQ9BllQrycQHNxHZ8DA3SVcZwhdAwWFXmmjBj
W33e3o/R7QWKOU8Z9cou3TE+XISmTEUnxpAtTUFlMQ52Kqb4SguV/1GsJGAD
9RMYK/klVrTCy37vDup3tJSoHFEabip0bDCBKJgwVPvZagojURtzQ9owi1bs
qK6ZocbujC6VJR/xWoZTgATWDCC0D26IFSnsEsysNYQykVy/Eu4wMPW2BLyu
ZpKaF5D59g3n9zk/he0LAcc+OcchsERuwQWttY4ATq/oFDp+HTX2vJsMRuPr
DYNcKvSyOQfMbmi5XP5tgZS1AmNtps721DW3J5JGhIOjY3Rm7ikVa2f7MnMG
+7r0iKcmvtJvxuzny0o8DlRvhHgkLVQrXy1oHyXOmhktn3Z1yplvuX+EgZmu
VNJY+Iyk4unzpF/HsNRANyrRibwGm3pXgcyz4hSkjvAZP+PtmlPqYdeAQQJZ
iOtte2+cbAQRbSfAiFKIxw5+2ho+kE5+LGC3uyuD6pVQEAwpG4VhGpXdFvSk
qneTI4dzGevw4jvfwaU4iq7oZ8VyExoHjSU/5IgrM6qUeJdGdHPyAdI6KrsN
nDXpFea1oUMuVl6u2XvS3UIKtpmmgO2GSquz/PyK765gWHKj5sZV+Y1kLqqE
8BjuHsJ65/Kaee7Zi3J9LpVlHbLjktUN1taBUPZuytV8J+PYOT7fV4vQY/GV
33nXeINEjVI0UZ+vP7ZYjlqtpOyGiL2mFRjrf+int8qpIY4smmEWSD1Bo3hC
PZZ0bmPUiSKJTwwEkSI/+AfwJcBicIVclhzGgCaMBOA39Ku85cvsUWwIXpCD
knPMnfGrLY3TfDK3C98Juz4Vyok+6FQssGmlJOhv8bLWJbWM0HElFZRG6scc
qZu48q43PxMhxLU5iHqWL4t1dJGriwStYF/JSyC/ksQBCUxWUrihGPmPvm+x
Bxzv4C1WQLAhSoKdoIEa8KS7pc37Y1oD55Rg0x9m1fWpru4LiplBP2F8H8ey
H27QwHRNcalnWwPcEvmS8s0QsdH4fIEOJxHGCLmAY1hBs8fd3RzoWrNSkLVu
byWmBYVGrONMN2nYAL/BVD5tqMx9la4chUFhLi9avR86CpVjhrgSDx72PJr0
If2P0ChhnZrX3JgMsL8NvUwsvagnlE56Zc3yQ0UmgwPb0Oy1tla0S3Svtr3p
Abfw4b6zMJeWbmhQ1BwsMlpXXzVDNF3QP1W/VF2M8kluLYTjlJoFmknb1xZS
86EfN+ee+4xqTzs5cytsOzR5AVLl8FBTjPxuFuZIDVJClWz2+N06M2RY+LhY
0BpA7IzLJYtTi3NS5OUwptaYnoa5diPiWfv59FiUWdBQum/+7KjDCr6T4X9S
rFR/3rJ1xJ4pEu+Bocn06B8lFM/wh5D6l+XTdK7EIpcZBdE3WJDumWGncsUx
qHAWsiTLbBFVB3PaJiR8w6pgByZa6HiETrXN79/BzIIfTaKmq59vYaIw+iQs
vsyhnmXJOImduO3sYK/UqOVCNbR7tQe10KSgRNutRwir3BjNJCdC0CaZy8n2
3uyj9L9Fz2UdY+98f8e9fMcNwSkUrz7SWntWIfoWOPqyeaOp+/PBgzu3f3Qg
kzN6gg8mUUHGNoGRvUDSchRIO/rEo8FhdQKid2EZQ5VACp5YYN6Ntsa0lp1i
aEuHz/wjEWvaekzGHxNvl8hRexMsSIiXLoFd2nkNO0VHFq7NR0JuaTUo+YT0
LlvPbpW95AE5yU+9hKPMaKeIP+6mGNoyPmOlqkOXKmeUR4dVCYfzCWDEWxX0
63cT0D1X4V7+ZmJejx8TsfUUOedQYWMP+Drokk4y2uIMi4jio/WYZDdCfAZ3
nz6ZH9XmOvhmM68Fo8osqvQJ7bbWm+Y4R5exB9U5HVukXXU5r7f3hNVhEtoS
CpT9xxxr/cQjHQ23mJ6x1tJ/rsf5LXKacHMC/IfKQvW3f9VL+3fwvAyGjnKv
/uAeOL8MuN7imAb9nxf+YHAr0R8tc0pZS1x9YQUUUf8/FOiUuIGgL9ToKukl
HWH/k8cX1Krz4mPYtM4EzF5rT5aAP2zElDUNX4aUMIe/4xhkLu5iHx5d/VHo
W5l2Df2JHECoRyQydJRCgUbMmUElqSjJVmxy3wFDndTcPWxNgiRo+GQJGTSb
u/Lg0TUo1CAbhDtCmPQvA6093UGvu1Tr8J5ZOfWbmpNsjrkfaJz92ijUei26
Pt4kf4sD7RJXKnK1a/tD0CweZ4jTGNNdA5zVp4U7/1BEAzEytti719+MjDEW
ii4z6QQ40EauzcSETv2ilxNMO9jQ7G2MbW1jaHOITlxOeudzZ/5rhgUeGDaH
BXqRcTVxxF2n8RNylpFI0B0OEQoH61zc82Cyq0DFA7yfRf34hLPpV7KRL57i
mef8egOS+uZ7z2yOZFrxVhiMe6/WnOkTU4zE2/IZRKnYoG3ADLAohrtrJGkP
We4YHwnZ43aetU3/uFrJSdF/78mjVSEloeGUiFSoNJYxBPVzcenZGUBw4q2u
+F6Jfn5lAPVvfK9quxQE7PtP3HcPAkaAycOM4fAz1jiEn7uEQqKrbh4N4TuC
72/jc0wOqUYoZ2XeJVS/fydES4HwMtH6hxYiKVWTlNwFKG+tvH9DLc8RB6JV
5zL5L2i3Wk+2v3xeOOnolinrP010L5CNaHU6tFzL7T0Q3QiZceryoSkhraE1
cVrQM6JureqOQ8R6pcUL0Sq2w9WeGoCohNNjrWOdUOAApQASO0o6+P/gHRmo
tCGchJWhImQd69Bt0I3oLt3eUwTv3EyliwvQ9saZTQJi8UmTWXlzZmSEkbmi
8iOa4Hu40ThDv1+uGmM32HBDNdgKbaKIX4UjVWy4nVpyH0jbVLQyQ4HuCZg9
2XlwjeBjvKlz+vyjlizlr2jihAXWJp1DGksPWQ88ChgOSycfZsj73QPamsbM
5oR3sYPXlJLcKJbvcdjXzsBOJi5uFwXzimsM5TynjmrK0Cy6j0g2+cZGnNWT
AsT4149Q8mcGlVCMZPWwjpCOoqtsyB7rcqZ6Fo3gLKA1yfKdYjg/rY4S6a+z
aaDs3U/vwKRpe6glLTU3s3AvrFMW+qIGPDlvVb2Xpwzq4EtJScgITL+o66gJ
Bxc1OeavnU8g2mM5mSsac7g7Z2Y7jPGB62viH8TT2nmiB6FLQ3jZpqm136ix
EEXS92A26Z0VQ+2jItj6xeWVXqJmla8mLOEzoLP5AA/3cPkx0MWe6svCptYq
EA7jDOi+z0KtxqTS+zzLBpTHW4tcRjU64dcp6i4z3m1PFkWK1Sjh81U0MwVW
zoKM5HnmPe8dwuZuInYXETEeamZj91DRDixAZhZ6r28eJ5wlh5DCkb83F42P
mlq3SYCnfAGQSB9lTAGvP18lZdEzNpiy3rbyocoajrSCPxVRiNgd7vpMWKGP
o9blxiD9uVAEpgK3spvGQRQrumpbDc7LUZqeUppEjEJsIsFKGQXVxTYh5z8D
W2pgbvfHlP3JUfCL9v1AuWdW+HCAWuw2zV+dCXqpf5sJ9DvJHYZXkbS1i6TD
nuZ5D9iEF+I9//bKIleIeXBS5PraJaQbWWKDgE/T7RdGnbuwqJ9w7GyqOFyR
AEg0+ADqVjLjku4IN3hGvVivG9C0Yq943yfcZN3ruCpX6yqqoWpU44RrS44t
/8bHM5PUV/HeXSV2T1axJbnaNFxPeE/8nFfOONdGKEK383FXcio+UiZc7iNV
9HOTA2uP1Ls8kGPSNl3GWEsXWeh7k56RpFtUhuN91Ar+6FqFrzN0KWZsSeW4
gDH07DdX8FMkV7KSSL2d35106oLC9BoZwAF7FAfI6nOC+uETk2YADYNMGWv4
TNV09FY94fRchOBqOyOmNTw3a2VWTRhC98BexIUHfzkbHBk6AA5kokhwroSH
Z+N7pJcbozkt+Hvt+KiXV4cQFlo89H+wSCQhbIjcbpacr/cdrFvoIiF+P0ap
aChxdoCGe7m7IrHjtO3R5+EBhM/iqgfBsk1DobjD/LSBIVdjM/2KK0ZPDbjd
ksVzGAEb5JsVdAHfxenelwxrgsFhQUaFfJ8z+aE+hURIzbrIyi7kA226zqTZ
VCSO0SEYNuHmX87Uht/OObbmj9ajl52pV+2RnHc4yvtbpvsIogMRIpfDC+/C
Tb4XRKb0xJVpWRPmvGttPV2FRUeuVdc/8qy7sfgXxNifLHXIc5+sopmjudgO
WImyCdJVLE/Nb1zmjVVL8BaRVANi48afgp+NpqeKNxfglyMUJzlcA+2JkXmR
kUWXxYV2SGexkV4dql1SfiUMBQBgVj1w743NVDe//LrMXPipvs5VpdXGldkV
lIdZcYiad0C2bcyhvpprzElbFv0SGHlHbKafejr+SiWf300FaYzDomsljcD5
gZN19or4fu1uPRFY1tl4EULFP0b0oDDJjehqXWdoKzYl5WmqyFSsxhBspwTA
xYeAkF6mzDhfCN7grb7DjS8bUfZV9PIKe3hhu4x8ow7nwR4MEqwqQHwcuYyv
80zLdv8hVKfBJyu9SiGzEG9fyNgWr0kA1iJJ7IB8vxAUWRQAWNk/2Jn9lK5W
irdcE64SbZARk3SbS5JFWfnNFOmssnX/n4Zt4rUsMG8L1YjP9mofdlwtOF/7
opmOtYsVge1KcoSp3KUfd9W3CqrkPeZ32ksK5ns1RU/O3B8F0eu+utvtssyl
Ld5x7XDEdYKp/cADGn53hGx0YUakR7KP1qyNEmYT1R5jwWcUMmIes3enMobI
PXUOhEla4hq4HGsyRkZJwI3NmOiHJ5uNqPJw3lnI904VErtUCXMN1MUw8EYu
0yZSqYHygW534BbJywC8c9ADJ8lrptFt3QHwn/fksqB5/AzvAPJXUFM9bV+F
38ZbSfvlV2zw5DjUHsDN5zjx+vMKBGjv8i1Dy1jiP6bicNSEj2Ab46nqbLDq
NZmGxUjiDIAInqTGmu/0oC1mmkpKnwB8IYRa/phUUEcjmVmWU6GrOqnva0N5
U8SZdwMMBLhHWnsD8rhQKSlUGRD94fiW+/WF2FHC7jMITfFGYXXqK2AkV8II
Cd5ghW5ZC8oaKvYHy11pAhhEM9pKc11cNDpF+Y8GjZfa6He4R8Doci66DuT6
BdcS3cOLa+Czk4uxMabmqVYaMBPcZpmn188kG5vWQU7aO9uUmxthYv6hCb0Z
lrsKgekko9zAXRgxdvZL6c0d56Ykejd3gPRVmiGON8U1m6kHHhXxGkCz5qk4
Y2HsMEwZg6AWj42jTcRuzj0gyafgawpiqaY38N9qZr+f6RZDVyh3NeKR/7Dk
k0Y8hzQOYDj94tPlB3GmFkZ9qVhsaPDr6BEAjA/90oWHqEQxKbBOIxKfe6WM
8ydUaKjryCBWA+4SZMlBzt62ErMaF3jrznM/CNJGWkO4wMxVrd6lxx+hPocC
BBCq5sJ0F2sVTaTqPEt+6tDAho5uTVwjz0FJ4ame5TSF/+qRa4EXdAA77Xjy
vBee8xljPemPAn+ACVB1ykqmkFW3SXKz/OeQYFyl2IAsKBzpbCHMqqNMRyS5
h5wpLPNEFw628lXndp6zx3mGY6lQ6nxQS67UYkOYSc0VW1R1NDDUAA6XSPmN
c6N66hECkJIAUeiSNKw6TYC3nVzcJjmA8eAfT1nEr3n8rc0QZsSbcihAv34R
p+tQTu+LVEGoQaQUAgNCvENCUeJ2j8YiGNolOkOoQ9y6GOoeNhad77XU71T4
uV5LATYV9FwV7ybulSU9u7MCKsgO39InnOAugpPzcosr1A35K67C0I0iSo6Q
cwQgRN8ASfsxKIu2wpabqhDfjamBUU4NM927ex/xqkkPWw7ZCdIgiLV58laO
r4UWPiqBE38TJqznhNUMm4OnZYt260QHbiVY4AgLs4oBqXILmEhKzRmRd/v8
0gQmIEI9viIGBJVfDZnGkJLm42fq8wMlmG9bECU/0fB9RNO0bZ44pCHBzI3y
3wZMNibDBzmmoIe7vwP17i9SlC99gkL5SMffIpZkvIhyavLdPME7VJlXIFeP
QOc3oawxduiM85khb9O9EiGnyqOSHAyJZkJqZDUaP6k1gN78dpvpue5VF+3e
oHKOGApFLX53XubxzzfrqGcKpLA6AWH48JVHmTYZHfPkcFjnTMvvpodImzaf
zxMFigzzs5IWpfwm6ZoVEljv5tDamsIhys7CU4vTVkvm1ErB8TOS6+nMM3i9
5V21s8vpianpUHQTHrQbrR0IYXkgLmpLJQ04x6YcmKsVz4UQ9BGlSmetAj0Q
7y7JM9rCQYH3AmNHGZy9nwbqOgs8b+4Wd5MhOQIVlZs4NUSknDjV32M4U3OP
VYcDv60ZXIrui7ZMp+bttFADTzc8/4WdDEcANf/ZNr0hyBRb9QCPz8n9ythb
gGYdGenadDTVSbEPVXEYOTfh8YLq5SiVQmL0WaAhXWdEHWB+GVA/OkW3Cbi+
FeQSgB9P/IHbTsNQh6LW7J+8HcE1CDWciy+8rrxPnov2oJDLVnqYAh6pCBPf
vd9SCG7I7GTo/kcNyYNf2kLpK75VGm9BTvUtGNxizUSzN9BZncTtHqTTtyIC
qQW5EOon04qolgDnvCtsZUyYnjvTPLkPtL9VKH2IzmrcmPyHDF/QFAXZxnuZ
ilYgph9ySKyr27bJNtw5I8kr3UeeAydyxV3kwpueuPDoamRvgg5hatXFvcFZ
xO9+mOJgLmyUUIhso8tk7roSZd4zeZRr51IOS9Y9KAfxkdOsu+RZXW3vCzpB
nnqbiyfgR8v4PaDvmtGDJ0HoCOtI/Fbo+f6pQShUXa6iXbzrvCGkN3fX9sst
s20XjJauPmIQG743I4vXjKO0LXIhELGtNc3XAktfnBSA4KEyslvJEWAyQUSr
jXv7hXalwElNoynRaHyL0PjNYYyWqR888+VykZ5zEDbVtSTPEPnZUZKoAxa6
24zfYzYhSGvpPW0idRj9TKNE6UqyE3NOjQ+g4sM8CAcufTkovLt27yWSkG0Z
49mK05IG8Re1XEmReGzuI0n3EqMDufz32Dkag6PXyl7YNGo7AP3/FHfBmUeC
6S8bf31oYIIp710tgGkSoGlw2KsooZ13iC+Pn60uaG3Y4ENRKJMEjngvXvOb
ePpLTRoxyraLwdwq5d+zrkCUWw+pspHlM0SnJV0Rngo8HB0vAlNDzqqY+VUK
dn+kMQF8AbJFIxSeydV88S+FiKGcVYZdxJG+KyeNwAcVnO0s1MqHVKb3Aa9v
ihqL5nMrQ9x+gij5MDwBlrPwYhsvI04CGKeGW4qXApm4Ar1erbvJagb99cUr
ehpX8GfIIPjCckyvzENJ7YLslChVOkFZrtWLfQXk8ofzrihjWNlcctavkZbd
jdzfU+dTktdR5M2tOGT1zuVSBUc2aOg5JUMfV/qTFIAMp0tPHzPCX8opZIAO
yBNggw9hho8H6ZUmf60p66muMgxKWD1fzBuGQI7h2bpnFXoFfIjdzOnXh9WE
Gq0eJCooj33qtsIXMpm+ID4Z6EGDNOwdTLf4uDnLxcpJW9yIrfpH/zsuQqEv
Pt2rLWzA+UOe/bRi+cvs4zjfN76qd27ycld0ppG2t9/bI2J/kHIPscNHbP/T
Jv44N54g6UU9XU6/yW3cq1YU/DEALYaR5tD2EAZJBQPwlQtEUsKlyE7AJ2In
aR1pyqO4WnjqVUYBqGV+PP6bVfLBojALwxc12m89HjvZM0F+VI2wkxsgB2Qs
1sD2dpGaKgtjWR4lwywGdHn4f7gcXU9i4mLAX6sIXDOygqW5WMMWqIZSGDj1
jCW/Bb4rbWMR+UD9crpdtLIvIodEbhzDWuRHFQZbXu8ldenN3w3C5CWgM1b4
aWjzNloCTheHt0CR6PD44lGlsdWaqSVVqSK+S7/SKc/1ekGaiLXqxj2keHza
UZBn6IBllf0AANoaptdHhhM02ny1ObOFnMsvDDd18Mt56A2WrK9Ufkk+gv6f
xaWMBDrezJKy7UZaQN/V/yzVmQ2grLc6k+Nk1ZVVCt0lYWu1UkLJJvdqaRBn
XOEGOLs7RtTlDYyj5yUCF91T+7o/B7/+OnCYl2cpYb7/wfLB2S6lhHxaJjp6
pyOx8T3I8RzhCIEYIV1tlsbSSc8x4EMEWIT0jmJ1JoHZXxy+yTJTfqBzK2uQ
Mp4DsCCHQ9xIuGXM+6XNDGIGCZ9BTD15RAkhwramIP3EJ2zwdi1SpkDBfKR6
eLH/tdrk+dRyI29sUeg81GVHhjF8N3lqZF0Cv2X3qxU3N4+wlTR/pmU3WMPD
nIDbbGT4HyYQPxWfbl7sz95+rTlI/EIdJ4IxGjLfhP6WLrvNQry/eelJ4Rnw
JKI288QxbdCsH6VWwJu5/8hWTpQ6gp0uLDfY7+wuxAQ52Q7xfXiZA+A6sDFD
nXadwJzyoSJPrJ3NDGVibMZcqZBh/YRYkppelrhUrhFJ+bNt6PqBih/yJTfH
4cw5tlsOKF2JLvj8BNkMP17uYGU8Bswq5k0JgB4VENu+xVZer+39Q26+RdqR
kRTelubuoAqGW48jmVP56fF3s7A3QpVoqYVaMTxU7JVruhvEQTwDmExso5yu
KLsK51948Qfuj7JXWxv2aGyFfHAPxZxUhA93dXi71i31JeICasFS5EpieJEi
o2lOYlTCe0jt8nnyH6Xo1XzUvjcXqmkV419WzkGFoI4n7Ahnicmo5ejpTE4G
ZfqLLKmkCPbrmraYXISaEuA89yZ4GCoXfWfdgWOJEV9UO4h2Ot1M6SjpHXFe
cNwjekyB+1M62JWetoJJZnYr0OsJY6N1koE000Ud5ESQ79COLfPzmnhPzSGF
POFREuB0YmNqFzA80XR8Q5F12DBpg7q3CkRD1d7IRuU6PG4jv730wWzARx6D
v7QYKqewXIQfUHDbur4UnC9XubSfkoP/nekTEHRdFF5U+X058pvHovjElQ5b
MxVj8mNE0UCrjD5xDEUoODcEbdhW1+N87EmN7AM1Vf7DegqPg7Xom3zdGQm3
DVtWdCitaHWdD0c5SQaQiN+WMYhqo5l6X+OtcZG84+o7qAy+dkXfbotOSVcY
xZ+SLx57/NpgJHUB2eZWCE3G2u3wQVPOqU5AlC4irwYUviWn1axlx9JlavtF
4cIz+Q6BcgNRSnHt5hsff2KOmC1m7JMplX2kWBK+JrAFPBeI0tWIu89C6csL
bhoXzEtsIAEuNFOkDc5WLuArRWtlWU20fAYThxv25tWHuP2PZW7eMixxw7Pt
PRDP0aew9js/1c/Rdd9XeR4PMDkXJd9O8WPw7LndJl6Sft6AEPGRJz71pDg0
S30JOzcDwrL8PJamYDiX5zFaiII5b3dtUJg2nva5BCYASo2n/UPGzMhZDYCV
EZwAAACswoQki6/7fW5BfcJrNgBxQoDdgo91LzjrzPDsG6ODMohEP18PwM81
pxAFWN803noTuEntYI+jSqFYyWhx6Zoo5QXykNYwVinQRaUgyYpqQrvizcKr
wZ8Qc2wJx/2ANFuFZTSvFNiMMr9bWeVjD2knuPJz13ZEi4Lcq5rEM4Is1zrc
OeIV9q5pdoWV83TKOEIGq9ub2F5OoQmQMte9Rw+Hs0GqrDo8ttSMowSnJZdo
QioPbXX1MzJNqfoFvsOoKU2g5SKSZtkcPRv+dG237NJRtWuRPN7MG3BIEXhT
k7XossEwR8xoWarIsnyRSulMisbb9uhc6ALxBGWwywamjbZy9dFPjxL2MLk9
c3DBvy5+AbpbCVyQR3ybLyKdCQwkfuZkHl5R/qe3CQUyEcMKvgArbFw46Z+B
hiU1QqSONZ8PHMHoTcxie0eU7v2WvBdak3U3Mvv/3bOugL6M97VHhMWqDMHI
5rv40S8IfIKzBEN5f3106nEKs6peu0jXs+ZIbDoL0meyLEOxwBfYJ0bNKOPb
k25wnlybsc+pieHfCzXtgFE4R7BeIgz+kxv24n2AopWsKbn7ZqfnXTKoN6O3
AF85hSxlYr4gsVdjWYnSxiSPGE8rbcK7T3xY2kHT8R7ZpWrBS4J95jih7yJR
2+5hFRjvlCrFGABuE8WNrbcnXXzIZBBYuX738k2dbu8QsNIpfLe64MSda3VP
tTzB/OJepYEeFxzopkBRqVJTCq7XkGRT5ZEYrqsstSPx9TwoxIIqwbs2lHjy
0AHN1n07SmVbBmIY8tV7vmjSWMCYFz7zdbB0IP989u4MqjAUWftVSD05Wfen
2L2BJKxv9z+XyuBsCHh2bNHZ/a6WG29N/1naUGql8fOuKI6jByLvtncTFY2M
5AJ3e+26XHDY5hOMxtTj3SCeLm5KcNCtxyccUahk6m6I8ooeNEpp8CmGM61a
2MFbCfFjwRGiI8KX6l+rQf77wEZo8e1awgjQgStdAHHRpN7+vpY8HLcqUv6F
DD4xnahOMO8aZNSQuWltVXmWghk5zjYP2P8psTTDY8DXS3C1ORmQsmvnY9U8
5P7KhQk/eDNHI2VvY4TI+Xx6oZdWyC5ZTpiLaY97wMFedNhFuE81iEO5a7sp
9pqSC/6tiAdKQZTNq0Pbs4bayq8jIegE+2H8PKmMuPkxqHMC5PrgaBvOTuZs
+inNPKkjHLAHKc9WJagJ0WCntnoRu08zKCXHh2e9cEk+67EyIE+JdyjzbiA/
cLdfYa23exrEpEd+Xkk1zyTBXGLwOuAvPa99sAPLhhC9qvwMMSBHjNgmXmay
DLJGL7sZ2x6EyfdS346y737cIHIrxgYng6RwZ7bgQHxQdTWsmxPjcroa4zsa
Zjbh/mrfvYuu+bh7KmDKGieOfnTJ3zh90pyS4UrWHyriMcfIEgcYRCZ0abTS
+8XOkAJZuOIfOOfxel1GJgNav6qMoUB75rveCKmLRl1IIdUdgwGgcemMh9DN
S7Sl8hvf+u/dnKejY15A8zyzWIpkOtyf5FKG1OoByC0NDckWaO6ntyU5Vvub
2+zz8CUcBiY6advkfwrwspZPf12F40deJywsD035lHw5EWZgQrTwIDO+rvk3
s09b+868eVi8Ozzcr+c4iekzL+Fp39B0NFwMqlGy7mGo+cpdQx9IDXP4d/SP
Xb/7jAdawMMvKPZ9t2zMGvDNcfm5gW9/Rt6U8iYG7K9ynKaK8aAtV8djVJMW
9qAbn2J5zBiAVh+w0jQFbnLncSgkLVPdrUyM6OePM37EN5U/bXBCR/QF0vTC
ROUWtm1NAprdHsG6fqBL2GsFcSgIygT0ZK9hqIaPLda6EHJprPafF9RS5nOp
B2X/G4iXeLXwE5v8o7DLo5q+sz54C7YURVtIw8dT+l8peDl5gX0ZqNQQmXxQ
uxAgYvxwn+3k21Gb2qR6D6kE/w6A8iLfi0A94mG5h9O+kvND98KIfWSB57Gc
EKXOB/Bn1o7Pr3JQrZvGY74UEoYPc0mSP4m2A8+34DjdOtep1dTkRubGsryh
t50fgXTIvGCGNm0UW64IvZK5kaM6++D3dg86YRJ1i/Z3eBQL6QPYbZSv75pl
uD4B2bq95ltwpxleUBQkryC3VIIAejBeIgBa203jIfQLcvQmj7Ho1v0tNsbn
S0VgfomKascJTmoHGsqIieap3XJpdoH8HyAuBAjI62Pmoz9+9mHOlT3ebeqa
59jHXUf4Nn5EE5/z1AU2F+enhdGW2Sy+f0EspJ9bqV9wiUGwgZFZzd/1S4Zo
4UhdmkSqsQMDWa+w6EoKBcH7QxBvSXhhVffrJEJTvFxkvgqfIOzgx8FsWe8u
DwyFfxETjbETLAvpZLXlgWXrRaGJr8DtvJyyBJF2wBSmrFtbcatcJuQmB37N
uwxyUSntTOldKTBNCorWVXn/jKcczzss0VjNL4DbBMzmKK7oK4fW43NsiCGF
p+uAf6HrorJJT2yOa1eqk1sqoDj4MCdNpIHZVpDxQ4YvZ14iKOwSgzNKdMqN
opY+50tTmqzbbw8d/FnluNdSIpdvBsX38n8vsmrm7O2Hi6McQ6Aki5N83Ayh
Eiam1AaSYYDUlRm7ZCDsShPEXPWWCQ/U8G/ieidNjPYiYl4z7CLMfVv7TezS
8/9FxKKZWlsqHDDA2qXKrMBZ3qYEfU/tgPbIuVu8qP0fX4dOgpmfb0mubh+C
apcf7aXkMz7haOfaM0Zs4d3WKAmmN35yHgo/4XOnMIvOsNh8FSjKwW6HLvky
9TqfpJdT4Rp4AV2Vd9s38WdpbbMt2PN/E5LyaNBzYsu/aoKLu+U0SWBQ3GMq
gZMgsGb2+oeThVPXuON+qJm7UcbTBdCfGMEAW0lj5sOs1djkG6rAsLcanCZp
9TfSMuCA7zUu2mk3tovP5h755EeZtSIgsJeGpYEef0N/G66Hz9i603XcvoAF
xPJqXI5bit/L4k3vDnw1PR7nnzpuJgdW8NoZADMx6cs2ckDsyLQCijm+5R+i
6pHJPgx4wTSQnqiFarcG8Jspkadapk1m0V9oq6rLXJxNrdWG/S2krZWgI6Kr
vi1Nr5nI+eUy/cy5lo98QEFgla9xwPRDbGwHHDO03i4jMEWISwsINY/JXXtD
T067MOFApC7YnRB8O4xm+mGazbFUnHhsvSGlg+XFMo0pG1MxZjxr7yiqJdVc
nHO7qSIBLQTmiBi3+1m1SDYr7lv0XkRURpw4yABzvWwSFAzyqV114ihm2Bdg
aHtYPs4XrfNIN6nWOzp9cVHsAdQqMMwdY/cg4N2cZoSXopDgiQF+cH7vB4Pm
KuSdlwnrttCtRqQvFSm9s4KG+wMTvGdTwG/oyPxdEa9wAU3VTBt9TgaFWgQr
sb/eE2QiHK+yFNDAbVl2+QsHiWSkB9q6brXET+dP9DSov81bkV5NX3x/0etf
jFJjMiDMUMttkZtoFQ3wBIPp1pKCs9cyVxI3vbZJ6Qw9VN9sz7ibnroXkV6t
f31s4WlOlR9b+zB2HijRi5AH/uoCoIhhD4+5mHEBUSS+E8tqGWC3UzOC5COK
/lEudfVGRzYy/v6ZYA2EWdHO4fQveBjcUfQggRgnpOEezf5y0q/f1eURhf3c
CuBucbNPx+e3qSyl3U/jlAhvoya+fFWki0VBOqmzA4QAYkb7j2vonBNRfKGJ
6JvRt8Cx5Y7f+rk0w8wLdTRwuOggxAJZJZ9VUcGYDtKOKsrIcHdDRMbiEsx/
LtAzW8O865Yj/ptMrzYFw0j1Aq7kv1HQoKOCvjMjzbLWeGXS4Wc+R/3bImE1
4T9CHLISBMTbTXUv0XnSTK6+rsgNRJ6Ua+ziuHHpADB8Wh48qkZz8khxjGWt
T4McAYF/yuqW58JR2CFbk/K6/cWrG2EsL5EKX6t0iglcPQFXXydB/ggGFliC
uCqokT0I3HBURMVGZkxl+LX3Ei31UWAup1RmP/NwLkKgDkMD88pucunIWGPD
g6IXr3b00WfBFkVWX6Voycg/RmJeYMiTLZ0piPLrQXbyoL4JteDj6QzuC5km
BQ91KksEUtiJcBU2i98xNbsUxyheQcIBX+CBkMopQj7wD/PxvNy2o9qxfHGm
PQW1PPghBarEz0wFr+RvXdQWvYdAewGBg+glXLzGA2nXA7Hq02w8bWuwi/Qo
YpDWaZ65EAqiQIWKh2YYYaQaYsSvAvnN1nXm453fN5Li9QgaOLbSEs9zqkeG
RD57m4zs5qz5ItOLwZImb2bBf02p1WM5WksTtbEXBaimOVhinXpkxq/dOaw9
a7VbfCRY+svONlimW6++fEoBKME5YFPexBqeTJZqdboW7hSOKanWhQo6fTXQ
AI/7jMnPJJ95Vcqej6sXfxVpICrKTXd5IybWjYiCtkADczq0+b79vZ0gfjAQ
FwEs1P22MLuFB/OvplcyI/ippg2WPuskkY36k59DhbabilwL+BEkpXQ3NpEt
aUUhiVDsa/LOXBz2i+rWNwpqLE8vc2ZIRxHjoP2/1Zc7hFMAgx3nBOvInQmD
+xPwXEJxj1OHwnOfibNUGF0HlkU0UjzdSYZfnMZ4NNAw0sy804kUq/dwwyMh
M+e1FUiSXlWx0FSW8UtF9EqAM2Ew25Rl2oopdwaUmOSQaF09oVgKBsfA5+aD
bEbLMji4R9IUdPoF2eEe/fmnuiYH7W0iwBFSG9fGiK+jVa+O66y3/mdiU2jK
qnbCSlkADPOfP/Rok6wKgxDfPXsH1Qpdq3ByDzS+RuXNu6fNGSkuxFB6ZtsX
C2cdP+d4/7IogWuARxPyEoh9MYgUMWBmCjKs/yZZgEVD0+8GQdSFg0XPYujy
+DNc0bkNPFK8MlRsFAEmmOWYnGQ9ZRxNeRnMKNlBtY3kRsfW1LVoBL/ZvDkn
7KvG0tfNkJnqvoRUIMibNqU3iaNxCddgSd6fyOIdtJB/1vEpefwah6iFI1mp
wy1OVd+61WcBhTAB/SY87HDhNbI8htNYHu3/cGLlO+uwNtZTdMtygcbKUY9B
v6LstSYKqSWgt5PD2LuyRau1Df6azjwr++vaJj/AanlJbe76w5HjFtLqznQB
7qDvKY27GQqa/EB0szdF1U9X+5/G8dsFVdbfrCL6bkijom9JYVrFwAP51JHl
iYycvvOeomjqnFs5tG5gA8diXOkNei2lC0CNuK6Dn+pCJlDiCb8evwpZh8QW
2bvirS7J9TGC8Lohkftzdw+tRkuNNwOoq19ZltX0TxGYLypnoZNspvBVdNXV
TlRIzdkY3AcFdZhtyUonL/wS74YksRxlrZG/SuLi+EOFrwzOqc2UIBbaI23S
VdZSJ+pafAkAwxLhaHkrtlwp3PZXSJASYuQJnLv+NH1JR57BPn8+1cDQzGCe
BYf3LuSAfBUPrU77KTSJtb0cla3+SyFMjPliAa1qqGJU7rseDglESByNqT+1
3tguLRAaQ/Q0h20cwe7MR9JzfLfIngc6TkRrTwp3DRty8DnRf3i7tuNSn6vN
60dNEn1J9xNTpfxY8rhirETDuHuhp2KZMPcckZMJt1/tfWSaYl9UgaQuT1GJ
4hg+KUkoQ4xEWOYW7S2VPVK3iBNf03mCWT8J2IK/VYTe11zb/AbFmaM5r3nX
+D1Dq8+5svFX4VtdssfBKK5YWJaZLQvvIAWIGRt33eTe+fSAsmUD3Gm3LSYa
67x/JmTJi6gWunzRtQS+8bEbb2zHFwBNBMQCfab43dI1UUOs/p1AP7W/cF5t
BJNBQWgPy9qWybiHa1ppUxEtZUNv+Z2u9c07i9+2Lw9PZPGvm1kZqgIvlDjk
qMG8nSU7ObPbkYZj+DG5YG+uLERHXRRtKI+veIeRiWArbsN4xlsw49QP3fc+
J7rsREfCzZyNB57yyxFuhBHiBSkScfHeQBczSMA0kHoMOsYIhjDJ4fXt1Fg+
DEE/CVq8kBeL9uvoJ2uMI0t1TgmJcwSlpV3PWgp+rxPI6ZJ8r9Tu+8JPk8fY
gDsOlHZ/h8mbeyUsMv9tMTykIKphAgxpc+nO4HecG7avyqBtoeUnHQcN0I7I
6+hNJSKy65MX1wf01LBpI3YXBF1P8BTDb3NwUS5IOxHMi2qRdAmsDYLY4VuO
GXIi1yIxMk5s+fsMSqVJ4HTCP1YdnLS6CrMB+3h9qhXWwE359iBypsYS8Cok
Uc3TQy9JHptS6dx5B4mddV/vct3f8CWfwZdHcPv8zESrrGqu/JHxEriIKm9v
FsWajsZ7zX2R+rCAa0aBbRae0/VeM7t00tyvbKv8Q2Xfuh30k0NxlZb3mx0p
d9vGr6YcO/gcAWjIzBLAmbYjtFHSlBGRmvMLvZ5SqLHtrXFkoc8Uy3H48WHU
i5bcySi4Z7JZbPlQS6TEgC0VTkcYjRD+ylPqwzrJdsLqpKdZfbrt2AH+BnCD
TngHop1hIO+NrgCb9Bug4lHWuRfQXT5c8Z424D4oWo8SbrDnrGuD+Zz5AS6N
scDhWtZjQrlSdhLHGn7ydCgw+ogvQe2uaome5ip1BFE0cVns6gftqg40Hob5
nx+E4WETLVTjY25UqBMsc2Y2XvXMYwirN440nVKrRIgHHhBewVl2fJvBkJvR
jVUdoiTK7BTYpATG7PDu7fZVF85uCwboxLs3UGzecrLZLB2Sc72bCrQKVi8A
cV03429VahUxTFhGNaZtEDe4E/rvjzBx3GH1ntNeFgnNHMncQjUzmm1BCWA3
J1tLM4KT9YB4fKbFAzpTiJWO3KiB2N0b/Ia8GZcvyd7xYqlfoNkRAsFqnwUU
XYKVYoOESCcjcrIFlbzDs/vshK9b4OoujUuMqkqq/6OrbFdB5dSLMMcbVKVm
+7UUdvKINfn9JOMMo7tU7CK2ePXR1LNv4GHgAxg4QcUEQ1xHgaoyUG3rdx4e
xOHpmXZDgk59JZ12YlRdXeLlLX8fhXxbSUeIYK1tOVT4xRiJOJ1Tgc7snf4z

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiKycLouMcEe7pHd1uY3zQwEysFHdUDs1B29W/e2TnKezpQZb8JHgtnE2lQCSgIa3jnLNaESq5U2QepV3hiZETDBITPdQlH0BzcCdpypBUnG2PxkolGJzhQsshnAmv/GlREQeElr0ZwQsFb1X1lGhKqKurz0UL47vDjGJOEivhw7DJYVyA3WS+Vjs/M4xXxUQOX/vCDpiKPbQq/t/7W01xA7UueRr3d0M723pqNBc/3cyL5GMyXML2oFUWJYm5cRyTrD1oogbuLPapeKrE/zTBinBE9gG3091ZJ/9K2VdZCgcBt3PiC1KhUOgYY/LvGmpY0OETmNQ3m0bmLIUguCmb6sahWLWQBVsqx2AhnkjELD5AV/WL1Tmx3voqQgfgPgxD7wnDx/pgUiCyAxQ/jp+uwiwwlevDg9m6DCcqc578GTNyryAOokYvba65/GvEa/2Y7fWSPngcrx+ooQSFWUYyZ6mLFY5IUeIIlxLYpMBXqZ/JFXvA1GUQpZMvbJlckSo+mdc2D5jofv83CZvLZoQ1dRWG/3ZfP4IBq129AT7hubjYPSzG/z7HwSjJ3SWUk8U91dWFwNwyA4NeYNs/KbAVYaxhxFxbkbyKNSPoc9HKN0ROVd8uYh54OqvVMX3XBQZrGGD0DgLt2WrfbQVg8d4+5e2F71W7+5ALinVBFWRjwryHIYWtDwPx10Vaty8jlonyykOczFFyvYqhQ8KL8hIRgRR09GB63aedD5mg8IX+hJ2jDly5GNKrKhIkiJJqu5sS0oBWDKq6aDwCIqaIvTCz5"
`endif