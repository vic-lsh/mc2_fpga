// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OXoV3naBWN913z2AKAYNwxN5JTUYkjUL9vEYXJ0M9K9YvT9vP3jZIPIcAULJ
V2gawvDJSC+cSWd/tTaf36LHF/M74ufwCqKPGfMu3SqnnupnPE8+eJFwzImK
tCsGP1SXaaHHsFklExpXm9tXpYGDnqON6CYsIIKhyzMBC42R4MIJuNync5eY
aePbZN96zjT6pAVfd9rW8moUIovQPUeG9NqD8egTuyjDeI3ICh9eWToYI03S
nN/eBsM8QKmYeiGRFwuy7CzVSgtt3vBQ1R988Rs9OfeScBoDGOqaju2ZdMih
k2Zz5fSEj+B2iEbI7ais/8fwOr+jFwvqeJuPwD8oTw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N/wSx3Dxa09Oz7z9asVuTzGnoLFRJmxPZVym/u4nX4CAlOip23g7T7MBv8JG
j0kWl18gOv5XXyJG8ZsWGnPC1y72oX+a553vtqHfQ0VM4Z0X2BuAQl+342hJ
aJqs2uL7RdV7BdUnbWkjDlZOGUVsqtjysSAnTcaZrx6yvto+evGi+EPpiVq5
nUExyyxwwpqPj9zc7KjvggljOEKUvD0rmAXWMxAJHiJRDIpWP+U5MUISYnsY
jZLaVppQjvjEeBqFHsgOI0ZNV2q3GpgBTUpL/VWjrdgSdpMZcOwLYfC/zyIy
aDslZTJaFGgkb4290MLN+XGy5X++b6MYmQe6mgb1fg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YxCuSukwG9vp0LIFGD6hnwBfOSqDpyXQb63S48yLdjEYRfG+fSSLEaROtSb7
snnafKpNYMd+hrg03pVukN65bbwkQzpHNnJe7WNVrFo1QKxkrraASX6bYH0z
i2BVpPyOzJZUNh2KxSYx9S8WagyVdMOitzR1KVK6Cl87GHSCcDCx9swvBRka
WivdPpJx+uSJD2ZYysFqDIrsZiJrsy+BVxDQUYZOAZncX7rhSMD5uKNjX/6M
8HtIamhcgZYeWu2rLZvzbAfnUY7CYGedUJ+UcOHVi+q2fcvIKpzYwZrr/Rnf
1N6QWpKGm/H6Uz8HiC9KK9gmAma1uX6nxrnfVaq3fg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WA8B5j7GAr5kGAcwfRPw5yd+2eWRZu+hVYuBKk2BQBBSRPewm5UxlJGuW2+2
XHw1mWa94UsxeZJCVSBnRn5dL6ZWE/sfmonQX/b61PJ2CX1hDN8YZiqiHMUO
TZYKa3GzqPijCoI6v865VSVxrPfOFF3DZV06gLkmjt+000CNKBRDWRhWhEo0
QLdKU/txhKdsVroXIlLLSevXZxGcBHvOnCjVJGrevFrJX9SKUqjY7DScfxzP
oWSI9saLJSyqWcfG+vbFadUQxlJ7ybZsAr7WoV1YWuRjRhyHKuVxOVlC+vxt
9gABzQZ5B7n/CN5id99sOwVYxC+wlY/ee+IKIqeUOw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YR7Nbhjw9R7cwQ3uf09uCbmx1WKbYyvSMFud/R/2o4WUCIN1C6OJWwYKtsZH
jbBKxWU4WrBJvO9ZXyje9slq6KVdbvtayNec399OBh+gAK+/XuiaYffo2tzh
02h8cpbXiiEB/oar5lFCElc9XQeJ5q/i71IUiSmf/XGshx4y9+k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rZXOUmzVdGqIcSndxL9KTya4F7df61NXmBewwr1UPER21MghoDF8G0j/Ptkn
9bc1gAq6CEglvtxvKAclnb6U4KIDwBoE992wf6QrKV33fpJi3IP/CllKg4E5
l4lXnOWDn5jabsdDH3PBL5QLjWWHok5jJ1ISRlMeHAuTlJPQqUnw77LIpLZQ
wZyE4QUUzlU7rNifgC9bDrXrh8mMbhTcvPf34aKqd8YiZZScJiDYOtRJLXqg
MkAhMdjDHzrTZBlr89trAUqD32ziLQ6d8uJNUZ9ONUh6UfSSxlCinCaokW3Q
ZVY5NonSMJU6gJ0DywFN15tAng8yNF3XL4D6CudkAo618rJEEOWwduGmgkxN
eALrH4JN+kdLEeKitwvUR2ZsED2jGAFv1CiCbqpBjz+ISDascQZxcv2oRb/K
+s8DQILVkWzRsG+cvu9IcJauc60IbnkYxIK9Rc92RJls0qiBuX2DjbMSh60g
VPfLraOEnmfcDEYapk+hKBIhh0nCol8f


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZRWcC6DtdTsG6+db/FXInORDgOf4OkO6jl10xNlenILqS5V5cKvZGAXw2N+6
vJUjT1gqTGXjNwYN+wOv9OAmkFtL5dptEn5BF44J8hPWFJ28UBP4cd38kFap
x0MgCbtNs5HFoEDGwwCROJVtbxA2GbTGZVz5cDrot/1oEjgvEjw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
StGxXUkaF7MQXwHDe7j6CEKuv4gL/69aJQ8KjOPk8lF4XMIVffhwCSa0hPpe
7B50C6PJaZntZRzV1Klod5hML1HKEB+jgZwdBujdrumUcpiSWRET0nyHMsJu
yd0AL9zwpW63bLmHWKmIs1LAWPJ267+77AFr8FFR4d/RuT+Q6JA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 281168)
`pragma protect data_block
ypQJ9S/xpFSrnbJdzDJHtqfbWiyTcb9bq/DznhCeZmQNptFsgai/qmlpIuM3
FlzW2iJYk61VxZJjrar5Hd4OnTK6K1PAe1XJDCSSZnJvcQb+DlXNmcTI98/x
cHWUQb1rGvvZjdq0AfW1q8umbAiaO2DB5xY0pQgBRZpXd5agbFq/KPIqrtBj
Ybfatg7xRAFUSnZ2tqpCSi2x5YygiFDLcEkjY3cB5f0bKLURs9h3O5/QKwRP
RKoetip7En00g0FLAcWsvyNIwXhoFZ5UtAgGoD2nkzbCWiOQQ4nnddH9HfVi
WVhNmzfTyZFldY4OB+i4y+t1Qoc62NK8tS7M3Knohr5OGl9BgU4i12hdByfx
xTLCKXEaAPJmMiTvUdchOkN0r9q5MkQzi2HGDdtoIm2xrxQ+9WCWB1j/5p6Z
viujDfveI9LNuP9c6n5SzsPHhCBoeciIfhQbulqc3WtRvc+3hzXg7VzXoO9e
ag4m9C0QbeKv3b608xT3OK9yHSKgfuKUKDOJCsDjGvPZkipGUVW5pcT589wy
CW7qIjHrDJSHMMEIDvimE6mNMMVEi/2q372TuTTvPY7porfJ+QFUP9q6E/q8
K5OJHmocXfiMJ4N6OSMcv2XlvEFqRi2QG/jEiQjnoP73WLIgFOLitBAU4HqW
Np6Azv2nBAAbHH45F5zrK/cc8p+SNhZTJ5k8RluCGKht5W+mc2F7umkxg4nr
jZlAADKyw9nVN9czKMsOlVGfa+6ihOJrAuZy0vbk5Pe+WaQ6ljsXV8Bp6VRh
XOglNFTH4e2wFxLDNZ9S+n5qX4rEhqRIaTnJt+b1RBAt6uE4h7f46KrnU9UH
oWwhQfvTQg0npYrjOVK3UlIAdiUylxd151f5zLbwrROvt4b0NJAEYsO6q73U
5Z9sN5qwhAzpzqOp6OVb8xaSIc+JBMV7MuZpN7NnwOnb7mVh0HpiYtBfFthp
Sq1cvEevNroXvn2j4lHttRNYUvg0KwQoxpHxBRZqa8MaXoXpmt86C2PCC4wJ
WsyHGX9x1nHu4s6rx0t3bQB6kYOqYhMlv40ZztfDRmzF5mhdONBI10Rc0aA3
5f4zMEhAIBlLDDyd1uc1ZSA6FHWZFbGJ+nCEcRfApA7FFBZRB0MzU6sR9/sd
UsxqitcCYx7Tje6aBaNSIUtPxMos89RYPbWxrt1aSabDWLnoV/VvJcqZy6xG
/n8EM0VuLDYy9Km83NsboEiQbaroe0UvGt5lFZkaU0Twp1umxFQ2kLJn5YzX
EqSeUdpuGjKy5ekxf6IcBMWniJtkdGwYWxdm2XKcMIVhd0wRGfKC0ucsPl/M
mzd3KIGZRge9eFEoO6TKccgh9ubnQTucP3Ug44zVW4wccAvN8TvmwcAw/N9U
zJ7ZLrIHiubRz+mhTIEcjVAURBOnE8vcEAudUvmOrWNefV/Yhz9fjZwZCcaw
VTZ/k2SwkSWvfG/lBVxGWIGguRscQrYSA7WEIQjmkt8Y+LlhYn049jaXbRMx
PSF1Os05y5Ne10ho+qad9hna4kxBxAxMDXl84D7ngJ1hc95OwO6UPN36URCM
kmHOH3HDM4IPXa1iLeUdAulca1mQQ+2ZUqEH+OFfgV5L1YB2BM8Eaqhv8P7S
kM3Tlr5m02k2UQi8ns2hQq+EjPHGKubk24+fZXCj2IjMoNfZ4zLec4IVLg0m
x9DWRUKausGH2pt/V0ApR9JIeWcbim2PAfghhFtQ0vOYQ7QXBMZ7vpC7ecZi
Pw3/bCwGIWr1CHMuzWywdH4Umf/KyTSGA0AesSzNqH7Oi7ABcJ6JnFMRUN7S
YPMrjxTJcez1cZbmNnLfPqCAfd4qOGYfy1GjwgOSGz0eoNgzTORG3umuZRdH
wRLve5IXzEcyenFVcKLffdHAeSp7mnOkiZlSZPmHJy5KevnOInDMGlUxNMl6
RSzoO0aQrOKRJlwszznaO0hYgrdLk8pKfy4E4sHp0QG3tD80tAQ9ltTZ4sjL
DNfUDeL66GmYBHjgf5s8joma+sDFXV6Yg/S4TQwlcqu/zP02WTj7eE3rUepI
+qYaZXTO5q/e/9pbawLuwnay8TmewaG+lTURQCDupq11C2KQKDhBg4+Vt6xT
k2Q2rz3ngSz9I6J+/U3l3CqaDGsTkEuQElQjQl0MBYd0nB6aMLzNs6TiNiCs
eQxFe5ClFFP56+xKY3cF4xGLGXQj7KX3q/y1ugyy6Ioj8WJUf4xaP2TevmCU
BrcuI8XhQUuaoRGX2lY7wf0QyuyTgkqpyQqWgrzPwkd93hxXCyuHuNvbJ6wh
TDmazWtT5Pbxn2LQ+pBbSHZkLs47MLLl8Jehofk5nW5iFIKwzYgnTrWnjDyf
gBD0vsWi4GdgcX/wGng3NOvOSgO89g60BXEpfrDwwgN/g8HYRTMNR/vmDXGF
BaeT2hOVEhmFE+GL28UlM4nJwcGj7Z7VOn7D5cCco5gRal834IRuKMQwvYKs
ZaSGlp2tzNMX8+vTIT9mT19zATzeA0Cu+xchl+hRqvrYeUxGF5GqvlpdyBbz
8P+F8ggRLj+X4fPHzblrCLOuVZAUj5Sq7FYjuBb4sqiHbnaDEEUv74YrljbC
yUP7wrUMKjVFR2n3Qf7GRkn+ahMO4ShLRp0N4qBKpRkRM/9zNXLC6OPaCXGB
zwSWwiu9EZr8R/+UwcAZWSdDYGv+ckEAGeqmilaRbwCjD2Ck6h6kFY5PF4ET
JG15tnsckm46+IjJXJl8ZDDLa9ZEO1ohCxsqpePax+8Na4K49lI0ZMzBH32j
yzxX57T0ZksBmzsd5TNnwF3uKEuSsdm7G01uNZCCsoA4Rxeu7xS5qQC3x9qd
TRBH2OfbBTpFoFS+XQ6F8OSnR6+VwaMgK4acXfEZOh0xzJzFAJIb7gIJ0L7k
CbebYNLbRxnGA2jhbxJVKGPxHoDuH425TnnxPOkJl2zAccsHFKyGQOiA3kEt
TeF1UjKiCsk7GUsVS9TZt6LYGFkynQ4TmkSBtlfHoZ49icAFCvFdxqyljPzT
wrAs8BnHN0esKIUtmz3wZWdgiN8+34fu90W4gXC6MW6Gvkd3DpaBBU24U4rS
OnIQjdJDwLX79qRtlLoUGlgvCeYy1nNggBlucvL9Wy/67VxpnJQ01WSS9sjM
WUjal5eT9mHDO39yRc49c8YzCwQ0Ys1mIc/+keyDsIkXyd0+miTSKGLp0crZ
yDZLHz1wjmtD6v5wqJCfMEmQTiefVeroWPorQicEPtbmUaqQFlNDklmqBakJ
dUKxKLDhEA5w11ZbtYH63MasjKYGGPXY3VaklshzE7tC9xXtiB9NA1w8bV/P
XSjoPGRTgbx9O6mbnXuUZ8DpWbyIVFpTM81xzwzjm/sNB4m/RJJK8WAjeu4g
3bLOhlGfqeZmVUD5RxVQsy7xbWGtENsrJG9L4DNBRNu1DV/uo5Jkh0qbM0G6
c9l/3uhgmW1WBKAK+j7jqYLywGy3cXqOT6YqPW9JFWuZEFfN9bgOymTYE7TL
+XM8Pn92GMw+3FLEN1bk3eSH/ye/aq32Wwnlnh7pgSqnYISg9quFxJ+Vdv2c
yxPSKALa3bvEBYoQ7pZj+zPXF4uNTVzVTkcwavL87PBP1u2i8m0aPwsq4F8I
fR+BlrRoaEgp6DzY4Xndxctlr5DtiHkqTl04Akb94EE2d16IsyY0k6klKeNa
AtFYkhN6NzRRSr4bk/DCYXvLByDVFEoDRhqIamPwVCh555A3nhL6cMKnPXIW
7A34AszLEXbPNHlntoorNR9A4oVCYC05YPbpBe+c/GOD/9A1Z1uKxiV8HbQ0
7vccFcTpe9Pwaxw+lWIrVETeREKo9DJ4bu3FsqDGAhBw0lSP4iaVuWQzS/vq
SUxv5CXI0SlYwDQ7wO/fz1b3O4c3S/AGr3wgMMNv8AIVQUJujMCzBma+APGH
7Jz1q96Hij7JCPPoujWR9wBdNcghB1i1ZQUQ3KLrMocDLehmF3nAhEGfHmZC
6su24LLNz7DdOUEG29/eLmQqFXf3f+9gwSw6TWWY9E0HqVtBkQ4S1zMt3qs6
umKDA6Sr1a+cJnzUkFpbpwrX1YHMFem8TMnrV5+MZfn14f1TIEoksFmRNQTt
S7XJA7m4T+VXTsGYQyq8Crwfg9uRADFq6TNhP/RyVX2nEct69Nax3/7Z06/c
rxJ4LsQrI1kGRJc8pObuFilbVgvHOAsfFg3HLiD1nrqgh47BAFlavbdDGak8
LopRkgH9UWxcy9KBJAA7MXkRZn3qY7PbXcN4GkgGow9jQ88fCjnETJf0Ofsy
i8qkk0EACu62QVYWxmIwUTK8jjhtRnw8wv7CyC8P/k99PSW25BRZb42q3Caw
on+BIw7mB0pvT4fzKoZOoW9x4DVuCzgi+dhIK/T/WHGrYYTfb2Y25mTSJVLz
3MXfhuKwNxfVarmAGMQU5D7I9TFFX4Ywa8UhTxm9h+5oYhMGZdvGOmR12I0s
CloF3AMdsafPBOTREfjC2fdI+bxEEfwXrWeM7TxYXp/ki5yQQf7ZL9t+xDzw
1TkWyQYCJJ2w5eNleqe5msj+psM6SitDeak3LDzeUTQhA2t9Y3iskJJXFbX6
lXWO1NgaH9KuewFekNGqtm6dSGP3B65+Tj/I0kvYJCpyXTA5WZw3lq/NCdql
sfv5iX3OOEubL4b2YLrFIJ00/L6dZj791vwMETrMTztUpYulHTW0SN6LJEgI
yRNjhg3JFvPOHZC4H3rCgQEi0QGCR2N/azQPcxGr0RkgABjt4z9JVnC4661k
gvyMH9kf+tiYK0/q9P32RBNFO+7o0CCzlvX78K6gpdyOcPyBrsBjc8gxNZzx
jD94DAJV60ISBtoT8YJZOJGKXFAbFIplfUTqFsdC1KuF5YPdNFUuv1Uwdiut
MDO74AOalKBXbLP/Z8I+pyC0054zLel4L+nBTG8+ct4VVtIlPXlU5Ch8FQee
eMzcfhpslJ1sG5NT/H22LEd/R3mbw74Z7KlwsrtunwTnAYQ2G2TFtyHy7U4m
PXrUXZt84Emc8BPo5lbd2frrtydlkoCs8gn/uGtTvgl/XcKSFWmhmy3f40AM
A6d1ruGk8AqK5y0aeARXe1sBQEDKp9E+/oLEoFPhgsUho/GgXhKz2TwndH41
RMlY3AXiWmjQAibNxKiODWRXyQSHPIk2qLtIdoPUJnA6+vdHNDycoC9awcHo
4k2xOmDdTxu1lXSZgEBCVS8sJYGQwB9PkeB9ErJLyi0yojNrY7sboEEqbTqI
oBI/1qHHc3cXk2tIKqgp2QwdMvLzq9GZvVO43hMUHtq1vZaU7tjiHTwwag1s
41Ddqxz0Y4FP063I0YP7YgFdbohjsO2S0ao12/fJHSj1CnkfXQFpJURM4ghB
l+NZL0LASX3yjZW7Lqp1nrj7xv5uyJC36eeP6IEpbgE2vDXjm5ToajRgBVwu
kJ4IsUuW8ChwoSGD/92TyxuMgjeE/3sr5ehe/IozGe/pd1VyI80tJKmVts7W
pocO5LH81zNxqbdxECBD1zW/tKL+C9Pt8S5nb8O4WzX+lV3K0IkCG4Imh+Yg
mHlJJXoqY67gWtCWNrsW1udo/wLGh3VlCL3VlF6JIhkBteU4SqnY0bX+g3So
Iqxrb5J3ZLap8sdUQtnpfGtfE71FmgDNBpcn8NO0rWgJ4O1a6u1H+DcG352t
7pX4nQv62JttxKCVycMTEGqPEDd2ajhw7W56p7kabe2IbpONoKWesXCuyv3N
MLO0s/2Ii+gsH/5pPoW6U70+0lqpGKYC9+er+AWTkSSoG3Wev6IKim8/mAlA
i+kHy9LEW0wLDgHrnZU2rJHcLu9GYYY7rn8DbJgd8V9ORS3EPV4bUTU3R/SV
rKb3kZlHslazwEGQ4h4CTdFpN4JvkdUJl/lxrigqkz2TWCpMXo7Ppk2l2dis
WATyx3O+0ma0aoW6KEFjpoLnhw2+d8IOKK+A5eFe2Bhv2uxMLOaijUpJmBqj
rmaLD2JCjNSeZowlCQRtGPs6gZFwZfChmebd0DK1iBWvT/ntcFn7qiXvkNGJ
EUw0vNVVv5xWHsMts1uwqksCHrsHYVn+bX2KXwv+Vz6LWlLy+/zh3sT1y3iF
oWimpZTfIfOXPvyau1/D8u0sx4O8bMNtEd+dJ97Ahh25mnwcKKnkNLBWnPpy
fPpkN4oruHfu9PDdNQD1J4fWEPRWNLlXHYcPDrHX+aXc3IwUKy5yvpyxHqDt
fCCA2dkXegnLg9Q1MsSBO2mGTK0XUrWrPV5D6q5uk6E/4rnPdon14pLYfpYf
PPIW6PcltquWHaNnh3eV39hOzrk5vmC7ouaoJk/V3KRmiyZepbSDa/A3FMQv
8IAPIB9M+Syr9UErrSYdsDJJ2dsOSn6vUEjbvhGLZ5VG6lDIonvkY79POQgY
/oPqF/g10e0zeNBOoqtIlF+cF2XVTZbFlFSBnyP/ug76IbI3UaU7lFvmxex7
CA+qnaRohJLjKiL1AFMsfORnFpLBV5H899purY530pJtPQv5wbV44784J5bN
gPLbdBi/jYEte5QjmocbJL9xCDQ1j62weizwJY7G3y2gd28zSSwNb1IXh93Q
HZmXpmFnQQWy3END1s+CcnLEH+Zc2DpuWGzHmdcPyZeUWNp/kjyjPjIy8jc+
XS1MtMY5/fBBjlwd1Wyrg0BcnJ6ZuaLqq2fm4cusSaURWM60+qyXSyHoGTb4
MXibq+fhTHaUK3XxpC44Xhy6X0ZHLfub9NO/JkcdWe4qdDcQoJcoJgm/fd9k
K+rzDV1eh77kvKs88DQACmatk2BZpnEoMK7WtXI+w4NFkXXmaaZEMof3XQGJ
iM1Ehc3lc08fRxIIVmZ+HneFW3umCfKdYM3AH8M6FBS+0jtmTfw53FZCPAyk
g0dW33pSVDfyPf1LThpOuGcYdr48VX3ES5q7dmnadwuPS9NHzhIdOlm2UAyG
BN3hcM5sb8flb70an0LM9Db/meSdUtm5AvB3zFnuIJrN2Oe9FiYDkeTZzzmE
k6SLv9Dc7I3vLouFPQgng/jNVLGz5XFTwZZPANTh8xf4QFaaUkRyE/5BKBLI
pOOt4JSixCrFhmwbXPyrqgW+GPA4KLG4cS2aq9jvtC7Z//z4gBYpa0C0O3U4
OIUzeno352H5oFxRpoj6N/qDUbbXJjUHjRRqUaBR9lcu4HLYhD++q6YGPsp5
obC0YyYgI307mkDT723o0O7PMF/UH8I6fEKMFaT/7E/oT8abfCCo/yczJ8ld
nMLYCgdfh4u2zzg0tuRUvdWR0UKMPlt2UxwRdZh4/6AvDjWGEyVzHx6ZpZGb
5Q2FKZm6rwzLpY9iDf/JsN8c9gq4wV962fMCEnnY8tsvYuFPkncg4qGHIQ4k
DzBjrgjK3kCZ8D/TagzyWGy2kbLL9KjVnVOxipOorYkaFgwu/qbgPzOcsd24
XUCwK0FR65e94Pg9vrnNtMj24hselzPc1ifUtE3lC0enjFIb0MGOMrRhvitq
doviXRjLv9KBZ0rngX1FRqgAQIRVeEm4SCGJ11SLUzF1CBqUmBV6ezFT2ix9
UkQLaP8Dnd1zxZwk7qpMpn2KhVWYlQC972OIJptUwyCNOXklUnAScnX9U4a6
reYh7Oi3Ci9/BXiZviPuz0P4aIYYuFqON3zPvJW/uBOKj28p+2v5g5UZy9cc
0ISH9FMz6bpSsy+yAOOx2eVgw9ckzHEuAuX/wMOCqIWQzU5E2dK9Z4p4aj7W
keNWXbgzmX2lJs8kmx687D8qG4zcLkla/mv8roR0i1QS3kt5LuoGi8bWFoTc
RqBHZkEq/xnDywZvBLo4iaSY3zO1TL1KikMsNroaduC4WcCrIBIEN54pJ3ZL
lVJGSVqXpkkKU5Vti4OMnwwl/Ov+bmMdxIYC84nPY+ByO1YiZFRV5A0t+Ue4
kzSJHc6hWdFW6C+QQod683BBJ8bZ53ssKnBgZNx/FKQPaeb+BEb4hWKb9xDu
ZmL7JtOZQJqccanUzFEVz8QsqNJFlvsYCwSaRWunWISF//sLnbWgyh1a+y+I
riZ/EAEQhKWb5IZ1Y9X/WWM5cXm6aVtaekLN+LKIBrHXhe9Lv+7Y5KOEkNBa
DuEHqNAMB2N+48vkM3DcXqof/uyerbhlD3DdXrXGhdR5eZlTVubac8shKqet
hKY2LMy4+Q+91vo3GKW/dI3E9kn5e2RfpPVnYMNJijIt83Ub9Gh4eq6B1FH/
2hraDahwtpzOYxPohKqPaqrbMsZ+u1kMGxtA0XyzuhH2S54+hcYgP/TQUlaO
McE+UtctpN0+fdbPlbLxIsoCrexHGc+rCA4HUZ/867XQ31XcfLkuOUS6zcCc
/nyH5SYpsOes2Au4/CivYpxs9WyZmvQByQ+RhqCtD/E7oVmItLVj9CISxMuA
Nm+5WbCzppUcQ9ICQ+pfMn5GYYwhg6Zn2Qy6qni51DNpcIaXJm8OHIbRtE1G
yKoPmlMBeE2rotgToNIAHY1Df7zetpjrDOTJLZ4Eru7TS3I9K7ehbLONhKUT
QvO+qH+eWS2r8M1xVJuFw3G9+KHQLHInwlpmX8bC0CqFG4RRiExKTN4VwZ14
mMUbY2uy6wVcEQwO7d78zmhSixB6nYVOeiogoAkZLLbnIN4yujpgNouAclAt
otg8IBwtdGzfplUIONwlpnm/l8hH/PE+Z2SE7nOLV7T+2XPsggU/XecTFHqW
Xbryo1lsoJZlkJrqpAw8uKVSAAHgaVarmpqbVQRE0CMtUavVN2idDtHNDc53
kXXlKgGuabg6xaeDCTze5iefyLc6hJSVLVFnwihcvrPX6be+LLp6HNdYpyry
8Ob2fPt77gzxJoeLpLtqKo/ZN+uD0v8M3LfqQ4KEKJlBDYtrLyc4dc0r17N1
5TJZLlktUTQmjZCbTF/zMPr3+Oj3oSt1SpXkw8qNuE05fCXK21jVqegERgBs
MrBGx576OJ2mm/wRLUwg6/HyzGRfFP7FOxq/1/6s9HcX1ajRXY84qSqLTZ9o
dCAYqKysDwEEm90T8PXeEIEkX+5zX2un+/pAGQ4iDKMkZB00K/Rt/sRYUF7I
38t1LJexlA6FwUU8uamxEHXHDkVhgwiHVPS/V0vozcE0O3wDgf19jGuKdtmW
/ywGPMNuRO79M6RAm0g8WVKetmf8d6qyRPSRiD3oYHVX4eeaDEY7whgvq1F+
1ynBbXUSs+/bGSsb52q931urUMA2Dwxi1APaeA2z5rrqMTOZ0lZnKMJpdeP8
KxpwWZMoRLQwKHUNdu30f1focf7TLM9Hvngp8qhnffyFbEz4o9u7+O3ZAuiu
P3bkllBGmGrLWY92BCdyLN/JrcqqaIUIeIBMLiGEReZCYqfocI5YaX0ixYQz
vQD5NGPAho1yd1gNAVyI5xSf54vf5jUaZlsMQmzmcL6e4QY2zzlHquxp7wss
Pi27xnGd0nmfer5RugfcniqWeLub25nVwkini1VRerd12JBTi6Q4Qzscyc8D
45u0VMyl7XHjK0h0e6tEsoKz7mnXAaXMQ3qMqNBKfoQrrFnbAepLzR+lzxdX
9Gflm4CNtx6otqxaXGFZyyZHvjVvFaSJkSSHtiJYo1aZoWbI7ggTvX+CO5MQ
onJ5NGxXwJ7FvZ8zdIZgzp9jvh/vZWbCE6hry0vtJhkhL0KAuQ5AUQm5sw06
RyCauO/kO86QjLhtCmHfRA6Enn+7awzpFuxxWtT1HiH1KwleWyM1h7a7AbHX
LRLvcffwMYnNpGGrDQMC6DFCuIFGGbHDoKbGuLs5vowF5mnDE4ZrzhtgoVNb
KcLbIJqZ3Gks3V/LertrcLKv/U8astzudVl5dlltoY0/2dPQ2DHvmvWCnmwq
btmy4Z0zLDCIAJ9o8F8kqEEJdL5yBy59sxdxpbRkwKTiq6DMtmceyH/rYeF1
civQIM6ALBBx+QS/ZYwZE8FQYuTjUKBrhY1a4JoTpZzsoO/1ZXEt8rLK9JUG
LYamlnEqSBokhEZP9ZLPH84a9WXaWljoQHyB5sFupXgXZlALFvu6MUX6Orie
okkoro8wqEHbMNX95eRhyUjl9QWT9jN2g4csqlP3DyNtitjhB9HIfvMdma4N
6737JLhMP+VlB+4YnFC82VtMwktG31a12/ZB5jjfAZeUdqypnO+0cRff1UQF
k2dq5WcKSWNvn8A5bmHKtICp5pWIfYAWrXYXUMQ7Qfhvjg3YD7nD2YYNRNll
248HKhvizyrPOe2anCUrXgpedH0M30rK7Hi7B8jjtgzpxGom00xAtUO2/bY7
2Nl+zFh7hRFODoLr7AJN3J0ORReoBpoEDA/qvvFuKoQAONKzYVKy2EPYrx5D
06HxIUwOt2TO19nAtEXwm/qD0sdU1EOPOBmc8UCCEqvzFWi7iyuC2Iji8PVe
j3o0bfPdQD6N/tstV2mZhaX6y+Zz9G9y28GnsTWFWqxeZMRwB0PsOQbIftHX
B0SzuxmN8M+f3H8vug9kG7/4ZjS8KNzLZkgwujnQb4avjex+R9/Jc2FmHyQh
sP2PNRvee0VcG6gt964ILJ0NX8abxsYHXKnwgQV/IBvXhFfAEpvbwmPLxSZ1
3cJvxiNDQBkf5/WeaKtg4QQD8Kv93YL5JMwIb+Nkaw2QNyP/2Rip3XexZeK+
MmgXX59JY1EuMnP0kf+2pn0NgG/3lI5CnuiqsCjRETGrRyRbW3aLRKxAQvZP
y8BWyhOeGf1Cd1IKOk9dORNRETcdh1b+b/31x0vpz5lU/hMpLLS4tKtUTAuI
3CD+lduGwkkPrgEnUNb+lB5UbmJ8zyTP97zeDhYePf9Wg7rl6LD9jzSbpPJB
OkmTE1anX4nbliKklvyQvt/SKS4CG5yUpIDiZ3OvGNpV9bqPnIk2DUJ5A1O7
+Ej1y0o3J4vwqs/EYU/S0EZ3UkCa1FuqUcV8LBS4ixkfA/bR5N7ATEf0BOfK
GpIKcyTiiSFfkQJEvcbybWM6vV1I6+hnVUDh2NOIZOVN+QRumf2h2xvfGYSx
fo96gVfSH7SffryMBU82x8sqVDahMUJNkQLzYM0TD9EFGvc2gW+OSo6tj64L
68TBjn2pik/7NZKPdkPq1La3Ww8iEH8kZnhOs5fQWKT6U8TKzHmbCRkDwrXM
T1t+ro9rsXRF+620SYEhCKE4Wt7EiLzAbuosPFcTXYOLBuFuugCvx9Zw2h5O
+2HFeMY0k13SlVAyscPA01IBvila+GaPOzpS474kXk+D+7jt7mMSvKRAK9sf
U97ieoVN+vX2MAfMrxLidG/yd+BTX/3A0CkKXkxwx1e5gy97YoHn7Jn1DFL3
zAviQjY/EO+sNpKjYpFdL86KNA9u934De0Rm0aoXEzIK9d+AOBsdZnEluqBr
BXD7Ld3eb2+yEk4ds2eI1Ry7wkvffUstyfXY1iS/rmc0+ZSOJdSqekMmUcPr
w7eWvFrNrY8G6NvA/AN5yW4B1MKOrj2y57xlI6PMdKoswKRCsbkNlE2LEO27
DDGBV/ykOmTetOZmWfPDvI3Z7ADmaYEDiZKLalrKBsGjsghzGD+0BvnSTl7f
tAmnFMPutzFNXvvqqd0PS047i37S+t5vDCTGfpU7JpOmwq2UQee6Nk0uIbDF
LaUx2w0QMtoe3/Qw4hmRE0Cna+qHpGQB3HHsI3zJr2vfjZ/UXw42wDxRGZQC
iJOSwvqz9Sv1rMt2OMVxPR77jg7eS1Gdv/5608aeWKPxXsJATILVTcvJpKOh
Tgxg+9GKuysqASrP51TKfhis3Tl7HDJ8Bmkw8rf1JrS0Oa4Ef/DCA/ma0d/3
A16eS1t859k2OQIxXCvc35h6t7DSjY2NI6eULIr8cwv9GB1M5XLV6er2sinu
FxHEjltpLSSYo+HVz+XboTrSIjIP7IYYqNA64jaUxESKpOj1Ee3a/k3ioCPX
cJMdHM5wAz5JhFWMjTetl1AITkDbh3TjbJW8EwVU19uHQlT4igNT+kExzmYW
XeNz9c6kgPw7psIpxxZTJ/+jcqwPErQ82R+AcK8h7HqO3BC45O/RGEYICEWu
IXh7zKzU2e1QlXJlhAVeDJsLkM8J88mVvHrG0Dc75rh4+W/vmJTwyvUfRqXi
TPCCC+y1KJZpqtIIYd7krfJApWF4bIjocd2SpUw+J+CF8ZHTMVtkeK5TVHkm
U2mj+2+BPsMtPEXl+C35peMLfK9vwqz8Y276PUZkLwIMw17InFfmxi0zpWRh
hWhgHI/PJWWj6E94drm+h5cTNSK2TdH4ZIVpFil36a7VKs90EFkZIeMJrwXi
kvDhSoFjgPBcFRdteTi4T30XIwWMp6ihbptNBmOYsVZwuTbS+wRAKTBBOSRc
/f+A5AwmevQyDy7gPt7kYjmlUUml+3lxaVVQoqY4y1CNZDi687mx56Uh0CrS
7qhbRODbRigaa6xcEYZcBicnuV8Mzd+xqhkpynKfmoiYoktSZ7wpXl41yraU
zAg4NyPboRmKBtwLDL7hgt2AaVz/fMxqNLw4pbSvRuukrRLHVYh+G9Pqhi0L
fof/EM47Um9g/J9TLJDlze56u6WCI6SgRSipLMOrpNi+BauvwRom8QzyOsQB
LiTyYSGEcUaOSYTfYV8EktCzv2gpgst+ehX63Cikmd3NAV7cjmP50NgCBgd3
2AsLemFU0fQGDxQlMWXgCi9xCs8lnfppl9HqmkpHkrg70KsrJDxBVVWB7H9o
lKaz30Bo87T7P/sFu7LfC8lURiRL8CS2EImateLNtd49tmOqDpuVW96vjyCD
0LN68WOVHRGBKz5iDzy+1ipllFNWVda96qIKeMh7fOmwWCHNoKYc2SLwbU4Z
luKVp/t8xpo8lhp1FK+RjlsTb5rIXMEQcZW1BqADbNKI1xk5MJjUCuSSDf47
bO/4FLkyLRRrunJOJC+smuAsWbHsiZViBwLED+Mt6INBdPqCjfstEYkHb+4X
nS/0lQsSOBaBCs2rrpgAZqnO4Sno0CiDyTwTEpaPs5noOFMWzLhjhpD/ObR3
1g/LMWo3rdA9yyAaYCWQRUEwioYxyrdBjl7I3b0tpcesJ0N7Ayh4mUvnEESP
OtyvzQZ3gXtjsaR9HJReuIjjYl81LCHHMEPbbhw1vNhfJcpzTp4wKeJ1sqV2
sG34yTiZoFm+Rvd3fymWi9w0PiVznW0+u2OqWVclRuKxg+cTqjLql7+yAz6t
aQ8OlM9z2rcZw2tYEYW5Ew/KBnaXgVy2bn/5ojEL1TjZZBECjNRCkfQy6vyi
MbFtlX6bkosFcIztxIX/v6+aJbsvf0yeNQX7a7gD61npLrIL87dlNkqG7cCi
vEae72fn5UruX5is/9pIhyBkWPkL0bW16OWCmTr6DmLPA21lRmD0ZFYbgamI
LEs8x+ORlwn3/FQCmAJVep8KRkaPmBYunubaxNQ/B8RbQZsNqYZRJfSjw2de
mUJgeooFtvd3iPTuTk6ISK2yYlqoU4g0ZtknPgZEPhSLkkYnhLjLxPJXxzw+
NX+CElWSAZr5KoYefl0KezvZRXjjq2zRb23TjHB4L17xmr5DbYBw9WzWpDzM
2uX54w4iaiEFnTpg4olWZ0bTVvzHY9549vIA1gCPyD/C2eer7ldIpYUnHqal
RFs+wcrTDqtSZDpWg7mT2Am64eV2pQ5hDLYWAPrpmdTsm42Lwic3VONuXeEM
Nr489+B0swbunz0DHbKB0ZDch+UwiRKrO8DZgG9sOp8xJ4O93IlwzUdvBEPe
7/gSKtdTGcHu624WJG80fN9N+vNkPKgNEOj25VH8WkkgchwIz37ftAIfW6gq
7MAQnXdac4/1QFKwLn7s11jns5ZsK4FaRISSg01Ackz+RAAbLHSvZ/c9sKAy
NnWtCVGhcsmKMZa6eZH+HdzbzmNQH1Bn37GeClxvL9jvo9CdPAnLO/P0rTVF
DRa6XBtqaHX/Q7OVyO/krgwTjAbICsSM/gKOt8f3v8sCAqarFs3QGVXia6MG
/Ir4y2oSzKKDmaqgCnyfETwh0nkXvGeQCZgopL0vGqUMxdMdOGlV4kbphhnb
uEoaDr7kY2PDLjLffOepQYAf1505VnOSFGbZgxRBhc+HDVlwWJdJDz6CRd75
+5Y+DNWbjS2y0s3hTTx0h7oS1TcjxPz+ve4w0BcC+9XyP7CLwEbQqaufXgKH
FuRpaaVo26r4kKTgZ9GkZT1I3tHz7L07lhRqa3/3JX+DbgFMhnrjAwh6jyMq
rlY41FfMTrth2xXl9D1OKYw0r6j6/hWDjWCAySuZhghi8D5W43u4axcNmyOE
/MygFrcRbpfLp++1qj1yA+vLr6OO4B78M37ScyccMxgkFWAw/9cqzyQDduto
KdNLouepXV3Ch3QSqY1P34T773AVJwt4vpzK6ghwRE2/WApAa3Al8uNpeJC1
FxUFe4CQDulc18QhGVWmw9sNoZI0sL9pPthEZrU50tPiOF9HCuxA6SDuO2us
iZEzeFU6139gewhdsbArAWHmqqEA/SOgj+1F2nz4MiMFkhJbGzqrzcWQM9MF
rOl3Bn5r6q/V5gb8dORavyl8giotXjCxV4bBblNkEkCF993GVFsTl15bq6pw
nrD1qDsPdt6vSUO4/pOtHZsCNugpO7gJTrLvVP3dV47Z+yzaBRnd+hZMDdKw
sK/cY1oIIIhc4nH2A2XKNTdTDx6AyJ9lFRZ1JWbRyNfbv6Zl28/rpja29DEY
Tbt+3JK2+mygFr3T3f4SA5EqxbKdAjl1zwmXkW7214AA+wd3x3tYmILX27ew
r2Ob7M3rSfcUj2qfhMPRAs+uaSDwDbH9LjalNIgvst6PuiPNDuMu9BGyiqOg
umaRpq42xl2RIaLOEXposnlQpKmKqyHUUPnwDtXnCOguBEH4CmsjcczTZFXD
2m0T8w10omMXiaEQpoUbweWT4kJJ5MxAdUvtBD2rv2UpSPq6X3PwoWNP82Kx
res8DWwPNDMskM2REl+WP5jwPD+8pfbulT9gx46EsLhtBt35Dt5t1kZnssps
ajMuHFgUfq5x15g4AcgoZKgGRAkVgUCfu2oeSEnLhXNkWppAi0gDcQ7B0JZ1
dJh+zgo3WcHZFekdl+nQcejOUS6IqOs1JB1OIHu4MttFJBSBLAY63A7IFUe1
lN5dy3uhD4hMPzBkV/JqVhvjSSrYbUWB6ebHtqnDp1wMWapf4npFsJxDb+Cd
9W90d6M8Gn1RX8xykJShbNSx94oeuQFqfxWPHvXRt1ljtGWxv8cenJJgrPR+
wQVPnKNQkFYE+43XNdMe5pGSvugMQZqpR5w/K3siqygoBZbLCwvxMRLItCnq
Pa/Z/T/Ga8cUiZ0kOxapQIhae1hWYzt19DX83AtY/dSq8/ddNywJ01tS5/av
dC6ChJW2TVi6R+jJoN+0xX5Vh7H12FyWtH+nrZ66RVSo8U98fOcVIhjyVOow
IK8WsV8KBgiaXnvtzkVRROt3X9drXK0Kht79zcteFRX2I4iqUXvoZjGDTfRk
8JVkh3vfnKc/0R/oYfhe76jUKWc8aayz1M11/Gg8BRq1oYMO8Bk6QCnOSEVE
92xI2RsXSEe2XaId1RGuSAtW2Ou+GLz8SrTIolRHF7eDk0AYV52bMSbAQaEk
q1i1gVyc2cBFT8PiKrV9BuLp81mkojTwEJ8+B7U65vUqmwddS2sYUuyjpwEz
ybgAdEWK8MTDsCwNJFSUcjNicvUXdhfyhTTDO2Vb/yatFm7cA4pud3SeFUN3
Wcz6enq41Cnbb8S4OisOzoa+xaZ8SVtFDbcdp+FYrFmQckdTtQtdJtXMvzGY
QMegJYQpylc9xbsTGyohQRfJL7E4BlKUviTv0tvvixYMt1wdLvWHeRMxAWDM
b3E/Uq2l6zV3Zt6/k/xbOGInAgYPGeB6GD2TAs0kcvjnVon9y2XsNTvsVJsk
blSulW9O28FXvEpkh/7oNoaUBX+gzENNPZNPWbqfpJC07toPVEaz6tmXz+wD
PV+S3Fkgj+h6bUtT++Wg3m7UgtquEuIROMMjfLbZgebR86zMXXFm4GKdMeOk
Kxhm0q5Urpvc+QHlCduLGFzwhPoiRGWsN74kVoxhzCQtjs0RCh3sTNDru8lW
EIG3LnhnO+5lr1KWVD3kc3awYmF7lrQEfI/PxSlUp2iWjkHh1rAGyk4L+QYW
HN8ydmm/AFxTTfovvcUAR26VITj/NlIKzEVZq/1qM4/6bFQAxmA0wlpcNsXb
9k6O8lPb4An5dVXYUhSOzLx1vZ0GVBsX1rnbji0HbwDM7j/AjMn3K7//nw1j
8vxUaJpjvsp8CmzjdEvo312MzGcsqYDT6as4V+1xymuc/nVWK6O+9StmLR3J
EDduEFrXIX91iHgtxVU51GSrScdcaghbX4sQpbuO9cphxLB3Pr4h9F3f7s+I
HvzVPZ2t92rSaNg0Jn7AGYgeah1KO2exQJj3oDzpsQYYzX081t6fbTDVDGD+
pH41Kg72HKZz8QPNHKB0Yc7KGkVuCokzltxoRZZZHH5YEBzp4m/NZZ6fysfb
+Or2jtmCsUdzCtLzCD5lridlTq608vIzhmkeaZ/ZD5S7CavDXEQiAWdyLxeA
1r6WRVtQ+pLfWOaUwLTHHPA4pz51BG9fNDL6DuKVPv+guwEAFnSnL/v+UP9P
nHIYUKFqEW6kcXbRgczBVGoDqjPmoi6KXugTwK84ZchR9ZgjR5v2q1tArq0I
pORw/CdHNMwu4TZgaEDeoo5AMSqxarnc5cJTMjG3w2JfLXwchO9b9cGiIlLd
LLRtpS2IRmV/6HXwHpig2UDvhPWa43LyOHY//BGHMw73YM2X9UeumgGo9NcA
zDaeTYw6YvECP+MwV9chZpebxg7f6vmuWSNBp/WGqZC0uEICnUzX2AtRw5R2
QOJPJfDTJGXnNWOVnNHu/LL9vfolEx3Bj/s3fawOjPK3xRClR5ER94aWvUEW
yrJriMlqwUB5yucDsbYikJwXse5lZPCdDsu27PSlbDk12DDFjngJDc9fLe06
f8OK8gEhZiL9Ky/gRyJdG2ePPoNiD/HF9K42ZE5lQPSE65rnDIF0ax54BX5f
rriHv2S+QoXkXWhjE5zhtDZ9YnP0ERHeear/uPpyWv0SWgfiSRg7dmIVNRTT
Y2N9lWb46A/tVZIT0TzorWfmN2c231zWsL9JTvucsTY8T0epFodWtKK9QqY2
b46JMavn7sLYhQHGd7P6EQu6lwZJc8UPpyZJp7ogu4Hp2aJwmw00TEpKBj83
kH8V/LJhMtvR2KJaTTbWDhcCBw3Pd+rWDmrD4tj9b2DiO3SyzsjtOfFBgc0a
myG+GrwcxHP8wDHGXPYLH2731kqX1SBgSlNtffefiTC1+nUz7ItbD056H/zt
6b5EUHG/XfBVLycd+uvlm8TSfieoEgGyHSlaApifAcj6c9bvetq1dFgWS7Jj
FFOP5fKIeY8qb8jLBOJUfUrFuMIL7zq7w6Al/zR/XVKU7qnGVICKnnP4hh06
ROR0b8hCcUTYaLqaWJJA2Sj2yHaM/6QlqSiWKPZGhUndSmnF+1ucRfGbljiC
rmDBvMmXtKlyYy5e+GnHLcKksaHR0Ysg95JdATmMvu00+vucYJfOgRtnQSXi
Mlt0bgDPJ8bmo37bQOm+Mm3H0oQuvtxzAeymQfbKio3YkwgwhBC1+hL1c4Ol
2Fk2yK7jrLBLwHMLO/tVRKW5gjlePQs4v11Wqwp5+BPIFLSXqa3jA4oWufCw
sJDig8tibzxtQ9AoGSUcxx5xqAOuyZJ9ufTn1ZNAfkcJgL6pCM0xz0PgLNop
RxHk6LAyy/Ua0CLoMtUOOlQIIXpyWfDKTAbjXMJLoR8GfY3HTD54AWC71K+B
KFNZrEa81vpjELWdzVD5RspaZNb8bMjxEX3LRG/qXs9dY8M5i1OUQdqfzdK0
MOsy036P6IMpoAJ6fGjSHAprtR8i4g0MtoU+mhrDi+DwqFs/w7yYcbVlcRT2
FZTJA0BC5YD4EN8dNOJ5Btsk5KhwEblzlFUKYWzma7k1qdixFjedeoCwbUpS
x+JQet0EK5yJyH+8+lu1s5mGZ71/lJaJ8iW2K4IaCeYPHoRkbXYCVSZYWkxG
KAsGuiU2qFn8xzIgQp8wpMPi8SYOKNMVKr7vtd+oPgBTEKkaJFxPLAd/+jMD
tZNDagslUZA5iuP6Mcm4U4JrIk1yvgFVLVoLinLQ+R1idseItRb1ZHeoqgcv
zrmPmMMYf2oObuOdM/QdSAMCWihNwR92ugNtZVxh5/9joFgvH6mLFktp60Ib
q+stGROdLcQSu8SDgU3mbHRzlxXfD2ajulhoCbOFcEW5f1SRUFKRA1ZuaPkC
DCHJcZa9YU5F3mFHdpeeGUVMAy3kgZQw9cH81O9m/Gc23WUYxSW5DUSpGvXu
fpRIDY0zsu6wkM39qd4sBQRdk84FtAsVaZ3L8nLgsxVjOX7XHL3xuv5MWRoO
twtMmOAYDxlETxYxm6jBComh00GoizTr7Y1UqwL72vrvwkjVszC0pS7qGFi/
wrMXFOAjaO8/46OA4g5RvBmJqbKBkV4DHMFY1SebX7YSW5EGEs7hf9MtSjxN
eNyRMc6G+CvvqWRbOZwEltloaK6oIY+g/DUlxoCIzadzZJHkkAaGz+Y1XRDg
hbxQqVSem0D0AgsKDrk6FYBwV7ChyE3TBvHdfBOpDzI4akv3ANCav1RvnQyj
k2aG4pN6FAHNIt8HWtrSPniAPM5+ICVzkWtWREw3lGH/C5BHZhlAbR/qoQ+M
ASVxgFvcM97pVw2NQJdU4xNA/f4gMUhb06wHOBJq0lOuKFG+gUAcT1U9TV2i
Oviff+jUFIJmAXIfxvaJ/2i+1bEUZAIKHF+zy4N8ne1lnLBtbCRVWql2HLSA
zYBVT0n8Eq+ForPFSP76Ddng3EO0WVqs55FvyovjpzIWfb5FmGs2UL06iiON
CFN8Bcmi+iPrZI/FjJ9nIfhG3+r3t5jTFamdbjd5NwJZCw6WwWv294tF8vOv
xB+AEdQmpoJjfanXl3O7+esnDMw/rL7YsSmoe5L0r34sItdN9qKhL7VLOQRm
p1x/5EseeEl4RuNCymvIBP6RkstyYNJp2wtpEOKu3jNkwvWwPFHnVnS+t/JP
i0wNjO4y+/3v32nhETZk3jfC0rRJLxE5Wj984bqd5Tw/sgDxClFSwVQbuz15
yzfD4CLfp2xghjb1ZPO6kN/J6C6t0teaHIZiC4lcQG+N39WzjoHUr8222LRB
3WUFrugcruyvDTPpfBcAReoBHsBSZLxOqwG6/wIJwOM057YQCRK7Q+y+3+v2
yfMgO6H4GdH559KhzMiJlNoSHOmQez0fFE9h1rLS9e09LUJpAJDkB1m7TlbB
D/JiB4wgFkzkONenBCByAA5DOl92OUEYPLvOVEGx2pxH1KyiyXiZ6cXXfata
B1omE0V6zbPCCAnAUH+e6q69onafkhJLmKAyOHoJGr3tWI6t+uKwPSvCaynf
BO0D0bt95XXIHTE8qLusPhJ3Uxc1sCdMjx1SvI9Gw626Uai/Bnk4EgSbkFWS
VlpMdJtxvwo3dEXpD3Iux9p6pKE+h0QWzLUELBSoouLy98Q9CSIXg6VvXbCE
fudM+rubaFIIpXwAUoZqlnKSFD5ZFsuLMgHU0i5kZbqr9Fekv9z4k3GWSHGp
Oe8uKwIWlZvaZnzY5vuNfdJ0sO/8Gp9ntlkLhbLNVhusvtlDdZ5bPQ6Nz7R9
HlJird3w0uo8Ilwkv6BrJ491TAe0Hwdos7rcT7/Kc8xpYUCkQJraeC0bItV/
ZxNSPUBOupwNWu2hhIxAehtN26n1V2+NbrU8H6RxvRgnd78Si4GqhH2Yo8KZ
LpGV/Fuv6orM4xo8ou9F+O5GdDHr5oyx9YBjGZT+1P7pn+W7fA+dxnqIPLmI
rcQhx5ltPMiux2JNeOexj8PP75qfiYD2D23Sy7xPTxWBzR+iQCaCZF0dfYeb
fsfuMoAyheq7zajze1ElrzjaX2VtW1JGM7Ijzhn3h6vDP0Noypd3/0RC93YB
xa6lTnGDDPpwzbQQVkSEbqUE+Tbo6NXq+5F3nw8x1NQ/l6ewKo5G8y25GPXI
VfNkrMkbeIqe2d2ReNWWB1VpOdldMOGTQFTZs1+refXgF56rfOfASmfhT52I
pDiRzrZNueDmN1Sr4TQa+3gQmUHVdQ8Y9JlL9OPT7XSZIUN8RtIgKQmERumG
+LS+U3rERquNsqvro66AX5PhhkzzV/a7c9UYwwzRbLxND642cfjeUAuP39oF
fSELKRHALFYkA7KAx/po84M3x1p7aCki8md2YLY+ILEBG3QVJTqgFVovzjZ/
YarUgH4w/eMqnjgen3AldQ6Pkh+BpqlQT7/PQWWmHPDkmiiJXtUl/Lcudor2
iO0GtSvhJQdjLVhJwydyV7zxUw/D223oZ/CRTF41MI7cF76sJKOvbob4fabn
xeGIn2xyIa3xnHWniOleuSiHzczFFME2M1soaPB+OV267eJHkccZ0HhNXRBT
UUcT5lt4eFFuCTJGf7mdRyQ/AoMYiaoM5Oednjli9qLAOE/nUZTz1awC6TP+
9y6Tqt4tTiCHqroOabaEE6sQEXKVCwe/uGxjq57l8KKLcHTYPL56F5gytjFx
n+f+eh0B269WeIAiBduW+T2dgwuWP8dM26GAb8QgASF02QZJ/xHyVQD0KGX8
9nMFxkW0gUcD4tkBnBC8CikqphI8GbA2U7TghTrkQ/l34rOjN6YJYFoC6H6P
P3iGgxkDdLvyVVLXmex4DyYxeo0NDFmqB4eduglVUnDj6uEdLoDN/povWs3q
9/TXXMlVk0seeprr1Nd9RqiW79DqLHQeN6KhgAokEBXAS/aht1XVkSF4et4O
bPAjlfyn1YGlH2YYOuuW8VzzIXGlgw9xI19sqFG0LrxUNx3pCCYHGGe0W/sU
h8RapUlvNgQjt/6Uq03iNi+sxE9fwA8rmg9B3dpyF7FFY04JKoEMRov/PI8D
C7EdX6eJqMRHM95kWVLACblN/Xw/pg04HnI9AqFGV2fPlSI2/ZHG5hIZECIe
E0d+qfdx6C4PZD5CNNOq8sE0FkQGJT+3/FQLqMRUkQWQvGOsGDKaEfoXdqjr
fBR/hLNbg+Ayz7q+z6wVSuaQyGBaL/9Itif4RCBWEB7q/60HkUUIQLw1HSgM
Q7okqwueQLQ3EJZer05ZQPtiUpJBmMvrjNEhJ3xR1NfKumY3A5CjE7UYO+kf
NPCbqrWX2vj5Rvqc3s45m7Olj4qc4qamsyxeY37XFQhDivdd/49qR/5RzQX9
nZbn4WRDdvssMsaq6/+obGFJV9WW73ftZ/Vc7iK9vN8vvRMyL/iGMXue9w2g
E2BlrFmHBYgb6gFpeJSfQH+SaVsnDT8HQx6LMeE6NotFVQ8sadnUbqJPmVrt
pTn6oYTOokbyhG0y4e/V4b5YFlm/v+hZUxjdWRGiAiktnwZtKGoRA1NjVIFh
N7+8vV5cQ78yIPPnEqyrDveAOofzDxRgeYWgC+xshB6bcAMXGiJkIkIasph8
6pvUazApN8ypp7kcul0uvvJSIFyqJ5oVFkaBO7aV7o3tidMsLLflcrc5fIby
XmNgDoQ8wR7EkBEm7mt2HzEiGPSXZjXYWA+wugWFhSUhN4qhP/GiNPXYBKUm
r4nwhWWdo1eHP72WMaDaOo50kV/JWdaadx5FMVUvhj9L4jMlT7861esNianV
1POgIUBOc5VhWj0NqfNkOv9sZxItX/Yj6OymLa6x+1/Ham4RgcSMVjWmRWkD
RDF4bqq6htyPWaxs38FNaLHD/h25ceSIed08jhmqawpQMop7a3cdwcHBmRi7
ewQ+UDISSwTD/wcYjlcQEoBsI4KvbeunoWtqENEfnBJJrHSYW9A783blRNWI
pRJ7CRBAAgwp+aDzwFu+54t83fUD6lVH1EVBB3DrRSruhHm3FTuQVlOVppR6
VO7EkBtmdYcllSwjyEYM9w2WGvr60eGhHvVUaxj3FeLzNU+VvEVs28Mho8o3
l/Ddk3857y3PMzwrDnlLf9qiyEeM7CS+UyJfZ1JbLOKFTiVtLvnpfB6EnUBP
P7QvWD2EHehYsQmHnB2GUwPvQQdqK5F2XjVu+uqeGmMSn29xu05T0HLY7Rsm
tsSvkKdwW9LY9XoUwH+GnVvAJ8wcwNbs6tdtceby4+Mm6XlMsIDu+iWAzryL
Ao4sMa/ay/ENjEUqYQXCM23LrwzApQp2wifWbP2ur1XF9EKO6IFn0xjlK1DO
eQ/RrbZSQ4oQRGEQP2gstUd7JldAy5wVJDI7zWxr2pd3i1aZkUTxlTwvYLF1
BqngT52trxBlfG1YaU48ploWSvSjSy1hjX503IW5XXk52Z803hSQk2FaUFw7
FBpsUI+lr1tyWkGGfbCg4spII6TR5iZxeIVzAmOeHybpjpHZ52IVrZ8Z3oe8
Q+dLz2tDSysfxs2LcwTzF2htyBlFGAeA/gFT2ztaauveisAxT9Nb2mP4RP/l
TXYqE5+eRqNXDe6ac9X8+SDK2iOPu3uXXERQSS3a5Tf0l3xt+jfYI6u9Ey+M
zSw8Jz7uXnbpUqIVqg+lmYKVrQT0Sa1qnguJX19ukdm6doOtvuSup8YxGT1h
cXqVbIXohT7fBfqW8bOTeSUMuGoUJ1zDmjfc2CjWBh/S1nj5bO5r38NmE9tj
wHig0qy1BFoMERN0rxXUcbfOevs7luvmckA7y51l2efa7HSVxxJ3B4JoWbox
6EL6pTRIXUcENNekM1KKf/fIX+pM0T3AZrY6uyZ68gtAqMZDwLFZrd9yhj1k
cy3h3e1zsetwizzztNyzedV64JLdULkOcaxwtseXAe3KbOnhNdRa8r+V4CNF
YXocU5bYExZa32ujgBYWFCWwlwhP5bNsqRjZ2SZttMkDlDNHUYfdgPzpDZ7P
v+MX1TW+C0tbUYKeaqAf5h1et8Kt9y2+F/8PpDaIkIETg2jt0zaYEOqcbx3D
SF48iQAbh1cBsD0We8vHUXrDvV88HcEA/K3eNQwKMwYKiAK9K2xcE6hNa9pA
aaKFyY718ul2uojy3EHTomAru8eGdZy56MSTSXQFn+N60u7rJOblDlFcMPYp
x914wMMzGlApB/mAU6zIsQEzMMtgJwkJBO/smU5RkAoKoYFjHiOfyR5LMESp
H1VUiLpcUXqOEU7ZRj1Xa4MIV+gUnCxpbX410zGBEbGj1zKngl20f38T+nQK
1eEtKts1cGevA35L8tyYCEUJErdJkLYtTy7gu46kXebLRh7s2j3jAyJNWpWm
5WZIkTdIb56sEmQPgy11mZdPE+GiiTHp23Dr6Qh1jAig6mDLV9nIsAynjDr4
g0oJs0+3GlGFB8BATaBFSzDqApQTVsm6DsIPi2p2XcyY6L80NV/FqIWgcyEx
AaUs0/xneRhKzRqlrM+fA+LAgIgiUL3ho/jy2as1WQNjTUOw+XOhqSjEypN+
vul2el8MozMIttqEuwmJJUTXjrRfzEcATdoR0PW8r1zZEJeaViUW1DgHEJ5D
THJIPN8j/+dEtasIsVPGqPmXaNd1AHSNAEgfi9Qd5gCDR2FkliCKeAffHrhX
891Lj3bBwI+RbrmsAPKL/IVLplRjAyZy9G4sZ/g0Bxxv7awQgesHHlwHaWBf
Pgp/Snrd7dC47aWEkTR0k0xmM9z/JcGL03dMbLCSzQ0lxYyFepBlaA0KnGOB
Ar8VOK6T6erWayzmC1MrN1027qGQAeBOnHaMqRvF1zBhfNlOT5ceLD3DGVmh
qOd+8mQWwThvqxhl+DzjS8yp+VYI9OAcMPQdbZiK/vGgXJVWvHI90eo+p9Ed
RUHcNn4Y5himUgyokn2uThOEvqUVN6PIustudXbNal/4va6KzjNBjZW386VC
3zEkpEP8P2G586cdYotOpxmXpHtMYLffSKp3vf7+ijKCdklJQQVpnDaRkdPo
x9h6eD7l8IFekfk/TbtfRf3ydBmGMMTOsKIuFMXAXkR0RQIIzRsDgsYqpVQN
9lLelan3onw8z4Aq5SlRsqV416JGWnpadLNnjWA4iKjDvuh/zfbrFic7A5kJ
/2FvPli4y8QkhUp9QMh8tkQuUSov5oKKzvb7kfNFGZpVkYl5HwXbj80J1EG8
nfi39Q9goGoLcso7/eqrMGZdC4WzUlxhx2WN6pe4nTu8OIsnIvQJZDRJCaZJ
UyFvc81GNhGYAHKnKdJNlSKNQwYn6OKcQXgaovKF7NnWCWWakMpeYCa1hjlv
byRL5ZVtZTkae3sui3mwyVeX+lfolAXsXhq2PzYDR/KsN6yxIYCGl3iS6jsa
grQl8gDl0l+3uVED0AI2tgeEK4jHUUaOeOr1eU/83Cy/EaHsyC/pY2LBX/5k
nTDxFu1hZDKK5kGiXkkTdEV8EG1VxDILsYCTQnIG2oLoxeYyEkNyycBcH8us
634TbxTR+rNwnzV9Bh7mqScw8LMVGlMLNTb8YxrdvdhvJgzdW7d0rNrOmwVH
dXeBGCvFO0ogvYBw3+ZvskmMdRmzEle7+yk6IkFc9+Y91p5Iji4MlXC4snx+
ii1A/ZJtVaGBAYxYJMnEpNvYn48ACuTlUJ/ilBoFXJdKcumziVLudjTsfFF/
jOY9xzlne409J1ChWx4cAFCdupuPLpfZrhgFcom+t34wPMP+vASJBDpV5uEL
riWsfTMKEopp5Nmu7o2sgG3ScLvSKlwX8kbKHeJpQjRGtbibPnIZ5o9QhMvs
cvkg+OZLhfOvi3JtzeqBpNnCEuKUz9mFVLhMaTM1bBLslaCRlBrz//XEq3xx
y2l2DQspYmDiqlS8O67nPZr6EEumV/62alxaIkQLzDhbLXwoufbemCJh2T8k
sgn3d3zpfmcQu0quuvCBSAUmkdvVj0kYh7EM/o1iFuqXn2Ddoz4mZDYKjem3
QhVUaj3Ue5k3t76nxyn9dGxfCCdrzHxvr+R2mo3lAQaN1epa1nS7GdU+rf3E
3q5itErLQ4q8HfqLnO8dDWrsRBt2AV45AzFIXLbvhJPgPn2sRIqaYuZXgbdY
g+dsVytjvbGNby/i1ZHfxUPny3zw3a+xCAn85uLicpOdbfFD1f+LWMBnkQeH
hqp9f0gINCXb8gjLV9EuKwbr54ieUazdTDn+xQS46Y3bAtRxSo4BD2tULEmu
57Z05tbvQRc50llO/ncaixFrvuxF0vi2yN+xaqV6/Qu1mJULzBk1Ufx7/ODU
j89JjTwrbHXd/unBmeQ9ZvNH9UE39fd+ZhN9fq8lPB+b0NjnHQys1PMdv1QO
hg+T4ylxduy1aumIY9pB9rHn24x6pwWp6s2tRke8EEavBfTrs4G9JcxpFCSO
K3rR6Bgi/Kt2U0GATqlJK7NaBygBa9Zf1BdXfdZmqCM91OrJ7hZIw+PWQuIz
ClKPjFb3Ke2SxRdvmWnQIYrxbTuLNbpZuejQX3thKdQy07QW+uc2Zzoee2lP
Lra5SciIOyR+tK4TYRL6HV9EPtzVrtv+z20WfY8DIpxEUiQbJ6Yu4sDIn/qG
uqNUu7Nz+7HUv6C4rsGWlNbhD4IjH6GKMADf/tZ3wTxx5vO8rQbO6tD6CSMK
kLHS7/gCqa5uCg+V2tg8IVgF8qQEXetMONtDttg+CXgGf2IzHoWTHgeVcn/q
8w5mQC2uS4wlayw4+zqK4KBsNdLgF44DeU3hBJgWUtmmJMME8F6aoqOUFsS/
H2q8rJwb8RS90L9MHUvaCsYz+c4mxjm1A7yO2q0TMLYbGcUx5vGxns6qb98n
IwR/Jy/m1y1kqLfX2SCCPwyuPOrodQQVAveANOLAUuQfOAUSJ/gpciWnKivh
+5cAIn/FwAicCa8IfGb11inAj1dAi50Z2VA6svnn2aFkSdoC/r6J4ZHKSomJ
wmxBr7IWEPBX67saPsu+bkidHehvRvbWWKbzMcD75/ACNlOQH+CoxEAI+wEf
uxpkALcOIQhvyMKLI08J23Zot5HLIp4iJyQSQsTH0bUgs4jJ83vXiaMluAOD
e5N+dMWJUbPy8zIjj/26E7UxnrGNrEUnOxHjyzRNxfPmvkfsfb3LCydaecE0
Ktwt6mMv3yEwLRKYF1/IZCPyG/I8HM+nCWZ2qBb33ncBm16nTK+NjhVadsXW
laLhxJhxz0cLj8I0UVxGUex3HBgMBdR4hdHyPR8bbSNS9K1rb38xOtWLtT9y
xBBqie+n0+FY5ZBxk1XJyfch5laK0Lb2Dc2sbd14+2kO8GoKvkD6qT8MIEfI
YM61/nbdI+gc3eiCupnJf9tG4D3uBtoMCoeR2RYxfT0Oo+kZNiWOE0Z4GHlj
VSeZVzY+swRKoqKLtGrBM2ySTtY9CChLIxKr3p9mns5uxidrPv51LZStUyss
OoQE/I+DSsr010K+QZQbYJk4mKpVDcz7cizT8BsPgYAiwCYPwEODiMuP33Ws
YiDoQN/wgudHtBgNqCZ8XjBDIeUN7b6O/k3Mj8o97gF74O97dEZmMjHV9sti
46d9UmSLjXIDnm3VF/E5if3YKkT1qB3zKDucFNwN7gIEdZ9Z+IgAebcNQjOh
8ZZBsZnFT32xUwJhiCU6yCOAntuHrL3YHnJRgv/KE4swwELvp2uDGlpytlDL
fUlouyCYuzvkBeugep+9Q/vfIdqQfhVd+QqqOxaBf2qb0b4VHDKVGNarML4l
L+y2ffqwvLPwQyxRSIVqxZqX7k3sGfSGnh8ntSA5oD2NoJyqTqpyx9h8P5DE
EXDDrtYyS05c0kuVYKkZex+k8O4fG35913kACEGx5UylPmiXdT2DgbeLnSS7
GDq1Sa5CkD1AJvrIaKKH5wv90JITtWCVtEzhrPyEAQHGxnR2YvN49nuWQwqb
1SfvWTH0jgpzdcKKORSr8Hgp17htzVrRAWjZpWo3ekIPDb+SSJ37lPvY0R8A
+5DkGNNJTMq2LFzgwgTXy7BBgb70l6ADOL4T3GUcIiuoJ0I3Jx0ERVm+G3Wc
hviIJXc0TL8BiM3jAk0D0fw0U5r0eRRELkvVtQHwN99WKCoYl7DYZf/Aau3f
WMVI9y4w7YzlQEOdeH8HqRQIUcBKKqfRYXLpconjp/kYGCSIJWdhG4RS1xl+
ZZ9bGq7ckjmiGG8DJoppNQQBsLfyJTdJoy7T8udqRB1yxLz6997uMHyiqXRF
DVD9kkIrlpizcf9Tws1LxVieY5/xXwMnqvDt1k+OHjDko+yvfD4nVGXhwP6f
6MRHg3F7c1Wko/htXl4EccACHriIbgH49VRD/5Av5o0BY2p8+G798D3ErV5h
//kMKt9WeRULb4H9fVoQQ5vpCrgqGuJjxhuUF0JKX7aSqlx7K3Bf/AijOcJ/
hYCCAiGseIRQsC7/28NeLayK3ACXQxcSV5EMwiA6lMgcoZ9MC6CVzfnLb80l
Rw9DvON4UBhfM465wNYeGBItUi5u2XpGu5Itr9bKZQsTKTcH061I/q8gzifZ
A59aLVJ1d6ROhKzRs02iHU4VxuXQbg5VpKTosfZevM2TUtOPwvII1wIl5zOW
xaTHbUzDcJPQcjXRipMQ+Ygh1BK2n4YsephMt6AWRvzMROeShdOYSHOc0rtW
OOzgK9aahW/yH/r36cnX+3EpYXj1LDpdsID9Wt07yiJgq/GoM+zAWunNavCY
yF9IwI67Mu7KpTrvapVPaDBDLAQH88UQwVZ6f7md/XWDbndatid38zsdzyZk
6fAx7znXi/h9C8C1dElQ1mPxqDuk98QmXt97FXfNYHDcoiH6Dy4c1HTjG1Qc
SGwHkgiUNdBvbMPygQKwmH6U9xjATY9qbdc87RhAQNNM2p00IQFr2Ltbljus
QavoGllK+AQrqNR/1X3tORcIiDV9m73qYd3y6gEwlISciqCfxQovstkk6F02
dX+VTY4ryLBJPoph23u08mbLFNh0OyHn/O0C4KabgBWoFRWCkfWAjAdBSYsI
mZe0lEkDvupvfQQMHLx/LWT+TbWpLzCTGdjRqF/17PebOswgvQHmzGk2smM+
O87J/N1ruq8XzuE0BOTkrAxCa/wgyaGJ7u5E0KZWc7eGxssQ8xP9AMTdsUis
TMjMinsNfLsS0TRg2QIKouc2hn56CtFY6S04MHLTIea6sTiYgPsHS/0AXKQw
T8Q7Vwz3Jc5v5w/SRYBgCTZ+fNmdkLmRJ6kKF5jsy6b/A2lbRy9tTw2gQGOX
f75Tacgz9SoljT1ndyK4x0KBHoBIAz4AAPpQMul6gmoN/wl2+1hHI803Utjc
3bZNX8KylCm1miX76PVw5R5TiycGvyIYYy6fKuXEO1EG4NtXhvVBrupWc5U2
x3cHfdBxhqrlK6O4yiKPXJ0nqtl3iRMCQ8dRzAjRKHoY2/eYlPkjYmBOxt17
s8uq/v9CY53XlB+dz0GjsSuSdOOzZIcyyI64OhL5bzg9aktxS0u1DofuFiKX
gOLyMEdJY/hoDFhgqqrdU38M+cQQQjxKCs6I93eSI/E1EsRa8OWdx8vLLLJJ
4Yoh2wC/WBgaQSNogIDx3EcD8KGlw1Bkf9k6SHy3WjPjzVU6kW70p3DlaOh3
h5XopQzpF2PW3GFlPWVQsxXE/qnhUKDR8Pgl7F1HR3NrTYNZnZ18bxUVmxey
omawC6FBEql8AoppSahT08lx5tDk3TnbdzdtuQPhEqcsYPRziKJVP6Cc09VR
szW++OaOnrk13C7kgqJJzruyT8TusmbPhumr7JY61aismvK0jMh32j4bylan
chkRcdti/pSS5izT1VEKLenl8zn45huABgv5XAdKKyJdZwjUETfJBeG0RD5s
IzX3yLveCk/mw6HdB9kHwW/mGOFlKXVxxh4jUZFvKnLGripUu6Z6EqvQofmb
jpr5rNwEbY6bx2cuVUXULt1Jq3cWXuvwgOSQsGx9IrfiEwDuZ6yzm1wvkjqh
kce6NHp4cR7R/xGHgsbDjO8A6DFr5aOpVWfJ1mOw+I6uAoxNK7EPKJtpreXX
qOKD5HZ/kXe2/j5cVq/cI2ZTB/N+igl1seSk4UeZhgbPjSlcKEmfP9DW3iAT
8bnj6K8D3Gvhrq4i/CBdH5zbtQ8SOnuZ8jDo4BqM8ImlTkTjaVlLykrd6fdw
htw/QhWZmx1UGgzau1/ZOEuKhOeifM32wPXycNi/W0ByvtsGu5ogvBJTqHMC
5lZdAHlPfpDJZED3vomxIBGHPyNZGVlty+8YslYD208nb254zz0IJySlAYbc
D5Xl/wcPiWvULTE2w6nO7Cx9kB2CIRHpJE0e9mILp/DPs4v2KiF36mHOCkXo
yU3a8GLlgQBYTILjcbHPufUCDXm9qJB07NKL1Tu8lI/TdyTuUeNfPAf3MR+U
e2JMiSYlr9scrNEsWZXNzOdvhH2T6TObPRD4+DOV9eoU9NXGvFGCZsXNDpLf
jbUkf8ksx2ZQe8RIiSyzKXe1qEcmoej0aS01TEU/g/6gPvNV1LduF03r1fKl
6QMCJu+86U/EK6aQ3P1M7SPOlMETYpoeNWM5tr5y0FwUr3FHNRQJCOu1Asuy
mx/u0V28q4mFZiVpUwV9Qpo2Evdeq3GblIIy482nnb3ABS53YY3B3EFgTFsV
Nba3iCVMGITIMxTkdHjYBx4lVaAhFMjdkvDngYBsF2uDNvT2w2JeGVHLdWli
FWA2w36OP3Qc5eqeUDR+EaRLoo7wTxvVevoZaujYPggNqzIg2fl8MIUn3rdB
3oiY+kr4jyRgE03yjbSyNNTUGxl6vdDRDapvWTvE8wZmTrjcwjpi8B3mjeED
gaEkUqnIgSW5pXPhP+YCqLtuVBeoAQDYPzaTmPmjk1rWBZZY/vVGuXHvyELn
t/7ax7DJW4KivjkYuqNGkRAbZFI04mIDDUITVytVDOK/B5wlIOcwFvMdkC/J
zWcPoULzwcCSGzhHUXSvBohVrp8ZGj+odsZVt897NlTxzS68aR3Oufwllfus
my/q9hJGaqBG8zOhtmy4KFuCj2Q/nMusrrj1oqBit0aG3a1fjlAHuX0rowof
Bo4oyGg1nTBa0yFIB2DCdD+Qfb5Ga0EcWBHM5QBOxrATgWOV276G8Pb3USz5
2aeGI8nS2jmHraVMMZpx/MGUwj2bzYCXlXrMGoE6VTscmUvVO/uv+D19mVou
1VXIMaZxDKJ7QRKlEZERA/LLfpjA66RQ2EXYGzzQaXxAoeOhAYydqF66deHt
VYdKQ6pwchvugfcc4hRj/Ux5gVTVe+SSYiNU4cHMhvlevETWQz0QBAtZJpEY
93DLtFu/3hfawuLvJHOKtsr7AYXf3n9ZfJDXrEhugRBp27a6A9O/k9AezweD
S0i3oQ8d013a12ZM1SQOC6iOd+5vFDkTALgIsHr+vQ44M5UtDXY11EHbU089
dMNhqQ5qowWK1Iv2zVofhsgf5zK9KES6/C9rzJ72ts4q1WxfJx9mfoK+amxd
e9eP8+KF9X40iOJpVbtPhQ5AZ77YwPuErOLnJ1tDbJD0qhEPW6wYVHImhzFC
q7+wrrfIyVV4EneeJJiZxOdx67pwuazYuCarqXxmj1KSvOLkcH7HXDuPpRMD
wLCCsHrduqy83b4o/HI+/AgpYHen0dwuAA668kB73DU1h5FECY5acf9GoMlT
nj8KYxwWsU1kmJELAIWUPJxWUkhrSpSvRnrDmDw4OsGsE8V/r2XJE6FrEnCj
GQMSLV06vMFb2t/gCRawccWykqrq+/KAnqehG6BLztLogBbMAa0eUDiTQrxU
bPCnROP7e711MmvshcfRoUy+L+8yju7vKxRSXoLNU1zKtpfoaEAzVlXOg+W8
As0AQSA00oZ2+oa4f2MUXPosN3g4HVFY8oekBpULQOVdovawOctOJBCmpu2T
05ME99iS+YXX3KtQnK+p8M6e0MshD9vuxSPaJeQnj1Uw/fNg1Giqht/Y5tom
Jj9TYGuIBR2pN0GYA+HhzvF3vuqNu9V5FKjaNJYlBSx6NakCYqhDsvTPgcZg
CRNjlK6FwFwFfREYGK3Tak65covl8o0sOp68J0Xvi727C4e/ipWtwCzcoonl
tmIJmZK7S2lNCNdKAubsPWkLmnqMAi/FKf+b1L6f1D1cPSARDINF2bSMZDXw
8zjRv64CW0WoTk1rJU6Ve3ekK4cqJfMbG4hHNxyh0uLJFE3d/VPBejdX5okr
0ldvbYbQxWEbL9DjNb+EDowxst2HyhGbQ/c1WhKqXt1C77gDllrL5WXApxx8
Wsi4HRdbjuNp5CGyhrOdcXwDREB+eVUE20MgBbRexf+WWEMnz4sJZ8LWYeDq
aq7G0E4SCflloWIUm8odGBs3/40/HB3pYwC8Rfr9Hs7s6LFUsPQFE2aLLDmF
QQFFRByM1ke/Yfp2Qznb9jgOIaM8Oa8WWBo3s6rNDYzWY76dQDEFE9cgG8xw
tabydxwsRvzAliGmCGnTtoC8CboWRk5bjon/epoR3gQ1u42S9Nh9rIhIDmh1
UQqxQe5kmWGADcYhxvEYFvJX8y8YGnfMJPiD8oNaDWhN+lunSLJiW5Ve3anj
MWvYYe+naeYKBg7pwEKzC9yJbtsuFmvIRaZGSVxrQaDIz8sLU8jTpRG1PHd/
V9Bnq2ekxg/U4HuqqkqNQv1NRzjjyIO7rwU6u9JnaxtbR0JHNecuS/oCoW7h
KV8foyNV0f2yPVlNYpm3aUXnmbZjbCfgPFd2h6r7uewyCJn5RdQR5Tu5rlEN
kPxHxFED3vOsmre0TCWahxnurRq0qzeFiHhACMY5/rBuwWlyGyLtqdWDHgaf
VTb+5cUw5LPxqc84pjlKj4wvjJjsJW3X/mmZPNjry7V1JKfulKKOPw5EcnzM
6t8z1kitIoRjINUAU5dgKbvUSItaLScwUVfzAwkvYissKhm5N0mlC5VMCXaQ
VzC8naSVrgP+dvBcusCHjzQGhRfuaU/n4G0qiCUcZMyG4p4IJ3CPIYffSrHK
fMnqfPGttsMDzE4kj5RpDEhDh5ULowahA61KEcTBlqHzzh0mXAtJTHcDDlGh
jUJdnj6/jtgQCqpjAQgG9IEttDoRCUhMDkczIsLm3KZu6eKaivBv6x+r8iZn
mp3hMUge/e0GhBs7nGoDlpKy9nVxA/lE1imWH2pgyKRNnT+r89xt3G0G4tod
lJBDhzzx7IY85ilEToeLtSKh3r/cY9IL82l2jFpNtPXIjwLSh/clFBbKc4Mw
m+xSQLKcbcHFR+68PIra44n1USd4pSZLFHOwXgcnxXETyTE43bdFsErTKaaO
ovTfdElTMSiglZDLXznxCzMP3PYGqTbn8+Jg5GMfCvD+xkvMWEKzv2/fpOmF
aDceEAKhZJ/YQKlrWCNcUXMgbyt/WKZQuC+zXDPv8wpeJBZEjjt5UWhLiJrY
eqPXowelbRxIPerKT0GYpDgbT9aR14pyynvvnCKKecU37Ht1iKPrqpIc8+QB
gBKSKZdYHsTZXgdoM9nJFV0E5HtjoFpVNL83SfdvtNn2iZPHX1Jt8VWgd78I
gW3goqgcchv3rWC++RFbCC+OKWh0HQ1wLo9pR2fHi3gn5QGaPTFzVzSHHtXu
E2Rc0D7Lw5wLiColKy5XNsdIu0mGc/wC8++GIdg6mzHpfN0l9WwFPs2mDRQm
EKksrLSlImKcCv/0uuKWfz005JHXThNCIhfRYZcAg/l7JMt9PqkztFcERTqE
bMOdq6v1eDaFQ4KzBt8Ipz+jV7e0GG7Wje0h3G6W+5Kfp/VexasNjUwpWox7
yUOjGaD7hCr6eHSiKfmHzWpZXLvqaUyltxigoyM4wi3mqBlGaGltLmICda96
JCmI1cDx31sp9dMcJ//p8vUYkGlqr23kYZ0zgC/3bZ9bSta5ed4xc7Vashma
VFGpCP3Ndl0LNV4J1EaxE+Ohm/6r9S7GFhXHgV7clmHUPFcRkDtw/22mVMp2
yMcnSdCaCwfJo0iWD2WhSrcsywp5IXJJyD4voiQhMDT6a71F0evfUzjcLah5
6COnJidLTXV2FvTQnTxXPVH4TluM9OSMV6/WA9XT/Wf4yLmQjaPMcLavQ36Z
j970vx7rFDMM2+aKFvPIlqT9CBQTyP+E5XeduclSQieU/6aGk1GN5u2SgNY/
PmCyqzAKpXKxhzykXyl7RfhxgM55Z+avwZGEROcQ/relmahujoAJmvDs+9js
KU6l85cvzhjIngwhU78c0LjAZA9SK0xNhmT2xzzGvkZZyDvJBilutuZ95SdR
lF8ew/7c2vS13gN3AHU5J3U6VICBlppsBWdm/JGwdnbxt0JWPRC5TF4cieWE
zHfSIigoRQvVw5MI/MGhq58BOIbNtaiIZCiAuiCBGaTpj088t8bh2/rugTHv
I8E6ppf8TEqlenhzGdzGvtairihhXagu6Lk3yEeXI91HmVLLCbHk55PRNS6P
NuXEqAnF9ILlyB0hNhhlWxbUK2LiCbtF8vTJrjxx6M/rN/FgyHh9hDutSaNA
j1Jp6qsN1c6fAfY1sAnnc07ziSFonOVip56F4hYj9TRPqIG5P1lgJCd+c5tp
iTL4EZZxVYGDPOiY7cC39iyraOrbva080iCscv9yQP3zVqjq2XfnYTUnzLO4
bFG/S25DuxbLcx24OOf5wT97xz+x3+WpffAgs89YSumik9PQYw2Jq7j9Tkuf
IdURSkSg9XB3EapPtAGfaBoOjHS/JGy7H/L/V3T6qU1PTB613OBE3UHCfWcV
M28jfMIds4XaAPx6MW8zgxriUYpNmZVdsKTNuZSGcx7kPwNzTTt4V67WU2WH
Im/s2BCBFV4U28oXCFnqx9rx8WIbWrjvZtDk5IODSvq809lEW6hvs1LvyCif
vkLV/Sjkwu0D4ghTbzON1bm/npdnJQ9tA2WpHBXjX3T6hgUwBd7faRKX4L6y
M+cusJFJQei7VsZWRtc4HdvfbwfwgyuDVYpq7lYsQ/uLqNjodMwx4NE5t9WV
HLLik2pMxp5pngDyI8JiZe/chkz3V87u5dVm1VD7SGNNnEnF2ovp9cgUFhDm
JzyRFtM86izvj+axrMHubLRynG/DlTuaBo68hCVIkFMVtrsHcMNCOwRvWRXI
c8KlQRWRxoTtLerTjjT2lxATniZKuKy6TpQMYCAHOxt/WW1njGghTQTmsgsH
nnjIqerzjgvCiWwAX2ptQXkMahGf+M4TMigJoNZvSq7Rd63VyEocoiOPMcVo
eczz30fvnl8jqZbuf4C6fuBVxAlKopPLIjqdDkga1EApQv4gNA9CO8DerLkU
RiwtNOFHiuKUOWlU65LLRfpTGXD4Uk/xTkHvcTxCzESNqkoIVMhGdRSmlYci
OscR3cjOLCV5Z1dVEtvKVLY+3NIo1Un2ejxlAa3OOpIDLOZwGofx1TbkwIHD
twmllD5yCXbZl0+2nDbLmMwLhAQE1ZT4nIS3vSKKjKV4fZmuHWxGoyO56Gbn
9iv6V55kjn9w7tTmhcBLZakEe0B7FHX3eizPbRt9U1MZQkc8HLJ8JWnS56kB
FfgoRtREhrLxe/0YYSTNYBGAmTV+keQQLSLI1PYiJSKfszb19NN+Oz+pk3Md
JM/X/VlkAavtPaBY8DSub21pMcN2hSXf54uKBhY4moId6jpLB28T11id4iBp
Xl2zAly3cpNn/6wuk0S4SG18BCyO9a7HOjc8519gV/2xwEhMZ6vxZw6BgLme
phs38DLa2C37U3PhqkEbR+yTz11gAOn94Uo40fJJXWZQWTiaD0R4mF594/CS
HRUm1fFvPZ/xuOFDQEttqa66R3lxsvctuXOYFRtxrEJNjQb8xXqaVWR4OUzR
hjS77bk2XTR7m7lWPrZLEZc4tkmU+DBpnjsGTxusUdZUSdGC/wZS/gSkbwaR
sn8Mj9JMd0tZNdwUABbTlHJT8GqzRKrueivIN/zOwl6gmgJwPvvyr0TGXYe6
maXvA1oxICctWhxZOGIuKqxq3qabkBBaVsAm07PjNngSMsAf7KOtltlNVTdp
bcZbftDrrggRjLmsvSsTbXNiTNjhmnIX/ppkZePM2BlYLEiqpOloM2khcwd8
e+BVVE1v4c3zdtuC0A1d+vACNTrxOrvwMvcMoskxa+Bf4zL1b1ixov16XLHX
aTjlW07sAGPIq6wNWknkDV1WiOOzv34JVGUxehWkZg21AWC7HeHlGilzOmWp
9ryoewHHTo3nh1AgRuJEMb93YJJYgVdQ8cyvBFl0/usprxe5P4tAvcCKP+N6
3ubNZCalAcTh6G9MWc/UbMfNSQd2qYwjnPHvgKvH19W28pzWROPpifcFBwrO
UpjXKV+zz1JfDQWdgocD2KZmVFtFgE4IWgWXa9q0t2tYLD18hqkg29ds4naN
UUzeWsidTf71D2etAvZzjDB7FR5TsNwkMIUed0l1ePN/HBpSrzZQv7LbgQ0/
kc6VIRfNz/9AJmuR3yhTyQaemlONQ2keVEZbDe3cVixIAwwrolwvubE0Kfea
c5OQB1RoDZJsMDv9gbUGBeD3aF4Z8IacYA01YTFXA0XFpMhDfto5wzGiaeL3
QyLJMmnJK5/a9dkx7xB5Knm1cmu74m/I3Bn0nb7v6p8bfiNPO68pZkI8Cj5r
cdOPv9BXjNh/mXEiC4FJHqfURZlrBFUmCJeL3txVd22+Q7sksStuxonqRRJD
SOqtG6eF6H/YF4i8hkDl2z3hSH1/4+cXpsX56nUzD7VnLucWdEZEPoUMEedI
4djY2JZ1rDUxoMu+An7/EBE6YCi0Pzs5JhWXu8zNWen3Nwls9Pf5EWAxQnLs
Nh0c/ZZRHT0+0pTKRo5qi7+3zX58GEWN+jMbwM64icCidltOaqPP3KoS+vrO
dxZq/7A6i+EqYiNirBUzO73E7X8Lv36XLp5mVB5xEl3bUsB9P+C7HyX2kt3A
Y5ClC95r7P4ccK8z8MRbl3pzHSFJIYWz4ogbO5WvamzHZcp4PkjKLG8+f8gv
WuN4RARhU/5hqo6U046fXC7x+twXlOyRjQdv/RnM7+uyF1ePeGikxZZIH5II
7pz02HauQUMIOt+DVVMsvUPTQ53qTPX43P57ZDK6mxK5+Iyw62GL+2YnTJTf
5n27hw3nb4Z3xJSdjPE5veVyW9PfUzWbS9kVvBVXuBu6Z+0G1/TxVqWBKXKK
94bAuWlab6vEtEKa9ByjlX2R2qLT8JB9faJNGXiMzNj19LZM4etDv3jwiKil
YvuNnCJLFsrnHSAoukv6Y+Kojlg+ySwmaXAwMhvP30kJZSX7ouyA5OgAL2cJ
vJzxAyAL7AeNrrFziT6VFQph042tFiBrruqzTK4vnopEp0FTQOZ11FmXDowD
KyX7Q7YiZVL98dMln+n+xu73qq8I1UQoCUhY8jE/s8TRHwmMaFvytYz+bTaj
v0h75zAOjhiS3qzLq7ztY9Xo7gIS8z9q9ZJjSf83pIDyoL/CM+8iOiI5ZCwX
2uC0vqvkCfwiLxD8dkdry1L9oGjebbUzyz/c7imjtNsUaPeCRmHGklkwJKjI
3QIbwnvkSwGsibEzxr9wutmeeh4pOx8zbVSobo6VsUWEDXVNqDZzKgmjBckE
pkDhjHCHAnE55SKSSGW/Pr0ugcaQCx4ZTZvrdJpVFozae5dbjjYVa6iJ+V/y
IVaswWb6Ql03Ig3T07rQn1x7wh+LHaKcNNok3010ux3AN08atqMOs2m5wd7i
r/9+zgdyQPc3K6E6cEiuwrIq6k7i6HdWPI4vFBfTtvgw7FOssA2cnQMcvDsa
a6sx7HML9C+896BF6ZJOeEHT0vmej7QgMn+CF3h5nimUw89qdij3wnnwwc8n
Uh6N0x8Wm1zVE0Sy7AvkBSy/BZ9ggXtKXRMCA0TZn3hehWvFcY/Sx88khXcx
yjCfRmrZZicZyOi5b75SO6ZBhATCb5YiZyQAmAGqEZeZEfXKVZmenBs7tTKe
Ow4it61rwJDcy822WcVlcTKIBgaA6CeyWzqJylVhEqJEG8tcHPtyJckYFq5q
ohxxcD8wk6pEXCA8FlcSshOQb4PHILhS0TR3O8gD3LxxuTX5V4Um+HgXyTfy
b6PfG26Z15+MWtXTyij3BtkM47vZdA35+7nAd4EcEpH0bE4l5e4rd4/xnkOH
CBF5lyqpaRbTVOxYpWNRq3k2CUXe6x0uOUClo4nxoH77oH8KfweQFwMZWvzZ
nrtFh3yIQZwArRdVvsB7lAXppboIbe0tPzgjzJUC8x8jRjWzwdT0WWoKoADY
07oK3EUGHowVLz8hjyWiJejxGhc5DOcgb1Tl4f45JuR9N0/7a/fB9VEgeU6+
gy4qaw2gDeCci8xgMHbGWRFekcjzbqkj5bkr6WSzEYawVjHKfWZvzXeslAOF
e4QPP4BF0RyMgNoQqIu92740S0SHbWf3VuNFaR3GAvdb2luYpePoexipCDBE
D7Bm7PmdcSVgfp7Tg3ItlNaz3wVq1yZiQLS2pShsYU68EYLIJJqrMXsY9sRa
G02Tg68YzQ5kI22ZIXdf7EL2lNI/1F6i2frTTkCelUg6RqQhC6WAn2HlYTOv
HAbo/ZBJRT/NAC28pxugWtICcoUdsdR0cfI7WhZXNKnZ4X2DLuFEFqQYCQxD
ReLE63LwlpHVT2Gmqbw46/UsJbPZBn+s/YgaQVNKCq7lVF+VDvOLvbYU3NlA
QxNAlQsS5diLhR4qcgmUlFa9Sz9dxizJ9nYq2SOYL7H5Q1SFmt4Y79Zi+RI4
ypHupAM6Cxr4uzrgA3chi4vjtpXtDN6qe7XoIJsKTtiwclCHA+B+P1orLc/d
nCOxQ3EEm09oCZ4nNbrHkUxNdSwqa3pTYCmMBLp1PLuaXKJZP2nkR9+Lreun
FDlBJfA1MKPa9IDEPj+ypZU3QXwXSeMw3kXAaqWgpJ1Uh7ZS+KXqK4d5ufMp
Op5hME1j6EYfYA5CN5psLh30SJKyLh7+/JhZg7A/jtbV3WZXH7GjkOHmIRmL
6pbgpE6++4Q8JkrBj2saAQE1YvGv8u3332nIqmYNanfkGNnnx4Vmc4QPVCLc
w0tqH2R6rlu/EqKcQEayPi6uctDttdIHWSAg2CGCp2kJAR4LVcPbd/u+lnuQ
1qGY8p45kQSZZVHVeUJWVFZqM+B9pWb703+t6j2QiTBGI1rNzKlFCkpzDzRw
VTu0NEuO8NPfSIgZYJQXzgmSU2dIQ0cPKPm42F+s0PBhchDQYzvK3rZsORtq
iI6G/w77dx+Bn4F3oi7vvykX+Ul2+a52ni+erDYclWLtKO9Bf1nN4mPICzXj
o/L27c+U71q5JR8fRlnPl4GnZtbGtd7QoG0y6fKW5c5Zjz4d4has5REKWglB
1azPHMp8UxEhi33Cd8i5a5xg2Jo38tEtlUSezjh1wqnKOO+XU7qsECDHa8IT
1Mv9pbLu99qaBUIZsjJ9aznAWnJK7PiqyatLGfQlmuiC+Fpya+lxEkVe8D5k
l1Zng+OS22i7iaofIf0FY15eV/ZSFzGqOmmVd4ktmo+HHo78h5dFO8Hf8uj8
WeRhRYAb3m7DY747I2VUwsURzqEbc3KR8DIFkimfh35FIPCGPl/2Yptlp+Oz
ygNUZD7qpTljoxA4I/TCKgA6xSnWRdXVBeRDLmxMomvSfZ6BijaZXA56uFdl
Z80WBapfRPcehfhnVL3Dx9qxceRE2OXwmi+c57Ks/tld9335tqC4q9Q/09z+
JSJ51SQFddn27NYPUT9ShIMKh7LI+YY2IOHzno1XtdMxo2MRcuTiAigsv155
4yCk1n/JNHhCaFl2/1ggt2rQEZ1lmuVnwdbMglzOL5ywLJVXUx5lJ8E//ocm
O73j1iPo2osA5Rvm48X7F+9tf5cu3w0PSwXuJC7J026vIyZQqrz+RxAgBIN+
mvUkSCHCJLzNQvZgo2AWzoRSdh1zx7CK6jGbKbHjsdaK50l0qys/uCvR316U
Qe6XpBvya3+toqzLOLdxIEew9K8ChRvkufVXCaBxa1rIxTdb9mih3bRYLJCX
l1sRmzrD6LMideCtvrw3Jdw2NUiPam/PRx0ufwiwum9kNZcugnRly05uLLaA
oG6mI42Blp9eWza8e+NBeJorHYTNzNwYNv8XfPyzaIVzk0A7wN3O3Xc2Cj40
ahzvwl+R4wMoJ9n5YGAIOS9v9RjNKDTOx0jXcEjNrVuvKL6WWsOlesLsBD0F
2vjZGj7r4aqx/kLngOgIOhQyPf2FnYwzYw/4TPq3yQ7SMvkhOlNgIAEcDKHb
spLYW7fPQGTRN9O7jvDOXJtK/Qnc/o/Z9w4ohrhIafOi46FXx4Op+5kKohHF
3NRJESyJAeAAx+wfPWZzVT+jUhrC1k0pq2/kGB0scBHiS693ULmqI3zZXoVM
4AALbotPD2ICiuv6e4NmD4sfboPGpEVRppNXRwZiIF0Ftc4UCOOI+ObcgP6e
7xPaWij1sYB7RFfmfXXS2wABRTbHSCyNwL6sz/pRefZLr2V7AFL7SA+MaX4e
4y2J/Fcdg8KJ6qWhyyQ2Tf8EIvO7rwRaf4HDNRwVdhC9VvWvVD2zCvrvY15W
WxZY4sg2qaF3Yhq7U8XLlgVFDspCGnzwnsR1m6j+zMKqtMqM3GWQkhlrbFbH
AAMWHJlkaF2Qkb8dxvZcb0XzptGu/dwM1eQz7vGuEvnnwTIIhMhlUGLS3oN1
DFjv1v2JiMotSviOLLMFflZo2nIRiGOU5pfrXtvmKSeXR5R4KvrpxerdXgOU
Y3YbJ+9zgvCmGtmskcOhNNgvWPPnICSbaD48lvyfTUvRcS68/sfeaRgC15Dz
QUaSoZu9xvResSG9JY1lDkImrZ6EH5c92F8WA+WNr6Fwxtz+RK3IH2AYaW0I
hBLpCmGxqukM6ZghzbqYio4sRL3rQcSYuyxAq24WdctiO0OuRO9SppxwUqq1
pnKdoCW3jrozDtXbHZi9YdMwv5fl8k+0sMjHVfinrpy9bFNoVb94hSF756sh
Dee0YWUooFFGnOGiZ7etwJRRPbPz9lYe4TJaBUVtgqWmQ04MgJXCy7nfD0ib
IqZVHse2Yg9Q1SbdJDJGibu7R5qOb+/9DlnkrTg7cN9f/jroKOk6uSI1vfuM
tmoP3wzBz8rsWO8V5Ivx4h+6gH+jnLpxO0RJ0upUDVF0kC+2WzDmG8ZRjsNK
HKDdidZDkrYqEEBn8vA/Nsjkq5gZEHUiItkSQp9m/cuKtgyRQW7A3qbHpOGe
NNAjgwYdUeE9OVFrEv/3UC+R3GdJuZnF6eGqJrPnNsXYYiFJPN0UsJQI7/8s
kbUUx+NOxWDspyBbLjoHQmvDSBAypmIc8Jf7Uh2R6xcI5+s9YhAdbmw6vg4x
kagUwMTBhu7i64+pA0hveJsun9LN82UQW+WGnZ1f41vK8OUs/drgpeudYOuU
Gpab1pJ+w8J04jzMJAs+6eRvIdi8N7tN+PWQmtf+i4FgVPrZW3TUFG02/nfT
V9lnMwNkYu8w+moIkd+Ry62icvyYmlXfPoVkFFb+8VAIWSJK+EuVA4fC+doL
aPvaBUkPd4UNr6wpO5fpFaZbpAdsdoxbDHbKlJhc7XnisYoM2ybgTFVlM0tz
hNUUKGunrBQzfzQrR99xU0Yi3JJtlVlt3VXpVzTx2kqglT/ZZteeN9juEJqv
aHcaVzvlZ4LrHDhKF8kL3k6LpL6Vl/VZ6QEuKacSDEBeYwvxJJ7u25UutFjt
k/NPYv5N4YLyxsrEySVCYt4g9dW6rzBKGMuMtxPys+cl76wsAlNcVhFyEMP/
6DLn6g2SMZiw9veu4W7yPUeVb+i2thsE87UUODjS+eH+TJgODzcNzxmTl33V
7rkL13B2KfjwLI9nDeMpcrguSrkEcAfaITQTUvJBtwkht5DV1EwaEAiQdeLl
oXZcp+EpP0g0ts1RYpFaAEFzbt7ZKPqNwI/dHqxBwQrAN4MLn5OJpHfJNMBl
ZLcZdi9RNjrn1MxIGWFmvfBAygeowdWHFElU/oHVJIj6TlsByEaudkiunMmh
wvO3CwOYFTcQ66uz3Cy33ZbOUwCfSXsbrWsphZsJCATQadPJWWN2/KZ4FBH6
nzt9ROwDXcvvBu3DUY3939qdvfImWHkDXT7Seles4M0/iLda/Hp/eZYP+M6T
9sVTwqGAxK3oghgc9jj9G2oN+rOHWaVN9kwpgiozHug2rxZu8LELdG0W+Oly
Hv0GNi5o5vq74h3UAveIJe7X0N6JozsxQCKbK5wJljAJ65+YJa5Q6wllV62f
i82dz/w6xgcbckj0aITUZZOC1gxvPUL0O0aSYxHt+hS6k/wurhqUO+ekWNeq
ljjUcUmqZIt5b6DCJMK8ct0CICkR5iQ4TwVvuZsB12Bi8QRtQNowQiQ/Wu1R
xc9QuTlFzwqwTQgL/gYYX9JJuF5f/0hOMYci/NyCYc/2G/8uM+qUqzCQGZML
/SEigGajUKWFo82WGA/2uzSO54LeydIJ6jZ7wFvasDTzI9Fkw1p3UP076f7l
oUg0m1IiFrPDN2qUpZVFRRMNTibtNhgMyv6yhU5/rA4u8A+O1Kgyfw4COB/C
0RDD8F/fm1U1rlQA4lWr5S+GorrVOs0pTPmI47Cq2df+kxSSr94bE5Z/eRnI
URXIh8U9XzQ4qUN1MjjYeME7+kglimooojIbPxcjlx+V4UL30FIQLMpR0aUv
HUGqbxim2itz96ofxpyY118Agve14StQgYu2FkRCwZ1V9iTIN6YgeZnarxF/
rKdaFC2SHp5tKcw+1ZFqylt8MbMOM9TrpKaAk562VtvTsKU9/62+JNQCgztT
TFSvsg1wONsKFSsgWIerT3cUjj4/NK53T9zDyooxhzD7Pykhj/dQKNssgm8a
0ogSnuv0T7JEMZ5xfkMyycM1f4RnJK8+RQUY0hL1U9ySuvkWavPQ46228RPy
Av7b7b/fqJOr2f09ObKFeEofPY7cq+u50GTLM2ulZFKJIF2uhKmKCvILuMgA
UM0TDLMTQwEuwyD9w5Ft7Ek8TqUseGWlK+uetdjZt7JpMqXA1IpRbGCY1IHt
KWLY8wzoT9kAnLKt0753l6qE2zMfleQ5crS4bDuOEFzJtmXPUlJ3kgZ7AWHW
BwWSHbke1zcmf5+JQowjR9YNMFySFJcT7QcXjseosyYQj9YT71TolfuVmmOM
+aek+ykCtR4QQeAeiwBfMgFORfGSHviVxS+cwpaCAW1xBQVq5EtyDVsQlr+u
lQnwUMfypiz82HrYbfibpy6KYXoa9TeY2DMNO9b+ykReqXwOSEsOgFNCGJ3A
yGHtjXmKZ3WkOYzZPCwIFOOiqmTk1VH/2KGzLBCnWPXwdWkbiuXqEn9blxXZ
o3pwhNO3Yxu+2F8gyp71O8IPnpg6GJuLDw2cRxM5SJK48G/5vzdULWn48brt
jjUVQgDNy6iOgPtmnWt9jOmsh42CKCgNZiLS+Vmip7l76YqhfLW5BqgixW5M
vIyGObKOljQNlbfcxsNVFCjgeWMRfh+Dan5yQmkNzxhXa1uw7mfsUkPZeQU3
csYD4DdWfIofqDnVphMUVhfsGvelTNNry8G/KNRHWnnyA+Jj6zDLAkglVeb3
45tw3DEQr3xJ8LIrPgFucY/630+qQunrh9Zd6awDd1MVsrIVnc6SRg4CtpWH
BxNeP4IkrKvrDycC3dlF5kObuWYgJoHI/17qXvWQYk3SnKJ4dXXQBuebBWo0
Xs80eRpT1bjkWKcJ9D6QUNbDW1wfir2K26SOLQtC2cL+SfE0AqBDMg+NagqM
D8qm14b117R13ooZ1EcOZCnTrKOVX0+5fQeMyDnw9FD0fQCkTt6Bnq7RSA1N
4lJqlYwxFNjjSp5kEz5I+qiyCiub5dJgMXNHxRlqOwqGPKkUbI4ORy2kDQy6
N6Xm3eZs3ThIseK2N55KSAyCpBQD97/53k8vevEMnXke7y8ffPMUSCRsvSCj
BfRRs8MRd9K4r//wwRN8O/o/oqp1QP5Ct3fLZXFH8mbvlu90VJpfOkNnPV3q
9fT1f2GnFl6Ex9hqk/PkwH3qXzMAIJDfU4uHlgPnqE/QPNF2yOv6qtQxp6yO
NLZUgc87UZt7kxP70FpAHNsJWFiJVWnuqcSwk9hDSUB1P2h6iEF3TAvLZu8U
DXqe2BJqnVKdOK3p93I+vNZf/hXOAFQX0/m9CSOa3Y3kN+/ZG0s5E6S7clBv
EfmQ9RjqhKuHQnqFLACRr36mcNRhcCEN7VSUO+G26dAaFed7fSrHMXduDgId
XL8nzLB6zUnS8rJTi7BQPK+ioxa1EbtVsUiZQaMZ8AEh8tU0bHjZBB+SitKH
+m5qEkgN2fO3X135mN/uNbW1SmuX1rHgBT2e9fnkuRySyfzxsB0wzqi9PuY3
qtTp9ViyqCSI1QSJqESX/LH8DnhYmsIstsMPCCIbINjKTEWFqgirh4VDd8YZ
vx9Meb9KhPHwDkqunq75+HDk9QiaMepPtv93B1QuXUUdle4a/u6yzUsRowG0
R5iAYQ9aEY2/l/DzWgI5KTGCpg5VReO2fB1E/qo5Kgj6sxrxdoAC4HuALLXn
OeN2nFFpeGw99avKZY98vJbBYvcjs6NFPMQHwcNxDVBsHzU7vm3jzWWql3ub
9GpXDKP5rBI9BVED04Du7PvkEL/T0lIy+1mq7lwR51JSyUOhglvh6Tt7tUz6
SuWO25cLjlwRv22ucXSvQlJ9X3QEB34bgS/TzQK+/1gw9RYNBhQCkzM3XgV7
MTWl8m61SR4LsHm4q/GPuAm/astlP/KiPJXKPVFgMJ8j0PmwVVfVqGwetZwE
sRt9Dj5X+LOp5eORV38LJotJI7SyR5FIFbgWngzMhP/sK///DO8UpWnEhxw0
7H8mEawYNlz4Z1g6UwzNyKujjLEDTt4soAlZE0SAzf8utoOIJZ6tv9GkbmUE
2DUn0fjnqZCzwwd9RqOnJ7xj9wHPOmA1YtqmzI3spxFz6mKOHHpCo6jrAu/H
GrAhgvAzIsvnKcGp2pBnCGKQpR4G8LT5lNTGv8UeAg/zrLVMQ72gnv1Qrxas
t1P9EjLkrhC9h45Y/bcSAxLom5Nyz+rqkA5N7KnfCcwepqsJ8vWKBucCJQ72
mGVebSF7gIrZL1E4jq6mgzFfE/kbTxuPeUPw6PNE2iDc9/KDM8rExoWUNy40
Z8F6Obr4hQQfDUnxo91faUitKMfYdDILP8Dpk45WivKXeobC5W5gyCIvLBfW
bHmTdxZ93x/IMzP99N2A61hCDvLRs1HJzq2Z6NAwQ44mLAklkGVGGPtIj6DM
+TcjaYcBDuT7x0AbtJ4EeyoDXj9THPTuewmon8zoF9JYkJWQXeF4leXDoTlG
YbIYHkDa2soR+BEvfitiPq8rvfeD90vhxz719o7jS8rBFmi8d2xI2saWUTGp
3izZk98c2O+5JYoXl0ITiJ8Pmk9//XXz0hUjX+5JUuR2s6n/JehpH8j909bH
3ckSY5naQsRLeR4lX+awPiTDkhuYr8Jc6z1wVw6jjoGCCpeNbvSAhx8qnUeA
2mzCBN1wwF/OfjhBHUnWKUq8IMCyYlQmmxfPKOCuB5/C2tR8FndOlaf31Y47
U8WxL43P3e3IEvXbcA6ToRN5pJWVvYV5aD/Ji+UHXJemrnI+VKxg8mSEDUFO
iKhdafkCNtZVJVhQZcVeKVogEjwleXd0uXmUZ/j0YJC/BJrL+Q8rq65WDYKW
+BcV3j9c4E3b70hdgnOj86b85CBAiWOqBHRj3reJUmXK8NCql7ww3+x1+WO7
Q+YfwA2rcFveu0SL+g+QcxYfMUpJvY+TPj1efqG7uOyDVNIcTbgWucpmEUmt
JPd6bCWq4OBzEQpFsC0pr5NRFmFcloSyUkDsVYqaThn8ETFr/4gFmA8iUU8z
KSWeQP98QjkUR0ZqSGQaXRH2GHaYlc8OJILfM+5VSwla92JRLvlhBdCzRmrs
8MAzqPq3UQn+BkA2N89oZRfQ/Oy58PrjpHiEoy+c/ZFEAwLokW3FK2wq713W
yu4hczuhsx8HdfNr3I5KuQL6hBFXJ3JNnCOjWpcjns8QE/2C7MHRLIU3mTv1
hwbdDTjO78t74/QLWvjt0qy/AbY/n4iC5/qJmnGyMP5mr6T+Sf8+uX7pehtM
RZxioli4n7yBZrRKYl6Zkd0nT4F8idqQya0JG7BDxAH1lPBKukaKDcyUA+Dr
KFRSi2oQ6hGvTr9ZwZSbrLe+/me0fGfPPtVtL/Ir/8uFcnlz/j5E7D/EvifP
NuQgTg5x0iWqC4I7dF1rdHW868XMcdP5xmeeot3fylmJzqloEFZcPAGXciNa
nQvS5g/Y2ApVxZDUdRwpgBTnF6Gev1m6tUkEeQvhFoTAsliSpEib1gGf1pL3
mPNzskXqX7caKz4jxEoC9q7CfAcEgN3aIdPW3QJPioDqA2iG8Nhq2AUNCXC9
PLf12tUj79kyhvPrR7MFesL+7RgoMNsZZ/lmkR8/KF2aJsm5VZvqSxL7HMHK
XAwL7hneJ3ffRJiqnEG8TQzoBsOaKSZyVBT+PSyV6UnHfdWoANua35gKYoi4
xhOn8tu2vGzTgB1viDAj7tGuRhC7O3wzSNQHW6eryKGJ1tMKSYG78xJFmBHW
MWlWYrQb4FDmV0VOEEJqcaqR1FpiJO3fjzs4dyKzn5LrWZ5yNiL4BPsuXedV
Liurah5hjE6Bt8nBJy/dW6IlYxFNff9PP6XGBMpqfo34zJmtJIrkBucmnBcj
qvonTgD6Zug4baaTn8EaukmzcB/RO8e88XBl57aKkGnFeEpO0Wl9eq04sPnv
A8wDC4cuNFjhurZJDkHPBaergICjLQf9zjOr8g6QvQTZ8aP340dYSMuVKCV6
q/Ley7fosmM/V9Pr6EkJIWKeDVmZ4L/13MYKZO0KQ9lw1+41L9mHhvZ9YorT
OII0ggonb3KAvB+f0Q6UGupIEkcWRzy6xMte78tBfcxjbvZKJKfI7biGYgS2
xfNzSaeres1tdUP5XzQLXG2BpfCY2KgonHzDJ1SLajwD/RDJN64cEELe7+1c
AUEtwItXH4mjNQJ/QS30fYo5ypuNjwIUUo/ha1Le5G1/G8Y1wWkVj+HoZzeE
GYcriR+fVkya1az7npoaByKngC9WOmqE0Upm5cd3yBaGq7YTxWd5nxefIzkP
xRwRwDvMao8kk3k7ViZAYQychAeqTBtbzmldWULsyNnfjHQyJUthsUJKGQnJ
Ar8MMqGd6Wk5xqXpuo8EMCx0t6DGNayb8s+74N9FW/nTkZa5whjLCcu0CXFa
wTrn4TzOuv/majrBo/9+kLU5stU2NXNqsUM89rD7GWcXE1P9iuATyKzRDjBC
h+GJn413rN+xz+fXoygoxt4uLX1xlbFRN97BdflqRDsbDaTgghfQEQg14Ruj
hU7jf9DP6bfksnZA8guTwyNOCdsYU3RGZu8XXnRLCIa51S32NTV1GCsCdrEa
+K1wlgC/eIvb6Ic9IAmrX1vlDjemo6QkI7lO2BVoNDpoh36ygiHUMCR8JyWI
4W/1UvkKpz83RDppQyP5U37HcYF6LxT1GSZQiXCkfFLKS5pQmTOGIwTEZiqD
P2DnBuQtalc/0Qe/yw2ONk3iHFejBLSA+3aKHL5EtnlXoK93YGI/BDAQxDIw
1PVqv3VHyaziuPcfvSPoJjg+3Z2boPtkDt8g15SBPx5q8nGbDsUJ6J30fjpg
fZ4Y0mZ99H7AjL0v4swCYH9Bgz0Hf6fCfXXmDj49Bckv5oYffmlQuNk/vpJi
LTN3cRsc2pofMbVQVhi9Mdy5VZay7OfIFITnU2WAzB+AJbuBtZ3+C3wRhiRi
XOE1+J7+WeRUBNFXuuByjje1f8l4YEUC0RV3xPP6MBhkaUpNa6XEXtnhcO58
3fkX0An6I6KvDHvhlLd6qwMKgmXcZP/XynpPxmf2GS4WSFHvydB+8O9KHGJK
XhQHELYEv3ZDglCu4H6Mh2DW4iKw9QC2ZEfLdp5FStGha6wi2WoooLR1Mfqa
sLPNIxpshrKw5nuxmBRxAbcWHLh+vUwAi/oOg2m1hL5/7YWGeMSZanPWNmz3
Ph+DUCwXZdnSMDJtZyubV5vl019bapWTKcZ+lvsp1HgaIMUbB6i34pSR6j2m
f0jqunzGrUfj8QT0mfMWDLgK9KWmWLkaViUeMWQzgkQ8akMsoz/i/ELUPoBM
Tisl3wM6GhUirQ0wD6E1u2lgPh9OQQ+crbkT3Zh70VuFbe3bGFclSWOR7NKQ
f0bzjxPNqJNK0WG3R+Gn4RKVFQPnmkAp8RirAaEF1pVJ0CUk3hMiylYIbX+j
jnVbqX1Ls5sZroh3rsbW/E6F5gvDXuHdWpS/SnpRYPJpcY7sSaOKdVoCo3N8
fVt/pLfxHTIBIvBpS/qj1PO7dZwSJe1RjUa+ok5eFEElvaZt047qeiJQ/OFQ
XgD5gTcYx2N/rnrh7zK3TyU7ry1VOPZiyjWKslHY2MChgMeci+kCuOwsRJHg
+1oialOFVvzb3HcIAW9XKH7NPDb7M3WYx7cHqzs+CYLSnp7JeVfnHiqFEWqK
YwP4WO2qlRgWYZECxReA53OutLEwqYA0QJFocpO2JqLikrPxjIQ7OF9By2EB
QMCxn1tUF6UkJg7CNCrFvJQF0Q8LIFLnZZ5mJwYftaw5Ak9tAdOBdwgA9ZQG
hsABXp9unMOsvbKukrkqvUoYsI+RjhNAPoz/iDBT5IIALoDiLUYqo/Uas+gQ
3Y4b/Ljk+2fi4fHeYfL1kK8AaOOkhZn3L6xs2KmO4UjiJJbQoSyM3SVWvtOB
+Gqh2uOio5gBdAVlp8FiY0S1/zvD74zJKijCum4m64i6n8y2DykoabWaDX+I
zi26Oe2cLxHDG881rzDuNwWYe29ttQZe7Pf1w4TiTm87kymctpK1H9cUpHIO
pXpzAaRMWwy3eR/arJmWYHwdrzrXjp1ueddHW1mmZ4eEv31raxrCZJXEwqAK
tPhtkfbyju9BFm62IV5n7M/OT1wWOnv2xHegBlbMIjrA7USCjfcYHrQErIZs
qH3h7L7QjnSMVqbXSs+LQrkRaHkf7H8s7Wq+xiBby3Ec5ZpRkU1F+/rBEIPB
NUf0IRfmbLLeQRCkJoBTgvlLOQnpAQVijWU99FDenCwnMYYQODYTjF6TARrz
UojnVwSUlDgkNL4pXAjTEVkQDQzgx6YMod1fa+M8j3Jys95HTe8Z2h3WcTET
lLOrzvg1FFjkdozGNyDaXWEXKj/04XOdYBfuWhUxn+GRHXejcJDdjxrl0wpU
LXgl7zV4GFMhz1hyeTfQXcTQTBAFi3tqtKfTluJgzjvuriYQ4rpDlIauHJyZ
/ypyQ4PPF3jm1Pf63eH9qwQtb4IgGZFIlvoRXQR5PaZ+65r+gTr0JXZX16eJ
tjE1KBM4x0AN0Em13aATnY55KXyQd+NJqOo1TLjoZDdQYY9dJ2YJW3U5h3Xr
51tAywWz84Ikt8SzQL9fjiB2HWbBD1SwEjIv2+DZl3NWgP0XSZZpAZRP9hCQ
ve5KYn0dPVHl82jlNnybvHzbowVIRgy581wLLoMI2J7/SS+CpBhqr1VNKLbq
12+6oFJcDt2cA55vzt7ftVr1QIRgNu3fFMF1UUWrbiu3U0Vx/m/N1NvJ7wlP
GZMTQqZMz3Cqg2KHx87yhLj2KWBivNq2QhD5xyXpOiQjSZYu41U7rrSUao7z
ktL/f89Ld0VsnOkxnYnQeIdS99k9hN01+v7iPPBp10WXv8ADuDGQ+2tIab1c
MvO2Jfz1KApPzBqB4LXESJ0ks4D2bytirUAKNwIsI6VgL8sS68M8kjil71y7
kTshSYQ/+FdlmJ8v/joWjYNdT/ReiHHafUqFfigl6RzrGrixdyjIwcM7TbNI
SB0cHCplTUT/3jP/WD8LO5iJ5DruwjylBHDGDRQ9VW5quU/htht1cU3pEW2l
qDLM90fT99sYKmSIRJ2dUur+rmXo803+8QdR0pPCYVcFfr/l5uM8ahov4cIw
hi8NmTtNPNfIbgkZLSBHwzPkC3TVcQ8EesEotoQpJF/KL0IoDdH918s46O56
8OwRkIU6KOiTmzZjCeEquz99QLdxTcS68lp2D0qmZFX1Ltc2IKrSW144A/il
dFcHkSXe2IUyZCd8ZXwAgE+a4FHGiXYydaavqQaQLRLWS6Z0y0Qa3iOPT0lg
Opb4TRe0ABGQ+bXGTtbc2uz5ZHuOEVYH/rpeEF9gJb5paI/nWY9i4eCSE1++
YIuE3mMVD2EK8C6CH57Xj/GYlrbyxSrGKVH9gUsTIyVn6D3ES4RsH9/GobTz
/SBZOmE/FknF5cPNWCBhdiCoSxfYkavjgD7lB3MM2Xwlo/1m+RZQBVbAlsUM
w+7AAezMrHRPf8sEXm1MK7mOsjGLbJnAMRC6+tfK1gc5OxZMM5sZOps1WXRJ
wqSjySWLBbyc7N+WmHIPAH1TlbpjCkgDwzwbZ93/seEK7y2CXItFmNRtN44m
nFtdcySTtO/vZGKaFEJ9T0UGuz/pNkZWxwarHxSWzWbDoLYSii7z5CuwgziI
2vVaVlEVjSQP0R9RaojzutAPe7w+V8bUB4igXtjZ3RiUy0UETjY2TZ5Bqvru
0xzAdoKvE4V/TIAlTTLaNxBQTA2u8b5wwoLzpdZHTsaNNJPMjIp0bI3xWVRx
1ZnwLQ/x4D211NFEqUCfZj1jl7BWwGHDiIV176rxEcxI8oSiy0VxjBzst+Ej
vyFZHwIY/Q8Io7tJDuLzTfqSADxA1J0vI2JfM5rCs7O1IxrFvQI1HCIds0gV
59FskZu1TA0Yr+PWJygiGJEx1qHzpiqzJ7S3dqaRBg/cCpXSKOIDkMIMZGG/
8n0A3EYsUBfnudYOx7TdIHGOIp2hrDy5W9FLWfYo+u45QgS4OLL3NvAXhJIK
KHMErR2wslvdCiWG+53TNC+/hIux18rEFkAGtGySPgY9XgPN+9SR2JMn6IiO
Y7xbNSKWtnZJf6+mqbTCSi4olyIfOu9+KjBxB32Gzhtn+9rCMJREMTuELNT7
UiSqWFpbaE/hwR/EKL8f2HVX/Vkmbo3Vuih9nFElrnOtgkxAskYPJRcGHT6F
rk2qIemX+TbHPbWiNjiBu320O7hAvQQrVgJlr4M3SEK1MazGoDl8oxfKjXcw
z/oSn60Vhj2gHCkicpwSrWLg4iLQ61+d/12kCRc4TYIh3Q/AqjqSPVMizWm7
RooZnZphW3pufdHHhoH7+n8JSNswckxMeLlBuuJw+zTcI+6VeIYhxeuMjy0y
oPlPKuI8Zz8uXdouwDuNxS5BqxJ9O83YNr0IwU+TLXaEBKO443s9Xa7pWHb6
IdqlSydRZWOL0/7RcFr0K0LRQ8+kNh88bwVyIYkSNh51f0WXKghdiugZIYfz
eI1imn4DMYKa1iXCxqtxEZwFGkoS0BCxVlZccat2BYk5xc9okiV3RXTn4twL
BC+VRvDtE99wokF4i1++CWHLNbqCq7E3e7QV4APiTCvJO25gcGlG/efnNp2w
Pdh4V1zT+50ZMX/6+hsjYNHv7UqA/BVUDKIltmvIeNU8hV+ye8Nz531Tc156
ywkXBvUBT1LMUxnlVITeTUNz/2HLvVxEVWHDnXjnvtkHrIkC5Yi6hxzbgSFq
wnrWpAvqKWWFnuPTDaD96Zv8rOJMgnGvn/BMnVEJRZF4G/RCQKy2grvT5w+e
4zT7W7ECLlHId8ctjHPaaTDcp8SOKkr8a0fXVjZq+zmHGuleJJu23rA32N+7
FtRIb/qW5kUTCf8zC09TkSsiFxZnMCJWsKYyWF5xCjhPCozOsBMMVGjMDpKY
Mgt95JbbA1dfYw8zGY0tokz3imdOvf+U7dAwFt8PINRXuOTtAYmEXCKUk3I3
J+6dvuU+H4wERi09aDzOjTBoVu7yc7TjnIBZuE+KhVS7DyWxxZfKB8FSTE/p
iRFMYS2c55+gHL6d5DB0lgbaZwggMh2/iZzlXvb36tgQXjNDDB+s9bNGv8VZ
JNruySdSSFLvRJqd8acal1BC7N6n/pAcYEFn51AfDQdRCC+47V5QZ7vkARQ/
hDyLCCHoFyyv2VD76Io2knTaEY1mhql6ngDZf4NpOl6+x64Ef4n6RzC+tCEF
RvVun4x3D069vLPH4usP73S6B7eSa/DNdZvv6le19S3xfEzkbr+AsM7ibwrf
/EuxsGY//DyHX1SusApD6KNg8zjDLHQWrhXDD2sHM7/SsEwoCNGFWoooyzps
ojjJ6dVV7QThn+KMNPqih4ZZjUQNlseYYnDqLxIwbty1MM7QOoN3avPARGl1
wd/rq9if+D5rleRY0hiY/tMkFYdkiiVVVAXhlvk1REkFNU+/VRQyfiSQ0BgE
N19eJvUB4erUzjgYmPOVfsx7Pjt5tOuNNXG4caDBCGaDwINvgZDiZMZmMh9k
I2a4l56lhHXpR/HyZOtive0UaBI73bIGlGFTPidDQhY8wbourpkAuYhEFdv8
P0WjL37Fqh7z5ofVFV1yhOoaD6Jwr8uhSPTzUKdhfpD1Ge0b4tuiuC+qA4TE
NQ33za2L2e9DJb8twW6QTvTCzRr9WmCtUMsMa+eay8Kl4ViSm3QCPJCVE7H7
F21yVNLNKLH0O+TCjW48H8GMlkp9E9v80o5dns38Dd9tdFuTEj+C26/dh9hc
goeANrp/8nq5xEG963NmzFoU/CqiPxGSJHhR0x5glM+mm8R6JyLdjwz8jZxl
v/aDcvdMaeU1mKvRNu8mTSWXguQTIqpW9H9YERAZv0ezYRTDoAquY2UiAYzn
oSzqFLQIR0z9NWxBaer4pn5Ug+0bne/64etF7PXT1HUN9St1hPMKifbeRTgH
2dzI6gAG1Cp1EJcph+oYRzXaF0LF9Js8wX87RgiuJuO+8brw3YR0rl0Q0m6A
WWbRTl3qkcpQ+GlKhtihBOzS/PfFXntKt4QwlwIhYDvWEoyPHdUL/w3pjRw1
7pR12bNQCzO4MZd5Z1QtKRp5oYroJksRo6CKFhJRNVSlyRlUtm+Eo+9W7gnU
lHZor8+hCSGK1E4UhsEZC09KjKincsF/moIh4YjxoVD4MPYOa7pXk+mfyuNE
12AR3gnv8TtPsxNenwMsCVnyr6H2Qt+AGMLyGwS7LknWyVnP+k5qzn7N8OTs
/Y0vY0jdbd/Uy1XcIcMww2IWc4HC2IOrQ7Nid6tfhDdgq0g2dLV29QdN26Xx
2VbAcmlOcRjattZXu32y9rHzCMQpjNRYTmkyJY0J+W8jn1w3DVnwDQtgFlZA
T4Pzhk4l3S0vVcryKavqqqjZTsqGCxsj06B/jKG+Pe9Rp+4fSINbNslEhdmL
SemWhEAe4fITiwkn1MX4FSQYXCUUb4+IU1NFn6D64rWr6qrgHsI4jj1e9sry
cxyY4KAULaciae0by6D5lf4zBnxeCo2baixsl8Zoh8UAXTTATa0nhz2bj8/k
g+y1C+PkaI/NuzHaAZO4eEdLuSutF1qrxygm3lPKuVGmom2Ag+feG0C7aSxo
NnJ1Kn+JPMsf5sn5Lyq0HRs9zK6gzeNajHHB1FKk6HxGMLvzTJXGHRKnjY8y
R+AdlbGJHWoK3ga69xRVpVcUKZxiCKF8/Jb0lprn8e4I0kvjSZZOedZDVxn0
zuXI2EYy5imSlhPSTSMQK6d//5nynkqJeN7xMfD0hsSxT38nd6k4IilxB8M4
ryKZUw/226znq8U73p2jdqCvjV3tTLMJLXKswjiA1fHTSr/xwuk1OE0kADCF
n2uUh6VGWJlhKoF06FrtG39sSRgOWBdK1BrGaIyLKiRu5GPfK64b6g2VxZWf
i5XPhIqa0K/HrAFFRfjaSvjvXoGqjIrqL+hTBdYPtFweDgCqKoNDtoZTpwxD
Coa3DfeImNwGH9qWHghorIsYxHbc3Jt6/dbAp3psb1L5h8g3eDTYbhWQvZ3O
uD5pxe70UFo2r/5VB/KDARbvy/8+ojZ6IJVIQw3ToFvQwRxUSlG6sTVXUGlM
PFy3yglBTAVynEJcmCxA6BwDOgH/rjEuPenvXwS9d+yzNT/14zKepyDSozLr
Ih/4jKQQM3TLrIPSFGXjLo+1D6EkucCJavghFqqX1DssO/+dUG8tdAr1bZME
p0wwuHkbnLvueHtT/YroHAuHioYQ8m1yeDvDb52izQBrGQ934YIdu3Skrr8q
O6nANLSU0npgt277ApORQQablJO8kdLfFRJD1Y783rFApemSh4aLVXaBVUvE
DohHrmnTmOLFRlO+A1gEpx7L5WAixOD35r3meZQq/j/AGJBN8hhhv22yupce
8WAyGTkusA0p5Elf5dMzrt3i1RLFb4zR9YcdYSvnxBaCv6Uh9TcENmiiWqER
8UIxxlOhsB/kyJY4V0vrlu8FSB6as5xHmc+KJlD0Jv6N5aabqWP+VEJrVed6
UX5wB52FJaxpxSHrB9sXyKR5t43fzQAFGeTfEmn9wUH+ab2npwa27qBQ0Cuo
WgI1tEW/8ozvQGs0enPimlWcKUrS3fR71RXh3941hPrJ9JYxSSxpt10VnvzW
En0lxGy8nPt4iqgANQUOniryZ0SbVX5YZu4nSD/6BPgF+6v323Mma59akpA3
1mO/yQEdIRzsKeoiN4Lo6Z4wsQcKAugFstniEEjM82ND/Lq9FSd4lqi1+7xO
zwiEvjkkg3j47Z7thHAQPWhtbVKIBGdmwPaEfnbJ+2WbCeVcXmoizk8SLcbU
0jiR1En63gtx1bpaMCBN0TCuxuEPW8gfrCBRE97b16dzs1oWZM0nID7MYshd
smCyfkrnpr/1DLyjugIXF7Cy7yabfa8ijnWjbNCC4ETKczkc2npxxcKJzV/S
ZduMA42RAYccWHAquNRET5yYWyKwzYnoWS3LfS7AxSzK0344+abGW53VYHPH
q2lI9CEYOmqR7enpS5EFPci6LRAg0Y4UKLsrtvrlqBE4REoKPSelWe3oSgGR
0M62E8r1pbCNNczHws5/z97BJUpAyIA0yKqepWYm4tf89TH/ZCLVaPe29R5T
jdVPUJKruIw2/5sZKC+GV3aT0pg0vYviSauCJLEuIfNTCuse0HcI2s3exY3a
0cDjYwWhNjfbTFkT37+N74j7uNZK+W4+EJhZ4t8BeOw28m4CHN1PrPSTTplt
MnztYg67CMkdqyIBuMKaclCcP6yS0v1hJwfSAfNKzUM+p+AsYLPtnSkXV1kn
AmpN8XVhqbHKAIleDYWjAAJv8KZom0Le5mtYC4A+nhSwYpVa0AKVXmwpuyuk
3AwVfPAIOE2wzBIS0Wh9yW35hnAFJjEIlzXo9NvSRDOlAm02+0AbFtnOOXfb
SPT+aIAfypQj80oexibB++pfq08ALaIhePgFxSuu7Jt5ODAWDxqOZ1z00Q14
Oghc+DmkjCowyWZXxdi8cgCiXa5TEvf5DIRpC8AJcfb0pF+5GbwOiVcVikMh
O43m291b0IwKkX0Ny5BeQ3/n/wKDTafmKrsiRForazKt0hF4AQGPQVVrW/aE
NdiWyoj7IXw9Qumfas+DmnhMF9Mg2i8w+r/QYFajtHq45pbCE5Oq/kc1SHO6
LTHYyKiOt+wDlEoQougOrOJQDpeQxXqNRPNLBslMuXV0t7ZwILy0uPnQExLT
qutjvSDv80Hjl+EcoDNfBGtZbbIhUAQ9E0nWi6WYEW2P5eXlCkXFbTmPVAfQ
UxN9jLW980bYcYThiAdWh7PO5u/OXQYiFcYilnta/QFPCYs9jM5T5Fe9lWj3
cveur2AxLUlYVqDjv0aXIrFgZT9bVWg6mv4fA4S4AWH5Cs+4MQIVIvp+FIs2
Ltir9xyoAIGRUBVSMRT9K+n/BrXRBuQoHHaDFiIq5i+vT84rONgtZpeAwRtu
iuHZpqqnTaSUMLc1ScJJ4dU05nd2/bZJWxSWgp9pUMfSHbu1u1U+SQ2NO7ez
zrANENv+jy7skCtRnM+bvYmkqiwFldQJGYAPPuZ9SwT8UiWrjMCmqDg8rzCD
8PvESKNDL5MSpJ0yamUIzi5+ZKpFA4Jat/lXPIjP8TtlNqUkDPWJXDABI8rz
NpoE+sXbnSrOCKIqB8RVydAwQFK0id18onDReONJbU/5dlJ8hFmWzsEwabhg
Y4GMRo+0NGOt1BfxuQF3OGua+Dd4QiPM/GTEywlkDBCclFlCwDsm2NywP1/E
+JTuMKGvAyZksbBwaHREnec26Jwwb30J/HMOy1EENrEvXzDDZPV+fmBu1CYj
Z/VOzWC4NgaoMpkjVN5Rg5ozOHl9yNCJmEzNsj5EQulcClo3Dm9utf9lJDQ6
ie8GsOEKqfO2HKUuzkqbz+TEUHRGYLGcmOJejIkUo4uVZteugJmNa6IpqgXA
qkCHS/Mkpz/Jgz8+KBQqlubCekCGbd0peF01xjtDIu7GjGYogno1LSPk3SlM
DCnyXb6bIgw+ldIJqriYejh24qjxMhGkQ7dg0FxcG7a8lxw1WOhh5Imsc5WV
OLti+Qu+xolOog1t+F1QtTqcEeb7U5ZIXhiAVQOtYFnI+YORnyl3kKiMhPmt
MvG2n0X43F2ul1MdUrlaHqi+3Te7aEkKs3LLOEFMORq5yF4zgj323zWyJTSn
t5klIIBB97kAulMblHrsqB5e2ilMnyFO+XFYh4htYAExq4EHoFN3uzRTb/Zc
Gp4c5RPjIueZ/Nby0lOZbcOvzVX4FcgI4jVvfGqfxp3pb4tqEcHo+iWOcXdP
vwAWgzVmiA0NXrtl+0H76qMVTbWn8NLBQl/4IrtxxKrKZ3LEOIaUQTzR7u6e
cM34AeXqvC42wqce1kQAIVRrd3Tx77MMDImnVdBKcCIQ9WX3HAaMbbyhAMj2
MUpCqgQt5+XcjeOloajpq9hH4ctrxCJQcOSUAYEw3IyZPpsRoSx43dRP35+W
7KTtd5fnTTknkHARp0AN/xm8DqCAUH4U28N/Tw9hgg6TksUS/hPbNOna5L8/
LDa5ne7G9x0t7Ydp7tOQAW+yL3ZktDJ6y4Cguixxmv55LXLcW+4v3rXQ+Na9
aaaAbnhGaGduClc0G2FFzd+J7MYvnynAOEGQyMzIS439Yq06CUyPIOFFA9GB
YkR7qr5CSMw9qDkCD3W9K6lYkL/Sle1/z35YzmDUhXWRa45txmVsDZ8rcc2u
K7z8RHVxtwdR/hCR7khY+0Hgaorec5sXS+k06RPxYlLTSI8ugmg6IajfC2ft
ayK5I9VKmNDkQr5kMrjXzix9/KJ9lHnZT28zzk/RVbyMeBJ+dM+3erSRhIOZ
+2KeMUMQAqS5Uu57XVsFFB9KI9faSlTXtJKkdEJrKaw0ENFStzTQSuESmubT
+l9MQYel7iaUuUpfIaWALP/H20vCMceQSm2Xbnn38t5pUnT43am7/Y7kHGwP
/pTUrYanbkRyWr7zlem9JFV1DR11q0Rat8kHwngoNevwfAZqfAIOHSDP6Jm/
/khKdnaCTcbEsZpINL/9VsYlsTnxdkEmRQCqH8trpkDuz3V7cPaTzBxaUT5D
o1e19E3DYA6L7yO+GamzGaq+oIwiJWS2Z21oLFKJMoTTgr2sEjOL1DOO8zry
vYxHILb8ISSOF7ji3jh5JynqEcP05jkLXxfxJ01skNMfOKmubOtmxZfEXwfg
f2IX7xi8gyO5ji3cFlhoghr05wbpM9wgAcj4RNKoK2AKLpBnM4kan3lLx3cO
BnIv4eMmpbZanThvbO1HFbbhmtO18TDC5v/+PmE8w/VaynfrLHpzm+jwUdCL
bIjNHDSAkv4qryEjYIbiqXzTmXNGA1OJSQywrn+9YPib4/yUux5zT4Hrr1w4
JV5Dl0JUuDRNsGP9Bvkm0SqvMeZQvGUJ5sgAJg5zSjjbqsdwJBAfYokGNqCU
eiwyXq7qfWGo/TVLZDWjDUb+ry2MZ93WJLcMDUl7qVuRoDwMXZOx9kMCw1Sh
dc63tAc6gkFq3MIybxW56ajjyiBliRLdhlfg9mhF9IyA9fiNmoc40yi5xH5z
uaVlgTFyfFr9fVUtiBneHUcr1OUdwu0DmvY1iYIr9suD9fMaNSLcsy0SzjcJ
hGSu1nM+7ZwqzFWJvBEfmnNBuetBlaXlDx/x+0SsHnDP1cNpXbv1t2QB6a8d
sglKPHvvo49GXKTUs/JHubOfRSZYT5AHhgo0VTHI+TWfZbiO2NjCt70MvVac
qXTrY21odI0yJNMF9LNP2Aku0e1gdvMeaKJnb/fTpJayeeJ2shHCMJfEJrNy
C1HxwkHtc+YTFp1bF9RGh7XS50YRYwdd7tmKpdteLt5F9BniCTBKLDEjD2Hy
7fORqguDeOZtUfm9GT2aNpFMSY1AvZdHIKVdCMes/3Fc20kGT14QTmobziFa
L5fccsMOSdjYRJSEy2vLEnfhDiPa0cb6sEe3JkRCzNQ+JgiCrPPqExVExIWF
HHakC4qKbIrs31GVQ6iI8BPv9t1yMQramsUWXlZA9Hr7LDvsY0r2qtR72bPU
EfPSzdgiHCP0yIRLS83gDs++/x+RWiD6/HrK6UsyYUFX1VAaSrvMdhgx1cDh
abA4ACQWuICSrvHvlbhpTvT+KAz0EJxWF5Br3TXZ2KCUIvpyaf7cgyHlIBu0
7i1kE1R0HbgdgAJ4kEUrqM+L/kO/m3wZco8SNBIgrwZEdsF1HVCXV7MPXd44
b5wE8e2qxdTliiDpdBA0jx2B/slKvOIIBm+ZSUqbMBLUucyMniPrJZXK4lGQ
3cr9mHMl6GDDgmjJccC31sFFHW++Ck1H9MWcTKBf233z/dkIb78m8mdgIoqY
Lt3vdpdZTPDOldT/K1wsCTj6f2nwPWs0S0Ov/6/Be3wPa76qzOZInscMiLv9
9AGjsOqKnT6MeeKsowMn6ptOebANflhPbf26UJU5JkDwU3pW5LJq/zs3PogA
oPJN5FoN6LPFJctFrNP9xzD3nbLAfFyZdxiqy2XqkN8ar6qVELt/JRYXz8OF
BkNC0j2dBIZ4M+tlNR6OcgcR5garCnA8rw/rTGoHAbxoA9I5USDGJv3F6RAt
vH6Y1gySiH6tcqw9clELthwVkWpCCVF4SUB5bvcGt2NmK/l3GR4Sh07M7TWD
aqeLfly6ewymClEN2vLi0WYv1JJzgp9nGSPhpuS+eRGrHhisv+D7Ef1ePTxi
kHC/9ReqieU9LdK2Wl9R73AT2KcOrc6rM+KUUC9zJOP8NVwC2r46Rd1W7Tb4
cuDiz7E3T6a1eRRCA8EgobaxJmaM9JYEkK/tTx9F+wCOqJBrG13Kn6BKo8TU
4ifhDec+nesh5NkYadCgV5YLEZnI2GUEKk/jCKs9SfXmAsDyUDMfIk17T7ME
oh3vSWfglZBQatJPoDfEOu1+m3EAle7gRGFdWCgOQEwLvUwbEqeJKZPpB2Qm
2aUp2iX5NY2cBoTOSj+RVsEBO6AQythsXpf47CBgq0gRXDUf6/cp25+XT+Cz
LJH4qD1iaQ4q+HeKLNNavu17z1BWA56oOZAIue3xceVc9P6tv9y3xpAo7nYc
q4zRAnKCXc2BJ/mArHLbnzfnfhUBS4qEeA89GHIiPUeiY52uwQ0O8Lpm3ZJS
O2CTbqvbuXr1PxTEgFW6xdpdSV02teKrC/UoOQ2M9v8MQ8IQgG4NwqLIdMLR
gWhY+dFu/4UjLLV6rQXbkaQwLnmX4h/DqJDR/HkjaGccqXSpsG0SrnEfEN57
/OfuHGDXmWAbBN/kgaUkeoceiWOoRyHl27pPaoL4hLDd2h60x2JIlZsWm98U
1xvMMw2Pepwioz5LAtoI8yanWCl1XNpa9/6uQdRifciShosj9l3jUgohCScg
kzUUnQifYscSIobGFUnQY3IhSejdKai9l+kRBQoVXENMLghyyDUh798+1SQt
sAMt9jnC6fEhgatozoSp1CF0/v9K2M7iAvjHhV9d7pw+cqnEs1+GSHVTx2Xy
XhqkiCyfu+0Us2BNNZjmtQSBevaSgEccGXtJFBFhNMw2lpRY1XLvZqHpAQ8m
2es0mTtrVyIXHdrC5LYr+N02ZLucS23za9XxXj/06kTbMwm4kAvQCJrLFXkM
EB42SofiPubqT811F2JMA4tEPBUkKzn/BgTXRMwAfQuS5qH6gWnif1baf6h1
cj1Ed/l3jRsgcEcXy8zFIxuBg3lYLa8ITThWjOVYvdYTmglaaPBJbYKklNWW
0inGwyo8ED83M3tvPLjKHbetkVJsKUfv69/uWMm65x9o1sfcvVYnHTveYu8F
vgMZpYGSqZpqEHSF4fQMQALnJsVE7pq7zUn00q8iGUCSkab9OMmV7kFaHF3D
BWxZe8AG1ImFB7UThaHYthCZevPd3dLDSm9oUW9bzqNy2qoz4hlA8zT6vQyH
yCs7PXB+QcDiY7e7eUqQyt6w+gc5j/so8ZFYger5JBlBjDkqVnJBqM64hVl8
7mtpkqUMtZ9iwZhH4UMwyB7LUWM4pzFdsDUqu6NjGAcr+XhQpmK33unfC1Nx
MfIFzzXfAMQBrmQy0dXfPgA3akmgnhKTUKd8dI3W32KIGMfwX31lstQUH3oY
o1AcEZlf18ypsbw4+3VvJBjGzTkw3W3+uCzj4WbiJSNtxnFQJOIlbq4RMx1t
y+tEFv67rcHOVjfaCg6o2sRnVtGorxdFIwO/8T8/17dNAkRW0Zb/5UcrJDPW
ZfYcTRgOGFZWjSkfS4qdlP1KbhJ4y0VtgdqDUoOg6KuKJF30csuPuJxreA/K
XD/5SOmt8d5YSDc42Y8LjHAst7vBXCSYKvacI/Bah1oioJDxXpVNKyDKU12n
V5ZdCRRD9UPg5vGGcXBGoUM5SptL8RQBC5d2SrDFufBVV+p5TWwoDvGSPrDj
3HePNOHg8quT/rNcf0xZ21rDDSNXcGkAivYEEh7pnvMC8fynxWL3HqmzBiQ+
VInDEsRhDziJf3XL15pj0nrRyQIMTek+hjR4B0++fT6+ZhaAP00y2JbbOGba
1aR+dCKHpmxLXWQOQeDUZa2tgfidbn+3c7VZc6p6FMEzF7rQR2zxy+JQ1Bak
mK19+2HTDO4ERfFKtSDowxusrhuyyslCnaA32ArGwEgz5jtMIJHfonxPxCfx
KY0MLfvXEPiILGwd/8Uubh14jTU/Y1MeMZ2GclApqffbaJB4yExuXvNtg2XR
8ZA7BWeoDGWrroH5qKLmIixGpljMDT3j4Cy/vLJPEcVW5SFKLlcoSavhly3n
IEZqVMkCYfkKxCqTYUubArhBtqT8R9FQxjXiSrqkb89bhgL3bHfHu7I/nnlK
6yhqdj57EjFAeid+/Sa+J68TTJhk5QoNxGk8qLo5goXPrciNd8TYPAOPuGEg
cUVMqI1aJ2GM468sqbJFRk+0hFyvRruL0rD9ltghruS9Ps8AI3q4LYtR3qCN
+vtp84oAS/CkaYLdfIM4DOicidPOIvYRwFgDvJc9g2bGWkWhJDKRhcrYSjOY
Y9XPIuXpNwjgAcPcdbcekKz2OEVzDsip/UslLFo3tEwj759q/laxqNkfNKwZ
KqaLpGzMCXzWTAqcmZPxK1mx41yLbNUqKUyRmTExfNkoBym6f8x3jieHomT2
os/d+jTCM/N5O1DkVLsdH8+FlTUiu8rmCmNlch9Ru//1fCyTmRPHarZI3Ev3
TzjMMSRcF7BqURKHcDkca0J0YAnB6B16ktPoRIeCqdXWbP5gGSiWNMhyVYXi
Z5Wr+iHwjnc/3zo5QZs2QRL9027zoGT5DXLO7NA8wd75KlP2G9RjuTsfg+oU
5qsrTvGoebC6WN5GcaHWS9r8yCcPqosRWaDgrbggqnPCBdTEnH8uUBXGaAf3
HpslZMmCI7L6Qeggx8SulA81yItiiLjtHL691SBJP6ARTlEo77qQARERUFtT
/c/G9CqTXFGPvy1y2I9r8dwQT4N+DW6zHznVycgkHUL4dkniq9NsuBIL6bgW
2uQ8mgNn8s4mTkLirULJfdirlqdAfk0TtEwOrfDsU9tkzHHJIV4XH9ZqCtZr
LrOc78BT2VxVHf0XJWE1HHptjLQTLQYw8nGObIFOm+AHGPTYyoFGbrRPyLre
KinSAewOMMj6rM4PpWDB4fYSuqUZhujdoSRO9dot5ahuVMXIS77gSwNxT9q4
d6YbrrbArBlvBlxT48YQt4ukHddcuvccBFccOfL3oT0JwvC+79PHY9sgbGGG
EYIOcmPGKK/veH1JXirKqmd6bPL9GsQcQ8Bp/z8dzix5LIylJ++YzWfdj/Nj
rGg7VwgxTPH8/4Irk8CohrJcHyXQ0ljFpwnpHCNvcZl4dUnrsF278hkrtG2s
aj/EPNkSbce/Dw8OxtVdp3SYh6Wu4APTl9H/SYXBO9z1p9C6t57ZqyNsaglL
053TECg7hU38AsfKXltb53a77BzvJTmWYLMPDfRSQ9BeQgglvIUFxxJLVaG9
2IsfQgQJ+WLc1ikfAB4IfNPpNax/GCjHw9X5K8J29EBBBuRgIgHKxn5LRmy2
gN0Bv7r5H/QAr/PsvYIKJ97UPmp1ABVQh2qQ403OFLupyWYjwXRdBtNvr0E2
5WcvFGsFPrZFD6pPrM7cOi040C2XhWuNL7dF+KnjJRuG3VshGZnFj++AO2gl
Yrb/hMU2g1A4oywh/inDmBZbeuNcrW8fY+wST+lwFxMTifymaIjOJGKUu81b
ASH64botwU22RJAb78zFoCMOBsWCyc+7wWNyx7BajmAeUWUZ5mPsTRmN79/7
K/qqU/h2jwhT/E+t6ewonTMirEStUF6MAqs5AdUqkmGNA7P1+dj4oX1E+o+t
g4KarFRPS/nZOiXUETEJdXeysLPWmM8KNFbkRqB7tqR4cXsGWmHAiEyGRTLz
gWGJMQzfHZ6N+4zyBeQ75NMVBCR5tBfbVYyTFG2ZdyOmGnE27JvUeSLLgBpt
QVmOh0+LBJh9yz0tvEDBe1Oes7JsTqSQoLbhFG/NrExfNuNk4+Qw4YkJe4xI
SqeGcNkJNL2kDv0dZP3MPLmvY3Rlka6kqJolVhVtg6nJon050x/s1oHlXm0E
TcwVgkEeJzuWUVzfHUVk35H+o+UmAJAaBZpqiG9ABxo3knoXDVw7Z+XOBgcU
fvlzXLqT0UY0Vf8WM3AoKJXNdDY8UklXDF/uAzcpi2aXOiXpr+xVJatByZRf
/liyKfji2fLNm9qX2Mm26ns2ItcqSm6fKa2qZBmZbOxTRNWcO07v5kTJ1AUr
XDp6avRUoAvIE4ZJ2tziLV/Z9c3PZOOtzDe6HAbIk7h3tT014P1NCAh3dMJ1
FbOrZw+SrMYpUbtwxEIQ2gt6GkhBAX7gflBLJvk3njd8XmNDU6usiD3E1E9n
OTL4KlRIGawMgGWJa+IXaoCDFD8HWlQ/xb60SNMYQOOXXPjsNyvc1aTvu8yc
fRlg/DOIlppdwVzkib1JDgRTal9JnsGqt39AmHgw8pmfqpZDZF4hJCnK+WAv
Pq08LPMQmkj8XfB702PBparLOPOBSGxP3FrmwQ1vyv0w0HUB/5qpe2DlZgaP
GoEYGyMNDHNC6Qs/8kgYIaSIw1aeCB6CmRyYvwbZMdOv5aKs1Jio1Pit/SSY
3zqopanOzTYHcq1UgIZje/WlqVoQEVCwQ9LopJ3q8Ufhftwd9BQGp+CI8URH
sYy5Rt0bk+5GgBGrVzfX7/9wG5QJhXJJhct2w47BzPNmP97HPC145O1yOFd3
NP/iT4A8hpsuiqIYe3WGejR1lpfC9YJxhrOT/R055WiZFdQygoF6OCF++C/o
4KmtBSsXvJ38ij23Xcma4E2eql/A1CNMcxfgP90CMsh3XJ8J6hSpukUkzAda
JJb+zwJvNMMgtGys5tONf/b7DSFDW/TzshBQdR6iZLni19pGnAlHyP3w8f76
0tkhQ+x+u18E8lWmlKt6pbHLK7ZvAU0j9dNlznqlpwFQkQJjDdBB52wOT80a
w9IVuv8+58c/+/ruvRxw9O0DmS6fKMbq2WsKtpRmCe01aIiYppIHobkBmZ9/
8fVUT55X0nrlGsK9JrRF4PUprrcyyk8emES8QzF3Nud0QpP687wkb/g0MCE0
9spKYxaEvfYAZmpEq1lzrwK5Ogw+7ddlD2XGGPXeczn0VtTDw9garFgFajZb
4604iYha8IGvSfJc1r5JS6ttXKYh2DW/NKc6CXeEVYZnAWlVdaE6DhWn5Unt
KEGGigKy6OQANt9ZOsGD6GVGiRzRIkcTPNliTcFeuMKlgZneCXPm/8s2e9+N
zNodHab21SJOkZy3kDFHoHAXwFy4c/iJc0NyUOc5YLS4yWyzOUZqN8egzABh
7Viez/AQe6JXyv+MFcO9MYUWrNreCgj4tajJFvv8FjKJnqU3JRjmlHntIIsc
NMryg0tKmLmt5bVuzvzWFcYjTAorXBflS+EIa9U3wrPV95b9I/zfkxrMMY8/
RjgXNNPXr1nm7eagIvYbdcGGDJQL7l6j1ANBJimSbgEK+crxIs6r4fqAbERF
srhHZqRuHWBRc9hDu4ATMw4nfRLWSdcWbeJT7L4vNDXBSSNfN9cyHZhsOCyX
TsrX95hazpj+qONDRIm25xl94Z7PGxk49pZ+QnuQFe8W5wchxqeYJebZ70l9
hhWceqmtFaWyKM2OduTNu9TRo9tYBM2Q9QmdTK1XQ1nvFxkrD+neJ0w12ZTF
uteawFPNeB3BMYlMcgVb3A+xM0l/2vZZh2aK0zfSRGlpM+cPe5ytJZ9/TAjp
pJnOm+nonPyLZWmAioPJeNgP0SiUMCC+6/yJT3xWEawkYxrKqzd3Bkd8B+i5
6j3YTi7WOg5GZqB4N9YdqzFdePTBZjoAifD1Jco/6ZwFAkBp6kooOiLy8c3w
wTe55pyOcdcShbW11GyixRmp2XC757gZpyykKZq1ozfzeY/lZU+WAVr63DbN
nPIAOiM4lRFYQkiIMXtCkvDy0J2e06QaiUSmC5bHyy34neJ4J1bXn7/LEmbf
1Yw0SGR2Bse7m21vR6w9fatpBlVCnVnSpJnKGhzM4C/UStzl/BdINkHUM3Xv
ujyHcS9ohbevQpAmqY3lTQ+oV5HmV8dVrLy/K5eBfeiHv0Fn5ymhK+Dc5ROw
hWmd88X3Yh1b8g5jt2eSWnogmvhpxMoCcrUgVU1Bwbk9MSNCPF+ZKShqw7bc
rB55i9QGZhyeshqfmMfBmdSBUje9caJrVKPMpXsJ5zHAhTsRD4iFwHtvXOFn
v6NwAriRxVKfyIa/60f3zGjwCZ4Ube0Mw/qmNntdaZY4sg9jt5WVkIOPDSXK
wZ9XL2kdbQw2fmj8QyeBcrmRgLusu0ZSpd+GPtc1CPEUs479ZTecEGVbESvr
CdWrOK0X/EIMOnlUqYlXRWtE5qGMjxTbEOV7DkApQBzWpEq6+gk+PkVcA+aq
vpvKrVULHV/EgUsSEh+IGcCY1ijbsDv86Lkp9aYJ/NpT+Y4W0MVCQuwd0l4H
fjgFG8kbIN5SQcxRHl70122RMZ/e8H3KrXi9kHV1qftoTrTAfVl1dZOKU0K0
ljHrZPgi8ohatf4+DLO+2Dpa3VazpBK75jTSsRKIDY0skAq2mCKuhQ9eaHPH
aZH9aiiAExFOm6D50SpV3hsqJ+EibVvnotBSl0frfN5ZBlrf8OCgCjRaWF9X
/91ZQSGfAltgwGbRHgavP2BCE54ETI7m5sgINr4/J7FuK74rOPPHoZ/RDKaj
MSw1l1P/4Mb99vfCD9fGA1Jzc3YNn7z8AL4d1HGRqHbYCRzpdxDquEFcpRIk
XbF9iFSHNypTTwtS+xhP/4CXX+99eNDu2aSgEGHE1RagPJScOtrh5KbSmlTM
wUpInjM05QzUn5LKSagZ1hvdtxMzpYU2OsGBdvt34YrkE2kOLiUW7qJXpL/Q
umCP1YwzV4chGx44OEjx+xeEjpdmt+H4AnoU5peLihypFC4YiYx1np+F1pdL
TylSmva8JacWIOsZQc3s0RjIiL0voSttIFbbm36ixYuDYErAa/pfS8+zO0X4
gWFw1e1XKaiJQtIV9frVbGzqNZe2WX+py18c+mNZMV96Y93LYoUwv53//S9g
eYdmgT6AswWDtJJ+taj+oq/QJfet8vzfvbdI1mkd7YdejQxI0py76CYoBu8z
rxq9bS+KwDTAd5OoSD72RRhgDaMVC1JuUJM8fHRZmtNTWplmZKmyc3UYqGXw
TVmXFsiIAhvxtp5Rpmr5t9Zp8vhKAjIbGc0nyZiuS4nkrm+3YU4zbZUmWb1n
WENKl2lO86WjXfCq1HOJftEpizqM4/KiApIG+fx7pXX/NqUs8P3b5c+5TENV
YHfKMyAxfvVMVBcVkHDr/JipXUH9u6P1DZNqpuxLehsKJ0eiJPwdSao9LeWW
oY83+gJSsFf605jVl3ueJ8E+IeXSUZoppvHq1bnMsSFJs1rCMOccpJNH0PZ8
IXMNfe1iLkvEGjxgOQEB67Y1siK38P0jQkNrf8JNBBp7+/YTYA6vPwuo0Qqf
0NFR4Ex13JlJLeydQWLOTLwJChQgW5bC6avTpHVFlv+R1zjSOFylhYg2wHCt
vDMShjIdJFBIaPQp/xBIbeoBxvMQeRT2VBQYpb/iZmOV6RSVO1rOnspaYgTh
Fyd+wgcWSDuXsLDSZAsW6GVFlrStgobuuX83cV/pIK7HbRVXIkfB5I1zEGHM
oP/kvwaTT5+hIvnDCZLZFcBrADkrVwjjL3XJpopkxTQTqvOvXyUcupK8LBMo
U3Ugy8pPeqdXxW6gSPZRZKq98DfiPoptqZo1BdDZGDRLTihDQgaO1ijFJU4P
64gySd8vnOUa28lKGHQ4BRNgz/MO80e634E1qjMjsnzUfjIgona2flx1Dx30
9Gt/Y6IaYpA9W6D9jqkc2Bczi26wyz+XYugBYAQojhwJri12/YkeOR1clA2E
cOFxhjJqqxWM6rnZTgU5lloigjzjSFt5dTo4aqNRhPvW5AS4U3PPCutEjeSO
n8oaHig7etL7VrRPvnuUTPXTpxt2spGLZ1cvbi0ULeDBCrCkpmkiaG0LDIIh
+QPTUEKcXslHJb3xZtri9OcNDMSOXshN+NvDyLpTjwNJ5K4C4dquVjJ4OKDx
CEoBW+SiasJYvEBPbm2pesatmGkC+JlRnrsMiXZdfgABm7FnHdQ6qZNt9GKN
IbIqNPY8Hvq35ujsiEOElhpVH3tYwXsF1mlgflwDwNK6rtRYvVF1ABE1UavY
xhVe9qHtFHGBjIyYrVuXAzmfBEjvrIZE7+C/GOYYue1+5g+Kl5rxESVZo4Z4
K02KJ+MXgMVlhI7qwWNyvyavPIWtyb2KO9qo9xWyzaydVj4jh+wxWabo5COA
tivgveteLVkqSRmPoaHso0T2flm/YE3TWbbIz3LUljhExMuUJ76htL0jX5PS
pf+AjerAt1ml5yilkciWYt8M/dwEZFKeUUkYJEb5JLfAxBp0u06B/Mwxx6iU
LKqpmbQSuzqfAL4yJ2JTf7R6Pl1uTFTaqkVLdYcADygBaXvDF1MJA8n4mWPs
4opaPFS/wGDn9/WKRoNWiH9pGyDsVd7oPGh7Rr/ofEFuKUxBeIGizfsvFVt4
LXlOYUjHnshCCh2Hi6NqNK96SvPOd1VYjn8dKAHOBgYyjyWJaRoDmzhXgWQl
bIezrq0Rnh+FKL8I5J++1SIZ3Kr5Z2zm5RP8rPv4lPhIfunktF2Ho69uoADS
TNPW73AIUQdordKjcxfDrCMJHh5UQ6EoneQVjNe3Uh6KplJQEznSm4Yxe/nk
0jzNCU1uO8El6Q5+AboQot01wMS9z+jr7p/ULIpBaeqOEIe8h3t3mBwVQHil
ajDY4nZJxX7xuxNC/XApk2FzYO6mV4aenN/ISaLjueEBdHUWdnE68tVnONJ8
5pnG+n8zDuAoO2QCT5aQ9mje6Em9SD+jbG/J6bFVXzfsnUjHSc08ZEype4Jv
4YbMxSktsYM0Gk1j1WkNK8dLgLptuQkqPVl0r4tN3vVfDjqjgjPtAnvh+hJ7
JFW5Jqi6iR8V4qh6BW1x69I221XZDI2/iUiV4vzAOZLJ35DA0FmMv3/5nC1y
76K7ITDJ5L30k754yQaLqgy/xvlNQHhNhwwT/p9zhRjnbUusmxskXB72agKg
/mAF0RcpH6/PqGcASri1W09q5qQTtfKudFQFevI3qdc5fKssGvb7M74aj6l3
WfdB0svjoXpRpWP7GOrABPbqtWSMWHTYSqnQUnM3WwyCidiZ11Iga8kotXQ6
DUOq9qarroiPUqcfvIFDSRWxpusuD14rqbCJj74kFW/ga1HBnwk1J1UxywrD
dtSxImvabfg3HJFlj+tu0BbaBVhkBxOrHlO5jPEcKuUnZo8AtUS8aJpXCmTQ
hJSIuRVFZOzfpRjvVEd/KmElitPr7CkNdzkgc+fGiR8kTeQitTFersd8jiTS
kyfYJ8IGPf4kW565qbD3kjxg36cLjm28t2GVF6VqR9u10bHdkdGdZssBECvW
jJE6eoDp3TTqlSNpBcAWGckHoHb0aeCrMHDsfsENlmpJuX0nzL6OIAk8QfTc
18jno0y0UKUwk3qFxLOnfLKIKHKxCRdJ3nmg9s0WJE/8kHR5ACixUGWQYtlt
roSwh/ApJP878JG83g3Kyk1RDUGC6QScsrxVbJ2vvGpaEhFqNgh0f1zA7n9d
CmMe3cNC6PDjxl+QEcq7lXaV2LvhVadfplFmAWRyZ7gQ7I1pHwCw+DsWYttK
dXnp+YpCCF/20BjLBOXGVO4LfkKnBwPWKHr7l/yje70c7JYX+yUoAac1Ny+M
W5JogSJr18UQY3rCqyeibifLUsiRn5ZV/EC6uHR8FpEMoXcU6VvSetgWzCV0
iBV5uhNuGcnZOWqtPrbqNQuv9hrD4EghXsRqFTYU5oioRmdiVbck4Vd/P/n6
Ux316tyFDYUp9WaB/Bfq8DEDC0Ijx2ASuk+6MLZpK84hMSUCzwCAZR9/0dJp
F5M2m67YFr3Z7yHrdQ0jcu4CJNFYafzxWtx+05YS0s5JBla/D3GaAd//+x7+
xNCYW/i6/mb4dyEdGgPwMZSouLzWFKPSOn9IxrG4JVOCpLWUiVpsBHw2RaKD
NRVFlEbr7G4+VtMdFvDDgvX6vCZ8PHy+wvFGS4PGT2Hozu3NNALKGNFBx4vY
f2jU46Jzl4uJlO+IL5toYMGOf8ygOwnceLlnUnNeKVjGMxRg1c8T85zbigV7
voM0Tksab7aB3vW1dJHtHBa4/IgybGfpgz6AAWtKjfLroe35/5Oj0Xtm8IVL
v+pNb4L3cCs7zklr+SNdJh/18kFKZAiPvf0vAk0/3izHMq48BqWs3We8sFKu
+OFv4sOXcutTi4KR3OG84E8aErSuqVZGOWQS1qFw0rALDBa96UVS7qH/Cy20
Hlml+F68Za+wcFICeCSwLb/PnJv9lH4aORgB5EhR7h9Znjf34ueHCh5fIKJh
blrWO7jQrYqC8eVs1haRdeBki3XgcZFYvW0JnUz2taNI+olvk5cSFajbAD2B
2GQrZkkGW98t4ypIDLySytvd3WKVWAdfu1cqvpGPoZYQkamIS4p9q3GD741P
dJzwPl5mfZ5/GL9Gk7MvojRcJcKTAjS24XxtcZvZviJQmAqz8QTmuoYdw1CU
CWHheVuvgGA93kruTZjcY+fJjC3gqHTA0I80T2mlhloDc812oKf7DbS/4S5A
FAmFoJSaOSRuxnsPoC4xXBwQSN8/dK6o0tI5Sm18XUdBZ1TKL6IpGIjclzOB
Es0Qc9dbeoE8LfaeQC1SffvQNYZTYTB6NMgqKnDHyh4PIPp/GUsz0xRGJcqF
pZt4/qT1KbLyx6fsDp6RwC/d+zgLLgMwewCrsFgElAvpsU7f49HydMlPA/Wi
FoGN82YZqDXZeRBYvsuYhfWteFTCaBkc4LCDtw2dta4zfizZevfybViZAniJ
I2dDRdN075qSKTQeWu50b7MW1PuP3oAm1kHp1qHCN0HPkAh96q1nH/SzQXJk
9qZSQF7c7/5JZuoqKGf+AadcMC4PVHugEEyWXBjzTeGgt6go/8y4qXA61WwS
+FrcR45cJLo/cKBpjL+jHx0N6wvc+yxyfwrKtbszYoTsk48I70cFVo+Xv5A3
HaleplhLYcHCkkFDJcQKU6i7gZmqjuaGaeCDmWxPZPSZTcOTsfoEziIqZrnS
J4IdIUsAQDqa0IU27VUJTuwG7IyHgu9VW4yiI16+P4edsJgVW6edIOcoXy8B
k3ZQjV6+GccWxuHodZgI8Vq9qjYvXBdprXjpppNpQMwFZTem9bRV30hKRU1a
/0RBkYPXdk14GmpbBzFBF4akgGDUp3Iyw/VFxB/2XRbIOrOpMIlFwpZZYqnB
ZU4FJKkqw7e4gmWH3YUIuxZqx5CVLjHozK9xU5syUvfZAuI5v9yCIRmgApQf
1ejQ5pPGzUUUcpkcjhPs0C/eE6MvvrVTandQFFTkhxpWcgCkTIIUtJO0zpN1
HyC2KhgxNZiEyMkbcf0P6Vy3jf4Q8G156ed5mRhxndW9ClT0hU9+VtMLSChH
bMqK41qPtdTzp/oaOQpmkj463H33ze/2lad9fz50V18N4CzA0dspZPsSy4lh
a7p94DLaf2agu+9wC+7/tzLFsVaG8BDOjqQc07vZ3VNh8/nJ/O1/0jRIqrxB
B4ASC2R/F5RY4pKx9a2DCVTQoOIDX90L9dW651IAVs75UsukpQPnIJOOl5Ku
Btjmkr9memyYwso8y40PmXn45nHZ19VAcFnHiitmfpSU0lFI8QZz2brQ8uk0
g5iuV4YcNv12CizoGkZonAbF/gt511hDN5GZAogZzR8Z5pVULc/Nx9DTOYL4
NeFOGC9eGasvb6Z9D/egrQRePFyp9znFs/Pc4SAjG7kX84PItux0Kjzl9VZZ
6wL3UNR6uD8uvvot8lSm/dW0/hrMUI0ToSlNQrFlQgaI2T7DZuonKmRHGkDb
IkTj05jv9EXzbt42Ssp2Z0KlVC5hgdwltre+lKOJjcfDsE1T4HqEU4vp6D9E
0p8U3kywPOsdbq2lY2wVpWO+R1E9ZQyyCdS9tOPmNY9TPXp2MF1UjRE7e8dL
d/IxelBpfGso8ruxZk21EMVeixTVv52Y+Kb7JAtYS5eo4K+BxcLl0m3yyJ8X
b8mkledscbwS+Qqn2ZCV/x5mp+JXy6AeqXQzA29JLlxIYdUXNw5othySaB2U
hhj1pAufrN6n1XKN9qQl6JbWetAflmF8KrADtpwNPmV+GcYDN6Dp1n85fS4y
XwHJlaAd4bfMU18GJJR69f+wDRYRii/81MBoCx+ijLks6jDtnrhW9vsrFCu+
tXq/6wcWSigLzpbN3HZsRn2BLoQepZYG+4P4Zr3JdU33ZVwMO1Saf9+fHN9w
Y3Oo9Og/KiEahyJbkwM785NIftIAMT90CPuTAHphXThxD651K1usS3zcDJLF
v/AAEwcVArnN5mJ6QdhHDysW24TOH9+oqngHnGqdhgvEGTxxp8Boi2NiNaWp
8ShilaI7wttneKoNE1ZsVX0wDSVP+8ibfMtOWJfy8ctTcBZxodrvjGkdiqLi
b246bIc1xHLTIy+gNlUb3xoJzGd2a2+ghnaISaXBBHyyhePZKi68eDZH8nUb
8YW2qP1pJ9nWvkll91NqICCSPey/R/vjdq2h+EbdRuCmxIR2+tl28fyy6aiI
gBF8NEY/Z5Zt8YkeJ/qHLacTdOcWyDfG5XQIsDpJ5pWKf0apW7hmAIf2DqIH
cmrmCFDMzKkZgoPWUCl3jvm+ARPmF3tnnXFkt4zkLE0xEAtURRgCf99Ojm0i
OfuZcXqCLX6r/okZTCoRQ4pe0WLgUGzjZnlZdJ/qmK8aMOk+uMaUyy3X+myN
+U0HbTa/2J3t+kyFns1+phymBqpSEIFs9VlNWL3+6cYUkziM18C7fSRlpj5u
BbK2PKsfilatbK6GVOBGb5l6l/yrfgsRaGxpf6hi28430F/oRurjW0AECIGt
3frQXIhhS2frRFcOMAo/2O44wah85o5ZTf0BMRgDw5RwgCz33TViQJLYbCy2
oabNoNdDxCXCDyn2XtlqlYE6eIk+UpuSBALYGqBJCrqWEK9eMNnGVzMwJXdy
U6fVS800agOz+mz+PkZrY20/Oov4B4AtjHBEsB6RvFjZTmr6LD5veRjuTH1m
3oYdS9mboX90LbIipRXtUNf6h6pbO+oBvxsj4srmVuOGZ4bhOBjYdV1o264Y
A74XQY3xvGVsMu0nMxHuvjfgPr1Gl80InFHA/lgHGwPDK7CdaXodR3f3n8V1
DBNeE3rkbRXQdYkrPubW5YfLuDb+205C3jTblIaT/jNnXPY2hVSOCGxmKuup
ilvHeX21gn6pGzdlhpiK4TeVGShgwYzQ2FgrwQwPW9e5cViX0DHlgmOg1pO5
waIfiTKyEkX9phP3xv+xJn7gZvkaZDob0jhe8quFrT1iV7AK20bvw17biBKx
OPDQNvNgp0Lp7Keknx2vUgLzFJL4YSVkXRhm9UwqRr34GcYfaaPqcfhTDFLd
6bJ0wJ7sFLLNKttZyBMXeD0MZB789u2gr58Aj/OXTUuHpGVQuoxCoXdALgEp
6H5tM7rfVTpGqtM1xzvKunsspsR5aH5tGpKaJBIQJI4VDLbFSluSjdylnYgM
m3AW9QJkrO0pa5iz/LVQ4mAVaWT0oTNwPF0Xlcz4bV54+QeMVN7uOaIYWSSv
zZmDsi1hosl1/xFXheOXkCg7Z6Nr0ZKLTSN/8Hg9XrVVDhm1PkW5tR+HrEf0
jYInNR4XUT6EkmDzOl0/acNDxDl4+7GWB+GiN7UuBpaLi2Rj9Xng+f3wkx/p
34YicfAY7jl7M+mU3G/6X+4BHLshSWmTifRUeSBNRAqcdeIZvjaH1JFh/WyP
Oscv+EcKXfHsXEvhhabW+1vuHdVUUTt+omNT3B92Uat9rppZwvmUWYdnkxSV
9w2hzHSFb0FyjP37CLmMKnmApugYz9Gk7giU5MbsILpNRECl2MDg/fVasXoh
XxsHh62Bla+diIf4/6RRpN0E/OYQGAq+DFg9zo9vWmHa7/4SGuXR6D9BAkRP
qZWOBapESaTn/niWR6JyXCBAuE2I7To30GL4KlrGVabV4+hxuU2h38XB4cOM
fywP9j0s3HK4+kQiL+zgZIiSWa4dmIoHI/PWiC2rS3doPpHDpELNP2oWBPh8
ucX3N3qg275/K4m+pjvWrf9iETJ4aRzfx0L83YRENxgFInhNNxQrZHEoGMUb
unds9EdgFweq8rxs7z/pL42S+GQX/xfn5x3RHCXkEaPuT5657Py8/eLkHCr5
UoD6avIOG9QymfDjoYHpE36DWdyqUCQEiiwfSfygb7LslveBBJ4QK7BzcTEu
bkDVMpqDzu7TbUImhJ0kON6hsS1wQfKsOYzLFq+1qZgrSJvobC0OyfIT32nt
L7H5I7B63fot+L7flDfn+GP7YAJDY2GImWzT7XTnHJc/wSdc4D5f6YOm75P6
IzVh7WAU2FFw7W8jvIU2bX/NNqrw8vf9Se5StCOYheULUqfVJUFQpev5UbhF
iozdFDcZWac/yV510yAJ8uAkf2DE9RkZK5mdLZ7ZXpjIFt4e4irH4tbeEqGf
pQkoeADyQNFBgfiQAFpiBlJdvZEFJbxZtlYtPkHyf1olYRikmcMDtygWQPTM
i8R79rRtT4EMVCajWEKvi3EtyRYdKZZfLIrC6HfOKO//qet55ZL+/4wN2VYX
5u2E/33AWB94OOsUj/MoAm5g9nvGxPDnk+q6E+gbarDFfP/GqJm0uN+xhKkS
IRlZsNqRe5NpqW8RWSrNon68T4A+U/DYiSXCPo7aBPJRNcD51zF5eAe2NtLv
yMF+ZRVVVpyKVCy1FihQxj+zI4Ye7wtLbYPA1l54vOUzFGc+nt89CHwNY3MF
dAFbOCrlPbyhtLpUGjgXvyoy+kXi3t2Lq1IDdOVqY0FB0wDiqbRY/pjC3Kr9
D0PhKtWFTmvPgv1elUxTLR51jT0OmUtVYUfjgQa5pXx17/BoraNPIwB9uvWL
RZhmtoNaqFbJQdrCymfT9sBe56tgYW0RjTnfoabsrtXB/Bq15QaVBRw9XQIL
6i9qYQm04fwG76KJcB8X5rGinIGV6cw0yZf+FSI9KMofu4pi2ufOj6rNXqqe
ak/z6H9cv10z7a4DQcYl1oT/lAd5dWoZi3Cah4+O5H1/EfKBC1B/85iy+JIe
qTiIxrahrrgPi98kj0hExWXBEyK0r7x0G+Q9BkmUFP3YcUs3EC72Bw2bESLJ
SJ4PQioN4jWw+HkxXTPjX/lWObeK6/CcO3PvnmgwF4S47x4pCdoRBfRJqvrD
c7Irzkagw1EIgiTbvSQe54ZCBhM4dUzWn2p9VZE/++ruAH/J5ujvNPd5WJYM
VbncOkPhfHoStf3ZGHcNBc76LvGmkDyv/QHaYLpaNanrHCTl1ImT7hIQK+/M
uqFUBp9gFQmECoUWOiULY2ZHp73iFPYVNFceRa0vljw6yEbiWMlxmSLWg5T6
vKQe0i2puR3gBRfjZsYFvKVxb8EzkLEoShGdia4WsZ01XxCFyHzdr5ZQQ3i4
XsJzqLVyLZyj8q/wzcVh0/li29VkvCboloNHa9UCrljZA49FaJsRnrTa9TV1
6D34BmawVdDlzZEpqmb1hYLg/nsQ28ym1OtEqvJ13Pm7+LAim3iJFotBeic5
j6s+HNUfRH3nCPVB4GbFIwiV7E4OMrxnd+vIN+/2zgJR6izQgblZGycoOZYn
KcsW96QEoIz8+Q9Cl350WDqS5zZmCxzqB4TttkpLhhGE5rPo0b38KUzHpm25
jsdcAbkG12S6v/Et/MO6ajxWXSlPepSu8WXBBVwqTT39Xte0NvXMBVyxDyaA
4VxnDIoyh3n14tWIn1S6160QGU8Ko89To1MpRt8LrTIhrteJWyAQOcjlWEQL
wRYfc70enNpuQCDAyM4BYV1YF0Q2DCm1YKcU3jLSsXNXlX8RvF9o2S4QF7kY
2Cr4tsOW+395SIHQGdMDGGKGKt5gybukD+wbSjrdDz95oV6w4mZi05fVzr3c
J5rUc2OYCJuhJYL3HnKh4EzH9jIZRmwDY+6bjTFtGf2Krw/I4YEd2uYfesVD
31OE0c/3LkpBo+vuan8FzM53mAGh02zlsZWCAviUAZuDvz6aTcexFjED1Oq0
Xj0n6i19QWYxWc2zFifummdJzKtjvUxM315OvBQlrWXk5CBISg+Kux3V/cH6
AG3ugdpuIKFGPRFc/+Q93920LZIAVKC8eCBXZEEec8ZiHVO1VYMMla5PidNg
qr5ZJjEwarma0aPemO4RxEle0sSYpjMJqU7MHXZWTFfPDbTltWDXqfNL1L96
6k2+HwotNmDPKmRElV3hd/bWfBLS2YvkEeGEVWUPRzOwkYraEgr0IIUPOJuI
7OiV+PemuqhY+0Ad5iWl6vWLTFy4pfBjB3o8p1DuthCd9jP+ayLM8Unf4pBb
KWUxKNaexxnGEvy9SiL66KFY+TXPGRQOxvaJNVaKNQD6FDgND4Y9g0dq7wOY
dDONtTR/sCVoXfWM4pZghrbA5bhEhH4e/47vV/+ciAw6cqwRMrdXRdfstwSF
r5EG44d9LRCziKXUN3HeX97aoQ/Q1EETdGLY8/7b2m886dFoQWWu9A0HtReX
BDgb6QTgp1/LC073OYmMkXVz7ufSJ8zriPewVfIzY6s1+5wpQgVq7ze4KZQJ
NnCAo2JRQRuyQiqWzwYmpnDaezE79n11QLh0iZkB86H8JK60K9h5VPyQRE/W
WLyRwZIZjF9vb/1ZZ8/Toc9RoWQqzo5CF07qdhzPXiGcJk1bqOBnzXGg+8h1
2AaeOEObJ9mnVbOMfLe/m/rG8F+Oci75UUNkTiMguqUqw3XAgqBpPLSP+W11
P7l0ZF0cX0LqGTLqQ+XlNcL2ytrPN1xgIsDHKJFq0sXqsLVT8nVURrKm32Lh
x4iK8zXRwExM2A8EFcxzQ7zlJ1pUdpuz+PYpNNJvkpvg5o+cQ2ZbpbIhB4/S
JZ0EYg/eGq3w4Y00RK0vABdf8k9IPUs5mwPWs3/ngJAIyR8ms0cd62tAysEX
aPiCsozq0cCw1V6cw7gcAi9B8RxADSdVlGNJbxiI9JZQq3LK9Mu/j0NwJFLd
/wVsZ9a//lVS+WrBijmTna3xA1Dj0bNWUnKOf2ujN6ppyUmoSzPD4Vpk2PoZ
cJpVC0HoARMo4Q4V8KmmAwM9MKSs8ymQR/VUvmdEfb/q4E+Nktgek5hjzWet
EBkgRdRrV7s01kHy9nL+1cjlrnug0Q6OMOUItx+LilWwV8T4J5MkGu/QK54S
j+LyA32GOZNq5YtczZ07lWM/zIv591ci6rcHGeKNq4GuW06cTPAJBxTf1ZDn
RGS6Hb99oE0vH1nXTnZTnP3kX5LqFvHDTrjEleQMMU4rjfqDmsJmlRX/2j1X
b1MKwSpq7dsIhRtHJG107Gz3gAt30A/MutOGF2hiNxRbDMg6JT/DVlgkNUy2
98AFZHfGD+YaPJGr6E63FHDW9wUytvFX09M0vLsB+KwuYqA5EpLjLxngBWg/
vw3B74P4GiGLAErtSGx+3d0FH8jxGTB/F7YIPqY51B1Pe/HASxaTUm7yaWVz
nM5hA/pHEuEYWafXz7xjhugSi1D3TKJ0JrP1atSansGo3uyZGehb+NzQLecd
d+CLl2WKtFnuptrvi+FbKk9wU9M9fEy/bEzwfSEz+69jqK3P0aB3Hq+iWE6U
UrAV4EOfMVo1w2d9gpfYpCJhAExb/66lsnTAzvuozF9xU6ETk6ZJTGe+2fgX
Qs7O4mwcmBKxhNRUmMIiaAkLnusIlhX153WAdmoz37Pmr/N7UPGuxVWWa0kW
kJ2y97VuVaNAixvoQTROurVSBxGagMi//NCdi6lm4wqNUATD2Acd0bCBAnKQ
I4+xvKPtth71v4IEx44I4MV1mf5fgmhKgd2PlCm+CIhwTDjxbdf5Hpu8d7BT
JnSsdLPJD69MWJSzTtOZb9LAPthZpGXOlvJZyx9dz7z2T4ByUeWVXAQ/RPra
PT078mxd8fAqAlhgIYW/avj1+y+RusHvHzsf/c4vZGn8rmCiw2SvIia+Al7O
fEd6YbOjgl5hEnslvEJ7sFjkwM/Hj8JaZES2jR4P6dh6Aa4B/+vHTcgSANE9
VSAjh6EgqRYb2VpwnyFK0EG5QD9lQ7XGtEg0KybV6hxtuLZM+GhibE1OlbKc
E/mhW3rD8kQW2ZGC+ho5RbdMkzCPR1qcM/X8KlxJve51HWX9q3EY95pTPCil
dmsKEi6CMkbLYQh7DHYLzKFzv3wy8jQVK6X4Sp5q07zayNbrtxoa0s1oBYqM
J6hbid13TW8SC/pUF+i1lj6xE9WRKHhuvKFlZUngJ/TUk2Y/5VyWtQbByjBE
fzVOPBsr8z+6wFTSzbGmKEzn5D4edg8rINrBKjOx1xid0reG8c4UPYjZuWK3
WPREuuXYpnGV6XDF3+mVCAQAazyjqc1/FzRdJUF9Xx6esDGMqe9lo9FeaQi+
GRlfNR1dyEtO4nuONoB0+Iw+gFvHEGyEXuzAK4nMC+IA+3IN5B8OM7FdXTBD
9ANsxKnUlMCKzJXD37lUSv9pObWQECHjWzZqjTvWCHSnpIh4o2vtWKaOY4bR
RkVZFE5fI6NsU9Ek65W4EZGGnrhJpV3s10bk//9rOLwIdVfSIRugdsiAXh2k
l6nVW000VA0GwaGz8AlQacHAiSYV1vj85GJsGHXRjR/W3Le3m7cVrl8aEwbB
JtMM0oES+4/FwgyuBMSUyd/dSssePWZHRyuhSxJVbytjZJt4hp/xCcxnL1Zj
k7PNW6BddZ3A1uY4d8PEEcM/kC15Vg4jKXKXEm7chDvQwGMdB1yfXxCfeDoQ
jv86oXOJtUpejl1WyDP40+U20tqJteBmixbzaUMNs+dVjOohsVh7i/t1Vm+t
SW51OkR0nk/oeuI4lVWIUK3b2RCUVKoQUOv4GkaZFa9QsqGtMgqLfQ3ciXYO
WTo0cOn9mOhl+eb/1hpEZ1BvQJ4l+TTIY6W6S0LfA/hsOUBVPrlnaJjsYiqt
eRjvBavV9XUPGm7LIXEEKaZX0J+OFNhGuE4RvVv/9BndK/T5YezMV8ezuQD4
JXahVmmiusmdYl2uNQsn/Fd7M+ASGxB7aRI3qaGM4N4zA8sd1HrtV4FKUzhl
u5nwlE4be+/6Yk1fM8754yCh89uYIoyBU0ljt9UHj4eQCNaTyZN7f59sYQ0A
bWFLWT7xkJF3j5R4wAPT1XULk/wmsru2YpoXvQJH9eibDL+FWmKAhWzb9z8F
6eWn1ip2n7XYqDDbK/Wbkhgkau99bpQ9nA9VbsnY7eiraxxMdcJ8C4GmR1yJ
UgJ4NjnXnPsJPAy6ntObPb5+TKmBcfOatdsSez6cGfIL8+lpIYxdpvj+tsE2
HoEgmc7D8eG1yxLm5r26ugxuNrALqICGEaSG4fU7GDxMqfzkCPEKfasMzHt5
sRnMLIKo0TYTOcSt/q0CWRsaaeCkoMT5N/1tKtLq7VSl6qVX9YhKlJaoVrcz
tW0QfbKsfxqRCBI08Xc5HOEdWcD6pN6fp8XD5Yu6575s3shZPC/6FjSw6jkE
t9HXR5k7hTnwswNWyq7bgb1HSt+hOKASmjEl5sa17JWnlzdBoHqTgwSx/vCG
5PVAbQqpzAMDx6+kIb+bR0wk77YC5B5FN0p3PXWpTMJX489i/GD/1EC8sn7r
ZQUZSgIHoOMfSkoPVVsFcx30IN0Pk9z8xU60bVPYugpePBIvBU1Cy4SE0Plf
TK4JPwXi7VupV2IccEteimejB9SRy9Js/64OWQ7poCn87+Voeh9t0E47CLre
ipqwJncHMzw7PWFRjWagceRcdyA4/anfX1xp0KCKVVj5DAdeDPuCMGszHWmm
ZsvzSCPyGw6vcIa2it43SC0rMM4cfVRT2V4ukeWwehRmeo85JzfzPfB+a0IB
4gTuCWwrdHZwXXymZwCerG2d9pTWv8fw/i6jIPmQmIK7x4Dnd/yXgzYfLqTF
UfFOqTMxQtJEEB9kXrPoXOZ9caI5SlWV7XCKZ44qhJj+jB8r/Wn2Au3t18xp
TKJaLIZYzWoMtkDHEt7oY+Y9p1aRxrO6NYXoNk4KnLP1N780fTJeabvJ0PRk
Cxv3Ciy/MXbuyzVWiSpkBVnxMHL7marQxLSvzM90JIG1+IFCZ09xIMXjRZnh
V/LWvao7QQH2eWt2LR6W1822F+iQD/pVmC7ktEzfFhKgkU0m+p2Y0MB9adTM
Ky87uyNJHol9Gt9NDnuk4vXwWecR9Mz0n5k2L/MYvY97D/6mR7HyIdALRFq9
QGMcwJdoW7J5lUKvIvLHFbDi0zJiPnqbn7mIS2e1DCWuH4emXzBPt/9bm01j
iW7umBW3iwZexhPVzcFbm2mHqifOaLHgyI803fA3UquY/9k7jQf6O28clZyM
kNELQn2jdhvNyIdmhGTedgS/I1ETiwymizp+xRRmp7O7oI5y7//8ikc3VF9L
Ku1Av+EWFGoRp7S6yfuwUa/JfUx5wDSFjnRmBz9LOFnUmYr1FNN/LUGg3aCg
xFCLccypzeqG+q7YPyjEbceh8oW9pK41TrB8oggOP5C0kCQfeGVpw0IcsN8x
q2ywRARoGK/KLYqnTyNdut0U3aDkGWQuz6n4e2kJXYjpc37gdPLCXXrtfodQ
30MyeQR9OCZqYpYKPJ06gYmZyYMHwFeQiO67OiFsiZ+l3iV8/ydcdaP8iW0Z
sU7NBoTYp92vqIQIJn8ORauSmxJBWh5aXy0YML9Jml3zXDzJZ5QF2e0OnYY1
hdXIJeMc7toSnZCxeDm1djE6uuA5W8VGv/jlYVhAJq+qMBnwa+DL7gP2uvnt
pA8XMFWbO851dUXOBMdFLRti4/hI1/W+3o25WlaG5XA5rdDP0d5CNzribxLG
xz0P0cif1A4+/ozYCTzrU0KgWi9ntraTRJLeg3gvFna32tuoyowx8Kpl6yhy
FblxgihmY9vNX9bszHIj4yGIFk3D4p7qDBvYffQLc4vJyHe6aUC/e5Jn3ryJ
Oi8TTQvqEPTNqZeV10ASG3fwX3sDVLrGppR6poVm6JZQf3p7Bm9WPofoZ2ft
aL2QtQIANMBcRScy6IIunSPAd/Zg/k5vOp1Dbrv34SecWsouksvvgukJnMP0
tHa0/AayFGwyZlOtDr4t78T/nX6R+sbBanUHautopSOtMCt5mRifQCxfjhmP
bS6FjMgS4c4Ds1KSgsf9Zz13dcakHrAE8O+fD5RQLBw+7aKwmLcPMBf1vCg4
ouqf3J02dTTv90XDhGbnzky4c0r9OltAdr9jYJPaBpaVrjLlRJ4I3WwGqNmz
TawVkGLRZ7sY3oWJxWtcrlpYWX3gCQ9RBT7rhMv51xaT9WxmWqDgwCbuLjkd
8FYwgLCGPw28XK7G3pXSJzbvWxbJUkho0DMittnM8iea+07iRJZs+LkJXulA
n4me8JmUPgfvom0sm7zGyzPtfjjSY7Radj6DORigVZ83NxL24nQiHIfR/snu
56/7atIj8N50Mb+ttJMjy1W1NyvobTJf5NqI3dUF1mNNlcrt+IC9HO6DTRcb
I/ag2fOlbeyNmCL2fDvDXaA1Tf0hI/HCILepJLr9D2xVohmxWLWaNcvHS+jb
3johtLbj+xikwtorIj7vMLfIuQN5GyWU8zGxulyhCZNFsOKzi8Zyc84EurHk
qLZuawFG8mI/5K605vusZa1hZBxfpreA1ITUhllot/3B1iU9snCxioNObVjn
Q8GKW3WgdPzsrmO2fg3P8paOSRYGEhUdpsmLXY6Ga+Xusas+yggcwMlX8ONC
gfI+UDiaIGBCNhU74T0tL4an+ufBppjG/m/6y8jN4CdeVX9AiHnH1aOh4L94
519seLmK7qoJTILYOjXRqZy1jE1CYns+bNjpPzIc1GZmzZ2WJJWVhHvK9l+s
2n7eHpPeE99y8ZaAIzjjsHLvEDaCiuzXa75AP3j8XauhOt+cxTJaKDJ581kZ
p08xSf5gV4JlGex07DLVJddGnv/abJy1STWbZV+3mEvGBko7PnAhQfR6AYdF
dNdgcOmqWr5bO/bY6NUwRJw4waf5lgjv4GlqVXQn3y3Xvcsfgzt0a0jGowbE
zFzZ2bQbdZu+ziMYcA2MePqasBNlfd88Qiq9UPai1+gRabIRUrD7UTPh+PE2
/yb2W0y3h6s0SmLmP0Rusctk4YUFe5ygXhqDm1DQVi9aQPNrqQYjYk7pG1MN
+koJWStlxv1WARIuEz2OqROtUZ2snMhlW1FkQfX5iXB1Xr+seIy+3pwpTmFY
FoFMRRkztJ74IYrgUKgMEMupjU1HnbPh93mW/o4baIiW+kYC/hZujto5kO0i
YTUHPVJW33UQ2uAXQNfI2fhnjj7Qaw6ENeARjLSsnS/59DbPCB12o9RhcJgp
FPvfTZgZ5uvxNjQcCkGCAMhHJt2DgglSySCrKOJYzS/4/+R1C/Xvjmg9pYKO
OOpHHgE/BnQV8pqfZGV5xNKv6FjVGmYuLbM/lQm+Vg/LrPUCCzodW+3uCdTb
gVHLaaJ6DwLeG1AIyvcJTQQrrtNX/G1WXLzjzT9M970120Duw16sQjpzmyK0
+GQAQNCtQajLOEwSibuBmjucE8hJAOjKFaoDd9c8hvqaoX4z3MY6oNiQb8a9
s+9TfZjB8P2/vOLZ0bx/NQdWY1N6QI/8hIQ/zH4knQa6csVOq1bEDkPuxHwU
ZIaEJsCuLVzY3X+SilzRjZzRpbJ0Pj7uPY49wO4FPpQrLQprpHPVN936X5md
oL6BenHthD8gdX/jcGQ+1BK6EmTGvzH3O9Sj/0F9JRrcvIjjyjHGQiZHP1tz
6188bK2j4PgDhtGK8I82C817TamvimLtS0PV2tNYar/kV28YUHUsbKRPSKhw
mbEiDltE6mHuDa1dim+cHBj7G4jmqmiyvOOWrS0qNYupeVxvJW+c71rR12Ca
rs/o9PbSYgaSGDVYddUCR3TrSpVipvksueqpDm0O8dG/9VJ3+dIz88iltx64
8OVGPlBiVeGPiq6Q84jSh7BHG7HZu4fr9wKhLy9Z/KF8XyUdmQSCo2Ko5UwP
uRZgHoYrvgtNxpXy1oZE4JzTVckeVvU1ev7QIFqIiWBdaYfMSut4TQBWN2Nn
KImx31WkxF0DeszXaDcE6aKwgI60C5TMWhvN384mtt4bXroeVbhfilmGXXwD
JqixE1yuuRZylvZepNtdkM429gCMnQG4/BKzvyuANtVftYJL44J+GZaIlGmB
+PqrwStkuOKHQolh8f5Gs6JRUqArBFhQv7X16dG6ZAFzfAOZwpvKMWCbe6H2
QJf9kVnmEGG3DWDT9l9+BxOt8l+WKADPIDhG5QDbFTytHYgSnl9CTl/FgLPF
jgvDcVanUUFzfRnjSeILuP+CbbEVAnwZtRq1U7dZA7kWWHzKaromcprIrzae
fcve+H5ExtPZ2mId4n+SYhCKVGCfOpeME1ZDhqMiKZ5iMPSwkal3ANFRwq92
aYzOhWVTI8/9K9p2zufQg4Rh9sS5u5i3O3A3OAcuv9s9CEwQCHObbTPMmgwW
ZZ3BmbKOIdT0jwo0QbFw7LE3bFL19ejLdW3F6kw8skSpaKB7i5xp3hSj3kaK
oe5ViIv9Y6vJNSxr/72hi7auxse3E47AHx5HQ11hUJrx0vsXnBNpTjzN/+D/
F9/vlzQzSBkwV2+YM4j+2qjz996mZMyJQ8RUaJHM+Ycp7KxyPoysiMAQq9ZB
3GFlW8v27E282YNun36M5d4sitc11fQo6hoZmrnv86fWSaWj/EFPMW1MxiZn
XDXvp8ObM3B5DMyPsMBTkm+e5v8sgN4WRPfPVkMCn4DSTxyNGcvUOsOm0tlS
sV8o7S5q9SR1xSCtovZNu7kfvnwMxGmAKggNn6aURDfI5L+jg0QQTpHzuIw4
oovW7geybo+8xrHCcR/x/OlIqeGgQPkWdSrcZtHRQXnALEFVhqa1gWjqK2EX
WL4p4061rT36WrsI3eFGXfj/oIH1QH57r4TQGZbLIpJg9gQMkKb+/DIs/wBc
jxdYF9Jc0t+vVRGJZv5dwy4t/bib3Pv3oI4dB/QNy29lrC0MT3nLFr7musdi
Ia+eFnT/lhIsm8Ccez4ls19M2/g5CG8pSXhmQIzog4ZElvUuG18ZXfz3rXLh
bbXW4AptmKk/OzUBhI0W8JWOBR2fWwNamyxjOn+Nsw0JLmfBRb9xdFUgrZMJ
Vbygu6RTQycbkhoqrpcdak1xatVCLrjNoMnFJUZDZEA9Recs4csiA+RvjFMh
GTM9wxKb1Jr+z+VT4SlIa2uVRIHp8ioy0b3J1HXMYo4qBYJ7zVmTB2MXweVR
48z+MiwY3wUcZy3/UTZtmFXiDuSXnq/9I5AzryU7m9Oq0Nt3BuMQG63ft94S
meClTscJsrI95AHAziHGasLsl/7yrsvwr+XrTcEa+riKL+VKjUAoeq1940A7
eFhtGR9Y+BPQyZYdtzZs0OQr+amByHKwYuLUap64uOBB27jp6mVU3CQONk2N
L65lSLtDc//fta3YfyUZX9fULivM8E9CnellToQfWdbh4APPw8hx7d39UGiK
rRJOD29fRD+vTx08nqRnK3vxdMjJQG27IELBVfqonmAvmjG4wPcDYWz2Sp8s
VyElUmN0/Zyoe7aWNeN/AYBUuyIJpNqwjIL9T5c4KMw4zm1eeW1SM9lcjBlx
gP2r83lfiHKVSBJXC5qN98r2yTsa3l80T61wb7EKyUvSkbPJDNCV392r2ooJ
FM1wt7BxmqpikEaCETGZdaMJ6ktSMM33DbWlJVgxJjQ2gi2x7KbyhZUAA1zF
BIrnZkRkRy9tuUzsbClTo7yqQ5GEFKIHh9V+08Bgid+KTdI+mzdC983w3oOA
xa8Bx7wy59n2cwQrE+QwogBgTLH5V7xF0VvEuKfzJirsSkBBi2a2l5HXhbTF
7vm0sLURTCeqqCqnnJdXZ3w45lpbuD2Eekiu+vUWeBwuJ/k0TEAoDbzlNaod
IXci801qJkFSa1TFVSNKpLMdWcxF4NtQ2oQxTnbOsY29Q7SvH4+jGqyJjftw
zBgbuJB6oomXRKM8lA/aNnauqCVmbQkTg9C7HwodlDvv+pnb5stR6ISENKdq
u2z/MOL9OiyosnMOpsbm2iJRCl0RtrApOotJuFXPreRvQM8UHywgtsqDtBQD
gi71Gj4I2nGQ5NRRYS+UdgYMCdfUXcopRAzMVSFC//l7WBNyZtEMVqdebKRs
gt3l4IhmmXu3ikE9kif14K0EIEADFFSNOGWp0Xo3IGZCXXxIvct3P0eqnjg5
l1ZTRjYT3372u84EWBdbhczDsfADF+AJNL/X+StC3lwuy15jJV4/VERsp+I0
+A9J3szwHd5HvL/+2LHxBtM3BmUp22k0BqzxSnFgS31K/F5uZBE1Kj+R8vDH
18mCpdoHdhX1KSgdQcC6u3aCK6Q8KR9yOLk2T8mqcdEi6Ne0Y1HTb6rJk7ao
gO+CJsbJllf1gVYAg0lce1WX4Ag97PN4zWqbk/4U0EUU0DGLywQMHrqPhSvi
Al5vYYOh7c69CQWIAMfyLmaV2Fz1/z2Q0gsNYwTBM+nioj2n0yz8eAAObsu8
ZjKsYET5o2FCSgKgMyKKPZGDIvXZtvUDgT6856B6JExajl5+yi3DjCJB6Tm2
ygujyiPDFesnei0at1sgrG6IP1dymOukWfR248jUnt9o5lCNeOu4Zw5AWMhg
2Ru25xgzxZ1+tYCQI1mz+jiTiXZrZc4QK7ZIaGvSQTJDvvqNJru5uw38gvxm
Ir7w1JC5aiCFCv9aucLllMtin61V8VUqn8qg0bCPDabd4/ioyz5fPauH2YEQ
cE8x7Ueyy5+r+7iq/pnrBMJfDOM4qV2w+gnCDY/vA829N83nmJh2tpEqw+/m
OG6UaLsGuer8Fg8D1P+6wMjXVwDWYik788EwstCpwNDW518TPk3Iyiw7p5dG
0BbSTvjUAI8brn0gX//V6PN3ajCMPOs5J3DFuL/x8NqLlxkttLvZ9eZyx5mt
8CTg+dfohIBjnYXzUyKZOMqlAQvAj3u6W44Q3TYEN3Ki0S1VOGlr946g96hx
Eo+zirSWERnLBBBaPowjfHT5SX2nfAdfDtEUWiaxCFGvyESeNnL83CCxqm0a
a3Db5U5WRA1tcLujTCI3vSG6rpBi9D2tpIkAeFP30q0bAQxjc5aFQ6xA+vtX
K7D3noRlVGVi/+v2aOXdf6qCuv8w+SaKt03yC8W+m74tl9RyuS8CM50MH85a
jgncQa1LJyoz0JtajWCWe0NPXMztvYziS4zLtjpiq+KEbA6oW1qcztNAgoq9
S3QpXx2LQdMZ/l3BQZgCl3Kattzhxyy5dFarcoN8BBXUHxalcb7HIldDOOlU
BJVzAoYjNjB4e4OftdcVsa0tMXQgHzELnhY0wl/rybSj+kgFB40iEMSW3Y4v
A1J01MN4+2+5tKOwCQxkqFrOykTam2u9MreR970p6Svwv89PTP5CDzpaqo5w
eaVUwXDQt3JM/+1Fup3RFKnnms65n94KYoLesf3abb5IM0uA5xGNad5k3s42
KumiPgYWTrnFmzLhQ8ALOpM3YXT4Xs8HpMIA3a5VQ6b2MTMEA2hBjmIlRo6R
TboxlSnG5nSFNbFKv8B/j1cSaDuzAYdwhO2MeMcrm+DSoTd6Zlqj7mEgmv+g
UlBzjkHMiQtKzZwE8y3Y+rO2yXzafgxFZqGzUgGRsAIlqtzypbRwhSRbROHw
JafSbTu4vus0PFZ3MbMWD7P7PxnVcZG7HmC0E+alCUBasa5Uk39UuyylfrE6
96nfvuDwzTz8vQU2fZWPuzgYLYwWw3yxBli6BDCrdLHkFhfF4Y3eZQ7+LEs6
rLHS3y73Mznhl9Vjb7OazNbm4ZK7rRlWFlpSfKxQv0PrSURuh2vTeVVmlfFB
1zjJPF6W3zKQWLOj7bFMQNsBL95hwMG7azNyy2/Wbr28AUYgluTqzlgTdTm1
6DlTv6bWDJmkivWCMTQIsqHHCwsSgvObb8ND6Ozab/ojuzx0MvIKL9phd13/
+VVjCwOqMVQNZafZz83n13Ovx6Y8Iu5D3a44EmqT00bLom9UgIaY8uB0tlOI
My/0KSlZp65rI3Yb8BhKRruAQYeVAuidx4cT9/NPNhuHBqXatJ9tFjaeBCrb
9WVYZ967KMRS4QymKm7vbEz1Z36x6bXj7AOw2ZJnNxfJ3aXbjc2I5RZqFCjJ
IQMRy4d4lo9rKT679U38U0IylIR2SxflKpI203rPpOBMskpk1AXQiaIa8Dg+
rbhKmRatSz/nJe0TcURH34q5Rf+5tcBtAxdAaBqqNbqlH+TKYSEE8NbUl70m
D7IxDzZDwm/pE8lxmetcr1ujFDM+ElGPOoo6v2KdbeqV8o4xD7nRoqFxKeQA
qJh6WcHtOH3ZGYO1/zN7LqcY9rkckM/wuULRmwY/WgMSt20LQ9FazS5pgkcW
cy3uX521Eu8sGWrMOj4Q7F377MU8wncaBrA1+3/DtL++xy3GiBMv8XlcTWWh
JOQWCg2riWiLdxnelI/reJm6h3gyIWhPKPEsIyfOxDOgL7cq2bcX6URb8/NV
vuQ2zav28FN5aiRp9B2fVLPb+A/JMjwgf6NVZxiXgvqW3WJrRybbdr5mfV3T
zSGdhP0XNZbPJEGL+m/WcVR6tFkgTf4ZesKO0+zpxWjDdigZdl3ASDc96XkU
ZVtVVTjdlMYQERT2E054wQfCPey3TVVqPcMHy5c0hqGKNGqo4PO141/RHtha
/0w69LdxmVHSzCQC4skOh/ETpUDuZc4orvEiehHzcmXzVsFHI5R748PNGBP9
ApU7zxc2AwoCUr7Gvhl3OrPdhmH8bJ+c0MT9EQyYvfupalSilRLgkVnTziom
xXNx6Mav1LcAm7pGU/BTI8btP6EqAaNHKJciqbWpNo5mEEi1hh+4mcJF+uaj
WANAetfeY5zZgRrXUx0MG+UPAuaAGPgF3arL5zs7HayEKjCadeAOs2+8oi67
/Vt+PGPYbxw02f7FMXeBKhkai8Cu9Ok8b6T+vwnz+BMyfKaIAlHWL8RQbGfN
vSo7bTIqpK6080C4XXmOfMXsCrvYlC4ZZeVvof/m9IHI1BY9UIO1TG0L6CW1
MwkfCvKH2j3sQ1tvnreyaPjtaV6xqHCXRAv+PjgB6usqcnW6dYBlSH3TZOKl
iwMJRKvWOJiiaPCMMuttyzsWNLC4z2Tphf4xfd+oSdoBkBnRKRJEm26M2dmx
PxmkA/X9lNb5Cq5sew3oA/w8NcxjzzEsR5R8dktPE903E5ge72cefxgLZiQv
9QRHMTfSyRxwCaWFFoJcAuTUlBSzbjGbBPXQ/GmHfAg/m/jl/ffkG/wsWzPy
yCrDCb8GlK9k1rORmnoJFfgvytdEbUeeJ/L0QOzxNUvSGqWbxQNnuBOLJ5eH
4AEvyFUIJpzeR6D2DobnydQHai/QoEJskvhfo0Rz7oLpyDQwAhVN2kuCW64m
C/nnjyXP1Rwz8p0bB5kLaQq1Uo9+sUXL+Ww0cjjaBS7VRQyP3hApUe8fhhKu
83KtSkv1+k3h8WWPzAB90ZZiexGsfGeF/u7R3F0rep4uXAU6o8CVTRh5ppYT
Jh23VQG1HzTjexM6ohnjBJtqyzDXAUa2QaRtjxTyzdObjhtODupExXx3pV0A
2hbsA3mOO37qgN0WEXRSBuvdvnyIH6qbpvIne02HFSNyLpROkDxbkDNf+tQu
vDRZnLjJP7uzuZ3JtgWNgMqu+NNKQIR/yTAZEEqqJfI/26sH/LKwaiZvb8Yd
iZb+WvGK+r1cfLSJtAOovsKqZH3UZindQvRIa5on9KWz3YxpdKdGf0VVyqfu
U03iKE1BFDpYEM0YjYyO6m4SOpqdiTRRDAMLyuIkLKyVM+kM0dgxsLB+FH9o
fUvu4ESVgMxmNOdL3ItcAFgBnDch/HjNdJKGLtvjN8pRWcCF1vV2o5i9496W
CQYBUP6DoN2LAaPcfx4OIdAsvNPBSKs9Qm6szz7JpXFwlhFk56PowU9Db7xv
hzTvtT0VBWfblcfwzYIO0jNd+atwQFjIekkOUlcbK46Okz9XiF5IHogOjFx/
OVc9dVolJzAijIITBWnrTpPpCoN64O2yiGx9AK+VP3u4NyVcv96PnU08RaVm
KUQKL9fZrS9vK3F+PGk3RuMNUEyj0DNWuHRMFPfnXifSLO1CwvSLXkunq3Jj
cDVb5fXuuEh9h68x9lW5MF8KtjAPQLTDAWU/64XKF0CUYmwpt0roMq1Sxkon
UQLNG/a37WE9HcCfDDjy2Zzc4xAsr18bvIOQpV+EfxOsEpmBn4eljKL0/Uvd
s+ZoJh2TWvPN3eypNa0vZ+oPHul9Sh2gCvpupZ8hOI+k50SdRAzxgOG3sY6Q
hVlEPxWv7J5qE7TkzShncAMvpDI3Fyx2zyxPh+HR6a8hhszAkW6cx5qB+TQ6
Qqc/5AiUw4JDltAb7+2lBRC9O0MAAJpcxUW2Sdp/uHJIShc5eDG5iV2yEXc5
OFHTQ300fYGtBPBR9WlzlNwd9FDSA8NdsgnjkptYkD4Lt2i4XfMaVYKi0owi
qUKLEJ792qLT4wz5X+WfvLl++a+qsq1EE15OI6mDut6bbVp4OyLsUzLiFgta
DiQta3vwPhIPee/O+xDEIUyayo1EB8eh/tAPDssHm/SM1XVp21Qe++PjapA6
KCvL8/d0hhQxaXXb73FN5uB/T8i/H0wnXmjp5gIbT40YA3zMStgeczkp9DaV
JNGKEJVnlxUcnjbl9RaoTLmWPcwkOzSC0AhHw5BoEp2kwTPhV8PRLlewaQU0
uLpeS5Yuqnc0hErHHa2/NjDDAB9L54TTOvohzvZLyldkZpfBCf8up7Q9eQKH
3KAYPPb3yKTtvFFY0vl8clQrg0T7X9OL7M5QkCIs1dQ38vWDtXiDTVsssv4z
9OZzO6FvA79g3QatUuTUvHLkghZDm8JTN1sxnKYoWwMy65ZNCZ/59lNUM71d
fKGa0/uM89noWUO7LZLy7nDTGXb58qQmdSHWBrTMLRVTyrY8tullQVkoRThG
3x6qxyS79SF8EVFR5HJb8MgjeY04H0tjwPMLf59VIaBUxakhjCm6K6BGBW1/
rXYuv5K0SYbsJVjdXMSACccivfhTr7AUGPFAhn9bTZf7DhhOMgO2NDeQCoO1
ZjP4mUs2SLyAOKypysooaK5QYe84qA9WjAuj7lHuX7gjeMsiYHAqFTbWVexa
1uLZv1ZA7dFrsFtZQyDdptWJ/VKkq8bHT+O5DuBZrOqUEplGowLv/mScDAdk
8Orr25RR2QF6e01FfQzRid8DiufZSIAGKUfrOc098/xSbxl26jNMmJtsW9tV
xoUWadjYJ3KwJswHXYZIPpDTzWy//KKLe37Q9xUUPjxo41eCxDCSQdmr/5Dg
za6qSHuxHMqujq5rCUUn/Dbh9Etj7Lhh67yvQe7HUQzabjO1pyTebNf+bqMc
ZtTEU3uCs3XT5XXYC6Bua5p3ZwWR9uqeWVviuo0I2PyhjYJrA3oC3vD3e4bt
4iLLHEI8kzdcuXsKhjtBgn+/ICN4I6pr+uGwH11VyGazWT6rwWcLy8T3spCl
94foFeBGrOXOU00Sefc24NvsfWc0I/cPEpooH8k1BvVVG+0v2LkHx7467vVN
6aWEZnCU4YecXmlXu+EqkrybrwBevNZX0wLj4t2Cq6MU/smDxZMDcOd+szia
h7UWhYIaDLP3KnhKkHwxqBom1W4WCsM5nlaqdw1TgFxjIn9hmMLoJOxOkZ7O
P9OWBnINwAri3abq5s+J/pC5LWWePPke/3DG7pMYtFq5RhjIgmu2WjeerGYk
jrJlTXVvyvzKTY2nqBwJyBfRe3r4WdlUuX5sjynl6TUY+1kmjYgODJ6aS+q4
AZBrcHCcWsyYNM1VzVeIs7ProUvQrC8UKZhimnmvF2Mc2mGorepZE5A4X7+w
Dqeeogamen2XHgnwHQrC5lOIyXHeqsHG2FxLH6yqJLFHDa4BiLyUuKJi6W6j
BXNFTvmZrbU75OG9Gwcf9j3uvcy+v87txR9GErqUiyswl9TewHfMFgLbLKz3
GzrOXXF5fNIYcqtRvZAyWbtqKuvLVWp+sAZFQX33/TpDR/Bzc/RAG5wrq7Y8
Ny3byAlbapLZUd7v0WUl653ApsIBj+eVtbyzn8LkkNuVnIIqohYbqKggxyxy
4yL97sY28j7eceUhuwb8Vz3S5jWztoVTPlI2TYIdjhkBoxF03hBLtj0vwxGU
HMl9aVe/9oeZgye9El3tgw27tbNMIXlyA3cevq0LO5RmWLibdwMf8pLluAVW
zmNyKVPmvhik9MmsxUmTwRYwK9/S7UW0QHi05RktbE1gslA2hzdDvdP4OpFf
20QCCJyZ03nWXqotJ52aB2uts5AIa0bg1zw0qQjrANaNFDmYmhdru68OvqDU
ypPqPSBCG6KtNJrjOlpus5QEIHYQ+oIrFhsMUht9AAHWdMf7xfcJhmPlguOy
ixiSlNb9TjO6odR5frvSDzJJ/9Bzaw9QQjB2o52k4XErIzwlYQ88eQE0tvEk
0eCnX4FHACoJ1YwSq1rZ2dqJqiFTLFCHKnrQ5FLLJgU7WPea/nry0qong3/u
RYZMMUxUTBuYYVA3wpuddSKcx0+1jhpwnmSp6Cr7DwW1TOQnZId5gOuzN3sq
N+GkHZj2DPuoTzjDkgeq90JfvTHj14CbnysX9nnUKZMZj+AXcsMoF7VhAb6k
KhJ7jTrvVD5M0BVonFnvQjBxvHFmzlr4l9GdhuCXv2UuOtw6V52G6hRaKjGo
o6RkOtVkvUbc+HVSBISAkb+GeRmihFMwm34UpIBjFSmifIGmn7cyQ2ljKuc/
5bRbIuXev5owfK05WMtQVrrtjGjt9Ol8vumVP8/8fbV8ot6ujRsm2knz0NBV
FRv/apP36Y40QrbsHzg1bbvGajqxM03I7/yfFBPJ8DTo++Hkzmg2h05HBzz3
GEO1TFKEdQ7N50coU/WZWgkBMidpow3tz8Taya9I9F3HlzlOk7pDOl+Nrnf0
bxohaWx0N1S6Yp9V9u/JuFIQnPKp+/ZczB2qsZsJZLeqKVrxKA9Y+LEy0Fbk
rwKOQggsV+bhBIOF3R/xUqEXUlGHsz7ZV+GVrM30k+ikjg+I0Sion2fUKJD9
qCTvL3G1p/8Thg+iktMbBtjHjDUUZSlkz1IHGCymDrBNGNNCmhhANdMWGNDE
NMaA2TA1QcJXsqnO3aM+Fc+wKJS3c+Lm2kiiL/ubtkjU8xOK6AlmxXRGFMuz
cSNg14NWIxUibvG9oFFVj672+UfZrW14lM0/yslGa5YWxApnw1Qs3E4jBY8+
ztOVRVV6B/ELFftKCdBSNpDH9D7FlsHnv299tssYoe2B6KfGhUtqF1jKetL3
rl8MgUb/LWpWazRnb7Gf+U/S3wR+PodQzs2hFE4wC+QJHVCXpU3WBhWtKDLV
af5GLVStcj7kHgIsyJDt+5sZ+RQBWiGT1G3UhoIuj9VtVAh6VyOipBPpQuTZ
Rem1XRT2+/gwJG7jAGIcTNj5ToS73iPb5uK6nfNepStOE65bODwGdmuizF0r
MHqTZibXMSKv1YvKjajQjr3xVACVM16WSACHe3JmkFumqRVdEKqIrffoy8mI
FPIthKBdFtMhEzmnnFLDD/chCET1DEF5OAFeDGsxFxvwAuGSPE/ABc1vcf7i
F9LKONx2TYVZ14mtkOm0ZNgHfqff8H897TR01u9Piz9zonJwlagpy5+/Re0X
xXAv/Gnx/CoWaCJk/sP3C70US1QivsVHq1ttN/5XU498+vDvnbnr2wGIWvFV
73D19QRqHe50W9LtM1301P8UGKiQWBlyXCf/mXpw/n8MrC4f3uJl/Mx0RFR0
PtRaY44IrfXqrQbQSnINC90exThaXpeaLQR6kQoohIkFYAC+Rp2grD0IzT/D
0sg3iRWh0ev8j+S7/oZEpENKiYuaxh5kJjXLY+A/CeYLBwVjpcV/E7RmhOwp
aS/B9yTWKgeOtvw92BQPh6+FjWQ7Q+FK7M+InyDlUB+/pGJPkXLMGxKdUEJE
dSQAN4qSQuGVtznnJdzFXIxUn6oR5r/ilPsDHoeLWdFV+slgFxZ8DW6Do9YT
h5fpjbHqQU+Goj78Q9ENHodt4tTO0/5tkBluxuMGqBi8y71rfh5VMsbcR1Z6
sQ+R3DQBT1T3OGO6ZzwuxZtPseB1Kd7pWhlTFW0Cmpk1M8Na8g2LF+oY8tEz
sexjtgwtUD7yMRI3PVnJy9VQaX2Wydp/rwFY9+zEaMyu1glH3IUj7BrdK9vV
3+g/Zbd9U4obZkvMxGfirezBEanF/GhZ+TQqLav8m9/3t/wrVNYPRjrjf8Xx
iYyby6L33mfLMVtRsNPo2jF5du6eYtJKnvCIGQQpuvKXCPx8FqT+BI8uiqGu
3yMaVQLzHIxCNHHKoA7tTn+gPOOpjBoT+GbVZqK5arHLAC90GTD0YSFYSOU+
vW1AKaQBeA6uFfu/S973UHds6pE/K6RN0079sgSxdVdBXF++/Su6LkR+aYri
zSE2HLCMiiS4os5g/5jRXCpXR7n4jJnIAsNj5a38KbPCwhqMdDN3PR4mEjpV
HPyHnYmffqbcZMUAueeX7vYU1HiJK8QPW8o425LoxX6Cvd5YA1PSf5WpfsiM
zN1GvZ3/9BkO2igvVFoFFrOuJ/ZWgRXOlhA8MbNWiZhrK1LMPrAN/3q9xigl
fNZnuJgiS5P5cFBVooC9o9jzNT1oMeZaDPITtsv08bWN4aLGkKS4fu0+bD8j
0RDdg5U4nKfJI7uVTk4yqTsrxbQXD127EP8Wppc76HmP9fjV0piI8rGFhe7j
u8yRWID/BmLGUdB6i4m2NyfFigro8JKAdVIGc8se6m0ALWdbjPmswsqKsOhR
g+HSjIWcv8WyM68FIB81ASQF4oNhpv2/Qt0myx+TrbKONmmMqf8jK0Ei/pU5
O/yAjv2oInz184SWSEbbpDIVl6iQBQO1PjWAwISPjv2v8bRv9Hgkjqw5xzpn
M6660GXbTN95g1iabS4EdKV3T7Cqu97UCMi5enhPMbH1xezRlLtykRxo28wS
4HVp+21CO6mRQvG/A5kBBZzFSNY2au5/4gTFxCdx3tNuth+LUqAHqv8tTaZX
uV7Uo9NZ7MpLdprLjwfDQfOgg2q3x+qLmsbMLowyh26CtPddbjDDwhxa82OK
o7dct9kSpmBAUyH1xr6T2uli8yApK/tszKXmivq9pLsZaSSM1JpOqeybF+JV
UkyosTK27UfJZBxaMnqjVDMpHpbXv9XnE+juAcMPP9DAXUWMaUiTt3WW9HGF
Fqo3FT280KSY7YaRcTj2aB4c+xikFHsP6N0GGlGIEJPa1AQzXDJAWFlZYZAL
kJgeDcB4LArYthkwOWu+JcTxswul+PeRd4OJ4xdfB7C+/7mN3qSF47Nd5oi+
bBE50ZWSWkX2QVHmIUTKICQ55IyCWXyXmV2WplLZq1VQLKRZbIPS4wOid+2I
HGYnioikiVy+ioAlw/FWRkdnu3kHPno0qLis/o80GWwrt9ck+jkYfrA6P26R
jDRIxd7C/mtQv47iioXy7flEp6kcWznsNz1dYGtt6bcRelgMA1DN3OjGG7oX
f6BPkLECOGL/oV0yR1VX8YfH1EEM1zX4AkxEA2tCa7VjWC+6H39813HouFOt
aoMOMZA2eeQ1p7MvNNqb/eDRIRLUyP8ynNsHrFLOdbKxJkRhhGu6o2z/I8xv
YTjKXF7BgctimlrnUPs9+c/mk9jYDcidF1uPRFZl0IxBMA1tW1cQUYaFNuXp
j/6ArnrZNwe0mqEJ+OCSyOfHzhqEEd0tDxdXuUyMv9+fKj985DUWx8BJFK9i
Y9rhzNFAduITIZJkNTtg5im07NXkjn1PIIi43d9Q9WUbQn4QeyT6uzvrh/CK
uEnTqc2DE+RzOs/Am/7gSqfUima6LDvysqIoIMdZ50p4T7Q383/QnZRLxhD9
kNJKoS7+m8asnHfzZWbiePjI8oKy3McNtGNQtgA1kDn4SKKVnuKaBiXiQnpv
4cJKI7lWjzyukwE+3IwmRjcns9+fye2313CyEByATsYIZk07T8NKIfFpoAsL
nJ/d6UI/bBdhnwGPG2abqO93P2x4f2RHqLeHeS9gtl5vJdMOVdVSDwrQDQiv
Iehu6UD5BwXbPQA6YKvFOBTt1ZdRnUZZtxeHk+ifkcAjUVFnNC0tv7OUHGtd
lGy33MvKZfxvpkG49CSMKka7ACV1JG91WIqbbWsa0o4r9fvDhhlI36J66UMZ
da12/Cv/OQIK7dR/nF/Rvs3R1cPj0tsVstTlysuF8unL9mJ4wi1iKtSUUqA9
LEZWleYnDLIraU57XGmKzdkPT/69b+insFbsWc1lOWmpcU7YV1BqW0Ota9Dz
eDIK5Zy6ZKY7C/JpC/QAsvm038KRHqH3hXwUV7ZI4cyET4FInWXaqHh8mitG
5yCQK29TMUl5+VaP2ViA2AlUsNTe12Ctdq26qG0CQDz+HDfqW4kdspJa7QQ1
UPBTt1ribUM0YicqGYVipnBR5zl2eYGa1ACN1WvmQylYIzJ9oVQLxX9wVck+
1ApLGStasxg68EPFw0XHa/a3OL40q2SX8Dg6g1hG03W5mslEhy1fJbe7dMrY
phbtX/+OZjaHU3AZoRIdgeA+UKCDYdelxss+ZsvqxBR8EqLMFAkqOCcZyiQC
JMN1gGbyqztuUy5+qX6d4HZSekTfBjKxKlZHHBVESrls/rOOuHqfcyDLLwtS
YfbiuV5w0EiJBHjY2WTUNDZCJJK2cjKKb4j0uxlVev8uU4fFn3ZjJEreRfj1
ZEAu5SqR+NbItaKYAFuiL0+ODZhC05rrEHzAE0ZBXulX3JzwT+ZQ8qf8HAmS
iEGJfvGuwytC3WUK4IeJgqEkT4CbAp8GNn/8UyGS92/skS+WopvsQ75TTCO+
dX7S6XDgWNrhbKFMjTK1+9PkBzdYoTDe4f/bVrGmQwRa5wfoF9F3fipdwte8
aigfKx9jyrUcrehU8LIt/S6zxhTqty299EmMhjWlwj7Me0heT5vBGZFnwypY
UCBpWFvaIMefe7iYFabqMYJMilMo2DWC3L4Da5NvZ1g36TsU9ieuR8LDZOgh
UoakqBO/xxn7hv/zLUD29fIVTKPlXcgf3VaOmcVFpRQS5v+FC0/YjmHFn7zn
EqE6pbAMgNHj3tuO8APB9Sb04mf3rBMx22h2brillwTDMUmRTkBpfaguhC3O
cvq5uE6XEV1XedbwKLcP4ZzYHu5H6/37B0pU6s3gX4wxsNLLVhrCrHiBOmol
52IpcM5Xa/3ckbjkNlBfZJoKaReXKTo3/rsa9BBNpjcbNgy4317hAfX0IEEL
QcDomcB5C8pIJBnZul8s8bG5jj8m79A8cq7T864ZcnVMH1YJcFIoOg8EVDEh
b3/ScmQNqBNlLUZjmxw6YVmgKV+KfiXCZbsgoch5cstuCZoAxfqsF/cj/T9v
5+qlKlFHpL0b0l7WNchs/GIBUi0ZBNRPzy8P71ssFfXGx8Aj7euBsZTPRqEU
2lOcCvmRuHJMqiWj3yXaoxtZ5ylA9sj/HuzbPZ4zYUj/IK7tjLLSNnMPxnlL
CgcXPToeYZUEWtgKOdVn5b3gHxB8Y9XZxQbrK5idQJQkO/SyEPfu1dENV93G
3baANydT0FOtoUuF5vO9r2cuz72u9ZqZqsxMgteTh/vrY5wlg9sly4Wb+6JK
L/S2eUdPvFWcvfRZWNeDGvrL/dsOF0v7JlWusncszI5DZAivyFqg4163qq13
8PRSulgc+s3zn05SaziPhNQAEDQSBJvR6sjsaDv5ltV1wy5/NtDbXFKR26Et
xg2v456wgxFWgGDOQSKKZ+nNhRZYgj3HDsTpYeajhvI/hyujqNL/ur9oiBV9
X9Rf1yLogcGug0+t3Hr8UDEON5ojnAeeNMxZN5aZJjZ61hgMaD+wTS9WZaHz
Kkb+jRHZTmDNdZJmU8wTFvPWR2Oxla2K8+64z7eS5A1eeZ+7Dk6N8K75rULe
VlzyNttRPgtXm1/R7/c0uwRtsSPJh2jDGRoWprV7bGGtYQIdBms39iT6cv4e
J9OW7RdSB3/PXbdOGdAnt4KlBTYFOlZIQEFelmaPaTpToje7bjYKAP8aJWF3
f1gjmNmVwdknNxu/A2hl4vtryjDKkcMEP6lDQVXxnNgJzyr+9Hp2T68d49+0
k+S7UGNqZOmlVYpbhW22F1vv29RUhTIPuLdUosOWkJ4/5iPr57sSkR7k2QMd
iVbCWTYZe00x/lVaqDadEyxoHWxWSGXNmZdp9hIxp6+6ySX/YDdueGdA4rTa
VtvETCkV0jx/Ga0vVmuznTSTIeHrRPQnk4W1lRXH/dbX8890pMJfuAkN7zCB
5JMuanI2Xwa3FVKgz3B7VpjNgh5Y+DTiiYPSOP7a+le5GX//F82T2CDxn7PZ
OwlrmCCt9Pvpx9h3J0YLYMIJ9gFnVmfynAIOIjspdyVZPLd0QRq/j5dtowec
TAuBtikhE6pPCPfg9Kng1HLcG35b72x3nCmuvaTNxKY5vR2KSrPD6JhQn0Zk
AwPaxIEaLfuwA8oW42/M1jgRqUoUB2R1zxY0T+OgPOn/p4H2gfLujc3lpKc/
x96dvksxxHVLqzUTnxEs6x5BqTjUinbicZZyf4QAkaXXPLwwhzOxLlPkZn1/
YWNWhMXpaKcZt6+IqGFZShL+OWYDjrKhLB3bYdSSpYJy/idxKg06Xd/3xXjR
3eNOVf58yQr9An8cnQMcciaLFTVAxPcgTFpvwDkw6PfMGKhrMkTrQeRN3RIc
nMASF7C8WrX4d+jUmIWiKGRQ20SMAVx3m5HECZNFrITOpfCnxC/zgYvhzaf7
8nc4T912KMKnDW4hWSQ+cliOYrXfblM4pRglE6nswK6we/vE9DxbGgUn/q84
BDTrB+DYCTuAq0REeApvQvL0U3Q9xLIYTQ8osIix0bA38H9aQ70JoZCiB0vc
9siC9xj5bIKbkZrRzd8rSudTrUOUlqJkx6axofJf/DgVWFhqW2diXoLCHK2c
wLJ+aSZMspM53+zHt8kI5Yeil66aXQc55KanUgZsG9ftfHlUTXfxtpX5n3MB
ialYh8DZGLWIKyostwfsPfLZ4hxEaX4l/AWZrCyNyh+ZunWZ8O/X6+Hzilu6
ratjmCdDuLeGUPhIPYKFxinNwjSyQnD+5swqVeWeCuhN02CEf5p4Y3e8LMR+
vyyaFxpQaQlCFiaXnOrHKUsLuWk+srnNjWw4E2wjWRzy4HOrjfvwTtkyJTP8
RQSKSSSdlPZE6xrdTcPtH1KiNXwM85MkqRutPnXi8ODCEPFsxLa5n9kAho7y
nhd+LnGBaG3ntZBF0sKDr1IiNjjD/oNZW1GP/3/2enQhizcS71F+g/8khlPj
l7qRfAWeRfuAke1+08BXT5uXTs4j9UI7JVlxkSadbDqtDcb/EaSYmA+6yB1m
OySPrCJ8foksnMdoAEfImeXJdWMcW3rxzKlYLn8AK5rJwgHKkzObIiOZHwhE
Mo3IgGZ+hNJY5pdVwznqUayGOFf6MagbTarE38l8Fb6g1ebsP97BABvK/Ydb
hyRxsz/OdAO+7qHkykVft+HVmsY0MdMFfwAmveEbpmPIRQ90DjciZDY751Ld
aclhmohpIv/sxdCsc+xqpNedS7kFVTQTJso1NPROxfggppUvTTxRK35vEQBX
GpVNmadLb5JTZR5jyzS3GfC7b9rAczAy7UFlts57ZN74L+VjWMvBl+TYXEuf
RuocM9e0ku2oqUGDhwp60O63Daen9Tknx0xZoNFM1iBfXW80foSNnk8+O8+5
u19vOtiACzAfkbHdsiEqIv9Y/YerkfFmG0227xxmp+UptUpxiJxad1IbRbOh
sLGItHBe95X4wGK2uHq8fxEhM53ZroPWREajF3cm35+qKgXLFHgrYfFx6PFB
eX7S21drGviSIS1+5duo2Fd8r8VafjJ5A1e0QIPzw+doqEE0OqwgxZ32lvtN
b0WebhrexyYtDW1xJ7aINwHnvMZ1SjZFuA4hhHwaSkURfZfqrIoF+NnTRqbZ
0ObaFFfqGX9qJqxtPc3gwSbQJOGnnLW3g9BPFN7EtYeLx6GBDVilaukzKUdo
aCPzD8dc4LKUhT/j9nn74UeFicPTulRZxjCWibFRseIgmNQKmjdtlLzZKOgf
fW/+Gz2zFayvB54FenLJyu6oIs52A46FnW4XOMqM45tLlZ0++GBbvd6qBtId
bY8n/2bp7OIA6Co2bf+OwJ+H0dKGbqKPCXXiXwCjJ8VJ2ta5R67msCApNSMR
XRkrCjYxm5YYrNIBIm6gTiYm1KLcQDs3BKVdkSFaLcJdSoEcV0N3Zog2n9ee
BnO73EoELyx5nPxRMLqAriUhrn/SbvA0SvYhko90qfOqBB3c+TyKpN1rGDzX
gTL9NYiVHZcJDFP8HzdWI5PG8unU6rKJ1F5i8UiXrvi4kRsiDObseOCKE/uo
72eaKrNPUL8k2N/XD2S29eCrwIDYalE55A3YlGK0xM2+cDtpwL8bz4elwdxh
lI3FrSclqCQTkgtay92fz8GioWXmE50FYfZS/ZqaIReR2JKl3QzmuPyfDZ08
UvtzDys1FVwGl6fhwycGPlCk+aD8F4Kk0vIKd5G3EN06lvoMr4Yq+1uNLhfy
tBglP6DH1E8a+jmrSArymkZRkLzja31blE7D38rY3MXyWzEGII+nAbYekXak
BVW0HCzTKAozzlzxRdxc+vfDG4H20iZZMy1jJT2wIMN0VUE8tfY/GAg2uVnb
t1+UGoLcs1YrIR1lFIT+UmgSf3XWZXqZxrXhlo6sqKlAQjUgR5R/JaFHIHvT
RUhhhgsD5EnJKxME8p6/Y8QVlvIdtKm+1Q5+f2IReb+DydY8MXmeZWYHZ5kl
7PY9AOrg2+JTIXa9v6t5uBFrQ4+xaGS9pKd7XfSrMaUvrpFIdGZtNRHk5kuF
0cK9Akh1wWHHYhP9PVX2Ili0p7Ab29kSTUlCawU8zI1SN4+CKnL6eCxFw+kt
CyLU8qJOxVn9TPpbr4WU+CuBsO8ng0lNeQJTQIrlshR/8R0X6Z8RnsDVzKWJ
L625Wc/T9FN2Vp/1veBEFjg39cNfk1jfatia5Y/GdcX92TTi9fZlM51A6r6L
z0pEPm1+OnLQInxLnRYx2lClSGmfYbDvYUiFA+5npT3KUVWBJ6Op+B+GZsHg
NbJQCASBWRb4Kz8/MCdGXUKFbuqSwKP0MZIa2ZMzVcQ40O+Jf+vhhizdpQKp
GL18/d8Yd6bfVAytwzPRadCMN9RDqgKoIpg3LZDs+FqVkYvgqRmsSstKn8HH
HugZ/l8uXE0VGZCp6XYKrEHfEc8TjGc7Qi5ZZeyliJunwjzWfdEJSWsdy/lj
UJLw0x/BGbKifbx82Ve2uRNcfTCk+PwQqFzGyudSs8cgyvRSt/kSVpm6kk+X
wnTs1SS5V7mqy91kpR2Ygh7aoNNSkRiirk8YBr6TnVJWqZGtRUBMWdzm7x9Y
QqdTKb4u0PYh17yChb6bHRT8UFkZjts/nvtwTTUY4+URgE2MiYakqjz5Iw30
/gvMvYJF5iDwxVUk8GI5V+1pnZPKSD1sMHsFmMYyA71g2WWCsVdv/a2FsKhq
kiY5dqSkbXzUMsk4anZWPM2EAPT6ATZtSbXyBHralH1Bcuj7SEMaXaKIv0xi
/upLkWYnaaD1g1IRFYPNJkap/c9LKw4rQLaR2o5AeMJ8MkaMZ+Z5hurQ5aaH
YhTJ4i/ww5Vnl9xlRzPeiXCAzsrR69ZQN00GBoI1ZJcosqQ9Vg3v8s9TdE7X
6SdgCYw+CNQpoAMWzdI+wvCGOwEHu441dOuKgAFI1zqHtF8at7xlXOGypzYX
FGg+fvdzHe7Z1/NDmxuQiJ9WdqEhBGj1Vm1tcIiDbqpM3uuvRg0yEiKZJTVN
QgEimVw/1aBGY3NisHYRM7bG9mKJBJfZ+94OaXjAzH3rQZ2UN0ItVdAf7kJO
eOu3bI6ixLcEv0JJmGXwEYri2QPNzIPdNVfcZZxhUv9a881IqHGnOQXocDNW
8dGPaAdlD8iShAUDV5+hkHGcI7GGYoYCD2PYBnddy8fVor93h1dEMyl+IdDa
k6EcOG8ldTt49qVEh3cQSTtX3c524Wq8NONQija+mlfoPoA1tk7zG0bxn/+D
W4qrid12wfw2gjvKnNiheKvQ7AGhoFY5y/yVXAH6APRs+1PkvyMoI7ubrZBt
UAgtoFq2H7nJNtZCJw9KuqXEZVDXWEKaMCpFZvDC4Bb3TVTRU+JfjVvI14d0
UQtjez4tO13Lo8m0uBPY0yIXMMCoiHyN3LfwzW6fmb0y8w7QqFmwxT7ONDx4
fZWrUrsv/NqQC87Tu8jsGTW3GElnMf7JXY+vw4yaixJ55wztXcKsYk9rHZXb
U9cuh38sYPup61wzE9qzD6C/87HZEcek1BtlremEkp2iyiCVIJBwwPR3N5+Q
wv5B/asJQilvWSku/f00RauOPneG9o11LBM/cdt7mPGlwUeU3YVoJKAG2Qt0
KyFqvOyky7x42ow/UThZUr9VKpd/hEYH/5HUfjPgGOx3hTETQmmWZnbYIF3v
99TVGIp171e53voj9bFRTqvBWKj7S6a2Bjy1bJNxZRjIlpDpIe9QIx/25nKN
FYvmOukCE0GWv2WEWKRY9zMoHgq+efPP/B3LVY5v3dzAlAt53DBYEdCB0GZt
7k7eg3/PUa7HQuYNWR0r/Stgn2rN/8u69l+1Zs2a6bzTf82rrfqnJtFw6GC2
vwLt0lqGiJud2kvpsODer+PAxUUFLF42HAVz49AYpjRRI4W5fMPJJmcbqazQ
EcC3i99B+4GoopZlHJrsNnBBwx72CGmpWvNiRLAyE7x+p/enHQ5SWXC6Nova
btI7CGr44yL4AJ+7qJr1ng+DKicQ4vgi44FKxq858gEi7AJcYYtxT9rlg1+r
KvyZDuZnFzApJqQKP71caCwMOjUaH3RVUflGbo2RP/3BBwHbtbvGh1OKfSpZ
LItsefBXoQieMekh6326YrbVRm/TcfK/ARBLF9z7L/5os9iKWKwt/+Ts/ZR6
OPPH8XEqNKmnU6ay+0nCK925TMWnIbJj3OiDrNl4M7o5IITKChw26nvJqMbb
Jf8jd31zd2XwYGPyPy096rtKY39VfYShyck41SG274oot2/AMrKYYtW+20dk
zBPyyE7Z1ehrvdZSD6GxaFUYxWjq1F08dCEosA99Ev+fkn42Xb4nRpk2MtQ3
6UViJ4gv0VOL70xK0hLC+dVm5QDQR1pcYP7G4h8wUjhTDXrSalMyT5cxKLXz
9EPQjUOfq5zc8xU0lnpj9S3Gqx/tNpbtZDb2CP4o90XMNcVRZ1K38xOfzO5J
bAERsdvlLF2qGmZ1PL3YQPKtQ+5S4TigF3lV5gAIjx1oEosPYb2KfBcXagEx
hWqQF1aXl9Ug2CfutMgKHRllO0eFgssvnrvI6tCOrGEcPCYxmH1JBAEPvqaT
GHRLagh5TnuaaojW8dGE9u9WYiv8w/nEjgizqZcw+R9wvktiMbVa3OAlfMyk
GVV/Uqjr2czfYLBfiGkXsPQvjwdsViIYbRCHPiBtpNdFu9g0y3+slyRwlTDA
i3dc95ljC9GWoKExlfIJabQOvgsi2rVMaHOQZO2LUTHqLIgbztP3LvehauSX
NqwlJ292qq5i2ncb5/WHDxemjlnueZ/LZ4gj3SrNjcG7OcXCkUyncmQSRgTm
+xD4Z1JT9p2P4FOwmWW4laLNhEgS83RhbS1WEZBtzIG3IDN8StSEEPGSik8d
3KkLEsl7N1dw26XtWyRT2RU+FwuHs10Sj2/mgW7NaQovVSkHszgTFVvZDnGF
jc2oVHaQdwnr044c7tLkzvrBr0+qIcEt73DraDpJgvO1GdhuOXHzUU6KuveW
S6AZ2OHAmbX4kyrl8Ng72FGxS7g2XAq+VJ73NoT21akeLOb13rf9tDpP2XH9
IjpInn8Uz3ipv5DHUFQRawtmi97i2d8G1uSV6W39UAXCgNqhN9W0c30dNuZc
xjInb6GJz7nin+F1zHhSI4y722Gnz8qLSPFGUrGUvWSx1mkb3supe+vYagUH
vsvddmJwb+/k6bjLc5nG19dsT4hIDuycifGXUWdoMskX+iVxaGget8WWLf/+
+9Q9XQsUGRbH7XNThNIObKsdvpnFGh9Q24UTipIe+YGGGg+utYB6XsBGd6Pj
Emxflzfa91UnGpny0ivnaKg3O9DJJ0lmtxXYUZO3VKs7O/MzJEwMPpok6D49
03+Z/XcwMexC3Uwhl+0MHp9TnELr6j5pugNrbTOqEh/lKCpKSO/uAw9YBsWE
qB3nbFHHR6UfZv/Yk+El5WrPz+zrEy16BEPqsT7gKSm8vuFiYmtiCMYjrE5v
tBpgOVNl27VCFYkegR8wa4rC/1Op2GOrtvSTLpGf+R7Y+KU9o0fG4agQq60L
ACVdEiELH0atIXQqHmnFX7a+D6YPhd+BxzUa05unLqnxdRAHAW6D8lata9Ad
chOGBIJaUe5sITGCLn99nMyeR5WlJXLOukJOu4TueV1WCTMo2r7BiOMNy6aD
4D5qoyIpZxT75SGzkVIlLpBTebow3+i1NEEZIhqpBajeoWLTPU4HoQQaNFaB
qED5iNzlBzBqZ0/E+6CGoJMydzk9NKfS15YyRP+aqjQKfWBmbGdc7zTkoe9n
1FlggMbnDJA5t2ll+uoqR/gjTfQZQX8e/RM3uXkOEFIM0g8oM5njoKDXJJQD
Vsncfibep9Xsg2HAhJeeNdsFE7m2CQl5QzVyCWOuzWo1aWV+mKEFpG82G9OP
T64+EcQeHfdaJ2kb6nPxpPR3Ah7umaLWaarSuL4BciFC08DzlgbbdpJ/D+IH
QUEKXmDFK9nsNSmGdCmDlgjHpjVM7+vns/DYkEnJvA98kYUPEb9ojJlOVQZP
dx7xCxd5W5XeI0sieXJSK51MXzqmzISs4jw8xLTR4u1ixxVJtY6RrQ0S6JR8
N6Rg/3YR3v4+w8IVofi+zUC4D6YW/src5XkbADchCIFM4y895rhst2gQBKBk
V8dhxLA+vHq9ehKS2rz2B3RS/bqRszoTk4kN6TtGVwOrfT4SSaDGC8+rJ80U
L1XeJ5Kzs/OUYsDk/bYMXgIxRh3dGkMlxcrYJ0KO9263zfVNOLFJZUEIXBx/
cU7+a1xVYLERBmf1Jl/afkw3Aas7OLCeOlt3KwRpH9WV5IV61gBwcQN6Xqus
8gHl1tjhczNS0W8sYX9LLu+NJL7Fo+/QbATfaaYhqMaB4M+GSE/PdFiCjx1N
vu1XvlmMJj75Fi6VkbKFtW+BIWGwPxjfvwco0KhKZkGiCB4NUWLZydrkAPPj
xiHASs/hkaKlb0zlzfsAbeiZJdcoUy2dCiCJDVF9lFWaXhkywErIrF9V6zuN
PMUBQB8LRspdVoIoVBZC1Tj1/BPSeRmazm9KrkoOmmgt142p6CU3UudELGUq
JhdLVBFs6QH7Yl7UGvLKOclgk0GUXOwxekyOwSI1elE4u1VLNe6t59BsyWWh
SRfAShR79yB3oKJjxjKkQeXohwj40oq+LWbDYxQoRTM/wjEXdBsdyN6fqBQX
hs6PfZdKF2ORcZbExGi1f7pljVM6JdR+GuUz8eWvc5lPMF2JIsFwv8kH3TE8
aliq6deaIeMSKlcyfk2o0RNNHmSh/EQlwazAmi0wP989zM3xqQyEpCpK0ugG
E8ZPci6FYdJd2t0xyBOFzL4BnMFVXu00bk0AovdcbjQGoaKCiuhg1I+otlsB
F2jNYYwQCpg/ObVxEHGWCqjWwCu7bkkj/nD/ZO6/ANOCvyvR6jpC2vmT5VEu
R37J1RpfQycmL4+/e6GqfDcBm6F6pgApMfxAM5JtzXTEfybLB0V/w9jgVPYv
h2tcqhzaXnJtETwPFNPDuWL9qzMQvE1CtCbOhWTsvGNAMM8g2aNa/m6UQCY7
ZlEgUSoPzChlaJx9s9iwwbOdmUcOSijkisHFt1+htfL9YCtPNYfTnmErDSlD
FMomwODfiolgq6w54fVmXmnYyjKzLvLxH6G90jk3g7NfFQOZRjs2Q0yLw6E8
798hZT4uh9jVQjgkhZJK0OwOpi6EyMA2By6UcVd470VlHVABUPyDDaarwVm6
QgqkFJJ3eJIQDZxuJhxPumM0ZCr+P1ix0nsTc1eWMm5mMjlzuz6KglwRab31
DVv8Fu2jnwMgUKGc86zFv0fsfO5OklARSVZRq5Og4BBwgiC5A562c+1RUBYJ
JnYooEeGqCf02s4BgrWX34xPNjE7egBAOlhUO1nu4Svm2TOwHCkCvfUlGbTo
Fa2FzC2WlFZhCA+KW1TLOVFSo5fv1YLkMCFOuax453DIHahMWYwrol2mXM0N
R7LCgRdjHs6Z3FF4L54MvZqOFhSuM5140p1YL0T6SK18G1RHCDGPFkGDC2uC
y8AW2E0+4J64SJ2t9y2UpEA4TZuFqU2k3doFQf1AEQVqRQ/8V8lTHdnkUUqx
fO86oOS5S2vMmPkXzmgvY1CIzKGOTnp2Z/6+6p0ehWaOjyaLObHO4XiSh8uE
tHhVNKxIJoxN4lguE0lxPUDWM36QSQQ5rLYs7VeQyOewgaUgtU03WCm9ACcV
UQqvycLSe2U39Bty6z+thUk1Z82HOFAvU5pODkuz3GoJywSy2MTDP6daY6Mp
2jyqfRiCkq2wUUa6RefG3fH/ceg85KT3EwTNcDBtCBw8U+VtNco3s945wLTh
Gr+f14eqqhA1BwnQ5vgkMDu1KUJeRJOw4xFqg0JNbrpdnojd3Sg/OcSdYG4T
bbDx5nNR+TasliM3ItSk0PWadOsFwZUQThyib4IIhJdLQxId5CGKEm54MtwS
YiZvW8r0U261XLJZ7Id63BU1wtlOd3AO9l0X2pYLQMCFIM53APIlMJx/pkQF
XRlXJmoq9GRaAGIdrjhs6Zw/8+dEgM0PQuQC7JRWiyIwTavgpz6Ml5gTq484
2ROLA/JQ7P6wyXd71T3SYkkKvt0wImeCX3VJq+Ij9f6FOobq46zEzpXuIvJn
JFgGjsthh3MirSj12GlGpyUNoxoX5mh0sazuuhMEQvfBdRo+a+b3uIp2hb1v
jve7WxVlZKT3b0lKdgrZTz1vgYM9+3bGyJMtLP0TXoz/RtkARiVklYpikZgA
HAeX3PXo6aBlbULhfJzxl3QitPQLt166T0k9tB+IsdFR4yjZQaBeEZQhIGeh
HkNDhae6bXnT6YzSmokblTf1SJUgvYynhWSkHf0SRx11j8ha0VCZwPVw0EKq
5xBgQtAg9LIbZBMUS5MbpYa+sPL9T5FxImRHIhlU+1Mr0Z4E2zySuZt5e/I6
5MoBEao4Cy2IJyZkXI2UwWMpQjTqwZGAOHBqex6KHuYTvcUWwehczce3QBhJ
Uc946pXk7GhYKHGXNiimkRtW9jGz2KFSd9/KFlu8Nxo94uoxU/h4sIrGcLjc
AMvkydaOWFORV8gJdEcYoO6g1zEm4ec2G9haEyAe0//DXDCG8Qlnf2tKNBVb
xaVuJVZg84Smifu8V9eTz6WfuW4WPb332SGeWStYxYBlV4vPSP03yuQhWuGv
JqHmkEahG/jYTs87rX/NS2HiBtP4T3EJS9eTXsVFPDofzy3x3ZIIprrinW4E
fsLfQqnmJPlRv8hy0TAj0C+zAjejiA59eJe5ZIr1JYL9gZktVPoeoJdJu6nl
QZonOgmbs4di3MIsKst7OQ7y6SWjRK3Uj+A6JJQTWWULzRYSVS/lXljinaP5
Q84frpG+Ea6qEeBtAzuAhftPpt69OCb1oCiPAeGoxUR+TQwU2WBH/7UjHiMn
RQRc2E96Hu3y705TMhI5WTZUKnz/URS2QfYd9UKed9F+sJdEkxUbW3JmG0W2
sqWwLC1rMW6255WIuV2tDyA7yUGK4ln+4dDVILgFBsWfN7ZjhuZ0N0pY2mWk
9dblQE3f9PC/qid3/41I7CuiinSe/ywtYqgsmtMIXr4MysC3/nZcFJfKzhLb
qcT+wRdccXGSHe2KfEU1i2U/8CJCkv6L1+i4G5eigfV1nhLxQ9P0K1+RzUEZ
Nrhgo/AeE+TM+FOKHu0qAh++bqYAe5PB5bQ18RvxLfLr3qCjNjYuUfKrfuMZ
6IeMX08s/211h+fubDC8op2OXUlx87G1dHWbcmWlgDR04T7CK9Zs+c1mqCgz
ZhBEoBiUSBtaeeHK1hNEkGGTmOnJXN+X+W7lY3Kkw3YwAEzFMFdgs/4HSeE4
0F4Haqpnieddg/VKU5xCn4gZOTIWM3vvCZzJKAI5qd7r9EMYeaA+pA34eK0z
AVuq27ebhTlaa7SkjJBAD4sA0PvyPXSQtnd+FWsKglNq9DZ51i+xzfiA/lkN
E5OAclbzJcMCgOkQ5zfnkjggOig+YhFsB2gxkGReaBuKFNwJPM44Xw5xVwv5
SVBQ06BxQz2/sVi/GjDnVbrKxxrlR0KMmstMCuRRz297f5u0FeG97vlyUzWl
EQVqTxprXNLJPDqySEPgw8MK66r8N82Pwni4xiLCj1HB3kLV7uqhg/6cXk6J
k7Qrzy6jn0ckIUxfJtDA9Zampq9AuYVWTDGRq9OJYoK+G93DsbNLnFCAvjVN
2kpZIkeD94MGuxv818I+x6jAEuKzWoRaef+y60iwG3xkNkwZ7eEqYH3974LQ
t1srSBlL5WerGwyWo1lNFPD4VEJKj/TXIUXTHF6UE69BStyM2ANqY49djMDe
aZNzWJOleDRb6IjzpKfH2ehAarf2H5x/Xk57pNymgGV2vBZWdy4y8Xo/cJ+e
Lwru7KgxGknLNogHXSfjTKUBBCePOzxKWY8PYR+8yaY6EXH+Kj2bd2Ka0ZIO
PeeJJQpbm9STqHvb+6Wzuvs/cTYf4/klYPI7Ii7DgFNnhd4zwuX2RyZLv9eF
QekLZsZmTsiAf0GQkRJv8xc1DyEnw2zRXPUyP1XnGXsX+3WbCPVz7ceOlpHd
5h76q1H3E75InlFdA6oeZlSkJSvSgnrI3gJDAN2l/yXslWX7btqzd4Io90uE
cdZDhWnRewPLx+Ocm1kN+Mj9vVwOjjgKzlQ0lJsYYeSz+cfs49jAEpu5glfN
SyIVQh9H+IxX/SYMvqiwlOnp2gvl7vZa3c4Q/lDQjtYxREDOnBBPkBeWYjVi
mwfXxNDDzFJyoQOLDHnRaxOJCJ6/3lTL+uf3Z9cC9WWmaUYoYz32Yl4Nw8+a
8I28xLk6FCUmvDg7OZ1QRQ5ywzjdN793FrcKem1KULGihEGZD8fOL7IhaqJL
K+Nc8R4+QrgTafaFam/Vd5MJCz3oyMKGE91zhgvWpw89GkyaTQe/L3BBaWQj
/+h2n7kN2ZwRqVjZ56u6VFaiQM9KyhdgoH9MVcYFNTR22dFcShCH9rJLdwjA
gWtukRjf5yYXEpkL/OQaGiXRNWoDr189Qfp9f5HAg6ZVWFdn2w5pg9pXxx46
jLAD1k3Fw0MzVxIOLY76p+MnXycZnX/wefcETQRU0820XtqEN1kgAmBDS5Ci
jlmd54w1TgLY0vL1OQdW1pE5hmJJkCFr7wWgmyXkV+ibfbBV8L1FwXW3Brqm
ps/c2V+EXIXlEPXV3cqigCqOhn3aA8+kZ8Vfj3Ll5Gek33xQD6uwnnZirc+s
KTFpFBll30M3Qeo9uAr0ncfLYTLcvGiDjTcCO7gRU/XhN0SXR/w5IbAFJmkC
5nlf+FdLkGBqXFLckAbPvX00a+x4z3RfDSpu87nYuyVjA5IwRezQmoXNeE4S
FBSS6+c0b9O4pc+Ii7G1erPodtn4eXQursJnn3Hs+1HGgQTHTl3yS3cqet8E
8lGsWzJPXYMZUoHsHT4U8+vX2ZZfbbeVc7ya7Y6Ur2QhNDWvkfe8vUHDmZ+D
v7Dp1PEZK5Bj4WeUrmZMUtvttPxrSLzfaoEz9YSjSFGKo7SqNYLfqA6JGr9P
4z5NS6K/e47AtfB7aa3slDCkaDNzURLiYX37bxiG9WUMcH2gktbDti3GoQdM
W6fNc9tkAxP9EmrCucqI0wVRFfk92iFni3RHIfkBUqTtdEkz0xuokkkWoL42
mkqax0qLYBvBIZ1FfZH5dajEEkl94wl4z1J3Jg2cHNFxoB0uAhU4DgGhmwOO
HUC+hVVCviPOYkaFm98436oP1jL+0SUm99eznwLNkuj/V4QMazZcqmx/XetK
k3zU5aUp/CFpVNqBt707Tr5YMr0qUUQeD840/j32dmYNPT0TUouwB5fOnll8
otRpPwAs055LqtrxpD+Uc4Y6X2Zc6dXwvtBNVO7a3ymzUy8NMy/E11eBPpnc
JPeNYe7bv2Farwg8BwXd81RK2bQ+1qVeoDmdFpazmj1gyC6rA7P9rHczF7lW
6GDcvBLNZXwZ0CFzOJFt6bwOo1fZEuSKqbfacV1XS6EOyCDbCY5EX/gNBY7L
0Z3KJeliUfwCdqQyyBKQR+F8Hhcz1wOmFpGdnDBTt028WdOO81KoK/7vysEN
7P6HPT61zGfAzy3AMSHEf8X0h12B+rTmghI87k5oxrr8/Nl/gQaOXmWHJR4x
QypYV/f1gf7wClJcIs5EEii2yA/s1HYVdR3tdYj3PcdHwnQA9t2BqXx3XF6m
346aPjz85snhhb3EiRuTn3kuttVsRO9PdEikAu32VTNQKN5u126hhABj0h8o
2mBZgHTPByrVHdWOqiTJFQN4+S3sFEbxkqcBBzYw1tG114BxZaJrzr7Y9fuF
kzsmwNkuS0L/xwc0hQtyQvBU+wEFw/ybC+spLW/RUcQf3uzx2Eu31SlSLcsa
UcUN4WT5uXWZebwpOO3nL778x9WqG3/Y8wm0i3nwZqGa9aUZesxMb2PNObBN
cOEsKWA5S0AjgzMQOfyJukjnn2JG4AFKDpR7CD9lH5/JXa/xRhAGzxynHsqZ
gosDditHM+G0s6j0Ieh/PGF+lR/tHE6lpYBCk9Uv56ligUcy/QeWB1o3etk5
r6hvu7ThlRS/W6Vk6YMQhC+cYgMJ5Sch+HZyZIweTZZpZ+0hHE16XoB7LuFQ
YoVoix1gnfoNCUhVNWpJduo2Pdxrwv5CnNO07TxPja3OdwypL/WUMbfFaIwl
Svj5tpfE9q57HjCVTNuOdz7o9izxK1wlq2AfhwqP1S6nldh4bussFMtCK5If
h0SWFiEhYZjKXenYeu8lzIy+gmeZ2qbksGXgAK4ZoqRdLqKEbqtXuDDZtTL+
ZIB+CYnz8shlDw6P2srbiF9SaG4LzQaxsnBd9M96Xkr3xDG/2qBf9TMm0ylk
XpQMTfIJ2oLlC2FJ94RWXI7ajXcYm7csFKct+jGAUANxZcmxO0Yh7t2wjJn3
/JfUZg+8BaURlzs0avgFu5xJ0n57vBjuCAHcJS/PutxKoE5Kra89SQb1pBKk
hR0pluv3EXXjHGSa6UCkzJPvYpIPBmY4s9KWwPFIbjSn+AAcOTvW6yoFWD27
dPY0yys5EdDLL97uc6DVPNI6Z/ovpe8q98AZqQPoQiey+r/pgTJhjUp5HUmd
UFf6acQJUpqQAXykOT1xpqsU/jTVttj5+eoCC0swwPV14eIa1BTtqq1N0vTs
Vztf6Qrw+fR2iFFrNLHBRxCLVCyQRdEIZJSuj6D3MNUjpbTYjLI0QKj+EFzR
kly+hgg1rcx4R+jYsF5Q6Cv73jmDk/27DW3j8kik3atQZHVx5wNaIlzk0g+c
5YTu3gQxkXiCVJg1BeIjbUryhLZqlRTYPXM9PW77j/CVxZolbxpOJKRg44nk
oLrMM8RnBMDy8f3GNdGLLWD5tbyilsiLjQMQxpTiOGz4ulKqCVYSn7+JYpzw
+eS+M6+uddSso03NEGOry9Vmy4j/0i/J0bYF1jqnPdFWMrx+zXqONBp7WjKK
FSUJ5K1+4QmE+GkS/oxhIotTZOB7cGcE+Nap6Ihe0PS7V+cTyT0MIrbV0SU4
XOqJXyaWz9gwAUpXjbSRLFNinUCmsEfGHPz0uweXZq/HOqbGEE6QY9OOMh7Q
Y+aCs1dhMhewaibr9fxGovcLbYqikw41HS634k8Ap32QiqZB3OV+mZ8xlS8d
MPcZR3aO6758N8nNaPoynFwffXygVzJgqdnkx9MzRIir1W6+axbjRyZsJLK9
aNFAiNir0M5ue3b8Odx1ZJ7JrEK9/Cy3ZRARV0HVXW3iQTPCn2NNyb3fjqGw
FHs1mJJUmxq3CATgLQmdzFep/2PXgy3qekQTej1YEkqrE2Ssl6A+Y08Nfo3+
wDwYkvwtwEYY1hBXPTbPOGPJfpINW4od2Xeu9VA/hPS8g+P1bcr6Qfp7m+vZ
oLDnZ+XHDRF5RpC2RB3dYdnA+rFB3YR4qnsCY2whXMTY0DVKDnkgwx/OH4dI
uH6iqzM/FsSQUCeNrZxFf4QDrsO+lnX1RkV6R7OLG4OfPpOE6YwX6r3ynVaT
jlKOUKkaIzX2/fMyNRweXIUq/wUfEFrPllXwUbcuOjl5o1KdB12P28N9vG1d
0yDuyk91ghXN1SGhCliD8+cWTsn/vxLzeGLXUtuHG70ZLewnZmsp0FUrajDS
zg+k24ddWt93eCrzR4UOIHb1PfnyfuzZrOW0M5EoEhEFbVI1YMwP1RyQtEN9
TfsbuicAW5HKwMel4fj1MDhTXo1RNvK/BVEmdFutSEuOO0JLhyZUfW1G0r2B
pGWNlLCeAYTRkOrFH+cjP9FF3xV46UBrIVA/ZgrlHq9RXhBafuke9bVbueqM
P+B1cgMULE74GaBFs8otdLhkrNOZwToIgTyzm9dQZVrUnWkddjFba4kZoMWi
eLZX/mcg1neURiWqwZhbR1SsU2trtnP8NgXLIeMuhHafX138TA3YVZbJrjIL
NnkMH7GQVrdKqmlcsxDwDWh+FMxKqvPIaC1C4QHgGaK4W6XEkaG9tJeniqOW
XRnGsVC5WQE/y7nXWqb0F/JUF9e1Fk2BahvwzGZoisJ/Q0FdXPd/AbybemlA
Hrh6Yc26b9e3JZHe1NTGfbJbCo3kxTz7USnohgWN9/9P9Ilp9wuY82vOOZUr
FRqNidX64f/pYMH/pe/3AOhWx+8iJkVTdovqa38DgSbeHF8kZNmDDUe5wxfk
rBFQ8a+5cjOk7djfGxXjn1cim0M5OXa0JdsUD5MrLEFmrIGTOvLv3iufcn8r
6iMGw/GSSMKV1a2a2a/JEN/r/O77Tb/V6poUyBsJlou7ury29IHonOM35JmY
i9KYeoEwsu1ZHSofy08bSfzYCLjlqnIDKvu69Nyh/Zi9ahAIPCHxZ479xbMU
ydzDacRoxl9iWQJ6lvf9cM1l3UzcBvngFAXOaKphjUuhkFCsP/LQit7nQlTP
FPBYEcpDUwdvXgBd3E2aDybzb/eVwfExVFI9CanzZfC0RTfWc0U2xfiKrqY9
Ng0Qx9c1NpZ8sayWWQO+lJAUyWxt2MhkHfCq/P/g1CtfbJG+fGh16GvQaiE+
LfdSl+x69HZiw8PLum92G59Np/X3mb47elzfOrV1LM/dQX4iBh0JCNw+uYSI
EORGb1DONXn6vJCECiTX+S6o1uis0QKb5h9aSBORZ626Dy39jRG9ZPp4Ghnh
Md9Tb0bCL8vj/BEPpJQsa811DIsAYL325Rmo4EoOOkG+oV+O5CwkMN2Bi/ZK
7fxt/U4jl8Q3/gKVHcvmULMXsjPR6Be/GsEyGEX6eofCuXiqGrJdEd8315ea
pNPR2nF+YNXoYFmfJp7qjYwaQpAdMEEHC8GZPv+La3Pxln4IMaC0dSb6eTYf
2lNFJNNfamkNzrLVjn7Futlc3YP5BnGAVWcPIyNWBd9UXSKgYd51qgwQdjvr
u5B+s8yb+PtlXWQzJwYzlQRh8YNRNvQTd7HJsapJuGy9Lp6D8RoXrNge5ENA
Q9Z059AHxl3shQTFNpXip1EginFL86gF4pGBbfqiDWhIuHB4QBmgv1kEQdVs
ohBgSLGTcjHTiN+8jUl5+VZvBZAhk6duUOZAVCcNY2e5leDrWCsvM01Y8WvR
AhcjO24snhsjxpCPQvw0Hag7RrA8mLlBB+sjf6e91RfxG76kG2Q0Aiv7wI75
NberhWMPw0Vn+UH+m28eyyM8EiDY12XU2m9vIDinFIpTlyYhu+1AC/l2OqWV
rDeH3yIBHHDW8Dc7Y0GTvOv/t9C3fAR/b8BCILEj0ny0qZmiWJXILmp9RAPr
QTpqdjEAt4WP7Z4+90iJf8aiWspCQG5WdCitBJvjqglPOw6DcugcmkIzIHs6
huFLDHp/N+t8uovdntgyXf5YZleRp3vRI5eHRxVa1e+N0J5RNQMWXdiaRYhY
sYq9IUFO81KrWplmbRUV6uHewMFH4LqKheGAfQpYY6Aqh7D8iNY0fHBGQeKx
FTXpsnHnIFDLJy0w0DDSk5ORn1yznEttNSDc0VKo0uekjZYHDO6hcF/lsYAr
r4J04OSYIOTG9JBPv1EP0bgYWx5QMgI6pRI3yymjDz0dpg7VH3onTphSiXBB
s4EYIpFtMTJvVSSDyWmcQw8AegIrPqWf6nQH6z8wfyuTVj3HRu+KTjjMELTG
VwvLT0xwtLnRh4DF+IcH5RA0+1+CKhL//RpjwCTZnyeZoluxFksbsDU3cyzL
nxs4PCd2r5X99c/ScAAHAPxkNMNmTsW+pjuczye4/yiRsXB9MzEvOv1d/Y4Z
eyfcm7oAfASOlGo7G/4p//EObyLonKuFoc29xt/CEkrVqb5U9cPi3o5mlctP
reyvIVz3Jwibt5nsnTj5q+xT46geH9Ys+XGKpZJHN8Ejp1dTXMkqhcHW9eiL
ylKK2HObH5tJKn6a8jajFcAlyvL68F+6FgTTloeny3939qQ3G/Tr/ixYlouv
xvbZBIxLx/5ZclV13q1FFjAlLqf9rXz/yzp8PcbJAFhxYaqfcgeyZFDfRj88
T2BM+XNjdcwTERq9qo1kAEJc+gN1eUFbvjv2YpxXgyDBMll6QWP5YGFFxrsD
sUPEmlgl77RGqIDAm/EfhctUv9WZWpe3SksrDpFzITHq7xEi72K/B7MeB8yl
Z1m4WhbmTAX9am8/yG7JnPvTmHAlB30LXmSs43JSBxKPBWKQuIRoexETimzR
rI09krTApg6YwmNfK81D3fzl0YlbX2k1ux6c9YT427ltCv6BYOsDi7jw2Xom
rKf075eviipg2MB30p6fraATQ06fVP6iL9JPVarLTBCBW1JxB06wcHCIs9AJ
GrHf7AFDk7pSSue7T3S0cUg4ENAV5Dm2j8RXZBy9dEVHU3SlUIXbVGm35fWq
q/4Zv/potL4IBDyA0ZeoHH9J++3pAfcSmm5e/zDHCxu4y48mnPVRWrRYBEDe
qg9CDWRO1HaSH5e/cMybRWfO5X4ufj1jC8QFG1fEOR+45dbdaIaqmnXKV4hi
fkQBs4J1q/EGejgF8PYiP7Pl+fWUGMeQnf02lkz4SIjgSOhWGlM7SSZjFh0u
9e1wL5vT9ftLMRmupha91Uk3insqgjxyvwuG1UdxXZ+o5/X4ej7KSTK3mvZI
ipB3L7Uz09nwkgCzDB7gltKQhqTW8PkelYRBgdDVjGnsltsgStm7oCYmvBOx
Tip0Vj9V5Erf3xLQHdHGr3j+NIkH+GGjDpOz9DcPhj80XP01NBxMIc3p8ZpO
pJAR7rLptkwD9IKm8bmEQs0IXbEHeuue0BcI9+xOF8yN4hmmLToHd1MRNYJy
o5heVwDc79vIVYeL0h0v1InV3+mE+K7KdLaA7VT0RUfKWx57K+51z76z7gT4
22kmJAsxziYZ39ZWUxHaITHcPLE7M/HOGVGM/BhulXe9t9PTm9dps216YYfl
4p22S1A3r6l/UEgSgb4SCB4F8R09SYMOtuL8Jdu0Ec64kDYe9Ln9/nQpupgH
oH6si2zMVkS21dA3tN6QPdAMiE4FJ++wZfJcdJoUx34YhGvILey9+XxlHwbW
EetS4h8MD0WSo+PmV66KK+7D3MtmFkCRR+s93wn6jowV0XjE5jBHol0nMSjc
4KZhup+7yv9HRvgVxFV8r0CD0Cp+TH9hjeLzWdaj5yhTpDH2vcVKezmBqElg
mH86MbodLYaBr4rWh6FzPVUd/CDcU59lNfWPJuO3V8voZtYBw5JLPUNxeaUT
0W7MvRfFLXESG1KZzQEFCjtRZoLXsk2HAb6T/dqOEj9a5VBfTT6COXtV0zHo
rGDdiWm8E9SDDVA+/HS5hShOnl4Dhw5nPXpwn3jFT//KaDii0fzuNxEmJEvG
NC6uQr9fpPAeWjFlgOsIZb2AoXaOoU9EHRteVNQwk3CNs+uoX4ZEyk91UsCx
z1F+omV8KoXoDqCMJ+bbgxXqzH4IGWRzHdlPNXa4Tf3EcEiNYZKSovtKW6/s
OoaKqglQbAGxbSZAOt1o+rfGgWeFxPM3nymRDU3pq/P6DR+dqiAjwreHBXHn
knrRhamooGI43+P3a1rBIvfkg83EJFd22Mevkaso3Z16hZf8cpU7+5r5PWy9
WNxRDc4bET0bj85SpKOW4AT52pYqMbxXSRB1FyZ6YpSHAagqBNMVJ9NPxwJn
u3lxAzIF8zfgvd08E7rO4r7RMTb8DRA1SevS1nYBf/tQF8trxT1H7Q9aqy9+
n2PqOSjOfsFf0KM3QPm3kO3Ihfq9asL11OP5CqB6FQvigdJLx99f+ux+kElA
H5ww2n0sWWRsHeTds7OqzH2Lvlmmtl2CFnjiLQEDExmW8UiLdKGjsqCJbaCl
xOSYhxZU/QMnY4iBCMt5Y98RpATdFRZg7W+IwgDv3GKI9/ER87TYf0JzdNSR
KtlL9KFdanlfVZx8zbjwuY8Y5GYAiwQmoJ8ubr+y7nn+267UCvr/V9hMcyxv
Xu8PSQTedg8O21F8EqDEHK+oiKxSq6nusGQ3BJSMtmb6vuDtzv64k86na7E+
D69itU2Ts2KnCx1tLVy7zPAlN0BUA0iCkfFttv0suBoXjF8y2p0RY4cbjFTm
P6f4bshjLJjafYENSsNzJ7/ecS94YQOPnVAcOWi82ft7WtbkcRVAhl3VcBTg
jXNOgQHrDHX+JFjjaawIb7cFkgrdFfBWRaTuoX65+9Em71vXQ4u6aqLMH69G
E7y0XDFGty/XqSLohmB9AUMFMdNtwPDOg0vLGBkaPV4kQSzjLr+Z4fg2aaaH
jeQioPEQTZw+YRwJANoCEjmQjiI1QH605ney6B1zvxyTMsjRYq0qA/VCMRXA
7JlONHisEVh1AvnUNETNDj1OiRgzVze3CIJy/ATl/MwWytbCQZQat6J2NBYN
IH4WdJa0Z80JS66i2r0y3BCsTSdih1pEJOZd8ygU3ah6Bl+N6kNK9ksWXhzg
mks6iZ68R6Ga1vdq1cvAXVqGa6Xu+FOc90jVXgqyS5cSZ1vMSiBDxNIMtfcn
xltPn9dWxmj7oeyOwbPMsUNkwLOLCxHrPWYKjv2pIMiXSCrQTDO8RtAIOLeY
fw6wj8e/PaDN4ervk2oDZHIWUWEZyt31yhcGIoIGiV2sEKjESaI/wJ4o52OK
lSmk1IopF/6SnRdvSG96CLcjpIFYaHvRUOHXdHoKOe7os6zSMfwplCXtx006
Zulh27xCAa7MyJK2IcNnM1xvJZn8UlYwJHbyY7t3VNdc4Kjyrex4As5rwBjY
QmxBJit/NnqSb2ZT8LNJHYzrsV47A78BQLjvPjQOY+N6xt6mKq2vnYJFwclw
8pFm9I2dZTsZ1K8vxbvk7bBPKqkIXZ0zkkguKsU0jlk5jwZTMguiubloy9ZD
USNUKD/r2A+iUEbArRKTrRjG+pt2RRQTH4HOeWN8sHhwOmEbnyXjslinihM+
YLNmaWUID72KbpiSdR83MLIuHpzh9updNvme7mTQOVOOVusNWux99lTQ203n
3cCTEdI65TD4dt+Fk92vi8PAOd5TvQ3EEdng2QfkmS6HMOitEy4rChe8WPKT
hBztCuh16s9A9x3xL/AxrcSMeQuvDfIljkqbn+DHIXW5aZOCsN8k1CNrAZ5A
3On9xKlnODpBzDC94X/ZYY5vAIi5N6nQkmvhv4MKXSpoA91XFPVCQdMevTxt
dblabUerqOodL1RXR5usZmlQr1wv/S4jGyOWhyOVr+fJFATf78aHPbLDtI5h
AEwXakWEhGmQgEnrNfIcmj4+MC8ZknjzDbELYP3JoMdcW4qohTKdCYETzvxo
6UiWNByPMnV69iovPZNSC712HZxrl8G3wKN4eesNw4JKiXI2RzdaMdMKn4BH
/T8OZXUC9mxf0E7Wh4NRJ8ScJKsa3rkHIo2VO8GhZSce3BBpUuQkn0cH8iiA
AaNOM4Tht7+Xhnre+hF6aqWDiz9cmqVor1mFevUUMDG7cLlDDffzsRrVnHxi
/ni8YN8j9217T2TQuf0OdS1X+N+sOaY9940PyjkKDUAdQrG8HNz2n6EAwf0t
MSi52rKOOvFVHsZejdAgUXpJB0l+NQdh5PCWT7BB5ZrxzAX7OXkA0o9Zy2Xv
Ie1RmgUlmZlfpyqBjWtklQDsL6j/PShAz6G/RyW70+cqxj1YHqxWRrR0JdTu
9ScMKnYXjJ1aKOzo4mCpEMG3gXKCLZ2sRwuYQMnJnAQwpl2AGncJcOWCE35d
t+NXuDVk2JhvU60Eh4CxOZggzgWbgKZ4kcoulwnS9/deJ2bHp0nA2ZWjBdFG
26FMcGZ95Luh9gf67EDaH/edvVDu0qs0nAhgYbLJLXkNdzoOA0ZrJjRelHVz
YgT7y5svdPLU3412iXyoe+sxI6kldFz5PRXjb2pGr+OHQxyw6FhA1UhHI9mj
10aggMy/E4BsqdTPoCJI9igwFCRXXNVbb4VTT0U4vjDxt/ZKg4McFPt4Znwh
OtMTOXlw05qvCRSg1XoGQaeTeZpxKk9QOsEUQIR7Fu7XWl8sgxIBbX50QA3B
qhN6eDrBZQiTGPycdLvTiyU0H/XrmOmh24e0Ue1vHB3vPb2s00KduYk0OvwW
rcyWCQW4A4dZ4CTcJdH/m5p59YV8xHj5HN+qgJvbqXFEaIWaw9YMqhWES/gf
wkqWZhf/tgDyFm0CY7hteH2uhdhMJ5ebbOnnx+5JT4067fm0lGoETGRWJP/X
SZ9pX/u/r+sv+HEkFfeTQVFWpBLq1sBWn9DKQJdKC1YVs3WJHpy30QH36je+
ZYGBhSXwPKjLQ54lDawuenI64hoXTq2Bgy1IoNE3LwFA7S8yCrPzhkMF5KAY
cTaL8+oZSiVanVCd0B40aRMT+zPTQcGMSoAFRernYSTM4Swu8Ty4KVGcCPxY
KTFtkLDb7peV29NOD3m6UYcmVRVo11nu7XvByf3Ng2bAWOfgmnroXWTgQ2kw
ItJ0kLbvb9hPpnHA18kH1UO3H511TLAk1CGZQVvzWswUZN6YLcLyIJv0PznS
K8aPFjPJNdlL/232cKU9cd8r/XX1doztvtPpREPYOMbdW+beOdqZ7W1EeI7l
20wrIYrD5Sui3MDo1SLJkfZdEZXQKhvZJcAzITJl1w7ux0S6ZtGYu+fJlOPO
qVwWXAQYA9oFI7LhNQTAKTkVZ6qT9rJbPbOyEqTeU60Pfpy4pQsEsMC7TdVq
IDZ5Jp6O+jzw2mRAid2u1NFEmZ8m351dZPVAM+lgsKqpPwnC7tV1YiuNQtyt
mxT5wvTXcRgGbqetcFQjvjzOuZ+/GaZCtygOxWIAUbjYs5h0VbO5FMOssyok
51X17JP/cTpFxFA3FoQJSS740X9pU6DbBKmG2M1bSSsvuUhz1OoyeKw+iQj9
B8VjOVkR4qxFg5NPGHHBOJzqw3O4jskdoPUI3ffn8j6EgUFZpayKYyoFpzr4
Vgnscn59/rfTP7e8+M60728UL4i/CeY4bVDTNT2BwcsaZbBnn1CK0bYfG9+i
lgjbrW8w03s2A36GHtUliwGNM/O2rV97GPoejvVj9LhF+RyBDinbTo9XcblJ
RohZO6OnGcvSzxX0jUeBX0HaEzzKfz8wdjNKENhJJ6UDweONTHDa4OuxaBTG
9ckCmjczbVk/NC1ekApz3x1otps7uzLP/rWPLJ32ZZy9c2xjYw74f4aV7Ts9
05FOrUTviwiOrvtAvIspTQf5D/2LVLW1JXXiWwo8sdREuD9MniON3gQKksF3
swOS2H1hwPTb1QT6QxUkx3S25OX0dwKZtsphO8B4udbRhY63CFepHWIwNWa+
xfN9kHesxC0USRFtoC76PvtQn0CjI3QFm7QkBLB9YfyN9NSgXelJ0TKDpr7D
qXofgDKfy7pGtuVa2JJ6sNaaFfcLHKWJ5nOSnfy9LXe5MBuLJGTMInMGJAyr
uK1xZNM6g5yaTAy5GFVCdgRiOUBl8I6H7zvBWj0MkArpvu9hj8reENEqP56V
bmYA7vRKe7EYMVqxMClUWzedrzaddf3tBXbOqQ9Nq3nk/+hS4tecUObB2z1e
LrrEy2BHb1fkL0BtYUHZskNHWSwUFvG9WERALMZBmOiU5Jy1Nw/5ikaqoNQo
YH5UllVW2f7G9WFpC+qyd2bA0bMK/T9dtxb1NfpKDdHAwCFHK2mmEgfGm3mE
mOn4M9ntF1IS7KdILrJZSs9Mw4r5L60CbEd2YLwfJFXEtSQfDlBL9LrfJ42r
cOsr0Yb0bNXcIdziGf465NIgI7SSsf0EmN79Na19T9SwoAfhSOyS0WIe/JLj
RZYe45WZAz1kdprJE58LOZuObe3Kq9YMlgD47DSYiVRzOy6je1wO/wkuAxLp
o9NeJai0Na+GBob2fzFNUzdlmg5QD3l9RqdoTHOxTmVGROhVujwRZuG3gIkH
+tV/Rfd03FrUAD+jJZvD/MELC9tV/BKETnaf2NZ7Ndi/sHGjovKIavkTquBr
sIZpzDFeCUsVZOOVWRMK+2Ah4Apu6oC7EQ8r/0XcCd8T9hjfwU1E9Vcky5md
vSncKONbLXL0OgVVGsIF0TyVZ1G5n8AAkCkxXHs1MRDgufy/r7yBNZsPNAZM
olEJ6+dwVua4XKS1gg4ouVxnJszl55A9ogSpz5yolAaniJEltKBhgJPQLiX1
JmMnN6H00wXJpMVzvHel3IdRmJ9jvHvsBMYlSXeKpLz+gIxD5BRxCWlH05Rl
wlMfO0sqGnzuEkrUa8+UaHZSEpW6ORTscu7OTs1WJn0gCywMKr9cWzVY/RKO
s7qVRqLmGDtXPyU8byVu4HmsuUTfH/NOcWYifpjIA/oGzlIDVx9tHrr/BVjR
yllaGDEB2X/L06O1CZnDhc/bQa5FumYPBdtEidN0+xEOyfjoHqblAaGHuqaE
zvaRz4y4WQH7K4iYKtsgLWrpTIqzsa4yrheN+FXvD73wMy9XjlwT7Q+0zr+z
nTqla9RHi8ywILPtMt7HI8LtyI8oCJyqMa9OvmZ42r0EJb/oXeLNkIsMdgcT
9rbvwUXKcRtAIoFrm2UiYjFDVYvo1tokl+j2Jn1MS1zsSkszzFsSXTHgQwe2
SrBhMrImU/yYKRTKjGsvnbht9oWFyH5722fmHF1HYYaIxhEjwYq55Sauexg2
l0XX53WiqK8Fem57Mi4gT9BpZhI8rjAzbUDj786g+klTxbY3o4QCgJZr/+pH
/YWveM/SmdBASzvjwAr003VZN6k4FwhIAhEQPx4Zkage+2YpPdZxEPJ4w9Wl
rSczNCqb7cxiaRxqpLbwFjnMVztzcMkxqF9SFCzvgKIWH92u5fLSyghe7PEj
mjRk2FJxJBJ6vTemO05UhsDHV5Mli/Yco0tycUxPGcIMYZW5MKD9xaLjmVH9
Mhk7PGmfc6WJWxQqzXA2pLFWjcU7l5BjUxMQTw8PkXPxp4ORV5pCrMj0EoGH
krNEVNCvYoVhm+whfzDZVB/YhZmPUUSQP+E4SLuzho5jHzEeCnJgXWeqyEFD
zq4xZWJhM5eRTCGidbsjVcgLNzfwDiomt+l2vZQ5DxllRLpg2Cocwwhs6xvb
doFRUkD2ppKb56nlCkmrZ1123iJ96+nN/LM6DJdqByqWk5Q19Donn8KSm5mq
Za/yK3ACWWo7j9aqVRdcxUqDOB/Ji3NNkQCY3ztn7jwvh1Rc/8xwjHv1Yr8l
R0urEMg/4ja/6EEmYUxq5sGB3NtvvC8Pbeb00jhBvzTRJpVJ33V2n3xYA5K5
DDHvlbReQUHD3LyhXgmSexwtv/s9jtVXaRSg01wBz75eNTd/6Jdl8b46Ix/j
DxnmMgSbTosiFG8yPVY9mLm0WRm0PX87iLeoaT0+2DbVZD74++7zb1W3rHPT
uaEEWZjlyQm93cJzlPKQNS11T59rImgz8VgW7FzNDgs1+7WpeeFl5S69F2x/
m1v+UjzUtLQxtP94ygSv2EcCq3yndBq1Ca+ErsHdpVpaii2ALVHeBf5H5nJU
Gq4PODl1PdINH4OaLvmCSnLiMWXuaXUrN8TvrwAcQh1tGnqSjKJf9BH5+Rte
+CKhuSEOmDkR1ZwQgLLaDDtS+ziJ/NrH6xeGmdWSISF5DyUOhhJptMosUE6G
OA5zRIq7IPnlxNKy0dZha0nL+ZG/gUALtEcGRyPdjbW4g3zohsUIH5/RvDEt
8LJK/i2jhCZKBvyuLfxSi6guP40DEChUr/5tbNaRtbAFt0UJT3tOmRuYNaM6
xWMZLGGHYCmunqIBB5VpcEfliU8lRFMJQjfMbN3aTGpbq2gDrzW2kb739WFN
XkXPjQZyu9Lx6jF67uJ+0tar9mNalaIb6dFJ8rRgyOm+a6N+T0J76hDUpZ9f
oK20Txt22L8UUTh8x4SFgulMDV0roMPYT4666JKDDuHF/j01SLxAIWzBbcTh
8KYwPjxYrBWwVxCEULEoR+NGXFeXy3xGbNPVhEjjg9SNot4AXH8buU6QfDkF
F7NHHDIIKKG7/dqWxap80rbfbysBD8Vp9rJnAn+scSzmSygfQPj6UK7B3jPq
N7c6e8rhzokKYllgl7yxOCES56PfC71JvPqqNFyzvtxq1tjLaYXEj0l3EFnf
38oU4n2RB7vOJOWkR2ovzj0Vx+rG1KkgF6wHoSMf+fu0TEbQL0cjZdq7j5Tx
h7YDTeAfvNPyIFCRM6cKtSYtCyeRmh5n9vEXi6FLXunC8va6oJ+igI+GLQX4
i0/a3MFUYhw9NKautGiQd4xWz7yBC424mJQtb51675xkuPiUE6FliKEeo1nT
DN/6a+Gblwr3QDQ7QX0gB3dJFkcMOyIDoAYGLt1/+Tutr8GP54bPX+YmGRMJ
+KtyP9uHGyTLWGj8RyVsESlwtvaDQCJR1ivAhE4FdcMJq38BNVE/6l0/nfn1
5kqTOSb1H/d8bxK+FuqBetSpkKwAdDJ6g2ZZoR+ECzCKi3MCmIrXBAIOgIdu
TXhF3/xy1Qt4S+Fh+eex7DjiZWqla8tCZm+vpLW6XPzBAHYnH57eijLGW3SL
gnumoBCJVDQ28mP4r7mojqT+WkK6vc2Wlxleb/qR5CnnMXfzZ92zR+MtbM0s
kAHPgQ2UR3PJzg/H0RFyiYxbx2CaX6DyIdcmfwmtXxd9EcJ2YjpiQEjBIQbz
1iy1qqo2XmLMUEWOd7OEgFrrQvuWvTVuqjUCPL0Tr8Q9ovUKzO6VfOqgtXCT
VF7opDmFNVLl9wQgiH4ryGK7MHXoSd4zEZvkmQ2MoAgl8mvgsyCR0emy+HNM
3y1qbNLWuSLDzLchgBHCLxNImGb5u8wSCzILtCsM9Zo9OCWep044htgIrvzM
2voTT+eZ9qGe6AMkUSyzoHmBLUDMlwQ7nkGJbm0KR1fq4Dorj3tIwhUacxJX
2m7oTsSwPOR0HcVr7GtgtKXApmiUOha8OONf5660xO8faopaKVhBnkvFcJpl
BBWCPsGeCd9c1LaQaC8uceouQueU0ext7TjVs3wqPOpmuxlEredCFrnSxvGy
Y7y9GP17EUnewa4y7VcCEnhJy5PXta4gYGPS8VTjecNrdxO61riGkV7ZMDBT
3qbeHu16AsG/AgR17F1XAd9WgcS1ueYLsXYnGX+WP5Zgk25vMPWZdxUIRZXi
OVM/Pw5FKTgpKWbTLI+TbRI1p0gah70422CoUes0QTmVPhub+jLkMHQYXiF7
gqgrqRGK8o90Nqo/CkcX0mNk6+mJ8cI/9ANNqXbf+HwqlFaGMfoxmAja/c5S
5rS5Pk0K4Uc6X0edlgzymO2ELkKbGOsRn4CYNRIeRTHayFUhPzAXADhsUynP
fWEos0qNEr67yAtoJ4cQjX79w06Wqpv6/TNQsv9dw5EJCBFhpURJRTAb7LL1
gTeAX/PLWO9hM4tNyQRDVDOGVffTLUuoDh2WFljC1XG/LCiMUvtvclNSmY6H
hWDS4LUaCBONGEoEQDbI7YhG4d2Ppl26jltcbJGeUIOwwsaJgx6hOG3fgEY7
1Nxfs5zTiIS+JF8GpU1MzBKghrrmWIAnPwzVXq1Uh+D/VwcXAKvhA4reGQxp
95cWHW4w+JnefJAmmQxp0z1Nd8FsQjBdajJxp/7+xYJSLYSvBVyiIoxO+Yv7
KV5NCr2vBbM490o1IMpdAbCQXCaNF8XXQI/24KbsBTUelyZdLfDbgoAES4Z2
VpfoyYr2wtMHjDmndkxwyiS+KgS+QKIGcyO3B9TbY3UpyRcM89btRGn6+oRm
nVfwZ4tTqPDFgrtcJZFtT5LcFq0f9l4laEEEoWSMuP38QF6lh9h2VdDDdPaL
DOBmv0q7s70gJJfrmLibyjJVATJkXCXAE0IdbhVbIz2iu/Qbrz2oDTixeJl2
3TUdLyEXBOhubZDH9Z0h9jk4CGzdmNjx5I2VpQQiN61E+SlUTuPOQI1b5QvH
98J95zCzZ7To9hrU9f4qCmcz1HA9N1gA/LwfDcMyfUN5ZmDeBK5ZaOS71DhN
AdoyZQPHCy82gyDBp8QVTPax3+LtP8ORVvWz7VKiZVGFEbodQ8qTmiDMKGw2
0NTAF99Lbfv1MfR25d9KWkh3LOZHE7y9X0Gc0ILXcWSuhm0kWTcDPH3BekbR
I9itAbM/t6J5FHLeRQwPOkffwhA2By8YGsJ5SDDRdqnIcnHKjpcAzHefOwX2
AkImKWGVQjkE5WFUhp81oHPqZkD3mnx0csKg/Jc7tofEtvfh6mDOLebjrDjk
Z/J1dc3SzmkuGXj+wzD3uqExaOMA83dSjk3Nfrp7mvxxuiK7qAy9i/Wc1WEs
nVdi9YnW3nqmvDp0mEaHHs/Yjxso4RlHDzTmtV2ifFK6dkAJUHLEwrMZrd/N
h1s0SiV6jon1cvwnM8MEPJDC7JtVhhvTmSlQFP9SvGQ4amKBZX+4hREukCZg
XrOCv12Ci/yISAMXIDJja8+a0+r5nICBcq9g3fGmMHobeQFvg+ze5kUXh7t/
LGuT7r0Uk/c0knPI8IcEn5Sak/l2UKVO8JTXlGKO8Ahgbeu/h5TiXvO8pN+n
nx7lb3MpMiocNnfgXwLepUK2v6HxkA3LO+MOyIXJi0cX9ff2o6jc6wi+KmS7
C5J4JQ83YjGdavOFfYInQuNx6MoVcgpSrzL2Sewt67jbMrh9F2RydsWhgItq
LVe6HimWEK2A76ItmskqgsQ9uq+9WUOwTubXxXQKpTjm7cWBLDY8lvUuopYa
emck41Q/vCKRiynWkup5tZPB9FjLvQlFCjs8DNDOm8xc9XlvibX7Rvm3rpQb
nHjR4gC9YXF+6QQIzq8BuXFUSDqVV9OIL7aX8TfY/vBQNPZrum9HoOBe6Afi
KxO0Me4cpkZ/Rog2JjI2EEMFC4U9M5aOiSF765g4nL/U5P/TRcaHeIADWdj8
Ij4yCcpFvkUvP1Ng31+YRPZwSQnRKwC1MhSrvior+S7oiA4CUNXgPCYJ1HyC
3g0Fl0l1jt4/obhpc9TZc+q8YshD33YIGy8xJpKzhGoMCTTw1M/SOGjT6/N1
LSSS3o7o8l7rErszsqFl4lQh53+YU1TY1lU4co83PoAQzMEsIYPWJHb7Q6om
C17zs790uB5nPccuGauRQ1FeUDRLNNBfChNFkShWO8lFxeh9ViDsagIYGsQa
GB732vmmQXqzow7y1Q0MygawMSs+ISUy+zo0vOWtpeOZX0dqr0I1bLiZsbCs
TOh+W4H4cjo5vmzUvqW26EC8a2E8XM4rtagy9nL2EWx7run3LvjnMWmq8Bu1
qd9p+HlqKVe8kpsw1vhcYAG3m+Q1wLPa+9YOBNoSB+znCpooetRG5MSn8t3a
DcNKoLJgRDTWC6TBfujflQpjDH+pkvYsFOUUGYJ0YI5bka8Em4zQPTb10ppB
zdssFuM45lYwEapV4LgdarTNWoDTywi9kv2mAp/RzkdrHmqn8ofSTULb7Jf4
n7plMZjQenbExTTr7IjSAC6OPfgr5YUa4ct5vNRz65T2Q/i62bvWbWhXnBWc
5oTQUKe5qe8RzlKOWCq76KGUZRS4+aj5TWbQ58XMbLKY9q0SOsx2tzvQpW6K
T0w/EWdxYovvPKoe6sNBZO1DwSOtI/JgsqJ9WFcHDv5YCx/Z1Qz7hUQbXO2Z
yzZDRdOwsFakh1zP5ZRWAeJ6rX+VQuDGiA/G/XveBdsSMOMPfUZHmfDDquLp
pmV05LEdGazTgHqWytDQ11qztjRoH7+TXUPnB+H4jfUeJM5ZYfZuV+8pgvAW
XWOLu57rKedwDD00t1G7MJOlgLtZ4DsWTbvHD2zDne8rX1jvJAC2IxtGhZiU
IgEd6zi/vzb9z6+zwXO1Mxn6ilvqpRoKvQu2MDh38p5nRj8BJouMWisyHrQA
xs9E62q81B1ghkZ5lwb0T2d8PYoi/2q+3SRu7be9oPbJ+bG9J/p5XXfe0fU3
fLwexHo46/JOkrPMmaRGVsOWNn7+ICYm15uehrGYbXGMPI0YgOhD6CR84T7r
zragTURMed/B3bu4db8f2cyhKfgODI5XDU2i1XasnSiLbP+Xn9RkeCP+Ygcf
qsAoEXzROXRUKM8tZOCpozYsFl7RHWyWVYEXUPCvCQc36+17mLnqnLzRYzAC
H33YxipSbIvmQfZLC0cmLnF8RscAqI8dPWK5maWSHjJCgQiRr73DVqDFmqdl
+ow+1coCEK7rjNOYhkzn7cgJUgdNRx7srS2EolzCPBMt0sHp7poFqVgDZc4J
yaAFPKJTK97dfmL41L/wzsn3jgLvhiTrVPedb+krOVDd98L8CNM0yHo5h345
Q8XWhnrVZFWePERQ08qrB2JfAOLhrFBynReEr2OJ/ZsBieRogXNlYZE+ILpP
xp+JwV2pZj4Ytawx8xgWQ07/T7l1D5ZeuWDdNXgA3Z7c9PhimC8P/n0moRxl
C7yb8yOTatpun+5fazYajFVSByViFoWX7mgDIxJQLiXxeJDSSfNYtG8jGCvW
X39BmPggDpwzpwRL4gv9hYsaj3ubcyr5HLZ5ebMvb10HFxxKXcVGFirb8J/k
PNSciY19M7QszVrZIfIJKIAS7mrHbV1cugsOohm44UecyBS/JMYM/zDCH0FN
4fTpnZhfJ9JjREN99U/epssVhkNSIbOWh5l3H9EtD9WBVmZkemNu0ESccZJh
XoBw6fkPd7F4cLOk6gWT6G2owT35b2AnqUFAYNftr7RugGa7PjRr4TwWG7iM
IOWj3OuMUtgY8xneE+JUdDNILDD2THU3EUJM/N7HWT6tau/0Ep5pLmrwMwmY
l7X3MGTob75qOcACPQiopcsh93Aoqt506oUBPiBY8ShGCblGjRUDPVLXReft
2h3+sdpoNjsG4MJ2DtLE8XlY3pXFIsUTmwibfba7rI+4oWXZIUHX0wxqYQQe
ZPYt2PMVIEqJ6UtVO5JTHCPt66d68fzVfgimHrKhQ3ZS1xp1t6AQK2BT4NWk
vqCbX4p/MDwheVvaZU81tGwSO7dsDzJDTJRM1UMtkF+9R0gOmOSQBxruEdpC
1vPP377vuCyqcUzoUrAng2WTLrFo3vKLihSSR44xoa2V+/EkJoDSdKRcybYK
zTIkEMrfV9HeZXhjWRiOZiv3UTqBNWzIl0Du1w8E48M3AhxtPp7+E185PUod
+HGMn2sXmdcG8BrRMh+AiYyidN8QTU7wHm1ze3IqDTpYj1JNEj4HvpNr+Gco
kFsTszUDK1sFnR88NV2KPHHVtt1LiBQreGtGCo75s34kJbP5W+fWcV7LFkcm
Cpxn0JjeWo+zoG8bJ0p/ezzMDX41Moce/rF2Ib/C4IiVtnsbBLdmKngeno7w
2u9NGxeFKlJ9mW/+8bFVUAQwhJ4A8WYHozhVXkQ4fyczH5FiCxNL6mftoQyE
xA4BXYkNL54f4VVjqCeyhubCc1KJheTGdILsn0khA67+qJFY/DS2G4X94HIC
JlWZhk9ZCtZcJf+al+otfLb0JRY6+i9GzER/dWleJrmu1My40SuEsEKp8vq1
pecVBu+g8DWAN5alrtmdKaT75DmprRycZqLKx+6Sl9mssaR5Qr8TOi+/8B56
AmYTYzmgrkFhRlXDyMGiuQa7Q/NJL775An5hfppWZbrncKaSOc6sS/5vmnrG
UMvmgD8KCDFXY5PI369f4r+oBB+VrqOy9ze8bZVpM7lOF/6zOIxY7S34V7L7
9CfqsZPx2N65FSvLESxuboQsqH3t+icZvTqU7drIEqO+xoVP3qiylDywszdZ
zFuk6YFAQuJTCeXW296GYruBmCw/YYjqz6kQaaK08snaMJDElVXkdQH5lBBS
DAO4KW1qqjbHDEvoA7KTBYGtHjSFJEYXWmxLr8au67HTywSMUoLHlJDErWFF
z/e0pwfY0xnT3OMJTgEoMqQc+qjC0TB/ug0Yz4+FvuJ3AttJ3TJSFLWoOJrR
dNO2s2Ce68DOfkiZt3z0xIRFcrh9bXWjIq4eny+Dy7blk7FbjJZRSVqIefnC
jnc76FtcjHJkDYD0iNPjWEOx/nZljS5IVQj19Vx7qW2ibSqGoeBRGa7ZgHAo
3nDh2Hi9mSsedj9apX+aznbJUz8s5/hWx0TNtOLOAVaYRKUXRR6qBQ6Z5Cez
/EeENXa7luYiqySAxVv72AH2vSIvDbx+5YuYg+ilwolNUxQVDDF1/VntGRNs
MQSow9fQfa+dfHqfw1hCNxKDG+YKYq9aa4e1xUd4NUpF0/Cct1yvu+iTuTkX
hFY6wy5pABhQDa6aF8GpQsRvzW23ai+7/7BGeEbnB+OzXCcId9ImTHyRAX0B
+NHHI0owQereDpZe8JaUsbRUbHJpbjSxIUk6ql1PrWkTFKL7+nUs6QkvpPPR
wXWiV00dI+YA5cWMQrnWRyc0KDMnhU8rR5AF/KpD6+pHFiHHZdYpztBYFeqi
QC+x+x8zclv1KlESD9D9Dy43KDfTGcd2pZ5FfxAIgkWwnjCrLCtmDUed2OD8
MK5GkoQjJH5CUo7t515FNCMqh5I4CwCzWRqp3Yff6Ee5Gf6/CAFrnAzWsf7V
kgGJ3AlXTPTTRxwVlj9c7D4ohUxjFSt7A9uGelTlDj3E6sL2xH7+O7+5EdIR
OGZn9bHEV+KADb169/x2hB+QwoswYXbLHJl+gvcMLViNFrWFd0BHIa5lahlp
Zeo7YpKS85HKeBHp20ThX6gmIqjyFD9yi7P+Cf1luNONGe226IGUMKO2otCz
jw/uSOK1Na60YU3Q40gEOTBXmqRD1V6hSc2/C5c/fhsCkT3Hn2QIufSYNsen
jH+AZ0i8lLwNGoDEN+3VaiKPAEKpQndZfqvLWJmO7nZbMcKCoWRa/C7xdFA1
IBvFtXcqWhR1m2wy4V0I4KnQas8sn0SpbiGwfbFwXjtxV7TeTE+J9p9/mxt9
dZMXSsksH/tvtgm+lZktOe75i5OPDM7AgjghXl/6F/z5MJyIwo7zMcLqdMEc
+tHGNpEjECKOnsR1FIImK4ut3fIjYbc8/3fPqgLfZx33Q2EnlqZU8rDsmDw5
hggIRK2Dypr2dCPcRIRbq9HoGtsUiSNTkabYktiXM081GNdGfCcO15oFIB+/
j8pSzPwjTDaIsGntPrzqq+MU5fu0muYijXq+jon2MaZ8Yb1dICwggZVM1vTb
9YiHX1oy9zYnNkf0Qhq2pQiVGr7hsyUbkN900sdyDakkg4wPDdjkOWQxrLEL
0THDc+9wrnhbjaluadp4Np7eTYqqTw6Vxgu2XsmPwGasJXC+LsWsS7Pxu5ng
iWynrb0a9usiZBHjHPtCdgZR4LKR2qUF2AlRqcZLD1nCLm0q76qrSitnsuKQ
6XoZf7GHkiXEl7i6M/eqGBTnzQAH1VLHE47lwONguk5b3aPw6cloCYDvzN2T
n5bO9xZPg0MEVx2qeWXBw0HSR7XYtwX7PhxWMlTG1ZbXzlMQKuTxO2jnBazE
zRe+wiNSVs8LoX/3QlwbHPakMWJnvGomuTyvJ1pxq9uHSerxFiZuZFyt5Jc4
5DkLFVomuROoP1XSZn3N5jMHDZcLWtuwXojSF1Jfdfv0tEmE4aqiEjabYl0o
9axP2vr55vAC/2FyEcZE6uTpzQORpxGu90UBi0KIAWX01YMAUTafOD7rP4Qz
d559nr+AU3bxRDLPLp6j2ILyuK/FA4/4nvNMqEpQwfWa4l8qZ55fLQs747sW
0ROK4nuziVqd1JKr+kyAqjuIBv2F8X1RvFhrcoae16qq2ehWX/ao0tucbiDT
DwS0RHHKmhANwo92lU+CkKfMqIkxZTRgKVUb/CHYlQ8Lr8s4Pziyy2gL1xqx
eRV1Su7NsMM0u9qznVp48RymYw0PQ0X6TZ5xK55Z+hc0sZd+8YrDo+LBpHNe
ked6Jwy4Mupr0ffC0zI9nRIid2KT3CICWiGpeilCD/fVDfmk0pWdLOPfSNPl
ziq6buvrtdbTIuXm8LCxMcZybusPwasWdOjkHXF2iDyID49QpeBy+ZJvWOrM
V3rEWneVbNFSgtqQLKTg6i14GZLn9QQSvenIeqFm3C7aNu0S+XhcxwmJfLav
u7GR/Ds5nZwN1SXfxqYw/3pwXDE1OP9D2E2fUjoT2/4WvrmfS0OVHF5COCxv
nOWiF0EBMSrrzHaZnp7/ORg2rPI0btFMxs88PwAl1K+0Vs/NJrdYxZXnW3X9
be+BhcULWzkJ2e4F2Nae7n+1duulOctwKUXyrvWk8VQvhaCj26Bs16aU9H1W
JRmk3mifdZkGdXKoiIqWvWj9dMf+2rkjfLkqSz/PVUtb5xm5E3o/aR2BaMqj
MOTaZ6roLaZI+AFu7p5nFrITrgBdsWAs06iz16MujEMhGmzt8DSdlI4GCaNJ
lRnOhs/mYG03pJufp/Ne0O/8VuSYIfFAGP6x6OG7Md+jD0GJPcpofdI8PF6I
2mT5gQjs+QzH5uSZJA+mPWtuLcgNVm7o+ZAlCI03LK1GXt54/ZFDpTp+O8hv
NYwm5cGVJuhsLL3yE7AMxjH7QoU7IH2S/Ltsa1Hikw+4yDQ9TQZXKCErGyMZ
WjYVhiUkfbi00Cr8cWFotsEbGbxPUinYizRyu4tN4Pucvr6tPdr+wfn7WVm8
Z7tGTkbWbeq41PyMUO9pzIvdziJIONBx+XFD47A76lznH6uc80XEyZf5Vbk/
FCclvj244/S6JnTnfxzLWukRteXby/293poY/DFDYSB9IOPGiyUdClCvTy2h
ln9c2b4Uy6H8UyqLb41c0OTMWJhIJXIYVhTJnv4IGGHfWxokYuW1SHg3tgjW
3VHVnb6Gt9+8AF25lZ1y07AQFJoDaJ84uQjTTSHQ0pNzutYI0L4bVVjoy7Jm
igO9a5LWHdooSdo8Y1C5NLGT24gmpkBl5Qwwx0N38PTntuDPI7dIBF9ougBl
lzvg/ugl1FgaU4PO+9ZIdjAo4VLiKeXBlWJugCIzmnPII6hXomX1IDt1wMKh
rYY/Dy6M/BzP703QiPg6RzfKa65WoHXqJkEon8p5Hi9stu/f7BUv0a6wKJgJ
Z1FEHikLizsCPzmp/uG6+wt+nxukZnaiL4UOWzvYaZHYOtIh3vFbhraObjjp
IIaDDFmjGDzPyzKI8z5bHk+qn9mZSDDIIwzqs+NLvruZnkDLhd+hBiIrrIM/
K/KG3ar1TXpBgH0HB3NFjvC9KDEZnDdLNJlFMI1l3lKQv0HzDX8pqOK0Cj6Y
gDVfJmdibiuSENlguyuPCtgKM+8xUmTujWzVOS8VT2c2iSOMjICpcVPQ2/SN
gAfOM5/c7hVf4pGZjNw0gpRuFFUlpabFpDb0YxU6jVi5/Z/Smfwf3O6bM07R
XJ05RrLswjonb+o58LRbB15gQVzuTS81nSq449/xdIIYtVS2p71+kMtw8gZV
nDZ8uN5ICIOUfLsQTm2MprT/yNU4l8LEY7GVxkwr5WCI39tPr6WADINb4TTr
cVgMZDhOE9BW2afTOd0jpyP/+cJZjfUTTmohFXAk1N+4QHdplR85J5udjRSq
8DSkUgWAOLhdpqMkGQOGk3UfGTK22iG6iBryMnssYTvMI1xYgnY1ZQFWX0dL
bnWHvABCazpD35CM7L0qyrsO/udKSEkx1re8YzaaBjnhMr4USLbpPbmwvL69
4kz49pqpsh7pmdfDsb9PpbzPxUC8Y2z4w847K7EQrFsfr1GPC2NhIyM0aXxM
8Tuxk/fwzvu6TCNewF5K1vkGlxU9UQgrMTF7UfvgApnVqPzNF3x71D03GfoT
+UG4YAeuVPyZlqRlC8OjOgXYAprSLVihSue2sXS4k5VnylloGEu66vLrUJ0H
kMrlKNdJ6I80y3a1MJ5qbt1fd1AKH99V68h/UfEv9S4LKGiVSrdfsSaGUsuo
RNF7FnKZWIl0Yop+2/tw9CV4i/qa/xy/4YVYPsEkZ6LqHVEuWJBfCfFhkxoU
KgdkOkO/vGdg1Noa1blU0VHg/YzH1P9tC5PziVffMGdsjUdKEy46xHBZKzQt
3T0xlhvH6gq2xlgPkaKQd4jiluDmFuYs9HFse86H1OVjRd4SMbK2h/6ffknQ
j9A3j0kk+/T8KAll8gy4uB336uIXPwphF6b/Dj1y+hv+XDrdrMeo22/cIiOs
r4ocu1ce1sG6uaaRKiozPv0rwEixTQmDLNj9pJQIyOO7bB6qeBmvXJBMcG9T
MgSZB8gR1d3WsIIUCoXl+Rbn3TOiL9QJ1jXrsEqkF2gR5NZbRYQJGqmAhdXt
VWA9KFC4ARAM1Wq1vzyKnpUXrR9kFwyv66Zcr7kgSO/o/gfkNDt2zK1T2gyE
UsZzsMginVMgsnYQSsYOwpsk1X5gOPlnEHWNbNyrLQgS6hNttoqF7h9KCuRY
hQwdw6cgm8Bj4vLO+dbCSyypVeiizZoI5lYmYPj1q1SZ2g67vm6OIkWdDESu
rhp+sfrxaEnd3SBu9FVIA3eV9I6u8rf2teY2wPaTLxIXcv1mmfauuPLCOtF6
x2tLn8DrFhOrWqaJ4/aQi915Yu+AAOyfPHGVnirw80FoVw/t7jm7Ui/Ni6bU
8sj6qtJEZHOMa1tUZk/qBeJacIFazF0cGIm5EcrV9BskKCKzMoFSaifPuVme
JrfA1ZUHGU5z+aR4s5p6rOnaagi1WXL50nEOqUSK4BMvhNTd6Ms7RsKRw8Ka
a2ny4BepRdby6H29xV0gSxOoK2qw6JHG/2PBRxE+LKpHY3iMbU3IoWbbt7Xm
E0S6817tvCH6vFkHOWbqkdr73NTu9BrezrarIO8mVVWf62NkkGraWCYF78Ps
Q7NhRVRnrEMZ2FeLNDssfbePltyPfC31qvpaw2+JvGi3mWUVvlR3ZOyt1Bpp
uyntSlPRwi96e143SKLYDaB/NEJS/Bmpm69q4inLHHEaiZavSaaEAIl0ZF7x
1bsT0aTTu9z0DGkAPOjQdxnBFFIgoWjWjOAXdtvSQvOupA5sFkvCp85k+GAl
vVAL0O5demsDYeOw4PD9NwfuN6HCrD4BPcufW2pjmPVgke+Mq+oTrwnezc21
VmG+C2HmR4p7X/D0LIMefoXdCzbE11m/B32fB6eixaMZfnbfz/8ytuqX0OF+
fJyXe7Ev4y0tlwOADbkFzSwbLZGg66HpfT1WMztthqlEObRuz0kGvssT0J8v
3/yWXA6lJcLr31C0qQimpnbXVbhfho/N0g37oPSGEyY0dyAYxQ/M0PLI0zYm
rlcNWwX9b5hpTB9ivcfnGp2lFa81fvkAg2ck62ecCTt0z0tu8doNLgw2o/cf
QSg77cZHRxNEN9JNbOyUQGGOHJtNXau+87bVDt4MwPXdIYn+QK6RKDm89sMP
H+I8U3n2BGG7es2RkFKgo9B8y6uYpzAhgETCoXjPkVBsa4kqNVPogqJScm7d
/VSAzX/ECbJkSoS9M40MkhYhXARW4VnIjGDkvsNi/7pl8OmYJr+CYwPXCPxi
tJnf+HONw0Sq8F+QVF0kS54EAuOWsdcwRfzOaSpICyhVFWroO1eIA73YvzbB
MvU9HNwBEiMoz7pY7RA6FC4r+sewAY/6bV0ORxq++UBp6vJVIp1SBz9mgkGa
3CL4wBYiuMbksaZtH0luh+w4ymbO33EsmApT2W5aC3hFy00ZZKf6SQe9P3o3
ptG4fiVMGj5TtTAxQfU6cdp2lcaIsd5U77gLzdoDamvNK3TwnGnIgcCfyg7a
Ex2zAUlp9+L5pVwIgvVNZSTO8NNOo1HH6VrEMwA7alfIVujnuW9waGf+UD3+
7Df3yPfetWPi//Mm9auNsRsHZpTLrUj1FsW3V4i/ZAPO9UxMpORk9ujQRUN9
eBkUqTiRPYbV7oS3jkNWfevW/QTmW0zgdZMULK8tFWr6DHYemn0ZH6sgLHHO
L6QTSwZ90aOZHyQOKXkU0um+EXYlm+0yDyL+tpHTfzgsZlrk+5NeI0TwUKu/
LJ7ZAhmcRLh2fvv1P1ejkiubugwZg0Qa2XnI0CipV5bQapHC8DRDiVRqMLe7
eZUtMHNet41YsrE6PP5UxJtRpebO9+Uv5ruMDYLctHoFR9Ak3z1EAHB6Ac9S
sFQMaohLonS6UGPn7nlBLTupbhr56bAg/QRD52hvNZV5jATQ2umn0S4C8KXk
lAoZa/yOEpWnrMm7wYTr44juBPMdX46tPVEDIo8h/la+AGG6srhnaKt3GYNa
z0FhiL4AjPpZyDV8pdxYGJJWHGDhY38WNhF+wB8YliqrWf7bv9FopOCmEzXK
6c/sjGM2luZE+aOdwOxG40yYF/sCxSB5YdMXYQ+4YvPM0R6Vq2DZuXINzvyA
wOxirqWXbt3zN39zDCP6vKBYFmdJuF5PejXHdzBJcfhQLcihn3IwOnUJ94FX
5AUu0rTZCAK+ccBLGqlInpQ2iLJRrm+wGDiKFrh1OiBuBFx3Jf9E8QKZFT/8
Y9+ac4h4ix5vGH4kIJom84zKNrEAvHiPkRyQSvosxSuGTUhN8NA3vFKnRB4u
ID5Lkj6qqH6vhiXjTSvX+HCuLgpYkfSJZf+OSk4lM0f6x+NVozJbNQY/Ows4
Eyy8zBpqzaKJ8+GPpal7FIIR3ySoKLZC52LWZq/whjR8ln9FEAQb1/L2qSCr
Oqwxz7LCxuVJyUOA0SVvmmEhyqXN+lkgPzE4i0SJ7UKWcf2nKmDytd6rodcN
8N0QObtPiWhfIUO+CvwhsOSNT0Eu4KSfzdImYdwsUUFu4B2yOWZYECheEu4M
CcVhYlqYpRDrWW8/ivLj9aqFAkW23vH2yuWpZusnjuoxqpFlfXaBpLnHHARj
G/5Hifue9aXZqOb0FulCXdQiLRdwcIrwG7s4Hw7TjFr5JJQBo6ssTXtcEIb2
y+EE5ooQikMdwTNnQMphy6aSonpTPw2vURRkFupwZ6Wo4NSofaw7O+aZAtGi
Ay2ccOJocAvlf+xnCFcUOIXcAMTPEg3ZECvX3Uc2prH8O1hAwDAUsuRqF85u
d3cD/KdY74aPxFUszD8zYHzNHEQCh1vF6mHlxJvP7+ooYRlBhSc7JLlA+s8w
sBXOeRpV78CcCZOhi6OBcbEZoc3JybMeitdtFUwDEBBzvE+Iw5gnCTHVKVr0
8lz13MQON/it+vG2xBFG5jDq2AtYcieVXqr16Ec2B8g1LWV1xGtE7ejRLyKw
TPWO0Hg3Ng1/EvRv9B/pEr12dhmgWoM/nkAf+NgS/ZMNaajKnPXPHRG7d3qT
QWL32YOTjYTwJsFX1hKm6zhu4LlWZKaqhsZLXgXAfJum3psKtcopoVv0vt9X
8GNg856KVVDvpYK0N+s4rZIrg1Agp3XkjcWJw2RQEAjN5rBMGJHDb+U7lxqm
JlyAGQbAfV3kkC+p4zCue75105av1ZHiU9JI3Z/B/Nsfv/cR89zxpMIc4K7m
JZXP72fqZLKHeSwK1AjABnqB2j0Ulw5bl5OH/xdBKTE6i+1kxYBIhZkVtFkj
xS0Qa1zPShVZU/4aUH7pdDRN1cwUN1/CH/bFnapY//yMYsVG4eSMFfhcVLan
YT0kFhVy6KFcg6gcTQ0NmV9w9I6YfQ0mwgAzi96lVr7Pdp7VbzLTOcmBOSgg
k1/NBXvYUt/J1R6W17lmfIvfFq4ntiqcb6pxOPRP1t2f9uFNZxLMNBnQ9fGV
UBELMjlL/nBGOuIl7yh+tGtmsTc5X0LyY8gDJp5FXttx8u05QIrl3lFiL7Dh
EZNqJDoEfBmL6XOfcMNhWKeFeaXiteA4cc1PjFJLlfHA1Wn7wgaPt4Gznk1m
loxeWaZ6lRzlsxiISQEFNDECber8Xmdoj/9DTnIeZaK0wRmNn6TlIBV/atrc
DUCM0S9EvFB3Tlo7ENsgJkEdC57iMIWPv9Scp+7aTybURTWHTCFSzvory8W+
gQcOwiRMIhrvm+I7oxdYjae06lPFmL/HZJB89QSa/i02+JygGrpH+OwqD3Zb
CLTNDs9n2b0tatL/ne2utO5nunK3dGIH6KJmoF5YhbDngyXZqk7JhCHGI0Cn
EwLGDIr2LRCUhyMrlC0lWcecBRu4/KLmn9+m0R2CwTHHwZdTc7L0/J99X0uI
v0gT+mTdryDDFpGXUnUZqB4wmedMHx5iMCt1zphcND2+0SM3rxBJK99HPx0K
QHkpFUkqW0+SZrwmdKAgjiAUvwdyZq3qOSc27NF6j8Y36oR7T1QTygtS3TQ5
48MygIlpufslf3uuKtCfhhVTetyN4Cg9ony65OVB72TqJreigEF3Tdj9tTwi
1Ptmr8qzX/Fjnl52Vgh/pHeE2HSUe8ZW+lmaLk8Lm5m0KvfCF/aIsZ0XJEZK
1e1BnjzyCUcP0OuRjDAx4XCspQTA3mTTS/C+AVbr2ayPm9mcFYqOdywFpzWm
K0v2fs0PmTpnt1ffmOeawhRPrPBh9t5R3fjZFcKResYGCo+LZZxjLishtzXn
0aJI0aYRvaDyVCRVZNJ6nNB+yCRgE8QCJDK7JYzgkm6EXnyjJ1nHrIPFNHVy
PHDVthkVaocnj0daMyrB5X0xHRlzjfdBaMu9703wPEgACr4ePFsPIgLbRugq
8MKG12au1q9sUyvMNAlTCy9iXeglx3HnaVQZF57z/KPWya+YYaQVF29vzl97
K0uQm5dcVnWbdfpexExOSbLH3KCefqaN+MPKKc+RMWkDlgsK+gH5mvdgSlY8
SfR1HXBZYpu4YiHOr/TpX4vULTw3NZtqkC9yk8co5wBQHaPxD+ebLW9nGODB
iQbu1d1tc9TMGxZoZSY68NwvB44DLy8LUbdzpApNjjCeGcVpA7V1TGKAe+A/
MotpphLni2sAGFLurRb0OANNQNWUvRuJCpXgqfscfnKNyM+ifiUeGWPTiKA7
tzPle1y2fFRaR9Ag4qgfMnSABd334ULRHAktu3zMWwaJR/PlCZO66JKFnjKT
8LMCAlu7nrTLxDNMgQzMYmiUhcj051gl0+lRlLfAD/IOyfG6TA2fyjOhjkwK
8mCZfpH0YmlYd5Dn+BXZdOeauPslsAcAOGJMxCgeetHj5jdPL1uTyf+hXabA
FTHTFQBkeQPMAkjstS0Ivy3W2klqrJ5X4cexWo4g1pF9+9d/SFicTTg2BHaJ
t/N76q5raI45Y4gEYyeFMNIFlajHBNhhP4+BgILFe67LF+YQbD+5z24LugC7
PoHN+JN/aX+5KC6v8upolgpgUH49DVmjVyK0FoB/VBkrJJ4UZHCHvZn++Ytu
/kGRldRU4pkx0AMpqnJoKs4M3wu0D+4AqZWn+eexzAP/ejB04Byl9LY0IR+j
thIgOHrVZWxRa+oxuer4u+/CnFxqutN8BHQH4coXqlqjszE/3ObTtDQia71h
/GhKkJMiS7DYOMDg1gZsDAQpfO0U1Xyx6rfXJ/zFKaJ4ILlMZU2otBy/pmgd
38C8yLT8XQPvgK6pSKf2AZFp1w0yTze6bFQ4H0po1FjfXsI2J2Fv8Am0M5fG
3vSLyWSISM5XRWY7Rv3LhsY5Xx3061UwgC8QRtM6AH+IytyBXdY9+i0iT7O/
SSF1FrMMpnXuJz/GCvAm5KkHKuZbt1LUOcmAm7Ol06VXn5aGU1bX787M5+j0
WdaIZIL34wAXHmpj0p0sj550S572fT/GtnB4Oqyvo3Njy61zafRknuijlapi
FzSIJ8Jppuchgg08oFkByGfgSkuOwrZWcFZoaRpCOwPTfyapZpyYstTCdMJv
uBpwkVtUKtvNAVWPN2U7P9WjmILIU0vCLvEq7JPhUmsTTocKJAdk+a8rlkPs
Nv2TZOgZ7dyHDZTtPKLY9f2asMwY/lyHnlN7wreeVbiLFSLuFYeYDcuFNhkN
qrZ20fAvD+7iK1DoaWg9OI9vzML7bq2KNiyWfszVBcJvcyBEHHK0LK5fQ14x
b8ZjimWjXUzs3esN3KldBAD4Hc19C0U1g5eJyDhyD4JM2uvKYOJDmUy2EBfB
J4XsVxKj87ObPzBopxRaUBOtcRVda3MBe75SySkLlkae3OPd0vYscSf33yj+
fkq/X0EXQIzwYsBulvWoNNFih15oPqRlQDJ+muYgx+ZuvC03WCWlOeueB0oA
RT1vGdFUOrt+NaPzu1PIhMlWEoBmdjV9odvNEDQuVRZaxraiNLMdIk+UzuAT
0acxAhFwTDeSN7a/NtUfPRYWAILTuWrfF9bLiosmloijYEf12uEJwFNAHZKZ
vKw0idnaaIJg1pjj/DcS5kmTbMYN3SOANpvKHUolI5bMABFY8iMiXgzmhNxd
zqd/L6hwXVvUJ/JywKRjxEUq7jytMFQVU4u4Q1iuZifhwXMjo55VE7/AsCGr
jvRie3uNIWMS/dxKkXP7+c83uO1cdH0F7Hx6hUEXeyhKCYDRyIV7ec26MuE9
PK32Bnk5yJbv0I6B+vkbk7q+TGZb/Id+ON3g0CT9c8XLG8Cd+x+nuu1SbDFw
tiLbKBuN2giWkepBqEacwHkJr7tKu9W+XKYBLmxcaRU5RTtoYmCNcPzk2q9J
vJiSlgzsopU0U+f6ET5XHphPCu1bPf0M5jyzkkjOmDbmiX6ZuYYD5Zjc1Otu
sBQYPlC7Get2oCv9W8KRpLfO8SK0qnJ6ymH9xgJtvek3LCHrmjC2VY/UPz7+
Ql/RFFA4yrEj5b7/fxKplvStsban8AhqjjfK42zawNgQTEXW1iEmj9ebk8bO
nFNSczodGMbWbIfM3LAfzI8yVwu5TZDGjXS5zDUUBUs+3LLIWfW1coAacY3t
VjmLVsmRWZnucrKyD9ztZuV3XgIyB7uMj2xGE68Etbxe+gR9e5V2/g5kYezT
ec4D2RyX9ISwC1RH+wm5JUc2PMKYXwuCir1rNIJ2qvAdxUYwqVvpx1QSU43V
nqKmC5niC8UFSHoRXkElRvo+aHbhs702KMXpcXYWSgAObFD301HmTHqPUU0j
0nRxHe6xo6VCk1inPphGDN2WTxPWLrG8DnuDYieWcKNjrBgaP3m/Av6+yPGQ
y4xVgevO2khkXM20eVwcGowvvqwYgCgKwBJAm7GFVDobxM/nYOlsyDuNoi23
vH28wQg2xI1+Jq80dbTdsEElOBblSIA24EEl0py8MUq7ACgUess7FihSlpQm
IgbT8H5+o2XbCUgo0GKBocs7sCBfL+a+ymmEIP93DfW73toDdgpQuTsMWgLg
SOgOv8LifFX2idfNhJOQiKnpM+8AA1SVm95JI0wCHnA8JSwWRl57MGpjx41H
g+c9B+ffsE31jaqSpSiED7zZPx9/PuSo1RPsrNcjKQi90a0gXfQGgnORfqGH
rxiqc1g8rKbuPx/VGuWmenJGba8+lBOiKP/HvYf4piu+y0AIyP0u3/YKoPqH
Ki+07g0HdBiinC7kjjdeRdHzef/+n5YiK0BSfCN6PBQ0WnK1aUIciFInIAkX
doTdfwGCWW+ZBht1tIznEphzq6Ub7/QnkIFG6rWsa7NR0N0Bbqst7IyPu80L
TWnPFjzuX7rKTNd1+iYj0fOINXhHBYDWHvc7dKKBeFEmObJueQkVyTXfAIRV
RyVqEFmD5Q3gwcQjWlaIE3ajU8Nrg8NpNEm+fYvwAAoz43i5lifayRwUlufG
SlyLnAZ8RUhrxA6+y+ufzhVgUgF+Ny4T2cxmc0GtEukeEdVmzqsf1um3lvUT
iXF1qwnqk/McK1k2SaRYgbs0a2pEc+Vsia2/mhLzN1rtPCSKn66+Uue/2ImS
VMiciXbB8D4AYK2bc5pYX4iH2SOacBM3Eoi2lAsR60IxOy8HjYg9Z4ZesaeK
NPP8DDZCJIvWuVE1Wmt6nF27nHzZcveWNpUjmeJkm0Zv1EkWMvaiDMW5xGi1
5jl3V4Rdq6ZCF2rAlTbMYYAsLqG5N5BHOhln9VzE3h400uQrieOUoQCkpLjB
mJWJU8tyQNhAy5XCparPPEfRwouJWtRW84fe46UWxnZlIS0aWTG96aK88FoS
jooX7mitdJeKjG1XehUNrnVfyx6AlPRc6QiYeVaXIT9SH4y7fm9G3Lo9bVJK
hwOFkF/atsjGdE1HvcdrIdRSx+QmGLyQUq6m2YeMGHFLk+BI/1Xqc7+0sRDq
y4RPH/hsXN/9cPuJeKwBywNVDrRbnkqOvTfuj/rfGDHoNb5JiTGeiKFCjsoN
rYzub/aIHx9HTKEfEHUqgqlxtLJkDlB/czUEntU/QsD6Vetx+Q614sXy076E
1CdPbrdQinlTcjtA7GF7X548k3L3RUbnFnMmZc8CAmjbh5ySC/9BnxiN4OM4
GdO7jPejstcQVBe19BgOaIJDNURVgfAzxr7YFflFyj1hj1ULb9BMPJ02sTqb
DmZvrltTwSY5uwqxIGuZ2O4T9qCtArn0PX+lKdfGBOleIe98i/QfCjI2iBB+
iDG8ycBD/vTCuELylJ3XEcPi3vKEsjmDetQR1Uur/tMA6X8yXRmAwK3wSBGD
QP4eMpTiu6hc+nV2u1vxUs/WauYFitGo6LFsU6dI7dAMx29KjermjkNDpTYh
vNnw/EKyXnzy0qH/oFUu98Ztbw+easluXlabnO5B4HfNlIdc+QbzeKKWM/mx
zI81vXch9xTL88H+XvhBZSzkEJhjunQWJY4uxU8buLwCfC9kFKfPPytIC4YB
2lOuhOemy/GJRQhtxLo4wef+8vEBD4NrILEh1ad+OcWuBZHKpM+ezdgEApUj
u04z51+5YNvBTZyWVsntrpFfa+bIpHIK2pcRHIXhGR2CvlflXYlqJQ/yjmIx
JrQBEz0ALEcTUkoF/DcSDQEtZXn1HZAUhqDu7LlN1TpJHJHzCktjRivIMsit
tf5x2iWLq2qz5U6jATn1fJ/eXoJbkb5rkJSbtwFXcUu3yRn5anfnXJXxKO7b
Ebi75vHBAc6WKmzyxxHMlcqkeVgqct6d561gOPKyMF4qR8j48aP/XKQ28IB0
w4EQ8Eiu3kHXVjVoebkFVSndSrWVduXckXXsYK+OORy1EYoSrLx7Bhoa/H9Y
VPxfgUG1XJNrhD+yMVhbm73yc8NikIH2tMtSwQmwgdXhTC26Ww/u/+yAfwHy
8iHAIQJ66cMDWNTzHvAYcMGoJVDC3YXMkeuvFT1kf3MfxwfZ8dJFDhi9krTs
xUgPuUfFCu3iG9lv0Frryjtfv3oBt+/Oqoz8S9o3iAFUst3g+x8gC09Uzt7s
iNfymufYhdeM5n0E1h4QS+CSm1g4YwcdDVhTahVrJ3L0kqA6aafDVABAX3AA
YQzzSKM0LchVtZryY0XXIoEGth1qIyZplLkdyL9gnRpDK5BQmRBG9F8PwSFn
ShrX+ZHx8dHQo7AfTkxzWAol2mg7HiQqLIFBG8cAkohoMdphelTIUBobpPXh
dyKeaxEEuWSXYnfqEJkr3FP3unh47/JisW9hM5da0AH8h97QBJQqxx92Pha2
a+4k2gg49XPJQTiL1Xf/F21uhr7cwLuAk7yXa8BJ7bLMQUvmtQ6g93bDvS39
GhAsgtFNuloCpgTcfJbSR0aiJYglEBTnI24ucZwvU31NIPxkkLEzs/3UoSt3
EMc5/H5pVuNHGYwGNxeMweqE0+Cd0Q02zwGdzlavx6aXVMI0hoggiFCoOYXf
GLlz1e3XMU+QbElkaexEd/7M+vxwZ1XA0AWQH5mCX209TVJue50ageCSaraT
CyX+ZyZo6pjDmINRLnfrDg3qFcpTR9zq9Xh5wIHRlt/UONMMcSmPUeGdWWtH
yPan+Q8d5Uk6B8qAX4WNMYn/gaFQYquPgTbOwOJ9ehYjZHpfb0n+pki5oMFl
r8aBvtAbTo94pm1CxRnWakZILpuqxcLrMZ5tc7zoYXlZCq0krpIjI9UG9wvE
gcQYk+p2ml07UAKHgxK6w+Zxr0Clk2JIQpO01RJMcUy8ECRIjQC3nw5X94sd
IfmhN7whxwj27+xHc3/76vabRx06QSEmuu+zpUs2YT4uLNvvHEZc9EmIbSc1
+t1Gd+vgFsmpy+wQ/JUBkw/DLhX2XcotC3WYWEE8WQ/au6LLmxHtwXtNihlI
vpYzbQT7GVRZhyrh3n/Z28xxSfA9ffUVUwXuDi+XhOSSkoJ9R7EV9kaFj1+3
/iZjyR5QvlnhmLrcMfS8Sv6xtp51OXsh4VdgZvxA2yHxXACqNzrQa2a8qG7v
jszNSBUlEngdVR1NZdVGJeU98CdNGNvsDvUIUzMS7fFJcRxKXFMhpfnKsMd+
8Rh1RXYZrs/JQclWbMTGUTlbaXoRZxA9KDnN24B4AYS844Czvp0yxX9zNHVE
YJBIGrhMKVcePRW7e3AXhndz8SbIGPW07W1btfPiHhmag9OpgJmA/DAQPwHV
m8RzY6ckHpNaLeVbI23iWFhzNFmXYp1nefmpqbR7ClMECsA+sMwFVwsema/C
J8oEENAnPW2TeJTgRzuZJstWu8lPSPP/jYZ6wptC+E+K4MHt7KlzK4VPm4C/
3QxA0t7ohL9YjjFEF8J3kmQpYIfs3Q0auF7oMNfQ3g7BjoGdFrFzf/yty3KW
wGfv1uJaSO4N67qj2f2iY3CXLjBkvO6vYCpb74P5NXmRXJa77cxHWt4wSL43
pGFxrmym/dduDYNIBasWg2jGYaVkaQ7m2juxYurwz2HucGfhP6Db80/GPmJ7
7td1Ps1nWuP4YhV2pnB7T3PIKaUeANpExN0nWqGchPBm7cjZz05e0h92n72B
QUDPg+eKY6H0uXRfdtYoE5Ek+r1YQfLU3WfKHz4gcxXOIsSmqliW3G1YBvmg
Ly8bDStLuCNiWiGVIunZCpTzTBrIPfv75P1IC+z/AxQ/4t2UL4GhBJ1Bzrhj
GK5r1IWNjAoaJP5f+XfXbo8Eu57hgdVKPpma+XecM+gSPVdpm4znC7f1hlFW
Ok14JX1eB/VFeEuhSdya6E39utdduNRsjIxxMnJ4r61TBYVJdEImo0y503oF
TwBFUuXVizcDMTeHQy5/uoxIGeqY5DQ95lannMX/wo+3RIjBHUcnid5u2+jz
0SWM5Hg2kDlkNebtbER8agxfkQ/yCXqGVmUcs9vXEwWPFcZl+dLTVkmsQP6y
+1kgWoqywz46AsRYbCf86Mui+idAJatflUaaX3MLjZQW902dvqWGBpV/ZW3Q
UpK8p8cGj0OoIASubmysp21IB/45SByZAxXS38O78GuNdyZl8Awn33Y9e5WZ
8ePCCpGkCIuuk12fm+7aJQtpmyjUsubroRrOpfMGJ2P6wvoC0s4HBbWzQq5v
XA6ewjdalbrLqxUM+aWSupKWWveRCjGggu8v037x9OmKaukTue6bOrqAUT2q
PBr0Xcd1CxRX7+mpC7yGaN0OJVlKfg1rn9luxR5yFbDQo1gXZWkx3KzfysB7
4wJhA6vwGzrKYeQDly3ZnqQ+f+YMclGZqwtlyD8EKCWR/eGdQyvLNWhWkfTi
IH/Jtiv/+2+jgBU+lt5h2BGc9VhdDCSD0PMA5NKiWY26Y8EetNZElBnYi++y
qiYv+oOSWM4RMJAvWCJqmPNhtUDDwH7I0nZteFqLPWFrRY6puxflRPwHvNRM
W2R28XiOOmhUJRkPI2qwMloVwD+2wSKJYU1tDR/uKqNKd3EtOG4VTO2odiED
EBMqAe1HJZVGVaTwrjro3l93O97oJJbRbJPhZmFs7UBGVC+mrja7Jz0vxlEa
TpfRC9UVIDWBq83NgVMupsFqmTvJh2h5nxqFrv1XUXTVczXmY/QX6dKNdcac
PCbUgyw0JCQGuasWjgQWgx9ZFhArrc+Z8nqx/KR/eipKdDdiQqVyCRVx/Fg6
d70ssCCHk9bBavODhOfQyJqDVBd7T41MHSxY2lXmGMRaaXnEeLYtm7SZzKQu
dAXIYLHxcuvd3v+sImKswjdXQaIXo66Z/bykH3iQqkUzfUjZv6ZalJxTyOpP
Xwwv7ouRdJi8jR5J/sfx8Vuasdmlhil7U1g+mO5q0T/YJtvDmSq8ebyFwaO3
RUjWZGCm1FHidKVa6dVtTvVdq4BjTrQ9NYL/b/iUHNcqvP0CqdJqDHOccfjf
x4CHW5uggKVmyOfcHIZbIUCj1Gs/z0u/VdmdJcsgd285muXjDnB4nkvmk7xI
9dCrUsLMbnzUOVieQUcI1wJJlkZ8/SSwfUwoLlC8cRHy5HzmVAwkehLa0uP7
dH1APe0jx4Ub9KNHgPIga2Wp94pDKNhGIPvuMmi+XADDOI+3mA9cC0moDwoD
2tHqdg6KS8eryxmWVUoek+ztBcn/9LsrFgSICSGGbMl4nZIwtMvj9FkcD+Od
oIgxM38RnxPyGdAHgNg4pwEuWBfq8+iyFdh3ITLik0PpFVLfdaXkh/z3EXDt
Q2wKImkZDyzq7yHDi4o3WVteqBLe2MLBLZKmA5lS4NlfmVkynR5FKBGdaPGy
lBVAVYe0yMcKef7UlYfYN6kyQYKRh/saYBCLRcsEfGSu0jkAg+qTW0x6hy4n
iRi4UCBTn+5iVXz1b9QsUilfX07W0qayfceFycjlZQyS2GBNNaXlXs6FwanI
PP4i0HFUpGqtPBmtS2dkAHva64n8mInRcPYnTY+fiKOEosbeWlWFoM7v+n2h
sJ/g2WFbNWMZ4+/wGnM9de+7o9NnRKyQDKMX5zQRMrglPDtM3J2/69NJ5U8X
9U2la6On9yeMw6/cQLg4WZ9o82N2Q78Np4B003rPT+QBwPLH3/HWrPWMDAj0
VTPc5RtE9TONMngdL2JwYiypqVas46zddp24nH7VzQ/PGO1dHLMEjpY1YNJ4
qJaQt8m1x7k0rwrUR4ee5kKc86nbqZI3ma27YgBva8qyDseHLOgFEwnHRUnQ
hxfCre5CwIwc01wqHHi9Ba18vCm6tNielF/ar7CuALIvLP7PfYdCWQYo0WXV
hJbV8jKj5VMsU9iTqiiLzuhaCzOvrGCSTbK30BqjCo1hPiOtQtU08MAPR2Rv
Z7PQyx0lqs1sMcp3BT914fND7xov8q2JmSqIK1L0qcpyg0E/MGQWh31uP34L
K6rswZ502WL8PJc2D6h3+mcSgjikMdD31g0GHs5np10EhBDobM9A+SN5zv4/
zqt8CTHKtpUeRwcwZQADyJSPO6KNEhzha3LJXaZl3830EV5aj7CY3VZo12jU
un0oiyhZbkxDJ2aMQI1FRacebmMtxE1L/LIvchHH60tve+AhC6UBYnOpTU3E
+s4lZDAZz2eiDSOFfSKKrbT6UjAetTOpdmIWKXSajN6UVsiyUfrZHa5Ld6h/
wgDzzTaElpaMbqSqc/kSL5zxBG+8CU04lkJowoWokL16Q0UpYDG0b97nS7vU
PD781OcK8s6N9PS6mvUcRcLI5A5iMBWH6RkqPI1y5NNo8GN35/A3CDg6SJCS
Ch9p37xEQoHV8OPE+fETlY6fe6vjyAD3tzGstlI5eTBwLHu6a9MU88v/PuRT
wT299I22k33257K63NC2iazoXodGKFVG93zP0PMFazusOM0otIvwZyN1Bzy5
1OA0pvu3J5Cl1WUlX6eLOk65zMGKtarRhFtVyIlIxqNUhOyE6jVb+eOiDf/i
9dPelIMaGmbQNXC8MyLrkM+tAop7Iw3FZAVVcHxYDisvKrgBjImmKNSM9ig0
oBfAv7nV0RIR30oeLql2KzLAWOhZUYCnua84Qdr3uwUDtVpk2/gtXW+m4KQC
sJT/yk5L1zVOtyOYNP+AEe2wboums13XJtfA6JmnbQJXcZra9ZVK544FxeNL
Qq+OXJMn2wubnh5RisTcD0MF1UwKAhlTQCubusCjp77mmpVvvgs0RSAgvfG7
F3e0rFH3cUEaJxfXaPwe8Q1IZJgiVZ/TsyfsrDUoCm5uRuHXHYowEPlwb6ts
Snr+Cm/CJPg2PDDsloeKnNJFpH4m3Pgy5lBzJBh7nasHdT6oLkszWmcD0sfp
BKcNC7sXnzggEzT2Ly8SccgE6iK0I0YBgsjkphSshAqWkyFBmSGniGfZDz14
Rt7RpqPB2rwat217B9BCBMFkoKksVu7+H6oL7m/FtBmMyH1rTgZLftxzm9Y+
vea/vyIGPO7PuBE1agN0WkRRXwy0TlHJvTR2zEyh0dL8spXBQ2fFmZWYBjyA
4jMFEtt6LeOHn8cxUbvhoqzXEY7NmcSsxBsFG6KdEzJ42FHbUMPKqDtoNQOO
IORjfO1vRTG3OewqlfztZJz+hLRmi52Vm4yUH/7tB5qtUwu3aUf9ighRLAr/
R6EiMBsTWw+kkr/z1mKCO8RgCcUwcbEqkiwVxMW7lCYM5TuJCQ0bh7xC5uBL
Tb8Pk0UlfC9OnJ4ZL08RyIgUhJOtPwxWTk/JjVlCpC3wRFT27pAUr8ioBi6Z
WK6BDr1iponIIzy80UvKwoHwohEH816UTYJXtDaE42csOewDIiEqo6OHdsLm
elQBk0BeuJMEGFk235uMqroNEmKwXx9lATnX39JkB890Zi+oY6Vphf54jHi1
2xzIwnonBMiHiDG2Euo66sGEM7NY/zkfqdH5ZbNcJIsk0Xsdilb6GlEs4Gyz
qgOZ4yKXgpeWOj8pfLLXDTenJTj0nQHMtLDa2VAaagMlqZ9Bvo7gY00KRklm
RaPKtBV3bKFnjoNbMFEypiAAMETtuE3BRHMxFUwFKm/2D5e9w9sqI7svxnPp
S+0fUCoRVjP1BwOyUVXxwdKe1PbJD2ZuLCqxU6YUZFwt/nJUkGfr4cLhQztX
KNXYGs/P3StfOw2EdHi6dm2p4S8Ce49O6bWb2bg+93WFN8dUdZqnPjtSojin
M7kQ7YyN7SdB0/HJvk7//ccyiQad3guaFni+JiVW4fmy6o7db1f5rYmFRJk+
VKn8+5kOdqi5HsL96E51NZvERrtMii0Dghy/MCjIxJcMtWMh3fSto4yRIp68
ZVKo9p1fj3jPZXCODZhaCPNlyB1V3QRpqo0nOcYLCtex1bNP5w70j8DRIEhK
jHVgbONkzWHk2ldl5+x4c05QwJ0iHg0JK72S5SmLlfFwbu/CPlgqlvBqGuj3
/QMrTCcy+0rwuY6WRWK4NphqnWIKXKcvO/924fymxtUKOJJvC5IqQQnQjTaw
9fHN8CTuDO+UnWwiul7w3ylT6bBxx01eUXfSTmosxutNOYx2rF4g7ogKSm/2
9vC67BNWt0qwS9S00sBdtzwatl8x+isGJCmABO1nmcWC3r2wgQUrzzf8CKfb
Y4ysNYmNkaJsnEUGb05kfDOKZZ/LTmmFsUz1DHlqbIGmo3ifIgy2B//IVlCv
5iKy5e2McINc1AzAOFNsyldqcdflmHLMzzoJx1gZJifapt92CnwsM8MyQcj+
e+bDZwJvfGL1C1jGclJ/gD/DSJJBhhRomtnQ86BerIxNLfhTPHfV4UjqWfq6
VFXEbRLj9ZKckbFmE8Aja50DPe8EPDRxn0k9zpQh6ILsd3lB1ewQf8dNq4R2
S6buqqXSGTwB4+nJSKdVHZfy0ZnA6aZJQvr3VZ2PaX+hYx7sitqJm8LzJlO/
l3Oh0UJxl5LihZaRl3Q/PnPYOM9GNveHhmgevkqPXpHpefYC/fVGJpCH83Ju
p4GmWQbw0ZAFxKENGIKwvR7/36+WuwpY3zwijcEMz5cs0dp68Qy0YWq9JORQ
UknhjWnlQ+U0oSg/Tzql4odROM3FGUi7RR54LWZ7ZZdAJpi8xXmOe3PaSAxP
fm9nwoCQtOjaP3/oV3rbFx9fncyQ4aIb58UMxiPtfoLbJX+V4RtFCV3meYe6
pBlz3OuI1fWwn9ol1+YfUY8D5sXeZzMFsn0cxsNaushQR6Shxhb4coLHZRf6
JMts5xQZypB2pBa55twwGX7Dt4rFda4LlcsdEPCYy4qji0UPrRwQ6f3p19t3
rItCPrm7CxMcbHtNxAd0ZmffdQIueLCLKOf2qRk1/PD4yGgqdNILd3xWWFyy
w+71rh1LSE5Dz2fund8ImaRRGCMnA60nFTeXsLo2qWuyVaLm4LU8DdIMJBh+
TtEK5YxbV1gZt5f2sQDw83gPOpsdeqmtxRXMx+gaPFqGA4TKMrOZKxu64jsB
FH/75eLJl257ZAgR51OsDkQd4+kZWah7MbrP9sTo7Ba+eIWOejGmq0eaqqs5
j3a64xRKzmcTISjzfvk2R1iUsChw/ciIwO8Kb18WEW1ORISDqLDOLaD+US80
GWVyPZQbZ85cO4CvK5wwnQrMhJ16gKKLeU2hZH9AQV41Z7YB2Mm6QgBth1E9
OCmwty3PxkH207EdaQEJmY/iI4jgfBJhL8xDUeDStR0kSVe9QxHWouSSEssI
7nPQ2TuHiciKwEPsQUATUau9MEZFlDWNr2BpQEPK28PprifkMiIMaR8MzKT7
es2fDEHT055jthBitV06hLkzGtlZ9sEEtqsgktCm1tdJ/gV6a+2fiOHmqZqB
L2eqHuJjWy1VmETwJVeA4sAOAUNyWtLrWqmhwTHLflWVYeqO41x8KUqN1pzG
AjJP6t0meON7SIldS5MPwoTZ+ErqSZCsNJw3Vuyrd83l0O3+ie2/NI8NNGrp
0QqPZlnfAYirTpNnm5zw+uyKFcUW4Q9J11ulPRSs2LADulw4babfyW1vLe6R
GmQxDo4v79I306SDWCc3nq3krR29A2HaejVYquGQLIfMCeQOLx7JpgG0Gf7q
N9Es5gMFzRT3eTMjh0EypUPIOU1GTZ8CJIWsoYNy4nGiaz0Z/of9wK7MYtBG
fcxdbsUWklKtYlmWtGmnY+8idyYKH5E2xMB5auV9NNsB7baV9h7bCN6o+4dO
GC9lHtsO4LrgIy4ecdP22FqlbtbGvkHFrx7UHkRrTxHSOdma7Eyh8qAGUCtY
9mbA5hyqKpXwK7OFLizgG7Qbq1WkLCxN8elWiz629hicgWVZiT4eaWB52zel
oZisWwdo3azvWkdzzEU0icMLfy4HzpQBKLlvfdIQxZkmmQ0K5ctrlwTfjfZe
6K5rigoiDEicgwI4PLzyyDwRmIUWnHBpWkIO/HMZyA48s695yNJgr1/GVt7g
J+C8e10i5Q5mIlisCYOqmLg9htGeGfqEaJbSvKlnk6hjP0RH5uqYET+K6onM
Ol0IkJB8o10jyxHq14t/t1kUvhWJsjoko0M/9BUs/SvZ/qjLvLC6V4yWPln5
1GnvfASCIE82d7Uazt1RNNVVfI0JlQwsS5yr6OH3mXHob/DNq5rdAfD0C3XY
NkOxvbzm5iNEdkhTzmvL5Ga6Owug+I5ufhWuBKmek/BNVtNBzH67yujmo9q0
SMJpfCqCpGtg24ggCBrYmxkI7PDueBRk05dcT7zGyWu53Ip/57Q+ek58GKBp
jpSWfHa/TZGxQsx1cyvYA+x0jn13S2WMxYp1gVGCd1Ce6DpvR7iBVmfcZ85O
6Q2RXm3T3g6ysFCZzJJseHEXkxP9w4JKZi1FgZ3BDG+zE74dR7+ZlI4Ro94Q
HkaMxsmzrgh/A1KpIzyjPiY/Jguj+6LG31lmMBS0xlcmc74rnvloblZQ6CNG
D8nIpwxd6jnxURPYkJPErm0FCVFVAwSCISsnEOag7hGfs/W3mrFAV77q4us8
5T99tZO9OeZKWu7HqHISQdNSbyT4P6+a5Kw6/ob3m4coqbwnuXsA2cyKIk3J
63+3Iyuj1GrysqKssQLiKy4jdwX1ivcIy6bll4ICIDiNsEnU3Bbz0wLLN5iw
hZfp+1ip2p5R3My04c1cza4aGhBIlsuuTx4rH6jk2dtDOcxvSfUtP7YX2zPR
5qM+j2shp7VnZnolH2DTIjHAdYmibVyVWAxSV16jXLDDYnUTNuTO/QcrdjTc
SKd2zZEB6DfgUx3W+etAjgDIk34TM0T3M9lTKIoBYDdKtAIwEUHrJmC2fSs1
tS0riEOoZDgC35dWh/UmUxEkWFC9xcsO3grIlKifHCa6K52vE1vamSYgS/3e
hV9rqBo2XV94ilv8bfApVoTt8weETPiLM0tvwu5p8FtMeJMBTVfZitySZYHj
ptgiM4WdOtxnmlJVFQYgKrfqVSfqb4b7Xwzu4CZyXr+REUb+u/j/1lVabKOD
9I8OHqawMVFc7/WdWPPoP8zqayD3ZlZeywQaCd/uewOBqXUXwkW0E5DsxFxS
Q/wSu3ktC5Xrl3sNvIIjrcWyAihgHpyVsDpEzjV0FLgstIPDlvnQjeF7uWbX
Nyq+BlHCFwoYJbIE7870jJTu1fBVIltsbCk4qn6osVUCWcPHcthrJt0EBSNE
r6xhspupNgQgxzIvtVh3yM1S8y8lDjZZZTV7EjjL4OkV0N+xq/K2yuiPH8KZ
IsoOe0lx8iJD9xTR8V3AyxIlMttO5sMz3UKT+CoQ38gBpP1wnS4hi/eG6gAC
1W74EQlYKIqnkqUyiH+pyyRVSuILXrg5ifzq8UGr1axTjNw1+GwFjMEJD19x
jJKaRHr+DnGC8WQ95wEhnV7CuilEju5vzLJxUcs7bHsPI+6TdArwyPLIltnW
Rm8FwdYQ4SkNd6uGBE5Nv4wEZcJnX79mXARSfvYLM4K/1qFLrlo4rcM0Uspy
taWw3d263Y4z0o4OpIWRmsHsUgjSFsSGGYNO4OzwtVwU/FhXH4DVo10qIZbI
7GFy/QjHOBaJUf9fQ1eoA5h1pRrFUIKvlRNOW4ErpeqpS2PBhjPgye7D5o8i
togBPTVdtq/gnTklPITzZ5eSVcyOxHJkHySGfgJ5ef2WoykUDj8Yxm8DFKzb
NNm4IWPs4VK4tUSzEB+/HlDQxLWKR2JTZ5hLWy6jS+FkJYF4R8lIk7ZpXtLi
FVkk/e0TaeJ4UZSVs+seJcxsbIxijRXWVzKf8f1uJBhmSP5VaJ7wiN3P2skd
QyqAHmWGxwd39THlH/z7swf3NM8lxUeYt9+qrWaxO8MFmNs+pOI7rbPPXj+z
ht8wJMc4fqHxwqBWKFBuz/KnxjSW48npUaGrly0wQBddkUXnU8+2OAbAU45X
vh0Dtfv8tF8v6lcdxKN8fcSkwgduJbJz/P7U3eOxGOVQ51hSslXdGj/+Pp3N
9EP7Oz/yMlnN1KKRMRIeiYwhJNmDS8S//4RJnF8OtrVd78pU+4GiramLUTQG
4UizEe0kZRtzDWN99M8azOlgHfyN+6HXetmysIxTa1OWsKCKTlKX1V/8aJwz
AMa6Lzz5mlu8qn0xJkDvQr8YMLUFFfKqJmOEYPLoyOaWKHxvqqecrjahpRRh
U2kRc4RMv/ucDtBXlGpn5FgzDBIQ7GTmYTaXK8FvHKjhgcsrtpn3icqKK7LT
GESveHKDaoayOO2ExXf3pXDw2TY+loIoWhLvJijkwJeWtX8l7eOtZYcT2LP4
wi9Y8gNh/VL5iRWc+4jx3JxfU+ouk0/EGKC6ff58tDVMnRrBbXGe1/8WbwWn
BG06gDjCiZAA1c2SuEHsjzrKK1WklBQIBntPTSEr7pEzEkMaNI1jF467i6w7
ReKtNq9KLcNahZfWqnWgMTf2x4b1iy8HUXBUTnusnCSL8C2uMuRQLmcVEVSi
ELZ1Fiency6cuMfOm8EwSvn4fNyZbx+KdvSfs6WchSTczibwqurqLJSUtu6L
RaHiPmVXqaKjKD5tCKgZaXeXmuW7IQHA10dLlC34xdUSF/slJzwuWN27owju
bR+YNUEKMr5aNx8r6IxXnuLfgqgqlHB92/F0TmyZtW4MPw3DE4COZvI6R4lK
/2iyR6yKy5eOBxYxZsgD1gvCy4uSGZdaNQvqtSmbmUUjxNnJgu28OHBGu1gd
lV3VaYjphVWe31YeWn8AI/VtKneh425f+NIvGB5++/DdYI2JAeIi1dpjp5C6
T64IKec9dyZsyxTuO12l3UDCX9mCk3pIJMx8UoCesMgLJkqRKGTf9koypZsO
8Bla7Pp7lqA+EjL9UkLQ9JikzEte97T27szlA2fzpqqQ+4YfmIHuJb3eVtxD
5+72kbt4OZCLCLJs6v+GL7n3f9jpUXOFR1usoQeJdcXQVzb9X75zEEs/FolA
MzGnhTWnx5jsxvUB0NKWSyFOMSjxoeRQjn55DDgPBqwUAELPxi6s+9jdTINc
R8fGkZQJ5afh5CehEGy3KI/oQtrW40BKpikPjJlhfKX4oATGJNJOUediCn0L
+O1Yoqq/5Mqla/8A/nYszg51spRZpevE4mOqnmFbiiZQt8SoD4YkRLxp1UFb
PG61VV2kHr8cxlf5D5fiMJenMj/+bKZcRZtGacRX9dcAZfuOn9N3QU8dYF6G
1zbZudHrRCkOXzVCjzMdBYoafjNSebBlyOsREWPCKGWb7mWyeFWq0XcuKEPW
KCRCP09qPzvipg/IJ0FLwGEB3qsBp0ML3z+betXQ6XaXky37NKAv96cthz0Y
Kjo6RRiQCkDNSdoUTS/TeJI/h1nDSSAyw1hEPDC4JmpzxN6DkZQOTjXdGEdh
0C6WxrgJw0/JdYlZ2LxQk3HerxppupGQx7FuXfiWO1Gt8oOYEdAgkLp68drD
HNw9VRfSA9lnTYvM0/tjmJurfYGGtWJ28aE3Pw+olPLkonldObsRSzFyiFQG
VpCF1RbQt2VhGP8Q0BYcp/4iPYQ+xNlmCfHeYbX3boZVds4kxlGFhgf15Fy4
zmfivuDSxyOlnjMxuRsLOGZ8+lFCorEWO1WGGoxARLvCr8AEyjw8vK71xHER
lmcYGWSqYQFrIvYdCzvj1t6+z8h//odzFUaoTL7shByRF1NEg/DiDrN0Zaas
jbKWwJ1tkGB+xQuVqOpvOVlOVezB59z41O52CFRxP6k1/pPJ67mNmmCVBSAT
qorV73Fi+Ltn2E4xBO5NV1zs6DrdQPXIFSfQ2HbyUakJO5s8OLO3OgVZXYDj
zyYXeR18+Gvl3AW9fM7pA0Zh16DiVQjppd7TW+LSyUv89J/bXoPJv7zYIjgP
VXpsfuGmP2zRcO+zcJ1GWkMlwZ4vnEyzs5W7luSxdKx5wjYiBwhOTs7GhRZS
tEGYm8CadpCI5jY+6WtyRrf5NOP9cEWi9AlLX+R0GyuYguRyu4EcfsrPvEVA
ShDdnbtCYkRBs+4yie7RzYB3Sl30nwVtH4hqkfpaBHHVCB6pe4ohCqCpPWNN
JYzFMystTna1dUSG8sTj65eCJv9VCeVb/q3QFZw/j0A/8Qfc/b8t4h+153Do
3Q4ZjLOBciNSmsaxV2qtmLH0QItVx7nQhdVbDgnh+bYScObwprcrPK1XlBMi
ooNVBqvuuxNWFfWwv0F/cIFNSp37Tc4pKYXUe6wPoFNUHEL1Y2CI0GNDJnwR
mHW/mywqOjZoZDIZv3MX6xSNRCENYGXQPUZr76cQNBDrwoVwsOs3Gh2ziPdp
f2Miq/Ibslu2q5+5VPYg+K9TTArbZ5wOp62BooZoo8HjQJgxBVcQ44eiCT83
+HoEymDLPwpKvSR6sFO+oiFVQyPVX2UCpigTS9dbx3jL/6ft3ykKpVaOAUGR
lj7t90c76NUCUt1ons1YBFNdnTHKGcINIdolM5BL6D+ozV4i++OYABa+1sAv
+4q1IZ4OkO7TOkfYf4CRJG5uVGOQ3HHe/8Ilym4sxUAlHuphTsxSUOzvORfS
bXSi4xYGAerj/BrwLcQCK1IBBsZV1OZkViXxAFKfPV0WgDEOSNUbit4BDs/b
LenZ8qyXYRACTnk7dMpSib5/jIWXymyVYvB+0oqaj4EP0f9j6+29sccDiKDH
JO8c7uK5WRFL8MeKtjj390heL9vWuebWKSEdCq+6ymfXJ2UQ9S58iClIGmap
Zc4F5n/4iMSZacQrMmddHe+tXQK0RQ01yxek3Y4OD1nNgXztf2VxsjdgMJj0
dBVdT3XylfMslyGOO/VxkhOWCmUOt7C37A2msCDJoEUEP/We0t2kAk7xwMl2
Cu/204qUNsfYnyOd5bo32mf+ZzjhF4ePZJo2MnXYCK0kH0zcOubRRKeopP3/
c0AHnlOIB/o2/8DuZZ2mUm4L/Q3Mrfd/Mm65+Gf9xbTCZYYZ4SiBKTdXr0uJ
Kgjm/FxoEg8dseuMQGEErJD4I1vMWUAZow7C0/eBWuYFvzfDolcDkW5r0vJD
hTG0TGvkSw5zJWg64PtldQpiw1dRYvDlLCQ4EFOtHBOiKY57+W9P9qCg8XKO
AtVV4YN0cEOiskwlNULHfcIWO6GuNnGWUJWicbOpdWM4vRQhlpZWTikvDwH2
nCBJW5kljvDryW+lN+5LYyBlCfH7Ii5iBJ7sMWkb7zK6Shjjhbn/R/s5sa6T
Z8+OmUVRK4yRJ3d+eIWROMDOK+UuM0hoE5Yre2ZN+Hxz5+QamB5gr85R+CS5
4XhCSoVIoKbAgb90fRWd/ndx1zUyVQyp0AJVn37PvPWmBGSioI8exDOTkyeg
/2V+EURlNRTwtlZx0xNqGCiSDJiKT4ndsSn0X3F4b+oF+LtiuTRwj0Ut4kNi
x492oi2ajuOI5CNFybWSEsC0MOgHrw3reGH8UXp2WgDoA0GUfGYy0yDP97AE
a22yo+FzAYUMfJ6odJgKqtQWhdokg8plgtnMDShvfZtjM1k91X7wc/5iGra+
YtSANi/wl49t7YIsU7frm3yAs508y+ydFeYxU3E2jMdJ62tftB+qQtpt3rRB
4J8NE9pu+uSDbjCZ8SwOysnFudTihVsBfxHgoqzxHeWjNryXnlPknHtq6G3C
KsoGkiUGLOMMw5X4SRrvkVYw8sfjXTcHNx1oriPLueww7zoR9uWOvqr6puqt
kBM2QeaL28FJgReN7yPVMqmV9ump71j+a8/zDj1HKgkd7PZS1auZdtj4lxmU
fLNgto6Nm/h8XWK1gb3ACo6h105gsDEp1vbldpe7KckW3UFClhcjSI4ougSD
10I9uWsqkWptu7cuwxaYrthsFJW8CFJN3ImC3VKVhYc3B+Ub4764kIXiSvtF
oxKALnR3RZZnkNKFmKF09ipyX8ir+BuoZWUJj9NgiqO4FCL6PPBBRRZLuKRq
FxcQ8SstCcL/RVALdk4HjofIomFuEVpe7Qb5VL8cD5QLAUHjGC3jmtHH0id9
fesnEgt7IEwpVdWTjgNumf9Nu886E9fOFvMToilq0V+QO94o5T68/A755M7e
G10WXl27vTv1xOS1HaBGKrWvhDjf1q9szGHaSiAVdryn/8OKFUjI35kBH5TU
Mi++K/+x+IVx6Ug1ua/lWVLryM9l56tnvYZoOoFNY7yjCzkd17tupTpitGzm
oUPG2WV7X0f525sW7ff9vVNaP1sC8m0c1AbbfYz8M/0eTyOIh2mTK6tX8zmC
r5dri30m7Uy5YaZI/Vv5T98RPPVBjnm1vgqckUanEzrrZXNyKhGIaU4thlSo
W9cJzlv1PJMYxM5iiEDxEU5U2aTiFdgkbw1CvpwaABYmkqHu42c4sVQ/QZZ3
yzizBgyLZ5RjNIXzM99PhbhHBK3EUAOjERHZayUPV9n+cCAsFevQEm6Y0TfY
zun6TrxqVwV7gic10qSqdkkD76veMYjMCmOH81vws1dtMeG6FAmuhUtFa/0y
s2fFjOpv5aZLaH2zkqutPDdl0TSh9cMAdSzLXUewtKaMV6oZDdNDKRrVirHA
cBjY6Z+UXuxpuGdq/MFPpuCutC+8z/cWoWGXocstIkCZiLhCgUz6mBsZVFML
SGrQfE1hHvCBrnR0VHUyMkF4ru8P10Bx3o5yj+gy2ZRkfa+1rYWVVXir9eXB
YIziII/WazfTlBQNNCpBCRlGzYOO+Gaow0jmJeTBKSsTQAiXeIxyREKQou8s
gFG4PqloP1h+kEBAw0/1Mn9QefXbiW1S2ElTjWDnjDL2xn+iL7a3Au6r0oTl
fR1IqCnDsyh17uUKONvu+agxufZvl4ID26R+8rxlpkKE33f/ygldhSaA9jhk
B5T9EzTEPb2mr9vdzgnBmlzTUCk78MGBRfcUVr5Y3xhbLKqXkjGFMTmtdyuT
f/5ZTzj+skKGH1qhB5fTHJOOOhr4IhQ29Lw7DewzROd4XWVQgYmbKgfEkGEx
VLJgqnMnpRUx/8x0mwKzva+xQA4dUHG78EewSd7oGd/IaXUq71/uRbDD18bf
d/pSchgyVV1519caXrw8spcN177lh+TprJmOWrftb+bwH+v6RxasAXWTUkvr
a3CaJ/Lqd9hbRGdEZyJPQ9QFgybprqLh4rXWqR7rd70maIwOeHHZvNSjUe7p
6BPe05Ycl26ow1R5EYi/j2zEe+3Uj0dvy9jzWIxpSG/WguZgumGyAMsYbPQm
5VtG9MmMrO3KTMuL7OvsZ8oqIaQ+2oueYme+q1WNwUvmdb/K5+TnSxsX7ELL
hZ1wVSVrWCFrmY0JUK+c2tFrYdK0Gc3O7DGYXcLTiwEXs59Z5Qe7ZHCkUQsc
f0HlZqPZLpLm7rTNqPySfPCwS1Dk55/1xUyXOIvOmc6/mQVi2UiGR9egUYws
RYvzwwJ1/4skSrXtGm5sC9vye4Z5KdNpjiPvV/3EbZmlr7ExrZRGHxE2rTqy
/9tJEv4l5/IoclcgrZzXnQ2G+wtn4qkqBiboVvauIRxrb5rRk8tNTVjYim3b
1XTu+had8/xgTGQo65C4kUpnlbGbo3fEvLgrT3CRwREY3G17SjfNizDAcVSK
bFZAx2TROFxira50I7xW7ry2HW9rJRb83+taVPiXhDdHEQQLAYsU2cMqemIn
r0WXIrfwcLLwSmJ9u2XwLly1Mcb8UBAl0RwYcfkTJY5YhDZwhkSlf/62RB3B
dZt/oEYqO/bk390MmhEHxMSyAKXbI8KYnmJIkEgS0w7x7/7q7t/RFPOnilym
A/vtXQnVx0sfB72OpUhC8v2e7wO/uy9OS3ZWBmHeiNyk9eRY1ft9IpGYOy9l
EXOpvXfK22fBXxBMK5Idc/nINitiqvlyXGeMJoaShdkM4wODhkd95xU1ACam
w5hZrnChoPyv71xI7eXooyL5WPY7jBW6oCmZRNiTwXBEduvJtC86pzCpzozQ
RtbXMigFonWRMSzka39Uy/2A5Agsj5Ev42eV68V1tUna9KBcmIrnXKUP2vJW
wIsN3a2pxigaco4jPDAW+zFzNr53U4LPUWfn0e5KU/u4C+HquaJCuX586Bt+
gelA5AmcXHAkmMHNaNYLCtgPY+IWPbK+lf6ckV3qSnwj+sVG4qjOYvPZFzRW
o/lkri9QRQt31WjCnt7PZPi9v7Rra8uEUKLtZrX8H2s0ga30wMBrqel+bZrC
mWxiwPpcd3dhNvyLRLtlampTWtsPOaLoLtPGO/kk5pHsmpWaxuPzM5LVBPQ0
8tvEpsgD+W+9hm+uaNJKw+qT2pvVNDH75Kvurq4k/x72i6RH/y5DgfK/WPNF
DYub6fqnaFpQjFHmJE1OiimfHzLeOp48xx8TN51hQzjt7EkMZ2G42mbL5r3z
wwE3r0cBX510UtxGuPw505wMoCdfm+gnzuFux93tH7I7BYbA7Qj0FtttV87V
2B0U8zOHDx6dxEtWvgnKGRn0PFrBO0pV+V3PYesP7HKImVSULT+Utlvo+Gwa
agIMS8hk+C9rqJqlT45hudbNYNVf7jW1Q8CT3YvxaPKvnszQanH5MbIyKp4Z
A574rvGIKbPJsT4N5JZb1K5HPle342VMCQX39ByyuuG7s3FwTHo8ynL9q2RV
L393CmG5qfBkJaNxVBxUH0/UAcJZQPOPCC/g3vpC4qLtWljZVyRPAhgjZsQU
PQwX/X4AyNXk/VGq6S94aP6ciWXi+berEdNwNLs4A9boxBREfgMDM7ZmLIWg
TjvUxQSpcYvGdQTzKblQ348d/qTc8qSZwkkTOkDwQhrDXS4DoOL3I8BRu6pC
ckqLQ1ObCHIEFqL1UkfXIdGXHGbZ4wtNlwz/abi5hYkfZOKNqk2lRCQV3pSg
sclR3ucnnRiQu7Ammx/MxpXqNmG5Q/HuGiqeaHsbANsk+xVpuW7usmv1VgkM
Nue1r59+pRd1gOOUyCRSIpOlM5tr0+Mp3aA89fjRdhURcTrX7TkC0D0TdUMR
Fa/W3l4CS6C7UeZ0vlKqMmtB3b5bU8jz3vrBk66ub0WUu0k86CSCuh7i4tL3
UqM/o50cH3imrIISToq+9mrDpWqh1qrZ766oScVsZcu5r6SEtXXdwwKRz3DE
o35Nj336G/+Q5Gi2fp16yr6QuMCAf3aNdCP4hxY0IgdbLvP3VheQe/XJKt6M
wnGKNjqsb03E3i+wQ7UNWCRe1rachr7rj/43rx2A/+A6a71KP7YdzoMasdJh
ceFSNwoDLyZqZ+RsNWdAeHeT6iV1/9Q29WlUqHmtLTxmJbUWc9W8NySa1VGL
ubrrjleqjgfSefau/1xlTzi4UEqQ+KNFcBFwCWrofI3pHm2q1tcO7vyEXuKr
qiZHaeVxL+ba4YMvHkPqyJ5RjdgNZnj5F8xzl86VKjIQQleNI7a0xe9k98xi
hK56X49bj6yjJplNUwYGhnz6mdIn9uq0C6Kbsm4PKUc5VEZeWAZrmJohX9Kd
5lcuU84NSrXhb9iu9MkOci38CVoEyNxQchWZscMYrS4SCzadTWrlyJefV80i
Pc7lJu6hmjuJhdlk34GLYUMjU+rkoKb/CR34a3MpKAJcDYilz+vZjz9TvJYs
MahlCuEEoYWwOqeRr1vQ5kGgdoHQokbDAm9sg30qKTwymjrAzy4Dtsae4X43
ne5Wa/bZJZ3PE4VZvmaQRCV7UJmfuhT5OxPlSYuAWymTWB1g16xPwJ380U14
W7cjvox9ZCMmwfRe4ErWykThS/rXOAjAl9oYKPnsMED6zckLiy4xG6JEMLWb
67tCFt20Afudyvtvv0vQO6hTvZb2z9ee/BJR8Ywpx3hiD9ZdTboKid9atvvC
moPS69YaGwImgnSd9rQyHLX8kyzUf0ZWROF1OinIFiJcGxFjda0Hvzcp81Jx
rjaSHXRj8fZZOGYsCT7W+mCvNr6kAdRXC+Q5xtuD1sRZC9Qse5tiRbTq1XWN
lyQnra+KOfvvQWMr6t4HxWEHmPVdEoyWEORzdPbPk0fgTo66K27LPuFO2H8G
R/49akWsej4X8QKcTdpr0chFS27mQH56p0Ubb9kQh75NdSMqiWiaGlAL5HYS
+Vf0ZvsT3AcZvMN62Zl6zfFcf2wQV21t3g3smjqYViVv8dO/wfZJ1d6agPOW
jQsZHxjo7OUR5b73BuFry6c5woZ5IZyuqgOzw7qexlpVFUuxaZ73dmZUOTOd
3tCBVt++l2iRkesV/0KlbY54gGF9QWy42yhAQVhoVwucgB5JCIDm83auugzy
QhCwiCMrcb+Z3gce2W47vp3+JFaYCxiNWvWfEcfu54sAMNGAVoiVX4vQrUaS
3yuwRnaW0GT286PD0vrorF31eotmeJLvwqxI7J74EjR5XWPj50vuunlYKr+V
CKTuO/sIrmMVbDrPSN5mFytG7GXwh6jLJB5zteRLOCI0Q9dxegcxV2vBnKXC
/mIfP2WizRC4CmRyl9LzX3UfTWfVn5770dClHpilSGrOj5vDPm5LhDuwH/ws
ID6ajQv2vIv5MQSEWYxa9iQthsUtkOH/4HmcTnAPdseFMPgrInLIo04uijFu
gCcDoSPlKP+SUThaol9A2z6y7rfwVgSWfAQ6yhbcfq8hyL4dG52sotfpj0jJ
rCXHeuJlCbi7fqJUrmqvpZAScUTiM2tnTo3fswmaggAnGTSUcEtza5n3D4r4
Ps3PlBsXiPFSpQjas6/io7PnThqRWtT4PboCNGleuf/shcFp8D6g2y+gB6fA
Np0FduuEOkCzr4qiZ+HffCenTLtCTXJsRSGmNhKIj56xdKjwhCBp0yU2kme8
uHGNTHQLv/3KqTJqAIOmk41CuMf0wEgViQId3FCT+7xh7BWQagzm7FXCrer+
bo0cco3HsK61lrIst9H3Dsfp5WFqCRZRWllEZdJ9to5pqW3vHecj4F/deNLY
yBVdFS4cx04pTJLR11kcwpmpa1mdMeVj1TOBrL6zZ5bvUJtuYTJyX5CcBfI5
jM4d6AxfZqlur+U8EZjhrSd9oQ0Peb6ncG9m3RDsTYNJe2F1c8qh3cICwW+l
w2Q9iT8+kIj+cGsEGznQ19tL94ZXWoXB5pHDxcpnEbHXDtagix+Q0VtlIsFM
YSg31EMA+XJQ+s872lPjSzDjDpm8e+jmxQkhr0X6NqwL5145x45yM4FLWuTg
zrD8d5LUo38V7IUJxliuhiO8QXjjcJIE4c/nH67XGGjcXWbo8fEEzyB7jdXU
ifuaPTQPyGayQGX2o6rTYHZW2lJL5k4VSCchgAIbEWzbw347Hd/lv4b6azfZ
ZtrFzVawXuA3HhEHV+WDfAl97/SzR1xOQ174vx6h3NmvgcdMQkgqXPa6Ed0+
H4wYbMUb7QqZZitdqqB/TJblYyuuKmLe4u9Ecch9YqLH1HqF5xzhcxZ5kHIz
ElsYeAFuqxKul81l4uPq4cXjNACmekSDg+W1GIM/x30oZ7hi1s/9Bo6AY+FB
vBBxEEGR/fhCR9Ox2fzWDGuwOr0HcHqDVzbYomFiVPu7YijoJshEqYwzNfyF
iuIqCjdcHrhv3kqf7mmcIomCoSkNbee9t4ezIL6JPcn6v3dPMUaW9L7rnfRQ
HkACcxQWOadN+bO4INvTG4XhSaEAiNIBdAy3ZSEg/CUoDBbOT0JTZzEuAIbu
1tftAzk5aEdDgVLv+sA0aC1lmOId1e9m5W5tRMmfg6jtapmiIWV0+5EXKtJz
jKbo8gcm2V4daeg6d58JCE3BxXLeoaBLMl/ExLVp5v/149+Y4AULgpYV4ow6
MVpvomhy+QSxlRTcFtFWzRasySEhBoMTqrhGnxzo2pdj3UNa5uKmC+YfQA6g
xgniJ5Z1TtACOTeZw2hT6dX8kinUIPf1wPMwlR+PTL/QRzrNmk3GbLXHk6/h
ZtZRKPQNyVHz+jvD6M3p8D5O5h26va+HPx9/o5Nkxs9WeRhOup7Z+2P2km5U
YVnvs5BeZzRw+bcimwL7VRNxi4r8vp4Ya9fLk+k2Tq/4CVpoDh9KdUDIUpVj
ijMYyssUQ3FZYGFd4OSNaiOlDQ662rw5Jh2j46U6r2xvPwkpI4XBOMEtv+FT
Uw/2oJDjsPux4JDPP9NoJKGcNl/ryxW+OC1wOmaNEytFlp5UwbP0v5snE1m8
QeBUZsKHcUz03+RRO43StWv/WTdRPKrXx9klCrYZ3lwb4dpAdNvuhpf+a95l
joei1UPVYxHz+fGm/g5VuWKkKIt9PiNF4yChrOQUit4gCMuLX/G+OrGVYT9s
ol3l+lsZLJXnfN1iB7vDHATJtEc2IZhXhg8PwhtfbrqU8EyhxURtLx3hgYvG
c3eVFWNlfLaW8Vt1YKhvUlbm3XN2NRHzqC5zwROR+CnV22sFAax8RbuPG/UQ
r+8QZWSGKEVTcriJX1j8Dn+32fYgcZw4IGmBXDNiBxyJUpVOCM/SLKK6Jajh
aOFBdLREOef4CvcBoqbxOwVtnNiGAY5IzgyOa1tG/7w2+jGLIbZeD3YPe3wC
r4CqHgwdKmCWOOl28dbKMcWwOsvLjv60eLbEiPUaimYDqQQP/HN6auwaB/t9
+inoGfrLaHfOOlhHoEdf32L7kxmiugxljn9YqiNcP+K+QMJCzZGhFX6nh6CU
vjZBSrESkbzdr0yHP3C55IuXodNQnnuUcd5VF1tT+2cD3iEAE1ij9XSAnkQO
UlfDw+8OY63eKKtnsUUJAnd3oPptaa0oS0rVyI2Fhv7L1ta5sYXa0HdHeRG5
sQ2aVQEIAZ+8nBffcclZXV64aglOz22AfRf2PO0f3ca4bT/8V5C9yeM53VWR
x0Q7cWTdnxi5AvAn4s43DEPKPeSvy+2W81nSIKd6n3akNUdqx0Nz3QaNA5ST
HsbLww0rtBH+NeLC0dvcWUCWu7rTlQrvxBiRhOn5xRVcCrt7T3LuT+eiRSUk
g2rCwbbvQj8xStgowkduQgNK1oVBL/b3NB6TgHg7za1TU98hGOL/cq7R7gog
mUhTGEO9geYYuEOdf2bnUtWLcUXc4qZjRHc2Ts4Y/D+6p87As9RxEUBVv4d4
/w0Uz///uXSMBN1OG5FE2VN8RRSFqr9heo86MiTq4addwjfY9n6iBdPNBibC
4vziZg8hCVs2Ja+22PvVliV+VP/DSSJCB6xJodA5yLM3rE72Br5ZwrESQ7h8
XSW1OK5OnuAtXnCJokhWtHE7BT7WRps9Bf9QPebgcJxyv0BpJv//XLtOOrlg
6OLC03aGLsFJdQhGsgBp7Dj4iKQpP9kub5wC3tfpbAVlilIk3wsZhJn442rF
ZCKTkaFZldqdiU/dEtbaP60oJy0xFc7zkB04IrRki4eyiqrbbiYFwcZ7Fjb4
gXg+2JI18/c78ATbk8kaN6bFoNT4490Co1Wz5coyzZD7hCOsqschUeV/bpnv
iIRXQScsbgTAc8Hqdmi/PROi6LQoOj5J99bOfQFTyGLch6aZCXujnlO4MXi5
5bvCJrG5QXclxqX5ctpLfOZprJVzj4cP6gV7iEewIuKZe6rw+mmaIQxGWD2/
zSA/kyYP0NnKyPsDS2ArFgLqNLjOp/WK6HnUsm+s4Nbp6wkxIRHq7vF7hT3V
Oa9tYBg6chLFC/6FxAzQ5zjSlQzDaxe8mN3niNSuev/+F7KZWNRQBcsWmJe3
xaykSMpsP5hx+5s25phr1aY4eMwjDrSnmeFbpQFVqioJ6hZsuj8EKc9m0JU4
dahs3YI1PAnbC3Ywv61scAgm1XtJ0Kh21SF0DOpCnqRFHnEz4JvNTzXnpUB/
RNw2Hdi5kZSueRzFCHJczijydOruoMAkUGig+059qzJ/ZPwjVruIB8YtwVIa
jk8CC/rutjrDK+ZNtESWTY8/ZSDUNLFHPHm68rNlEtYRuZuKkXQUSH1ANjiP
017Q/6CGWD7catLy3EOzKBij7ix5NoXKe63KLz9WEZsbFUCq9Ezfi8qZEoKl
URX1XVs7DHk264FdF+ManDFkayVhjnmgsEihqmYsShLxWWJ0/fvJF8uyjbn9
iXXOO8parMUViaHXla0Xta7zQJBA6iqDyZ802+41+SEAma2zrdB+F3Vf4OWz
m4L1ODn1yeVuEkA+HqA7dMqYUfMFe4rhXDZKsFG2DCpWNtBgubPi8wvaQMA+
oR4rIo+FBOdcogMTOF9Dfctykr5eA7ZR+mI0a/BzZ14DTRP8iS3go1ktOLw9
0CQkMhyJ/ztYXz6jgRjR1a+dFYDLEVuYROZTj+jIy0i8rK4gY0Rdkpp7kjXs
4RgmSLLx0dQZRBHlQx8UQqtVuHwQmFbEiwZA1ilGjBeZoNLuBLtxjXraGuyD
QzLZrG3o9hVwhKvtobz7yWZJYVpAWUmTSPEky0k+MSdvOD0z8ytLAw0ZdMEL
toZqtJ8Eh/naJy/7oDhmWhzgecV51C4YwBHYRBSVjVZec2bRxgYtstgqLDgj
F8STtJq8gdTT9VeU9+ighBX2i2B4gn2YCLfW5D76fvm2kqPSQqJspxxruS13
FomKnMlq5SsJgdTsxVlfeShilQn39+pNHEbm/HOVPHyatlvm4t7UUhqcKnY9
EpvJXSs128qQwOwC2SKcctwXlp2AHnEWjsmGAc7iliNEZhFIiM5BEjY8qCC+
i7YIudyr9am3mYdPKUwkLaCTm399iBfpHfvl9vFA2KRqwZuyRb3VJ1ioqqme
PpZwgd90pKVR5BezarBtzIepXt4zDe3+zxptMfBXilHJN/MaWK4d50hEKztn
QzPq1bm4WNC+9e+zy3RHw8TmvvpmLu/C5xW7pVRdTQP+8tEnuxzh70wkGudw
0A7uHZUwwbG3kmLobx4daUYIP6rqqsiWTcqpKubTKR0mi6/0yXFukG0FgEU4
NoRer8O1Yh4xs7iUTh772MWg5jCl2UIyeLSQ8UGrCh4MqOmlrhSiC3U7l88E
acC1Z16XCA1TvfSid/DftnvEjIdyKqTbrvqG95tJO7OEDh6eabWX93/MMMT5
HB/A/g36/E90/ib9N0UPr0ebTjcjL1HfW8Wh/TWHF3HDZlL5eu8r5IG5Ukjz
Xr2OeKtS2/xBaGLUgW+j8hhLxTXqbOvIQENU0fFwk1+xCTzBDTotk1Q2K1lh
C0PDTVSBHkmqZavZ99GoDnGfgkLMebgbntsRwRkt4WWHEmDfuGyLZoRgVS+p
1oI2G5BDn43ufiWTlWqQsf9z/qEMcbMfYSvX6F/bu5dGXw+RXDjTQQjGCVyg
6h2YvH9VtovxEuDYrZq6cu8//6CcQTnmxapsnfs0xpM8kwUWwZBES6MHX6no
emFDo8MyMgvPdWzdifUKtVp/+cP6OSELGk1i7g+rFoHxl8jZhpRra4pRB5bF
Wi1kEvPcL56fZmAk24nkg2hT4YFQc0scJQTy9UmdtvtcOhr6PbwQYqNJ/rxI
mNgoMwQmzDYllchesq9PugqV86jAnd5QujnEKFJEEGi3Pfa1496gIJ3GApBn
Cm8DvvoeYAnrUio7C9L9eMTeSZIZO6VEP6HTSfxkuiZEkcBb8Li7l368Jja2
BPqlYy/yoc38L3oIp2wIw4XL480Xd730aJEuyIIGNZAKVMebAWlwIE7QNbiZ
UWuNELwP9+oZxd+kiY3r/O0T0geeo1Oy+5uCnsd14AR210MEeCZXzPjhIxUO
w2JtNwuGyczzSBUL/HE61ZIYBsViww0TmwxvTtoAj/5X6lGi2opxd7OauN6m
pcBy+OGLeCIuXPawvsUM0NselJYvDMUGXG4PoLdrLBqzVaZ5V3LO3kNpPF7l
FY++eUlfdoKRpKL7WIwt/FUjTvxl5U+kT8SIuEk6VTRiTSc5ZMIbWHtLOZIt
vrWKUDHSavvzJ0VAVwVzekOFJgPuxH9msswFGqGx0PghY4q/9Ba+UgwMbGbG
cld13UTeaeD50eDqq33XqP7l2Fl48ZnFsVXiUrx96AlrX0beg8Q6yESAgdqg
BvpN1Z9bkWvQkPma1WKtQUT3F7vjs/nGeso+buUhWzWHqVb03K7sZ6FmjBmB
2tQGsA7ZNiuBh8I89UY8rz7mmrXJU6XcYFQWdTT9XWJLCKgmvc9+/sDsWzhM
lbvPCcr0cpzEdTTjH8d0HuoxnrKgriY32mXwp53FG1nPxLC+VYW8wEDGUVKS
sa6sOIlRGoyd9Q4Clxl7+zrQI3v3qOhATTSEFl3MVZ58VSQkjiLujIIIUb3T
nAsYooKdePg1Dr1Av7MQh3OuJQEh45LdPqWieueN7qmMM2kWPaYiBD/ms4//
dN6Oxk2cTgjecFeF5sHZ56tjaikqPtsIhifHjlXSCrjEBj4GfebFx8iRrN2j
EfgxaxQiDPHoh/xtRPZ2B42r6qNiLe8GvKcPF3yfspaLNnmkwiJqzlV25kTl
0o/b9WuXzJYgTjU3hwLWGAQn10Dup5hByEUDOYcIOhp9wsJmCYGXok0oXRsB
BoB51JbZ/xFcnIQj0UB+w+WkOm0G2F05b103v6eKD3bppLPqHTb0A7ZlyLsk
k7063+e1wVrK0tagK/W1j6kvbiYI6TDYtMXOKkKXpyVzbWg784GKY/vhniLW
R/B8jWb8+ZbBuvcyX7YH6vOFOgzFOSD6SLy/IJNwDeN6PtLy4qGbbPgrBT62
AuyttwKvncgBJcb/VtURLGCdZIFVvmp+kBLlCQDRl1+UyReCdo9nZhzOIEsA
hjOcOeCJYUgeRv+MyEBC9u5niDUaDBqN/QXlaeKEdJKFnHQVxFepLH6LqTvS
VYZuP7dmXY5Xk9qIvx9rIAXAYxgPcjN6vDe9CuOc9TRuTCUkhJr6BL2FQGUW
QcrbraU1oU6BS9Fy6B/2eAmAJAGNSp50E5Zm+CaABvXR8bNe/iSU0j5mpOAp
BnEFLkwNmxorLJZZgBw9BBsT9iaUe3cD2tmmguS7Jzpc0eist7/gzrA6AC7p
6ybXTCOLsIY7jwRyRq4O99nQ+8IaHCFKSjCNSj92gZ3T12QNoE9E1SI+9eTG
tMnmkGO/S1dYkEjgP3J24/nznMUHcjzcxR9K2kFxmPtVIxjfJynRgra5eaI2
jNkN/yGSzRzDSbTFgHFxHGEvLAlO5f3+0wYB+ngifQHSi0AJlUX1ERpNau+U
UgF67VpsLPSimpE2tLvUxAq0rNaBiiOujv7sk+aUW57+JK/YUkI/kbKpmpWt
gaDTgUY7xCsrPLnL2DgHrlPOzxGPvOwI6FVMQ7qnZd05idyGybXIscX58H39
Kx5MjB7UwRCbgPF9vFbzSYeiX1gc8oncJigc9Qapn3dxi0KfavhvQdYFM4aH
8xTNRnHuNNpMMJH3rKXKjrZcoNCFRDzPfUHbPBiZn2U/3EfVfPcpZjQGTdsn
SetrVz2TGKxx0wfeXKfUgbyBPWzkz6iKGnpoU1q/cWiuAk61VMpd1np9sDCY
mFf0mpKwXVlS5dcaeZyy80aHz1JP1NBlqeK4KxA8sow6l4SO7OvSyiXOu6LO
GD8XQJkuC0ucWvUGyVABFOr/eW47lUqrImZ0+w5p9YhDGdNB0LbKy4vdPvFa
GTUzPBuAWuB40Y8hSKfD7Nx6CvR3lyAZg0/zBR9TT1e83VP2CFzqz7PnEUxp
A1DoDQ8rwQ9ch2v4YbK4tXMkD/O3c8/xd7CU18eyw1IN8gUeqkFpyaVFA/PL
kU6+SMZlPOC8EHcWUr5YoCpyYANE1Vfrx6ZLyb7Z97i+qnpSh4KeL1HFLsgF
uaONhwNWhwDkdPUnfms8BRqnklDz4zelQIHhQDykO46Qz6zE4VkXmMTqDWPY
f5Zg250nA/9p++Irh3Y1tPSyECfiXkY14oD5eu6+Nz1tGKYFwRc+cqedYt1e
xAsTEJTW5A1gJu8gaQl6Babay/432N5DN8LLUoW2E3UkeerNkZOqO6GzBm5N
Ib5VohmpabipyGy66aHJ4JjAJZt6R8n9k/roOq6bg5Z3l3DfFjZZVtlXEfwp
eerPpTVL+i0Uq+aMvfjayYPoFI5AIoLkY8ZbernVtKl4BcuOP02qG/qAK22G
ZOfZFBFTuY7RXP0gFIKxH5GqaQ24972cy7z4P5o1WJvY/4Qs5zHi7LrslLJn
Zl2HdsW2f+M1wh1UNdIz3xy9XOWnD8NtIUQxSZpEkzhsGg3nvPhvudytq0WC
FYe3gytfKwdNrdbD0vSt02eiZJCPZNvyf+wz3LMCAHL9mVs4cdzFdnVnGkBD
n9EJSbeg/wa7DJj8bUZ0guNGIDkjfsrsgzompfJwdW9AwfgktBHRZFvR+zY8
Tch9mOXGc2oJW8EX5LwZhEIpJ8owroulKJxcdmnGBSxdOx5IDLHSkkL5sen/
UAIEcdkD00BRoDgtBKfxFq2IkI/1mI3nMK6KIVJ8Zh+xGtsaURiQ+t7lr5A6
6VQidjQL+ZUD3NakaxTXu8j1LQXZdw9z7KKW7SocGGlfD/vu5m4giuutv8/L
ctQdgLe2WEwe63+E0HkY7ztIyKr4yvl13gQv+pGu+orB/11xGucEmCDy8Q5K
oXUKX+d4fUpEX9jApHsISawqyZdHHX/Wg5mqwkzVuwbkANKEAkSHPLwfkXMn
Xyk3DSTKnDS9y2WnSUYC6kouuGQGGSmSVi53GktukhRazYkSUKiNuJI7PQRh
y82vg52TbQGZnUztu12KR6Wf6uuIAMHJWGl26MXOTwWADkxLY71mLKD+tdQz
mZbwwXCebZ1ooujMnuQpP8GPB4u23YieJ6YUCMafAJIlebdtv+/+q0cdGYXf
ah+rxSBWf+jUWeX5WWTWVkilFVvnBwAiuEMdMVrJiZ9gdDDSFBigf1HJjJtp
rSm1zseXendX5vxoWHgNXm/BPreOFAOi03ITpba1fSEOTas0AZza5gjSa2Y9
2075HaHKwMIEpDfU1vJ4iYcsP0MKJjdyYzKKTLF30SeVX0Ovs0FWwl5ZwWus
mEeKcnF6OwaiSm+q69UxYt8i6266y+tU60MM57XwfTVxbG+Icr7bX/sP2P3v
2YeEqPVat66wl+9p3e0e/mDnm3xNsjM//KMUaxmvR4J26swryioTF77cY4Zf
tuW4dJfWMPljNUceHdWQ0UjxTVHnlhNuFO5STLWAAVdb8clEbxrlfMJDHDGy
puzgy/RCK6U4cbk4AjhyODdbApPd6qNEtAvG/0NE8WKPvBfKojQdG7clCbti
xebgQ1E7DiQpGPdImTLpgwU9IWBbgFuVYmAXTkB2Q8pXCX1KKp9c9cjZ2t88
p1UQcux+xGvyZxcNmlhBoaa1fVkYI61CemnKI9nWwTbnwQjXrNyjqqSB11K1
/4w37P/Yw+jTeSGD65TfKGbtHm+G79BEBZIW0c8dPnHwTVX23n9CZQO5bJi6
FywZwzrakzfwlaR9+rU+2AoiK2Bm4aTdbTr+quFsvvDlAiMqorMiZ9gHPmzY
m+xecSsYqi2hbh6FtBRqky7FlV5VNuYUYqjhlFySOxDbdzO/5qpmL1N1wd9L
yc5sPiJ6Zfch7LMkBf91OqAgaA+hwfDXaifFRNBkLzsUmOaS3XDSXNaZDUv6
8UwR6Vuvqu9j6bhtg09Yl7vTtPEPQfI6ekspV4SEDfVqVBNvROnsrKtIx50R
sQAUNtR4WPxUDa3ag1p9n/OMo3vBJ2CG62Rve1LjuSuJeDWGAdmptn7RkxWb
OKl63Q6iyUwZzBoLSvnshizjzxfEuEml0/FAod+BCmtSbAj1F2Uhe5jgNwz6
LJdb25OZwfixpyaWUSY2ArVjWPwtGa0U4Y0iFEeGGL4BQt2UJD02Fn1FZ6Bt
jUi4VL3/dJgC4Rh2ipkxXM98WO3UHgbToTYU//4LUlrRV2AIzAdwFzHgmIik
fI/8ZMx9credktRw5lr0J/dSz5eMGBJp5DMuESMsCrDxh6qjWnHyGTN2/dn0
b6p9eV7ppntibHHCzyUWqlhRw/A4z/+kvaf6XhArgZ8oJYe4TodOTi8qYnjf
KhEjJ0mRZ5s/+F1eS+oyXndVD9ntSDiy0iKJ0709kMeJBc5/GQLKAupthoZu
ch8pcET4rXHu8wgD8T2T4Y0aJSET3FXEGAykFtH1+Cy/8mcbqw1anrNQYqFf
+w1Zug9ghNzZrOwr/cC2USSQ/5yh/j/X34kjYisDAMZ+SwCM457rfm5ttk9g
LM3s2wlYQKyJLBIbm0G6iQ1UVbEEKudZkYnd5Umvgc+pibeLcCHKP0TG+V5E
q18Baq5z4+jZ2McK03ePBTr/Oi7owT+Ar8l5sTxCaLk6l7xiRG52ek4oFqrt
nKXs31jN7hKTl/XTvlDkuQU3vjXfYK7z5C++b6shlXf0/hwpIO4GlcSgglVA
uaqU/tRlCVlbcnZIDNHiLEHwwbgGZGnCPRCttOG/iieCTpuqhMKWgHPtToG7
7EgtEpylyf3LoVKfHPtPGAalLwMENO9uMXDNETu9jJs2AJip9C9SDgdAM2Z3
rLDdOJefxOAQH5nr2LeKbkuKN+hvY6iSB4FHVG5CMs7FkZc0+laXzN7gTPzB
SYIu/1BS9Xdwft057jhBB2e6fg5FU8rGafSfWV/LPT7j+VKAIFt1RtxYiaYj
sAPkIJIIoa4n+ZnT/W84bAAl0c9/xHteu/ReWXhdscM1G9n6nWUUV+VL8qc7
6LQwKAWii1qfuKHYRUlPRAi33KXzI0G53qVUdmSw82TWXAL8lGHjlEoGyz1F
wramH5YdFNXK2Ew4OJrbgRz+1vNAswfbJxHxCMohmXb3Tsv+EaPHFqSZ92bT
xQUX2hQfG+8XzCm/3pVfyahEw/BYrTdNzPG+bn0MoghcUzdHe2Lqxbr2OEuo
L8iYufwRFnsz8hx+uDA3dUodbPFF7jlaRzyyD+8U2TlhSaXrbD5f4OyjB0uf
Qycw3voNdlUisBZYk/UvGb8V1fBrfSddyhPEsIC8+UIZ8fLI5h/sfzd1CAF2
qwBqyrL8gt664GUlu0DTl/CO0HJkfnIqYT2D/3PIiYj0WI6IFmoNbQsivi65
0pOsU0CMs64VblIaKNKrBclHarF3Hq4ObkCJjV+t4czloelljh4QCp5oJj3a
HnAD92/taePOLQKUxLes7hlqcMM95i5e2+3WmjlWeyHGNwiPv7H9iE6KpGT5
uBfunRAgbxHunah3KoqkCdWMtJoxkQ8neo1eBdUq4VxNZVUZ6nTf5tclLj3V
vsFhSBxzvKtJoawDExgeSqfQZxPtbJ6X6IpchIW/eIo9/WfOq8/rqLQQYidh
5ESlfcTNj0DYPT2AYXpozF2ziooqnVje5HXQm6wDyWLoTa88cV2X300XcULS
iXqnTIEAwD/snuqcb3i8zPC7JYEZu4iwcTZgcVFaN5vDGNC+6Ya/vJFZLZT1
+gkAfEEX67qg8onvNc95qQZli5THY6g3uu7ZQd8Pv1HJC42iSBMLutKFRuOD
ciTKNK7YQGjBReDtiULw9EzqZiQFNIgUL92ZqHjJYR3nR/Xw599197uosKtQ
kodO5Qq3Tz0C/CyBCz8sxXnofZGqLzB35oKE6B/C5mPJNIyVMqyu9qYLAm95
AIVipweYsWODeIJi8HpHoaHpuUCjlarvCNrLLfpZVAl9EmvyByv+0CNzoQ4z
RzpvzFut0RQx6Ke0UDa+enb1egyCss+pI0ayixjs2i++9XyTrHkNzKe70Maj
/86ba9E/SYrp6Axrts+bL9IPqbHhF5BVYkoIWXDwEnEwDo98lGBMQsbpRwFy
jm6ltu+L2NXBUMqDEwUdxEBIf6R8YkIopAY9pM5tlDTVn7N1Qvpme15ilhlD
QGjHw5dCZKvd9mKlOPzB103luYzk0lXsHS79g1VIZAw7MYt6XS1xQ82B+5s2
0yJ+QUN7k9KmrNIT9n9mqynkbE8VhRHEEhgRiYJWtBjpTpFLTQIeHvQYU375
uet1Ub8X1sKax/4nOnGnVULnYZcodZ3lWi6Y7ABGPuHfKt8AB7Q9O0KyM1QR
VdR+l6ysP3HN9JjE1xbFhjQXBPHRvKhYcmQgx5QBA6FRs9g0mDJwXlD20b70
NSuiUiWKR0rV8ym2RggCGyYXqb6+Cw5bCuE+0V2E1ulLfL/UE5Evjf+Xn9Dw
d04FMCsgJOXtIBLwfZwGlo7unCePyoztaCC3eDYxK1LpJpA/hPa8IYU7msnz
5CVL3YGmflO4EHL4w9N05Vh4PY/bvX/PeboVSYbRwJ7jt8eLW7VoI4UQluIH
HGDbFfhl3FO/9E4jgUmQ2XucuMnEqHG4P1YhtC+r89wSkPLk1Fa02OlR4VbO
iHJWVXt0v/4bw3RhdJm9g3Xm8E8CA3Nr1YHCLghSxxw6dzBXWYbvRA68QX38
x/RKY2HR3tNavsZL5MUt8XGVmwrCgLXJxWMf/RXy8mYOSeZx55zBGG84G9j/
3CurkZlC+rTDwO+uojTsV6dxgUYcOsieYTkIf/TAqquNmvIQBGukxGDnYYvX
i1e4OwUfwoL0sLcnW/O+VExmbbej+8IeNU2NxbkKjf8ux9ttgxxeI1mCrZoh
r+dLQ5H7zrW+AVCmXlF1AIyuDxRpZgkygIKXQV34LWIjQZf8eoX149fRQ/ym
Pba5aIt1FYKzSFHIw6+IwuKxbpLJmm7Z+z3NCh+p6wrXGAOOKN52w3AbhRn/
12+Epn3RHD9qIwBb1FsU9rN1HJbbDKT3rQOs6CqNhuFFBgxNBIM4IaqZnF6L
YF0bglglZ7QzESujEToLpSHxO29OXflCx7RjeIfvPTOyZoAkiOdzkMi/n4OE
T1CKLcV6e//1WuFtjeKHlJPe8NBmy82B4VTPEU3QTWMLRIvo98Sj95INn8dv
WQm0XbT8PEPfR3T7vQ99UeLO9pf0qSz0jy2kpUy6bcgAfZg59Wkri91s89sn
Fa2fvF0SZqtDDXfHxiBMOQh95T9mgvNJirYhqZeCnnuZMVt58d80USgl4Bli
clgMGsPvR5xe7x0ctiAIoYBcKo/AFLcze4lpj9WANRaG6s0/Hu7IAPcie6fV
Y0M4I3cUfiblZraRMexxLB2X8x6V11K4lfQu32/LsnzyssRzwuAi/0XWO6SB
8SIM3HKD1sBBbR/Y1NaYu+m+jqdkPK2jnj/zGbBSHk52FrNlPTbuY5BXP4y7
qVWeZW7GWiUaXZHg/LOAjtIKTlWOhyCH3GRh2FRrlpFoyOOpsIZtRjFGeHSw
zCtWxUtM4cvYM7BWDvWWUbVEuFPmlnJeH6SivmeL08yNErZgizSTLaFuOcYy
bQKuNcX9ccEMPneMHJ4QBE+K0GZtAwjSmb7jhXChHouAAashJQ6uM+rDUP6L
qL9Y/xs3qvUOJpp7/resIlj+wteDvHgIQWbs2WKnBa2oahADW3O8gMDqgJ/V
HrB4O9AAofuEISSNQsefvrx1F6+RClegwd0RzN7q4+uMPeyKJDMfbzKGX7QR
ddDWxyG9x+CtEMLEKFYafo0gQpK/537s7Gw02VAmiQG1vpiuFCKJQqAKzpkQ
5qzYdX17kd65J9K6SCay+ZMnuJMBICnSpAyaWv5mHwJGB6xOm5H3en0VNdRF
uhbg4LztJ+0stfYTw9ELau9tH5nXo4A+tQfdJthsVaRUiiEs8ad4m3+qevn1
OzFRQiYy+6jHw4KMUnbEzKL4jWrlKfQlO7h9aOwK8ZM96KJzsSaB7RryPNya
g/0Va+0WjnfupOnwuwHNX4Zq7JRMBUsTNfKaKVU2i95PkWa5M4pzNxXw+81D
c4cy0w0RriGD4R1FDnG73dv23z2h1NFlCniBZXiQSVI+X4y0WiWC8rEGukKR
oYDTQQs2VWastbZ6AcNqmHzoBY2VOd4X/SjHJHj0Hy7a/rp2/pXf5fMxfWol
O3dr9D9Nk9wsWKQJRAas7OjMk3HBFCjE2kZEnnPdxLYxj22oM+uxE90BP875
4xJr6YuDNm/66hDcFMQKGWMA9x6QKPbeKPxv6gdCNJthDs1MleI7DEVzQ9vM
z6BZn+FjPDg6TZT9hlx0Zdklg2f1A99uJaq0jLs0gdm25La7ZSZXtgcjiWqn
Kz7VJRTNrvXMjEHnX2aUrF/DXUWyAJ/TFN9KKZekArAeRLKYXeJsEQPQUkgJ
1MlA0PZ+CBDxt3Wy2O3ibZatTCU7KoYxy7F19d/U3IUh6BF0X0LyAiarB9TK
M1loux7RCOpZdlRf2uypNzxu/lI0xbnISwXE/Ag6qsU6qlsSh+d/TCol27gV
tMRns0vesJ2yCdl69GSGmcsnxJd8/wMFtPkQ2k/E70S1AcEZJvJ9SlaCEBQb
Wu6EPuMoAtCP+a9GeiARbUWyZRTgD+FFnlqc9LA3MqqhC5nfUI7FDXpPZqIV
LI7EQOUvdkZO5XIyHlyEEI7IXaOVp/P8al0Nv2y7oxGk8MmRzUStxho/Euv0
gbetjgBzifwYjabJwbtSbZJJCxNR/U7z/nLAbjsRwpFDsSqEU1TAzSSjhEb9
RY7WawTsJm6yP+NM4QpJZNasl3iHwNOPh+hOp4TRZfpkicFB8rVRQPJTfIzC
hZK3O90CQc9ZPlKNge2g0OXLNS5kZ/b8N0p/i/lEbLruAV+LVoIyUFZ7z3z3
2BM1oDKVO50paPJR5LO6mv4CNnG7rTARSxHWqm+Z6ATqEr8VlQWTg0jQHsB1
qoa3u0fzBXBwYCPZbMbDNI61AFg7LVnDSmP/lN7sgtd65GL2A+I62jba8egf
3SWh1j5rDUFkWtAXKZTCBBMouHuRWbeKJOqlWyTS3Wje1H6X7W7+phOE5FBB
R2CEFuO1mgFLgBhAJMCFWiGyq8VBNovnZ8IWbEo3yj3DAq1sY1XNg7qnOUWR
hSix3xpN5tKsk1Z9L/RVkhys5Xj75eHEfxKPrIapbx3v9MiWaMz475nO44nv
LAbgGYJW+DidSnRHOfc6ruatJD4dhXJw7FAYqh+UYVR4Dq2TLj81Jk/0Nxd3
zHKq4Kodg+wlp7qVvrLAVcz+wuLC5mP45leTvBgCxaqFRFtxiSPTJZxRR2sy
KD7rE2R/F52PL3VGVIK8lU8SbRAfKWPHBJksALqNAsoOmNams2nodo0S2dbe
bMZKmvVLM6amrd4Sw2zFgfx4TW2GQSm4OieiVfvrrDV3FSen5+nbhLKftcxy
C092sp7z9ubj0rQaJ+c+zftTCRDfFrJMCXmcEdnwnI8maCE9h0gkG9rrH8lJ
eMTcIFwAKyliP2aZbv7ZubsiDpKPtUGfOBJAGklXC/ew26bgNLxuIb8ECQXj
ZxhsMzVkiKb4VgEX5KyQxZfG2ZfEF6avffFFO+KQirP7TxHp5rfLVPKDoEnO
VmlPe2mwIfeS2aETFjdrU6uGdCGnpSnqRTDaEmUVGSo2aMc9K31QhjFq7i8z
+3snlWL1GfD/43n93EVd7F/6cjbLlg8jeLBzL+X8woTNNPhEw3iVJm060358
W6gR1WkAqVfF25ojmSEf+bfNPBHAFa8xHwrbg8BW0FoSV8ZFAFVnOXD7vZY4
aCd5pjC++hKnKAwv02J7oVeh/Xgs780Q1Kj7hdpdLU0dU1MleLJO8+m0xaBD
+aDr3oL+mRO4d92cjG4qrse1ldYijc/Ld5dME0+szyH2TUvONZUl2i2iMU2m
6xsxyeSvL/jIsGcsiepZwu/Y5Nh7Y7rSE6igDjxfIlZ3Fqn0Bn7pBfdQaSfs
wx/LZT/eSUQO73j5QZHA1SyvHp2lhSvyqoINMw4fD6xxXwJbRTOWZa/bTU/a
D8K+fC05H01Dv2oVqEcy359Sw7oITZA2RvmqXQlOaNPvdGaQlr6XoEDH+2tP
7y1vnK1PNSChOYXlefQMpJLDn14idqWunugEO+1ZA0pSAousNkmF3YwQFEBD
RD8YngR3UZHiQthxs5ZWWPk631s3kcdjMLkXzzo2aKZ7QLFwGBqnirbbC+ul
+o32515LdCiF76OoRwa+hvJU+YsYmEiNNt7fo4s1RwQpy4a3aqyr4Laj1o/u
4NYicyvnpcfpwl8v69kT6o1Xl8gWjkhLIe8R9nr2v8brnLh9Qf9daG/O+ZUo
xLVLkWAFeQ3f/FmCp4X3CVgQvZAACTnzeR4Iotvs44Q8gSSwr0IJlwgg+NUZ
ehILLiD3xOG6yOmMRUN26cQ6VtdSdsdg2JdBxpY2ETAlqMLOWmtFuGL5+MAC
GRBAoi923SQJweGBJVmOTSiMHw6u3ZG5Ju9T7ktvRQjnjNcG7YbAUv8Je6LM
YHulhXeV99UraxOWQZvx+mKdbFw0DpkiTS+voIpy3gr5m+34up308zo3mF1W
x5UQQ1f2VPwjr2q2K2yPKQwRIgeaKUu+SqkhU32BWCx9Enr6ZUmdocYNZ+Oi
SOehXTntr6TbPahpXsC8yREnbqtSB8dvEBNHDJn0aCRAOirHlu9IIsUMHo6b
Pu+JKlTZaDj1ObCsGGbXKS7zNmIBt0vx7pM/QEFKLUWIyOWL6HyjcAokmoNb
2t++A/GmVG6iUnOyF2oRe5DyE6c8+uw/Orb/Wbui1Homi7CteUZ1rdN2vpG6
dAP2IxTvVkwd+NN+VArVL8DaonNZLaEXxwCO7t4pwtsSSuoNEbgGQVqd6lml
dA+h6F174JE6kBxfqWkXXOsBOrJoatstr7hp2xQwQdMW9WHji3efk2zQ9Ghv
ZpmQz3Aqt+vOCBc12NFZcHC8cMgkZ0SX/02LmrKuESH7ky+5uoJ9pOMxTPbp
SWJ4XpCEep6R+T0cgaJYG8yMPk52Ga47kbWg5EHPkgHZXL0W8gdEQOMZkvGz
DNVYAyu/BU9xZI9dmHmV+5//oQu1jw1TTHpVvLUQoKZ6M0mGCZIhKjTan6Dh
hGOD0nbMQ5lFZgi6KjZx96yHRm7EU4UZrdujJEQ5cs1C+Q9nWbu26tghMDYj
MA260LHi/epu3uGjJTw1G6oattRRoxRRnBXkG1pz2SuPtH8dcT2r9Nf48J4A
+2I9LsFYAs8zeO2n9nRq9b6aOHpMFeBMPGXoXzowArVuDVJnyXRTiVpN5R9b
qJyCc+PikL/+C+Cwj0NMmq9mjwaZBc3u9ANinZNsO+59SsRiTxCdqHXFPZpz
tIRcjJBx1BwYcYsKkLhCvT117m9xLfPgYKfu/D3ThBuTidONXma50M5cP28e
VFBBeTkHnmRvChtdK67FbnkUWcUdKN8xdX3fAqrwlQXf5QMMY7fg64KODtJA
2BQgZe1fAy83auJgqqYHoECgBX5k/tLa9AcYIoLgsYW5nQoHIIrQXAcJWjx9
Hn1cYuFeRisL48kAzHlBjN1kC6SBNiPMCZznuYPhJdDbLQ5r2WODMmFuAdR2
k6l7gzGpDUhldTrKwKtYGC2PmnHkOtkq19ryulacUan2wu2Aaygn4xRg5xqR
uzmEjtLRUGit/tpX6/1SWQgXTBrogS/SoYLXDG8PNNgoi6S3ZpfCu633DdL7
/z1ZvovIOFTzEZWksk4hyUL9iE6GV+rDUNDqwKqJTtpP0fjkjkVIuE3oSazr
WDB3sx8p9emQ5t6CJZ8zeVmlv7zMil8RM/RpdDvDF/2HBXJxqZHiQTK7JEgX
/m9hX9gH8dTGxTSd9plgjwYvDCwEH8JxnAJB0ACoT1YsOM3wH3ZmLoLW/kdc
66WxbmHEURIAZqPSXY8d9NnU/Q+7/7eACRCmnp0ykoqJq6pWdYDa9cA9+7Ka
eTgCs/jIWmZlnikuftzUulabWLtWIuQP5/CeUR3W0AgfjLr86+zo/DuAPApC
rtLsCN8SQfR5SREf92BaS+bhv1OI30e3jq839Iv9EEiXkAecaIP/C9wyOeqh
rKrK97ob+a3UD17bOHYQF4+tngAfuEH5kxDKZR81S9RcG/IyIC51fi+sW+76
yzFqWs++Qkx7N3TCvOGqd7B72l14AkVg6wjTx8mYrA6iZmLOvt6WEBqjCWq5
dWqXdepCCpD+bpXyfDUPdQAH29t6+2NcgFsYseeHvbUBAH8Tzb5N3LNGCYQV
qpYZrpveaffofvFhJkivkVdXCStPIxJZ8DPimIamxR8VvMiQoOpQxVeBJxbj
U5FRivoDn9JdAAT4tW1mgqhLTf/fEqkrecHjruYDofOZSLPaEBSqmvAAxjf9
dU+EHhH85z7T8lWgKrV4vlH/nPNgZLPThDmn1HMj8jBfPAiQsOIl7EKHpxyr
IktLRqo5DRD1/k0YKhdRAFzNmCtvQh8XRSvGrTr/sPH0IuMpzqMsbyIozMfA
RXhxcZqXnvHv9ou3lOFFsh//furSdFhAoOL4A4xJ68ID3oYE+ME15Zdc/Ntx
8rkJyQeifPop1VtdDLHuzR0EeVLp1Adb1K5SJZSG0bur2hyCAMHQ8MtTYmUR
A4svAj0yPBZH+eIy74pCWMd9hFFIp4/9/X9hyfYNzGuJBEZ5t40G17NpYfjE
+/ymQaVUMaQxvT+yU+2VOEwKiQfytm/lhXqNjAS0l5w3RyMLFXvuetIBA/26
SUbx72a32ZnKkPk3YCsTVVfuTiEHTOQO8qnLrdh+7l7Nsvykv1xKVD/djUfj
Xv4WMS/k9b+gKj5924K7LTKHFlBCNDrrUoPzk4NQeyanYJ4274A+1gJ0qB1v
4NzCbEExVbKY1wF1De9sbHvQSIUB/6tN0ZIxQnvCTQ3+VZmPPUrpwYuwP6y4
GGxEqvDfS8EyyPrcx7EIBIkdaVmxiRtvCtc25Tbdx0C8vDQvSLblnBLPz+ND
OTBaCO7drpoSsRrKNH1YR8li+jesFE57n26o7x4yV9pDqY5C9jXGZj6E6Tnv
Qh1IU8cwbxz53Ixxrb+YayQRlBamMkllddLUMNPATKEEDeAoKBFRcfenqCS7
eNhA0zvZiZifnfPDnYq+56tcYiexplqznHU6LHSLHixElbpIjEexCaeZ2/6T
FSMlHTx7ikGN1G1wzilO81etGMwJS1i+7sKNSe/QFNYDs7hhb7Uy42OIJBpV
5ugidMsSlaw2HSNUU+QtY3PekT2WvnJlIGuPxeno9GY+cRkiwZcnDd8TMTA4
kFbfsFIHpMseGZE/XbST4AQKBZnjw0MlO4hgqxrefkKiq9x2iooNnV1yyqkD
57cGWR/JD1SPl770+2C5pKa+/8vhJqc+qusnPjm/9NCloIFW+vxDpLx7m8Sl
cLLw64RD0Xn8weeBnRrfM8rExQXWdplzRgMrcCtpRQjExex1craT6w8KZm6F
O/ZrI7CHctp/SnCwN+lvCv9S/qF4S31mVs6y0vlpqm9aJ8ZrKEc5CDNKLFc+
fj5+XPSSRefJJ34dMs1uL4NunQBgr9gOvl2ryJ6MfHE+2akN03Dc8VA/mpym
uHTN+RJDSGQWFSNt566zvpkYqHKTzhMJewIDCCL3vECgV26h8q3W/fThHYBM
DeWVqrev5FOODd6PGjGh0EpxQkXGfiXIo3i5vgbJxXv4jn6wuGpasza8io7R
yJDb4FzcULLsHcSSbdf+zQ069MW9NnzfdjYBWXUC4LGVVb8eJdL4B0YfPha8
2fvhryQNAXZWjRgEi72SWTK9C3iwovmr+moU8DaHoLsAfdDtQd55VwJgWb3Z
zcGV4gAPIt/lX+KKYvUvDDXZUH/zix2MmicWDciyzUYk0WMyvTK5ms8te1BV
CFEtWDzsQjuEH5D9kvuAEvnaxguFZKICFdI/NixtNy17nFKffUStlGX8VvHt
RcKGIDij1NwXC2HFUzjvZ/pPZ9lK8XF/oSapAmeRveZeXR6NEEARSyQZpTH9
OHUKmOXSy3qbkjXDR+IysLOBnNphmk+CLNKxMKTyE9ozjKOZioSlkABQC+gy
KOojhcKPsUtjWgXJE5qficD40RYYC0eiJNJ+c6UcItxrGKeK4bjZe/BsHfxn
pPJAgaTGCa9VLB1R2exolh0mnxXEf2rivJAp4e8bKz/s2ne/ySRRx85nrFhR
6h8+CgteNSccR05ciFGlohJIjieDAJdUiyV1aReGSMXod8t+lC6k0/BwDMml
S1PgBjnNWZSrh1BJHfaMfUnFIF1rpH4D9+Jel7CRvSFf0biYXv2qqXAKJn7T
gUow4UiI7e34eFyFW/rOqGuzV5WaOiBoFBb1ayb/MbLrKk4DFFrsd7YRSPLJ
T8cqfYbfaqtKQ5bgNF+WEZVQc9bOXTYiuXnwR2aVDkePGk5amu/99/oMvqaJ
ZHu4hbgAiCMkgR9yCLM6IsZfquCuarVVLZAK1gC/rfiSGPf3p+ThdG8C4DHE
GrrRQuSuo5dQOWc0lJJizLbpnjdXsIUFkRZ0jbz1Iz8+PbXRk+G6dQVCtO8g
m6HPV0eSmLn2pIAZUylHqu1wk9LOFec0YMr/mnBP6t83uDhKoCXt8eaKmk8k
iPmLKdEgpp6SR75TWi7Mb2p2Jb3lZTCsppr/dy4rTltUJpiGep0Edl0XkGKN
jX2Xddf+Vvj2dQlFY2326z5+/rwEWi+KYLJTDD6yqd9eKKzumwi9RmPt5tpq
0kYn1lpeQslQNKSeT97kSX4HpQ5iboca3SbTGR9M/6zt8CnlKnzW4TT3Q0vO
b0JdrjY+B92U/xg2cL0yd0iImCR+LOzPfMdeuuqJjckxcJAd84M+uBAzJ+rp
uM/DRtUSzzEy19Yv1oZ7BLyF1TwHRjTq8o7f6RTXPaBWmrLGOhzXILcaaH5b
4ucXIm1RN4hi6BVTBQLP6+6/revQG7SIeJVHrG7JvN6ZVrmSoDTqCLSmhUHF
lfA8ALcEi/i2RSlx0d1pPM4OEYcCn0DbpZ888l6CwM/Ap50jAaUXx7M+gK8x
ybeiuyUguXKY5y2BXe9fPTomSf88qcbalBrzqQSAQPXDRC2MTwEplaAaS5kJ
a1mrr1DlWh2zoRgtDHPjQQQTdppXijkykDPI+AF0rhA6bB9wmnbvgAMkvEiZ
mWZvOSc+gXtE/TeDhUFqp6G2G+2i82kLBZXf0HBxEnJeYf7fxJGhrVaktPaq
+1bFo2u0v25lXfXTHx1gHGlFej71ea+w+24khLq6rn9THGlWYDThHSBM7BVO
Wj2aZBkW5Xehwz2Hhz/H4dM2kwiwcmcVRpUMpNnHFaKBoBe8Mnd6VsD+41Vp
bqqTlrRSo0chDML4TywiVC9ojeJ2Eq5iu9/OGsa8zDY1xhH/90q+MMMvBCJi
7+KoKAhQTGKbOe1CEQVxYKXO33OC8+G4ey0TChmpk3AR58BZEQCJXHg0B5eY
Z7JlFOuwSgaWRcy/vTxB19kfUX0qx0qR44x+bMryhBNrZgjvHmAOJG4ZkMf2
afuuH1pN4ZSR88u4AApiVveNguSPRNL723tHM51kvATGO5g456FRv+ykdChn
/FsL7Sp90sMpGBWZYKHEbSBBgqPUn2kZfRfG1PHvhPLDXX5B7CM0YNXwyKO2
118vm9k7cmsI2KW7FbLAMyvtUfCPU7hQrbaGxbTmwr04NtHu85jYcq5pjHlN
GIMjfjspnM5g3c0qZu19dMknCe7v1aPZuXoE0X2rpzj0wkGmwjDqlS8X3h2r
Y2rOGiBAn1CNRtUzTw/5J5dHhxz3Ecl/ZCjr702K8p0HV5BN07/GpgoNccpy
LuDX2M/zMS79sEiDywmgWqcrnLkx8SI4+kCDZWkvSw/NzpPvou3wBLCOQJ9m
3Y69//JcW+imidrGoN2mympas57EK1W1smsSl3jQI3neXhIF9Go7zdrVZYMU
WD+1ut9RK1d5jUGn+PURcrfndR1XSK0kD/ZQK0xs/bVeunc7CTVkX0Va+c5a
cyclIsfaUfM60LeE5TpsWyiEpoOxWCxyGfkeWHbER360+B/5pnOI4QAqYkTh
iTeB3oEidd3aPo9VZhAjo056urOqq+bZu7pILsAvaNDTFQrWJKVOmLcNrM63
hAq2FODWW0XzGhzKEJU2SmJTWQkWc80Gri4KDqJaBz48H0Utq5zmpeUhBjEN
Bgz84JnTXW1EPtvFyKOGP7Ys/F63AEc62FU+zcs6482R7xn0cyO+AlXe6G9k
csEFCRTxgJy8EkMZ7qPI56buCF8GlDsPi6whqJVpI5uSZGY8Qni0LcA/HY7D
l1ULvnQiy7EbLbgy0dezKtLIeYC1AkHt5gWHy2zCDM2IfR0bpGqX/Sew/6GI
wnQyreHo0p6+GjlRxseVdTWfbYqtsRbpW8a0ZCgeLx2NogFmTJgdzqeFsCo/
zkM4hp5/LNAGUoR5GzLyVcspJpgJrMr+EjfdMBTJLax+AhSd6LGPh1c/HZOa
eow6hm/Zkth+2C21rrwUqE7vR1L0gvlGsWTrOunm7cm4JOxa+vs2FgvAh0c5
uQ/LtR5df4XmYV+qS6XbxH3gSA180tgGeNk3QiJgXJSONsmwO34q9K+RIoAi
d5v4QKxI40eZ54agKYqBdpzMyfz9F+uqPJ8+7rsuhgVZHWzCb71TrR7ogz4b
oPi5W/z4KiKP00K41X7km6DBk1CseeqvPV7QdXGs8gD/g508Ln5dsqwMPZtE
JIEfgppAFWea3lQxRW+nSkuLducWVXgMs++SlS0EA8nF6EmS/dR6RGfDrt+H
IbXeekcJ9AR9hsG/dfMWbJAkf4v+JKfxbP+1BLxfYo0hi42n7yR08rCzOLmx
qsEawCWTt6qN5LJ9cWMCk1AYE4oArtPO20aAW38GPXfeSSi76tWlM9GwpFsn
Td5R3QcAW7q9GRsXQgd7E9xf/BXLVm1OKr/Dii3U4ZuBbZd7wgITsuamjpSA
gpjvMf081B7xsjAvk9cNzk2TSnlCqK0dy1T8XvjxxxWguyd9e/AYXPr6xF6O
FtlsK5uHw1hu1BRalkprgbd+onLqyxEIXx6qqPvQ8OyMgAgf79wIcgsuR1vs
yCi1XJAdsA9pBjB+k7yMPgk5XNoRqCDy++8MWtoPVml2yfBs/rkzcq/lY2qp
aJpRoc9rHQXh8qiE/rIHy3tDL1OiCQDiJ0mVsc0zNcpz0ZkT9Z2Voo8mB1xA
EDplBR43Znxxss0p3WKUpEi0yCbANhCeFAcSv3s0ngoEf0G3P0y3+JKXOvME
v++E6mQ+G6KMxwc40M1ud6tmCeFIY8vmqGFIZYZ2vWMjJYuG0vNwnlDBnlWD
o+WT47acrWu79XbBJFV/HsRI5s5imyW19UYj4Sukqc/aQp6puICUl8UcZSF6
7DeseNmBkM66EpqNJVhIxIFRiODtZTc/yisLuLfTdewb8BoajNe/ckgbDEIi
5RdLbM+huph/9+9fJ3w9Z9qUwq0yP1gnEjW8qgH5oCN850wU0xLhb40N2zPs
U2LTYp9GQxXRbeWaNMWmBY+iBQxEVvX/+f7BUqsGsqIkHSsujjs73v2CW0K9
KketOKUfNSdZZt9CLS7lIhVYLQg4fXNNdk1sk8o3evE05hED14ofM8xwbLZh
z28ljcOie3aR9dD1rY1H7pOkWFWO1Py1ceu371SJabt7POCbm2AS2M8BMUfk
JbpgKpcROHjaZmxl9jsP0LcOcjCe4ppeZ7RnuswAWvWJoYU7sa86aRJikgQQ
ueroDk5sePW3D+XUGUQ6xlz+6ZD5TpMUmjpRul+NTCqzdtCgkuyaBgC/jLN2
KGjfxUvNHV4k4cNRablgpY32TZBWH2tIIYDsonZCicmcrHtViqqLaNDLII9F
g02tnkYsn1iAjlnlRTm6fin+bwxnRnH5R0aYxiJPr39AxHuTMAiZcEmZmg1H
0S1Jd6t7YTfJ8avux19eY1nXqFNbtzE7MbbIHrTLcWct19lsYZorr7gI/ajz
/dQIBs6hocN6R3qPeMK8zXjGwF6CgPgXVMTanhW+sdKC9e3UDbU0zKwYWD2c
iuAqk5rQ32Sxg1dFQXKuJlr4PxvDSK54e4kh41JXhID6hsjymCpr8lnqsNoa
Bcn87Q9D/0XzVM626mDi+u19WLI4k/X/svmVFU+xaFirIqP970P7TpzWvYte
KibVzitAzngt2p2ay3/tY3OnsO2/Fapm5WK2F1YYzbR+uHFRmBrB3xuPA379
uRCZf+xiwAUmWBQeWt4ik2KxoDcl8wfC65kV3M0dvaFZBBJaQ4xej+AmK3hf
UB3akAfGgRGL8WmP1gh2mFnus/Bq0S3iUfatmgxcsEYQENGF9f1EprQXmYl8
NneMtrSzph+tp2lpYwd10H+aEsRf1xKjt3x7M75dOdbl5nBKiUPrPicptMAN
nmxEbeIs9O0XYes1C2d8mUhD3MgW0eZtJ+Bxf1Os9tKITb3l7iltdI7I9989
+FuOKVBqrbBknri7J9EUaW7Z9t3N0sC+SlrDRdpzSKPbwXWl1BKPK0Xvbqgo
VSbzZTpBrtu37DX6aaRPWFruxXzrgncT2vAmgcCQL3dScUBpV3iBqpXlpkQo
mej2QP7iC4podsBCV6obqs4RIJOHn/fOeBO48FJ4R/+kmaqWl+4aYolFGuq0
Ki+5M2np8JQMICsskiMGSvaYIKSeTVWZ7MqGF069LD4BuXNxhI8UF7AgLxNA
HdVebhYcxuUIkIBq7nJa8hB9GXMVdAxaobx0NQEm0OQxY82NnyRkgKxeR2yT
J/CCHs0SOy9k/F+UdIgUZ50ckW6dNkV7WtQgADeD6qVyjIej6yZ8E6+w1HxZ
xXjAUKdFMm2+if+ODqHwogsXYR/K/dBsr+gOa1GJM0LqrA6CBErrwhmCRo5C
C1mbLsSR/BDArxa9r3qp2vm0oaX7Mv1ragawKSpHcqcoVDDrPYE6iz0ETHov
elcoFE1owHz9RdS2euB1UXGJm8gtXURRGx1oJtJoeDNyHtRRB40g9CMXmv+R
d0feS5GUc9YnWNnI0D8QNdaSzJacit2SqkPp+huIyy2MFIpaO4+OObKfSY80
6w272d8NfWrUfpCPEx0nUFVKTCR8YItdI6SWY2p5brfpu/oHqSsTGYr3RFZY
x8uGCtw7avccnAFkQomieEfSA9NnT1eBbagN7ffaifE/Q4LX7YCXfCaAltrO
WC4Yma4lxuQMlzU0IXPFxhm5oZkvedszFOd5iOKHRWuxmMBFSNetBEd2VNXY
+SvuDSbWo/sF7f64EZoGRZgFLdQZDOYnBAKKx12YENVw4i5tz9c1/NacFZgw
qagX3iizjDUHFnWAK4G90oVWjCh8FVkPhsYRPvcGGIKdHkqgGp2xaRNAR77R
dngqRIS4G3g3qhXD2dtc0I+VlPlmY4GAc3ZgO0UODreljThmKr/R6D9ut/Yb
uH6HsiRYWdeYaTXMStoQ49a9mfKH7vI0onhD4MfUOmCciXmTzjYeAsVC4T7z
c3EYZyOUS8eX6WHF4hNAuVDpp3vOOK2yApU0OO5v+88c4wveSZmMiITxbZUE
f4t4p7bsKrYkWkyuPFTXUnXeT14u2e9Obsfkrnvm4B0rcNIaIveekiTHi/W0
eo2tgn/99+u/4WacjqIaQvKQMNnMj5RxhQqB47JuVn+evc2O4AyUJ5ORqO5J
NWepjd/PRsvQIzL3hV776te10mFMiXMwTvgnnQ6D2KzviovKiYf19VUk8Iwj
wnIpu9wiMpm3wpSPSvxopor8VlP3Xf9CtGrQeMH85tWa8XTqdJyWi585QBtm
tuJBu05PEPQvyh7hxbUSpp3qHYitvohjcq6RH2BvLpSDoE8MZfvUSuoU8oKx
IEFCx5CkwWa7egnrh3cUT2j7prJIK8oisP6wWpqx7nItzNeQTjHDnQy5iBaj
ImyxHdFZf+ZbB5V3E4sRPR3YVUmCF3qHo8m1E4k15wlYSYwySGWB1jOQ0YsC
qdShB9iC3qdqx07rQcVzuMxHl6AhDOg+Z/ljoSYwZlK9cbxpRVM9hfnUGQ9+
h+eLSLM08pkDAJNCB6ZzqBqVaYgy4YuA9BwuKCm56n3Plid/DY9PAXKzN9wx
fpWRu5DvGQmtfD5nvDGrW5P1jJ5jf6pv5Dv4v8CuB1WZeN2NMVe9cRUTqKSm
/0o2X5I7rEqJ4nuFaCGjjJHlgyPxxu5oRRDXWvwApAtMlTdk2z5O0aoB+xlC
2MT8VzQjdYIrpDIM4Y9e5Qf2kTjAEXSzrwLA6ra6gW7Ib0ioHyuntqDQYAHN
8I1/T4mwtiugsfRDITR8ivLxHXEJtYq4Tyd3hStlKE8JEP/xGKMx15kfplmg
PE7rswb8kbxr5FIR3iq+rpeXvfOJMaP1SFQWFbsFBjn8rKHPO8NGETW3sZq0
77hvGT5JSdwigaAO1z8mAbMJKQWodPXabgpCRwrF2oppIAGSvXCcOJBVIhb+
YjgsMeH+SYlQME1JGTi2Fhi0briGTDw87Zxfk3l2jbbEe5wtYf5MO6sWBWsK
zPp69JbIx2KhKTT40TD+XYmtBvBVhYfanGMnqdpj8d0xwYJA+p7syxDlBlz9
Xsf7yIplqwYhkLg/RLLmHvXK9Alpt6Hqm0p8dXSzdIeIt8OS9TnhJHDoC/Ks
m9PVYO5AchCKm6PwRVSipZisaHp2+FS/i7wnKRXG0qsooeGaF6H3lHEUaLMw
VfJ69PiiFg759A/A8lBVVyaIGvklSz9M4EPwuMZCbHIZ4Bx2QJMzCDwNM0F0
mAbkVrEVwwEUbUNGM2w0r9f8NO/yDXg+4+b4rMJTxDTV480RwkphRlJof+rQ
BgluIr9fllwpZMdv5cG4zQT+nO2sWqve9bVdmVJO2Ly3XifdrGkNmEphJKx/
ATltl/bV/SrQnSxQ7CNorHFRkhJW1qF6IKAKWFKqPWyAGfyaSlWebcO0G6vP
EjDxSVgzA5PYcHhLpqEnzEXrMFHzSiL1CSoJb+Sv27M/DselFpXXpbNgv6/5
cKwEt23xYh3CKGOrn8CbglNOk5L80+M/3fk7cdNKhZVOahK/q293J9SNerXR
fIZ4NFiGdBh27Uodp5x8odsCtbmFTf5/kfmAwTCdwwgqRBtU3XeLGZJAWGf3
qhoTNCYFl+fr8QCxXVdqlltbC/KFLDKLT7Rl4bgal+ljyrgl/yqpvcHc8fZi
6VnGgxIkF44649IHXaD0SARydkCpzxwcPVofj3qF3pKB5kCISVMuerfRgV6c
FdRoqPi/BUNWhXdBWKf+0x4DDHaHfI3TSL5qoBLhsT6YQp07L3wWZnjI+BcE
OGNgWgriabVvaNV8pRnqqM1YNnpGFHij5gXVBCAvjVda+uqfeBXDtwMypHPT
02M9dTRLylI38liCDUXrNcVIvYJGMDRY1XGqcUSQ/WFIktEeKT2HvK4VB8B7
R3g1ZX4YMjhuom8QMYC3ddLtmnAeo5OaW1ZtQb5S/c5qVt/+7raEiZh0baH9
bafv3g8r3oPNosJc9CKx0MEkp3JgjMrr6xYDymTOqX8fhekVMrReU1WgO9r5
WfcqEBtXXcZpc7y3fcpyK0fSJ1nj2JzzH1lJIWCIb0LKUadXL/6NfllE5oy+
YZQzXR786kKyz85yMnUKqL9NTcKV6e7OTjUXy9JdgpAN9hY8/hSCy3ro+5mL
8GVxojiAs2FGuhdHx/IOsqMo74Ggk9b0m99hgY9bsPueCRM5lMEUUWTAVfkD
+nvqRlIpL68ZJgfRPf9/AdVNOnSmYqZPU4/GO4RJYDgMduoRgmZMSMyzs26K
HcgYJlnm8kV1ZRZRuUgSo89+Y8mArAgkKcPDM43WUY++wkVcSGKo9K+0fVSw
iVk91OMrBsXR7JWq3L9IpTu1HEJc1KrDLehPLrF8cSm0W8BJxOGJ8TyjERUW
TiOJC0ViLTa3ersuQebfjsUE2ATCUJAI7ayKUtFPR9FVUNeIkfU0loUyEfH1
6l+9NX/zECxp90X1TEPRx6cVOwkmNMhWc2BS3NzPa9auQFTizZnkij8GNcn1
77Iym2LJhPImP67T4ihiEUSr6mYoog923mKF1pAOOtR//4riY0I75swFbJr/
F06jIAzHDnnp23UlnQouqt71XdFnb7m6Ug5VIEFH/PDPkcTJ7NkZHQI/fOnE
98taB+EXYAtMl+HXm2jtHI/90bnThNOhgCZx8rF7LsaVbsveE8HDarED+rlG
nWMFiWxC2fnpaA1jHgf6/VvGPnMF+9BHqk8tfH3kNSAg2n/eA104Rk1QT89k
T7uQrUjgax8eh5ezAb8WaYmcR86kOkjRRNhPWiVtJYQHHWmvU6eSAEqWForL
m7lT+3BhouMk+g8z5XfkEGghLDufp5HlLv0NYdUkn0NXRzIQ0b1O/hyI3gVi
ZPgFhsQyoaqWwX5aqWrrGScuRERODE72v4iSfZY0orJHo32tkcDZ+t5QV5HB
BkKc/yycc2aQ81ebsrSNv8p1JkRMnqxYxncDdqrHh7hZ0rykCkn2jEOu/uuF
MkeNrHyRKHQhDmcQLAm/Ucct+HGxPi05EWS1VeMmJ55FGVwGtpPPPwS7xc4P
hIh1KcOot1wVLxBgxnaV0UeNObrRnyHKYaIQLEi1nM5hDXu7isWuzpgbIRHi
8yrAMZ7h1Y3+/KbZxItwkZeKlUYDPPB+wp0wThtwj/BytgDani6NbR87dv/m
53rBB12rsI1jaPl/eGYM6xfb3BxLSFBKfOkNLqyxJhlO4NZNFiJbz811+fEX
i2ufRG/dt/BgJBDNUzoz1VZX3OIgkSxR0Ut/EeqKjpkCrcNJqYtWxrh849jh
zcTxbHX/4ZvKZhf4OHMwi9rNQy8RbsSf1vWpi7H47qhZMLRX4QdF3VsKcOBv
bgPqR1l5UdAMjWjtbrXB8qT+Vg+zV4CimbZswZrHNWh7ZA/J5MgB/VuvP57q
Fy5Ad03P2H5HUFvzO6YD1/eaEjbabbBdT4nkRYs1/ZUpoXd9HgUo6FdBdU02
EIiNNMLI5dt99/9s7fh8DxByLUzkBjlYUGp0MSonCPaxvoQxnrB1mYFKKkPL
ox1u0sN/NY6FyDyqaF3pDhdTLFHSEuPBZu3GqrbznZoZPMt7ZpQH7cKdRRBn
hGLhHl296ytebPZCGRuq9/SU23M8+bR0h5mmY7ArJHhjf738Aj4wG0dZ1QYm
r+pNTim690Zyk81NYWfYtazWkehqKDyThYT2y479NHjyoLceFkIE4VY5euFe
Vq2HZPzDtaRKmEY498jKSQ4u0XXuPWQr/wt0xnF+C+6/emrZOlgI/dgOaBJ2
fwaVWNLHZQAtgI5HsC8MOCgOvEcNQUoFSyms6NQPeADVr+EGjY2NbqzfcPt4
mryElN7UoNItAfWakL7fb7Em0dGK9nBOryaLZBhTCEGPolFa+5qvFQgiway1
JpL8LaNXbxKbl42WcfuT7pvfWLheeksK4yzEoCY+X/eouPpjt/x8SdRKqMSk
k2oCNl88qO0B6JFx4Mcy6tuopc//CV1vHaLnDB0sNmGEXLs4gTWSK6gMPvM9
PrcCngCNZ0evwub4DHy49N8VPf9VOOAcvY0vLdZrvO9zLp9p+pud7V8ls/Sz
f+Bhk32lzBTd2Tq1ppq8coptKiYNQgGm0kPKFmrdiBw7uheKp37iwuJ687we
vfE3ss/t6uApZV25UxPgXAOnLqSOY6LMBoXbQswoQyNyfy0ww13CKM7+0etb
Jvi7b+ULPb6vPrc6JS09h/sUJ2H+Gp4LNadWM79AdhTE0XVOqHKrcXVasA3b
rw2/C3IJzyp5jJlaUgMVojS/ugKzgjxhk+yrk5ZQfK9C4VcBMwObFaBDr5Gc
nFAzYF0okWg6J5LZtjFyeMivhwYkoGSMBtV3Ez8kMlHqr8gNA5hMm6jHQH89
3s/+zcPkkxBnts8VeE/DzPWBuFGn3xY1UBPCUey+OTfjK924fph5kyKYARRN
yX3A41dEyiofuxpKlDMl6ZjWpD7f1hueLrnGT0uwaM5NwF5oLFd34foldg+P
yd/7PEMX9LEy5u6HjmEiSohk3CVUUjH9kfBgpNwRoNutwHr+MNr1fDud2k4M
QGyojSZRsVQP8gKnlxTnrMmdWh5RUyDqiYD7B6oZXAu1w/RJ1a60Mcr6YEAr
kRqxbKJkH93pvKFwAhbhxkEcaId+ovvS68KWe/a3s+T5konfOsMJsOkPjDiQ
P6mtMGaZdELNIER6D3wL74gmvj8NWIYfVt2MVGzznBAxV/SDD/WxqB9uAvgT
twL6aRF3LxJDwpV2BS2FpZdt6RJOl8vBHysCCz2fFgDmkVGui0md2FEkoj/F
lOA2ZGvGKc3s0zAxnoSmcXP86zmFt1rCKNZcPzd79GLpo3awi6V/ai4fN8D1
4h/nrr3/yECKULTpfwWZgrIgDt5DlRuLFn+reP5TkXhwhd6cvdsJgOBdVKJv
HcYZgmI+tNcB2UJNjQtbtd9spQN0kecRwezoKwdlgDDYOhnPqYXsHQn1KT9Y
eGNtGSfKvVQFR+yj5Wb02PNTyxKgLSayiZpwVxFDHT0iGhh6/UiZyj37/TEn
Hgcpf716EMNZ2AdgjRehFM4l0iNcOmRiBIJ4KTOYv0gRFSAw+6ul5AfxUoX2
zuakIQ+6ZpY5y8m212Cd+Z0okVDE0yxyszpvvrJEPNB5fhFYHfyvnnPNx7+r
gt/kPgbgRYeaE7LSKueZBWfiw+g69Q8vsl0+OBuan/SiIEaa1J3rn74ohWO6
n1RnArFdgSFFE0nBxON/ClP6tHQopKcpqTFPyb3Cb5J+zQtnaroXC9+W5BPs
npBXN/YLxzAPdwYMUfuyavPKh7l6D3ESfEfaNl1J8hlbJwub3i9I1e5cFsqj
uOD84cWzFoJ2+7xi6DV+yJhHqjc7zPPVYrMfimH5xtSiq63D2kkRcLYgYJdZ
rjuM64ED27pf/E7QM73ruUA4ARoVYie6SPylcEQTq0gUEu8s5ZMWW8M88ws2
1bY4d84gxxGCpJ4V4mPu54Xw7z5PF0nmiQFKwXOYj3qAONecGFNwLNNBhqKR
6MjAp/uL5CL8dYB9H8rGglShKeIQJIc98kXJ83P2yKO4Ij59YAWthshySUNP
D+AgacUfONlVnqoAEYJ7qu4GrhjbX2GAyXm6TzRq34e+Ie43ospy79o09y1I
NoEQ4NfrRO2GNxeElHbwG3SP0QklTrWPySLV3F7/Hg3WJUN1lud/Eny9PUw1
nWcLJeTgN4qCAYZkDFseK+MRopPjRQPwplbQ18hX+haUU6iiiFainbUSdSvr
/oMPTP8+ShUo6PE/mBPVK+/SSMOM6UUBYnbAbi8MraqnmnRnA+mtdFzMeq27
S5RUnwsge8HyoF5337M5OjZnr0cbro/10aQLpl++Zjj8xchF5jn0RuB1k8En
43SWPOhCFGajsQjNGtdQtkkqbCf18PXL/CdK0jho/YBehe/6L4vhjkvtYSXD
DW4ypn9SeBhmeJCiWFxJgaBJn0AkS1kRPIk6VEaeJfc620V+N08qkUDKV73l
GzOhYkbiRFylR+FGBNSMb9AklV7KaF4dRvnayT/sBXImIl/UD8wmLHFnmnkF
7VYDS4Bk6iI0gBtYqNNsCYtWkJCzp+mmOuAd+1jTvMmsr6qoWBcA3S9joJ9j
/9FeBwgYyq7lOTR70J5As/MvR3CR4smlvU9RRLARV1igFLU9hGXeTqIIRWn/
2yEJ98Q5EGsMYx3wvrUo2fBq5wmzaEeh33MwOIGZ9nE03IR/sxzr2BiWud8p
3WGgxpfGN5y4IuJ47DaeZRUvnkbBPK4071phEvpWU2ShQBhNhrWbKF+OpQzw
20ws+Q+RoSTOtXwqey21jDc9x4MWvukQms13E+nvj2PWDxsIvSxd5bttIGG/
NQJvDYW16P+benUvVHbBvObP1rGobiVRVJy19StojSoFbMJOCgLFJuBFKtxM
epVotEl+vvlvHbTcjNyC7KyikUJsOE6/iqV1Kf6oPfWJC2KiNvmXC58sJSCW
Ej9RIFRvrjl4nhmawfE9V2+flUcvmEIlxyzFXncz+WDwCUU3ntGSPFbygRF+
vGiUPKY+HHr6LtIAPXYSqL+U/P6zWvpj0+fK+NOhHvssiJbc0ZIOH1N0wuzw
Jch/Qd/WmCxTBA+f0F96Oe4/OE+XZjW9wEkJGjLBoKfGv53SiUXpXJfSBkf1
wH/nxk8StBR8V+Jx2D58dIISyIxlijKUmd1LbL016Gi8Zgfh2szFfFi/Tuzu
w8Cw/Ze0uHHYVHg2qcOVa8qyGrfDJ/rhw+Qr4tfe+9MYjd5TCW0gIKdGPkQl
O+dGV957YB/5QIbfaqSZ4AavkvTR3qmOovV2xZo4FwSBtmksyg6Zvz9uckWv
FprKaezHHBrJeq/X7Tfys0E8egm+ljDPZfI/xRz2uu9/+TUcvlBW1BY30apY
IHkI+jWYS+fYFAGnTVsupGa3By4RjxGcosoXeQ/7tivvlCCVma1Rgep+COwp
OKAq5F9LL9mEgkXWmJYkHaH1vUbEFlTY26kw3GiQujyA+h9b8+J68pAoHovp
SSvabKfxamViUShfaVa0qWI0DokdZClIhdEFrKi9ICCZAhORUWPXSxh/kyYn
lk1ckrnDJr7BZFV+G84hH9Yei1O8Bscx3eM80wQYtsn8J0RtryWeU0t29QQF
g17/yYrb0TV72AQ8BZ4Tjz7fWbPKPtNoZefCt5s/4ox5OTcCv/ja5DlxThxm
SNMr7ov7w9lnBWdWyozepILOcOcv2RLCmkd0oHNTdzbDt2QcaSdEzq1XzKsj
CcaVz3XIgGwERWMz9T/EUzZMySUUIf6zLLgYVPCrikoV4wHq+sVxrr6SAjON
Qq2oQa9onFJyHaM0J+v9ReVI6BXXuaj440lKi1sfDGyddu8+CPwHhjvxBdX5
SHyv1ZZP0jVev/Hrj8W9KQFFV5E5BwdM2D4165ra1MYtGKdBi6khKmECGgDF
7Zo2kY/o3Aa312Tez3fwIzAohT7lftofHZdxl6WHD2yXBrPOuWx+35OmXHoN
fpVaNYgPspgweWVAtsJLYCC+67fYNfgaLFZdIECSACr/A3ZYOf1bMQ7QvjmK
Bdj8VploQJQO+TMcajvtsFSDgIToHb2q+srIa9C4+Leud+F/FVs8O668IpzG
4wAkzuiaCzOBkATfTnIC9NWrPvRK4S+26OsRt/gZIfhOcydivmItUgyDw1XV
s0VN25YIG9notbxw5seJ3aijI2ijRoTt0RupqvAPLh9Ag8IzTsmpSXWPty8V
Y07vCPvOmTz8BVPfeReh4LET8iu8JKVePaY1YJqQQKFku5WO3q4+CkzfBuwa
fsbTjeF8aMAMs1WbaZEU9n5xeED+XZJu2Lwb//03cCYSWn4HAAs5oxFvbFcd
NLRAjJLI1UymzP9QlbHh1M/uHKkTlSfPbQjaVCJqDjARWW/zF8d6qTNqKAx1
3AuTx6fdygDBZc9PovBX0s9pdwGTPJm/SGMZJt6Xo1Nd4U3m/B+Ez9LovBQr
hDr7TWU5LuM9LMBaY+lGeLED+KHtENBK+BDoZhrcQg/UnesEJfAlWzMjAqwj
mxHVnEPkSYBFG0kySDf5XvgyQ3i/K6ErH7AEz2ysnc91ISc+tZaU7IYgra+7
xcD1aps5I0MivWc25N5WQgcf6IZAT951sCQsyCESUwsb7b7dNKb8nokaTg6Z
bw49HErEaFTRBUsA+5+FjiaeOxAN8WGLBHXFmVToUQGpXBkgmeroJGpTjM0H
NJv3t9zOeGSTqtnn+iMcsv5jK2E+N1C9/Y5Mz+zrQSWak2L58gcgi80QEGmK
j33y6znBn4XCzOkWyXBZfQ0dh4LyujQ53/9t+noew1ULZT6DxshfIaSDNxxn
CuBQzz6JYCIBCv5k+UaXMyqtr7gPeIWnpbsXeifjRJIwZC9UT9AzXr+yZ1g7
u8yecRL7M6Dq/Q7bOlLvDRQCUY8PbKFV2ipHli6jv53UPpcTHoQahfk4O/+p
xDK6WMMSHKFp8ckrZ09mGVwxkTWmLGKznha0oeHScS0RSHYxlgYt39xO6I2K
/YZB695e2ajffO7TX3fgHIgReDoMI6B7QglVu0rxDvMZDrjcN/qiuv16Hxjv
vkzcWyZNyhEoWmNp6fhT9OLSiowSLq5nj0dqYlPThqLaQ94VdW6lsh3jfgV2
espIN3qTwZl/CwDhiGT+Sfr9UEZFwNhoigkooWoVmX6X7MyuuPngSyMrl6at
ZIZ4K7yuy2CIirmuKwd4jqkcE3liiaXfl0RuVNlNhWnmjfxJ+aun3sGqJjhg
qlmSr1VMRVfFl3ct2yHFKljrICH3pqkDUthqlF6RRDe/3li225kMlwUVCz4R
HmxVeeC1tzECEFTIf54GMBWS0IqcaB5VbPihe3B+De09ubug+TdOJBqVXbdd
3AF7tVpiLMxu9sa5v0OC8Co9KR+ho87ZLWVqSozdO0iEYjL9me0fjyKu7N/s
dkKPxeq3yC3O64UGJZnY8Hgmn151/n4g79iCbnkblDeZjbix5j/pYRfpDaIB
vPhJh5bobgvDRI8+KY6ECI8it+w4hWytnAl/wpz0G/HVioJOghro+FvKdCQS
sM98LG1sc+CRAw+KGE3XehQ96Sq95sEIJFiWS4BeguWe1lWLrXz6FHghRSmC
4qi6NjtjEldXY7bQJ0gaiEMbuFejxByXi85LfWGetYuNFUrZPg/vZuc/rHWH
Yhx3q99qYW0wcpOCalvO4ySFyIQeJTqfP3pQUTdzw8FjdsuBJ3KbYM1RkBSH
EUhcfHe+gRoVOT73tf1XQzWMtOUdQd11lSEc9belEzbjgU+FILKg+BNIn5N1
sw5NnTGPKokHmWg4ZS9ey0S5o8LcwyIRd9VUUNRDu3PccNRI2NkSYQ7Mal6t
BJcfE51K1seLgRsf5hUi4s30HPfVRiURFzrJ1xrFgvFal8uskWwlK5PaEMtG
FwzGdSaRLVQ3oxjJpeuJYafRRtBw7IWg7h1vzvaHXmtvEYIatsfb2H0K93Ao
c45d7S0RR7cMy1TcfpvIUPwt7lU33KHbLTLphdmC/sYRPSecZ8RaKVTjIl0E
Mqg8b7k58edGM9EywF/2+1i+P60jqQMUk+1RIW6WGcf+BR7aOmNa0AWsZbvS
HF/95Dbxmki9CYlvgBlun5T6Daa5XajDVdF/8Cl6Gmm9BH19RBa+jnsQ9okI
VDQxVE4+JAD+1VnXQ11HmvRzbg+k+6CIRM5isigEXUfs6F14aI+0St4bXWyn
3vfYMOYQcWSajKIO42WN9wjP3eSjt1EvSYbcfGmNAoS7xGDRDKEaqA9cDwMm
YMp8ES+u9Km5ae7DbfJTNCdy4yDuWjSdfdOfm2JuFiuj9ERsmuEHP0y6ceDG
kl4t5m79pPGqje2V+tuhRagzPAQlQ2DDDmXv8IdjE4TJBRVrZr3uIGYZ8Q/Y
ObSF96+DIyZLLz5T26S0cw/JHcQnq1uT6cCD8/jn5CgsJ0Wyvk1LXr3qdcjq
9JV3LmKugWj/Clp0P5eBfuoQ4nY2ABPOB9MP739szScPhQlgYp9JrddtOGOk
wrDJ8unRKWnIdkFo2gnpt9cwhntyNJ3k07+zGgj1Yd1rBFnnANv1HiOsKWF+
vN3BF6CjnLFi5Sel+bC/uRgUuPQIjmLAWaZesgIppVmI/Z5KSuCZVc/No7wj
npFr9yNQ30+B14B36tQhia8YaXtsdxQ8r1JOh2i21Zaye5j85AN4edwSxMwA
56m9xGUp1aJwUD8/NOhb+jtsyW7WTlRHnF8V3KlS71ALdVMpD4JDWlu6v7Lj
GTClCi7A/6ZuWvfwVFn7fMOWdqGErz4Tb88GQtM2xYZCb27HJPAr9vAENsah
GvXKMG+WS9HVpxwGSL0jK4Teq2Z2hATWcCrjvZFe3ViTlnk6crx058cmHlO1
ibO46iSmaicnF0vDNksUDsg7WYOPIb5KeypGGKSMeTacNmE7aSi4ob5Oqfv5
qiYj92vzoomSqZ47InNZSalK9+YoBwj+WNllAYo/GKzv4VWWgk2SRiSFVJ4n
WjFvtw+/Y0PSprt3HcNpcTkMFDVUlR3kSuqzt1FxpcCtF8sf5H4xiFKHlv/t
LHTmjgkTNfaQAFk1uQKBJ2RzrHYpI5mgk9vLaM28RNfARyPH63BCeS7engC9
q4MbQqXlOge9hJcAjwq0G4+DAwb2t9+8j9p2oR3Fd3E4Mbkk7i51ZJ3O3lLD
L9LxXCsyb8OkHFbmTUYf96SnvBgasYZZf8B5mfUmInfL8q+Dgn+D15YzXGjZ
UDH8lgM/on4Yo48PM8osTIniP3xjR9HhaO2U36VUbJNyFSWrJ4NqOQhxuJfk
1AxbgN69fXcKkF4dWmQN5X9fiy21KJ06pJR+wJd1B8cfqK9Np9JYX/iqNnA/
yibcFvYLSa4y6So3HB3WjHzD23QLy6Bct0ZaX7ae1oUODgJvarS+mef+gbEj
3NcCGGlZXdIzfHsqf3eVoo0W7TDsiRfvQ25jnaog4I5u+gp6VCARh4x+Ynmb
Iu5DbmZWY2eN6bsoDM0UtlvB0mtxQM4rxwwQBg5iyN1qrOQ6T/Wllp6etApK
qphVwDqtIuYiHBp69ePvSpgpu80otFf3xrxz7GxeImPM3dktIWY6D86FlYTg
N86s87VBsAQmxYASRRWuhSbHsjj5YsoDxBp4kP26GHQMl3iZhuRdfUXQkEY5
RPsOvvy2UPqZ8HvQqKSTj8P91mT6dziiSzp5GWU/oPBxmAG6hg15+Ohu9uf+
JR+HrgQALcIxMGf4+Yv+pMT/MOepjIX0CVmIqfMQhxomDIqw+fm777tBBtI0
37hD4mxX8LuMBnHqSLLS8asab1wYgRKNtdYj+Zh1ApWNy3Ydi9MYbKdpQHlo
jTdicipQ9M1ewHdQjd41FcwGQ6UvvMaJgXyBDtrBUH/6NZG8uUpruYhdFZbN
fxLDEdrqoLM/acMGGwzMbMuQEYHjTYDpfIdBbx8pa6V1+Hns/qFK2dntIzCC
bm1ixSzdAhyG83KpwjrMzJKtWUpqk8bseGcPuKU7o6ath9yG0n1hc0bz/hx4
tVdSs/TKSNA0rMBLC2fOliShLhpaclQq4NNfbQ+GLgniWo7lIbuC4mdJs7IJ
2pvVBSh2zsjtdX+XMq6YlQNibsBLsMOa8/Y2GVsBK+3lMr3nhQuaPj1luupq
+MW703tdzpzs1HG/fqXx3db/+NI1m2GqmWe+s0scPOVf19RkjXpqEUmG6Z4d
mkVkkbCTv0EnnRUN02vwQt/qlhSwxAUKhpny2tkI6UksvdXDqOy68TawGgCG
u/IUKzjxVUtvKffyHCk2xgR0cnA0FPYzbYr6btybzsxKBMCMXXQxrETAYyRS
7z673ZeHdMihuMDo6j0szkjPYyBrHGyPaFk7pMJ9n2m4WG4RAf34K9dbX8q6
/JnLBk6DiTKG4PVSOOAQrTQ31pdv4rOmB0vzrXhYTy1TcFTAwzKm9TUM0FGK
WDmdlpcFFNCy9mdTotWa3Zu+gzIKJXJJtd9OKAT9k4zfNxjf915rorGURMD6
PEqmbGcicrrOAAzvvrh21FlGayDJ5jcp/kvhjjwrXniYY66QNsX52vDYUQkG
xypIufo9DdAPPNosC7vzny3u3fLqoxikohSDMQzXTavfCm2Tcwo1FGNrmmgE
fQtf7wI7kQJX+AoVAu34pnlpvoepjH3LpYcYcKm5XHfG1yIae46LGMn0i+UB
iJUpIVRAYz/lLmoZ5NybncCTfMXoBtQoO/l8JphhayXpuCIJ4AulZg6+vSnt
okUzw8w1wSPt5cs7fbD7oYe9wD1rvGMDLg5ygmnd2uyweVkB1C4VMm5eSL2X
Ei48/bv18lxUZzJKMZOQ3Q+ozEHiq0S2PAqh5xwlWBmlrfYRtRYfddu+Srye
SIHO2F+jyZO36Ip35X8d5CQ72+p6bGr93hT1vEn+HdWNFjpOaJQ2DMKK/fsY
t7Ii+4Wj4R+J0/WSheAW+2lG2Op/C4PYOB9LSnimrjJoyMVzzF/2OFoIOGWH
iGC2zzdY8law+9qgwumUw6uUCuNmcK3eMg/OZvyXI/RugpXN5RNIkeYr+xBH
JG/3ocSOwAdHynb0y4k8l81T7F/N+GpwUtARmX4KIzCDO5LvB5Jx3HLmytIK
p3Cb44kqYc0muQ2+FhwpGtgGtnyPq5EvAf5EssY8NOHxxmSfjrlMMjjQYSo/
hxuDR22cXuvBLmQifBHPuQHfVGw8yWzpqnCW7L8x5/HJq1kJBp0d5NBcBQSw
AjeBMEMLNe6xgy8ZgHuF+6BF2yKbBNhHo6vsVcUiKSK1GXJr0y/rg5MFEhDz
+UCLngPYxTgQAiF4YDeovxqTqD4vTLrhe4zOFFR8b+B+y+HfVrNtwdMLaEMP
woLwdzIW/TD/cXt0wC0e9nSOFPaTVMqtNx+M3Qx3Vnui8+qamyGUL/j+6PTZ
5p6KlanlaQ53gyU2+X2abQYEzdYALU9is+b55WH+0oErhty/mMPlybwyzQni
0QXPzm9bxyXdfIMbACH+3Fjnfecvjy2zomF1jPudNOYL3Z6djT1tui7/GAUd
wycBIEwE3Kcg9bKW0pCu+Zl5HU7sSLxSZcfHWDhZI7dDuvcePD3x6YzYzDb5
MUrpc2xl7LqLkQSyOfSw7r+H6k2yT1rKzuqD8CAsaaXZD5YKyk+MvWxWyTDk
jmn9r0nVgYQPpdJG8NpiO/3o+utdeGg/pGts94Ky9/R16GSSxDOBpSKd0HkF
Pz2cI1TepnIPGPcLaWx2uhKSOz8Uq3ol24ie1wh8s0M51sqn2uQHlfhhIgA2
5b04dvvPeVoPDVFTSGvLC8i63uyFx71AS1bhmV2GjapPFBc7YN5dZga+2/g9
opvOAgNVAohOCD+39auS5QkNcziLxbCe13JdUcNfnAFlpMpNUki+3l8gND69
MpGCteF6x3RFHdRCzBG1mYOZlrnKI3IJzwjM22j5KECx4MJBFYwtA1xZ70fS
47UvaTzuU7TN2KPfEx69MDlyjvpS+R/j9+CuKM6PCOg8/fjrttoADpRaYsCN
r8oR4SkNy2Qj/XavBLbZwEJwLb69FH5q5MXT0caNuIXc0HdKxZvJG10FzQEF
E50TCtUaaOmusxb9k5lquYPe3jtuszPJeF6wYJI9VTxvX7x8z0v36B2up69h
mgo7mOBV5F4Te8cgqMq+WLy+Mfq314/HLg+PQktaEY6qiW0swbT//GfS3/Tk
T3B4Z7lzcO/HO6agYZHtvOXBdY8dA5l1imStiT9q7z7ryar/3S1e84vBm3I1
WGlQ0I9v/LQVB5b0GvPLvj+w6b3TEhGDkmdu6/HQrRGX0F+pbsLOaCkTM+4R
JSvPqV15sI4P3h/NJwqiMyOtzAMW3vio3COeldk7+5JiVrRZeLw1IUAra7eB
2WhhNPbrZ+ZRiFbtkC3mkFiwhXUliXxFsIslFaNF26TgCaV5xdBetFQLLQO7
azZVRTktn7jmpv/brL2nvOfcy/HANsbAFiyKmEsRfZi/lQqXS9Ge9j9af49V
f3Cm6YOIbIqSZKWT3kUK4yfPAK7lKRgJd7CVry3KDUtx8kE2ONy494waswDo
bDz7Ym9zCHx0bRXWO+T8pc2nJnwRPFAyB8KHlCnqmyKHRm+uUer9Z2PrDTU4
QwNBmm3xuFuAJiYqsyjkBkpdl7QhiLCcB9CjT8G677SpGMoxmzyO7bdkGuQJ
s7F6y3IyqaY0WHY5Co1N0XRMyK3hUgtU2tTwSMaIXV06XF1VnUyL/z3MHNru
QhThp7xfEZusLSAN2CliGINhj1B8VzpfsxUk/sDLYnImzyeaOmO+D6bWrlxO
++qNbAxyM3ChfS52MWOZFwbPXHha25aI01mGCc4nFZ4dsryLIe7RzmCuamqN
ynqt3xKI2xJY4T0+dRJtiMfG4VQNJS974AZV9s02ovLJfmggZ+IBeQ1nel7+
89C9POAVMcpMbexKs8xDjrqAj2+qGOEMTZk215v9VI/W8kdIsTAducOp5H9+
GAc888l/bLC7UDlWA3ZAMy2j2xaur2lC2pgdnw2j+9GOmOKC2r9VhpERA7ED
bDDpjV3u8UBp11YwAznNhWtk9J811yebeEQZ5tp7n/xKujRj6uyeJCfK+6Dn
Cpa80ArRT7gu9fA1Nu5o4oJUmnu06Xd3EBA9qsBATY5jpF/4v/lW2Ztdqz5F
r3qx97attxzFy/hVxmbPNdB6eoKEGFjSLAhh6eqtDWANdiUAx68RvIoT6fHV
zJKSrL4kznv5nKvqNUp9tmMcAlLMEHwKYT58Bgc6KTGMKZSmCm7EyuMAxC+a
XLReX+bMvTVDJk5NHhWvQqCGPzLoGLLPgiDxCWkakPIzFJPNByI0pCYGmDsk
7VBxd0Dn6KN4lIIDpWmWxAySFofRFp9PEy1O8YOItVAT3FGly6+lAVqvwOg8
FuFHPvd2/ghDUVu+nnQWCfN7OqUSMfhdQ0AHvzcMkzHHUjD69Hu254X5konA
BLfC8yRR7Rbfpr1mdz2kG9F6DqPFWNUfhqvNOM+3eoChQkQq8OVLQ/WjlNab
eC4TbQoIblv1uEwvmR0n4Cw8lQ06e+VkfJ/9SNOr0cAJVQvszIsq+SfS3ZT9
qqDwZLwFdY5CAMc5Bi8gwZQOY9vXGeGt9h8aKRz8JOmEpZhdIP76XRlPNZZT
Gbm4OhIvhh4sC/FcgA1+T52SeeqypVTrLqk6fRiUGzcdB2+KxV7YafkQUpRu
pTxrw+kLX298QdmJi27i+TllHQw/rYcd9T2TR+ujmPvqsMszyjK600OzOKX0
yzx/erCLes5DcSXkET/+6wVsq/16lu7VVLAZAbZJKKwkjMrwNlazwq+X9JEE
1Xr+V+TR/a6AEjPFmSqGbdSoBsMqlLXA8mKuXwk60c2vTOIGT2h6dgEMw73p
xqxmlpC/wHRv1YU64t16rIJpPahsdwrPnKbJMelYC3fNj+oVvTiekDb/3eg5
2vlU7pBvXfI8OCMLC9QkxB6xorTTNPXj/P/OS9J4W7snKOLrEo81h4Atkofl
vOIM2d1WZQ+B55hlv9WT4AdKSDoTcDYIpof79FJ7wcBK4u648eB3sQQG+jEB
fkJ6hhOgg4unfT1R4z/9pGNzqQ24/1SC7zXf+I06suHKj6wWUIKbsU92DaWZ
o+OVkzzBFnmbuyCBXEuOLuBOyv0XpB5DpPuJAyYTyl7GUEM/phuB5l0wkhJt
PYZLqW+CJf8Y67zptVU2/cL38m/kD/VaR1xkBt2aXw7ZXCrIIaVr8y36phVH
NRen89cjlAIJX1Gj/S0q8gvdp7MuSs0VHMJvwinolOmuGL3fm9y6ju0/KVwd
FF8LOsLdrtjQRM61QO/hjbNhuL7xaMKIsecam3BOZC7iNaY/pI7CwPL69ZnS
yASh0eC/c8qY3Ob2RGLnnJGo228dt5SP7zo4dRPr13NVa0UqdzN2I2zBfdcc
J30kuW54/eE49mMAGaWKJdiKPIuwjKxuHvKQkd5zNbrOz90TgQ1nJy32bIi1
J6+4l53X/hMRS15cxwtDsMmmZbjdUEcJ/k5m6t0NSmv2BhGYaw1MFqqQxuK0
/qrJkPddkm2n4TiXYTXqIA/Xl1gBcLpahNCA2jJf1LenpfucJDTvSM3UVDHG
0R9L6UZnWL8/lvA07o2fInow97ub0zhyuveJuEAmlmmsMvY1TNyitLAga4IP
MgB2G6VCVW3XFvz7TTq/0KRtVBBnTls6Z/NmAYdR3+cdue9EhbDFVm0Czwpk
mxyflvI7o2aY2LUBDDTr9p69o9usk4/LaKPXDzxRjLs2JgHnlk2Z+boqPR0m
isstgKOnOM5B3iO08BI117/sIQhw43r2rEbXfK2GfSI1lMHMejfmVI1wJi/4
Fx5ghJenDbtDGqBKHa5UEe7k2bJX/O/I2EiW3VZw1cBM8M+elATFL7dHk9Am
h4n2rn9vwx9dXbRDq0TLmj+crUkGgdiSCMncisFRFWCq3PJx1LPqUz4dswRw
9rUQFDB5JoncylzQoxS0Y5vNFdKMqvxExiMlVX93nMekZnz17y1/+AWFDitP
G8tq9Q6LPt3zI4PAdHvGrHpyEcIsRzy4lyFucKGy7UGfOorsUbzzjfOw61H4
UMZADDJaZK37IjE9cI8jDqEpFUsHdB1AwO0PkYIA5J1SOdORcoFhRmM99Nbh
JkQlBAnZOuObXMslsv5u4iy/vNYuqMMrmFr6wy7cAKvM+4HOcehXsvZNGhoZ
CMUZlBykjmqkhfEKePC4+Eh7zZUq4vPyze+V+Y0zlSL0wPjGf5ynV+Ve3lMS
96555lJvvJW0O/58EDy0whMswY8y6+TfKMmhSGOQCNySucoQBudq/y6RSQpL
SUxq8fAnC/pth+gQ3TyVXuNGWpEqiPbeU/NydfAVSMWelY4wa7Z3JHSH2KOJ
EM/6Szdx4fU5hIrO2B/TpIK+VeF26iEZcoSy9YuykCDKXUe/F0mqBs3tWZgF
AWNQZgNKaHYno7UZLK+GIooToEK4CVl+aRM5yg8ZzW66+lKkd7fuszYvcymi
H2IhZi/EvKsdBZGrlta58YuI9jEe72pzzxccnBpgC8i5OC/2haFotDWy/JOe
3zqnkU956yaIJqYZ8CaElUpRlfARGDOBUff+B3LJctQ54cr3KHoetjHMR69i
TRGQPTfY4ZQDIIoXBedJ02W5CM/kqARboi2NAy3DEIQMW1vlW4U8g9PcW48G
nGc4X1GWYlddIHhUP1m8qy5/drS4GkQXrl0R9/Jcppy0qzgQ9siAZE2j/0A7
AyemHEFOSYcO9iu7UnGbwhvklLVZFyghDDubkmIqdmYdSxEEpmloxPPR3frm
FAIgMmD7yclpuIczY/OY4jptt/xhjSvXCBhApfhOjPTRVkzLpexfaWRUB5wb
bRdVoJd7DEbonEHr4lOnabDTNuyUBQPZFrOxBTrYX6TWcU5DzUPZI0pvKIPP
JhCg2LBjCGgqHVXdcTZLsN2kDM7u3G+mAhSW+KS6tS1NfkTMtjbrDBB3lVT9
rA9pnYnrEORFcEydd8E57cGkbcLZ+dL4DJt7/cWitzsXUDhEX0yhfRJrhtY5
hxVkFCdNN6MO2P3X+k++OuoNZAXCg+JBS7Px7Atol7uHhnQAoAorwoRZLKe4
aDB2+f8Dild4HwSscKL9vpMdcIG3eluaDWeBjSnbxoaLCPaaUcV8IScf4Qr8
LYT1E1GQVkNDntxjkwOp5AX3ZA9K+1Ws7MqgeBWmiJl4JG+kI+qYqBxRnF+K
+L8WN9qNLrKvONWgwy8lcp3PgzxRFev5jZs/WbI5Q0wZVdfJaxsJ2Zw3l49p
aHdR2BVY0ikE+KNLLokzvYfjxvqzwiA7rydJFKtkjpiKfium13ZJI7511cKu
/lAFItFgHIlWextBLj2rqIREAeHXocolOprQVpCqm3RHjWUJllVIwC4Rw1NU
aF9LJXVE0fvUzGlEevaqgyt/HnxYNj48pRsf4ulixXAUtP6I4rcQbiiBBSFq
zGOpsz56DqVOvPAVJPXBssaUR9MmE1vgcLZmculrlZDqPZQF3jjhX2U6Asb6
W2MGG+KwXqWQWildNWq+3QyKNs9IVLhcjnxFYl0ZEUBXkOfCXuxwJe73WaHY
Zh3+LKoptzFczQJZhZd0+gSbujE7HLNNA8xMXU6D6p4/WHcUTs5HKqOrOsCJ
kwJRSOuGwuCch5iK99YVJV0k9GXNCSqiESL8TmvRNTXpW5F+sNbOHKRcG0fq
92yXwLFtHgreDFdhn28mkAYUGy/ZTGs4nQ9iRr2EaLXjecN/0nc43R8OUJeg
3lXc/jzNbyaRdb4IEXkvWbEO6cOyEgbjvgVS7ktQ/nClCLmsLfqg0zTJbu6x
1pB0s4AVAa5jviTFpo9eOZJBzrToK+w8t0/kbCJsZwxnXVEli4aIJa7rHLLO
Tp7/yMqtGb+XhmBM+83wc0WvwZ34T7ccKK6DMpQpBd3SNZ8uXs6TrBfwzhEU
urSwp8Rkbho7mANjpg+KEenJTNlMZIJAsCfUtWMRCH9vTPffsfYxMFGlYJxh
NIxkwH9Txi26qX7/6XDy9yTG9mWFBmO6mdaHboNXpHxtnM2vgaIQEiZzTNSV
t0vx1NGQ+IuMFGdwPoWl7z9moCy68Zef1m3qcM4awv11s3HldxLEQ6VNisDZ
1NqVsZlGzUKjCAgSLSfq+ZMIes1ZU/vYQ6umplytjQyP+it16vDdQyTg3/Bl
OtHrDCTr1SmOcTpwelNIqVZtn2DKt8C1kIUJaE52SVLjIUuJ5Xt+HoBXOZse
hB1yzirA7xGMz0bfQBCrEVTiiBxGIvIqqsYnFLnvrjyRTwRtQ8y826vJcjX+
/jU7QW4D9bFtKhIK9EwQ6lobNpl7yy8VVShff+NbUvmgjPT6r9+kEja9cWjX
ElSOmy0gWpzkPfTL4ad8B3+gQbLsS8uR0529RpLdrJTmKh+RpR1aO89rEuGb
dj9KUK/mkWUxy+wWEODgVa0yDRhEaetV8i7p7arn5XkP6Mx/l3/lQrwK8pN1
SgsCGLI5K41G4CPfa+OxlglWtY+NqE9XXJBUOJP2Jz9punQwv8ccyspqvLLU
GhKvLiDClGNhrqzGEG+Ygk5yQ6ED+kSxVpFuuiuSghrfHmkhY8dTSSqjTJUx
8EAZ0YVlrcL5gHNOTvq9gu4jY9TWKsatPAwK+po0jiKm0Qd60Yr6HurwzeEi
9b5uomdsrKeNbcIVpgdXxvle/MozTM46/ceSEuhZyzaAVc2lMgLiKxHalgn1
x+SvP7AK8Fv8+omSPqnsQniiCN3+d6XsMoq/3k3N/ec+HSVX5bNfzDzKm52d
Ff/tBOP+h/F4GfjtHhVK9jty49Rx741sUrodMZXiPnKrVNiZ4UgbgijreqKY
ub2Tj+TFw20OBXcz+JISkl4Q8VCulRRq8xe95QR9TbV5XRFoAF8MzDS8AvNe
YdpoJU5dtdYAplkJtQltukc2xg3O++PF9EiI5uogaMbWRe/Xfk33PZ0YhnfK
ecNAE6oBbCR7Jjqedsb+yumfvHa01fd28wUl0Ns8f31tQrZYOxAO09lwY20H
N8YxmaRDh1TuM1fQSlsqHiZJ7NnTGbcpVIUBmE+o+3XdmKZI+u9OjaaJVg3Q
8Bc+YHdMqcCg5GLCeWZMuwYykqpyvAjcobrXywpR7ZyzJdSMpsJ9VR1fz9RI
c4Lh/DcZ3ocmvSoi7/dHUYPKdS6vHHk32oxcIZcf2l+cAe8zlpIvoYiDwzKI
SVkit4mOpYH0yQTp0Dyqrg/ky8IFKCNOJpVBghGpJBT/u4z0sRkvhnTZussl
5xg3KWm6VSXINZ+xRxqemMwLokdkM5VoC78vn8/x4HTzE3TKbiVUhfFV48Q1
RRwGMyT9xmFCHiQZM61RB2PmtivZzPZSIOeMzA8XpV9bPpBbt8rKElqC9oI4
h7J0boOqMRZpV1FHLcIp/KWrn2N2aXtFPzCHBRX/o2ieSY2qFspKfSg+zai5
6hKAh02quTviVk2SuR5sTkoIKHQSgK070stLiocM09yCszXFFqyYmJH4R3He
VQaEitYIzKo8qGBij2LEdUyN6PCrNyeVatPKkRXKbtnvlIFotrdzJPyNwt8J
RMbGVMjIScXRhus3hMTg9qMIB59gs13FUPwuAsd1dkU7WBHpTWwF0AFPDWjF
sm8HmLB6StiH1hJ7xrdLV9h4UQmlLFsX20R5ai9H1vmcooxjS+LXY5K7vMyG
GHKm4OFs4NMkVqYDQX0rGOVGTYoqOyOoYCpHtZt29M8WB+5xS7qSGYpSueJt
BGWXLwKmzvOw96C1YfHFY78jBSu3gnxMiZt+RaW9ZVF/iKj0F82tW3/H1Z3B
JttS4Hy/TCtC1IDPdd/yMkPMBT/d4dNzyrZahLsSu0QjwvGsIK//DmbVbZ4Z
WMuyu/xNs5e/wdunWzaMAmUAYtJ6V/p8LK14TOx4drlM57WtdSmdFARrTVQN
/b5ZvVb5xJ6hJ/R8esK+rjAPxI6FgamL5ro5K2GZ7R3c2L+C0iELqpZXxevI
agVvM25J/rYaYS0Fqvfn2kas274koLLDhRXT2zJ2t49jRm5VCzVWIWm2A+W9
LZcONWGpbGVNCOkTYJPkz6W427qwSBBpoHjFinmO8ZXG9fr+/kixGA77S/eq
6/GfgZ3nkzqbwU4L56KFbHcOz/kRRgk92nAZO2kW+NdUU+7t3xZmbqr6MrD4
9GPf7W1v5cwGOUBW8VAzopuSCZsM+KIsxh1BHFAN9Vg8N2fN8vUd6wMVr9Bp
jgFi+0uEcPwsMQx12hiRgJtwsIKL7PpU+xcoTaJRQoXNK5iffM84Np1UXEK0
0aCcFD08k2XJh7ZY6Z4BDx81DT/CEHjFf050V6AgpNsjKxBvuNfWdlfP+xe+
iGdpAaT6p19lODM6RCDofQKqEZW+voFx0jarm/H63ppLs7jlMONuO1+BCUg4
pHfbkPysX7ySfFRM9QRL5Kk7KL7QYTIcbFxqnPZUk2Ud4uc6W++Z6EkD/R44
cmhmZNsMyBVJiwS9iz+ZPLdxT5Fm/lLOm4v9uNck0vkkmQj262vM8tzCvs6I
fijUxYlrJa5A8Boib08wuDo3JOP5UzrI6dDgGOaCgSM0BVhFy0mrxU2iMVll
QjHaP6WROIDOwqIfr4zFkNr/KihPK0G+w4N9F6tvy1aKstCPiqAbSvLgR+F6
c8mZoL1GWMZC2AerusdAOJL8rWFBBak017wlh/JhTDFwNxvYRE6EHaEe+Y0I
NgJZRrzjUGEg/QKjP7h15DJy2B5gvI76Q8lX/qjLHTbHAfBF/BbMul2s9T4j
nV0OGvrIM3U5NLjgc6wVqRabDXzldueCKg2ukpNGpgcY5tl+YWy63jOK2U3A
YXCD+yGasMhzIUaq/q9WAT6OR1nLzDg0h7AThlxJjq9GlxKMesTGfIZiEuDW
KwLB8uo3NRBoGHZ8fYrDM+uh+jmUrhnmFWVbGEwfpXbTHh3676mNMsXsPhUI
j8l3TYUljGExE5VZX9jx48Hjq5X7IgzXSOGTDaEZxA7TtJxnrqZLkcW/4J0X
2A5ruNokYSCQWJhpbZjDmckGUi94iAT68kiMner++lmLAOAWrnFESgps4cJO
dJysSWnG3vvoCKQyJRC8bkm9z3jxuHx1seq8wqYLawW33dUXXUKsdJc3WdRG
JZTUhw7IoAuxC0l71l6q5vk1HpQc8RApDcCh2h3UTwX1hbHkjsIfqzpKZdMG
8jzwY2lF/gQFgpsM8KrWDHZlTNRP24k6MUrNq7VPA24c0WX+Q9sYoF+9aXtx
Fw7cjDrjKNE5JkG4NSjvRECuCTRjEH9QnJ0e3t+JZ6VaBmgvM1+hQn6SbX4f
e6QJbFN9dWVtpmacQZxbGpDJlyRe5JPVZ/8HN6c/23tEk6AILKf1E3deYSgV
xieHTvYIeG/Aeo3cpF0TPdEe+7rJXJq7sxPTJiv4KPkLk+2JKCQGrSGHYDPz
qygkX6A4We4GuQ3nY5jBxCXTDqtUznr7uWtkwI+ahvicyVzvynpKlgpzcTAn
T+n8HoVgk3TNP4bL4ijOA6ZQfM3KhI3dTaUbAxwKPZJ13clIwaTSH33Oi1lR
O8bt0OldfJFBkqiEZdqXCXoeMs/vLXNhWCzbfq0zYPAoZSN9st/bbI9EBo6L
eAOGXfSXbtYczFg8oUOfK0ogB1ZHMaOqenJ8Aw3Z6hGYGo3zqMnLIeFtIRCv
jOxpnXnO23UBmUuzWMI644QK2TvDa2LnXXeX1EnR7XEe8ltySWQUi8fL2Xkt
h8fuu3C62yVw4wUer7Zep06QlQMNfuWOcNvoydnM1bseoDm1UakL0KDAOS0+
TuUayUm5NU12F/XE2LtOEDGacUcndR/16bh7ufTwjM54DWM+8rMYBh04jaAD
V/mBLV6Yo3oLyZ4+WHqwqIhxOgcIwKVhYFbEztH8UwMz+DB8x68/B+CA6Fue
OM5P4k8Mh+tZCjhNvhKCRyNSge2y9X+ZUXdGvcJbPMGN1M/02T5eIrNmZMR5
QEwpSu2Xb1F6392lcJCFIpGqBQf+1NtVNtVDSgkW9rE5BnOwlExEHHsV5JlC
2AXXMZg1mPr7YO4/XOjm0kABdWEI8r3wHNdgfebI1wmssgSYGNKNhY18kxw+
3Tm8IEx00OOM8npDRg6lHGyg8luy8sa5mHzidsPTXW5zoua10QdOeTxOLbn+
mYNdJZkzcY9cmwgVqFLucAKUhuLHNQxQRimMPdDwCoA4hqpz0ZBwchIfM7nc
XP2p9SSAPEfLCIfRQk9PDA4x0hL25b/QsQSW6MwnWdxOF4kwG3kLXQbEkTUJ
pj9NdpHlp9TZziuMJwN6/C5C5rooe/YoOaGTLvBGJO2ZRIRmM7VdmsWU1sph
v+f8hbWMQVb5rWXIFZMDccayHx3xt+oHZETrrnBpfhjmjAlY6kxdEKcq0Z1v
R/PhQ4hKN5dirUUNXSsl5IEfenEFRqET1Zw1Eg7BS87w1mWDGptdtmrNngkf
CiYNozrftuJrXQxJ3F6JaM1NLbhfiVJyqx5kKC6Yy5qJ3qh/iDvCFb7Pxt0I
8w5fzAA0VMwrnyp0esJlF+j2nSGZ/x/xgCAEDzKI53q6IjGvGRkPupXWFLNM
OMr7yzA+hsQPhNz3B+l+Xoumvj58OQL6SkpwH3B7G8mBE7S1LNefXUm+kunk
peE2fdWChy6+8dK+34obVSkgLsmsayb5ImGJjF3eb5LIHJeX3/7zW8AF/v0e
jlbLGClUYEitfNJld/1eKe6rxklh1OW/XzWuh65dopKaeXMLM9ZFeWNFzK68
vWiJoupW5LPzxvf1FWaDVYSAaKA0EAoXAHFXUbnC0jz+JRYUnb5bYZY5M6mF
fvqmWgCzQJHXRfBBuGbpQ8+Cp5Usymrbn0+GZNozAgNfzI6qZriHc0E6RVbQ
KBG4aEvJ7Zgjmvw0BuCHITpi4xSsbYMIC/2TNtiRi4XF6skezJJJCjqn7kPv
ZK6/bZj+TKrZgRzV626rjCIP3rkVU3m8iG1O1GjLXSHdALWrXSeQNgBxBqNf
KHak/HkIKD/8kc8Uqg6yH9xf6+5bZmpKSVVgQrMTjVTKudGyskIRiHg4+q9I
3V+mBBDEHDtlmCQDtJSfkxAOQXH9MkmFtKgYvNtlOw1faCtrIOFMyPmYbWDy
er06RB+i3xyy3xQZTdZ6WcoSQKQvvPPspehcPg4jdIK0DbZ3ssISaTJ9RHwG
Zp5ZLp68DrG925qLd4LQNgVx3Y5HyuSu38os3eo0fFWwTwKTHdCaOzwlFGzk
PANurzsjP5izCKDox24302pPD2FZ2Av9StSXvZadbYpDlBL8vu2PH7Kso6hd
n7NUjVZXM2Ke1Ek9JROHpMWKB7KS2DHbtpopg+PXCTBNGLSUj9+Jl0WBpwNZ
ffrBvR7d8OxwBBRslDlw4lipJdXwTK0+l/z7Mc4W97m+ffcW5PPmO/ZU8heL
YfhZp5G4R5jUY3JflfIEj3cjyS7B8uH4R8e6ANc3Xi8JLBA8F0dbgM/6FSt2
kmZ+QON+WxUx3s8WMG+vKVlnDlL4Y0VRC/IPNMgzc8VQS1AA0FUQuS2OBUem
c1+lEocrcbPwif9KfcoSF5PH9nrKlBxTX6hs3bbETixvqOEz5nBU1CqkI55n
RWQzyYz6htVT3NSCNWZv1sSDZqhDBDNu1bKam+0OSvzQw9HXtJkZuhPeQI+L
L/xXjh2xHo6ITwbwPHbYv9QIoBODzenfgPyqgmF7TUr8BRHA/Q9x0Fnn2nZV
HjbHziFnmIQt5GuZzB9IsoSjtsOCbAJA0qxqQ3HCunoR8fhbc32ET2AhdRT/
yytiKj+YtY/sBuEkt16q5zrnTRaw3Cr045jzXgw7w63OFlgrYd3XoRJx1Ker
XJufMTOa6aEey6mZbidvPDRwdePaqIvEJQLG0haoV0ph+v7RNrcdP0f4+U7j
8VfAsRHnV0So+VC1JCesBx0829cjbPhObH4ch1EQA7YnASZigl4bntsgDlIM
tacWGNdMwBQggLrj5aZ+75qVA6CKT6Rrfwfzgacyy1ZDhwWrJRR4mfJ4Df3f
DSQ5QWD8LIhxeLUAR//5WQ+3joT2cu05fUzqX0wqeTKu6mTMPyf/G+2mrmnj
vYpHEc/rc/eYcirBdYrRhKwBp6bX+8bb6Wz1ml00ASC1Uai6WawRXVa61DkN
tptE6kGFboumGqy/2PF7UyO8iIu+D2TKu+7Q1UfO6ot+jTBkXkG4142FRdiV
p6BS1WGmltyBY1r226htVrKStHj7dv+alJp7LrOfa4/sIUCWzgWdOwGO/5gt
gzGZ5SvoHo9wPuRpROVDoV31qQIuQcwqEuWO0iIf80e4SxZshyljUcbEhSph
IiqT8+oT0CYiHEt2aFXtLrAX20N3JmJPGaptUn+U4nezh/4e1PmsAMdcphlf
bYIMMQXtxER3UX2SMjCYO+qFBankm+FRBpicUc0ROM9vDc80tt1FBh9gwHMw
Rhumtb8g0TYGoIZYQVXuT/ejs5jKs0G/PTw334cbeXFmpzN9Ql/God6nJBAw
J01tFzUSDt1mwbFnV1olo5EgGLgUZzR8eX3ReNpH0NeKsJOH4DQwHD9R2YdK
h/oocAF2OoTN+eWFuZS+J7svh++/+Xlh/zwjgi3C22n0g124fE2p5idJUoZL
qMPaEIjgbk73xbdUGJd//z80o5VKkKZ838WjyOzVU3Fq3zSq1fvuCJe/4thY
F4k+6Cb65nhU2rxHuFDLWQS8iPWgVRucQ0DWkcPc4fHlNDdbAEQvc3/dNobe
eDikV44vgKaQhQamtute3HvXypMhz3phsmuNJFjkHJ9PsbRsWWedB5dfI0Tc
KXF6OYY+KWW1Yb0kQiLJilFj2jZm+EUExHCp62yy+YBv0nKsWDiDpET6TnxW
0W83wVxJbT/WuyetROF6i89jzIKCC/ySKgEakDY2qWo1nBT64bClWO51bDTs
lVnsoREH/tFL4MrfN/x1jbLBuouFq81TDw37/RUbIzHLdU/L8+h2BBgXYiQo
9fZiml6mDEnrll0Qw6IoJikfcd4X4adxLplGevbo6c2Tjtu6ax5MEh4rLpQM
mul9pPe7dUZaUED4D8YU3NYY6vwNhOY91nHBOGo4pWV4J6XReJc9X40G1sNc
Tn/PoYO1mMCHuFgytNLtlZBUMaCDOAvXf2XGqn+5gFIiapTEfgPGrKS4I+Gp
54h3I4IJNZ6j4zwdb3ybANu46yp9Z2FWgAAoJ/yDW4WM62S+hXezevFfDTOn
RXAYumhDX2ZxLssI68dqJoPd81tIH8AhbCyLuxo/QHvnYJQFWLmAazfu6l/F
hMtvzLfMk2NkUbdhOVT+UWyhMDgvkIu+RRXfhLKSTe+DtRkSia6kauAr0C5r
R6r9L1hw6CZOHtfCx+JM6lgPkE5WUcYc4j+N/HvoK4rtyT/yBp0JIu4RONmc
k/jJiErbB6Tck+sINi9MZFI5C+0jgaG/rPwz6bYqtUof2b5c+s2Zl8L/13EB
+jROoE2b4vrd+9bSTHoEMPqBSkFuBN33SYmFYD9OGVGwo4cYUg32TsJx3+4j
p9Ttw0THk+71C/s5iRIDqlSaWpk7wCnIz8XnFvKnDDdzQ+ne9ixdaSK1Z74N
zwW69Ulnq93/FwsMJZdDdtpjOXj+YFaXBW1fe9f89aIi5x3gDxo4N7yltl2J
auKDcLT8Kia1AhJaUzhXOvk6JeCIEhOe0nq4xRfkm/9kuy3lO7xVW06POwGZ
7jOtDbv+oqzC2By/zD1eApt8egBMHtqLy4+qaA58Emo8l0ZqHbgmm0D/E+Dg
0m9jOCrEywMO7X9hHxbm+E0AxDGTadXwUk4Lrgu8ij7zGYauVaIsIe5aeoa8
ub0OOJ80dbInOZ2wW7jbXdTduoU/wmRVeMPltzHSPgPjk8iLX7Nz+XYA13Ai
/24OR7AXuUdLrkpzlSMAISfQMdzAwdyKMcVFDja8lICtCWDFopFRclZ5UdFU
2NFD7MLJ8NU9n5mWx51cn2OQ15QZ7yYEJhinmzddf8r+E6xBLR1RLbY9Qd9B
YeUTbmVsHujSqUIpvtLIWNX1/gDkKODihVduELoGx2EfYVNPVG8RSrQ+oCuU
D5YoQAJTKfXWBsIDePD8I9bcqCs3uHg2jlVjUSclSG1Gnb3TwwLejLyFvpqR
crb+16F5FwHHeNWDVLfWb60glBP66SgcfHH2xBwVCUYbguIeTUP9kuy0f+NH
88c0TPFDg6hYNVauESvSuhZCY/qfYltpblk3fCdWkCYZdkHKAfYRpI9QF2sG
5G7PHhqQWWY0+oEpClIJ8pO9eJSiCrzyntaFrhQM+5pz8qQBXuQ1fEA005LS
lhx6lmVZFFfhcg0HzqELAzUOra6ZdznLgVhwmcIsCU311aU5BfxSy6BsUwAQ
1NlJxNPH/f6a7RTY1r7vjqJ4uZ9wD5sooonVG5UYwLNA97W7XWOCHD8V4v8s
bUsUCtptGwGIUY4hp/jg0GRyTZknBoQ0T3LHDzuNg1IR83TKaC2dJbVpOjyp
+70lTKx+ybUNW/u8wAuIrpqp+ZBNizZuHZeor0lHuqortk1LUVzXAGisqxLV
IH/EfHHVtAcUDi0DIxLHQs4zKxwRExI84j+6rIrDqtA1t+LCuFtnUuLBkOGf
Bu5qn1fCA26NV5vramL4lCn/mNUZ1cnYaYLm894K6m6S4WsjZdFV+8L240kO
6aZVoWPbyCnX24Dcp4kwNOzJKTWdrR/jr82CK2pVlqkhOXADLsG0m9UgeBBD
MfpAHVgw2QCGpB/SuhcU7uPBzhze3/pE27HeTAGPMQcBIaBjhpnF1p/0PYYm
r/mgt7MldOds9SxK++m73r3jpJmmPVJCyreB2oLTzEPpAzqhmPdf0tWt0GF0
LIK67cnsvrRF6ofomipINAdsCUZA8nevv+P20nmKHCmi7WTv97/rWqfV0247
JkUlSRfOfGS7LKXHViC7inJ83sxLXED54+5dwmNd8KcQemJfa3c7vr5upL8h
95t6x+S6MNs7zi/wE+3M4R1tzT6u41U80EMg7Nl3+nuVsDUlx3iZXXWVDRrQ
W4IbF02zo4plJYrzF7Mqhdu92TKlMCeP6nUZnFRQAc+B68/ZjKtAR8zXpi2K
EkE9/vFQ+sltObudSsqRlw30oufLBfHKLvWdh1x1aj9cK8fEXL+2Rqn6ePnJ
yn3f6daqT0lmHkK55qtf9wBmhqS3rGghhT8qvfKVZZPelEtIY7xzQiE8EqIN
zWPF2h6ozToU0xHZIXx1akybtPc59QVKL+MbSuUecWhtu7YEQFAw50wS7xry
OYrRxvyN09J4xF2zBkuKUO+d9mF/p4kT3HvJ6d/jBTwacEP93ZpHu8ZzjQDU
sAoyXU4YFD5nSyNOE/idWOlg3bSINfHC70GRSLNeH9zEWG4Mca/ctTOVKc1H
2DFpfvzUOtAdEUZuCoxqQXOhD+TWeZgqrSJ8TPKJm3JzDVnj+eB6Un9H26hQ
S6WkqJ0pkKC9eOklQqEF6QaDVYKVelMGkc43TBHkrKFKEB0X74cqURF1encv
9Y6c6Z3+uPW8XMt1iWKcHlMg5glgVy8YhkSmY+VcEJ0ewKY+tP5PTvRsO4Mx
CEprcnwMBWAtSs5H7Tr8Crs+J0tsHqaYNspAmyCFCk8X9yiLcTxwWkTDIj/H
hWLGoutTOxUfmArkgEfAJHfFyN9IhTZwKPgDObS4V5kHr2w6CgOGElwncvJs
cX3JbiyBGDGd5IZ5JR8XBXBAqzTZ5mvCREolLReEaWUa6HBRYdenAKtUubz4
ZSVU5zai7WOSRB63dhlE3g/MJkMDyro3EWxV5s1aCUq1fJQjqTClMYoTqK11
fMoJq0xe+nUGfe5XIZMqy+Y0zV8cszZi8pi0wu2LtulYvMHHCflKVHf/y0tJ
KiIOAIQoSXhaKgMM6tATr5nKK9GbWIxotBZkZuEYZ3vigGa7yOP5GjiLfFuA
40rnuWw3gL8Rdmlw5/59i7ITLTHjgAHLpKhXVxMK7W+XskotMDh+MeE41Aoy
N/Cv89g1t4OGhbC03OB3QUvttgtvbTaQ6uvfRGVdcwzGHcMR/1xv6rbTIUT5
V2ZwBZASIcQLJXSiYvBfJTKGROvJoDBY+JQ+Sa5QZPeNIHNXwO7loYvmKUj8
EuFRkj/iukaBNbwuxid36bTlfeGGkxJpSeWmEnHu8dw8uNjjj/Jg6XxypLiw
43V57Nm3A8ojjkpYz3yG2QkekUbXsT+E7PMy8t1yNxNUTm9A4EspGPGiN57D
HQQmbXosf+0SL1HeBrza7CFQfdUZ3Lti2w1V++vSgaK9obvCBAag7/bBOvHA
Q2kzEWghs42LOARyvRJikOFi/mN5iZpQo88K0IY9hLSY/79EZgLziTm+Adhs
jZvVEJ5yQ3E3CBJp5LiJm4FwlEGK6ZEXnCVkZbYMpL7UnVtNyPklLuwDEM1q
Hy3pSzMLZWGqPKePLGXVuh52aPn3+/9TS1NMZvHfHACVoGwfXyA9PbeLo/tw
EPYodiI9WTdexsqK+90iV9OY6EsI44y39pwtRVlYgh4rq+w9zD/buac3P29N
T3P6Lr8PC95lM4qOeQBKe3uAocfIwZN1Kias1qfPb8hTQ+Qvqsvn+G5YDmcE
FseN2l0hC5DWYLFD0DPhW4Mt5E7XRBR5fhSfEleXyLVb5NcLJppuulVwU0SJ
bUVCRphh8OG9oFyUYjUfZUratw6NI/ZP7vETGyWTFx1QrzU6II+JC6H21DpP
uWRybgIHNZukrUWOY3SMlFKvpfiGDjMaoa1ETZaaAZu0DZ1P38onwF5RC9dT
rqyQSQkGOkJcGw77vz9iknysbrMkBjJjiTvPT9Xx9fRNYFIdPg5GFYCMnp2y
fDIlVYSR3FegjnDSmCcAJbtDmXqsc6izjCIvEYu/lC6YFRnwjowgemEcA95j
l0mnULUbY/X5ngh/Iqjlh43s1HSb35BpPJoD72IcHxRSwbEjp6Si8YDfCOl0
15gba7RZHKonmiSQF/Nrg3SAMJ8KCnuO9q53JzpJ+YRfHZFKyA7XjmgBta01
R96d6m2XLQx9uxbS2ggsG8d+lfks5xPLx+mxZYl36ujxQg51DOg+WI1Iusx5
V9qRQnUzHWeGAbBczm4jb2Gp62zu7IPfs+DVFg8BMAYuzP5MUPQgG6dr52ky
QATP4EcZJiIm5f3ptnFxjYojFORjfTmOPpN5fTBnVShO9LMhUqwaRAoj+Bhg
yN6JXTGxgFjunJkpLTExSWimuJv5Lvb/gpr74AJJRPBSUQibK39icACrdLeK
x8PNqNcnMcfFYQUCDSKMN8Ua5dhbLTRaKhzuM1u60G/00sHFrJCUsePzG1Hc
PhWARd0YDa1WFae9Qwsw13PMWWV3vX9jaW70no2DJ0YpvX3tPE9UpC2ABOq5
0kIDAS7qKkGrXi+aVXXuEMORdHy5lUA0Jzdi7wap1HmEgbTAxtsiBoI6cGSX
yxiSJb5C01vEUuD1IYYFRLCsWrSyIBQdfQCOu2ZZ7q9JdfpH3qRhCdBFJxFM
BRSSgweIpZBf7N+0G9uRGCgU/hlV11pCS1RwPn4qzl/svnl62h5ZrI+YC9L3
9sacD9ceoSNNqG793FslPz0blZn3vKNJHGYTQJOt6n5rijKVvW7OCPqd4Zta
00Z3xcYmpPlzx42EqNjaYF42wGUlbeNQIWwo556zgK7AZeOWhEB6CEA/69L3
vPbovpAYyWrR0txYeDtj5Ywusw2zPvAUQQT52d2DFEz4HUJYhkBRUil+OkiO
sNg/DhppOIKMgFHt4HVv3YZ8e1R6kWbyB4b3CwzQpjE/9uTcyxLl0GOvAO6/
kq0cgYTgAko17vUAA6Z2h7PNJURHv/1THtgwaH4D8NArxE6SxQFhHF2McXF0
xYG37US8TMTzy4a9vQbzr9o5VFDkbCQEOae5wyaLCPkyB3O0RJPOlnn+MGvf
8To51IYX8liOJb9dojG6MRvKYWexfvhh+wArkXGRzH7r50Njeqe3/mk7pmjP
PUkQck6syl9XoukE6S9FcXVc85rUQBqkfSffzhAuFNlNJ3bq7EoRn/3HIH4c
zUVUoTMnog0lNNMw5zsUZHEFG9f8tA4XlMmlu1eqWeWFijawQcy01p4dZkBS
aTzfbpuJqTps9W5YEHRA4j+dx3Z3oPYv6gwlPKKTpo4T21vjE7Dyli/MGiwQ
fTjXS1J9Q71iFJ/vfaF+Cvn8Y9p9bSoabstd7X1K5vdG1XtdWeZDnQe/eFtl
ZqJwPef4YO/XqpL/+aZrTeP86fwmyHGex6OVjIDp+kz1BWgAzoorzWpTWoO2
0rrDOPt3vg/Rc55vhQUsWePj2c8qMlOxQN1pKbXHchVH0Xz1waVenRxcm7z2
y0+TDUHudZATchYZ8KNAejXA6u2QrfAAknqlj63bSrIIwzMNeTXWgm9xkSTh
sS5gkC5IrRysIghuMjtjp3VNNyt6PMjVBKx3zjvdNdfKa3gI3u7uDO2yiWwh
8WPibbqYeZe+vT03T+dWvpoO7PvLIzOQjhRDQ5Oh3Ks/tV1YtMJaXBeTWiH4
uMhpCqTZzzbnn/vWiKGF+ZqnoKdVLxuugf/wOb36AZHYvUc73UFxDKPWNHNf
DXou7qzOF6L8SEvodPoeWRgkCif2d4rSRSXHTe6LQdPX3g05vA35dXhF8zA9
T5AUJ+0Sqrbj6jS32T1j2uLKRZXRaJhhAphRTMucrNdJ49IPs7/NjksrfJmN
vTqbjAlOOBruCKJTA10JwmjfsKsDfmXH1dnt172kPOj93wUZ1xkSoUqNN8tV
ZYTOuSekg2/R0CLAUTfzWg/Myx1mSOYJRys4qB/Q5Yq4Cq7N7oaoZrF2wIj0
/Cl9wiOmJ+QFrjJATuknIzjAL4w2S5IfUGL47bBPTxpazr8+gPmX5wpB9sO+
7Oao4TpWhzmiKEQpiNf3OLB6Dr/EnWMLn2zC0cin3Tniz+g7COsMTU94JD4d
tYHERmkG+g37GHVKvTcOlEp8HXqRxrmfRPXFScpiX3ImxYyBrEKPfhN8xrOK
zHr72dE5TqH7utGNCUuFB3nsKn8Ps2yN7JpDzti/HIM0OxpD9dOWrgwngYIy
CPtzGDr1WgxB2NZqtreKqyCW4LS5kDLcQrLmfzqHVkGvzKMxk1QIPQoPZKQG
amy6lWhO7cVKtMTg0MK8CKIxPAnyWoVpQOU2eI0xkDQ9MIgsxO2pQLh1bEK5
ln/Rx6l7bFK7oA2GCzBnI/EFNG8YyTRRAHreHiB0VHIAC3c8hBW5sXgH8emx
s56AgeLHcZ92TFL1wlvWv76y8dcvcV1nHf1cH1bYWa3A8etCSI8srtkXsBUM
lE9o2tfySGfhxOVl4xC+VR+OIMJD+urBCdMteXjml41K9NtHDbdTB06YKsEp
bZdlHYuPzGOxxUQgOEcV6tmQoHnQskmEFymkp6sMoSlYSfZ4/T1htfhDMAJB
3DIKW8xUavsn38tbUp3cA4kfXQyAl+MOK2j+uSBPygLo+Du9JKB1OVZ6fPAd
jAp+Pv2UOWsH6g9hBfZmazTuNe1uGUp+2SxldBxylqJr5vkD7jxxDWOv/n7q
Ow4+eR96msytiTs58MhI09W4L/4+umVHfosz6PDEgvKL5dzWv10Gj4mly8dr
FrgNanN/puQuZnKC3Moa/EqoT6S+SDuWVNrDQia0zON1zf3n/+oUqEj2h1Q5
EOEqtjovY9AH7Xs4w0W/rz3P7y99sCWdfknaWpX2BNuZQK7d+OthKbQQHMYa
GfcA2949myvKzgzzGG+275kdC+dx+v55gGN4QEfKCZEclxAcJnnUTRto0+M9
m9+E5mY23F+4hhA3uXg8fA4D6e5KX07q8YIEDprRwHv+0V0ShVoDumSqLl2v
NnBjQwUoRVyKR546uyj1CgmleolK0BOv2t4GOhjvdj5eecirjrz1d1kKPloH
mCmj8HOtgCROvDw7GV8Tb4uuWr0FoCtv7sDgpUXvL9hCBvPEkVMFWofeHatl
xlK9nuRgYnb+EYK4TwPmRpAzlaYl7xUqmmQ2WlZWa8XpVm+MMd1FGtKQMHAQ
nALymoIyVAxUiYlLHR5OVmoPIhlGW5TlAz5NqLVMSRc2efxkGVeXTwYGIYwB
ta2hEzXp7rv96KuaUcezDHcCUZKog3gGRfrEUaz06nGhub5ecOQV+kZFWsLY
/9E7Hnyt2d1CLBu3ih1IiMceZHtUI/kG9YL3vyG0wgLEwlMVtj/LmUMXZAjz
iVdt2x8jIX7dZQTGKh662fUCLVmKHMYaWGV367zheSaSwtzk2r+4jldTb9J/
O6zdrRupo/TakTgB0YkcZi93IenM3JxEMSONshuedj8XtwY5Oiph89IMICc6
yvNDaeC8gcc7hBMEhSxUszYTnX3RXM0MSJR3VA8weuRvEvDqywtBdncu6IIb
tZgPr+fpd+1zWKCAbxoG+d0+8W5ByjsLZndXLX+rSXpeezxTEFuc/JB6CFo5
NUtUwz6K8YqE4cEF/bQAqX9aqqmLpWP9cNNmQTEfFgLY6BCpIPRna+7TORoO
csRz7tdKwahqUkWluO13ULDl+4HJqZPij1iU0eANbK7jV6IIt0YnPB2QzREs
bkdoJQPR8jUvx82ZlCHcWgqHZ8BF1sgofagBawhEb9NyFnJLZdKfN6vxzQnK
2VBl6SHT6FpT6meOk+w2aWfvo1kE0qd7fg0M3/bR1yUOgB4vmf4KANcfRTmP
pVNyC6fdEf7E+aHGKtWemg/wa1InoUm1X7eJwwdgxojEvJr1wJjYk3F3NQdp
bV7bMOijcM0pXbh+GRr1YLK3tywcOcvNaDbOuvjFhJH1pKg+QYGvjNteD9Qw
viFOb2lzOcNGxITRuKCYnhxaEMx+3+rdxNgC5AR3ro/yqFfWReVIHPUpwVwh
54DZK4SdyscpzJ5A7WbBnmIcCRRgTvePgdhly+W6UYi9JH1t7ZHt1tFZG2Pm
CaAnJnuwW+Wuc+fx0O8lvNu7AXct9EUvhh2j5ZtOsYocxtzf6u1aOX3LmYdz
i3OwVmkGSHOYctV6+G4hgf6r2wHSUKORRySyY9kr/+izE1dTeNygWxHevljq
1rkc7rg7O923i0XsuykGtEyqpiN14TVBGA7Ja7SDq9sx+Ww2mbod0pnQEaV7
jHfKOnh5yD/e919SLZucHsJV6/s9tR/bvu9jS2AsZg7SkmC4AkJNaZ8Op6r2
VDBV46/stu0e6YhMfR2UJbh++IOGA59pZ75G+bdBkxrgVidMBkXRloKYexAm
E6IsVd4x3gOlLQ0mF1ZxDsx/mu9yRbrWBQrYJcQJ1OQ8+hj/k+uGealuZ6/J
eLhVFjfULAhinBka0oLguK//PRgGTpk5fOP2fmfFhLVSg0LE4Ee9u++f7pM5
LnzehHb0sYkFyFbtzkuIGC5IOQMoEwEVBEJ/rpwYEgAOhOuf0K+L/EF3OM/r
Kvoy0MZ0PIm2JS6gaIgrwHyUoBkbcl+K1gt5SCdsyclfuk+Ta3EfLSDYcV4r
tVdcV1rszkSIzcCZUT/2Jku7KZanRhWu4yeMw73oHYcc2tKnh74k6j+cKvxo
ml5R1UbuBaL/ClcVqPrF7MOfUPnQZeIm0q/r+Nu39jlbZLQbIWO3BVH52hdO
TYR1LWsEux+DDNCCfq1GlZGtLx7Ptjmph659usU12LbnE491HXd2FCF6eyv+
d+/XPpBZNN4TJntTDzRY2lbZgCA8+12ggR4P1jPq6X9H2JnUkzAYKoi4uKpg
Vm+5RVlfv0rP9NGRc2YxjZ6Zbb8fFBjaQ3zSTjEF2GK7nBo69lZIKfTuhmdB
vt2TTjD+2USsfPbgF5jWDYM8iOnm6qTZrm6uNVyKm10Ac5FZKxOqllK/KKJm
V1tmbVyuvJ+3z+wGrVGOknsGPtSeXFTEl1mmrFYJsVrXkT57IL8uOb+Zy2cz
/g2eRxb5mjL57X9NmLj7bJrC6+xNeF4Gs/IWp3S6UgmEbQCbDY0ILJtX0pvv
Fv3/USQC764aLctXGwKJYyW7sFEPLJg0WNyjdWIBkZfm9IebTFjTu//V2Rzj
0XAOTVcm32NsLHw64RQ+PUpRItyY+6pL2YKn23BsF4K40PlXkWUvEtVdclbJ
sL1f7G1dDfpLBJi5lQ1iBdYNNcZiNUzxWCzfjAsw/cqjCNR7QNvplebloGnl
m/rqjNIv/fWbVSE2hahKe21fjo9hgqG3LBmOJd8qJGEbGsYkTyHu+8E/XoFC
Rjyedkfet27b0H2i2NcVwWaOMoov0sfOBFpVtYFSy+P6Nau0gDLIhyRym6C+
kf2NUygWyCVOhx3vDhFLn4Op6j/4r1SrEr2AXwsnKR//gJQYZLPX2IAbqHeM
PWGA10Z3LeIGoqstgEkYiWVpIKvQYA/bOHMxA0nXi/DM/31nlr3sGoY/4U21
X03QScrb9G6PFB6wsN2u2AnFj+9kozFIKy1mvde5jzg4PX+E6qiRscQJoRGX
TmKp36UBQchbSXPcl+fN9JPH5pD4Nw8IJpvJ3iGD8zK3FN4K2NdQ9LfSsIuL
LTKmuHPP+ggC7PeISzwhQJM0nozR1o8TbnX45CaK+KYvK/dfVVejRs6OIWS3
ry/0gWgATXg7TrSXjexin46+arSjivsca2nNE9Z2pQ+HrfD8DVlpTOBEkje+
ov4upcGVR3VgtYknJsl+bJTChFuNtMf/ZTQXHF51TEGYAUzIuENedyKY/j3e
mvdWWfzxaMmV5n2cUEmr/OKlUEi3m0H33P2E9AsLjLoSW6STeJaR3/Ay/3Ck
8jXfi9x9NVCWobCIOeE9tHpCGqa+lFpiCWUoyU6LV7YaCrWYiGxEzkkRUIJ5
WMIZxMZ5EOcO5fLlgVUhi7wEsuktvFpPSi8+iR5bfy89YRqjUSFwxC4CL6Hf
hJoqn+g28YZMXLXSq7hF7wuPTqABrNx7ajL7LN621nORUHpB/oxs22E74ol4
UxR8CJNE1ByXypTIJd0Vquutaf5LL1jxYpHgspVYgcuNwZiKYLjP9Psg7f8b
7UMfASV5drAb2Mc0JEk1NdrTgCJ5lXEOq0V07gBNXJdDipegh86eQomPwghl
xhUuIqoF4/95nUg//KZAJgtZ4S4YTjXKDogqpU+lTQ2CbQ22pggjtAnze7as
84MC2cEAgtJ1vfSJssltH4uJLJDEcm32CgEnmGuTVADd9xAFxP3kESuutZT3
svmnipLKTniijCP3piJKGDJPgmXMWh0KY1qJpbyomTzU50dtzlClbhiJrhf+
DvTf+LPK1yCL2HSgT//NU66kGThHoSTpneFZGwRL8uqyTKuyn02Y9K7pHMCT
vtsU/9vi291AMoi7JzjWmTbY/ne/J8n39My/xfUATE5QUzQp028Adot20vwV
pwgUbLhx87hD+xbomleqR/1HTfGJvhqaoJQkiFKB4ie6mEW56DRpQb7Gc9OV
SKmdmpncfRmT0+/vwrCs41RSaJF+Xc+cuyqONp3z9o6cnbUtbFDNwpaoy+1w
iddmfuNNSLQugkOGnlYm/bJZa9qH/BXzeLEJZswgkVpS4RK+nR59cGnDDRSK
nvlRaqIgfguFMcFbPjecZ1Ep9oUBktpyWBxu0XBAsh+kMaOcxPFEHqE2hq9o
lBaeT6REhXNsd6Ogiabxj4OXNIBhoCTIXWFqaMjVWtweIxWwyIL185T2O+kH
zW2Az3syO6v6m/Z0rBvXlY9dJk0tmOyt8qhUCwoizPefg6DIK+WOwd2+z+8C
TJRwJfBYUDhyeO1/RMryBc/KnIzby1aPSD+oZyFpF0aMmOXM9L4vxKt3pG8J
CRWvt0v1uDeFVu49yfwsQ87J0v8u6spUtm2J9ZmrTz/PXsac+dVpQJ+YVh+N
8obd4XqH8tlxAaFJHRzMabmU79HbiBALthu/vIkxNi5JoTQEVAAlS5bvcafA
oyiKHTEmaHCvdd53eSJuu/FbC/3IJoMRudXr7GrxRk3/45OEDYiAoTVXDcAy
kiNFN8kh/3zNyvnAOfJM48Zz2Yg+QJNciTHUMDFVtM6dMTe0BJoPxEk455VK
/GzoYgRXRa5yhtx57yHvpMMpNRa7CFNSt5o6QWotHXx4pzARpGdNngdAcPc6
6UtZjyDtyz9zL0e1gZ+K/fU2K0Xj863uSrbVQdlpdKBeU3EoSdMCVHtd+IUV
UTPKwm2M5sKZr+i7ivLXzNJiMiixRipfV2QxJ6fU77hzSiO0bHeEOic44l7T
tDupBQMKa2SIPVMXzI7TORYOE2jrTiQC0yTUiPO4KRv2Ux4pyEDHG3IfOEHr
hKoRKD4uJEnHWIJzdE4mB4McEM7Uy8S0YpIh1WI6Na4Bm3FuyyqJORt1BKen
IHWKVpM3Hhj9Yc9h02btfIzBT0gtnFL4EdqEe+dox5Efciid1griKuRmqjJR
6U8fRdTN21uCuaIau2q7KhOk5vGxdwiF7VDdtloTnlXS62ihJuXLeaUpGvxs
w64jY5MPiqbf6auJQGQtuMeDop0R5TcWQ3ND0UYb4tlr/NXanUiNsyFVZcW3
i7tS8E7bySmxZAx/N02IziTyXgJphYk9f8PYlmCrQoo9ClFy8XFc3fROJpaC
UBRndWyoNw70CouPGHA1iVsZefxSbseBiXNBtnuMTZCIZP/WlaUUu+oKs9t+
QlY/N/YQ+s2CzQs93maIMlyXDRICK2o0ETxuufZBIRQVwjpAgLzE8MlxdbJZ
918+sQk9ewEipD6u2VH2XDHX1G6n3iiaHjHncu+MT5nfaFfzUOwoQDvMRL5U
KNNqGshbLx5GTZBFMeR/xAVzRfTMlkDcYkFL3Hr6bpnLc8nyLlKWyqe0KUXr
hk/rXJEn0eJaivaAmH8QuUKJT8ImwIaKKD6Z1gn3dSf7ohFg02cbV/z33Gyt
tDco5jn+GpWzqlhZnDfT8D0pyTXjH29a5Hx1PqoD7YWBwCC5YCdo2EqxkInx
cR4jmqHDKFNxaVM7sQJ4TA+hN/Bi9FMpJb0ZG3lJDoYe6u0ppSJ+f1mEsvy9
3DYH0U6RYV5H7h8p1iHbtydRXp4oce3SutCsCgWT8dNHO3kFqwxtzVA+3idc
5753J02B+VeCgmtcaviRGqajuvrqGVFDqHxa2vVwa8Lnq26EOh71K+AFHzSE
DTbAxQ60DOTfba1zX1Bju2UL7Rk5lZCHacrEfkkiqn4Rzgrl5iBouXCY4iko
/CIX485Q0yHaNOAA819z0fVEQGgZYpmpr4BF5siBWVLJm/vszuA8IfVzYMcz
0W0N15aHtKN00Mab+dYZYwf7MDUDNLbzRUZ9+uaf1yRCdXA0Y+Ah48z5phsp
rr39LnKENEFOwnHBuz5EEy3dMq9AZXLIPXqgqYvwV0MNNMM52ClRVrC6GE0b
cX6c15Sbj/BW1sUYnp5nGMgx1fNiAu/5rqybaXu/YNZaanO+3bsgi168cUpq
D273DpZyAr78sx73c/CV1NO3GZNhoUmyGYc+IIxkHooz3YSOKEbK11crE5Ul
RznWrThBRMYnPFfQWC5vAjiXb5+Q6qrYMbBiOL2j2lE3VzQN2fODHFg6A1bU
s4Jyc+CR4e6tZXpOvjZ/AJLigP6si9WTQZaZFq/OvLvSEvlVYlRQH6JGWZsF
TLyESMnFeAROFV/PeqzZ/lmLuJUjYvphmqkQgFQ7oi3+Kc2XJgkbg7cH2og1
bPdhuMdFaAzA9dj2XFQ10la5ivsnR+nfRjzFK3umEUtdk2L1XqHwGJclN89H
PScmOoC6jGL+ge0BWNaVja4ZAwZm0ptu/EiFx4PthrmVmUUiYE2JI6Dsnxp0
jYiLYByg8/i0KWvWl1Si+9QZYRspARjeiF/KJNSY5AQcMo612YW3QVdrziNX
gmPjQ4dlKASNylOgoy6Mwg34Ldcw2kSHsiXDbWqLXQxbli8iLVy4fbwBsP+k
keaBYUUiEjlDfSUN6Ru1ffcWc6UJEL+8fsLhNGI144x1TcyxA8hderOZw8Kw
k8cGz60BlT1rw5fLbDFkk1ASp5vRHhC1Gs+DgSi4NExYWu34FoGXFKyJMngg
kESl4jbUIk/oZu1djn5Z5G8BwTo3K38IvYkFm7ZK53ORa/KVq57zVryocof/
ViU92PaRqXQcrLDMMoIxSyGvDyiMSpG4Jb/6EeWFZOLpnq3r4gKePq28fz6S
Zg7aJYCWvyM+oKRoUx9akwZ7L6UrC8Rw563I45dkXmZiXlDHrO4ctbGtcZMS
/wHcP6DYBBQ4KMAuEXvNWNZZUOm0Pn7ZqXA6sAvWncDsFHFiCyFwgeHsdiDL
nUBfy6X9jBeqXzy67oho8qmlBtkJSiSYdJKC5h9y4In9gWSzIAzuQxvRKMaT
p6dWFVWUzlJ3Ryk7asCHs5W3NBBNbpgfRHyE7CUkYJ6aDb/2OCCMNv0p/S+j
Jby7a4R7G2kvGbonSRpLYSUnM6OYd/W4p79bs/iJFtW95tDNwMWQXnF2O8f6
DXkDLWJuOeuf5VOEUY+nnLP0KYTfiRr1xmKj0uM9N9vyXluBJGgIs817VlSx
84F8BV4wom5dVVL1bM5b6khSCgjhVFMo+lw27sexvOgvRj18fevtktjihtbX
lzAbTeVXRdqjQto/Em9rpy3BusX9eyuRfWotWd5C6Nh+IX5CZTWPdjAvg7P8
5nEu11YZj1kbC83OsZZ9lfBNh3LOL30gQcykeoUC4uyfY2d3m1MTDvzhHjG5
RcGn/rtm8zXLvlFkwGxuM3vdontahqqgk6YX2lFIgX8KltSpRCuVRLR+gwGZ
OTmaE3cbGrCEw0k14JPRmi0Q/vvK1neSIJDg3RDMuoLy5bAMkgRikxeIb7ST
h39L4n51+xijM6SdHxSNEJn+oj/GkJCGJ6p3h6I1PmTQrJfGHVQpFihIZF4+
wvtBQ0pizgMIqHMIEm4r7SaDzIbITF4F98sJ1CjeEgKQH0cAPlQVuAgAbwuS
YE6eQ5Eoyc5y5FeiXtOeyMX3+Urv0PggjdUMDI2iROKjJhDAt1S/KMVmvcb5
P9MU7bDDBndDmREYIBrLiLx2iHmJmpWZ3wTb4F3J9DoIuJLhJ7vVV1PP+Rb9
DyDgBFsr0zPUNhnwHcwUQ+j5R+VQCWPWzL+RYjL2joZWIoqohAEXpKSo4SR1
TaiKQDZF01cZgJC/7qP6cjtW9SkQiPXoKvGlp16Sz5/Zb5u8WBxTmfq/SW3V
zt0OcsOSGEGM0UByJ+xbN0s19TVaNgUQRWXiArbIxNHv1ELijbZN6JBkkrTq
tCb2g7TWL9rh73Pzq/U300bbzNHJOBEDZhBjGoxRqe1Judt2QFFxYEOG/Fif
v9eayoO0ljmJMIS2idoLthoOVWeHHjZyPT+Ikh1UQhkdRUvdlSDTInKbK5CM
ZFwjYuYkYUIHsw1fOCXgze8nC+7boPJvlD5woM5VjYta/sgMikuScVLKXzPH
iEAvUKRTjh69RaWa1yZbKmbb6odtLh+rGjyfl4OE4FrekFxDrSt+PpP7Oo55
8nwDweozvhmm2VZES5s/WuYeIRWBUE8L9ITOUpFhrCBKLHJr/37u8g3aRz3+
dggGZ5V5hUQ9eVKddh97Hdv2q5n/VVN4phjtUMeeROcnfo5He58vVDEUfLXe
3ObvM/D5paMmnYXbHgfzUH03VrOQZN1bKR8Me2/KvcSuyXdTYTTVqQzvriDZ
5zAaKcj5Qu2UMxiQqAuulXK5rRLdPyQIhLta+p0Y/DhnRydeNyeJ/6ghAqYU
CF2BPOOeVGzEx34PxI/9ZzNmpDDHypHZczloCz8z42cM8aon0OvA46x+vF8E
bMvNQROtTuJxiTJTiXyJ+5vbRMISLe/1knWOQGU15XAW0NpV4nFHQZThycKf
gngWl8ld1VdqnUvuj0jFjkYYvuMnVwTw+n7fyieBLvb5e7vTLbArRun6UUoK
P7zhCauD5Irtw3ibkypdpJqsHWJNPfoNZXnM2UQrTDamduCXkwqMjLS6kCMe
U1+xxIbZdVlbao9wy0K/nvLY1lisE1mzHKdtAm1IVgpUboBOyo1KfAUaMIwz
Bigc6gN0zNB9rj6NHHu+X1OuyFhaqQ12J/68WoeySlg2nqH43nDWWbfNxCN8
MMBeYqRGs9ubmLjW2LclseYvD+ilQFrjdx9kyFT1zrFwSWFMC24Woa2CJDP2
1ytu4sQ9F2EpnM9hqa8tMMPI6dzfXxOEVS3KDR75qfM0ukaOFdLzWI+X6wnd
bAkU33U9e3EKWKjSSWp+Xx5RRxzOx0ciZiXT3t0ZufO3X1QJndXyaVV8EZls
x5F8CBpqKl71CZOVUm8j2ISlvT6zkMjPOJqebtnrdtFOBEn+Lo1jCLsgrZLA
G7Kn9wtxbFQfGpOYBYxdIw7CihkOhSDSgu7CzfWh0mDgei8Lxe3UM9fk8vcB
Ts+S0YFts0bi0Yk9TEPuXp2n2Gsx1DF6OIOas3bfgvhF87bx7qvUtwHi+GEJ
KPdhfB706x5m9e1hwaAfdQ+uqmZ9WcIxrIGPQMpqyiPljdB7iW3sdPguTeNC
KtdF2ghKKAOtkcnDfs00D7C9h66sK4TlF+ckmCekKXmttXtweqQ1mKYrNI0o
u71w6NEKZnI9vfAAc/9c6L2eHv6ugsfD35NTsLhzHpyDyDEgorF0uiYJlWZ+
ggCb3/3XpD3JlMbcNDf6bI94jSp/HHmCVGvHqW53BeIfLhILUu9ODy6am5Gf
dm4py6lpVeuKdgjVq2sdHEtBReepm2uPAbpD6G3g7SShG2Wf/qBvVN/tN0Eg
cQ9ixNvnzif5xM6S3gTjUFSDiUU+GjB5qjOyjQb++V4ExwM6wpJKW2Clnq96
6JJ+hrb40kOVP2igAimRbEUPZMUXfs6Ns/8Ht4RTOWsQsgvQEE6uMv8jTxVu
EMqU1tL1EameGY2Xp1sGdLmYJNGQeGTPBv9HVUDCGlGcyllHnI5Fq+buaezU
vDfwDlWBo64QesB07yRSoBEKCn8EYtIiphIbX8KZ/sH+RrmG3aDYZKoB5cQ5
27DdgZFOGyl1dtCooXha0ZlIdraZvRAjglwgCBzLxzAOT+SJQ8u5GJuZdgiv
A5axN0h4HiOordi5HKaqiUwjkEkj4ItykYpkhXGE8I2Catxz0LzXck4n2SMN
kfVVWm14VwXktqcB7NUhkd1og16hYp5OuW+7QK1TnORTzasAL4GQq0q0712H
+a2rlbURoDx2kImHRv/IIIrvh2Dg4IyvxEJscRgZODrb/nJkCiw0tsK/2Kj8
wKbV569qEBgsh25wpSwHJtRmjdD41LyqO0tzjRbfD9nOsOyRyf3A/MbogJs/
8350JjpN152zjUEwTJBSucfBJEKJutzo4VhnHg9sDEyM4BXvDl7t5VCQxCYC
3YvvpDwCJFI2uzJ6KZBCs0CQ+bxn+h4RB/StInGjZJLj7vxtxsTy9hvTBLMI
ZHviySY9GRUGr+dKVN7yxswYjaSWHAoKNaquavfwl+QOVj3+B2IWqrQtSJBg
7mlCeggoKHM78K3wlzTR7nQMj7bJUGto1qrVBaH18FfeDNbkMXNsrip78ecT
os1w8QgwHtZWpi5i0x9DReYJzxE/URXlUekOqI5K+btPmKOE76pevSDNPapg
HFTErWJ3qESlQiPxrRvo8/56r/Twj8bCUd6czotgIjU81FThs+1958F34xiS
LqbL7M3m0iYZ/amBfR73Pe9EAefElAOksxFcXzGH/OFu/3qKHbvgPTdPrw1y
pyAc+phnZPHaO1ihqe0h45XhsDt0vwarzm31BGVR+aUk804+yDMqII8F/K/O
57nqO6Bz5Npvj51EgtKfdyO34LLiF795RQB7tmEC+tfjRNXTsAERw7Ep3tJX
VLRdwUE17ewYbvsD169ODMZ3wlI6/DP5stJQt+R3Di1scgy6YKg4AnsKUYlH
Ipd7kH8m5N22RDtqRjVCxknVCVNbCFzyuWCpOXyqJ4BxjSAIVj4UbXmfCRYP
/YF1RrR2ps7JdThSf1vXey2PkvLXHKhxTcVorgnPfpnM7fC8eaENkUcrtJm1
mZmBl6u7kJw8DTA2MRBsVUMY+OdRNDNosUN4WT16MaPy2U4J4IECqt+xC/wh
+UJZbnYtJ2OyPqtJWDCat1IS0F+ZsA3vGgr2q6+USFDGOZcazLsFdkrjXAaK
ThAdMH+B+zslWpkJyLrisDHlZDM0sJGTXV3DQYQ/2+74Kfrv6uySpCVwRbG9
7xfzOZzTbMnj8fUrkn+H0tkuKm0Ts97tXBX6X5WyU5SpvtTik6rqc+ywr5ne
gvqSMqWRXygAKbBxhtkpDjmR1ft+RhA2+MMmTo+83dOe27U7QmF1bp1sMube
emu0WEOnzudkn0M7yPXR+bCnb/I2SZFJ3wCMnnMvM+ydPvKbdy5qCcr8Eie9
hhMxa5PAEojm0Q2PI1fPubhp7GdTTJqoKKctC7B6/1MrgRkXEwRY+Jjxibqb
a2XEbuw0GNt9oYIuaCXak4r9pofJ0AOlR66BU7CtbKQng+udPmHNy9JOPqdo
BfFz64GdolFS7PvO9qsSiD1CzQEcWf9PTOTjlNBrz7dwLmxf21CmTT8bjBkS
5b+Pc7o7mX8jF3NyVa0fdp6AG5IjoU665B1jAkyLSroPJOQw7N8lpODhPgkw
BbBWTxChxwhwkaqy1w6WCiyZFOLYdpxHguUK5Px9FKPHbXnf945o3Rk3Njlc
Jg/YJbuUsrltovXWwwFo2slsWaDWxtDiwOxE+oKShGvxWOZZbghogXgBp4Iz
HZIEIkK8IRtc5zonijUZaR5pWIeLD6J1HKv/DUhL3l35bmx+T3I0B5UxvU+Q
x6PBTBK96u7IDxK/Rb0fgWZLcyNkNjoXL8Vvg42aBhDJ5HnTaNzRZbg8Kl2d
CMT4p+EQTMCmlc435PmrtU2tXB9xZpqTSpFT6PFjrSo/qzPB0mWlNfnMNBQk
6jT9wT6gtJCpz0vycEGf/XeF+hyBxJb04FnoWQm70eudRjzdM4vYMwY4ENS7
YQbM1t/KPXdO7m1gc91UMr5QVUzlMDgrI3B2zoP0j0NonK9tcdDWf+Gn9sbO
fT/2nJjt/sHz9d8HdZTsj1f5BTrDQc8kNP1X//lY46fDyTH2YdFu8bRbT8wG
e/5YI4sEybQo+uzaaF745/tOCu2LGTa3C3/4rp10JYfxwq5UPvjaMtz1aTjJ
xs8bK+jDBK8mG2348FqG8TnzOvGbaDVQwWEcci8ad8xmK5+bfcgNNs7TRR+e
mdCOpwkEnDSkST646eQxJRV4DywgmrydCJd3aJDcXkuyQJt4HaBZZ97yOk8U
QhrWxfFTdZLB9RSdxGpYV/UXUQObRDBvo9Ks5R3uxG12/bulZiLfQ/NrcXbP
Je/VNozm4SK/MC3GHrUoEZfN7tRcekoF1tFcLctgiVJ6men0A+ZlMRARg1dg
cHe9/gIFKy9uzmGQHQkH1B+h3kSyDyywNQ2Z6H7gOg9el5HxzUAcULjIdjxr
sThtQvF5ngqp+/X+ef6LJ8NyODJ2NbfclQiy1qXbMSB4zDj9DfcZif2MWUou
AHlbpbEAEpSwQZ1EcTCB/xazJeav1yadzMvoIOoiaN13+gfW8iRBSK7fE7jA
+PCDeajWTu4s1sF7HGB1d/0AX2P0lHBfXoXfTHpEgd0P2yHrdmMiAoaseloX
zr2jeUo6a/9JHi7wHlq1ysLEdvZRvLzUCW8zh9fv1xG1wgwUsSSGjlOklI17
BmH3g4aS1FXTJXczmGpaV8uZtgoJoWJRFCvUVATiw6L8TuT3T1PqA8cHga0u
hPHm14sLJxpGix2uJ4t43Q6RxCmdOgUca5YTNzmgJuw3/Jil4Hl2cWQOZEH4
ykOIe/kB4C4qNl6mLlJafk+jTlWoHhLlx+I20MHs6zXNc3urppsvn56n1VKh
dDWGogVa7LF2n1H0IrCT6cns114zQsC6M6+79Z0hpKh1e+8wcyhXEW5pCVEx
RrYPqfsYe32hk9UgW6vditP6pbIVWivzdnbFsqdEPrBeALupJqr3jadUvOat
CwmToDQnq8RfE+We0Pi7Cd/31P7M7xJ+cymCizA/6S6rI8ZCnRPwUIUr9O/3
3BF+UZogBTXGM0MypmVBiTbFmcLTlknBMOMDSc1Zk9PcsRSH+mHkUYkUPW4w
NP4Y2KE8Lw2Vj5MOKbNLeIwRRzcUppFC8FKqUThKFX+/1YAt5YWU+Y5OtP30
aMJmqDaHJK9PJqU58K0JSJJJue/Vad/V7PnMIx0xfFclha1fCyXTRRo8SIcV
w00Fb56V+rub5zXLJUZ7qsDZ34LtCSrzniCIdZyq6Zf5XDuV9EsJMJ95w975
3oEbN5ZQLzEoMBlMxl3q1pZulDSrT5j9sgnUEcPZKaify7HCY3IhBKhJKWhZ
Z3Y8OxpDIwhuoqxHTTSQoCOCxOs7tCBHqwoFyCO8E+LmvPYdhoQ3wMZPEXjN
sax+46VhZQ1phkonWRjfo1xqRTQghlTgngTTinAGN2qE1x7FOS4xFuBP7rQs
u/D6W66u4ZkCMYJRUxeDOHkuv048i65yiGP7U8LLv9HCNjw+CzraAj/FbMsW
qj+djJ6zSJjbDoVV1pml3O3H8liz4D3YCvmMt1CngtL+M8EE5qXsOM2Mv4PS
ZctxKvhbw10B8YGKdq+Q/LvVWfhWEqqONPgeuXHAyBl68tsCXyB8p7DKJOZ6
SAQ83F9tYbn1XLAtQq702DE5DaPZSuEzFR8gloVUqRdkSLjAJBTch+9OtUqo
E4GtwSpFnt2J9EgdwEcaGx9m/99ZmIpA+VheoiBgLS4pWAOsZ6cgTwTzpWWh
W3qzKiYUmSqRS2xbESNxdalXi8NtX9cfVn+Q8SwYqqi+jSstI6UyOWvtAGKD
7fLJPTTVbs5oLRVSo0bwPJ2HgrPeoLr8X7XgUM9vRvNe+EEfrHU7Ooae3osY
xqxD/Ydvs9qX/TGdlerYYT59v8LqkAEXynP4wSvFHFe9qilmV+YvFHRsVmbp
clCyNIrffNkO1YWmBlWrx16x/ox8BvNNgKoL8KWHHVeT5+384aelbVkecKA+
o5Ri81AAIUH0i+f3RQ8L4TLsRiwvP1Q6FEN7HcLYfuj1mCBD5PMNfhxr3yu5
3+Ic/iCRJeKwYSxw1vaRXr5fX1Syd1QXiwXXyBW4+/i+SorY+H/a4yuA8ff1
n3oN2kmkwW4QC4g0WH56YW45qbDcbLLiMk3riaGOoIpqW0VHfz0idU9rBMXZ
V2J7sBIWPo5JMjyAzXOFfBEvbQ6uZXjLkDxlURX/6kjV98vHJlHQiRDkikux
RbmF8N4gC8Zbd4Wib6KSND28OdSgmlSX7di6Kjw171L7mbR02xFVA7YWvo1M
uPnP/XDycyLUnWmnAEEwgk3NvzlC3/sn20LwsJYH43R3172AWVW55SIt8t09
/xBCgi/jVHLlCh6SEBI+xe3nzEjQvrLt2rvMOhrT5Kqn4lYWqvtv7ZOapUPz
aPnohTRte6/Mi8baUjfchCPfzMJjSJiP9hKCqQ8lazLG8j+edQMeqQd67/eP
c4eJXf+/HGzOvRGy1iSHlJOvBBRTa+BnAoFUoCjYycCvfv91mvG6atgkL2TP
KnpvHuQjFdylM/LKoOXbEEpk0x41pGm/89jABiQrRdZxlaIURhmfZP4cCKh5
GacRM+UK9OKzcXxoj4JcdeUjrrl0+uGWpEunFjnVPuhac7CIy1ZuIessJxQE
653pVOn1omkKkoTFOXuDKHBLICCzBVBX78dLQXxv19n/wRQcuCRQmex6O+q7
SQtCeSzZ8cSlq3rnoqha/IAXxAseOdP9PL0leFPLwVV5C+C7KCxPyGtEUNce
lVOAOpEwXUq0r1aSESiAUOoaGwrItW/sbrLxFc+NCuK3iCYDy0VqlKuWtNO+
QgmkZyTEBuDrrXDCSFqXRLAUNZYZdYpdTvITa13bl8UjeBezXtT8pPG11gJV
DaQjL+25NGge1ypWj8GWhUsmz82ov5yrZLYuHszaStWx8Lz4hzDn+xyMYcVK
t0QXMuTuikF2MbuWgXc69y/R0aAWny3J/NdcU49dq/H2zdXZ7SvuGNHXyaYi
UbAMvPgCfRcMq1m95BrcNZTqwj00xv3U+7K9R8EDqw9KvLubeExTQYqY4HpZ
EirK60NqJgnvt7FvprMbXWBOymKLwkR8pJiLw/z9/ns2OdcjEHAYK9BNWqH/
HIlfrTNfigZ83CHwgbwYdPMfkI4XDwP7YZ25ZBk1MtOiXFN6UhSYyq1JVFIT
DICaeTJuUaAY7TsXLEkvjMok4Gegm9kKndKFFXYYNxA8Xp1q1FWe5A47Knwy
N1cz2tjkQcVV/AjKS2KlzuOhMIUp7vb5T9GZqyZOZwA1kmfjMIisw4Rb0ZfR
H5Hjtwilpu5JLxJRbB8Xu9t0WpXF06W/FKNIOKu2bH9NucNzXG1ccKUcufVv
NFMhayj1+KsSAhNMGYiHpDXjifGKqv5ec6X5STv/pUvUhgBPmzLNPrS+kleE
/A8kO41kezzEE5pGc5PY/HKBNp+cxT7mW25GUL8UaOzQrrx4DCMvj3C2rH6y
U3HT84Wa8AVfIBaF0gcCLlHhHi8tHekbfPwVFboYryndBeJHedEZ3A91mFfi
mmiHdJYqC5V/NNqRIMiYVYphYN5xcb8OAxHaWXsjJxhZDK1vNM52yGXen0ps
+QZvxxNx7a5BuPFnpZNtOmdwuwrWCO8FlYCS1CquyKZ/16Zt7Rs616X8SIhj
6cpPTJmsJsaRyDca2daVz8x6J8w+xW34LW7EeDgYQJzv9adVsz2fVRJYHpPf
gx7GiCOgYe0VqHZxKLZuV/87kncm1Rs5KwkqyoXXfxPC1PSt0HyX3G2IxU12
CthQ8FdEFCA+k7kdGcKhPstnPMmwjCvMNyhrpDFK2EsAt56HQw3VJVWMDusV
pZNJl8Gzr7m/FdkA6hPdKnlLuyIDn/RH5VXTg9X30BguqbUbKKnbLjTlI0rg
OZB+OZVV8MhEtZK3GvWGv3NYwKIzAHS1TB+ks0gz2pzJqYf9frAU9oktAFZl
ISN623zwNJ4s60db/L6aEVYlbkc+NVMhJ1wBAQCUgJLrhSqgpQlRMEC53cQG
iGw9sWe9U1gX2OBAOQEz2PwA75s288NbfQ66H67f3HiO+eHplhbcoVbpqT30
dRwHIwzo+FeW2cMd2Eyh6GFNHkKHTJe7RnfxCW3jN5OlXxHE9MOKZSxsHRrA
ZERNPcD4lGbm1hCYZ/9G4UVvG/1Jb07c/MCOQ+CieAD4xQ9QDaZWGIIeFdyY
onmW0yimbDbr5NOG5wFD+pyhAQIADc5NIfhBPhabkxpX4Qm6F9qqZBvfI7UI
VpDa/FdbsIgVyFNv+3Ix4JEfR6IdSQE26QnWZwtlfoMfReLWNYTcjUT2oKlY
DW0NW+tQcaM48pbVoaNYJvPQW/MTLJ6Bd5ti/B+MLkae8l+9C7+Hl7LDwq+G
FkDDbfJbP55dADbt+QRdoRj6XkWUhXM2z0U/vWnMnrqzKKDbQX1PVkPmSS6z
yDXdtx0yTbMjDt1AwKqcFwP35oS54XPvNlrF8rdcSmw9Q+ktCno8mcv+gwaM
tdRZUZtXJDDXXpYh0acr0ciliOwOBJAGRFpyvoH/cymdsCcv+GqG30pkj9vr
Xa2rTbnStJJ1HldNWcnpQOxh219NrhK4gXFsyvQwFY+JlmhbIQmEkdfXTJOp
79N0Q/hh7dtf0x1izrXa9lXeWoK1VAUMVmENl/5DG2wb0YOQ9yxgdaruxaT4
iwGhdzqNV28se3TZB0AYBM6NM0MhEWReGvZvEnN97emGr+uUmEgF/DLXcnSn
n9Sybe7RuDj4osT/h65ZqC2DEIAcokfMVqe20xU/I+3F/y1h/lYvkVPgPvLC
hAiFz7G7XRsiKXvworDekzcbwfFnvGzsVCCcJ2QSi2YvEngMm4jD4zOYWm4p
S/O3gYOLWNLfJC7aPwlCRnmpPmpZLkzgCczp0TDdnBP5+e1NoK9DZtxEOFKK
kz4RNweAG09zljgbg9Qye3Pe3H+YqgA4dPyyEWhOMIBegQxcYuZrF5bhQ6bB
FRBvzpDSo+qD/FEr0rzGnimz5R8vI9gQXGWMXio+lPFPkj3+XDKdJMNb4Ocp
56D0lkFfhtNgXHyEzL1pnMiZeMbNOe5UZ4fBWJ7S9Z5vbX1BDaOETDWQltUs
S8RVRJQR2bH85221R0S0i67gLjstUe9TvoRRWj7hxI3cWeVB0wwoLE+GzLeq
DrDGbPNgnFPgQz7z43zrwoaf2Wepr+uJ/q8gbaIPVGCgisbJzZrZkdNKTxo0
AQZTE8z1Ft8NbBjFo8rt1oneWoh32je8FKsfwxmJd2QE+RWuwGzER7bUIXBA
m62RlMITPV8FKwa1H0RPW0RctPSmmUMaCMxehdW7432xfO2I7vZFofhCynOV
2NPv1sBxaZZJV68Uwv4H4qS5g8rzcRiMV764jiIj97LCYpzXoe/VOBDZUgai
xLTw2lwHV8zWue9eRaIsL2jpFLkW9N4L+rSsqm4BmiBZLN6hKnS3SufVx3J2
eOLYmCDFompWLqKZQOQcX1JfCN7nCEt0hs24CW+NVLO1TyYuh/uU692Dn6nC
iopu+WQVPc/Ha6ojRIlzDl6+LXNaYj5LURvzdo55el3BLbZB7WnUku4eOgkl
2IMjEhxv1yA13GqnAWuE+UG8WqlVch9Eaed2ge7/kx772GQPXqbVpNoa5Vxj
GZSgHXQjifz1xOIDfikW2XkJBagcuwQKzt7jJ5EUVeq+R4/q3cXaEkBSSF1Z
bOVVcfFb3aFHt7HNH8LXQxExP+R93Phd0WzXbfHH2fdHDz425RQpEo37pc57
TisqiA4tOt4g7YVccysftmGSoyXIjGdpk95FktCJH8N+vC5QboUvqGOISssA
sIL/h2+A9BdvQrxmMtHG4aXq3X87hiKic81MpDDJ+DMfXMjkGHMa7YBFJu04
sfAXc9q0qIVWMXf2bggvj1BUIashXNVfjD0OPR6mrJNR/q9dx5ymsQ+z2FWi
pVMT1qJtk+rBrd3ZtwXN9PeYbRrRubGBac9VPcvqs2nzzdUVv9OOiM/cuFpG
K8V0+XaKNvAhwkXA2SQ4pkW6X1XQVeIrM0IO74TXW0b2RXnnH6W6+LWF3yX2
pJYW4CpzLBxBBw+c/MgM61hslsN709xojXSLNK+pYiHrvQIKxZfWY08sNt6N
73OP7Xn9cY+TNfPjE+wJUskcwOAVzrRDQ2MT9ohDZLdDh8VWJ2WfH98rzVVF
f9sBh+ALR96XBhWLA2FchgwnJ/rgbHQyBCXmiTjQJJmV7h8/WVg2hpAvl1XK
jzCn+Sb0J3fdhSLQJOc5RZ7iQFcsrT3nKA6+PSwAxP8e0UEQxNsnGuel4kmB
g9Q16/5iUGDkoBZ0CluS3oZSl3yU5Hltm6pk+Ug28ZIebC59LC3IM8pu3hTJ
ecAaR2rILE6y+y/YKnGwJV5AVklueO12ELrdnS1DHV7wy6o2qyqoF7z3VWlO
bwA2QWKrEWPCtN/yqrB1RaNC8lOzycvTtv+howkDACLeRZA4uPCr7tzZDLNG
5jvvdksBLq+IP6SpIP3Rd4g6JFUqtDymKoE1vJuV5qq7D1uQDiU9w1qQxnuu
BZWWsiURbEutveEU0RHwRlUyZIRreDkJgb4Ra7CN77NeoHq0Bzqc2M1ZLEjJ
hRxmLw2uC6Gmiq3O7bQehVNEMSVe9+2ksPbkkrp7S7BE1qFsOV8652W1mvMd
W2mrDd6XBJ0wOiJ0lJoau7aLD37So3CNU6tg8PhVWN9G/FdYpLmtwxyOrHtQ
jakMuqGaOZEPfyeQ9aVAoQk2VZV3FWZ6JfCuPJWqgOVQbW2O60Un/KO3ieAd
IiOA5z23n7i5FIuWBwYqR6Sgx4/g8oTtGldbOEfYowdfviFydogNpeVAybik
tfgNaS5nI/191ZcdotroNUiFbJa0ZUPXDBqxzn8HV82KhPKO00P7HXaXkpT9
o3Bu/ySITC2CV6gs9wqPPQKXvcL3FinX/iY5LQNwhLsoGUp9wiwP/Edc999d
CIUXQJRRb3Mr24VcmY5tbKaDuPYhTEZF8CLoVAlorEXWsovGiBDnSQMryV1m
hydfIrXib5TlFdigrGfXvBvz/DEZrU7yIvgvz9unWKUrP/duzcNu33IZ27e/
dJIUqRIbJeT9ynqlWTkbbX8nbB4gTyCfPjHFnAxRzP5zAUc5XknQdfFPLeNP
3irq+N3M0iSa6Os9caYMn/ahYhIInrkNVjKI/UXzkFl6WWOmY7Y5dPRA4aDR
mqZ7nC51L9uchPw3M5HL5LCCYVcw6DsftkuMkKYrR2o2WTaWrzQyDWLUTvqd
xeHFaFwStZFXFjIkxyzftb+yIKqZtcyQAfOXPEkMSNxZhR/LZBMXLKVqhTnG
g8y7Ux0QIPtB0CMcLLSd4zaL/pPVHLgP8zieDk5zYGVIaVIeCKMbJ+Um98ur
VAvPGNk8yOBkdBtYyDiz+S9wnJ9WIhJWhb5hArBbQ5zT1FZlWYIGMYE7wAZn
mlcffoFVgJlCOFCnlOyQUQY5KQygn564cQETiUwyIG4nEaPbS8XMlhm8QsAs
/41Bdax9kQewl/NKGN1qAXeKrtvDmy8wnqwbUDkCzKu9FA/jmxRIlQ/7oRnv
4GQhvJfti9HE1afhdXa7zDN8PjBqR3Kq+m2if7gsGjbE71DoXhGjrved3aWK
CfcuZcOoagoDjp8NOEkyjg72i9bue7CqzE/fVUP2R54TYBmYTPP3Er7BqoLW
gppsydR3GsJgS8O+CweGMrVon69SiYTri7BGGYZGOWQH5ULJjgjFOe+eAEPX
AoYRwfNwWAkvANVsFuHWedkwnDzrnmvSJg5uJ/cHeO4+Ryz3QBYbksEff+gA
ktGuv+y/ZcHRlhC4WiGI8Qokjzq6ELVAiKmQgQ8hg6SJ//wSlH+EyToYE3oX
Pa+9EORbXPho9uOZUG57OeR/kP2p1MHoHGSU3DxCjchfPixtREZRACOede7j
MBzF3WTtIhYAMTEJzmzM81v/bjMVYfyb1XbHjC5ochZbojEWbQ2iTLFfxWWV
Ahu1sLuQv9kiUB4Qh+cP/QI9wpt8n/DwsoCwcI3mG5jp15KxORmBzzQN01jI
gdoUKJwcQJuELgU81wpzj/4isd8aTZlIYWm8XxvwKd2KuHmhZNnvS5nR1TiO
k/qRDXHoahJ8zB3MnALLohmUHsGuOpuDe0y6KzWEhf1VJXCN7pKYmpa1s/Wb
Fuf/XzE5T4wCfB20kRdhO2IAHtpfUWfs8DFzpGjdxX0vw+cJ+W9u48m8V0gX
O7uLMBZ2OYGOwyWXq0Pmid8ygSBTjjDssQgaIZ1aSyQHbCCqsTFacFyK1k99
Pv/TA6m8g3JBBKIBhlM5cCxNX7jId+3slk15Kp6aWtFZY32Vv+xAobHohQzC
xEhUkc+O5Wpa5IoTEaQoYqyRC4Ub+zUou30moq/kTd9w+A8RnOuMQVOKhOtU
gbeSlv/Rz1bfLMymu0BeYk2X24Ek3hqVX7yqwGGUVJU3+3cDYa3ihP/5qLjm
9XtgWfStV8aBDLPc4mEt5JMtXGiVst+1EaFfKkDkXF1EEt12b/Tu65Kj5Z0B
zflaX8QgIBDgIbAaEnrxAzcYFfJtrKdZtmVN1JthD8hu37PXxIEDjSDVsQdz
jBKLjMbY1BvnBnNY6IYrqUMbdGVa///cygMCUPqX39VTFzqfj89eVDRP+S7U
15q6oHgtW04bxLeB2U7hif0CNip+MuNU0wH8SEzTpTjpbOBif5DY1LLfQPgF
q//r5hoZOpymbL5RYR92O+xwAPvI2/H158ng/789Tot037bPo9oiTzZzA2O9
NV9lnbb7Y1r5xS2NveXVqB/Zm5T3q8jV8PLxhagak6rpIw3R+gm+2VSE7AU2
hYdtaA5y5YGL+HOTi+45ZuEZOh9H6oZFHCsfWsw9p7hg8tX4gtHh23VzJ0Z/
r/PH/bJqXwhCXr/lElB0WOyuzmAN1tDMBED0ZAx8ZIC3W65r4i4zyYNvMkR+
1OtMKvi/JR0NQnuAAXOIq5TksOEytORd2bHAAuF/9JognyyrE7FqFui5iyNX
dZYRrTIc0CGhLYFa2fZTtxWyZ9J1NskVQ2DnO9+EUKSOn09JCsgKx+hGCXrM
PZim1j4OnKkVfniLuD0zy/BKtrCbVF4/7ZhJxFbbyMZ2VilwpOxhWYRuHd2k
Q3RO5vlujS/HeTpoZZxmVGvY52/oV4ugx6SIPjEzesuWGnwt5IKCZcnW3bsk
jCT8I180q3fC+rOCCg7kATBTxnCvq9yTHBmjBEPenT7HGMJ7z0DntQdsUDPV
4Qd2HH5pRcux/4jp6kzsEPYYRuIJK/Sx50ay0qo65DOrV2b24O82ekaguV17
xvJq8v1WOHSVl6B/JFrIWP7AvmJEAWZmLV+m9w3g06L7HFrWhg3PdbZg8MwM
mYsqEnYdYc6pcjlZsOwPR/Z0lhf8nW9JuWkWnNNGFVvfoKFDPOJfPG14/WK3
5uqHA0BEu2JabIlkQeX6tA9B0gMhNuR817XupTCuZ6kt2R748ultdAFuaApv
3cmgJiBu/xHorUjzCpnqJrVjOmDuNv2ca9lbsYvKM9bFAZiJZHWL3Yiaj/6m
pe5PldsGIbCyPoL8ufJ6eKaizr530uyE5ehL0DebqLO5woPVjeJ7rGWyCu0N
AG41LyV6c4+fI5MeQjI+ka+5Mjlm1PoPI9JrOV5//tatgvlxKpwcQ6fu/NdC
Joyz3I/FDb7CJKihcW82PlszqzuuTh0k0NyDCeGKTBpAm24k40+RCkQqe8XI
amXkwM3IzD2uDwmJB+P9QvKKDi2nShpflDq8uSTB3ARo6vzFlXEeVIpB9186
lJ50pI8FX01J0g3WgaJK+3RiO/MU4X0tNIAE5Z1EGShKpfbYHBFmd0+pma2E
HmRrYBls7m6RaQFbx0TQRFYxfMnxRSKUFUij38QNk1fsxydyE2w2iphxkT2d
uYDI6LArjpirSlvHr2Ee0mudHwTFvbIwv4os8XBRmVib9lILCcSlle1UaKQw
F9zi9ztS7O4pjuMGRlsz60z2od7h0hj01tBKP9+wG9YGh22yTEsqWtTpJgOp
tOTRlWPZ+lrVIv1wfNkDAqLk0fF6ceaCdu13qlZ+K2fk4cWkZ9ebpwMGvcPR
WNznBavky3Ia0nKn8ePEgQ4ogRpou2Wusc5cM9Q4GzTfNWZR+e6Rk/52sukb
siHLUk+N/0SkSI8ghMy81VB/S5679LHI2uUpyvBi37Nge2MKhsY4FwDaIRvI
dYbMZpQMoQEIxPogj0RagL8Kp/Oe6O6FjaH5NsqGfUaejhWzze9oYe9V1WCM
8bScCmsZ5mUG8y2E+dS9Ch7yj7bByo4J1U4QWu8etWa6SPMhRIrI/vy0QC5Y
8NJLz2bTlomnbHIgEWFJbDXcJlvz0COAM83V8fALFPtE12ShPDAWzDukVWxf
lrW+KDv2EdYsDPALMDsGEx0Fy1x0TnvHi9RL8PfALk91YC2cCS9E1uXbEueb
/Dlh0V2RY2hY0Fg6mw2Q/DaJ1bUlWHb05UGpZq/NrYN/DI6P5FP/XMkXDEuI
yfD0v7TMcl65azdd+YhRUFOhMVuVojYSyewwqubSD7cHaldVQw4vAxcHaH4z
MVbaOOnwSxW+zvd2dnPPSMMRQi5VJK00FRHyetSatA7HFe6I7w7k563ovh/Z
R7dkX8XW4Qi3Lb9whAJX293JWbtKNMJsp0DOTfzzYFJ9+3QgTOFUBAAbYgbl
H8dlV7Fc+CQPTkTw3/60rpzJG6ORkoWfZ2APDc1UXiQsg3cbdTQYquBkSFEr
VRXVVo883yLuPMN7cViIxVNGtNqqzNzNPusLy6oe3sCEMilrHaTZHlHaeoms
+kZ1QJou2fPam+unxshSfpr4hKDhQCJqQnlrS22XqZi1OQbXXbpyYxka5pdI
TiiVHXvh2rg9AYao1Op0Hs8HDupWjKl4g4ZxnqHl82u52ND/MZRVaN6eHgiU
oyFcGnQHC8T+/2nohagogGUpkGP4ve/ZcDXNNgOuMBxMYwBG85EdOyeyqdrM
yj+0afbBWLDh2QHG70uY/UYeZlwXEHTif7gQgbsAx7en3RyXDBx0m32aSRV3
w34ihJRB0VXhiYPbPj6R2VicJ//PJU4I9SZFm4VdHYLqGdnL9OB6sDpbKbqD
0/5ZNrO9hUEZwN2Kic5F8meFvyLkF2z+Q8x3ao5UTpCrcVflmxBaqvAk2x/b
N8qw3wt2TZfIFVmd0b21WCRnmXkdR8jZK794DZ0fJHZskBiVbiXUcinYB2Sb
gJpf66WtdoSRivfnVLwrAvSwWbirYuVJ8uFaP1Rf8yH+VTlVs+Wvk+Qafv2t
8diWJVyEBqSVHoCb6ADegsSdQ9tv6Omz8CeNQM5rC12iCgONSlvR/sJdrMMF
9PMfgRGSQtqfZEQUfSQej3NZEcsu10tYN5l8S7IorAyNrFLZamBe7Kgmj3dJ
+nLo2tPe1NM39XZ99sC/UEoriRwKB9WuGTLcO9aFudfh3oB5HTW2jhb14+tx
K/CWPwEOgisTK9b3kjb7IEN1rGdRGNH3l92N/i4pWwLkhhA22ETan20k5/lf
vIe8b2t1m4j8HZDaXOeAnnrNQenKywTgzxYXUGlQRjgH40yC8xGC/nRTRJ9X
K9ZuY9EJPq09Uc1PPmlwtbWVW6GJ1kum9u0QcXxM70/Ku4lvcy4MmlIuTVK7
Md6jQSpdiz6usQ15sT7LwWvU2tZO0dzOgj6FMp3SFyFnmQIDW1zuEKPcTp5s
3u/VAD1aHQnyMBGqoCi+QzCxaxBU8rCqf3C+v6f/CP+7oIHTRoSwv+7Hre/S
ZMpaVpE8XkxqUk6g0IuNSlvX/aPwjPS78KrkUCKbCJQ6dsePl4cFSJajwWVs
T1rgJ5k6D+Kcd3QLpvhbRBhimyLcZDpktCd5Kh4Ya8btR9VmVfB7xRMxj1g9
FuKpvOIyg49hi/x+yyQWU5yEFixAFSz74sE2FSj14TgWumhP3GRRc9ZpsEhS
9tvwOYSFvrZeYNelbnhRyvgR79gpa+uSSUkybu05bXovQTd+PPnld3tYnPpq
bA2ODeIUyF6HnU5/2SnzuZ1pjXqaZA6xu91yCbj2AriOVFjJze5BT72xcw3V
Z84+SPKim57ouw9brFw3i37bqRw0/ZD/3vQQFtw3axa+CWb/sjFwSKODZBlP
FXZKWBsnszzWtkON7q86laZ1RVMLbHupdqlhwRbxe11Hm6ie66HOtCbFBwJ/
5Txd3u0S+NIwfuqYRdp9BlEB2otXiFF3nOZmzEhfUX8+2QOp5FVzZ7UprGwW
BoFNdoeb6Zq4zwU6qYL9QlRPCv4cjYT3nevfLA6HX7mliv26wXrSaX5AAcw7
u5nOyzr3qvpGy2GvWVDIE/bhGZjRL2aqCa2w1YwX7UXP1s+Sf2crvMbru6ul
uNkWIrLQxRUeHZAD9ZaWjXKo1TX93EeeqfGkSYunWWXJ21jbC2mDa8lo5zY5
sXynN2PeWH6KxheB2DC8i12TqN3udD6+weihTG9ijJvm8gD1d0xCaH8uxzLH
GvX7OQdM766yMCnfg/Z3sFpfeIMJ3GNshvMGqnzr5gGlws1NAl35NxvWqUAw
hCcxt+O01ezoG13jwcIEpq46zFhu0Mqzg0AEYc3PNhsFGHZb3kna387zILD6
+fMOMDyIp/kEBci1JPePPhxIK9qCiR8JLPGo6qZPOW20t6Am43Upz7b8v0L6
ibatbS7+A5qf9RwkFD1vD+v7Od2P1FaLqNbRTGbtQOpF7K7xAmPswf3Cy/kn
momI3xznjDR9uaJBDakmO4b3H0I4FvR2sIeid/wmv/d5bLGhh80S2mtlvD4C
4x7q+wvpxKW+egZcEiH1r82/9mNAKQIp1sv9kww12XWDh6I8JdpUAF0RMJH3
ENDMM2IV9ZTexxCQHFWr1Yzy5zdbM/SSgc+MuK63zogyPi+6GKmdCFLZykKv
jdlEth8NjKLYvr1890s5qAIH7xAkMN9CFeBlKCBJnqjH5X4FxBqdwjJXSumH
D/A2hw84gHYKoCJtw7FQKy12E9kJ9os6ZX9sEnQaUZndKiHrcPUpK6BH1FRp
5YwTlllEbUxeBbUqpJAArj70fawPgIICduTqlnVq+RaH32TuVWqkQIL7mxYU
eqQP8slP6gb/tY5t9mXtjChKx2HK9qbXQxfNYhljVF1wBTJR/kEG0KFEq5Zg
42VN79xrMzObJu0AxntVHGGA3QYo/qqgyFGJujpYUU+04V3zTlSNCJJdxlXH
K+hoQUuluXYgRJOfmMcaBgIZf0MjnDi5yCtf7HhXJTiKNElAtsFYZPdTbaBA
MQMOtGehr46gw/xpA1GalROE0wRvFOvJD3hMIATU1tzhVRKIwptp95VnlkCl
QP1rxaqoSzrNpTE4rBlOAHUIDwPdTkqDeIYiN9IytFKVfa6SyScYEyw4WAU5
0uLKXtkAsVXMXp+AEIfSW0cUfs40bOBPItthi/KFzrp+WtcXBvj7gI4ZsU6x
XKfradFFx+0ISHdUG8yppK85xKsw//jqV88pD8ZZ7J8rVGHdiendR6WMeR2w
U/GpaYqXHOIjW4DW8yHy5OXMXnYtEU4dEbZMKhdKpPj38gsELeZFT2qx/7Oj
dwIF6TTCSWirZdiwWi2Go5Fw1DaDJ1LAO50BOlCWj10arndCdvmGlbnRRG9X
nXL4/pDVWn03DAVrqJDc2dGWwiPIZJEKxka/YdHx/P1l5Fw1Hp6WW6hNpNKr
juSkOxP3K5agzWAhuk4qiS99ny0rs7QRNDDDRAYJltNSKRLobDL3X5xAG4Zi
dFp6SycOLx31nDTrTfJA/AL/kC8RjJKqTX06MbD9cMioivSuSE1tUWXKe9o7
EOIIujfTIFUCoQemkNtBBJx/qgYt+CmRvyVzl6WmMV4ShNIBH8H12JFGGEZR
wgs+9jjnOpicynQfcqb18OVyQNYh05ZGAyrYYoLsPe3ncZzDTk9Pdx7OM44d
eTUAHgjDFv0AxwcA31UAoHv3Q8MQYYSpxeFn8QPZAcD5TJujCZruB6ngoZLy
2EUnkpdhAMpqTlmTgQSpRIDLL+Z6vGWSP3bXPjimBxAmwhSZRGrMyHovI84w
ZYO9X1I1mFqhyPbFLPMnun2VdwxrE/760V4zb7Y/4flVhfI4k9BfbAWAjQsq
xv3md9adEvuB/4pPpNvHlad4hunwnV1EZ+VIsPrcTcddBLscVgNzd6n19wBr
XFd8LvwUL+5YDbeFT3oFibdHgJAPpTjwX97iz2yjQTYok0TCCvZFHVsOuIkL
5KymJfp9Ltj9a10dqv9POhjloinivJnGeA2LMz46Pcj+9nfxurCZFcL7+fhf
WAHEaPpl/LxX0W46yLTMn1acFrV7hepgSI+KtqAKCaPVcyWGqZQ9cgJJmI4s
roB8/cPcbhCY/8w391sJsdwTEH1DqZaAISYIcqLYOcAhAzyB1s6oFWlJKIfo
7SCv83BI5CqMXD4UERrIfd2vPthrDG8bK63EbIqjBbO5ACQug9fxRp73LqYx
ZMEkOt0G8Q+e5OgKx+40+ST8sOcKUvdelCiq8+mFdDFNpWmf8ayyldh1uTdN
kiydzTFKJHjnEtb5iksHrhzFUHbzv9dkYgqKUZYZGl+Dp3gSFdZgtiuC3+Li
GgraTfMDDHPcNvSPPLJaYqcX31jDZ60j/856P1w2JEkYjcanwqY3jGpujFRJ
6GjfVhGyzl32CYX9B1ChFYOapTpbeO/cQtSQOuwsknU6DAGmzlIsVwq63AP0
Jej6R/NW4eoJyF3f1iacRpUMh1D58RiPU5HEe6RJ2oadPmMIuQA2oCn2Xkib
rVdPLHsQyKO3PYw7J03ZIyuLMIp5BNoZ2IrM/lfCq/9dRvAzhrffaUvdTQ8b
dzR3loJoL7shmPCZgmXDo0lsOHIj+JTgmRn9y+7E+T1rL5S5vznS4MJ2oXWg
gv6CZSXW3HWYOkoSkpoHk5yt8nZ5OztzbyozWfBTuSwpFAQYIIJQoAyxS/oI
/TQNmJic40Ca1G9OB7+fj8cd5ZzhdFVtFCnBdlDzr+NnAmsqnqrlW/9cJXRF
mFKNpZNuaS5PJKAXURUHVhBProLinXNB+dggXDYPkm/83QTVSpdFi1lks919
ykW2ZSAcyaT05iuJQJjQUqSpyuUQbv2wKOi01WIDboIEWTB1BZ8lLOc1xK/H
eiQ9eEJXVS80SYEBOxIXRAwKIkFLjofGbpZ44Ln8t7e62+10CPUy50xSa55h
BanONSM0ule1XXjS7/4ap5e0ZIDTa0paCpcoeNMmKj8BOZ5d2AcM5vdj0EtP
G7W+ARwWeENLJ5kh3v8dOI9WgE2INmftHnQh8Sw4xcvTPUIE95LimvrZFpmT
LDDfMmgDCL1BTgjbDUIl77omlC1bn5N74xDnpitKsGe9OLfUDMqX1SQeEQH3
5TdhkVyf+6sdCCuI1osjPinPUD984NgVhYxw/jM20RRqRL1bdy+5BCD9Kn63
7pJEQGP5gH9RogGiG+HzlQVLixAY75vdNixAc4mPrMMsDBGhsL2XyzJKdnDK
F8z0U209qFZvuikblPw/pDppVs4RjMhGMrgawmuRLgUAHSDeazsPUBunHfMg
x8q5Kca4v+8e3ZPx3t3GVn+CslXnOJZDXmxLmapd4BQ8NkbXtwdN1XUroOsl
FDrLJpohC8P+Rp5fC5QJImRUBe7qu2Cv/yD/08cF66OklVDNkIC3uqSQaSkU
Ca6CPvAC46hz45sJ8wgrYlbw6s1JMz6MD3Oa1RPz30zpQ41hBlzLzlLZikYO
RfQ+nGjY0y9wlhlk4I+RW0dOzD0Rwik+R2XkrI2cZ5kqV/nbck/lrK2W6gsh
4/VVFWUgjvJG5qOzjBdOAzcM329c27GkmCKeFkuqGFRIz6odW6VV+YwvFWgL
vebGPECZk7SBrZrsDog0ceez/zLORso5Lzk3/Jzq+k307cAy5LMmZNn45C9u
Seo6sPE8a9xvonPg+DMyyD07EtPNOt9sRlamRiG4UNUA9yZj9a7B4GV0X8G2
CnBxXnnNiLvhSkQZ5c0QDbhIznplRNFSMgOSirK9iqSBJ2s2tprmiU0ZcGKZ
JA6DvVnl8KKyQEfRbjUyBifDMkD9QZTL50B/bIGdv/unbkpur7b6lobRFgYk
yTGbmH1I4CU+7QJuXjTNYwgx3d+KB3siRyBkxByD+W4dFNHbI4allxCGS6qN
7n1oFG+xEgGX+37+J7QF2W+OKBgnbIpwLh9OsqN6H0ZctzH7j8rSUsH+gBZN
Xoi/rWti84+d9yvWpO5fTuh+zMGxXGXgy3SwJ3IQvU5Dj0B7rU3xlYubJ9TR
Fug8yCnUJHQNn9bRR4Ig1Ij1daDnnNE8IfPY8/F3P+SBLZrx95TTgMipe5RY
x/7/lqdD028/2r0m4kM7J14gLop5YGdoYJ3RBbzscSqg0GEM3Sw7+aVuv/1x
inspFA3x+DqvRjEu4kTMt7kXSM1KDCSNwq7VcP3pBcrd8BYI0ZiTasL9dRyW
r0YSF8A/gixpPPuO7obVk5g9EGlGBNQQhI4ON8xhVqyd+2+M7CbV3rJ4siFz
R78KpNyY6i2Mf4T7DMkEhgLj55QwvFAY6aIj3EfAWT3XJOINWL9nH9m69v5f
4nNElV6sYAm7scvOEy7BLsOwmmsCBEdAmC8IdhB+szlWFaLNbJrlJow8vygD
d0L9g3S5XiU3GYf9Rf5fOdhMEK/KIow0tPtYSrESrR+F71OuDnFPqUdv3NBo
5bk9nzkYcCkHyNCbLWbLa7FdygQGG9//6flRtfnN+/asj3otKuKjjhSQdtjy
DGDLm/dRKmtCucsIsqkbQyG9aalBVu2X3ZV1hVQ7aNuBbGJyxNdVNNqaqhjp
UeycNAargqQGp0wwm+fWuIBAypaFKnpjxDAEaKRoAsrSO3NTD8pB9CKVCNpT
rRXm08zyvWSAIHU2on3tRbCxs50lwqh0n7VtwKED4FZ7pQtSJ5H+QyNfoMDo
Q2FEMlJ7wpcAwRF6ZxgROhcFrOPUPnzZvsNIiZ6ADiUZnul3xuIRh8U3d4jW
BOnf3w9tjJbxMXZEtmBQ7yA3kYTl/wQUe6+v5/NzHjC3OwM/4nZC5xxKhOxX
nGb2lH/pL0fu1jeqkTxHWWghuiFoi6eg15868+h1ttM0C1kOKFxuGcPkhqK4
eDx+d3zqYvr8dVHxmiWb9wabwkcg8P1DN2HMsfa7r/AQ2tJYNtIuVSyPrAfl
nXuEB8Zd9XTmWb5N0g2H7Fq9s7kPBiqAzZt5+YLk16wJGTp6eWoUJo5F8/ML
X/wtZKIdJUjPuX6zlUZXD98zEMqR1lR9pxhdEB1cx3uvRHq+zsVo1uXuTDgk
fABEeeJY8wlFPXYKUFKYEyVO5JLt+UdAr/Wt2Ugj9LPtbjBnfc0vzDDVPS70
/RfTnZ9JUftGRxf6dwfz9yVm8uyUt13ugNoShxQEni/RlF5B1yBQVpqP1EU0
i3xdFV1oLcqSxB/m/Gy487OXWICsWmnWpQ+z4w2/hnZ38mhlkmrlIdpxfWHJ
P8b1Yt5NrhH7v+THxQiR88GU5IFks0Hw0VNeqkcuJsJ+yP5K13JooB8YDnGO
p7vKPzR2BSuYC5r0bKlOi1BSt6t9ipOu/N24gS63WX8DT0BeJ5hBhWzDVchv
F9pRgjhX1gg/g+2Qeov57sNlnrmfW9iBP3SHZ7VCMIz3+dJXewgwtwrhiwBM
jNASovFUBbynG6pvyaiE8qOpIS2ytoW4BkCDo2R9K4j8pHr5kV5+l3Im2stl
7y+bphAxDL3ciPW9nbpQUsa8641yugaX8i7hy3gNh+xWmBxC37kd942t5eWs
U8cDCPpKJrKQCTCrJySWW5bV1SsXw46bVpHDGLdvbmGlGtanq771vkaOHeHi
Busz5SW2JJm7xf+iSli5sSsqw7N4hu5D9FRQJ0gkRXbKvJqTITz4fKOSPsiR
sDDxyPTNAy+0unqtTQCGvm/SEcZzobHEerHdxS/ECS8wWbRmUVMulfd11nOY
ZjYxMiOBQvP04uymRM+VwvZntjb3vvDHYv5UqiH/iKoEl0pjfMPlxNyncrEH
9IgUNw5R6N0JQnEBRaJYQjNm7fRFt3ZJ7kcXAovNt21Ggsqblqkmq/Ph4Jdq
nrQi++n70YEqOq2E8qe8FZaJHx/p6wrdWfNLteePcQQIMRWChD/dvSN89Pzk
ijzwOcz8075fWlvAd5/QbYwCUbjU5ogAjn4p1LKhIeIsALrJnGS4Zlrl/8c+
EpFYWXaYRp4WXeDrhQsKQq47yG75oxRMl1Ousd6apTdIXNDY8s5yCwbSANBm
MncGZj//yIpTwPvuftnATYFu7iALen1+UXUDLzSGlwfgxnKj688UgbOG3qnZ
0JPw1UXu5ALt1tF25kPCUvkILETZqWtyPfO8O/MEi7Oe8Jzee7F4XBPNOmW3
lvBfu5FGfdSgicsTdhudZXJYY8obmividpCInoEK7nwphzdL057odn2bBjYr
VK1g4W7E4dexgJp3LyKgP2gDtbazmZOeawnkGElsJLKdv+djpLegnNGdJAKt
+UqKpUB6RSosHqbnTfSRQ48cVsgyW1gSYN5vqKyYkcRhhirPbe0uCTWUr9D3
5Y6NJCR/xgquI/I18jB8AfPMOsDZkY5sonhw6kz0fWUZjO/X24+sXJuKpIAZ
vvs0zrdc46siArOh7H56TfCKbvNVbPRPONlPDuhVXsUjpmKlMiesp/lwW5f4
LQ34PvDwgRLdtwd7klRoYoIuLCrkuviGwZEtZQUvjmyeurzcC/fa6x/op+Ms
YJBnBTFc57kRVIxCvaLEKi5Q1Em1HkIRl60GhpDOXD0apC7OX6vJJayDlMxx
oEdE0I+1y1epsnJZrT3odJdiX4e341646jHYncGyWnG6ZB7iohu6R+j0IkSc
ev4yY8B1RgryPwflATWuUuKvUck14WmF9gvlUedvcr8Ktnfu0FbJvZmeZRwq
kjcIH633xlNk1Igmy0+PYqRZkLljO9ORO462kJdWJ6DzdGz1c6JKxXyMw7QA
uCBL82lL29HsuMswZH3vNBpCcy4+BSIDmIDbs4NuCkjDE5dhitV6rf54Ixqr
RarNAX0XIYBMjn3o+Ct1RMT8gz0aL/ORliO82aCRZoKPNl+56rTA77M3Hhpq
h7iMkkbnAP3T1X0W2sDcmIgC1pb5Pe28nrX0Ih7jnXDu/FusesY6qFXOHz8d
4ROGlKSi5ac0pIfHiZlXkI2O7zZHLsrPnRsezc5vPKNT2eAvoE1EAsK8/2nL
ISTPyC3nuLNfiUIL0JIl12rUpT6KbB/HuYw4d+1rNgifijyymKBaUL8pbxvs
hCvWiDVnb/QccuZ+rK6TOY0j0Qf5HYToGXlyC2FX5e5FwFOJoW3FWr3S4R2b
0AHzgMqpU7OOUE+Oavs7yEIYohD2tQblXUkDiv8DxIc8sxiYVv3WVlvO81jS
3K5/Wn1I9Ld/FStGB+L5tHfaWGyKo0J4KWEi5gMk5aDqAlb6lcGexTHbuJnU
B/BeA329UfhRPK4PRNVHR94DelHTcLTEaWk9wEMPpn5IT/T5U/F4wt42yNxD
J1DP5B5/ejyhjisgW4YQn+f4FI1z9lyX/QmDiz4Pm8Zjv3v6IVDK7BPZL+EJ
sH1SgdLVuJSE+jCsNs69XL11rQAQgMdxBXnyyejcjdmVwzCCs+vTLAzjhZuV
2TO1zkXoe+kKUHZEN7Bq+goQ/JdjzO/zEN4SLYf2j0uc3aZjQ7muZpaquo8g
eyItX0dxKx+9N4slH9V1n1zxIRBWUF7dF+f61vGwWwY5MZ0MCU6kDRag5mUQ
oo1C3P69P4t5/dXME/A4Ba72yIwyiCVrlqJ/riCAFslDHCi8D9Bt5weLd2l6
emx9xp/AmzKxRY+T8i2PFcdS+29oJiCtPpiaLSfHeju0WvbXW3nVcffttiBa
iLijpkqXSZegFDBF6i5SMQzNb2xPhZ54ZPXpUH1r+f701I1drm4THCWMspeC
N9iHsMWInwdHn/YMC1RSaSVfq/7N+klw/DuUEbRfArP5QnnUHM2ox29CBmLp
Ly4OPU+j0uc2X9jEr45FDJqlmFj0ooQPBD2Z8kHjmXnmBaCvViglwKBDXhrM
ZSFRXpoC8R1GwJO0XMgMNSwt8IiRW7o32FnJnVfdqe1rGDzyvs460P9t64vK
HZfQQb1/KQ0ihtmUWgPx7/6oCynLdjPrGzSUlYk6SH43cz9CIaADeRLZh0+p
XRfiz62REhY2ZvwHhI9WhKfOk+juqDl8xr9KF/8Q4sW77HjFsnMEtgx0HSX+
+dsbEYANZ0Ey+f04CQtlD+bhpKYMtsDs6Ja+nmJp0QtC8V3gMblmclfIcBGz
0CrTWXZdwXAcxVDICmc2dsL1w8v4RE9mHrK7sbeJuYfpTEEBvLMXFzzuSMEd
vWCTpWcpH74EcOQQJhRpjzX8WWzX6J9MMyc9qWc1FvMqFb6IwMRJXPSU5yGp
OgnAHPSmOKJgdE4t5Pmn2fyBsb3eHoU29zp4Mngpg7/4S0lijRPVf4RXVIlp
KMC6I/5wLrKG0DnhSIukL0M9TedJi0zkmTx9pA5P1a7O15s7CY683r1IMSaa
aGseN1IkwktiDC8/EZEe/NdNtQwk5YueISue/UuI1UDO+AvcDqEpzF0VgBy2
l42CwXRm/053ZBJbg1xlZ6ISk0aY9QpAv1GplNPIJUWkGulsWrcR2U8zQ2VQ
JUKYj6bdXrgrAAxVYPEGLbOnYFMEEypoGYjzW5gLZRa2l/hi8oS3NS0VOXAt
tnY1+Qd1CaL9QMP1lH5Bw2MuYRAxID/k2TajsfGt98uPp5YAqqVA26BDSiob
61W6RD9nlbGlnwY75XVXo7io9kVxhAYfQ/7LhzT43czS5rJqOagcGTrXQ+El
GiOSMoAfzi2DaAia57FaIgte7UzaAJ2vX4e2RbZxbhIClV2QpFQf5w3obp5i
whP7xRI0Oy3xFggRzELjsm64rtradGbmRA9hkxXvp3rRgInVFR/G3bnLn9Om
iMCVjiwBLoQm46elTL2l2Z2YqPn60Ge45ZUt2I5r2dfeHaTliu5p3KzFJb8q
RoFNrBIL2xKFbi5hmWDyC6XlrrJaBERzk5BBBIBxAKNZfue3yPjniiqJbdav
F7ELEyhFlIae1qtCznC5N1BeFku3EzqHz5iHQrS4BRmyjqS/aHzx7wLF8/J1
yfeHdNQp79E77NmzPE2r21HlmuQ72QvtxceOnDBWQzapBibGETpn623l++Wy
9YMVwtkh9tQFMa0T/5OylUsMS7QnxBwvXL+cLPpFv9dtOS7lOUYzJ31PXY5y
pa2BTKKRNrFSShBSDuLe7CkRth0Fuw7MTMnoLSLSDjLJqLCoYXdlR3aPrYee
2JKIoiBPb3paUkQoVonjbeOH1lP1TXVTQDZaxRRRF0nXkW1Z5quRsygqXhci
9k0fxIG6itcLSGU3h4XlwJfzI16Q2bNuGqeRNFIZ46fcI1+nSNiN7rSXrwaE
4zPO/lnJkh0YtYmiHnCHIwqqNw3CbO15ig3C0HrjQl+WIR/5ul3XZderbC/f
6vC7yla7VrGSggttxqqv0g4k3fNyBxl01o/a5oXQ8I+TCaG9/cEEOCj9GOmD
TqS7wUGoBIxjoU+sSBqmOCrLefDfYYu6zmbGd6umz4B8ismaS4cWA6KX4x07
AH0onrG1b0UPXo2r2zv1NeT6bDIfAfzpexGU/s3gd8CKleu5/VQW9TOlm9PP
1PM5SUQtSxz52la4Qq5n59Fm2nypZQ7SdjwzTUCsacsogmCaVD1O2NnjaVr5
zTpIx2zd1HsTjwvH8DWCBWkiARG/Chr+bb4SZCSY8uJxFmMn3Heebjs0jIoJ
1bavWDpxmoXu/q43btD+LmLx8ijeO4eY3h4oj10yRTz1sMLAQmb93Lrqj1ho
ivo/2U+2D3P2BYP+2+JIKRd4sKqz1SYGvy+Rrv2MjhQUVI5DIcwQaGdGGMiR
0oPqvvVNHhmQE7Dbs0m7+7kAJVQqJvL2hRgmGWsdddmquQQfklu8MNoPu5z6
VqZB7V8pz/v5MwjmYoP6xfGMUpEMigWR91o+bDZ0j2TmDZzSKngo0Wv1IDgU
tqun2bsgh6s4Ky27xt2zhgl6eCNGKyjVUQt3YkqWBDxytzM3EVgfGCYew+zb
yA8O9RwJWpbk2F++VYtdNzbiIDJsC+zHmBM3GYWN1M3qdiDpE6zAzTVC/smt
lomr2kBRhOkLTDePfrHlJHUYjJWd7QzIVj/3Ol0tx8eczYNt7AjR/L7JXy/+
B+EcWLdzY9ctDc+xHTs/srCxiwIfISgbSh6azAlbcKNAxjSb2TDTv3Y4f6qt
hfRW27GyZI6rfvCApWshWMWfw0xbDlXl6XGb7HSE03YKvoyspKdsjoOMAHaY
Zn7FjrHSdpg6iJD6IgBtMO1Yp7J02A4JYDot7i62zwBfa7cKWpwxKnlfRZjf
sKsBtXwAokLfonvGl3g4aH0Wpk6gX/mO6dS3X4SyoCm0Q5HbQ4M5Iu4mr0yH
HSd1Redv/pTJi1kRjNAgyakDB4wV066NMVn8ySnd7WzkAVYHyW4iOHwld2hP
6gakDK56MMexvU70qQXC3xOupuRxYmdDR5XP8I1UEO44ct2zyw3yBCtUY0lV
nGOIXuLAJAqn9E1mlT1B3BBdT5lmERv9ZrhS2GC2+h3drR9LPGA9E04AJwN1
K/6OzLsKt6HkbhO4zO//J/Pxg0IZMbdFjKTCYsBhg8pS9yiqqz3+yPF5MIpa
+uL6AI3/FC//WjObvMoVfLqbCOfVRXhTJvqEW2VS9o5L5MqhWj5/n5nQP0wG
u/gBfuQD7mx2GBWPZeyWxP+0yFKDK2dEWHSDIEmyb43/pvEHgPUkJiuKkBwv
3+ns40GaG4VSUkfaMrFfhIzRtbHknrOhotqWLFTuqs9oaCf8m6h3bseedfKH
2O9mngrysX/ezv7sLGjy4l7GhEkqlmBeooRCa3VvQJ/plUuPK4YWdc+gqIIn
ljNRyUnULtMTSx0jdOKA5If5sNQzJW+vG6wpdbHlKxmARGUDQXFNkUbSMvRF
crVNlE5cOQzQJXXp5mWINuXp1M/RG+qW8I4gzkQaFgJfN5kam4Yk5FAZ5CmR
CqB+n7uDXscwcquLmFW54WXxd0fwVlKLzo7fUhBempK/mvZz3MYhmKn0WBXF
Pnmu8XxHQ4PygvAAVMQIvNPmWnGaHdn8S41oRtGEDzhWk3tDDXCrAUyii40y
v+IA/DhkF1E3kxw06U8zAq4apQ/GCv6/zCvuqFTFxu3AVc9Q2cR/cKJv5hBZ
LR0K7U16Fvo+0zECUseFM341LAiMH0opkoFnLsLvZoYb2elaqdlMNVb/rdh1
66nE3E7cFTcwfrScztALt2ob0N5AobKPp6y5ZB65sNOWVs4Ua9YALcc16zaB
tX9HANVih6LUukkIbixb0Z7mrE1ANiGz08tT86Zcmp5dbwy48+8ig7z9kj1i
iwBCeHyh5w0SKJVJD8fBzXX5p3xMAnwlaYYgNs+vFkXnZQJL/vzzKCB8nRRq
ewgAX7hhS7oFKQNL7nmAQ7Jce9xdOxvAy1+aIm1iCToUhw5XBHCkomBy7Pxh
J61KW9yUzygaYUXLsuggFecPDnrs3dTaHpDwLfkT5n5OtNP4O5VhcULJig1G
r4EcCz/LKCBf0F0eLyV+mmHuw6AZagE4P6p72/uQno83miFBP7fbllDqrzac
mjFvzwmHwEjc9keXeK9cCHna8L6FGDXSiSxl8qXMkNduEI9mSa6yJIBwWXQq
3LHjzCoQgaR3Bk7HP8xv57VDkJQ1WydiQw8QRsNBA/2c6xApLt2QALH9qeUW
RJc74wHoOHPZtPIyQnG0TtXdUP1ycjdFEVYZi7PPk71ik3CPlgrocFXPA/w+
r4bwK0oQqVzwp2PESM2kt6VA7JTC5LWlalBHhsEKKFzf/BNiBQK81dPqyupI
sj2bWM074qXWL9FjrpHriW6REamdrvZz6pu++pi94D5/wOznI+I25aruylIi
znkBc91dehyzelFz9R3FTQYuzJ1H7+VPFxlNbKkn5vc8NDfuZW9H3Zy60uX9
MKHYGbLXWOSty7i9rtCqEhOggXQgI2JTvEmvICN5BG+9NXnZgA9I9w51I3HM
nj5s0xZraxJZYvP1xfbX8iNsD5pB7Kv+tlFiPwhTNwjf8/OJKkqj2jBHiklw
Z6HULDzQ89h1Ft6YTV8L3KeD2s3jvL3fvhim2lsymCoVzCpDJPcLbqHWo+P0
4+LaY+nbkZ1dWOJk0WHXe65bY7TfeujROvAXbYOTzixqGx5Fe2Ts081zwsIY
tvdHDupCmm0c4lDPS/GBDLiLLDCY68mRIcT3KypzrYUqVqVVRhSVioG6c+nS
sRqbF4lVCjyOKxHL+3/jLZ6EKkxtiMH7ehKa7uWRXujOuc6mApcjPqRRHC64
KovA0nHmioSb9R8jxQ2BjM/f1A6AK//GHBTTvDzCVfqveYOxildMqjwRmrxY
78e9UlMjArWrxbE8CAKCHMFQVynbC1atbUrdsKKGpN2n8fRm9pFTEHFpl00X
07MRZLdZuqJJbfwuUt8TqLPv67YH58IkdHb3wsvxfHfbecEiu9a38MVWcvP+
pTLh6SlPYJVCh7ynjlAA6IH5pjUJKAZEW0hpDGRjD5VClwBH6y5v3sWjiG27
dGoWQTHpwmm9LAYwnptEVkmFXRGmFCNTXdeh3X5OIW2A5XqHiMiLnmGddvGb
25H6kryW93oaZ0bRkbuNaLevsk0LC/5+SKnC00IKeso7NT3B7FS1ayn6LKLJ
VjdfaEvnkI5vjsIMjglzWnQADi2/EijqOr9zoYTSvty3gFCjoN/Ieaqc1boR
51iBk9BEjw0Qnl/twbobzzHsvxPlVp9bom4yDE12a9XdfloYj9ZsXUkYoc3P
gl5KoLx6zp7w+PtLodOgQvqXxUeLKWe1ilpRqaY8TBZD4mTxZzLs2DwxwBDu
6WcpZe8G3Pncg+tYfVHTse9GsmQp8wizMKbNc0Zt4DFsOLKmnGnp1RFoN8L/
tdHNoIuZ6skPKcO+Qpe+OUfktGK/NGSsdS400oKVltci/iHyCef3beDuSP9+
pj8GWlpTAs1K9G5Wq0hk6yQ5u+ba33oxDV42NiSD0SB8cPoCk+4dN8f/1REd
yz8RdVDwxR24EcaPsHPZ/bfEzH/fBsaAsJH7Or4UkJmFkEj0fVu/+eAM+Me+
yczRKyKabsHZ7uHCECHWuOr5/533ep3tzishzGedRtRHJC+sqo+iNzIN7Tov
ZIcat0BlMM0t4L+PIvqOCeCxNKnOYLTn5W8oOlV+vHXYZ/IOIbfUAASK3tPq
wv0WqFgg2kUp1acCMFpv/qN68qFIykvS+zs/n8u4nGhnTTZtqHt8aaULD5sP
E+CYcRNX1dmmPvNN2CctOR7s+DBLs7F6SLxPrnu6tLU3908K6QYUlQONOrx9
RMNKJUs8h5jwmn89NhHOVtE1LqZHsOvNHMtQsW4lzRRTKOTzco3+VHHth5oJ
EkO5aOEai9ezkHEuV/f4ihYoOhzIbHwdjU6e6QkWLHYK9UU6/y1P3GRIExvE
QgFzuuyaWV+bvys0XVTDqpsUhVKV4Fx8ZaRS2BOBTow0oovPx30BawZPVnqu
4JOCSLhbBnu4lCP4N1LELZvQJZVecI8psCvww2YEvkp6U12fQcjtlPU0zTqR
DiUWm0v7aL5zAObS+1Wzyef0YTW2NMNG+0afmWP0JV2byiEtStbNBsVM0zLJ
DPFPSrPdya86gfMwHrTZNuhkrMvd6fwdn1Or7RreME2dwSI+Qr4ucGJTnm2w
7wito//wPmcVR0FLOPlYSWTtHRZnIg/mOpeLBKPGVJDKaXcYlEggEuMxZ/LD
xL7sV1Vzjt1iphYlNtTuTYFVn11b+SgDl7o1b8syugdyo4putr4j3zxrBXMJ
nA0ZuLXzB9Ln8qfQxItGPxmwMmz9q+tl/qLY9GauznL99k0GLA9muw2Ha7Ib
Pg80LjGeizfkRgGjMsDdE4sGZbMLYe/mRGtDjVrlNW6d1TEL3gIRGSYZdo+L
sEogAx6hvrXB5a2/ocC30aLe6JgPZ6eArcQKpqqbVrLJjICYm1MMfmWkKIwG
kPk9avEcQGVDvQ/H3A1x33utRo5GV2kn25IP0KbQTUG5nwBbGjcbzbogvZAt
5pUqOV6Itu4cwYs0CzYCiReDs+kAFECom/D8YBy0wvXZ/InrHdh9QL4vOvuv
irefW8NtQ66z+uJ7WLBRogD1lDcQX0+D1hhgO+XcclvPsaYgymh/xuR+tup8
lAUmQrMmiJZPiC54nzDtCmTkd46hc+9nL3vW1skmebh5mJZyMK3hPn+5/KLT
vcUBxWZJGkoMsXTHnzD611YRsYFCfbnbyZ+45ffY5zSJOia7audqAtlyXLFy
h8SGt9utWUQBV1P6xY+34YYFpIYOPzwoI4JBLUsO7hD31yslbia/IFVsnq5L
caLF0OmJA0FJZtY7U6w0M9biSJExRuqcLiiAqfr2/ePThHtBt7+q7N1xYVUa
6YKwfeoz3kmaPb+O9sAQqPc/6tWdgnz5B64wVADrj9Pd+Q0pICjA2njSCkCJ
fCKU1tBCk3M/ai1zzTBAkUdAqPHTzZ8lqFqiXP7u3BGigZy4X3dswx+4wdv7
d4TJC/L3oP8o/UJwzmDelgrUgvB7Tg3clsvj9L4lCUuG/wgpULiw3EcDRMcC
Wr8/JLTnuI/nw9fXVzqST8HQpZ1TE5OCbf8FQro6KZREsWrGjRd2TUPs/A0s
net0y3vFdHVkti4a5aK5a/ULW7saCWhzm+KkuHtIeS+RdLSBOGX5MmcKbyUn
z5W40HHwNOq07TUKBAgO9jcLmtW/snSjLUMiYaOzg4ju7hcvh84vOcwLWg/L
YicvRyikaElr2EV4AnAuln8FIuZl0gQtATUkRN4RReVA1hBRSo1dMb3rHYJ8
HZ4/QgTP/mZejmiIvEjmonxTM41vOTW+BW0O8A7H5Jbuj4iYYmXt128wakJq
hqctXRNBLsItOqhI1ZIX493HAXH7y/KmF3qGPVlV2qm7DOUNBzJOqa/jMyPe
By7sJHubfrVzXuKOlCQ4z7icjExyxJa8RVQNmY6cLSRUct0RJtldbdMKwvOG
nl+M7X/L99IV3jvLZhABPx5y/z3DctropEdexHLyfoyjgg1thw0O66WUG/yL
yNPE5UKWM3M3GLhrPQgj1H8rLGXm9kyMcBRXHSQLt7Xv5JQiizAy3rsw0d7J
H5G1bTz2QxIKPzsrRfcwc1kw81KQFNaCtwWc9Zm2MU5u6POnsv3YRGWrQbiC
bNZilvzLhC3usA10Hu8Tdw6bi4tRHjYqml8Czq+KcDqgW/LlQ2KLNH49JKzD
o2cgC1EoTYgzA7IDzm49/E7Px29yFo3uwScO2NCB7gxO2WX9jH247+3+9Eyw
4TF7MuYQXBnvVl6Q9iUTpfrTWF5B9lu28nDO6amnN1GaRc2rPI3x9rwO0Kig
KxRfm0P5CBiKHtqFX4ZRXwTjiLgPg449rLLjPpQcNF1+vsE4d2TrVIOJDTbC
OoioFFgwhjQVqdiADrVog5N1ywK/hAyQFqUs3pXsX94u5GnjqR7pqUpXBDUX
e8JOojLoJPAFJ4W3RhbqKAlFbdHyggeqev96DjaCTLLXPUpqnQM0lEA3VnFH
oO/7XfP6wsry1S6g6NP7hNZwwl49WeLduYKWNJ8IReLlGiCBC3BTiN12bO2r
EfiV8K9H6vCt3si5w/zhtn8vxBDUysT9ANnJI/XzAdC2rAxQe/w3USMcnXj/
4J0uHziCsfSSlKwCYaonpfPWpt3C1TRvMcHEc/ieGWY7NcM78nsseVpoZh7Z
uoRiJuPzuFaho2gsBsPwdCwqQQ/lqVlaeow38iJUZlftuCFMlgxR9hroX3VW
Y4hWCXHbGWM830CVaHAqJGzCu29us8hMVmlze92rz/2uIavTfJFknjt/KYOY
HCvOzUzXCaVQ4Ri1IVNu0vjGP8BhRU/OFMRGcvMqowoIoiK/H03QyXLfvOTt
uv8sipSUY2mew43UtVNffpLaHDDKK1dShKYFT9+HNSTESnVQno39D2MkvJKf
bDurfS2g6WgfOxpLZw7x5XgDWgi24UntWzDpDBzYd329jPSDuk5hkRFhk4hW
0gS8ghKOpunSH4gHg3AdqIi0/hunij9AqJOa+lfZ6nFob1CAXP6RsiVuF3T2
k2GZzVUb1TRPKOVpmcQIGb1T7D5UKE7cup3zVav9Xy6qmyiKP4pmZXPgHkU6
mKXm88BdR9m9xwomqve+70fcU/JUS+p7Zg2h7RgcS24q5uCrI5dndzToXEyF
UrNBps+BT3asoxiH+ruC+sE0/d5ch9w+jXPTtMZQsSGQgonCXTNSQq8Pt/D1
lA8XVWFhoNTBXBHmwhWMQeNbhcctMVm/aFrzeFVJ8mmNalejOROmnszZ/AuS
x1MEGx6A2t8ERIdH8duhP6kUSxvSYdIMhS1x5EV+dd8c1nlIKNCOO24hi42n
7sKWERhECCQDApbz+shx851PztV6J5IqScGg49qrJb0NeBrUP2McwqqBz2he
2iB4zTtT4SQeQkTBgFkAa27QK0SsHBOf7ZwfBLXFFPoEGkI0pYSP1XEDkpwS
QnVchOFABZlit6ynm+P+KwYNjMwzkIYJYTfYNktyVV8i0EDksbwtYfJxNyVw
hbYE+bG3xK2cQIc2FpL/kJJTw4lDFF9y5rzp/UxH5pYD2dzLaZkT+FKYPUGz
AYEzf9GcCKiabSjoZ70b+RPEhT/i24J0DiA9ffc8Lcg2nVeCzPRwWd0M6jFs
/dq/7lXxk52PTMtorwXB97jYqyMUdc2+R1Lqu7OIOLsUhMqJeh526Xq08n1r
D7iaKxecd6UapXkvbokMWwUUTAyAmu0mDDwaXdPPAOHAwduYv4G0zmIILyRZ
Hka6wJMs4K6hsEz+HKBlscR7dpxOWIla0UlHDEmJeTLjN31LIJBFMbvllJ93
19Ub/EVMNnqxARptfowEcpBS0J8S4FdVsepv3OuubgYzH3Cmg1df7bzv0448
x6salHDohZEfreazkKgMZIOGUZsaZgVuoEZGwNq4dwBLw4qzg3QlQ0NTCms/
x13TuKD2OEUacgrGqQuBah60nQ5uC+wiqf8oe4+n7MsJk23HZ0sBChwsVE+M
L6F2bQRW1t18AsC4aaWgazVZQB4tej7BK4054A/izhDgtCMSjEryC/GRpdN0
9Fnilso5WWcDzWjngG/2GoOQOF/bOA7JlCFnl9il/Kri30sCekiURWdVpidU
LfCpBs0IaUIG3jCWK6pMtwzQJQ8AN+c2ooWNCoKFlf4sHCpErlKywtoDFUNB
xRMIx1pX4XFmTxpESeVQgfAR4IXYYJvAgwA2A4M2Bz17dc6IKgkS6EB2fAfH
HANr0sU6htdl5c2P8tceLUg1DU2i0JgHJaieyDHmCROrqKQgu8okYnVC5Ym4
kITrbUg2q22LD4hvxwG32VPHzangaRXUNHdX0JhOuUbgMxqbqQqxqZ2nWLvw
42bYydfS9mJBJPtiSRmviQDoUl96Nddee6D9Y9urYHYH1rKYKgY6dZvZGM3B
QSNn/bLms1HtSjh984lnClpEL4hE0TS3HV8FoyhpR57PYnI+qwtfNiI33Rcb
bKUdIq+QplVlhx6et8WKWNOo1s1LrqtsMBcu07dTm95psiP+LhnIIiu+e3Ly
GGWiaMQcmaFrOSUi+nPUefFrzUN16XXOm/RxP6gn+gPIltZBVKF3srZ9fMiM
+gM3RvLxlD4A1HkLoTCSInIklsWZIUJM5zgzHIkib0HLHsha3e4j+YT5O9Qx
GdEtziRfIl+tatwIDkqTp0qI6rvmJWt5UriOprrWNATEwF6hN82WkZS8E+4Q
BGg0QOLpAnCETJc/kbLaGs9fOcdzlVYl+is8HewR1p7CfVfO7suO2SVjzjyr
AWEIOTkHc6xnIRXy04Ma2QPRj1sat9XlSv3nycEtnFiNTdJdBv6m3dIN4kzm
3mOYPKmaKww7+Fyv5K+4/v5uC2vOTcijezGIMFl67eThOOF3XgzvtcRyWdGu
nCtwurpcxwyoJRaas07lBQmFYlzASYQMdFMwOjydB5vbeki1LDlAxz9D9KaS
aq7mwx8WbSKEMy6Rq4t+IMXxgnqCUOhq7ZmXgBKbVuysdMQywO+RSjBFhdgC
lBcLDnV5IiQrzOuSgNiUOXSJQUGwsgzypQkJt5hJlm4l62CoRvau+8K7Nxbz
bFyXiCdUZM4ymo+VXzi3niOaKVT9zlgzpPWwUfoI9/gOZeELrRR0fHZFG5w1
3bAUg9sIuKGlWX9g0tJzapSxtnb/hdtcImLBR2n2P6r7FQpNXK0wY0lw9pKh
UJHcM96gAKVUa9mHhKgAmLJ9sDsbbZbsQuHCVNufWkerhFH/OEOFj4i4fY7w
9cvzQ+1S2tHO2nuiQJHBkWg1EJ2pJHNdCMgdzapXk5Cd5qmk6SM278SYpOCg
RdXbAh9GVfXOMfh9ABw9r8mmIgcWf5ZAkcB/N32kZ9mICJ/a23d9+a/X6r3B
gsP9UFvh4DI8JABUoGtmVg/aq5IE+73EPptou20u8fabLU8qY8d3Ii9pumIe
PizuNGkXRA7t1XTDnSQPaZjQ1LbKClzvFMihQLYxCDqfCsGz+O2P4yWFTQIf
VFCswVrrW0TvOY0JMcMWFO89P5p4NU9K8Hp55BQNH0qD7Ksl5tlFymE9C1hR
5KCDiNX6TKzfVls7HO3jNc9y7jkOOTh+xkhRDBrDyBn9rDsxx7AZJzNZaUHf
/PxSWpfXIs9h4fgNaCz++VJQeQFXp4cRQqUBWHtmAtprEwOjgNdM7Nn390N3
Q+rEga5QFj0mziH/7AjmMULt1ebmV+pnqvrv0ulGDPi/aEju7OrVqcKGtdKv
KxfzytIFS4PQ/lxwvYFp6hi/R2ieh7Qd+biLRaA23xpHcenEKUIjYiaD3cmj
l+jQnm3FkVZgWMGOoN9/ZwYzL5Sx1RMSrz+aSFnF9MJS4wxLe4YAv/KwcfmD
HS0oYpTG0iNjOroqyrljWa+oaEmcWmYdPRn/CsfO8G43WqOTIFnh4oYFD2Sm
WGAnYPfRQh0q8T+bT6zMwH3/vbz6zBhXUeCe87vQsO4C3GVBduoG/YEuM8RH
C0869iZd7ewx6243ogqJRuirkck3mHeVv2uODu4x3lNzv7YIrfQonWez2Clo
D8aK7Y0Ov/8NmvQS6mQjye/apZGnma94C4YN2R7EE2DolbwAQ+1rmymqcd0G
LWV85/VPtV6XE5AOVsKu2OPIPoCbqo7W/EOoJTbTFSCSoKS0WaRUAWoiv6k4
fXCsw9eZgx0qo7LPcim/J+aRUdw1ansTu5wn8JLb4NsKDdhaisIiYfhWmbSV
hk6z/gCAvhxU/KDIXWowbe83kC5LM+PjpJ4DSN36BhBYeGp+styErPWWEjPM
hMpIpCpfku0xg24slDM+GoBUBKKr3Fhx0d2imKubsAXkM4r6zuNUZ2X3wQKh
gY4zYo/Cmjebjw+Cw3pcr7DxUkyFFfpyxVmh8dbbFknf4bhL+I+/xjn17XdW
H/mFzTvmaiZGqBB3R/NwquqP5rOQkzOlLgz30Tr92nYQgv2NgaTk6D2KlXhD
fESbxJq/BGU8wroY5Hub9KxuFLqIsisWrbJ8IdZaF8xxMIjGmJ3It+TRAWZx
yTOBl7LGXI+3jewXMTDIjoAsaHGTFAHIY5YUzKJCRWEaJcv5ga5kvzkgJyZZ
48Si2T1LNaRmrRHLKM+wLGA9aT97LKjRi4wfZdW4wMH91ydtXYZ2w5iVNnvv
ZKOw8VlZe3Od+olWgnT8p5iNues7PR1b+b3wW6dgbrvnFxMCFUwQg3yTSSvl
N4kDXQUvcC1MG/cKN2NjhiueAC6SZcPWHEx60H3uv7/P6sHsGSSQBhuCBXdo
Q3wSfLaBkwtANk9FZ7vrLsd11NtV/Dxmi8pCPttxuS6skAMRVTGgQh4sgIZR
HU0XKeLAG3NHfRp7gUSDs91RvlPNVExfgmCSxCX2bZJJt/h7J0ZCRPCSj9m1
WwGyIvSPiS4KtyJzcB5D791GlM1SWqgOajgHecH5pU2YimjblwK71ZFr610+
SsAW0kT8yuRp9P+HJG2vOjttMk5s68Ggrm/6g9kNjjrsupJO+Pbb4fbMUecX
phYrpJchBa5rqKzsv5eKxbZpbZdHshwy59KJLA6V0pNPF0dlH7aX7ln2emHo
TxpA73xZiDj2KplItXivV69JSgJuJ0aeFNDHh8r0gAsOGP7VMtOt6FOWyTqL
K0XupuSqGR4Ob9Kt4ERpoWfJ/G90SIqErjlelC1/V8JI9FMSV4uW9xOzZ8kR
pDkK1xRSWhLEtfVkoSn9Rzw4HallyjsVIwk+yYTYJmsHQZONXYPcO5+f7EAV
AGDlLeFSV9rJzPP8IMWZIpusRO5+Uogoio5H6mfuBRsV2ZeFXuf9dQhU4NNH
gZtjhcQSambm/8cKze5sxh/GLLErH7EYUkf7/XyOjkDZA+XuzALgvQMUsLj7
GzUAj6erzvzzJJIhm84QL7GA5QJKaEiQ9tGdOyInWgMUKMB2woGt744ofU9X
MDOd8LfMPbl3x35UWLZ1Xu+5ZTv+b41tk7oUaPnQfwRdTaHdZ0awtFefY1M5
cCBoEkzoUiXKXw3zhL2TfQLFuSzOU+WMaRNN0awGAhEGwaNN6Q4xlz+k8pE8
2EMkUKYvArMYzIg37R3FGUaFCOdCmuHOkQ7kvMrVjtbdJpDF01/NyGCeAewg
aF8bfYkHCOFm7Noe2r+jjntx+E7GuvPcl9ITLq2ti+kBGIyfGRd4o5tCnHVT
8/phT6oMR+IJIZM0nlNXO8BKUH1u0d/fzThMHQuIBbtQnSqFysOLvwpaOlrD
lvKN+7fqTdXqws/EgH44/M3lEG29YaJJIbFRvmQ6SSe8ZB6SGdLl5G5r0xsR
V/H6xBiHEf05aBZXTi6j/jFZX97nEcrhLbKfNh+iv7s8Wtyy11nAh+aaTVVt
r7tKBQU8Y+HyhNNjy9lc0mVTSZDmaEd+THA6TnrdTMrIX5tD2NZSMUzbfk5M
ZKYPQPTmjz/g5l6tXmBcf54Kx3A5SKlQVT2EKAT4WYLHE+9TaQfMjcmMc9wl
KlcI0MHm0zmsmdC8aC6V9OTH5dY/2vhogk/hw8qwN1YCO1OhUIXj/7D6RPUz
XUFD40gGSq9Oonlb9deEv3VPYCgbGOitiP2/dSaPqx1aZMUizRg/gdBbxKaL
i+g44pGmTAfa86eDYKzjD4/xiObfUockyaPZQ6FhFTg0/YrsZhIGrTOkfaE6
othYnBl1P/CgfdBtEljBm7Hr6hRdQz8Lwy35XVK96+5uCMhn4BhcO7RMRNDN
I5eU4ZGFG0+fivhi19QAkgHctPdzu9Zqk7E4W+pMzSx9LnVuTjuzSrUDLw/M
MT0IUJ2JfM8LdGGsCu0+gXSckpa7Ds76X+Mj2JXhtptirTFfmdNQDw/uangR
G7khYAX5X2uCpvxBGufNodhbbQ+bRld3Dbvsfwy3oZ5mxtjoifNiyrlKxHwb
OtpZAuoaeJSLcvYDmO9tW4VmqWEWoZuOo0back9JJK4WMerpLBfDeocElwdC
eQk7oXrMAiweSpKi6NGAK1l9rQ+OMqfZGfuP+RIeP/0R3SxNa9tZmpq/eJc8
mOJcA2pff1bIV/9l4zcL+/MiAm/iwEySwouVSAUQkY07Wd0/b/eHA+QXq71n
KYoZTohdahAZI/mCCeVvskXInRlwD0A3icgDxfr8AVQMlOB2671Qa5p2i3nA
0nGu0jl55COksEHHPBWfV0RJIb7pQfzYeG3t9OOriiRLYCX+y+YtidJFqPNI
H3IjUmKFLWyDn+obVC8c/7bqdT9e91genvy3qHrcMZbOn42coyW5tnvXC2C2
9gHcICKm2xfAjHiVJid4fjLQp5L4jxDG6VFmRR1eMlzciNo48q2BmrL+R/C+
oP7PrVXKkqa+/AmJnTbwsF0ZBfWBMRxxwuxS0Nadf+ajxUWuVnJp/fdoNNpz
vmFHifJZPvLGW/JMlmtqg5TcXGtb9YeaUtBC/fBGozOZ4ZsPLoMjrdEIDZrM
AO2zTVRfz7Fr1BJ2rA4VewdrIr6kiaXGyVz+cqD7ryrzNRnfNcrr1st0bDbv
4UDI5FM1RcvWt2I3iOhgroh1HCgp0GxJC2lRfxdoAcnuwUR7o2XQj22n67+r
GlIgmo4p2Lz0/NqZwOq40cC18Y1+08BHFJe72VpAcQYgEnAfv6cxy24+LPsb
6V/CQCox3w2+yDDfCGnio/MCdN36UBqdnPgZe6NEOCBkkKWrFrFadajRgHsL
q5KkZQLivpRM49ev0ZGHVhTzsFkhN+XhJMVI+fK3T8UsxjkOsVKD/02J5hwo
eaHlN55FdxGvxTmIrciSUnfNAgZLwPyXeRjBLYVWXi5CA+w2RQ5Es5Q4PFjn
7Pn7qFzvo+0fbiFl7SjVe4FPCpIwagQoGkAMUODROyzs/ruk30QCxADxUk0t
lhgLyrJGIGaF88JLA+65pbdzMeQmog0Pi9LLcntq+fPtqbaCgyF9MUh2YNOe
o+zB2KO62naWEI7cC3Lkxa44mz+yuSoIpfpz9CQNhtrD4c+Br4RAfSzgMepW
hGzwUwDSfvkgmvpx7sTDzeeZf4kdeXPXcyvcG/IM8+5y3B3KH4eoyvpWraZB
LhfVYmL2Tv8bs9l76jbFmgJu2chudLX5cGBOT4x2oj86sQge4M7QBJOhJPf5
01uMeodfBhVfjhZG1Z0LlCjqdAZzEIgJK+5Dem31zRtdAfmpAjIznMsp7etx
8vhdjnEB+Gi7EsQSvJ25NvUFsHbVqnv4QLHGX8U+SQZoiqPoymS4yUk8+J7l
20/cDbKHaLlRS4QX0a2CKFxYa5fGmxdZwGXMfPMw502LbgOSU/HSvqeIjvoy
ZHZQxduq5CwnP0DttRn4EP+EUBqZW0xuf0F+PQKTVa8oRKoWCmp7aanuhHts
ybutZmlR/CHK4rgSM0o/ae+3ZhKIjgvlgnQvV5nniAiPAHQ184i2xgr63gRX
SIu0JEpxoeWbc8L1e+qMmMlYexz76mNlOFKKbFGAWP678uN95sgKoJWfq1Jr
2WgN/o1otqrIS7k3rtopGqY1uTEsn6ydKf46226zEVK1P+xrBwuolfoAz+JU
CCpdakAhMzJGk3VK6NXnNBqIgGYzn5Bqs/zIY/CzzE5qf1IAkTRJiKr1LDvT
jNd5x9/KnWwFDx4fTiNZ61e/avpZnkEUnC5qWqAsqvgXZumhzWpIfka5qWd2
kFOl/6jfDRnjrywt747Bzt+TYcd8KexJOIlAIn8OhFzS03Eb2oiwJCduV/C7
Jp6aGBrlf7H+caqbWCYoyYx6UW2XZdKIKdRdfveiqgdE48pgR2nao+HOACIY
n4eo44cnOZ2HhRLQkDQmkJMwcjNrfaY7ccwiHYdJDUHBt7rXsKB0ryQf+v17
K9w+D98tEWhujKVK4Zytrwa8SzqrdB3XvUkASVGUQ9uB/mWXBdR7tcQbqKRd
oiGFrQQ0eajGSvx87Km4FwyctiukCjBySqz5N/54Ee0kC+rqHAkS5nz1eMWJ
Glc9qGf0j4KNCaxglHjsCuv3QeCLT5QvsXNrGPjXIGpO1+COP3etvWvI+M8u
oTV5Wnl2CgvcPKsqTOmxwD6HNngBLei97YpagFRGaJhuU81hs0h8mbKc8NYl
BmEIUFhpGB2zRzKXty3whx9+YTMMigXAMjvu6mF+EHZNF+6AHwd948KZiBRp
sPRd+nYStLr7VyzWI89YnXYsApoln6hK7tr3Q3cqBSJKdbEuN14wyK3mtHuC
TWVLCDkJzW1le3eOby6QaUt+MC7ryT7tN6i7iAQDCOBJH8XfYXqBxKcKB0cH
sz5sBhNxuYToQVqz7Fn5PAQqzF/xYuP0DzxffYuHOP6TX6Ethi8rH/alti0a
z6XKD+Re0VIlGRqvq/i51qTd+OpJoSUDitnG/X/fA077agMUriIbm85eNPQd
ADEFmlxdbPPG0hOPMonpZUaOiosDovY3M2RJNuh9QXbUlPtPntBI0aXZ/Nnz
DExyoBUU7CKMi9DAdoPLZug+wlnlDtoy5GsDS4e9D6JoVtNXmuqPtl9fM+kr
clZbq902pEl7XV+vfrbxAyZ/rugIk9WWX66DYpmF75lEll+TzNXmCvHNAgdU
MsxiA9s1fEUmMRbOyDzaYtlL4Csq1UE49x5HJAd+5ajn0hnd7x4NETzhBbIT
Ni3LCbRgaUUvXsD1Eqla+FDxJqfN4ongaCbWATv6XpBnILXT5EBMeIzZq/wP
vTbnUs+ffWv53bDT228Lugmq9HIPKpAFe6Rf7zv1CEm/ZO3ZcWwoYjm+Pt2S
3KoVhw7t59Nf0GXbWDSor1jfue4ZrBfkCyELvaS0k6e+RVxYw00n2hOW2fgj
xLAhOKG2J7AKfJSE0YvhuwDS7PB5aQbKAZZvb1coHa95K6zemKS0uzbc2/4E
+unnDZpmcUAW9iCBmSLHrTQrmlPxwRq+S7w4ABlseiDD2Zq1BPz5//jaKQqb
6G8AKVtQRCW1ctxuHYqpxueIPtUIMArxOnPX4922ITS4Y138LMBTYhwbeQmf
1Kc8m4ONFrnfa58pNte3WV/UCx4dIfvA9DAt0kBtVlUE8LRm5Vcp8xVcU7We
mR5pJ9gP9zgfFN9smkFGeY3mYl+wlsE+xaIQsQCt03NIVb96wBghVWLEl7rL
pVWKmzCGVEQKMjOOQkX1hmKngp3/ud0afGO2AW0m689LsJL7Td6Da1C6D8ra
vLdfnVas/OYr8TN+cg6NbzDemW0bxU/KjT1hhmzxt9fQNOKJMz/iLNumKqRb
YL4WzaFZvUs71q/ZHtCFTXLEEJhgrRx3uP1J8UxQ86p6lF7C6M0PEUBcJkLL
mx45unNxSx4E6Jui5C19i+vgXbkEbolRRvQDQH9+/7bRCUh69HElv0WfVuhL
retquDAjoU1soL+jeic1iY0ft0TQ+8IOAnnXSSGUc5rVcrRG6bjJqSMnT8Bt
DNJdkorNX/UL85kHaF4G3sjev2Nk88OaIjwpCeLzbbwv/xjqxbJb4k9uwVEk
XFcyu/f5dQfQeV9OnVzcHxc6scuZNg3i32JNAQVtHxThynr+DmVaB/C+fh2G
FxyLAk6W4Kbtea8bEtX9WVLKEzYZcepMdNSXd92OxINvL96AoCxvkQkgDkQP
db2TA3qGB86gN/DxHjUJBdhegMAo0zzzTsExYVW0G1GVqUCeViV9ht7RhsLL
oNRwS6IQqykU7SAtn2Lyk7cKvka6xZxpebKvJniDnQR5az94G62+3u9bHU6X
K9aj9hJ5LYqWMDgPoWaLUefIyBaFt4B2QT13kZUKkSuAuZYdIWN7SYkOzgN4
ufhCSrElB3+Clvr67XszpKQJvQ0MeXjzzDXLPA/aJ7lACnK/J8BXEkanBlsn
dKBuIdJBb89k/40PT6NuOj/zkk3dJ7gy1Jr/6D2pcDCUY9Z8Olscawt+w+pL
p1eJj+IcmKEtCVRXaJkRXMJWy6FuszHux8Mshbjc0wyKLHrRlR9/SHVp/CKN
CYG+EOzmX7WnA5WRiKoLPkbJB1WDnzHNatX7S34DRlC8SZZsRFO3xJEhFZiw
Ats+4QdAvUFzGNARwBcj9fXEwgnxIf5CoGCRpHDeF08uIKqsPdnEyWfLB/vc
e2miPtuUz5M11XWQb812gdeTu113h3YXoEcs3c1AReIr1viU36M9WYUgZ39w
RBxpJQvHtkE6I/zBsterOHbZAjy+XXCH7+ZPv1liOtDOdLGO0tbvfh57uXrk
aBXAtCr7lTxS4hiGIwE+bR3CEOHSbcmTYJiO3WFu8OdkaLZoEKHiVhP1kH2H
reB0UWMHwEwPhIDAm2pIz9j9IioSYe7PJJEaiio6p5riH9F7uURNnb6pni8g
MzYBho/2Btl/C6YefXLJiDbafO4HN7sap59e2pJznYr7q2qFKrNH5Uew+MJm
E8xQ7m/ZcCiwjYaIHGUOGYJ8XgxLukJxmRiivCCai3JzbX560ZMy9QcbR+s3
P/Bk66tpy+B7Uss23aJFX+fTGQYFAjqjh5RNqWDXaqVmC8bf4AEbgqcS4bKY
lsnD5k1ZXCKQAvBYZIrMsU2FMYo9oi5rRwthfzq7Ifg9EMeJwfLlHMF8HjM/
a5dzkujj4NhiKXBcXl5w/YAcnwFQtQlagIwjuC2lDHXm9Lb5riTql6KALT2u
UZnCbL43zkrQ2qCUjJGGdWKmlNkhO+iOpw6K+TZ1VeAmmbCB9ZHko8BQ8qVr
JwwgZS/w7NOg2r9V5CpTA4E0SvsqjJA0CESG0qJG9puqmopAyObr9orAp7Me
ro0sUiW6oGdIqCFs3F0qwRHdqlKAYedbZZEm6BpEaZT5kTRHAuCvlieDO9LV
wNqmyoh287uxYJA/xvWWXHXS0EAcH4YWNH+zQjCI+lWK8xrIlJ8fhmvLQYAx
6T1C2Zlx/BPzkvXKRHN9awX457caq6d80g0GAFH+u/+EeqQSx+yAgb1GuQvT
yfLBQewia5DqZEOsPVoQ0Y37AGQlU5t3frUVAyXaQaYn6BmEAj/3UQQi1zNG
HKNEj6BtH7CG74l46UEHhKLt01VKQ23SahQLDZUV5L2sxwjKG0mUqHo32Y6l
hYm+pEfy/6J+xhzCrsiGrF6Q6TPmHdAD9MYRwtaq+Mi28pngEJbgA/1PmPGk
cKgaBFNhmRBeQaHCmshk3A0yk8dShHuV0PjXNM8b/GpJ5oJSOkk2pak+fwWX
3b64bhdsRy1Hf3hq4IPcRB4juZYM7jRW8bPVL0p9GGciJc+3akcNzDGEWMlY
G1Wv50cMHNkG5D3EWU1vMm0RCQHiYitHznmxXcGzIiq0K8hnAXJ0Nj2PSGLH
3zMOzjvtdVrPbqPRlzKSXwgeZrTiY5rqrMWqy5j9TAmEAOK7GGUtw3+p5YxW
3dspLfZVpejquwL4fFx6Bg96IY7wsuYUoXFdvB1nrM/YRIZ7yrrVW4RFkGpf
RGfNG47hP1P5QcNLIjKuCC5AwHOosw54/Id+z3v1lpOel94A3yV6vU6Q2mvL
BttCM3ox3khtED+1AMLjdn3hby5nYkjZokJH5Sd2pSZ7xPXyDglOxX5uxcyc
0MTv4NY5zAp7FhZ8N6DNYf232Lrtxjv/zSUwpqv2s1rHoDDO+z09BOaeMtrH
iKUIEKXqzRvOppubZEyEF+H/Ph6gHo3frDSYG0JFmn+FLVDKlRiahKceacXv
zAsJOZOHmAthVXxwyak2AbGNoQBc2PME3nUx1HB1ODO7rP7F7kYiQ2CgTgpq
bp+SUAPYVfOb8KnsSMPx3LNeXPi6KCBXBlJ4XAmX4mEHfhU3rddn0xXt+w04
9V6nOs4EEZc7iVACp+Jp++3xWtPafuFP/Mi3RzuvODN5Mn5EWQDw2nicSExk
7iCRUW5AZ5EHovWpcf5P/5IqbHQKX56cHWlXC1o+GDYH/88cvSu8xjueLLxY
rnFP4VYnM1zhgcJmI6YCrOUu2i+kLMQ4Zv5vUkdZlTlIxirf5xYNQmenwFSR
rP6z92jFk/K7kNYSgEQiRRida15QnX5eLDJpQhggnei5PqfwQyDznGD72DbF
diS+Okg4zCbxGtE3gooxoIWaOqL2oY9qL8BKmw7/SUlj4vIK9SFXfDqHKDtU
+WGFJ0rlaO/b8EoVOjS5cYC6MQI7OwmjRNQZwLMe7lAOzhqeWP4/VmhoUXv+
Ts/gz3SnB6kQTh+00bDMaQ9zcDiW8N57HxegcxtE/64sAaDSbULz8rPirrPT
aU+ViscyuznmJ4JOrGpBgiGEjsarMRivqlru1RXunWEtxns/QCFvCE2TX5br
HlrCEXnfFp/g+QswU0s76Yta8XFBetDcXskTxagAyZwTWCYMdkxlhCZcnuVv
ZSptgBWViT6BnElMo5kfxmhrbzUghgLnhOHqVuRugyOMfZJoTI5cptCrqrUA
krMilofCEFWtOB3r4jRPqZETcyHHFc7egH+NBgAcRcaPxzajn3GdSax21NYp
PidwSdSgzNXBqoaIrSEwVC3K+5DfUj78KpaYPLIhTP4XaQRfQY3jgfq6AjNA
3fcm0GVmeDtnhvxR3l1gwVVkslSMT93Nc/5MktiQ8GPfVCSDbHoU/ni7cphG
cisspbsRU2NbOxZjSI0VKn6HsuxMYEbD8h4A5pq3p99AjW0ggRd4vILTjdfG
clO1yn6t23bl7fkWZ4dc85aHLGQdAHWtTvwFxz17HB6nFubKNcFzit1lVBS1
g/L/mhKqt+TQC9r+uhFhYBKssslyclpkvuuuXMG3KHKanVvjVXbEZ60uHLHj
rUrfb5XT7Bracr41Y2aVLM3wLCXd/gNTNQm0XYoS1hC2KvcZoe+4+LG9iIvV
HXl19to0UY5dEeqtbBdrPIoFhYDzqlel35GGjV/y3nBH4PmEXq16olqX76lt
kvBW4y2LwUmLSLFtTCjI0Rg61uJP/rspkNHzaKDjJ5a5MwLsXlZ4vaSxePvB
xolfjrhNUbhKtlB5OMwNotnZEJEMVgQoAPC1c4dOUh4eHJdo+Z7YGdu3Zfhf
wd1dmuwy6WrdiXxeS+2bulqwIyxT0Mdt4Ibu5/LiEA2aYK/Xt98xL6vHNf3M
x16EgXdlDr9QKhU588GTGz8g2/ICyAOTHatYQsYYoC6sUG4rh/MQ7TCPwGMs
9zNUD/hy9BMd5hYqgX3xbEKbqfR4hEVzB5cPJp1WkxJRX2aMflzgavhRVhXy
jzLMq85v9z7B1O1WX25ekrdCwGnua0bSh4wuJ9mAJAY0b7tc2p9omgVo+1gF
0mMnErtYKJ5anJjchz8B92Yh3fMC8JZGMDUjj5rLwENC3bJO+2PPIMzfF7xN
dU/cEOWAtoR0Y87FcavWOt7oSaIVAbrAC0RmLVZvyj0qfM6yvcqN6/cF0Iti
55z2LxVyiv/bhYBByZr31zeYhI3CBv2qLmL44KdWtoJpisMfbe5Hpju4Hh2b
PEqvk/c5AjtIRTUW8fUDX0GnnlTHBUimOFfmPQ+3GKHCkHA4VkFHfNXjYjxK
IH4kyEdFqZu+PuawMn7b3bhmm3oNlY8Y0smsi+QPS/nEejt05hpVSd4BDKpo
jYJWJ/V+RN4WI908CB9TCncyvfDnhqTv1jztGDp8vy2kw/y7fUmx0UYkNi5q
KMSb3Ios5++tTMEyrMuX5E0kU66SMSGilyfYrwnQctL3cefBAAPBgWlu9oiW
3KPQ+Wmw9w2gnkCwgTvG4v6/8dXFJ5EhUwvCFz/cS6zOtFF+X3RwIazteDXy
HYZoTl+sGxVCgnvG/ky2QrcymrGJVS+xgjHrmek8enx5/t9NN9/IANI+wVnC
NUPDMtwDZ5ZPemoKMfbmdSyelVZNphLW5uBv3+GgpH/Mo6A5trKIbFILnr29
XgcCIZRKXtykWRj7NMubfZSsbgcohOeXSIMraoozmjFDPsLx5Ryumzwnw2VQ
1tUE2vUN/Z89s9N+8kkkt8p3xHgF4kQtvyTa5dD5DwzmuqAcut/PvZiTtjSU
8JVKGtHWXHX5c9XEFCDRW2NijaOY//WEJc1n6VC1oQNGWi3/4yK1GumvsQbU
PvMpmaoTzH1tQxTcYXWKEg8qaNlC7S0HbCPdgSEDsTY+1G8Jvp3uLJ0T3POm
InROcuIoG8oh1/anmnulBuZz9TOrYmYlH3Ed9Jx9F9XgPs9boKEyRFoveJ7h
R6ifPRYZ9bFgPUqXUMMx7MWXNZmxO9yLwuYuqEJY6ukw+9QLif/Ej3O37L9o
SeiHz5mMnad0SD6MIJblmeo8WwXMxO7w0VFKlSi+0FU43XI+fNtUYeYdvnwX
X8gLhu2w3kGn4EF9qoSoDPK66FE0zAQDCAXox3hFWeGzL1rhpZPMaRFGA2bX
HTNCV//iOd/dP+k50UL3IBN0n/wDgzsrg0cIP2Oi3jKPw9TAZCeDvRif8EN0
88FnsIsWivOrK0ge5zKPNtHOn1WPP5ylkqmxcnvSZrplGasI+lzPQrRmhN5R
uC/W4hCOyP40IV5oBZcH4bu77qz0uEJ7JWtcL9JZT3oYVGDuogIcQqyh09Mz
usrmGBdHLX/rS+IqKRIBnz7VPXF9hkGsUEQdjS7Lb7PDn2GSk3zL8dbKwW0q
C2T6IZLC39s6pigjN0wXOZfZ7tEkzkLqHpp3ptbkJfTdBzxZFgSn1SF/Y3CS
bzSyg8kCIZgBzgc9PGF5dEhrrRHeo53LfBnwC2Au4YfQ84VQNnCbhAiDze2h
PV8QZtjmRAyxzrPSgJ8ixctM2vgyvP/vLtgkCFiGQlbcIVu/E5P83kxi1YY3
CJFkSDHFkQk0lHR3/Eg/XLIkQDsKVndb/I1JUxjdBwopYXpbT4Hu0ZMaDlFT
PV1xuwyTote/IhZ8VvnStfroTj1r5lEzfTHP6QCDB8ZexGmo2mPEsB3ekUNJ
EHHw77LNY7jrUHpQK8kiSTsjh0BwLH3XD5Pr4Cs6QB6JCC32kDeu/RRxDSSp
oh8ElEPaocyL1Q7Wn7m6pGb7FOSy4i8ZFKrhiSy+XXF0UReYDmY6VrQpjnXk
BpG7gKYkAjrElUuKt09LwgIRg/KrwXZCJNyBKJlqGUOs2rUkpCGkoafmDDNI
BV6R5wqRg92uaDfZVXOJn6a8R5MIn7Q7at0aWPJi251XwW4LOKuKP2Oeh7qC
D4kILxcUrkca8An+VJ+aBVHQMWeO6k/pNUAKaDGrU+68S5UPABquc8FW6S1b
NB8+sVQL6ed5bCFIMaSReXgQZhZeC2Rxo8h6s7nZkL3kn9oiG6Oi45wpRovS
dmHWpdxUkN1ckQegCSS/XFXyFssjmFWfRvw17vpASeqf03fhnqL78bSehKQx
u4QIG2Bea5YqzX3JlVGEoCAEjvj5BDgjLLIaSIisLn7B8VbFtFupcER4ruJY
Fo4XnOoBIy+947WSg08lOKQeOCcnrR/q3D1P757709u/+Ju9ik+kt1Mr613f
kvMnk/DNtifIBHMgN/s6+hCtlOPMEQ7T3gYhJZD9ohVfyynlh1hLrqZn1HX1
A5vZxhYXvKHWHAIbkRJELSDGR5SnI9NbCyzP5bJ/jOdQv5kqXStW7EkyoHXG
P8IrdB6Fxhm5rmzjw+gL8M3gzktssEMB84//Pnmqfvsgvc1Aapz66Ow9qQoC
UTN2jh/EwcBj9GY8pK08fXrtUZEMM6mleFOmqCMqBHwPFMb5/XiGKkahlXbH
ChcZ3N8JVdM2G12087yHXyGtpAmKNr5E/UCzQRj5GxIqLB3l8Fco2g5wHr/X
qDXkkT9uIC4qKYYKvODJUdD6V+czxqfw+YpQN7GjzV1pH3tqJbnL4+LoM5IY
+7wOMLMAHoKh1LFvoW25BjhnlRazWWhOTVuuhOY+AW9yO68mTR6FWS14Sv22
eHvPzxdVpAxgQTf5Qnl27fQUosMJqkVRgwF05xvE9963hB1yJ0xBU7Rs0HqS
uvr+eCO8fMpYNvsJRxr9d7FGxq7KT57/AUvoP8Dk+o2QBn38xpkL0BtO+OnE
/YL+Riaeu8C2M/+nk8ciMQVSgu+8L/knRJKoFM97Stb6KD7JIQ2L5nJyMez7
9x1vN7YB8sKpAohKwJ7GVYHsrngD53jQrxOhhfVGF1Ps7iXW9LSZppRScABD
geNMTiaxvUTCHdG0bNVqv3Lentegpd9+W1e+zrLIKyv5JY/XMGi2cjkQ++qV
Le2TbXkPMCyy48+vkXaWR5u/aKMyn7gsjXV6GFx4C0J3acnjnLpUhXe/iuJZ
a12xHXC43W/B/htNj7OVNjZcNtJDBjEbetd0SNCjWdZCB55XsHpKR9IpYlWw
MCqXXpzIR+VrEQPEkI9lv9jM8gjj6qaHgB7/gnJfV5RJuJ0ynYTrjZDNUxxr
NIw+d3o8av9WwdWMNKV6cl/iM/aG9a4r7gka6BjzhdpYa9PAzBWLdEApsGVq
fKIMcCvMS70iBeey2DJqFpRdx9a31B9IDdufOoqEZ34zXR25rX2lBqdCD7tX
EaPiMc+DGyLSVJjWufmUaRsqSRtviqEzJ6U/mEEpObTwZOaxRn525Dp/BR+C
co0R5PNRtRHRxV2WoBsEqggTbL3Y40N8oWbDnSCqQHVnXOcqLSPl5An8RU4A
MOvhgPZXM1FSNL2O7ouVTT3lEQeV4eKl5ui6YVLLU+bYKIXr32yTMeKpSsPD
L1PcMerYrOX6ndda4xk+8MviWJUiblk2eiI19KhmOey2aQ1ttghbWaeXuqoe
2fuDVbciI3WQZ71D4fYEYxPRm1YN5H2RwjiGq0AUe8axTXSE4XIxNWR+j4h9
MDOHADC1bm/1fJaExQop2E8ioBD3UMuvGGXY+CCRTmNwgFw6S4ArK5FCiUYR
ou4ldA/RezHTXw842He3XOZj/hW8K6hNluXJOd/JrIwKDDuo/r2f/eAsGHc8
q23cIyY7ax25uEdAx7r0Aiinw7p5yOecS0jnPOZCuYufa8Hzcrikqudb/Bm2
/58m5mWfnN4PaYzinD5FPB28Vjb/WsinSzC50xD7m3bn4I161qy6uv/r+raZ
BCty0nrl2757XgsbFfiZykYrLlhNfD0RMFe1N8SBkYKXCvJFQY4zNPVg/Qbd
Rwp/eppA2zIvKDcm5SvZuWGB+O/kBN1/ONNYSspbkfMdmqmQwYaDMqMH1Iqd
pfptOkoXeFsd8YXmCrl22MMduRZfXg0ptrV3KwA7u6SIuSQ3blg9/y5zG621
wFJIIUuh9YULq2itxwP+OK21kUYUtm22eu1ViR5z40Y4ED+Ep7dSCE9MGN4P
vm6ZEkl95ZWvJURcbJ2C+TigVMRJ/1FdbWHmFcLhpvTOADo8vkZKwME6UCLB
uke9Alpe9O/AknP8l92PV50dk1bZKqeIH4FtKo2YJLm3QdyzExRjS9VEecm1
p8b4TjaujsMPkT/nlB7Lo83JjRDThYmgAcZAsGRLF7rGpXBbvVbjfjYxYU8a
kZRRqgiyqI8ELSw1DIMHvHVzttA9ySK6gkwr9OS8s05Qufhz9HFn/btDQC5Z
dr7QiT70TwUsewmDIkH39+rnmhk1DJMRv+sz8bprheGLXFBeAwCTq8rWVO6q
lXrHO/fKj6VVYWXNQiyklR+ewvbA/MfggoiZx1P3AP08JvdiArku9zkbwkHM
1xXKfmiIDNoXeXm0gvGLd2j1jxyVqEl3pNrv2ZLq6ZnLcujyTQD1q48mi1wv
KDairw8S560f0qdEjRh2xeYj8zABnnT2hmYbzheIuISlD4NJSg4k1FDAE0gI
U80bTxTq/a5XPSOLQFUVJngIXuxdIcl3T7FURhl2oSLnSnrUCbekruV68lU+
6nwqE0lEhP7INcFOXe31QCrokm3mzXMOz4YsrIDuKWLbHb8HnXlzolfkqNLL
ndrKWOx+0Eb6QZk8d1yAKHnC7K4t0vK9jh7AJTT8NRYZ1eBKSM6wj+oiu4JW
beW9zVQ7xVjWRs5r6r9zSa0xZjx1Bn9Gxu2RxI7/vqIEQfkSiiGD4AD9um48
2W3GcgusMYk0lFE/ml+gUShPA7JNYL8RKJbba5u/1HIHTV2v6jYqL9AvoFGV
VXx5LpJcUAQOouGCISZxAOSw1b9eSg63xnrxAxah6N26LAK2tRq2CHn6DaQg
UtDVK7f0Vfy2czPo208yTTJKPVwGwzaCgX/fr8+QLZdHZ+IS5lmbbi6f1j9E
JrqXNcBY/iDF7ZXDtM0+69DrkA1R5ayu90VGbcP1+KUo/33xP7HSIsvbOf17
ABmwVIarAIp7pNK5TKnize+DHfVROPLx/6PV395gwu8lmKb3UQUvr7OeZWgN
7rOree3xTJ7UgRzB38OuT8hUh6/DpLyykUdhZziGzq1LmgCz+2F/uF4EYNty
BcL0QqXICSH3g1Uws0fkCRmkJqWfhWwXV5XrpnFJ4InOrl9ZK+pyq+jBbfll
Pi5mbTqVbpOG0r8TolhsM0El9QDHk+H5Wu+ck2xqFXMBl77n7llAxhwvAvZw
RJW2MUEunbTuSZBiPZNInBsbdvz4ruYAD8QK1+yPNtRYPgOKLqAwdxahZDcI
c2Ga4YID6i9P61JI1++VfPjMX5Rq8LpHfJTsNhISmiZvtJhUoTotzYkx5xM+
iaXgEF7wIrH/319bSzeNY0Ejx09wscIFpsVSFmyKevcJE780bBaReQuhKsv/
s2BPyZ5ukOwPHFV7dfufJGHne1Oox2XuCLnhpvvkcyVLeuEmnF0AGRA3Qp2n
9ACwNnouVTn9H1Fa6z37gVIVyJCkNnj3/aMgPc5HY3yDGYjkC2hZACSsY4xf
F9q5bjjmVQ3k23ixCDQ7VEtI7szqGpLzmWizpmInL8m1JfIQP3pf3QsxA3ZG
h0EcECYWlLx1tqgdbhlvx8r0gZCgXCKGnTiGUmzKLTNvMft8ELF9D8tzVVd1
fLed1gZNXYh3epX5UlczfNnaLLJLIr5/va+Iqrnf45ERh/MYJI6YeFrjWW2L
Fo9U61hW+BgBqthLtR5tJYV6mZqNps0dRUX+Wm3crXDXZr8JCm6vmeKjqOfV
5UjiY/m5F0+7NW7gVTStIRm7xI0LMW1Ot0vhsdJG8t7mqxpqPj8Oxg9ciRGr
yqR/od5Llxf7eTqbZDFJPGHaoeKorByw00rPcbZ7KLTCg7gFV1xZ6qG/Fe2c
WzIbilAKDPEvX0qjZtljr2UyiLz4/06pmarVRlsdm9jxgxNfBSkCWj3Q2cHJ
+C5a2wF+NmbV8tK3tvkGeOJ0nechHUJF7qYC17uM40kXJWg2rpEwqwzg73Ly
mg3yTGUw2ydofblenTxCdCYsedAuWaPWowDmjYiiKwxnqYz7Tv09mdaY9nQ2
aqe90p1f3+/nXo22VGrwUm79L8m7ZzK5aBPqmuDObJjGbXHHY6C30uVOsDXK
Pj4ee16f4o3tK+DRg31yMW6WuJuoE9LvQzLYwgbNfJwcGv6A83iVIYGjV6bf
RBkEyfxa/kF1AYQSnlB0i6P3ZRF5/rKf/MlQwF4NmPr/fhRGI//q8qus2KY4
ZWOg8ASdbUbqqAI4eRK9j1KLAgSJn46ydTwKUMk8UvG6OMXBFb7CZp8i7kcy
ERLeK2YZHlFpJTIVJ8RRJH3bbBdlSEiOL4oxGgd/FBy40o3siVqKSohm5FKw
U6btDCT0aLlwWv2LDprEFw7LEfYGi96VaVzdOsYEYhFBLgjbG56taIjUGGLr
NJNAMlysD2dr1608i4kO8kFarXMI3KtoyKhckxDDAgYMJTcOY5xVY+5qRkSN
reagAwbuQB/5BD/VOZozEUlrB8/Rx3i7oPnUR2jAYC3sv/qUWFdLIbUPQ6O+
8QuS9+PqdifrPIOBkwnipYRk/WxM0wxiQN1+//Zt2QKkddma+MSlBNinr0R+
9kD8Jx6JMdmt9A0ivg3c0xssCNYhHQ7jkmHc6ySpwEOFVxWZzuIZCkZ+7UCM
ZcsK5liy7CIhZLJMvxmUyTPDjytil8vKEr1wUptECX60WpX33r9qwoFqOASV
IDlf9001k4lAp35dtISidpC5rF+II5nh1yz5jsWXaGtHdWSai4EFN7l+R9Dc
bXJOwg+ygh52ipF6Omesdp6IBPl8+zhQ/Ld5ITYVFkL35CVseGaf4l58dcKU
EDPsQ9/7pDXP35CAuOyZUh+D5ukR44otjfr5FzRBFE4Q5mjiYLBM/tIBMCwJ
gnbjNUgTqihqRodGBI0hI2qjQZ+8HeZxSj1qUjPZ77FrdsiiE1rzuaRcZXL1
B4fXcEDnS07hB4spAJYyKpaLAHEJVTHRWSKJM8T7vej2ldt1rvjhwYbEUoYv
6CsNr2zm22vqn3/73J9gzp7YscemLyEuFFVM01yLbLpumRoMWyTI9pS+I3pk
m2L5KzINW+QpURAimaBbYLr45kJU7Rd1DnkRBYPd8+NZtf9A4jXZl268zdOW
VyBQN7y1LVXyU3UUhvunFE+P61z5ISaV/pJLaYokvFutqB46yInmXlLexaGh
gHaTDVTmqOQm/tF+cOBO8ZN7b2dEcxrvCILSiHfxAS/GXEGSxL/ulgxOHeUX
wQtew+lhTU58KHlHDIWpwN/XHVvasBajQSO78x9HphuSEsW22T/EuFXQYH2u
T5HHmQq+e21antnwmM9bQ5grkKzIHO8Y4gOcaDJj33rJUh6KU5q+WXhQA0UV
pQ3Va45GYxtDtBUj8g6CjVkboCFWUF5+fOCyIKC28byIdnCgAw4WqHHovyHv
VU8hwiomTmoTr8yx9aHGN1rYWT/d3ubMATvfHb4F3HB4rKc4QggZ6CUiqsf1
akSnGtbsZl7QXJtMTN5ylPrg2VwnASJGVRQxFzu4DRScAlnvWf+iQvsNVqP/
XtyMgZ7SVOd0IboDGuUdMr1HT/bvD0nQwvdmLmd+kj2wuFXp/odORo3GcNP7
S5RcWusdrl4t1F2bGOz5X2RCzqLmjvWoc31yXCVdr1jGZFLAiGwxneoTKVyh
lODesSEBt2Ua/m+uENTqT2Rg+pOUf4FkeZKX7ykeTkVZ+395WG5ANCaauB0L
9QMcHgZDLKWeFkjT1tR/yHWTOQ4DLGglqeYS6wBEpBnJtd5ym/EU8dngSHrC
Feh57gKApeZdqQFbtdVmp6RVElWBmueKxt5OMqW9PUVozK21wfxlp+5zw9oJ
1xdNWPxxp/sq+MQdMG6nz/EWc7VsrRaQ41NpSfgBWCC2ibNj5gZHtZGqJUnl
95QbsHF2O3pDKOJ88JmwulEdAoDuuz2XKMeXDDJa2JdCnR1eYVhFIIdo2Oe3
vyGMxXlpO9Zcdb+ARMH96TkRiBuZQxzPO84kbHoDjc5ylThRWYNuHXoSl6Mf
820TBw0In8CArSV9V1oJvCWoCT5VSOGispKlJAjw//0T4S3qnWLu/qhWOidr
AwmxQnxlPxilc4W53kAQsGlqscQeDujdY6WATGMp6VEwn3NwZ3Y7RHAuO0Yx
uGyfBLE8+Qz2go+bKQyDSUsaa2+RCvZbWR69jV9fyawq6eg5KH4AsDlh5b50
ENrO+uSa2UObuAndJcz8Z0485u1VUR43ABJOZ866dPErmRcMXyGwTwyg5EEF
6wn35FowW1GtntwciJBb3xCjc3YgMbp9zG5B/0aZkR12UkKvBIa9LQUyo/5o
a1v+g6kaAg3sQgEzbKOPnPKgooPapIaeh7/KOE8D91JVGgPGLr3Ty/6seMqz
djDCYhDeCuw9bxTtSv6EcjivOCCiZAqZsFE1J7I657hvCB2qO0XnMvaiMVmX
aThQciGLvg0P+VECLnyvlfgYi/JwGbfIhKkZ68C8S3oOEk+4WnJT6dD+jif8
WD7sQiAJ5hOyOEWlZUIWwXpXcJjHqjHmO98ahee6+d1xCHq7nLq/fheNvTCK
lLRDvqTw9WelxnBJwiFhGZxt4AfM0X91BixG2mG84tR/RyQE+TEbGmacPoJZ
wfsNdcJEdcmREX02KBQSw01pijzdmxX6QVUqEBQEAKyxAaFGUSvOYKV7uLou
X4gIFiJnhpaS3KMY/Ur15VgBt9FKxphSO13sTs2q5ZPzTangNDGGXKKH0OfK
hjl4aF2X2NsJCKd9458X4+FhhL3ka0pZwi6Zl0Yc6Gmq1naghb1f8/fApkbn
71zbvW5tUn/rxl1xWRUcwiStsQOYChPdTdgB1yqbgmd/+KTIW9rrFaXJ1IYp
0hztHkgIn83t3zr/c+NXfWEHs1rurcGhlC9jy96yA3K4qiSafgMiv71cyuYH
bhooXpNM/knv9cB1JL/i53ZXPONxloMq8/nuEtKOf4pWNd9Rv2RKwnijL3pI
pBBoGZaJzzXlpwzaZ6LlYf1LQXvU0tLLf8Qgnd48HJy37+qqU7+iuet/noWo
kV1vinmKgu0xCyT/kDtjh91axr6o9b+u+VMeePw9i/kZUObrtuPMhIbFUM4w
ZjSJ2d9Q+uca4SPfnfrccjocI+1mipnILcN6r6E+PoOMZO3XGqZ19jwhN6zQ
inqWu6ywI9XyB3zlE9Xflyd2j2Uh4e+0hTV3x4gT3Z/yvZuUEyXhPk0dFEin
Lt0vuAnFkiFpYB13wMFCWbnr5dChZy2qoAMFR8bFai5GJnSMw80QK2dMfJhU
JhDbz7MsDg5Z+NQIbLaROijW1mK7tdIdD/PNslE64bMl4lHSf4VDue1BN9NV
zhfmPIVGF0iPW1wrnZ4sw6Z/ze/ycAIc8QlG9NsWD2dsnKuc40ZgS2t8WYsw
bISFYJ59CmwOjn6ZC4n0oV6Um/IhRzZX8kK69PHpbR6IkKUdAWZHZWGcOndj
oVotu7l7rCWF9x4QDnAR53uAf78DD1JoDGlorMNjNkpURTM/y0MJJwkBbZtx
HHyRM724/c/VJgbG1Mz2hvV9sZaTe638VgtzRPDsaTo/kQ+0YrT2GdLvW8qP
XOOTWUW/A1pPX0WVPTjfyB2VSFhBDuATVq6W/M6pDI2O4etyhUFSS7hdBngE
hdePZLY5JM6mP6GjjDIYfT0QhDR+nhEezL/Zgo2YFX0VIsb83ips1ZgXhQVQ
zdMVEUa7YK0aHEEawvoOqLX7r+Of24e9zqjAddTXnv06g9JEGVjKHlIAtjtR
lPdnTti4rpkmi7Yr4Sp752avzfPNnb4Cpt1FRVftL++G2JsyfZ4/NGpXlKx+
bqkGa5cCrBJw/b77XaDZRnGuHDFIZwkrSQqHACd1G7gxUBcDoG5h0rh6WeJ9
mOHnzHo+SujkK87OVm6k2GAPyvl3vVHUKgZi5xlGARW/sB+tvnfTZ2D8jANG
MeP8fhFwlkgb9oZghgdpnPGy5hlqfH0u8AHO6tlkGo0DB/zR5RkMqtYVpyb2
Xcdoeydp0k2FcIplWCbHFNXHcEt5iMFLThZ6UCbAYmdxvFGqqR01+5KJmMxp
L5qi/gP/MyhcV3NDM2JtlaNaQYS/hJvMSGXflyPfgOcP6hFRaI7oqnqKJaEA
XH5GJJKWzM3RmIb9CnkMHs8ltpFWyghiHF7LRSMKDxfLynOfmYyYHk3MfadN
5tTIUUPW6pizOZdE+spjmcY+ScIjr2vDYWNYTfnlJeCcnGWs1f/l+0+GkYhI
x61E4mE2ImcqKpkhG+k9fX7y/hjz0ZDXUTPAjZrU2dJNXY9KOd/zweAAkw4k
R1AXoVa56UcFHMHSsdhbr6wNH9MJUMFXYHQDXcI0VVGYH8mv7WMn5ODgbecW
u8JR4RseD/cxa2l25b3WE17BGHXJhpmHhPzCgLNE2D4/lEJ5HsRWDn6mANHB
6+O6dal2Ga+74q+ouZ7/YKhmV+Gii/vTGmV12Sv274Sz9ge0zmQItvwqc66V
BwUcUTb0Nskd9y2Q5MdY8LwU/GTuLV3wo8au+5JVBjYgvLcNr+1eCANKpNC6
StmoZiNbO8TG3kjKe1wqlfzzzOHJXDI3riRc9kwwjpPQzz2MVi8Ticz3D+AA
qlND3IlPqePIj649NDSIu3F27zV1mXpLXNzVXGo84loEC4Np5z5KVH5Vr268
hMQ86hX6TMyjf8RXcZUy8qaL59konPnshqLqeD1q3ZJTzFIoGkq3doVJELly
EfveoWYUGyPan+YYMzrBJwePaKymcnVNX4WJ5Kzu11OZ7/fzrYLrdoMIEFyp
tn4rIlF6uKXrGSXMrAmcxW17azgCIBt9iU7I852qyE1lxI2pIsuDmrnQmHh1
455fcTZyk3Mr+dNCFatOB256CkOuAp0jmOOcTxcuDl9qcli9QsGg1DpBZWeG
wqlQrUuAiKr77dvYBOFvucEdEvyg13rwN7/YeycB5E0PjNa6kmw1X1W3H/L+
7Uvlk0q1ncHizl5jKExOpJdg443FRvYaWxx8hfHYZGxsndG/rUweMX2cQ+bS
wbu5V0kaB++SQNW6LjQONtv6tWbvwHVeQ9A94PDrt/dwUmmfMP18Vt9l6GhD
Tqxm3FQp3z4sFg1wPmDaRVEn9HMX+pt3F+bth44gjIzxlcr4Ggid3lcmjf3/
emp4YUWUmBgrevpleXeAD99mSSrS7hJxKD7t1ZNah1QVBxuSCTVVFOGflsnY
mlOMQARmidQ3F/G7o0OL58fcJbfMgKFNPlmhvCk9Z4kgd8ozM5+PBPUUZyq0
sqqb8pfxvHZ4Nk5cvSa7xD2VQl81eIjMELev0Qg9PEwYTLD7/I7PBN/UQ+0B
vf5NIsn6oXAnOeJpbEukx8drIy8XxFLl9C7ACLHD4QCOjsCI+pyarr02fGOE
YSpS/pPK3RRfLQBz833HrwSEjDOECCkzjchbo0+xru29wua1Zh7KTs9bBXNu
2aq7s4d53EyhGurnb+Dy9lRVoxx6YJt0SmPk0g50ykeZDYW+24qmZtkkI6xd
FxXJzeatJ/iKbnRn6XneaD9S5hXCY3YmEiljcUKImZ4o7wmoeaVsT8OEGDWh
koCHIE0oQCDiw7yBrCM7bRVrEaOWX5Pl/uoxTxctaAlEv2Oejx1ASpxiKZBP
j++DX2F+YaNJoUQQ+1ee0ndB5MGcOlSSjlQKx3xwvfHaccWqJPQ/+ma1hAlc
dDZvcGNUAZWKOiJUuc16e5Jk4S3TADFMfOdgzfUIFCkFNLBV/zZKlcEtNpnN
Z/tlm2e22Z9oLGaeC0cpF/qSw0Xq4diFDrrS/nkhGVR3ZynN2nRa2IiV7cqH
i2DMAI6prbluhh4M/aBafJTgVusS8OkTgysQDlvXCyRkGtXJwVdgAxR6LFLF
NkRh6Ue8I+sK3/Cg8ig3j6LhPbuDmwUQDqGmSaKqbLgGg33foW5OuvgmJjx5
KKX2cDXKJtxRfyeSqTaiP5g0612J2LBRAQkCkBsPrx3mZBO9bo02/9W4aOj0
rIzIZMS0wX7Sp9by7tZ9UkAG60oktJ6NKEkeG2u00Rt1S6ie4vajzRHETfBN
cazDNkhd7p6y4IJnenZ9/6zO/haf9eYB6FU9AEFCTEDZLPBATSt+DG3ACD8L
T1U1yDHqQUUSMq9QYQAqtbQPxorU0tCqRXaLKovAVaCkb6yoQjbVhtuvMNye
JzZt/RTLuV02F4snEOxGvWvOR8nTeR6BELw+shvyYZsX9jzhIHh4H8oaAj8F
m7DzHmkD7HyTCQA1i4/rWDY6IulB+Fpw8ORtDi1lUAosarQf78GDlM5Hli5t
yxlWLjjKJadcXHP4/t1U7n9Nq2Qw2wv4bfnHRWsM3QTnGKo91ylxdELef8T7
mI7TKKtJWYge/0WIomTCJHthGpOn2DABhruUMkyVHPINW3livxRHjlIgBbSD
0vIznOmxcOf28TQxFrL0p8orWEmSEXhXrT02Lo0TjMlyzJXByOkgZU2UNUZy
lxaMHrFGYD5lYuozgQWcMwCs1vJc89yTThzUnHHdu23CFNrU+zoHN+k7ZV1I
pb2yAAX4iihfvLLTJ4p8AHniTzURgIQjrnedEsXxnA0evVi5CB8Yx2gFw1AX
sNCxKSaYoLvoRe0cl0u/KGRS27yJsG+llP4s9PzL1nCPFZ0TYdLVZd99Eyv8
aDYNsLAlPvTLKCZXCroJy4oGh5iZbw/Xtxs4d6DMCtrTYAjkEWAXzhZNqoB+
BSBCfbZ0HdcoATasU6MuUYOz8XZzcY65Xp5aDREjIURbL4vSd1uv5bSpm4FL
EsxIjTYGGZ5R/X4nByRoc4W+SWUgLkwHb4MYSJi3JLz4pOHHlSJe/pUXRh1Y
Wrfsky6ucL+GLEby5qOQwiSRWfhd3YvFFAFH26eqGUPMjlLYUa5W20sasi1w
QfJnbYqCNKQ+5frv28VyHf7/UGm/OyKjMLwgSvNE3T7e66Y8+OVf7RCEs+4r
V2nnj2HqhKy8kH4dywpsnL6ZYYMnKHH2QtRBy0b4Z94n8oO/mzJ1Q4oJ97as
q+tALJM7aVCRKVl+NuTIt+h7mzWSwtONkPiEiDW2GGIzef1y3kKzUuPOuWme
zwPduQ7R1hPywd3eCtInQ0TVHy78be/ZcukRZG2eDT+rmRrv9QF+6LC0UO+c
ywltLxa5t6RFq0Y8Rjg30fWtI9vN7LdHd9RlLPF8YuDckB32AvBE0sOltEFs
V+ieCohU4rQtt9BvddO+SLKgrR4gztkvXx1dqbXyxmlDdqpC9bycGCjr2zu4
sFZ4aSXu/SswRO0S04ajZZWWe+WBR8kKA3+k6B7+15GjyjYqU7XLPaOX6jVe
zZpl21Y1jw7DfFSk1UCmeWZBGN98/dNbrUI4bwqb+iWD9R6qz7C9keEqYrR4
9bp5gig4Mx4OEx+v/F/VZq6lTKkQr7d3fvCiIrxIRISqwPHxfXZoBAVICuO2
1R8A9+j67LirWEPaeDDOYZ3ggfoHCq67+Kzw/DMQ7y1uYn/BxUsVbBeyxqN7
GH478CFHTn3y0kdf3/C+rW/vT0VPOUPCDC86K/MhpoAO8p3VVCmf6RJ+YCdw
gZcn8/SWj5ummGhgwm4JBOhVYJAq+jdrTMuVpQnLMPgt+3F9w/Moj84iFl/v
NIGGub7G7eqdPL4XBXormB14gvzlLWCpHGKl7cEDdByLilOBrJKdky3/pEeM
uuAbSryrnuPERl+M825kYjUsu6S/+AjBv9Hrpn/lleRRgFPQ6jaF05nIRX1f
H+QAsk7XRQYq+cK9QCDBTETfLkSoLBWt3BiFVqa9SmqQ6klJeiCSfzGSTTfl
us5Xp4tArEZEzXBlXCG97nwovJabvymI1fTAdOsxvQ9UxK9PlCBmpgxAhGM7
MFY8ByreSPIP5YGLGyp3NWA71qc0ISD5Ki6aMtpV1y1FYldk7iDKxEHgTFQq
s/Aj+eGqz5l2wgQsSUkhtsQm4f1+zYKDEpeaeORIEeNXXmgHeeNkApcPZ94H
7oZXxLiyns1FnPaPVZMqqtMo/yxQff3K7PJh7aIcea+dj9VNVa7yS5RbXj2z
pkhOZZd75pF7EaV+jsec+9vnTmw9tDfTcI0mL1ArmHaMwT5S/zj+pGV5aAqK
hfYhX+6RGDW+vbJZZx5YZCP5kM7CeHL+Dewo3Lm37mQSR5aY9YahPAcKAADT
Udf7YgoFnsTYZzHBK1N5ebpe7sCQmLa/Qy54FOvOu/MyyNQxUTPzt/CABA9a
f/DnTnDbJK6mIoHV9HRVR6eL2XRZYStFYHibl93QP0KNI9IXaHFxbfdVcjgt
3fbo4ctPfFtOd7qKVhMD3T9jblFC/Rl4Duj2jjC9gBgTthVZHIBt1eQrHPwz
+J5bzmpHmjWGifwM4oov8IwAzj9U/fFwgr2sEoGJ0OAfWj1cTqEHIflZsyAU
EkFUYD733ZzH8f0m7XHStyiJuAz5c/uZH8ORv13X7lpNSI7P4G0o4dhHZb3U
lVWUPS3EXLa1OD0G3sGMSGnj5Gur2fYn6XTCDalYjG8jWBpbnBBSiIarhZE2
2kEp/+EBqeUP71DxGypxX3tMQgFsaqqEutJUIcEbcUtrb/PxyVPJhFPXQl0q
e13gRs4ME9Lm3lRFrE+7kdwKne3sN4/4PLbktCiYkoyUhZQxQ+C3sSCDjbH7
41jYFf9kxXillCIdRPRSv2bNfdEzwbdHtKVV544Iq6t3GnCeqmdKwLYp4XBW
uae33Urv9p4OHT4k9XDgvp18Nw8lmdkGH3BOjLWhcw1ST55obMbu/g72ObQY
Cy3Cwwt8l1TpRTtxlQIBLTfxCjROP/3lG5Kdf+q9brZzo7fV6vUoXrS5zAfw
D+4u3ogTWq0FFeb1ZeaxVH9I833pSXCHoxveONx1UgUP54xBOyLx4dg7aVgq
RYhU6bBf8gq83saxZ8gwfqi0y/U5+9OryIcVEP2O4YG2ZjUIsv1YYav8q/Z+
LUohWP5PG25cNU/D+7+uhOKKuqVH0jalNuq8RDTugTcpyW9968ZqVDAxqc9V
4vkvGY+cXPZb3W1h8M4n28YVyF13ceQosqG/B5QNG8dk0BP1lFLqCmDalNey
NbltEQ/SoBDRzONVTi2gdsn3N/EtIbwXv2HRHBM2x3dneoJvpAnut0eHS3xQ
z5TJ1XioSR6r3uXSVuQQRA14xDLO5vwHbCc7HVK7mnptbZZF++ak02vyNbEc
x4QWVkhrh0sD2JsD4s3K2spL8dpyhRcbSsf6D2Uq9MtLnVTWx+QDJIMuRCKP
cp+yI08vujPRqAK7PQx5alkdAhyXQYUtWP0CBFz1JHiHDctFdVumuspTJ1pk
ICCMoVpwygsLNyTbgrLBS0Ehtwtri2sjOcdxQWlYGH35WP3ffXOsihzDvKOZ
1V3tJZp9aWw9jhaS4iu8fDZS4cOzxK+E97+ViPeZZWrUyF7WdFqrifTyZiQN
QMmYYRJKZ1aozwJ8m+TnU9BTE3gbkg/8gXXaeWSSN6gQsPodhthd3vjUgEwt
oeyBxhIJbSuoZpzJUBI6sIW+aMM1/3lZPHGuKBwlxAHwGGKa7xL7Nnqqx4nd
MQaCCh+UsAWOLio8gmshnuwNSKGts7UieHBv6y07bgp8BTW9GwwbvE2RA7d5
n+hhT53JrghQxbc3kuAtX25G1tEK27ZVlw8X5dUmAgSZjLrL0O+Ods62cmHF
nyc7giukW515c8/k4Ywnf4LAxKs7hFa29usqtAxqsnxK9ti60sVyLxXT6muv
MyS+vfMGgVJL9TjW46H1sz/wjzSQnsFmyjRVoA4mU5VpZ0ATbu2G6bIu+A7X
w7P+XpkTkcwb2De3WJV4NwQGktTdxP4XJY/85DtVEFqJyHQQ9wxPNwB9MC2w
ZwIiRnxzo3S7QWHOSnAPbxc5upb8IPeuGqTr2ySiXsofS4MXkO0j6h3B7AbS
h4TyCNCvZW6gXfnrMcmJqELJq2h4ZaFNnlFQpe+HZIwU7EAcNAdamss7Lh3e
STwmubCS6aBUiMxUzSK4N3h+wD7WLNs2XGaSEADlahIAOg1UpEr+VQmiB4TP
63nohlOIIip8zSCD61gMCoF6vhmGg6ZCcKNLkuNvjUN5WvPvkgesPmcpgUjh
SkhLq/RmUFZ0VHZR7RXg1DlIAxkjAsoBu2GaLr9csjCbnvoG9HTPC3GF1UwA
JkUy8cmKrlDy3RSNHMkqkptbLR7+hEBFax6CVlAdLezuND8WGoPYiezIgX6q
O4bbsNH/dlZP1Ur4vvpHY7v2IHzoOCrsf0XPLS9dcg+blWi6728QjAahM3tF
PfZukPXTmA4ReM5FhXILzY4INsoMIm2qlemY9VlYenqzcGyTBJBOKmNdDKyr
iFthPYYyUY935DW9IjVHOuuqA/FUfSz3bDTDzyc+PJLOJdRx0bGAkZj/5+5R
93Mn5o8KOEDXNgM797O3IeoHD9uKHTVykA1MY14znu8drEBtkJEA8X/5zD2+
sU/mgZY4Uof4V2GljMxxyC+tzvLG3rztcQZq5GByimEWaHeEfY7NZi9xGZPo
+6snk7YrOnGSTkJp3SNDG9v5n9mOWZazCtmIynTa96asMpMhfi149HeeqVyQ
/JJl7RbtpMG8m2DxCORb0qna7BkuSM09QYElTuwcGKaYYA9ruV+gG8D9uM68
xiaROYZxUA1zJwxt5ywRBEyzRStOnI+Fi9XtBy66CUnkPLSu7bbtIdg4asPa
5zAFbx+ykh1UrOvUtdYsjUO4G1AducAkdcgsNmp9bOxk+0NHd+OC/pc7k2GC
TKrAq0T5fWqS2x8v7CjW06p2SJmc947X/Gwx1k6zpzXayZKCviEQOga8ztGy
Klc3h4MhTVvPh2rpXZd2C0NXFGuQ9SEGCRiJX+gyYXM+F0Wqt1b1VOIci3oU
8ULWzvl5RhiMKminAAy1RJNkE3sPAZV0Zkbvadj/m7QLIhAgk3CojWBqtP1Y
OpEbv7ENamQtXSYjlXc9f2LnopAHFl+mgbsgfFRWJEE8cXiBfXjea8GcTyZg
I1+LfYVkv7aifHSqmqO2x7eLMQpa8fzOLL3VXbsBbNM2lt3L1Ad2aks0pfjI
Yrt/GlrCTgMNqlKK9+Dk9QxKBdn+dYsLXfymYXgqErANosDNVvRuZ9UzcIf+
0yUQmvQGrZu7a0rKSCQboz1VYL9+AekNgXBJ+XSnB9kJqyIrUf/3KyJG6AeW
/HoLFazsjQjJVRpgxiYPjnasenM45Swq9pG7j1e0A6b7YkEpnWhEItMD7t6N
W4WkJDhpmjYhkfDGp2IiwUaVLMcXP6b0rRpAYEGEEeJJ0JhW0NbhCry9WkxS
W6ykvxxw/wC8zUh2naWDaEqtok23dnZiNE1580LM2KFPzKWDmYp8hUkGgXGh
NdvGBjVUCKdc6lpATryD6dh//xSymuvtnTXY1D2yMa4jhVWJyX3JV91YCSYA
w+CT8kTVrw1DaZUm70mAFPIYeSqfM5gJspplrK9SjgzkdaGU1j7i29ZvvNO+
MgTq/bQGvQuo9h9PlKLF9UjpJPIarUJqcFYM/qMZXWM4S4fUJ771dj494LhO
udcJzE5bcITVgMEcbgUNTt32kP2hTlPglbbqwi1eFyv6Xz+GLtSCaftsGroX
j2CihTVJFXkhQwAbZ1HHAcr8f0rHwttz3nzNT8jXxIQosMUegP4Usvl/mkw7
2tOUXKSKG96aMBlWnrSoNaHZoNFKFMMVT40lC6xX0+AdzrG6EYHRE4hy2eiK
6x8d59kP93r7wWKc/XK7TViKWIUFqLqCwIeXUP9qeVQmiPkfQkawdh2GdkAg
5wFXjftPzimg48M7AKiMUA7YWZwRphZjP/KLexvkFhCgFZIFeNgN73CGiD43
sSFWEFxzbgVN0w5eOq87Gy8SIdOZmLU5NvI2TA50pxV04AVyKYGApm+y856T
xrVN6Wdy70cGWbKrUQ/SvTEH3wD+DbzdJtEkOZ2hwTIHudUDDDxSmbqL+hW/
VILhtmW7LcSRNdiIl6jcycdZqcpz3wwMeASmjT4mspeVGqTHo3iT12wfhcm+
ViNgQ4i0nhXloWD1NsP7DBQ351fmO5aEbUQX5DBDywtovv8DyfhD6CbuNs2X
B9ma/BuXMIFLDm9dsUwWRr49aPrkzGlNTCUVRerIaO6gJWSgrwo2P/HNeXYx
MrIaJfPundnJsRqQioacTyYydFeBtX2SJwIWx7srdBLbUgBDdC6pz+xtwEXt
bbA4SG+loGEEidJp3l9qnToYdVEulSVLymc94YRYAbqnSCAOYyjXN0sObGZp
3vbxS7ZurwuKwWphNTxlDKYAUHz4xcIKUN219tJ9bGccI5XfVTiKV0RwnY0f
Yd+OqviNCg2HCLQGlsW/1RQfCTo39HihQxmMFmihFWI8G6G6W28SKlXUQMTg
YLbErpDGB6Cz8wtPIWo7uUJ8yWBByx8H2MWdTRqV5UR4TWIhWqM7AwJLOMa/
DxkRLyxqBrL8iup0sfVXsefSe57NcyEnC0Gz55JED+RIegHEig/XgGFuVUsw
38fPPETEa2jseompS6hI2/jMRec5aWD/GpqWB/ZOwaHgujE+YVQLCkkdVKdz
dOaWzwA0KSjJSc3HQUeJSALtjuriz10uJIZP7GWD4fjb9Qkgi9T6sOESAzzG
/x9ek4azzGNVUH+UIxWz0T4oLX1EA4lqKwcqwV0d1Qix3sf7WBFbda/LqWyA
liHQjIUwOCp95f0o4nN1KlGXW1XiVxGuyIEoTDrQ28tI/OhRFpoLWDE9S3hF
ExSXOc9GTnUGHa/wjSmP2lCVm9VpcbD7KssriXNxcFmMs2WfG+TPJancKFDl
3I8B0fGnEDiqNcn+9ibM5ritOmmAoilZSOra/zilPqizRxLP66QvrHXnMH9a
DERed+czKrTTwQm/xzaoJEbi8BwPuF/mNm2lI+fAdqbiWjIXOrGYQ0VlMHxW
d/vKfv/5FHklGJYWCs7hejBtbh9qwdebaeY+Gb7H0BjjcrPKggv7PJWZn94t
hCnAsrjYucoPoDwXGotcaYSzFLTHs7lS0XuFvqwrNqICHVcWnF7CFtw43h8B
IHXGkwKwxVVNjmpR7v+BOD/XBuRcBcD+cYvHUsKlNKJDAt24UrhGiZ+rvFr+
hWWRhWsB4zhU8/mZgf229pfgpp6a+tQcqwIEfFlt/b8m+sM3zdLH/BI5RcZn
HtaccVJWvwj8SUYyCXdk2AmP1ec7SGNHDIpD64Wamaq5RKt69TOtenYcYG84
1o3+bLYNWzV1BsamOac9K7q+89GDQX/P8x1f84ATK/c0ijDaLgHI5Ex9lOae
eqKJy7qXcVBShUTtxVc0KpdnB7so6uwQO3CTDEhs6fqwDEr9DytwKjIvZpPp
BwxW+a5JWXaUNt0P1CzrI22ItWovejuB4uydzDWY4AMCB+9NkEh40inIlU8r
YtIHdn46PDFZ8whFnl5UJfWkAy9dfc1ECB0QAvzIeRpJf+7MLI0HFFHH/KBt
Bvuu+s1AN2NsrEVEeE1dtdjqZHFn7YUWzxt4hrVvkQ7m8gK9YITMuCRuPari
lK9/YsUq9+7VxDGyLtC9JRYh/PdWleVe0y8fbcU5kw/rqEOFtFzMZmzNYl64
y44WqAu9ppYdfl8IZR814N2LKq+mANhEbOwuQSC91I/mBuM1ObbTiUHF0QPq
UcyRjAeJSmb4bpJ08f56eztgZP/Rh+3hcjXaegZJhMyMIAMXmRVb7V6O5V5X
4ekc6JpJI7kbarfYwzWMLSRLzGTL8wV9TDaO035b0MIhI25vtCAlmjzWt4Da
vVDO26XSsAdMqzhHLyGG0mHd1dTosAHfc0ObPO7CGPqOLgDJtMZgznVngKRr
1PIWc1D8AUNHs++2gLpRlpDyUZ60eAa21hDxVwpcbdhKHrJyt6MFiP26uIsP
ksBFC4jalqTZFI44GowKgOIKfCHQ/cTSCq96fLlwwBt2tL+XqsNOhBbfStRa
1JIofEhbXok4nxU6lB4rna+nWEnH5Vh/VUug0u/zxgWCpPJJbnHx8vtwj+sy
NpuRi3ARmj0nxhTtNEo0oLQewT8hATHqS3VI5JlI9QsSN4WF6o2VZI0KJ6fc
JVVlqHaAU17psyIbvnoJd5qAJY37wxUvuKkPsFShyGOYUXQk7GOuUZOp/ISI
7hoAmGmjTDxsCXh12VJO2t/Z9pjMTbiAX9hJkJG1U74AmfnjI6UgZI652RGD
9a9TZKxmSd675yGqg7thvA95OTnT3KBXqoN/+4eRGwlRsVGnuH2zID1cnYB7
JtvsRi0x/R0Q5rAB4bWXPp++zJKAwz6XJ1V50mJW0le5xLHhbWiCLYB1byer
I2IKwmZsJDhe+ef8q6PyH2FVZGPrt9jp2CDsohsuUe5AlvAwA+soKXzQ99Dk
V/Ax/AFLQAEGhIcxmOMWZZVnjpnSoFuhtVZs7N4jzUaHWBhmkn38HCLDUopo
SFliTluAfGXEEJewTQ8GY5iUjcvulDuTuKk17tnKabNa0FnRhSrsU/dBXHCU
gf7W+vj0/9pDnlT76uJpVybUkNwTVFSZJs+Ah14pnqjX7i6knLdHWyhcEf2l
7emgly92g6Dy2YI41kTfAigjD++V2wPHqL/BGeEadUUC4LpInoNm5mmyexjw
fSGKxEKcrJNItLOD7jiDZLEjlq1HNN5yc3nADywU2JiWn5IYtBf2l86Dc6Wp
qPgywjGeW2fX+Sq7HSr3wKn1rc2ZjZk0gxEt6lEwtKLOo+J3vKMiSsr3YsVc
8K695wwLAIKavhg9vejS15PHBLER/rdd4ZruOnCe8nErVY+I9kYXOkg/KqUP
D7WSBbwBw2pzItIW+hUzHoam+g9guUe99mZuFnnHmQ40KMHzeCWzTA2yIHHp
Chw0mpnMHbyqNK8jhEchsVTWVpf3zOqnu2r2i9JS00tMoncS0Bub5cN50fT2
bx5Ac3nd1kv1h8/CjJEjRVxTxcUaGmIIt09qwHRSSjIlnIgrvEqmLGM6Nezv
AXFc4Ryg3sFfMOiqCkswyGu8DU/S+VzZNqR007kGSIRtlDfa2ktWIkArGvcY
XxG2dJNnkGoV6kb/50JmsO+p+Kt1OKLKzaXaJ5T+iuB9GOREnyI62xlv2/Le
MA2Lq2lANMYHWvNsY5afLw3V0U2fxm/vNZzcmB2rTj6Plsly62uhIio+ZeX3
tCId1eeFPRtTxDDlM+mYe7vis15/+ct/Kw5Zx81RfqjHgZyjPF5s30k96wxg
YRie24tXpM+fkVWAAMLIb0vLYLnz6f1aN7q5YLy+aQ3LX2FDm6M2EXnrpFTX
IV8vmWbONF+WZl98kDjZe66njAz47bJDhZ/RR7s78mgRiGg0icA9ABr0nrIT
rz3aNwp45Xn4wgSjDqeYwCq2uYW4ac7Pe+82IKUFcIJOw5mu4zoJ0ma9KQZ3
je4QzZXxEVjWIGB2QMZsOUyzD/ZWsWp4odio0WoIUHA4Jd1f5UnwSZYpCOCH
UlKGQitSW+iL9iai2BpzdSpFiJPJgtOtgNwAWMbxtpRISzaOqfHrbHKiNAAf
KWWV5vRXDZggxFVaxhrvYRnSEccJSJqm8Bv9DtuzgusbEh16N0tPsSGBEc3a
CG/10hfOLRhiKyh+vDsh64vT1PFHlzGgMWKfwnsA831DUqAz0OsJuw0qllGj
yeg/9POQlTnZVzlj5pYb0wWYJOnBtue90++uqw2juESsX+PU8AICTtoMTQms
1K7gU3dpCsjHuzq8hIMVGVyNNl8pIXrm/T/VqjZG6hY6V3iim+dC55lkjTje
TI0R3B1z5q22m4u5QXsGBUsOs+aSVDTJXWPlKOTuzMbkQejwBVP/9CoJgJ7m
Ke76KK+p9EwaHhgjQfEz8uwldWOCIp7HAAqHQ4s7P6lmHRehB5XUfEUMQck4
GYMtwKCul13/cuvujIgZYegD//sW0tldNfAUx4E4AGizwbEl9eVKwOmKqkv/
EpV7VjR75RTd8O0p50cpCmp1gg1o10VRtFMNeMUgcLf3fnzis87QaFTv03w+
a/dEtgLObdFUAkwAWl746ySBJv73lnhWItvgazB3iAN4JdqwO++XbalQm62K
mlC7Y0Mz4OT5KtvIz2pcq8pPHeblwoOxMThrqTNWc6cCuzmoGSXwjokxZHnb
4ZHth0aprp++fQoTECWV/zoM8aaEakIR4gNEu+fVYi6mTUE0hGRPZS04L15D
OqMPrco2X/eRq8Ld3gWWYYc8RK/FIQBaQGVQDlOPiYpdsJCyB2mSnAlOLTln
pc5+lWY1uMnFs2HrgvPjq+slXFuuQahtILyYGCcxsAftO40ACriB+gXZOfZX
zg8rEn/V4WDuFJiYltLJQq8IbleqXmXuuA2vDQZv+tA8IwSXmQYjGlUQUinG
dfUiIU7zEeurHxor+yyQoq6JumX6o/ne1XMFUeqPIZuGZVMuV2YV5HErQqhe
R+80JT7WnJ3k2ETjbqab70+J7HBJ3S53E24w15w+WiM/DeRwxohJuV6I5fEm
BlQB1UZtm034DDMClDo72P/i/06DnZ21tiwoFGEsOg5pslj0VH5acMODB2Qq
PAidcEPvEcFOBy1HiB43FcD1D6j7zG9HaKy99VTsiAzX9ZmG1/SJn86oDO+Z
yYYMsY+tX/Np0Dnz/5OgVgrDT0Idr+WR4INQe2pvX7CV5EP3oJlVqC89S+8e
IFiXVLHCQwxPS5epoiwupMPOVpMXv2b1thP5SoWsRBaN/v7if6QdRVi8LNCf
hBoY0gUPjd9gXRDZrkRfJKqOyhzgacUc/7z0VsT3w6ZiHkrl57ub0TqB2bZI
sYaicsOfwY/toeYQjD1FFkO/dfamsM9mKwQWXwlWTSb7Tc2IxYv7kiQHIHzC
dkSiwG4Ds7LF10G1NSnD/tJK0mdXC9jyuBrzK3LM+tUnIimrfBy5ztPJyUYl
0KUEOw3kzIXdprWhpa9uHNT1WMw08rQJpQH4bhtKDrZH0IpjdBvFajPVK++R
T7v08v/SLvd9R+cpPam4CabYlizLggnBaeBbA3XTPku3WI53hc7EM3hisd7x
yI/5d5pnoRBEAtvzhvrMP14g66jULiNc7zm6/pfVTlJn9nLH+MiSbS5MEbpa
1M3J6SKuF7N7JwGeroqBw39gRrlvpGMVfxGErWyeVgOYWFbQwadzzaY7yLEk
g4EMkl4n5+OLV06F+Cbj2PbtxLDYOZaXttBvlXzqCPoVsXNkm9HoaYKDVJF3
vXG7CA4yENikuvotCAvLfzI4Sti/l28eINk/1ZIw6J5KnHpC2NNgyZM1VeKj
fqKBaTd8h6gwD72eviV2E3AjBA3afhgWLhOlPEi1H7eqgKl4Fx0Z3oLr2pHy
YoBmzFrIDd2Xd+c4PZoZQTIeh8Y/OdcT9v9hHTdI3OOit86fbyfdZc2FAu+a
mV5pUA4xrkfqP4iKotYdxTGOtXjKaID+l/eAZt6UwRkAVXgfdZRW3c+zPiwX
1rGBklGELUCPPSz36UKirwWeIX4K4zlql8AGEgdwFubqzzvIO+Q+jKfcUY1o
WdlIMVn7x03ZPqpImfNdcDJihP5KJqlKeTAOWhv4YKGYn3aBrZ//4A/iW+Wk
xFX8B6JHNP6S88oAZa/zRG9+q2/jL+Bo+K82Nk3mo5R/ze9WZaEaNnwS2hp1
kjBp3utX2jpXBkDni/fvvRgBI1M3ahTvc9q6VLsuVHOVu7zDX+rsRlSt8PTX
xWQwsmZwSRfp6gQpa8mBDUwCbPyrm7NRF3qf9lSqml0Hd1wKjQtTDSCAwKJ8
lJeUmEad2WQWE4WjcOVu/yruETejsg8ML4dVWIk3GmJmxaKnF4KUN3pqMZHa
3wIYmBo2aW6kac08QDs7VFmu9nDWPdIMu+/gBfIdUlMw71ocjd7vS7fQ0II2
I/l8uVrXyjb6i+UaKe68zLAdrzYYcZP74U4LFJjY/SrfT0l33FgmRQhXLtCH
oee59e/oEpYMf7Jlca+3K8Qv2z9o5vXi7wV6tAyftAi6hHlAIhC27M4mELSD
fMyfi+18jV1tLijeWQEqtWvVdeZVvNX4WO+jZj7kjIDfA0o/2DwWxj7uJRIT
OV9BhJKUC51eUkWLIqU1Hdd3SMdOKrjMoy1kvpa1n49OG9pXRfWvSvC7XKlq
qf0POVYvXwsawCIPXUkCI5PaTBa6kr+SVpV45TGvn3FGxdBQvcC3/ZqHIIvW
GUQYbyjKEpkMDBhDtx9jInLVfPMkWDtuR/PZGhFtNm+ET1YeFxpxcUhXNKYJ
5cKg2bMfOs3tyStKrrjfWlX7Db/LouqQ5G51z86oIYjJVN5aG8x6GTEjMjyu
M8v6Kscu3vJoDt2UTZYbn/cuW5OAKcramlZmDbzF/COG6cHarHFa+Ger8622
9uybxeaH50zd1eeUioevm5wSndSu70FvZrIsewSQH/5PpQpqS7jFvcCiChTl
7aVR7tz76Y1XG+o7gjL5rW1DSYy4DuTC7/wVUXKklVqEmsOzTOM/wacP9fjc
1zQ/oLHIcOHtB1Zfael0Rany9K3drPYl7enotXM4MoaV19SZoBUuNobiBYoY
pE+FYKP82UOGgV/k4alf91VM1ZqEAuRRl0DdoTKnBubhQgSsIsXMpwY/Rztv
FP7bjehoviHAiFoKu/2k9ZjxxpXR4pJyW0DDXrQXOEcZtvPdRnYRMxZlVBiD
RTISud7/MFmUaskK5ojYvxGE8SbxBia6mCvxBnKW30wJ56eeokwScCsJbwJv
6NewMzE2eg++vy/KGaKc67GQLeVDnwFba2bpoLyqJ9dBlAWyUc1aP8JHt6sj
RcSDY9HKVOj+cWAvaCmoeRwnKjtOB6pp46UIgKvqBRaY86/yZJargJhIpqjs
IUE3v8pFqcE6gGBjMe1P6U5z2WgQYh4qmIhZnqlmwQIU0AiyCrWmjCx8iDsl
10IZQwwVg7RGs/Kz7jNaEWmqn6PuUg+idOKjmm34Zc8lpVRpG/SspNcMY9di
/naRp6D8/GyR8dCS6qvNA+TbBCS0d1Nj+38l3NWZODybWQo4fP1SelRxyIwi
x351PN9/d/EcO6w6kezLXTXZlkRZr0o7mpVCSInlx5OcJXQh2iOJTnIWotE5
4NsbMtk1wdfIVBcFBb+OnmpE7OXjuHwSAP0Mr+MCKV8nYKNcsef2A8ILBVvV
lfydKCJ1xukXew84PjTnJOcYwxuDmWqNRekDOPtm+PAPijidvKG+XvSr0lpW
AlPU17smES8LcIJi2UamNaOoYo8NhIqAQtSt42DJT3EgS7TS6m26QZQoX3mz
9usUClYh7oiP8vLSF2Oq6ZuAsmv57oWTv38YURARxaDEcIC/S5SLvLF3NCGC
I/OifVGtukeJkWKC+Y7Cm6NWYlkg4Y4BM8sCCYzxaGvu9i/QihfVEL4RLkFp
lh4UVtsSHcextzk93/fryTD1VZlX6Dw75BGQxJjJrbsBYG4GRrLuhMGTULnL
S1KX3lDQprzmIvcbbba928treO2MdjYWnEU+EtQS0aol2aJLwzYf1bVkYEtt
C1BZIWK9tOnrujhtkyvAVY47r5EuIZr1s976TeJkhoAtv0kGm6rHwfY4Pr8f
d2qyxLZP+/bCxpypQ7pLaImscr6J4ZZjXlbOlu8z/08ZMFDqyU9GlsgKY9p9
VMg2+VC0CwFgQ5oO1CsFvJPqnSLMJXXFoHg7zscyLL1gGViVVXkCyfMcIi35
0rNXNPrY3Lq+dwEqg4UlZlxELo2O4UPpbD06FHVcpQXyKfb1zrGn4N6e66lS
2a5yAaNVD0hNIoaBRaNrA3XHERXj6U8i2bQi+CKayda2nqnZXK5k+vO9OPm1
B/lj/R1nZgPMki2J93b43agGJzty8OIMByG3oeuVOnHzwjeoUIHKEIkenq82
hWeBFkfe8OE7oFg9D7Q8pJofFS9CHl4Jz/WZ3dyA5y4ZgdqBVPfsU2iKQT2s
TtJulKwQ7yG1ML+PauO1+8BlxmHTkpta+8wHKs7qClxzcUdHbIKQwg0GKqhy
qVWYmmLBK5CxuNvA4VIixqdgvIoP34mfaVRnWp1U8SX+73KL/kvaHrOg1p79
2P5v9NfwQEi0QsXsdarqeT8PrUQI4ORVJt4etl/zYKKOHtQ8ESHoBKXbm5mz
HTljMfQjjEAoo/Hce8XwgUiw1GgtGCm4jKJfI2ONVgjInWz+02IVBrwH432G
yFqVHkGP33lN9o0L4aIUy9R+BRsS+xXW9WjCgkQsoo2FS/2c36e/mkZPIU0e
qPL7vlDxwwVxJsB/XFb9L7EO+jAzlD9b/NtpIXEtG2gx1cK1/OHszS+xanZM
zz6ddNayk1eaYSt1bgFjU66IjZI5qhVxfdSjgDEhST8mMxCcGdJjLyUTf1an
ER17Pm9iXqqFfNDNaL/xPWMsit1760gYZN4VN1hroHWMfHFpIHw7+o52BjAJ
qkLzeuEH7X/Ay4Zrxokg3yH55d6KkKgf7R7zE/et6Phw/E0CQFJ8uFNZa21I
FDyAhfcdHylzAQxM/QzJ2FpcNq4nI1LlpNzed6/z50W2N2EtFroTmAY1YFhN
ED0A0L30a0W703kbk55dc4tP24kg2R5LeBgkoEy7Qn83IDU8NCDxi9HPBrHr
rWAEJI6AA1d6XuTyCITrLxXTh0qIR7+XQOY9adyz3SZ06zwY2W4Z8JImAgdb
CZPF5Gl7Kcz5sIV3RRwIcHlwCBJwxKXLaxgDjoMx//u/RqthUTrwqt+bEI3b
iBTF0e5yMGuv8/xOJbkOniEHwY32GCLESbhQjV9O8wqEvNVLnd7EBJRedkVC
bAYbTDcv7aJVoiz9LwilABM/NQ73T6rtqwroPJAoEUQ3OsKRjqzqtJD0vtKu
tTjnzFkH7s3GUHuw8OEREarN9C8QSKz2SQ9ID3YOQ7bdf1b3cmZuLy9e3duW
H23VrDzCj5041AeW0eHD/ArPjtZWnXbt/D9xnamZ4x3a7x8NpeyBvRK5lZ5M
t3eWXmgAcPUZFv3PXWLEvhSySkr/pVjWnHIjLTtyynZdLYszAg47YZqkR9lr
uJEx1kGLAl7XXWtFmgmp6CUqMdksjItuu9s4n7eUvsKdgIOuA4waojiyXe+U
pUl8OvJk4BDY6Y+CmEecxJUL1GHd0u2DQ9WAFk8i0ERco4q46jRPHUwriUOQ
UeMHHgkvYch9Brb6OI7I/aVUNYIWAkMbC83z1N62X1T138O/F41C81lqmY6e
PnRKimwL3Q/1Wp9wHe5cQcTBf92xDlPIc34Y3WmJoUEHBWfHkRC/PHVd2mal
ETRGgosc4NxHv0U9olGSFL5AiImWxQfpj2/oK+gtTO4Av4UdH2wk68NeG15/
pGpzCZmuBKCvZ2zZyiAKdzi8s++oQ5FUW91wWgKPqFjdzTUR9OWkmalUaUn4
h32HUsA/9gIjDbmfBwCq2qioPFNmpbcKljQTjQzC1e/ZZtv4kFdQy0l7P0hx
s6fCjE80M1LTMjT8LZ2e5979SH3RwWPtu5Jet8Ib8vkWjz171MmKX7hsUCRp
8zBD1eHSgs6n1wcKG05nlVBA4zxoz6xDAI9hoSEw+Snc5m271gpeRNhVg87H
K3U8F1r63gr6DAxRhhvRSQ979Qa7viUpYpdIVFq+z2zwqCDDFEDQzHVHLZFR
1qIgRDKrLin+a0PlZbSd6xfNy+MUsSJ/5AM6Q7cxW66HjF8hXM1qR++Ul2PR
UJWPbaLYa/c3s2oAr2NQOJnKw7UlBGNHTJ58lq79kn6Kjo5yvUt6PB1SDQH/
ckzWLUazFfFHgtbeDPmMGsEblUAiu71lX9aCeqdLlcX4wcJTEdC917Re/QtK
V8qbAu3tg+3VDmn7yStZGYboZPUTLRWga2KHQc7bSzR9ZwuWLY6WoCBRKTTq
0Bsdm2K0iHoJZPEEpECzz2OuRsPGZNdMGCtx2acSIu8Nx9z9ZpobKVAjN5xU
+pYgR3j+cAFPB8BHMhi5hIPxAuWKBiHYAjAWBpfh3GgT10Q6/qRLJCZ3HMP8
mtnNt2fq9zdebsUR09S+iry7zTFtmNxpjxCPaWZvt/qGzjaCdXaGZ+31BAYC
BUtK+tXKjxLe5IvKyx/s15OVvE0LAZOfvqEA5yFiL5GIBZbMrgSP0cVVln5I
3fmgzK5K/SeiQW0/JCAjisSq4+tKppYnZWDenxaXuCeONQky8391pEmW23T+
OtmRilkFAFaQ5qVOa32kKn8Pmx9VxtHAWtFCFtu13EZ9oaAMWggYcpqCy/Oh
PokK3M95zAdsbNi3nu/VOLSiemdPkoWczUc8bHUHDbeP/ZKHJx4AR+zXzHy7
0GCPcem7rnHDfEKl+HwLXtisGAT3fBHumj7846itF5BxZVE6uMUrVMM4A9Li
ZdlkqS+YF8Nok/BwE5vqFfsRPgMsxrDFqa0b5N9MU6wyMEn8QIL90nvEt1PD
ZbnCdzeCYhmGh4fMvpAxqgzXUCw52cD47fQXD7zBBsTLdAEn5ERI/qIZ7kpk
hSo2OrpxRUygQ5LLenHxDPaPPiq/QLl9p1J/pCF6pVDIxqXt1aXietO/KRLS
65Cf/7bIBgJYYJEsHJcCvghvYs5DBUQdOYInoylgncteig73WBe15dK2QY1A
iH26pcDSP8cZAv8ckfDy+Xgas2kMHiuXirFvdLcEtNyLOeYPmlKICJw6bcAS
3DYWpOci/iLneR6he5bkJtUUngNKs3uhBMjVsPS1n8R3QbZ2Y14quYvkFcIK
xxQ1ah0Drqb5a7w4WZWQq2UT2oerW3+GmXT+AyznjN6Rp7bn9FF+7bYV6tCC
iZZqVqnAnwgVbhGRQJ5Bbeh9djeqOdk7pr6fB/60iMIZBocPY1buCQmgoXUS
xX2X3krmWLbELrbkoQCNjYnUT7Bo7x5rdLg3THhvbyxFQ29L/OpNJzyl0Uby
rpPkOY0vl+tM+LC4UotcPNaRm0VtDJH8QsjMWni9/69lCfQyYuZ1SFZ/CRGS
39d3bDS4lpMiNLU+378LO8xh8NYR9zd6cWt5rVR8rxo2Yyt+kobh3DN3HYu+
Qs0zDteO7cvJPitSupYs79Cl3mKOdPjTseo2WFxK57JKkwV2cRRnpwECxlCJ
kWj1MvRMhU/mPIyuZqPGgQUP0Wf2nLTkS3hFMS5Rkeqp/Hap+L7HJLRuf/cB
OlUJdd90j8sr4PvXI6GZOtCF8ZwLL6n1klX9nUyxAyHPkBcAbc50RroiSxgd
Eh4wnAUUnZAxtRLKgUcx0379HoI/kQQetkdhFRYJ4AD/Yqgemwseq8UW80yV
vo4/9SxSBpXrtrBnOcNds318+jYd0LTrr7mCtDsmqeNmDgV7OAxFagOfCxhU
5sBUQxAmgFPulEQlJBmDYhynqkmNtCXCoNk037oeMFAU7FgHp1UNfcddB7ki
diCMGZYtnIedSqx8VnXUP8kAkJvdsZzYjTHCfBwY2SP3Orafwc78UQmcDaeP
VIiD0ox6XmpsQeXnSRgwFetB0VtiZZ0U8oP7oHHT8eD1QMknEUAzMWu7QvQ4
mH/S14kZ5asADB+xmJzaCQLCJtn+Q5p7OgKCMA2wolUrOp4oQTR58tKWmJn2
QQl4Fs73r/gH/huTyOxKxd5Aio4G3vqvOJJYuU3fCt/NgkFHsjZ8TELSwUeT
GfYVeSuYenqOHJO2Q9e+AYtkhZWuAJb4SUkjzytNNbg9ICzzNNW/zTxGZbJM
ySLTpsQLvL1ZqbIWGwGQvFxIXCQdxJWvMFd6AB6xGwT9j9ZG/QML9XegrUkq
opb4D4OE28FnZaRaM7dpuLYKwV0CYGn971JddiVJvp7E1UDoxiBo6C20b9Wx
PKLQsiE4dgmFE907F6JiPrLr4RpBD7blUc+rPEV3RCk3aN2sMl6ErvnBnpyh
qL/KL+rxWCogRdrWvG0gy/VfPnWZ+ZZgy3XF9laN+V86bVPO13uv9VpZgfDv
kIbTTPJHZpSCNxY9B8ILdNexGYy374NdWGByb9rZ5ts6XFeIvAzHcL+StyMw
g0I2/yJeOWDBU0CqXRL8RPUWAcpcv0kvmMCb3pBb8GyxItdEjz/C5Ql0D2cK
uXJeubOzueIo1t588Ae3Ukt1AIMk9NJ1xX+wuNILR1X1qALwzvzq3J2onBL8
cObfKyS6Evrb6Sv7hNdfQ/R73q+0VdvA81+TcIDidtwzv/D6CPZT6J9ykkA2
PPyLxxjVRX4iOq3wmyB4Ue+dxTB0mgaGNxS26I3lC+226Q/q80/qZm6hy2aJ
jd/zWa9Fvs5aqyVtaR5e1sC+i5gpMhCYN5VoOvt/FEF6zaG4t2nFNicjdZD1
c6saWoGJiZaX/RzzU/l2xafxDbaE5VedO2/sEsmSEL0LTOJlgwU+NU7JdxXz
iVCHgyju2MRlRea38EHB2StD7WHeuVNPBYJtB3t7FsuieaniN2DLitxupZT9
orihH9ROcrlPtANMHXzQ0hLdaE/OyauxjI1PaGjH4Qf5DOnhICXJEs0TNVai
TpzR0O8GWJNhTX+5c/WfPH6Hr2zWu7KiJJt1vHAmr3Gis3t9GiaRDWOYZh0q
6NyAc2QdGdrnj0xQG6/8fS0J3vJh7A1hpp1d8w+fNfjmREQS0aTinuuGID6c
3f8UGImFc64mwqPDxvq6FwXHJQUCqYO9yhH4MGKvLfSR7r6lD+BrhJwxwgGH
c0iE3uHFzGdco5G6r+KgXpMy4yF/G8NdoKYPA1iF9HYcvV1M5zIgzQWmovFE
6Iy2EsD1cT0JQlOl8LEOEnamUNyaDfOjRuGFEZZGm9UVHAAA5wT/To7fXh/t
iH3cbABU6+DBTeHG0HBuvR7VBM3lcTru0UKID7yBZI9A/x0hEZoj9r5klhuL
TtXavr1TRYbJYqZ9XnK09PgJDMuauyPrr2Y/WH9h8AMcon07FoAT09WJyins
EZIQWo/zRyvJWQdZitLIgCYDGlS4ZE5DCqRnNjmwdFZus0OQEjdLdiAr9Cbc
Tfk2Ekvo62Mg07r1YBCKvwQAA2ifwCr60F8DTbvCsWt746AJYP3zssZg9SMU
Ej8u1S3kQhUUilHmOfMT3Q30HBFj5IrXD7hWcBDJtaIuFSewFihBrX2KdnDz
m4sM53ZxfGgmUPQT9QY6vAElSXeRqf3Ex5DLpzHSs6tISZ/Pr6vh1fQsrLkz
d9lqR+tXb1lFKg9YBze9uHEAo4K24YgB8u0wwh6vFp/XVeXBtKXFrXy9M9qB
6vZuvmP0PL9JZ5K+eycHOBjwDYx3sNKkMFtLwVz7v4Di6rW0IKSRmp6mdnOw
eQgWO9tAbDzEDR9263FhCMjuIgooUnjyojB+30f+pLrmbT5HLhOUl6J+Tuxi
2WoBWqdLrk5rqog6eWOsnrWpRfU7TWv/wWMlM8HmXAezcpJTXuGUjOMpSlYI
7+YDwot/oSr5QKY8x85ipy1CdTXpDX2bFg2RMQv7ppu6JMOv2Joj/bsQxV0x
TMCvKHIWeV2rtmS3g9Di9NHpS0IwA5XsT8Gvyc648M0jvkstklDETAlWfTbX
oWNHqmpjwyHXdOKpA+UjwPEeZdKRikz7iPsLMqiesf6VX0EIcZoltslY/B+F
tYcBYmLbPvS5astSXwz9BAkLm6puQhUt0u+cV8ol/O5g0DxKIX1Zcverqn1X
a6NgSqrUeZQi2vcSbXcjRuu9NgBVIo3C/GebP8qkqKUMduSSAeYDaPE7T+qp
ViU5o3BDiRqfWDhzodnLuWmPFEXOKH2gw0Fav8m8MGIDCBiF+RjNzBwE2L0g
UJByeal/qG5DTzgXKaYRVQukBqS1O3s+EENfUebdVw5sjbq9NuzelXh8SoGG
oYmHuWh8YESMoDnHzp/3Xqt0vXMj1Y6BJYNJCuiXZgAp0OphAUTYDwF3Tkey
ITx2RhRZ0UVrTmWiKFaTo+Dr+OG8jWOtSASzKBtTWJ1Ys9EJffcTscROlUFw
a714N21xiRfai27hVN+vOXE8sgDizBLyynWcCioksV5Xg5dinDLzV4f9c3rP
99hnAbg8yLdfhS5L+pJoz+4MXwoKcKa6gLqCshtxdKejtHie+H49x+fFym0x
/TjNs8vM/WeYYyi8lwqY1vS9VZeYROLvP60g2Mb0ZfY+Qg6vJPdTPyFLxMN5
B8jSkAeBl10NbFJl4dtcNF62IDUFFhoHIt8UOWSxDST6vwCJd1EyiiZ2Tdvy
WbF7lDRz4XZmlL14rGc+/2htZdj6+Jzp9joTsJQPgP85yxsOUi6xLUrrbO9/
dGeTjsMaSfHChIkM0CTDXKkq2Xn32e8c4JjjBTtf0zcJ0JpLiiQWyu8ImWCE
bXnTN/98rc4ddPTbwpCpTGu66sIFzn/d+hBGeGuQE7pG80VxAifil4QABgE0
nBQxKW/TEbPfSAwy1Y/whtHapDBkWG1V8Cm269WNiup6PpnsvJ7xjv5dyySf
BoEgw2b4/xxJ9fNdkjo3+q0mqE0Ml+FhGf6xtAGTZuPeUnT+wVdOVBGwteCa
sDFtg7SQV56ZufwnQkncnDaJyUzHTunDRWhzV+KhAlajqG9bOxLWHxvMy/S5
g6PjCImBJbIyk++dAOEBulGVH91mj1GuqSvaCVLzaPSPibFE+MapEfEw1Xkf
Pgqhs9qGpsZ8VWZffr+2o/JbG2wMn8te8Ys731QSTfyjlntDfynoj2PgG3G6
qRmwGsTQckpE9yOz0czWeTvVx3RdHqN6egz04FduNXOevoWLWS66Cx4fTTf/
jjkytLnnHXdidOHzFpZAXPLK6h9IULTc7dqaKUmm6r3vD8yEr50Kf/SFyrFv
Whr+evJBuNSAs1E9XmgdlTJEvncuEfs+VKo616RSsDb7bm2HNt1WITMv5fOq
eut7dk6+Y4S45U5h3wM66S1jl5OaJd3rikty7zwNG+T+NkoUlnWcHPb11rRx
HEHSWwzI4lA45ZbeNYEGWXetC7ZnF5o0oiX547LTu7s4/rKjCDzUm+1pKvjW
biYkGdYS8Q8Y4F0RUX3A0UcEhO3ER06O9+qwd2Qe2KdkmkfJAirVqx03u3ku
wOYJ2K7UiP7ZDusM37Z/DjdbL70uQMYYAuFKnSrIVfEoZHhQ30CxljRNgEvi
HeUeOz9YBJ3BnFW7HvCgIiDtmKv1vu3d3Q/gVbNjHRCwOguTuPtiXo3WyIQ7
fOiT2vLNpgQLQSDD8iBrNeN/8QOfksYBJlxsH1PtFvS0Dw8hrCL0LAu2LULP
yqCyr4p+sB9iqbQDXpXJRU2pic8dIAwytBX5zg88mcGm+HsPKWMOYMc6P14U
SR7tQ+O3mNL8T0UEjSn5Lxy2jPGSeA8vCFAVCp9ifi1Im7eaNB6aVkw7tnSz
XpSis9anI6ONyvw++eo5g3VqPQPxDqF2Q/+woJCTlOTm81plN6DFAjCjuer4
4Vtqkj3uOMndv4kDfTqsrWi42MSopQPHh/x0mCw97k3Knj/7/JMUQvBf7WhI
qcARg5NWKd5djVV2L6rI6E0R7TUtN2YRwQMSvkiZtVnxH2W9tM4Cs8MjnP1D
CLIiURgLZEfQWKyxMRTsjdVQM2RkdefI2s/OAPG7rYOqtnos0Ot0qJ0btNoo
oFttewFGgesUuhS/V81SZ1IM8EOlpSgIESSr+ZFEt/APF9tX/RIn9f+jbBP+
JrbhqAbJDCdygwwdQ77kQwsQIF6tdzT4Xj8+oP2z6j0fPwPulnZlLuMXG5Gm
bb7hfTcjgCstV3IKlcOn54wVVRs00fzgtKaW2y/U979y/++6rCsd5/aoPIxK
XJuOG2V2xQ0wH/ug7avPmdc+NNECVX1mmpYD5YGQFFn82eZWJBiFXY+qW87L
LqCjunRRhP5JbpZWk154ApYynZwOKBWvpxdFGouNO9BbW16WcD4fjlRo+9RR
ne5JN8zo/39KL0AmRa/E7MGl33Aji85kklWF+audMxdnynbi+RRpmKw8Zr6B
puMr+Wu2pAADkt7RdePfYYaGN8qAT/1N0twEDIG49rV/FkatwN5HYGMg/c3f
T7g0zV8o3h8K8JyP1h2JUq/LhBTbdfpRGykF95dwBn/ejdJ6I6d+U4ll/3z1
Cp93zho1P13LYJLL9OWybsxnwUNCyQQ8YnPXCfZI7DFHhfB2lN550418Uqh6
eJcv2wliRPCk2YkAxNvTaPo16WDLjqECD+VbmcYV7UbxMkLBaS9l3czegdmb
ErY4SxAGY+8gIVk040M3QFTVQdTKNeW+ESjtyQgKYTR/yCOYqLTkdmtx0hCe
Tf/la4JjZXCu26MC+npGItAQ5KnYHEkCrpQ/dCr5xq3u3CKA1lYSpIIcYSWQ
sizwpmfg6ukrQkZ88tRsVO4kJd1KwwAUN4cf/WYSHmYADU32us7v2bm+zW0u
KSmZxo+g2uZRDzF4NoAlgnFws+XB6tEpqzElzAEvo45rDf+XNk6Dta3LIxba
sXFgFV+iv4z5cs714T5dVSBQ8N7PjYdWvzPKt6UmHNLRe6xX6wsnTVpeVOFx
0nd51RG5GTWyDcms+3+frR4tR0QA8fJFASBjwVIxOl5yPs1yIqvEtUCKaMJP
KD6jyMJuS7iMKskHxL1AkKgX8JZ+X4958rMpD0lr01K/5a/agYBUNC0hujoA
Qz0HKamrUJGXasJ6y4XehY3zW3GeEGlxVQi1dydQ7mnr5MPiKKOyAwvhicyn
cOGMPmhywnXXf/qgZvR6NCBJ4PPAeoie5AD/Ff604tJrAitMA2bjL2qnjuWa
YHrlMhK4zq2Gltjg/JBhbShlTOn3ibkxP/7vuP5tC2WILVLZqnkg7suW/8DH
EYoYTcUWtrF09P2mNqJv/tVrz27IJ0cW8e12fUAmNIywORNw3qS9TXjRxK0r
j4cGo6k7nJtE+5Jq4i4tDEAk8TOFi48X/NfliICJVW7rM6l0Zz4shtbpVi7Q
3s5NEF0CdPqQcGlDbBytG+sSX6oDsVSVuLpPmo7PboU/rwTdl1UuhW1ccHtU
HGps3sEbi6QGPrTSxIfNwEEXDTVV5PH+iMA7RbT+StKFiSgWDW4Gov/l83Lg
Q2S+4HRyoZuk44nSInJmn8e9Gz1eFdZHrWoyx8e0adq6y4hs5IG3xcaOllqS
5B9CKiwiSKU2ZFUTSYEtgPS7+CQpYdeqG0RxcI9xVbZDOniPqSq4h0Fv54e+
QeykcnGNQU64ObMNoyl6MVsyuVmY3s3kwvNJCIBZPQuazGXR97AkPrVhyPC+
QlFtM7o8tmXd5DLqyuxxXdGmXmBnMQoGmn0aRITnVVTfhtlzdr/7xs+xoWFx
ekdFkz/wg82HI7FBJzqMcHf22DwMUJWjUJ+zu6Sm0Kens53C4GGUv/qdaZQn
6gig178okhjPfDms9izu8Bau1WgNkZ40tCzze0ud/t5DNF3xy04prPQQfZwr
8FpTpfZSCyCNGmquMc/7t+aJsQblaJ6EGZ4uc7Cw44aKkmD/W7u3QQrISk9m
sqaHCMfAWLlMzYv49dZdBxdOSkkZee3U86JDtjzVSfQgAVT7YHVTX5c4hwFS
N/3f6uvnin6I2x6+EdbY/lByADLdRNApCutANwp6VB+18QbuNv+ytrHGlINc
Rz6n+YV4D5ATFNIxQaP9D0gDfRkjnY9XLOW8zKNfsoculM//ULSD4Uy50mQA
xtLXMzypnX1WOMtSi9RBU5Of7br5eE/A+boehLhDCcOK3jRGl86xi6h8nAc2
GIzMMRs30NccsLCGL7iDqIJiR2DHS83M6iU3wSC1X3cul3ygpfdBu3B5C5th
xK7/McuHJbc3ykMEddJSzKhgYREyacuqb9AktGAH1plHNgGbPgkILem2hnpa
CewQWS8lJF8j/rAsqlTv6UUuuxJXnZmyxiELm1O8L2ZiTnOcEjrICdYJh+WD
e+efm3OD7euqobb1NU4Ff6Hp+WqIupZMfdEjyvGOg0th0CjB3sN4Sm8lFP7j
UMNWGvLSsX/Pyl5lpShwfhGZ2EyuGBPF0Aedd2G48d8QEYRdeYfmpQY5GxEg
w6A0etRihm9YuHbwc4lmgPxxfDVuoieyL+jdJHINZo/Lvw9UfSEC54auWZnV
W31q8zt5o1R+RHnVzwfjHeK+30rENWiV4ibrOx+pVOxSVj70RA/xq+RmipS0
RE+4Bu/v86S9AFbN/k0YtPnyAm4rMAh3qJBi9tZaYCMR0tlDJ3ojfANgl/Yn
aaneSKTTynukl6kKMQ5bkQbTci3XRfIerv5R4HCEOIGo8U1cslrp8Nqg7zMH
4RW1v71GhsWvn1B1537G0FuGxcw+qHPzJ2ry5JyEMQndqdWuhzzA9k4QkwU0
P3m5eyhP0p1QUG9jVavJsFMkw46shTEQK6S49V7tRRZ29SIt7TbjG0h7slpQ
MLgFyBIZbZdEO315m6FTdzxMNbVc3FA7VZcvzkI8J44mS8CghqOzVIJQMruV
rTbnbZJgG+l+BVKfWG+MQmpDQM4Qwtsvm70cYLZpVNDmEBTVn8/pPjHDSu7F
iedPc2Ju/HRdpFi5IiPyb+hyr+QWY9SV2nzG1PhKpy9EF/nArcQtJ4V2fXW5
2P8jtpGCfixsVN/yySql8N15JhGf6D3wgwCpDZF298XDd7r1YKKXCs94qy3v
CNYkacEpDHVKCzChtw63DMR6THd3WAtasLk8uRfGVbO2LwtFu5+N+feR/XVH
qMTBYHJtwPpYCYT3f8BUJGiCTc28uXwXVeCb4nFpzyLoFP6Vnc5J0fQuGjWI
pJt6H72c68/cw21AXGT3PqtzGwuXY7X/5rEkhKmYrpAfqaQOKDgjGd4Cc+WW
G7fJ3ML6CDFf8dBU2qcsleFxmeb24SvRdnfOyFsmopGz+bJ4xCq8/jgRYKEQ
dba2NFRFR6pYE+G9bwmuB/rGGo9P68kPNLDE4qYBEwfnzPj4ThbWBMtmxpfE
Wkr9lMJU8GxhgLb6gKo1E3TZjLOezQReLCRIQtrxe/B5FnKQK0+IZf5Vu8/q
yMTOjse2FWOYg+mODzbtyy7R5WKAU0oljOOOTBF15PaAc/f5Skb35Qz4p5Ri
GgoIaNtPcL2zDtTvyZIIJFqratQce6Q13J3oAL/lL77jVS071abUrieR9Ftg
g2E/G/iLZ8ghHYVfsh7ZirY0rad+HTtQW2nTxeJ4CWW8oiExGAqrrY1JV5sV
PcvbtCflf1lqW4fstWQF9z8Pj4mk6rBBmFRWVZJDcoSjjnyxdQoU2F2GDKw3
rGxTneKNkJwi8CZPeGbsyEtEuQ3Y2ZT2pKvNIAvmXeriB4z22K5JPk/U0h0i
d4tNK/Sw6ToxAdNG+jIJu2IaZYC9w3f5iL3PZTFLwx7m2FT2LSHpv/9cbYBw
U0flwawj5hWQE7cR+YN5IiYEijFFUHy8P96qgbIt/y8r2Jq8iZOvwtubkUZw
T0eU5BvbNLu6/SIkvhOnt19MAwCWm0ujXUL+zfNEJKeUby4ycA7WzxBELz/H
9j6WkdDrzcjzUXNuljSd0Aa8FXlZ+HX1hOLpcfvPAC+1rwiRoqmOYzmZAW86
4SHCL9HnNdLoh9MznqKUoyysVI97K17fzn4xN2MwrsbXg52ws0x6YkdK0CbR
q2W3SoNWvGLtAPXXLPIwcYv0YvucQQUidWB5nDOuuLs+8mh/jr9PzfJK6fU1
QqQD9wSdgvpK3vbFcY5AEI5hduphHWccA4Tq6/Lg1q9ZAAZ91EPwOUMotHXU
KYVjJbZzcnISk8c5zHO+Tvzq5l8IiebU0fwJMMW+lqjsAIa+sEq361gv+sI5
79pcD5FPhoQXJ9vJUIW8XMqYYyAu6aj4zTSJWDe+bs/ZD3V1olPF29wspDBM
XdCJY/VIyghoBXDE+ns+rWwWaI459WsIsqxbanYL1D+2jvU/frDMEjTT934C
pS9cy5ZsBhm7/OhtlEO/regILIv1XBnVBNeOihrn8SGhY62pUyC/6GDJcSBk
AmNpQTnA80u7IP5zoC7QitRPXmGJ2NK/v+CLLP/7y2yogAFNY05pVDBjDVZw
Px+nIja6bGYBbMhZw30Lc6COPr+CF6NhBhiNkW2B3y/9NTpV/YzCzBxuvRKS
5rLwLII5XdSTGvCtGgpTh0VuUbiCzkn7Wp7jL+GFWY387HocL/n7EeTyraWm
EjwWemiJtUhJn9AmnRAXcKIKa2GzHSBVD42D0vlo2iWfx62Yx3M2bodLT3a+
kWA3cHUpPA8mcaqND7hQSbEiBdWz+KvtoxTQaT54dTcF7YCSm8qL22fruCXB
epgwRb0yEUQffsDiUHWY+KvaWE5Pf74KlmcpyvQMgFNs1W2sZ3+qnNqWgStC
vWoKPhNuu6Fr+L5RAcDe0ZhhWDmt/zwlgY6r2CwFbFhYTzLLJU3L+zYofesw
3DnBTORO9KVWzw4L+Mt0yD7bEqNhMs4bCPSh+X1TuhBrOegafZ+U+V5yliMH
1Qw1vtyXhl5WSDrqOIkWd8j+1FmEZMAvi0hBF2qmMwdIYWntxADUCs5R0VMw
+OwsbQmj0M1ZuZW6FziNxQQzys8arDWN6cOkQokETSPn+g/C7jVn7QT/TAzB
L3s6QgUGOZ1B9tcD1gq3rdFiwhtYd7X6mEiR1aHuTdfObDQ9iwgpQjBBNIWL
hVnrRl+rT4f+pckXv7v2DMaHNVQzpwWojp7+fGlyxolYCV17kL0E/LgThakZ
2dSgW5MCF89yb+STjMaKip+FZu8TsUzaiAYWQEPKMWCd/wpKvGA4z0/f2u0o
Y5deVT9q9kyvv9oLEapZWvji7g/zRfmgrRu3ymD75p87tdE+/dmcc4mEJffv
eCRLcq2t8omkSIqzGRBMjvjkTkQj4RcDCYfAJ4CrBNdJ4/28Ei6n6im8jJUj
+h/f30FUYhGwt3nQFySERFPIhBeqmzSsX3SClN+CGTH0933avqTnyvbwWfpl
LsrZ3+GB3RmUH5ipbmH2UeJGKhxyl4J0lSsfbsF3clgcN5bjdOgT8IAfqN2j
kzWLFLEdGZ3SAW/RILzZ+CRXl/XqahqiWE7ajMh3Uj3adqIR5omrG9BAzisb
iiFTQyJ4PEG/a9gTqIDxO9YTL7We2/i2kXX613HIfL+AfsrXfiiGlqOcaz9q
WNHFcKaSzuXl+0DmYL8Zmj91Z3J3ffBVk7osmvujjhse5Ndq0UpR4gb2PRYf
sIPYXQ835RYYnTK0uxYS2nQkTkKejBSMd4UPeFporkLo+vh3WzYV1BIy8O8B
D9Nfucb377NHo6PO/ZKJgNNQWItEFHur4TBsYfMmHYsZyAMmrKrP4+KnZzI5
4uVDVsXR/TrfZy7VavZlFyBdgzI1D+/7iXLmotciHX16iPRda/dHfeH57fbQ
i27ZZNa3lNgRpZjU5anep8H/+qVIt97eBH2qelyX9W5xKx4tUyTxB6zFk8Wa
W7KFbujuebtFmVde+N1yPxKRFd29Lh8D4DMaknrcSCEMKsu/1jIJ7pzjBS2g
jrQ2XKX3kfYJ5ruTLfzSIrLSmEb18Nim3hqZYDfHWB/Asrfr14CG8zBGFMOA
ZfB0jIbiOH6aYl9Le5IgnbSTl5XILzRjLkSrtqRExxGDjRLQVcHRsvxD7Han
UTEeEt9vDV+tdfYECTwQ8uVDgHlMZAIPw73p4bCBj2fl6DwI2lZJh+cuWvaB
qulPpBKZxrOSJu6yOp4Ae5DLS8XCDzEdgjzSYFDg9p8ndzCqZ+ta9EAOnbOL
rdVLohavyATL4QNjToif70rZlY1a8wPaXe1Aw9ADY/Qm6DeNoFrTtFAQ+Qip
c1P0jdIxbFdn7Twzcj3/Hkr5D0TX7ZxAkq2nTHFVVUD/dSPYt1QZrmNj+Tir
vDpy2KOjclkxJXp0agRre+VSDy1LFST7sXSR4IxqSwPWVjmgC6b1ArJ9QPvP
SvnQ7aYbjTKYiGw3NguVfpBqzju/az1YqdYW34TY1JKIqLuQ12z87xBEDSqW
ul0syVhXUXlLrrZLlXPCejXk6bNaETHP9uaAFUj6co2nDjc/RyHsir8OFidE
GVroTquUT7EBELHy0/i4SG8uPF0WrOpzxRt/QP/gm9epcaX+XlNbKRS+kpX1
7MwNSnPz/b2c9YKysKCzwsdjaExDDjlgjXRtR3/yx+rqytz223o+dZUA5Ie2
9PUHW3AQQ/Y/fTUzPYkKETXGHQ8VEICFhnFtdNVbV7jC8dYaLBrAkAi8X+Hc
1ZCUgD0fK9+Iju+LVtkjXoZwzUV/sRxqrXEubwkBEnfHvekzbVPeRvRYpY8+
4d8iKWP+ZpLAGHtoeJq5NY1jMIF/R7JT4zZZKgjazK/P08Js98ueQ1pQDJRO
0Uk4iGqsLGqrVpHKZKxII70W5OEQTL8n6nw5qAk2wrh+K3o6j50FOyqruRPI
O70/4Ou+KwhZz7bn7g4ttHli7nqdNU/FGfWN1lyNjFyr6hv07yuBMLdK0J34
lFMexhme92jmDvgabXwJZJ7dIcxW+coS/rACkvAds+Hx1FT0ZLQr0UcBrg3p
eHY+pdRER+xVTzLd268wn6K5d36zsCny4V4ih3D2kUxyBBCnW/EowWCD2O3i
jmZfKhyw9YpCFJsBmbUcTzKspm8Iz2I7uS7nJXbpc73sechp/kf0HjXcZjJe
wszWrRCvIwVBIxNamWmxF+VwZr9H8ndQJ6+8URyCLAKcTuUZs9Q+zEf8H0zw
tsKT+lctUVdc1nEg9/jCKdEx7uvHQsIHLlrn3VHe0YTUvt8TWltEDJ744L5J
JhtemRahStEoAXoNg9qcjLdjzbaT6k1fKhp/6i5RxsyhhmL5Mnyf/4NP2bpS
0aTTLk+Co8uHHSgeV2lCgE/qoAAi14beXL0gJpSkDgBdis1eZxuOCzF2T3HS
S2AAFRYO5Z/J0/g/5xnY46ltLdY9QKEkoz+eDO/LADOynstP7HwG1JV3n2tK
YzYzEQrFQigewQJnPOsiQubnOLWbdjZVW+eE3mxPNzRi3xHHvLoZOxk743VO
HfvWtQVQyJLuxV5F45Iyy5d06pHPPB+jWL+YSYi4OGBT+o3kx/BxjG8UnMsM
+lgysGXFbpUn0j41wEMrPn7KHhvLNFHUs0MZVWNKVgwpDjG+bx8VyF+M8hoo
iKIZZUrcYPzV70aOsMUArV1BXB0UKcn4TZ+b6WJoLCa5PyQhIm3+PN57MRwv
sGEAqRI8rfLYEjs1Q3/VnS9/YmP0IIUnS23RyRY8A+oQfIF/heN3+3/W8EVE
q2zlCh8PgGGTZgTldBNhZiDHSdG/vieYvjqSZj82+HvpWDqaFfcMB/oJGH9I
OujvX6VPIszJ1Qt4B4qmOD6STx9IExPtxRVRht+UE2o5cizVcDc808HMfVBu
+BraAEPuL3JmDSPHpEzgjIxYm4LVLnOlYtEmRH8CFgkgZO6idZq17LBYRT9L
GDln3cSha8QL2E/AHoZprPNTwunEkTcrml3GKZPeiUvs9HAs1OYGyFaDtBZa
2VAgc6aURxyQPBYmZKhhNJYUAwPEmcocEETnp8et0+jUEIIPDPKfzRE1CZcT
eneqdBVhCTsjplu/n4vLrBAY/LdwSi4UPbD/5NazA2M2yPI4zAzaIuUw7c2s
tgg/HP4PJDSA2pGRcD4B5nc9FGxR2g3cGxlo68kt9VzVX86YgBAlYbi0wzke
AVCnFD43JaBPPPcgZABiVV76RL59pDl0KgrlRI4pslq62CDVO5qruEwcIOs8
dnDF84cEFNDjpFYwZndskpgGJb3Jq1fQuX77XZqGaSjIXSrsR243menMc8Q6
xxqh5Sc5w3J+nWGReesWcWBHhcWFzuhvC/FJhvyefGBZhCO5rSWTLngADpxT
SfcnVovMcWTaPFlsLqqJf7TZcX1pW0l7hAhBsEHCkNjSDagAFQGsHlLBxSr+
Bez+eLFqWICzBWECqxvCZ8zyRSfM7c58EEjQgsjLKh965Nu6e0pULLkp0+Ae
ieNkKd2zdh6FupSU/rkKK1vDfhgi77LexDNSQrpMnnMQiAsMHSTBed0q6x63
Xn/53ypnGiPu0PgQ8ufOYH8PL9yztgDT2tRHBCsJAqWb0t4nyDnygbPrvXT3
0fB/PCg44KDb1u7in6nLgJ8Tz4Em8W3TLuiyv2OboJAvTQ92Et2BB0FlaEDi
JfGD/CISz4wa62DPJvVzcVsq4WtXBPAOo1sG6erArYe5ozlQKgtQjRHojimW
4KjnssRnQJeql8mkTEvVxttBZMu85YA/zEXD0eXomDQu29ZKyeO2/tSggLdz
1o+xbunf9zJ0nTyqayT51NqTQy0RprsyrIgzpK6dVxq9kgBMxQd96njN7Xex
aGXQlq7lOU7IKRLk5axeRtGdiyn+nfDrZcx1eK9ALC/kQlXFU1/PB6NOPlvS
EoTwHGKaXRJDbiuhO96WpRKLbOcOSBo5nQgzcgx1HH0CH8N1cYUMZNJ8HfUK
1XCKSBnHQqmIi6gY9zq5/yPghDe4XfprHZqJjyhM04ch/Pqcw8rdwQLB2x2D
PczQL+hE0UUfwZK99bDKX/ETBzUP2YELp7zKcYCyiTeGFXbctJMAj2vHUqPX
48BvK+CbMoTMQkBfg2xOow25dduhKu1yajPDrWI3i/cq6EH8xhViOauxXZmo
Vo1QkEth/tVXmII0Bsw4mU52UvcgPwbz4JT86UAHIz3tycoN8Gdtb6VT+vSW
CrRmrAlhGoEg7SD8D/ogs+wogePZ1NPAysLwpzb9gHkHc1nRiIXmXWHsLRdE
5rbr3ZLfpvbK87cdO1cBIVxatABgH+bhu448wbTJ9tZ/HF0mulAaZ0WwB47r
XnfK66xRiCaBVSYw1Gt/05AIlVBRQJ4npojZ7xbpIGq/R4Q4plldbPwUdRmv
BtbfWOdyQY06Dy/+ZgrDwrnXuEIQOCVseRsSyZPsW0Fy017K22nIWUe73SH0
T4mAU5WggnvwCTCVf8RGksI+8lcRIUZDrhfX2S3xmA30vI3QTW3lm6QrfjRA
idtPMfFiwgfWWRcpHiYyjc8U5eKVIaNEKpnibSMhm3DwlJlEbwppGk3IiraZ
uDrhsoE+N2Fhw/0zbcd+CgvHL/oT2ckbZIdIRcrkMfDyqdORqEFUy9+kLw53
1Ssh+Kux2jraLZzaANwLKHcg+HAbFHE6u+Be8MWhW6Nwe7ipgTw43urOAgvV
SBRwjrpaYUtNEaVYKcI0alzNV+V0UrK/mmjfU4WzHiKvf9xPwDIsPDlnFCVP
yqjTm+YxCvVR0uKHro8W2Za0GGEssidzzNbGWMEPkgYb0cTE1n9e/YyRShvo
/OhWRK4FSHD2VZLt9NNdooAov/+DhK6Y0FZCj4ex/c3vxvQz+1nPhY6LqHym
ySTqfBQEVs8xBuTmdQ1CPcTqIt8AFTNRUTwEhMrO5u2igUM41fOJ0IE6v039
duXoBkO+uXw+/NbzfFuhCEvo+SvvmFk+ehHfZDAeyiOMArrIa9kqo5bT832i
cM918rpoEsi9qaLoN5Aw4L4Es3Kpit34ym4O/dZDirH3PePvmu6p9rpQZCIC
UoSC5BLoKAKjbbqLTLuzRt1lqJ1E8eQwo+AiJT/7ucV0fH8Kh2vfQ5VM6sTZ
pEl5Z0h8dW+XZ5NPqao/vGd5t1soa3sypeQaGbHJmrWGeY5yIoaJ75F1FokS
tMuInr5hUJCrsZZggRRtHcLWCK9l/5NYeFWbVjiN9tITMsAZPzWKwZZXJyTL
ADl6YF9fuf9Bo4hf3XjSEA6Dra4nmx2WHY0CP2B0Vs3BnWW01SvOrDaIWMA2
6NRiFFe/8FygomGDOsacD/Dl6Vhe38Qc8xs6pc6itY7icsM43zSkGTzzV614
t0xTbwCAXwRWaspMfD4mNQ0eFNY5bjAdrDfnHSXTSkrZplpMMdHnNAsbgz6f
qR+HMa6/rEOholwcx4CO7OkE2tRD1yrNhjDGWTHdBaHFJnFdwl/YnlsPM9KC
DrpWkFKekxrqiNqiozfbekDuOC91f1x398jmAqFwxMBdMU30don+SSfoVG+b
x7W5irQsamxmqExA6jPqIodNhYfDyocNPeh19OJGb01zOSgJnTY4otJxMiaD
hHmo21EpWnSI8B6GtjjYGWfxmQWSSRUCHH0m0Q6MwjjvnsOZGpvlmTjNZ+n3
hl9HluM7G56qS9jH9zka8d1GtHb1tZ7H1naK08yEL1GJ26XOFgtsNBM+9Dmt
KYBn5FgsgmkbzcSsWT7NboO+awbN1EmedPw+a0WGG/IC7ugH84X0GZWmK4Md
qz7yAEiPZNQM/XN3BKWOFrja6RyU5/G8P8CZAieOf3vc9yu/kFJrjV7BLYh8
3PMtvnXC2hPCcexUoO7hKrG1yybPVsGoXf7lM6kIqxRiSwtQ3M0MnwvcCtlW
wAtKfWsB6IoGUL5CL10hhXHtyOofrmtnc+dIK3wVXzDFjdwQmHMMOoJJYsvn
d25U06TYDaUyxZ779OAVEsWD+GyCnvUxsqdu9nL4bw9Sp0i80L2/hZFAEENC
gz1QkzcMTqfdVChRngYg8RwJemmSTGJW0+fMPd6U7zyNdCOF1MUBkK+KselX
h5GAPEoifmFSn4UBwsAbA+GEVNkq1WZdOsUhpjlkCxOX30TRRyZSYyWAA/i9
o0IS/QOo9b1CbE3Fz/DzoJpACmSc4iLGYGRSRvtbnUz4xSYQZsgKELm7Kj/s
XvDbVEcy3MRNQsN+TjDojCxs6nevW5i0PpYCXmYoCO5ODZpLNX/HL64rDIRN
2rMIbLKhVbbw1IjzbdkUDKUDYm7HoRoxUEySIHrXpxzl2QprubKaRAOHmDxT
4s8C3FbvHqezVHbRR8S3J6YQXEsYklNc7IrRqxlIJ3VVTg4mQ5gPX/IBBGIf
w+rDtB3ecdgFHzaYkpla+4OpSOlCvJ7pHBo7oLnCuqp9ia+PZKbHk027FOW1
sscg2b0L1Ad2HQ7Q1c2xTt5CsFjkRt50xnp/MxDoAxfHjsoSJkLr6UThfCiy
yN5SIojKmsqZQhC9OJiKZns/xgdOcXEsGeVQIBWRZ/Cf2dXqYEtKzugObB9Q
j7nKg4NCIMsT8OtYSjUX/NfaWgLr8T4epHMmq5/B+6Q+rXBkYXGz1vrDN2q6
pdGc3b2j4r/hPtp3Fe4BmS+VPu6BHeb56sINSJLoj05ytGzzbGccuZz5PdD5
XOdOuTtaruOCtHe6rGRiZXJeKTqA/ey9LR0dDPFgNQ+nSxgNDPOR2+ow7BCA
Y6KZZXF6d8NjJe5mkR6xZJFJy2SSLoBmYClVHKXZy45kn5kgxteM6L/xTjmI
5SexUEmcPMQytl24v+OwanuXDG5uQWXqq01Ayy/4UoDPY09qJ5Wlyi0ldcaS
vB7fCKXkvt5ogwSzu9lPX43vemJWsdN2DQMCNI1HdRa5R+6lARCmSXK5U1XS
sse83luj3ZQYyj5QG899/ZYxf9d5amFcpeE/l+hMhlADBOlXIwSrU6l8YjHi
ft6JqljKrY9HIMRw6Yjt/nPS7yPGje92oHA07oU5wSFPfwBc4OLmRl/kKO+S
MqxtipGOsDBlzx1nTOxHJG2p2S2m+r4qzPUJhiaUQ3JdnHxOsZqQMHvsaExu
cgaRiWpMNFSI7em/LZ+mUSSsDYWaPqiedXwmiRNUsWUdEEJOtW5sfwW/MQiD
1kgFmjexNT2SlM+Qls2zZ09hMBVJJ7gsJhM9KxLJNomBdRBeoRUpYOBGf3xU
Un3DvB2PywIwN72YLAYphJZUP/cRrN7/1s154FnBKp+nSLHjLUl07MuSbSnT
KIBPis+QWq2GFQdTczV97XkVqE183tfTWDjp6eBC9SCMpTY8GEC//6f5dr8H
3HOLCO4iyqAKRKbBpjtmDdMrMEFpeZ0zyJiuIa3csbP9iPYKEferSS8sBxWM
UlwP00L4UUhvConDGm4m+xJ5z8/fXqIGusZUlCt0NOMU+gO+BnLyG8gbrZOi
PeNDhHtkh7DppLqxt5mgjHZtFh/JVx0stWhICy9Z+1a+oAVJxQTEuLoKESCW
13HdXMAiSNtdkkIOJV1XXummK8oCIndEtDeSAT1HLvHrL/sPucaOD1i71AoM
ha2CUDL637WNN3ZcAn+Y3TEDiV2BnrTrdBIpQHVB/i0BAZ5ZbIzEp3LGOZNM
GpkhRUC4YNHmAQsAtg/SyRCKkHgW5YYAAdFPhRezKIYuciHMxu1fQSzIvBWT
jPY/9bNIP+ddoOBMX3u3dn6xMX4Fo0HRHKhcQBOOrYg6X1peUU7ZqhM8LfMH
CKxVQUTEAe5QXQEG23e6nKM4inT3Lj6Um1h/pPKACvJmE/KkHwa0MvysW0jY
FA90VxmiLEyr202tnM4K5coD1mudZ3yxed/FcQjuwg6xpqfpDoXTVt01ty0+
sBTvnwWQ5C/GYmaZ0bofupupVZDYm09y7tAoO98KyQ9dAlZuuK4PPT0PXjJE
UHGXLtNyA77ByqzTnwlRoQ92XJ9vo4uazduP1F0TdA/Ag8WwrGepmQ+5ePX0
prRmE8B4mGdcUtMTyLDcPCBp+4hkd0bys/LodUkLYnbTOrkOYrb3rmUEAsfc
tz/Banv14DzSuej6klYUxPMfX15KSeYmR9tcm+petboNgrl6hBcP+tFNK+4M
xfiVzwfE7pe6qtozChaosTcJywsPsdV92BH5PjisAot2f2UtxxmTmOPAOkdq
CY26csbxMRW6M/hxkLV0bdBoGtMFxEZFIH6aTqYIsa/zaekEWQmh9dN3Z15a
PX1v3XqiUFaF/SKwD7YO22e4krL4Q+2xv8b3y17UdovBqRpaVevY32NCUVw3
8U6V/xAV/fNZorvOV4SxrAc18SyzSF3/5pkCvii6lzYetgq+jgKwvm854EaU
rUMZx2GpBeE8jq3psIj9Dap5ghLCLn2D7qNU1HARRn3dWhscdxiKki0riM9W
ekN4uz/mTGlSsjQAs6QhTJzS4Zkqf6cIhlngvsrJ69ihBLOTJgPxQbLm0ZbU
f83/lmLk7CPp8iNRyxgAIiH47PTIHRou4m6xQy8y4qCFSq3i5qjhtM5+P0g0
qQC34O6iC9MU+sQGKbY4YXYKH73eLml7QoVLYqITA73OWXt7vVkUpWHWOBqS
Jt8A8o25B3hu/kY6iBQYmCldKglie+C83HnBkbte0FaO/EwzUYyf1J6nE/7T
H585mZdPeGG9x3PWOfeqUa35j3JVJIH3OL0I7pU8U6yqPqPjMr5q/TXfD3ot
f1/sPT6I4VTf5tzlpnnHPrFtI+OfX0k24UoSEU9j85pw9GuRpjF14GYfE9qP
OF4TlxsAlOSf7FHOx2/sEkDefGdilrl7TF7WwI1EvKF8UgUNeYDI3HyITRAK
1DFAHsmb9jUpgb/RGw3BvjfMTa/nj1qbVwYPymfcVJDeK/W8Vi9QNUwD2d6l
pAqXe9ckFimiHJn5GFTP74fQzBx3FUhRLAiTKcI5ML/r5bFDCpXrMmE+4kYH
c8cNlXTwu6LGe42NrKpb7eVmG2UGKqQoTuIWt1Ua6V6qbPGrcff3SHPmjJ7K
HQFWQ4oJPizIvwjX4zj6drOutcIFb1njBEQMoxBku1U5UQ8Hzkw0lZ174K6U
IXP3pw5aVORVfJf1yMmclEuzHMpijmoxi1vy5uIOi5HRE/RThJzKPLsr3TdR
3Fy2cYypxM1ABwgcQWY3k9ieokAmJNBlUo4tVOaakd3BFOv7ObuChDmcRBIm
EY4oDz5n0e6h3f1nuGks9ffUBOfynv28wJ9R67Vfk0Yez37cmJs4JOC2AbD9
xaBjz1FnosDWDipMVNRXxdoI0pp8dteOnqA1SMOEyM64DT97bEbGahNfCSCq
kt1qTVsu6Hxh6rMuNxcFnh+ka+atF+VlAvKO9JMh0SJzLeEEZmsTOFPNEids
sCGEWV0008pM67YkDXr34ebfyj+Bt8M82Futrrk30CXukmeBy51UI6EYThhw
tadcR0XokK8+VsoAxqUm90z6nWt1SSPC9hrL7SQVlyG+cdBCkSXmnLaqFHZU
DVsi9qLgIhOwP4AeG6jpSmR96ZEuo69mWnMe/81UkkOOh7RSNYMkt5x/jzdr
Ol+leoq9x9VgnE+0ICPX5cCCuYqsPd43hL2XvR+ZJm/TpehFzvTtUHefiOn6
3UbBq+cSejRhnPIKXS2Djifcp712g9kMP1DJen0LGX/03DZW5vVxgDMYGbbw
8p0t1aTVpfrjKLQ50pPZNpWgZZ2x/VeBlQYAFNfvM5sGPXWCeTAO/rPEC5ir
gxduCuDuetudTIZnutlkfaFrbGVXvZChBtNiiyigOJjXG2ObhtPApMz6Lleq
3+TuDq2cwowK+UIk/y8kZaCUxW5XLrjNN4JitlIrn3kdeADiBHL7I3i9izuR
0r9qPzifln6utBIj1pb71j8Ibkl8Wd5dKkVGoWUboYjx/0VZ6eANtshIUIOo
uX9yFrgnyGUO3AfUUwnE/emKd+aX9pBHie6t162dqtqU5JrEofz+zJALxnEb
P74fUXtwjzrYgsw2Zhb148WWExbo/69qr4JNBBqzQ3WAcS+Udy3bJVt1+whw
LbXLkyj5k/jXvZ9wWL9jxggItqN4wofeuvWmL0HegdUaU/U0NhFUlpk9XK1L
LJ4pTXFn6luLa3x7pIlLA8e04E4yaID8MCLVBMiEHBL9YlLLpCnMZqhewz38
wlN8X0tGQdNfoXLhheYYZyIvEGwYj2p1DiFnjm1Uy1wuKsKMApCwstdFl/s5
JfgYqOQHLZ9uW0QMQ3gnDY7JFbpUT/rQIZmrclPM06JfEz2suzaUcs1jdpaz
3IEiqI8Z1Rav0IHuExfjDugaJm3jEVLHlDHjVLeo0ulQrX9r/ZfNOYr6INsN
NADu4Qjmd9d1dy/T8jcZQC4VfijPguwphnswvlv/3JG8lPN4caminIXsqv4d
Ml2cezEuPUOJNuzSxe86+LonaKCBSV2ksUVZ2F1cyo7JUFDlc6AFgDp8HdDK
aQgGvWBdy/lF8a9Cjlux1G8JGRpTIb1QuMDQ91axdXUCjT3DvYsDfiABVZnA
/r2FZtzXft+lap4MZryOcjAmeWh4Mt2zh3LHp1cFRN/PAuPZ6o8q/0sCAHS1
AbkPKbXanmeF+GZ/E+N+PKQTOBEWCVOzVdszTD1kCfl8QdENkozlnDHusCqm
i/hb5szn5nhNvyvGbqYpKuKNA2qhR7ViFi/jCV3xONKhYsax/HaNt8CgFYE/
h+O916ulj1IcY+LCpt7PIozy5pg510dRY51R8oh5D7tdSPyt9s4EsIBFU98S
1PyVEFICb9TkOOAoKTWpn4TZCd30hT1B+ttID6oQydd4owlxq6pOwdIls61s
TXy7Slt/C/O8oehzexHSXOIajyePl0rUHZfWtaIhybfeflk75LANJ5wwIb5+
Vy7NTdYMrTU5/TykHOfkHwm/49BC0nmqd32OSpAp+GUiXRzOUyeE8tpFAUuV
disrSI8TGryGc9AO3XugvNKsefo0hTe8fpqaOJOx+Wxw0Mp+4oKFeKWBfo/i
w+ra6O1d7p7nqdCe7uE+42Xfz72grWIoA5JL2ZXp1Nkq/bgOfbmquWuuCw8O
oK2w2fUA01TRZTLrFuXZOR4llSTqRkGhtXQa5+jiCAfwnkX7csu6ysyQyDrL
W9XFDq9X+r5IP6pkKuDn9/i8uNavMOuey+zt75Ze9PVq0euVB7zcK7C8Ts3A
UyY2sr3uVfC14h38JClBo3NzkrmR0CcG5u2MxQxn6U7yaSPwV6ufrLuLGJVG
8usnQlGEDT7NNlBamCEPK8yCqRCJtz9ARY2GZXAXkqPl4BqtM7/5+NPrtq1T
j65uFbZT5Eky2LiJ7HIBxUFCYA7GpgmcrS0lXuw1DLNPHaDAD4z/y3sbJAxG
yoUqr1VaESZE9Qw06u+QPNy57rugdo6aUty1k91lH8y3JMRfaDTKwmSE6vyx
30Oa6NMqPBDE+YqderKdXE3GfSGPJD9lg40M+UnMyOAmSybEKgGY8SSeqAm2
x+AAsPDvcQ+vUmUnsYfJ5lP/g92t51u+MOg2nqSd9yWKuqUv/PtGqyuDbw3M
JoCdQyRtAkwZeOWgst0loajG8KYeG0o7hCVPLPMjcLhR6gZavaC2VtQPdEi/
wDPZo1fHeGkqY9nkisBkCajIQOHhqHhp4x1TjtL/R+ZZUIZyeTaK+/nhIQ9J
5y4mapkV9T6oqI6iHoLRzmLR+2mj/t8WYuysHPGWErh2kK908J9Nh1Z5BV9q
G9EuV4RkyDhRDtf7kNRiPq2z4TSzqYaXu0sqRjmXaZJimmbQgIabdTDpUail
vhFjoy3kZYZZs+SPBnsHy0Xu21VO1/U6vCSxlZkhjCfPLquNi85f8ON7/cQL
wrATk1SQzJc4+TQZ+96O03NVTCLZJCGYb/Kt92tvFeoWHbtvvKUy+dt9I1YJ
u/0O5oGSazS4i9mkeHhEG/nx6Upj/Fi8zzuTCK03qJH/5RB6ReLXiYg2GChB
sVsIhSakFUCkR5AQvQfiA9NDU/09Gw6KBQ23v6ioNRnbaTE9C6veCdwb+A5q
KDOrarpYnciGKEFBkLVRj2zP40JPLirDuEmV9HpnUI30oTdsEBIlpyjuDhVd
ge66RYgicKHrQN2g6cWSsGYLZEasSmHN48u7eX/QyME+UjMYWJcb9gaGE5OI
znxA5YyYDt5T8tDMTfwYTH2gpNxbVBBlLSBNLAz7iTuWEght74NvoTLtt+hg
QRclZaOND8CfQSqqsB2j2DwQAIWgb+6xvu4qsjkfRW/yoT9ZZLqmmsDKQYLx
bzlZom1LPddxCLHS8tNhj/VpERl74kFFKs83MTpiyQL29tI5vAfT1RCjAZDW
sZL10SChTN5i5wXbE6+IiYa9d+stKsFKvdjojHo0CB60rO0L21NBvpRos6Y7
f70+7TYKF4KiwgDMIVE/6nwZ0R1WojlJyXdRifCbxvKqWD2RUHcz198s4dqC
hvFhgmStnpMIyil5AaLgpWjaNC+IYQzlSCXgHz1IlsmN+Pw4g3+uSrrtDXVM
lylkMiq2dtS4iSYrxBW+ncc/cdXhKIyHPbe3r/OPIOsf5x83FzTqDvBJaQTO
CJ0w04dHi/cwFBctBTBU91cwf3b+/ITD4Z3l1NKnO4D06LXvMcUke0y2xV0y
aP8M5U3B1F12dyMbwNs9ffel9Ss3BNr2gt4DghN4tPkYtcqWqryIMHlPXPUv
iOOSGOU3r0SBRYh4UEvV2A0+bUVxuSXdUSzBSf4ZsIgIxJoDWX3de2OOM/Tp
xoZ03IzYnl+hlb5RmSsKzzoFWXPljh/FobP7vV0ep3YpDFd9PMRXFzwWjWgp
jzUjf3cYR0djJ7TlTTOJQINPKb47PZDNsYDCJf+Z9QdZGGMs09E94dBSJo1F
Ou/0rRGP3Zlt2bGOMSaRjzeYsN78mzwQJwSHJoaCDucgcReuu8kvyB/ghQM5
L71IHdyt8ZgQrKBE6pGI08fVC0z73BiN1LaQknpI9ossl5NeWSawil9XCdT5
5ddDAvHemkQdvX/+Yl4RPeaX+4C5dghhB/Ds7PeasAequ0TSbcMQ/zXSgZjh
f9H53aor94BnQsQZChHFCyVvGd98rI31IU1dBq8Fr7gaVDB2hHSnBTSdrYQq
4FtDVDaYmVZwb5WBo8QG0CeuGNFAO6ImPjyb+SzO/rFvpbWYTSMWAfE0JvgR
kIDU5Uc9FH673JadJWooM2KalRQkaxObRZZiHdi8CGfDCGUl7043ad4JLurI
wcsDLK5O6l7GbHZcLbUn493PsHhn8YTOosJgVfKf4HDeGlkLMhK7j/3inNat
Q/vJIFgdqcdJfvBRSQ8zpLZu0dRoQbGV2TPKnSXbdo1l6aWXvWo2ylGbsRB5
qFbm2xVexhgjtdKjQnV6DPLjgjC+GvURQGE7Jel5rI3uxg/ha9toCPaEc3jX
5z+brgwY9FIqnjAoDqEe0BNeew2EeSI1nE6s4vh++kUeCkwAXKhU54fqkcBQ
8AyB0sxtQf5nCTqZt5zCMYRJx7cs+nfnaCsjbTd+gZIyeADMXJjSzzV2ciMe
56CnL2yxlc9ABh+j2OWPWO8CksZBPkItTTSwnimhvPVIusVKbBAO5h2c+Nbr
LKwNwG782d8RoWaqn+PWuHnFnP9j/0KXUl1fTWSBoCjRrs04ri5kOJZ41xw+
0vfL+1QeQby4+Zp14Lhqqpn2C9hwdZc1ihfqOGoazXxh7mdhtESzKix/IX+h
Dhm+pSnamDJTmGgwICWlTqoif846xoyxp4kpF6FvzXsghu+t9+KaQxmmj8x3
m+vWjrZvezar450iMDgHpnH0Q+2SLMrgEilxkbZkLt457bjGWP1GKAKnmmOK
KjwU039SYdWTT5XHNwzNdf8lXbYslBizdIO561ez2RSvsz6+4bFt8wKlqoT1
g5jrHT8wo+6FI5VEVyLq2ZgcnzXkcUKe3hgbobXIGD/VSPqkONQKAY7MCNYg
yJni+6mTgYF/OWkKUan+I/+qdsv+NSwVySj5QP38VqIrTTMzgUnsayp/5pAE
615x2GOpEL3BDxplV1BUxbOyeb7qy58rTQuAicC4Lw2qXOY/QwxEQdp6Bgeo
6g3E78xx63V6zFGJqujpx78JrP0msDRYUzlP2gGIiQf8Vu53iMfM9hgEQ2bf
RJYiJRUCLqN74R94CFGM75G9cqx2ZqsQb/Q0yGxvnfobFy37zATczAeZO1zq
jkV+NKcL3dXlp5+WLD80y8cSUzWm6SGc031naLynUrieLXmTavynPQRIaK7J
RnUpT51GXd2OYWaSHrKaDqzd+fc8nggDARoeP+qkwWObX4Dp7D/04SCJOtNr
5Ye+U+4JYmfIap4SG3kMc+Im7oi0fhZvcg/4csShQqs67Qjvg7qysAFDPTtx
Oj/ES7Jgfrpjk+L6wyQeq58tpRGJq/blo+x4vam4E/bivY/ukv0iiwGbuLCm
n8GWrvysP1D/kMK/88wACe7GTX1FyKXjZttxaz/N/n41CgVAwTOYNQsaMNTo
krGnQuzLFTwdjqIaMLqT9/vdEINnTfom+ASbhFEuHFXLp0ZZs1xYtDS06uSo
DAxQJhrqhyvIwTFsQMnP5xFn/XIqgu82U//U10B8drVjCgE1+MDTf27tobG2
8QKGGYOcVofSB6Bfz+49Cs4d1qBFEXodQjE7yNefF1A3FbaShdtcMJsx1PmA
/nJWS20NvlonOFwTemqpw9CRowzQrnk9bf6L7pSE/ee0zcgxB7FoAjoJ+76n
j2gIB9HEsvHfw3BshK0Va1QfjNO6oXZHVxGB82K3VkGl6c/z8sbe1Jzod8fy
m/PIcQRFCiOskgdPcHc2NoQyuvFHjJPFkv6FGQ0zlW8At358BCEoiOIC+SKg
4PS/9M9gjFDghZbGt5VNPpMKZpBW9WrwgesAKMc0NCnCeFQxAf78u5al5z+i
pn8A9huWS4XscG9VSI03DbMGqNG47sFa8LeAzXDXNGWcJYiUZBcUZujt1Okn
0rWbCJSJ8orN7if9/Zl4UiCZ338dXKdBNy/ZoHwGCzvZEmrFlSxB4ZaPaxyw
etfNMlxpnILicFZ5EmczO77wgH5sfNFryPUoto3oh2tZTtoaeaZqfmNgpPp2
U4DK6620OTcSPi88WtBB1ijeh4GOuUCxNmQufPuuxzg8lPHqyddDwkQLXIq/
I10kzk3NE9B6s1g7NK4RGNZScf4QFRtMxC8OF01brfGwZcxUUHHLSj2Weyud
V0fbLvhtx/C38s+xsf9UDDwYZYjfnwYtKTWkoISHdCPk5HBA5GlUbu5euod1
dhvGyHIDnDwpV7lp1uljaMw8bNdmbn1MehaqGBgU/A4ZNb8nazsf3MH280Fq
QFsDUOOzojcOFdVdrWxS3wrnlfwC5nJVFymv3yhR/ZY3fJ4hLR5fmsWcpoJ+
Yhpj7ShNF38W/AqVf2tVkIYnz8N8pg2CQ3eGPDqo7KYd8hYdFe7dwMc9KlMg
ZbrRClB7hLYCrwfqWdkp54BlJg2ZJ7ox1PUVcVTgydStICEy7KYoz7k2UYgV
XV4FuJ594AagOMEPdX5O++9v3pkcG6HK4pijXIvFwF3J4BW9FuyqKG/c2Epo
qHXOysQWckuGzhYNRU5Xp/4zyNPyx+/vG9iaj1QP+XNwnhXG7kd497GWUKHG
uFpPjcAssEbYo47tnNtE7z0M892/MQAVV2uK5EXYA2RekV/1WmhTqHq1y+14
WSLGLIn9QNgRQ4OjbE1HTfBMEipNKK29h9G5i7uVNj5E1rz/w2Aoq05sQy2D
UKSKV6c3zLmadJVZUAgqpk0mJC6FhXxbwftHGrs5r/t8DIC5ewbbboFQqZ9s
WZ6pjfTG+3nDMA7f/bzQoKAy48onKjW9ohf/CdTbBW0NeYySHMjKv/y2L+xv
Ev3gJUcqEN4Oy9p2JrsEiElv056MsjTZSOfivGT6kaBgv1gvvRrMZZqlg9vE
Vxq+fLhUVOcCs0CVULNn8z+SRmK4llgt3f1Vl2D4E3zCnQWRGnNrYm9Scmim
y1J2ErCBo+Yy6LIhYHlxbsbW6XbjutFUPX/OWXULQ47RAeAgd+wC/CzMNJ4L
u0+reni46WwkN1XRsgO5lhK+XiuxUd0d2k5Y9OtCP1fzX4vk82WGHyY5eSeA
4lvi5ZHL0Up2TTrdhUQD6tMHDK2/rL4/KoC57Aro7iJDpx83boFhaVObRWxn
xCnnwFXjclqlJ/bgWbWasmL8xOEfj4roChxYMgU7KhspO5mZp17BodnDIPC+
y7r1xwlK0ZxjFv6hb63WrjFSHWccKIwxf+M1csaAapdgHcVtK9/1Y35Dp4OD
FyhSv3vczb0C7MWw4SyJ55PzgUJd8hxmNP0QsQT3DL3g9/+NuTdnkGhJcshf
q9uujjaQdDFAE7X8FMjrh0VANad1nE881e9+lutiTFYg3yB7nZKI8ZpF59Mz
VO9zDqtc9z04i5YMPMaCRzjlMGyJKK3lIwLyM2LNL+u9qpmKtm68hWJImSIz
xvkpDfXF382rw1XVg5Swwq7lQt+F8xA43WLxAKfdoxSJ+IC7HE42NdnyitMm
nAZIBmVrpCihHt77TKBizLaAG8Nz4t9TR/yOxbURh9+JjIu90f3LlsiO7q26
oeFuwksycbzpue9VvJvRZJMvHJiCjUkcP+rjWQZXhxc3xrPgr7TAxQlLqS35
ibezdFtUwgrc4eZTx5BJsdMB8Kw+RxMbBQfRtPXblKf8NTam1PFVOxflpEPE
yY4ePH0l4MwkE8y/X2Yh8joe1CBlwn1SxgJf9poYMG+ZrqCZJFIpuUnQ3I9P
OjKY4Of0deFXA5i5sUPZVS2c+pmPbX0ryjKDifDy0Ke59HDL/rnChhc+tMKh
jbvi3mXfIgLHVv4MAtj2saLWltj7oNCG7ow822mdX/6ihTHM/adA+0qo3we8
9W76+iAJ3vnwuXsbaW0d/Ru8FVnpqv4txuxruo6AnK9Dzjbevzi4lMvUzVf/
/fSzQgUGjtofAvhcrEz6kB3iL+qdEHCVqb1r0BK+zeok1OxUudS2jgPPhIH9
OeA7RpSTkPH2U3bIqMzO05S+CDP17cTuB1Trz9fjOhwHioRP3/MaJ/Ot+Pgs
ZPXVHhLzrgXlmFNmzVe8GxppZY5zO7ImfXS4UL3CE1eSYhh01RzD8wq7yCYk
chktfzfSR0jJ83xPqioVOdAwUdJp7t0Kwuu/zdp8dced28YcGiu7bwUt9RIA
wdCc624tGkmeaSibSDFW2YvSCte+9ff2s9aiXUTQG1W9MwSL+5PAS3m4TCLh
HqftSQg895T2A7PUeYdFtMtMtOhtGcVuKdDuB58SWfl0d6eI5ctlyHLmZ/it
CD9rhYM/O44Sm3s4UrFbR+55eKCbky7P2vVpmAR4pHr0BuX2c975VDpCjSBF
9mqZhA/1a5ATR1hR7F0y97Pm/IIb+7xqZ/IJURIqFEFZB8H8F6MTSWpcbLOW
bryT3o5JvOaCJp10TYHue43bi5Vp3ECCLCVpsUSHjp+D8uR2Y4UB3K48FBHY
IGgZo4nfUFismY0977Ur+P/k0FJ5DBDFPejjEKgBzd+CNJN5Ho9YoZZQ66a8
r297FhN1GnhoOss+l2+N6OjnvlxDgKc0sTplB6g9wwSDH6CSrl0dnFT4iXfg
QAtErjm06skIMir+DBJmI+iYfFkGVwsywe8DQYNOeAY5FkUVl0r4prl7Q3Ar
vyKyF9XkECSCtM/CXwFZ4PvFXSe0CWkNc2/P290rDqgE3V6oJgHxPyvvNNav
ZmZTtwiQJU06wR1tJsG4BAOTzjK13BSDZhF1WZpOqTxBgFmJce5XmVRczs51
nkPEX38fMLOPbuPtpVBVtW6yKbypuixTaq3H1G2AVqBsU7RFdxnN/QSRXtda
JuaTrQwY/jHM10EbywJBQ3LBUVb8MelIed2YTMCBAtCP2sU1yGG/MY/QjFxM
Q67x6EA5YeBg28ySfjtG63lSxzo1fM8sSWz+N1ennlCFbLPxcnDEUasj9G2G
h+/UrnfhTpt0UXsD4O3fNzcdrO2UjxGYZErCnbg+DV3cB6rTKQwzbLpQGXP1
GpgDP1rKqidEMTLOOoDYKwVaDGnR4a8Cr3lmOeYgHzHt8P33w9Nas+ieVfEF
hcRyXDKK2Y1fHLjdUmyRoyYZItYpq76uYOU1kSHQ3mXffv3GNGPK7fyqfMQL
cOPhhJJWp9s8lJmWxBGIJ5HH+9aBFlZlu8x12/nAUGoy+DQz1Ex+VlIsFONk
lyUYTiwprYvBKnpG3ZnR/mNAjtDBpUvJu0qo03gu9Lnb1RYvt0uAouPMvC1+
dt8XriYSv/47bDc0JvnIwxLlMtyFGBz8FwOdnEoVtf3iK+fMpp9iHxc4Eyx0
4SkDE4V5IkE87keqXOFgJPCAUgwZegu5Nh5B080zAW1PhfD2iRHvYd4OeTCD
JMDYM4LgWl8ASfbNDBxsUGbVzScS8LZkqlu2L4VuxFLC4rk8RCeU8iJfOORo
rL4QBKraf8fk+DTvy5xpKvj8GCAn9GwyG95+KaVEBmuUsEJD+s9BB8IYitE8
dRmwvME+C2LxzonUI5VHZxBVQTebHipXlRctjAPby6lD/Ph46YzXCeM3EVRU
jOTzYawLSxtcFiamfrvVbhZKzSLvJr28r+dha5WIXY43qAUbhn8YXp8s3qSM
eY48L29oOdpU+2Uk2L6LbxwQDaDFKSd2D+UBAEeXt9dcgblysFUZSKZUym8+
mcpU1o5FRHaHEgVfdPM4zl+y0Xrye6R0WzgS2Bb1iUjrj4V4M2JN2eV+3inQ
96GeASh5X+ddr4nZrY4yWFUbpbHe9Uc7NnkXLhRukdgid8O1I3qnz+PuqxPk
Vnc7lkLPp9aSl58FqBFvjQ6Vdrm8pWJpRlfuXVtQxqgE15fm/iNP/5za+I7+
Mmm34oN/Ljfof3I5CZNU4vDOTgOpR+7Kdh3mDaHafa1f+tHi907YXbvggmUa
MAcTv+TFeflNMUY3vaBlW5wJ+/mDfmPTi79uEEJR0rL3pcQcQGxZT+GmEpNv
AdhsHwVKBAeZeW6CXm4yv8BRYLldvx7ixPH3GlxtoOgqCVtjC62gSagMOT3a
LUbA6hw/3/trS54e098RElfuSx5p9VJW2IO5/2O5FmXvmN0JN8eQIF9Jn3F+
366WebbEfGSA6KYVKE7sITUe+xE/fkkO8vJG2aB5qITk+mTL6y2OcA+y1gyJ
wQFLcOQVIpI3nHbdYvRiAALEhYGuymWPK/t98w31CddxZqj+cGjck1u4yfUD
jsHCuc4JA5jjNo9RdS9J0tu1/mnjKLRZTyc1XQUA/OVjvoG7fvLpE7RUJeKf
vLD9bYjcrCMPhyK29TgxxtNBpWTrnuhkKWDppJt1vi/h8zU/YHeUlgCaGEn7
YPmAH9sQOghfw9P8F4SkULTMmiCHlKT/5Vhla38XTTkPngv9TXNPcTdiTVBT
gehSyH+xLuU+C/9CFTiSU9+RxpT7LjhQaEAW2DSYgXz6v39FnCtXWkIt+14V
+Sdk5Jiizvsvz0wmIB3KAaPDGLQSGvz1l1bCZr9TYOM/WQVFfom/sjCeeetA
T7TeYkHxkcOuWrzwd6Fk5DM+EtPjeKqKy5lW125Wcjvsyh36JzKgmsLhrX53
r6jPCKt0d4pgST2la8QmRPXVYg+DSbVF1UnN6XuQL6Tx7H6ZgZyOOlN/MhIF
pNaeY3yISNeUAkepeRJvV53GMZZvtXtii15kCCw6t6CmeOJNQRQXPvnudGuu
oPW7jtyEkRvBhCuEgplvskop3EJuMbDpqotZ8M5sDMVcq0NtwV0/BjqjFR+M
PCCbYmzI3pQcErKV40CIktGhNKRwvBMmwPu8nY9Rw15SVgLQx/bTtjccGP9H
iveFUo/GaGZCRxC8PHRoiamUSmvyvNDZDoIxSrN+s1F2MwmxuqbnO5uAc9JW
quZ0OTvsNQ0RmjJfp0IXBX5ErLQNOSKdU2DxYxdoBJPBfqLiKX+bRaCiUEu8
lliPCzPgj08cSXR5JKIgaBvvOi/scD/O+AbixNSAw3fvFkY+wQSSNWAI8nKO
TkI+xtQca+wuw+rmJAhMyPwqtw18XUQfFi+X0dv1EzG8fT4Bac3KuBq6qLRW
6E2Lf1AI4aXUzbC3N+jSB1AsWIzG7eXa72auqV+ZEHPy1TxyQ10FUXxde7qS
KUgKlxt8MimazqNY0icLmUjuU0XvBrpf4mSTGm6wfAdDzfOv3Vjb+kCoOUq2
uBL5suesqHhj2gqxQBBhKj7/wyGJGDQpBl04LgtyY/LlthiO17jCggONyDnC
b/PNjTWJ3oHwaxDR49xdwKKziO++bkEhk2fgsWQ9iN5EhGniSC6ftITR2nRT
TwVZHkBjs3D2Pppaull9ukG9jsGXvSapJtNG8ToibJ2AMzLGWUN9ZAwURhy8
7FytXMaGh4VyXCkRvzzHywMQmzYBaKYV949xshfHJO+R0wsfhmPC4LGyo1IW
kM4WBHkgMDBcF6rFf+21LN3ogecKHwXphV1IFNOArvgyqIBw4Ns0e1cshVK5
m3lGVvxKxBqDQhiikJgA/+r8hX4PwyN/Kpn5V8Dq2GIl5Sap43VNo5n6roM+
3fohhku++kmK+RcLPPr5S5m2DQV1oItYsw6XXp7sObVqkFfXlRCq/MqXNpRJ
61oMYjDdmum8wk2KwktxDgM7/fZROSs0P26K5oZhoxxLMX58ELHj9TMJb/st
Qj0qRpOMjnlY/HggNtmefm8oegZdNFXgHeoYuGUvGibCPSxj1RqgKgK6P0fi
h4I5sQbmt0yH9fiDW2X3U/MM7R36hjcsKuN9hcT1Ze25f4Sfu+To1o/jcTQa
TprOvEbIHWMSrSRa/wRt/kF8+xaz5iHk78ZJswmRaM/fd6Mi8I6NE8yGTIEj
NYvO6xG8lqUO7oeiAuMkVZ6/6E0Uz90na9Ah8gpBQ/1b5vaXb79Xtn5mmBYU
jiUiLiVdWSacWNv7jdY2o57sCHBAgkL7T15uQtCe41V39aG3Ez/iYHQx92sR
s1+3EsqcPEhk18yycOJJVMTFZD/dQ/KmGHYUi71D5AdgBAIVfCW2D1WgTkx4
eQZYN8pJ4hD91AICuVqsSYAIyhiUYIo4cXd+QWvejc6Y/cOdNoJeZstLEz7I
PwjJuUVHx95KZva13mNic9rpKv0OqpfL5humCCjSMJIBZc+ue51ULpp5ErLx
RzINlnW5UqC6DjL7BLpdy50nm/ayAbcNpdvsfm3eB9Ii2YAaRG5R++4O51Rn
8+0GAqdUcc/eXMLF+Uhe1bMzfwc+MRC1Ds/ExVggoIGakzdyjRHMGqLEvgqU
p8EjGFngrvVL15nD2VPWHTcXC/U2dxBpEuc/obm48g0qzZLQP0aB66y4+RHr
RKTs1PRJjd3eOolMfFnrY7zOys/njgYkEnj6ptOU7ONF4QF8N+iq7wDp28TV
9QLx8h3yjm3Fz2jEEs0wa6Ow4M1Bj+rud6v/sAeCPab0ZkHsVinoaQChx4yP
8rIiTLGJaO6aDpcDU8y2w3La6O1dv3zi0yiPtoIT+r0ktIKWlOUORLnz+vp6
rcgjqO+BctLaIEz6Cx67vb4WudSLlrZIbAghll6xci9e7UauEB/D2GlUNlxV
Lgl7kcOCqZ7Cw4cOOsIhkb0uqJtGb4zIAP4OGgpSo7vTG8qDd6a7wsRdnEXs
AwbD4kF9Kubarci2ytZRBlYI8wg3xPe/U83qCPy6ksdB4hLW1Luoxwpz7g9a
bprFgQR4S17XTRh50FqFcJpfNe/J9hYrcoJVgJZoEwy5ajKf8HcNx20HzVpg
Mk2PPaygcp7TLvgmDjmK5rJCe/ScREyu56+Amfia+4RFVd55junOE1ahRE8F
tMoKnMcz7gJZqdA9gLOyqVHJ1V4gO6cceT1GHnt+/PllutVX/6NhPGwvxyV+
zkHCKAq3n7UaO05dLi7R4OaSCejIw/UmYQZcO6CEZ9CNYgy4kLuUclTetz8Y
my9zvlE85jws5qVmoB9ut9tn7YZXMVqJCo1nTtuqG8NSOcc2D93tH592TaDa
QDAr7J71RO/N2ZDkuo/yL15Jq3NFVgo2v2NP2QjghJilUGZ7sqk/3yEuODKN
ixER6/+JZJ1Q9eGyfRxIgWpyAGAZia+XpdxlnHo5JiWaG2sd9GLO1H2cbKNf
AsnOo4sBKfcXNXhd4MOJDDp40ME/rR6FgCC7JyoikqY6JGQcN413/gvDYqHU
kG5M0U75xBRslN0qRhxuZrzmiGMHP3IDZV2vobMUUCbwWDc9BdVx0Wfur63V
mm+DVvemDE7SuJrlMd/qi1P4B9WBon56SioO5aeWhu/ZokgjuwpVe44GMqun
I0KhJVyWDk/pki8g6oGEoc+GwJx6yFubUtV3TIwEqLQlseNGEx94FC7DpkRq
alSiAl3yju1vz26AErOHSl3dwAe5x075ubiB+3vbbynLmrj0awkLcQ1D5mby
A39nYOceNdsIg/z6JGoE0WxtacSgZhvwNBwCpb1wGCAEH1+VPfvmxoa6NgI/
+YGGft0fnSPFJ3hmTBnwMiV5WblgInoQLZV4ARDnUCVl4Cb4iZSAg+rsrl/E
BiDDxlKLzCOkP0C+UEv9dHzPF1OFzWzkNBNVIr/jjiQ/045E6PClmDdjPDZ/
yp6DgzEu3Ojd7XNvLO1oJBZoVxMwuo8l78fKqWIX45g5AwxPUKB5MYc3V7Rc
VolRUlU7j0I36F7fBBqbtxYyfLLjVqo18/O3maJEMCgH4qoH+5FZVmYL1the
9glIHIJNnNT5hBgSk1DNDpe+qr/9s7ErJIy36qOP0Zjqx1OTXA2zEBMbWtNG
DF1c7I/lkzMWrPxe3sy1mbmLe96VNMFKJs3Ssbf6QsPbPl8dANRF85gJ5wOv
KK/bsM+3SjIJ0gxrF4RL7owbhW2+5qwxVSp4odpC1v1EBS6twn9WRqseUa63
tui1AuRvXhrF+qd+jtYU6JcNFJyoJqQsa/qNRmQxOwwXOUGmTQRf3PwEJG/N
ZcwvrzhC7Dg0gY6UtnPQPfV25rpbrZIOKNr7vIf9iW3bkjDeXSc502xNC4Vs
ksFRDBEAbAA0avtHox96JF8sJWg0IhdxwnwXn/HOUARF2DNLx4J7Qfb8tDIm
5sUlSCBFkE3oXI6tqNsgwB7e7b2V2PrkR4Rb/4UB4ZKNeM4U25d+WjB5wdVm
OaLIklSkzF0vlyPxdFmS4o4BkYEsdCCRKPVsGCINlHZ2p1Ou/Mt6lXAvMklZ
MToSGTl5p2Rhb29qxRsAfYP6e/kyUxthBJ4e7cejnk+B/Dw2SekFQoPCPamg
mzP2A6zhKZT6lKOxg8FsAxmnCEvVjuAJfs42cNC4AmtPI71jrofQvuGimtw3
N+n+rR9eBZhv39Ao1ElQ8SptaM9Wh/ggM2CJhof/lHhyq5gbTiNn8H/8VGVs
ql2/Gu64zJFFQ+klAfpWyisJV+bErc5XvGtiLDQbTL1uXd5QpqlhO4ZFjwQV
LjoHDI7nuvIMT3B6R6gt5L1e14MikWhycUtjrl8QvneIA/aHKjfRTLpo9u2N
2ptJmrNaS9rTLEiye07Bl5eXjWw+P5LaI3IU7N9WB9mvXwkLTlMYegOdKhme
Z1eYpNm2N/x/LLPXGkb1AC7RVGml4oaeBNp5ovFsW2Hx31nNr9tHG6kqDguu
bVkVHf1swqYedLsRO5C4CdpQG5FsfgoEC0wCKwxgUo3/NfSfz2Sr7g3nFpS2
a+H1dyT6vT/7atI//ncmr0uOkFNtFO1KXY3VyxFK+E6pOsjmwx0h/gSyeMD2
YEodQY/VZdZibV0J0GvwSoUXzd0PI50Jy1Ht2panjHYG/7RPG55Djvrc8imV
amCfkc10VTyO2Dl3JOOimzongfeIYqvywZSNAj9d+2GssEZDMG0xaDDsdR4v
WphDygdBq9ihaWn97EQKUbcc1PBqxKXrRk5eU/usdoNdEJiL0bo8g7Jll7vJ
EJ2MupfWhEP29OqAljfHRQRfn1HAv9AqjIM2jLQjA9RAeRYx1G1f5LA+2zOp
EY8CY5Vcjo5EQe2LqAmvDrgyVY6W2LmxnQf8Pfe0+L0snRyVmhH/+K+hMJHg
gbO4ZmYre5XmyjkFhka6nzu/zuTUEyCQa3RSTn6ZdCwdi8/WrqlOL4ZICJJM
vNh8B2OQ9tFUjDaZHyJkmgdzqgpxKOU5FNMFbKE8OUrZ7ohoylERvcw5nzIg
eo2mtHIeHT6bVYJ8fxIib2S2Q9KMwQ6NAaO8hEgE43cTSMYB1FWOf5pHdaUD
GpZXdx4pRoj9D82XF7vAsFv8an7LWXuxoPvacEM4w1+bbDY3qAcrJJy9VajZ
fxYeNGt7tPvCQ2trtZFh2ekxMDmviKR1nYrvoWotmg1zH8ccD/OhouUO2Y05
d2V+vElQfsulTwWUlZeW5JSeCUH1Fbl7NyugR76d58sgDVh7X0jVKtQbE9/4
QxJFeb1jP6HsKKWEvt3fNBoMSGnPsLYF7haFiFHH/a0oAqjj6o0wDa++fXRu
xOKdeEbx7NSUk4qiX4fSVFNoQOK43HFGXsTsQDgJEN7fIuQCH3TLnqo0eemB
suKg7A9RHffoGmmW4bGLhf/4ZC5u8AUOmep+MfChxkKB4lCFu70MDduEbKG4
6ZJKnUEMPvOpX0XUeYO76vOyPCVAPjOzetAaIoC5Sd+faPsu20n0PWnRTcgA
jolKRvWsaQgh73av7CY1/nONljuKH86I0yT0A7jI8bH5/r6B3qvBhfxvILWx
jVsOZcuBc0Oah98pwXLhsRnx0YfrYRTDFHOeLTg+357jMadbRBezER3ZdAVd
/Z7acNzVkFXFxyulq1v9aLZfHOXm791Co5wO1ARJPfqn58ji0r0d82cVtzDP
nYYdYNk6SJp0wK/72wc9mKLd/KnnS+BtI6M7kEpz06v5SK7w5RU4qrD21Axe
y5khWpbitBlxBnpa0hniupz8gDxLvMegdMD+sJ3N+K1m9zrPLq2Um2LDGglL
pUYVjCgeOljmYygX7CN/Dl6mF14IVX87SXngkvM0mM7YUkjvmWV6GXSiPhJE
r2VpdeqHS4aOMEYcKSWNtjKnqBgq4s7CBhBqLqwz90gLVMpq4C4qMTVC3Gcu
MqtleO+TdppCcdIDaKJ0NWDvP51nsfp0tqiZxcOvKx7pL0TNQkrs24apu5qc
Mr865EXBMRBUdqHL1jZDjXFYk3hyoAy3cb+cGhmGKEyNivXZ/dgJU/uIq+ke
TeiMeEs7q+qFmAtnSCaTmbuF34FI9TUVfFGvPEAJ9Ocqdk6DcjCwMQvfWsys
iEO2kl2zZon1ZkDfF4zrmzNL0aUDLxsT1DFid/Yr5AXN8j9pVafFjmAVgejY
JfSr3fyHtdEgHpyw99a8bUe4oNF9rx0ciVosh1Gg1FzPJ4Hbo28j0HmHbCVT
/b5h/+PT7/RPRD4Cpd+JXlLHjj4d+uW0L0nqncFHCxYZpaIOOzhhoV6TQHWV
89K/EulOBRemBucju8wGkqlIAuww6l/lM+jKi85zSfl9EvO+Kbebqo8NXMkP
50XjD/KlaHzypIjan4DWF7XVOg+4fFOdFi91SlNvrZ367O9vKoYOIrr8DmAb
HK+9KEYJFDeHC1PU1iSmHTDk8L/P9tBIqAextOj+JklWVM9W2/irXuXvM8Hy
NMx1HJNXVMmPy1AAsu6Dad8AH3h8GHnlg9PdwVO00ZWXlWeDZx/msVdbiPxF
1s+hBKC5UQ39S2rkptMhKKjBKmQBB9+ZkYvp1GEGXYjk5vSlM07bD9KkUfDJ
Xe/6+evQdHM1iMLHmzh2PNUjW6t/ZHQrtgjxe+/JtEkk9STpnIkh1y2zFC/Z
yaWBoUKTtX45bFGCc955DbDIrQuInprGZp4m0P1tiWg17sG7Y9p2uS3uGJzQ
FIBELPnhrwCT9f7tz6V3XNrYSo9Ob4SVjlFTAqWYVDxbDkAeSanI+7si5oQj
pLbc9KSt/5f/zEn2WlnVke0shm1DTASuX8b8TZkrYW3CmTWBPZ3q8rJLNa9O
4+wHdoGpceNlBdpUeWavdxE8PwmidhkmA4is/3OhQlKrU3RRC4SgyVLTDH9f
Jj/r+UOfp11pmcHq+NL5zvB0v3ftNCrVXOQcMRPkaPc6Wy9yi53YBwccmqZk
vVdU+98ebMb2afXxvHkijzo61PPDhUeki6XLzfjNUGsYmCYTm8wBzwbLXBsQ
MFeqFj8/JkdAsN7hn03XkmhzvUavatQjW2Q312al5GCga+z4e6bld1KsuqB8
n4BMy2QrMQP7uLjPI6bBdq98z0ylrS5cWVj+7ay12dqFxQVgxO7yD3DvR4ED
pbMfiPdx6LgUW85YLDpq4zAUPLdadQJl0mJkqnKtVqcapLtTI86LNfoAGLV6
uGaSeeT91QHxrdQTd9Q8HrZTCUL5+33BjAxz05hrbnQ2cb9CBCCF4cFSPArF
MYmu9mCZtDXQ7mWkhK0qX3aPBmvrSzVmYcXuWqqVQH54PSwULcsp1C9aL7q8
AOmn/3s0IPxZHwFaRz474yo81u9E401/ZMfaKSadLdy4vDhvImrNLAqsjCwh
OtXtM6IRo81fIFZeuGUgAm/ASl9B+Xr/rY5Q2hOzwWGR1Q90UtCmCj9dUoul
4aFxkt03CCa3tpxIJiZ6qb2y/3ak3xKUP4UtJAVqUkwGMEv4tICw0xteTKP8
EqUcuDfIcFvslq9bdBU1FVi0ZlfZF7uywQwJejEVbQoBAi/gONUmiHEMkpto
kNwZkvyZiOKH7qJOiz5A5DnOWsCIk3NWjf+gSDp4gdFvufORTCXQJImslJMV
99R8hwnnCdFTiujm6NETtWC32nu5+dT77a80olV8ST8eRWsyJbNZDm4l0kRy
ozNwi+Y5vK1Jh3kcBJ44RzH4qnuw81CrtQqoILhz21mN5Y64SOzAeb8NvJtL
VtNL+6Lgalmq4fdKwLFsTpnogCLwz8AZkqx4b7QjU+rlWIZ26Ssn0XTS8Cjz
AWqeflgJZrABXFvk4sNH94+yn3EUwAG8bvSRFa+sQuJk/ASaxS2RoKacG4co
jM5U6iqzz4Kim1ogCIlwjHLt59vT38pEf44KNKrilgguZq9bOQi3GJzmGPtA
TTi8eF36jdGEnx4FH2kF2tkDwIiF1znc5nhncQSGmTpXOAb6rGDKEZCmBhFs
ffW8fDDvljeTvfo/PcOFI+pEoSPoMU24JuRwgVzbMM5GQ8UYh3YDm6780n7T
jm3zY1Zuvp/pDlbbv04Ym8Ws8C827rM4t8quUxU3bRdVswN2qpvnr0LGT19f
zsa4orhR+NyAZqRjB68MC6zO2MA2Zk3oFPc4Ndv8Pd88xeXft8Dz7gGMjN+l
FBN5J4RkBakRrYmboXE16OOFoUdN0PYJ6hcBz5bANoPl5mh+Rdi3430ERW2x
O7uU7COFkfkTpxhaq2UqHyPCx1/jGyfTFqGNZltfMKj3OC1oU1/ZPGDaGdR2
WXtUvvUY85bwgxvwNAHnAOQrrg7kFphQcfE0xomx30Qlh8mg/QYyj8wjZFZo
aQtvWFL06JVWerxjgHcTUxJoNW3A01bvfHWtDmrve0nbP/p2xd2fGZl8slPy
5K9FuUkjuIcnNRkZWhV+DlZhGxdI/hc7hWX4F/sXin3Icu1TzUL+Uqt1XWa3
N9YiP+BnEu0PM7d0hl5TvikVKWReFuKb3488QqvdQNFaASTpvSmOhUq+tbwG
mDcaC1J4r6v65YC3hrtMXxVozIwP0zetIZ4Ew17gdD5SZZBkuKVy4T0YdXlA
DGEUlVparsO/RzAq9vXy5B35wvhhQ7HGHpcZjGvxj2bUs9kOiV3lPr3pNU8j
lzYjzQSgTbVIJbwFfTjA9LchWPQGLCRDjUNOptaZ0qewhWYjeGhfGCuTa5/i
d/mlNJ1U1ao2x3KUfullOFkz+ZGoK/f9C2kht+6WD/KhvXAvNiqfMCPtZGJG
M+NLc5iE8UsZ3B21ugsvjhMKGenalchYjvpFVlR9TE8eJsqWi8wiQ/JLpCpg
yA06yT6NVwJgTeZTWo5igK9tVPZ/r2SWyJc8WKG+e8ov0V/xIPGGOh8kBU8o
C/XIgJOXTh6ya6dcpXr5Fv30S3zIIv3jnaGTZppPHO5InypiqlfXjDRnhTfD
XC86zeaoBFvRHMy7GRnziQ1MMvu3BRS6iiTybFrnNOlhlaxSqxaO1WuhsVgP
UdcAw9iU8bnb9iF0dJMJZKUeti12QiTNqOd1YbYX0u7V4m4poy5tZqJUmwR+
yP0UAMT0lNgvEmh5pZngXOhHme384q+n7dSetY3Xbksssi+18shOKnyPnlim
J760zmih+ICguzqtPzDVceXN0U2rKg6jR+3tdEJZgq8m/EVkE7OU8yVJUGZ7
CORH0ptGcR+DEDeZjqegG6+COgiaFYqxg5W3VBxDBiJzywXLAYbMDOdQCcdT
awq9c+0doFDxQ7TGP7v9SckCf8RMn7d2O9+hdIO+Ypua4E2tKif58wj+q0/e
oTgUI56n59fnKKro29mDGb4dww5ZUnnR6VLMDDgAe1ma794EYOxuL1peZvWN
UcjuqmkFmhOberQbOx0j/YoheARrbCoKzEeWiOvrYpZdv7jt163kJJyrB91+
NQSHXmM4IBxRhBkmsI7QSWndW1eYwxEpuSblGpc67H1VImlIFkoBFd3vNMe9
xKLlqLRoAK4i/cqk6ggX+8riUbF/MDNq2v9xZ+3nP6AB5Q3+7BKTE1GW1L7+
DIELHLRyJV7YZUNu2xQLoui04pMlcRTB5PxSpHJuD/IjNsOG2j90si77gfBr
9QJsRT/VWKtFn01m4N5oyE7uFyULQjdLu4I56Dwi/1MymeMoQzOi/tnX+xqw
HgxibF+rBgkh61QFcp/QdowOQqNHw+iswqLBJ9Y5bmUCJ9Qtqs8Ksa5iKOii
fY07BptkYKDRSKr778W6q8S+/pBa64AyM+vRTobjeNeLYVL1mPzdCFGFkqSg
zmfsXgU6rgoZciWQZMujMkAe6+mOe3944L2W8dCIGXGtxoEHHu0jD1/pwhUK
IIrXDQpU7HGnoT+gSN3QGTz+TDjT3C6YTYCKAQEaPaJ3zlwpSv6Btc84Y3lZ
s+4o3WFjiU3jYBkdkmM3HLhTAx+H9trxw1ffSnNLY2PWKfttrGnPhu7GsjHe
cIoSZSw8ebX4y6WhAERvAQnHejzCM8KgD+EG8mNMOmpJBVQNEQa2tKyC98HE
bDWWg4I8xWjUZ2Bn9PaFzJQiS6Z80wOBUfNVy+DVUIkMpKNLJk0eDOkIuHMk
4EWQDIzPKhcqOfv3ne16z01+WvTXDR3KBxd8DcLTE2rS0IoP1DrtFoAJgdy3
vOafFOf4KV+0cPmlIa21CL5CfiqyZ3dxFv8HMQjsPaXVZ6rVgh1wJrmjQQrA
fu9GCiNB1dodUFa+uFA6rdz7dYLx0bih4JmpM00Er4RpYyp1yv6+4fJpkqSn
q/6LG+4JRj/MdvwwjYCA0/QeJB4YztsidwONf/SBlayRxJdnp0ha9zFK0CSi
uOWfaE4pltei2nWWFSov1/CZKYv3tplw09v0kVRI/sXhRP7xA/jBWmxkuz9U
8+2zd8OdW0IZAtDG6swB00tVDAw5H9RTUeJfH+lTmZ93hJOhGGsCo7e1iI/P
TPfoewz1eBk18CawCFiNtiK+Ndw51kBBtJ08CoZeBsOe61VriT3nWGX7eZFD
XtYNu73F8MxA/M5PNaJaCk8VGKlkNrlD9J59OtVARQH89eDgSY1BNH7HMq4z
6y+GQMzwTGHyhIKIFe9diD0qiTLTgX+FyyTZ+Mc1PDgndPlDyRIsW9hd0zQQ
dRkbT6ZEtVak07wjfI02lVpxC24/qw753GinBFJsndEoBlpJeTICiZH1Nhnf
m5IXxs+S+i2KV6F1rng/KuisWA5CEsiCdy61yoPLNLNry/32Ybb8bUfJZzmI
18sT+w0U4JNh1BRaad5EvtbFEtmyx57uVWMP4+K8yuHS6pcHI7PcEUJv2+kB
hliuzBJjpqiZktgwr7IW0WDpu14ToF1uWpk/5At7PArC5XnqoQJ6euZXwpRR
ofTubJdQvro+vC/HE/WML/xGm5Z/EM2SKN9lEUCtSCmr139RBw3NrHm3oYyj
qYTL/VKcBgkAFzasNodV1mXB3qGsmxfDMedBTtDOr6+DpKpAFIl30X0ybBTu
YG+GEIhKCMSa22GA85Lg6/SCIl3JKvj5J9P5N2zvSl2/pS8QTkYKaDmOeOF1
ZiGaYTvp6ytZkXCE4w7jz4TgheZKgu2G3sIOwm0F028WSuKiFmWibhDuF85M
WhIkaX8OY4XewujEV3bXegG1VCR4mFqPYlZEmrGNHddxu9JiW/1+/whNNK2t
czgAsditsYyP22B5I2wJPTv4eplJ9sX1ZXzj3Ar70KZSR0YjxMzba8oPaSnP
2/JtGdZF9yRH4iLNwzt0Rz9LlSfVqznBht4oAFA4HpYRB/sOtKiUm6wUwmok
mfJyDd57g2/Wj+LeY7ERciUJtSQ/Z0YuuVYW1uVmTNKEKwCs1GSGUIKEyZId
B5SJ1uHrFq62HwQqIMQ4fYrfZAzHn0c+YsKG6mZmw+f69OJrG60r2c9aXNLw
c1WuBDu3iqwkY3XgpvyYo/0tpVEPlGnDybZ+StF6zIkNdu1JMi6tuhfr9rFM
vOm9rZhvGcfApQFAV243Wa9I2fMTeXGl2bcOk81qp+sLmr6ZS2BNOYft4Ev4
29NZ2ol7PjAcDa2VMAC2qyjXojPHIGc95JcqbTmjoeSGQ9XLAd7gQTUa/Q98
BCdU3fR4BJ0ZA+yy9x20KQQibu6ZFLpXMuaD/3ocRfbJv7PoXS6iaAAtws+b
X6P9BHjAeaOnRIsnEFBSlM+VW56R6JkjnP7vhNgiGr5HJd1yMvmMJjNA6h2V
2i7VCqg5nYoRQV3vaRj3+ZorXFW4SmZI/wP6x0O2VTqqD/qNHUdATLCAH9Qp
jWZYTjKr8QGA34B8jScUsg+cfsgeMPGeowy931xWWp9la0E+adwOGPtys0kv
uz+ZibSe6KRonJ2WLdL4SH+YgjPMTYtT437wb+CGMBX6f/YTokXZYWgQBE9y
nNRorhZU3G7uwRlmPCG/Ge9TkQFoZNhL8yJHyInnCIpH+c95nO9UOqhl6h8N
SDfbd7ISknPhwagqjEx4cjrXl0OK95PUHIeupQZp9tDdMHL1+X1nUvvReY5W
U6DqNc45OvsBQEpNVN1orHqE8huWxR0wHxF26lvCZlECCIS2BwPdLe9k2uaj
Gk1zi+DOtOHlYHag2lh4Ijod/Q4nI65FosQNTT7s4bYJVsBi3bWb/AQHrN32
3TC4vt+oNYQJvR9AkFOw4slE/IVJGsu/gS9MSIuHvMBh7E8kxR9rrHD+EVHk
Hm+2t7aBiQj6OwtBaCGxa8vywpWnjsPdghfGzfQ2iAn3cH6MH+D6hwzyLHb4
T9x7rDl0XzzUg4lYPp6easrQA/Qqp+FGjZ6KRyRsR/2RSytLxa5bfNcsTvon
J+1FlA9wAfa96fd2Kk4tzFnhi9kftvteOU1OKecE0UEzWafgog5TDnndI31+
W0QK6SFBfc+CZCWus2dwHgKH6533IfpoX9qdEOKZFTDuEpHrLd93aAbtz7Po
EurPBbdvkzY38OMLQW64CSOn4K9wPsJokbqgF8PoO2A6jVUjOboZ4wsX2Vdb
AoRO2BJBiIetscfEh4jOWiXJqJ4zylkkxNcEq7iR+3T5zt3oGsywq1XnwrVX
cAAgJoGFYMFJnxIyckQvvvhWnEQCdua974d5808TZEAM0AzB2KGtj9scS6mP
uTop0AwLa+Z5XDHWy+tB3Q9+lhSBZGa3nXv/VuUOuJt/LCbvUNJ5sqvzOiIs
7p5JPm40y/JY4YxsIVSxUNZkTFLeBYUmHAQ46NuPcqCZP6BscwUzW75voXVx
wq1sEKOOQvaxXkhhuh3HpxOb2hYpxeSPBu3HAItk6qbtOmqSCUu5RKBoRnJB
/ty0VntdHfS8lhuxwlOgAXYKXjnD02ia2X/WuUYYS9H2ZJbLMkNtVJKNjlru
tu/4sfIFLvmYp9/eNSSWH7Ya7tEVrvw5zDQ4uuMGNC8NcWuVVCA0EC0d6jFz
DsQdD4njk0h5R2Qxkr+6I5idZWQ3n0VxguVUNDeIVCXfULHM78W4N0pyMkuP
qP2Iz50wPcDqEVCruQ1bzmEjjwnmdIViuR7LYThhDdJFOsF+B3jqqeruVEpp
zzO9kB59rCyKb6S+MKm4d24A/NyvhTxQsB1+KDU/722MKGkiLGVo03bI327x
n16bEqYeq6KUKOXkrFeXGiDu8MJ8QDX9mvIcpDTKXwQaSQxpvlSfqxMhv4/+
aPgqDP4jAyKmkM8lvYYBo3ldj/LszJ8hcbrElsmgTEvhUs6Irs/F3Fu8ONxY
ux7a0arHgPdr2KnJ5RS0duEPnhOpWaPtImme3h96ji+BAoJwlSRh2J3zfx3G
EcEvIfqOqmurarRIElVyHgRzq5rI+j9keX+f3Iw+FssNE+c8RJQaJghavOPd
aCTyY8H4/0iWF4OnuHKthJ0ywmQLOiMFMsQrxjnVC97uzC5FiHzFPECySTEz
IjZTPt/YwX7meW16UF7S3/aho79mk0oRrXOWFZ9OuN211R1wp8qzRkbSeB2w
PGiP8SZP+rUA9HDqJLiwKuzvtY9LI7cTA/2truV0zZ6Qxsgz8SAURt2qdAYv
9Zkuaz75VyQ33bdm0qpccFlRFHt1bztLosj9oxUgPsMfy+gOn7kvD5l+hoia
GMJAUTqG80qJq1LzoOsjTl/YDUjmZXWUQbZjjhAq1PTebwZf1T1oNha33ELq
Jik61URozrs2kG+P9+xLBxBaKfOjkk+W3y1aUp75PR/lABy9l1b3EiUwvkgC
M5Q6Sn7Z3ot34iPCzALCHaw4v+k7jFU/eaNUyS9v5aJabDC2e98/U+RttnxI
LGKaRJipBOr9kRyljV9BNBWX/vvcsVc4eodOyIfk3LnI4y5bXBDomgyUiEzk
RVxeQcBbvQAPOCt3DrwtB+cDTLY3/jgeEefG5a8gqJvPkpcoagjEn7Ds7Crv
o3KqCdxfWjXLh/GcEv4zHOMZSE107nWRgWRRclEtOVfivbXpmgCfPpKmhqha
Hvzt5a150OM9J3Bia1WXL/c3eWCACICRFarn0bEgZbv5e0BXOhvn6BgsbtoG
lAN4PpeVq40wERHQrgme7S+ZZbc4teRfeHzPRmzf1/bASD/+PKxG2KvJz0Kj
YuCDXfQ+8bCseeFAsXN6ol3fqT6Oe4Hu6FCLalgAHY2Mo3fd+Cy4MJoyPJb2
AWUzQLBlpa4Ao4WYVhlBozPtn0eytlg7p3zkhwXY3eMi/b/8+8h7FKw7ZRs1
4TBA2VDljtqljEdCd3alWSzmbW9EnRgr7cFrLRJzRHjBm6YPsHCujIQA0Nj2
vw22K97/HvH07HF6xm0y+SKCivJpH2uNgp2k02HXXF8pIlQeb97v9MZm2DTd
sW601zSq5jrGE48megA8QrPjDMLQYKvtFxLrWy0qnczCXJSki17DfV+/59Ey
2/5nJALEA0iXGB8AVHfiCUQLMYDZMha399Ka01rfTyuKC8xhPCEDPHC7AE3i
b5T2wxU5PZrbgZaac/RqFg5G4JrU2RYom5qpchjcXyCvaq6ewy2I7VrPWZPm
NAPfJLpiuxYdr4KKVOR6JFCB1DqgWVfK4QzFv94rrzkw/s+JCQNZ93JeHBb7
5sUFCZaDZH37FeQlD7F6ftx0yNXbLYpq/FETfvxoVwNQrMXHKiw9c3uuYUd7
CGE7LK2Wcd8wgtz8lF0vLEnnU+4cEqnQEpxqg+5fZ4dmkUsSqxLEhYqP4kPd
CQtdUrxW4wMIXvymRXzrUbrx0hNkQ5ASrxadrhtJsi2tB5mGaN6FW6Zq72PY
LC9hPa25pXB5fAA4tgmW+xIKOsgU8zspAlLWl50fOFFk24k9293QafULAy6I
5x8L0YcIQwwBNTyakuyWslTrUxeeYVg7UyKauvZyVnReM0fHmvtIUaYLMsh8
tU8/PvPSWJVHl0QFXg7GeRx2FvowrZM7sebUHI0k6m+CRDu5CGfprTURX5jg
O93VL7aqNe5oFpdtY+fiot6ig/2VTq4wYlVqEiuVtj+v3RO+zrX9rTLl6v/I
44zf+j/hulUJqfvjmEtk1RLE/AiPWzlZUSq7B+m4nwM60JsTp8sl8N7YdtNd
biGQ2kse4aFtIVCBbC7STL9m37Xu3AY/SJCRQaP/SaPsH40UwfLmtH2cgakc
niAWfDgkEvpCV9yd4JAyzWX5aNazxdGrrZIPnJOsPr1PyITwvb4zC0fwOOch
r8vSw6AQzPrX7xM6/pV5HLXFsarZ8pzhLnrmDRcyDSWJaP6lNgC7SpdvYIFe
M3P3xOPFu2LbUhSd9ZMnUqO/hs5fGNEEcH/34W8EbO2Vqhf38GX37Wb3FBcj
oPsOxAYmjqihGWPSRcx4dETzVYJTh05vHgh6aRT0P2oxCcVz28eHjprJ03Kz
0j2o4KV7c9n2pM+CRceZQJoHJr7VaDTF7vHqNtSZRInGwC+3Q3nmsUV0Wv/m
JqMVG73v2oLlDH9LjNU+81CT4WVZIWxXWF12zEdvLWU0sEoK2iHEQgSOkgcz
vvLJhrwgSL4RyytFRpEsTYFXbfl7zCAM79le+qI2RlSKG2iD3Ufb1/ciKol0
cUefblP2fP121GCHPig8CNqUWdbaCLGqFWHXmRB5ST++8dGEUjDqe2mt1lVt
2Kjxo1RRBf3c+DJfeXkrYyVFHKwwTE6rezDUo/xHpBIhgOKl0ikqcLvFawNi
hhmOT+TnAd2iA2EkBMcUU9pgC/+NZsx7dW3oPac5RP8tY0ceYOGP7VThSNE7
Ebu2eRPILgULkSL3XeZ5vaoUAvKGGEITb61xssIx6cVKe7KDgZVqDGZI2erQ
i6peXyzbblGRrjOykj9RWWRTemPD7EXpLM3+fNcLAfxd1EiR5x0J94mvbZUc
CC7F8LN1cP4X7kXagAMkYJWWxdCQk38GZg+FE+iqdIz4Jl8zOO1HBsY0YLkd
higyoATBZsISKRt2DehM01/0Hw7aFoZJMGdbqS+yjFoJOL5Twd7H0gWEK3UE
jER3gCsyuR6G0Adoywtgpi27DQRgt0Gck0VKXzOoEHeVRvEtb88QKLrMoKdJ
zngbgm49b1EOZRBJyTMIiHIIqURTzYjrEAlDf8Z+lQ3K9zU4k7ZGQnVBkI+J
ytJagwlgGy/vDE8cHdLeschqJmCmQSdHzAKn/22SlwK8Cg0OKLKKkMogVz/P
MchV/jFZdJrIRS20FThtPKHKuSDEX9waRxqC1HN4Y5N2pat9na8FCrzpEMUH
onuq/vZZVpb61XOodmNsRNcLzSWS4CM2phSKbFE/fGajr7WbqdNWHeh3NmfK
ulU519LApfkqHrmAZQTOELXQ8BTA0JXCv31gaG86wd4ng8bD5CwQNc9eM/q9
bhGOc4U9scq1EVvdMMgHB7sGDdS1TUzs1yGB7FW6rzRHfuMEnb7Ty0XSS57h
WORBjwb3fjnPrVQlXudMh1woyoeGFsqDR7UHsdphW6m3EBNurTKRo0izGNSt
/TOwkUXnpDtVM8d0nDQnHyOLbms2FZb/PrWiag3+RbQttr3QNFH6/uEhNMRj
P00dRQM+aM9jLHB+15LUR9y4O1qR4/AuJAv8ajzB+vYpxW8UJ8oatXjJ8GHB
+74al+PjFf5q/DQ9axvbyj4ARyedGV1OO/vmhGIZtO91wGWEaPHY1qb9QgU1
N+Cfz0ctMpPhyMnewByi+ehyBatBXwy2/AOt+MSdxpS/eacCFHRI6kX30yl/
fm+4+J5F1jEmed6luKjsBTl1pT9Z3UfS63BGdB0qm1meWx8vudr2Uygpq5GS
Q7jd5roIi3Thy+4SbuSpusJQ2QstIr23xKHoVT4Nv763E0UFt7uyMFXM1Qbk
XU8tDuGeAsRb/mE+7iWDcIuIcoDEfGOYi4Tj0o9QSHoN7MOEi3evPJMJZp+5
S/Wu8yNDrL6MV/YQbh31Q6Z6Iaq4bGbv6V1qBwaU7M07T4KeMzhvz18Xlbdu
eLQWLdi5jXnwOq354IlrDQICXuEnynlELZY+HMyKUON7l8igUM5mNG5fxE2K
ypUS4aN+f4K8+S1OvZSbwzVcqHlf8d8MNmt5kR/L9sVAvvtkiy7wk5Npoc0+
B/vIk2GWc579R/KndyRNV1pKhbDX37PdAagLAL8nH3UDem7wzCRW2tXufwBF
phETxSe6YtcEoo/Ic3Hs5q5uPVRx3+WaeWl8/XbsLR7iaofFMpji9PoSfIIO
Bm0vqStEb75gwjzP4W9/orSCakxnnVvHrkrZ7YXi947PCNNNK1sm/udAVU1T
p6dZOgW+7QCwFXwvG4VlkD+BTUq2RvFcNqfPuqRFN9zM0Vvdp3WUH0N3r9A4
nqZ9HnhlbytPXxfWAlvFZgI0aT86UZQf0L3y6n1IN7nfvu1ptV57J+scZExO
bHWhTq9p0uSIFf4apO4UDfHXAkCm6Mp1rnuNS0qaNh921gKca1ozJz/B7jYU
dcR5rQX6P/yFeLSN1v2MbdflNAJG1UjcBAxm6h5KAmvll63eHFddNfWPOnWI
rhVNH/89pi4uwOePh/wZVRqleF+ITqrblxFpIHUpxyxOLcEjfDWMA8spYW4u
ZtotFmZYUDdE0Z0pUVamwbcFXT8kg53ZhQR2yGl/F7PTZ2nZPVZSKjNdl758
FADd7ghPZzy7O4aTvWOhFsU0BpMASTLdoEP83bSPnai/eIP68SXVbf9q7EqH
qyfNdf1yvgRpXL3Qme7noMG5ocA9aAc1GY3TMf22Y1KWAyueysoAM2jh5CHP
MHlQMq2q9t8NRnG7LQy8PJrlvSL+suRqtisxjLlVMd+jYgZClpOJF9j1txgD
c+DeH2mhHcRAzWeGdZTPreMcHFwr+UKi8+2ralDAR+5lNdAgkOafdMJQgBnV
XMLbCyYien6Yq4/wQ/cHqfnw6TlMeF6sq4NsyMWBHGW1jvO6f6eNHk0OIiY3
jLBWtg65+EOECLY0IeOvMd1qwAn2EHOV8g2D+lIOrHHe6rXwRnXENmMDP7/D
Q9Om4/pZCD5fOuY61iG1DfMeX3LjPnvRz+rgjxBRNFSlVdIXCc5KS4N3QsBi
zE/ULCrN1xVMHFyxmcsLSFJNacTzF+4XJtxQK1snAlVGYjlbPbCXC2pBOVFg
l1vFgvGrDcHsgxGfGoXSMAtPHaalfsN6PZOUidZ1VpmWUPyNHf7EpR5iRG3f
+fdl8Ps9c2hdWwpjmolTkvsB5bH3B8veWzVt7uoPLx5DS2VVQqVHPoUDxg6K
RxSlmXcbJPHnN57gjMpsSwiydu0J8rhtc9Vgt+YD3VRzuRXpacP2AtUrdOVM
ThMWdkWJroTyNh0RFD2A0I79ZuKI5dNudskhGdqT4Si7LYn+0loP57YkOZey
bJfHsF4xi9peIT58grya/U0TqjowqtfvpDeG/KQ4QkEYRJh3J931uZsnV2iG
WlHtUc/2kW28p3msqUM8Qmf7TlNP4ypkX50KNCilYY3mAV8F8kF377YhG8Ks
aHltTL0Wd9b2JsTC3lQ+mV03tsfUefqyLJVnUDvn8+yV5T2bGcGIs5kwGd8E
M8T6NIyoGMryIE31iI5Mhpm3CsDXHiRSLSfoWhVNZvhboEmSmBvldlGq0FJ6
oS6w0FgV90tY9srIs1okQDQjPKtOGTPRmS4pjBlxVjNsGGUpSWokKGws648a
VvlmgN4F8RHFVNi79/SbQL+T9jZy+cz3+ETsjvImCJQllLgV1WUipwB9k4IU
ErmhrrEvym24TiSSgK3i5D9mQD7rUHB4tHbtVUdlWlej657Qa2lwAehUyyo3
2ymGOjXe/49SSH+nnLLOyM1d99+ovYIYZezfwN0RPA8LzIskSJ+VE5vkmgN+
is5KOoHYvwXGCJ7plHbLI2dMK0fkoOG0FaGAkWPHL2aVVTpjHGpRaw8BGOzO
zMMHe1vN3A65iJhOZCFG0nfa1YwDKhEwLQCsPk1IycjiBkad8XYULH/sahrI
pIOv5fULlIvsyq0cMqpuJ/fOr+OLYRSZ5PzilH830geRCpPWH54FQOWhwqzd
45TCm5C4FTXPhsAhha4tDbezQN2b6bzHYHZ8fVH8jCDzXL05QoSrXoBz0O6K
HlG2fUJeNWDWH5jpDqmHtq8FLcL4yksIXz826kN986Nm/0EfjEaRCz3xp93/
3jRGsJcr9E1yX0APQSFz2AGdnHKhPqnoz3acp/YuW9mEleRYR+8W84FSJbUO
d91lkvy9xjif/wv3UCegZAsBCwF2vQiOS4NrruxgLvdjtfwhtae/dnnK4s7v
sqrRuI7s7iJoU5z6T61Ct8IeYPMEpOgmLa+V5eMXZot4DeHb0bwWoP1w3t+/
KnIrsDyhLERJVY2NkPXfC0Ru62b6/v/bwNmwoIphJ8r5MaS73XmM4wHb49pb
q9hjhqmChgEf3uJek89tvHjtr8Fr3LU3i8RUz/pzQduhlDbFklqd6PLyGHMO
XYKqAvg7BjAhhJ55K2XNqB18dsjXLYiA0KGf8QBplnoFGIL8rhyY9vU4kdit
zomGX6OZaMC6QpMYQHljKrbo2/AH5YUUgxQ2P2OYvv3DsIsfs34TYIZZnp0E
2XsX+zF339GAAA47+MW0O9G31tpIht46QHa4Ozx/Nd2aRAVCJ2Brs05qR3Pc
+Tapa2aao8Wk8RkmbsieVHurrdUlVJr3nvbf34TPQxMVX2oqXdQrPhGgc41k
S+ypfa4Ptsw6x/1v5PMMFci+nsiN9HAdxOdzXO/nPe9S16MdTVuT/3LsIeM0
pqczbPAPCn/S14dhSCHDYkqqvVcjUS03idj5AJsST/f2CK3t4mMngJ4RkWdL
Lh4mB1Sgh5FCimJAu3CA+7taQeNoqhlLB1LX5FHFqTp1HU7uATxQRYVDSUwm
26aPM8tJZD3i3ALHj7UpXZhPtklfz1NJazlBpzNM0yOwi1XFD1bmSqh/lWfk
wGkiHffcGzYN/7pkUoymTOh4tZzUq+4Cm0gFsbcx75IalYINUYBEZwHj4ela
frJk2avm6S8ugGjXRxkEmbCPU/50zHTW2H2A+LfMESvaUK9nyUiAblJbsQfF
X8MDVm3LYf1s/quyGpVhmdDPTGLeFwaCon2wURQi6Ykq/9Qq7SfF/3mmCnNn
fpb3iLeBY1dON7hUTyargD5XGg0wAQqmcPWPbybmk1KHGdfNke9SxKw4gLq1
5BbWBPqfMX0JDWLsh/qDoViFY33fGJt3mANdLzXmmWS3kxAYYYCl6DtG0iCN
ncr1DcKi3Fyj0c+RJ8KZCu4x0XhVp//6DpnTUWGliBbiUAUD1LCecNFPM4ZW
BrPwwBRonErCT2s6f9xbzNuRv1HMfDabATjDo5VkLGS9i0Vwi5qmQS7GI4rD
IcHi7P9xtxO+94Igmk3ZAZvTkHyu9pvibabLr0juGfIKmd2vo6enKN++UC5a
8g4R3vbYSmB3jzR6a0ShYzzb52HjZixhU6scAmtVu4WVimF7AdF00Fe2b0do
2lZL6nXRu2qU3Gij+OkQKKuX7aOXWRYSY0jw+4S+PpEgofL7yPuebussYioM
mrFPwjwsFlwzix2DCijBK88b+27EL2YnxyZ9ID4IOegC3mlwiJsal2YVCixF
hyr5oofZC8iXls/EoYVsNEhffihg0hOkC2q7lcpBA1KycHweJXP9xjALPyK6
OZU+a5D6nVzLxW05zrgj3WfXR+12m5ZBMeMcazv7fC1gtZf4Bte8wyKgUEE9
sqolMV6xoMcOEEsHfP5dAYekHJStxBW4jBq/CSPC8r9QaQl0lfnzBo3Q2xxk
PTUS/Gm37mxfcaoWT5yCEFKfyDy0bpPKVzfh3IBUHRYka79pxtj2eONc91nx
d55nMNTKX4hR7EhnAhn1lmPpv+pROXpRlH1mnKf4riKSgPqWgkkjNzBpgZyH
jf6/C2SWGH4xgWsw/pVXpaxz4TFdqP+SzTPKm1nZYQm+QmtWBHQFdIFnOWXb
Ms83TCvIcXIDKp6E2gbSnR63PyzJ5zl32ZV4/JtwKbE1vLkwWhPawpxA8DKy
db25O8eXYLmfJXINQprA0mv1a5FWH2sgdGGh8MKpEDDaiPevd83vbYPJ0Vx9
46VIPYN6ylw02iqasK1FdR3lS0NpYSCvQV4ICNFJEalUvBrskc/lqGENJUm7
n9AynicOCKLXKUlp/vRGya2P+s5pyw2QB0vm6eO57NHJVUEGSalOW8/G3fwM
VCPBZCqqW4xmemIn3koQpgnyH/PNegghCaiH0vtEIiqpbYiSSC5acVPgAty8
WiCeWbFnItvJiC5br9G4h/CGmOK2cD/KSQFV+DMH/kDGkfx9e9GmpSnW1AEA
SdYbvRspwpeiyzJMt5xV+7qB82sNtNhAlM3+RfMEQlolBPNihGMPy91A7u+Q
DCy3T/FW6DTmKIPExVtdXBUwOhHZQJlqiE8+wsJYM/1c/hjvHDioq81LaHlv
sXxjpfkZknoRVIqS+gQB5mlVSwV4e1jVmVQIpjGMS0SKTB9MGCquLzj43vBN
iXUHiEzo6AbLBJJYjMNB/7WwZJraEgFh/+vgkvlFDLUKeuKYbuOVc9484w2I
Q7FCw31hHGJPf8PBLotiMG6wSCHIMhx646QMkPzQCq0oCEGKqGxlCSQDwe+b
9WwlKCDxNeA7duzfeBAMV81ZSRw3yLIcD3oI45JduU/W0SEfHxS8Oow9D8wk
lZa75cLZtACaiKyuUePS8lzbS63OVn+qZNjOWoNaIn9CK9nud2r0RbIL5RV5
GduMdiEPUCMIf87PgmRk2cY8w5EbuFkYd/TPmsQRaQAcN17iQaixk0LTwAbt
BffT8y3fAuZPLlkaHUcGH4g4nrevNGU5kUEaOLlXet1KXwGuWnBH96/lPPNJ
YdEceukEAmFIf96GlfpvpXDqvNnPo2svRKXvqVRuaUXnEy10UlWVuLyR2f6h
Y9sTPfnSu1mE7piVgzB7BgXu0PJgBCGxU6vev0Si0hoTN6ibDi4DI08zICIV
A6Oiraf0YfqvPq0wlsP+G1YndLMdXlhLPIBZyJr0kQz83f8nUZ1XMsxgoA2e
3I9y49sabJvfnjV40XOG7uBAv4aaNNy7F7idSsowoLatoFmJ5cNMqtbaw0DS
2Q46WORW/0urU43/I3NI9MxUEgDAXyG2LJogdo+O1E9uQKIavlro4iDreIOK
/KvK17LwzzeUV0DuO5v+z7+ZtVzf4vJ2K2K5mkKRlHvJ3xhqN9oom5x6+p7h
jXIhfDk9EE0mzwJFzOOSX9eQ06+7CL2vfaqbXSfO3IpQ7SgcYIZwhlOjs22o
GzGepUFEv+keAOUuM0R9JZrnyXhXFQM9SbbGtAwQROY9ibAU9LRDvDCCrYaS
mLbS3lZrlb7SqXkZ8GOgTQ4FK0mHtce5Q3hMfLadWMWEtUV2Wc0/bhM6VJ6t
aTClUz5H04tne4c2gppu47EzSDhiGra8jvL0P4XStpRwAw79YJM+QA2Y2nqT
eh1+gashWDx6QBYsxVHROECCohWPSrk2djBPsqD3qfZB6+AIrJ+NqGuwcHBs
0Lz8EpIYHlP0tyvr08WG51YoXi79Vz7XVhUoRk1G+jo+ycjCw7oP0R0pRr1z
54cLbDhp0bsjcbTH/do2h88d45PsR4zZyOEjdoXp7QzbhNUSa+nkfVk2KFsn
USYQsepsKBagMrD5IXiAjepYyKsoqI0WLlVsfljvbx9A2wi01LNVQ63W8lqi
iRvHWjg6WaQTpZJp9stAGr2E6W78HMFe7z43ScVnuiJVh8HUQn24Gk8Xw6sY
PAi/4Or5gZGnYm4Dc/4RxWrhh5eKUTge+6jLCiAbomu8swgQcngTT4Zc0PLV
5qwumRQWKNFvqoNc2GWjEsQimauSQfI6ViDHUAwEk8VBGNtqH9xO1Vm4cWeQ
9/hDVrCVxwQoIDeW7jyCsMOtZPcKk7ghNRxAkx1nAh7cVd7Yb9Rr3OTD5t2M
2fv7/4uhP+MQUAIlF8Lw1ZuMkG9DIGU+UQMQIwcBZF3c+kawQkrm6AhD7vXC
sfY2iJkJradVVKPc/QlNeAeQuAanpMDWeq8DBO75PHX6WFogm92/9kUQC0Jw
9TIO2OfgxmUy1AquJGD7siT294XhyRQScbZZqaX+beQ27TPFVQCZMt++UnE9
Ew9ZCJYYXAZcvXnVutzdkgZb0qJWMPlNjYi1v+HZog/lpPPdcrueoAS5m8Qw
km7ideJrns76QCGVfTaK53dcmOT+2fxusonpa3zdKGmrkMD6lPk5iE33R59z
K+IgxsXnfy1zDqBgOu8PKkoQAtRvGROBo/I5af/w1KJdxX1E7gVqEFRdrDQU
a9u0d+lftnY44WfN1aeVPcOyM0n34bDy3OpRHBJq3pH7vrydqlFISxrSW5IA
rUcJaR5itHGs0fei3rSW3kPXDju1RqS3fawcGze7Jd4804AgMI760Z0ilUEq
nFJrhOZUPeQtTWS8EpDLIt/6IKguIOOTM3CIt2QYsOULfdORCpiSHcXgdn5W
yRgB6lq7f8sxpqqUPFnuuPUYf9C+KDbArBNDVpPUGTqevQ62bQhNEvGAZLFp
SV7xQPNTMMxFezIAMlk5BdkGEmBOSsj7KEUyuXkFvXDI3Bzzo6ctwUQ0E0Xf
efYkZKev4WFifD6mzVaQhGTdYAtuyQJZMdJd3Vn8CHpV79yqTfJWLcle1oUG
dVHvJaAqfopYG/KQToBkYJ6fWXc7vL4PA3IQurX0vgEAEpzXRCeaZU5PgeVj
oOSN5kLvVof5cAiOlyY/62uZsd1kboXo+ZHd1MhjBO58QHZBvsjk0k467mNq
50pbvu2yc4rGd4VtP9DCowuvWzU3Z0RVIZvT/+dv8Y6i4q6JgmEndBXFui3l
aCrhIy1+4JY7XV21ZjoS9eJJW6JPDGeWigb+40t5Y/Nvukc5oZE6sKRE+wYt
8/eOb9wgYlgqGqdmBXoWK8hC4oDqzNrAouCFj2kXrwr4yfVHJeR739cr1WHd
2LgWmBA7yjUiKZCYCgmJpeDQ9ux8wboUf+HhKh7EaL7G76sLcE+EKqYtM7hH
asa8PkPXvICA6QKf1tZpJl4BNAzivlzuyJmv9sjWiSS2/3+j1lUEfJ7MniMx
T6w7fnA0HUv5zfvyVHJIA8WJexbHXaUGhgqYtsqQupir60BZBy/D9y9J9qk8
8/3W1VNEu2v5LgewFwwiMP2If0inDZZ2pYS5i+T6GlDEOUpC+6W08R+V6S7s
PvIwC7QzjBfFCi8mksa2STm5XCCSzXMhrnh0S5cHRnZfZIdq/20Nv+1zn21F
+MkRZvZL4jpbUN/Qpwi7iSqTsd0bNdcxRjH1sTLbO2XEhq9h+fc2vUAHF972
qaEUK/SZgXuhLeu/YXqtC6xEglNedP8Kk3lPH4leHr8ogBoGitPnuAmAxKGM
x7ymIO4kGhUly2XD4jtoTnxdt3uaKeIkYhpzYlb4SsJ8OZNYtae3flLqQ+Tp
88OsKYrr9q5hcc7JEiW4st53FDe0ohs1LESrSFaE/tAQXxpkwpXCij4ciBOm
Ljaa2du1kpUP0LmBtVNQpz47pooIJrvOzscK430rT1aTZFQ90hrIdi6Tkkcy
nUCFE3iwuvXhwUv+n94U32onqhNR5jMS99AuLLbt3e5Hn1AzOOiONr++RnPP
avhcm6iyA4FmDYskjIwBRWMAwVQSBLwI+ea/c0HMhg+w08y7ehfsadr50Uk2
qHMl3iMGpVOaPGgIWyGUcZD1QZnhWimQjwDZQqzO6Y3n3W4tsyIgfrhPyVIJ
Raj4AuKRROOroUbTBDwxICIzxVmt0HEfkTEaGsqwglA32MBPx0M7yMVVIde0
5kdiMPiX/w1ILuVsyprTNy2LzeoBPXDkLIBHL8KTp7VjTpbldMMfFaoJa6Cw
yn9AEueWrHef4b9HPsARjGQJHzNXFXhMNFqkyqOccq1RelYgk7BfvSgeJ1eM
6LYEMe6n4BqI2qAYsnL4ZWoypIjr4IOZlFsOncRg/803lAGuOuU0AlaT7/s8
KHmkRHrISMZLQz0bH/3dOH1YyHtS50XIxcorJJLZRsnJu1ea14NpGiRf65Se
vjDQAFtDZXPqb/DGcz11mv2utmAHWUBpX/sLiHD4s/76vBfyiyra6Udz5Vxv
QJLoX6AuofCoN+H/2NvNhzZu/PUj9MF8Qelcs8vDfsCxEXYdZthuQIOiGdNx
7pIhNrBu7T3I/Y8uwibFP7vxZVPB7UqiylaUOzlJQgZWgVq7LpAplwwvOuD1
y0UCRG8zRX5s0bAkracxmhYcGNPFq2uCQdTb5PBF9qduo50tHaVcSjSw31qX
YxVTIMx+nOIdzdtw6F35sxwbtEgdTlj4JsSHTkIR24Xw0/GjqbL9FM5eqldo
sXLjdXSVAe9zCc7BXEnhbDw3Jgh409U9LYf3Osyt8yDEc0Oo3r4r6dc0UVkY
/zO38YSSSF0sbhI5qE7UyxxADIQtOiYFic9OuvhOjL2T+5yIgQYwrQegYtt+
kn67eMOPV0vsYFIV0N2GvXvw+4Cdb6T2fkrgXAtbzTojFT6McyZbXkaLscHE
BI5KmRRaZcsOMkjaJRb9wiS1sOVZTW18LQ6hxp2cjXSF93ThRC6BlrJJGAnR
M5dUoE0X+EHS9AEh/ovW5A/dfIyNU2UozMCosgLTN3oHOGjzjIVYF2FR/o9+
EdKp680LlY1cRoy8sErB7MGfybtGv+2QJkGqWndGU32BiEXW6t6r2VNL+3fg
p3RYT54obj+aAA6mmnGrkim2UpZnTfF/d9I/udlIwuTbRM1ONLbzgQNEFmue
/z0Un4BWxmL8yXOSuAqwOG8gyd2sNqeUIwSt5QyHuy3bXX0bXETuR2SoZnZc
dtH7GKhuBGzpwwKpqTbAekvA0Xnq83mxNqB617Z/W/Ey7JwbSy1SEICZ9zYP
WBXxWIJofNFS9lB9x5dHJcMOA9KEkVySJ1A4tJFlxqvEeX6ZCS0UY01E/4gY
8bBGtuDPTBkdQVBnMzpKZMpawIiSWp62peyulzB39D8JmvyXXH8y+se1Ughj
c+B5b1YIIRX+JEhE61CHFExQPEtG0hFXsmQItv7sY7tjfAWlgf0TacFBrybk
Y5pd8IkEmaheLFDUEB3s5b9HBHEywEP99Gt6lPUFZYwTMCt9x4mbzkn/6CTy
MCGbS/vepgfttJcFJ62t6C45MNeZZC+5CkKfbJcOStjGKArCt8BhiNqoVM2n
wocQHIU2syoo4SwqrqwOF98dFOh8USrJpdre86f8vd3GLU9wrYKGCBbKwjuo
Ahty2HsZ7pTcrftXDyKAvV09SKmvihYCGSBKiF3tJsCayFyKsMj3D8Ml4O1h
3GO/NQOcC/QYBH2Fum/U5arCPkDJwUYkiRizf/tU1nMrriJpCDKyky0GMzNd
nQRF/BNL8nJIkddjro/5Vhe2wMOLWM4D5HTGdL5lu6sL/pmQbdXgWtLqPLsy
/r2ymGgRHteAKb8KQtESIQBrUpOwkF20tkBQG4XXHxAbESDYy3XOW/AuLzoE
vIMOi6/892xm2KgoFsilD3y/0M9L450YGH8pLWSYtbJb1EG+AmmNkxBb3h2g
tMDL70kVCCtROsD4svT7uWegrhSCm9OjLq9kTlm2PVGx7jor+Yv52Tr1dQR4
wP3bsVMlcacT8LI3/8WhJHt2j8OFewQ+R+BadCD6AZOU5NbZqd68Lb7OskF6
2IZ1bfCcwPEXcO/ZodHXmhxX5NA7Lih2NUKg0gLA2Xp1EEmlYs5LmTQH37Q/
eD94KWbReF7TOhXooAMfjOjm6NGnrLntIffstvPKLS9oKcMXVdxuSA5R83QM
DbKgIQQHgy593oB1P+j76rYdNYN/RG8kP3AR9iMF0USYchbnK4AfvJEQe8KG
+5OisLvMwKK30WW+1EyMYvq4gMm5L2y5hw/YOwZt1ysJWe/LvlE75kLzJCFF
dVYNi4zYftmNmfXaorI2mFpA1FhI9mh83O43ECAWBOniEPl5rEEM9jFFcONH
Ikq6/NNtm8/2W36wUe03kZXl9IuOZcKQT1JFQCuLuHeyQYs5pjv/vIpwNaXP
M3jiECmkOxlhf+XQEMGSW+AiRyL9o8jVCq/d1bIaiFBeJHREvrWUY3OJjBvU
Ot+ZkiGuBxh21Q7V2YdkRVNPGMp/wTG+8HbjupYeSh9a8icCfscfGQfRWk3F
ahR/Oa0aLDw8/LLgmtDKZ5arhSvhDqiQbucl4TjJyPGo2IgkPUGlT63LJjJ2
Fz9JU1hZiGG517T9gfJkgWDW1tyBpxRIeJhaaAVH6TS9ALlyUhzWC1L9C8wi
lhfEzMvderbqbSXtaTxJVADmReIsgKWhsavZypQaqjhLhyp1Dy9kBD6/HGT8
SYK1/MBVG91niSh9MIxtExVYHf9WQLGfKkX7sCTZHopGEusTVRQATTJN/ueM
C6AvNKteoQ41mJ1swudhxC1uy/xI69l7UTSuX1mB3m2SHnfXQaw74iWuLcOU
+s/5b1+QRGGn8jyB6NZs/GMgrvTV2hkMBQG3qso7sVNsSOwna9DTjQvpB8Ca
FunbnQ+aDujgQwBTVq0bW6EOWE9PN9d6fOd98M9z3TZgCwnR1jh5Y4PxCHxQ
QkqLBgnnqVQhSmeO8B3OoOu9+OW373eQPgHUbyAkntQIlxu9+c52EQQi0Rko
hwT4VX65c/f6VT4NphXKwZhwso4N+aIvl4hslwqOh3yUtRApjmn9K0hYiSzP
i6y0Z9Z52RO6BbSnsY3I7Qiygm9Gxmryc+LyyVwelKZETfknWsB/32w9T47F
akS/COgcy/3jBcnOP6VQfjc7n5tAWMDWnG58jnpFIyRFc9MpxrNGWgYN9uFZ
RCpe1v7M+uxE+sxllQUwsXO0/K7fbghx8LlDiAeHCxxX3/oJJYfrYNy2zpIn
g+miRfJPfdNvW/KBoiAqFKVunrfTSfwqF/CkDl+Xia0TP1neFzb1rZULvSdZ
BZFOh63zP944yLD8PgpWId1YtFbHi8FQ5qbx1kCkv75FxIixKblYyOBbtJWu
cOLJphh+SAFevnCLgmSzsS5WPng3AzIP3WcIMI1XQ4apnHBUPB2615WTqYsH
1bILDzOzj47k7DHjaga4SVkSJUO4EhXzTxxEWbE6MkMIyJwvckUWF+4fep5R
MMWttSF7ocMMBcNcD1y2zl5dMn9/pcKZzl8rLzHASYJC7XrDE7zfiZl9cKy0
e4zNNCQqUVFI5k+VRT51bdhM+4i3TStQXNn5aLzYj4mqDsUaHw/+onEuyZYv
SErcwIchFeGnAoFW1OUpnpJf91Tqn95b4G8uPoszbjYM+/SisNTMaMkOrYBn
1Meu9HHBHf+vqbj2mfnWpQhjbvcXATF2wxuMC28GKPnHKN62v0X/TTHqKnxR
G6piwo2zg23babey3eU8a2m8O+KpRhrTS2r0IUOTDhTX1MGsaW+OF25Kv6Vs
z1hqJes8Tn3eNUz6VUtxhgR+PLLKGID9/Dv41glsnVNSHAenGJOBf5+k0mVY
NDzQVlDhIz7+nNpw+EnlJ3sGD+pO2Y9kORjcF70KvzTzMaBC4bWpnSq8yjOO
SdspvFrrQGNnlNcl2NAqMKr57WbUZnzIbOO5LuUKvz92/rmOyQSf1J6SzyBW
qmHv8vZQ0VCkRhzd8eUC8V0You4iSMbp6JnxN1HDZVVUuGcO1kbZI41ewXYb
bh5Py+TEzE/ebgcJ8RptlfPt0Ci4t0zwNAgB6UyHTJO5Tbe9xxsBgRR7R4BN
VAiHmEndBXIW+d+1HCjyZq13933o0jWrwCGotr3sm/VPPWqEK6cUivqHqBKn
mW3kVl3ZsN+RGj8p/5awxH4KBl8PzmixIRFoMrVB8h8z///K/qsLFovDqQD+
9j8dcQe+dkd/mCE3ZZg/Aq6Io0DXHBQyO9I6Kvoq6KDY98T7IR/oVK41oHUN
eex3V+HAfuLVW0Qz+1HVLmY3RcOL2i6w4aNyPEUwd89CmmqBCX4fn4UHW4rR
3XuO3mI1SBAvHUl/eMHSWv9JRGxQB6giQCwoEsLhTxHprM36MjODcTLvlglX
NI7rNFuE+TF57+pJoVJWk+5DF7RNRzB0w9RbXS22cy+rr445QDu+pf6GAF0E
ejuC9GxLd0zrhAGsHHU2thB2kJTzFvFcip0s911ob/thZvf9BXOT+yRaS9rS
9zCI5bLe6NrqzY68r3S/5VgJmd1VTPZIwVlCd/4NBpkZBf/Bk64MYtwnoFHz
GAFRL0tRbMAl5C8qwGjd7RonCC0puMrrKQMdpbXYUPV8tz8nFvKDcEZ7HmtA
+ZsLoC2rOJSLwkY+SI1a9wg0uJn5IgrQJP6lewR2URwqhQ+c4DIJLQDinUFH
r5rn6NN8L2h13MDZgm29y+Zd+ZyZqws4q18SUYgVDvy4cK2XVuzyl/3ssDHt
V7OcKWG2RMMICA07SEN3b2zQqLKLEhbP3qN+25ShQsWeFClkcyYo7q3XoKuU
HvhA/Md0GTnO/+W+j3vQ+i7lgdl8gjjWwaCP2IKnE9qmdShK+saTp0vYEQ3u
XEZRDStbscSMOOteCqyufZxbdVJ5Gllhh0VPX7VMWQUf945bcnDKAVoKT9C/
AAztyYxoVAAO2DuJCgT11S8vpo1DEjACMBmdFEOKd0Izbb3ImDPlt2n6jzrg
i88hGxA2nI020QPW5riODcBMRhePK4ToWo5vGd7AP7orWg59/QmEPqMsukhw
mI5alsJPOcj/DwQzhuflHH9BrZWv4ZmL0UVfki53h0hUxsu444nA58mIqQIu
s8LKWyAsd9xUp/z0o97dPkKRGCxkS5BOe2jR3400TdGttQRV5MVePxhHfPix
BVVhayvYYnY4cZCWmtq0CsrvOnAFk17onGZPMz8P4m7uQoKZyFu1HwLGM3lq
guNHxfybOymkH9/cos2Xia1yckWkuhokmsNFhrYNKLm2YLnykOy++P3ZYy35
4uY2r1N3SgHoiQ4Sn1mrMSnMUYghlWFQnrFp9vDSeM7H3YypsFKnXhXUSBBo
i5Z+rALsUjU+8El303pHMU08JSWjES0Te2vyxY/yBvXS5Sxr1HBRI3VujvEA
oecU6bvJJ+jSuKVogHCrG/5JLdJPowK9eDig9iHHNMQwWnQH6lKlqgBEP+h/
7Z3aXfS5+zwFguRAXpkMyZQsyOGVyj6g78RRhZs79k+X3rO8YZKKCuctB7mT
wT8SbyxLPzKR9ZlE86VT8FNLtNrY8louYzauwHlarxO/AFFVwtQmmLIZcySw
opupDYGi0IUu/2AH5HhybowKI90kbhjOhnaaO5aA0Un5r5+D3jEdi+4dFLht
GPYHRc9xU38ryRd795obtowSUt/E9K8bip87yqA27Zk1Rf88OcvVdZ0zlfTB
3Gm9DLX6yRlhlM49fXe1AkxDl3Mqc6zUIuhZQmkiXPkIJfJaAm+cEH+Z9tUO
OB4vMiVa8qRZEdkmlcmm1mpE8tVq37gWOs9O3zsGi1PFw4FdsNQQq9JXk2Hh
xvKqQ3VIZgyapf6P4RsnnQpdnyD2AfQ2tbYyqy8GqNvbIHdgFUheJERYNQRE
JyI7vOE2NXi4dvYhBvAcZ4XGaZg6eK5/HIrW8hIc4V1WiLMEPUH2a4415Dlk
soyUm3qUcPex5xYs/lQw6YPu8sgYe+0kuu0thHr2OjY0e65cx0mRtmzCA7BV
xFjJdC1XfEiUjvhj61civlQS5Tvof3UqHxIc/aMePv4nTYpRSsBvCKY3aQFQ
mVdsXXLDG8jRoP3nkx2dpkFbiP1MzMI31KwtBF6qUgaWBU/8oppMjFOBhjN0
n0H84YWF7TdAD4sLm18R4EyjEI2uMdEFZbmUouMrfRuXLAnLQXvcEuHqAu0t
KI8CnUUJOzTkPtMc7JIgdxz3RJOq0fAwutUGjhPFnT8R2/kaYoVYBuR0w0l9
LQIqbA6UxZtb39VDKe4Uk+Dy3YHaV1PS6WGY39WlH7/b2yNMdnnFGYCfzeMN
UjTBHsrEo9tUJbXttpDSBFDejyDzxQVTSJELdQrwYIXF/w+s0cHErR+CcL7D
e1ef4Bpk8j99heIQOlbI5Sme+yPSIC9M+dNkdohLaPz5KMbKD0fWRAUUcgvE
5aomMkQ14PvaUTiG4NgQDIRMXA2iMeWx8gPbNtr43262HGXjkZXOIuy9kJGZ
qT/O1UG7v9P8CW3ww6qlXpbksfLERaNip1uWb4Ypj7lLhQGokpeZLNN96xRd
1w/rV2PnhF2/nO3o9wE+6v9D556hLHG3urCakS/0M65BORqdKR5TZ+ZqmrSN
gZ2yD0buLbqInAfcmjiR9ABkm0MjlweTpqz5NT1b0PgzBxjkp2EIHmy9U1iS
wo1V+iG69pM3iLg5AYPof16G8gkof4M1ciTkIVGq5hlgqy2ijwt4bFXLCz6A
+TYLKrsyTzp1mC8aHNRzd2Xib5fC0zXSAhWB2urE57eL6dIrlnu/83jVkPuR
dtg3qCKAtKrwXMWWymEKQ2J2JL9G5DNvX6VoJ2agh/PwR4Hp4itQAbmg0Hcc
xx1EPpOPM0rms7VRz1Odh2PqaoEZwR9n9F0ovVctvbBnvix4fxHhZzXKMY8F
IpCq7v65mj1DsntCDoR4zz5CFkDYzVQkNMdldX76p675VK7FXzZ8Eayok8/D
WlWEtgTF/TV4MonxHvl0jKQjhD2uTe3R9UxJnRx6bL/dVbJgUsVtGgIEmC/V
KfJIa2jWNDIS682qyb5KGSHu/UEYJ55dmAUQ6nqvmD1f63TGzPAPH1LH+SCI
W3ZTvoqS218CT1vzTLwvb38J0UI+YAn1JCXiEfW12dZs/CoO2DDeRPakEwz9
qw/grz0w1VWrYdFiA7mBsWkRI7Mwn6g88FAi9NSfSc4c+DKul6vgWUr0IZ7l
yZi14VmersJKS9XJsv3orTaGiLwh4rmKzWcqObY0Og8Wl7BZby0h8Ub4kD4Z
SZdZMCO0HAzce97nSEsBUdf8hMvMo/K5dx3b24nZ8yhBcL3siX3sPVPJXncy
9130x+Q1F4eOkl1kOZEDjeubgWG3JvyfFX0f3gDZpWsXVGN7QLpL5mson11m
ruaIKjKOUjjKJg7DDHtvf80+aUAPG/zVRHJzfBv/CGPw2riLcuJQcxfGZwjV
dQv/kGsnNH/UaH/LslhblHCO/E2rAgbIR4JdMyeFW2oz+xJ+mSBkbAgOQgDB
P+WCWqU6vxBIQfnEr9WefGlvNpYztyekwbf4wK69NVDWgldTncyq3cOKEcyJ
CScEDzD1LDfp6ydyb05FBpjx8wM/olDy7K02sEQ2S+Lr25vPB5W4tnV6AQ1e
w5manXBuB0JKfu1fEhXlUedw70mYgjzbxkvumKz3lR5J7BtxXyWVp3YyKF5r
w302gYiaLXZzu43201bE6D0BN/XbdisaW9tlyrwbEmymNjnNKN1uf/DDaV17
rzzyvus0SHvQGCkwkTxHoaLA5PVH3cJZHDCHgo5Z201JANF+obwCXSlUo525
ICYN9XZXcv1Gm4SKdhVJtbIh9ki1isXOWmdnLJeKibGiVQUGoAyofAVJMEJd
QnJoLGnwnwpsSEKCeOSWlLaTFr7L4CIXcII7jx2ZZGQRD4afd7lo7IlevQYA
roeYPjxpM3rylmxSySQWw1qE854FDhK6ezhwV+JxnKnhIORtTiqDE7fAdE0m
uwbP8BgeXPCvNpHtmGu/t+ANAuPeQLuVzldoOQjTlhyu3dzJW+7q6zVYpuJU
imgJGGn7xDtiTDCSBYS+nYaksj7LmV+2ksOtUwUxG92cRKhYc6Abo/Q93XJi
LA5a575M3Wukk5T0DXXyJHe7TA/ccvlmjyad2uKY8bZtWx78XIzl/1H+lqL5
AqfTqakF/ppER1Hm/rc17Vdhn0NYcgDjjfi2VyKlVQ44GMQFFMP3n0eJ+kJq
FThTGYwpif/PZU+xBF9vhlvGESA+/mhAPgzyZdCSqNR6WaPIhAuuwlPT0SGd
Yiy1TvfCa3W/xTfmfT2BpTsRMX9azFg83CuYFRyK9tOCs6wpobw0Jeku8DF/
+YpOQjVtaZNwWSPCCqj5CnT8BtiQ+8CenXZO/ASoABwlQcBf4CwcNTeeUKPN
yZtCm+g3Akpgwv+8q56toxVm79sBCG4V9HxWdQmlYdO4941IjLpAvGydFxVh
ams/at5/pvQTzlnsxlHp9CuITh29VLLS5CrKwpHGclvxRmANaNPRTR635Ec/
4AezX8r/0QiKFC1wqkzvKTUu3IQcnvydG2mB8KcK9wSXlN9+AuTs30hzVQFF
W2g1LS2xhM7CvjrgUelI1MA4Xs8L1sFY0MjI3sxrAydc4HIJ4WRgB1i7gSDa
FTIgcWu1jVrcbPUTU6sGbds2FpJLCH2d8W2TfcS8vMrFkfIrzhwEDpl4RNKW
zNl999rxjz3sxp+TLmnmIwiKRUvaWFJ+DxSJLRQuaUv4Ae6CleEVJT81ntB0
Lm9DjdbF3xbi7MGXzDQ372Ml2yav4MX57jJqo28Vq1kHkbYlZbYirvVI5a88
jfCq/IJBvjyfByPXPSl9uJ9uMX0d1XV65APtKAOLdNCw2qmM9klsANirL5Wu
v+disxdHjoFnFxuxovuzbNp/mPS/zYKjYviNSygxdFVoVMDf2CcKeIoC6pcl
vDGq2ecAte2S68gI1Dr9hvolGlI2m/TtBPRNrAW7h/sHkmbs0z+PrrECJvH4
4TIrHffyNUK6c+V+gdB12466pjeCpZ+KoTqNNxWCccRTBcpDShnS/Oh39fdG
Jy4hFCejpc1atLH7OERcXFuFBY6fIebVNPOrRSlPxuRC8E1vJs50yuGsfvO5
fXeIM20D6RZbqgTNVRuin+wL57BhvVIwweyFwgVNViC+oRiKaSjVbu7S5NGE
r2nNXTWa664OkpUQHU5LRiSjS48J4ZE7BvFDmj/+pU8iKFm4nRB52tGLzpzU
kC8ZtIkMFIyfL8DBxLS2NcWgeQP7WCYnFqfLccjCiq06Rnw+CuOXOl2ygmU8
j7B4AraEA56tfuf3vNpJNUROEEzQL7mnjSyFMdp7di1SwnC2mqEUzqnxWi0U
e1grpAh0ht3QOYYdjodM9fN9keHqgnBjQzOo+6tGMS/m/RtMVa1LAu+y8/JR
nSq00fPao8B0EcL3vupSSqBuCnkjbTMgRkYrAVjtVDRkiFrVd5XlMlHyvmoe
wGGA3es15Lr39KgKkxsZWD9uRrF/vX/bnqm71cGEL4bKaTQE4XRzHjSbq/KA
KdKfAbMbU41eTQmAOtAFD/WI7XXm87LOSj6pyq+RssaytP3Y+p569AbdhLAV
pDBarIwalsFm+Fj+boIsdSFNPmy8AC2UGv2a3voiNk3mhDcP5u31PAyjOo2S
0MbvAp2s86nNt6JUGui86kHVBz53O76VynTXP4MsRgHDJC9o2w8VXJWDvmnY
X7qZGmd6R1VbxPuPMFhExw5zSUaCtD2aPhm7BkVcmUJFKIy/QKn1T95Z8TYr
YPPwLFxI+ZCOWq/vuhgLs9nNj2kNxUf0/hZR0KRgZOyvIHYLuyuNacJiAwOk
xzzYFW9drMKPDwGYW6sGygk11cKRaLk23KahcECpvQDPeqInL61pdzeVjKon
khZlTTYlagX0s1VebD4bp1a0cy8BGN0gsZMWxX6R7ybqXzWvrv1YjPzk4S69
SY7xuAt+yKXiPXpXEMI8x5d4n5JAbdGkK3YEuBJbyeVTsh8wRuEpgexsqiLJ
X/TRAavkpepyrJNx2qeqE211mDYe4WS1QLN2XxpsqDqVXG6nGxYXl59vsy02
raEJK6zomKfKH2zaugVKdJuMojgw/p1704HaiVrbRngVlThghFFSiH+53Zm4
30AILFqeAcbPM6J+TafMuaTyjxZvlmFstonu15juchkVOrVcdIvmwxdT0MLn
ywAcFRkhByH3XG6pxOdAYABsySwaQdqHHE7evIgN7X/bttSjyZwfwUpmrlSk
SMJ14GAxp7lWFU+b+LlX1KAfpRFQhO0XPQAR8eBy6Ij3ePeyIn24l9Ah2dBe
fBUXf+qDA2vPqjiSGHyUnGRGHqbS9gvSUwqvDbYR+fmSdQvpz4IjVsU6tBpk
UG4WL8fE0genPmrEXNujXU0anlbqDuBv/E9Qsj+fdjpiGZjdwSM5A0BPecmJ
Gn4ufSFY4tYGJL7zKmDUS5vji39CdTvklIN1ODAlzCt/dcTHdUOmdDCo6fy3
hF7jXzAivPH6bsp97KwGbClD92UvmUdcJwXYLNVmJ1uEPNp1LdRzHSLBzFHv
J9hZ2QhHknEF/sB1+829iroiz3LB8jlgmuHDXngPJch2eEKen+El+i/T5Rlp
OAHJboovF4XtZNFG4QY9g+iYnzJzvlRtyeZUSFgE7yv/TbllBPWbvAoZvox+
qiEcE27VX6TpHx+gnmV0C8n34odjZXrXyxenJN1cxG1muTjoGB+RxTdSRzrk
eNkVcOQU7rvzix/yH60nRJ4cVAJO8CYORX4yT2LocQtuZpxVArNzg2TOjdq0
4+AgcOuZDDj+2Q2+xOgSWixnH/d1ke8SVZ5KIKgHgvzMPi2Lg0ktgLHP6BPV
W6ZOQlAaHCBcc7RTS5HwkJn76OXNO29qApTN+Ecpw5hsw7ShuJKS48klP5hA
p7C/0RBGdPHNVeXbcsjS74qezDzjxmTE5pPg79fz29/FNczqaiW4dG0CefDm
nVOBIJ72oLz5LbwHmkiM9AAr20ePMl2PuhN1ATGNaLe4kVGth3KKUbkWDUCp
EvK+fXtjKgl49GeyFAMOqlnxcPkwVC2emoVTQ7vgr6d9lJuI0TeMEuUSQEQE
Jvd2uKHyyX0aqZd0T0z1X1/pqoolbOF7mpkRsU8DTcPl9532TusQP+qeVLbY
/XE0coHDV90mKphhPIYyyHQyAkYv88Uy/Wbx4C+zuf1bmM8JipleVtvOCvsL
wvq0P4PtqkFvE7zFmo4rN2jHD3p+XYFanyEiX5g6r0y96PctVBGIE7VLYghU
swTYzWEzNBr/VLOGGV9AWyMcn2tFpJpJYuxcuUMSrYdUwQPWFDyCqhzOnSQi
/0nDalBZnh80Bxa/tOSlXLN6C3GT43Urrj4936RCPFRuAvu3+PT9veDEzZWf
ZKgMk0Rt6s/enOVp5OEIVlSZHohBtB12NM2wLbQUEm5wqdFvTLdVru3RPlvl
ikR0pYhtSrh+yZsBR6/i+DQekJWpBpygNy+vItI5RWas2jvovHrLEGOjmC9j
hUu6Nrb5n6A1yQLbFBfDbKlX/9K1Zcov3VXx+tUywwDPJQjscmtenJsurbCE
P/1w14c/5isp24ZV5T45/oRv3Inc9Gaj0PbBqWvCAjGkQGA4a/zKsHH76oBs
Yy2NDIrj2L7zV9flH2x+0NpSouhxzD5C0bpi+bSRmaa3raF5/Z+NRfQknitK
Bw2yTBS5mS8ggbSa0+l5/HZ0KA7El/y6NLSKFqApstOXfL+N0CGG06VgQat9
Egkfthzqs7foysEe5iavBDUu+Ppv77ZKRjIpa+8aDrlxpeTUl2+DB/MBQVZv
DAWREeYA48ipQD2P2CcPhDSLUfjtDg/lR0+Um+eQln4KCjEc89pHarEzDKlp
wZ4vCWisUk7IQfdj3o2DEtoF7mBYWXzKSfwKVBbEs0VOtbVa4bwLSlbTX82T
pvgccgUoWqnucljezLFv18hos49cxNUly2S236mXMlgzcd0+vxzX/lfEbFMs
Cv5LpfgEM5fFffwxIiVQUM7VZ89IW2qH1CN33lz7p7N+u0FTMiMWnwf57IJN
IaZ6LMPgpIsyQ7CQ7PCe5wlHYL++fndzz2lpeHCLNJt71Kf5ud8VhGpZKfaD
bjX6Yn8WgOg6CNI43ucJvjPjivjxWTfN8jquwwktSyvmHhIK/wHJPY/rKgUz
K6V3KzFl4xJK+tSwiXAZVDRfKneG53ZsbpYpnaHfQoSSc7DO6wIlMFp6dEvS
mN3cfK6AiK8Gz/nAE3T7SOlzKu3DPJ4072cUluBdMy79wVXPfXWvmvWUYd5J
Tdn/kDZGKRJWhJkxcgA7tEOCXkOqfVdL8ECo4mOXzYaboSWQJDURfZXide6R
X1qVXJtGvW9pcE0F5zD8gAdlTv3Ffe4Fq/jw86J1c7fdpNuPRWaxBs8WIEqE
KrH5/jmwY4Lf19bxJU+FtaXowUtH/xktnz6Xyp7uA3pFbo87M/yRHjB5Sfkj
WxbPL68O02/94DMiHGlOFphmA0ok1MRMdPCtLokT1feuRVyUR+5j9oP6q0F1
Ovz6a7c2wU5L+PM588FOFO3qXobcT1kCT4M+8ScPiC/qQ1iVIE8lEv4oRc9b
QAEQOcN8AgMLLdDewndVJveF07RwthqL8wL5rWbX5y6qAZRDXh8daLSkCo8/
xrGoZkR5b9hyWRHR5TyqwJxoA9+FsiwTsmkV6W86nVVw+9O6bwxhPf+DvkZA
3iSd6wd/P+/fdxOgO/3xX4RlU0qHCltaA4K43KhjPb+zNPEfTwYZmjvOJ+QP
w4ZvJR5CVlZjo4M49Vd/8/fRGjaUzds3pYkpvXkXP/8OlrkYamY9gYVsJLA3
cG7DzqreSlWM0oerIBdMh1/1leO4gY11Hyz7j11reXO5Vz25lF/cMQaieoaM
ZEpCN6g9cpI0+RbrGTU46TCLxqamdvFYEAfKbHUqkfkX8gJYLriUyZAfZrMD
e/Chl1nvB1XbVv+abnui+t5CkoNRK9rsEPa23Ra3HqW2/XqGxAllCqIkqiO5
PFvXa1ldBg1tCoB+Yvt5JGxD9nll9GaIqmy2/aZM2IzoSv5ytn6F82UMLc91
nWyNta/ydemJN9app4Ag4uNWc8jrYZ6VuXdP4KCxTQayR5hMM7tSGJt0Wyq5
99izhh0s6YEBiwkWMM6VwPcnBX8cg3RF6ea6KTOKG1IwAVK+HT9yK2Ks4F/M
CqyZpyhvgMmXH7Vl3setQEf4Hkv4B9g8Kd9XYFxpsg4maaSllsby4qIt+KlA
qKnB3Q+WXnAGc1ODTCFLdUP2Y2nyMxuqiNz+U/AdquVDHBgSPqoL/fNmvuYV
/PkQ9eg5JpbYkNkrt7v382FiNmyHKuNsKDuod532DvpUUeDRweTO9Pfu2WW5
lhYi9vRkti+b8Hp0yMKx1ybz6pd7cRxG6w9hq0pBqN/0h8Yxkh3t00eiSblB
wkGnnPL8LAfG00gmWTiiz7l+tyTK9NL+SwYxfqWYl3XPPCIy6HV0eskfc2Vo
IxRuvAvHLB027dFjeyPuMeOu4Yw8wVqhmv05TpI4gtoJJUN75yb8u99GTYst
2P2aCs4W+pmo1uU0EkJbs47/p0joHErpaZys3VUvyUn22OyE+41CVxaYo5wy
jqpMAA0Idg2iU2HO2nd4Q68y/I7OaPU4JIkWoHt/feQDrzqFmE8ZCaq4+PMA
8pUR75BXD5+Efa++VPIDrbyj/l9gq2lwjWG456pg+bcNu+H+h/x6bLBOxrEl
4fPfS3qY/OasiieCjRaVKnZupgW5bgUijceBaekBf5SeZchvlTS6fdEpqiLd
XITz2+CY3X0yvuuOpnW+x/IYxk+WAbH5FK39wlWE1zXJ9RiOkXOXCPZU+Zf6
hkHTE+TytqOuS62REyN7DUk70n9saOJ7ZF7xmDcBci5BTCttI+fNvnwQ2wIe
jTqPfcNkq2fFu9gFgkhrLqUn5leQafSKIrOuUHkk7nl+oPrXJJ6EuTEK2/HA
u6hV+ASrGc1qboKXkYHloN9h3QFp8AAXP8gCjg/x/DqeHonIWNJx6x+Hq6uZ
OXw7tmWmp4nJLf4IF7zkq9XNpMRvXbulJDBhraIoF3SbxKHrW6JFRt8Y25Ei
1TpkXwG+PiJJlYrMcVlsZCajFihLGsKXrZn/jV+GWBOHF/Llimw6am+BtcLX
jQgwDO6dGH6ofw8w2a8OmBIuUeFvT/4TnTuuT5HWeDareupKJhBdrllyTPy3
Q3auQzmxs9VbhqzgG1xfrrSlc//dmD5BQSZ6yPKshMgxpZD0pbMbs1pSYS2i
XcHD/I9WrgTiodz2NU/HIJLJkvIgLJN8/JmRLPuWmTKV9+6jibuXi3h0fFLh
effxmci/T/xVVeXM7TPhIbg6gsqL9T+lzjOwu8nyvi8J8aLJBKYrB+iNHP2y
fjIR63vi4dB8dVccdsoRQ5S8CnKVt4w3Xz7fQobKNYdhNVDWJsMCsTH8ZibS
zjgNifjYGzNkB9KkUn3zXnDwtOVioBIIrEgCuAGbU2LwXxKFzqGsZwjsYVBK
9SGQwu/g4uoXz7J7aLW5ftOfF7TUTW0G7BI9E7md3CXc5D26Dbb+1qdYB608
v/viHnYTSQYSu8bivDVGQZ8aBSlkYLV74wTTrZa1eRCM7Dha8CukpWv+nO4k
kxToo15imcFD3NIcWRKwbfjIRvxVULaFpyoATdKoM980i1X/XuqYSPGwSJhz
S+grPeyDFl6WHG7FERTohAqRAVRvPqa3gVRY1qlJZBdM8JU6fqcDtR/BQJoh
wepkGvHXHwAdYzxG7zRlfyfGswWTsQYjTM/STevyeefdK0KlFGaodxUUNmt4
aHXweBVhXqKmNn7fXwSgy/kNDlShJw4cu81xJ6NyYZnDWzIou5r4efujl/52
HXL3DKm+Xok2ivraA9P6kPQsEWtYxsr88hMcwx3IrDwRfvCNYkUxABsJ2PMb
yN523mjoF5h0nNc6Ivf6P8Fupo/ccwBcB9gV1X8kLiWwLBsbCJtkQUhu+dHe
H9thA26BC+ZPmJ8rUxqTxBszX+KkNNIz+3JokEZiVha5t4bUejLljzdKIaZB
FrCLiuBuxAzbqax0YSdigt5ZBc6hVYQbGiaOuOWWWINkYuVafR5YSxsVkTm5
q4SuDR6WhjGpjjOWJE4EIiaeylS5oj6/M86OfDWbdPaksmXaCponrtLaUlEd
ICYe8L2qMEU3ENXPN+gg9l9HPHqhDIFEDZZqo5oXukxH6UTfs5ECfZUnkpEb
Tvi3mFlNhz1xGXuECMf+SHbjBovZnoUONayFlq8ZsWvqNF1vy/7vizPODsBz
E6zwQ4J0VQ709PgsSlroaYKrDnm54xJQ9kqCG3TAI1+gPi4fwjNwnNGbln1p
hDPggaOc+oOYPd+B/1BeM4prM38HRDSI5H4/8TqeCKlSLCp0c9AnMeZJEO3r
xr0OFTIHyO+XkGmGPkJro4DLdLPpnIYqybimywuW6tINvXVQi2nc9PfVh4gf
nj6pprm1VqSd1JMyGjDE63PSsx5XXnvPRqs3tTkGAQmBfBEW5LjkvBboVKBM
qFWrLETv08KfiT0G3TLaBHc2X/WgMVBX4uEJDpjSiIHKVN9BiX23XcyWM1Y0
xewbci80Rzrm+v0YAFT1YZMI9OJBwNeq9WyI/a4sm+fSlBfih3mBbBSg8EHO
lTS86H6CqXH0FuvoXi7q+iqG2Qmxlzec0qkABlp/ph20VLTvUItl6/gBn7PE
YyzkWz3lztbWUkL9xe7hImc1T5C2R4o/J+oLdy5sqdVp28PgNDN2VJGGWErJ
rPPLYZIBLtHeREh2Bo8Yk6QYLwEAFHZTSEbFeu0tg4bcCZ1ncjkunGrgQzfc
/Yg3jWNAd/S8UhL8IemTHaHPXonZcA1FlSvCeWnOymFleOsJ2Zr8wN7GFGiw
qRChJUa5aaXdje1/XKsVLJPN+HtPdDeRV8EQaEvJ5Fsf/VmUSgIcXLEOJsVs
WTBnd1HOngLJ06zrvip7RjAPZWnMwTkZ7EBOgYzDG0WTptjOr9bqEbh4/dF4
4qO5h6VbREAkfgX1wP3NcMMm7SOezR9hJX537cvztNJnZRoGwkUIqWFScDdC
+LvNgAEPamGy2T9qmroxNo5xeass++yhC5npi2r2oym7sVyz1XZV3kgasWGw
OKhaMCGwbTyhldRYEvzTic2zfzxBULUL8ZHr99mh1MdDcPmSbyqIEwisJVGL
i68WnOEX12sh9zmTENTJCeOGF78GnhOmqPxIcnO8NMl6HnA8fFlRr2JUCt7F
Mt6d0wY0Pos1EtB2RTSYJW72cnpkk2UZXN6+kbwNpknJXTyrk4+inZTe9wbl
vbpqdV+CtzHY+RSuPnXHW7Dk3V899trTDMMzt1FtmRbPzWX0UdxitLSRx3NR
8RM0rAmNCdldzyor15YlLsnI6sS3gepu8W9ukWx+BIpoR3acIJOC48LGvty3
9mxJPGUsppn+2E6Zvo/d18En7YOHtw/lLDV6POgzfTijIiGMlxT1pWK6WEIG
R0TC33TgwXPCAPSNH/S5ztMLXNDytO2h4GxoDrcN6WfTPJZZrvwjoclEOZni
lKVtZk8qGmrcFDJ1IL1BND9ckoStttpSt6XJkpeOeTzr1oXyDKYt2QCXSs1f
Y9kI6SnDRYXSNw5W0SgLuPQwdEan2vGznn5e7h4meKnC4cJZ6MH9FXS28vlR
qsqDtVgJjhL9MRTqlq4JiJbqUpNF11ozeMeVdHPXpcyMd5gYrSnOknX67Kbu
W8iynWSt6jtp/3jJpoKNXUYDkd3vWw5eaPxFylGXy4Tw8eQvFfspAJjPygTf
uUBigyD98/8U0L2VAfm/VdVeNOBYpY6FLsfabqktHzu5583b6+Ti0ZV2MadM
Drwvh2TdHBeLFxA88S5TFN6+y47hgbR6IwhZWdnoXp8qHqSZIiC+3/DWHOMj
nwdysEkxlH4rmpPqsOjuSzUx3lV2p7bxOBW0yLQHt2hzUWGgmzCUDFfTVdn4
2+dsBCQkc7SDK0uojDb24kAwsRMSxbopAb23EICmL47570FLvbpJljH7dDwf
d/+8VyW6j8w+jcHQ2iHvuXVoVSfZTjRSVSDOW15Qkw97gmaM7HhYvpGH6xh5
gaYHyaoZhO+FLXqlAmOfRAGekZ4nhjtOKDlzJxpOvc/SrEUbShK//SEdyDGx
WxK1kPpz/aXqOyJB4JRFFGhdFDsEwyMmNFygreQ23N/2Tf1fMw5Hkzy5sbFk
IWk8KL5YrsdYudz05DbGVP+EevaHBAPaXXdAcP5zm8y80uvFkdRIgEk6CZqz
F9tr1YVf5Y1WbzQa9G9HtW3KU8FH7RuJUg8I55cde0YeCUVEeDMAGCNt8+zo
ntSpbTxLY1SVbdUa52XlL3dYlTB/b41v8ly0Vx8CLfpxPqgH2PkNZrdIiQGF
iN1FF6vKwqEzXjF/CIuPFzQZjyzvs+WwZol5qyQvMg1iM+/G4rshmrkyfvrO
K+tAE9ROPBgzbOPgbHbwaZLl074WqrBkW5SjSvtL1DGcX1d41ErszLHGA+W+
Bh68wSdLUfbTFDDV1+dR36TM/zMLaO/FqraBpj+leUUrmDRGxmmrU5xIX4TQ
lQk/t2R+jsJ8CnOeyZDrv1+z0doM5ez05/1nC/F0jqrVXtDbgtmLeAqFqvOK
TKicuFfjPrToziBmO7p42IMfF6Ib3KHv2CNOYR5/mz/KGbrpr+WtREFGUy9O
aSEgbN6ETv4ldBFj4MgRq+ayFL+Ff9bOUoysRI7fw6J/Hj3sVaS1ViVp70Sl
iQL2w7pv6cbQDjWrOfXFVk3lTLhMIlxs3UYWfhGQnp5oTJnWlhEr3AgWYBAd
RVyukok503gvc/2uhbv3CPDEExb+SYGE13Pa0mbG+Nh1N2T+ZsGrbLsEc1J9
zi0j+D+vkglhxoI6xXGEH45+GgceJMi026xaT0HgMsmsLBN9ONGx+KGgqJ1k
4OWifi8WbCCK7NwwisxoVRd6awo2sCvQyXXvdxooZx5aAygjd8Sh+XHwSnij
m9FEfD7ybBZR58K38miJ2wxP0OYfGIqUA8lyYgD/L4GM9xr+IEkBIThExf1o
mSmldhs93VqRujxRYpmhXpQtv+q7XAcygS8mXS70mRq7teN0bhZQYKojOGHv
gXXsKW9L/AgQJlwyr+qxYT5Y5xeNo6gE2M88ZgyzIKZy51+bYDFphW8QPLH4
YcATrs2OkBAjWQuK8R3Ib9mi/WO2sE030OjgwMYlqf4Qk1egR3oWOcZh1lCP
93gkrlsSFmWeZ9Kzp8O15CArcoj2ucsEM4p7rseoLWlzpiKVmoRK+Gj+INTh
TwRjN9dbvd7DViW3NvQRhBs2cQWZEBkAGO8T6hTxhh0mi+dp8vqQ/mDzdpE+
6gQMow/qYQQkosAnUclPv3D/pyt4wQ/ZmQSkG7j9VeHWaiLIhz5XzoDwOsHr
w8rrrtJvldQisBKrQ/n+FWXiJ452pgNQ9YYUs4uX8cDqpSIcVuGhFixBITin
tzxQsBFm28UyI+172w9sZNhCbd1NUnfYrOtMMHmE8BHI1+29P5fWP0GBlh2B
BIGWXuqB3Vg+qLg0LKO6penIsrj6pr9NMCx8PaScPzAO/auKxRkGIboBwnTC
SRsCiEUabkQ3i7b7/IpTRMYBy8xXyex6hlPnxfUqC9jWE0UkBPvoaOUb9B5b
vTBaFIBQSa40jrycWf2I8IxQTPDD3EhcmmfV2JBz6ilJQpGbHUy8uEPXpy9i
qKAAKQ9lcg4jawoG/B0Me/6kvCSwssQcI79e9jR9mSXP5irKqHrTkcrU7Srj
VZCreXVNWLVE0NzDjXNhbRGRcLcrv3Q/HILPyo8ziRsE2KKqmpW8oguX29Qe
q1Zqdd82c2Rqx3j3ARsDBIQUUUai9BXc5b+g0Rz0dHBIM4UvsPi/rdbA44OQ
rT/l1imuCq5zfombc5/k0DM63UhrAlEt9/qK3g02zzxzsVp3IYxaeuHy7Az2
oVEuXJhF06nsMec02qf+RqP6w/7nIXrFXuvim+5q0NZPLW09wsHSII4eETvD
P5szKMKtq/EpSqkiVgb4KTwWQGMY70E+9mOJHw4BM1WiP+PTyojgnAYITku1
3OYfrr5XACN+oQDFN2DVpgNzpfCvwj/o57OPG1M/4dslwpEGXt328ZHVuFlL
9hJK7iQgwZ92gTrLcZ4MLNhYxohfnnQw0zN5Xgv05eo13NxCz6avee8jbNWA
qr+Ht5wRloU4ppFeaxTzsQUDgzKQgSqvk3eGmw2fCHX3MdXUxGtCA996PLWy
xpVRA4LtZZi3vg9Mno1vs5LxqR2cFAYVWxVoWBsK3g8kvv/MAmUCm36ntsRi
egHrcpcxfxOhApt6hUmIr8Dy/oyyiSPi/JmtzmNLsAKqjw0c1xQdhgSftU6v
/MXu+ktXgVkaAIj22YtejModkUZp1/zyXlq/NjKwCvEoQ6QBtx3jb1GhXrd7
jeRlqd/lkg8+wSOq2KfooPxT4d0odHI+5yp3dOJP+cP9JhCRI4axucRi8c5e
mwxYsaoQkXFSH52TQEPk99e15XluKcTQYL+5PXy/gfRpjsFqKfFhTTkb3mSP
2LfWRUipazUB3uA7ODjU5Kg80gJleL3/Mz/hqY0l2dZNwB4m75GRMtEXx5DV
n8xDmnqLqhmEHf2rA+mmgPMFgwbgdHvGpzdOxNl+zi5DRKo78s+T4tx+M3PM
0ew1Yt267XBV7SotamSCGcsBhXgbZnNxe9QDKsgbHElFA60gesVjTXaeoDVW
HRrNgx9dcvISkuxVKNkh9+jO2r6jfgiR9hx25vkbBP6DMBXiw3Ih4t3O3QyM
L/ted+234T+96S+lC7LjoUnGW2+gdLJ1B+hdVOebkgjeKigTZ22tVjB8a/Mn
UQ3J8BNa8WsKLsfUAf6zlLSkwO6dLKQK1++GyC+U5DGhYzwtmu3s4YqgvnKc
gk9E4H4Qn4xK1Zr3g+AUmbBGT44fIupIy4Ci0eGHe1dWr8iBgByawUGDqS4h
SZ241RJMf0gfn8H3MfGgVjAsgvwZueOIGnVUfL3ljhHXsHKJeXFg+zBdZzd6
//ooVYaaV4poJOyoBAjoalyCsAFUQsVVCDl2TZD54VDs3LwXRisVQi1VgAIf
Zm+oUbHQeB7hj7U4lceVwPbRDAcVLsGTy8ME/91gMP5z7bKsMzVAgxB8KohJ
MzWi9Uo95CzTC0JysyNv0QT847yu3YX0sRNu6tErV+tcvkOqcnjSwhcMVeKa
Ekh1C1KMPG7amqyO9kIiYA627vrIzauRXFE2k/MmGQ6gFyx6D6xibpxPiMc/
Buh6o2BXWID3+Ab2JvUx3jIdk8Lz4b5OwAf3bCWhdb07hZZesCb3CPXBRzA0
J8fe/+4Gk8kETjPMwk+qmHldMf7ylE35dLQZ1XfZBzaodp7FFzJIJ1Q5QT6C
ATRhSjLdqaEFV9JZLkSM7YaAD3R3RH7d7Xg1iSU58s+umGq6VD5wyob87hv/
6rkp55lOcYaaaPEb/FEm5NfmrwwIkH3wAFD/t5Me7exwrX8IE/J8Um6J51WP
QYxQvtrSa76Fm8pAP62dSK12KVPuTwUHCtrr5fV5ViP7vKv2Sp8fi5tHSm/p
BP2OXgW27qhCj0zSexHKz/tOlGCngCHpQqt6Xj5/I8Ga2wIUfeshBTHxxBRE
SRL+aAakCRwZTwB7SJPvjlegsHqoNPMzfL/Gfhw82RF+4uE6NF6uNr2t93YG
+B3TtIhT9jjMwpLjEGNqvKoymJZXcD11iIMYOHw5t04hs0BS/FR4bN+r50GM
5h5IH6JjNpICgCMZcmHEN6hoZ1mGSefejcD+1qZoqnJPtBT42t1IEAB+Koqx
HpKwdeINJEaRyBmmhxw8OOWxSJUGercjDt2PhUg0CeQAMBOloL6nP0BgrIW2
FAkOqH4o6M45KaU3pD9OPnXJmAFYMqUAPDbdIYHVK5YKpOIG3Bp9w6V8iTVd
OduZOIM4ZIYlSv25X/f+ebymi+bCf0lAWD/pK8b420K6L9KdybCI9lCJL6sH
MQ1X3FFSILtDWLbolXLIIUen3ATOFMqkFUk4qCbpmXN7AXxe2Y94d1JBQwqr
IkeCT5RxiEjRCntXeXxVFK8PwAiU74ZNIsg7Ktiec0J/FZyqWTazrqNbBfRn
EVwrrJ3DjGaypOmoCVFTjVnL4k4zuCXFyrRd6a7VqvzapwWe5vxK+o3hKKX6
Z6ldatKL6GGV1lMA4WZWBvUdkQe00LpMq62RS/4X1u3+geDgDVTiFQWuFBVL
3KUN6tjByA6PojwxAIVrqFP0VOFKhtG4V6HfVQzH2VE3ewAE5LnPBXGXbQ/v
wB9JCDJqAO2SkLGK8ONPB9vfeQ88DQrCnU4OfGecCGjqi1O1qOe9E2WOfZ7C
h/fuMEQA9yMpoxfYSOQA20dla3nYAyDiuhMXFLd4wJapKSEcbXw2KNbRcZ2Q
qukEEE2z9/YUbXparCFQCpFEMg7hiqZtJymkoq6A2P5pMgEpociAVhIKPjuX
+axc0M339zL/Mz2oVaHi7ma4Y9vsGywhH95RCc3KjJ9syxScAdQJq/Ki3YyK
4EjCIy8QPpTX0uvnkdNPvprEo0kGE74U5ScXQ4FQLRT6lVsbE4VvAhLlqY3m
LEJNiCIks8B1ZiOF+W1OIgfzLj5LizgwFkpxrjGrCj3OBOcLJjjMYWdeKLth
8v8G9DobGBbYx/QVteOtjwbAPXNIwD1bovPylHu2n+rHcfccDftRUJ9nToQ/
M5DAHjntt2CiLwwS+bSAa1sXNaColHG5EQLUXAe8cWmps6PhmzaYDa3lPdQe
Cgm4sk74kUYmlQZ2LD2jkeJNPB6KNwV6m096hy+pVGYsCJ9Zh/5x3FOmcy6L
jxnrwUEg3SAPIkjV0cuAZU2C4Pvb+gOjRm/lEdWKLo9E2iHfAuhd4FaDBVdJ
tJNR81eBKqDe1FzZMbGzbFNxq/UVOvImksvfHjY6KS/ifFxPXcTGWc77bREg
i4HA9KJU2Ow+jIVS8p2ITHr4U2bUwrJoyL1hXSrvUD0Gg4RwyDsF5/XyGFWG
FbilK2DmEGDfb4cHfksdBlc1svIl/I5pdfyi/tiGGEzsYZvKXlitSW9QLpyR
st2yb60HW1C+uP9O73DTiUVeaA0YYyPKjNNM/xmi8n1HP52GXsEq3Dzju+tL
qqD05zBC/QblhRPaArksJD63zGfsrU3XBvnXV5R9C5Ol1tfU5kZ5gB9Gdyli
PRa4mDTqYdbU0hdkgQ1B86YLO8Fdiy1b/TRLqSgswSuNwefX7HKKe/ssvt48
GFCHtGaJlCXYo+VsY/71sqbXa3rx07Fk1sh/32dP99o81ouFNRwcIFRxajwY
P7TT6uUyH0nQq7jDm1hDrwZ5IniIBRC7nP5L5U1Zv8cT/xbXINBEE8rbGg0j
UI88C2cw2m7af9tjq5QPPrMDwqDy3V4ETv7V1sCjBmuz8ENbULEOfYNhsYIP
0ooBxyifUIQju9/Tt0/FYr/0YT7FZxJBraowua/iSIUrg9iqtz65vWGIvL/8
4gJ6TGA7w53KehcQ9Ll/DYhDn+0wmznqP4uDNlt45Zq/rgKRqo/12U+FzWKr
YA2GqFPyzOqWJnoNKehslbODLM2L5ICgiJ4mUIPqXoklb2V/yBkj72lrgYKX
P13idJPgQtm+lwRO7JSN8Tpe5o15is05HhKU3HVi7Bqqj+iaEGO0lV5OpYBS
Ga2VyRF+WeJBJvEjPuXPFbGSLCGGU2NRBonM8hggtqDLkIDf81iIX3A3jc5J
/aPXlN+JAFLAjUwV18qxdO/ZRhU95kq/+/9Egk0jnT5JLtXMbCoavGKsXf3t
/Knx+CmqQGBZrEPVPvtyTHysaiT7Rn+d/eduQXRCxoaZEDRTrqJ5AHNFyyaK
qri91BPhThMIwBlao/6VM8+zlQtjC7pyX2y5CrihUYDzjTIN4McQKn19Cl+5
GToFPJMNYz8DfCr++JPsI3YHH/wONXbwcLzk7e5e7YeRr8ejkiboOz418iwg
8kzDpAT796mMNUSM8q+IX+D7BpuMs43dgX0GyJfF8AqXpB4c3nEfcrz8cRQW
vfFEYP+C6VFLl8pc5E2APaG5MhLxO/Dy9vrsMbA4YSmzgknjnGcNB1LgXV68
GztKTaEVOVM3YkxbgMH2UvFaAXe1VSdiZZJu7WPp4U7Ro9sZqrKV7+E4csu/
IvyBS+TPZxxNGCAVwHuiEQygl5Pty45jXAi4x28ZyT03sMzqHXX0CsrroR20
VwktJLC//ig3MFbqHMLRJg6+kJIqzM9wXw/nJnC/E6iLFc+3gMxTuSs5k9hm
MhJPb3fHdj9r6esYjRKMv6R0hx0C8dNTvJaXYUbvjwrGbhMEsulLO/ZanWtN
3FIEaOWX6cGp8X8+rGT51IEjQM0d6BCqsDF+fSmWX2K98VZ2b2lEOgj5AqXj
XpjkiOS39fhfgV5NMvSwPfJtoSEcZyY/HXIqmQDItp3P8W0EUxBLc1ajS+MI
V6QyYk67ahaoNLK5DmOR6FSbksoSMiM+twfUZlhOdg/OmqzDIV4BMJuN5G+O
hqVvZPaUoPaGe6ax5I+pGWyeqLGV9L9bDSjqaRuZrYK8kGPyYX6WF8RIJbyM
boXNwbrzAZXPYOtS2tUOWjGl0XHXsbqo+dFdTnHfYJAEsyjRfg9jzt/A9XUX
cv7nVsg6Og//08TyGbsy+u5CtBHsh3ZiMIDBwXDAuC9bafhCBlXQBCc6zT9B
ibNT4IiEyYiHYbrFQ95tgKeC5UHAI1V3fVyI5ar7lSIw+z+ny3O2BhRpExKW
vCxNKdPgA+wSA8d68D47PDjO0vHW35rEjNcnH0HfaTJC2BRQJuWUj7eHphdf
RYRq4Ls+OsEVdvQ0rUEtj5uqPBMqh1yqtelZBejgd8Wrj6RwcVwCX97eyX8a
nLjV/DbolBGs9W6k2GNpseTwfqUOCvwJaZw11FBABieTeTD3OUsdSV79Dfd7
MtuD41zSs3H2gvgScH6cF5HQlbTMjqvQpKh/pZhNo4jSeY5eXlPsb1SlY8RN
Rl3siTCbvfeRtFtTX6ZtykpEhAu7pVtZL9QqyoHCxY/KPmskmjjBYfrwFYdh
RdCkJEIjoPOeuXC0nemhaBFS3MypdXGSAl94CbVxC0hbMv5styhnXVrq0Vs9
aIUbH0buTUH0cK7QMrZkRMoOQyzSsM3sVcJQQJdnCQLghb71Y1/pSJ8YQud6
gvz4aku3usW5DFys1I6VYmrXV2fTcRcS+FbaTbvfb/ry4XXsBq0N/xMMhx1V
az1Pu2oJTYkorC4psidjFW7Sgc/BylEPty5IRNil3ihqEPGrQ+tEoBlBxzwl
nUT/kvqVnTAMYPtNGrUx3aG4KataYGrvcihk7ICqUTakVUFbyOdPPQIeUrBp
heyhDKZPaIiZY+9DxdOEYBYkv6d0i7NXH3wMY7LsqyHlEpavYRD3aT7G1uQ7
v3D7W5/eNCQiYcsKRXGcZHERVc3U/98zXj+IhX5qJRO83v8RWQ/1jJSh/OLB
o/TdvsuHa1qxxKh90X/w5fY75rYsiVJJlyu1g6Z09OSiXUfjAzEZNj3MAGgX
I9Ps16wq6dKruKkaLpWeR7IUjiAiOBDvqdJLygBXTt67jYXZBbokgJvBbBaW
hRiTF1IuJSxn3PI0FTn6Lm1jbW2a3QZRMHxyEsmJMeKJA1NCEVA7AwGdc+Fk
69NsD/iF4cjhVWKU3Jvm5D1XJj2FPT1zCbgDZeBLuAeLST75gCYjzLDCpXB+
fVqIzrwsvbnnq3v/EEqgo+D7pjMt89au6tUbx4zi4gH64tBnouRqMnSwSdcs
DFeoUwqKhVtbJFoCSVtYKT/Oe0pBJJjBKk5pIgT4H3hAXRHF5gEkERAFYb5k
oq7FqHeS4q8Rw3AP9F02FX/cfkD3wvLPvF5Pm2rATII7uk8ytiuON8K/0Ky2
vHqpOJH0AehgUMZ6dyvr6v47BYHs7V0/Wr4UwnT/M9cmp7kRqJjoFBWhpy7u
ulcxlF7mivtmCQzvVwD8EYT0zxSLiUtBKPGymlraycg98YLuq66kJ6xk4WfZ
lCxp299JPkkb2Erncrq9szh4isSOmZyZeI7T9oKzERc4ATc8CWe2fRr6Exwp
B6+GcJP8SImxh7CxoKEwvkn0hZXVMNhfA8vPicZo/DXvcP6hc7oSraHhdnUj
eCTdZb6HVbzPFg8oKRRin5jRH1K3lR2QPhA+u3d1gZeSsjsJG2osHEZ34YVs
oENWkfzYqnVyXlH6+7UJ9EAG8CCZOnxd3aRoec6E2BfAex4ra2+r3N9nSHJb
tfGenOWb29w9ewNceyRBrPoyEs5GUy3rD2+aW7IaqqNDs29JONFNQEeF9p4d
UjojM9z9xFoNxAycX6t/XVQLs0OlfyWbWuBgbZDqmimQqv/BDZawcJd04h+X
8HAP6hJulrNCc+uP1Tx2H8jAmySnB5d5VlfEALZ7bhr3Md7KlMf1/EJXr24K
oqMA+JbEddR2EbDg/5T6LsZz0Spe1UAeATajSJu/bMaXr2JyRsdQwfmlJ3wP
UuEt9VOHNOt5J7NJWdwQLT7K38D++XwjL95KJGgobbGMh8G8rOtKCoXWl0x8
DS/HtyU8kRdWhj/z2yGaf5qSWBmIEoQsCt8225chaGICUTyiQvYxIgUcd0L7
0y0DaM97/dy6pZoaC405ArONVSjvFs0T3o9smoEdNwl57f+v3AQClSFMUps8
muI/C8z9/otxtT9cAm/HQbrgYXyKbNq71mpa1ajLXQYVsaUfW6MtZV+ML3TJ
lSFjXl5N6wPrYzdRGFVjxdAPQYOank89A86Zl2D09HBZCeSg8PLPSybnAdjB
tyOJnkwLLvrIO0orP+tkHoyO8mNp+RWogzrRP1DA3bTZiodzYV4qmITokZAo
TZpolIgfgcLispBsxtHXzPl1JDxkQwqG2o2BdsPsb/9K3kv+Rjha5G+RYsZi
0EQOaA7c3tJDiyZWYue70t4xtt2AXs5UqKtmz/ZQsqGUlFj08f+66qIYKpLd
aMDx53TW6HttjidBm+lLv9B/x14OFE2eUVgXcPshewlgyMlO7XeaHR0l2ke/
jPJxEPIZ72zptw5Fmzy3k6lkkxZWEt8xllHPS11WhgOpZGmd+t5NbnspGQ9V
AvvaHJ7DP6uCg5KLiWlrIJ6txAWALZbE6tR/WOxRkkkBDFQ+8FpQSK/TgShs
bAhusGAMRtPrn0D/aVKy01aG9NjO3ZvynjA0t4hi4vyaORRIyzLa6O0NBRhB
pBzPjJib8I/cHqeWl/ovpnJzliOzUfbNrg0oy8PLhymf/877dRekGjS4yV0Z
/7EverWarAuKt43uauxktmWYkJSfNTkGCVeeH7sly9kn47j6/GaiaaIZiM9i
kSYUqE84KAPVNCcqjRJtSTGjIuYdidveWtMsGMDd6VWWUZ3j6c2pImYpX7Lj
1nfVZM9SfBxiVg/kJ6idtzY3R6y3K4Xex8NZ6MSORJd7C78ieRWHyDns0uJv
LQnxPBZj2OrMpL0AyAyLjRv00lThjLGU/zNc8Og3nRshLsXScFU0dwMP8EaK
34wxvEzxCs+QKeoCsvFVBgUXA/mUqLSFln+Cblwhyd5fbM+f8nUUxLwz6Qzh
eI8Iq4Qzfov9eanNVPayAsvBSTy3ZvsLpTYZIek+Qs1bBZSOpHPH+8xTdtKD
wkKqZ04Y8WX49fzltUAMgCPxQVZcagtVxXW0Rg4aDcc9wZQb4EWv6TbbMM6l
tKSxT3f0kjZnQEZHyqXYewRwY/vIW+aCH8z64E3rU7XZ6dICtQDUCH8RgNCl
4JF3L0VtR7t1s9kOD5+nEDTP4yyJOUTqjy+k2gZq1cBbnigQHwkebZN37ft9
D6Mb2a/3dD1Roy1sJ4gMc+TSccvjnZjX2sA+J3lGElbrJNJZKObvuQfX5aaO
S7mwk5QjccYy8V721SzPz01NvadNkBwzUCio+BXSWPInXbWVrtkBGsyjdhFI
g8pWwCjzp1H2VQJHOCkPKS587kyRE+Bhi7MQuiXVHMKa0hsrITJoJsqIVUxx
2e56FyZiwMSmVz9u+YW2l2abEpWJZ1ob1TKfrZr7pu3bWHpWe4Sh0bmIzHBW
PFlk1TZjt58+pSoOrR70GXIO/GMqDyFA2Is2rRH8gyZ5QFkfD85xRDCt2GOW
QDWHhlyF3pWHU5afP0XfvDf5xTB5OK2R66LvEKNqldosOgJlrXattfTdCYNB
tbFYxNIHyoifgVJUWxqs+0jJAcXH/4b4kc+1ySsMtgHW4Hxt7JnMTaO24VXE
O2wZYUBi2hLuH3W7jMNj2qb3uUV69H7szrphz9UvtGDnP5gwsMWlRUQKSBU9
4BeOYEVwY1xbnvRrfYyL7JCY0qKkgPNyMx2gjZU1wj/DOcBzTEMnanMDK4hL
eDIVrjNNlpHGcR0CWvCxkxvlRRwgYGhpUBNtsyJhybAOD2HVqUFGDHtmUISs
hmoCVtgx2uTXk0g95lMBUgUU67yqT9gudUNWwpuv+YgNVZXfStBuEUHWllo4
iTkZKoqgiVpSzDz7X4Sr37V5KABdN8ndwlxXTA34NNSswHW4iLDbgvH2gefw
yQnmha/MpNnpYubxEvlZpJTSshBaYBC0HApsLF2sVAzjDmn8AhY9dN1uECr/
aWWcmA7LSqSYWAWHveE4qgw9ydZR+qOKB9grFYmuZrGHqqLY8cYrDtEBG7eJ
cWVe2wHJMQJJ0Xyq4CXbmKoedbXU+Ua1yCGuOuhRn/xA8fTX8EtadYQ/5Uib
3c1aq8edrnjWsRN/Dis63WG65qljFBuWpAtDsAMzlFIMmv68AuWEnkz3mkxf
tEDjcDPl7esuHFgZLQTFdBmCFoNZlnHPpisw7H3moL8yDsUYK9AkhNNhqVRS
q870ACaELCXGkf5o0TYfpSq4vcG0FUHyMtOXky1SkoQs1wj3bE3d11kAtr0o
uG1YhxVshBMI5FANeKLBI/xNCg/OQrCq+cE6Y8yuLGe9ro2QK2B0RnNnYXFm
DOgGOtxtHsjvxeNUdjdlzodPLvFdl4IUbtT/PghfQXlyTAeIf+SqXm7OuibH
mj54njvdJxd/K4JODYLoidkb3kdIxDwl4d9QXEvNSU5dwr1zWrkY6l0rbhIl
xrEL6cgSuP5/kdIUmldCHqZuHIq74sgys/KsMjmpAFsS54nDvtwHMPzWpB1r
BApNHKyk06r/SAIlFMIoQWC28eum3gHHAim6/RKyg1lYVesTcQPRrSRbQhFA
0JSZjUnurs5MovkEVnOjE90hFE6DXaPAwlzDY9PvdioYAGHMGyYY2go5MkVw
ZEdnFBBS17luNOEQDHTqJgtHhmTeGBmvzJ3aL7ZdPnq5Q/cah1hA/XETZXgB
bB+INC5LbPt1YvUxgopcwg44WYHq6g1ieMF9u1Wa+7Jw68q7fH0JpikaIThG
2lo2W1LvCyKqWzUSqnmGll3LXTzdETGBMuCVX67SeLLivvIaJF7LDKund+NY
N2/qJ/QmcRtPuORIkNp7vawB08vNPZ2y1JzA8QSWBM0+loJrOTSZkAsfPXAR
YGAkcRqmHig=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EqTNUlUVcVtCauP18sPa30zaFB5nBhfQTwCN1G7pr/4KLzXiwmxFjei3uvWF1LJ3330FoYhbRniO5STV3QCHqkaYArc1zCCu1+1TNe7Ea0GDHFOsA0x6JOdcAzCNFUlQsoLPD1LkGUOYK2r8dFg3gGTlGV6tWHSFLwF5hUDvGSIq/sIu2tVkKMKyKyGgLsVXJrUXwoy7pxsDIDo2Nk06H46h7fONdXtBgR6h+GofibP62+01YGZ0+bo1BdHvQdrHDPmxWlgPneN9I5/yo7PUpodHw7UcBThlB5/2qSZbOKrXJD+xkJJ0hmZoZgH3+GxtqGcJXRCiM4NJqzc6Ionfr5y8LerNC7TZSGbRjhmDyg2LViv8pf3iEPcHXxlFGrR7u8ZlhqCRxZmn/XWyKp7QMi8d/nHEEFVACeS2F4KFNRjpEt/mN5ZbB9xNGHkB9IgvffTww7+YdBKcGroBw0F2m+S/7ney6QufZBJjWLdIJO7FGLo1BvFi8rt0xasJ81Z7h4AjNA2RE1WrwwKQdH3/TXXUX33m4lhJDNOXmj3glxj5yHvNdVHUPjUFJFG9UVZ+t+KJrp9bN7/T7tlDtGmEDkZIknxy7kZtEjJyynLznETmivqqEoVhB6tPnf6n3dAMkxL0EXHZc+QiDJjGjlNv/OMd5jJIWvuIgOXSSe2HeocG/YYIPGhuzUvvHp27Og8Z5tT/6rlFPMIz3hsXEkPWt+fklYLrvplHxuheMUACy/I3xg7lA4f9ajZdy+oTlZmBveNogm63+FMAcz4XqLKZtS6"
`endif