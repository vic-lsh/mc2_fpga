// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJkcNnACKzROINnizsHuHT767X18IwZbmZZPlbU7+5/ehAmuLd3qjVL7Ij5T
DTRZ2nljMNwgESf2IeNsapyxM5OUYPCGfI9tujJSHqKXhYMrkgVseAp/VAyH
smRu62iBNlmzE1aQ8eX8t70wbD6AyhuQ+YumFaGlV2eJ8HmnK4Cm9MmnRen9
m8UEDqc2SlT1p/5qMdsZJDraVVuInEilCyY+shO1f5rHj+e2eTya0YBrlHWf
vu/0J97orp+yuPc331J0lY8s8nEZGcXlNnDCHaP5f9J42ey2oPHvboaZ1xVC
tx1iomsRNPdi+EnLiyjZtt5yRJTPSDvQPAOmykkQTw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YxSIB/jVyZCOsf6Va7qENwIt5Nsi2MooBV46sIsXfdviGRzJeubrt/88TzHD
ihXftJkqVgW10ereuFYhM9Y15lyCBIOaIVZmAD7PCOBy/S1Gb6nEMVVO+gj9
ii0cawSI91Xcli8DV9oGwJcEE4HN8Fs00LJi/AXDqgmSVOWQg04IpF+yjTgK
VZGLRlUSlQPsTPBHSwI2Hie4HqItzMWEXmBX9lrCulI9yLCjzpUmQBFIyI5Y
Ro8SFk4yCymIe4cz8ZUnVUKXTtGedOFdDOWtjvvU3XvlGGNzK8pvMv3xqwW/
UTKGoiB3DbVZYherlENk1hUnQtmLle48o7VncxK6Mg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AXx4jQBJ732R3+Q27TQAiKpfsk3gCqn/0n89dVIJUNlzeOwzQThoWfsJvUo4
XfkWk0p9NJrPBihNqPPchRnoqRhl7waTxVhmcmZgaPoy0go3EWQJssa4vvwY
QAgbLyk1pq6BHXHNJqBkne7zHGvfjgc3ibh//8dJsKtn9FtnyLtJnM0Ozbu0
zZJBvSw7SHhz9IytDFmU4KC9CFjZdNHyCGBvRk6aoZepgRvvuKU9SKYxAjfd
8jWVA8ZyGj9zkmWX/GtdWvMlVFESrPmVEXy4t6BIE2xll7JRODJxrVv1WT6a
b+VPEP+YruB4DFJJ94Gdl2C5RLvsK+InK+XjIvgxuA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nkemEbaVJb+nPsv8juCMpaMcV4aT5VnkxCcUvYBIfW3muAM+Gr3rCNJYqIhd
ubJruM+wmnan718y8Ip543ZDgaC0LH3vqug0Jo/xbTQF8K7VU/5zezDuJMV3
p13OYU9Qzu0DKQruCdAdOyNTtkAK3YePdrB3a8Ni6BM99naq+BlEomk1XPHM
ZUkykITGTKJu2OOmDF/K3b0+L1UpUXSnSll7zETayDou4KyY+2gJAUH080qY
pNT3PA81fqSGkiUdXzk+Yri60pCykBPI4NgmAULoDqGtY/KdYE8wBMviWVXn
ecpBI9Z2glqMXNTm0VyT7O0/mIy1Bs2iCFQxtB2emA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I3UJNfbJ93Fl4sk2zrwV/Ea7LcvjrKTrS71EqzjYZ3zG1spYrMPaKM0SnU/e
zw3uVgLE9ONXGUqZ/vYLJF8RbzKV+rPUmmV5/yl5k5JiGP1rlsWbk8FDW1T4
Ky/6jdfQ1ynyD+iksNKq6z4Q48x8Zdolk1a/AGUKioV4NutcR94=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NQZKSnZcXKBU/KJwg8U1cRXmF41G7KWV3C4nmkiz2kj1j8sYxORMOAxD0sfr
NYkwx37C9IRi03oXsKd7O58nDeDI/toAy93+sL1iLH0YaSyOxlqCCSurYI9Y
1c+JhwZTyUZA1vTgpGhp7fkNcP7xv/RiylyLDq3pVOoFj50TtCkefzbwuJJE
wDOyo9Je/Z1FFYZFXm3unTX8O7PGhTp+5N6+NBfN0NcWF+CqLBWU/Bz+eg7r
QAr0PGGGnFB6RBI0UQLlyR3xopJYFAlkH8H+LAiaYFimresmFccp52GsHK9S
MOfLd6CsIvXdjyTuhZ99v2nBCiXEo0ylgfZ68uUJQG7zus0uriW0uq76Zt3W
ItDs1a6llbu8eh0imM/3waDwbJk9yYsZN01ETEoemf556+qOhxaRGJxUIuub
Ko91gwk76PJRlClqc1WSem+OYg2XPD9XcHEq45Q6OBnF2bhftldq6ABygsSV
1CrurXDBN0LayYm52UXfhBCAkJMc0JOB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ExjuxOX+0/9wJJG6zCCY5mXVKMKaoqmbIYqYtBApheNkAtrZwf7UGSvcbhfI
HXpBauLpLbFHFtl+fe+GWe/sCSYugLBRXm1xMnXSSg8AIUE6rGPmKF1ZI98c
x3sAUvYRV/6n7ZTEhMm5G7uMwQhwOU++iWZKd8yzAq+KWOU6xCk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bWdqhPJiWIFCVw0m+7zkqgbs+W1YwP31etta2Ui1qCYmx4M/PjvAeRtfgxZY
XFi4u44TNP0qR3EJPT+RcFH4KAbPFTqgurzYIky21y3yofa1Q/8IVSulDsy6
gF4BJEwrS63JhbjlCwmcOZX/RWZce0CxQwxB1unGYCy/Ep1kQwI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10608)
`pragma protect data_block
ZnfduJCIxL0ZDXLPPzC9Sf/xvizGpyWj+zaLkuH/aKJIsBn73yf25wWedT51
OeSamTmmI4dPc5diJtr6lhENE/KVMJsHY6dBZfpacrZO9RLXERsNsDRQm77D
7RzyAz1FcakLnOg4W44Eab/GH0Wnb+CKTq2BONlyr4R9g1GU5afgTQ+A2ZoI
/nFs1diLB+gFinuwP2Gd0h0AitseyW/xEB449ThWKAEOXlsScVvftxaBVixk
6/JNJWU5dxSK/FQqfczoIVdkrCAklW4KyfePrfrNyTZWyJ0MaC83wfxtNsWj
01lXmkYuzcogsRaMKLXW3BsN2FbYS36pNm7FFUaFWeYP1SV6bJNQaSw24Z+V
FbTBJJdNxc3bUaTlyxwwXdA+F0q6/l6nB+YaeEH7dtJEmVqwU8hfUJ5XHbsM
exbQ9DvzjFAciWqUz52ylVNOXvV0fDsO5CBTlUtYZd/ZJjt26oGjpaIMykZ3
waktrszei52BonJUVJqc5f2Bub3CJsjcvm1e6JXL3FCEpGTkBfDsyFsRHVms
AIsmwVsaWRL4dJfbIo3/x4WhgHRgjTaQ5f4LXHZRCdgGqwalCIyzziB4qNS2
ef+FRcOWCsezbyH0SvR8Z2eA9hezrgKPeaa5ZykY/Jzii9qIUOEZ1+wMwUIT
77UgTgBNamzaEcuD2+FCmQrQJKvfO6JNyP7zEhestjawTFdV2gYkqOE/A5Ro
ueYdd1b1VKRJwJQvbdhuB7ju09F28JQQjqOBN5slCgkKPmHzWqT1V7HW/zBR
KXJDxIxvlq0IKG0mEhOk7in3x3lectIhb0NoTIXZZhqRZZtumrxi1Cvx4gZt
x3/p+J6W+V+wlsvsJu7ivdPANx8T/WJNJhmiVw2kUg2EnVyPkmZwFu3y9SDx
Z+0ZIXXQE4a485HFRypmsx4NlGTDLtqBCrcMyRhfDVRyWEFS4H7Wa/jV7uoD
gg051+bILYAmnY9oemN6ZRGSfxVaEYR5zvnZ5zFID8SqSE7MSsm3IBX5Uo6u
Nw+pZ56+depDJ4XGL0t9QUeUaNRf3jtoW/BsDpAFOaOb9vkXmNYr9eU6QM9C
NQsU+hWUdPx+VJ/NvNAOsMvl6fCpZ47NEmFDuFzVC3ly3+LCJv06xSQQDga5
kyFFevj6qaJmF+Oi82EgZ3pLKMgnhlcb56vSqZ2XzjldCUpjvMfKtfOXUBAO
hjeoR5bvFH5BYZoBvhWCYNCLBIW0oHBKLl3Bg7Mc+lJ5PzbdU/0l1u4fR2y1
NOnYAza8enn0kTw572+GCOwFJ5SN6NmXZqaf7aHCLFD1NYYj/q1EcLtkYuiu
MZANOvpNGAqBBVUADf0pVpqgRGJZb8dtGF+BSOecusz3GFwbxLepw72EOYFO
f1aMDXuCQEfD4e2p0H2UyGVNHoPopgbifneEv/Kce9UbSKTWss2y2n+mGNRi
yzE1mNExCE7g+UhGjB9OOz3P0UNVXxGputnN31gBBS5Uh1NQ4nYViTyX3BIy
bSbo+0fJjt9fPG7WZBIN3iqpdKLsZpGpQ+6umiKwuujS6ShjS2YTcQk9WPAB
xd1rLTVtwvDV6iQdwMvZztH+3v942P0o3Wi2L4lVfCwG3i41Ak35Sh268hdB
j3h/rsxC7vns+sSrch4CpLmMJQDLnXsycgm+Rcg76TT9ymHH0pLQ4+XEihZj
HL9r9e5uhCipR+XUPMYUGor/3GhE6VYhE+gYWe5INxN4zU35ZAV92Pr/hZKR
L0bHYR9nPEdTpsgNT6KXhHzoahIYPzsO+RwBFdRushEbgeZD4Fvu9SSGY293
YA9QLy0Afd4uJkd9iV/Now/xM+SIbNNu80yFFMNTSmf4M/+yYePvgC3ePQs4
JHYHQa0sdkhyRBwhU98UDDTfZp99bA4teyzfSsdv8bqFIvik5b1pKkXIApYW
Vl8FFQ9syzexgKEzv4KzG5evvuxMwJa84MSDSHIrVA8v2v6uYFJE3laYyOuT
PLpWefHsC5npPUchS8ZaGRfKZMb4m2zYvpsHez2TADQjqEOU8QTRsKaG2NVR
P5YqUIa1Z9wi6Hu6bz3ttY/t7HJUJc98rrjB83avSsvK31KRNm4GdIyRCPyy
Vlm1H+a0rwx1xycKpn3xZnhz1oK7kE7mSduwzQ2Z8IxmHxQf6ViDmXKsaa1i
P/+HC9UrCc2FVJk2oTRREsQSRl+EZOHBoM+C4HtDvbEtpKEYm3qzcIfwpiLE
IJejxdYhIa6i9lEghF/MBkfg9cPojqMro6sDLfgUQBt9Z8qnRYgRG+CltZJ0
sxgYOSxaOY83jXI/TkqIPsQu46Y0IAKGOBcJhKbp4Hfahk+kR5txdxsgy7pv
eVvpAmi2yTLIEoc//tKadyJhYU93hkjtx1bq7uNyG/gM/y+UkTlnBLdlhBEJ
9nk35DfKy5LAPfikeDcN5Rbrchu4/8D3clMM5QHC5o1B9eGS6NievoDeJ7va
3INmQ+delAN2oE+VxjpLbvKGmZKiExj5IQUL4PMpPlx29ARg6o2bzW2597Wr
bAUY+feG079EDLngUeWEcza+bTEsuTHEA7p8in8qeUgYJg0eW3/hsW1af/R5
dCTsuSuOdtq7Vqqu+jGZGOYszZkkHdpuYvLOuy8IP3sJNb+quWW8eoEst7R6
v/Ih8VujAaFMMMcLqKbNBPWIgCSJM5IxDkBQgW0HNRFzX4aOkQ8E9lxOegCk
uSbOWMOFoKc0laonVKYZqG8r1UtvNpgAQrKFDYnbR+/yKpWXHOs88uO4I/8w
AvRQ56FTImatztHEkO3j9p7Ppy8Fa4f4NJZnnxuIP4bQtM7dkqcN17w+zwQo
PQGGqYR1GO1GXS0CgmAVWyrgYqE3e03Us6xhggjwjTaDl8dRN6IlxuN9BhLe
TdvyH7xbEYyrL8qhpRsfrdsf6v9V0Js+nI5DbRTmJhnRQijPekFzssp2AS58
Ol7AyxB7EdDEzk3qCRTwnZ5yOPZ0AnIQ+yIT/sdcFq2idxcVczdOHdrmdTwH
LW8vyKUB7YpSsouomAkCtcm3wMmfrthikd2NhcSAFQd4rqP8UpL9VzopPrKX
exKy+cAbuwErUE0XmFf/Y4zoYGt6NrI9htPymmB1N63tITgEe6dwPd1U9LNS
nsBCwArbyis1BV7LsfMI0BQDLEnNFavdiW/EkWVYDSjWkGReB+bYb71g5xVM
uAsGWq9ItipdG/03rx3belBKytLDLRsMeYJFpBIlXkk27Vsn8VrcPJLHqwbm
2oajtgkJfda1AohaVX3wgw9gPA4H5WMJ7+YkjlJ0/+1HoL1TUseBiQ0WNDJU
8iBfU/BuKYx1ClUME0l1F2IdkU0vu3pmETcujvZcITmD6ktCsxovn5Lw/uYr
VwXM5u7OjDb01XBIbdwnPb6FuVwJSp8XceSTkGbUH8VroxRNB8+/srhIfhwx
htgHZerwZRSsJyBIHI4fmK2jg3SqRjNSJKquBtqHkW2SHRLvpcFkSBknHp8M
dZmWyJwKMW3U9RmrkFIxk5cjrTBPPLl8RsGHFRY0q8fqCL06G1/TsVGo+laj
y5YXb0FYdLpkbTWIgXQ2Zq/G+vVucuipdk1ZBYs/GBpXquVoy4O13k0wd7kj
vpS8SpDIV1t25knfad3OyYRJQaRIlPH5o/U/Y/joqSfc6NgLiRoYu2SJW1F1
jJAi13x1gcrH92n1pHKqA+jsTV84IjMR5D9B3IMEOrp6VeRJy5QOev7YuVx4
RWGCuUto8aJ9xZ8XYnOK9unpBoSNe6/UCY8hQkdTNzjOWOEN53GBBFs7TQkd
mGx5jsLKyjfTx5D3xE/jhbGDSiLq4Ka7ypSbBhp5SYwBotsFeIh5T5HDzP6D
i2rX2R9ZbfdbNXyX4FVz+biTI4ZxQFBWuVVaruoZ2zjM42pu8ewvGstTITmT
0KFi2u+ErTXpViaNA+AKx0kjawAr/kLwRRfXEzBaZR5NrlPwuHjQEA6x+waQ
LgrBMmLtIxPZ0MGcGNOjngwv0dEsuuCLi+cjJ4KWwQXdyZUKyLCCIW0woGAc
NtUY2zjBQIkZsyCabN2/b5Q7al+C5fH1z/x0bpQ42edK2t3NRde2/C3wcId3
HGnlgP+In+kErIjqw/ty79u+56z+whC0Ob0mkldwMv/7YVhxtpeDsUgZ9yAv
c8nMj0VTAxxxEAS6OYNJvIoUXg0hK3xBaWnPYalLqRruzUrEfoULHuieaC7x
ADIOMa8jFy+euv2fXpbjvsWMOCJ2d0pBGDNVC2O+HfeXIuN8M9pp2XldwiSg
j/v2IDZWFrfBo4ThAguH6B7PGNC7RKuSZ3cvAlDfpWaAqcfBb9R1YSPJbl61
CHISJXgtTT+vliLgZkuDxwQvmLp8n/WeKF714noxkvqNdUo583H61tSQQZPO
YTRXoxtiOEn0NG4WxzJCPJj73V3cqmCO5X7p/fgsrMLnav5EbrG/5m2R8ePQ
b4fQoBH5Ffj9AAGOrckoeNpTN69hEQcEQ1svJJ0pBIr/IM/2UGnvp28DVuWd
YHE7e6bh+Bf4GH1YEXvmrJ7wOdDYRsh3/PuP56qqCt9c3bPMaxPxS8ZLqSIa
H78IXbMN13o3mSvPkxqre6K+CKkK0p2fs4WGe++b/iaEFCg4YEnU9+AosI1j
5x1jRbwvPRIgb+4N404RQwjupIO6rHdbtwgee8iWRTjakl69nJWk5XD9h6oy
OrGmq5sdQpYc+cMX50xp1F1szAbvxqVK/BXjtv8zUdnHoS5AO2mV7ZWkdAcO
1K4Tscs8D/he/yoCuszovjUSVgbekT6F3Esu/ZsCKlKNk+Ugi4A+vB3NKx1I
P5KQG2lAg6SKg+lgVTeOUv7f09eQvNPsb81942WwHVYf++DHbJIyzcyktMkB
qC3kZ9I37jFrt1zeBBK3RFANRs84bot00YinNw422SQQGun8HvJwxJgfTOY+
qYx+DRRh3SOTX9cZJm+Gk/F1KS+NKIiUBmmojIf8C26ENh904bAUhT5rxunw
AAAJuhChtFF4Hqgka08lt8gRgxtn8UqeRmmbOUo7Plz3f3yBz7sAxV9ZJEHP
li49qqS60o18VK5XFRVfh1u18CpasQ15B6XKuvs/vcvTPGE5bebM5jl72bZY
X51MrlURhzIDc5GfHEWJCK6y5XHicrO+lBIBHxhbof4WbU5XOF5yqiYla3Vo
d+RdFmnEYeTjzf4brOzo0MTQau3Km7mSGcdf02PrYDWgANgNzmoe1ayYTvL4
h12V0MatKdKPdqLmAKo4frrjsYJ2yjJcrG1cAEv2GVhXx4tB4Gvqv/9hovM5
xBm/NgA3khq/5VrmyATYHkjluFEisnt6+E0NYM6SiQEdgGG6CpAwNydZ0iU1
qH+0UayTBV3pFqBx1WNvNMwsr2l/VVgR9mVHpsR5MbEFGk3ZjPAmiTLD2kmy
Smy7Wbi1q1pVgd7a3UoKSAknyJXw25OEkzWHsu8RtA3lBZVFtpdTOxwtN1QN
AEivVR1BPrfnUxms1Y0L4JVSr3M5DkhXGkKTtBydte3FlvwjBKzqnrN/2VLT
Cx3BuMS73o/OmEHC735ZM8rSEYDzqIpxa6pbW+SnnzjwbtPDC4GkOj1jZXWZ
vPG6ZsHJUNC3kxb24r3fTsMe/9HWXsqOTIRKAZCGflTd8yPEDuUl9F3Vfcjj
C3Yq91SRPOlyPumpYnpgGFkAiYEijIEH0/hYk4YYgAykRIm9UjzN3VvW5VlQ
0iru3k9Yz/JG7rOfKi0on5KlnBtzx0+ki+9HJCQUyjSXJ9Fu5jXXxFnkeU9i
THZJERkWMBdbBjDgSfBQMdnpiTW0b+J9k5+HmGxk3H1jSHupndyHqQpbTFri
Nw5lzv3tC5TTIbX3hPGbFx13/lOV1p3O9J0TA8TUCjL7vJkk0Aw+nxraG3LV
UsStLd8NYIW9oX0zdlN2WSiuSCGUqKuIfDcO8a/sdddqby5CoBS5BXHU4eqi
k4LEtI1CjbjoEfuo/r4zB8crRhUK0efzwvXvLSDSm2zNbmoHp6cOrhCCc1HR
ZFy4akzmHD36ZUWi+14ycbIOdpIalC98EKNX3eto23yuLAdLY/ETAtUzfBkW
zTCI18bEtxDYvsSsw7JcwTAZrS304l/G+HCn2+k9ZixN836BU7HziDce7kBH
KXWKUS53e4Ub0pkcsCEjiC5LeqfbRNdlbz0rWDLhE8zNSjnkcz5kIBLeH+Su
GHKaHNueS6ZgPUwKKN1HKpUwTfdQC+3AztjBVjL4AAvIwnx4LgZjKCKg5dQF
jzucPWhR+4i+Ir58HFxb0xBT5v/lPAhMbrjEc3fSkyE4s+koVbBraeh45Vcz
1TWm6pmecnOgPKGxR4WzeqJLclX9+h5Vo/XQPHr3r9tLiIfrV8i/vnhX9YZ7
W19p2jWbwmIE7hRvXeH9XmwVYgG0O5dz2Dab6t6mD7ztBrT011AS3SOakkB8
b/rH5xOzin/7s7oU4sOB5SNBs40obRB9yVjRkRRveYDK9EmTMnGy24xPSjKD
gfUL6nalJgrjOeapw1dlGz9NQTXlIgru96AShAVVNXg8SnFG1y7hpT5/aYYh
V7u/cIOgD3KY/Bq81TcXj74F3IbjXzCu4L6F8MV4IYpGrUafC+ux8YA9d97r
RgJUtwrA9wY4+MQIWfkIwN09khYeeTJmOuvXtgf99yGAHTnUKUppxTIkJFqC
RbiHqWZO9BwAoSPkvfXDw3JEfWyrFzRcTOcI2ijfQSyGvFozLZD0GbtrYivP
jQzFKqTgrYVB1xbiCPqn1rR2EN5erKmX+MMxtOdYLUPpNxuBbrkVCZmCo2su
5fTNVPP7rmPAV22tbfjQJcpaV2S5ehqBm2nNm49lW55+KCA3WPrYm8a6BqHv
OLmnZyde3RXiWvQOJHcPfIczjMVmqd0OpdxUpzo9Wy0mSkrRW2ByF7joer5J
9Ngg4pawBgkhGFJL//5Z/PooGLJnRIxZGICtH0lycbqS6X8tjCvFXp2gHU3n
IElk53FzqbAvDZQRKSD1FGZUqj8CHPxzK/CcfU07Ij5aBvQktPqNmzU0iezN
NHInt/q4J3YqflW9Z5R3QkfhrjZ09+D/V0feET9q2N30SAJjP2MLVLv7YGq5
NzAjZ26T2zo7hMCS8hvEBHfhdOD8Xv9/L9eqXyqSi5fUBAukd/PEN05q87oI
iBwB2B1CVuPSLwJOhOkE9h8OQRrt9QJynHrzDlVAJh0tjybXAjbaCwsJZVVP
RAQjutEl2KMRLQcMteiuxsr8eQ7dsy8WqbCBMbSDXMmvRAcwheWSJg7yZmy0
WZBmLEXN0Mg1ERLQC8jf88ux+ojPq/gaYtcKvXiJPYNlMWVvkqA48cSF64KL
OGUTLy/+TgdBJB5lxBzgZJsAKnz4uZU0iV1VSuZBLXbjhra3EAvttj0eWrD5
4Giojb8olifDV2JbPTYUPlzI1LJsz8xdiBmeU1DbbWY4XzOmvmuegyL8ENjz
NcnQpETkqKeK9j3HOgn9GDY+6kGH+nIQuhaOV2iPv5PB6TQ3IO4bNiIleX3z
8au3+E56IStL484ckd/rs//6TbPolAh/RPNESKSy62K8BTLgMdEBgCJskAGc
55FCZKnYo0wf4HepkYdufimzfZ3LRBYXKA9dcClKBGPgQVaw+4TbJ08uNNub
CDBMTLqEahYHayb4oY6D5TPrK1VUvpqgL3CyqRn6x8c6FSJJDjSSZ0o2J/l1
Fvduqy43M8TE141IwJuVLx519moQdDIi8M3S9CIdnfZGGjMq6uvHYezWWv3c
ezteBeIjCP9+/9slb4BLaGwqdhzLDVR7q+dJe38g4viqVkayodYCyBYaJOma
ewh+bFhZ7AyWcSwtbCzCnK1Hhq/4RTCBK231oSwkjogfbIZWn4wMXAoaYTFJ
9r3Mn+69dTRILsq+2hm136AT+cbVLRq3n1+eYnVEjVjTZq871qBxfZpbGy+0
MEr2jnk/jEQXOlBYd+Z6Z8x37Xa9ymKVUOSn/8XpBQjOr6w6Qr5G9FFP+U4J
3T0HiQcFsMuyODKPqLlL2EIpAdt/FKb/p/N/gHCZE7DdF8mMyPBHV4hZkx53
oNZjKdGewbnDJCj/H0sncpwHomLbTsHkPUbTiB+oB4WAk3zDvp/rGa6SjHzY
C+f2+SGFVHGi2s5jo6LCbld035VOYZplMWtR22WqvwzKMn11LWvrVRl9evBt
So3ua4MEoOCpYEQudHoA3aJbksPDfevvSDva2Fwq5kBsfMzPE2S6HnY9adbm
p0O9Go/kOduABbDY9g5hdzuUuJX7+PoDIyGr6peiaw30Gw+rj+GFTPQ+0NzP
kaqqrtZP31Yx+PPiG7J58TOKE80oy1XFi9nsu4KlpKKjiLfKErMuyVU29xm+
QvLFEtc4l8XJ6dvKeZ3mxRR/Km1bLbbOvDnUx8YvoEomarMBXwgFvmaXDya0
1WdPxmdNEZu2GFsanhFKWzHAaVA14OHTl1nhJCR8+WEksoJ+/JaDTAY6rlSd
Xwc15jWKuemgAX4S1OfRxFc0gidetJ67hj368hatkANiqTbEvIXFzyGB262l
hir3gLdeyaPgkQXziUzIHfEEIhgosYnjA7uitwRTegfj5X8FBYOfCcGeM0KK
7URshXY0sH6tYGCAGF7CuhoMTFbrcgBQPc/jwrzlqscguy1kjNBZ3PKZbQ0B
J3q3gceHHYDFa0/JcqBcmCGNFQMFsM09JzAbPo7P/NxvTv9vcvD48so9zS6c
pQuTaowGcQtgRVMVmKmmBRpoYoTKSWKUJvlxDW8/hgNCt11yEcmzZ1aams4S
r5SddyKvDMywCMbozaTHQ1/M3nrXRt50hR84sMYqNy+zfVvSN9JF0LdDjzqt
KVqtIfTdQfwYkG02NayasGkUnlTrXp1V+jFB4HrObUDfKoJwkuTHuzfoIc1t
ZZCe9Kd+SrUDotVwcb4yjc5pcR3QRBdrC60aA5+FRgAmTnSO7J/u9l4mXk+w
wDX4oMknsIyJYw2Jj6pdcQM0shQjQXvHaf/I4TXWfBl1bd9q7zXM5rxyfuG7
vz9Io4J95/JRleyYyx6dSnKpIySmo3+7xTuod2vAumS5fk+tZszSBK8g/q+u
f3loyrLJ9lIzHtt78hO6Htzx96v6r9zba5FWJgDgBKUMTXmAyRlMk+kSWauX
klgfOD4QovWZpU2tyGBa8VSR+CqX36yWz8fmsuxNwNzTVr1te9JJhC6CEr5o
iye2S2/FZv60r1O8riSbbSfHvRGnG3HMEU2Jg1aLqxrpiQsuCdahF73DHIn0
CCaJJFT1/bkLJTr0eHp/qLt08xUVHUqwl43jtwEIVt/aUOOPpFs2TpX/pUYA
2wy7Q1NSBLDoR6ztDY1Qmi3MftDVo8oI62HbhsUvF2Y+Lm5E/vthy3LIa2pG
9vX//1cdM4uiByZt4lDd02YDuayzuMJY2eWYBZwVa1otpO0gSdOEgfcpKL1A
VCmHHJz+jOPUS6ugCH23MctaNcpO9ajhOF9KnUF2wdgoV9Ex4ni7k6Pzi/Yc
kEsdqMZRjBu9DX2vg/4/DO+ZQKvnu+RkjQ6zD5PBriGSOfC6vSuoV4ucrSd7
REJh8BzAof96Y62vHocHdlfdtzzIWtUYG8JMe/Wif9sZ7cb2MN3DVbys/Yed
6WFXhY98HMaevFu/WKriXRc+jXZFYZvS9XSm4dry+w2GXsK3hcjR6cWEkBIW
rwomSmNfzIa6cgb6gERHZzIdhxM/Jlk60kzZMRtjM/GBAyg2bjekqBBZy0F5
g+VkqwQxngPSIaImwCJfXxLq7yHPloTnTOOSQe28i4KbEcAMmuqxRGAaTf5I
wRf/EJjACMyF8hdebWXstCc7HLgWtY16RDcdsEJ8F9NbY06SunCI/scIzAGB
qd8svAehU7LQ2DNg3gyQZqc07YA9peZftv2+/sEat5seya5i7Nc+/n61yPCW
AZW464e8XDaRqmFqnu2fyIRX528C+38KTd50YnLjEm1NlJEjNy/Tdn9oI4SB
zz423aZhj7pmTn4MiLdiULFYmIVr1xLvYWbmEElBiTeNJAqKtoXyWP47dtdO
pBued+VKf8AxWnqeIggRVFGNiSBeXxsoAw3MqcxJ+jfBmb8f2PKJsxfRxym4
iLkbNHxpwsHttxDtTCkUOpGwDyDryLTn2JYW0DI+EwmcgZX2nAt88P8g48LN
sg4uVOCDxvLkiXQQemJIC+DYc/GM6fXZvq4bm6v6kStsYGstXC3TRQS0z6ei
x6XZH0YHEI0HFu7aDxI8SdzY4t+YilIQ+EfCSSLC2QRjAv78mWGO8uVRv/I1
57+quavyODym6Ed52XMqDxfcUQ82eZ8L9OzlBmAv6eWKitTv7F+4fkK447vC
b2AgnFSr3VfVCsPTyKaizS9v/ztQgYgoaou6lZ3KUQCmmxjVqbXd+jfqJ/mF
R7nq5YrC63QDQVABVpLnGyELMQF2XFuhA4mC/t6mp+2bf444amjY6KCSf99i
R2/16QNPhF1KI4oohLsw4IJvLW+NRoKZ+z/4mTgcp89JE6Q9mzlhtk1WwVah
m1IF//ORZQu+0ks+2yjKBVcw+7xPTqQLB4D2vrtXzKKlD2jUrmbI/E3V2WZ5
+VmllcE5/D5kCgtLVDaq2b3s9MkxRFNJF2TSgs7TqpmUyRQVkCkzM7Ne5mQE
CDqEXrGGSgYkmjX+ZPWcvBsk9Wnu8Jw2hzvHfaFvNrOOuo3FAwN6LgbTt8wh
aaVauAz50szet61BuI7S4nnyDT72czjNNcpH0JyW56XtPhxE8nT3bCbLC4f+
yEYoM1A2ZlV0d169gVzgR+HyU/KpEjQm6LtxM1x1tSqlXAne6dchsDHfcTwm
w1e8PG5dtvlKbqvDnl/I1dHvvwPVHZCemN3ve4T0BHKS5lNBn194J38ptv8p
5FgO238VXTsGOmzK9bT5z5SC2bT1zxPPARpgKd4UkiNiYPTgPwgxu9bQ/MR4
Mdo4T5thwT+0UuAqi0WROIroxaTekkLHzTKN8vb0LAYtt+55peoMSOUjq20a
pceTL4FPJ3Kfs7XRq4j9FhBop6jeQuZUO4EjJsnz8Q3sbe/MQ/d2r3pJAUPd
XhJZM4Vj6AaZsVCNFRc8Su/fDeTvQ7x9zWBJGXy4pVbAwOzztTNMEXzk/+NA
9uleXEhUXuew6OM8vtJzaAfYzeftLKXU9L/suPhO7BpufoH/sbSzlz09XSGl
gTndGX2DXHODBYzNSea9SUtLeCsjNO1uWPVBGUfRvhUdZbF+WBO4Gha65U85
bU6ky/YH9Ov5v0OyT7xCniDgtXXc7wkMWPYG4RzlV09KqijsSBlULp29acxj
a5nWYrt8fVA8ZzYM/Cbp9pB2yNeGn9EBwzhdb63lqX3eJVUZhVlPKrJ267gu
sXWXAc6MVXHFvYpjLmadJl0iSNtb7OHnV504DMUOX0dj/UCd/xcYm9Td4y4/
XUEb5E6VAOh9jtG0Hzv1i7SN6CAfQX70E0JTT8fcwfPD+LicpEuYcWmSeA76
b5w6c+pcDQ+L/SooKmjLUZ5JVGqfaGikzTJnDpymq5HEtf1k9yfX5IIPfTHw
Cpk0APEf3STAEPRcOyb3epBJz9+3YT8myxV9OrUS8SsNMw/STikailKZ0aYS
hXSAgy/WKynAv8YPqK2Gvet7bBG5AxL3J/Nu2hdl736Sf42rt/ddq1H97qJY
RPrZ9dW3peDsj/jucLLxdTM1mFOkxpqeB6y8uL1j0nR6P6/f+tffh/Z9S+uy
ueqNQks68dpCdpa6b6Y9takITbWQMIts7Z0hvSJYbooXDL4wm6NINvQAHXsQ
cMxZPlHs4HtgfzOXPbHt+97Qs3fH2UMmDMRNj/MJtVdC1XmWsy2a2SA6+zT3
y5lrstT2TZAimQRZQiK5XQA9ggecIomqhFvrUbM1P6HUHcUWfpDXrIp+J9dc
ZwqbWGSlENdfZoev0dcnxusElJAgKZisstZFbsRQP4QCU/p1GQOYkFZMeK0e
rX45WY84r8615UYAb/QeLg+AQrUrO1JV3KB8dfQMKPoD0kEAfbVJ5YXJ0NYB
7iF5CnjJGS8ixzo2nn1K0k9eY7jlEt0t0RuhqmaXsqTjwLMbm0dtf+mGmFH4
xjogvDggJ8cIZRNMYGc03ynAhsILBrDDQ3g3aCSlNcuFfJtnW7kGfgc7nDJ2
ysJvqx8we3eh62sQJI+YeJCdywsdzvEJGj0d1XenXimo7xFxWq42Y4HtOiZ2
VUpeHnCTCXJT92/1bXoB4kU5VY9C/oebL08JhDLS0tyzASU2jcZPtyqUM/pr
VwDocVeFiUtoKzrqRqef7DhQ4/l6fsgk+574Hs//UBDav9tsWJYJxRM0Zy/U
zVhSlBrXYiPJ9+LpXS2zVt/KzrZkjnGomgoPM/JjzsFHOgrtC7f0dt592wCz
SOkgSBA85g5TaYX1VWynKWexaHBs9BmunWRxONn5JoC5L0jX/tGS09pUHfVw
qtS1CzeemSQM4aiIfBfcr50qayZFs1z3v1tyBNjrBQvX8E5at3O7uorvYkgU
1pWyVw1mNG9yozUq4G+9S1XRhdao02d0iY+xHLCYGXZXdw6CH2gIrxmimDAv
6UUJOQJcqJIvgGMd9AX17e2G+25ezBbL6DKKOMWDLOSB7Z9tkFrUFPcxUCm2
l8NQArV+Yn6bm0tjG0Dcd5wBV1iv4t976C5J1ORVlNMlAHG9DJOXa0eHXg1b
Uw5SAm16iHjCXJ0sSlCmIt1H1YboDBjbI7jeB9A35kCKTKC0LqmfOpizbyFz
uVfG7g5hkpc2GxbobX84nPLHgnOoNJZwhWx1DO5EpwnD0VkQyoB5D+KIn445
bWUc/xUUUG1mEJw8vQieUaJBY1bqfnovkJ39ZAHfKlbInfUeILylD5YBHrPs
77J/sCQLVy+vuku29ihSLcOqLW8CjzQiK+TQoVUUX9bq7A9pd2K7cNV7H4aQ
/4IpeZdIyU0AUd5U42Kt5pL77/6GD7cF8TXbfaihO1SQmINCjDawZHv9siwQ
Alv58L5wr3TxCnjOr/iRkVd2Z7O+hFdcS1mQeAIpxl/BmKPD9KUdWodngWkM
x/GLWXJRFXD6RMcXfh16pDCvNepLUuYJ7uTtwv57cg1z+b7e4aNaogq9t7Z8
Nh74jBsLLUXWpCIhmPG6Ddw7gSMgueBArX8FODzum7ltREZr3zTyi8R6dmte
2sGTrr1zv9bGDAHfbkGOEUwn+ISFl8ruwn/4bgae0b5qSmXokBm+FOhn0T80
TxSOMyab+CvXlh/vjdEax05ltU7NXXGM6G6CAHmLg8ngtdz/NslaZuy8rBtl
4oy9zLfKZtio5b7W+AzwQwtRj4ZFQCrDo87k8rpanSMsgqli3N6wK5tRbUSy
A+UMCJIGMANM6Rk7aIQRFn70m5SRzI57LhzV3PdD9XgTPnDanNES9fsgmEw6
j2YwYTHl8t6dWpAP3AVvAmaXnPE4CPKCWc79A9dRQ3X/Kgj6JDveVmXJOQ2q
6fVbsU9YM9HjYTDO09VK5UNGLMyeo1Sp/mPoHgPeZhi5KaXkPLxA2NBKwG+b
xjkOGuVh9TJHI2nb6w2sc35OF3y/iC56NpA7N2I3H7u9Oou2I5DgzWAiVDI9
xoZmpi1980K6xmV07DUkyOnYBO3K425JIHpx931d46nVpX9eg7UnvQ2ngVaM
+XkxuiN8qrF/mCpBFSLKaYiz66WEpbu4xW8+0ojn2JY+k4Bqj1SG5tpggwK6
nM4qd/Djod0lnVKPNie+egMbLxuNSbWGpwkMvriFuJAY+c0lVRcGhZD5xrt0
3/hQS+KAl4rjCfMyOAELdTLFV9YCG5WEL57RJcLCV8rHJdd1n1TpAurep2ti
8zr7gVwgZG/1FbSCtUesTgnOJ3MYi9QrVzqoO8jwBlkhpl5A3dIQVs56PjJY
t79HF9DjTs0P5e3s3GH9mWKwlxg32aBTnFe225gebL/4nwaq3ad+njKOm13R
9aMPpi+aCgzNixvxFDHvJ9UpC7154VDSq0TEnKI4hwUCZaC4AnGK5LtxodmF
EAb074PEWIsAlxKcYIXP8mRsSsmYDRm98z8sNXZptKpMjw0m2R4vhNXv34/4
EBZCkjYjEfwk/PJaPOTf84n/S7ME1mM5kWCxNHq6DkkB6DJa0gyQsfxj9sIP
S1TIK9cjOfo/FrQS0wVuf40hhrMdNJgym59S/SQYxM/J

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eq2YHYVWl3pPz/pBZaSGrYX+Kjrwz/H3WkG8XxA4zM64BMAiMA/fpRUnUf1QZZRa0IUqm6sFVVYanIE6w9GZSPrYuVOYc+xM1ddiaF625rACJOCu9u9zC9RBfrXmdl/FDD8DytmCUFg5ATNi0MW20jO/MpJ2gSw7/fiCerGoV9mWLCHu4srqIzocwfPK0wqaZLOa7AOAELTjc+7IxKNB+bgz653YB4N9vjy5s5ogrJHbiqiJMXDKmzpO7PWnU97p590jnN5OwoXG6PFBuaq0/FHmvFkUFBx4H2nYdfzjWyY8z8ysOmbSNR9AMLTwgNEQYKxyhJgI9LrNSf/nRPsgjX32wfUpmUYdnECqao+H/raRVKITv9EOGs3HkSkW3N6gxIemG2ta8hAqgbg+NdGWBCAg7FIApnnIRl5nOJU9xudVPdJgHe/RpppvJ0I9GV4MoV/4VGSOUKdtnLAjxdjAU4IdSDg1UBaj6QkzuaAKEsKpU1RY4eIs7x+xaexfX1pNDhXJD2B4TYjjEi/pACRhIw3/KOrD4rTtuso/3HD2l1RadQgVq8GzYKK7S1EwEaOC88ipEVzg5Xa//z0jdqzyj5kXm7x58wkbM1iFfo5AnC3bel2qdMaLs1TyhS3bbgdouCSXWO5nS8BOvv0fg4TQWhJ0/nV7zM87xfzt+cXAEbW+DjUYxIl/Jabbd2s7gZ28/wnuL+z7izOykilJFtwD8b7qysLmVPt97irwvlwIcJaK+5GEHFbRmMsDq3MQocfE10+gDr+db7zMTfi0Oqs1Fy4"
`endif