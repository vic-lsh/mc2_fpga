// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eY+d6b6N2/tQnyFYcvYSdoPw8ikcepO1agWymOEPOEmcSHE5LeLvXsrMynY3
B48yU/Ga4wpv2oLQDMaKiYt5IjJ6CgB4docyLumyMK0nMH7YSLdnVae/n/ah
PKBVfmH515OwClLNiT5I86B47hVE/dq9WCP0K9MQDWDRlahok3KQWyY8yPYS
O+iqdoOVJi4Kz1r2ZWcWLeApVaGeLGeaY1wtCLwrswdxKFypluByGkWIlYNy
7uh0RLLt/Rvb4Kt4EZ4+/aaAZKApy8HTHXDtPYhxcEP5rDa70McP3U+siFxe
uhnND5tUC6oS5pditMVB3MhtqoDHNcVkb4qfLD3p4A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H2Gw+BvqstXvgT8h76FCLHFyBQbnukRMAK0L6X/w+skP/ehkNcPl/qN5Cf53
nARLAjqMe7CDmQZ4ktipt2GuaOQI1NGnqw6bMv21+XFrxuxAafpy3UHG+9od
jZ/0mOhlnRsNMHX4058kr/kVaxFa/LHWypspZ1f0de6nmQeLd5RpET3j8Spp
lETSzlWFFkh87C40mF2UVIIlI77SSnBGyV5I7FRc19MBuTdn1DF445LTx6K9
jzNtI+C7QZzG80ExtT49SEUEX77s26Pp1P0ZfPOpaIRrhKuVUiHIdyKcFmAw
cSQPCgC09K3j8AHjyd1OpSPVzjESwwWcSLoA13wZ7w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bGln8/xuPALgG8/qqDgtpaixu9EX9TcQ+mV5z/ZqPD7CK2X+6H3nuw0lE+XY
F9FH+ZMWdI6jS5aTXehHIgl1wZqju7UC7BrDzTEXZGs9g7eiOPs4gU/tiDgD
CfhByEZg9IQK1m0yWSTsu0UBMARuLWOby9T0JTTVloYoNK4PUcHZLDObBuBw
fKuMZ5MgUw4qyZ9DLbhNqZYx7KI8jbU9M4FUEhYn0/qKyNNBfXc6QlYa5FWn
uthSCGGJz+EG+qsDnTVdxwymR/7BwQDDbPmcmpSJeWb/Y1fxwNKlz2UGjzc4
2HVAFs5VvwIR/R5a8Y9I5P4LPDaQGY8lVwAr0jrXFQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NR1DnRAHGKpyADal6TIYiZpn1hUtmf5jbaVom/G0BXA8+TbHUeqGfA+0clid
K+eusI01AhldE0TaJze8wRzcH+Utp4VGai511bnEbgEUeMMSzR5H3+IPFEHu
Tf1k1jYqu11bqAc6WJHLGmL3wcwqHS3QdczOlrKpCnGaLOyILaKzjbFw9PkR
lG0PTvwF2L3E3bhkYwAqxjV3DX7rzdtXlwBeDriPL1fii4/bxu1/vsylwxar
nL6TSPrgz8ZIDab7p3bPcvzIxLPqL2w6d1bTq2oVyjM0INV8Pq+LBUJ1EBFp
A9x9uwm0vQryDwGM65V4G8yhOOsJkBhb8Bw+PBKl4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S+E97xq+fiFShz7qAlxiLdKA4wkIGE+xmrzw9WtrfwsUj11he7AMtVO8sIkv
Nxx0jv1R1Tat+BIr8/BS9xyUkoqErSEjbQUegC1STxJt+k0c072cUwwYbqa6
h/ZrYyHTydBZfgWDkw2a3UbS3ZzQMhfRk1Yuu9fmaNRUHT5OeQQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RZ7TeN54YZ4v9QMCJqeNFuz9ZzPze/ldjeBubP+zK5sD+8s6B3Lg3YAL5BRP
06/LPr49Owt+ekjuYRs/X4y6ooV/0GGzV7hWLMpQe8NzEDaldrY1XSdq1DWw
AMHrEoVIafcFhGR7J8aw0UxJeneEwLZbB/YKVjR9rhcLsi5SKqye9raMNyJ6
s+jN60EucY0l//PvsKhXzsGfSENjmaFfqugcVQSn7LXuVDM++0oqn0aG3Gwb
WRvFEEd+YeziGXTiuXzCG5zwbTvYfJzU2f75utktlUBEdmMxI0QzFkc+dH0L
lXQO7YjOKXmv0D1uJ8luIBMDODOYQ0AvWM5cKjyFFmvm+6RWaMNoMrF9s2AW
I7y6HCwCy/Zv7tE9/kjeuW/1lh35YljCcgkKnMiaxE3muY8l5ASN+8zGZmn7
il1d9aIf4bUknh3Q45Xvi6kqXf5TFnUxCIS8hIyd1FSXoZTlR4JzbWK7K9Dm
5y/FGLmM+KslSTc8/VNEExgN+JtJrylP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qtr9lKbGgPhG3O1zz5hiIFy/9rK0mDwtqPhfnI9XPikM8VRAF4HvlyKAfeUu
OvQD4ZSngt4TKEqPhP1WKM1Y0daeHIOOtfLZ9hue7jX3yOQcBXVLxg2kWlvx
4kSCih462Rb1PGt2TBGT3oF5QRqwfBRkKrKixNS6l8N7BZi4j1A=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oYI5zPdaD21sFIVQq9H0eE4898GcJwm/zc4O5Q+lmh9bdF22iHQnZb+3CWsj
Za5svwGTms7rC1u3d3SqV678bFxKNktZHK5DHB+/EpXidAKuVyYRuXC9HmeV
hSuCc8OlScKGMk6Pn6BFQvKbqzFwipKJl6ubhfuHi5UlqPHWzeE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8976)
`pragma protect data_block
Cf6uejXvEa0qXRm7XBjckwVYSOYSHG+sianF3JEWUqY75SI/+9FWdz2lGQFA
yt+UqaUevMx9nnDKtHFMwTKcubNyo5JUoRhg5irVr+EwrCqj+08+LesmuIVa
TgfOLlb5YnHvdct/olyq01sNEHvLS9a7OMJS3VpCnKXSFjFCynq7/4uE5sX4
LhEhwdiNoYFVG5n4azHLE46iSXm6PiroEF1XNO63QD/xdCf0bXPjOUT9PSis
E/6irGodu0PX1QMBzZYHu2GlMtCk/qJYMaQ5KG/Mzh5dnav2g3RvOYJ3wpqI
koLJ4/g/KGZGxlmiEzCloQb2RaIFnaMnIc7p+f6890exYE9za/nDPrP04bsn
LnEO7wlirVd1NwuUyVW9KbPXjRgUr0lFYHGclk8NXuDSKa5cd9VEoMIndkcf
m+M72+WawxsFkSCVEURwMp52F0gCMGEs0kYhJ+FgHhvpnB/V7aXlqEx/QDsb
nJ9Hskn7RzbQFjEWOOYf6McCKYGPzTnbGdrPUAk9GgeMsg+ygaCSwzNiAzyX
YBWOzo++tW1iOT2Ku40kNFc4IdcgFyyM8ZKrCAlBugtBMY6+1QiteW28+ApQ
pffHGlPqR9yTsT/sFtNHWLRfC67GKB41CGJUv4/amsxHjoBSnAG8i5h7Vbi6
76Tseu07OXsMyLhuC/hXqXKjH/t7J04F0Ph+hwgfLHjPVs1QUAOgm7bK5s7i
nhpRGXKF7/So7uSwdq/p0QZcDRuQ8bzJsxxlrGda53xP+qtz7scEEpiHzWaC
tJWaeXV/lGLWRecmW7BnavjxkEVfeULlsK8avW2RkcI1xhlDgWVmwR2Vm0Nq
LAHrKECAxslWRO2y7290yaS3wzaxjgZGPpT48V9oJ8MJKIdM8v4XXF6zqCWF
1pHJR1BzrtnRH30GNP9eaR/eo7PBjILUg5PRlL1yafCNA7/Hl7YszdjRctYx
CEZYWD6s6p3kqCAkwXEGZFLf+Dl3XqKlZV9wCUpBoZC1Hge8XJUIANVxKigl
lImY6rUOHsWLY6ULnmRPB+h51iU6sPktiKZOobZESA92djufXYO7IaL+OQar
aq1LyV+zoZ5Og/B8seha9eQ8/R1nnRHQp8t3ahAtWSZddglki65Bua7+LSzg
tRuX5iL7yrERN4Ewsk83wyiEI5iexoOB4sDv6BM6OxdEJOOzKARB8Mf12cY8
Xs/dhOfe8aKOv6pA3kY5OQ50Vuvk2QbnSHez/5Sjl9sWRbCUXA0Kz4f7od4A
iH++kdd8UJG9J4MQYKzvSl+1Ruxqc+AkkmJb6lI8e0SDsEVVy46m0iJPCk46
4dTiKKSeOT6T7kqwnfZEFM/mPmjwNEYZLgOn9SrN7vpEu1g0FtHvLoTYVmz9
edjHBS4jrmDGzfObCpx2SkxQmZT/EmTQUAezEcL7jv/uWgCSPQcWQF79kKrs
hwT513WueeWWFHR8gyjLln6yMu1SOF0PDM3F+Nuizix2RzrLV7Ec+BkBGa5d
guYCaqLpITPCimN5qOM8imTK+t1VmtmyqEtw0cTQ2jdB4MSqbt2tBXe/q6pG
g6qA7MbnnLs1QyuLVgIsQgTQzWY4a3KYPXHBQLRtgjnW7N2z6hLHHN0vCO0l
2ZT0CS8wCvPoiCuWvDveY3SflD6nFn0ntWMQ13xuuqklx/1c5NQeaXZHfaMg
57GFX2dtzNvEiLMrYcYq1/2jx2GYN+8/witbjVmLbfxtJ4vuMUZvYxuPBba4
n7TsDBQKgG9OfFv3Bkl9FBvV3k1YVU4wB7ZyzrxhEclwUAeO8tKdPkd3W5iZ
xScfg5tlatTm2766Uusu9NcucE/PSRUvm6KQjRIWxg+iHG7xTowL+mzC5cSA
WU6tnkpN+u/NK7RyYMDNX1RHs6GY4jS4i/7yL0o0Al1epwnWihBm0UKo7qz1
fKjcpcPJURsZ7sMSqThmUWMh6fWwAGAxHB+Bk9QfXfh6XqX0Lk4P5/uDziEQ
P7amroCNoAIJXtDa/lCBKagL+hq+el5dM3B3XpvM8I3EIrz3kVF2F2OLVBoL
IkP1tsRHQL2D1DMpe9gB9zJ2RNEhB/3x1mOCfc8xGUs1/lFNegHV2qusci83
/y9GohcGI3pXUVz2uGCrHkeX2IM8nAriABz3yTDc73OmK6mpJAsRtON/GtSE
D5prkIU1rrF9huTPfE9XMe7ME7aYa+/jnk04Uz4T5HN9D5bLYdilBYLlKvnn
9ZhSOqbuQ95cCOC1GcT6ojiYp8FW5jdFmYk12yNp8xm8vjy2k7Zt5gkzQpYW
5v6z4X92kIcbXS9+IS3JtKh4jRawkIZDj6OQX5WD5Qe6kqt1itEu3ePAtViD
jxzPgaA1pbRuc66Wf1lp6wsmMb1xJa/cDUSgejqb1euVA9wSY7w93h6dmeKx
fSpktzoOzuYw/LjsRDANrxsoKtsWHtZABO1MH72zpHxz/6KmUp46hlbwFqTS
vDmaoP4dNO1BufGXA4DBm9hz05ewaH4qDpahXSTMEUl7kOn/3JZrivnfx7Ap
SlLzgznZWb49Vd6WakIcHcVWI3ld4DKg03zo4mzE2IWKeq81Vur85hUKKVKz
27bH/s8i06vq1xq1tlXzi79ttQd6WPpfU8KYKfei4oMQ3VE4/Sv9GoLem1RA
Vccfn3N9v93+lzyWUCvSVkBy2E7UVMShhAA2GsTJPTQg5HUZXazrjmkXKdne
X2I3rIcofud467oiKCNiFA2KeH/xvrh4WvTZej1cDWLCGdoLJx14l3kUENKD
jZl3dRIc+SI0I/m4muP3VxaHAtEuanEy62j7sQ7LFQz0ZzWzKgwK3eOwlvQL
r427/TU3jFkZUtcCn04kpLQXBt8j0EMoy5a5I5gxaZiNIvFoBSkXaC8aHGI3
OF14BBlNZq/7gZMO5y69VAgB63pL82/ZipD+79BYvJJ0T55Xa5YxwZnd6Fu9
aOAS1edOSnBua+Wmd6LCbhvC+u5eQoRNcTYW+FUA5UxqQYAMlD4PVZCvXiW7
IZlSqc9MmrCjfdd7WYcnZCg58MqSKGSomedCjo+f2SnmLWBPxRKyzcGQZbwD
8JEXtyHphKA8IUmzQ97R4IMLkP4HrB+n1EM++IfBoQUMge9ogzKgSvCtGwZf
wtS11WEIWT7375ZMFTTU/nWQNMXTnD0KvB1YE7bCCDxCwv3ruM/tMEg7irlB
0lw+zo+dK4AWxI7qIC2E2iKAuFgrHuoaueFv1etOL9YkEKSuDPlAwdTecgcg
7ApZDVAFZeifNrINwWKNAGH2b0OjUwXepPNFzJeyS0R4aO44sUNWQqbABRMh
QLGWd0V9YspEUG7tsPfvkPqpzflOr1yEg/3913g1mrkm41d80btaanQ7Bu9G
BNUy/oda0v0JkwJYgX82k1ZOe0bQLan2oJMI4fLNDYoEFMHqKGk/VQh4TtC8
2eCVX1sEJMEy+EDtBnzTc9knVbRjycwIgrX5DOZL2oqSaMwfuuv8dcQoA9UT
jL/ZutzTG/+Bz9dnpknQ1iB9Uv/lPmgz62h3cDtCeQD8WxHNtZQE+lwmrA9R
y63uQCgEO8Bmvov6yISvCUKg+q3r8dz7tJptoQUfKvBRXN3qDAhGnwJs8NPS
F6+R3yhV9gWTd2Yc+J964KGxG/coX1aQx2eGCjY5efRcDM+H3YpC2nKEye5E
Nz3IaFmWRzy5V+bHEabW/fev6z1THow7NXVyne/GRHHFx2VLD81QW0tHFzjt
8+fB9eNZLfde0w+rL7wNDxF6am9T+cQfdPp9T+yENLewaKco6DiN73Qrcgal
aEb6rhxAFsxq2hDREe2twK8PbUPTCKeva1imSMdgSbTNku/g8cwDpTMWegqt
8DPOOSBUPx+i7L/F6WYGM6ruAcsvhPNB73KSPh4V97Bscajkon0P9kSA8uW7
jIViO6GHWp1feP0HoyG3czfaQkfeObx7pP3kquiunifE3fHK6NbIgdggNP7W
VYgwO9+U+iaGf3S1jAMXJW/Q2kd3pdU6ditL/GsRhVPd64PWX73Di0GsNHr6
DUHCYQ48k5T+1sw6B9OT03LqwPciDtpmw9xdM93x38Zt8W5fW6ep4jreSNWJ
4CE2Dm2nhf/Yr+dj8u3D0UAV9YnZWVYUJ81F4Sb6Qwszn6kZ3vP3GjOuSrYs
RfG/EeOKV8EVfC9by0W2M1Pclzh/H+uItGjbowl1Ix0oO4WYe86bBf8W2i0y
V0SXI+GOdNkWKIR9ao0U7tfi3DE+aaIPfw1b1gQrgokEEe7gZ4D2pB6d2dKp
FrVqZz9k+pWcsmrmqvaViadteD9aUQuDAN5RmlvZwBUYG8fuzXTRZ1YEQrGJ
Jb90wGXlwU3sDiMfIdOrU15gZ1bdqs73VluPpDV5kgGNR1N50xx0uc2MnCmg
Ked0oxfCkpU++Njy8Tx9A/gHSel95GWpeQBMO0IKNRsPwGJl6sjh8zVw1iHO
VflB+wsZA8W4aO1bTUoqsj5O6KjWcSRFxYaz4W2EUyPVnISaQM9F4XIJzpZA
6Us1hwNf6JN0E0qbXAiLGMcUJTrSoDYexMsI5/BiryYAbu26H5NAFDeAfCV5
XYL6z9sZKr3Hpl4Jj8knO35dJtvlY19cgxrglkUnFelZ7hzpw5/LmckQ2EjL
7U1yWCd+0RhvFSte+/hDYGF2PR5oK15rgun+2it/HAVYM5I7GrCQBajj5JtB
huVh29FKjFlVVYQjh5seCf7W/QGZn3nPCsxaxraPwtWri6mlLFP8ajE6nnRs
xaTAzOHhgEM/+2+6v0MkbJPL4rfsbmV+l0AucgjGYJmiBGoMWg0Mpixp4jFh
1qorKteJsK4P86wr8OM3ueU9a2pMxPY8fYy3XRLPnGf554tfCMetqR1GgtKN
0uqzXBqRW/jEtg50Z8z2EgRI2Apo2UQO32VF+E0tVMt/8XI2Gcrapbqcnz33
TRGLu3vinEN2D606CJstVxagzULsjAxnWGs03Rsc2dja40bW9A3VMmOX3jBg
1dliISUoprlaBxrKeqXOzoXT2EOa3d1m6TrS9RJrN+V3vi4hxZ/V+NH9D8Jb
XVHsaplYQ3iuQMtZx1cp7MkFF/hEBh5XuPjVUcEQ2+BxkQtbwzqr6yxBDvaS
VqJWUqIOaou7ErC27frbyCGoet6tY0R1p2SAeTOC7VMn7qMl9zsMPm4CVB+U
YkinDMPgM/rNe9YO1i3ANI/IrsyG3jpp+LKl1iYrwl68n7XjxewYTEAFjumI
uInDJs9MS5+DM4CIW73pCp6x0nA6+J+LGINzNXXiuVOGOmN61GNaRRgtyPcs
riCDMkLzpRhPAz5xM5+fRBRnMQ9zy7Vt1vFvf9jx2v75fOvbI/TR2BTbdwCk
G5pch7H9WQITn7rARfccGsFC//SekQRBXuTIvmMhg8OQkCLDfDkb8ps+k1eY
wK/rANFdRyajConyCfBwiAQ1HrWX4BRwx+6utEfF7xC1fFlJOSIdSY6eqhlL
N0ZRQIXE9kPrreYylZXdIp3vk7hJ6xCflN10gxoKiOXlaSM3TKJFUxCGQRRF
21Boo4wYKTFpsHSzNwzGpj9TC6Z0F+gO0+Rb/ocEM673IXah/ZixY0SRLcjM
mJFiT2e9em9WVom6v07cZy1M8AUZGw13YZNahE0vDiCt96OjOMfZBYihqiob
zefuALfcXdpESeq8OB/xAP3lIqgBkj7EAIQ2i51Wr/z+3H+jPUri3A+VZwdZ
VVptpV4PY4iswPVEWdYpMqp0djavMOeF77UxLNUvBAU0ytyXQzUt3+97ehHS
DjJccELZK4+2COuQpAacNfu1x21UWJMxNduzlWyP3UqHRELhn1xf4FtPi3ri
9lpYT5gtrxCLbYTStjYbwu1gG0c1kdFgrLMYzORl/+KtM6ncdftif/+Y7SM2
iGHUY2fQe6RX2/PrQK2IM9WHTR465sR44rYigX4vV+RoCtYEuHRpANHV7vT3
asER+hKN6xXgW3RjMqllBiDhoPkgcZ6fKfWQ8IU7CSrDd6lFoPw2SD3jCYu1
2q1mWON/dCu4HZzGJr6p2fwnY02Xlol5FhHtvb24jYkcCYIJS5wk5ciYGFMA
EKCsJT7a0PwOJZ6k1MNPsIId2lrw9F6UDrmr1RYVPkXiboKEiFWaHA6jTLML
VgLyJ3iqTuA94Bm1ROdFtGSGZQj/vy187QS164JQ0FyG+WSolav67bUNe3jk
eWJnA51jjyq9Bo6yx/vj7Z0ArpqWmGqqPLfb4VyCx3YGibRUSR38kWIfuMDh
EXR9NqExD3UVh8H2DvBcKpdmeKgEI/6C/RlyyM1iOipsJLVNmgvw8K3o95Mz
PLrLbJVxJMQGy64t1KqeG8p8RPkEKC32WHBkCj0j5fIMLRAGS/EycByt64/k
SzNeq9iEyqe+9k204zHMftE6cYvcv7Ip3eZEFf71YuzfUVQrQJE5z1ro0SVQ
gq5Mx9I722gAD9gssqL7UPKHgvMHG8lLB0cVOvOxCjAgq+bAO6tBFiO8f3IH
JfPtUO/QkOsL8hr33uQBbeiRgY9nKmR6awmEi3eE7LWktwB7n/Ut2XwiDZR0
+tre9T05bAtUm3BRuJN8yVZaeI2lDbuupny7kiAiWkuwemZ36tviyjR4cW3F
/9k15nTJM95TnWYlrxwCAnCFvhzj/ielQsyCTe4TrypbazTJqrS6VM6VQQ79
jFUUBUfZeAVSlxu0O/uknSPWLvd3IUtGmRqR+s3YnXgdq1KzU/gvnULs0BNR
Pob0EVfwu8kCSiwkm63H2PnlCPv93L5zd521I5+DK+HeUW2G83Kvt/JlyS42
AAz5djupeA5Vkjvj3mhUc7o+NG8vQ4eN36wLmls3m8uy+yKOPjqpQ04GP8U3
Zy7u/FqYkIL1+lLCvasOMf8xS8FZ0NqVAznq5n601JDzdScIFJa4h4FNg2es
GypkC856kL4FL8DTVvEliFGh8mUE3v3l37+W25idbfJwt9cLEa5jYF5aJ0eP
PrzbRMTUvRjCkNGwhwhwkconVqItsjw/1gtvOSCwqLZ4w0CMHu+vhNTptCZS
tUg5OUgd4SYFlCoAo+6wEEVPsQMGJTPzcw9/KhwhOmTdxKNmmfgfPLBhFPn2
FgIa5F3a00ep2PUsugdqKsv7sQ7pKswFtCgk0lTzkL33J0UY+Jqxl1DyK48R
r+mWC7I4DXEvMdvfNGGhETEwaACYkxJvXHRkHNjiz3WPVHttV7FxNSksmpQY
OTYn6nlBVhjhJeeHepB8VfsAvqTujBewU3/Ma2H9HSw8MNgPdeegwuB8222H
wI9jS8VortreCgAIX1JmjA+57suC3kQaEDIybkUbNLa5cwJySbH7t1EWTnL0
ZraLt9X7H786pWt2+7EcpgIOhjHRCXSNzJogez0pcKFCXbnDq/XdQU0S8nHI
AHA2xi+XfHmysOAAeEKAM1joP0cI3JBzgHfIrK/9kXXxMr4fg2zaVKMLVxXR
RNu9ZeSQ36ioBsi5Rpk3h2lPhyGcQ+rYKNCfkrwBj0wSkBKhWrAcwlTQ8VvV
+g1tARBDoxqvlMEpvB3ASjy0u1VkFjIIpc7CU+Ch/wuA540BzQ5hOXi4rgv5
wUBuThanX5q242Oowf41tyVzgrEhIhv7FDwecGbNboR1R3dAvXeaFTYG1FrL
7p/nAC2nGwDrYvlu0oRpuMHY4pQ81wjyymRZiMnu0y/ano5P20eNJK0gYvaB
S/QjVaWcI0sRKovfNvM1ymM2BxflZfLJPLRwBpqtTa21N+EW+UvzqQGpPRMi
zyFE15ajJsDPbQ7aZw0Fbi4MifRri3tqoYWcFOBnPWMW3m8gYyvxrVlYiYUI
LVqGGbx29PJxqi3m66DGGyZPROyR2pBmhTqt4zwEoFhy3/XiGQbVbJAuUR+p
Lxvs77p9Yx//oJRoBsh0sEmAwILsWCJu0dovyVUUxF0AmjJvbFGSFw+99/Io
rFnxj+PWeeux0xvIUNyfOqkzHlcl5hkwnGBUjxbmVLKqyBZpPQ5GWMb36apX
WjFTxfjeolb9WClK+YpU6x4ba9PVlJjmBDRN2wNk5q8c4JoIEvvoX6ARRXf3
7geZb614dKl5HLmWVWO8JSLuEL9CHtf8yPSLfqEznWrq7Z/ZHCrkYLuZhah0
HVmrr5WB4EX7IznK8+FLV1BnPM9jURSW9AZzyqm/klcqrjGunAKzDWD7lT5B
YUFs1TVUUhDqrwQb0aKuIf1k4MBLPOgrLia+45T809yWYdXGUgAwDK/0fiur
8nFVcCI18tzX6jOEnV/bEyCii4GS0bYrDrYfWh3Fen/pm/3PfqHJUXS6Xljt
5/COzbRnW54L7/p5MSEn2185AE8ULGEcd3VdrX94HCUisRcQLZpJ0mYP31kI
xiUmYmrq9bSvZcZvDAEe4G/LMBgTEjBObT4ucjxapB2icGPNM2NwU/rxzM7K
3PPrGs0422GOqgk3UlnDWEbekvpRVXawaxxiF7Mg66HYUsoKplFaJ/xPxOH0
fJ1wm4vg+PW8IYBybbouVwH9VJEC3qmogR3Uuo9ZsGq37hlkMOjzGD+KpdNw
1kh5MAHW4ZA6PmO4JjbH0ag4BXupOr7UKnoWCYSM07vBJGN7OjSwCzHRvww/
5YEAFEIE++ZT6NDEpJXjFvEdnf37IEHsEgbD8R/aJ5lmJwW+vgM8ayegU130
6c3OJZs3JXhRUByqM2cRshKg7s/jk3BdHPKi4SrNs25i4cx5IaGgogLavENc
wtrVty/FRKlll4sHiV57Ek6Sn0UsqW78j9bjw304dr+u0z6EP/s9wW7gpx+G
QT4rT06vMd+jAAI4/bL5LEMuPFY4Zfn7BH8+W0um5ovJvl5sT7gB5lylI4RK
RmXhn6rj0SvxWlhdb/+5V48QcwscWVxvQGNUmMLdtH0pNfR6WIIMeAQApAi8
qITySY/CWnlDN48/F8SMnQMeiUBbG0/nuhmFGGLFz4fCGrLaj1W3BB5/jlx/
V2zeJMCanair8xDWB5CCwI28P72U6bMFcWS7tpUAHm+HplUkWXldqqPiOxIm
YghsbWw5XbQvgHlm3ylZbLLEGX4rL0RGcwvhAUJNl2xsjUaAWUcpd6hQmcQj
2EEKpu0wkzBc3EWvivxriKILO9nYUm37m5QHeoi7KwM4U04VUmVod9wu5x2T
g9B/HvQrd1OAfeUeHjV3P+DhbzU+vCtNAyg9HSoEiscDZy471D0EiFun/qmo
yF8gU77hrOornCmNRHrsYUBiqR3d8YnpHzhTMMlnu53Qb8b055TfyI84BnPC
xWIZA2W7c+HAVYvo16Mbnq+xNG8ucT5zX6YLQ2yA/NEqDqmXmmXxmLFc8r/J
wDOWNW300S1fvlMV05Fv9EX4iCp1nZp9I4iAExxnk3QfXKB8Bepf1TavESFD
efmuzWdxBdXgdvOpvkfat5PfXmqQyQRAwjaippd4clIMiXNkYFGGu0Ix+TMm
2CBPLVxnbmuXC8B7uJCmv0srUpRnfuYdWqtWRrHcrxncxd8vkxJq0bm1+1zG
E7WEldupteYT3w0DidLmVxHQsDq7w9c0oEj14bFc/ZyLGwLeKQOSyHTZsy/Y
k4K0NFgBjUtN7mjAxv0W7ElYKXBu2dH3cgCpAqineCj5BFt0MLcWYAUkPYKg
v23jrBi0fm+rFcILJJesVy2xag/iUP5fGAheNYXsC2awm5QV+Knw/HMebmv9
d+eIJSlKSZwzNTlElwSpJLgZH0SQjliL+vmk1pHgB7txz/jOXNvAHgkVEH+2
GxZBPlZRKQNny6QjAsHGrYxe3cZurTR5lgHoCFJYa0tlydjJ0RzisW1F2kHq
xBxzWRH7CHF6G3IJRbsvaAeFBFvex+Q1/jBfslwJ6M5GHpyOU3s4MmJr3gVe
4bM5XYFelGT1DXSvFpHEJ6glnEP29Ys6Bnjy7GT9b66WshuEEcg+0ZMQxqOX
xGP1I0IeIpTZSU6RjzNJNGPAoMBTTBtaHffQ8CQzScDDWy1e/vJwkxzJZYRQ
ZO/RYMRbOhMfqJrvm/3lwWODiH4pJhOLbCwUnvVLGHsc0SgL/Lras5FUesZV
ehZ2z15Jqb4JyhS6KhRBghgxwH2bVTOfYRJDT2ouL7pTOtapI2vtTI/NRt8a
Q5+LYgRuthU8p6W5xJ4HobzEIpZ2keUkgoHXk5ebq77RtXFDsFJN9RCJgc36
krCSdYF/H5pAbFn+oNnltn9yzvRB9X1NOJFMx2R1D0OhToqHVvxw0+pL2Xn0
6rHwMszFu/M7S15i+2Nd/NiIR7pIAN/bKwIFZBrmbqv+K0P2hNADZGVcjMpZ
GbclLQwCL6WQL3XXEDRN3CoxdD4A4qOs/E0KC/biLJZiX0PpndrHXOPA4ium
rHEqHbD4RLRar8nV9u7eXbrK+Jc0qTXg4U4guaTbEoFD1BtRfNMB60QJrM+Z
hynR7XX5nQCdBUBoA/PAb1rPIv30Wroq36+olKnG2FM3eEil7b74G6ryXWZu
HZL3PvwuSHoBnZPV5/0lcfVl0A/CHgZtFqVjOTOwlIHQyrSp4Uo6KTWP+pJ2
dZbqTxa6w5QbTvs+LqTGTNnvsJoL2PXeyWhpeClVA3yvDDapG8AL+pktyLfY
HZZ+OhgSU/B9b6b7FTQZH4tHygOOKtiYNO5jq+Wj0dZeG8JkgTrXx6k2TbLW
fton/3hqnRq7LbCacDIIpPtClcLRXHvUTnip11uREy+qn9r+6HnNDcM2OLHY
WQc+/nEUpUW73y4yjJ8vjCAL8Od8KsuE7YXGBBKVXYJ/9wZN5alP7s5l0v8R
396tC0Oc3m4kHKsTEN/7THBigcVO8kBPiEf1VZ8FwgIRauXWdnU0dTOMRt3I
fQonYVo3086jqInSkQjGgGRnZMzRGc9m10olZlFwg7V+loAJVtwxK5r7tXLd
d4q3B1PkSucTw2zFqznxDg7c3jMTTj6y8XQZLwCNivAyiR3D01eylRz3R3/8
JfF/Hd9FZtQYGtsGIqoWdm+5eT5mI/JG9zMyykoAW5oYBFMb7gulwihb+bds
9XtlfJvbQGDdkICRGRhojwryEteIKSDL1mKhnmjtAfC/R8a+776VbV1XoM3R
1XVqTyCryRQTZQZIDwlEG2QgXH1CK4wFsQ/rqAET1vosaqI+V5pBCH+kKpQA
n7+/p7DOctNBAl+3HUdcegA+8RKs7sf2OIdDxnbCTq/D7JjEbX7zDLrWvF+Q
6cgg3IQ/f/fFn6a9rifgM43wDt/1AvHbCte8jYnKri4xvJxJh7ntLOyJ9liK
TCzw4HOWCuEvXK2pttVJDvdubrWC/BMaSH4Qf/jg53jxxFYcs4O1BApjr4G0
+oEFgE8OMUdAzIjZTzWwNFmwYn3cuF1Ngvm5HzTkwlxWcSnpAAAmCAYzY9mZ
OvosG7vC5B65Sxujr3xEWJodpGq6g/e6Ek1WzfrVXolVQdJMqmQBnI7YAjMo
lMXSWoZ5WDQOwS/74J+n71hP0I2IABOk8/KGa+jKfTaU8LxANaK2uoLSjmjR
hUQnZsFmfny9gTYEyX9mcP42NkjusU1kVURtcuNoo14g/zLxUyFsu1fcQO9f
LSkaQ3FPZX85ViVJFANt0yq8hW6Ngax4tHmyRhKWHkqGhytGFpC4LZg9XVqm
QS4FvClUtpTpQ6o8UiOZbXyAW99xaVFq+IdrfWPLGAhy4of8r5TysWOeF7AX
rT4yzsdJJoHcbCNYWmFkUq0JV78dJq3BBkP5Y7BMLZvbWoa/9MyL8U0Z5b34
2LBmXMZ35xjHATmZmU2S5XvoIzus5jS9nGa3JTBdoU4M0U+8qGULVGmRemm7
i/+3j3sVg3BmwiXTkyaoqc0jYFD531NfLL8C/U4dDwOofxUpabF6eQ6JHgYt
ynJCeV1rW4vtTthk/QDIdB5S5pANelHrQ71eTmZKL4IJEIkfAoFZfYOflimg
rgySItO7eWFZyxri6yje04pWZYGTCyo1JK5ox8jvD94t9xWOc99cZlofLZRU
aIm6BUjSoB45UhURS5BZpzSsLaBh

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JUjdpeWrcOjupJW+UMMufP49z0b6hImiPMaq0zOf3k+YExSM/UqUTZYxDEEz7eI/rz7b3ao5fAY4hEQ9B1tCYHNeWgpkAECxrD7vR8DimfUUwRkd4Xq14kq14goHPD58CUaekayIS7W80vsuL6HSQp/pBTGlC9FCvAAYODe4pbvoGv3nyoYR0Dd9m4nA30JGGMKkoqLkUzfS4fDyrwqnSfR9ZQuzAclDUbttO3UiezFBAps18eoxGjAd0V1ab2VMqAqlX/v2lkoGLMzfWnMHX74EC9/GrWOocHm1Lhl5L+XggbvbJxH8lttN9t6+1jUVIzgVhqoLQBfVUuGHPJT7qivLy5jZlE4gMwNjmVc8qRAyJJmXjEeC0ZIBygAkOtEtqL31zpwc1TgDRcW+sNm7h2RQUEpRCsVRP7Ja8gOL4EOY5SUdy8tK1JodlZNjSTizQ/yJFJ+rMHXr2km9hC5gvGMaEJ3GpTRmCjc/9+hnQ9vcNHrdNtihOsdHCMuCox5rFiYyi8asLi+FVyHqMyaXGE0ZeZxdWLSx6OP+a3A4e3TAUXAlQgNWRtx0haGVVc99JztIy0XIhE/oJK53smg0Ks67trKMU00y5gi9Kz5/7zNfHJpLSKMAzlGq/N3UeeEj9XeOCweOTZQy8I+MhBZwjNztP4STqdYfgOXMmKGqXoKwBtKep63Qy07xsnxcE3cmyU791OlKmRvIiFfiSfADa9zgE549lBMN57qBsSZXQN+B2+a9TacriB5lTLpNz16XsdEnT7eEPNC7n1tdvY2k62"
`endif