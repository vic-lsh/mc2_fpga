// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sGXidr/nP1nz0F7drEoGjboapNFgsSEUMUxY/S9BtD6gAQrl3Pq1Bm0vK1I3
/UMlncSEbmhrFRW9nzVKMQVHVTheDuq3Uk1lz/Gu2oMr2CXt+otmoI0izssc
ErI+0LGo9m9kH7bCajn7jUkTwtPd0VX6NHK6ynrBhBt51jLiJidKp9oRFqNV
qsB4Tj9kfLzDNlSTf5EiCwe/Lyh6+PxMI84wIBiBqQnMqk71Orv8sGXT61Ke
bgTyN0Wli6vgNe0hojLul96V/hK5zfaTmfCWlT85v5GPN3frERoFqwI4TWi2
DuezAOkFcP7NECYf/PuPqF/LK5v10NwqdWOyaBdPDg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jxuOE0XGB2AT9D7DIslrdysxCg+gVkk4wk20QCHp2ywFNYu1dxaCvjWco1dr
y2b1cggStwk27sbL4pFCFTa0ekedjfExRwyDelbqE3e0lQhVq0vtzzo5z+f+
r20po35fIGq6A33soxQyxwqAsCRG8nUHILucuEj/xo5V9lMhH0QIa/0ycxK8
6hGcSj/34v4ozv8kXfCONb8rpfHUNLWs8EZXgGhMWsfq6XSR4UPJ83mXhqFQ
ETMc9m6CLqMvSXPzyenHdrC571f7DHfLqIuxli2GGIMtK1m0INrEQLbQCj0B
uDkAipZO/zAFk9XRWFLSEkoAw8M0R2G49oMxAom9KQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UImzTAjhPQjysD5X74fDdqkkDA9/6kVM5Ircqdm8LWUa0athw5/FFVIBQT6u
bVpvYUnvN3FeT6yj9FDfWWqkZof1C2CmVp92l/hvTZBSYrsvV04KpkxT2SLO
vkLa8FOTZ7Jo36lXpFkYlnQXwWNW9/Bzdfy3vzjeGG1k9oQ+SluALTbnJvAS
eavUeUymGfjVEY1Uxxl/7aFmcORMFFDdlbuO1IA0ZF2k1HnFR3wNoTZOjGcs
M+EjTTkYfewzCLAShFW2VxrwoK5l27ngXb7RGv+SEUzfLom4yne7WFbSSleb
5qdPKRCUHHV6imuMLs+C4Rkx3bw4l7wE8Q0pSQRejA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nvpMpiE3Ltu4l+KwvH7Fx4w9+f3ez/cqBiQKt685UEMdDU2FUUqbXl0lj5DM
GSkFsB38ghZn3QdWAVI+8nx6eTM2+Ma0v8tySNXyOJAz4NdxUyIEXRuxEPdU
RPgciot2EfSf7mSRTkGtnOsE6y0yhXmdFKo219vHoa15h6UpjVvomWR+vitU
nBCOauMVr8oeUpkz3FMgVY7I5lw9AyC7XXL9vhDeLDo/UyvfSkP7HXvSgcb1
YNQnkjPB7Fm80lhO95ZvXqjyr8pd9vel6tlB9D6mnN5IJ10kAeAwzCni0Xyl
6Ee4/d5hOFXfr2pSC5Y9NjY9idiH0fwCptnVvm+TEA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NySgqI6K4I0eOxNWy6uFFY6jrWG0GZ6JI3usr8HAinIx+yz2WKgP4VVGaPcA
bsfd02hAErSMqMuWVU5D/XsKfJIxf/TIgPz8dMxi/pQvCftC/+e81Rw1nfao
K1BXtSr+/cSeVQz5BeAu4u8D1bR1kvEHD2MT6bzjUzvnuqrS2Ow=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HFhvUVTUY4x5RsbGL5ZoiW7o8rGukMiM3/ouQMqCsMls8Wwx6cnao6m1+ayD
eNZ9ULV4SLi6m9kod+HepIWar2LxrYfpjtEIdSES/CZhmnGocayAZqPJBJsg
wJL2fYRIuZzE92G3l1lp/Ue3zKFL+nDYdkJFIwgmBGwpd7y7Ai1JReV13ASI
tFskVj0MmrKSZTdKaZoQQBSlxasB0xkp7DDvyXxUgirSaTedDfoba2s1EZfC
wAgIGy34VmdIOky5uLL+A6JYKMzyxm6iLLOKH5Qbj0mO/JNXDoG9f9Uplsu7
XrnGeoJ8Cuof3w1S0y97cKG5OiE9IfLK7y+g/3HX88EEZnI0ziEZ0GA/5m3w
qnmTV9ZDMzJVsqST7FBEFaEZUc54p+Shg/0BEy6PFW3uxHeR0WBqB43zpZtO
q3BAP6ya6VMchdI/8ptrTfanh+tBv81ExrawttkVtU38W1Ot+8vE23eksR79
BzlMF2SXIPBEIaqjVhUiPFcihpjkZuDq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TFHZNUPe60wGjnLy0QV+g/hmbyotn9OPvyOkOP5rhh0MDwB1dl7hYIHJLeAQ
MaY0Nxle7jhkC9tBRa9WxyG/lZihsAmLug6fAKx33oi8YW9dM8ncNDwiDlxG
1VYda7v2lFKmSLPJwmrKxFsnAiRueG69ac/xQDAtPH9OLX4c+Oo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DpwFWAuyK8kcOI/B0m+Ovp1OZ9hXPQhVPkaYceYLJRXiihiNFdD3IyIaQVst
g8JbziWuyfMV28YnFKw1YSGgU8nyi+t+e5gCHQEdPabtBeExTShGTEmMpECn
EuGI0FK0c200Zie1fHaZlpR3YqXYINbptFJ5btMcIqIvMmM3IuI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 53776)
`pragma protect data_block
kZkllnCZ13QpIE3fF6OJ8VCaZp09uVUKdbVet3Q74hoqsawJcrY7F74FOJ1c
/PTTFdXf9gwhFHjs4rTrxQTFphG4A/UAqoYog/BwtZQDZnc92jMoYSnyY+xY
f+T9bROKl5nSAiV8BVbvNQCnG1ddnDLETQIYiJGtRAP7PVxB7IA39IlBwAm1
ru+09/hE16PNNdsOhEb2Crtlk78oGn+oIdLTC1c2hyaHRTy4ZNnBA/bV1X2q
fmxaJ4LhnYvipYr31fOZlRFb4tR1LWI0f8syjCJRXHPoidbPCkEnTVNW4cPI
dqRzRwmZbvlgsvlAe7gmXMNmBLiYchFOPpUpjX7c+oVIs0x7df7/9qdfyAJT
8B8LaovyE8pyeIgMaT67oR7Rjc3CgiIo+6kbwxS+EJegUDiK+fgRm58nEpmH
huezqbQdZyKccXlHIMbahMV+58b6h5zSNu/r2ccAVA0HtBQ0CTcUmv3V3Phs
aMjKZdRmdoFyyphUYT7PzAW09+6rekQPg80lb+AdajOMArWya9C2zK+TEmaW
pdCvR7yzUtbs8IGO6Lss9VLFXK45x5IVSOfU2vca5lOU6K8ezraDxvbAObRq
Mw1kOJHowp03vhxm7zEOGxHsHGB+6LQfnEiabKKY8ob/7qv8fibA05RnA7kB
kHqqg8kIWdNEY2R5dNNqNprD+RJH2DEbzG5zibkYqIQE7Taxn+NChPjxIvsc
FYklMVqLin5VCeOD346GKz18Hg+IomhFblGAMsMCc38+v4S44s/TZbSZkPeZ
5u1qiTLnUxMxo+oZHPzwO09yOHmny4lxg2RTALt65iQvAPdBpg7df0oLYgxo
ReKjjxzDPSi6+B37jEsdzsnOJLdV938qrg5VzgIEXnsk9tgbK5+n5gQN25CY
ki1qM9izhrMqpBIpFTu0/8oCI+VXdByYTujm+q+b4Yj+Ppt633hTCrHepl27
21gFas1oHjzCSJzm+FDTmGYIyfZXqzWpzIa2eemvDHCPdwzZmfssOxyZ2rVC
ySktHN8KteS055xRcKIrNrCWwXgnPpdLgUcDsePmdqVeoWcqlkiySr3/iuHi
ZeVWNh8hZ+FTGXqmQfxdzsrclZq3Dy+wOeEcg/FWqUtrjVJwDgbd63WEHr+P
nQzdVmW79yXmAf41IiCUcIuYi/UxWT3G3UOJJMxPFQR5t+HcQRKSLr+ADhzO
8WLpzYVOqDRiU3BwGfIdh/CN/FCrYECYimMkPHCLugFmHhNYtQjvbichCmCv
p002IOX2sFM8I5eOxl1QUrywdt+b8V23oXRuv5pmSOCDTLU3AHD5fVri8WDT
wIyuJdvxx94AGJcY0cCunGSPAakE31GURe8v3tzkQsfHSydFD6sii4ubAVFk
F/lEQZSq5TdHBewT6UvEXbUOuyFHJcMakE0+rpC6alYDOD/qs11B7674Vvy3
GW/5Xk9oIi8bdJKxYEoYVX6gDxW9+A9N5GvF19Nxgp0xUvjWD5FavgB+FW6c
/CeROfQCSXibpO8cfOQanUKA158xwQUkCR9m6ArHYTEtPLWYBK6orY9EvDdz
G1EWrZxYXnarCOq5Nl3GzqgJ6MRj2CG/FnmpYLc4HZiA4UBIY4EiPkpeJABT
veov09WLZ5u2IRh1AfTFfJVOLZYD9ofWaZSio47Bem3jc1bMOR/gI6JBjZyp
q5UbUFfiZXTq8tExtUWjHcpPxylhf5g4IDsDMYTV4oCfEXuoa3n5AfCAgvQE
SOQvu/WsfkOfkzHuuZA/xwnoYh5+9vzUU8KqbVsSUpkjBR+6TGRTbkinnIWi
BovBvMx27NImGtY+90vq/YzAckZiR1TBaw4qqgx3EXazNc5zHdibEplCD0P2
7v5Iimi1FlQe2eNykxZu7j4qTqHbbiIMZjyjxpXGQmBXLZAqQDEGel78kN1s
aCsw3WXt3JxdNG9VsR/u5gwBAaN2TIZNXksfrwwvce/preFHOSP+VVg2LaTI
n/Vh19/oFa0xpN2E9VSJ4FHawAzxhVY68oB8pqL82Y2GfR2iVY2uFSCN3E6x
wJj3x2NDELj8SigjC+ulvCrYz73iQnD+0Xs6heLb0O2Np1Xheg09otAOa1KZ
FVPn3WR1tpMaqdSQvHpgh65jj6y+U+zEWcdjLrPIgjnD+nhd7UAo98wk4aAJ
FDzsWdKzjUbxl/zcXT9/fDDXtDEYkKrrknrvxpHZXFEMjua90P25NG1ynxhy
kKaVSUy8pBcxumtptJF0JPgRtMFvQF2WwmRy3TMl1iQ3YNCuzeZ8XOoESeLD
Lsam7XK+ydABib7h68AMUABk8DiPmhKwjwN2V+XaiyE8uOhdw7sNcJcMWoPt
/UvawD6oHes6Mc1jQpxTwZM7zY1i8Q7tEJ7+dOYvBPtu/qU/5qRhttKw9dE3
zqqq0nsvYMKw5C/0AlknVx8MAhf+zVFuQCmUEYNiS1aOn+XVOkdFzGFdOhyk
ve41lvuxzali1MYCExBplogSDeRYQy8lfBGdu7Om7BfKv6HDQ4j/twZTTz92
N8iFMwiACqQ9Li5eGA6RBXLlL0mWEelGShmXvftLZHe1w0PZvdriyki1QKE9
pJzW5hNDDMPKdK9wIRFtslXXgsktqxG4et4mWS/tjKQYHncW9hcsUo6hDeji
adHuKYTZUJoZIsrjufCg0fD0cWFqFj5qAB2E0uVZqxFgvweGOx6HWZdWI4rT
PRPzexwR4kcMVLxYu8h/d6sSHbmCvbtgZ37VJi8j6tsnCr7pqRHx8JdsSVpC
Ki3pSjcD5kzbnjU7lPxIORVYknQ/6Gcq8iwc1jbYEo04Sz6ArjIccqXK9dDD
OawVMVicg8gQNfAWW9rxpfvs5CfMGrWqj84+IKyXptGa0WzPDW4wtRli/jF+
W25a5tA20FnMLnJyudjTZRV57QtmV5bg/xnYpjFlU27wzL9Hu1RuqECP74cV
ezPUCNTkt1RZluldgW8OlifCcHANrqyl661OzGfqnJqgPcqvt0+qk6W4TWTi
RAEQsBIvxBQiIBj+522xU7dV58CSR9fJ+87FGpwmfeW/eczy33AQ/xHNhBYZ
vOEi4XXzSc2Ki+EHN8AFfP4XYkhPwapIfE9+PpFDzKwlm/1fZpYRXqJCC5vj
3iqWvyceAaDQogUqaDBTINDM3BoOUqcLHAr3wBR2lYQjX3b4SwaGgh/Vgx0X
iPLjFsf0yEbLO+AgSvh/kRPNZb2jxSDRr3neEWL3RvCAjSDUhvtetyO7VS6u
3R31RCOmWqB/G0GvFSY7bMi7CREzvKewqxc4jltx3h4O3ovmRDAlyU/IBKRx
pVHOciC5XRVJ7W87JdXH81J3zA8+SNCwwY796VLDXpDeZCbrf+6ZSVvScH3K
nWNWPFPgG2MDgHN4rhITWPLkl9+UB7++zXWmDmKohmduQq8301TmAQkakAkB
+ctDiQ7aDKdZ0V13w6xwmururCe+Y+8gZt8nRKXA+x41ajhIgfMQ0AexXplw
79BaWirF/bEA7YDuntpmiaiR56N+80WHtxXumYnz/5MbXDHees8lN6l8Hs27
r559v4o7wj7Twt/IpMzAPAQqr1vbFo9lteTw41WT/n1kCIY88SGefo1nSrao
Qjn+rXPr/Y9GlINJ5czLfQWv+6YRLh79R9y8bX20ck0jx8dHIP+nsOSKG9/t
WT+jhhKZJ3vejbYOcq4vAHxf5W8wbxt2dneefKj7DaGRshvGink+fQpaeVH6
9eFHONbtvF34pGVOqrOV2c6Zo68fF3SWo6+0ngE3xdZQvVzRxXH9wskzyxhs
J/tEEIhfb3ii83mXhyPq446D1PISqcxtI+gq0/fn0+oRpGbdEaGL9KBkT7Tr
ESKMthUV+KPjPdbWCbnf8lMkDUv94Kzd9kmQtHiQGHdR1Ekqq8yLccGHMTXP
ITXJtk+k1uICj4m2I4baSnq9f0wuqlyq3/N0O7eqdbSsEBg0SjYqETWtWidx
NnjELUcHe2MK0zBoRQU/A8Fw3SFT7ZtiPqrsqZg0eNCV/Zb1Q43ln5sJN90q
LbsMOVX+gshojUrYDoxZxAjRaZvRLnVfFDdJ2VDe7JkZrHhsbgjIaq4xl2TO
gz1j8we8b5T7weDFyPQeVjO1EfETsO8a4LjT7k1FKpaVhPemtwMNWte7ToBF
kWudvDk44I5hgrNKnjpnnoCRSTlJIEHSpxkXFolX55MmRdIOi9w+WpQMNvCv
lsRUA6bFqriRFTgLisRhsgLjCdXLZ4KjJfzPN0Kj6Pu/YuXXw3vQAKoOeAAf
lNHaMtPwqfcip6cGKT7FBhbgF1qRV/P/npaWE89O9H1omF76bAQAYMwFvJpj
kZe6RsGDVYg6bCnaKUsP75zHApuOocWi40PH/Az8He+seB51nRqOvwzvj29n
YDHmdTu5dluOtyrQcwTyakADDa39V4OKm1kyCnTvSoZ/6M7U9YWgSeDUfTYQ
IWl4GyeY5cL4qbLlEv9UxhV0kmJk+UzWJZarNBRORuIt7KcOK5GbA1ImUDWV
1Z8Kz/iMe8tseEpRGVlw6LYq153T9Nhxa2bO7v6W2n1XoDumB8vMJWB6c+M3
fdz81Zpta3cBQKcBrorHSrWO0tXvGrVM2cORbDoRPy9KaFIwuRMmLAUf5MvS
KSZdQbAxZ5e5MQgazC5s2fQSihiZgUMWE3N38wNdqYjjUJmd1DMNcBRFbHqZ
y6U0BPfIbB6aZ/hkt0tprpDwPZ1ikjpgPv+X3MtS+v8djvlX/VSgBytJPvqm
sI9cOkJsQwgd+zdIUP5eLTnHIPFF2r3kDtTC932g/7A2xOC2/B/q6vK/asmJ
EY88OuJZCz4YaKpQ4REUDc+Ego20c/jsxEyFuRhRnFiDnLyFsLuVtFxjmaxr
KZvN6WTEgZFQ2oKtrECHIE/AIOkXAWoRP2E1Eutnswt4Zo8QZFxTk8n+XVEu
aM823iYMjQMqfCqe9nH2CVTgloBM3Fk4q9/Iyf14Bi8sUFrMq26Ogxr5iwVX
OvL2lPcsJCI9bjFnMtosFd2AaU41IgpO2CsFOUH69G+FkxuoQoAjZM+Ga+jz
EH6Ng3ttC61N8R541LKov5VeUd/uFgXKNoGqBuS663GTYq0bv4R3hCoTJ7ow
eVgvGNoU+YzEVMjSmSi8ZeGIxIfiazvrwbS+NQxAVRqV8ZT1V4hj/ptH+cdS
Xy2E3cj3ritQeQ/a7/MshAly0qbCOUHdxS5Q+SWblOk7EOtAEBpkE/Y7yoaH
HwNDHG+zhOHFtQ4afypl2QpYeufEHybv94zpxasqmkhGTYv09OXZ+YyGr6EP
FAl746mq0tnyyf2lSomPeGQCbfld9a/pAbVVirDTLQ9463NyMfLly1OFxs99
03rRfxVH/41d6LaKCs+a8VXm9FteVFtFAKrwBs/1SUC4cCs10CcGX7+KLm7A
krrhHLPnGG8hZXlyQju7yyu1cEaUghcQaOaVokN+E3/CWpyJ33eIXoSFN+SE
zhzzM/PMIOQoX3YOATjpznd51ez53QMp7XD0JrQAKGIQs5z19hZyyNiLn0Vn
QM0V/GlogOFQIdhhygh2V+zVnM5ZkuJNIoBfqqDCYyM0t54aip8K78nl8krq
fb0TvIaQEr7ktkr98PPCcaYktrHT6cXEO02QiFnhtP/Cgub0dLKx+v3an+0Z
FaZFtm054YGKnC+GlkXHnHxUbnaUMH+K0MmQ58sBVKC3EKZQvodExWUgqvMU
3/MrevbH06Vj/1ctd7zk2rBX8D5Pinmhj0e1XPaNqvmtMyb2KASSVN5vfWYa
0ZxS6iDek78iqCU8n2CTlyRo8FYHakBQ1ALxX+4YXBqLeQDJ/5aBOnA+4mFt
+yR0n0xSaQE5BI4cxLDi8zemfZ7ySYee95eLcgH25QBaUz6LhgdMvYl/j1JF
hE5fFmckLOtSBYJIBYEhDf9PdI9ua4j8dKd0VfSvi2gv1DN6y1ZTG2V6onVl
LkZ1qxEnpLYF9lzD9T5bmLcMErI9ZdB2PLS6NGbNY33AZ5x8u598lEahJE71
i3rpVUR7oKVL8Nw26njvb3YpIoqRB4G+QjoaFdvMdJWeurErjXh2jAxOpz6u
xcYs6ioEtoyGynB6/r2mdGMnPpwTvfGEjOC1+0/DpoxMQV+iaJl9iBJnjfTP
nGULPwVl27lPIVTgeGwt1m6tUAV5uZoVvvnduOKO11HNjZlyWc3ncmGAnjWi
lpdSARSIcJ9PTfUEf2S5D9gPDiUAX/Gd0XeHWo4nIGM8GNTmjyfNeZQylAho
fjMV5YHtXkyoD+29dP903Yzxt76i6WGW+E5Ao4EJrpZ5ZET380GQVO1Es6Yf
3SC+Xc8iNEQn/EtZVnkr75g95H5WQZO7a7HEi9SMAhgcBatVb7KuB99dN7QU
rBWHGRFXe9GuDBuja6QqrKEU7Xx+zsFKnSqYAGqoVEQZCU5Htr9l1AXAX6l8
NNl9BewUw4Lfg1hXQeFw1yTOeq8Pj6Ft58z7XL9wbj0rbuCCTw8Rhg6asvMw
B2fPJqKoGYzptc75psdd/gKR5rsrumwnW+UDEiDJPXwDDB9ITyg5R/8KyVvA
B14VQT9HYDdnYt0BBMbPE15AtuCKDGpYmRhiKKbxQ1hD7QH0eqqh6jyUwf03
CnjRGZrEr7eRr0yrVbyVPAQHhKgYuMlTF2PAS+m+iMLh25ibt43wb+yrUXm8
n1jhBHtvlTNgNd198BEO/kJ6gTWDronv5+sI53iJH3i6iUvyaNmwCvkhzl20
fxunicSpVocnIPCZoX7Lf6nOYZFr4FmBy1Jzkliwo5DWj4+qIGONLU1UhZ4n
ZWXgYzRG2+l6/w8pyFPo1RYPUQlP/nJSNSZcy17SbZLNog2ORYUmd9fRXNiL
+yJOz/R02QhDO5lZb0ABtss1L9AoyDJB5gzPhGt5DaQ50jmTI1C8ALE8Cd/m
gscZPYHGzYKMOO4Ym/Zc4KhOH6HhOXuLo/RlJnxmtSBljZc6fwTHFGbV2foF
+NOpPDQdVCk3cTm5Qs2T4EDbY6ieuqQHn44rXxPOxQxia/ciq93N4/b4Zh2R
rUMBgIh9A3iyG6eD/JMC7RuqderiQNDcEkoI/mJ1Gyt3LD9BTmoCCT4GgePC
9G8H5xej4zy2N8CBFckea8FkgedjSSI01s61i6VP3jHZ+7DsNsAdipzpgGmH
rnCdF4rTWJRgtPFrmdBl7j/KwvyCqJqorWkQl+UuzImkHtRPyW1CfY1qz22m
x9gX6XgYQEr8H79zxHtixSOOqFY/Yo0TA9QEvanZAUjbA7BRHFZApAlgWBEE
zR6SYscFvwK8VXhETHXRgaGQFerNUlnhs/uJd7VG6R0EZQX0sMPifCU5X0zi
Va/QW27T75nbsLQOCQ10MrATtC5yE5giVa5CVZuJDWwdmMAvTcncR3OIrJIw
RChjCN36DGklegk3VS/PxaHowmVH8i3oQgHeyObyrk3ntpLrwyObCcilvPa4
AC34oeyS9N+h1spDjAcgz0luE0TT7j4moYWQyr4oz4HXYMLrAlokPik71wYI
vSfQUq63uj1aid+GCqLKjtbcZqBlezdX6ftLW+EC9CsgcWlZgC2zXEAG6QJf
BnnKWoeZckoM302mlNK5ObA3Uqz2vx5PzWd2M/nJVZ2B+Y41/ZCVHN8L/zXP
NpDL2HGTQHyZQZg2Zk23Oulro1pPkVFzsTWB57x72mIMSIizwjHtMTWSbj+T
+fPH2M3YtA6Z5EeevI4qNagaC/qOqjwHYfWdU/TAlAb4HvnpvqvC5DY07JnQ
3enY6ewG1VPx7cYSNagrOQmG32u2PcP3uWY2/gckhA6WGJjB+ng4g2vZJmI1
lws/YiYM9vwGbd/a2ySDjvBYixEpn0H8UU6uHs9PBimgc8hleOMa/9cPptsA
aipl1z3b1U8WSfkGJSOpAWRYG7VfScJ/EoMVZ48hrgEGc667uUN2Bxp3mGn7
JLQXEL370fNygrbEgVOEC+CGbb4W8MYMnzkXV1VYCkXN3sZJfJM2yd34aTAk
adjZGffrz6o8LUvYIEwFeabO2IYC/dFYn1v/9n0omHDbhAGS2a1jkZqo9Kmd
1AbD9HGZPMl0RfM5wR5c4NYn232bj31rUKLYkmwbSKDjmok48ETIt3oI75y3
hkgBlYU28uavQ0iZowb0xuSN4gDH9r7EvToagjZ2z24Sj7dU4WfKUm55PUNa
W/HtPQf1VDxWixbvNswrKWfWuLd/i9c5PboBsT9lv5NQXSw17pRRHvgKZl+J
59dT5mjxzm1w4USC09L9fR81NbB6XbVxv80kexUrd0E/oaGZU4AXzMUvhQqo
V4IzWB61HYtTBHO8Geyf6GbCalgmLgz9O4JLe0QWAyYS29Z/mpCrfG+9bhlp
1+0bz5Ef7pQHZ0XOmKtL3YdfdOKce85QmFPZoNoZ4X+ChnqIkt+YlYu/tMrN
mySW5jjJ5uGZ1FzivIzBAMkhVZ5P3f5ANQQTg0PGFRhYWjjak2FrsfbGfBc9
pjo6ze3dGv86FlZ7yRu4NF5wx9aXMNvWjF0U6i8dbU+3kcDiIGEK8dxolu+u
uW85VM1sTDMl05u7021lShQMMS51mfq8zuqK49P5MvUkyvDfFtF6UJtrt7Lv
iiW/HbAEKJqewIujl5qsB0cnDTca5Z/Bu8FaBWaHVe2gNK+CbWqzm7c3wc1/
XZIKBxj8yYaq8nvciaDCld1QcI/SEhfkM4xCJGee9sMelVivL/lWWg9+9E08
LJ5DqqUMvD8SEPfGcuKpTX02QsEu8qVnv5e6IM7uKNG5Y3LgokAkZbXwHMl1
zQwcccoBgy6oSrWu9Xl8oHGz7ZxfK50QCMtYj62jVP5Kjjx55z2xkn8WbtFp
SrkgSt3YeOcNy0uzwI0UwT4+XiPyb3qM1MUoTFBaMOKShJVpr0+01Bp0QhKO
kGrJ1oBpwcvtALcpxqLWRRYL1VM/MGleo7jRDQAyiyBdA1xhAmW6LWYB1K2b
3sLX8X/hF0ipLrkZDNzuYepnTskm1aFbVYehqZLhgZFhA6x5EtOZdHF03OAo
H//fjTFhgQw6wGp2h3mOdUVruKu/n2918FykiNvpmeQDGDdmT62Nrp+vyEeJ
21zsKZXaNllH1H0H8cKDvz45000j1WMFxRAh+cIh6/LIF4y5nJT9HgyjS+iA
N/ocMEO+3tNXU3hgsOdTGEuqpwWQLzkmgC/p6PIA60zCC85oFozJ1uvOJfEo
WsCdW4wWcqBPZjaHfejJIufX2231UMp6j2xKQD/Rm+6+V7iOA82Qh6MqEQXB
IbUYiLrqKcWJUb1WVFGDOa817u9Tehq83NiA/QRzIpqUGywYCQFFXPCIRKZY
3qnoELpZpBy11dHowIfww7Sg6PAygkR98jVzx3g4QZDR7kWqqCnKxsjG5tmf
7MNrJa6P22soDzHh5Xn37bzXNOhODqXC+cICViD1gILm1fCvbiVj8IMWbN+a
psqQoDM0cPBOvdEPqPJ10SqevdFh7ig3So3jfVxM3em3Zz1mCNx8PZKRkgep
ZN1GBDqlHzOYEk12Cxi2vkXRS0MKwJzzNQtX2gwBak+JTG6iTO9yacz2Mr0z
BMW5a2HSZAWf+3Gmm5GE69+fHlR1qCsxqXnlooBdyOCmLHYBB/mhgWGhmwp0
3/Ih5hxbA0aE1/iBSJTX9HZ2vDXfFbHYqPVv9xwyPMEaS8j+X5hlcDrFznta
Aqyxyvhd+0K2VwKxPUtsCYKr9lINL5bX1QyZn0f5ePZ1rGTiH9onkY3nxQ++
R14ptdFGJbeZVS8Z5d2CYWLahQ256PYQWinSTcVGuWMCubbt2Zdv28f/k2TD
DfH5zp4TYlEjLha4rXfs3aN2HU1y6+muEMn+3qo1qNPr0qTaKVBtFFoRNmHC
n/SzrwC8JsVlJ7laHf9RSVvs9JKz9sDNKyw5PTYPMozQ3zAliBqMCr2tzJJ6
IN6J3QJEF6w3cQAI87b/Qyxxru0LRPi8BFkBYon2IWRAy6FPzk97j6IPNUkH
RsfLSxh1MUN2yTpiVFr3oT2uSCIyzf9UK66pFdKsEDwVj1jsGWIlVnp8UfH2
N2oxjXcVq1ZYq9mdHJ/9G8dqtpBEJNa3D+QyekZbRWxz6rmm9S74Fkze3Fym
2+MLo0aCRlWGD2CV3094cpUXJLeOF2Y8QN42Syx/wv23A5tp5a4s630IEtgI
tJFqUtnhLkbVyUAQ4nZEZflASD9ntX/4RPUiLlCap4ug3Vj1p0PEou5Ms1W/
Jfg+N8RKz9S7oOOxP30YlhDkxR0vq/jQ2fr0lV47Ls2gHhtv8zBoxeGY6WCU
GLgzxbeILQNKTqtVRbtM41YqFL8TvlbxEKwU0AWDlCJwS929mwzxMiIeU0LK
1BiGJEFjPovL9SfmVkv/F0VbJi8nLvjjpWKcMCKOtgM8g2ENy+aHo9bswJZ6
cSbnaDVKme+a4WFPPyxkYOVEVIxveJLb/KKFVhaJDyDW3LC076N6qnyT7qOO
Tmr3yS8FVN6B4XK7Bb34Dh/aYg5D7TU54w2TaUf1c4Zr90Fhp5pXeLoGswzJ
Kmd103hpHpvxACkx1byGBJ1knjp68lizBAvlKTrzqU4Q0XXJ02GNuZqXGqH9
FEICpgZxu83lvMOo0dfDtvpi389rLQpYNlsKXfY8b6yAp3xUtzblJ06VuYBu
QbbhcoKw9xlyFKXD9HCXOoygAeBbZoINbpVQWiSE+vxwiF4kl5aNT55yx8q4
XRTUuqF+MEvBLYJCDzT/TzlCcpoi33tgvgZ9IJehAva2pj639UyzmIaT360M
mG7tREmY476/UlsV7i1x+1ZBbJ/ZphpPk3WJEF49DLoTPM5l1QFxoMSWX6aS
XeaFOFfpMLoprd32RGxBz3Z1XFUaHC79lMy9n5ffKRjKCCusH8HPmNuYGkg6
fgS68KVm9ap6eFPnVg5MMm4aklDC4e0OoTcK1AWPBQ5ebTE//vmMOEJ2K7k0
8T7O+jWPQ4Ln0i4peAqS4rFY5fRvUHFDGqhQT5GAAD2jf/JteTUCmdr4ElnG
Hl38/veeoVVzvKCdbaw5IWyoO4U+wejklFobZhM/9dsI31/z7Wy36qrM7LKA
VP9xj3Kivdr7ivEKPk0nCeyFR3e2BuhLxpSyM3fSVtsl0GobvDIuGhDC5NRe
puj2bUHihlSlnCW/cR4nGgid+xym7OezrCV+es3HZDmKME0mbfql/3LBitQH
hQvvOBeZQ77556rpLJOAQulN2NAZknvA2j3Z/CfVbfdOXobpCVUB6Bvww9oL
1rsY3OkkHR1Yk8lhgp1+ijigI5MCB18BDC4c2Qv1b9NhAkGB1pk+2n8r6ZPG
uNqXcseKy+FOUoFudw5oGx92Q8gKqztK5nSN4B8leZHZIhwUnpY52O+iWsQ0
Z/vIuWACjYDF0s5JG+4JLyL79v7iOHz+5f7zKBFDY5Ud+2nC+bioImx3cw+t
p0yTkxl+gzSHq1JfKU0XttEiFoll4EHnbJEwCAfi1/q7jn3uInlH3UHP4owg
RzzFkaYxy21SRDsxMAfWhQ1t7YbLeTgjkReGhxuE+RC99lQE3kU6hV7l9/8W
xntaxmdYQ6lowFoVOIHJGtr4fAqEgIUotjLdrQsTkAHCTaOl1LaSCF+hH+IE
q3YwLOOC1ssEJFYRYHcIRjepn3KeHwkcdcCXyJPXEYWEWMkvvbX0/qqf+K2s
JUUpRztUW4Pmk6lpTCjaoGFFp8f2owT3cs1NckKfVgxpRFFStgTSIwhXvRwl
L9Q79Ib2GPHNuYdcFtcLU/p8UKh0JmX5yrUs1xN1e6UwyOldaUuX8hR/Czg7
DVCn7xTsUJqvyEDhMOr1KQyWdTGf5EXpyGq6lJGYQojuvQ0d2HJ/vSb4OkXA
0rMY6/HvNadklI5GdrFGcJ+CtQO8h6si/QpSoQImz+9sRtZOCxaijiJrJ1bD
PFM8FrtmdgwBJgRRqaLS//tKVgUVioljQ1z+BODXUbjZoP3RlMfLpaGuwfDP
QUE3e25xbOhTUJaF9dGD8E/c/LaBq9rsSipAyh6o2KTz6wa7WPrk0DrkCCz/
nVypthB1NdjKOlwybmaucZIPn5KQS8ZSjx7iBJOWDb7ddjs9sw98iMEw+qB9
EOn64xVJojxgndkqbFYlCcLYpeRmN1R0iwbFKI9v4VO6ETQ3LxZSEYH6taPq
jWCGmRdwPWy2R/A/HMw+EeklCBsQIGeGYSUuEeLiUG59jcLalEcORHxQzwQ3
WaimMkl88kR8rgAmV83asLkPQb5Ll55Bqnz65caST5jaI8HsAo/88VwkOOfC
trPQXQV8WoG0v8CxOAbzPcDUsuTOf8JaRLjuFCBImJ8mN57bXrTMkCENotBk
on3s8CDSKuC2NctehXQ5D5E1rmxqOj6Vm5RyUbYgOa/dZrpfz9IGsXc1LdRw
7ZJ7v42ClYfTp1M8rmq6QMFd4PI4bu8FDQCKipFtMq/p1mfqiitA883Vz+D8
QvhFhtkkHN61NB+ihpqr7ev0g/hU8MrtnLuK7qhV/kL5A3+wXVFEyYVcyihZ
IrpDLnL1cBB/WSfcdOhJfKk3zqEy40vdMshU1M8ppwGBE4KflN++RfuoL+cP
DKbDArMcq4xG0nmjs+YdzFkW8pfUbRbzajPINL05w5vYRIdSr+jCHIfxH3FL
kptfv/a9mXGAspvalZEMJ5sR0lEstAufxihWSm0YMreujILcSv17l6XoKGGT
NQ6sq7hl+y0qf15KAsURZs4tInhc1fdnBumMl0RwCnYvCCpJk5CFkM50rciI
WJdkiAhMDN80iywO9p2i9bZpFXd5+EEC2KhObsf3D+KeX+x0T5nPZo6oN8Ty
k6eYMfr4ZkJD5UlFgHQqJf1uRJrhDnysGLpcltDi27PTWOcM9bE6aWm5d/J7
j6Tjt5CHlRLEMCV7JGIfC2hE1qmamyiGRSep05+xK2RzATAyIrjb2c9cP7XJ
V8P47Wys67a1EjhF5vMET5J6jIaGtW44l55ydP9ZuiU6sgI1JsM4CpDsf4dm
uJyJ+VggS5f/D/8XACNZrvx301KCyvumHzhM1aeqqUSZkWkrMmPMxJzW5kIc
BQkFEyaDiOxlrL4Axtf0w1Of1T91f3Q6Ei1KrVR947iSg3CPk3VGPQD5q0Ce
Jo4++loSytohJKFSU07QjpOotO1/HiWeTwPwe10DzwdPzVYhkaoSo5krJCJi
9jkkyJT4ClNlyT1CTLdOpJKm+Ci4t70iiU7MF7mfJ1kiErf4L3Yzb2JAGWsB
BqLMRd8bCVNpTGytPFQBc/7/esNkPlUzbpfnVRiBHWe+9McxzOL8Z+k5NS7W
nqyhQiX9xY1m/PuLyFf3g1c3W/rkl/jkL6AHWaIU9jLi1cqZZu5MgbCythlA
1dn6knEPFZ902R5jyBm9jTfMFhcgyuaczvOn/leRck04aWNYRT+Pt41UOb/3
dnH2Q9njDkv4wVFRPRztLMrwjIg+HI00OMBlSrRqXMTbvBVgwnksJvH9kCw0
IprL+K+RMcR3cI2i8k8kqwl9HoT+28UBUN0/jKsdpcu28+Sce/f9gNQOAfNF
IACKzlS/vC4dnJDFH9wCz8W3EPXOR0tKeveEfk4k05jX2sOkIDWe0od7H+kc
pPNznyUuWjkn+ckWd0bUbQF6DDWCXID1S/dYeQlfOfNmmVCGWqqc7DKlf0fV
1NJfTlStFbMU4JgvuXHsW7iWNKuzpIleKOIIhP40Wp/PoDGb2IT242RVVCk7
oB0nl99kDkvpqWNCMuDEIp6kcjeigrYjN7fe8faaU+ih2B7zMQz3m46dlnMC
qM3UIqm/UM+j4KDN4tNb4pEjsV44YdlghqOhf9QMj4tYv2+uuXhaOMtLg1gM
9V3TeS+wMQpomfL0hFH9JQrnNgRprepJlblv4l3II6N8kadXEh2FfSOSeHp1
0ioiCseNfZkjkfJuT+DIyNJ+Bphq1/QCHidamD2QZX942NnXN1dEjMwKuspw
co5OE/rpy7BiMrVC9QGQQT26lGDI9OF67XGgZ9iBb2qmvo67/Nc0CDUcj3Vl
ROnNEGsgG6dnm7mA7GrgE9Sh2m2OflpPTqsHJqHN75WRSFYCnMWo74GJltgi
XSl87WV8V03fXGLN8FIqv/sX5chLgxBT3VJIKSh2/F4NBx+CmTVmAxikfzYB
n+ds2r4XR6ghZdf8WnlH2gzk2lPFZkWRnsnWx0QpK6v4UXnrInYcJ67tkwTk
YVDyFbUed2yewtHs4q0KI+oysfswMswXRvnxbPWqN524+x6/fOgvkE9H2gKr
EGE6zmNBTaIRYjGu4vi5DaY3pnUllz0PaETi7z865Br1tVbJyDC9n42JxzLX
lFOdosALb9rA/073B51X7ucnJu4CCI1nc4OhFlZp4XX0k8hAM0qsTPMSB9rw
9bKF5dcX0MH4KAMk7qhVZhPZhV0Tuzb6tAXxxpRLtmY/CH7I1mI2paNQV/C0
Hm/CdERE46+zaTTbloSqklOS1MgKMCmEYof68rfI4gCm2ClpInJsCCmSHwSt
ms+jNCdgv/kiXBoIohtXgEMDe/SmjGSwWHjaDq/NrCPCkXt9Uv3u0RBiwiqA
kcMRUtwtp+DQDO1/fRo7XezuKipGUBSxYTEWoFIN+wTBS1yjxYv/T9FHUMUo
hBcm8ck+IAavvT9vUzXS3r20INbpgNypA6RrlubD1iK9z/TCZOgah9/ujn0t
+PRSZxzNhKXhLZld86Xv2GUJ0suuAfUG7UW+f3KEKe1oWCMSkCj70wBnOXLj
7Gqhfnd1agirTYmSAF6SEiC7Luu7k3i/08ERKUv/dGrjuUcdeEfo/dtbL8qA
qiuTKXbdysLfI8VUTF3EZuZc8csAszarsL5a7HiL6MyWwokDbk17ZdxE8oMI
oqkeEBEFWmhnJqHO05GyVWkTLjIusakK3cplKn41DNlBwr7KGw99Ng3u+PI1
7UfCoN2zd/1Foqkz1cKVDB6GdqCU4dCcW5jMD5bXowxqsMy4/KMloh3ayNFi
3NaNFOkuDs9DtfcH5tAA8f4/T4r6PsFEjonhPr8h+GUfVFM5g1oXeLbXhQKL
B1OerHtNqQ4Bn5XatOkDDKpRAO6+Vdlm0bdG2aya585C6Zqjxz7kKOvtBaov
gtPtA3Z525R0hBElNDrDehhxJUYc+R5HmcM1QVOoturuKItx8crmsJ+5wbJk
LQNTWnS6rXlFBJo8FXkNXBVt037dppvjGQcnibiQxggEbn9UP3PANHEjznjY
1M+Ag6LHRFRDfFLzv9NoCTZX2WQDz4+DlLlEtMmCpU7Mstck6P3FEe8lZABX
J6wyVfs9QVtAl8ThBi8vm9t78Pw5bYiUS/GEbMMRFXbaF7nAq3+JSpGo2HRT
AynjD3iFv5Wmilr96QzydZL7QivONP9TdoSHBwPYmLiOdODeRIR8tAlFORPF
elhk0fnQMfBOoSFTgcoyYO9Kk9Myt57ZCef/ULbnp0/Gg4Da4Fd1bM0/Ey4p
pG1Jh3yOJmzH7C2pAYIY0B+CYlDdMV6/094xoVLEGAdNkA7SUdf1NBePP2Cc
njAhsW5TYmPJ+Y2uXnH7H8CnGuRa8YdvZFs7xRK0ODUbgJ9Z0ujevL/FmeB9
nXEF8KBfEBsjRI/0cBYb2BFpFTPhWfsB7t3cipyBS4ZEPDOjPXAxtbme9p+b
k49J1/kwXacRMbP+CSTvhJN1vtmgzQSjWHPpVwv1rdZCAiedTU2pGJb4CV8V
wPvjzlwjDxT/mBOXJ0SW9o7Oni9WwckRBJ6ZIZwpDJRGSNpa5+5mCBEIZVPw
ePCNeyN9Pto6bhHNzU7rjRWhAln2pZr0+8yOPEJgqoK/hscNbugk4SNCY4wj
vsLGvV00xQQvTVbXfvI0f2EwT0fyEaK4nSHuapi4J58O+zUUTxoeiSqNIcls
93Cy4MkqLvR8I1R27oP4S9GYbeiJdr9Krd+gZWSVziYfiZBSiJoB1bsjpFxH
SIbtBvXORtwdZoZGYplQUaKwBogkzIFgIwdHO6p+c7JxiXL11vFTGgja1hHl
ZsRnzXI+dxqpDoGxgIFaeDc6/NxrMU70FJevQlqfGTRvuJhH8lh3aIrk/WDs
bMllTu/c8VxTnomhHLJiDfjO7hx5bH0qh61hOB93o+TbutMN1zK9jAUWNPZW
ARDyOJ3pcy/oomIBPZZRJsjk9HXh96vfAZiUB5Rx4n11oIYse4QgW+p076xZ
isPFcNkrsNGO/0IPohCnn6pKQDnGIdgKF4uk2UhUo9c1wrF8hjOwmBTZDF0x
yAuTjiiqelX5ssj5ABpSFw/DBTu06E9XxN+VnUqfnOuaxP6wfKw9PHo5CYDo
ncG0tnGQT7hmFBNzevQcdvTpvOjdd0S1nVgb8AMAdi+uwv5csIh4l/BWgQDa
gBPa8y8YMgqOWmsbHDqquG2dLkINKN0wOCPnvveEcy3EwNLR5WMaBr8VtbGN
2rwQJpHcsbZ0yKk4ptwcH7x0WC8ApRWhJbUh60GtYrBB1sRmGiDOEErKYKJ+
hkoaO8J/y8cEijS8X1fNytED5EsXurmoESoJt+AeBadR0av9GyZeg4OY7fcj
t4fTbMrt8WQhkxwCAypoeB3CipVBkeRl44jzSPeeLR4vWFVfrWhrC/CYV6wC
dZ5IbXjbW9IheFgK8XlSihMu3AbZdIKeKH0RsjJWO/c4jVZFH652VAip7u0N
kgMVfcgKCQpVzYklrCGO9q7NQz3WJmwHj2WjfbWuyu8VJ6waf5g1RxVEixht
0aRi8bpAhGjmVoUqQaiyzvsgjPnY7nMF3SZZ5LBylyUmFGodCRKpcO4rxq+l
83YBDlrEM796XxLSvnw6RI2pSBcci7plSFsqtsQDLw+towKs1ft1y5VtTt2Y
ZZSYgNyCTybAf4MQoqMua0STuzLUgwtqpEbc4YLTErJrBOpVGilwpx1yL6HR
uUSRCutz8iPjUbio34QqLFMtpztVVwJ8nBCaHemRIakSApKwt2ps5uGCb6oa
QjfENrUPdT/s+P0TxVXECb2a1w8HGwafvB6pO2lFXB06leKsTYPgehC0Lbdv
DRBuaWH621pW0zSYJRwMk/pknSLAbQji9YMP+Nt8ztUjFte0tOQP1tuU3vDm
Zexv4pOZueWnPgM/FNkKxErY8PdZ1L7P+GdXxC0t1On9nDwcbQjXIKHzVxSw
UlGej8+MltdxXK9o9+K6RWctKqwS5ff8IwfEM4E1vC/VosgkA/eydj2lhM3t
Z8X3bD38QzMNnfmGgovxQsGjF2CPBAHoTrP6I76XtYZTywwYnapkzvJmQGv9
u9Kp3z8seemVCRZotc9GQPIoF7u1Jh3m5hLo6mrG5c9Bqua5J0MTYFEydrgV
iFhEftj9A1I2TNQpzBqC9J/HF62vir2B8kahYxrZ2HZ059aOxgZ21EDoGuXR
TpgRWpS4VmPGF2ogaEggiTX77yWeQSUNXuE4GsSODRszvGIsxGXCe7PE893O
EZ6WTZKu0FKHAQ/+SXZkuNhDJb0CiOLNgZLQ2KvqIiAhz8RS4R04wH/NVIYg
3GejZahqWhOj9/xuni25jl2XiwST6v8OejmvZK/BYvapuv0p/BdUAxRhWbNx
XIjmfmS//9OhQLHZkdjAGmo6WPeN7MHhE7rNsghKoKYnuORRqljQbDSwVLsS
o2ZXCe3M2k6BC77FKLhe8nRPYTxAdRF+jqUd0OSqSIS4HX+UI7+NmqrByFCh
AUs7Fbs1uULMRubPmx+19l/653Jggd+oDBWrgOo6c09dIUpuOtLTZAuXT6qH
vy0v9+mBJ/HSqx+xqa9J5sgp1LaG5X5JkYGXGVDMFzSArhtWVnJ/HTMg+Rx/
XLUzaf0ETJaHL4Td+aMtVmWrB1ttrg3sgt2+P08s8rgMlyeb5lbjfNhKFazA
MIZuO3OipJyhpCoL86eJlRvDP+V5rAwH76CWUekjJ5ed5FD3ERXn0VlHqUNv
TJKiLGtL8CP/4ASyvAFRBE76XAmowTMnrn5H1NT7XBvOESRp0ZrcvY0i4IsP
S9samqyDPqH5lNNXrGzyTobPo0ZowyyXsmIIFZTeY2ToI1Y+wTNJ3+q/h+sg
ATKnB4E5PKqKOfGbjZeeby1qyU5655o3XURfw28Pt6fYRoz0UVAmEWctFtSK
L4MRCi3dvrgj1cmsYoAku1v53Owp+u/Cd1soX/rqic3qEsOCnrXsa9VGMkny
d5ZccC2aL7EkawcqNTnF/01mA6ylSImDkkz0JnzAI8dw6pCIjJ13zAF8yDsh
9oHAXwE3b/IdxoDG8ngqaAA2Z2ijsi3H0m9+S/BvuN3naLJrMG0sBc5cVGgG
5V07Xo7/STt0pKXYFrjjhpucLGzWblG2s8R+T8W3HIyBh96fGD2F5D7nPUkH
JbDQZTFGlzpQpwnSjTBNBquDmF6zHoA+tUfnr8dspmRMk8CgOQxvsxPMRAyM
5iacwtuZ8IGApmMn7sKxdpdUeWKKIb6kruE01Sws3H7pd/I6oKVTSUk0YDit
xvFh6Kkr5saR7FmL4o1YMkmjY18UBl3SiTZaD5ahNZRCYIIz0qHQiggqPX4a
BL2Mf2iYzFkAMbd9teM80lT/MyVO3f9OnSM7TL1PmYcHWgajR0yreF66yr8N
GVZlUpM1FobhPXsJFffmCbZrPS6g/W4xrpDIe2QuybVE5eT+eU2Sf14gBUT5
5IwmcAzc+n5rom/oK9NeB235DH3XZE2nX9SVE8LyQ8pekbbFUAtmoTJurnWv
i+mPxjIISkwKEqaKTz2MLfmyaF2oOkc+y5h7joqzzBRVeqRHDeoNz6iLT3sI
vUnT69GKoBO1kj38jsN/j4SwlgALl1p8TWMs7kCpUuwzWLQoZWBKSwIYAq8D
9tgP1gsjAV9JCVc3qA8yaPR73oHEZR68+uNeMCS+SqZ0+0aWUf2eHqio2p3D
px8uolcfsCj4cSXmys5wmeK2o3/qPPufvWa2gPhqGaemwyODtPkLHrrGlFsW
t4drLXCMHjm11wNJD/E+5ofSeAFj1UhVOljbXJv4NQnvX9jqQLouou6QliQj
cokHvTcrZdPIGBL9BUT7tHCPieeHCGRy7poAM/dzqcXG+p/6GHFUoY1598/f
o67t3txfsgDFPUJ/xpfAP2FF57KHOfi/vj9uKESSHxOqafMEPhOKB7YYAzEK
qMkGza3iR4KyQ1pyHPdzXZ9DzDBKGFdzDyeQP1fTxTPQ4neSnAu4Ri1IUMJz
QlSSXYK0l18kNez1ysegEMVlz8dSLbbuwW209P3lf2BBRZNRGIng/azSdotz
JbHfRAQMS3CtSSybPm2H6/Xsi+NQ9IqFcA6oQKfjRmduvvwzz06B9K1b2ARS
AhCfaBTpf1AMKUdqRq6ugxmy73Lb5qNkuOn+F2QIo/jdn2ql8rInWCxPti60
F2Sqg2NqONqwAxBTFREQxubkZEsb85Om/j/BzCjGj4BxZYcpMGSrkqHSgK/V
B8mBLjLlFtvCMUMDdtVgNO7aD6ondBvqqtzYiGfD7JLJ3fzhbZ4p0tgnDAGA
PWZmfxy1pf+uRTUJ1xgBt3CMMspaqqIJCdQMSp1TYl/o+DGZQGJ0XoIS67Tm
Ie8CBOIpXtQ4tFARls//77BI1Qo2VC4riqeWh6I48osjJzsTf9JMmOpaLk/g
Qkm324PffwLQTG5xmVZToWsEMkyuOiFTo2iMiu2A+NDd6jzcyU8adM0ozO/e
CvjhziexbG3VQr8yFb3M/B8abqJHb9eySEA2RjfDZK3U5/62Aenxjp+ybG7x
pleyaPGCEwYhKZij+qfmcWe2H5K+WnuI0V2RmTNZObtjAogrnxuMV9nQATcE
nEUgLlxcBcmBrnjL3cBOuYUYnK3QN/b86SWRVlqPARJy/J6bIhk1izZ+ytDg
jxDo6zVdGQ5mEG6OolGU7q9SO1b4lS5L3Slj+wzoKh4eENDXKnD0A50fq+gi
CdmGRQJtx7d6mhr1eUObEA/Shm1HmqmHODwFO8hqXWAmCAFwkSgMCVMNj+je
qZmGloho6ZFZ+pKbbHijRGTGqPmDU8d6EqY9MX9f6/Ijt8NDRuifIcW+eCyH
EZGo3gBIv7Jaa7MbnIxQzDOoDuvdUq2LF9bWcEhryerlsv0taYX42Io+0RZF
kOuwfGBWT/F5eH0gmMLE5zUCOlErT52p3PKP63oXVT15WsEdgVGNZQinbSLR
+98EYO0KiULDGfDyk8MctpDTAVddrfhlLbnxFtSR7JI4VatGm0C7jsLS4kEB
q6AXwsewm7e+so9vXngfTZxcOQ6Hlc/eSV7fSQ/Dh+6hjPyJ9975xdYc9spt
piS26xhfZDeBtq5GboQbKLTvsTwPLu6iYkaxHOJu4nn0BkhWrvTu+JBF+I6P
tl7Qhn/hpBxdJTNabTofBKdjMUMPcjKL8uxMNJ6aA2tmOxPsttn6g2o3zLWm
u8Br/SCxJ4G6K2+tmaM64GEQsOJqDaxbCESsmFOtsmh0JWSM2GtqOSQwBFwv
kglTNUAN8sLMooX8vcnaNb61mc5Xdnq+mcg4+RsVF0+ZUx1l+KbCw9B3CtDQ
u5e/MFnP9137zr642t88EsFniFHmU3tJxcLvPFw/QVGqbCuPzrL58THohkf+
/rono+yd/LpLTY13771ZY7DzxqgutITi8CDrn/YuqET54jyPAmAvxNFkBXoq
vu0HIx7AQwt0XDED8VRFCrfI4ItjpBYJcalX+39cLsiciT887QRy/YZxDxEa
pLz9nqeF8JppflRNRPPMbQzCzgdHGXanpeDQB0nRd9oNIro1awfOED1oapS2
+mUDda02YlvkUpGeAI7WW3I1xXCWoPXuJJQZcijVkTRAnMMTmMhC+UNTEEcS
8Hb/RBHjCHpox+x9ZUYiNV8KO9pZPNyyxfee/gM3S2BiDo1zjY8UWLf56YNx
m0v92NSmvuG6gC3IERtBJNUZ+TP+Sq4BrRRU7i6KL+CRSvn8gz+/eaz3kua+
pg+pAKArjW76BcwOC0r2wOwZM4I/b5Cg+Xzgy1lV1UxCbMiHaSqUcrhP148V
Fo2C3XqihFjb/afLV86ztvQFSsacxMN2bPGKQA+yfPh0/HJbGxgi3sy7RMQC
7BqHGyNVrfyRxN6G4LObbccstSZWwdCiQuTcKjwPPCZ2Pex47rxsPBHQJ9Ui
j/JBefu97IMSbOtqQA10eTT0s190WYif8kqmuisbnHuGQcK+pW2LKdk5WdF0
rtycZTM/jOl1EkrXhAFUIhc81K2lo73qljF1l4h+iDl0D3AHxaMxnBX1LmjE
ZIy8mCFY1aeBZRllku441gYpmHt10caRXhSdodLlrtxn/tzMx8bY4z/vCuK7
4wSp7GKB5wif5tRgqJMlwlDuFbhTQ+X6J539ry9YzHH6Syrde/D696fTgZrX
cYnA3VnzoXrIqpvvDlgzb6Mb3t2KjMB9nvyrjj8wdl7FNgAv7jIhefXEHulf
x8j1oVnD8G/r1Uh+GfZ3OvKryOLPq+uyXXUA7lE10zRcBBQFudLqcfgBt+3M
a+jLC0UJAITkHlrJZ4KvGBomy3lQdqmBR1zMlZkOsUoOGPXOlV+/jC2k4Fo7
0o1RLgf7Yycs1+GgNcbo0f4KZJaxzKuoAzmlcb7oLStXNKWF8UusqrdirQLY
fVT6E4uK4JMgVP2Q9aBRrXg6I+8glw20l3a2KWXCQqEfWf6MPHTYcJVY0xXx
i6cRnvQFFweJ9LW0nyo0hCTeLWjQYvxDy7ESf5LaeboivNV78DrEEeiGKa5x
Z+BZLezrSjqULYxf1yRfQCylpQYsG9jgB68PPpwniPbdU0ryh6DTHGGTUQVb
PSdrbpswDNY/gSuvyLbztaPd1rBPNwQzpLphuyTg0Wz+oQTSmBP6MyF0Dbjh
obv+vMLdJPNAKGNhFg+JMZnspcCmyfqWZoAExU0JPBSZ2hVuhAummUjTm+A5
oDHuOpGKNZpcA6k2VYaWMFpRufMHhJ3rvTBnhXnoh5STPVs6Mw8qFxWXFYJ3
etKf+yeVTo/mrKzKZyNcFWD18mtufHC92YzxBH3SWocVskY0WqYY6oomGu4C
4l5+Cs10gnaLeXNzUUuYp2ned1h2+orZKSExOY0g+0NV9bwgm3acBClBsowo
bAuL61GwJjGDCJswTjce6eCp+b8OKXeyAkc9CdCc19ifSlMXyAKJs/x1GMbZ
B6U4/qN/OIWjBoyIt/aulMk09I37R8+xfOvWw1IVST60ScOlAg9QkzzrMeBJ
tzFw3eu4UI1g/O5jAlWZAITqTh9axFOfldKV5nbYajI10IBT+gThVCVgkjr8
Z4ghJRp8wqdzf9ucCBVD3xsU+aB49jz2we3JCVA/+hNFNlf53zoHT5UYcCF7
mKKRczrRFItWS6LrAp+ABIOX2vLQ8QHAVlAPkfQH7rPq9ARLWm97utfKkXU8
VpsfRRuigfTMUQElROYaE8Q2nvEB6DmAOLYwGtR/mQXjHv0rSNKQqFoJSk9N
OKCE1T/eQQTM7UStfc2LkBDQIeZ86f73E8oT56QMiQV3WGWL3SCadZSe/CZk
PEIFDWHz3cTKgLs+9w1l081h5QZw0fsPRIPU8Cz94288jJuQ+81YR7ZlS7tY
CD+2bvsMhxfO7DcMO9+1yM32PFgHhQkdtR450cOYI+wfNTitOIDJv14lMbu9
WHXiptidO+UkkhKFn5aatjAVM3429HHcy+wqUgKplOppa0+oiimW11seetMz
m4aRlZVVwH6PgwIm3YNdJ8isvrJsEt1ZJhL1ephTE2l3PM4OmcOKEmkpFi2c
kfjlfQEHZzYX+aFWnm+Jc7hjaGMWgOjja7izkl5U5rUJAadOdiHmzBK4EOxx
ri+OwUbewvgsWgwC9j51wmuneGfNz8GAbIvEakQGgxCLGVSttV01PlYaQkpT
dLWzMX1WuBt9A70t2EhDaMYs6MmGKdkocJzXgHRQbrFckK0mAwplAL2PH5TU
cJgkh1KdrNF0MLFYgFmTzRYo7t6nvzgmbB4a5wmXTV4fUhtHRFLGnR9mzTyf
n51oTjhIA3cy+C6pSQkMb7CZx2vJqzSS7mwO/ymWz56fEf1DGH/M50ImSTee
N+gxdneHuR0NusTKOh2jq/B4qs1skBenwIEa9eEF+tBfIksHvdnhyOLWWe2S
Kt/zK0nb8txcN3sjx1spRKDAGnqKX3KkZSVgRb7Uo0UyPp56t2HfqXeS/RP9
i4/736IwysP/TufCqMFhQb1IPYyknuVE+YgWoQGz8LV0l4z8jrJd7QWtDtd0
I2584B+ygax018e+mtAKyX3BKmvDSFW/ViqRigKSc2MrFVmgdEbpFxhfC3Bi
2qgkBRmMw24/RQxvvHqZSzjPqNLRZ8jbFJkOjzAaFrHKTf87ZO0xyicJBKBy
U6wwzuPtmOESIQg60EDcbNO8byVCvpaAH+DQAt+3qFJgTDvgafmTKKGX+peI
+O5ZicLVv6VDZqq4vyoz4r806WMHOAqfDozkdRuIc1OCbeFigxXkloMm41Zp
OE6zckKAl9kRoDOKld2RRC/bzqdkdjVc35ijPDU/rajKQeUyDGIJiu5tAAGF
air5g1UtZxBtSWaaZL9tJlSGliYO1SNuOD5rL3O6DIaHsxsiWpBogsnN3mD/
Uz6J5WYhILc4l9JCu4LGuUL/SbjnEg/VKxT+TtVHgrddoUcbIbIG7juBwIx9
9VQUQOKAf/+B6o2omAaxN7e8qsjdliAb8V+4kJVhlm4ejio9ARNCHWErx81h
LV141PPDHvkBmjtBcpkTeO0S2zAAQB7fKg9QNxq/axB1+Y+qwW60ttAddOWI
jEgDkd8qINlqy5CoKvf1ywSF4rI/aiaFl+5mq9eepwWjQ1ECUxECS+K1Dp1X
ISqREsAYpiN+FwFZuzA/pm5NwR1Nc8yJFaU/VOq1hNkV+QPuS5LYQrZ+spt9
cdRKLjEarOL27ETKBIFvQa4LXi3O03TvuBPZVgWppS8uBWnpEkjm/Aaybcfi
fIXnp0Cu7QfvkPgNpx2DgSbcTvG0JVI+UZlEPv4Hu3SAsIOs9lu8c+5mYMA2
r014UcQF0LCnPyq/w97tha8VRk2sJdMY5X0xTg8/1ynFgkZJW93Ncdl07qs4
LRRH7u1GwcxHZgH7fEzTHQqOzGd8CcuA6ESHMosQRTZD43MVQYjTSWMFgyth
4wbCQDaK3S6dSM2jglvJQ8+j6yesEBtiEwcCGPU52hmdNiDr8ImKNOPxqwyD
0auFfOeRS4jsGzMPvlj9hTXtta4gQ19mBqNzoqD2jw4teskpg2zVX8jjtffD
J1ehKEKzC820kopzoakzNWm663Rr9UUyHV2LWoJ7wOM8CZfBj78MSETjwv/d
dYpn/AA1UsLLjGSchiW0YU7LjDHyhGNuBlRqh1ZjrMnAb2/W/L9GVk4wA3O1
tereKoEcXN2aJyh1hF915S1dvxb5IpCmPro+OhTCx4DgflSPp+kvARC0oRxV
WH91pz0BCgAM/r8TNhIoHQYkcW9bESMgaUZgx3eArU48VHCZEb1eOTHALUfo
/byzQT0tw7VOZiywkJ7q3BVouwP8za5Kk7OxxSovb3gMrRy3W1r5D1Bu4KqR
F28Fi49J4uvcCkZjFBUcTEIiK10k7It2djZtashAsCMj3mGQWCrmwCkI5AAi
w0h1exYAtULCfIjCrPvCvbn+0c+5IHOhvHHeRbPPxwLOeTsABFGnugJ+Zo7v
atrXskzfDbMcdq0QoZBM1vGuRAP+VEj3HMcItrv9ikf9znXga1MUvPL3Vap8
RRbVWxwCkFy/acv9Vxx9bXgPcJnk/aUB8XrdP10FNKrWpXMxB1Fq+Bb/KOqS
WAzYFcmsU+Qn0NWZRX8mUtZq7vKd9LJb/tjIsUEJfPtBV2ux1JLfs23lpK4a
DyvY6d5DMC6yVaNAUgnDAJucEpwBGaHXwg4MFlv8dvg0UQXMu4T38UYLjCNL
WW9r6XI7wZnkT/+X+xTuAScOqyGa0mfMOQegvOAzy4dNB0pFLK17pPQ8HggU
CuOTHkyKp2VGMs/CHYdUjO7pwoRBTCv7P7hkNGMqiXIYCMvc85feiufSEIdM
2z7Y25w4N/MuOCrOpTOd0YSuWc7887C+B9x4+IVR/GRuKFMec0ce6Sat3Af3
K2xIXeuCRATS7MWkENTPJoraw/6u+zTLrJuWdXhdGMCWEaxDxOZNK3yKmYDq
nNmsvQnHGFiKbBPSvMHDOlYpI02rOWW+m7yt99wQ4RUY008dBkpfrpNUv4N0
vXii9ptTy7934KWvIbrZDX1rdex5yDXz/xfYmldl9jsF8axm2r8OzSV2JNdL
jCovRy1rz82kueRpom82ciD/iH9oeSy1eY/7i9V2eJKJaulbfPoBZYq3Jvdn
01lr1ENy+molB52JOX7wtBaQSyMbwe0FYw/JDeV0dPFueLo71j2e9Sudk+9V
22v3hUk6j6SckqKBk2pfHSVeMPPAs5Y7GE+bL6M53QNOIaJbm+aQZIYe0mBG
3ygnd5XDIO5kaZQxsHFfkK6zJSUS4595X537NtmuLG3HP+Samf7C/y9WvRy7
+3bBMYx6Uf7fZPM/KdzzZ+dkxu9Ht2d7+AEvM43L4zHepZe235HdaafUwC26
y2G6C339xiRSnWSV8kIHBm4aHfGLigSxLHutf+unUeFxuQPxFw9qrQzhgCig
+eu/ThbYfJE+LcbEATJNtzg7qle89XWgg1wS0S6sW4Av4lrU7xjTksReEBl5
0FlZYi58QwSW9DL4H+etgU/iJ9dvl+B53xE49AmIJfsOtcWLwAr4I7nMp5zd
xpfrqxWMf3JbxIhBBHzCZp4rAni2nAeFLhmT2eII9/LHGR/Cyqx0ZdAYu7bz
vA05Rwj4OfLwK2YawWFO1ZoJ2IbaXbTK04qcHneCpr0DMUs6FhHNiwOeoStO
Eqg+tIsaLuKv211zHBsxNzEm6CFX2+aB8SOUEPallQXPCR2EaQQsL5Ok7JI0
owW4X1YPKYUZAkBRn6R0cPf0EI/Ss2n0tYve5WqPQfXHZMWTlR/BOOcRAIMS
gdMQ7NV4lX9WkyrWBBs2IrOsO6ohyjkPx4DmrxBZ9t7i4pAJ+IM2aEjWbQTn
9fjAxbItFwddvz1rHiA/ER8T6u3FnR5v4LpGNpotOjj8OiO+yMQH20R1zufQ
Fhqv/7XITMvdMY/lA88fvjCO/D2SWjL1cFvTpILRUMfm3XdY4N074XyK+93v
FMHO2EzrACRdxYDr+wtS7ywXbJcV4b8O2iV79sk/V1Vd44S+7XHEADkGpQDu
XsuBDdAbxyHgyib7nVxk9FBrEde77HH+TgjYothCQVPH/EOpMjqLN+dJYKJ2
+um8D01Fb0AOMXfphFmMZSI5o4rXpoHSLFQ8iwMKwj24bFScMW2emUkIKKaU
dj+LYeBMiXFZnsPcJPu0Td+E+20io1VItbgmY9QV5H60xQAClmF0oKzJRNBa
R3iUzfpvhkcxEx7Ba9nogxu47COYQRRFBlhNEU43LiOLvYCEuP8Fr+v/Wd3a
XSlG70tLspvIs8PdAmP7lzbZ2DF0ZdjywBoZbfv0Q1oIRVYC8EEnCDzK1XrK
YLdtXJPN/hVQr4b2Gb3LqVnwBmA3NGIIPNVFjGwV8HpMfm9i0vvnxdxArXNI
/l8/DMNalR3En63DI3fkAhkGwqtZWV63bK8/s+Alf1L+FLXkL4X5j/Z8x28p
AllxxU3oGuc6B0RbNQmEfr5RsNUWXMoRF3scJYbaRBtO2TxeX3yLxjOCOaHA
iwP/TiNyHDqT0yJgOyAX0XQwgfVmbVmeGEqaIK+6Qb6EtLE8FvTE7n2UtQ6q
ThCh4Sf/NWPfqRoFkdxnCEtKAGbnKUdI1k9oZBqJmYIyRPc4vm6iTWUkQHDP
Hhc+CW/eeebcd74kGpOLvFOow6o/76v+87Wcovr/cv57hSrIqcGrtsL2BPPE
SNwWSKLC9wfdgnesFSEtvX9B8ONpf5kfj34BZhqlEqN/4ofJdOED1mCilkGo
p3qjoZQMsf3dhQXfd8ARfGsHf+3mnKMEXgkOK7u5hbjg6gIPpiarOznz6RwC
HKNsXfNcnUwSHfW1IOAglI9zwrQHhFz69Gjb+fDpE9xSIvah6337OgjFxKh8
CEuPFJ9RfEMgy6WWd1rc5PO8qNdAHhNF1UlrrCudba+ORZowiQecbAZi9Her
mO1WOLxRWjL8tko5vrN3bmOdDQyVosnjk/DbB23T+22MjlkBezq6U7TL6VXF
rm1ogJrKEMzauN9NqeseqMQKmctl+rT1Vzwt5VbLVVycUYiYwPqg+BgRYDFi
NowMjD/fU+TwB7IfSQBvRlDVF7df9LPCt1gnn1CQdpzc+2pcJ3vOJNXfUs2+
b6LAKPtPTi8vn83jgvP2sYX+oWaqtfhKuMHdBxUzP4lkr5nbZo4Rm9ie+y+2
HYheimd4f+fBM/ei8jl2HSFMIniX5M3LgJcYN1zlqwq5nPuMzbmV95Oh8c2o
S7wpbe+iSm5AMQoe2w/hMQqWfWG2UXOwDQ2j1NmWyyHAmq9f+SEx0lm87RB8
x/kjSEUKZXv59CENXAYnu8MVP7Ml3Csx2LtfAXOWxx8p5gaqkf2Kzr4XyjR0
ErBy7y13NoulyGV1wci6Uq3h4GxCjLpKJ5gLIXhbDu3pvW9lPEuMVTWan2YE
DoQ3TQoudr9RMMc1resmjiZJUNi41kN0yGAJQYl4ZU8RNAdHvQJQWI7zOnHw
nrZLq7zFOElMCzuOxlUCKhsWumFwn6MbEphmBYTrOI/mXmfWOrLEfDRDQThS
oYq8vjoq4Qkh8KYZme5xU4WpRqXcQxsqXHXerWY5bsGgV1I7MSuQwjDNUuwf
32VwBM4njYqYRCKpVEmA5A8eEGEoO5JvdSYLc+UgaWBd5rlIP642I9MDUALv
7XHsv5xAvOtOy7BrKmzngZECg25QtuSVOw3msiWaA9JVtm3Qcqfvv6ffJrcU
63dQFMwqEnSOVdUdklPyDuqBfOCYSlvHxB1iAmP7PTG+bPagxo9avsVmvu6/
1ibb/I07so9gXZvBw9VzOHsvpdbzx+SGpQqn5dRwuUH5dss9gs/RE6Ke6RZM
CCnKigdqRluedsXecE9VM+12H9OFXaJh6kQPyE88DhEpz8olL/g96E69KJC8
K+oAxRFyNa/okv/n6P5aWHNqgr3GAHDmseAwIWtus9XjzBuYw5fB81z3mlh0
Cbm55MlBsQ5fd6FidH/5R3y5EewA8I7npkT3TXEYLyMlRbA71zbBCwvexXhC
WxCptwYoH9zYjk4vlaisfWuhiFI9KzDw0/AVtmQy9N601wZumiYmWIRA0GbG
MkYiFBTKVlWyEhA50CsPtn6slh3+s31PSBbsHxWNrnlK8CVOxB0qPcBhxcel
xY8jU2oI4/eZCHSQakHSjBr+R+5ayhIV7e3iouv9G4Hw8RhTKUGGHznhiho1
ld8Vbs/+l7CjJlwejC45jiXTeHXeA9Entm0reX5LWRmqIImKvBia84NNVaKV
HiWxLy+zWQthD7VjXpyb1TJBfMlrAVs6EON6wZLQ91kW6FNlB1Yz4Sj9RZ68
n5VfAZsYUOCxsq7T+KaPDVLsbO8Rk7vEnHNGUdihg22tcPn0mJ8PTAApw/Kp
7A/UQRG+fShJHEXIkEbUeYQoV9+kxVy3C+vUgTwouH4HkR34/Zf0kQBkR3da
EJ6HYcEHvIBeg83oMN6FKFBRF9z/c7lE5ND8qnWVCX38powARZv3IsjFO9it
6UsUpn9wMKl+8ygaUSj2Q3VMx3DnqxoUc0xZSw2nmhJqRj4j5ycoRdGGuTxB
3IYpdM9byPm4KMDXjWlJBXTaZOaSNTmtYjKZuQimr5uDULoJf9Po4PFZWtkq
thaOizfhTTQPzossDM0L7JS9W198VYHjIf1L+kIkBbNPezJJIY4Uu2/e/8Bq
08CvEEkXpxNJvY9imfBvzk9Iprj7OYFcSbDb9mGY9lwRJEjh8WqoVIU65Jqo
LSRtTlK4/o2ca7unTbzyYfmk//EQpSekHFkPFSpvAh/B62n/qyBUgCFJcX5p
BrFVbXJtzuyGy0fZeOyk3FCw+nVbfG0T3LS+LgNnZffz5VlfWzMI1u+JRyoW
4YqValkXorr6j/zeh8+cL1FznjU6aAokybQezdA7CTS9UoTdSCniZY/+74CW
xgX5Zv6JN7TlB6ZBXQdsrQIRNiixCQXzxcuhBvJBlisKnriclr4hS4czyeLb
LWP/+6pI/EdpXmAws7xs++GjXps6Jy+etXSHCUPXapFQUErgsukBGvUvWzRe
fhG4d4bTa78KnXTUkbhsHFAQsN+gKRWKhOXH+P85VGvFeMEJEfLL4i26rCF1
BYr8tZ23cpS1G1nsbTMGMejy/30Ak6qEgbFi4QgfLwlHjmCg4e2z+J6kDQq+
UduvbC8wDz2GBz8W7Iz/EY5HLk0aaHhZDmq8UG2BCJkSoZ7y7j0IHCl+NEWe
kcZRlVZTbBVDDkJEswRY5RSGtPWYySpbnET9RxT7CeqFXKSYfhn8agx6WHjm
GtkJ59gQA/G0vEuLPPC10QPKIB/i2c5y0uxMJ46ftmywuECtMV5v5R+461uA
GpMtvxW+sbXPsLnVeBHivZQDeIsOBFjr5WEovE+FPaQxifk319isrGsPPUC4
ZWxSjV6bKnxhZsDyf0Un+aCSBN/mdLA/G0BNcOn46znTm8vXbq+E2ZHIZyRi
46FoxE2/uH1MT0d9bzxIrzK6iNe2R4Kvlukpx6r7YZLjjJRw6jub45BSYEi3
bTRN5Qv89WlxSvRXzlJ7tE6xk34BQHVWQmV881+xFigbAa933ntlPvvAwFIV
xRN3ZP2WrJTtCLuyp+5VQE44s7FNYlY88kkj7aoZ6o3H6OppTHlKhpUZVLnL
yPymKIpxp04KWxY3qkk0F+qOfNABl4PsjVU6QeJEAdFAv1Mxcn7fc6wu4W9F
OPnUN3RIV7FPGJAfK58d50zEbMg1MluLEID7Eu3TrNDWmxxnIIIXzbwCEQPK
D9b7M5WYC7IZCGawBawgiWv8/U3wHbyCuDgQ6OMpR/Fcx2Zfr3o03P4wm2u6
HnSnIt476GZ99OuuVhSDyNY4yTKDLb2Vc0SmBofvsrH+7UY4bV6GfFIYrf/3
dMh9E8FhtqAhOP4vM48vGaIb1OqkVY4o+EUpB1NWBNrKDV7UZsiFaDZ/o4Dt
YN/qBkmuJiPKurYxL8+/1GP1lCV5DHLPT/i81x2mQUrPCcJiItHoh6sGDRLK
vjqhQO1quFMz1y1h2Cyz2zuEmSYij7SahUVkG4BXP8zvsDU4aYr+RHhChfGF
UtG4PIrunvKzYaesQC1eWVZO7des6mxk0Z0lQn+/aJX3z4exqaxDbfbHX+Dd
kJg/bButU3QfBotQg8kBB4o26bjxzUnkrJ+uLD1au5XqkcGghmjTlnHdECUm
G/AE19lS2OmFLJF/w/MIRl8x7HoaUIqJdAFp5nWiMfm2NqA6OzeyeU5VKzeP
s1Aq7IkQl+VLpg4VyZ2gtpsCbWDNAwH6GRW8QGzy/fVJhvC/wRTokHBF9/Mc
oYxOGdIsGsLmz0v0HRTnJ41kO2QL/esWZwqbGgSkFM+Hit9OmzGhkv0+Ojp3
VEt0ZARDwI+n1HzItlbX5JjF7I89qZ/vaynn+75YX9OXzLLLOCxNYjN4XWui
5BkendpkriYoDXSfJULLBW/67tOHq5S8poS3TwXSZUVH1YYWCyDoB9xCBL4h
4yduQT0OEyyw1/DZtxG/8pT/49kcdmvTuQteHvbNXvBX/riZSqTz6tA4Uper
jJPl97JY5mMF7NCeK4k57ksllB2PnHcEIBButeoaQHef+1ZSywhNDy+62ZV9
SvKnyqbALYwvl1+4h3L1LOYghwVoXguDXtQJQBuYr9lSuhknk5xBlRhBFUVs
eWiGeMRE6l2BsgSkKI4EhRccmmrYOymMm0gIbLvJRAWnm8aMdf7q2SJDRPtE
wlKuLqqfuOso905PUP/R0di9cQlWVON+0uzxDBJTQoS4n+SbdM8QSb8cxa7F
JmSfkPE2Iyl8GHLOvCgvBM2FoC7OI+Lj3NaYXF+0uITFdQXPVcwSMAzJwIfW
iMVHQM1+ayJYVMgehLFculW3+CCVWc4FgzTLQGv6lPD8sWevEArM8u7i6bQC
PRHHIvAP5O5G2K3EkBzeyQGhDPqD7xjmG8fv+Pe6AII97LK3kqPNtPO/4sN5
fVmdQXMbrYoy7h0Bv73OqgMXeYPtpdeG/rlXEHsBNiZGw7BM8NB5n6bD2ER/
19aCahEtcGsNl3e3hzkK/C8mPQaeSBKNitUtPtZFOYP1+Tqw6pQE/ws5H3Jf
+n3kC9HMpmmUldzdSQeGFVacEiXSiltRcRTVtsx1Z5cRQIo1HqgyL+DyVBJF
7erxdQU8PGXwSWWZqlaSHPl5woBIlRCJxWbTe9/svzAADdVsDMkbaTxrK9MA
eNi5CoW8HPAPmnEgMxbAqa+nTw4oJ6BT3/EqGrwig4Ijna8XEeW0/0AC0YKV
Q5PB9vEhgxVupjpewf8t1VmFlRGVnqqZWYqHVzakGmWyh5oZZeNEJAz7dvs5
MdZdt48GvyAHaXGTZ7hb8FA2U7vQFc01KE0wK5XpBIIra0b8ZCaeV+7bnS35
hV+53KFYngwmpM8v5YX2500ra2E7C+rjabJFsNAYUZTZGmoqNO4/JxsNtrwi
Gtw3CWdDt/Kl4SL8jFSf/YSlkIou0wCj02uej69CYZ/D8GLgn+lEvxu61PIL
wnp8aexooLKbv2EPOlR61UAX9vdFrNadnbwEGwr0Urup1dcaTU/idNJTf5tS
8vmeq/Be6KukFeT4dahgshYtIwN7+NliOi/t9xT1uJZjQIw746OqmDPAJo1F
2sIeK1PCIAcYiY8W27DJ4Xuk2YU5hD1LbWu6w8H0Lxh1RpZxaPti15uxgLe0
yh8V48jDUUDCV4Lp3+fpPoIYGfdQt9Co0WKblvDokWtLdh8n/cCv1cD+JkdO
pqywlhqdRyo7O3kr+DIIC3CCKhr1rfR7bnq977wMlqyTm5OXKJAxuQZG1k0/
dNcPV197Zgf6QsHZdfI5k+8axZ7R34sparxLEKTFguKyE+R49BChvUriPqmm
WVtzaXv9ri4ltAOxUzrVm9VAh35yoQjrrosivE5MFvf7A5AQlhf4CFg66uKL
lWQ66FVJuAHBUMzc98BfMjoYuc0NE/FV5Cm+TOaCbjAnlPkpXqUx0Y6U1B9e
CwGd6lnrr41cqZZaXtq2kabgUdxtYCwq6Yd+3fnPs467jQQS+9oJ5VeyIOpo
AsRy3+SPjhMdZ2SBlU4H2WAnmuA2tocJUTM8/D4kCNAL9iDvhJiA8uZf+IR4
MZLfFtCtAVz4zepfuDqUIMe5Jw2KaEhcExYiW1n9aIHadSy7fxCe0ICOvp3L
XjrSpRseu5LooJ3o+Kw9Jji+slelgrRqFdEIBrQoa24QkPvdOEQnHtdd8vLD
b66msKayYeRQ3bOezyTB4SDL8ZhfjyAk2xBXC1QUXUaIcbErzN4G4CBQPYSy
YOD5kOC489mK6xmQYGcz99MPg1+SU8YgaSZpEzenvPcpyCNbDB0Ykvagrhb7
gfTS1jal6ON29lCjr/uSzrBLWX5/AadAyhd9E+KWYzOwnJufjFA0vrZiVAd5
E2FknIY1WWTH4MPrNQc7y2si9HfqEGqN6lsQkdACwN3arn9kYylDTUk+rpnl
bvNOxOIVO4xWVjs/s110qbHH0qCsga2q/CZ7pXTIqDeGmUdWemVxZKmwXLLS
Uq9oUcTl9CGgZV9gumlwVV3ocrgeulagDXJCaojjUGQdJtOfJ2EmQr57BvSW
uUAhMWlV3KH1so33W3AuBPAqs5z0E3r/XICOpepnI2xEhsbmJEPUSff46jAs
OqUz58Fgsxd3yRwxQAuAfYwvWriw73FMnZXRPQ1FWedu/MFPuVHYAFGWb1ra
y7k/HyxeipvJTwCH6LUZfQVG7g/c7J0br92b0k/hebncyrCQImuVtA+pbnIC
F+JFM68dmMIso08wbW6wtq5EWCFHwYY9s1ClltZE3hVZekYHk4FnVtrei0UX
7xee+CU8t4b7Kpfrnq9RqONe1VNlTXuq98+7Xnd5IXORuHqhKVk1bC5nq0Ex
SUJDys48D4hJGyeINdHYUQcPKNtXgFfTIjsugZH1zg1vE4QOpAvFQYuPFJBg
ZfwxFM66Z8txCKcSIT80JNF1uvEfexbTa0A4GIrfJ+RPE6FpMGNSNWOllJC2
lWJ3W3B/oY0h64/BfkQCf7dTYNA2XgFlhR19P8Anrk6h1cwV5prZLWnEtrOD
9kRJIgI8vZ0zN5C5IJr0KDEfFG/20A4tQynoFDNvw5dYaSkrYHBan9pYYFot
y/7nr0KaoIswNINQSabwWP8K1tBUnp2cWX2unfV/gaJ4Ph7vNkJmbp0uhEwi
TfmIhRGXXxSit1DbsEWkw1e6YTKenFMIBeLd1GTdgke0B9HxM6fAn1pnbwOy
jnlFMCGT6Uvg3D8qwKwKNJwzgflsD5VazmWYHla/asS+dyUsXjuWUWp7pSBG
lk+25xWj76k/0pU4tFF3xdmhqYdhY86b1G7VuyeSE6DtrmbL4+A8s2ERh3eq
t/SONMShx7D2QAhqmi6cKQsEMXclTziOceE2FwHM8CYCLrCAnMjQrNrkme09
L5UrAlRF3WXIOJnJGjbCfv5KS4ezZNOuCK0Dt1H44NBY40+5qcQT0kBsFvCN
PEaGaqDBFrUIYpHc52oeHyU60OWWTJXD9m1H/goFTO6n9xXW44IWhXEEqpKI
ERGrcMOzfQlNHLyrM2Wll1xquN9BTrzu9cH4fKtjj/T0WZp2bLI+0vwWSg75
Lsggw0zjkTkDGjT3UdNfVs+iqvgxsXDADGL3h3NUqZZDj+O9vsu9bpd/cano
sWMJmVXODGIavJLQohJNm58U/0U/lKYaW1HLzNCKHtvoEiQJUm5qPD8eEmcC
9plOQISakRWpIWezOw187f165xyNZCC740rWLyhDmrBxjFODskg1F+Y8wrx1
YWeE2Qox5tvPtUYjucux2CRHGit9VEi82udg8jyxjoA8/IQ9s9+l60cm6sbU
xxrcf3HYgx3C5LsmDpEtflymSXAlkFVtRNYiTBKbOlztsg91MKMDWLw40GB0
uViE4EiTfC/3ynlpdv/YamAbyIfdhflM/X/juPNIm8NJQoAAyEiZfmTE7hO6
aExI0XsZ/wkzsZNZaWR6tpRmHoRdONFdnC7XByr/DKWLoFYdr/P7voT4h6L6
qKF9j6ru2wFYvSPqKfHAmZW4GPRVBtPz6slD57G2yn0rF/5Qm/p8Ye37j/3L
yIHqpAaQWe2a6OKaDRAxese0+ZcJ2y5fpWw3fOlGlFHsj6lbchySfFyhFkX+
hGJIZyOGcJ+1F3DbIktiFWj5H+W785HlNoq3XD/KVahDEbZyQDn+027zxtOj
qG1bfagYmm++YahCu7WPQg4QRQlF22F/xUQqeJME4MmyEYNBEVtkdTCF8A6E
Yrx7Nky7xJStsmlb/uFPaOEX3GMZGPzEF0ccE0jDTmoMocLecYbVfCyC+nKe
SSxTc5JEN71AxlX/4YBlXeu2vYJeJEhADxrbuVFhwDIeQjjICb/7SG6oAcI5
8k5aHcc3fPaYXGRICLhnCvdtJKltti7EKpw0GH+YV7wdoH66kdmYaY8tZ4Q1
+qT+RLHPU8cNYhgXUJKmHpr+3a38Cn3f5wIIE5rgcUmEmpeCBLGQjTUSIrUI
5sBGuNFkiZCc5DJIAPMwIQHyA2El21a6z8AmBZrjr51gKP6JYJwHK58zw1gL
bIpIHck2qAys9ZJI/54/U8G1t/JrHObB6lzzOyHx2rsTtuaMuenwxRsJ7NBu
N2dily8SozxWtueVKFO86DUlwDmQfovg3yBGxTxagSENeRMLWSZZ6E9vPT36
GMqgI5Hbmjmk7eAFCQ5Eu+p7hrYWVMjFXYGyEtks/zgnOKHBlzs6CGwUKnQy
U3yYCLWA5o6T03jedRnQYF1nzuhPDuWJmpCO19AWkyEZ3NoxdEDrRjMm6LIP
UNI7ngov1wLlDAKDzOueJeQDedYIuNWVF0b1A6+QIk1DVex6Dvvylh2PcqxN
uWdfPYByc9NB9JBv2RyFWcZo0l3fUKLA8wMmrA7zEEoe3NtGXp/4Fh/22Phk
CzWaodTgM8B/mIUgGdqQ8aUOmQDX0O1vZuJB8LhfGxmQdSrNDYxVpRGUJDht
aAwM65Oa7UU0fKY7W8G4Z9riooJOChQMEnG2TWWZ/0rZth0YIHaGNWOzLWtz
Trtn18jvPgC2Gvm3r70MmXeYYNH2DULyKQokI1xrVbCToYWQw4QsOnQV2El0
cP/VLQPQXuphMShs6Gmoyy0sFyjZHjNhGnBdc5DVbkoUwzfdpNMEqLq1cl0V
rPBQNRyy/AQ2380Lo1e4nZNehSsY3rRX4aHgfms+DjaM1kCHF+pWUfE9uhdc
/XmGqqGJtmYIxXuFbtz12sr6M99Z/OfeeusS4gV5NTzgYqZ11sX9leuBLTve
2NEaG3cB6bSR1ndpMIqUW3ecFdl8w7heqSczJWI5bG7OpnuZYqhXXZBotdKm
mjEbp0/HEw8EwawchgyN6VjOtpBLrH83Gj5/MJdJmCY82CmTdgGnKFXmF69W
6UZ4DBtQOe5ZPfAofwkUZVE/VuwZ4iMCKSlFHft08ZowUYTF4puWLfXhH6d9
oB7IfE/QkwrvqYuKUFb86DWOWcGONIVz7rFlMqUS5+gu723hf4idKCfBdg/O
Twn3LMcKp9Qsf6hmqlRiPAWIhFjlzq0glxzH81NCAmTdVQt6ZTxFDBinHkSc
zfJB+ewijfhmY7Mq9K/ImdsSJIlY5/HeT9F2sjKCEMeVDb7ND/luFSQdL2a9
eNxPqGONv/Vc/uLFl2AbzGw7opR0gc1y/qrxBxDCeC9Mh3DHbQyWLK3ae2sZ
7YId7OFDIHnX0R6j6dg3z6iZDLrzmdry48nH2QU2cJ5Y3u51NhnI3uRwn/6B
gAgOenM6xrQuuZAwLvCT2ZS+7yGBwJl9JseIMiS559F2Ff61rQ83MTwuNqlv
ml4omOeUpVpelYKOOzV6vQMTMlmmIWSe38sWAY1pNDTIuRrRlekNvBAbcg7K
3Tqw8gyqhSm2OMjc0cMnRUYdj+tCDNoP2RcSuzmZIZ4ArlKI5fhibFNw9o47
SefexBtEWgWHe3RiNLkjRvcgmP6roza7ZpVQXojSKe8TZr32jUiR5q4Mx9sT
Z4EHtuKuqCVR2r677Y2O/IAkNV4mRUFJwRGdRoeBLXoiAOmT7NKHvU4MaLwI
BdSVPMSKXIeJRiuHX5iTsQTLrqxmuIOX0HYr4WCUW1TZ1LcMdZ8Rc/sG9oAY
LJ/Dcjqfd3pLfhbmM4n6Fo+Ba7h1RrwcYT4VMW6dJaTv2drA50cgN11nwGsl
UJEhHkVD2JvFi2XDcSSuTSjf7aT5TYRjuQmMH86xUKvjqeVY1acKtvtoGppr
3Jmi68KFMegb2vyDBw7e8BOjYYgi4RLRN7vnCwOzpmzp3LmKYOF0XpvknGOE
Rrmoky6aeX9/+pPtjIYiKejM0ME/RC1UphKiFSjOo7rmuSnZU6Bi1la7ydG6
RbPAuzpCdObbdFoPA+2/DxSr5KXtgJGoLyNQ7sBT/tHN4OO/gvpEpaRuvdir
vzYwMo9jDGKA7V1auECfIBBCz8znZHhSStY+x26cUxgKXcZ2wVByALLl0ghg
EQS4eLaoCuTxwm+VdwSfKHF6cyGOMufApzPvY/xiJ2a8UCVm16I9pgEiaInR
2xJaKWV4dueIDJ/v84kpd/upjMQmCsnEeg+ik1HJQp7h0lX2nQbBjS8DR3cv
oWFSjvISs1KLo1nMiH4VCaozV2A0DtG2SxykbuuW9gkRJRydIGr/8k89pc5l
ZqSG7keC2hV/hRkeDi38MC9nbtO0iePesg3mK01TbhtYiFmzoKbQpM6AZvLW
zi/baQDA3EBf6ABOw1XTmv9CxIR0ImVeg+drRSxnRGP3cCzb/dyV1CHGt0Tc
fPPyd66F0dTwxkqzj7Z1PC9payZdzHtj6kJCxKDTSWCz03IdxdChgxT9nvfP
SmfjUTPyPpYUTZ15JNN3TRmuDPOdOsWpAvEk2FKt3+u4votjVtQJ/EtP0M4f
+Xr46kgy4PHQHY1F9PojKjeiQOTdRmOswwTmU2GBERLL3614JT+3TsAlOJkO
eYyKmjAIH3kw5CUQAWrKCypZE4LaWnitU/wM51IteJwUXgTpBfrtLufBUOrH
qRhehWR3ZrZJcEWdYTsdQcuGx7FCOgbQAfmd+vt2NBTsWyDlOBvgpNooRevO
7KUvH80ktOprJEdxR/4ZQc10154RyyZlt6AzvB6gx2azhu/4kiAOLKVnTJMY
YDUjzHwt0h5RHQ71Z85hufImJP5NDa/qcGmaNvzJvExB+ENLViauP6giFLAs
Mf8I4hfqGsQ86OBIly+8Y5SxB+WrUtGGbU8vuaowH7IdmjQKnm1ibhCMRST0
jtzGn73qLpe4j+1dmtx2mTSUxVEsxpBBhehG9XJIiB95pNVeeJIHF9aXTkLe
x50Vpu7XbwZ0VtMBfpDkrDBEdmzSSQwZX3JG88GCNkzB0WUYzZnzOGG+Xedv
w2srA11sNT6y/0Qt0iAMAh9epIUicJhVyVOKIyW014Y6Ec04I3AhJnjhVctV
/09I1lIEweEebMZhl7wmFP4etUe7Wqjfhll56/kDMZQYYTVSsrQcL5QdNb0A
Oaob825Y8/DsCOi2Mp0UdVaDWjkgpbzOVGgNEc2peSh/22+TaXVH3yEDtuoR
qcKDwU2uLiQxaEiSB5Z0qdKCUL4HucaC8t8rAs0FbaDX9GZVB27fSXUo3jUm
Qfi+GK6z5uao5EIwQh7lNAZ4Ngf3u4qKPz6NMttYklFziQWO8RsRR8hvWDeD
nDScdLX8mxBgojlXpqayllnYhUcvLp2dHwg9636CivaZ1fsv1Pff7u2JJ4/v
HunfHLqk3r/GzJqmObPR6DrQJZViZFeCJ0fkj2jfF2ZGrdYpJ4v9ynK8LQSq
nAfCYK7jy7WYbWe97h4wD5K1ydk4LGGwi7MMKnUskRgwp58xs7RBefwfBsLe
KawoYZau0OAVYf1bET7cX6YHrM7b/JLxdUrIPgEEMGrPLPdDSMbkiAQVHLF8
20EiNkFmqJuHZVtPoMZPeqeBvJDvS08VBZkJMhWm/iI2PQFftFmh4/RVN2t3
ERzRrEuCsQml2VAP0g8NhHzKG0ZFqRlERk0uoTictikq6lGHCp2l+UxZIssJ
g6v+af0qE/MKQlC4S/FJVrZZBHs3dEznPcPQpqxjttexnbZN8a3uK727xj/l
AeQxZnXvLpfw48TIH0aWr2MXzMSWvIsV53o1b7JmdPUJVR1XrC5+ExlJMn35
1pvKwQjd6F7EAU3JZ7HE+wgYM842T8dPROO1C66uJ/BYJkwXmup14qEVJIqo
9vhSYBfxcFO+3SOjoY3TzbMTxLnkFEjmHWJr1l3WHev2IdINJIp5cAhW8RO1
gUTHC46hR/h0zuTmSNLjYDz6eQLN22FQuIeJKY9cp58QlkcgYteDqdd5l1eB
eIjBAdOJbs/92zTTj4pOvqHSQj1SULhRzKkufCwnjnNLB1u1aVvinPQ0VMzA
l9ZZ8gKmUSEZv9+fxEzZ+X08TrRYbaUpflUzTM/VDuhuZwwI5lBWw56ik1Tg
WB87od34ai5+WouBYV5zryzJADWc0+3LhsxhMRhSlBzN7wsD++3hTF23lkKO
SFnvKyRVGrIK6GmCqAN5Q0Dyt97o4N5FVE0o6/ICssy72ccOCHSCgFAygUru
ODT1u0++YhTFXhW9EvFpnZ3qvTyzd9px5bGz1bSdcc/AFQiV9KvvsGdg+sJh
Fa78mb7uGXqKpwsQ0Oc7pfBtJ82pEjuGpnoC3fcmKOOZX6TuDyfS51taSji2
8b+h/BXXq6Y6jk/QheukuXqZLV1sq5bzxKSZ6Nh3tc7h3MbZFS7Kv2GzRYQR
/g8oKhnviwln0IKtp5akj0VAtu4kpo+76KlPOpmevnL7wetb/krSyIQAkwbO
uuFpdCiFd48zMcFxLrVCFt7Gq1W8xet3eMQsXvCzUr9VahFGfITGksBlBsWN
ymcA2MdfQUpkPLuzV6I74w1rFM183kKI9VxrmbLjcyBtpiYDFVj80OeIRtvJ
KggGW6BjvHRRGG3GybptIODCBAbZmBmPpw/5AA5UBemaeO8Skpt8rWXKlcRC
0pJsrO3YDWrDaTUalIM16F+nS8zOcg5kujjnjxWKPZBbdVDmEj7EvQvALzrA
pgv8Z6f5wOWA4wBwroyJDPXPtE90DtJHCEAYvLuQi9rDyTFGTVQbh7gPDH0k
vRVXh9L9FCtprF9rHkXRjw++lBE8WXMa1VS4n3FWbgYDVkYdLcgRTJ17WTh3
mCJ641DTK4ChfsDWYd3S5z5Gstb6+1L9KLIxantUXyDnthJsegNWAgE0pD0W
mq4Vf/jc00/T2Y8AJNBmk2J6j5OQrOUu8fV8wtBo/bVcnI6U1MbDkvXTRGZq
P9l6N2iZlUYcrvKxmyE1g1SDe9/JbBtiaENeGDuLNIg3kY8S1O+YpCn3BaLD
JJ46E6D312vLbyaEpoqAmEoDewkSKjTZ1GIJWaMcLCQStzSMOMZnmV1M/sel
b1sxQQonzQc9fXZ5AuyRLyDjSDQTwXrqnKzdFRJYxOpXCkvJDNDK4HDwdPl6
JcZ7280OUZ6XYHdCySsNYM1UoKI6OH1gajEv68q/RFscGOVTyYRPU/anuB9Q
1hEmjfjwaF1ZEbqsN03305KGQaExdHLWbpNrTRSRdWUiqtpzCDbnJGjhnQRB
rG0xTOkA5HVQW8m4m6QEMPM5rMJ8FFCSwSfEPkgQdGMnvSajd9ETEu3Q1uO2
7gBTtXohJwOmp4VZtNAQAa3xIjFOCS0G4SH+eKJgMlgUaTZnd0nljpmV8egA
3ufWznzsUxcyjQfHPjPKgCHXfxntyLNXRqR0J4BW8C38fcBv6D1lsuniR8bG
gmbV/hGSlNqu33FVU3GlY/Cl6H4S9I4cOicYvtRrTcTnr1XUBDiY5kDFpUGn
lRA45he0WMtKIuZvreRuzez3qoRpt6TkSen14vNND+IJCMc4hS6AJ6KSK7X/
+cZBrCtl9bDewOJTO7BgbJLoNuhr1WT8F4JBejf7Ty7p+exJnTezAQO+rk6O
JU8jztq1fulGdfdJ13uyUhMZYE0hfbvqXoX7uxNSabbLVzpxuHISAOdOMJY+
Ldyts+4UdnPwAk3m670h2Q2//RiPbMj1HuG3e8189j25MZKLi12gkBcNw9CN
NxAAUccSSeYeT7nBwFpilejBb1rlbZ5mo5e90JggEwQqMEPR3F4TQ5TIH5nG
d+hLyFN/c0cJdqs/FVa9zDrKZaqKMnGmHqsr01Yahx/wO+p+X51S/EpoeA74
EcjfxwXaq5Kcu+xo+V2OvTL1ZkEpYCwjakqHZh1tZvd+Ilckb3uEEslaPRfD
IznAjEz80Yi4hdMIeR7eu//EkmU/Bz3SvcphzAnN7Y0q2wEzaMyE4fmMW+Z5
RaX8hroJJxhQkOxKqp8xeKuTnSJvUTnQVW6FYzf3MvyLJROV+XrSQnP6No2X
udOKH40E2jxwMMBMG9U4ZZGkdzj+FoPwILp9QvPwncB4RZyGuwbZKVS5VeMd
kki+91GX8AO3GBJNqCfXb0BY4ngmG2aLmGeFmc0KrYwENCCvstPNnURTTn6+
znWG9o7jyA+QtQ3dJ9fl+omchJ7zI1IERAM+uLR/bj0F1v+nL8BwZpxP8AXx
wYHKLDZZznx308mShvDOeL+Pv/yu0bAHRzDQANMXpdnFgKNXQsstxJizK/bE
cCWaN+ZnoNLtPFZZooQ0nhIGyUEPuzVaAmD6Dhee0qM0dqNaoHVpsQcxNb9i
0+mog6qwNc/oTN3qjmX2Nzwu6fX8j1ik2PBfXG2P0WgohrLimu92ar2bwijo
Gt52mbTzjDItlQgFWzBitPIOl4WNaIoWl7hDWVCYgzlk4lCe1P8SmNbntxLL
2XIgJJWicfrZShMRnUq+b1Pqn8TH9JeZx6a76XhyeSkocoPmVsq/WKHCfSTr
uFhZvUHiTTnBXmV8KyFGi86pkQXlBpai72/sOIIBcmA2KM9icDhhJdhX7eJe
TPixCq6e0aG6jD3z3B6QvjVM4JQWcKAI+lGz/HVNZkBy/j3utI2wm5Du986h
pzBA/QK4FsNjq+k7culOaRWPwy/bRczuAsFqyIV0eXRc263JweX5qxdUmzut
TM/IAVlv/leCNaOLbnoz/NILf1yu76Du9Uu9x4QFoqAUBcVFsUMtU+HBcNW/
XHo9HQ/GDIlyGW13eDluKPRoRhGscpChqMz5pS47HR5e5x/Etw5n9yG5tVYk
54wSlF9c887MNYg0LiPMD3qD5QZFVWraEPGO4E1CkPH/08lpVtwC389t0plu
5AfCREgbfvk33IKZYXNkFZVhALek4wGpKfYPZeEEPsz9aSeSz5/RQZuF3VYV
zzqnZ97/vBi2pNuLrHvb8Ed2rTmdT6R2IUNKNrJ/5Dl1zSA/hOVdeJBZ14GL
fAwVMgHMPiVlpVP33/OJBOdgHKEjOi+bS6LvcwoVEL0e2BflyHCIAVxcosbV
SDHmhNjjq54a9iwG4FsKC5i2qo4Q/kz9dApktUrpITeQtGw/g0YK7zFx/jJ0
BKSdax08bXXwX6CkZb3it+k88cpji9X116g3xxi0JwJzb4Gi0JZAUY7Cc6En
goHKMPzoW0/jZtEEIVmCQRqKPQxy6h0w/9JPYcNV6482cbv4vi5WIUorjLcw
zm4X0WFH/irIwadRPEuG6OP52VU1xowYbbQpTWbqXNU/NDCeQDov2i3WvWl0
DcljNuuthlM4q1klfbPFY2tEHjtyhejBxIxhgNPEExm3AFoxyIR5gk60TLGb
Vzhs3V0C32GQqjUC2haSM7ZjNdjGnuYudtViBR7UL+YjWh3w28Cooc2F66tM
dDqAP/yBKlEhLsJKo1pt2OH4o7ex+2dpBanTY/99fLq2eaHduJJboKuQlrkk
cit3wvQJEyra3vGAAbHwnVphjvfAxBv7lGUNckkoqgRbXWpN9DcmvAILte1w
SDA2x1xpKHmEw69n0KyHFUjs0pEHtBJftAyRscAlQGaNm3cUGqmHvAkodzpm
8Y9gUpd0z6GA1CQwzC1+DOzXnMPPZ5TeHyr3kDF1ROIhDskzkofhs+JgYIhg
8uycDO+7t+MyrXXa89bop2DZK8VZIWmLZv5jFvaXSSUEeAr1eEM66vDIyMPL
QZ7KliXK7SzxzsCUdl4zmX2AHG3dd2mEG8Fqz3uEWGDAdm2m23bWKNVFOp3r
HuFsbca3oYc/18kuteEPud/hrbOhf5Q0Udo2FfFPVVbSwXGn/yzxSBY4o7iK
8Blw2qLEXgSLgZgl0l3VhpjAYiSLRhYtTqKTMrn4n9xpj5MNlvnVsWALtfmE
BOnaoVcpYSw4y3vbGYj4q/BIbHspVNaKgOnd8qGGRqWRD01dW9nWoSycVHjg
mCh/LcPI1rtwPg1F7olyEbdm2RY0/vNOZ3qR3POfeuL0Ya3MUmHlrekkoYsd
ar9THemdBrJONEWai8gZ0cet4oU+8cyDNJAIxnLfOAhzlzaPKmKYKjmTy6j4
Pc3L5SGy5Qz//vD3tY6p9zVtmlrwreeYPfnYJ72SGdPtftIsHlHPGDsSMvOR
m2yy1m758+wnHlpy5M3X5MTBEbbiB3oN1vw9hjwXO8vOG39KZzHsxvR44YA8
nPp91YklAOysv93hBZg+LSH38zEWln7XX7XBoSkw1zrgvKVclqa6I8dkcKN4
Rvr5ymj3gKGbDAD6yOfW+UHGxQ91IOCzvNNY4FqCSl6URcFiaZymY+9T3W0l
lMTEuB1y3wy9HPJocptgzNNfkCqiAkgz+AAfAu3ifIzKzvJpj9nfzVaywHxD
RLUQF4FKPEV8zQAlpZMHGZt1jjJMLO60Ak16ycFKmDyEUAXN+1cgVVkkk9Br
qtbb2fM3UIsz9+RG5Pfm03EZfGxOJCHXWMtRoN77VGymrTeyFcpmZ855nlEQ
yj81b1SfZxWD61erR+2AlLNbIV627NXksYGhyCM4t+5/EHVIWssMee3YMDEZ
lYy5B33T336Jhqrb9GxlERkQ/mmYGx6cBN0nxfoBc9P+jGFHnPgebDAJkUb/
QNav5WhmkvKcBLc7zrGRvBFSKKAep6apGU8T4sNiNNoJYasaAvVQyBm/fw3d
DxPeDONQhkK5Xoaf9XOPmcb7OfFhfG19N4qAXMQN1uIMvV8flmqnyxdUbysA
vraoLx4847MQMNmgGllq3Lr9HJHhM8pb/8aQ+RpRoI+xiB1VOn0btCR/L0TL
CSXJ3ENZCAr/I2DfRij0U/9RlYOoVUrUKET2l1mrDD/ZNK38MNrECkohEP4J
RupwVl2DOz5UO+582ycSu+BEYOZNMOxY/EIn4npnkT0tSUTlYnalDpLgqGr9
eUPLMaVxEPEDwPkYkZgxYgK/SWjW2/+IIaTRxN/aMBZeuPZUJ9WzTCKRg05m
Z2isiZvoioZ9u8cDxHAzMmFzYuF2gpWrY69OXDiU+Bo8SgEH6RO8Yj51Ka0T
CrKi1tKXGtCxfC20RyG8/OC0PWX4xFJo54eYsUvQTm3rOrUgmtc69/Cl8MCL
LNNeFmhI0QDuOS29BWZyQ1/dQNky1J2Ei3w34w06puZM3N80/s97QY/rJKqX
gr5fR25ZH5hv4sXUYyvcG7dT1j50hJhxVdfTsqSQ1JnksqwpVgkVAA0quzVq
8Y3x3AiBBwL5aate3bDJgRuAy+iFD8EXb/D+5I1BY0dnACWMpB5YNHSBK18k
YGau0U7ZLQB1YrNMk2hkXBqE6xhLyTkMUrexmuUswKXSkPh0+4Pu22pfAJMG
Cu2YRhU8Sx7My6l6DkXljNZcbe+S56WwqSeDRW59NRUU03M1CfpLKOVe0u/s
LaFSdtvAQRBKHaJ4zlWcEm6hB0L+dnkxNyA5jjkQVW+Vzx9afbzqLWVdfwnq
5rO026NiWB2xO9F3wzAUCR+yPylj0nbwAT52MOGyW3BhC/BnFKhxvXijYM62
ixJwzwfnVIhwK+1fJ4X1hNjXXimhE5dRCZDkHFtnExeKYP2sGXH8W+oOU6Y2
3TVxI300MmHzNPx9po7nFpHT/ss+7jUhWOTlSBdr5/m0R+1ZgDuJbG5YRjuQ
1D1a9rwvkdliEXxNB6a4KZG5ahVRI3KERLVZJjMxdjYMNSNBXnXxwhHOR1Mu
P+OZRYm9XNbOWKPgZfY57BOMBXgeKPHDmM6aa3f4sZRMJUSgLHJo3d4liADm
sXfgLs3Y3wYhZPn4lqK8D2RiOyZmMnR5oAnp3olfiutqFGSf/aMtx+0KYz2g
ZtntKfWzA1oteCC2GOsSnGZi3IhSbzXh8wRsrtiJSD8aCGg0tDV3T7+zx+Zd
NJb5s0B0ZFZexfl/A3yKGnKIYBg5adwQ0vsPwF+IxaZAoomVv9+yVn5JhYNh
oQGojxXvt9e6rJIoYQCMVFLbMG2PtmmXf6iR5TzdrvDG+MIRnOcbJjvS2cCJ
QwOt9LucmygTzCByL9gAmGzGMAfSTrgEMDtwIlwyBQG5dVCL5pM5MDnem3H0
Y8Cl+rycl8t82CRnOC+vW2n59xhOrVsK5lNkmyj97NylOZXMlRImF2JPbHJg
HC4BaNNDYVROa1O733dVxkf0b0LyM+cqIg5HtcISseSJKemm3LNZN4iyEPKu
hQmI8RqKEupHmdwzg0i3B8jpDIROWtxkG0p7nOff52hcsXpjcOzEHW1NUzQo
Sk8aXjG/LKLjkgap44CIwhrhRE3bQyHrh0Ti2vS0+JBMVpxvoCeXqN0ZNh9h
QNYkOfh+1wtoorMK7q+JvOA0LYpzOdaJABZjswcDO8TObfyTBBjyVDDzhb+G
GcS7Hsk7e1lhyGhrPjNpcgvOYtueOdu5QlX6s8oDIktQXoiSo35VSmM1V/tX
gMiSIyUJKUiJLt3RiHgH3lYrGeN2Wc/ylvidyFAa7kCQdOSdtlMyBIwmpL4v
iWqRZuTlGJ4ajERpiJcwQz5LUXatGPJ6AuMGtb5DPi9HRVvbHiePS+ZwWhMS
nYuAVImAmHANx5wRR/nDBZ1KI1pAZKPXELhrs/Z82UViUl3u0arYUzYnjdU0
DtwWLDisU8NRKUEDjMC0epL6PcjpsWCVmL1zHJ5aU9ffmPFArL5Mc+lPqN7i
8alF+6xTQRvhe8Cns3TZBv8Ovc+VgmWtYVXiuYMe+FttN6dyN7EukXr88aDw
gl98TYfJMnSmDyTpWHuB3RFtZPKlU5RyGa779myfGi2wA+kFT+pxYXPPaFAf
n2rqWGMnOyZK0B8ULWbvV0h1SZ9jm2px6+GAwJs613zzJUgNwq//ZDP1K2ec
pGHqaKCnwsdHopnwZMnhuZXD8oNN/Ou0Q0Amd4UGoJKhezHJ8SffBoVT0w4d
pafPmbcoTru+aQTEXUkAyPjH/Vkx55m8jiAMLH/JRDk9rtSREga71puSw0pI
nA0xNgvj/eY7SFlLZHyG9Ycmy5qa/XfRNZXtjWUDu3Mvze+lLKlX8od5etQu
Cmm8mlYeMxPafhAa1W9ukIoCww1lfEEWLz6RUkzN2QSGf3I26wP/W48AALt4
vzOUNrpn7/Ghd6htFmKy4IhtJNCBzW+jrM5kRZ+QBzsWrs9rG7qXq27FimBh
6fNj6s/jRzOiv/2GwsvOQ6G477sWumqJQQPx8iTQ1qWB1FwrLTt7jVd/2R0k
k1MsQ6LSVuGAxKTOtHswNuyWTJ6SwcXEYUMPdjJmtZAnZ05AJp/UhN1Qpr9q
z9lXSa6XEq7YU4qICvLIAoyHHDH92pHKRJ5afxrDUj4mQ8hXTDLsAelL2qLM
XBoDTtVusTP+pGeDJkctxfYshxRvIGfg/DJlkmwQEh2k9Cvcw4Eq+21jvNLW
eUqxf8wOneoEjVb3E4fcYcV8xz/ZeG5iuVv3RKIovwxcx3viTnHo7pga47Pj
1vJPDgHrcPZULXSAdP+dYxckxzUBzxgHKYxK0i2YrAB5cYbvRQn3zcn8XfbA
cygwxdH92RD5e2fImcHRLGhufsUNyMGj5+SiL25M7WrguSQzMkL8fNDZt/c6
M6GAd+aIcolQhww8+n9J7UcgG8+QJ0mv9H3XQmddOfgTiUNKcD3/zMBw2wT1
JzY5qL7SihuK99jFWWy9PfsL46dUi9dbNY+58oFMGOtSFpG0V4wtmqp95oJg
nys6B+nh7Z0hAQJrw3EYSVPDPW9I1WK3gHJzI9IKBxscpI2I4oHTKzI+Z3gn
E+ol/w9nXntzx0n6LxSOq8NJA1NJAz3+HeDyoFetSo0YO+DZ2b3fne/hxWME
otxD2++wXfd5msiYk6cdVT6fRyqQH8iaAB95dx5tvgOEt2YidWZpSjeG8r/9
Myi3TL6yVrmQBTArYysXwMo0XTTgohyUAF72oKLC+17AN7OZeOcsAvuZRTj5
LwViRkX3dTPK62TuBeJy7DNo06Oqb7GH+gJwUoldt0c6X7Alpt6hXSBV+VN7
gPmA6YzTYD1fAe0afLrdAevoldUkn0zF4nDxKmo3NlFmZCsSCH5wGfYiGV5q
0kV+KJFE554yiPcZBaYYjLnXXQtGPmxy6alhOyJRrB4LR9/PFgdk1tzRnMN9
ada/bGq2OPDnae9i+RSY0QvuyuF6ov1DxYwh0GpzPwnbV3LzCZpoKJh1dsc2
DYH6PmoADCmq6oSH1s2qKnBeSk7zMMyIDYV9CG734EDUiR9dQYm2OlB96pXu
izlABPpqRbCz8rv5HjAcJpLlHL3xWQabxAXSI4Zel4FvtwrPfjprbBcMRlkS
b5qvRZVfdltx2Y9/g5ysnP+g0fSewGKFxIGrOwdKt3RG7CAO+0pd8KXws8s6
0uLqBXVfh6UngGyJS4ZApCR3W9hb7/W/8RTFsqck6J/YKQOQwwivhqVYFHHp
fF32Gd3aVmbxHSUQMVAx0z+bPb4gn45Xsv1zBpoTeUUAygmYQnyE3xHoU1IX
m5oL9QC7pErKjU82vtmzlYRZOlUjPzjwNOOAkT64P3klLnlscA/mqvkAHZFO
Q8zuZItC/DJo3egMnGfMZB/qv/FPUDr1/IUeMHZrVoq1DpUO3TJXNYEcZePN
dA1nRvt/903K+ddhAE7/CcDdAbh0yvKDW0tU140I/AWudAl+DgTgeW8vyVnn
541cGnU5L/p6Js0TIJNJbM0pepsjiYahMZ5q9sYHMUMOO/Q3IEywIhbwYrCF
h3+Me/0rT0rdelX/LIVD3aYqGFTG+J8E1/ueowpHTh9L2QD1uBpU6LZuBAQe
WbtEj5+tySdT/cRl11FcYfTJitjd4TjEGrfY9O/MWnjAN90NoFPwhYDr6QeI
0R6I9q+A/40/yLJ4f1AX2zztt5odzeS5y49mrhcPVH5vHP898yqcK/pOb1lG
FKcA2NtKotrSu+L6cA3TUWyNnfnXyTF+4HHeeoOKMgySNH8LMydCUKiz15nP
V0ALj8la9C4fdrwFPctE2MTf7bYEz9IjQx4FaBdwEgFDJaV6v96SSVjNLBtW
xgL5Y5MwhOmZuz6OePW5XwWrrazpqwERtHWqDdKvLn2zJpY76NVXT4CIHyoc
G6ffZBJWbzK66w2VOgJHQUs5FcTIS05QicjgnbkBQ7COHJLEupEvZ7W3iUZ0
lVMZBkY5GVc+e3HHTfuOJYT6j5a0x2YccdFJF81Bxz4aqNvWeOSfqBCltf0r
P9PkXK62TEGIsUfrVJB/XQ8N35m2Qv2O4Cfcvy012rLSE2xrsSk9FtB35ikz
+wS+k0T0WiAiSAQykB5TcCIjYqfA70tQUIBzkHzKwqxp+Ngmh1y2LFhRZKWu
EjL3EpxREBUVM2QzfFb9ZAL9D1DrF+A21pfRUa97LfFB0nvK6uoehUqjM3QE
KmhLWRSvKI5KDiyDacBBz6k7+hw6LEt3jbUAVv4ZIRb9A6MFo8jJGZkVdita
IOpkMPX9p7y9IfnTNSzXQlOHJj1jm5K6gHzfw/roGwhMKZzlUsnQRTk71tbM
9Yi2yBS4zzYY16Pl5CJutqmkgaqmFvD4PBid7Wzdi8XcFenr0kiwAvKHhvbZ
Si/SxacXh/4Wam90P7yDnQjOx0oeVIhAbGHaPGRCvI3Z9YNqS+cty9WZi9qe
zGMYpYSwwex/7ijO0FTLdfHkjtsDSDT2eUOEwFHobrUsb2ht2R7hkdlwOV0i
9SeqxriWTI3VgLlATHzAfHYCARZw51Jv2wiA8ntvAmk7Zum/u2jjN5CdaWyl
I3Xqf0Qihezhh0f2q24Mje5DKCRBlFiUvT/rQbQbLf2H518C0hxbIYazMP2L
pZTqSyGTMymnjfgvE9R1ndKIFZ/W4KOSDTI/j7pYB+ikWJ+H3Lq42VLykBxi
zb9gUX3EdfsL0PicBpf3pmCFlgKny0UYcnYIZIscRc3vDVqxQZWceC/R/xxe
2CyCbMG1pDpRMjDUC1owaYaGHVLAJmWljd/Px7dGd4WKy6PP4ExoUJ0vyvz/
+JJOITX5YbPujkV9ztG77D3pL7BIedVkqolsX3myc/Dx4waB5wa+KOsw6yzC
AN/ddVwYkK4Wal3zt3QE55oZkIBcP8wz7r+NW4DvoUvxnhwk7PF7t4k3sFF7
wLahbhxBxYxDtwrZTky3WhJKpadaTn2Z8HeLjaLpm0bf9vAKqUOWezNw7PSH
9DBcdpPwqNKsitgb9XIRIiapfG+Oez4J6R/vC+/aYcH3ENy/jJ31F5oagJ5r
NkdklpxcZzDW8i5hbrexalAUIp05x6faUdUURzjDb+idnS/o5JNoDd01llRa
tE5sbtCmxQunQxjgan4JenZ2TbhKYlXKKKQGEIiDt20orwWaNfJRJ5CbX6fw
xbUZrl9EeMvjmbfbEhooVaRCXa39Sc4ARvIF55tHBckGjw2shT/6vlAF6yOq
NO3ru5lRkbH83DSnA4uVXuIyluCbxYOrmyAa1cMD3R86cUUuPFkJaSxVJzml
TRC7BAj72/ysQkTnTKHFjMDgnVERbnXr9EcHlxj49VLyteBoOGS7cOdDMK7v
jq5xwriCLCS1T4xtADT1XlD8b3f8rs/a9ux3pMC81Kx73I6VetKMa908nPc1
ysQGplrleZnaHCXvmto29oeDUWvWWCM+gBTE04jJCKfg2YrvcKJUcCCz3iOD
nF+MDI+2fP3SnQwBlAx5cRaDrNC/oCwVc+c+xPrk0USJamuICO3zyxAvR+Dc
kcoTMCbLpcnPkK97DMAT+qWwuKkZSkvm0sGt+Uhu+UUwp46wL9lmYsfuGahb
xF7Ki2xhJBlAqk2cX6KIrmE9MUu91mZXYXFkq/bHogdb7kSp+WIFY/1SiHpN
nVwQ76OwoOYm/bxpkQWe7/HpnOrWzWq2hy0H3GpuAhMs/NqoI7QsE1ZwrzaJ
B0Itc5DYYjjOD1ag2ns+wP7RefETt5Aqoae/7dHBfBN5gHXnWhs2m8uBmDbS
4pult9h14MN5m0Vtgfs3rDa1R3PiS8zbEExColc/BfXcM/b4MZR6nzwMepAT
fiJJ9CHwbFsEIsh/WiztSCzywFPLuLdXOg4qtU5kJURp2vs1tSuIc2zMjXBG
vlfgTbhGduiwRTNTIAfU4PHeIwuW8mCFMfKv8TuscgoNhe1KvXfD7KG/5ZfD
/Uc+Tb1yzMZU0vgPRxxrjlEfzgDoea22mFm4UT+mHhj/6SsxQMulMayccLv8
JUvBuqYPpblf9ApFsCo2Vvm1nHx/eOlk24vUD4MaHks6DxisuY6TfUSnSrsY
52G0mfc5DVNtRL+JKil45pQy1xQRIOox7MFi0/cwCUdy2nZd2hT4Hv1rgdFU
dNNsEI6SiEfQOBUgK0S3lRbvEHzZDZpgJ4fNtRYWZghq7UB9OJFYmkqMFVYR
/MOv4glvJI1hq86lNV3tjC+j2tyalcFQdD7Or9yiwMIXTLVhEzuHPpRH/wI8
rUNLj0gpKSJH+ZXkTcS5COeNZIKm2ViQ1RTjRaECaRM6MzlEhphxGPGV2xK5
IhaSCdt/eW1xvdGrvfQNtAQ5AEmaeNW++Mk+5VTOnw8F/nP5UTO9rzAdeisg
hkQ8FFar+GzQhajuDiiY0PmOsHKiKQoOVuxQOWMowEDo2H6B52+1BtLlcz+W
/CrIVTTqUrFjTyC8SU/ZIBEwi/1hS9bOG27g1TVKy+QmgZjpkCyW5DNqkfBr
i0ko5UYWNjMpTSFkVwoIHkn6WMOFqYtX23giACy1jGgdkCE56ta/UhzrbfRg
ciIMgbMsDby+Sna4+cK9TfwmnkhlwPDzzylzjV4+Pw3pbEauoZhbWPAgsVAo
G85aTVHmLn2bm1Pe7tgwgET/qOKA0EIgoDGH96gv2HC6AyFjZKhyRKv7vA5C
9iY0Tl6TM7snzTAU+ZbzFssqJ3psF72/uPYjGz97A9Rkthfac5+kTtF/ekPH
r2uLRfYby9sK3glQCH66GvAgKISLahIlDucKASmQmn8MZX+DWzplNL5mGz7F
OczgaLmEWCDELWJ5WxdZzwElc7ZF3okEiAwDXRU0kWQ+FcU+RGis6FbleaSX
A5iFtMRpzdXtVzJ0Nerk45N6ZmIBS9TrBu1q7C47InlA1es3Ep3mEeXfW8b2
EhzZ0LBMT34qRVzqq+r142IED5O+I5KXy+cBb6nqwgGE9vc3jehHG3rInY50
gaQPZLDtoDDbaw0j/XopZTHL/Ule/Rtbppk8ImxRnaqYiXdSkrspPv3l33ss
jvI9MekcJH0UsAZkiA/Oj9iNo0E6A9b5BgVTIJbo28reue9/iDjBnea9Svyx
pNijwmpuJMkS+WiC2wIka2jE8FC7LvCn4TDPw7+xKqp+pFRgejb0G0IG0a7Z
29NNUwI97emS0OssrhLANhA2zlYA7bhVWa8rgXUy2wfegS5B0fFT+LluI9dP
Lz08MW3vvmrqTTl3RbViptxVNZQzdIIBLFTtydSkqMInK7B7GDupM31pnoXl
VonFvM83qzWe9UVrdPwAJsE8XL75TZgn0Q/mQ1+Ot8PrpUTtmokk5PITEUUS
bilBpm17tWU+hxbsBOu7tbY7DljI0w7IDdUeSwUAh+B3yIEJW1YoaLjxNd6n
ugJpOcsxpWq36CIp8szeUmYo8oedtfHt+p8Fn0uFILcuwHVdoOMWDecF9zRO
zGs1gAeFvEdP1KNIBQ0sugBszv8J2eGs2B1KzvW1mSC/wpW0EhpM8l7spOwp
Fz5mTGIOYgF2+Rj+XmWXeSRyehd9s9v49k5NVHoL5Vw3DhdmotuQ8evQbnYv
ftVIxFFUX7ycnq9ZP+foKfkHXWR6MUXkzEW0xxuEFEnSTzOOMhOuwp/B1/ly
hnEO93H4wv52nRDNO8lQ01JpL4FjWsf+Uf+LZSqYutomrDmSsar1BWQAOQYg
sRtRY1jDGb5aYVczH9GWi20kMB9D7YGGC84FlNuxZdqcTGRDZcN+voUUsPhh
hOcFCeXboj7siPfswXlqNE2ZpQnNLsU9NbLz1nLlWf1qEgIv65exvf7c3+jg
5nTNoySmVaXEOLEQsm2TxvvtJtGCRdonqu2p0X+4em1HvDo1IWvpSAWxzWh7
fOdHSJKRUOA4HwNQhVYcyi9NcBy1/HC2E7HKpuatSBQqj/3xh5Uigu6fLzjf
XnxCU+gmkX3e000FzTscts0cs1rfRSE71b1GDtpaR1bs2dA8iCjO/F/reZ5i
5MUW0OnsbtbLo7zxvABbRIF4F8gq88iipFijB0KK9MR/SFylUAPkmTuh3IdF
wcHzjmCsdjtgdldtzPZrk3IpfHJA4GmrsFAh+uHBcHXE3drxVe2GDeqnopcZ
Vb43Cv8TI/b5WaD5d1/RFU/e7kz+NHXQ/A+krT2Bb2EXh8jRG/rBTx4p6xUS
QMSYb1zyl2SMrmOjQDL4cYkl+txNw0zXr8Scj38fbwI4RdxDHWqZEGK1dDeD
jgqCDT/OOQCgul7CJP9D7ZweJk+wK1pbydic2ZMbUBYO0oANOpg+13xOeFZ5
y6edfvUqzYZzBL2g5csZc9KshcQf6b42figxmWhLyqB4GndRZOihzK5pGrAM
DEqLCgPViKHMJl7ILd0/FVICUMZvZs9UVwrD5MHdHnCjoxE9giWomL+a88RA
cgq5gJXD2z7kCcJPH9npimVyL7Yn+HQhX1evNYbRHafMeEkbkZKJxANaFgGC
a4gQiDznMSEAKNtgYKHq+UGYWdmCiKhS6skhETgzCEP9fRuKmyE6I3lKuNXd
o7Nxe5JZ8PR8ZbDBEVj49iReviVxInBoZdrcc4FKh2xP9YaPAoJdODWNENEV
zRM573sWp9aHoO9knTOdMXbP3NctEzdZdIIvKK7Q+4otBmRQ1p4fPHmPJM9M
/vVTXXHm+PNxc9+Ol7RODjgx5SFvqlIapwUHfLpE6jYc2cjvO+2NOQasMHvg
Yp6uc0fGhoNXxA0Vy8FDPRTT77DHr7Ih3iIlase2uoWEiuqT73W9Nn/XSRUL
BrggvSCwxVMCDAHOXgIZxzNs9NSItRBQhMGeXhjBd2aRW3fogv49R+hsFl65
JZsW1xULEaCEoAIF4NtNfK4mt5saGLQMZLSN9bLlzdVs8fjR4xutIv709zZO
rK2/jBeQvdQzSDm2PzshGrv6YvPEHhFZl+RYJ62kvJtmAjfKN9CVwl4k4KFR
NSweDhmIldw4j33AgxwcrE2X4wN5KaE/ZcYPyFmX1IoA+yHwx+vRifg6jXxW
VYXGfF0+/MTyFIVmhLhH1CXqISl/O34S4JUJEWzyxW9TqQknhQx7l1/lU7zW
b2sHMcmBEsoL75/ROIwtj6l2NvqQH//m4+au3tw6BFrGVjhNP0IXsAUY8snh
UUMriIiFyEGWQm0swtWpfrRthJJyWAFRQ3lg2pxtxGJjh1e3UU8qnkOhE/PD
WtspkJhaoec9Tb5ur0lecESWG52G13a84X0Zbt1sXybZzVcW6O1nWm+HapG7
l2mWs50Em8GKduA8AXATWeGx8/0mdME4rNfINAHMG7kUlmnDqXeEYWlorl8B
A6AEgZCrmQ3RiqvUKl/cRDUD/XfzGWCVmZJANcca164OffqpeQwRbDZSDnFb
USzt5F/4PSe922bag/j1Oqfw+geRAzuN6REtsUjxk7Stl3ZUxTUrmohLXC21
+jy5egKWdmuwZKroMhOR2AwjRp37ZqO035zoo5Ky/PINGYV6MWrqu8Q5EiIc
/6abYAXFRfebkZhritFOQs9fnK6YH7nGabx11vLBiETZHTVWbNlFtaDOYeE5
gJ7PdjDZIImuyDoMV0UBzkyU8GgBiYRW42dwBj62FktU66BY6XfYIJez7tHW
qQ0R7RKfaqNwa1InJOZcTPAnlhzhDEb/ULbASUtfvvZ3LD6XEaIIkwUFQt3C
OWuXPv9YvBC7XjOcYFSO8Rzn+/mDMP31dppqZad7A+Kbel81AfobbEcptf1i
Ob+nSjsHGf0dQ9vDSj91UdYXVlbj1RAREuLdBmKvPipFYH7AwEwr/DetYi/8
SVD36eJZwN3vGRAIxakEPSiOulZ29VwWrF7dfOJtF/xR8dUAAiEqXr6ou5k2
R/Sdl4TrUUfRWGoKlqJv8WoXnobeE/lybOPUZwmYrA+y4d2VpPia+l0nN6VC
FA7AN1QDiPfPamSiMuYqo9sMX4X4m5Kqc0k2fgJffcU91hB2k3zK6jmPRzSn
T8uC9FyU0PkMxNHF0MJ42QFZCiwIFvnvZWb3dk3knJtTMX4jj+ZUoY0G/FE0
Uai93JOkCHYzN9LVdtjMAzxU9/Yp4mGlK5ekkZ+qCkm2EyXj2rdK4DEfJaKV
PLwPeLr8n/9R2kXMpsuoYmGUvxSLyonj1PjHyKngSZ7yHORuaboLnsxrvy5E
Slzs7zTG+gYP89V3CZW/fjo9crWxz1M7tqDbWmXsT7Kc5Aj1uq/ZW9cYxURT
yXZY/mKjtbtgtGmxPPQHC1IviHwueRs8kwcz0x+dq1O8IYrpTSaMmh109tey
vsHhdfmXc1tmXsK1ts50zQrCCcDXwhrE/xm4kgpoXjWgDgjJixTs8kNjOdh9
U3Pp9Lwp1pZWTwcwITQIt9TxW7E9VXYOo6upKtP9nhlWy5vHrKrt7OYG6NtG
45FyaFjmrPjFTi/y/Oeb/baCy7oBlNPHQ2dVWifHvpCX3hOpW3/YK8hzeSfF
uCiVkgUE/ddWpi48CwabE4hp2QS27XZadllMrU18wbhHRIMxd9kAnXW55Jv5
FebXPEozQuBNBBYiEEpTM4JVmo9cEl8l01OhoMngbfsoFqnEWC8A73YpYSsa
mh3YKM8iZZFFsUOvlQi39uH3CeKzB5UVnc8S1u6GIZNdPcUO4MyO+kyCGmmw
iY//SPfKW4pWag1xvH6E9uPUUBr2nh6uryP2+uwCIBkxLUt2eUU0UrKWKo5B
/dkm4zVZNeZNP5gKgsvPBerrZR3k2xRK3ahKVr6h83mug3Wu3Z44lvDowdXg
AQZ7Q+LEVamJQXijH1imS/k6dXAinz81AryOujVUomNIz9AyiNXbuh2Cpetv
yDbo6K4HnQPaD8EEUA16xf30iLSt4wpEvdvx0lx+4HohL6m9cp3oMkZmbvRS
uQ+vycM889IKYcbrWSwrIVUv0yewwXog2AVc+L9IbNPudi6xoEl0mi37TFio
h8Qp0fSq4mB+3YQK/feJ90LdZCWLvOesjhg4ty5WjtzjAkn3yO5LSAlUeuJ3
k8mFjraPvPcLr9zpC81igGxMuyjCAyjnFmR9HoaLX4nBujtcE6uO5byalvH1
4eAjbth00TMK9WDlOvvp1PRUQuaf8Fs9vapXAIZtAUMW32WiCai0GXcVQipu
IBv2uHnNw6sXyfp9vKtpiOneVsNr4awKoFwgulDSMO8eOizrvRdglHxc0OIm
Z64PNmX0C6vnayF7166vtioOgVG9qfMDtZJrWYjcJi+TF64HDWlWTrehgfyM
+I0pyRuIw5L9wxbnPjNlUfszNLx22456T+FujO6aI7bvX/9V3Dkor6Du22B0
NoOQLJb3NtoRZcIqBpHtk/lylahJq8k/wQ9qw+rF8thyNP7I/dEPh4RuaXaC
exNJNpNmC6VgJDiCIP7M9vLdek2VZShjBrCLNc1Q8xrxBnLK2JJ/wLoBBcsz
Oo8VIyHVvoKmDWWkqVzmejFEZPBCDMUXeuWav7CAYUnjapfFRcguVLZvQ7c2
DuadqoCkb7cvZZosTkdwA1846NB6s5fdYkLMcObeW4pAbRE2ZGkhkpFVM6Lv
8qKxzuUN6KTL3eiZLYgBaN/amfewqp0YTmS6dtQPuHfM/80O8rAo3XxxaI8H
NAXNYFUJWYvbgVDGZ8ufQMwbouAW2yv/hLjxWTIkwsj1dBkkJM383+o6r9Nj
wH8RhLG/63xgDupLqw9RGwMZ1JrHydnkWuK64aqzOT7vt9ZGOboNoav/XsdS
kuVywOALuhhU+5qFORZL16jxh3eKEQJm248hn289h9ZMIXHgNxJGK3qkMvzD
jueaIdteXU/RSeZqUOrrgdJLSthgk98sxjPLnMgwdX3lHUe2EaQ+9r39cUDu
wiNq20cXT5pWYYXOoUQjcnmNQJydVyk1VtdO+qGJH/1uSl8/pm1pDjmHxoKZ
pyIXVMIRoi3KEpFMvEBXf527V7+9CS8ReWir4EaHFPNpNl0jrIOyReifWE/3
AQvQQrQyzwLTEqMvagklG6SmfU28cn/LfOQIrc90dmPj1fBoCjpTVH/3N/qO
Y7u1N2OyedY8gKNBHZbFUTsMD5qyehIfpTc5k9xytp+/ML/oA+rw30RX7QlS
xi77Qr5N3L0TDUkEaKzF7r1mQUaIteGmt18BGlPNFcJCtRqtcJK0i68cljp1
KXsC4hNvTbZSwn4K5fsY4t24SVmlk0X4lZS2hvuG6Ovl/92qAGAsoNl/WxOj
441PzP/kNUrOqojBy7nOARYkmB9/ibZr1YMfA+5G7E5Xp5XyXHqO6M8MyhIo
TX754XE43d3Dt8JCyjnrXkuw+tunEX1dDOh2JtKGODjJ2K0znCohTEN8/f5h
GR8UHgtytlFkhOVlAJ3PU8v7QnzZwXZeWABygNUkkyG3AwtaWidR/IRx9xID
IRc0EdMwHEMhsvakxmY0YPok4d24CP5IlYEpIoBtiJ4UZm6qtJX0GSzs4qKK
pAoBQDrZBQuKCkAMf6CUZwxP/KSPQ/GjKUdg5IKjJVmAWmqQSMoheUMLyOhd
hNsu8bipCUAB3liwmHQ3R/6W1uhhrFSaFPGRTYpo62D5SGObnqAUDaAr0r9B
plF2MYBRGEeAxLetW1xXnZHDNz+6PwuM5mNclWVXI6a39698GXtWC9nLH0AQ
8ZW6Dm5D6UiCGAxwazxWV4CCY59n2gFL7wPua+T7zmoPtHJG8NzZS97zAkGk
wKkwQExBtEBQjloehQ+74CyfMXbGENoIPcGUUrLk5IWFfGadL1Nb69QsnkMe
iFpdXFlmGgYterdk4BxdK8BCetI3Z1GgEtBhzFAYw/LwALUtuN74zPhZS+To
N/wfzQWc93cQZtsHI8/PN12CvX9Dc7NA5YGc+BT2gkALtPLBLVv6XiXTh3cn
3eopuaidwTYxnHNFQ8wNvyIEgVUsT2+/51Y4bZYIG9tm2nkREtsG83JONJUe
jkglo+AA2FLlBIhVZSuZly/9+KPdi0+cB7MqlL149ER+7HBypSjSfMHzZ1he
A+zT5faVafwkcO9KUWBbrroe7VNZ7yGcErjphZlZmT3zIscBKwRmO1NeMGjP
EvmjrIW1zkYngKVP2vvi4gaFVrvaOdV230GsvfUnzRewlddMgA2yDx/eyjHp
kz0q0MBMaQBG2Zw+haUqi3D6yT//cC2AqT2nQrWXDc6ky4EE4RiMnbtrz9RI
MmjKtnj1TthYuxffqTYoVezGy4LoAWjCULAqz/ZHX15jVLTuUlEhmE1iy275
4OBCXdjaNSQ6/Z++905UUFSdd+X/sKNuri1LJU2JhE0sFyPaEOKjDeDAsIug
qE5AeUJp4ly5s/O0BpDvpnjoZfPT2ssxnn8NHM0bUC4M0+YcIFh1HoHEhpOm
k/mD3YcUd9CvXSKx4xLCSpZcGh1GZ8PXnEeRdTux6qw5CTxDTmyxs1XUeOX2
DWuQTfEmTXbyi1tITCMWWc40E+/tBeTlKyU5NDB/CUcoT+AABEWobD098rkd
m0LJ8tQhYg3ZPPTg4+WzBrpET//X7XLSDRFKdyvgZ1IUQLfIvFAaNFXmforr
jKhUYs0VfOPR2BiT01qzefHv7vlV86sOiRN49k0gG8s8Ki7Msar0P2y1TTNE
/ZJqmsY6LZIag9UklFpD9T5RTmg8zf7c2NNRkIjR5ymYntoxxgGDmvSB8tfG
bSNV1ZYwOZ+NJT1h2vhVpirdlu4c7vT8U76QCL/nBd2PBNfiEVWt7UXWjJjn
ycEqdbCixj8p3ukziEk6Mpnyj+NSu0uJovOIC2MPNSt/pks8gXKYcqb5IjQt
5EHTCZ/fHZJgOliXR3wyqoJawmPO72hMZ0npkxGAkFHEGO13cBUSI18C0XRp
8UkUDgXwH1vxblLUEl3aH0MDd3NHKKvt3lIAgWE2GlXr3hWIftjZhXcjW80b
93sB/XP6ABJ9m5Kmr3zcsx+Ze5yrskWd0kM17AsC06PUXskCDUqLbCehdK0U
GVldv6H19Kn/KuiFlfssf1r9Y4Ztpkr1NcYlgfCucM3aVkRsvKIXFXa9lo8U
rC6CHDhqqDMjhlvzgjlmM/i9HxVYUTl7za2XmPsC3Qd0Sd9YVPiFa0Zlzzsx
jSRxPLnnXHwjtevB1mw7a3B4/rVQ0jQQUAU+Rf9LGhJzEe3TCOOQy4tLrQrP
pGbQ4Ifj7Iv3BH7Al1skFuyfCAd5OngBbl3YVC90LGh7Gsd8IFWMWrqJ5y5T
57ncQRIoxa/QVJ/N9z/j9H/wJpgXmi02kBsf82Vt5Q7RbroVP5CPgyuhzf4c
QJPZHW0AaT6d42A9aaejUd0cMJgTu3Ig9sLO6Dv90KgbEirRnhab2YKR1WDc
i7mZ7rH34fEcGi0WMwrYViTCMDCFn2p4Q4HB19+w9rHktak3cjj5KD0DCEKo
caJRQSF+rc8nAU+7igykOtuM8MzpME2as6ZTXAGNtn9fKDl+sF3kUnXGiZg8
klE1owesAwjizCoJYA4pDSAXCTUS6yWz5xeV/XVB2e9igdS4WXOrNSkbgnFS
YKPtSURF+jUJ7s19TTw2BhuCP/BGtb6H2/rmyMa6sKTfG6d4GzBaK+5Uwve3
rh/jgCAgi+NcJrLlyNOcfhO3EiubC55dWvtvcjAS75ZotGVXOEB6GVqbg/ZZ
1G0pcyA0VdfAfizaOq74n/VRkeEVRb+61GzmjmMunDz27Va9BooX2PkIb5Aq
DP5BdRN61B6+u73O8zdTSiDYY2wRGmaApVVDEa5l3JU6XWX7+24nmV7YUHf7
H/nbLNMQjfKozzU/fiQgltY2ET/dsgRTHrorVgjJQNs6W9pRVTjJjFN7xCOt
/fivjKj29ax+kzrJ2dn0KxemhVS/aWGrLdzb06m/RisVLpOuuvdXeezqlmYI
1og03fxXwsJbeemcSCLpA38XIh/Y9b9Y/Omt+/0o+4I94XhNirhmVF9SB7zV
DHcbMg4J9gYzN2mG93jIJhWKcSlJCyAsKp4O5mN/4qmEHAzBuuRXZfDhqBdb
9GLfyglbmZPLOQi9Lwg0i5ZlEtOrbbMkXyhQ7SIpw+FVQf81EduKFi7vMD/e
0KBGCl0yxLliUdKv5Nkx7pS3ixmNJxqd6fJrpVZ/hV46OnEzatk1yEenBcPU
P5YhyuUWFTfhjh3dvc/XN4QHDaquUCDHq1/gkmQpvnLsNw5qNW3VKJdh2vfv
gcw74ap7rWZaFZH6WUP10zIkWiFw9xedHD19412m0kIUWYz6vLe8xNv2UyxV
iBeOgZz+GhFDE9pmgGezhgyVvHKPNAczWY8ojTiIC0z86uig+Dy/nBnkkiCt
9My1XciP3nOBuzdo1O+ILYSYILKQcGeAdxqeV3IELe5wNG55H9x09loEWKll
UMwCUrjltj401CI4fu+gyfDQYQJ53Yr4BLkir7qBMFAxdOulYrY0/dRZScSp
XRdyp8zujFmS2xWLoL/Jbmoox+/0iEba7VrgCC/w/QtCqUDY5dKcH8HOdoh/
993sz0W1UTUY9sjiy+pHykDlRTNznphOnSqYbkvw046znoJMJBnkPHMfy5ni
lWJO1Vzqe6a0ygkH/aO9ATIhSYZM7vnHO/t9wdrLz8V9DU03EXGOjmWRipqo
XmfNsi58LHTF0B2mjV3URXKsKEeJ3joPItvTxF7JNZ7h+4mn3Gd/IoCTfqsm
WDk3qUSErt+WsRY7s77dpjCbrbedTIRNpHCjhuS/MXVdCwx6ac7SsDE1vxsW
iWHkaF7unGKCh5N4C4skMo0QXxpb7+b550Xs2KOcRQ+Ab7NvHKI1zTXE4aq+
fQaXYiqxCxgbL8WrHf5EG+vk4y5I2MfhDsnUdDjizOEJ/gyY9OlX7E7my/Iy
7AHxc7HrTl8UZwSq5165I7Ek2CdaJFE5X43BnbQ/2I1R0goQk72JTmgJHxA8
0vUaBiwYcPnPvMKpeNWsTJwZyFb5JTHeSh8V7iljdA/LVmQ2Ac6Frc8DNYA9
S+wcC36If7YJOXJ4h2o5yLLo98JpSoNj1KgBcm6YZhhs1Rqe7x62u4pk16kT
Pn0mK7NF3Biv50yXsONVboHBzfQqPJf+xHFlhPakGw9CuMrhzEhX00WoS1mH
OIf9bUsHa67n99eVINQb2C71OfgCSm4c114o2hsiOBmiVl5Ef6blRNdCSEFY
0Jd8+MDP3G53vjarzhL34GNNHonrQC142OnEAyMq4mfkB4EO/VsUiEHyd+ri
H/Zg6lEBY+5kBOhulAsO/gz/jHx5qEOeVXBquekeF5wJq+cBero02DADcNAR
8hfuWCFRYg9vdJM5GCf1DyGueGAp3cNIL2ezUfzdE32xuEsGoQrXDtDPo9UD
e1xmKd/Q+o7celPezW+CSx7DxPf63x6LtJlmIOXJWcFM7bNDEuhjHhPqjlvA
xixRbvZh1BMIjQoo03pwM4IxJAkUewc+TFCgvCnjudtkA/YaT1La61qHmypn
EhXGOOlO/nBSAdnM3EAHMLfFU6qGsoFqhJQ/8q4ILPy6MTqF6yqaqUhHSHmx
FabBgU6erTfvazxYQKlarvvGy0YpRlcnbx8MOB11szuyqNQRHo2i7C5QLt3d
B2qCWikCqYZSjGwclueujTBU+fms09jbFNET6aZ5ZCAhd49x0YgPncBetKE/
J2kRHvl/FGar+UmUNjbTgiOy57a7mSkyMSHfZY/ldyiIePH06JSBM2hA7rp/
9jP9ir+xt3Ob33yGwAtfjB34j227rREnSBOmOE+LFHQxA74Q8NR6ytqpopLO
6z3PQprxIixtTturZYJUfx/vbvbMWj3qbl2haIz98YMtzZ3nnBW8lLSsGbY8
dGyOMO9/fpVMEeCJZhWjqXeviXdtPsrwbf7fX1XunfB8OtE0sgfF5zk6myMp
zyz6d0WkkdIvokupSLAR5Ekql6ETO+hLfBBwe18PGudg0l/7pAXKK7UjS3pP
Zba+x9kOHIr1pFs6xJsSQwJq0DuWkzQr+dsPrYMIcktvpLkHdtI3GklikDdi
UiS/CyhrMGuKwZWyrnI5M4eYYwIPqOQs6f2OJPGKy5EdQpwMb9v8CwUNEJqT
aAjEAlFDbvQb0AYR7FStGvYelPf9ViDhXKDnIgoWFJmcV/UT/f8shddAYLjM
vwoddijEvM2Khq2Z9fLVU+7BkaBepoKn+D1rEhILcF4p8TJX1r+WyA6QkgPR
zON1dP7U9J7wnkyoluQDFz1vMH4emvYbkPH6992vT4bb5Rq9kal34VMKhmlM
kqCw1MlddOrn9MXxIqKiQmIS0yCvTMh1y3cE5PLBKDctLXvuEfyLQI4g2eJT
zyCheBgVIVHlIuqrgH5nwFFUj3hMitdgQX3qaNsCftyFumKbJOvGDtGJ9ZtK
q2nFEhfhv29eLTjGY/ea+lmismM4XR+/CaOPsn22fQCfKTUEmahMJijWuWFr
MoOc9zodP5bU9xNIJb2W3kGMC7S2yycWRk+nA+7XZNKz1TywD4nM7otgOOCd
mT7Nb/ZeojGXrumCrDXSmZrXEGYxcB1tOevDLNYQO5aCjmS+e9DjFm4tLCff
0ufWrucSGLNuT+REZPui/A4fKTjZBudTWFeoYVJa8NO1lvebpJ8k1OJvRAMC
XNIz3/yI7Oz2m80G1ppvO5vBVF2pv/NmRu977QMWC6me/loXDGzmJJ2W65ho
Za2DN8DuSr9DVtttfmdhZdsTZW+nYWOP4fr/VhByGQ5D3YCrMUsnQzGhL7u4
eatXVOM0ciNGiwfGKKh2BEyRsIl/9KLyMsW0NJizifWzYm5VOgTLoG+YXcnY
z7BJsPIL44fMEZ3o/gdzVRONkFt/79zedIaFzCgbFfBH47Eap9KzYe95GU9T
7O1d9qx1qKLP4JrmAtrUQXMwYGNY7nA0WvVJAXkpprIxO1v5eudcmGExbdhw
0GSMh/FE6wZI2TmpiJbw2fN2rvNPuk9FB7q2FO/TYMBTpWsv4et+YW8cku+t
dLM+sIT2SfQPwNyXKYgsbkXAXnWslRE87pYqNvTMUQMjO4B7gFFprg7+ngb8
yYsjosnTFSzEdaCmzH8CYTiM5ejJ+pcKd6Kh/DXtaIy+I7hpOLHohbboBY3e
twqhLefsiUj6GOVpzx0Bj+MzC7WGl/xJdBMNXvw9LvYeRMbmckAL6lhdI1IX
C9r/zEVBvYqFapODLWGLsINFVFoPF9xeXAjE+R1PKcU7rChqHMt07IFm9mY7
teFRnemKwRIx5Io64Wc1CeScRZOGWRlzxFifQnrlKQYZQ6dDJk3jeUh0VGJE
4q0gzHi/hjyio+sK6k/m/P6CUMkNqyJvT7N6YLlgGBH2yntJry08ESOpXNDk
vDOfCDzlJXW/92PfUaUI3IchQ61KSMA4x68Zph1b5VD5B8B4FIQkF2pHPvhG
Nv98AhpifLDcthOQJq65m2q9xow+xXIaxGQg/+mRxwbLv3TZEe3CV7t6Sv5J
046eh1zJzjt+A0V8QsfJUVl3qwIIopFwR0IjfaS4cl+7q/XddQjf9744duNK
0yx92F40EISORCha5T9q1ErD9aQxNmoSJ57ab82mOuR9dBA6KgKUAbI0mjNi
4ib3zndYBcHws42y4WqV1xH3ds/kpoCDaBixjaX+IdNUuD+yv+HegnJ+wt4W
p2TfQXFvenoX2YY+BKRLucFGB3L/Jcr1jCEZ5b0rFHMOKE+ApywjCwgd03ib
VT8nMylpjv1v8zig8lALuE6YRh69AtinoUicMMeXPbXdcdGbqjRn+tCrrXzJ
N6alsr503hd6WRMCroL2MSo2fCcTZ1/HV51w5gYYlCX2rbdUH2N4LtxXk6pA
ZIXhHYXvrJ+19nLcVWOUt0N14nGtkaymeugeUEE0o8hFdBfyOb3qfckaCKEo
2xMmAVAkKtnxZ3MKXdL5kJ8m6DmaMvgXQgWqI9TTxhRD2mErkWtrgjIbgh6x
Ie4Z+hLAH0K0UHtdq9DTjPxeSga6jhMJWs4nGFrmKoHK0dbjbqeGqk/JYxLD
uWPQuFNznNdrm4Wmt6VsxXrnInkQjy7D0CnqXldds+GxRAOCwiOARtElnU+g
bBEwBdKqpC3D4xQOR8ekNsDwOPy475AGzlDq3KDows+5QJ57h23yFFrSSRJs
/yHx7vDtTQXo7yG/aclxS3aX+oHDsawXd4uqfOh1refB8M1x/ZxfE0xLKq8U
pCbIBUZRHhl94OO+6gTOMa5yWE8Gu2qa497qeCv8Kp5c7XKYIo935lY+d/0/
pfF46mlgYgWg+HvVS9IBKQpQWtM7oq+OZ5soDguHRU25IqfB6Uv/V488hYXA
V5i22SzqD8o0TthIpvbRxsRH+5zy3GZl3I/sOrMcgg/3mzBJ7FiJ/JQxeuU7
bkzfvaNo73WpJTV2Bqd0qgrvYDOR395FWAqcZQwFmSWg7t7KdY1ydakxgLgy
ZnkdpVgdlMIuWd1+ZXw4351gqDp5kc06etjtAtvhPbbCQroXvTf78Hl0qUPa
Dury/iD+etTPux2JPhA2Hk+1FtZfNr/QCeuzYGZ4CNu9Qfb+qlFPHhjaUndS
a4X3KQ9KtVXf9OiNNi+p5+WsvkCXfOOs/jL/iDJ4ksnAyXmYzI+XahgYi+dP
wzeYodpp0UXilBCLcIAUVi8y+Qszmu7Q2YEOKzbWsPgPIcNbKylZvOGgHt0G
PJfzgmjt7zhQRNIBRfO10lWKGke8Ld6BDVz1/tF5eFK4o1z15gcoptqUiQkF
fmFrW/WVLEOW9zfVmMtDLqjYsanPzXBYP9HNwadsM6oSruBsNlhuOwbZglEa
MD4Upai26OzSFQEJ61JhB3BRbpaN1lCWIJMhvO1j9prrPaU3UpbxXF+TwyXB
mEc9Vqk1jccCvqUOvCae98uIE2nYfNk9Vx/Vys0Ahbwd6090QEGScFipoy4N
2Iwf3qIF/4owwNxA5vIzHBYiv72HVTXczkqvgXb8mNQYgVWUqGkXCSkS65LS
yHUXnwOTC9yOrwXakVQ1XTEDK5WKAaG6U4LWiBcLsMJyGTps59uJ99KsilcD
SB/9+L6KWzKjYZ2rpZIpl5db4sFMZx1aRqNerocCHoYWUJWgGL7qyMt5UIog
1b9OVdeOW7X5XzujduysRqJeZ4lcPjEtXKvGmym/MOxO0h+lkzR9Evgaxjdg
s+mCYsDoNNP8cOrfkQbvoVXyW1oZPtWm2jX5XthFHnikVcib/yFCuryxDyI7
1Jz+U+Pf/8pm8+cbGT5tac1zVnaR5RRxz80Jo3LUVlH/jS2TKGWvVlbdvgmM
nTDXbxXkUMJVvXaNRqpuDaSyjk4xa/1E8SLBfEGUd3oj30gkvyd7uasbdbP8
b4d9sUm5inChqUJlGPaNcFFcCXbHvvcsBFFi6EtlwCCJxNBW/9O+YJ9frKbO
DT7mxHE2B2JpByIvcgrz7QuVp5glEEHo7S9yNxQ2h/8Mjx1qw797vFHGNfRD
yISOxh7MA5LefmrMePL3iS/82ODxrjk+I1IeFTKl46kq5vs9gzT3324PMPNi
Ffj1h7NADwUUxWftcw4IueF/GljrE1iCo/dJN5U9d2ZFELQ4MPs9Tqb2LWFc
lXBWGN/192B6hGIkjml5aDueiOiM5sSRyHzsq5e01QHOayteIYewMVpAVLQz
XR4mcWqoVgG3X/xewXHFtF8xxMB56CgImZ4pPnxurzhYNgFuYpkXlTE6IvLw
NbTMtUtA+7EE/aL0SXmTz1lq93uOgJdZXISo2RGX+K0ztNGc3CPeHsqwJGhY
2mP9d7qAdc+x4Mnth4wIQf2ur/mXn4ogUwJCvJgr3ngFv4lxOcc2QXObBJOe
3AHGgH+lFEsFN3aFKNTGdVfgCfpEvnaNFeJILTrR/O332IXNU8AfDqLlS9wr
dZzAHdHimGWc1BNJkX63wd1ptvuaHBL6MQYT/78Z+kVhPH35TCKEZw8GHveG
pcr0oApe4GANveOlRlt6WFGBxDlyowhpQ0Lf7WTs3KQjkrpubg+e+9ijFueS
NkBoCuFVuJcJJb+U5mbKt4V/UzDh0xkyXvBPr6dQfCe+YFt5J24x8FjV5mIs
Eendot8qh906aeofO0wdJZVZHHInj03VaoVjjKDaTEen4JtLF/4hWx3ujMNw
XQE/FfiJNd7gXObDSPjpAcawwMtOt4GSoFXKNvLyZOWdtmofUi/PItmKokdB
zLXXa1+1vQ4l/kqtZxm0YEuGiDLHq+gSpfaTbxN1cyKns0vtcJKoPnzchSlw
w07pnvlSEKvGSz7iiE141GzkiVs0Xt8TPopxDeSAGJasFN6OkLzmfiKg6uVr
ZuAn9b8Kjr62cSP1zmR8EuAbW/+svx/8zK8lalHAE/7FRg2yMWodEtGxzSiN
bfn866l9kORO4KR1yU+FJLA4lCvr6ITPj/gLDRL0t6vsu2JkxBpZnKyFXBlh
C5vyjY5lkBiBJd18qAQJmEpLC95eEbZS0HCFc1rVCh5cNLi5nOiL2q08X2Ij
+WhUN+LSmSX9ESuQer+KCOGG5fdUwoqaIaehggnZL2DKa6rgeakhHj13pLvL
WMpsAdQqyfS0DEWnrFXikF9oWq+AIAKkuKtTZv9mV3X7sLsyFbuN1rnzRONn
XVAcOAR7uDJU0McKhYyFWS5QFiJGL8pTW5bV1c1VDhUF7qJGPeGremp+pKlx
REQiLNyqdrW4qbmRAX7ksouFf/+Pm0kiB62wgau5CByA1IyP9kfo/g7ZF64d
yE39zapMqfvQXieU5PDzELrOW7Kywrh+gK6sso5/Tu3ehgCbf3NhHpuFzsQ7
gE08Xp+U2VAl1d96/3/dnSXvDj2yKyaRnSZa1hr0WpsOh74Aw2AC1jw12WDz
unybg/l8FrOPcl64SpT7PsyenS9Ewwwg3VOeZlg292V2EmasKdunofYZpw7n
EOn2v1wg8Hep/++O2oSfYmY0/rR8CZ/0iHvnHR3LaG22oHRRfjDcls/14PkF
nNneS9i5N3bK4jZjiut4VxbXgctMhJ3MlHhFCQfj2EhATe7NhiqfMlIpHJqL
rySfjViMcAHSy7N0DwptE7tsFj/OKoJISBR4bNdd5FsfscX4+YDAoLuzxyXw
HYwbx+455lbl4o4ibH4xGfef1r1+cNK8iLVjVYbJ8+3FVb/hoZWTkHRo1pPH
uOMbsi2R5h/mROo0w4M+XNMcsN61PzmK1wLQG+F2OXf9mESjfXm7EgfyvEJS
J/ZC0cFPzw9qMd/zDFK+e/anbSjr9BdnN1tR9ODuGnP2dhqC0eYx7qWBANU+
PB5IhrTBHpr0UqKkds5r1dov9otluPMuwMNAmmp+EcZr7Hbl82xB6LxRkkfm
xHalpQJ28ICPWdvnAHYZqbucKTrcxSvIHjIRSroNjsbPYNzn0vOefVPWnEeQ
HSYWA2WX/71c8wkp82/kjjuWqe9IO9tSGGcoLe5GVpMwfhqj/IqpGw+qI4AR
gSByK6Br+MfBdCaHgrJXZzpL3bE0/rRJbWra9g3WjQz2UP8Jl+Aic//+6fI5
+v3aeG2jGcPXfWgm4JxKCXpIxCoao/YPRwu1XaXagi8suxax4YCfesKB5ZY4
FqAXThMfTCF6ashUjnusjMV8po3a3kaxWazGg4xxDlpdqqac9QBtdH3E1N9I
vWIFPx0fjCQNWa8PQSMq+rNqP9BKboSSWyp+SDV2cs7mgLH6SNrbiK8UJ46E
MKSvaOOls3GG5FF13Zqpun4BI0dey0IOprjvuHi12Ye/fd6S30jEShtJ/2va
ESoLi0ZSwkrIbXWxyvoZeJqNaKwEYi/m/N+OJO4RPDb5bcux/VEAwrfky38e
0BuZ1yj+LtZQ6msUIurc/jsMPlJ5TH0Mu1OuCitbA4NJs6MMSxgXpq7W6Gmc
83zRYCVTtEeRot8kMuW/bvL283qj//uPU26a8g91cChklDeWyJLO01dKignS
CDfO3OU0viQIAh+9+5k3OILvcPArDQb0daQRQud6hbrYFmgXRQ9Z9vve73AO
9evr9Fy3ti+FYs1keSCS203X+t36UbD2JvUkom/hJHCS5e46Bb1o77dehOU9
jH+3CSJi/lL2oKsgg+haTx62flKjG17FN9uuTojWKtFn6B/IKXvkSotxyYmN
03DRjCxYfsgkq/AJZd8gqHSYje/UUcVaCeGS/yAR48RVYl5c7I65mlIXcZ/y
RJs9G8gJNvAHEvBsoUmc5yFSK5aQ69A7UbTSbZ5v1ykGN6XJcwKBJR3KepyM
i6ppWEnRh+QmQ1tvWIn3csUG4SWGvetszkcxD7gYvKFBH5zVv/Kk3PCirkby
Z6WKFL9aV6JfE35VSS/LIq3Uz6TjAQYPVwEZkEuMMTl2dFItmCZuScKWbvoh
0tfUQkf1W6RxNPsSPi3Lx440ikTH55NxOZ9nABQS2Ra6AelDxE1fFn85S2W8
qxLdzt/hoN8Nq/N3QsHDNi4aBIzoX2zj4oCqaUF2ndy6fK0iN3Y5aEbIXac9
Wa29vbieKgrRNa/X7pb7fYP2Ua02+jkDETaW5DS1THN/nU0RbyXGAX2ooyM7
mysEsMTY/ouRTKjCf0PvmzZPGBR/7SgHXcZWWid18vJx8z1PHAKrghzWlYmB
8B3JFaWeiOJ+w84RTMdcCuAGl+/BNBpIuisd35XpyDVD3gpfP+haXjmkc9pr
+wf0N8eojLLEVWqRQf3tsjGSoEfKsvHLVkkKXlGkp2h7gUj9/9PZHiAN0WwA
y0t1JjDT2/xCn+QbogTwhC+KrQqxC2eyz+dFlLl1+3fDFs9xfEi6yn6Nq+pw
Gll875lEXmrq6Bq+Vr6vwoAZnTE+KNUXdDUNrTBYyox1L+ItqL5cVaXVwAiC
NxOZ7hHdej9hhRR2DN8v0+ovVJBgLCaP8uu2c6iAjL6AeMX57J5TQq+wM9se
gbEFdLjcxJkeR9oucr4Q/zwdRILq+S2Nzrzhyrftr/w47TRzOt/3Xy/umP7q
WSGWcyRNPJxHb9iG96ZOXjc7bBzTKVnygKpoaPAEM6dvu0qWY4+Gxtc8j54q
SSxq59CQJo7NRk+vZLCc0iVMSYHVxtAlLO5CDvq3SxUSeOrTqhxf/qO/DA25
UI80blWHWvY5FxpTV0HOqmBmW3nB+TGDKOiny2j86AMUE5adEmwYH9AaJo7p
ehQFkUXHz+QjbsmUD+cSIEyaj1x0G/wKbaa6idATBDOp3rsv5vHm0fR/3bOT
0ZdIWjR0gJrSwAs2LSpv1TuNueMXNWmkV6SjOX/98VmPuvpx8WT3M1+NZtmx
5dQshcenvWikq80evlvKN6lA/mLmAN+2cUAPjkkyDgxjI6KFKwqqNF5WqaDf
Ui/qtELKSp06wAqNuIlPTz89EYb0xbIm0r9VaQSTt/PHkGl30Df0SBk1RbMh
I+6af8muHTrK62LwEKJgCf1TmAVTAlMXOt+5u3qmCYpbxCexuKCGEacaKHfq
Xt0CZfG3pM16QxXtvqlA3+jwopPZhDUlNhE+p2HZH1V0nDdNjfv/DvlPk9Fa
uolBzHlKkw7OdeO9YuvoUCm8FM0N5fRb0YtX6Dtqbzh8Jo5Lg6UEE5860ft+
B45tmXkYH1CcBrpmZVMnzBEJEwRrOLH7kjEoDV8reAubJyLUh/N6biFeIb6J
QJoK1QszbIlBM2PrGVqNaMa1dWUp3/P0gvhlpAlmQGqG/zS9H3PGnfD9RaHE
4vhYl3kUYjMSHf5vLNZlQT7kpfNCoqGsGQDJyXjxRvuhL1Ggh6ajmryeJslr
GXrSKauaJjmAWlPXWp8LGMr3WQI/mU2QWwYux4dZL+0c0sjEML46lbBLH+ng
8rwFs0YUXKXM1DPd0C1Cg3cpC/6pEFXj2Kmkiz0IrRY56RwMNY9vc0DIDMDF
r+Bpmsvh9rjtuUi4RxlMFZ5NrQbywx1qPtjwGYJCemeOCP5ik82ze5I7Zmtm
wRy9aHkqO6548OgzJZrWDOnKFToDNccsD4YT4HwXXZ8kTIfOFQ3sMZukDCHA
2MMAAQCziHmNdJ2L6GfynOoa9yN66f5egZGLmNSxGFSqz9f4OIY488AF0y9x
XiTBlIUPVh5B1ezjLxVTdf1gzWl4vZa7xcO6ej98p8SaObpT5nC9QXhRQvXe
9jq1y0hT4pyKVyahJUe+miaCa9shsAUDI/8K2+15RG1l1RHpLHl8Dao2OsUX
nAZ4DoqXwUbxGzrnef1toK69grkDBH3HyDukYsFF2FfQ21nsHs2WdvoPwasA
LLDFVVax6XJEreqfjOvBhnuuKQ52FJrp3yefIaXiVzKg8VvRa1qtD5eVVp8W
pMsQ9QvEh5+5MLH4TNIkZTo9lqSaYf5SIvlGZ3gF95U3zXuIYR59/gNKdK3O
pi6DyC7ZnCQXkffnjKRlJMiDEqP34oVqJl46YQ/X7FG5IR7+Hiwl8sq+dzkg
9b3CfArq0U0lf0jvb0rrunywwIMGXj8jz7tv6137dui/DnCPmoFAOeQ2bKHy
cfLSNzn/oVjv15Ua0k5iUHB/IJ1CmHpkvZkLKND3NdZ7BZrQkowo2n2RPJVt
evv8ELgTm3fo/b79D4PZ3IIjnPQDYj2lp5zYmwWl3Hewz4ZNmIfb0XGK7/H0
0fy/7ck2XUlIooAiib+E+71xgE+YuBB6ATpy0cla6repDpiNCICMto4W7JvV
Im4AMOsLQXaw2uLuATbxr3czRVgZNeR2q4L3QnphELYt4B/oLySs8wzJK/8n
NBb1h3bnm6WpdxFEhdBoGKWejADlTSH+smLXn1n266Bb8Wrv4oCKpu5C2moe
GwntqZv1JeeZ28mZWyWTY/qOuBicnguq3ejWJmEkl8u0EXKqfXW/3KfhFL/g
KNyFnVDRbtQ3MD/1yIf7X0aDhMNXCeiKzyozY0hLdsotj2UX/EB+0LFiYbaI
wNXlNsrer1bUrBfNX71BJTZ2VEG9N+TnXOjYDwW9qZGfwGYQ3ZcVIIpJox5r
6qjC91+Fp748S5OwuYGZvobtn5QOCH8kYYymCWvLVFnGtBfFiTlGfC0UhdN8
BEZFTMEfaBnUrdfOwJBI3hSSBkO6EcCpIz2bkO+DzTSEJv9wR78QOwTpuDYO
jWS/V5evytxKDjDWsfRsu5InsZ5tSzz5YbHbyXEFQlqq4F9g22ZMi6FvEm0a
Sxd2vZDHRnskC3rR4msQLb6NvWeB8MehSBi2zjydckdsFd9VqYXaQLyaGona
hhSTBJ6jb05xwyVR+QWq1ycoHW3r55ecH9h8JVxYzCBR6Y79EsIUiQNZamhE
H0MuqL1iCLyl+fTpLa19zbaXeY+jcmCkyOZGVE+0kesD1wg3ZtXA2o5mttdc
RGCCV1GVSli2lBQ9Jw/zVRdHAG2w/EfMgC5ciIery9tfZ+a2Q09GeoysqY/B
oeBRnFtiny68GdpYJzO8j6O3mpY39v0k3kmwQh3iwdV1nZr33AyL8GMtw4Rr
bIvcCjrUBQY4XAbkOpzJuig2iVVBLKKcBnvruM1acy0cqr+lUkfSzPal/XXc
zYiOw7QpfkIDtq1TF7tN8Tmvv2RKNt4s9Sl3lnzER4g7NHRzb9LykCt4YDU4
iHVG7OO0JCT6yHYBSfAWA1vfa2teGmSDhz/mNNrTD253CtxFYD+s78ERo/p9
jbTiI6bvWB2xxjUCl4MF9OksJ6wBwLk7l7KjiZ/z74+OHYLRu97k1jdpjHgI
9nrliAlAl9xlfjcGav+7esM72FtcdIhcSxXJnUInUQ+vewxTtIftfp6BAUL1
3swDb/5+nBkNETsnpW+KXO+XTQu0ahNL3zO4dOe9JHvzW93f+8W+ChCRk9IR
2dcZxxQJoZU2JF/lYAWdvm4cB1P13xyyQo+X80Q9ftWhH6YFp9O8EsL4D8nH
2MgygM2bZ/NBWAkKfeWCY406ohFDK7kjhWkqzerc+Rgy3bJeDieRbEBNuHij
aiXtkng29g/atEQvPCYxPZL4Q14NrkaqU09teF8IWxy0cZ5WdWOJAt1BCTFS
nggIuStfhoImwmm2wYcxFfII8WPsgySytDHm7KdcUqnA9352WXytzX3iK3gk
GmDwR/JXoYg9IfrxFPCPrRiKp/86hzleOe48hNdFeLhUHN2N0BmUtOEW9k0Q
/HxjMTQlmZowr/luqK7ZAl7crbdXG5BPF1yT87YCgdOds+pNB4g4BmFcawI2
J+C5MXwSHjrTBdZkMXmQt7dzBcsGOc2K5/lD1PXs7Le/Ukbzb//udbqgUTwP
8xIe8xmnAAYfQYumRrugulSf4WSwgs90+hT/l71FZ6WQhPyEJl5tRKgA8+zB
vQCu2HynZoYPVgw1b8e/gmOLI0kGdCR2FUVRt+k23XZzkIlL4j5jw1zSGfKq
CL6oAv6GgROjNH4Ut6N6CcBfJdJelweqCIpFzlimLETlCPpsmP1qfRv57yBH
p/AAAhXuAGCDlzL9Qr/A6+YKkcbW8+QggbGfNPqREwoylJcyBeXr0TJeAQFU
KicOPqPnotDuCmjmCT9ToV8C28gNbUVWi9uWF7PXj6D5FLz/CcHpY50KwOjF
Vsw0ikdX+UfD68o5mhTRbcpw7rBbujgPMD7p4YeTGXD0aU4I54IWcaiMNyoy
6oWmRVKBDDlzQzBwqOrmHS5eO2P2z8m7xwNiYFjwiVyUxVOYWGDNJV1cuXv5
28r7f2s5C8sXm+EqbYduOJcmYiVSZCOTXLTmlIGmnTnwG3T8HL9VU5Elhh9F
TeCSzobzf6R85czbFp4RTvHINlvuG2lDK9Z8lSfUXIJD9OyvhHbzvG0eO3Va
z24h8TDc8D0LbhY+CX70H+nk0tz9w6n0zDfnN+8f7JzdwbBBfOtLzzvMEfrB
5lARamT3DzPDAIAg/k+nfe9u+Qnx10HZR/d8tryC+1ifTRO/GzEHOyEVs+o4
E1KoV55m7mw4kjvoaJx+SMGkvEU6Vzek5eV9hPNr3fnEjmncK+bHVrgeBRSz
RQSENWOIpkYmIKgVFtQDkHflvSuouMQ5wCvcco5q22Z3WESKEPF5HhsLrWw9
5f8TK6Bc264mbarzYHV3boM7Tf50pq6TyeT3XMfmFfpaNy2h+IWJGmqVLj0h
wQ7d0vvO/qgwvk7ZY0C1RddAX6EubYRcVbs1kEXNhrS+BJhT2t8hRRQHI+pS
+CH672jSN/lUr1WsuZV22uronvg6fOcF17aHfjMLKpU/QcwRr8ZC5pd+ucpz
3LG7DTlR44Y2htTJGr3PWgmxib+emuXIlubXZOSWST1AEssXkxdYfG6vnGvX
bQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1K479AQT/oDTSAEquK3Px12zpVnDfpNzhmvPLvgFywyiIaC7Xq5uFGOEFPHOfI3BuH9KGBio1yzMwBFDMaCwJJLZnljNWd0XIBXxcxQdeazvc3hnsxpSF7zVHznSJrJKTozB8f/LchN1L80OlJi1eZqHwP8KRTcukKHF58tCZkOHIwtvIAXBMR3AMCL5ybmkGxEXxL5GUb/FNGI+syDYTcChOFx8o7AgVNo3Ok/xxKFmZmO9D3BKz7juR5PU5eQB7zUlqdwaTfySJ47xdxTbdHSSUpBqtsajKA2oAsEDvKoALvXIxhHBYwU0taCm9Il0/cOQAU++GTP7SajsU6znubhP7RA3DlZRdy03ujmgGB0DsFV2K2S+Lnkcry0BYneUgl0Twsqg2Dx3jnG+JKW1n0uYdiceahtYC2aTHTWLi7SCJXBdw9zxD+fia1F8mpkAZ47dV0OApD/WL9kAN77WXgO0Ks2Wud/Wxm8VoHCfmVcWE1px/tdOwvwA2CktM/zXMDHGEh1hzCfuy/PfW0iYyPj4lgOxa0y1Ylm8YhXQ8Vo8RrWkOJgUanhaBHv2bb+PvnXrzfWG+Pv8/BwVP1EIrQTevoihlHxgLYJmTEYbx7VNSz2nO/3UXiDo3jRgu5giVTD/2TRwt+svba3wR74NH3YrDrxJysN/Jiv59c0lyD0LEhcKuQxdoUEzURKdbnmbiXFOXsbwHFujspFLqpK7AfbaqVwTX99HgUU4bea1d3jtV8cQQm6WKNHrIg1u1Nnabp61ERpOH7ifRmJDS8e9Sg3"
`endif