// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
boKeIRrKn5X1JtcqudHNSya768hgrP+Hw7u6mZEWn/BDLy4Ik9jAM4pkOlr0
n5Yd08U7ORgXa56pb0xGcn2VRS7kb5FqDx6wHUWOiJnlVS0RI30d3NZHexYJ
XvrfeDMvegGVA7qFtgceLeK9nq/QpiTvbXRBQabjZKrSeGqZVS3fnsZuSZKj
caxxGRCIFFdAMGybHT5W8FauTp5AHBOR2YLFCDpNIxpaT4eqansCWP6pYG15
6ExixXDWEh2q95WEHWD21yxZKq+JaiMJTey9feRUq22f2itfn0/0Wp64DXKu
fBNBG6WuAXLMPJbDnuKCKZ5KLWwuIsD67hDcPpl+GQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nwcl9WzTN/z6qwQFxSl3jUSj3uEA3GSCAuNU2huec7Z4xhycmTrb0lZb7Owu
QM6d5RKOZ7QSLEJCj+tHkK/LQB/klEIOCClGV8rEGe4lx6+ggLVmMOdoROG+
V5++Ca+WoYsFwmbby6iMU2QDvNYOYtx0g7ClmEx6zaN7xDwUHvOOQMUyFwLu
QjytrpdZwNRBESCpybpW0XRh0/g6IbHo40wmbP2+ZsM7S5QqknKpuBHrO/xe
yoe3RDqT+sEx3iyuXzih2juAuDNIW8bIv7958kSKalG/6s0ea/GiuCBa501B
O5oIzFhJsEBvFchScVJTOu+AWVPIBZiwxXNH58l6Hg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VczSf4rNpYYXj2D0irNwnbe6rx0SSy/lwcupUI1ppCx+VzbxNAyzXKkXFvWd
IyP+6faU502ZnExu9EUcp2B4bAWm0Gq9ZESrFpQQbSRV1iB0EQ8piRLSLRLN
ACbNYKHnyIYmpCt7Rjzf7kg4i3VtLxq55AOn28ma3PF0vuiqJimx74Bs2Pys
2Qtt2Ba1eeVneWvXWKBKsBmZwYzD3qHTP7Uaj9zy3ygk49U/j28HdEZE00eq
PC9m4j+E8jXalYIOPBsQZkbwiX5wANhmRFXCoHRsPNSimbrwZVEomDbDG6Tt
lF05JmOyU/jKawo0BS+ZtxQqfOW8whasepiWQxfPTA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Sw3nuSFFA4nO8AWLD8WWiHz0yPiQKkHXoyg7JpQuo+3p4FjnhnL4VlciWr0X
PTX3N2dgHXb3htxvz1daQbv7tpXUuIVA+44kI/rZaL4KQlgtPiSrlaqTBpnp
KMNMVNsRSl5SQcqVeY2tpAvQ5CVizJZKEllJT12b71PwkmxSrOerryjhutXR
x1lgxBCwgVJwCZIg014947R/uEKsT5DiCEGXQEuaMMpWNiMskOc7OP36Zcsb
chp5pgC5L4XLWw35oUNkkQNC6Epd8ge0mwVYlyt6SaUSx2Oq0TuZRkLJfJh6
k1BxyNK2k6DxdI9pOIbXCWp3q9NggnAM3gIzyZG7MQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Lfw76Ve2cXSCmt3OF8q+lD0W585aZ0E0tABStPn5w8r+jqfFwnXfZZWJUZ58
w/tJ1LC71vh7Pg8vsBwVcjDgfyekEMs/qhLRiQCJgxVtQQhkP0dKMjOlEH7X
bu7asuhbo5YnVyVEINLFKiDzQsZZ11k+MFEtKJANgfgQ1hgUGos=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NdZT7xPuGqfdk8+krnrdkR/GVwbZN8s3JjdAtxQQjF+VKftMpt9HhFnrPc69
m5IFOzZyfHEfLMVAiHYZCI4fQ/J6l0TD2d6SUAfyIAsy5BrczmEeTu4VdC1G
nib6DNhaWVvZcP0wzgiDRKNTraE42lRZ/s5os2Jpfo6FEXyTc31fvj98RFWV
4mn9j4B3+xHUXA+Slj0S3Y4oJUyK1R24QGvO+yxnTiBBzEsb6+THzC+7GUvW
sx0WMz/vjd6zYczh6jRW/YtAlvUAWnCGXlwYbvOWPx/NkXkE7FrYyys//XCx
xl/Cgebd9KIVo8ZIRnWqEq+d77cMSCURt9xwIz0sTT0Mo2keEgNkSzz0MKgx
lxExwGNrpw5LliUmkHIeVdHbmcFHdFQgREmjyviU8XE8jskHZDuKKHK9H1CQ
nbQbrOWSOtO8qVX2UGwhvoMEDAln9w3F4sZjj859eYHsZqn5mqxkCLJ/oGIh
ZL7lXyV6YBovV0RUVSpVDfP3+z9MM++t


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QIqK4mVmguvKVSobpE+dnTJZpwZSvtMQ9tnTLzsMoAeHMPQsMGhau01QMtMF
TyloOQi5mQGtrWD0Q8eeAnUDxtTuTNLn0KsMvkZsyw1T71/CAZWvtYdSz3vs
A3xj8sX3f+0t/wokuGOeh3y8JmcpMdu5WPYf7yL0iJCo0TmMgqU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L3ooGXZLweVtBctGWs8xVQeZ/bzU7MFkE5SSoK5QxveRCmW5v+XXtd3NIvH8
YSYSOsYleST4LHD4VyBG/VV+3VGiw2FEQZt+pr9bAsTMir1ENseS/Ce/kssD
7uuWO4g64ULhdlbkwKalINoFsr4dMaJoIoORsDWJPjYfF6sdG2U=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4448)
`pragma protect data_block
pOFAW0byIAr5CR3ebYR0CiqqjGM9lWHUYgQw1PCoM6IdCYc81gyKSIcvxieU
qVfRmqRrSO3hoHEOK+I2hRs7gDy6R4yco7WjQrU/hshC/VIypFtUUYjur4pT
HWMYB8/deBKsjdpmA3DnWxNGYW/YJfg86EZidTFjentzou5WQ2thYWuJGHbM
oW+weIQrR0+D6WRmeBIxTuXtm++yfIswVruxYojOPQPsxbD24+m3HRV1UIud
f3nFSx5S6cW8C0he6BNtpT7lXCvHjHgc7jC3yB3p2mT6p7XRO+MHIaTq7NSR
+UiendGzRox7kAxVpwcmxPv142SKeToQIcDLMfZwcLe3JpZ1dsZLPSDI5JOy
sxUyXxYVHRtbH8L+6bHCglmZ6ocrSqaWSClLTKLAug9jPkpphnC7vHc1rAKh
86AGCrM20J1vFDsVRQuq1edXtLUuf/no5DON/IKRjdrknRfwUjTtkRdZHqZV
T35P8QdxjgbeK24ueLxvKXdKi7Fj0sdYAJs1PfDGW02XYKaYdjHn+FZjZkae
FsWXoFeepr8nUMZoz1auto0VMFlVOmfH/EWDfnaLYdDbG7jLMvX5yq74SxVG
J7rMEioe8mKbNBlParSIx8AowikmI13MnD825JhjFlY/EJ8NkhghWX/l0WaM
Nu5pVdNygWTigyu73Phd/raQ38P5aR7mBgOLbQ45LNfnbQ+Sm3rSr9JIgoYL
I4inBBpjPuakDzLlJoV/76O7NQbm7xZ1PHQiXC1fgPBDTMRZnRdmZPvLi8gB
0xISIvlrl8BUslLxE52pPsK3Kv+PShauzCBEa9XCXZKV+n13MCJVkvAAlBPJ
CVQxSc3calCFxw9Q7ON9Fj5rydBpzdzRu38H7jlE8DcK9+8GX0r6kr/3LSfT
U4SJ3a/jIsRfx9H+mGI5BV//AenQe4ugwiq90EiTgueQMtPAgbJ77rVp+BRh
xSIHboEk8AbnyhK6Fd3CTB8A7QktI56pZc37zbFPYJiSmzCkTnm3/gjg9ZEb
JLUFWK0AZ28XCdq6xgVr4c+3tLmX/3cu6FPx7Ha2An3oGaFRNqp7hqmklDxC
0je0RRF8prFs5qh9TBfHpKSZmQZWve9PqzzEZ0LhqkHNbF5apH4SXrq7eYuE
+kn8Pe0dUl0us1XZgHMfZLJuXSutYkefkmAFXUA5ktP1h7OGdTbcKGUBtkAt
hm7+PPidDcaLvAOKbX90mwtK4Zs3tlv9FnTHUNzOH5UVBxCSx+G4IEhVZggl
+KW0H0g6W+ck7/8+gfdOpUqvcDqjOOXA8gLqy4qMAdj+OT2RSZzetg6Lzj9m
+hifw2glCHJVauNgLWkR15DlDFjBTqSRQKbwGhOXFu4o33BQlMSBvH9PvAug
UUCp7BRBZUKsgWeqmYg7370+wBFklWo2KXT9hyle5vop6w7TmwLsgUQm2A76
Q0KBn8ScrG97rltjSRwh2UVkdMh/mWA7lacKPtmHaabwxVf6Jl9SNvaPEtUE
tMiE+5Vfdmf7jYq/oJOvA7pLMHed2DfaiNsjkX8Z4doMucyRgZNRdNXGYTxp
UXJ/FA5NeSi/EXZCDoE6t6rtMNgoP4MnNCEFARV2HtDRVDsQ6j/Pyx2YVyhZ
firpi4wAR4nFw7+/R+5QqTuHvkCaALtidirqxrov/rrq5Pf2puVf3KcLtiic
d/LTF/JyYQDkE0SWgdTFJ+eTlB3l7DimuA3q1UO9fU5bKv8NgF3yyKW8wyh0
YyUxswzF7a6m/7+s5recSol03IGYD4lI9McRRkzINWF6vXyoYi8Vqny/hyth
AXckURIoib5hxzqYvksquANiZ1IWzjU1SH/RU9sa+wzIDmE0IrZQ5lIa2jU1
XbeUi/FtqKXiqf7BlwcvKjOAsT0SZnvyGArMeaX4feJOklGiB+BfZQaLwn0p
KKGMj8ChodvHTblIw2jD5S7ffspibg6BHjZ53Dbn79ITHC11N5ddeoE1ZCjj
jfFzZPUQI6VMT1bK2znPZBTUjr8AjMdfROAU2zSRnxDuF45Bd8cjijnUyKgb
wbBYeuud/jAwejgh0bYwabYQKrMZDTZX7iWOSKkqMDJd3THgDM1Cs36dHBBj
cpNa6lVb+77zVmyr5agG10OevTbRD0ndYgz/LOwfWXOFOyqBwuRXujc7Ixuo
yNiutFhZS+e8PHjeShZYoMUY/4NjxqPo3fE/BMglb0GFYs3XP5SVudPh9h/c
GQxtG9Exg3go9TjHhOVyXUOEIfcpRv3xISpfCEHKD1h4G7avMYezaeG5m/zV
5LFAuhWbDEsqTHWqLMX/IX496zLnix4Lw5Qj+h8cTKNoYYvGl7EihgAkzYuH
Ui0YaGoOWKhKfSy08O+oE7YCB1lDT6hcSaK1RuIMt6qorkOJwEHjAzXtVarp
cu+xXfL4NQRJ5CtM6n8x4ycrJ9oVVQSTIIZ1yxQtn/1uOHIxBN9r0+ZMgvSr
BWd7rXl/jOxFuS0724SyC2Taan7ArELW1RHpMlKom0GBmsYGcHZCInftj7/e
bHF077X6QI/azFcUItPRFpAvXiTWQCuiRivBJchXXq6Rvzmv6Sx/WX6Svmc/
be2DVQrpH8+D0cvHcuDal04EYyRSAbN6mrSMtrpEZv/p3TeRXckm9xg3u+Wy
5iuQmJ4n3MU2nSy6Jbf0j7NAAviBTjMdQLAuKnlBB+r+IMkAQzvzYv/1LwTE
5Y0Y9Ho2brh22mCZ78lJ+gJhsUDdYdE+iLCU7ecL08dohEnnSLv/kDZQrDsy
0JERIWJlL+vY1MMSpHgHSbSchnhnrCQ3JktfLgS1n51uYU6evAajPD6Ck2Sz
HNkchsmNAUz0a0TYtpsGy+WClMLJMEsD2hbSW07btcRmBrx4xcVqKlAoMrQ2
23iN7FI67+LJgy4B00hn1FyevyBcnKo/GLqfUnfUTMhL6cq43P//RiVKOIOF
PTQOZteaIu1bR2csZf22SlTajGQ320AAYUUN6lzMFrqK/lvWjlFOpXHFyi40
ViSUfgy7ausUIC+vKlcO6YhUO6XPYxA6pLRLPn55asCK7UpU0G6u8TgJNyP3
JoB1L1wjau31fEny8rJiVhpyA4zVqz7O8ZC8zRiddsvYkGsE2y1SmjJe13Th
/KonMCPlLsK8C3S8nuho1+UV4Bn9ZG+P7dZGnmU5haFfhjkQEn42TRoMvNR7
lEgjolUcth2TV1VDQk3gLpTm8a6+B/Q5Czm7VuTLK9btMY11efgLvEL0NJdw
CfHrBfpGW7yF9J0YvpMsPIqCMC83L/yeJPN6wCQGdDwihmweNiYPJrZ2WfAh
Ngr3PhClzrranPXA6gADAR88aAPXYlXYyZ0bhQC2yrhT6TJBpsnUI1yCWLhJ
VwEyO/waRa2CmdlYsne9I0fOSvTIK58kQsjMc6eaZkUJrVLFCx4ozw54+/hy
qdojhoZ//2w69hmLjVWGFos9HEOMLXbNGm9bwxmxLI1lbyyxPj3q0WmlG26Z
IZw88U+RCiLQrLfRG0GdL5bldpLtcOz3eyOkAPwLqWAXyINi1T3wjMwnm1HS
Z3FgRiE/Nq6EIdJzOcF0qMpFJniyaNa0XePrABO784e2AR5vfOZvKMJo26tZ
Qpfd3JFDZZtJfNFHVtVZIDW26JXJHjtRQx53C5STd52MB7dXVJjKT8eOXdU9
kS4wHVQCMvuneeHrF9eIkSSzmh6ke34BAeGxoTLAtC/C4rsYEN3yJOWxawbE
N/T+HgTHfkJ4x7KKjSaqyRdzwrI0cC9dDSqUPsu33FVMN5gADilmnBK3rigq
pGb0JssLxKDnldos4PU453OUmQRJEaacNfVNXnKFY8kFHZGGMKwdqtbIuJbO
z0/EM65h3cLLqxcQp0Y1sG7bMTk1DdrOq25qhj6whVJN8a7sA38pUefgruA4
hYvd609OjgZ4rYI34AiAFXLmlxGugPGuYrU/Yzk+t4UDbZpl/Fv7wcxnlEpH
ubpWtFGMd4xBzRAf06fCdnkOIae8ksuaZJ48FqijhZwpXC3GJ/bzYcmzCygt
7r0BUOGczC1FjA3vKzp/UO26W0GMF0aa0YdKBDuZPFDwcFUklu17kYBd8fPc
s3Q8p30xt8lxxtcMzyH8g3DP33CV0CgTXMuVb+pi+gaZ/+ZF0Y7v1zvclzic
1sTS7edANElQ3OBVyPJAVBHKqq+MkK7XfdmoZN4jnIroVwwW5aVWAavc3CU4
evXw4RSJwfHDJ5BqpAW1vpibWeIyVbPulLUfW+uwVaADhFbBiQKcHjXfMcMe
6UzEjsGoILivpWLY/ob4cfpSFDcmCbNghLOg/X2iW6tHB1rj4u8twRqgvwv1
LiFqIvbVESGpx54X4JNTTIDkCa/JnT5yBVgqQTXZ/Q4glZ4oC5VfL+Nyaq4j
7xF1F5ajFfw2smOPtsXeibSJ2jVZD1rLaEmFVC/eD7uIp0u+uqXfv09/Ak6Y
odxQLWYosw5P5m/jT0IJDrP7wSK6Q7pALIm6EXtwTMsxmiLXNLsxeew6hkAz
mfKc4qLQFc1TZrPZSk2+qOx1D7g/t/+Tp7sSRBxSyXp2ZoPj5QBvz8t70rzk
6oBNd37HHojDDSQgWWtvBTVN62/0cRhW05jWTbCINX1jCARPfGMvnfLZebon
2TQqEfBI90bBlzdFECFL2aTXJGfNeLS7pvIkrEzxb+3l6mE1Ys2DrVAdAGPj
NCtwsA7FgLxo/y74BKNNppYTjrkcEpfT1j8Xp0rFQxiROHrqNpdkWDcvJdv8
x4yGASdSycdCQ1Ur3xVAe7Vu1C0V6nOEDluovDBuHbI1ppVx/3vhOaVUfaOn
fmpHICe6yfHH75qap3M/F50qoaaM6zISPJdXOZH6Bx5Ocldc35aqOR92UZL6
aw69gTlmKxGQz/+1rQkxAPpjv0xZTSwjbav67TrrmnIpyuIfcqMAQmiyQL/U
/TJwZZSzWTcJEhyXDGUSG97Yy5GuHfTO+WaSvBHuFLnbiO0aQ/e81/R3P+7/
mSeuI2MHD/ymZk05r+o52oTAuFG/GPZ5dMviqKDHIsRUd4edSOCHzW22Ibns
48fos8IqvnGBxoyaAiM91rSL/SAXdQLXIi9glBjtvkB+oqCEnLy3op6cUgOv
D7e0WJ2ESsd+VtQShMgnJn9kWtWOdCGOPVSIJW2EDVAqcaRXASu+AQR069fg
2mILLpCMEy9SAuJ9kISB9mEJ524CuHKKlmqD5FNd9Rm96cLGGI3g9mCuT1NM
YQwvIfouo3bp1zbYdAMu6507Wmhbj03+rWIE435VGCQcDMhgpFzSJmtBgsem
XBfGbY5EU8nFPXUh8SsKsjALIly7rCzC+6kTyfQsG03CwF8p93o9yfbkDP0a
Du/OIsfzGK+KDNRaR8KHJ8ldFI84W4MBuozj4nAZXa/xgX9zyZYBH0X0rUXi
owTNLK5kPuydrRnH2XLIc78C5aSaheQs2yU1RfLkPFUV/QoygBk5Rhe00BBI
fzaNzx3wNxjrhkS8zJEa5KT7SVvcQz+wjCrKvqMSdxmV2IifN1mfz17E/1w4
7T0NYvCOFk/nih5QW3isd79HeQA4RcrZ4X6kd+05xaDjoaf3iH8gWDjWUOGo
g0bp8DulYNSdFJHDnVIkapsAJfwUOlmxGv+yTlvsk95FlZvsMCIsEe0P5qOQ
Gbc0Na/7zOUsQq3fBFcRj28mtIUYa3b4EUIuLjlMms2zrHdpMv5gTCJ4+m4u
A32WGm3Bwe0rMIbXMGFXltygtbzTYf6N9vNHNgNhJFSdSApZ02lbQ2hkKiUE
NapcxrtPIzxOn6c5i/m0xCXyYycAcIwcxk7/B7R/w3s9lY+Betf9+adr1B+4
24VSUo/jvFoASJsihR4Er8HPE1+JuViT5qZ+iwfHXOfx0H9sPiU/6XEITn8u
QxyDBw7FYJ4KIJlGIuckQOtmsq7ST1RCPamparSCqDPXAvpWq3Y=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyJI6h9/Q5Sj8DBKTnqZu1PjU+hig6/zcixmNin3xfQfpQ6hHvfvN3FDqFyLEiT8EWW9ldtyFe5rHLvIDM5ffHdwtQuHkjCwGOi3qnzUuv57dSG1/MqplMbofMC3CPmwIJc+9PoVWtpcrILhPXZVCWK1WxNgYfaOuc02+edDwg0J2hLxtA1oIAZ4YxiPKV3bXaUMF+VAlV7A3AXmDWVIfhXbRv7D8tBBeKZ1U/wwBjkbxnoRivHjAD427KYi4ZXQ59z3a1AME/fH689w1hsQiE+72Uhn8pV+hFu12oiueb+UBHH6NJOUmrOFR/u5qlVbkPF8dOxsfVjHWce7bZ9m0teaM1N7toV5+sv9xrHnRhVuOKOHpEuKEuWSdjnJLE0hS9Ecjbk8f6oFwxd+qO9JWFN3yorbfePPvo9yF3JaDVPI8xWVuEk3JryAfqZq2aN0Ce2A2FBFJwRzqtfySf9JI8vNnmsUyq+QI1SQHjxE7Ee867NzbRHYEUpW7hL59iSd8ai+XBS6AgnNn9ri3N743ev/nRccCA15KbC18FILvRpa0Afz9nDRr/2otOvrSaMIa6gwJqPWpUkRrekZtQ5/adqXunZWJvWaW0An3lg66TYcghE3adQt2+ui8kjrh1QaTGbveKGvlCGedBC4K616Twc6kLZhX2uRpHisGXI9qlNWiNfRByRxKKb+XhqzDnVZE9pIpV918QZ5hODsqBMj+Y6/dk9IzReI2S1Xgw/mIjrKlXH0NeulsDo3a0C05fp4g3rJCVozxQYwp93sRwH+uWsg"
`endif