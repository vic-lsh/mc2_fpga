// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
a3pryPCaJCAyqcWhexdnvabcrNkAvuDP/6l7L7uhaAh06VlPHiDMory30FiL
KR1icCcQ7XZ3hLox7+WpVdaCWy6a6HanQMwiqs6n+UJlvfqSG4QWVHmTDQ5S
W2Uiajop2lpO0wLD52o4rhAHEE42ADJgqYK0b0u35vimAmjlNU8kWemzFXlR
Sg71bEJcK/NfRXJNIe0kInA1X13EEgreb5Rk3S/hY2rQ74Aw3+d3jvyvvczA
pLv5K5UbvYG8+Of63eT7kJmnH0spTOJiT802ZdllM0xxun8WDkV9lW6xMDur
bDCvqFiDmNilUA0ZKCYvtpzfyXEgp5yTSFZGExWJ7A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jYPVH2EQ5b4b2oOzhYSBbtGkLyNVOVd3XGDjsd2xJ/ynuTaWXQHNJh1odCcb
mKHSuCPXJ8B2fLDiQwrfm00a6Vz5Dc9yIzdQOGfweMm5jcDmVVgq6R/dmlKF
/sMUYd+Hn4lphTAu+34kB7bJDwybEtoUygtBwvmteJxVE9xRfFo3VHNOLBwc
1vJS+6wK1qMbSwcj4opfI1dQZFaDVH44ZqTZb6ygOwH3fPXT7NwRX3qsJ7Gf
mMtcAHi21Rv1C0KruU0von7GIg+Sww3n/bVLG7kzNmw+Ilu4PnHOphZxwe07
Box75rGUSwmFcd6ZC7nOT6n1cZ6z2RRj67lpRTIoUQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dBZs6Qo4eLzSBXLWQG/sL8YQiODQWFHb6Bb0bohFTFXW1KQnRoQzbJiPKO60
A3pGAkh+iGw79MY+HsQbKY/DtAGTPmU505lxARfVPiUa/I0f+dE3jc2gW0lG
dHtDozSaOnoW+UKFQ0wBdf5+CdKB2pSnqv2HL5pn4PKRkhsRf8sHfutp8ihK
8T1ZTy8LvfU6HVQ2aOputVxoMqtqO53Up5Ga4t/LosZBWv3qVDjRalJEtxNX
ix9VGruy5seV8mPY69Er51ffrS5pD9patcbAthu+4j2I1oGrGEeVBLnc2yyi
+KbOB29wUz5Tx7POybqKjCIIEvLgWKhYCXNNbAcjVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BdWSTypUmRXsObKROfAh2QYVCauFcKmAfDEqqENQWWdqucwBpi8kFMmnE03v
Xw9Q8Z+W5IpQZKt3QFVscyvq36s4/C0Mry9ALB+Zj4x2tdKGocc5Gg0dwOB6
wICwR/N73wO1+/Tas3JVsqGCi0fjvdVpv9RIggpQmjvGIQj8n4/2d2FZAWdv
qIySlJ53bhj4U1z3kWY7PWsrT6IugGqdBz66dC5Yn9AH2QC54Y8CtG7+XHFH
kH7K7GJecL5nK0avzBiDvs2BDFwwSjK/tDHbEYRkfDk+e2hdAXm1/H1utXVe
5W79aTdtyvLbgiqns+6VbPtG8kxACxda7C08YGIlSw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rSBDZmhCPAcCSTtH6Ve2jYVUp7KMD6jRn9ydQahdyA70W7VRRM98rAcMBRNO
NLbFRwtSVu9i5YiRQ5KO1yK2hd8rw7rvULe1SAFKHafD7fgD6OSUN0+qtfwS
Fi3L7X8a9nzZ4YdbYglu3u7D9DfkEQ1AldWn3X3NKmhmmI78xl0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OacHau74w6soQh98k/NceX5Oi7rGcU4aCvHGbFpxR74svbzLGsr/JIKG9W4r
IA0WD7XQ75GRc8emo8DuhGJSOi0nKFvuAVEvyh43ZqjUQ3angnnvfQfHLi3q
joc/atk9EmoSjUgBPxyU8aFguW9g/5HdyM126rTQicQJ2VnMFqi0EDRP54Yy
laJG0EN00Vb5HuQkIrPtOf8Vf/6M4xW5PRF15Ojurv65uNgjx+dCdGzot5IS
vvfNzSdzer82JwVigv1+Ceg/GyNLeLy3lefrUzUwGd1ywr20endKSngFhacq
Lg2chdD2ZABFRtI7/apUCpqhIJs+ULrsFnHQwi0LGppD5n5jrd3l5gKPv3Rb
ahVMwdtaZtUY34rAn8abHlQ7EDQG1ADdTGPbPN2YICES91TBrxaBVzu9stOC
85yIQ9i/I2hMkX7RLUsSyIbORHzt7LYOl3eq4kZVscZxBVPZCtQaAPHjPJ4O
5QsyX+igFZ19/nvrtYW6ScQsEnedRw3k


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KzderEs2dstksPhIBSwTPEBXvejEPTgha5YTlnNT58hiS4/SRaXS5kD6sgOh
qbi9JQGRiFioVhPbIQupySX69krVgG2XVNaFIYoRQnmkSz9XTiFTBLug/SEv
8Uy54kfAf3jcbN53xOapMdzlY0PMjzsq27oDGJFT4742kqwOmZo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mz/4jWl5TuTHH/4naojpKrL34EbTt48ns6vwMZ6ObpOtD5Nk+kW5MjOY4xsa
IVqky35NSCjBS8iis8GiqenTXiTNrJHLmyfXsCfy55OZosK0YEvkTTnI8nJC
rOZmU7hHTWZmw69u6Clbfx7zT2AKYEcr0318JB86abKGQ+34618=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8960)
`pragma protect data_block
yugw2IhbkrrPjHj6oZizSgLZvRdX+HF+TmzDkmwF8i19S3eT6dn3Nvbox9bo
K9ZA6yr9beWQlwPxC5aZH/XjRaWfN6ipZqODbvyxKJjr68scqvMoiBWNPCOG
P2Ko/Fuovb93QVhaWUlitODOk0vkCmUeT1yrWrQLdmVbo4yTj4rN2FWB5Z1Y
VSDHgUaqTzcgJ7IO+v5V1gWfc1R/7dAcBzLJQGrt9DQ+G/c0F6dRwjvAwLDA
Pr9BBaDJspZDSeiYQNBLLpkS00mBlOj4GLcDgqno0qFusBIl4m000vKG0NOW
M9ICn5POgupXuGEn9yAgG9aR3qP+GwgZVDLJdi19jr3TnOOuj8t2o7rsEzWe
arcRGmrUh+D3vLkMTgg9vR6cb5QZmywGoMXOrknYmxM/ghGJiOIbrlEqZ0oN
1soe8hK+OsM3lEPZCLn49MkXoY3OrnY7HAXfkZZzBqVS1qt41sx7N4J6s/Md
z0ldWCuGbcmmWDLYsjL+JafFBgJF4wPohg5bIWonhGwT8sYg6TYi72ESGbM5
rGwilEZIdRiAKQiLkvwfR3VKACv6+knFi8fk0chufb6fCbAP+36mK9QI9VDT
M6JNhby8GS9qubc0R7rdv08OINbuzmzom2VCBPzs2CDRjEjGmM0F1dd9/D8i
q9Y3zN12SmEZ0NK4Mpw29PD2ZCY1oHjT3BfL+djlqpIwuovJJgyw5kYu3L9N
b5L7fJ53POSec+r68k5iK0oOf0n3isuxIly/ZjQlFViyIqubPIcWbio0pwlN
GZ/GthSIOzTC+sNTPps9nOyCtj7rC9RHk+jCcHi9tT7vHVSXQgkOAq4Erui2
iGqzDh1EGURRO1/JM1RPrHsmBrvbcXD24VBubmTiyqhax1TnfZCIX8w+E0bP
u7EqFrXPdRCymT914aGUwGgYNxvxCxmFduV45uBuuLmhY0p36OH9Ies5sLLc
aZvQru2CpgU6dmYs18NUwNUkF+ADTu9mCPy8tG5KXsMzazIFs6WKydojLGYa
dEa0gn9MkLo+Gn0rco1OHgBV1XP50p2dAWK3iRjtjWJzH3rlrHuk3VU0vLQl
VuhKWJZY+GiFD/dSiAXIrhCng1iFH18TfRUOBqWkqCHabzUtL1T2rhKgr33A
/HnPi5260jXXXBlCNGvB2Xjfx6PXOjvVN5eFN7x3R2xYL98DaK7351s34c7a
XYztrD4mImo6A+KygAeMoQa1qYJHoTrYjpNLB6tsir6gUfUlBSOkr3NqHA8d
pKEXni7ywOzMJPJzdV7rZgz/gbWbHcPdjryAgWGM7gY7ySstISqKOpwpifux
lUzo/g/qC0PjZq1HN41BWdKzrT2qr2bhU5CVthLh/QDn16Vy4F7/3MlxEb6o
eOZ+NMnUy1ESfWT12qOihWqHGpLtYV62AuY66pX54NzGx2xvke9jOGbz1O/m
akRe3uolDBaR3pz7kAdzJ9S8VgftCsKISqHLIYlQSvDOv00rFD0RKA3Iowjy
WODlg4p81kUa3QXbGH+qlEmO50l8cVLJ0uxGnnwQ1WSmFoAKW0Rb6zzhLMkw
RansXibGkbj4xdMGfGck8KZEePIgw/HRIufw0MLL5f5LO8jwMMX41E7VeRFr
lnv2r4l6Rcq88ES7HvXXTSoFwyCpoXtR9UYvIoNzGQ3s7W1OxgN4YhPY1zwn
H1njoF52AUYXCwURjibGegvtGAsjnI1PFijFDGGFbEsRGw4TzRRJBwG1Pen4
VXCUfQo9C7WrrV0hKCrRci1lZ44SsvkJK2L96Mc+2b68J9B2n+MS/BuGgFD1
ZysjQm4JbLWV4R3GGrY5wtlLNrEFaovmSEdtV12OaS1pzQz6zPH1QzNkXazb
IepATtx8MDffEbD0VMhdakUXbhu7RLlCMoOjJbVv3l8u6IMn3ha8iwgamSAz
ZJ7af6CXCfD0UWaxkRxs6+CpTx9CA/li71AHjvZkGDad7KzuoIQb+DxmDC+n
Obq2EDD/FwelGcjGwNBRyzSLjZebcJo5bfsxsuLYcTp1nMmEgtqlghYq9pb7
bWJJalW/Tf2Jy/oTdGouLiuYOMAtmwfIjqeGedxHnNl4p/9S6vkGlRVZTBgf
LOpfmdx0tkE6jIXMSzL9JYkK3Y4dIRVpFjbZIdWXBoRQNmRRGhgZ6I18WCRw
D4Nbvz6fuIzbAS9Y0kAuIWSKB+UPo6jGpp6/duBcUVEteLoRuvQHY0Xp2fav
RqETH3ThK8gcv1WPwz2LbMMto1zfJ4ULazRNgvfv0O7IQ+vEOL6VY2UGxN+h
uv8ae6MHSpIfC6GPE5XqM4WQRKe4QTNJYgCy3UxmksxA72H/QzY1sd9kCbxZ
+JHekpXZ+504Y3+pvq5omEFWtyTxxJRHuLk0fQiLPH58WCmpelmfDWyJk0Mx
Z1tg3OFjgUY+NuB0DP4H84GLvfg/109qiZkAcSB9u591kNMQ0nWMInxbnw5R
h77W58Sd7avtGjCD3xFF5oOv1dx4qDww0Cy1fWke/QxaAXmOPMYn2q2hCrjb
4ebZfXNniMkmOFAJ2Zx0HT1jd7YqRH7whRakdYNWiWPLr/TbCT0q8bKYV3XQ
xhmAIhvyDLM/Jya8vJ2vRfO/2OOq34LMgu0FlT2dJXGjcl48qoDzItckURjS
7fQo3iyIocyPybVmvChzbqLJg0dErBrJQHzfynCWsQqo+AO1P9hWtqbyeHHo
v894Ojjvmi6Qf4v+Bt8VOpY+a9DzsxKOAr6nm9OH1gdN3NtiYQ1yERFYLiVz
FGP9Z/tVL2nqN20dXWK25U+HtqYjqw5Q+DVPV9hcEaEYzGqY6yWPDiwTepsI
h7JnZ78b6XLPXh4/AECky5aYgHvI034t82q/ySaLwT0VKAXINsgk1SquWZ55
K3K0k3vUGDNF1sS9EUNejttwLrVO5aX/bRwt+IV3uTjVeTQV0N09Ux1ThKSQ
gIw3G6VQBNnJR0xH6XkGcpaZJBRobe038sWBcr+YxOsS1Qxjdp+TqYyGuQMp
xzDIxys5Q3dBVeqHHnCOn3gkITyJVAGsJmV7+BaVatGhy6JdpVn9HZsuaQ88
Tovrmw3U79OfWw0Hq6cRlxlsJfi9MrHk+0W91BZYkNbWjs+1TPx8mSP6ZzVD
TtQnQzISVRWtnECfA0lVBGcnMhi2L9PPZeM9VmNCLeKxs1DiUqcfZJWIplYR
duZI0pM/dWVOCAO8pxbponD0rJGnXnBGaDbOqYEx7OB1YebXHlIuNaijpGOT
jgrP2pxcsHSfxJgnmmGCpE9K3JKrlKVjLBtR2QMhMWRPNgpeZoxpUk2TjTAo
R1OwNrvvIPCmhcxT3X+hEI/tei/d3rXXIDwYQYvxt32V6tjCe4DKr9zZxfIN
UiD9etxVMNFXNx755wYnk/pvOGlG1XlWIrAb9fvJAl+T7PcwYFOfxqffWLBm
4A9VQ6xaGKX1nl5pX40wE+4gntkiuAodYeRYO+AZAUaEtCM2QoLw7EGxAF6z
Va3ugTU7tTRmQjlE6ZUeyl0hN9W5mb8q/I3gyBBKv88V5DmpBZAOAJniJbJV
Hr68TZwOWt3H0sljumChnPZR9rdZVd+7Goe/hU45z99M4dSVIG2sSy9cM6Tb
dP1FWGul9ZHH2TD1wS+u3C8/9umXtKMmzc/vHEcr2LTOti5LVvSjWyRNkAF1
ulk0BsWi1FslOqSuVqpDmiAKf53DR1oyymVDMu2+4Ly5WhgiTmd8nLIRIdrI
C/G2r258Mo9VbtvmA9mqLpyvw02bssUuBsPnddWt+KZX6rf1JHMLbrdnDw4V
+y2sHacEwLJAiacPuiRgu1mJnS+SlFoTELmuNyELKSGfNNWNS/3WeOgYoT9t
Q0q56hHUANpFMapVpT5FzDZi8ut60ESKz44ORHXgngdRC1K19WdVrVSffk3O
8rfi/Q9YWXqbrEtZTJekxOdTiJTBGqywDhR7xVOD1oeaZypuFd4jxiEAGolM
0Z7j3iFtkkBc8hCkuk8jAvMgHUou3KiTDno0CGLCSHs+RGHv5TD1pIq2o50/
ZWgzL5agiUpqsZ/QB1QQxFJniTJ8DZug1Z2Jq53HewJeUE94hU51+BCvqJjx
XbnJRAf9f2bNWsFyz96KTCG9PUoZ618cv+bVKJ9damirA9hiHbIQMtA795NK
w4V4FSj+56suZEeKkKO/GCVT4kd0epapw5P3FqotvS+FpMZfhuXG/bgLLeAw
TtUbuDZTVFRkRgVZsAyXE+DJQYxfnM+MVexueVxJdydPnbhGi1Om2tbpBPso
qq93184x95wmnD6KityjLGJIl8kVMAlh8ESV3IbaCA4dp5lKcgvQa/t+AdeI
d2NPyxRojKS1oHNzOpja+7TOSXayhFeAtVtChSF+piETmdkxL6pQ+W1tu4Cc
HnWR70hhoDpfOyw3d66r4m9MZedyg7Ox+rJ0IRqUxdAxCRORJzrv8/WIE93X
Z5ti/sNGGyVUw5zop0WoqMiVpPVms132hmcpVzsZ0w8fP2OTrc6qXM0Lf0M7
URlvW3vPTMVKQngrU5KABKnhCXwwhLGcX7QTvGJyAv5gmaurOLDyHJnOLQOU
V2g6D2q56zK4tAgo7WmY9JXrwD3AueXj2cnsAvVtIvASVnaCThYWj6o7oczq
JMeUAAfdF8P9baNxndY5UxXv2xgTGzq/h+oZF0r7WWHiyhFv7kHrZZNKq1Qq
KgmWTs/qD3W9NmxMzlLautwXKdgyzRwYg27MGituexK94Cpy++HmdT3zZS0v
wC1Ybe1pzrEzJ1Z4KVl72MP8mj55/ITSAmtBhB2RL+mszayoEZjRfTjPhC3r
m46WQmCG2MXe2vZh13VppHFjws6OYvuMMYor2NcmsIaOhF8zyQrqhPD5zz7c
hmIq6jEpUI6tTzuX0jFSz/DUXeFYrbul9sqlF1XkQyynI5dMQjV6I1bBroQ0
SN228GYIrJXnepE7UHIz4dEgBOGLjswjUusm/XfB5KlqPHZuixKw0wUcNUN9
Kq9k7E8a0s0gbr5U2g0CVGL8YG2+jzHcKiI/8ouZlEH605+p/4t6Zk4ArOoB
PWgj0L9Papi9HzonFxoZzuuW/BgB8TmEusOpZJclBKimhBwcwczLNqN62Am5
wkboP98A4otEN7RDboRgOVmW2Y78xclOHMdSQ/GJUuEsSVoHLeuyNWrqxK98
pCcZrbq8Wph3P9TRArpoI4MdNE8x6C7yy6DPdF60GG6PSG0WTUUG7KkRFSvS
12pw6WZBLAzWQEtoCSaHNQar3bCU6+St+WNhnal9IuOFiRKEUX2pmQZ5O5A+
R6/0Ne80Ri+m7579qK9pAztOd8fjZkz98MliS5Y3avumkwahLLyolKvtabHQ
t7EuB1RTU7I8g0SUqL1RwjBm2irDYYrmGWJTti6dSJ7/wV+wl/HlqDAtvn0N
IaoRZQiDTytbRke7SwUxBm4pWPHp76c91KDe61qyri6VDdMRZQjmir+rRiJS
YU103HpBnzdSkjJShvUYLLcpk44KJ/Kv7/tX8lM8ezdqO2eDF9qB/pM57VCz
Z6QtJwSmV71W52EZKF9HTFnFEH4goUvp/GiWqyZmeEDLYKEQ3uawhiK1KcS2
PJSqbLnfoWM0JGmzlYJfyPDZm46EENqNQGzdxLDgIfhdzgiej4phMjGplqml
MsIbGM7XY7N+NhyNoJgov2/rLRF5Tue/nOhZKa9a29gQ9TYfrvI8/1s1z42N
l+lJ34c2WnFCeDcn0Zb9T4wlwJHPokIVF1Aq8bX0kIbPHVHf9YR5b3GGA1U/
3M2cd/babxL22YGeV9GnmQFg5QUM7Z/k4AWZHXjRQc+KscuWShQppbwepn2u
NFzDvUyOJyWQO40dhLp2VeR2lE1Zx2INEM+y4We1yUJ/4ngB/NqEBZgr9CmU
AYZoFVkN0IeRqJHLun8gOokVEf/CMeIOgpaj0ImjhIpF32XcossQrofzU2e1
i2B87zPJL0AZ0lE3zFyKeIo8FA0qONOUAgwIbeoTpK2kP1GpNHgW1Hbjnb6m
FcrSHXpkXV6McdoK08dlPJmhSC/qyWyyXZm24Det+vkGkwEKwyBVFdWp/A+J
9DJKQvEpZJ8L3XMGfFlN1x5+/wgIkS8/Zugb0HEhoWFHOV5+WG4wzFtka6Ra
EjiNSlbQYpdnV/7ow/ZqG/08rKy2Wg8OjYi6nj0dC5SnLDzOG0gw+zgjq4Df
vGHXsYEl48DrbA35y7WOyy7X8A+QxKNUql9wr2Guxpnq7JOAqokzCD8ggeI3
OpC+SnC9lKhq5+IOuK18ZP4YdL+VFRh1bZVi7lEjVX47pEt7Y/0KMrBdjzE4
+KpePoRBJvUlEJTXsSjASif/l4jYdzGfJRGyBfuIu8fiUgkwOjl9pTcCaMId
8hDsb19cI7PMvUXV+olaZS8zC1OjQBaS3ZkFQa56rq/asWkMyr/ExaRXzjN6
dTLH9GC3yhIlGpWk/cpCS9GIzDrIYluNXXXkcnO560TMI1NPc6uQrFWWZbW5
YWbwEY0spnGSNQY1EqJjTKXFLOXVBMO/Uz73Vsebg1MP/Fh1Qio/1wQZ/vDB
1dWt4pkG4EIrgmFEUF67WWsPX4jABXHmvurkXwvyQIIbxDqBD28+vosk8Z2t
0qT9UkQYrGxseCyPyOZ34VUuekSpKQHOx83XC+0o8M1SiR7IepkSHqe6MkX8
8/HCHsVOxiPlyUnh6HDfWYhE/K0zlyonLJ1E6UYwTlTPnrgWuzwWCW3Ybc7X
aVHU1ik7IJTqe16ZgkqRGlpoPBkaYE0+nZOTSaK+9aLNdlk1UiWxOIXNnzPS
bluRZnEY4a8K8W3oLBC/X2SWoNgpU4imQqrM4kbsOjph/6Vwedon+1U5iZMw
A5QQ5p/1gvS9gmu7vD9TP5dKyRX71JW+bPy4dXA37hH1xKrtgEtDUjqCS2J1
ptqcSt1ntHhsjtmIrL+s5lXbX9dfGGWUWWGW8U6yjsdFas8D731D5KkOc4N8
IXkDN4I/MT6zYIN2CIJo5v1vbPbKoT4N+d7QlcjStn2zCSwLFi5K5hOXiiD1
kFV20ZLgUpxV/ArWSRico/THbM1qY1VX2jIEgwrRDPFIkjMDawxFdh4/MSvN
Syb4h1NpjpWRH7+TjkQiuA/qGH0FRy7UDn38/lEwSfra2Vwaf/EkUb7q0NcC
G/rtnMZy/BPq4EdTowGXS/4/NsTXts8DvgbZ87IFNgeoaTCqKE5LQjW4lWKJ
RD9WM3RbQr1iuQFf3IyJQRAa55sry5BoUMhMIWPvlOdoaAc3KnblKZ0KhqwZ
/BvbkBo3ExCPR45jXozxhZPJ3EsI6jSbr+WrZMI3L1ojzmi+qTVtTb9VMZ70
rZ48O6CFJy2FfrHYEF6VCn/IV8HK9nOxcNra0uNdIzK36A9X1x2HUCnUB/Qw
LziDZ/62PccCUm9rv/QJvIb3fWr8rO37y4Pyy2MPaRr9gwDQxwG6rfrRiRSC
7be626hmvpxdOP2LEVjZKgK+HIkyM2W8GIMmHp0tc5rCaM+1q/CW5X2FpFcr
hvqswPpqq6Axf4HCL9CGdcTIg29FwGPatTeJdgrBgi4+BvjNtXTHZTvI68VV
hscaAdGSCwx8yQISCnTch9cumayGEJqHnxASXaQxNGs2Xs1l8dsynLR48cF+
+2I33vtASa05M3Px1Cw6QtqEQTdiArSt5SxJly/J953MuSBPdnfo4mphU2Zk
AWT+6ueJ2J0jeKAUVZvsr7cBPpd8SY9reAEKtUh8be3GKn0vMWr16582g3K7
7Ym9QDR5zOcy76hOiucsLzMngIlsQSAKfk2l7uIC+WCGJmx49J3Lk1Gq9uBL
skjRD6yFFXRdvQkvJ/Kva1vO3NXSEtyeLCtQDamNmJLLROiN9S3JWC+oMjEO
XGmnLGUGtA+4Utob9ot0BbWgljOlnFvxsQyMTEQ4vE81u1IgbPTztkcB0/TQ
5bbL8MtWdNVfErA6c1OwqyrMSpt3r/cJCG2SQxelAB09SJRzw5g7++rAWEXg
0BazhaLUofUnYtj90p4UM0AhDUJZwJMJxd3+dzp2w4NTiyv6arUwfSwVlCLy
ORRpytL7vEOUyc/tf3h1cOMlEu9YxkfR3Y3B+ux4wnIOqYG2BtQPAi70HQ3q
vPhmA1XwagYyOQAjhtRO5AkJUWfAc5khFkUJAVjTpE9h+GIXZVVMdawASBLp
SsMqFP2yhFdssVS7fN8o1v1SIV1tTtXyrfZgnqsxPKkCbUdPhDvpUXX4tuBe
2TYntnjTPLdTp0ZNWxK5uqtvQViVthPvfS8zlOA1aDv3zzhtXGA0n8RNG8ow
NckkKQ/rNcNJ/wyMgso+M618iHJOWQS0mImX48deARaeb2AhzatgeHXq0pcz
MhBR3d8yX09vARv6tq/TvqbHbmNrRML+Pv1iC8xP2sALKH/86ZeKeHLAkPHh
mG1YE+D1u6u5aJCRcFj/i+Y8R998VAnkBwHo6HXwY9/wJqJRxvrOcRDCRlKo
EAjrHiU5Hkin+ACJG/KDigVuSh8EYFkpu9Vp8old8/awoDBG21DKpHdZqdg4
KIJkt3uOlmAS75b3ih6GZnCpfUSyr16nRd6IxP71Kqvma67gDdPqvyEGwLMg
BvoCbgaUQGxTn4ulCH/V+jryx1NcogoGlBq0PEEcjtVmu7+NyJ9dhlsLqfvg
RWlx8kNTxJ+Pd+A70Uoe6WYygJLISyznqobBYGkV6ayUm3eQwTOgYcJeRSOY
vNXggfxNQi4rHli+WoNR64JIxTmbqYYaDZtD5XdlC2LhGc1xcCKDS9a2F3qy
7EQLXjWkWjtK/o808g/bruVkfgBCf6b79i90nCKFvwyoCABmmw7Xi2XqK818
5OcQjD04uvV4bI5fHieABUjDZquIGpUSg89lO2pUinEEscAaGDYSFw3XjD3n
INWa+HeldyXnH3sNUPiwHDr4uuiyGXEmo9aNiUodDt4kynieq/aH/Ov3JCFH
rBKB2ykqd9t69KlOh2cQ05t9EtYP/w+o02h0b5/qAvnUXAAvHIURCM/JzEt2
Gto6I/ks0E4VCfV8SWyhNf0OhnFyI70DSF4v6iPLqVdyqIQ0FfNefdzFbUPW
3CgdMdw0EpEic2FTa0ofgvETSSlg9lV2W/ajrqi02XyAYh9NSd2i8ay/5jqI
pdz9HyvgJztERMRLgiTpSFWY3id5CzPYK19UR41EADCJI48aa7wf/ks908gA
Ugjk25Sks5+1CcWASQ7LraUKD4Vlf/+yzR3v6sv1xcFj87JZqctD+tFHzRuu
i2hbRkT83U3jPusWhOrAMbQBHiY4CLUwCzWfB42k/9A/u10w5aFUm+D6XyyD
5h3I6jEnXEkJrtEp0QktA4mPuOEeDrB4nFAj7VJkhVvhnDHTOjxMgsJW/AnW
69VA2ycwBmGP5ignNZyhThPuacG9BVnLdxxyHsue4PVMXAEc7vL576bMI22Q
nu+DHng//bJaX9G7GXDuQaonjzuNw5ojrBu1akcGYVvdKcvdN/NYfviZ/bK3
8gCxQsqZ5PpMUFjPwJR+/3kPS1HKy/u06oDVZxICiq5jvVHd1P0NvVwmA5T8
CZo2sWV1eQ68YTxLW6rjZiKlRZnHH+br8JHbGnSg6gAJZxDVDQIix+04eKbh
0CnxFR5FSlChe34gx9JYqQ+x1HVBVwhylxMd8yVVF5HfQzjyM8UyyPgqhZk9
p1Z4m61G2s+M+m1uouhKZEvEIopyfaSS7QBuv4qFbW5+ls8iIcdsWGuto+7t
ATT3FyUP89+p7rGgzjA2TutCK4C5J32VFmArG0kvlmQXHtgB0flytl7HOWk7
w0lHVxt85G1yAPkmGbVw5Qm37zWX83HBMLn+O889qzToGut1U74JHzhJJDIO
c4WBXZdEXbydSbItCGmeq1NONBdOncIS6Th+wCCZbbpKNzUZQLuXM+xVJekg
2H7v3+PTB9QYBL7LFvksuIi0v9nPG5MuRtRTL6Hye2JpV2AJ/7kT9LqsPo82
Dv+TUk4hLvJ0UDsSmPIzkmBcvJLpWE7A8SmST6+ZC5C+DfHEf7Y2GB92HSGa
LLG0A+vy0VjKBr9KYwNIvbTgM5K39klD6VHZYKW/Kd+fOmnA426+RuylqR4m
0nJQyAJ2042iPBtFORPoFjbWN9uOJkGOyQoast+k+iMi5VsZsvdqbUZqS7XU
iRHJlZ171MsaqhBGZ1rXgygjQ3wBA6h/KBMnXtW4HBZdP3cp3G15yc5vqQ2P
zZXWB3ggR3KnzWVJ9hr8tij9xQ3Tl8asklsvhZjrrz3Q7ql/pM1uUHW8vJh9
aQWsO8NQcYf7pQ1xTjtbAsFeef1KjG07EJZtMVioZdenHrS7lTzjHzhtipSc
L9HN2S55gBAyxW4JtBDt3A+urL0nlQnlpblqKQ20B69zxnD+rSEM4m+tNrEA
fGBoRmUjdP5NrF2gyKjn6Ilbx2s0iae6mT4qLokT5mhBvXEEsxlADM065f//
QU+fAXKaxxhqTOZK5eGIoVwU6MKMPQ4wkMYtkb0ZQ+2e+fgdpo8lqjWw0aN7
Nc2lWPB5Js0sOqn197spLvEkFvvEEvJHGyOdDnVV+boTgp9Ox9FUijs2jYkL
G4o48Q3cd2VANKvnEOgQTKacCFA5SIQQa7nfwg6/nO5sAXNR4SVpY4rPSNe+
msJ3NtmmzRl7DemgObvoMsI0DAxyJogwYh9ICC2PBZy7qFQ26LytDAgy3K9G
Jo3QL3+0RVLp99RfHr+yS6vePd6lCxvQyxRvvuFg2Kzf5sz24i12QU5uR0AW
O4Ac8OG0K9vjnYpGOg4LA2sVgggxpIQ8okYLfdSLBfD1kf05Hh7FrdWk3zj7
9ufi82inYpDd3qRx4V7eMHGagcfdMxG0B2ntv1KZji9DoH5rlDXc00af7P8m
ka+eEFTcbKPD1AcxtGysb+jNjuNkBz4LytNkzWarMHJvTngDKj4Ilv9PwnUh
RxgdU7ZXF8bmUxn+9nd7+SDxeIA1zvDmGhkNpXjkYIc8Kq2YUrWSNBOVJ+73
Er1s2JOJVqqUaDM10qdiYgYveHt4e6CkvJpwvN3Ph5+4xrwbrxuC3MDYpfI4
bBbnv63FfsoST6RbZiFXrBMJUf0tlfgX/OJRPLhoOrw15YY4/PLzwUx4zMWT
floy/Yy5feS0XnFsVqSDSrmokMpzkK7V/W4Xiaj3lWOlcLB0nADApbIk6oTr
5KhnXCep0GgcHXYodlk8gcyHIJZSt8/Zc9yocBoFZzydPwJ2SBLPFGDXiMB9
e5pJqaCUFD3IS8F6R7Y3JViRlljmf8WsMG14YRsK5boUKj4om0zWRokblI1F
IPVt5pp9YPO2Big/Zw5Y+tgrxWd9/nbScXrr33t09D9yQT5hAkfpJQuxrh7n
Y5jr2Wul5kUFXjPf2wXzDPh50qs2pLMNUycAT1rEhB1zl3n7liZYYD9iTIFA
2YqjY0chqGZF0ljeoosVYLs80Xxzqvspr1iVUvvsaPnM85TNwfmjYRFXtUE6
7qk9YzO7m24/rgLh1gThimlL2j8qHs5cmOF9wfL9Nwg9gMz++qC7zf2znrfV
zHGv80M+0VbNtsl1oD9AiNIcMCdUQhLony3669qcrNUwiY5m7FpNWosz5UmU
tgelcbEqLjn2Gktz/Yqu+buCSBLJWJzxKCmUFoZhRMYk798IeXwuDRKVIV2E
F4DbIZJEuvdcnxp6XsAGUuMLlKY8AVtqbUc6UgUlzgDxrdlcBjrN0BqQ9gNp
3HKoxXtiepufljM068HhfV7RUylbZKmVV5PDEH/ihOfjevFF8ehTw64P9h43
ZTyzhj4NRGABn23Wh8YZEMeM2FYy+JtmvH5bTSVc71+vRiPK7K6FL4+dJIwO
Rqo4GNAtVj4GL+lK91p1qaewhspO3R/ZcJ/4ZBzPSFW6PeYP39pNMwa55Yof
CV5aiod82OwjJpZb86Ed1cYPyPkBSige/YwbFtUt4y+PHNBXIh09Hbl6ft8U
Ti8w57Q=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGPjJEV6UaXmUxfmABRFD29BOe/rF8D4k2EYCdvxa/MjBMYBORp/yG5VTqkXstZqaiJumadqxohR87nnhHl7EY0rJJb3gAGUdIOnbQDA/eLByWV3ukjL7/measXl70DL6sofSM8nOOiDo3QLVLFirCg424w8k6Xs5tHnp9QH6fMz+LNImKIk5vG+TcNRGBT7BDgnY5jkUU+himhN4OQxOFWI2Z7RHSSTIdD7ncD1Cg66FufPlSJgcm8u9TYNBk8UjkmsXhcfw5vq4As9I4vGdXMTa1BWFI7V0zrmD8J+JTIhOT+1rOyWPSOX+w1Q1diqqzP05ujSg+WDV0JPFl1B1CBLJ1NmZZLjYduf6pbUKvA+ch3PUjdQkQdPDj6lbXMQ9f4djU+TowTBc4dkGr7zO31HrSHDBFsv6bWOebx5HSylGLi5MBweEv6xRk6YHJSKUCsfvZS+zkeMQHM53nk3dBU3c3fHW9SoNbzpxplm18TFmGlfucbnOAM8jtoEK0JwSMhdAu7BYDv4MJ1YBsDHN6DwlOBm1rgWmGvS74UTH328E7VCVnlw5FnI7SGyCXhuJlFtYtTdEN0rATp4DigiqIp8FvQsxS9GLzkVInV0BzUz1tPhzQGkSmCUApNa2YsdPbxZSZzly8ylNwJW4CkKidJHQphMoeQwdHz98tSlD898If4/W1DVjtn+vlN1vIfk48x9Ox68Z8hhO3SysPvUrtjRKTHNBkopkgF61hzac/xmmbN8ylXZL51kjeMoGNIIogJ1MuUyoHAIXPyItbAQI/EC"
`endif