// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IIO4fXt5728zTgwQIu5i47I/PtfrF3W+xLIOfDO1lkEfv/OtvCarAa9r5023
ErZ/7Y+1dQMrA7AS1K9WeQsuOLZR+v9qJ4Ov8m8gNZ/bAXtI3nWTnRYdQ6eC
RyDW1CRJapOYwKsr/ZOcPzh7bspRA2Q2teUOszPl65wYc4I3QW/Cs29WK/l+
kLbnxK1tX5l4dWVwe71Wfp7H5emqRqULgwX2rSKjXthybh9ruD4sGtgqHGl8
xRDgy1PVlKcWw6lMIYit3qc0OQ1ER/G17m+eI+ZrpN+atbCD8AxzqaCk+LPP
EY4+rDqCwTZKRENHvAjCl8l9Xqg0JPNVDkiMrHg3+A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IU6M98Fjp8aO8rJQgYot7B2TamY49UtFAqpUEMTCm4T4gr+xSyfvBZI8iEqg
eSqn5FLGnsf11JiS7eHXW8RrcQw/S9X19frcW7/nQwYtJ35UyKdryOL1a4/F
/jVVD9EvpmyBb0lGEy2gbs6005vkLcPhsejpzgA4ZdtaphNM/V5Xcc44tF1l
DyOqwwtP8bpfXPmnpPjlCAXctiygtsst+nz2A6gdd5aSHcox1Kg5tcuEM96E
f0NX7ILuOJsMrBtf2AAcx7qh9oC+POCa2syKVFdmHk40o6kIEZUru5NyXMgZ
t0mfz/MMg5WrrOrlhD0QbU0BcMBMBelBwHtF+F+Clg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
llgyqHpQLqR8PIs/na6Q5op/lPhuXa2hznOjw6BLH60Spn6Jpb8sO3bOqSUg
wzqV5Ij8sjTOLA9s4q2GOR9mMvDgesyYEwO/XRNX83cAyq6tVWlm1oem1t6q
h7pdbPMOKwgZs2Ssz23Vk5XAov/i80Jl4ggom4zS0h+EYUf01b/CcsL206to
iPYRyMIL7FeyDTnzA4f3tGzm+FI+7d1ViSL7s8xZ5GyBkqnjBFtiQhuOy2lk
ONc7R6lKMAu4cIU5Cw/VDwOZXOFQ+1zc+L2xxZMk2e8L10mBD0UvNU6h3wNB
wWJK7mhgcDMYzx+NeH4+9zkxfOqOvNM8tMfymCTatw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qLvaCiu1o0CEKVUof5iKVDy+xOltlbR26Zwjo+aHBodTByKzIWJaRHFnXAF2
h7222QJSSkflEeagIIw+j0jS3m35HLG5UMda6YlcAqoxqZ+rCgbk3kmoMQDW
sOGvQuy0aifyps6RiaGWkUHfkkiv7tyTUCqbrOD8YXSMfqr6eRtn9AvCo/WX
dZsX8pFaTKbkUp8uS/xc3wYoOxu+cJXqbxfSr95veMSeQVJJVaOb4VkWufLQ
n3Cr0g3i6TBAuZLMEz/yJTKyzKJUyUgXHv38C3nKrZQAbUASLbamKD7HGidX
B48NNy7kE+aoC67vKbrhCMB6BsH1Ai6oSHenvsOpAA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UMRWrjvwsMudL4MuPe1FXknCeljmoSo1eErs6Focb/GSodQJrNQCTos2wmGp
/frPpuI9XWGhtX+M8Rt1ZuPRk1Pv1jvjIrsF/x9JucA50byYMmxhPV6QBoxD
GbbJ1i0drU0Haojhei5uYZflzG+0P31AXoulRSXNHT1zGPvuwUw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aN9Kw4N/hY7PuvpKHyo2wVVyGfSkpLPen99fd9BwdL/DDRYUspw5jzi+OZ7B
+I5f+dIWm1xG2DuLlPhO+R/fucHbxIF/im3NfgLN3iJKE9dhA1/EGPxWTz51
K0QEBY+Ev/WPBigGKIISfJiNC0gVuFsBR2sM9VIvxv84JMcB2l279D/aJIT/
cFGt8x11KKbD2QOv6fv3nnfp7BQ/RXhN9gD/5McD/qrDxIAvFUsddldG/GVH
tVeivpfzb8WOguNGzDltKpvmhbmHIBJkrat10ktxuxQAA/sebBO2KzDfKgdH
b1KXg4lcjBGkWrdk2M147nGghnhKLmH1c7TJ24rGPi1CVVdtJREmZ56GQNEd
sww2jbahMrLTdlsz/bIeEp1TlEfEnt54zN/sDF177i6mjeHAXHEnEwnGXZ3H
gSz/PrhyQ42cRh+5iIR8kTvPnoi4kDa2+I25Lp9gXujmM5pJIiam09UQeBaH
8MzWMZ9JF/HW3WCY8sucgb10NPVn4GFi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kUGwY6VyZzCqF9lxCahiage7ej23pYmos4qmuPX0sO3a9tK16XizC12d+PKd
K2t7mJXDV2K7xt4ohBPiTaoAncU9qOOL9Ma+k0/dPsWOXdF3kodAL1CX8UHu
dhHg8zeLbfpkoZx7WaQzr8fGzm5dGD/ZDvcwY8iyJJYm80itydo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pLOOH86+T8TLKwU1Yq37XERQvCe/elpK9DF+BluCQJs8Z75pJuC6Q3uyRYVv
P4Y6DIGrd24ZafV8s+n7ddIaDlIErEjVD07RBDvCmPhGitEOjLu8qmHBYfBH
VEdPlifMIBlc0/4JED7d2O6moC3ZpSgEBPJTm1v1EXzdj+6PKUk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28720)
`pragma protect data_block
475XHyWD+Wp6zyy82TVUA3ZFzcI+z+ZRlOZeluy5nXYWIxxPPPBAP6rpqS/y
nNv3cJCIwSVEwtj5JSdluwW3nWt53dg5CSsN+aMxw+u+vzW4/Jehnke474d2
Hp/jGOklWnnV9YT4F/GZcQSbSkJKr6tzzQEvpWscVL7hX4Esse598yJU7BWO
ZlGt7BLMXtRqYa/j05j121x4Otpxi6ygvtDfqhVBJqcztkOBgT/+O3Ecc5jb
GYGZVp1ajMmX8mbaLO7Zl15TdU93OlnFsIAh8yt6CkHwI+0nOcy24mPxtNFb
QldjeyhpSLZRIUMIXLg2nQ8YDvxy4u5wifNe9iOF7bC9G1JH1bM70zspKseY
mEeBpk63zDzVmI5YgObjOqYKL3ncQwCH6vPnjpRZ/MHdDnL1FKHDAkiDw/qp
fK9ywDIcwQ9m7Yn3qYvMeTQPtJGjAONXPXkae+VjazGWOiMKjHrXo4zSkZ8q
G2fALYQqjaNvQMKzkbTP+fdpCn9GDq+z2EvFJ7crG+A/Vwv3SBxUET1rSROH
xLsW5PxpJDIJA1aKUiluBJA/UPNOEFLnnk1RgLCqeTzAfwI7AqsUm+o1iPmM
7Vvn6qLB0Yvu2J+67OKNhm/yqQRTCCzTRj4Mxi10EgwTm58TT1Y0uTHU0dgb
V+4pilZoJy/aigpqT0QvZGdl7YIIVGVWCC/0iNLaFI57QXOIryaxmRrscVdZ
LsoPcPa8YuGT9eejROsch7UOsNYby+tNKL828FSZ52pJyJgccAkgKv886us5
/VO9eeRbfP7QDn9lPO0rCp3HJ9fPco11TTPl2IsJ874f21pij4vaDQJ8oXJd
y7OY3bW5YFSK949aoUt0opOZEDjXiOem3Z8DEb+LOSjlP7PuPd5Rb9N/Xqgs
JtwhdWzuZbokt2ksOww45yV63pBVLU1rw02OH+5CW/fi5j82ZPZ0ej744FaV
NERncUIBqadBr8MIEIHUqbG2WNjjFVAOnoIMR//GK5P1hLL8SI68VD5KSRqD
qvacRREaXGflwgaOGF1XAUTr5tcdoPi8B/lQqrMPShQbvFf8xO+ktGgF65me
Ds3QfJYsCvQwSQxa4UvTT5kb/iKF3eI7fqqnY2GV1shX6LHzuJYDPPAl4oQG
tX6knk1bJ6RfadrKpjZS7+nXeuhBYxx+ektunw+sKdu6yu13UiLjkxoaNenX
ZkH0olojUURtOkFGZff0G+7R7rj+nGLhc7QuafAil1mNq2OxMLHtl+Wna070
d2EczLz9mNBGj4hcpzP6TCmxu2UR4XORrO9+XJyEnlWKs8WLsTrdfdvXdx8T
dsGpFaqY08Xk/6FHo63sIDjSIZPSc085s4wyWCQhrudYR1sOLcCvtdF6A1WL
NcZtqhmXRVjtnyaqIQnhxm00bUx+O2ThM6cwWPfkoX1nGCxQnPUvdBGOlHDY
x3Kq7Mj636lSINkW9OhzvoNhC02ririiZXwYq+nOf86X1tNAVNDg3uIZdMU0
fZ8U1aAPlSvHb7DeW8qyw10ovaSlmEdWdMxsA0zWFMtVca/MQkilTYMj3jem
Awk942nKPur9pMXAEfaUNUU9t9LZ0huAiJZ+0BnDCEchCyWvNMYh1wdVURcQ
xFysJDBHDLOqYkF/I7wvzbS2MsjaONAi/L9Wa88/lWPBh6nKN+SnW+J+Pw3Z
xf1k9rcYoizOOCq8bhiDjGHRR5rOhNsielOp5HXwivrdRg8ug1R+ik/dnxNw
1xbh8nklvkWyB/r5uM/6VSXS2gTZJgVROHf49gtT1l8yVV3RmTLg5mSvu49m
rId+1T0fEI8LlGomJPBn27rwB/0cvH3Ty3snwo0yZekZRhOnrGLZ69N67wbR
QlROZ5k3HLlqU4PZAFEqGMrWU001tMHsq/tKHxAszVKVeNtvY91JBT3CplPc
7rFhI/ULbqjMGXjn/d1KFveLsWGpVLwM26EeuQxkcf8WampDajfJFkHEL+6B
t46N0LUubp2sDsAcWuoaxrtM0+L8og0wN12gqc6BCp2E45DJbaAxZlSglIwO
b43kT3jgFyG/bsbymE2KfiTbknKJjWUVLt/XqlEpMH8PB2FFsDCGIHun8hV1
+Kt3x/xpAc36W6rUslhbufjCUWDXKv4fihc8qzcz4RPitSqRYSQedTIOGWzS
gbK5GMyAi8YwvWC+zvDKdDb2zlBgo18Dj4lb7+/pLTGlA0lMS/42rMysvrd1
80vqI/MbxyKnAdeVNGGpQXtpzMkf+RIyatHUBaGTc8AFLsz1XaoG1iZD6szU
BFn5eG6KEHATkg3+NkrZa1TKxgNxHMKD1ilyV4yXNoQ+dmhOecgQz8KdlY2k
+a3Zv7QktKoVgqpcM0pcEF/Ohpac9rKZSMekHrhRgHjpwShWZVIHlirwA/HF
JBrnThLy+AzHB+SNNgMTRcsOAWSiJcscRjEqFcqP43+H22Gihpg5DFAWCKJb
Cxjpg69erjlo1ldjAs5j/gnWE6aZ4Wt9RdUC1uJAtRdL3t7YzqOJLvsmLRAg
EBLhyY4nvNUVGIcZhIKsDQU0Ap3moiBHhlbJxl/5iNTV55MB0kF5xcactqFS
hch3xxlq27dNFgxqADv2qehA2drber5k1VrPWcseVb+5hoN42DG31Gx/hqP5
QXVo9Vxo5ApFaonBdlWhHOu22a5xKKohHhA0h1bZLDmmT9qxjNmKQmgy2zKG
UO4M0jkl2oywXGqK+GZKSHXakiCOjzsUcyaok8FFXrsKiGZ9gmqaLzZGxiRV
7K62rE0rbKUgzy8dOqSUbFKtjsOp4LueNoDsLHZPDqV1ukyB1MUaRGJvf9hp
hphbd7QtrYtT5TbU/n3Waz5whnPiauhidzyPjJxLv5IEVVzJ840mFXa514rD
YD5UPwqNa9l+E5eq//au5WTnRScx7kE9Akr3Tkkj2vASpcbfJnxMFDHtwPz9
oukp43qR1l35kF0yvvyFZScVoLhsKoIzt5+UhtxoVnPNW8F9lkmCXvH9pOsC
Z7uMuBPt9LfaN4IQ4cCqiklyVhJbPPg9In0ludKqfd9jQdJ7coULl4BiUYbj
rjOC+jowO7MGk4AaPgaZp5HIAXXWn27E2QBN4cQ5FO+XAOe1nqM5LYotCzgJ
AFHQ5Xw2FvQVvWiFPkFIDSGrFmM5e+FanLXHi8z5wufWg18q7sxz3uJq0Yf0
zt30U2WyvM+thR3wU5uX4dYrIZU9r68rAo6l1uuSyS2qniCLum014ZP1P5e7
o7T8IKxf7UZzOhOmJqCEBFqakEeyyRPp/kRo7pbQTSk3svZfu6B9trTRd7am
JYii4OHJJYMzL8ojJ3SPgDTtCijjYTmkeS+RCV1FpWw5cQ7SUgR6pigSfWOp
QzLRi/6SywxNYPcqely2XNoPWI+dCD5XNP0vb6eNlMURTE4QbBalM08HN/eP
JEpfRHT9pfDsO5cpmS0Ddl5/PutLauVcr7DVLAEalW1DjlUQlaHU3RxUK+V1
3FjqzhXq37lv3ZhX7RyXXyuTf4JG4wM4NuS3+/v8X0gONWxW2BBhjHSGGXmy
p1NRBDsMQYnYehTFCpYIW0nzgrWRbnF/2CLSentWKkL9dMoG2qhPHZfpM10C
h6wngyTVTj8unP8f5W3Ar8WThr+23KUF5D1dw0h33FxLkieICjg3zZez46Bs
yrptIB6LF8P6x1U5SG2EyXU5VqUbyOmNfoh5w9CM+nWYI1cWKulx8I68ehSc
8ApLhE9BX8lV/IJLdZgImAnda+zpiOyE/BkS3LNAk7TzwnPYYs2kZnGus7Ss
ge8uC8ZNztNqA2og963+1qDKT7XnbYyvG2v0T+q3f4PN/D9HCC90J+7NnKUH
gKx1oyWsc9FXlvdPThUI+kaJjrvDQ1jbthFevWELXqqTK2j0uuPi6jz6RhCt
p6VeELIpYBsPDlVIqcUEjwZd6fRsZXUliJNu//tgWKEkX1GcrX+o6eMC3b7U
Wf4drpXUM13r0jB64ERpGba05e1H3O/6WGNzJG17WoQPR2c4X9kN1DBZuTwL
CJf6maulaiklqDqdYHb7c96JHrt53sPQ9Nqb29CBMASXrOTXbmUwe33C1//v
ALd5EnFqrqgT7q2neHM+qJ42NzYb4YMnZiGP5fAlbOHNR0Au/by5d/JCAXe3
4idqVpHaCpZrjm+/GgTXtd/GM5q/OOzNXoeo2KLYFqXrovOuFPB9zzFAueWG
7R9BHl6fnyq0rfymYsnX1CWsXhxRNCtlfXAKNg+G4xPc3iLNtXyFhE/YWWKN
Q8XpR/kXpi5sNftS7ZVuCkHYCpQRRXV5ngnqRMsqPG/KW1eI7ht6Cj0xO2mC
il3mNVoc+1SqSDGwo2vCjD1D0HWs3o/KCdP4FgYZpHUP8ZK84hggyKo3nrD3
mOR0LvYwmY9je3DmTg0jsjC7e3CgXGAAFXIZ6ZsCGIqpnsW7owDgqIRfJlLC
mvNTdjgTehXmt31mf40r55/LEUZQWP66xL0fld7kAhESIr4E2E1YOAMotstc
tcjhDwAbeAxKCoMShcKqCzUo2yRAOCCdQDxXpRYttRBnskgzvkLroYxHAQua
BCXjoYg4eEyVWA0vyI8YNIINkaFFGVTj7W97rrqpD76wdRbR5fJ+UQg7bj6D
mMTKvRwRxnoKhiLaaEUbHoufu5LW+gvWheTSYqBDSWCL5LDC995YPEIyc0R0
qtngEBMtXwi3nQEG5gVnmAMldbqhKfWAMlivuRl7FMAI3r7PQjrtGqphttAv
8UXJhF71S6n2ejFhbhyozqe7+a1KBoU0t5TxJpgpTIdmz/worPvojQVKVM/W
jsNRn4J5X7kCPZIlmttGuU8X9ud5cteZ6r9foK0194NU4qIZSzgbdKN8FX2M
7Vo286c7Yc8jfTDwTaYPEYyhZskFys3gS8LnKWVHoECd4AAA5fnplRsftctt
Iw+ChFfLsfuEimrfejV8YzQhXnIYGlan1YTvKDykYKK4isPvGpfwtRxHIIbw
NX4/E9QDhYRMUxeO5Yw02e+etwNJTVTDwt/PKepbjRl3mkQKMinu6gxcWB8S
Nu+uYVylp52Uub9cY0cPlQRavk18mp8nrnRD75daKGj8iDB6nwqR1IaAnLb6
NtgrV2GdXtTz0VuGttloqHpYORSpWskxHuAiCHJdS1e9dAlFDmcGPmaK282Q
zz9CdANuOBa7uFHVLdPq8fkp4tg/oZJKqhqClR6vw5XwPvXavFWgzK0+0Cv6
bvSTUO8Ec4eqc2+8NnUJSOYi8iyg4RwLoQbhRz6f8Nm8FwGqltjPRPtb/9c3
NsSYIluiFy7BXcWLgqQqevYEGiNBcdLhCvbMBwkTxr5otjLDQsXoHasKQVtD
bussd23KXu8CUM1Zzt4dH17J58r/kAvPwXdIHQIYFTuZ3xu19HqoI1x34zZD
U+3uPttct+EKduGYdMBMw+0WTdt7w7ugtMfO0Ad+e4rN+Yzu22eIYD5xU5di
Cd40Q9nR7zDFx4qJ/fBxgiGSMB8C/WllKSnevdJl29dQZkycl/gHKiRfQyeS
QYVUfRWsgexMVlnUPvh9O0IIyWrzAX92w8SC38wbptDI7Bj2L6ZM7sve6+jh
KkFvHnvoYDZ/tkJF31uOVPeKbw8+in4p0zy923pBuwafLAYCc7b6IBotrdTM
6HeHlj5PhF9B6xsZTDMH1pZX52Ma1emHEBGndKCE21dI2JsfLxwezBrJ3mPE
RGLDcawqRurxdjG/QHfzAfGdX67ESWwuLotQ1GNqe+gwDKU5sr6+5otkoffP
4swZNR84K6v08jEUce523BlVsZieiDEbOa+npCJNPM7VaapmAjN1zQwW9j/t
MogF/2e4Qvz513c3cRfLXyEWHgOQcrzAFHGCnRtoeGRkmN/LnQDIqWrspDXA
6neSRHZPoEjUuhokwjHZw1jQ+6KMawFIwsPgjaAcQiH6TDw68+b1haRiwv0k
cy/Q3WgzAChqRNb9wlNcxEdfMgP0LmOU/rRREw/jsVC282/RdhuppfWhjxtE
l4q0Aa+O/EgfOMz33hiMwlzJX9hFo6sfNIll+ISUALByx300be4WM0qrc9x2
Xj2W08tqzc7r2f/fGTuJiqfPauYgHdXf0FcP9cjr10dezvL0kJrctPSqbyGs
/hUMwgo/l3azuopTmPepU9mq2CiYgQ+no5NRUOE21IFl3E2Bw43oSCv03Tvr
h5ybVtV4KKM1z5MiwW4mU7s5nF9ueOM5U7aiVYfDXda77ynkueC5MjkjP6kO
n6M3+nl26LRFZmOnF7J2+8OAo2kPdPRkX+J9Big38eg35080gwVc8G8ZEsD8
x0MPnGDV7fWJoKrVmKQf3N3AZOtE04tuWP9RTSbFVhLICGuGHF++ciALFFJl
rxvkZtddpnEIeyPFxOBpI/tMPJB2WwZ5rH11est8AiOJMNQqlXSqfLVeYtlS
SPTVpk9jXF5uAL2sJBWt0EASMBm/JEhzwqkL8Y1XwbkWGsmodyi2CTVkbsdE
eJB3zW1SgJUxoZp5/NHQNCooR1tGQdCvnuEUoKLUEUvGAgESz+zhjfkDLvBY
0U/TEWQFOSEtPbnSBu5ivJVraZmVBFZiQXqdWrU+E0L8odlkodKI6lCNngCs
otIRuphMvIGGmPoRhLhJh8u9oWrAoaNOIjJ1PVhPnoh1Gfh9iCXi/hBEk/gB
VDVeCfzaaDTUdnmRYcQZT0oc8TUsGLreRVQtK/jTEaMvtXmIe1/ni3TfEkqt
rTKohxwL5lsWGbuhud1D47mrfS2HKcPdlq5MZKDi7uUUFzC5qvV6VufUA5Gf
xzi7YnC26fUIBvYc0SMxDm1IXBVaYpqQV9AvQXRXo3GHSKg4pkfrfaYYc5o9
DfnT7DpQ948jhBdf/GwGL8g0e0/y5tFB4nSZz5vSXxvl1UEdhN6RbY5ppRfz
GBmfF6RsYnmRPDIcU9ZjKi3fFRdrcwPXTkqeAE0lpglv+/V8JXwyJiz0iBAA
tLk2LYgPr17hVCqT8otKQdRVBfh/PqAsDZlWjYq7D1GoPvxf4mFTatLwXBUm
2yOIXCsekLCGUmkaglXkV8eoGjGWCHL4nPLyUX6g1gMf5nT6lwP9DplnVFjB
lRwyAguzvlj/PO/9fzKydjWso+/lWAPgRJAyz2GghjYg4/aR/CEPo7iBrBL7
Km4UXEBJJ3wdXmBORtWdh13ToDzsnJPMMdPbBFreyVDlS4/HJ2PD56EEeFXb
nkAdQTNUkIQju8mKWvapm+ayrQNHjoPNinjdfOMO1nlQvBo+h+Hnbr3TFn6Z
Qwbwj7XtRrWExytp7Hxxagj370UV4YJdY28xwyoka2BZuYPyzLK76zrvlwd8
u/x7a9LCntoPD/Cg7bFu7+pAj9PEeeBDImW6QThEIEao5HvDq8fnCZ1QXLzV
iy+QWssakLtV0RoMoFympkuhvboQS4L1MeZKgg5qrzrS/FiNpRAagrM1Su2S
9sWd7wdi92QqXXJFNSuwwKwByIXynuAL9wJ6AveRm2fxzyeiRKfMbKSfBUxn
cIzNMvFM751lAa2IK2FmVFuqkRcjxBc/Ep5ZXQfnSOQ2MWnXgTB4zcQKb6Mk
sCDZ5BMYRBbuAS02Yym1JtzDL72mk6Hj0bDBOFtpDCvtO8dSlzD7rBffY1WS
H8dNHHwH9v1pgTvpKbESGXqb3EBZG2uMl1J5QaVWU+ENIMkoC9/3cv+a+Nyg
4hnIbv1KLuMOks8589M2YC9PrU5Z34caKvG4tqQ9oM5XoAzmCf48aDjDC6J6
xqk1BOCae2gSpaogZlwZt82KCASV8rdutkO+0djDZwz5LiXQwJivrCQx9dt8
DL9aGwq984K0GTpB4NYOoY1IJPAWaFIXO32bUttGssgYeyj/Zm/xIXKgsgc1
ejdDmMD0EWVlHZbFRwV52nbhyve9MWSFqv0GndgRmJ9Uy+3Acu0k2IZebF9X
nIqvMwtPK6mup6jr2L7PcYkfSDb/fC++siN09zDo+FbGsSJShELFrvi6uzns
1A2aRHG7RTWVK3qnYipfEw0RhK4OEmJbPHRy49aiq4w16ynmvbm75i1Rmfcd
8uCTfzYtQmpDFw+gmP8tVi1sJ/G3fhUb4sGGLC+RA+0vDN1JCfyMbOX4mLZ4
nmL7YQeNFGJJz/xx/rFslZ4VoYISuXTw17Sr9fG4QOfOgItOKmEGKrI7dGXB
s29aaQ8cnKL1GdT7+QE4UwecaCt4mJGfHc60wTC1gSPZ9miRVh4z8TJy2JIg
AY3wCCp+h4jwCkvQJfoTWlzx9Wu7HI+puNu6oITaduY54XWx0jhlRpKcyYG0
+yS9lNIo6VWXVySY/phx3qzzvIyhnpdbixduGSIfUeEqHCgACVgAqgcBFpBm
g/QBObWuE8dAEHvfUpmDp0d6c3E7wA1CyMhkNezBxAO0ZQqe2QPNkaF/Cfzu
ltx5xXXxVk76WC7fGEpCY0bYrFBQurcH6zbDwI0pg+3GMviRCLLS1cQ/nnpI
lwtTyeSsVDFvW6I9U2wmuE2hxdU3/9uz5cpQwALwtBcsUWfwvJ1b0mjng07G
Mu/KSUjILfVNbjcSxhI2AEJ3vw6G6DxMP7pg5QmUc8hg3htzFWXilsl1MaCB
u2LUUh5+cjvxhleknHQOpQrbZBQ0wm+KVsuviz82dhUYXQu+3PlQHaC3Tv/5
eriRTtZJcHxRVQ2aTZHFzzA1MoOvdv0zZUEGlrjdvbDie3yNDqMHc2FeG1tB
5NVfqohyMiDxpBpPSJ8xBQxCqUKbMbaR25c08jzSMDa5jTWw3ppkpeOyDu01
Cck6qz3M+gaj76K7tvbM+BzwJTDYD63YaB99CQ4G8B1mSwGTP+QuKg5g70yc
N9lGsm5FaQ4dL3TBKS4GttcfSQ/u8xLBGwczQ3KoDmF0euph2HUYWFiaJXsJ
F3Mkn9ZrXw8N1IHIk2Jj9Hu8Rf5ZtS7U+koXfoiWAHkcx6DfqVXcOjhU2IbC
VQG/tS0OUULzy9+uASCSt1QBv7t4tYUgeG38Rruk/k3buoXniEjQNvMAIl/A
6EnkugTmFHm6+WPty5x8ku6PICTg46mLJDpqUxR68Ha5R288nFmwedTwD4qK
Bz2QoDiywIIs7goMx+LOYw3OLXcN+Cm1Q9qr2U8DWZRLqZlrSnHZ5QIQ9a0g
90BAEjIiNVwjQoNjYu5pPM8Q027t+F0omBwYjJlVo9YxilTFFpyklTigJpxF
hdMiR24H042pezhi2/ZR1Epk3u37IjjjSD0Zrr9goDESL0EehwCrX31+gXFw
BgBfpDoWGP7yJJp+wAQS9Rq0utkzC0TjbWeU3J2ViWbFYd4FR18NTJOJ/hh2
aSFgLwsD5BaraZBu3GQ9doQo2JF4IPTC8Rpc8lDRXNQkLrsscGJyKMX+WEB2
RV8MhqooiFFIeSaCLzfne+1RmJxngQv8oc5hRJRgOX7vfxfCO7JUxK/iB009
PN/R33CiqAe2h4h2OK1njo77w315Qr7YfGhG+oXQPEnMT5fymZJO6aKWpTHJ
3IfpfrpHJ+x3+NyPI2gyRFAKbH35SiTuQq2N7uFXMqwNER35E1KfHGJBUtM3
80DQDAYEnxOKcEG/AV/Cb8N3HBbVbW6ykZpCxDWKhvqr2TaEs9d2x3c9xF5k
YgCV86b2Ig8oEbfwxnMPlB4fV+/PXUslLVEonQID/cyOhl7rcKK85XKFFHLP
KHLeksFoOlePhhPu61Y+S9uHd+REFZeaCvgEackw7JNDEt1SRMNJyI+P2rBm
O6Ou2CSX3AYbp8x8mxOp+Jjl6qmkAZj37778pQxWa0+svX5CLTtWAE30+SCV
qcMhd3G3cHZ1On9+M5bSba3d/5G/1EG2ILHO68dsxd91XYdFNo9xlNb99+oH
K+5vZnMxRK3Y3m4J0XMDunA+uhCBPHW2kMQVSaePTypDQmFNo7qqfqmgDoFt
BkGfbB6l7ztyaf9MpUNnekp9L4d7ISbVURxwop22xivh4mNfmnN9WfnZwGQK
3dWvKVM2vzKMs0Jdw/FlvpLPVM9IJpG6kVz8C9croSaBE0aOx/kiQqIRC+Rd
lRZPOWdoDb0TTI5U8xIBs7MnCj/HDSA2fR/S/lQKjBc2DMNBD8gKBJ07j+CB
pBL2dQ7xiMW9R2zZmq0G1ubDMQFRiQEQQxP1iJYEysLEg2Qbmyass4QlDnHg
tVF9wTSNpmpclvFcWPAiaJcg3dk1E2eFZYFQtUAL2pap3bUQpVO4+ii1nXKA
t+6oU5l2vVxn7rX5wYsGbMCHx/LJhCVkRzNf770ncpE4YdXVzrg0DvHgz29l
AHIfdAxOiQBAb2tTLyF6kYnuivEluRN3eS7Z1VjQDbjM0mfl35uiwC5jbAqn
Gx4EW3fGmEJ7VMsnLJScq7K7hk9nMCi1JXc75L/oLSgkcaTgTV1mzYVnnjFt
xzOMYQNeQYIM1nD0KzhX+s7EIXNEonuHuc9Msx68LEXASm4taVzNr66gIIWy
QNB5X45SJ1ON2BWX+AVwdjGdzvPpF6bDN3Fw2mT003Kj/8m9X9El4ElEZeZd
PwVWclBjaO9hTDvZR4dn18mSCYrLckrPf75vidM21FCyHzCI5yqgVlJ4ES6x
oJ6qYiDnX/4a1p443j/krXsqN8cAnvOAwOEfAL/iiMRAVCE51raAbBxnodbi
syiC7KAhoApXv6oqxeG4hZAGYog7OnwaC1RhWjzL50zlk3ziM0wWhnPGIrq/
b5elfX5R3c4lvj1dvcXyyG9rSQJjPU/3daygzlZyrf6aqD9mESCf8zTwY16l
Y7quY11z5P6WI/fEfGh9iPclk/UQPLUr8Ev9bndtXHfnU5XZHe38m6Fv5W1P
wDEDegx/8ebCqrQTtlAZECkb9IRkuH3PhKp9o87uu4HAa8tbbMa7MMYkc+sD
83Ut7CrU4v0hToiHQvC+VBCioret3k/rdy2lsh1Dl03TCnCfhPKKSOtDcG3q
DNfzqbuy8JkSMo7K2bSZphYsGCeJJx2KegsPTFM+dTnEw7kd7/OePIJORu+y
uJcJKK39pMFS1MqG1EILB/s7B10GcfBFebmTk+4nmM0sWsBGiHRmApG3XCD2
hl5wq6iOeullViUKo9xXmqB92/rGrRkZj3eTetv+68IMUCln0RY4YgCl94UO
0cj2zjtzXYDzMjIUTkayKm6ZufIhG2gWElqbACMQxcohCpJpu/hBQf9h4j1G
yZ81y3BFgTduXEaDZWHiaNGhMkI5crGnWKJh51pQiHsZ8t0qZj3xTpGs6PKl
x6MGtjHZlNqT1f3/pkF8Hy1b5TO4JNqVlszDrNGuupoPZ/OkRBxRDTbv1IjN
qo9SNP8AaCh3OHtlorGbnHJK69/2dvUfGze6B9ghWOrGpNYRR3k6KqVkgpX3
oxp/meNp5DYFlhAE1yua0mjQbMv3WJEWVKi0QDZioZoBCV/eR1ggkZ35bWv8
qujRnTR6UjXagmBNmjDyi44tS0iIBq4+brY2Jk3Utnp8JQ1L2u8nT8N7MN4C
QfV99Cx/VhfVrDr4DFWzqXmMHC89j2LnGEKELyh8ijHTH9YuSl1JfitQ0uHb
e0jFVmlgq33DVizQFbDkdmPZIZJ6zUgydKK2sf227ybSGUNm46a5i+Xfp2Tm
tiqtLxgiQCXVJ13brVKMV6kXWvZk0p8WpnKOwJSP0XmwTK6SSExE/9u+aXAs
1FDexR3WsYVvgd+DYwcIwzO+2UoLHqOYMIfKfDj+i9JhwwfM38ia49rtknc6
xlrBToyy9DpHdyENjHCm2HWXqzIznbmE8E3GRhvYUn7LjYbSUSpr+DpMaEcf
jdDcj39pwKNWwV3E5+/oWP9IsqgCHfhfhr91HPW2fJe/0Qnmewte9jltQumX
MF2T+vAORDOU6KOz15Z+Nm/7LVV8+IldBDzzwo9pOi6vSFJbddjnbTlOdFU2
sjWAV6apQD+KAuoR6iJYDBnjVPXMgANPyDYVjrPyVTD54MZ5KJac9b7D0lND
oV3zDu1rggFP5OEseklCZW8XTzO+BBijP+2JRFRR+mHCajL43dXqY1lYnL0K
ceVj1PYO0U3LfmYs9E5R5b2bSd6Aapta+yLzU5+LpjMzrNI27R6QEApqkWJS
UAo1x/QI2bpYJ27TcpxihsOjNOsTztxsbVfYhryM5viCX3q0wbB/9Eq3N5Dn
EmuVE/b0HnePnrzUc+5wrU5r4m6kyFRX/3AluPajdVBqIVMuS0JnOfJZB4jP
6j/GOgn0x7ugMCika8DNA85Oq0ZeJLKGHK4LH2eDQz+p7Nfn5u/HTBvGes5n
F2VNk12vvr+0odPLqUOyZnlBTP5JNYHgZ+e/mXEKTbe7NxM0DWgr6gbVEMFK
LxqOqBNWxE2sAjfPmfM07BrktAJ3YSf+8ycWs023ZyDPRabndNwg+mvbhy2j
CMa9W60xtPRdVZRjZHopjX/EzTjFZW9LNyfszZufYCRu1PAKzaNXB4jAZh98
bGBZOPb5sNl6nFz9R1ffxM7OlHzs7bJHvmx490S8swsSLu9I0ZzrLwesSzcl
4InuhNsuPY/sOZbPCR5fGFdUlGypZ70VAP3ZsHDazLDFYbo86HvrFyiFoNbX
rarUbrZGoA0J1U++G+/J3Ghv6u2xfT8RlNLqZ9xBKMChnL5at3LnglEHSLDb
Fn4jOVSxleW4lBxZ09yrD3ZNWs6wK6SvKpiJdw+PGlOXaxnvryTzfMNeaMfe
Eky1zid8PL+AL5//Z1up93zJWynGJiOz+G6f9nL6YVerr6NIcDFA62Y1F1ws
5F8rKko5P6ir2bvV4I8dFCQllqBTJ0M/T0LNEq/xxDezzOZR3Z/50i2yANez
vgqAJagtmHbfeql6KxsOTZuHQMKL+3kqn7/SiGma2AWs7uBiWJhesaYVtios
DGl5oKv0ny6MKQmekgr03YKSUYMmPzTvbVHzb2d0r2p9Nad6RpRiKpdrO+/s
KdmLoar3sxiq8ueH2iDIy5DwU+4AB0m8d2rm+VqCOxXvEr9JeVNp27gCclh9
QNXsVZsmGS9Bh9Yo/eT508JRSCQ/emJt9kGshV/oMZmXh/HUHPS5Y7RMfL1m
DQBzBZgJJQuw67nQFhHa4zy1iqqfa1FseV4UEFuMEWY6Ou7P5gNd8I40UvG1
vixOYFKQ63OUp0y/2EpJps3+ECcAxNmITY2zMqnahv+h7UbiN+6knWA2dwiB
G0QEGTYR7ZzM0BUAHsp7z8qZb9LRFhHLXUA5gyYKzNQLNZsGJQRcPSXEo9kh
NyUJUlpG6ilQynxMrF+GIsXShFche4IqAxamIuVm38X/YsKSTFZgFF4encCA
0pdMX3ffa+VYoOwNw+xH7zSs/a+LvdMMG0kr84eEf21OAOCTDi3YmOS/w62t
+FhZsBIPCcHyZWspV/L6W3smcM4j3aB9kPj3vlJS4akGW+4Fo2ssRTUu0wbK
ne1GC8YZe6J23QRMyvtRul9xsaT651LenzcnsoC26DabQjrnEv/+C0aGE2jD
dGOjKQJKVV8gNDkbkh9c9+YwOtR0I7oPbzOn+TbkxC81rSfk7+584X31/pXK
oJO/aQATVQyxTbdwzsFZqYbRre0pFECmBRK2AJxum3q8N3+dj1H9ofWzEIpH
nxrt+yG75QEGFk+lF4qVGOH3gSsJP+jbSf+mQIDocSRWb98XhES2vEY5nkPZ
meFNfVk50GURDHXwwf5o+PfefM/L/+35jarzRWkbADQb/q+XsP+KsWsBBgTX
0lrXioZxnfKiexc3P2Fg1Q8pjcY+UOz8EiF9jVKsbgkhAR2ikiYYYqT5KXUt
H6fz7buiptekwU3krDh03hDNwSO/Mrqvyn0JL+TPwGosc6/U5yK6eNfW85wm
j1Z3OGZ6+KBRJ9hxbZbVtetqNWGBlOeTuaGelupk2Nje4M1zS4JvV4mOcq5z
Y/yXvxdpCanoip6uHLfQiLjIVYT4561zyq91nehV1NzyR0ovOlv0C/7MD9C+
ir1Vfk+zhU/CSvVl9sp2J9TAOq6yp5NbtrqYlKCUgzWdblEgRk20+wk9XT9s
3SfxAv/wUpZ3sYjeIZY2Bh1VADAFlfd2tgg+nr+y2jBOeykhdNEoZQWYJF6I
tI6RKjMfrk67lF/Fg7d+XrRNVbAG6jV86QzF3qx4wpt1jDq4Mv6wl3gyK+ja
rHpNNkWpAAujVBsY7vdB0VCe2yBl5z+eIsUVyeSqaAJBGupIAm0oTghEn2ID
NC6R+26z4Vx8azWVoBvetI7XqohMqlmuAGgFCYm/VVeV3i1tlxJ9zgaKLyQw
U+wdtTfqyBdqilWOnruJVQtMEPgNmBds/RnfkF9naCPA9su05EawbS8cmupD
xE2p3azm0DfBPNQNvF+zCQO4iMR8W4AhS3zulOoPXA44d51mKS8gOax7Tsvg
lTDCbBK9OYevcPjlLc5SHG2+Ic3MqwRJoyev6Wp1S2Oa2fXv7ASZIH9W2thb
s9xNX/zwa2PTlhEx4hSJK2LwwHFcpmTu6k+vA91XSfCtsMC2kHzqDB1LjEzN
XTWO4LxA9J8ouvoiGnVSVXWLn/ivWS+nLo29OG+pGW6ReJvaRSDx8RZhHQhf
uNC7sjsy0D/cr1CJ55G4NdLqYqxDacwzWGaTgeYKIgClUetBYrlojUml11qE
lt/wPseVjhpDJcRsaO45KfErvlAz31YhwWIAMWivrIZYDOW41b9mkqMjmKv9
c/qAlikCSCROG2VZ+zKNGVEsrhzlmBo5KTFqlcAHxVxiQRXdOzQqzGFxh/O4
s7dHqf/O5Px078+8Xu93bv2wjzf2K+41MgXGi3MG4eDWVeRFgY5z8CsKVrMC
JSw10OP/VzbE5OfrTJEHQ6WsU7Vzdr4PdPE1tJHb2AcGT+P7CUg1uSDZ8GVa
6SmRsByKsD2ClmkRTmDZblm28ufeZwgdo//0rBfhrsvcNzVy6HWe3tGtyIm0
/f6hjhJF9yJogoM08iiimfvFcnk5jGnjNBnXD2ZKpXwRuTcsYZFLHlWHEoaw
1SGrsPfZDDpauzFxFEC5dAGzTtkBJY2gkbRWxItCdeX/P6ZvkqdJvj3o5tOD
3PIhob2UR2LKdEI/Rs+bXwLGCwPlhjlYzO0yPYsLtJ+3l9ldn8CTO6VYGYsC
ZGGI6YMg7ArVGUlKp/nH/hDQrEu6X0ZIWmzATTYBIpc32qWV4Vx6uRsUVsKH
G7pPC4DjfSeY7bDg7+yhbH7NVQqvhFgVnJz8b3G9SuF5CA/RrV7AwV3RELel
8b37UGWlnnWR5wRzBkGkJ9/Ro+5E2Hn5vTsfjKGC0PU2Zetv17A1/fK9dmA0
YFnljJU44t2/7OECEOh6JpV5S+mg8cmLwzR8cbNJIYRd1cY3vIWLjAxhktnY
lFRRGkPl2jI3INTn6Ws5aE3IonOiTpy47WgmaXTFLndyvdzhgQOo/fPRd06r
rTcPm3T4CEXE0P7GK8yQWNjfMPeOwvd5YGIAueRE2lJ6r2iG0zU90vtPFj6c
MECAcUVMzTXXXqSIxuheZEoyu7vIblk6JxgRZoEiBcQzTlvF1zMqxzeBiKzc
3mUGRoTflOTij5Gp6jN8sykWsKpsf6a93HQzZmVSCLXwMedb/wECsf32sEst
sRcLFxOyyvCRVgh/RFBSr9irU/16v9+xgRdp8FlAetkwg/EliijbiKXNwF+a
hPW8FgMZ74Q2MbcWh5/ve+5wzseMl0cV20y/tIMnNGrScqCiwHoSeHt0s7Uk
tf+LOPeWpB48OaX0WjG1EiExtBqEqppxMh+p7gERcZl54SyDqP3D08gc33fi
HirbIeUcCt1LQd4CpDgEEMmrSS3irK/uUf1ejPZg1zF93e54H9jYO2JGKeZe
EHqroXCd4GKr4jWJEE5nxfhSH9kNHJHPg4lCCXu7U4iKXJTcMn5OODM6QuOL
Mu/KLTFKb3xMzLEqzzrLJLi3ryIoW06rXzv9CX2SXIwH0VMjIf627FtaZ77W
FVKmBusz3pYW5XnlJqrXkGkltUBD/oirjv19VZ/6S6/Q2CQngOGrhLv3VHvs
uy/WjQEzN5jpfn3gH5+5w74n3qD28NWbc4GS8YfEXb6hmNlRS6QTRtXBS/9E
FjhHut9DhXk8plTDuNAncSldcWNeNrIFSKWuvTRoss1UE2Kwx6wjB76PYXUd
KIQc/OcM5PYQzSIe63wKRmnEvsu8UXkQT8fFxs0SIFgcDmVGC/Bn/ACC1opP
gGT/5jBBYYpa72OOrSw3miq0m8WxRIuPlbAkxzanY80dWKAmwDu2TWZ4ZPdM
OdC3QsNP7XVbgS8yoamJk53P7tiLIPf4bbQgIhAcYw05JYXPW27TB3ZPzr/S
lnOwYJJ2n5wNXl1sv1wYFJkezU0r1755Y0GorvNsK3O5o4HC/UCAw5Q9nISL
jqntQPltKOOHT+HKsTC4G5EjInT5ui+LHFS8XauOlN7XqKCveR1+5JKap6j7
ULs8nWUbDQ+HYTrknl3gLQE1FRqpsdsSrjPTi5le+Vg2zi+9ax2nI7IIWNab
WBfMTwJiknGb7f8X/oticZlfFTM0L4gXpLxdLf0v8umzjWNyCjXnGN6BrI4L
+7T3carHYdIfox6A1js5YQpQr9iGeH1UUON41N7ERlloJcrPpEYER78LkLGn
RtLcUm9mHvV0+065Q0K/4tz+X6+v1SBcYsU4F+e3X0TCJVeG991QJPeRIoEE
52xdwwa2IuiyKBLzMn7EqzXIw9HR+RpDZHXSa8nv2ACm1oZtvZoRbpp9DxEX
IQYtUSMei8XbdxBGdgLR9C19ALAYy5cqAPhOu16QVN+U3CQ5XVtIb/cjDmkw
z7W+oh3NVrxPVnwY1rIveKRIUAAtKpMjhh3NjBZP9Qblwb2m9nxXZBlrmqs0
5oDmMpDcJ9+FkpN85AcIODO4/SFR9ZImhfOxvS2RxpgzW60HTGWmAdXbIgaL
4IqKtUc53qD+dU+WgMLJ22t6Y33Fuh19VQC9wlkqRVmRUa6fDtXlfcJLPv0o
9brG0sNOJh4ydL15qGMSgp1q6tYgQxvPZ/8eIm8RWYIhfyRbg1MT/lu5dZZD
9+xyA7thP+qyZWTPaGDXiego7rMBxxZYb7nPtpdGU6XL/Lwh5IF+k/5OaRkG
YB3cKavBreDxULGviHigSXBy/zkKQDKBr6ZccmsKsf1fHuDS8AIVgG/99mBE
81GbDMF929iMbu9zu6AKuA/YtFJ2u0FlN6nVLfp9P8+YdHA0k3a5VzHnJtIB
fwzz1J5EZVCpoN8PB8VSYCX+YQhSMp6syessxbAMGnjLlmLYeEYmpx2PZqDR
N9YP+yY+DSVZc2RnTommdvSA8c5bbiy/YniFz0zkthK0OhWBTZfsThGtuH4l
6DO5Wjsd8p05i6vfChcheQbEhhqvjsqurlPWb3q+RQ1R3m9Oi4xFKYq/E93Y
uHc8XYm+PUcAmoSfTXYFlh0dahZ2+n17YLA06NdndUrJXWH/lOCIaoFCtiNA
gus8QAkzQFgoUgE0/dXjo5Jfu0jvqYiKxTLqCjkaFG0eK/z7iAl57vtdYkP9
0/Bds2Bmbbt1WmDevfNu7hpwVKR436CMQE8aI7vqahsQqa947zZgdEUAb/mK
sNcNdISFN4j0jy5HqFo7aVOmfrQGzW9c4GDeFABpCARjWL2KFnu9pHg02F2G
nIthFb+fDMbKGvlyrV1O+79F8gj6A94HWmKI/O8TvUU179Utwrm2jIwq5HcF
NukP6/AFId0lku+xJlZLVsxVPr1nQ31W68HvdSNmmv+7cOLBGFilOVzzvxR7
GKrSW3uoVWjwx1pzF/cdus+b5NXEULA627LMzEjf3bp35NMB7z5IyE2FdVpF
bfNGGxXi09HfB/DtaCixFwAPhdLCrG63trQAZyTbxRRz1J5tzWXeN+S79W9i
HyjBaoMk0kub0T0aPFW2fiGX30mMnsracz0yUVhrU8jzDN7Jqqt5ZtKoaSZq
fi2LFdWTbbYsw7FE9q9XH+ehcaKtNRGQgNyC7RBU8tBIYqU8IR+caQta0n4d
jtOwSUjlTm1LnB1mGk+NqOjLY77icy1x+zGh0/skn3395V4w6QnJVkhDvt4+
i497HiEERUiMYPeDyAapCGG66tkgWJE5SnKyouewK4HXpHpx28+RlM1J19ir
3DdmpBfocd29MpPY/rSRJWGFsLpvz+aDIr95b4e9MxAybmAnFosUZRcC87cE
CANtLkGkmgDCoMfGSVZW4t7F+Y9Ax9E3AoDVTtIMlVELSRSr9GTs6aiPvap+
hmxoh69HevJLUqODsDnBElRul3VmMWJytIJfxyQH2/6eAE//Wd7HwS8BsVPA
8wQ9VGwOZahBCnR/XaErSVzht0wtnjp07HvXpxs6008MB9OhOQ1qk+Z2d/z9
Nub7sHYAs1eixHHzmkrRCgVnm3rEw0hOFnMsoBRPC+lHSSAOm+N0R/L9JcGj
FZQjl9Yqtq8PKoI7HAFtGQk15TDkv1Cvctb6bU1an2gN4Yg0MdQUZAJMYMra
rKuBINY/d4ZfWpheEqTebGB7sE9GxiyFckZJR33u+unCj6cAdf2nDmhC7Q6o
RkZDEG93/f1Hm2iJyyr/LvTpJ4zE2jo/FbcAFs/yFLGU6LL1sLTrPRK9QQpu
sJBGG0z7f1qfJ239wQ+tm9mi3GobOaYXpKbLI/MCLT7OHp8sYPVe9ON8FAyi
0B+/sS1tjzRl3wPeDZ7M2pw9Ivy4vjVNAo7u5YNo//G6tPI2jir6d80mfLWC
4LAHxg9BLUy9tZ3TI63bTiCbUy2r3H3+Tyay6bY/jGyIhFlqu4OIU1RW1Ve7
Ds+lLw03Qt60q1axYyiU90WiQAvNkgtgKycgbxvR+D5ubrEjA0OeZn553I39
ZSvtt3njxiMDh5kd+6MMt/oApAVEq6EtGox0FgiPmF15j6DiZag/BOuog7MQ
ebAuslsZknR1n0xZNdR7g2+VSzloYdez8XxaqHGCPzai5nuagzOobasKr5mv
nM0X2ppy4xvoCiRWpZnUgiYYkP5y4FTsBKG1QnIEWb9WY5Gm+FrMFeVMUHpg
9QxKp+JZ4W81xq1iZ8q9aQBRZGR2XifdZa4UZr9u+k9DJAvLzdEXhkfQILM3
nMZQeDK0EyaD5pzJrG1clCAfi7L6w7G2Zb4KFwyU70jaBzANYIPg1sG4uD/r
ghSSuXjx4kRzZjWRV0oVgbEui+lMM4CMjejZiSBcGLVg5SlOj3nbIxq2mv4l
ezmv0bFWNoPID+Hn/f6i56qJcsA2U+G/VppQFR5FmrxI9ESiXcU4p+abGHmA
xgBdhmpGEZtGZQ1hnom5a/E6b7UOkjpqH2iSamEsRxoImyC8zyFq6eKZvfwx
zKSri/pmHxKlx2Feo1S2LIh4vliZsKdwA4mcbR2bQrYIHwz8xITgfMPcJOpv
9/V07y39PCdO4Ig15bp7rgQGWuPBemCkPiwnQ7boA8fZSX/6+jFnFjENCwV4
RHw+cRvzEHpzc1lrqr4abDcdT3aWd03s3khipmaddLMafmATi9eAsxMWWMEy
hc00F5ArySJ29B9iQFMm/Y78Tx9u44nV4nWdNpNwD0Ek5YyXknPflRwlbrKd
I765ZsxBqVyhL003Sj7ORST7jRByLr+3MxOqWnekdE2Wxpnd9Fto8ZtYfoCn
IoVpZFw1Z5KKola/G+kVD9NERtsb9z9VI/YR1a+jJj5x7F12uFOLkwoU2cFK
sTTBmbjME9VFvhe9CRFqlEKl06mzwW2f+8A0padZxDuBrj9KkEpHxKBVw/wr
k1yi9lZ3ADJs3yMpWNTOp6FPAuWhlBfAxa9EkzJ0RNTMVQesGABxhQ9Y/9xO
YnymNPjW1JK/SuHB4Jxuv7mORlfKrilvbrcIoBzyKoGIik4rJeqFESHHp8gz
ofy2HxILF4cHKhv4Xij/dRj8I3lFQZ3CW/AGbs/BzERmj/HExX09hIi537LR
Yp0HZEeHlonTHuHOvG57mHw2lQSKTrBRKB34w7rv1s7pzigcvtf4VDwpeZSo
FeLq3O5DijmU+w4HmlSPbETWRtMPHkQdUqgYbGvxNT0Hy18d1jwK+Ac7tPRd
NZeTmTUJV5x25a44X1tBkKBs+WHDbmM8qzdQimsn7e247ePe/72tnkJvK2rI
dRrhKHDCw0eO9WWZp89W0vlPQgzOsoFvKnAdRpG12H2Xlqoa6chDspFCgMnv
+tUp65Cyb1Z90XX+/FaNgUw82cTlFK6PB1C1NPI7JqrRg9t+cWGGLofUaXnv
nPuk8CWySN2eVUR4ZGRO5zVU89Ph0CJjY9Qsym/EBNe0VZxI48BwUdscbbZc
wCikAsPPB2JeepE78men7TVSIV2l0p+kNB2hf5Kr7GQ15J9HYmfD/LF3TbHp
RUzMU+qeMhZXUFP8xVNwDTiwRxR+x2Ys2EfvgOA0N+BQ9wbYTLn+QQ4vn6Nc
6G3N6VhHv/05/E/nHIqXtG8P55AXAUuOCGJr57yc513ZRKO/Z2RjU63Zk6G2
tIZPGYAc+bnonapVgRr5rBH/isZZlE3Vc2oJncKu3tTvlut2CqRr1DtaRw8w
Q3BJ6QgDWfEdLH/0ZxDXCXx+fILkTILV+hW49IUo7cPUpxu6w7O2B490kmkF
SIeMD9k2tfL/NQJM5RqOcYLseGx29HyKcLJwPBHxxHZH8Up71enCh0sep+di
54jMkuuJ1PnnBWxGe0XZwC1u/wPgUFwQbKTpsNsqL3gueyQleJMe8EzgBIrG
Vy1G2d7DG31odZoPMc3VRBGewkIAj+h03EuJVKKUmfYayNzoHOmLQz3gJ2VN
OzAN2Df/QRhKoxby4TJYmI1qDKKWM5rRHLWtSWfLbYMtE1QVf6BIma0S5fVw
hICBE6LNoz5nfFEKOvyqaL1ohlbPJ2CXXfeKjmo1pJUJ6N22jTPBCIwY/1VL
09r5y9ZB1p/VhtxcKcrNcFZZruSlSUUSXOk0oReWuITWLkl8VaKtIBMLNw1B
NI6mmZaxUutMWTXoEU6LPvXh/ZML0wgcU36PINoTsrfoIWafCliPY1BCXXh+
AJ6wANPygMXM8haIzsUOwu97H4h1dHRMiEP43LrRHw7kdiYn8S3wrEdH54iI
ksiiHHoH+q1N/1q/YaJuEi7lJq9iUNHybhNtoXbgjGHBRchrk1oHwp7Xs7IC
1Wx11A/PZLspa1GDnQCDOPtqLDfqNqDZqsmtyaeaDAm6p+JYVn+6O1jxZnwo
Y/qPii6Sxy02Ndi09vbXd096OpHoC/GnuKwrJWR7lFyzhGNISlm7Rdd8UcCh
LQcPo86paxcwmagp5syZ0fLG849zlPPy20ia1HfH0gtF0/qNzCmGUaNX1/ql
9hJGPiYFg5NLEQkqT2jP1/fJTp61mafPyi+/W4f7jZFUvVxxhLkOqdcJjDyP
w34Bmpe6Y4jJB97ybMwEW6V8uyDhJcBVbR4luTQQKEoLQqrpxTMofFP7azLp
mssnoX5hCcavT5Vb28xnJxpGpamAyg3eFHrRHB0al8dQi+4y2xCHxBP3+Mcd
b5O/bvAzxm7G2boZvAaX3bykWo72Uy1K13pcIQ4deEROEoxK0l5SXH6sU08x
HROgmTwAsk8x6yjpKpn4k331u4PDdV19YkSeaCnK+P/Q2UUDzCN7uvopOrds
6JIoBbuS9+9B7AMW6ElV872EaMpnxd2QSmmpgVRBTZbyRo9ozHvQ/0eMD/Gc
dI1KnUhdcCFgBBX1gCXLFDnucoZ/H/tcRMCcvg3pKSY9Mr+ucLaA988j6m1e
QQd5ygZ00HNmglVqtV36L8hz9R+x1qKAEOfHxCiXdW8/5Je2FayuQhzZNSwc
k88CUrwO4WMctg78NuMO5/3KQAuXj287ky0ygsElT2r4pbNlpYFbs5GwsucD
Y5C8WXh2dAneeokoryh1TSWo2pkQytKIYFQUGBwqs/iXCagNdba7Zfu+p5bx
GxjvTFsrdZ6cCv/S391wjqEmDfj6zBkt+6wldAlQDt5+9D67kHGwXBEZXd5z
KNhO0EI4tlJm/Zd7u9Rhh+QNqBnoyR62uKbkRO9zq3phChJwOy8E7QDiQrFW
FQcqnysPex6y5oruFvt6YIO+KVy+mTctuxkeTQe4E1gxbdTXn7HlDdOYaY5A
qhPXQOTN0RrGMMfZp89VhkaM6aYGPFBZT2gaYOkRG6zOpomH1O/AJNLuLDjb
QIiES5/vqrL/GjWAXxy4FelRuAnsn04r1wQFiKe/MoTdtxht+8rpajHC4Y4G
py7mmuNnoqJlR3nvjUDdqIUNLmQE9ZfX1v+11T3Kr0IFNYv4Dk/8QnRN5GFi
QHyo7dbHyJadd3ciYom1lsj1xPPx/ohWXzJD2q35RlCpzPwpNjrGBPgQOKKm
hH/GVb4BdiSv/Nkhx1PxFi+hPNzhfT6gnKEmT3RaPo9lcRIEheE1QKb4IvKv
tT1V7BcyjRQNlGSOcgfRrt13bsMtVeytvi7Z3G8mUIk1FJs/gbf0T1KqtmBX
k1vCcE0MrCj1LilsCpFcrWpqT+F8iBycqBOhI1awYrHR611U/JkrKGxxoDeM
cAwjtKInlu1gBrdFe+bmNZoqukZq2L0WOK6tT6CTT2p7GPOuoKyHYflXfoNu
ZmVPoZcc0zEh0Naa7I1hEIxj2pplOwvqckcr/fi+ZFMqSEA31kUtUpNTHV9t
JV+TW7HqnLbJWQF4AZ8bD5y+huAPekoRLG2LDX3MWCI0wUh6N30AwSPNbP7o
vZsmd9EK4U9Ud3pWklQviL+mK/LW8MZnp19fSVd0Njh1NDu7NfiTEawoXb1Q
nhCilANbADTpte4nFFGHfAegvEz19/8FsnqXOc+ZOHUBDu686Jn5Vzcsc+5C
9bFNlFllmWCE+4JgTkKiTeJVg0wjVWkgzZp2y7XEmZsMbGbwVzbGhSNCez9O
8FzCJ6Asnb/OMoVsP2b72O1Q64WtvJVil2YmsPJz+eMUhLOT+AeFnJ8Gwxbk
F5wn8VWKc81okQnMlpi5qIU/D+gG61j4yLbCM7xnSaPtqQLUMTP9QMd/+w/3
TXXIrdPCVV8/X1NjKnRwaENVkcVExn4pak/aaWGEtQxMflujRu8XbaOwnIiA
6njr/Hi4xVgKKbAdIk3841e4nfhrVgnAZDLnAb2zQLp+LKUBiWL/+TFHPRvU
iqdVMeVEodWv2+GhjS0wd+uLYeLDo4li1IFJ2nUJEOxu0aRsdQJsGen0Bn5B
ZE0hIFNdC0E1jjpPf7szf0nTkfpT776+9D5CorTkfuQkQ4QOiv8U8vt6qzRJ
WcXfwdA6/iPNqlGYG+CBZ0yzBiYBoUtCEchGZctXfvkrByD6/ifL1texRqHy
XlyVqHA+epNrEXLSmoYaaTMsCJpEydWN/OdUD3jTO8sCaltt4ewHIkwZ+PT9
ShFEzULy3wpIjPyI9bdvSnX7OWqyTnGRF4vgjWgr5pgeT6uFQSwWrmQrUfdN
hsiUZpq0Br4TofJdBi7tVLuyymGvjN7715wD9k+RtqbgqCHyUW9fb66Wlclf
WxnmizROQyifkvGaRUzaKS65SA0Be0NiDiZq1nPQtguJgfyntJEalO9PSJ7Z
sW0UTm7WVDWSeXiPGmda2NvjkFEWlfhBiJSq8Br6zdezFOTwNmwyXQt5u+/N
UvWPTYbxMNPCFmivICyVHhsHQyLESfOFISFPecSd+TDs8U8GK6RqOavnBshW
t13tgyc6rndowORUXqWoBa7mGNeMTHN7qPhBKlOrBeEiJ0uCulhJF/ePtOcS
Zl0tNa2sGZgl8S52JdFoeYsfEtf42bR68bX+54/MGHe2UXOkpotl9EqZ2tIa
cppP5B/cBvjM4gZIKT4rxdMzcHp6+zluV+uZ3r/2pyt7lLTpPLF3dXJG+1jC
Sf2UApapx0J43/+/RbkBOAiUB4eYtp89EwHY60k4kqqfvxFqSf6esv4RadYj
zBX50ndmi1b1fqGrN/u/VT2oyRVDyAPjNv/ZIsrU2HbVAsf5FWOOFnoWDplq
wTnijm42YghWe12WMAu0KDUymQC9dqksr33JLuJvhPMYY2qirG0TYmRH/0FE
KHMCQrNFc5s1gCcSNzWJSd0c3MB0yw8k22d3f8qWN7Dzz14zowJfd9qoZ+jz
bOepCFNYf5OrR0i35uCEGb707Nzwm2KAe4FKctbeq8IdW3aS710iGAuP8EHM
DKg7sf1yIgU2eRYt5wrS5/Aj+WnIhwaKIaoDn+zUN6UsrXMCGJLcEej1iiff
IHII5s8NgF8/UrZppQuUef6raVW05EvVWp828cCOUOboHY+sGAdPuMZEBZPs
Lo4+d2MGSjanmamMSjfWwk/6F+zGwTRKzC41lD82bIdFk0wI9MaAMQirBjMa
xNPwaJz2Aaoe9wF2C7EXzVYXAjHxYZnohhD4wjfoDFLiaIAI4swmJRy4j8v0
PWOadPCK4V67FvA/bamHh/VVOSVv7tXNq2RMYp3klP9hDNSpXVxUOgqgJMF2
nnFpeR/Gqq6/gGMo1iLbFEZ5E6+z6y15cqbFgGwLj4wmY5ew+dIKP/qMFh25
ah8noXfGsbmzEkd9QfyBwaoYdN3GD1+7DNQKfnKEm2RpKYDRlidYKkG9BWTJ
8U2UbVrJBTR+tT4KGOU1aSTiAYzKqQ12XpNpoI2kJXMAxULXlJT0PKQOqK1E
RarLwOm3T/28YnIByuxlTXrPNcR8yHRgqX9Y/89+RxMXUHUWRKcypK0K+GQS
VheOLHsfAWXm2Vn+NZWq5nUsc/SrD+/lv2cYI+N9WithitYtBZFt7sSUCjwY
mv2wvoO3vU8QNydhx0KWuLKLptDzpLgQTdFKFjjjxCHvz1e0Grq4Zw1P5hLr
GS29HSYWdPwYA4RggygEj4RTN9qMf1hfp7WPoPNDB23G6bk9/0mV/HukSGyC
wcSxXmC1HmNKeiG8Ji+/RuKSjzaFbiDnp/V9dcvQGPRse92M59lp7v843bOM
z1WRypCm6MFrMH3fXZCzcVhKpAUAX0C+MCLYRNojtB23CkD+sSuP94xPH8Qu
cICrwEkdpj4mJOafiklvtNVO21QgOQEFecWzm5CTPGuAYFWlcT87u9k267/V
mKjb7PMy+7BvFvRms/H5DDbX4n7sf3j7O5faPqPAqJ4zSW0bty0Um58urmqW
HtOS09kdSmuRuLDgsaPWPZzX7FW586TRRsFzcWyvHaDqg/8TT9NnY5StVZSx
82yMc7hVXomvZpRmu3IDchrQkoBLD1KXvU94e9UOs7MNi3FGzluFV6JuqsYt
uNEikSANFGe33EVVqEnTlc3PFIMGiWEiAweEq5X48f34sm2l20IPP4gmAkcv
jXnKkpjmlMPsWJp7iZMbMPeNRuf1HowYHF430ZLSiyCJbZKo/Ai9XZCBawed
IFLuBesS4F4kqUPKJwA1vbxJ8YroJNMN46/oIwWoIxjsQkx5NvlR/T97IKC3
AmOq9+7otgl0HqkGFtiHU+2vX/m8byXSFQyivHM/KxTMLPtQInYIZQPbCF8f
1W1QN5ckYklCksSqprH1TVyp9Wl3HHddwerq6kbow/4o0jIqfLRR4twFbmDi
I4QhGHlAHwqwG3e8YfReCS/dQvri9i5CtAWabNTFhm4Bgz12SLgYpcs19G1y
+FkDi/CqbquLph3Tv/UyfmjcRyqHdXJHzy28h6AQBBUTu8iuDZf/mfurO/NS
hsf/j2r+zoEPFa8D6WMwdhqs6izigoy737zU/Q+rQIEYzGF3OjmzLVlOhm3M
b1ioRyz/ECdSQi0MyJdCvs58yaKr1Vg4G5p0nnVAPqEFZYTY8pZPZ8Lhzw0+
aVvw2gr4VU4AfKFenlEEwTKUFW/JsAPpaXO/hIyuzFVLsnyzO8VdymBMmpLw
pTKNNxn6ky2mHzuIBjwXiEXKOQciQFUWGdkpUmCP/5qqopWS/GN1vJ1UKc4W
LhaQfuKJde2EzvS7v4lSJye+Qtdz4rxPImZC2GB2K0BRddpfjGvRnnVLSuVg
P+ItNKMGBLGTYC2wXsODDIjNAcHAP5KRMluIvWV43aZ8kJYRaDa4NFkHrBn5
qBSILOMNpwA0OslzT6NldM9PI6ZCcNgHnkEEtTxYHQUOacJiYc5ikwR+9fIl
DRih67XES+gHHvMX2s6isEQG97F6Faio/gKnFFqBQGdBxVWrB575JG538OBc
p+laWL8ZKxwP2hCbYci+XS30JvvSXO4+u9htHwd+UAh4+3TN2CfG/Hl/Y+4b
oYKSjIfMdyA2zYdjCQZ3DKoNV7QcGagfChv6pZhv+VJzv+t+8xwl7STaQ8UZ
7h4OQ+n4LckjxaJNxGTZsaUWP58nOKOqRYnaFrf0pCQLfnR+RvZbXm5uWHSw
gIaZGO7tlHJt2hjYE2nPMfXcKCeiPMmbUYi25ErQAm5JQY9MzXmXbgH+EBBQ
5WCVQxoNpQhmPOdUvgNb+QZRvqYDscLBODKse29//C3o6BdHHJkyHd8ZsvDx
m4m0cA1qdzczDlaOmi6hzwbrZt+CgJq2faaPndtEbR31jxIF+g7PjynOxsTe
AK5CM2LcIF+Awdso25MZLlinMnRMrHrBQnS5kqd+9ODtjsk4cGYSFK5iMMrK
YzuqjaAfK7IQjmk5caXkFxHmTutnsJ3TtsZuI0QArXgegKHrj4EuJDl9ojZS
W2O8tH8ef+l593t/1Zzb4+ga1/BQN3tHp9xZhGf7q3c0uFq8elRBqtXueTz3
MNcECigRozlLVZaCal8BwVDQpQMVARSdBhrx9yWCYbNq5weE9ySlHkup2/9r
9OhfpglRNrZZKe7rfulmr5dziXLD8Floi7hWJwL/Zi6t3GZTLYanAo0DQLoi
Jk4bSRKb6vqYOo2Y4rvRDGDCuCgL6wv68b6yA1CpubMsOq20QmBggwSpuNzP
CUfgZDQlnbREtPtz8Mis2iSoRJ1yFkdUyYsIj1o+el6NemdiSCmyUJRiFdGc
JlRu4kbl1Tzm77rMAO9RHCjAoTPyXUOUt8FtI6UpMg4/N4IsqnPia0xj5ZNF
aMPoBXZY4UckcC0Nb1Hfojzl2lppFBTAT3QlfQYwk3Iqf/s4tBMOVAUxwrMX
qgyAK2ZevH72jOu4Wz6u88AGsz8168AFdb1yoYoRy9Z0W3aUw8n9tb9qYPTd
ujsdkypUNXiocLTwdFhgR7ErxMjIoK4WtWCe+i+cL6AXEP8KB+2ceq3wlrCH
E/6P4s2prGsF5t/VAQVsF+hWm9+SF828BqfXLFy6ih4BhCGs7gA3gp0ZgWh/
5R7GDIo5jcBHKSMyr8E65zl7Nx9d5zrqwsha+wk58caC99SqKyj/DCeiyNMd
XO/7j+QcNLF+5RWeGaufFRCMLihlXL0o3/LxIn2FMA0pqkW9uiWogcGsCuoA
F8QUiFy7E+/dKYdS28X7mWY3gfRotaY9EUY3o+yVLRIvAlrXXxw0wGZY1JZH
UsDm7xbFoikOmcAClyK94I25+jrBXRo3oRjjBNrwwxt1TV1tI+PsiS8/kNd/
hPInebd1ltBvbNA9filnJ+HDZa33ZDG/RjUmpwyEhzBVMv6JOLjk3NFkkCxM
7nwVaCsqaJwYD+bujBMMSdnKOveUIWO/ROmOcpZatzeOBFH751goPnTmilf9
rwVdgaIgz3reZY0L4TBgubNL6djjSviWwsNssPM+qAEDwOq6gJM4fWQTJXbv
tHp5rBcv1U64at0QZRfIvckX/ooMFcDV+n8GygoCA1h7oz89M04fuNLIL57X
/gDry3K+Yw5JVMldfaFA8cfor+Q9KmrPBOczE7WchH6CF+9zW3ZOVbONyQ4A
FgHzb8ZaNbR2MYt6VQaV+Zhq43K1Ikvtdczl82/Kep5+tgw1vTIDIBfLgSOe
RdZ8P90qZhj2sgOMbTaibN6XicuDwxGLsgVXd97kAPjUn2HFMCpBJpKq3CQz
f6uh67mvaSCqm7tAu5mMipMH46M+RXiXBhpckqqyzGa7kBwPquBrM2OPi8CJ
4XJA5S/b42Pl6Ee/PIblvE8MNZra0t0+6Y4fXi31h6LmxupAm9BB81xuw2bR
tS4rdiHDj3k0Zp9L+nwp39CX+VDQNHWOLISo9lWSgSjzpQjzx79grIO+sB+K
9Z7aH7AtgaHODhiUxB+m75bm4FcHfMiqyWEoHbvZhtitoZTDxD20evtdHmlz
VYTP5DJgIvcDS/pjJKwA0a5bw/WyPh1unae6Z8NUP1dZQw0q0X0ViG6iT2Fl
8PSUu+gPbzPMcvccCIacVWVobLDK4ANJPYn6ckLrcGzZwUW4vHwngNgiKe4B
MrPjI9UhX/35wm+tG8YMYzO3s3i7o782JFWwlhkEVlx5/3MHmYT3t9BqCA+N
Qq2Xvb+OAQs2P67XmI0pPLqruPnb8A4GdvjsyrpJcmaHy0/Z79sjmampJ2gw
lZgbvubvTVZ4oK9puoqZbKT+8P4qntmrVeQ22oHo+z9FZZQdCq3g8RxJlQTR
4ahEv7FBPqz7DYI1fOBelrVytP2k6UwHd+3PTI4znJAo15zN2tU9oQ5EdDdl
md47d1XoNX8Od5Z9hu95g4yCR7QA0ynYW6YFuYUuypap4swwXunE6+5lYcPn
qdb/8r4dNB7mNJpJ1iRYNzezHlzijmDd9LxDsXi1MG9NB1WqsFS22LNPZKOh
1D/E2NzBPcqgfte+PVRRPguXMcT4nJFFsiVRf1v5pyaO0GbiQqlJFTyNPcvr
L9USllgIEDXjiThm7+qdzEhJ/273+eKdLLnkSlD7e/GEdw6rS+BuFqxPK/ZD
qWZ+mWwIK3qHWshT+4qnflii/KEHLQji1cgyH2+n1RIoV4w1p8ZH6kVMz6dK
SIV8xj+au5wh+FX5aRdnOUsXlNp6ts4HHSz/G11lEDH4VGnuUEyp2INeDYYX
NyiXE50wmoNN1LX+ZfLlFbnb0/Yg6WgkzKp+ch5nxt0y7k/y52XUgosVe8To
GRULEovkPK2BeOJ4We/sDnYRJ6mIRFhKSAuwkZVHdmjBu7T0x+8MgkLt3aIf
dccVm4HELnPCQQVGh0fUVjBm/6KSIrwLAWRNwcyA4x9U+mXahibShHYsKqPA
N6CvGVPAbSPMfMQ0jFRJs4GVM9Dn6F4xaeSftyiMA5QwlC59kLtdfSz0R+s/
sfB+yqXObBOGSO0w77XZK/U7GJ8UGQ2uE41Xes9LLT5MsB6xf89FnF1J3MRx
QiKcQW+YbCLCuD1+usLrJvKuuflGQlEolPbEuLKoWlpSiBirpULp0xIyN2b0
mGjZFyOisjbF01K/hGmOiHzfWudP5lS6DJ7NQ6AZAlYGQwnuPE1PTDG/WDMD
W45e4LgMg0EsvhboGvPXbUCf/Nigi19irKWRWfu7UXXkK0JpVnmqDcJTgOqH
FMcintI6KMm9dxZghoXkdLSxu8pRStepmKu7y2hbKFyMceIGYWaiaTEyhShe
5E5F87VyBJOlkONIyPBR2paFb8k+y9a9TYQJIp/bfEDjXARp0el1xpFKvtdW
pLGeWpEWXfEjuxdLuk/gubPJ+7+FjW/DjvtJwHSFG8ATlT4wNNB7CRj2kNfd
g817LGszxBPxpP7O7P9YyCrSuyfOMIX5ad5rnyWE3mmpr89PCIZwfUe2rUaL
nHWX4DzymxsKpRo4iSLJyXcIth2nd5Yt0zLacpI0XZDME7du6YTZ9cXiS6X/
ss7zSkadZpRT7GFOfPO+OEMKLU5cizjT+4DCKDHJbfyeq59sgcDv80SFH1oO
GAYfFAUnO3mQJqBcKArN5CIlePRuD5wYp490FNwZaLoXotOMExvObSeHiBxl
ptJ6+1YXoN2cya0H2LWbIEu6HxkiYVAbSdcJ4qEWmq7jlBsT0lrLCeOfWbQI
mJxg2vWEi8Hf/W5WnNzMaNLNLHAKNoGY6IWy9dibUMVd2YgFWnNqYaeDNvsn
cCNoqQFSnNivlVru9IU1Gxk9JnVp+oy4ZZ1/8YjMjTHLSojK6BpRVSWrcYqV
of9iFk3VcwjtUPnwU/hWhIz6IHn1cdLBFuyC5pr0J3zmj6jNR0Py82uW+Z5z
Dx84ivZhisgI0/P1Jb2Xyj2GbkY3g36EdMIQtkVROIEjGn7gcSnThRSzp1Ve
N8AMkE2pxI9tf7JM7J/yJ5khfUiLzmL4OpyMhz2oJDfAuA6uknDwl2y2ufF5
CeI0Qp+0eLnNS6UHSuJXx2Qx6TB2ftWLaXwgvCL8zD2hq2nWrPc0WEVZ2JKh
Q+KPQSpiqJCMN3QvOXLVYzfWaua/sBI3Sp3kI0/XV94eRvldNQi8kDTdEmiO
pFw8JCtugsf8Bs//+WqOgW4Ow5kUr0Hs+z/V72R5dvnxR8UBMBo+NW/jlosd
h3J1uG/N1OaXzUKfzxV6OE00OJtVbs/2rvROxW1DFdmXnIZboC2z+zDlz7DW
Te7mPDwYhWMO+O3+7gIc6+vWYk0HvSvpf/Rm0GIesetV5jMJVEA4vM/cEco+
gGDPQSBxVHdoxrIWdi6ReXC+n/6MtPyUpL+MdBhoK6qHla+vnokZRLeBpiKM
3tsOZ7IbD+q185BBg9MFmCAnlP7pX2IH10WvmqGpi6ljW72aWrp94J9TeGHR
OkB2B7nG+0Y7WGaymzxFUCLiyLxzhMyYwT3eMRwy1HeHw0Jtc8hwoHlKJYoE
cF5y3FKre8jmKqiN7lYuOGIFuxTVIBLfOhAzD5Ezftabnrz125vzG3/i6Ol2
zLM981+H+7xXxvBq2fFeX1yncL4XCZFEsPrefyZIJxkWcgR8lgjHdLBNENms
gwKxiS8CnP6kgQ1abqk8Kt4Ly7IYY8Zvw3iqoPsrrVaAXwjX6Pee7K/MPvKU
waE4yVU9ZxE0NHNFhPtC8aJIBgiZ/r22AAe59aw5gHsu35uS2s2Zl1IA/Qhe
zEZkdO0lH4VXUIju1IKNbL9ZFemYTcOoOvZ608ubD4UxP/uUgIRc8TOb/eVN
2EW3J+d2FOdabVJ4RE+p5VBW5f1J5vaTQp1E+tksplHeB7MYL0ZR2A1Y/3Zu
isriXYU8So7tKNbFgeFC3rWcAahGEjillKDkgIg3cORyC1VOn8qfvEdErscP
U83D+a6a/ETdwISO4XmFTxza9dtt1++cS76nZm9ixuf8CCa2HxQHSnOABgKO
03yiXeRviuq5xSnhgB88tMe+JM+h3eS4/cJnYjwEpp7NG7CP0i7Qy6Ab0qwn
CtNHq10bx2/gzsmLmgemFXds3SKySTyjVwYtJMHf95Ln305T+Dn2nYHViDjk
k7be/5LB+2VhhrqQVp8jJVlWVmhbHBiCDwnfD5GzrWBzX4Q+xmqp4xY3nmsx
PrQkfFR+BokM82e2fNkMPkPTLMSdd4TDuXOtx73V7+0zPf0Bd/fsENZRubpB
WbbaPLKBAMvyRE6uz8wgXXNSdLVRay2Iv0UkSY4qrQbwwnc27YnGeNVSv+7n
clO82UZTtZVKWhAM8YQN8HgtighdV5dkHUoMrOFaB6ndU/vFPogRKZCPjsrh
V9uOxsPi8iADlF1xasYBimjAjCMzi3JqEw/TZ0AXVAwCKb6rp6+/8iR7Z6IO
9UQ94emdKBMoDG2V1u+/YjqzRmatF83K+TMpV/TXZCt8cVlU0306fWlrypi0
t/Gx0AlolgJutSbByb0RSe86UYkaepqChWgIFn44HHBa346BBU/VfDCPXxeI
TA0KM4YZey9NbC6D6Fjor5+ENOO16JGbYKvt67u0k+Q4w5EguyuS2dWvpSv0
TWgWfBhNuGayqVXmzcSM53WGsz4NusaZDmNEFR+jXuo4UDWFXVn3waHrDs+l
tWzTRhblevXGIFUOA18S5UQNot0W1+73q/NkiE9+N3As94CGrjiVlJp4q1a5
yYW0mPVL1ZEO3vAhQ6zJ10HmberYwuAOJFqu/1O3BdAIPQC81sCicHN/2QM7
phN64xuhzyb2nM04zWcaKWtGDtPuNtUsqVbQKTg199c/miUThfnzT5NRm3tT
zyMdj4lSQGnvtMLf9vSvXxNvcTPBqoq7fw3itBD1qwBL21Kln+SqRXuwBArC
Wgm6srgo+q0q6IbvGuEEVzBxyp9S9ElBjtsWpslqU9loqqCPivTIzsXoZiju
MFamVC0EF+FttbV0i4exk+4pQ9WybSg3spDd8zG0GdrqsrQntps/IbtGrDWK
uTDN1O9UqjcKhcKAthVm9jD8R9iBnMN7rOrYoZFqdHrc5K2y1DbO/x6oP4/l
7VOgCDxyDVpe8imS/4O51ya22sjmxjioELS4L3wb11H6mzHTtlCLtAFkPSbr
hKoKbHDa4oc6ZyPNKpFtUemByVEjBctKhViTkm69N4eeUxdxjI4IP1C5oqTT
IwN/1JhukBVL9yBUbZqqR7gABzhld+JewCTt6Z8MNUyC9pmmlZohWLSZvj7v
jaSVbz1fpnu4n7GhalBj5CS5ovrAiQd7mQMR/zpZ8M050sdcQq6ODr4mlstn
8NxUOCFtaoM6RynjLnLWEyVaza0vmIlI6H4+Zt/aARltS9l0iMcbu0Wcg5mF
vDKQU/oZ2+CFa/cGr2YRk8VendyFOO9AhYD1hxPHTsaREequtyzXGUCbFB8e
ykzuAA+BteJYQ++yzTeCjdeeQsNWDkradfOIHNkrPdr56ULZPZwUHPzzCWcn
eB9yBlJEz9JACapvWADgHg8LlJ/jUsUwVLcXaZMrNYOWT6LRNZa1lfe0nnB3
haief08wavZPTcL22mCUjIWwmDMu1WAO/4JjzEug8gHq0u54OLejbYJTsSHK
AOGViAM4btWqZyZ+XeVFVFosUhnK6EgiQhKjE+ZeS7Fe8xkgSFdzO2ARZqRh
mjWBkza2gs70YsiDstErFmSBR0GdauHzGDlDJS1grgpoA78CBw8KVbCQ5Ly1
ChZJc1PPzwX9PMuNj4yNb0MCfZN9sNJdURQ7ZuLBQqiaU8/eqgZmKi+p0ZFU
tsdfI3F+I/i5aIvD8wK0TKqfVH8UskItX9AU6PeVIe+aldoGgziaEnHbSF05
5H7R/mqsqZw/ob+wGMrBiXOAV9QWRXNDHNT7DxOiYEnEf7iKsq/1m28wOp7s
E1g57L8ENwn75q5frtqIZuFaluWPjQVr0JQ1QmPFwS+woMytJTMX6LeogHLb
HjhK1I2Jb3/JzyhXQuf8UCB03RReH2InxWQE0hbgyj9VlZv7GnwfAnv9dgBv
ytMZKFakciNxI4BPOuaIMhpiYkiJks9C0Y5QleMYPe6IN1LttTwtRhrcY+xh
e5HLlcER3d+MQ5Z8dN2i0qbkB5Jcq6UJr05GCdTB45lYeDTh9ex2Um2NYMrW
/VMWGRDTtQYh7/F1/XibDchT0VQhTTEN/DZGWLHC4ZY8VEEQCLLY6Mfk94hj
cMVm0CGYONpc2+HqxlH1tsMNXYiK82CzFdyQAOLgAgyiHsoh6GReczBHEBxM
DejxQwnO+BoaMfsywa6n5MM5DMgdiGQsbplpvYYgo9HT5YI+/kdBj5hCa/bJ
/bVjHiyQV75si6kEl51Ae8fTSD9KBysPaA/4u0FM8iCxGVZ2II27Ok2HECdU
mZbU7WHq9WYTCLhKKvBbfKzSV7EbdGRKxu5hIoi2NK1QQItUMwbMuIq+DqLY
wpO8n3IQy1cmOwdkXc0pOHM4ZMWUPi6APAUFBve1UMCoByHGaQXVwdKsfHjK
AEo8wSYshLOCEdZibnyowsWRE8kIRBPxduJghS0/qiMtuS3gCNBRkN7OiYoh
ltXBYwbMV8seAR0m04bmLqeEyAQSxpCInhXaqHmGa79J1kcVKGMSuovCxb28
lPCqqizKC6lXcyN2US92lyCokxCH3Pk61QQ47QvB4GPTXoZDqfqo6Cf28k+a
8Jwg2wTy/Y7Xnw8q04Pmpf33OHVYCAwazBs20v7pgnKcS4yyGG03+qVhPEMb
U3XfcZV7Ojgu4C5mC3wcWi1Pio6O0SRlKprLT5ocR/laRo6eKGULhATlyqsd
rILDX4BDAF7K8kW83EGmThbMJVA+uDYKt/AKm10G0J4oTACPdi4wmaYCGHRn
kr0SMU91FW0t2YxBemtwYRW13gdQSH/GbcdlDIJquDrxK04e2W91itigRlZW
WEHFLZFeHJECsgjnBGvCc485Jkoaw0TUs3haKF9sMyFyCYx044Zvipc1xL6m
Ol65D7TFpEUxeDMOeR/9UXCtxXTQoCTijMFyLisdRb5JFqZAYE9i9dcLB0rO
lMUaw+LZShlbIQYUIPZOh0yAONkJhGHHbgPEp2GE8eyt4BMHdUTwoI3blwaD
fln/2EXALYMyUIA05addU+N/WkSVc0ZuEidZ2wLhYOGAJ5F2IWc7l3fFqES8
QROuFhuBNpWkNLSVzSfbz8n+q/rOfKJDxLCN22FgPaveYlUXxcyuCRbhA/3p
TsPSc+adIIIOtyYAqO5BeFuCCXRevxG5kCNyr5V0YIVYCDGgKaeGUV9G+4nk
9gp8SJDZD0pYB39vYdBwfn7Rv6CNUXbdG1AaI8LkVXnDICSmaFdewfTHhHK+
f0tf1HkFa1jHawumqIKJGMeKYwMptA0C1xXabLxbPEfNgaoGeJoXa7rd0jLu
shnGQqRjsfvnsToiOCWPZdQuChlZ9wrzbnm4nDAEWzrGJQ9Z/ebz+Tz43MlJ
4Asgy3tW+o7YC0UMfglhVwuEmr3J8NMu4bY+cL2vuNftV4PWZz/Cq4WVKRGH
gDF1gaeHM+oMssQ8sek+cZJaejP87tfWRTnNik7aiTgGUjDDdXXY0xZbR5c1
zVrdPquQnrJgJ3FKE+50DWvl3GUbZUfX1vOm8sju4s7lVv7dbTAePyfaPtwt
5vcA9p+GVOoldkZQb6LH8yTr8kt34I04BQ28c1EIAq1t9TJWeMYsA+S8KJ9W
CmTEKmB2OrMyzIBgAckz9atWkhqZos1JU3MRyQ6mQ4VxYAvAV0AXOMCwc0sx
lmv0mD8mJQW8743bYgXDb3cbyApPrzTWD8QIK1mA8+8oa5unGE1FDODHTD+x
/Gr4zjSqcaXcIT/Aaf2zsbpr9T8Eadq8HyD0F+tuvEoBLmKPdO/051FQaYCd
S7hv76+u8N2RJ4XTkLJSm5MXieokeR9uHUy67wahR5tqPZBQF3I8oDQiBEgo
3buiowGJ+hhF5xz1H5QmyLrOH4lMRxnGDjNy/hO7Z7SNGi1GrU5X7V6W+ArB
IrqbC6cfN7EYr6YzzT8VSoOu6boDAAAY2iq9EuT6u3MXl9OGHsctahLBIw0p
K4ePBHArma3Yv+Y/fEVw+XPUyVvMkqRWmyDs5Z5pnXhmQiu+1i/GlkUB2k1/
xa02hA92k6773Tj9wcSDg0ViT3le79vdkOO8e2NaTwaYMk+DNeF//BclC3NN
/GceYTOvPNOU9YgoxZoAXiP2tWZTICf4Da50qJBNXOgMFpUgNJAq66NK/sRw
GzgvGzaNxLtyVuQbkJjmrnyCFxfgr3Svt/C2nS2Co46B76dYJeiofGxWORbg
MwGrrUGrVGPUkLWT7IhWFWaE2gdZa7p14D0JG+xMGJ9dLOVnY/R0P5y6rQ5w
Dmh3XO8slxpNu6JUxBMyCs3dDsf7JE3uHcdTLuMqZ8MjcqfNNeAIKizRwVEb
YC87XrIZlqXF9YoAUIw8ZGt3mSm4v1puCpQ/4CkKS3n/grAlx63l/7swl2TP
2ost5k9+LeFWIr2Hc36owXk/+beqTIolrLrJijDSXAHVE24E8jrcNBnzgdkw
kh5I31wdA4knm49rQ5SmxkgpjDoH7cV0HLuTBJVRrKJndoSJE7WEZ0PhtnIb
PIWCz/5SgI4qfEtnoytYigtbsX+MI4W2RNzD24Q+gCkdIymyBkrq4+T6h0tw
nkAEBoe2BkzubqWrnpHdpS7dzZ0s9sPAXTXiqJ6sAXiEjY7g7g3nziyG5U0f
gUsb3QiXG86lMApTtEWiMAmTYAZRogbSXis+/SHJv0NKxgpsqkZx7YI9N/im
K+jdRbLF2Cfy/r7iE7dWm1kQx8Cg+F/3ovK8QJ+8taJr/+EphEr4bzkBkpYN
sYDpvCRM9Qp8r8dIyKKHKbdQkE7N8NQ/YrG0cHe49JouoWIsouVNUp3U92FG
tmswBIcMAqc573l8QNFayFkLKvrQUsMeQKEQLKnVH/oK35PPXYlLcgfHP3UW
TYfGNz9cd6qJip9f+x9P7dJ6JEJswTPtXoVq7RwkiWO47GLGBnAXZsD/hbBI
JoZ5wbbDvFGNNiG1UfaRUeWSEYsLjaIjPcoWpyu0hmrQpZwArggN1uUISKad
dGHAG/wNOYDhzIPmqcZictBRoanqOypdjlgwzTrQll977wzjbuCugiaFBvvM
fsszwRv2qxbfJWZoIEznXxu0bxHVeKZPPqsQOIDkSt0Onv0G4GoKNP72xYaK
0+5aDyms5Am4/k4pNTRKOfHj6Xx2obc/BbbwofZopj7XxkEFuXDRyRkk8Auz
wDu7Pxka1fGhjZiIHYfS2vmT5O7St6agzIrKsVZDJDuhRKso1K8ypz/MFFUf
YfLr9hltN3cBn0UxaIBWycv/Ew3R1nznFEnefgsjpsMJqIFcrTE24SVTvAl2
HVXmbRyQ7ZRH9rU4DA09K5TIFDjrmsLQ6q2tUgeBrJDJBUyQsKIyaAtyAD4v
impdztWnJzw0dXw1iK4ETCyggrwOx/uRoRLwAGpN/LMcTvgdgkFJic4XDbe5
nI1mGYclZLSmVPZMsiyhYlcqAPcJ0b5ecvrcrfyCWDtkSc5b7+2yZTwJENxJ
qC0D2XIJwnErPW+TJkgXrcJ7FDHmCamLCEj2l0Qchy4EjPe890K9FII49KWA
eog9oFMovZ9pC6QxTDEfpTzV72YW3qHUFOVw966PbuJHQFOcDzsk+a5m89ob
674xcNAGN8M3JhHVS9eptzJip5ZW0L4loK6kflSqWPSXy5Pn1ax6Si2FYxAP
8excFkeywvO2XCrjW3jY17RNabwIKAJuiGZFYqIZIE/gHxm3HUdAcZGwtx3n
hNX5itZ7SkNGWuvAemaoNXmIcOqgdkhtjXrIAR50sY/ZDZJb0Eo4QO6DKqXI
q009a7EqoEHoRlfgAkBSR0swaR/On8zZ2dyqanLuagdguNLaQGbzQMf6iw+p
N4XvAKknae/+uO9mIm4nwG2Un1Iv6+SVrv7K5rwErpfgtFKGKEVDwfq1RxNV
U6tzspHcytZJqH3QPv75m3E0joTQViaX11NUf/nE+tLx8HzMZnGP9E8Yxi29
G33P7x4WBqgI93a0ZW/Oidw3+Vj3AWTd/WxDRITMC2RhaGnkX+kQPmEFmfQu
e20xVcuEh/cXS/Cduz3CopMuWLoVeqI8TOwutu+nzf+SVXPLXhUOM/FW1QTt
FMaHJ+JRhcfbRemyXxuQ+Wxo+ocudMb4QNIDT8ne41SfBCShE12hHhHHrgmG
XoPf1PnSxp0nCGz7kZNaZbpUGrNZ09M/ZntXIB9BkCtZH2BOkpzAW/x58kUk
ZqYZMEioRlX8cHDi/3wJRouWaTHcN5tyHTntmNDu1MN2vWU8SEhIlmeDtJAK
7D4LK2TYvkZJn1E0VtN1SGkoROVutHFobUujmF7heeEjpkNS/c2oEANJoyf1
vECtKZvib1lF3+n0RXwH9hWMAABnBavRKohZLljHLcZGWxBLwb7ZiWqy0f9U
h/JDkpVYsorhRKs6LCkgQkHe1KUDc0BXGS0IrjHaOWnIOnIHAJI+bhY85/6Q
flS9/WzSfUChaT1aYS7v+GnSktOydUR60jCPNEuxMWSUbDLJgU3579i5pPHq
GMcNPZa4znAZxnMVD1FFywdQRuDs3b83gX1hLsWQxmFCuhck8F/4dg6yB7QD
vMp4v5LJCmTqUmSVicrb8grrpNcK4ACIPXf7jSaJjdEp0PkcgnWlhC5SRD8j
vtFlM4VZ9E5YUw0+rONpJ0mGetTb21lNlJsWCRyoxpowPRVp3a7CwuYaqPcS
1aN7lSAh6xEAxBz8kszhalaBkV1F/wepre+UlRabLUN4639L7FWISRIFQNEn
lAiGjzcvb2Dd9CnHMM8yjE2iSh0RIzb4mQhohbD50GoN4vZ0FwACd4zyJNiH
0mziJVO1lIr5ckS6qrZxMP9Km2Ghl1RrM3Qgte8Ym/bDHWO7biIlwr9YFPFF
5IZmnlF/x2sZohiEikJ6azznC1qUtW/RXTi8Ga4j7dDRXRQHj2GTEWcJJGz7
tvri+QqUx6516gMP0CIg9B8Vd2ojX9I51dNqiUKRcgpyR/k9+v3eJ6qCv3S4
w9MeGXza7XcnXF4rvFHV54wdjfGwE/2DoAr6fxxaJDfHanqw2svZKveQJVJp
e70qhPsyk+JI3wFNoV31+ihOURnBDnVdtGJtWGWdQf65dN5RXjt6gqNv2WOo
/Tkn3LpmkwrVhDQUptoidEldcwzVUbCew+Fa6vjmC7adCtO7ey0k+TiyvOg3
DNuAqIq9tLz3WqueTk2HAulb8hLuQ1ygMl2BfmIuLLPoSaBs62NtK/F/B6Ma
eBZuEWHj05rG6Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1LHMC5KmKW/mr/1u8Avy/fBOH3q22lJl3C8Aa1WCzx0x4CQKG1bOlRz1HoPOQ1SkdJZPQnUONm0clU4i28Knr5YOV7rk1E2L/BysdfRaT1JLdKpCGScqgVqCQMgOd5dPs3WcMnRSgRVaxU/AXDqTYboiBpm74FxGcpbX9Ji1oU1FtJI/LTsVOWT7Gwhv9bNl+OK8JTPhUmLna7WxS98Qdd7dhZx1JfxsSYxP2DOcwQnXlpaB98CYohCz1s/nuhhmIPhp7+kTitmYBADfqyhwnNbFeuOvTvJwmTJz1NuWCUPcl7dUCfhrB3aYprIH1Ap4YCx4f5XbM3tdvM8QW/goKJxPhTLazXew6QRApnRGNgozBKQ4uWBpuFZSUSRSpxNEmbcFCzVxOc/yv7C91rm75sigZ1jT3sc/PFmbVDz/ppoFh7W77EUAnk2VU7ODfQ2UUh3UG8xwA1UbQfAbyAPj9Pb5NTnbNPwLC46mPQJobnSpgtPdXHPeYeE2OGv2aTYyyt+FH5eF7xG8Lxid21MA43XajjXzexthtatdCfES+239Fc3A3O/FyZ8cJr4HJvPTZSh/wZ/fM4DXKNjzfvOgJjeCUWn8WrtW8b0pwxR4MMeB+d1ibEAxRVpln8GYNBfuxdDRWQAH8bXdElVgcPRvvL6ZzyxiHGHKlYOus6p3lkwFfFlLurZe2LLkVdfqs/aabY6NJyEVCbvHXnAMZfinh5ko9/6BgINLuMsFGvDuhUAEd5LTnO60hrOSSuWzT+C3RUGheQnFsPFKr0yzitLoh57"
`endif