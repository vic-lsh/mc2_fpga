// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0gDsj/x4EBtUQuTFgaKdSQsZvMrxBdl/vod0+k702sTp6n/Ox+Mmyz6sT3ri
pCIKjpMgIUjfBENNN4vhkC94p3esNJQDg2F4vi6ALlMbs8KBsMqeSopEWJ2Q
yFcc/eqw7WRWR30MyzqQ8TEQ6VIEx2DNDgyD2hf9zUOPrWbrazr6m8f5f9WU
iaSjyKgGDjOcqqDmUgokzn/w9TH8N8UrtkEw74z1UbUzBDu98F3jnHpWrsSE
Ac4cDAi+ws30oLxLz9yKE8IS9T/i084W/hKF25Q4ry3Zwz0nEJGu8+OGHk5w
iEWkLpt+fl/S472xk5Ttku+zC1jLlXnZd3GCZW+QuQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EkdYXxX7xG38c9VczCZesEIRy4dy8ntyCo/DwvSEJy3e4KwDXOHLhy9g/kDC
Gh8rZbOAXsoAJzjMMiFFHbJCQz2q9YStwdh3ErAkyN4tTlx3GiDUUVbSUqqe
4Flg5fkJXBCdkW7fmXPjS7ez/BCjfqmanoNSrRi62JHELb+QQr7a+hUZI6RD
BK0EI1Hfidrk3zOoEbiirGZAAWdgAxaU/rd8UD5O2px7dcPQJqy8t8v9kifP
Cq7wVsTJ1LxBBEkigiHnEhuXap0dHnC6QSHo8pM1sOwVFOv4SHW57/+FdYu0
mizOJ0v5aMq1wQiPRhfGqggqeRUnatWb2oKB4CzHPQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fq/OVRSKwj4H+/5E6hyQImGR7EAlUQxgMDj6WG+1Ba++9jvb1+pU1KgjIbAf
GCboovEBerxc/EAjoae1lGdjMkEJWBbmV1T+RTXVsAy1gcN2xstw482TPcHI
wzfFxG3Ovt22w3rzzcZcAAOPEFcozYpvAVD0vl00vqDWbAkiLlX35gK0ZbLS
6Qg8CVSsL2b57F1lM1isJLnkdUk2G04qrxyTofO5zhK1qJUFuxl9CaCIlFgI
8GlMAPKpj6EPjLgiD2aXDAKM/GOfSzccsj5jLpnnJUeQiRCKlJroJjpfhFTH
rA3n7rE9rHw/psWppmCPxmP87hFtD2BzOgv9aB5d1Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OXJskHjGMiz51u1QrZw/t7w+X3mrBoEZtx3KwqQ7cL+sp4FLI6GTE3qBQrCE
1xx+Thtgj7ib8+ShMLxJs8IPzOPRlAkwaEf04z+hlPQ36MjcgROtcKFhaJf2
1yx4dAk0VdvhecruhjnwKXOL2QTY9hP6KI/xsUqTtwrERDCLLUa4MrAOMage
86ia2Sbr/U6teHHgYYIwcSuDMgW6yHOgOWOEasc/IrQy614phroLoxtNJkRh
HQntNlREj5S24roBtUpJJjaAiXqWSQrOjQC0n5xU6mzhiVJiUgXnmpHDTqsG
dnckoC7QTQb+5V/Hio01iPv9ItnQ6G90jUjhPhE8Ow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B8gQkrnln1FO3a4oPMAX+e/Qt/95y09DzzNfFP5YSr37m+5Wdavz0Cx7Uq7L
4xeIlLO2fK2wvKMaQFHDHxlY8FHmGjSr06z+oXvbsOEfvpLF1450lR6cKDVQ
fyuqHZ/803ADtgbMYDI9MATeWQtB9gYOcemFLRWddAdGuXfONfg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZBdn+K9+CcJPKCT1j7Oq/d1+MB5nRGrGzOVEKiYRzu+/NuX2dsda/lQD1DKl
GwxEeWbJwyu5go28TRmuG5oQE2mPGc+y10ZxYf1Y+WL4gABCjaInzJ00kueP
LnR0lBtprTMATC16/kTCgBDGKd7ak0Ep3xFwVTFYKct9KuQgOov/hnII1+tD
sjiDi6ZxW8myFhgzRHUF2YChFABh1qzW+48kCDwOYdWCvCS857jAuAXyLCZk
I2npKIJXd4h0FLH/0+L27JPhb+xtVY8gskuvBCI3XWe6bPHZW/ewofBJh968
Nycy3Dy9w0NIKPsPCou6G1WTt2euvLhH83b2NR30Q6bB/UYGXKJKP7KViBNY
nefhuh+G11kNgp8zjF4qFExH/yUI7vqfMhKjcxRgAipaO+McxUxHd4iJfThe
VxSFUICyShU8aUCLUv7ogF2Ho2q+XrauC03chKnNzzW7gYsXbDPR5LJNWuNp
+ciE2Tf3BGdRdAIf3RHZ5E8v9ZgktuNg


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LAMEZ3fnynk0nNn49kWfKFM5ajOAq10HTydaXJYRVfasHT5kEYQUTxJZU4tS
yh4nLJEOpJSzHy9Vl2r8Jm+wEx1glov10+fA3pr/fbi3q/jTNVy6yLURb4qe
wWmBOf5DBQg1hvAt7GPAGmyI09nscba2bbIak7XWrsehc0RROds=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hADhYrCSkTJ/Gih+dX5+g8hNfaSg734CZhKSvQMQQNJjVadBehiytBTOkPIb
fOcQtbNugmZmyUg1A2bg6+ry4ZerrCUds1jBubzds9I2wdRNERr6tfLUxzsE
zo7aN+DQpEOc3ds10JOd0P3n9Uley3hQLcqDGvrt+CSarOwXDHE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1248)
`pragma protect data_block
64F3Abyod4tuqUVo/rnE4rpZuEEt97VXOXXGVEhQAWSHKdpVZClr5smp4K/q
IJZYcGba6CmLQMr6HU7aG7mNbLvA4catcH5CNwzLR06ge7ah18FB1uBouAqr
qpV9/SJK14Jk8Y8qUxz5PcNunro8ApJoBvcd6DgwXhB4pkEf8ikLNsV6X/+D
GO/y9JcicznRvnTo699RMANLP4AYZCg5XKpyy0HWnAZr7iK4Jfqn9LYHhLtq
fAsYAJEX1OE0x7hiQxogFZExDGQakNHDXkiYH0WV5oSvR7wAjIu5JYtFtqiC
IsZnHjAYtvOB0yQ8Sjy6oHT903ifeaDYl8CM35XMpZo5udXVP8wjePewjHw9
/W36g/xDQL8nZAzOIEkfB9pXNgkaHomxLr5DDS/jSipH32J2Bh9jUjEr3fY+
lGQm6HYPUkxXm5Sbjl8HIdgtpTtjyzULjpZeCpU+4GV7JBqse8+1uHFdRnHk
NTu40MPfeDaUzthRfOogHlhsHzWO125iKg4Pjt2EBlkt5qutpOjEafplImUn
0379oX5M2xblzRgo9xk5WB9GSiE+YPYDcQLNPxjFNm4VOjImZUKxmUc1CPiO
wX5KwjahEhKce849ZwauLldVuTtETMsaLd95UWGRYSRcjxArUv6CXB6g3iO+
dhlu/rVAmjLsftlGbrsZ1LnY4VaOMsY8PADowg+zSRVRdqsL9a7FsKlw8F1V
XTGByAyIqLpBRGw0JXYX9mTg3Ho1KnIbsMix7IfOtzN6JmK9YZVcrx4bSuTZ
1unK50u/jRaAzsJpcFCr0aLrJt5xvOLNOsYoeYnBcWOMhZz9sqMDogP40gh4
nclDGMxiBkgE5gcukTL8eyWmp5GGKOfod5CpNE0ZUI0l2R8YDzrz/Ls0NFKt
f+HcOPidlDlO48MCKrL0BJpYrvtvT6SVh4p604T9IsIa5Kj2Edni/W9IZePf
Ag5eRkszj6nY91P9pS4xMWuX15UgYKM2JrCEBnGcZlhtz6NLXTPsTZE0DT3L
iM3pfgqLxG+OWc+W3MEcmt0qG3X3SbYDvIU1yZQ+oOb5SN/vKPEAPeCnQ2mk
mEVgWGODgZ9gD48Sh8QaPpd8HTIUbDBGehtQqqHiQ5+x+4QdE+MbBGv7L88W
MLODCK76UEJ3+66zNgdBtyxaDLcQ0b6wmZSuuuxNsnm3eBLK5NhHQ9wyKtV0
RP0VAQ/tRm9X9rMDXW2Qq28e4asTOU9EpjXERjY0yRRKEIKHYm8eypJpKHtt
IcOGhRsv+ZCVzbJ+o79LscCmDbusTqRbdhoDf0DoHkzVYWVsv22/8sYrDcKq
GdoHSnbRP/C+eY2dPEg+kT9gJ9/VivVyZgvHF8E0cY3KbOvpFkqv0O5ZbQCT
KepDVLeLlYAUqyZOVJB7Cr5YVDaebKuSsGLZUhojhsijVmJhAUfJ9G5cfn6c
PfXYXvtLjIEULoVsu8GVUmVA/bVQlzJu8kpodggSFGU39EHRHhzcyZIXmYuh
n+LwIfYWd+g7k6elON9Iolj56xIKvdqDMVOdq/YPPcoZjdhjcyExRLiscnDU
Iz+rBs+zc9Cb3pdNpbQXLqXFSn385WMG1VzYlIjUN7QMYmln1qxieCDhMxLX
Ara5AM8n+HsySH0I71mXWjwpCubKkZXyRDx/xpwxX5du

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqezV6FWcEwJeTZDcyYnVGDciAOVFOnSqChfLH7SZ4C6xFfR4KlxAhBfWEelxggifArr3fE5OE+b3UMdYy5Ca1Y8pNMKh+RJ6Dp9WY60qtzSDYlopX9AkkZEJgrBK6BoPyn3W/vzJMf4hW6LDOuQnZeoOYTJKSTbXIzyL9t3MEFlzXgwo/+iaAokVhSCA2txkIXEgqOL2lkcSTp4wC0qjUhGwzxRkU5qQpGuyuBDcyQ4uQqR1uYfHZ8tUqFS4YJ881jZrHYmVqItzrmGkxFU/whstSHN6xVJh+iWIy0bL19unbF2iJu5hSSDUGRznWCvAGm/6ul1+vcEODhsvgCivUjfjXNYKhdbyIH3bKF86g0poupZz0NgqiHf2m36/afEd9UEkmJEcnZjoHBUH7DryrgI3T2v+O0VsCM0KSRyi5FcMrANWNFIycKA42s6f1Zif16nvqgWXb/fU+tK5RndDgtDkmnXrAvyte6fZCwLCYS2kFJa3m+8BtgtuOzT2UzydoIBpdpfWKBuF9kiGIveJpNZv4U600hxtVJDuEUI7/1aEmxZaTz5Q3Y3wzIfmRep4X3JAR5pPW/HlheEG0GJNnhSYdW5IX4hKFm7Ed5OWKkWRlZXGdhtHmEYDebXueHtxsntxMf30oaeDkIUGhG7TETWbjRTp+0MIoyLoq6YVgarkotcoSoibBu3DaLAj4H/5GsTbTM/Y4ru64BJw+kjHdh/ns4qwoOaez4nkNHO/LIPE1efb7PA47H5rfhNmJC1UKF5B766o7bF4mvY62+3z7qo"
`endif