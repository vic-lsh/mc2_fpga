// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N+lY3nC157Z6PC7glmdoR9l+97tfsTDlJIs5Pxqqx7NisePtuQG7o9HKGM4s
7MzvLQBoQMR26BArAz8TAqwemPqnee+wQqIm9rrOctWqns9zZ9/L7NOM52/e
7IuWXgMyNPwuFgQnrYsiccJInUHXNZaK06wP6Pewz9QF7N+10XBI2DGe9G/R
faouW9tYP0wxL0W+k5BMOWWwnxsGC5j3tOkbeUJh4rcqm+S7RwlhfHByWZk+
7CYcOBAbvYMNDJoPCh1FzA23DYWUCBhdhIG92TLw/QrSWy9nUaC+yOU6sceN
6D8cs8lUgqZDtgF/wYjdi9Pk2u1NsHGOH2gLnqYJDQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LVz5vWwsfuFBX30rcyTtOKAluOUzYbv6GhClo4LPDFXpyXjuluLsZAbZCm3r
+TTGdR4mmBM2WBjI6YQTTRceL0xRlpJdZrQiUB1XprnlUHXB4kzTmXaawO7A
z9xZj2XIS/9v1cb3DBShqyTZWICLWWybEr8yxgtuuuheCZA4B4tKJzrEBa/H
huH9yqMoeE/u+d3B7ZI/c1mll1uVMmoftAqExShwGsGXq9x83mod0WsUeTf3
VlwTdSLkGFmApTJO1JHLX9qBHmD5brZ+IS8I222EM0hnNFRuxlLnjoe5HQ2/
qiv/mb29a2qQKTqDMLKr3XuYTwhqAPhrL5bwZwHXKw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E0sUg+rzPwwim//0VQ+yjajs07zrj9IAQtYSqENjR/azTHM8p5ATVjDfmpz8
n4yDpnNEQme0qjAI+WYTviGzNX2Wt9Jvpbcn2efkX6O/SVuTTmGnh0Vu4jJK
JBbbEiFHSkcPtSBpwYD59jT19TbGTX8wW5HUiYHL0pVAW79KKcEOldH8hMJZ
9bfQk+Sxaz22UCp8+FLTRg1q/1224i7+8FK5fztndU0j7B991W6kDkDp79pE
VaFCEPQ0RJ9mi/HbvyZRSN9XG7tt5XDV4lBlSvH+coLyKpInNSHIuo8aeC7h
ZYgYZEMKgz5zXjd2KDmrs4XwsQY4tswKqTQVipoFTw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m2/Ps5rnIM36j64KzDUh8qNvt8F9bnsQlFK+Oz9lRme4P13xuq9JJmaxM10N
5EbLyRvvHG8mmoDc4NPQ7fmxzWbIGijEsW+87iCxQBWfE2GGpl+yGs+6MS59
FAXMfQR3GqWtMVujbVj/0QBdo1vadob2+WrCF7RPnvDIcPPWn5vlR5pcm9Gb
BYOkDYBiFja9GbDhtUzFGsIuV0avWPf8LUHRu8aSLuYNu7ViP+7HLQ2GFqMZ
/zXEtqkIyWeUuK0eVJqUQ0oRSYrWYgc/vHM8XcYhE3HCiOzar7DqYPdZ+iGF
MR1N6H57jBh1p2wsTbjd4teW9WnUMqdCbEvTj8Uw1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r0pr+2MMoe/+M2/PClLKz20Y23N9C8LFuHl09pvuen6/WdwFvqQ0I8aDrrkf
MWEEsoxfFyJEVlF9dR8H/p/7r3393EJjUM0okd5msISFymcBZJhGR4HzITa6
IcpDxwlgm8gohU2i/HnDix6Hd2kRBK8qSxmiNT0gXADb9e4gKzA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UjUS2pKjFapUlWnw6O2jNB7N/qHL1E3s67MAQjJuZ+cZ8yRMz4D6Ohctfz2e
pHbhWWgDmL5Ah+aDGFUlSpC/+XATwsWyrxWZWnmo31cHFo1enqmoCbK789x1
K1H3ZY3PB4VzzxrJsGfsz9tfjtqaiD01zHblnQWK0O8OXVQ+Q7nRp3FaHhNm
rX6otWp6woYzUBIUJIeNrFgmTkrd//7eG7Df8kdFbIs0TAg186eT5+EPgI1U
4lw7zUhcbCWwuuC7JCaG0MNsJlEp4ALN5AtaxTjlcoDoRTrzEl78megyZO5E
ZC0y1NHF5dNS+/nyvHmgPVM1j6C9ANuE4Ke5A6yLvPHmTMmR8zquHtuvgRMc
zr8E98Q0GS0XNaMY+JNmp7/l/PLPc7tZA7EZNODqmjFLtojZsQ0Ys5fgEXyU
mXVfGuMyynpHo2Yx8y4pmxEFqm6Yqi/HGJd7tJHZvbo1BUfN8ixyt4EiVnDA
cukAzNgvLGy/fTIJQsG0gJdexakYj8bW


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i30ZkgmYElklHoIxk/NoWOHWz5WNdjZQTk6Eos8f8VfsZwIX6FbS9Ifhs04d
WIuR8JM1/nQMvnY29U2BdLnjq0H2vl3Ebwgsgv39bT9dBL1g4b9yNjq/fXvV
rDm8CQfsPOLqumoydQxZ85zTgdhz/8j7sgGdUMKVUNUAVXArZ6Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kRdQM2GtvgTFAi+nOtY6w43DvKlsIjJOyDLvXq8OsDRQB3fIE5rqA4zn7Njs
KY1ymLz7r0LHxFUKFsDQBi9y9NBs1QfW/2faIgtNa5CFAWWUifgWvYOTTAdj
3TOEpnFnEJfLVtIXG/IwfQBMEID2Kkwn4PClBbUofy2/KMnhTMs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1408)
`pragma protect data_block
XGl/lBCGni7xUSGQXFtlB7MTvfTRDUuv3fzuK1IIVgevSnj6Y3UJFEbZE/uZ
bIDOQUS6+6gYHXhDKTygxe/98IxoMMr7IOK7nyYYIKlHvn44K+Q7BhLNyyHe
zlpUgW7en0YRduOBv+W8OJ1Oe9OPV1wqb5CWgBTj8wVfeyhpXPZEKxb2uSE4
iayJVigr0vrB7XNNetlVoGuYU9hHM145nYBe4Z2qZ7Z67cSDaY4wjaK591j4
mbWlN0bRLHShoeHRgDV/jm9EdgBqcH4Iy8tfzirHgDGoPy1pQ1hvkMqhjs/2
2/3VzvEAQlFV4M+P4kf93tKgj5A0lVXHf7xz+41AfCkbVCP/6HbQUTM3cYy/
Yk1N/j20HPm4XRCws7eMHJR1wRXwbkDv7vh7jXk228aml42n0kK0U4hZAzOj
8MssAtiZY/KHT0gnrqoiaBh+FHNL9Jz/cd75wvvqC6iltFxyzY+s1FeOFsnG
2nU0n/TjXh/d4LpHm+Lf8/QS/idA5jr6bLbCEZX4o+SyActIJnVFcepY4x+B
iks+l7xQdxOucI2fpFxtxQkZ03KHna8vgCW4K6O4UYUbjhRbVFHDWq8YjajH
4UnWNk7FOtryO/NiF9xfIVmz//XyXHUscEU9ULPpOB+XRCtLIlSQ6G4QALMQ
OJGMfdPzY2/rVs+3dJoftVG8NxBeykvlQ6qu5lKYvTqJpDQX3Uq58kn0BC62
fB+q+9si0nsCZqbxHMvijYzkshmpK6kbCEgdmtvMQwE6aJ9Zxdj74EsZ1IbB
UMD86MQ720hh9CQt/GwqdFfRvNy/Z90OCXqAy1xmOx6cimHaFm44EdtnQs9j
mwxSSOJLC3QvCggBrYiK4+qZPI1i8sMaoX9Yfj9Q/DnYkm3N02P5mUdfOdcD
8B28DlHtPfpsrCn+xk7mP58VlYhxNyPWm3ZzC/5lG2ofWpJ/YJue9Q5j/Fiv
W8dVFGRw8/lSL6KNN6SnTIgwFF/bDLfwR2e25VAYV4gVHOrqS0sAhXjXJxma
qnbHSevum5ObBLyOowuHm2e1T43boRnmVDjj0puY1rMhaKNJC3NEWsLdIznL
Ik5KsLuIF0Mlg/TWqYHBT3kDN6y8SqYc3qy8yzUZFfVfp5i96dAmNpFQaLV6
7hvUSD1YwFppZGHZKKbgE/T58R4FqQVCskKgnpksHAH/oK9HF7IdrGGQUHet
mzzEl5XcluorpxSRCHFdTNo5iicer1RlmkiWZtOzzOh/1u3T2bpBQWXL/P/z
a+HMt+kXFeFmrfF/5l8W5eWD+Xyxo7lxmi4h2UUmyF1AzXT/8KB7WdGkc2Gt
RXUnHkTs70j2DyC5uF6VYyDCkly1dPHbqlIDhXgoe+zGb2Vtky/q9ri4YvXg
IrfAfDoFFtkxWaWVOXezIbMyMW2B1msxQfLVy1YJEjnOgLzI5glyzFP4JlI2
k6ODuOMJQwuJpLWiPZ8syjYD4WT2H/7TLdjLYrZ2t/i1C/wL1gttIXalYagI
Us/vlvcS+Uj0flfjclCAeKtgXGDXTB/8SF72F14Acn0mVBOhZxP3uq2Ti4ZF
bO1aPEHHoN9OrVpUzO80enIgcB3SnXG5qsixCecY07WPOGGvecPLFn5WOUf5
A1Xjh54W6la2skfoeN60Dxyg0oZYSpS4jtqVvkNz2lEFW2nRtQ0nqiqq/atj
tUNxtepkpZLUehP9K7GdQCy9lmYyxc1IVe6SDP0lWpikrximk0coGDUSRItC
cEAfVyZZ0g763koty7EYC3pfFpAzRSmmV2Dqimgzs8FqK1z6d2mDsCrTFqdl
K03j+zMIeQ5Bqwc3Bxtv3Fa5HM/ZUsQWyA1NNLsK+Uj6Vkf+CC3ZH63C4XdA
VRffWI2DxguN1zyqmA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyIjk1wSJgTLdLbnYZqODRGurd0anyI9waAIbUL3b/OeDbUBYaBxqzCJsFTUmpZY6556jqs0CF7gTEDfi4Y71+Apt9kIozUHhesk4MZXLZEHQnNoAiwDBfXLo5IcHA2grxqQMqOWGqpqDpZTkCqFL3phrBSt4e+Wnf2X6yo7ViHNmOQ0Q1Q/pRLu0XDsTB5/KbYCSSJpD4MDwD8MPW+LEDVCGThaHAFsba1IF7YEPtF4ydXsYkH0RrTGm3ufunvc4TBziAc7Qxu7HlDak1qBCzSGtoC9VyM3/bPazLNupgfsASz3S9k3LQVVTwRyq1OU/kRojguT0P7kMNLV+Adz29ihXvxW9uyoVwN4vRANm3VkkTSINXDkDO73PMNQN7drNrGPbjAZi2HjbktUI5eefBFSKokFNNcS4WiHDxWhrhgjkdbNs22FUK3awi0lo/Yo3BcgSB/OUOaf2tT2sD50ZX6ZZ46YGmC2GMypeOAWDbz0244Ba3XKUGEnwAMWEOGFP3wWNs6CCq49WOfesr7hQzCPeDUOXqMf3Cvj48v/hMDbXOGcj7pjkBsmDQo2bizsl3+3AEi9fpndKnMskb17P4BeW1xJALoul9BLTtJ2CrU8ruYNTkSynVvuEqaqcQGXemigW3TKKJHLUxW14VrBmmI1VHMwTPDnS4QAY1qdWfp1Xl2YilVQiorz8lM6cWIEBeYmf6ijIkia+KcU7W78YmC2Yu8t8ACy5x8gYc/2D/MxDHSrTgUOxDLHlymCn0lMktQBG1LBOMtB8XkW8Sso38w6"
`endif