// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dX0X7jQNq0z2/r6orEF6QhcnJ1dmwGNHwPSPZg8Gwu3gA7F+OzE8Zg5RUbc3
gsczDnsSmL3xmQJU5zuIyLICaQTszzuHuJE+kiLEemB72PGB1lKcPYthrBGK
GHFqeOa5Z8e3CkfLu8R7saoLW/d7ut3loW9gmDCbCj/Fu3CDXWmZKPDXWpIi
wmyLz+6sj7jOckTp5u5wIE1jIkqyyPSlcnefHg+GRyhDNd6AnXXh7Qnj4/ma
KHNCqdSVFK+Rv+uuvXj0+JxkX2huOXuiXxmBrKIBCubyxCoM5l2URrD+wsd2
DZzT4lZq6CC9C7ADwWuHEd6GYqY1ifZWgygHxatndA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EzqnX+org0URf0PFotUaSG1Yvdmj8LtXKVBAeUqmGFWdsDflInDIvIZKQJzJ
1t4Vyx37GY0ms/jQOUnNQQKsLYLvtp6lyTaJcSdmXCzrsCQnXRydX1q7i04o
IgO+dJqvKMmt49KArViUqXxFNDtMr8spdfsFh2z07OTfhsfJVzvzSEuDlALO
YOJIoyvwU1hvIOKfv9/X2UJAPsPeL0ZolTADo3Sy/KIIvNnHA2CQ2FCCYAKb
X7ADsRKzh/Mv0i2KnrpP9H7777SykpZB2KdvMxUNTBrqjSOuZ3NZjbrjtKHu
+7h1q6+BeZGHJ+h6QIn4Bs7HK5xsbo0ZAgwUhpaXBA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VKhY2uOsSg652lvg3tocqE1tVdATt8+Vt4gyh4x0/+A8P0pYKnMFzT+l3vaH
viy9/zSk0eSmbHvAu1qRn/bLGYORaI8PexCZi9xuf/kmrEq6M6IrxFKWtv4/
Q/4biMNQKfikrwTslSnauNMoCWIMKLjTRU2agK6RTB0Aujkb+aHImBR4tAyo
EYCZ/GqhlBEArfgiEFX8BAotIv8GdC+Di0USJ4t2DvFkJErlfA8xcDZsvo//
KN86pHq6Iy3a7SoJb3SlgdsOctRuodW2WY7xbhnHzoaP1rJGWsn/SlNqMERx
j6iGWWqh16G8KzrzFEirRlo0L1VRG50BWa+Q+Iu1kw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YzB1NkqKgiGqcoArWlUoijUHszVL9Bdspy5UmuBrRV5l4tg+FyQS7mxUsw+6
UwqQgK1jaUJ16eeg+Dx8PHvbcTnnFezlwQgsbI7lAiMuF2Duk0bcOlz6OkHm
QUc0XkS5LzLvHQJfrGDETxxffrf0jm/5E2+fZkltfS0V5RMgowEGpLQcmOvU
VczVMlRHfYF7W9/R7Mz2xnJ5EYiCQr13v9uYICW4RjOQUdXd7sWNvXJP2vHk
u2XLpUxNAwoYO/1noarpwPS1FvLqrLY2u7i7ImmxwEeUK+On/wIRbauOE4qv
T/6ENa/F+pbMjKHE4c37Wpaqtc+EEE1IrTOXzcP8Zg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iJoWmbXawmIUy3kBPmEIOvfVSZPLCY/CbbriGtGLBrC7OiTMcTvsZ5gEUfBx
OMAnhPGhHVmfMgREwzsTUCAi84i/2oxU8rimSC2ITkBqigQaXLH0hSs7KWSq
IUusO0enbnocV3QzfNromwVzmMHGSdqZSJkV4UG9RDK87rpqSAM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
D/Vc0ip9Sq8eZw0b1IEPgjL1paggxBwSlJB7+aQeOIlZosmlJiZl8WE7hoVo
7TXJiFpxbcxESYEGWZdvICiEMoDCL6aqLLYrub5+ICmH7cDryovUdXRFVphT
qESR1J8bJ964+K+IVOHwoCfC4paDQRumh+h8dLDBWO9sEeF0lm2zM8iyNz7D
xgCKyafA1kwnB9fpd+v8sTpEal1N3N5JwOFuL3SW3yP+LVdI6pWi26BSXD7W
+eVrdd3sKzthgN07DhHakYWKxo+vD85BxBrxrk26BcFOntVWT20g7F8gpBH8
ZOW1qyCNAJqR3gl1AG+y3UULtGRGvJXOrZtLUuaCUmjtBf3CKo6BkuMix/fy
xqTvlPstCzH++zUoEMqQauixB6x1XMoyZspgk94QIfdiS/yJ6XrBXZiBGnew
FSxSPlLwqxMIRt072gxwaVMMSARJk9FLa+mbn0FK2xlPXvGMNp5iv/bWTwYq
19lgk3p6F/+mZtJi2j1Yz+SUEzR5Ar2i


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H9WShb8cTFQ/co8dYlFPkOM51ygppHomfdAKfv/I2LD4wrixVEfBC7ZX3nK+
89c4+fBLceodvv0AnHYpzYyT9i8M6QnsUrdNoJEgHju6be4hw6pJAactuP4k
0FYt/70xrJk6I6iM3py5aXF+Q1LX04DINKhk2naJhipPqeVCNIs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sY8xiuVZDcw9h0Kj5upz0v2VvHJRUG8g8icMF/0vO92rvYV4y1bzQ/0fmbCH
rZE3mG1kVV76B0Q1wJYi5kwbzhEP7wE0+vICPnDnXQOlV8UMEQ6cJgXNECoH
w/krr3AbPTOnn/4WrQephA/V8IoyvFNYHB+kXJ0Yqc4D1gGUIUE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10512)
`pragma protect data_block
bAdxn3pUCnP79UfFdzdF38Kom+zKpPGkJr3pNunubfOnHxYW9gClwn3kQzHA
WyEARFG//1B7lPBRLSeOoxR2GvP5+z7soJjXgdRY5D+nmLeybWXxHpER6qhk
byEyO2RxQWFKaEafM5w9mA0RtIiZmcqvCOFM1N9Vkmueu9zyEE416VhqFxCN
0d2EeIRkiiEs9Ru1IC9zYDjSl4O7untAiGj15J1cbRgD8crbBELBWOkvzGnU
ynL/6b6t4GycvKwoYlcRsOYCwGzVGtzYhWnjWr+Ms69NxdszF6d7YHyM6b6a
pYf91D76zDNcoA6c6UyEbmGYvu2jFJGAkA2ncgtHQ6L42sBrd/9Wtt+Hx+ho
jKngLlslwtLfgd93D4ut6FmGkMdYE+fzmx/RSML5IfK9lp+EFKE+t9iCc9hF
nRVLeMuNVpM3VAg+Yj7LJa816/VLP1+HxhR25VbnGgU9WYX8PD4FxSt9hHo7
kgup7364567S/O3pDqRsYCobuMbbesKVEEbwgMrTegbjf/EttPKAC/6wFD3t
sCeaBFtX8nzDoMgJgEcLRqsUwuUzMb98eVw0nrei+6aP6atzkayzI8Rx2C9c
+iwnzSCCOOOdyBXOSnRrGJXxHdCGC3jS8kSRldHZkU8NeRWcTuxUi4nM4Tg3
ciVgYS8aUWeoLxuChOhGB2Sk9BMqU5XxUo2ksYYUeGKt6S9FW5NcDOXpmEN/
3DxRvTk8KT0qzTjMysaO7p5lAphejGoh09EPtECLwlyh3k09VxXFe5dToTG8
n1+OFz8ae3SlSQmeOPwSUmKzmXTgSxlgrDcwDnjJtuzNpi0c542swhEAgYwT
A2cXpKn/I8s2q1kJL13oGdGAWT+ubIg5k5bYpnZLICnKG4wzvqbhVqMwPC8B
bWD2LM3fX9kCi7/OBC3mfn9v5lAdEFpzEc5GfVAKOTWH5pTrzmc81TmsCROc
SMgjif/pgKQVNli4wMbK2B+As34o1nzt8IUfAII4pCvBDrMI4cb5Xcmz+v41
ZVbV2ExmWXse473x7UEQos/UX9h9aARLbMr4nrWfLSuIrwOTQBFm0HfKsoq3
LXN4PHX4MSj1S1US4rRBJP4COrspFrNvuQ4SuKfxZLx8Just/4426fQHlcuy
vkRvmCgDmK6UpbplubiXvFjsaOLxazfggrrbPI0BK4YqdXTrS2VZi8bFt61O
zacw6GufBFQ7VxHM4Dhase/qSz1CLk5VJ+vTVnFIebQksmTM6h6nDPPXpsmn
PuHbz8U66jw60v4uRgt4S4w+BYXRdIMjAnkV1e7AWLvKjDpO9Bx5VmUggV5l
SmBevG6RyUC6ni2lDIIDCjxpEx91m7GD/oDMTqcGEPITuiV0MWatxQo1Eicm
wwMCoWbtBamXLgL6K2weug/PldtGPAmsidnIkTs27MersKczg9TVaH/Ec58A
DBMftwXIh60k+G5z/E+sGWGJQteC3HIatAg98v6GxxhVZ9X/OpQLvPGHKC6K
W2BmToBDcQXKw8nSPz5PfLGRJ9qJWSFGh54NmQRSvFk10dzipQwm1UbxTTtG
arODPzIjKspjAmrSZHZ7J4QwDEAFUHz8eegZ4mOIKBkea5oaATHJ5DYvcJJV
YvK9PgdRATyWSWRe77XQuu6nKFluWLYjnLn1wedF9AAigSDXXCX2DvocqMvC
jHfcSu9G3j130fg5RwIW1IEBRl8eQhLs3BKH/IzVbw0jVqVrArzSS/j3K4OT
L6vS0cEW6igkmMy2RQEBJoOpCEcc6r02eG1+XLVnNQxZuBJoPRNHmVb1+L78
HT7JXV3PsBuix1FYKjszAwU9kEk+KHJw1K9/nq7vWcCKA9cwVfP9WmAoceX4
ROZ5gyXwU99Y75yUPkAC0ymVzNrYDfmtdt409ChATd+Ub6Y4aAVAUG0Qfw2r
rCJkZrV9VGRx74LZRqegupII7vckZPhNmPILJ8KAo2TnF/1apIe85Q8CnnUr
iy0lg9T81b42ilBE0JvvaibkSKA7EhU9uQzLSfskKtP135lbRTtTtOiXYOs0
ds93FnGvWZ2SpxkLB0jPpPkRkT6LrOIGq6umpi1b/wN76QP4unw9tGYoLVNY
h66Zv4AAtFCdEuFXnGF0wW7MANLprS6I4CGVSimhjp8OGKJJN/C33twTHnLa
Cn4wcnwxcTLIQkXhVVLnGBlC51c25rkY2VxLzJO7ejR7j/2s0IrRJU8aUnom
2SdVkaE4kzEf/GWAEoyHcDunfgxrTCUbGk4gVEQOPPN3ixmDO9RMlPE3h7L7
R76WCCdfbQ9wtyCveL4oNJ3HVVwu7fa35IFw2IP+DkNRkcGJg/+u6jjWuX/A
SNJ9ZgyfCGnXj4w7POZ1J9UVNy0MFgVw0I39LVfmkW5EsatOIesqqH5wgIgH
Danaexk5hzHCBkKGqM2S11NHRw4slkbuqsDUm5f56PZLHH4AW0CFEMJKrzRK
RL7WRvrP0DuGOxeRD7zxTlIHePl6jzwSHuXo9f/cTMPG8TAWCJYteywlGZpg
+3GaVA//RjE9dR3zI4Ii7Gw65SkSOziNXj45J3IV/GfB0XQgAFkKVxH2D0LA
Q7u357uvCjWbOenj5R+M8DUBmuFHiKZhPptNSzNXF2iuS+Rbh5zrEP8zfaBH
ng3fSpVuPxRTv+aB6qkF/0vf+eZM0tydBfZT8yxQkqwrIDiys/PsNj2Tf51A
qbPLDbkkzmrwQvpVu6uaiUebIdif8NL+8ni8hmM3619PUHXBIinDqErNugn7
35Zh1XOgvOtYrOh1VBE7L7g4tpRJY1nJS2zkwRPUcDJlIc6qPCH6T49A27Mz
tw3t3VCZZ3WD2DWSnxjltDlstiJF1uq2EX61c4P2wUzIdNkYta8D5Kh4i4iF
1NvWjhUntptIatFNAcjfVa4eTTaOqeKYpKpByvgCPnOue83s3yXRGofYYB4I
2SzFR4mS+w7aWQcULu6VVLlTtzKhY7RsnNk76Gt12aMnGIm2TTwRcuB96nWx
xlo+aip8ekQZ3uoXh8NStqMVHOnHOI1bhGJYCb4L+U+m9/Izv1pXmiWLro++
x5WvUy3RCwOoiuON/BW0TwwdG9MZIYAZ6V9iq7Dho7RpaFyp2XcX5YmgdX5j
08MMTFSgkmsgIyc8DRcVEuR6sUox+YMl0nGYzoJsODfiKUBW9EPFJO3m6x3Z
7lI2qv1umMa/ModpDTfJG1l6ULd1GoSkzTf0TRP/O8pEwb1Y0Qo1e2Mtdqox
0nCF6uhzdkfVKCFMuWQLE9JLwWRHKb3ZHCoIvWI8LhNW3Om8+/329V37cvTz
kWtTD6qhZB2Za0QpAg1yTCj8XQ+0gwzcjMxbqjnuO8W9qPM5PCVXIZkuNXa8
1ArdkkHDGKtM4Nu7uQAF8ENOqUkg3GE+gaUIQXpwMFvOdBAQ06KtSRIWZTlO
hFf24MZlj3Uyl4uxLucveMi0Ux6Jz0RFz80os9oN9w7BvcNcd+kz0krzX0n7
moKIf4qHx8hl8ql7Bvlk2fkH5gEiovh6OEMIBliYvfdE3OBo4LiSwgUh+Fuv
grf3VptXsXLT10xyDbbr7STZRG1cav+rro2QT1Vmb2at4w6U/USdHhhT/6R4
2qYU6MdusKlT3nVpUCMNLHZjClPHqMRNL120kJyw346DAIBYsUfFyI771dXd
O/JXL3GrNukwYXbfm3Ygw5eIgE1LKkGXxnjMH8nx2XIl/TYRY54nDYkYaGsN
0KkjAPSCCnGZvuinMxMbpkDvhCwF1lWLXZkDw++rUKuwRINpoEmBL3aYZgbp
6xp+LCGndIsasRH4zAy1g4QzSyyoLjiPVxyyJIHgVAui9EFBSv4ybMBBl9pZ
VhwiieBBzC+jmiRswYLTaVKjL7kB351xhpMb35Wqu+1+N60nzkFI0H+tkaBU
o+MXg8WJbB2vboPKAx0QT3+aNQfs/6GexFHc7pw5ARhWAInPf0Ui7cmBwkpk
hcsNTomZUBjhUN9WuaLnNjJQnDNDq5B8S0kFKbYa73pMJVF63Fn+L5wY0/Li
p6gH3bxGMmzm97C84Ugm26MdhuV8aDb8sIaWZFzkylWWuXF/QpFE32eRyLuO
FihIKOm/7gAVCagM+ODYIpjl9M+Ltf0MTN+Wm4otHMo5da1XXS054hJXbNEz
IeLc0osO21SQYWBVLk1/C/yzPqd0Ddq23URg5FXm2xLrN7PxjeKAxCHfiGK5
IkHBnRyC2p0FBltrpJRHzChS+C5f+kYSqUQ/Ox6RVsOIogCwztQbU+F6UupU
gGRJOQDAsvXzYli/MqqD2RujjEx8KvL2nWmPBC7OenF7WOxTFCv9oRF5xeGk
IFsb6RY7FETlU5IOTGNVZ3HykZAnJKrCibJpltjcUNnNFUld+1yi3iTFfwvh
CvcFpVrtvX22wBm6jBLQ8s3w6hY9WHN5SDPoruBgyb9PQVChQNg6HgCmxr9m
uJTudx0/ARHbHhx7nZzlwx5aeF03Nd84IR3ghwKj9zsK46fCQ2zQlPJLesRj
YkGARzqwBm8Hl6JFK/l84yfAj3jmG2+dqfuYiWC3aAULsbf1saAff8AIX8im
t1ZJigCzT221COBWD2f0Je+ZZ+FK+wcibZ/hur9aweDBNKT6awlNgAAB/gWc
iTQX4/k0Ko8Uf9iWW1fgv7f7kBVFIb2er0W2UbqMJajyUOblLQ3+O6Xu2L3a
LI3xfjVKdRMsrOcPhp8uxQ554DEtL+QVar18u62rU0jTkr2Khz9oJnJeJ2CF
jfkfa7vGriasxBoSUwyuXV1hxZwV+31zRYBdlK0TkDgbBDm4bNQ3C8VzMWUI
6CLQr0z88Sz36HjvUNqkraBDCbZO1P3itxSpA+Zd2fHkRueiK85bX4cZn72/
FcJdMwt8TT0xnorz37v+4ccDsd3msFhsNrWc05l3MuHfA6QcqQBoOzo93szf
Uo8V7P8E4f/fRZiLeOVmumZy+u4SJO0vyKU51QmRyFAkrXQR85L6uB9yXQg4
fX8wz7VJdinugjuOeXxGc7qDPyCvrd9xKO4WhNZHkLUtL8DBDWtrQ+GY1qMS
aQnIf0qeBz2Xhz8eLEMxYaZobSAM97IHb1XM5FCLxfx9X/imf6LJpwLyDg3a
dKvY97fnHJSxFDbT6ax0V42+Eo9xSKKNlqU+aG1iGu7UJQbE5Z+lL09b0pMr
F6XT5k4uDH8UaPt7JDnKnJLi9E9gwjqHGfQXZLqYvqRDTcPKQej3w+ZTksuq
RbHzJenp24kV+B+DEqBAgMcJaShTa5YSAqeaNfyDdkbfZIcVAdVP5MzuId2y
/dR+PanqHG6snBAwMdG5gjZZ3+4Hq4n+ZTVO8mrUEsCwwdlxhybl7MsVmopT
Rj5joGIA/KRwbUGCceohqnxzuq7t9lj0fC4gRBveBSvclG2G+Gi6O/8hMdRz
EK19yp8dyKLnKgK3Bw0TSwdlw0WlQiW+tyV0N3SGnmxs0pt9Tz5zcWeSdcpH
7uYNPM1Bai3DQ0jIjJU3euJxdVYZCeFUnQiZrSCBU8UhmwtBd0mre08Athea
2XWxLl3BlfFR+Z4lR+3aRsQzxklow1J9ATqiKCOpwKHw8lJTETDooFMBAoMM
6S8A8bkYH8HiEBhFBTYENnmxIcQhCSGdfWPr70fe9P78brRHd6Xqy/sBVoo/
17rJfi9pdAKYacWsGsvwpyA8xNopUfiW3xZiKlC1gUdw4kDeQhs3dQvxkNFR
LAmjrkkNSccDmDhuNo9zpfkJ+moRSkdDims0vkoVP04evoENLkGcEWUg73nR
L1fp8rbjIKdPIpnibkT6tF82aAyqklOkA9rcmxRzF6n1MlGcY8AHlhJERJUK
Ti5xe7uBgj/Q53yXwR2y+fCISfwisovF+V0Cy3wtWdGnXFjsvY2LIp1CgWhu
320L1lFpHkCG9fHTrnBEJRy89f04ip+MRt+dhWzaI9jJDem6gxfvJcPqervO
b0cRrJ5krKphmjpMdLR3NI6nP2jdlR52Q00ZKjScdkbBXuKTaQe3unnvBnT3
4d1XX7fdWiy/9EdQceGnJvkhnu7r71bgkW5Sa4DmptzZOgnCrt16ipVS4fST
AhKM6jcqMYX3f07r9gFTpoXGuoMnSGRPex7/6Spfl72P6XqBDI99fn0oanC7
0fTG9g9VIflbjaIg4qIzFaXk4cHtgZ3Y1LS84VxCfcoiOELdd0+uoziOJj0z
DhPgV1fzW7DxHdFdTO7mj/u2ZRWD/KzIPhcei/iIBvqaOt3140itPEHAAj20
2HwI39we9YT2CngY8O2mGZugQRG85uoSUTom48lArEZ2ujdbbwqH6KD6U9bE
ouELEX21ZyDEf5A/NDv3LW88OWNp+KnncqbZXwAvwyeOA8hF2Q4pctG1LegQ
FcAthbhMO5AwJhD38oaX2n+cnd9MrGqZMe/QnMgRg6CVwFzkQWtYHnj49m+t
I55S9OWrU5WQeomlr1tpyDuzP7IkCWPFhuA/hUY1+6G0+FCqsOqqXR3kALY3
DZhP316oKP7QieSMa8WKCgUUNBZzRcK8puPXt6HQUyAPD3LZ3jVy+HY5g91L
xvahifRD/N7BdrJRxbQvRdqT0MqeQORigsHk9JFQVK4nwLjsoWwWRRCe/CiH
sf7t3q0voeE72XIunXUWSelkOjp7fpblIqJA3pOLH3FIqmTrPOdozquksDnR
9QNUPZJZ863En2LkpLL9Q+M9Vx1JDYKSHdz1bk3d2shPouBpBSpwwF8M9xPH
3PcR3vNKdg2alQ/21FIC/KL6lYWtAlyE98kZYhte5xBUeSxlk/KpCd/L8zF7
l2YIUk0dEaiN3kQJ0lOVw3YvnUpmbFEQYSYT/A8+wsLv5a7fBzECdGvgZbJy
FeIk7PEbTsxN7UWlmXbzNfbpNhu7ReJrBKqpBaHmAHBCcgB4yLCcW0a633nC
1vsRcX7rUonDpIZZToi8SBS97/+y2g3lBRutQ7Ogd3q/800zP02M3USLImHc
2wV8535Xgds3vGUgRtyHzk+01jbOMWnlWiheWDZ7igwb9QIdzlX9YejhkPd+
HfhlagBYZma68tM6CHE/UckU4jZy1hyPt9IuhICkkn6ChsUYphXREeFS/K+Z
q+nk0iBkK7GrYdXtxukSL4BUBH01amkpVkXdrefnWXOkVYcVTZYXpDklk6n1
sKeIavZWMUb+qaVab4aV/EMmrfu1SpV1I9Vm6n3pUnearcCAq2B117oTJqIW
HkT5FgiEY0yVAKv6kFqdtbthcKEhZKfW4oD+oq4Lp8A4hOzED+ZMzFWJNU/9
di9BoqvixK1x7W4m8tWeDMTgBpLlZI8Zo5LQZPpFQ5NFMPZHCknT3E3kg/Oh
pVjMHc54tUf/XJKADH6YI4XaQaRjELvdOpBJtSjv8uY+iGDxjTisXS4NL+Jz
ITB5WL3oiO2sayv2FG7fiEYUcDOZu6l71r5PV1JCBG6R3piSeHu64AGK8pkT
GrmIZeC42caqGU7vHN7tEUpuW43+hYv7GYJBkqoy/FHVN3BoisuIhH/knHU7
aAm0DCAZ8iQmvHpzudTFeeSkKkCRqAQki3cJDplS0HoE/Dgky7zoK992KQMt
N1X/hE45CadeHyiMCG3h/TZqq9P334LRTiNBS5OtcLv0EBdBqn9tl/s+Uyp/
arALFpGhkrHolDDaloUK8fvxZ06LEe4nBFEkm6DIp08RZMpIbIKLH5lJXfvc
YStWBB/4MQnh48k682timtKlaWtX09lSk3htzVWRGmp0iEa0g5UFt4e1hpOi
LcrQZoYUFSLzVJogtC7v8g1VWhEKqQVWpU+jBfRtTufplW5G/yyVJ5tHFQeV
+f6zJ69OONsP6TwNmuAZudJH1OnP94FgHpxawXfVPST4hDuGzkiaUDu56tcd
bVIMW8oa9I+GhoVvrV9ri7TS70VOJVhPZ2b7yGWZh9GhwAr3rkzLG6tkN3/h
fTZU9O1ZJAIpD+2HAVe1pxi5QT4SU12yIonpMnoBG2RinfAwqSOrKk9/wteR
J/tZnhqrOB46KymitXM5glsYbt5MqfjXc/BmPRdcei+jo7naW+mwgDUcA/K0
1uX4ZrrrQ0CBs878aOcga1EcNPLm87U0MRJV0ciyjVmEaoXDS54pAArraun0
pSw9T9bO6GQwpQrmpWVWjbIMsN0Jq2uz7woK+mLHai3m39xBwjqUfts2oXhL
csejZ5rYFKw5+sHxw6qnORqT8PkneXvg5sD/nlaBn0xJHa49sbZQ734WcvBp
FsiEgxl47uEJyvKsymzxdzTRyFCszPULGMl0WrE6COn7e8JQggz3rQGLA77r
DxOFsNhILWg1j31Oi9t0TcrBi0hIMzZdZYwiGqgeqj1MdSSp5El/Kql5xapw
tdQlytHAF5c6cc992sukRo/tRNq9nF5yK7Qf7xiZwufpbQAp2deVFVlX79uP
ZvBN5/ds+JRAVDM6gjzYDoIsKE3tOLOx39mD34iI9Sxxs3hqb2HU68E7OPMz
0K8hYDfVBf1vNVIWxChF71vTwT1O9r7nIlq261WKzmZ6dwTjW8D2ZXDkZ0N1
Nkc4d0kbxrEB0ECu+p8wxBygryHtPPN+UY586sWVSpdIGxa3oNa7i/o4QVwf
Lpzm/VSyfAjOxfRCu8ndydd0BQjzgOUtdsRHRxG3d1n/F424Q0aCsrf2ccWb
czFWb6oV+p2r1Dy6ieusS/b3Vop2V9Ie22r/eQe9GaahoRrGAtbhFcf4XOat
DwdFmu6VZEJ/lcRwMOrcKrvBVOHJNLHIz7vABjdB4L/kkqrPH68duTCp0E2Q
j3kyiZQ+GZxZcM2sSWJSZE0PmJacFdU0/SFC65uFCN3wT88Vxu0KYPejVYs8
lV4jrCm7fLEcu24sLd/TMrVK08aftfZ9qVGQe94lTeU0wdVyx/wd7SIrS7iF
Tjsu/uobQwIwx+BGCBNoM3ClwVdr/0wWsj5kSSSclSWCNz5mueTYrHwoAtWQ
PO5Q/lNSYALfMGwlKAvuRqrUnjfSW0fpQr9xXYfVd48j1N7dsJot5C8hzCfN
FbUk6CUs6zJkoQVi2p2nAAR0/AOUkERVY+APesGUNx0Zf+hMrtHbrxMTD4XH
oZc6Qor4MPXRldmZ0EeMAeBWfR6aLBQBHVd62h+5Joph7OtT8j0wU8Wq3jWm
zc6ucNDqec5nLsQHDSYbUtlu0wZC++4yRQzi8muLHHavDMrKvmIBtrfcCLsC
EhU4fBQrtBoQuyKTqKRs4wh6J9y9m1auPn32sZPieCVM65dz3B2vdTvpt86U
nLBKgnMykzZGkaFEK0x3fcbjtiQ8/6by9hWyYoWN5zSpMvAQNeSurO4qofze
rJCsoIZKB02VP/wHD25nKPu8tn+gnRyJtcbEGuwlQ5K/TNCAoQNXSfBZODJE
duCJknCDym26r2dteG3GP5dYkHzY7uwaiPXgyyUf3qk23Yk/96gL8CGoJVAF
ZXxmGTYfGfZqhAoBH5esc7CJFU4n+nZP7wasm9OLGG1zaifKUdassk9x04IL
kcvwnjjvhoXVWIJqnrP70tPBUL6b8uJiT5mQV24PiPbFkMjqmdTlFv23xt12
dI6W3ZQSKPYi4MOhOfK4Npolc1bYI44zh/qZlUk2JCmbEKIK8D8V4W4tK1NT
jYyPgfvIAqi+4fxSJH2mLA91hVbVleQ0yIo9a0okiV6IlYjYMQAriFsJ0l6d
vaccX1QH1wBgwBlInIQiSyHY3S8VvXvuWYwTEOSi/MUAEVlPdA7NHHgeZi23
RQERQ0k/iqpwdpICq4EcZZ5V8795MYRDJriIKul23SMdUZV7M9WMYV7wUJrX
TYcZCivNq8lyYHJEihzR//+2on02ltq7pv/WmRsx5EWyRpI9B66Kljx5Xcz/
246GZoOAMkx33C595lGlNXjghY5SCUNhX43p7c1vtOnKP3knqpZosKE9XD4W
OHZKpBLg2MFhC4gUqBV22rRTfRlBNCqx6ARUEj5FkFGAEKjHxD0qSXbDupcz
qBrr0bXHFhQjR73z/t9zj+ibfjkvv8nEMk9Jy1EPPUxSWdOf+/9Oba3yfLxm
bRWUlSqca4Ncjb6WRispMtjkC/Lzw8p0/wruwBvMdNr4bR5fuj9Of5ux3NRO
xhgsDs/bq5pNnfYgVQQjETyUIqpr38RyALr9EK/NN1fuBTKiSnUlxL/C0Rkv
OMG7WByjcPAz9PY+N2i+YtISQWDutvKga0dCj7lTilesiy2e8Qyc4Tkj9tGd
cXxsy0P05eFkZhisvEZlbSZvOTwdBPWTh65CDzXjArpCnIk/EymrlRrvAKRJ
hR0FptN7AH1+HByRSR4gtphLxAE5DlQXA+i5LaMTtLFlBhKYi/AWpsfRa3Fb
to04eWXCb3jBwMjYkhAHc+iPQsp3UUtU1MxMi7A4DhoR4LKE7d/zO+paqXwg
BML6yofy9NEl7TLeRdOp1J+vaemhITCA397+7B2hPNLsDrXy6BIewF/wYumQ
2SVTpghkiMVIY7CXgzFlbfIH/So5s706rJJL449eTefT1Ojl09KXaDEhkSpd
fG1y2FRNETQOnzZxUJ/ocxi6johO6ZVci7/G5p1kwWEtpdFqXCqKFEvg4eqQ
qJrpTulWhN767HntAmJfYO4SffTQZ/8kHR/QA3Z5gt1pl8ojN0T1T8lfLhPi
LCMXcW1OHJzbLbYyQQdV9pzEjW6sBK0KPOoG7ILB9AZ0svwMGFmQAutFC9+h
K0YoFqjPMV2yPSUifUDjiYND0uXbgX5hJssIvY8SV99V5wb9lLXhkOao8fyL
6J6B5XjX12D+pOg7KHGVNJJf32IqCJ7MA+tjbeV2HfCQ2GJJTvO3Q4lXQDhR
7Nj2ZeuPp8nJsqc5DxjkgRHiCjpksCXqOEeB827qoodbmbyE4OYfy8uTWK43
PgohjcBWmk4A3H6J36UsoonWFuq0CqW0BK7FIAr74MieazwvO+jE6JmD18z3
LKAkVTVWeRRDDkPMzY8mhWQCtMQ+zaO4CsrBF2hlMXj3EUTetnHab44XcIF/
sJ8+flyfVUc3i9u+7CF/iviWJJ2lMUO0eD/3fDGNP26rc95wzHJ4lN5w5b6g
yR5Zw2ditS7NAY0bb33YQKdGvCLtSTWxUL9lRpqngQ6BMVtGj4M95HjPr4dA
RuNDUTYu9hsGZWcLCiO6yHYy+iH92M+Un+rqXfdIqzWB0nqMqn2/i8//CjM6
58RKRvxnlxQcPszOg+q99aE0SWXCxU1aygULuzWG43YIu0N9aKd3aarhbbJe
wFBtvpL9h7dcMAlVXOyeB6jD3SB6NAVAxgeAgEUBVyQ95AMupMR1IizISxHh
fgXKfOsN33g66GgefSaD5lUshvxpYPyAxcHKCPoHsxdZDDenvxJHm4j93DWE
My18P0TCgcBOF6mXbrVOAdiaED/h3C2JADkH3LyqHx0RsKyzkqR2ZQusiNFl
Jmzd18o2GOpofSy5Lb4TkWGROhmj6AzuXWfgKJyMCCAayctdvG91tUYTVHtf
n5KMSojFdrL2H6KWRi6pDIQAR1kwXPQn7D/7irWSKwAox+R8sh+XMnTuw7hf
yBs/vWk/bTQEdJLIag8rXdy6oZlACFTuuKdf+jQvbbl9OrPD5MKXs8sRtCvK
lDul8uv8tNMlfE8JoZg9OOECeRHGoaSyEwl44D3BR5saWq5IiTuEtbgnJGAc
E6XP9yw7g7p2wEEEY7r4wuc66RYF4OiyqSEbtEzaGRXgedo/0x/xqqNHzn6d
9rg6wyzst7jddYgFNPyA1jX/zcjTZw+1tOyzWpD/k0tPEHRbb8SAQIMhgneC
ortoraSt6aQ8nwDIWE/TBsK1DxpQX+DPas5OTdIA3ytK2Hqz/NdD4ufx2bSv
CCh7Ogcu3ui9egcVhE4GAJXCnFkcuSgSBjteKv9w5fL492B6dxPg8cyH5+Bl
VIHeznk6yMaiNGx/kSYKwNf/3QkHJc98X7P8AY1EymyEOSr75Zznsub49v3u
miUUUsSy6feWPaFtQERlRlltHcfjABNuMBE2SRHqVTxHavCkcQv6pavR9NRJ
FkJdwU9kZ5UoeJ6wu5OiiyFt1Lh2FMpt0aas2QXzPN9Jx7cSin5kOwNqt05i
G29kvz+pAxQkE8V2e7wt4uleIAByuGnlDOXX3M5pUDk/Ji/C6wi5XpscE/hQ
HtU/yhoQW/RrMpTtm0y6Dsrax9UcvSHtRcQnVliGolquohrghudoWZ7p/hhP
fAVV39xILkGmXIIq1soeHOBNKBR9/VCTIJue4nxmb/7t4t5oN1Zw6aYyxtuy
3BPYiw74Ix72UzatNPnAkouoZXY7nAiwNqiQiIUs6TVCCQBWH1KOC9it2r8S
p4Veqgwr7nfoIwrZfkc2vKUptkpEIs/crcZR78FrI5oez0H+5skaNw7VhrYx
6Um9VqeySdzzHe+UzF5nJbCgH4/hgjPU5/6Xef3044t8kTVcspvmqoaYlLVW
PVXZv2NpW9ELyaL/z0E8lzX0HQsll0vzWaGU8xKGjOFil41596OjBUxtfbPu
oXFlIw1Cpkpbc9tN2OAG9fDN+S72ADm/wnqMvqKX3XgSEzG3N/RTFgunCVKw
KLYmqgkXAcPI3mnaCqtON1n3v5WjP4cbQZQ/KBCVf7fXnTJ919+GA8YHe7F4
HX5CugIOgd3r2t8IgLKmCkgmmZi8FpmLqX22hQ3IWkTg2haAxcLw/6DuOK62
k1NRdLlFScaqhnWyqcQk7fF2Gz7v88uZRTnSbltzO4oDI3f2i7X1yIhFWl71
lM4uoVr/eY3uVgzArlglfBZz8353o8Osy1AVyCCb2yLS7EYjmUt+oMcHHGv/
y/DTHFeLBB07lYpcUvqgH/F1NoM8TNUE0kCTQMVzUGThZlN/wg2p+PAaW5cn
F+IIEOC2PIuJube60a6wUkes6fw0iei2M+/cSlt+U114Mfj9KcJpBUunNp9G
Q4nnddtawRq663qmER6WHiEqOzL2uXALoFvl0AkESMWWAASGo1rTEuAkzLm9
zF0vJmq4gNdy/qSA+fAS/ZVb1nIFdDnb7KhCfQRmjDXyk+0BoYqJqTA3roZR
Y3CbmFVntEqeG51Srs+J645hCJdheU+t4nOAXnd+Gn/okzd4JcjaBoBUCLAk
Prsaej44RK7zg5K128JNJj/XXhVPGhATd6F9BbC2pZwRA5RBy0ImSHXBZEZW
cdRaPEM191D+GRU7DJlA8ql4ltixH6ZPyFHvUTKUhmWRgvY0QYhTcK0denvu
i1QjSmZ4AUoEcPZ/dNwTDZAF3tYGHeDRhH2eWUbOp+r/ChRXXtSU7r2mCete
4NOXL6WgQyypFSzFshWcOF1QDUXU9HE5CO/RLODMM4+CB6bG9JNJ2e6yEGDw
bnUs9wGDn4AZxPwx717dVcAQIdVxWlcbltPDUwFmzp69mKYjx+udmiKYSJNN
utlhnBhnPA9o5otnIvubKgrmHG1Pw+FvD9QAlc5T4sHCZnM8CNbzPC3YNr/1
7zvhdnc2AR3LhRWm+EfZUDXwk7k0eSgMMk6m3NpXkQnuhzwGmllV5/VDnAuY
wlG2a4OMEUFv7CY7cuAzfq76TrrBqIRmhP6swBrzvh+QEN4LjkyLpWXTjCPq
owCTJB2XkcTvIUTF9t/XDvX9t0igOJovNlbc+Chwkls1eGjL0xgMl2vY/pHf
Ua5MYCWZT5ZsoHxTwgFWlW110TO7AR8e3IW2gg6ZEFtEUsYdz0uSg4dqL9vO
YDrc72NUhMAy4bFCtDkog6Cwp1Pxcm2lYuXM4OqvBNqvo0+2AfLvBifmmuj/
xcoaH7Qf98qszZNPm+N0uC5ET7VrBhEUB1kr5er36MGfpzQA7ky/Ce8tgz99
oXl6RbkiGXIeDDAzV09DHeHVL9OQ0JBU01s1LWyDKVfgwo/6NSImU3TgydQ/
0RaaEakVPl7gRBe+TfzIaVX4e6FiQc33SSRy/CGbeiBTP0ej7b52BtYkHOL9
cqkv71BhwR+Zc/DYSQ9d9hQZACfQwep2iM+0LVWFaAx8W3HZBj8RpV2LZVIn
ZBABT5Rl1NxtY2DQvWeskPnXmzd7cEYlsV95

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfRBMKzk747n3mUQpBftifGoA/ooBtHEt4LjmoPhi7nJGHZrzjwxYlf8XeDi2LO+Ip1BLCXPqQQ78otCc5mDJ1Tz7tq2C3zVEtMeXFO2sGWMiyV1B1xoeC7B6W8T+pO6RYdmaL4pZYihbKLkyhesTkWEdGRQVfV/2fRD0dHiCG7yxbdyhT2s8F7kHcEaGPAIMYLYPZzjwgIKgwYeqeqXCN/lmkHWG7kGAXJ1g3a+bBLz5ieeo24nWxhBPP9YdP+J2f2uK1HA7ev1OJeqGAslMI+KG2NLcLdSel+GF98s6kfrtfTiORlk6g6hoxzjPihBXgcyD66dYyatnhrMXls3tOEfHwmqQRvQFSvTjvaA03Y29ZEq+xpmbpsVZrH/oftznwXmqpDlVXVt4dxWmh0C+2u49y9RKg0tgQLDqM5ruMBKh/KuuJKg8J9BNgIagk9pVbM20KXS5OtwiHJqgpuCeXE9KAok+S6jPG3/s2PZ4ExMmapV6lJ73HPtl86b11F0JTKjAJEzUW86yJ42s+cgHJoebtedTxznTwpKFEeL3q+l4aPoICpfq3Jrz6ScTBpPHVGRdUviaq7QJZ2/iz8wseBb1mo1e0c4Pi217XHXN/b3M+1x9ROIjYPZRFtaVInpH2UToVZpOsP6TM2fxe4BLJykGa8E2bxLCK+J6TikszwAMQHQT/l8TcB8lEyF6l1TvUoFY3vWwOQyScBak1GJxAftYtQgWuhA9ggJAK7MGUFbV12bHl7SfoFDAzfU3KMmvhmWX8QEUBqHC3CBfUVVW7y"
`endif