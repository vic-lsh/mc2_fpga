// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LQy9nKF2tJ2uo+cm7eEIuAUcGYmwKMx8heXkeuJ2Je73V6XlV/gXzL1mbPNy
vSBun+VHdAMG9zPKyxn9jeYvsZPG+jA96YNgqSt/mI90uAnky/cHgaLkOsUm
RMHS2vGY1UUiEVwfvIGGH0FaiDpAD7IS2a1NL0qO673id2QOctjF/31SJpeB
/eaz8H+TRWQZKfRR3QZ57rbA9BfMFjmA9jceamuv7sQ7vNLAAQlpagfh+M/B
u1DuLO8qOp1sc9Tc4bFdEOm3rDdXn41POhWaLgGhs60PdCU9InQSaoNZuWQf
nqpMgV/YJEf7r97WeBkiT5pTeNIx7+fg4KeQRtD4uQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VShr5nSM8JqjT59BJd5GN6JSD1N91CtATBfNYcv0h7xvtituJP+y6DezET5z
d7ASxkFuloVNbpHSwzFov7g6HS5hKAlk3ME34eEDnKyyenvr5tFnQ6H6O1Bz
D1/pIaZqieb28Gqp1JBPdNE/oEAmtwEqNfy79RIRS1imA9BpsOC0gSGKGFHV
5rmZljivZq73RTU5QaZGGZ6XEt11xux7YsMohapn4K6kDoVx1KeVHRjH2j7K
hJqjlmC9tcu/V/TSwWV4XQkEh7HPLSQqdPOccE8lAIHOuYqv8vBh1spw2vT0
V/ZWVx+ePOfViMGx3xLVWpboN/F/Gj5Qajukvod+tw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VV5TC6jZ2zlNO+lDjs7lvlCAKhJdHby9e+qTbM2URXrg+1lR5eQs2fyR3gnf
tcfvkdaP0qCVtqQoaGfRViXUDYwwEZvhiMMdkcFBCZKsqiZnttKlXGbXMJRj
42Hoy2UGzw62UJuEhN+nhXN3jLnVLGAjig0cZ2aWyRR0vq0pssTSg3XRq2Jl
nDB0udVpgrh0wdHFdb/4YbQbIUBPOjdYrunsSAX/UhM4yZ4z6HM5Ro+X3VpI
q9UZ88CDFN5GmOUsPFIEWae7BQZFXzubyghI+Kv+UpwP3OTEZpXTitdqPA+B
HdH3CpiTN3zzo1f9qc8+Zmeo6yst53+1d8vX0uqlEQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ho9luW7rJZOJJleQDkfNdAyGUFc7EaTfuGYNde5M4SXgc0846ixYVhjrmQef
/pe7HyzGchNFDiOoR9ZZIEmkF+TmpQlAqisePR6rjiC5/3j8TvRBNuoTkKUh
5S0+8oSEPCoCkQRuKp0ShdkitaaBLmeO3J3xgBffw3geaxbDrlTCv85YHW1t
tSWVlBREr0F0v2krsv7VuLPH/bAHNOo/vlqIhN7zzesssZ4CsNlzFYPFrahl
i5BX4q0zMZ/ltT+FFQca1kjZeMBbtFJn2w0aj7zOJuaGVnjrsD8+8E11cvbu
iTPhKLXIur8V0NLU2mgOl/1ywlxUIqX+ftdMRGNU2Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VlFcF2Po7BlOP24j0ylePA67aEsk++49C+BPKNilsn0kXmTfUjYlXHqOLOwh
HUA5d1bXv2W3bXiSedIePbBA37o12wFnynVxMpqgl1ir6C+V8+gqojRLMkDl
9BQOXYx1rbOtatSB1Tvkr8UNxGrdhdQNuiqMZBwn/6Lpe+h6Vcc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wgZY8TwdCzWvmWCOFTFX7MkdBJyIV0AtqKw7Mj9kjSHIh7ONZtSu0dQjudI5
RuIuE841QERpqS4g0MRv7w4F/67ddaPbfjfqp+lB0n31ZQpfZHKbiR7C8k32
LH+mRRoIQ04Ysv152iWCEtGRb8ogbgWIFwN8nnKprSf8mmrqipxkIv76Lhey
MfQQWcu9WJF+rI2qdzkDVsMM5fDLxcX7MRQZxrwb63sFbZK0MQIy0oObGqfI
55tYJ4AWR/eWGH6gsRjo5xh5jbgayL7nK3X8CnPNFEiYsz5VyARXPsYTTOIX
Bq7pAqVL5LiB1vqb884tDoCpvgsBfXq9R2KGFgFimu9SBb2+FO3kD+CprB++
07X74SkIWM/mJEciSPiQsWZBGNvnIWAGTCfha4aH54ReYIsotsaf+AWPaocG
ylGIcBIYTnKrDwdTM7V77kM/XB8wcpXf96MEH0GSMXca0/fE+LldjWI8hcub
pWajA2JEt365pKNhDQ3T4MyDmyiLQH+3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IAPVlVy0hXs0RGQDO73SvwM+MNtj/oC08TxSJStmETu2ub6Tv8oaYGWWuEyz
InMah0rsCF68f2l4hG7EtdDLMUeVvP5xJmYpng9bB0myontALNJPkdoiigvP
RMJdMHXpAhPhhFhCB8YU793ELpM/pMUuYaQg76tVwJsutRgesCA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TPV5e0hfCmNsNywHJfnsGo8hQ67zYEsGXeLWnpMNx6wrfKgaFYCZvuDGCPWX
n+B7X++0M7JieUFq/VpbCQLL/BXCqV3bc99LvAS2G52KBr6NTFqKyvs9ggmR
I1HnDcmcIJafgRnjU3SSlHZ9rQ13Ehy44fyakHtTH0IkxGAqM6M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 133232)
`pragma protect data_block
skbCtHKceu2NKhsDGfhSmIVktKlk66Bb+mpqFaX+/Dwa/oqF9bbNQrGz3CqA
pn5o2sjVLkaZkayy+UFDWCwAD1DCPE3FVEfamhLeaMZ7P1rTRd+ULxjjw5jj
Cu6QdQx6U5LZ/i22tk4rtb3O0ihpVIFMMGcBvG1SegnYo54SdMbLIP+wQBUg
M5CvZ0KIiuNHvLKG3M5OjvhRmdDAxv+Uxz+Ox7kx0rOwLkWARi+whmgiK7K5
gtbQlwP4IV/26bIP5NnAGfLQXa3DZfRuxFLenUOLhSdAqCeD3W/s+GZqLkjc
SbWCec3zmB0nE42w7O9dd+KPdzg7nE2ErDh0FZMgHQ/iIRLW7m3QFzGmzeKZ
TNIeTfDauJciw3LkJ7Lo7D0VElh+2Ps+MXvL32ag/yE7hofMalJ+6qvhQC1y
PwlQnHK1w73GaaNaadvG4nNVaHVWzblppEMLlMK2oVPOtMpsTK0gFCZDQ9uh
HeRXp2T6yjcniBpzbTwR1LhNQd3GtDE2oEhQKZRnh78CV7KWVtvezLdp/Df5
0QUrbk7v6tWttKN6Uyg8jNHSt2dwlrI0vQxgaTPmHp8vaAc05/yzuk86JAte
z4XJYOU+Y5AHGJdtPZMg7ORRapKb0wV8BsCb6BmvdF9DVcJDFuX5dTkuar6O
i0eMoFJYu4OzojamMJFJYjiSDQchWjJIEJ0/h8nrvmlzFYiLHMCpIiE9p6dE
eZo/Vf4nWwNa3YDxu+IwaMr8pD2LfkEDV8iuurSM9iaeiYEyMWwWZYYj4B1M
X6ARUFTWWqxcnDxG4yG1CSIKlprKf650PwmcRg0VGif3WOgEA2lewA2h0FSW
ILIssjNKl/zmUgcAhYmTjmcn4KZsB98IS/oCetqS6L+68nvZF64fb5p4Vd4D
rIHFCKZc8SbXfNyvuDnMxoqc9HG2fcucEOBvGfzywnt/333f4TrlwSAizT4B
L+CIY8SpPPcrcauMZreRhaeOzSxNZmr/jsTBkFH+qEgNL3CZ136v0D/p70ig
fe4XCR56GA+jIiNpKCGJGAAArxOEK36X6PL8MC0t2XfgMe6MFQuRK6cTxXfP
BLgSDK3RoWDgt8YjsHW1sMVX5x/3M8qQVoBiEnq98GhUQisz6Rkb82sOjqTw
OHrm/s1ivsDsuWjFzl3tjrT4oq6KkQI37E4kwzXkDB8zhNrAwWnrKg/eHJ5h
4mLnjXR35sAMmvs2ML1DSRd3bi7M3Ru59j2oRRO5Uz6/LNzx1ofr3dbTR3CH
A5pEO45DWFez6KFr6E8Z7Th7yR3AhuJ9b49t+6q9Rv2Bd9CLbBQJCP5R2527
2Grdk5opEDSeHfMkurdIY7z/QupMXBGCyJoAIacllG+lr+SCf8mPfYIMt/My
ORRCoyCIi1YaGWKTIxyQa7/S0fRKxsi0y7e4zk/yHI9ktsm7KjlBNBl4LB9S
Vf7v/xQHno6X77gA2zNSWRNHpQFa5dO3vBTJrf9L1lM4g3H77LSxevgW8usi
aRoNMa+ahMl50hXf4p08v2ddVq3OyVK3duYqFPsVcpRXy6DBcW5OYgDpEFPu
ooC4C7c8JbEJJmgStP7+HW++fD2xq+9BjaB7PNeoBYjr9eYjxVmlatyNvz4D
56Qq6uCo/sNavFtio7WxmvBl1jInj5Q1uBT9ejsIuqt1mYGiPUUBNyRsmmu2
XrIU542q9sUppAqq0Ci2AV1g9+oqrUXd/fIlxAfFMLfl5b6ikPeAbhJ71ha6
mXI5YAeGDZbviuDzRdONyq/wtCRUZl+JZ2F0FAdaL8JpEj80aBlYU7TS9/z3
QZIqFRjKAi2q22KLmU2KJq633evHmdwbUyFiOOKQn6NXc+LxVMieWIBkOCx0
fpB/AUasNprU8Rv894F+4/Fu9wClNqsoB+6VT6XYOgyI7a8BUVw4E3QztBWI
qlV+GvRoaPR3y/dVEIpM3UDO7LiQcOYBYcAyBOB0X+EQLCNcyblpV4Q63atc
egkE99+mpUuMHl/5x140hlZRoyVZie63hKStHJYZD5MnZVwzTvBqy2A/9Lql
6vrsCO8jzXAPMHSiQ7PjanSOhq6mKNhGYLSYBqZg/X9E1ineK2EmJn4dCI5g
Iqh3RSvrlEW0S4u3XBTs7VGWxwuuDY9EAgvAGLyLV0X2P+1RaBMus1oPDBg7
Mysq7Tfd/y6V94fCRWZQBSohJNfgbOC7xKn9lTA3P+FduT9mH+IExg6ty7pB
9djitfnLjNnB8HW4GYkjo4WsJfNXm8BP/Lfz20I33MqYOZJcch918YiZeRtV
kQ4XnzTwsgI4ghvNj1UY4b7/rhyXI3nTn5UPzEzpBl9tGb6GoO3pE4ZkVeXs
7dVtsoxn9YoUpeN5CYxWcSgg4fxJf47NGvDfXzkJWwft6TzuiyLSFrS6Ww5L
EdB+t1jUR6o1SlvldgAgt8SWxd1bHZWo1KlJ+8GvSb9Hl1Z4lkw1EPKCq3kK
YZARf2lT8H+nQmpLrNRHVSOSEd2lh40+nhpSh573RSoYSy3EF80E3NFU4L0i
aFslJ4idbMXe/8RZZJIWO5VMuBzvyTiHx0RGVpY+5FWaq0OgI2Iyul5wctT7
a/f58Rl21HgktjOOj2OEFtqrrLvYBh8eLAsb4PQKbTJdX6T/527Prj1OV8fY
7E9/gQwVLi2fWQDmlO1o79zIM9l0qrXOx3+UE0byChIcPjOMBORfHj1iBCrg
9wcdKTSXV0UJcGVFtx/usagQU+6hcQoorNLhija7P8Nuo6uPC6aRsJreT88P
zDVVcgD3SDaBq714vzvPT2DO1SZo4IK44t7I/4PY//x1hLeIIYoXEJbSJPoD
jNtIeVXHBMjiefutuoD8+C5LPX/oJ7Mir8DlVtHx/RAAGBEYd3K55FKJxx3M
oA0psSpzfKWl1/2IS12TaHBfDParWKUQhPw7F32j/FRpI/Eh6MdEiNcvPUSj
bLgf0Zaf0OaStyNeBojbdKnEtKc0BdRCeKqHib43Gkexc8zINuvg4Gc0Iucs
fO5Wy/qREp9kRAhJdjCaYGPHsXwTZyAOQOITBptpYkeeul3U7WohXWBmf1N8
mfhTNR1i0cidPQ5ITbHViKDng3X+cAEzFffaZ0vR4ZkV7Khu2KgKBzmZjHAw
3zbYWBNxard0t7MY+kkwAzPVR8IioGOKGOif8tGkneD1IiWEgD1BBidvn1JW
9bVvHPuZvNXn+DCgdcY2vAZglMe5DK/69TdyeHP0bel/0IY9fkPjMY2Q1Das
9zF73Ee/8ajpGDsyKQj3v3WnhO1q86eXRsQ/KBsWe/BiW6I5WMS5DCeQTjIz
8leJaXFERwBuxnMr1SlArsSyKLWEnhcnCTI4BQvI6lgds+SusHnXtRJBFvvP
4QUZCAfoyr0+v2bSKEXoyIjetqXSRrT2/t6LpD71m5DQqzeV6nPIARd9XNjV
wZ2+zUTU08zeFxf5k/a9qLAo7a2rUHnr0YTcXZMPtDVhnWFLTz4J3qAPa9gm
/SeywUiKQ4aeEIqjNJDQtefJ70JmPcOTzphRyix4r79y8pRvxzmMEApayEUA
FZLzDxGIpoirz7mzwWYoBO7AP/2K4D4sGwAvZIrz1isEd10XcZGJGA7GfIG3
5tvNnp1xfc7aUCgXDBhmT7Z9y36/lqzH43VqnttFSNrXbDulh2IeUX0yGUV5
O9q131LJ0nxG3ALGVkEYY25kAqZoOuN50+N++268wVq1TXHdnIDVb9s7MmH+
dbjf8X0QaT8CEGjo+36dh0+f/HOplJO9otFwDlFnm+I2fsYIMMWZYwG20kIF
s5/zb3iwHQ7Uxst9cjGUI8GzeYm1lksZYrRWF+rfpC/1Y8FBifXUVYvZZQwl
8j4UbB0pysvAWeo/UZ3h1pe8Y9X98bVNpp7jTKagTDOKrQwDtS3tdoPf+WgR
yZadMQYS/gNQFF6ebP3EXMjsltC0EvYZmjCffPrRhke92lUpEREHU4TI/Nmn
JK4zWAwoH4CniK9L0/NktVcf15yS/QjDOHPGXas4DXhHQ0DzopMGRcJ5+jnN
sUsvJFThrWnp0GQDXzlYDGwgKIwQgZpT7/JBihk/dJppn1r0vt8UFrUUk64e
yq8LgjMDRsK/C+L/Ute43V3UOsvVj1YXs/n63M4J8nx4Ns4riV1CPNKblzZp
bvI8LwJVer9OQC2gtLiH9VHm6fu+0FnNx38zQ4TaJIHfLWiyU1Xgja6ZcJp+
sCmRvx4q8nVubCzFaqqfGGgFLKF8iAbFIQ1bSGQ6Sp7AWmPAcLUE2bLifDSB
v1oyoHVs7PduStZKPkAIymCP8Is4IEI+RuM/2bacmsJVXkOyWMP5dIQg+0JV
1Ej3eKkyySZ7JV01mYDbQ+8clCsjNYD82nqNa2KAq1W284ATyTFD64UwWB4P
KS2FDuaxhE+hudFVkgafDME2/mCbisAB8Dodc1aMpQErOLSNoy61xfCbtuhv
0h3VOKl8i9DNbwRD8+JtgeAgp5hz04vcjpBOs738dz349F+kleEtK6ilSO5Q
d8/Omk3fAjX/59jvGYJ+IyELV3OZA9G3d1DEtXs8bPEoxdJEc0SHeyqmfSaN
1lCEHIPfB/GFDZrN2YuC8eT6/ZJXBcEZHdfDRNimvMowPOstA05MS5H8ShAE
jbM5D56urJ3Rd/XVFesKIIGk24LUk6agiRmSWxsydRqnoGD6yePQeWtP/SvU
/vXIW3hCGeF1w6wxuu3JyIk5pcOorggYjNeow3j5Ia6fkC5M9PPh609qTIga
mRC0Xqfaengb5kkax7vZi0OWH0S+CazYTvkbezsfK0rfIg5dfLx4+Y9/btt6
uZNSZrXbq/iJidmxLfIj3l1SIhPSzGzwYoO3EqPfYITI6Fmeq7TONgNsjEkW
lsiy0zRkpdQ44y7CsUhaGzsI1vN43eZtjdCN8GMfhJgEvY3Lh7CicX+jrGA6
eWcp+u3egtJuEndLU3OKEmMEkDnAq/L781n75JtryVXkfZ2DhO1gx6/A+cpa
xrgw+Xba1EW8fFZkEDipW4nlOlwSvk2it7ascS+YuWlPiwBa7OUDz1hbxz9n
n/Pe/NPZWshaGpOfR/imSTieW/8NwufREPNbjvpIg/ATtaLeDkzvVOGWgSs+
5URWbslbRDdFmldm2p3Lx73IBl/UM4N4h+ahzsdHQUNGP0zn3NMdju6N4itU
hhNHTnsd3DkZyE+Jwlnckbx9ucBXrGhUE1qOwNfhqRFuWeMQOyqtXkAyJUgQ
dj7YKOGvkJz+qjkaDY3PfZVpDm9hY7L6Ow8PuBSryzWRqcFHx2nLsMTnfr7o
Uu2//apLtEfsciDrw4rSYCgnDmRLVrHoTo4cMVkNOXeRRn6PYLNCIvUfRH1+
fhbIlcZhq+2drYKU77Kam5EzyyhXT1V5D8lDjFWrDsMF0Q6lIzpWT6LddgD5
55RcuR2ysPk6hddeTgLTUfRrXGU0YxI4cVKcn3ROtYgQDp29rdYRYa/bv5VN
9gPFhRI9XmkjqJ/BDYTJUFrATE7ETIuIxEbbB7uz3vItT58k6bffNtxMLym+
sTmn9yyYCj/VcpJJzc4dTbmUQAUEPVjtLeUpHyQN1JNLCiYTP+ECec4OPx7G
m+LwTlRvCwL5/WpWbaX1s1l6srKsYet1Pw+uOrB5NVuyIK68sqoRNCPhHmxG
D21uUB7Bw/Azc4SfYXcC4fwrnZPWJgec3TCc168FI9kAfTSdH+67xTv7sl7i
FTYAuh5BBL0+tj+5LMaD2kSw5+QYfjGkx7VaowdIq1SfSbJjYaJONgM6M04p
mzkOchRQkknCSNySVk+36cMirdWCbVIKpxAHbnWKgYq77N2Sp4qe/80YDkZs
prbgNJXBy8CXT2WgJ/08OYUpyXt2aN6wVj80I/O0oHXEoF/ksBqYjviT86Ep
eM2liLCzBOkRGdISwTDX0aMPHC7KNy+lGlTDqeyZgv7D9Zf7v/pNeIaXLETC
VCXs5lgCamn2byMn6EcU5ygYQf2iB2giCNENJdfAxwkfQUQihi9LkgoA9Ppg
vnvYT6FaqJTlVymSTJitVri1I5yxZ6lBaAPG3+xmNETZzjB80vW6RYobPIDj
qYxB3x2A9sW3k7/lTy/4XoamwNyUno8rMYVtTbQ+AxXD+hpGFtEezoiFvVhQ
r+9yp2XXfNrtmoqzlaJO9JopzE6iRhw9li9/MLX7SIOHkNVpwP3AuPLqt1UY
Uje2xbfQkGqwluWJvM3HyNZrY66BP7/ALgcJpOJqb1WIcsiEImYeLrfd3DRy
6ZJ+P/UMQJO5WPcSc+LyNy5RNTUQ/JH2a4k+vCnLCpLrWUzRv73h+LVlG7UR
kHSIzoV4JBWlZZnWISxtcCW43Q5s7dOhbseI23a0jC1sYlFaBMF+x0/kWYSx
p3AmGbPEosMWGnVjtLMkwOdAAn3t0RyUiWTkW3R4umEAPhmHUcBwyWVY+Lk0
go7bOnluC9XYMh9usVByCL1gosuXHQ5i3yfecMF6Dd4F3ObMuDt1BPvhwmj8
S8OEN/SIDRqx3llmbtBTyE2PCizN6t3aaxbPvYKj5NEobANvB8cir5GS0bKb
pMHHW6tMXh2p3Rt57oMaA9vg7236EJU/6MODmnIpjykYb1E0MScMLq1M2tRC
tjDtzQnuOn3JT39bnqKpR5kprhz1fX8h9TXMJBBKnzjT0tPnauTYimlq9yL+
TJ2YEDCRH90dbXgWw7lK6IQo0jPboo4ln3ln5LkbpFf8mpYgTmWjm9cBcZ5q
3fMG0xXaeJpMU7uop/rDULtX6AIEwdeiWSgIng3FPVLE3/qGrZd4T6z8RrhL
GIlFhM6NMoxQJBZZ9ys79vY9zJnFbdAzyq9kYiB4DaBHB+ndwsMXcXiL7zz5
rMVEzfV/ZBdAZpXg1AS06KLx3+gH/tQrjR8vuewAdWvlMu48dJ3UqAtDar7F
TgKnJxjFLvwPYxTZoXXhoiW5zludFoBRengElY+uvJT8k4kujtPMR6Gl1ywq
Vj1sTw4LK6V40tVfL3o+fpEFRPZrFl2Vfs6zf1SEnqhAVCcbHl7jSSwayHYX
L/ax5Kn7hIWuny+H6TYt/05tUfzmNW7M0QnqkihT7276lYRIKt7T6mM60UlA
hOPWMZxN/fFNXBQMZIJBfO+4aurTVJNpVN1njfjXYX+2XeZ6Tfy02UKcEWgJ
wHvazxOEb5xyjwVVBb5BJu8Ijqk+4kDaar46EjbYhFRT56ei7wOraugDhAu5
yiVF9Adn5V3iWqph3vDNpMT2IMVFnT0QYJODb8iPI5ffk/yrAykE/mhZLcXK
4It/U5KaJ66my/4sl0MA2x/VdC50kXwFXP2Y45X3qcqp0+qkm8HDnzx/rbYY
S8mISBqYxAdRtkRqCPrKpiSpMwd7q8Lnm7KPJRLTlwPXDiC4+UWHkwJ+8ZoJ
yPFpxSMZkYdO316bv+2lNEageg+8ZDCj695bBuNP4rvwz1IihBbRp0+dIoaO
sLKXOxRB55iseI7RB6fhBqI/PF9kYbHUrhbswJg0aBPrGYVpd9gD2x4YuV6a
5yOT+pdPTwpeFFMWuhbC/QFR27wUZdncvSgJ+7h9H9UQt0CX6ewoGiaXd6Af
Do9mZezI29mNQa4AquGxMcHl0d3i/aCSCSLsxrzfRlE810Le5nFpQ7mZFdFc
GD2AjBiqd5vp3ymWASyILSTE9XnODPxYgB68wmn+7sxQyLl/XGAGZ6TTDMr5
jnJ3J+bwXPzqBcgl+RY01UGcaMEYgJ9c0/zjkkHhAkmoXAbO4q/19DBh9o9m
ixP9882eXqJITFqJiOdKvzoK15NIKz6UAJP33Dijtma9Ag3+m9hJGU/sJVfN
u6NgG64Gb9xMUpj86bbBTo63SUfQL0LV0BpqgQi1/G+qAkYy5BtcgvehJVv/
4O5X0HekdqBmrWRbYxjtF6H3Y4V1uFfzhNP+aFn+kAxy2Wg1Q68bhwFRi2cM
+uFRixGwOxOaDby7ZTjlG0u43cR2KtwBQMJ1/xSg4diNNEs/vpKErX1PUuy1
Y45Xjh034b/v86awJ6EW8QuLfm9yDdyOCLBE86vou7Deb9N9t5K5+e/whTBZ
EalQkndTzwskrDGd+hO19fU4FQaPNHB+dKT0FOcqkjCZjEfPVJ+jryarl4z0
WLBRx+qXabtL1mLyA0KmosnyYP5Jx29GT/n8Dj+mmvdEUGFBqziVzWqqkwjj
fo1MNB+ameU7nBcTCxQP9KbF9Bv2dNHHgfXpZbbgxVQEZXSIXbsmFYg27I54
ThPh4bI4a3EeO+KgFcw6ekktfp3/0h2Kec/VyIJcefNGMZjIGkDrRmNjhkPZ
TwSkFYiehECscJu7A10xvpiq662KKBJrBGBZnGtddgizyUO/ub0AmgUwSd+v
f8nHG0swc1wZ0VSrj7ZC0i68hMQlgK1UPQVKfR8UsQfc9K5Zh/DexvsfIVr/
3WrFqzyYhGzePmitNGCHUpkHWkwaEDpF4tLpJqkf5f9PKw/0WrYs+Xb2IgGo
ULXGh2wkN1BJBfdqVSjEX0XzMPkJAfeO7c2MuVvO2e4SCvL1ssmu9JLfudB4
N2JHxGxieblKbB4jTye0WztXN92LbfrmU9enaJiDXJStr6dbLZzKnTyHBcuG
OGsf3HYuA1+iR7xXOrJ021ms31sFw92FCrIE8ydOzeKzs8oiBaNgRbv2eWJ/
Ftibz30kYbswi8NPUUNzHm6yUgxqnm/rw2E+a5Cqe5NWDj/aXASAthm2Hv+d
UlRx5tHoQ7U8eTTdFsQU0XQWBoJqjmEP0XsRpay+EyyU6LJztyDlx3RYSrGY
m35o+0BI1hZPHFA5zoKsb2o2oMf8FmCIPRpQUMvjsDTuIUDBdry6oLzvq6ot
qwDkjbqVXK9NTxljRST9mdak/HidXsgqAR7mUfLf6WrFZF3Sw1tRWcZX/e7S
EYkI7sda0tIdv9ddYAdsDWIxfjTdAXWGC2yayvnNn0tvXGVE97MheJaajp3d
hTJdSUp7gS3RwLXHxnI1KdfW5N88w76YbQkQnhtfI1MteI5F3z8zthX2HD9D
BzKdthGS1bd3X7Bp4yoLWlPDpPMXS0xJQXlxWJbw0GMxPAV10QBaLzSX0VNJ
RPHhs8TVLOUeY+SHxTTgairAfm9lZEH0WDm1pjwgBNcJWFBsXU6FQNyXpKo+
4+Fyl8B8zFzoCvrqATbYqefBBHnRplO9aySHFNwIj89cXIY1v3lPu2mLqMR8
CavQYhaslTrd3Hf503I/X+k6JFPcfWsh5Y1AdRm9CrPNwC1jyd8FDs+VtrM2
wfC4+NFNNjqRIDj/ExcfAno1s3bRBwBvjLGOlSouCP03nmo2SWZ/UThEOs/1
tW72fYwB5Mj9cNPjl/eFGPkwDbOdUcKKDxC9ANrxzGawqBxlBdyix+Aw785Z
YnUOomJr101DZUP094flBCpHQQfhU4i38iv4LK9m9CGC5elcA6it0EBN1+Ke
gomLrj4YV6mZ3c5sLN5ei2BjyHeh4mHAdGXZfq2w+A0ALPDBuMPiMwnCb4Cu
EYWUeqW3dMFb6v3QgDq8aR8cSNt5QDCDaR7E/pmYZBvqmVz9DIZDVERTNKXz
t9MYVs4nJ/zww0EeLRkG0SsAG1kDLsaJNAP7y41n3M2ipz057ieoXzSzGXN6
YiXOgYUDjZlZCedy62p3oXJefZ+ROd/Px4cwZ7IEvgG8lp/2kyH+LsMpEUPx
2DaxMdaReqy45qZSg5VxzKiYDfhXyF6UcsxwRaZaY2yvIKnoc06fGxBSKs+H
GwBmT9G/w6GUqNMFPvKO3khr8sL4fqzQPQE7cuaDr558lAcZOv624+hrczT4
tPUmn6VMKGHEnDAykCxiTbAsbOWw4J5UiwBw2CCNtZdROVsiOM12UiyUXvnR
7dlWaAuNaz8L6d/P1sFFc4einpvXuYMJuK4xs/DVSN5png7ipgRegKUaiL7t
SqVLy4DG9YjiiGcKVS1nH1fyJYhvtWo9lD0BXvurfnVyCbXtaxT28U6jar+f
jxPxR9JdraobgNw0+2NQo9Va0AvKAaiurjGJNCC+iMRTN67BBhiIfF8hCJmm
A37/jIgUVHxiPSDSuBKiZS5VVXSJ74H9Smdj9VgKWWcVRLqiuD4gp1kg0LHm
CkcqlQGAXkn0FVV7A2Qg8M0++G1Y/lna6QBRaK1Ty9rzr13yEpZd8qeKFX1U
SCH5SECYnH5CQmgu/yPOkFs4rsvCWovryECiCaKGKtx/Kxh/m1xN7Tmyw0rZ
Be02mAWDdarMZlCPeZyBhm+nYuQKfPZKBFL1hYD8vr+P5xqGRe7IIQzcIBHE
g97uiDva0t3FHi5qcReXF/7y2bKncIE2X1858XD2+k6I0wGQIBCqNMv3vSpU
Cblc82Fqm25cNB5DKr0MmY9fDUpfEO4tyEWkSip38p0vq9yiOeVlUUbAMTor
69/CH06/Jf7FH3Dzx7VZEyPi89UuToncAQ5k+prNuDhvERa4IKaPCbnlgTLo
45MDfs2bXLm51iIVDn/P74THZNP6/b323+iMZiWpUR/R+NE7gsWB3TNsXmpt
UGPPYNKCOW3KQE/j/nCKNN+13OKVyp/wc4ni6LHW4sHhuY05ZTyp26rIcfdP
6wyXbQ+hz9aeJvyNSsYnLiKkDXNRuySOXu6jiFHxBd5puBuh+7b/Vy6f65mT
1G3PXxWK2LmeYZJFEnRBL7HeYyyLgMw1ayXRU5QIQPC1YKHIRcrsVE2KmS4O
x1taBlxnprXzRSKSoJg5J/UwVK9qMm2vKCZotMa91NTyAQZtVGC99Uc7yhD6
sqjQOOVMlxaTrsoFXuMl87yooPEF44HUWfzvbPRjWn7iiZri8QTZPLLqS6jx
Zd1he9RGWXahnk7zXwUCcWjwiynzqvcafTZAiiHfb/CaYs8T5s+bQBWbWOMs
diqH7Ce8TjOBCMH75SQiJxCsKLmm4LnTZG0I7IZwELrqef7fLUDe5Sz/Oa+u
IlHFlsYLcXRXJz5F7tepOAkFkMeDKvoL/biBADIauYN0ZOAiW4Usy3PLcEY0
1xeGLQ1lsOGvDIYKxbQ7MekMdRJzeMh70NnFB2hsYhVac88uS5Ad0M5A56Ug
r3mV5DYFO56lnL7U6D269acJ6dLFo4PugYS8yfvvpqLTYTnY14D6L5+151gD
0cB8ffY2Dfk9kWgHfIS+AKs1T0X6uOtHdDSalJ59EEtSyTOfZq2Pq42qqqqQ
9MyqW3lshS7KNS77wbQ7z5BDNx/oP+mr/nG43LSHq3UpDllMOLAhfNYpTGK1
4JaPHPz+S5loCuITZU3OKNDfbmz5CJ55TtQwcMYCdx2fXFk0ScgqDClJ5iVG
OGgeA+FSWgnI/U2S6eQtkT1sQ+hWw1Sz2mrvzV5uNBQCCRq39qbgoNZhzs67
1sSjZXfv/YhEsHpcCj/7Sq9C7pl3ZlTQbtvELsDJtjpMB13/aQ1uzc05DyaG
//aSJXRM3uVl/fIIP1YpdoKY/PmF1Wjhqor07/Eq0XwSAtkiAJ7HOqSfarmp
J5FLL77+LugXplDkbiiAVbHWg1geBR7Lqbs2rDaaoCwAhx32GNT/4LzSjRrM
4VpY0Pye9z9rcjPMFtHEc/s+g6U3fCM0m1od8k86H3pEdQRNYzpOSbJE5JfE
HCp+eBzhUcVzEpJJ6nqUzGAkmFKfjRo7UaRqmFpVcKrlK9zvq2no2xSyiI0Y
2LK7xtcEIgxEPAer4FEQyw8mvHmeZzGcX8hRvqC37fDSSmFIdD7Ey+yI36fF
t+j08OvO/ytTa4I1EuFXi67Vkwi+r0ELqAWngC2wL/ivCbDFIAGy8Squm1+w
JoCIMaI8KitaglEWmYcoA+zimdBZirjcJagdv2kCOgjzHpM7V1iz6a/Czndp
y0KnCrrsI90Tk+e0fPlV4LVwIpMJCHcW09tE7vUst9GRGfw5F5HvGvZIdwyy
ZLuK1ZOhOa2oTgVEfHjhqZ49BAjNEiCko5EO0yNoLJAhEajw/kuGIgBqzCpL
zj3apshrwSrwtSPE3p8CPCRR5Fr/ZsnAopU/rDCIpxnh/8psJ55Gq97eGTvB
H56JcuQPLYe3yY0a3VK1p3HGEGr6IscodzwJD7ERPqaeoDvGcQegKaihFo6Z
yL04fo4SmN974JWid5qZMej510uANnuz674bGW8toS0a4TOpD/P5Z0Wfjdoy
KdTeTESfnAw96WwdBzBeIFSfyyF+qrVFzuraFIGaSssek7GfGzP4BB2jAD5B
ArTieeJSJiMyWQleTvvz/ME6EBFMhlbvA8V0AhKNp30SGuUQs98pGEpFro18
JMU2x1sn9fVIsA7HcA1qxC1wCdKpRwuB1u7GkF2gO3annRwHacsSLKP9hzO7
IYvPKoBxZ9X3mk1UyePyC6irKxqPlfColQYy+6PE8hvs/ZXrOPnZXCUnIIwg
jy0APWBs3ffK3NBiG/dRTHskWWO5DqrkCwy43QrzODWDGglSxFndYqDBbLFg
dJUebgL63MAWW272v7pCZctvHWAAV2YWU1ObIF+5WgV/0GetdBo/vypS1Ztn
a1xTd/DTuC3xwE8jTyA2s3+43yGa+BxqbgeYdAD1L/n9uWNueLlQWyWHaVho
mZIe6aTU8dr2ByOisiXW2EAoMMYdvbbLmaReB4sF7KkOw+ETlkkOXZGm097H
ZX7s6cEGcZl2Ti8A4ct5eqjeEpcnW/odOYRVSSJiCZ7qL9pQyJvLy6nPA9KA
oRpeFBuc+oHKV19FJ8iS0onNuUy+n+jly8NA15efNkrgXSou6P1zDvz4+Jg2
iaqpLZXPp5p7yYblL+uSfW2O+g+pWt4kUsS3vui5M9t8kufYQnzyW32YmV27
fbS6CZFcpYwK46tEhjZK9aw5WqeKWM9e8M3pJL5LAYKjMfHrTJ0eW09IR7cY
PAfFrDn4YcD2lZ9fF8gQrjl8YdkHeLvV7I5x9MZR7LgDoAsmv9HvnUnTAp6C
f2fdrEYVwS5BxcZkIoHK4A20EttI2ZyUUMSVmwYzt7utp55B2t4hIhtSAJEE
w4+0+1rnbwFP/+FbC1qpyl338p5I7NbdDSSvFZyDhORUBMT1RFDKbRW5bAGi
TY2HgE1uAi/zuRF/ntY/C30ii2JhKiSBncI+UZTVA3mZKoCSwIcmU+Fkt3J6
tckWjXE2yprZhADFhxO9bPJPWw76rnFTauU3X0Zv2IRNSWNlPDqlSQ9YjUHU
CM810ggeGqQm2Gl+oG5GK7fVZ4HPL36MwT+qpuXGdyiUn4bIKIHqcI8WxbQX
g3nKNpeeUY/jR9aHYHGXkrZ0zZ4P5zwTjcqUxE0ByLOPXifvWoRU+99ERXEv
qbIJuEvyH+U+nGR9e7eFQSe0ruxBnKcEE5d21NLkha1AURxoQpVTt4kVE1mu
ANQnJv/Ex6MYLTSnCNOVF7tZFEeMA5/1OH/VLYqcypqR5z/IvX37aMosqEvY
DCQn1BClvZ5n3Qr6fIe4ALhugKV+/UYhTm9u2ZmJVd2GTXEX+VTqLWCkuqe8
4tHQ6RiO8HzZm1+G3n1UHB+QdHWt02OzwlWD5+KUCsZWHVaC1KPlCg7gQXx6
j0SzjN62vzs9VfS20OpfYs4c6osBPbs5Uk5g10MIS8LwYC+DbwdIlWOWiZVc
A8n4cJLAp7/jhdCetSPGki2n9pT41Dmb/0f2/+oRz2j5cnq3tPM2oQ2ReLX/
xDrDpirqdhdUPMzqr7oXHvVnwS1J/fUCVrsSb0jshzgmVCZloexwLHxKFLLH
6AYqnl3El+y5U9BQ1bSkDqXVlzcOjg2TWLoU7rRTWFgiluCY2NSsTIOVzaEp
21syF0SdIx43fFEN3OnFH0PqDSQa2uog6m1n6uIfURAtwx6maO4+7qL4jqZ7
ih1ioqciflH4BWVZ0Sh9Lz37qpYZXQBmbp9fVtbb8FWdfKX53kUOMMpJ73yc
+eFJfqqMm/avtc6Q/ANj1o7cYp0FlBl4vtE2YTiR6wdbnbr82ts2zCPuMEEm
GZJWyzXJ/+dtzq00jpuJ0kL7XHJ3g2dbMgWvt2r4pWl+kdxd6ZepH9vOgzxl
I56caCG8wNZQdCaQb18Z2tVnOEPmemDV+fbzB8L10OIAH5/eBAjEiUG0aAjX
oTvcUmDK0MzWed3uNtdil81C7SvOHlJ2Buw41jtiJmptHVYPKDO3T8ynueVD
Cf/cZTNl6VWg9g57x1e/QbQ5+m5S794D1BJAJHyGth0djsX/psCZDpU6bTyj
hts7rU2d7DPfqQhQQCrdFYR+z4KNkRAtmveTs9NJPKUdcuGwKTz/WZcNNZQr
3dpdDnfNeAkFTtpvbIkP4Rq+kiiLIQMJfXa5YomzWS/uaNRpwZsKO0mPW7YH
pPEKu54pwm4PytPKIOSrcenvPfWnLgbVX7L4YczTlo/PxuzFgWu1cq+pj4LO
gBh0ZRETv+uB+XQ6R/5sMLhDiZ4K8TflMR7hJGPzuq/75sfcVw3n3H5x3htk
NSjjLIuPWBiLpyKFx3iM2ODLC8PfJHvHySB6PySDb+FYTq0EXd3JOO9cc9rN
J8JrMfcr4Rio6+W8chcRMxjXQ+VYsa1KFqlRTMcCIG1wKhoZZfwX1Raq2Vi4
tnXo/0F7n4RyPc/1MqHNcbAfYn+w3g/8BsN8XisXfjskmYC0O9roiJLwcr9e
u+9K2ybtOTKkKcQgI46aDcbCv0RIcqjzFCv2PpMB+bCi6/Rm6NR+XUCPDyMP
pczKUn8M8TupYzaS0n8wj2wFuavI61NNPoGwUJZXd9gkyzIsS5/WcojGwkVM
xaO+BZIZcybVm2JPluzCds4TCLTl5xLtzcLAdXT/Qf10NioXgc09ysQVT/GJ
eqbjdcLWVTtP9EmoN74gchg8E5wHVTWx7YEY3yEQc/8DTXFfGMnRONP5026Y
ms32d4mQxw+296fSxnUV0N0Zo26wCa1p1yEr4LbpxnTjgnkTfdGvLy2cVwLE
KJWtE31hBqD+kfsBSO3k8OpowXPgvBZ5VAXOI7rbD6TbK3Zj2yU459wo5wAz
nwaP/9GoK/gU1UtTfv7yoVaAx/Vy6ZlVYWnGRlbnbvLihkUi8FtxJlMWsCNJ
8MWzK2xLm0fAcj4VFAIWGKL7VzuVIT7yWdHkOC2Je4gxUtzs5j2MKvc34kSF
jQoShwwZATVE2I3omVHPPrDOUUncW4k4YtCW+i0fP8KesJ7Ih60uizzo/cMy
KiJ0Vf3aNb2xH244t5sBp8Man5eknCpxlgl25X6RW+OGkrjUGHCTeFksWFpV
sEKS+jtwr2I0dF19ZM4lnunk2SSI8TlSh5v7Hr/YhCfYAR/GTZlFVz1mWnUO
Q3oDWIu99cXzbjtt09ElHKBh0gptuYdT2AxRU1N4LB1ER36XtRoyE6Kn1fLT
36R6Yq4iKW92cjKEx4DhKvuHy7OvogGnZa/mzZPaZ8IggFPWJBenTP3AguMc
bS14AWkhYeqFPpWKiqI6FuI0+YBghxAexIpxf1fzgwCWw3ARZkzT4lxtAk1A
lBGhdS5vochz2K5c+Sg/yga76J539zXoTKf/kOCTyeKL0WDbwlWbzKmqT9b3
BPZdgxTAV6TMCIJ8AhqBUvC/wBbaSCREUqTBXQb+ZuRB7YoVnRInvrXngH20
E37Gexs5h4J7xEkk0iUPV0WeHBEfErW84RvDeeYOt4TPXY11OhhOiSd1PvL0
pbLWCDlsmQb0n3Z+gPA+lxGva6XBXEJkQOgHA+4Z1Gwl0UHwnLewP2zMbQjN
sXUvPWaqWo1vFwGOeNHqvHWZd763t15n/M1j6VR63I54YUdoFeW9ugbTsLEY
whKS44vIMWMEDPAYopqajKqwmOd4e4pV8WqN2K31F4cdHEr8ruZgWlLvZ9hU
52YcSO7RaUZO+VU33EdVtSISV7VNSKTBt1QJCZc/yxeKJxGTwgV5h3Y5Bjy1
FH3sDSo2fxS19i5McMo69k4gZlqFHUdXRkDZejtSyAYqAf90x8rID+i0pqkv
BEHwu8AUcqDiO5SvyRWCKz7AFecZ2OAAmhnWEup0yOs08u8Yog4dUpZRHiZx
Y9VXCgRZKm1/VLU76cOX4GfMo1SL5DeVDQ1GBbGXIFNQj3i3WaImTtwjyg3x
uBm1BunDmkzpfwjg3Z1yRe8xon6ld46Nvj3Bg8lB+hfrgH40ObJbsY/L7ZMa
E1Ift7KAA0WkeIUW0SY4VmVfHEgrGojunQJlEee9gAV2ZwFX1v2Y8ieZTroq
8+nwHbWACCAcNyf55WuRsf0/Btcj8iZ8J8gRn2BAST7ssroRK1EqHfskoiGC
G7Z8tMlw8EHa+GSYZmW2Vsr0g/Irj+Y4KC3JQNFrc4ESLDb/kbORBc/XOL+g
IVPPwb7T+dwKXiEgjOLPPYdn296Vfp6qsfkSf9vE5ky4mgXJj5esgEc8lFAJ
mhlpQdpwdJLSWxkzUozdJ2n8QYxp/p/gL/dUAc0WXChhMzL8rwruq81nyBuh
zlSB4O5cMEWB3/KGgK67i4zP98ytFUzagNI4i+h64qgtlJGP7rQUNrRfw98Q
pwnuuEiTgMcQ3tZwYET4/K2iXDSLtu0Xy0o0xpcozsNMpp6FcMq33X3lI+Ld
8aqaN8wip00x6GOyRDdLN3I9q92S86rhGKnR+rUaLoyG/wnjZ7k0c9tvkH2P
3EXSM2pULs3vPXGvdaZKSxkd4PJbzZNHIE3oKJjinOawJjxwDWiMuscRVlMp
Bq/NKvqW+dT3x2DdqtVHdJPb4jAjeQwi0xE1y/L0DaeOYVCA186DPD2BMLOU
nX16o0ReDwGpa0j6C2zhJkcondKOcGLx5YyukjBLmryO4NemdVdaQJSVa9kT
NpkQINi6Era2nM9YnA1eJYyY9Ho/M0qgWfaxsJ3YaAPKm41pTbsyJr1fe3Ri
ozYJ6PFxlyyy2Z6AWlICNuHqqSin9h9PGX2BbdgblTIhTc/yccLOTxo11j7T
OZxHxb4RUW8s6tT9OShNIQO53EnouZijRUxvIfep7P70ctmaorFNEFL6vOOZ
NDXgZfDrbE0cKdtCdRQOs2I2i8iKAgYzt9LbFVp41NswO3ZXjAT9M5U988uy
4DbE/2wLew6clYdhioAISD+ilXFzvYGfoYrazbOx1AIm6B2WNaKiXa330a2k
vqvWxqPTNI/zLveA500TDDnTsehm6AGL2XN2vrLrCxwKd7QKgrEcwxQqZk/x
auFo+zlrGOx7Lze0BsCG6kurAgV0xwAgr6GUx7tRplR2tuluoRLVL57FFYTV
LIAwloS3LrjslvBeTdLYOcneSKP+PvhKOcfYVRd8rcZTLh4YMF8t5UUzZ+3h
oNGkn6wQcXTFdc4juAb9hmQ09OQagMSork6zT2s19+ytc5fhSFSDXAl9Gn8V
b8yp3gB0s5RzCgf8RfgtMZYpCNChUiPoeZjfvya8ix8noa9cPe44oP2p+MSV
YryTFbjTt1vvpeYbcRl/xiaOLEq5Z/6g7d+uvQJxTVlkWtOFK8SwZJJ2cajn
rxoEnopZ0aXY7iAFWoKBMhj25sgHOaBO/alquffT8zws5KTwaH/qO/+V/jVm
U8Wir7vaWu4SFHSYGyBNy6JtLTk1MCtARO526ir9Cl5agCzK7k38kfeaGiz3
9YBbW0AfjHIR/fJm5GfuvRfKThiZwzxK2L0q9Rj3LAZds7TRuBQxxPhcqHyh
WGlIYKrOUs97FkvE+WjFv1XuU5ZXBlL0sDmGEsPXJEzzbrhrbi4Hcj76+QEx
ix6TcHXc2xXpxH8Gxl7da26JMJG9swnSbBctFaPYgRFao5P8yeSpPFP5OVD3
zdQPqO7lyE51bbHzc5a4dzqz+XuurXne2nkfWoA+c09mqv0k6OmEzpVSX2Az
LaTboRn2ljCd1WFdAQrEO7r8usc6zUfgpzuGweNs4yx0qKN88z2KAWgv3Ceh
Rhl/umexo1z2+fF/2roQVY0YddYx6W+xk+g3Rt2gq0mOTUEBxiaRzSUWwQYX
JSqBfCO4feh62BbEACWc/golDndKZrGnBjsTjhdAI0UVDbasUVZ8Vfwh3Em8
EGEujtYqkktDPplQkbccBGZ9ucyxiF3lETPL5tSeUKoJNZPykGdCVnh44CCD
Bjdjl8JEfLNf9jGOCJYcmTZx7ntTc9RcwXpLvAOEgsM/KUkm7g7n/fGf3E/X
YKcHV//umywKiozFgd1MMijt/6YScNbZn1RcdMZMAx3AUYiJeslhjxtmqofG
rhQ4vtdquRTvzR9N5XvXVe75rCR4r6oOn+3KTve4Xad4kaY2rVji7hY0QLUI
at/5rocwFxuROBn28h33GfJnTJypZI4CdIll/TKLiZ0h8f3mhtS/CMzhX1xA
Llkp4JgAmq5bzJPMLTNe4qNZEnalxvTIrMz+G7zv3TvfbCjOJ4X4vWE6/VAx
tunhaSy02wCKBGSuwV2y31AdjbgjWMnYT+yxV4MOZOISD8jE3J7psk0mRSry
ghKSn7c154/7GVSymz/6eh+AjWaHCHTDMQ421brbZscnSiostC6/oxjHy0OZ
igXA6Lq8p8AN59BiLglpgU99lDO02jENkPaHG3BHCKBtjdN3cjsTxsZ/fE6M
ua8MhRvUO+A79xVFh/PPccrZLakEWuqjWTTMrQVdmEltBWVPDcb5UDldM5oX
ndjqEOmJIMOaeQA8xBWwezQaiy6GhL/YGlc0cCbhuorgx0LahkgHvPHXjnMH
sJstZTTijcG45I68QLuovBXmJIwrlQca7Pf9T4ze61sOnBXAJ1T3cBGCScLf
NFg/oVkRO0vnENPUFkf7psHCHNZy2nvqp1pLB6+gDmoUJowxf0FxJ9u0BoJW
JVxokWSvMLGST+C3OVuh16MVC3yP7WKsPaYqNLVln0NJA/seElgXq+GCuLCS
xvi1RGT3KIkqJjPuBE0JAarP383HK47I6L2a7vhitVfj23wlsNmDYZhYgPqC
Dird8cooZyOxa+blTMMpiyRPJUxjwPMgkoA2v8VNsdddArUtMr7bEPg/kPKN
6TODwK5dYRwUCXXcSBwvIMeBZFx9odOomJvkBg6+X9An6cgAqr2q42dMYWhg
NwF24FPpovtT/YzcMspiu/L9KfAENWzkTaZkyIIVzCZIKXAbiUNX+NHKqSou
v8NOyn6NiLeBauDeZV/kdzNile3W+6GqvwtPImsjo2kQLlKtfWgPiy+b+NMp
SQYHxlUTiL2+q8e5GOeZHXjCed+Iy7WnjY9YBBfNKsApH+u6Pfa4/OEXdsez
uH/KALdh6Be6jpKgzak9sA0VC4NvSjRh5hwGj4DNwebZfmx9XdVc4v7kn3xA
JRnjT3lB6stSW/g/owDebrWre96Fjl5dfT58dj/m9AMPD3G+3xU6WINENsRZ
4vdPZtwpOaGi+6lN6X74Bp1xLPPr6IAvoZnoP4ewTkJYrmcjCAe6Q4q8fCXo
R/8GV6xWkkQ/xI6/swmrhZIu6HwUC9YbMSI6YINp9ExK7z3caMOFDYKAyWaz
4VzRyU2afL4Bfa8hU5qlbVZxjZs2VBrolq8wKRKBxMqSCx0F52YtEW9VV+rF
2f33+m4zgQlKZ/6+Bs5LVcPZvXonybPVh+jE6snFiTe73l0qkTB5GRYV62GR
1DGEynbjp0BJkH3SdsczxT98ySjOcukCAQHaXA5QBQHB9kjcTP7sSgt925MK
ENpYHLP1RZ9MubEJrjSp1Yv0kSV/iij/8jRbVokqiBnj3rKZFl/DzeIXD0Yd
O5gnqXjdzcUmJH1TsydcYBZUfhv595LIWqLrZ2nkU/Qdm5pwvXEbfILSgjSQ
aLl+F9JDS8LZafE6OoAoGxLPrPj9kgy7SQgvOIm9bbjKaQwSpkjNjcE+ujg5
G30Q86WSO2FFEXNY3HD/DNf7IUHuLKlePmc22aKm4wme8wmqxGzi4A9VTaLF
BnMevArhKBguO+q0tO1lFdu3C4c4+F6FOeRQvZQ2wF1bEm9Yfdsw4X2soE1k
N6c0IQcpBTd+tj7f+/ckxgi4zqut+bPl66WvP6occXsiT5bYnfeAWFe9iuMB
7VRQU6Sqb2qDC8KdA8rujK7XEJrB0d9yCNTGT/aVNLLxd6KzQL7KYRh76M7X
kBIaZDtINGnPwwRt6u2nkqhgp4N3aN26qTCQekB/wmZgR9OKVdNbKLVazN3J
xgeApCQkVzGAA0NtDAghcPxaTgVtPUKJfwv+DVgVVBKK7d0IcBVUf+38h3jR
/ZylL68cAPGI38ZIDW7XWMz1u7+0rkaDDZ0Ehu0H5Zwpise3F0w4qaCZ6FnX
oUFAZuQFkenuGzrEextpQzFiyIuY8Q7+g0GwIf0R92ryEa8IQUQcSUtO0IHj
P2X/Eqa+fGXXRHOMbKLYAQbi11lkIJelgHXc6XnDQIXUbHmkicVcOOAFq/qE
GziHILy7j5NWLCfBa+R+dLItFelTRKo8bKnSHaKFHbW5EfPHDlFVFfS3MrLL
mfdGWMjEh+E1lb4SVuWzWO2s5slDR4cTtJsSc8M/LCFvaca0cA3wKUnuLNmo
Ekcig1EGkgOW1XuwqKRN8ZKI25xgQGrLWLJBgMrlkOxdKx/zNIvnpX8Iywub
0ZJWDKOkpFhqZsTpDjkwCwLDJNkC5LrtnQhI7jZuXgJvPMlT5tnQljdG+ZId
jphhKyl/5rwLmB3GCU4GVunfg8l61nLrVjXmu++Tapfzbgd4RIo86f0bkGG0
R4/UwvjET5IZlbrayLLDb3F9Dq8RAhOWCK1wd9hHToFSiIKaD7bgZi8RTNSI
pA6T7i1VE+jHHs6yxNJ2+YNhxB6tLuYhjewLfN1ZeH65OV4TfvZqrv+N+05E
UVT8BKz0U1pI5oSUNhcmFpcGZ337XcIwjLFw13C9YdSaqrM3M8DXfp6rGqKd
/Mqkc6TzXsfkIrCmmxgtnZUyRPcuhZjq2AFq9pHtzPme5XuLbLLtyTa2YcTM
0rS0iay1nK0sphDXdAima4YTFEa69PcStC9Icwtl7ORhVhVuNgV8DRmr4jaV
wlz4csefOKN1eUzmXd545A3sr8OYYornu2wtYZzW97SQeTP6wXNjemB2Mgx8
ykFqU79iSlTzASybdHnMsKloh2k/MK9yrGQb2SbqhSwm327YN8lsvSVuPOnE
BAYF5wfdcJBfe8E+CW3HSiRRdsgtW1Hx+nPeOm+sS8OJeOV2htb4ysPEOxjh
B6xe4T7993sRxe+02aN6NCL5FmpSAKDyh/O8FES1ytu83Q9cA1521I9zWh51
ExMTEh85wtYwas/mNRaHqyeEGNQLW6njVvV0WBAj48tNrM3xwd/ebor1Ammf
CcAAwux5dKjNQHskGiXXEtHh6wANHLCBMhrDhvTFvEjbrZeDzX8bNKC0Lb0m
hbRRAGfDz7sSCimLjpugHfpTqLo1ForGyVsnYhU2mTxBn02eCBJJLEmTS/kk
X4UbN5eEH+rLKooZPl9q+AQBVCLHM5s8hNgTSs1YQbi7bGJlkXhExRrsFQZk
rKHeiclIihWKJtujhEO9KM2QhHxgyZE87LTVpYwP4xBZXuf36d6Y1ii2hy4U
O3YjIW6hlLUX6NpCiTqng3j0eEFHW7dHuHPD0BOfASR97YlfURMEICK1wLr7
Mi/lP5JK5ewwSGl/h1avxMv2c7ioq7O/hDoUZrNQPKMbRtR4csCRWJSAoOwp
VGNjlnHipX4+q69OI8XhXmEE4pl8ckhChjy4V9kbc1EAsINVy9x+umsrNH48
bFMjUMVGkpj4DsbT0DzImR7n/XVBizaQDb1MIOitzdxfYUpOykwUAJbMmzSz
gxXEmebsRtPlV5LcZ4Gk6X4g3RfR22CLKjniT18QUpBhunQZ67RFGUD/jn0j
qCIolZwUmamLzzVEi1KN6ezZH3MFURtgl81by5syqNaMR9bZ1GFrWSCb1nHB
4NrfSaSl62V8fFfejAITE2Guoo12PeyZGa7pVPfrpIuoZhISdt56DrLebli8
pYJutjMqCH3B7kcfYhhQ2qx/9YfQMJELrHWCgZAoMIMwfuGsimDE83zyclC5
WWZUcAcFFYDHNgMcwbswBh/tZkJe132t74cigc9nNbXrbnKgQnnFaLt4+AUd
LNDYmeCaDzgImCwpluyanQ9s+6anEVXZTdYOVzlz8vyZo7Nmqv2AZmNwmew9
0/9TKMSECgD5p2nD/NOjKKtdRNiycK17F9wNCWhWFRprCGkRiRudFu757Ye0
5J+O/mEtw+EI2I/f/JbcqklK21nTQEYgEa43hf5ROnQxze3HzpZ1i52GXcsW
LeAlEJPPvRmyoY1SskjgGSAiDglxBFCvUIQDkoSJ83zZad/1SgXBTlLYletM
K5uTjbrAZEzQdVQ3G/08vXGcetL9+SjuarPBeHqDyY01uxZSI2L7XrEegevC
NSt3b5hdPxQx1JP341+cKO0POkrkRKU6CsXQGMB1TRFhNVceJu7nTKPCs/7w
gGw0uB+wd3GvA+CqgrlzgoznitQVZv+PNZ8bh5GsVruNKR4gklq9rXcpwx3j
gkWSszszcS+FuYJzbSkgN9kBj/HMLqDXxV/xKLr3IhmIXr9vyF+ofrw+akD4
FA77a8Srp6/uwDI/bvBv3eI+8KN2ZWGwPIr45SavM8yV9gee37pdlx4iGiN6
QgQow63GfxFhZohbFJHSlYDp2C/0vSlWFC2crM+Mofd0bayszRC0ukF/AfZs
688zJSv3vXZhtKiLdPUSizcRa+Kn9PGSamMhjn8sxolYYnpF5mHtauMIlncC
61OMw5Xmt+piKBcU6TLzqEbmQOj4/wH5lbZOKumAgQLuwt6SOx8cDRSX6doA
X2d+XwjSHaiekvKPzIdutLvaMBpaklB4qd6Jrj1FuczEewR+1QLzMdGGOr6V
LEmI/q/uDCzlBsfGOdgKsBgCYGb1t9iyN5SRmexTuTVF0we6+HqWObVag3CH
uzVIULcEdG3ET50cX16ziu2hwZAaqRVZddDCclaEnYLdlpwVGUWYFzsdeeLd
BUhaEp2MPxWbybzN0X6vc6hK17ITqGlrvrEmlNdnyLzGqQqE5pyG9PcSmo3d
l5OZg99pDFXeADorVbb3oQp3zxV39adeBwBaJ+8M3x63iGhVuzj6FX8xJAS4
13hu/x9mc4qCFFdAcsHH4Q5tTLx9qAPhI//vTyLqHqNHVsZL/Th0duclkNOX
zNlrCeZSIM84sn0VvhjW5aRQ8V3oK/9cT5yh0Lq5BIZS0ljnTuT0E6BztTSQ
V+DkiQYnEMNvw+36GKjRlU5RCGJ9YM2fea+B3Ih3ZskBQIkLQZu/fsk/3McD
3Ha0PMoXvun4kczypZBzNHFsWsJ9UiG7cG/9klGEe5C+dLPy/hToyAdiyFgj
LtovFf70ofpFntszEaAZctqDZRo7W2L4T+XYlUezOdNhLoT0ia6aelt34f1r
cZ2eb4TvziglwgkNSOoCyivTQ7lq0t4BssiNej/x0vqpVLGS89GyehYVPeGL
2ufWNcErxzcjP8LjacX9e2cUUpywVWgg85BPXrcEuNFlZLxrBSXxeJsqfRIB
gLtfFY8tPtogf862ohIYmnHX9GUpuXWEhqWHzFyMVg7yP0uGQCZzuFI6aoRn
OzuJlo2GlYbvaWulM/Pvw31oIkFoOttnd38s3gf/CzClqOKOtZ427tjTWcUU
hx4WD71PCWdQ4iZfZx0/4gBgpgih5kh7xSeCZnDoxNhRRhl49mFb08xvHIVQ
F2zOOfTLxVXoD5Z7YZhj5i/Gunc2W70FKRd+ZdRCaJxGEX8COYVrYEIKfqrI
4DKx2TmbjvKmUp78Ky/wqmRnv9XLoVbRCbMGYpVnLsHp3rDNPPBvyLydvD+J
yijjfjGEehkqu1RQwq0Z8WYhzzB8Lg3zGTyy+aG6mAxJG1Gb3MYBABzW5gbT
T+9FsXHG7AUK9r4qo5PtnCU2/XLV33VXQEGP5YAqgTeY1qwf6ICAANkunGPY
I5sD7i0fjw3CiJnVpGBaab04vFoXEbxiVe2PFKTWbwZzn6YkADoOndyMKEus
EhpfyQYJAqucJR/7xf2qWYlOFb2yhV9H/q2XliwKzuCeGJpKZpl/gjUFOXOJ
JMdVYJQaqW+MvFUr+zVgMBCXE0DNeUeZC9T3ZW1LnuNTiQSTnf7T8i6c7QHm
oZ/VcQpJ38BtDJVzNhQ3espVQIY3HPQMCe94tj03JnRaZI9q5AKCGepDoXbR
wduDP/7G/6mbeNWOoR3Msb+oPHX7/gj+7P+95zHg8t94cHgAICawW2mrpuor
R2MEulDyiapGKGKdYP4xbxxTHxNPyOvOsC5q3KYaQyFzbB31UlGMshZN4krn
AdJfFsoCyg8Ev5qhtkmcq2tIa6BwlmspxIrKQcq9+suZfyw4/GvdtW8EnV1s
cU6NDqAMpp37XXpL1zbk5BMgLdc4wuUzuWGbhTvo8L79XLc4at7zd/ae9er4
2nkst0ZqgxlytlPBS2JQ16QvRII2B65Ov76TQH2DigEtFquddnMpNB7wkA1u
8gCMGZdXXpjjmp83szaihnEoxEO+nC/52INgT+PWYRlpz01yuzuEoIaW3Sr3
PuKL+W96Xqx8AHYMJ9b4wN9QFlk7SmiMXl8wmTb7YhGRlvw8W25JrDcaBWTl
ggUjr6/+qoXfQ0ypxEErOk/nDTz8vHVaSJBRP+4HXCE+xvuaKP9c5Kjn+oaV
EA/4dhoppovl4nnSNIccYqvhmkY6SAHylKSrCG0K1O9GQy0ujBOAbzr3scnE
hthr2HZ+8DHVO/zlbEe0QJqxg1w2VyrvHeYlv2Gp78osY15vF2EPiAFLM5Om
vWXuO3yyyGkFHZFoSf9ob9qw2oXu9/3iTZsUDadQH3ltAiMiVHEBh/5AwerM
yj6+8R6NcBqhaY0jkS5T/Sp066LQbQdD1O3txtFLdUmrK8oQyhzRiggbany0
bhRHGzz2P59NbWlSR10yawY4QRIw+RvbsI6ZElG8MgAZlkKlNAMPeykl0YcU
pjr9zL9L3vJYfMPzDWbI4DazhmUpIoiH3leByPtYJKtMD8dvQtxlopbhZhfD
YRXyRaJj1DGfFugUzHd4pUlxnlZqWLkuorj+1BdDCR0oImYtcVmkVHL8fbyZ
oGQKNkOEqz0YC6PcbMBrv/jDvAIhebXbuyQHEDttgplhHV93Ojr9pcyIrs/J
RgmfCK+7Dw13GZhoMkmWRpl5B2YLcpVrFZ/Hkrxw8XGbKK8Ca1oH8Ichmmwn
p28xjNADfs6JQtg1do8zH442Fqu69rOaVlIrcubsK6I9glbsrx+fstMRjl+k
pcptvKWul5XG61M/kXvXiE7qrn+7h0FqZjRG2djcVrx+XlDESBsv6u6fXpAj
AYoq4ZYfNsjt2cc6/wJ/J0gqciMlQNvFoJW2iRV2P49ILdlC9O19bbHMc7zo
1xCBzUtyUc3scRcdc3hbaEHq10wAYt1/gNlQBXJbr04NoO67x1L/jUgpny3E
mg9qnQ6a0B8wkK4mB7EJX2hDTzawOfbYvGKNQXKto3eaFM3nY4FUOAckL/gu
2bCuH+s1jsXzoCGCnx9mIxNQrjiKqBA/srXvtSzJts82kPphP0FsfRm9CvYH
46FcfEAZOngzNagrWtROVTGgDcws1qsxbBODi+Epbb1jB70bCIDnyoBZLcS0
R1fAlMuLZIz3m6zRuv2GilcCVW34OCet2glBd9Zmu28f2/N8iWjhC1/7sWt2
KAsknanQJ6rmWjOz4tHIIINoGWa23yPxVq7I9PhS3QfhrBNkampO7o7ajewg
34ub8GUU6859d8V20PBZWgy/eI21c2Eacde7M5DxILXdUzK7mi6BYQNKhZNP
+TV8TZamBVead76HSZeTE8ofF5Fug78eZXOvWX+ptkFryDxN1DTUZj6acyDQ
HGU667mOSGqYbeu7ysA0+PgsCBgVwOh7yDc8BckBe7mnMB0OWZUEZ+s4/SN3
NI3c3PE9DiAJ/wFuGSWZ3woFqgP4x30g4AzwU5f0mzwoYIBMMW/j+eNz3xk2
bapk5s3MHXmxWFlsMTUV7L6YExnVUKxuVfQ/QIH76eRMG2tpVXV4Y6Q4Wju2
YC7ZMi/Z+y3Uj+l0Pokbw5lTzTr0vgRaOtskX2LleCHsnGYxgbHrGXeT4TEe
cyGlg0OJjdiUx5aUcQOU+Al3+vAcRrmInYw6AcbeS6RR1aqPBOWltEKxVjbr
HUed9Lg/MOTgfGb/NPu/Ude/2bxpB2NlwdMU8N1uFU0XuAXONY64Z1lD1MyG
MEUIJtd81ELOjiJ36IO+tx3QS1qRp4lHC2mK+XG4tS9s7vvWxD9Fmj+AVoB6
ALDViX+g0RzZFkzZxAvfZF4IF5Hmyut+OG5E8LvikFrOluYgYpVwB2UaxJVV
IbGDlMw+J4DcOfN19+Xg4WM9n6keKMGnJ1N6mY1TOxnV0rLd9s9LXlxfkMQ0
/8tw+IxGBpkNOtbu+xjw+RD/BmXvb4IlUltIi/UxGcMXRZK02665Y8HHduMi
+RHMIJSRl0nBynUsVHAaVNsSRy6jzS8knt2LGadXxdP9B1j1Tm5PfVRqcciz
qwqVAOfiC3ocQCsEulFZlLRiOBd1t5IOZrddM1bXpoVpDwgzTu6Q0e51cnol
AbDlPFhZB0FwQYeQ5nW5OzfYmDYDJSSKTag/7OYLPpeo76VldBzetnWQYppk
8qJ3Cnu26/+aWdNEYKDYCwnfcqYTrk/zkO4rxje9Emm2PX2ysmpKEbmo4jKS
+yx88PHBYi5EOzl7b9wYxR3nymo+ka08Vihcl87pkbQRVelsyyNxtsr7bhPn
jMgWc25JFXvo0XLB7TRcg0i/jUvAo094HRSLlxoMwPIL/0fuBjRpU+CJjykh
AYGCbJn6t9y/J0kFq01n4dTAM/7OdD+DOKmgU4OJ//wJDtHe6JGa9Nng1Sby
GAp8rofFYBMTt7lnh8PPHhJ8gJgAMbuo/i5rLa6laeAWlE2X07iVgxBljuD9
7YAx5sZLcmHDbmxdJ6Uf75Hqusyrc8uzx+sIiSTLaqUCDE11uGClfDjFpDpk
kTXMOsHNChGaE+rLKVjSXABuvqKlZ25UpTWBeCvPwQXsHsYc0SjCEDD4Koq5
g6joGbwCNqjl4EeGED4yEdi3/yw3exzV+4oIBaLeIcgD+jHeM+7iC+KEgGeX
N9A99AFPAYa4HrXDVh1ZvbgvJRnxLJ8yLwA3ZepBOsMLvCHccG55Dcq3culE
l8dbVwNKTsrgvDThi3BWfxYE3fmwzfTVmLRCdSDVthx1v1Ay3QoZAkkOB6zi
urUYUy1Ee+JKFAGJNxTtCE/yDIwEj0xvQG4L/4tA3PQ+0DAsaawn7BGPMiF9
vpT4GTl04MDfqpi2VZHVI65w4GelWcbnsQJL0ct6x0SgbzcerI1/rSXsylBY
xDn1xkkdhwOrXnfA88oFiYOh+3pDiM4iW1/CHn/GialogDvanKTkwahCev6W
5kWmjvzIYWX9VxRdRabJjQVQaYZ1fdR9xKup2+aLBHi/d0Ty+iYXitxu0l8e
XbX9cTh8KOqIGMUkMUl0mQ9xy67RVriCR88NAzwYCiPw9eGduZ+fR0rKioEk
eDXGWBFOzMxk4t3Bs55Qkpfy+a3UuK52w32B0DeCSYsfzKrK6TxDyR3y37bs
Acovp8BMReb1iCJCc9InMAiT293jhCxtU5qVnrpSAskzQvizFzG/zH9UEKq6
XFRdbJk5/TfKWkKLrNxH49XJMl72AwZgsrWr1Lqzw3m4nRqLNAr/BPRzumdY
sOZKvN6sAur/SyFBUfUhKe3rXk8lgV/nkuzIqCldPhirtD2Mvtd2M36gox5D
10fAoRyqwlUtHM4FnPpigISvw20K1HHXCpqZuNkertmPqHfhNO3i2ihSPzQw
4+4ZiUcz/rIWkyoAenmXaeHN45DnvR8s1pjGZLj6kpu42lB+bWSDujueJtZq
IrXlyRmUSmMEDoX7K7G0qKch0oA1Tggd9YRnhrRkZU0JHgu+Rpl8vMB+RCYj
zXcLC8mURx57UTotRtpx/H479wjTcEera6Jh2s5pzTqwt+QDlN/800UR8od+
mJQISK8wKPJF8wMrV23gUiMGkYkFr2EtLBrttWFzR2ofQdroXs6Eevj2w+wg
lUlUavNaW+G00mUttq3/xTM6eea5redu3irtAdLafxJkHhcaJns8RB2AUDG6
4T94B+tUIEWPsT0wZZOPm7YXAP4XMa3dP9wRP+xpZdGImgaH2XZXUZ9BlHpG
gSOhkao/m06+mLt74e/zxmbUiHYWFQLSKGaWhXhZm83g9aNyuGtIoyGmgzCk
vH47jjiIJl4+Lrsr2gR/yTyIyP6vF40KF0uvdvuaqAEKWAzXKtLtkomecVtH
hULLPzyFQO+7TDLuDlqzXs78CvJez64KIDgNaBL5biEzma0y67I7dzIT2c4p
JWjcpO6CcC3wxKtlm0T1RRZ5Kwj7XfJwfnmyhDBJcfTLzWNFpNiJFWCWojic
TwMA4ok0f3wliGRr1eKMppFxmLyuf9YS+2Q8pGiC5bTjrUETti9ndmvS6i1b
mNPw3CGv99CeP0avudpg0vqQsjnfiMyENeyTBhxCiYS0KMbINAiVttZ7QdPE
K19mO1FAtZOmy2ND/uNaeA6FrGKA6lBalyT9zdH1IYpe5v4kwNcGHo1ugwI5
aoOOPRQxDCCdolzmAtu+Gc6EGzks1j8yvTrmgYr5JPpabykyrqwAkMfHcyCR
a2BMu/PuZAKpgefYFID1nPiQeRwVNA/XIwqJ1aPPL3eoRBDi1prMlvZVZGS3
j1o/+i0u0NJgMP6MQjctRquu8Bbj1m7+tmL6Q4ZS/cQoJk0cZOINs1f+9MpV
/786xnKdeRps5y3eb0gXP5v1bq3wjoddenOgOkY1LSUxiO4/RPYbmNalEaH1
VMRP7ou/J3Pd+XgCrflPWpnHn6oYVLoDVtCTuy1aWDpmoAxS27b3c4rDKHCM
TZPgtQme52fZez2j7Nu2G4ELfu0+5OeZLzk1Ackh89KzwYMZbP+TF3ztk07d
lNdUmrJbSK3RtwreAapFiYdr10n9drfpMAyRomKdSOW5j3rkTtLbXDq68cLo
Tfw01HGymEMCDkbEWyT1Fdh74eyqrs21eqBo9FpxC2Zpe87hB+kRVqbDOx+H
krzW6+0QNvSKfjd2MX9hDQGRnJPy9u+CJbzVQbJJwC3VfWQhCwLaIiCSR0CU
jCmOPCHRuVVpnDKvnT7Ci2U5VgxNN6wZus5NKJ4ocwFvdWF0QVud336QuwYs
0Sd3FWonO+4T2vQ+pZcVIAKa7kRAthKI12BePp4ndrXKwvnTd3taeKOaorey
6phwFvuan9bQ+o5HVwJM6ViguGo6vfwz2ipFq7JzDUDJBe/SBHqkQ7T3gLB/
opL39l5uU88DMwWD/JWsSYl/hFYx8w98PDHcv8tbRhF4Oy3yvBqBW0GuoaS3
owXBoOjXkZBawshLsXLmB2xeRqlCUN+y8vJRDEAi394OI0zSL6uKEV78X2+d
BKcIrREuHgvkeIpqMNRlMnW4fNszCNooe2cMMaAnIeuu1yVWdrWRkp/HdR87
IeTxMqjAJVB7gJAbIsOsbe2QQBsJ/JtGGuLJGL4Kzj/t7Lg/yle/hChakeHc
Y8eyRic3cRGf/ApsFkgb3mAXKR6RW8s32RPMhhQWW3gPQInP21OkxzpMYtLS
cp//WWg4K8Mf4504yPn8jP0yeKJeRCAudd89BUiyJHz0bjhdhZzn2Dr5vF71
mb2rixphIBcXZ/2r7sc2OTbup1h0c/Sk9LdZKsY84+rJ2HF1g2e4ipyPdAr4
La5xqoVe69qn7B8yjE9mT1rOj/Cm61uuO7pi+qrVpCxrXsPMsmptY1GgVsXX
QjdGYwxwbQ0S0lQsCbVX8l9+O1TgN1X8AWASp4FOctCRd0PHML6LYYtVCIYG
epijwwr9HD45TclEKAYjvZ6iPt+HfccHrEEk2ZoaWQHZcssBwXvCF6eApDZp
OV3GbLWuWbQBoJiC+QFbBLf2I2hRzlcEAJPwjRqKVv2rcleJsl+QGQs8oyZ+
mhef5RYE6JviKfS0wtT/sxkg1bK/goQL7nLaM4qIjYeWfPSpC+WBWHoxUpDu
isC+7hmSAIvl4lb0dBq0h5IYT5zSCBshP8kI4tYu35SwHqLAloEzTm2eIlqe
BY+ifltDoa9I1ovHVn8Ij6f9Oeny8mYUofI6TmDXsPas7unKAj8UG4NqfAb6
puov5D0PoZYFFtF5QmRo6QYp+QA022BhyVm5Pz3hKrOMisY4XUoeseOkgMoo
LyzGMaPTfdoKu0UWohPfcKAEomJmBWuK3UYJZpWS1e6e2rPTGbsFai9yjUkV
+yMkn9aclS72Iso+0GBaCaff4aashhSgJTxlXs8VmXWw5I/DMr5+MvkRP9qp
I8idWKRBmlrAMkaLvm8dtfgiYXEx20dUZDSVbzYquvlW+Z3hmQbn4nxXoDAs
GGVv9qugKVMYyrqEq3Z+OkovzvpJqZnwKVBWsRrpRMKlVWtGpPT0gB5dTaVV
KzyCQo4JNs1m6pbf4tf7qOMxxstff84f60ry9l/fc0ogRcIlDueKFZQEqNha
3Jp5RFL664DGgO9Fiw/9TEUGl6LzY0YBwp7Q/wf0vCbgUZlwvtlQky22Ci6O
enLHITfE1SEuu04whjwWDJa9AmgG6Z8+VCBZIlqxmpQuDiW7jJhI8P5TfpmU
leC4l9pkgQH3rgb4iE8j0aatoytoMTjZTwUuAwBiXJd2jyIWgL/vJrJzs1U3
s/pP/wOSH0GI1DYhpOIn+ImWCe+3t9wY0R/tw30lMabYrIpdKGX0CHfJfVRe
nQ82bvHltEwMrTfn1U8uw1XkJMGT2lFbQycdMnWwtv6tlbnqOG4NlBz1vBiw
Nd9G2EAxlIXOLhl0stloIY2Ahb4+8q3GPp+OSm11OnBA1SpYosIuctUAfUI2
wRK0coc8yBHpJiV0V4Gmx7E7MFJ0emUibDEGGHTZmNBHogKj6thAnjnBkBNv
DKzMKL7hL/ms/v2PQtk7ed3nOa5XlA6gHSu40W/ERZsEHG5NSs6++cNZY8mb
c71LxemTp87lA2gVFD6JIn8qT0mAPwRIP/x55plKH4OwTL1UQ4ZKpj0yE9g5
IPdg1KZQxDwPA9DhCbUjALnOiR9Z7I2AhRdNeT0tVfEiw5Qu+WFk9n83/7P2
5MHyp66/KZKv74gTe5i+Hhgi+IQSiGBoKJizEp3fDx4lsT3r0UMU7ONwpX05
ONwt+374LKfGiu7zWkDQiW1Mg1GPrRedbFGUNIhkwL9fxHrVLBypTv6oed+b
U4Zbd/nDtsC+6UbxhXcaaojE3osXtTPj1HuJ3Q1WI0h/YbBu15BlVFSwntsi
/IgyERDEWigyrQdD+r4A9//jy5iQ7hRZiyv63bM+zKRrah11tTeiS/e7ZkXa
TdEV64IzNsEVs9MBJWfMqggcqkwSTAaJ7uQL8P8XXlNTMpZv0Fkj+Mbpq/gL
XaxPATgD60zwRDN3T6lixqYyaguWpRYd+hjqxyk8dQiwBKv0jqaeyAcQ8Zl4
VB63BWZGmc/rv0PlwMqgvHYseV1KCYEHaaFjQlmkRz6/SkCxxqdkKP6M+3ew
bpgX53+tkKDUd3/mgUxPz/LiUBK42GLW3V4ynzeANGDKKg1+LsYBdTLIiwnq
zVnGNRPuWzIZRjx0Jhv8SToY0gGKnJzEcUU1VM0m/NGU12/1/qD3kfS/4UHK
PMG5zXzURHkqWrkzXk05D78dDBuXLny3e+W1YEkMUWYFcyili719D8U9fO7x
ZyIsGnFEtuYsUJD2Kz4SJxh0FnVh3bbwEfW5ppfzNYZ9Y6Rq4JzYcFaRNlO8
vchOdqrvEHi1B+917zKVtf7e/xtEi9OVd8n403+cSBnz8mJBMt3zTh3Hnp9D
yLzXt8eAKa5pUdjlBq3eqOfDvJtYSjMc0lJW+fFcN7iCNI6OneJToK8lzG6k
rbGPH01IwUD4afd6SVm7TqOwIiRStYhPkxvrr728C3mPaMMrOOqTy4Oj0xGH
6owpTF/mCPjFXDPKf34qDH2SP0dj8LNLjhRQbgEFe1l+6xta8tMWz98yQIcq
/x0uBIyVE6OITFUg69LmOmWlv11A5texWPL0PRuvf631sx3C1m8QFMCyWgBQ
35o+UqNCZe3e6FGSakAUohk4K0O/AdmxKid+eQBRiWTWmENlAgZVBKDcfaW2
tu33kCafFTRH5Ebnr/uIBTz8FQDkuaaQz7a38wFhThHr43/9yjhYTe72/4OQ
H4CHki80Q2KALraDUHm/VO4dDcy7DdK3t+JPd/o0MgM2pM+XdruQ1ClqDHTn
w+EWJDWrBfn38wBTw/v9rwSCYPjulgDu/2kzbJlZkvKIsEqmIjSaqZIkPDvc
7nbNETa7S7cKdnB0/8tsN8ViI9Woh0buZCTZ0bvMHu3lyHooxj+0ngZs1hoi
FXcdzOUa4XUd/2AosR3z9WvOT+H7knxVHwN68Rp7EuWdz6JXeOSS+K786IsP
v/rQsjaknyCs6g2qaKrU1MIUYjXXyZ4MDB5bwCQUDjKAgaz556TTgiPheXg7
O6/V64VrvNkqJbXXC8niFqkpr69tBy3j37nvrDBpG6W1wKjl+DtDYv13IR1L
JuV6q996lPQ7sJoSeuvHgEsgLGI2Wt2chScs0xx1y0DHft9NvcxKTcntgNSF
P5jnNvAXLFVj0v+J6ogiaFx5cjec5IPIaXgLlKcVY+SL0l92xEYbUsAsJjrq
4xYovthOIWR2T3lRnI2lJgvdT9PFBfvMV40YuEzHr4chBM2WJZwjFSn8TqKD
0sD3vqG/dR8XK1T9r8PsO3zc8jCn01o8CYBSyCbzTEHoe8m90o8KQVsYIXGE
0nApR+3TFGn5IHdOd5tnbPLFj0rd7bRBvg8PPm26QUTLAgjWsCVYNU2M9j2A
SM93lWFpPDW4EuOGtT/3+OtSZecChbBidDN2d8sEa/EQye6rx+ezTtG4NVHI
zaHaNC70UCv0FNp5INXiP2YBYZgS6btr5VJW6Zh/V9V8u0gjzi5B631OUg9x
WvNB1txyj6dEChJ5ag3cOSqxyOSe8+2v7mJ/P9wwOJcn5nB67Yrq4STULt2b
+FeR0IqCZT91d82WmH8ItGtnWpnAMKBdIf8rXGeyXJEy6RqtMLzJH8Jye5KW
2Y8dx3G3uilR0Bf0Vc1I2akdqNVtYvXKcoaT1wwcEjM4Mn0G+9+1sTUj3PiT
0oWOUI6zcbJSz3pHXJS/EECt0jRbR5PegZeToDkvqZQfw4jWXllZKamxrs9v
2NIyfkN0SZS0pVyXV1c6zI1132QDTJCoWDl1/XIV4HzErKAtzwZDWYya5dis
BaYtFuoLWA9+FpX4yUNFqQFOdwJRttyR5vy1QZ7p9RxHQdF8S6D8sbXNovzF
NfmBKGQVWGrfcEL8E6amzI/7sexa+rteMuulLQ3vmD2SzOodIK1CI8Rr/2Bm
hhuqlX/+Hg2s7t8FFmfcWQpxJN31KIbwEsgqDnIUS9sJy8ZwqmN27klOhAX/
vqeas6tdWfbV7fCJX1LYXuhjEaSI5wAC7OAxLtEnRleblHNK5la7zWhLSLDc
RRQsSaPaGK93drNKDvxyM0KVjQbZZcaq1qSOiVYcf/LaI92BQMcZOtj5X56n
lJtcTnRPfBPWbIq5wpNC/52KOrILpb6hQQfB5+Qix1Hitkzy43F4InZ5jWD8
PhmXrSFfjm39gvwp6y/tUxEb7VPZDgAHHm3f6aXMzAiZjakp8f6DIoXh2r1p
4onUFBKzf8VSMSLjNlwe9yEaM7SLQLANaAn7tmTwoaXrFtLgUXe0AdwDTMHu
lecgP+A2tJxyjNk3/OaesyZL9MStoiPxdUlvfUhy3kDCYfp55UnVBgI1kL04
HSPD3Pk9dlJFNItNzO9IMsSKNs8FtElU5XuEbuRWVBEw9i/cG3XxgyU3XbxP
VaUQyXVaNl9eeVHmeMOubw+eQnAzzjaBV2hKgAU9TH4Trn8/8zae5SZ7drv9
TaK4hq9rp+mOMDGITJzE0MNRlwwcQTC/UJlvPJtJWVGGb1CUK7kbJJFV4YtL
rRVCxyy69hLirMaQr6HIFn2Qu6DwNt8rDU1Iy7yy2ydBtelk3uaXLgYrFiDL
lOR0ZST/1O37slPtybM3m8AZX5b13U0UL7SPa0J9KuSL9sSOthAt+wF8Nb/3
eWj4ubR6qsHkJk6hAoMZj+V/oKUkGCDmJAq6V3xp5D8qemr2dp2IJXwnB6hb
Uo1NLOxdAEUCpp2pPXKOSnKuDRsdAqm2y23fsSB8zKUM2uXUKyEMohSk8B+4
n9cotRWNOcStbVeQ1Z31Zd9ipLqfQsgFTj6SZeFL3Y5ZHy2QhLJSKkQ+e4oC
Jbp8fw34UuQZDWFN3zlI044PfzGi/5SBWaqAw+WL0Cmt1dkf2RQz1RHj4KCD
1Onf2FsHinET/22Rs7MFRMbvLg1tFyjXvW065N5rBJrxxmJBz5rKeXAl+O7G
uimqWZ6Q7v+zjJC+IXpurstlWs+uq61o4XEZqyhwsNWctAnq/FdqoMsPqqKu
I5/i6uBArfa1T9kff1Axy9KgZ2qtOYihEsB/D54zCLEx3QBwrYPGYtubnJbL
YR9LBKnJAPOy4q0C+UTkt7/9Ui31wYOBfZt7N225NVbSZ/QJCtYuxs0/r/dy
N5ajWUrxHhLxhPchZm8kCaSssyRMui/rUmNTvUQ8y6IqO1tLhemsHBG6VUlR
jfmAlYRZvAb0nCxfafJdOIEsKYK86s5r/0bkRapm/M80yMBqgqsB6V1Guf+T
UzHOXsJQ4SlUu+rAf0Z6jXOeoLrPSadBBP2o1Y71ov5CXJjLXpesag6mnnGD
dTeNk5u6fHJHkHqGoYLKPucmhj1HkrAZdpz57AFqrpUlT/hYa2OhyIbFc+3P
xztSHLXwQs6TF018HvVROJXev/siYeTWfWuCGZvBzsQmA+gt94IAt2hq2Xt0
3gGIsvsoonVlaxGF1uA0Hw5UXYKRBHRlXp06UUJEoU+7jZJwKzm+xnUUsUoE
swgq8rfnUfiZkeDs1aKErHW5HzsLvQK1Pe7RrFj3EVoVXObOMstQxY9QtHGN
CJBf42YN1rYN/p4rH+a5nLoSzEsx5G7779m3SbYvOlx2/IWdMAkkDz0h/Xzc
dC35ImcRWpZndMwri/p+DPasSr3xcuFe1DqTdG9EQxdGbkL8z+1+MKksDzZ9
LjiUG+bZ7qdyJRiz0TKGvopE+hDSTVgAUXBehrCJrNStjxLbCM2vcJNozYmI
acnhPegPCFg2aJFLjJ1FTYqcVVqW3LXr67/zOrzYw6S5uchfsSpNoRpK5e4F
/18LKWpMy+a3M4nh+VlBi13LsCO7VSDpcK328WQgQOpWCYKXXeQFP/xOJuAc
BrDqWFjv4kqgz6WaBPbbLUDAB2ZfwutFU3x2mHtzbpqMCjGWEpcmeZ+21BdG
wClU2DnyAqdeYPD2wpx8shd5IYq2sp36GvdFRsEJQ4i162UOJ8anrD9JPYnZ
t3NMmpiIbChDi4ZWEc6f/CxSZ6XBaZeCQ1RoXBh/c/L24uZNri21o3NWPza+
CMcAqzkmsHGb+qyA7WOx0pNGiQIJY7YXgerj7Sjm4Dr7PjOLsNMJr9WYaWkx
ucElIbUuRMTa7f9YWgllKy0sCQmMLrfRIbN/BI/RPzsHnbYpbQDXv5aUrCPI
5Kj1hwmr6zJRWVoK5WMUJkxgYRtjdf0z+ksWvTJfDTeOEpBwOsTD2zi9Ce0a
giCx7t5IOIrED5HiH9I3zsSExmlt77TDP/+ARvfXZCefWaARDAjSOAdoDmwG
qS+6Di1Es5XUF8w+35v2Zcl2AfR6YkekwOVfFz37eJ6SXOTfqwHXvEltnTHT
TlR1XMcTitN8EAx/EP5xlWkcX/Ty/z5O+5fDXKDb0Otuank0HVaxdFYkBR2o
aN6nSEvNDLDC9WmFQRwT2cCKvxaoNTiKSJYuN6YcIONIl2JPZIQiWlsz5XJ2
+yT2kWSa4f0rPN4+T4Nh0l0rSnbSTOK3B2sC9Qn+79jepJFEiDoUOSmEIvdf
C2ttH9IcJPTztP54NVHHa9lCnaZTEQqd+GJtYPEY4gNihhXJePT9iGzr5uxv
3TP5ophXC2ClbcxUOHNHvLmz33CsTtCL+twVJraBe6KSJD+z8DL47saSUU35
7okhm59niVHqvjDZbOsSJHOjvBybM7Ob2y/2kCtnoCt0AleRvbdkg/Jq+MZY
uxJ+5Xh3sOrKj3QcLt5qkThWPyHDqEuSd3T5KPnwrX4q6rDYUms8WfoWHsEf
0lKZwv+s2U7AhfdIL6Xn9DDCIs/4PIKux/vHIPWH/ZUvdGKU3nXBbHN3FIQv
duT4C5ZOBC2JhrcwanBrxReWOehsRjkis3/NOLNEJ8guGGgkbq4JK0wgFVpO
/mf9NRTH2mzrcohi7S/bcsPElZQvsFVm8f/SCcuTqWC5mSvdRnZAtT8hUnqk
FBoHjnw3WB+LNQImjYH/yosGanHNbcq//nvDZrmh9irmT6IUu5EWmFvwNP9P
jCm0kln9IjOa2No3TGA377mSjnJe7gh2RPwhgJwLM31a2wA6B7MYj5eTQG5S
yp9FjaidoFVZn0x/FaSIZXaFmDbkDCcILYgRbWY2gxz+j/Xzx8oN5UJOHhz4
Hfn6kh7ECUtiDm/gkPpYtKq9IGlQo66B/Ib9uyISFUU8S8YqwwBHv4A3kfDn
XpuPwHNePaOrxnQvJqEE9UQy9FJQCXzccUVCmYQUGWcM+AmlFLPbhEqU6j8a
egOFfTlJLwnlczEnb44hh9P5YT4pYDnSGgl9VFTvLG8O2d67fhutG3mx+25c
gNvQrd5Qvnp6iPZz5PPeqMCBB06aqjhQqA0mtI+KJZupR/SZVQ9uubbS7J1d
Rot2YuxUtgUdEDlkJ/2wnT2T/qY9a+gkmTm6nqzU1ZNJtri71h8s6MQGemQn
XFA8jDf/FUAlnZDhMysRFOuUYtNbtn4bv9zOelfwM1E4XQMNZwWlPXuTh55Y
JTqcAiQ2REdTCz3ALwnhHq43A68x7aGyxtvZXTzVQ/WRtSD/Ge5l6Zzm/YFT
wvB4fLTizYgsOfcmB+HzoUXISG7y1EkrmQP4miltf3B+FfTKx8TrnJVbVwvq
RunFTLAPTRsRLw2kFQh+C0wZoZtx14C2b3Y3LSNOU/H5gko4ikG+FlNOeR1M
Q+1jhlo3C5lAfIu8ocBKODJqOOjXIwypZp6AtLOc4kjgPNJzWHN0YePMx3iV
AY6WtEkbl0uT79ki4aKaMN1UuLOffIC3Vqoj3i3OUEWmyZjW7TVpZbp6XII/
E1VVQNcsZbhm28b4Azl44H69Rt0E0B6wd94y9kGunhO/08WOb3fUGVpqEmv2
zIRLMFSd2IT8Lhm30ln/92+BBlt2S906Dn6D9QsO89ne8JbYPaMsE+nUmrJc
w5CX2zqzj5TrUIcK92XZhrvp57m5L2qK2IWT1CogKLAlzLhHyVcXMG5ooEKh
h2h+1NVHLagZLySg13DXXfarjFU7O1pZiMEm1THEYus4vVLLGzyWPB71bHNE
L9ehzNJwqMvJ3U9Zeg12z2h2V3Br6W6YEVNkCOU4f5TXKBw/2gmivuIArsub
NdD7//rhWX4ZoL2A+0VNQ46g9Q/olM2bL5nrY5LIhtxUQHDVSBfgrZm8Ooyp
12S8MAyI/qHkupiE76QojuYNHatelUK7Kd0zA3vHQU8xFOSQTHjr4N4nRsdL
hHI3KclVEmTdndOVvkyyeyPmYotCUvq3PuZBKHXgxsWN1Uk1RKf/cTietl+/
btwC1eSzeW8qMwgjzyh2iZDH6OBU/sr6nskYkoXqgMvGsXISPxEBSNtlFLx6
RFrQydWoW3j+VFIhc2gKkHdeTRGOvaxWLYrpoWV/8DDIVqpOf1w/SvqEuqyK
VYcjGyKSJ79Yelj4hzpLZNBfBA6OSIQyoq9KARCsZyeB2gzVGitvjYAdyAR+
LdkMaXrdAw2J58Hbr86nX4ybTTozxvwAO8kAzLo6JrgukgXXXOzXfkZaur15
rfHggBTF6R27ztRUWrFRLNLtu3MlV3zK3d4Lvt/7GxoDHJJIaASrw/XNJwSK
6zZEi6+IcxIjl9NkGBttWn6JRo1wWibJ+OrNqij70mgMSsLplZxm9boO+Vdt
6etEj1KZenDSDlHknDZTn79OLd9N0Tu6Lx7k9YvY42caZfaHEm46eskv2gkz
u9nXv88R/NiBK57z7G9/AzMZKDTnh67kOSY68QuH615kzx5QNfm1Jxr9GYht
ZI/1MjuAi2dUptpaDWg+6/JLThtk8Q976mIgg1tvFjz6gpI77O77XSSYGQ19
gHW+xKQ4vZxNDsgEKjIySinpHv8eLfuoEqYx2BHnuIonBg1EVDM7rifgMhos
zcglN4Ml1YhGBuc6HSP5pRVa+YQj4QSaLRbIXpue4mxJQtfCl36WbctW0T24
elqmJtJ5QYybemyD3s6YvbHK1TS+AznZfs0Zd+uRypq5cR0dFBTPk3R8qFIk
Dx9Wt5W1cH6DnGZzCSZdrOTOeyThP6Snjzm2wzgozErULwUtKmuBEnkMcj0f
P+4C/Mqs5tg1WpFHPBZ2Aaevo7gQYeltemoRDE5PfEv6e+V4IOIUOouuuiBG
WodLQNzrREQbaD2Lid5IMPnV58zsq+9RufhRoe48p7//GTcod2317+bI8bQa
QNsK5XV60+jvHARJKwyyNRZNknggT0TtYYhcKBdJPocdUlW2PSPDQ5GVbLHj
vz0zPJtT29j8tCxGf36SdAq/K2BplkN840bXmaoTbHKo3Cxt8MruQ18khkz+
Py+HMfM2QZf15cIJyL/6464AFWWDNzbb1d2vaRw2lCaqgZrSNdbtKBBUdLFp
9VQDLBNmpGnMbDKCLpBMNkpt9RKo00ODmRXG/tjsn6e9OXzzRBpTOps84roL
8LXDeatOfNuevJN+vn6RZqRp6untxc9g7EOAW/xrwJMUBKxBoW2erBmGKtg5
OzCePm5FQhBXeV3YdfAI4+j3RUZYBqUX29r/pb7yTnBz74WeDrKquKFpPL56
NiweOfy6CEq2z4pfkRoNKw6pemJjw0kMncfKX17Mq4/FfrFUWdWkIjz2tabQ
27zhD/ghrxW3dU2U2Wvy6orWClrkOyb28cBsyCS27ipaDNM9cywmmDGcR9Jo
BU/rYNeLuZHfBvAd9EcpLbkZLTzWQbRMEdXhPowzjwdFyXhk5Lzmojvp2Gqi
1sQTiJ/PO1FaY7HeeAVt45mZare4xYsSJN7yRpW/WGTMuEBwFGeKNbAT4dAP
88UtbcQo9iifk77WZY16GqXzQXB1sqI1gG61lSqs+T8aE2FpoHl0eKkzL46l
Y8Rjd1Q9GEnqWGB6nZ04RzcjDlq5wnn0nTjH8+vv5bi9BvQfEEINMsWupV8c
rhCe0sXLIyHS1dKTOGhwvknYx31I29ceYx/NwDeGFhA7O8wBdEsT97gBUf1u
6pmOGmenERu6C7gPvXsuvWGZkamyReKkVFODNjlCzrC3styDxHED1hsFSA1y
aISrchlS/U1SVScvXetZ/P3ZWMPALKhPzMm12g7sifxFiL5h1sEFhNb0RfRw
ynna8uVnoKgnWFbzx2bB9QcSlrFuDFvAoZTBXgowo3ehDSqEqMBaXNTCaBXg
WINX+8CsWIYwCzy8LxYUmtmQbTomtJ8VfIjTmnQDlBsnqR4jnPalWyg9roAP
qmE2ifEk6smofRLjGFiOs6Q/J3wIX6yC3ns2yWhwSyDmb0kOk3FQZgFEY/Fm
B9AeI1iU0Rfn3XPfyEdHQq+tbgiyd6UkK9R4kzu0Z5o/KFbf66X00FKZeIzQ
Y6MnjV9NwAwFFC8NgsTLZR8gCyJ39wqf8pcfIjjLyHCyR0gBb+8YgStvlj3E
xI3leMT397dK9XgO26JvuKthK124Kl4gRD4Pj9IGESPBIrbSErV2lECKXQxQ
puiQWl/ezvcZxrvKXnnLGf3X2FxQUOjp7dP3B504UjhR2u5n+Ekso7WF5P9d
7v9N+osIWRqbYkU1FzguS5INQUs152isxoJ+/pP9zSJwYtv/2jzwcbGp8HCZ
VBhCeWeyp9ALW2EfsUmUE95FSMp4ytmsGAd+2LlWxNe85aOrPJJKlcxRoSQL
ndj27kLMwkw5IleMSGF2/l6ljjkhGof8I4PS/W4QeLKIzQEH2q4gdIJVoSgS
+3bZbsdjYJmIvuGLNFG3Yp84LREbdnkoldy0Cd7eawMez/B2ccsAhX1kkhAt
TIalXEkTMFHiBiR39tZpiUKiuV48mjKraBB8ocHKa/2fEsGcWYfSW9tDXvPU
VMMQtIAWXDfqfmNMl54GCOxLIhQ21KawiEMehysP/UzouCnGrXAlhrCPWWEg
RTpJlbMhIuyddW+a4r+N0dcvTg8JLqO312Q4LDGDV1Nl5ks50JKrLLwjI8SK
jaeQrx3Wz9rBhKNcImraDDOdZfey8SmLtjO5pCBL5UJ4iJ4N2mItAcxS7e+K
Q9vaSsS+7s7rePicUAErAFzH5w5KzfaNXQuEqAOTlI/72Sw0uy2/x8MnoJfg
LBorlVhScHRQpeVf0UaTNAbQtk6xYR8xAshkjvxmg/YTMTZiKg9LYSojvA/+
Fgsz2eSgABAl1xwrj/ZBi/Qi7va0guzJli+f9B6B/ISuLMLN810uqN+o/wno
BteGp+lU1CtN62RKoH4dZWG2pxEXDUtlaXTEHEhweK2OiUkk/tHBEOiHWeOR
OJpOHdKWrK+IGFwjZS5o6MMyhhd2BsaAZtlkb9chxtLFLe7dNmOmupeOTPi2
/W1y4+w4NFvjkFZGxVj/+GPjJUJAeu9PZcA4hc4WBTzwp8Y49kfsCA7S65FR
PgRO1wird6fTlF4YAh8cKdFkQ3Uud/kXFjGxNKgwCG8IEpXjn+RrXw4dghwE
gfgSl0Es88eRBtySLzjSJZhxMjnPF3EDSwhzOd17H0UicDnOm6UX4WAEs+Gw
Br+wfR4q6zDXr51PO+PKlxG1BsSzzcwZg4y6uMleL3GtkMkUq8YPRX7gIBQE
0yk1SDW51/nqZHyZIceuzL2LexesNsAY03IWBN8hDVyTGjAgy0GKfK72/DOq
Z5VndWTUNFs3OJpLn8EexltY+HHuEQIOEXKoYCEHpzBoiZ4cEsJxVjfA4Bmj
341dPb9Ga3EICaW9Qj4myyV1clxmD3KGa0Cs0XqD4U2Mc+3tZGQnCntdNH09
ORmO1BpZlXZbVJA/xNarw3lbISZh5ZLmm3F/7WqdRED+oYwDJNpUptnnfysf
sqNYCDsRj0QyrkdGNMxuPBgJhOd3/ibTLflvRL5gZzLXMH4w4J9Zi3NNXIxm
sdEJnV854Jrg5JUp7zoHxxdoD0aZ93GHecnT7AOdZIjmiC6Q0/FAtpnu/V46
CsGbAE4i/K2YQuDBkfJK8Zz3pk4A4RRXNJldgSuzisnSL0OGiOAOmVyPD1/M
OxTEIY3T8v8dWKIpz4qJ1b0ev2CesPvCBGHcVxnpa3u7Z6CES9OotGmpFLq7
RLDxk925apuo8swW+7ZKUNqGbzfFiKupC3MbN44SNcfoWCZm7xVXUBBVYo+i
seBEizRCxmOVoME/cuWL5Uy5KWQWF2en9aBWC9YOdyXf+iS1xCksZSsLlFkm
KHkILv/HOHcREDtfeFQ8S5ppYwwI6cDbRNSjSNrkF7fIkrhGD2dxC2T3LIHH
zyvg2KVnUQT5kGRH29bdXDdy4O+c8a1tM9iJH0Zrmcj5rrhhJYfakCQVi3Wv
0ZjUMNah/0KMlqCFPZ6LoXunpMx/c/KkJwVlNt85FJB445VtznyyeHSqkHbX
AZ6sw/EbOihXVK9r7U7IVBp+4VU3yFnWsx+cnvAshW64jjBgGtdXt7UOnLKJ
8rjmIvhI77rAMx0etoOG65s/MMrnWYEtXKGtqYW1d0VPw3KaksFwFlwxwi0w
liKfxXdW7u3MkZ6C+sbkvVf/YTsd/7FeYwWcZdL4adic2SqrBeaZFeHtABga
60cohFSr8Gc2agp1meZEKKNnnaOeRvNIVpedY2cC+AVE810YLSgcpXmF5fAc
UpTQr2H0QW8Sjw0sdF/5Mzn8nW1trs/SMXggJC+l6i3UcmiZv/uL68zEGtIv
A+ViNNzVwSFqAKdPnCn7yTaxFrqXukgGr67bn1ZhuXDGWc4TMPju5UjNAbZ6
G9EJBfzePbtbOxcZqLJpqYbAyExL9vqnaVv3kOYrKCD+kizUe49rH27u5zeu
eWNdf2cQGuysWle/nO2SwN/2a1pIK0CDUPU1YF/mg283/lpgrYVcOaaSvWPk
bF1U/3Xkz7pFLIGkwyyRSQFr68ta0mU5KfVzXMGnWmaASWE1QTPqbsxEU4kO
uoltKK7Jw4vAODPv4BNO7KgQXj/gMQXgyP26wAhtn/hPj9irPowvHxRipr8C
r9RiOT4N7GF3AxZIfsKhSLpvADrf2dmxXsrDRzHp65sL5r4CL9SA9Uy9GB4a
tm/NDyrutSJwb80tmr/72lY2rVJzPviZX72sdpqMvuLjLt+QUKYqLC1rXmrt
vtolpDJ3W9hoHc5SFY6A4hUWzl7/n1iVsg5Y+XcX3zsz8+cIXVdxv3Zi95NP
Ks8Cg1kIXd1C1uDmPUy3S4ikQkJNjYVX7FaJ6ZCszSKUaxwI8UeBmPFAUcDH
VyfuKg2DnjLzlO9EwQPfI/1gdrVEJcDWtOLtYbuNVebcT52SOb+4rRXFjsLi
9EG0QSeaEZNbBQ70GNACNl0gmR1zb3frn6cO9x52zaLJQ1WgIl1HlRNzGfpL
EGtC3pJEj6yrxfDcp2UxybKI5YYXz59L/ndAxaoZAFaYBFmnXb+uodBcEJVa
y6pXjemUaQouGVER3VXx/Mt5cHRqYhIfUcjBH6qY2PpjtzXFVgWt/F96K4y1
ZpvPCI6bYTslbn/KCl173VD5H1AdTu9hodso+7FfW71I13BFgke2LqFHyizW
F0ZticNajTe79pA7mUHr3/H0LcI7EEQp3J7KEmuWWrZAZwsgOqFlRQY+tVF1
dgTwBOrJzmjtwi3eKXLTzLGJSnxt7ba4aGsQ9XTX+kDSt9qYpRJZyLxKp+Y3
TjnUsrCmTrXJk2XOaxA8izcHD6YZN35qj7w2a6Ao1BRQKZaB34tj5oRbVHeI
eF+i0AoQRRbLZU/GTrjkONDp87zNFe2GnarXFXTodf4zipcJdTOVzrVzgb8+
xO7pzI5w9We+5dUvSVxk3aPoUiP5kj3YkDPoQRCxm+3K6ihrlVofcewQ0zz/
bLXgf0xtkrIi0l/vkSogHBsSse9xY3f+DHJZg11Y8JnLocZzXr0RL9GhURig
ET45W064zq0nYDI8uspcMRIFVNb8WLDzSEoVkSM3dNHxx+ZZI2qYVvZqzer3
SxEPUF1JIfq0onsnMAOgz88NA6VWanG29P882oyvN1kgIBEUavv0cCTKZqCj
b5ofR6WDSNeBglQZ6qpRUZ+9dqPh37uvzimCej7pmPxJ5xWox4K0ZTklMdye
ZxyYIrjZd86Qe6QckqRDOCVMkdOTTDptSR+JBwe1vw3+wXMMUDkfmRei6Rh8
3/aIZmsmPkXSQSn0y6M51pflvTpET9AYemwtlTQ7iozs0sV6iOMg2xS2mNmf
SX+XIAUsDGe03XWD1F6fZXjGduefoDP1kt/W0zDww9MTLhF4j2ij54Jugou4
2JZsdqFVb14sI9h40NvUOcO/0UIllY4kgiFRKflFECLubOUkktmTBFgmyXfc
SWjojvAqOr/GdlcUQu9iLNfGogQ+RVphDCDYm6V6O3hPR5cXV2N8FGeYafQc
YkR6wvZ7Ma4/MVeC44P0BYEmU/ES+wGJwHyvLTIHRCz6JStb2qN3JnMA4awa
rInbHh+5SYJ9nZwmdPN2fSQR9NmvGvoG+3qQWk8kd3y97EBXcWDWVdItw3iQ
BMbc9rT1KjEfK+yYA4K/sUDog2c/ViRqFXT6LXFxTNyVg82zK85cdCr4B8Md
Cs6Fql5bfwBRuBWlDHL6Mr++NnYzURY2rP1zFBEInN0wrLcaOWkdWhvlrgvf
glYoIFOanoO7NRVMIocaL5qEwC4fyqzjvg4SfL7B4o3FNcR9XhEfcngXkNo4
05fGNc0RTxWLLdrFeRRp/7b1lP1mmQ3bVZkG2zmK2/ABPEHZDOfTyxEmRhF2
dGrRCG7bRbamMbfPrShbVph0gD7/WR/0BRe3qh3WVmF+SO61TWx0LxlKx/y7
Qv6mskH+TME4RHetI2JYvUbHBp39ca1kiQzynuPf2POCFOzZ/5hskk10d78c
m8f/aQ4eHfrro68qUYc19v7ATue+QZtteKYKrzG4YWE7ogtqmeCYsz2V0Ats
SOWJuJNJW/rULHKUBpW3KGegxZw2cijCmO6SMXEsNNMCmPt8ypD3bqyryBxp
lPLzhOzmJZSPdGgL3bGVj0+fQDzIo9Z6ifswzSCHFrMcm/CqQaee3kGDBzeC
SIJY8O15yuPKLP4pRFWAcJnN3k36LyWNAnHTl+YCsvmqOF+qw9FWCkLVOITq
2CmdagfTSWkLZZG/Y+2NuYFNZTmwr0TaPjmguMOiG3+Mja5H8x6KesuzplbV
nkzcLwajB2sTAPcam8hP+XN2DbH3NJOBzs6OoHI8s+PGRsCMYFtNDOCTCfpY
hvLTtj5LSOStvpPtsjDWGMWBhk6bHvX1RnfVg+XiPtZmaXuM1elupyqyAyRQ
skClUQqGy+VGQ7aVIZXg5kqdbm6k/AbTpF+12ey4DgcLBPq5h4OeMg+hj8lE
uxdRnvvp2roiU6R7qAtLUrHi011MbN2GWsijgtW7Jtd8/f3r6DL0Wp2RT2sr
sP838PIE74kJPmFjQoFNVT4qG3EWsyMR6iAOEcTLWDcDr6qPfIe7onv7+xrG
MWP7dLjqqpstW7z55dJucayJSXZa4iNTQVLYx5fwt/Ab851EUIereElAz2rm
h3bs6licFIe9XnH5irxXFw9QWxO3zYaOLL95c0rumu2b+eA0aIGJ/exJ/Gh4
hAGc6zZv7zSfJojBr92tsNmkxx/uZpmIJaqgELPcwQdk+ZEikbuB33Znco7J
M53ujkiUqXmH4TGsK+s8P95IGXHmgOoz80Gg+NrhZMplha6rd9DbUesi9Ult
p72rb+mzux0BO6gh0V3M+xeaOBN701WhzhScqBoMR/rFeQNmxaP2Ld6lSSKJ
jRzDf2Y62lJeYpywvRavmlsFU2262wdWh53uXVKLhT0UJNk1WgtCuWZT4AoW
JJTStWpGaI8QuXpRoZk0BS3GK5dlDv4hnHPzITi8/3WATfVxQTOdv0z1Qcn9
hnM9BmN8gpToYVesq3jHPQPK2ktGcAr7vJdVLdNQ1GH9rzbMGMj2Q0oURDA9
lws/387hgHynsjgWX+QlG5tBri4r1rAX4gPCnKfHV/dYckeXp/+9s8W0tYHs
VGBLtV3g6sYQldChtvDOP8bntcPubQAwMl++s+vMy6oTjcfzaTwPm/USzpd9
JYp2nPh88vPzPx9ynCkQ4bnCfpDNBg4EGhsf1Hm5BYuADfLzboVPWV4Ck+ey
4c1cZ7KhWHQTGRGenTeorgSXOE4d1ts/RPc/Z2b53ZXSH6n1Zs1hVgkIV/4Y
GrmYqijN5ulWzJ+asSAwMFyaffFRxm4vdesrxwiIC5ZM2VFwcG9tXGC3q0z9
zIrcUlq73n5FK1BMfVug6ES7eT8VAmY0CTVWhkU3eRfwDt6FamZLLoCIAPUr
oYHpIH9JAP+sdyCtvhjMM4cf9jABFt0e91B8PJn+lDu82YAaGa8F0He99z/k
nAkM7e4J2Fqffq1M0UyvWxKpe5QQJSthxv8+o0EyEiCAOB8t/O23czDJRxfR
4FSah0/yCVuUyRI5OUSM2ZpMAEY3ytrvqH1W1dgE8Y7a/7+FKGysZm7oXRkn
G9qAz+ZNBpKOIPha7ZMhf4ERMDYFjEcuz9JBQB1fCPRd/A6hurH11p4Ducj9
HY+T3OoFEEyHPvz82Z8iY5LqBt9L+oVfW3ZP8OGcioUmk6GYrVl4BzVEWAP8
en4CkRRKU7p+ZxpGx39ge/68htd9Na9/OzAeYPjoOqB0EZ3jHLtJfyV0uVeR
uDckVIoWSN81O/rcKZGrF0hyw+NyTlEa6O4j8v9bvnezLx4y9RmC+mfvtYp8
GxFsm7q8meIP3ExJdltleaXV2L4cUUFc8btPUln4TojFPTsFhYH1O0M+yelK
LCFjsDfsHmxI4/umqazD99jRDHCMPT6IGgKcw8yjQbgFMvwlENgMw0BunshO
9uU1w34yVJ8RbOUHDsU8HKL1TMNqYrv4qC2H15rPqJ+yRcrTVx4RWSGrC4aC
JY+U0zvEpEsGIbzCWzvxO+8NcBU1+8nfxDFi1iKKEI+my94d8Ctw6lYxIc6t
5BRzeq4AHdBbqYvAnhrGNkTMeWPQvHcJSleUp73Of2BYtszFz/MSb0Wet+HM
hxqkLXHzZFAMv3bFWxzNc5ZI9Z7GjVx/efRkILzqq7McIzK61XkrdcfEwpKF
wFMYj2LMGT3/Fo/JiZB68TjoPNXYomsZGta+yI1kiXRjKFdUmQteBySLlJua
oIpLoAAR7Hyk732rvBQi8ibT6BujZgRgX6l5dFSpcU2vw6k6yOxgLHw/MmeY
o9wPKLt4K7rzJR+/tZ0K5cdNKbfYGQ3Ltme8sRvVmNCpDzn8gDWO/1tV00GL
kTuejxDXU03aBnR1ULbgFKbUHmQwqio430PgGE61vTAxVhgUhDJWwBcR/lIu
YEfbt0lpHE711mOzWGaOndmbgu2nf360Pp5DoVfe2LdH2YfPe0zMM1/Hk3yT
xFFV0q/lU3+CVWFwv3gM1XeqKGG8pgUgdJXaM1noGFf7j2a4sPrts9Jse5ry
6rGny7ik35yvD8iEahvQ8arUs5IWW6hj2UN1jXpjG9yr2DIuOdEapwLc5tB7
XoesSPHILgdAnYmhgOSQbeIWgSipvgSMbq4ojceKuRNliHLVSXLZ5mb+SpNi
fjmhyKF+o+YMdryNy4anItt8nrdRcFvz25TKd5uqrlrjtLcP0shUfdy7qt8o
l5v8MlS7o4CfkK4dFrKmbzxvR9f2pg4gOP5tiNuqCImkj+ytAdvjAWEIhHW9
ANKCaFkLvBXQBGqf0pe2CsEnosfi8gjWfHUzmBjYlAi9U4Dz9ya9CTzxRLDY
vYmy6Z44B7hqj3gJxhGTXprmaeF7xEJrmp59enaNN/1PnSxIIy6e23RG6B9m
Il6LPZRyxJMAGiHMnzBFsxMehnGk3MFM2v+9ESH4h2A/0ruXswlR56Zezb5u
BugPe/hzWIcx3IOdE60xZWEAOY6WrWzn1IZoSjMm2GL0Hk3ecWbS+J01bVHi
lGT8ZK4CsO9I3BBwZhopZ7h4Sz+r/l3bVcmvdkHbs8dRWYrpmEmN7C+Vxf7Z
NcIt2c6XRw+sUFLAPl4QMxMj+FFrIp/MqIlq+Qi0h0hAx1OWKStIjVe1GKFb
07q1kp6TunPJ6yV1jusgM7iwdpRXQnbTucsUBZBl+VgLWQ+MPrG6JnB1b6H6
2mNi6BdHwh7imEJWXXBJ1o6TcnvuVsPupSiFubbe3LM3wWFNwFHP0SNrGy38
nAGb7JIoFtHGfHIcqCIlsBxXHvwzsHjqj+yqWJUYMOEeyCoUFz2uGPMOKVP+
vxpu6eepfi0+ROd5FiuIO9tFiKN5vkL0RmiO3vnnk8jdbvBmmmD/b97+Dnv6
6sdfjVZ+6IexiFTPrdZ9jfQHT3KLb9RjPxS6VVUO3aX/AFEqRJqiXeLjEnr1
UfIQuF+mdBle0LqZEmLNM+16TNDl/efpOaIOkDHnmFfX+/0IqZp9TQ3FSQer
B4RmcmszrV7rvzKT0qEFI8BHS2+HHO0z+29jPp2GjATqB1GhOF+IcHk0jOWT
R3jkv40BAsVRrUYSy/fusHDGhhkG0Fy9MF2jpLSWcoZTDqErBnKuQaDReixO
l2j25e/Ert6K3mg1W2kExKoXk7ryWQDtj7gd04/6UrPTyDKxmYtixAkReG3J
P4llhI8sEijr18uqqX9IQoja099qohYxR4tE1vR+/C1IRvsgTV25+zJVvaat
whtcG0c6xZ7U/Hz6oZTJer6LIAImSOgJWUEWe3BWBZ0ahDZduKg+jHl492Yw
7L6CM2mDeky1HLoQMAyupQbSDuWJ0HNgsB7DG8bI+sHxeGcAZQ2l62FEXY0n
J30Ul60QaQ5NqvQ8N2ON+rX/UdJ4Ryx5tkMqfNjgD9KbE++mgZCWcoFX+eXs
X4a3HCOc0pqUysUQ/WWQ24Qu5nLcfUXdpNsef1dgPG2SezCon7lxf4aMGqXH
p2MHmyBRyaURT4lDgWy2YdmKMLI6BdH9Kf2BiV2rPs83Pk9I0Mii3OL7VEsa
TI1wduxl2M9FtMxBYfmvbIqLO3uc6SVQ+yGVj3YxqAnmOYxm5td7+p/MWBRj
rGyWUncmYYhr+jNSq+tnTSrjy+fMZKssSJxKeqTGqwoW3Lw0f8TnsJL8hSLa
olcEoWfWYatFiH6S3yuTP1q2GZTiVKwe0zIU6ol/pE6U85fx8CsgV7U1TSr6
TtUqbAms2jSai5tQkKAwwUvt7+dFIaX2qS/dp48iG2G3lFgTdcRuNNCz8D1c
6/NTthPp+JkaIQcf/FtdHFLUSJYy1aChpvgEwAFeMMFs+sE/qF9DIUNjl4GC
95RWjWL6evsFldIUlqpwrF+TLtg0Dd1zxpQAIP3TAti662iGzHXCaT9faSSU
aO2uvouaPHTXd6rSh3TjZxurA33InfksMgMaOhY1fga+QOU16U13nKyLTlHP
c0no9s4nXfspX6VPVh5j5daY8LgAS2PfwMncDNZRIm3qJ2rAE4Jq4Hnj9DYV
rfi8WvKc8FT7P2cfR7ioQRgXunL+mth1pqA3TanP6GKbn8JOmGMnOJS7DDYU
tRZQW7v9y99yA/apJw2kkwglZR6o1AfCYILNj+WNprzvT0CuarajZ4/GiFrn
vaO3ZDPeSAIh5vnPvSpoMPih8mSXltVqnS7/cAYSx+umjDsCOddD97uyC/5x
FSPTWmTUb228KJUhFNEekoaPIANx/Ly1s+2TVFH5q9vSt71+0vqDAB3XAVof
S8ZjIT8KMiqyDYSAXMnzNBYucWmXb1wFEVt8x3CYzQzLZAauAKLX7eypsK4C
X6/5FncUZY4hPyCRvTh/+qg8wO971yA2wICyffByEcKIRx+5lqixdYIMZ+5D
x4EcT6L5i4GltGzW+WhvWNZzjKS+5dalYhWhnq1RKdrJwoyo4Kp5ZJHMm0gF
VQNV7dhPN503RJOsNr8MLQkItCNGabkt6w5djgJduBgHeRwtabaz3Ilk2xUz
xFT88a8LCJdn9moF5WZgnSAHqwCggjBC+lzbrDoikCsmFTiPy4+tNzhyG46X
6+OhgwzS8po3DYfd3wML2jaiUjIBfXfWIeRgrTdTkvEXk8RrLdQAV4nufBm6
QNufa5z3DCjxAcohZ2TDV/+3f6VgjexWzhm7GLeD9cspO5q3g8Jue0IN0dpk
KL7mSqDsUzvNlTnKLYcjgSdOO77F0DE/2Gx5xsHlAi2jO7UgCCBiU5IBtA6J
YAyzk8IW9e1xotxPSH2LqSHpzsgFgGk0sMkw1FUQY6fSD0+AZnAE7rRrc2bh
sZjj4Gh6ZpCEaHD8lWgKS6JqDrKR3iE9ou1EXgfl2Q1VQsRfbaAVBU4k/hc+
QRPdx5PqbVmyRuZSwszhmLrWPgI8+YIIKrZqO7iKIjZJ5iCmu+565dlfa4Nc
eQOyU3EtTgTzNzJEte8Lslhcj17ji7/GEKDPT1fqJWyzYNM+wWIadMp/qIjV
gcjTRxa34a5HmA7FsFQeLf0i4KaZcZUodKyOCZTqXZ+7QzfRhPK8JdOSYSNE
YEOH04Sh7O1tcQri3JPTTcvA1Za8bTTSR4ScfeZy4TyJucWEI7XH3rt7Ff0S
GYffZaDkviB6xw9UDW8vvPKgJavJJ4q8dJDHplBZzacbtgA255tZL8Smeyyr
q0G3fr9C+4YvElrTV41edFv4Hg2dDm7hssVJIfmDBuE4F7Cvqne6oLv244Nh
CUXnijz11hdY/z623wqdHMHi4Wx7r47i8pypC78v/H9NsnTeA+DMFkSl/DQ/
sYXYDRKMKnsRLLr98xo0bmvww7SCf7muZeV/62t0l69oeQ1tDwnrtTDsOMvC
U2SIdGD+zMqR/2+8bGANfx8pvhqYtaigL/cipPFpBfO60eLedJaroEF7uu/B
dobjEqtehkymS723d+Wstt3lqhHnt8zJRdrbsDG74C2ToRkjGuKc2T/L9cEB
M5LpDky6hne+Oa8wFWI+HtG4BpfA9A3MYdU60SLfCriKRcF+E00aXj6RTERT
Qw9vK2vXgZuJTWIda77Owvrs7uqUnFcgIrpfpSoJxfFVKQh9hf3p/kTdvg+W
yXLcrYpO/jSqUbZe1G3oqZWX7Lmb2i0IVu98+D1GWhDCeSCk1BfMxFrLUBsS
FKrZr4eVFXK7Gg4m94ODNTexUJr0Sil4AYMUVM0sUSOEKsRK2bt/4ecLgCTz
tYHzIrPJuu7vkSPJqCyOzS/YeE3+m39WZx8JlAO3jpaL1AStmHXfkCfYwM4R
msbTWMu+WOkEJMYnQtlYO2eoY79lQETGxGAdW/Evutvs4fPkBWTt9dR+UDf7
oNyo/sIZdnDst52Q7rvQ7gpJvpbo/ndJOnB/1AG3vnH2q9Au9HKhXAaYs2PA
KH7cjN+F/j+YcdRytNhyOaWSsNksL1ZFWRYDDYM7F/RvoCn0EdEEl5YdGpdq
TYxg++tKPqKvodb+FkfPc47OGa0Em3ta8noSSEMsj9WcD85kzJQI23pobiuN
jVwTP2urYrufXClys4JzBj+ncCRPeMIYTF7eMz7FG07ApFmLSOsGijq1hxwI
iwgcx6yYmIevN2eNlGxTFuwoD7ONDAQ9/s9O7q7qdPnek8coCQezgmuJM1eK
li+kYXpt20OHvmAqgZBWcEbAp4HqIYk0ksjPzt/+flmUdXKw3U+ljhxfV/SZ
veCSJ9PbM8vI8BLNeoOX4W8ypV68L/OsHVbdT//k0qy3/S8AEABrHIQSJ5Zh
HcmTmkcXSQN1nV9gZONtIg0EibSAHa2L3t5sOQi21faUp1E0iRk3P/6pzWBq
AYdMd4BxO8QXIGyko85yhTXhc8WwGqpNoz/dD2w7ysnb4fJmMl1F+RvxUXPD
hf1lgMr6QOhJloYnZIQB/z0ALnc9FOvlacGXk5eahoIkhSp4A2vI29vBb63X
aLJbmNGJIfOCYtpKIDlf0Bptlb4PFecQweFAo23pzxq0gucaJQs3lcXfWzC7
7SB0zPKUoQ1lsut0oycNqXauGzrdfWKDC3QOOWJvaYHdAMeBAuCb8UZNPNJq
4piwFVmfuRMc0Ni/jb90hlDJKu1STrqBdpcmFqICJtTL1dTGT/SKX5fWQJyU
2y9CNXZt8vasgIB1d4MzMHbJvf5/PQshtdkEwCdL1k8JoLjtHDph2w2klUXq
bOJDydFX5VXCfOvAQiFjtZvXbrnR8iKslOC9BQjC9CUiNnFl5MVAvGdqLJ98
I3QN6MYagQ1wFNETHxeMgYAKqoRy5zvK6cbcxJHEkj0LTQtAY/1fOBw14M3d
FRS3INPRkXJ/UBs11d/PMZQzztJ6wXnDCZqYNFI1AQw7abdmBAJCx1V+uOpl
+vIR8JrydRoB1t/wEom8dTDLG0QjSDr2KWZ2sILhvGLF9Jb6IH+ciynt65BB
N1ROfexgoKNavlO1UUwU8tKq2uvUC2MJc+vZ6jeIWDU9evzjyM2sCMmcXjAK
BejRDGN5aiChKc/Z21GXw+//sqZAU0FYgDy9J3l5le4SwR3A54Wv3c6wIhNW
8VXMchDAVso59QYOXdms+AGop0m5+dF6qkdF0n5Lr55Q5aCkFqYdGqUpM2Pb
4YbfBVpmBU+FSZkEibSv2hSLWHtgeMt4Gmpet5v/d66FxrLPcDFrJc7qxATZ
UGHYg4DQqITEB+tO6za1zTL1Cq9eY6ufyclAccUcRxgjHGnnqPYTI2nfJexB
h+n9XmpVLtLgHncgDJUSNvtXlu8dhnvXVa7wYOseCkhA77fhGgzFueK3BrRC
QQPo2GXKVfy0I+jLSZIBCWs7shSnVoqk3vGJXMK90IfDX9c92Zc1uFWnkZCH
cp3oqzChIUNU2LTCQfs+HYTp4SEleajOLC4T05IH2t22duatp61JJzJidH7G
Lyaw6uy0/BDWsMBytTFI98bm+DsWDhue6KblmgIfrP22cS2jUfI6OqmUW+hj
XctKq+KL0ny+7xMed6U3YxZd2A9mqZK8xcA8m9FLVMsP0CfQpB/0pyAtiR10
nZ0mYNto0Tvl4ZmVilyhjtEpkw1w3B2nw130cbKvi63tI9Za2sn9pUn+nOTB
6041SNs26RyUu36bvGP7qCJmZXnBNKjfyLDgh14L325i6Yu2VteU6aC+wCoI
L0Qqbun8Jt/BidzHeG1yn2GoTueVXFLDNqEVA0mOILt/gxrQQ2fpa8i1IyRb
Mht/sa5SWr83kpWQoaFCvKGPPVDBvv+oKKfvurWVuKVAKSjgH8WQf/kJU4jn
qxzuckSNnv9vyDxRW9LtdFXzRuXCZLeIv8dNg4hBStO+eromNKlFuhyimmDD
8aW99k/BidaIFDvP/yqLXcSS+2yv1L2Q1tYkrRDCgCjuBebSzFSW4V0dZl+0
JWJ9qL1pUcEmkE2HWgOCPHeLSTzkyWtuujYTXqXB+KHQDseqG4cNV9eTfHCN
DuaiqLO6lCeubhchD9OeY6c3qe+WftTszlHtvhAxG9Aj5S6QVkqfC+acF8Tp
7Q3ioprjfBBYbYN5dAo09ty/ZuqvxlF+cTAKriWz5YxgWrM3y8I9N/WaCg1v
pGRwdqQTdTEwdPesNd0/jvwPFIHlm3DAbUiSzgmr6hAKfw77Wc9fU4Wpumbp
gEC7dK1f2p24PNPOYVtAeOdKeFjh3lxjXNkdRyUAsRpYeBi5lytaX4i2c+bR
Ltutt+Rxw+Zv2InDhwVmWWzXuKQ+/0wVsXIZpQ8AhREUwQkWoD0kvML33KWh
9/YUEceTrSRqQynlFTueYFNYtyTDyjPcNvfa2HqibxKH5VkSrEi3D5ZWdGmK
P6SfzMx9AZkTyMSUMa0CVOK6TbMyv+V0/hpTu1iXqjXkEMTscIU6EJXg8Scu
h9K6OU9S7jdQKMPvcrqst+09cSTDkw45fI8gkt/COZTkIRYQZdGwMmEHbwHh
SV9uy/tHHTttOLdOwFuU8v7QWPja/CffudpvTf1yw4Tw/7M3ah6UeFXUHiL9
my85nRV2UgmyM+0ks1/jboND84rfuirfzJHEWkzxb6s05xjM8mEjtgex54yR
UZEzglRWbLhcKmbmuGM2IZOgVdAK3iInt8SZAQTBDay1zkY+o51a2LgRtaun
KpLbjXYOEF1tlAeBUFq6wBLn1RJXjGTkOfNpGvVh8bdR5zK0W1haK9TJ3Kck
JxfSsPURtYfs0quCtX1s0M/MyDEka86DoaPOyw3nvHIOJjMbDSyAFOlSd2Ym
m95jiAk9YyCBzffjCZsBkDk53u7ZxaNeasXzrpxaBpixvMFzz9ysbnmegHx0
lWofjmbXBsW9xzS70yG/7bfQIKbxKEtzEfLOmWanOixNA9Auvh0KjTMzMLq6
ozA+zT00WrCveEd5kEZE9YJgfvxU+kVnHaMn8lS0f4mwdMmjd0wpen7nLXXG
W670GaKbY5g74G69Ri/8u8okVx9198JPX/xI3cmYZvXJXgDZeGpzTCvD5ZaT
YIOQOxBWdXBNMOjc9UYgOBAIoIseIHViS1eHd+SDC8VbTAmHprkxaQF1g0Xg
n6opkIldOYWtL2+gRDTZgGyrq1Bz36eJbZWDpxGW+8hDy+RTYiM/8PoDR5Mj
2rPj3T5At2f6lLu8ReedUp8R2jwuypxbh8CQ7ZBBuiajSqYTK9ZF3RSHMN9r
0wVxCPpfc6jHqxgwp5w7v4RRZP9buCBqjDRkMwYi9iKiLsTt8cHtLLEslzKc
6qmD3HyV+TmNC3uVaLrfvzolGMManDdLMYr6gWhq+ll11PjiKYg8JOnyUhOP
8DatP5fmYTjkcXTGKv68HZHAcepE2Mazj1E+0RZMqRAHsO4bh06UyT358FVG
bvQgkJYkeppwO1MseFO1v1TokTfuTkxJzd58bInXZD0gKJT+aK9jZxUTSf4a
LseUP7FmPMNL6nUl/TI10V0RTJ6whHGUGoSZOBcmlHUE2KzkHH5Q1Vz5M1PP
FFnbOJMwiSZPkizMR29YPsRnEFX5Kbf/jcR8M1mDL3Ls6ZqlOwlWkfngEAt7
9LncBSIT0+UJTsjrdYc830qTBKv/rfvEUctgIk2AkJ+I2c8Ib5nnzoLZ7q/S
uHmDRZTUd/4pEIEswYmEX476RwYbuAMhB65YWd4RKoX0vYS1JQmxGc0XyI0y
Vf5CPfQH8iytgs9uwgaW9bOOD/dItkgG4qf22bcYm6JNZQiLrQsqFTbXea9Z
EMYBr+KDFb3ooT6CN5xsxEW8rYnTxHeynYZp3CuAG87ObbksdgFixopMReJJ
h0JdxYhvfjvTmfQtOHKWxxEB2y3tHEXufcXSmNEvBsriTHLE24DrSAXjpL64
Fnea/c5GNZxDT/kB+FnOuOy0gAJTwNLXDBUdxHWuWB9jqAWdMfjZ/HwZWpGI
2NN6tuN7HOZD1VlekWYbvGJzcW1+xhtGKPprpYtwhEucr0I42i5RnHY2vAcm
h1/U3xmwJ2Sfc3dIs6zFA26kvuSb3ygRbaA7seiomqjoxIYUDFo0m5mowMIO
dikmVIE+aB9t2EQdOvHsuuOTCacrEDgXBgrvaneC1aIevKwTAJKwH/BBayA3
WbpcQIp3jEGk3TqJGzz6m2ITOKxGRbm40qv50SWDCPVXL8C2s4qJWJWv6uQC
HP6RyodELNKVEMzccJxLEr6lZIoT2wsTMSlPseGoD+xqUAGZIdeBTFq5Vude
8ag9Lr/hupMeBTZXszRGKBIhsVa9TaSNkrgMFxVxKUVgucZNzsfPUkMtuM1V
6icN3svfyW3sgWOitZbabRAGUm0f4aF+1EYRd15nW26M5iAL+xLtHsKv84sg
kC35sDC6uFsi/s8vu4s+b/SczeWjzSLoYnZlafAe96dj7mQKEemZfkG8BSaY
2w3EPassjiEWOXL7TM+KyluhRzbZdmavlBbWYbXjmbPCBD8Ikzg/PV20Mm+e
rOJJbHEtBeK2Z/Zxiopp8kRNeVynIb0Qa6oLIR63v2vZWh52JfzBigcNW1IH
hvVEU3S9eL9JLW0knIDChgW1VCZCJ5FBvao8Bw++TAxlU3fYeWyuw3ciPHO7
/EVGDEur4LCQkJMGJeOeTLdeGjTRxr5zi05yUaGGksDcq22wfLDXlwWE/loT
6lj8BYhVVotS0DsgnwEVwFz5gCDqL5xZnHM37Wpv6bTs4pEIrVkeloBgmSQM
vQkGb/cJ8Fwt8yjWaXhvy1vOLF37Ayx+aC6Yds+YDrl5xlTAMWQ2Ym0O+rNT
jr+3vRDyFJYY4lDenBur6K958GSG2ZFbi74d+uHQL4JsT3xWyj8ecb5ZFEVC
yMNzJVQJZspkHELu9UyLRiiczW6TI9GWtr30q73I38Ap/Fx96JERMomsYrxW
d4r4ujWpIumU51JtAAoFgYPTH3p34O2sqt0OCNR/Z6q9O6vTA/PRjzT+KdkO
wUuunI4MrUR8RUkzKo1aXAVoolMYm6bQQ9DkdXoQBHZEPS63zXK0blQRXIOx
53hUmK1ft7+nw/ur72Gf5ni7qh/Vrvbwv1AjeLJxMiNOGaOuxj5l/R/Qwzz2
Pd/oNWXO+u6eEBeNm++HxStpVUZZ424/5/smU16FZxdPCRGjMBImyRpy1oHg
Oi1U+plTvoZAnTaCUbNkfU/2L0CM4eXR8jconxf8/TrpIWKylRWt6uK5QQcx
fhDyTYnvTPyN+Ut9ze1WkMvsJaBFOfJ8x2GdTaHp5Q4frxap7Daf440+p8uo
CWlYtALuK1Qf7TEqLe8C52Dme7dCDQMhVOSKZzRoGHzi6/d0+Jt8g/7rCgd8
DP9sywmb6AMoVTV2kVpXyHVMsa8npzsbTZh5htFChWa5OAcSUeHizIT42N4D
dl/StvevL6+2YdysC0qp7J+vC486NafLyfw6gg4SecC+bT3BDPHabiS2krJs
YjBes72EuhjBfgEVL6p8Z8obIHOHeFKzRYKO0hey7zv7Jz78+JfGJ+YV3YMP
gfslGrebRm96EO94b0BZ27b1mFk+UsapsPiP1DqfWJazTSEBXG0v+F3/DcZq
d88jqDqM1ZtHPgfpe7TTjVCmG7fBxTp2eki6kdHsBp0Ww6mqSwT75np5mPbZ
sJHBtauxdPpnZL51gGsnKlxefXKFLR78FmzXRchN/UvrflUR4aJefAznYaM0
mQP7qnZRruNfmeiGYyBP711EBd/WQ5Yz8MA1elNiEEMbczySviNsbNCV1FgC
8K5dY+GFov14yBiNwcQMS72l84PuTr0Is9WZ7ZYCRs5HvkNoIOfJyksV8Q0W
ft4Aexy1jLTdz8m0EgC2oHakWlW83VukN8iYx7vvt4uOoeas/CqTQDXZ3sBQ
F2dgXrf37ewLGjhT2GosJU5vYiXpHlok8ZBrEWav34+tIlDahZVYGR3dTmFA
J1r9Z9aHYPIDpbej7iGvfGAOOViJoJ4dlIP9ybstcslpQAa20hhVy0fiJFEO
jFjLGCjoViZqgYWZrysY4Z3yursKOPvl0DatLF3vRoNylOg31AidMGahsw0Q
npkYBwdgM86iBqp2/u7lGHa5AHe+a4AbiFPXzrte8+2tYm8vBSh1G4Qv4YTR
1AI0wXcyKV1gP3QSPLXZkjvprjvsHGW+SQsUE+hgMC6SqjIpmI7qtDVEfQyI
vZ9e9mYKdkqP8VwcPPpVEWH7mk1Dma0uCWpK7xHc0pFx97WpEVlRJQZZ5N3I
IZzTXjcDx6kF4kUMWt0w32mv7pnWSfyePrrOktG95I7L1q42ZgyPaEMBNr07
xaW2oZoDS7TLD2/+ba/iQ//nBps3sw9Y+npTiexMV6XCF3Na8/huceKaJ7r5
5fcFSXMvSZq0jvxfrBKDnXCEUFCmZ8TMC5LFyJJg2SQ0uTdsQhUYaPTgWQYF
f9tHHhscVl8JohCeJcEvzj4Z9a5x1Fl7Bjc4mBI3ITN0VycroNphXdj5ZKWD
vnrFHp8fslLj1By5Z/r1WAUGvFUKq2Q/mLyvyJohR15q6J8uRe7ilxPWY55W
ogyUiRQJe0UY7LTgF8LZOLfe7Nzii3sl2C1eLzEFbGi5ehAD2yP6ZkJJdrjY
6AmaAKXJjaLi3IkuiUhw7U+egibXS1WXKPxwRqBW+wXltqDohfyJaS0tF/b8
PKEMf416zG0pTgBRVrC4ik41JaYhN38WbgRZ2rnLMnTxQ8Q/80EK5+zXecmo
OzOwx4uNiBYxvVo4bnXb0edOhhbZEIJE7Cr3BjxpAQ48MrQhgRZz8NjXUKFC
VE+/Bf/XAe6fbrcYHAc+y7qpiIqo0jpXTPJJI3NNdZzKMZYNrV+mMgWixh7t
UtdhAvRbl/kXI+1jC5K/Tk/Fx3qk8A+x9+ZG0Jvge2UdYBJqTyLZbEMcxVEu
3RzycFJoMdWw2/LQ1vqDfFpmaxeN+gOJGUm/qxWfa3pTEdF7W/oOQobFeWNC
nlQwHHrtZ6H6VLZ56ahjBXPWTV4Vz9CLuxLRtxK+cdoEupxZoYaXs28deNQq
gr00oi9VuIKhaVPiAjQFv2wjnelRB4HvojTTRLbmMARne7klBHf0+pKi6rZO
ugjOI/6/616ApZ8EBD+N5lpNHbi3gEA07i8kvSKFN0NrVS3cedP+z2qIQ8xL
jbhfXIUgqtsv1vi6JkBkPwNCv9/rzAGGxqm6Lo/LBWrkeAUT0r7JoGJ3VUm2
IZP7XH5pWtKFB37kE//aPz6YsCMjNHN49PUrryoXVDR8BLH+p0P5CuMpTvnd
XpXAK//u6DxKQxR8oknMXu1YTpxKJv1ny85vAWWMKtrAy2l1IueKXLFHzP/D
h9800th+WsuSNxNBGzRPRVfieCVeXAgEY8+VUsEFwXAwSDXF8r4V9gPNGmgv
1CVG6GVEDtDGdfsFEkU8gLBfA0HFcPlnfy2eErDC5J0Fl0NOXkiEA4k4TQkD
Nf7glf4+GsyiAq8OOBXG3u8JjmrtoneRnXYX4R1MHa7v2sJxnQhP9jhswMVB
/nsSfsi+vIv42wZFyOPjLh+dxWJNTRdsGA+Icvnh3cJSyF3kfR42aUqaymZ1
jdxGymnPOBEM+XSUeiLg0gOL7luz83IsKehQYz73Zf8BvJbPL8hIc8DtqY7B
AVjEg40DdUDBJqD3u6/PlOK6SKaRIZL0hEg1Y+XoeyIH/D46xkHY5d8dIs44
RuxnXbR8SqxqKYiBU46jNqDStrFPupFA4W6L0EhgHCFQFNyWFvBQcr9AJ1ec
6Yb9IrRil/mnUvDvX42nbFbP78ZaCrGQ7v4sxR6SS6prMRA5FEo6ofmt1fHm
O4fbJbHGR3Bm8jGVaSoNWNPfGpyAaQGrhqHTyBSsA3BMFPu7CvEBYcavy0TV
y/JBuOUwvizCb8LvsHXptYCjytdwH+zU3ilZGzQGMTgTRskxifWnmtyGsmHv
yKE+1056P6d1gK3C9tacr/uh87KatQaf7ICjnb4zf5JF7z7xpMcV8YgpicEV
9QEOXjF4l/tSh2w16+KuyN4R3apLMZIvY0EI42fd5kaBAqfrmyO2G+X5nPVP
xaQe5JTXvPxByLx3tdJr/TlG0hPN7DpURJ/UHHMWb0wc1HpiyEOXLsc1Vlfd
RVsHa33gh9ZwJZXBujG2YbKpRI3QMGW3QVLcvknV2kNB58+osHPDUV8dcn3/
hAj4FkNdFd2V3/+xaghW2NVajnq3fYeUj2pqQCAzSD/Sn/MfJ7qPJ8SDzLtL
WD8DyhGbm2orY4EnkDnLePOCAKpzA9EYxFWWycDZ2kYRfQMRhDKDYi0vKcol
RhOBCkBr29OJgtzMIp6jXLnhspq2X2zuAdUbT1gwsBgaZMyMkWb1K1Vjd6qb
y1SlVGh2lPj8W8Xo9uTsHRnwGBmz2JhIe1L96TWPlz/4IgCyDQx58UUUl9gN
TSitT9YFxcmPGTTFIVG+yYJ0ivQ1jay+YVHmdw0yYluEzIhm96kaPRaV+Jyg
+6lBM/JKFu7moRjboppFLg+mqThWeQd6lDQhAX/BhGz7giUZCR61d9xqs/pV
Dt4lQlc9YM1SaDVxEMcemyImXST/SdQMCGnwNGuwtm855cJSJZ2h1/WZTlGM
o1j+OWUS3hZG3fTqAxoScUU37RYrd6GS4UN69vv4lUCrwzezJfxXOwQ3UK0k
krYdomNu2XOqGnsKzXeFeD0WHUVDAzDSDGtxMk6oQYFrU7RUEgQDyMz6+qp1
G7lNvAMGLMaMeg7lRkpl5t6zcWue0qotDGs2wxBOICfYTP2YO8rySTkAPom0
Jjhjh4VQZLXeFYsIsuDN0pCWG3aehtG/sWLqGseStkCbl2eWBgZj5qayCe8v
mkx5lLpSwcdT2Xaou98mIap7p+kL8i+qP6znF828C0WuGxCZNWxT09SZSnoP
wq55ticEq7ej/pzj75K79hIowoYJRuMaymXDSq+JjXds4cKpCGSW7ErOggjk
57Ld/YGoKbYYX99x46N1gTf3ODqljHobwmQybyATUaedGLrFKtrYZzElEWZ+
Y8JaykhI2ZzvckG4bHJQtjd8DITZG9AKnVR68kvEmYlsXsBrhxwJzJpjg4f0
quBap5loDzW5Vvn17RSrJCTGsAfIU3wzR0gNo9gHp/fJE92paNULysU5Cm/5
s8iuQCWTPYQ/d8BmoqDnQ+nd09ThVpqYuouQPYPZndjS6PUEEro/zNAd3SH8
47l+RRg2esFTxVOg+ZGMKysab3O7jZBqgrJyk7nRJcqQWz6CKntORHFJTZTO
9GRNrz3HV2GGqyKDKTalshdouxn5ePJDZeYN6Rm+RwDYMKg97xhKGvDCFiUK
oDm04fx9mb2u5u5Y/m/Kq9fJe5UHwPofKXQ1HA6+fmVOrong9RQlpabcMNJQ
Fx26ferNfKD+URDUJeZePBHzQIEqyz7Sbdl/qEgi605Z5mOiqiP0IGtrPWW8
D+ZmVgWq/WXhJ761Lj0rW+iBlef338Etwweg/arOrgoNBNdiQBzy0tvMhw4V
BEUZ8d3nEI5K+e0rpYAL5moGq3591P47otwwXT5JXUDAYwH+0TGbZ1w3Grrk
v9zkE0UyO83lkDKspnFsat1LaaWY10F4y3EqzKD51Vp1GhMBVw31E73jSrWO
zEBsa4F85Jf5ZlXd4QpGNSST9blGFnlMFWnN7AexuatT90BR+3+CU8qNl7Vb
ePk51oQxLTKo24Gg/v1jGMPjVVslQzMmQyC5vMXSN2Sf/kE3S0pICp+ow9Ra
M4AKbel+wyeYzBeE/vPjngt3CcqoApBVilFIfU9jI7aJLVOct5Mfd8xEo0PH
12OWQk7r+lt+SiQQPmefKUslCieo/zJxc1vyA1xYFR3T+4B62jYxaeketwnB
RqS1/DcLPJ7JhKi3DxhgKauGkS9BrgiuBvJvRtxmNt/DS6pshs3NgQq1qewK
a6jc+ZTVJ57EWPfVYFE4DCi7i5Eb3ORZrgE4xkqOpJU9Jtvf+WyV7vMGSn+K
jodaruNhZ+77QPIVE7o2aldBeYn6yjKsVHfOPwvUe3Ws0YB/taC7+RRQ0IGI
LWzKPGL9LFZSVcio4TWqg3QoAonxaCyn3zT92UICd07Ny8I/ipxNuwM2b2oL
j4lsvJBgp/fPEq918r3Ff1VnirijKGnWeXXW6/z7qdER6xA2w6etqmSaHNgr
k/1jz+8S7KFtae20xMdQFb8crLq7A0WzOi0fkiRRpwt3OfZxV6BSdC6kMvL8
lZOVqpdo1b62ujlFuVqAMk8RtLHRuO9PEtaIb5+26iIFOGvE5HTFH0ZIPQaQ
CNgJxnOdfORLsvNHu7xnClxKOySRvhsxxmdz0PXQC3GjyyyP2xHmACF2PbET
Voz4B/dl1Ea1zcxLM8qMG6QrDHYrkgPvG1fp8g47oEkub3EWsmLGBYxOyGrM
eJ6h6lg9kdbRh881BItPXSjMQ/NxcN3Su2Cu/ahAwbCKjptJWivYQpdJEzmn
l2tKC9i2ARfABd7OFe3W9JkGg1DxJ4JT97bPEPXFG3QKyh/c10bYHz8+cH6S
ye4Np73dFdVuOohmfWxHwILkExPPZtWbb/q0Y4J0m5LcAi9RQm8q90YBFQR1
QwI1XdsPjKK94gfC63sHPBeU4wWPfBw0nwk2UsrU6bwSqpZEZYUvxm4ysaWe
qXuXNN8PH053hn2gwfNbX+5NsrmyadonQ9cnTT/RoJBekN5rVOZNzznS4O+A
69xx/kW7iiITV55nI9unHKl+LHFshuRS4/Ud/nUwEy5HkMIa9zO9/BRPUR4q
lthrGQama58S3pCjp8jnu0dlMBN8IPZWHp5JbXDhWuFfeablTScY0atun8Eb
UrMJylb9IdDQejaqUc6G5oLKRs6taUPQX1l2Feh3hCrbfKUPtE5KifX3yEDw
OS58IwG6a8tXQaQuTwNgh/IvZEIPos5QPR8eVfVTJ0wHFf9CQqvUa8r5lwJD
LZz6wjNfCAh2lQo5bgWAwRf+6rbmLIablnTGN9MJGTvT7mk7sJvvRguJ7okQ
jMyFOqjYDWoKoi7d15Qbn+WFke9FrZILZ2sXY+6XB7IJCJK2IEahFfNddZcY
EhwriYmTQS+xVbIsvkfUQHmwodefCPwr/FeqzkRaNpeyhztiR36JTeuXtZch
gv8Qk7WLJWWpj9pHtQFBs2fVg2rkNBs8CGotP4vYFLH4C4lLy6lRaiEckDu6
QZ8w+MXDNKpb3ujf9zraZCK1BYJlIWShSC/13Yfx5ORW5j2PHud9O4VHWzOW
i7O4/BuEremiBlLHxeUhHPBUA8AtdzCiJq46711eTgFzrlX1GqwLpXV8d7AI
kgaxiwmltlGHdhs4F9yTAWsZXrhzZTf4SDdd2DL92hFXWuQAnT+y17HRnnVI
Lwk36d0yJLe8MlK0fve1/puA8BggKk/zrA7fD4CppWBH0utEA9/26g5FnfaK
6lFMSMj3ePBC7eEdhpkrPp7cArWzw5Q1M11mxbg2NVIOV70gFgQxvkJ6tqBq
xViwqp+M4JNel2xQapg/MPGK9tod4Xym9+is/4fy4frOw7kYG/LixnlSmQeU
tOHsdhP0kaVZBArqfHrVwCAQ888OiUF1s+IUEJ+x0+c+zo9O0MCdL+jBNLEH
jRsw9ViSy7R6NAdP2LeWRCu3l6s6rdhmZN8FqCOWm796gBkxOwbY2+VQb4wB
Nyp3x3kfBSe+7r7etwPoVwNa9LH6EyoS/38NKMSLaM7AaYkQQpQ0pikYeK/A
fUrg4/gY2h9k/9T+TTOO86xopWcu915v9Er4C0QcTqQqPdowIk5bB9WvmtW6
/IQXqkx4V7iHJFUxA0lho56Vv3ikYZB2gkJxrXzz4rcd7yPQCvQuLS3AeEH5
WZ0ZuAiYSdkquR4Xb58NvmDKnFB/oleYQWIXFCzsIHlDrZsnHtQEDx9zQ7Zk
0vVZaUp93uII+N2s9yHRSh2RJqK8H2bD+X9g8Ek7zpNxLcCBi/H2GfvP/NY9
yzuPWv9GHtFGe3YT/FLXpEEPYWZvwSYX3IkgGaD1foCkv7lxXUPJVwJd5UBX
S7a5Q90w3jXM0gDt2cAsIOTKkrMlz5c6wJQZsyK7ccj10FKhYYHyTlT83Kel
t7wqd5tb8JXKjGwqQAMne/Hq5ZTJIDoX+ebTX+3qA2+9hYuhpDfAWtQ6uswh
jkIC9aFVwZf9hqK3SxPUrubR2sk2CkVZjx6gnABcNyCAU2cAxUF7s0mS0Z9J
cAv9nPICG5pY10W0z4vgcHhY4pBcYB7rTnVoOfSFY1aC8z3I/q4DQOafHrHu
L98mrIARgIVpkgY5ZApGYw0xnJ7EuvKxwMoH76N/W5NlUC6mzwT9+hTJLWeR
JG8cGstpLwSTH2DLecyO4ZYzUVNTb7NX47tmHM4PC3jhsppgVObJFFgop18I
kSGKyFGMUUQX10YWLGWmvfSawLf/twVBg1jGVVJ4qa8PDz0w0j1LX5GD6Qpp
rtguEMFZNY8833X4ivObZ5+7EoqyAmoO4seLDRRGUuiM4V8yBX+x/0Ed/HPe
2o7Tg+cSmSgh2S+QrXQ2bBk1LVUo0hGUOBZHpqXCVPy61l6ZIqMrdTWhPL40
dMC9jXYYcNCkFVOHVCkxkLAlCo3ZpbJMn87HF5FrPxGDnFRgp3dJBsn3zeA4
Psurkz/hcj6DTeSpQBgMugnjJI3Z5Z9frZIgvBBAZCF9NICXbrssSN9IGwHQ
BnphS8BRVDaqDwx/xPWH7s3KKI/pPnln+iCrD7F2uKK9WPZ8qJiB0Amlf5rK
hxwrCJIpk4691dHrx5IqImCiBVuRO1+40U1yAO4SA80fZzhBZK5GBrvmeolW
G8tQ0wS8AXZqZauIHqbYwpzDdxniqfyLlCOny/Qx7pDJ+Uf/MNPvSeD76TkG
ZhPMiIIivBKu8CfUuJ2kYWINAlcdeU6wJyLutNTLNwqXcSItujcTZoj0+JaD
qL3ZgOsHpggF3DbWmHPa4N2g+u1By5fb4Ip/jvSKRBQynnWxR/RNQPr9wN/u
qzzLCNPZfsyOGqF/9SbuTdOtZFVgujCd0pPll9nO4jrhE857wsEgJ2SLfEEU
zqXFknH7edv5frTw6ui2MlaqvtmJoxbIlvvxsYO+TwTMOhqrYo2IdcetZ9pN
e4EBdPJ1Hc1WW0sbb8nwr3nhtNspADfafwdslax8L4Jg4NTiGelciu1wJcag
Qqq8Vm4r+jO/EzesHqxt4D1jYG+puaXgrgdzUhCxtbpUN/RyEr9G6RMqHd76
WVqhhyP9ZmwgrXO2CSBsh7D4vBM+ovEycnA+VNNKv0TTGQLB0VRYctyCnIBM
7wUOl/99yu+0oxSERsAhJQypGF2T7BZfxtjneNoBNsxtDOte/rnc7lrEFLh4
hCNXlHTtjRBo6NnxJoRZMFTy/0CMvhtJTFqaBARQ4ZqqUdbwmtnP/ZaC88pk
WRLwkweUiw27oE6i55Cm4mSWWQ5x+Jh1f3TRqWEyNnqpIAPmisk1+3JtbU0l
ZuZEvx22TDV+UGvBkDUNUZqX3CzgSRGUCFhnSDBdmkYSINR2zCe+m/ulNNQr
FtAqfZN636QRrkcAFpvj+5kN5+tEyFwEuhFgxIYUiBhXOLAKtURgBmCtifuh
XRmlvofyNwzxlOJFEl3IOc+8YyMN/Pnd3bIHfaf1fSdJFeoPri6rsYB/BA9b
6AZAQi9bB+jV0TpQTaqkAOxBfd6AbfKTs6lPzFuhFaThRDPq2H5XfDVYuvHD
bvFdtZZx6FYsjjxFRlwH7Q3h3GjZLRt8cVsQ4njY6kLzlO1GKI3Ga8Z3deRh
kw6pQWPVY0QdRzUQSwWgosy48thZmmsKncGjSgsOIUk5Lt8aHIr7O81p95HU
V6pu63Gittxqg9uVkKJhl1TK/ZNlZYgZfDfOtQdWTlCq29Vge86CJA2Alkic
FHNs+eXQva+Rnuxe7uH3l0rWPcRJfU8JEVbyxfpdFYZOnLG/jUvlQV1J2Ki3
HGeQkjIfEKGBCHxS9zakHRBxdXyOz/HqjyEYFPSuqnH34j8z/NM2YaErrkUg
fxGzBoRiK/pvRiz8pn8GN+oatClUvuOL2aDbBI1XHe/OJ1kRBv7zx9pMAAxw
ef/kuZZzjPPgPn1athsjjE8QSa+ecgKj9ejh5GP3b+ToIWF/vqoEeFrwmIo3
KG/tuOUzZkX93Fu9UqpmpNxfFHbXQYsjPntcfNvA0EcbLmW3Lt9fN1qhB9EY
wbWueiboFhwDsrxUNJyLIPKpkhude6w/p3rq85Og7WW468QKfvEFCX2AVsQb
T6Nbs6p0NsEz+Hhqxq+kcC4r1RwC0HeCRLtmMExxUIpurVaBzEalzxpJRr/3
FwN8xbisMIiNv93517QX9AixUu9VOqq4zfSnSCYRWhfMP9S4mpt1sth3fS03
jW881qHktroB5mxeznQzJ4/TsCAaQJM2C+4/EI2jQCJyvPWB6tDURpB/M/dX
se9ms41S560QDBkvFmiimQVovhUPMANqPjWkWz1t09y9Cysh3LNcdN2TKkST
bl88AJtDKahn8xfw+lbJVqedZhjgO364CXoz4PWMTRFTjbT9CBoeksDBatJT
wSfqWqY2yxZxK1dj6qIPGZ+S/soNSPuYT8KUnoN9AzGQQzWjaIhfCjRkZmPI
npgIhehkdvNCOnmD8nHVbfewdWSVV34W0queP8uKto5UVoeoRznSLbSa3oW3
KI5viJlICZp4nM75d0Ry/yHjT/WAUqxQjg8FHGEpav3pWlPGGEyLABqQuWEt
1NgilpHdCIwZaQt8udz6vtHuRnib7ut9NN2XVbV72JxDJj299exqH2aavMR6
Vn/Bz46Sn7c5Y2zcl6zZEXU5dMyCfHmCbbG6DQmz/1vu3qSmNmVegE/aSIpI
eBuMW22Lj38gJfFER8zylP6fhOqkgYqUrO+Ey0UdbDFcPjbpxH9gxlHIIOc2
P/LSznKSpSFtBYv/Am3qTAdrfxzeZoGidXs0iZiNPlF8/2+gJaZm2QRJh+Dv
DQvJ81PwB6kZu6BUdIcYTO1sIMlAR66evs0SeZHJ6LgnHfeA1I3qGIReS6by
Zx9ArJ2hGxh7SCVelthY0lkLDGhhQG6MXKxanAB2WzH1kKxJsmzAUnroF0zp
QJMzU+T04Dyo4dTmk1lJ1SqijF7EuOEbAGS++GRKNlFtDjErG1lOBAYi+Crx
B2lu7CoqeN1SozGAWCBe0LGo7tA9eQM+eSt2jSr5c+Lv7ywTeFHm4ZbHH4N1
b31zXrNN28Euwby9gwjchrtXeEJwnURDFc0IWAHfkaPGAp/gg+evLDsN9ML+
8YYQBG4WzfRiRvz5+lo44r0ZOwzBS4F63/Wc1kPmf9evVCkJ5DcYPy8pXNnX
sE2r6y2iIHfimi4VHdQCFS0P0wbPMqd15U09fmpJ0tDJtUO4V1HWdbkvz9xQ
wqkmqvMS97GzAlIb0+YE8NxTUBuiFqY2j3RiEywZ76xIrMw5Xa0RcKP4/Eo3
8ZkiIc4dK3RPyta4xsUmD1PwkGoZyx0Z8gXq+QNRYAD2L/y9FU/CsabYbjNM
jdTnPdaUCEKxREDW2jxeE+RgmK0GwhF1PwPC/iEVdtT+NnTQAnbgwIYHpSKH
PgZLcCconyFr0yshw3pZRMfB4HpsuwqyInb5GT5lrz1jJR3tyGcEnxRT+ib0
Z5lajgZcJt+Gp2mRZXaNt0Y8ofSm5LFmHbKlZPv1yuD4D5rel7/04dHXkLzJ
enpeiStAY3Q7nmVA/CqW1EDolmReIa5Qvm/n9nk9PjgdQXd/5dQwtrkECE2M
H/xJmLIcz56ifG8eU/nkOhv1VAfCWTOjhwxT3fMKSIwhrfYVuLCP+WcNW7CJ
U5Jhx79u27bpudiZxO8aRXFX5IbpZBRmJhs9FhzhHbWaxEfI0CAsmQgNtuR4
TiKe9kzUVIxSNYwGT0pptj8H/HXXOXMyQioGnsJpRBSRSUDGbAyTDEJdocmn
4nzQDCfQD7400mijH/DjyrlqK/jDVPlGaosjLTA6lVBXO/KkwaL1FW8ayfpQ
FkN3qUU51txzXMrTClsm1WrdBOA1uPxRZ9eRNFnqofLw9vWx5YS3yJ1ojt8P
U9drcT/PLcXYIyGueFDMboGJQ/qhhpXTdGduiMPPmD3D44SlSIAWkQYIlVda
XOvtnFMBhaOabTUG3wj/NbMzNXUk60PTYXlLea3xLSdfb2QsYWQEt+/oXqFt
Ya5WRBjcitq69/7iqMaD/3d7wwLs6SIl6icX5Ubn+UR7uAF9DNodx/fA4xw/
6Y5V+Tog0vPN/HCSpooHCku1URFp7cpGwI9yTTiKfxs/vhHzXybdwkFbWR1h
mtNILH/Qd473Nj5UxWVrqgXzqNSSXp/igDzOVeyI/Eq8PLFHZuL/Q0l3zHoi
5AnbKZOZMc5p2letTnLGx7asKpQ/7oeBuAroWnKdnVZA8Cej8bkBecyWQc0u
Z+8A+sH2+ExeJnaEOOoT4ZqcRXTdK1NXiQNHSZ4Mbe4t3BYFC9dsqQkBKUtG
ABmx///my8dnW2eJwo8BrkBqpfamh93T2kNXrZnfgTfiIIzKaL94VoryEPuh
OcwszTaO2Z5Z4HXBVJ+phbEpXNwafVHY32DLv4VFTV8nl48zl96v/HR+lYov
x11vPWOlMOmcBsKS3SxjQwMm7/W6HFMjGdXsZ0Lu3bl8n5xC+VxTQu63awmN
2M9vhhL0XikpIyUxyCQXKg8qaeg/MtTJqoMVKPkGGbdohoaMcyCCwD1wIH9K
0Z5FDUDI0qZsg4HA/9bBxSFjwnfCwQju8J4ZUzUDgw6V71E/9o9h1VuSTOZf
b4k0wZhQ/YFd0K1BchodBZPkW63FtCBeam4mZ/2JhRfgJnQjrkKpszl1twp/
aTwoDiJmLPxHpEgmEbcloRnUzjx/We7zAYkQZKrzbhdtfp6S7BCOu7WmJF2Q
DjuRwrhpSzs/j4yV+VUm4Q9ql38Ko+McU1kG0YnyHG7R71bmqVqydrUUgXWE
bKmNP4IHjamc9hWzH8LOS5tjmDKV7woOUTYVbCv1QGF+E9Y451+Yue/CrvvG
r4YCufnwn+/Az+uVpBMlTlQeXZrWu3a8jyQ9i6bzYkINeK1kLZ6zWmKbviiP
rYKRWtzKXxle8aQxFlRZpL7YsBU6k5OHHv4H4uRBgfvak5IvI3+O8BNzSbKE
pPIIvUn/EonSkRMZd7YcV3jUvt5pMbrys+nqASDoZH6JQPhi0CpGY95/PTHc
IgukEkcaBB6mbyUdISPeSoxQ8U6XP3Yu78peR54dxJ1kHosNl8vIYQ2y9WbS
wr8bLFh2h/NASROK86wuX4ORJFs+43ONHHJHnRgngyyPcYaSqDJYOzYKgliQ
DGwUOODV0wmjST9FoPhUGgeATbQsifIfurzc3mJvByS2epaIz6IpJIh0C9Hz
s2IpomYVv4Q6SCVKOZrtUCPjQN1VSyniSA6AS3d7NS8uBhUeaa4lyzrrt98U
LD4x+Inn0o3EaHKpMv7YhyXzp0CjrWr/Hmld7eiZLcDqdjYh1McsCxY6o+ri
9RIEjUbgB0qnVhjVXEyqM4HOVKiPD7rgWpg7Mdqt0xG9NNkliUULe4Q3n9Qo
NVpGfHliQh8D6aT9LjMLcbA1Fdqo23N3+Xnkz/11wNz2bmD88BBJ0H+exSX/
4Z9HkkQ683JVozbg6NBMZ2LmeYeyVlL1zLEngpPQ82VNXdQvcOZn5wht7oXc
QZUsx769MrgdeT0QsX5PH+YD8ROsThZpJfcizQJQvD4Rg7/WvZefi8nf3H59
Fph7y6EUVeYhIUic7EhZ7eOogR7scHbw1ptUMCmAfpVfzi+L5IbKFOSqFsnm
Gbox109SSjkIfgDNNTaSxo7dNKwE1c4QzYc7wquS6w0cOkUsgIiyYY3lQGh+
4D5Dj2NMINdB82/r1k3237OJTpLz9itcvsn5sZkuVzr67ZnrgjGh6wII4O3q
cUimgUaAFvY9k7bxb0dk1sNycPlX+XC99x5ISVMbduOgM5aaai0+La4fno7Z
hfPBnaas+Q6D2+fof/4xuGSmOI9CfzUGOUyqG/+Q5sTz1cJtRzcmLO2zqqBQ
AugU/ldIeNdNwGPnMGxYkr4XX+QnQEICfe6bsJcGADms6Iyxo0lTHegVaz29
RzLy9nuMkIwknfsSdPZWbNN58jq3a68+/XMyhRKAH7R2SF1l0OBkcEsKCikG
VmVlCtt9L+8RFTl8CHmmpFvgjnX0hG5BkhE448B2S8a6HRDQMCsTfsShEPfj
0waJym7iks5DHL9CO4OtRHUOE7AzVrPIRz/MlQiYJ2BKqx96b/8BX+lVljWh
eP371xtaC2i2lIzxHj1H4L8zJ0tLOlgEMGLsKEjX46keU8vcZnu0aeCR70rq
VMP2Djg1hKNMATK3wYUaTBdp+nLZ6f6UnEuZ1MQqocfeZs/l3Kp2fbn/m1ID
ffQUV3HvtOY81fMJkadzFwse+F6fz3rRPSeuHs4Ji23XxHHU94H/+tqht5+I
/dtQJL8GDib6bWb8lwQTfkArVCyeqB3q1lFZSxCTxCnV5jftX4Bac+r3liio
3RvDshT9cFC+NXdDnr8m+szI+aPE769s8fHMGsKMT/+vg5+szg6p3+y9vX6e
dBsDRMBOJ4UoT/ecLZdN7QPnRUCsOUoVDsYKxJRLupDqeYrGArJ50BQVXpXS
thEbDfOcJpidjuwPdrvmMdOhkhEXsXTwWLuvM4WBgkCuOdT8o/QoNjdTR9M+
89bowTt2e6SHV0oUEGPdb3sj9iwxt6+iMcTtRXk3XHHGXpFEIr5wv3L4T5ZE
wNlqcGEmAm5NbtzUgUfPXXJw1hSodwhc/PsJJhc66+xi0pENPQeyRL8ymqnU
2g+/VKL6Q5yaFNE/sIjWK65/KaoLaqkp3fL5bVU7xZvqgjESht/Ffll7JOFR
umPylvLJUEK1Jsi4Q34GhVDMs8kYbP6wCnnqfk/5pl+qXtVvJmPYdZdicmyJ
CpHAyDoScWZp+azJrhq+xeD+5vzf5JCA2wsU3IY4p0R+sZMQROTSLpeqkBlQ
bfH++TN9dn/iHE/p6nFQPfWHDlEUwCk5r0H70jwF1F9uqczXFOdE7eQKwaVV
f/hTN9KzuyWF9f1dBXFI0N8jwQZQHS9kPNbi/H/9hOQLz0ynWHeUpsqDjwsy
l2V+I6bMmQj4ePVa3HewRRYjHhnJEGOT1Y1JceaShhTzTP0pavasTeoq1cxA
MVFcYbZlqPK5JiKkbLb0wu9hJ6NboCumZNMykPjsvdxKyR0Dmi3qPQ1sXzRu
c36rO7R9OF3bDNIsEqpahKgaEHuwKMzrMr1z5S7+yR/sNcHS2FA7PRyqY1Ok
7lmycv0fUZsR1hzdf8TSS9d2OFn7+h2riUk3Ij/1Mco9mj7oVywqrobTIXPE
7tIWdoA0HxnXtJUV8Mg58sXYWmYHJPBokylQMpGzqZ6HFRl7NEhkfw/TwgQX
0oSASKwdNJu0TwlC7chra/eGCtw2oDH7bMdzHUndaZiZCxa/gAgtArTtJTye
2P13umnjrI5PE/7yalI6nUJhRGKKtL7J91BucXX8JWoICXGzil6//LaZZCpy
GqPm1IBThDkNHiQ5qGyo5p93DoC78Mmq3V1KRR67FaFeE/z4YFogZiUm5aeA
ygE7kmB2C4sM0sG3LoZqxRcTfydyAX7tNKOofyQJ6vLCCcfNLhMZxwU4cVql
ZZOulpRLq7E+6uG2CTxa/gW4yIry76evtROiD4XAFxA8NONvIeH8cD6TFNqp
OmHDOK5TXzGsukQ69eXVi76voCeD3SoyWGzSKwaSdc1EJRhoIJLngiMvPRKH
KaSpgS6vOTDBYyw3I+76K3aBGK4Yw/tzmTBQR5CqfwArnZ0ulj4VREjK4ac6
5igepykFKdFteZlN027MSoK+7MS2/Abcx1Fofd00CgnLU/Z989k+R3ARB4gP
C43LXHO13GU9Lvcirb0ccTQSxvj9Q3MC/jeSMcNJpiwH9F7SZfO0Qz+Kl3Ee
ytf2DLZz/jr3QWYlmBKR38ZBqBKpm5BCrAkC3+7oxEz1sb0dNiVRLYKfapi3
PK2m6ZTiY+4lF3ALIhHyVXhAI6dthbT4dlcLPdz93i4ZGKLokq3IFwn+5uCL
NgTi2PGnXw5rjQStd2w7UaJa1dx1KAyFiE3r/H1W2jDNFxISCrO0Z3A/ZCTA
WMWI/qTpqy5iD2kDvS37bn8wS4T0RwSpYLTuBUMhdk5yP588dtASFxtpGkpg
L7Src8fSdzAan4nn5tfMJ5V4vbHEwT+V8QEvpyis9dS9bEeIZzOCh9mogk20
logr783LdLFYg/ywn7980TyXygPD0ZFnYilnj7R9pF/HkY8K1lWTvWyC8ABH
an7WJHqgdwzYVdadS0in5wPXlIZ0pQTSY2etNjZ4DyzxUwSGyzaO/GaVZj0K
Mg3AZISYhBFFKmb0BJjhf0LKxgXzt9QzHiMA2P5lBThwpPlSWbeCyhZ1MoB5
a3sCqB11kkShaP6A/JLmi2IOVJn/Nkk2LmvSAvVRwddLWFUGk6SjAh0MRBOj
l/2suLdp3w6qVNG6uz3jRQaonGCigGPltTcoR6YK6LCM/R1n/QfskBXoe9yM
Yvz2ehRrMr99ZZ38gAXOQ2qq4ZVs8Qt58XGLYPYpRQPlYZ5RimrvCmp+Fbmi
GpC1jTnCmo6o0kdbCpjH08BNEeZI8s8HzmotANUlcXMGM4DgmnGV2Z/3R65y
/MQ6vMDw7W9FskS9Gsq7tvSMa9tcO+54g3mhfvtWCJcAb8T82nlmol5kieCz
NX/7BSMOkLV945fhfVQ56xVHYRe4RnQVpK+bgaFxKSQaAdZnHpEn5D1wkMKR
Z0TerPppk1gKR5L9qfoD8+m78NKBjrQxwFI0lPf6/GakjNqYUHKQ0nAjUo1z
JpcsaBB9rXllE7w9NiMwDBkhE9Xs4U0KTWzFCkFptHrsXcNJthXwNbRsZpKy
cxCEVuo63RmnuI1G4OI1MBUjwXhw7bUV+KkAI14YCOYaW91GsnWJqm8aISRE
lKZ8dEf9pJpWIbxXTy6JbBGA87RET5XA9nLwPkJgIKQDITArgkvPrf4ylYQE
I/+nwnKEsQ7MbGOurcma83D4LADXP0KR40aZZH4Lqp3BLWKVLSbDO6W0caxp
WfhKAr7IcfeJKCTDg0xCNp8k/R4TlYYsjinbhtwLfOoZ3IKJaRCyg1jxBJQQ
mWp39TbPxSP0xfhfTjXTYE3eeKBROUaQXroQpR25ALlvalq9ewH2zmTtq1IO
WvjUCroysbzhgo9FuHoyS5DSNwtW9i3vR3/TiK+pMIK0Wg531UTAM5cZuXbC
oAia7i32+oh/8z1k91aQeCBNPUpWPtLuy4dayzyGf0GZaqo2M1ozt+ZtVM0x
YSlH2V5KSr+OgMe9O3iNFmqTwuKNn8B2Q4etxE29RkFdu5mJ4I1nWxeB/Gj1
xgKxaDszFWXTNFL2F/uis89MsHbd5FBu53O5pYJGJYLLXREsdS7JybOk0buq
OM15AN8px4LfY/uP+2vyHQo2PbYUDpfNxLAtNiPMyjykqZEN77zzXbeD8Gut
p2we9uLOZzlKReyuW5guUuqY4rS5D+yMej7SeQHqlbuLhLpRshYUfx7ninYg
ibjXJkrrUwlox5xPUytWYokMaI1SFu+uSON00Zl5obnRpvNM8oso06ZaWrT4
pAL56S/rRutldxJpPRbe5T4MHxf2JRk7xVtri8GTJAUL46eTLAeS8EI7XTaX
Zj2UZJQmV6EK88duoewlZEPIbQJ/zRLjkrE6r2gbHM7u3+LDIfbtsfwuAYqF
vAumtRSglp0A2/UBFkogXgA8j/2HXzRxfq7gWH3auJkXxHTBX9k0WdYC7eXN
Yd6PmtDze5JD4owt/OvuUEQem6SmzlW09BdvhX58moiuy5/geHwDoMIiYlsu
55EowQp1L4aWIP1Cuww85ge1Of8SwbpzHw1WSit+FL0IyuBwUIK/MsXAkgfp
oSCpQIea9wwztfkEk2hWSz+vyX/exHGcMp5surLIsh1Kr5s2HSARcjQsCh1h
0WO0458AhpsvgFVs2/GWkYVWJO27YBGfhjmx+KcLPbHj4wGyl3qPeBbOCyzv
xlZ2gF4Uw5W47jwPe2jQN4wkKNcV9uv6yi7jbJNKAKbDPxEhrDyV77Wd+gjG
ogTuuNfrQSSYQ5PteRUhtVBTptuBByvBuka+tfZs7gedrEF1pPej47qyGEWs
pcgxyLZ2O+vKVcXRbCY2cMHYm9nnlwN+cZ4BMjLN/28GoH5S1kZiANSgWgVP
GV6sO/xqE/spC7WtAvOmOJ9EnXOSBMCuXlukkzvpiv23v70ZuTLK41LdAxNO
ByIcsUKYsQs6oVwMda9fdInx59JRJ9qZOJoeoEbP0fx8p41E9y9Qn1axCS1o
AyTBWHzPY18DMYNZQLiVVrGtWS0aE/8uwYdL/PmymX65xoUgU33R6zBV6QLf
CBkRKjQthSEs+mZ2AVMYXzLN8H7kSQcTgLso6d1Pmj9mdK1HM+deIgiBemU7
oOgGSLxbS+aej5NMiWnuO4LmWKjSI8+0vtm8uSZbkyW/cnIM4M9KYmWIHMIc
ONFupmY27w9+fFURmChHSyCK8GWWopBTdM/T8Dl8o+NQhePqiZiVhIjBf+G9
oTQX76Exjdn6aix/mDpm89F2NPse41N/znRhdNEL1tjxWnD/l++vcgTQPSxu
pY7A150ChEjPwgwqTPdqaLywj9IOq1bfKBFw7CPdUyOPO0HwMH/yKuJws9K+
AkgeHpIKMavu6/ZabN7UlMxl4P8qe4ds7U1WYoAr4wlJf40upmGoUQiNQ/4P
L//zLb2GZZdbxVPnFakn+ItkKPHB+QJ/jBbFyIoD9nRW5oXNplxS7RF5EDou
Rcu0FYHdm/KNdGnNMV4+m1dkB0UNW22meIje1BaAmmaJ7NhmvbQSLFhKqkOd
OxgvwBtOeZJ7VpJbw04q+Y4nuf6dPliEumWFIc6rPJ420DqINe8Vb18KtYDA
taUVKJq3Y0IYexl4KuUILM91zC8y0QedLW+DXJI3SDMzMmKMPs2xqqYjgn1R
mIG6eOfOdwc915860f4ZELWVADVMDfSNJBCApZ/ZX2Agqx5mu/6xQiZm5DGx
pj7AVwLz3hCcM5KnFHLw1GjR+soVUwP7picWX8Ed6S0gn6AsJmvWdGtYvX30
weE83dPyopxvCrU2uHrFa4vrGwP5D5LMuU7Tn8uvXsRMkNza2y94BPhXLD1F
y3Kk4e6mWNu9HbB4KVEj9ZjcwUY9g6CYQTSyqUaz2/T4PvP2NRfLaG/bKxxB
6i+ifsiyDTlZDixoEP+4MBZkYwbttiSi8GpHDKBe05xbXEEOubbmvULIeu1z
sqP3sgjJIq6qrxcn7Bs2vi23XgpTERjWCi1R1bXfrQZh6Qt5nr7dP830pCM7
YvuqmNcNpU78BCqmIsin7s3AhTStS65aTH17y4dm5BtalbBaVs+22vawZ9Zo
eBSHR9KRr1Mr/Y3Mf24UUQwdQWSd/EkV8OsAhsJil/KZRsZMb+a3KORZp4I7
JZ2mT1qcACUPi9H8sgFdbGwpYzk/o+ePlW/Be673d4sPWa2CXgg0WZL90ewe
COuv/x01rYHbVmkA5btf72pxDrf/6GK9rl7Lfdx8c0FnBQzCjr1psO4DO0mn
laao+dul1nLE54SM2hbNPpnvRP0DOdOqvXF3PZ9qylPSNuYa6F+Dihrb/UU2
rVhEEMx9TwwJDZKnL4IU341byUgR5LI8c7uca88wlKCQnEzXES55ybu0tUkD
rHz7jPNWpud1ONIsm7/Ltx1zBnJlsvUp6CHg3WoK5M0zKyeSQkCmInIuVH4L
O/NrO3XtxfFGIzl4corhjonvybUvv3eLxBDOSiISOFBGyd4CBTPu1TocJLSO
99mCRV2XuRHdcw1KWNb7YfmL8b1XofS80UItZDRMeXUClMgTS/zr1K9j5Iqa
xUc5y5EVlufGEfNzm7k9R74RAuz1HClsr7Ymp43JqDzVoGxfRH7IP29qu2Wc
/goRgfFKwwTzjoh+RLbo8Qtg83Tbd94/TDLDAaZOsyFu9er1KTwVcF7V0RU1
mpypFXVqXLzv2hGalWZseDdRyFDX6fMHEv310dtPUJ8M3rpZ6zD44cvrm5YY
ZqOGEc8R2MbzLVeIhRIV+n171JNTfiPIVzd86QR+YKfrrnqSMWHfQNiJyIAz
k6JV5nP1bBx5DktjJezMdwsFyHrAVIhDGB75erFUAJUZCiPTJ9kiaLll6ocr
kYbglLQkn4gHpOQqbhdbwx6Z2Zd09nlbe79b2kKURWfSCzgUcLG5wZWOZ3Fk
1v/wTBtSc+xrGrLLS6tGa14xp07/cRTc0rMvqaQGR3uJ0N7OyFI8OfXn82Rd
xeKy4oPXXkKzxG7qKXgUebZMavkelopKYot2ijrKn0+nPBFYqcSLAfbTuEWv
Kcg7oH95m2Nq97Cq7lSuLGy8lY8zy3YXz6J7bL2/oQ5iog+CsQ8IaIczfnyN
MV29pZpMBkrLMn7nQXrvqt8b5G7VFsdtiskTPHRzbgqKOVfnU8Al4oNx2d2r
qwyZxrepFjMdgMZbhEaJeeodCs9JxSVzrQzP/NJmVN7t9SwK+W0FxOGIVkVU
MV75I7PGUDkf6FsHi2xv7FL/AbTeua4DUFntHWunDiiJwALwq7KqPsHs7+q+
wX+n75MBH5BGONvnkCP5RhwO08s/LCJo/w8tY9LQDMG+KdFECr20JARSc2RV
vrE+1cKTvMrJk2mpnUCYlwxpMPeSAFtSerPFsUdZ4iXa+Y9yhVq5zPbSbccH
6Ss+Mbmsbe0n0MGyE86ezoYtQsGwioOgu8yWYnxJQaiH+l0S7VL5S9nBVunX
7Pwo5PxcVnZqiMigu8U2okBTHUuLe7bfexKRQRndx2ajcsOW7qdidh1VBlVE
BuuThaXxeoYgkebNxZRp0AG1yYrV7YLc+YI4vZp+bkLy8npOHcAXMfkrN+eG
IBmB/83D1u+qrULbOagxCZ7n9dXLcki6r+ATkXDPUpLO7bqWtSvPevcMvzFH
0XaT28gpxzr4HB3wn7FGrcQ5b0KLZqm1JplLdGCN7F09WoFggCjuUiT5sMN9
KRXHms0jEwYDH8fhzW2YK7HPB3pIFXXLunAj4CmyKmPQuMJBj8ik3ZMOluBe
4rhhTYo/SkKQ9kg7bnkyJbKgqrurgxxsayq5ZrKvuqMtk22joxzjUuAGx96B
SeA+JwNodFiuSN+dmiegZq5o0FrLfhf/ISy+AC2ctyqQYuUA+7CInr+/PXGm
lNA7eNVgGOH9JhvTfcrLOfxCHjEyQw7eVhwqwO1HL3jAa9mWV8kOQR/ySTRy
ZyaaOoUD2x9CtRCKUlwjmnrJwvEtRiT/aL2V+jl1EPWqtTZ2hmTnJlvH8+Y8
TtJkPDBcz+/jzFDyBE94+M99fZ4A+GzNh7sl2kVyQx41qW7+wi9ZsEU6tdFI
NEPyVpHYO82EJYv292Z9W0XAS532POkrErfHbRa3adPMYPfu9PBaQe49ptem
WITbbLoVsK8SWzWmGnZDoExiC+k9+n92yw/fRoKE/MQ+8csGNK2uhXOhW+lX
iqeuZhgIycO914PZ9cdfMHgjJXkLvp/QpW4Qd+WI5+1DUDHNMCZWaN0h4hYy
E2E1KBQnYK8qSiGzpQ1g4mZLcCul1Nfm2Xh0ZA+zo8cYMlm7y6MGbpJsRG/c
/pWSRtDGnlgqZTZK6QwIBYMW4OK+svnVBqt5sp8jcSMmSZ87FYyYzgTJ9gX7
WmhLnzLwyffDAj8KD7gn+W52D7NbSJnCZSw/+pnWuahKB10P6+PvxV3aeSbz
w2Nzm9APBe9R1wKQuLIPQK6rKdELlACmAFhqRC0q+GMRZy9e5ZNu9jCLn62Z
zyZbSeGORpZNTldEU4JI5OCswbVm+zC114XghKKsKQVmRhDy/lg27wKV3WUh
wjzoXl6IO0tsjxq8wwpVScaWYDhe8mT/Cm4SrQp6BIkkjn1OgUsdOP3kpG9U
8NirkjDbDR2AGIoNPcghkM7eyHgMvrZIfo9tJqNdhOQ6Ema11btLr6Le7sF2
ZFkYk+8X7S6g8Prsihp6ZFdAoa6/ypOUEhwpB1UCuAqjM0LlC+6Yh+O0eyOj
3kXkyJsO0N5p/p/YNltNytTeITyKyR1N14dxBzOfHjQz6az7PT6REJ908Ezh
eHKJQnr9Q/+8TTJC9gzNMjSvHqeDOjiNgYvAuw7NlPvvPrk7jqKvdOh1GAjx
lKdx9/B8otTDKB4NCMe4czq98g1VQPCHwMP9mjnJ/LJlFsFozsCaxFX9WQYy
hybJhrlDbMrpsn9xQYkynPjAo4czMsxr8MXP5fC0T6vQKUHA8RwQpgk0c5Pm
emt4pjPtMwGFDX0q9pUuMpYE4GwbWfwJ59myKn9SqZKxJlhzDCg1P2ldXh5Z
oiDVWEWzAumNnBI9shy+J4wE7GZy6dQQtKlLHF8p75oHCN7+l1T86zeRP2NB
+LncKzzLsb2BAnxmgAuqrhnJVgjy/aXFug2X9OsQ9srcO8p9ari4sOIVTEq7
nlSY44WP5JH/LTXb7o6UOjLd0y0obOEE61yBg5ibRK2JNAhOAEUbQdfdr3Dn
sX/zap9vXUPtx0N5814m/hZnA/wwgDNma96GaYJS7hEAbLRkzTLPEQPzmibs
3XelSOecjhUIPPasxaeP3BcOoN4Ox4uuC3aHrrKCjJf2IwY9H+vmqlvFbVts
8N/JBLMvi7AtaNvPFyFAWXUN/9Uv87CBHIRIs9pgJPLEEgccopvmrqiGz74A
EHkWYRTwTW4dNeROA0qHlseRUpmI7HNWr1x7wm+Qh85I1273SYEhb+WXDGqc
vsTVWQ1glUkwqkLMVe/oROtw+QF7te9iFcGFlCdLLSUDyc8pquOB0/h65BLa
IRAaEiwfk+KvCVjCE6r5bIgvJZjywjxBAjSA1qFMYVWLCM/QQNKMo9RGgI6h
ITcQHs0U4EqFlcyBhczrLmlzgXRiygfELxrDANwMtfBeeoukWUFB4QSJrxmT
8Xnrp0e7Jkwttjlcw0t+kN/Ctd8PVqdhslQEyKfrQ2CKmPlf6Q7mLGrz36so
YO4hspBcCQPVsuGkY7uASZK+cfWzzNB7m0YBOGGLH6k210M7N5agE4RBXYZ9
HLn62fgSUUjsDnCATuxeRhCLCiw+HyeVr0oCJ577XGzBjGbm1Q0P0zlMypNT
g1BacwNUBz0RLMNeuXFPWeDUNDOFUkTLtHMEg5KjZIBLVkidzKbPXm3wpyNj
whoouZw83n0i0Kq/W854D5P/DaYIRf+nksXDg6af3GhMI6fAyVDzWfzIYLIg
tPB6qwN6s0ca2/nwj8YS7FQ3UMkOeNvjvblcYQWhzb792XQq4X6lCLLd09kD
lqUCVGBvRr/CvQeFicarbWEoWPDjqFgdT0n92lnp9DNG0sFo2AF6Q7t+KX+2
/A2bCMkLftpGQOGf3H+z9bzPF4I311y14MXvuQIjwk+nYI+tpNP7j27Tcrml
UiF+HBuaOqiPwNPQNCvqKuAHnCh5lSmX/irt4bDle+3SQimxk+zC0Sy9HxEq
c37lLWvIZg2hbcQewcMBFv8u9Y4YFJmAXHLJfcOVG74yI0g8QQ6xuRAUVlLo
UIXJjVDP9IIjl7A1KaPibrqXbnm32NYDiHHzTiUzD96gA4F5iNCF9rH8KHSJ
HTfQBaqwkQVRtauR9ciE02VMVuy+KcwU/ic2E5Om1iQr8Xdvj738FaPnPrKt
ov6UiNStDCOm+OpXN26BbtlONNoFXMvNfcEi4Hnpzml8E3C5k7LV2UD6tuhI
boTQS2ZeQL84hHLGWPd7ZDlk+UCDnN7GGZWaLOIwrAkEfr2WuLK2nX6YSSHm
Uw6QJvMAt55TIRP+oCwMTCgbPhl5+g9tbJ3/x3t2tXIc/GJtcjBfCUDV2Hkt
4sTBRtegEeWTHOufdAx2vphK0Fo2bwoYDufn0mfi9BdCQlVsAcoinXovOc4K
NiI58JWeTZaO0eG6NcjJb0sQVOrwsZjycIzwDTr/hq4ZgbWo7EWQRqUMw0ZQ
8pPmr0hvcP6sXwgCJ97f3E9SHuwzDSJEdpmxYZFBKCSY57SO7pHxXOzbKhSu
b4d3LnIPPXqEwGxOy6q7jP+qLOAQey35Q8t+2Fdxc8ev+W5367H+uM1cj0Sr
5PYvcJDincVURzJrMN1XYmzie+SFRx2nAR6xh1ouhPnC6hEI4tLmxnoanj1r
1/+OFySe+SCPxcYlhdmN1dTPd5kChPbn9v3H6n1s8QvuAsXmwaSrnm3WhOMO
JLBJfguiNdpURT3NIj1KGuE+kMYDNmzgdKIP9WfcHTtxExcRbdQC7cXVW6am
0HaCvrF9n6ca4Svj9zI84Nv2yWdgJMDR2C8bfqlgiTOyshZNMlTjjWDoa7Pw
Yzev+6+/qZju3sBPU6oROZskVMaRXkg6LI1YSbZob7K8i7/Da946yAPDQwAT
6EzGx3VTvTqLLb4UZAeScW54N1Z8vTvw5cHQQvysS+Pkd8V/cLFlHbszHXPa
QnHqSwS0RPw/FN90/6UlUQrLDE4AGJAmoHFrYiTUAwJHtKsg0Bemebum+T8+
uJF6BXlYQAvuM52vsjFDWgjkaQ+pHA1goyci7JX5gb/6eQQ68p0Yd9i6Z40J
vPoXmgeC5VcF77uFjoyS3oR6PJptUMFVBjSmQ4bo1gO4xgzq33hsKO29tiMy
75EM/ecvxWSwjm4w7gR3EC+gjhiAe0GeYZYJkKf3vWQaP4gfPv0j9ys5L1F5
j8vHw3twXFESbVI/+zTEiWuqGEnC+DFOx/+hYCqcx8fVymFJvnmfvAb+BqvZ
JVzQoNnnnKpzyLq6Y+B7lZj9o0u/65Z8tkI7j3tWEMfg6b15kcPdi3pzfKVF
yVAh1Ss0LkdyqpGzTfL4qoWnel9kKaLTNPczwCyNzdVm/nL8XeYc1LjxobWQ
yPG5hLv4Rhjy3k+kbm1ucZyHGUD5JwTZ2+Zb7QsjzSmQkyBTs/9qyjO7deUj
iNGbIVmx2YC/Y/sW4+nzmYC8g2bNtXSSsnrovXk0qy2b5NrYbmhxx1xOOYaZ
eJvuNnY/g5Nv34LRylg/MPWBkPduz2n7u9p3DuMLG+wtRKEgA/+p4fbh7dJZ
oAIUYT788GrFXxwVG7TDPhE30UTzgn9k5ycUZsMagzrQTusbfMHQPEBwCEtP
uG+OX7D4/76E6H/unperHQgUkzJjV1x4cSYJc6Y0BcoUjKb9YK/VG0esoiuf
wdvO5WosnwKeDrvmhWppMqBLu+NiCmSZlZmM5hCbufDAM2JTnWiHi9JvA5+W
UtHRlAhKfs9LpjwCOgyuNm6uEsO41Aed9bUnL8qLyVDLF5x/Y5NCf9f6d5t9
dYGgGaIuKjlZ+JzMeFYHcnVuOlAPYQ56sTszlnkM286phpO/webm3rh0j6Qo
/o0eL2ygkE/Th7S6lhlYQobbGLnO7RLDHjKIYcghXhp10NoPZIBsSOTsReWR
TG31fs5m/k2pftcUoE6IuIXBNM5p32ihAP/qy+0O7umyKr22hXaMvaO6Qx1A
hfMe9M+WD6ujSDI3E4+xyuVepTktqpl0AYiZBLHsrue6HWLxgrUOl0AxSbhb
gQ76enLA6dJ9JVu1LbOEkMxAOxElmIr+diWN39SkukjOautmYnqJ2w26iPlx
Mdclh+4e3qEG7mbYFp8ZHdXCgKPlokswbaMejegpnYGEJwDm7PButMadU07F
ZQ1hlprJgZTTOZW5sq4BPh3aW6aR6nqIv2kq1c+FWJIw8OpbS3NgnMfHfbXk
5xO5VqMaUtJP4OrJPWW46EnSk5227nFukK4tk283fjPyF1H+C8N7aoq+Or/N
U4CcRPjBACVMB5X91il/prEwE0knBbsqlKLjxAYiZOiFl2GxoQFgImF01+UE
VWt2SwQtsJaX+1mwaLVn3RqaSrq37reBAle0qlwr/T7GElDekF0ekm02iZZJ
AGlgS+/XRy1ETpWkJRQA4fkSBE0vhXhSi3+5M9kg7+n6D83PrDcwoaPhRrs0
Ow/hT05FixFo2LPM0naTjs897IeL+3w9IwxCArTIeFIxYUj09YYMXhplgVBn
KDQVVTKHPf45S7blRUlKJxivyBVHWgB7b8YcDrcZevho5H20L8hoSVGcDpbz
1x66dvb1R8zimYrN+S956JWWMO/sDInQTDWoVZRkyirxQEMlVEqZz9NKBFOx
0UPSX64UsKPwg6eZkE/z95fEyrpdycC/Jywh4uxmiQ/Ha+X7VMJ8Yrs4WuGL
7inMbHVHKcy0z5Ws5qkwriRblWGTbut+woykHtELcTzzHt7OLo8f6hd7AnSJ
GpuFFEEIOcvO2QZQ+bx7W+huF6n4R6tHKqCotKn3XdM3ivM8gguS5gU5x9L4
LSXQF5vvxYWePkQksxIvsG6vVwBz0QOS7F3OxkTnXtmRwtavXyvDuuNgbvYu
6EAtxRGwy7/wJJ8onW7sJVLOxrUnjJsp+KW3NaY6b7waXkGOdsypzvICLLem
9vJgiMKJc8g40gfTnXdIeBSHGu8TqcPh8iF0CFphCBSTxZCwBzplp+M8IPvo
tG5MADgZCFxHTTNTDcjoj5JVXtaJfUbQlG1/BlWL+vfQ8QaPamqz0WJQ+13e
iaCNLh5Kzxghp+9eey52dovMSDQ3suDCHdMdHVl7BziEOBK7N9H8SdMg7P5z
qV7sZSJQriuheMFuEWQoAlzCY7taffqpyKNd4fb6VhEo91Y+eA3rQbNH6cul
mP78xS1lINbBb+HcxJaRWwIWkVjdiHBzJXwS/97D/gHNHaG7NvBYbEbUQ9FN
+tFSQXHIJW8Dtfz1G2GHERja9XvIPonctAkgfHbpCAtj9M4MwzbqIYIt+A5O
GSMS6KZ51/uc3VWW2VPyimsofs1J6/zf3/yKVUS+y2ZydFnyXu+X0dzP9z/n
M6r5au4YZBAAgICC8c6J4h95uHkQXcj1vXkNcwoNElKEiXvy8FN/p52cnhbh
vlhgHJ/YHLIAvv+BJCgO4U28KkFeoWTncIRZ2pKNNDup852K7mSGYniEIIoG
OEA35+HBOaqKMyMIhvKl+6q6pYwAHeDWjoNW33JlMsbWCzwBef6q8GYogrsa
yYE2VCs5Yv+FQzDoRlDG5rLIO28zMsJFj7Z9Y0SacGHB4ntq8WJI4Hz6aLY7
M8WI9JiBteza3Co7l0Y+SX+v9BZpRky1p8BhMWVT6CP3y5RNqNuhFnzw/bkn
t/gk7pU/xYGLy+GUfdNLn40kTPiY1wWFfZEPd1O2LYD2UboEzOqVSJgEdrE/
nJkDCXxp9sloXAgkqBVlYILZY7B4NHZz8Sb1Twx/kZtH9irZDyNBDLdqAyis
weNpyIJrsMmJxjmClo/+NNpq4FXvJViqRH+j+EOuMj+9/gr2H1ajONvGx5dw
X64EOmNy2SiTf3VhQaqZZ3uzTfkOTAYVO+wYq854QsBUd0zZR50ztJsf+pp2
uE4HWu7v66Qo+Z/6cUVHjBH3z6/dwI7DLdijAdfTF7QJygEWfqbdW/Mc9KH2
kW791X0W9pvWbPibeHDhBnlQpWikoPbIEfqXAU0foWEoRF8fbSSuap8eUia1
CRBZ4KaeXkuMeErQmYiIeITwwrI0wvIYIjWUhFZzlSEwGYBlRf6RiHVnAHRx
/v6XvBrgjleZQ6Rdvvr6n+nV8hdvgKXXO0lpIXr0gSbc6pxHacsYOzeFycQ/
4ezSzZ7Vk5SN41JY9uTVgpm3wQZ2mpgsMb9ZbJb8guIQ6eKqBCnK76ctEszU
C5xH7rB+p+sN+LL0wNpF+eblx4w73fM+FZMFjRbB4l/o6Z0zjsLjYm+bhHQU
41xFHFvbXgOgUdFFYQir4yTozDT9BL1saKZ/vRFJLuPlw13AAu6R+xi29jnz
GUZCEV1x0tTwtJpW7yW4QrMUo+GQtkmgPDOzEzFrtf+a6e37V5n6wJ8RMrdi
qiFapPeFl684lCzES/bBIkpRqv6G95aajCoa3/zB0yxSfjD8S0FBB+mt3YcT
UuiGERfB1tJR81mfeQz93ILPIru4j9X+i4FzxtX8qWzvqR7Hct6SLEBzPRFY
/uigYROd/KwE/UCVaJhAPhG9x/3mERVLUj/xymh/YW6WXbxor+2UEQDj3pma
/3mFp+auHpBxgJJhwG4PF1D9NSgQCdm2uCOcnpRIZ9qWRXRx9TAuoo0omcKV
56Yq1+6tW97yR/w7llXAYLCLZhGIfVseyitxvLze6Inbxuu4o5iAS6/ZeGbP
+Waop/y/ToYjUeBXnTWXxg846J5K4CAmycuI53Qe61yZ/v8b5+q7dR9S4NRI
NJLu/9ll+CRiurBad4+AxzxcKVFV8h9IpUfEIMP8FlcsXJjxV6hGWX4jVq1/
ZgoXDAvJVkg3DokDTKpBdbwbcI0XZyS+Y9kAYY0CWgW2pZK44BUpZtvaKx6n
sy95cR7/YaiiISRb4vypIRV9auS6WAIiLu/ynMe5XHCj9Aujg0+VcKAChZjz
9lEoXdcAeStl1TLkkSi5li898kaBzHbppl0xReANQzt3uVGay+fpq25zqffU
CKdwr9ae9Ht2F7iPnVOHtvCaulY2h2crckhQTVQpJfKkIDJOgDSBKIcneCn9
cJ45o3Pj1I4azCxkn+NGfzQRFExaUJrDXOJ/HMdNgE3zkcODvklfdRx8eGOM
laL8qTK/KluZ1k3IfkaigLU8Km55Q3YUN+o4my419YNd+iMD6JKxI5vcLxrd
CSmadt7CpIr8u8phGTB3JDOpqoiC5isTUxAzNpUHnoJq3uKUmcpEWzO2tYw3
e61FD/4V8Zlg4JC+R84CnFB49v73S5a4D3ZkqS1qQVzjS8pyr/eGZ1KD4CTU
Pa7PuoP96N0Axf91pXbLyMK7oCg2JlNcapmpUf1dQXau8lSUEcS286YgprXu
QmNNlsEmnXB+Dj8+ram2ssGI/LrBUqdWZwiWHrGDDzZBLO9YfTL6qrt4Wlvl
dezy8pQqW8LtbSIAMUq/BwGkYMP0pnWPcuWRg/aHW4MBQiDb+xWwlffxiwYj
eED5gpNWhpksZAwhSuP2b1NxZr5GYTQ2SE7Sm1A00PBxA5U1lw/WIdc1wpMi
cORnCilvXnFwoR5gb2MiXWtQ2HTobs5t/UZBSQLnuivna82WZbOouelORPXQ
ryHeARRSjyWaZFkFciRZDYGAya53NLxTermR5hm4AUp4b9yqI6sr+65nWrX3
a7nmAu8kypfLOsaa/gwzrk7jw+wD27Zv7mkSNqCh0BbgjKIbyLMG12NKOvu6
LJJ3oVCZqXpztqD0rXpbwSRlrrjN4NGM222Y6zG6a4tmGaDefBK+4MgGQn8S
jK/3i3z2GR5C876fynDm2LqaKZtVEsdNZOrtxqXhPZtXuUuIb3abrtL9/XZR
rgcUMGGgpe9cF1MmM9dX0Lt1rurcBDyb8/z2Ei4vrQ7s9Gw9UkO6dsVS/skV
PdStFCjaPoX+HUp7CSxxhPS92CE9jPdOjWPr+i9QbVeJRwj62cjL6JsO7zeg
ybQxzPuXfA0LDb5efG4kjiiDFldt6a0j3esU++qiZBEXS7949PA8DeXEjIaK
/9hh8YZiIxyUgha8SCpLsMjkBdFhUcQ5aBzUhEQrmrkEsZW3Fo8TrtH00RJR
hxsfIdinxU659IClbWsywbYocOtPx3jLZgUdj0jqtWpg4zclvnmEsDHUMv9W
NBM3Y4p9kHSaAWhBe1wEsadILEsyPIz2mAGm7nnxjiJMOVbtMw7lqSWOAuhS
B0/lYCg2ElBHZeO+zKwLUrL4q7gfnhYwrV1Ik7HcBZmFtAzjy+ZtiZf5qNuh
fW8cGHILH94IFAXwMKMp9rnCl3WZQlZ2uxWPas3IDtQqaEz93jRQnaAAQ/9y
VvXFIjGktwPt+AfaOpFAJUx6gwhcioRV8B5J8YL/KGd62VZzbGPnTfLViGFQ
FBYXi4n/bU0SpXcAX5hRojtejeUlaVMzSL1PMVaSh1q9+phNcX1nFQVUFalW
veAn/DVZeveo3ZB/+XC4maQQgkC53lCSjR2PSeYb95LBYksH/fTF9VT/WqTJ
q9CgYzBW4Q5QWcasaKMpyWA7tKy0kIsOj8pcIPUZRpNTNZ3uW9a5uma6hpSE
o2w/imWjiXxLdbjg7O5IYgv/FVr2TGcm8Cl0q1uCZN7OJL8nW1E4sJlA8Xh7
JkmIfYva1ZS4U6UUK525XdfqeI4WeTZFmGlmrlNroHDbXWvILMGWBLQ8T8ss
ZqS+fkPjNzWHWPhe+6v/5R0/1rlqBYuKF2QFO1nPAcj5PwXIB6RBVaUWCYXQ
+YaBsqUFi79zdhPCNxh+p3WGYhtqsAuhlUR8hcYFB9IfxH+5qKCXhpqSsC4r
0Ct4xMl50SISNYtCBfL1NoOqjkIb+nmQoWVoQZ6hK8rt8TelR6uUa4d0BLmj
z+K1xR+AJ7XCCmebEX5Wu7ozjoWN/WcL3ET1/Z1jrUzqrJZuuoTJr3A18Rp4
wh5a3JH1ddoZlO4JReMKGdw58w2g2UxIsuj+ZDOPIcmFjazSBw3OEHhpVL95
ZrVqnQaZUwBVJRZ1poOb8uLqzJXG5oQTjQYeUNVF6Vea30Z0vkN8E0QYWeHB
Csv6vG4IbtrEcz28TG6CY8abDzd5UDZIrm91bf3hBUxES0PZb7jVIzgZypoz
PpY6yxbQRv0yET644yjWEt2TbN7aFBMwOHbysOOlkoviEQIeiLzbrYiwGZHF
BUrm1yo/efZmVMQ0fq778eLFHAwHTZyhXRh8xLXaSb8BRGGg1/5wj74HQJCg
kNHPTwS4ttsYxPuZ8tNjrHQjiX/t/QPovRaocYEePBZWKXvsLEFVWC+jHwku
nC9Q+eOlQdF6jkLD63rIs9uHTs60hR6JWmXFjvlyZdV5EVNsmBXE3F7TliaD
8RD7+hmVtyRi24est5SfX4TBWnRKvuYl/wKxsBUxWVoJhscSvo8d4MAf955B
xsRF8aUuxlG/XjcQ95MRC3UaJLI4xNr3wt0RVF5OmaZdcKOdnSkjJFFprsbC
nuwlwVVp4VZysLyigIUudUhcvfCuNdftDGlKHT7AHaN5PC1URR3Xse8MWQfN
4mE2AslWzeOY1nXONrzUTx8EhQBIGbTrVgFPSSPMLP90OL+O+EHQKIGXOHLA
Szv8379/RJILkmBCj1CP6jSgGh91C0UnzdfpsEEefIXJNBFvFdK3AAOhgByD
i9FQM4MWc1kVdr+x0nndLUJVacP0znrMXAJkQvp69PAf02bmeihPGi7qj8Md
4dpQU6YgBgQkNtcRN2W9EvoBI+lGT4JcYcIeIfuV6RDRZW8ftTjXVL+IFhLz
VTv4sAms8CD6iotbzA99EAamdl2rE6Py3AtcOmIZILpJjZ4oW47oLxq++uUL
N529hTGbS6qnIumpb62BGi11fKGhSK/pR8MBg7sC7uP8EZ/2TSKIaSGAJX6b
TenfgzzT8gt67y1a+1C4N5VSQmq6eDkCdnmQvFaG0BI9tRg9bjeIStZqvyN2
aFAsF9U41/VfBtwu2JAhxEMdUKAm4uZswquwmqer/WjUObpbZhhVs6YhmT2Q
p2rZ09CT2EO8FE1ZKpjBZAC+r7hKQBtkWq6QLgzTtbZUh1gxEiW9TbMT5/9r
M/dJ3MPRN+n2ucqqTwbGmTYT5JzujP30WyrD4ZkV2+3TiChQTPp8i3/OVkA0
4UGZGUHhYcxdwIXNFuPTdsGPvkuJy32bvJYZbIYoch2Edl79gSjZitcQkqvm
hhgwBHgUNfMdntXanNwVYlI3T3ijBlUE5iQNOkfiXb5N03bZEXZhhR0uljnE
rlEr7jusrb+JYSZrW6aRtfzdXUtswu55liZsUd6woq/aLlk3DNCHFiGRNpgd
5eqZmdASRD3ciBL+m5Eh5pT6qA126MwzAr9eBqXGLjikrUm7wVuxMXAddFOy
zyRLuWTGK0YEKGA5sgpwvvaWCb7frb/VC45ZJIk/HnZluSGDzlI0Hdxcis/t
qwGFSgJqET8j2Hx1Fzb2L9H7aGT/o3Ze7ReymaKGITWxnpdBZELUNmUiuXBm
M3WsFn2dWI6mNspFm0jpGhK9Top0H6m8TEllXBGFeQz0FroG46ojpvv8Rd4N
oIeHcMVWCXWohqqaz/ouv3cLvdEBn4r6BV8ohi2HKRbxvUP1mbqI5LEubRtg
lde0BjPcq71JbbuWvTZWwLSlOGgWBtzrRc57l/tXsAL4fowwkP+pCbKKGu3p
S7wp3eAGxqeP6VVQbyhgkRezPVJGBiNIg4tr/8p+Hu4dH3Z2+g+Qa5cqcg12
9r1RKPtwLR0eVMYPvcePODclxo1D3pVZCszX1vbl7AkR7NYreNAHM5b6KjgQ
ZKwVner6QOazVzAfn6WPC2LpJWgPTP2j2xcz93rNBnsQJRRmWEsrYjyPDKva
lmLpIzILv210ijpDll3nDj0KNjf5qBOiIE5qWjCBY/BL2KXH/V0cGwMItPS7
11KVO64ddNtUlVjtdj0zLIIoQWeACawwXKzCLoT263mh1IEbat9F+wtyottr
NEXc0oBHMWDBT+Wy8g8K+iH49kX1R3XbncAEx2rnPCXTNueKpjo9Pue18ILc
ttfjwo0bv7bv0RIHFPRW2wrslI0nYez6Uru7Qe/foTKAVgNnwe7nn3h/hx3r
5OWQMPvSz/z6cVu+k3ODFuGg8KL4BuLvhM7OO3i4VjewDLDsoNSJIkACXJUA
yF5Rfsdpmf+mYY6Kaz+LUDxR2OnlYSoS05bmN9yUSAmak0zhY+kR43d68/z8
xlV68rns5PB5T+gwqegpdsBcCLS8qVGB2qix8etAndz00MOUKwlB5DxGORUq
UudeEqjoaC7UeaoNZk0spa4HAMZmfKDTujwTuG2auYhHQvfc37oFHOWl2JsQ
7Z4nJwB3eAwxkKqypNAAi0hMEqggDu/PJjRIbifXQ8GkaQRmmrfMiy9DTwuR
gbTK+iMH8RjGJDucocHWLxEhcmU6/rCKm/ql/YUyM1BrKNfRIf23QJzNPh2t
1H1bDK1514S/doOjC1UT1AKWiBTMCMY0DMe0kk9drDrMkuVGfC8jHNNkREa7
BONobha2QUd3nNGJxrQ7AxLGpaHfvg4VFHJR5Ok/j2Fs2jAoQDIBcvm38vnO
yMzW82//yuwFNQGxg/fbXpZbIv4Kh8FZjsGcCHGK1ItsqoDRkXHhD3aSPMHM
UYkFwyYg60QAGIk33QGc0Sv8qlBh/FOyXqOV+dix5z15AlYpHre2AaQtV4fk
fl3G3ScKnxLjPByYEYVnMwvoYVKaC8rRh8KjRqvOz0oGpEQEYTAuP3JxIo/3
VTG2WJRMLKAvlExPjHY3q8cimjdDXF2AzlWlQmgA5LJ3oAoVaVa9gKFgQa/u
AW9CSOu66/dtUKeUzw9P92WOUat4HxFHWyyx2l84O8IoTACgOZSARPf6uxTE
C1w0NfSQ8DBffa/EGnQkVzl/frNeiqj5SuzmILihbIgRL30BzhMLloQqNdOG
qF/Ka5KShGUQp1bOz2CSskSat3w7PCntXJAncek7T3rnGNRBWEiT/ky+k+2k
kox09qxQij3Ds9cEaU5efTJdkyVlINkqK/QH0qNfAhUaQxYr+5sCiY8qtgra
yCpOfEShMYeh/PZcymJbJHE6usaRF0xNM1TAFJYWN/kY+kpAAj7dICxHJJdU
/ORKKSGLiTt6IIsqBRCfT3aYH7gYjYF9zmrdcMBoSlBeoimbpnRljA7OVgfM
SojPXl8dg3mrqC8Rfbfv7vFlh1UbTJp5YA3ZR6HT+YpDdlGEw4gv5qKtcdzG
vEIE0a42GQmeeE2nJ2cVPtz4Vlwl/hlSudZ67HHsDolFYpbYqWQ0Q58/rzpi
a2Z+ewxinmthcQOte0jWNdMDXj4PW11TXN2Ix0gMlWUGG3tbtR8PjUBhBnAy
A5LtihEJ7PzYj8Z5P+E7NLC6eOiVNbZOpRfkw9dpW8FTjhrr3w6szFFf6U5S
ygjngbjg1xd6C9yiNIkcLCJC9rVz+j6uthD4N2ovKiJSJzTpXpA9iy4/coTs
8/pqIMGFGIkuN+Bx6OINmbLplveZBauvgk1SVTn6OxpCyYyU/nLZgE8pkJrA
ToezYrVV1tknV6mMK8n+3jdFI1YJoegammmIRVYfMYD5v3Dh4R61jVzq2DLs
QImt8UevUdsb4/7urx3eFMJLJkHKJnpDkVUX6N0pycn4X1RZfrmv363sTylh
MkcfUffAGvh+d4RtGx0iICQQPk10YYmfclVNJktThWmHU4ALwYN6E72f30at
D8DCTc+FOy0iqx796u2neLMjYTuvc4MoA17L1KWUHWYu1S2SwEWEMMd/uAhd
TzMsnqJqQTgMo0sBk3bJFWrxRgy954f3Z2oBr5OnFnvJ4wdCbvX93E75RFBk
v+jEEP7LlSHjm6OZBqyvxC9T4HqLWzDX5kwR1N3bGOxRh/ZEUuwjN6Pp5wZR
bfWe7dGyW+NBi1QhvSqhoiINbhK/VRWkc6psN8X4WJSlpv8YFYfBSmSKt53a
Me30E2OJYP7xoy+pyf46iYolq3PExd1fJDyEyyIxxxFOQT3l3CHgY0bHlxco
m7cAscjwRkMpybiLdLNLajdP8To6EsiSnIjHoZ1Nc9NPTT8LeD5wt6zqrSkT
N863xn2VOSvXs2mQNTZsvkCtQbZXsJZH2tPUAVz80r476573KIA8Mka6DrHC
NdGIsFd1P3qvwrIegO0G8rpaRPe2F4BUv2HUfJWBB4XDVSds5e0+Q7HPtlRU
tncEKidBFiAH3X1B0JBzPbVTKwij2ae6AguGvPYDiaYsWFYFfBhnY9XTxHq5
6EYzwf++QK0W2IQrvSku1tIOzZXkSm3ZKa2zL0fiauxtdWO6rTzwMW9bj75g
xMMYUn3Oq4SxowSEdEAYYiCuEsn0TnIlzAISYXsOpmh1mGTnTDY35o/P245z
Wlolb5T1zC1Z81i2mBrQ0f4v9nxVZgznizrwf55Nre/LiIQbn7CdbiN+e0a/
zzLZEXQ9IkO0Ylqp5/r6LpWhl2VLx6H7lTyi4polH0+tksB5XqqliThaw0G9
tuhomISCxGspF8wmEUSmbxq+WRQKwWuAEPhN6A+/QCDIq7A/3mNRAJiKavhX
8zj17lW0Sa9jGxGT+S30GATsIUthq6LeawV7oWeUByMymFrgL3RwU7fEuojP
SuF3bjm9tHJpYbydGz+H7szZY0aFp84pNCgpVVZiesl7CdMuQkn6W4A8GZCf
mMMXfQo0GnXQxM6Wm+VIIb3T2EeMkRc9pPEnWENJLWr1SfT/BwjdXQQZCG+F
vMv62axUZJ2DUbPRK/Alq9ISyW35Amt0Z9s1TTduGYHL+g+B6NOeGL+D1bcR
+DFD4OvNSr/8NOo6mmenUoU1FVglcO1kwxzcbM5/xTdwu8a8AUxV9xp3nANi
WJi5GjPWsKKMGxeHJTP+YLkx3IWXuGXfzoExtEyCHVgZhhCgPtwmewXr9eck
9TUg+Ec7UAd7PohoCSfP/69zn38Z2SYbniLqcRcEQY3F13Lgh5MM7YjfOwzK
ZLj8xpuDgNyjAv2w/nz4Gt4OwI6XPYt6Vrp37mxvW0LyUmdLxIjqBeFgPti+
2pLIv6QF7isPFyUY6+gi7fv0qSNpJ6PddDhFlXLw4kGf4gbJOOA5acvFaZrp
uyA5G6mq+6m/gkYHVD2aTKwd0jyFDjB+W3WdbO7MD1E0k0/SrSMjdDvqC57z
yqFlt6HBF8vo5QHpUuu4o+bmsS8AWsNsrY0XnL015VRLWIDasYq1pBMRVxpY
QotEB5qoS63ypmYyx0+W+ixHc9clVUFtZC+rBQ257h+YOVWKTNpou/FYElSC
hE7BIcML5W9yblKwKnXC8jciL5rzpr2eVlVfoJm5w1CemCXmAvf1ndQk+EvT
lVNKPOw5+yTY7+NwsBW+RVAXpcvnjM9RDW+Emfkz9gs9TW3+j8sqWAjFLApy
vB+ncuxYdCpgRU0RyPTo+mPTbvsHwu0mRdu6ierQokK6KTtUSTM6vo6UVP08
iEQOmApBKI+irG328sObIu3hkDftsMIEAjlnFZoP+tukw6MhBmvtIMtYiD03
V8ldIFBUnT3JHN+hvVNX4eYewfA/v2udQHhtLJ/IAhP0glVaANpVfLQAVwzm
eF2WRpmKd96MxUG8sTKrFgTo6hjoJjHIC9r93YoQPClB/gsgkJhdxlPxqr24
DDkx0t76OGJcAUS0IQ4ShGtU3hw3SM4BZkdG5UtBNovAQNZ8OMnxRS86aFZT
XsJO0wLhFyfCoPac6W1A2A1y1yBKkASC8h3xSEllOwuCufTbUC9Opf6ocFXP
3iREv93cZbVc3K98upcUGk3O8f3o7LxPla+0Xr+7LnEbAGGyc7wG+DGvHKLy
s7I5vJ8s+3Unt1NW305Y7dXnXskoCAjpwOqVyUlYfd/My2eoyn0E8BlIE1OH
dayZcCyJ+ZL26Or1yb3K5NRZ9spDFNYDDvaVKPAqSFbkaSLVVrLtDOS60tiz
IFke1LlIY7G9EaeNK/rEf81RNqvpzXdqlU1/cJ0uzw5qLnv6OvrdCAmjf1SR
ctNMJmC1gpYZrxI9f4tZ7DlhYVYetvcZ+nvKwTDFnyjUVwF6x+fV5pPNEit7
ZivHL8EhgxlBdi8lTfBF30TAqNfYus38GtaI2t1/hDggSVpoTfPCxYTGuFlC
lAZpDldjwAlHwwibas2PGzF3Ktq1zcLvmS+KhleD1tFjbgiZ6lHwuLHiAZnk
QDq1EYoh+iJuOanWy7i8NH5wcOluqwnPxjLY8I7E6s5UdUxtNWut0ZpHTsUQ
zYlAzacHRP4LDungrzUOcv6K2T4FwbeZoiI4r/JNhJ9nVZ5mpbxPI/fLwZQM
31fu881NyD7d/Q/19RlVYj2YhzZbXYvtEjrM8ImoG3WyRXlYmYENXZrLZC7M
2yBY+kX4derhV1C6sm9anjINawkQypHi4dEjs74VnFsTVRQMHhiQSrUOSmVp
O3RkfBM4leClqfda/j/SX+vbT+dIJT/CA1gkhWZuT8MrR3dN5zbjPO81J/9r
MuwcX8Y9wE0MxhbDF1u/Jal3D/dEwNCsYbES9KpNzhagojBEV1CuybrYgHgs
4FWYjQ0F5BHZg8zFBQ6H0iS+5Tdf7DVygh+NT7UGl8DgBZ4El7WRGZ+Gv13A
y+qKCjG7RrO8/il/91gNSbi+HqXMqqpwb5cfDJ+o0/cprP9bOhsz0BjJ3966
UAINGsljXYJ8Jx0sN3a1gUAeNybgYA2n6JP2Y0M29TispOCRIwad489icP/m
zTU63JaOXpskS6Y+3lqN0nj9MWjYJNIi3rJA6LVSHE06zUu8CcDqFBzIiVIL
Qepau4qvo6AJsIx/3+WTylnYxLU+wVNgAiNlVbgeopVi3oyieUyLmuMwF11n
ctLsfxDGtCq6c4HrN1PKiiX2GHrijhmQdLqpXu7bhPHx/MslteawpVlrxtZQ
CJfpRDwaE5wXypeJ1Fs8nvgCekQC2qchVw6w8FbCaLjaenzS6UKDnZVm0bYk
4ntc/DGYMTvblltHA/ihBOyM5EtrAsF05026kiYUtypU2HDSeafs9sKpWBm9
6kHEO0ArrwHjcNWf2KFN9wHGe0ZYOqcr8uI50Ywj1qjQl360rJZHH/GuZuVj
nJY/FD1RzQ9SMId7FaJUnVTWT9x6lOTWRqzGd69MgPrxwWFwyim1RArFMY9M
iaGGJNE8rt9AtGvAgOznVtktQU59wbGXpP1HLAmPH2PPdRBt/rMt/KSbhlEP
UTyC6F1i1NJwJ8W3LX18rCIA45UiFgeFS1tNrAhSagT2GxgLWFAaKsCJfu7L
UURxRs8zx92qbDIRgAeYqPrSDD96B2WAmKm5AfE3nOmRUG4bc7hQyokW9kRy
Rk89d5JNnwxpGQtPktEbr+/ZWD0AqBT/4ncaaceGYcsfIEef+ZctFh2uCL8L
p2s7VQqsO47LGy0ATDMdGDQ6lvs/UzE+1bIu0jnkLOLkmxj3s1OZuQ4uGS1i
xkj6/yhJSt5/6sSCzKqdRt1OOiD61mE3fOHOGIbr7gjaLNLHGUimkakBAi9s
yRG6io4qebq30Jkl7yiOiN4qVvUK65/IQYOk2t1GSHt3cmXU+0+K2JHwifKg
K/vDFTizAtCmnOFt2QxcetaYWMjQ8DABArlg/T/wkAhleARSiW0flpA0ypxd
2MtJeZmi3bXVFh9uUkam6r31c8OQaR6BzsjhOYDl63xmiSpb7KwPspGFAJ+w
lwQd5lXaE1j24TVlTdMzNEtxG9w2I94qS+8JS7RE3PMGwidcetyaCN5eXJiR
hxoECaM6yF19/WLULyyWs8CpphDcffbOEDlSqJeywFt4ECkg0Tv61RPu2msY
j06mPc3xEmppt+sboY49TazeRibUzO26zc3Na1VPpgDJ3TqPkbwqI7PhzdnF
OQ8PK/H3jBSLKJ8XrG703cJ83PwPqbx75BdqDsAbfP9g8FFsuuNp5Fi+Isqt
gcwoKPTtKz6K37eiVugO6MZOAmBmXe+1/3PAKKOcx7lEa4eCnqvXiGRZLj2X
wQs4zwxxEtrvqbcNws1ZH0YSWvtCMhIEguTFjQPCsc5Kt5MUfDL1Rr1iXvqU
a5p96LgVxbtDZBaqpcx13nkP8qTxZpXXcLCxxoK7AiqIsV2asUbDKFLS6c98
wdfj0yZqksTfX/rmcBLHfMF5GCJJnqvssqWhr9Irgy3Of5zXsBhU8NxhAVx7
v3TtRIfZYmqkKs3iic/xpaigsqRktKWxWUXoo2IlBZkDFHXD29vFyAkX1xxC
uajQkw8QISJYi51kivrLK+2Hb/6xm//T8Hs+D/vkuhJrmZXOcJFInxPs6+5O
QDOHu+KyYz6TiIBmwdvnmBZIf76VD3Ue6ysngAM+e+hu7eAxZqIRv9+ap/fO
z0F2mX62ybILL1IYK4ywM44X5w7KexLKY0YUQLWYcim9LTnlgMbOXtlsNb2c
ZQ8cwAJDpxL3UNmaaJ/jrG1WWAyfumun9AQDMORYn3wE/D2NHwBc0mP9JqIc
ZxTJkNk0EElOyB73mXrm5rceSmJhmwc1wq0kA65CY86cYgfSRLADBYoZzvrd
shb931ExUSM2gJJPlxDyzSlYne08KWb5/FrnKqo97zBl5fC/UCZdtOYmuFNQ
u9S1HNQCn3AMltmLYeLF1KoXQcHoBvQ8sRZxuHnLlmn/FBNC+ZPdTWvWApiZ
w/VIU/UMMTOTKMkJb1+d8OpQ8dpNylsZalK4NDRDyl3jyA1L2WwbuwEuyMCI
OfSMPu0Y0jsNVU5Bvamx2jvMtUXz1crNlXxaSbKeXNDyfTtp6OTXRtMQk5p0
02sEjKAnQXoSQZUITSvec3b9Uzzy6qYfrd4vAnngDGr83maUioGGwLPBaVJk
DpNr+5jeGSv96XBHew1oh/4YB7CYpLsTb5Tm+m2W5ZDrji7hOqpF8x1NFPVf
mDan0qmJo9BqBf5VyriOgugCkH5gWoDaLeyuKqwyQJ8fz9J+LlJIt4oZOFHW
IpkK6lwizhkvirkIZNBpTBw9v5oZqtgdw11nnqJqzxk9NuSJu+ecfgohmf3y
Hjhal4WR2YXpsORG9Csa36LSgAOHLDgF6g4Ryp5EFbUsrIyur2428b2VjYOt
zekCGzOW7jNViggytxzoZQyP3K/HIgusjOpQU53sm93wwjE7xjqYyvU0lKQG
scvy/Tt8IgVxod4nyg7a/WKNZJ4PFAUPyHdC0H9uwSE9/FvR7PPtPu+CRofw
fQ1Ac/2F7bddlh/pw3CpiT0MGIIkn3pTO8A8cZGa0G2+qju8RkXwN2dZohbw
G74lWESDlO7HcXESwUm5CE6dMdTSBxiHWxJoHM24pA2w44qVyoRLrN/7we0B
OgbJQa5VvuXFEsrwkwMNLDh4X4T5orrOZ2k7gHkjzySLkEkPsOwL9r5wpYus
XWKIDu14dZryUlfxv250XvLvORI9xy/gPfgkDH7SJG/x493y+KRihjvQUqtt
sZhnlUrn/2tvtAVknmENVwJ5nuzPZUKEushDtEeyokph2u+4q837pRLoIjeE
WK/4Vbam2uuNhGxFratJx+M2ZspmIJ3rBxu12+cXMyrCeeNzPksxaoy5vz+s
gVnhxINfBuitG2baDwIpNqBvLksX2Cte6YBX+8Y8fyIfgannxd4Vidt5U/z5
tw1MOZZch5SUptxO2EXzdGVEaJqcoAD2eo9gKYaqb5t8gjpFggBwDl04+E/B
HZk13njW8bPeahngcXzg4bOtzazPbMidpaOMUcm6iSBQzRAFT2j/7PNS0PP6
ndR5fpWvSb1qg6S4d3esSXdM0sBeL8nIBskswAWGf7oY9oQi0BQU5/SHLWkC
Wn0kuFp1OrceI4k5BbWUuvs3v9USa2AXXA6al9wvxo3FBwa5m6EGUbFZezYY
M+4EHqZRyZTrrlTT8wzPWKzB7G5rTOgGlxuEKqMDwXAxZNxZ97UqEZfSYdNA
qGoF0xIsb4BEy4wM8PAINuXPir3+05iIz1GBl66+kqmyX+ZbjhvowK55+Zp2
uVB9ws/M9yZVQX4aTd6ejX6rq0im0nv+gsqbi21zr3NiISY5x7SiqWQQ/xcw
uWdbZRAWTwlVnXOoaFrZgT1BVAWj9Ora1vQ7soSz/fs5a4LyWlUybR4bKMGh
6/AJS4Dbrap5Hxu6to8M8CZd0AVin0gVR7ydNp+hlLz7uJWnERPyWWq+LiOl
IeFB5TIJj2thykmOi2b46HHgMf3Q1+/vn7L9BSDGd7/KMBq/seHt8ub5WH/Z
jKwBZD+W33mtW0VdoO5dI+/j1jJxTTNiX8d6iMG48Iuq+MhfjBzKJWrWwxc0
/FEMcW+67TCT56WGXl0mwZ5vZmjMUPF0FrWcEN/YgtbGbsUEqPVMDc4irUGd
GzpQXE4WokJ+O2EpMhrw2VwYqdtavMPIZLMz4JxtGLn+gERKOihIFp006ith
advridC+dTMtt0fPdkwQbASmyS3OJKqx7ia/YVFMefigzQYzoNFezClEMuak
mxJP5KP3R+NHX5ZYMzpA4L2aMIPyg1/A5+HdYO5GtTK95yMKkWVuK/Jg/VxX
M5VCNyFpMqzzQYRJYHtxmDNjtqoBSYq1kg2Ic32bnytkr4pZbJ4FuFFo1U1E
dClYY4qywsO5DnBu5LPr4s54tCaU2ozPd3p66D6WMGVIsjAvSZObmcK4k/4Z
73MVI9MPrVn956ys/RO4QtSl3vD7X9W+UpZx4C+1Mfg/pxkTEWNgze9cxlG+
Icu8ss15565VMuM05JyCLZjlLkYa/+92J8k8j1YK/7cLpgTlRv4INnHvf8GH
VKzuv0bjzwqH9N27Xwxy1qgS5UDjjagkIyhQ7eksB25rihQA4f42/UGFFPXw
kViEuqGeznzCIHQpPcW10b02PWQghIWye4G4F/x9dhd0IT6eqE/jHxOQCL5x
01xoHYDDkmjqBjQNsPO2085NolOiwRcCcyAvOGwbnx94EoJkdW2Pw01P1sfY
obiy3PK3JYfx14owC1I3JYmaSY5IOsLZA4Vjo2fl1tOLOR/GRNbOHWeOnI+b
UtS+oVRKbCUzrj5AZ9tNDWPh4izgSbomctVDhN3sIXNlPzhArSFWkAUuG4Sv
kLII7t/9arf4ACQOQKY87GzTSbk2SdnhJgLCGjoGep4g0HsudWFbVzTjO2Vt
H7mXowW6iNVzBBa5v0Te1Pu3/HZOh2QR1lwksNcimCGLw+i0Q9p966vc7/Hr
zcsl0G+ZVKKv2pCVXidNnpigz/NnhyapZ8HR/08cfZq/I8g1YIxSrDyMKpuc
kjV32pA1OFU6ACQRk8GESLfpVybUDCtQo85X5dlLs8DMVzYx2uZrkEyCE1Y3
tfcsj5oFmOiWJOYE3/yF25uNVXKZv58ldW0XgQzjiaQ3PRUcnZOugk5zWeaQ
798k3amljRNhtgHoktd9PpxMmXpSn6/RI3lTHx77fSoTg8WC1cd85Nn0Vlr8
dJ6degamXTpcXWjQOzstB5no4OXQskt+eCS00U1Bx5Hqch3VwzT/rXGw0YUK
zMqbpCAGIeAPEv52BxRitpR9/pjRlfKk6tgiDgEawJsEXprBXjVk3V2GHZUl
z5JEazX80VLjqoyx+zc8Prr9IxhmjbwnDVG3lAkv2avHpHXyu2XomVfHx5zn
CbiqbjUyCJDT2xT5zKenVa3SvmdSzPCa1vSwmLc16kKMdxQxOUOR7K5S+HEM
3JO/zxCphlEf2CyKVJr+PVMGMpC4SG31P+R30DWWq6esKeJZI0N1I5njRKQ1
9zOrClJTmWJnysU1oUJuLJJSUSEt0ruj64DOyrKGu6FpzTuiO60sevF5G+Zq
zM3c1JfvWsoSjd1m+iISAThfuMrM37UCiFA7I2bsRli0fAPcFDNMgxGsXLAw
FCALI1wtnivn56Aq6C9Nfgw5NZjd+UvutLRk6u8grsvuaJmHeVMIxB6Ija5e
cY37LNoApENTw21i3PTfioV+ZiV85WqwKoh52xDXP7yp3DUDySza8ylTROzV
1rBvNFPnyoB/QnRto2DQXRqljCbT5OmuFovr3aDDUq7qwfvcB4jYPkgMbgy8
G1yQ6qlFAf4bJv/vmg0YSCpHWIDEIpcXUqd54sg59d+Uz1rgV/EvEI2oHIgZ
TbAM/4ZN0CwXS8ZGZJur7YhzyJ487oox5nyEV8uLs94qDaLTTobnRq3hellm
RfF414W0KQxzkBZjknRYkZuwA8IKLUiua4uxg8fiqSEuQesqUTnamkHsZ1fp
1If29ztexVL76OxmzDhIUa4jPeMncK4POPqiDKrNpujWYrxvaM5kk3HiIBuZ
A2OM1hJe9qLwOgoKbIBZfiUa0OPFNQqpapX/EQZDUBVhn70QxO6xlz3itIY/
kifA7zHBl1J2giOm8i0CScpU1fFsgaKDGtWOZBDk8FaCG3JEz6kH4jg+gj/I
BqDGd/qENBGJooQp63dCZRuLzjUMhYanTq24ZEp/mqH9RRewGhK8HjMCkH9f
nnBxaLjo7ZmU+QJvJYH83fP0wuDHNQGROCj//qiLU2bc42sWeIHofPFVSp3P
YsbnENp8VvDi2j0rC6B8XaAiUeUdJfhr4x2fk/sCbANdrciAxq5TxE5k9AjS
nrJjQ816mlLdJlKeTAhdT5+IROe5vurYM8OlHvtAXzE4+dtjW654FkF2NC6r
fqm6DLAlYGso5V5IFFtrj9J1vL8cWIfdwx2QciCA1ecgnBejXdKoLyaO2STd
rIym6mPZazr+aRLWrgHgP18Lu7H2fnUYdvV0l4zM93OHl+d0+4fTbO/6m/Yg
td7o1s7B+H3vedeSO2YuCApxWTWOUPQ2IejXUkLndGOq3Zz8aebcVYnz4kIj
3moNA5qZIlotxWAlNhL5gNmX5PwU0kSK0dr3gYfBX0NFrXDUDkqQyW77arxW
h9SAAy3eMU2OZWdPyGBtFI2pxjezA3MsxPh04Eb2FKUiLf5SKIWFqrqjpdy2
6ZI583y0H23V/xxhM8DNW82SCrMlnjks7qNd2O0sLcX8fCnstk8iS8+orWj2
pNbKdtRfH5VYWnXbIJvN+jKDnBfS8pVcAKKDqGWa9i9By9G0BaicrabHLduc
Wz4CuS7RYaxRSesjj/xPVcyoG+dNPzU5f1MI/ouczWCWKfG2x2eaR2KSynA2
emRD1bXA6BT1p2DytHmfUeype8rxhoEHvmYH5R+m4PLbKT5NlDDXOI9ju7Ln
beGtd3S8w7jxYW4g648xAinSiNPWWarhJOYcsZgjt6BHuMq7HGaJzZarvXT4
5/QnvBOP5lMr+XMGVDzujp07ikmvnFtNtbqoRkgu51apQqwISOdRbPpHdqAY
w4L0eG0aiPlGrDxYwHuZvDeKGxmFOEcmzlNSjh6nMkTU4N3aQUsF+CBjUZC6
8jmsclU6GzjqZfAt07yQcQTKgfPRnQphMkcc4+zB7EgHOfN4bbkBjEDjH2Bt
WpczozH88+H0yGnWBaX0IuK/q1NlRaNTjulAaSc0siQ4DnHJPbdjYg8wCrX/
/KFcFJJIvv9YJQbaoV5vaxwxosElnZFSIrRS5I+o+O72PmHjW/VhmY9NacVG
FpyHXE/5EdgBKhbt5QBY4NxVUAtRejNrOghlhxq2XPMAkI4R8DC6RZqre5OE
dK90+ZBj/HnBbu0zV23X82kc9rTam3U+oHpe3gKhF+jPd+I7U19whBKlK1c9
8vP92MCjpX++ZDuu2kPojubcdy+REYkOc15UDsZOvDwGnkNloa1fM0O8Ow0U
W1EyX7xm5Ta4ODjFh9AGFlzC5XxxvD/MzAMxr0jVzn93kGYkggQ+Dqt7XI/C
ajKVLVge7ffXKy/dvft2VV5BqTVMh7yw/2bRDAZ61tn7e1ix+ONqT9I9lGNK
FkCLK8e8Clipl29rmLE7M+WsYiBeXQuMSOwlVGa8CSpFh4rbsEmfsfp9FBQI
j1mabsJBM9bpg5rUSPqOHEPe0MxtBk42/URFNVWTewQ5vxbT3uWtVrDNtkdY
RwbS9oExFUbDlp13jztF8Rjx084FZj2CmABIt7ShHqRTT6YWHcy5NF8QiQ+2
XBdTf80vGgmhvVP1rBoMVz/gH7YjHPzXxhH3IwOEewgtHkwPNICF/qnrs2wc
Lc0ULHlkKLUQiH5zTBU1DmTZZVYfaEu9DhhDbha/KX71O62tLSP2+lxoUCFj
X2tqiIbGTY49lTaiEJmNs9VvMskB1sLv5v+/O0Y+Lx58/AGf5A57JvrNqVjE
MIfRKZaPYH4ef+EUKvZz1sgEgLjbm41JVQ2MRQ7DVoLBzwD86gaHucPFu4qD
CIme6UQtFpudEflbEMRtv2RrLGKzPGL3BoShaHam2jQgK6PQuWKEfT8hEoia
bHLoUFRt4qjSlGF0IGepYfHBoAUBbuFY5TH2NRvzEu1dii5nDy7FGLrkGOwD
L3wTwHWbUXL263Ot09hqcC10sZjm6Ry5UGHoXktzxE8I0ue4vY6mf6NZ0LbY
F5qtLqduNaVKd+2DgyTAtQmO2aeHn1c69xH6+phNNTaKOtg+XnfW3MQQ0CTL
M6KzDVTJOeqtDm0os1oMxdfcA9vZQDv3HtSe+LLcTils0EL1WTcNiN09onZM
gqP7ZWFHo90sskA9aDywphOlW52+zZ5Wqh7c9JMu0XAg/TtIqY6RS6ziWRgc
4o935beeOqptXWj9oEaXO45omOp6rrBuN9pIA0q3poTXRHUaOfHbpd949yzH
RZvjbVKU8ygGLoIv9BjEpiEAbr1GEJWBCikY2VNXJzJ1BMcd/jPHaPkiBYGo
BmAeE3GU9NKI8drVgSCwyqsq50hoaqre1uh/ZTagKmtl59Pfuvguo2HSo6cN
gOgjZ+O+BTE3rDx1VGqD6foRzti4MtSfvWHBbWHPW/3ZojX1R2dPDJRB91+x
GiUbjU4bxq6F3pg+3k9WJDNH4AlG9bnr6NrGO2rocr8ypkT0IUpnsngh3KFV
ZtLkKby/tSXdHmFVYNB0DS5tQDvxVKgaksl56gHNdlG3fTam0HJzDsz61M+y
bFfa2YHIq5oTotd5ziRahNq0KcOYEJBWwAlqJnu1BpPWhCzG/8Lec7wkT9u4
fPnuc+PC3RGMZeDvOLFKn7uRtwjukAXN/PxQdJeM4pZfomzcA4YDxGT53d3Y
WkckZq664sWXZulsISeY2ApoVVIab9BykI5Ix4y1QK3Sc9iAKHkhhWadwbnt
iXLuUAfF3ZGP5pafKLunL1+8rPZGtRHYEFfofKC9k4WWcMfj4RkL2oM7F/pM
OqH6ULrZuWAu9gYx2XttjjzPYBGhHMV7HmkjDs+tKBEfKdpzemcyKgFimzch
5S4rjgDUy979ArIfHlmb6Nnh8T3df3rp2g0b12AoYyiFtDd5x2ZrQ8J2VCeM
h3VSRq+EjcUMHyCw4i3R9I+uEaw0IYV8WMS/LHlhzBlf1qW//dULVcIUBGWl
Rh31T85aEOqgh92OyERWey8EPOB5ueTomh8uEurbx8NS+7iT2hpxxBVH2nsb
9BkFSrpsdyiGGSl7yZgehYWAzAISsk33XLI5WjqR9FmE/8Ud/jZyke4+q8a9
n9kaFKqPOKOO8mtcJ59XAryLMF5MFfUBD1VgF+TbCf57snPx2pMYQrrd4QwX
puny2yFyh5zs3cGUZVC2q1sImsaCAlYCVYYMF6VP6NKN7SlTRRT4GLu1iwcM
vTiz7QGpIRI6DMQmVqLmoGv41jdXJJKCEJRTaG3iOvhu1fuBZuaTW2J9A3bx
Bzhi/TG6fkM90JnNC0D7lR5+Fi4sVxvOa8Em9IHBdwi+OeGaLzwOXYUMl8Qw
1MzLZvPgvL6cUhROQxAArdItiz7rJc0H+BoTyh3ONMhuNdzWQRI6HqC9hkCs
AZZo8q0SCOlbzBc+2ANuRGAhnEuAsMTTIAkXcQqftHJiwqpiTIM5DB6tMSSc
i1XO7Yo+CSVCDORD0TWz7ABTZ6JJby3zDgf2PC9R1HkliVT3ITTMMrvnpQg5
zIixItcg2gny2FK5XuTDIH7e8JIhx07ciF5XU2cKxnF9+Ue82OP39EgnFOTM
PiIaxfuGSE2aWoX+Z7JJhF62zaM+yEGEVfRIE6k2UZI7kE3wf/QknrZYO2Mv
nie3sWimm0nX7ppaQ5W/vK51gTNHoUUL3MxpaywTO37yvvm0A6c1gOo8yP3R
MiT7Bntg9I3lOsAy/bGQn9WRo38S36jJIZEivtibhWx9aozmESXwVw/q/mDc
exPmRS90EzphIhqdLaBIYezXx9VvJW0N8O4gPXOaBNINVXA2d0vEHw/73B7j
9mnDiPSkrOsa5ZMGcXWjinmoTNfRz8rZE9VyswZKEnlh1xsWPGd0JTpicmkG
NJFSxFPRGJtdFle0qwYtGUZCA8l+HrT7zEv3h1D/jI7D3Mvs42FIYc8cFwwO
vrHiGg77cMMhP2/BghJOLGAvdY09VdXpv8ZbOiQXZWmvnxxkZXHkcAbpxr6H
Ptz/Wx9lo8INLHu2UbC45PcXJ4O3Jrcpqiega1gn14k6/VBiPH4heIxW51zT
wcr8T1NL7vxwKv7bQTpi2kw5wYM6OPNGwo3jvFjP8h3700ZVsKAWND5b2BC5
jCf1VqI23U+rwTSLSgdYcjK1YkLvvrZPFNYJXawUSr77/RPTjO+QCZPwXJR/
76vNL0rFs5CWYnQEPQwoEI91XBupxRCci+P72fJzbEmXmWEAsiCHGLJLlKfx
9ijkD6I4oclIZgkBOK/Ty/ZjqOYSEOkJU7Y+O0UMgG553yTqBrXqTnXe/gL6
ZDL5nxDmGsrbxEggWAoelK30hcV6GZT4ED2FgLHDJHxntb7jun2Gq/A1ZfM4
QyEf0mHeSTZcsQBTjatEo6A8lwQ0HlBdLT9u9INkvIj9bsexHa2eA0i82/bg
XlEY/jL3EmXNbnWM13UwSE6wt71Km7fl4CzYDlQrdn3tVd6wMpOVjHjW2b7r
drgACpjjFLVjuJtlLMXAdSMGK8BfeXHOSaNL+zt6Qyqt+TsWKCkCRU7PmO6q
DpbGlU45eiYgXuu3uMbYotPni7TfiiqZ/oWDmrTyRLGI+bgoizoYtgyf+Kyr
Dqgh1XGnwvwjp4gXlLDEI9aDCg5/XK70N7RR9qvXrkoFcI8FInfK8i7jRMhC
VVvVUgamKgcKzyEgV59lKAHFdPSXpv3pyCBry20CYCkm2e0rIaRdvTuI624A
SVd7d8YbomeyqhdEBcUgfFmNTUiaOoaP6Uztrw67ivw6Mv9yHdTy9J3KuTt4
dicK90pVV5TVMKd1ioX5QBerieh8mwefmBQgcmX24S4OLitdMmeHnAYI97VN
Jy3d749k4wpjddJHlwg0kNhz0e4wUjcpAdHbDUnEPmyH7ITCHhphSxfCg19q
qiliKYXaJAkwaDcdoimArzyQl9N49DmgTjqiaB5WLJT+0hg1fXklToocDxJV
/5ssyiVsCbx/KDVtDxdo4BJ5LHAOjMI3EyvZigGRImXxhiQag6k/U+m2stRI
7raTFHSGA6bgjpyRCBqF7nc0d8oPSxGMh+81fvxycjvhZkaiQvX0YA05X/VZ
F3l/e8vifGZbs3Vsv7IhgCsSdXziuCClypfj9d0Czq73UE9DmNZMHgnProyQ
/5cIhLbe2Xa1s0sZy94FlS3bNT2Vv/86e69guF5d3MAdtNfaxsUenaHkyQ52
7Yvos1QN3vjIL3E6W8ewCA/O8l3K4RYXRwJiyf5rwXjJn/9A3/x5v3RfpBNc
fBJweiqpjU0t2tE53aqUMhZYC31KVUe5MlJSBvcgzKGmlvdnldR/8RNUf6Jg
/e8D5g3Tsfia8weyvacoxKyghevdaL5JIAGmURNm2de+u0wPIUemXCAjABZO
30nBNwxpnOFW6frG/hnvG5z4BMAfE2FYUM62Fha9X554mDwHHSX7TNvR73HJ
L/iJrDBhtIz969IyRI4EvUBnBg0R5K6xyvcOhHPaMdY39/o/9AEAnNDE7De/
4c+kuzfAwMdnT7Otwc4M9gOnchazQ6TBSa9l5kwX9v1IdP5JRTfRhRxG30OI
LNQNwdzgm743Yu3kgn/shOWcDRMFdMwmZX0P1RBJBvES5z+qQrw4Wl7Uo6Ei
VNlWNQRT7oYvUupgEG+O1JZw7k96lq1Vy3XfrIpgfVF/xjLKziwx3f+lG4A5
8oRkZCWuH17Jybtqf8fOkvUS6bQGeLug81x/tNa1mJv7dIN2Oegr9QarhOg0
sC4OU4TDcddQ+W58JFAc/Jd19I/B/ean2uVp/MD35I2LlWh3Q9/fmrTeS3TE
NHTncw843pz0GelfqIm1NNjXSr1AHWLb92MH+rTAgLOf+4qhzmPD0wJfa/Cw
6dL/DHBwzEIw7cxf5+Bcf82RBW9v/apY3exeBh3kWLucHsifW7mKecI63LYO
em+aG4AjeZnqvCCLeRokCUHXikDfm7sbnU46uhb0mcGBcviPoXaHznLoevnU
lzftmnj8C9qk4JKr5ptm+M2I+oRzT/Ko/LkN7859s2RCN86Njp0DMQgrWifA
FutMyMfcHohV+DiTUv5rBBEqDfnstso59xihY0Fe9qkweUgRijpoEqCyhVf+
48UnBP49JXRU6OoBHwRgIuOcOZFpxjaCvqBqVoc+sH57lFL3E6aGGWShA4ij
iieBZJ5gdeIJA7VqZGbF+dhthfnref9xv1mKeqPXvjyaTGiH1tCzEr5TpQIn
7h8nloL7oVPIj1NVDA8Zwy3f0ZDq8IZ28WvG1M2//AkuWn4z/GRUn5iipSwB
uEBLx5YDjDLSxlWIuN9n/M4HexscO0PDho6AQ2K6uirYKJ0107wh93yC4mat
nabH0+B0w07mDAi3FUxyOXITU5hh5gDHQYLToEFrtjoimjCt6RCB5QgUsw79
H5ley9QZnZvQfoRnVJj0blsALrwEKJA0MryS/Ep4z3PoOpVNkgqxFMra6W7b
XYo22CEyUBj8DSuc1qACk4mczpSX020U8c3utrY9Q7SyU61QuI4VnATjtI2r
yFdXZaDJTYzoI+obAfZsv4YhT2AchPtqUWFnJW2/loMwQYX+wbkASvXXA0bV
/+kK3bSQwRsFz5W8ScAPCyxKAhYCt8F+gaC15+PxcZ9v/2Us2kHqjKlH/ZBL
+aZAoCDHj/bM/93HhZouXSHUw2hSd2EgEPfcr8ZPHaToDYmrCYYikeRBifAK
8Q73jqzPmIYPuoZjfUEHZ1/UqP/EhUXyXKABO7qYXlg1j142DisJrlPV7utc
8FpOQHTcau7r463xZILBFOQ1o0/nLY8D01KqtaKxZTCTgLv22/r3RJQaChrh
IsSn+9+K/ZvWC8FgVnZ2q7JsDXzdIwsfs5euNmyWBAUnyRCPggD/vuPJSgB3
MEn9p919PVHmw+wyWnCXPuLOVVgGG2v6q9qqMdLxZ5DH4TH4Fsq7JZrzmhjz
qfY+8PhZODR03gU3R2oHirHfPY8KQ7kXY32xOb8xXvmaKfhbAFRWw4AXJvSk
OueWHvGnHOCKGdM5cPuPIlX/BeqCUnKAElP0gwkiZplZybHccxPpnPNeIcB3
fxrICpt4i+PezH7Nlmvlhapw4JGOxBEKXIAOTYpYxpwFnQkU/vHaoXX/s1e2
DVqXEjCHyPSljGI+QtTgQ/DnaK/QpbFguBtDoyrsBOFigOrl7ohKpgigpnRp
4PLcNraRLuwYUasM39Q+Ft6xHzMtHEwKCh5h7f1pl4YdjWmQEqwOYNlmKTFS
bklywagbvX9jYrxTXkD/Bloq4uHQoQhkYZsMQtx3+Pmv3fGtk0qzCQujK9g2
tlXwqU3WGig42WgKC0IaPMmIoiTHU3lkVWgxQgH2L36VJ3UDq9jIjStuhUpm
l3LjdNfZxBIpUOusYcB17gtrVoB/XS91J2r9+EKjmgWgeLdxDUwUpebt6ydD
6/EdsGJV/few6mNX/b2fTskeCwi/2BChFFfKlqX6DNP0gUWw5AVWIUxp9NMi
qFiZgDKSvI0D28j7vRGzQAvKFiOMbIYgXOMZBZ8QxG3+ZL7ZYZKOPLzfhhmY
gJV/rGBTc/JHi3AnX9N3CyOt02+VDoiu3P64Y125w7XmLh76qrmuWwM1atHx
UDqSvgBVcBZOPlf0CPnBaU5NPoIO32u0a1SvPMdiBlqAisuLAi2zwVylQeLo
TenmJKV/XIBAphYKhNnHRTzf7FhkxCZbKg8lAMSZgWMK4vigMqWL4KmwLAPJ
/RvLAhtx2UjXZI82QxCdraRphEQ/WLxseotqoTv2kPvUCfrljLypWh/b0gff
fdj9LftkehSamArUGMJ+mp3ZEV6kdoge8QgYuWD8d/VsXh7BURsjDwC22405
l7yJvnQQMSZrjgRliwgHjOd/sdqga99GOsH7UKAym9CaEcgUpf9D/JeVpLo0
UD84m0q667EJSHuXK6p7QBpX0BeMcd5ebsLL4G32VUC1328JUAzCTQnLqqrR
ddsgo6DPnR/q/ejhJeHteylt3Cqd+SvCUxq1snKf9i8yncbXQ8EgEzt+gJEc
ex4wca8TqqiPsDlpuxie+XyAgGERyGrfWc5uuB593p12v5Vu1jJYHeRyZzGX
Q8Ubm82zcI2JH7ZCVcmcmb/cAEsw+pVGVC1+44BBwZo4kJiYkVdZTRycc0pf
QcXwwY2Fz48jIBGzYEwfUq1+F3Q8hw+SUxVWGAI+kuyASRouxKanp8sFR2Ze
Qzm4Enkd+b7AwV8LEwb+tuqcECfzPFLco6u1e/4yNMiO2+lyUgpwU8Kro/fd
0TfLFrVRah/KK34JfxbsM2Uthnu6tl6yfKDewX/WXqA8MaukFp+Dd/z8h788
i9H4C4ddBNobfTyJ+XQK3FLauHo6I4FTAlL3ayLYOBGdtZHX30UzdQKUZWPF
JdTlJhscqyiuVEfv2nNg3nZbGWJXoda9+tf4Vum6xnsAz8GWftLRF+mplNnc
rSrnuy6dT53JIzE1IXsz7i8K8s75RssP55kB7T69FTpfPH9fIhZ6en/Xi5Eq
erketq+EsFCMiNotiQb5FWTGr4jayU4cIbuzt4M3Oj4r3qDKh5GhnqXWsHOi
8hGo5mfrMDPN4YjoSTLv1jyWJ2zf1uA5bgpvpD4pnFpiYClwnGEnHabr35kr
7w2//ngDHXcknDJs37+ftdLHVWzJe4hxJxNi2/RDAsKep2+4+lGARy5o/Te1
bAFWfA66P+RA1cIMwyFA6Luq1kOALgmgjKCiBT4ss5HqodOgxJjsQ6eK6AjL
sGTnjG7/s1Q1nW6n9Oe8Al3c7QShd2N/i0xVjESj5r6mFe1T7UEb1WODcBIG
CtMIT3ORmLKM5oGsIFA8H7hsesa8jo1b/B5dXipGEPODvJlXZVBFN/ZwOAHb
ydemGq9tMZV5xI6ubtGdzPBsXAB9vRDmb53B28t0gly1YBBF/tzVNHT4mIoq
5bHFzjNVaoVBAo3LfDWz/c3PIJE64ksnNC1CLfFDOUn5QKle2V7r3XnfbqxN
v6gIDute9655jAQ6/dvDsbV1HZgNvmeChjuczFqCX/1F4NxT6d/Vu2SLVf0K
s1o41qhv4a1+Zkbhhlcv2f2+bLQUAFc1TA0OSHODQT5cbBVvidihgUaVmAxV
1Bb8/xixXtCVSwvN6TjvXrzoilDGIWVdhgEmVpst30m7BhaFHCc5ggF2ehQX
JEMqoLQtf6ckg6RvLRZYWr3xWkCetPp32J7+ms+mox0/EufIUvR+dApnaoTC
1ieIHVzXRMLFxn/690jgzrTxLr6ai6ALGjFihe7a09n6GaygQ0TNzB5TPMxb
Tqqw1Ta7MaFx+CpPuGVX0O2Rr0F7IPbVBnQyi3jAUHEpvEwPd3Uz3jHCwe02
PmYSRHol4VvluyMCGs9tutY+zib9LZB1c6ukqNN289D+GrXW9pzv1INq8gO9
dinsjlcm1YB5ya+kl7OhULz2m+Y6zvfhet5Leq+K127vSEOSGGxW3kReIjrN
/ysmYfwgxhzersK67d5MHt7YAKWnauRXb3fuNPwp5ezS2lyObwvn24kRVmZ8
oJlehzRj4cdR5MfVJS4L6I/Ldi5kF1ZG0EGhHWPpdbvqE+izhN/zywt12e8h
83Pi+0KME4hp53qicnnrji3L1o2VUc8RVSQpkPtXbgECjAFjz/bwrGlqoYrP
4sXutShwPpD1lTBxfnB3qeXukS7YA9uuLzu+9af3NJ9SHfNVmtBgJSPg7E+y
aC2fBlzo65Jh6bVOzkV53+l9VKWPgJdgMCt4qWWnu1ZiFLdwYVzbz4nq3Tjm
42t8JBK6sSRYgC6/kiss3Wmd2h9gS8czh6lBanvljwYr4wP6BuQsW8Ek+J9F
f9y8dFukg1B8Li9s+W8bkAG6SHsVC3CGlp30dY/kmtmXirrh/0CqAZb+S2Wf
g/FlM3GKyaGdIxtxmybJftwq5kH+pWQzBkZdaj5QlHw77cfbLO/OZjHgOI9h
IXWjJ7cvrpQNgiRfffa4YbtVYeqJ5w8kFj2xyzFCq/ATXn6To8cw6nWpiUHH
Fxf4OUw5Y2W6LowqsUapmU5+yv9pOgIse2w3AwUDIMtBuK7vuwdTsF3DYjLR
4KfCd9Rnbuq71R9DZwkLoQwMECW3Ly9/NlAjSHtcwASb9aaoff/+FY6NebAB
y0MRdIs19Fx+5CNjqRjJuiAcOQQsjgU7AKTaTyQUxChKW78txsi5iUPgfAew
sqXwKgGSZO9T7ZS83WkwjxO2TD+3uFNerVmTLVMbo2P0fCcWMQ1un4WAZvli
7tNjLHlsCeXkvsrsv+DOHL85KWh43GlaL3oGOGnETvb/bA8rDP8D2R4WiCMy
yy30v6/S5Om4c7MbIlgGvw25cvmgtwBMxoYQFRmk5Ct8zBL0H2YJLorA8fuO
TLUNnesTYe/7pZebJuaxBcJYZW1x4UQ5WLbaSYgC9MaiJWdkGACfrSMq825B
xGgEew+qkZ/RAn+m5+YQEl2mDF56noCADnzO+4nTvXxRq5O99qKFZ+ac5l/d
9W4WrhM4DocYOn/8Ha3PR2aSKWAXeTp3yw5bNJWdpb/pssXXieowiqNpAsK6
+lg/sjEio9Od/ypa+Ed9I1SP41oBpPGyjtIxY9A7j466vc7fg5kRiCEc5bJx
GMnNDuwI98F8Ed82Sd3yUXE1RXBYF/KYn5iEWMbvkaYYrj6O3TAvUS615oS5
Z9aMyfb4oGrCly7NgcyEdy4HRfXmT2u803RiKyA9UdaAjXngaUVoAUwgjBtE
0+13FwzV+8lQCBx8YNVm0d4c2IvrQfT3U/Y82KSQg5GNcqsbhEIr/w29EjN6
VVdTiMrkuzPnmEPLQOjQ5aVmyk03ZZyXH9Tg5afaArpkXH9inN08jTihO6LR
Oz7rNIEza3rP1kkJ2yTyRZTIBg/fcls2om8vyo6niN4FqoKd0nBUhKgtodZW
I9kigvbHg5amiU/Zf+XInppx73Kj93WzKCRCc8xVT65fJuScgBefUdk3ZBFc
eBPzHGubgq+0TUGBuGD7EraawJqyV8Ng5WWZlUEq6CjdpVI3Yhe/yxX3Ciz/
i8QWD0sn5/QRnxqDQ0mmgnyZus/8XItcF51XCp8XI/WXFhb0Ep26/fwT7qxh
zDz9JvBAHmvq9gTlrpgRX5jW0u+FIJenzqH7VZpqVtKwfNYGi4LCoSSBlgLI
Cpz54rqhfFsSOjFz1ENaXewW6eCqo3Dkz8KEHaojxg4xLUp8hphVvz0Nl7vc
PdZDKziAhtx2techZqM4mOB2uTwMkC5SkUV9Mse4gA8jXkLgvbal6xQeypG6
iEgcKvZEyQaocgOD04elib9gHif8yU6MWxR6wDd4eFXjet18E4xQQp415ca7
JSL5mJw6nuWUOkZJqWecKwF9o+2xjmDCKI0OFUx8hfy7/4sUoH/MpEUZMpx2
tT37wga9MhIo2N0m5fdO80g14tvcQyuImANc6SQC3Jy5JFNdMkMvJd3/sDGb
7QdY86sZr+ox15ecoZ2SWYjWd/mTiDfSVYWJVfDTNAh/wEyE0jqd5NXv7aHt
TRmrY2GddPp3PB+Gai1JYiDW5MF7Ka6ZzVnR53WJivgS1L8hOyjaI+qtENfW
DceN4+PO5EgZsaiCQLyibm29WqUMWzsLYuuHNufQRWLbPOQcUH24luQ3BTUd
fozdbBHOox3J7U9/Afk5WLvCOFGuljntzhnTMuracHYWIufeEfPwEm7hlZia
sZa27UYYLCsmzim1eCkKLggiKngc4JR4aNhBPkD21UgnkzIuK6pWz++mSwly
X2XimZnPyidQx3SVkfU+wzsrGK3NB9hKWWYWVsLMr4Z+KxCLcONxe9cJljTo
ew5NtdemgVvNchFyIhIRmlpw1Touo7Yzxs1mFVbViDRHJm1j1qC9wIUpaqVn
mw7LhxW6LDtvPTx0MRa29DTz1Al1qWXACqQnQpckzxjc+Gb6pdLjMKIjrMk4
CI/fcEZyctIl8GP/RWVx4CMXu413OYeuXxUJz1XyRFNEYQI61RL0Jh03AfpO
tnf0a/M4lirXzN0VtCbpxCnyChDbc0P+VNPfPxP/7rXK1DEVO6s/Jir1Dvi7
tAKE+3SmbfeTYJoz/eRNUIicXNNurxHq+b/fbaAQund93lDydI8jA84YCn7G
m9qWmaMvvICAaBGO11ubP7YIrYzkStGpzSeI769o+vr54cXmyKcWhz6kZj5t
daHNTJACK5V0eX+LN0uVJaQMkWESGFBsYRxQAoDtKNzvOttgg0o1j6QM6+LK
2HshTeMDqCVTJ2NtlUG5ul2XxNTGMCrcOprQBag8msiz0nqJ25mEhiEDZzlF
Wc9f4+q9gCKOEV04ZotJeGas/YzkyurBz3RnFyjGp3YFoWpvtnrQ2iSANci6
R8/luOqLsu07HmTX3jU2sZ9n5ERdE3TGNvH9qYyNM646X6DVF80CIoEJHbpq
9Vx7zuHQx7X4RVxsNmjn5lBem6HXszj5z8edd4RxCQfh3iEXy2O3JmD3dVJf
9EsOCe92mqXiGmvQl0Oug7YBN7eIR43JDUNVsscTWBnVsgtam7G36069vrGi
dURSopbMUV4qcV+M05DR/zhPTY5/obJZZvcQepwTzQJp6NJtiNRrCbM9km/k
NNYI1BMb0gsFGaS+22WKFrkWQGxpxN2G21vh2xKlM0ZQJ5dQ5pfkn5gBys9J
gULCOwVOCVOZiMU+kQod9EtIfYDrkKwtyE307cZqntN4CsC0f9E0C9ZgJgso
l7INeVN6RUEqtrNy0FpCPJKWjQhGT85RU78xT1JyKoCETgHDXuE/1QeS9P9V
43Z0PENgtySzb4mj2q7CHXaMBAMKkUAsJqcrlzpLy8bpL36dBA950LPaNP7r
Qlxou6wQmz0Xts8HCZU7JiiABov4zEjDW14jSbhCkWMkOvqWdWnhHDiipz4s
MhxyFWCQS5SNdSPoIzVoP3wlar5KxwB4hhasSPh/51uoqlr9fSlllxw8Thso
LAQb9HQeBryaqn0sS+shqYEys9SzZckhL3DQJiNWUpSGNaLcwVMh0mpnrOek
J604oEDfgn7cjp4u9Z/W7bgkmMzSNXJHPOBsz5Hv07Skv7uIMY3e7qsJa0rt
f4Itj/5bOG00fWjU/tgUSqWH1SD/Y0ajAjyuAgJcoMWJgCNaHV3pg8gMUtQs
eLz65NKtCnGD2eIT1Xb8Dm8szFmID+MlS2vvLstrYI18FDfMde3lF1U6lTr6
4EKTzvLejgf0WWdp05LGq7qkcc0PT7fZX1kWiwHTEuZFpl+730MK4K6sL5pR
5IOJUKIN9XDnVXDR/1OOq0DJbfJMTeX/CSoHDDBV1MN6UrrAil+UtTe0DhkE
airq+gYoZKftSEo0RRMZ7Y3S6FwvFpYpfl1DkPDUzz6tcHjdp5Z5Nou45oav
Lk5eMOyMb/Hs92WWM1PzcvjlFxT9YCLiPaWq4ZtJIgaHEe0tozKiUdZMGxN1
1aovuzNXjXoktfxU+RquVfl9fjdcITyMdwDo9KO01kJJq+rAI8LSOGF/B8Gy
9rY+UJtIAKgbAqnBIqk1BBRKfbSEMqAwDO15V/W6bU0iCJ1XiaBhHstVahXr
6pDPowLKlA76RCy6o6INdWHAq9ExSF3fQkCdUWzlejRB2wYHSIliJzqWx8g7
JU5/d8QjvUsd7nQ0lUZ/dT+ipLYRZsXmaHd38VS1x/PlAk5jzhmTUmx/GuOm
4PdZAXfuFa061/FZQiIz2/86APebw5rAicAEcCAEtSnbEt5jztRO4LAKf1Yy
ctlQU2V7eSt5YGT/bWqPJlsColzhe/3Pk879U2e+YAJQYAS20oetFf3olPlU
HN1o4NbG6poDGZeNGENNavCTQ92cPFusv7jXmANt2LWwFeDIb7/DFHHe+tGI
L5aFUOPqjQ8qFcdqobsHRRu7xqGF3bzUUwnwTMsunbMA5ykk8E47CIHe7zE1
zLHrghjrZ0Hm/XJyIyUhJsYixiafUpDLO2ttujv6yj1lGvZ+cXnW0nTFvYcP
OSg9C3yhQVe4iq9DQ1nCjvfyQ7k/VvS8xAibrUaGzh+8aCUsqs4ArAfLTXeM
+rDm8KRJfxCJJbPMM6pqzen7pENZL0F4amiuEjdDAldpF5zL2+1vYImXGBFs
54e3iUq4AdaE0kpoME4FQzx7TFxjFPzlb353/h1vD460ZcoYNU6bZQJJJ8Mh
w8gd2pRfSjPfGn+Xta25P5D+4YXRQCqXLXDbVPWNpzEL91rfqm5gL6JtujLs
AxVhjWR2WQQtKHaRQXpHuGfqyMCraWpaxIVdLRK/yneNQFa5/91IgeZF2Beg
Ts/2ugQFge5XynYW/5Pyb9byZWg55jPIM2qi/2u+wOU/80ae63a7D/+SUdem
09TGxyRuekFGnwds9T+gT846nDU0TaBcvFIubvqHhVrh9tf/UbMeXpPaEOvd
QQLcyc4NTaovmp+7tYxwwsvxT5P1kTZ7hhdxSC20NhZT3LKG5MNlq1XBtqz1
ufYXkgBrF1/GaAuAaisCwwXDg5FH3Qq67DuNM+s/YpkIM7/bMWfYR7zNNhml
P01IIcclH+y9A3FyqM6z4QE/33emDnFxNlCD40b0CPEY3ZfULXU0PUTNwiNS
oTFNJqaCchi1k29dA93hn0pPrjaAyyIJYh2MT7J3jn7m/JHveM2vdqUsoJbQ
EAqLg+jzZM8l7XdzCHCZa399AnR3i8uQbCtoWsUTOjFNSPlJIiaroeFIP64W
T2nmn3FirzpuggVsbfmXOeeYGJsBSkqkrtAr0Hr0LDgsDbqtqWhqgWCVsWTL
SGCD8FykelALAJ8L5YLFYue0q0bYHFz6yZ+THNx+gDFXGooiR5qbAzOm0494
INDzb5Yr85nJMxXsPYhaWwNmnojoQyelckVIYgeAXDTjUhbROV8M2d0/96RC
2rTT53BRWlwg0qnf/FSOJhEGiOyScWzsaO0rC1MbNh+kr2oXWnyNjP/gKbcg
ptsY+BL97WiM3VOjphGhs+QMohF8NF8Nl66yPbGKgIfElu7CFiMHWc2H6iS7
hxnnqQVXUGTwQNX/xTAye8AnJMS4ZSlV3uf3CK+Mf/vYZGB8mgxFEjnBS5mH
jYnYUWKhbV80JiXQllLYyEixPmrm3f94HZSghdGdHsfI+v579Izyo0YxUwuH
LjEM7q1FCwTsZoFZzh0IXxazMOFPO1U5M+PCKsdjSZquZWsXzaVRz/cnesH4
YvKFRVbUJk+1yGbPVhQeo2OXiNAUJS5etFPOITjSj8CDylbMaNt3PLaKXqW7
5JsePv1UOyplymh1HQ7JSykFDmTWrxf0Q/PwvazzYsTNGJ4Zh+Lcv0PCKIZg
8g3cRsWr63UyPff4q05ZBsEgvtZvXCkS2qqYCUTazNQbcC7WyNhVtaoqvjbj
ZHrBnslGx6nnkUUGzYNnH4Jw9SuQskHL/RUIUyqOQvekhytxzIOyq5EsJDAO
rK7W4OXfjpgPuBZ02JDIUq+b0fCxJVUvKa+Hta/1AVT0o1Al6LqKyUe671ef
zx6JBf+oWG9sb/dJ8cZl+x7mE20GgT7oq6+r+qSoY0bm0lVzS+5ENNIjPL57
ad2RQkd9Y+PwKFAv7JBnzDM1JQC4MPBPl70We6SuwyGBqQoPi9fMKX5W6V0y
GJvlibgthBWMaeMEKrkptcVggO+Zb21XwPspj3UF6K4FDkWEPpd+qEu4eqwl
hi7z3HKmW1Qyx6TubKZ/JpmD5vAwlHRwczDAXN95wxt11iOBtsge/cMiZ52/
I2qu7YvnergMmp/K2eXj0cY+DApSRo0dyZUP9hKNUGkbIvpqqoj5g+Vs9+pu
vsr+xCn10oc4ayUdHpGZMvBldx1WejK+SEXpZndvPGMOmXzikkKpzFOlnN11
tTEbLwBM5j75B5+Tciu3VgWW9EVEhXdsKP59LRxFZA44iSSszCvPDr7fAlAH
b6SMA/nrBnt0e1k4q5iaUIZRadUnAeC944rdymj8vL4dBH2sKHAeMrq4ORCt
Ynph9TgXWOQDmEk37J+vd7p+jFLPy0MoFohKW3XT4PGpyHdxFryw4Jvo/77k
bljkjKV4iZ2ulVCtXx4JLo0DEtNV3MMCLOdjXAEJhnm2jX+VHeCZC2z39ICX
01MIw0NMM1q9FIrdC6vzvq2ypeE4fJk9jSeVQgo1nRIk9X1nWsfGOCXCcjTx
8QUtKX9aJApQTwFxUIyZlT6P33D3WxlbI5pgyB20wMhZ57x7OY2olVWcFWas
x1g/ovgZCkdva+gTsO1h6VNKoHcwlLbZje3pylMRuoG1qoxmgC0dr/kr5iz3
TZ+6QoUniW7AFLRwmRyfzCX1uVe1eBPOVDAdoWw4OP1arwiwsfZ+NqxFIRHz
T8RRKb05rq6SVwK1Lnsc2oTtzKAfUZYQLMSB4pzIlcukX8EkdeJiyGgB1USa
2DgmUkiLeIfHuKaxw2yXhetXSHxQFBdCgZMd70yBJ1erdUL1T3OLzjccB+9P
8Gb1NGraXsXYy9X2VB8A/gllQAI4uM5F+ueQGocedFUzJByRuN1T6ohmGCS1
fLyoJ2T+FTsW1H4qYJ0/EYbmT5WZdeS3S9brymeSt705nigKdT+t1M6fKMFL
O2uQzJ0mLV1axVGbyNB2+spYXE2OFLgvYKfSN1Nr70DFY8JDTDyPu7dpeXUP
PtB7HwPF1YFJZx2Qm+vMGIkFoYqyn0BX8stOROpXrWXiFq+zBTt8lfbU1D0w
xYi57MFMEMu0Rjzwd5BMdYyKpCPY5NvVlPKmu+0cKLcfQZtjffzSt5RK+C5t
dUNzRh/7D3TlRzEtvoMbtcwzeAyMPMSVSZCEe6xNHE+RLsTd5aTLnceCFtFc
3nmPfuAUqGTtVm7DYtADEQxdZPV/xYFUSFIZQLFyCAJy4wE07pKrHBF7h2pT
1VhwKc6ZAELshM42+9zSU+mJIbQTpVisCm33WXdrhDLOiI8S8nURmCT8HbzM
GpaFy1Lc60vkqf6Xdxi9ZX8HGlB42Zm8NGnUTi88GX+P/WUd7LCFyn0nPwgS
e13+QPREOmvQpY3orDqkFs/eff+6b1o1pfjvonp1OQhn6E3+B/bB9nVU0AWD
14dQkG/MfMETw77WJW9uIFIcAExLmdA5MqVq9Pz1MUfTd4GyKKv9wC2WfD/U
K+xz7Vn4gJRQJRMxOG1dtxMv0aZTMNWF0zjxaXn3T6bzeoYt+JV3Tv983YVr
5HlV32z5TdWsf2JlxPGbTePPsIkpOdu4yq/6gWXSbK5Rss8qL+EPNxSdkp0+
dcTURHLU3O64lrmfv3UBHhH7mkTxNKI2AbcW5TWDwwWyu7r1u++jaJpaluAS
aWeD1c4Yd9tyTtxkE0a4TAFXe/mS2ZmMWpoYkQtUbqqySgFECZG5RdWJ6pLS
519MqWE2URr0pjsdzuZg2cAnieFKBlQeYTEfw18fvOtDzhv9EeQyMSt0RKVB
pEGO5CDqSk9JtpV1m8gT11kp3+/93Nn3ZgI7CLtC8iKb5/zI2FvnQYB4K4Z8
KqHVNTb76ACgCdq9pWeafs7dT8m2g2wrhXSxVdoG1AptheIXChjZ72ySezzL
cAw3VuTwkMJyEcj+aqbjtyaiE+Re94a2cad9SbUh4lxdTJ9BLq1UvqnZ1l0R
0ys1ARBtlk8pcBpeCSxuHIPRT7Dk6zPNcpPyD2XOSJMbl0os5Q2boChrlt5R
kanSUoq34RvPLcWMJCLrF6Vlow/zBWGS9dJxRqxxmpUquE9xpmZ6vf6MApGN
pXYkfvGvFpdKfFRr8hxJU9vEocpynaLpyBDG5/mILliq+KtFUzOpnC2/hNhB
1aZGpv+aywRxoDSL13MCDGKsMDQgYDCft0evUwdTdD6Q/4foxQxW5bUrtdre
t9bskj1A6hU/C4eeVA1eIuErd8Z1iNuXaYN6H7HW/ZVTwFQf4Tg9ShBSvPZV
9fYuuD7M3cnkqdNqB8mkmLsgqXyAFec+PJtBNOKArC7XuJ16Tg+EWkmQYku2
jnPj3vrzmHQX0KI6+h4Dmo2lqH6ugt4NwfzGLqYO/IMEnA3W6WrI1iOEEmBP
9QeiAMkx0EuKliiOFVVYQwKlVn4LwQJJRX+zDgzBE6Rhjfon/LBi35FBuyJy
IYjUpFc5W6CkrbtC71T1DEySgsTOYWhXAbfOU44uCWujLR0HY9qQlsjyZwR8
jng24XuO0sHEsEaSalSYVg84RsVjqw/Wy0tGLdlvYkhnS9k+uuVPZiqpKWTm
XNPEVLWKieTPoQhYkRYPAnYrv8KrW22tjXgvG8f+W0Gq1nkluBv+MA+COu5p
dkbX2Fh/XaUf2zToZhCEg/QhY/9WyZsPeHp1SLSn3K/yqYtWkdxTkgyu7mo/
pf9mdH9a9eDFDqJtWgIlewiezHmQzAXJrGJZC8GbfR60XLb32ITSIZECVKs3
/NAH47Sp1fwmsdx304rccOdS4PCkJMFWdkytN113Uz+JoiIKArdd0+w3aL4n
eND5h8+zUrIWfA816GTkvJBqzs9s4ymSQTqk0TO/uXPlBxLFiPUUQC8rYJxM
UV9EQjV5QEE3cHaPnlfTmkW/BIWuHBe/Q9Zgvh+wP0sHGhzDNAKvkeI5rRSN
tSyyLm67MEeRspSl1+l+QLSFdiH18+NPjiCv4DANnW4W5Z7+j0SbvyhbEYiG
KY9HNVHBrCLx8ozOgruzr2fwY+6c6cNVN9fV0+m5fzcU73imvgDg9BrxDEeU
jFCGvHZ/09+Qy4nvxbEoapYUJ5VMe7Mf5dCG/FvpNsdA83dC5E5CPA5v63nq
dX/tCBNjYI3of6Rd9zg+2I8fD5W30riFQkgLUj0wpl3nV91h8VHY0PmNAfae
Z8p3uEJriOQgedlLQqJ43QFeWBsqW2M3nrZs2d7zm9BytzfGe364RweqrpQA
P+jE3Bi9DJ4lLlOPdGISXhMXg/Z/RxHhAknsGitq5WHRaGDBZsW5twZJgoCS
wt4raqUg0XzDO+LR37ac4WJf4ZYPXe6h8px6E38jNmwMxb9j2gftYxdBo5Rf
Di3q7PKF5s61+hDg+PaeHkXN9QJ0yGtgGsK5LR7DSlRPUosAASeDTfzSCBdW
g4o6lySFg+t8l8lCa/+cXz/ucfNDA3ksOrXvQlxd5zbVQU06wNxbiWgJX09f
+ZoeZMeWWMDgL2hlgsX+7pgWI9TUE1qV7LVBX84zQZZD6oLuFZztEuLMjhiK
k0qdAJ11oyXkYaHzt/TsMH8NR+HwLXGixN1GVsIxGhYBW5SOPdIssiL2zBdG
mPqQNq/cmmL2WiJlp53c+GeZPgNj49pIM1PYlkd5YiwywhNHSpUWCDkCkb0a
tmlLVtO28Mm6cIrDQ3P2ayMedzLwsY8ohHxp6IwOZ9ByVcxMwA+7DOWEWe11
yF7IQPPetsR1WS4xQY5VYVO9Prz4ikhfQc9ZIPcqPftKIMrazLleRgaciME/
YDv046QW39uFTmoRNjwyhe69ahjjJnL3A5f70tFYKhsw122Ht16j09VsOlsd
DvYRXf84ff4aihX2fcIf3z4S14swr/VPRrjiq6WUSXbxS8eG5x8IhyeZBk65
qIhlmw8FXvJchmPwvTHz/kCz0kQSFV3iMpwRx/rmyxGk3BN670s3m7aLmP2O
uu49t7EMfDxlgLVeTyrYDv3ZEShuiCmdm2rBNHSSdAwlJtXMWhBjglpRL6tM
lWr8hbWTb8h993S3mt193sQnB0l9FksAvmDxCaVLQGOIHxRCv+246S+SnO2z
ZehQ6LRLv+o64dyyYNGlr33GLfbTzxZOZ8MqfBP8APXdXrFQJGbz4FfhC9hM
2N4FEhnFXX6IXJpbEdQm5hprXBCuMM5x5gx+xRGnp3yMqKvQYIVDMHJgnHoX
nXKqsvVIwIVk8yyQvtxMmssFfwou8FbPyMRMRgF0c9oxiamhN8kMI5DINxBW
O0wUJu1R80ARTEVJoZZ9s9ECINl51PjyRE9oJIexzmUue49O8dPEeZwgdXVB
TdZCWzP6/ar5tf4qI/tnGJ0wdawnGVLskaNETq38Dx0VLPmr/m4qQIoofCQg
lN5/iaxXFFfaGza2CwaFHAlMwixTJNOb9hdFXPijSM3o34cB/IsYoPXs5VbD
gwJ7AvV8XVm2KXumMShgr41uIYgACfsFx4ba+jmb1g2B8Deu2mYDm3NTEb+5
bNtwecBdvxqpkHQxTugVPPco5lmiQJlkllwcu9Ywdt+ij8SFB7n2cdbqxsNJ
EdzZ+EwFmDSZ3MrpRV0Cn7dZSZy852P2hZcEYQytLFWXgEzqywrfLSP0z4LW
2Cb+Bj9YLUSYdayEDnGiBDDiT2Fe+bW/o2ukYe2qqLCw4HXYcdT41YnSyaDS
xfd/yzAvcx3EBFJtt8ftaDv/pYBs/WT275MHhwBkH3bJIqZJDhTCmCiRFb6x
XBiwgFDfnHgKmkuk3PcBkzRoVsO+1X3NQY7KSkz99CnUOj/iIc2n7Ul5IjJ9
XySnzLIsF0T2tcxAs40Qt5g3FRejqmVMc9yXg7yGM2Yz98PE9+WNCLGOeca5
siCExRuz7k9QHHCFxPpprxswPySoCTPPbJ1bA0UTOIWJCdLfg1n6ggUZKISH
d70//5ih2/dagPNroY/6UTUVgBQbriUvhnrIdnJpnJA9KWg+WdiEis7Tadjb
PcYUHle9qn+AhvmGwUZywtK6KZDX9oz0YjWa2wA9Xl7fXB1oOPhf/UfM52rT
ue7aftbHyqvSS8hSXPCSnMaDPJvzkHz7ylqsBlAcyhIymDOaLE73p9kLa0ET
J40qjqsNIxiORwkTVJ8TkGsB96U+U4+xQLvU9sX5HG6uTcfGUg5hGF2k3o60
1vcsyTVfzxhvCd2RxPuGs+KyYfgzTUxbxsTLlPu2lHf4+JZrxJUS6ZwEsqou
TRez5G96RyCRm0Szorw67mzPtZHFOxWgC7IgozLx2HRkbtAtyZG86v0q4puc
0jTDVRRaGjSQ3d5aCOAWD7toENqNIp1WPnv34Ah/uQZ5NPq00g/wWFI9KjKj
g/Fo8Z9cEPKeVnJvinXp8VEO17aq/Z5Kq6TWh6tsjbmzSryU6ODdjm2Z6sTZ
DXyuFFiA0a6MXdWYx1qVi8CUAvXfgHmpEQsU3DYe9G8qPtwJDx475UbCGZRO
mTnpJVzAvEqcTSRKtusniO52eW02b0twIRhjx8Cn8Ud/WTHQOWWVp0h7Kvzo
GxP9Ei3cfrnbjNhgEl+RT7Pkvo+ufm8D1SiNWm7iJJ9giKCKV7ajnU4Lqw/q
5QnhdvKyCOTvPo2Vtx7WFd3h27j/VIoLLkbb3a6QPtgo/03Jc6E49aLqlUQr
aAnLUa5e2C9lb9Y20SOGZmNajbo6h54z54G52cKz7IPc/K4SrJuae4DxJ6ro
Ybywb94zqkVcM6iZOSNL2WFEEMa8D+AqCZK7H8djT2jNv8ccXPlJDgG57wBV
71ImkpnyKUo7FNLS+U7G7xy5M04bcReMmd6LfURhcNtktCZ8vYDNKTtA3HDf
dfuahbO1lYw80pj4sZYzZLrx8rLLBqDpG9QSBvCuNxLFHrdSbE0jblAbAfeS
xPa8BywMb3RctVW9LnzBRjce6UCJfA/HswLHrewHnrQ95o8V9KyIRNupFjFt
H0MDbTgp+9VAuBpiPWI44Jr07PcXBwMai/ACnJ2bksFHi+Y4osHrpLSx30uy
hrtoO0h2dmeR91zuvvNxo251mFr2d+0wwYCv/l8s6J0/L01ShSwCfQrN1c1A
LcvVICIm9/eDYUYEMLlnl330JRpL2un6NaZEgEbJ+G01mXqffMQ6dhXxGEKi
Foh+6ac7UcxAMFE8/baYdLBusG88+XUMvBY9EOoFf+Z67816VFrjZ4+u0/VH
dZrjZ+8wGQ6DR34KYC6BCtN4oUhBoQxY3Jt7NIcxjzjQ2AYEhD/Ujl676oY4
XvrXWgHLzOdV9kEe2c8e0DAXI9jJMWe4QhLT92sXgofq+tIkrUoPmEj482z/
LcF5KWvV9TmOXKCWgq7VFQeE6J9XD6FZTzh+GyLCBFUbmar1xA+zaLwmWfV+
RBVSjXx92KbIhX3Nh7xDXmMT/G8Pshgfo2668Yf7BqbuPCEzwZzobAnxaY4f
qGGVSTxiCHpF0fazJ5beAXeaURx9+QM4CmXwnOPVo0YRYp1p8PGlRMcoGf3N
1SSHYH/fpKEXhA2LQ1NnQ4yM0b73SToh4lYOAet7DMpg32ks929fY5NqzbxE
Z3+dRem2tsUKX4ZaB6JzcahhUssAX2kazsZwgYkuvFQqAyqvimXM8qM1DxMs
gniEmQGIWiby00U1CNVOfOWRZGK5KEIl1KsOT+xtcIMGBiLW8/LTLxH65x5B
OnMGOCbZi881j2a6cJUj4THaWiebT6iqCQxfCa2CGNegpKpBPe4NXFfBXSTs
Jh9qsoAdrD3VrSHuganWrhInR5J6f5oOittMSNTyTLx6+IiRO464dC50vanW
vP8fRiT2voXFNoHsQN6pyltmvkQ4g8a84cQyD52jEn/4xPZswIiTpE+kw5MJ
NILPS0QGEFM8Z0m5aPpuKQq3H2Z2fIT84q49wTxDsJjEkAdb9vcZd3+iU+UP
cRcAcs+XfGbDTmwJSCC8m48E6kg/7JpF5CqMxDalR8oQgMDRihd+aaVZBYGv
nZ1+CnTeOp2oeCcnTP6UqJH3HVAQVt+Fmm73XJ9LXoBSFJBFt8zt9vloBsG5
lSz3uODMOkRT3f2XXUStZP7pE2tsNKTwvC4Oc08+wVBjs/FY1x937XF+LDvA
aUUpiWl4dgv5qCXWOUtoixE22QC6goIa+sQE1MM7tP8E6cgLYr7pr2lCEFyE
ghTD7IqCC82AB08b7eRAv1aCyvbxWTwG5Y6pbC6cVWiP6GX3F+4xrjzXhv5N
2X6vaGdrtyDAWr58CyRN6kr8UZHiSFq5YqYWW4sVvoaijyqkyJ+77TvY/geE
w7swU67hYbQ+waVZQ7q0aBovDIURFDHGhM1Li1x/oNpDUmnYHu/S86GeM2Ci
ab9JYE5SEtJseO/yz8GNl6eux09NkgZgVZVqqy55WtQZSYBZ4qFbR5LZQBD6
K4wkipBf87qveIrahzu2OwAiPg+pRh9rJJBtiWwnCYixOVaAV3YhYZTaYsxO
bob5OYg9zWWAa4ld/pEGqv+mpaMA0DoF0UcDF5qsi1AjtJfiI1XbX/0sA6OL
Ir9tlXC9iEstimmgxJtO7CpSbTR+XojlNIiN5PUFUKMDuiKGLe5SxEz7DGUV
mr5ux0a2TrupX7vi3dMwsaGQGNP1OMaVnZsRUsJ10srxWED0ExZCa8lii/xH
Kgo9P3l2+gJlaWszbbBiGuTrOHPoL9eaUy+oWJb+Z6ev1aVgqXXtUBN3q7sy
FWPnDGPdFzroDa5oftACN2kZ2LjUFdgp+tSsvdBAwasAyBkIloRDMuIHqyaS
dZV3ViVK+KQfGzRhY0U2cR06i/LfKpM7gKuV9gz3CkoZmbs4njbe3b1EgaLm
3OoKw+RrAnxbK04Aa/Afgl4sY/UDOSGOhHqC7mzy0abWkKC22XFhDE9zBA/U
ALIVhNQPgC/0q/TIGCLKVfMMN5NbnKoBjvtnpQHZ9gzGDz1ipCkBLc2KxPqe
fLxP96ROunYM0sSW7dVln7Jmrjm22OYLcmXODXzZztVEjkatmvFud+STKRHK
i0/wvVDiKrZpApbb3JRYPMjvycpSdDKIP38zEUQG6Fq4KgoMpF+5LRHbkW7P
wAQ9G5budFpZJV9DBi7nrwwV4qW/qSM6ERXrLV2SCe2wjD20zpG5+eXin17W
m2MJDbTyn6mOxIP/tBTRe2kA3RvSQoUCsF+lwDUGrXEorjDJF9Np8cM/l+7I
rp7Xwfbl6j3ULFIusZ7XIh/SY4mvVTcqBOZ9cve2/85ppY4cAPrZZxKoBLVi
g60a5d6roMMWlmiECLR4IRwsUCObp1cmojeHKZbhLIqysn2ssjMNHtbRHdh6
vzQ1wTaafoi5PMKOR01qiXmK5SkS+p8sf9OO1MFMwdbpW0ZJ3KbtwCnL4vWU
MpkkGXshRD7ixwEGkC8q5QKk0t/VKywgZ3wISiRcqeOwWpJVc+odBxFR37Qg
nEb5fr63G3xKIe7SDqfxk4nMT4jyd3nGcj0Nlsp6cSn6pfkS7ryOWzq2j/L5
wu0Ahw3fKe8DQtLpwszZ/oer5nGm15OV2xUHbllfpg2KzFD8Mf38xr9qXZhA
J0V9nR9hFFXindJ/PF92si7WyxtLvrGbVCXQFerqIFkRS0xf7OE9UQixSP/I
yWS32moJDA/a5Pxf2OD2M0oMV013QiWIzOPEGpOqjYAM2NlvtRdEprg7G9Jj
ByCJ8aXbfEuy4Y4ntuXkpCdCp19OIGTnWhSlwbY5UOPztvqxdNEiW7O7KLlC
6qcv9kt0xOdieHyHVyxIrJvLpvWWYhU15+PmJ2YYn4jjI45E8OTR1rEYfMqQ
+bs7OJXUUifGpEk/5kXkKcGg2kw/iejC7zB+2w7xsqqrS7OTn9/VA1zEoBHO
cxR0HFkZcVTGhQ3JQM3OatHW4fM7GU+QJ7bbZJRnpjp0NwOSCfjAFXf7qQFa
T58FlWTcHW5hCxXaFzEVSKXwdGR07QQusRDfKB+mjOBCIpo5x5USZ+2imo8M
xysaQl+cICBkCU4zcRmmwm5LedDBb3CDHAEH0u4FXFG8KYI6CrLSaj/ISvkX
3n3LAZe6MdXwxJgmho0U6hkldljFxH8ouw5TT0JMKg0Mm9HkAyXOc770wn2m
c97j9GsikjPeEFGSb3yG9Sp2/CATRVMXnqboSyXRk+GJqaWyJipW90oBlB/J
vGnqgFtGJJTlC2Qqv2efsS/uaUXNrKvVml+MDCsKWd/sJMWzXvDJVpVCPEdL
4TQDZR+nxaJ7NJG6F5eQMf06fIp+Fc7jEQQg7g762ulbFFpPfk4ntI+aJo1E
miLCPvGRXiBrWW3ks5RgvkAHNOLqCyrUVMnSbXojqRpM53mWCgZDmtmI+jmo
oZaaJBvDu4j5D0q6JuqJJoQKYrm1WHRzFNIdeyWiRGLdaHeYVOY9ykbvUdl2
PMJOuuTtytN+J/ohCpwCgX4UxrXWDskgR1emIgFqfIhYyhOGCDWL4FjkoWc+
qWVqFLmg0cXaKQgG3XZWLwcTC6c7WxrU8Ox3E3K+zE0mkhi9Rc7Ifm1W9sU0
XjO5r3jQYE5lNGv1cs9yM2Ruqyrm7KICcy8FsxiKzpbQxWnWTQCrqtSZncSs
+rz0h/hY9BAWEwFhJtiJcHia0llB+r5CmQL5zkBT7oQetKezhxXz1btRJmPe
IqpRxi8n3mx5JFtqiMTujT78XLy7bES3mkbYrfjQR5fELLR3LFjEGgz7wttE
qmwnuQWWcOHQAI/k34EjuCdi8bslyDZUaZF+0K1YGxRxTWFm7mITnYgc2AAY
4kobXzVtF9LUDYDFtzFHZaru5tRUxQjZK70XUiW96rgBI5q2cVqK4kcgx1Vc
anrKRV+Z0LPYb2ERVHDXOI3TUOEeBZXVnuP+eFZwOHrf6V9eFdm0NEEsbFvX
LlKDEUMkTPvIFp88+1CGLOaebawHCk3ZKLYGKfwKCe6ajhAdy1suN9HNLaLM
4l1q4AoLrwt4dzg18GsIDCvMs20SCH3lpm1qchD3u3zLHVc4mL3fml24twGp
3Nr1OOooGxyhK25a+HGLpSQHxsn4/x9ABt7/QZNyhDEFduBgOQ0EzDNpSnqu
4YMJOyUzbRuBQVdfogizA1pDXq9mvjOFUAeWymGC6VyORZcOOSCWtouykLDs
5JY/qz/Yk028vKLdXypHWmd55NWD7RclKEU+rvD/bpM4/LCS9lnPpzg/ok5D
GVtl+gi5N8Oq8xn1eCKnfrmBAx9Cd26J8c2aB+MJgTYgvhXzvpJlLsNYsYGm
QNHo6rRgBOo7xcl2VrnL0zMqtN3oYPd2oKbjv9Gkt2nyuM6hkJ7zz1gX1heH
KqJRD0gt69WW6Fc5eXvbp5wLCkxyZHeyH3Lkm/XPLfIUpqlEDlC7DBOIxcvG
u28R57okCvK4RQUQLl9YbOnd6wEE/ByfATK6JVWXkmpcZg3k4jzcdjfldQnp
eziIRAfgHn9sB2tnGq/jQFzWDOWTaK93BIZXgQvrWjbGLpYjH3ILYB4g+xAB
st3STXSPiV5b38q+k75PrYm4VW5CVHnqsLuDgHkjtLtnt9yzPSF2JV3bTto/
vtdt/jHg3fzzgQWQbpB2IktteiDijwWiBxLsELJfF9thgKmMmYX8Qfnj9Fni
597p79WhtP8EAphXDHnLcqj8JvzJetmBvBNOng1mDKXLxMP0OJBCEJcXNKUE
/Xg8zG/I5C6LGeSvzfjgiEf6dTQI7WI/TSf4piuo+7DJYhsYutnortQzwWdn
lp9pyVC2qUJPyU0abeT5t4uPM4onFq2Xa0+Y6YPKV12SJ09MU07aidYmnkGb
joS7oa4MP+ETxT62zc20UbonUEmb4JkTgtiYglhYAReZpqwbqW8xlp24OJlv
J7Jui8fultQyxkW2HDrdU2leKzgxTY4c1zUWmNcLve2d1A6WVJ10CQ268Zj9
R1sHu0GmOzbIdmDTUgKC2bR6Dc28Rol6H9YiwBmTBKGNEbLE0eNyanCdLgSC
AogpCSCRNUCBn0Y50SAE5eB+45ss8TNd7VWqTpmhv/+OAZO+oerkDhs5i6HZ
suA6f2ZyE7UATw2/MCUotorxWs/6MQM2bRaupZJ2yPCGHhXZfUU4SZ6RpfZO
4EM1yM4BOj/mr6kfYITutwz5s2QPmEZOCmMZJ84CLR3/RZd4xuhELA7x/3XC
PY6x79WYtkwGUAktDEPU7nJbJrRBRC6AxhVB+ymw+lBpVMfduHnsgAmZRrIQ
a5G1+eZUNcMAolBAcm/HyPTnWRvjr2nr+94LFpy901iQ3tiD+mncuj3CNkeH
AYV9SjxnNaH2uneqBnsrtAMmGjEtOET12mRfMo3VkjUzIgXNwx/JXKi67kpH
CnEWrfoMjT+PjPRtRpMWsoLR+VSAUKdLRT4K2SpyYy7l3OqOI6WqQ0kxwXD6
suv+8oosJ4p+GfR+h9Y3itueMSvlsa1+rWRX2K3aYZuprIZrl4jakojosoXx
MVEl28xu330RL2JJi7JHktTGSEIh82fQpWCubjmB6cyGCSqr1tbdU3MQI/Wn
sa64vb/vQwclfpQpcjEvfdoglMVPqWmlThxp6OL85EIVyn6cI9u2RNVYVrDY
mjGrayPuAYFCEhmyqenenicUykPseXGDjn1+f5agKMX2eNlG2WDWJghA8g78
6QwTVn1mWZB+97HK6sA+Vo9tZR9kDZLLRJwC0VfGqgvLd7GC/Zk6btESPg2j
A3QoLx3uxHYCY0B2XZ/3BaTjHXuB0NoTpOw56x3QVp/b/2YLbzh3OsaQdeGq
3EfgZ5NtMCvgGlf9aQCB+NJw8Vgoz5ZKLAvJtaS/GC4nxfaKXi85abTDY9TC
85IwZJJr+ura48Kw/npZu26E08tktSgL6VADENJ7C9emhb5qx/KQtMQU40kJ
ZvFipuTgttHmBaanaDPlvHSEUKALADsaAsNOIZm3oShf59i/Sng9Fei/Vi2T
TGFSa41G347frfZON/yNHD5O1v3QHSuvv1WSKUUHTsQCWOkbtdj3QOjaq0UH
CIJ9uWZXffD0VuW5nwjg+8ztB/FrqNJXIqBEn4lV4P/w35uPZSUX7+KU+XZr
HCl2swMvVA8CS0YCaDD8Wf34W224yT77HBA/wZk0C5EUVT1oyEnBlLCwa+9p
Z+JBpQ0tIrEgaVr5Vj8dH+/xi995BwpURpMkWFwSHhYyFvQqtFa8iYndnp85
cS+e6ngYIlPWWkFfgO5YieDcyxm7xfUz5knzoAVPfRcN3W/1l3qOG50fdF6Q
GYhxDHKLHvT0TZA2fsq32QbZxoSWZJgBTjTDdPtf/tOPzx1nMgP3hHYkS3GU
72uN7ess2FmICwVACgCbAUQfGzndH/13y23FlwJqxFm4B2AlF+wrxpOKx1Ej
o9U7QJEFjMn8grRCm6MEzxbCJnDMOASZ2c+d4bdAoFprFDA78KKLyA2M5kq1
JFVmP4anXtdKvPcdg8hqsOiZFDBBDRq4/71+2zteerI/LwXeudlGrcmPoEhO
hNP9yEP9Zuwzr1eq8CwQ41AyvatHsMZy/+rX25XmtH4XmrLW995pOYT0t5Lw
JBzCKt3k4BIi9hQoZ/wiWUM18G6UfvSuS08C4Tw+nvdlu1OJeMH9F5ZoHHUT
SggqJRXXDHiR8aOockQU/gXFLchc8Q1Rt62spNBLra9UtUh4LlzFxwLLR44x
Ae84btF8JMq40uzJW5JiezMwGzcygDeFOeMfeWg3KN2I49wm+JhJEPzkFksP
TBKdDqoBlfPgjmk2Osre61Dym8ChPvvij8wXeHs3hORVgJbU/EbxiqIzDlKh
0Xbof0Mc0sencBORCBe35tgY2NL7i3PXnyTc88BsPdxlfuyEmiFCh6vPVvWb
J6enq105rF20zJoOTB+zmwe20UtpRwQeYlhzkIQIDJiG4jTiOuExlIt0xMkJ
6HXtupLngjGSGMAZ+6Es1+sYBXjP55KCV47RWmZ+EuRhmr/0BiamIgYteAPS
PpKLLmaAMH48xtlHBb60J/NEt4wl711xIX9Qnfb7GnOjudJD/yeEx8d1Bpyq
89sBkqOPVD2B42jQkBIAkVcxxtTS65zt4MvLUQCmmfEWhjK/fc+QJOVVhPI1
cqivxgzeOXPJpLbwR8oewrbC65JMQ1SnLajTAZ6z6vfg4xUKvsxFt0i2uCZH
pEh1C0NQ81i6uuiqL7EON2Xg0K5txz2aw44phfJCDxCVKG0iL+NcrFbSGAzf
v63bndnhkDfDsueZKFMGE6JTsYYuMESUcIaLbc85eqB0oik4Epcg3Cy3W39e
WzGPAUS5q1kcZccDW3Es1lRZGhFEQJ5+L24w5SPaBWRDoEZaHqcNIJjabrIw
j3lDb1qH1MvUbO3u1hrS7UKXIdENy+2zqiBSE/c6ug0pmknXbBPeDPEHDLt+
KOUn44ZqMBmXiU0ohONjfwKvzmkPEDiW/XqvfeLGQn4/l7ldMEwm0CTP0eqH
zwE2uuu7PPDYDP6Y2073lZvy+NtrMg9YpDg2qD6IHWhE4uOkNzYYA3F71dYU
JwTXCFl3rqotmSZAeJbgYN8QdYn7V2Ykl1uCjcU03MaJrDqvo7roV1rG2eqE
9mi0AB/1sZbZ69nu9vqkGldZ9kQO/v+x49ept49LS0p999PvQSYUH7fxxNNT
Eb2i9ueoKn4FD4Wb4Cow8K1CsKDNzuOcdNYMK6lSjLmi/YWAq+Nk17+6MDSH
EhtBVkkTUoIdV50aXIB8kvhv6kwRIE3/T6V6Mtpp/znxkF3HSVJVjK+85qnf
xvrnQoIJpe0umraf1555s61F3L1hoifYicH/cSBofT5hDQaYaq0bYeWFXygS
okBzlbkrBacT5irDHv6F263AEvIX2sxcp20BOeCP5Jyl6zAuwkBsCE7qs4v7
sp6lVUJ06ZM7MnenovS+OS7kZKaS9X6QqxWYSGHFsW554jeifWlOZZLE/u/v
BJjCPwp9u9UtShVI3Dv7V1m3Gexrup0m1yfLQNjHjJMwHaHD7rqjeVOU9YGY
3NDT8M2FS4/E0PjWSnfUzGCQ6ZO/5/Kv1QBWHqBT9r9d0d08O1BYupYKf9zl
bDwK6Qixf3DDQSBOuaZa2Dt2wf8KUFc2v6s6kkivt7isWIwMeH3I8PGEdIfp
lpAcB59Ofg38DpQDLQZCh19JmgmowNtjkq8vUgPKGO8C70OkyuKgRnPnoMjF
aiyD95gCuGecDqXKml/XjW0xyTCLH/v2wYKn9mm0hTjIk7BS+2gh3snjQIno
7h6c+kdw3y6Z05en2k37uARi+pAS0rx4LG5+fNM+H39R8Gp4FMKSyLVcX+eJ
RYhQsE7tyrR4kgQIp7VQwzV0Z8P5JJgho+8ZFskgsZHfxrenu6vtcCWD/EDR
xnwkurkoQzCfa7QYgSx6kVbTP6o9kYOFPsMC5Xk0+MwA3HYeQ9TjHjwq2HlI
vx6Xq2ss3iGhrfEqlKNoRzgxdXuWAHkECQhemlMdvF6+BdBNz+rWWhITwJ8r
fbSNtrTRMgBTBc2iDC75KgoAuXE5mKfnqrSHfdNYGIwKxv2pNBb896tx9z0P
JZdOd3AncmYvAHoMsFaCACPCZ1thEhOI3v4Lr7U0oWWIt2UNyvCqoQUamb04
Urb+/qahpvVwbMcSS2IY8RR5AZj68t7U6xg0tMQENpjwn+uVeTKPdqAkmtsG
ZDwXi9N46VQkckI4wZkiRGXmumDvvk91iIbcpZuA5XyBJ5ZWcEShkANEXIy4
eM0Q2aT+0J8mzo29Q83LbcOpsI8WMd4NZYWS7xM+OafL0wJ2miaQm0nJt2+Z
XYnkzZ6TWmlshXEyjJLn+d86WseQ16aK9KlMRL2nF+0ONxrGSZ/5zXFkb9eS
lICINyNGOEOprodI1itF50wutvfduiskJSZFtxkTyEE2UKpI3/NKJEkC7Dol
j6qp7+5LknYf4Ze/emBSG1yUGgfQkq6lEkB0rcnvzanaYCMvjOcS6fKOFJjz
5PNi2tph7U8JasDc2suc8xrfNYuaYnQwEVMDqgePlZRha8DNIuo5MI3ukPi1
kLwdTLTyf/7foik/o6GWsYFP+kvs9di38wzyQoUa8ZLrkms4ruqI2XewyHj/
9c2cVRxj2EHwdzFFsBg/4Jy1wBo2rhC12svCbuQ38YrX7VKhgwlVOGSLVE9k
IIn3dSTIB2HCFFd3KoY0OM8kqMfYCAfbxvzEa7wRF1762OsnCMZdRzCN6war
o13PHK0rdrupx4OIMc8WTeMSyTLrbcG46EqsKq/0rcKLtWSy8E5gLfOv+Zj9
+bDLoSFOV1bpEFgC2AspC4wWxVPWMgM/8aJSm6Bh77J0LEJBH+f2d4Nb09yv
nn1j3Rkf/AKSTmoRNQ9kjtYECWj139Tp2+cLCppkP1pgSRoLqo3UbavXo48Y
X/JaHVEMRytpg/ZHb814nbgO0uX3HG8VjWf+ud7m1t/ONDOi02T1avs8mrxN
Na9RwbB7OW9xXDrF2xAtUXQN5+MlsK2UvEsjGE0uvRwWbEHOELXlUU+E9DjO
xrN2y6r3CRQ5bv39pJSWgQn/EY28t2QIPJvTZpI0aaBkPAeTvMNuJrevoSiU
AE6jc3jHYiL9jpnD7g7QWR57VhhsNlW48x2qkfJuTjavlOVyppXIuObVYUXW
/+AN0/Vs3lTZSLgG4iFh5Ew8rUuyO9G+aeoQJNssfC3Pux4Bp0aTHMgV/6f8
HA8RxCkCQrIMe/g6oYZAbJl0A7T5umNRvAxMHJO87kXvbng85VmLEGhi3bS5
QOKFPFv2213/YX+DdW5RMZ98p6fyoF0oi+FXs/skuulCDkRXZtSQ1Qc1fPO2
n4eT2p8RlyM+Ejl9NNtSI2V3krir9knUoHofy8fYdC8oBbB5H27vdeSZjyek
RDzS6tc46XRHB9JX1edoGnMCdxgdfStqe/o6LyyIVw/yNXT8Hkiv6LlH27N3
pODoK7pxwen5xNi2qEht2b8LTizCjCWU/peZFCKKAfOgzcOdZ/06roiywKyL
MkoAj8t3h+wHjD8/afYkbI5fB1oaDVFa0VhpVc5etADZqBc2zAqRlGQB+wXT
ZM16R9L/TmiO6n9V+shT0G3GBxaxtwkeWV0ytggVmwLoEGpuaJzPg38qE5NN
V3gbxYUbv5tFhu+jE/Sxn5tCqHtBryoiNmvcd2UHqai0lp9Q7L2HN0P4s7AR
68s5S0SEEWsUZ3DFIPql9pUUsKQHr0DI0Jp9z9Gjt/jpEjCKRI3Xn7QM3Bny
Yq8n5u1dKHCLNQOWDX8xPIKe4sTaDU3bw1N3dc269mby8ZJ9qvAHC5wh7boy
Y1vLkPch8iG8dLNHijXhVJ8Wbe93HnYDGmxepnolE1kPr4UExBYlKrqYyLTM
lJyIVRkhI1OLyKaWJ3uQtGfj8REBRqp4SYzCq24DM6ajXBpWZGxj3yj3pjzK
vCcKdbHbN3RV+vGeMoiUDYNLn3+2knmSrh0iqc+yANmHXZVIGyY3WIepk09/
dEO7tHoYNCDrRWz/T3gddbqbwAdyWC2J4FZyQyA9Vdtq1b2cjrPHvrPV8yB9
lse/Df3gQoeq0i6PJ2EYwf94EKuKgATO1HbgcEI40LQbg+fZePgQAnLDkBIh
EK7Lm60Rp158CP1LShkZErnbDgsRP1FfDXaEaHv1whyWatnd68jjU68BfO9F
CcEywPtZUX71RUeALeAuTaSCFc4AtYquyd49jxx+HQGqQl8M5zklyO5TRpiw
bNrDfIadr4ZrgiFP45Ky39bp3u1nnaJP6nJXmyk65PXy6nMp0Jb60iTjxYlE
6HEMGD4OHUe46NmPb+0AzXKZDmKIB34wEQw2VnhVxmsvp3bwjVJe+Pf00cqX
xD+OJg+wkSnPS5yezgzYrpN6gpzni8Y5xaCqFgbEOIKAWPezgBLitCG1Y4/P
F6IC8tp4CrRYOzc69pI0gZ33vqI4Bmtg6qAUbL0b8KY91LJtc1R6vSMV5Q7Z
r6QMP3Mg2UkMRA3T//FtPP8u/+zVbEYbK99NwUC3iIxSC7/m1HWJPkfrkUHu
bXRTa+10yCvt5vh87f2Evh/dA/2gzJcHGlgkB3XXSHEH5n4HgDxbQ/86zbuU
Kc7Gkj57agGV3b7aL19wGjjb8IKqkUJt1IuhpgmXh0E5Pt9naKF5f5CcCxu9
a+zIV3aGqF/gzkodB7o/BLd19giURiuc5cyD2gO8cq4uYNbcxIbNDF0yAgnl
E7wYF6OHZB6Vh68x0o9P0PtYGbnsuHiEsdxrUUROaGquwJgr2sojRJUWwHSD
Nq+4tECHeUpCYmJWBalkXJqpOU1d1CODmHxXgLLdH+dMpFXxJMtSmMgJ1zfB
lScnVfRM+6E/7RD/hZM1ci5uReuB4CCibd43C6LpD9Z8rlEPb4jhN5pj02pF
tsRNXB+hw2vuM5PbtnS64yGiaf0tflSvAzCKOym8Ev7UXyid4b86fEhMB8bT
6upa34OL8hSQSryCRHNVQ1SlNKVYn5BlPL5XyJ2k6aOX5keZDDb8jlBMJhha
fYpufkXex75O9/ilRCi/Qp6NV4pn9kIzOjQsfS/uwiE9XN2IvFl2Bq+OcLxz
RMtnmn5dG113gQIfCE0Ph0DARCLcafL8G1nxfw/gYZpWnilHsbADcFXb/KRZ
fFfb2Ht9in69xW1CvAleA2UWpWg+WjjkGdzWj4LX+ze+B+V4ik3slQ3z6r/W
KNyvvUcovs2aDLnQFKq73E+YCNPGP4u/a9ZnlMr5ci09EHVRy1isujeDfzj7
voHCRm+x0mHynxWpDv8i2CMXhAtzc+0Ju0GxBhw2skUn7GIhjQ8AMdg1qyDq
J3crn8r3NQ76QCc35GS/oT26i8EH9So99SZuAsu5z4E89gZxAK6N40l/L68Y
dLmLxP/IZ7KKLRamnzsDDx/2QprxjaAECERKuFj0li1/Ibjmp+RqNFdJqTVZ
sLyY2jbJxaF/cXFcMZ8DBd2Kig6s0QX8WUQdg7aoFEXz9fLbiE9dqKvUiYBt
Iw9YQeyi2Ezq9X5sEEB2wrDkGY8hLYP92PkwaikA1wH685y6/ed/90hl4I6x
y6l/G0OW3FyJ87XdDv2FSdFZ3glDCCd9iq5jyft//B6AUBVWSCEbT2Sd9QMa
9iOh/mrtn4VgtB7NJEZLgLAOeblWb4mF3YyDzpoKj7VsO2ouCp1kubUzlYXJ
VAZKpMqRZpa9GluqgvtiItJ4jYixJ1JbCC5DFVxnRIInuLbOBA6/ByktZOOb
2bN/9JzbSi2fKuDHFFG2lTVnrgXq38xxpAbT18TezNQyjpuxQEgM2Z8JPgYg
d4NH+Det5/3Atq2AM5Wly0GFr1SbNrmPaHNO1+tgRyjFRDkjkA4HsarGIFeF
4NdkWnuzCadFvheRRToq8w9iR5IeXc7GTcvRHsEYTZtbro5A2LNIRHVRIPIH
9iwY6/Imu3FbtDUeCvcagUZ/7RURb6VS/8Jpfp97CfvI0gaRAGOgXuKHYnVL
ep9UzQrEdWiubtkRAzIJ/nZtuFvrHlH7DbquQV7PlPJX6T58lgHn6duj8Zt5
TzBY5z7ST27YtooHHR9JSmjYGGoeq4zrKO/KJmEcnrvyg/XB9pzFnMFmFOnc
3DzR9N1SfbV+pgL16kBw1ENz9yg7+f72/mXXGSkyxOHxBHRY0hrrWBDn5N7v
/CxyYaUmTmvn4ZpzQyfxPcuxRLZKVTzGJnKlO9f9RJzuk6+UlvgRerDV+4wd
BpowKzjP4ZKmQhSDLlwHULGC7+/thQuYcfBY4tlmD5TE6Ji2eXGXgvbAUx2j
W4V9oqU9HaAabpDbnXqcD2NgeOVCp7P9vbeEhQN8/HbiFApM9s5OtiKwAGxp
DwogWppki5epMtRocBnLBWI3xfD8Fcx9DxNsR60DaqkXvbxxkI/KyAoTdDwT
2XX2NW7WVhuqe/VnqWIzA3GcPMd1Wg0KBhwkbvQ0GUvigIk46MXDI4HUROHC
cTACLgGntAy2KvQZH5xCP0qDCpoDmLbB3VLgu2pts6RQpaPGkVeNb6TwvYXU
VGUtJQLR7QPg5zLsBcNljmcxv9WJnGk6fP7h868GsNApma2Qez1CFNvxooY8
PGTWvxKwjXAIDHSIOzYwxHG8EmdqWQ1mpchy4orgC8gXroMKLrTSO9a/TZ2n
RJjyI97qwFX6+yb8jHi7L5KMCs1XgzSZRLupObriWwN5gR5vns/0ZtKRrk8n
IVBWVAiSsS6PK9EhEp8h68IFbHuLIPGBBONCMJstPRVON764MM35+Ii0w4tm
KxcekbOWpIXJrV8KOCz1xKvqdpDJo25GCweXoOFEIJoKBHL6sPADpgZyxwc0
Dd4XONU2LaDyd5aVMv03PD5EiwABL7sQvKF6h6mXghPWyq549mW4LcejPleq
okR9cG25ytpP+MfDePYRWV0g9c0+O0+5U8leFPfPSLf48tv2HAhouaKvwff1
4T4lAt/haIikFqUczwvXULYYhh3kwIv3XZTgNSjRQs5g6I2PAEfauz6nJLS+
fzFdbRnjcdTFWsKFi1gpm1z3qWwk/IOZTB7Cf32naAoHx+q8KM1b/owL9Km9
wBzqePb2Ukl2xrmWzhsk4pTVeE86aQh7TsGihNMVA1ix4buYFunYLbl3q8uc
+5RpzX9sa7AunaE7JC/+Dk6JFxeutWE0OOUEjPFuqr9lxEznQFGJkrnTsAup
ZRUVp0tpE9ffUSythtUQMS8Ylv3IkAIk8NlfttAp3fB+67qui5OZRoWKky+P
aipXDdQD8++89hjKRbvuvYu5JdUFJnrCHnvMUkBX17q0UeVvNS09CZHx65Ef
6wdKEKBkiKauo0UpX9KqTywzFzhATjh1uD6o54ceo1O1ngN/eC+6Rv4jbkGg
AdfRR68CjrSaz9t4rphHGCFDeprqDre65ON7UQjKFMf8N0qhcHdfPuvci9dB
JvlXW0NlLhAj2kfLt2a4g7sqiAtOLeylqxi40qmTOLzXD7INATIQrCeY+dLm
3RX8aSUrYjTQL9PYpM3wahOyTyrAJDAXbd2/A/CvLCV4/aBM0HYnUkQQvchG
QFlwDdZ6XuTB4JW3Z5aaxojPNzuiwjkwWcW09/vKPfnv+Q94/RiDFnOA02kC
r2MU3I/5pQVZHhcOZtFNQ0u1inW/S41R0rVYPjms3kv2ldpjilTh2KILfAMj
YYMLW/FEzwMXqdW2HvXI7zWC060NXPKb0Nz6wbtuXf6K3m2mVEYaqjYuEuFF
3VyFz1i+rLrTUHq72gh6ocGj+GtPcH1iCH3DrG3jQtRTIrvJr4GpMouEFOdH
WZDcubqgUCg+xIyDEckbvZPUHKR6IADImH8zCX5sTa9tG4DBnMLl76Ueib4b
qaZi2iUM/U5uxl8ODdsxpPT5hLE1CAHsPlqr+m/BqvIIqoWpZKo7/NiZH5eb
KC38bK82mVA+gTju3wxDqlkG6N9Bozkb3UcHYNjefpQrYEHbQtBxDGt134qs
PLQJ+hTBp0AgQEik5FwXuPrYTNQ6IIkCIfOzSRoe+TmPMlRKfjej6t6HUxPr
09dG3kw1LSEYNOd3svJ0Si83EWWXQfE2hJZsCU7pLX8KjRpP22hYAtK2Lbsc
gThvR532eAuaQWFviB4Ap2I/6djXRs2qAhOw9jDv26lAYBdPWDBU9smHzUvo
P+0nblIE6XV7RsHOdcV4WQzw9saxNjCzHAIPfYIcBJXMbK2yrdP2BDh4jWar
UdWannBHqF07KLfU56MZVfqb+zSatgYbJ9DFM3eWsmrFPEfwtowHJHlOvNpA
Gqy/jGB7AQPMgrWqsZIsKcFaMUwOjpA9VS/jqcUETOW7CiHZUMqrx4qNqtV0
S0YceXWOz3mHeNI83OpL5q0D4wueRnHycOfz9lkLKcC3C41Olc/BnvUP2xB5
ATXK4g4a1nvZ22jD3X8LvsOx10D6gemjZaCkMya+BacYBO4Qp+IvXAd8DuYS
gdCRphYcp5fPMEDXL/87hVJGwqc0ci/IjZqofXhHsEfZojtMsQpXitjFqBGU
XHDwS2si20RoZTc49MT9oVE+VB4IKyNulYypMB6Bhyy0Pm6CjMjg15D3twoL
8V8UUpOk1C9hVTczsmUQjISvRDRu3eov2Krk8Cr9b24WH0e5rJnHHcYI29pI
NcIT6yHWawARLEI6zWk4SRpgQx8NUeElo/R0jKqNy6WXi6HL3xnI7zkcE7yN
zjSa3RzbMKTZA+v2eSWehFCctcHK+xu7becrJCI8duD1EwD+vk/kxfMwgml2
byqih/3nuZt43Y9Y4XznTmDAJ/lVjrjo5A96Nq+4e2faEh4V1shdmTjsTw4z
1SfuhG1pvrr5lAV7VmwY0mhvWqSFivZyc5myBjHFNRdoxCF/Uluh08EkXWeI
E3fpnwmHojobZnuUF+zdALyTkdNXWzcIyI4hKyhNXHG87zbONCd7u+KrvhE5
uwLglDsfaxrDsnN/J7HAm/cgD+19dXfpXIFcU4UQyELkPP4dfs4VuqNVLAHx
3JuFd4ajUUtfGbZDP1sJRM+3MAHgEId88EtbNK3e/dA1UUtFQYQK6Q6n/TeP
42dugXB6+OVzvrJoqTquFhgwCQx7vsQipaF0KRCQaCxIX2t4WajT5scvD1IS
aWTxwL0EoxrzQs7Em5NUg52/726XCOIs6xtDurP8k7B6C0GTaMrcuMtaiNqh
qR8vlPMLtjFJhHkMb89N8JFfGP8rY4MBXKiMxxFyDbwzbZU23eRNXBr+Plwf
boHHW74AxEgl3HB3LlQZDEwynjlY4rzPb4GJul3YRwvb/hjodJgDDf/OzP1d
vWz00lVFsrDe3F6ixafN9VzMa2ei4yYJKS4ViLZtllroTXryt+Bt3LkJ2jd0
VdqdFdnWeVxuKSmiqjUrZtWXGcOf/qT7R0gkyWV0dE4f1K3aAOZSG63M1YQ2
s76neivNUrCHNJxqQGkEcrG3rCmhEpYOXxOKZFINZLbFIVBNhs31AKvt9geX
sts+FaRwZe4AHGMV1rFfqMMwLUCUJv8HjWDfoYmFjVP9Rashjxnup5CpC6Ab
PTLpimbs7NeHXPAFtfMm7LRga+GcsWVX2VXhbcsYV6m/nIxGOobKyxvwWjyL
cMT0/1DOp38YR3CWTpBRVjR/gqzp2/bF+3WIYmYOQioe9zqX3pxYfEQoBbX9
2TXYAIbB1CdtQT+i4EhAMl7uIeT6FCrXnKqut4NpqX9V27lq/fSyc6VZxNgl
RvuQcKTfXrdykMJdciArHvUeJ1vsfbvzCDF7/DqGCaChqLnA8WNDih6s1QYT
4EgM3N36yCWa61sj16OEIe3lu0hJ6D+cIg8jCzLtdWThReXJ2gM9hgnsENpL
TDhQaruOQ87nS3PsZ1jYAVXqjJb8npka2KavxNSOPSvQyae7tNTsNAPCvVSU
+8CgpFPSFlShiGdAdVxTmuP2V5kk9Sv2uaNKKvuxbTKTtzBAjHjZTQhdspvT
AOP773Goz75qtLXLyA9zQLzZopnq+ujdnJm+GE+iF8+m0dz1aqB1XW/1+SNL
FbCfR0TVCeUuuPkrJBhmxCb8ARDiIkY0FPJ0HF5TG6tkPUj5ZUoEa78NC0dP
i2YTcL2aGKp/oc9eEoLYscV7xTxqj8IO08AaTspZuvpxViVarUekFXLy8vvj
KvUNeIEBmkrN5mxu/hwJiiiTAGf4ysum4/1DRmoqQjSDEa/rEzkuhg16tWvO
eUZX96u/Pb7qfZRMpRgS0uYcocGL1Rjxc81ZzLw6rdr2d9twLJwC/2uakwgY
pu+tfxtCevWnkDupPX1C1wZqYUX7NQteztcjKMeDhPTZkR5pjs4v56A210Se
p7rYZp+wLCQkiK7M7YSGPiSs0flPBpLK2zHI8OTPSyShC96/5DivMOiRn7wG
2rSdR2jdZzGnb7SmNBAeaqZ8lbfAK4i7V7seIHh+URQ95ONQZd9ER4bn57wC
GLzleOuXt9t8Ie23F1e539v8oz3AxxfOwpA8dttF2CyD1/QgyQ8NjQB2O1ab
PnpjEBpCTK8PbfDlWeKXuSmbF4bJCTID1GLlEBXOeQVBrL9d9OYpNH5amCaU
6fG+masX4vEiQxuXbj/dxePeMEDsbxbpZGSCAT+4NhGivZtNSg6D5LQvuTkx
TNM9SOKmsarfCKhZLBsq291YASIYJHfwyaIWZ2NAY0jB0YVMUjEBfvrNtyNk
eIZdKwAWqIWFNpECf0XnASnNakTp7qmiiZI/Va+r8wc5o/EgVPFkOFpeqyRI
1UDoEeP3P99rd3p+devEl7QdGtQ4V2vSenAFQiizjXygaNHuZE3NfAwJo/wh
IPv+MapEb4RxwnLSRvYhDSUCYajR5YgBvXEK3+735VjsJ8TVYfpGvqbNoyZx
k5r8jSKljt+95SoT8fXAkZEtZWQYk344eU0sA0G+PgpCA9CTakllampAnz4n
DDs9CTKEUX+GUrFPH8EvC2oQjHXy4WtTW86helU+bhLee3c/75zpppcO+nGC
LxRgFbIIeeoOMZBypL/pz83Dkn+c7lqBWg2vdt+yuJb8rsOvVnaHBJil76LW
kASEVM7zAbvXKSIS3gVFfZXHy9bhKw0OShXgUL2qmKKH3MtpOFsLhsdwTyok
Fl9kMaKz1vGEVsIw2xEZahvJnmyy/8Eh9ZfLvVWMrtslVWEOsSThpgneDlsv
tplluUp3TWLwp9sjxvhZnd2Rv88d00GQ1ncrzgCXKAERyDed6aTgeiOGrbcF
RUHh3UzS0gDvXk+nFNdaXMXM9p5t6G/EVSxcxjSqIYfRTuY2dGtBA5AXfju/
Xw+6RiSZFJ/Z0GfepYTRzTMeuG8S6OkmOjXD8fqN1+ybjTMG1NB0aWnRnDJW
p5KpEtdwCJxB8FSAKj/e5LB98eIgeqH7+f4/bDtmlDxHnc0d4IdT2S/RjS+y
CqqBCKI+B/WnnxaIv/Sg9cWrY20kXcmUEeDiV36RJGUV5B2KiLFmP/4+nn3u
kussEcIbq8zeqfKfrxuYgemZBta6XvCYhl2kfs5ZncK+UVA56UEQr5ETfSXe
lrZBwoef6gUbo2Y+P8kYk7S3JexdmlABW73HiI9T+gPzMXMXuKDkONrDdzY7
8V5P6sD086kpvNptCF+ObvuusC1I3QcfwcXy1di2g2nKeGuu2iCbb1NdmlTo
oS2L1j0daA1h/x/WGEbzs6JMUNQZaMLagZO3Ch8Q5KA0QIXJyEeUM/2EHj7B
IWcn+sdK3KZRhs+SMV1LMdwqeHOL2tF19ceLKZf8DyzDcgOJXs7IbS1XKDSD
avW3TDiXXQSyks7DIp+g97KyMCH7f656+yW/Mpzw1n1+DMpoEoPflGf0MOoz
ZFjfHLRL+CUKinZHe8eXBa7S2nFYPE1ylifLpelg/5kYOGe9zWLfJGm9BJrN
BT5+ExlTAkYjmy9OTnU3tnQ5ph86IzPunT7vkUqIqiKkf2DXobqeafpKK6n2
0HqYRw3ZhrSIIJZy1YXGx5Skm1jousjunF6fmpOdKe5PIC4NfgVuuH3chnDR
G2rc9JOeG4fFGizAFLYa7R7JJn6pC/XOHLdimdMPGHPp12ftTjQm4Vt65rkc
g3j5ximEDsnlyfwvVbPF3HLa1y0VrX6dLL9lTHisq06HcrN9OcC9xbmoJVbv
BhApuf9N6ywQsjPGk7wmQ+0zZd+ZCuZEAoyK+s+bD2NNjlLyZERftykdMEY9
yacMdhxm49pzSvD8Eco0WVK9+tjhzbS/A3c3w5ME1tgRmptELaFtaemSEuoE
rt3A6x81vSDlS9OSpxXSF5GhdAayqKCXJUzYopQ9uxUc1nOsFk6HSA3x52n/
aREwFgVZG492w/tif0Ay5evGcCxCP79Xt7xGm3FfAjGGQygCcpYXFFrLY8Lk
2Q0b3JpNi3fOUIMMyERMR6ivWNOd9CKDziQSF7WP3lNHo8lkDXbqhhGTU46S
DAEGPlLd3KnQ0A1PtDUpIYOPVGGgt35K+5G5CqccQm7X1LGgsF1KMQ0y9snd
FzVb+c5wXDf5ESgLH2a11Z+5yb/bX/httt64beKSIm7twsj67JEJEC+cexmY
3965wnM/lW4TrVVisQ6QBtzpIFpzT00fIwBFuboFghIkInWBX8fPlgeFGQ3h
F6NrwffE4SNBOmkWcYJBS1XVV0KhSsSOZmMAX0ygDJjus5m+/EL8rPS9E3ji
4j9XJW2TOZ7w72UN9UEUPbM+Dta9GWdUb63NrJUnBzLeAQfK70sQ8ufkiHLv
WxyydG2iYSba3vnJZRIW7aadC/kwpylyPBCglMaoxAyk7AFg8EWFwvwqhNRN
jMKFjUjF452K/tmnJtcTfO+w+F2IU4t3/92iwYSy6RpVN1a50FSbNLV5iHlc
3OKecOjIIOCW+83ajoe9XTwJ0mLVigv/C6xKmtRU/Tvhjkz/XhJET0DXauRt
CYSrhOf7YMw5/igk9KK7693qw/xmARrah6msKRe8JS7Eb5CJsIH3NosrhjRX
lriS9gkOoDrV6atM1x6P/P6iF6AZf8VmM2DDlIpSe+inVmyEujIbqsLQex0m
QGdRZzevIh280iCaBLo9KhtQOomzyQF0M+T4YKLZu6tHdpZVs3Z1gQ4dUPyk
YBA1n4WN8gzKzDyTl2Lc0/wIR/TW7qJNJsihKTh6/U2OyGvUFldoXGMdkLBp
g3j/USY+5/5pe8MJk5XRYN8REFDeukdwjfnTIXX+kr40CXJIJA5Fl5yZCCZG
4oeHUxQAL6kku07bkxRwYdLx+ob8MM+5aPpiDk1KRUlIrVPIfymI0kwaGyQq
/pt8rI7owqk3UFWR7knaUIWD5Cc+X+iHTMKRIEbqCMVFw1iNHMBnB1ZyXZRz
J99jHNCd9WLw0cLCVJt2e5Zgeeu5XhCRqgm1NxU8I0U4a4aPUccHF1abI99T
IDooTjs8e1NGYcnn+wtOELsmRypYD/DlEhP9Dj8kZFWclaol/AIRBWdyN/DJ
onV+Fj0A2eMtMnf2jgkoSZYmNrgs6R/ltH45YBf6q/Ix3qTV4oOu7EKt4ktZ
ioJl8d5RA5Ctlq9byKTrMJ5gD/HzDHIg+6QrwE1q1e9VOUgUrc0OTBhYVrzv
JCOJGTSxeoyKFVI3TfdgvpjFQhCJAELTDpQXVd9PCEsWr7nYSv7bX8nSZdmV
cYaS2M27JfC55KS8ZVYt71BovLNLYKGyDi52Onestk7wgNIvNh7io6sXI3uw
1s87/QZFAFaRCyk2G0rc/RHS0VZTFX2j08S2jspb/FrHH2jKXGb1Auqtqzka
DrKdkGmkOsmAtyF8J97Fy9kFbWTkzwVacTElhqkdUAq1Wq7HDmbjCxJhC9h1
yEY6pr2hP/qvA97VohRlQONb+4Dv+XIHxu2bvFhTnlqBptyrtOoqc18l4jzT
zghOXZT2dh52Cy3skfeHK+UlyERez5Skzr7bJt9rf4CeTQK/K6CHbYhZ6cje
YDyvUs9MGFl0n24JhxWAi0BouF0YwnYf6Uc1tZf1zlJ1jOBTL/waKFfqkQ55
PNaQ4NTxaSE9kmscRXGJfEWnRyGrLXLZIg0O8gFqPHIxW7EsRfw5PYMIMRYc
tMw3QMCjVQ5Prna7wNjBrv938/iZudw0ZoIMxB90j/F1lyjcb5MXS0TtygsQ
HXvY/3tCbQ5lYgd0VY9OpCGsglKm8EL4ZHEBV9eR7VcPtEC2qtsyXMs7jjxS
bG19UsQTXdm7xae8Fu8uFBhAuwNTgoDEZ5qaO/vFdfbu6AnWnbbi7azkhw+q
8SQDGefgz8YcjvqYuhAVgZkouNETJt2OHaaYBnWEorq7R2R9mnl3YiIZJJHh
TD3VEr8p/jihYyCKIpHK8PrjYrbsFg8+lWp6fI6SSRhH+JpJlrJEVwfGMiQe
XYLLaqX/g/AkcGFBsPVe17R3c6HIVu5pvKLFYkRElT8fRUfRq19m3fBF++gR
BCHh24EV3kAyrcj90Is1XHiUt3tFwZWRg34YhtkJ0tmsQDcajj/0iHmVIPdO
5FHjsbg+WDE3/hJM36OuFRDv1j4ZzScjYxjk+G6JfntUrp3WJmflpOHDpn8o
5PfwbYqjgE+3REFnuUxrInR5AOzsoP8VX1ygtwf6Zn4zwW1GOTUAUMsBBBja
DpTzmcsDlOpjQUn6mm4ZWcRJGf/xwoP/NPoGszSUcmoqhyHipGBSur/QO066
feCUbjASDlfXzuSxD2Nl/USPZHHTEhahCFPkONpUVDFh6jO5vOUbSxjNc58n
mQtcb7Vdvw9CbGnlmwPiR8Qwbi5618Y9AG2+Jf4LtrFXJLbo9LMWULK8YmVr
oN7WHRp93LfbhX8nQcEMH+hutyGAXkN/Y8R7ZoOgtFhP/+Oy7BvGOe0UmksV
Ar2vRQ32RqNGV3nlL92+x/XMJzoggV5Orv+729j76EFPQz/CG/u6KJmbie/y
cHShM4teNWnN0mC2zsWOSxAVbt0+VK1Lmk+O1VQx4tTYTH4YBBkyAbYIKjy+
84QAPtKVdC8DvV0mDklmIGZxIFtAc+e+izIucACyQClsVF3FLNdQ//woZM5n
dzm4xayIst8ob00VbuW73PtU0AGVrlPeahO19fA1AXOX2h6mHJyQ6GcLsuG2
fzTh1Dw07x8vNuGryJsEFnQYsV3yFOL9VrtNJ3UdV59k1zY/acy+sH458JVL
/XDGsOjz0AGUiKtILDpvHkbP8Iuf45d46bVUGtsG6QYW72aAX8xgmyeonQll
6MoZyuK0C2YedmJ2Cwzjny7Gvp4rye+G2cPf9wtzXcvKUmYn5eQvBjYL8wFg
FQbjcEaw8FSIp76Skjv05ftpmzq+q1XEoxlPts0ARmrXmucLh32x0T1YfXm9
kKm6IuOBx6wKV883F6zH3eQo3kXaRxVBMPnCx6DWARPnf0zKKwvJOx6OdpnF
gvUhJGiSu0qnZVl96CSDXIp9H1gt+eyU3RBHLbDUKsMPy6LzvPczMfNtSXkC
VYxXLW0JSBx4CN7WrowTHOXkuc1Oh+KCVupWAJz/dsx1G3MO8+KUMWy29yW7
kqL/I1DbdlaTtE6Ahb/GzVZ/kcYVKO+uSCbDFXBwvPDjwTE7WE6wHeAMYq7v
tY8xSOSyWbm+wE1QdfhDg/7kwj0QOLoEAGJBt+mnvUQuhumsIVIptnKVc34a
bSipbKKl01fk1IC6ro2YLgv06W9CsQwZ70zr8j+584TB6E3ykfpBBLljJLJl
q5d77mkcdEMrJpinA8kK9IJA51Wm8Qx/h0tz0FEJYoUvuk92O8HE9DB9dAP5
9dsOJG5Q1rQ5kDiEQ95kG+0xyqEm2rhQxOtd/rT5Qy2nq2GouGSzaJ9pfGjR
5du4Cga6Insqw5Ze1MlmQyX33QW/8CjOHx5y18HFapGfyDjaMQ38kI01yQZs
DOFbXoT5nyri56cT6MBY+lOrFw6UJQMpn7D/3cJBH8K8zzb0RM07iKGpdF2G
ezwmP34Zyn08I6NTbKQ3Yngy1K91XFueEqDT9T67sU49jboCZijs5uJDhSO+
pjjrvcPPlwYciHG5YL9KpYIS4yW2MRZAXlhcoZO7inntrJN19hG5qIK0bKAw
LGU5+hMXdUZyxgg6CIT1zx38IbgnKvBfVQpdGVB3DUhOqmrGa3xjR9cEEaOf
ku41XgP71VRw5ghWmzVScxmF6HzLOyTaQDRnzw50OxaD+H3oSLGmeCjyg1gP
OiVeFHfw7BIu63lbGcZAW6XCO29T+fz99t08u3qVOP/60tmsKUpkvRSfrD+H
N4QD5VeI5wdMrA44Z4SkuGq+CVCW35Cmpq6WI+viFrHi+Z2MFIO832CEt+tG
xZcRKbHBUZ74gKGYTtW0UcNmeWlO+HlKZTtGu9w2y/V5nGrHZbdcp3JP/O9V
RDTJYWBr3ngsQGbkKT7QZmfrEnS/FErkTObpCj6AeXKQPnpwnmdb+oI2++Rg
9b4wr6wE7T7BDclR+MCbOb2uvGGhjHtoX4HGLk4LIymhC7fmUYESMG2e3XJn
0PouvM6u30qN80jOVQnN4V32yi7g34M8htXmj4je5fdRI17N3AHjHC6jxADZ
QWESGLpC3WeFwwggdw2xITGaraoyp//ZUJONBPdTo2CQMJM6xofggJyr4ivA
Kd04myzuOS9QCUXczXDPgho0J7uwcbOH8v2FkUs3tSuWkdEir7cnNB5nRZhR
Q+xMlS82pR8UsB9+BdLN/PCek7rqOtXw6uN8qp9R9GaidPkAsPfcR7vCxurr
kl72zUG9lUVkVYWxjW0+BwH8mrx6BjxT/XhkllKnXa7ZaKmtu7RHVN1hahzS
n3idcKgIJ1JPlRbPDdjzgyVymckmBAX9LEc2pNCU2aoZstGDqBeClz6JqoVz
jXhzmnyrMfuHOsk6mfarPxi/PdzSTvPOV6tDDWS+sQHDUMlZPNB5uwzJVVXF
90jzZeyuuucbxaC9vGDiMtrNsJetbRov4RFG7lF0DWist9lJUS91i1V1x/KS
3GSfiZYP4bOy+3L4rf/gvKda2ucRUh10wB6TXXNXTOtsLKcrgacAbvwOap3B
r2OYTNcYF/tcWddt2jClfW45/vGp8ykiXaxio747rmMJibGARWQsGvTV19De
Ot0faiikR8huQNiRJbmFE9aKHLhfJKEZmbu2mvXX+f+dLb4Fj5/SW8VQbvwP
soErJHtnkTW3x9YDFOwt7NL0uA05qGui6nqAKNdK6tqmTC3RacigMcOq36QT
3qG0D+rp0EesWZtjbSzlyXwOSCzTvMmJpOTl8E+m6Kpp/cgE2ape2e2mAcvj
NFbKw1wf+IoS1Ir49Yve/4MZ78T7Trh/1QZmmpavvSJV+9LDVRIB76YeFF+5
qDDN+LLLZsT/G70MgIfS7aRcnuCHd+/YB5cLjdedsvPuVG4A93+XDd6t/i/r
/VBV+4TLfvGQV/u18gF4LTG20n1A1ZOhhoEfiPpR1HAZltQ0YbqEej0xAIU4
IQ9ovDA+SBsQ6n8//kNxlUpVWUTL10uUXF4bpFixQd3Rmp6tykkGmYvnqLOC
tJcIH/M47D9jNMDwpsXMJgb4/UEk3crkjD0wyzqAP5dmSX39KjiFePxNWvh8
aCsGtpQnrTgsgp7S69N5PyaGyG/OF1Wk9z2xQ1ejPNDoM/VuDAZZd8rXU3Wx
cXjW3dVSZuxamooe30q5A+J4kq4vF+zDAV7GSH3UOMH7grmimxwfTP8VO6FG
INiU/dJ6n1J9tsbK6G+UVNVEp9g2AvcLqZhLCy87v+MQMZjhu2JJQJ5aD5Ik
chfZggoDs/pOm+rq4F5ttpiDmNH94HrVX42aoW+eVlX5udAw2i6sEmWiWgFw
giFH3OElaH4GRe5zI5VigZxgQ8qxr4RTVQ0X8hRunY+Kqjyq6XInyLzGwcD5
y3mXZOlqsJOOkuy5+Y4/tfaZNcwrLiJYkP2m0p8Wn5y6f/YbeDluc+rDPR+I
MkSQKPsv0EIxX5P2vDYYkvwZEApfXyHFEpYEnfjlrmN46ug3bKChwRuZuRWw
q0l0JpekYDDGwwKMsMvwRP78/eUav4u20JGImuiL2FwvHWtdChG6IuRO3i/T
NHKSNa0HzL2PG1MF8K0rxhpxck1GVHXSMPGrkLOxdaqccJDtsAHjBzrg6g3c
TAlgQrddPL0TiwIRLSyIj6cR2ElFE34WWFQ/8suQi2GGOB8GiqCCAMAzMQWT
heOwHruc8ZlKSm8AAmv6XWRcS3SVR6i6LPrhZHU1uLn9+tLfH9TgDL05bczi
mTI7OCUS1TX0CuXO74uRvLKMdsR56ZP0M1DNI5/NJ8jQpbHpWNPC16z3RuC1
9r8YzROzA3qr0hhfHVHnmUlZmEEpSdAKj/NUvRjAApKciGlUCOwka5Ra1ezd
fz+PJhvP0wVr+wbZfwdN/u5fVuMRmJAmKjudm3DOb+TU1qhPn8u1pzWrTLLK
lzbUiOt08YLHdLbJ3Lr77NoMVE5xfdYxoTL3ZqmGrXEQBUEcOkxiIPA55smw
xL1gwrESm4UErWOsNPajYMImw/ZMo296Z1UOtCGfJxk8DvSmr85sCh7HZ1jp
+O1dTuu54fqiv1DnPdnAv5y+dyJtbLPf7yu/x+uk3WAIQM3GVTWrcPUAPISf
Ttj1SGko+niddK+Xu46aMa1SptwLDnTzQsK1lwsUhA5GT0gBpSGkd/QJjrHE
v8Bq9co2dZE5IMe9wh/BX4Ub3trzHewpTLxVlo8Cn7dgIKKxlalVdOmWAmVn
ut2bCGNg3EJZG8AQLJfe90tzRwMFwtZgEdFwoxgkT+emCg+bSIHcFxBOQ9bp
WJ0jODBBTpjIft9ZRmRKX1TcFm6d1h1uZWIJBpGzgARACgYwGBWcTsOq2Yh1
N6tL3eYap4ai6x8rYjjfJRIFint/ofREC+GuKl0QyvcxeRevjdfl1m1r6euk
qWWk6XzabrH3vNyEAocAyvVUE5CNPs6GvsMqnJa/w35aygUqiZh1peirolcL
bxWu02S2NkssAJSGXL6EgfUnpO/c68sZlmjtOM5OvSvTbBkDxriNWpGWdgtt
1STOxqW2Bp7uS2jN3ZlJcfKYjKJDNhaP5jfdYBjs2FJI9+hL2/GqYFSoSdHD
f3kuPDVzm97E6e9WqO6TAuGwh3SbKNHcB9jhDjsWgiI/wo4LxPZ3KPxHXVRM
38RPuTTCytYwKiPCfTHFUjvniL/AM4renIauPZJ6v/41LRS9q3bqdB1WYPL/
K9TQeBAaewY+dguVtFfVCZ4Rtsc8Izn7kMsVClrA3gmUcwKr9R+ApaeyXQKL
F31+JQrOFkG6FwEkN5S9LNBa7xNog6WhOFEmVkcoc6UTzgnsxe2+mNvCqex9
bvSW+IjcNoLqhB3qYx7ZuKtj5PWo86Vhz5SgENxAXyl4VL9WirUY/N/Zk1+5
DZvsLGEWHXhrV5XuVmI7uA4Sbpg41TAtH2RRku2g+8L2LkTWiur1iapJX+Bp
BeodYMizKTMNC5/081YhCdZN/yCtp3PliYBAh3XvPu8BHROw/E1IVsdDyMdg
G7+r2vttU5/Tkm5F1Yxnfmy0xpc/pnmnxBbWnN+MIFbt8v86S0x5ZWtUZwdq
fCRrMAty/Fsvkd2NeJYKn/C64LzkVZLxteZocxtNp227GqtCbaxGNMpL1Uod
ojrJG0vln2HkWNUDBiHecAI9mc6zJAz64Z9dwP3T1Of+qGRL4y/5VhFAHy4y
trdFqzH5JnYPvkdXHyZkko7GVnHKQOFElchhZ7CTPRBcbo8x1Wpfibq0Iecp
jhFBLio0weR6IQjAWaTgTeMLpzVBPVAT+axHVmD7C919uCGqnCKkE9hI49YK
cRQs6HDmr0yk0g3Ys0p/LGJEuMuAa/S7YzBUhZYmdaQHIZO2wpvzAPxcnHdk
xEyi21zMTeEHfejd6GUhCRJ1bnxuwjl8TfoG0snHGTdnmcKquYu5wf1sncFU
7tQgWX4j5bq4akjSJsi7Dt78fFXsxfeunMgtPowRJJb/vqqijeshlbSaQZQM
9FrKkQdn47hlEbsmiQrXMnS2yqmEb6fqJkzs8MFc2o+NaUuPgjbeAYQAKrlX
5KbVqi4edJhLFstaA61zYNrwlB8Ln083xSOBmBlIOTGH+3OYfY223PryezFd
Uaehw+igAYo2zM7v16HunoYDfiUAGzDs4iKOfFtQNRxL7BBO0DBpwXNrAvcP
gDUcmpWPPzUPYzrEUHp7Sd5uXLspXZjl1/z9n/J348NdfBVWGz8fe5PESpoN
EjyYwOmRpCKFq83Va9N6GESOfFgOHWzeI7crz7uvYMugyZZskFwLc3820dxV
aHggyCOfOHGBq7rxZBtRPk7GPOAnaMUpWWWZrm/K/uSLvwnDsTLJjFDa+GMc
wcors+LWQbvw/zgpKowG0NzPmvT52y05yfmhE3LqdP5Ljhjl13N4uyRHUhEt
O5cxCaxmEKTvIkfm+UeDdZSAi3bUs075UYvIhVI9lAz+XCGk5J07No9rUhNG
uNmsPHOyF2Mm76xGMgjZzwzcSrRsjsK/ShVRgdpYmic+ppQMmllQ9g+OQYvZ
2n3Pj1fXShrCCXHMVCFdD8+Lie6MyIMumd7lSAa6UPhB83ZLZPNRBykFqLMv
42OwfOX2tVgd9kulAcb7+SCMGFlsDIkQyTaPYJ1nWS0J0ntDBRbCcU/QMyzz
7a+8/J5YopgYVUgwPg6vg9cUGv5Gs58QMupAeAhInMHBD3flEVi/vsJA2zqB
Y1jQnMCjbwSnfePwjWXW6o6URFMnzOzp6W7wzm4tIhzRkUTktP/BdVCrDoti
pAhx3BnP3QGX9rBN8Nl48+HMFfuInN56wwq5XaeXvcdetaSTyVuEqIV8bWvZ
WpLFf0r9luziSpDsdhj+Ch5Wi1knp681a6nESVmRbAIS6szXjZkEkQW2nxY3
7ob4sxcGQIG3xRwfZsQSwl2Q8Pb1hlsni7hNHG0BE5oXdgUbFgs3XRGyG5d1
xXv/yv8KslaFuZe3P3o1GoZQmnQllL6BYkQcbSHRz/mB3moRaSKDa2uVBPvn
mPpcyJ1m/MMeLVKt2uornqjrKVPMWzMBGo/Is7qBO6BJRAuBMHRWjiyVkm5k
E/6ndPjaGDVS9F8d+oRdJEsdZjT6jiEPxaVqK536IxJvYFlvJoakxyoN6cWn
8CHot7W/7xxSLlpc/zPNRpZBK4DE2F0Isp38dGJIZX62YimKSzLlYckPngI2
+MqKWiQZckYtmDPvsUZXFpfXsf4q2FO47JHKWqx/4EObIVOW2leV20q1AECS
IoHSLC+bAZwZOdthcLqbOyNxILNRJEkE0uS/dHo+HKMU/DX60XJXdD/YyDzP
xkyrephDoLuVpJgVayPs4wLh9G2YzJhReR7nRGJwcenSJ5buY/yubjSPeeyE
NKuENbYN/W9Z1tRuzmFx+8RYsQ9blOybPCuo1Bd6jM6LL7MmhuaZnwHAZ5+f
zOTjVrun4oTDVZNOun1l9w9iQrK9R+xbrufdtRd5n4Jf+RJZEJluXvABPADI
HsN9+SKvczMO3Wh8sZAGOgzJ5eS1Z401Y+6w/Quy9sTT66r7O6UybJOoZZgk
zwJTLKr1L+HE19XH4grByqMgwHlg6rMGiF8GX5sZQgQ5RVBrJwnMhTlk2N/R
Ux0GoDMtaYO27lWyuvAGDdB39vJFJxfGCXKdW7yxm3efem+FI4lhfTTvm18Y
/3M8nOHMhHGK35f/onAfIV2mM8d/I4MsomVILieIeEvWzX2ur+5Cpiwgv6w6
fTaI8QYkTduLevpqc8jiGbq5xIBzumrwshRW6k76BHu7XyyKKML9+EH6oOyX
F3fZ++Mt00sanwU6DeWQ+1AurO9p0pKhXhliWLykmWaQ7ylBf1dTx4Vp4fRq
RlZSisbj2AWOF98BzPZ+a/7CCH4kQ7o+dkaeeVEtlEs28AU0rfvZdVc19EVt
eyT2Jtbw5/tUTOtXhWC4DV2207SLvSUP+dqctdxuoWuVowhlRyUjwEhyI6Jf
PjhoFlA0XLuJe3Mk9dcUainYN5kAWFtmGLvkExX7Wd4Cc4xPEGdaV59/bPI4
Ncj5qbDlmf3a3JXCoQpr7VItjyweTUdRG4z6wZxdxzmUBP3ArG17VdnIJq3u
zwD6M0MXav0DZPw8FfE3tB/krD/HDYZrjleYTjTTNR+0yc5LjVTYtHL1ABhg
LkqS8bSIk2/t4pBQQPmmcbQ2ukNQ1RUErA91bJURphAMli+VPYqiZOaHMX5Q
vVuS4gxGelfA/Ssj/sXlMa+Vs6dAPTouKThVoWfklkJ+VuMLkDk5M7dQwzKL
3HI4QgNL59rFasnxQ4XHrTI2RAjvj5CNCSUZPtmixdCljPP1/r0ViZ58oSnl
2ExWdfQ1ftHQLA5xPxtuI0ZbBDiSiG+AHn5z4fqe+q0frCnrkMC7K9RfQgwv
peW9qsOGS6HUwSu8vhpFdJw1S33yknnUQXEK2EnpbPOCEJNh2Z9X04yTUx4A
G+GktC0dVKelIQutu0J/MHdbs3JvTwiio/bWevH31R7UGoIb9EguXgZER/NO
ZrIT3RwuqGVeck+Bd+I0rQc1WO++lT2NXT6zh1AL4p4a/k9r9cBuwtDqvoQ8
EK53hw2CBjvxQNAYs0r8SnefIYnrymHU60gJqmZorm8YAsQNRUd2EV5hQ4Xm
T4BvqvFZR6kdlP6yzVxFUNPMVkHEqBN+W203n3fOLfNW55P1OZyouvkkja/1
XxxWSlFIoSQfWyVdIGD7V903WSAqfTuZR/7U66MJBOvTHh53gjVVfosOU8mi
Unq3lnuwCtoShUEPNmtqTbmEzjyIElqTOs4lFrXSo9Ekv/heXy4mNaaI62Wa
UGNYX70NddB2dQi9dLkSByGUSGhdDkL3V7PmhZo65KrIHbtx5EPq2F69nJX7
Ru6NJAzB5ycOGvslqkuZn9wDYyaidW1rfUEJkZXmbRFJDlrtHLYL4xHs50PE
d2eCvyhaln//MtnnFLc4Txv55NsXH3jxBHrEURsA4ssTVHigHI+yB5qaHfyg
L3micRplGElK5FxtI5E+JQUthCwNhvYRRRH4OOKYsONFC/ctQwcdxLUTeLAn
0RdW78LCpwqfb2IxXce45pB+FxOKRXA/u8O9VOthJYlieE71iiPgdmFKiXaB
RDM05Xxmc18J66aYGcGHPUoamCv22itiRLTiWbGWYynvKFGGomCg0tZUgMAS
claZYggi9l1z6z5cpjJJAvHA2GdqxOMSWmSLZIetA545Bls57xGb0LUPmBF1
xg0Ghm4lxo6GLuUesrmrurk8BcM6hplWr9M6NreldnSdHyRhs3A6vdyWzr9w
NWteeja42FziWbWudFJS4c9Xg+AkLKCcVHvlgzRuaqB6lcr4HAkF5EhydHAM
YBd2Rs/trdr/9v5gpWFvmjZafdBIPey9wS+LgSksBczU6VBJ/uXhkFaIUpww
v3CUJeORBD4vxiqAg3rM6lOfbxzVdW/kicQYeDRtymeOK+dbysrG8r8UJTjY
JP3jp3c/1qML3m8OZM2JgsuJyGbrUXJAhWZrVl3WqBxzHbcs6fk8ovZk911h
X+OHrcw6dZ0XA4dYY5/Ap+mgZgs/0F0M6iaTGwYLI4U6coMvWpxnEZ+Lid2t
YECWxOotCX48xPRa85v3UjWGBUUzotTKzDeLN8EY23IYx1J8H+rThVpUeOO4
ubHXpZ5+hbb1CJxHlEAhQ0ohLabYDHtv5ASNfIQHbHkd5KcFzLfIRZrj1ZOh
yNNkf8HdzThPR1Il4sin7MlgYnNiAcoZgoCzvGJ7NtGXX17Gw6ljCVy5YcUh
Dw55flOIj+uTu1mMvHSK5pzK5BFFTHP6/1xiTKLtWj7QsZDoPHfPPbc0eniX
NNY0xiljSho7Q9n+PdLbcW6zru43wsBT8zXxwL3lCv+7T2oU/KDij2+tSgNg
SCx5KhEoeIOIIYSAJ1T2CfEO2tw/agX2pNKUKBNW3xt6mm6E1yNQeddBIpZm
0Dr6wrBuzPpIfYnSRPXo4mG+YNhnCvDkrGfxbVoUMulGulhCacpHIY/rQg+D
7sfRM0A1XtfB6sPraJuyZ+gfMCloiRgEnx5OcvFS3XS6tuxfATkT0c3rK9bF
Sic5uuai7HtXUstBCvxaRLcevbl5wAIwAMUDsqFkJd/pKWc/VoG++JttGo9G
UMLG0KHpUnzFipzSFI5Myu/k13kvXVl6Tm3fSJPM2eKzq4T+kg/wsRLe6bX6
EIk7ZUTjqgDZQ2nR1eVz4RBB1xmoUwuGLaR8e1s7BGRr3/vy4ukFFqv9T9gN
LD4B0uI0YDcMhqaNaTwhmEaQ5pliNmuG6b8hxhNzbKLPoBP7vBhTCfs5ZUAT
5Z77rW19LAARJf8t5WyzKBuOk54HOLKWs0qPzXyf6TyHunMOO/l0fD8lveck
t3Pnyfv6njpAq4jEv8956qtc6g9Aq1Fth94XKxii3YQBoY4FDXf+AnL0jsHJ
u9LqzhOhz7n7A3OxiZmyYEHzVkEyf4+6vleEcvsXs9aFFxQv1mlqXRGjA3Xh
ahZVh5ouS6Gsph9/HiPPglGd8wdUjpirQuF4e/nziAd+XyHVG/VcStgiJ7Xg
n84HCI0Pcb567UKDhTAoakn5xE82HT7BXlEG/7EDxuV/vJi0R/5q4d11aaAH
a+pITFsd/0dPPs4zf7EhB4QckY68bwmDwLbgNzWD0zDNR1uTC722+5Q5vweC
ufHjJ0g0Al7wmxQxnoCvTAXZ3tLHE+V2bmFSPkZoowrjMlDCcGsFffYTh2Gf
3ZpP4z5CTf8Zk/mILHISDTR+yL4p/n4fDreNuSGuQrGnNvaGRUZepa7bFA3s
jXXYSnz63+RogUV/SVbv8/mE9ti5zqEW3C+HIQbCzyu9teGVJCB35S3OSH0X
urAJNNAFIlBvIy1RadLHMHcvuOfmCo+o5O1X89FWmjOxRZRCQ1k7zXBGNI6f
8WBfvsJSXu9fiSfzP+PDEa2AETRw8DDQaPZrafo2t3hxlYpjuf3ZLG3MyKuQ
uGa+Kitkzt4QqJD1BexPr7oiLq6qI2+ANJB/7d5WXHA+bMVfYY3h6khgy4rg
/MUF8rlR1z/YpRu68EkGcAVb63GWTPwH3oa+vbDX0qZQwlD+Br7h7T44f5Uk
z3/T7e6xC33GMsWU7VZFXrJto/pQMyV+XZDgsYVdNMYkqy8TMUSBsuO8iap7
QgkBsu8aPPVYn7jK8lC+Qv8PDZckaIdvh5pEOTMMfciIFbqezccg6tesKo+F
Uv9DHz2jEJknjLEyGj//EkF7w0DrXrulKJOCRdNCte0gEsuzXAKyX6wnUEk3
Gx+mhmcD1/+C6B6OXra+SJeeTfGJgfC2KHrljdw/jaKa++yy7M1+V6lLjyc8
guUuV7qxAX6axe1mRdnwLtzR0LXSF2H8Cc9MFonY6ob4ux2Kn/oF2oPMKpz9
+3qo7qZxpIfif4WS2A2+JGXuyOFfgRTCmdXDS4oeDCO1l8y0vVERzHjnCdaw
bzZKzjjtFkzHYOI33nb0yx7d6tuCmeqLKMRLqQeC0lC9Wihh8WCtuQSuK0Xf
s7PGGHVxcf8HYpmJ3QsKdzAGviuCKzF8aPcPr/P8wOUAovrBczYSXBP2mvPV
tx32R+d0mhH3LdvSyULO85wcDHOciv1femOJSHgpHNODYpnS7rBkkDsC1jMm
sHazGb9/qYYInRsmd5rS8nIFgas0nbgzYhxEwKzTF+WDNZI7v9e1XI+8gUYW
rzwxLfkvaUlbxfMrh5Vd7cNp77VD96V6wEVbW17sVpRBX8mlzu5J4SaibgOj
GJ0+yqpcVFtLWJo4xYPBHM8zXOL4g5ZyZWnaoWyfX5mPVIbBrFa8MeqEEksr
hhUbwuCzhQCfYWcKKzKZlUJi2D1PFKcJ7KybUYtyuiViYCxPIRlEQ9bLOPTV
DmMSHXfo0LJDJO5xII4r7C8tuOvqQzeVYPDc8k+IQaw46hT5FAodf6+iZOkh
J5dsxfJ5VGD8FMKqd8NzhtYe8MGVJ3laRdyKb/zaZSEsmTJ480yfXfEdBUhq
Pzx2RM+1ytPZewd3K/JZrZPbqangZySElMlVRtcvVbGO1kzaHU8oTZHC41p+
dEh0avSTG3mmKvuFudyU4t+NNaZN1S32v447XLhyZNfh9ei+2LwbBlit/com
Htt9SheaO2mRLB9LFvGXF+/dwLZD5gBzXVApiJri6EmNHso6XJCsx4J/e6Rx
c+H0jz+SWGxUT9UFYSIVH7+PcizYxr+s9EE1BNfIP6NA43XT0oVwE5qGHBZW
SfwnrpNOo/M68qcvTsFG7AM7UjCfYNJlqrFRn9vwWQzl3qwzM+nQohR3YEH6
Ts1KorSs7PpL4yoiTNetRWx6czFqoeRFAtPGM5H9aEkpxqscHlFi1PL4RE9O
iJlRpgwa0j3NeEV52ytweE+4DNlkw3R7VvdPGqkgS3Zyc6qyI1l3ci7Zlu7X
JyONfS6z37K8Y90PVw00MGNHq3TSJMd5VFFQIe/anM2n9igeOz5n70bMVTIL
aHBM0gHujB1kqarkHKkvGG92QpKMh++1xa3xNGWYiPJR0RBEXwvGI9+Tc2ue
KOLxA1UxTo87CTHewFCgt0N9+IV2nhfxvULom2Lw/kOJqAC/bmuFFNcHBXkY
M0k1LiR2nRHN7pBhsfgmP58w+LE7QGyWSWo5i0diz6asijQUuiVeu6PxIfuZ
X3fiaY/Ed/4EI6UCIntyju5mKnqcSnHL/V1JtnkTvxKSrtmEVhl1mvtoSbe8
1PZbNUUAlmEGS6SOxhCVo20GLNPG3ruuF6AntOxitrNoDNFin83Gq5RK7ESd
XAkBUP5kpt6A3SHtnwKFReb8b0+rUiUkzzz4fMtF+uGYICw60Nhr1xWl+f7T
zo+udgg9EfEZD5k1gksy98kwNwKl9S3dNiMbfPAYMxmW3WAW6ZT7blmhlG1N
uDeLdaR4k18Zvg9KRV7LglvmJYoDpyXoI+88YXI++nPiFbMjDxcvbRQZWmTt
9EyYeUJ5Z2A6bcArc2v4wQi+gFQ7OG6v3LSnKuNNcaUADclmoBUIAyDd+lwD
SMbx14rIWZK8Wtiw9uDuVLkMRSXuA+ospHUEr/wXuDnib2Fy+3gjNiD7Qmsw
6ouOVoxWlHR2JZKcrqlkiwJ+bbwTM+q9uB68H091R3Kc5P0K77rnDG9sVRd0
xrKj83y43ctHSzi94qxyE4SqcQpGO31cCvb0QYCLSZoaPquZvpFTq27VvC5a
Dkbf1YkDPsljyg2b+u0Vs46POBYXBbun6U5hsKi/JpTG7XP8d7E0CZZ6R9T8
0VCooKXosr8FYSy0x0mURuUH/Bowx2Hgt4VZ2jUnkLJhEDO3QUxKey5v03rR
hNBfFwyz+oUOXbtuUl7+cuHtYT1PpKTmFi0oL/w/URI1h/qMqmS2p0HxtnER
ursUJCfZ3bjpnSgF87S3Oa1sY3a8xClwpyZMNfDbfm7ldPqldu95M0OntViw
q7T5ATZjsLm911sJux9j6wAQUpsmTr58hDLKHJKPSsbnfQxzuR2DWl7HWzWE
2ojGihpGSw/rTXZh8PN08+W5Ifx/A7y532imZ7s3pTx6KtVaO8RvOthrfv2x
AuyMT5LtlGbjwh0uPnygpt1PVKcUhhsKOusknXgn2E68oW5JPoIAgU681Zp0
n152WibiVL8n7wcqDzvtLDQ+9g3AFi+n4M1hEYQXPbFrQMmYtbiuLJOiGNQz
DgNWYI/4SmxWjZsSOWVvm2JN3K/jSzudl7biMzdO1hnJ9+k8dIEME2tyqxvV
2QuBBuAdOsuXKoK/SFo+STQRrMV7nZA3DLnQVs2VEYm7mMuYMIfPu1wXiR57
xCKtaKj6P0sCBc/0zmKb3mOMUJCQ+yapZdmPOpLicx03tWzP8OKKpdLgnvrd
cTlHfDFdrvJU3zh353UV6a4jSlTE/T0B18xjNjZSH6KVSKSruyrSDSBddzFT
zL6I613MLchsE4mvUvWa+P722icGaJEZxnU3vRv527rMldn68mcOm3x5IlQ7
aN5BHAmewrtAW4dne2RuH7PDuIKpkXfik35V4RDvFlLbONk+giwIq7geBxFm
bK2BBj5AOe1/l/i2RI4dDPhJ1oG9sHnco4OjNkLjN2dqrb9UYP4FGvxM7Gfu
nrwS3LiKlNXkdum4lqNpAvdLBpw/uA9O7dFfmQVO9QsjbeUf3Yh/pDbYReGU
44+N8YMgFLL3u4UB2x1ZOR9d6O0HUBjoAvi9zVbJAsaSAr28QPsATIcsVQSj
sd2O1GMXgS6PeeITSwOQWO8ULRqp+8skv7zlYEC2/5N6unq/BdVwsMXc/PI4
zc5Vs/CCypoNARtPhtDmngFsK+aODA5tyUTiD1ed6GpcCknDDIhGvRnOTy8V
xwewEScyX6yAyxaPwtJmnJfmxjttRZC0rGBWbEJwdkUZvfq65jZ2M30M2hvn
GeiqnfRixXXNK2f8PxZ8f3fPrFZrr+eoCGWYCfv+12UBHDwRWb9Y59Q1tWr+
+LAgmGPSQLirTZVz+HosSYPmaFYSunfjxg6xVaArgIJw/UTadtNl+F2C2/01
K6PjyBOIFK1+pUIzNmk35ABWDplOtMWF9dmomHW87tflvuLqlH/7pMwSGNrQ
wUVASXT8X89ik4K2Sc6NkhgHgOLY5oANqIjdHZZTlJ+MPDBea97PvlNAVjN+
Iw4X8lVed2iHgAqxqqQlHIfkfydRPRC33UYof+7mXMU3jvYEp0sg1V719asn
ARQ4LivkRhtY28AzJgeP8xtIJJfPm1o241C/BYP5n++yE8vAb+gWpCQ3xqfm
4dgOZOOHSZrNvJfOB3C0sJGwbaJitn2mH1JvUxfXJYHcLoFHhweM12O/KrBh
n6MMV5YaUN/TM8SO0sS/EbR5mQUmh4+32LF2uM9VSZgAx4P6HK7OZwR7X266
7KB4lMUxMmZ7u3Ekg1T+Vdas6C001ieMZI3XHwpHkFomez5Uu0IeHsmMAr8v
5pz+Xj5M4W96TWf6Kgx8DRlH2JN3hLiZ8JuAmtOxxPm0tYT1Z1VENsoWKkC2
ZVt9gkIVyLjBLxoIAfxJ2PcMmTM5E0xkGDV/0Fp1Lo76508qEa9ulBR7EaG1
iYDguagKtbiHd00tEZn224/xS3U63Rcsh0NAtihdtAB+PwaBQ9keLi5NM/cC
HOUNu5WLWue00/glFeTCELEE/NzIfMLaAmHfVxq7WGZO54wzhtG0IVMGCMcT
a5wTHuVQ9SzlXnEuGQO4ni+5R9AknS+49BXrpmiRAcw1KcqhaeHChTbROj6T
rrhl+7YHigr/wb4Lg+R+dztdhS1OJXgOcq8wUt4g98b1istS/uNxBXZzFnik
AZDI9Vdza+3A3gSdItcYECbRJXeZ+2RmGZVfFNwOPtjLqA+HwYyDjnaoMzzE
5grM3mI1NERJOjCpNp6W2m4BvGY3htpZM/R8OCpmls9E9SZ/4wZyYwaDWStn
A1D+k4rXl8sWNiDOtxbrSiiHqlL7TMBcj1DEPqWreYv5rK02JcWw3EQY0dYk
ANvvVbrsKcxxe4+6GcCLlcM1uGUm79NzZkpg822W6Pkn7qPiuubYhUU3R5EM
UNIvYMOGTNtpoljGwjbzt7/fn6jNzsMhhoU88qxBm8x8upheqRYIqQIsNquo
VLOO/j1w62PKW/0lwd0RgNjIZt/iRIsiZci3rE5/o6NBByVSi3YlDVB01ctQ
uzFcd0AQZqDQDJ0iW6kkQAhm6N0bM/oxYra3pbrYE2VYVVaRbaGL4rtEEQ4o
yfnzP3USfialgDY+zE13CP58iQdik4x0QOcWwH2p+6bdrlP9fU+Ak8NfDmYS
sWCRxjc3J9jb/5KXd0Lt8mBb42oTBDaC1Nw4HhCQQP680q8jYyK29edDQAko
ol3SOMP+0lZIt7StirjfOE00jbYfYvxFkCMzpzAl9HcLOKZQb4LgN0/P6oe5
A2hCKmMCYkb+7LgMsBN7VXlmuM/I/XaeqggQ9kgt8PjAR0AnGxya7P9S9+tI
eZ9+i0tb/uuFm1gsMPD8cRnsJEzslP6U71KVFU8E8dhZrMtJAWWLlzqoGdbX
4NQpuF90chqm3hYfufsaJK1/dzCMQVRW+/DMc1uCV43v+qbSDk4REliYOiqp
KNrZYSRYdRf/E6YB/Rqe/Hg3aYt2RONnTU68SBVvxqF69REl0P2JNfH7auPQ
HpBKE5Bmwv5NB5js0lgyXwC+kFof88al+0wWRBJSdaoVJH0VOwzgfijKRUwn
swuiNAmPlh7Nu92mauhCFTmki4q8Na/fzBlANqbtkaLIFwR/QJydModAhF8Y
aj4fTouo17fguOPDMg8cFpET4zC19Li9LcEpFilXK8QnS0DcwWZfgFM7iUPW
l0A46LKzTf8/XAXEsG2zydF4dBgKXTL9lPJ18sqOWEK/HmIKhsSVJJ+Mv1Qm
KC78FnsE7ssqcNwWltwc/1dp004Q1nMTbYHtxbIN6J7fh7PQbGZuB0gffWfS
mxqtAEqJ7KHx5+wtrXngx8aahMp1G0NweKBpaZ/7QXD/y368H8XPT/VDZC55
7q8fqDMQBGI0+mDXyUowNTise8+kh+nfdnXjoGICb8iZm1lKwoNymb02a0GJ
nx0QzZT3cBJ8beUFpFkGtb0FbQzsNRwHGnaX0llspWlL1ava0M3sDAvU6RGq
LXH/qoDE7ZZX1hgottVDHD1391AbBX5itsR5fpzpCYqlrG4C07s/qFz33Y3v
/x7sGE0QJGBSylw5AG9mo0bnEe7Lo6KzA9gYCRM2yLK8aXVPcV9gZL2dRUVL
Qz7RoF84zel2xg8e3v2m0QcdYjr1NsBv5j8seMscQHNaWu4Oq5lCxbU9PKnM
R76dj1SBu6CeFHxggLwN3M2IHXFc0A1cK3kA+RXpqNnRnYD1vCHp/Bakvryf
Tno4XnLlTH/uhAClYCUeMPG2YucsG5DkIcltvPsyFaJQp64jvUB+WrbiYy5+
Yb4wGb6QZ2UujzbFBLH0OYatpOiU03uRJrdKVJM5WZKFVcSpnKYnVIvAsCPL
2GSUbWFHyrWMCkCjZSikOTZPrbnGzLss80CiFL/52AAW2AhSEP8gLeXVxkaj
9uh0e67a5Va1GitE8EZ77pQyDPuHBThNuAFgEB2J8vrN9YEpLxCv5ct5MWQj
hdXPB1fNuD4RChDYV5DxFmrSN0dLqEmsVbxKePCgrL/AqpObRiCUY9GkibAV
Yehk7lcT3kx2ZlgQwZYQIROVuF62752mc5MtzFO4T/R1MMadMAgpnOD1FrgP
uJpbU10mm1+oS0ycnp7WXiC8VwlKjlwYrrwa6c1Rn613LAljKbZKozxDaNes
YHa3GPxjL+e5ZHi+xt+DueW2oOl8z8fPJOXQ1TytLBOzeaCVcBd2r62JTUmy
8uBDs74gD6edI8Uo0G462uKNeWPkHorxlGeas/2McfthkaL9hE8UPSOrxyuw
rGcKwzSEsqp093+RTEgc6L/ZjFHw7VkG8vvfoZtTEpzUVHkJnBliU4ZRo8mi
GBwoHyEIuXdWfDNodIpkdfGSlU8RoAklW4w4c+lQpEgBHF1bcBfHCPoE4Sm4
E3Yhd+DMF7nkRhvtwFFkvJMO6BwVPJ457yxFBi75dCLSMVzLSlYbQuNP8uZs
dKpjmFO79IioQZQmFwWABHSl4wB9RZ04/3zb/U0SAHa+yGSfQN4RRSWGp5iO
67535acE5Wj1kAw9bw6M2C9o7gKNbs61OnfC9HstBFSwbEGfdwE1pl3x79ib
3ejzYRu3tpX3drhCGM7wdWRGGlzXw5SVVvBuUTbNvl/evPiNxxPyCcSgfg9C
iOOCjWwmdLE1wC8EJ27XG3ox4Tma2/d8FRKHbPKTMzVoDx6+k12E3EZNTpML
6xL8qRsSg4VCO/RBigxvi15tB+PK8+vFRjqhVg3YV/o4cmuECgYmMj29ZJJv
Hly/TjysB7ik5M7mPq/8AmElRjcqv9pd8++lO5utkdeahbJF00TrY1EOyH+j
wKhFzGLMs98/TUg8e0oMl8a9yqNc9sdAV2huAmJn94vSS68dk0jIHK6mpLk4
JTwP4YBDKZguJm/oK3/13h41EwLbJ5jwDNheZBG9vEr5nP+uYTeqwkflNCBW
quGtTEXWRFsUtwEIFKLzM5YOf0lnY4qH215AdH6IZXQwzuhaMpgWPOcne0EB
7MT7HWARBtLwxiQYlpu1EJhsjsBob/pLZuhwa2YVKd8uvB5poRB82y4MMaHg
Z7GR11kavGEErDUkcfN7iM8CrYW5wso1XlxNWiPtK8pEd+ZBcw5zurVddVo9
LtcwTYfDmnjc3TsITqlBLmLrNFxhJkTGTWR1Gabdh44ft9+YzI1JjYz9ew8p
bWGwvSguFTV2UEa0WYEi+dVfJht4AJ8RzRTo4NAn7WBv2gtv7oBL9oIVv0QY
dk3tL7WMsnLC26jmdKSwQS8TSjF5il16EAb7wHDZkSbJs10LfiqsvxH7FAbE
ckcVx2snuMkb2IEY+X11fe86dn2HyGqay9/7vtlVi20qiQKBJGmyPvnU4AtW
PTHxdgOgDsBghBS9OFwAOQWSmO8+GrrpVQ6ph4C9Q3aWjwNpEtpZH+LN1eNu
3nTyXCiB48nBIDvX3WRNoDDMr+aexxSuSjY+qg+vKUIY1+7emoQLioq+B3Pz
LL3gAW7+JwMe+BU9H27C1ZBh9bdjrlxtkiTZhQ7gQNKmyJo21h9b5Bt0zZRY
cwDyKjzVymbi7D51wxGJlrqBYqEOVZtMbuuQz9jFtEq9rbpmPyj/t1Xm2CN4
HNIWM1ZqBQJeanwP3oZZgjv9R4iDQ2gP08Ubin5O1g2fTKoce6xtdRtwmIDv
qUsKT5To+/Fjfc8lWtxEBNZWN+9Q9hCVoUvJ0IkY5ivPH4ZuyfsyP7TxGi5F
2jsICrwQ6iQs8LPMcrl7lu9K6g3klWAeUjTLqJGbMUGNsAoW7IHeoMhdIDEl
Gla2AyK98Iovs59nQaHNB8N2F4fwECDnt5fTdFKv0vCKgW4/gvcOPnRlYHJN
4i/D04Q2OdvNtt4iJnGNIjt5Er0262koOpFpdTQPzWPqIOFFJX9W6VEp9fWO
WrkPJnYxBpmNPoKKH4OoWOeCJE8bRXQeLEvvI9IGl6X2LrGMr5IYyIn3QyIx
eEMZ/nbznc8datXzq0A+G2YkJoqkW8Us/dMTDJ+1wzKnNYbN+1C11wlRIqPC
p9TwKR50ikl13748d92xU41zkXT5lOWyaFEdOF96tbv9t4hhMaium0b+o8rj
C6AWfnr3S0ycQtPCU39k3W6ZzByz9DMlSm2DFWQfEVSHQlK6Uuz9lVv9Qfdm
RTVdunq6ovKF6BtFcSt3oR6pvzDj42F79RYPQixnHoJKJ3bOUZ7ILUEO3zNj
IKmGpGW7g/yTJHwHkwq8s5Af/0/paYgmapVLemPZsoH77i8+xwhJY3DRoTHJ
1bTR6jzXg9GZuVhcaxOb3s+9pxvuCkJvG9WjMindjcHOO4+klswIccRKouik
yVei165kspmKaEQ0G9oUS23AOPX9xSqmjwLAb0d7sFPbBwPBYP+4WTFX9KI6
IVsIrTAxQTnRTJij7SkyqsH6Fgh1zcD799gNpJzpZBe856i4tCCCbjNC4ceh
XcqwyvbWw9BJV16PEtlOrICHIeCHfAMWII5SeUwMnFkzkivOpZGBE9ta72yy
vsTG7Blqe7aZpKODr4EXRn4GxnoAVzfsMgugJJhj8frhCkdSYF8qATopzoJa
1Y4PSiy7gg5ip5klnYNcwRoQAhZn0GJMT5iMbhlQnVVSzkiY/prH+0CKfny6
KxxQm+w5/X9uSd4SA8sbUYyQ4vwvWMHM8svPZapT6IsBNXOm9fkLD7lCGsnI
FEZhTqrS7+y4F7NSxp784K3ax6/OUacvNJFqkIywJlBrLqVyV/rMDJBAvBJW
g3/6vupeL364ko4ZH6yMbOBISHa7C+0fvgbPace2Df7cED/ENYh5mkaYvn42
PZs8RZ3EfkxfSbponVmpaLGwiWWl22ZOPUimXwvPZheo5nKVZwhN3fw4Jb73
J8guM/kB8VJjy0LxMXt98CVhTvhub8xQ540ZKuJA0Gu2HQnOVdAua/Z/tpEy
sIiETYzFbq4htrPe4e966bRAhT3JmDN2AUlvN3RTH2PpeaRyf5GG2KQ2p59y
2wNz2qYNPEo3RFrICBK4IS/g1GOTcrIbHtsjOYUVDI1qd2U9C2jpivGbjrlh
mYWNiSbROaSt/AkFcGkbQBtOSr8j6PXutTZAGGTF8d8/22WUSQ9KdYaz0T3m
p1ArDXglTGKRwYNqa3sfsfJfQ1fn9u2Ssh9H3ytNm1nEZgkK8RAGGK/HBF7O
L8LzXJaAzuDaRKc5OsI0EpuQoCzl7Y3rSBu0tlgNflG2E8yQwIrV7Eenwbsb
U+KM49ma+83WbBSY3GWPustahhEbcxHV2IqXILZjrfo9B7ifiXuEQ6t/CwnS
1krCOs7FZrvr6XrBjfh6vJDarC3i1tURTfxGyCSK/ZWQMImytV3fAtRcmdpF
QIDCaAmF66/zqgtdbaWvzHDKfqRbe7FJGmCUzak8rdGu1sd97KF1P6EIGq2Q
Q7wBQOIQOcBPVtQpxXKjk4A84YEACxyknhDcwU2a8UF10xxM8d693cbgytTC
Ah/EbywNOLkpSdkTd7DdDgXBhtQC4c5nqYfD0aALZHwZy16Fk/7mRl+qV4R9
HwHzJzegXn1COQMbl1bH4vLWluiTswb/ZAqZlNA8mup8/Pw9EdJUegWmIMus
NMW6Q2LMZvlx7ylpth9UcsFIxzeYbv9C9u/ta+UWstucNbnhVOxtIoOjHcJP
uNhkFIYJbyVCVn+t4W7WkQUH928so546KKFiaRNdOGqPTTzmBTF797cSTfss
Yae62A4W1VOtIsJo6XYgcT+IVCvSgGFJbR4KI8hMu+8uZLU1G6CTs1Fs+k4s
t0XGj2PF/unFM8Q5XgC7MGpq/gz3ThwQrwApl+1qAldAhQvpBgCJm2L8IDBf
+8OjZN7aiC3/cUnJyaU04H/wr85ttUr/OUO1bEws4Ch777qeNkZM/BxiVsWk
YSWmUFnb7U5jeF4ZNjnvoPvHKjt6z+CnLsNwKjLyHsBhDL50M/EuwQkQZNWK
MUK9zIlA954+diMasMFIhyYJd/JHf9WABouaqUy7JS0sfFLMylb2aFlQ2d1P
q6wp/HnusuhBQLYIjnKVA9t4cLlVviMrqsmsd2Tgjml78wBDQ4eufeJl//fz
hRrMv7Odmu99EH67mlssZXoslCttJaSY7Cl7l87fQ27aUmvKbGcjUGczRpz1
s+rMZLXUoI53NON2Tm+0mVrRykLSmBlOr0rd5Zmu1/o+f6hD60zj1m7Gkl1U
J5plovi+XWJTSqYgkxz7MKMBiYzbV0afsUqixbYPtCM8M0/0EKfOKB2lSyd6
V1YvkhLtY8ak79DnXV5+kxuWa+igKwfaf67cy0DPhCuepKp+xRme1FhxQ3Bh
nJDrrfDS3zrw005zPO0FuWfnjBoANxCekFVIl2cUfUF1FaJ5FmUO97HXN17l
FLpUdR/R3Fw/yTDYesZQH1zywWWo8fzEch9TICTiECc1M++bTb2OBJDYJ3+t
uv21guOqYMHl1GBkEmC2O0lAaDKYifVp59Y/FtYyyljy7h0FXtMdP08M4qJ8
m2+ziYNl6m5zoyiCmdnYYMwuYMfnbXjaksW85DHKAP6iXbb9R9pICjM2LGYf
e8OgVe3SVJS3G8ifBOe++/EVeNevOkHkMzfEkLqC5N+ndU/nsIeskRRspTlP
a5ih8FiomJgRq0QJE1xR3VI5iyIpOndrhkcxzrNkplw7lwvl4Pkmzk+gFx2/
PblkVgojagLKMVM408tz7rpfGHPgo1WncZ5mZOlRTAEnAdv/PQpLafnHCIEv
3DEwwz/dw3S1BaHyGzcKo2eteieLTeOK4nmF/sY1f/k9X1ChhKH09f0m1sbG
0fqa4ida8OC03kM6A6/nXDhXvcmze9dOnJ5gMwHI7h2nTL7bCN8vwcyn5qUc
vDO8pVEhvYt1GZqNEV129m9QyVvZ8CX1pDrwVyssDqoPqDcln9BvzeoG4+qq
4mA9QjZXw864ZjkH+AIJGAD/CkxoK0eaaa29I4qSrumbvbJrHZwd1frXANgC
SaP+8UPIw61Jwp2rF222cHYnEVgx3g7iBsjDfQv6eqCfJ5e/ZBBJA93fcQ6w
a8WtTWgThnHpd9SG8OVqZ3vsKFU3E4tXngEONp2Un64/XOF0nH3njxjr2Zj0
+cLvtYskDSpwjCMvHBe5r8YpLyzBFwgW6K68yYvjPRamtYyEa8RY5hIgl+Y7
761BkGJyb2zuWsjGeroZlPwahTrNFFsLzImsuZCoXEP80b/IH6GOUVpEHTFd
MP9mmihHZvz2P0B9VHjITICbTKFJDwYS3XSAVkwI/5zNaDxCwIGvhVNmMhY1
PJEFb+xhKYCZWTZbWJIxo8aFU3/IuQoSjtqbkTHqgaEfAMOGb9UCy9OvZMc5
qd8fQsaFexYjA4UVYjIMdFz3j2GG71Uw8VvNYlBbE6hdbE+e3X+sVrzPz2VU
9jmXlp7vx8XL3wFJMkFzi06R78oAa9Nb92CVhpL+ouKHkVsi8ovKDJowRG9f
Q3/OAJE7WBxASDb34cxFl6lQoQty7o2jTYgYyYuAqWaLm3+Wf2C+4+4yytsa
CkksWEjDulj2cXJGltGHwredS8j6sW4u3n0qK9XkfXRzBRJosky80KVekvGI
4j3HLawyqOpJtuf56aPHAYaAF0zv5+12ERUNUl3qnkRI754kiGv+NI6jnzHb
uC3eJ7tN5gYakIuQ9ZQQZITDjwslR53MjRA9uNFspp5jCxzDtewEJqNbtu61
ALPsS51rUJNuCM4lrZiXwD+vcCrWpNa0x47bT4KEoM4wS1Pp31jLXRa0/omv
CJN76zISmmD4AEGXeboy1+OhdUYIT/mp1F0iW7GOr6oPCGxZtc9ldDjUnXvU
aWUC3Qj5calckaSWa0MvFIqR5ADMyyx5Iw+P6yemEs27C3kSrrKymGxFBdwf
u3xtFqkmBkEO+sL5LNtgTnpxkzqRKmscr24dCmoeWOnNR+idPF5arf0N+8kI
Nnzu+aiyPV5Rr6NMDEn6bk8zsF18LmEx512Z0fMlZtvtQ+SryxuCN63Msnj8
kEBDgd+9EWsCDN3A2Za2V/u1n2P7CJukoU4axzdcTyP9I4mkjpnIrSnCP8Xc
a8uaXSMsR9OdJ6dTcRDzm189D9iQRJaMgRlHbHkLnOVrQA1JOCvrn5czOyP9
BEiolL5t/vZdSrtE/cIu0wiv3mmwaOYEhTNxtIsYpz9iuKR4LZl5VZCDGBJH
qFma1elOMSEk2kt8g5CVsV9upcrMFMMeFMPwrNSK7z6lLsNKrSTg2A/lFvUG
jDZCCB/DG3oRoAEIjLxtRDtu5iAG/X+pOj1DumshHBgl5spTVRCuz+y1bwRr
hLX0HUkgknJVmHFmubd9WVKEEHCejWBpzMCkoBLd90bD/1+Usk33T1i7tF0s
oDP0AJoRzAgUbnCcVa6OvhsB/adjod0ZSsWadCY4V5o6gaIrvvPchlLpnmrI
YY3LKSfgJYBr2mtGEIo8JsR7g+ZsHS/jPJw+e3L0/E/5K2qhdJn0dYX4MFd2
dXVCV1WTFoqf0f4teh36DA/lOAqIIbaaq6mSYIBdriYaQJYKQwS9/ZeT3ibv
AvISXSgY+7c74sjqTTUjrjar10dd87gS9e1xrym8uGPD4+LHdy37f9fJ1I3w
2cmdQs9VF/shZ5hMJICqJWXgUp9gm0yWl4FhOik5AvmRztYDvqgGFTIkJmEc
NytBYRpWDX4rPlmkWCptjBAZOARkIMncaiT896/THk3Wiw+YoSD/Oy7TC8UJ
FQUgQiRtInFbIEG9W7+l0rfQjd5Y6X6S+qbHdpy0LsdrimfEzptISIW1Pe3+
eJMdnafKTq4ZdNJchzBiWVJOTz29fSIapojo9t97OICIOdULFbj+B/vONFOD
ZFI+odH0+vCnx362Ll1mqsDr7wcgo8zv7aTvtlLMtkwgQJOBprT5Z8HWiTUo
lN+WikTs1uyE5HyxF65riRX1L1KdEUMdBwwnOuDgaNa9lZftrKcDeq/w1DrU
OV3CSIk6qaVZj8qMb1BM06AmPQG8nneX6hZTfm3fEvIRTdTTVR58mjdC3W0v
KkSuFYT/rWPpzbkI5cCp/kx5E23qZPgZux+7OT8JIO5EGvI1LvJC+1rPwXrC
G5IHyBMQuA+Q34AQXLvhWDNJ/P+q4ruLJFloEK1kf9yndb+1AR9F1u9jCtC5
228XxXLK4D5NElVXfT3ueRdRWroUH3n3hSuFspx6/wU9AVCS+QUv9T3zEjMs
rm0JkMml9DTSTJ1g25899sck/XIQJ9nGlENeRhjrr5pYWLWq4WwMS82Suoyc
V+gX3iEG11t0Mclqmkz0u3hoiDaeo2fuONBNErXyRjlzE8yp05NTLFPY5UDY
c+qfAzerjChsc5BEixpquzm7G8UDH2aF29vTz5KX81JHjdLbmU4bRWarua68
IJRYpcsB4fIdGWFIfLLdICyuGgaSnCZz38fN5LhXhp02RM3Gj+kl4C/jYiHi
WadlVx1tX0tPwlXpH1bbKXNWkK+WXcg1wYd8kmKht4Zf+1+FVs5X6yRnvgWM
oiqlzMdaCG/DRLy+ao6X0oOFfHfKG29u6ZweSVlp/aJa5/UZYZ+YZtQM0UCX
7ph19HKaPK/RFDtDs2Pcns5REeQbh6JsZobtdPzLHQrhpXk+D35e2MTdOgGq
P0NMCyVj0oFmgstGBY4NxpbGwnn/NnvxJZ0RQmU7ofHYXa45FafvHy6IYeO9
HM5UqyfLzcPG3rPFSDWIinaoI3xxvoPp4//lLmknxw/htFIINOAe3EWKDSUw
tLzicDZj1oiK/bZBszkOaoTMsoPDimuPTbuwoVPDH8QPHrO1jES6Ile+434/
RHiXxXiQVhZpx4VuRRv209KxRu0X5V3dc4O+TonQ+hJLNMK05RWiZwLVeW+R
puh8gdSNGTkqeSAtkKB7ELAtcSj3xtLP/Dh51tlZ7Tvr5cemMqmnhcoLmwrb
1d7nTsSjg9Znd3WLHjmV7pZO6/t00VZXsn8kkj9MRREfRyGHd2MF8YCaZFmO
pdYrtXCfXcn4wVXUHg7BnJ6cN+aVxvMeLQPztPrie4jQN+35tQZKP6BSQ2uF
dNwcHYn6OOdkx4cF2EJfcbI0bnXXvfNNLZ+QG9A91undXlee6Pyl0vdX2Hlt
sCU3Ott1TP30aMzmJaQVVkB/shroHQIXI2fgcydd1iSR0WfQi4RPzIc+qotk
k+FjE8+cKa+eccKSQnuMgVNhUnDcIfhBkoGQZjyWqwV5vLvJcaV8AdY2wP9M
/L6596v1TtkmZzRWDveF1xq1SWwk2kyVaI+EQNw+vynopxFM/Uzq0Eu8aRGO
0uz06RNZ6pS0JFwTxxMSHxxBy49OvUEAXEcOaDfNbWKxpPUA7bVCqtvwEXzy
uvhLlR+tx2k/ti25Q/eWWCaAihGRQQ0Oo/gPQbLMbE5WgLNB9sZvsq06xvwL
5cYTGe85UHnguPRCkE9EEyI09hX254GZQmkLO07XB6eH9bpL9BnfiLfrtXqE
ACEbZwpdjjKsDc1XI1egWYmqxVBK1XsgnDGjPh23ZmDJ3FuuuuAHryQeH+3A
60XrKhHh7G2ZQ9bhuvRLG3xUd+H14YpXY1LLCJ8JTwBaDIwNSd0ebaqUQDFy
5B0NR4Z7OG2gPEjTkvYUI048SAsAOYw/hV4K1uATjZ92FzAARd4RlDitMOGE
5DEEaNdX6rvQuh4T4DqZ8uDhq6VfXvmwLMi9tQ9+/0NAUOc6wAMhWGkp+ELV
8gzUPjtWJGsmLvB56WtX0bY35bC9XkmUVHSGppOi7mvf6ShWcypVDsg0kAAZ
OhE1ju/JdBi+i9gDFAizsZF76NqPcxrNKsl6SFZfgpdSsu75t0Tx3I6yYex+
SJjJe+9pVg9TXAu5MNQ1fgZKHNIl4tk/s0VOO+w5NQ1964FOYfYzWaJqo0rF
J9GiFws+ftYeEG7b12/1OaXjbcAi/q1O87Y+arHcbq7FLUtLLnvmvDLHLIiE
yQlCr4lLFXhWVYn5Rz9GOsGSB4S92xhNxMF7Hs8cI+ckQZPY/1wDWC/bk1tV
XlP8MeQ0bZLIIa8936JWg7MznwkdZveRRFdjtVLmkTXITmx2epQeUrf9CNA0
8QSP3EmZG0igtRb/M997AFNIN0Nh7RI0po1J8FQpOXH7eS9p91WrLOCWotPK
ncKeSKyoUPyPw+AsjKXNwe7JNnQwPx1Art/t4421fHq8VEy0JCuXYqerlKYK
56dsfUis203VvFC63XMhPS/sWOVfwnUwDJmZSwjBXBI/BqTqrZTY670FqX8X
3d7gyomPqISJPftzd503/l+6kUyC0r8md5KrMEEd9Ct31d+NCZwiiQ9uJFIa
jABvMXOuxRWl4plK53kyX5AXymQx+PM1aDNR2Ikvj702vXWfA1HHSyi5Rcvy
5zsJ4K1IWDjcD6Pbuw6nSYupB2UaeED+7KiH45vWC2NspebiYH8BxRoSD9k/
SzF5BUGboFqhumbbo0TLpNmodbez/ZyauLb/USh8k+bJrAZ+hTZtsY35neWT
qKPKLAx/rsktpQrrobpu0xnQ2zd8fJQeB08gHhTdLVQbeho5gZwXeUwilwKP
+y33fn13VgKLP1ytoIpo4OtNQKndIrzRjKmQi6m5U5n0rPR5Q6NQN0tSXtAZ
DTtufVyKQO5kDOoaF9eUC8yUH4b1JMmIpLHnk/OYmE6ouFgeRdywkXoEJgJi
fqX9BSNqzyorA8qkTk7Y6/XsWJ9CtXV7w4Xe3iO/MXlGqeVNZmakfAeQ/L9F
NyU4t8uL4HkubE+fffOck+TM75vmuvT1+0oX2qv43MlmTN8Oll4xGikLCQAK
A33U33wUEBPotWQWd8sOdzjszDpBiv9nOfeRq3lqo+NeBlpJbA0AAFLvhInx
AiLMomM2zvswngomsl3f+vEmrtCEdtY9EBAtCVA2/CsqskL4nq+meR9StFQm
VR6HVxITMnBLze1XkzQbz1jpDC2VGeZt1v1efaETpKw3u7GLn8ZDOgcYp1bl
+5Ac7QlHjuKwBtMlDizKYe8/TNC5TVZ8evQfpOC87tnYKdSNSppdE7ENOEvm
F1U5j8LAXiSNZ+wHtIK+XbN8cIoKUXNXC5u3US4buOwZysCDv5UO9EUgQaSb
lmrciRKpPAlsnq6uA5hONvsfvZWspvG2VR3I1cwIXemIGPfGfciMEtIj2qtb
JEU8a3NfTyejTF7RgK+IGqVj5L8b7Bvn0N2y+z75KucEEC7xSqNvKb/ZyRK2
hQO9H33ElnyoydNXA+92cllv08KOczmk0P9NyRRYyDglQCoLnT7Oq0XTYYyw
bq6+jLWjfO48nNGBHU6/60IArr+3lE49tBydMviTUenYekXSy/1YzSbR92w/
GAxZWe91xV1f6KSXB0iyrUzOETVm1jIaHWZs567wBrTKjRcDvmsL9YDl1Nmt
UcdeNQRnc0yYvzujdg4qWSxxu5BJ+X7oXSyvNl0N8YsbnHfj/fzFj786wg3g
FcCiS+Hc/97TYCU3KNbBn1CC6ORHG6ErJl8zdCXBllFzx6vBr2aZ9isDRI2T
YJ5zu2VCWNJGQJNeJ17xfa6MWhXnTM0whVZVVBKXZGlebLopURl+pKz16BoL
TrdNjo8VNbJma9+pIRye3/qDJB7Lv8mQM/r4ufHP8IsIonQC3xsgl07j0RQl
0p084F5r6m7ijGwCFRXRRQ6f2umJM97tzBCaf0hUH7e/J5fPcRI70tXHCuhp
t9o/3VGJgJSHI4gvMAIStRK8ej/IW8ecARnP+rWPWP8m/+41p0VLUxkhFAgy
GDQmw4/V1Fgyq7+nT88qHJceOCubF3Mzf4Zd3xfGLEBSUU2gspfc3RwRcMqT
kohBJpDOux6wYcPRAs8123769TJ5bUO6dhbZYV+wyIayoZwyng/4wjrupXYj
2AuE3WxA6GoNLuHcKCDl+yMHVEHUC+f6HSJtUnP9YMMEPnTXC9sWD7q9prB+
A8uuJ0iHkNAfGcEeDauHYz3qZi1+zMCC7kC0vvFQ/D+X9m9kBRavbVZ6tEiB
R1ZJ+5ISCpVlUluLRhiyeZPARcLBNAjPHegsmIymu+wIJBdjqSdL3yV/DlSP
7AzGQQ8KfeNgw73UYt7cOZVK26IcI86oFNrSQtfmIyBAoatAZEa366iC+8tg
bMJU9BkRnTdQPXfhkb4IX16XFzQh3mLQsBcUISVXJQTXZHCxyMzk7Y4TDYZE
HqK4E1m/llofYXjKaNKJnSQAtFyg2EgUzKh74w3npfNm9vjl7iFuf3MDmnkx
/j8zHUGAv6rsEVP5u+RS/rXXiRrAq14g9bNIKjyDrGSJyPvs/dZ0cp9UfxY2
DgWsQWIeostdq5PimR0iLozfrNmZoZApihYtxvw568nwoUcb1ZhHhy2lWLra
1qrAfYbznz1VliSZ+7txhTfcqZZPMcQVq42RG7PxCD16hTprfNPPKXFxu1bu
XaOp/RJcAeSx2x/Kv7prlLoQPskD3086ylfrSbDbS/ukm+FTY2GzvwJHj+Ag
cH7E1iRTYyWsyIf8ItfLtDN90ped+2cujceB+mvGgqneo3i1F2ts69TEHKyP
JvR6BQW6GnuckSHI80C6QGcBHWGS3EzSsnpJ8io2cQ9KZh2nuiKks+WR2/8t
9Lusfv+7S14x6baczxsxf+ZLXGNq/vyiCWDZ2u8b31egxRNNs3IwmLSSyAbp
7BD8/x0IJAMoee0Q0lMLhBXTAxi4DRGSjXhxzEVEutbosjIcWrpwSIfEcU/J
SCsFdLBRjZhLHVQeSIW6UaKlfhK6sIYyX+X6OS7bAwvBhU14rL2KlFv+nk8j
lvxapptLDZSHcikGcNgzgDzK7FtZ5ornXv810k9Olr0hmSjsTegIln2MdjkG
vsIm14aFswvswmSgs/B5QPbCFVFxRwRYdLSt1vHYhC+2PaU7efEZ8C0D60Wh
0YU9/D4pGfNtYNvi1JdM5+i4xehFsb7beHENzZsRBqxOyJGVYHi04EkwQJDx
Ok7YJb7Jht69hYNCdCwnL/oqgTKQfdB/dMss3+YVkZV3LNsDwRZ1n/sB1AbT
Orvo2Sbt57At+pTZawhTvOrZ2WFdt8bfaJhh13Q73lSSQXJ1gEiTOMrhojsn
aLehjDa/vgkfklk4d1Sd1Ern9XGv5F+c57Yx16TJUg0DhEiV1exU2ihj2b3i
aqXKWUKiHWgmt2DyHfTjl/0cKvee+uOLg4d9ykE4HMnThd5fj7m2Ago3vBIX
eCHXYz9OgeGksnhqiHOmUCfaZc2qKJ3YmesksAkCGBCkITD2S+ibJD5wbI1S
5Ogf/WlPzj6c4wx/O03vbPBFNFmZGY7LmzCz4fQkeaANGZMnD9KqM02KRLyt
8v11w2DT6XfjFPS37YGmaPWxgY02YJhFqY5F5qMW/0htaZBn5YvrfIdvMYkX
XG8QLkVlfQlLpCTn4noA254F/CDjrAnr4lkH/riNjwSD9SevVqRFkNA6Nihx
PAoutAXaNgzB9vujgZiIqHqcVyA3rMx+pR+c96VtOQeViWiW3L+Jzv8m6zc3
hQ3HLPMUXVVuryN/BUmlVMtUIF0jc2l4EwhDQVXua6szXNOJ12bhrAhz2+aw
W0RhJC5gbT/uvfL1qGiTKQx5rxWBldRu4NDZ38Y2Gg/7tMa20yQRLUlY6JK6
2cavc2ssSYplTYDu10WA2BmtjE9Z6hRlrwpb8grz3L4qBK4NLlDnxV2wZCjA
Q1QvVOjtjDJZ3SGyqRq1aMo76agZBh2xt6TBPr+hKKIr9bh1QABkFbuZ8qvl
i/5W+FkZVv0HxpKiw0vym7W4ay7Qq8VAAcRELsBQjiGlY+43yJ86QCehyQDF
LT1yuNhXYNXwxiwJL9K369U/Ruv4WnUto2kqaVIU/xNNp5nNgMMvUzs82kqe
bKhBtCCMbWifgqgXyGw3I7lda6Wuz4NYeRvMu1RgeY+DnyNPpB0xlfjua2Ps
R2huwqWbmKvbwYik3QAnmmp5/sS6ni7EOF2cV9OC90a0EL1dhz9C4sxfjrDj
5LC8vc9WrRQb0pdxVhSsuRLxGLXUoi2EMZlNkEpbH4I7zy7qyzsshUjt3Dx+
XmC5Ul1gH6NsCxO3pPC19jm6AZPzqtI9dnpMghwpSKbyCI2crp6Rq1AxPbHP
8TEmtwJ3owSSKWBssgCx68jYXeSqMakeX1KCnIq/n9KwO+lZkF7RvqQyzrOT
Elq9UQhpLkmCETdPyq6OGt59JKn2lYXW54lnnbsNjOPYZSM5om/EbEKKTqBG
5q2UMqpNcBbHd06FN0EpghVjUx3R363bDvJhFl3L1mzuEFis9lIMhvtHjhuk
WvYhXsxsqzBnhObkPvMW0XXuAX5H3I4uElaiMEV6IeZrzAxCKfD8OocTgT23
X50OoghyJ+GcVc4pYaBxAviHwHpsZJpD6D1cdJ6EX0OVvUj3vBkFDyh6MbXh
DlG8U0erVgMhC6S757LOSqOzXCZKUh9Hah0mI0PXJFCl9WfBFb/JOOhIfDhX
/A1WX+bC0k/ytGrrYerBwP4HRvX2xK4KarNA57rABFmv189i+6+3SborIvud
NS/9BHaYxhaUuzqH04zvnVTXEI3BjE8KHhwv424n0IJ4H1yajhCO8W8EMdJU
Nab1aPA4AN23Xo+fqrgRLTFwiu9bZTSqv66ZzPW9jU+V03z2v+NrSy4mFzVS
CuYy4xTuyD4lSSsGbgiBx2haDwzpD+8g0CPyp5Lmk4bbKm2b6pa4v8Yh61RF
oP5FTpD+xgctmdUDT5iKOG8a1rRDaCJLnIx+XAAIl7KMiwGNEnqkLcsFssQp
Pd1wgbhWL23EMnQ66fznm/QXcbkaWFWR1wAanFkKCimSWEWZU5V6norLmVZP
dpWP2AVvTF4x6AONoRFhmRi6YAR3Q4HY5y4heTuWJPVAgEmCt/trIsYPx5Gz
gM69PPN5EARjSZn0EIUegL6KAO3oWF4GHKGh4h7m9IdbuwqUDV5Z55zLjiC2
LZqTS4VVCKEtNp3fPL0JJU6btIpFtzJTpeVky/1P2+h01TgBMR7Ob3V7ELOU
MjYFXtIZI/saQQFo9L4qQ6pMIGrAhxIgNdsb0vHG4zolK/sgBIo/u35uR7/O
V5BPY14+RTZ7JA57t+aVOMWAq8/6QJKO3urBknDmv3bUAstM7Fwx2bNQaKPp
gBvGlRy/UnfoNn1JcWhYRNoBY1zPyrrwbxcpCNKkgczoBZosJPXO0GiIZgZp
Tz/b3zbxYS8fwm5rG3SMPsG38Fqu0Q1jfQvxkSSzjXn19NmCbGYm7lHjr7l3
XTmrI4RySWJxdhT2UrZpEvpt7LFqOzFDvPXTiLRTdtRiD/tH/sAvzoFj6cqw
rK2u1ZwHk1hWVBBHp9zECZSugP/XhUj010kDC1U0VJSzZyDBAoj7a6aYtc4Y
ULR/akEtkQ4cnDfk15HeK449YDXmATnnGQGx+trWPbsj04fDpPOqYIYrdIiK
0J2BBs/bs7sHFFACUwL8FMCRhuYmhxfUK3tFvf5zj9bfLMEHEg3GPqb87c80
AMz6g895Qzkv4eNjQgBqBc2DYMSzcFbnBuovfY5wceFOw/yUGrxWIT4u11cR
bh/pkiLrnF/PScqEWnq6AWQHpiGyYl83uw93nh5ORsa0uIxoHmxjG8R+7eBt
TsFI36+ZZLpjuqFaf+VsfEyQpWr0LSUvaJmGl4DUS19PImm15qucJQhH0bzN
ac385+n72sj7nUiJB2wPvyoVYMXsZiDensMvGZE8b0nuMGytHwMEVgZOKAt9
QpKy2mCB+X+U2bLED27UMvIeyjOJ18YczxwUXXyj5+j6kLoE2DvsW2t6nuC7
TZyIhVnGll8wkjwJYa0OtCEk41Jtxj8B1lb2jna3tih7pdqOH6kKhsOEBq5v
altDv35C7Jo5bdeQopYQx4qJ7h2WkzLoSVXOm+zEa0vChrD3brv4um6Qs/Wz
VNjh3yWG9wo1zas5d7BoMn7RugQzUwaGBqykj+LIrGGlbHDAGyDMJriYmQaH
qrW+oSv8F9VRzRVambonwfP+tKVNlU8mx+YK7iFrQL6I2eH/0Yyp+HFxRAEl
8C7PNfFE4yIuX7yJ0okpeoSqyuCtnZ7jBeAqY6tfzm9EgnvOI/kQupWYnInG
nFYu4ZISsD/5ik1dUWXVN6KF1gKtLZkq1lQdAEqXA0z843d1ec39/BOxXedo
oVRB7yZ3i9xRaiZrQW0pXrPaBleBy3qyUsTgz185Kl9ZTvCXlpiFGrTi/iH5
IMbLLgbrfzANPWS2Kz+gA6ITRA6YHAu4CcrB0vFCj1/vPALc0i+1dp3mYbKd
qGZu/70CsYZgHbGwJ2BtZmsYMaSWdpIc0024G7liCWcqXkF3nxoPmyiSRL2V
xrJeKvPRGQgXRCwNvIyeZdTGOTJO+qQjgXaASExURmB5pUASmoZaGk4hVjFD
k+qrlrRdgnjxuxj7ysx5zizVreRXGxEHMSXBigsu6UdC07G7es+YjvPRpGDK
BBB4jthp+hR6tlueWhiueLkoCaVHZCSGKAbqOBD2c1soudAlfprB/ebZ7QYs
yb7XFcoYKhSMI3XiOOViVcwK1kvxZEnDBghRxhzCfiwuhYHqgE8R3EyiJTa1
ksxSqen+/TX3EVviPn5+kP5VBQF2d65xI8DVsPZVizk7/R8L+9IQoix6LjWk
7u9NTQZhbh6YX4sMyMYIpLnsbeY4ZaaxuOu1ke2gutZg+3jevY+zGiskjyVZ
2XHf4OA9JVHHF9dwTIy4A7GuQ/XAkltMHxFdkGh18rMlzfJo713gywl0F/x3
HY6wXBFj1EWzZ4nOiIMK3N/RH7w59A0253C6m4MumH/6q98xspw+j2m+JTpB
Fm9XmWZ5nZz7yr15qgs3CqahTyrD3i4p7zKnvHjsJ/5Yz0XI9yriRxE9y3Cc
z2fgCQoAjbi9BpSZP91ZXNOa+IKvUSQPRr8GVdNu2630rXmTkdw5l1q/9amo
SqcWoFSzFSYGjkZdY2Q6jwi9X0JZ6u7V0UtuGy/8MMmGRl3ofEpjpZLWkzyX
2VUpsPeWKznZ4+7e5LFkTtpHidVrzzUleSzOkEWOyvtYBEmqrzOUwwyGtsfj
YRbmk7Iyu2j0Vf6roCdqoumElZEov3mhoclN+SKhHEdFkeKTkGX9s8CCcGuG
t01wrXhXJX+Kj8sr8ctDFsO3Y8OoMicPZWqxfjBt6YhRz+QIsc6SCdd2PqDH
hwfhCOA16n5d144Z/2G+GhHx6cijmd62d5lf20m9oLA5Vp7fNVvyff4M9qaC
OvqHh4+Ew8+XdNknB1RHSOm89f65lJgcQOYaYgwvCx4nFjsuQB+aJIo4bhsy
SCoKfhQpQB2pM5VBJccRGU6mia5s62GOfijCs+lvEUC6s+X2l20njhVvQR8i
Gu+YyBQRBpqi8IYFwCR2rpsx8JUfXJrODr60E4frNrL+7o3ZY11cgnUYegMz
Aw+B4k4SQg4Z6EwQvy0HfXshccA/9nnAEDy1A70uN8laBuVpAyhN2EBuV21A
SQlp8afPybHFw/00UY/CIlCE3Yr2/Y8Rj//OsVau9kw5DNx3laD6Tg6jkOno
d/qGGuj6hFtDEzuuJfpsPG1ZVNQodFZtAW52l8VCzAdPEywjpPKipDtPXhs4
fTKADLmh1smO6KXJWxuaP9nksifmK86TE7qfjOVjuBbOoIMqYtixNYmrjv0x
t4p6+qaokBzTQhf66Hz4h4QrtqHMO8jKJSkcqFm56ei83/wN6AfPeSSiIzIw
PCua7J+CZqTTIS619j+CCbBcz/N0he+lNEgYJdaKk7iVnP8JWAaV99kbcM9m
8zFUCrjKAgPmbVY6A7m/UdCKFDbJx659Zr4CnVkKAbPFDaHS7VlFn39QVDMl
Mb9YpZBL81fVNrkXLag6BbsBa4cXdHDvccJVCojxHRdiET5MFqYSYrlhAEY5
qFD4uAoHFxTk3e3Cl/sGc2QCAi7IZxog6KRozPEKiswe6xpRa4IHoy5AwxKR
bowoWyFi8uGhhXidG908Z1fXoT66bq7nn3Bt8qaRAPsfEfMUApwMJ809p2qU
uNxjdhY+bDv80fmE7pmjiqwioJI5x5AsKqLZqAHPmA6jBAWbC4SypbgbLi8B
e8993kCLb+aSrZ5hcKxrt07NwSfdkESi4q0DkpdB8kwbLcWrqZqp/D12Pm3/
4/1nrJ83g+a8e3R8i+Xvncx57Bcs++fZT+QgxYJcQILT7e3OXjXItTcH9/WT
EtB8Yc/5t+3eBu6JCBL5TeLGQ1iCVqitejQKuUsK2vTE9D5FvyNjiNfDLz2p
7xGXRZiMNbAePKS/IeAk/i4yUwzUKsWx2QAEVEzQ7TBtEaVF1fRBufKfbyts
dTmaNn0Zub5alSdFS8boag/ESYEOjGHHA4XEbHUcVlYObVO83bygsXqD67KY
Au0lRfg5PncF0HKGP45ilSWrBa/FctyHQEPDJSUTPB+zDpUUKYEqfijA1cxi
93NVqESrUZ0Sp0bXMlz/KfHENSr48DguOTXGwSXC0kfGcVY+yCSc0LXdoDYX
KBWJvoCE+2DdnSsSVr3CVrzOg1LfMj/Gro7x0A2o4eytZhYyzRdtfQaJ1P+d
gvliWXg/B1V/E/YFfZvODJCEitL++jdTgrvqTMagEf2a957bDiht5+EXKIt2
8rHWjdITS+m//OoBbChCDpcl5dozsEKN5QwAgLpNw4iB/XAMHXx6/mIlm2SU
uWBm/DfgSgQNhhNC/HAjap8WoMo/7vOI7pIvMZ8UJ3aL/oSjiquEBliKjFwc
GMVjp1xNEbm0BDS1JdRZgrbVIXcQ5EF/gQUpJ1gJfxpldXn6iFG5sf8wCjQF
Iy3wHg23hOTqxU3iz1ELBn9aWScW9rkEHN9VLCt/ySjEj17ue700TFNy2Il7
ohp2bRVXQEX+lEqEc5D8kSAdcEX9ubOW+hu812qsBBRCcoIwbWp657woOCbq
qIl06661TsaY1Tx11beavE+WUKAueZz6pK4GjQYR6A8pqhABT65A+mVU8P7Z
VeeSJirqu089sYyvSy6kAIKqBJFMqGj+e2VML/jlVIPX/JmzZDuTWizMFFFz
T+x9v/GotpMb194pfPCFPNgsyBsJzS3rvDlggNhzW4CStarVZ3QsrGnCcfRF
MEVU65ZJ0rwr14jkKGKepdxYWx8NJ68QgKYVoA2HDXLS6GnIkFOf8Deu54Sc
Qfmn4sc6PDhTBE5MnVO5rPRDRLjThzQy/RQVE9Igr4e6ejnkjcqMgaSrcElj
TGZK7XkH+BaeyPjYCpC2bN/BF2XJ90EhTTWtXmeDQXRu977wLy4kGKi8qQmR
GRzFT7hW+Ml3zFZs5NFIO2l+X0J3dNdEKODg9cglrNegsZw6gx1dWVfRNWLI
YY9pd7v+ETvYv9GfuP2X4vXvWq0ou1rensuwRqAcSJ5fsAmt47fCB1jUsFTk
vlbZ+m0mdixggiZUlTcSznAuuJBbgN60SQa18tuP7AeDyv8x8sWQjuOkwhs3
G1f0snSrWstn92RoSQhaPDo2FxtzlYIXR6fZ2nxNsD7NcZNIckIZ4j7LJsbJ
d8T632rE85JzI4385686YYULfrNYx9tnccb9x2ZzyPwtlb8hq97aNVEZtzlE
0Z7B6mGZhQhgw13ZOF94+00citENoVpaivZRe9jx6asSxh7tOYsUQys0l2ZF
crHQJ4x3/WreDH3IDD715iVJ6PtAnQaFzDkdSwBPMkTL0RsyD/R2VheKBdJW
KRVZe9X2kv0u4t8DTXjWCXzsDxhL0Rt58ZrgwtRIGXV+6gebTuuk6bAE/eei
0D99gcmhAxH9SOD/W2hzyfDnqXvCoJB7z/y7iZvcYuPulq45I/gu5d4uTtsr
VkOe8FWykHf6bA3/vptmcu3FI3mcUKDcZd8BdAs+S4RGX6jrsiacGsVyZ8wX
aFDZ369VqeH/02hx5Pg/X4J3VNLIyzkw9baKkFf7FoKbInJ0PmfJEBuCGM1+
qM+wR19qstukied90R6BMh/NoOmviqTOav107V9+FL9cxVMEidK97BcYvQ+7
QNfEWev5LyUnpvNj6jT9Mj9/MbQON86Lmz+6e3HmqCMdTK6JZoyb0A3BY6XK
QTs/tRIKxBYFsbiiF7tWxqaNwnh4hJas7vXGF7wKn66LqLeF6GDAkbg8OIGV
zSoZ4v4vDqkzjbbw684hB/+nHFxc+xe1mBCdpmD1EIgd8K5tRDH5IijIrpSO
npVcK6a8/5/E2tV9N+t7bmCBrDupD/yy9Qy3YlFnssyDA61k/XVDTZ1swSTX
0xIBXVB1UVLTOkCfm2ix+EPUrWRB9GMRYBZnqgos6bsTilDaTzEo7PP1jarN
PX/Y0jKBkAiEUlHjR4Lnc4ptuf+TbDE15QevUTzZj0jyQj4JlSe7zAcM5Jw8
dKOKMQghQwDq+u/gn5Qw03BlrH4ZW0IQWEge1j2GeVF2NGgvCW9rqRytC7vf
W5G/tCXVSTgoixljcPQQ4oziP/wspTjqVhhvxNG3VpOt8PvJkMhXHJneVuX1
CkinRtUyUJkcuQaOfheKf5oR7kerQMF70gGb+X6sxrKfKmQ8gQlqAMTCRRFT
vkGZGCvE2jgz/xDtTK6LFOJ3zxdH/tggGS29C8Qf//d6vW6fv2iGzAVG2z3K
hbjnFQ2Ac/qiwRKDGf6XAC4mMxfGJ2/b+gya1ULfVTfpoqgq9QO2e4CzkrTS
3VQomNj7esvU23ionASXTG4o66jde7NkhxwJxz+L1nROGjB8YGyqfyDQPb4V
pGVQyQnHwFUF/N/MwinoWZlwTzKK3qw/LE5oQ0q7D+uFzopTYT9qFjvuaTFd
D8NjiO8R2Ly0oY46orPKWMo6OkjioVRGwfyE2kl3ryD8OTZga7BUukPAj0dH
6p6XSvTQtCJZt96tV21pZnB4NU8MFZZKDTYp/J2sxOw9UEKk6fYj1Xhavp7X
beibPrYbONqo4lAtKww7O8P3jNoLMtDihgI2b5wrghfftTG9Ud0rGqCUhMay
5+z7OuXf+F5AWNRqJWZaqnoLYiTYH4RnRRi6lGuxdTLAlyWr/ejspqu+BzVU
VPgVNhThn28JrsPklv3pG352eI+Wnrng6iTOKqGk9WBXvu1QVe9PQ43R86tS
K6SYTlyFrZ0ulGdVxTa5BcD4WbqhLq/MwT/wol/DpgwYlR57o7gvFLFOB2T7
ImVfJBbTM8l+JgtoCLd//bNHMLfC9jkvuIx7mDs5YWOwgNVjn6WPJQf16Bxr
yYpLcSpyjAGR01fv5PFs33L72VgxLGEpObcfyJ8ccKJ5ZneBm6MGZEWg8BET
Giqo22fjygZH4QOmSReeP9Zwlv52uw0dYd6LLokW/Dlw4unt+r+ZU4Tf4gE+
7v1wfo0rzUhmdOnpWfkLkxA+6hJgvtnFJ4pJKzGiNmDIfozrz/S6uwStp+w5
hKaW4Cw1qUlozDGAj0oB+8a0LtxoMX+q8oEkCg1nXiR7MuY26AP+UzPZI5b8
xvHqifK6AMl8tMIcNw2B1GTtqaOzxWqlcdpIoPkGwX2Vsb15JBPsq22krq3O
HofKobyEfukj3piQ/mXH/E0rfMbc+OWlQbrhEQtDaCNAVAyy4k/SSLylM0H+
KEAxYs4VHq8vJ8bGb5uSyXMzk5foZKBDyZpvqhGDnQnddB75ne1i5YDsoZHx
+XHgZEw/5pCUBezfG2QOrECyzF+nVJnSuW9ekHnPdFrTMMAIv7Bb8UHQ4ysI
2QRBRrqAdq3Y6QjBId6uvdMhBfnZmcwGwqY4goAQfG0hxvLLKCPZevf75/7k
7/yC/Ung8s3ua65TPfse0bstZVQ63+vSLQ2ToLH0tOBc6O7GNvvwLJiL1uvL
yY8mKFh2I9Cf6gw1ejeWoTbCR8A00A1z9FOenc3C0c4fxpr+kUPjo1cXU68h
IWygGirbSdF/pev9pt0/jrm0ekYu2H1dcaBJLNYcVNK/cvDl11Dd7tUULP+p
hW9smJtX4H52zEY716utlXWuU6/tVFBDeZR+XmKzk6VSTpQHTLD8SCKVUYpU
tUXKoP+2lNJjv+YtuD5Y8ue79J4qYXbraKnlMwVcuwCk87frx+lZPeL/OZEA
W9EAl+8x2lvNRf53qZIbeREro0AsJpsf0LeiIl8VEi/k0I1t59uKSdITmriW
Rk1Ynep0HFlVaCtydoORi5FaxNqRiFzvhzaYpgg1norCBAhPrrl2egtv6u7K
Rdttr+jZNkBXrPlNbH6KTKv6rDivmdTBdknbBa//fKqLMgGgpavwk7JBiaq7
DQI10bQyQfhUUmV/CPkw0Borygv7aCMA2go8mGskUdGxShd7/yu11IdG+WGD
sXQR2B0X52tA1WO68h2m6Pp8xTaOo2NL105Mjb4iCUcojSDZNfupU446oKiP
FaTPKnh6tJTQtCBBlnpductmeX0rIh4ITBgOK4Bxlfc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpei8b+64qz5xPa8wlrNzfgr8IJIvN/ooJepI/llP/1H41EFZzAqKnNINmHsisUFkZS18evdf2U249FgRN48Z8uwnEnY42rwIr2ZKZYBNI26yAHBvtfqBF/vMuS5WVpacvS5NTwsMj4HoIGdpzfXn7oGZOoC+d4NGsudTzr/tn/pMfhRPGoLFDecDdUFa5DF47zBlwDD/P8z0bXQ3gf9W0oFAhXVhahk9ThNz2m09jp6ST0VYeSyFU+XKHhMNXTBJls2D6KUCfIaGi2tSiYn1X0M8U/7A5DNZ2Uh7QOeoLf6CqU+aF73y25AXR+Wh3Cpxd9cAqxH8wbmcTT3x4jXtahqEDXrmksoh3ybGtjiZ55LXTvCaiq6uYxK4jRGJjOG2uAibDlq+fio2VKZMd50jWI95niDar1KDUpae4Dvq3NVtuPeMsKoMZdVH7Y+5gD7GNvjLLMKOWCJLxaaGRk9oErLpPQLBU8d3MMCVhw5DhuGQF4LL2i2GMnwD/edothiwH6EAYIIJ+uIoVQaIsCDkRLphvYo5hCJMU352/lkKUWM6VCwFMtDuTXjG9yAJieAHfhWFJmKlZv6xhaDUCKxBlN1s0FwhwaOLhFc6Xl9qJRdBchq508ugZtxYTMJGo/7ocYUxQltSkevK/thQig9fzJ/iGkMi0af1+pGQcynGzkLXFSwluhah4MqWWmVxHHq6Jfjc6uhxrnRP1hgWVnHPs+wxL8zelQf52epDxT9Mu8zqoZd3/jS98qZAZPpkLHzrqA6XuCSNClBu+wP8+m6MKu41"
`endif