// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tVb2UH0lljZ+idUJQdVqAeQml44Dg2eAatSnabVKzYnVNfgZTuO5/F2Sevct
HsCWtRxCvCIpKPBeALrpc4ioTRtbcssFJ+BR2Wi4VYlbWwPUqRUe+3v5cMWd
OmgFmaXum3HlyNeuceRU+qKA27mjyNCYG5GkBxlDl8ZiMMMGonqRwsFQI/jV
H47v9AFORsEOIoIJc6JGZtLzaP5MeaA8eS55QMrPB+mXz5PXYJ1ENf4A4stx
8kbgO7lzaw3ygtbr34HmpyeCwoM/Slu8/Rxn+ebMwdEiFl7GlQn/jAfd4v8G
ms/uG2AL1CqZtcUU6hnvoGOslfkHiUI+/fsysKv3Mw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GNgRHhQWT6CDhcPS0NUVcejg9k+kD564veIZg+VIuEbTgVwB5apvhCAljCoo
eAYnzCVUDFwVdgLtnXi3xBFH/ccaENeie1rkxBftDj4RzY5ADbq/oeodAXIB
2B2wa0O106ambhrdOt9bxWppKmOI7V6/aB//5+RQGRX6yn8bBpXG6bnKSSl5
UoCqFjy0GLFn4pPNMbYaZNQEpTzfsq90n3XIJ1qkKmaqChTa01lkLDmOZdr8
zAhvMQMP3TxnVpudvcNoFUbT7CaTI/WgbvBaa510dcOHM2yMt5qSL+Xnk2h6
+MsiKi+tpbDY2wdKbDHaupsTkzj86cNZ56mhU/I6Sw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hI5ZOCuZ5BJo95jzblzTyBjPbIEM07pSAAxVT4NdedlXhNyqjlKYiJvyefC2
xKwg8hiSAVgq49bhQbKSU8jrPnhyZ84KfdiB7m/rYQBEwlMn1TWGjNwYOnPM
3G/VxDAlU9coo4KoNKJCLOiUtpCI0nPlz6mXsyqbUurzpFbrEFZXFJua299M
WmB42XqHvty2AAOr86VCymi1i/fmysVPgVewQpQTtWr5fLi1F1RpbzobD8Kn
VeB+Qtto6HIVMwubD7MHqoNomBZaQiVl24+zfNCrUKHdE5yne98SG/AGWPgX
cCtZciE+bEchAM7diN/11NErS9dJxxKjH13rS1s3Aw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Io0Yiro8DpbbkYPitKJ+DF53DyYE3885n7upbhXrSu87BPMBWz8gQB/95PYc
mdTBOW7SPzXaTvg1L7lqOpDQzmCMPDQpU2L0ZSGMpXSx5gyEtQqKWlK/MV+8
sqXDevB6PK8vfuwU8rU1FOdju6HDPtunhLO1c2jsxcaub/jmIc67OOO1qDax
bOua2z9wMDG+n0bJJh/AFnFgfUPg3QD/2dM8PlkFY2YTqeg24dq8QX1v4DaX
e+bEi3gDPllHfbvzHi5rfyYErPMhaEQQcoBtK+2PYtV+HalrqLvQYWmf3m9y
IBmw3fIrmJ4tW3JteqgC0PgnC2C1c5p3QIYlQtWmXw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ct5XiDuBf1mmLRnFa6t5F6xwvK1vxVld0TmyRPk03+CD/JBm7AzPHb0azkLR
9BqVOCNAi4ezAVaxevxAI3uDOg47f11TTbltZ8ClPLvt9ucqx2hiHQCPHsga
wFMriRAE/9PZBQbjqnhxpAr4JpR6hetRFds6JhWzG8sJ+pWSbhg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
g6e1AERhGe/A7JoBuB/sYT8dbw8JIXAr86j6AuKI4i4O+Llx5CNEIordiWRi
RI+tRSJzcj5vB9o8MRgAd3jMaGYQpW2fRSIx/+kc7IJTkKBqQMEYzkr9DkZN
DXa+ye2fO3uOQJ47Eh5Bj75hQR6TZfJy0l01Pwu9eL/q/M+5SQH/YbsjFl7c
ILomhozlpl/RvRE9SrkNSVXLKt8kH797Yu+K/oJC+7Oj6PJ0UL+udntinN9O
CrJ/2UbjmaMQaQfJs7CxwRifUnzxlRYcYBHLBk1iKNHYSRufaqsXcS+iaJdM
aqzAibJxU0AOGhzpMNQDFmrMjD2zWmLebHoMxFBKrTsIh6i+2EUHf6cVV/no
j21kCBGQuhW157GtudPhkyStiIezJjfDXm2pDiDEcCjMZF5BXtp25Yeo5NOP
7bT7lQriNHDw079aqAQdcQF2xp8RPaJ85+VsXBVr3higZtgTtNB2d7hp/8vg
+l5leulVMIDpPAtjLFQn3OqCqDd/wsWh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Tuai0PRSA9GG7poX3mXyq9OXpeUX7G3+VCZ7fCtTUH73a+DoenkxZz03eWlq
i4Fm5mso5U1zwpxe1cLIPTdWlO7ezq8945nPaG/KKnTae99qtNwDCrqYjVSM
qY5V4Ur4bWWTzAXzDUxZ+tj7dull/J+q7EOy0b/TkvV7R8BgOtM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MqTYgc9Q0/FxlLorUJq0hmVoAu5Y9SEyF5UDM641KQ4umKPox8lLeXkTy1hp
zHhyl3pvIEu4TBvgik7RotskUDg1ExH050noetQgckiO/Yj5XhFrw8OierAy
BZ+9TmE2lWsdVy36yc7ushCic76bVDG/42X0NSNwxtf/JffXxeU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 77056)
`pragma protect data_block
Y/SNd+r7SzkffJItcyHC0r+vLk4I6QmjeF9x0Gz+z5FWUUIFLBPukNb1rC1L
0vrmIXIsUdwzWsYXphkvQivbr22TMCP/3VheYb/Z0xmp0ZKwUmNP/oABAM2d
jC0MYxxOM1bh0NVPnLvklF4QyZMmnWYpnzkhboOdqLJP8fWh6QhUxooi4Y4Q
jZFbcWo9wUZw6+gJF/Z8o2+cWWK4kc5UppeAyEczcck9MYP5tRQtGi0Nm7eD
paLwZ8msY6ComULjoplD7UFQdjmiCFz6dLGvMZqs4ujWkHB/SZnWGhuHyRrL
fpexEzVTB7WtAL3jjyEOEo0rKwctqcGJ7ruyclZWD3hF6iiKNV8dOSD1/fj4
DsMTBUYc8OlzDu1gX5egzojIxH6OsvSv3Bz/BubvrYu0Zd0NXlz8Kb3G8UyT
/6jVlJ73AqGgMewQLd3AayqMGK6A+kOgNEyqfl+j+rwoxjPUxOhaHHBK5ACw
QNifKQ414hQxZJ9o6bdPhx4+Nl7uSC9oF+//6dSb+ilOwhJEZWPYzADh2fGA
wzEzKlg8fSIAvrhSCnQHCfrUW6zyUAnVRYqPFp6su7Yn1SWKXdV+9zWYZG+Z
AoCdk2WP+H9w+7G4Bi0cX/SEJSz86P+BJqCF87mONO3o7dfHYkiIBgn2BsFM
jyEDZ18vBu9dok7HuiHx80WqTw7TKpiWWcnsryLlS2ImXS4IkOGhfTMlYy5u
Vjn9IwbbzDFToFHpihqvW/RH4wpsh2z9NDxE1hf4ea7U9dN7N5YfamxaBCYx
ypyx38Z2SfjP5SjPG/CnPVZfAB6Ql+Xnrz7QUxCT9SbyqpnS8hW16pc3nXV5
ekK1+bNql4B27XW097VULK8mCFKbztETu3h8EKGQmtAckcp6ZcyP86zQPr0D
TwPE/1vWFOxbnWAb0j+v6bhhCr2Pr+hz4/6kdLi59+22MHodTrwXHigOOhQ3
s/XT1Aqyhfjru9QRs/N4KV2PEt05Kxw56WW35mEqbTOdykJyTgR+Jy5M2/Xr
4LE8tUQoJ3LyAieagO/vNpWX62OBydQngjLce0hfwXvRKuB6BbTo5vBi0fed
wHml8C6OnpuwHKJ/tweokmrmwJ1dR+WmZIWltdEigJZ/tKGy8vc6oa1VTgzx
3AWEyNx5fMt8ADWKInh1JFnDbLdft6snhlFdHih9OFb/7c/AO1lTlk/snVNl
CvbGQgbQ/C6t1CuTrH/aQtZ0JcpjVMfofvxJOH5KLgoJhr1IOYLNT2LHITWD
GIFHwAW1FzNPs6PfM0fMXFI65AtN5EIzg6XBnCnKulpdrvZIYsBjf0+MrFVR
4F7o5PqC6NPv5bTvBub1qPYcIOCGSXPERBZ3Y0zL8Z8OqKN8D+iifgC4ZxA5
Yx5NEFpeUZIWcfr+F2vXeVSJMbvmTcvyqsAdoycS2CoPICmWFulRxI1OxD4m
mjyE1LkmE70P/gaHdqG/MNHLfxogUlFn/RahViaeDeOPBrqv5+w19vuuaDXt
DW+vCirTWFwtkTQwx4ChzLYHvUW/30vJPL0bedWYm16uvgCpTooVvBYyXrwi
PWnNY/PdyqhVnyjz0a8tCJsmTFUkdhRYtYe8HOJOwoEltOf3F5JRGMnjevTK
2mhY0+0UEMtXrqq4D0/O0b+Gh/Jjj59LlQ2FdvulcxUkRF5xX3A/hp/FYmtK
RcwIwZriW9QJrezW11h7rSfJISnJ7Z9n3MB5wYJSc08K5LO2xcFLHxqkIS4y
deoMKLxymNUIM+Y+QszmJrEmFzkrNBYCbexyYx8w26toRHd3/N9MSAXgR/zU
r4kXaV/MZlQsMJPpBJ378q2f9s9mwjYY4qS10SQLPf5hg4NDGYC3UhP2a/+P
oJ9d+BoC43vBgBWfUQ97vY6eMo1zEPEM4prh/aJFhz3gdXSvzsgX9hixQ10s
7zgW5KBCevLWGREhjdqyI95OGER/8Yxedq66vqlWrl5xlrkTgsDauc8YZpg0
d6EX3E/ha4nQZ42d/vyXjzjuKQNMP44gqhjlIs+v4w32NRnlC0N8h5ebOH5M
xqaJ0uLBWzQZ/ZSremP1IlFkWiZ3DYR/KF3FOEXTITuA4N8y/Av+k5/SKdJe
nT2E2CcvsxkyCqJEaaZ2M6Sghgz1ItwvWtKeuGGMN9LD+8ymhM8He7Ply5d9
Ehtf24NAQ4E/1QdTTSxUD4hZ9RJ1PdWRYgiZlWsz929eHYFlv1n4lk+0Ww5E
8MYx+OeYsRU3jX+ZOQtOKFsJCMI5b72MeBz1/3hrjHLc5ni7tHyJzWOB0Dnr
2w7bQj+mezwjbOSgQY40G7QUHQByU0YpyonnnjOhJ7Y4BPl04az/AGa7Mkz/
IOoUvsXKD+65mKBiQCZCcTBXl4xlekfrkDD6i0sKjykscS8T+zmpXv9LSKpy
J2qiJerdeIWMkoXNWsGUycm6A2FmFBL7eK3VqLcOdvm5mwbCNEf+a/1aHGsE
+u+sqDDFjDcdaeV3o98WrCVt73/R5jPjID9uOaRRIp9H8alDEbZ1vCuVk1Gi
v/fIP3rbHDeVZOViOAYAbG8+K651Dk7L/4Kr0CggDhO32p94BPUqwyN2nTG3
ftAMAlVqeRt8c2bjbVF5riS0KS6QJ3FV0pVRalQkmmxcuECemEy+WJMT/Bev
bAjsGLeSZfJjWhk/In4hfR42eIaD+j7VbpqMF1nbllwPB8cPf79MvADF0nH2
7dJ/QgRZ8iXFptGRyhyJpmE+JJiELcbnQF6FpgsPVG7AehzuYWJiMuMU+kq+
y6omZF3FOWzSYl1fcAUF3j6HTWveAcYPSrahAo0XQ9sRcHjqCcS1F7PI3vvc
4Q5BRA3Gf8+VC3oNEL/25EsPs12jCB5vAZtFTDRb+lVS6yG1qGDnoQZOdtf4
k3L4P2GTcgnLM8fCT3NtLocnwNKkTHoAcbKc8icuDjd/xxcb0bp2Vpp6mPRz
AKN2Xs3wEHmvkkjADF3AixBJlNtkwUtsFHOeRgjThCbV6H/JoLm/KYAdvgKn
yUqZcWPZ1Nbk6ml7I/Np0OdATTQYFsesnwOAudTF+4V6lq8/oecy6tjilfYr
UrUtznbxTiLj80ST6k+D4ZDYDjNXMGzjGqn1K9JNf/QMbZvBUxm/YOrOgY3A
uuo/6a5ppYnDK97NDavesg2H6EP3rixZe+vosN6XjrM7tbTT+nqkZYWLMOCR
2ReaHTraCH6fMRywuJW6GcQ+wRDwbBev9sAJSC4pElTo2kwv/G6d87oAuqpF
GRty5lkyV4LOg/5IgysvQ7OaSJk5mkQoDaz9Jh07HIpMMExXuReAhVaptqha
uPstlozz+o76jBsnMdyn7XaBOY1mRrC2+d5SMaGY6dTBWIMDSKgco//EhjDD
z11zR01MokyMu+etT2Xh+CFWu32Oi/nW8KnXeqXUTyfn3DRvyXBAC2rNK8nm
NzosZSTV1//K1h8eZpLm6bFQrvOkC1QQ3YXwAjVmwANIP/5Pkah7R3ieO2ek
2KktZMreyGVtdWoejJ4GqlxlFV8SBldaxcnBz6wHrsTIhEdqEVi0VuXUbv/Z
KE91D3M5GkdJiDjroCbHhnIkVNtLON0G89wGuDaH0Yj68aZHzhGruu1XwN30
z3it83uHS3+Y22Cg44Q0xF3c6KfH8psbeFuP7/zH5g2oQ3wxWC9XJFQFmppl
s2tfP1b4QfpezmF46jY3ZiwldPpXyrtrSeFG9e7N1SKOVeZvDoT2zQSXZGzU
3o8AwgRF2bqLZBy7XaJLldgIxmXhvBXe2hKIUxvhKLX4Ghfgy0+A4Ur37NfU
RyjZLNO3KH8rVFcXX/oQLIlpO/yj13mDCxNf3NHtx17eyVxYui6kK9pT7KCs
vDHPPBTyNxXZNd2xO9VwbVRoVqiKWsOksBDAT1dGMS647cjR39jyl1Elnaki
UCzFqMXVRgzzr798/ByzPuxBlkGDTyA9o8qeDA/ghTsWYLAa8hKzOnvKw45H
mXEr2uAvC539aINg3tsb3wW+h6YwHfsmsPI0pWXd+inGxQSiv7bXtxL42tJp
Cc8CvG/umtnT4zVj8X5LP+xZ0c+LYhXtmMkGdCLUGpT6AqlF/MIMVwQqKlQJ
yTQlPF+ED08/xpc6VDQ0NebezcKKUkTAXVOyu/45VK0t6izCo4mZ7GxMY3RR
t9TTTadtS5e52WifE4BCWSnj797QZJGO+UB5iE0W3xhfFOPv//V3FI01KgBD
xEmygSBRqq7oXB/dwNspn092dJ3u2Y0A4YO0Ntfb74s1JbFNef84urzLU5Yu
fMA/cfXHqbt5GQVhySuPFSoSit4ji31DBenuUsfXFNOdyruMgqXMPyJHpeNQ
vyIF2DtXievUsek89y6ItNvH68BR6i6YQKD1JUWCPcTsdXEOjMbt+/KusRR4
VTrBzPCUx9iJ+xBzkOiUTQirlJDHfj+yAww4DLgJ+jMHl6JQAAeluH2PXkBW
/hq/9AIRf2tGztQ3KBRSbO7T81KZa64OjSKmTza4vtCgpgPRn43ZcdqHlfVV
scI5PwSE/X62Cwo6kmPFydKRfRMbBj/8c25OQLZ/R0IYDVdXbR7dc2V39OAO
sXp0RIN7JjEvLOrsL2Id7i5iRxBE1QIJOk8Z4P+Z1mCPPxNf4jq/hweo9HMC
M/tsv2Jzs2a1RVPx4lHSqz80PURMdgxp2upxj6ix65VCt6VTyZiiRVkrZbPK
Iq2vHYv3PA7DEuq74eqejebf3JDRWKc+YoHNX8pJEtHODsiOTGLUVPnPkChQ
DKdkdCTji7pAJMuZ1Z2EUbO4BkRSM35Axry9yQu0MR1tEyg92s3i/bcLCOsh
t984OuNlwLMXJ1J8VsbEuz9qtbHu1mEWG9gFtHjiKv9df8SIdC9KnMkUo5bP
VH9r9xK30T+FkwPRbzZu43RaUjAkJuT/Y1WyBhLCL+tEzTqOWgUWlZ1Ogf43
/IdGb9jCysoVdMYCJ6SwhU8MbAt9t5QGE3ltwNU1AuQ6sO2+WiSx16QG4HJv
90svQDRb5P6r1L4a5SaDi6eOlrgZoUFtQoFjvSDjtIV5vGTdl0l4o9an2XNJ
5IBGbbbiWdc8kDPDsO8r8BISthfUsGrwJPdz20hxHyiFN4YkiNehqXyRguQW
V3JL4MuuPhxOw8M3AOdytQC5kE6xaZd2zZJPC2MYkWmfN789F3RuTSYF8lnE
nLF9ZuJ70zjT7QUOInwC0KvwbfatglRkP04DzoGigkce8cTBuayHjzRsOUXe
9U53qp8IL3OATzJzK4H8CiY0gfqeGzVnJ9LMliwDM0h/Pt0D2HgSIvJlKBLt
s7JfiiBMu1em/x9+f+u5Y5YkyPLN+5m6tarFhRIj0Y87nkndgh7lPZIECBYV
BDxhtjb9jiidIkvVkSXfBiCafjjwblzRX0G2PChdh6eXmYBp10mNWr7zVkCg
5bS6tfq5tekaschBaWyTjMAme4PrOikJOblQgYsoWYavXt9VDqc4nn7oP4rC
7i7wso0Bc//+WXxSgmsSoMGTKe8kJcmJWP3RSHQwWocdOV41GH1Xb8qNyaYU
fbjdYSkKQ8pcRxIDQI+5Y+WA1KY5NXRIAreQcMe4+ublTyafSbOcCiga58TS
SkQggysvSOnc6G83rqXbS/Mthv8H/w0aWNyC3guaMNSeG9G0PfETdGjNhC57
DTx7Ye5ol+TpX+cduG0KKKP8BgNxvdeW4sEfpohilLCyiELmg9ev2kqf81kE
tTOHnc4Ea9snRbEtiwiKo+BjacigpxG92sHa5mgnhnvNWOuMcVKtpFZxOLIz
JpPUpxCqJQVofitOJbI6hwJTAhUCxpbNI7Po8/l1slcD86YgGXmvkMsxWMRx
pfwfkT+cUs7XlDT46d0Go1dyTb4nLx2IPjAwq45TyVqBf8NPKNHfC6eEz1/B
U9n/fCSAUv2rMsCNW/lh8ojYuyuGlAIE8y0v13iOzvaCtb9qRfiOYSxD0JDV
LydhOXucCGGK4p0LvzCuNXaBTSVYsurHoKdIw75il8HghfScUtHsLHYH2jkb
oXFmw5NocS5Q1juRt0CCnqPzeK0a5e/qu/gaEe9Iw7eHZZ1Kdl/iaeeYtYe9
4b7My2aYEojCf+1B2x04T833igZlKhLEcdXgu5cyh1dL6bZy+L+8zdgoysJF
UwqQGs5m5Lmfgn9AzkdutX7AiWzQyo1RKiiZm8UiPLHjrAKYbzKQgUEUa2+x
mgcRFxUaPo8X+fQ6NfQqN28xgPbz8VaeNPIaJyoS8PuUkHOv7n0atGuy4qo0
cFT1Go1SgGtjlMLEcGtxlUNMRWze6+PUVrAgtuJXXRloRG6GgLCqZlG2KHZ4
4VsXwvG99QB8MG/RzOSp4IR1p/RyPArsZxlhKS9KwzKCoBBFTAXE0pNDRb08
o6BshdY/a6zHTy5We23QY+XtEsqPW4n76111gZbsvd0MK2Fcd68NKs8dZt/Y
Kv8xItFGOm340Nbc8PMopLFf86uZZkwPoklfyF8d2mqqJDXfQoLn84vuemer
JUY23Dl6zHyk+u+8mqjWLG2U+qDMgnrOBjtysnbnkZE7jRGAwzO5GP8K5BPt
2B2LeIsTfUUW7jtgHIXDawJucLjWSLV/wwL4fjx3W53WA/oItMxeA8lRiCTv
FyHC1EvMvq87xWy/fdK5XI+rOULMizjE6QeB29FfjdhZyJW9fc1cldgbH8dQ
0LxMIZdqRStEOsAa2h4x5tnepKR3MOshxnNHhXwIhhduWaCAgHFdpzm+L9Eu
geR/fbaPqY2bbhCA0OCEizbCCt66d2cQSuYP0djqGnAyHFepFe5I8MKLuUiO
R6Cs4djTLJlC5MEnv3WN4zrMUgcoka5LqpiWodt+K1DZsIwsvIh/EdOuIpfp
cHJ/9vb5vwr6x0npp0jDAo2BAbqEBG3hhSq5cx09KGGm6DC9NVf7u0VeUBIG
NZFwW6b+V9gGfclAgP548jOG5pBXw3/2v2ZXS0vhhJPlMxK3vuxvLdV/7MiW
mhQCeLbKrQZEywxFqtkAU11NUjRpq6o4jOcdW8Z0mRRNeBJSbA4JOC7yerZe
iJeYNBFlTeyQ3YuOMS046zjJTRKotFJ0LOa73J+Kmd3PL+FpWZqEK/eXdrGr
kHvUEyZ7FJMpF8xuFlE/EnIk3u3Du1U8cNkTYC9P++WsKGtCCQHUsfg4TxvE
FQLiuBwbqx5uFx3541XE7pmCD+44Dtbef7P/tkJKmmh0xnM+yzD/978gZDcG
1ZOGkUUc7He+MpdxS7nN5Mh/CE3X+Mf2i/M0nUzQDkJ8AJBVAUzVdgnYwwfF
zIsrVMRVtML2miavED9M85XnCy3p+vfVpfbh17rOOuHfNQTvlZRmbIAG6/p5
dAP3K/T0hHOlCG27fo+z1ncN01eumU22vkiToqOD2phCMBshivdx6IwnzXQO
369HbsfWRBBcfAsa5DPzzlllD4aDjjyDriDVWv8FwnBfBhQmufD9zhP95tXJ
jAhGeUaaiXpfNQev6Lqps33HhspvZY8QHtb/9ErrVKr4mI15CXLRaD7luJwS
Yrq2xgC+u2zYQecd/6OYYGLx2IS0YvOeJZBJhphKnXz9FX3Q4dZNrcQ2lgJ1
Fg7mco75zM8hLDgxFp3epWJ7Shk/827TXH+/jzOjmKrhwNFdKE7mIutifmL4
6WnWcGM/UPZAwpYG1Uub2+jg3RYBypzmuf7BYSWPdJRIKiTIXrY7PlEgTkd3
f9O280nei7bVrO1N5k5mqhS4aHu0CkYXhJ6lm46UXF8HXTE85jvj1Q67x34t
HVfuosKjlqEzeuCpaBX/uudGH19behwGyp+aP3KNWGTdC6x+gHjARZw/1eiF
DzFJaXcctfy7V6tzfAELZ0BUPI10+Uy9DhR3p9OM0CANYz2HC9mPXNdYwyM6
h/76e6ToPG28WYFoId4dEZ1oZDn+v8hbuEHbolCMNRQDRacMJF3Lh/rfB+ks
OCP6or4W+KyupqE4SJDX3So18hLnycQahzjDtVjs1Sb11Ldp5ljFaIUFx13D
Z1JK0JOkY7g6uKz0XBoteaKn5wG5vkDkgVqdm7qgNBx0BamTCSK8VPBPdOsz
bzXEHp+sBIPGkFI5kQC0b5ATMWiIFcKGqFsVHURXQ5tdz7e+6Gj7bVBisjfx
3ZMAv9JQyDaQvdOJesH8p9slXdmqa0qzBi7BXQUvtDbVXnCC2ZUa+TGDROEg
styqNJrXEiRQsoqk6vXSoNc6m7rcYlPGuQFjw90ac5lsFVA1qgDeYKBuKgXe
yAtmC5cMVI3JDctB5yaIp/MejkARM6PsFprNwiGNF89yguWCQZ5Mbf6ToEMI
l7FUUIqqluNddf7/GpjQ9z106PV6B2TSVDjMUOahWWBFJV+iE8kNs9Nlx7d8
wQJHjClRTWCIqnVWKVzno/cq0l9kIO2BtnF05kMDMh79dj1d4aJHCwlBScmz
D8LsYVpLAtPdQc9vA0gLMtMTZaY8Wbbw7cgTilimJ+oS9UQmHyvR5lrxO2O1
nVbNvJ5oMIGk5oNX7gfp/SP37qk4+/Xer8LNrQ7MJ9Hl3NqQNZxnzsI9jAn2
fqI+tlUIJgDpMKXMtISnZFjxfm7qXj1H8EoAS/A8H7mT15Uy9KtqJHuxaUTv
Y1iyqx1V4BMGjJie1nbtzs5gAau5ZCCtaECwlozSqiTDXqmy+UYCuW0GrxH7
n5m3pIa66jaCpp6rqBa6EFySCwP8MZUY2HHxdPPbFNHJeQtPpf6B1NbiemMm
vbEjGFyhigKdXAbV4gYKa5PLn4flkD3P/U4rJ8gSrp7RrRiSU8ZVomUUEAzX
SubkE8qkXrnraQn4pTh6n1/FrE9PyqekKCFE4ZhY/wLs9yZOlPIGVZZ40/Vb
O9qQn/7aeYUVkALSYYAPrb10hdG3MwDZVnw6NXzj+qOcGtZ5siT2wh6HkMCB
cUgKXGO2bdgOLY6ul/Yen8S9gNX7KTl6UTqkgrfucv0dyZVfvZXO9SkXiZ51
Yzp+DobDM8PkkyiS7woXcnLrCnqgVclUYezDrYxTP/CYcvIQO6ggLL/B+S/1
PvPZUXL5U6vzs4Kfb0561JoLeSq6fmYMcmCqlTlDRZfny4OizlaDbuuCtRhw
BRURHZRQW8EE9s1IDgJ5nSnQE4nLh7x0bM6zKUKF4m7zc5LkR19owDsY1RxM
xA+Kx5+/JVtZCdoSZE+9f1CWfM6bbYtTvF01hjbug1AFPWPAGo+jOvh4pWk1
6N35CAX4189hw4orfwkBv+/F/irHQCg+xYD+9Mnsr4jVuzZo6uuPo+YeAAeC
tqZ/mk/Eye0wojuwvD/ImmXV6gxiRoT13J6KkW4CDOoneiVGQXpupek2wDC1
L5EC5Kheu+AdNN9MaM+4WfFYOXYfC9OpCTYWMb1qcLszKF9C0USzzp96z10M
LmT6k/ytm7U8XQMGOAR5+Mmgv7CLfHRTkR3ttQ07G2QOyK+Nz1Z0FW3469qR
h6umzBLI7MEcFjwOqGlvhwHtr4c4OThQd52/St67LVTSX8r7Hoa1ln+EeYRb
tYhuNh2HxCb/D415CgyCtO/xD3EJ4ij2f7dFg1TFcxBSgDNp/hTOsurYIkaU
DXDlwRQmKRkegIF/RUIRJBcEDtYbZTdesO4MnWfMEjjbkf52p6jQmInN3Tzl
8NvM2Y+VQP/fvtsvYIlBrv1BUjyI48YR0PNek8A7glROVQsrcuLtCtkf1qUP
StAtxTWqOIi+XUUDCUUOaxNbwkVSP2bI+xdBeDGL5oklOpUAbtTO2Kf92nw5
/trlEbHNDejjHFZMLZeVY1mKI+YuJ9a/LFMT4WYOOF85gyHFlopH4izbD7Mw
YQMkeFdHo6zVQJNPFwpH6XnBvqowmo0Kz0+r+oKLvq1UTnyTiv1hPF4DomTU
vGVtblXGIjNwBqaj9/7uoTs8wEKLvHAuKKSNxT+hH7fbqu5s0BxdKjnh8Otb
WJVszTXjPr8vXG4LwVEzMKd34uVk2qU92vz3Q+BnKVy8+/8cd3rcX919HvWa
wE3kAEVkMLPTnrXw2YaYW0tmn7rMel2GPYNpyPUS4/+4jV/x2U1zMzrMI8mc
2MfwDLFgkOxxtZFqtUZ4oLwlKXrberJSmuq2IB0cJMXG+/RWSTBtRULdNLf5
pFjV4wgLOv/iEzbQc96R7VSkGDYKfg10VaQBqWEZti+MRrE2BNjYvwTu4DG7
tzepmS8jypiV3ZFNP0+OZQKgbLO+uCzQOHaAIgfSfbmuYZ0jAzC6uMxiw4LD
D0yr6Fpc9ImLx3lZW/d4RUQ3kkxRiRDf4MzBWBAkhfUilVX8Ko2GPqnrP7CC
+GcKzrFf65Pw/7dN9mcY7mQ+V+IAbmGLLWQeU+FWg1RiMgQvqQjqFM3drS9g
rJYtKCOd/NYO8ZLchSoi9dUFpyxpzWvSlCec0qcRuL/12w6N5l6PWBr2DruL
LUdEO5D6TCjEO8+WKSZOqPn+n5ikJjCbMVveWCkbAHEbVmSnCGQ9vkHyWzXW
Qxq+xjhMGbCANWdDtVxOfxxtDhDlriUyk+7gcweqD2XC9URVjELVX9EpBl57
e10kB6iQE03J0qrVK7CPrMotXSftIltS33tJWDCL0YTVn4J5KnsuFTYH9GUn
Fhv9+6628a8SJVkMpjcN949l9Fyn+lUO35EqbccxPtCwlQFqybWTgF+b5R9N
+T23NzMeUlg+/y9M+wdY02u2TOG+Fm6LTbilO9MTtAUs345iCoWZVIm+ChHP
iF3RwYeacXGFG3SAt2OtZZE0v4Xlbqn592Yw7JX190RbqYkqqIU1aXiI1juD
VGWouhuRNXoB0Y3hQ2leg5WPvr4v4LkcT5zqgI4YUf7K7KFo9nDB1IA9w+sK
l8rXb/4Y1f00vt666XsJ5WnhWaJk72ovheAf+Wt8ZKibAZxcTHrAzPNsfHba
nK6rqVYS4eU6f8vEsq/t/BFKM4ZvHZRxB+C7Nwo7jVwOfRKtaTVnUHQIa+sg
6Wuo0vILf1WwckmkWg925eET348O0f4Id5KDIukSOmFtMJd9k0Lnwkzm4gJY
0k3byf87Z6WnPrdHgi8x8OlaYJ7MDojhY8KtPHhwrZRjdK5FKShD/MaM5Opx
xT3fuSE9yITQPDSaB20dCiV5deWFpmjugYwYbRqIAJJGSk/Hp6dh9dBP6ZAV
h3Yb4Hs6fazV0vNgUiZpFed76nxjY6JuyF06z/HqX32yefahSUd635v9tk7N
LmI7yV24iNQ7S78GC7uiGsZrtDyrcyCQMG8/DTY1l+zjM7gWOyuqwyFinATp
AQuEJa34sHOmNnNUwSe8ffaEKQ1L/QZqqLsL503qUZw1iMiE835sL8996MoP
9bQG+D10p6VQ2md05h9hMuygoU+Rirm9dTCnXwoIXQP3cQaUisQwGi+oUwbS
yAyuLFzSyQ6BC2WhCygekqYmQlT22FCFG56LYfsP1WlKDo1g5dAVK5vCpYwB
Dmp+Ss0PJ89aGmQX7c6laY8EQ6JzUDwJp/K/ePspYN9p9qsYwjcaob6Uw73i
lTGA23OpRX9TRFalGlGERxmgoz8WwvQoJLSNAEXEQOx5EqrrO+HXzXkp/jJ9
pA5bUjtMjUbDv/liiyiAxv82zMP1PZ1eFEfpezZLHqVXorY7hFPvYnlH/6cl
RrgNLxyuu0DWRnSvwKfo0AwPPgcZF0lMBlgDjsDoHhh0ilJw4lnKeUD1vhuX
graZbrk9DcF87nC0QqP51TTZtf7x0rB/k49H16g7mY4+xtpUq/JffuhyHIno
OIIe6igx6CGfe9adaagXmN/S01QpVCE/wZC84ov/xBwowSnXBz/AMMQ0zTNx
IFZDqvD8Je0MqaWU16Omowr7ck1r6MYEGRTCtjYX3wkVkOCYffPPkrBoYwS9
VbLkXvlzNIFg8ogkdTbHycXpam3LcVk48vasLvBTQKyWnTRbu/Wp0kj5TfO2
FpMQh1JOoUKIIZlE5QubkEMozdqRkj5QOX2vtPs8N1yNmVtewIidazwwzLvl
+ttWStUyrJgyFVKiGETmrLVvg8gsLrS6CY8b4zKjCRsfeSJIfHpfUqZGThPh
WjajqyP8bBqIk2n0/3wgviImbChhMSZITkKqvrSN/CMHFk01s/5bVAihdFXr
Q1z8ecC1e+6gfuLm/bkKPO+6Fmf1Jc2or6HJQTDHdKDKmRjx46JDAIvhrNOI
e5K5jkK5ey9A93DNHdg9pSKBbKdXLuaylvxK6xEPlw7ZSVS6YORa77nlNj/d
LRaJWGeWitD+cTbLQUlYcA08SmIKuVNovPxu/ZCpVHJIpA5Ve0j0LaObAGmt
yAeFPfSck9MgjwxX1b2z5/XJk0TC/3niTRNEG9faWqFAeX0VqwqDCame5ngy
OemO6/USNdN7nVpb4hQQfUdJvE5pKtGGvhXfqtHAWwr1DFORyl15xM3if/l6
9TzKYrttRyBOn9rwggT/TZ92lzf+ObwlrjcNK+2wlz4RrXrWMCMLEw4+8Xjw
cYu0mNj654/I2ackC2Mv/T0nU3vgOOI0QeHTEKRLBO37LNONVjuIyp1Eq+9c
Rv0EguoMlp34+Sb/Usis3cY7RfPgzqOiuglJNl5vUFigZmQQWB5loNxsw49b
wncKr4cyNnE8qxzXS7HhyijsX9q58zv7yBIXLSs8pYI8VBfhZsq617EidDNM
Et4OzuqSl0uShgqLbhqXhmfZuuc+MkQObMU+KkLF1eNqrXUBgk6fSIasaEbl
aHTWiTW1P03XTzqOleKKMu6ustfmWKMb7EzQxGWVAIFexc0+gQU2FHsreDRQ
MnXOzdQFQdvYcUrgLFMgFTBhSTodue+dpqv5WvnMBMwSyzkAzGH7ZhzzBKpW
7grH/DxQi3bWxq5BtFEpF+14eePfz6r5gvS0jxzU9Wt3WKkdE3a1uYqnZ8DF
RdpgK553n9qxE91BA5f/MttwIIkxY5Zz1DXCUdqYd9vRmgl0xHvw4a1qOGAd
Ix7O1HAP0eff98WKp52RKqinwU5ChaiaYPk0qJrkmuN+DF/G92F5cQ8a4n0a
nMapdDvzTAbtfWLQDmCuk72LVAmPgl0qynQYIBtQ+yhKYpXfgjasDk+tQOhT
S/WIMbzpAoHmGiSwfDRku8U9FOLkycczQ4BiRTeRoWt9U5K1Nr6JDRpDAJBJ
D/qq3cjSih/QVH+pGW0uO1NT61PLVm72WjhTtljpNH3gDKi73NnNLNUr8vxR
n0QHg1rwIDgOHsQqpbh+9p8r1iXFa203UiGjWp1VzwyEkseP6lpzfdWiDMHc
Gxlg/1e3qUcCuVwZYyfzduQnwjoDWtFKF5lC1Egyjlo9C5yma3RRf3o4YKjZ
qT9ELRUbLpPwvJosAqEp5sgior/F9Mf6GXTBCzOPpip17P5MflfUtvDqD1Gp
zx8VzWYkS0gmvHRAVQiVzkx5gJkauvu8f5KEx4CTm7tRNnFTiHYgzLepLVEj
nzo44M+W3rQ3L7cVANvqsjebHXJ5d2bSBPTl+hJxc33r9vfl7cxtfj3VlA0K
7Xt74VPgHMQHwRRkkABlkAZZPnV1seQn6ahbBqnp7wT6AGVuxe2b6uEoLWaE
GPHE9h3vlCnlWbe0mjiOmTKhwjZgL4HrLvi9y7HHZl4WCaayPDMtu/ZP4yuS
kGCE3Oj7vzAyUizY+OGCP6vzutpdF3KrtNcBIkttOnPkldQIFrgiRZ2LbdtU
++KXj3l2KZw+qQuJOJULLONHLA9G4wjC8BRhRcCxiU1RIWhgBgRit/RHKH+s
lEcyI6kNnPiR+MG7lQoGCFkOU6AlHkK1DWC1yXhguI1OP4o+z4mUO98Qp1hx
Jo4ERsSkZsljId2WEqdRKA1JkqmP0nRgPDYqaF2EfVaMw3QiDiKKhjAUhe1g
4WsjjcB5f7ZdgQ8InuJF7SI1mUdsdenhOGZdD78UbriQTC/vfW7i1sxUt5WN
LbTnSJRrDcl3CFl+22MnnzSbtnAQbvFRcYjAk2Q9RrcI1hOnUgAO9xWqqZIR
Pzhg7ad1M8Qtz8qLhXaRfvoqdOVgTDyWksvubA/2Cyk+GpQ4AQ7DPJMtXLIM
SRn/7aC4cW2s9KSfdO/pNi+ayjyrWswoF8emLZJhzosK9MRpGQ2SHr+HgUv9
+3DZHd4+Y0c44I+HYv+I9lYxk3X5F8GVj0vDJKXuREHSrZKg+B2WlNbN90L6
H1BARblZYDFk3r19IgbpRSvojnqkhQVTHXCRYzZtD/gsCOr2yhIxNlJ9I1ha
xv9xb2yTUJeGlJGmGRxLXa0VMqBaC37FIYFznmPGu3cgoJKR9tPeH2R060Uo
4fnKgf4OuQ9mx+mc4ZRnvlQsM1ic65yYQ07EMVR15PSBsV2Jj2pMyhltGnzI
6JDnQCFjShBIoHPB4OJyA6Necm85l1N+wH8aiav8GQzVlnkMEu/nqT8Qdkc4
qE9sgBMa1iSJstsEQ0NDnlCtaR5vxAKSmnvMR4hXP9x8y9JpvKLtEh0ENc4G
WDLduoWzDKk1+aZtyRb7TIBsjnBN2RoCybp/RgnDn4sjDXN+uo2yjn08aNBt
PlsdiWNGfWt+pSr9EIeluNwzGTgz38he4m3TGDQEMTII92IJZTS98u9qGbFg
os7F0AT8NgYW9AtxMi5dWYvw44HzOYF5z5WYg60FCv7av9EiTeIWkw4mLiCN
5VQyUSiZU23Hjfkg+uq/Uhm0N0iohJQTKDeTB91YKAKceCJMMAXW8+8diZoS
8Le/6VV77x9YuatuQ4ZIE/X9JmC+zb9OMX7U06zk8DZSJD342sDoUEHmhIJY
HOLp7FksivhWFTXvVTQxQKqx1hWH7F4yxNv40MWLnuVF/9KUlfB+cPqLdV/E
TRklbCOM3qboyo+/QBNGhNlSxd01fadIi8gPUeXROD04r3OwVmf1icGtg+Ji
nOOVttp1LRC8GCxqz58aoTOc44BWyTlJg8M6x/Jvqo+rpwjLzGccXQqDddkI
OhoKALYdyeughYrEuoZFjLejiVxc0cOBjoEGVIZ19GAV07u4xYIXKJkpjRJJ
eMOabjqRxiIsuUHgzism5Tivr34GZ/beTAnbSZ7qF53ldjv2nW/OqnzPbFDF
QoiF1SPmXmvgkfOIQr1Y3/NY1Nvzu/AjtTW0Dgqw1Ja6nx/6q+DZkGxggqsG
MpwcDMhZg9iRS/4jwjOOvV61lQZ2tOz3OihVuucoIrtAF2EZAOzyTVbh8qST
Vwa8VY0+2PhZq2SgzqlB3pRuoonh1fJLGj96Bs0zUgvyODBHAj0iOyeJ7opi
h6JHnnrxKNcLzRkW2vOdfYTOPsHbGitRQLYd5LUzpIFo3bQ9nHNvXblJb/If
LroPT+YWPE+uG/OsfdA8+oPshN3p6SWvCTv3R/0CuTuGLIGLQ8h5QxYxAJzX
vJzLdPn/2UNT0+TXV4SjfdK7/a20zKPUMf+DcZ7nkG5EwgIVOy5YYbLpFQLV
0y3XtmC+/rxlNWwvI/T6H8Rhud4NVP+MvqrJ9SXs4YVOQTB0l/ueJIMQy047
zlQWrmrKHBNJnQrMY8eoSN22fFcWOgSqTeslEN8/95VPkfKBquKFGE+Z1Dox
48hbWjMqoOW8ob07IRkhyFCdRGsMgkFYQqIOMd4fxobRIGQvIVg+qoaRxihJ
WMkkh7PFTABSmo1HgDAV80k/KsBEqLD82dFnyXRlliJaaUOLlUBLlhBHlTYp
1NeeIumiZQOd+qm0SKCH/dezrT8kXQi230jU8pSXhEzjLQFgM2GnT9HRI93k
R3b5NXgKOTlLSBEeZGN0T4k2Q5AUF/F+rqIuAyo6w22yTpks8AegYQQ6YBBi
gBJxsILdENdVgo9fpwlnfyU9Ym1QrRZ3OmFw9Uh+VyMIohp9zRZcgAziCvyK
sJISzR6jxKwaeKau7qbUy/LdC0yET5QD8+fhwa2bh1w6JTcK3o/uzxvbrnsY
dClSKqreF6lMQykw7lrOWwo/HJ4m8TFMdXqmbyjw71ZEqxRUNFQ3jxDRES15
NyPlMtou0KpCLWG69vpBpb3DGv4TglS12w9vmmptjvmdmrsyPG1EpYfTLE7J
7Vg7f7kEYR+bgx5JV2+Htk2vanDJj7ENLK3yTttk6S/Z30jHMN9cHX7/QtCU
W9jPT2t1MIM7nLjq5kNX6Hm3OxEZLv1ZsHV8zqii+WkKkJBJAM6SnQnTvjld
lBG/3vRLfHkOCZVcWYhCOhVvgWE4Nq1iOZMmG2hYXGcxZIrgMxx8aT8fx/mU
Phddu76e1+P1nBNo2t1YR8VJT8PSOE8gpLXTChspiEgXoYQIOigkjFdghCQh
g6WG8E1WM9F8JJQwNr9okASZ1oyCrMfdoMUiuXidRyb0r9kbqkKcFwltnNri
PCp2It2p7qAFv+WuIwAIlEjhUQDamgYn7KqErla4XWhZ1dFy2vB00z5uSB5C
dCGfNLIsRFeqDXAd0deBSYMAYpUD+fPJTgc/H/5f+6aytaq3obMs2XySQHcs
ssJ1NMuxoxs69EpR5qw+fkFm9uLi0p98sxDfRixx/1rVSN1PFQSyqcWZahQx
EjkchdwRQp/B9aEyWQq+TIHZI/cQmGi+Zcj/7fdoiTRfegH5Qrs1BNZkjzrz
jaP8BCmpNUIS3TreAVxj7AgRrKgjf8eSK74qEsLq65Zn+FpLct2J2p4eACMS
RLVu8hNJhfReqgDi2vGWHmJUc6hiKFO1PjLJXnOYI1m6goBYE1PejpIph0Zb
QwPw6M2wDZGeoOjbQxLT7/vBSiCbaslginUEmb39IGL2rtlWBqK3IztckWfI
Mcji4YwyzNGNo89Z6EeBactP9qrgb/NNkCNaD7Y1a1N+bMXa1WVlwrrHIdna
Odjf71iL03Rn/WjtR7kFYfIzkPRmgoHxsubVizWBBQRkpvpnmtiQl1FAiW9e
j+6jdQ8itE9tDSoXOGhBmazlHcwAlQ0++1l5QFpZ7KkyJ0z+0A67e7OxeHlh
7qi8PNf6uIPVMYfmbaATLaFT2IeZTwf1IpYthUivkN6aw8p4hVV/eYC/D4KH
np/S6yCA2cgVCv5at1tdkqyXceac+7lf5HYAMvtwPWvSsy0hZFBuVJ3Xm5PL
2IlJ9Qnfv+aOVs3aSN3j0prmu+tLK3k/6bV8amU+Lb3cYndpLR4Td1C+vkKw
WOSsX/vlexh+Lcr6x582eKNfUQx5k1ANuP0zA1C/kVfsOy5gJrMJfyDJ4E85
S7Fawn+FfeuNFxV1mzmjKkg4ktUIs6F/VKgy3Y3qc4UIUg00L0QXHv8eL0/q
GfMA8+rnBd9CU5Mu4i4yKUe6muon9s/0pymTGkE/D5J2xklwuzsjoztmTLYx
TVQJbH8oc/zmqWtsdhrZ9RroegjPs2/rxJbjyBhL7ifwOsKbbWLP2YOQB8pJ
m92lpmjpnzD9wlwgwzQe2b1SM9HnTAp8+smkW387uFq5sOiiJP1L/SoM+u5n
iY07W3zZb39+di3GOwQFevhB+SYyygetnilcR38fORdmf/MsyM0WiVHKzoR9
xaTDdA8IPaIiR07bvi2G3QpB58Plsgfw4YI1UFf6JwyeIv1I2ytk8R8HYs20
425b4M13dWIm1QZP5OtJaET5IHru6+f+SSj1u/bbRGW5tNP/NOLrAVYU5Y23
5nAC/DTjnjWJ4c97jY6gUUa5431iwchZle9D/Ea31m0ORcjhw6BEUMg6df4k
niwJwX40s4QmuhNQIfvqxZjdbXF3rU+8foE7aQ+XGyNozirhBmGy/9hGeSLk
KzZ0UGITpipsj2JVq+sKoj4bFDRD/hxNftTDe6M/QV6TzV3QtnMFwkpKLE2f
4DbyLbxavmqwnyo+BlP3hW0HWtMHt0uOWuiOiBAVRlIeUZpZvpqz/avlAFTp
4lYpyQySojhWiX1Y4Z4LEl0Wv8PfJWwpLw4KqTUdVRILX82WKID8M6fquz1+
L+Sn5wCdaptco3ZuOht7MvK9At3zy1+blH2vBkB4p1mleGdT7HgLmyeDgQl+
DL3LtfV9LJU3i/zP+OOCBpH4IBfGj5NmuLqRSz6nBqmz+lqsEI/Rc/VQotd9
f89/GSAHJnz39gM9qA8ImUASOUJ8kmg9fnHU/9qkna6Nv0/SG2kII1/sziK5
bCIMBWkSIQA0w6rx1Kbao4xNh1fFNE4T+scv7CG+22zZuyGJer1Oh4vSS1op
MnnF4aoNOJMiFVU+h9cvlRZyQjiPFtkBrDtQIgc2MECLfZugbJv8KwTy51yD
5hiJrz1KSobX8WPYSGmygNm9o5mc4wwaNqKOmzR6tMCSp03JshAoXozUyUI5
e8P2ZohQsnlbPQNQBRCNJKGG2pvXp+pLxNDZe1v32/0HxY0F+8gw7UWjkDx1
66re5ctrUXCq6zMo7n9jIzzlcB6tlObRl8TNdrFV/SUe2Y8u2A0/vKDbt0hJ
bZvEaC63nUCrz6R+XTSJx53jgUb375yzcOzPCZyz/72Iu9AaGF/TftBQsQtj
2mJXVwIuy/EKDEwOjSxH/2IF7LVIt7jbiGfTT5Nbkei3PN7XvGrY1F4pv7tC
V7a1YS+j90+d9ps37x3Qt/VeHCfFfu+CyLrCctu1kQEinjYTfAWVB3mhtlwz
J1mDpkSwYFzwQq/mpciYb7eXNu1YeqhVzkQ3Vvfn3q/G1adFaVmWR7rAsXhO
SZVubJon9q9OufeDXfdflZGgRaB+sXp89nUBMXMtJy0Boil0t6P92FvjO4Vy
U4AnBwdE4ppnWAn6gpura0sRypnx0D1IqDrpd285F6yo9/3mo6sTuTXs+fL4
iSEZ5hpVzljl5CwaO4MRkBrkmsnmBb2kog14Cps26UTv2uVRfKekFLOkBMzF
myCJm585Yj3H6zEl/hvTq736QH1PBOiNtPkWdeK0JW6IY3iVz0y72ef7EOrU
H3mm9voAif01jK/m1w9TPtob9K3sc8BrDjBzsoe0eSabi17e8MgXAcLh2aQW
7jALQURddpVXie4WGe2u0DWkj5wt0Safvls+6ZAGW9ug4e3crAtpIejSnrQv
P9oSmaPoHUO6NMNCy5eCPswKJ4MgtDvaPCKAGudsY5VAGhvBtz/vD3RjCsaa
GPe6TRfbcUY0sXVMrBfHXgH3sESmxYyLKekgCDEDOKRv0HV+yHa/nKASAgJg
mdjcuZJ2VLCqC3DRU1TcCaSwnvNhvNA5xkYnzqB8nBBFA78OUGO7PDcVaUR5
IpFBz2wLfEJQP9thpstqz+VJp87cjAcRA/H6xGW99EvV1YXob1HBle05FqW3
HQpOTSeOBDXPND9aDJ/mY338oL213k4ZmPHIxiZBP6E5yRsgFkcGtTSAiy5D
AoklcenFQgZSOdtNOCQHHDr57I7akv6Ir/xOakYpnd4CCCVceppYZ6pJozQ5
isF7YeotsiDlbNm/bHrc9ZXvLP5hOu1fxkgLWtWMKr6EWYkcqoCQtLCmmsO6
99gyqhvIqRe2AfmNAlCX/oZmHRqtp+sqrygakdm3L3k6tVrKhbxEUS2BcSLp
I7oeq9tG+fQ12+DXbMBliv9Ul50hEGngsMCjrQsAClwhXg2DwPErTQY/JEhY
QrDoLne3D17Y8bMQyas/UmTnivtbAXYMjlfgyqrfotFQFZ6pR6o4OOmZ4ZRS
KpRhGL2sFalZEHCWqXx4J6rfgLBr/3m5M+8W9VRuxNCZHQJF3HW65Cbn0fF/
drBH/QyQ8IN8BCO3rdg307GXsULA89inOCrPvKpmljM64zcbyS+3yFQcDEzl
DLmOoA1BkFfCrM7bzGEYmesVhyIpg6hVu1Qu6Pq5iBz3UK7SLSd7l+Um72ve
ZJ8Tun+KRIJX/DwQVM50zRwrEoDbtWdGDZTE4VD2IOi2li9ZTSspAi5kEDlG
Q8yRxg4cY2/HLI7PekC4XVRr7QX/eSA590iZ8cJq2wTUZYnZY+bcIQmdbe9/
DEsq6Brr6vgHW0oULEEsBZrhBMoZdnDis3Q788/Vh2AMqcbJ+6neImRkNDc0
51TKaypc53RGphkoE4G13KV7PTne8hjnkw05aRryiNjF2yYaDFY7kjnBT0sm
qUMQdQ5XtAAnEczLuZspuIziPSMy5ooX2ZHlsgLfyBK2rqgyqS14ea8HKGBL
ciUVtCuUzkFAgH2Prp5hNvxEoki3ebjD6h27HlpIPVG414zwLw3W3HSRYKzx
2XJuNarwK2TEOzuJCAPdr3eT+i/WTXuAxjoSpneV3o6I2hIw6Qzi6A5epozX
Xq6vHp3KytW9wvwqjj/RrgJ7JlcpJTQnqs4rcJHdb+cqL/wfbLjTDBvCZRrR
YGykdTK5yAyIErNkOYPu+l/MadLBi/c3WzHE9dMRt+z8MjZsyvxjSzohSmKB
1v8VzNvgyQpJuAa3sKzahwKyOdX8X3Z0zMBQDl6qAVQ1BjOLfurj9JLPywGJ
Sv0WgXiW6hyv6blQufDtc4yBddbsJz41CrhI4B+qllLA7Rf6cBNWiZr2OEjr
rhaCmDSd3CFNQvNkFlkzDv6uTfVZbDOPC2jgP4iTDhkfC4d4vxMuLxycwVAy
9+jqiZntqowDGSxEoYufAxVP4mK1m65jweExC0/41EsDTtgfl6gOCEKPUNI5
pU465cgJdIWVrQm9GBbIePRxaHbtoHrDqMg2F12yy4WkAmvBFqcUrzeesv0E
cFhx6k528f8ffgP8NyNIORpF2ymUe7ssMUZhkW9UlZL1j2WajtTk4OOnLyHb
/lNNz1FNmgGuTchYuvIL8JsxK26+yeKVLuv9LBfbcLWik3APB7xdIlBHozSn
fqbtNHRHlZLS401cGr5e7oSt2aWujkMG4PfNCHTnt31oqvaufH3AfSGI1R/V
GojlpvZsxhavxAxPV/z7b2kCTjA4kLnF3VShYdjBD/svXfV4YzD6BeOlp3lD
QNxV8+ISKYVp3RJN3xFW6tNAqb+7ISpeJPDngHk/816PHw6r2X11FLedOsFl
R/V27mrrLki1qHJ5iMw+AxV9/dekShJK+zhV/zPEgDSuYT+JUDMk55SbLGU2
10gSgfp5f8OmbnVbvmss4rKq9tFx0lWMdx+SZ3+KwxqNfYYoMCIKS07csYGh
8tcW2zjSxAejwYJ7VemGRPR2VMG0UDBTFKB0CxGW4R0emXCnGfH6Lh4HykXT
Fxfske3uLRvvXjVUMBjtwV3MdIVf7+tBXbv/nfGXMtzaGBTQes8FYiNg0QPP
MV0FLDPo3V9Nc9tZ/YvQZoh/AXGmY5qXrQkmn66YOK9jfA2+GpEDfntCE8U0
vsDkNmX0XRu4U7e9kWvNtU5IR/6xqyb12UQMF7d6QicbyXnaQPHXnRv4ywrp
srccJSOQMielsFYP1fpa5d1gmzwko7WoUAa9qdDDGbO9o6aJN9iSf96YBmpE
HV2cC5RE7tRKAP+DDMZCcfVH2QOFL3q7ypm9NZuALepkt+Dq4ljI4BdWAAH8
Q2eeBbx1AIRdxWY5kB30UK1+VJFpKl9SYml5q3G0aqAHK8MrATLpPb/d1FmO
E1j/m9T2cYjZOhF6vYf8OliS2id4I6rc/8spLjBjIUVWml0ET3jRYmXzDSSP
OVzqB1fMw0IJFOC4DtpYoN96EidSFx2QzGOnZl9zFAWfpeBVsA5ypgbMwTt3
uUZ/cuv8Ni81vEF4+P4A1WhPN8jMNGQra8Qi6Nj/0tdmYHM30KX4nDJrsqpZ
B3k+LQMsjA1UHwLIcgDerff73AjNqTyAXzy5Jm3/vdPXjeL576p9ie8tME21
7Vowvo7DmRvkiqS2ZYYxDYqS6T0iUpJIrS3/jgLpKcLJm5Xjb9Qka7a9zf84
lMiXTIXP8NGEzFTIMIH+FRKjX5iBOWa6DXerLOX1j+Pi1T6QSd29mgh7WJks
enPKmsLstNgDyx3r17/2WfJ+2FogUmUMX8dCHAlel9YKtVL3xv3w48teOKJt
MFSVDYwXscr4gMh4FVm210yfZLa82Gh+VqnY+ua9GcxlvvEXsFyrKAmJppPY
a4JGbubY8FTM2hwUzgceWPEE9/jvx3qykdoniZC1EPPZX/YK9lDUixHhOiqf
21KmJtysQWyC5ffbOKz0q7jID5zKeKZyYpBPye8NINddJCDRdioqQy1WjBr/
V5DRck3B9MniWxqhY8YsqgN02evmmNV7P8LvtcJVVIfIsYHtDkZqOGC4JI+l
Mc37O3Nzv75NXK8pJU7UBvHhIpf6UCJW/fqith9aNklWCisbdxAzgz62gKkX
Icn9FCXPNsgjrrYTvhZmKtWsXrWchqlWrv3Gw7iJZlnFl+2FQ6CUAT524xwK
C1yKe5wqtBbVAKvrC0k8/gM+jd9kdgRf5eNY94FXMJClxD5azYXOUAyjeOgP
UkQSs7Sxc4Ci8Y91WLkl9tkhFiBVw42BscUoITfcvS70c8Cga+FhrUxhNY1z
j9b0FJNEZO5tvYN37BHHHbRaY1s06V+1+GSdz2KPrOIQfz4X+J/6qACv0RV5
OOtgAFku9Uv+IL4UtT9bpq7vkD8XwWKQYYZIGfKlvJGHNGtw3IdQUXnRDtMZ
8oEzFwYOmoKQLgdYsUFFIxGvEQiTmdGJUK8BL1o69GQGLRvKJVZZncF4kWdl
6Z35TS0ElxxvEW9RiqbTp75HX+WYMSNMgH6mWgromVCSd99Gwz5w9LdMx+3v
O76OUUIDM7x4ugvXx/1Pq37UrVoH3tSZwIeFAoBOYKagFJjPk3+KQTFwnUs6
NGHtxya4kovYJJ2nxfO6iO5Fi32gFc0paJhpRHYDI/ARITnFfxcyd5KwGIex
2aUCBvGhiVX9/Q6wU+RIp7M/YxZquvLtgkCseHPIvkCTfjrdHcAMrDRcLd/j
XGcwhcYeBPDvdKQ3xAiXCE8u7zMt/c1F6X55XzEcKFsVN9sWsGU6p8XtfQdn
UzvZe1JCDKxNIpIei4CwJ//6QU7Uu2C/M08vzOd0TbQuux4vJBrK3tUcHo1S
8IJBMNacXEHB4IhPp3I+n3E5e0CN2nh10e5BOTSAeNfqXA+07TP+mMCZvO2y
sX3VfkCTjYqC6vPdhdvg0YRQs0Te56BIiSoAJjb0r8o2vrtPK/JbToiQbGV5
XL/xQ0maea+ksrYqmm06SxVmumgZz9fuWP1v4aF8Sv3hUeLP/cPve6jo133A
n86bmdzhe01nGNk04FQOz9WTWKLmw5TZTzLBVfoVUf3BGXSUhLorx10WnXIa
PFaA8Y5Xmfyweroxnq+PRVlgLJ4NSPK8UQng3JUCMlsQL3Y21p/eS2SryC2R
VND7wou+zX2f8pmZ0anIfn3c33CLWHCA1qkmK165SMzHjmROY3v10CzjMaIr
mAhg1JKZ9VD9qsosDi1pVoKYsx4sOqEn+UN0OX59JJ7MiTLGpNh5+CYtkjyr
F893rR9NH7dvoRT1zUrjnxaVvulrT1OspwOqsAqFHCUTqWmjFu4F23KxygvE
3pYNCQFKaqrZPDKr133r7+Ei799VuL/sWhWwS8w+T0147wqok3zyzUl0LlIW
Vk5ni2/qjKPkKqpePQ0AVd/AXFxFHrLQgnSgEj3LzsP9pmedWkI3LorKz16K
9kJ78k6/TO/FK6Q3yRmEXWPCwKYC1NRtvV2HLtWSCNqciuQMFl1Iudh6THDi
JALUAVneZeB8DC+mCwZfA37WQ1BwL/1Wl1Hd65EkOehx90YQ46bcp2EsoUWG
lCubMFcVmA4DOZMeg9ZiqerHwlEbML1+WZlesq9dpMsNxexofK4Kky8NKvP5
tnGy71Yr1hKNceNtBzWS2C0+w7V5599WDiaYVKAocy8LehIm1r4M5Hdyl5or
5KBkBQzHN/E7AtuC/lxhXh8Chihp73Z8e/98NRYhbdS6LOrhSyOmuiqHM2ns
XJg8P5f46TxcOyrh31azqMm+9cdwV/oNYLzYjTNaasG3mEIr88/Yab5QDJ9F
j4C2Ao6NI47EoOPjWtX+YueikcH4ek5iRFx0PDt4kIZGeSr9iDOFntkMC9Bg
QFVKYjC2idVfxWfz4IRtWTqPwsdmnPHx5wqL8IAVnEfMZtPyhakA8aGmrIFz
tltpsNWWKDcvWW65QKlRc5qpQCUld9ez3TqcF90JKD45v08X/QMQ+1KGMyz3
pBFOeRp/IsHpLPoGJpDoBLd4bqMppoxVQa3mHybeLw7+i4Z6S9vwMiZrKcav
6GY0jmSd1HLlK1FooWo29R+bJrI5a6PlGWPzwehtuq3D97Df4XQ+pAL9uoYg
zDEfZQ2fIkJLoiqgMv63ZdR1LCjTT5ytLe8aUJcftFB382hysXVwy3+dHfiQ
+VxIJN6s/G9MAbnU6kzl+qj4kaBFeVdGZWZj8HZxHzsOb1zWXLkPyevCAPy7
0AzkQAZWJv2gbsTLPbo1mJM20vGs9JgAatiWT5qbxkXr7PErm/hz7XKw69Ap
zvFAJrbECIOH0N8hmnNOprSHJcXKTBKn9cx/T87TlJRxlsQa1tXQDFbTlUhn
D0qVL04++khd6WNUtQEdH10Fcymz38oW0KEKXie//FH7gNJa/8cb34so6gcP
4R9Z1TiBhjhDY3XQCLB+8RyD40LfF/7dsb/Jd7YBjGBdkU1Ia6MAi/nhT2vC
yUVpygcLS78CH1Tvgoq/YhWDS8PsxWan6nuBfk0ZW2YxnNUfjTjR0bK7nY1y
Gb5hXfvU/s/a0iJJ/Caja0p5dC65yxXUUFeIgZyHFmf/tjBf+zbvOSNtTx2l
UVKT8gnGw6fDsFwFA3uA2WETLYR0aCiQ5yJn9H9gu/CfsCjNrUj8A0bu9AHJ
gTAJI2K6IXQTEqouZtRr0O0D2FthCJa/F7dUsDbo3BXUzIrX3xiDBP6o1oB/
qGHIiWctXh/teez1WhahAW7kKYLKWgCPi0EvvkcAEIy0J/CwpoubNtqE2arx
bItHXnPr6uSnJXF3DWmJ0vp8WszOIOMuWmf0LR4p619OdEqrgMUogwF47KYk
3PLzCk1eK86wdyjrfSsbporBpnjTwt4BkG3J9PZ8w40yJUl/wS4pcBkgwlyi
xDwb0TAWzCtHwyoQUt2SXbIFiBpVNx0tvY7bf1TAGJatYDX+8+aTEd3DiPua
Ao93jhj7F76m90WcmQMOk2YhgNCEZnZKWCayUWHvOXeBsVDLkBQT03XZLVII
NSR40oDdbeYPxP642c09mqN4kfX7IUafDerq0kmkBWKJpZx8+dwvJkBST6et
cy3ohuh5KijIZGwC8XndKePj6vLQuVZscqJ+KNnZ/yokXU8TH+QgPpX9aqMx
tqQBMHh6mWF6i3JD3JnrgL2xirrep6oM9o2Z1DCnzRIeNwftI1+dt4D1V9tG
kkg5EsBflT8goEpu0H7OBEFIXiuNtEJ0dWwAUd4GbXU6E7xjhlB9XMILXSy9
dwVt9UuZPFFnRzlFcWVFsSv8HK+H61TphHtmusfp5ATwifUaRF6rigaxkier
bulXk/QLl0FZqDf11aMfVM1MhRJDNHYkI1heNO3Sh1I4v/X/R8ClTi91y0Ra
8roCCWRfauUmNGodcD0uwi2qdF+IjDl7+/LzSaK/22y8yXhSPT/A2+bpJkIZ
NxU/LN4XFFnOzL7v/1ifg9t0yAzMhSZrJgQX+ADzpt1+NbZrStsbZXz51urG
byJAJASrzznZ1zYDxeLFAV7UL66j+rdx0DcOXYwmZGwtEASiSzkdOU72yHi4
Fxp+8uvjBrV1S3WAC3KGu4EjFWpucu10b6yTF4/rkPgCEjNxLpFuowmnXu2h
Pe2AuqiPd76s1BpCbHYMlTbfBxiOJIpD+03ffhRJUSqJsL77x+8ePH8wdjs3
bJWHrWXIfG6EgyIAUyXvak6SUJsj8dfErxD1H1KMiizTyYsxr6wzi8PQPUaM
5Q7HkkHE3s2m18cASOkAXpBgBv9i8Sgl0WAHD7IHrJKZqUlUn3R2m7tOpeaj
wW8e1yKGJEnrbTjpTtfH2yxx2ywUjuB3tXAXBlOPphoK0P8OEjsvyhW1VOfi
42c1IIM4ZoHrEVUab8emrRPztGzITLbbvNM50Ar1kbQaXuV1kSC38R3Py3WL
C78X0qqtC6HfZEaqYVWg8IPabZwE6uNJdz0YV8Op6zfmwqsFmkhUsYKrH5CL
oWdzHbcQBWFYpkybHB2hT331h6nfZXlzb2vvltRyzekcT+B10IGq8tWICJ3r
OCwdaM/cpiDOljSCP2GEUaesB7yuZkiR+NLZo8kkTR1FP7W+D8YRn4MXDcna
5yf5q34ky7xf/ZSqH4XYVx3cA+w9YT/iHE52R6Ej5McUq+8ZPXpBciWc35UM
yNPW6mcAVrZG3e4eq7n0M/v+AUKdTLS9bZQ7UuM2ftd4LExdRaMytDHkxCHZ
YnhUffe5LVKnDk4paqjFM1xGdV4ucqJNt4FiFEk8sZ0srVEORf0VvahZyZ8c
rDzErFG5e12yglhRSi9AnzAPoAIAlcHzn21LoHe8OxFyLzr+Q9TgNwV44ALk
vfoO7UQljSNLuX0qhsZsfeGLcqCquir6w8OSpspP3PYONZelOVu03F+scX99
jAimmEDVOcOJeJSrgcQRdzdr4fc4YeBKowber/7WKUhfoZVovjGSx4SukX6c
Tnz5fCW02n5CYyTqvZLimlS0B9AV+Gu701ksdLNBNzS1Sc6dO46XyBPr2sts
C+WhyHNJAEXaAnrojCgG9Ty2Xwdpt9t1GB0DlBf6f7Z+TihQsQdgpVfJfKL4
G1iFOLqAO5nvui5pQMUgL1v73oLhtA38SqDdatXTsnC29KEKkiAiMv/qoodJ
CteFJiHDrbdKh3/RCXAtYzBjGL3Z7otlj/xhQ7rx1gXNDZkI7na8ivljjz+/
Kvelaowg+Ve2BcvKyk6fwc8LLLLKLwDgrADETCq6FEr5dgKeYQT4/GDBpmy1
V/UhZdbLIAkfKE/7kDxazeFLOC6DjvTN+lpSuN5P9iXRS13aQBia1FjdKwmD
1468EFEj6YpLPz2EtM5PNZs4vRW4Jz+Z0Y1cAKfzJScKxy4u7a3axpd5zmpR
JtA0CRlNBj7e7TIcRFz/KMzYf8lZ0A2NVqJ4sffNzMVpk7f7vGcGprRi77ix
TT7FSgbbmYPnRnHzNFNCeBRwV2Llg35As9M+zrWzazh3ov++39OPQn2rYo9X
kw2KOt/zl4/TQ/fRUDT3IakIhklbjMSh/9BkPj6Re6gCYL0ir0ifrQaoA84W
KXqC8medM2WO2/8QbwKlL7/EE4dE+GINaaRmNKkLLyj6k8c0q9KtRu1VMpFH
J0mCZKfmRgd9zDTgS8zWtvFjG29o8wH+aZBfnwft+wU3HHedmamSnaW9H4Jw
BkrNcZAsRatf3FokEoBE43gJHVjCuSPXGCCa14KPAZzlDdGfsG07jvCacP3F
9UcWL7D9VFYufR15vro8BNL9w2J8XhpIiWh6+qKYjlcu+KZwLFuT7/VOeYAP
diNE/6TYRhYxXABtox8+BgjqZpK9S0mLC1h0Vd5acmi0J8dpL1ZxZuqkZ57H
yrQN0iXdfz1Nub9STi/LJM1DfQuLvwHf8yOYE+Yv+yY715IeLPZEyen+eDZ8
eVhBNgrPNLhF/atKjFL7eialyao777K+akEsayNHBHp7+YcANDe9q0Ls1j40
YF4luUQ6d7WjY1JPY3HOKv/tppjzLdfyh6GlTDo49r0KACuuk4saOllnl4CJ
59EF4mqKUvkHCz9yW7gcDQGDHK/NfuFTxboe+m6/t8S3Qi0ZTgo1ZZEDwUQl
d0yV72rvsvKb4DXcS3WxVwn/r72qge6TIu8m/4gPAZffgvF9TbVo1W21jmLZ
A8hk4Yken1n1jdjTqBZhbHe4wuZKMLXGdN2Q19AGY3q8M+hoUkqYwUH2Itd3
W23kCRPPdoM5J105LMbVtAYyXtCM5XG4ZevGUq6Z7g0I7pGEqBLv9BVXaMhg
fX43AZKlCDaP/hL1gwgvglZ/+AmbUstxmdzpPq8VSvnkzdvV6nbp8QVXKTTV
qgvRpf0ZmkjMt/nl5rsZrsJxp8ZHQwZLRSUj/8rV1fiQirjqNBNNZ6FxebqQ
tSQZSZRrKdYua1QY8MnBgjXObcVA3f05ismg2AKVcvwBUqwAPY2LPQu4WYm/
UCkjiR7iZJ5MRIi4TyUDaM52VwIXwmORaGx31EEL2eoLGLDcf1gOvOkciyec
JISrLm5vzQBpnQ2r5h0nID0sHoM1+muRVRdGckQc9AVkQMAPWaIutCaDB/yO
fjlx19NusFwG1NUseEZITmPt9fOOwY5z2UJAIOdgZ6tyeWJx/VcdQIwqbdum
+ipqbDmWnrh/obI3EYrLgMuSEz//QvAwZcBmEOZKq/Yv61kLNEY3htpr3OpX
sPZMLcC1mqA6hDDNK8HP4TJCVcl5UHXe25ZwqZwRxobtZTyTEeMtSHvm7ZKx
61teeXbwHQcU+M5OSv3kI6ZYjIh2zQGdCSnLznSwqNRIhDkkc5DlsYonRXUR
zIgcCMKrn0KtTCOXH/bJWgwipKwl5N4kfrZXuwF2qZos77sRWPulKNkUi7/8
33SWcq9bL212bJvxBXTshwG1DiCXnMWppQchd670NoR57DqtsjUnIpdQYP4n
9VNwT7kpNC5ZoZrlNo7hPqgroeIgo8W7q+np7LBCEVYr6GzSl2AzHi/2AZam
b43m+a3ktuPOForqK3aOt4vRQwDvOXUI1muSog7TZRmmDcnrpG/t+AQc1XEt
SP8npemNPe8xp1toqP8Fg7kfqdaizrrK4nfPXVa/AtWpBnH5V5WsyK/iFqMo
Kd6pK0zlr8iwUMk7rrv05OrszZLIMADbJim8iE7GHR6n13ZNVkDZYqeBO+ST
Id0k9G7AoQXKbNsz765caTVojA6KNPe0Uv8AxA6eJE1kMrW02pJqoE2kwP/f
hC3t0KEGSk8yPRPSfY56sR3YqjcKsSF87Nyo/++7wvY0DT9c+UB22gT/G4Mi
GkDdcsWMwaeWvP85vKmUek6H3I/rutVDs+3/GNZB8DAyb2t/xTDtSq7pxAb1
5kHeT/8JeG5qGFnjxfa6ZR4A1VFNrGx+s5iS4d950Xf4kAtdcSch385oHCt3
UApouHLVh1W3HN09AELw00NtTVcuGQLZQ2RJcbpYUoXrOAj35sgIyw6u02Cf
9M03M1lChv2Ju8GyI2hHWfMNckSWCswhwGA4G/OlCEutkacDw+CM3Yo/3HWH
zlo4fak6M1sER5pWHxqRNYxEa6orKv34I18mh0QJN2nsSY/s31190pMqt7J3
+s0rjXvLgyA/RIHIzg6nhlZIyyhoDCK9OzLUgah81NmZgRPnzGgfirozrWXp
kEIDgP2L7Cu9s05emZPDhxaC0ABNjqN2JDaMJQW4m8Bs80B86AZBRR6F4eg7
lsRWw7PUOdIKtEepmVq3v7ncJTc+j/IhvwuorkdWf/xGfQzxBX/YYane0cjP
ztfb1CxNtFGTqHIr8f4/eZueMjKJ7wybmbkcKS6qpfou2vc/KAGCK/nXnVV8
O6DJ98JincRO9C7SmLG76SVevTJKumodhoD3qMOHqiuhFQIKL12s7TtY/QTC
US3V2AVZfJkHDYUu8K8TAfao6G8UxAe8xuUo90TKqwNdGJKf+JQqlhYSQYaL
ieIdP3QPU2u0MYiALBI3+RF6lvphUU1tuQRT5H5Y3Daq90tzayN9bmuv8mkf
bxgSj8ZZdQ2DvQO/YugWURBKVIBeFG9E//FR0jc3jaNRxC7yw7baFIPzMIuT
D3kXMVmLiShgvZL7MnWK+eLcQfw8w329f2ySPHqOTrRcdvhdbcddpJly1MWK
R6FRQD2Qf64jMulcOzLYODPw/4NJu7TkOOfCnehOkMeqfMHrqQrkYzwNMT4a
wPUzeDR6xLHiq6YbrZ2JM3LBNfjhye3D8pKvO29y2JmkHWIlzG7oV8EL8Q1Q
oBWFgmMRztqSso9KNHtuWZVvVYT+uYi0b/KXS72cg5vQ/o9ruvT7QRFZBjp5
wEvyC3prs8J4djbmkgwD8qyB+eXXf+etjDlXNLu6aebmPh2DEmcSXTs6Qzcn
9YddFIqjJ9WXw49dG9yrbluq3dE7+vYc+cyxPWh1xRYAEygwd2UOx1PBkTHU
Tbjyy3fHMKP6HFZtlHiAEkzH8KMxSqadhU2v8XhMUwE8c2in2CN5lFmUIkMx
JG47j2QFP9pmv8Mjf4Y7MNHt5bvVnPLL5Ne01v+aVqbvv6dNmEUhQspJ2oja
xee0rh99Xp8z832IRvOAXO2UlnxnPIzbLO2Jwr3sN0kAlE7S+8nWxYFVaM2O
ySdCc/jY8yqzbQVHmRUJBWutS39c6p7Kv+fmrSjly6kHmePFYsy9+cX/Rkze
DPS7qZrfQjClI/7EldLAgNtkxwujMXJD7qtwVTw9U9k81LxEcBG8qO4FBglg
8G/R521NpdRaSB4pI6+XG8yWTJ1OK2tmR1exwwe/KVrnEzCLeAnVUwrJbJHF
H+wgfcUQ9iZgkp/OvTjPaXpOlYcwxF1oSQ/dJCXrC1LrOZIob9qh5iT9VueF
myGlj1hkWap+l1FVwQJvKz+s/lHiOgZ66EwpVozJd1CNyOHQz20GsKOn9oFX
KK81l668qq3UgTd0dXphHZW6OKDTzgMTKIBg2x4zuxg6I9jWVjqivZLdStxW
VqLRXENV/fURE7gNhb7Bup+tlE/k7EG262C4fmkBD9aLuzwSA/h0vC1G/1no
eGnsficbzVk9effsnaEbFkqh4R2HMWZJJXzFbWuTXNoFIUUx+3YFyJIKVTpi
X4FSLJ4J1nbzRNeKJXswhkxsDgSctCOuRZzD17wZfY0ilJBwvmiRsaJ3OBhH
hPG7G8jPjSggtpG+9jh/pTnecbIkcm5PcbBJRRX2xt43wB0q3oZvnvY1mi1H
gMojM81ZJ3SynaAm89dxHfDzT0j3wfy/2LlgD+vX+ekRN0OYuzlER9CIwY/7
anCUdWixPo2xFrFVgAHG6FRnwmyJmku7Z2q7YPIdXnNhhGDEe+rZ56l9U/G7
44Sz5XGnuWzgXrDWjPNAejxAgXgSMi6Lr+h7KFuci9GnE9mCqGxoS1Uzvo0F
l4H+UrIXN684OvAWOrHtoouNgD1F4NHjqQpLOK7B2bMdbpsbKsWNO3WR7TlD
bjehkjf5F6QQfjAhjzvTLGN3nJeR87sY2lOAnqlq6orQVDKyYzdGXCJOXR/4
RH6NAk/gxooBkM40Cvjq7PPRCUBIz0Nsc8amL+ubI7vS8KjxbFroLlI5X1kU
+QsSwGR/fDCXHpES+ku9Lfsj+BNSsmEWnFEXTtiUmt8R5e8nJ/TuuelO/SlP
HwlokeRTiMeW0t2uA/59D/aMxFWJUDiwKURX3zNN0O9vF6c5w+Tr7at87fEF
TUJxwih1EDq040U6WOwnlChegPOQs/nSBtxSDGgl0pcXsMVzw8nf7n6H57s+
dI25Y48eY8zakL8O1pJ2sQpdy2jDwr3mS5DvWdFMvYyjFnHb9ZLQuGCeot8c
0Ysa5MBG3qXjLNT0jkuTILUla2lzz8ZYCBxuJjPC23zK8j7cuO8nL59qSXDt
CRZZjByPPnNT6oKBOJ+7IfTSkjVXnbdPYGjZrag1CuLIG1HEZ/P8g8eKESFD
imUOAp17y7h4Z7fhwa8HliDUBzoLyLe8pu1MBuH2QJHUtYi5F10lpLiaRzSk
fOmMgtuXh1u3/XbFd3RjRgfb1LC5BF8G++qyxCpLplz9T/NUPQC2q3Cs4pu8
c3FreC8M+jo7Ca5uVvpVKdCSy9F2WHX12cmAEYnZuu7/ngknmLHlSJG3tZT6
T3VzmNAlNYX5XxX+SZHcQzxshSRolEftzXGOwntb6+w4B4oNkcqEceM8M6jE
evmJMAY60LwsxX8ofwLid+BFitMC1yV0eWmmk/EIclW3/Y9vGF3f82+IgiST
1lzFNOeydFVJNMKc/8AC7F2CzXt+gAXIcF7X+xsjvDo98iInQVlcA0j6QMyp
b/yPTVlE5+SWT6Tk55phYvgbqh+NYvNWFEwLQzvsS3qsEOnBRS+shJJVMomU
Jftf2XpKumxl+yqc9DaPAjFcquwdKdiKBmpVBIz2SJFniFpACM7j0K0bc2D8
AwFL4/RDgCkXHPpv5Mrx7XPv3fxQpyRA+cTgnk9yAR9HnGtx0pDa3u9TEbhZ
2R5oOE9z17M5DebdzAcImjElSch7HVXRUuhIl6CEiNOFfwwJa24ZM2M8DDai
/ceo+Q+ABG50rfwVxLe7C3NO8O2HhUe73EkMWtveSkCd2ZZRoSeRe92fxz7k
T/DnIf1BvSZSYtMmzIpZAhFsgr9bVvhgaejr5cJW9ncWgvIL01YXMd7aHHaC
hIEsLDzOizUnKUQlw5xVrb+i48sU0adYlKM5giJeqctJGP4AsTr53V+rgwJt
VcQG1FA1t1/WrkCDEkknP3LHVD4qLoDLHJRFgOs0kB90Z4xUQz6xWhkcFoOK
teFTwj7bTccjiV3sXMSHDwpH+rP5B7NnhV2Dk5+EWITlZ0iHi72T1vyGKRHa
VIUzGhmqObEwrouCB0/12QonlBykQUhc55ctq/bShDvAzbRpU9kMJrzejBcd
6CD2G81P2A57mdTHazY43AqGA8gjEWF8b/Z+kTSoiD0uAkj9OZI7y+AtmMAw
kOPbYM5xRRFwdr697XV6LZxYXnmkSg1TfggNbpwrlcLgZMEHvUZ4VuHv4Gls
GVab5cmhF3he5qZZNKnJtHUhwxKgW6F7So8HcxbBLjo82gIbW0lqoyc5ggtw
UEuWXohOfgQ1AtAkhOHhkw5oVa4ebDSnCEnwVb8fAsbvXEfwDgomcWXvINcZ
ljuATtNuJ0WQHKD6XqBWs/L62Ab+JglYn+vTJaqWjPwXkPLaYvn+SBwUJymV
7X4OX5JcpDwDlX5LhBOLdGLB0dpgT6B27n00Kqd6hJsEhx+eWduOLoQsW6+p
ZjmiUNLAJtq2Qc2a/FLsjOgrWC1aavAOs6zyPbLY8G1wjW0dXxD6J0SYAfyc
/y9/8zOfaZuzLXGb0+EB3MpboIvfwNReax3sWu/+zJzL6xGBmOdHPbciTVqh
TkmFyQFiBfgAIwVI4dUDXhWCqbnsOCl4h5BUvtot6LFWu+QDfplVnTV3uhNO
TPsUEvZi5yQgTMPk37ixj0eGmNuPK9kko5ANCHDMc5sNSeAM+nksr4kOSdxe
ydCr7Jp3gU4csOxqbwQ8BIvN0XGcvR4rRstGSTt0HO7gAqpxwYHS2HU2kCQc
O8lCKKa3uw4Tu5MXXc/Oo/HN1exSIZ5K0aakEq/lOqzVAOK1dB6ZX8VFAA7a
IyPewBccvLvJKV/uY+IwbHlBKa7I7dHPXfn19JDf+yKUN3zd6JM9dwuRGoMO
Th04mSXAS2HM1/Th3JYA+f6rNsbpHFOd/WT/BARsXe5tnIeALRCgYj4FpYnM
zMrQ4E2i+2m5Y4gRd1a7SkH34KWV/RDgsqGN9nnCJOaM1ZaFUSBjLItgTNyc
NSOayAAaMIYad8fNqXbtFC8CsYvgFfZmso7sHMOzVbhOp0yzSi44guYvVK86
iQSE1lYZZfpJcj6EdKrHltkKZstD2chLHShoKJ1ob1BKxzUKA0TxI5KpEUoG
aiCsBVZujfVpJxGaamFIthoe/8sXUnYICqZDgIFqNdvatYL4Ec3Pp4kZLnAa
suxFPRoLye2qX2mmG9ZyZKGwkefm87aCCjufcd1AVFsqMetjqK4n9L5ivqw3
kecjZwTwCW3m6QSgA34kosmC/c9QrsYIMN42+RXGT+vkMfh/zCmymX8UDYT4
8sNmLWpauR79MZt5n1ya4nbG9MU2aua/Nge14oFGHp2HqBQwWb2t5NvX9FQe
x3OtIzmfzDcS+4Hr+HjjarXgqfzULAv14TsDt4L5s7iw3IAM1KbwnqPlvaM9
BreFk3mjv18nSM7rsExNRxttlyC7jeU7+hiKpzLblQkv0uogNMnKjXAad1EX
Ahk/tCqExFCtobfjjWQvr/IqvxqBeIAAC9KHWH+tXzrE0g9ewJOMYsYVmJe5
cthcNadOPEllZUGc2dZdEYvN7UYQjLlh8lRyUolMnxaLK3c37qrYNNIMqwCJ
HbJMQP7pfiACJImOHaDpzcPz//n0Omqahp4eL7H04W84qJ4VGvYGqGyUVu7r
yPwr+3fDN+7yF6iLxAHAHTh3ura8xcqPGwluP+84GVd/AAxggj66+zz26fux
cDliXp/2KFsxypb7ehICCxffctKjNCZ10bLJ26mSn0pUWbLkIml5sGhzaXQL
YbZlxf4Ba/OR1WGZFVU3Qe3CPsCQtTAvUIYDBwIADuP0VRb1FOPuU4+M7Aae
GAqo+QucIAgA6yDRXMQPgNW/0WUQsCKWNJV5ikc+LV3kjd2nAVveUuuovrJ1
NKg37Th8umt4xLaV3reWDlLcrrsO31yBgrZGmYcyoEx8Bqu4+7ynWb14b8H8
oW6y4lGKaUJzY/q6LKp7Wuk6GGfOyV5DIyM21qvAuadqun6rzqyt1+ihi0A5
DdRKeUUR+iyFmZtkEs+nB9W+iqyreKU/M8dw1DBrZk0+s8bQRNPa3K6Dr3Dr
DPAZNFz1tBH7Kl9UBHIEfdc2bkLZnfGSPEbQcIzp9nGeCpHkVpJ1uS6VyuNG
UCHPBXC6TaGvRDaEcU0wio85+du7u+peYLJNR6WV4QpxVYPAUnx+xgISbISw
kW1yubKjP6rAOBvcAY3ak2+EpUY918I2ZVJvi2dbbEmkmJ3DaqdqoRdjO8rx
tlxQpAmigHcpipfiidsRH2RgD30g5jrHAKLBUhkI9gkawQrFQEgLLAJi/CfM
I75ph+2HsE2QVqMWs/rOVDBURddDimcB6UxKHnp93fXtNjVhReQ5cJYREsr8
TqFdhJkQ/lTKwpJMFdNLdz7jY0lk79O6kbzK1+ArJDv36pkrpf1bz9XLPwFd
epIhqbIGl5nD2LWSvfUWtgDKYXo80ql8/6NQtt2/NclaLbeN7iRrK1OxoHkn
9B641dYNm2nEbTgQPc9TnwVz4oSTZevrNPDZXQWjx9vSj0AsU041Gk+Te+r7
QBH07hVH7X2hjKqwiThtFKNQDKtIBDAcIu9dDI8CCIRrnyF5RJSpO0o3tGQM
A+Mpjv6i/kbvZ8K1+0iAIUwIMUMDR4M0ES+3lGPgSZumwdeX9jtZJHa18AHX
PCLCou+r2z3amqJGqp+56ol4IbfG0CJ5gSfIrYVxrEar2t2YT69n67tgFbie
bvb131DnQaZykX5z17ei+entb7TjwVy2gv2E4MC/PXQg+UxoTX4Qmr0jJRnB
Waz9cmVFVgc0Gk/2Mgjij6O0oes6MzIIGsh4hQY1jYIjtuioXubyemtx4tIY
0n4sTBrhgjDctjk65MGGDaOKfbJKpNkkkGKaPG5ylxhosxvWEFkIwusjLwE4
NOXvOfG/KBnwQKxci8DWVMs9X8Ng9yNkoelmnr87i6LayRDpWD0NHSVNqIh/
4r9L75oeyUttkidNWbLo1Qpha9QT2CTIn76LrcC2XcyF0JfQV+EIIWRPv3sd
p0FRsjXOctRoFsXxlEjVrEp5PmaPXLLam8rgw4CMO1vPB2XNgtIY/V5P6N6B
hAn3MZRd+A/O+lCp+7/4J2SnsrLoNLuDo673jrhsvf/eFT4Pq4HaPMF2sRCi
8HIzLk/ScoDzjM4abmWldUopFpNWE7FG9VzW6hiahtYs4IgSNfOiS7WKAB+W
65JTCI8J4JGVjMwo8xH02tKisc0UGnPPdnPEZdn7f/HFzGXeHA0oLX3fMCd4
2/rjddf5EaKGvoMkbl/1xY+BjYJbreImK5XRSYZwpt5C6EuPwvzN2FgUmGB4
HxYbKMZ8LcKA352Qmzup0sXxXNIG4xPubYL2QA7YNWXZdGTvl/M34WWM2DRt
XeruC71zb3gGwEj427l2hR+LK71O+IcDtld5r4+YoWYpjiqeEeieynd8EA64
2UhcE+GhPLiJmtIYwUDZAgtWKflLfblQkTrrLje+UP6OToCnGSNRDWpCn18w
grtIjo8I/sr0xD1U8iVRCD/JKkbNeNTud3hPFNsToEZ2QKduU+IZSy21nEZv
Z0b5n79T9P46xtoC3oi9TAgoW0x0d293cLWHQ6g7SWtDrJstDdJ3XN09h9tQ
YpZg9M5kLPJSjb46dANGb8kdQROhY2Qiu41EiJ56tHA978VgbcUpu5EYSiJP
1ZrUZcYU2mfRzx6eZkXFmzSTNbNwTcvrWaIcQ++wzkN2y8fn5u2FyGCmBMz6
w+67DtAkYlbDiOa17/Emso5p6q3RWNOoc5yiMqPNr6tjLFzCPFCfBlfFsVrv
F1pZhZzxeuJkjKHZISZTrMcZpXb5aBKpsZrT5chuD1EmkJsQWfieOLNLk0OC
n+QldiTctdD5jGJriUfkl0L0taqkO0qFw4czbMRAWVTyewL5/httCibLOKVL
XXxp3x0Kc2BO/00RTTMaS49aw3KcoKxFnvwPqNQaHba4dAdf11zwPiJrh2cN
2zoRFhssR64ZoIMWAxP94KzVMxA7Fwi5yjW/8dftVTmdqqtKoZoH4PlEumFZ
LZH+amKYxuSK+Saj0UHUDoOzGEsHBlOf0lY2MNJZTQT70S0hWsfHxp+5YAGa
VYRo3CapEp/zpGFjVVX0c8o+FkMkXwFgPmnr8vcmzFjCqc7fbS5agK3BSkuX
8IEdzLujE4M97cdHBxF2HMUvIfbgiM4B3c91UErsz9GdIF+efJ1bKimcAt8E
m+mht+tui6Tn2vtynSaNcH2DyFNWJxlKARjvSBDUVVfM22FCITff3nQJUl3c
Q+BSQ3gBmKIFkoj6tPaPjkNBQdv6ssNwvRLkCtwIiUMc54Pe2W5oEdIj5VJf
d9pXPn6xdVjPQClsRxaJxe37ZRyUX5jl0m/F9eGZFmOlCuQ3PQ+Ps+egPtZr
aRIyVNUkG6U4cvVEQQtiOyr+owdEQAD+TK3xaF5TA67yCGc0WlkyxjitC+Wx
MOGOw8sXtIeYoQx54LF7THlt3xeellQV3hin5uSIkykI0YwNE5qAjYr94A26
j2g38p9LRYgMRKas7WsU1DGeB1ptoU70Z/0o2Iluy22zb8o6Vpi8vUXifzeH
xpLu4CcX6bjgtBYXGzc+z5mMBKmLxxKKS0ACNAocx1kHZJTZgss3IJwdRR1l
appN7EQf4sF7Olw6n3/9L8I/DgIPipn643/BRq9SqQ2oFlTZUdKDT3JRsbwT
GTWak7he0GCIRjU5oSFoq5V18gq4qp0csSvigs+yUOUFikgBvgqkfnDnnf7a
I/DAdwiIuMXyCvZTyWRHplWM28H1MUOPbTvjLuoOsiH0TCQ8kEgzDYrenppX
GUWBsX5M1JBf82wlFG7qp5qyLpCRfY4+RB40S9ESuvEUtF3aXbmF/ereMGjk
WzXygJT4Bv47TGTlLtEcBOoYLDSOkmDJD5x8EASvGPKzAh2Kp6Vuvf6IYkuE
09dAwt3pPixw8/L5eiNjDn6b0N61OIgLe8NE5XOEzsGXPcks6T7L9AEjCssQ
t9nkQBKw0nx4SM3oBKAD08BdkTbUsk155uGqh/BvL3kiiZA+mcJP+PmBzAEo
WLsOWaBQQF7iHJtbVn6z0hbUoGj0opLK46IKPm2ImrU4VHrNtxu8OaBkWg6y
K8sjJ+VP/MB5zZ7ibH+GGSQ82I6lQVl+g516y9liE425UzjRQwZ4DxFD5+4B
xGqxXMWW6/9MVtEcj2QNHoLpzDc6vEYXmfPLk3d8WEdFd/nq22+LrO87ai0g
PNmz5JX1Zs8ZiJjUJo2UIE8uKJASu3N+mUmHTXgveB4frEUsEyaj2FYI+CWu
4/RK0Aqq4bzwGHHoqO5sVOBRgRlBTmUx9nUgu410ha7x3FrAcYZjjXmkagoc
cjQWGy1HPhj7Y0a8JXpgqfZjrutIy+grQrKy66rEdmqXQY+DWokqAzjbegUO
nVVjABqiBp039zJlFeeD3rWwB8U2i/hHdLuWRfx2g7bhIvgBb6Ww3vsFunXk
xG4OFZjnomV/IMKiqhUithJFcnsUchtDmfIsj5SF7ppyEarDiktq2AfBQeHd
/s5sTSQfBpRBEnhYbTuwjHkJp9iPi+yUEa5hBmS3BCp6wUaASosSxQtzmWYc
joof0z5AbTwL9G3Pvh5+bEEAH0b8/AIMYXqnNV5uWTy0KJEqH8dWOH45hTIg
yR2txLtV9h343nUq4v1oUrBYc+E1cO5DQOAtGXZuXaT+1ggRp/lySTRpj0EZ
q8f/WJYA7/mJFkTFjtwgzWT3W9zi2yUlyi9gUKjJv0O4KSjTd8PUdpp+bVQk
H+pcZ6+kF8mZe3FbOg5w/3i+TeGJ1nP4JTs2OWfzmJMV72StUiMI+jEHbDyE
bYGRDa+UPDk3poaqoP7rns9Bx6SRkY7uVGVmfC+kjl34Wu7hAB/FFC+tmex0
ZXHf9ZMKhOGR6kIYCuzReymYw4+eBUjSq0X11Y7ztdC44vY/vyG/8xBjD2gG
Vg20DHRJmC4FYTvA8DEusKw3uSc0DEh36IG1oglPnj1V9PrHDQJLckTu1+0A
JQ6VdqAsSom/A9sQNiDpdJK32rQfimshaA0hF/pKJhIQ7uhLon5+Maxl2hR+
xuAkot5+6ZuVFOan5/EelRzYFr7UGLWtS1oTTjob7SK9rDHrh66dIZD6qmtG
ObkEVGqvwnyBZq+wazMcNmde4AUdsY5H5MwSHk7Ib0IZx66BeVP04/VP3lWp
lP5q9Kb65zENcV+vi9HMj4ARJF72jYr6p2O8rOIw3wRxN5cjmf41lKeygTqm
XZG/FjAJImS3wSi92FvGQr9oPKX4IX0vfUmoXKvmzwO2dSaxPDhzKP7EB0gp
ybDrpi3oy2q4BkN+98TB4LOoaOFyBSmhMwAlEneRfZkw50WmfSq0TRRRzPww
jNvp2+pnffsCXFtD0estN10xskDPIgJDDv24TnSGnGPMAEGoqNFNVm48K0l3
K0AfdQC7bJ+kgs2wV6Uq0yuftJ0Shzto2Q7E4RRCyLCUqbl1jGOCa1CNEiIO
WYLXPY4/azm1wwjdclynrsUoJaBh8GMXDyH1bqxzb+C0aitpyveHYdvq3XWZ
aEvtT6w18lKo5GKGkKJU3Yid8AhDVR8e8R+kkvKiFMLDPBNodYZU/TKWegNK
KXreyAmswHNCNRh1jsVihfcNo5jrVxJYFp3cF7Yt5HjXslmUbC7ktGpwOdoS
nkVBpnVfNi++7yoqGekA9vHoF0ig07TMDBdr8u/C/Mg/fyXqN/J3J1/+Dkab
cohUPPaNFJCVl+Ajpc4p0JqvlF7LnxkcE2IEXFs1Ja17AWQ6jwmnH0jk+/rm
H2wEeOjtA7ocECBHNYqpCUzi1Lo9cfYcG7oGYykfhsYI8CgBsk5aS7PUqQWv
gUM7gXuyMK4QA6idTuM6C5TYuq6OK+pd26vWOlcimav+MUHhtsveE+QM47M1
0PBl4D0oTECELFqnL5qu+1olhl2j5tT6FAuthsj1D8khoBCCueIbM2LjFc2t
HDLI3FLYyGCjhTaegqj/bQl/mks+6XaxkFHVixUQsaNT18t7dTyXCVcCTwQ8
8F+XkEaC2p1zzEX8jt4BOk/VIu3uxqLdb4u4qqvCdOBHixCh5ESVfuKI0NkU
sDuJG3KPbwYNWoNHOGY7jsNCcQ2xRsOIwTuqsiiYp46OV3Gv4ithpVNL+5cY
oz/FnSwgTDt2n4uUcd9wpfQ9s1LPbndLkqajVJxlLybOjUBH8hHNliEArXKe
6Fh0E1QwQI9MJG9uXllxY3OJDkkfuyqpPOj8SeiWu5AsWBmseGBXLFSf76vQ
6dqsCDBTwaTaLqkJ4RuIUF9br/isGbtpqWBjLrU5Y1dUHPS6VmfGrWqrRsNY
itwIeBWkNr3Mb1yX9OP6dsH7e9QD85KacMCCzrmJypogcG8M9PhnJMzb167r
uZEM/Jd7h/tq2RdxYFrG8K+89dV+8oVdl2A0CxS/QMXDnV8Je3Mpbm6a7ZgB
QgyEd/efYGQBAjQDIeYvS/6L4ABA5ABvHmAapPyjZbD09xkvPmzLOqOhFJS4
Dj47td188pTBiYOtx7yGRhhtjhTRx2SA3MCd/92Qsdwuq9IkR3zkVDl0enkO
pSjrC0Krk0hvtoXXq/6CZuIK4cwwBtkbuvdYwCmEAdCfd4i0LGzVOD+si0Bv
4I4R6dDmfiEyeyn+UEJohR9m6D8hu+cS9JC6o6ZB+AZpR44gLZFnevB+j8AS
u9C9sjzYE0YAWmxuVOQiGNzOG2uKuSGb2GS/9R3OYIlVFEaUSQd9bGOStvL0
oOnndsGf0kieGxl+CNArDo1dI58EDh5c/nKa4aaistZkiEGRvEpLSWO+50Dq
0GjHYiq06FRrAyKN9Hd0qYi3i120HBEFxYCd0M7H0dHARqfqyjhrQTfPDTbM
wVn1GbMR5c00eWGb6J02m0q8sNUjiliv3Pocu3IY+KVooYkrjVpo0xdX/LZv
JkRZgBLX0OamRsvAZ4nPi8wv6TQZtHyJ9SmzafrfhiZV3+wB4Z7xllWojm+W
ZgUUIca4Acn3dgMsqBk6iwTQ/Jq9k3zDQ0CGV2ggKxYUco3SMrw/9QvDf49+
DwikWtbdsUtaRaoQrBSNzWxXCp7YeUvHUK+TEXCfyS0GGGnMePLcbqJyTOpC
oejgD3EDb1a/uqZG+Ann0OEn5gdfA50BKqTEEbpYVJwk8tobTHl42Z2uOBUO
47A1kZEvpRiAehsYH3xeZbFB8cNFkDknUV9Hjk+agCc8hFYiwhJqLWx8q4iu
ahMIMTmrpYSnfXxjqbHMurjm8DEjoIRL2ZOWVi2r1VuYZ5CF7OuLnN4JaUMU
jZzJv82Yy/akhFWfo0dZ9jx4eZQsKDAKJS3gFNCRchJA3nZwbILZahPth6EU
hIwkUt2I3N2fmIY+kDQHU6BRnTB1pTTJs33W5WYgSaHU7k8XSdJYPmcImt2W
aJE5sgE1VuKEzvBbrRObnU7c4W5J6YRUfxxwsR4BvPaYTl980Mv1dfkufcqV
IhQecnS6eoXvR8A6+Tp/0HDj1wjuVOFY+x4ozUqbJls7uShESjEtBlmuLFVW
/RAv1OvjujatWGrg+W7lNhq6Ge4At245P6itYENtS/OLUwW4IBdGzOm1XuLv
nEPfEGb8jcFMHUHgAvNQ57rpkH9JXFru+uODEZ1FSokFJTKmD6AbgOOP3MhG
2hr8EBl6C8vTuC++wiBMh2hEj3IKizxNRF5+iax9jFrjQicusAOU1UzBuV7T
08/iovEMJ4PWQi6OxS+O8sxy64X3mnhwM/GlHK/If/MJGhfEiYyE6NHmYP1b
9w7QG1GDqe5UYzZMPt9N6EAvRH3wyNjgpvA7sTuwJVGsEHzz5AyiVv1fNTmP
9VfbzXknXf/yylz8XkhFlCRPnHlj49NeCAqbJL6S0P0kFPrJxRroJV8p2I79
ei3+luRBJs2JctHEcrtwpYUV4fUEiIN1NjaFn4NJrxDPBrNoCebOiOH2yalw
46xJD/l7nYXnuTww2B+NhTct7e2+xjnyBlcx1zrBNJhcCqn7I4poWYYW+fnk
O6FyPsr5ZmnBRo2FA5jeRo9enirygob1OjvjgsyMJ9Ht13ohmcMq1uz3yrML
yWXG5zYTc39S9qNVvzWhZrM0ZbYVOGgESNvztBmVCsXQg/Kw5PSPGEzKS1w4
iZ91laHEjZlpRrlQkZ9i6CqdwDXBSZUpjjUX/0f5pL1y2spoJnO81FQRlIGn
lEyR9tH4h1i8dcgz2BWHVqu9mifqTE+9JmD4DWPL5SW7knOVKpDNcCwHjEh9
AXLRWkQB6sBtjsqjxdQW5o5EuKq8b5t4uLKHFAwSsVed4ELIV9pxlyQImP0g
nQwUOi8TFmoCtD1CPpkJaVGFaH7OX7GIBjx86f0+YPrlF8/j83oINqz7ZGWb
yKOEN8FZTheKoepxxDPgHimML9/n2b+46zqED2yqyyGO3SEADjHzeB8NRN1l
3aLePjeoSXv+7idoCi8d1/DugoMKQY8riqvItVcjxrAyBhuoaWKxErSjYbGa
fLo4UKQUbXh6SOA2BaO7mmuFP/shPvZKxGXFy1nwck92aQOxSL71b5YQ+//C
MehRbGzT7iMeUBFpv7Q1aoy9qtw4YWbwCqN40HJNeIqDc8wqZ8+wpBuJC8Dh
MQf3Tu1Ny1TKNgb96qIqq9cql238TkIHnP3bRv9OBmyv6/pcf/WU2ZtzC3kC
U61lQhYUYdX9MJ71zzFhjupJM79njF2usEQIcqKvGr+mOq6p+ZcFAxaj0EVy
vRmc66GZsl/Qm2HQhTG7fgdD572Q61RI5xe6Swg8u0AuC0EUsHxArF3f53P6
Q8WHWwQX/YK2XUV3WTsYXdqikULi6YXELpwIf5Vsv6+IdzOfMmmXPZbMJXgO
2wTnkRFwXgli6WfFw6DVnUh8pahV7Z3kYno/dK7LphiHLjAEnhRQwf1S5p/4
n4vxHuCqpeEHIi0car8b1Ze5akxRKsGQ2aPS4xPSioaIJvV4WbeYXrl5YWVv
ugk+CwdaEJmOpfHvEYF/tzWBu31boRzz6RBibWoKRtc+wn1rcujbQDdUJjdA
9CTCWoYU0UeQl/MokCgfungEAMB2flxngt+CCw+gjwc8qV8Or1ZT6y9krUVr
54H6Fb8mG40gMdUd74YKEwoy1mnIj1dOmnzdrLesteyzbOW7cMQhc6b9GchQ
l2vYM6hl6DbY0RJWq3tzrKG2wY7tbTi/yRpYQ8+5wCDJKb17Dd4AbJGVUboY
c6ZiUGuEYY/LzsWObzA5SzO/yle+edevxC3R19kt/TVij0a15zxQATe2RuKj
8iGOd5FLbWc4xbWrjzytX58/dKEA4P1IGg3LJaUWnH61TC5ssT/Vcv62PvM4
PIWmPUFb9bk+FS/1V2i4Vdk9WRJZ80tWzaEP4sB9px8rsfJ5uo6H7WQMeHj6
JSXKvuhgBMlimKEgXVAZtaxf1qH+Ewup61BB/TTWYbrAP+C0SRsfCvRgZ1Oh
JZAu6fV+BGOvSNwmWqIohiGcunPQ0EFY/MXZk2tjowv1pJYVRMXOiq/2A0z0
lSMfPfUa7ZNEehyzOt9dMGPCJiwSsCVbKZuxLn+DlFSXiI8HDVaKOekhfH6c
3qto9FeUFUI1uV0I6qz3cKwlTCMDfFXyQk+/RN8FL3QH0RYSEe197qqeYAoA
jtIINwU1UJRtS5fRppsYDOxdIM6lA86e8NoieAgUlEOLxvOjajyS4u3CO2HS
0J1TBRP+s1Rn0RGi2p/RrrdwzU350YfExGr6KNnYuAriyhI4QPrf9djE7puf
RG8U/uFyBwj4LMHUZQefkxFYjht7Z5l6/eT2tSupYtTritFAFN27+yZ3KL/Z
+8ZYghSMrkHFFasFS/kKyy3Tw2It6L6DZhHg86HkrqIK6MUi+R34la2yc4sk
M94Ex3zqKsp3sTqKsu5rKOKJTlwnlN8XkWnDpyl+mLHupO2SpxBI+9/XjFVh
9IMYyVn3XGSsP4k7/LsXtac0vy5sAODcJ9WSC/7WY5dDCsftilzSvWFmZU1m
SWmHXaE0a4W2Jzz08clm6kiL4z842wvS+o0OogK5SgCjbXyUq0wWvPbOhvQG
wCEjxBY6nFGUkLu907KPkCPdZhgWPE3z1+zYcUanUCDNcZc/EcM1K0HKfThJ
L7zgwmiqGzsqCIwvvPUEePwcJIawyP0dpolLNwEV3yZmBWGBt2dmCAeIf1Qa
4lnSBxPGB0mXDcq3SBI9xp/kc3DjmfNC7sedqQ0aLnz6V5DLNSUG5jo/oMwv
Rzo+2/hRhPL1iX2UkccUV555KJw5IQZmjDet7kR8ILiQN3/WybRsx4WF8fEH
QRyY6zOhiTSAyVAWKYOfnWBUoz10uztgC/o72dw+p10zI1sKmd8HC6byIwpx
uMf3Exc8T76pIt70CX46jd4Yg1s0ic9+FVDRnEW+u+UjwMyOnz1g921w2nit
0DA2/Qxa0vKWRmt0ExkBfHNnOyP+RWheVw8U7r6YGmhA9q/0Kjl6P2yDteL/
4kA0SPtkhUp+v+vAV7hQVAQ+gff4KyAaJSDajizgNyGNqrriDuXE7Hr861Ug
KsY2Zf5gRIXoE8fwec23x+mHPZrYlQRjh8q+n+l/iRUZxbHTkNzPg2g0nUuc
VeImQjXwpTapzG54XvslLsRibmCs2kcHboJX6M2al6a0saS2EMLgmEaDPXSp
hzFUwK9S6Eo3XXVYivH78QxPPl19cyVHU53DdpTV8I2Dkx42QUI2Mv09KnAl
BArCKkqNhU7HQ7/vRbZqJOWZd4xCKcVWMYDwo51GWnG2w27Wq2W1G1dKmvOR
NOxvGlTOkmayxPv77UQ7GDEY9WUyK9yBAc5rLa0/QxKbszePBEJVHE9Usw3g
TGURbv1YBmDXxFEu3S0BL+WcE00u0nC8d0AcmUj2Jod1vuraZr4zpRsHJCX0
7Nj1yx1vsEkn7pg6tsviGL9ckbC1lmm93I9AvqhgAZRTC4Cor4FhS+8Oe3Ze
a6UrAKoqUAXWJe5dKDFKeClyDxVgA+vok5ZA34zb9iTcdvpNPhxzLXT4Acij
N/g1UhvIF0g3QKEaBgJYgjW+j6/8OFjqME/KuRDMHXLC65ebo90SWq/kY/XZ
swPwCZOg+Jg5+pe0NP8n+oLbxFJdtK7A/NFtcQz/J+Awc6zwpQvFwpglBJaf
lnHXgHhzQ5Ywz0D++oHjiegdr5PdhPaR39aSJ9MpFJ9ewhv0fJJpmGffjWsP
+QABQ3FSBn20+BNuuEO55/0ZC93u2Fo2SrDevHsA4gyAri2P4ERtXiw6VHyA
GzY31XdPy6lhmOxBvtCn01XChX39hutIipjqX+6PRGeE/IxUT9Pn5xDwTgz5
ZLEZ4s1/Zs4uZ/MgDsS6oDTgbDGSO2f+fH2YIAjylGV7uaN5ZXoMRVbvrGpt
HRTMg2XVbPeRYN69RBAIOM7MsgC3RmiIDRtHlAsGaqr0u5DePbAqTDAhtZlE
UcfzGbYfNam7Evf/QGBxxb+InTnHYmUWoMtm2pXClA0l82gjEI9ajyzvCpIq
D8jEuehKC3XdKsWjk81+B3lEXQrf4Aeget0PFO+gfPFuLuLJVP5u3a6RjwU7
BVVH93koiNu/Vgz2dvzrvikUcbFTwjCPQzFJUwezy8HzAL9rcx27MF/bTub4
0rTvOAC5z8s35JEBrcO7/5q4vWNmw2iwbQYXnLkeYlR1WuuCOPz8e1kysRso
ilXE3KUMRuWjbE/TsBizBQPVUTwR6sL/o0hj+YUA1FxtstYqHvvXxatJrEqa
o/pJCttstQtGdQpWft+d5mx1Z3ZRuUF0HkED6urigjaXT3zKVuE3KBur4xPs
RY84+XrZfLKbCKg/E6GeSm0kLP0g7vg9j6U2FAWqN0LFT6zn4j7Tm/3R+IIw
yjm5WFTkHKD7EHLamGwQ7YA+g2FqVukCezscyAgZxn+tkTtFwoOjUz9otoiV
JkYpuh+ltFfzhd9Qfxx0itn5JAsqjxDm2LrN5mNZr0w5TNe/6kLIVoWL1NyG
3luRMA8UR/JTyY4Qh0NHkHxMJefWr2ITMbMxwoSVFIsSTnKTCEc6VFBIjXDI
fNNSvLiBVn/32NqXV02iDKwmNeBFTLDZ0kiaNf2FYVhTK0w1RBYxk0JdaNc/
N28pSeePgNzoyHjzyM1UPTBOs3WgnmHiKPIi4v6R7aye9mBM51/qjlxO0VuI
7M5dgqXmcaoG4Rj/7nkrTGAE2OD3QL0ReWYxnRTHts4r8fYqcYQeOttQGa7y
q9K6frhplT1xfxrVKYvfHk7FC863fvtB+vlZ+tZYdYLh+yixYj8dCNNvnYiD
uLiZEZ06ZBr+uB/WWFzC9UXI02ePOLVB1zYhMX7XNP5TSDrgpYdmt+oHGKTL
2DtbdobqKv74Dd7WLbL4GOtQLbhtt2oHoayg4zgKY0cS9U44bgaGKJADAzLQ
tkRXiqWVf5Pd5OglcIf6yUs73ob2T70bkmscg5/ziO/8btu+/DKi9FLNhZzv
2fkL6dAG1W0RYBmpqF1x6CjHC9WIS2pxENDycJAH4ZqdwSeF3/u4wHp9xxVf
O0YHpM7G1k+7IrXiw38OjVtSb/TXuiMRWfC/3/vDzVn19x92N9r1696Kj5Ur
TxRr2uF/V6cqpugR+YpILGNa+qVtsWaqI13UxpQN+U7lg9++qvuiv1UGpFjp
0fZPO9OnQom3NNMz9xeZ40XHfcdNBeM5AKehZJw6B4qTq8pQW+FhfXdHZQQx
DehDLl4gj1kP9vfMTxEE/be++nh4VKbrfDpQvXQYrLKVaH0Fz1dDi0t/7h6t
zuPWOJnIaFRcL9/cHboFAnM5vZ+lIJZa0zoDFS7Qe/dEnd2m4FTZ/jzh/uLa
zRuW8G6W00IUP8lyqEJ7pLstivkDn2EY5jPafFxeRI2i5cIAg8IyjMj3vu2w
C/GLyZjLLiB38yy+2eVcLplkFII2pimwLl6L8nnwQLyVbJ4B4anIUca4XM9Y
74X2O6sWNwnFfnqpev46itmhdqR9QMBoKjYw0vDRcV9dDztzwuVeO24VomZO
W0tA9yLROzy2to+3si4/vyzAghYaSAu9CWyFTXCrk4FSO7qgPM8NkMbkixb7
bRLB9Irv/54LkKcpYgsKyegI7+356drHdD2zkiszjuL0WvivKMEUs1wecZ2S
kWionDPuQMK5uvH95OD4u43Bq7u03NjMeWJIQTuQVkXC6VRXMVo2H4JVOkhr
JQ2ySTmQvRPJIl9S8i/HkR8nKll6R+pGwWgP2IiJ8LnySk2zN2gQZ6a2po+z
jk8T5p0NTlyWbZiA0/276ijDaQbh5fUxyPAiiq7RoYLQa2zjIgo7BfFirclp
ohC41BRJoHDF2kxsA8bsbI34gUSehRk+FA/0DSgXqNP9ntT7gAEr42v4QEt8
OZLPKqQI7ZE8tqfNpJMUjwNkdTX7SfZuS9O3Lh3aCrW1jkfXmk0aVWGNKL7A
yCr9BNtlpnKI4It5tTx22IvVtDEvWEtCUp17RQQNH/qYg9SS5ozAP5Ms6xEK
JU5u+U67I0B7PvmyIkioXgGzu5IquXXiFbUjigLLG8TQlinIkLyjBMcrAl/r
uKBEUh9SMG+bP/oGchvtXiD3c6/a2tWsc7Ab1XbgwwSIrg7q4ZKsQaAuFsbx
huKyPlrlrgQw8NL6ECGGDS5kW9mNGUisTalY2UwtXCEAEOoZq4iDtQ/BGDws
Hd2L3cTPRsKs07NFh19twYRymOHgIKhH4j1yIaqnB7xcH2QlQ80ENnGaMgKt
tvqkuQt/m7K3zkjL8wJsIpRwJD2vqNFYuF+w0jX5gph0xT+7i0wLNJpbV/iF
1gBL6hoibImxLMOjKpWRTTOTKJFaKbDbe0RfImKO/8TFFSuzEDnvvkoXn0Oj
k/jS2LF1cmlktCkHpLOqmnfnxrxmjOHiH3ExPhIG29ZgzMKhcnxmRFhgJESN
peJ+klIY7ZLxYm/uUBzJ62FKF0brMsAlLjiQiW291aZgo9bLlwzdC35cOami
6O2GRQzTQPSHMD/dOOT9nu4Y41AW5tZD1Yg8bT6SYKXMwVhdir+HLrRQx2P3
eTm/KJnYBVw9l4WOc6lgVAnMIYDr6a2fcunDdQrUs7ARYT//h+naC9a9i8ei
vVgSyAQyZ96sXgkF4jROlZDgvKmpECmMACcSwba/sO2mXcQ9OC5PiNS9dRT0
eKBNqyorwSN4WwecO1m19PrjBewiRMionvoOzxjK+yxnn68DqZH7JcWSJhWr
kCJWMGpMkkMVo2EIAmUBFsY7DfD2veJeF6q++hkMmLp2szdsTqLOsqKnZEGo
xgUwOzuX+TLtr0woR03mmDYP8R1KxE50cPYtHz6fQ8QUseEEVUHREU7NMW1w
Br4Yi2lLrZZN2hWxLg85MuO+vcDMItaP5kvKZ9KYHACmVsMI0daIg2QH9B1o
4drsd/E6pjD1M9q9pbH6AHF4MgOTPdZP8Ueen4kQz5KWojUSNjFLzxLMNK29
6+7mg3kb08esMbFss09jMXme09T+sSr2qOH/C2CfHrrKtlzOgLlUxXhPVNgb
hvpIalI6x3nvQRQ6pwx/YjRsdYInFlPQL8nHiMJUbv9dQ87Xus40l1PXBFco
c01LXx0t6G+0Z3wnh1wjsw+SeGWCZZQwqxKt7rEDseU86NcOQE9QjKJYJod0
1IcWFLfvdrMIKGsrzF5xP7WDa/QGY8uNj35KVoQ0e5CoMxqYJEVxIdo0pL57
avZxgzl2Xc8pwvfNYe0aW3tFkYFqvplODKhYoannhGGj+x7z0VE+uWsu1iT5
sm9VNUE5dQvUYf4kAR4WV9lk41gvaI9cC0FEoPDTcJydJQc4TdhbpxFHADAR
3utSm6qC7PoiLpMGrYK99I6CorYXPTVQuQnVKw6+AsuOyiG4dOmEWcp8suIS
cJKdEB+7nwAqpoJa1YzdmS/D/L9b155o4wnsJfpjBet1jIr3v7dgkrChdcOm
nmFKnDv5tLtVNC5MR2nhh5kkAp27cuTs+YCI/8S+jKdaVMK2yvX2xwj7BV18
kNXklKnte41wcyWvw/G/JhVCvyKuO370fzZeEAoey6bQceAorVDsh9GZvhtD
tvzAfWsLy0KBQbCduC46ws4pPf1f+qLX2gmS4hXo+ka02RJHF9lf+cxmZZge
rAJJaFXniIoqiYY27FxAg5tMFJKrlebfghpF7owdNGYwIiTZCtI/fJ1wl4hT
xMBGYQpSF+3hMFNfsbV7ontt+/vIZqhwu8razawn8e7yoWl9GGyEeF0VukxR
jhYO+8KIebAyjCia/RGTXsJoFKUy/sb4s3EgGpFFTBNG4s33d7zpS16w2gET
BOykjY5WfITv09i+NtlJUczvOgSWaMjmoFtrfMGYJsfqha4xM1kLl9hEMfG3
dOBPZqTiALgeXzwJtiDVfKyj8TBlxDYPxhJ7hq/8Im8GTiqJXMv8B3XaiAnv
lZmJwH1fFTUyg3klvBGpMtGVyZTPZ1vwa20Bwq69KIB1b7/LhX8z6JchIU+L
MqVZEaHRw+CF2iHldFARlOdW5iuHJTLETfqtmKj3RYLXsT5DPEOnSz7iMDic
bD82kX9oc12wuYW/3zunMolJf1F8awz7JQ58niAsmJg5l4w5zz9XNRs2dleZ
uelqUG03dcoKJozGtliXpdRxvnUmOPJZCWGt6z1ZDm/CLwlZF1JREeSJPEJb
B/px6ZR8IIl7jlAPbkPufhr0ZoQ5B4h0utOMH+5ufu3vHTKrPkTZZkMGy9JO
LQFSzSj+ROo96UZ+NA89oSOIr78hgrLIgoPkrFEROLCeQkCaTh/qIZ5qG8UD
LWjaUeIN3qWZT2YiDbQipc3sQeqjf0w9Mf+NQLAr2Oc/Wh1jF70HmqHXQP22
IAoYh93l4+mgV3q8oMh6YmI8b3jVtirjK3o3qw4XWLofS8kwc1pA4VTX+tls
297qBQMCNnTq156bxMYnlOiGlJeUV79C6lEwdGsV/OHGlPlz1hBawbYeoe9Y
6WsT6tf2TIS70qaLNv4CK2Vt5+k6I//h24eFVhW0lVZu8T6PZk2Dayvie172
ekBVyJ4TGuoYdVvhSLPIIAmEeq/XYmIOPT85XiDi5wmJcJkmYG/0ASx7mp4v
O5edeDQCX1/yuSy2MDytYZpDGNSaE1w08m5yHeEn/2k2p2RdA+q7t2j4q8qg
hXWOcK8IalNBpXI1JpUsjQYe5nD1Fi6M0AD1v8o4A21E1uJNaOg9H2xLmD+X
6vXf3GuMHLthx8w8Gkk22rs2xy3Kw63uqxQ5XFWCbBOY8B1DRGU/wkCtZxpe
Nj3tQvfKF3RKjNuJPQexr1IYmbjDm7J4t0qSzEvTc9T9/DwB1DhFvntDmOx5
TMy+MBx6DWX3vz2pkr1dI/ANaSiX0m2X8JBfcgLJ7eh7V3WThtrbFFZFKnEe
SxRw0bCJRVQBzKmazDZbcWCfdyXIjLwstpzeo9iiuSrT1WSzvzloSCB4H3co
c6eSgyEZdbWSjhB64MEyBgNMFMsoPElSShM8o1rAViZOQXILw0V9ddzg720u
PmZjrXVxenI4rZNMVuKEEIMZSfQMjStSK34ML3zfjilzPkjSLek3fYuDXM/g
VJ1gxuGFj7RwbKRjgLucGHTFMfQa7PFBudzig1b7cOJkE/x7WpX81ju94DBj
y0m1W4N/UJmp/TykHfxw64vomRdWHNr2Q4fJU8M+ydb/kwTBUz6PiL3hCk5O
pV9uYGWCWNHWuCg/lCg7s4FBUvAXmPk4OEyD1975V3gCnXOkBLGNyiaU6uz9
ZId/RJvrt8B6v4vAdKOdZlg0xk45yJnoVnp0UZYqTL4dNlKAGEEur9XKsryp
X5/cDjG0O85K5W05QnwYlNIzBWErYqWMbBDCuwyUohkkKMPDPhnU/Lcyftjb
f0zCFzmGjfh78uN1QH7v8lppe+l1yR2TBiYFe2RMQpKGRKWz+RFJzjLDlpLZ
yRgW9yXXwn2VcR4VCQnA+CM/jyzzISr3IkoOz7Gy4/e0YmnZeoVktjhz+x4/
fKWwL3mO8rQPxugcnJcNj4dPU4SAGA776c4xlhkRAz7GRZuHByYfRjMkydPI
ysbnZ6stqEnPfwAEaFj8+MQZiNlhRLqDpLxVkLdiUFezbIVv8duRgXcRYEUZ
j+MMJGB5UZiSXf0vrTIRGivE+UAwvcolgahl3A96SAozy2z9oUWg+Lsu/Pgw
osC0pAtLPR1vuEg/uepCVpEFfZ2VGq+BuxJMMTs6PNfGHUvXU+9pwUmvRFuQ
FqTgRca2ph+hL3BtnZsr6gBGEHIdy1YeL1bxLGwAw1eh8g3IULhq71HAV6Wj
hRPp9tbL0pL88aLWSKs07+AygyZfRj/TzJzwGUhtc2waXUvHNm2jzlV+/cwC
QMaJxca/xzjQT1xOOy27BLJEfEd+GrQ3nH/Lr8V/erWtFEW5eK7F1qq115q2
AQ1nnzCBYM+fdoK77v030dg7j/dDC/gmpYlvWFTy029tpkVLijFbY2nzFnAX
KATi3BJMS+4YA8fTuJAhEJqRh7lWpMZGxnR0VdEHRouipzQcPt4PmCRwlKrJ
mQaXt6OlJ4fblZ3U8J+cLAIzdH5E5vrF0VgcDYxFjugsgFLnsqbBr9yhzdts
d2QIdCY+6YlCbL+3pvDyWQ6i/2J6LLcHYQacQVZOasoy1/ZcwTwKN5N76JTc
DaeBr6Jne+ronocJBEu4Jw849yhSBQWRV9dvrckfDuXXIl8elVcMn6rm2Vd1
91XSgxjOu/GUvE1FaQWUMRTFypqsIxDF1GnXTWtIILZ1lVs6l+HEvWJbKEIU
nao2uk21XflpocTdCXC+d/+Li7UaLctj8tDBIuPZdpomrbMtmfF5MqMJn5Aj
1pz/DqtP79yWywYO0K2ai6hNv/J9na5MgM5rI/7rTtLuwD5n0IKsUvhIP4A2
kbR1PSvasYsGkjAlWgHHC8LpXjW47yQs19zg/PNkcGXnUIaztPCjQhpNEnWX
U0JqfKIdWxMclxkT0J3FXBLU3msGevKyTwq1Xj1UsfvatxkFiyh/z6LppOUc
pj2Y6KdzQ2gmgttkE7GCKVuSwaMOYBSXunqAZr36Z2EqAPr+Kx7taCTSyGtu
HSN8zjCLia/AdrXisEFPMqXSKOgrhp+eSOx3jAg5Pda+OGU/N+TT/Cl2Bh8M
VA23oOW8q8B18nchh28diLEHG+LAu6u4ImZHDoxc24bVSbByYRGZm1RV3dtp
CxT5kB9V2IVexiP+sh1WQUAa8ASuBU1xd39Aa8dxuKuxprNtiCQy59seO9EZ
xfCI8PvJCLmkXj79aR63vyjZ0auK3+jsrvBwSdsWAgxjaMH3AZfh/eHZVQnQ
BpmBe5kXA7bD7MKOuO9Gu5f3f/MrMNnluyIZHiWzgXAPFcjUMwfZskgvqoNU
7nFMWxoSl2jYc6Kw9Kw69eVdtQ2JQTXlOjOzkR338KefQ5Hvi0FSUuEySNpm
D4ZLgQ5zKJ3yq7+g7WvxFFpVmtz5+gxOuE0VKnPawLthPoLQUsGqAIpahxjz
PG0Iokmd0XEVq9wfxGAsaSrpLyaCrF+CXkWWcdc21lmr3YilCR2362BI2GxO
mvwgafjs86cO4WUTA47KHZ+nOSxuBe+/1S97Ttnzw7xsi+ZsAHT0IccOoqoi
9MSZDDNjpNWMaHN4FpF9QmHdjL3p5MnoJkiUE/i4CctVNV38uWH4Q7WbJcMO
vZtk9OEX6lgzD4pmxVfeo48YaR3brzGjKBbVi8iJD0ru380VFwIK/UfukgbK
EOoW9ApdSxJaunf9J1tR6lDOa3WzaRzlxoGWp2s4T2+Q9ogZDIoi/+kpepl6
KCU3pJX2MqxLvv1bZOLDV7hIzBos4V6H/oRI2p1eBqR4xefuQNn7M3t0dKSU
E1VOQ+2tU8hnl3lYiD56ISATQXxTnVW6Qsa+C2RiBgoPP1gbOIN/l2Y6vnfs
RWFK2p85goMfWue1i56n0z7NtUgWc6EXaxV5GHc5DOiRpry/s3VwJj3BEaYp
J8pIxksntHS+2P6/pjcu61RWtiLXSkFsy0u5B0kFH9rlwSnjf3QlEJ1jMbX3
CQJEXdT9Y9bTG8Q3BOqZlgxu+X/ClwGbloUBe0x5c/vQRe73rHolet/uYY07
Wy98xbbzBL3GvEAvaRZ6Oa5T175PcC3pcP/4t7E+jX9q9Tnuacr69jYnwsl/
alDU8vKvJr0C2yCbooFH4FeXzTNd+uz6ozyWzeQ5iC1KevvDDMy3Pw2foBo5
nZhpw+JN1/pV5k4TN4Rac45FX/NYFO8IY92DtuBy4q2UI92hvqjV8LEzqRWN
027B2otnKzLtgoN4PYy8db/ygMG1huIQo5m5uUl47elG4wSBLF2MElTqpfCx
/Ilc+QmV1A5/IMDX2a6zeSdRihZH5rodDWS+74BImCkSvlWTTvWJ9TD+oUgu
SJCK4Ic3ktBsbJqabgLqY+IrzCdNvNO0aQFBGUO3tDkgw/CQKYLWMdurY49P
LJDSvk9JKMbltmX3gd3HiMJL6taW9jAj8P1MldGMKrTLyZ5uEFrhTPlVk+26
Gk6ssSIEjb3+KgaaKFKmq/bsYX0T/zqdRBov7xJehhvmCiJtTgRcILau6b58
o0nedo3V9F5ZdFazcdhipt97nLP6dyynIIBdC1HzT5tk2YDXRwkEOvgO6Wgu
NYaSnoYhg8VibuodDBkfAyTwPwOYggQ2SXe8ALs05gePLA9zf9fFUXZmJZ3F
k3bj2kIfiCmiOZ2By+l6/3tHYH9xrVeoJLxQ4h4vbuYPR88jU7/DKpsITMvu
hoGnifO5XiSQynmgDiDPqLb4wInBzPNfXZrtHmc5NT99lfIoxm6V86JWvrs+
38tAAQanCFOYi8e7cXPdIFrzip+MH15Lru1XjpHyp6Zqn5mePErt6faT196j
8VvNdQuDcThUgYw4vyFWxtyLrCKuvbmEdRGuE0e0c5ezLn3m2oktGg2pGSLv
9XbA1RL4yMKgIJrnSDphfJV2uFF8XPmYGH/5UtTMR2qfFXEgNYWBpzAOiq/G
80Yq1t3uGX6LMOA0N7WmToNzkTlTi1A/cyXnjZp6tybk01lVNR49DNMQi2Km
6h0CoDmkd+3vTmgZNHFqeMHt6VKFoxvF4hUDzpU1VGyVtbZraNbzfYe4RZ22
HWxe95Pvor4nYjYeXnleJwYIwKNvfqHyC3jurE9Fk1uL0I41upaIeg4jf8F5
I2tby32Pm1qxYFzCjJ9yK05M7IQuNSHmjfAV8uT6q6+fEJsi56fms4xA0fCz
52tqUXguNi3Q2oA3MiuCSG8V6lkve5Z1t/E9CEyNrMTu7JQqSLLRl+/6JWfs
WxLSAb9tgaHTSxNOaNK7yd5Uw3S5ThpXXCnYkOFhc+ne9zzYZsm4UzQqg6We
SEinthXdp1aP4ayJdYUbt2jPAQEBYX3LMZy0bcBVgQps2S9FLDJRCgLggYyC
Rf2IGpPM9/+BPyL8sh6vkyGlFAf8cMYMwUCTxou3U0siQ1zM+WBfxQ0MDhfS
9jU/91d1Mtmz4Zf7q7Ygks/zYlHKdfJRHIbtbJvmeAge43q5+WPigTqNOgFy
J2ZFug7c1RjJJmPyf3iK5Vcdc4Uv2Jo1SkDGsLaCLfHW3O9JAjIa028zZlsC
TZDyK5Xj1kkmuraEWUnOoIArOgO91HY17IM7IziCnYaOQMwNuNssI7y9Z5Z5
auhbH36RG3T3YWOTXqZOreYIDeQPDFgkbJqbxGltFGQG/w5nBmcKZ0zz7EJ/
fnbSfcJX6qo/mPlzTfTSKKVCFZ6/cIVLX9vWPovCxcMilxC2+Nmcd/GtHU1y
dgXoobOpDzz/92o3GECuixTPdCKSxQqkxPa+AK0/oH6GQhAetjbcsqvXez/m
+RVb+7SyzLj2eSEzybZ3kVo5I/pNxgF9bk8DYwZThsKMokhCKMPWQoU82ASx
oGJwooUUVlltLQ6v6zkV+RruUUN6Wc1yY7MoxAy4E6zDNN3azGf1nIY+3Lap
yuzB3U3oaCNir/AZlz8JfPYWPRhaQmCMCfjqh3Nr3OPPDAhN3JP9fipuNmuX
E3kuhALJt2InmW28AgE1vG9oORVRLsJ7YgZC7Y1/leGGlp48BICp7MA+uxff
4MdsdJv3NSTh6Y8zMQiBPCdCSdturcweTPX14Mw9O6l7Mg66v9IuBIkDkWuR
b1c90cBQGnHrYUqgy6lGpr0VwaTgecbZCZZujGe26U+IcbSiNcFrQi8jUUEW
tBHbim6B/TQ0dW3L1kM/mTIV2XDQe23FH8C1ezFeB/og6QEuhCATiJPBzX+d
wDg35IITcW3C2MF8XHv6/50VSdLtaXAutQ5H3QEtB8yMHMWgi8dgcEuZ/Cia
U2fMRbCvhyxluV2W1aJpm/lC2vE1N5s3Ox1Kc1sQZbF7F5YXJd/XeFAXPHiv
0XR0Qjl3SimIHsymcDF8d7sLwOhv1hB4f48eEL0K/QvfbS2LOnvLQ7qyQJ6F
uxC2kE+5m3Fno/eQmsC650K2OA4vw5yr7NX+pnrqQTP3WMqDajqIrawRKc2J
4/9jP+JkgYfXuoEeQYXCaqKDvM8XjCwwYLfro5dekPKdVNhCADmr2ItdUlr+
VslIWGDWUDaUKNdpQ4KQgpeAnfTgIZH1e4vDwDOkpEzOJORzh/60ePUacGqY
OKHSV/6rwRHrNGejLgASIh9Q1uZzVpJDX5wOBoOGq853G81ZFL009BkYOht6
DFpwdeyaSJmDQb1S2RaLYg0b6IgipZMSgAt3+AnqmuBOqRokLbIkihNLJz3E
tQmcTyyr9+wKpxNHTZSvyjwaQxlcKF9vvo+TB8iT4eG6vuhFaIZbX24qyw4r
/jP+e+L1D6yvmTnSWu58SEnqjVF5c440jOPZ9OvY+b+8lYFpeC3Ehr90Ospr
g1KNO4dsoptXlK2iyzUKan6+mSEuTX8f/BxZeWb5xNUvi+UoO6e6EO6nPhRd
gRuQqsZB8R6DEhyJtnsAkLx45mWthHxOGo7wax2PZYp7UplELAWbxwF2U0hP
XXs1qqhzrPt6fDxxx+d/cALIpVbKaQURglQlb2M8G1uwjBSfsVoJAPAvFjCa
9ato77LzpQ/1i21rEH74MS3Pq9CRhD3/B3SutdHVLNVzN/9QyefaGml/bcli
ob9to2VQB+ogXRC1toyMuim8OpgzVW4NklXuA73ZnnC18VTJ7f4elSySZCld
+ySPFaWanSsu31+esalzwjfu2nRV2jL1EInaYNLjryI7S2Je8omMr2YrWhNr
O9ZQ/CAkQMc4LZ0EfVeQHAUm4077gSwSvVlnDWIjm+Ih/kvEpdg9RcApBRMn
7UqAsBNAVBjsc/l+atQeEfLK6ZZOoxmSzpUaVydHPkZWJ+Tkl0BINVJo+Ib/
fakFMGGMjoQqOQXfzEZ/8zu8GjSmzanZKhE3edJhX1z+ngNecsnRH6Wof1ol
BR0o7chzLARe0hXsurNsULHlGZ3a1sk8Fl6PwzP5X12twz1RFVG+TCYQo0yx
5tHkSVwuMOKwdOXy/T5cOq9NlOeLOtrpxQlnKQ6lg/CdaFYuxtJ4TuQaBqGH
Vm57JOC913HZObAUh+W30ZLA5S888zSVCKTdXyQA87FR91n+wGWRLPAMQgnH
5MD9kW32UJr27hyEANaoejpHF76nWA280oTfi28DB3j030WOPNwhLaguTYMH
1TnpA/tEGT4FaGSSxtQdjTttgx56cX0JKXtscFS2fv686KmrDMZd7N5K7oLB
pXTDspjolI25ZgjR4VJPoLs4pVFDrQsGMAvfBXujg4q5huS9HzaELaoykPq9
ZZzpWWqw9k7ieFi9RVpAsrm63GRzIfMj/n9QQ3cJoZ5KJHNZT/4WeVE3cNsp
/pnUX5O1kXPtXg4FAJVnYLflVn/flBWlJ3YE+wxbF76Rkf+5mOUXTlOqzNHW
6qkQWlRUt/ot4pboW/dmvTfCFLXDtnYySc31BLIYJE5wTtUc1zVrQLcHfIF9
igZyjVoUavCDr/PDTRBwFrGKoIE0Ps5aIZ34xpB36mz1SdYn/hVGbpGOCbYx
7laP2a72BtCCs3Ls26EKX+Ge4y/qCt60hsP8cQu8L6LtHCiCKcWcQErU7jEd
+b4D04ojo/iMgjeocjhV8fR/phtbhaqkRkR3IHCybZRkPpMtOByq7kbKpuxw
QER0u3fBJYIqft07wi+SSY28KG2JCmT/Lans2G5+qnE3CEeXonG4kXEowQZe
WklbPVIR73y+pB2waaG3NwY6RWK+4o9VMkKDaVoWn2tGT+PPeh1rrj5mtrRd
SWDzHLnEVfeuJO+UNNAOdDrArnnzYON6nexJxN7Y3jP6yi29xn4XXwsSxTS8
O0hysoCYN5vmjKZR1WMWR8CvAI1F6Clzv8oIYUCsIvDpcid8ED0xAaEFOUbC
V3I4bYjDRfE4QNgP8PcugDloD+op8Mk8urkon/9R+avYufS32AMn+SSFuspz
NVr/GzdL5HH6S6DOe92j9jMotouyc8GJDZYRQ73mKgDZ1uwjdGruLdaFQAAW
0yFIJmAmInMEG0Ua5dLuwb/HTuVZw6NRPPCAu1YrlhwC/B8EazKjNneqVfPo
uhBzGoOwVxJDzP+PC4AAXT+1k7mcG3Y5sPjAyemYL009oLhm9Au8a3jPI590
OvJvMaZEg3/A7qRmZmIUW06/EafE9Uby9NdBD4yqcnj+D+LSUKDooW7ZojVq
APfCUTyDpWCze0J4mzUa7VWjntuY4FhsYAqoAJlE29DoZHYVHsNljqV0TjSs
m3rBiDpg0KONaEuhSpKB7ixARqKulov4ZmkT/pYvJJlBprYMSg4s+PcVui4m
PHzNkbV2djs1ZcqdnzlNEVQmp2KbJBZwX9nwlme15jSy2B3mYyP3QVAUVCEG
5KrlGQiCZ7R199FifyifR/kD3kH62xdQWSWr9DG3GQyKcrMtTKmOzFPw9nfm
AI+IfdTK8//Oh3Giw9qL+r6IkNL1orvSQ0GinwT2AnIMgB11GNomNTCwRx7Y
2ULQtK72xU2REfzshiHptFCG2n7tnv6socSVaap5HA0fCWwrkv9jCDytKhCU
Lqi9CJQUYymOHK5Fe070AZbeAmjQZaeOa+D0EDLkDnVYT5vRgppu4gpQxl8e
Y3LCnn/hCTqHi2dugdRiCGdBgxYQE6MQJbPH7plCuJHeZGQDoP0kplqNt+46
Yb4N8TZbqZJfWDDH/r7xXTPGGA3o6C7p1Rp2fCyxWNKewCetyApeSiruKSqZ
dJVUb7o+vdrosJuGk7rqFy9jjbySNyHLzpMeQKZTpXZc5IcIxQ3qxBqxESDH
REhiZMKX33bizAZTEE4Ww95lZnxHkB/p1lVEdom0zGov1F/uP2I1YJ9cX/J8
FRCUMnsBRLOLqqjh8oJRqY7DdjopZEDa+/Nst085AJFdqLv/crTkkRDABmVF
oNG/Gv5jMa1ys/nME18+Zg8suxWr5ajsh8PHrld5OkMzD7TlG5Oh1NaOUwhN
yZ8tIpwwI/2t+sClOPA2lhnmRcuv5CLYeggsIPQ6/au+MkI4Iaknm8T2CRvJ
AocO2waXo948WQk65UY/5sekHb/7qYe5a6m4c5zlDy9iGxmcLnWJfCnJuZHO
APbpgzV35zTEfCWLafG/vUMw42HJuSbVsUqGH2c/8g/jlYUuKHgKunnHWOFc
CYVppABVht8wsOs57rE2LS63XPp8UZ1Zu+7tKQWLVzoVTwHJuCwXVpIKGfJk
1Ai92FqFJurM3F308ThDdjayh32ySgHMQdpWfGiBABLkTB/vTLWiHzSCwNLJ
P0bRJthPIYBOU043s29X4JNAxQi+f6MjmPzjZF6D4rTXMdNvogaxa475bRjQ
K2hVZWZZN6Fu96efkCD4HjnODh/VtnPaJZ6+8CeZLlczupGBFCZ09RJBzNHZ
62P5x8PlGn3jMb0wSEGNOZyUW+Wok39Vt23DvmGpThf5PXo0Lu0dadwVDGdG
p8NfcT+VPQi0JSyeF/vUnXcne5kRx4eyX8VIiEGo6y1duijl2+FhR053NUUh
yecAKaNsaccRF2qgEiYRtCzh42aSuN3DIyCy35PtqHPYJ6vHBjbmUEEPLyK8
c5WNOHD3IDXKvhyCcUXMpJlN3TVMQk9Pgu8GmYa/HLp7oo+dgoPo1U43ukQ8
pw0JdRfZVY+gyBOQYSzBXESohMLuVHUjyesDNYu9/sfyi6Xw3LY01TriJuXI
VS7orocARXsHKSOC8exyac/28fJQ7VYIq2XeUwBvrq1xxlb7q/FJAWxtkirT
kFE+bLAylDp9Ug1KtnKpxRVER/CnlNRXpPHMhvyK9R9FJp5FfqLNyBPyoPXj
NKb9eTsuIcZptC7UJsdzaOseDIA2wlh2kK/+qC7mi9Ywk9tLFEJdpqfi6vaT
hk1qydlSq/6AhTEjCkdG6VRduN4jKuwQCqrwN8CaJCVqvJBnB9wUC1RuaiQC
Lgyq8aBcqjh8wouqnjOIjdfJ+Jyo67eZGbZ2TEEQWNlYtVPGXx4W+DGadZz0
464+Fqcywvrv8ozEXZDaj5jVL9GY0TRAoWCqvFFl3KU03K1quBiablSqqe7v
HNUcPEKYble8KlPmoc5aYodjfR0x7kuqT7t6huUiZB0wLj75ztG6k/DVh8eb
v4rkLoTpW6Q3xKzSP63FOJBAMu70juvCWkBuOshk3PeMpMr6a3juIpHXVXRI
cAwAVgpDXmugS06eAogM3T1rFzP3bZI76XwsGFLCRMadBozEOjFhwjLn1NZw
QhAB41m3mB0YQKF8mB4HdIK7t0GYBKFAXjVVYZfeKveA06u7EwiXMd+LZPwh
2v4Ru9TLzk7z1nJFYSDQk52aAbSL5lhRpOUogovwN9H6gcix97e0BUL2qjT7
mHY/YtYMkBmva2HN8Um/RvopF5j4+3Xl+J9h7YMMGMLzfXpWa+/S0vZPz8MX
oBC4lyDAfP97qL5XEmnA5DT4PT4YTlG/RX8B8liCchV5a6531AKzB1szEj8O
oOlkRA3R34IMYNxhjRGjK/jUzmqNmQ8rGO3JFUyCyr5a+mzB/AKTeSDwkdVl
iFqhLj5PLhVL1uExVFLyenYXPOyO2eWLsRK4IEzTEozTrEegNhxd33GiMuIt
on6NBlFdmJGrRtxwrZ9z/Z66UAMUoiuEoakc8rZ+yRnyLBgAULLj65/0uyqn
twOtYWVOm1vJ8hMN3JiQyr/YLHg1r912XILMTSuXNWsXqDBgsbF/PFzbxE0i
5pjNPvydLfflWEH9FbVLbRteNmev2/Sd9XRVkelMBBJWtiU45h/hq2ieBr4C
DjJLV7bO1rVTHdvlzlhLMlCyBMfZcYsR/IGSsVlKAG7nvpYKMkiaa2ubEaOF
EJPj64X1C49ICR/sH/DFl7+z02uUk8wuRNoLZ9nwFrtF6o0YRAVS9u6cyQNN
zyvmsE2R45X4rkqNF8vi0WXXEGvylrbaTirH/5gkBz7oRdAzVnat8PJClIDF
voYh70Ix3MzItMtTwAvTR9He0kyCytusWht9tfQ/9YqQT6E16sDp+PywQtnH
vRKEa6vQnwO/ISmdwCDyj672kGwBHrC6TqdUK+XTPOJyED9GHY/jYeBNNlYF
5YimT4Dky3Cb61hk2hvJarXMz1nKdxuqeylsLXYQBKzQyfU+5y0vHjHXks7Y
y9Wfob8KCOoqXpfUrnNnd36MrOwn+6GXadP4KnBxphwjFPK5kS/eX/f3GC++
ARftKBJOpWedsBNVS1/b1FzX7pLyDGbWpDJ9dVQKHDPWFqlPEyYmbzEsPcoV
ljNAk5mned8pcoZeBmKQhqB30DHeBYCd/zspNZ6QBcjZxgf2lvFQhNTzxCLz
UkTFUor57Oz0mfe2S2wGfGdzzvQyi1yqGnb469iOv1aBbCOhzg3z57/TtSJq
G+jGsVVbDIEYmXWWrDxGHn5Eu71JWW4Ty5iZ0Y4SQIZBr4F7Anglw7A5PROM
cpuRLpgCJWqDdAHX16yoEJNKr8Y6DjzLTr8Wn3k3lA1cjOgbmUNDUMuxhxEC
WYM4amk/I/XitxOwKwUD3eXfVZbtXZIPOY75ukzBWcJUY0IEHA/0q8JGKi2u
AbuUdAOHkIuE2oxobKLyDDyTJsnsB1fXUtafKvKnZ9LGcCPcZMTLmkUKdVIj
Ev+tl0xRR3CFgUpkNQz9l9mLhSEdw1jYE1U40ExUy5rvyVE92PogrTtXTJLf
FVRhThf+jEpw2BYCR5izO2A1qVLHKv57wNi/SnFKFgqXWLKQye7Iw82Z+x+y
T7I/MQdpogo3oTf0uaJHuVsOWwCGxIDv1hlHs7wovJHIf7t/c+ygQm4am2vn
7qRccR48ZjPgREHQAI83DiUYohlnm/SmGzgrv5e5sXL5DW14k4mGpcCECrbl
odhEtwDcTvkcJMhyymhDqLhaisrRohVlaL0NBaTZERHcGZa008edFvh/Y8BK
MkHM8r5zuTy4jfBhIdWq/RsRA8SwBMjWj4UBn2xzihlquE8S6mZa/3L8u+CR
vHnmP3zcQbl+J2zUZyhYGKNAZyY+pPMnWf25JXYrgUpQto5mqtVRZ6kLc9av
2bXdw/txDsb4Lr+y/kU/v4GROx0DGrWCUwGVJ3w8H2IRc3ysYqzgapNbZmCG
8Fv7jjPUIvGPv+m0y5RLlAWV1xI4JqX1GnDyUULo1rPhAflqPEZKJs6sN06G
sRpFAGdNAWsbQw1KAwDELTJJyA4D4imGr/eedifoZxUHxbTNBXQuF0e8sqYO
Ojy8b85OB7e63Ie9HqMP/ttjeMiyt9y00WPES9rZWGzV5fvPaTY0QPskqexT
0MRg5elrLeftiLo5cwAh5AajAXKH3Xp0kOhiVdchucCI59bRErMzcKcJdAJE
d3CivT3lzeGZ2CYo+eqIk3TrU/11zmhKYENj2UR0z8BlnTdC8R054KRRZaio
IrpgN1owABTSs65YlY1W6V7j/CjFnOfEcZNVzprk6HWGMDkWD9hFH/nj+/Mo
9b+6EKcCSlxWFrur5CDZeWpAJIcmNxnLfx0ZXJ+VhdJA2HdejRILLRRTYKat
cyhMyjgQFbGawYcjenV2aaMMouEe68FpWA32iPQ7+zLz/NZwhEyR/aoZDTpk
ZgFgLwDjVZuOLXugT70/yBw9X6vCs5txrbqAT9aA9vvs4TW6zbiw3xnvga3T
xhgubaNYMz006hwnSXzkQh7X4arUeyVN0T1eyRtBC7oH0HfF1lE8QaGZ3Hf7
Cc4DP0hWcR8lWe5SXcbQiVxPXY5V55Dtdwc80AfGKz3jPT+TXD2OM9bDIWF8
nj2AA9Cv867IVxRHn+/6KknUkMRgd3s9yuL8yRDG24ROZLEHqwNWIMXlQPO7
ansQUx0yNuMrHoNCmUs74IKodmMJtHROTQm9vqONSaPmdqTaLb4ZBGXvHqbO
q2K0dqLC/eR1+3cIn7aRWdT1Hzw3bea7PBhBHAv3zuHETWymrZa5U2j2eoZ+
hPB4o+Nt0Zy6tMheHsyaU5ii6E/lzhfKT0a4+AkowIfdohLwEWWzRLLbyJRD
lRGvhfU7+/UwZ4s3qKF0crOB9m25yGcxXSNtlLvp2kVOc4kVpk2BkbhSO/dj
VEfhgEBcHUjVTGIUlfcfSiUJ/yO99L4+4cq29KOOCd9w+bZXkj8cOUA2zqc2
JRu3QFdQilscDNHLh1mrc4OXtiG7TxEvFxhTiC68SgsrZL7vu9shfp8wOq6K
DNbehk6OCXevBIh3JG6K6klB7FgsjYlrddOnw3kpZQNeBxIXtgx350kUMG6Z
iqDQCj1OiVberG/8gr8P+AqCIhvl5LtM01YQWUbFJ84LNetiTusxXi+Jaik4
ffVXHyipsXcu8pcJuYuCbD2EaH9PhxZAVDiu1LSVpoIGeObWGibXge3hn3MG
uc/oDGaqJw1GI1sWsoVGTC7zVnO6+0e4GSNeuENuyDjcETF5bWvD4QI0ogtS
SYRE/lMXbuZu41hM2Xapot4wG8VxcpFoN1WjXgxV2IirL46//fcTcdB21iOD
G6slfhOXpjXZ/1IbYTIvkALUCsHoOWsfCjMBlqkntdktotT1Phq927AK/QXK
8IEaY7bkFHgQRRPo4v72kiKdLIgc2aZB2h88oDqHUUpdO5zhAJx0er7xvrOu
bSnPDXeQDEkJO8lYyi9JESH+IBxU5KRVSep3RpZQn+T8/RXM55XdLJqWoFyZ
x++Fbf9mCfMGNdiyy3fRT+JBLG5f13VwoipiufLOby7Hh9HSQYlU/2Z4uHv+
qjAqvfEMQn1pstF2FJqENEaJbVbwOCss0+BJNlWiIXO6y80nHnTMz2XZGAFM
BT8LM3m6ifJfk5IGXkuSGZKj+oNFLuceL8dyMm90gWKTeSQWSNux74lNbC8u
raNpZ01R7DpuCiOmG0YwARvS0zlJIxzC6ZtbGxtiqvYPMt5KthkliwB0tvKb
MhwC78G6FFFwv7VKKpLYqwoGdqwNY+IiLHqW+CI4oUBKJPxTJmy5uQMFSJjq
kvnh0ImvsQx+OgTUgYe5ktp5N/eB7S+uu18DNmbKPDkouumukMjUlpi5cmaX
3z3aMyKkDrvvrpDZfQqhWcKtIBSXgj2xAPDk+tjiu/+xfNdZ4KVNDoRh7Etv
u+xPQtXFokHli6nAdvZGYgG4QGRZ/p2ixufS2dNUvSTfO/xfQ1awZo22bYeY
1DoPfZgXtfcJ2U1e08OTmCIK4KmhIwzKZWsZdufIobkVEDI1EB7a0VWH6Yfv
mbhsOjLbjADVTuj0ZK6eH13RXAZrZLdGiSfL0AuO/s8NgTUYN1hRXe/vduWp
d36enPq1vvvr/9v4ZqKX/wL65fhXo34UdGBgWLQhbz91pwf/p/yQf2Ep8CAf
Loxv/nS+yYZ59MJukNbqVIK35TrVL7uLPIXFarzpJsvFM/zgYYY2FSDHLfT4
HVqOOj7Tud/FVnC38HQzvUTQ4s8XTm2TRkU5bBfpWjiW3ExBqlsq4I3RWMBc
jiQAJDDWySO9LJfqyDN3RSTIieeGfsI6DpFvJ1TNuoXh1jfLsn+VCwgLVkgq
VUjaz+K3P5dg+acgDlQM1xph3tsfV8lEnHTxWgI2KRGEQYdElxXuOwyDmL0j
gd7lU+LPjRHfeXLwBlattR69kuHHgGfIAiQEdDrsaAmuCvyzqMUQVdpSZLcJ
XQmriulOOb1EVmORmQwIprVYe+AyL7x0XvLed1TzXjb6ZUFwEYojCfwocz82
qNqymaGH6xfDFoZSmd995YGZEViSKhJz29VwN/vobHOHNKQF5DLBRrt8kB4c
agBNsU708XksCKwmKstofH20Ko2a7zN2J5vkjENtVbG8r8B5PwqL25x2q+Dl
Ng/TGFNZz88sVU/02ic/4V7nGR1bvxXZGBri1CLaFZaaUtpva7+Zh1wakVqU
xxanc9jHYYS7I9BG8dGh+b3PAKgMpiEdFzB/L4JedWn1GyXfjA3hSpL+qU5U
ZhZ/Hbd1OvqOEa/krHbnU9Yy1fpmeD6nzcKZBBClPzs3PBGoC1dGoarfCGVy
4AhhR6AxxMdIrdduB0wlUzCWczwwJGTPfsaD1TtMYSB4GbIysNqDjGJL1WHl
Z7NQ+eZoFLrL72+e81hM98Xet2yQuQo5VLIPNcftkMKjTu8G1lpWiHZpTDKO
PSEY0ZR1O7k0l+iu9ztn5SY9x/ZzcKvsijAmFSE1hsY/ilExwDJTti1lwaZo
qVBAb1nXSLFNy6fqZrSj5IjLN6aVXIq7A8tZo+rPpgqQGTIBkd1r/9EOchQi
/D/C/mg0/JkbQzRC6lfR9GyJKrrhDwfinuMqdU3nqDN3Unn1fFBR0J28euUF
7F/QvKxLwsYoFkLXWC9JJ8uMjCsVv4UWjUTyfzXTNrvPJe1MEpKH8+JtF6VI
ULLdVPqXq5JSd59kH04kP4fbhfmi3DD22JHd2mUofYrMSec5+oxs71FAsL/S
F+bSGvDnvZby+aVof1EGwvFEt8U1SJWgZe4Mahrsrw7adOkcfICig29mpO43
D4TnY6Y8n0Y2ETmZ9ZBP38nF5sN4UWZYkgGoLY4yw5uaL9nwmww1AJUeG8pp
Tu00/20yhkC20MdB8J2DgQmJv5S1eoRjoWWW4cikd4czLq75ma2G/AMcGuHN
Co9YXgPQKIl+VtTOgmKovGf0Tbq6z9srSKKNFp4zrLHFuowAqVnkM9tghmGq
sOfa4Y134/Lqybzq3JCAQq5jVPzTJ7zF2jTLNb0fr4cBoAyhDul2TwmQpmJU
9vQ2+RIBDyaytmTu77SqPqisCVY+L9cie/TLURidLgtCz0ahldVAQfreP2xt
7jChtsYkXNGFLjVcAJ4ZMZ3q53uEBmuRJgWGyCRe38xA5OgSQ/3UWZ8DHJwW
Ct8VPtxM/cxZfAk5q7ITdB3M00GJSsLgVWZDQxAmBF1C7I1E7a0zqXeWkWoZ
jjjCyj/kx/GUxJt9ltF6/FLGHEOjOlu/JOQoivDgnCi5OPMhRkEQlM7d8/DR
icLwuvJvcK/3GEq1oZgZhMbXfJF8tO4TvKugm0U/sLLSrgBBC9N5E8/t6kxQ
3brvtR6xiTkHlyk+7Wts3iE0DZ1nxlTaZmVPYfzUxmMDwAOLAMIGJA3CpvaL
dDEc1S9IbP5SHi0tOl+3BWIR1jyaFKrRX+4ek9fLeiwHwx7Q9C8PkhuXt/gu
B7DRoMAKf5oKuQKHsxoBkFbzqxH2MJ8T4YuxJrppa6Fp9wJDXF18CSmyChSg
gjFK/sVZJcnfV3/xwzsFUABXmfghWvtYsMdWEl6Qwrsh03bowQ/9MZXOQ1zZ
Bbrdx9iQHCYfF/h55Khccnmz8uaiwMYmEV3tpWiywgQPpdAu99HL7nWIDv2U
BdgN8W5IROB8u3uXpZrXbwAX08qQlr5sryGQU7ZK3QhXcppdOVIdBXp9dYxf
iPIEHejhrMC9Gy5QPJjU5fD9b6QvALFr6EdxYgMbJkhVI6cGh6vUjUmXFz+m
QrymhCWsqpq4szZsn3W1Ymx4T3OX2Z5eelQ3t5vX0/5U2qGWKluYoENJ1pYG
dL6lDhF6m53BKMN1DCUp+zx3cmJFTO1U0nav/Kvw5wAhW+k6svTWP+DbhV3H
77UDF3T+2TbmWdbNycFL/tcxKxZHQZCJUjyZyE+2OasDEThKJTwdRCO5K0SI
rKe2JRfnQv6FFlFMCWOgRwr0vykb8RQOQnYMoapl8Z4W/g/cXaJaHOTBKdix
tWTSVAZuLXzOZcZS5pk5DAFMvNSHLeRYsB6cSXduulhWT8yDkzgh311MnMhV
pVLi/SwluVgqfvqDh9ZitzGh4VOqo931W3StYgaV1T9U94gfX1sU3Iu+oSrY
WwrMAEVTNgvuDhzw6iNqF4auQ3JS8+tVqUTWHbs7RSlmJ0zMV6lojKLBmZdQ
OwLReYi/TaZp/r+YiifV5Wo08jCEECIz+5Z/T/mlWOZ9tNkoxYe5nJrYLhV+
/SQWM8Hgx02uPz8TYeMU+p6vc5F7373VpFYTvGUNUyR5uJzxGQmFDtT65Kpx
l8VZkUbXJCtBaqxk0OiB/IpYmmOCGlcfYgvq/ybq0Cmse2u5nvrZ4lxq6a89
k5YNVt/jEvKvSkFM7OMAHEzeXU4qeJrTsnxPILk2+3k7ki7EnS+gDg8zOGD/
p3pizDZXg6UxltI2jPe5QNNGuv3kR6nKrg5tc0szrQkvPyYgIYnahJx+9Llf
vZzhWGyreJAY2DSzRjkRDUS8cHUn87XqCwquw7dY2M1+Gv4hGqBLDVSVNv0X
gQKdiXpT5Fpaxx9zO0yB4sIO8jbeXOZPdw6MWNPWiTNI65sU5Y9esw0TUqQY
Gt3Sp/NRwMgzrYdjAf+IUHFulnooX3pt3CHfLB6jg3t18IT75WWl0hNUfnSx
u1DwPfUlYu20Gs313qLDmagdhjYg2SSDcGsqB1Jy+1hsiFRD06CNDXYib58m
DPwVMZ/L1wS2sRlwwCOC78S0+fj7FZ4KGUk5CqFWS5PV4Kf/Jown19rDo/j2
FpCPgc3GOt8NNjTAF/oyug8joOuFDNXJKEGA+WzFno8VIRZxFn1iPqzxYxlr
A0XGkxWoIfEUfI+cHBXc+NBqf9F/mfXA7tDUB6idFT+Sfrnfso0DdvrRaImG
tkKrl/HR9VDQHnzjW2udpRTu/OLMjA9FAOA8WkOuRa7jYC+5fOoOE+HYzLFU
/uLLLlTJQEzaFvkDNF3JzeqQyLCabVUwtC2HW48gyd8waA9l0xtQfntWSi5M
+bCLKv804q40oNdrIdpGJipodFcT2LpetM0ytSvOw1WTy5ZsbNAn4R/t3EWR
0E6lupz3WlvDPENRWO2hcRFIAqf4wIlJuYSb0Nq6xTOA2gJhh6rJdx5ifmRm
w3IWlSis/nM3w0IwHnjlz9FItQADsFytBGR2LOP0YS2S48jaMj7LwgKX8RDr
4KqqNPCgLKlLhvgVqjyz2MRUVf5S5p0Qea3so8UIU70+wJmIW1ImLSOnR/Cq
44jaiLj3tSmlLg/QHz1Mnm4D8OzTm7TigvcrLfLRslPhy6v8v/EXdw4h0oGa
249tFIdJIKpCb469oeWv5EWjJJ8ngV+/G02NnByDxaHItUupx2PYoQLiyw29
LLUyYCdPwVWCE0r66nWyikzCxEuJdxnw51esSmEkDSZB+Hrl+y5xdRAE5YPi
4eqG5dDIP12UkHkNYwWcfgtXvHtIhovF0PACF8fyVU260WIwr5kX/KRNGwys
ECTBZlFIvygFgBqIL4ZOpnklDUKroeGwU4QrSgtzhQssiKKskCs+6wKnfUx1
sHemkIZMsBHJoWHgXYD/D1o0mt4j+zBBt80+AzKjJ+9IK/qMiFgy9tKUcfll
2wcUqea5zlg5ILdV7+Mi+1itmfrkoTKbryhrTSnj+SKnILQJo3ekN1DwS6la
G8jKMcuNMSFPAAFt+g9s0YEFBtgaAustT9JML8+3Z6AeNGmvF5eYK7DN5FaL
Dbw/gJXWIRl/IJj6O9Dr4I7ICdYl5dOVmR8c89qJ1+1hLM6dIhUohSm8BQEd
na0FGMOmF0uetwXvgF26GsQzBrH7fazPZjN1/++9bJlEin6TJx6rNId/FBNl
Mr33n16oR6gmNY+fZFS74DTFcZ08nTWjH+ngXb5BFiyjmR+J6+Awk0Efolki
mo2tgIKJqhmv1mRJdS+WSpRcvIOYG9zIhQ1iv6isJixAvkQ1CCbO1UUUpChK
JrLPey6t9rf3byIrg+iT15LVYO399VYfuKcX7IavbBBdqnih3fJhasDzC9N1
jOhGm7tbXMS9wjMV/DMucGVFN/RPPych3Q3nSKCcLgo6PFRjo0fA4SdtujkG
2TeHOsjX37juYHYMMikOxURMMxawlNe2A1mX8OoLqLnD1UH3KovM91QCsFSB
4rCzPcMSUFWLHIcWMIbD68ObQJMOtZCClWR9+TxB7E0ufvoWmHBbvBu72cRU
HUsBIMqcdgSftY8vIXaQxO31YdAhSfTBshfdfcYNW/RplekemRaRu2TK40Wy
/M45H2wT/z/TIKD2sCJCanBL7IZbE5eAeW/K/8qpm0j9wZUM2uLon81w2R6i
TblAtZjFoRLst7i9MXUMxzrL/jAzzQPg/2dIWYxSrRnQNchmOAfqx8hkSsJh
wods8swSodv6mmCd6b9tQ+SfbPcgd0XeXvwYTNr6hLLvW4n7FMu4exPDNbqy
K9fms4ye0oreG92qUJfHkoUrURnPPrz6tSwoLflPnvg3GfvVUXOGuJ81ucRx
or80pJgU20fBTAnnCsReAsW4SZjaNGaQWmpT4cAzxNB6hoa9Ns3ewdUNjuQ0
rD4BQ2Y+TXgYYEbh9WG3XI7YTvVYrS2EE/6H6uFoAMx0NKD2eFeTirGoHjJa
wj1R+R2YUAgE52O185UIirkJ2ldp0EsI3xkhlr+FPCBFYqkFjtdZb5XB1aS8
qemfQdQ73O4oAiiRSpe9lDHJnMvEJT0/zDgsB/hSeAHRiC4W/RyHlF32i5F/
TRtas+2Bt8PFUPyPCbeUR9tsrILIzGrBdZ4qokAvqMHJBVWPi+DFETV7pFKu
1Dzt/DPHgxTaczSMOc9QgV+nrQ7o9aDQ0QNBDNat3dTjIHkOqw3iNx5SRnrw
rY0+KbjHq4J5WysSkuoMJcnZb/1md2gmxzCrtBOqbgZUNYRjrTvc/pP78VUr
5ABUfd1uWN1UoIenv5OsJRI1X58LMQ1XAn9PyTXH+hKVL+25g+XtnrNz59sb
pdYLhxZUhMpXrIrW+3lQnBmk+1pV76GeUIWaA3G25/c7SvtdJvitAu4ObhFr
mklK6PTy5Ug4kp6O4Jr0ibjZm0hs/oV4mg8BC23MC36PNC7lk2lzXnJ0sOKj
O77UYo1En9ysGf8WFrhOIXD7oTJR7eyTcAcz1zHm64WQVtToy0iyeh7CEPMo
q3jenCqpeHqeDyIUEsZvPqh0u2RF8ihpZB7VLlS+U8bi0MiXyZm/SyfQgO/y
UiuJTAUYmGEZ0M6N7gzUHmCnUlkQrNfxDe/cGZygBDEPaVkmeOgXuW8njVgd
jSlckc1gFQTh8BZWiihuezss8t6cVIA6K3NYhOFdmX6K+iu+RhTUG3VoWygo
hMV62x6Jr6vRBq+YOy/BECC3EuRLHt9bcAeKLwfsXFF2QGcVSPuFm7BqF7Ut
6xNAbcpTDbpd32tKMJ40HzFK7Ze3x0B3NM2CJtxf7z6IC1u2Ija5zFrMw+SU
AcTlwCZZY+9ihZCKjDlm0P3xNsE+qHvCxL87OONg+LF+ag8pSGl8SChKQ+i5
01pPM+tvJmn3B2+Z8srdq6YdOBQplox7C95kYkvJ8rGw3ph2xIy0SqrcV6kz
K9vfKXM69s3g8RkyZCCt7giWfpNa2XEwS9lR+1ZWWRu0cCJf08rZsLgW2q6g
7kZMw6wmjxz5/cWRGBEVYxjDI5MajqimSUmx0FHMLvJ6ABgos6R7LDqjoEhz
oOQJGthZkezfnccAx0/Rk6dg1wGwfRADw/YTkPAschKLIjhvhauOA2zalsiP
I96v1q5WbftT4UNVKvICIDekm3FbhCeiMohMkxjIV3AfPrj9Vsf9Wj97RD16
QMtU9dIqL7Ie2Ljkjo9P8QAw/7yodFxBJHREYLzPiW2Tc268QX/M6jTxppzT
EQLZkw17S12GkDhn3r4j+r5qdiQQRsnNfXVyvWiCDDiMdKlPtfUHNMtysHFl
IGn6j2MK6X+fFsBcAC74O99cxu893VX8Mfdd6ewy3EeQZID4cec4iGXpPhaN
4sxhfq5Kfxjao6+/pjcIeV093AN0BAcWJ20l445lIXogZ8r2Fkw3fQEWvzhL
OIL19ZXEKdUHnKhRe+rhhVWDEHqTmH/+DuIEfNUe87lDwU0yeGlNlUenr1Nw
QNwj0+5niyPwlxh16eGgX+ucqzJgceqwlxzol9UMTqPf+2+etleUO8YmzSiS
tis0qisuDhDxFWptS3t3KAGqpaIaUAw8UkP/UlMSy/FAaViMJ3NV22C4MCWh
03Z8ThN+GEsaV+iwPAAdsZBvm7qLfpNYDZ5KEV9n2dui+krbXCu/wpCQKnbl
fe8AtNXYReB8MnnGMLdK2u+KGcwx9bEPG05Z1vFsRFOcoivB+i/sbhQm57de
KrHJv0+zjejursgMhWZpnyos4W2SU68sfj2HqOAD9Lm4Yhp+XM2ZmZEy0Ybe
2MV+l1YAMLYH6FFyNaBeiyxvQnsybXQ8gZ0AoKmEt2/58Fn0ccVYN5iDxnWL
YD9c6DbKaYN4OMKMmgC40pj88++AAVZ6TNVZfQzyJw3lhr34M41jClaEOMAc
rMx0MLyQ1Al9xxmrXGCveLtRFLm0r0Cemc70DKD074KSOXU04gHFg4bgCfsk
hfZ4jQAChUVhqSTONk6xOadz8J7C6BtVvIkgnj4G2NUrVtzsWVTlszA6WH2U
SwCS7VMIRE1Rel2LkxPl1xC4f9nZxOByV5LFnQx4/9SgWZV85AiROsYvRmeu
2hiAll2qkvviK9Bc/VYNUZEyDYA2GxXQiTSrJLNcWwrP1KiMZHIdcakOrwQ3
Dh7yeLmwfjjpG8X6wx4rH/YJUiFpKHrZVo4pyATV8urKYN05ZZUvoFqLNmy8
X/Cl7VvSejq/7SNEsALH2cavmFmSb3FW9ObKsoH3a3pAcP6KdaC6RmQ3wULX
44fhEqRtZWeJFAQtFX+nhEUmIT+PTOmhB/BYxSZwBXSbiPexOo/p3Uyhoqee
1QpQXrmSFAtFJIcdvllblZ03D/meVYxEwZp3H5mztV+CHybsuV5hHK+Dq/gS
gm4G/I3uYvnB7lA1YJs+BQi8MElXZWgX5EF4jzuGpXN38gzdVVl66cRgMJ/5
LeWIt6m6QQJ1g9tuVEsBvOWvt24kd4UXTn1/T2Rnfwt7JrHqkoiyQ5jDTKIT
spkLWPFxyKcoxk1EN/s4YtvwQ7YOdui1Hw/uLC8zMInNJLCpavsWJMS8qJ/e
phtXMVsPdl+/Uz2DxaQctr/rivjThE8FRt25AoVPAWEnWSOG091WpNsnWpj4
fnGbpt40dg9dIG5mOUbEYO5fWLltRrKShqcehirlLFJ7GK55unj2f3tc6YyT
WG21SxCaUaGhdK7GJIv8HOd55BItUL5Ik4aSCkStaJkggqtXGPjcbc4WXuRy
M+Xj2O2UowtqmBqKWuOtzNxQJ3J9K0AB1zikgKUJuq6jYJpkJB8QL5aFHCZ9
/okzdMoFHakNbFDi4TJ5kw9LWH6yEf93g8+tDepj7TrHqjF5TRr2KzaEAmzy
la4k8yq+u3cBjyYMB0nPE93IBp2/TMVkhzJy3n5+7LbA3KfA3rkXuwBDbihH
lTI8DJl+LPf3I1DW47LZaDPNXFK04t4w/cK6BmvVAMUOSUUbpDB4ywNmJfNX
ZvMnnwmHxccP2uYNghZk8yEbqmQArt5+a0TKTFYhD0wG++BRls7OVp/pdZkV
PVBiZAu80y/BqTrqVxeJSf2f64RXrsyCDwAaJsYwE9tlOsClJYQE19ZMJ+Ht
O4GIlWBSFs2jZrQeI8nhqluzi8bdQ4Tfc0vmWyq2ybsDmSBhyEP8CSmJ+Tt+
9o5u4r9B91OfOKf4534ldLAVhDfpJJ+6sedJIhPT++JlXIBRMuPREx9AbOBl
s+uDjtz4qzLOJs8pTwkzV6T7vse9xKwaowhtaLDlXQhnXqoQJTCzAmTtI1U/
bKdTJlJYtpTOKImji4TC7QzYo7S4xcX4ZPtkPRcgGa65VcO4w4CdMEueoVoa
r21qTnG3EGBtM0D6EP1uTT6N4E+8IMHNrJymDB4uJqFs1vH1a8rF4CM5zs2z
l9/oqyIbx87mtHcBcKDIQC4+2Pc07inZa2p7NpXucluDUMVghOuOStN1AVNi
ACQVWhzy//jTLbhwBtwStr4AwD+A7QNs+ZOJHlqpbuMNA1kN4X4IY84LRJYv
TInNKMmTG/H4ztByrqU91NaMru+qyoz5gsSGUKEsVd0Xj91aAQM97MLulmEt
TdLVct+hOXcRYrCRf3t86U/jWnkFkvfpOW/qeh3/YFaV+ptR6fV+PoHJgAuf
IlPW57rDAFPA6JWxeuYpHCza/GP/2gOHlQIM1ZwS8bfwq1HzAs0UVLrSY1vI
Y6fKVswKeQdAopGwubaCw1i5XcKw8270y9WhWUtc2M1JvynLK4wizxDOu4dp
dxemkW7Q/D2FibwHz8rv66ozCjhNAPj3OJ15by+/zGoLUn0xWJ9XoX5rFUvI
DRCKT1vUw865p2VzyXUtUPAGeUtwm3Wcb7XZUfq81Y0ye4aDjQXMVY6l2sd2
S8fNS8YOcV1FRpWZvKdK0CWeEm+bu52XNFZDG0lyHNAvCKPehsbH8L27crxC
XPgjs3M1YSEkYoiTp3UhOOqVD/9D7fqku/MOJw0gvJ9XvbL8gMPlTMEbL4vg
wFyyd+aPRUF9DbTrSzAMTWUrfXTdmTdc95WF6E3+DT8v7aYBnSxoLCl8p9Ma
ZVFzA4ENpg4B3WNrVfl0gyk86hs2WDnI0KCgQ/FejfbMQ99XMevu4eUfbfqg
7t/2gk61sniHulOc6XiG+2ryC29GwVmuDY+FO7iGGfnyoUXc49LplxsvgWJZ
sf6bVaPo0QNiHkb7Nk2DK2WzTtRimU9bnzJh5/vkt1mSufXDDEuNWr5OqSfX
OGO0cS+MxM5N5uXUU9cEyt4uRZeSllXayXVeHXQNYF5fxXIJW7MOiZn7N9rU
MPNvqXnMso2+QhMoAHFvOsGQQmd8i2d2x+6H1kTcixplOH1wA2kOletNl3qO
20f8cyMeENnALlkJrzZQgjMXY9LP9Cfv23jPUADNJYA99KElTksNwwLzakXg
aW6o4ADnAaodpcZJjTQw+Uvxrto8ntOioGc7V6Ihwf90HOS3oNPC9CgYfENr
d5sFA2KrrJXGZZfVPoQ6uuj0ZZE/aThujcyZX5Ksp5MuBxwENpWcHXmuKrH1
qJ+/KNyAuN/nOecQoa3PIp/ugy8jXmm1xm84ELTYRbW2tTHHrOSacbJYIYYL
0yUUsO9M2mMHHKO9+g3ig+hndVEvLuZLZrxTaFB+ogUAXYVxJ0K7Xxv++ebx
hTPXM36z0hWn48SM+sNpUFaVEBrvzGC5xqPiv5Blt5vBODUi/v/TwxAsJZvO
rXJkLeTKJBEfq4Q+r4QmiM1HILl4ikZWEBYF2PsLADZty8zNv5tqYOt8U9wo
5oVoaZZ8oX9T/bDL+h7CTInHOcqbLCh5iX+T5aN2ZgnduRJIrK2EiIy074JK
uP1KvhTcSLuuk92n3dnG9d/ngeSg9jjJc74/MVBR888D2kOoMzKVUDpfmFC/
ldNp2BcHcHmdkWeITu4yzBn5xFBe8+MqJRKWJWET9HtvFW3fZTb30pqhGL/I
Z69W92HLEvQ/HdOdvxCgTRYrHG6RMkJV43kNoiQg0hSj1ZmcbY8N/aWSMyG4
gKGwp+U5tjJbyU9wXbvd+MuP0AJLw92VRxSK+e79NLmxIHl5QL6Xo104TUmn
L8Qp88oRVesAOngS3GQjwmLEhZSJ64Nof/9XyBiAFbSWGZJr9V21MnPKEsCB
9HuDBowaYd6gr2hTkFyHJSKCOtuA1RNNnPViD0rpAVRxGjOiD7Ikgdz3+PwF
l2GhEZHOcZsN5NS5ymW485uskI3DBlQ8MfU7z0qv18Ug/9hZmfc0gLHj8Rki
Z2Se1pRe2pN7YGKQObvVyXpkECT5cQyG4ACT9P2nlhwYlgVwvst2w0rIlgzA
lmIJmk3OnLQa6+wDNtsU7MxWsnrmw2qr0PG85NDibOjJ7A4IBinSQxpyvOFs
fNZDU0OFs93kfv0EZy7niulTSm2BsZ25kFxUhPgOrnKiEXU9jd7D6aRw8Qm/
9z6nnewDdXVZ9b8HRNSO2A4fVzpPMxZXMLXTES0DxCgv/OzAGrtu+iaH6DNt
WaPrmJooB5oHq2FewHcXQ6jipAMr7z3c5Tu4ptEPNocyDHUxhjE1nflxf6dB
4bXFMrFUUCCi0ccNTpgrHLXUVjR4z6nx0RHVmNKWoqBWwc2w8qgYs68GcyEE
CNYbJkwDmunwMmjDRnfiyg2Ig4UyZblQNhBXCzb8flf8S+VFwijGIaB/oMW4
mk+laT0JqXKmUg0lGQIsW9XGt12HM1vWGCt5xrj2NzpxRvIBna92UYocaChw
MZkyYbkTFYe0/bYYsCXUWGAK03GVDQVA3NvZBHZD9QwqxmFuVs9DzcPCySPv
Jw3tHLVRJNUTEvQnbOCk6T7dMIz5fjUMrtaiGu3ovRSMLwdVSboCNuGyhxXq
nJreMpeQq6mlnJoAzBzMgf3qXdNaJaxJe6Bu04lBseeUzErobtuM132T4hv6
vqTFMIVbpdUlrqHQH7IHKJZlw0lzCakVLmVAdDMcLpebd0FkV8Q8YUMXGz+w
3+LLDhuTsaChwsh8RVYMTgVUuS3Si4CwApp7DnoF0BZeHZlJGu2nO6SkbsSE
FJKndzfRCD/bh8ilVOP+paxHgVmkx0gHLDu1RkNfeeq/7rrMXOSjzTheDfB7
jQ5q9ErHFw0ZELV5ALRUu/oTihNUFp7Fvu40s6hhvRTgIeL0P0E3f+bHsIwX
uzJDPKuzFc4Rtgp348vrOsHjU8N83/FDts8lV3B7C0al9go4QfZk7PXTJCpM
J+VfBQjcRagKH5C/uBqREQc2S0U9rFGpB+lYMS8b/VlHNnhpxiBaj1rJZy3D
9/djhQgV0AgJxRnUi7i8l1iH5t5zsnq1ctbUoSJIov66m9YIm+pAwF1WMFKB
MlasnhUJsxDWkLvmnqE3AFsPVROy96NS8D6b9x8CSiht0PkWYLOmdje/3Yam
PZGoYzezLkarpJ4Edfq770CV5b0Jqe/3EKiHkpJNGXvTQXzM/Kh96YU3KSso
aStciDuRMI1j6zkpLYzz5KH1KILShkg+3xyra+cnuHpVfjSgS7BhlESnkWhX
IGOQSGvvC+cBL23tNOSHD/QdWcXdJoVq20ImmbdnRgn1smiRwWwdZ6uoyBUk
JtE08sZRHhtuwKQLn24yVlAkHGt7LHr9938yCHmmoXKeB0s0urkVSBX9vQwG
RGzgfuBerCPeju4JW5T8DwJyOQw9vFf3Nw+wPfNm3crMEhp0BG9K+QkI1gab
NKoubrvUU9J3CgyPQB8thH6cIEg/mpldeWzp/W890adlgdk5aFvkear41JmL
VPPoPGPi5jSaFiOQDuMbmtweXRzRBDfbNzR/OzCauNBCNvCuNraJMUz/Ww1U
vBmbYk6IbhOGoDIf4A90YC7UGej3V7D77yjAevn30l1AT7RbV0vqx7gLWw1H
EbiUfHNxac6Bkd/AqQsCYyKaovcTjoTd+Q41Vqyf6L+cq270oqqMOgbmAxcu
S45wG5x56Ajw8P6ovxCSx+3ZLQq9sRRhJBWWG4EAGi/8EDnDgaHy0mjpPB34
hsooudUoZCObhD+TP1ejM2nXUApgiNGxc5BXMtLPAbFLI4AjhcIJ0ybVC2YZ
HkRBuEXxDiBEG72CxAZr6zAwXbDUBh7WLa9mQoDpGDfaNwF8tNMkrQWS0gVW
hJ8PSrC0rorfefRpNAQuJTi8IQqCaBduzEUs6Tk6LciAKc7ypl7j2qFvxpYt
7GOZ9HNxwdWNbonjokbQ1Zm7+TU4ABEcFTZx/XkrJV59O4fz1g/JZ20tQSX/
R1vd2h06I6tPQLki8rZD4DFcpT4igTfaqVXtTKJ+I6wm8DBKI49eGomnDxZY
QcwuJHz6W9ndrU65nPqBK1FibcyzG+c3gsTAM9CS4VUgUIQjvRZgqsynq6y4
53YdFgr6M+We61b9h5C1Mgq3aLX8uXad8SeLw7Z5VTEJIsNNEVKee+5bQpC5
uUohv1SzmGh256B+I6ukALuRSTB3pbXK69XNSOqt/izJkd7KxPk7kbevwl+V
f0hRkBGQSXvZa4PU+I5yMsSoIB2NLTabzATvSYW65iscENMSbS+wxWjRrKSm
vX51QEswJiDKsIoVQXccVH+umpoGZXzhGgJq6FgBem/8ksuQ2vNgm0W/DNbS
xVBZmuHbNHK0XKkE8QMJTjhCFxYJYCjy68k8k9l7fiQ3626AmfaDK0yyozsd
iLSgKWx5CF+pGAuuTuhCWFUdQgmM/F/Nx6KjXEjkMXrM8A8GVAiZHrBMInV6
z3mZDQSjq9npDMFxjWtCt6NMxfoHef42f3pMbQuZwnp5zuYfuQkc8ihkgxJl
QcOykdFgrWPmBG+8KleJ5/de+1QJT/eejQHC4JiOdzlkEOXA9f26TGhA/HZX
XqzQ4j2Vp9pfSFFGB0MTwD1CsFkOjkwnDwEBsBpYgzIAu7XKgBsK2ZcklHKO
LZap9ch3J0EWeukuyLerWFsDEqHqTanRvGGUeJSEJMpnUdN3Zk3QYTIrbCps
B10p5iwgINxXKYynqxpGKodLYrExDUPMLyW6Tosxb7uv988UEABOLIA6lAYe
4RYny591s1Xp0QF2ZUVSX/lS4VYJQaEDgwUqvi5fMK5NGF6SFXobeClhXv/F
z1QJodyHCu/q5UeCWTWnG83LftCjkZYqtJB+dsSKltP82k/4sMUhHkoZntIK
EZN6Wk0TRLwdq0pA/Y/Thq9Bw3wDZm0rCWmNDT+f1bnuSTx43Vp+G2vRgs4R
PU2S47ReRtNbtM6fsaiDa6Qu5iGW1XOgcsXM4gW7u3EKPeqkjFuVM9qmJu08
NzMu3BVpy9hX0MgEYUTlCMRY4XZpq0XJA7H9V4FzgCug/FtrbhkYb175CuK8
xCLkTvrvjJPtucrq2LkitrOJWXdNQZgNn6PDyrV4t6rUZtq4L3qCdmo2GZV1
qfrqHdGJHWmK4BgP9PX3zskxFZrbDOxCwaJgUb/k62vVxCD8HPNrvLaxAsmX
HVL0a4TnZmgS7w0MhVpruYWQI7htSEge1g39MQT3nTJhRPSTrQT+5IclMGgZ
Ks1DugTmE6npdX4S2I0Q4Qv8BTmtk12L7R+z4UcLUdaCw8DdblVOIqIMzQNq
EojaYSGIT5X4GJ9qXM9SUG8cmSWr4jH+92A6kKUzEB6+swd4eAt0R9zqCnsk
PIxP+b0qzYwvATaOkEuhu+dV8qNcdqTtd1GIcfFtznqWgGskIWIvl48R4sCY
DVG3JQFaqHKTvEBVELfe1iUH9gKUSZF5OTZutkfz2hemwcZMrzRVIhh5jqfM
Lby6rTEKFpg++ndie1AadMcJTko+FPunSLXET2o9Awx27i2tPPSfC4WamX7q
e+iHzp20itiGuoIZMvUKV/mdas/gWvfh5yDMx/WTVTXtVRFkJVkCZG61+DHb
JHFurDyLlbgs9EvUXsOohpCFWi+VkuDRz0Cra+apS9YXLnOkqP1/n0HF1yTC
ow8F4AKGgt2Mj50zssQpKP/BkqCkaPQE5e6KCzPIqwaIXUa9AzKTmN3xZI9Z
ei8CmLHbmh6dJ/8N8jqp7RcfvMCtNdzHXIaKuCKsseGAWcPX+pxmnrJCF20k
Y5nIoQjwup3BzwTV8R93gCPpilwBpSQYeO3kiJJ2auqOGc5zEokwY0x763xO
OAzbC9jGtV+YwxFu99SHkKoX4Ik+BILf6z3PLP4fkgQASKddzJeQbFV7UskW
1+gXxVhcuh6PbF9HD+z3PxuR5QXpA4wEizDw7nlY4WqVbSgwbMLssfs0urml
qeCJxO+uIHbF40akN2+7j8tU2+gc+GqkjStx/T7WVn5TzYWLOE2Gpb96gUEz
yVo2fpHNdGZ2x+/bTuLxifqpu/86aH4f754qwNrS4HBq9XSpUWTDvUe9RxRJ
+qZGDqyRygQ1XfiGD03zg5xjFeAPEEbs5OlIBvtiPxS0GRoE9yeK6hQuikIP
nrrfNoQp94XT15DN51B5DSu41w5eZJHS0AmfH8uBGF4UjBT5/jPUmaoGM3Zi
oLaFuBcRGPvIC0QwoNFbPpocyB5H/fbqC+TOjvJeWG8JDdVzYMEKcZgKyPSX
EZOcNssbqqovpUytyJJnLo2x5rDVYRDhN8o/Yt5DI+dzr7xQn969eyMpOJqW
tKkzu0JWpMv5g74LpLADXBrze1bIA3oQpCraCcuROSHuS5m4Tp/Ko94JTmrk
QJGCxoqPLrOrfj/do7kaUChCNUORRdvXqzr4pp0IND7a+wVqqVXIR91Fp6BP
MVGBfGCD5sXH6XVAGXlmadrqh+jdle9awd8rshNPJrcbmpCv/9aXN3hsN/Xi
ArjzwEXxQjLuhV9xIVtGczo5XVjvlquU0vggVozzLS1sPGgstBmh8RKU/gGL
Pgt7dYEbiK2LP0gAGmTv38BDoyOPIX/FIJ8msxqqPpBsEZNd8iP0lyjDhF5f
FqEEVUtpVzKk2AnhH0U1lkw9vWUSqqozS1J5WDeQIKN+g0RPZDtUAqpcTK1w
npIVgyABYNuyNrK8PqdtE4ERa6JemS8qCNfNWVY/wwqnByJhuSwjsOT7YwDW
0uyW3ONEzC9bE41nTxbeJYbiPel7yT615GV16aAUMD3uRNZusQsWLh3gZEoA
VqL3DDwcm3GX76CD2e3wC5qLnzlJ7SmDPomi914pQ9FRGVlq8SsmcVKWSnw0
tT6NQrj4sWFgKihKsOZvOrPRHv8SwqDEX8G+HDBW0YfzVHezL32bJ9g7E1bu
vK+boKSRhuKf6ZtJRaygRGXov0Plhb+SbjhqhJEDaCywaSY4QxYS+RqxrzUU
EBEDoXR6F84enZpN85ctYzEJKRiAuggCE1CSWFg4q2Qk8PtDtnWk4wSa7EtG
4CPLPfqucOsK4muyor0xjLq7gItvELW3sZIQ3ZBwrG1df3xCIg4sCW0KBhln
J15v7+GXFUGdXSzxUVN4qVr6iDpGYlC352/X4j+S+6JVP/bkuhgWi5T+Z6w2
GP49d7jZTERS59Q7K+0J0V948i2+KY5BgOtTlbI2jtWWiY75gVGLeitmjo5d
zluoMIv0aTYMEbT/gnyoSssGi+iB6KOD/ZF+cLnU0XrUcHzF/8qTBnRGx0ri
Tw9mGWK9KQeRz/I8FgT831I/ivXqrSk2AqWUjjYY2YhaKPe1Ziy10ZdjVX7h
rlvZHn1/IebecaP1svqQ6mt+uLc+aC2eMtRl3wIBWkRmDrdzMRr4UnJWqEYc
ft7DI1wBmv5S4DdAyMkiftZNcg8EEP6MuUvCP9K/udKxY7LasCCGJ635IUZG
tCS30jHvTCGEVkdpFyBVXLthjNosWypQL0CVrRSw88m4raKxR5jPxBDyKZqy
Ct50O+H2k6pasrfbl3GUtyZrYjsNXMsCa5UKW4P93OM5vaD42LOfgofo8NI5
xxILmanZc/o5WY3ThRKWBrVCR3vQCBB6yYGAS5Cgs96DrdmNrgTPjx+2vz4k
HZQk8nFOHDieK3ywJ9i5DgBe3Y8sY7idZFRzXdpqucqnCpl9ECQJAcpVP7Mc
r1dvQuv5intLByseWOQM03bjdjHVDsOmkxqqyyqeIZrH+vmOkHS8RMbW1Naz
Z8hTEYT+jSCGHefWYSdfnOr1MUr02Prtk1ts3ADbJH9gAZR7aPUYjVu2YjH0
DM8grN99JXPdtvnKCF8sapi8Mru5qze7/VLWlHMORw7Xw91xKfxd1cb1EKza
Qj2t3xavoM0VXprYNG/kuMyzJ2FAt9wmAw0Ra8KvgewSOc0vf9hs7VOTLXTO
0ttlHM85iIFijvYwwmSZwMtVCohPDYhKADT0P+IWIVbNFt/QswbGF4QRLHvN
gQdXkLrVYP37KPUrLdoX3Oy26dljAQNXvn2mr/LL0uJAkX3Sf0SwKwtuirLU
UVbYI2dxkZBR+0f4E2PuWGYKxHgB7zA9AZEUo2Z8aV8jFFFoEszpfbTW2pr4
fMfCRKJOZ47HZAQ+SQDI9qyxWYOLNURITu9+aHlWDJ5Jn02NDoP4tRugreeH
E5siD3q7idvekD5aAQacj/rUFDT4aJq01S2pNPygrt8fml9ymxawxgyAlX2x
Jupdi0pr3Ugk0JDnE45CnNF3Izh9lDz/dwSJReQoHCJQFzYpddKT1YQxsDUk
HR6M0JJ+HoV011D4+2sT31H1+72x/+2P68oliJYmmeseohh98Vz/agJLUrys
kmuR6xtzl14rF9j19GbtyyMzMa+PKIsAtwNICgz1Oj15B3DEuuy2KCLs2iKJ
QTYxAhOHf8817NYmNLFD+7Lpw02i5MzEuTGd+U8wATLLAQh5ojLai1vBKoQp
ed0P9ilQr3YzgiHUFdAnZlfWQEjD4oatCC43/XxKcg7OCG3nVBn77bcrFAA2
u6FzTydOSkho0hSBDI0c0HRlAFVbXNB081+qZhlL43dcdGiOCaq793AcOE7N
H4SsveX7yqWQUjP76w9XyTxL0ipEjXdK/48NBJCXutN65T6a8p8oDQhxTOcW
HEV10Bq+rtJNqGNldQfsFBYyQV+4y3z/qVG7Q9a/kfUXlhX1vz7TuWSI1l8O
xhOT9t8Yms2Tdt+iXOwbNJVl+wn4JJeB3aN/XZzuivsulG0lztSVu1ePs4zW
8eIz5yR2v2dE9yu+nLw821py9OC8rFU6dUuul2e9M2JHI6NqDXBu6TKeQvfj
covzfTRZKg7Y2KKxQwy0NUwpre1DuzMT0g74FjrQbGT3WmgmfZ059b7MZMU1
diiW//avRC9TSqdDYDvBYYGmOnhzH+aGkdz54rAS6h5U8pOCN61DbJpMDvn/
DEo3SppTiXNGWYnN1GR51AiIOqMvYd8K82QHnHDG5pfhGtI1WEyf6cGem44W
bqtyP4G8Os7VlB/zEB/oe5IJCkzhp2mTP1XP8jKkE3aeXaBv0jRc/ruOZF1p
gsqLElgOZOQtgYA46VPJIiEIF20qs9p31QTKBAq7uXNYGFzdlqfZY3mgmwMI
/PrUJibLDWd2dxw5iIP0Y6ojt0X3w78PLIDM1u0vRmautpJMLyzD/1AxBxcu
qO60zIKKcD5O7hg8km9Pv7eTKbErJPkHKIP6g/iaqbbTHPrkU/1XhqMXx5Db
sXzmgNxptEZX/SRi9tFqlCc5WZmcdXWRPITlYgTyKYQDKk3y0R8anpPVPJ0p
cygefPXz/P/5sKj5iUaFNa88U5ahO8RgzWsBCiI+A+Tjvtf7tmVIWwNnhaYP
KIMgZy1dFjXVe5bTOMoovmtQmffFO8p7bX1bEj8oQLU+CQNrxblTzR7IhG7H
UKygqMfPL0Aw3UuuA7wttJvpEhGHZIMO8Z1pDjwekcZK3EL+ZP8125qzi8yN
kyQsW3Bn6c6HatGywdLk1TosK4Xm1ck8T6f2sux/1nJrW8LQp1Z6Rgyytz6b
J5t8I6fWSq2fzMPUEXSISRqjMpN1gBMKo8kxwlOT6cYz+OAELy8OcFB5YsEI
gHkCrxMp2qqLo+KtFG/jj6Nzl/kLxUBINKlmOU/c4AozfmRD0wMGsCvpsr06
bwpu2GuGXZg5ieS1G2Yn94e4ALG8iLhYX4XgWAMd6HeeWbDxBpDcvBswoVSh
RZs7ezaPrE4E+U9pefDtXnBeMqFhl9jhXe0rq7kQpCSHs9i6sltKQ/AywRzB
xGRJI7bzNvPZfI0aJBsjgBL1AEmCLDX3MwvNUa63MajlMUYfRC3KSShJfXbI
0RKV/PbJBLzIQ3Yz30gZU/AYeOKKrR8+bjEx/iVt4Br9wig2iSLblhmiSk/m
DuQ3XlF3ojOGu4jXmBmP/qClDTXE4n2CeK0afH9f5Dg2+ezrWM9UPVn+f42i
royTIKoKtHStZ6ByuL9QLw25hXS3tBGHuTH0tmmDF68J5kUMKi7pS0eDzYSZ
HvRqyhGRPcGRFw8aSFFPvXxv+hHlNHN09H65RLljaPq1gjWnK+kNwepNFaPm
o9XHaqe8Z851kjGUhvEK+d9g8RZtUUbg3q+RwfcjlXK+Woq1fUMGajAsWJM6
OPrrWe1rJNF77WeolzHol88cODJK1+Y/NPGu0xuA1t+6WAoReWqAv1auMrFf
H9O6Gs9TacKjwdXArU3CXh6dyZg7MuZubuoS6LF0Z13pHJRDxV5u33QItqxl
FO2kBBkdxZ1FZl7pfEdjC8QbIo7WN1W/aybAgy/inUC5EPvFCL2mEQZjoSmj
xdroaNvEczfY8lPSKsNMYRcNytEtQEbaaXZP2+MipyzKbDoYO5Z8XtMqEt5j
91U1Ef7iMKyC3tHkj4sWQ8+pEXJrpnOVmV1JEXoNbK5l697BgTwzQEMk5paC
XpiFFFsH7tGd+Afq039DLhoLQ7b9GrmDz6X6WecLGB71TymAlW85qKZ89j6l
73BWenlq6Us3Heeg0L0yjAIkVhMUvkiFQapXBGS2p6nsO94SaqjB37MO87pI
mv2j4mSXyR63LZ0XLoaDUKxwJIVw63dwXvIyPZW2q7V04145cDeV806WkpG+
sxzxTZg1sSK5ZDJLT/y8QkPk0jEgXtubGA4qpBkxwfcRxp99IYZ8wlYR4kfa
ciVFgIkQggL2suse/+K+pMEbOTjlODatHVO0u0bmZue0mOW53+17R2Pf8V2X
sQGjlbDEvBsLuUL01qBLKAQNiov6CIniJqkMu/C5Snj5JAyaUDf0+2y4mOhT
btec++hnFcExYwtsK+0XN2B5XibZ5S2/zM/1NCXPmvs1FumxZAX0pOJNRaHs
RZLC8HxkW2GOLQkUc10T3wl7fwLDanWGC5zvRxDsBl1jGS8f0VB/ZPaM8iF8
P/Ofbu4zppJUK2N7jTWsTwP2EpNHBXVAC5ogdZn63Flu4znBgIc0+zZg0LAK
er5VotuN9TI+5LxP5UZLgFPjpO0haGhrW4IyFG1kvuuWvVPnB0wPFpz0lbuX
Q+NfdR8U1u+OneSeRcfqKlk93wreiteL0OVtdjbbSMN25tU4f4m6UzgnVDzO
aTGubhW5cSlTzcKE77QIz+TUHzm2lMIV/41p6C/vjA6ePUOHCoL4+KPaBmYx
nON0x8mlsMnXSVJ2Aq9gYHk3NTmQb/ELmUTUI1HglgLEpPszX/HCuxEyxHiM
xC8Ra6pkVcmpZKu5NRmhYB+T5PZRvoibkyp6+vGfXc0LKAjrt7PHAV+6pXNe
fxDlcUEi0g9rlLaRsJuF9qrI/V9utJVcMzvX8wuiGynfRwgagWZL3kDyavgh
ieTs9MPTtsPIihYYOw5sfraUHeKOK9ZYeQqQ9LqjeHFMjhxFwDhUbU3ez09+
lGgNzUHlbP/KBr38w0iUumT8/3iz1/9UdrMiZ8AIUBFfWLvQl4Q7cu0NZ3h7
3RDdG/pogfg62uRF1PJ/8dks5sVsd5x7wLF3yTuAH76tyUK8z9qwQCVrujgZ
Df+atOqHplzP0gNqovBTpQED+I+7Gm6H/uym4mAPkfrdA42qP2ZVBmJLnuET
7k/6FDH/jRSQpzGY2TZk1DlTj14uzgsCXk02sO+h9x1jP3sy1MgMZMgyLSx9
iuz2T3993V/1pQv6CEkgrW5nRdHwqG00haQ4ZA2QFD7HGGArIdt57xJK5tCd
eERKbfHLdmTzf9oV8dFtwFzeTbOG/OfHFo7GffahguMo/D9Q8Vqn0sqdzJ0u
SiZsN3EXnrDHSlMuDQh+Lab5PsJVNXthK6oVuIyLFcefsy+FXnosKqkVqfK4
HXKti+S/pyfa4h5WbEOfUtX3zTL7uGtfcmvJJCmGO4vkVFoSChOUYctbD9CC
Ubxik5PzbgpVjGTXB48KW0Yk5h/J3nHOd4AO8dAKvyRp98Tm+2iZhtVvUi6u
kbmZvVI67klSAaPA3nIHERiGcqsU+536Z5GgtyOq+G9E/QY9fNwkO7kbRlC0
gdoOcXrdsO/wBQOHnPbrRpJ9c7hTvHUA3HS3EXFKQWjx6x4yeR47OvMkCyQo
mx+PP4nBAXrD1EQy0Y5mWyK28M5fBnGi4ElYtsot8Tjdx5uCr5L9EAFjE0Wa
Xfv0XulVUCWZwG+cXzYZU6qQxLq8kMZ3JAEruTrnnKb1BlBZLFEzwyE1gUwk
q1ZridJGchKtHkE7iITO5Ni386+B5PXzWVofGbHaLe7ko1ZbRn5kHKdWuFGa
ZfkhMWEx2sF3txgg9JVkHHl9ifi/Cp/VGcn9QpEGfOyiQtkleL2icEssRbr9
UBRamD67Ny/cHqHzT4l9DiNfAv9TsOszOAhThH+UQYoxvMGQrnzkujyr+PdH
YpjvtC4iCCL8tq7qA4Ls0J2KAIN5UcL9bN3UdehBQo1b1b2aaVsLLK8VXh+q
Lqx2Rf3+wV9GK9+7B66t3yFv1/cPbITwD1/yOV3su22QqRAZJhN1bvuMdGyo
DNN5zgr/iYQoSRrjDUAPVLgGbMUI0t4xnB/nHuPIpPeOJryBCkafAoLoUo/H
/NB/csDY8UFBNe2tdQ9nrM8FY3KBc0pr6Knz4vBra3HN1mNC5lLQR+m/o9CR
RbLbMfcyRTr6H1ROcXO4mjFlfsT4MbokYxFQjxQ6SVW9Ivea+5eDH6la7p+2
BasrFS1Rt476fi0hoOZMyjOGP4t/oGfjCMn4uG841h+CI4A0d32QKMW8VUFg
R9fzfnDZrsHbncdXEnpZi9bgJ+nJylcCBm6A6EP1ci+gtZ1ypi0dKHDNATQB
x5mxftZfyEWQBY2fBKrwacCD1mfmmtIe/yNl7/ah4EMUls4NWQmzBtNauruo
HPTZDOGlBW3WurpkdqaLGPBWV0m67X2fxxP3+1ZaklO3/+gcWwBIoXOy6iQB
Yty7UUUPGuclyHLdebWWxPvHT4Gd2nwWIqHuw8CGLFN0oeblg6Ttd7UbbRuR
9dil5SgSFAZzpPlDBI/BMXbNjFDXvZxQOOYxOIMd4eaPwJuAjLlpeSrYOYIX
RmJLIepkLSozcCb6cF32HTl1EcHBv+W8ZvvQKmxEomalJ2feccTSiBWGGdEo
YoXs7iibr5nmSINtXLW9hxtcFl130qZIPQKDzkiXcnMUYN1lWNtnMcmU52th
G5W82TEGJBeuEF8iS94a8hx3w+ORAKMpol5M2Zp+YPCtjqKYXDw6yl+W9KD3
ReCXvjrAGxi9rMnv0bHbLZerEpgpnSAeGTrCcoCGvZvve4R5qciJ/bij+Nxv
1GKfbY9TEItxfZUBdV93eYDVIo6zDMYIKKP5jVRkFuhMnnd0ukAbGPFybrpi
1R6sMYD+ntNz80gebq4D6AhqqO/n1L07V3+WU8ZriAPorVJC/TsGgO5FELYX
0L76KCRm28jv6lxKiKqfSbMeZ2ZdEBHnMxP5Yug93Q9v28XY23UcvA2TuhxE
k08numjctaO17h54DGSdKFefnD/9tWHpLUgmwzBx8OK5Kl1VbUpuB8MBlRo4
j6ZnUId5ZlC3iEovmPId3tX0IVGJGfRFB8akj6CD+nYMOr3r+EnOgsfBsdfQ
ztcwv3TN0s8BsQPWSOfO+Oq/4l802Y1OA3Wc3P6HN1S8AYaNZPospwg+bkXE
6sZYnaoP5yJQ2mnYuFJ/RJNfEbL7HV+spQzmHWpE8mB6OhU96KAFuzu9M8v6
kB/TutWDrLF/9yg8QgWzSyRbxaawUXDkZCW3ACTmJaNobhiqrUDHN6NdLw9s
LwybIzDv5mhJIPX4DokNKq2tkbhtWoVZmUHQAEL3Sr+9+k9KZob+0qQ/zefR
jv/7F/32JnyC+FognijGJ9OiwwihL1Ov3O6kYh36xMGGEQOXSulm2zFJBZKz
wYJ69VJYZq3joME+xo+C+Fo45pzZcDU3Bm+8IRsPgzu0+USqmYjoy524AABS
+mYRs0p0UhSS/LPs91xScMbcpYCvOuQze7+s+oxZsU1sA4M8PbHFPvYQioj2
VUnM1PCXEeB2qm8KWID/3l4sm0BrDQ8PT+Kg+l2ZKh6WtN7ObOc9yiW64n64
P1FO/6ZMbrdjgUxX41cXH0qbFIfoo2Qt8WwJXmLbtd5jcKeXpMuBZW/HXP9E
CkAzL9v0rWNNFEfhXZ7f+oWcAwqm+JL1Klewmbpxe0naIzTz4C05Iubz1yJY
zmyEMSFpa8V+kdNvvo6m5k68cDxTayoKdtv/Sl7ht+0E9ObRZrAmbFDFiR1t
/vufGvFbBKcIzJ9QpN146zm2X5YwS8dZP8SkvRhTvlL7gJsIgU6EWdWtNLN6
yRCLvDqVucoAf+hH3K3euYHZkgpNBplY44dSoVPDdqE+5gXU5JjAW2tB6HMM
eovxxlsOJthiX94eFFIEPrBytWIlPnoBvbPFscZyjK+T0SuxpyEyUB8FuCXu
VoYf+CrQpUfMXaSQMwgT9ryTYEkVYSr0XJTyOMUOFwIvpfbGaCgdiiruc2m+
1BitnftwNpTPg94EjWk+gISJseHebDPmWuPy3531c4BbltnyJPr2VA5qTHiu
iFRD2+MDjcC3ZcCiEfE+3gqpxFdBxxBEhhgOjBqsLitjlmGKNLkzFsRG5y4I
k1N/nZCkrUL6Kh1gkIu1gmD7vM6DqiJQnuUMz0ad4bvnbQgNCoaNHQOgRle4
xbeCfZZYsjZdHZea3/x+5+nChIAff96F9FGrp5hMrEJUO0ssqhq61fXnM8RO
mkSRmmFmA8CckZWFanQIxPFlOsG/QZAuOtwujFvN+GJmdqrQ5ztNphT+pAhR
7jeF3pOsbrY/3asVZL4rl3pMJJB6qoNtdBFPIa4g9vltjXvv7TPTuGypqyB0
1ek9u10fzfxjKy894ObtQg100KEGMADxwI5MUSB3+zYBME8aOW0gSxGL0O9i
AQuAthseO+8B1bfJAAuPwrN7JuvmCxZm2kfW61HXKFDFa9SKe5BhC+V91pAn
RuLuxawZF/t+8QRBHzaCh0yxYK50SVanTt+KGas8KYOJ9X3dQYludmufpAXc
BmbMwTVf3zSiyr97mhmNhX32HbkArZLmSDxDNPOjxc8wHkXqu7hajGlMtqLx
AKt9SnLTyIMNDvt6ETZ5I6ibwqNWgaWA/x+1VZndeqP9uJFTlVE1PRi4yvbF
3/xrIoZSc/EmFUnG0YSOlo7NYNzJZz4SfEQR7nBQVgVoSCCldgGd6F8w2V0C
ecmphzHBAcxUMtcaOWcGhb/4mCGOHT90SS9mroRgnqlzo/rWFNOb/uIMK9kS
q91MP5t5ZJefI1Ri1f3+fx53Q+9pj0LTUVMx/vrGvh1H9gTSB5YdkVVCr1Fz
RbLSnf4DVlCjEeUKhj/Dt1ua7q4wW5Oe9TnKWBq7bt3dfoykAZqD/MlOqAh/
mcYfLRs6ptoYS5XbcFnBJRh+PL5eGz4xloDix/8NjYVwKtFy4f+OyP3xpS4E
lwMHvywu/cKZk+4LKGmNM/ozaCVsCrM8EIXfKnL6wjGCY1zb2Sib0Tb5GMXW
wfjr1cH4hLH5LxlXb3h6QbnlQJIAwF8246X86DDcYP+a84vI+PuaGXB0iRuy
RZuldMB7PaIDg7PR6SNGqTrx1bxeWrdeChROHPAD9OszFVxGv8EfsbBzgk/4
ht4TiIuUSjZ0NIBgRH/a0ESlwKcYJXyL7G0SueLBWfwPZ6kZHddQhBDdXzHY
RZEfpaoupWPAGyldXidRoxJhzZMggovtoEoQUMZqIU6Gx24rA56jmKO8Ijcb
Zvwc9v1PjuFo0QZ7VOF0DmUHUSN1zM0E7Wtd9YPsTnAyF3Du0T6kZ+FgwDX4
AbKU6fOGk2y2wIYXmjbllhZMwqOD/xS7wF5n2OLr2JdIcRkr1qhZ7Jdb0O6N
x6wN8ZbwbG/FVUdBTqPqx1LANDPqjXtfbKbcyExRI70+AjZ+gLpukeFgcmDx
bivOY36Tc0cFt6g8XY/XobXSXE8J9eSWru3m4LdC8b3Nh+mCFX8y64nXi3tu
qg4v+4p+J6SYjFr9CwJWh7oKK+heCWaxA9slX7BURIBmbOWmWkJ6QXQcY6U8
NMBMtd+wXD7/T2M96Gd6kshfxzRgqpCLEPF1Y6LDeLwt5OGAaR7zHfeV9xq8
8ODVJMGh4mO0GZADQ0Y/LAnd71Audm5j2DuvHURpK2SJVdgeuxn0Z1ZbSbkG
uf7IoKmnnWu88+jDv0Ye+cTrwhG1EG/UHH9w63Zh5qGM4ToxupyHUVJpBnZM
WxerpqLkIkGFIU3LqZ3eoQYtUIP50zqoz7AmmO0KwkM2pWz5cDG9iQm9UyZw
Rt031xvfc9pR7ISSwBeuCN8ZTVd3jq/2P/KhTGFaWsqrEqU2mCwxaaqVV2ux
sSwTN723/WtPxl9aLOh0q+vmJH7fG5MyxYCikSjPEADvBXBfCjS8sggfv7U+
rZdpCVl+SzBnlMadPoZ4/HKSHbttN8mxnCRq2DJlgScEOmeKo8kwyvt0vFHO
QCYqzk4aqFzzYxDCDbTy2uiTapEx0kaMhRUnvp2jBikWXNBw1KnWe6PTszxt
a1vQetvnZw/1CtExgx/Pe3XTuGmRafc2u4cnyLRaVSD7Eppq45s48dLcAyYm
Rqrl+OPMFpX1d6Ct+zKd63kgBJAxgBo6NxgHCcFD+tk+a5cdaUKHf3ousfXe
v4alBzq+cqkKhKyRLHyIRgQyPk/37RnkUQ0XazXFIqMt+mu/dGB3yK6ClCpU
Kdme9xxNxXiAgXbY4S1ZmiQZail2lSQvak6fRwsaNc8rFGS5MrOUJBipzgDx
m2pigZyj1QgFQ3/e1vQ+4ddx1heG490nLI2Apd0HS7kPVBwDAtMAbBJOZBgn
BU4IQi8rvcJL7RbFh3xz0vkNCUH/mRfm9P0sMsuID0bd+4SXRQpSHHpPjCsN
jXqn58CJcYaPQLJupWUfRmYgiRn1puNJ9ja0EkO0xf6gwevC1E0S9kWYlsnu
adsfrjA4SfohpaW9p7/jCR//NOgwiuRsOUfl0rbxTo906xA/9xuMQJZzotun
IcbhBilYZaHugos40yrvVkiSeaXGO6jN79hgeN3k1Pd6qhkNSesT9wYqcDyJ
rEjWgzwyYIsPVEpbmsPYMkX7uITljuHnHHF5tBdmRFAlBQoooNsnoiqzzq86
FjadbeshWFXu9gpRAEz/kXir37yDuWdryVZWQ6kXl2IqxUeVkws1V6uGyDfU
pPhlg5/ksUgR2xkozWSbTaBPFVcTp5zggWvDCADHkByx7eYl/O48zpyQUBPz
N4O20NHLCnBJdIDgOkquQXeXUxGm0jahKICoP4YMlmeZbEsL2B7J8LmOmCLi
liA4othedDqhu3reok5W4elNjIiuczemzoTxEvMHTbgp2jowTkHqWd9Yv5u/
vK7KT+3b9r+k3yzTda+6n1gstk4agYmAjDa/t/S/H9EqY4BqXby8oGYHSdrf
eAYV5msbt/al1A7EH4Sc0ZN8yiPEvbIPyzZnqELw11Styigyx92cI0icH+cn
VEgYjIuKIFoTtHVMAh/nPzfMY11iXPXezYY/yHw1wjzXIHzrE6XVdQ00WDnT
j2cKYU7Pw01a11dAuLf8PYXqH17ATBwoy9utTZrL4jszWEC43mdVngmBO5K5
1Bb971H4Q57mnkmg3VMaLM+jbXZrvAQlArPCMHmvsamTSVBoR3QG0aHwkqtq
g/MClaUfmtiWCBizXDPm9bCJqXHgMJIFD0j8x6mKQiv7qqbb6DX4kpqRlbtd
ss0Dn2zdLfbtYAwALE08MFnuNU1JRQmQPoXnHyT1Ewi+BqN1No5LNU9DHmPe
ZB0m7teGyQh0Exti6CqzRDIGXLbQyY9Y51MAU9QpFBkPJhHBk7Ydb954GrdK
vqXCaDakgnwRfZRIALJgbsG6CzEkqto44H6C2dSlFv9N2814jgA/C4vjtq0O
6LgMsUsqCgPt87nUsWq+nE9J4UFS9VESJWLvaZpp8Laku39jZXWyDiYfU6xz
WjVsBn7NRecGFFg/CCySZKfHyDvUzP8APA4tHa6Dj1RS7jre+80vphHJPp3L
SxajJbVH0JikezmoksCl9D1tVqjryPRmTK7uoX8KlGSpV3JoiyLErQzsizSU
v0dFEPSzM8jUROQddj5kXSz6Y8NlT1nDqZ9uEZoEKf34a7rN14H9nDhpoUNO
mvOxwUNDOzmt4UVjO6iI3MqRBimcbfsECfYxXnYuL9J2hxNOhsmfzNAGYL1H
ncP4H36G2FARBoXoHaml5n75VXQc38G1mUWQ5DJVz7UNwT5uxywFsDkBLn82
3/TSaQLKaw5tJaVW8c30+7qeY5Z3x32/KfRVnK5BdeABmphFKJW3BLiFtdOp
T7IozJSliri0/fWMB87tWgmQR4jezFvxN4NAAm4dOYoocOjU0ner29xh+Ync
3KMSToZvXViahVbJPAvYTnsEx0ayw5muuOKxPr6hibIXXWHnCZWbloAxz8vf
9F2TFHJ/ENzooqmPK329r2jKYpxwWW/A9IyN1I+58QAzOVgpI2AcG/vpsf8Q
o0F8G0dJUx+IiAMwNQXRrx2CqpU5L8JOlPf60WPvkjNVyxHU1ASnvoYIoryn
i54XDzQ/dA9i20trXufZSecU2Ds4BYPiQ8VHYIQHGYYWJzc+GTXcrp/seOn0
kq0NbvRFUL+gaMo/izguNxLNY7SM46154/chy/mCuEzmM/J736pXUZQjjOI6
tYjf8brL37yaIRxj4sZUncUuWv5+WuP1A6OgNi6tcsuuzuIKb3bq/ArMM7oL
7qgD7gACOKk0JQyQPYjHYibXok+dMySRWUxYX1EZi9y8f97k/uqeWaZqmu0I
M7zZ998NMl8nK3pi/cYhY22m1Oba3LDktdsuBqXgjqKM0rC9VZh2Cn7wgf3C
OipsvADeNR7VrW4J+MapDMxVfkdBrWqoE24oE3UANe1lRkz4f/wpbhnkEjKu
q48aYPqUOsuk54AzEFvfVOGR4lpUfotg4X8fHEq8dCGbJkNrYaFrDWdW/631
D8l7ylfqIQ8pMKv8duOfhhlMpP5p1gLAEu4KJQB3guSJCMUEg/azf2Z+V0JL
R3Kpvv0WrqyU//lp38ddsvPFShdHH6Isjfztm3zuiIQ3ZXazJswFqhJqAqmI
v46VJBbkaAEIgn8pt+Q7U2yySYLwH7oO6r92hi+CSqkSjRi3qUAoD4/LAcoH
2ns/8EpaG6WzBD/AVk4AmtgkEzq/OsD+D9ijwvh/uiRprZt5BGVyL9DOQwgN
uIfSX7z7Kl4QTVvSZWNQfg6zhAuiSlH99Y7yeqpJeRY3fh2gQ13E3tuhhIyU
y2Hv4TG0QzvDJPXr+95+33cEh1587ilfFhSpBefnltn1l3/8DF03mUYA7vNh
LASFCcAOkTDIXNRwej15v1kTldVMU4FkJ7HJ2WMdihx+iuRaA/vDArXmBsh1
6VJgsufW4F15q0xA1cSEPw9ClgcSWAXBrSi/B3RIylp3cJyd8lC3/4LOeI5j
kKt+VFJ44GonedrjiL7vly1I1+7upcpEz8wDkT+Fvd7mfDyihuUQIb5F/HAQ
ddCpi0nIMdau1ari92v6Qm9kqpikqhWXXeKbUVWNAE/4tRJPh/9hEzlKfLJq
FvAp4j1ckFN1qe6zsmlBQJx8tXWTjccwk2Fp8GjULciZkRCZl8lJLSvj39QK
mLd0t8iyM/gejyXPCeFIEljO25tqm5ZVqedDCbY93JAtZoCw4qjR8tLnAJAH
nPlbSR6WZOnkW9OLKYN6su5zyDd7jyfG9+0TZroz8LuA32IZ6uT4AopXlVdP
32PRoOs7m+KI9mHObig+pMvjJ0Xm8nnrb/akm/imBTF2W3OEjHQGRcreP955
uwajXRdfq3QJ2dkEsmfZIEBC/7KgVZBV3VfUBL1XiFjNR53pZmE/Kc4v2yPj
hN2zbpYxjvQlOXZo9ZQLiNYtimbRs0j+AwbUkkOcpnYCB4q+kwf4pNZbm5dt
UReJDNxaUucdlvuXK9NP5oZB26N73yFGO2qFfNZp76GgISAD4XRKpG4jraWE
Xn1pJ4Dj3rOPzZJmDAwrMtO+nonKczkWwIc235dYeYuvWR34sXX9crWQZm/J
kix4G559RlRlB//YtpOVrnJYnc5hXyaf6Qj6vhxJzSzHIYck2u63tLp233Id
7A0Ih5fv4qxU+VTaImi+7JAycIGaK5twCo2Qvn22kD0EL2Mu0xZwS3K9KcBp
sUB1TeswLxZo4zFvxA0unH66rUwhesjno4pRUpAYGNr2fblc22rMqf0v4Wj/
A6Geq3JDwQ5JD4PVSRKgzlfiv7K9+I14oxnuhAeQFanrJstYVgGoAX1zgcQX
EB4VOmIoDCzoExpRXeI0GtsDEK+lufta9kG2RSiaaMXDnj5EKyh5gTj+3Ejb
4/eEyFmOa2uuOz6qaWWjxm3CEJmY5e24HFLOch9eBLMxbQyBhMA6EJ/BgAjS
JzhuwsYyZdg2xAuJ98MIgNQZzxObAM1YPJUfQgxdv72kYeklYkO0BTVbQd9W
L/Qx28uPk59JVa2HymEs6Vw0atkxHKhztdnv9YNh5oGQQ9X2lV8ogDU7wkdq
pHdBdGuBjUtXer/bzJOzRb421Ce0+4idQKxcVaNtcf8EX2pijTB+J7pu+bhs
OyB/ybkK6sNZ+ONw8Uq92k6syY/7WgEBevyb+5HP2MGRdU9UeUovNjMgsgBH
sKO9qFYnVSv8wphuu+zR1+fpIaVOCVQMoR97HThRiuJz4v7nOA+tDAB9uW9i
7ci5bULtG5McEB0ceaVBgRowceZbov9KC9AixUYAN5R/SNLD7pGK2RGNS08u
QgaF21RyV7j70g8tD1+aiUqoW+Sb0zalSZiX4f+2cVE78b9HvVdNjZsF9mgp
iea86vJjxDeuDQM6gZZ7gSI+sNkhs0q3/qK0He1ayYdj9JUpwYF21ggBogbA
kNfktnm6svmhvbhFk813Sde/W5KSfxXJf9xTf6kGwaPIwQoNgnfUaveQ2Aaz
Am0ZVX6hHrBWXxsgc7FqxhVQO4tpXiJrxEGWy9hWX7QrJ6oGQcCQB8bivrAe
uiefZYfCf7tD0cl6EvCc5b3rjNdie6XRuLJu4EdGiPKRKdiT56eiRFSsFNDl
GcArsDiYO82OQ5GkLxza5NcPXTLRGs0TZNw9hUe1YeO358yZjtckNkX6eXUu
FHVbFzLZOEGCFYOVgzSPrxz/NMR802iOynrZ/p0g2Ht9Hxzdo+j6kHWPHpRo
KjYZoSZArDC+vkB4hf6qtEPZRsOqZk6S0RVKQrg3OaR8VpIzg2AHsaj8f0YC
wIkn8E9d+pYYS555cnrjHCHlegloyIvQEzB9FMSG+R41Y+EwYarLbr2D5k10
jFsyQgavE2g7qetVuvXOpfD0H1XINX8aeHkNdH8M4RRkHfXEBFIIZRqeRhgS
Q81dYh+QS6NSwuApst+Fi3mcOPAnhkeyqzxOlKrwVSRtlamp4iEDQkXzlW+9
ihU3wBgpNRJ87Yg6dWWsnFtVcl6H8SAHTRM8k0p2zJ662LOjswsogr08j4YV
KTfXh6MMFP+Sw8PJGSc7c60jkfl4j36aP4KCzRd2v3kwqZ1B7e+G/xQ1azRL
TCmwXtAdKM56dh8rAk4A0EQnUPJNKsrB4Z7wSAjT03zyspystx/a5Tb7+gNG
AIqn5I3usRNuV3orV2hExVb/ymJBdgm/oWBQanL7iu3zJWF+x9MtZGOgLeG5
Y82kW3VVxgn2tdpSsu3AWg+4Th396Udpv5Uol/h2ULkfwFDTIB2PlLg0FIy+
4PTySWZsreds0GFSRbkY+PVWlZuhy7WYlkL0kBb7bDr163vZHPtnJzL7MISw
6jvZp7O4qZ2qWYcrQLRWEfXl6zN0Du96oOZ/46y7Dblm04LIZfXTvVbbZhuu
imEhHjxItpso52rrnc9Yj6nY42N+1jfvZjIdr10xalOCWDZp8xLrji7FKCf0
ZI84R693t7A4HNrPcWkwOBQgjSBk4T3jXyVlZceHwmy1vgtDCELNeWfwb3By
KDX28DXJZO22vCCazSZWDPDUM3LbYQf8Lnab0XPJrgi8I/HBsfT9pgLv/MKE
tcVaXm2+HrMtc/7ukx62vjO/k3XGDY4H0qbVYsAECCYt36iifLHSYLmaeS5O
SDXREvXitoRimx6KhtOc8iGvt0/nwLmkDJwquhgDYZOgFlDRg+ciiXt9oL/Z
ICuVPBPqO1f/+HtAuIE8KHsKM3YwCsAsHgy4BBqv0kJ3fy10PAgyFxbUqRrK
exO3nVUEgt3/Cj8YTcFyD0wDXtB17XoU79BPHI4h7Oq9e3RNi2n2BlLN+YP4
EvGN3S0mi4EWRxPE3JURXg9DuMCJPhJ8PYJy9S4UqNGkYyB1zZq7xrqGxAwc
bVDhgbD77qqpq/Os9VLCiFQdQ0hvw3zm40MI1NKsyc9a1/LQ06RXwfEFzjwO
EjnjYAZDYzjZUO24L4pj0hLjig/V85TC35/8+5lNj69uZQVyPPiFNNt2+KUr
AkpGmSsStSUNiOrgGQ/BvAZW500Gfasq+8whGpSajoNi6y8V/Pi7Za0kgBTy
JYOt6Mya6W4u+oSQt00UM5SCDKO18Jh2wwxanNspFrVzwos4OAEK4NGkVLh1
iTviHmHclNH/7SHdNvTJmUJ96/CKb/KQnAwyFmThiOlTfahqqfAml2UUR+XL
MZjeJFtIHi5rPlP6p0OMF+lgOwGWTZJ+7hT3rsMZ5T2/rG69HNC7Ct1O7jzr
KktmCbUDPTedc8jtsF55HuO3Nc/16oYDSsgjIhjs+wIncSbPQlFc13FIa01M
ReQQwfbC3M7iONSEXjLoECHBB41CBfM3xIWBCdaP5e5AYj2vMUoX6h9/3Yya
5YQRmjvby/F/HBA20al3PO3dEHjSzjHdR35LL6IJMI42WhQQB3wglnrnj7cc
D2WPg7u1oEH41xPqethiZyVW39dPkMMDIcTm04ZX7aa/pRVgE95UlQj4sYjU
BGEOH3DbuLjrAvaMAKdlerEhkIyt+cn59shbcmSW2ne4e59Jf5sjeM/kSYdE
I/2N+byiBSv0DJYQ48f3gBsWHCaY1rudOK4otOD+aHpqpmpZ8TyHOa++KDgV
2nLifMigjjn/kHEdcye4GRIt/a+dMaEoiBUi+Rcd/i3XsOQy4wjF3gfwIOfI
lZz788Yz2Hhd6MAfC9mpSnxToRQqjRleR7c2r+jkflGYX1eiH2BujvoM+8O8
zH6rNKbNuRnDezPjnM+nQsOR/aL7rxtdAkyDI+Q2QVaKwANWI03wmwhpUkxl
Ta/Dmxem3rDXhhICnkADlrdDd5fdotHxrkGtI5UCv1EFBeJSftWz2MU9h4YE
p+Ca1OHfOYCxEbb+iGfTzTHobNMZK+wiDWzj0JXXs7j0sTDbrPDW8axvSOTh
A5QHA3B6JxSS5Qwl+jEVnIv8C8Rs6Tn4XTRHXYsURZkFO/bf1kTOQi5cUW7p
Jl9aEMfYtOPJYDeOEW53aXs+68H8EEUdSebcnCmc0XK8xG+KNbSHDi/d2QiB
px3q0fdnaemfpW129pI6sTAx1zcWhJCU4EfX/eTFj/o4xz5L3LmUr9/hNeiZ
zlLo0kb+S0qZ8rFYqROkohnsGk6GmUdHNAxzl9s6nDbHC8UFfn7g8Eryw0yP
ktVpCXOxW92X1vb2VN7dotZV0JbcvuexLKT3VhRTysCBKDtiOkbnxQPe4PfR
YCFOw3RLWMoquRt7abYFO9cM120EvlX+RFtceK2Xm2xfsGKM50uxnpEMrSPJ
MjXwDj7puKXiT33rqAmEob9VosqZf6Hgj3HTEheEjENypRJbXu7NMIUp1mcz
vKkDavr1ofaAMtcXyU8C7yQYXNCRfm33ODtDFsG3Oc48TOQmcFIeCyVW0bcC
mOCUIJCumpIKQyqHrpLtLPWHJbSgTxfY2OjrmowVVFM8NXhk0Ov3p7StXi33
Xzs+D/QyUQdWTJF5jNDY0xH5MDs8g15g3nsyNe6GWSD5fqT3QJLr/KsNRp9J
Ma+koP7IC0gnr8ewsDb6FgxzSKt3jXS1wQmJVOGC+Q1vxKdVMaZfxcI01OWK
ExNeEqOCo2zTAjVTxIJDREroLaLI12Uy6IBvcYz4YvgNxtCDIVSYxrupykmw
Y9cC+I9lGFhXHjmReRmVdzr46P1QmLd26ipNjepWWN0QK8KgW5TLMP6GD5pO
XiWVIxPA7ckzukv7aZIfrcnLCvs8Up2I0cLvI895l03Zmb1uM+tnM3oO4t7r
tBTZg1v7SWmMkx2Pz4Uw94l4wYVSXo+0R5kkLLdr9aGwvjGNphYFkk0rLVqX
Q9EYJdo5FRm1shiUu9CwCkdY+VAzybEd2EdbLgEDJ0+8f97mMJDQ03HsugQH
lJ2+Pa2rf9JfDWWrt4DVPRgUatRkYnvM+IBPG3yIRcyEtNrMS7RY3SJKBPQG
swbhTl7UL8t3eX+Y4oCszcS2QRZ9HYpP14W8MLKFKlNB/7w4LuBszoMfPl7/
LJ7ia0ryAFpLVOEPcvTMLBEDzDgk3h8GI7SswpQITF02Y5wLTNqCqEmXYLnp
8OOLcJmg66S5gP/4CB1JtpuEvRCyrPHe0cbMEoZm15uO5pD044FWTnP++Zhv
d2FM1oc3P9YH0dOK6WRtaudBCDEksNJt5QF28OrfbYn9KPn6uCQ4tDuLZWOk
T42D7FapQFNarlEKDFNWrU4KYq+uDgbw+8Z41jONO6XETt5jFunNVCN8w7DM
MKe/bxH87+sH7+RELKnnby3DayptV4YHgHDCtysdvq7zVgSzY9wfQ54HnqxI
VNE1xB4Dac4oNqNG2gjnwRuK6+0hrmjfdYESkrtGxp/xsKrgEzilgbe2RZDx
oA7/IURyReWSbeUb0tGDu4ubVFh5MZx27rVs+pIVBC1kRDsU7xjsCyTkq6yB
MfGA/yOs7ZvWIcD0CxYFc33mHca7hqfiVcxgko6GOZSHyvnko2upVL1lJkkv
fWteL9O97GoB4xBm6AoSzsMdJCFjb4fBGyu4oIDLCwoCMyryjIR35bi8jTpk
hvtU8kguB5LOyYQi6/gBugJhtT4MKY5dLRKqxHKH5tdGjpMXUEd498IcFHX9
f7ycvEfXf8BzV9mcpFkYx67E77K4MoHi3mi9OaxLUSEixzC8fk27O10DujIS
j5kwu/ZNA+7MvovEzkSNVLjY4QmCkjotsbVMoU7l3G2HSki9iLi40SQvhBWX
5lQZC5Br5cFLJMMhV8h+FwomWhUHyCbT8C8tCZ/H7AcqTtX1O409rAwg8HfD
T3I+wONOPSG/3o90aBuLukEuiEUPJoT5UzMQBNMcipsqGSHPSjMQKbpvRGgE
KoqkDMrYLs3TXpVDEki/q3oMvws1L0YpO8hfglVuqaFUoSgjjoCryNT9722+
mlmbkNHoLDoAcdbRxl/qFKODEqrMQyOwWLG12Rni7uVSGer7t2nLNk7pLGPy
JhUBEiz4DSkummsmToSsMeZryYI9J+XAyM8S+Orj1U2aQgdycjTRqfPVtIPr
mBpXVXc1xBEuev0y1JSp9OWYobl6uPXUkOMhspEq7+jcGW1L6W6dqEY10y1B
v9Ne00tjmimHhVhdK8zMIKVtcyYvdMkaECYcGzOeOxqxXytpyhoqCCIA9hAZ
Z9BiLaZ/HQ1vchPs7cAd/RiklaoSTOjQuXhFULQj8jf4wpBSe+IFFS2/69ak
ne3vn6Ikk4N1lNouTuSBNdHIkcekiGQkVMEjdHpgjnt+dlKaxE5xYKI1Vlh0
JtFr+DSkJzj45M+xYdbRXWVnLM72HPl2L43E6k7uEcgyK2XT+Y9FK/5M+Rqj
kw/2GYMiT/bxfItfnBqR//yZlPqfXI6kiBDm6qOOtSJL0Z10b6aOiqoYrSFK
9KPJEQYEYqXJW4Q5+wz6+Nuiq/K9FKZL0aq0UWhHaNaoAQ5bn91OrYqb2FFr
2DZKL5rM28X3X1C4ix9awsRk1pC9mBPGPLVZBAAItMZhrcMsEQ5oKCNBEEWp
Z86fcVY1iV4ZL13Vih2Z3qLUPcw/wXSUJrdFryG9BfrLnVcu3N/NHSqFYb7G
q4sXzQ9m3QnsoXz8fbDcwf8lA4Ui5S76cqFqTn0sryxUfpQsQWvQDPQNF5Ar
AbkZlAQ+la2edyVMI7cHCrbR8VWNGMwThlZt5ciTyWe17Wr1NHx+Tp0npMXe
L7CoRyhv6ohc7bVD68jwB47ryWWk3aXg3+rAS0PBc/HdhKxcT75ESVebB0L+
c93lVLN+LrpYeHlrWbno3UKvOZlNlStd3hFZsYS/sbM9mb7fhUDUJvBA6Auj
kqkSEu+/gRvLYDlVZL1EQF7nxaG1bFN66Q9tKrafVAQw3LmMWVFhfiKVdS2B
WmOXQ3paIg/0jmcnVApve4GdJWHYa0y9pxoeucotLmQ6wnrC/JLkJxRzXQ/K
7swdkpwxMFZoXS7i4Ah461J3rePmzCQLR751GN4IBHj+e3DqPInzDUr9bISa
mulsuQIIdThhZcM13iK7XX7cEA02NgQDtASaRrZ7T7sOOKcJ8eWw6jx2ZsqO
SPDxqbXdaq9ecKyt5JLhoj0k0RxOacOFSqsPiGr7oBVoOLstkzN3rKmuAdlE
K7z+hjks+A3MDavOBuPj8IM4IzkJIOxTQZI8LpoVO7q91iSTqN+qrzTJhaRa
gSXA6kXz01W0zj6H1aqqN031Im9vaHiRHf3OAK5rnHClfFMr09DWQp1hQ+E8
OV/p/O0OaA3WIe8mkMO2nqisBbKDRjA241jpMh7toJLoPC+DB7ne6jxNK/uI
Xuz23iHncUi6avTuFkVDIAyUnwu+rx0OYJhp8DUVtQNrvkoJc97zwIQ6Bbbm
VpCbknc53dDEBR5oLs0v4TtKmcdOLARiIJdIRAx1sRNp650PCLsLDorzzmnz
3MnsW8B7OcVEofJ4lQffVRkwNcBmitRo/AgK6Yr/7Ab6k9RgrdJpTj+ktlIs
6k3X23fYtxGYvv/rXQLGXmjfdl8LU1hWHw90grlHbshke8V0qImbtwymlBr4
0+GqbOqwPUunv+4HhrqUoPCpYUMTdh7cV7WFef49gfR7SvgyCd/8pdEy2JIA
iwZ/QYsD9vOzqTyR3QA92Lr2fVK0L+BC3t7gCN5xyr22FkU8S+h1NhrdJdHU
QLIcewhnxCVxndJbr9p4FXRGE/XExjVFta65lGMx0a2MH1gm37wXi+0X2fCR
hxcauiuLRZ03sevsyK2oBiTAEIP9tg4Gw61zVs/NKZ2sgfHrWUmeU8vfYNzb
Z427phHfVNXgkZZ5Vk6+0spK+Q5yC3vRTztKyB+zAqBP/UJeQQa4yr/lfrK+
BmmU1BW0/JZCTI21TfH81MYOrkh7NFNu4eeUzzk7FFUbeOieL+X7VvE9kYdn
j4pW3zllwzPaTIKr2UoHr2Uo1eaArh7lfvNijg7B4Mh4mOcIHNgVGts5mVIj
Tx/AmwMVbx4LAxDq1JQ5RHBUhEPpL2A6ewtcLTZrMCgZtBUT/95qR5z5WKgT
3jmZVCeE7w+DIJmiLY1resHHD0DgV8i8IzJy7GILCs6xZ7jaZSQxC8fVJmtQ
TnxYgwz0lRRNtoKGilCbxK44C1G0bcTfIK+d8NCWYVjBlblw3SLxrWTZPfSY
L4518lRT+HtEBiHAcARGvUWHz5RaUQ1xQgkCYRBHn//EPsfLVqz6+Q7OT2Nb
b00ieXXYiJ9v91FkUf92C1pzQ1DZZDWtAamr2Bp8Zkeimu7UHvXWtfs3HPUc
jav7nCNE9wC7NZayj1QqePF/VOdcifv/7n5okL0EqCDtphV3UolryvbssGX5
NuvHCFv4Q0i2RSceswPM8eKW6Xhzobtfddn7MzJqT+Ko96+7YWdo4eixKgx9
DE69d+flzHfHgSqYpLoLPQcM9pvxzpgRWqhiqitBYJK6VcL/syw3wjS/ewyu
VwpGpxCnTjxbUjb/2LahFGVFFvw+ETguR/6+/5BF6iHFSgB10/BNn3QfhEnG
wzxkh7htCOaaQsM6/GUUggLgQ3txwU1k0T4zUKsJWfGaC/+dC+ULLl61vPpW
5oKyIKWoANzkYJiHxfjuUYCrzHkEPM034ddOeLtye1chFD7vFrpheFox3tyz
sb7oT0+Q5do1My7xCM1MJe6GxLeoBrYrbf1DpZs6rjWigWAhJ22x8haepgPr
2s0eZJkaiP3Y8mG08f8ZBj8ILlupSG7D7lU9gS8pkDIEubc+t0SX5X9JqdmG
tvFylc0z/imydMlCi4knIg8j/+Mugft5LFoKMWCClgjf2cAbVtOay1A5e9lK
riS/9dYygWPHUnRrhMFrS2LbGF/36xe50p5KwtftLi5X/q4QdqUiulOTj89P
nf+4yi1SEn97yH+ZHO123nF391MRpM9ks3Sw60pk5T11/xtZRPahLIwaG42r
L2rHUF883hO4fuhRUnzKQsyzZJxOWaqJMq+E6cKDjBUwVNnhdi711Csvk32G
8GsktWcOh1krBRAGZrulFaKQfRaVMHJGPEgihOQTApQv980qr4w7ogi3VPXI
0nn4ZSKxy/CSqJprFE0KHU1pLuuSDTnd/VzYFobHA4QSjB/7l1RMVh2ZZLjs
1HrfP8DJxMccjRp8mx3xVWNS35EeIHLjVmlKbn7kYR9bCvy/2O/dnaIA5G+O
ACIt6Kh0O42rWTvjl8TJjkcqTxGbDgj4ps8uy7QuhYSsjiuLygOyyjlOuzZQ
+jzgSxy3o8CUEGYYcQbzFZngY6kuLRLGFQOECAB7cWhRUG059z6LhlshSjAb
7A8anefiGz1xlyCQCy0A1uz7MGoeh8CB6ZxXeAc9SpjW+ezgVigF4CN6toRX
noujo8nVCZhNQekkgMsqQDCvE9GYyC+hA0Rk2+Hdu7MGb5p+ao1s0I6w8FQl
c+OZhuKrx+rpo7VhtCst+KOgQH0TdkjN2J9zLaLiA31hxf1yOijqO9YB5V1z
RICoL1rY+YlLYXvvR+pvp9yydXY3Plr4ZjvqmKntS0G7KajBRh7tI7IXPDCJ
SArdpKjKcTMhbM2SXvmAAHQ/QgKyHIe/TyrGvortv0ovgrGf9OGC3VZ161ar
qVSgqlpkSGKVka3yHuSAzEHETpg44PadtEz5CChxhjgVtk8mrX26/yadPpU6
ujV2+O6jRV+rvIPrAeNNoopYClEZ0F+xlC1FKnz78i11mlqRQLhayVcTWea+
H5kzK5v1NIjT/rh8tgowsRTEvPWaUgl+JV+cU1AHtuu/GPoRt4xOBrwXvuJJ
6cpoqj1TklFCr/ukUGPG+gBtVyvp0Y58FhjEsBm4Jn7/Ckl3sBpiM+j6mWkn
OOcOB7jUezUkc8Gl/BBAeCswxdqInr+Pfz8Ob4xbRewzG/hXNfuenxZqLsz8
fye3VSv/3Vgb+5zzCcHkQ3O9WpwvZshJcPiVOotm58b8b7fBS6cRUZDHu8wJ
ARsA5Tpe3romfspya8dIs8iwqygmVMwk9S71sSKJJj0raIUeb7HZ4ZLZlQQP
6YZEPwIR3Vo40zQYkDnldBmFJ0yPdO6D5VSw41WHOV3CrfFqOMhDKS4i5C4U
ngQHCZ3iewwF82IMHPg9P4k04waQmn9YLTVvR/VgWZQAErQ1SKy7qfJY1syz
n3z9jnkZQ/AZP+wiJnPMlf47Gjg210lpLuph4xHmpCmXTsOg8Vv0tXFyg8+E
e5SAJB5yCEfx7bsvnHI8tfIn2z37qQkSgVPddaG/qF2rvbD5mmtA6isN96Ng
LhzVLfRaTZ6lC4G6RPKLoU7iUiI5MQLbv0/+mxx/x9zaQpQ+tNpetkx7WPcF
r2i/9XMHmKkEygU0n+10F4ZL1SwzodvrBBq9ANbNm0oHzYswbtuaiJV80V1T
Q3V6Kzc8+cjluANtRyzEpPLkYERFWZj6uaGCwoPn3XG9PHiox1+o62pIvfzy
oSk8NMikBo1uZn8qFXEzlsIdEZtQKCPNsFux8jfR8KOgJZw8hU0GkPwJcO9L
yZhmdhyou0pgH//e+tv/uBeCyx2N++rTKj59+uS4YQbpo8NA75hOnc1Jm8lU
Wr9aAxINnckoSMbYu+vuVHa4mjFdt0wcQP53ocnkEk2AfSXDvE8JCm75bo8V
annyezx/Bfd5/HxKQKYztAoe57UJgANVFEl2DKh2ZAP9UoTfMBoG1XkjXWpK
rzbarK8qecIYQRxP7w2j3cT+N6ykea9bqETTE26qTSkBIPPtN5q/IW0yksAW
F8oJWLHRQksVUsJ3B3Q0cuSDl2UJUqRdWG78QFZKxC2P+6O0WcaluI9xHU7O
E6VUGpY/H7DRRFLowCoR7yfJtwNQ16QBZGV6eHtVXazu2vKcoYzGsaKzaa53
qEiVtUYg2H0LQH4uXBooI1+MQ4SiViXoDKEU8gJY+KGDYY+ijGiQlmxcJkdR
fDOS0NUBtEUtneB1y9+DVNM1fDz/bzhYrHMfAObzAsO9ioSuTcF8Laq2+Jmf
yi3EHOy0x0ahkGToQGOWh5tUEiiXqNqvgdUjrEbWTI5urmUG9l0bIaqI+FY5
AqasdL8ESW8u/WNDbbSyAuKGY94gZXQ1WywoPYirx1mS0c8Bi92yT9DoHd7g
64b56hYqVHLfyj/gesGzjtTwTkuxlfGear+rGeOW5b0XWaK7AVxCy9Whq9oa
2KyeI54UcpFpXWco4KKiCWgm3P/8tpNqr30e0CAbjFxJdoDVW8tZipI+sJEw
RnXwwn5yRRjf1Jj0BeIrfgmzCIYGPo4WSG3+JdgUNb0Qjf8cA0qNTbWjSLh5
nyAYGB1EVWuwUGGWdIIM+ahee0yIuK9w3BgWNXX5WWIURgn+lgYP21BDahrW
DDLxDoyXhnZbQ94bLd9DcRdogL4Cd11vbH6ASHULeMA2sUGouf6WYCS2/3dt
uQLhKXclJB6ZcMocVoV4gi+EvnpG4njcBmqflk0cUukzgxdJNRqz6INwbju/
0Z+RiEFbj7UDHl5yo6mFmw4Y1Uh2JoMb8aLlil8Wo+ESN7Qn+N3ZqZwMT0zK
E0V4bIVqDaz5u6D9i5ehXJ0g30BnzZTCHOgPLTFF4GdKpc1akk1wOnImxwNr
JdWx+P8euPei8IK7fVB3ab90glVO4Y46wCg/NDcYaSEtXTbCZH7bnWrnsGon
WjDhvcDNRHK2U2l0eAZm2Wiut4gTBsJ7YxX1pNP9Wni2rHqxwnbnGjY1ZT5C
8cJ/pYIgjXJxc05hNl5zkU1XfkXvDDy9pPt1iG6uKkzHC/lnYhASDH7OtNK9
eSylv9c5CAFC2cAEwHUTTf9MT4kr1kz61gHzMD6V7CYV+26ezQpsTRWrpdMC
8myNFHSAnbWEUtPRcXA4GXVVjln6l1+cRilQf1JVw3+nkn7S0vP/3NTk60Ly
YwGzpOyqigywKJXNZzicOpVx1MWqRHkDTiYI6vLVShg607z/pLuRS/299vCa
QLYAH+G2WXjEqPwt4ivvfALQOiFuCeWGZNnXroV1x5gtWxlAUZYw973CCCN4
enWSdYqTQIFTZxPr5xJaCH4qz5qVES3gPk1mvRFy7jaEC3yJt0zxxnJHoNWc
RfJS6ugYMwjJndk+2mrrRw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTwINGCBenNYAbjJExuvgKdD750iqnVUEc6YEWoe82mHnTMhax5BB3q3cbC7fZqNOUdt05xIZ2Nvc0hc41QDLASARTU95XZuiWZQ63NNQQicZPThECZO+FTKFOVtwr1rtnNXTlMzQ/PkXBIJyjpLmKPBv3PNwt0U74dRpPYqsCdDF3uBd/flALSo8aUZ2SpvbPKOIhFR5ibar/npB0tOa797Zjr6DzXn+gq3I1naS/xDm+jrWd8nIw/hNxObanQNsAbkETcNwXUtVZu3CFmncDV7DeutHRcQk45JcYLYUjRlHbWF791z8E4VhRus1Ru2aly95HSnTqf9cR1IVAw9ZVVHAsrSjeFHKA7+uYOjJhFAdVU4cnbJ/41QcoiAIm4/sLcvzWei0MFRBi7vLw2+pUvEY+YFfig3Gz7g/lCL5FvaYAs41Ddlf555r7m5P510RflHVhoT6C8/phq7xYkz2yiWj4vwHZclwdbbGRMd0Ta2Y72aYkJRcx6I6bT2TX0MgGw2bYddq1V0KUIZ7K2sB1DhRX7xXXuW9LbnQ09Jbet/buE1gLG9d/Oa3tIZkV+AMGaMXmBgRZFVlSWtDsokc03AolAwYsOwcTww4f++lkKU7vGErn/SeQkft7OyV8echpyc8qHyiR+gkApA6tU+LuPG8vCY4cwNZ1PtSwgU62/XH4xv5tq+mhhb56FzdVh4kadcQax9frABOzNkUJq0opNAGURj9TgZ9XeiuHxaMa8lrIYrJ5qrqcZYfyU8qIRzxQBCxrRU0RqP7ykXJ5oGyqh"
`endif