// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GuqJLhb72+Ug2RFi1HT0UcqdGgGPjIzDdVIXPX9bimRT2HIgxQTWiFr9EMhs
E/ZJrb0XarrKJKohI94eNLH7+r6p9fWfl5NwxU0E7G+s2e66yXxaVcmj+r6P
0av+UzCLuZ0/DqBXjuXQDwNH51Bs+htlzYEVG00tJuCoYrDKqocOviP14k2e
9o+SVn3hcptHXCPVMyJRc2Fv2X538YIiJHjtNbi0+7E+i0+F9nQLjELsjwMb
shgOV9yN0ByvZwB3v6ZvLAJFUHpcjIak/lLRY2C5OnVTrTxT3BjruLP/Fa+j
W0v5fQ11U81AVVt9qbTsSe74XOD4mv0i5TBTKV+DBg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Qsp8JRl4Ch4FjPRsJloktlZgR8ZhzbJYxwoPArt+y9Dk34PxpGjWe96wd4tM
6uXNDhnh4xIuQXBC6E2QV36e+XSE1JSxomnxTuVgjaAkZ0UjZhDlfilvoYRc
1O2LUXDZW0yZrjeHfTOfGfkMk93AToQq3sm0ljOvyjPIjtkvNvS+HLPHaV2J
4nvKhSn3FDIsRE9K/zYtFfx6AEK6NrKMYh2a2rAmLfZlY1XjT0qSyFqNyYgG
BLWzJHLLTYlKzETaq65JtJpvecOacnByfRaYCgolVLuusK83u+Eg7rWT5ER2
o35k4oAZMizGLGcKHqjUybN//FG9tkPHBNOnMdVW8w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qVi++KUc5T1njTw9Wu3JsAim9Uc3y3Kh07wel718o+JAJY6kJ2BdnlW/8fwJ
c0VGpPqnCr9lTiJzlpDaKd4OUgAUoVvJR9kgTVUJKwD7TTq/fQlWYTT9lS94
QVke5D6s4uRBYKBB6kZMNwBYWW9KEjkSO2te3qIxmlnjWyypi/U9KOResEcs
ueCAfDRd3fJv81+KUOUFmw/VNipBd1/aJZmlJis/dgVOs4CmC8otO7x+oonk
WKyW7U+UvaHLCkgaYE1kx6bamHzah0qMjNr0VlbMMhMKk8ya9bQ0ct5u28/y
t3a1tzQApTilVnPc0IdTgWHLj7KL8fE+odra4Jlgig==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bHU4OAEnLMXeAULk7jYSN8o7HAqAbUsQ9n3MfLvZO69HkFySbXqIEbyU5LzA
jezJV+ZQynvVDnySkMUg3oR+yjOpSE0XYkdRttx7FKnSOxfXZRCI5aidLrNU
shZ1qsy7RR5+DgE76PdC1rCuhU2wOtAbOgBUFK60A5qbbxeXFeADqV5nFsb/
AkFQFc1XtRSbmnja1LE8gktNZENGVoERxX7+y8/8pTBOe0wNv5zwz91SIKBd
M4Xlw8/GEyHHi6Tut4BbwAf8V1Zq5Sap1ijCB4EQsWYNKGZaODCfti+8uMx1
oGeFOW4ipgQJg/kPoCM0qK7QH9m6Tj7SMvqXHgzcTg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d5NTmHd38+zMZBvUConFkoEREV1TaE/H57Pr+eWTWhhDwFMbRhc+UxL39HAq
4WIqFp8JPv3A9roHjqDCkJ5tcB/JOaq4T5Ivun09n5R1zRz8h/7cr5Ibckf7
slHSpSINBNv9R1pvntTl/ROkm7p06hwUmHuQbhNf54XWyRNqv20=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WPyApbsuU8yJCnl5P6B5iaB+TatumtfFfPHm2ycWp2Uh7yF27ZrJhC63cYqf
aViD6Uh5buafBNxBN6QiBBDgv4BTGJFqOrNJ9T3mDlCguOK4nrZqgQORDTlT
AdaIICJKmOD8sshWpDynBuqmane8MBQeX/sdlRhonvyqM8iT43e9Feb4evRU
8kQ7MrYv5LEdYE/oXi+h0uHQrbx0sVpEKEDXmuigd17AoqhjlxCky8wt2ud4
WdUFMxMI8TPq8b1IHki3e9ywU4pV6RsepfP5UTaerc+5T1s/2YWCK5zLy7Xa
18JcjekkQ5MkpzV1tSFkLMreAHnmmBXzpBQ8Z4xWQ8jFphjbNQeamxG2+Mje
8pRd5wl3fRFyCpejFMlmenI9Nh1dRieGSYXq/rcYwZp5iFbrsJf0LbRWxHBh
zbKmxcUW51O+tY8txGmRrMdXGNJWdETN6dNyd24nPDYEf7nJsYa6SmXoiMR+
LDL0aPxcg2+QRD68/5/awyTFzAPn9zhl


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s53okTwYjiyhz+s5oBzWaSfl8jrIiUlkIokPxG1HPLKvZTu73PBHHeREp7xH
hsh+UQqRRtNVpO139gGHEwhOFyuCSDReNrn4NDjkpe7AHIgZ2ASGA+rzWEif
4IlJ1kuf7DNJdfMOHOlMvalvQBMQI9qZrMHnAM5pgGLFvRKJxzU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NFiKhdsuXnr8mZgk+RsVFh316Mc0JB/SJ8t1coyPVEv99w9zFDDVEWcLzo4Y
02GunT9tHXm8ec+HJ0IfODcHONxLU8j+cNbK2k/q/lpnOGGd+XbNtJ9SyOCQ
qIezVLQliF59ItQsOlWpiDDBsG87RPjZTMQPG+CRuTagj/4FcFo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8768)
`pragma protect data_block
5bRhogg4x4SXkcp2IqYsyv7QQ3tlQayQ/vxFApjEp3pxVBvULcUiqOs30R+N
urYtIH0Ky+nfnVwuUqu5K1OnOBD8X3yYaGzJ4G6zCXli78c66hQq75uy43G4
gDabXDmnh1y3SZYxXhDXjzCP+/Lv1EqTvjXYlyMZM7MPXGqRFYfpP1nIHBHM
PRbPLtOD12D+Fu3zfnDT+JJ8Y9I5Fs7BuwMHJH0BQpC0Gs/VNViouzOE1vQh
QljiCLpc2A/tp3FsIS+d0Ljllr16ArzzHUesWdYhzkRu3C0JYvqRZXlufE86
GAphM5T62AtGE7VwKHO9jUmMtddy0m4LE0FB8rCLjyEqXsEmxEXKxgeDuh3E
LyCwv+ZgSNmhMSyJLP+Bjc3mJ2VjBbYpNSP8aocm9LMo4o56VqYtKS43d7Zc
y5NIp2Wy0vjEDfPothr2RSdXg38SLoxyLdMFKKH4T+DKlpvPhJl9gnt+mZhR
pVrlVL5fMf573Ah3EnoC94SR2jb0+1+kOLux9sGxVfwYeFktUMGBjfhK6AQL
FWmaquPOfQx4DJN4PYsl4gZlLRDOCrIc/vSndhyr+QHmPg/1swVR9AMOi/0F
XHWsYuZEtifeL2aonRRrhd6VaafBBMpscUDbk4UXV0TiUlUhdZUoJq5U9q1D
vFnaznOj5nHKSFmylrm28fu3KWgko7jPNf0VxM8RIU2loU/babAJIvl6p3oe
zikSG6Z1dfgKmXighO1a7j3khEGo8lGz0Wr/4zQ6Yg83uXlMAgp9WDLNpWcy
ZKmceWP9/CvLer5iIkIlKh/jqmVJsS+vgzpNVe0u//+qEmURWOQfxeu54sU5
vNq1LIsoZo/coTZEKiuaYWURQd6geSye1KY9enKu2S2CCoKbsF4xUN87yetB
Mvs7n6bPXu3v9nXMAyc7PSwuLrjFzLKTYwmJmV9hYayQwpQV/7EOb0FGxKx1
PjFn5SVnD2TiADOv3rpD6eeuLZhCX5658Hm2j0SjG660CNI8rnO9nHlbsU43
wzt3bJyjrQX06A2/ctOLAYnGzJirxbqvDtVhw3J7taophxiHlKz2PIBKp5Sv
xBJe56A8qubOhUpoRbbdgsCSOlUGtKBX8vO115pFUbrjmC5J9U5Bblp0W+rI
oAlWFV4t6qMJKVLmYvxKkGQ5M+0ba18qv/f9mvBP2vuam4CqJX5ZzTTtEgUo
3rplsU7gHbtR1/7JJcv4iY7iCMu8Mg2Qx50ub08nuswj7F9dl/vCZT9MMhvN
X7OQJtfKNKpcgkyOQUKgFnk7nPAcrTXwPgbfOx1h7WZMlD0DI2fL5P507zMj
nXNgmi/CsrNy/c9L7fotgNRfyfLyufdZpaMMJB+Mfbw6VhsU2gjaO+7l1opi
sQWrP3I0Cp1cJvJkzNitlMsULRkPFInGuxYoWY4MzFlHKC7JHDHr4XyQeSNh
JtzkUwLgbH6kE6bLTOAfpJotFgfoBvasLToaXjNkTVU1s4/N/WKh8WLevzGS
qhzcu2WvBGQmyfaoD3+MHs0soR34dngn+uz2jG7sbS0irv/G0nvuLMiEV++B
VcgtNpeK9R0YHRsXaBXLyoH1+5IwengcgaYO7uromjTsAgp+jwE4Q4a0K63h
lDN3/s9j/jEDkc5QFMVwrlKK3Ah7lG8VJNaWDJfnvc864Rrylpsvl5q/fMUk
HZHVKgAzwMomPQ9eIzRzWh12khNJqRa/V2/t3GY08hpou1ZhdYCy6XOZ4y7m
dPdISs69ueeY+GAWlP9Vl+FuL3v8mZ9B/ruYr46Wm4WvZrQpcPdHIoUqh+72
xei9plgIJ5YRQMrIjXVQfnmU4w9Gs0GUUqvsp8aHe+VMbtMwANgUVsxJXtx9
PnAKvBSPVQmYkzPcB6xpX4ZCmUzbX4TxSiYhkw8zpum6g/Vr1vBzV3Xm9dot
PlMiKdkmIIh2SjwA++tvq73BhMalx3ddQ8vZK2lS+2Zjl9fLQdLJ5AteB7UJ
aatpUboQZCpmxSY6fd3KEktvVbzSrbBMho2sa8wgA48F/fM98YVgzNiJdYp0
Rbj8JjHLrTQ4mh7EyCOQLFxnatWCZG6TgVfebtsUxIaAMIZHKIqPiXbJjXgi
lITJr9JihIo8oAkFtXfivfOhYIhH/cECU1gQtk47kEr++YHgiRi830JygWx3
4dauydASDbct7iWWzCJHkci4ojngFUUIipgjjaDo9Nq04wi4fTK30NtgiH7l
fDUZvCGbQtwQdka2RDS5T14RXGe75XAyPnBdJYB/ii76w3T4HEKeI86ZAtsO
ohMymiZO4/SUwLcAt2eUczTbo3JjUmhTEGAdPPZ3NBevP2scp9sl7uuQy6pi
bQxXxRnnFFLAxEf1XTvpLTVduUJ5kjJaIlLhocvbzjmpo6c3RrpLXkUO6mYN
1SW4+daGVnh1F9AbMPznelfeFVkNO6aVfxaUBUrfIDcAF0RTvAldQ4TjZ/qF
o/RC1pD1zlKmtkGBMQKDWUD3Dfmdl+G9W8KASsneZqeV4YD+PS0nMVXgdCBy
xu0o3bnqmuBjS45vC/9swXPipGBRCE926r3N6E/q5JN03c4fRpWTHXoiU+h9
vJMyHn9RQMj7hCafY3Q2B/67dW1XXqaWCG9BaEEsXpeQCRs9QFsh2VA+vLwo
Atw86k55g6HOhLIx5dagPD9rtg5KblImwS6vHOG+VIGUogjCIC5BWm23EClx
Wa4kEXcmQXXO7G+3ZRuvM/aGN0MnGDU3MlWOilg09k5UO0lcwf7dNWNKGRt3
XlmINb1uB9xoimGFlRSFjEwNwQIlYwf01zSv1n/yP9yc7phJCONpHYF2YYIw
fsIh/IWCuOMS6ePKfxBQYFSnfbAOzjHJRbhe/ELevzEOgknj7t6Ipw42SDld
Kvd/cdbRLaPaWsfub3zyG3S9s+5n6m7jmEB0fSzG5RFFq3hdpw/0Z2XRSgqK
J20/QlX/VXWyosjMuQJvNRfSS2QB6qXoFOBnb1C1PK4hCxYM5QXuuuBmiJkq
xiFdfeYkMyrYz13HffVcjSyGBDVzqg7YLIv1fCSeBJjmZDfGu3nC0nHfjwJL
4jP77lwLCDK0Q31IuR2V53u9iZilxXfJFFA0x9BgclpW12iOpygX7LqtNVfb
nbEBQezDA9da2pt6q0eaj76v26RfFHNwGgJnP5o180/0Gm5R8qsdL5GZpOyn
2zTtuPlwLpsM04EkoyffPLLTzDOV3UiH2oMshI6uWiy0AHkgFYff8aWzEVq+
XrLOtk4DAl9hmpHMcm2EbU3Tyv7hBT0WisGg0dhNu0nXqGyDPdX1kNFG69RJ
7PtngmfdA2AuB4MSdXmr2JxzU4Wq+uVLgm6+/Hw2H8OPh9lLi9suTiHUjSiV
tXbjWYOgCDlFQ99RJ+RLcIapr6F67PmwBlqGyv8lJsb8UWlmm5a1o9ev95Rz
bFp982X42D1N6wz55ejmClWBmdiQf07ywtWlZ7fhjrO+AsOVr06rGGxYG8yA
z8lBQwWZekHiky41386y1Go5Vf5v2vDmObNwL3iFgBgEMITE0kRpZ+Ympy5A
32z5pqpzovc27PJ+m41RXN2+cC1HhSQyawv7XC8P6Dnno+Q1hGOhMuZC4Agg
tuIttzJ3rCIZsk3Bg+Cw4AhMwbeeQt3xyV2/GMWaE8Lvps8WkfrGjjbHuJSS
mSqR0hnVm0SZax95IVsPxsbOlYp6fabcucH4TMtNXkJmYh1w7ZPBXVuUf2/Q
4Latb2vBSwOiELzZoByCxiVolu1I971FfTyvxsGowY+iCUzcZ0HNx1S8fUd3
71M5E0WPL/Vm8QDaDpesiEulSGWuivt7ONocZ0fIJ/rUofoFtwN3QXnEX/CK
c32t+7Uejj8Kwri06aKlQrx3OUY1XYX/hqMobjzEp1m5UQMqSR4kuGSbb92f
QWmLSinT9NcO7J6SyEiv+e4L5N1hbuaZZP9IQyvkmtzOUSbslCiD5FKpmRKm
ZpxoLKGsS9vVihDhxMnmztxkeEiWcT3GndBV2l6Env6dDRUKJa2yy4h6b+52
oBbjuf/nikLYpUjVJLKH7VnF839UDAfK06/BG1Ex8ZnvhuQLt4EbTJu3jPf2
IV8MVfpbwpH/mB4WvklyfFpb1aCuoLq63TTiuGNFT/VRXUaOM8a5ZKtUw235
MIGAfiYrRIxJmzkhdYqCwpNXEGky1+Ko7NnrZM6XU/cL/hXUB3YV7QxqZNGF
+B8omhPi5t3WPoNAcdsgnleBQgRDm06wvE1ZO0JsHWc/IYM4cYTjYg2J6ur3
uymrM2DwV3MLSvDmYcHQmNNzcQIKn+UXyl4kB/DieYgwfTHbhmWtOHseewvI
Vcf04gUyOJ0PBYV9ZU9esIbHHysHXQOcL7q7Z9G0XEA1lbuq/Yi3rGdxBEKK
Bh91P3cYxE15bXPMYFPTwzj2U0wTxCOTE6mcpABSS8aFWOD7WwM8so7aZsZd
JBEWNqdF9mC8oqSnGr3mLpm9wyrjl1o/DrjaeZbKsZ1JXHWCPmr0xbLEz9lY
Bxel6sIftr+siUmYReKvQ74SjxyHxDv/FB/SIqwzG0Orw+UY369M4onNCFHu
XXmrxDWpZGZ3Ep7Ikxi+U7ouw26adVRH6qnr2tqc51YfDVqf4BNS+z6aiatf
AgTT1+Xt1xggVsnBH6aNf7PJ98rOfhtjtrKcc/mzpX4K89ZxE97ZKhJJv3R9
ZaIbOJepxLo/S8ph2ICMJHY2FpxNgpvhUcxWGXV613WjB2+DbMVxNYN8isDI
wNrSiC4z5hN6RB5KiDbbgKl3c2oyMhuA/7K9ol0RR8gqJJw8vcEc/W8KUuG8
Ax+W767LchUjXlWrMQ8jPijxctL4BRaL2Jr6SGNaofA27X7I3uBoAA1gcief
1Oyfr658sCLAT/Im7fLCJGnQx3xMJC3+SC7Bi4Cx1XqLJfbptXcWJxNc5BeP
RZ8Fh6vV7jxoe/jBGYaG2//Ae5jnTbZz+DXr9yrfIqaVl3nssNQzJ1eCZ3dl
XgUk3W2apBdH688S9a36xj42RWhfhetn8AbDCtdmG4Mg31/cQfi7JUJmbLmt
42sOWAPyILrAiwSi3yDZ3pf73UVusJM5T7egREXlliezazbHZ8fNWeavHGO1
pglqO9DkE3U6K9FadlosvdR9CuktyeaRjkg6xChvr+hn5dvttAqLixtML4Yd
mlXuV0/vL0wlxd0ZJUQY7MTcUWDFGti4pOdjUqqE+/P+oK1wSOF3GCX4h8pJ
3bBoMQigfFXvjcYuVlMSyJRjlfSB2lMIgiawOYeLd4hf2Nm+fd2DnPb+av2q
uF3U3Tduwmztkh3SL5wcwNuJ9DYZstEszjgm2GT7IcPTgGw1ghEpwmOHWydT
yxldn52+TcZ3A1NkiCeI5yo5R2ihBmOz7rMSIvNZvEpNZXiKzHcE5uVRdCgY
VbjwJwwNbn0BG7VOySryT8aEOqIjzmMcSXAbNfY2Xg8C/bOBld8mew0VEA3R
1Br9C1gNoAUrdMpB7rT4fKD0ymhtRS+Dpmvc8tAykcRPjS6d2hWqzoTCWDFw
mVoDJMAx1UghFHl5euDK8BeFJlpL6DFYGYp4DneaBDcyUdMSAojzJJp51sN6
Gy7J49fhLsZ6E+3GyRsaqwVeTvNKV7uXQPCkw6VvUh36hNY6QdVqk0bLlwmJ
AadJP4pUmMMqoDiC4ImA4Q3qlo9R32exs3bf5woSmD9Ik77s4RQM7Sak5xfS
81c567ocVVX2iXoU3VDng8aNWXGoPvwlhPTSejHsfyLVmO9cmMTDg2bFWyAO
mrIBsGFng4Nrqz3F70W0DDg81ZcSop8mE1y2dTmE2l9NHrHA3dKF1st17ESq
EiWpWpHDC/amz8ru9VWM/WpXumWChn/Fqex6LuIHxMAiyaxg8PD9MyspWnxQ
qJxsPYx68rXM1bZ29uiesKmvnWGzDfW1UBUfYaak+gJA7PBuYlbqcfbk9W63
yta0wwyCn4j1famA8Sk3EWTzq8wj9DoKciFyHVKd4u7PPN8jOGhx9b6YxvVZ
CZJJ8MfsJH6EaAaATomcD2vRnrjUWpXLWpRkoOpKjYzGzSxIG4M7MJSk2Lph
ne1hLetkvZ4LZOv9QyxmlWJuI24OIJwVhSYCsG5SO6x4DG3L2KTDDCWLYtd3
3txNo1cqv6Q2H5eDhcZU/7lcBjjw8LPfytQjy4KKZ9oXmgWJ4b7mLsS1vCpd
I2dQCg0DFvL3FgoFHF5NL3uUfKcWIwUPFeIk45VZSiNP7QIksgtd3IaZZ3V5
V6tjjaCDEUmWHgSp5zj1UxT51MKkpCA/6fwKf57IOWQFm+zIpgg4F3vChFNT
JcCEWmhOjQnArW5ieFwKC8+1SKNUFhho8BtCvs2QfAHuwhzj1q0phwqm0vOA
MMqbBfrnukKgKmR7fjbJThX8Epp0hNTItVoDJgS+nIUOxbfgxKuHagE9vgFV
9tuveZkQ2lRb7zedLQxaPw+QP5++XeEx43t9fOVfmqhQYyEffHsjL45uYzjO
X4NlwpIlqS8tWOBodsJI3eNYlWJHrh+nVKfqRj25AQ48VR/p5pbNVaMWT4cr
Vfr8bGPaYgfqyxlD7tCf6atao0o/MMjM1Rm6NQ1k4WYZxy1J4bS8c+CkGrwB
r4VXulDmGBqN+haZqzhHX493/uXRqbg2vHEoC2GNyNm510EfxPRBQh9fqmfJ
8Aei69h2Dq+bfLRcFwzwNBtMYTcm8QIEM5tqG6SnvBhqgwKwIoKTWApn7J2n
VFJIYfn7qHzu0myFq62odQvm7s/I+JK+VMA901gZ2mjcnp+Pey8nL/AiQ3+q
Erd1ZcaABUCGuqMeoufszIpGgLOvZUYXBdJ2X3eoN9/smmT8ESG6HSShfROm
yVwPGrDkYz3LdJeLKtqH/FERKOKwDAXR88Zw9YKIDqC2RZxEISn9hdBC4hjC
eY3wXGiP4/h4n5CQfli++UW0ZPLLmssEZnZA0rkGsJTtCauZXkDnZTA+SCq0
nJKtkv5KkWTdcW+6IaprupxhxQiNPRVSI8qQAriQwio6+/sxTm2bKaSebMIR
ULuauC8IluoSjFl5xpSIks+4G6L3SZwy3KeHPfHcRxY12SkN2qf1PrBpxGpp
evLSzuF5rOmn2CfmXWavgTkfMZEF+n4+Gb7aIEQF04/ejd/oeKRXGos8EVGf
0ZyFdBHxHDdA5++rV+9rsmgvXs777Q6X2ig0VJLKll9qB5sl7JSAYRsOFHW9
cO3DrcghfnRv65fLHkBhJTifAFkv4UaZ4qxcGJ9z8X+wwThnMkRmpTSz0hzq
0GmcewRo2PdNvt27EMDVl/YR/XweZtK2raqkqC0P32S7421Uiw3q5c4B6iPe
fpsxxrvMNDNxGKaM3j7c1DkCFLjisZue3y4ZF6yabV+g9ddnEQJHPSLbha56
78aDFkWeyUW3DSVcCZ47XmyiYUjQrFQ6KrhTOaJsAYx/SehEqa2uiyDg8IW1
uCGYifcxeu5t4TP8Lnh/BPMJ54GwhCTSJxtuknCuJAdtmeOKzktAHwUzwbt0
/9A7A+5ksqzhr6Zb0xi9NaSbt3PcGXIlN9uKU32g3mkxev50TD3TDjY+bz2M
A7K0rF8l222qgabolcuCPhcwzwlceGu8gYuOwH0C5zYOyoDswJp6PzkDpKOQ
xMyNN+hayL3rNDNkpLcQQl5nI/kKh/ettBCVUFCxkWL/b90GnitjlUKnRGtV
6xsxaVt8leqhAvHSddOlHfRyr4bMnB29Otf8UkEZ9iAWeH7c2ctZnJUIiVhh
ZQowHgqBecbMU2OAVOYtN9BLhTSn2+uMcotNY2muJ6iebZIa1mcjsOlD4xzy
WMzsnhVfeNv8aadBK8P0XBRidmiZXS03es0ZGqd6+r4sNXBqI2sSz/2gKu+j
zkic8I3Co0SyMZB70ygcqSuykJ/Vlgax9ptd0s2qGO2IqKW3Whxj6TxDkS0d
Ck4LH5L+HiYxmmIW6+iytmBdqgJv+DDPmyVFtyJ/OnPM/ACTndiJYTuqt03J
gXN22skQUZYpooMj/FSS52/iyV2/58OkFVsagsGqnTm+lGD7G9MXpS0ptxCO
S6Vb7heCLsbG3WLhBD4xSrzTYBnYlgd47p4N/aYP62QRexTVSuJV/fCJczI/
XJEP4bntqlx6QnBiNoFamf41mpHn3JvQyVdeZhwSto79sO7cVnRYersMMZrA
wrrc8JY5GSo2bUdBw26OE3jQXk7mOxkCqRZ68iLnV/19SGj9S1XVGfals2s6
Y5ED2X9wM73Nyo3RYroiUm28POiSPEUoG7b+lnms5WaGV3FZFI+zqPXHoKJf
FBeHE444gqZxoJgLtaPio4ljEQL9N0c5X+KrcbM3RHaobmXzxTQ7j2CW1r+Z
weTPXfIMfHzHRpd+o4sl0czBstZ4DEnkJrezHy+PSeBfwHfooc9p8ZZGuIMl
Ag7p0IWX1Tp5c2wVVDqO9Tioewlw7JCFbIkjM165mb7lhNVToNN4tYSEyGNP
ne4VrrKQsVavMgwUI4HQRQqFaSwX3aEl5aPV8sqC8mJC1nR2QSIWTmUSZaVq
XaHV1Jd2VQZd4hEsQ31hJWQfkjM9CI1yV7Hj4BAmcmviMVjAp2DIAtIYZGN6
zzw+G4Ota5fcKbSM7D3jqWFcyHDtKZNyGKm4CSBOWf91pRRNUxh8o9ZKhW/Y
8CbYYxlwJ6NlYE7xBEkybDMT1VJQOEmoR+qm2AQee1BVJhYO4FCjxatYnSG/
NT4PbE09kinMGP1bYGYyTXxRBu+IdE91rPxi1FryUCDykRRRGfovrcp6kInB
uHck/ZkK/ot4tPXLsWCAEooGooiokgknD5b3bnkx9bkTTFhWu0waaaXUFbLt
TAyTw7GJglvUXuph0sCc63SRw6FvrxnE8pygNpKEIlyz5mnDFMEbOXA/9pCA
hJk2A6YQH7jGOHrQl9lU9tgEv1409xwEWVO4ZmbA6lw6ZHIypRAdkLEDYcXK
PaovbkuflhvoMJ1XkN5XC3MyMFu498GLTdqfVmDlzpe1ePAGOpzmutL1+6Re
AYr1uZxceOGsSIwiDwRC4G+3W5CAqXsycZtsIfio89kTJiWEhpOdlSpKShpF
GG90lDGz81tM0NUEPwk911R4N8aXMLI1tonG1xRtE+G3Ddqv7C0cvICiFmlw
BEwPadFZKA4YjFTsElH1/a5bdV4lAvn4FiAWHDTZJ554v3/AxyIE5yn0G4x3
UmiFlm5fNNZso10l0CD122OOU8Jt2gzx+wOwwWV4kWidUTHz0+/yse1sLFj2
pQSybt4QbSdAn/Px30HXD0bjBy9j3TPgeuR3kBU1NO4q4jHklJXHsNkmWTLZ
OgCcgJMTKjavDC5vYosGrC4ujS6hScoCIwmcKby1TWcQnt0BgKB0KdyhxeKi
aRnBz4Hw1AIpS3cogTQZKNFZdm3hQHGgXLcZ/mdmtY0+P9M7j7dzjk+CRPT6
8LkjTHYAM73/juxVz+6jihRSUre1Gcxb1gYEu5MzFxcaOjDFIAqrcMQq81mO
c5GAj1PsgiV+g8AkB3Xn0VI0eqtSVIxinDrf9y6DdtQw1CRsYi+rZObzK/eu
0tLa1pjTB42CQe1BSr0tdAGyjLDZH/mH9OVGoTs8Ffmx019/7u0oYbKG55/b
VaLnk0iz6tZ5opecN5VQYo6nEG30gZi7EeQcRGLHpCg/WZkbzTsgv7ygfLx4
C0/XN13dRhqz/2ZFcxg3VUGM8x+sQF2EQAEQO5BZcdGwLrUFmlxLslXPG2SO
v+vD7MuOj5hw+W2tuWxTWypis8K+NNH8NcwGo13KFgT4RMj00VDHAWUaQnjW
HlT9dGsdOKxg8TzG05uTF+hJRFiu0F0gbvNjSQhJDfKHvxO5KNRtuUnc2wt6
xg7VMxTYYylVXJ+vKUcybiWbnilR7strPnCmR6RTmFWzjDI+thd7rtR85ha7
LMSiftvUME55c7ya0W7HF7aRYCr0cZHXOW8e5+EMeh0/PIonFa+BuU3TpDRy
X97Nsaw+/bFi4hz7uDE296vHCtAyShns1ezOELbSHX/Q3cRt/WSuJf4GwBUY
pHmCwEIyfUXqOOD9TUN6UNFGBLGTyhzd9p3TWyYizqZzon/8uhZCjUNwPpF/
BEDD7pBHR5zTu5t3Ccr7FVYiaQgSugu74ZS9xutGuMcl/77IldIXTRLop9EH
Ai/qSaIlMqDTLnDdbfx07KEBIjT9FSFZq09CrUWpYAvnx+Z6FgvEuQzXDEZt
cEFH/rfw76QYSFnw4QNsEa+9CekDRjr2iQgUrKhtRtnYFBKz9YXKuhxrMPRn
qcZN9EeRsVJGnYM1UYUAWdyIQBUtJEvENCT4kDRb5utIuwF4JyBXJzD88pWt
mTia2anU4403hkhey3GyfdQxfij+2QMorXWlwcuI4BbCKY9N6bB1CfQ0XuPY
yRjtDUBPJorAzVHoVeFpOJ0S6MtpnEgP+nfZAksAWbLtvU7QxNV1NdJjSuh4
ayqK6c/f/42JmoWnKT7h/IV72K6YZz9f3n+6pPzXvNeznn2CpLwD+sRxPAG0
24mcp5xA3Qe1Cw4l/YcNiJjcwS73AO890PuDB9L6dUh3QogXQm5X69i8L0jS
56g0oZEwuq/Wcmd0Y4n608fTrDKNcuERqzLOTz3UPUM6CdS4THkRT4S8iTdH
AZAK2xdVvphYmwQw8GX9+IX1UZ4YEHWvZXg0JNGQyuIuX7AnEA+PRfDfdL/l
psQK4044V8SpJcJ9eK+tYmlkht1F4Uxqhwq93dfXlHh8GLuYIG7bC95q9MQO
pRr5Pa33366eE3JqVAM7su6kdK6OCjA0+ypEBG1bJR5A66ccn4PXB/ki+LO/
YkR99Fh58uW8Lac3x8qOTjKQKbGq22vU7wteJYfuJZ19RxLUebK1QFv9zuPb
lSQIfI6INdp3O0UXQSKvIZEL0KYwlyJa6nBSj+KeQXuLSpbA1PIbkJ34sx1n
Qtt6lTYP3Cm0T9dMFteRrfx2w1+MD9VEXw9gAOOarWc3EnEK25Pg5h0Y1taC
ZI1dDk/ejE9TFKHncuuaayGG2JlgskE/QI+P9PgWLyXGd7LtxtrJh6HzyRm7
KJ8NcWX/4xSPjwdspjLvzAnWwjylqbiG62ZdTP8iW6LZAuQLzco6eat6ZR9F
vzzn3fvK0fp7ke5W5tUKD3cv1uX8eh+JCxpAwyKi4SjQwtlVrw9DwAAaF283
MFG1vKhCkglHfoTawCjbHDjdytLVDg9SUVKYHr8Vt5uO4TuVxElG1bxdt8//
mzwyZtukXP5KDNDHnW9gnJA7ynRSlL8Gj4+9TkoQevDh3+f29N4sUkrkKOZ2
mpP/k1+zmPWB82tIs6NAZhxijiFsCBYfJV/p3ET4gnro4DT5DwNoYc/JLT+V
CeV7EHPLl5ofpi/n1MGpyy/JqR826mXkGNK76EsxfLszUYLxifFmOVilskzx
Rl+ljBlUQ9rAYHBWOoifZWPqix4am1Ns3Uq3FCMrziOiAGebznfDapuR0UmZ
4XMBiz5CKobgXFxGLyC3Ctu27gxfxErzR8xFvtDaw+iDs+AlNzxrO67sSWsM
kDOBx5w6SdredzoSN9WKjZma1GIoTnEMuydEOsZ9/gm37zSDWA+AiGn4fSID
fYn3nEcTjAtr/JxkbMuO8E9FBz+oUTrDDdizBr8uKEw6fOa1cbmiYFqD5TK6
DqoYOSS9DTGywmYVUNtl/cjfFFlcpmrUarALRslUwQx5xmQ4A5U=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzdnrtleyAEAO8Ma4Z9M0aiYs0+fet+XJ4fxPTluKXE0Yxgij6tyJ1icHP9tDTyMUVQ4onK+JHSMYX89tZsPSqPIQhCsD7yJAFVTTN9/tFF5ugEkx9RVK84oaUrzmwGzNjEwrQTVxGNdPFIB/lKTMVSPPRkPkLNu/AViHlDBfJL927SzouGV3ZA2buhOGhKgVmQc/e8mOEdKf5TwzfS7Ukqwh0pWJ5xYAaukJXZBY4V1xMoJWrlV7urysKW5dYLf+Co6bKkxST3QkIqBU/IQmgDjLAYZ8x2gJvQcH0GtE9Zsiq1EBZt9q2tlGBVQQ50uRC+sqWQ2CWBMq4MNbzBBOvv8gB4ZKMkHVKQS0xvyOPgoggeADMJ5lNnG+8JtYIkOFVFNTWZNHdO/xbZyqERl7WSZX9DwTT8HI7o8Z3xZXCC4t2ug7dsLWkFqacLSqAYOaOTLWiufVMrns6p4HQ3EzXOTNFnMJvDtxYb4/8yP1CioagQRJycK+OVic10oS98aATUBTnwBLkNEHzj7BeQjhvB5ZwOKBsIzAz2JpEqpJ222mGwd0qLegOVnA+rdLLFWNWivP26dlBGb+omxjgUrBVAuFNwYlKLC4bETfCx1mgAg/dhhgX9sAHc7g8ur2Ihs8M0XebaG0LHNYGUzuAFPO0QT+cR2VRLlT0XCdh1Ln0dhwEn5nN+x/cXnd7G6O6YnED+G50aXSBcRTRH0FJrQjzyLRRN9lz4bc7oJIT9yEs4YawWEg4kA7896XcWMx9ZSiqWIYCZF3PmnUYBSpf+XVw63"
`endif