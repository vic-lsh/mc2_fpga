// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TUN50TbHtf+ONYhRkLVmEd2bKUz1qa1WcndY31zRLcqh5N3t9ReU7b5FVXjr
SLe5Pb8Zcw4mEQrIWDv4GjzzbX/O5bzFSAl6xqLKmhGkH/ZLQqGRjqJ5PWFY
l6Ex1NaU6kL3I2kER7h3/x+X13ZohsGbJLW8QIAai0KS5z+WcaFjy0PPRr9x
GKIp4hh8LRuBbsiv61DV6d/SpJyQCNJYx1PTR4CfUpV6lvXTXDd3jiHahLU+
YIhg5RMub6s+Tt7qLlRykwxal7aBidooBWZUnpqg0l36tXji5c/nixYi1DSa
Yf95XDZitQlI8rE5mBnLnhg6pelS+z7PShD1aSqa8w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i6+fwf00xPdboF3RtrH09nfl3MsI6i8APAnxppvQ2kInHVN6PrXOTsARzzp7
rU75+Ox/yWStfWW99e1nKRgoFvN8+9hC+DwVj/JQ3RBjE3iRoKxro2CsdQMa
M34pQNhxEj4jiN5uOURnzZvfzP/jf5RtDP3Vv2FlDCfsSQK9FE5UqGg2WkOC
tgpAckr/GN5/hPUhqrGMTHQDJrULCeWVm1qw7JTUgNN7hyNVYl7ayJWpQnVf
jX1jQEKBKazp7HklTCahB0AMw1qpud3vwXDjtIGJW8OWx/AfT8AWw7DstA4L
jb/OylREpjfZqp/ROYCMapqo0vGWmVqII8YgHne7/w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hvyr+xMgoOhAeHO1Xy67q91opBJ2Gfq5tJv9poB7tjOaiGbnOMTXR+AzCmRz
qsRk0m0f1cFpOoq+Z8kPXYaHjG7afUPVKbuXtI7mDGF9VeI5q/Hn4YXCZwzL
wBTLGLn9vD0/exCf98Km3Vv+p/5mmkrTy98f91NEfkFR/ugTO6FcO5yugl+B
rnmHLyptlHnOdhWqb85pCDn/7/Yl/CWrY1mUAQta67qg9cR0cxS30viqb6fV
aCmzwBuoPMXTGL2oDIAgedYfvv75cNIn2+edvrQF8YhnHDMpi6Vo/G5Qw+hj
wPfbqmDPzSv04LAuq3T1ayo5b1ElSS/oE1m2foJtwQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d3mmaIm7ZCInzxNhhmtzBTxmGLn+Lwo4dJYF58clTxdnWwsJJxa8ZDLvZzeB
1/17rZa7ss1iCQo110oO0ItLyBd8QyVuL570hAVsY0CEZwOSC4nwJ6xusI9X
GU62heVYQMkkYDddggCjGxo1qf4amub306QjT8WYO/a84nRIxg6fJ43Olkyv
NreCtTH4ewRvDsWun6XuheFtCIvZGKK5b0gZ/v5+SD+O3IshgDUBs/n+EegI
A2P2fBOzgQuLw6rx+4RdnVOWrtMmaCiV5GyLnNmngp/WTH9iw5ZBoKhLoofQ
/ebdLlF4lju3vPeiYkRunag1QLfKLFeKxrDHQGjfoA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iZUdu6JR1PsDasHWxSCRSRaF3ttVgO9Z9vMGLhj5bXRy67aJtRwufddvia7G
04E5c/aMoa1DT2hDMql6Qc/Sgg3ffDbAkxL73KE2jRhy80SGeJKXgsdWpGCI
5gSQzOVJnKcCuEY1JB5Rap/6HT5vHQoeOZpM0uUP7cxGE6Yd8Tg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gaaZrD2W8P9Q8W96zdHg9ZmB3XBDS+BWWQyZc/MJLAxRTCwotqO+sO6Zk957
JGzbmOr538wZyOkiBxUpbqi4AKgy7u2f5gL7ZQiO814ZU1vxVOoV7cMnE0h3
bMVTCJAlfKlKcs1t++QUusme9w1+/UgRDjaWsHaIascad30lI9zsWn7rMNdO
0qmC9AOs6scrWVdMS61IWVuQxUW9gaIaKt00qeLsJ2ic+J1szqE/I4QzifTb
ADPUfWcezh6SDolZyVfGfkpTRSgAcH1ZvI9bZ07rEw1VIvK6NzPIX0NYI/fu
bnhcG6J2+O8GNz2VaKCqX/keq3rgPS+suICvXEIDPEKBu8lGpcWRHUrOSiC5
xNadPRSdVKv2A4i+LQ1tMe2R3d+hio7OlOZPGKODzBw/LUq8CLAag2qBr+DF
CNhzrE/IXCX3+v1PxhryNjWRoK5Jwug0JyHUd1da00MgE1KffTxDFr2T+Q56
IOu1rHijTaY6oq/kIJObcnkVkmL87XYT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bTDGWANrsqW3Pu+6k4jSWDaipXXHigCEOPW7rpYhHTa2bK+2nmqjh0JAXeWd
rmCYJ+Atg5sR5Ma4XRpbMKTRQrvVX7RHiYfJF96FMwuNfcQhKBmoiz8DQlVZ
1w0UO5MnPl6GIF4THwNgjZvYjv9ao9RUI8BphhNnDmTPe5CXLT8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ncVdTHiRghX/dzwqCoxb0X4L9C72XXQv+xA1reM4PTXxZUzsfUI41pxkOafG
jOAWGfEN/UiroctCrv03xkYnWC7/A1vZrsIrs1Zy9NThs+sUZwnANEdAry7B
CCXQwh0v6WXzIShEIjqG14aRom/bqLphtdtqiBx4d6KA8Km+CzQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1072)
`pragma protect data_block
GJIDfcEd1KYZGx9La/TzR9+moF9tU1g6lnb0vQYG7DPBZyovxhY3MGvvlfJ7
xIBxF4n5v4cjO7BO2lZyEMlwRzgRUaYpFGs3ufbl6+uw9woDk4WJrWhD78ie
eMsWrk13QbDAn2MeEX3PblpedxpvuwW9HPLVyVeBmPA/Aad9ePlEiCNv00kv
222D12GaEYzNEIBw5yU7nvbxQyh3GN76uacJpSxTRh6E5ITCxBDaHuGmBFYv
VIsETIzFzauNcsuR0A/ayErAvhVTT69g7UpqTxKkYi2BpSdDEW+0HZpcnXfF
77FEYSkAbz3v7llljAqRqJQ0Kukb3k/YXGX2gs989I+nnFA/NJ74A/RNHWWD
lNBfLWgYtMp+XK6cb97B4zLlgJIzob6bOAFNqN6HTciHoHQiW3vz3joPrBaE
7eadpXRssqek4zK0ggmsxJDu3qFsxYa9IYdsqAVh/0nDbNtgUByNCsWUlqhL
sTUOUbYrzD2znKQOggy4JLgr/gY+3VYf29k4egnNy7AKbvKz9h+qm69e1ahJ
QJ2Vb2Yi1AX8aCBbxoqvZbJFUgBJLMP9uXSMiaf3uOwRhE5I8zsvoeue/8ch
wMduBosMNC2QIOdcMrT0qi7PUMJadbplG+ctKZs+u37ixYh3Xzkvozosv62C
7w16IPsouJDZl+HIFXd6szcoeo5lwxuRE65nyy3TvHMvXdZwo69XiD4HA+Rg
oRz6Ib7vj/SKGJv7bNy89qLVGHy3Qf5HT70lbMMGd3t0xEix/8RMRbpbAemJ
GirdQIb0xQJtNeXOs1GqSTpIWin2xMsKtj/KjmfHayWIv7vfO1vtYy6tAJpD
nlLt8TKpRHymqrlzExiYaBoHjFjKkR3fwGAJkByChnP2/frJNHmV9Vuoa5sM
FUZdzutR9DVLOohq27Fz/LGMPJnrGn04SEjfDePGSnUfzvDG/NHp1OYmtdQ1
/zcJJrQDzsUnIGUwbxLSmKeLasLux8r9mi36S20wQL2vOOeVbMKRQrTq2u3H
10nLgo2V55nRWBHJsjLKeiqi0nZOaHW5t2ziDSoqj31PFoP6cPDfJDC5zMNH
cFnuO/q17qZXdzKUgwWzrlZsKFKob6uhlaD7cZM12//Mu+Iu62iuQjZADj3f
EgOkmsPj+r06pY/nVMS4ND6TmCUNXBcGpCI2uAq4BtHNbXqoTkpsukLbycW/
g5TDLrWLVKO/meFi0EIaJ1gtSc9lsANVIkcc81pWRCVVQz0GQwRh4vg1YtOu
KHddBbODB8xv4CVxx/K2PblwPFmJs0DJmiunw4K5zJv3G3HrrOiOLWoVl76m
HG6j+p3IXtb9eDBTgdxfHWK68gsYApEIjrx95F1eNcZMH4zBx0AlYPGw6gam
DiaYMS5ZRJKXx23lUf6SJcYBDSks0socDd8/TZzebpRGenp7pQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqeX4D7DFK2g8lOymgG1VAniTa8OY49AvFyFrPX93FTnYZA+8DuwYtWMn63Ku4Jj0Oq3OMbMXTYmWb1ABs4t2KmqGgd3A0NzrX93vYy7WSD1Iy3EaNl7S9ZEq0v5Vt+0IWX+bVK9O7Mtzf7OVmkDMzW+BcC6ti1jQd+NtnyX84+uKUwAd3AbQODiC001R4Z+qZglFhvZkgnSrxWjh7Ev26c2r8L1R13nGm18J2ednuSr8xyEz94BlzANFPM59fWFDdrYHrBskDehs/CIzO3aOxx+NSOabRjpnb/1MBezxXjicoCWJdxQarjrWU05/NNPNsz/BFLWlKjOggspLuXo9B+I3mJwnCJtuBHhW4kj+MeAmoxdusSJSaXWu2sLreNEyrz2tHYClpLo64TR/ovU3hPi+tQLs2PbdEnJWTnvGFD/qJXWZ/t7fGYJO2BcGOz/PN/vzTy75j2jUNkCO5f/tPS+YYM5h9yagG4yEu5fO6rq0J6aKouIjwkVOtkVJWJxNSIA2SUcdZZMz3XRAwB930VWFD1qB8MUMqHCyB2UU+T5q1H6rLZL/dHVUGLACE8ro+P4KlqYJfyGeKdEveSExEatHfhAWIsWHhwvv3U6PxHnpuHXjzSUTRGczsdnSQqEOZsD9t8Fs+3QXjakuqtQJvc5ch0RaA58l4sEtlmd+BwDoDH4LIVVBbGM5nBUCD1e8steW+n1F1DvsYgWOya0pwkO/Xs8U/641cd1Hm05KBJB/E8qqKYbTFngT21dI9g2DyjboHzwGwq/bEuAde0eL5fO"
`endif