// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
v0ExKNzRxCMto4ZDRkv8HPBSwNfKBExL6TI7xJJZKnWoNlLzQyhvN8AbMbPK
aBvWcPIL2tCJ+GFCatu3wQmfP2yUEmEW1n1Pg163fo1aj+/0qwJFqxUBVmMx
uN7rTV946LD5lfZIVN+lganUV9OZ8ZJkLnUcFVQ9RZL9xx3v3Ltfp+OuF+1Z
uxXN0mV/BY9ujCyyu+3jQRB7bXVaLIw6TP6gTmn24FOan+N1cwDFDZcVhYz4
4I9uXB26Af0dLm+ZcMDYI8q+ZZZMsWgZokoo7vzKN0u/EXkcos0J6SL2//BV
LsMtDaHzbUqt0mbIO+xsgNPPCMQ8sXMcfylqFD881g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fwPM1hEhsJ5uT/SonYJ4h04gt85wCk8OYD0jF0w5J38UGC7m5t+wPx6HfVzS
9PzweQJLUecM8umu6AHmAEaqO00RdobI7DCddUvjcyDZFiW1wur/opohuk+8
zgrwN+6Js0XPL3o3K+tlMnS1Ybq2a7VfIovJcZi6Gdrf+TEl0hoRmzN0/Bui
kxw6FPe92W56IEE+JM03MGJnbPwARS+ukBQTs3JJbRYMGycWcIOPsqFV9uru
ZSkkiYhMl+oInhNxIMtreQFXJSI0WlVcpmDtv21TZkaTPYtFg2UEUR5ZMYGq
O+HeTdOLw3ROwGqT6Mg2UlgdjbWPL4pjSJznn3Ou/Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RCPqLITjG6PUqqyy9N+ncNJMhKz0XHvke6kB2HwvBi3aZvMDGZ7hFRnW78pP
EF2Q4+DBs9me+Im5i6CH/rYonQR6wki3hQWR2mPkK7Q5dGqq9U3jhDGGXTTS
D5IU/W4I6H4xg7WEWPrHx8l8AYFJ7EllagsZvGc7ESc5AkPrggUPNtfaR+RE
oPLB89OYpzS80JCbcFMvTk7F0M2JO6KUAsudYdhgeoEWv2n/U7K6zpqaDftj
Q1HW2PpwDUX3GyKItdGBfPVrS64HA7UWACjokxXLatESXoQSc7fZGy6oYE7T
ALBfIXRtmiDnkBf09p+gfOl9O6+OWqBmOhY2rIFwDA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mFmOmxELz4maLd5ZSzaxPDUABQm018IQWxOzIITqieQPEU2Zge48q50sT/Jf
NwkdGhUyrkxJ7mriKKoZS4x0zyLR3yuyuQSsTl7wVNxgF0cXN5ddcolNxOrW
+S553On3Iqlx8enBhcNV7J/ysqMy2I72ndyjlNNHC9fjmyaAceM5gswO4gIt
wqhtcQjgYbx3UW8QyAxX+sR+jao/4rBPEzemCfMjBGqIGDUBtIlXcAcXgIoH
b1Pzk28MUzgQsseC99o0C+xQR5l2l+x5v3WVNeuY2RtLDhofuVgcOD7Kigl2
httO3owMFIXLem0VO95rfGrWOzAu/jbO4DWK2oSe6A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QzQ5on4eiRm9hQlzj2hroY8M8Y9NlMPHboB6X+OUIfznIKvMOdYSbzGlGXKP
+w4iR3TXKrTuMRjZVG7g6ATNLVrgFssJ7x2eleoNk4gedQYth9lW508Mi0ta
vDa8oU0M+4pll0HBkE8YOg3xFjSwTFBi+ye9AwQKrsRBtnrGGgI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VQ1nNB+kj18cBAMeNf28IM3EMu943vvw6OxIg3YDtK34LMHxBetIYJPA4iAV
4RlHrpAAiM7XNeY99Gg5TPM7UGTnJxOVIyQ/PIeB6BGMRXvx6y7SRYFSHS3K
s0Qoqgw3ubXPy/3SP5l5KZFtEHMdpsJz40DqLeho+ihqkhBtpcoCN6jc3dlH
mWrgNI34tG/eu8v4tLitau+hfHAQRA7fgfeV0kn5PXp+/tWIKdfzspixLydA
ANxGf/qhifISc//NW9FrERWvitdawDmz2dY3g5K84xkRTnU70HXOc5hFw3QN
OqfYciMBWjYVp3TNkKbGZQ3cNt1eXziVR5xSf1/Cdn6NEg7JJPuYAKLuo/HB
PF3vbA4UKo3qSuWMWxkWtNJpMh/3CziT8cNDfz8u+ElcKsVRLuMAEgOAXWt5
0cTSSB2TXRvoWjbuoapkWbFLO7UQWHfkrNFTtdPNflwxzNl6UA9XOREa19mR
T37BZ6SsOISN011rQzEKqKP9sa9QQQkG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nr/TbSQI2PJ1daVG2jPh+pZPz67n0QTkLYTD2/JYzWVB15qcsO26qmiX8pKw
qefMaO4YnBvVa1/eeedCg8h8D0A2xftYgrKhinS2HUkfz8EL7kLm5GzaGq1w
nV4vd3wpc1gSLnGkYrLPhrqFgl8FYcbGhywuV247mPAWIVpZ93Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O4MCI1o6+TRII0r+KykD62KqOuZ9LuWBjbsIPRd+6T27gJV6cx97cBUQhS4d
HoxCBbVJN2KGUY1U2ymPNWihDDDS1SLjz734umYnHppihXE2uUTttlKKYX5g
bLcLQt9IctSy7lAsssiL3CO9DsNgLtw/UBZNtt5KJIyYk2yhFKw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1152)
`pragma protect data_block
E5fjctfOvUeKwsFhfkKLZtw72/WiZHQU/MJvWDPGJbtbSfWUllporF4x8Mz6
RJDgTNPTkzIsP7EGe1YZQgIjyWRyq495qqqQn8UOZ5ViDHr1Q6nRVgyxobJO
GtuAXlTapbytR1YVn93hlwjmSrlaYQBC+qmU+fC0jrz7HNBBb5T72sLZM87s
56j9KwF/zVtxxSohCtc768T5RYZsMBo/OC6qXurAH/ra/hNT8XAsOTv9mxxJ
co1TOEhS9Yrty9MUTuj+NIsS/BM4tvzuIXmCrGCfC33yP+tkxTXfoR2XiXfn
6FCgrGN6bBFbkHJFQBITAeerBIpwQ+yJl3cF/0t3m2wEmPCPCpdMPAXibfhw
di05dfuO8n/24sn6pgiMHvDGMY9W/lyV26Vbt82CAwIxz4cUM0cq98twj53S
hMsnwQ/1kKH1Ra89j4WlWiBgikROt2UjWHwDt/gCJTzwPDJbDn+md4ttxRm5
6qfN8rQDENvcu6i3X7VUVe8+Cv55Jx/7SgHK9Ge4tKePJzfPtQMAjBg3eO29
VtHMV6f4Ty7vtFo5uAyRnNLCma1SnWWEwvSgMx1iVrA+Rjfow3u+3g3YONW5
Us91797h4ApVhdbZjm7V6ixsMv51oiyRhiybjn1Ucb+hSunJOJ+gvI3F9W01
xRbXQukcpeJtX34U9Jv5JWs4+DevGRXR11qfsDpVs8VbVvQ5/OyZz2JAxzPQ
POR+M8cIAsj1aD8bpWvJg2cxOxGkanBSjQtQ0ukkH9qhFaH0hDGzBxbjC2aS
yQMOqVO5F5gB/YduK5mioiqv6HiJVPb8NLDS2YOvvz//ZRMJO4kYG3D3yEou
AIr4Hg/zt4UPX2Hrz9bQ+zckSE97txn2wcjdx7Ukf/EfAFlItysUMN5Q5o7U
0miEZekercUfoBqMZSXba83ueOD3EH7fA+f6J3m7WSeR/psxHFTH/KXNH38j
oy/H/QtN7pXt4vmGDnTi5SEPJBCr7HCGwRSEQDLZHHpWbZss3kTbuY3Fqmlt
F+mfuAcbmHqfiPiL6g+PtpM9I4vnUE2Sv0w2YqTswbwNTlYYBEy1E5D1JaJ2
qM20Yd1QBOt+e5lHw8uSNP2NpvGLV3ty7iqiezC31cCVY7Jd3EFakPWoat33
8x9FfSvqkYQGGHqGus9R/+Kprqa5D/Ymz6tqdmnSHzMjZcSgr6dLMh1W0CIQ
/bnyWlcyAK81Js3iNsBaLm3m0n09GsMz8RHZV+vy4aDCDGyLYWv+8Q5vr79k
zrTVpZuqLlEwf32PlLiMs505IXty13eIgxpV7mV1jgui+ROFKzz1IvdzEsj3
n2CwICjlyCNryF4CvfuBwiWy5hQcj9bTzsxPPpzCEwhxjv3hwoo5CifP13Nz
ll94hKu1u3/7zA8+GWrgCrG/g+eNsNgccXq/Q2kWygLa70rjg0ur/EFZgSAf
3P7S0lYA8B6+Z+IlliMlQeBkCoAsts2zCk4J6Ki7xz6DKkR+SgXPYymkGeZO
ClMYbv9jIyZHxOH9EquY1hFmGGcJz+Br9QZc

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQozsYK6159EE56uCf4+5SbqJmm6TRzSr3eqLhdhBN07cuaRdwG4xzui6DBbAnNcs6gDYFpQkUbD4LmDBhbaeDlmgqX/8mmfYfgnF8BQ10d6fvmbh/umBdClXFJ6SVK8dPesabLvZyFwKh++mDmm9F7h8wRB62xmG91ln1swj42Eb0U0MN1eCOMRuOOvt1LnWHf/iWcPzm+JC+f3biqwk3FudoHPeaAveifW36nqBXGgSlSYZ4LIpHQWRGIKrDeZLcIYKuhvuOFHzTBp16X910PVeQe/3YLhe7LxuAUzVIuZDarf2VAoXr4zUJrBSJMhJkQNh858nAcIZOnWS4GnpNiT+2S+UdRG6eLdn4JUopHSD7TKyaWiE6vHSd52lQn0B6PgM1uuoWliSnzo6ma4LUUMQd/hDcWlkC9sbBGVpuF1GeZZfUNk9sA1UJXMgHesUfBMGdeeK3JMWwQzZUVrQKls3Y4tV2ixae07COGhOajWyMZpkrIjJXtgnaVA7e5lydLNZQkSfeFkXFxbFAAW6WwNRH1upCVFDjZ9Gestyv+9pQnEH2TEeHboC32Y+0HBuEOW9EF1pDstPlSMZDsCXB+SSziuzS3QrSfWNVtcfRWiJjH6sOkOEhNg4qn4ofsJP//aj20aw1Du/bBTlTODBMrnwTGY2qhF+v2zurYHC9keUg+YNQtC2QfpP+DU3tylE8YLiK2iRmlU5uSyw3GT2zueaq73uzmMZwWCp1gXKzpSZzYs5Dsz5r96UpJiHH0bfh3qD1M03IX7QgPexO5isNZbE"
`endif