// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ruWnOapMfW9rpkr3qVtiWgdNH89VPWjc0jVuzMegwEUKEpYr4bFhYVF9GEn1
xo+0nqROvAoYD5DdC3aW/YVZy1ZXZhkOboiV+4UF8pX79xz53Y8tlwNPPSaJ
u4wJ/OpbPpfau83sBW6p+1c98coA1LdL3SISFqYjyPfEfeUPli0ejTq7+aGp
NfAcZEc2NkA0rsLd/rQSk2AEgSnTjD0l6dGj4WaGMLQvOdV7AGvHZRCvd8E4
uqpVlfRimPZ3hnyfJkdoWN+5+eo4tHilr8M3nAIwEyiaZtV5aef4TuOcjTwA
t7ewP8v/C/NI38852soJAElmrZ8GBzLi3a3fHEypaQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ique06UIsScvqnTEvyDDaA0ja7IioS7x0NyX5KCW1hsy1+rh2BGEiYWRgINq
IrIsS0v5HskSAC429I7Dfn9qJICU0kV7LXKpQU6CgeEhqtA4NUxXUcz3Elro
AFDH6l1QHEmP/H9+VoHlsUH4t2aPRkLghIGH6rGnE9ecJ5q8ZHO2eNr9E8G5
mvVgP8nL5gBJ/rJqoSkrDGPG0v/xktc3lo7dglCkvCv0D/FB0ZvvyOq5MyyL
H1t8/9mPkJ4U0GHpQDT/0yTqW3fkd2cXEXVjXJrEmgRnt/Ehl544FW184OXp
+oA+Os7iF7ZJu+nPLUbk0/YUI8fBJynPGymawj+aiA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J3HYVme30nR0KXoDYU7QpQPCQnShi2hsNGs/WqDfpnSQpc2VthzB7wpDatS6
b6kmL9O2jLhLrKwFXGpVloelRG0kBOa4DSXlKlWHXLZLVSiysfXHqlDBDwob
agmz0HgRDQveQeaq+g6HyHoczKOrd5eABTqZ48pXa8NlJMF+hxZybLTOiVwf
9LTt2fQ+qbaz7Gfus78Ai4XdAliB2JnGyYlSTo+6iFHoT4DOmEDCa9IcwP7F
FXoEqFJVr8UizjBI/aHO9Y59Fe18XWMGpXaGIv8uDVjTC4OP7KzBOpatnY7i
gY2GDHgaXAojgiwhj8RypYx+Pi0nXHH3aPDsAR+0Og==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ebg+ANDHQKB69BzkpFDo+O8UTlYsgG/5RJ/Ms8w7XaR6pTQCGKe2q0navbj3
0UEt+nXGMnIT08+SzBWE5zGXg8RrRIOzeB2FNDoGW6neYG905fT47YVqgB7r
SktLrY/L2IVO5gfzexhMZGeOKHx95d8KKViwhdE0vNcry48DCE90J/uCL/Iy
xEyGh/QuaMbVRjCAIFYg8a0zFs+yos/yJzod3aBLWDOuxS+s1wB+g1YJJMhB
E26Z4GDh8uKq9v6GbzQg7ecI6ClWqNEQJqgTehcfj3xlhvjJslubdgw0mJO8
5YbgNamalNkMg50+uNUxPxGv6gPpiDjjb6PZrHaVtQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MGQqTXnTRUF6nNYWP+fe+HDbgyF9ybv/7dTAHGh9mCJtskiE3PMyMujJV25j
N7n8pkx85PDX+E14LYL/iGJFiQDN7tAfZ5fz/5bOj6qjf6ZYHRp2mCh+p2kV
AWFsC+GMBMimCWLx4COqvxnu/u1lfWEp20HrlQM7iC6sNWWP+M0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LRWAJ4JznQ7QigL5NwzRXp6NC7dKcdsPiuIF6+E7AB3kXx3j22kWrS3zuJVx
jBr2MkQrlZd8GnL77/HTllF3sOmTBj/qR637pWY7O8IwXB1vM7E/iK8ONtqF
nq51s8VU3Az/ujb24A7X6JISiOX77E+JvZhYkoTa9ABXGKgSjsN1HRR/zCHF
jShdvgQXOQZIP2A7FQXvCCdqkNgjUUSUvhjrDJ8cVcapuwhjbkSNCj29q8Pq
5Zp5lN6oOpYapOdUbA3y0kA2rFTPDiz+fqsWrtPF5XGREr1WBXjzTgWspiw/
uhLBI3ZhvMTQWkGF6WEE91CAvsCFgUoKBxLXGazATNairh7SxM8Q8NnV3BRm
CLjpGWwtXllWVwoROnLzcVW7tAlHNhZidOsn1z7Ibq/az5f+BhCOnbygs2yj
L9RoXRlAsbPuhzzmnfbyLF5ZSYflvjhE3EOxyYPYcNn4FFXwi57VRcSc9vdq
r6OuEovVBUup+Xivpo3jnGfQAM/KFkYx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ui0PQR3ajD1ku0eTLmGlU+bUT9Tt/0qwBoP53P0PaV5XhQ3+LQoZquZIlbeT
Hvr4F0gBDC2xOneqvzvqr7K+/5k/5hgLmgDL869VJcpjy9SbenXbEnHoQa7N
7ZSth6GbEx+Dzg+7n/sVp2c85F2NJ+eAznPX9sHg99MqSV1LYKY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Mbg1zZvJ25Wa9XIA95y2eEYgDNHiqcNfFXHNVJjKY7VlaIHfZPz5CuYn4G7g
rvO2wTVtbDBmHL5H44qpvlQiu4vnTstf+fGeo5DPlF5i79bmmKSUcepNId48
pvUZz/zgd/OoaFFw1ZLPfPCcsDRt4II6b1JbyjqHAS1Z7LTNBYQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12256)
`pragma protect data_block
6Th7MJzrYIFQl7gS2QoFuANBuF/D9wkWKSDMJpUqsDmkjRHe3uguPHWQ/+Ci
3kJ0i43FBuioCrYhHtYvjbbSemzX24t/xRG9noJxyp/WE4xxce+6+Z2b9RGT
2+C1I23yUBuJAlRnuCo62ADIQYdBodpplLn+2+vots5YaaKfwk2Hmak9qRsp
6bNwos6ISamPdEOH9S/uC6wLNTVWw32QIwmLfg3r6Pu/jk4rClsI8uUYM5o4
4kce91u6ScX7kWNriXnzuSe1fC2LakXTVaM4wfWt+Qf+Rk1bv0AIpjULTr1u
2DJTmRmhU2S6iujXvAGLKmv6RYQuODJEMbC8P4TFUswkjuWf50GoKP2Fj82m
Q299zGJ75Fb151oWipg93GJRa5o8UVkGxjh3a+cWApDiuVGyUr8Hs0+Aws5o
F8T269Dn7wDDFIB6zFNnHRbHh44/8LypiHpp0a4YWPn65C0PumZ9gmk4k7Y7
9AwtN1cwENUmxH8u4ngkbk5hEJAxW4uayK7LMbdXTitSlHFDfyThcHJ4dyip
0rg3xVCPTnyxtn8jlBRqQFEc/3QIf83iFAVL+BT9viiz9QsbX7JxyJwB4H8V
e4cXjEf5HOa5UWHnbm+S5/+cAj+Qyrb80sof/cp/+eszuFRYztHH8aYsQTOh
F+d1ALOYcYjdBwrxORZ0miG7Oqdwrc2ZK43bFAxCR66FldPobdqMuPfZ5yUa
rTRgBd7tGJnSwOJrYlmKsgaLcHSsm/LetJL625vbtij2Luv5qP/N4vHk6uah
ojkZWbEi/fRMZfSZAd4p7vcdShsr9ygeu1gDX7cBV7Fg/6QFHHQtH6H7Xly7
epXDEWB8QNRgAklRD2AGn4Sf4Q8KUElPGdCrd0bPkqH4zLMjlE8yMvPC27pS
K8/YJnf0W0WvlFzA10xnqsIhv4KzYj9nHdmKg0Z7W9yAtIY+deHhfpTuutgb
/A2x9y7iPEdCQ+L77ZbUMLvD5OlihNoqnxbUrd7bm1diRnfd23IFA1jqY7CR
Z8NrH6mwpAXgBuQDXLrv1W4M7eaYC84LGtyXBhakDXIGX6rsItk+bTJUpf94
DXLOPNwiGoR+20DCUubfcxIKNM05SayUPJu7aR0e8ReFxyXIuGbwogSWq2dD
KnDnlfZPVmhTFaVCRZK6NpJtclRwZslzTN2t1PArRhYJCHeVObOlSM1VDalI
LTGy0BD0/BE18Sxl1QkktEBuvPr23Giphf6Qogxs3/foQpLU9NNKErB8eHYa
j9e5q9Ck2YfiNd6rJppjuehthQ5gJsUidC5nP+TjcdAF19loNqZBag4ZVIo/
i3RtlMp6d4W0WPrgPBZUjAdEjENaw/x7Wj8o6xyL5XY73LO++6JSBHYLxE5m
jVkfQGzI2BxYsEeiarr2knr8xyIw/E8y+Vmvwp0ZJCFD0148oa/F7Xs77C1M
V0aI9wGT55AvzgqU6tXUzDUldDaunzYpycVcPam6TcAYqSuCE9YJLQOnRa3A
SupdL42qTakk4SWyhIEfU6J2m+xvmCCH3/cbprDRucg/mI5/dy8DqpDYFTb7
RWKpewA4bf6zPrwtT2y5oTeJFEiOOI3T8FVtk52q3yfC+1dJTnbmvON388qs
GOhKavB/22cklBt6sxrOeSOsrUZO4Y7GUzdgRUR8pU/FMZD0YtDAjL9OwjSc
VMYCdagolyzAt2g1FzKWvsivh/AfH/RZ6YVqGhqGQYNoB6Q0mn4OkOWmmYrb
Y3KCr1uU/wjas2xHo3Z+yPXFUFq5EwTcXbtrUNK1FVdxZGaK0rnUIN+b9WA0
hap5XG/kGqZASO1mXRUF+hiI8VkF+C8BSBcVSzWaKg+0xXXdtxJcAu3I8qmn
Rc1vYUtdOufBTLm3PUJF3nsJMlhEAHScyKu7R/dO/YXBHrAcai0pzhYpSd3y
PCfYYIZpEytPfOMYPys3m0L/tIwQfdm5fwG8P4AYwcoulLcGmxPzvke4f6DL
78OJn9uSSOGuVU+6+YZ4hUAPkEbiKfd/c8kvOgtqGjcEN0AnChJfys3U6/Xe
EUEyt4k3rSMowFHfAjqiCzTetmaKi7Qg0M1pRGF5Sn/cOeGOR/PhK9jFMLE2
+oOGFiRSkBn65a6MM2+6Aon9e4cCtDADpuCKGjOyRtrHmk52TRVoLZcUqjK1
/E9Kzja2Tm/5uHHrY8izukMKisIUH4uJei9FKnnH0FPvmDwMVv7o9oOxqpVS
FPuRhac8MvIsJggzGZVaPdkPioMBQSsEyY8F4JZlz0thppCHJ+ihbIF20/TV
khXUF0uhbUdVbq+l28DI2wXUAyzdAkQp3a3YfgxCdjIzzAHi8dT9GFal1xdh
eU9vflyDDY8QGomyM2R1B/A13bssS+X1EI91ovGAiTmCVXyHNnXglchh6cc2
mIKfqr8W246hMsQ35T54BKYgOv6aTj7rPbywU1d10q37WKgShI99GA949poM
68bxrPGdrRIe4i3E7FtYHC0Uq+xTDQkYQU6G3ItzO4IZ3K5HbJ/dpBGdW2hN
PLsESIqDPYGBGeqtzsH6peBEVMPni4uZt+XI9Aiv9GknghdgyDwct5dhclyT
D5L5+/3lni+eUzaMC46ydvVrzZsqUOEjyrWNQRUW/G+L/o8n/PBaCyQHjYCn
wUxPIHbcNaOLTKK2xU8RLsMzRdiQX//K+t7EbBss5igM235B4f5yKYXrbL+C
0hnHKcN+NMY7PgCttO62KRNzew6rXNRoGl50weJG9YQb7Y1djrPGi51KHXJk
rg2Y8O0zdoW33mCudEtNG3fhYdIkN1/9blvwl+qxOBY5Mkx5/XS57PNaZCPv
bGPwXgX0KWsxfh3Mbg/FjTOvzJWfp7q+y6Qy9sHFLWtpr1138B9X43O4ZLYZ
JuksWVtJi2VsbVNsQlPrXtDCyeb+tUQlfRTfumdimCpDCS+LWhQQxLGWfRMV
gJ7fjcciNmxTJWyiozPbcXZT0kzKkzbBVhWsLDYRLrHRI5N+d47iE13Q93ej
koFN/uRjAspFtpj5sjj4TJwqe9PwKPGsHIhgiFYpZevNnlaQwYgH7+ETYXik
jpZ5KWjwBNsPdXdEU8HUN/umAbRJu+Lrpy/Fdo4dMYft0xJExhk2ko76NvMo
w2UPXjVOPsFK6Ukh5hBPxvPYwEd3of80GBYvk3/f5C/Zu+EWY8qQaBASw1YN
7nbmYhqxFztVs43O8ghBQluvW5eyROta/UGf8cQ5MCAakn9WudL86w4fheOQ
Fn20pQC8h1iSnnvLqZF5ZI285KPxUnSMp1YE8m5IjqtFcYLHnKUb+sdcRsqT
ARuhvFfAVFoN0/pwXvb4wfObe+sP8e3fCMq+ddIiAZGAKCV2HQGS6KEB7FS7
+UYwHYrIC2C0H19dJ/SOsOl7uypfIqyav+8eecYm62ACsR8cOZbKbNkwn6Sn
93fPze67ZcpmPknXTuoxGt6ZCpv1CG2enwhREuEizqSQl/ut2/STiXCnQLlG
DzTADAWu46477wHjdsVz797Dc/BlnQNG6ErFTTZJXIdGM45rnhWs7/cttCI2
bHj2elJRixyBA5IOfZB08N5LJRi8nnM3MbE8FESJN2WcKSb/81rNeclzvo9H
ynBEYeso7t8eGx8u3RXuLzzlGUrRQmnKySJOJ/Swg0JnxjWtAuSzkCFemMk1
ezU5MHSVpbFk9rN0MoIN+X0A0+MmTVQIsg2r45eVcbx+hYN3hLFmY5zyPOVJ
6T0SfnQxUk94efR2W8sdz6vDx1AuM1u1EHCJjqkWQdkF5EJOLTfKXdaRufKG
PpqExn5CPhHFps9Fb+PiEuEzX9EML2EbbhOTrYJlzPNda3GrwgMPO8DmWBfX
1MvxY2qdPtKxmRwZwNHrWJ13m1gnBqJEyZe08X2Ruwd2M7IFyC0K2uCU3a01
jPJAYfxQIm9mKsxZOMGXYQBI9QSBUFCxg0Lhw4m07M9apcGU9p25/00gXSbB
c5yb+loeIq6/Z6foCQ60WEcbU7/03t9ZrY8F6SJ7a//Xr2nP5frdrjWWpmxX
5FpBBNmIyJuzTx4vMB4E3gbE1ZPAhNrI6jOnsOFIC46O2Vlhwlk06f+BT0ay
Xr4rPcS4EYnBqca1LuEet0WAeZmjz0TJOuSv/B7d83Yp0faJMpD/6HDtbg/b
j3kDUE6Ijqvnk+Ks1YgOi34Mf/vbgzwbZbb+MBy1P1acX3w0v76GQXtaGD72
ZoDdH0r2e7y+0Yt57Jfrx2UpbNKE82e0pXKdC+eYvMhWq9jaT+j9shL/VdY/
lU5V/OyfxmfQ0j6mcJ1wyrzPSFjRQlUqIIJcDtfN0hcGtpWf/Pzv3rk1Jjut
nIQMpldj0z+cU1Uo4uZWlW5VmZUFRguRwczOoO3tLr09UVTz3Wmd3eppWH6x
ymmRAnP9PcEWo6mZDhQRcsMaIQxeCyzTzlmWG4Vx7r2wCJr/+eWvlPOzJQm9
MVtCXQw6IO9lhGzaP70qhblnDN2YFoOnv4cFnwXHg0u+fRAQ96YXRXT2dVeu
asz11EL/clHZKJjKzI6pqDtHNKrPF7kG96xe3pHtAiD3ZI/OkrttezWOZ4Om
NqdSeRuSa+opWdUTdO+pRXUsjUMkoSRf0jT205O+tRMGJZzfwBBuVszZjuJO
1UKmUNfDkbosX6V1DGuIj93wQ9t6zg8HU2pg05/1riX0z5yXMCZLKgjDioVa
s+x7VGfFgAdAHBVkdjt4ioiCGNAg0FdlP/jvAnwVV8xoPZse21KgHBmDAAIg
XfqAeDPqZ+bcQwBWEyS1WcHehsYILQ9NuwhePGTru+hb1sGSqKy9U+MTvBEW
snjuyZLoG6Fnl5HG/P6AwsUdp/GuOQQoYk/3a3l9vx5mNLdZWvMgJHFw4PTx
5AJG6aTPKU0HZaH8pSeYwwvLBGEW80+1q8/aP4NOf5gtrn/TUYdtoRxemVXK
4G+C6YUEIJGi0Ku4xeSVv2XjqCVfJd9vc2kuncvt64QVt00g4qsM5PTo+YEb
BVlZkrDJNAc9BSzb4xOmWDQC0rNofxbLzl1fOcD4ickpzRGipHKG2aA+u+m9
nNVbZG9TbKVRcQ9vNslPD7dTFCY1zpQSZ+jq2QZgwMAU0lIAUqj51b4+AcUp
5CU1Bxr/45RkPyS3fjF+vtuL4mt6V3bhJrwrwVsudsYf+O3Pfk1BEzgVQzUr
R/rPX4xX5ooOjCSA1qfGqFwKE4y6IbR/8BubUSM7wXW5jCn/4zh6TIWmhLCV
2fzfAwcqxDCW0ujpb24zThK/b98zHW5cpBzojEUOr0L5q6Fg544JPRPMU8d+
YSqlM/udP9nNfW1BZ/dpNsNK7FG6yqXRB4/eJXQO+S0v+TMQFuIZ+O74DrUA
IQL5ar+6I88qy8jKefDDznGf21pHUTdOq2qtkA1n9k0lcoJ3s9YTG/n149ln
Cr0oWu0e5A+5dSuhVfXWa//8otW7bGYMlkxKUDqAG/aqaAF+oQsGuQJfl/wN
6cbHPgY2VkmgH1I1qbQv/PiPNmfwinpUSWquziXxMPtvqERcZwpMAPj4rkVa
0+nRGYX2szSkugwaW3pE4jNHOcOSA/03utTdr9Au7bzea24IeO8TKg47NHkA
x8e9Otvim1RAOrE/a738DCwVaLsywD0vTCl26g11Sumw8A7nYMeEX3ji7IKm
9JxYSfKkS8EAVfNq3YmxJklNgL6bXenfrpt0WqbIVaNLZrKZgZzdr/N/u9cI
NDfbVARClm0mgvq/FyjsNTV7kqjkUuUy0Zo/GLubmQsyIBrZeEL2uMGBbG4t
fSYEwuLJBjhNisnB9zKN2gBRtSjg+GNd+9IH9ex2DVN+WH0nBAyRysWlLvRM
oKKzRQEopkWQxXzpUK9pwHYEXsoNVQNZQ5OidBVflqSR6tbfKka1tZk+h59U
73r64hA7hOfRhUPMHoxQFt41Xu1YGMx5VaQuKqtzriyuYEQ1jZh94My64pSd
E+x4GjrcT8wHdxAXNzxVs5X5uh1STHqYHAMrUJLteMMS3cyiw/BT6qWTIuPw
LeFZUtpVwajP0RdbM4TaoE6MsRhrOlBRFFbHAWQdI9Tmmt10kC2BtuwJqmJE
3FzexOcqjQIDIJ1nh7RPsGBTDCqi9o7lbSvbuQt7mvykJDieWlYbxwktiJ5d
irX4XVRLVype5/73keIT5ucMivwZFimbvPix7unQISMcVpZ+fdWtNVuUO3jO
sZ/M4W+KUVStFof0jRr22ZoX46ebF51ADpXNdXRCWzt4N/UOdiWMj/uVSiby
QgUOnEMNj3pxkjmqEgZWrgxSlCCrRoWZeBDyZKvZ+am+/Dgga0HAKJUhqoZz
crRMROLI+fZkjxjE7j2Blezo4tygSqGcpj9cJOdMFDLeQedVMA7Jcnb8yinJ
UowYyTnu8h+aKalMgaYJQxvlL2BQoGfYojdU+Au+IxvY8L+tJqfdlB/U53l6
k5Y1tdx54QibmLv+rk+oLRCLSJQKh0co8rOiK4jEJrQuhD83NeTJgGyUrmmp
4Jnnj1fTZjWJllk8U/U7yYg2+IBzWZiHnl0sSZIw7fvg/6iAbxIsBfoeYTjT
hl88lB57JmHvMdy2EMxn01NBEP8lLS/6nKdN/axHt88Nd4RXizU6haZvdsE3
ox/M8AL/v9rU7SfnFeaZg9p8NhsN3n/Wo26f9+UX1p/itFSlKYfCv3Tsq3Ki
i4Ke+bgpbqTLMbOphRqm66/Dwarm/Qw75MTTwpf74FU7mQH6rUz9mLGGmine
Cc7DHTvqWEE14uXEbSZnnSGMHiRa77Ye3ZtpnSQE26YYxqnpnTSavRhrJqpx
5dxaZA55h7NFVgxYXLrJGA/8vVnxaneGWYqiv59OqRvgZBXv2sl3t8xZxKVe
ZdLY6meQsxnNcy35X2SDFJa6blPm7HXdsOf/dlZzB6CRR4QiaRflouna8yJn
/tcizAai8v8EBK4B94JyAG1hDcLNMMAy1GXh4eRFf6XVllyOAhgPA2MnqqlD
GAH/y++UE19L2dPuzTmnkbf8fCtuDalAeZHwvwnFe9S9C35or8zORwh1wiiY
yZ17brcvNhAqPOsotZ4ShCU6QJCNl2vb2WM1Jf7MSiPyJea+Z9U3aekm4dN+
JvmEo3vlpGtie5orGgS0WwNRTaM2G6oPUyeLpr9GNCCCtDNABOCbht4k8M4M
ebhfcXshQYaUKmPNQAtmzxaMYtbumo2qMLvH9HD8g2KD4DwXOVxohBCZyRPA
CHb73po2FX+E/VvCP7xi8xHVAoEnL8bWjFjr0wbeS0WMudY+EV+PRPJu2Atn
/0rzgeGNwUiwDclpkh3T5ODens8+Wokhvp6oQvs9ZnuLOX2WgQO9ITDhd/7V
DTEwkhitDaLxaseJdSg9lZ4kGXWPlYr72gdR1q+Cx210+mPbNHcOh6ptMfLf
qudY7+ZJ6dgtOt4KbjPbbmYusyo3cZrw9HTnbzFV7N7Z9IaOc4vpdwEyzNMR
MZ95fO+mcW9Orbom5zctNsGpnLHsjKgwjONPGOc+oYpJY+WOlqUEE/aSbzrH
Kk3XFrvJ3Z2Mhe78riJso0vCav8O9hqdGbP5d/8rasF8HGn3drXR+yQd6DOh
XxiDFnDjcb34aQp/sdGs2Ltd5SSN8iEnYXid4RdYmJLkPGOHPxpEfVxRNf4m
bH38Ok+2n2vYZJPKsT7nOKkNM4qSHPUz1bea+DxFyaJjj+ZfH3ntegyqhZZ3
oOu6mqF3HaA9oiyT4AEXvq+0dorpAn4bwI759tVXXweIrV9IJnZH/vtl2m5L
gqA/biekciguYKmQdPjv+qwfFam1MogXyF6G560aU6snBd/uVDkTuObEj9AW
yWqy5P+68xfeYZtkV02sv6VfEvXRccfr1WQusDLJJ4m+oTcJ4Xa10YHfIH7h
Wee3Zv5JZpNcbUL94xci5fu6UxeSMnDULUQWPxx3EAsnwr/VhSIAwKD1fC1V
8v2+Xmmkz4OstzAeZdgIZ+FXyiGtQw9mSyUBAMvL0uyK7agl/b457sKy0wp5
MOUJ9pEmzVJH2hOeo72Kw0r6On0CPyNLd5TY9ZmkDVZNxwWAtgS/GOSPuvyz
lVFYyiZgz3q+pyqN5CW1GgiS95AOO/rsT2AxotZw2flMS16rcQ9oRoV233Aq
FYAO1ifCaeuiSXqbO41VVEjiqAFqgzyWmNEE2j7tdFLjEZNaftfstJ9qYAIU
XKgkLPIJmQEMpj+EGwMcUo2ruBSaMyJN9hVoj5TNnGrW8PlDSXttXPLrfk9n
M/Xrpk465pOauq8XqzoIKm3zCwgK9lVg03rpToZ7CMq9D52CbwtA8iTwRIpT
2ROq97P/LABy3kvggWW6lI9sVotUXdif6iprKriSNYGZHafXe7EJycFmKbSU
ybbUPco6NLTEzjy4vhPmfoUxq3j6bMU5xdSDvGe6/UUbv5w/kKTvZFbWwJHz
rXyVbHEgf9rfrqVVukCvXSz0widT2V0GEgX63qeMUkGivinnNH17WQ/zzVIU
GSDzTNltnm4tcTv+obnkSq1QGF3K6on+f1hlfQF7GRI2wQ00++8SCj5iS3m4
oXmTICx6hrJXtftiaRvxraTz+2IdAP/rXfZq5ElO3v2LIFcqr+x8EHU+HOua
VngVbz3SvHgSIxu2oQs9eYk1rHfv8KWf4BJPf/6pqfplK6uPVhtbfG52fK0G
SC2q3zqF4G/fL7tDE0sMb8dX2/1yRK1Rr3XlMv/Y4KKvsyX8tLOT0tTzYLpl
cYp2JtjYpUzVXr++zMmciZ0uQXaUEH9MtfjnIEkFKXqB/yFMCxvpBS8xWM5I
k9kWq30QlPpumRtoq48bskaUGQ4emXtQLHCx/MVPuH0JHgDO5US8qC4tDZiF
2smU2rGAx7Rp+3RdATCyPnS4HULZNrcWItUaJC53znSR01uFppevHf1BUoCu
5ywI1MAizLTYfPH9WFiN2Sp27j976EWofepsHdRyY9xkxX7iAlaTWvnKAN/9
k7JmRuPXg6HkGZQU7/yWRUaCVb6HiRiK3+nrqO1/hLXEGTiEBj615NXYdpih
fSASzSKYr85Tg2dAsOvR8ah/80Z6Bu4V/GMynuQu/ZHGJqAByik23MrsFKxX
oQsBVRlxOAqYqSvRCoF/n7E7EMNTIFMKwMAJ4SqA4XSnOHUZrscw5t9kxYZ0
GzL5gq7VSSL56yfu9fdm/J3mTYj2FgWSMdf/vwk5vAx+VvItfZHobLACOB2Z
yHqj5FXXrJyzBt484EBycHg8ZwwSikFe9K4rWLGoe+NV/99jN9uzgTARqOWq
nqekx7k8kWMt5Rv9xjCFIlvwEXUubUxiJ9wTDSJRVJSxXrNV2ul3friyitSM
5qy/RloK+hcXojBclTlG2wltujYAzOEe/YtiDaaVjBnD6HciE/5FNRJheK1C
jWKk2tdfn5Askf11RE/qAiCPQCQFkGulmjjZfQf9763GLPk6iBGrGSd6RIU3
O5xesmJS9xR46FaODogDzGN1+or6Hlvhc0o03jcyBjiu1ZJBZ/DJai/YIbbu
97I/gVC4/AHEaP67HLIIPxuzyz1JXa9XeVAmB1Lk7WckJFG0yd2Xdvpoe48z
TZSRal3Ps7jBrSkvcw8UCSByze8n2ROqlpaU2zRZXLPkkiSsiwULz+C4+3zH
bjg8PbjGsNGohKO827Pgdfd88K7O7KXWZUl/bC0DtTUQE2Rndiuka0S7Zida
rXDje/1+BY3K8/lXcHqJXCG9nujP1HwMbp7Ro3lgurLFq/sKMCH+Uu23pkmD
S4XWxYbmCtDeT4AIULeWGdsb0zqOyYCvkTXuHjOYTmr25SWqqMWzYwq1VJTW
vxNTFB6VhZK4fUCgPSP4RJ7OOsd5rBTmrWKZGhaltOVaBZU8urv6jig2D8NY
cnXMlbk69T6cufG4MSlhU/bnx8/PcWzlqEnWhh4iqFLnrBFAU//Nv8qbFXkI
MwdSI9V6rdBO199rqMa/SEqEYxdQZfjid+iZUsrvmd9vmDQ7ZKPvhfp8JKLv
3VVnWH0Fw4urSND2pQs6E7xjudpkGCffJ3mS8rQz2JD8mKdc38oQduc1ZHs/
gIgW60Q90330pqJKZOZrzNDXYaKq04WqTcr9yPTKtacyB+n8oV3ClHhJBMgD
b/q1V1x6XtbKf2QqH1kGQb/zpufpIhfMnGzS9nRfzV0vm5SE6BhqujVYqHxF
05zR22bT+xrmrJjdNjRd7tb49guk2rT0CBmrNs3GJJw1Auxs2zH7hvTIVQM+
r9M1oBUfBmsX4F5GkuQBrJiKEUAXEk/Qq7M3h3H3CWuoKs+TzdfT0Rt1rZzU
NYZANQ0rSu3WPrsl5CYaJn0FaMXOjm8J4gCzlLup5wkIuX+5i2tTeCNmOn5n
9c3iEjJhcEfwxP3UyBSrkIGsadwdZ713F6/NDqAvnqVCgDXPD5W3cp8zr/A7
ctnp68FedEO+WT8+A2PMoFHww76r9lEHscEg6ihssv0omomot5dEkhDbZMq/
abyVWdTJcAm0lW5klv2ATGkTkpc0+nntqFDY15iQRZn/ueU6iWTVJZVCD29i
aPTjjDoaK2uL9rTUapI/auta3Rb107BZ0aT0gdnZO3CApvsYpPTVZyRZV+34
UqHvF1W/K8XLK6P4pxqXyR1eciLIG6a+MxscFMD3UGKS6qNQhkB8cFHXO2I5
YuyUBj8J8HVi5ZN3reCc9IU7uLYKVSnB0q6G8/VlDEfberVXCaaAkUGnNqLQ
LYh1/EASpjhIi4mFjBfHNWrv/e5qUu4zRn8mHoNL874GHlM237xYI8bGC5Fq
UsINCrCzN7XD+hfTp1k1aEUCfnUCHaiA6DVEfsR9mTBHJk7B+MiCRavopU63
OB4gN7Z/CfJlpz0XUPKkvL8jRGWXPxH/Qm2twLghXuPt+soVP1ZFE/x+SpbF
Utk/mlWCvRYMWTOI3i9vpF5DitRItr3vIOzyj3p4ykWqo1Lx2FmP3IzCB8h5
mSFYOpVnzVAkFUye4UfEU2f3FhJYspID2+yi+CkR0Yx3MIHJg4SCzXeO8Pgi
Ay1p7GNGV38igk1oAfbUfpFUPbPSyIeT3SozWvOxIiTiM4oK0naRHXvmiwT1
VJNLfrH6Nttj1rCpaue1Bi1sD57GleEBNBrgU9ByxOGOQrwaHmgL0ASBI2Ak
7pF/uMjm8dodBTqezX9FulhN3x+2hYsXpW+J/vCkJFZLapmfTB/MFwygoK2r
P+j4+N7wYX89NeqGlQBZiGY+cTQRsXDW7acYzft7/u+Gtge9hcJpbPdRZgBk
OqJBMCBu27yTXpBuJE1DKNzjLbtDWE0c/SKsDN5Uwm8gxxlpRxSfbyEvq5hO
z48qNKTKECRC7cyHalc0wU218MQLjYwR6OHRAIVKikH6dLoeKyOA/jH4HdvC
Hz9ZEz1rkaKd32SLewD8Cx9O4ZQDAtNFbiBxEM1rVwYbDmkj3eTBw65Xsxrn
YxAfxjjZgbMbewvirUc1ETYp/eM/YBKibUCIbqWrAX48lgBHJ/BmjRNNAVLV
izhO+F/Xtmyp3oqhxlP4vYc8GAp9RusMZwmANbVR6T7EC5SnxOurGOZjiDks
kFtiIs831O8gqrellp7Vi2lTLGVY+cSvdfumfRqGspBKv/bQuFS2TnEHvfuD
yYn3QDQ6yQfH3oCQ/Lvpu+omQjXgtjn+8kYxlRTVnjkgl6EVzT5W6z2QlaQg
uKNFFFChOP0fykGaXxWJO59OKiPWQCcfDEWEvzoHA5XH41Iw/DJA2Of5WMzy
ZeGBWu7S27fIQr6tR7+79n5QzyedX7+KlLuHTrXaa/YlLDL5M+iIEakrE3ji
REoNHuh+a8xAXikdZo3ARZlvKK15YPntlMsiCyg054BI7OuuvyiXB2u0UydJ
pFa/U7JlbLIw+0A6j9TpwSI9fTpnC5UbbdYXssT04X4sJNiOuMlqEn28pfRA
hw4Rn2ZXARQaevuGyVGCg3dEVOdKdFXVq25MpHvjwy08V7AfOyAOQPAfBvyB
/fSdasl8prKtqQano/UsTxNWrQ12YCRgxXRX1iSlec5f8PE1qp2EkhsHUGJ5
E8hp8x6XZccydfze8fVpCye9g7K88H/TBUORLxBGwzHcVSK70H+4IkCax/6K
ErhUMFXR4r/EiSujUE+MRAZplq33kMweqM9aJTnwsxfr7bNCIqfPSPpoe8Y6
G98Bhrt1jM3MskZni/eN6TA6CTsMzE4+T4uJf1b7rE6CydiL9HPf1YYRhGPj
+OqXyH6Jwq0t/0vo00d35x9EMupUrn7JXzvyoi5YCpMeObQjCbyeHFYI4LUS
0sO5O3YNn/gWPjjbGtq3vKpvuhcS71igRO8x5lVLb3rgvJ38b7FGO2T4JgQj
EKg5ZZeyBDCkNQgQNFHgdTy5pi5IqlcV6eQRX654/bEVQIfb5w/bGMlKEhmm
+VcJ6gh9duIsmYMaBRZAv9gmgNfS+BuRSyO/G7N8DN0cGfvRLRWdrjpudk7t
8Is+hQfHOeInZa5UMQ1X/dNP1j1BDxstsTvuGjYjbvU50orjUlM414ArabJ6
DBGDYslsfI7Pcc0GQZGvBJjs9iJG9keSZK2TXAB5ng1wNb35vuieb2m0IqgE
3Cljv/G6BDJ1S0TULIgMxO2CEIDYKTeksY089QUW5P0ZBdEmWpQAzI0wdnPZ
GkYslzaQAE08LY9UcSTy4dJ/gDsUVjUQ1pzd/fRz9xITSB9HNaoO0sQ/ndQU
1nk8s7iPuCewJVN3S/+P7QU/NX45VcMoV6BMsrrz+OqETk6XdfqRC2C5rmYR
iesbp/Nx2a3JvyQG4rQJY8rSdYJCuL9uH4oLVvntwf+OTNljsXhBjCjfDM5K
dSydBu+gtzbxvGLrlxnnPdgX03atqaW0i+hguMrhbe6CXz3b9csDgflfOS0P
y1v3pUBlh2ms7bCA7Dzz5Z5DRRImKAx3udCezO/hBbNYeBZVFLuxCYI8gHAI
3gbQxuqixQU9kzuTn6dujRD6Te57UzftyeikrkqT2GkcSS8wWDIk70jjP3dm
QavAh2er0HLOw2rLOwaY1VIeil/eVuoM998BfEBGsYbe4hnyI3MlUSNii+tz
Aer3AUDHEOJ61tUuJb2I9Tfndh9kkTWqMuwnOlru821VgkONg54uqwrWAj6v
eGg7TG941kjghe5nKCfZP/lrw3q2KHFnRBK8yndR/DjaEmmVRJ9c8xTZgcgr
hCABIwilxtPGNmDgxsEuREDbMNcSlkUv2I6GZ0WG9Ai9qkWh+wQNESbOnP7E
XHpKrfmTskGljqzGsYzzTATWOMYKfKv4ClHV5jeRqr2S5JwMD+Xcu2J+Q6Pp
KQ8rX0MEprHjD3r2ca+OK0sDwFH3paKcD7n2zqbAOYl3mNv7QgLnROqvAuDa
5lVsqJxSiM1SZ920//FNhtYH54Zbk36C7UNJwpzCfDdMdvmaPwjK7Inr/Wz8
KZm60uxfs+0yD+GOvwu9JRErAlMzLEY+chEIbRVkDN4bjwF76N/6l/Ax8vKQ
0uGIBuMl49puJz4p4JVJa4Tdbv0DLQIt5C+uDQO8MLnoRr0FdGpjdVOcojCt
rb3Fw7j41lyeN6K2qK7ww6loirXpvmh/LVKu70Tz9SAK+H5eeirR25zLFrQs
leCDSHXaMY82i5LdSaIRurP7VSxRrwuErn0bigZITys3jTPghHqqY6+9c6KH
GuCZv/IBLLzcd0af05BWS58/gHYq5ovBeS8YyRY3HXnZ8Mttd9kLf5wUb4Oz
70fnSQ+rXukcp+kbczaXgMtYR+WEMUH0LXyU1Iujy+BtasJpLNJ93YBJi5DS
az3n1C4SXcXNJ9d9U4NWlATB3RJqwtw8SwYClNpuWdTdTeDz8GDc9k11UfHw
ZXpQrKqTDC43Dcbf4a4DxHskrAnhBCupMkZmiwM3ROVdhsFuug05XtpVUcay
U51ZcwtzAd6z4OqvFloYXbtMUvD8nd7uUair/pxhMOLrYYcl+fkI57rPD7h0
zHvn/SVP0uaGHMp4h24qLimyeR100+mbi0Dxg+qhXK64qqTT950qoJS1JWNF
wYouhq1lba4/6p3Lx5yRIX2yuOlBvY9F5HrU9aa9IqXOFBjWCF45n/C+bBDC
vxuY46QnkMLtPAts+4dQ25RILrfit77JStpHu5I1lIsHnjwUVmZXpANWGGBn
rBFIZqJo53Im9il8Dhnxk7C8Itm1AdKvAtPACjacw5kvfo07BEkhQo+U+f4o
4SP1hxKGsCnXBDBuixYdkutJbVohM5RCPc2jH+Gb5o0nmv8qiCxGLrmoYvq+
zBUv6oNnD3oBS8/zWJ3SGTgfogIxccuUK+Of02fggchA49HSL8fww/Ly4DvA
q5i8tKzHsenmemconfbDbrHmpIS2e96EDiwvc1BYIt1N+857Mq7L2hKnUa+3
57sHUpEHHlaxDBbR1xHfH9TkbWotvYJZpClizweiFfN4MYzMLZwFQ0GRWa69
cAb9ZW7hG1myVvMEk8WYjBa5RnqZx5lLUEidGs+nSLiB2yUjYvcWGQtCPBA+
cGKUfkXnfWg8s9ZBZRZrajGbM2z7wZs/TaUGrSknto2k6THg4gpZbO9vkPK8
xd15CHs0EgtJGzPT4naBhN8LwmoZhnDtupegbk/U3u2CNDZbTDOGdkMrSNDE
RHXPcooR0ORhugEALkoNgQoD+kVkVw65LXOgpjZBO82CTVCCcOrTc58t9uGu
rkkT+q2frLTvp3ub3Ya5T5UkdHAYEEKMrnLPUkaU0RJDCJBOo8OgDVW/LD9P
YafjfsaG5nQW8cMMgKDhFcVoVICzFT0jQjgXUjpJ0j2uSQx2UaEZ4ksBEz2V
T1dhX5F7ERMr2bnGm0dJLtXE+tpB8O4jGUdVvMnpDTweXCt0KF/hCCdJyWqq
wfjXF0v2FdcQGRaA2L2tPcTFAoIPwiVBeccqR4iPyEMFJqoSVZAq99hnCeTs
ZIfJM3n3IkO0LnHkw7AqY1tKkl/GG4v2nrKUGeEr71WUP1hDYm/WnRSQlx5I
VjJcdBWmGyL7R3q/sP0wgAyOST3d9eWsl7SOMiReeKkC5K6XO+qFOOnwskl5
IvCnDo8tJ0zvuYuqnEiUKCej2ruIpOi62i4gKC9WqGyxHsKvfYeyLdjmIhpo
N0kHkT+ZzjZ4tGHrLdeIkBrptTQCqhJca7g4ZVyboZVdAbxkAee3faWpIJNW
lf55xuLfvQlG8NJ1Eo5a5r/vXXLrqwHJQKrEc7fbHh0xs639WsB5QKTqMkLk
swRQPO6eKjHyxIAsteXa3EHHvLCimS38HrHmlAgT9QnpnNMTEdAuknSKEI1z
u06Avr7f/XSyHSyNXtjc7NMoPRq451/7wHQQaURrpJ5Zk167zT/VjFQhFtyo
uKmW6AEBfN3WcXrLT1zOo5HJUVb6CoAbjZPLFRpSBUSpbFql+sqgLyWQB5lL
LSZvKjHuhLsszGLWrGohWfWOaiPUg829thAa0XCj3PgmDr2cbf0Hf1/qBphE
Vk9DmMeiZRt18Pg0c9pGxVg8uLYMUGKrbdCUUGpsB4eJT1k/by4vg2cGcYUr
BpSBX5x0/sbpS9V9F1T1Y2CWoGzo3calDDYaVY1+FDW85yChcCG1nlI5VBj7
Ky6VRnfi1Az49lJyQe8oBNEzsXhO9AmT84UfF1E6MCrokpmMqVDo7jvHTp+4
mXVax/+1ZfRGVMH7Ux3QczCYEWREFTlDax733LzZ+9JlcuaeSWXPwfgexF5E
LICeoO+R3pRuR3HaT9b8sjah/CLHVgRWe59ExlvWwnrS8UaCfs43eiDfVrvJ
kGUYbIeKFG5/wBYsknVmH+CEwOYKNOyk7SSObtHWxIPzfWeA2NG8HbxNaScv
muEIKKQokBO2BaefeBV4mr1U8zijk2FtfUxf3L4GeiP3SVj+wRq1usTuNOMZ
M9amit+nv//CjzBPLRLt/QEudRffhrO3unLxuWedZnw+1kY1CXuNgzuPmSRp
wa/gfVFJX18d3fUD0p+3hUNvGP03NFiHYG6DWKtnLY9mdyxVAnF//PABiXqq
6EdApNFuRUvbWI3voICCzuK3Yfw2xc000bs/eXPGvkxPgchZ6oTJciUymOII
CrIrEaOnJ22ew9TUKfcSWEgLggjTmEE43Gw/H3sz4QbRRj4ckqE152NPbh5P
ayFdIH5Nj8BTdO73yZCyq3R3LBfVdUp8r44qnWvw5oK1ZocKu7FM3L2pTOjg
SDn9PkC6NgxgAuD/z5YdmX56Fl4nnYKVMRn3ef8jTvcq6DmFVBIZY1b8R2Ln
Hh2LL3MOyvK8/gXjz7adtIGyf85y2pq2l4yVDJCD6kTBiUcAXPLqTnNmja5z
PDiG6zx48tAvOOOXi3Q9Kj+ENWxXzGuMbd91yM1SvsCRxouYGklHjbEIlm0+
1IZ68T2MdFP6eRUcEY+j1Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpejz8KgZlkDttimm2xt3TiKdaJoVz9+euJRo/RlsnOpDSxwy1p9TkoortvCK8kR7IPF+IKW4/poYmj37zx14cD6rYsMSWrSHu/zNBAelXPpFe8/en28f6m1PSh2I9KV3z9qKXCJtKRmnm0wglGk9Ny5JKznNhMJDV7RegcOdJm3GnGkOMyDjQOGv9mJk5KWPxGEuQvnUSJHUMEUDTswwssziPSxUDt9yTquzqje6sPbr8HS4NEcdCz07tZHMFHeh87sFY+wltSESLjcUlhCOYoeMJQhpyv5G1pNMmCxZfyNlcOtqpW3wo/r8uDS8Hup5R0xKq4tUbeq75BpWM1sQVHHNqlj5h1bXV++41MmlYsVNsVYsIPAwu5zFls8UpziUI6PzJObKRq6zUHCjPGJZbmtXVFa42kX/fbzeJn8WlnKDr7GT+PJnmBVte9a2gAnU3Fbn/VieiCBdSWDB3IQIpVs3c9qljWuTvYPjvHahbrCbt6aj50b+d58H3Rtg1kmrg5y7WMeMYkkKuJMzlF4WYyjlSIPDlc+Hbc40Bavcsm8LGv8qz0qaC8Y2OlrCHiapf25a6LrgnNkQIatn0JUUnD3OaN5XcXWNI1FOfoCObM3QtwmZZDpgLEMOVFOgGdxSYdW0Tp4ClevTfUQc12ALjBGY9Im6Uq19O92zSH1384o9F8k4+dtrzp+yECqy/mnAh+g3E/g/+qkRfMtvZWt+v+liTl/JhpiJ/57g/8AlVGCQuV8GBW8vOIKGrioHLgZiIlVxJpe4zmAFHsDhAt+gEsHf"
`endif