// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J5H1YN72JzCgnmCwUHHYxFopAjdmYevtoYFyRN2Igl8Ug8H7N2NwZnPFUqxk
psSiBlCeEYVewztz3pchejXLNr6YEMmh205XToRYUS51f/e0q6MRautZLRxu
rTsXMPZfhnZ1MHbFDGsgtkBVQY3+4Rv+qm3lr9O5aAwgFveVvpcIOca+pn9q
Uptb8wK73+o/QZvEGRA/t48hX8rOaT4E7dncCv9TiDD4EHidU4Ok8uOI8WRG
LKcGV3FAqwLEx/a1+WBJ2E/KxAP1d9Xf2c28XiiUl4ck5fqPfOp2gw608B1T
wcss95chNgDGB4JTTMgfv3rcKnffLZGZag9IjsY9jw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
myLnYyiWeKZvnFeWIAoeg5F8+Q0L8QZpWk+zm8jgoCFalSBKVDn4QfUEqGl7
C2y9Vnet5QgPwBDrlYnrWDkBblnq3VXPVfe8nGsetFVBpDp4O/eNonOLAbUC
oGIKoTyermmTwCusD5RU1mZ58cYVXgo7i3jXjj2Y/NRmgxpaAqcufD+N1t02
yt5LIs3NRO0omorokmdAk4WnZgeETKkg3AhPbTivUxayYYPnwdXZYg8H+vxt
nbWAJ5I5+fD7PjMm7FJDQudPYpUJim97HHiGew3Cyeauw7V4rVE8AtEe0UXu
Gkp2VrOp2pqO/6OFAvAvaQR/Mdy/8Nr0mTCbsLBCsQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h/U/p3tJsp07brDpdfZqY3h4VR+XdoTQPUkWcS6xO/gx0p/3pQq6NpBaLUAm
uX/C2qe3M4p3r6W6EXt7cKBpDKV3xfcc6DamUs/qvrG3z2BPfXYl57ynqw/5
YzyUuce3pRl57p7VDtLkkLBHr6/YgL7u1rmtARCgANsR+FnJyZftI9sbY3nw
8XeCghaTfV0i3YMuA+GV8RbJMFMVV4Vlc8J2Qu+4SC1Zwk5IuP4qC22q/gyj
vbpRI1nLM80IWghiuYuQMny99FYaBwKxuT6MLa9ShjgaEujWwxRI8Frf+TKX
gCvpkgQXbgOV39cKLsVZCtDuN8WJMabb0H7b8UHlmg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jkYbWwOaOBKVLNnZ2U3lwxR44MVvpkCGP26DwwraC+OywkJBZJxBVUlY/i66
oAV6ZLLkyYjGte2aXIU9jkTCqlx1k+ewz6taQMfhE8uO+ydMxtRYaYZrbBT6
w6eRHAy+WhhCTMD/B47X4lMxWLVC9g00yTGb4fxKUJPETnjhA4dVPYDG7gb1
LwjOi4J3wYruQmPYUS2DWHbXudSiI47PT+kpRH4g110ZMnU6Mo61Xu782+P0
9qFobeo/+dY4mINFNL+nvDGewT1mqpYQvcGg5yLrCavfTfjfbM97IbYtpklp
Ge5qRMXnVH6rkjXF/7mYeYf5rkAuXXsuHl38AKc8nQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
atluIiNcGUQQgwFlw0Ho/4OuLwLsAKCFshVODUJsTI5KzTpulGWHhejK4NCZ
OJ7FoFIRNoXxFEdVcjCJWwwKPpRNXyLvjYhA8TQqAeamRkkTbQr5t56B/r/o
PG+bZ4AhQljGakW+/RZekez0Hxl1I3m/6vRmy+nrZHEKJYItbWw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NCUvManj/Yt/3Rv72dfS6nsc91m97eUItZUVvn0x8cxOgBRMjQTgAa2P139i
xRsMiGk6lMAOzGzcz4DGpd12sf1LeeZf1dBRJYCUW6EW1NQZjz3jCMIwccB7
WjWdf19/6ChzGHMhhrjTcDdVuE3KR2Z6EHi/0rG1/F3dI4f7pd3V0vrymvLU
qW9Xkyd/F6XJy6rkKYKG2sVt/OAyiJamMkNLuyexifBdfcAreR4VMTV3/6JA
F4PG2H5ROEwXPxXzbHR03LmLqxikrWr2CHIKC+lU2Br5GUwzW3VGR5yc6hAu
FfLQZcixTOzeV4cOj43UqVII1CxRbjnFLZUxxzlb/XTsDa/UE59/5FbZmgcz
qasSDkkI9SVM58utBtt10p24p/AppfLmU878aas08DmugQnBDPWRPBGfod9k
LZJrqanf59CqJPyPIPMNT1wPHRLd1+WTqOQJKcEY8+LJM5rKVR7qwCba1JMp
W72WL2WyyptohNyn1iOxw4pijEe2/Nk1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YNGEE1lFPGAFtCogzllcKU6gt1LK2F7q7OLhSgrj4Ht7UPAkiQHuLPr5WsSt
hmRWWix2o3HiiCG9pYzUQpnD1ImKqUGkECmC2HQ2DIYQprLzhmx4DgWa657k
OwgE9GussEkjD+FfJQn/xdoLa8rzaf7XtyJ3zVXZn+edxaACNPo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eu3+XAHJKZ9aWPFtVFRy36KlSTyQHW7xX7dpMyZGJDTavVQO6swsEnp+KLzm
04gepfdole4t4ugivCwW5RDF0IWCaLbpdmMXk1D5Hb58112//sT7+Yb1V1n/
hjp36a0UeFoJG4JdL2xriIgVyUQPuHNhxWVYrf3sMmjFU7Ykowc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12976)
`pragma protect data_block
ptLXFGJtPD2YGGcMxDiVGviPUlQc9xL2zlUqfu3J4qD17GiE3Wstg1reww48
hrj5zxB3J8Ts5JnuNGOTfVzDvoRzRovHJQGC7Rq6z1wjRGNePi1YDKQ6RY3B
wBYvgFQIwwslgYe3E1TLkmtjFjtKij8s5bBjPAwR15iMqZHosD3WVJMcCink
PfEyoYSgAuVHjX8ub7Qn0t6brPEMWL78zpXVZNSZe1MkhgKWF+ocUcTa74uu
jSb1lAZD2anxLbkR89cyUcJ7gbRvfG3JcdNe+gG10bCAg2PetLxROXvBt0h2
01/4Iwc35pLLICnzS5Rl4KW827+dSkIkwkj37vqOk7aKm9Ll3z62xFL7M45d
6QLCSBxB2AK41OALypIB3xHKWZsPyU3VRuC5bmTtAW0v55pvYgboZT/evGdN
OvR9dI2/3+gOXtF230Ea0mqBhMEfrGq4+Off3mJv1do286hW8ztxEfvQHU24
UZ2/n4lRELbrORIfDeM7bSD/UBOIQYqa02pUgswghUBs6cRHkI5+ae11RkBl
fVsEPawEmH/KYtk8wfMP54xu/nfjLCZ0NST6IVzTv8eL6zzEpzBqMUQY76+P
IFBwJ7kt9Wn0eRLKudWtlNHOTl6GR9UBoKZrrdQ3TyL2nQwjNRMU02I961Fs
UJ8jMM901ohoIdZrfXER+tiSOqk5yfJeF3gt3lH2qMAIippuwVub+TRBLYim
GPWjMk3iJPb5UmIzP7f8fUdGdaaHO6da/KLnmV3IKsOjfwY58/M08TtJHck6
Zh5S9Wq+3nY0s0fEZm8A4dVGukAjSGlRBiUPvp0Xn652tCxdHs37wweyEaMC
n68mldpA/wh39nimNlKqDnJWZ0uoJ2JW50uwQ8/kORDV3Iyasfjpvk9lk3Se
80XwJ4k5+0SO/tZwS4VXl5N2p6bZwKqRZHdM0t1TgSgaIDzc9yPbzP776wu3
Ni0rxQuhwuopyLonOORujLCK8rNJSBMIIueLv2IxydO84faMO95ibsxegaQa
R5B+K4NXj5mf74bVLI7/2hpU6HDtksOpbqp8Qha9VIbvi2QcgELrMORyms08
2CO6OZQOpEQ2k7Wv+l8dj5zc5cLZHtAVlQ+tLs8qKmpYOYdFXHRA7tRPB+rN
oW27BEzUKSc3QcNpYceYT5/+oz93PGuiu5fcMthzTgYVpvIuaSlfDvQz0tWA
R1b3OuFf8e7/Hcx3RZrn4QRQdmutYJOklqexK2VuoSV5o0veh8md7Dji8mtF
zhe8CHmU0WOg0lV8/hTuH3SbcoCW5xYElQzSDwcl/OFZmYyuV5W2zrnHuDqE
0N8RlT1MeHx6tzQ25dIHUBGYGiaHdjsbT8saq2jIjryqxXfyfcftqNnVSXM+
RYjQJh8z3ubZiCfUHqzl9do03bKv1FQiHWgOT+hxCA6bzp4VG7CAO7/+wMi9
83Ku3fuCE6T9o6XWZvlkbVmhsbChVL3lmwKnr6xReb7c+BX2/T1IuvbXXzFE
onhZFJubusTi1rhgkNJ8kip/zri6XDguKUV49pCePb6maSXvP7S3lSq7Uasc
ur0JX3T892ChgZ9b9nuaEqGYg0rBVDvl4LJSwEoU+8e7YS+i76riGVVaGn0A
29TP8Lpw1SLZi+oLRrHSEiLhfa0CTXBw3lDw0GFwyktUZW+gKA9kt9mdqUrb
NKZQ0fFuBJgECHqxo29SUhsERyK6ODuJZKpczzBR3jGe9Jz4fmQyRXTDccf/
lny82wBG0ajQoaU0PfCpcPNHJDZ8fOY54lT/HfKMBQi8Qmr5tXJgCFmHNcBB
ha4eXvNsLpt6nzAbgjeWr+yS1nNopUV5jHfNZyB0WZdbRbXQbF1qCxbLagXv
3OZISo7buc7Q+pZYTtPVvcigT1qP/+zc91cvqmbj229Mv1RFFVmyDgFiYF4i
lowuIAAs0V0oRdwH8dg+AYgYwHTknKB4s81NFoMN5ALxMC32vqk9BL2qtDEl
8lDT/qBUU5tRubHuoLgGUk0b+C/SHZYnWY+zR/9G+MIXQ+TAGt98RxRma/AE
OTHxqDSo2ENlQVNQsVqLjurvaz1kiHbm5GJn2nbw7Jum0ReHX88kh4cFy2o2
p9SPmA/Qbpa5RWJ8u6KEBy4ReUwrscRF6RWaJ1D2cz5N47V89zDSC1YzC/lk
xFkb8dOsMmiHUlxYOVbTYu3Dcfz1y2tHDz9M4qBm+n6w6DHHqWHmiAnJnEMd
hgEft6PVKgWttxmgFTx/gIrpuVdvlw9GCiC4YgmUdUqvZ/NJHv6p+LXqTt2T
LoAjzlEpXKWSHIcLWRNnPfFecOOFLmooDHf04EX++ubMmJMc7rz9ggjDduKZ
XG+Pye0+TFDMkEz3OkWQ0eXAfQfyI/HGB8DEMS2WeZPcE47MEXIwQgC5HNEz
+DQ3ZK915iejzee/wLm9P2cUdBKorM8XaFl1np95fkY5tCHt4vGQbDSw2hxi
01YB8cGuMB8vbxpZq0VffJ5M+1sNDPUh+228X01SO0BQc/LgOdBEyd1LPRdK
Z7yybArRK7T5qUOdLi+c2czMNeBkuVLAo5U2wLPAcyoq61Nzc/r1vt+lirw5
jPrhGpF6TLW/lkRXuEUgkl3MFgzc2K4Hee/leDOsQEdi4xiWECqSBnSX4DrY
lD5J+/XhCmDRhCWJvU2JDgG9NPL93oniKWaDIEqFeswSwchJvf/Sg9M3G1ca
pizK680jrVnaZr8r6ygFgDjrUhJRI89D6yKQAbMGnjgOd9puc73DVESrReOK
K7XOH9JG+JAh61cIBG2ilHdEqBvrTnbapEOAAwZFurHxZ4gdM/elFh3ZQjFR
5DPSjOpjRNKvoCBFPTKRmwuQEN+1J2EGt2HQ+5E207vyzf/7N3KmROi5Jb+2
jnWHq0VZrvyIMLMenGNRWc7cts0q5n4+8ALt5ubtHRd9BP+m95N4GiyyvzKM
pHvEQP7mWQqTModGbsjDawS9OFRfXhwvnGi/0cYyspWFnxGY/qqKJ3ZYM9bB
9BBoZU42tNbsHUopj7aFzhk0oeaFTZ1aLbZ83KsmvwFoUQKTFnqBj4w4tzuM
4suULo8ZosAP83GGqbTH34XI7TL+rJVVLt6yRd/+gKGXVeWGu/E/3MZm2BlY
PMXsp7kwMwy+usirnFZuLxO5U4IpYzB1hr3+K7Vs7v6Bf9oWuQ3leXkhph+/
Jom7otVxq/ydEFwtOg4Yw0J/sGJuSHzuiJ2C6VENLxBM9OBcheVkSp1Kp5sJ
m5nUnXq7pwFIuI0z0U+bPykC5rKJODxvFcC8W7yB+hWC8BgxRAH+E5mOFnGg
uGWlUhURjsEX3IAZg3GNuD48Lo192gGjCnuGfcwJi+Op8mOIkkdPk+GYm4pT
8HRijk1fnPNSNAoMq3XmXDVIdvGtL+DOixc+5HByVRprWt6IlRzNhtt+LPn4
SSjGaSw1lu8PsFXMWk73TbEH+/C3lbDfHZyVSWKpjObm0u9YcTjyVHXyrpgb
7pW3LsyAZIdQdPVDHUvlIyjXxKRCpeMccN0w+Nodbx3K+6ud/FCddepkgpE2
lJRadDutmx6OvjxC++lKPXGNNuUQ9kAIvQvwnz8peprp6+I5yWzXXun5MOUs
rqSrQv4TFGuoSTCqJdy/xJvw2++tp+fpnEjVlPei34EhtfmvDRxjhx6lAEnJ
Ah2K2v8FtThpE5QV672/60cEew1utAr+YW7eRkgDZYXInxrWteXQcip2I0a9
yUj/Xvxt21OXhaPr1tTzztnjULQBWciQKLNj8Y6RGPrvNKBDx64sX7WpQFo1
hcTzPXfs8W7SvfjVlttIb//gJ4OUcF3BNuZ53klHcR64vkyAZ8339D0lC3V4
fa+a5SGCAiL0pnyXfXTWSATQXuxkMb7L5hff1zPSOXNjMSQVjuyYRr19+Hct
CxgJnCpTgRJxs5FPf8oWe13RyIKlTZwpXphIhn0FImWPRyWlRs/8A+SHxJDo
pO/9mKU0HczIvV3i45nDsZYmpUn33WZamtJCdENTuGLYGPTDSbird4cazWeW
A2VmDtnOtBDmHZgcJzN2LFnEmH/ZTRW3E5ofhJh4n2wnmZzDWMGLBzDa4t7y
VrBjO8F9HuH8IiAbtYUJ10YL5su/yyNwfOFVclTcvoIk8IQoJQoY17HN/hrj
uuuS0tYFrDLBDE/3ZL3i4AVSYxdl32lVC1NuoM9M6gDk0KIKB111vl9AAbso
VleiZbHdkmc6Za/ka2SdFsd9D1YxQc3/BlzTDED/c8FzCcVvVF2nl60t5ixU
FrxM9dQXtN8903isKsCkvVFrRIa5IxMuF8dFMY4eijCYM8d/eKUetaAacj5J
RySCeKkpW3X51JpspG2F4o4onmniepyYOgvChYmdXexQlfUIk2Fh4RBEnZN4
K6F6fEoquRcM2GrigFnaSJJ5zdlt3TBCZER9KMye8PHPcJdB6yh8fyMqwShV
VMRDhn/gjaJuwMVIYRQ4yz4Y1egPxzj1YW2CdJxGTtWUjzocIXOO2hQ7byzV
in/OC+O7YeLdOLUGgK1Q5mMJCpnd0cibs/YeUeI9ct2PIe7QC05TTFBlpRaD
4hkvFBmueUZcW5BtPUksxkMlHiwEA/w0i2ReocKmfLvcEpDcE+1GldVeeFmX
FQvSVqu77xXkwpefzof+/3GRsWQcpz0hh6YDQQD9RSG4zyiT+aWv81xUbiGb
Zz3MF+lU866FRoNyAoR+FRr/kc+iXm7Xlo8Z5vtB1dB6GGAKnBvaCZOuiUH1
qFaAIvF0TcGDfUJ22UTxlm8SSIKrACdgzRb66lO5e9GFLWvpXwB28eDyf72d
So5FS8jOySLnL+V3+vXNHojt1YUDRe5oesEcar+u6tI7KniUnyfpN3S+4Llh
Yy2nZI5dNO5LfjeDWZsTtdzdZmRR+ykETsHS9zkd9/qWBaf5mHWnvAfS3DaN
v6/KtKX77cTb6JEs+gRHbmdyEigikPXYxyQLZyK+j8e2NW0FNOEvSOKXn0sh
eKnAeenAeSmPSJ7V6b72A5o2vKIe/dO4sc2OnzsC1hvIMam0kXqrsYLRSisb
qrCpkuor6fdbJ/0901udxEN09CMRijMipCyT0qxNsvJjqiTbyKlpdxdI4mFb
jVKHot3OGQl2QjRKinp9GRjEKgRSXmCurTjRePEWmLz1k5+ZBzm6spaNgFt7
c41CeZfWut6M04kyK1rtYcs8FoltTBCnTamLAfK296TEB+DkubbSKRcFbhjn
3S0A9cB7YJXMrpL3O/XJNSo/gRMVAZeuDMRyhORPdVDPlEUc+CgcIAuiMXCW
mWN//AqLXPZwiMFfUfeYgQ9kGlK0aSfcCG7iLMSoNl6Ib0k2fciZkzMMQnYq
xpMhoZ9/mG5T9twkPJa9pQoDRMX2UySGkxVXAmR4KbBPv4DcaPzQdE5Zs6su
vbjn4EBNogLNQFzi2ZqXAA/p3QKKz6Ts7yBax6I8lhP2oQ3++oSCABDPcguf
c2DNBMclJ49Yzwy13BoF393kIX7/g/MH/2mT/+rc1kMHQNt7LEL+YKJ+JGXQ
nord9MH81db2ehzgWvMGoykpsJ0hhQwxGpM3sCdxp1s6D/ik7BVUVCZwlhZI
VXHBXIwUSlHZZcQJZxzSwbBXXrhAMeCevvQAlu98bxT+aJhjVHzVnSYXhVil
+aezGOj+YiLDOsXr1W4yX2fBcU5oHB5Xy8XJM+ADeFqvb7PYn2sGscMFnyBF
1eRevp17weUk3Ec2gtxjXWg5I74FJd8CIBiJX42t6Y8yaWoOJjuMJXzAX0FV
u6HARw5vuwHyEFZZIBo5Xr6K3lSRButMo3r5kQHL2IOG5zCCqZc1+U5lLO1e
qmpoE/Nw4HjjCcej82WIvialzR2TcZF4GWJEYlk/wcSSjA3jmmxR5d6V8G3a
v6pQs5as+VSPgkPzTzmoI7E2I+UNkwz67YPgTpueSC9W3Lf4gDIcFy6T89q1
/vkFLGJc4js5J8PG3vKTOh3nm6Dso+RMxf+rwqMqIE0r9gW9M1wAMg6bH7oU
Wvcv6x11cPC3AzLB5iSLoNOsLFcSyPFFiI3YmsoByB8AJP4gMcT8h/2T/hCo
evewYNIDIF1UI0HIprtmcOOXVKBO5I2HKY3wHYG70iA/+38noWwCRznz1zZh
K/huKNZTF2+LMRJFST0zcH4zJFPfKvuglT5ANYwITICpt1Jp0NhmuNRvsPet
qIGmmQg/1V6w7MBgQzQ51Vqw9XF4rWYti+6VQWuNh3fdw/ukLfAMRufkIQwe
39H6V7a9rVPF05AIXSEZvW3uOU87bPnMwjbU8gwmLMuEerm+hTzkSpuMWhsp
qjbeNFrbHVrzTsbeh+p44+4EctQvJQ5ee3YjPaQJmrGl+h3X7SclUNkVF6QP
P1U0K7PGzrh39pjyHOPgPO6cSP63d9LQ0bi8w8DloXaW0nAn+wbelWyCryK0
Z6P9Y73tYRLL+ngQRSd8HRcM2LnsOt9YEhKtXsMQi3oQC85Iq338Yf4YWSvQ
CoZhILNy4+zOoexJJQCxaMq6Gp2ip5zgtHDXx1TFx5MLpK7XI6p68bXgQUpz
Y5J/LvrpgUF2P6E5ncKdY6mSL+Atyvh5JI1WX+MUa/BvNbentYCG6KPBGSyb
KIWj+SZStLQMMvSoNIgwNWSLoc99Yw7YlqWwj4zaXDdSK9vjzG0AAwLTStYb
xzVgu456/TDl2mP2C8GieC3BEsWkymcJ8extgCX0SA8TFREsiELv3uckIedl
9yzAusEXMzoJhmuLCK27jW7Qlh+L0pVaDHrx8SSabvn5sWcUjSoqriWd9FQ2
5agLoNA4+1nQoiNK9lqkxsHR19Fg4ZBFt6Ew3eHlddse8Gr0UqIGMp1/mHWU
tzTgZ2MYTSPgUdpCO4gBiEH7PrAmzRyEP+HzBGHXWBKGzAOXN9FCbdGh4UyU
qIxaezIjtqNDZro+0HSJzH/6utwPextO7US5RzucUEdO+YMtTFLbvGyT1pqK
CahvUmtwkGkiLVqqM9BDWx4cYEFBGhkheCsWjBh1PVVTFfna+iOZqRWRsM9X
LZHiwT2PX8LDb0g1ofMOl0I6A0P8CtxPyNKSZmgpdCcz1FsxMK+uflx2huoo
scfC4JWSIh/xikcJAQJ7C2bxvVkHRopqymbdOWyabvhAAcuNmzlp4kkIvKim
RP/Iy0kPggkzHLW1Si6IsrBgJXw1wpjEH9ea/7R22MhCc5qUTsUQXBEmJBm5
4GxQ6Hjsq68hwb4aT2cNyBStIghp3gnGeQVrYN3BP3W+O5Us5AkgkB24admE
ssvqSZMR6SbGNkTTwln9LFS2OD5qhVMwrrG+Qenrhaaizoweu71IX4mW0d9A
WXQ4FI0wp2GE1u0vltotTNAkMtmDPTxwhm3p/VMJ8TYAq/zrlbs5sR6oRK1K
rvITeJSU2mf8SordnkHRmANu514wJsi8h4/O63cSiU9eEN3FU+MJiG8CWeKf
ugh2qNmv8emX1tB8smZPk8qQd7qzoEFb1rI6ExBX0OnDRfDk8o2cBnZ1kdw/
19cjvnktD4gIT9Lzv8D5WXQAQLoK7F/DHZJE8eBFVGWGLHSiDH3I1BvE/+/M
mS3esWTx/8yhHbqkzWVLtITpf+/198NqDMa8WhAnusqXcse5LNoQPxdRq7uJ
fM7QnPadcPq+KLIBm2Cfx6nWM0yfdwjqPJ9F8G5TrtzvM9BMSP2aqAiuiZO4
rk9LIPO+t9xXNfUmTv5zkCd/ck7YmSl73bwHheKyMlfttX+g606QNNW4HoSZ
ZqcOpan2BzvJWjHrYYpKH1+6w9BcM+LctCXNvkqhE4pM6EzWoRpIvtlDLYZQ
M/7m1PAocZcw2XhLrQuvIZuX455f22d9TEfBxAxpsUxsM0qtUtR5+B2CJrq+
YWfJG/xgfea3dvqjB6E5Z6wVpY+p0jhtCoh2hcsU9YFrmarlnjYBy6ndyxHR
IrbmlY6jDeThEb1Zl9i9fUsq7x8llGFz48sdGLSL9+CdeqQolnMvfmFG66VT
XHQnjMX80MoFf160BXr7v5fORLLN8gFwETE0zLk4lbISBv7v97rCCcQ4OTXW
6G1XxR0Z/0xWoFjVG6/48nwBZUFh1vgR9/js7DP3Zk1xz9klQEGhJdflneRD
SMguSAczgjTyPCxAO2j8PfmXAPsJWpc2fWRvymYxsvS9a6zs8W5DhvkF0pME
TLkxrVaBHDaAFp8WZF6MGBm6ipyUvOLJ6itWnF7/1sVwy0tuwfzYzwRgwqiw
Px87k+DlAGBEEfDe4hpz7Q6tpcVdWoXuxp5iDZS9jQD/jMXWcKBImJH5kEGU
r5C52wuQZFCvq1B2TlvsrJiJe37z7KCV0EuprZ9aGynmMKalV35dA7s/+uTz
vJmcCsRwDqG1lZDWT6FPAcnXUcVbW39k/TPM0Bpn/GMHiOsDF7B8wardSk3+
n+3unousgiuav3inE2M2qRaC21UtQd3ZbtLuli/euEuNWi8gt5c97kFcduWY
Qb5TOo5c2jxF8cbF6epXI64kLDfG0qFGwIRMEyVjBIvv6948y/gRCY4mqJd0
ADAzhkBo54Ao0RirZF0N7KE6N4WsIQviraad5eioimMoLs42jmihujBkWPFP
/X1iv5wQdLhazJJoW7ocUn9M1GwZLTp/Qp8PzxQDbvD1DKVwVlfwMPfBd9v/
ELdNTB1FHeXjSTO5tSIc2AfZZK8XOkygR9RBz9g6C8ZBZ1A+Z6mmiHFaJKZc
O9UxoIKDUl1QAqGWmC55y6cVDJ1YQl/hiFiKGQ47Ojiz8NsnwgjCWF6z9qPj
kqF0SU0En921LvbcaXHP91wsENy0y/wNgF/2ra5NTxSp7H0zkYt30HdwNmIr
qb6ugdXkSHHD0xiYnh2FON8JAiQuhJ7KcDGae+ffKARoFgtFg7Tub8BNSmYW
VnGjIgYlDb5Anv+xLnfR3KmHJI6shIueOxHwWqOu5rpkbARdBm7iSfX9UnBZ
JDjNS2lro/OkwNdIWThiMyREbKYPEFvFHEBs/nCqhRgGMxJw2GIeYMIkQT4e
iAz0NI/uIAeyZnYGVkghXqPVZIc4gTA1scV4D4mvNWdnuvAQhmmnNArjnP99
EbKUG9ymsRb/vdpiwAtA+Zmp45zJRYy6OWJm+FIQIn6m6nNgvmSFI/hHyM24
ll6N3sYYGCH+qSOa7CeNvQUdFPs1dojWqwjwVEpy2n7V2LGaJOTQG/nyagdn
E02E+OlxsPcO44o8bycEITHEtAYZRno+giHXBgh6cs9xYDszcnTCgpgQrD0T
JS4jT7g4+QNzu/39e+L3UUfip7e6hqfJfd93wyKB00ylJTsIafAI2JSCrSFY
H5Fjy/xuY66hkSGA/Zoto5v+5VfMdaDcLJP5lisadE/lowl3f2DDILiBlAUc
bEQSffPd00idMlrhW2dUAQTbP9j1k5d0vU8wU+HPtzqsJ1izXtXq0MtHBVbw
HIxmdfGzso1ypwK0F7cSI1ixcUfx6yGWJzgcYNoG098aCaJ8i5tRyaFPCSZK
N0e9aE1t75c3DncYfY5bgONMmweU0UZOjFYVGSrb9ZFsl0W9KxXOVf3r2LVm
D14tZ26NOkRavClYYjkC3cS/f6xRKYnnzU5PYnaJVC/g/bF78V/tXo110JJx
1wFmHXjSx1biCReN21hfubrVTKtHMQ/lDT9v3J7V81C2YqO/bSASAdaHA6ph
VSjnpRHjTmCzClA8Zi/0nWFWVWmMtC2qNjd/bpwaOvJUe5JPeHmzNg8uL4uO
Gphkeao1AiyMP7GE3Lxt0YtTGp6C4eWoyAvsSKTOgMreSi7Qrhfsto22fK1f
6FcaVLdx3WfQDeoKdGlU3tWru+R+FJAd1tKGltIzHdOnYzei7k6NTAP28Ke4
+iJ6BqrVvl5YWfeRMoGnjb5aPsrvMNleB4scIflmSRGhq9+svCC+ioQAKuyS
AnCLxaFjQUXSkOSm9yS5WAIWuxfUk2fFM9l80SEUywCLuFZt3iOwStYLNTG1
lfEZMccnIoU4RlS6jE5XLeO86NYfgmHhf4jVlJY1FqNY/sHYwR+/x/6FcTKf
3hgaWtOmh3unME8dJC/EG1UseQImLCIrpHIzWGqvQGJrPDWyic6al3lo+ePM
LMoxgVa17QyRx9wuKQeMecBzzR4JJEI4txfBo2XEZHyyhjSV3kHKYwXD+XCl
dwI/Jv6gI7RuIxpNjvkkW11xKHPZX9y8gQMAR05DimqxjxKyHhhZY13bPqr7
pIJGd8lAzsmo96eM7Ax+p1kpqbozpAxxDOujZWkItfi3dfHvtzNHUco198Gt
D4dbHBDXUkuhxFPDTDbbnZ//bCJNkeStiaBudGnMcGi+CNQ5pLM6uQyFK1Kb
KGbETT9I7dIbrZpYmncZZsyqtykVfFiBRfhfWOmfKg2T/B2epFg8NR5A+U3J
TPfDbzeGhOs28uKXdpLPNVJ3SjNVM14LMvpI9J+Ah0PIw6FsgYwjfpFfY7Bv
m0dpKCbFqMebTQoxgbsfOSaqOGkIwlLBs+7mOiSqzhBAHNWlrApr8xlXAaTG
iQLHz4IyA4Onw7Tv1Ny+K9q+/a5MDel1llNWa220Spv8GMgC68WJci1tu+bL
VBJ4vOOPkWjAqv1ZZUG2dFtz0nobOZKx6pHY7oVzJrFfG66KEDL5RJUoy7vk
IYWzJJVDdtJS59Uu4zW2nMe+pCoJvK4uCqLfaFxra37d1ExVbFJybSeo1CI4
M9jGbchrS2GNyqAo1erq1eMReYxd/1ymaAY6R1VoEMfDxEH4FNnkkBXwE9rx
tOpaTLfx779PuMJC47FmF71+bAW5q33F1nDy3v1TDnSJHwrfBdQeQKaJr8g/
doTpspOl+rCwgLYhKxnhpTmahnHjk05FHGvVTxONfkbgu9tPG6hTsWAfoceI
KMBS6Ll7Q2NiKeeOA/XhH6ErYO0O9/WhGofoyvu981dqPpdjwAff4gjmytn3
n24tzEZeLryBPsP/85xYb7wWJpzvfDcEQ5ZDSPEYiTSFhd8XY58WBqzBIPXX
3yzza8fGAdg6PEL86khBAYD1pXKA4FV9wbTIvfPUpzp6uzAPr4Dg+Kc9x1ky
lheUycyiRyutqu/byfIRwO1j7etvT/+DNNCIrtBT3UZnD9s6/Jmc/YK1JKvK
LGiM+Jq3DWk3n0rHe1YOy4SpXQCV5fmz7oC3YotynXesMUEP980Xez45tWZ8
Z/js1qrCECi6lDuB3aIQoaqCXOqlqWmyl1FZrTNusp55v2sEGTwkuHO3EFMm
tyHp5kQFQKkwMcQmM2yKtJDAzaPQ5w18n3hZLfzlmKtNyNIe9FiM0WuopgHQ
yGhWYU9mW8ikUuYAb6URskOrOzvjZMh1w2D6fJIstQGUBOSE0VbtAqCiI3Sd
aLsifi1lRPWx1mBJGHhx5+7dZL7QNBVk5cNlFthtxYAy/nVNoE0oBKc6kNgT
GGmoSVsDFxF1lddfdZiNQ34IZXnILGZRaSc4kvkZPe5X5lnnbqlQXxNj0jgo
tBC/RJrEH1R6A4VjR9XVEOdaHvLjzp8sAh68zGsGk6D/HYnIv98meiWvvGQG
i0EHn/6wt6XJOXmjDrmv0yBQVrisc6jBHugWaxih7zA6EqfH3fur9XCNF5ER
a87z193NnT2sTJj/B1GrXIIk55i/WpRuRbqEdgptvyXmTxwczyOoTUd7gmhG
Qcrvr0H9jP5nmzn7XAuBrkTDJBAsxYxweoK30mmoOIjcNKPg3uXHDfMy0auN
UgqIxeqMycNsmsGfnXrZxkvwp3drOhhnYsb4vgy25sYZeeDWQUJQPZv9rGiB
/WkP27jMGxo9Yl1mb32zHtKW3BehsZuXR/FpvLdmlfGc9tcxKNmYACS7Al1E
qNVQtKPobCtynDzmbRcH3Fm5oVQK86neC//fZ7bo7Q5u+eObvYZPOItI+IHc
YM7Bld41MVwGfC/5WGhlpDdHCJQWnQznQC81BJcATvZb753WRWsLyxyohcip
YwDldAXtovlQJc/5e8+JZWTQ6XezBHGAR/uDZLR609uUUPeLf90C/PGq4sOm
6m6jvDUYrCQ9zTyXgCyIf50YDPNzNrPHA1pnzK5iUmJiug5W/S3/j+5PzJon
vuU7UUlY4NaIMNLMaj3hbbKNrxUzRa9+p2bea+KmIm6DpFg2DcmmPwtldOpW
gdDA3pvBhev+1t2NNsgqVF7Q9azdxHPfRd4kl8jjtutt3OBBJf6dCCpvoq5Y
LceFaLCRBorfa7YD5/VMqv/CQWexPcQdmiNUNCKXpogtaz6mFvA7BXFSqWfi
5Xuwv7PXSmZtbuZWaCTdiHdb7YP4e6erGP1P8cCXXxJyUET92Cv7JgFlLNQ8
tkoLV/UgzO3ny1/RS4s2yfuGi32v0Fbyna+e8f0G1T5mTt11l5YphN4QOkVV
LiPH/jMyiEdk1v26qCtLxmRX25XQIBBhgDVgHIVOEeeF2qC/imCOiJYnzLqa
28RQfhgIsjmfT5tlPE81WR3f5erzNrUDJkk7LB9VTVJAstOnSWiY1KNb0Wfd
xwrRxEwKgHKULpwCgBFNWsiBaxMOoKHWebk42hT5zbLpcoHIXbNiQBpm5cd2
AnjjpFpVCJ4GE16Lo4R5m6Mq6Zy1yxvOdXHpnHO1YFccGnT+iWoL745Id7r+
AgH5hpfKPXVIhwxGtBZFdVntDmNvvEjA/woX+neB4D8R3D0BUPM3MO69W+1s
6WVH0H+WVGo3mv2479rxB761DPPTMcZU+AHOOG4B75FhQmA1dPKQUB2t1APG
+t6NZk1dwHLiEaxTelqHSVA3t1cD362ZawtjgIEpEeMFAbkhM0QD7Wr2y8z4
7p4hUk2tDHAZOqxrpTkXwyT+Z1ePbFlYte0b+VbKKwqTY2FzwBLh6fDw5fHg
0PGfo4nv04V+xOwFn2gSQZ1K3EP3iMUS8W+NaIxnFGKijo8zQfw8W4Ut7ZUI
YtMagQk//H+WWtLv8NFFYX7/58b4v2q5MlVlZFr0bGeD7WVcjRKbQDWA93RP
XuBB9ddZylD5DsYFwsB/QMzL5Ou9bk3uos2X/aVYy8OQPT2u4wOoYWPtylf/
0J+b70yPB2Jba+b+DDF6MJ4LebtXDB4CuX3ccWB7e1hq3IokT90yNdmuuVkx
fHme9Y43KJAt3GDKwBpN14g9Vpcr1/Twri2d5jjzTbqnI8/VMHwUE9Y+7KzK
aUPkgAXeSajMXcOSGbzt6VVewHrjRjjVBn4cPSZOICgO3T3n3lQ580SKWBpj
IzxnKCQVWa1WbVG4ZNbVGU9/ZhEIEol7K8j49dnNU5pJJSnVNqpUMQj69Bv7
cP1clm1haiWjF8oMk8BJLGPYZcjyni62EMi/0GeQISvf2ymFNBMwCVJKntg8
eKVqzxzq/uppFfOVXJ/9BgmHMjEAI6KgIAlNpGPw99kA7oR5BFjEN3UjZaX8
nb2rz9Y0jN8bOIfBV151oy4XU6hKkPuy9gIEMYI/t2DnEYDxr1O+qA8E2NSS
8LT1J1XrwEAn0sOI77ou6DnvQweTtdBh7yoSb+oDQke6iILmD8bDiTdn/eDb
BjjAl/c0r+vcZsZDpAklCBc08zz1aQYT+VV+C0f1ruC/iu2ne8zqcOy/fH3a
JIc5ZRDFgyHmqYBLpOQnc6qutngPIXk0ZN/NfsFowhI3jX0oRVY20k3bl2s5
v0W/8ZLnm1rZ5MhlZcb5qEutJjvk6S1NAgvWZ2cfOS1HP/mk/+/xXlZqKSDb
TD2VLoVL4J95sAfXC0gfQag4sXOIVov+aYPSHIr3edYwSgcc8lSxUAGB6yGZ
iuACvk+JqvoxpZiCx3a1i9WC8Jj9cHTX7sI6Nvhgd/TWpqHcLaFsLU2W3m2f
rc4aWpwjV8FYC7x0mRhWFbktTui11S8bWuPVrGl677x1cWdGKCtuwS+n7pd3
KDvYv1FFPmA+OSJ2D/g/KQOeBYloc3St88uk9M7SwQVG79gDIRHRxAyAJwWa
i9UDkowrJXSVFlSYYdTuwwKNJyL4xaoo+ciG8gr6QPcgB/b4JbomVUsW0nC1
1UM8ns74YTLU+f/FpAsYE+ZuduYQW4cMEGKdkAFUV7O5M1HuY5wrrsYteag7
Hdg9kKOpkx/nBu9iZ/g7Z4wJUWooC8ycd53EV/x8ci2nUQe1+nJk8W3+W4Ku
azl4RMk5l7NUDqz9WZijcLW7o08eCtPEF/lRsmwhEEnxnvLFfbh1FZOA1Sob
PMBj6c+4MBh6XaIQRPZ96EVoooelUL104hg9ui05XrNmE0teWUqUKQ6ZkraJ
A8uFZyTZZ+PMjhmJ3YzeVC8eAF6I3x7Ei40nu3ANC0OzktOUFlvcr3bh2ZeX
RxnVVvWckim0r0I4KLOW0CAuLSGLmjyP4J8LtSzdqVky7pnE2cGMlZW8Cvci
1wEnnyuOBH/+/POTjXOzFR5+o0CUBPhmSZ1GilB88qZqSM1/g3CB0I/NoVB9
nz77Uswo/adN+7r1PI5ONUzUTM+NZqlAksStWbrt1HyYPzRdzHAw0geijZh2
hdbyZPeFblxRSRjW7NzCtK3x8W+dY9pKmpG87XUk+nP5hyxjIshmuJLE9mPY
ex78O30LH/oRpvQFqNdVZ754PMcq+kprK55dNdyO5Hpipl9jX5iyz2k3G85f
Dm/1NhIERNf2fYGl8Fk8NOdTTmm6uru9kuwWn1JKNkZ03kMogxCab0AwebGs
FTeO+jEY7ImZ/xvZDytAvx3hhHV+FaPv7lXR7jQMM+UvgT4H2bOqPFp93UKt
RLadRYlWv8jw+Wz1hryTO0Yyxja/6H9TfH8bj99cxfYYSfDBYJezlFekgsyu
SLrCSzN+7LtMsYYEoS4WH8PGCtLUfIqOkDut4cORAk6ecXOt2k2X8HMSI0+U
eyf3f34pyQAKtVMDoxl9uFNROL0wPN3DQZFHvOK1KIv2CZgWpA7IQRvIzhCD
BvsOGUAR93S7zhm/zmdfiaJp5JV9O3zxbG1GnHrAz9jARS8S87CoZCBBpf8X
4TBR8+010L+2w4PzHOrPorF+qRjE3U4a8ujMsymIGD4LimnPdzbBvdgSKCZD
y/DivA4gdgjGJyia7xhjNMU7BOliMjgRj/+E08vi80m0mt68IOwtd4pVL5fH
IBEg4j4dO7gpiIMnEaXXlYtRuOTPeDPuMKZH5jbR87tfvi2mNvv9lwQtZJmF
++2kqeesv+wrdmCmpoWymJJhO10xwK8aWfSk0AgeeI96u9QFR3z165jPHbnr
MC7+rk+stlr71qG51r9c6kl3h0Punp7NJpUnKiIwvs6y6erCPUGYLX/ioo9P
QvePJraHRriR/GPYAIJ6Vpm4e3kpG6kMnpwWl+DBGgp6GhYm0fTgqs/Mrh0I
aWYgkqnnQpiA8dhLxBXyzSwDhRF2pLqixRJcAGLmBUDbrT8w6lrYh/xHOYEH
GN2whtJnLdDLhDgL6/2mMZW9IfExsWVO80ezKV1+XzB2JNUc/J+wJNjkgGqZ
Rh3FyGLljC6wYauFCoG1nNO9zlQsKLWPLksDHwLCQ9WUR6zggDOAHsnX0YS6
/GX/EDB8wtBxn032aX294vELD0nMaVQcWk0pleWGbAZXHj7zfXHcFq3nBfeR
/22fdBVmRDuQICy/Xc40dAfUAXH3m11qUBP7xMCX+7nn2DkJKcoELEXNnxfZ
HyNuHzI9wiBwtibmlNBoIDdPICVqXhaJE2a09M8A6jghnVU4Xc99u1YlaM4b
ASBYGIZtuM8Lma8z184PBIZm6OLOA5kR5yuZO9VeDyuDVBuhh4Cxm00ENXEO
CUNA7mplLe4YaU1mLaaCLPvbUnq1E6SE5ypNwAyJpcdbsX0/gIU4VIPMGHZT
6pXg40AJt28PxpfeVY03AvyxUbNmd4QK93yrwiB7aWK8n9YR8idQRX7xQJEn
zZ8uWdbWKQFAoWS4u+WsNI89Hhz0tLmVhXFd1tH1GdkrGVZzRW82CydFmy1/
raDiZP4XSZUBcnqXHhSdB3GgEMa7fO/t2L1099Do5b55AOyAR4nlKnKO9rnw
k6vNhkdPvtMPf1EEacEq9Z08oBD1SZm8pgVG6TSlN8QllqnGrwwNOzv4K7Vt
WEi3MW1B6HAfvIuq6sx0z8jKSm3FlpvecaV7JaD6+oDh5BT6eh96HafR5dgk
aelRG8qYmUcmeYdHko8JXZildccQhSAQkvjejbTmHrXMJ1h2GgMngj4Ju+hd
K2QCpp+ggH6lf10Wcvu62d0J1d8OYrHP5P8fArx3sMva/dH2IEThzo8jKV5+
V6+LMKa9Iy8uHtmorVJ+yO/5eexr4013CSP3qAPpJYFnEzLpy0liFNI8IaGd
QYIR4Rg36slBjsnM3IhF9b5vtJ+Xy957U+7EF+JRKHy6SjAdLqX8YfWDRDba
Zp3wh1mmon29qXEGOz043yM9j2mQ5saockFKgNjXGqwN7ZGQeD5Nsn2yL5zT
kcDqOQRGsTTCi0/qIONTREHitowoE0zooRIsjTFlEiwsAKx4DGOkW8OEaXDe
aSddApBeI4K0x7XRnuY3TGG0Cx3vIqEU73e9/y2yHNi94HAXA0tVPY+9zqGl
TiUK+Z66JX/U0XLQLPOCNEpcOhzpXMD0sMvuA7Cv4SQmQfP9bXHWZ2WPd85u
zOBvi03m2XuD3m+XkbI+Ntwu3MRDQqVB6S8PO9rTOERcKWxRri5MnsSegjsp
aqn0SM/7Qg/68cL4GgO1Rxkq8RTd/qHgk4QArkrBWet8M7uYiW2zoQQ9Qtu4
Mc5xcfSa3iCJ+W5AMHQGT4cw7aqCtvpaK6rEd58cy1a3VOQZT4PoQuv9zDMG
/hdTCu4E3rjy8GwxXnOfiWRTmgbUPtq0EBEryGapA3fHjxwK8KkGiWa595yF
5j8dgKSEkP+EFA/8rCyp0vtsP+FdGuB+RzigfSpy9Ljhfti+DTScX6AJwn+W
42VRHZhYgoW/JG42M3YgSUUU1iYWvr24pCC9ML7MmhE6kbg/qAELxFu23BNw
pSXXrw96RQFXIvZKSNptt2iFAUbQJ7x0e/xLakLGnm419M8iBkMkEO0WhYjQ
T57Z7P6lQs7dpXwU+mrd20ACjZRpP44ZtBcv0t0J8iZbqFFsOs9r/Yz4SRbS
d3lSW8RVHIEGB3z7BLOCdgxznaLUYJiGzraeU4CcSoyGWXeZp+fBAuLVa+VC
/EQP11Ct6UkTGbCaboM+0XbL7oJbw9gfC5IgP6UyuG2kNEIct4iW5zv6Nx3v
jW3q5fVN9s6nfC3Ev2Pwue3Pi+zRVAfBhjDz6Ndxt8CxNMyCGTmxH2D6+/gz
uAW+YVKEqiX7NkMgDeZgTo99azrP+jdvROE1JxVRw/yXUg+bA0pwV/9n0lC4
A9d3viJrddQ95oXgfob0nw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpejtQdBy6jLSntqxEdocir0hBUxQjI6XvaV7lTzVbdOFk+Exz5KLUjXsy89YD+fhX9aeob2A+oZyMsnc8kE/59j04FpIPtdzS6F3xgwACBZ2l30IqvAOXtsPZ/leOp94bJvnkdSOOpbQUQEv5kxCRtmfSi6m0abrUnyzxUTY97d5vW5ihwZuxbSI/r11mtEDqAjjWv7josDR9X/dRbf1MKVikQFgmw0qu4ebwtAYiAagsR5XjedJYcTDis1KZrjJXi03/jz/WbVGUYKhrKNmG3p4iatmZstrPhZ+hr/84MahAYfLrKv3S52pU9BmB7+/PQHcY9CPbRWbkRqXWn9VTxTu0lKmpbBKsfj4m2ZPBLu7a61s7taoObudBqODZVIUbcYNlCwTMsKyRN0nO9ZdHm15jfjqAylgsikQ5Hk+Q4KP9aJBvCeix66A9tdqFgnJNcflDhbz7IBr75tekk/OyF1IQuYix2SOoq2QzZ/Ik9/1xZa0nthJ7ofuDG0FkF60tgDHPY1biT/zW9d9MsGlIW/iAlilgx7tvMH2byfeY1EVibLi+psZKjURHclHKvOw4km/CTdqFw3U+z6GbmtdhRpJHPEeYfmtF5UsO2WkI/Mz1gnD1f32c22it17pYKR/2HXzMsn54AlVvXRGQ9BQfGRTuJjBt1Dn6y6rPXd30eNcYj0gcbzN3cHqrjFmLYPSjbEHWpABDmskpaiQ81+jsZBvO7F2BcUQgdc1W+FWsyXgTy5pf2JZeolBIxR6N1o2JrDey/ct5WTKsXZk/B+eXqej"
`endif