// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CYs6cjB+bSi/5UI5esKZu2PdJYXQxsBnYBbAiRWSisgea38lD/HM3D+CwAob
iVWutKsW8y9CHNdYKPMo/zgQh3pOYK+MGYtZ8oznXPXr2e0bG49+inP7wSYj
WFOqsWVEW9r1gBkXLUXO20ExdJEC3QtkvqEb+vFZcJrNIGzyK9l545UkWeWI
kI8QN7xpSuHaGt5ySDrN/xOLEDp+FQC1Cw+6cVxckeLrNkNy4Xc8I8EWeKnO
GBduo5aBkF0cmC01jcB0TapH9MczRpqHDCe4OcE1FpzKXODlrBxXtfn09+Bs
b2X1Tqfptv9PkcB4A+MqpSwF36InTZh+Onuy5XNlOQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ABM0QdADhVzDAyEzx1GnySP78kDyba6bniqZ4WKjAPwhv96QdRo8b7PaL8V/
xstqDRqZA+TQxG+39M3uJemjsZ8Fg//lnjjNbzKqJHjPlHv4U+U6PynYFDWn
M33MoamkkaQ08wWe9i229jTGkGjLu2MJDUilRwl+j046K0SKYQP9XHJnCEvU
xFJQar/v90GwYJfXOERLYgbBUReL52C7iJkPYsilz1dWAGAapqCptuIISN+D
4nCs1SFmmQj02jhKjCmsh0t/lyweawQgenB8Bf94xIYtlUE1yrNNN5pF8K2l
uYoT7WjZGWAA+i3vRhfrZZ2rsLtv13OHFydFsn2d7A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kyQ8SHNb/kGbBU2oQYfWY/Cwrf7bXcftkoDRzjvqvhDjHQ6V7ywDDFz9d5P4
At9XhD0N3k+P2yX4e9bHZF59RCjnekHszqc1PChlrYuhPPfsIW1IEmq9jLxc
Pua+FwP3y/jkwh2a5HniorKyh/yz597ZvKb8NCSIJDhrwjB6vCQZlvVBjjQW
eFEnpYkOowez6txxAehgCKV8wpoyyUVRFQFnGsNJCAvttOCT/EUJqfLZolzv
vLWjLwEKqoZX2JA3b0hLe0n/HxlwN3ym9zF4CsUo1HsZd7IxiPDS9gSHV+65
RUjlRkbWnfcADNf0Yo6Vh65vyoSCYap5Z6/XIqznZA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cF6RBZkVW1RTuVdJWT8pqafsoCIR9AMvRbDYu04vAklH0if8EtNoj0FaTuEH
B7plWiv4DG96oUan4FQ2MmRBUQEsP8jjvqY9cFHmieRjztNBfZ9lhp8L+SrP
keKtQviKz5eyVxl52ax1cvX19OEY4Qx+VgNJYrA+lstrUM8Saq6vMwnGupdm
OZFQkhkMKbybDvpAtXpjwVd9G1a6iqkxGoye4es0AYTQrU0ay0koVl2g87wR
HwgCCOORaPUdBCgNP5gksfcxkt1VKdIsi01uky9IX60jvzywBiVd0HMRhd/e
Cj2Ljf+ZwfQuxyRBojWn+En6SdrCE2Wvl2a/E7KHTg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JnyVnKLsLq6yQZ3qbNqQzHJPNzSmy4tDWzNUHQZBbbRqtcy1PR/4kUKD74ZU
/XmxoFRX12yGeMytdW3jQwXeXPjKXyboQI25eYXz3Mz/buVwUlbOgBa5acbS
EMB2m90QdUafQp7Z2qupX9m0z0tSVoGDwec/V5h4yk3sbRDm98k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SKIEDbeRNtmmp6BDUC2ABlHbZu4gE7TWJJix1lWw5Wv7NNJ4nFsa1IUqkzwO
eunajkotjWJJvSohqivm7OYtivIE8InnUQ5kmew46qXjoMTufbKbJRfR7LPZ
XAh9zbrn/ePawqdTn/lmgEI2SbBHoh/1+GDJ3H/sezLDaYvirm4KDXfLLw3N
/mc8MG0PlbrIDNVJpolfVSRIulm1ZXU8xn6TTFxB2WGwBPAaYd/hkmiE0g6v
KgGK7UnU7UtBpwScxTIB8khoUQx9RJTtpzoguDKOp0fib8Hj1l8exAJ/isTf
g60F9pVadWUiCPTXeTUbqsEfJ1UfL8mEYSCI0bcWYpWRs0cTo1QWifStSbRI
ZGyhiShm+V90dJaLKMfRreDzb1hSMyBhzvKcDH561IMaIOEOni7zOZIixt1k
V3QO/pQRnycf9WKobttaB/koIWRpilUns+eeievLjsvtiG2V8k/5BqzX7QpH
eGH9Y3KrGuVimQ0JIZNTD+Vl2x8kJ3Nd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ow2h+/wJKNRqrIFYIIrjaQhCT0nNMrgeRQM8cd5mUoffjvxDfa753CwCzFSu
eGY4V9+PVQShSqxT/HVDm+Gl7RrVoc7vWhQKkhougMbqUpjupA4gLqRE5o99
TbYUdgBcbT84Rmet4Tl5IPeQiwyx78gd8iQucdWxh99+Z8Zmp/w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n6mlvOiKdTwxxfsaW4XtVmay58een0LrjTOtGg2427m9MdwNVXsktdR6QJ/Q
UAnd8WsSFiMoQCfhrmskHjZMO0BkX1zEOAyN17kyzVOijqn3do4OsWIcQRDI
pFEUAiOIbnOhLZJtwNjPttCkKLSit5YgG34WHJri5fkUvVo36fI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18624)
`pragma protect data_block
m0kT4hOC6c4KsvDrmFsz8rpEkzl+mHw7QApQE8NyaiINAdLcDlFZOhIYaGdN
9WlRUOoeRbudNSwb4+JvkleT6qbgO5OzG+EvqPZGBT80b6XxMvU3EBtcC7tC
ID9510ohhfjeqT84gMSyCONF0AvDJlsj3Rb9PrU+C87uAYZT6vqLB07Sy/3m
TP8IvsA6fHLwoHLqyYeRtXqmeuPsI/33Q43d4pprjJol/zuG4wHDChnBzEwq
uMbQeqK6bUeDguOon5kHpVJPQopr1nnaF3Lgr4kTAVVqCO7qdHONF8/jk6QH
r02hiC3zOK2HTtYpgeqo10d9p8I+hxPK1IJ+1+eOF9eyTtak6JCQRognoOyV
+35SGVlv41h0OSVo1URKuA+UnOFslEoivWut3ewjh30jwgABzCvhbMrohfC8
wG6RzyMto/fpqJKf6ZgJPKVOiweOgsL4vcgt/rXXcIefOrIXTIM9wcWXZJOE
t4DRPDiATt5VBKSHQ/EuaLSLM5j3JCbyOSyxoznpJzXOVTlI6RGQB8URVb0p
YUgpZOWVjNs+CWkIZ8GpuxUfQ0YDZZkxkYwwUS0TPY7QBX7BNEwuTRi6M5vi
mmWU5aodyHBsT7HMGMOhFpkTX/Pk1jzAbqxC1jiuhA+MzRBEDuzCw+jJkJld
gYCQ4KkISdfhBwB1DF3uc2b2/mOdER9mOkcvOr5R0tuRcH3wiyTBjB+Nr8se
weyRIvmcClPXNoTeg3J7pxA0OIpLoe2UbjtYkBzRGmh8mtLy9gKxu7ChUHVk
gKFcAfXv3/tFXczrQXU8C61DB22ZEZ+q49Z8IaF5RmSaldsPCAetstjJbhn8
iRmfG++f5bvBnm/x+oUr62mHxEKucc1tbUdxcJVDlwx7VFFbQCGWRJaLCGst
ijy2Joa4BVQgcWQlnfMk1rUepr92npTsdYUuMySc3T8LNit6u4wTljAw7LVT
lH/xW1CQCyNYGuSkgLMPl8lD64k991BbdcQIaroqw4/ZTGmPo8tTZuIoFqh7
pDMeEFeTiDSh6OhOz5s7T9jy78SfKzBYPhFlxliJ1aBYOjag1P/27wGLbTUq
lKTbQpq+I0ZJayTvBzI3x6I6vP4uoE1t/fmSqlahijIQwhR9zk+g1V059ao2
+yNrkA1NjVCQyFVJPWgk8yRzA/TsvGgetvkYCas3mAOCGtxiQvbCoNQQMP6t
CxGDZUDCLOqdPvdrMb7dTkXVbAAiKER+roSAbX6ZSuqF05qNXujBfEAVFjrV
D3BUfE0kygJhoHtpLNa4RJxu4xXZzYXolnNPI/e/bg5r+ZeC7PY67TR6BN8e
OugJfX6bizUgMVAceEdRvjA9mbHrRm7JSKgdhsNr3PIxCK9JoliSa+kRqd8n
xAtCkDc0Q3RfJR8ZXfoY/mZmNZ2FWaWaMK1VGoWbILUp24me4rDMx1JjCKWv
L7z6Vjafotzqk0BVoogzrBfePRbQBkKUpQDWb7l3n76jEmqmF5VmQRf8om5u
t5UcwM6jA0kLgtdlq7PbqocbPgQhmRSUnprlHk8P/N21OF3cmAKJQ7mZqAip
WcwIDKebGh3RuD9BbxxNo1Owk8QolqxHxL6RDBB7RvA7zvERSSDXTFJ0cTEk
/OyagnDxMDshQpzGeKljj1FJQU5NgDO2TdSnCvKyleVcppfKzqNwvyNSkDHf
vvGDjB6gs1SZXAS5eNMV9ZoYv5xvCu2mRIy+outJNHjybizpYYW9IBHUp+PO
NacD9bVnRGsDPFsDePxO/MPEnVEmkjvFX3bkhR6/gxUkEfJP/WwSvuHU9Cpz
8SRPKAhHV0plweXSt7ZdPTSreWbjrE3J0j9sJwSN4SLMs3ZqUaJoN/FRchYw
JLClOSIkBFhCSCHklWtk8GUzSVqqJqFoGacde3Qm0AJsxa82+5algvaIQUw8
5X/qPGg2oTzNc6ovbXC26aLB9T0WPuZZ+OPYL6erRy1Y+CFBjuhAmRE1uROK
wEUCPtcqEHKBDRJpvxBpvBLBv4gcsCkIM0QjL9Q/EiylIqpT3Uby+6YkjMim
PLW/wsrLswKDi5StKppjTeT0JVlb3MfahefdmmrOOs2ifQtJHyWdMLTLjjh4
s9DZYrbTM6U6PVIsS/0vxV45zjzwjuPkGcowDROxnfUsmN8Wkjln0NfQuI+S
D+b37bR4JfIw7yf23hHj3PI3FFkEhVdMjE2WbJBO8+W3ykwlAPGcI0OwL3wp
fCwT4JI1HzUvwUZ0ej5mF4rziaaelAwJF9zEQxc4A0xRe1JFqDB/OZMDDAvE
i1XaStvpO7h/UKL4B5guUOcF1YBCdrHEOgqhvs71xc7mfClqUc4Vgql+7sO7
wjThax4U6Nm8YPlT2SdSsHpg85fV6lqxEoGby5hm9UeE3fWDJiSghQQi0rUB
WFxd91GPLr4vTRlFS0stKs5scR/MwVccVLwBekkm3C1SxnUajz/9xgykNsFV
jH7EUzcQZmKxVXgTyC+W6vfRyaKOt15ljxckpBiULhCDwu9km/zjZ1sPvWQJ
3/KmOJii0AUBJS5AhG8nNYtjqjK2VvGLyVU65O3dGZPPP9WCqfUYezHy/QAq
i1kirV/zBXuMGcgLgz36CqD4lVc7xw/qL7XqamZwYy9JBJ+D1PnsWgL1ADkJ
30sJ56TY5MsAUiTHYGnPpIIqLILaHaz/xU/P0vYWb1StWETd2KpImn4ozKQa
ChFw9mnU7udTTughnZ06lrsDiyQDWQVWme6XVfFq5wsmR+A2kpPX7FOqXTXe
nhr8+nrQglSdru2J2e5SHtKUGSgQTPw77xVdX+VbIpY3Ig6JbGhy4TZSqEqi
xdmgUueFnbz5tDN3xkvOl+qhL3pdwehMnavap0s0TMwi8Yj3uWMDK4a7R4iF
rZkm8hmgHHRz+pVg6ZBLx8XwHdnSxpUj2ESzMx9AxWbKGSgH0UYrZz3gmG6Z
+gTupf4VZsMkjcWlRG2S8gBUidmEUCgjZ3j6vRypJhE2TcYIWwj1pO2syL90
lTeZ92Mkg/YOyUO5yUhWmPXhrIOb4Cw+JnGRYKe1X14QOj8aEqrxWozeEgMl
iR6kg1NfxtPFZ13ppUrjhmmahcgjQ8yVVl2NTZoupbuc1hXT8/sQzeV6wNiM
oTbTsw024ifFmmbnoIgztehuR8gwgu5rxJcuwgpUh2P9HI655NtS5ryI/Zq+
sfjVmoVnnU5mDiD8+PearNpGxzQN0SzGHWRbXUumormMiQgk7CBG7GsFXaR+
iTIUH11r0XiOcRhaSRqvnjHXkLLsRjhkm6+EgS8D3hrKJP7uEVSJASXSCBHg
N82Mkw1dUAJFqVLmMSLSnl5bTcldSrgA2z0hH4Vmjz3iT6YBpuCGZISWgaH9
3FjyHrR1ftGPz8mou900AVjgTBizFALjYA9EPsFKiHfa/xOy+1gsptnY8vYP
VStowMO+RZuL8vCA284NfLfiJ5hyQBZA8cUxPffoZG8TL3qLOZktzsII49kX
6xO7pTGS9vHzXzgNhA+cbqNyuZn4b3sUQPnCEoXzig/qpoKZgpRywN1o3Ipq
0QGtV+TF5hIBXQd80VtI4Xt8/kHQ/Gr1EoBmWhKqcFSnLy4Om+8UKbOmAnw6
t8RCCviBshxDtScOhrY432hTqfh8aLdfDHQvXFxFQ5hjMaYNHAHoXw7Itw0y
+HLXwl02B0IC14kO0hMPzicRuxP+uwdZ1AJwd9bz01WkadXS4haCuJCbuVxG
Ls8seWIhJt/CBjpTt0hYlTztTXUskwVm4I6yM/eE/GZpxngNsn+17hVTtgWg
eW9ueRK/sK3ELfDQaWTlQz1/a4RsnE6U3RtDFyc7/Q+xZlhiGn9lHX73QqEk
ssOj9Ao7aZmCXxQAlnHoHg3YPP101D5PHuVmyOHkZ1/TsFFJ6eTuOkfjHQVW
cUr3Rg7PYi3LJkS9672+O+Y76G+rZ8/9CpYmvLGlv4TpdjfewvGVLtdnDEc0
rLu6xHoOLWrPpVWaRZA4YaEodjIr9/EqtwUJ+OaR/jXkoLLYglRo8ownMViD
vHet3SJELK1yk2zZc+CRijvq7Qx2HT8U+8FeS7KZ4q9L/NCx1pWKZwze2fc1
w97sQR32QYXyp/VMIXidielJhddEJMCXMZ/E5g1FzNWTWywC5Ou3UsgkvTIb
fK0vUbEDwjGpUtlQJ1JwzsJv8iahu8tdriEF8vT5eLmj0ZSaPxA2aduhdHLG
6JDghK7wvrwiZD7pqQB1yjTo5N0FQgY+RYPimunJ0RDK75L1pyOHMEginv/3
qJAEM8TffzQUvAjHHaEkbyzTzwlF5QMAP8sk7PJoTHUCMVbVr5ZNqc63KVtw
LGM77S1XX6TMhTwH5nwJWnNcIr8AubUnRZQ0i2ZOEZuvUSGQmadEYUuHQj2z
50MWsPrmZ6XNyq6KJZnlYWxLtmJoy9Q90sv0G9WfZBW8MBIoUytw1hjfrMHv
bOGew54DRKauJhe1NPOA8Q3ozvinPtdXzEsHKxJ7ot542rJHhzum4UQhSHCZ
Vlmpebl02gdWAIGSAHXj1P2tElBgxRmOZcc22Y22Qxoo9b3SPP5PLfbk3Gce
5XYd+HKzvzihOZttY6fnD6oFBcYUR8yXWCcMK3SOoegwSbn9FA7j/hMS5IsO
j+l+b2KNX5iZoJj7oV8AoNrP+u+b0AMZ5B381JPyefoL5an3Eenyg/YI2cWh
d1b6RKCyhTXmwYdYJ5v1jMLJODM3Z6Pu6ZU5iFSgz9rJgF5Q9SwmejOdxYtn
3htZ983PNs5hKtTqzuVDAPhJZTVejd1nC3i/Tma1P0X5paTANnqEmDfUTrIv
qdLpSfHlfh4cgIHieFHxInocAS0xoY6hEF8hrMaSfs0whS9GRfAbT+GfdiO2
okaqbQ3u2VzBjaD8Q52wFZ4nQPZknYVOCw+gc5VCJ433OeqTr0VRfLkNJYtb
tuR/s9YHlwvLzlV4mjwBS4lBtcZZ4FKVXngKu6KfHxTwE+ypQyy8tTjJQg+o
tODOahwVKfPCGOjH48Bj93IVckA88hRZXrjX1WzXOlDALH+f9XNi1UT/TFCR
4Xxk6TjK69Q2TbPlCxcwHArkRxuAISJMrxtiDNfDmD+YUY4MnWEow7AtwLHN
x82LPzcBsMHeAvnUY39Ba3Vk7tcVd1A7yj3/56mBtLBZh4rGHjYqFHTFfMym
Zt2c6Fb6Nz/tDtBSTcOk9nRp8M9nt9XlahbsSv9HT8FSr6zphy3wYWUmGPrU
0Z8olmci1dH89ccE7aRlogob+TnFWcMbvQDjg7XGBNDzSQ9QwvFduxTTMsrZ
RjmWGvHBeD2WPtXXNesZYCAHpaZXWbwf4Yj0itkW95O5KhRP/IxXOlMNiNdM
mlIfdy7Ea5PqxsyOd+7eOlM+xt3ctUxrWu5nIxDGfIcsS82U5XLy63nfDmxw
gbA10jwI26T+4L/gtzfEitucU8FgDfgOCvV41CYIEE4WduVKI348KlANcDLc
QArERzaxbW/fU6/VrJXK7rYfYEspZyhmgClSAO8PrD0NQvFpNZaOeX+n1P3A
lXjvMkrYS+JX9zL5Yx+E8QmyWD74lPL/7+k/IbPd3/ImlxLUhWxBTLTbMR22
PL37vdbZ95lmB5zsoZR/TNVdWhG2AU2Ri3KXXA295U2IXEAh5Y8Ww4b7ymwx
DAGNS2igwC8Mvz3W1vkSyrF+XHd0EBTUmPITaxzTupF3DAWu0lJRxDjm8V1G
Xfb+PevL7r5EPQUywV8h7bhdO/0tb2yFnVMRuLeexsdm1XY6BU+Q5yVWT4rL
B10jQMWUsMOH9XUHZ7dogiG6W3Tnv2I6xQyvj3pHjxv5/Q7nD2+N4YB1VJPY
Db6wjNZYPS9a5nE8gv+wCM5IwEXGxwXT+dmiHJY8Jrq56nrLlVsy6JVrN4Qx
A3cZX+DyHgfYyqWALr0EeNyjoVGiAerKnvws37933s/yLup8qROsnrwNFtfQ
8iZJs6FCZCs/w7zqnDjcPnUd0AAuuH0ljJE+CgsHWrw6OiC6iKcFaN0eoQVp
i7LkxnL54uPrbn+SyD5M6YOrrjO9kk8ixJ5hHTxi2N8BjihRbbjpWWzwESVZ
+ORin4Q0FsW84BxVsWiSsRJhWxP6XOwM8kUItXBBQSGrvuCsyh3eJRD5MvJ0
ZeBaXXH3OTkhjk+yjSq6RkCswyjmmWlcJCbk1MLi7+gP5auflAdV1/XJdast
TnzJgVtcmX6R+zLo92JDgqtQ4zFVHSSe2/ARyaVOcwXgVjpoZKkJcbDlz9F0
/aeVmGnhRzDUEUbhvb3lQIlgRFFhvd/yU270628dKNKuX0Da48JERQMncyZK
PSm2BRwbQCDEWDT+vbH6AoDRbGsKP4+96DuyFJkL0VCeioKTxR5I6VFgNfYr
Vmi5SsJQAduwT+dRop2dk7JSrGm+AYdMfcqosTjHZmqGrNvndJRqORW9Lex6
T3NjFlLNjmM3cmyYi6kHl7Aw7KFvK0D26FYFbSTw+OyUBP8Vo4k+Yx+Cn7FB
yUCl8NpBpzy9AJ8T2+szxxoOAJP+8FOYjja+SnW7574DNrwZ71p6kOKAzy7M
pNEYh66ZXNIxXH9z+zCeEASre/g0o3lEm+su5zM18cdv/5qWh5zh4leCDL4I
mkeTLeKee940sUFm/Z4CNMLkI0VFYZ3L3EHCy27INnJnoDSOHNttXasFmLMh
EL2Lyf5GYbM6t9yB0e714wb6FPWXZg7t8ucsbzEf1QzSL4zl3wQgaEwtzsCT
B/GrlTeEAK6IXIE6RCRjSvYFLDZx4rGoVxL+l9GqqD6LNqfsrczn2sSjLxiS
LwL29dfWeBUDMpatnR2Q23476AYhprPGCWvl4/TS73MSrtX9xWUpttbUrUWw
PJ2Vl+lrrM/0KEkbCOXuwVKnDJqBUa4oCtJWo7PVvZPJM14CZOWKDbH1b47P
/DcLj53l7Z1j/Y+dV4xFvxo8c/yFhV2o80XFhOkNvHVQDBkYspvVYj5sum8L
ZVmeku2vDeJvpyYxSC8eVjoeWnDsiM9DmXGgAiwPL8z0R+DJ8zhkq/JFjRZx
5w1yzHf3MZnQRXVGA12zygEL+nxjgVYRgo+eifvyGEs/Q85F9XAq9yK2C22/
6PwcmTK719nVH5jXiColljvfg7Lu+AnHSzyEgOpk1luJwc2PKeoucuio5dhG
0u0xquLdMkOwExov7Wf6174cHGMn2A4uFmCHnBu3uozvfEx7orvF/CYyIGvQ
3sEfUn79J0MeyLlWqR0ahTARP9oX99IBmdD235OwfXWZ528j+9S6mtoeCEID
zm+g6jQY5uExxDKluD6UEROx52ZFmto/8zW0aRzk0yrlDeSpMwPGMAgYrpEG
z6EdHMEqsAWiVqQ11HAJREXbjWAkpu2GQ1KRk8pjpZEZ9DWG+kyrqYwmc+WV
bZyFwYuurI1OUJvn0w8X2iF1SudOAtHzFE+90JY63/8kRG5luOoo844pEcSI
BlsVQ6ohHmu/chGO5XNQUhHnoLtzBmF+Kwk9LP5Sd6ekkthbyOOWgz2Z6Y5T
OSdp5Ib2Ll+JiEjBqfqF7BVIpLCFv/E76hZl4tX+bnB/XUHBfmJDs43iCw5u
ZrU04LjAeAvUPtZk2CzsrYY++JYC06Z19ZS7dEfejHqlx35nQKc1XhdlfvKj
GBiYZUwS3iohffwTaUK2V9wLgvTnQKUJZIzI1N5zHohLVJIZ8dHbgShP7ymO
61dzZkIPw7LJZtpqK284x6jjEqVNum9XKa9xmDMUKGNN3T9ukoFsxtWSzXTJ
f0p9tXuH6ofEK2m7kG1P/QP6Exo9/S6fwX3nCIT3UQ1TlUR3zhqoXv/Is9cV
tVMitPQSpaIxm5UDjlEetBqRxyrtRG4OPswuiL+VfGUyFU3nt1UwUlP6HBHW
1EgHea/JhFLA0NjVCAv1ysBNSwBNTZIBOZJ4JXuE+PSn57K8Uh079vd1b6ee
CixaIPDEiM74llQLYPwGFr0p00acHOw+LoRxRrBjj8gQYLDZMmKvK4zSbLsy
kgwp0jFGvy7fie06FD7xvIkiPspN8Ldokytz7VsekMj42l93Dpq4F+OdMo0p
0G3vPkbSRSwPwX298svsrHxk3VhtiuXwuvMXsy17se9DqGUL6RiSaF6HHEBo
uGJESDP1+sOsUykZJpThdbUd8LTI7C+6msWsGkAgBC3FUZf1+0yFAFcIZamy
iXZYFagb13eHCDWDSQAV19M4dZ0CMQUgLdwe7oJXAQnDGKmkW3c8eOF5aIr8
qEQ5VuZ4olrx951tCL7Rj5iPe2ooZs7/Njr19JZPJjZRgubWlIY3T3ghuVgX
FoXmzYAE5GlWJdSjsq8ux7Wyj6dpZHOBtx36SkQ2EFGYsyP1oWkqmnwa1dCJ
vhoK0iRpF1XsMQ4oNs0bAxd3i4Go92W2fm/aVS4cRX4ZJgry8SEXAXumKAZr
1gEM2j0n7T2cWKxG5pPVWCSUhkIXuhAQBtKL4BxORrnMraGUJEbmV7mNLy5w
HSoSxI9LV6jpuNF402wRFMHX++vEkR1mKNiQ5USDVLfRHZJs/tdJfNHdnOjJ
MPnX7Et0s6RHgQq33RxBUHne0ZM8K7PBWK+kMF7WWLmzBvwrJpUJwR2zDFT+
uZA4hu7vyMtAA8RpqNdRJAiMsR8GFWnY9b/JXDoxg9+uwsBE4Q4p13GudAox
SkSBE5ZM9I5h/nW1o+1+403iqsw7M+8ua3bDP18op2ZJNhdjA1AEZoLlxvME
vPjpHjyNTYNJczy1HN9yZqSs9l01wrxShY7l7UqVba7q5mUEVmKcJ8ih2xyo
rd+0/DUqAd5qRKLeAydoO5upGB4vOddOJZmoYu+zQC5rPCm8Vuv9ofzflUIG
2HyyQgpPmcoDJrPznc7l2P0X0X6nqjYrwJzZJPqO/6kDFcD1zRQST3Hl3Uo4
KeAOEGWZFgnHZAKnmBce9TguYz4jE1P8AtDMJ6fzrvQmlsEODhYz3dY8CUEw
S9JviS2UeOY2tXA2+0RgM5nf9bT3YI+ohVoqDi2L1NhOOeSMeS4O8YZJ3DJM
LRt3Um5iAUzg5TQ4sIeen2iC9WvA5Cs1Haz4CKGs9Yaxb8A7Ca59spvwKDwI
MW4Wp3DmW5Kn3jStVPJy6G0W/f66PYq751k2HE7Tn4xg5l453t5zIx0rDLk/
TlKua4YSbW/Y1eKV9tBet/4CQ6Xran4tMq4j9QqwVq/laP5CL0hctHXAhnLo
J+4Y956K7O/r3SXrJunoHxOfsbk2OeCdpa8pqQBdlc32agOHXyQ3lF3JLoYd
wiToy169m1ScLH+eFS4JR7Oev3MxvHIvN7uUO3xnte4YIbWafqfpsukgar3A
zht8p8Kh+v7+1n1slFGIE7bkfRooWbA+dWcbsgO9glIkqcsD1u0fuTiq6uaJ
siZ9WQ1nDm5uCruwrz6+5wNx1/kt9rZQ/I/bEW5zKJoUpNcUhoU46Xv9Njk/
xkdSdiDhTXijaP7OsmNj3PeCaTPigAgPQnjt25wsd65UbCqC4+VwiwJ8Sk5b
iLtHyvamlBTbreu1336acej4cB5yNZzGOJ+6bPUlh0ZWH2uGTzmLaWiu65Iv
s251qLsNY+NorXFmg7PjBKlkjB+cPWUY9HaKYHB+QMQQrgXXU9lrHtJe4onG
w6xPbbWGtqhVk1EClMdmZ5a/PAl8z2NSvHFiF2AEDuqVi940Ce+obZPT9MkA
ksxKoQaeJ4s6xPJ+q8nezrTWUifMuMOE1qfx67FZBoOOLrVL6aRJY9f3D2cP
1NBX0IP6898ZglP6DiMZnuVXalNHxPy4QEnTF8LDhRw3guT7KFFfZ+cSynAr
Zl8er3Mv3sLEV/mTKxvHlkca22tlg30HiNrcAgto+gr4bqTPa69AdxQlV4ZQ
FhAkRrKP42K2KE+fT1M4KiWncja+i11t/Ws6ucFXbDMNASlS/nrT6a7k97sL
wIwqR5DOULuQ9d1zD2SePjvHQvgBZ8CqEnOLhBKgQdAn2pCsUw3FPmOJuVuM
HQXB1P40uOfjYvRHS9q1rjtsgA3tuKIITeQyqkXILpkzNeYghA4D/4Pi8oPo
hyINQDlTWAvLudTcpHmr3fE6e3oH/cMDpsfAw5Skeyyok5DwoZMFoCGsESHI
Ok12yz7xZptz4H5+jfYCt3gRzoJ0zLbRTMc29RKSzno0CgxE8VocgJ3Fzy6z
0h0GrokJcmmz+6OGI04bdhBlB6cjlSm90tOaBuxsltaKRAvWlvUD+Dv0vLss
Kcdx8GUEB5QXESx2w0TqZDxEON1opbYSNNm9qV54aX22rAuBEJ2tfZgUSLCk
PLaXJsbA3ptCF1Zpbzkhl0htE1HaGFNiAeiS9zOHwc2o3dZbtdM1xk6Itz6A
dpAJTyuC3r0Z8O0FIRBQx5TqLH03N4kx7nnnkegjh5BWLRlB1WNlQS7UX+gt
zHV9Q7/KcdC4Nk0STAwjsHxkZ02dDyaEGyfMfrO0Uf8TYTVlpYaBBZWW3MJ6
JadnWUGyraFnzraVbB8UeODeQI6JFLkrGMWFagBr/ztyyGpzIvLVxlIAdWzh
HiaRwXWcSfxY2O1Vg9wuLUR+usr98UNd4DYZdWl9vAZBF0aiu2+MRQbGExB2
ZVytfBwCBRShcAoP0p3Pl2bBzAGicTclT6AJRFVHTTPk7QC563/s49GX4t3c
PIT/UiNPbKf8AD7Z94BM1YawNStWDE5mbL6feK8+CLfMSUndy7SYbb6dF/bG
D3uwxSxHOhvqeqcMFWgtUrHESVBaVti3cMJl9fI01EepgEp2PzGyNvqXYGJD
rXy/WAn2Ue0GwZkcEfFClc22WPMCAGQ7YPTofTgT0bAo/MVUNxLDMQ2Fq/kb
Ro+b0hB8CXzzrIrrflo1PHMznqPn9iEsJ0TPs6ZrMFaoFpbnpkCaguVeeA3V
UCsYpi86qFtoYrrWBW7h1i/Si+ERTVal86d15Eo0/g2TdBd8trW/amqml7Ff
yCYIZyTE/NF+XbGQmPiTT2VOR/udGE8/owPLT/pw2XhyYvQwz1cK+JwMUShl
RRJ2YfMSEZJu4fRNeaykRfq6m+8TTjEGWWsAyqdqsn+TMtjE4fioQhAe58Lf
Orn5HDi3BqLGBD/VvAkJ/ma3mdtrBelqPmVo6GT01cccsrbJAgP3hB+Y6RW/
YAuKpk5dla2wxHjIUhng1mHzT0dIPLzRdnX20U9Yj5Wz8X5ggKBGgmelzDs3
2Kf7p1I73qdaNjnzjeJI4s2ttN2QbppUzkfLxI6Dgv0z0gTe3DT2KqFvZmxn
zXR7estuKk/oTxRr+Ktzhu0D6SNqhu8q2heI9uUW1czqL5bl2J3JgyoW56KA
pJ68UiH63ueawNauJmAgrvjtQ2HSz2EaZnQ+d8PJquA0GHGRrYLP52gobL2o
tzlScxgQsY1QB/SibjMvL0dHypp5qtE4j/u+wPc3TGsRWiYkiTLiVxM9h1VJ
+JvtlWOC6d02ZsEcQVQ4jbcRXHhlJT/2W5pYa52xYNFUqpJwPWkG1bueBv+R
MEyQExR52+Fe6bdRSl8XuLcT/ErK8thbKnmUm8n26mLHLHj28QX5LqltZm0h
LQHPjU7TVOM9HiihRhHSogtFC4Ws/ZYAt/VZo4OlYFEp92lTKDUV0m09c2q9
h0Go9z5SYARKR6qJWeIsmCk9Oiomhu4z6cssUo6h2unaUvthdIPU2cEhNNtq
uSuE/Zt+NV4tLK28xNDbKe/z5KxGUgBpbN0l7N8Gu9rheX2sjizHEx/wqfvh
+KbsnhuKjxhjVjcTkUsTu1kSCNyQv1fUFNMiWMeE6sJoLW23YkMDLuot3xve
ailKFLW1ZKsc20BXDeYyRfx4gEqJf80tfW0snN0OQw4Z5ZggR40kW6luK/ZF
ExkLciU9+3DB0pjuy/2oC5wbIFWcYgH9EArNySi58mvYTJYheuZWpf2yjVd/
jLyvi4232O/vNnN6RxBcMzjl7N6SHtp/SXfijJA4CbaAaUlunzhzEC6hhu0F
C+nI2cbMN13uSsjPtQrvA5TCQIw+c3PrHBM09B7TjgP9bMWh2kNkRr4BL6Jg
FLVyh39pXcpHNR28SoXgHCoJUfMFTaQQZWs8pXVyEvbWWb4JGlqNF8kTf16r
Fj/yL7WljJXHK68aQlXrtI1ddNx5LC3Tz+EOb4M9wnLAGn3PxFcAuKY+y/GU
5l8DGCxxKpnsA+3j6rlFhuU8sAeGvaixheWfkBAVnVliXPv4VgPhi9dKfxhV
P7x2oKyNKxbCPzbLSM0I54+hKBQxLy2G5BuuEYNWT4fdvBtRu3VhQMyEYcU/
CwD1PqTtEitAJ5LKyCpS/J+L1bWk+xEbJyDGk+phaONRQnoY5HsuM7EhL96x
Xs2VPTdM7SMNSXfdeLIvKFn7avIX9PE9AEqH94cOYxmWPuqoy3Id/CVmUgd4
906MhbeyMp69f08/xSXFpUTE07vxDgXdcLZ1irNKEe3Lwk3dsByP2gYtbXQ8
gHtcY27L20fcZ19KJhMSnSBQP9LdXB2yh4yAKyZMWfdC/W+ArgowVR0i5udz
FrCuj6t5R9sMeK0CCvBrCCGQvU0D9h4S0JPnPi4wx437Icxbdw5Ian98Q7qH
hH5Mt/msrDRTPePboaC9G86liIzy84e6/UKLRrxkVHJVYFdOc2sqodrUcUFY
NBbxfxFs/aYtLcWDXkrtO554ThTb+7xG16zcysOhixQXnUeAO31IWrhFNfPS
GLPFbazMgPicHkrjdsVk8eMdgu3s97Yd8Fm4jwwQVNXXT8pjL7KmC5Vj6FhF
BqvxOhv7UKvNkldNpEfM9Qv9iSFJ0eeSDczcT2keiXk9jOToB5fmJckDTN1g
tlrtv5i7gXZRixy07VEKI0g/6F17k3zSWcLLVUZsIO2LT5VkFboB6g/aUr8/
fNsVYFqTLnszMZwepegQK+AlX7LX0Og0kXXaeHr43DfGAu1VyVMh3DpBkc4F
b1rX0T7rlZs+glCstH17rQrjD0vufR2thw0R9VIZYcbq+Widhd0fEy4pRFcC
Zos03hxNnp6EPAzFUyNQ5Ycmw86f7LBN/dIJFab3akclYHJeqbQDYlLf/Liv
0GvNflxrB/fF5FqtC/FiZF5TjfW+aErPGASkK3b3J9hbjsyCjE2Ek5ROxPWx
EQ5N7kan1SBnLHtJECqaXy/gVGRLAOgi9RYJWEDpMOfi/aWlKjajcCIxO/dW
PBhS4usLVhbo5+SJtM7oWfq1+tevK8obMd4NB3Cq+Lk9NUqzdRtSP1hfXtK6
Y1axIsVbhKNSJNjFlo8GSN9vUJcNBFNh5Iq4ObvTqHR4ADolGLKtsgj362oH
NkoWs9VLKttSMooL/5Zb8peZXr+FiMu3mbGYdaRV8RywKGwcX1gLTPZ/ZTgA
W6yBPn88n8zrKm+p0hUcEOHflCQQqQMCDWEUoXnzsAicG23NZ40QA4j1lMam
7No2nwEWxQEcCEYzvCRSdHoSerwIQlIvGhQRJ/zqj/p4L2qZYpADXd807QAL
yW16qZOJHaG+3diZ8cvtLR3FsQzEHxMXEcfhVpl0pIyqoF2qZxYnSrquhCrc
5oOhbcTQOkXvgPJ1/FasPQUOy+POddoQ0/3t1gsA0a13M+2d61Huo/KYfwCo
Y8L/8lAgs9LpVfVIizIz36u2o9zH/JCCS4HaEHbKODS0UT1ShSpLnbObkq7Z
R61kuMEsiTadhyed5whKlDLiyLZhiQJEm9rtOQsilR87u36y/GTyVLjWkbgy
hzBL8xotrCKOISgiwo32jJSsP2Z3/hTMaMtKQp4+GHXoY9+c3yQ5N6BAthye
pWP9xKZlUVmWsRf/eWWk/AumRwgQLoIOVF3DFynKFnIVJyD1QhB8VGzHdYvT
Z8Mzjw0ep53GZcLtddNrNA0EaMlZfMT+j/+NGncO+P0vCf29gqZ+yM7pjc1K
NQ1u/Ljedq7CvumJoqmI1ierLfYZVVt6u6NlisLm8b48HOMuhuJJPjIwfr4n
+C6MtIIcEEL6AcfNRFGcSgc2IvYmM49v7ebJJxqTWLEpg7lfuGGqGmSvWC8o
Oc4PTeCK79SrvZvE89JpbPk992BX5lzITRGV/wPfnGN6IPNx4S99euZxiUAh
hwO0VvtN53svbv3L35SkKuG3bofsFpkVBk+C02PBZ6vXSBsJ13n58T6QZYy8
TANkUpsqBqoVop+SzCZbzUayNLR1sStDLY54/C+m/Z5FlN7RTvnqv57Av7b4
qsMp3otEnjZkr7l+ZBUMLFibe+GPLW6Wm52B8+TSXv1ilkKMOKpxpgFjkLMn
v6Rv1JktK/cskKULZB56G87IxJYDLw0OuaH2CbiWw4pvRnZvXEMNJYJ1f5vX
4CvqAtQ//j9YaZ3JwchtC0/lATo3utm2ub43T2UxeS4Sy/Mqk6EuiPRtgzo+
+j60ZeugFu09z678M3Yql2WhUOCJRUoidVXVEdWeJi4RwLnLx+p0J2LP8SWP
Me/Fx7/6MyIdWbLnzFrWHo0MwD0WahcKqGqtU6oSd7Ey0G3EKAJbiXllUwcn
MWA6aB1T2J8iBw1YrQUpV7l38FjyPSwSXVCBbou6NcB/lXGaNSk/robqFGY2
OMzE7GKI+WOfaYiGlglDF00ieuYka5xOzemRAfnQxgPaIWWfkB1/PInjfL/x
JI1ugg01HR601mhzJl+/fNwr9iLxl24J0qXVZX4oFHMeg1V+QHdaZGx2fHJ2
AExAoE6XJDRlotKP4bOmLb2EdlGJ7KZHflwXJsQYyjYmtq5B0gE6ObkCErmS
6TQPeaAzdP9Qn/84wrfhpkHj4IZttOozkrzLf+hw5z1H/N+a+1YEsmbEubiE
bGbr+m4jInMzvqS/51dSIPnSZQ1RhitdIGkuXM68QnIITrACY1ONZenmqFSA
bwZo5LLdqIUHdqhqqkNRC7rxOM1oLwJZRrVSkhFf9LEPwRpQBQR5oaZpZ7QT
oRnW0hc1D6qzEBFQw5sv8xvNd8s/5lZFelKndbeCo9MId4xdkgbQN79ytNu2
LLdjFq/o2ybIpu5hqMXpenviwsOry6St4S57cAZ2pyEs4f+K1ncYElA+e3OM
1nUa3hWXVnoQbTVH2kQU1hcVyvAzVyzYFYYICFC1zN1aR2KIkY7/v9iyjoCY
qDi6xz8qGcaJwrU2KfEB3O3V8hdMGC7ExK4rtYAILTj6zrfyEHFpxgcMKnqQ
XpzwhG18tcwWcre9L0UWNZHgqZlPi92snZ49Ww17AeGFP9+/Yflmi+aNjFG8
htQSa96Jz/6PjkADw3OiwO31ACEII6JQxyfjkB9njmKazXQlO+dCougy6rxE
WQsFcfh7hXhKxH8QaPQAMUwoqkWy4FuLGMSR057p/3YGo1xUfYqHzFqWn5f6
rhjKk89vPTjv4GjuuxQjJO+obnABctK6ggXNA6gKPSRES1IiducrfEW5wJ/f
JC5x3dLa0hn+Tklonmi2PAnI3Eqg6ucVTwmIEjHyUzQGmy2XVBQXBFMJuaOa
7WMb3QGBOXSx4oldLmnynyeqfoLK4xcREpgK7tftk/KeOr4GnrCXA8iy+9ZX
jlepFLkF/AvWXpfluS8A0X3FRFhJEg5SDaKty6pVCmReT/JSFgZXYadq/oma
oWmzk5JRmRzsKBXmMAfhQxrJzN/rHy2GPJrb12yaQhZmIybnJx7DKAO+LKTl
zuPVlF1W1sTyatoFQptHZi9isYu9FT1aNZrGzq3DGI5xZVWsWG4cBAm6qD7X
yEpfXUBJCdhAT98wp3G6np2XO++kGuSaibBPZwyEDCJCtgHLqqKyOzWEpaEs
Gbpv9WfQ752Qf0fcq+KdDaddYGrekVbTFi9CgUtYqZJgHu+8PQ3ZFPqkW0EY
zzYHVLrfQ9HzIXNwNtkYj5jXSWfKOwULsjTu383qc/doKqRI18BdBnIXSSE3
wjxm14aahkVqd38GSLIsSysdzwiSBD1qh2A7O7ePtUjNLoLctZJ+CS7wB9KJ
fDQKcxdtiqsNv1C6CbUvgWtJxZmiEj6LhlpB6AZ/pL2qQWN9f1EI9cIuNjTB
BA3UWNnEVpv/SfE8IehAcoun9BzPCR8CRQbqR2mDweCV4mCfZKjF3ukvpaqP
A0+9tbdbEB5hL7rYs72VeNW0SlV+u+HX/Kg6a5ORmZqp4ds9T1W9QJc4eiD4
0GpMIdMF1DBf5acOlTflLJqtU87FG6ib5rw4GU6yC91+TdS61WVYuPFJ257A
tXwreturWjyllX0pJ/gj6Q+xYiiR8BR3slXYuMB7WQ9WxsnN1J6ULTGb1Dcy
DApgKZls0l4TMBvGpRH4l8gVPMripYlEFjn0aK2sdAAQJEQlvYrn1UIMic33
bF9L8R40lHrNoIwwjsMmfyyzNj1icRS0RVaEkxZ1gOxmiUIwHSeTFCdECZoY
G3P6T60e8HeB5lBM7GsKZwhDUFwU/eZyQW1MtauofuN++lagoM+4E+0cb4zb
1TcTwjgzhyKLVFxVI+bB1c4ZOWfzMwLimhzCouH1XAQHhNl9bxzS/mOgSp8u
Yo30mSob9b8X66P7k+Vj/TXiMYTESeSAINkwuyAK426Ag5CZtCA13MdKOe5o
VvG7H5aJPY34aNmI4yfv/uYqVPIIHvPUbtucFEqI+2eIcmFldJp7cucAhIcV
417sbbbjF/rshhGM+sPfsEi8XCkXqIcTZrpKO3Kvt4PrJ+eTsVrP4LOLeQi4
38vAQWsHAFwAxcK0fq7vKQmv6/RGccn4THQB7IbTyvcEvwtpOWLLRYkB3lVc
4VS21QJQtXNekPGldZhTwiTBeMzYgWz3N/ikJyG7YEL/+b8U7E9FbjNgHnfX
/Kdih1jxBXchm2LrQP26FDf0HeMooBpxqcDquD5I2hg9x8zbJZNoB5Unxpym
3IrgF4EbUwV7Da6nTWaB1dQY0ywflAoGAagB+5hEf0uOb6tuQdEJ1rEr1b2t
OQ/XlGE2Yx89E7sZmqRuSriw+xM9JAPKWDCRb3mW6yQLaD5KmXTnsXLxrqO/
tOoXxnN8Q3Ex6gEDK2uuiAJfn4ENo94DBpl7nE7Z+bDe1Bu2OcCbdhJOBmPY
/pErp70S0E5Q1ML0P8TL0v/jGz11aQjv1TWjOhzePVSZW50LPGc/cmAFFICs
AVH+yUck0hFjzhzAGKVdWYJFa++Nnzg62M3FF26xVft7pH9XGCTVWXgsGA3T
MXGv7D2glM7SmtIy8t8axxALJKVhIHHkjI6aMbz5XOa9c8uJJrbunNTSMTMl
jVDhOMpooRhOYzL/3ETxZs74M0mi069UWJ3sdHk7QzpV43Zw0ROh3HfV2Z+k
ky29mFSamLsCzybXci1rrDM34Yr5AOCUQdPz4CdsFaGMPfRpKWwavoagFLuN
SyEYzs7aO1TTQh5wAmvLmJGy+PIa1Hv9Q6MmK6RTteG/QENSK3C72K2JpNxu
+sjvXoOrn6LSHISqgVdfEEv3Qh2MXrNIDAanrBRY6VMUgrM5cYF3BxUeQwt/
3uB7GF38dkDcieVukAHb5fpmi7fCLCWR0H1CnDAYEpHn6MxfPjVsllZlDA66
7S9PgzxTo0D5I3eXuVncwq3uX101/trLslJe5rHZwxP4YrXM9UCiZ1oZuoaz
5N3rNGb9Ph4C8l2tsITQRw0QJkpmEheUAGeH5yw1qAbS4UPUyUWSenT/jWTy
gL3xAX5VBOUd6qRY/Txxk5Yl+gKvqRccLk/ESuby1RvtPk4jLv/EVo7trIaV
CtpPQwhhARN45mKvh8joEsvIKhdsERhx9Ble6JzhyP25KMiKw9uhpoGfjV0L
SqNgqudIeB9gaK5Rjd+Sjk0LMehaH3PyP56LW8c1KpWgQcLbKywAjRkUGoq6
+/wxR945RQTLHNjRH8BbkYd/ha7YehvmfUcVmVQzmiWRrfgElAegTDprMIXE
cqRautcv7QgprLT3z5wVPbBPtvUhwHou14IXm1mf6rGs5WgJiYOzkP8g4Dbx
TTU2d4EhJya96ACTIIL+u83H1RqugG07vTfJ7AW4AK284w7msb2/har9Puse
BJGMzkwDgg1Z8vYcUOVZ6AvJMwESfKZ4MBhIJ8EXw7DqqzrinxCEJPOzJLSZ
mGhJeQ95It069bKej3A8JtnqYPHRvbUGYMy70y0m1SSNpHkag7DpqyxA3DnP
0vRleyPhGNChp/PLP0nlV1qJlshDfHWEH/UH+5J/ol8T53OQGtknrENYtFyQ
6hVrIrg05oLqZ/49WqDe3LqBfYF6lr7XJ66Bwz9Z9SMvkecSwnZtyY/l9WMG
dcNVSuv7MsRtKOVPzF6w4ULrbmlMe0U9BZKBSuw4+9OyXggwyRhZD6kvYuoP
KfsGJbBi6araQgDvHYc53zfHjt/rTfhtSnbjRczgXQoVyUyIw5VN1evIdIHM
8kltoUVQd6cgCZc2godp6JHfyoWpSVbhlB0n7A6kxQcVMKsBfqkA9/KoJhDm
yaUQDm4UsUoUuItucjQf7sAZMfBw3vAYL2GKUQTzrA7soLztpMpzVlFdOziv
nakTL9qpTB6rH4n6Xkjh80o06LMva+RDGp/oYBr0PiXRGrB3h6EBLHO7jPxQ
7ksfrM7qQRtoWcw3Hzn0bOqQz9MBmoXp3gbYLPact0/xCla/EX3x8ZGuvof/
pr5yYYgXGrRmSfu39Bo/nyXj2hC7I/b1FAx09an/zwhfiNcrP9JSQmkaR2Nq
krIDHPVD5g6spAtq4c+ButvozcoCo+LH+/tFyjjq0uUkO89fI8k0K2w4swCj
QLQzl0vpX5thAWDmZ+kJNGvUQieSX1N6S1KR0A8vTc2hlierTcEcA2kp84qr
fRNtMs9Wio/PFvztTjeLZBVF3GId6mcs7hXhUz7YZwQNQ7pceXO5AXlLImgK
ddNXob7B2uhjSN5exKP6VJJZ9Jffzgcoc/3jfMwIccLbY/rIypFa2Ug5i2xj
sDb8AsLLH4biyBwfedBQWJPkpJo2LsTwc5Zw0ivB83iD/91lMvXaWvfYxd6z
VInMNO6VviRa97QZ5mYTchspxIBuTkLGELEj1R25UCxO/gmt3YcJqsYOwRhM
VuIqe/itCZpplO700+ijlI8HdKuJktA7XGm1LXbmymVX3ps6CmskSSAljGm5
97JTICiVA86bcXOPrWlrM/Z0eBYWOy9G00Ac5IShd5DPPKlpReYfCouZW+mW
DTzhg66FFkZyx7hFSx5yK8WaXcJffThsrPuY0kMJvV+J+kxOcDrai03xNuNR
XmBYNJgT5xah8a+EBiUcnws9CPjE8PzgOmiTC/z1anfiKct1zc4I/qhj+Uor
pn4c3ZQcd98ffGsiWQqdTBGbmaWwyZTpu3U89UXoFmEiyDDjFc4OPniTrmYG
T5rDXqpQA3InwNijKikYyZVYAEbZGA/CjDrPqaRM+OdVsvB5TfxIN1mFUgI0
XE3KJKBvBsSNTCUgWb9uqLdMpCFDV/jMgjzIaA+e+UePsHS2P4/j83GvphRX
mGVNm9q/unZR0/TtlV5m0etlSZDEy5PMBkYd5CRRsmp46I8XxfsamCVy1l7E
GDYj5qgBgXZdSsMMG2PvHBqdR51hhVKziboJTQ1EYF58Hay4uA5QloZ6bd4o
iuovJBETzEf8xEcJvLkc1GrsAXChFxBRj+NJzMIO0cqplTH8VpmnAOGNatq9
GWGE1YA97KTMmPF1RVqPjQcZ3Wxl2Rw12OuIHyVA5l0YTLNPm4vdkz6q0gdR
5nwkfwdrMCFBXp5xVrbe3OZeOeVa4ObKWpeD1xhONNkEMFTsH6JBM5AtAHe+
CbWjxMVSnm36A5PwHNnl+sXOKCKyfpvBFPD3WJkVaUUM8Kz34qs6lbN5JUSC
3dFuBM2k8oC4tQkxN71w6Gmpk73UOj94Td213suOp9zppdVhdfIbcsvqWKwU
IjD+9xf9angB20KZ7KdYSwowlyZSi8/pcDjhEQUUQKnfqhHyA/gM8P47J1EG
eFI8xWhIOtDsGNwMPd+EVDM+G93HA33Bh8E9gI+3dj0rzepVOPLOECGET7Od
e5+4uQn5VUgXBwrxrJn92KYQ9a6wH9dJhQzOT96GEKtLqFf5bh/IXVrgE9Mn
gnCdBX0T5WZ6ruHWLiElLkh/9YGJyTunZ4fzHxj1oAFKKH/eIqXpztzXrUla
AWLQLrS3Ge/sBZMAMo0LxAV+03vmoT/ORP0TOE4PoFJS/wCbZn62nOt/ZNFE
1xhG0IijyOyQNhrnfwMo8O6QH+PKpDUFpJrqjMAL8mulV+yDGu1Fz4wy9fhD
wJS3uej/PmEsnxWON9/3TV2kSgkwWqsboEEVNjYUz+1ldC3wJC3WZE2kBvzm
fULo3vlsSc2iYewwUiL2+1AmIujzGamINHcsDEMdFNhGHGGJ1rrs8coEnzwH
/g5EdnXNfPQg9pgJaQPDralBJSNyW6Ai/AaVOjpzLQkPMn42tHyQTQ0MJggq
bxqcWBJOgHIMbroGzQ68OTr/tGeutUkJ2aCwBAdrjDoxwdHwFnhL63gkUKt4
F8nqwma8J7P3oQmBVNJSVLYRZj/6NX8J1B5DAmFgRABsmsEN7cVfUOyeBW1b
CrwrvVHnLnkkv0+EoHQ7Zj1rFg4wQVCHlz8tnLNacjdBh9IK4fhLw8K1I3f3
pbIQ2GoNPZyejjROPzeEsCCkNSn0g1luimlY79IZDpqwxlMAGTQovqQutTuk
ZOUg2G3ya+d3YAjc5V3aF80989JJWE2N9ZxvL+4KpzJ3KqZsM9dqRWc0Ruz6
APuxmN/CufhIooeMBZn61a604jmQ00IBPRBNVLrtVKDnGJ27C6CUMs7v9JRh
N6rOW7OWdBoqPfvp1uKQXvkgPJFthHUo50cRHLRwXMomoullEClW1pX57GZi
9uK0ssX2FCMHDI1K2IVTLGSvJdLqiTa5IRdy12tM6wFl8FCgTEtVWCqT8c6V
/RR5D16oZwD40L0JB3Fl4o/6jeiM5N20Yhk/q1kUV72TRMMo69gXKHl2v7pD
fGWaSOtMKeJRgfiENfLtuwSnzwta4P6/82HCaI7Dd3WdJvzWv3eM/OaTuS0W
MvywJY/x0IUDBdFnIEU2hmXimHbLXTSKMy0BYRI0JVkJCxyhUi9tlgsuE3m/
c73Ma6DJ34Q4kbNV04oVYAjOOkrbjnDQ9OFi2J5f1Y36ucj9Gfkj2tSLPeJC
UXM9gKz5XlB82+Sjk5+2vM/L+yO2Cdssa9oeHTL2VloIDx0/kDCEwiEnxtyP
zveHJ15oZFxYxCKaWhl4FskRYfR+csY1yb4WLDSf0qbZGvANLDjztlQ3qB6f
8yiC1sDLvhqakQy5NQFo1rNOgKQLnYRzFT4wUu5UbUlpH8Z+pSv5XxfQMW1A
vvxwUN0scsWwqPevkUYR5jK/OdAkz8lDjiqCwroCvK/dlfXlY6cV3qzvoutF
8PC3B0W76b6oDv9Sg8k4+0p7TqMq5wM69PCubx9lvCliiRuU0xBSjksIcRM8
8uokecewWUUZRXQHjpDS23xG25pF3TlkF47KrtlYTOYgujL7hQynxI7blEiB
+mwAmPBNLffLRzVIByvJtYrln/W8ZhtgdIhJ0kubIU1diFb74cs1m5uBS9rc
sC5v+Eqpn52ovN/rB+x2uFQDQMwBBBiFUTQFnVIffkH0XRPXywiJEXWkAZS0
7oXp7zwpxlYaAhntDsAXTTrVkE6UHlyzVXFZW4nVUrBSgtoPaqgbgoAhh0c6
p9I0I6b1Xce1d8GEWmqeDqhq1NtZXH3mtTrAbZfXRV0YBoalKdJIRk1WRuh7
IuD2A/n4dLaTymSLY9nR/C63+x17tHPDe1gCxDrwUwKic4nirDzLBDAKQPyW
X6NUXcr4xMNG4XlryQ3+7Y9HpPTYR4oXA6eJZAXbzVJL55AqeED4ky6OSvpr
8Iu/vOj1SvC+dsR8eaApnS/g4n7AUXQ7LqNbob/fIVwID1I5nRFEhMmiioLv
TNgA1HPQ0C0qnv7AOy+8clECq6bzc+Ev5uLgr45qNpGLuXyXHkk8+HnIq9AG
qdYe4OfM7hKRLzvW+VCbRvrnDwo9OcfJ76xafVzeJ6LACkPZ5nguXNUE6zu5
2+TRAwyY0X7lnSpzAQzOX0VNy+G7lC9On6/XOZfwNlmODWr78JIHxOjmMlDY
8BQIJF1+vLKDERfQ+fUhQsn9Jkhk5cf4Md90QubE7sBgiaXD/V18Ipiv8lCm
12ruq8A78jvjjvgrGnvkaHSIXJ9lJ/U1hlloQ9LHV+Vu+siZ1qypru/brKYw
JUqoafBBDuunDKFPZYmmfbcMnbCzMtBmosZRfR9GTKHkuXT22NeJIufEi68G
Ab/zXNucfRqtRCliNhOkAlPokkG3XSB92KllD0VZKfsWk0S1B29Haa183Mw4
QiW4WHT4gGhH7vJaGUU/W2rfEAyaK/1shdQJDZJtvayZaUmPSsHmH1miZT0R
yedM0KzWhNsPwFBg6po9gHUgqkCcOLZ/QZBzGfaEeFR7gEAUiWJ+xACE3VJk
N3cONFIE2hjcgedymibqAL0d6u+5JZ6lN8ASsGQBasHp8uVORgfV6NHCCaL4
VSD3nsHgDTR6Lj6Vc2fPGLVS95CHEAsfTbmtOBBJKtO5YLZ14UBodKqYZPuR
AxdGkoaLAOQyFU+0Z0RysHtiQqcu08jJq+Co1n7Z8A5OlFXu5YfQGNsah/Yq
oSg7Cy4oBB8T0bNE3lF3GC1S8lGuxzNF7wos70YyPmgW5bESoPiwVQ1f6kXd
M4EwT2M+I8yEPZ+3Q66SKFhC7wrN/a3CseNIU6v5BpnxHa5IP/4ebbHdCCVb
CbIGoBc07DT/7D3sE1kmD7yc7UUc+RwiU5ECTNZFmDywLf1pur0tHn78cIUc
+mkIeACAxyjpuCByTbnYHiB5ip/bhnOzcIxzXHLGHc0eGL5bL8zAyKQ7mgcC
P+YtI37+Av8AeMQqFmz/CSM98eD0Ik8P+sP2c9yrzT5Z437qzfrBGDnHUZbu
mtmPO+Ijavh8uenEnGEHNgFhf1G7GdifkBHLLglOCb/hsxgGvruGQSPKj3aV
5CKLDQ1cZ6+/y6MupH2Fer+XGz+GYKl6/zr0dGXVGmyzPL5P4XIWdZL2J5xM
cuGmXu5dzV3gmZpFzASFD5CHfb+Wl8KZX3L3uvgVVvezIupsOB9kI7LZtK6/
taZkxqPGBSrBknvGRFSaQIsSWBugAZbL43SsBkKp0x4eDeMPDsRDooPFpVJy
NfcLnAXAWpY0LhOYNMB56wiwdOVLwjcxm3ud8C6ZnlVAPRiIrP+xsM5zUqQq
jGPvrCsvH7v8InDWKb5Jetj+y0q3qxiNhgXMnGzvHRphGvq3757hvtqwZU6u
+3PU+gzI2RJ7nWFujI5EdwfUkPQCp+DGDdJ+wBzwFQEhJqcZ+W6se3ldUaC0
YcEgx9QMmtECEb+Ro/7nzzANQbX5Qbnb4RAP7rdnWmvK4Q7gqjcSRSXWqt8M
eythZGXN7cIHXpYbu8m4X7Xo7ADpSmsXOG9XccOvaNmr8jfne7Hvo7HYBmf/
kwyyLqAJFNRX/b12fNFXp0ghbis1EO4cgiAlYiK8Aq8ua3JEju7i5NNbAsSS
cEyk7jpsCTU8Afu57W39R0+W0Gdv9TcExBMZo3b7Z7jScS5GT50Jhajy18iC
ugidIToLnoxyvcz4r9afHDw0X4NUlsF11krjAkwTRjBp35+rcgQwJRYJTi7Z
vCdcMJtHMxoPrEtNdkTJaDQHOWgvESdQH1GmXCPkGYHmy/PU+N8tTVnvcHtK
0pn9LjW7KXQSoCUgOKIfqPAhRGl6bYOkg8LvXP0S6bqFVWJ6BgD6FLyzYaxt
ks9ERw5OVCJx6A0rSk4W/PFUES+HzTZ0JNfZ+xAphhjjUQwtrkAL1rmwFu/+
NrJALIi9tzRPCK5ZpsOqfv1OFlRTGQAqWljG2ZadQLNn657nqK5g/YO3RJSD
gai4n8S0dHKugtxn1y06c+9hEFfPhU5PeVZ/XilCjGt6fhx7hg8aeqz/PvZL
vO6Fpy+q5KXVKv98OFdLSXBjsvhx9OpAiEmC7bBNIruE9lTnGVW6azA30j0d
FZRjNuGYu9R8wEMgWuiK21di/NLc6GtR4W3EYQxVt9INqf8VA0sIF4tdGP+B
MuAMIOBfSXnvdbKcUft9Vo/IrIjxEOLhk1wznG3NC54mg5ioEA3DKzJmOuwl
NCnCBCKenOgN0V1hefPkWbasrxUCLYsJPD323xXTntpZjW4D8kDV75qx4xkS
TP6iHMMEp4JsMNhO9HliLvCbOKLo9qkhzalPjDmCA9gYc07hCF9+93xhcrUC
6ULKH7qLYFHBszjjAcy+CEBj7pvdPdgbIDud6oyKEQedLHIzxD+a/bv5zaog
kksTQVJR74bARpVYCOBjicTQ5j3O6JJHVQGnBA4KU1FAMSu6cE+SpirVmFCR
qnV6qdkAy37w9RApS3QvbnlwMC0W+w9Y4Y06OzNMF0FoTWlVVikmGq11m+CM
sAtAvVGIvsjpR6/hAd67OwDhsUZ2WuHa8J8gPMaANwrGXD4pLo814SH9wBal
1qWDSL109vXITlW65DqpQyB2U7k5JVUefUuhLNNFcyViy2nFqD9byXXUhv19
VAYCyb1LTpNOJHZWMJ/9n8hw6qcnqc+hEtOLj2ut9k2EPvAzZKhXL4vythNX
rnmqiwXrDzCWBAQhOtMuw7+Ax+tgDpLWdCTxmQ4TjL0/8VNKbueaKY7YFUBg
oUcNk6LrM6qTPsRIPuqxxyLgOsPkcBEIKrsuoHC3fxYcUsAS7IcBla7ITszt
IrCoDEGWD4ktICM+Dbebuv0dvQ8RPodcuPAqZ/U6LPxY2gzFRb3Sk+pZRVEY
IlySjqY5h1KhEfNUt9hn1OgdFB46M+hooHBWSGFlMXjQnVfr0uUtsWVAi0zw
KUDrfM1v0tWy20Fdcz9a33QDpr7Irpkb0IcOISeXIQkmXPmb3+Yh

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6CFQ0q6dj0+vxNyYPd7wIa4yDYouM0ewlOAiLygL3BeHxBeH84inBq0OTn4uzWCLyeczUO17tTr76KhW/m8a6gswVr/mJfUHgVFBIPKzn16Y5Ff9ejng0hDsom1W87ceP1haTJ/6lE9uDiCQOSuPRXy6HLlXQDowP7oHF4EJ1D3iTu3mLtD3OxC/SqJzGZnoL/L0SUm+WLc0eSNRgLVxhQZ/BIv2rZ4TPV1biwCG5C9EtNzXX6cpg2My5CAvERYrtxrJWbVP/4gtsgV6RZ9nqlAs+s2tMrkYhwDw6JA75wUyEgnhaRjZUmMjU8Do/oxIHlBF/6DOiQoEij61zElOSh0ueaboouaw8kobd8Enw+etslMLwaH5NuctkXOW43fXL2uRBrt2Mq+XES5yiTngvCPuXDqQB2pLT3j8ib7dr0vGWzf46VGD/zByMdZDGTRZLt6zy/mTWiU9cLLfuv2cBfocik83byxt+1cWhycpVhMhgEwbqcTPUucKrMyDxC8JQXwUYRwtbLbaEYPO99Dkr/R9+u34aNa+8bDTa2grep9a3kx1BUB73G1LOV0Mz9gH016ERcasocCO8mbcfwfnoTRiMQEUNRuHmu/AHBPrRt4k/0jshMddUqCf/xHWvrUQaV4onJlbdIfh6jIQCxyez/D8UHJWLofYv3kPkE20OCfrv3a/TypEcoLJQhe7Rd9xfLFCR7rCWGZI8Jwg/b/ePkXMM547440q4g1pybwCYkfHgC3EPjFiRD37Bzr3LNTi74c6077kTVhmGIjLsHqhKjI"
`endif