// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MVu+2Te8AyF9dHhjHesMc2JowdsF33tCQZBR7KPYu27JJHh6/drcfUVq5m0c
pfc35zHwCjGnyFexx7dCKLR8Jse864gC48MZ4PSEogGdMDe7dB4TkTy4GD9i
WAnGgNMbze5cHLsp18KyyUzuG4MuQBaL0zFfROFUJDCH5/xjCgpsCS872VMw
bCh0NvfB+elDY1pobSjlC3pg1flYL25wovVrVF4r1rv62Ms1zpmVOth49tY/
MV/B0lzw2RZ81JqjyUAbgzo8v7UbwolUHS1YNzCJah2SE9yUcE/T4HujDsga
E5RbPWf4Ke5E/x0q0z1LjFpYkJk534kRMQswEDdsAQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JB/EZhTO3UUwies1uwteSV2sIkv/bOdcLfrIPzMQf5+VsIzECLGhmTkefBvN
RtOax3cGEhOvLbdEHntJpSTm1a+RH/XNjvlVZrkfQl/4U4DUi/gcQVnpi5Gb
V1u3IU039Xfm10I9tre1FVAPLVHAY2VtLEjeBo/W+dFwPKyFmV0nmtrNwOlC
ZuglqQ4PMwka+PRbQeRn5vFUlxejsc1Ab5boYAZg1M/nKxDJddzhjAN6P6Y1
WnzZolARPmyzipbz5P2Hq0IJJculaGbOKO4u3emrKM4zs20rO2dqMVlj1Hlo
67KGUbDv9ECHuW+uR7eWNiFv8UjqQRiBJKetpB9a7A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qq1VL8kR7fQgQtzw5QwDsKAGRVdbDCp6Et5/yvVMzwprSGSzb6poB56NcX6r
Y6etFYnQoqby9Cz4eN0L2Q0H/nnNFrQIVEiAVDGbyvhO1b7xq8ecmZ0LL3iH
ZtlmB1kdYE/lVRicUA6zUa0LJiSjSqV4Xw+UN1zBkZDpUVpirPFILdfy/uIH
i5OUf15wCewtuRkNzX1FpRFVyDo5WO8jgTkmCF/Y7TxxB/j53C18fnS7HYnQ
ltkPjYHcWbucaQf5o0txsnu0g4u7qOOhCdznIP6jiSrjVLFLSZ4Vyfl3IwuD
I7THPWk2W5CukEPEBYCKrjI8SEB+2+fVsrvqf1eRpw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mwm5U5Kyinzm8nbYbAMGGgO/sSllhmRd0fg099ypmJEpjPN8Z1O1AiWnyuWf
Bzq3Kg/arAElot5fuo57rp6Pp6luIXq+z50xM/qBUv/CXXLMv2CYcV7tjejd
zSrdMmOoFIS0txxabBbPQTncPgy4oEr7AhcKQ+4LFhZxJ5+dzxuaQGK7884W
dZy0RZ8VS9e8F2RX37qp903N3M6dka/87Llad0KtlZrA0x0M4000elMBG6Xq
k4lYeVRtS5QyDr8uhoZ3E7etV0O54n5XDVJoZVxl8SXL24mEeyd0U6yWPGB3
b55wgYOWBDD2YVtEwT9q9y2nDgDOnhX7qs5XMvsjOA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MeaBb0NjBoTdCNXIYIktmgyqBvm5B4NHpDQxidU6XQ3P7gNKFC2wG3GnhyMr
nJOKTUky0PUCQTLooP2zEWnuTyGa78V0Kgoz+GYfF7x3ODZrdtu39+I2P9wv
A69Y4FK7AiJRVcs3rdOM++jWRpqOQ3jn771oqsKA8/por6eDi+E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CyohXmN+rIjYUozgJLdcSzwWfojHgqAi4JYe8Xeo+juKzALFZQM4nazd1VLu
U1PVHTG7QdYRZrXDZP8Y9dejdu/tZ7ziIrNZP0nUYa0Ojhgzi+I483fkBVH0
AEsnD8SKL06yEDawv1NqoRMRBDm+GjrAvhdybm9DOZwCqU7l1D5YOocbHOhW
RfjvJMrR6MscrDHFBrVnzCbuCWK5swvHj/lYXImZa0QZexUA/OD5I2l5gLZ6
t4Hnq73zodKJxn3qXd8jD2VMl8HUmUOzrOyvi+lfwfVdGhjRR3pY8jtZXl4K
IMcNItLOynVxxeW2mWp5zxUS2CSNFdhDqxoR6Opi8wHR0QCMm2Fn8w+qiZsC
25Ai6501pzp1sch8YiuwtSjhUCA57bGCT7nNlicxA1Ck9MGYtvJWHzCTZmDv
V39sIjMdYCPhsYiFxu9hfrsEIemOJC5RWhsvBNmRgexp/2O6zRSbC16BFB6u
hEqXFAjie6gZL4gxcd7B5aFNkmoZvLyk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BWaM8Lu8yKtFD09qaoCmdJ7eiDiJCmDI0S5jryzl8XshfQndQyhKcuuhr2ng
hji42phCoKupGIW2frRGOhrYwqQw8KkEG9lEd9vy6hL16zidsxaFHqs3CIAA
e3F+NzUB7FH3gbsIk5js7ga0l35dirDQSsh4Z4FIz2wgFNwXp80=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LQFduALNwt2PuYp1j/i4E6PfqHcyWAJIK+4QVhKze1ofaDA/m7FGbmf+Vt7w
Ie2dJBIxH08kt+gkrFzXI9Ma8R/K8UD/nxzwWrQXBk8m0OrZrOLSznDU77+S
UGz8S5JwygC+kD1qxzOdDAv0RUt5tvK73TETY3QFzttE09iYa2k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 24096)
`pragma protect data_block
uvGwH+AKJnpG6ahbMbL2rFk136f6+yoH3/ADeOb/xvO9w4YrbdSULqZ+T8I6
i3mBPnoLRtJ6xrU/5l5IpVpI1/8o/vA7cbcUxH/q389fcpVQKzUM3PtBGKze
sHZ/NQywsop46ExM6nsY+c/UiL0cYqwKYt+MyNs9a6edVxp3c4vG+wcQ1wrW
tTVszQibcuOd1e3T9i0MlTiDXm/iyZ4npPG4ecEgSMyX8WMoZku6cv+qz8qu
Iw4rSdaycuwkVHXM4yyvTng1WdZrtHxf0zxM78Si0h8GuP+rOr5Y5ULcPgOc
yYHUDLgm9haqr49tpDD1nUMsJzLaFsdH/aEBIbA+84aGV6rjFbTxbvRZNYDf
rJj2inLWaMWgYKYn5WLw46/fJkNLlWriICVPFYCMuOlsfd0xma9O6yI7sI8/
PIDZJSBeyd6J2ra2Zk4hajFQCIwTs4SG5+kiQFIa1pp5WC0Fb2JM5Z8hicIi
IkdKgg1WMxddWlmSMAUhVsuZKKpq7vtpCS97mfNrLM7uKW3A8rLHREFtx1UN
yvWCOJB6pcf7VbhPdijrH0o0aRSztk/I/hYWHDjo6MaIoeFtABEB6bob2Tza
w52nkYEqocMTVuichGX5WCrIw6im9F0Gk5Y1LTRG1hAiL9XCAIZ67r5bl/Pj
5iKoqR8cKPRhjKavMKbHvoZaToBY9rBdERoDV5pI/BUqAl6fMVodxfaxR/Vr
jAt/kDK8U8BG2Zi0Wt7j4x+YU8k71xJnXu5nKVh2Eo728cfFArwXFjpdz8Kf
PV2siX0ETJbLq7IvZYrZmIW2D9886jkLyyIDkHtSNjPSU+s2DX5DP9NWYglA
Mc/cne4X4XMxPcKgOO0zLkC84sybHgaDXZIYY5bSGDf14VhrzEO5jS9qX8bP
3wq0DUQW/3VOtfmVBUFc1Xm/WX7OrVgdMKolePqOinGcvPeWMvjfDloLxk4d
e2Fmk8brV2H7U7pQb2+YG8ug4IS47r1rkKUl8nLSwhHH9+sEafUewgB16Eql
pG5asLrQgLP5Dx6K2ojbEckCtXUMyf9vIdQ8ZdiNEENcDvYwZ8P0bmQwXaeT
Tsc1iIdw8q3x8LeE5hg/EZay4iPOLWRxcqEyboQy1wdd1hGccNoPHtwdGR6i
uW+Y9zz2FDxmxw2Bi98vitbeqSOQjNRnasFa842E4d7qHJfb3iSiAcNAgLCs
dCzeiMBpqcIs0l9VYsfQWJhSD33clG1nN6DGo82IFz1EX93g24oR9gBtuD3C
D2sUkzMfthVHamLKrr9W0iDDvdbKHwVhxBipIr5rAR3jUEr4K54+yVeME49l
uBexlMp4WBypjepUzfSIHLij+oOuxIgerslWOeOeaFEBE9T5GpqHxgEGO4ep
fhJj50yxa9qAvMtaqMv1XoBBlYuQJnyUA7lm5P/i3coteoj4PbSrOfvYRJWO
tvBEwHKJcWlaHwwhCqsQUXXCSYdd2fTAGFno+UWyAUWuisIfwA2llB0m8kCV
J3dbLGwnWCsCqxmxeRxq2g083K6RorWE/iF2hM+uiI3XXzjDEEdPJCdzbMbR
PFaFdY82SwVaN4CLVzzW7ja0T+Jnvi0CER/wgZ6CddVOO1PI8O/u7/97CFdt
EuP4Po1L3j65v8kgDkr7HDoQxv3BV0hehMEAHGKmgJZ055RC0PmD1IqQQ9I7
SChfNH0iQPNaSvOi4g6pVuACizKCylVQoDJK/BnFsKz3BppJYy7AhdUkKSUj
0HBEOsY73xHuhrwzEVhyV6RfzuZ0lrTePb3DkuXVEc/Cv+/lUk0C7ld0U+fC
rPvGCjC8FYJSl3MM/10h/zOdetlUlEgjPuScdWdKETre2J1UnGIWBBlL28In
mA0WB4EWWRmRqiCIMs682qTLGtNONCflcEUP3Jz4rlpJVZVoP3779HEVVNsg
j02pKTTa/6p5GEyMgL8p1BfaBHxnHOWg28gm+Yr7mnku86G1uEgrFGAgg65y
fDPCoJwpqgdCqYMous7OLU8aM+r9SbWpFvhCXjTEynlu9qKDsC9toVf7MmUu
pGuMtb8KBAaKJERxr1hZ+sCMHTTWWKJUg7OaGRXDl2u1D71s/RnwxhyG27/j
i8WAoVesgr9prJ4e2LJmOwuZdf05xx1DMB48qrvFuoU34SGcp6tqtUTnkjAc
dm+IQltKHEtq7FT1gBj90jvXMdVc2UzIr/qQWc4AOr6LPP6Q0pmoKhm1f7E0
GXEA6R7gDzlSJKjyehpebX27qXNIEq2YND8i+WvaWw1icduJYDYjZ7jbQ/Dv
EEV/hugCTViEBcIeBImvCQGTN0fM3/cmCT0AnSsoUiTA5aDO6XBQNVUqV9eB
BH/GzPY4vcwUiL0yChka7bvfEBVI+tPKqFyY5Ze/uuN6hQ8fAm9jdC2ZP3ZY
AUTXEInQu7QaB+1928RX6g+ZZ2YW/vYeIBwulu8EyUiujIT6H1ZU1p0lao4+
YfvHftYK7LD4yFue4YCjWMqV/ggbFzTn5Ogjuph8hSk54qi3i28zD/Hpm/Kn
3JlTdVVT4gm0RTRUwCakn9ez5foq6nJye1Kmda4UWMXxBHUAxBKl1fXo3xOq
vZ363jGrDsspOqQWm09yo3R0MezZSvdZgurWzCr05LnXGAzo5XkDBNWIMUGs
0ucOPikM4dxGRZ0uc/Px2404ku+rQ7e33hBmt/YssQEbBdAHZcyoH5GBVzDM
0pG7WzT5yLisdYERE35hsLDJkAH6L7HPuPdNvJhA+TfCcsUBhJuHNY94/OAM
4bckIpL/XuGhs89e9y342Zf7RjpOfkHJz9ec2xZ3t8X26N/qQr/M5v8lfT4M
2jOGJpy7nINg47xZGeJSTFxvkFmyuO0Yk7dgCEsedVUmWcPt8e/uO8llyoRG
uejY9xoebD6GxGeUAha4TPJupAe2zoUFNruwIsB3ULjLKxKeQJoPmWwE74lt
yo7PiKnBQI87cUkdwt80vKAXiKiIoF93pIX4to17xMdFmsu25Zb+iHJdjiyg
JMbP3Wx2Fn3E3XLT4KZq2miHIug4N8PISFzrAYDvWrZ+iUSe53XiSuWyf0/M
qxkUkE5e/BudrzSdvQ3zYDcCpizneHCI0oZKCar+N3+lAPCn4SzxT2vZjrtu
E6H5v8HtLKGz+MOyqSz1aSreAJFzHxtZjQxAprMs6pznRn8zLfjqkKl/gTTj
+hdry4NfOAwUIjtCDInDcceO/V5GH2pRrfeIAB5hj9EQIr9V4XLmQGRVTKBp
XeMDEiKv8WtynQ1ZO1LBY0adKjIxvWq3l4cpCwmGAcAOOLZYAg/5aiop+RWn
G2Dk9Z1k/+3deyeDL/BG+J5wkjBTECfeFOIYGR5YYETNMwBZcxWDfXqdIWxK
eonm09AOO4xsgHJhWcBCJWuktKrNh1oWzhloS9Pr9IudJ6saAYl1f5c3oGrQ
JKeM9Ek352EVJnu0xzqu33eICI0gIIfjUp0ZmdMXYD+vIy59xPzLuGod4D7h
Tx4HPvoEDG6FS7jpAW3UFUmhgQRpTe2Z4lEytyG5yfbvnJYSX/sssVVinNtT
0hEAqwHWlvZfUfVvYOGVwf+yLfZf/OJmTAZyw6aDGZ2Gs2uiFElbUxOVkU1g
6YMyK+Yv36DFfhwhCbLGlNvI1RAWVS5DWTpOR7Q8/zPBsdR2avMrcjnHjYJc
ACYwSYFVKJ/ocjNiZecQaf3LJLvRkz+xlpssFKtmJSDww8ByjftU4HEZ6P0P
o2yTyynA1L2CPxmXneIKtoqFKKY+voWDXWuRxLDmBWme7aGDUueDb5IAaKC1
gWw963S/gqc3VCw6Q8Z1L323v7KGj/zdk+WGlthsUG29eMH+y5/C2wA/deIG
Yb2n53rngTjOsiDTluWYjgy4ShUlSW0rOBQ7sZGkispX/PlNBameHJY0/yc3
NsCIAeKtxIzsWmA61aANjKtXEO29vr9mwEsbG4a75psnhpeypfE8UDxCcoS1
v4lD9I2l+HZw6xv34GN8EmTdI1Yd6RONkxKYhO/mITllpdYZ0/wiyNGbKP1O
w1tPBmCSO8UFfnvqhl4aMsuv3hH/DD8HVDTf0mGpxkGD43KgR1eFknbQ8SlA
yeV+7fzd3SPPJVGb951fbsft+JarxFQBviq5pVSBI/KsJ2qt/jzjJOREbf7S
4IW3HZtr7cmPhUW0jWyLxraJwYAOGaJCCS7uZ3y11Iqik67wwfHmTEwk6rj8
flt0jf4e5uqpq0i8bUElJRo/HjYFDrrLShYhjBoFUqsOGF1Hbu5+mICheoJB
E7vEJz4nw71THxEg1M0ZVQBkZDGQEqWBdCEAvSHK7OGmqXvILDGGtUMRsuKb
zaGHtGkcGLKfH84xo0g600gpIBeGn74POEnQFAuZD8hic3m6u/cepOp7k2Y2
s2baUEHHsdJg6oAPuIrqkTRQijdaX3HpxtY0YgM0eDH0aRG8qi8YRLu3h4QO
na0Ip3zJ8LznPIEpLFHCbK0wr78dRZm2m3y7HB35o4kSQOYAB3nUUPnHuz7b
t72HAVvS7isfslwsb1NR6eofoRBcM+ZpjOs4vVrCMk81Gpk4wE0KKG1WAv8Z
leFLpNNRz6Q4OPbWXmdCST1C/JVvjQTeNkzb8TMUjQQTz9bR//sz8DAOuQlI
rJkjUgJ3X3f4zaAV+VusBwubP6sXlMaLpttymX/QyQQDYNwpwst8SgPQFvqV
KXHlGpQzXNBUGmKCyPiwX04hdJqTf8sGDmlXg+GuW0C51oFmoiJQcoJcVX19
8ooUg9X9dTAUs+aoJXsDw+C0gsmguA1t9sevllekSV5/ztBL/L4/WeJKmma3
rVbjdKuKqaSWa7ATIAc1s24q9rTyCeiC5gBMrPeFJl4ULpwMyWU1I4s7kOYy
KNNmzoEblMkgf/xeN9wU12fvevGxksJSxixvqGfmxyBPjMh3eS9tCab4pdwQ
9P0aWOIwfVRUCOGAbmw4GP8o5Q8mWadmoZlke+yXXYG5RD4UJDE8QGPUn2cw
YkXJ2+tBmcYz90wqXgeUDYwD/JdyIABAf+PDaHbF9dvRbhEBe6ezec48idBx
Nq1yRbk4Gf6AEqID2QmQGVcmm3R89jRNAfP2O63Aytnm25867Lir5Ld/50lq
TSd8P6RxzYIo+UD7tog1wvVbP0qHBF1AmWgtZn8Q7Z9ntUREZRO6Nc8AXHCq
GbH3LEYiRNrK3NXj7yMYpnoDwHGkMJ/iHljNWMUtdKJZXvNEWb+vAWTxhz2A
kxW/T5w002v3DL3uDwxNcJp//yw6TU8is6pYxz87GTNNc4JaC7QQweXoBggH
o5/he21sycdfaY3UfFEAMf8MFi6kHLlBAwCL+b7LVtBokZM4Amj/zcH+AKPx
zQKIVrmPKw4opFqsPxRtAdTJBzDADfccWwMerO5nmVjejO6Lq9DRp3IZiRPn
0Kp9ZR0gdNjdhCPh4UuqNFZw+9OjnFxleVi0l6WNDNixIGwPVwOFmdJs/zZ1
Olr4vigd505Iv0mnVAcBlYZfdrsdgXO/LwB8bCLD4XhT5Z1x2Q4WLBCNW39K
0mfCgumQsIlLLsqIZmUoeKXaIFkgy7YvEwtDPrpRSWChXAEJxdoG63QZ+MR/
BCy/cRbKl6FA/lUg7aQhCSUjaantIYO0j8xXUQBOC72ziH6OEjq1akPNvA9U
N1qC1KFlw58davL7AOz21rlMgSFjZnTy8x3we10YyA9sIHn7iELLWdPy4u0n
nsGIntgZ99wPpxATFPkmd/TPPNeM4fzGqZ+xfuTWuwIXFRbWkYf3dpA5J6w8
ynUirT6gjHeq/ukthK4Gnx8HiDNXLGiB99r1DR7PPuhC/jrI1q7T2UrXzbN9
Hwi2obvPZOQhztc8rurJtdNtrqRZ97Vj36r9+4nefF8IcdKYq1bsQlbdRboO
CzuHSk+SfMkIAkfIumOda/zbapfPyJKuUfUpNU4UGNpVbPiGaeRIy44nFoiA
pn6s2qecfJdydkIGdm47BYSOXyoSJAR9C6LAqOAJw7Vu7lot19j4ykgTFTB9
FludhcVZZvpKWL2cMolQdvLiioXFYe8mYy7gUE61Dw6zqPBlhRgYjZvJGBQz
OikjAStXGoi2Egn2lZ4Jgip1Ib79y3Sz/0Ile2P2l2joOzQ/9RQWcThJ7v6f
Kv1ATN98/mFYPqtWDnRaBPDIZme1KRIOnUms+HCl9tSON84TG8beLeXgk5/l
f9LAWuCIJq3Is7xvp/u7rM7RZ6iIhirzNhpyHHLGfRkQiAPIQ1jhLWd8KhMU
7KBnRV7xiP+cNn5H6+leIyGAqSMciHmSvYt4z5eOy7RF3RJUpXEiCu9OvnqO
WC3W4PcZG5ERHgRhl/WESdB+33iY6CyA8tGP+CbjxItaeWs3bl1WjLh+jlSd
1bQMjKgnbVikyA4Xq2sFZBEs4OSbPHlVm6r17fCW2gZhneptVAYiCZlmljTZ
YrF7SiAkhuecD92wn/FXGNV1TJj9IrzmvI2+lYx8I5De1MK+gTksTUiQw/Vd
ECzsSljv8vq0p4QmAZFqtkLUpS4+pjiivImk27ZQ9S9aqnlWcILTSlYWQUIe
yG5zSPi7Crb7ycAX+lU2cqWbia/R4/tVEO3rz2fmUmpvcZL1biM9eFxoDyae
5pZc/CrcsHwxdCwKlqoCdvIs8XfiMYrIvGHDx5jZeIC5z82t3L+sqVCpATio
If1/bCniPLAeh4JMfGjXkJh68a4ccyUdRbZLurv0jpB8uPSgKPMlt846zGaQ
+Lz2stb7LRYtg+4SSbB92Rj4D/bcaq0QULMrHB+DP4iqrKfUPu0kJHHrPtXx
/8usNABroC46omTptPUmX6BS7SuqYMjnIhmFW/g29VurA0cqPznnZbb1BQ82
pMsiKCc/zqb6KIjXkE9F9hXb6Csvq6a9DQ56iQ340ZGRsSGQQYJ6QUnek7Wl
hv/BV0A8bZ8LoSXp5AxgVIRGnPuvxPFQpYg4ShYB0eSN812eimOdMdbrmTK4
5wDbydhka62olz7WvSaOhqNaY812gsX9DPw2YkXuuW9WRsI+9uHGeyLjqMT8
kis7lPkC8RXLg0AG9V+07OV35IohYRGG0cMMnpTSqgfesLB4x1aqrvjLn+Yi
RlGmYR/9WFV8aLbS/OcnYTvdnGy7Uh8+eVQdVJPhEtIdsldfy3A9kzdyq23i
U+1uAEFc/YttFJyGD3T4f5zOggvZXNzVC+xT834jEhAjf/QIP1KxJTxA3dZr
N/8TMLd2Nb+qQ6iuQy0LHPY44hFYUcc9yNukLjG1fsnThJRwg5OdZhoRWP62
f3U1R+OCzV3WlKbHAX+2qoLkUSrf9XW3eCSNZaeBv+iF85g28PCGqpe5rJZn
TaykIR+Ck0er2nFfNVpyZTCPeD+Ane5XafZhDYv65IE8UTthGIlU5dC3FqVs
fK3dJip0UCfEEkDINhIxrEOPT6DfK6qMzUNO30OS93q/JcC5Y9GH6TjtQGda
G2x62AkJxNxFcSqtf84/Ju80RZelCvGaATn1wmaTqcY6JRezl48N/jvHbdlv
K1Gx4j9Lyg9ZlAeMz4+F+koAycOoUdR3OshXtBuK0ZD+6opG3NGEE5fY06lT
loupxRRFkzKogEyiCUXATbwh6s+hDn/HCngNWDfhDur3IFoaJBjJsr7BZr3/
cOwK5AVA4FXqKv4UW+G+KYTvbbW8s7LuPXyxFHAxG3xsbWKRfPapvyCS8uDw
F4oPBWce5Uqp2WeVUCM0rEZMWrUgkW7JZ57ef4BK2npwJ1MYnCJhmYjcVQvP
hR4dDT4N3LBkV/niKuiyj0hCPfkhYLngPExCobW+eFygB6dlsGV5WAG9WkCG
7kx2TKPjGPvhsn/0R3LLFPtcSZ+06ejHKBTmm61AQdYWFyPurJwS/RCDpN/1
qjPq0aSly5n5yiEpCF4P/fk4s4SY/C+3ywrhYR+nt00/6i749jxdD47bUVNs
Gxit9RzgBY8GbxLdVQWnS0J5hRk0ef324ji+8QxjKf7Y7CGZeQMu6Ou3Hdgh
S3LJ6PKpRQak068oTuFJteEe4p5cMnjveXrLur3vHY1aII3u5VF57Ufo+r7Y
uVv0a0gV+lAGXHx1Fn0qSWPlRl5rA1QJ3VpLg+fWZ/DTE5ajpkBpuSlDsmd6
+Shfa/IFiHJA9NHLR4btkJ3ibZLkmqPlboUlX7GVHJG2gz6XNZefBRZc/M2Y
ImPcWqYPK0rGRAWsUH9wNTmFr4tJk8tCKG5NJFS9bA2rhH2rBjJybttPT9mb
W23B1VdnexD1qgdqH6ollnzNKJ4ms8qL5VL7dFdWI0CAww7+FOLNXJyDCczs
TIOwDVyU+36dU5+QtATfIsdizB+Uh5PvIkr+zBw2Fcvje25a/osZDcu6XPLf
t1wOQRBjY0ChJmPUnlHGZ7O+95LmlilVa6ok0aX4XX3RouPklUWj6FjosAwf
KvSTINURxobjkLTlEDpOqKyzWvXx9Q8qQRvumesH7upez2zwBWZGCKpvkjYp
puLHJkoEtA5Q2qU/u1DxaxvT1niaL72KAp8oNtlU2nY+s5QkAZp6Gu0KDiaf
y83D5dqAHYCZ2ooPAlVL1vrICxWX6rNbXFHTh+6EW43AntC1xfLQBxObKZ4i
sgrpGw+zKJYGvUsjyYb3myLuy1446sZYOTO6TkWKNOGYCOh98qla7LH5dUa2
stbzerHn/clagrz6y8gEptAPXqi5akEW4rfJ4iP+eS2AioWmdxKrACvvIArG
tDwR369RymOigZ8f8rgHALtVteaXDCQnQhYVs9aHHvDQMka+JuEhL/Xq6EYx
bD62GNOoGpIexJzpI4J/NH/ztcmk/sHVU9A0UXs4sCEZHhm4pZyVuBuU4daO
Jleunf61OiobVcO73/rOCRJu6cjZKEPCmZrAq7GUGGZCpQYR17+XMQqvMJo9
YsUAfbOKJpJVQ/EVaJa0oqZ1ns7vn8L3NBW6ZlpdhlH81s6AD6Wi5d1H1uD5
S8BhS27PrY1v0FDno7Ue8pWfgTcRH1dKxbBYP0VkVAF28lGJpKzkuRpY0PJ9
exSbODjpyFipPLSJFZDamaMxjUTbXCKi+M6VrbR0THlwWU6KPALB8+jL2VpF
lYYJTpJ3EH2ubvPycwTopx7isthdtEVlAPzs8a38lT1jy3ge8o+9AKNAQ9n5
POw2Mb9ff68kAEMmt/S4CFSvJYPLxu9S2Q3QhLtOVEXDCANRor52kvGnU3Yo
M9b89z3HoyzxGwKzaCnB4eAENUr8VLx1D0b3eExPX9B78G1y+J5xdJTPHRiA
eY1HeWnruivD+4IsTXkBdT7fCuExrO1dlsBrknL5VZBa6x7SpnVDP/1gJ4af
0SzfWaQlYbGr5x8uUnxgPcN8LiYOIi3zEIutkQhhGAGmvd+qeH2T5/VpJusQ
Gt6hEWy/q1h8lggdfim4NR69M9WIuyqKdmCjxA1ymVLccdMSoPHqG2EAIc5I
OOkKFL95YejxJMGqdz0JWbHmuyjBLT/Ea2DYifJ47NXxvuZ6ISj/f22dml0i
tA5jbHL84aEJ335oVRCXTHHEc6/tWMHYBtBCJMXU7GLhrvzLDISmSaehjB5g
d+Uw46oUcXKF0a0E8W5k0oSjRB0G04F0JVJhnRweTN6g8YfFKp8ZjPnIkWDD
c5qXENrJRueu9sMXEjmMdzxEfWa2EmN0tkNBXb2unaRMQNhmTlnol6tGvWj0
nSbydQ7VRN/sTm8hNCqMVlXX2+a8gyDA9oB+axZgn5i3BzVp6WWw24NlbdjQ
3EiVkW2RflJ44UOlvtrKe/gbnb4Tdm1irVnTPi/mnhEXF+2xnkKkCo63aZeo
iM7B6quA3EL7r7CcQYENdvayvLCJ7BkAM6hxs7Bvt/1jIKqmyufrja2EtDwV
i+xGcKtCpe8EMwZNMonK2orVxkWDMVFh+yeHyH6QxDhanvP1u7nQaTOkWJiM
qiNxf7wkpAInnk0mEMNhfKW3xnoZoqxmI3Zfq5WlQ7diFPUQclP4vsWWKWjK
a2saETd1kZA55PQ7TkS9vyAgtavRX4CMIRxqxKykUA7cuZKkc1Kvz9CoeIhO
hCvfJdejj1aGYbMntAoYeKlDz0k72KT4L1Wd9utXLasxNwy1eiLNVUMzkpQ/
CYXKcH3ghtPfJo8WYB8L9X/X3+DArftpmka9BYbaH3dyBcJ6K8ilVk7rXYfm
2SvJ6HZQfpKfxl2ALlrjVQ3wzzoFmi7jN52hQi8fou1LVdAa+Ht5Cg8D1ifU
lx/rZU8XrWXgoQRZ6bigQGc5Kv81ZGmgF/h+00IpW2kE3mrv/fV2MLEf8rN8
gWHEIZHpGVTzbDoYz2ddvXaYHF9eL+IKWFcsMyvMmekUdHDnHgaikVHj6Tdp
rnpR4q1dk9HlWW8ZTbspqzwYPEfbXtfLgihRdDzeCQfm9iiP8C2OxZ0B0gkP
/78EsNFQ+8z30WeN49snzwLDBwyXxGzmeXYwKn2Q9dtPc/en1CRBcIeoPLJG
Ywa2ZeTikBar8TqXxdez3yqA/TFd9CXN7KRX1feRl1fCJBxNO87uvsZazqQ0
h1m60HrEnDEFO+ErwCGX7WhuYE/+a14bDkUQp7x6RKC9s4iguqGIUJkdRQHe
fWks5vNl7ZOEPLL0iwXSa3l+lawP+x3SOQKxcA8XrtXpIdOZS6DsXUYmmMLm
K/6LpSlNjSwy2ByUBl06Z+OVB2q0bA0GZK1B/Za3vIXy6zq6GqtwIowmajem
Dy5mcrjSaz9+Ynft5zAMWwFdd2VlFGU9+U3/G4rRuRC7iksN23NdYUOLtBSh
l5gm/WBam6s9TB1sgtTWqZ2XZzHU5kedI8Ix3CuHTkHBRHeVHHiV6/lzfmDm
48vPiITvm11Fq6hmihtItGJ0qFjytlbAny86kEO543SogmQuofpNKfpZOJdx
XbeuDkIJbnFXqeYHIr0xaOCd97MsM+YaZCEoyEjz47Dj578Ol5MjgvjC9Zxp
9W31lF9LLz1Fma3DZ9znvio4DN4KZYrXmA4cmaUjxn5ywNiVcDcFFA8OqG2p
z6HPil8zKI1a4P/DBiIXxaKTUbmqzXprFbCfxVrxNvLFkos8VhzI48R/vF2m
W6TIP0w2skL8KLKjjJd1pJUSmNtWKgo/iI1xMYf6wwKhS/kxrEv8kSEBdiGM
e3dhlSKYAWi3ElqEXitzahHPTragksARP0I1MMl+62Edt9r/32EiVopgO71L
flFxlTRlq3x8NY4CJNrarrsG3RH95Octc4C5WqZg76U8+dE6P3SsNSmPjWGg
pAWwl6beCboGVhHytA5JfKb6pgCoOxR/rt0kz34KNBRixazpYUZHN3Q6gu3Q
s4w0sv2SyJdaXJ217zfG0ChHi7ALoJ4I+thUx+WMpBsDmIjLQZSSsjMetY6/
n5rgoiB0aLeMKZTAPI54Gidf8GPsMEohKlh3udptKVnVcjKJKmQ3f8Wb8JJv
ttCy/Y0N6Q5BBS9/IK3RR62/2I1lEHDIhpOfV0f8sJrgTvpLtXznTyhBxl1g
P8VVLGgc5nR4/qlMhpL13QEf07Tzz4bR4rr7S3Ggm2zrVGlbZyFhV9hwRotW
GkxEdC/gz8u2V0F4GmYIpFMvmF8ilKmL/381PczDJ8FNvwQr/qFYu6MfttMd
4GyEQeuRjzDFmnRZwX/s5ePnb1XJqPhw5H8+KK9vcDIBdjl4ZCUj9o9AN5iZ
g38mRKXd0KHRGVeThYEAPSalCBu6Z/HoAswH5uyKtErwJEqhndDxFuqSDcG+
BehSU5wDTyyDgHgvkOIO0oewNo7ZJGMludOE9CQLRV12fxnY9coKD/o4vGx5
vDdH5WeDs5P/kH/4zDV9ocPgMqxy9IAHxGCRZ0nlGKMbWXmu399SWMnBWpP3
EplbXGgGIXMGAZD5uCCc0wltORfTJREenmGEo2OEWfHbf6x0bQKdQKZqyvb0
X0KyyRL2WMFGXDFlLYhpKfw3rQKv9UbELsMr0MrlkpkQHwuGvjF0tJYDqTgr
DeZsy2HtNMO9C157seFseQmxNshcLAPwStD/rHGyIFzzhxZ6WAmpLkKpDIdd
qXAiqROIOuNb4Afwv7JR1tBOokHL331E0SFcIpba4jmNrnNbUsTvxJ+0zWic
3Zth/RnnBNE1n961h7DiaRzKGv5Je/9QRvbcz9HaEIXyNPzu3g+7uh96ehTJ
A9eQ8ZMbskQ47bQfud1vnWPQRW1MA3Wv+IjNPXQ6y7kCRDYKXIvsKJvyqVWx
R6MlLU0OpadXy2vpUgAdDoPvZ9C7CmmlNd4stoMEf+OModc0Gv/MFi17EjBB
Iw4gWGBEGh1wWQHeuX4Y3+ma1I6KQMqMZNz4MSfdwkpoWvrPYLtUGI8oLxHJ
DzfTIMXwfA3KS2/Hswcwe+mHV5+gIoMXQdglrsletdD8THyASk4RhHSryD/c
1gx0cdwCK0xQmfk+CX842sQOqx8vPtDQxs2Io836SgQTnS4zh6onpQWf+WGF
kJey6SMa+hTf3vVkExu/ixx82JLWMFUpBRl3MNjH+LXLyD91VGwYI1EHJfQX
0+Mdl2SGrU2Zts3zGmospmiP3D3rw15utDKgLzQptKRc9PJRCGIQ42K5UWjd
yiyV6t+6EesVxQzhSgEHeN/dAC18HJETMt172HzA4wT3YbJOf+vyWkadvWGp
7tdKvDWp4sfDbOXQ3+qrB/kf+SaSoFFHnCGyTkotCDDI7eAuibPPqe2/0swQ
bjVsoet27wM/owRpgbv60bbzjOMYdk3a30NfEl6VW7l3YCY8Anrkh5BG16Y5
KN7FOwAWapv6f+/p9HtlpTolF7TkAZ3ZQAwF/XjT0nLgfZLe9AxrLOCWplCP
1DB6ZvL5zjn0JU5BTwA7bTFZdVZuY6cg2DO9lWgAcNK/luwRadMmZxJz69Xz
0en5d0oLf/nzYTmHxOfEeKbTTPxnSUJd+TRiYb2WUqpBvGJkgR2xbZGbgcOJ
W73i8Ke6FU4h+GlM+hkMLtuViBKY8NSOPCv9c3gkaOMCkyK3NMPq+g9jvMnj
eUKtrtNRxIfTstmyNRHOaJLPA4CqEjMtqbZ/wqfQFBZneHXVrnuH0B3j4YLL
WxabjaOobY3sn++zNooFZQXWMbCEQRpVilhzPUuMMShFxDZgOlyyZqxtEE1q
7FamNJHp6N10bdfhURtutPrrw16DjBdwHqC5SFAPtOcZkHh9kuGsQ7MvW6gL
O8nqB3EP377DH/n19Wt4Lj3a6UdlwIy8ztjiyoAwX6IeCd8ZBDutND8YqMx6
SahCSq9EGv4UmJEhFsFyDv+0+U503IEkHI9nbxZq4TaXmLpNOWI/R77t2nP9
AEtShgTp+NDRjvCWiD0pCHx5Bk4inubz8byAboXpxHzvAgz/o/NzqSt1hw9b
pAQ4sVVWTWJ5Ns+KgSLOQBy8Nphiq0tbPlhmWQ22cJEqtkw/7TAiQNWNPNms
pxWQjLr8glmbjKCG1kwpNYdlebQEvcOLrOuUYuT7gWw0bV9T6dercwtQrLec
XaGk9ZA151D3YSB9v6eUjiZdkZFFOaCg5RdLOYSYPEsGBgWiFd0xcQJZRgtL
91jWbTpj3cZEQCdpYu3ly9JJAmx359xqShOycvVbAoEgPF01aQ6UUrGKjWdY
/y+icS/Xgk9iGRloGA02qQCDtHB/TlXr4gtI0EbUZuh8QUYMk3tJ3cJzcvdP
ILG3SZ9rYCNEtcQNbyX/KhGZAQ1AMfUDDsQgXhpSiyWCFWp62mo+x8rsx5o8
Si6cKdcnkX4qcetndtM3ktrWd7okeLaWvdnI5d3q8bErNt/mk9On63meh1yL
cHkNDJAA9tpwylFRi30SUW1Te7dLVZe1YATVjRwVOXrH1QNtPWRzZgQxWFT9
dMf1rnCii0/SOjAvW5vs5uEo9jtlHrx1IEbz6YbvHyzqmvLR427qIhhUgZRZ
F1AfFJ3V8rBqJPN26xCB0uGeJLgbHz1gtSLef81gSKMxLnVMdY9QLcEeVETe
gxbLk6j8xtkdm2MS7utyCi+EBnpn8Pu+Iwz4gWTdEL8wkeo2guz1iN5tIbD6
dih8O0uSuLC6LgMgQG2/SaB/K/5/tSIUz1t8Iepb1V9w/WLApKiVtBntnHUU
/M00EXS93IDmNfl29LWwuPD1M64B6aV0NBxZZxCySz7v+qiTEpdv/zKbpsIi
J1JYKY8Un3oumRAHKip2Y5ev/sEMn1Jm5o70Qlyv/Ml6nmGfpnSV2AYnFRuS
8KefGTNInybUb3TLkFx/OO/90h9YJIADoTFNh7Lc0QFxu0Mh6XvZnAECZova
7xj+Cow2l+YcdwmjK/ArqELePLonzk9hzhvp3Ima/d14ckpHDM+SnOdBlx0N
3eVAV+m9vzk6E600zqYatxGo9B/9CFlps8cXvBD0SgYFLEo3sdM8MukOase+
iI25NuWOzieSQESgiitDvsf6I1MWUb3noMbMZRCNb7uzD9KqkesT3Ou7NTOr
EADCSKTdh+VvhP/Ao9qIpMdH9S0aTwQgltKkpHkXGJKDIJP3qts1ZwgFdmPo
qg1H1S+SJsb4+axOSd0ykYyC2Rehu/PsyV1RQjIiGQkkRkeXHM4YTzEWCKhE
qKOAra/X4H2OPP02BJ0BFE0X02EcC2NAv9F+jPBPTABdDF5aYXHaZgibU3qw
K0BG9QjdYl61K1eu/5HhH8YNCD7/dQyAc51qHLqRsnyzoc6sHCaGsN1/mjuw
B0bS7bKVavKORyJ0Ze5bxDfTCn7Gq4Y1Dz0RSgB8TtjaFPEFH02HTr7wJtlQ
5OPMF4BV/Jjh06/fq5GDyIXIPpPFRKlvY3qojrMBezbq7fSJeXIfVPqdHvJA
gmnYntUhsZNK/NC7+IZJOIbiRnVHz6KafSFusDXLXa04VuRn//RIrfvJO9d5
6cHXjXiJR7P/RRNf8GIfSUNMtnG2z6oP/qt3kQIRsAPmontQn6VF66wPF4do
ioecuSoKVEves4BfJFM5uVHjwiej9bTNES9Yg6VMCRiQW1y9Vmy6ruOPXUrW
uqsI0Wd9nRYhCMRVVnyzKj3G/0HlD2UFBLDeXDEHiuLrnWTChE53MCKISfZx
5BECwgiUq4r5zS5GBytUp19MveSn2uzw+RTTR/TNA4VCOOeVOQExR9LVcy5Z
pTp55thiqXzkCSBuRAHlBoZRpPSafD8ITAf2UMHSwGyn9ADhPoVBNj8Czn9Y
sZ96kFw9JTBMTzDdPB9BhaEdgsgqeuX1WytTrL1XFp2pi5jjMkJL9MuSdT5y
5izhx8uI8lboBoW1c5dfvGIMeYaCwObuvMaMP2gcBAOElMUx2KifaafWGaZC
xUiTGr2tRtVo0Nka3UFTC4Co2kmvgjnbP+rm01n2BY0FFILRItocwQx6dQxf
0VCs4TBJ8S0ME1dtdsx2aj2HzuTRwTyAlXGSoKbLrI+viQTstkruS4aXhKIu
yF9bJ56T10N8SFFx4tVEVQaFYf4kVeSUhIqf/f7CMCOXu4fdUoq9bKsl2HzQ
/I2fDZ0WZtMWLbIhNqt2UOtOOpEcQNH4lXIyAfU6gW22cEERjKTXtjfA5IVj
MmpnrSAUR+qBz7Z+r3iz4P5W86GhRcuJ/kCf7x5qWCdcofSmumYJxjfoAwHN
yT2pEWxWawTz+NDMcLBIqx2SBsr77oBBrvHVQkuYP7hA/tlGuobF4V+NQ1l9
ZYNpW0KfU59LV9mNQ+gvwMQnolsmEuR4WMlXj5jMDKYu0xd13Bw6aUFQAunp
P7pxTcxR12zaEBl4XRZmQKE7B2zhcnCePKIp25TRFJQUTcfxjRM/bB+eCMFK
A6yyhvyCq859oQDv1iRZkJ9ED7xGYyn60x9N4Xkze5AICkhB7GguIa2gEPLq
BXbOZ+0RVJmT+3/AbzVF5Y1P5TQNkkTjujX4nTTqEVyvDt+0OxDIcFbijBzM
Lzk3Haw1NMA02nPQ7I3YvqIpE21F0WM13mfsuw8OntWsvo4ZUxUrlEh/1qNE
2LnIEmDcK1scjPeOEIu/QV8/QdFMuj65irGp/bZk76RKn3/RJDcsCc7pSQNI
DIw9XA1/HjhGTGjBBCax3TeOsi6uYePpUP1dm5vp1GhT36huFYFtebaeIhLD
CJRe49AYBy1Ry4AUAivcpr+PR1fZimddsQ5rU93pPW3IymOAlyTlit2+NX2n
ICE0gVpph+/dw8Y5tZmied36SUc2OEzgWHbuQBkHiPYRLpmkGi4X0NBDe5hJ
3zWuZatz+Cg1DdxSR6d30buLvzJ14bolR0VSD0TuO3nUblI5ujGqyzimzWNs
yCgd+Ty2eYKW+Y2K355FHO+7NRCtsYQowM7ne0AJ5x2XWpxwGQmafwBovIMO
Yh89S7qPr44WXVdVRjcpsC/r7dlbYaJCTGuWMO9QPlsZ14GyPm5HfyjIGipw
JBGZ2IcH8pfxZyNs6r3BOu9syFe7Bul2QzkmNRVub4xUMerlkSBzVvBJTskx
FXCVmGz0vkGbLpGUYDCVjDpFl11YxsGh6x3QBT1g5H9AskSApXazkGDBC1OV
rw6ID13iwnHw53NW/ZalKSA7TV1DN7vBSF5WXCrBMr4Dm0Sw2RoNsgVPEtRa
ED+iHCOXAyGpfowYaHrh0JttegwF6qPknGmu3+ZZvZ1wgR/1OIZhWL/7j6mZ
CfLP/qY74WQlpdsRRjga4OJsdxfbYxWuV43ORc5ecnfiza8JdfbM4YB6MSsT
ZWqbmL0Eq7Jx15tyjAjAyF3FzCohmvlVFSWUWsZhZ3kjBguFiGNBUWqtAfRL
yQA3FT9TKW2MLyfDgonPT4YLRq3TMXUqx+OcEo+xaDBYjkOFIqySiYVekdz2
0nOLi7vVrWgL9syN9kgWMBcp9Qr2byB7gGZQX8lQo/pAz6sJjVtUvK9xMCVt
IWrG3ejLL0mso+H51OQgejq97EsZzYeHmi4xk8/Z+/tDVWzbObRSKrHwCtPJ
g186zLFCyBbGRBh1HsMkH6+DJVivJ9bVwMe6Eg17JZxZGUektSxJPtU+/XXK
dG/xgfgeVIavBrWrozSDzAoG+jKtUfFdReUhEoUQxVpQocsJlzqwnhCaECNf
yLZpq1UmaZYoOYXapFd8tjZv5MhpahoyB1XolEKgbrjBPzNEJzmLaWFKB9Gv
+7kd5EB1wsb8Ua6f4EhKxzSqn1wycXspsQNcURnxLdWCDBvcX0eLF6BYPCDO
nzWwar3zkbFjC4FoJMuZN3r8wHJE6dTwn0e4xF1D5myUFtfrFvJzTofuU7AE
HCY/A0zlUIlEjUEgJaLS0K6SUlF8Jijhg1bITld86Y6h7PtsWBKLyJ6zAlCi
64y2CGo6QPTQkFV+clC5ehXX8EXgN5wC9sjnaYBhuap4UCcYTD7S5typJkDO
fq2XmqXHjbBK/6g3LxviXgssi+Cyi5VhtM3xqwfrxaBZ9Y9XtgAP5oj6pP2Z
6dT1jvkqy5eq1Mc6niMrYANhKUAQDwWt8LYssibSMKtL5qyOHYLkT2fMZxYR
9Gv24Xq7s7plPt7YOyK59E6zuvv36+Z0HtBn1ozEhDqaz0WVraUqowmAHSeK
ga8TxaOqtYlYYH9sB69X/Y5Cox5FTbC1VKcU60Me2Krq/6lv4jUgzMtCm1xo
+9hjC1TKHl/kRMtlk/EAqofBkItUi5KIVOHwmICItp3PJgzx5DNYeTi++TAh
+D9Fzhq8aiJwrD6tKm1SjxNrCkeDg6IYwk4Drq6WeDcrzUsjmnJ/sGQ34fXF
wMaz7PDY3aGrtXTDdASRE2dtjAbLoHdfRVsCNoZyRYM9q89e8ssF7hv6eBqz
9S3yz2dfOsbludukZzNIVc/uPQB3EzBKmHwSOeP6g+DoSyGSsnT1HDQESMip
Jp7gy/GswnuRo0OunAz7mKxqy7t4qab9vb1Xs7joJKpihgcmdEy+xWE9agan
uYJ/OrVYcbTX63TxWOnJ53yGN5ursfJcp3Meu9aYsy3vDvm+127OTbpha+UB
1zB/3TkEXT8SDwoGMQDoYZGoDNM7S+iZtFWhLJNe6MyAgDhQOUDLGp4Yh6ab
0qzXPjHKmwpZBchh8O46AfvHsLG7BOaOIyrZG9B3tlSb7O4enlqTMu9UVNAj
fwEKksdkLKUHhMrYPwc2/dAb2+ibLSYldmmkdv6QPmSB+u6tV99EzZlnHAZa
/icpxyYG2x+/qjrNL8KNXjtxgMur+fkOm54JZOtvZOgnIEHxGGyKszwko4Si
g3sU4gjdrz7N5QBMHv2/MUuuQSPz+1/pXpjrUkXuI6sF2qU2livoPMcszFWi
yphfEuUeM9kPyjn9qDc9fgdQTw/0BvLcvh/RCkjrTpTOYXNsEvOBdycgldxQ
mR/CtmLOuO/vN2CqA08/F+HsxNlBxtvcDjralg0KXtS7ZHXYDc0Dm/kxipD/
h2YenUH/UiU+WiSR0Wy9mLCGiAdTFPfBMyzI3o1hB1Fkq929N/RFKQwo8r69
c8263bHBJzMJftTPOjmhmIW92//0O1Zq7w1BX8JvOu7ZoRCb5/qOV82PxYl1
cMsVd4BbHhhY3XBk2+g+x+2pc6anezJ+GRPVIjKNXSSUYGvkrJ5hQZb+Wzdu
+5jaTbn8ZXkIWv5TkL8LqWjP94NmXIncymqXVgNYUs7AK6AhG24yI2mEhkqZ
yT/79Yi47CyAr1ot2W12EWdBFan6ouDNKtcL+FBbx4m+5NNPAaUK8xoxqCsn
d7gq1XW18fD0H5A/NAXOL+F5Pb0zJiFWj7JVBcDbVnKS149X7id/wg6bBFbQ
JNfh0i1KMDnXuxzLuilinSzFOqOt9WBurUAhAhehJxDNYOxtDANfC3wki9kb
ELu6wv+4EV7X6E+3VDZZnh+rP6WbPFYsBLraI1KaQrRtREBkAWqfD4qDxGo+
5mhA0pDEAgmVYt4/UP7WUiOZi2AfzsfmoWjqkiRpvTepQ9p5kuFOBQqIpjD9
XMXGk3WvMggpSih2o7d4nej2yHERGHmhxBEIeFRJQo3hVnh+y0ZZJT7tBjdX
TkXjFymDg4jLq7oDXE/0Q7BoA+OqMesVp/gaPF5tpsFAjE8ug0hHoROU1Qar
NsABzLq3M7Jg6jglN5vsMezLQND/38ad1nbJLA6u0BiNC2KNhbhs1oa8Lha0
RL1vBlTrSl513yuZGYmvTgTjnmsMXdvGD0+9LfeIIduKl5S5bUdKnSFRwKSG
p4eptGrdM0Gf6qy5zHb+kZPtCeO9dTgagAWwqCS/MjMYiJLnCtSRZ8387J9H
GRUy64ORGCnmzK5TPCrJnVQH6pvG6eoyO2/RKe28mnGBnajFDC1CJTCv8X3v
OTtq+DPKf6Xyf/TT2lfJPWGNDe9V5ZqDFoMZ9Psehd8epwP88cJKnd9lCDL5
YNdLOmEncVsR+mDFDybZDvrPF9PVjos+6Kt66heaJfAj1AW4Qxs/jjoqsW+m
MJgz1E2pbudkgsKwJQsyuJ4HplZtJCAOafTod952e1gWQGWqk07xkA481hcm
0TqVbhWz2BKIXUjwEmtNW5Oeo8X88qUQ3iM1hjVvqVzbINEs8reY9FHboLpH
9o2DyruA/ElGOuh0xuwaf659uHEjAN0+1AEBWWTChuWxlU0ZO2MANrRkbwlw
PMAamrpu8EFjVcoBo+qxf3VDJgLF6Wdxe62H04sxJ5VCAAfUXQan9ehLXBP7
n4saN6M+VmGYFUoU4iJleWK6b/wcPley+Qw+GcT3AsZaUHhz6qe4bAhWNdjU
SfcG1XaE4JEPY/rw0q87lajlCfEvFJx3QbmFVg2DwbdLePw4swm24QhbtCO3
f48UOBUN0yRhNj9weVNw1IdQN3eY1B80ArXTexm+HgDLSS2k6Paq1YsAdDPS
l+eFW3gQk2JlF64pHoIjf1G5wIVGc4+Yzie+WFUiK2mHCLhS3jO4oAuSiS7+
3uCbrLAkx0dwJdqkDxPKR7/YcBKusCVkUq15xtUf2dk+FgKbg9RYQRIA4RTi
Thx76XxBXNUN2wOj6nf6QDG4An+0+L5nNcisHPDcebvcNvMnSNBhTC+zKR4L
HQUkG40CiC0YYQ3/+bZW+7mXMs6qXcfu6CXvRbMDVZeo3V3Y696Wkcr/a4W3
InPVeGT0KZdiYjUvyWH8gnw17cJ4Uy3BLp8J4c0dFP0On8puyscs4ObgpmX/
oezwhOZ9eSZvRKAkmqd7kqxWnkCazcpBmOYhI62Rde1jFVX2lvagHt8ekq38
bh1gvl7ZwUHkM66JZr4MwCIdPYQvmTjtkHyWJd1n8Y1qYvVJlwd19/CbWGMv
VlUlPLHrPYrFVQOthEgOFnWZ6BD4bbbSuSpMmQGR1GypMos6f+0Ts9xu5KCM
hkB3qHjO0dgQgaHS98T2Tn0fxlifBpeq8chSCjjrDvbagm0OFH0AtjtiLDEO
FuodFIKxSJ8qeQJLCXoaQqxvx3yUSXXG8lr7lP3Cf0W8OgDSsSab3BFUyARN
28j54+eg6ARXnIQBsp2frxD8xLcThFCJAxP2oaEns58J3kIko2p2KHdgcOeJ
dw9xuVcmfSR5w25KbuuiUCKMj7r5tW13shihUu6Yyty02gR21yG53KW5eqKH
wa+78AX/UnNGmNtlH4yXmHerNtkxZIMQ4sIo/LZSVA3uzPVoDuDP8g7+bPPy
l1wA0rV0DDuuy41BRQXDaYdUOpSWL6Xkul9wVb20rnjd44z7oceL1O1Xe6zY
SOXVwqOUjGTiuMBeFf8fkZROacahEtfap9zMBGpXxI/6sa7/q62aDLs+jeo6
KTE7eFO8gPGXTpzHCm0d2aS5O83xricHWleuF7aQmZgp6oXuOIhN1AuOMo2f
22TlEDq8O2OSa7E9YnPeKPlgW0UH6wrTqEFOJ25dgSDYitTpHCY7BqPny3Lh
Sobks+y2m0ixet4sESHOI6rNGsio3lzMDMIUwnvRQbAkgbmS8yVa+SAuhY9c
+YbT5v942ZaF0LNE3SHqIp4xsdcwiPqVpRUr+zTq6FcuzLu8G5x1yux5xzII
ZcFQBr/PNACe3aUHwPa/Rsy/N1H9mlJ3YxSvwa7VhXaYS11dD0dVxNt5p4cT
Kaw9faeJU1GRJC+O9CW5Ht+r20CMvOfLud6JcfPbxvkI/Z09RIGibz05J9+D
SMnEdJT/ak4uJ0z8IbpU7k0wy9aw9bbrVqY69hkiv7TSWRjPmDRTPf14irNf
f9qbixjSY4Ps2FCqKYvjwpeRsrAs6wgp3bcdSmSA6Gg4kOSPIMDDg9q8q47N
BChycH+A6tsR6SwgVQwOMGUMxjkFQnhMkoUc3DqZihKfh5wC3xVeMsmS/Zdk
tuYExHGEyrtL4+pGUgwaKAgEiWmsWzC6NZ0cMKp9KLmyoBIeDSMugieKGfwU
CQ0MEQu/8MLBWcpyUaFMavYrdoMJ3rI4dRLTNffe5+tTSvmr76R13b6dJ7pM
JSPbDXV1M4a5KhAAW87TRULJry8OxrJ+LGvwA4AvQyHPzEHzi0rgpCCxzl3E
OTt47dbufFgJlLsUIPvFvys57jo2oseBMv4fVGV/g1md9ENqke5g/IsrrjbX
Jlv38mFrKvHj4aDlXos2746c4AnWhOGin5fv7qspswJw/+ncaN63mxXQdVQE
4USB54oytoHrQSS7Aek0SNo6mGzw9Shkm/YFZktAb5qTZPfVfcCWRW5KUJJ8
0khg76vOOmFWO3d/Ee5Y7zdUyruql4C/93jVoeUfu9B6vOdMPG8wA+tp6JKm
ivOIxay0oK2QdUdT/gmP8aIzflyB4V1Q3HT+v4By0V9C4/++lIakv2zWNVia
5MgV9pDi35KrAwIodVjEmS0uljXyMEnL5rkTD9pUus5EBC2o7/45ghR9f2g0
fVeq60Dq5eWGXQriM5tayhrH4LZxnqeJ/6AENeaQ68gjrAgfLzYyolAoOu2/
gLF8mxiyKLUrSsOF8T/QmxzyAepsCuXaD0eB0gM0VrAkGvTTkYJ0B3YbUkbf
KgNdipPAt+wyj3spWf4YXA3PdFKjykLj+Gpr0Se9o7EtEugsojwZdiJVExVR
C/mRJHCdD7o8m1poCMbiBMpyU1+mrTqhMib/C8kXH4PTUMYR0YlN/hoAQnCV
fAEPCgIOHpMasm6kmHjvRA22e6Bsiarcvalk1giG/S8SoE/GoVP6t5XywUaa
2zhYx472eQ2pzqn5+f7JzYdU+nwDvB8/I2jOUYzMRrANPZiL4BYbLR/Apd4r
KAbgfz/m3hKofSqmx7/IbSAifPV4H5Be3f8FQx6J2p0qhYmrY1eIpEa05KCa
m4lT3N6LYItZ3jCf4uonyRPEJRdu7ixIIIoQbwyIX0HK860G+BIWfxIPMJDs
Ygg2pdkvibPabw6Okbb8hIZtELIvyW48A0txh2ZjicABJVlrFcYxrpP4SaAk
GoM90ZGJmYofQlh+IWJqNenrMmJmPOhwJJiXcFC9nSoIu8hl990khmjKVb9w
Xrp8MevnwOlXy3uNAH997s0jl6xDlfClA/IWVsY5AtvJmd0K5E/KCmXi3XeK
yCwGUXFjpqHoGmC6OOw7/MBEU5uWjfk4poWxCLGAXd1bX/noFkThOtR9GaQV
PnsH/Vi/VsFMmY8xB6E1v9rJpgX0A8Pa3QzocK87rg8dQuKKMtPjRbUAFawP
iIJjtfynb9/PpVXdoCMdv34ySzsRvSRJfe4MNxkdQkg7zf5E8M+ssHqVcQms
pWUCj5/s0HVpMzzlypvXlmkniHGtivapjpB0nkQ9IN8aLNid5a73GplDXaDV
MafOIDyrnddS6FyuyDHmVF7hWeFhvRfr7Hjb/Hr428q8arbkI8HnTVicXBTi
wrM9boXDkgRbD93GafLutCudKcEv/RpjH+5ISWDtHWgBXVJRLkQ1uk1/LKoE
200SEaofrP/tCYCi0Kyhh6edubXsJtD/ESbXEIGlwV+M7SVGsQ2ffsYEryzN
vb6ldUhGoURMHMIT+AgSKhTpnlz0Eb3hl+NVzgJNijqsFOnRxSooHo3xph2X
L6JIHQy5q2NR2K0PP7pjrYU0vjBKc9QgmuHPzhmppJMHOn5TB6a1uodCaWzl
sBSAyqY87iT/J6vwUT6u7EyYf5G5XC0VO7iAfmtfbEESaq8aDKQWQCRgOJSM
yAhP2Ng0q0sVRnl1LD4eEAZEsph+oOUFlXKzNaEYY6XJXFjdHDP8gjT+8bIT
VUcRIclbP+L52PF1A6Cb7DRED4yJ9FcYCaG3VY/BNWc07wTQLmgVr3coUWCf
PLvYO78KKRNCa5iDqt4w9cq0zZL7oe14Ebh9gzZhDfMOeM7f3hAZdXvouzhj
YoVYDps+R9B5gImXIU32CHEVfuZLD45OgChdRluPk4cPtgmXkL8QJnqiiqph
YkJWCYdq8Egu2MupbykqYgFUliHShuPQhzCJi5why/VAiDpnV6uX9ctWNBvh
sklz+ETpe2tYGK0wY940SvEhwH0aXxsMuYityC9z1gHJWLu3bmYIg91QVtJT
SvFeB4J07F6V+atZ1ChyOu/gUT4SqAbDpDSStnkLZwxD2VA7XrO2TzCPNU7Y
wehgcqM7QkFSgtoa4bxX/hCjnR1oBRcDbuUWyDhjcDalsR9kxIb+iVjidA2c
7aazAgZpY8TyD6SsusZzPLuE1Tf8r4jMBH39f+5vUoaEqVwwmERlayLqf1JO
cS0d2E2w9IAN90+kHtbB72UHknuvpzfpwlgZZzkcLk80CrXPqJwjJ3XrnP/K
Dg9zoxRwhjJaaJSThfcx+ICrdlcwahjfghOL7GiJ5v07dTfKQ0vUPmluXa6a
6silGonRQHVWEfev2EK/RKNs/0veNWe3jex/6bbqw0gPyWVRQXIUBClZhntT
kYupKtkP1ppijoaf4ZkT6Ox+9NxgB+gmUL+ziLZjzBwUVVgEQsL7VmgvfGsC
eVKtyjOccth3f2LmWBfMfWJjccCNvnlCqvWu/cYQGvT2EgIYidCy44urmRZ2
Yqe6iwaIA18UIL9UzuJOGw3ebEHuIr2pXBqpnKoSBfKbPGPqc7FuHX31R9BI
BZDsSzhBcvkvUcEAy6Ppe/RZQ3IO+ZVsP9bqBnE6cPy/IMtcTe5IaVa6vk6g
I3BgYwN6KKWd3eHnoVKmDyNyUPrOmNgmT8oAiYki8QQNvixhqW1Ls0s8rIHZ
JHL3lZluPDBVya5OzjDjjtotutvoXVh2mUwpjMJT3rB7PqQQ00JmJv9BTdft
afdnTqtAalBb5U4n5/18I+yrnI5GrzcSUe9XL9fkUdIVMI9ZgcyOaDbycPY7
1ytKbxNBomzHOw6S8NIL7HsLezAavykVUpEIbtD4LfPZdWeVuHD1HWlUqr1v
SBuSeCh+gE6epvo/nDLoM6bjb+mFGoqweQ+YTqKvPlmOw6VVJLn57LcOrWTN
zTAlslz3RthMFWbpaSYF7TnpOlRmvZLrAz6JH62daHjfSgI87H7hQTZjCHXj
oTTuHNOR8lQrYFgL1VTmVMtJMIgZmkEKzLCV4z1g5r5owoso01FV9M7IbFPa
O3OMBHZF1x2eNtOMQVYskdbcUlHyrWd/D/af8DTvSo1esNThJmmnNgcUX9Rp
4X09k5SuycK71KgUgSh9m48nifLwQTNtQ/CzkgwmjDws+Zd8wGPczrFtXHqD
NEOkI+hC7PmCF0hdNXG01a+62V5R7gqUvWzH5xtbmIgKndBLXmOT5K9fT/F5
VQVEZVtk0HX1eGxxHRTzIj1vy4UmqLc9FV0m4krhxDgfrDrm1WWJSvwYpqrM
qGkiVScMW8rWY63eDYPKAEgDn3VDSSUss+6XJ8tmrfEkaQfMHcqzehvWJcSr
6eU75tivc9aWQfLHzHgnn9Tycqd73rVxf285SHVuw1IO47tjNYw5H8Dq6rM6
EKMFCGiIL65KDZ1BF56zzbrzNIm1RiWMQVUSg2NE817ER67Sd8pMAxW7SlUL
kXqbiZHAwsfZ+AxmnPaGT8nVloGsn95VpPeeg6VvVJ4hxKk0ZaFQJ6XX4sAI
Ka72viqpOVELCjSe6Ly+qnQzFuprnQaSsoHH2ZXzNNczbr3VkCsW7br7I34/
OE9LuBI74pMozdy7UP18ElQrRRUeCShJdTWwBtnx7+hbq+ez/flTVWrfkqWt
5sGnQgibFTiBbx2xmUs4KYSTFBUQrVvKXCvQLM7iTsKR57rzFM2QWW5Q2fbv
J+oplKj5iQkwDdm5fDklkl6kjaJ0jn39s6rEO220IO6UJDH0oPnsof2aRZLy
CFhsP9weUL+7ClOaI1j1kAdPHrMNNdUyHX3A2nl5uWJI0fb3wH3mTJjE3Txu
Cg2kyXPMzEkyI2CfAOdrgMXsOvl5gBLhIhblEOFqLVdZtubi6K+Qh3FSTLlS
5iqGRkfgO2+N9YnhRZNEnVVmsWVe4D0JJfswYn2k95dnzdsuqp5nyHOmilyu
7rgGLOW1ZrRkpF6cjluIPn5vSB+Q+skHfqIwQxLnF8MQQgCECpWa7x8ZbPlG
IwdoT6DGBcanJrDxRaUTTzVgr1eU92H6NljazAbNlpNBalmYKCy47J8HhfNX
dPpSqfjtghmcDCPXgEGxPiF9UemJxq+vlaI7AmXEexZTJ1in46w/2eDp+n/B
5VvLce0SchaWTH3EvxKHojnZjRY//QatT7pwqpGY0WqFHaS9hAEiqVWJfu91
nffjjErvrq1Edn3Uw2k7IC8VlkpB2dWrZrwecAwaWxkMLTH8i2zw2P4cFETG
TEWAfRl3MjpRtAEz7eiHgpVh+6oZoKCEY/lkCOifPSnhpybiT+StKZwXiR8k
993eBDFjtsiUqrv/J2/YPb/uy5bZfXrHXxlSH37a4GaJwv/58DwMOwim7D3Q
xncjS4yG5UY44nboj9eSNS2uK5KqOAXAsevZlroJrDB5LN7Md723muKmGkxP
hNjXKoQ93rRDg2Sf4gTEdW2EtSvQhyL3zdp9FhDzoo8GkBBQgT6lABE+3EFF
l8oNM6is9SYuqzQyZzseC7J3LPeWECjrqXO3Li6BoeH78bknyz9+vyqZDA8Q
ETRM75Z7f0bbkss3F/jxg7f1ugdMfwSzQMWFjgi2DeWkNtLYWk4ngMfbgJOk
J65EwHA1swOUyAU23bRmO6nFWCDnyukNloyBPGwWFTR2pH9MC5m/A8QSacjE
WpytBQ2N8bdDRwJC2ryOu4NEAJ7NsrvNUYxLQGmf1CWPMY4hX/MBQk9CtcXY
yrtAXZpgJI/YGt9OYBO7RO+cKoUbQ0UPXPzaM58xCubAIxyy68waoq9Pej+N
uTT7gnb+Wy3I8E+ki74Wu/PPDh4ZQdgq0Q9pYRWCPH2kAqbGdX6RRSj0pBef
xDZddYnWgmCa4i/fsxAHG8y054TteDYV7Aswn6RuGTUol1vnKV5bz4P8Chy2
vI2zymN6yqI2L8RLSsXsLhy2O+22tDmGcOQTwWM4hb4YvOcSgIk1/ikXFhJw
YaRy6Zu4KblvnyiwQcx4aH12ju925r0Q0idbxI5JlUJVqWOq4873hErrQpxz
rmZBUAYPsFK4dnkJiFNw3eRi56FwDAWkRWIfWHT0lw4tlkwo5bV5G1Fc+yif
oYFhxJBGN01d48JTZmakAwfGAS5HPqGpsGt2ECrbcOBlQTgLG0TOu9lyudFJ
LKd1EXQHy6BqxpaZEp8io63fKBwB9khRlBqz5Bwpx7W0TzgAsFX+BKG5vBQS
x/Mj5AlnCx6/HEby3kq6SKhaZBISZLSTRaTnOmL15jgQwaEAbXR+/hvedXhE
BQ9+VVn6wd6sc1Bo4VlfKhdpudEy/lEJ/kyZoTuPyM/Qg7jpAOldwRk2D30V
zaBtGJt6ukad28qeolq2h0+n0BB1v2ZkcZzU/U00a9hXQHYAJGUZlSGId8Dq
8mN4k5FokopgbS6a2Ct3avWgB92zd72b0yH2T+1ZD8dPtP2mx9ZYL7bHqpqS
QHeSM4i3HTTufJ/s79nLP9OtDbgE0JFhGu3LKXk5Nj5xycu7ZQtKHb3u+4IJ
85DuE3fe2WdT1EzDZ1ia26a1bDXLOpuj90qgHyUHf0sXYb5phdwMjfW3RVbZ
gQgLO4jFtBtQi100jxvcdRrl1LXErNCnweSm6QdqosMFChhJNhrIL0JoydqO
x2+QwkHjmQHuaRt2i+wkmrgpg4Zk0pns/yNYoa4rKJwWyYM8xm1q+9HXTNIZ
bKIG1hOI3pd9oGa+/GMaVGAXJVxRjHVJt0dk5+3j9JBxCO56uQPQ/dx6LyiB
wMWRCn/BsAy+eOJlAKDL9g1YBs7a3Ef5NnSktpusKeohdug7A/FYPoF0e7Tn
qB+G9ApGat4irzHzi61AOr+U4zdDxQIdfejNihxHBHKeNuwMTMH7NI/yo2NV
F/Y0ggPAOXncAEPxuuNLwGImLYuqbAttJTNEE4jaSTrdLowbUg5qldO3Mrpk
qjGEHRjo9eY/NsaNcTM6L2A9j8Pn2am9pmhRu116LKJ9Wtk0AatJTTu6Czla
CSffbZQuYg9cRYzytsxbXZH/hYE4u0E4jW1GiK7JVRJ7mVHLWSHuJK+2OX5b
EyLGvWNmnIzHREm457cZiaT2OIDzf6nnkiUG0xvS5IGlKZV/8sT09tq47Epz
bOVFOHFv1EMKEGxj64Whd/aQbinQCbPsYH3FKzDR8wOXjBYaJIdA2jpeuE6q
5ZufHrDSDRWG9OKhPn79Nq5o/fUf3+8GfjeY67TLEPIAyMfg4fKFJMg2VYCx
UK1MiYhpn1HqJugYaShcwTLVAgGROBvdEFUBNyd+M12KBxlfTK8jmxcSTxJ5
hPUFkkJkr/vrf91jjSQ+YEp4rJM7AydE2vrW5k9XJaKPXoUiyQdpxhlVfkTt
Bds9av+j7OGecf/lF3ofIHWXvkZ78Kh6IdzeRCMuug10fp2wr+St9KaunwH9
0zmg1TXOe61DkAqs09HBbiUSgGFpJld0LcCDVg6c2uZo8RBSPkROiG3HrDl6
VEhxOq7iFIVCV1MWHzZRAEEOxWWYjDUnvAFRGMdD/fOouXWeJ2PPtOPkAkoz
d2+WCuHT2qKzg+jbQKb50yrU1e17Jm4TkJHKilSL+m2fvo6/7PfDLu4lvFLQ
sp4pdGU25JLqZ2mK6bDPi0mFUlRzkP8F2RlCaR9j90ObBIJVm9DOSCqAf9Vc
/86M3QIRa1TQA0BDt0Ztn3P/Yk9hSU/fXWzWPJf5a8ckz2yesMNoFIJ8npua
TSdR464qveU2vymYYKTYjzjWv3Bns+mtcS/eFnsMvAMExMsgSnFyOjx+wvXQ
6Yz4TkHFI6nXnMOITntl0eSsUOxQYJaq7Vuzoiz0COuSctP9xYVrhap/e8us
JzqxeTxu3O6jrV+WvLILTOyHG95TTSxZh3mSGs4vrJ7iM2u6Qiq2CK/nc9fJ
imviERjTsHXu9Cj5eEJLAPQQtYon9ndW46FtL4eIuYPM/rqNNEXjUO6bQBoB
e7NfKLxARVkKk6pOPI1ei6K/JlA9bmMZuSgvNla720koIdOCdDNM8ZovkTna
Ol5X4Kc9BMQL1A/n0xunif8x6mjMgTrohDPM/obGjub+7OX5W1LE+guUeFfB
OGudWYO2MkfHKtCqt5O9JCykVq9OGRnpSfncuUuXXqcmGJr9bT3zZH+lixot
9T5PvxiOuhheksQepJPaJRxbkZ6RYdlgLUCuGpg8gaGauinge2rGtSkg6wLL
2zzRRblQCymW5BJJlS07NXq5QkWy8b15mJ1VZ6QyYu/kM/SJ19whCx933Fr6
uHD5hfID4kdgPkePWtXvgsWMjxRr0cOgLKSvQcBzUU0ODN3N63chpXogh1W7
HLpP0UKib+QgpHcrXBvv3L9lwE8kqsbAXiMwAb6CZQn6PIeJ2/AEB4NDgEG0
LviQ1INJ1CJIHGlIDS0WGxDWqH++DEbdPCeb3krQdb7RXb3SXaYW39d+yVUR
2X3au2gPflhvvGrOo4fCv9xEFvDSuAj9wHgBRiFqUmVtiIFNCmgzAEjW+Qwu
Td+ouSK4FBAzhAONDF1vtlyOiJwQ5PJLYvFU7NzTdyeJH3y3DOp3qpkat57H
hF4atGRiFgshfITcPb9RJBxQsQTctaw1GyOmh6URuBe5d30LPOu1WEC58gzN
/cOc39rIllIRTUnJ0ouiYZIB1IaDYCdsHLsd2LCxXbnwBs9ttMiQNAKO4ZM2
Qwp9VjTwKBRM/FemKHVm/mRwHbsqTdvfQtdD/aisaqHAGefk1MBS04F6fO76
wMyb7RC+QO3KaiUXS9x0S2YYU6Vc8+MYCjqNaxdeWT2v5i0dyWMtM9VSoUfj
lCgqkrZp6OWoaGFA8/xNyz3u/bd7smV1AISKuKjWqLTiY7xHtAlSmtMRmBzg
79w2G7smgi/XKauRuG8uoYwtdu5TrIGdcwQxvAxKf2Y8KbTdbLMtL/jK16Kt
RoTjMLi1ZohzmyREL+nIbz9I4O/LDfkPYWDcFdeX/YS1liELPPPevLXKd2+N
xlq3r+mhIfuSpxCyYer1E6ULDvoYziYV4jdc4s2Mzq/+jZfcXUQJG2vbFvLE
xLRK3WP/Ytq/qd3suieEFNuMOs5kGOteUkWkAdNDjnQxlBaLKJMTPF/MmCjO
BLwuTrHHk9l32kcXSldpK9WHjMA+qBHN65mYpv9UQS+vTftmwllgBk3dheQ/
Oblupj+LQlBS4ypif41gb3SuTztLgiDTTEDo6N9OAq2g7I1V/FmgwORxXMj4
5wDvbsxmc2N94noR6jSQsYEmKQtz3eHldPsx2Qnp1s3bHqD7MmIeRY52xVYU
wer4rZTkOSSgPdzozF6u6heIGRRGB3RKjJbITtEvP32wrnJ6N5XGgxOvGAxf
W+k157WbFZDoflQsB/nciPjP4Sq62FwPW9eaTRdh53Vf1NNGs0NZD185550K
iUNkpVgvCsgqTHPhCdS626C+YK05SaqdgMDZZE641MSVMDiIHqvP2MA5nrlC
4Ej2OUo6RFedkaUDSkAmvMEo4gpMjLrr3AntAYWGaS3rgoHaymrTbt+Z0QfG
YGpq8E/kPAofuf+75rCQD/tD23yy3Rpq1B6nMgaE6KJDQFekw9fOsxQXN5wD
LwYwS2NTBcBCP9ZNMyUo5yBDBkhxrziUTFW9JrEwrJYa31uF+khYmEuyhcsf
aHVvY3Ip8Oa2JN8KOLd1JSYECuGOYNMi8sY5SDR/6DhxkWImTQtCjkmTSOgf
70DXNCq+c+5+5cM0/iVGWe0h3s/WRNfFr0zY/SrZFuuE60s3QO8G8ASJlVdO
EYYubiNfzjfIppxDIWxH/7HgH/kpcYuVh3ycVXKjv2lw36raqjnsaAs1d460
7KHiok37iYkRJfvINItERHgZnzTEaFG2PRK9CbMpUEN7qtExEJv4WgDJCS1Y
wZWB1sVc8LPFaYZTxCgjWKBIlFTixrq2q3S5wT8PoLAPMljurAO7g5vgfKAj
q8YSs4JL/1aUxES0X/3nSw6eP0lraMc6aXRvDH2vUVoENWwRcE8MtJMIt3yE
w3clF/DMtB+S3FkMBzy+vjjIZmvkAgPeNslsJJrfNMe5NuYtsmtOEpcSUjZe
h2eyBOX0rHHRVdSE7FU+T4nHENu8ctNt/pZg5nKebnrJlTED+rpZ+Lgreyya
XG3FUqpuRYMTi0vVCYIzWqsxSS7DgKm2hrdRtYqrHZYZyRcj7dLFtYze9JBu
MsBgM4E0TfJCrX7O29PykBACCnxFPWZdM+/BKaN92u4BxMllvmpX3oTy6y9X
XZudsdsTiFz4huoXOPrK32kzRfTE1n66qcobBnKYg0JJykjigTkz1s+QlhGs
7mzWQ+pVVWBhwaGNKT5EIz11qBmwQJPfepVnjk6rjzDOFLst5YS9MYBdyBdk
/p/gU1nf8TuG82oXTi45xVzb/6mOqFONTtJ/5kgMnidtfF0szQtIg6ADA8mE
3FWA0v8We8AGvWbvW2SfQcMl8Fgk09CdDjb5u8/fcK0sozqzo5lNM/9tknsz
SCDuKd76LI+8Iftm5LGuN1o6iOdMs+zpf+ljrv4Pzx4DtMKFmZNZrl5sfVFa
XpN43iT57o7zROs5QI0TzuhpGVeJbzbdubnTLuvT0vkgEmQ+evexY4/b/I1N
65zGeglCHIh0hshBBLcU6fVa8Rs0i8/UXgXHyfiA0taJuQo0y5mOsUvdCOiW
niwbyyupolSdC6sVdbVCIuMfnuJawSNj6IWHONXT3IEMYq2kRrBYjJxlCLHP
z6ao+wQpQRH8ddK4q2Dj1ojdmfLjMrsSJN681/e0V0Yx28NMhw5fJvV7Rj2t
YXEWS1OjUmcLJUXEoTc1D3tihY4O8Najbv7CDkXTFKQkVA4oMGcFBx24NWvV
EtHXEBIwZa5uTLDJ6GgARAczGxI992ESNpzJcPgg41ICF8axZ8NV/1uK8cpA
32oF3UNv9DW0XenAFaye9P8gdeIiU+BZovtSFeDQ9+NL+mwlrojTcGBAl2qz
MW7iFUiyxVXAAj0YUPAbuyhn+tLATHPyQ3eOABKs+agE4cPvhO8UjGVEu0vP
ddq+pC61wh6RUqZkcnjMsBszeRzwmhpykbc+3E9ziNo6ps0YFaxjq0nBX5sp
uchylzNlYFIUUc63yot/RO705qjAtz3THJRkqZe9AtGlzJRkAEhc9OIx4VUw
NOBhTF/suYVFC152dNtGCrijbPmu0in3O9NRsjCr/XFjErHlyMGO8tJQWElA
maly6xjKGGVTI7BKCGuIjQ669Abg0fl1qytMCAywaxLbHAkJC8cslhmSZ8AM
Mvw/VfpQVo0QK7sr4GRYFr0XuHoKhLz6Qzhrq6DjJppBNd08GG7SdCSpuy/Y
+tnmZoCkTNA16cn4T8vERBFgZGkevAzh+slu+9UTTnBj5Tsjvcyu6pf3x7LA
kyNEtEIae2R4/ujKqunIVpXetDcZbsAxB4eAODAIWE6u55H9RjpdmR4Owv4a
BMWr7/j6E3ll9r4vt1Lc2Eri0siiown26WLpYtgLOkSIkdPlDKe3Cma21MD4
r3KGCubj+17Hh7k9ze1thw0eBModBjhX32WxK9GyV6Lu4kNu/tsNx0+TalzC
kkptYDV5/l+1yyPc7jE16CQJdzLGvZ0mjY2dW4Qkdcb5AUayTqZoNl3YR3E2
XBkbxOLpQdjG2GvZwut38GLr2w4USi2tANWeNsNiCg67BXi9PF8aeOpYt3Ob
7KOmbajUBBW+hQqgYXPi6EWl3hPOaLWJhKPiak8vc/IlfpSHJ1QbLTWiiW/r
aBDyx6EG6Ud/PIE20uv6tflOuPHg1VooLD3dFCWKHVeQ38xPL1KpBN7WppEl
dGZq5uMgK0ofuPXg1y9tT0kKOGSL

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "hmRb1hCms2kg5lxwgzvVC1ojkYPyZtVhUZroYIGDp3nv41l/XQfn8gMXcNw31HDDWBFvru7tQ/av+VlNCOY8CAEc3dS4tSN1iCLWoSLzjcf1An3u0nZDKunxPUWY57wMTkfTn6dFEXYBYGQG/cgNqAwhgy/sA9kmZ+yrzAG/xfCgRlDUR3RpN+hQPPycj5HNM2pIgRPAeD/5T2qj/frBFu5c2+SfDL19Hg79cXZFl7XgyQ4f23OwSN6iq6yMUOATqIlF6imhhgvYjqvGcFRkk5B8hs8U3XRFYQ6a3ptIdQt0lnoNzD4YUy/NOO+nv6qywGw8eB34O2a9LurKy71j2VqOZwNzs4kxrBWFEQPiZhPA5KLa7zvz5eliCySYfztEa5N/rOpUnqe5DW7wlr0AIA/Ukm1t/2wyq4M3+b1wGJ6y56klzn6wlbJlhn3NlUw7Z0v015PfHxYAPMSMUu2Yf2QLUQAV0wx+xmgh2lFQJ+ft3BtyZyzkjsFhCmka9T63LV/+sQueBoSSvqs5Vxqpfpgif8cHJxUs+2nxGDyxg1fYN0XjaGJLBgtyS03ql3VAsWv1oKRB+/08WK/2gd35zBQYZymeSlrO0Nb3miphPJvE37Cg0SnybDgoiKuNAx8W393Mw3+6rJllP05npjoqHqHPA6LH+vK39RbPbLMrdzmKUbyECuwzPEQONLyqQ1enMqk9yFLGR7yav0sWGqMniunBYAUvcAcZaD8y2l8oqC2WwWqlrcWkLrS00PqIdjhbpGMDW2HqQaPevxIzOVEcoF99UBpWi3jaSnejMTuK7neuNp8Z61UvcX+VuVVYqwEKvpGqg5oA2ilYxgkMHNX5YmOWjizGu6lIRCU4TU+oYOtmLhXjnJ7RsIbfR7EeJ6wgpl9mUeJyBqm6RtG3FZB1aUvrlsZVV9rhjxYcllK/oCskfadskLwr64rpmp5qZppK5kP9RgRC67QLUJjoVGCIlXYNiqq5gDmzhSejEQX1hukXZh1BIp22dP5PXb3ccAdK"
`endif