// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UtSNNl1k8g2EM5CNXF6x6DcJQ48+qOQeVu0TZRBAf2Oo7NRdEX9xSYMa9WyL
UVfjXc/BRCioDMIm4fAUg/3qbeLBMl6m5Nsfb/fGyoQp5bHIV2VHSwQ0bUBM
6fPOOQ9y+FaYK8WXE5vogUJgAFcCw4WVXd0paaE/sjJ/Z/74YRfcuiFwT5gP
Caz2PdhRgwqUlzXOWQYdq/wcOLkVSxBgsMQHXHc/to752zlUUv7AJt42Av8A
Za41fPIR/CooICDZit6xZgSDQ2IgvCtBUubZ3I1cUCM1U9WhOkkoV3+29SqO
wH+pugGIzqdUL7MYFIafXcdHzgzAo7Yrf83eW/HKuQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ghvET0qAwnm8Wksugzc/cDtFiaUchKQJnOaFCpuQ8jVyeZ8ZQo3LesnNVSZP
RqV4ZVvF1gtKWCVUVB5/FKYB/wvTIyZWXvr3AgsfXH32dDt0SyrF4lmnvfU/
RtbRTughwO0F9gX5KkZi/z0vasp2nIMk784dVnKFmUu7HvBHnfjVYqH3vqs1
gfCQieXnOowbx3b5hV9uNJZWRk61QDxlQf6p6j8xmi45jxowsYXE1aMFO3gs
nbEz9gYOLAzhiY8QrYCBYvfowj2H4yUSq3UOaQubpEX051cypctu1oeo2koi
iT94JHVeieW80+pqsl2FWFBC7F80lPQ51XSbJgvoog==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b2quZTSbmN2zWcatQ82NAukRxcMPdFoxVS7l5ZXs21d2eD0EgVHCGhjeu9U5
VYcNymoRMAFUAiBFUF1ZYpbCZaOqVLDco3Q4M3X4BqPuAxoaCoBbWpgqLoov
Nxyu6XZcTeY6qVBbegSymnlPJUk5jWYBIuPMs+VL4U0oCaURhlqa4D3ZTjrx
+fghFikZyHgO8emUppbRLLUyv758GkBgzpvaeYK+WrdIFU6mzT/fZYZStyML
3aJZLW3udyVaIJYEe2NDuSQw0THz9onCEzhRYPsR3Qg+vBpwrMrT9nqzF7B4
k+9ydp9SNg6YPG+PfzqUDYM7ra7dRG5hFOya/6LoeA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aTd2u50DIbg9EaBlFFpXjeM6df5cF0yv7m3t3Vz8WdWmcyJc8uw/DL40Pxxy
0W9yB9jfzYnaZY5/5kXbvYMcOBLqqkKFocT8dJs8/+mmxfELV5QKpak2hvZH
Yx3K5SMkD/CeAbYUOmvbx10sxtglTHtwvXq3GvpK7MNARHK4rdYuyNUkBKBX
BZ8RUL8gQXjmIb78AAZ1nGv2m4aIxpPgMEZfE6hwtMOqqzgUeXR8veDvCu5E
almLLSpegjCKSIql4JlfYvW+VNvyT0/5dm/rA7uoJ3xaW8c04m5XKrFAGwRf
c1iXnzfyxuCGI3hkStyk2Z6HFQtE/f/+ENAZl2IH1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jMsuRs+vxQwjirrImkhR/11WK68QAbmnVckHy8OLDdgq/xTpjkfsbnGZObMG
ojL05Vqh8Mk3/Er0DT+WoqOw825bnf0kx/i/O5Xzi+HwNrry/5kwpYii25Rt
Bz2jZp6fqxExw1fhBEsMI9zbBnu2RHL83tTfQVwAv2aPzCd77O4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
iz0LeZ7h8ZTJbyBf76EWmmOS7gSTzgkcmCjsRJu7p4OMnzMJTGlDnxi/dlNl
9DVHs2zIFJfAnNrVb3z7Y2MF8aR+R6/O4gXAHPUKylDtkdX3HWzgFIoBaEUX
4AA+NDlr3hDdTrouuzye6fCQSp9wklyAVoBcO8K8fAhnJpQCWKsa0CodimGc
fnmsdFFwoD9uUylpnPQydDqrindcSB96LnfSTrM+2HFCbvSPooG3mWmWFe+2
GPJ58HcBE96oupkjstMAt26DfEtEmJcDc+qG442Q64xSvzsgTREPzdeCzuxL
0LlAmQZKhIfya8cNX5iVhw6JhHKBXygJJTkBO4GYxhrtTH2uIZhUzGm01DIM
SHsrIEdc+FptX/p78Uq1JZ7kf+0i6bMV2XgjDau+STxm0tJgPtLMft+MGs38
Zdfc0egwTklSyz2dBkwQA42yo2S7zaOyl52ut76ltK8ygWHxcVQV81vBKPze
MIP19v0X0ogeG4Gx1EpcK5h1Ty+9rpSH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g+dNYk+ytjiSQ4ENY8t5xaJxlURRsgI94WEGQrFlORyZt6eqQJoF7PjOYF/x
NWPyhEgyCD43RilfIqXOgEzQ+WCSFN10l4tQcK2qBPLxqjf9Ju2u97R/cFAN
vDdBmZp9+t1QudUqmG/X5FYpMmyuPVC+fJ7w06OiXqsQ/L355G0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lCCn9YyDEk8GJz6IfFRGt/+WrU1ohS+rnyUbYHE0KZNSisbKVC+RP7dMuGdA
EICe8kYiAXXm3B8oSgjN7iYLzHn+XPTI61BHcES4wuxctpSPDctIWO2gb3oT
68e0jyp9SObeeZ9wCRdVmbw4tdHnROaVtZlhb3GPmbpuFF3aJjk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 94720)
`pragma protect data_block
8fWWJKCN37DSYgt6rhmGBhh50TmPUjo5Gg8zYYmywVXN3XvlQgvDEuzXA4PF
2vPnXdNPrtrNcCqEdhCw5/XABKZlj7I6+5d5VXclqYPnGJNbMklq1tEjVrzH
Lon1xB4CJgyoyyGaMDJk/UlptUAv1YH3SY6lGO3MUZ+bAu4fi26Kk9znddcY
KM06X4TNjL66FTGvRSayMllbXt4uMeyciwmnqk7jkSEo7Hti1BbIdZhIdW0d
TVoDF1aiBFe2DBAho1Pnzw7YNc+1ejg5RZUIIIwhSk7QU0H+uisTi1HYnS/p
YEiCUw42ReNcmStJAWE1Ix4K4ptTzUylk+Le86CHY8inaSf41pv8EPM7hV6y
OuDaBJTk4Mz81ZDH5hoEKJXtv2XZOMCTZUmwkZIe7pj9UTTF+bthL0MytxpL
sdrMwfD4Pzqjnwb+M1/9PkEUTdoBLJWdhNrtJe70ctnm+CWUlLYCJae5leql
ShN4IChWKH+uNny3FMw36peHfu9Y4aXd1+MjgY4o7MP1s6Pvu2AyN64OysTh
Fq+Ta7D3j9QD9hlgn+NwjIltiAKZjAHXvjSHDY0SlVAY8TAG1JPeWfjhD6X1
XlWzUQMhW9i+B5G8t+dg5l6ZZ1ZJRju3UBw5KOtxWzWzJwJA1mE9MaNp0dfp
7F497YOyBtGdP36kqAflS0a9kt2VACZ4nzje6VfvcSCICFX++I76xi1Zd5lP
ixV9OQNgIEkvzo1ns8U2hUHtrIs7AF08PwWsCUalLPSC5UvTmjob5B0OSYjt
Wn100FjCXie3yzxW7OycTjOH8Z8lKwODSH11+VDIfhUCfpGGhdnko7Jk45aP
Cgbl/8xbbDjehmgjsyeiMNR4qtryad76ukPIfvb2tv/LaszJrGCJziJnU2Sj
KyJUvOdXI8Vd4jpOr7Vcs/t0nBwmTjDN6o3ho6W90UL5G7ZnWawK4mhTzI7R
7RTkHCbpTGisX++v37Rk65pf/hqWrvB6HYzc4k2sQmV2OU1/KmQBVEFXj+I3
bOVheYVKUj538upojHdufcqCFovH2TA5rFWy9LQh2in8JiZNqDrh9t1xUlps
GN/s02pY4Dls8nwJfJl/uyJUCiI4/Kh3nai05w9mm+qC9egOnPlMrr5iBZSO
c97oo0q2Ua9drHVzTNNmYxBPqUmBdQ0htPSUfNTESuh+JyNlLHiHYqPwtzOZ
IXKrN/xe9B9IQE9n73mE6CqB1kql6lNZw7nutJ1PGb174QOg94P4HlkCDxmf
2vqqjelK9gprfKcEFaaUQzDT4NQAIpD8aeuJ0dksF9vfBfysn3m8u/bqO9Kc
0ldj0+be44bXboCvqqy+G7Nuh8VS8+jPq4sS+Iy4n8GkabaAHGD/6LMn3lCc
uMtPzZVxuer84Q9+3DVM8wbwIWtJSBNOXCQ9mpTp5YpNGTPXS0L9ZM/AZEk/
8xOa2Ayir2nqPNBfvElvmaTpDTy7JLOmi/XQ3yghxi6cjNY+AkEb/DdHGBhh
68GCil2uC6lqlxOT4um7RR7wqKO4RyIFkgAoj1hVnTMkRqoE180tpzwvKIjh
hdeuy7/WKtvNNtRyUvNW/FOXMkontZgKU+1/6AShI8UCN2MXKIgG3YT9ZRUJ
u+PtK+/Yf1EZvShm0ry27mWv3AVUOjOwIknVIqp3QSuVgZYk4ddodJUo7011
ZyDRgDHBvNTk2cMkykUNmKREDS6iufiZxqAec1DfXMEn5RnL7KcXsVyH9WIY
mmvVl7UE1kL7KAsQ0ilfagcVo9bRjFZ1zkW7AyUrd6xAb/CxSBkr/gGikqxi
m+4ko0CrX6yzzi3H3Snh/5DIh58q8IUUXmUVV8eOmCrrFbvtksJk73UcGvO4
55mdkG4xa0wBGyE3Cy0jp9TL/AJwoNim/5Ufsbxm1B6Pfw100+sd8g0P7jfj
fauHxb8JOUAoORXMsm/4x9YwwALWdk/NZPWMYaJ7izkojwBhqVKzb22orq3u
0rM2PY1TDpWJ4rNgf1vZ3bPqwmWJhuSghb1iH5KEQIq70FTf3ylXVbI/Yiih
QlS4v9BLrt2qgZfZGzRiDwJGQPDdluh21EtUPNXicydBKIOE+mL3xq1F+NSF
0XkDvgzhkSOBBKn5R1Dy/4FXQUwZvQk/RiHHlf4omsbVMJTUJcGxavgERrfk
IHMtqc7zznSCDJHoEK7Cw50uygP3oaJR4FI0G1c64gfAySmOVqiEdZ0KStN7
WXU0KD+EtVEk+QUJosWSVKTcMFFkNX1epVE8hugzcyHGrm8nU0AJ6//0X4Mc
ADD7cfMud5TP3Y9H6FANhcHtaTGor0Pk3Nc+NLjs2zjZ8uLLPTZSKkdd0NHh
xA24tRocA21LafycFgOBNii7J7iUpjGJm643xaPWMF+dJ6lWzUC+bCqGZ7ar
1E5OOw9IEVlgvjsX9zWdCPfy0W3ctINMGN3x3qKJDM1alnVequrW6BjLloLP
bfy4OPu60nbYCaSHlZHqpsjaBnPsNVjhsk71o+aQoy0kKZew0YQVDgZVWsGJ
5DPQrK5ZwZeWRc/YHUT24Faav4aVxfB9Pb2aNd6uLxST6A99TjMtB4ZtMZew
5onVJiVahIfRQ6wIoPxx9Pbh1wPD+RI8M16dPhhc4QrzgQO5s3gN63VnlHig
i5gdIzeSyIM4UKiPpnf6LpC5o74Ho8Elk8vz4sJvMsjPO6yBEqu+lOPQbaiU
YkpTJ32KsNGA6IGkrF2+Y/oDFR/q2B6lWeYoZ/vvPdIGM8OUJZFUZuetHem9
PL903aws+zDpyc1Iy01nqGHR7Z+YtT5+lprc7BVMnYOzKG9bQiVoTCUnAPMN
GBoRP5k0ktiY/OKiKb3ANH4BMsr682in1gl50AEDmUt4tQZ49qsCOKv/Ng5n
XMdmV6LtJcTcTNDE1eujETdZ/O/zIAf1cHB4cksBGDf28X+pd29mzN2p1FBF
Vve15nJDdVmSIP9N491wakUl4LY8IOGhx8j1yqr7oqTO3Ah5y3l9SEI+HCiC
W0T9OsFE+XzvJYSjhqdRwNhFZY3k7ehlduYruXWt36EyHEEbkFylUYd1TR8A
OSJpvv1/dwK2PtTLAE+i2NpGKv8EsCWN6TDe336E16wSiD8+RE5xpNF+s2Sc
W6DPL8LZ5TCNKKcGD2RithuJ0Fphhc7qYLbQcUUGBzUKrIVZjQYvH7Aj99qZ
G1cqCvUN7PZaT6g5cCBCZ8HOtVad3FC5mFCVKWWWW9UVBQHZrVQzZw7ssZNT
bPRncnhn3iIFlqXhwwbtJE5hY6NCfHwat3fcMB/cLr/L5Kpru2geln3Dsjcr
i7G2i9FE576hOYGdZVVXE6o2tkJjPBLZBcijVaZBgkMosOZjG8ogRB+T0O+D
oyv3ittNvBXrrMojXfBbJAl0tsnRgFkqKWDoBXHqQ9V38fK/2JZXSRu0VeeB
z+KZt5wZAFyRG/MSuSoErcJxNe8cee1J3REpRXaqwYYO1TDrAR45CFC/ImLK
PN2NeEpE9/ogXdvIAU1Dj2XpVgbS5tRhuqyfq4UY25G+ZTBP5JEtrZaZdBSK
E2qqzpiKA2X/aFnz8p/4SqWf2m2FrSwi+jtz7+koUlcl+B9XEIoCbMo2v0LW
CM3dPSXvc2CH3tiaKjnu61EOVtQs7GX8+iiktthlAJb3XszyjuTbUVOO7OPu
rrT4rXp/Zxtr8BhlkLX7oRtco5eWsMC4jbo0LE65/uOam0I0J4ihCJX7tWLp
qBIk8fVU8Vik8wWKV2oyrCp/c+StOn1rhel6GHlk8gNUXVlS5d4G1DuuPdZ0
gbZW/mIeV8cav3s0hfshmJKzxSqHS3GEbZ3447OfBp8nfRVama0uq5YsKtfA
pTfGWNpI7wdCWcBvPetj8gpkG21ThXLWkuWMlw9ZMcDN7UHoUFCEANxDn/6E
0y9QQ2zRNW9NMWWe0gltsfIVTvBJQyB+BM3wfGdj6bxGu/jZLkE5HySdMqWY
AUoTuwvJGSz7IoaVdkBAEw5plJsIfE+jWGSuG+fKMgU9emB/spfHilUOGSpx
i3R+pOrYkXZeE2VlHrb+sLesDpLteARs0JvFSuFZWWU7QnkVB40OymS5c7dE
13X+gI272OEkLHxXZ6X6LVRlYf/p2y9v39B45HwinlxOkB3OTFz4NyYPq0ts
GrDRe4ZnExN6i9ERq0DEY8fl5wMOyWMsi5rDEgH7iE2JNQ/I1BJ2MjULlEhb
+KaA9SPpCBaqtQOEo654ufH5+hXC+TUXhtZgax5NAJB5PhVB28iRZwKZMW8p
ouLwKQRUGYDdXPKPiAW0i50CYbSGsYD6VXrYyhvQMxc3hHOIdsjJEYbspLXI
ExYnSS8XXl3sp8Ozpm96428cl+4/JrCbpP/JXHi1lqa+ZenIoBHjh1lE6MHz
x6y+P+audyvH58tUZ4vZ5O3oK/JoH4EZrUF5kvesG7c84DXrD5cRNjv3VyYY
efk9rkxHeqW26tGHLapBDzX7DYCLsJOlRFyANovEn7oGOJIE66HJveabDSSy
2oF1z2/tfCoes/k+unIn1SExN21xROwddtPrGYACm+/u37UyUaJKOYKW/EWf
edRpZs5w5DBn2x9jmquP5zW3Da8N8GQMnFjJYESKXXkzQpf9SByGyleiyj2A
4/6F9ucySQ3+52ZqiKk+Ya9Vz1ME9uE+hcb7Ype/1ETL8v94fmiQ4tjvqMF/
N4WEHn+1VtXdBeaW6k76PY2V0oE/ytYZZC0y9fEHJouuxsq2zRFlZkqvMeqf
rasNxoLrPSQR23+iKO33etSqm/Dtr3FWW0gaJBQba4jTOf+8ZbEfPdy+GfAg
LP8LTm/bCZPzdh9WS2cs1O6MC8dzIIIZr/dNV4KGmJVllnbnLkULInIkiukP
88JA+DRc7gmedPAjdAs3vDIjQGE0YLAua/LNTvEFuz7MNL8iXyX/60btJrbb
iWluOP+TgPgsb+0Po0YGfDaHFnMyki5uU4teNs9Ti/nD/wmumfnDO9iwMERm
a4wXMyxMpkb9lTUYH+cikhZzMif6BNGUX/o9hsL8PQaAbp0ix6rg/GaOmOkf
vpHDL9lgfJfnWcR7LIDxsjU7uO2eZAPVeIaP+Bg2iFiehHk6BDCKWQqmvWLC
K6J4qOrwUCacnqfd+XoDdHun2/D6+xzMduLoyO90SE7Srif2kD08/B4Cr6Py
NnVXw2WQ/F9lS2p8uyj89R/f/JTern9PpMFyq7ke5qmk5YUi/G/eRkXA4RZv
LkxSZBE/bnP6wZ3IBDCuK/SR1TZdA42gTuR/g2WShHCsRgiB3Yb54zT1Aqdl
StgsmCtMLsZLvuLQ9Y5cfAa9DSDzGAkxVs3L9nteyBsHF4FbDvHB76xMhDQ+
TOKUAmUQBlD9YiRROWR1Uvz+8BiZpbNgUSdrDdcl3z0H++6pheYIBqNErJKy
updHQLXvLtcVLhEmSeaDDUYpP9kusPoiEM7DnhlN7lOK1RohLN4lXhFRWQQA
6gICDZHlhchndyN4T09D2ztGvQyJX9srhHkAqoL1D3BbcLM5Rs4+z1E6Ko2X
KbG16NipLYKTE558rVXI4i6X+1VKzh+0kfvSDnOFOaBto+C2hcCkxqp/vzt1
yk+puf4DPGNDtIpMw6+iVDhTEcKuGorlNXi5r/YpHtVgLiq+jN7dqoLQtaM1
0XI9LdJc2ul7e5up3/QwsmvVnpkS7E1HW4kUMkk/mviLjlhQEGYNlrxL41dD
AAvNRiJMi7jOJ/Syyk1wB9dP+NA67if0elhRn+gqP7Rc92ws87FWqPx/qmeu
7jMPhKV1/xN2M5YOe9+e6mAvJgnheZ7mUUJmRY9F4HoRAuIoQV2JppZlcrJ9
lWVKm2p0eTlE+DeKdJ8n1R10+027qJLt2ZntJV1h+bzbk60FCwLZGK6gu1O7
3VfH9KfPjIxbS25JXp13hUI3Hi4kE4axHc4jzo7FUNgfNbJPTXJwHmm+A4P4
zKi6jjygKIoe9QAQEC7g8e7D9+0VRm/VsmGNI9wPDQ/asKxcBFKLGzkNx3Ih
1a652GYhxgVY8TD/Py8e48W+557NG2zeCQyMsRdYdyQTeKHfwjWg4nJo0jXg
OTBWLSmQw1CHN58ieetLEoPPZrT4K0CfmAm1+EtfwgKl+LvV9OktGqSkuJtD
4XczQ+qwvmL4t/nQFiRYOjjB/55o3QSaQr+OgyOx92LsqBI6w/DdeCMiIuOK
WQHIXYdhxkI+xgkT0yslGBIzLQyRFMRsXBILxWFRmdQ5z/60qU0swZeJpFwZ
BCCreXLmDbY1XKkaTu9hMKSk67mZJBURTXAQSsjlrG8klSxJCccnRZ7GG9Ak
/C4uQTHqc8EXrWYJiNvvY9xI30V47MpPOPHf/R+9UYgg0sOM9ICqlAUxfDiG
y8KgVU3tdcEbyPMC7hVif4u68F+/Pka6jg280wVw/vHw+FVfRnuHRp0jjo/Q
yQczkk0aKadrmEHFaUY1qZVoXTgTd6MGsSVOfR781M2TZxDlIDqBOdiClLKR
Xba/hbXxbDEjCGOSm5A6wWGFWePCaMACC098CsuPI9kE8bowfvxiJyEaRZp7
jLjZiZVx5hVNaOx0f9vpdv49QOdj0TVWU9IEHXpdQRfv9VTiWR04nTa1qQox
xKBabT9GGVTai9BnQsLRCTpU71lghTtEJw3Tqae1x/lM0OVy9BJT/3tSiXVE
xRE9MVUYbkAlHQ3lVkKz02o/s/U2zZS1op/SDc28sgd/NpDn8+1YGn3xNBTn
4dbG14GqH1gjCmZKtqMjY+YbjPBMwWA3klRn9c93ZZjbdMTc0d5snfDKbQR9
UT812SEIgKXAE4hXaNcNHwa5CF2oOLZ37sykqibocst8icHhahqX472YwvPK
2+iJF7YszXV7d7u8XWDuTS85pVCz47nVALwCyFVFgs122dIBYRBfTf7PPxgN
tsy8u+9d3mYZtwBfzRpvAAJh2H9+jfa0c43KEAqSpZRVKA4GtN8AU+VDsElC
ZlQ6r7VjaMaRlcNSiTkJM+N3XWasZV2qutBSXwxm8LhDsl77IGu5xNoPDRJm
Nh9/p5q0oBDy1GkqBoUzbtyqOwr2Oarf9VGjXnEu4hmH0gkY8V4z/e+rwp9R
a3poSYW2MsM9IH8TgLiP1nTPOmfX5LThYduA+lc1GmmvirFtb/UEBCxipDG7
4BcBzSeUj5Im/a7Xv0aKc++01kMz0kF+27QGXpXdQNa6WnDIbFJLf83Bwzd5
9VkS12wZZbRG990K3bst8JIub8jmfSB/UB4o8o5Xo9MRIP0Ml9jQxKBeOWnu
e1nFv/+MQdnrFLomZPCEpruhbfPMciVtvnS2C2HasnyzCZKA4lgQBycIXUNX
JNvTF4SJhie5dLxGLpW81BsCFpg4v+36SH177hgz68OBMJGPriwqX6y6sGqy
jVMzy2r5hXZw9Cdzk0dBlnRYZM9oWF6iKyxXBPqheGvOQYOs8mTDP9TarBsY
0u+kCJL24yS325O6ks3IMonkLmteXvN3WBbyU0Fhum2fx3LeJhKW/+2BrQb+
QYm2yjBiqmebnlOV79vYePzDuHtqysWKQzcbetpBMBex9jqt18D1yz7RcXik
mgIe61xnz22s3Bok7E25KXBnY9d8nFwux6/9Z56UzO+4JJc1V+ckfI8TD9qI
52pd0klEXplTNkP2aCGWd8HYfZ5LTiErFOvvdjtSMa+SDF0oyJgfVp13z4Ub
7CeUok05FOUDGUtOJWzmWI5rMkkQR5ENb0a79Cg072DC35PilcHJArm3x1xr
rSrhBtwsIq90BH9mQ2h/iTyROg9D6WzPGgxf+57Hw3zEYmykD7bz/wiz3P5j
FhswUP+tkNyf9YBzN/kVVAotbTIaucFN95LfgVfYGDNamErAaqAfKBrygGGu
2JXxq66QAZcBRWxUtbqO69us0xSngJx1C4HBMx24AW/QNWyH/Uye6fva8E+L
cHQZOoqvN74ykpPUGS3yrm+sEMXHzHfydgKnh0iSf4uwaLRdOilCnThaIvEA
vuq7htz3YuOaS42qsNgofg3Z7Xx21X7AeQXK+dlfYF7sCc6dYAr2LrZL0Z4b
5tTqobvaaCcqGEVffrZVjeokOTCb7Peru/ZRiwH1Ff5LvxGaXjAy/kCzKUsB
/It7VztctmIjR3YT5rye+wAZ5LkXrO2kX3F2K68b4/OtGh8Hx7P9JMWhETUu
NIxn61xN5Bz4h1G7KbcuKDqNHbha/htDUZGLuuu6YQ+WnXMe3GHLh7jAAKKb
CJa14+LZIm4I2BnPefA04XNwWy16Wk3iLkzxXsgJpkCo6xTURSS6HcHx2GjF
FwWQal0sI/IoXsANtRHoGrAqZSHVsF0+8KVBA3D4aMxtMjX1jp38UvwLHx6u
U+KSHVML3eDHpPL5xc9x/bHJGS6bRCTtjj48jkitVEjtuM2zTgBVdfDqEVPf
hRpaJLNf6Xh71BvFisFhIkE1qRwGHN31Ti+KNHEzTnU0H+xxWzSQJRb1Icdm
YNT5qOif1I9/HEEs091GpuiSbLMVi2u9G9UamuLPYBbglQzkQn/MKfmqS+z/
qZs0A8FaOwqbUwHH6lqq15aJXMgPYSt9MFknVweF0DLTRkPjFrDlmzhZ218W
wFgXv1jqOnP6PuFvJT2KlZg2TA3O9EcFG/8Dp4X/ncaEj43R3DQtjTAabnIY
xuNHigCQMDCH0ETPLxzSfIArwYwgkEtKc2BztaJDxpfBXF+JAu/rse0V/ZAx
sKUJxRBr267mAoJ5ajdkzuHXl0zh2YoTXf2tE0/+m95eJbPDwJ/9HX6kmYom
z1RyssnK3CgrlfznLbLHokJQ7CDWaQoBrmm5Snq/nH2DJWqEye/sbAL1YRNR
siuWR4dJ0U4+m5r3QTKc2hUOw3Q+FhwONu/uDepDOZBYMgK5agAy0L8ZiRRr
lUhejRrcaniqTK4tkYMHkMVa6dNvKlvhIJpKL7xU8RzJsuB3hQoE5ak4tgSE
+lfgd6LGIcOzM+wPFvF7rvkA+pCOwWbqVJlN8EKAFr/my6ucC8xqMP/B6Zp1
b9ZTGo2j0H5IEYQHp9MSQTl1UkRW/2ykcRPk1x0YFrRYm9zHRoo6MhhKrROP
nQo7UIxIE179WAZOQDdPst0Q6ikaGj9POfoi+aV3JmX1r616aSRwN4b4uPco
RfUDCxUpKdu185DxgfPQ27avqUWlxHD8cZWoe7U/C8HyfyMUhLT+zcl5f3YZ
A4ZZLt8AeqGPaZOtnUQPfFuSsTOnsrlij7QFGAf71bDGovwGjrtIimgqchaS
fS0F4CExhO4QMUr+mRhv3HrcJZEKW13JKLhYNwuAwTP5lDe6Ee/42TG95PBq
yC7nd32mRunjWqszMTMsQ7un7I/TuxjlFLTC6al/zOBGqmPskezj2XBwY2Pm
ab9djx1sFKRB0cxA0xvF0fSuKGPbFpkcxZZj/AxeLiZi89cguQu3hKLcFOCA
Ktr7muN9Y/7brqV2N/0G79HO/Q4FCj1XEmGslRbl3VMvYpe/f2ru3aNshcnC
XBvBIt2045U3NnOLdJoX7lbm9i4bA2fmdhXj4HastF8M/mm7wjuI0gxnhX2V
aFg2g2g0KWwhFCzjmvcqdXkd/0iZ7u42ETSjjjp/qaHA3KnPzRW2iNzLVThb
r7WP1vLZcwz0/aEXWNqYXa6IYd+uDickN2dL7mQ/5ZNloNKeQjq/po3Nbi4N
tCW71HPfJ62up6oJkcqu3EacH47MUhyDczqi12P8nsHjls3SyBBqUeeZx9fF
ENpMLDZ6eYAGTUhCpxUVtsusk5L/n8+S1pgRXXsoqGE9x+MugOojvSbDdCkx
J+hyYizceBIp02MgMEwEa1S51M/IBjMyAmbzmGmtcOX4vhC6p0BNmzML643w
yyLxYh0/c8aJ7fS0N1sOwp+AiClAKAgfcpJ7K4IBo4ajpIsbMhzof6NmzULI
riNLTQKAveH6YuZo70t623jTkXdM5W+3EBWb2Eeg/k1Uf7kkPz0KpOZlgMx/
ApdTUF2olSMlZneNNX7sRkBRa+1w7ADq7Ku24D9tBd+ifKMWzI6wSnWuI6bq
x+/Z1BGhgNjZkgyglDuK2Jey8mwWSWwKKQpr+LAv6fH/9ZEr+/QWMMPn3Nis
6+r1WhQVe0HQfyNs8jCTG7i3MmXuulznXDM3MWaeJHAVb6PnH/jzB2kDCcCP
c2vVl92/wNtw0lc0J0bNbBnLJJEzjNbuaIDAFG2XF0gKP8LLIlhVYv4hflSG
1mK47qDKuOY9nfUjIkffBNYX3Qez9M/HfrNfTKhgQyxza+ZJi6NSaKmOjm30
kuc/K7brcEK25WYa6q5t7qx/bmlr1Z7ZeNDhd1L+3LLfFWQpX2ZXdUqpSRnO
D5w5ofn4Bp8YHhOMFU8yQNaWUDUErhKzDdCb8Wv8u7f89r3wTbSV0hOrga/E
+c8gqFexcx0NC0m9DLkoabzmykB6pHEba6OGDsgjKMEcldLLSDR++7rnscIA
Jblmv8uVLhbR3r0YlEjuRR+vgplkZ6tNWD8OWdjN/DE6rIbTcH8CBlDlfKcr
k9/gxdwNbegCy6kfSYB7c0ZX1qsZI8DgE/vIH3HGYM9NNqbvrt/x5ImF0GG7
2x1btZz8xrni6B0eKGdU5LHqqnixgPjn+0bevsI1Z5dojXHlrFmDRPlQBJAK
uF9v/EnDdJrw72Tjxi03PiqV1rDZ6Bo7qM8rFaUYPJDIsz7jeP+QEQfl5Zjy
X6KvB0SM6HaQcyaw9YbtkwmSymVETA/GdU4AIwSAAWg1MRoDtVMeWDcAq01+
KgNe8CDIDaJr5yAhTLxyuSe3gXPfGsZlSYM91iGOQDLpdDRhnKGkDlhxsuB1
hZPRQ0yu4TVySjXIzed+thcznGSd4bv2De6373zT24yUoLQIuUBF1zpG6fl6
veuA5WVID3eAy1mRGzMSo2P+BpDqBSCM5N3N1tVN0paH/JKiaIKiGGcBYsEK
qZ6BvGEjihJf/v6bHNEXe44pfaCY0Ph+s9Wdfk+waivVSx0Vd6eYjg1el6U2
8s26txEqidYCag8EuzQvQWSgXxtbNG5y5a5pKzIUVB79qH/M/MrVpkgeXXT0
3H+r+jADGa1xITEBm1t21ElTSPMNIM/OAsqwZXXhzRVdH22Nw5jpIrE9EuLo
lX4kZI69RXFYRpO9rvC0h/psG/PVJT6i4rp3rj91OizQ/Cd+l5Kl0ERqKFxE
1wFPA+ew+/5/S5L0o1x8p9EkG3lAbv/7lWXaNkcO53ulHSgdDIGYkf5RyZdf
E0jcafwNPJYqR4puiqa5PejfaQJZ0i92Ai+yGCOzCReSLCrgR1Ju/4NNzf9p
EI0sl5xs/C1ggDdOA6YTLIVntnbUDvIm20UYBXUitpvCOapgL5G8icNT5obv
w7Xpjo4OB6VJuDIhiJk7dkRqAPlNMqvmvN3RvnEfkuROu/1MiMH74/7frf2v
N5Hqp4Pu1PiXNZOQsAO4xDs15ENKDBB/QvcuxzNr/oFHyo6SCZFz/eltnd2n
LPeET9l7ltKMduWFqo0Wb81qRvWxSBlf+3kislxceIwJq4K/jzvdmQIYJFWw
sRv6jbZ97h7ClesIZHFOCA/qtKvNj9vP8E26UM2H6vGg359/deHbdmd4rN3X
VActtIu3GM9/RVzmmPcX3OxfJjq871iv7j62ck8l5iKugQemvoryDNR1vlHN
FYa0Dk/QSr/JC7pUud41QUOSOTVsC99kDdMS6icJwUa6ysD/i/eebYZAPj+x
iTDrBFY1DuyK9W81c111JbhUaDQ9/039/RGGMEwmtzfc/ixbwnI41iXsKYht
G+fahnuxn9O9raanpAocjliaVJZ2qUyRGDIL0Tldvk3pc2HSsip8W3PpcMaF
5cNwCePnrIOS+q8dr53tSOmGAwa/qcBmZKKQex1ArAy5zyeXXK0snukjZduU
2yyguk1amil/43WZxyxo2tQ3ciwwTqObkV1xHXJ3qFs+do2cfYa92HVZeeZa
ye/ep1j36u+w7iCj8IKyaJUzVOx9PQXbK7fXKfaJUQkCwcPlNMm/ar3FFDHO
S0H6OlGkuihE/eZTMsOMbeRP2CPohjkAxfP96h2e960R8AaHfsHOxf4scdMt
MZuao3RgcTLm53Mjj6bemhwognykE/bnBjhQC+Vq6yxEAG/+FrC9ZDSTPKmc
KVx2xbAvQHYbuTt+lxKauS7ItmfNjllA5VbPiTcRurKJFFedBsOA0QoTc/JO
zC7ZhfjM+DRE1gwfWJfwlwb+yUGycXS5q/CHysvAAczrK4e2XXroo+Jq6r32
htJrew43rHM19BUYVlDy5UXFIwl1HVj+ZfUk8DAl0LXP39E19c8ee2gVGIAv
3yxcjnres1SQLZKThwBPIl57FpU7pDUmRjQvOAWRuyvlz4KVGae4iOIGxZCG
oNkOKObJK68TN2EE5nzLFHiG6/Sya/4wnd9bC/DqFNgSYKvkpGKGzeOBlvky
qs1tr9NZddha/NGYUGbITywPVJ6KMi2zOlvnZ5X6vt4uZo55eTL5WkKsNJT3
9K1Ph4qKF1FFv9hWGRMDn33JgodkIMf8tK/fyqm+3Bjj/dGq65J29G1co2xw
3ivm0maPF33AQwZkGntCaKxGcMRWm0xJulhqBwCp1/kB1itDlxXyD6SIXNS9
2U04VS4pYueQZ4K/BPV7BshC/FkyBCT+wKhu5CGa9M5057r6rgQlgv1MvtII
/8UjtBiUhJk/Sj6fB/B5ZhWTPISqq3xtquIrcJFmJOOoyerj/NIxP3tIGBFq
lafrMEmJYj0yMtbb3TNA6fIFhAXJDbmTA8waocGOdz/rv3LLBi7LAEHPwQIq
l7VX+ZoxK/LOCdq7wskZSgZF8ccpfKOvC6Z/giZ+3LxPt1PDMSy7xpca/HZH
tgnRVNHBCanLoG43zYr2XuJxkgguqxnCsfVSVJXN2dLW8MntFBENqs4iUw80
nsw6mOO+pJ8Abw+kRT9hkL349AanPCZf/DnkZxCxdSMhEqhbzceqBVJU7lMC
SvyGFyFMnEqN/WAkRvVmVp6wWMigPh1pUnzJKHeA5UCdSHgS33vSJBvjDw2I
MRfYCDnR2z68p1G1E2osiAqIPkfUPadniIa2A51JT8H7qGvua4fy9ns7Ls0+
3hkT36imuXiUaxihkT8s3QnZVUEwm6CszqgmeRu5iJ9O4121bR0EUoAUslRR
AEPAIgwqMP16k5sBsUouUOOAI7f1dyertofUgyXolbNudh1pEUcNTVGgDJOA
AwWNEyXpOL9M8QDSJKFGNxzc3QL8AXPG3iIwrAduNqq8/Nz1mIkKENlM0yMc
iRVrac+e9rV+1upV68b0zr/vtZW5PbRcgC3CXGaLGUCOMupInVGs1yD4iwll
V/SY/U870XRd9ivDDXA5boWIJ+sKGcEjBjxxqNpVj+A3i4An7DAQ8aT18Aho
XMLYhFErEkIShse4q3PXeLLIGtx+5WesDG1JroOAiUIxu4NXoPN4ROqLH0G+
qnt2SNfnaSAt9z7RIv8JIriP/KvqEt2ZGhg4UsEKtH32GvxGqJuShjvfkeka
TsSh4gWqvRilEtElRJUXHD9fNB/UINuBa6b46kff3ixh8cQH0Cqed1DED1PK
C5iefa2RE9hoq6TFkuj64er9qKvny+IeqS638vUpgmfM8U3y37wCj5B5vJ/h
0lSJSR1kO/43vYScpaZsCj0Gu1nwDON5KbZuRedwx9U+a5c/jvxSQa017fBr
mLu10Vq9II2pWP0cyxTemaFeyHEdi/9d2keLdh0bxcsBhXM2Rmnim59f08AK
Je95OnES+XD8HG1mJhm64POadJSqSFZD9kOFJVasEKkoU6K96WhpENhyIA1o
wg+FySez835vsrbPtlL2n5bi/v8l3E9h6t7wmBPhtqdusLktQlItXxv2rt/r
Eq1yzS396dvkblhGedOnJch/y1bhBlMBi/5X3sJjNtEaM+Ams6DR8tRLSJo4
bySp70wX8dWKmO8HhqcwSg1sR1XaxK7UVfhWzaedRq2GojleICayScFUbnqo
yisdrZGhtYvFM2X3AcgfHmq1cwqETk9FuFmGP6F7vgAVrgWXd2dONWsPgR8T
EYH5P8lGL1ouLBjCGZrOCOKEFa2us7Wb+eR/6PEcV6DezJTRX6ru/ZA2T55+
zDRV9SBcZ39HdomI+w1OXO8yprENZ9Bm1fqmnmysN6VlUzDKRXwmnKGerfwN
8ybUmEXVHlYWYvkT5He3TD4LN0ODd2Ir3C1y76lnGupoZO48A6507kFNxG0M
V+B7iFXnIwn7Ziv685tgPFBNxxkiJYQ40K1rKpB5IXM8+Nvv1DOsoQn/i4LP
v+eY5zohezApvMHxgvuAXPl1NmM0yCEKAUrMkbMMoCJp0fV8GNWlvw17qb69
6yFd/Lvul+hwRAlffLjOyR5BbYu7LAn4+C91Dfn6b2lRw6Hsd3N8hVswDgRW
5TWYlvDbe/jRKHQUGhqdaAfvF5KoVL9khcl//1eEZpbikTZSqqz8nSrvQAeU
iwQ58rCr97+OGdf/YWfci5N1BQVvy9r4KCcxdgm41arrWc1DL4z5lbcqA3Hg
u55YMoGyKiv3oTVpUX5tqq/YWh3+v842hzGuA3F6sfe554FBcomJ3TP/wu+F
4YLX4tuniCpD8W2L+V1safEmDchLuNK5Tv293bi4WE1ds3zcG8JZw+boypl1
fII9IEDujS/3r6sLSNLy5cxBO56uBW60iXj5PL6DF2UNZ81aMw1j4L+VKu+G
aiX/lgZuEgzlwfzG5sYiV67LxDymwlCNKLRjtaVrl5yV+huUV5+asgAASleM
InYay2eLPFwf6Qw3g3qWzjjJns5uw7IKwH7ckjbylrsswVA6uLwNs7OCDX7B
i4Lwsabbas82W2kxykH9gzPX9+qIDmAYj8UujWcR7KSzlQ8N92zPOXmwEYgA
Z5ZYZkWz38BQ/d0AU5y2YksUTbEISLteVlpXwSEawOmWMKe82szBS9vAyOcC
1CUvyDGFXWj9FnODBqUNEnVUTtstkZIstVFiaZ2bl2FgKXlc5w26f/Rl2rIc
nc9XGofpWn67yvfdwG+fGWFnJMRsdGT0niG8AacqLrYwmWEcU4eRwlrHzlC8
UZG84B/8571Xdr1Tk4/MJBRCpq0RoCbjWEocTRAd4kHLuAUXDTYJPdnnL7T9
Wrbv8nt+TbrCVZaDtUSh5Gs9VXHhPe8wkAKyxyjrj+pGa0ry+nT7aqGuXbkT
vxzirDvPhfSKQimQRDeAqRgY4vhG31SG1qAwB/u3g1xodLlg8jFsxfmxyl/m
tCK+QZIqZh99a7TWfuUm2XZGRehY8erA/yLOEJZlNabDuCECXVFSZfCeRICp
6fgzbCqE8yxudMbyhxJfBMBINvbNieLCJM4IzCAQi88Dk1xq11y2ryJ3MINd
uGefJdtSl+cTRp44bRrDWFPYvEOMi0XjtNutKyqfn/LBYk8OKNIu8DfKnz1/
jQ31felC2JqMbn12xqH5WQrIsRURyzghLLXLsNq4z33ahMkv/5UCRFlT860K
1A2ZjEf4Feo+S1zUWCvTLoh5UJlyPe+Ah++VlYjb8LZrwe8p5P0+6KwQ/6+v
EQsa7fbrxagIsK8O/ne7tugW/sIlqow3Tpdoo+9Fg9NWWbTNy8Es4UQkI6Ks
C7zkPWa9cHlSLeC5xlI3alIiAZ8WTCi9KibNdfMXXAY7Ia33f2ALDzV2PjKn
FFsY4QfZroPBWhRo4tXn2RRAQGK3AIbDt0b+NnQVNTBjzgtaim8bm9qev48w
PD/dZrFSL+lEzd+BAt2lejuHRfm4/F3UVI0V7zaczltGIOTTNzYv1n6uLO41
7bWNK6jUoRbfSg52P+FDl4MVa9d+FAJzITGYniW1me9XXHYBRZCvusqtfTZe
u+NdYPgGEZ4HRiBfkovg1O3Hh//M9eYwahOrP9P4XbhiQbW6v54NWwpwH5g1
GPOqa+QaXZs7KljSH7Av1/+WCPpti9gM0nLZ+G8eHoIxdL7b7mTfZRUTtZh8
xO6EmnU1rdAsRBpF1F//ULCOy68m/9U2rqaR2ETCD559qedhNXTqghZMjMkG
LWEP74j47Ovg2srRvOoED+ahxJBVE7We+orfnXJEulN3XKaZhyOWiXsxAnQ2
LoCfvMnmA5SYJeAofW+W7Sh0b6H3nOPlD+Yqf+AcQUhARWkRtYfR02x3kjpv
mYuNnT62MjIK9UGrfFQGWMUSW5ZkcVptr5kc1VXKoOPIUo1edCTCaZxzvXW6
HcA3jfbp1xVMVkt20v0jA5M4UDRmxQ6m9s57F0keu30hajfIoGZc2ApMCJZ7
+8FJROqrjkp/bf9ASmRVuZuWYEkUCfmN5RHQx6k6Zub3ZvQmfA0mpjoOUobF
17kVHeVENISsGiGml9LCZpJiHxhEVA9lFjQcF1wqjA69pNT4Zh7OkfSX3bS2
oZuy8FR57gzW97kS7QV8Kh20MWOe4j/gZGhhuMfZIX7YZsloq8BFok8zHBKO
EH1hXYorqVByMHzjIvpp6EUGa3prf3EaJQEtOkC8fWu4dd6jTj2lvbwsikA/
OLeGPu8IcN5ylMY2dieDDjHi/EG/5A3lOTiGeppmKMwo9IxM/TJFjtwAk/53
+c0Q40ISpaYBd4+etlBUf5A+zmvgH7ilLU6Q+pE0w36Ip7DXpiPpwowMnJ3u
qjr6rllZg77vcsdtBjPSbFe80KMFLkqgfMXFsV1kuG+wlNNr+ho+fsQAdGzd
LDPkRfPaXwEd2I84qur1D1tciSoT51P/2npNEdhOaKpA6ZEbhEwiAyKDvt0v
R9WUaupWODjJxI/pnML9stwVhvZkT8L7IbTBUrdTIA65WtR7nerZSf9jHlf6
2oGNFOoSmWjtk8Auds3GJFDY3MZMDZuQbK1MRsqlw853CwnDmTXKFUUdtYbh
xj/yAvOwJlHm9X6a19GDkbQ3YRjvKhYGusThUeqleDEvYyzqianKwgPqctue
m45yHu2It6vF7OkuU3/ldsDD05rVrPDn6vVFTaB8Lxox90nZZOFIIC2Wtr9z
5f3kfG9dckmbtnogQi64A91ZDlBgHItNQd0kZkJ6FqPICcfRrQut6nlzxwoL
uenwKu0r8hGQ4/M4cAyzAofyuwaHJlD7ORVRcAx6hPs+IukdWbKa8RmXNcgp
DhHJ6tKHG+0wzpXOy720moVOlbAYEm+yrNpeCZQGO2Yd+iidAR12tVR3+kQu
PcLa0hSUGvDM5ULWCooMHzMiD3WuS8W3c7VrQ4Cy1bODHd/yRPnG0T+S/m6p
WwqlK3iDnqvm33A8E1OWh8SiQNTXMbXaFp2GW65XYcVP8zwvpD8xD2CjERTU
Vg+TLuoqjHp7ynyYdU4CfXZUAKqQQGZueKu2ec/Hjx1LwPVsos6WXn6wJx1U
quFtpege8cdPr4MPcgElNhLMNRo/jFUMkrXgyele+QE9MdhYdAlhqso2HGh3
dVFmJBbltY0tTqTapRf2Ohjc/kJNYq2evb+5KS8eJnA8ez1f9bWmarN4any0
+gXrRp9pLqD4oR+vbYEpRI6C6zU3WeIAxrvQxJ8QLJK55LTVGnTdLYHUx+mE
eVqxqUMjbHbpe4FFPWzzw7xl4WAQJ8v5NItxDJsiKXLOQEfzgttERpPq7n8k
yzfhfrlz8sGZEeqG/i8QS7cZoIkLlMEG1tPw5/99rs77TvVFEIco9BticAET
Np0EvxOLbifryhH9TANbuTUu4SxvW+BS1M30BlNqQSGMsy/hz2F2Q3KeyyV1
8PPnlyJX/+JAqbiG9Eh1d5AJwb+H0Tnex2Waabt7r2ZJwoAx9TGuMa1m0f01
S+0y+7EeUZXjs8yuuYC+4QJki7wZYpoJezbwM7z1wAddOWMgcZuSgwStnkZk
7Eiy5eyFkZMAub7JKEirn5WbSbQ7fmmdCsKD36AFrWigfRJUku/8bLFRbsHv
1vQGLx4twVsTMCtNz75mlChwxa495WqDE3BHxwcu1qb8t8xSjMDPRkfvYaQK
+0lTCH5qI0equoaexxUSIMBRzQIzI2lPofZMXINJwm/B+fePM26SOU/GIE8m
WTOb+iA1z75fn/1NJwh/weK6beh4aNOPa46ODyf31x9fKf2OydpYnBNQvOM2
XqIQXE+km5YynCdwAhenYWn8GmjjiXDpjJWtz47AD0+1PVkz+9uBFtptJ/+/
lywRvO/h0xWgMspniwoK6SJXrYhXptgIS+p/MEoG6brinG4C8vWBqKCf86ZN
rmFYwLspklVN/I6ouPwxawtMcWK9pE5lYAOdt8M9OpED+YBLu1D/W001cvuK
O+LvU5sDChWXUd5RfVYiGfb5ElmQZ60SoL5FzVgQqq89bxXUKJ3R99/nURZ0
WMqtjj9tiJ4lrfIJ4gUC9NdPpiCUQvWVbOHjtNk59dWbnOcYL6x46Xd5SQx0
nnj4r/z9mixaOP4PZv4vj3M2wzFsE93uE7haYdW7Jjmd5lmI4KwxUM+URniy
RLtjYVgDpRUWO54Czhj0wShe9+dpOycERGw2OECN3MiGgqhrMpkuKDyk8tir
IivJ4F/w3i9y9JKTgDsKwyc+5lnfglzAQyVhOcHV3Xwr89XNpzSah5a0Va+m
aNstXHKeo8QwOhp4nyZjXDHf51v4/XKb7f2kDs61ZunvRZkN2NOoc0ag3h96
9GjLEDyVR4HSJ5AiokEIsHAVuqhJWa4WjxGYCIFn+3P7dSdZn3JkKXWDcUUT
AsQMfwALTITVXyGlBU57PRxrdw+LlDqV1k5DsqvEQnTq8RJoZQ+7AYkkZIMo
nxUq2EdiZ3wd2b7JeRfeFMm4QBgNejERLF+ZsAIApnBCBPJxANRKfJa7NuJK
NIjh29rm5SM0IL22qGBmDaKD2kCKoXmEHcWN2gOidbJ65/oOyTHG1D66NyvZ
TMbQUw9meYORYHl3XNAU7zegIZ5azlKtoH3Dl3DaNO+htTCnxjr9hIOClO64
NMcLE4urqG29VOoNroyEcNJIbLrijKfYSfe1nvxeDyD/XbbkoEHwo7JFiNo3
6rrwYUVd8COye47bpmSFeat11EKA3vdBPQISk8abgTT8hKn6EFHq6MviJiTN
K+9ajU4JukZ6Bb3O5pyK5kAn4/1yLPXq+uQ3nDrgR4Yexf1JPH7fW6CrvJO0
f4zKpAUIrIF+Ry8sx7NNM6/wQxGsUcFhdVrJtOOqUsD9yWMxQSr790wka0q0
+G48hRiYe4kcCPWYiBPzRS4clSWRpPZOS4iODFFJVM8RD9PW83Pzo9uw+yui
Bg99y91GsgkgAbfdu4a4nCPMf5o9NQgd7ImFb0QMqe5+oCLJeBw8TMRFdmVt
w7cw5AOOGZzhQrRkd7o56yQTUeVXmquuDaTjbuIdFoR1hxERooym515+aYXc
txXy7WRJjyP/Qg+B+jgpcF4STJjbhcqNfhHC6O8CiWtpJFsEysrGiRA6wl/Z
5bE1wEnXNmIcXE4WfN3TdokYoSMta6d2ny/41AYay2ZXNTmTdSqn3mr7k8Jn
6Hm9Sj5Scy+CC6yo1LTCQ2pwIprozWkk71t1/q7wy6FvDjKTQQmG/2z+Xz3B
pa8Zc/eKaPN/2qXp4kLqJXMbQPkUxiRnZqEEFo7jeCGm7ejBuooNQgta9s2k
VLZkTvoEGTRp8pYC93Xktleq5GUTSVV98ectVNpisNpShdptXn/iwkpymvrM
Qiq4LrFTYXvoTYLdje3dM8Ulu45HV1QnN6Lpd1HM2kroC+o/Peu7YKHDslhR
u0OHAJa1j6C6f9uL5yqKVnQBBtKI8Jx8qdh6T9Zq1xMYJxO2hsDrPJEOt6zi
h2Lr8q42IjXaP7lolgP329JexkNS7Z+1b5nRFdHo6um7QQ+zgCTCUsBQiWBM
SoTMQ82KJHSfFtcPApsNaZAwyb0qg+QzKpdvOwdnx0lJTRfFqooKV3oh++Rb
wRwRH/PNmmwI57jei30VM+32tSZ/3NCrbfzBowcEYRTM5kMnC2Kew3RkHeb2
ou1fL2cmoH6CS61q7aTwEzz9gw1syavPCez4G37/nkaYeqShkEbKFJ341Dfd
7Ezs921dX2laV+n32rS8NI+qc64q5b4b1eUen31d/HuJFa3WVgSKrLxPU34e
ZnW1aVpeDnz/jnAzLyI64ue+JV1sRNUF0yqODT5xDp3h+8YEFxNuKCoQpQsx
JlUpvN3D3lLd1J/h65N8WiEO9RdLaGH8rtVqeUJn99HOtjJd9wHL9CwPLWih
q3B2O77qfau3kaH9/fQrfyyJiYtF6nit2/wJbfE0uLlsPMkPKEcYDJh0jOvf
QC4wDyG9MHJMKZATeDvtg4jpGe02o9L/d+NWAu8AVNVVdcbaZc2xRQgZ8bKR
kULZBro8H1dwN3G7Pfdjz/QdtT+Rvr9pLtWkqzJ2qVTHhHFoTw1IGJiaNDv5
aI1zQw+A8Tt+YGUzL83I6n+SZ3jfQH49cvLQcVjqE6N3NHH0kqmjZzeKPUzI
zE2LyIOiuBe1rtj5kqyGxIDE0IeasIzvKhwMfe6G8JOWa46Xx4Xn3HkmrWGa
DM8IUXKYRbWUkPhlKo1SsPGaNzYhQ72WQlJiOsRQWjludLL1juXZGE64rrV4
Y7ib6VyMSMXLGnJl2UONoicsDh9posFuOsHhnsmxFdSMqQm2T2OpSy/P5xN/
LVmFY6VyCbwkFUReaTdcPcM6No2oenHIKXNa3+P6FBjVusmH+EekPO8MUN+O
fNz6mtWlenyAIu4zrVHR/8T20LuH2W9JugCtlNzHVS8Lzdfx8/o8w0GMUBtt
9eu3iLCJeCCNfEOq4uylWmtDscj4IwMSt83JC4y/X+aYAZjdviiUBH6e5h4i
FC7reju50MD04eRRqUYv8MFwRzfvqDnPqVBUMT8h/uY8J6172+uMZGYMMGLI
5BMy52d1rG3ZzorAzlqE+fFvEy+3eCVvMTt/57PcG7rg66xtSDe3rRYIih6E
gCxWVoLIgGox4yTJMKj2AzGwJWA5EETBoLhiCN+mesR1s4HROcnzSDX16LaV
0YpwviSPJYNUvgCFCD49vPhVfFeJCIhGrtzbMRwl1fO1VfMCtdaFhBUbi0nj
SBUwb30aTwdknSxtV2MKkL/MSXFeXo74G/Oiaktu1L1c9UkIqDdYai4UiZ8V
7zWEDbGack4afADrM2f3toXAJ6tjVpCvS3r25h3Exo2KtybwA0LrsLsDHCyG
NTcmc5C38MIcMq4ETYWgwBgtZKE57UulH6nZoiq2XuRErO+uPQu8UoG4WsHy
3lG9xCkWBd1F6xlEmVCOtZpxtSkT9eNIN+8qHoBo8e4y0OJ8SOrbDPIeRvAY
PGBVL1CbG/wtDb7yX2LbsWSM5dadfcH3QQVfS4KZ0kmYI8maEBqP4B+KPxCn
wf2ese7fsgubzWuayeW+cYUrI1L+Ayd90XHdqTuZyhYNXlNv/EcZIxIjopgH
GBu+iV/cM/aHJk2Y9peGAEQagXCWisZWHYOMbVYbPpEQLceGuICjDjx4No51
wMIFjYaR6pviorF6FGEMIyu+5vZXOxlsPe34Ex0Htyjb8+0WlIIiPlLiT1EP
5GR9kcXz9maEVZRagfw5ZcifW6FdSAHdq/FIVJidMw/HLWs9GRlBSYtoSm7C
JMOV4dZpbguDG2yjgzTMHBG6/sTrWjWcvvKQJq61ZlBR1I/CBVj1fald6qIU
anIAvQyJv/flYD/2A//El9YQhomiXoT+z7BkVwerd3k7kuqM9ZYXJNVJ6JjL
IMs0JH+wcQG52pBYrwxerV9Z46nMEqbytAIXqZyR+YtX6b2s1KeHny8ztG4B
NO4HmqhmE8F5aOWOIoOGf38zWDUCN6/F1h3JsNLDYV59bgbKmPeWHKx6Uqly
n+yer8BVXfRIDCo8WIYkqI/22T3CmPp7hqDNCXa25p7NhCxR/5TZJNO8P2mB
Y/b9DrXJdMFCdzioQ+Iw/YPELnwg2rDaM0Kor/zYC2ey77531OosHHPW6Ip/
r2XanZgzC7vtAkazvWjdu6Gm1tk6OZvhJBv/kXdKLSPCgp8bQH3bKP0tq3hl
V7oYXx3XH/tjfW7kZBHPaZSpMdXZj8EttWRrykjAMJG6BazrFjg4+7aldHhL
8rN2lN7enofpdZYc5BK1m2xgY5rryYSFMN602hOqkUztedG95+bG5Nb0o2Xz
hvtxeu05dIZw3LrezxeeZqTvt3Y7MnvEQ3HZeri/VFiodSM/TSUHCg4oADsn
TGch5E8G32I7O+hsPmn8jgjQVnpwovz/G5T/Tu/qVYM1QrnorihJqMBYfkWp
KLEJ/NxpIe+avx3tWNoyXY6Oh3UM4AxtduJB9vRka5zmhJCChyx/Suak84lY
zkiXk9XIu9sdHYz0p5S9HKNOq6DFSCbeaNciCK6x9Qd/SxB5YiiCMGk6VO3c
5r3GR6ukZlXKZF8zFfH3YE7nH5zR9zErC7Q5/BPthWV566qlYd7kDGys415E
sWNTVkaDjvR/hSsYZKPeHoXBhl65JCnDcctHwOBSRoKPBI0Qu0OI7tfovcEl
sI2qiVTlVgZ8ab6DAyz7TBXZUznKBruYc3t13+IVCr/OgPvbJx6VT3QDFOOb
K7C7Rw7UrjQdiHE5V79SJ8EEBGgYOD7dljG1wVhik/G4elwkQ+3UQtQnBWf2
PtVsWnkQL4v3i44p88YDoYjBXKhByVTX6imcrDWpVLGIoRnkNYYjoJN2r6K6
FBDkqa+MdKFQk0ZFtR/WMcbndI+aW0hUKzlgtPRvIsxyflTVYxGE5j0EEM/Q
NjMmgbkyb/O+uzzozeEIzr2R2kL/AU/d5SzrAyfV1iVwucw4O7kVj5OxITQ1
9bClAkoTMYhzVDy48QPpXWufhBVrQwc2HLx8mig9Qd/Cop4tCNbHFvdHMGXb
bHXuIn4xhg9BlGddtrt8RzWuvLSAjKHfI5bXuQ+/XTa3KbTQtNj8PBoMlrS1
Hp/CvonCQJkqak49l8pztrDE9OK0mM3RwiaK+Ngx6qpUrIXCE1ojGEroNfAJ
FabbbOMSeT+VQ2vu6ThNeHp9WtCs3ED2GF4ApNC2P0lehj1poeBKhk0xB+BM
4f/vdkCwQghPfUaXimPKlpoLKw6PKRx9/wa4SDozoSxM97/YmDaUBZLKDIG6
yh0hvZsl7HRiXW6oLitOmRRBHP6FuOUMFzQzu6Cgy0jQ+UVy1olnjLsS3Bt6
BIENbjSS5IV/51ZaHWpjYqSDUFsYhBuG39HCtyUtxXaCwGSiQG8+lXGzOSbS
yzh84xQ7HmLezs8rMOH40wZJlDXeJLCTAendlVCSD3kuSKKWzQFu9MDGyGgM
7IYcH3eULc/EWeao40ASS4aXNKWpdqk1u3azhJG+MVKSox5PI303fbSwXcAc
3oRLFR4OPvOj/jSN1ELOxSX6o8GuFzbchCaJSahrq1fZ8EShFTK5EKfz2F4V
9FaWV2jnC/4qoQNC1zrjPzTUxZnpblnH/9iahkySMZsyQyYpIxobtae2H4WP
M7YDQEoKqX6H4GNeBRm8CtJcVhBGBjNdeukSkc//0ecj/wtUKvmLulv4W4f+
CUL5W+IIyCu/8jCwKFlX7OcVX4aecgHOhbZ2hkuEez/tkt1lRzGzuWmwoW0n
FjU0JmheNuOhMiQk3W+y0Y3vERnaXypodieUvxbRTujjPHVGy1PssK84N78+
G0FopWwz+Y5pL/5HaT54/5CT5u84sBKYkAxwZ8dqZIaft+/YSrKxglJQUQR3
diTZTkbcrkN2LSV7dFUHEOjyTwhJk4s5aY3DS8Q0Kr7X4BwyijGZVnLGQJkO
Qkrg4+cwAJhOh9LYvqCJHtjyKv3rw41gHKGvj+3zgf+HcCGeq+FmU4tOcjPu
Vkx6JcWl/Ygz0mZV/pDW+X27Fz97iIEO7qwqM/giVDj3UpMtymsMHSVlVVal
fnS325Caf73hhntLO59VJiOn2w2QBg5LgOza6bud/S/Gy99doOLwLQ2NGhzh
d/lD7nAR7mgnYF1ruNLnOxVnZNqB0l2V+ylIv3k9+rkLUQeH3c0trentqLTQ
bMZ6mP6kp5ytf1p1iHGY3h421HSy3Ss9oEXuiE3LNcU5xYO7v5UDGivSi9hG
GXlmNMGA9ZElJ+OYWlzUaz3C0uCiB0QImeX4z6+9m6v2QCOg03cVUinsPp9c
G6lwFRR/7XOtl9SBBfEi2B1iNK9IOvm3mCMm0G6fZmR+/SNUt2tF5fMpY7Ap
fp2sioh36z7FSZuM8LZVXrWIZ53pmTh7F2iea8RqUq0VeB0xJzZOk2XkjSih
Ryf062ttoTkWQp1Svu6N41xvlvfnll8K/8hNnz44aH4Jaf0xIsvc2rm6U0CR
NMQRhiYn7WpLzDXy2huxvu3LVssnGc2XbJ2R/cF9hvhY739ty8tLeApTIne4
WbmScRMTuKXPXOK3yrcPa05kT6VKtl1oY/w4je9jdFGOwSJrVsyMEzo3li8K
68MOOUMYiVrTyr2dFAiBlJ3iG8axU0vbh03XOZ+2G/crqSCMNlWPo3nWn6zz
es9jnQqYEStE1m4rwpHMvuNXSlLfPKF3Qz007EZjil7Yw6IY9vLAChvrZxtu
YPy8/SgFulfjU8VWgR81EybfFnZrhy+XKdcaKUkTru3sGylG/DeT1oOlfuur
vmkis84ZK2elhJm9gyVsOLwVJEjRl9YsFuzXvIe4MjQSZDkGPwsJInQtBBt7
e8whLsuFY3PpqiN4OKBMesPzw++g06b4Bse1MZArxIZyYMXdSiNW/KJ8MdoV
Op5tSRoDWOc5DqOD4n+/EQTcf16DC6Er5GuCnomiCSGwLkN87VuZQwBL35+N
UKsat/O4slpyDnftWD3gkkEfyJtP0O6/Jm7xVZI7oX79j3+fqpGSvvzkV7OX
wFGSc6XbP+D391CXjdCzlOYl5b8rdo9n8HRf1jno1wr6xustCzNFhwCDYjAK
oCBut7GantrwDAxsmpBCa1WFJIReQaw/jUzpwz84jcS4kt+wHlhhcbXnIJ/N
Ufo+qTLl/uHHDzpIYN/xnupN1DcZAL4XaWi9UU8aJYepY5etRQG3MuNLzzon
0el7b+L9x7fJbp3MNpuFnZ9GlsUYggUzsXH8KCMT3Zaa1yKbCzXcAlv8bQWg
N1azUSXc6nMFr1oMj2HNZEakHt21w8FYY3vvdGj6D9kv49TsaKeHyUzB2EvA
jCaUyG0KXllzWaXMNgvif5eoensaRSvSF5dq1Hk+FlVxk/R/4ikXcXiiDG0y
m+RtDAJiDzJ4JvJ6EzmyAeZ4mxkwCSTuc3fFgUBWbpK4a/EQu3jSwlJJ1F0e
hBHMVUc2EnUYS6wgeF5JHWMEN8lJm7oelK8+nBP+22aYzggA8W0/wsCxjpj6
ikvlgJk8Z0NlWC+WmLrvVRKSs59Zt1Q846rfrCbZmxC8/7HHzPKakJpwTIDl
tc32VujpE3Es2mNokyg3aWjrNdVUJAT9UIVi5WYvYgvug1IwXx5QeQseNU5L
2/MduwgG4Q30k/mHG8lCuxTqhbeB5q8vctEYwcGB4JTGclIjaf/WIa/B0YKJ
JjnOZk0IVmVPE9kmo14HUjJUFzJXdwSmK/OCX+g0fJJWT8ytksIobJBIX+/4
n7NJ6JQyY1E/qo6Uyas7nPATtb6kpN1mwAQdgEBw9s9Rvu3mdXKTb0zul7JT
wep+DVHECdLsd8nQR9WgRP3JnCSHzq9k5y9cD/sw4yseEV1gyFrCnTJ1XGkx
UyS3xz5KEgSC0/RuLsr3IfzxJui8JQYic1MV4Y0+mKXGk9LvchbIH4CB8XAB
6g2VJTbwBZnlVCOPMFw/RwhF6UrAPbZk9EkHEEYXPp0I2+n3qn61KVn/ILKI
CZqr//YSK5ItZI12cDslFqTYyAHjarQfxd2WbGnAGi6DXO0Lxum8MsdobBGz
cl65Z1Q0JwHpQdXJS2rWYx0qlb7OoZTh/Zin0PW4jPxHz6mE0p3xqPCmG60v
9/H6rW+QP2YaO2FgGRggIHrWsl3Fqs4VgowPr/7dh40E3tRj4Tq1aMMVVzQY
rZ/vmOxXQS/aW5qqj/Joe9lpnqkUwlDJfAuneLtRa375BKt2Q7jI0P4vRfiD
21bVcPIgV81oRITD2opJpnwHIqyNC0jOyv3nUOPw/BCinWGUSuLTpwWCGsRm
MJb7dqSPivdLC0zVCsX7RGILHO1e2AFtGwpcFape2IDQP3ltFzoitCyPyqUA
O4Vvo+rMFp/SQeLvo6v4CcnjP3sRs/YrB/SatjHVgLhI35Cb/tK8BGP/xCK4
YPDJh0kOEYnstBHTQ66zrt3vpjwDh8y989NwC1/uuDZWdWDUu5amV4LmYRNu
hHFLMGyrpTK8TrcbdmLFgcuAMknLqbBXQhm+wEjOCtTQqkQ6rnIKXqLEi4u8
kAVr7A5Kr6mik/Yd7x5zImRZR0M60c820LiQsP8E8cQotYCjlQoBaHqFaP+G
aKyn7HbgDoKai06g4VCrDTbAxIzt3Mew3dhg2MsDgdA8SUG+gSKTGF1/t/cq
VkLYIRzZeb7lDDbvBzKbV3IZjV6CHd1vpKg1PfY2kRBRtVIx/1P7n2jEQPZS
byH+VRP0nsKIqVL4x6d672wPHBUmB4wNnQOWlJLc9zX7LWcgtP/qChw1fb61
pbkq+DcrOLMMUlsC4rAHed4jsC++lA3zMPhePcoyzYR7liBoCyYJPnXSn6GC
EGeGOEImPYYqwnJtfbFRyN/jnIwVBGCZL7vVOv1xPTs3Dk//KbHpTLiMfacb
JAJlPoRQihEZBFsuN69yEoctaX8wkai1lX40BPfoV0S2WNPFxFofOebzjkVo
ApsLyAt4OEre9IyOEiMYP/+mqiU2oSa7KP3eP9wUCZVLWhcGhkFOgvJIAFAd
5D/sCmOhsVrW8ZEfuXgnzayFTWvdbMnv/+3/5OEKNF6xjIKnsXjVDyJWT7r3
lc8B0fy8vJ1YS9XMC1EJopc2mEKfA5R4z808iXsG33QjJr5nJdesfXia6+2y
sJIYordbHZTh31PjHU0DNQSEswS3xfxHnexsqPoF6ah7y+xRdIc7xZNkCjD0
L6I43cVUb9lMvEuasQA5Y5yTweanpd5Zj0aYKH4DY/p4jz1zla5/FsFjdi1v
jvPoGs9dXw6sAXF8Mp8XI4iMEZkRmX5Xzy8YYpXP35ojkjVCln5PUgZ/kH9B
Rl+uIYr5boDRzN9gqs7IFqTCBMiFbQf9FI7hmP8f8aDdkDqDaSSC9zL5VmbE
g3CrrVnc90ZbE63esoHxqLX7elPPRIVCBT+qnP59lqgfKJIFB+5K6XupfJlw
sX+3qHYrpfgdwwi+y8L6szhSRYROjlL8zZ9jkZQ3unlR/jEYQ+pzBOreAnea
mmNkv5ZZLPVIIccCiTDql78cdEULI7h0JLvoZuYSpiyRXKvxolkkvRw3X5Dn
/d/y6Bdk+LMZbVW+TJNo07s6P0+9GE881l8f5paCDK0XbuH8HRfa6n2rV+aF
USX+oFxt+XOsqXjGUPD3361n2HJvzd7RHjM3SfFKOGDwGrDZwd7XWWD8yt5P
wRGIdC2fZ68NbYokGY48hn14dRo3kTP//bdHqiy4a8YVR1gBFmcI4VOnvg1e
qtfcDBJUlOvsOUvGzbV0JyeDu6oOJm4LsYYb0rwvjdAmjFZp0p204Gk07On4
qxsw0kKvxLdwWbyTuhWos7wfAVQOtaPrdHESPXJugd9acPaaiADibs684tQ+
AlgmCw23F6E5K5qKH0gNoyxOIp3qmfdFMvgc2gzqpk3Fh6W6gvXRlf+dPspY
3v5IzyhQ1VNMmK3gNysWbSVYAxEytvZpjJu3Lz/bR3xzoYwUup/LhqZQGc0p
Lf7xj67brZ9/SaZOKgNN7EVULSmCPhh4rU0JsvE+rOr1TfuEqgydJNnfgBqd
OT8JpBAjYhwbQQTExq33hwau+Tbk8DoLXmZTraBDa0h5fYJCm3+onYdGNENU
a2CmUzRhSkD5xggtbAKi97FsNKGaGxVc6marhZmZ7qvmsJPxpCOPjATs2/Db
NvudWFk0VzhP5mDRt7PTS1w7yz2iJNI79ntLmU92CA9M1qBXbj67dqiaKH6d
K8PhVRoI2r0C8WM6lErCoig7CEEgVWCfES42zPmQgD/FhshFodycgR3rsUUD
dXJ0NQfN+vTL27Njyq0LwjknzN3q26ZOua3/8qnF36UxyO9F1AEJA2wek6vN
Q78WxCoz19L6QMHvbkrjnoIyGHt9+A1f7yTEQuMqJN37V/JKI9B6vkHZ7QbE
uS8Lx+ReAspG/XBW6rZ+J9beIH+I9u/lr5VLPk9q6TvHAIF3hOOlACQ+6vqq
UmuJQErPHNctW75Cl1alT4ljYc5cCZX65I2lCLLOSIJujPdGAJryzonVa3Gw
/g5iFUJQUew2rewyQKr7SAmad+OctoC7aR0Zc/j46vsocxcPRwch9RrfWSmO
eEauPcn2tDPWE7ZwiTxzVG09khBdK3E0vWcP1L9Pe0dVgY6v+Z+HciX7ZJd2
C8jyhkXUQJn/oChLgY1GwpP3Tb5p1a0qRrYYPXhEwwKDOnMDq0XAXV77hW9g
Hacp3dohhwG3EQIKtY0xg/h2Cp9h0P1iG+nwFICOyFYl1CFuo96gAP5hMxaX
Vc3JtdtS+H7V8lDns5XmHHDiI0sB6rkSqRNvkVjUu9hgCNSGMxMq91f0Aeia
tTh9efY8+TdRqMqT9VnjVJWI0YRC1gYLN4+fukiElYx151yipXfkdRDeVBV7
zNhlm5GIHHZL3z1yzoy0XHqd6WHfjLakmK/jqCq+mEaXJ1KMV4OPNOq2GpF2
AEPHlsH1kQsZIKoUF4hAxBZjkwajgpXU1WZE3j9Sir4pAQnDpGp3YGZ/NyjG
v1zv6ajBS/1q5XnWPq+4bV1aFrBiJFhAu6oo8TN2JkGZQu7XB/tbzLKKXkp7
VQt+7tO2Bv8WVHbsqV4LMwi19bSFCPA9ZwB+Tftv08xj0/2X+wQUvctdFfU5
uWXMDsfHwYcJvnhVqAARhKTSj6SR+lIfjegMqtdX7GV48+RPtXp6PCKkgGPj
BW7CGcOZIEIhSe8jFdANXmaHUbsXD2e/qwhpvwMi0i14AZA4oqYL1on2v4JP
p6La89lDWzTFQVr7qs0wf0j6UTX/ui0MrTon2cjkk428RNFG7UQVqI7Atjo/
FM0X2kFGlS3/eJn1w3VPOpf5ql0YZZFyreOaMRYABPUWY9f28sPc/UrxWd9y
egZJGyKfmWl2sfIiSXOLleJOJ4jB8qqAmISzTbaZtgKU/DUWl+84zLY/uWJ6
oKsXgrtApr+aewj1GX7dQHmzHaueeYkqtMxPyLwP1EKYB72Tl7gOVk2MCbrO
PplgcrWCTeeSMiUBXTocGnedKUtBsJeuMMaaNsVp0wZO3JjZIyBou5g7ybFm
U+geGw26U4brNYBt9D0DJqBOtvd8jV9jWqytp8o92ZTMqr2OJWQ+Hyu9dwTx
gk7cqk1r3+47e9EhmAUMD6/qH/nTDpMUZgg26c6eT4hNfJ0EB5oyHwuv/aSd
E4CXPPDjfGTQNWQAibwHDlKHYJL6e21UNnoc68BwZkM0wN7AWPrijUwlkv4l
BTZ5Qu4FTAwkCF/4uv/OlEPp0I9iAsfZghc8l6k56qGX4O7gs7XP6p4jWfyU
8xFpe73+3udMU9cNqKHO2l/eT3Dq+fAz2iMmKaQUyVe0R6ABxXPNGPkTpIuQ
5hnuv+bviLUU582WuItVZFyx/I7uf/k6p73230N7VxsMuD1qNp9ZCJIrgfeg
hVkWy51yMLqKmLNNNTeMtejLEMO3/uTFCcqS+2oZ5JssSl2rNsNnaYCOqHeh
0AOveDYz8xKqN2hlvjwRsNqs+IRPmohT/75fKPy0ocXHTgzU/bo1RcLIMEwK
AlMkhYH4M/DEwU2c5dS7UHAgPUVaohkCwxoM3Mss7+dP8austQNQM2d2EyAg
ywfRvJ9Nt8kS9J8GkWarBipJPVmUK/w8dpwKzDZPKDT2oPG+uyYg26fgMfRG
p0fKSHC3tAoIRSSdRPR1956mhdqi88goC7wWQ8hWm35WixFlTCYkTwg2m5MX
2QZE60w4opfGvPR8CK7zv4kAG7otY0UQ3Cta/1mwbajWjW8xyAMrvZ97GFmw
Nv1LGPQ+v0Bz2oAyvWqTTYrjwo4wiyZiI+moqki30h3qSawRbznxSelhj6lp
T5BEM3a1B/puND3zFhx80sTmoWHNXgg3CUf/aGOlaE3Mud4b5gqAMDy6WVNt
j8N5KSXjdqq/XvP6SFJVRPb1r1NOSWseP9e1hs1k2qmYDoBU7DODtmv78Hwt
Mj6gEnMhfsJDqIC9ttOnOw9UwlHdGpcrWnYsHZhSwxSEesp6Ppr78mp7smcx
/f9e8mjri7RtbzrK0y40mHUNQqbEj/YaDXHGt7zMqQoJeHuxH80F3Z+D765F
A6wBm3ijrPblUc7KufeL8Ams8b69jZHN0Si0CfvwQGkcCTDRUVcEqquoZzHE
xDuqL7/ujVDaeFB3TswzyL3zEiIiLSr+It76VKz0SSY4e+a3ujyvK94PVYrN
ZAABj/MujueOB3D+ZTdW0rp6YPmtIvulyL6XI7UWzU8ijJrfBqcTgu9S3+2M
bMU3DbQ6Oy3Msw3t5ObbmxBKZcx7swvd8tni5uhRUjJUbnpzxtaHX3NnBqsH
gkX5kwST0fOOL82ToGa7p5kx/Ge7qwxewsyK+WWnjztdwGONT8wlM+quZa8+
WI9U0B4rtb69/jSCEydkFfLNR+5MC+PTcm5BzrmYBjjt41NP02lAg7wij/NP
3+WJq9uQ2yNa32zU4Nd0PJGz9P15WZFG3vtxpkKgSuTJC4PVKD7kATiw7JUl
/Gwqy1DodHihtDuV4/eqaToXmecJ8VqeBA7ErWHcBG3FgtVy8+b/4MyB3OeA
ETAmvGNKA6bNA9AxM+o3/dNtGCwBrTo4u5I7GSh1Yx8ULvzMwEFjaslqWzqj
TDco75vQrf0PCTl/aOJ+0tu/6wQsfKoSbFxUlOGrGipdC3m9WBhSgQtMXppQ
ukTF4ZbRLIU5kNcRwH/SmwWvy7gdXCvUUDgp4jEiPjw4w7AHH4kcw/HVeKTQ
1WDMicoFnmKV8/0blTBNIw2DOjng+LhaKyXS7YmnaIGWg8wWmi8oboj4BbiT
WQ4UzSX33OP0oIN1b0NTgNq5ZY96VuoPzDBDRqxYSYCbRK+9ukviOVZKFv9b
nrsAmrkOLYF5F2tI0OJSzLenvNtCYezpsRByufzzFIF2VKuwa7GycUQdvypw
Tip6H3RIG8pcxB98vDhbRY0j2QfnYTB57wtrN3scYJNV/EE+B+GkkBexNBUn
6Uk/N75ATilWOg9En5kYcsXbSu4Kiqgp2F2PATC0Rd6d/Pnxcf//SiUZ3uoz
kxhJlFpC8R/TVI4L6dZbBr1KBhX8YztpbJ7X5o38uRzmSiL/0TJE3jrkS5lJ
R8IBgZmeMl/UPp6T9z6y+q9qSTJFkd/z23UtShmNcVhpKhs+Np4eNfQjmwab
iIHGnNAAUvfb5HNOBuBXcCZ6SWBraIDwh5KtJdcOMWJZDTguFlAB1WVVw18H
Yvh/jfA6fHHoHfZqeAKjFoXSFZq7KC1m6a9IgAZac3EbGDMnUJm1z5kyf6W9
prIzbs0jVYdAmgmfT2G4B2eLQlzCtOcHz774C8QLf8ONDjm5veyzBs0zzrI8
Dtb58rcKV+iSFVXg4r9GF6APfIp0VEzsVXdP6QHRsIAm1pEkgK+dGJEPDDsH
0m9xkYJyp5nbjYsiDKu7z2++lgY8j4S1PoQd1NOnenvoWmYf1Zy7K6QLhY9C
w/osFBp426gtd0ygSpxy6OI1q2KLEtiY0Skd3GaeIT5naLay8ulfyQZNe12N
vmWdzGlltg1uVSBxgZ+5QvDKfakV10tfM9oRDkOjX3c8LMeBbw90DlZgAkSY
XtQ/YG1D5hqz7cpDmAW3HG+XVLce2UPNbLc3NMVVLBztN6voZjYR/obgMH4d
r0Kksvuh+P1pwfvwIGAxtLnm9A1dDN56y1rSy2+BGlg9HISoVKoCHImyilnX
I9Cfv7zCo7hbWddi6X6odhdEuZ9LzwJiSjs64GeoVrLrWpU/OmuUxytAOwOF
Mm9tYURUOrnh4m8w+aPUxiY4GPvrCX9kM17RlyXc2npkyse1AsiV37P53Rrc
nZQmbKrpbW6k5aCvf931N0ExKqKk2NduOBX6AYvvKexZiEghQwsRTmE9/Rn/
U4CQeevsyOtwdK2BZ6Dxvqv62ZEpwdwD4etPCz2hmIqdzRvufl4pkQJx2xzf
UtZ1pZQdsJ78hjI8OKarIuJo6XWNRL7mjkCWbc2ODsMy5a+lj/Qqf+iHbf2X
5ZaOHtW5B1YqyrnrioNX2Jhy+j0TQBbJbaf7YkxUUgMAwhHP/e4LAoSzFcP7
UalaNkpAv5fE9xbrfoR8oD24R+DxQx5XQzWz6aREd/otP2N6/e/VOvG7tBnm
5kBETYhFUjAaojQG6qx/pQgDSlGhKbA7evM12R6OUq5C/zauME/qdXv7Gsft
Y74B3U4JCpjF443rqTQZgAL0XDZBAhLLts2UR0sRjHjD79ezCD1hUu8+pcL1
+2weOu7m+IOHuK8d/EtuMsb8/EtJ0JUkjVxLG7yX0cY1v7vUxoydpM5w3LcJ
PA+n201pDwPb3ZdU8QPDtUN4zOe4Go2Pvc3zs+Kve2F4B1pyP8xr3V1T6w+5
9p/KyuY1WFVrPX/QutWw0yGbFJhCvmxHxMnEoRwHLbnPakIvDZ+r4MXbSWL8
PAAX7mONOZwLKeUhKQ1EVuCb2u4W6PrLate0uAmF+QCNH/Ilb1E718zScqr7
YaSRJMvhScTbjC9GQtYOjA2Z9mfCOU75sFa9JlOlSCUPT8lVLRE2G+Es1+A6
E/rPRd4HPiE/bkD4MZaPGuHDXoRLniGouvvBKN7upfqGIjOZFArviPKTHZEh
eacWcgTswiB8ZxyckEGyInFPswjI39Ci6JmS+H7PU3nvgw/klsg9eoRc/nCV
DQdzro0HvmK1s8aeHoiLJZt5jw2Z63H68DY0Dm88dg/XE4c5e1GxMnLkckmt
f/Ej1Zf8IRs3+wVXhmsyq3yx9/41wQKTliiEDUKe60hK/Xpj9/G6YSfCtVfO
Gr2uiYQt0Xs5Zr+Zx8okUm6hN/oMNMDnmq+bHH7TwDm93Bn88lMSZakEScM+
o1SsKcplX2LvmNDhoOT66R+jD++ElxxwxIg2TcR8sVIAloJ6J/+eZ2lvp215
Edy7RTnoZw8DydmKGUeqHaJIuUAwyFOF/dvMG8z5S3PbEdSkBtisiOLundaE
skjoIkX7fVCRougxNm8O+UrE0dJoXq+AKj2lpPu/25XzhFw4IguubI8Pg/gL
SUvxVJmW86+mS0a7Uo0S4Sg6DdS4J82NXnmyMHvrnRf8zxPEuBtiyDTjwtQ4
qtHT3AZJEiDqjeTBd6PWjFSsyGhGzqsb2OGTRDzOkxl22PIrD8xca2abybTX
Ro4ZsJbmjByySW7A8+m7tgE2ciAUBtDgWqtvwNkNNSeTn81PYYjeDPcoKwef
x42le2WJdhX0yNELpKk8KQnKiN4znHORfWenY1G1l2yjbyqfez9udIuThzrk
UviOUHjd6rci61Drd6xJ5fTSIqx+KqM+LL/CQAjb4RZ7waqPWxZqVAW13rLt
wYv7hzoonG/H55THUIg1jgj58RcTDvNhgTdS5Vi26evA/hKUxjmSMsEe0lGh
r/MvKEGgaVZGU0PZaWHL+BJ3R6x7jcGRMaJsruz6DFCsnFWXeFlomw0nXoXd
Vp/bVKJt4QaMIEvZcHeFQ4n50INE0oCBI8Ljt1xU8CUimvvyrQLI9R86fTT8
rYcAu3ThTDn+fpTCfpIdsWUHI4zkJhMzsUJ/LdZ6otG43GQEDGlCLgY/CzB8
ahDl4GqZt5TQtRsq5l5um+3yxNwG4QvHRjkFk5Yonlkk3cp13OjPePHwb7uY
htE35lOIEjS2Ujf2BqqjTeMFeI9LxHKXe1XOAY35Uy1XTJ5czv4tF0oS2cYF
flw1tFF64n8WRJU3PKMukGNj+WuixPe6+G8s7LdwyuPCYcJMnplWWpj1Ggxo
TZFLfp3S0CI9DEhe5QC9J2ykOppT9vpBGT0JCzyNJaabULNXfV5aYq+R0DS4
iCW6rna+zza8mGBdo4QXPkmCOq4yGVF0Ru27xrBP4wvRlaHgzZ8xA8ok8+hC
kwgxwnE0c9BLaxYgMV9VVU5c26d9bD7boXPPsAYFq0qlWYmOA7pIbdejzaxx
nkGrI2aXTpoXa6Tq6slzzzO8iUQr3eUH9l50k7AQUix6eRB6vXlY9+uvu4yT
V/gouh9g05irgTAxOjfkbNkRrF2JBviytuoKYU5oOkJQVyDGl9HBXHgciJ3j
svU2AwP2abS9mnf1LPyVEU+7pd/WxMk+QZh0BdsdQvauWDPuDOqew1gfvpKw
PBz25cd8piIdxzDCcwwzXkDJpLR0Q6G/ByFxIRKcvAtfdBXqASJW2o2WEfq8
pmiKsJgqBiB/YbER9MHzZHBMlN5ORuzedbvkTVjJ4f5IVRd0QpAY9pthGx7t
bBKXU419Cl155NrmMcN9dQqr2JSii1k03daCb+re+cxv/etV7BpRM7nWoQJK
h3guWaLU+crCy4yZwze6mAzQnBqq9u/ohXUudgEJGOtkgX7vKMqR/T76wbmd
3DUF80Hc4k+CGyx2rr4C3B1+vZDmYbxKk+H+DfVjBe0U2cQhSp35AmRVzhDs
ytpEy3nR72s6eGSnIs/2bjpIfbpatgmjQAUOt4a6NBq3p0gK4D0h2J3OAtdk
crQIBFP7audUVlN0Bdisr1mwEHnzxegsC/tAxsGUnZlXvxFmBuXUk9GXx0nR
LnToJpKyDF51Jwy8uyDxlUr3GCuiQ7cHrXU/6DYGD1uJRi3QHBXuBKlh9jnq
wnCVuHv4UPk59Y4pRwlFxLPEODHNjpQa/Rbgnb4iv1Ci127OSL/ZU076GU+W
HaimsB3Vd40ilIbjCM0/bzMOIHqkSpba/+wAOll1ZuGf+LSzrF0Ix9Sfjt6U
dldSRVTY4MApu44N8+95JPkGlYnn+t/ZPBit7MoZZ2wbfZogMyLiA6rjJ49J
niyc8jAO/H4KFK8kW0MFIDFIzuRHYpwsFv13TJFBZF3hoDr8dGgEu0Z7bHRv
Z6C47mLvYq/mw4V8/DUwSNobOMX1xQ2lmrN6bBP9u+3WwfsVIAtkQR4i1iF3
Dr/4SH4R6ZC92Hn2fcOLarZViYmlEkBq2NvgzDL4wqJ2ArPMvcKz8sVg0k+S
zfJkgXEXTJiQDRe/PbAjYamWSdQGM38l5HQnthjtM9bSme8xDbQWLk0+vGB1
fz2fQLkE5ixCITGDPDeGEyTJAi8/f2SjwuQU+MutttDT13wDEpmchy0SJDdX
qtcALz6S7dvitDRdNJGsLQ7Jh0KvQCMov5WCCFSEAUXw3zmVDV0lp+0WiaQ8
F+uFacOZXvy6/0CgcnoXMqFc2t9EwVXSfYiuIUPHaRqh7ifT2BXtFY6uoZ9V
+E6TfXallg+REtzJVdY36owoWORnkSUaTwNQdNW8zvNs5y23yiweptkXHp1D
bMELs8USopwjiMMga5imvaJpboMN9y26zZn2r2e6znC2V3W9AMcYvTM86CaT
8FezvD3hI5KLFhjAJp5TpM00nM+75UABTVy0z5HUPXVGyP/BKz/Rc7/xRqfJ
faTdUIIZMJmjauMa9PVdDU3Pko3uLCpuL76/uKYZZNkFyqDzUfYhGDnAfMt5
4D83fyLpgZndyPzlOhPwXvTtCgMNhbfprh0Cev2cxx9r2zeD2SoWFELr/EGn
BvhYqvmLabX6OwiiSxN5Lv2eKwHyBPKHT6lLLI0nP95faxQJKdldpenwg6Cp
62hyqLObrhA87hMJan0g0O0+ICcb5scJTUse3LTfeNhQjSFpYwPTIdcx1ui9
N0xlNAf8+j+nUPOirqVCD6CcwpZ65nATz3Q37ijp6Tnq47VYo0NbcaFODfl0
yEmIdBKfIAOh/IfbY16ahULkw0m0xP3LW12Bzs1Wcz+O9N6QWZhfkolpfN4K
4v6snb+WBHCDnUvzVQnHq11AZhgSlm1rG8QGHtAaEV5pfL9S7xvubPnEiHZh
1DibOPzj86PqnSh3Ncn78AiUOFTOv9XpJhIVlKP/+dACFEAs1FftC6jWzNEr
MKy7b+i2WXaOD5sUwqFp99lILOjzs4q7CxF1dsJA+NrVlCYqBVIq7SLZn0xP
mmBAki7Hfww2JVZYanLtnL6c3es4yD4ZHKL6uJetP5FZ3zuONNnToM39tZ8J
HpBZ640bVpTdlPajWKFkLCvaaZ/KbNtoGNx7iaAGR/IQDnMxU5UXvaPvf8qw
uBTD1xa35w/IZi2yt5sCPeoytYhPlKyC7gfOvpsRS/1wMD0sWO676aclNss9
O0qoqw8iy48JzBI/TArX01DRl552bLNzTn7ddOy/o6ji5907r3xEs8aLVEg0
w1bFgtkl3uRoX+hZXGIEaHoEAwZnX/F3HwonCW5sDgkl/XHACdl9vL3+wkMR
JpUCXMLCo8/0n5aG2Y8lav5l2Zhk8PUOgHt+Z09goEH31yDJwGCDULnBFRgp
HEVVeJKrac68rmvTn8Mv4h7tPqbrCdiNKtzJkAGFdCicmQ+d3zCHkHWpQ/Ol
XGIWSaFcMsPWczPq97iZ8xR+wDeIxAp8XNnYDQI/vbS207UDq4nmRiWjKCbE
5xrkxCeFuQr1QFP56PwxnvyQ3mPLEfdejL9Z+qtqQ+Gwp1unPYJXQMKN+FSl
9hAqUnD3ahWoga6wPVYOzsiw1/xsR+vZG5Epai9YtGuOmaFdwHXHbe0ptGLo
E+QSOO8oa2XaEKlpIBvh7YylUpPTDL6oBxRLzcJq10098EBw7rW+PeIs6CfO
iPCky0/tOc5WDolDfwG54Kg2NiEiHjTNOMI0wFsKphjgjt6F/wk6kbNo2d7o
ocsSA9n/IUYIQg4fwhJ5pbdJEB954i2dbMg/zcMOT1b9iiwMY+q4TmJmiWVB
F7vzPbZ1dXJscgKs3NWMWM/E6JBdNrNPS3UPCPBXAFiFZpxhK8WS36X4esyk
xulWTGwQh31TpVvkkjalqS0xJityVRsZH66hxi+oAmU6/nYZ93D5McPT+OiD
7KJliuk/dxSXuWM0fPPxRazlY0XSEKzhnxqp/Llk1/HLGPZ295w0+QLiZbP2
e7t5aFUP55xw0soqjPZTTf4Rzvn667NgX3eIh0KIoFPERXXKVvwV5m73Ki0M
gedbkhm6Y5PUx/NGi6MRPhk+VEouJZ/yDQdfSHw6vwo1xduMfsv/BTLlVou8
tRP0EhRXr1/G6iph2nBZ1TaU/neEPp2ZlHzbbxwXPeohn4EiQhhbX3oVEdLJ
2/VSVkPXUEjclDdbUzhgUxOtHk01jmuFDIfXlVw0LI9+o0dcYSrgD4aSKHmX
jdo91UO06t/5Y5goXvHCWr3mxY2XRSdBP2QNSfVTtqCyXbBlpp+7fOF27kwr
F5k/1qwr30AnXzgSGdBVJOZ9U4LsyiBug6ZH2ThJGbi8yHG0nXDKiDw1ITEt
F8AckEYgQuObJDDjHT0vakK02kqrSZ/QVJcbnhjzFbcqFApAbhl4c59vAFSI
idMaXtLG2fEkVy57NyCxRcZD1yZGgDJYo1rNaAKEQy8rl7OnPS1heV5SvCL1
CkKPq9V0aCdqNh+w9x8lofrQNGEHC4FUUHXUL7dcqxDo0DM98yyObxL1QL+p
/y9W7Saz8ymtz/TuE43KDtHxD8dHQbMhwWn0VLAmr7nfSI9jZizMAcJ29VkP
maeJVFW6nnT2z7VhZak1w6zrJzrBwQf7M84zTsQqo04QYL8L00lUzVmwtC/0
5PO9l3mbw4DF6wq8eSCGwx09heEJO/CuZ8d/DZOgG9tlvuiNnKGXGRCw4Drv
xZ97Qikwg/oeBlgdNR1Y1ZefR9tmZx/5Mk8WDkr8djt5ff+YsQ7MvAutJcb2
whahtRm3iBoXY0dIrtVdfBwvyCeHQyYRwYtWssR872BEd44c77D6YsLhBzDJ
v1pk6HG7VaDNI2W70XUtQ3WoGDjn6FXzDZSv4N1w2XyxbjHKImp88RMTj8hp
a7+l0qNvLlUy4QA5apdLPJfE+X5SnSeG2l4IP1WDFkTBINfOb932FmHt5PSk
3aAa9L+nmsdZL0cg00kOGz/Lqw6HQGy8JQk1fljZE1/7ggyjna7eU4QKYaQj
PhdmbuTCIlHCrMTI3RrtIqOur+8yuHu5u4JvZGZ15eaOLXyLfyb0Rsu3Mn54
kwPRpvVZ94gmOtIOmbYwOrkPraWWkd7dcAJjztJ3ARqvl0qSxIQ/IQWtWOnq
llkItAsmgBPXjj3cg5IsTImitwkx2ZmrMh5VK6LJ7XFJfX9inwOCj3gIZcfu
Y8sZZnYggL7zTb6TtrSAPLTqgxOq9o9ySuSqU4b+ax0MWaqzVVTPZhZNk5zy
ehf81ycwlshKiDCJzMxHJy6LK2tsFRnMYD5AsZ0FknGbi/+J98vON0xib3/L
6r05zJlH6tDIPr0Uu4CdfUC+V/XBc8nyV22RpGjLJyRSuDCawlh6q/crCg/9
RJG/SE4P4xlcJLjeh288Tq92dmHtVSykvheEzg0zlBgsyHb+QRM+/Lgx+Fzp
Ppe6YliqOHukx2YOx5GoDcSI9cgVBJ1Upmbfag8/rMg98s/49/w4WkMOYRDY
yAeG5FVMUdvgxGMu14sJhRC5ZJ+iPoHO+dnvbI9uTKiyAgs60Bn6TlXuYMt7
YRcR6I32q5GOMyPTLa5A/foiTvr77Kj9ErNs5T28uzTZElFxO0Vl1aDO9C83
pupSruChDSTbtGE0pODEe7L+EeH8ceGXrwebI12ESZlCon3ofJZDMWqjCS/Z
XHUpJ+EYYiVQzS/a3t3zb/m4AKngihFpQayDIlrWycZ4nWT5v71iZd0kETba
ivpG41QZVeCFl45hMFqzeJJJwYh8rH8Oq/m4a7FpO3mF/4DQrVka3JdQ0HEl
/30XfiwxPaeszFqYsC49nO6RM5J8D/xE83iGFFN4+rJ1SITGd6UJgQwvKpVe
aezf+J5qaKv/rgS/wczhNZzg2xsipQmlrcs5k6m+2YJuN7UW4l2PAmbZDcJW
ht3UQFvGgQrybfAu4gUwU69B88BI7jGsXHBqwNcjbSh4xZwq5Y6WCK9zLC9/
UtRnUKG5qLNybLNBDjZ0yilmqT14EtDsjWW2D7sAivlQhsvLZlRQTYhtlyAz
asOxLcEc9xyeUs7Mgpq9Pl6odpNd6WTBpoxhCOaVJwNQOMj2oeMROBwQpKrq
Z1MeU5t+s1npwTE4MK9RNQ4gQElnq54Us8hdoWY2OhdMREMfGVJA/rjCyceC
SmNaj6i0IWxGaLPsbwv6SX4KmAfuR3vOH7PxQ+zrvGrE5vUcGQ+Vo+msMu3S
pk7DRA9LG6p+h0OisWoAixMItYLiVAD6RYEj8DRBs9PN2D0lVKCPTZqzI2ZI
yzeuwxia+Wr3m3d2oKVFdKHnsDIbYmdANwCkhLx5IK5AIgdo+DAp1e5LA7lP
4NRI7vBTYto9jI6OqfrSeXa4qfL6CdLL+lBpYwaeTe03u1eJPko2+HjIZ0cP
rFaIPfQ8IcbQwQ/G+VVBari29YOR1uB3iCx4O6HmdeCxCfNw5O/UPTzZk4g/
sSETP1UMffFgpYhhyUWH81a/jro3y66fPsFjjqGCR5rt02JcunljAnD86uu5
38yOWcX68NIWmlWBHSae5wazUMh5yrDl/FF6DaJx/+6Gv/sQHvZKt7SpT3kE
HTXSmjgP1mqHrEW3qCRqnI7hHKVpaG2S8myzKzRI7rG368x0PQp0rg8//6SW
NP+VZs8iv0uy2TcW4jB2yf9pCRHEdfvxYG7AzEj+5pOn1HZEv+s+vik/BRu0
sOqDYzZNuJUyojJVdBtohvJJzPrvFCS6cTPuGZYEXXkQZrpGkT4YvK0peiYk
5IZ5oCE3/GfJMi1ju0oZaYhrGX862OgAgj6QTWA8iQNGYrP/hzraPp2VmvsE
r1btvHiMnQNP8Z2FHf0nned6981+sjXRqMoi7bJ+0iDr/ike/aNSIxtM8PNi
wKRizYKgIWSMgt4K12mBDGegTc3yj9ImIFTJpa1kVrNLYcyYeKXZhrAZqEnl
T8fE03HaG/4gAwIelNS91XA7P5XaJChdra2zI/NWVKVlKvnLeoHjg1PH67dm
6njkQ6rlsNBAsMj4HUS2vu9ltt8qxQUs+dpVbhNaXhhQmU/23cvr8FzPxKYP
Z6OhoQYp2hJi+Vl6GXiYCzgOGJR+HrrUa1mFXAGgT0olLFRESJOU3F1AQn7d
Fm9nKRouMsHxaGsysve0YrDBDei8HuNlTouBX1mI60xAW2HTizQY1FdLsRm2
+ZdrIVp/Ru4NptP4HATJiAObAZQCSXi2D6vp3OBy+Es4jGet+gB+R240dyjM
AoQbk8YF+gMrzbx9Xkl9Ot8MZ2eYP94qUuhlUaA1n9OQvBBGnUAoexuTl4GP
TFURBDRNbQ5yVQAsErGqID8hslz6G+djwnfc5Yow3gTKYhDj9OR26zckF4OV
wxZEsK0/K4DdI0D9gsn+OpOivgkN2Rvd+UTquvG45ybp+l8zpM7KgHIG8FSL
FV6RD/Va6FywD89XE8fQ9Zyk3cyGEjtlfs4qloS753VW58iKKXfRa18DLH7G
cBO3ckHJtr5wZ4t+6xb/WbcTSvm9IX3C8Pj4zDxMnC8MHhfK6vVVYvIgJhY1
MWH4NQxI1gleUAHQ5Q6IlCZ5WZn3HRG/+cwPgkHLVHyFhX3r5F5wCVTnfJgR
QtbN7vYKKUyscfBPd8C2sXoumcke6vbo5RgL65JIAIZu+eZRYWk4cDHowQoU
hBayXc/tGaWc130s05geGAOn7f0T/Z+YwhbRTA7pYeW/BBepXi9WXGOHyBNk
c2+6Kd3aYfNO7JPNId6bykBw94i9hK1thC14ckfbTH1abcShbmA506Rka126
d8kwHGxrlTQTsWC7Dxt12sXEoOqs0HVgZtihslTjvlgNoV5/eHQPCt6z/34n
LkeTNepfqKsvV7U9ls5lQyW8StKvsnyEf7mz0lwfIoBzpkIxnSuBOXY1Fczw
DXs2WWoNe80O4eATcGfGHAP/stuOyWo7gy3kxuDMa44LdpiWpOmW8T1qOYXk
DitKtaf5ylt6rDH5tOXCx71+Y7OgVhs9hhVOM731XkbWwat0XM+9dboblS1d
VMb1THYvv6DRBwR9H7nNBJh7hcyt1VYYPwAwSIlVJn5HFc4W0koxmj9yXwWL
sdGbkOgkEmvTPlHNlJptXjpnVYWXdRvYiScssRxR1BevXrQBEy7S6yKO4QPM
Kgna8/6/TG4RlCEQgF5ib87Tvdunwx0cF6PK/4voX9SZsSze6C8DbborqAzO
cb7OdY6eE3pV7U8If6F9/q2iP+jvotLctOzYUplSzlhuEF8y89mAtGmQ04hd
zNmk4BlbReXkc4Tt3yXFsjv85jFif4l3tY16+XR+qVgD0G6aIEhVzEIo4iOq
05J/div+ucZAlYbAxRABBFU/60K2oYp+xHovoqkZLNWlwlxw67tpnJyHRO8E
OUPZ81TfSUWtK386lmgCeYvXGmNUUxwO0lJfsNXIUOUZ8AQwl6VxwcmvPtXr
l7Z/CHai12UG55HqlO5liJ/LhIncLIKtQom//OqAtjMXHA97CaVTcow6Fl9B
1wsq9s9sLWItzzOW3EyGPH7WdrUwJLHcUhlCKJdPZm6U1uMi7pbRdXd9SGi/
/n4Zs/n6a28qnVP/umsDHPUW1g5oHkbeBnLx6POUpp5wt3ZHs1BFNy+TaUBg
uc0RS7vhceZ86bV3qysD6LWVewLrSjLYgAi3YqXIt7tGaMnpF3iS9m65b72a
LfCjrselayO76ZPp8ORxGyOT8Y020K0u7G/fXl+e5MloK0onP6iV5e968B/1
9uXdHdLmAwHv+Ho6bqg0sWxVxHC+/SwIfcY+Umuevf/Hg0T3ut2gKNhnFY+W
/du//2s4uE0L6frieEZWfsaD0XxgOMY15jeBu4mAzicufA7+tzWlp+tiBqZ+
V1fQV3mzov2pSnI61maPs4WLcpUQpzlfX/L+pRBaDDeQqlFabWUbfx+pzQP1
8OwsbWvIjW0dsGdwi0Zb5uxqfDbUKneE/Z3IXVwco3+fWjG4clTCItqWCh/o
D+Alg3315FxVAshc6u5RhiKzm1KoN3ks8k+0MwMeEhq752o8GHb8lnI299pS
0o0r8rGGnONxAjMRbvivRyKy3mYbr7d8TEdCwHrB1dMpgvTTxCpvJFf5luL4
U9H9qTf4n/M28Wf0b99e3EYOoEHN6AW11qGc1gX1sCs4yxjJRGBUxhp+eBYN
966TD5le4L6JXJagNc+Up2sGtj3hS4VbWMGwUogjFZIekCkpNv6DRnfQCNc9
3OSYs3rYjwavgtqn3vmAcB4Sc1n7TFuycI/In42hW+tEmdrt+6/gTDBANKVd
rmV6BDjndlyV1vSeqEbr3t/h1PcCPlPJOBpFkSm0dtiSRI/yVAA1pqHBPZAv
P1fhqTLBBcapCiYsR96FatSM/JeNsmEu1gXPimdS0Vnl6yLyry8dG/tV0N8D
KWpgoLwDe7zy3WSERNiuEaIoUIzj0La11Zv3AyVO/WahoXk2IqexIwU+1SMU
VmXOptEZj1v4riLvUVQg3kMMLxFR4E95L8Gt+k5ImO5tT6rKaQNuROxq7QHs
CMiFYc4uHUVOpVfci/p0ElffCa/1SnLDvelGFALptpYAfYw0yrsnFMvWlTYA
s/xwiVJf9kUilp8LqfIuLNSRPzjNMxQE0JYAtOA7w9ybPWmGlOUHYc0SYLVD
rDN1+1i4YPnCWgoE2EYfZfiIXZyNX6ITSeuWYDYXbCBgPbbf3tAUwOfwJ6yc
oaZKLxB1TUTFAzVwgBnpv6kdFl6cw/rpkbh0Ct81AVeTp190bdRdDX0ADvy0
XGidoL5pm9I1cfDD4ias25Xxs86ElCt0pdzTsG9pP8Ell0EKMoXwIPJlkMBq
88GdMrOhrt2KYm2aBvLcKp4WNs1+fBeNdIu5oR/z2jnhQsS7eICjYo5DdlW7
iA6+GKtz4a1mwg8yvxOgMK6DO+WkK7hzJuhYLo8E9pjJIDx3h0RCWFZqZu4O
JGutc2rUoRHcwMJQFViTsg4j0xi8IYq/+32diKn4Wjvx7RCSdd+0V4DWs2vF
6M17pWdZK4tbSdA+BwsQrG+TRXGII6iosT2igkxJHFvSDL0P24+a2CsPV1As
VEwWOR9tFWxat/rLvFitKy5avGtuee5mJVhiJApt8yl+jY0MbpTSr/AyJypN
5Qgr/9x75jMzrVvXfeky1DlijlGanBgi0Hg7jEsrlZcpAvbSTy9jlUcMK+1Y
PqNJPaHLe/PXB2KepU+seCw6cD+85BOOvM8r8Zb5hHUhrTVXXE4MupalOze1
bo66A4UIIUV2gZj8Ai8DcSI2fa/YRzwwSYfOJgVCu+z0Mh1NOB425tk7LiPx
NHQ73CZgvdYTlRaqPXaoD5iSkmEUy8xvRUkIwvXHwQLnYgSjXXM4itmxOSQ5
YWuRsD/xRPih37RI7gIbchHtKoLMtJ8ARg/X6XfT6J56OQY+q3eant1Qnx9K
v4TDUJVSI9IAu+lbufYzbQiYZy2myAnV2w7M/7i6DTwMzpHBkvtPD96L8J35
c93eA3bIj8lV1r6PTinNCoGX3+LzrcntJlI1iYEJhcTp71BIMXwvdXBDAMBE
UIYlLyx4sgy7lj7bJ5A5JGCJ3ew9AhW47BMQNQbfO4xibNJAYrrmqPFcTNSl
siekWHT/disX6fzTncM4DSuQSuJ19szcV3oU9sOt6alitOkbXGu4lgCnXCpN
ytIbzvvHXnN+Pa6bSHLb9+h3TingOuZlG/4eV8FYbLEFvwERbDN6IljqA3qx
68Qttu2jNUdKJ6dXV0Aef1IJem1UqGhAYOdZUfNIWsFqjmWn/Zg+QDzV7BT7
RShnksf+5uzTuE+hol2JES3TeM9zHH18+EDx9KchxygsemIQOzvCFADL8w/y
XWRyzleNiCC5e7gOW1xnx7j5/r+Ib2YtZHBEQMkcVS6q1YwhQ3UZm0iuWVzx
ETigjD6yZ86zSbcTyRIzW3cUf+RylNc4wv3doVELNpxisaSaok6XqOGKTh9R
blY85j0ndPC2o4x/B9njpLLJT8xYWZvoDqxWe12BM97CrxQKio55j3SADb7K
z2worgFONieR6SJ/Rd0Zk9R3qOQgnsxnwhaYk/SqWEpvgOvwiKc3DhsiUVgJ
8b2nFTf+wIkuqDSAt6eNgyX4TiGGg3E1TAKbrJ+BGNo/7Qars0DAp0UkFwCN
rIDepXBOQhcVAki3/1bC9mfQ12H0VNxsgAMRisCb9uQJ0cWy5XURMU0lQwIR
8UnKMB5wq656jxVE5lwbalbsYN7jLvifR629c2v0kBAWzsZCy79xMRYgbTE6
x//SDpnMCMUKw55opa4xnTmI1FPDR5wPOax8jGqePnPsjNr8t/v60QO23LVE
rmHWmonLcnMgH94gCcq0GlWjhIdJEunE884LR/OaZg7zNO1dAn81NEzzWVxF
STbAU/MnXFX41vREmpgYAqmwNlbN9owgTbWY+vgvcUMCAhso/lJh+snWUi0u
o9vj5Aqy22UJg9zsG1IZvpxEZwC25mFD0ThFtN4zTBlksEWgMx2utkOJs53q
KosaL5lnxm8effGq/SaONX7Mg+uIAS6wjlifC0kTjCHdOTjs3RLXPfDI+IS3
+Dhk17JRNNfxtOzMd1O0ZRuOiNKGp1htjD+gBThy1RQAKX+oNpTE/UOJtwwq
yJrFDZXZkQvI8hSCLkQj4VJcxi4J54VjANpJYRMM258AF8rjwnvjVuphgVkT
7dJNxqwzSiDlC5X3u4urLl2qN6tKL36my0xunEy2aUqSD57NVHxygeLsjgx1
S4UEhuQv+r5hWbWies0g0gp2OoeHPfJxEtPG3tqMT5slBERlvXmLEeSyHSKu
gO995f3Vjq0rAR4yCTqKCaS3ihjvrnHXsrkdeg9FhGCuMiAHoJ52qYRwIfNc
jx7YUgBfMK1OOrdNg17V/11HfCUc095itYefmAw4vSwf3YKCX87AKceMZJK4
a2ci0chtSWeYKw+gf3lp4VzcseN3Xp1raHMPDkS4A7yP7yRMF7Sq1/lha8I0
YsniAMiZp9gLW/pr2CoIzZmD2tRry2bcXhUyXUT/CEhNftmNV/1U4bTQ2tL0
TWqbArCN8Zscm2YfcjaipdEw4r+25NkLXvyZOczYvOzX6/QUilqg5rtAItjv
4+zaTL3PtqX0mO4cYtZ1Z2FdmABkdaTtLyFekqzAidQ8BqMDX1+yiIjVXIK5
5F0nTHQoNQMW2wdEgGpObQYm0Fgs1QzhqdIAfjHSdaaF6kgC4dBFG/b8DlKD
JaD1rFbraxzFZl3MGQ4pa6oZZ3Kq+qJ+NM1XTTFm1oOesC6SdABX6mV1qiwr
ntTFjcGKbrNdJyxUcBIDb3TwQnhUXGRTrDKYo1uElPJEz84MTUYQs3zjPkvZ
k01LMDEwfeGGTy1HdTD6BnJM+Q+P4wSLAoZfJ87MvZlIXjx2v8SkBk1re4mM
M6/wgPeGDtRzRKBZtwL1sC9aUW4gWDqDg3SuW4IcsT4nyBbvNrkAZoqyneO5
wZ9mdyZktV+Epd2fvoSb+UqwkwYQYeJnVo4gjTaEI15Wxww66jIxCdA/SDid
SoxZWwwagkS1dj+S7gefMqieCicTsQIhR4SHBza4UBhfFTHUbb8v2xDgU5oT
i0myqFAisa5xpmf21iV5Q3Cn3Xff9vkrp5l1GATnBeHKp9MfX4S3V6MwNwou
LNu30Zt6SdxdayFjA0zHToIv9qcu4oUTCStCNKYVNG8aqrxv1TPvtnZHyhB9
kbL+BhqMPFmikfmYCG4JD1v2WPS42qNnpmif4SHfVvmAbgvqq19m4Gcu1xuE
Yg4yURdUSUnLyB5SS3iQwVdVckTl5Z6Ng0H3PxnefQx+qRRRwrMHBZpEH0Li
3bT4CMbo8kjJuXsAAY49vDCCEA6zo/zBPg5scUVb7zzfGA0BlUk0WD1VvxPz
3hxlup0FJJnyeIAIdvJFXYLjaT/8hBFJ20mik9Re2q/FVpRF/3n1Z7GKVWLk
lIWVLJ7vA+OlLrh21LjR6KqOoajKOaB5qoRzN0IWv8NngrJlD8L6zCNS2tyo
MR/ifRDrhGknL+5iStOmGSo0H0cMwuiPHUgmlWwZvWWiFpx/0PhdOlUAOa6c
NuPcSPN/jwzgoqlgqNs6ZrXxuvDfP1NV8Js57P1Hj7CsehMhOHU3hMWfi7Wj
uw1UTTdlkiM1jTdSALATnW2qY8JIwGeJ5JSksxm0OHcDJDaoW7tSgfyxUpj2
6sEXyE+HaLqpZSTshkrbHK6mVaYbjWD5m5/IHUvf6bElVBARD0s0CfTSK5xU
Eg1spTJ4n7Isqna1juv0MOpIuYSqxYos4w/RUYtIUINYxs1bI5aVcTu2Tvpv
HxwAiWF+mRqTcbH46e/k35OOM9/PHbcM4xov7EIFEETOCtTVQL+vPZJie55Y
J7oRSZS/mn44fOpjgva/OnVF2bIhtge9PraXyQ5STGCFsGZrGnsJ+9kWMOok
VapLVLeeRcxqd0MO7L6WSXtWKYP4esl5jaekR3nzfR+XE3JWuCr02LthpNMt
vfy8JkIa6//IjFhHgE8Wc8CYv2wXDeNT0fUmMzzq3CebVn7AJf6p+LVoaABn
RiS7a6D8VLgtwlsk8wi41MVH3HGtGXP6rAI+HCqit3m69+ynsRW1LJyF+NpW
LEVL1JNz8N71yw9dEsgYM7yADyLGL1W+ZsX4MJTxGML0cEVTXqCICERbkoyU
DvYPq2xVkAoS/H5/sCUGffh+iKwIkT708QGyiGLv+wfgnKPANKT8AyAvOlCz
FTzvGlwp2ysHz5Ab12srBDX4VXw6Gl6P5rHhbgK5eqM1C0kN9QLb05ZKjdDb
UHCQSFPrWRIButW6B3m6Fb4RD/szXvgShZ39A67GYfoRvjedGia/4sbVwSk+
oXb+qpWrneaON/92w6ElW/ORDHSlKPxG1rdgSbmTTzl2Vc7UQKgu987PCylq
MQxNRXmksqGhx2Dmqdk43XXvWJpRb9syHtHPd7bACsOJ5RBUucSe/IzS2y7N
apM0oXVF3KDUGL3lw7xUJc3QM60tMnDcz5LSc1M7/kKZnhxCCp8oR0AaeCMq
nb7bg4Z0GDFaK8BmC9ttH3gXUUUWLvBUOLYjTQHs8NoX7dQEIQF96d/+exeK
8wnHnWFN8H8DsykzLfCgGcq0qT8CjvpZOOGnXrotox9yKMPZjZelzn9HUf7Y
IgB/dEltVq2aNP7pk/45eXSuFkotFuGzSHARYslVaXXMJYj6bCreW6hbIOlg
kGN8/5hlNnIK8WfLlk4+uRgCKPE5GLuyLPW2D3zn0E9bxVIXy1I7Nq0F8ndO
mzQ2uk7Ys2SuAgB5KTGNCN8x/7SAMvvmdyJsTF8mScqS7hAFrs/13YIFaepJ
RiX4Esn5fInfuXc5RMhuiOEm4IuBiM4TPSMj5eEjVyQEbDd6SFjTaeXadcGs
IpjcwlBmzOEaHkummvlXZv22/Ypw+a1C8Bh1Vy6QZvmVoGazuKDAi6UUGJu+
fbXM7AbI6Abad7EhI+GmKz3KmUzvyT5YVRBHamzB1039JHFpG/XVUWtJKpc5
KdwZB2Em8c29Ew8JO6SCYAOE/f538OpTjkqPCr6sjdtqno//4JJNi8W0jgqf
eBK1nkRIsz/cQhGS05H2O0B4iZAiyzTOe6nh8gZ2Stw50kGGNM00Q0QZSKiS
+7lnecqMwkioROIYwG5lK0RZSYJ0DH/MbIzI0nvz5dXM5aF0ULXFl7xShhiy
XbmnHLSMoiln1AxR5jtLjGXs1tVw7T3VOucN0xsKdX7NNzYq+gQy6mab6gI6
dchFCRI18UT+G6l5EKWmUL6sg10JriRnze22Nb96rXZm4U4nuvKJC9mdqopG
LrrWsylDCWHWQMIKXR4XCsFvGh7AgAzuIa00xb+UmQrnGRCneS7TdzS3fCNx
cFPeA/wAlwWHnr7surkjZISrbwHeikeERKDVvgfIF6sO+eFuvWwE74+w6Aml
Yvv5AvV1QmXJn5P3EtE8lcekMo3FxBo0uHnVqcz/trWjFH2za2y21Auu8FKT
vFxe2xDq0mWh2dY5bCEO6+mW3V87dkOTjR1PZoFiec7IM59xn9TCifU9BSKT
yOgosbHIQeYasCpHjvjjBZ6On7NZJC0ja5kCoegltrP9h54/s59QvUv5WFn7
BgyuNdULZ75kQGNkQUOF43nkbW836kSv0VvoQ1Od39Cs446hNPC87pL06sWh
2gLkBVCWGvdJHcllidy3rP+HqjuHf5YOvT60vkH1p2cJECVi+yaRG6s5ER59
CXzS3vzmoxic2tjsyDxej58si5YSPY9N2znbEpYX++B1363kVdG+wp9eE7Qd
jouuzF1eft16m6xUNK4C3P3Oo5AJ7ulAyEeQIueri6zNzb3zHVZ43CzogA6k
E1oMOxPLehtO8mTzIf2bqV6dmETAZGnd2Vba/1I8gzHjdXy7e+qI4RJVbgZg
5Tp09KTNWMVKdttNBd+jLHV1pJVLkjw2wy6fcsvmqeXEF/NPBU0SAbGJtfqs
kda8k/jPl3U9faUAnaCdXlmoEojAcLGbs3VUo3kBFMS9olL/aOmGipqtdA0t
2O/F42TNuDcdTWvJkFBbE2OjreBmhZopmMkGTiWwDVoy+WScHBFDB0Y4FrRm
nGpiSwg4lZbgxT7JPMoKxoBOncs5sLKDcyCzxAs6LiDUXi5qBL41om2cX0Id
km22G/Qde9XaT3VoBKzkNa6p59Q4D7P4/sbo/yRPd+ET1kjCZJEJqUq16Q8t
2PESTenlPR10bW7pD3dfQQTrvIqSrFSeees45ifGz9f4hKiG52t4fWZpoTbp
gySZfwiQfXk+rbmteTlOxcOBemNtgWWEElM4u5lAar+a9WdW3XVnvrq0fBoD
RPeNch7ErlIURG3jr3vuU2duG0W9a8YdGWy2Dyrxal+4qGLERoxF8OREcMr+
9dLeEUL7x1VY2M2anfohAvADMBUDLmzniKiKeuCHKUOxJDUz49jmDwAKzrVW
mMml6O/q5kJEk/hqx/dCrcVTT3DDFXEaLWgICTUaAA+Rj9/xc5pnlkPB8bYO
YXyQpE6eHpebiiuMT4LXnaZK5wnWA47AFqQz4e8or8mVGOzw2J2lWE/pl9xO
msTy6I5CBnVONcQ7I5YKOjeE7k8tlZs1tYWAR32/R8hVdS9lnxQVkz+qWkuk
M0K3KfVaG0h40bLTRQPdNK6HMeYS2f3j2ONYsgDIeYR/QxiNEUnJjsWrCrI5
wX2rwB8LjbkU0mm1a6TFBx3oHjSujfKUghbrtHckvrwk+kOZ7JCsIi55SxGo
Yvd6laYwwpGM7HDS8OJcnqynt2h0cbi+dgHntf1MpDxFWOH595rhWW+NQWgs
W1mn5Fa6Q/wXCf1mHjxk8m3N5WcvTKEII6C2IEymaXmQDzmi0GHX7+gbLrF8
oawC/YpiP1gO5n5lkcGQaWawtnmCEVpasFIDkpUCf1ttz0K2Qi/M1dVnXttA
Nadc+p+Kqb+/UytR9oQUjhLhS6aWqM3bhEem4r4eeXv4LQ+qgg0A92++k2NM
IV5W3z6O8/PFZ/WhsEc9OtajFdRdBqZJDhrK2Am45HzqxJU9GcgVKnXvXqcJ
ithhakQno4J1flJK78U3nRUojcqOykCwnvefQpFIGHIKusJf3FIGnNOc1k+W
I52IvRcJNS9Uf33Xk27VlLacgRdNj3ABTLfQlvL7rEo1PHylPtj9SEPNx4vP
6ldIlJkH9qwCaC2KBWhqwlm9ncRqz2vepVJBXspGc7vG7qm1n25d0NKWaVmz
DLlaFUMwrIVD53sCgxwBwgspUfNL/DTn+enm4z9ZaDqViKzHwD25PElfHRau
TId5kjrJ2QRM98tYR0gQdpmnHIssEctdoxX+zrrrNQw0vdChnDBsREMi9PO1
Blj4fAGahkFwrcN6+paxEOG1QbFfEEk09EshPp2a+rMW/LHqYnRQxDYIoAfv
CKnulLbctEk1Z/jcoWm/sWgmR2u0natZ5lV+CPpBXoNPoztFFYFsfhQuwR7r
d6xFdXdkD7FXEidojs8QJBIRxLRWezrAZETJOs6cmW0joza3Hr4nx/QkaALo
R27xp61sGtO9HFidAZJnIsAkinbxzvLFzJG+k3qb3MeG5Gr1/apGrL48aBYf
6Uo1rhVsp8jmN6juq4kFfmCSbZ2K9efgNoZHUkTqABL+BBHZRENHo5HacNke
k29fS49x4KAhBJJnMuIuvBC+2iIyz4ziWsjKM7jp4GeZS6IJToXWSgTOBz1K
yum4LC6dBtVVEnxpJy+84EFyQrwNhe0ADMcNGyXKXuzXVn6EdlO/1cu2tZ68
VK6cUhkVarNvoWtLnOPkCB+sjd9+vvl8WJPfL2RPzv4AsiBqWNZIc0AssDET
8Cqr4C89g4a8UtgTVp/65oWqmzAX5VBFbNSxUo3CklK52EB1JKJ5zfHRhnFJ
3+5zOzhrgTtqjgX1kdYsD4TXU9iXop0bgJMgqKs3uUX+NoOdDkp5ry44/zJ9
4MMwRNK1Lu7phztUX/cEhp2boAyw6bHluABpwbSJxvSxIpENNUdJ0HEvnRIw
By20JEnFRq5+u0g1xehpsKp7eRj1LQOmyfPGzm82pfVGI83Z02v0Bxfp2ZkV
2xY5uLIfBgkXOAxUkmsv62MD7k+jK7268ECH3cJ4X7S8IKeodUfI/Z4quzV2
E/NwT2bEjX7gZdhIp2Ky2zwAUB/H8TsdLOAQczXoVh0UeJO1BhIRWd08gS93
lfBm+MZsxj6kx2WlGbWFg3vNwPVvVE5Pa2Au7j/sozkWnVLMgY5LFn8FtP69
eBUgqC+HJXJ1iMKKKeDD7q7P+9Mnb4FtM6LXtm0X5ZarOV5Luqjs9COEm0Vo
F1ijPASbzx5IR6x5rNI76UzQH2fYR5/EKEPu2swTNSTY16N5B++G1+DdYT7a
VTgbHLO8ozkuGtpuKDw9JscMkUGHrTkf/+Om+cTBVVTl1w9bt+/hAofQx1v3
EMEgkbs18Ai482tNHu7CnI5V5ilwXaU8BuMlg4rE+8pHQbV70b5Kjc9ET+gG
lz4jCJLcbZgnIL7aEbbvStC5APcorMfgrZLxRi8Q4VpLfPg1HsXUvYbbs9yb
Kgx0LxfBQgj81RR0CH9bj0sdV9XVwYSTviykQiBNAWma4pAdxFZK4uiPADvF
QDRFPyfAIv7lgCU2yFafG/eVsv8EJfORe5YgnGH0w/xznBaEH2WW/df9Xb5t
HErVpbFdLwXin9OUpSJHz1qTIHr6y15cG9CKm2LvC78afxPAa1hG3jTiZF4J
1y5xWquaoNa8uxD4pmnQZsr4lCzfWqGCwcRCyhCvv0clxQwMzHppRNA+K2Q+
H3eCEIHcIGe2Pg89W7Co8jS9GUsK0sKonMfrqgulHaLjEoU4Gl8qoRzjetTZ
5ugN0kEfmyIruHVdX06NiOhaf0wKzWEBUQXuHDV/lMGPNw6Fu+4l5TIGqEbW
a2tQwEVh0+pln/zBRbhVgLmw8Ux39mK5VNQBGI3kyxgm6/hHRSKG/PEcxmde
o+JfWVcZVGm0IysXtC7ZLn0zrlgOG42X2p6eHa9uyMGKEYqfful34eYfwH3t
k0Ha9GR5Et56AJpB7yQMfa+Qy8lh44vHsWKaWxxl6OfVffF38LiLRG9tNZBh
0owjxZ5eKoIcBK4Uy/7LSHej+AHdi51jqIQi7y6x0jYdNYyrUiSxJjyHKu7s
BW7vuq/f5ni2c5g0pAaY70l/YCfqJ65TqaA/kEKfYzNwO1wOP0NLPn1QvcpB
pg/Kb0muewTjrdPKei2tF3WFJWRm8vO8bgGDZH15pt7iPE0HhW15YLUZhwr5
jJdffZu0rUp3/0/gkHZGxTUdioQe3n+I5Hfvdt0S/eKPHZQmsxCisUmVNe4i
dDxW8Z1zTVYwW1s9TqPaH3K3ZCaKAF3z+EvtCszwkJwXh/uadf1NxkUPQBDA
cyGh+dh760V7ZjyUQh840lneCrw21iBsFEWdIbPPrjngq16IiDdIe4SNRPKO
k+smELgelx3Wm/NItd/P2/xSeQ+TBB8L006Nsql843DCEUi79W7b1TeqVJis
aWDYrPmwF6kdzD+CAyycAdd8kwI2lM3i9Bui3iDhT5hgbl+Ed120KHVBUpuf
O2FNQUOG8rNZZe2xuze3XUepMKv4Mfylc4PB1+3TDMEdRZ09O0pGuXKqjCcM
NjwNmZkm7A659f+WHq9VJW75r5pApeWrvZLARmDKnDbfh/1rFf7mDhF+1ZVs
yqU5//ln3UF/33hUs5bLN9O6mtW9u9E5U71dE/7xUftVZm6PZBbX5NkaSCys
ZX5IDqxoOaq+soBZufHVetI/3pBLmoZ9GO86cW6qF7/YBCE5OI5NQc2ha7j0
v41DvVOBxQXlQ9mMYBS47vOiEekd0VWSlQByPBb2YG/QMu7UE3CGwOly4F1l
iC7JNz7y6WFr3OqFFUqxZa9eYRjpUcp9TNIZoXFzcbT1agNC3eh/ujBfOwQc
KfAgxpVFVXm+vz7uMnzzrrW6nuRZ9EibQxCmRBo6oFhMZGVjSLuFi22UF5Om
e52lsXQq45qjCn7cq2HRupQPC6/OFXzQGjkeh4hFG+HlbG8fB1R3s6/+61/z
oWUByqSe2LTY3bCzW7CmNMg7DExhx+4mqLZ0viTe9xwVckGqzVQ9XZkPcAd4
hsbb7y2zTqAfg8Zs5NbA0O/rO9YBSgvkxwhBvlLIEICUi13X838zIIbCx3Hs
FCq3Z1tA924TUrN1DDJ0mFxeTD1OIICL4Hzj7vCyly85zzOgafb/9uURLYxt
U/BlX6s1KQr0CW8i/mgpqNhc1G3g4JlVc+STtVD+OAQgM5JcqcPw15y2a3Fn
NhGIGmk8HGgN5LSfUB6jDdzeLRPpAs7L9Da0b5xyEubm714c7zk8JTlHYMHS
WcgjmpWS6QNl4XZSUXQ69cpYp/K9raqTVIppcbRGml2jsTVixz2YjUcOTU8H
aRrWCpmwABvJGmfqpjQmkjqIG58V1oMuSCMOyDOgs9x3bo7AIe4rv4EqmXD8
6ZVckMqOixRAqQCrl0pq8br6q89sO1aeHvrbIvNzFgEa2e8JK2LG06J/Pv/u
A0QBDlMqlnpDqjior3ka6s1uwJllNqxZl8r7LJXLd5rxAdDoB3L+hqmTWAdK
/+Gb7c+Xyq58R2JUQdEVsrEIEqaF7OQ/bD0yEoA4rAqwR6EtFV/q867DWCDJ
0g0BZhEMhkrXSVewFIO1kTmF5AvbcfqlCtITV4WH8k9U7Eh7Dzg1UtTVQSs1
G/A+Vs5QpCc4nsz2hEyCfeE1gHUATbE9BNAP6amXSDUyPGpMsL2DX6Z9EK2j
sFSIBsn3aY3KTltmAcQ8pyK9zXX2Z1t3Kg6iOV78frhn65CX0TDeHP+UrkAc
z15j9wJh6lohkuSBQE8B9DHwg14Mth5XAq7AHt7QLTXwbR+nTBznN8mvRh1H
Ym6izzwFrJim2EFsaJSqiOlQeQHJjgaaTPY7Ro7f2/5wfhCrmi2ZwYQ1o4KF
cz2s+pfU8AV4CwFa25kEJVnKN2Z94K4knA/+zua6NTtjdJllJKq1HG8ShoMz
PV/UGq2tTGHIdlzWL92/PhLd31japlZefh1vtuyWYgI2E46QSUrGF1qtT+5n
qVAuzvbrl2obZgzcWkWNzfnxBvUCFSxiGw1JzCFmb9j/RTFlRgn48nA2HAvB
SLzVmZiyFTwUCN/Ji1HZPbwi9849rV7XO2FXemqjm8w0lNzBZB9EBw7/z9yM
vvjbD0SDQgKMLHrLpcQ5iMyaRnXz96bunecui3ETAlYXWeEOz/3VmqUFqW6z
kfBEaNzrkwk1SHbAf0NsU8aGG7lcq3SDmPp+kHiLIpWQpY8/kckWPd7P8isF
cEQeuGH1uNkboEq1EaZch6IdHvBQHO7yaltXkWGzuErhLIDaEK74NBFZZ8l9
xcc9PdOYPAZUyKwdcj/7OGJQNdF/5HSmGLradZoumob5sSEplUlH3sKn7yXD
itdcaRdePt64E6Zz7cJJncxegnIV0I+Ihr+LgBrR1aWpFXv1DcV1pII6JhKP
HD+bbLXaVuMvoukeF4CjbzYt2Njp8QZ+LxzFN7qmGm36Ojsb0I7S5IKIuXJA
PbgZmTZEm37V5i58nOqB6gXY0kEqHRXLmcfjycVObuCUnLid5aRZrwKhLERn
rf4QtlPb9uVFXYd3v4QZAVvzGQ1fciMUCyLIpErs1aazOK9Isg4S0AcmHZQs
VZqKnm1A3KDayf9XM4PdBIHCuCLdXG+tGEM1kkieeMiOwsLhPeKdrPJqTRtU
ZH14EuXQEbvjQUcx6XkFn5T23Kw1yeIEodZ4y/fi6OmlUJA2Re4G0pyVcMGL
ExxfcTzcKFMKW/gZrQem/PxVmTAQRPAnnMUj2sQCSJIzod/lOioJU7tZeLIq
AjFgipOttsTil1ZuMrFtR45WsHEKpN66tGtoY9ssc5NvyVKIgmki/hiIme7M
LVdOgMBDoRAbCz9qWyuDotUx30WuCWPJfhQcquUDUDbwCup89VDcbWrG4sJn
QNGlgQ9cFXAH8YCdLGFYghjVq4I2YEoZxxtfNd0l2AgRmkKbo1qqd04gAkDH
zh0ReBxxKDnD2t1mNWNl7I30+I/Z7wZIVrt78dIebTl/IXNcGr3e8qdhus9U
pHcxEwLcT2uW4AwV7m/zq9iKaIGbnaYxIpNzY5yx/jUgGUpmmVpsBj3EaVoA
qP5Rk21GMCqR51URWV1yZbGOv80O9MKpxo5d7RKYgGzDGyWDlN9GhG3RSt4M
+/kuoQSd2V3d3nUgeVlNBPUPIvnYUvnlB9PKXJQ8/WqHp/lH/6Go+eLqQpfI
WUnDwIPb8m9oJkcvZ6jTNO5SMsoCaTLEcOMU4hra75kehYW3hqGwBpVx7XQ9
Mc9PNYmlA0j4edtn3yzvt8SJqDHcrDD86HFxBAsKlpX2ZtNx83kL36zaCJTx
tMo+P/OLAIvFKSEMMexyDPYlE4O+gYRgCjhMP5REuN+LVQN15nXDcnir3JB2
uzcb4WNyS2QqGA8NsQ/F3WaMbM68BGg5j2EM4fC4Nzh6kOiU/uEx3UdNMapc
avZLrBRuAHQ2sWEGZ+yeyVZevIW8MkLDw+92u0mHlz3hn6khZ5oc9FZomwrJ
JI9R0JA4XsP5pVQ/7oZBKlPzBrvYPZXHcSk99260lGCADN+ecpQjF99/0aHl
JogEPpFG+dU17taW0p2YhDFN5GEb0BcROjlqF0WvDBpM/kXRwAVMfm2IZSPf
SXhx1oVlii7eIVJER41dOumwuQY4frUaUzTMswr6TpfLbmhBRA1W6tqMw417
2TfrEre7pl2wCTuQJKUk2v0mOlcZevdQIk+Eob6maOXW5umcW+acb2fOKY0J
Lh/Q7MZILZ/5OXS/Al/tjJjR9gzXf0B8zEbRSZbY59FFIu5i2PZpKH9rKqry
9Xg/lqX43J77wqSUhO1nyb4RYJZFQ3DWTeh6z2j3CWw7hnlzJv3AELSWxiSm
BYb1FZHO2Ok41pq5A8xkTkdait3kFEDu4xP57qObn51d+a81E42rzUJNuN9Q
KLWsJoQ5r4mwuICIOtA3DLqD+c7O3qXnvrOVXDEDst7lP17dhn4Fi9yS5KMX
jdm0Bzj1M9U9SHelOQTj/+fpiPKEVCQJidu5jLHqweEfWiD3ExsASQSxyOt5
hwU7Z9CNnsxqsMKPS68ukFjN9A9CEbFFQBbdjtgpD3awWCt14octN98YgLCs
0ETWMBQdDZ/9Km1iF2IAO8zyY42e8nFcGT/I/q+5VDqSs9mVHKb3AGFJ+j94
d0SuZfOgWVnIdLQNWQ9p7ajq/s8jzlgIrnvVETyFFIQCaFgpn4qqaMRZjwqW
OesDDWRDhsRcBY57CKkGemC1YVzNKk7kG8gy2LpCk8QpMSu8QpDVb3J+ff3k
LR4pmHdPYdzVcfJ+xcn5MbnhTlCMljL31KxectDWbOBWQRcZJ/zMASu262KE
wrmZaS+q9fEuXTgrwUAXxnyoFK1uUkh/Hav9zel6Hyuht4N6KInkrFN4RP+Z
BnjtuxSarnutxpqn1Nabwsm92VAWSETXdk2G8HyvpXA/be4a2ucwDEZCy5As
rVbuwFAfOYF9OI9l/uFflhR5d+4YSIzEpNYjWiQ50PKg4K9linEqVFm1phVQ
m1v6+6hoQiEWBk69b87V6JsAsTHFmsG3vVvAk1OvVYYoP/CnVQqfXqp2MwM5
VwKpoaFvGGL/dn4x7yEPi6AReiRGA1bLE6nyq6/jt/6PsQyd/m22x7i8YL/M
LjPqy6LWVr2t4E3QUt041fxyJV2kS68eWJxPUMpuhZD3crWi7my01t+zFXsK
DoFYDSrAq8VcvJEJYBY+camCBK4O+6ogxQJ3brWb01D1I3gAKMD63EgMLlAL
vWSeoEmNrsM53tBuHT81KwCSfaYg19sdJ2rtUgacgKTgMGVeL0iFc6i6xHzf
Sq3QP2lEqX3uygFzdvIt+q6EI/BUNB7PBe4p94TjXAkxRq5e3JH0vPCbya8L
74ecayyeZeeHhkgO/pAwgiX0USxxXdSpBqejR2nwc9ViMmpwwOvMKahZIO4l
FlFZrUNRQWBDgIiBh38jC5IFvdBurtjHGIAGHfN2ckSeB1qz9vyxcdaTxvTJ
Z0qFHvVp40iyi48zU5U3nt+lZ15ZiX6AF4yWY18ITqONd5Ym09JNCvYyK0OX
X22yet13dzkFfaGgSc3OUky5juS1ErOkhfkg4qQnLynrYkZTWM3U6wNOmCye
E0jefvDT3tLm2qGv7UP6t5aKawzIlXi5rqs0tKXnWJzu01Jdg6F+UZY1y59L
qOmpOhtRluIzRkrN0SHNF5h/afbx8Hu/KUsMk80StY70YUuOiNxSwnpUx0Hw
k2UBPHVNxtG+6CIP0wiY4XTksK6iyhM9GPhFMx8MU9JzMIqRyJ8tTnrkSk8z
Ygt6b3C/F5mJnv2XaG7WGUNOq7YK5Ad+CFV+rkBdo/xQiJHSDLQuzzu27/OQ
L2Bx7YcBf7jt/tZRPo+NpIt1GQlI0/BwICK1Axs9dKvMw0K4YsVuKsdt7DYL
0qaDJ9GcpXBjpnPmSAu2WTMKWl8rbXNY5JBigGayfULULoVm9xEk0wxVY4VV
tmcVv74HkaK3EWdRjrNtIKNzBwZS328Aa2yq7u4kfxgWJYpTLHwl/nCnJli7
kLUJO+02HYR9RP9yKJPv+5CS/AkUw0iJpB3okRVXlEfZD+/7de4awriefOAQ
r3VV3MDIEAvuigM5iHe+e9vpw0e7baFJOarnAVatHefi7WvNqpQYtwkeIsCc
z4NQ15zH4+MmrRHGTJbe4MbYG7+R6TJ0AnqiIBsWu2izb10WB+SleKOE3CCF
MjEhWuS/VAIhIuCz3ZGnXZs6O2eSsMEqO0vGVnSZCVaYhj1p7PyBvCACXyLQ
t4iEoWChMhiyf3+Rj6/OWLskCrOmKkrwx2PzU2OGIL7bDMXY7D57EkTQNsAg
/JSVHsj6tc6EQHuUFw3ojyYS4o6GABkdY1rCuT9Ag3qoeRLAh7lgtHuzsmQA
XCe1JpdUuzLO29HY7WC9Ox5TqXknnt5eayHSWXc9Rf6sI3m58bAVKLZguWAX
noY+6M9K5D+2UWQGqaGRKnicLYMIqytSlLSIXK75IZjpED8B9xc+SwyQdWzh
Zl+SvOXyUhoxE447zUWZCD7b5Z8CJP8ZHDgLQbfmjT3GdICTu9cftAJWNIG6
Vu8LiM5hEj1XgoCqqOr8HOuB5Cy1kGq1552P0M3ymfqcpX5FyjwqVloqE5B8
vZEPEGMe8L5zZQO38Gy+Dto1RU+XkqzZV1Q+YEEvutEhchyD3GtSeLsCwTPY
FbYSpBumBsZCEV/O7dVwBxdr8H75xY32V9TK6vr+pmBHqG/+rpymmIWMW5SJ
0/pb1OdHEHb/F0F/V++k0gqvFkhyZzvoh/VyZOW77zXQWdRYgs/rLIv8tX3N
3KQH6Yq9Sw78freyNFR1fxq5e/11G9S9QncjLsiiLFIUxiIyIaDmUZjPwBlw
tIh4pIwHA235nvFlI5/0hi4QpZGBwBgEjaDT7Pc62Ctqoqd1Svk42nszic+I
VE5bdZ4DQ0F1UlJ7JZEkq9SkzyqdM4AeOXdXNBY9Tq96Qpw9QiFpVOrmUsPP
RIV8yisXlmu17xOPq2sYvR2AcNy25kf+UEGJHgbgyJVc6jgx14w0xJcY+KOr
i58ukMeZUG3lgEw7mZJyUFHe6mpymOgIzu51J/Ryh65UxEsIC4v5bAq1Gx++
Oi24l4FutnBX1jPuy/T7/ojOtt8unSabciLM7dgBcChSvO46R+Fvl/VbCg/t
vw4bW06y5RzWDPMN9gcXMieiUp9/q3u6m3LDJ2cudEa9VH+GePThqEsHBl3S
Ze032hoMRnpIVQlmAM0zXCh+r3+KmWCliH35K+nsm5Id7EizjQYsiFxBTTEn
FkgJ0QRTn6Cd1OUFT1iYkqteDCppVanN0yYxR5QXuAu972d+yURu8ftksun7
FhwBpOo/t6LU4p5RqRddbVzSb81Bwwd0oYjMgwCqCi+DQvFt9fL4EHUp9IVk
29yTLLmeL/V1z0xvepK0gqhuirH6f1VZVCAidb8ioZRfELyazd5ploZwMxEZ
Jn33R/BipgzD2bI59ukG4gGUvnYhT1ISXzwBq/RGz48GIjyYAH/nwzQ82PT0
K87AJz/8V3zYAH3bNd3wET0M5PhI/69HH1yY5BbvndquKIr/Yg+r0VW4ECoc
Vl1qcyeDwgakgz5EoTKyWqHgBwUaXtemQCns5x+aEvJf9q/08imKPrzXfqJK
nm1Jv3sGoetIN2KYZ4ljMDtXnFqQoonV+XNK1D5pJxH5Wv2rwnzAyw21Xrnu
WmEXQXSElu46Ku1kzMHVS3QUJQWkhQlQcYLu6ByMzGBwZN90I2nFME9Al4e9
0Q5SAsMsri/rgyg8FrkX0QD1bww9GLyqyBhSlEcD01kPxAw7k6yVYr02IqX/
WFXzhEXxB+CAdnV/tPDeSzxpflWGQRlAvteCJEtUNaYld7cT8h3RwnD6aerI
tClMcIreXBZ7YjmSLno5Ua6MqAnMtUOGGB0fujCdM96pGcSimKTeELVUnokX
/kSvxSzUj6yycaq3nNIn/VCvDfwDKVyVp4R1P3Ve/IHHEFME1zkA+3ytTRl4
GAGCj2crCZXc7X0qDTYFQp5FviBDlFg7RLv+YxdeZoZRCDmMzqIJkVH7cfn/
MGBpsU282UWs2+p8wWk/pn8/4kBlxT/fw6vpkw5cqLghC0oOe/HXLN64nQyh
NxYdXO4Q3h7on0SKIU2b++sJWcnxluXNciIPmdvmx5hCDINRv2hFzS2UxFTh
IVA3J+BY006i56G0BWVSq6GEWCa6+xgXtil+d02VBM1PVeTtIUKkuU1IRL7V
prxhJ5Z/QQ4EKNoBchMLViDWo5kUkdZFNa7KstA6BAVf+7vG1SC/yAE5unCl
ZTnowvEqFuJaWaXfWhe+xp8QvSoPTp1YIq0+ifuKsoQrsw37QgGdVer+uWTc
y3vxM+jzerTD27/BQ01kEHBIcAhM/Yz85NQDfnnjAbVk/RkOrvUP61MBLqox
0piPI1h82OhnWmxjhEQcwyULeH3p58Jq9X/UsZNw8vdsrCuvTp8sr/dVGeCR
D1A4c63lalxqNVxAykSBMs7ImyvHV9QmwartUcmsgSmN5XrnarH/Q34OKAKp
ZI00klyColMrxdc5GOCPzITlanyeROiLhSxKX+UHJ9yuIRigW/c6FllfsIcB
npwu89saC3YuDSmSD69rHYSvNWlbUZLO9NADVWn/ReFBWHgVHlhLH6cbaWTy
xf2LanBCKWWeM1dfwpVHLcPVNMR4XYG9jfgdxE59wHQzdIAotyHfyXMI94u8
ZbSZJtZxNdizEKS3LGrLaAyjpFBW4nh6kuyr4Vry/zI1t41bun5m1ydCOUuM
mbWpiQPM4DpndOfauKI4wptspQHU2lR8zhkZxQvUbQqYUIn+ddicBVp7juuF
a40SqhTDdYkE31cLj3ZfA0HxDJmRnrsOZFS84rHaX+Ylp6pZ51ltcycvgAPP
eIdjJABxlO6zDmXWoohvVzBHYNaoujadqNKVmy5uoD4xyHvYqRSHSNaQa6Bs
rGsP06elDMZLBJKlgszYkxnkDnVszWmcFOBRn/GbKKurefDmE6jniXC9TwZE
RTBdt0O70okc4CDBrOEM0ltgxI8NqSOycfBl4MvOVHbv4I/6w5CEKFn7djoa
di7VGuHl9jRGXZa/zxneFF8yBfzuZ2WyJpOffNUKZBFIJ564OIKyQSx5iKSU
Lx2MRpQo6W3QJMaDOoWvvjqOWqvlZWC4WvJVccwdHij4myVqR6yLeDrjz2CV
LflXswAeOKVrPx+WBEdd2sP6bBILcScqZ4Ax5ylAg3O/CvudEiloCVyqIdRK
fVuGcXYbq8BRjb5eDUIVfJAPPuJyLH7asRuEE/d8HxnhsA8f2lFQHo7Tsyzq
o/TIZhxxvHpYBnqS7pe0Y2rkXUSRVuYEBZNxJb11BP6hDLqw9GHVxCTCJh0A
CsA5XuiemKuUeWygsgngE/Qc7EeG27Ns4PjPhfoks8sZxymp8IJx3QQFhNxt
m2P6DcGJy3N58m268Blome80Xzu9YHHktNlMUU1o7jwxTcscA3Joa4Oqrbwr
WcXkLpKvZMbURziMmrqgdVGoejQdOhi5iHDssBKnDuxWN6WCAbW///z18g0p
SllXULZ6Cg9FhvvDe1bgSxmNx4qjUJKjIwr/F8ysvarIMxKrkg/Rgt6F7eXj
Ny6NSLTJXR3r8NnGhGVBWAzCq7cLrfDQwCVHWQ/bXP9eRGFIZY0zPhKanjM9
r6xTkqDtZ9DEKBx7C3VMbJ1TBnL7HBMAQQyy1+J+TOA1xva8p8h8fgqMTRHQ
WHj+czrS2vQ067PFvDRcV8tCzh0WJRXHzv58kSsDxeeqN95J4CCfcphv3TQi
zqFo3XIYdFQYlsUwYr8jjccwQzqopHir0VgLMT9F+/W1xnCfwXnM8ZJnmbMG
M2bg51MhcgBgSerc0nah5CyhAdJZp1AM6UDIg+OohbieZ7ylpaNdb00lFKcW
WEy7LcqjCeVBJXiJT2bTNeh6AevkNcvxt9V+BcV85hN6lcnDIJ4AsrXJO5d2
j/SIIm8XCZGafVOsGV6kLtTUOApuAgJFqv2iHowPNRU5nostCSOC9r5DtpeC
id2mkzWMwAABgd5+Kjg0XN9p7pUFYTeNF541mZja0WLgo8Q4oKBtzDfm4AQv
IOdw0lJ1q7znV+T4RfgfVYOlB5HOtcHg6nXyvh2qfDZVdftoE4Ki1v9IxX2f
AdK/kKZVnuslwUNRV74h+pjoKSD6Hql4ftm27GCmIayaS240o3RSpldIOES/
ypm8bPnw4Ysz9tWCEb9/SXFEJdfb5jBrs3OFvPl0wfBE3PN8ZwrRM3rAE5aH
rPrk/aF8WGAZRyecOGA1GBXwTEW58TZyy9i+nsc5lRnuh05Z0n9925SK38zJ
byqkf8nXdFdWRU1oy90XbfmBa/NAsDyBBaK7X+atxrwSn8HfzYQ6HtncdI6x
umjiSyfXbzTDadbEWvnWo4BxLmz5cwa6l9jv3X3iU2SUgUjXPVG2ald/ZX8f
roxHsG+EZMFVL/4jdq/Bb2PNccQ0RL2P2KtU56Ndv8+JMnCJ92qGN70E+KBw
dno45eo524hHXT95TPSHPtMKZD8YEopvYXUBJQQhkOHgOG5wUvj2RpHuADUx
apMEsclWofQFLRE7nZUyuyoZhLibmzQAXMsg/pCrK4bEa/bJnjdYy4mUFPBE
NofRhEK3lix8vASDJVA+U2/nA9N9F//7LWrjqgFIigD9XT4/BTmAVo1z6M0T
BcIW460QmP8YykxuS9tUHVZJt/plWRSg8ASeXFk9lhQi1i1GJmiTW3z3Sy2u
Ad25UiNml9pr09YLQc16gs0wZsWtASBFJz6usS9SN2fshUKk4ENE42cs9ODO
/qGu5WneFRI+s/vw2lhB27jeZr7AYJb+MZiRNPF7tS664CjPy3vF08qnNff8
hmR+X0gi1moFnVok3rbkBKNV1WdTYFEa/15fvuA4+OFcXMBalHvhLq9PaGgf
qrt+K0chSjGqkHZ4dbSd8rBdF4roRQ9W9yTpnvPN3AK/teWuo3TyFuKpGrum
7CfmRlQHuQ4xa5ocOsFGeH+e6byNJC8NDsfEceswr7VMUdlCwSO5CEUrKKxf
qQcoJ444x7E6AvWIy/UM2/exP57w9oLWj9KVLsV0LD7CyKgNRPFxnDeEwKdh
Goz2KwMJ9OhxOxNhovOGlNYRYz2+OjaISdileofLEBYuUCscebPmjZMMTUXA
dCwUXRAuJ9z8Fidn6ndEvw2YMZdEIe86GR5pWB9zrI9iGQtPCgovVLHcVqy5
R4gbAkrGTT/KzdG9blmB+9P99VcMnX2zKThIw0mGiuNwB83nvpIkOQRM6OEG
VKu57xBYAsINRlzXaROQ3oREPk42DCxC/NTELY69NiNul3flM5N5TstyLyO7
JVcIKH2Oz8BGElOqxTnj9ZrgjDollGtUxnI4bQw1MC6mpz/Es2jFqqo0RAtX
inXMx2c/OAwjedyGL5nCtTN2P76dVCgvd05BHbgDVo2+iY5y9W9bezEG9kDI
vGTAJ0mim/SrswQvT0IduZz+nsdrRN+DPw6+UqrXy1dcotkYVcd0MRA2SinS
deCtmXEKv0BqYxROhh34jDPSRNbbD1KI/MQT5wg4V6rLg80JPUwh/TUO2IPj
/vWsQMzAADlABAPl/wWgM19lNdEVKHLJiyH+bmw88hP5lFtX77Hru4mNyQfx
IbrP4ho8nl6bzTh7Ikcp0iYCwOzCg12AMgfLPrdyIVjCUEDEUWGk5q6F0baB
ge9t900uZZopfR/5b55wt4C4LeJe4dHJPwi20pUtjojFWFoCoWkNZHTWZYTF
sV3sLEx9cV8rUlPGPyPtCBvyPWhGMu52WLmCQr+tRCRyrcCgvyhEoJ/RTzVD
aE2Ljez24tRZeSOBrc+EOZg+nw+O9D2xBTnOgaYV73ItbfPgQ0iJH5vSttWR
mDHpy8yPoCGW7LtcV7elBqQOzConKYn/6puBbTzzclTnv7oDNqURay2wNnfv
nxO7Rtztir78z9JYlHsabUpWcTDegI9DiYjF66jOjbBb59rj/ELqCNx0Vlxn
APtOMOPcDbOioKj4nDLz7JYG0RUVYJM8w1VHrTTqTLKO/uA2EKB/MLPIJRDp
EHt0YOIhonpYy95gfEFgrzeoczZfZKW9qqldlt1R/eUGzvjJ+K69NeMBzoB9
uW0uPTW3SJa/Y3vMBHmKrD7TSvSJwCqdJXCfwzORP127AA3G60OZJkC+c00C
DpEAU3TLC0Orlq/te+m7YcB/7d5iby/H0jpIQBeqSyCPV5uf16CRfVXg7dFt
yTB48WDXagV6Sr7tztY0kBPGE4N0J5wb1HD+OdGMl+ahg/iMUPTaks0ZLP9c
B9TJ6bS790zosaaabASk/Hp3JrfqvKaiZ7+ImoAXei8k7V8/0qyZihwUKXu9
pj5PAqsNtFWueeSBHRX8f+zcw0pW+qMxRfjw0lYN7HCgTB6AnfYItHUkJBX3
HZmiRoLIzIm0YiVjyjIPIF29gbfwXa0LsJX+LwrVt8i7A/s+OQ18/LmJCVb5
LGjLMi1IF5dOnhbmhSOyeE2alAh8l+Vtri/PM/Jie0/gpy1mikpQ7YZdJ5fK
+Jg/uAQ9oWy0sYvmt7BG+2RDCJSrryRFirLTeNVmxtQeJ9O+9yobULhNRtmH
UAt68F+YWmHEt4NEFHS+FtTOdblMM5osSJDXxQZTh3o6vYQUBTTzaauE5QRl
mATpv64O1g8dPpF2TZ/saqJnMLOj2xhrW2wy/byooKUHyGpl1MSNam2oTR0d
DnlTcg4ddeVWQNoJsmvSqYh469bswlfodu8mTm5d6qZIfC/zsVPWEvLo91fq
qCTOW9VMOMGeOVsPluxPg5L7/mu62M7dX/bzJkksL5A0RC2XphFSpvSwxt+E
RN+7/B0ggPhO9qHBsdgiXE/ORztl76YO6F5ueEx+yQJeW0Urvv27/V93x+Gq
fKVCM0/eAO/KJ4FUdKL6s5SmBnmbJ/J8pmUclh0rAToAHFm4pX6rUX0J3xnj
5UGvTU8X7XC8Rv21bvVIgDkAx7C50ZhUWIAZMt7V0ZE6AemhY4SwM8iaqyPb
tXIBYN4fhO+RezlyJLbxrUq14SO3et3Gq5G1ljT0Voj7CHmnJxJSP/huoLNg
LAl1PdFgfM4ONtuIV0L209cc4WiCiygJbbZRdX0yyu42Ff9dXGFLB7yKjljO
fic6os5MNAXLyF7LkYgvlIpS/NbVRdgkPskBwbdDYnX7pXVMKXQ/fz80J7/7
YM95LUAxr0b3ov81WsYcNbDOrUKsIXL3Z/kcOmYVj4Dbl2wK6UMle/5YUDZW
AY5QsWHtyPNX0G6fVBM3kmwddBsg4tkJlTsdGBCoGGALJlT1N8llNUlUVpj/
SmgFtMTu/N2jVcR9hAIRbJhHBDzaq7Pcb6VznF0wtKj35ygL2SfgytKGW6+0
qZpEvsC5P8vfBFmGAX07FPcyv1qFN4y67phZ4velHjlTcMV9ZlBm+UPiF+R0
Wku/kL0aQoNZk+v3FBh96ghrL6Ejb+vWPxIK4HHBqlx+w66i0YD4HtNcHyz1
bdPx6SPEJhsQPOVmhs5HXbXQjS4/n8fMRYLvG0lDBE13DBlAoUdwImxeEo0C
8ohfEFt1Mxx09A3/SQq0Bb5603DCpgV5CqiEmdLgFjH0JmikGKUehH6j/L0K
LpMP/tSvbR6EIEw5gqjYSMbQexTwoENfHhsqxZsuF93yM10HHmX/HLfDmdVm
SWd1gHprPQHaFEcX9TdWbjACg1CFu3hCnXhceGFuskoR2/Q0GcSDX3fUoWhV
gP8iLXdvaZPRmm1aLutCilTCY4ZevHPO5zTXkRrz6ns4sR7GKvIogZCzcqJu
Hzx0wU6SzknM1FZlVo/1GHDaa6ozSA9nvj89URSBuxJ+2orreLPZhFGkHaTb
C+wDnom+jwBc8XziwqMwjRdWcR4kV9uMh4shj9SsiApLB9jab4PGGFU0HKCz
Hpdvjn02ao7AHIx78k3ghK6s+bxkPdjNDO4KdGBqClIICZEbfKyi1imgmSDf
thT7iK/ijZ3QkGE/wjL34GRJqq6rKK9nn14dezsn5AS6BCyYnWdyEz/FFm5+
PyFz5dfB4DOT5Lz0vfbYvDaAsTQAn/YhVeGpoEgiBViq5+e/ikyXxmpz3z6T
aUrp5NGihc87//wzSz8tnp72SArmngBo3J11+/HYvD+vLtT1b7rajMCy+evp
+RM6US23ZHgqdFNzAB9WCGemDQQeVhlgjYCYH8KFFbuGf6AT+m6w7fEdTgKF
GuRHeMjCMydHHD9uHbUL7OrVO8+hamMdr4t23IdeitRN9fvRFIZ3eE48kF5U
da5tqHbx0jwRFmiiXHZ1cIxlCHrJZeMIadpbvttT+sx6HwepKERGM0ZRpy22
JORFpALFtpDjgVXDkcoEKOQnO1bDX57Ch6ICybxl+KtfmPoUGg+3QnLt3d9P
B4EjbHVNUKuOjOcr0W6Cai8u6KGyKDf0enSVBznWCh7zh19QIHcczUmrWRhV
iEuLc8yJ3CsIVil4ALH4t4qLFUmPwmlg+N24L97aBerGx7i+1YIiu4VfBoWI
OKQHHyL0ORWzAcg8E/1J5j2By4UwthHWywMooj/gsIgJZlyS2gC7o14bwIs+
b0cvxqBNOE9ecuPyPoQxhaQ4vFQGfn8+6ReJGtJTbIfm8+sISZG4s/WvSV3z
FVyVD8vwwfi4SUzIrMDZJggd5wcHgLBXWcWur9VmeO9VCflE7w1AJ8yfb9kK
/XaVNc+GrRrVb17/YQpf1WmpQ9p9g3PFEgFlq4kmG3XAzIpEXsm90WKctMw3
2Xq47IMubKxp9zye117rAkPIYiWhyiHooeYLU2Qoz6OJa4dddylJt9xEBjPG
hIv64/tCFTrfT+m77ObAmPgGmj5ftq+EFuNVX/PNpSERGvshgIEWS7ZHtf22
llboXpXzPaQKD2KTCg8t56nIxrmifZcZPTtX6zJPgNSlECAVd+WYDBvtEI2N
I7GIVQAhz4ph7lh1mWy5lu5Lpmkk/XKwk4XwNeO1m5I1E8HczGC9vLHu8W0G
5py/u+MP9KeNyv710KfsHwCMxld1o9FLYNO/G15UOuYd3Zd5YMGb1GnTLmIc
CiyJVaOrQym4vNLq3coBAs+RBvOogDGn0tEW4AqozCVXbxfP19Z7fz/n8uDn
OWCRvEZjQEJpjgKQGWaYJo/Anzzg0shTrdEz0CAlq1WOpA/ppVY9DRhd1ou2
h+yaN7eUMnp4m4S4ofaNTTr8++zuv6pOXaIQskjXyaY5dPK0Wb95dHvfw5V8
vTzVlmCDlqtUu9ViAquEQn9frgTs5AW3U6U8gpeuoL68xeaHKr7OZXeA15Kl
LvXunC7PpX8STtetjmE9JTS26jJZnoIYABHs4D2GQ6SdFyxpCV1Ar9UCYW7E
bIHeZrpDIAVou+TX8yDN2hqx2jRU78aYKBJeEFmqq5NSSbSTJb4D2vm11iCE
xpR7c5zqpmK9mw8KKp2jufQ6zTCHfwCqa+gimC8ozBl9vzKSX5kQ9Lz4yrV5
sURMEm650j0sT7e+nS44r+h0xq0cx7IqKcZKjDG8lp0lpSSjRQc/u9rD4j6j
nWVhbgGcuGlS8baixJuavo6bX3zsF2IxQSFmJjjCEK0IHicHQrQ2mvA/GVvg
M+9+5m3e/bcS1OtlyTB98qAh6khWalRMQR2+zDkKGRHt976yhTD7HgSoyrIF
EoGDZUz6H91xqMWp3oEZEsY8Z281IrwB9NhYYe5AIEI2WSiFutPQEvpRnQFs
Lzd55G98mzjABL6Ilii6bQ2EjR8y0vNdLU2IggNlKv41Dzg7JowJ4CsjHs9q
riTpDYp3+Q+34f1druUtbGC51eTAQWWetTd3MN9+ObgWl2Ud2HJmTFa5HHa/
HXJC+LXianchDDL5ieu6WT+sV531V8/kPz4h7oWnLb3ax4engzFewtubuXCm
MHe9ssKA46PAzdBZmL/LwsNL7DkwC3Wno9rD4T09YzEwxis3NerVrZksp4Km
iPwkzS0BTFjA55AfLnb+e9y0JoKQD+MSxqjE6o0YKNro0QxtIxP0rg41TMZH
oFjgrUdAo0Uz8BTI9VyWyEzLFGk/Cmy7IjdqDK+/4AcZ7RwhpEBIlIDZAAPO
RGosYOta1R99hh3gP7/+XKpmBCDjP2C7CsVGHQebEyWDAMz8atsxJT3nm7Lz
Vlf8A8BpsRjLpx6VbzMdOfQxqShlbKQYQVCitmRx6emGujJ9Ufnu/HdMqpPC
xcNrwKrMIQP+NergoYm4EZmWCzU9aj9EuK+2IENPmDOwnYkiKlSO6JDu7bzG
Y3lsdEd+maKytX4pnbOpv9TeZUgBg4F+arQ7w2pw2T8oPxa6raCjI5nkhXTA
pju4R3wuc6XRjys3fhXcsawB3mnQZOErt560p1sjtcXSW5dr/fZmvX9oBbtQ
b5oUCDSoWlMfMAF24w4nNAOETKZeEezAzZHtuLCV8AZFaruIroeQuzM+lEMc
O/F33XmbunpERjNS0qaHlUSglTPCn2OFJIZgZ/4GrwKBQjPJu0twE/9+/5Ej
tMjX6v7/f+qABRTRaRpqCwkTDhsdH6rTigRo+nsKBnYjA6TrtyWz6my5tDRi
PjBmIfFYzdEmaecUAsTNvRxU/9vGe/p+qQqUc7pcgHoUDlstaQEW/YbCzHCJ
3Xjmef/s+Gfljm5oOX1PNKlBq+qrnuGWUaakuv5p1PpmvPt40kK+oYiK4CQ6
y8mVePcstBqo6DX4PuLTB3uHzyRCFVAiTE0RNnq4lSnWDv+f7+CssTqwNDf+
a1MiZe2e0mN+F7kaZkIveCNJ8e5DMQP3oW2wzcQS0d8fcLpL4Iqm1jzWst+o
0t/lTFX7e0tg0kdErvALO6UMmGZflgqWPZC/nRvciycqFMeroOd+fdIYfcL/
uasD82Pp/3Bkey78r/lL9IA/98Wrpj5RBWwhGhwJlYPjQAY+1Q3W5Xu5+VRj
beDPyYIFeBR7tKqY2F0zUNvs1UZCtrjg0FqAjOEtsVopqXcaKhO1kpbvLUb7
eV1XtbCSy5xKVkFuomxx19wUKXCVmwCANq018xza/J8utoHCLF7IqiGv9YHb
FzddaFBZMAN8NBO+PyS263ZzGolgaFb0i5HDhP7ALQfoXoSOuj1W/yD42a0X
Qn/H86Z0K0EVOyoWqQrCIfJrHJ27jacq2gupfOENJyB1rULaM69pe774C7+E
0DypWZIU/aonQZ3Qu8YwTDQ98PHdoObX3h073iuCgRoeUtaCnAE4Bz2va/66
wiofYD7UQ/sovVJUAd2KcU1rfPzV6CsQEkvUciyu+zw4rm/GkFtKa0U683uT
mgrsFZ1e+DSsIqabIPw2GAQ9fteCve+gh4HKtq13+XmNlRoa07FXi9z2lvor
HXAaRPvhI+rqgQAD9iwzM1Wiv5H1dlEgAWjxjvK1AA78uV4ZQ8tVJBcLWgYV
DW30Qwz1v0v3tfQfdy19ZTOSFSowRXB2vj91x7H1bVMASmzkARSL1fGYMA9V
6mNeXA6Hr9mlC+hu6NJhSEkcQkOAKNVK/OOUE5TJ+ndjS9JB5nodRs1b+htQ
amryfHJGBMXcV3gL2pM4zpt78q/zUIO6+IApQGatBjUXtVNh66sMbzzOGAkN
R+QYQhSAC28rC3h0v2EM1jSriqLq4XW8P+HnCDZBRS2lYPQmVaDPQE92TCUA
n+1rE4ZC988+hYv9ptBy7ruTUKev+yikOjkoh44IVKTy1RPokq0LwNzcX/N5
lU15Y1rq1q9z3ZNeRDlaSyUAw/kZM+mU5m9767MmXa9Uh2ttdqCj84xstEZr
r4sWq5uasqB7JEDC5Uj8Zf/LxS6Xc1UoTYXj/Byki1GCdcaOmxaZ7LtTcT16
Ambsw3x2bTI7j45lcbToqB8fwtKThdVKTarTCM3GUuDItJb/3Q/LuBVuEP1Y
ucmIWx8Tab50bc28tfjga8MeFCuzd8D9qP9/bo7HDUQ5UGrzn1Lnx0AIFYxu
KH37aMfpNkNKGmhHBdEBHq36PuSz9Eqad77MVAUYOhk1SFrlq85J4aMvFAOC
a59D9UB6BQ1KCh/biBxjL+irP+WDXhhGbRrlu+OZdMY8QMmUwcgSVdJeDnw8
e3oSXB1N6NTZJoDguBzIro/Mulk6BzsrarLsRcnllkN+BrbaZ8iz7l8Qnr3o
v+PN+j1XS2xtjsWUICaL/i5JQa4jMq3vilVsQt7BAerBNjhmwHTPyH/mhd0J
DyMXdP/ZZFtMvoSgvuH18ZS8z6IWg2rxf05T2/dm1FiwQLryBqly3w59F5Ly
a0RS5ahcyldF+5XG2930tRbH7XEAWYvv+McSAmqThgXsj3nO341ZcqosGWNN
wSnE+D9nTNXb3iXP7yJ0hYihsu2tAbKBTaLVuw9/jVNcYTdt6x79loEX43PY
bBlwvVQ2eelxuuqpbTwqr8PNIqjHmXwZF458ikWFyGxwtDu3eTUO8cADoHlc
dZ1AWc2woupZS7dFzC7qcJlZOoFDZYIcu+AjRjpMEhFYuW99O1BY0RkjQKhM
nfA0lBXQgZ2L3cg/2fKS88UNjLXU4zV0sqZVObMjsK+Z84QOgUNfpKqxfBjO
S8+36TR7fj3Lcv83WZ1TAXVKjdxjJOa1tpeqEEDBB+XsX2Nf8BOOkrZE6XBR
0atv4nLz6hT/SslEdE0raoNm40bAdtmAuzfzROr1vbp4IFWjLMmwaGg/vgYB
eYvdJS460dtkLKIGKXyfMcQEnzqXmhCGVYX4Syxmrj+Vzbn01itTD/FzA3mN
GwSHfiYG3mO+F1OYaNBQhywB1k5PXO1W/FKQkTqJeAVhpFIIuyf7OgggGnSD
1Blig4HZQDyznXLA2fZvXvLP4toD8tveZagbHXPBaFsp+M2lJy6fwUmKHIo8
jsgoIG2TruUYT8C+swT+XLjuWX/xZ0v6S7vBb+j8/H62T1X6DslvAzELtc7z
p788tZeGvsQLVipqL7JFPAyb/eaiZXTnM7QACtu8cYOXN8RZ79/WBp2Y0zSl
95xw46dBaTc8YvQOnEILAZvQ89qQlo+geJoi5BddpTDzRej3JvfxZ9FkoDKh
rK2DbqJkRgGkFCizkKpIGubikN9xPtNLxTRbY/mWqd3jCYneCVob+dxP4F4o
qoF8+CunKwyWWTq0mYSUZiK9cTd0P3HM6deFfn8eW9Y0ZCHXf5e/RNi7UYS7
sOySzm2YzJP3W7jDqweX81cySolB3M/ZL+EIPqixyHnxYJddx7a5nexzT99f
miskT+uoXGiGwfRfD0e5iJaDANJNrXJMO7//GqdEkXyEMq64A2+TSiUp8AJx
HWxz+D8xW2wqCCzylG35kijMcZE4KC3wiR50ygRdwXsOnz2SiTDduEkxiLm2
0ff9Nno7xVrgfb6s5Ry9MsErtJ9jyKkvc4DU3q7YJq1orMO27b8k+Cztx8Pm
/YaCyyyOzXSfp+a9HXcxaanAvT+JFDw2gLWj/b758iLbDqgLKverpVi/Kee0
mX4CORvooMKnTbwQpiSeEueQr2RFElLAIPERfayVHlWz6HmWgu9habBUFGGx
adb5IVU66Uatw3MBvRDT4V8x+iZSiisSn8hONjoDGOGTwOe2vHLsG8xEeiJT
1hXXb5uWAH5zwULBaW36EJ1TvgCfuUtnl8MD/AIzFCAZQdRVExu1zWEeup2G
T3vUOA2+y2v4i9ZYkiTekAMSSAZaT/pgCMq82/JjBQv0R24tW7LdKCbyZGlf
43gezZ1h8bTCH+O9uiitdqySccUz86WH0tgdGt+fpy+hfGGJNkQamGzTLxjK
GLQEd1M4fQLRHrb7tyXZGUq28xDMmaEl2gCxhldYeHuSmxS30G0+nRv8qSLq
CvCWyFT60Oq5OwS7jz8p87kcGl4wbbgo1Xv9IosWijBqc158Qy5FWjbjrt95
5tRcjPM2SEMQag7Y1eFwheqbdDZV3PyHtiYh80t7ZjPvIC1k6GCAstjaIt61
XFGjBoQvJTRtyxGVxZCoFVanPsBLb2uhbF8UX21ghUwUTp/0NHvuy/ef8HcP
gcE4XtHdmL1SV6vEKjnOVlbNXl4SbMtbdwLKGRs0vGXTagg3IeHRgvxCinJa
xqzoHm+GePpvrkvyjeObxh4rdDkg+RoXtxh+mb1cEcDwOOAVdU6jCVSW2qCM
dCiOtuxWlaJXkttkrHONdR2rMAqHb2TMV8Gcwf1/dTWbsnzrgA0egWkgeJCf
6yujz7g2XPO0Fdd4jzAZ2NafRjC/VkkEbnbw17R0nwRVlwdJsJOzG3t0mYrE
tbsrRB3d6RwL1hE/CnfA3s4kfvoY+stO6b0vot872J91peNOgQ129vEUbviu
EObylPU64nI3uC73Fzz6c74vCzEkiSkHdV2iL08sz+ojAgQQv6FJzx8BVAga
EwbQINAEBHK/aImmY5KTuYDmTr17Uu5ORDRVyxUp+g6X1Aat7CbNCUxF7gFX
333R6wKCtnHgDNUWRFl3Ak92uJs+xvgKtPbx3pj9LfFVQB3iEP/7cUOQDSNd
QZ8zaaVpqHp48fkwsieKqW8tDghCyRDG0xR/Fe/t7IlGpr6ivrzdKOy/jkcx
UxusN3RXnLqfSDnzQX6IZTs6pISwcZEhKZaLTAdJIQBU2bqkYiv07bw70xAB
I1gZkc+EYxCkCiMFNUj911ezclgvv38aoHlhw7wLGX6b2/UjDUl8g1V6/X/M
gaWb1vDnofztR2CgXDel2jTCjVYE6HhwecH1vkRxWy4UWWxBDsH1OX2sb4mU
qohPuCTFcW78GKxdfbB9r7YfbB5p3KmidfysC1v0sSu83IpXj2pUtecExlfx
y9GNE+aUeY0t9jXGBJm/KBBdtuq5wiZWosbq82ut0/CshdHyAoQ+Pl2iOstx
x3IoybawZNdglZJ8rKTrYwk93Z3XH17GEWMkRgsDQR6CwFqvwvFm+4t1qJ8t
xhQs1b1ojdfMEJtkZZ7oM8Mzb1VSs55viQhwsyBlQM+/wtiNTP40XLq7Fo70
g8BNSB78qdvevt5yM43Vvsnub4dDkl8Y7khFvTVCsGwgKd2KMegK/uj5B+Ec
GIfbBSqeYRwleGdn5GhoNosGVpbYtBFYIcIEHY+YRfc1/MKa7md3E1Sy4A0J
mOP8+kZLPk1deTxebiuNSHOzqi6tvAeMQumrx9BY7j/IVuitwCVpJI7DNqxR
habct3LliF+vi0ZB5UFRRFieHyjAf1xkTGIb/4Aber0ne8guG4UYXAMxH3Hv
mCcW6ABHLcDWuOgKN3/aq33IxAmBG+tH/T6cL6p4aGOTH1QZjiN3uWdwWc9L
MR+znFBQiGNJPV4bHy/q1ah18k4+WVz3AuLsEGDqivuMttH13esvZe+WDXth
1ILDjnbHNL8k1Po0M+xVQ1DvnZJWBe/VvtxS/8i8jdtB38Jn5tawn9LZXSWJ
nuUo6T10l2yUJkdNRg/9+wsgoRCHYtaV0c/efUE7hyGKd7MyJcMam+uySE8p
bjsnJxIpbiRQrp1+wDgiy0JMzyplIKLZgDzBN9vVjIZC9SmgQZ1XQpgBTWhe
NZWoQ7ONlFBwOPRbzsABIfO5W8LS9ztpvjzeIqLQMEFk5LVjuwxLAQaYxJC1
5LtzyaVCI/tVTNrXlB5l2TxcQvgyxBfH4KW/xCihiODIMuDK5tzgznpLXy1n
BZDtEDS4tPth1QKsHSegOqYGIN2vsLYRy738yh02Kq1lGbYwfNp1YNrEm3Ak
fdKd0u+CLRH1v+zr6MxFOXqb+16QP0byqfzrQ7drKMqFMIuaO3mT9a/vUnsw
ViJM0Z/CObfP2QJDoGnWRDBXswA7APLatkMUHJhGwfS+goaEl+fl5h78W4zi
s6dfK/O1CpQCnUdfUwKJWiVPsTVJs/MXXlz4mtQPDxdMvOkgpxsrN+/J+sn0
vOsnJEuFA6UH/WY6qhVi3Ca9Dp42Q6fNm0mw2VhsoLSz+af/qdd4xYIC3FOl
WVMVgYX8wjHCCcKZmnxDnLn10sj7s63CqMVEen3ZNnff5yYR9d7JnGDyv4b3
qauoFzQiwYdxUbnShC68+XGzlAxysUfw5LjO7w+ZyoxADph50Q3S8jDRPi9g
r055XXkYQnjfBg5QURWe1j4VayIsnYiRcrVBfXotLUxJgzV1VqbrdUOqvHoa
n5EEjpQMvWtTUO2Y5ZgpIF46ly1MN+NoLB0WTSMp1gv+ivVwlGTfmZI/LqpB
qMRFSgUfQ0lGxMriFPGD76nAfhEAsIYMTon59aL/jX8axkIKlShL1B/CcFgk
7NmWImS0eWTRQSShzPQpyzFMzQ7WJTOupQZKR7c+9g9T7VgGgkVPhvQW2h+M
X1APGKh0jRUqNSyqNveogbkrcYvd/ZdXj4yBsbe0CQp0p5ecKvvg8dXx+gI1
jj0zutNhucxys9+dSpLYtej6OfS7SB8Lxmq2PVY4ekAG6ajj+k2eysVXPpCm
XZVQLpQPyqQmiTNFQhmGrwR59NoABHdg1DXTF11CQw49CgE8h7KHCYfxkD1I
IERrZmCxAMtGHtd8urpHUVjIVye4wgKP1qPh/GcOs7R7Qs+MeZ3LQ6VuU8MO
8V+YhfgfLoIi5rfGC4V9BZe3yY2cgEtZVHAu5iS0wOaGUE7F2pe5SvPh5b3D
zOPPLrApAlN9eeL91rU/GeoU35W8VsG982KqD1+R7I8GD/ZMro0LxrLdnBdt
m/+iej8O2unhNP5+QJ1SINzvV8ll0+CmedDpQklDQ9MYfGYTiPMJGxN9Iu9+
2y/7BDiOU6qvBkQIidMxAAVZQXb8m0Y4jvB33lYGoe+DUAdUOI8SJAUOlP5v
UMnuRAWmS8icFRGct1jGaktRRWfwc2cYzp6olmlCzLwZJxpq/pNEAajJla/J
TOzSEchtxXFYXKkhQ9MfF3xNg7b+eOqe4taHZcFUuChXA+n9/AadD2YsaE9N
TRUSgV6u5XyX45UqQjeG/eYaDicahcH8YDfMo4Ln4tf4WV2yZoazP9Knl9IV
dkd25IQmDqcdLhAi8l9QzTXKuw+JGQRoXqUY6T8R+yy1QLWfFLYg4BsrB8jg
csJj+pXxYgaDrbZpmdEnuelbaOvvIH3yJ4qXd06AqKohaFxkQDdzG7JU5LDl
Z75OO0SGh6ejdFTcJZ7VvNYny91EKx/0KgNWOyeImfr/MWxo/L4zlyX+euKP
HxAAsbYkcEiRiMXOuegQyG+pZM4mSUTjEiXanMsB40B/5Q72yYIRwdTE4/qq
EXJlCdZ1qVqbFLcpg7TQY0iV4xCI7naPEJaZG341eGdfgYdNg9kiNfGWyq++
Eoir/zLBnXWo/c6aeJFLIKkAl9MbTFWUxIsweqKMLSKf4AN64536HiBn7wwY
uDPc1iwOuAkeeDjc00TP2AYoe9Pdt8cRPr2xi4DyQBWwWPuQT6336wLVulvP
mnVJ8GXdrshFUkOzwDnWACZwZp5/IS3jtvBKDD1GY4ZG/Sezo714YeJF1KNX
sD90pt0opWW4pLKoyxoGHC+GvwDCC7sQ3Xah0Ggrd3QrP+PZHdCeuM7yoget
MfAyJq+Eq9Hrlxy1/Bseqwn5jWB0ie/otzxeS3kpJ2UkE48y0+OpYM8MzT79
bicn01QSDrVXKmqcIUNca1bg99FEL7STDQM8n+ULqoRnASBGBnlb2boetYlc
Ee4m5oLDPbGtfMh85fvD86aNflGWFq2xSiG+Sb1niy+4xCWCxoXSWmrMq+4M
k35OQ2rdcQjHs+Gk0+DdptQHkv7u2Qj+/E3/quk95XNwF4cgQNNQGrkGcq1C
22t0E5td806FqCi88swyEsYEILhQiGVgbG2xiyvWxyUs2ztEhQPD5zupDGSs
UqTIyv5djMh3ioWzVTFfEzMtEnb/ahc5CTjKuSYjLRClM2MQZKSM/9jfW5k+
D4Id5fPpDlnTutSZWyN7Y8GL/4agC7Jl/K3gB0yCWB4TRr9eTX72ONzospUc
KSFV+a9LKg+YpZ88Q5+2jdSc0j4mGd+II8r5Gl5+tuANQg5JWwrJ57hfCeB2
xUU18jFfYSad5dEwreD2U8CKrRH6qhfe3ETbCzI1o1jQm6FcaI0Z4OnJDLo6
EqqjM9rGImOyLR2mccPgMdRpZY8ZB9SzWyInd2AI9dcQnp0kTnr5PgZMdU0G
IwVIPbhmrqm7qWbjVqhHd39rpOghZc+sUM/WQzARepJkyFxbKgLdwDAP6vHr
HL6pP1njA6IyVzIp6AGYqwJ32/gtZyvA0JLfC3JQBeso5qotBSINzaA8G5yt
DOaJkEenB0gRBT7Ma8bLly6IUjy2mNaNcX4mlP/6JMWg/sj3cLP5W4jfFVE4
RPi/XmxZ6HonO5cISKx72uVJ/ak3nkSewFEMfmkjV8mFO4YX+0p+A/nPTOaV
92noc+kcxnkfqioCGIZsy8MUAjmyowZxvYgsND5eJsQoeLZTYVl6tHrwdPCo
N/uQ3EPKMQVm+Tz5KQCkMvXam/hJ1qjVYbGa8aRUTtWREguXhJor+6sY/1iZ
Z3KDdwvUNG0c24VU8KPWYeLQxi6iWpvktpkUNH5Z37aku5EC+15QVICBtUd4
5l1XyjMrgSkBr5aWyVfPQHLtsaiZOxOWjZPsZuYrXZzdTl/nppDriTreQEvm
qaIKVxJB0sRq/j3NbUWGhIJmGCS6HjbB81WbmwWd/isostZAYtFvDlnGPuyA
jv+9n5kA5dkMC3VI3ZMfOFCc7hGFa3rKp8yQAT0t4i8gyuXnPLjh1Fpcfw+Z
hMJYQ9TYnQrsc+vNUbHt0ExjKb4R/3KUCXU0EOauoraltvwaeeRi67wHz4Ez
QpR1jR0HO4Q9yfhuAgCJYyiQAlinNbqIfd5ZV/k7mNotJIOyjSwoaSWnHtB5
PibmHWKxzL31YXOiPf9fmSQ97heSErzdZzT1rMrDNhuwsNWke4Sy8giJZoe7
pMQLvPB7fSTeV6vFZjhYXI97EKgXjI2Wz4uTNW7LvlvvjAham5SP83xQCWrb
oX2khdQar4gJJ71xKq9w8LDXuNnjWNmTI+c72VLWO5frz267XCXIpDx/armW
3sI8Gsx/rYOpBmdISkB7vxID1npjm8esNh/lZBQ+65Vov3KDRr6vpFRYyAlO
xxHu/e8cxZn3axlBZ7O6EEQwMdafkYOvg5xgrBCtgjG1rrn1uhYm8HrKtJ5A
8v8QMPB74qh3t3rXy5LMGoQdH1dLNHaLpcqf2lmmR23gDCCmG6WTdWxLCgui
3FI4NlhYKQkjy9+SEAxyLoNLFtXsB73fmor1GJSSJefdZk38OpmrTl2Qs8ll
vKYHe09laMaW3JYWnj8WPa3pSoB9htv7lJYgJKVE4OeJKFJ/0moS+E+6T6JN
H3u2UAM27vmpogeeK1cXEmmZxQRPe+sF54N0XAeQ3h5fVIVXI0qvvoPuf44f
GgP8/vCDIDEXxKli+vJdqmqHJEVFvsCspKyF71zKY/Cven276YsO7b4Q+uMF
CYn3AmMijkvbFWuTrHfGrtCWj24+jVRKAGLIKiXBv6ngZ1fZi8eO3K8FjDQJ
Bok6qRLF4ZmMTZ5S5P1w/AtJ/rHJot9sY8kChvrySEfgDY219s6BIoHRElHE
XKy1C+vKh0e3WpIjDjiUDXIdMpXXx5wrMmoUL9+pA9+Do54c/LpZbTBsm9ZB
516vaAvvAnoSt4WVlsx0iq8osLrBzzp61rvrsvikrT/msVGQiHfD91dMoNiL
NYPDK2isI0IWBqw6+w1rFgh01Ifwi9NlyZ/+B8loPFZkVs3u2fStPNaIdAmZ
kuVI3VVvAqWqULWQemlWU3WrnNeRq33JlRExxYgNBQDG98nXOOwtzgl/yZqu
Nhz8YLXALl1nheWUsDI8ovfjr9SMmIybX/s7njSGlbFrJPJveQUYSt/qdPW6
PJLZyoaHTWA0g7yRRtaAE+OqIMKRmT2u+abszTS6KKLqNivx6rN+7NLcU8xI
SXvKcS4DBZUeyuNDlSLP+2K0zvhGL7ub+HiKXBEf2w/NdNtbcQyYfxIwWkof
nnkQg71fWouysROrSyoc7Psddetqd7QbXSEApUa6C6jsI32aMdErX5HBzD37
VGh/SUg5vELHqPZFXtNLiJuVRiU1CrTMac0khBTvxEoJjtFdZl9TYZVUXl7A
u6Zphvpukft72EgkcUwcUqHuxM8YZOW5rLBjy11NGiZaIpHKw5s0g55p78XC
yE8dsznA5j/YAuFS3HEu/5dDfUXwI8+zsf2ZppTmuWbDnsAhR8aHiM0URo3L
uBzPXS3ZhXKgUqIj3Gisz80SXHFkcPGCw9BszywU0zNLm42JQFab1ZB4rMsf
ns+hjfi2+R1FEZyU1H/MXd2hcSeGFcYTY/p59WX1NFXw4qj7DtaYxOIfotTz
/mOqD7mSJRX//GMNRtjzBVt33sbjf5WHtFZ2wj+7gkcI96QrueSzyOxoH+hz
kYphyLdaP5HribVQi8gQXcaBeVC7LfM5thSldtcJYZkOFjxROI3/vGvHSmB/
m62mf6FLR4TU0/qzk5SphzmBs5Ex4y4LZCDn4x1PoSyd058zSmO6PB/AH1Rh
6G9dkC9XfUS5kURUSQGvZRd8td9Ers6d8/qHCaBpynQllctn1vGziZ+AKVsi
6jp9E1tQDCSPh4jv9q4ZTyEvuZVmqFWDKoW7IMMmpyjDAgX04neurjAsesFB
MJB6ZDCdylroBtzI+DZvLqRAbsBX3Nq2TSET8xGB+UCk6S/nBb2Awb1gSOex
Kc+oeS94rCMOad8kMyPjVKbinhsj8YZrtDMd30hwZnzC6oPZgXgQle5vyKdG
JClJWfChy4hhgPargGMxs9v7eyRMP9kzircUFKkVLFWkMec3oBWOZC8S6Wd5
Z49UGqvH7xzhpzc0o/rwD3GW/mcSETRcMTtyHOgCTUXA0Lmi4A5OweZRSmRg
oET4Fm3qiJhIa+QKalHCZ5fiXFeyBWlDCXxkHjUxE67t6XSvAYUaMFIuBdiq
yM88JYy8agqA5GB/7Cb0WD3Y7kYsuSr4LSZ0mAnFi1enaGqX08BSk+oxjX2u
v3n9yJFByuH4aK+9DtTodENNR5VSZgm3i3yF2/EmFciq6UKLlO5tabFUVfAS
Ue+I7lOiySaBOE3c6IJTLUt/NyMXO1rFF4wjlTIZ2xympk9+Hx8Z6ct0CAIX
umdQ5JFjat8dkvx1czaXCcHeKWJs15it/V7pYfm7c2k4VkP3zN8pRU3KSoMr
jrT+G9rj1U/6wFcMfQWIajNyd6fZN8DmWHr4g/Yf2eI+htnjbXV/dhWIVJof
9BMr5z5Mc+FZ7d9vSUqtN9rJyqN/pzhq7ZeuaJQ/lmtbNZQ0TYtfP2F5htcv
+CpGp2wYjt4HQonm0xLyFBQYmoZ5W44kmZh9MWJ+cjBEhqUEU9dRWV7r3vTa
BQhBaWhkma8N/G0Kx5R0B4MhjylXKFO9ORdUusixNKOAJbmmFgyoA3XAoCgj
Vw7zDcqDGeVdzczuTTrlkUFxuVRyrxYlCrHNcc/NicQqujnl3BD3fWgGLgnR
mhisozXuOULZetN0DGmHPrJN+++3+EEweNEdONqyT8zr8gj8PHPaBYN6hA6d
4vYRKmg/X1xQhTaf/Mgmn0QSQqHq9C+RIp5z5BLQwXkgNqfw3KQae/fmC05+
sUKvbuaPBUcQpJGNXrZI8un6WtADV4w8EwGUJuTOjUN+gCM0zJqWveG1S4fC
Xu1iB1ba+LaTyzb1D8vd0SeViP4o3RfzdoaOjVXAbPzd0B0SLUbf+2L9uR2Z
e2bbRtz7Ww6RZPP0yBJPi5Dt7/L64WikbYrM0UFJWcgImZvZgZuX1cpo9mMt
TpVJ7wWcUWVql/5uXBR7JRX+Cda3wjDbu1TAMAaFD6E3QhtBncJN9bL25NtN
2JsK/w6m9jsbWbQI6ZjvwPB6YtcsQZ/C1QX8wpU0OUTj2PpbpalSIKiK2gBM
uogxZv7D0w+f8DxwMBdAY0wFGRPrlSU2pvG+6xmUuZJqnhcvyg88A1GEr2Hd
8eGPDywdti8GPm9A/LfQ8UdrHv31s7AfJ8Sp3CpLySYwB/t8lY4AiWaQceZp
Rv5tNfaMN1UQ4geTg7HAAB9uoYv/ZZDzrC9a6SfJNhJj2wYIyaAuUPYyyOoW
plIsSStwcYiEobikbPB9pWLBLXtHDbXZD86kClBJFh2XeBJpnBm9OjQPVbI7
0MEwuEfsKlixD+zuwKtMQielCPwJNybVpUICMMRocl9ut0h7ETvLfWXQh8N6
LR/NCPfbwOgcTkkmYub+keGewgKTDA+950UHMpUNRJteGAyHsk8b0tspy+kx
FDzGT1jl3H9yGsh1rEQlHdG/6HweX4HL8q/saI6UOMPv8TKSFLxDZhhViwHi
HEsQ/hnDQLxtoVraNlO/UoAYRiB01/mW9of+Zd4/2iGCuRBi88xhfHao4fPn
ALT9wjttziYGqG29Nd6QAYYmISObHXDiUlXu1N3ecJC7V3gvnU3VytjXs8Fz
5o5btzlyTc1kMee//aDz6n8mVNkN3Rskr0IItnSK/Ay/+M2LPB7quUv8Gcuv
p6LYmikIWxAiSMl16nF09tEXLI4wUuW7e/HGXn3G3Ce6ecrHGVSyAz1Vg7NN
MTP89vkJgtp12KM+TuihWBiTtG2aOlBAw/6X3rEIquFBKn3kXThN9Xcqc5UH
N6YSEWsH69K7pZXXukiuJy+LGXwp5WO56F/tjP/sfqD+qUb9hhxWJKAt0OUd
xSrUR5o0vyFOYuQx8PIZO5t/lRk9KGeAnLVrQm6ttyeTMe8/0fNw5eqglPHa
CwJ6RxmExtpviV2j96ajm0/a5eaY070/CAyz8+zBKEBq6nnqdBRb5im81njI
A+uCHyC64OBQzpyZRb6qHHZUXeDvaT0bR46TFOapQBPhkPTEDGsUlTcfl8zf
apISaaxxffCHl5LPMjlt2JTjNFkSycYS1arWvlOC+iKZ0gQjRHGOwkslqP85
rLAnIm+34vgB4pVX40e4pkAh7ftcJxbW4H1YiCK71hNIZfE/3SuIu5Rt5N05
azXpCzJ71NmjTxLX0mEOdywDpXIBnDg9udeJ+X00uC7tTmGh82eCJm4ogksx
In+vi9CeM8LTyNpOaQz7Un29z04COf+Tbs8UtzobXwMaa+giBFJbmsdHaEpu
YtS7pQQ2CMh+akiRx6BJE59x5z8WQYIYKEX6LeKHaFmThgmSJ0+67FsHFLT1
GPV3nqLtTW8EWd3ho55E3ui8DieRYoABKAGCDYPJs60MFLYIE5cbcx0J2pd6
v2RNbIwQItrOZ0J+l7/7cztoMZ23WUNtMs/KKUtmTFfzp2+PH/dePwHpxY+G
7ag+UFfbc0f5s7DDhRkG924RAciq3xB56qrTFPWi7HoJswIsUKizou4qF5bv
IxXKhnSxzGYG/mPdhy5+YUN7aAjbGT84YnQdmGebss8s2LMNITeRAJdfNooE
5YDz8OWBRkCxDXXRqwpT7FiMHl9fm6XOH3Y+pmUYbCEaGx4vJBcpaNVcMFJr
CtdpkanUQkZ0AvJRlXk5XsSK7xtUEvsUDncuLAQZrMVzHd/oUP55wLKJ92Ek
u/Pev33jYq7f9gIviPHmoo5dRSYLFm2CCisHo2cBAwIpEA+p1XrQQcyFBeKi
oex8AEIck+biGw9u5zmM/Vqofi5zqjg1v14bLA3d0IBtw7YIbPFqU0ojhQz5
83HIIs3xD9xNCxDgR+HkaA2SNfXBaYZLPFIxcB3gKgnqI4wsqOmyEf9iBTNZ
bPATBVPZC4EUCIH7C1jHLxb/F2YocOFcZljO7lmgmrUKi+nVaRc7Er/oJTx3
fWwWP+PbrXKtgqblz/y9xgiuqU7x7hn29N9wijFU9izY25jkUBFWopP15hNL
8PqaGYL9+9wxRU/0SY+ylPXCzEaCxmFDoDI6lYWPXexV2do0y6img8b+HUdq
lhMfQ8U6FZfdDur4LyZOleM5Da8znEpqE+pQG/1YoG82nuPI8U3J1BfFQEvs
U01Jiy8uvF0ZDs3eHlkuuWyPEpYdn0ZKvIFENz6XCEAoAr1XhSx8SlPmGXIo
eWPFJCYZ8YakH+QVd4BpUE0hoq/XZkdOvN3A3wmEsUOFwrlJL/krT1+jdkDQ
WVpEfac0S1+LtqwkfsudFNTlas5hDeR1pL1u2HZY5ECUA0j3p+1RdGbxjkOv
QyFql1TsA0zielO6aeMGIfGn6NPV75mpGVRgp5kTKnAcZSjd8jtM8AvCwMuq
lTwZnjV3E53uXHqRW5hKIm6vSqqEqgmRXVd9UnaatUII2K3CMSzJRJF/eMBr
I0h3BUZ/hj5ohIrOBEjSprx2DnQs/trdJ/WR8PUAC6Q2S8RrC5Bj1ZXII2zE
vsz2Gd7MXh81hq399JeohUN27ymn6WoGQVo/5SPeG0dz/PAwg9w/76+3iGWO
LDce3wo78FStvSAjTGj4tK7funoKEE0DgHUv1CFAi3YoztIZcHzOljhUhYqn
6OCO16dRV/tTf6sahY4/3zMdROE0HunX43V0iixCpLGcu7dCHjotYMdE3ujG
4hpe/1aeoy8186ArAHWiZN87VhizTubkqBy4Kxwrrn7+eX6QsWllITkBk8yB
e3SjfW8FH4fBbbj2h2pmSCJ+oNO9lieXWAHkZtp3ro/dbL9U8ofvaqps5nqU
58rGXecGe5OlSe10v5ukgkLsfnBliXFfgAertWai3Hg+Fp076iJTLV73WQ3k
+LN/tPMzeLvBkZzF9uM3XXYHzBlUdWzQ3jhR48WypSgj6b/5PV5yN/AJRWFQ
hHK/51mxQdsxq5bOKndMaOPFqyD+2AMGhQJW3GAKAhqkf1slFdBCJAaLNGCV
mwZyvosJUSZHT92cdqEtPjUy9DIJ8thCz2VcDL19xWFuvdJ/TWO1zb1N2mmU
k2Gjkg9wgEALUyX8GB3c+rOEJecWPklUuGPXVVZB4R50ngpD4htbYQaGMs5U
kRQeHcrcOP9Pi2mB3edjCAdOx6P5KCHQimn1FMoIPS+FQPmovDjBx/x3enYP
dZurKFQBIe+hFZJdkQk2HyXTrbFpUU9CQmJTXQo5ZFcKs8pmsOKDHEfZ3EkC
qUsWl3g75YUPId/qH7Q0+SE91nGFvBnLY1KQE4MToeOk/5VxjIW1dFWimxGk
xx/6Ex24tCa0OdpGyIHNpLSsgyPJOPkLswzAvRztmhAx8GSFNwc3Cd5DNJgd
YTKa5QrtHNXwDHar0S4XIpwr4jpt5mn4UhJnDcJGAQCIhLrhDt4+ExnxOl9a
uwhePpahjMXTEtCYiquxzmJBq7Yv3OrqdDLrfX3K7ohWaRaVilPK75KmX+j8
I8phdnODzYWektA9zIXDKooTqOYBxjTY211ih3tmsq9aYQhdjM3x7RsgpTaK
zT4VehDqX+5ckkXX4LRMFhS/pc729OdKdYVlMaevJW3IIRRBWiNhvdaBS7aK
yxW1QcLc5UAT6AXTmv8YTFrJgLYO0Igt9wrAFws7VTv2iKkhGdWfZMhIJgfE
6fSMWlX0HY+kw7uffPGawrJ6pNKu4P8bo8Cxmzp9Vd7lo4WzWpWhtwA80ifX
1tgYgcoF9LVJ6Xf7IdPStAVN3VMRUNjXrMoFwAy/Qx7NhXAlmRlaPkF6oNkk
l/lOuc8sCyxmK4Lv6eQPlD2b2XLBvV756iuy8L4TFD6pvJ6OZaKBJh5ZxqzV
KtRnsolYby2VVRxaCMFS8Q5XmNQ+EGvtCjoeyq3lwYXzAHQlYcTLVN/SNZYk
nD2omLaBX13+yv2zq8yuX8STvj26+hKSI58EngI/xH0wILts45rHeEyW2ikq
n0sx6U/MuCSzTP5OflmcJb721451AgpIl5CYIfm8hyRBUmebYBQKGuDTTZje
vLpNZHXR8hXNvlrgsjk3o8HjWOtpUUYONQ4mzep92X6uUJ5vzXxHSjROrD7/
3h8SAnnCL+xfq4XHTmLU+Ll3085tzDJCrclfgajO89TUiPhdtXci6u2wStiS
ovcBW3T7EMB2xRdj0jliy5Xvu87Z6+nJFkZwQO/RVrkTPXyixz1QeONkDSDx
xnYutyd57ig4XogiVKtX+sfzWfBpJVGEi/RxVT098xunMjwA7uKx0HTr+u9T
Hc8A+FocccP+ZEif9r6/7su15NhjjvsVz1W8ZVsGqvuKcd7bQLqggjHlOIAb
iMXKhtQPJEejdeJuVQCu10+/yWUAGG+Qs25IWoTwMxvwtkME45FwaAFywAsF
3yJbLT6ghQ7lWHuXv+bkxyYZv0g/Yn09uQd0oe/2sytWGAcgVXTEgCd1qQ1A
lrGGE85+EZw/W3t9ppcNlBp3mhuQkX8Z3lHXMIBO3qFgjY/dAVT8CDkUM/CW
1SxOx5G1qtKBtHtxCrASrRp0Iv9yxcVvrr1gwJSLHJxVqtsdR/+v+EwAq1k6
/hF4V8dB7ZnjZx7Kr3iqNQyc+k2YWj7ATp2eUTF23kUZykn84djOqNWLhtkx
bsht8ZNkfGqIwnPGa36o5DRhGBLGIX1hvZZakWoL8k8W5TVC6cEYgi7epa62
LZaBFgF5IZitUTGJ5TWgbgzQI0YUmfZLMnzHNP0wxMd7KE6LwEqMXMbJtvcw
cSqo/gE/c2OlUwLnDL7nPPYAq186SPPzrXCXUvL+Bx9HYMkVvMalCDHDIySt
/LenYn5i1FbzN7oEx8fLsgUoB3lz/tBhn5veYuaj33wH9CmaaugP/YhtpA74
stmorTJP6Tdcw9mCpgfQEFZdi/cm8JWLgc1u+W+TUweA5SCnWQK9gO0Xir0B
pYRv5plduweHvGnOU/xoj03l4fm/806RuY/oU3k1Pt6wDXryZH7Dp+3UOtdG
nygZ62A5MJLmbn7KiAP73tOWHbNNSZ9GUvkSx7YCV5t2+JWPcxAJqSKauu2S
CGisbvjGTCQjJJEF90RMJ37q1hlfMfpvQYe8+PcOBKkIm3WjJ3sHzoAQzGue
3oMAb7mdOnnc9/bU+X8feIwr6RKsgfeSzgKyQFYJOe8ZQ8iKNLWmH18HV7NA
23ZFTKZEwX5WdwCOB3Jy+V4V8gjigZmk4QK7DakUf6SFYrrT+LOzYJBcQECx
GcpQOvsqo+ORcR5+owkxgVGW1AR+zGoxcKU1YKQeeTus5SHG12xQJafiGLve
na4UxsPENyfnF3fvZWPxfON2OD8yO+zclYuF7jXGFASO08YUbs34hW1nLsQT
wY/182Hv5PCo2kHUi2EXoIdUJD8EAzZ6AXf90WTCdtYekvbH43Nia/zxmOkD
ROGG9ZEJ6vqd/7Q1aT+TPlXjprqeYvdpRK9CEI6NvAZgkmjaZ2fhTM/fbh25
R212n+5B2vDy/d6DFI81V2IY04x/737MCJJrtlXbu/KewY2wQNpw2UAXdv7H
rpH6CqKPHhsEf8oJGR7kttvxsQns3VWwMaAZSonEQ3Qs5wgjoeTS1POJE7nZ
Jxzu9nPmPwKqniTsu2J3cowwpd/DMIc6bC7fBGfF6H6dEx6U9nly1IamouvZ
eKONQcV/yel6rnocQrobSHkfdlF6WOYEp40C7TTztFBeCkPPSknaKAP313fG
IiBF8zs/682N31VXgiIdF5HLUSLCj0K+VMF2HzwWyADNSOOc0bxQnPeIGccq
2XQ0mOELCzPOgpsLvyfcZWH69jC/CzViNJnCdiek2O+abT7yWvBFRnpoBnal
y6IpceGiaMzTJZji4tUavZa4aYfmZRRuS5FWMynAwAbuwkkSOv/RzUUw8rCv
mHN23lJ2tlRVwc5Dxr7r+CJtbcO+vPHcOz4IwAE23BkUz/8pBZFIxDYmrfV9
br7ficTFOpEiarRMK1t4s5RZmUJ3qzbYYLCO4nAUA5IvbBK/4u9VDOXfYFJF
KPx9TjTB344vM4jzVykput64WARJfuo2uiYUxLbc7VbztJeptHzy88rVSkXS
CJrScLt23gXf/ZZP8uMrOpMVfaij+21H8elOacAT4uPTf6O3MbmhtRm9GTY6
nEu7Fd0PZkBFw8a51CBE5Md5YxEl3J2ix5z2Zli2Ncx/dwKS5X7npnQFR0pQ
Kjcdb35uokfkzVxUiFh96B3/u++Ld1sN/nDcZPvAB0Mb3c0i7ZFsbdi5rnFi
y0Ue+2VDTNIzqk2wjdK0DBTI8RKpW8laBNBxilYp/9+ceVyJS8uaxfxVyWd5
MqqX57AdCPs9lzC+jKJ1FQWFgfx/zvs2Z6UWD4pGBYequ2s4h4NdfvrK1oy5
v9oiqS7m67AtNZiJjLWQtdZLi/Ekak2ot3PD+durtQNBv02Gk5g9tAjdGe73
Lw6QOhiONCCdTlpdSL/MJ41rzdgnHuJHV9gAfFzw4n8vTvcwj9rHQSr6P0KH
7lDx6c5DV8nA5kUN7jjFvZwl3hZ28WQIeTZmVGpKBrpBeV/6yR2FCeXxpgKo
aWKqbyzmsXHy2SxpDOHBvZSXysrnLuV3kOT8nArbkMFe7U5MrYXa39QSbw1M
Qk3p0d7DaIOTmtrIcmg7GsfcOolKIiYCvhZLT4a3eaLgkbpBMGgu5ZXkGFM3
EuXIvdCTDoejMnt6cZeys1xBSSo9NM8MOUBKQ6sqOugbW5qsTB3upqmS3AOi
8TjIdEy0OxuUTpq/SB9hwBXIyak0nj2GGVPAvvxcl1zNby5ObCbkfFTXouYu
OFNQO2Up907N0STEp+1nXV+CwsQIwtQTbjngk4soab1ZNiRrqqcG3Llhd1jK
r/ESx6njLRM1r8r8PutzQdklI/MHL9xP5tG3h5FsPVM1wvsUqC8nWqEODEtx
5cB+S7LIlW/KUHuB4FmE2HGh/Dwo34W4A/cVfrLlU5GBLZ1pl5uSXxJviWij
iytSLWLCH033atib6hiIZM2uKQoZd3yatW5lMsthPm+nSxJdBrSWZnNMlXlM
grYee/NqXQQmuq6++qwTyUenHzJwYeZ14YsCWj+RHZKINjQZBtqhyJCqQ1Vw
ZK/m3QZf5UUqpBTwRuc1W4/1ROX3t+EHDc6HIOHSLq41Z8HDO78d3KQSZEHL
zwXupT2iTJkn8GO2rSuFayZSczZmxbRGM/mD6Jh6hVaLSTeOXnkDC7AcOOKa
4kaoh+MloOtdw0rnMkcltBoUt8fznMN49xGIvxu6TGD+iStfDXtyOKlLHvxC
WJy9xGRuJoKWr5H1NdX261jnWIV8GQbPq4T4Mm3kzJnLTtosZpW1DFZ/8sOg
4E2GnPC44hmpoWUCh/JY7XwpaVl6W1VsWTxjQES64STBAv9AEiqKgize00MN
Ir3X14NG8Tey73Yr9/FaYAtscgl/tAz7igiFxpghPa/AyVDxS+LqU9Qo6QAN
Wxw6GT0Iby85k2i+X3dKeiKLteEx4monOVXs6LmPHoxMp3kxkdyWMZTWHtNu
uXmEgUeoxrGqvOfrqQygzWp+KOhNSl/+UiT5TrR4lhx52wkw8QFJbLKgRiYr
IpJTx0dw0HKBHd0s4zSOQEL2wsyR7Y9JkhftS1CVrm8kmWgaH8DLMHrs7dcy
Fzr5myATcLDaHpCOmVnTp8K932kYlGqDCUihdJJCEi8EGwU4TfMhLsIDC0Lr
cOIZJ5tgHFfI5zA8hwMYvkP1SnUVJuR/CtqZI34jQp1xU0NxEUDmLPoYJD/G
xQHobGwow0eN5l3RA+DJqTOA2Pz3EoamdzACoZJOEDBfe2pb0G+4V78mriRR
FsgmBSt4ZPV5rzM4nBfTW1cmFc8LBybAKr2FWuTZ02NR/K2x6eyHCEgI4WOJ
l17PQi+sD/X/MzwIOLD+Dbuv2gtJLrrEYqwJSQihFgo03LTm6km3k0YkPsdF
/2nhHf0/je3VbXTPtkTiqizw2x6oWf2mA9c4hedp28El9u5rJneZSPDhpe+2
pUkSh78XDVxuxVhUnRyejqCPQY0R22vigbCZOF6uXaH9GQOv5OF7HUGhyPUS
pXLXcHV2JH+EUN/WHliuw7xO9wp40D5Ji/DE1aLFCHmITZgsidsA5rTXn3ye
ye7sIC+YDmjzaSsAt/LpP51dU7kv9EOYLvYFO4vAHAlaF5DPRPchuMRCoigW
uyfS1nijGb4No/iaUMD5Hp6YmdXY7kqxfihWWOz2msQBNYVeBTaOc37KeKPE
NnhYf+V8EUZn68ei65GpYeIpSbPS6MPWEpEl1ce0GKiHGk5HNXWlBNhbamkL
99eZJQQZgjf9CR1acd5GmKtGf8gjTXDL8WFeSMbvlZDdPiu/UT3PtQNerG/w
intOi1TQ8CCI5K2U9p8FScoSX6Q+4al7FgHktkgAJgPk9DLMU45Kh2bwTodt
FN/r3dS8DmmBxl6iH7LmVt31BMa/e+FbEk1yKmq8p+kVu82CzZm/dV53cxvI
2qO2YJZhHfvt/5OvbRkP7rz+D8HUvJ/wgJkwBWpWwV6CzpugJuRSSnD8A+EA
1j/OQQ041PNNdi7YCGFrpnIeXB4AJgnS6A01YiiEdYK1KndLLOiRa7ZMQ3pL
AsBRW/J1rsIciM3slVol7n5+xODc+Xz8Z/SxHgG3YHlreK3QdywI9fTcHVfs
DEL2/AIpOnUiHjAJob3o1D+HqNrr/x7FabdBWKrwsOHWheX0HGyHDbew5CpU
HFB/b4DGVCXRfdT5GEo/fGKDnePa0xfxsVfJ7pcLwWpEF6h2uTb4GGiPCKom
Au5W8p1/hefdA4Fpy8ssj3pP2y3K0CIN2PHI/EJsn0pS7NHG661zUVH3OkaP
WVm1fnCp0FOT0ZEbfAabMlM3x1ceITiLww16+W+b7sQehpIELbfDYN8vB/ct
59vvWMa2WRAqGcjbYeie5upVVdnDSh6fO+fBoacpqRESrInCSN2QqHmvqMje
LmMDEsQJhkB2UplC8CgsnrU0DulAhsiT28TDt154z4IZVUATQ50Lhbh071NM
kDLns0fC1maJ5SEhHt3MVif2QqGsodvLY3D1oJ+HWIkDXhQrPlh8MmlO2TcZ
39+1WCv8xyKVn706UGOTTkF1HcwMwybeM2djt0Sbq98GAGbNM+4w7FOqB0Yj
zoMuR4RLjXrL3RJPrD24q7MRyvyb6srvd+n8YS/msTuxoA9CgeAi+vmPA6or
fcX1wvbWycGnZvtgown2u8VNl5UY4ELf+jPbhn1Ux6Z6eUkNTis7gyLJ12A9
LrjHyVRfZlC+J2aBrNLJby5d5w350t6bPI51eZ4uX+0+ca+XmT2cDnRt1pna
57JsAZHcjXE/ckVEUyEabxk+jmUFMDd1M9zcJ58eMxYYEdZ7mFU2xd1I3PEi
MDksW9TenOvNpy/fzVF7qCybXtUEQdsM2dP3ONwCostqf3hfHsrr9h+FTzmW
3MC6mPjLPp1tGWSzYPvyp6oTNAmmjW82xUenNfkMdsXJH6LMBKFLBMVK6cw2
+r/l4bpakeC3FH0c1WsiJapGmKmLqOkd0TpdZz/U3ewF8PqcFjqrxk8oxbbQ
HLUip0EQWrmtWYMjJ200qZdOvxVLWj94KPXJiywghtKlPBGteXQkwDpPl7SO
+dRh10Ff2ZRl5J0Pbi+9cLn5PduNY8rw6gH4obbXMYMcMkvvGu+JEFBN49Wd
OOEc9aZmTFFdoXUpMnwE/C7gVYYh7UzcwflNBnDQVZEiHQE+3CuIGdh6LaxT
YKuJEO2vpBJSzjgSftqs10mc/O943OErwqSEspKGlyquBlSQxfu69GXqcDGq
Oji7ZdfudRfipqwXTaKwiNIPeRxr9/G3brR59XyZBkINC2sME8gcX/hDln3F
wW5rbWNiv5Gya3XwZzByCQ8a7DKUx5yngi2obAtETT45+JLNQAgoP3O/FQ3G
ceqOc8PDFqwe9DmGogtasXKuUnMS/wy2NtzIxgg8Aist5HxC5AaurjvKpnIT
0uoUTSJCFZBujSJ3b9GhFY7xdIHxfbRjAE9XLYhKgibd5f8Xx7ijYfedZvqE
y7NpYtUdqQX+BhPv3OdlMfpegvLidjWzo5sk7EmNs24RrKM4XFpx8Z26EJ0l
IFCs6rJqfMz7r4jaqV902gQc6F3KIeX6fwuVrYbbyQpiaTAWnmUMvwL9LsB2
lpE77DQRwXL87dopfbTddHa87g7I31+EOBPLdmkaZAQ6RMZcLCXNGCKfe1Fm
EqkMTQdj0An0L7HtudDWFg5d4Tszhad5HmZvAH0qPYksMGmiM/NcY+USCrHD
ZVshH3Bn0YrAB9EkddMY0Q9tOzZoKEyXTnzLMXuw1xIbqKDElRHF54W1EaDX
r4gwV4SVefC8Vlbvqa0hzZJIq7SF0yCQwcJsjQJP6rSbOaogrR70QboGRx5x
moWeGNfTD0AdBCPZZud4BeBwUDjanNSdLcR4XpwEKfAQ8A+iMBueiKTGC1IQ
wk4mykx02A12UJ5jqRMI9WYL+OL4FkiI4v5vS8iZO3c2K8Le8B8soww95PI1
jztHgEE/c9ZdX9VvBTmvy+f7JDPz39YWfnJI5qMGopGcxb91op230E91kovi
GYPv9I/7epuWOHiYm+IQC5jJsDbPmTDtvG+SM8Z045j+2BZtmRc2Lj/AI3td
XKuwuIGQ4Lm6VFP1WV3UkpZkKxkKMNvxaNexlDAavYvuta2tOiOOwuUv9bV9
Vn+Wzrl6qwbGESLGucE+qatMy3QQJqG9TnmyOAPcKMDGHhCtvwUzmLOHyQy6
5FAmC4hpRda7M7NS70OizqK/Ry3ulaJ+FkRRmDpux1434SeVyQGGzBZ3T1uS
VUnjeR6rTAKLQXMNELGYet0VgAdg6nrQGUm5dHz5Og7ddMeAfH+rZQTlUw0u
rnx9eDMQMoTZbPJ6BhsqMQv5XPWy8BW9EMf4Vn708yoV3i6CDduV/hdTqbqa
ZY6iKd6A9UXp8IsOoiSKsqufXjsmCQRY5gr3u1PTe2BOlvEAvwaZeE//D93n
RQUiHp8P4yhd26LD44s6OIzcfbvHNKGcBtg8lFuPSW4f/Fp+h2r96VtTq+5a
L53qYmQnxMG6Dc6FGL+Lx9FIbcSIbmMk5WK5gzEru9JkBBbGQRIMewAL1sb/
ogrwd89Lt14L0HPAOl4aZBj4CXJl5xD93zXl3WTUDGZZiVZZ7VSoswS5Rai4
Jlkn2xJzo5QUWYqTs7MrxRV5oHfGs89jKBFt9RTcS/P1OZ4gwWJBl39xRMKx
NvtW6f/h1YghJFNnwraa3p5rdmqklCFAawC1dnOWYVTHC3dMJ6sH71PmL8zx
llV9XXCqMRF6R9qD99YzbWEAdNVL3GcI1EFARckFbN4ZN1LoYruN40FwkEVQ
AyKs0oiAoiSv1KbD/AZ2QRlQkjJEE+z3l3e2Pi9yPng0Yh14bXdON3HEKGR5
dseBrD3IKHynjKqYDXtPCtZxMjBfqGud3OjW0l065fTqGUjoqA5W/2yOxa6v
3cLC+9HRSA3ZGbsbmJxAtLZvHpKGQ0TMxL6e5u3B6jQ0XY+J8AW3SjZ1jMl0
6zwutE+YUYvl4anZApo/F/4FnxZB/whKgA/u67ImMkdA/u1wrpKBtfaqKqGE
8e1qMWHuWtJG8CFkLI6LjBvrzR6WNen6ZOhAQUeAnpDVGhdMwYU6xFColDUi
+IOvsiOwr4ChM2UpP8oNXYjvtLq5Gji3n1W+p+CB/QNB812yCrxko1U86rwh
cpSVvnoHKKxZyAIgmtUhTf8ZV5iccLrQPnvDF/LdsVLlvo4xbyAMRc7mBiPJ
id63f1R+LW33v78p+07TdT7qdaXBQ57qbDJvRNh5wNIynjjp8XdowM1ttFWz
CvwJ6z1k9/hcfOmCXwdHZlZovZTUf9EGoWTiIc3h/NMzftbbHabV0DgrEt8H
S7ycOCBu7wcZzVlPa+3Rx14bDrqp9fTs3UFhAoYFtsCWGAAnu3G74KT163+n
mGQGAUbXC8OxEnz1V3ywShxvB6EmM6Wyav6daHnYMZEiNuSqa/GFPGEoZ2XJ
dFl1vxm1FRsRIXO1bBK4cVgpVi7ccfBwqtxhTl4HL2fXYtIVwAWI4t7I5sy6
ETzWGULEP2POQvwfmAddbndOCh5XHHCAr1QBq1iUAXl8+Rj8bNsd/s1BrdAB
+fwQB0drrn5tFezwF5mb+EJyrXG5uVmL415gKWBJ0CqWt0xnGDHTfVDxtjFK
brXH9RbDwGkQO+vHqXWjFMFAMz5FxXh2D8PtDQAbKZgTIo1+owYieamiggQF
FjpP+cZgjUULqspGx+WNeOe6+HmV6u8LCUYQBsEr0vbT9NmyOLpm4OQPt/iK
YRN+kFfPrFbcZxfBX7ykN7+WSn02x365CTe7cmBYB0ArEAv5YVq7JmI4EEWG
p8v0us9ldtnbSKRtj+ukOft7QLL6udrKHkeijiBZiXSrb59L7Lr+YrwgGBOg
nZNrFPK20oAxt08NNfPPHBcul2jrkPiqfKVn5++vMoByp6VNK/tqbMxJFEgb
Xy050d5IAaCjQ4YzGNnlgm22fE+KYwCb5li3BcdB6T6wnWo5rBdhj32hrViO
wpngVbctB8L+WLAD+o2JbujLWGbJwRMDpqOwE0CtWvf5uwLP4/2q3H1+3JbN
52p+ShZ5oo6Dp0sLCsshkXMxWglPTeMPZjR/6143ApA7IS9Kj42KgVUG8LEu
4iTnteW7t95SKMld36Er8O7tOGmeuPlo3RGsGW3VIKmjnQtJYwR++/nJeXQh
3OnRI25rF6TR3yWaYcb+v0z89+uadHp9s8tFJuwVH4VLbKFlpANqOlW26IfH
reE0jT5mc8eyC/VCpKhA4yikw/bdy6mNs7MP7YqTW5z41f0ZhNk60fCVSFYq
q3hxGD45w+0Y9MU+4/8oqaYzL7kYiX6ndPm+5KYRUINx8RpQ1uujbc3d4r1+
hF91gAo9UpUSBzMxhuhKxBf86EqK7r8mNyKMD/JuoilCdZza6j04zbpwYsZo
cpSySzlnHx4DAvHohxKTrWmRV2w6PSQ7vIRmUNSWyt2juK1vX+rap8IWjux/
Aku89WKayX1DXa7kCn+ChXERac9dfxTZuTPt+BdrNVriGpy0V6f1ZSprFtoS
qBTsYBwuAd/YEbYaBKzGRPcihE2dYK8PfCSW87SCE9x8s1otcDHhaxl98O7I
cWWFHR9DdH480MjWpFmkKwzSU4FE3DaAJ7g/uX8tCKLXPxGnmS4WEv9JmdE1
+MWlYyBj55wgNa3P06NQDHGaYVj1Mzot5PPpvOVO+Qzk7tttRngH4WeGFWHU
sVnyLzO3Dv3ehfr1kgAI0LIUhRX3Ixn/s0nnAt5g0W6mjEiuIUoQj3CR1U8c
C7CavFJvh2FGA2NpcXB+1tluQE3JO+fG86rY/OZqwQsN4mxd8yEy4Y8v5yJo
fEzslY3o+S9STjPZLDOk8n4OdQBXa1jV9X5Ow9M03TrH1GQbD4pSGDfkoqgZ
qWbrLkmpvVjXEHm32b2c7cNJ4GbBDCR6rROfyprtzf3kqLai8aatsr6XPwVy
IHqZ1106jwBAXEAeMRJvzDGtBvInig7r/uqrkLkC6bIK9Kxnv8+CjvGbW6E3
KMx3HUYzPhL8DcnuBraKA2fLgBEwiNbFXss1AcZaxPU7nIwQo7d4nIh6J0yK
N59QC5nSH6t47BRiChLd+YbpRwsfQ68v7WTDoMdosGEG1/RQsjkm5k4hRiht
ySYVjuDHsM87/ujspd1pTVb+yCQFN/ugc/fYJ6FhJXxevRJiOwaVWzovVBIb
FAWy6XX+RPQXKNdspqz8kFJpf7KRcBpps9jDBm7iBSWS+9/X2gjs/Za9A8b/
b7fkJv8GJEXETCQNhq9MUkWNBtoRvXY4CHJptGAa3upbExEpywv+OT6kSCsS
qZb7gkKPw7vVwPWiw+qabs3HiqySFbHP4H0+KscRrHl9ZD5zyPN1viUZrVZX
3GgEnaCCIEtj/C80pbVsPwTUNQPLUfsDpwEk/ns9o4CPY4H9EoA6oI9AEh4B
O1W0yIlDACKtQtdlEbVwcN2swn1cJtOLGLm26eUtILv7yGTT4wtL8w88bo3+
Vc9v6WCagjVzPg0xcM4Pf+galH3/HSiu0pnr3xW+esSe8N5OPZ7iecxspLpE
c0Ep7VF7yCmPjgy0KdBCK8I8VPBMHke3gQIoEkuZGeL+7AkdDmGLIJh2XbNO
i4hZ55xppr/V55NROaz60e5Mg+656FwSC3UR9FBMT4ZhA/F/FJ0NPCLfbk5A
R5ojHhWW2wqg94cksr7072Fb+Z1J7gK2Qv9O0x9g403OjS5pmlqWm0DYn/Tk
bzAUstP0+sfV2Wi4bYHA0+82Ri6pZFa34BHe23wF+0hKtNSArlHxqNs1XE1s
ZW4FyYtCvMH35JUyfzOCJBhTelW6kLG3zHAtBD1iWeJ4N+V4OaO0Tb8h+8qc
tuH7mLJc0Sk+jK5H233mXlOkxnq4wqcRIDB6f/QTAWUSiM6e3xThhcTRAsvw
rLm7ozPP7n8TVaWz0NwJ2hhfCjWB6pal3DyHlzmSvLXdsWabJ0JjA1yHKLGe
eEyzhUUl8eEtzetWHa21FdH0KUtdTKM4cj852anXa88uPdRQ/+7MCYIFxl9/
lc7AGIQNo3rxuhePEFZAxm/hmYcOa8QUptOf77hsQAWKrU1sxhnTWeMbM7W7
7MQtV24RUcFX+XMqYKb6D8Fu4sPDnq0I+UrT5r84HsL9Dx0Hl14p8v12uOi1
brLgF1n9XXNSi0bw6n5JmAEVzXkkzW2PSpmLvTLZXlDMyT2JS+WXjhMG7bEg
RGNKjX4qAYyibsxrNxRtY+UXSgSMe3TmR/46pfZYpGnMe9oTrPgCQp3ykJJP
ArJUAXRfd2vBBlaXujCUrp7DFdlZZUrdUsSonTgwLpKhpE8cYP618vwMteLu
PukXua6zLyt25BkkylpDuYgwma1UfTLj7vaxPWBko2Hmdegxsy4jvD145Fdi
87GOk/ZXGvz1iD3E/TWFrU9VHsUHPAlvgD0PGXqEh9vEAiK9upSio5JesokD
rSoxjYV/jP6xm8C929Ylm46EdKjUFGLuOA4ghDMKbe4JGlA3j1TjD3qGplmF
oSHs5lb1b5GFax9RC7QzMqM3eemufxxSKgotKKUumpsaKc2BXNSj+yAYCUwc
DgrOsAJnaj+NbtqGjK55Pc+1Tl68xWyawzQ0An1wkWkZaixCPjgQt3d1OvMn
KqSOfccABf1NN8ClF9JOJ3y7MJJJI8t2J8DBn0HEPtgHs+g0Iz5zTaUfgJ4i
6kEROYSQj/3vKjSYdbwSkpSZBMD/ynZ7D+NhsRLzEVCr3JYHrW5nRakF6r0/
GL1BO5NAyk+zRgxiGnsQVyeSuKwfn83qSzzSjRv9BMWkHS8qXeXqu9michL/
LSS2LIvODC7dOn25zva2rxbXws1wG7T8mu2LFXP+xE/gWwmLv+nGwmIEtWZT
HWVAy+u82inhtF3PWG/CU9LjjVh3cDD87BCmF8AZAmWzBvJL41LLNM1c7Nme
wDs0LQDlBTZx3pXSi2iIu9N2nUgj/h4ZdMZGcLguBk7UifCdGzxPwWcd8Zzs
T2KD7c2DaCglgBkM3q3DeJI8AYFVwhNTlcKFPZt2ghEhNfpSiSn4Y6QZzSpD
22lj/2heFBXe/FQXmnlP5Hd8UxkVcBREaPU/bTwsCx3Th7JNmWoJ03HiZksE
7rujZ+2MlfJJLnHu/JCH5eq3L9Sw5o+b63dbyuuD+wEKSMSvms8CVDoi9Bu8
XLGGTOp4g+aCvuOSSeuHQIUFX96A/O+CINEN2rd2urN7WLFp9s9D7hNPKu96
pIJXeqbJCbls9JEoj7IRZv/nZ+TfnNLWaGQpyavR5+joFY+/RNoY3TiodbXK
HFiqvhaX/BvAmrrxo275swa2uJzD9acnPV5uQvvOMBQKdLKOCAMeyg48TnDa
YRHfEQV4kyBK+Vad3mcywAmyUhfXU6ilUWb3l4hp0gG0Yz8IZ2GaiVXzCTbQ
WeA3tSxn6ggQ6z73nKzTCSMkJqLJPeqdyw7G4gOcGyI35JguNGg0C6K1SKnK
Oia80qoISlaNTyyH4km0uVb5BrE2uvgsGRbWPJisNkzpVr6mJlzxNT9Ye4MB
T+PkCt4ttq8gxEcevhwxq1h8iB3MWnC6lYuHaMwRKGMxgehmClBN3kIMfkLg
y+Su19fGefjjjSKywVIkF9Juua/WN2bc/5R5JjJrIXkM22atxOYIhtdcC2Ds
MiCJjBsRvZmx8XAKtXNWmaRgRh3grwB+NlSEKsWkuhM5LD2FANMKIPoz018d
zhE1mKKr/rnsv4PssglzMyUASDK72+HC0XrsWUtOxeqHqWX0V6uNCWqG7UGY
9gHlSFrCKBmPzKDjiZ/g4eU6KU9co7hQgdon+ykTgwfCjjKaq4R++1mGRx3g
tL+qHnra07ZbVZV8zugokVsr2Nj3ahdoQwex6SLjYutMeF9HpNkZjaq/lmne
hSo00OC9hJJq3guXQPhWTNYlpNpe093upxb8a1bYuSuUICVsyy/9+rCv+YhK
3TKGZsROM01dFuZ2YUS7SjuM8olta5yueEQmWZoi5X6fStegPvSKM94Rk8tq
p+cNNLYd4+5Wd0frR8YM6VA1BvzX68PY2w5h4RrmDv3+fU1KI7vFEN4nvM86
fYAIJ21e+ruxZB2LbWbsOTjD9nyXL7poR/tBjLTR23vf1AM5THuWoeXGjYRl
UF0OOos8fcZm+0KwLv95fnhq+MzNiyD+UCJYATJahVL2L4WcyW+Ted1h7KpP
mH7VNMf+m/l66ADMyI5Ko1vkiTkTUzabpNa0yaXLtM5h9Yf0Cpel0/2t//5E
zR+D3ONtNXJSrKaBr3AlvwKg8lxW2U/BXLgTG5lAzDWU6BZXOlsVmnuLzdE2
xB6o6UjL2bV5AlaqbKaePY3EZQIeKchERLaSeYVP2gr9NcDvWe1/QWxlVE4/
Nfcbbp98rQQfFa44bCYYEA5zxI6I8kdVmmbxpdjTzqWNjWpeq5D0v4jhZLf2
3qpGK4BjKRPEcFop6QnuBQVpvxrDhzbeQsqokLYWgG26s0AwRPGenzPK7hnN
+1dvteuobQU7bB1fK7Ah/XOPPLrDAR/O5mcQppCAAZ8zAukvakcn0xkbFrrp
EY4kzxIkruM7lulNforvO4wzEnuB5DbBMVtL+bfNUSUw+Y/xwiq1N2KST7FA
kXC5ph5nzZqzs9auNAygJjgOtsQefAAMUrBSLLgQtA0REbNX9FKBfiEpDsyC
2SCvBnPGv/N80Nt9Glwm5IJm4A5iLYJ1shkvGtS4TaxjbrLvNjrQD1w5/CW8
vesworRykvE1m9xKGIy9byDvfp2tdlVR/s5YsT/9gWmyClKLJtO4ELzhdEFm
6pDLwMtda33rAnMbHj9a3xHGS9H01PhV2337I3woK635fKXyuBtgS3Fjz/ay
A7kwB2C40GWhY8tMWeK9fJdiW1yf7HgpCbexnItUx/vEEEaoTyIKJki+F8PV
DykEoJrHaGOP8/AxWKyKQasPT6Vuc2rsPwFumPLyT5UanZhXIfjmLnK7C2VP
/W0fNHyvjrYRJnz11/WVNOPyt2h0A8YnQAs7W3QIVDTIBLPNmAJEQD8/5nr9
R1612uClB/ovppMtp8dif+Dvn8JGeSeLoq44YG66a7HH6Un/q/JltHpDESSr
Y8MLdCVDeMJDGTBcTsvn//XIlsDTZknaeSsSncCc3FStcjItYQbB8zfJ0566
wTpNXNOhpoQ3lpTDzCV+e8i+MDZPX930woR4jOA0YGyuGzFxTEKCT9B4VswL
r9mVWZGp/DvB6R8AUEUEjY+O4E9jV2OVQRXBEu6kdG6ByrJ5TX9VRxJUokWz
UHAo56EKZWS7fgfZDhG4uSiXWsLeA/x2ncAfaod4pOapnsNzArOU8BiKcCw0
+2Q6mdD8BRfXcwyew2DQ7pPhjQ5JguY8sf/Rt0pi5jtxyIhj2GgaO6CsxP3g
x3N7EatKNJHUzVYHQlfLGGW3qsK5XSS7MXiO2ZR1WcLlsPaRoFaLMCDPl4iX
rRPEV/i+py4NUcbjlg0y+vmxxe27ok0TiifvV1TF1zqP1mi/fVIt3Dp5sSze
0OoZEDscO0fWO/gmBXWKXrBPcyzhGTYtuv+GJ5ZsMsTbySyl99F9f2qY0OWr
As8wK0xsPiDcIvka0GFeOzxsLwyN+9j1ZE9koE48xjRE3pKuAY0YW8cpi1Xz
w6J/FOuf0zbAspu3geKMdn+/ZWaizJmZ1NjueJNE45KZPRsPuhUGQOryPAuz
bgWhkpQ9z9BmgARHZkSv2uRUkm9Ae23Ymrf6VnvSQe9cFtHSRS0q8J+62foX
iMcov5D/zDTkozYBtJKI6CbWbJueKurAdAKUHJ8L+C/ufQWjCI5tH/Ad4zsg
dW7K6GeyLbUW1E62CqTtWBRwKWuJ/DNnPg3Ngd48M0Qr6eU1MvrO1EXE8xIj
Zu9Xy0A1N2OmTjem/yj97vXU1YN5uurY5Jnr0VwGv54RkiJMSKH9TtsTvbgb
zouRiVmaZwECZUW73yKviG0qhaffqsjbCz+oDvb9xNkYEloIKpkLHrKSM4Mg
4X8t123xZ/Pq0J8FBKNjvUudvcmHRFlflCvMd2uSuqFyYFz/GuxCgRcHTogM
JuTTXpUCx33fuLW9MrssXcfHxdzL2JStIESJlDF4Hgnd4lrtHoA22k8MUNdN
6ojfkwQAZvhlVZKL4p/AcVTQ2eKfP0oL+Z8KQJO0eQ/tRnd96Mo/iXxsvuBO
Cy61ZL/j+7V8jXW3UFxpw8JKpOqpGbze56pl36tuPJmuhcIikeOAzsy36FPT
II+MiBrKs6U1xrf2OtktTHK8IVlcLryVAbrgctdUVuXNrf1GnhwFllQo8AaO
3cPK9R9NsbXTbXRH6ahVsa/1IolM4CYCvdTy36IZ5RdiiVCXMwYvXOF6ienC
VfRjqJz5kOuSmpI2sbWbN30det93QoGobKOAURdEY+5B2SwaFny+F14mVEc3
Os8Faf6Sm1TsXGfy4iT5JVwbQUlm/153nQqF9n2EbCugZtptB6LcmaJ2OceV
cK9s+Sak2qGzMxnzbcji2K06jH5D6glW5DxB/yKCdVan0W6aulbtL/uic5aa
S3HzAiyKUZLnnmbcYgGIrSFZHl8K3vJZAV+t0ifG5QyxtStRcKLhcpuiIxku
fx65v+WGy6SG0cSaupbZu8VsBr6jXYr84fooLhce/hQnWHz9W2r7QV2EWFyU
WrX/B0yqPw6Dnja5IEfk+bKgInw+EnJwqtmwJT3oSrqV4F48v9n3HsJvLXjN
vZGegQjUvCayt/toHnXjYZ5sjURUWRNPudSsiD7wKJZWzUuREjt6rLi7vpf9
KiWcM1xlXd9+dgw4w7hG7IEK9gaTYz5KyX1gajRXwzQjQhHOSrAi+yOaaGtj
AFhOqyskRMp+JDVViAC+IkZ1+yooNF0nnjZ3z+WFu0PKMnzyeCF6iaKsjkte
EOOK7qGDgZ9oqO8VenDMuc75bkj+teiOUtYKlS4aFi7tezo2tfNA4f1bW6VI
adVISatJC2SZQvU7wkDCEJ5vIDIPCNGHrMSPComBbxI6QaHiNzHp7N3DIcTr
e4aeNOO8g/Z3qhmWcsl3XMb8tE9BfbPb6L9xc5fJxhGkysfdVs1Ivp8T7X/X
Q50f45aOaBaypjtfQbeZwv8gbfmnJmcATj/9S0qmgq3pqc5mNhBeXOenTfkX
re4XQvwujfGIYDYzwQfMu5z9yQXPC7WxElzaUITa0zIoj80E7CfjrMS9H6cP
iHanbLYoLqMdfJR4mCuv6Oij4gMExNlRht/aprzNdU5q37Ciyr6Kck1DoIw0
E/OICdB/plxvDyEtwyt7Zvog/VMDFcn9/0jM4v2/5BdJuWhaybLUhz/+ifz5
zbNah1GvcQG+6K9j7W85Y4TaaTUBMNuCozPUU2PmVufFf3T0I88/vu57Hod6
w0KgbFQYIsP06/xtbyJzGPYTDtYa7XpktEO8yWEnP1GxaFAWYmoQDHSIs1IX
pQKflurxEZN5LfHXF2k8B5b14CoJpciPc3fpy1mTLRvs+kNn42S+slO1DzsJ
mePV8lOvUK6i1Qp6BLRyYvjFBltSQKmotaAV3+HLbhhgRa+colvLio6C5K4u
9M3EXKZt5h9aj/PtEVMVVMcrCxz3+JTm9aUIKa3h67ZycDe0/k13n/sa6fue
XIJPD9zBMnOdnEgwA3tkzp/S3CXctbzZcZRJLV9DJKkSnoJxS3hrNOaLit0X
hu5T4e3gN/MTvi4VbYyQYW6h1gqqxtou9dPjufxPZTP4qktY+BbQKcclWcLt
mrd/XyvBTnHoEra3LV3UrcbVhwu34S40+uSd/m21w7kKb5n99Pa+E0w6f6EY
B6xqQw2llgDtkH/HEmDOEG2mR5dKX1X5c2mNOsb4+zu+ujzH/HVicvOlyoT5
ypHzESZS0zJ+l/+axuhT0kb5YoUiU7128VSImYfrYwWjNQ0C7XYQBoUvGzRo
Jk/k1Yv14wa6drh791VQGthX12RazOcmGvYrKydip8/2S/9cvReAuC2nHBCW
3aGwrxMG7bgmyN8q2Cv46EDytcqAqd4j2RpeQJYdEL1hNuS+lWNVN+4L3l8o
NDOwUwqeVcf79PbUsivC1k0qCfsyy52u0Nt+/dTtmKiEYL7qP1Lv8jYmPleY
u1HtdUXNFGG8HatAwNCh7+Vq+/NEUqi+CPduYb0ZS22rNRXiuj7t88dGXZiI
1pI/Xoj1h4Xwlgx+GBbfflfSZ13HZ0TLFuunrwLNZ8L4qrKTpRQ4Vt2UCVzn
BOIpEw5x2XzhPeacIqwsmRJ0fJOh2frpgvSaQfaf7EpTpPElL3oJwKtj5IwL
EZzslO6eUHwo8T9L/99TwoSOMwFsRdlSe8B0P3ih7jnjO9Xwr/lWg3mKqRkZ
fcqlqaDUz7nMk5FcbX+6U1qxXOOQUnFhfkLS3FxZ9iekQl6XdxEkEVWkrpKh
ziC4tFc+RFcl6SXs8J3YpKYV9LLdkXVXQYQ+34DiQEtp3bga2uwd6jcwr9lf
D2YqU/z95lszRKwnVEHQCR8lOj19po1SRzERcgs0XcjWN5MaObagV3ONZMiy
r9fDLgEvx7tL6Ia5KM4yUSI0/6rxe3Ibj5UaKlR8A8uK/CwMJ8kvqY4hR2lb
HTxLO3952tD+l4vDRRH+/7Y8a4atwOse0vwVUxieUhwXc8xd0gn0CI7Am/cg
Fd7xSfz3zmaRm0I/djbfedffXxX4BQrqVWaWR5uy8ctSmiGl6NHRJcc30JGQ
tA+tsSPvNYB6qGMajcTPBQLmb7TK9oqi8yO1nPvRv8mZ4B6OpvuXp7EvNyjh
DKT4LM97GqXqGaYj0AjAW/2L8C/cpIRRFoBcHboryre5ZVBM6Aa20FFsFx2U
XzvUwq4JjDqCQa+NSixREz0k0+4BJwba+MNHVaTWWfDcA/zYrWm0C8yjBC02
HNJaIFCn5wlW1eFZ0SzRvmdSewKMMoWPmaZK6jttVFRaWPrd8Xw21XbDcBpx
+QrfhGRoRmFUoXj++UZOdZ7//uNryayTiG4pHYcU61YJXsW6QdNKq5cv//WZ
TlGiFYVrIxi1RFn/qe4deR9jvCr7sFAVYC5Xgzh9FESukKqptGkkt2GfnuGn
htZe6Lxy0t/H7A0WSOMws2a/UzMGC8/FWDGI0j5WdQiCUWdLSVBVNrfc4Tdr
TTg/sld+riO4MCB196ADp8Mm9QmnZfYxIz1/SeHgL4+c+k2BPK/Y9+uhj92+
311YeMjLyf1X2QQFBsmpn/BgxzAls68N1PnpwqsYtEtYZCnHPPBeNE6Ria7b
BLO/vaEJ1DzLQ5RovNkPiWuCYKxegUagYfhlXGsegNjvrbcCAnWDKKZT46do
+JQFcmVF0Mf+vals73V1Jy3u4QhzO4vBt8Il8oHiU0fcUAL5I7neFSljP13y
2t33fk9U6mH++9+L+18TBhau30Tw4dv9Jw3r6INpsGt6ZSubLzp1RTnRvDto
MIpae15XNu57rUHlJJrMlPnswd5jRo1ExUepZWRWk7e/Y+fWkI+NWZbG7cV7
U4CzxC2wRUxW3c8nuED7RcREsHhHHX6WHRxKaf9rPQtHu92E9gtWAO5zBIMH
AkYpxnzbLQLPAF4nSIBJIfKAYgp+xmESR2kCnpRk4bBPPbGvVzmGmu9ZukOr
Kqn+1AJXrm2vm9QdPOhi2wV508HsKAc6UXDLoWL3IEEmuC76hoqouxP0rn9S
80m4+wPu+FECZI4g6wbyruEt9RvrTjLUffqaaV/2aBFHsuuoJKQYiPrtpJBY
cR9L7T1iVS9lCKcqN2Dwnjv1vPHjtQdlh2J3Uuo6tajZhVHdH2Ggjwe3QUhe
SR6PxjcwNpvKB+pKcPX6em6ZC1eNJloNsUgVWgKreFQ3wkbs3y/Qm1iO4sE/
j+uyc4HWyvuSUpcxEbmVDm8NlD4G8B1N+H5Bt8o68+C9JzfKXsx3LcFONMqb
ZROO0bi8XAU7UvigC9bI7h6UEwXCBUhC0AjtOVHGmMgTVBhwsf6UG3gCsx6Y
x4RABNKDibxMatB30VwjlaUnkKN3BUDAc2ovh7OP9HiXDbRzAiICNSVa5A1L
dkuSJQvBJmhoYe8LrtgKR5HikGB0aFY5aZTbJIGKzS/3Uoy9FkCu2St1+qDw
uOxKqEg9oZG3XFUatzPRU082jGdVnDvfftxFIpI4+VBqIhmvvs1kGXoHARsH
2lIEgSpEPSzk3VSNoTT6yX0DjYexd4Pr9jUJGPnQm5mK1Acofon29C+yg7S1
mFqnDbXzXMF68Eq6UIWsWvTnzpZ6S/nnAm72wA5wh4vVDXgavLsJtmdufKFF
25u0gFipyoUujiuP0xwdv29szun+SWp4EdUejP4207e+4drvqox6QIZ1OkuN
K53a+gicpe0/UbVB9mCF1JGGdwaqGbX5moVa7t57xlLtj0Oc4Pykj5F9BGP2
qm9s9acur0LQABmEgGLcJQQyJWCeaN5V8ZxWslwBXZbqRKlDe2s/2jIpaWXK
xteH1rCQDrzh1hu4Eg8M6uSAk/ud2mq3SYlxQf7D5W5BdFJy5TD9MaiBeU0w
XcGFa5kq9CS+bO2w0+6tU9fe8wC1ha7KIyeO6gYXE3ihkKh33Fw7Ubtkn2Bb
hrTYiqW/7zHKK56IR3LbFGAdzA8yG0pc4gBR1XKlQLP69uYMKVPiUAGjz727
zgXCiudLbqCiK6qn+10jRuyYNM3dEnLUzCD+g41d15u6ZrBh286osfQ/Uob2
vKktDrfxpP+up1vQcRJ40V8gafBvNkDRcJn1YP1ZaWokoBwf0uuvTw+OoWdW
aNe2qv5zhxM4g+ML5MBAe3bSTaZVIRLhtir6HGm/GdTJB+qgIInOrONOPzGD
wUSxFeQ0P4VSXWl6IMKjCbWybuWx3KA/dg+E8oDXBTgoHowXxSvE2T70S/1x
fAu1nl87kU40Id6QtVrl9VvZPU06oQqxrSX1uYNRXPGZdo56n3g7mDRnwt/G
T2eLilq5TfOwBVDjzoi7oJ9EaKLhzahJukiekZQrO1Rjb0mxEofy47lonBa+
XsX+yLn5cTp6Co4eQrlACcsekgW3TaB1BOFq7XO2Ny6w2O9mmlPq1o6/mZPU
d2DlCA47drgZJhKBSdH7sgP9Byk50xM6LSjp4xShDkEy6L5rkcjWBlShzEFA
Yn2o3HxdAy4vfUIuTDcZwQBa506TCBYZ/eMMkjIgVR7bnMu8fgUKiOUh5LLa
o96gks9+biYfy6FrS4YoW7hsFuXWogzs9rByn9sT7+xINfOUheOvHvbsbSK0
Te+CLf2bN4JMxCzX6FiZLVvdp8MEZejRKue/lO54el9n2lahO8SFY4koxXAT
dRyjvFMGNov+cqzC6AvVcSVyRqNILUJDUj85Rx1+M79+aVNj8jrc8umsHytg
K6EsUMiWRiFnqd161fle2UbccJp0Cw5B5Phf3va+q+pc65T10+jjdbLlgukC
A9MHqb6LurvmLWFw/6x9cGZ//QM7ivhW6qyhM4QM0rJPJMRF8T8N1pNc0eMm
eZhMx+XqQDIkP/zbYkib+TdmV0JcetRnsXgUR8/Si1fFdz+8/1V6u7duZb7Y
14IOJUp7U1ikbRoeQSsPUZzDHqksWgucBLyfGx/QTH8979aurRiednqfwFc+
rQ7W4+V5397N/ywGHhfQd9u7rw8JX8E/wPw6QN/gha27Lc4wCL6+TcXJktjV
oe1R1/wS6yoMIMx2SF8rIh1BS46+bxvupzZq9jI/TGxPKKcuapzW8twyhNKE
frp/gxuoasuC3nuKW6ucc2WAqYFs1iihdD/F7xFG4bvCuROO+Pi1vlgBo2xb
fuwv2qKboSqsv0A+bxumuMpu6TWWn5rW4Ox6qeUw0AxvOUdPwdTG4AI7O3yS
W+qp71c9DggWhXXUWRmPHKzFTocMHUSXSe+pdEqRbb1sQBJhHRZfJEQf9Hja
pMHNy7qP3A0PGtwQWLWKYegsYuoa0fAYElFCMh/gWwem9hXfjMdf4M8csRyq
6Bst1B42ma8x2Cd32kyjf57w0F66gzDYchIz8ByLuiea2T/kDuvD8/wtYuXT
+ue0fkmKrXpVu8mmIKb/09AaN+KuBsiU48u3wrDt8ekr+zPmCOOisn8HiJ1J
VbGCvUrBl2Q19g4MR061MwKOUm4sITmhyrj0Ev+tQRDn+WhJWMsTC5Wx6ahS
F9eAqzQkLapOr7EbMsIaJ9Cx8gYsTL6ts8HD3Wyb8qifGOpyPV0kgGChaclP
sv4rznsJGfazyVcKOpmru2VyHx1nOZLOBHNZgZk4D3LyUD9E6aJI5Z00GHnU
ybcafjo55DFsDOGGbdkgeZtm5qZC9I+2GMm6GC7u1Zzfdst5tO1xEWpzcJfb
7PJCD2ivrnVo0TDbpaos4mX1UrTwSNjJYFix4ZcOTa/OtSoChBO18kKMmZZ6
uNar/Vu03nDc0hl1XhXIG2L1zo0cp0grKaID3cNc7VwX+lNj0GQcOqp45wlL
HJfZfYWlrGfmRncxItAPfLl2wPR1sn7bXEc2dCVhnJhWwYHS0oyuIAUqY3mI
JueoWM3G5fJ5DHvIcjDA3jLEYFhF3MTfRUtvkRkk4cFrUq2BlJC9Pwr+K+0N
rcqppMJw+ax+vmp2D20aByjZ/pFBEwanozzvA4fCtn20P/skqLQBga5ajeXf
9vMMvORGW1vpondaMZUt9ndyzKNJUItED0UaWGwb7ooMKfDVXHCzwnkP5pXx
fqzhQC22Y9YuOy7iFHP859oo0PIKzclRDiVIo8JSBY52pE6Ys6YtGxi6WMh4
aACH8BL3x3+A1EYUdhSTKfYO8ChTSmRyxjoGuvfssYEXLKYLRz4iv0dDG3dx
dW0GwsXmX440Bk74jFx5UZ0stZqoXrFw1I4LPYuMDJgDs9D7e3LmJhnc9AEu
q77I2Oi6DQleCiY1aUjiRkahhG9v3/KllLP725dhR66fmgOKmqYVbXRi/P7d
+JPyjeYXV1anKvU6n06vPASBPPFQGYQgFUJxy5f+OHboIldxb1BpFWhd69Jq
OvQik9JyEeQ2hyzuE44x59wrkjP7gy+9NYfBtIPdp+KRibmRX8B7OaRzITnM
9E6ylfaJY90Ufv35FdyNSVjD5kRIATESvC8ggVz+Vshyxb8lq0WvyjKMyQ6o
9sG2Tm88rzXsaBF3msSBvU7o0dXmlC+kX1pQeNXugHeWHYo2+W5czSz6VHn2
fH+tUemqQjVXwt12V6+/jgtoQlQNJ4synlbc4jfBg2v+3HCuiriBrmksoSgx
TGJ5FiHGXuLAOZhuW47RRblp0wvg29wStJehb6tGGIJy7KTN7v9O2FpdbomU
0HxS8HdKYZCXSMnqDKgzEu+LRbwOwxoFlymib2tFcJcFaV2ok24uCdEI6y6y
icFtjaysjg8QWJI1lucloRSH6Mdd5UdRPzOK+ND+PMpAmaveHF2+ww/UA+u0
lHVCDCgMYqjTEhqgOXub8lTSOq9G0AnqUl3LeY6LV2otKDicf3VEHXo0INbU
U1L8kN//8W0JE/tgr2MFDnIxENMW/Ry/S+H8da4L25jhhdQW/JPi455T4OHp
/zAzOXTV1+Q6xhSHO1VzrvshOCtnEu2UhVNNPAFyw+nW+LpJW+yb3CZ4ZWxG
P/KMV1Hv//tp4cojy4ClvlbpGNAluHcLXe1pznzaOxF1khpKi0lQB9E/15fS
9bwCpR3LOrJNJ3qPDo7z1b42kQh5s8eBp12PWBZGc4aGK/DEA9EI/yw6dV8o
jYSRfXxSLp/GuFwIfwN87t5uv46J/yjstqsg8DUQ7ZjNatO5OEXhClwiH2Lw
AEx0HFOb9ebKzV6qjs2UrE99MQ6WdWu9kpQvzz3AVgwOLWaaI9YEi3mD9NQ3
P3ACsb5A0HuNtA85b6zqUb1xRI+8cSum4vf0gj4jQzUMOxX9HoHrM8SWjZuR
8KZAF7lLe/OuBl/Zaz4G6Iq93hjh+VHUmjmgn2ZDCI2eGZWSZBTAMC848B35
mbzO+JBqnUkpcb+GKlCOsLWT/QBmOY5hifSD4yIBjKfFZTM1OydPSEkTFLXP
Ie8F0nKOlYNpukRpLW2LkU/jWxV2iwaWhVMpkZqhqBNqB6tA2N07CT/oAugx
GRgdyaJjWr6R9BH7Ras+yfjyUdMEAJQ6OArbqYtj/TVVqAy2D8HNsAX30w/e
BPBgBJxafPkpgoMbLM4SyWP22DPxbsYgiCKbBf/5o9PJ/C/Gnl4zhJcpf8m4
/+JfIIxgZYrKFYeNX3py1YHo3log3A4illrH7+C/W314yJLUOm4Tl2hgLCBQ
xtH5QT2TVi0DECDoBoVLOUoZtENsq6QsUyVyHjPOcov7gW+qbRmPLUehJypU
kjKVd5Xr6xCX61efTojEeWRoWzc0mAT8LXL/3D5TFHahGAstpININVTwnCKC
v7wjU2soXTon1Ww3WBkz46p+FVu8EFd3iJsWjzHrmeDpg85vxFOtgGR3l2ah
eZe9Qh6zZLkIYT7PsfkcLHBj2QDciqM2eH/hHznfrbQh9oEqF7QR16ras6OS
QdLJQfzTDd3FmgH8vCwYg44hmFAWiSJ9U5bRIWnpXtBfbORHP0C9z6tmfH8w
GZ5DhkNSabLiuUBwSL5ALQDpN5hg//PAGKaAhv1c4tzRcFFMNy3JWoeAaPky
KapFDTLb5tVyhDKFxDQ0SHP+0TXnlDLxtLLDST+aYOfjzsXKQBYWUaTRQQpT
Ag/OwTgjbSM+aVEyAhkxJKmdl35QpcSYl3HZzou6fFS0TrjQg4/oBWIy8zk2
XFSMvI7s4iCt83V6VWNHSdll+H6p446+SR2jivZJMp7NrSALBWP96skR7yK8
bml2/WwUmicZNDhtRgUautB7y8ChG+d0R66VoAdigHRXMPxjhrGYxaSIgNBr
ZReCGI++ysRfOnKBYwY/c1D9fgQwyB/i0ZHBisZWnNgBwNum6/W6vNi71o/m
C69zrm0rP5bRabUx5zNKuJ9Zm6jQst4FlpnY0Hy/6GRDPqFvTl70VwqkW4sr
2TFQ3vlPie5wDCb1f+NJ9zXRKtDEkvuIy6ju40annisZJskUdAFrTDHALRbV
4LmfnRw860ebWemMSe2QvbRq3+Zeer0o5exsmbZlJembm89GoEObg9VSWLal
Tc2b0I4SvWRm+OFL0Iirn9qK6Ej7fCiXpLNa3Mhb6Bpb89/NY2d4n9tawvza
YZsgZ+HBYi4nSqQYV1SVf1CjXe/H/hk44UjE657mSToXzg65nJNyHlLC0j8q
EiwhuFD4rVCqAB/XMfc7u7GwmrmoWbki/nEzyDMEcNLXVw+4x8u1j2aBWhEz
Z/IFmH6hPOyS9FPhU6fSr1TtRXHHwEmJt9KOxEsK3Tu0duEtcayv/MxK+ymL
Rm2MZNBpM2EH5qY/ylMB8AqQdKn5/9SOr4Jf1BL84EqMtDbykPbv/jt9unMf
HHGrV9yJ/QHDKejgtJs1O+q7bnREF86cmvRzYyMFBooeBkQhQ+dXvO2os/55
Q1h8x8O35P0pZDcd/dCyRIIFn7q+XPB60sMsf5lPxK2+ArzV7hcaEZC6V2CJ
eXGPqqRPeUaqQDygZF6fgZdneNlfdeq/oJ+RcPYx9/s+euspIv7Q1QglUf4J
Y/QNSp8+xTcJPXe/ZQ1Gssy/HsbXCPXGB0one1CmBalk7+lLX6rBN2QLLtIU
ZuXA/sYMwCJjIKA2Gr/51VASHaab1i+4DdoIxMuu9xKi4COSjArlB7u2gsVK
ZnxmrsVGPH74U+E4SEzLCnO+QUXi1YkEdFqxAW2vK1Mof/nO5gG5q1jAtjnq
LJIcwljjAl78ZVA/MpmM4wIdxbrA2ITvli46rZ21gzZxvEADhDx5vZEa5ZHC
FulVpLlNfa4gR7PClJbSInU/Du5xS/wD5me8h5Ht0bo3cigFxq3udJoxtTRm
nnzHCBpEMSnLAgnfIFwZeIh8t8VzGnGkg3SvUWI2EGH0hrGq+QyP83h7K19d
aCgwv0pWx+pWugyFKe7hOHMQBVeWcGZOUCWdkH3wR1/crEgq+mUVXz4kt9NJ
W1FY1FYEQaN3W4LyTFV508uFg3GTt5vc1ZOB8SoFlG8m7WDazd1/zHm2Jtk6
tpupOJ9s9xYAsUonNU5TuCFh7sdvrrMXunFqb8l2+ww9g0AuN0B4ne+qXppD
S/W3gQ0AYN3VCGwcDxpsVSIFNE6h7XRTFc2hOUmZiq7xmRiO23cMlXtyOOey
CiZ8dIVW+wEplVJm7nXsU42O2EgMTBQqBSTcMzAQHNCc77Jxv89XshuQtxlp
xSJjvSebrMUBNkfcLTT5qS4KppBVFMHAQVueglleleJEk3dWWEsv8rLbUIl6
kOfYYNsH5SHYuSZ0x1Rjqe6cNExlQQ9o0Q2QsieGDnLWnB7ppoSYM7Yi6+M9
sF/QYDnawXLyHkGxh8nFtHQHmyT2sFrX/X07Ztb7jkJ04DhOrbchVkqtFQ0A
DestCwapl/I8S9H6ZiNDg6b4QaGfyN3jmeN/zM05nwmx9GT+BYc1Xa2317Us
8n36M3vXaoxBSoK7wSYQQ3wecKuA64EaHBAa1benSu8lWPAcdjc48C2oTm/j
bkDxdxGaryEZMP6jgNh7RI94kYRRIzP6FZrqOrQnWpXVbUd5KFfkYwol9unA
rUa/KaDk1aRGEsYmIPFNRWuF/mQrdDSYSdU2nbztcVcpl9u06FYxUU8tHJqA
S9oxNzeLNVp4mSmrPIuE540aV0yU4AAraRmvnIoyyFvq9vmzjTrC2toODo6C
sXoKFc2jVRmEQGrjSUxs3Fs99TBLbSaTAiXwpLvL8hgEiuyZdd1h1qTST54R
zv9FLoacZ1dU4jN2XwE4ICGmqIZhKer6OFGzWmrmguVMCOSKJFKijwQJx15e
VCmjS7pp0M8/n0+XaV9d/x+ihAfTjN9y3UNPWE8xPhg/zojkhYqhMU9o3mES
nIV0m+YcYUxEcL4zDBWLGn6XgRMx1OlMNuciysN31Mu38N2PJu+lAJ5oSrOS
s4hj0lFRFVnkIzRm5g/iwqf+OeV8ChXOaasmZJZ7wf6qEzhyTVbQMJZOsLpO
5VlRuwJCCpu3d/w6NeSjBf9fMr5SVTqYNSjjCY+/X2WZM0a9cGl5lHIMuslW
u87RPYLdSTkVNVZV4djr0YiYWIdxpThFi1Rww1VlPQB4g7OecIIcqfSFENNu
pQUbOJPtOHeY0ZPz1GjbZPKYmsHpPK/AxPkV+MYEgNI2vQ5pWK+UL1P3R6x7
nGqYjam2UGe9vB+sq00x1jlVxvgbh1SiRlLuJeJ4/IRT5U07Rk9NUEFG8+pC
kvQ7jAMq+sRMIw3h3nuK/xTZJt+/mABIa+iEaHexVlsGA9NQJRpx7GQ+7f53
LhVK2m9CqFzsRs9GTp//HSXDToLcTnqxGFi+Sv6asCWjGZU4P9bzWNIaHNH9
B4NRlIOKEMtOXaOsMhgaslqL36jCVU8g620bcP4jYHR1ZohA0bNjSWm8JvBI
2usxUmMaVsMxa8RVgWC0hwIh7Hmqj0MiE0O/Oza1ZOiIb+nTO2pa95+P+iVx
7HzHN4VQHbDL9o4x87IjTu+yePT/+P/d0PsoFmQuIvPexWfo0766jW820Ubh
vrGCwyXYHGfbCiMf+q4El/qfarsrl/oj+gsGUu2DH1NTHMwLr/6JE8O7FafW
mBsKv/QPCzbNs3DQEkEOgYRp9jMiTch3/MP8yI4ioGNYHF02P+At6c3jvevQ
vfeZOs1VRfbMAv5tcS7tXMuBRxAkJWXxSU8oK9v6T9pmx1GopOL8XFY0D/bj
3sTXFiAznItuwwI3M1MhFaCmxKyFBW5Ojo/v3+nb7+C93ivVOWjN9aPO7XFe
Dql/Fx2AVRqd4SSuURK8K6f1qhx8eYHK1iKgbRnq7aj7lNwoc+xzk4FXLk68
0OjBuKvx5sTUeYZGyVoaDax5qF7Pv5UWZ1S8HI0iva2ziXgMOqLqqvYj0+Sj
lsn6u9M7/hsuDjjv+amERYhquaJBy8YPfH7IRgALqolk+2Rrt7KWhH1lVCZ+
RmBqtg1MaySgn7/Us8da0k6HRMNkl2suMe3d+fe0GvV88PRLbSM+jCm1cHRL
wnzzK4Vayszdwa3oCcE6T5SDGno0ihi6SSwbUMk3JK30VzFOeKhIusdCmXyn
1IpPA6fQ4Uurx5HpX/a2JDcYvi8VYg0riXwQivvICmSktj+rq2gZYERRE3td
SPLHfqhJE01GmmqWjmCErpjattYSjnCinapjW+/aEGm9c55V3IWWCuwWCY7J
HVWV9JV/4xcnNSxeDT00cFRUg7ew+MAUU5JszDpdN2L71pFEktlaY6vwRfkO
EQIfp8s73FVPrYeKBQv9ewcqPf24Yef/3H5O2VhkQakAfCCPyH8QNgcHhTAa
PW329PxxIUdr+PSLygcCXPRfjzhqXYypXqP5KoYIpb0x9roCRsNo5bhRKYiA
2uOWS8MtTo7VtLOmwjlrxTRNFNv+NkzPbsiEuWWQsxfV3ZlAmm/P0chSfNs5
wydRLxc6wc6SA4RwAACNWHaQ6lWU3u5Pygu2aFcfDysaqDHdzWSQ0j099P6+
Wd79aXaboIegcynTGucngCAj2ZgRriyNZFQqeJlBlPGw3yDWGWCAqEVy0ZIm
ImXiucWo5aseCV0uGM3sKx7Afj+X/TxUvAhKxQs3SfbincCzA4pDcvSlFtiG
zqQcP9GQzwQV6LwPSJe64oTadF4gsyL+N2qgSwLKSLfG+U3fze5/JytsT5Y0
HXyHajHofO0dmRYt/yAE8XARu4ADDO/e7tK9qS25CMez3ZwTxLbQXXx/Tu+I
1GcUB2SvdDiWkEUqf0YJtRA0erb4TnqYKAUE4mElEhpGMRp4iZ/1z8oWjd7c
uZesyNFz3OWIDBGjtjQYx2qWXvDSjUnCNCOlo9GPn7eiLOP+ZIrzKIK7JNiF
ce0+TMx6RxQHAJhsJ/dFwuINN/RmQqi9N9peqemkHuhpe12VS7Prm32ZUv9m
wHc2BfWwjx+X48XBe5yA96T+9PyRVu7lZRH/i9w5K4M+rintwfeib0XK/POU
THFgEU3lzjpkLrVtZOREyz3PDWy7id90fpsjVAs6tmxzgYWgZe9zS7gyxTYK
rv1smw27zcZuU4yhWQ5JkVdmN0whczzm9+rBnp15oICyVozQjYajEwckmLu2
0mrpzwdm7S1jTskcFzfYzRtNapL2wugRKPvuzHUarki4NVUgrseQ590PXdER
dBw1sweA5pN1EFNIjxMoqF9eDIiqj12w6WrPmQeQ0aqVb9WPtuwD/9OYIRZO
upQRNNxI6wwDOtHJ22A3copm4qMLN5FqFLSraGxMVXrU/aJu4NhXdpJx35K6
cHFgDzbTlX4xyWOO8KZH2ZWTMyGOqusTCkfyLpF1/FMlpZx+8DhYTnosYRzC
LY0pOIknSNJoabC+6oak5uO7YbrK8modS9cNoNTyPz7kTzaWbIHIjwLg4EJl
s5iz/Ag+ipv21tReyCSQ4FlZ3AcOZsOu30s+mtzCDxRc8+w/5bQX1JZ4KxSv
v1sIUEFLfLnn6cEg3/RB4IOTj9pKelU7v4IKB6doRzCGa22qKVcEyaM8cqNE
UZGcE0U0Nkkk0ThDDCK4fXZLBcyt1WkR7eNVj8HnCbsYmeyKz4p6DyZ7hnc6
fXv3vPxrJ+6yW7FIpRtNfXOlZD/jM4m4XBN4AEWmf0bUpynhpqNeutHkpDsF
YcOTWhfXh36AGpgCKyBC8onT5d6N1TCnYOLw4p/aeG6LbWX9TV5eBWpnQ/qI
yx0jdkngJGWm5TlWuhCDFW8wqa5Dsp5Rckp2WENFxB0bykQITYjUrlaEZ7Kg
2JaRW/1/y2PM74hFan/E0ZDXFz4Y6Ozbk8d+JMMmVSDWXJzn5GbxGVYUKObT
NWDpcIGOplMJ7nNIdF+gyUDNUqCVlPBq1TosyP1KS5RieSvDAwdIR9Syk7Ak
eD6C+AE/Yg2CZV1s4Z8TuHQLzZ1WoY3MGaVs+CIIMl6yyk3nCwU5Cf42LpEf
IJ3K79RC73qi4pmjm0Ahx5NKnnBJuSLZDF+j+FoHO6tdV/F4eIrb3qYdUsx2
JVjbqx2mpZ6S77T2AN0VeK2v3trPt2gAyf7T7nlTXYGhXTpTlxs2rECxE297
BQcB4x/yvCZfSR9S7upFhvkYEmUGVZQpzOgIreteTMRRseUP5MUu+Mjuzm/c
i9bAbmqTvOLr/AhXbHPXjkyV+Fr6Edu4jCOzdiGnnBWJPqWpdIQbhFYlbaKV
J4gYiSvVDkrb4qo8xWAOhuv+8CHdmpeFO7495EjmcIXmwfC2a72Lw0F51VYZ
cYyRrxEbn00bEe22mFtNqBYW92NdJk2iXJxQDkgadCQQSGvFO9nwz1aXoetf
+JXm/ge55R2RpukSXGP0QvacUDW7ibtC5Z4Ele24h6GlWdKnKWYAV94q3OiP
mN3XxI4yJN/rOqGpTbKIusd5S1426+Ck3hsjaEcZcKXMPCSkyuB3QSzuPsXt
QslUwVG+DruE9DRVNFAtt5EfSOqk53/w2/abJkL/M5dUU09hYHK2CjfIOuiO
SJRFhpFEdUQliEdTdWYWEDnNrw7IClvX0/YDsthQDOpRcVSUeYlcOliiztNu
wnXKo3PAhJwoV7LEAdWLTg7pNg60nf94XjDuuvEIep0fGJzteJDsbqT5/26N
i+H19237qafYWnfSyhitMEQ9y85eFiW9Mf+VsqtYKbb+QtDQ5X/4ZKs04d4R
u/2wdJfEp3J/2wiPEguI+qqdEJB6gkDHZC+EhPOmhMVvGyGTbG9EZJQlkF5T
eaMpYBRuEVcs729ojf5r56j2/I9ezFMM+Q2uJm05aGHdjehJTNFROCHeydFv
FhESJWXYtPY5Z68nFQ07chpQUyzdAG2HK1fWAKo5jmy/RGYiG0kAtPFKLtLB
Y85M5m61Hv7L5b8Ny2YfMoihBQDQv8y0LzWFM28+E5SbQHHF2XOdO/6ht5PU
ZRaL2fcqsgUjH1SsEvv/IG5t5jhOlddrfBWarbAlUJqDO1FK8bPWLCkjum0l
VAMdK8OYjBK8bJxTPH2kxdc1RhvSL70pbEaq+AhOumTRmeIvupv5tgrZH6s8
ZXUjeTg7brJOo6wJERZAsVWfKm3Mv5z0AkbttN8LWCw4D66EUSolEmBtpj3c
qHNQYN/2YqbY7E46Pg2lOmf8hEE26mf9YtuNyO7tJTh9QJoaV+9a1HPrnw/X
FPiPf+RtBr6SW8CdUnuiSzvOYLqa0+CA9vx0/sveE1ssHEG/N186aIO7YOpC
4dyIzIorAuGymnGFIKufXpSTnW/ExMWBQ43VtooqR6606DPsT1SS/Sn9nahH
iwhGGCjvWISs8iO5yDecWjquagVMbgo77DS5Ab1Cz5Y+b0A5UenPGGf4Wg6O
ktV7e/LqAHbbkS/Ct35a7Qpppz6qks0U+ziGqsRyC9TDM6YU2AqP7JYfiGSz
bLMdoLH3Tgo5wEbnSGxP+jGfkTEXz7JnYbIdnPgUhQoNKwmb2LpRreCaCbCs
kzoWbhXortl6GvbQ4jlXRnk6n0caEpoHje/bRBbFm1wxPcYAjya0XxMd4kk8
YNw12cl/8INGFDFXWGgzAJdwoH27Gk1S0i5edqrfQSvWY+O8umnZSAeILZka
4fDD/hU/Z5+wqN2smnBYbDnd9RTT9VGQNcLH1WeWIPq0jUQjDmVMQ5FriqZ7
o6EdvnqFTdZGWPbJjijYxQplkkP691MOJVm0Ir6UZGVMyyYHaZW6AVM1WdzE
v24VRE3IHDnKQ6Kq5p0f87e7zD15M0pEibVs6tXeFKrqE8MNcDZl7OUxSSik
nHLARgw/cYJ0BVPXBgFfBL1LkjvS3R0idxV0zP78yILgJHyRorNhwgHqoQ9q
/Y/uLiM/RARN8d3+qPI499Gs4dh5b4gnYVS9Z5/wn2lQk8ZzBJLlxOIrDJ1J
z6vWAR/aXpjnXQZF9iMet02YnuqQ0UqUVBjowwKqup9UECyxFlRzXGRoJoi1
ydlFdZbldpt5ux6Bd7mTEF1+c/utMtUjnqmfQM1i1AbfajGcvOSt+XrEOfIx
Wroch9TydJzpjRBVHOqEIRxr5DI6XKpVct8uf8nvEwvrja0dUlOwAyzq3WC2
05JdXnEh1pQpYzecwSUzNoDHcE/FEA2ICxmC/CYNHfL+XlOk04hdAkNjivFG
RmEXjPWjyc4jBIORZy3T0WJp/s1l1T5RLmVGAGXCVoSLoTGWeQRD3lQZLHLC
29yupNp+Wq9zrt/BaDQWIseBzgYT7IMlpdgFEM7/HKREfu4hrsPM3QDyFawL
7U5Z8qB/0fPyJwDgNJfbaXBu5UhJdkLZDAJoeOVkCynFFmX/eo4nP3GTtuuc
k8nwC3xZzj+09lve/PZFe0mYHWQHm80HFJmkY4c0k/MSYh9iFIhkj38t93G7
1glQ8ea8Y07V0ofMZUackCEtRT8vpIDu+uY7UeGWeLDU1XBAC/oeMcd2fi8Y
sJekohweue9unE2rPnXHPSpsj2iDG4oXUgfZizwPYDxXNAvkCCMbHmWlkQh1
giHqIVjqGGqACv1PkcywCLDGzw0mJSpuf2jCBBycEV6Z4hoap5fZqfElv3/B
2iqsR/kdGV8iUQ4HWOCX507HcVGFAXTolFvX+9v+Cp9ScN/HO0k1AFNCPnti
tSXGafKB0kBOmy4kdpAdD7ULWi2dmpkhUXr/MZPQXkYBtgfagxr2J8xhS5NI
Di66ZzUtXxqBzxzRBdU+5Qlbuj5kfMIh5UAWVXHCcPmBzaD9AQeuGKYNn4CD
tz9Q1RDjsTlQGqkNBS0rs/vHSr0WIaqpHmabVXlu0JAuWDTugp6+yWfbje22
wcq0r6w/NwiEhz/6b/loDj+nyqAilAEObSzdh8WPdT/hQR0Dl2e5dfshrIjK
mePuwcgLJB+EXvBgGZqfVcMSEDAGjUv5GonV85CFBLfFLmhdsmRS9yq57CwS
FzmqOnjx+S42RZ58kePRp/GrBfzfb5iwyBxp2KakrqHD78HjyqBtF7PgpPEm
Ffxz9EJsE2nc66XE5Dqtmkugv5/mVT6AC7R/tiTIdF43romsYe1eGLpmFVgh
n8dluDHUjSLget7Ss4dG9G29AOFeOHSY8sEI2mtoaLETSisR1qnmL5Z8p/cY
3QPXszmKfPruyN9h6nwcDBsQNLC//zHb6OaLSfHr8PNvlhp0o8JvEKPN2lxA
v+LoCmIOvFrJGyRfSFn1YFdSmdb5UQ/7p3620wqoiWNsvC2P6mmApogIFuwF
WjzoGBg240aBnoM5TZpqzkGtwx1PxCdWuHr82yT9dF7+Rj1iMzicY2tIQneb
aY9bytSgtVsuyjC+4k/wIXmvarmIH6HQVBMzdyW9y04fLJiJKI3LNq6MMXS0
RO8Vm1e80zpLKXBr7GbUL5vtWYXe5mfkBplMVZzvJvnMOxmSOwtWg2prRTMm
oviZcAg8LqkfKOhLT7t6bzCmgUkKp5PoKN/gNy1UvLWL2ti42Vd8gC1wlzfG
pUF0DjzvEEgk6oByESBXQExTRSCN8eejAHREbLVDlKhNHgoCG055M+JScNDc
VNTg788eEGM5gc4w+GhgRrX4gTucQicyDHuO7ZOaQjFaMDb4FzEic4ioxix3
NjeDPKEEPoKuEelOQS5JO2UMQikRrJtUbNiOQrJdPEndE3CYyCrBOTy5OwNa
9jnTaxwFfbt+8a2/rEFrHxFlL8442paq+0ZIlgMCF+SVDbmrNFqC0EteigeQ
fS2itk2Wtq+62NbPXCPuYnfs8yfnfcLj63THDb7dzko1pBoqSKrzCnO4DqQN
+9MXO038QPQU6b8QX/TgWwW/NB8sMCtQlLecMOWwHCCuTLdFCQYSM988vXaB
rBW6CUklzqEsFivqxLVbdHRv0S7GkNeqDYoIJRfJFIkwYK0ocg5+KJMDJXKh
M3F0EXuKhb6MhNyWK2oqE+pdLDJjnd4wUAEi2PxrWcSfCFC9HTOWLzG2waFD
9at+9bbMSc49QzLJF2aWumF8WB/epKwU5efFCkcNIREPF0l7gifm42MMEPvi
cP+XDIp3ud56eZOkRGpbkcNDh6/0bzV867UVAxP4TnYrFNE02F48C7bz8wpC
mdnkzlmPJIFeKHaCeSpvZWg2QzPky9ZDB+qEqV0dUZI2HTHIXrJ5sXKQQdKD
job1Kq8TPZYWdV4NH4PF1ILbB2D97M53kBLecnwIYVx4hhdVJSrFKXi8n97P
ZUEyLAnVkzwaHe5BmMskZPkr5VhDYqrvoX3GYzVFv7dEr3ivydAnMseweHTC
0OL84R78lcEmpTmh0ao4FSFZSvWBOOPfKxZYW3fFcUc6/FdawTufnfDJoqdR
fjwmXSLCWSMVZbEh3M1FGcSwcuOrNoNehylmv4eNxeHK++gGUUWMHSpRIG/K
n5WVT2KRya/7ywATUR92Bqml3qPZLv0fCLL7truihYTJrItFayoX8pCYF7m3
zJfbsdr230x9F6xjVPDdp1EPJiRs+X5XhYzBv+W9kyQgPTyjH8nbjYn7mw/E
AKWVdLKt9BCSNd+dnds9Oan2Br5OKkLOhbh7490KxRAQxTaJuHp5bSsRsXn2
pJSSXuLRIsVDu0a39Afl3to/wsfneqOVZKofYNcoQTcF/HkgogaXcgQL53gN
jYB6e4TEX2RsIcT5GHuZo40BKrepF8brOWqqM9u/cgsuoFp2dxdSAHh+TL1T
j5oDJNAQsJSoY1YalIHNSdmy+yI7My/0Hi6lRM7Nd97szLv/ZGbHW52pWv3F
oWx/U97E4TQYIXBalRIwKB2O9Nr6p/UOvLfmlqC5bxtDRCFdy+tAqScs+zsu
IePPqBuEFgFq18wbEFTiVncPI4GO++eRmmOVdStuXTk4+Cur7xZ0ehg6jdgu
/h+8wR+wzb+leIQHyTgdsS5bqwbZ/7rdfrmtHJYj7OkYFDdbqGGhglPHZBhl
lohrvQk2ulshh1RZ22cHoqKDcGCyr8lCX4FTg47Oami2/OJvH8KoErtXGiri
PCz7DOYGdMy1wbCi7Jw1hisJKKaSYrfaLORe1gbkZBsx4wPSfkBKY/gWfhAb
wk3eVCV21giNr52/wAtfx8l4+w91CXOunM5oQEGmgc7DxgKEQD59EvQzhdbz
Lx20OPo5tB57j/H0sJFekvoppMGgkaVLjEGlCdl3jx/87P9vs1iAbw2rFgjd
NZgFAV2oH90QbOc6yQLsaKaXod5uZ5jO6LDTf519dQvD02ozBiQgLg/DwsW7
FiteU/q+TIjlXUa7P+x7fosMnXxUwuYdDCkHVBDSrR6iMfgtrxHW0NHXCWsa
bQqu4jcOnFurFBW07tAcpViZQY3AOZ0wEO4prn0nebF3DH8g+x+NX77KJepq
I9Oy7gtPnKyFP5FzmsLcghK4Ah3cRQ2cJVZEyx71Z3Id1MAsSlHFK/Nbk1Pi
ibwqjWhlAFr0Ptkwcv4K0vagYRDmEhT1EcLHajK5VIt2NC9sRECdC9dQTZoK
Py/DqHyWuVp047AFNOH04a42VU0F9ud1KauTmzdKYYzE73KWYMLWcVjoVAuM
ND+ISmsFpIwK6sMyu95xCeK7NO5RT3yv3QY0CrJzPvJEm3jE164L1N0gHWYH
xKtieWU9+RKC3Y7pSnkrmzd2lvCOMqhg5BbpJJQWfS+swW9EAAQWV3K2yJpk
P5wowhqowwQTC87TfMRxvRcZq3g3WtM1LfkF+4dpu5Sxhs0KCI5DhAV/sceV
Tixc0iNqZuS5QQSfBFrWEYarY0vIMthfl+LZNeZ0vLhnWK+SMQOLQuBPYwCu
siwXpspoP1Sc1AXn/Er7vFKg2N7RzPizNCeIWSspXTmIbeCr97HWbvVR1V/s
zz18ytsDE6IOy96XThEVXQrKX3PojgQNL5+9B+ygjiT7V1ToOLq8H8fZ+THY
lCdrdGWlUZBO/pViFOGeKeSjqCBqEfDNzqbDabcuRHeL0Dg1DBJ7+xvtoTjg
tVnyYuGcra7B31svCO0dn/E28xXOaKef7xFkKttsfsluTYTvVYo+U6fdH4ZO
LS222x2eZW/hn1/11CHiXJ6NwEwW+qUjqONNhCUxM9MnyfIyYGEyvVo4c0BY
5ao8gc90xshuVdVQqCmlCQSkRtpJEVdEtoq62NHx9DahyNe5tPKTQRT+SQEP
zR18yYQ0nA9cJs9Cj5WOMWVlfdH6dt9e6FnBROxkzepw1+taB3ApG0UiXasZ
4VbSfVNk1mXaXtFurUr9NEzaSqsco2FbA2x6p1AS5RCrf6+4HjQ89i9mEBg6
KoG/04ezpDOtES3iDa2QrybhfD189gWuS0Wn5ZhRjmNrxRaPcdevlvFhhsze
uH9MTUUpmSyaba/ZTw4DYUhRlmSIZdL2T7Fj/tdDr7r7sVv9UcaZ8n/oAj3t
CKL194+EO4XJWeOHm36pIg+Hn99DmjozdBHkLaEvL+/nHabNv3c8di9EFnu9
mzv4VZU8/rrqvS703zkc346pzTum9f0J/XtDlsRQmeu7Lx9E+2+ujb46ABdA
mSbFdpntl7TOiH7Q+TZ5+1Se1exoruwewAvt95OJH87SpGaPSTskIk+w4uIt
F2SAqAnloKam+kTtQCzq1HnKU6KRmnlIe8J6hl44TXWJhzmyY0fQNcmE5Iya
6KY/P0D6X59vhgs31XOl2ftbEdW9+FmTTP5gfIwwrXrHRTxV3PPh/GDLFRLE
9GdBg7Czo8eewaq2xXSSBvBCK2sRWrNV2BbWHQbm4BSabcmiCFpt0+OzvsGJ
8IH55BzWff+w3xf1Fy1Cg7yixmOK3kNd61drle1PwmGSnrpInjT+LpD3ZflM
fT6BLqYN3kxPyKkagv8TLudcj/0/uH8xsQdYqUXJi6QD6Y7DjKjCjwAMM4pp
5wOsYsVLMghCqKehnHkpXetUfZbxkvk0/ZJMhKByGFtFz/qdJxvulZPJ7CAs
sZyCEDNLenBcaIDznd6+zyioLe7mEhooX1sOoa0TCPBQaWsKnVWwpWsn9yxi
KdlF1N5o0VQcC6eTu65eLhNVlUwuMxDwRiNikc12tzTSFBZ4Qx5SLwTHvdav
hO1IdFjB7bjnEDJfjXAwoFJFA2vcgU6H6nhZ3WxQkYsOJG0B7mtbLhNQCVg1
D06Jin3oqfgLhh/wF2lWiP/+7PPOrYGUd4loMm8fcL8jiQcQGPKUM7nFLOWG
5ZMADy9YO25IRTQI4S36PSx8P3I2XDudhBXp9VywqZKIF8rOhdeuwr70oHxZ
tSBe2LJSwlpSEEPS0mmVo5oWlAiT+WgcAKLIt7Df+OrLLUr3oeNdgYGJrlLX
cLdhLrzhVOru52639Xzfv8h6KDoa9ii0PCzocSYPokhGllqi0i6f5LbNFl6I
GGF5Ta6tO3Xv5ztRhYOX9DRwDq5zVx/tQNQuIy42yLOWvgSXmg92IHJq3//W
H4YGIxe+DHCxGCu3IFIPK1GkMkaOjC8YQK7glF0MtnsMtaq0iM0Mx6R59J1O
cB2AxtmQtKkGXksvWivCQfP0nI1IKd+nrs7jr4V1JfZoqcgvlx8zm+D5yFCw
wIMfQu/LknsOzBseNeTVNxazFq1PurpZcLR0FQwtwt2Dl7tSb7NMogszJjlI
3bihoKBvoldvM/tbBU+bR/ee2RjdWB5nU0IuZ2T3PGozcUWpTVHL4CR4cRjp
kYb3nuhjURFShFtm4rRdeWj+/NG0XkkCggtTz6uZYpuYVp2zzj7jyFocTjJR
BYXxAtqIghw/d0X5cupu7vPggGk5EhwFrt/xEfoCshCPW0l74Pt2AGm3g1eC
nQj9wKuPHhirCqduYPUsFbMypKpMKqd4+IJ9nwTppWA+CarFTYRXw9JA1wJQ
F9Y3lUet0dCFySxsmTz0b4HOJfG2fSV6mssBtcCyt3d5O2X5VL/ayp6PtZQ6
l1BOQ+0ZWpKp+19e/8nODySbEW7eBy6PDqsp4s4WLtrRpMEmL2sPlnH+3Peq
5Qe09itb2Nf7HhuUIzfo6vqMa/ctZQ9m4/ArOXwJ/UfuMcjAbklII/3PCebL
4bppc/aXSoq9obv15Yj05NWchWA4jcxSi4mUNi+VSJiO01B/37Uq3dTjTln1
Wk8sni4JTngeTRH+LXwswgdplDFez/uOgNpw9O5UVqj0ghZNd40SYjBnO2c1
M8uWaoU/BpLLEwCOR7Zl1hHba7tmLlmSjcHby/C5mSGaFtsHuGMFSwsUxv9Q
ssdt36eIuHY8YoT34MO5uc9D9YC8V20+akOZ/GMN/7Kt/y+XRPtpv/RMtPvH
BGnI31i8j0OrDZ3oPmpdpf1J5PK/XUwZRHfOrQqKAZI5oV7OzPOtZzF7osg7
fQ+i/a5PNL7tcHM6nKN5zs6adLb5VDlLrMPpqqzvcG8qPyWsnZR5WksOmsQi
nWEXyjezZF67ctj+MBunfr9rzod99ODRhg1WewpN8VsY/rr6uZ6z7KQSiapS
E/MtGjdnCLDnTIlrhFWlUl9FCbw99xWvKwjbSp8U7smQgaMgh4aBVGAheu/r
bvCiH++dBCbo4ScurpmIZlwED7h4lpmQR/neUlN3rxjz13CLwvQU5YrY8aXr
55dZ1DgBcnyMFoCfnQBtVkoG1YEXulg8/zl2qvUyNnMEheUROd09ITB8tJk9
jT9QhDw5V4uU9lZv3KJ/LYNnRJSEEOL6/jnSFG/xsq9skK34ykYYw+IWccIe
4L7fY0h/GDpSdGvyau2OBXFXUI22EbadM/NROyOqn0z7xtuv22XkHehXoV+J
NBh1SFUlgz3wZaIh1PFH593hHNf+7M/WdAi+om9nKNmpEZIPUOYfZgzCBxL2
7kCap22vjP3qvC4uEtdM1//WND0xw28YTlbcHJMC9EruXp8LL7fIqJE4mouu
9BxxZnCbSGP2qZdnwqcsWFME0bEm8iGD3sGu4mTaGA2HlPCFgbu+mXvt2N9O
Vha5ml9yeNw4rHHD3AJIFeVLbDgafIPpYEM/M3HKkGZCLH09APV2iMGxrrjl
YAYgZEwP4onBfCiH9sRustApzx7+hK615tUF6PMhCTa+isdkGYnTIwuUH60E
4RSV/rfkjkaG+O6+gFtkWDIXMf7Zjv//wXzJYI1f8DtloATEqupMhlQZPESW
sRJBRZ40V7Z6z1k03IV2bV2cy13XiFZ63locDsZOQu6SqMeAS3l/e4d80TgF
pdoteEdNY8kuo6ZFzkHaG5d1E16MEWzMYZ09kzi5AIRCIXZbEqTssTZ7O4Zp
zgpMTzaGv+K47Z2avEPbDk4wzZDDpF2cScyh/PdJRB+Ow8GijV9uLSi9A9hI
WrBsNLzGYXMzKA3K0R8FsEJ1EtBydVXrTVSA+USx6ct2fXe8wAitoJS6Tu1s
vuwI9fy5camZ3BbpiXSuy7/74vvseC4bK2Zu192mZKZGIWMtClSjolNN26Ls
kN1lcwyo9EPNIuTOC13VlQ2e4AGoN7Gyx3LV+hQyJ460/aqnT+AB3dQNPn81
I8ZuNJAldP4yssmZnViDbVXd5t7iKZHtJuY5pnseiSoKEODil38Dmlct+oEw
YNBbc9XNazhkVo197FHWA2XvKXD47LtYHkf3aZHYTN7cR9Q8TYBTge0QNP0B
Rzc/Uc/hVSCCQQTCMBKPuQhHXelO2BTtCzlm5GHXLgGuJmx2il8/JRfO9a+V
KLlxY696NxwuliYYQOG4hjgjs7kp33qeX0NV/rR0/c3t1+uJz15u2AXOG+84
+VGd7BHHF72x0V/YXS08GXL7i6HZmJtosJ6Y1Cy6MHWRwxWDQSVnllaL5VcD
nbyfdG6YrZNDZ8w7dnvLFh2Ympv74xO6YDH/5ADpsbjqr8y6uA+pm2hHuGT3
gjQftqpvdf1+qF4fC3uNRjc7wV+3MrN0vIO2Q4EERlD3Vw8n+wyqB+cOrg67
CP4kGhk6nbNttW5Tc1G83xAyk7/0n7J6sCKukYrr/8FADHCdeSeC88MY8hqU
kzF0tNUkSoxUFoaGt0Rx/tBqoKkiNmcbtIWmjAg0z/utT20Isr7rM06nCgmE
nyxEGKHgXQcMfTemErjw76UaPsCix+USQzdxvlnLLzwJ910vOQlytXhHxtx3
8jZT4VYH7aIsA2tA7xwcirCyAtGz8pGR3yz6vWsEgxKFVZ3N8hHiJnf9etmj
Y+ckGQLWI5I2suGiPZZinegQhQ1aJ3K78Mqfrq478wrMLA2gSkWBPmQ1QO/A
jxjQvzegdaU5XvPvJ8y2NtJZ4tCcUtfqXfA7FFL3eFi3ugTIiHq2KbR1P2HW
yM5MRv6UCDFtzxX6RheAf9omiLdoZWlz7csDKn9uAxk/T2x/BmzMP1hmPnF+
1tEV5BEpPZv7jpKxjnFakwfBQuP8ShvDXz29rB5A+h/hCFeAeZkG8PXz/oLY
2XpopibkUWoSuKmLgHiMnuRso73mOoymqgjL+b4w8AIYAR3qKEWyDbfNEblj
tX4o/mTCAJJhUJvDmQdYw5Vx+iLjg5+o/WbQRFYmnC/MYGgt/m0LCTElpT8D
mDPG29BLINjuqeq2N3QB8JLb/szGzdkcVYXyjkO6p8bakM3tOFDHXuCejkB+
cM2tqtTnPtG7pgFHQ9cBxkScXka2ASp06663IOxZiuU8x8AnciLl8IPdFmeY
VgVpU8N/c6O8V/cNDOFpuDU4495a4G7XfSORIq3KrJOxXemaIOgViJ1zAktR
rHOQPKUiFwRrik0nxIwz0/8ekd6O6E65l+G4QITq54dDUpHz31A+eC3KpMcF
eZbrrnozL6DNW9YwIlRhtEYlgKtn1zdo+uBJkS0/sCgJp1kQTclgxnVQY/AI
SaiLqxgdHvCNWKaX1C0EIEy7oE1QKpaq6DXG+gcqSz7AwmCMZOBt7v8dtYQL
h0t8abLN1SiOzq9n7AJJZHWfuPCchLdKxVnxr5fq8S3r0Qw2nZ9mFAQbIpZi
71GMQ69pZF0x41VyYdBiBZ9O5GoLujfxJDVKCw1ctV40swmtGhwA5hsKmIre
0zH7Kx8nGGmCqSUOnC76sd3IDUSQBnyIP8NdLhlu/h5rQog9rrdleYrLWW3R
iD3FY0AwHJbuSweNXCmV8unHY00obpav2FBbOXcoOwQVRmXUaWABd7sITuYx
moo9Xn3sdj3twGtTm+vAv9X9AYxmN75y2sNb67aPglUNcrAAhebjb79Ff3uN
foKZDL6d7LtHDYFovHWvg4ddX3RDXHnc1K0PLxZVtxVPHJgZltxBfgwcRWxK
nRWN2VXIh3XlqIWIp75QCupGqFYQPDvl5xRPTWcsidC96EJP7QQFbD2UeSpc
1xGakcfOrHPpeoalVnrQNBZHV1RvFOT509cz6Pp5QasFGeFal2ZRmoE1ye88
zJAN0UGZP+o0dZlV0y2o5YDQLJirPLHIUlanmIOC+X+G69mUSWoQHMN3F3dP
eM8PE45jkr1342Ccrre3MayQvQvPSkTeOlL82G/q08C6y4Gn8Wu9lJH9FhaF
Hv/3nDaAmgOXLg1mrLUealZfTOy54w0pwXBObEGbo7dEPX4oQetIAxAS5hUf
MtRxXmWat248VT+XG2zk9rvMpO8m4hJMyeRBf1YWc2SK1Kqy0RMTaJJDKAw4
K6ZKs+cB5ZEnk5YdqwczZq0UQNCAP6NS/9OYG329M9nJyAWIYD4xl4L/lDsV
c6/gUX4FL1bfXHAJCqHZIBfsEIMV31iwxNTmymFIZRPlK9iMUvffFQAGKVvr
jXeTqTmXrGg3HLJxS4Gb81Nl3aEJv1BpeLIuHuD7Qk1HnKZkE9C9aX9a7a/M
wUvA3at0sue+2SuArdZ8bkt/qZo4tPccEz2XeXg3I+dRwOmFsnoetorx/sRF
prurkXl0SC8djhNI2c2t+GdaiMedmZoi4daJU7VgXAThZd9KgVZliZt3dG1I
Rxw8GAySKhSIKZ9JHv6Ku9PRbSpqa2r0jIyTqcH8/CNSvLTkYhZJ2cgLKqWo
8AhRIKbYorwGkcPsCc2BnDfLRDVjhAzeFPUkaLKntSiED9qPR0WgmC5gZTQR
HCXz4IzUXbTLgWqD02DDbrEg6miP/IjDmWbzpbcDQ/XPHrMmBjH+Fd0fVYqE
UaIuCWCsA9eRH7wHHp83c7jk74tLqdL/oyq4cJt2OOHwzH3IKhaExM/QjL0A
zLbqZkRy1hzVMbyL7+1BS7uMli1Ji7fuznM9U8eoevat96/AadwnuZ0ndPds
//1XRwLUQhSvqHDMmRELT0RzvQ6Lr0uAqZfcFk+lcAJKGuBdlUCvrZEnV+oF
Wen3mmW57PLiZR4/tx6o5ND+i7KMGXs1TCfc42yi+NIGRLCIQfKG2J8wpX3l
+T9hIOWnbIN00mOH2qHDafapXz2HlUuDog2UGnhlBRFJtWBmovc+IxtJegoN
znqh9EUtQH8l86QogmfMrC7Hy4wnlB6iBDWpk4lrSjF/4tjWhlhORHaOxXiw
5+xtcfwI8BEwRJzvRx+SYY/+nxb3yyqLCFGUUxDNCsjpPoFosOnrYY1H2oZa
bL9aAma7GZ1ovodlzV2TwgOq6l6b0YF931hsfAuphZxEU4Q0EnEdT9F7U4qO
PLWDyNyomi438rtGEpiH7JfZac5NPA/g+wZDhxsHRMJThqpKsATm8ugcg+zC
9H9miR0TQ0nFMKYK188yNEYb41tKvmTPf7lWVOfvQ8tqKwsxPdLIUjx5dTBg
jl9ZKTaIiCMghYKdnZDOUc/cZDZ6xBlKSe+uB+TjwXa6gojhlbZFRNrETRgc
BsLFR1nZgbdJsBw3Xx2VXKKLDC7tATc4kBRXfgAenbSSMKe9VrXTnb4NgBdU
Nb2oWi+3DBUw9/rSdQT36bKB93h8MhOv8fQWOBIWtQ8Z6pa6uMV0RNTXqEnD
mcCND1U0i1Wn8QzyxXiH0K2xUMJoadaFod/0x7MX/0GYPf7RzYaJsSS2WjQ9
V7+FgQYTT42gjXFxYVUs43eaqCifS9/7ZN3iDoEAn0T3RcCmgnQNoyV4xNnb
VKLXazruoifItBtlWrwUsKcNOtaX7ASoXSrjJJ75vtgBQMoWqDiyxcE80jbX
ww6j020u2r01DJAb0vVGUd4xBY9/D60ehHRb90H9jxei3z4E4Wkmix4h9L6N
I6KA1aG/JeH+UhBZ2Wm2Gins0NQjN8L9q5mvPBspM8SgHKANNv1GoBs/Vh7a
6cETn4J3S1zvBYYFBiI655iQErkP175KjIqfugB1rEbYBkUAC3lR6XOTmUZp
Xzb3OH/n+fFP0hLe4FW6EdeeT37dyaavW7zlUt4+y1geLC/u9VPpI2B6vAhu
teYB2h9AXNVcwfihSoIt7yDYlxzqNYJRYgmSFZGscQjFjx4wq+MPmXf0Jb9z
mng7wIIpfI7OBF2ny/NX1zit6sXdF3DA3xQIhjTULKOIDnE+/fvLqvHjqwFA
4TQvoRn+av0HqxRWetaf1dvxANF2z1nPzMJn9MRxmi+L0orKInBnQYETUe0u
OKFngSeTfSnOiTJr4L6SrsVW8mK5g/52DOkK0+r033TAiQLMWDUux8eZU4RA
IKJ5DoYihUeus9XVnGOmfl9a2NN9SlLRoI/mu52+pBQcFWVwZEhUikxFGNLz
cjr6UcsVzZlbj7CZMESiO7go1p4B17n3+dXQMSc6MxNprPSUNkS9LgJGWXe3
rr3FX8HJT3iirsWbJj2IzNFIqogTi0zlkcpcFz3eY5bB8ex6lxQssfQtCSBW
SU24f1oO+Q0XsTCB2KSqS1cPKlhFDGuKimdYcaKyoc3GaiJWABf0tB6ojPIK
x6xiR6R+NjuCQ2u62dl8fnKGDIAlDfefsfSi0jZ2suqkqRPlBXPHjI1U2BzD
lA9aVimA2y4JLkyvHUKdF3uhyNz+9Ow3BkxK4PUjR0I/fRSHTa5GQAw3bJn8
Kwh4P5ldoH83qmVrLpq8gZfdCmeKIXjG036TTHDZ1x2jpgoVcOKk7ztimP62
JWwdfiyV5d3fnagnml+0Oin51YaX0I89atfK/VInL2WdHDuyotMX8O2EU3We
lpdmMLUInCsYS0t47TH/kfT5Z63ynhF9O6Q9AIlQL7zHj2xxOd6JG8U6EReT
xJJAh0WKsI0MXfx7DfHX+K6rhQKr0XyvCOH0dc1/8TG4VUkKAGF/8sxHNIBP
5wUyF3Wqbumb5A2FU1bz9m25UXs3wrTQSJnuQQnP1d7B7D18tuVv6YRk1AzE
booFPQzKftpBiTA7iRuEBmfsjgtERoGRKQ5cNINpgSggZbY+ng6d/pVqxZpZ
6wqi3A6UAqPWbABXivacCS7QxHwqysvfTwvq3WmJk8+whIwXhBz05o2RMUoI
Mpv6lDj/zxT8qXW4P6n+cwZv4trkoCnfm0qrIroSZC9uvg6vR9qX1kUaKgT3
rWTLNYo+j8spUuBl+EuVkcEFgM7F56RpQ02MIrljHXrlei6TIf67CchAz3XO
BCkBu7vYN+33mh1sCb6UJgnx2CgOY2RH5dUdUC+52SIEiZ++QjdxEmwFaVPN
+M7hT3eh6X3kHP3t8NRldNjADX9GkPaG+HngiWjMRvf/B0N078LHiXeYBypL
2phXxz7QHgmQJztvyOB/XGrMDoSZNFbYc5GyjfP64gn32fYLIXNNIX2bOWuf
T0rfE2tO7DOk18OtClDXC7pljATQ+t0UgpT7ZTgYR0qlcoSbeyxVmcjNnWp9
paYPzogu/lftDgvshNc0yLy4/ppCUth4vA0ygfU1GRCboSJL4XKMiLNM8KbL
AaNsdVS5TVPvtdhAKBSfQyVDS/cro2KhjSlExh0N3NFRaVCVl3QubH9hjDxl
J6G/2moUelUoMZz5ayXOelUTLv5QwLGj8y+nfbnWUAA32FjDaJeilG5o7L6T
NtzhSVDLxNJaRz0BhyuJ7oio5TnpsUYvQWBESqrQ8ViuM6TVULlAuK8UX4FC
QgQUrMbvK5NX2rsoobbtY3TMmZCSZ6eL/Dv7T7pKlv+GE4mKcEymMImYxS5K
T/H8+/zyh27TzvngX1pDkxWlVAJQwW1v0pWRQXuVhnbG4J/0B/P0KQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1J8Q3byvF53v2sd4+6+D04309Txcpv8zpxrIycUcY6DKBjxjFkNxEznCpPAsIBVRAoa94LQAog7WOrJIRnbb3BzUzwtYWP+HRzJFqI9jxv83EIPeMZgC5+2ZF15Zddk2FcgIsADURpza+9Imkq9HauqOtDd7UQ4/HUGtwo/CdxfvRhUVxBfOkj0KWZQFXiO9Kw1dxFuwtEJqEoQfnToKecvaSiSsdUvdMKy8tOiPx4xGgPI8RPSdg8fpn0CRm5shK0l4Oq0ba1ZIysH+XfvQ0b6LG/JAfsZ7fHjU+K7luX3FC5gI7gewwZj907FEifoOsSgu+aX4C3xBCIl9/afUVsO3l5umdSCrtI/k5qEJLV4jj5gk0wyqfbNgw70aUGD6BcnS7bebfKElatnNqplSRB3EqXAGnF6A3I7b39CNyNXdc0eZioeHsoKl15C9ApIjUmGZeRZUjBoZydcCzDVdU2AJ6mTYI8ePej0RWI2jkEBDSujbeT0QpswxsBtxL7dvUChf3afXlrM0GYhq1Bn7iYs9uDp9mcSTFU9BBhwIcvuG2joUpYnD4vmTX9KAdCyk9AOW6w5p3VOPTAKhmD2OphxFAyzr7GOPWwGav/Eh4Dm21R++MRro+O3WrP+vM+jqDpV1RxefT6HoQR5+8nXpli1CYBLCRuS3h56urcS2tpliq09luBGat9mecjKca5zVURYUBME0RcAXxv7YE0KldAXOMOlGttLhAoWTiVMi7AGfoPHcQSTyMrXCUyonvNnKjRRqA6gc7uAhO2k6r9Qzxv9"
`endif