// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RVflY2cG/bKwaQbsQCpioqjr3fimZ9+jwOvuXIFuL8nyX6NSPc3rGxm+vU/l
fPqT6wiPpIASXIkDIHlsTloeyfvt0/kq3Up838juOV4idUttWQkia0m3LpZ0
Xrw+aK9LQuKrfwoHu51/mkF8jAVO8IupIyFLMkE3tjq+0Z+WulHSo1SptH6V
7Yomvijcuu7mhnfBTOh3Yz3H+Csq+XudSbUL91K6sldLuDUqKzdP9yo6sxYI
0A0N7rc0CYBuTtSoijsR4L5EtDLP0crrCuExJlgsDhcsLw+hdd2tb82vJqRU
u/6bOOSKVR6AVV0rstM2JRgjoxrj7ruRBhz3wLM1TA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p6e0EvC7H+RrBLCEsf1cqXNsjzMJ8nyR9nTBRlIuTGEt3NL+4UA0RFS+YHfP
FfGrwrU6VmpzW1zALVYN26VKZuKy/YI1FkU+qIooXXqLb2YA1IDT07/2GTXc
4XuHO6rGPGjnXIFIXhYZ484SX0r+f4OYn3N7aXaZkePxmVdmrppWznDrGuRN
OyXpHquwc1/7txgdN1wP/Akn1agQ3tI5gVQzxjVNh1zNzpMLpWqVCCpj23qf
TZn46Ta2sKzgvOKKQvpkFZEuN+pAhjbjqlg1QcS9xpG1c7SVBFJSnYgZntiH
8oABAPcJ7uECyQ12Ig3GkmcXTzxb8iX4c9/cdw4ElA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BtKkFFnlctMOSYF2ILIZepYed4cI19BafqvVxjWEfmgwNjx45IZz0ipXaFYT
ALGchZgaCyV2JnaIp5xqejsOUdhQaQ5hB6+eX7qFjjgi26TAM/rK7v+k+iOm
x+R8ByOadzzrgLVBc4+KsJWPKgAd0RBqon756s0S//iWSosfLN99/AuFfRPr
kaGaqDlI3NnmDM7YFcojgZDjBquLpafJIwVxmoN7ZXUnKtp1EDslTyVgxHzB
IcBbmbXg/pBmqSjGDVjvI7ujXnunTwaENm/zJQz1p/u3XuHtIehFvfrSehuW
ccn4GO4JcNJ8trxKZi/lqaxezbHJVqSz+KrJbdx9Zw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NKwuWyV7FnDaqdaW0T+fx5wEk0zTi4IcGcYQis1aUQs0JuAsSvi1r6QKbula
0B7L47INL78u8x4Vfs3EvTZ8Z2UVJibfqC4HI5MOcw5g3NBJhc+S7yUo3DP8
LgqiyO0uQ14w5qXBQtdlDtKRf5Bn4g67/lrkIUayVeUj8psn1qpllNebBh+5
1UWBpPSc5d8HJTfSxI+ppaT9cisqYh9DdRpMOf69tTdIftjlnKqHo80e8OB0
0xcBZ/XVP5uWPq6eRHCQvxQNU3OGavDs3RACLicw7Xa6CRMHWXpZGR72qmwc
iH7l3J+Z9Rr8SWTWMznZdoKibmdF00pmtomJAiApdA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
N/Sby0Cm72m/rQkBeG6RsRzd6vS549RF8iyV3Wgaq6FCzHjcmMYbBvDdUYcz
C21vakho2Bx7wS8n3HSHQ4xXfixoHAAGhNxHAXbrcUDkOLKGsNu1SPngPhnQ
ScSdS7awunM+SZQEbTLkffKBaNizzB4RQzgfRCsX5Yr679oWKZ4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XchDhxx06ZoedTWAmC5gP36Yuyyfxb5UMGKA6mA/pu+I5RcRk6h/4ajjCW2Q
5sNWrvCENE+/mQtcouK1kqBuBVjE1BQsNe3Juo8eW11r1p4XzhbXG7dUGcQ0
pW6ESXOOhN0WiTsXn9P3l1Q9vbpm3BvJJ7NTjXo3+RuzSjmlbruA66f8R9YK
eUPlwl0gRZBlJ05FTaO3kZsHoyuBbFVUtDFwn4AQ23NarHH2OkEGLBuiPVbY
ff/QUVPlDgY3Qnsx0YgIPF6M6wNHT9PlHzTGgVAZXj+wuyqHBoR3A8JI4CQL
cORM9Wd638g9SzdYoQ+4W18xGukULL2fVfqTVSj5HKEM0Qs/uF8X+k104vK/
/GT/I/sK6z2VumPh+puehFqg3XAvhZjCeEhYhq0UBuU2DIisfKfKtysuGS5a
ds+difaVgKYx4GaXJqxvqU71tuvC9Jsk37ifyTJZxRjCN6FGzGL3gdE4lZJu
uYbY7mcRJqFsUGf0vg434zi4tm2GE2pD


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cETQW1zAlFuCnoCr8tnHXuQB3YFsfc+L99NW3mxw13iuEAECF1BSKr6Qrc6f
2XNgPzH9r8eEBLnp6brk49e+v3TKEefKxgJ7aVZf3QEMoXzkauhRQNLIL2HE
rYckv2vxO8wNmVjckJ5bxwdS2yxQY/9oTMsjscKrpXYogJsNzD4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QKLzAWWqpoM/wqw5+ARYNYIiRKhCoDi5gTq8vw2dCe8sFZrmTgfnesmZTt4v
6fCZHsxsJQgsC34kBITaoDYJX2Ed4KXfqD7c/W+8tqsjr+B2Vwk0ImWUvFZJ
JGVsPhhS3Me7ZQiFIM3SeaDgLdxL5DOcdvMgyJ3I0oYYVyPN9Go=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4608)
`pragma protect data_block
qe6FNsx2QExp0kp/3m60HvPEP3W7bFf9M5NSNXJCy+EYQtLmFThjdJ1rNSv+
L2aUXYBSGDjhadvJ5MXCsWBKR54UBk7IXxSh0//YdsX0LFKpqjPRapPWYmb7
p4yGDhclL/EOfDDj0XpHdnMhwpw7W85IuPqSsPR/JedRfybPKNLhO11VxNla
TbBfp3KAIQBpP50Li8EA7O3MRvalCPxj4YHvzjBBLRzqp7aQoxoEaApTtIb+
pncGEA3F5lS8R7J9F/qGSbeGQp+lkFxqh0PWWmynHop8zl6HxkGeBBuJbv4T
lBESAozi5qlOO+vjXTRfUs1cSmVTARqYwFBez+VmFMNL0JqaIi9gYbJYvPCu
tIuGeYhhBob+7QHcE0/sp5ytOevjP3Bid8yvf8x1sv4/u1rfCjyG+i9vORzh
zFtqD3z+lHDs9e8lgN14VkktvjXJSDe/KZS2hOQVxmN2dqk/WzSKkdg5I8xx
s7kOr3a5mhuw0luDJmBM3Bppsdlh3xpMlFePC0ImZI/aTyiK8KrPWWoWzSgz
vFy5+VoEGclWJs62YSEbIH7xJzn9aQeJ2yeplJqO1iJmqLsJr1vFq/AVfcHE
m9sopX28cczzAS1uDx2dRM8xn4Fxli69Ht/UhTCOrOQKlgVBv1az6uuux6px
+ssPKoMDUYSnEhLEB923rurcqFRzcBcpci70RgfTsrE2ARyNP1iCNcyLOXHJ
sW+uFsI8VIQD8j2NFI0la2nq/8gNyCuBerLRJq5NDhTuQAr9jjceveI5P/Z7
TCbmI5T5gBiDwuLGfdgrAaopxTIwh+0WXNny5cdZLmzKM+wyxVfKx7b5DcL1
yi+BoYkf/xNQd2m5oFHLJX5KcE5GXBl/l4yLICPGcVfsR6UIBZzmXgXgoix4
9QKM4Tojb9W+jil+0ckPTUFQdjsPmNPGQ7pR2T5kDMr8o2E+orYdYJ7xXgcb
Tpk4uS1ZYZwE7hSyB3j/z/KzAlE4DLNygMbLnTaXwDfKEcmR34azJTTq+9uu
XTt680yYy6prGNeWk3AG//SFJfiOTRYBB1efXNSujxQjc7wwpuGU2dl7Bmsz
GlwswlCGzAlBHF03+oomHe+Ko8kic3cooVnOj8szuZkdKJ7WdjpDnoIgNFgq
8SFv8CidmjSAFIQQ9Mj6IPy1EqjOby3caAcou0Ld3jZfQ6bWD8BVK7CibOl2
RWf9AlHU37PLEsfY7TsAzbpnEfQ3WdxPUuCuKkKXWg+LX3m3CrZTdIIxmWID
suTgkPHOBYa5AEGIC74Ig7qJSTIN44Nx3u2zGBS/J4VeA1Txy0wpf/D3lgSO
YK3iQfZonV1kNmJQRC0ftH+fr36YS0e1U5inWLddguy+tdZCMHbsm4h+3J7a
Z5+28KfF1DD+F7W6VGG/oEkTpSGyRLewKfkuTnCiqDLnPf3bqqGqIj2TVmGt
FrwfXuyEUrIe+U1sDWqFsfFoJUzsLknjwYJGjk8YuxRmgiQwZKnDRUKZZ6BF
04oUN0Trjk5zBeDijj1O/QEheaBub4dCeXUliwrzqWvxbsED5xIX6LKM4Be3
xaLWkDv3qkEECAFzS6o7gs9ZaZqachv9F+hxOgQYqKvGRkPKNrj5ZXiA3I0j
+3F6EB3fGUqLCMQcDaWPDJFUpoaZX8yjrGAqnURSTS9YBXkdYs4cV46OA0wp
8jdfJNEhZo4r4YHxLb4ONdJKd7AQihnX/hud+Rs1aHytaL2359oZnWd/2rit
gUBubbA8+6+zLa8ABORTNr6A2nkAb6kIHEgZnyijeiQNI+j4vZBvjK34sCEv
q+/JAWrftOfimae2ETmdsEYmcgFvAFFe234deqiOjV9fMtqY9sJqpgp3Cb90
SkAPbsUbZM2nlU7qbTGAeSuoNqgTbFoe0+NWZEvgoBct6wqDogl5UUfNmXqz
fkh34KVWE7E3JNZXxf8kGVKmwSB5j+iZzK6KxxQKJPf0dp5ht2z6aWiI5EhL
pWWHU5iSXU2JYw6rKvPSAPNJmhFuoJpXOorK3D7qNttYvt7Uf8QWw+c746nT
eNCELJkZpKL2HKCHW5A18vEHDq9j6c2fVj4TbP+CVILe2y2iduBKYrBKbeTI
4p1hL+uNFulq/zBF1GCpGYx7n6WFcQYSHXdJT79Uw3Y0p/YpIv7alrJToZeU
bbEwspPhtYpSfMLTT2HO9V2JAPzKcM1tJuYPmxDZzEqG9q/ZQcsqcDqyzznQ
GrU29Z0bXJuW5A+mgW10MegNY6Vmvco1b5JKtl/2mRIxO5FOUpbUQvyyQ4nq
WaysEweaoZ38U0tK8F68jGVQa7+5GdcJW262FA0/RumI0fg2UyQ63o2QhWm7
U6R6XO/0JbTJEhMrgvqdCjnZOa+q3FbGFKkizdfRAj4+ZW99ujZ7PT6Ua3I9
xMFzRLDnH+sfciNP25U/zDumDeLiGdFL/tSqyk0SP2IKA6kutgeYvYbEU229
3OFQnzANpHalGf/mznIr8RhSQHUbcQHDsP1E4aVfxGwA8ODKrSuee4PWS5x+
QX84YnvLh/vyhxQVG/zoEEjuTNWFlA2K87sWCBoaTyuJDXhHZBFjvgitLEjZ
R10DQqmbcdbKyeaJRBetAwwSTORhO+1jnDtcyzEnenLdnnsPwZlNAX0wgsbV
j/B8t9zGT4fI2UV/EMucbaTe6tyieZ0gfk/tuOhWWVbDOdtezXgOJXV4XdT2
klQjRLQgzo1RMcQqGvwheXYEqXP9WLOFUaofFKDhxfAiDTKdeUOymNl0F7Y+
DcrQPV4rYQKdcWlZdztk9a/NTFYe/+vLy6jF3o0Oo9N/VFhhqxQ2Bzh7yJYp
eOaAjdOf4sdgsN446F1cGk4h5q9tzek6MwIUYDyfEGj9zjsyD/51Q+LTUpfA
X/ilWyDzGbfHYfJhCD4oWSlR+cbJessnnSrVw+Jf/H5MIJ9uAXAzNQWQnwa7
3mkdeBix7hI77uNglvBvEYn5V0B8Z0BDWpce7UmGrZAaMsvB2b0O8uyosyYf
pUcZMCQqJXrUV7nU1bu2mRyZ5JC5kPlXwh0DeZocR63QiZ17iEOPQCphg49q
kPHh+y/5iMBScCEshSWCEpFMA+OfqvVynGBKnGGcSxlYTc1M0JOBwDxBj85A
TdrVjxkyL7xIX6z+NhcrZ5luG2L9O+Jb5rMfSWZHE7FhmTkEc2nJ+5PazHX+
703Cp1CvcoiBlH3zILmwArGDF5sp2psTkAFP+AzsplseN/NrGw0S1pVcDNK2
Jr1OgKc53vXfMizY70KXTumMfckWIrACEjcV92y+BQqlv3a7fy1BOgsfvu9/
Vs1oYR7o4NXMnkPy5UfpoYjQYSx3kz2j9CVnvOw5b+DlYxnVNK5i/fC28vOJ
+0Pds9wuiWOY5aXKWjaE7SqGqLjunVGGyC3LtqxjBG2Iy6b3b1RnGkB258qj
zVBKD94hvhh/kVtxrzmKEnKu88FeQjfHwHk/Twi4SHHRFck/ZV+DftwtWoPO
Bh5WU5GqKG3XeNg+T2wm0L5qVjd0l4ThdbT/KHKX5xVth9PAm3JIemzraioi
S4w0KPkGBWdyULwiMXoyLLvOs8/snRpyEBHbEGiBLRLHG6Sib51Y9GN+rHzH
sTetsdDBvLdn8xpfXfGYNW+Q1YtsMiYDdp3gpSmqYX/SEXOHMgMjnWOZJiKe
2h0XmcclXhhQYB0MrdMSFSqK8e6iHH1YHwMTgihXjZhI+ZExlKx8kk2RrFhp
xhea98IPEP5Oaokkqw49HmqLJa8RVWrwI6LALW4MFwPbdpMLsBr7Nukx6ztv
35lhLYWPc4ivl0sQa9PJsIiyOO0F8uwvYeCpyCx9BeWwShuaHAVLqPiwBYXu
LEnyFVV4kTFskw+YJPSbIuRgwzQuXBGrbx8fOEOO9gVszFO/UUPtJKb8fD6o
pp4+ZbNOjWK06pkvRRhmlKT8nXcD29vPmVdwbda4NirPYz8m9/+FcvfsTovK
uOGEDpKGuMdw3ZoxVMSbSbWbIBpiep5DJ2xmYKmj8l0xdQplQkWzgjoszVpf
QtJcO1Wmy4Tt76NTP3Ub9zr7kd/yipiOzz253ix/IHstk4c8glItXw8TmcQl
Uqn14Yiy+/H76OTNypxPF8z9qk81Z6j7Po7x+u7y6VytPHpRU8Zq7xcnKghB
b90EZDEQATN1cqqU8yUUpK049l7iwvpPAg/bCZt0vhGHaFggwRVvDjIpKs90
bRzl0sq+61U+Og4TCV7zv8jwTIJBZ7Q7K4Amr1GHW9sgasLyCwZYm8UwKWvN
/Y98hB/8uYYD1ymPRgy5ulS3wyivIJ+i9Ml8xeC3nPM1sXt4XTiET0CSivKs
k8MiViiRqXmKk+jkdraEzOjPLZz50bSyFX9kO3n5EFWAPg/DMlooICnSkthk
RRd0b6beQep+xCdezFaATxrm2fUwk0/2wxYdzej4IDiNBisKegZ5qYFK3x9x
PmDRAMkmtib/1c2KIj6AD0FNTaQPSw5sf1sCMp3j0Q+E+u+yj+Y7X6hOochZ
kG/NXOhWoXaaw86C5Ey+AuJw8/jgguKL//4lAqUepN7ayecqxOJXCppZ5k7z
vp8fNKlEliANPwrZWC9ii4OZ4HeYoYAKprMmQznqe9fE2aeX+G+vZ8+xbFqF
0HRCFUh63Wf3ocbYn/+uq8O39Er+kkxKBORTzGklyciE+J/nG8nj5RGYpYcc
02uC2BN/ueqq7MIlzJJgzz51nmFVxxK8goosQUVcDWYozQBvIhiYl2gftfxj
imxGMjuB5Tao2COxoJ5ZpOwI7VZ6rwuUhJoVQJJtsP3Iyk4/ys1nKYr1K0d0
8OP6ke5jfxYXQwU1MPiQU1FU3cHgR7iYeFtyZEmytIDTEpHSiP6piiJk8VBC
j1bGdEx92AuaM3qyJx6VdjdoW7b4rAXxZ94mlOKdGi/1pHBvfBkCjMk3dC51
XWmSlMGW0M2ob+uBReoT7UUL9uN1kBNEGqnyDCOyIBGGL/ddB03zjVAUSv6Z
AwdxLAziwQ35cuYod67E7liGX2/5D7/lJ36vvUGUYhtvtrDQtWB7LE2gZcnO
0cXpQapkdyS5TnMUrOVUv/4BBQ4ShDA72s4MOfS9OOC3JhpqsJN5sKd+qJYK
H+SK0/Q7fyUQKrYIUBvFM2y+urp21bBlt3zF2XF0PpZOHbW6wrt4T2i7KnKF
a4wI2AYITdt5N9BlTK26nS1lrnvB2cunP4YYCIDaU741gHZUwONFlOOZpw+y
T4K1Y38JBzcTp5WvZwB3cOk2wvFtlskqw/qBORuF1zhybpQzqKLOOCBPHHpG
1eB/UlnVDc5/Ils68edhBzxNYehROR+2zEOqP1BcP2ZzbMtoqgjlphlQRjb+
Pvvyt9x+Ea47gcNzoR8krD93Vbb0NyGJO6a6Yhpbo/NW/lrYjF72qmAJia+4
Z0+9nq4f92SFJLtdycCsqQxd1rJvSUGMUACTxW4E91079b+zHrNh+9orwSmd
KJGYvtxOEewOM9HesvPV0MOPs/6b43nDrt1AIlktXXv/Qj1u1qvt7RVsOdUG
GiJgSjuppN+yhY8uU5p8ryn5TtsVtOMLZLny7WNxSBb4JAKTf4CnrzTaGSCZ
XedPk8lLgcaSOjsvPiwirzCRbR/NjTUfVO8qWz5OkaNDtFr94hG8gP5WBR8e
7X7V4CB/4ELVGsqBSjlzXG3zw8Ts0H6uBJgKni4XEnOHh7SGsjuoHvfrUhGy
UaBy7RTpELHhrZJ1pU7rzJL5HDb+xyxyoiP2298TwlZGpOtpv+9c5RzG8tLw
OJB2l8ccr8WOR2wzHAc+OK5Mb2uju2ihG/7p2dg3OuJQE/XVffVGEC0e8ny2
7MTKX2u60to9vxKOlaiuAagmEZ3aUdb1bDNkjgSXLfchi48E8H8Oxrs/Nibe
AkHeAFOQLsb5vgsQoAhMIpO5lhuwnps9OD0/oUJxt6HFXml//w/iipAQwuRN
LTuAf3I27DEoq8hKDeiTEv6jwrOJLMHSAKTQzxhXNBjC/2KywxU+xomKkPP9
K9qcPrDGVBP5Ow0LnrMnMJ3fan/uCSRrAw738WuA8OSWcAwk5DRgJXmoxy3I
km7tDnkMg3VPpv8a8lCSoLGb8Et0NDF2QqrqRg5+LMQf+4Hs4JP7Zr/sCfJm
q7KjYfwkZ0hJSdv6KmVFn7sI

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzdOqwUn/VmLAMj9NlYJ1zLukFsgqbr88bTTcjgJNoe2dKM3AjMZTRh+ONLGyyvBr5FF+Mm8lT/OopgB1SlaEzMSEitqTJbFWEz4PLPUzidH7nXgGeTTCGJCwIkQyLJxGkoM+nYhGWYGcA+3ZhgjaKKv2C+owhdtSbFVk6qtSepCDDq2yjf+AcPb/S0zZF/5f47lDDI2BHyamr8TzzM/2h+sMVotWPICB3YyEhgUhfgCar+9eVVTI+p7D9ZKcUIOwsNfgsncqzJ/IJ7Xcefecy+sNW5TwBsl9/arvyn0oP+jGzdvMMTEFlSRlRXVxwrLz4bRt+tvKgvPGTvu9bORRaVLH7b5N5sLc+hpQfzmUpovCkQUjE2VA+ojwBAzlH6x0WKKsdChbyFNiIwAr2D7rmPbezGSLvZQlJoMhJcTTEdRfcaDIiIv/p4Fc0qbJSl9mTBt1i/sksPK6EWFnXper1aX6FB+wUOjwbc88CVj4cE/opFgEL2/sZ1G32aZxBEB2h8PLozIbY8u05KSrtJHhKiyvzLlUCCZhCYtYCeHSI5naOH0aUHGanPTiOvKJ0T9RjveGCYQVNd7tKwybPYd5tPPRtGMYjaVyb9L7vBLcOASuGqD9t4WWw1dRfh1O1P6l4NDBhoK0LiIX8YALUDhep6WW51tcWWWb+NCW0foDpc5Bh+9Knulg9tSi0uZBHgRoBKWOsX312b/F8EzAOnAI014kvbLYHDcKgOBRQvJPtDfEo6FZ815BaIxY/7IKuw81NQyVw145zPGClRUTw9fjoaq"
`endif