// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ou2uGVPSob6RuzjUrE184YfT0GqPjWUwRQJKeYqNXFBWnL8zOonoKLpAGE0j
VmHb+RFTQVjXcAbLXXGRzfOacOB3k/n7jg8rdvWHHWpRsqCsmGXp2VzzRT51
6pzSR4DK777AO0ewVrJp4CqhjvFl26JWyWM3NiXUhPaipG7VaNmjPjxhDlik
gKWlVKWymHOcZeSu6pdVK36IK94osftQCAjF1wbSczgvs+Xhj0hFLLFmbTHM
gg+0dUiLQmkck7mGtolTfvN83n5hvJ5fAXmvOSoSTMxVMtnEmMmFTZH9Wnzj
kuz7aRefXJV8/VR1XzLKHwHK9riT8XJYQeLpyLBJSA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EGvcui4+uvDeUcWT6Jls+pNE8zmId2IFTvFItRZnnfV6xIMMJYKiQSm8bk5F
NhNgPOe5SnaCMh2B5T3ZzXSg5kYWYxJdm7ifLgkI9267As0f0kCri/0irU4p
kEa8L1VT9NJXFa1LkBoyVahTWVUeD5ZtAUFTxubOOXpC6vEl9Zo+v3VQEdYi
WRVUPM2owVoMUIdT6QtO594BeM5hz9hGoVfCZVWvYGRc6zakUo9MqXkj5xA9
KJ0kUI4pR8/ddlroKQitkOfTY6qG4X4RtLEbDWc469s3S/MWGViTG4S8dpF6
TnQ8QwOWz8CWCeooFYWdVXbChTjuZ4uxo1fbeFY0tg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n3UNdL22KmMyXpZPayWph9TJgBv7u+8J39ubUo0TfbJMBex/wAMHO/PloeMZ
MXMZvq9D598UNhhqlx2X50fgzNqdHM3LH5sK01kwQw8cDCnQyeVRmLbKwJLd
LwatlxbUhMH+GBVHiwjCFCboIUhmxnOOIuYK6VwuZZO5EMRwRQGCcVP7Ha+W
M4KZVXdR91OTJDhGBH1v8VeQEwZF1Q337L+JWiSR48pkhL/PetdoIzkqoz/T
QS91+RxvUPNZeI2lC/3/vcAGl/JCAAujot4E2mRE4wuLIzZMY+PREXP9csWu
7XJdojdUASdUCZ1GiH+42Oau1iTShtfLZ2akY5m/RA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Mf5mDP6nPc6CPDGj4d/qcXBj492MmbDjqJWlGqtqmd013QFZJU0K30Z+DS0M
XjoW/y2tYhoKV/5CUYDiDouYpi9S0hxdDT7zUOPsNBVe2jdv+4e+6pmy89fA
U4/DCwDsNyCLA95/+hsb3Ct2fKInPft0kjwm1NHTuGzqoP2Mn2C6fQpD0DxU
AFyMQtFWYwq+7i7SApckHaqioegVCc4kTfxH0E4d7iwibL9Vfwobvkke5Vp4
ePeL31ddZLNkWAjDtjvku5U2cC3jfwdshBCwQOGcZBW6ovJ50UsmaOM+M8s/
k0WosjjBV+1fsnUKsEeLNNGsm/zTKY833BO3Oep7wQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m+AHY6cghDtj/HNwwURKTEvzGYnuPaXzsD7awpIkEghewufcrSWb8VSEzqpq
HDC+8SGYUXtWxNlrKAjmCKAh2dJD0bKX3F8FkWO61YqF9blHspitdc4l5WGI
5Jtx0iI/QGRt0oyQmyUR8DWZB8Y7B3O5HsyFts1m7bBnBNuV/90=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vYmAxxBN+/DVyO32WKq4gZNLHpsFvqTvUgntGxeY1PwLea0vtjVDZ7Hr5AXJ
LXNBlWm9/Cs+0vHNuR5qcgAny2fpAco0CIsXP+ueypkg5yxQSmA/nJB9kN3p
TkPdfDdAA3xcI5K2a75H7JYSVJFAEbCK5YuEyh2f/Bf6yNyL9E1H045BFsT5
q3PpHE/98I/i9XGxNPTjXcfBGQl2rko5G9kswcI/5DD9TH4mo9A38MixnzEt
uMFV3DYNryavxs2r2dWbMCgNpYTa8t6YX+pMsgi+oy+FofucoXl78qAuwGRy
L9o8Ttq7OPGt/z2wRQH5sdj+Ly3EV14534GJB95mg6OF3e1qAO6ax9rEbmGi
oHgoGMR9yHPrUp8/IJsbAAXwgCSnZLg0J1b3LTJ8Pqk0aZzJM5RkdgxMSAyS
ak1BQEBpT9GfAUbygt1AD/DB8I7RlK1f5srEKdo49gUlf0FbeCTs56P08vEe
XVTS56jxfcLrsgEp1rxdYgoVEcfDecg6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oGPXUs5nx84jjsf5T8196WWS5tvfYLsiY4wo6x7P7oNQ26448nNl0Umzr8XX
tsA15ErLGoEV5nlr89qn5lFiDUB74Tgib78ytQAOl36VzNbR/c/HRrlbOc49
l8xAYpv9Mc7LOpXifiMWgCiJkhHKGGXYsARfS4Q7c30Tvbg2/YY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ijOV89x8uVQrc5eIXzR69zYMJm66rzITeYjsasGpn7UWKCro9eEJG4WqZwob
5WOV9P3GtYHTFTEnHg7iH1KZwVTkORwk48oTIHTe3LHyTOZLEseO2c4nc1uR
exAgllIiNTe7aFkhsrAE11sZR7nq6Mrqb3+iawHdfepPZKoRfQs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7824)
`pragma protect data_block
PIyp+N4HPRz21NHMtuOUjl7tE6WY0HMd86WI2w4pqx0NklPlRM3+e7MQA56d
wfwwWuENuL7iJha0B91nMnstphYZ0b9bM41pAHFfDwDopI0oCVNGGY/9KxIG
Tp5qlUGQwhicLAJapIKY+DA1n3KSUpX/J46XXgw/CPq4YwqBTwC5YO1oxQ1f
2P+5GJDv6YdyjmQFA0hnlAg6rXl8m5Q1kVisKM+2v/e+r2sF3U2patdmlG1d
EOgI48EwEDtl/OWEjqjt3O73tY16kR64gO+lI2MtUgENRjBlp8v4gES7TroX
x0KZqj8WpzCrFKQEENo5iezx41gR77qKGalhhBRGuxKXlCzKwg87lwk+K8To
zgHp7AVHqMP1oQLiUiIkMwMShkXqEt8KtD9keAsAR5hM8y8ge11pJkErulMT
Jv8lhBuvQw+nCamBFElWqiDHU63pV3+XpsMymgYHZ67VTbINBWrkfJc4aqUp
KYzP7nHpleWhv2xPXWhmyM2QxwLvzrYpDyqsulcQPuaSLpMWDso51/lrYDie
i3VxLQZeFRy52pAsWwJRILYVryyx8KoXk9fxmm/k76d+jTDbeKyac8+BCvJy
dEOku8/DoZVN05G6Dwu5Cc5ruXop10dR68c293sC9ncGFbD19YfSNIosMzIv
l50h1y7Xil3i4crAXZya7Cr1FwkpaxDlPFUOId3vdQvGCrFnrwzu5mUmNHXB
VL+LXkV2KmsmE6CYvL/egcIx+G4T2JxAN9Q7KeX8yA45G4sibkcJax4PW/Ag
nTxWXd7G7W8Q5GWghqjDBcMIQ1B9Qlr44h0ivTYI1x5HMP8OlJcNhgp7N2MW
/L7cHcMBhJB0wNObbJ+SwOynlqfuHkWr2Q8iNnQJNaTKzCd0jeq3maT4vE21
kF7TxrGbD0ih21tpNLyPU8XXMMFN+WwChliWUIoGo87jRo/OLPvA/sJcJAcN
OoKvxckbD54n8vTaPIYFvdiEiAbozC6tLPdZ57lmGVbK3sNYs1Guh35sKM4o
+i4xYqh0D3e2px/JDV+xH/pUENyXEC1v424WGk/iWSdAbv50rVa6yf1Ndzol
UcAkUsiE4puYQspr7BZNK0duW93flBZ+2BlZfnEYMqxWLzsIejjVP0lNbWNY
unFATZfdyN2JDuZudmN1HfHGVHQ909jHAvgMwXm33XuVuc1SUpqryFOLvdPj
cj/DUYn8LFmzO+Zj5NME/1jRGqImcso5KGUjSXz7qGcqVOQIoNShr3OfT7nc
BwOmEoGafXMKLX6fQX2VRc0aZNIU+N2XunYFFfNjduyIxpN9vcVx2H5yhrx2
YQQ6WgmWDAAzpFfgLabp7s+4bi5LCRTtCfEq/jdlH+gOCTnUu0Y5onbrhPsm
JFsu91sUGU0HEtm7ILzCisR7o8Rs9im6uBEQx34IPR7TnvysVxCfjC9t014s
9e/xRwV9ZS+fT//pTm1dX8NTr+Bxj3PhigiJt5Iq9kWjO7sgxjhqhIKDonUg
6tevWP05jmFs6dp/F7dGUMG/ZwEbfrmkqIii1KFPl1SJLQLEQU4qnlgZd1EW
8LgCZ9qPiNIfue3IBoz18tY966wEfIEi3KIcah4vtXD2jsKGYF/v5onaRXug
l1Bar/zfm6RxADnUq7fWVbZDBI+0937JmMSCCCjI4wOib9FARCtJ+hBfSLqo
8arWqslVUEIruR0u8HQcGJMqWoZVTmnXCQoDaUeZIKqjrjMvM5sbmk24Dk6y
o2upsyaqW7hqGgJtbsqnppnB30aaelFbKciVTx6a7zMtAVOyOY/LIpAe4+L+
H1s/3lhQQWLRqEUx8sXG8FP6kYCToI2oCmvEl/BkzosNa2qGp+Ix+I1OJgVr
qkMd8JWGmFjYGBArvBwdrKLFDanWrvRGkHWEhds/9GqP1jfbQxrGd0O/WNJJ
evp2sXB88rgzsdbos0/o0sqeJYUcXwdgYSiPEyLCpREGR/Ig+nf49/eBhink
jEG8xAUiWVcacKJ0mxRcXaIOb6EyH3lM5ogAeNkqRQwB1POO76MIZPlBQrTz
WlSc5WL608mdIZ/pd8rxi/voId9aQVoW/vSNJJfO7F+PHvjXyt41mH0zbDhg
BPLIppyKIOWfw42GV30+kIeZfxOgRo6uBP5YfhqdpSa5/bDNgLWeWRviesVj
ixelafeHgX+2qlUazbIYBpESn4AJd/vGW0EMiFUTqu6wXtMD3AsMH/OindeW
ITlX2roigi8LXi410HtIB5SZB0K7ZQvr72yyWsC7A6o36vYhZgJF4oWx8mKk
/5bwvYmtSCFxoJ63yCasffSLNeHChZbY2gE1oJ5DWa3uXtQJ7S0w/Su5igeM
es74iTibWtmZwwSwyEAVkHOFG/2V0nQTpCHzzYLjou358OHAD4nn0KTgTVx6
6duMRwI3AnF9uNo6CeMSoUSD2yrWRHmrHEEQbiH9emZ1hDS3AjXydH8enuGZ
Fo9nr7UaLnZO0WtlEdV2zWo96glRU7DNYMRFyx4WHL5ETXpb/eytX8tGx3oO
0PHUP9xYQximabpS7ZEO5PLDc8wYZ5Bksdi+aXQIzdzKwbIUio1S/JVJ3B6A
M/FmtRPDVggW7I+uvg15Doh80RVUwUhlp9FQJyCRbxIoxfZ+kVC8+uhWlLNO
psnVjAssXnwboMsu0ugdm/WJ6lfZiO4ZmlR+NwhXCNaZoUL3m4UbSqpnSh+m
SpvZrw9qkbD91jrf/CjktQlWIE7NeHS0BcLsTsi2iJR4Qf9HyKBH6bkyXC2e
i05H3LPjXo4Cqz62bzC3UM882mamje7kTyaFg+6Rtc0OFMlS1EYeHcb90CRr
m95xxWRjtwKK+NRRw57qhvu9PxbJPYO28hXfxKDVmmI6R1CdyRK3B2nNZhz9
M7CeiXsNpUgf7bwaPyhVhdRAG7+H6+f10EeqqlnOoHs6CVG599wMfKnXR+9J
K6cIJUUyIFLYsl10R6uy66pP9h8POBh40LooeuVZYmm+BgaVBldvKvgr1H9K
l+GN/8utPqGog7MVIAHx9StwBUPh2V3jkbwPxWXZmNpA4Cc8eA/eDsDOqQkT
SDW3fCAY30AfWsE7BkGE7snbsiAycIzPrbozNXDXQnEJPy/++G+9noNZTZaY
jwZBLc+HjZKLv4LmH4Qv1jd5gTiYcgtnfua7k4uKaNZ1Vko8mBRBAzP7K7nh
IXYQ7QhPviB8iLEaWIndX/dBX6379g8GV7F2EWajJC26qQfllSadkpJLxmPs
EZyDcFxh5c37gFxGhoErIvUXYGZnizi16cJTKU/lgIBw3EnP+v86jcggGyuM
h/ZRwZVB1gL0jvVujvmaYY9jM+I36mjHWxYhNF9wSuqrvOs/7Vk0pCv0oQaw
YFhOYPqk++rdyq6uaC2fN3+aaORS7PfGNmkBnzyJb6gm+o7IaWXgHXbEtQj2
CZD3EmuKBEj/62oX9YiicGI5CK8Quh9wV/PzH3W3a8Uqwg/Axkcs8Ap4Gf1Q
cIw5/3fYVDo12l+M2Oe8Yl6m0GjQp+EOEZWBjxB0SObO/N3Xj3s5j4K7gS6b
jdbALpIWCoaTgxMgTcXcDrTR46WeKfVZUR5nZY6KoaA6ucmyNRj71ONgqyRi
VcJS4Pu8iqYE9WtRb10rC2lzu66QMbZfotxE4Zal5jcKcBJ9Qe7LWx4K7o18
7hRUcTRe6FND1gai4uvpNSmChNI1qA5kVTm7yqhX/IB5aEKRz5eSG19Bb5W7
8omLxHcEBP5K33Tm7ktFoh9Sg4pWqqoeN9QOjJWvWt/9NPy8ql/eAwBlpQzP
MCBEILVQbRzHg7QDxg4psmJZpeRc5Gg312StKzzj3UC17EPAm7kG4uEcOHju
YKLBo6uF7Z7gROWaku0I/Pc87JhjW9grVZ90fjag9wXo5rdsCHRSbVwyoMVD
GbluQhonty5AwBdJL2186t8Blo1LOuz0nl53seSEb4Ne4PmsXuJRHm/JsMTz
p8sbKHyj3Rvqaggs+pulYE59dvu3rFLcwFQDAEwXNdH9gJNt3cNHGwJr+qlK
Ch/hwJTvWPL3q9SuZaugQ3xdTlSQkXMhezy/GOZRGT+Tz4ZaXuaYBq+dInzH
42U0gf0QbndL7w8nNffOvzvbPvAt4iVDNVVZq5OfdDeR2qDAxehz2Ir6CcQ8
DKayafNg6Oh9fDKAr4Ega8zwM7I9zbtrmEnchv91QMn51NuzKwXzg3cAij70
AqS1GrQmNMXIlTR478tJXIcjKVgmHqhG+JP1IabPRkB5P0ogkIPgx+8s2MhP
Tt5B/SHNPAtA3OxIVEqMiSIPaOUrHUVgEtZMES+8KICpN6FbIaLZx5Iu3G9f
vHAIpQNphdAbg38RQcgCjcGjOXtAji3lNNgmyAgolRg/idYaWMrMuBhUCzhA
0nioZOkd9Guzxss7vAj1cUo75B8DurEBWqYwRulcluKt/ikOpsVKkbuNhq1J
bLukcQIj43oIovMnxG7Y7JrkdJFCo/YiFLQGWRnQTNWMbnQDITFsVxGen+Kl
dH769tmBgpKuYvY0Psr33rdVL5tXMuzQddCgvRwXImsNoQe67N+Lmr4qDML5
7M+2Wh8/LNSH7naJE/vNQ3ExHS2CEZMiohEF8Z3ldSwzNfindS1TZA+H4uEN
nm2yfvG+GVXCgnCAwpN9Gi4ZoDgPuwxngR9kbKDB86ceXm/j+/YWI/CkMlyO
wqdtxeTGD14cIHanwSxBWBDC0a1ARGvXpqg4p3wOx8v9dLnxKhoCTI4taAWK
dskD/xf78qcQUnrMtbKoOIcOrMFHlOwERHCAt+KayLwQWHzIfwcJJJHnJdjq
MkeQFZ2dfkjo8zA1pkhi6r/bTw+LSFd2O5IswdYIdo0VducIXymyp9TfR0By
AYEN/Y+zltzmru4TDTf5SW9dNa/bnEIpvqwR/vdIPoCtCorwiquGegK5n0K0
B5BPnVrIrl7NWoWFFGP9Nu35NFZFGefLAB/PBKDhZ3URO6TLDzq6g89aqSUn
XhrlCLY7ZwFw5kEqAh7Yok4TdkAUt0dLATsgdLmJrZ9kPwAVNSXZMCJzxTJu
fgvdBxVfvTwFWyIGb30zwzEwuvlx+GhN8EgYoOX2nDQI4jAtVPqiDV/RQt6j
25r2lDdIzdRn52ef1tgIgXUzNij480OGlXxN0WFG9KSITZGS/qrckG54BpJg
H5rd0tBSlHEuB98k0qDZIk0CXOKibI85n02SeXtaIUTLU8sJGfpZfWtHWvcD
iOkX5AHdSJPnASRYOM9kAWC/3NiEoqRwCtBuM5XO1ejd9A6AcA+hRCTxR0YH
t6YYf0DFdi3ycLNHq3WFdDAoUDjYJokNHvAMG+pVToRmqBbjrRJuUjpLx6Jp
T/CwtpCZTt+fzLp6BoasL2p9KOkJkunTdmtKBSROwjjfVLa1mcM/wYX0ymsh
OZoDHw0V/ytBoAV1jd11UohJc8SHQDcU0oBFBa6PAfdFPS0RUNFeaS/2Exrn
mdVqPLkpaAJxOSXyUxTNvAIil4fnEzvMBsX8PxHd0b3gEpGfXHljsp4kYolx
LPGSPFewcdfgls7t/CTITyCxDHZHEjLT8UFV3mbQQ7A6l6suIPNUsyE27BNP
kF9RqWSWStl0NDU6CAKt82TPcYH8iIhXNb+CO3O+4kdl8L8AVEiJcziuUOgh
DQNcdpT6+XePi32I2yfnZogk8VSHrmEJJ7INucLRGQyaG/2LC64jKW2mS/WX
DDTfhLjvz6n/+fJFXb3LCeoKJTJowezSW+tIQga8E2EIdkP6fmL9NZunphYO
/LtdNq5fJJwBXDJnQg9lkpB5uSFbbxsGa7pYLg/IvHnvwz8fxYACyXDNbxzf
GsEaSz9TIvv7YagHuL34YJcSbL7THqgR5akMeKIOpXWXjzVVPqY7Ek6JSUEt
Ua+E4ItlG+0lHkiopZN3P3N02OTRHCURiI7itzp8Vy3PxqTd4PYz/fwlLD+9
8Qs0qk7Y/3U3TVFDhxuvitQtyBcyEqOubHRXzyHP2e8A2q5WvHSVnbT0n6+2
nlI4gMBDzF8QrvdzVwChd8VhisUZ+R/f5dhQ2ZOgcV4ctgzcoB57Xz9bho5D
97ehOXxEFC8krcSkIKmyUCPIXNQqXfLQ/dvaJmRNMAjOXjeE5qnJQ+nDiznd
mKujzWpdGNc4ifdY836hZ7jc/VXcSX3dF6Qp6x+mB/qvRNgGz2xFxfUvF4F3
cYpaUdYNuRKiADkrCNj7ipe/Ibw0ig8Y6X7AFYrwnKaQfu42PTMjcwA3BCsZ
QzRn0B/qj2f9SunA7t1cGgrx2Iol7YpktimZ/5zpY+wQ5CFYnEMpXO5r0BMy
C4o6PCisRduyezfRKnJVn44qgyQNPEabHrgZyW5ukCvUmWP/PYJalNkUAjWL
FwGg0L1wPAPA3eUwxH09y677vQ4wkqTMdlkI6FVrwHbHywW0WXje9RA0UoyX
O+0JCyEb5vA28LugeqRu/DBsD65ZGEeyeDf3/4dHkAn6GSrtj6saJTN1UbOk
G1ZauszO23JDH8tW7jHNKWPsH6ImcSgR0DvFFbOdWjk2jfA+jrWq8rJhTeMV
uRWY9/S+3o/BHVKLJ2jy99Aedanuj6UIwMEgaHfmkpTkSStuNC+svETrdIHW
2qNyaSauFaZ/7K/8G5GGFRiMAgE2fPRA+3hz2ZWpveT1fTlPgR5Y1bdVSXzz
CXUd+3v11o2tuC1XaeoNEeovBGyg9gednWkf5/vMAwN6M0yinliUqGicSfb+
34ck+Cggh9HrlnDyiUDouVXVjd1UnvV3nzl4IBw+yZsMxSQww/bi8LGXD+hb
bVFKF5NIPzx0x13JmqMUMLgHgKZhIhBUl6eZXWlSZEq/BRXkIRAV69bZE3w7
keMIprSobVLkDxoFlkCWCAetDfNp2dD37zRQgIuewTuZjOgi2q+tuvQhn6yC
TsCgSPC8fqgublY87O+TzKrT5M8ayhsWnLg4f+kdovIlAzCZXr0Pf4gvQh8+
iod9ZjpmEgLkZZ+KCZORmH8xrTmVAGI/GHjQQTUHZnkuq7x0cw1iEJcQPPPy
vCMBw6eZL0VdLM/xt/3nZf8M1ARDES/rlNmoGe9gBbvfm6hnLIjzeOIiQv9z
A/qgTyQh6XHlYcbXTaeTrgu1iqXAQmdt1iUQ9lEuNLEP881Iafbu8YdG82Jo
mI/JvmznWLz4w7phg/LhxhFmo3PDvuydscen78TIQdrvQ7YOvhwuLRjkJ1/a
2maOR6qKdFDOMvZC7p1CenrzeSfpH1mqa11R+wtfTC1zKoxoAwl17oxVKmLT
rgQOMaNC9pRLa+L52xzPyKQC4g0ybwV8v4PhoYFVDzB2Ck+biSDOycr4kOxL
w5UJVgUnQBIVW9usZ8sEmnlK/PqffHcF+lFEk0Yjzf5B/KpBcsbDuXWaqMm0
5LxGnh6J0hVJ3W2IsR1dxk5zXSRqMOIDelBqkqAHB60Gw2InnvIFScGTdL6D
QSpVljHJ8+vsTh0eGw/kAD55AKM+sDh7tf5MhCroz0K1dEAmC7WV2xPDBXDO
iu5tZ88xrsKZX8D4TN9LbDoAOhdU6JrG237/NNonYXFmoVr35H6kIebv1fYt
TDT14P+oXTTooxYOac7Y8fVxrwa6JjdDgadIOZVSeqpfe/e9090FRprN8Jkb
Nx7sXuuLuvL148DiDSjAehh2vwjCYUAQC+d0e8Mbk8Z9pXRuedEoNznX/CEI
pm0jPGe+E9HuhZSh0YB3BQYESI470x9VLIrpTFT/AXjdQfjeW4rw6aaPoZE8
BUcbNdL6JKXBo0iTDUp/xJGDEVzXNPB4+k0FHkVGeSdIdNMd1gd9ZsG9UcFz
FOOupTndUIhTSnKsxfFswas7SbX58jqHN+aFw/QuAjmrP/NrssBF1P29RwDN
AldYmJIQ/gYA32mPJapgmbELiQXef0x7K/fDlhjEX+WvN5nBDL+0wZNz60EL
z85EcWqdFXkop0p+pjS/6e0Eps3KIL6zyFO1EyFFIloeCAUjZG419YufSSy7
temNQZN3ysD108qYh9JGqa3mJLrFZubUuCQjJhHsvbi4LUPkQnSwBfmNA7fb
F/zD8fMjmfQjCyfB9KJK6k1hv8lPFFjGWDPfPqsM+iyG40YHXfBgEUIsz1Aq
PWCVlMuAJSVrRGjnDCfS/oFNx29gMzGzBKiu1tdgjagi6vVCPzZ/NSuKWdRJ
ZivWDvNHboVKZVgufHsdVM2V7muBdHGqvNo0A2kFC4znISjOwpjvC1xTk7en
vcT40Z35X7+iY1xvQvUDz44p3sw2OFHsvNnAVVbwKp1Iqp/vlxjy02G//dwE
cVJ3YXL01kqobZPTBfxJMI+utwBbYg9zXWFFaqNR5QwY9YKWhngUhcpPbOmm
9JaKez8UoDKs36l5pL+rkPP0Z2AtyzPIT6jnAGz07N+6L+t0izzJDMBsqg/a
N5RppnQ21Tm92Ba6r6L+GPPhKL9bxGzIkdDgDb70QYMtnulrIbZnQOaqdcoY
G+4spd3oCWwD+kHvFCZQGzIvYy+QjRCUmslcBdUnMQhWKGnzq8DeUPAsKqXp
nrnMTMcLrpN0FVWeZub9ofXy9spKfJ017FJdDjBv1u4AeNKhfr56ENV7f63O
b7aPs0J9psW8E6tQxSnIET2Mvgr1CpRk0I5C+IpJtu50SPGzDzW7Kq/BkDj2
U3irt1P9/4BzCY9BXOs3Miu3+P9XUAV7HvrPU/f4Zts19uMVOsZ6+dOG/AJG
MICdOcTJGrEsjbYEO0BcijnfbcrrtBwbqkJvViJCa2goTsjcXbBtLT+8l22R
KlOG9AHpLaCZ1Hv1ukDemFksc34JgKuwTrESuVoe+14G07PdyvMiTh+ZPTa0
tOAknAlCpgEpG1DhJOS/VxQdKAuCFA5PmTrA7ZDo51gdHZM8R77yyfgGeOJC
l/3/5AZBVsujxkqZuijhERXa3cyNmMx0kh5Ex4ooAE5BhpVXPHt8ode3niAV
WVXIV7tRIkY137CXZ4e2NWUA6lwhBfrxkKQ1T1CxojQjgPquNFkJRSIMxuRH
p5qqt2KqVKpTkwyWqc+XIzr4nmj4O/jP4yIxMnAQdN7W33KExnhKf6Qz7Yqo
XBcPe2TNtXu2f6qSO6mViTFZyKi2lgrLfJ5eV1XEmoJuPocS4tQ8ObIvk101
SDneaRJhrYGn7aq0ht3R54IhCaqrg//ofr19mKDb4WzVf+Wmo6DTB8Kufuni
VAQrJk1ojgP418JNBdwfCllK08UAXRmy7CZu0wVB7yn8JZYqBi7yO6DC4lEp
vvlsJ5THPillHh/vojIqVx6RbYQAolch+HkfhdigT3NR3tufE99T+NonwgB7
XGuh8cFwDDXyN+5Q4u4oHW1t30j5trRteikZ3yP40PGR505fEJk6ELrODznr
yhBVa9HLOGt50fnj76dKYqWQKywFceT5+RzYBFysM1Owffz7n1FB/RvDTZs/
iOwoTI1cpwoWT9jg/O0YQ/xLwaAMf+LgUjz8MECOMM0P+syabS21er02tAzf
9ciqPdj01vL1PuZDWQjB7gkWSyM1O/BYoeS6Mg2e/8Cduy5+jmZ114q8dMup
eP5sxxi0k9Zp7GNMKAkczfG4DYRxCvD71uuuuYJOaSWxxsZemjzIkOa8kKk1
7EQoBFmGK/iuj5qyD+RC3EsuQWc0sRUU06yEBTiAsADA1Ozwqt9JMujlfFu/
VKl8+EymG8xcya3d4UbPP3f45XFyak36PgJSrAsyyOu1rJVtx2X5UwSVNqEL
7WKbBxiybSa2qIOc2axif4pY1cicdv2w2epRQlwMMj7EarG0c92HWWSzQHAs
kKma7OPbhmkDwY8Q4PCmsuNQBp0o/K29vkpfZj3frlJLsqfsaCX3PRHvyNIp
T1bhlH2CNdG9BNM86vX/0dauj8CtBdxSa+2i29Db2eZkq719ktld1Sdlotbg
dnq+JpcLxV1k3MKDWnfdw0vv+gEigeod3AeyQeQqsKPL80LVyjcE6hm/P0Qq
oQRX2s3RTPirSKEDv8idTm6X3knfgM3v8CLi4PBVGBcoQ9v1ieXvyRPU/a9J
tabvjh9j0EOFCuVCrO1W3Neu38CtxwmIs8fDthT1HQLOXFGChz9CtiWsjsik
sUl9olV27QL/Lde1OukEJeX/3vm3fOMjm2X0Yoo6K6GWhoZtQH0jhmgOj/d8
7NL/uL9QnAi46G9rdjmOqXqecFdLbN0q8HK1jICGTcK4frA7vv2gX3IFUlcH
U634BCV7sVt7AbrfUCADuuXiFslhQVpCNeIiY8oo9O32hvUcFr77RSMEvLj8
tF1lgyqdW48QEGsOZw6q9wXUCtKxcrO1yx1ITNcjS/tngOY/D/j1TEQeXPqN
kGhQ5WwxRFUGB42cclZg0jwvzqNjgaDQ3oLNYBaPXWM+cmsXVE1UesiM6qQE
0qLytbSr7oPu5tBgLS+O1SNU+0j7ZlZ2IuseySoEtsEiGRtFnfnC

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6DlQtN3c58YHYHKTdniHBkbrNW28jGTCLtPExO/4NNl+ujYOzTQwb0AsrryQCSBDm0pTBg8qiHvFpPMOtFBbINplBnw8rsSyxt2056toWNLmKUgXhTpQVz3khQuSPACSZ9t4Cly/4WeYkSFIuoGv0qgYaBX9kKlU/7T1vrF2B707JMKR5NEAirbD4UIKVYQSTNLyk7BpvKM+sUurnwMLwh2nACR9bI959TmhvgWQA3emq2c7UxI9yElt6Iglgq8z8u9wZJI1mykcjMJyLp3dwDx4GxOjlrd6D8jnXugT2pOnW8D2CEykVUfi+b9iwXOUr5Iy8fBvfbpnSSe6Wuc5ouU9S5xEpREACkt3whhZHNnzgFBFr7RjInJYLb+pysIU2yzfj+sev4AvyP3anKp4TlgZx8YnP4sn4BF2I2APNZBYOikvnZX2SyC3Y7Lp1hdkV4bYheX+aeo19oERLJRhyedUQp1u/9uRxsa75a/InoojkNgvTO06ZeLViXycW6QFMNCx5KK3ZdiS3CcE1yUrl2cWHBB4nbxpbo0ZeLyRCQrghthsW6eC/jJStSn8wuV2fdpRGh2MNqavwclijfpqy2THROF2+WywjtStwRzpFzoEZcDsu8xCfZ9mBFFAfvvg3XRnSw6FhH+u6IQgmq7iOSELAfnq1BbY5l4vkqXhatD02xRiumA14U8HurrjvpbTldvLUNIEytNGdWj2YpyN/e+ao7B2w5jAKrlQVUel1/tMXkNoEYqg8QHIASpRyGZv42jTzyrlM3wZ90LrokKzasd"
`endif