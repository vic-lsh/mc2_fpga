// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eEof5BUTf+/ZtPzaPunbrrGKX1DUyr2zIhBTtIPyepoewAFUfphLhwRrAx5/
zLFXJK+JDo71G1bhdH0bpv6YSpNPCWtlF5ZgXtW2BMrhA0dwY6to9eF2woul
AfV1/PHk+cxdzIDgBjRF/vZJ1v26gLpi1P87v5SdUPf7wqe6E8rEaS2op7aA
v+o0z5p7O9as42jjfQchWqY1OTtaPO1Xng8qz9FL3F4r7emDikqOdOalz2yh
UiIfAnXyB3ZdEMCsR1jsGiS1mtiXBhYQQuU4wrTbb0xvMqKBMWn43eQJmNsG
B0uT0rAKUE/CMedd13vaC/EMWI7GAzSMDBTnDKMZgg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i3FTDnAvYdvFd/ZDd33cCWlAOUL75Gx7AwCQ/am+Tao4YlU6AGcoucrgyw2J
4ouJKUGt+ViQdi481gyT7jCkoAK/V7EiFJHknLrsUIa4s641C/rd3VL6Rbch
HYusG2fvZXpq7J+VqRAcCVLfW/rnsYXLo4xcIDgeyCEbwjlzzBczAjvehlX4
DiQNMJSGFla4iF4mOpjCPRbD30yjpg24m7aLf/MYoV5BUIsM7k4wviYMADT+
ScPssH4+WR6e7OxEP2GhHruEBsVH29deMV9lzHUq1nEKB3TfvEx/422T1Usc
hoJsLdlnNFuwTPhDO3nTomZjdjepedQhz6csKVKqXA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E+7ANv2qADYDllJZ7X7/tVrUCbMrFnDZngFxCu7+37ZbcDySRGzy2kXYNOzA
8fs6odmBWDezn2GkOZSDAHs8A4koh3xAG93ilvRlIkoD8ApKYgv+mIK9vEqr
uWtQW+xu/gdAIgBIyAt2/VlOdZ9ypgFfIvVZdkh1AHSQpb3mJrAzObxJfRqA
+inh6ihpe3obnJ8D4hXF4QWHU61n62l/ywEdfwpFm6c2jmrlMcciwYukMwiz
0yckW+JvM1TAzq+gsI25/B/GeaW1mthViR1RWg4F+5uMQ6Mmx9YeADzx6fKz
+jS2gL2C7vcqZUsmoOia5zGAb4r7HRVFBasm978vdA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ktcrmp5OETSRSf76w6qFL1MlTggxWeyEvAWwdaXEBv7GDq3+ysd3qmTgaiNW
wvQY3imRy5ms/M8Upa8DcgIjZNLMm4BRd+i+1aUZ6/o8Y1vBH7qLbnHkO7qz
ub6CwX4Aw7Fyj1Gb2BUcjJKZk2FG1Q080S4esa2G5dw2C7JKQ+NMgnaCXkZR
jyEtnlGQS4mWyYpCx7yw2wcUy4qHBSaSKKFnfsEWpAhM1UcmoMYVy1Kx7Ec3
tAuH7kbCBcZju+TIqWpWHNHuJjJCig0EgLfKUxDgmoBUQvXwvwKNhN9HW8s8
dR3e9cK1BKnTwwd6eUWFjbQCWs9T9qPfBbkQP/xOrA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jHoplY3MffXIk9sVpv+tuQWHcuUpnnQEbFGyS4yyHRPSCWZ0z4zZ+PcXmiK9
M3RgiqiexWvW4ucMSFwVu32EfyvkI3SXri2n6alyLPWfxXJ7qKxEbotv2QCz
ocBFVPqDZ20Js+38bldHXaZEpDLGSo8ee5oeX72SBmVAYXuAVZY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
megQPQEu+hnE0UbIJqjAZ0arVU3OTwjlAnoO4zPtArG891tlJYyeJQBKhHsn
WrYDo70MaNjzpQgLoXP1m/R5Roh/jEWBtMcgDkifS34fGh0Hjuyp3OpFQVg+
4KfNEHiGmmfa0raSntGb5m3PRVgVK+CYB885VoEZrw+B816FeoWq/4tu/RgZ
MMOuP+OxKR4p8UzwbMXxjCVe8x3cveFfrufVFmHwYLzzH75ccJibZoiclPPZ
fLfRj5APhCM4XOHAXj7MYvLP7KXRqEtfGwgHXoCNFhE9uFTEdr2bj/FXtsOY
EjF66xHRkLKkcS4BtJedE0Ulg8sUqzYzimEMB2wxPGjITttOdJnWybFwoqeM
ULpSaCZZIUOPOk0TiKBtlBmpEn+Q2YCfQxn3dU+tvJRbsmC2K5j6YDTuPs1Y
SgsZmYQRUKZNjWWU6PTcqnxEccDKTiXoVHQFf71scOIdU58P1pV5IQnaVLv7
g+XakhaCMv1PqLxqKh2+eBtbfU07Iri5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oqQsF/OO4YB3NJ7HXORY3P+mp3+MFnAArUh6H10LN9GMn5BiVTXg9GzHdo2X
UksxFHZtwGASELq6Q27rulkOcIYopsCgVF29i7maJCMIYD8MCYVRRmPMEdSH
9Rk0Dru/vTqzjJEJprnDvcYgDeIEnvyK0I6OVUgEIPG8v9y381k=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sUIo81OOx+8kz6H8p+WelUeemVyiQUvWi1Z7jcHaFf7mSvkdjDBTPtdjj24N
d2BYYxp8GRQUJAstmgfK09mCz+XZTONEkKNabN8DYzZyagBH2Efr4YWAZQOf
VYA8Ppn68E+1WEL1wgpbitMuKyvDzV/gNuOUJsjSk0KdeXX5nxo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 976)
`pragma protect data_block
CCUTizKO2sECxwpT+6KDQsmrBX8RHIkBO2aOBUBgM87BsZb9MeEjPOx4AU8M
BLHmfc3xHng8LADCSJ98SCJHCebYOUBnkCuaKun88+8u+nDP5qzwEJSiDZyk
9lkom6rSa+SGzAC0c/fKO/6bK5qMoyQisgHTfCfO6zT/B7cSxSlWlFAB3Jh6
5RbZRfEAqbrvmdB6vkYAZJyCQMu/GUI9hZkCO6AIG/ZjTyGlrVaGMAFQRi+X
MNILKyqStQKdAcdydtru1WYfSsrP0qjh8OJEURtjKDysOCT5g04eZcpFkZ0K
nSR+d3TDWQu2z1CviXOiqd0iY2fKHcVJbe9rx4kkrLods3qCpybhgZ0aRmGF
wU7HN7e8KwFs44bixlHK/sn0j45dId0RL6ADAXLXmm2ms8Uvwa22TjvoaW8i
yBcaPw/Hx+uQ73VDzdY7fV1i7ZRnMrxBkkf1cVp1wJTVvZMOmY4JiZ7GrtVA
puSl6UfO9k7Lnf+I6INoS1RLNROGCzR/7YUIvkojJoEYxFwu1LxzdXjQ5iP6
nzfRggkb4KC8FELgU+51OD+n+/aKDtaJ1EMELu763lLY6LrFXfuF5WNuEd77
7qxzkMDHltOMd/iRqZGdVJ8iak211IssVHDbDL/GGX69pD0NKrY3t15fWq8K
+2jvqw1SaCcL8U4HdXTYpIdS+TIiX4//vGqsSzA3ZP7ffSAQ8chrtuX6f9/v
fwiNyuZtW+agL6SLPgwRZ9Ogn5QN/BgdokqnCaiB477+oGILm7tBZJ/NMx/+
nHUXK8/W5T+c6/HQ7cGKsmooIlxwd/FTYm2DQcvwDenjzIyfFN6YmMiItCmo
y/XKNkowk7i3bklZlheltVbxoojNUxSuqhQ2kdv+EDc6dXt4gf59hTJoorDw
iLT4Og4cYNPeCUD5OJqANTT1oXI4XDYzlyAVNf/9AlSDlKmtQB8cdh7Duhd2
h4yY5VpcuDy/8RZ1VJA6YDPKq5eqbDnSHlSGqOMxFpuyVAsOD82TNNrjIW5o
Zf3qs5IIw5HcNmGuKwSaNC3Aj82005GstoVHmRYDc9sVNEsQu3dGRB70LaNN
fPEDXg9Cnl3DPQefyhkq5uibISbGuYxx7r/VKHvw099LMFpnC05EeqRw67Pz
bDgQql8PbedbLc4apfmodomSfJWxSTAAGX54yHbXURtKY4gfsGF6pmzF5vnO
RlSAb41Wm7PTjTFAI8i5t4xBbW1fhQuGuao+50yAR/VBqqo97vbDnI1ZaDrs
hnok5CZtO/920CRGipvf5zUCDkUr7EXX+GL6Ilh0hw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqcYla59qq9BXsEkWzzHMrLRhVkY28tWlDHnLgyFlBEfgv1ouvLUUBLeRNW0VxcNFu1pCt4FDdXovCFsDlvgibN/4tVSnF8YBLajSB4M/W0rxCxd/buPA4LEsA64BWTzi7C+BRmW5aIedWrUCMVPBVp7Z8B5KmRveejenGEP+aE2UjhOqvXqCoSix9rt08pyJnZBc6GamMnCJHDBvR1+THDC8LHvoogFuvBy7783pktDqPLMqC4zxTlonwp3Yfsv/tKUOV4f30ivQtQfHUUDIc+Z4OMcuNY0hI1qpDtRvsHyqJaxBhYc6lZi2GWXVF92cWn9RV+52EYBVYZRco2nur/J6ANuXAPkTQhrh9/ANhXcx4gNvtIq2d05GQ9XERSaIk2zXu3y/1wcbCkQY5uwX8hifGi1D+/IrGudfkNn6bK4Oc/73iNFluB8kfyWJwFWzRqklwjef2g7DQLB+3Z8KgkaaIeTSLNmuwvRWfvDn7rZujfIQ30R+CmSGCDKakXqSNIshmavB9DWb0psUhMkFpkPq/MnSfi9cAezu9bTbt9SEku/ED1z79GDGFNpwLRrlyhLVzWxEQEfr6K5+vzAn69H4dkOlTshlFXA9iszy6qNoqrwBekNcOzGGCBh0yhkEPFmDg8YESSQSkDPWSvVUanldk0XOqzIBKn9vxgzysT8m5ZBqBp8Y5vO8NdXPP6FITLq6JTjygH/7rwez1cj6WPlNX76hDfONCUBiQ3CaeAYJj56zXLn3A0Hq9Am90c7L9C7c7ZZrcLhlj9WjrpN86+M"
`endif