// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pgCKoywLrlCEOlVpNB3wfnGLxBo6qeJ/qePIHTnldnbcSqdXBGtr7zx9nzR2
f185jmu1dmg0YPuZyeN/bFt6gTKbMtQG1yd5MzX3b/3lQnS8E4vUkhpzVE1D
muaTavVBIqmVNrxl/qKKEGe8YHH3C0feB4Bsf+UmKuLRIVVgCgKRlz2uDjNf
HczGDuywGpJfFgPd5YtD2WebNDsnYTdN3zsbDFo4oMogpbwpB/Si4ve/Z32O
tJms59KJ8DWeatyEXZHr4MhrvripbYvBryqIKB5FVVp8KZdKNW+tLi76psCg
CvM/KDoG91KGBaUpWI9cPpBOpPo+tKhj6ZnlGuYWYw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dr85oOpxiSt+z6tjBir4GQxttvxFdigLwgwBJMNfK/Ug8SFUDDC4o0uHTZfH
xAwmATnHmYgxuFU2hVRztDd6jtrDPG8NBDF5TicvgyFUr7PVzUFhIH+nC/Sp
xBB9y+lhNmSotw+smjxuzgBEp6ez4STZQJiqiGbeD8R/hkI+7KoVEIyhQ8nG
rCKLTxUykPdimTFgFQNcBRzgCX2+9sCR5qTGAas2LYcnPUvS8Rxkexq/UZO4
/Y0SyfbL3RjXUol6tOEX2YvLIrquQAqnopXW2V2VaceGoSNvz9OR3QSvzCdz
Kf6QKeToaljiALmedB9IirDQ/1c/66aGJMauADAOlw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
efc4c4YsIKIN7RI4yWohusI0prAtCQ8uvQz54Ww6CcGjxvDvy79wDvzhV2Oc
CznYNLf3VLy3MnlghWYZ9aZGaWzB+Z3xx/h5sgKM97s6aCnW7DDiP6tinZF0
uKoh2tfL1L2h8K+j4DYS2xfvbTM+POXOJsCu4aA89A49/afCkERZwScNwLLF
uu4c+cmBRV7k7UcKs/C32mREhMCAd86RHXUZ8fqq48v377RCPSQqzyqnlmI3
UvqzlzBIhTI+1tIPsUloE7GBs6IpGR5RVh395DwJzLVkgnNsblSgDgnLllQ+
ZcFmSQxJw7AKhA+yYeJK4wEDd8Rp2MJVwWQqWcxGbA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GAwUBkkX/wAnxMDj/WQuHrDJEB/E3D+sox6f5VDaPA0pY54rb1+/OCNF//xd
fZEz5FTbeyXuV1IUuYtk0wxxtTyFfVUfkj0Vc8rNsf1HHvB8+lL70kyDSCAx
qCuI7p+4sIrGsN0Q3aokFjcy7TcHcIawBYIa8cOSzJKj5fFG3NTKWQCWjQIk
c09WNuwS7ldojLDJ/31wev67PcCWDfr8NNuM9NZBHKzyFl2AaAPnUOj4NV25
h5tVBVumB9rSVzumYGR4Q53ktwE2bXHLEmtLy6EEjFbQkV3UUcq9X/u6VmRY
qaaBU90x/hCnwxMwSr3o6S6AT3uevg+O1xFRqlytuA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
loPXQHRtE4KZH17IPDobCgYt3ybjWdffPsSgr5c0EBZhdzD1C+FmSaTn58gd
G6x9p9vHDG5iLrzKcxs6DaVyPzGKWxbzV9GVxzCidHDo5Sa2UlKO3fT+ZiSq
v79olHSaT3YUc4CSarSHsHPC7EvtUjj6z+qYDYA9CQ76S5PoJ3A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cHbct/gG/udMe6Z5byjbYYEYuErZ0lAJZ2E4QbTsakYb4xwxHUHniymU5/Uo
/FVpGCMLpBQR7jG0c5R9lI76j0ajk68cm4DIULrB3ajRjKCUd5LurCtTBHlo
buXsU5o8JgnRy8/CaEp5Fwev1UNvODqN++cKSf+BNPvcpFdA/w4eEnw6Cjah
p8t//sAkvhhGPaznLSJk8O36qR3JpUX5uFMM+KNjzxPggnE6WK8R6z/C3kct
utcTzZyXQpqQKPXdk7wfNuGDeGjOcFRfZ+p/FAazby8oT1KwtovVWzEKm/R+
jT/k4GTq+Z6229AKdE97W96x4WxYcDsazCucEz6mngPhJ/NxCtp7G9pjR+Vw
rL4xm2OD8inClC79mqRXPEqhZlBWLtZ78ubjNVFG5ShPZFM/osbhmhs1ZYAT
RhOYp/PN3aB0npVGj7I5sTwDgdxbDsp9ZiTK3nEIPjWNBbo51MYzRPGrjRjm
ZRGcmN0yVDbhSjFsz7BqZaWrQCYn3T3P


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gCjCJY5tOzQd5+aduhfkVkyaMNj8QduGslglIliehfrZ6KLA7J3jhDPU6rYI
o6yg2yqlfAR2v9k4AwdyhZIMzyknREyE0jPuaJUt8yUyHrynrh0HLXJBBVjk
uLfAJ+t87mT9nxuwLo+QxdRxSy6otVLqMHLKmm2BKlxk6FQqUFk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h/1qkWV/uZ0uLLT8ZDRBq0KQMz1ZCpHknpCYKq8gzXWB/dteRIdRQlA41yKf
ytOlTCdv4l5+RPSIZwEVu+du1+b4lEKzW9irySQKKQrJlqQBfn8ci6c8EUfe
9tYKbs8gAeZRkIM5kjde2I3XgVIcVrV5NhHsEJTuepgo2/ANevs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18160)
`pragma protect data_block
ik00xz3Og1Mk+mknyUsXn2oZrZ3JPlk9a2orzv/TLJWVBYarUFh+ktSfi/iU
WEsLFSTZwCc0fO2Xf5dMyXLjayJHqM6UVJ4Jwmpm6H7QLgExNFxVZMVRUWRw
mjfTAVOrIyBPCLUDve9E7b/anbPSjfqOBBYKYNOBbg4Sl5ip+6E8oGPKJXCM
LK9a83Whv9L/V4yk+BfstRWDU77qjnYA4NbsEb1DjQATd+tASB0FjfBslb8n
42PGVbojDgrkbcMy2SV/kUKTmTh5K2A1qknFni/agnokPxFUx4EHMmjJAlCu
El2XdvAfsElz6vSUoOwL9DdQPZUomFHSo0ALTKpYQz4KHos1L/7+1FTH0Vgb
4daJvd+YGEOcphI3yYMC3OpsrKlsz6tTiU4IDFNcQaXzUbRoo6TKK9+4TEOe
++RAwE4z/6HRL9cKBj8akvgdt+3D3DES9KUwCVzf2WAstcZWPPokw5vc6BdD
GtqsUSXRJQTrtEez4XCQRAbWaHKFhcuCihxwoN9cITUdWuivLfA/GlzkoSry
OIcQllmOFTJGsnVWJQ6ZUMoCj87C+fzCMweQtU4yOWokFaCRQ1IackN/Knri
Gw1+bkHbvnzpbe+xpFUjArP+KQcV/SXq3dyaRP3rfOBxrB4ppeR9x9HMJeMC
a975yJ8aAmAP40e3WE+JI6pirGDa1eFjPbf8W1vCzs7qJtbA5upnRdED6++E
mTxAa8g5GMSGwY0Hl50OWYJiQTcvt/19/Q3YguB/WSzsA7fX2bQY3hFlX4Kt
SoXP1uqc+k6T4b4uHqnyz3/yhZFfcVLAlxQVXqi+7MqaK3gl+DSm+UcBQXkH
RmFNWcN/Jj33fYb0JwQAmKoD7JBt52tLKcMKngITD7IvQfZOitNWc+CXBE1F
LPc9PpeRPdHUIEWZVIFs1XWtUoTHxuXKKrrf+jvccHbELDOdywqWBH4NyE1l
rn53XqtufjEe3Yz6cbtIbZkMVu2j3yIz93M1w1bNvb5fdwQxJbYt4sQRZ7Ap
SG6rFFuPgq8C01qGiKY1yqWEnoIYfgHvHrF9nK7cDYGvCOQWMS15elGwXIke
E0qjOHjM4qTPGmBYtwo/mfnG2ERiDJXryFzNj7h6yZxpGWvdU06LV6Bl/HeV
pAzd0p0aFQRH1FQMcqOWQvC6+TpF77JaVhDF90wIVJjGfTJAwoiD1VdCey+U
3PX3HBc4ha0Bdb17Lde8tTcxMd2xBMwwAbjTge3DhFcXE4gllCiorXO3NcUX
eYZ8nZ4dyzTBJD+6NVfZYwNPtKETVgblVKv0D6DwII+gZlOeoe8cbD9sJH9Y
Rlbdqbi02dNe/StnY7TwTWMjJ5q46/3JapZLpy3RygCOuV5BbCALq9Wd2sfB
b0uUiwJ79dbTJSwK0unFcBvrxCVJmb5qXGdebB1W1grwIEZY/VV0pR3qDHek
PaEGCExEi0Fzxk97GBsCP+/798D1gkQ9cjnF0Knuwb51xLtz4d5ng1kSQy6h
5tHUFRPM5edIWxJovX6GPdgwNVoS3z7ufimwQ8obY+RPaVZQNVCJKbApclSb
zU08Y1pZ6SacntGhLLUUAzV5YP/JvOQCOebznJaaqHcxO0Q5AJMLehqM+dj2
KqBRvDJhVXAFwy5bMcVoGBxaGJCz3al3wkxN626BrCeYrYaQEAkBnZrC7azO
k5pHZVmjSC1ANEK3lpUKlvCgW+U6a6bAW21lRSh5dSdbjF07F8xAYQTnkaGN
7/Zwt20R/9jvhSJ3pov/z4zvjuVGn2u4nI5qYlGOuHvn6yGbEDpAN2NnQU+Y
+oaxBshzvAZzScd+EIn/Y66EHNVSX0qs10R4FrRC9/IIps0Wt4oLePKvoTCm
hBWR2BSHFC9QFmqqZ0OYAC4R90lvkIBn2OVYQCEIQdoK5QUzug/KCPsjoqHG
QQT516QkzaI+NrFGmO27Ghf70NwVYjTEMI2hfjguOhz5GqIWhvE9LNoqFBQZ
1nbL/XNtx8jlQ82vEpOkXhbJBi5wtoJv999r95cRhdxt4EhUifYTt+e1gtvX
+MnEKm8r6Y6MOj53xqOb56gQORZwizwmjDWzQm4UOC2QVojSHUkvf3Ju41oa
u0LIsXxo5TErulapoZypjEcc3nRlfzzbcDExskEZM1EzJyU5dhmNxWT8PAo7
TYHx9ZhEUszA647IY6x6uje2SC40Zkew0IQG5muuHeLuLBtW1NTgqbGjNl6w
UWWv9s5/9YpaVDyXupBorZUdJ6OyJTgm+LI+l4GKGJeG888WmlbAvOO49rJb
rg+CGoCc1kkp8k/qK3wbQ9hrFCY6jXN0O6ZIRgrYQ0HQA/FHxRp4cdrX8/sj
mSOACtVLwToQzckYcK/wN8xNBYa67KlIP9dVkjyN2PiE3AEh5DcknfJTA7Yr
BNGmByuFQWNFHP+bCemjWRpCnRPmAUzmIk41vW8+ydBbtnRWwYvEUAVZhmeI
5qSFeB4e2kd6+ub7mqDLY1eWVuUCIoalzgwDjGGt1CUr/361i7CvmkZwzKwU
mQyNtYThkLnMjfugc66xKYB1F0MNnIoI5LxVrTviEUmrcy9MB4ClmVhbsh2Z
1IFRWDagJ27yy/Gfae+J8bFMZtC4j4LZvL7yWxUGLoc4pc9TUbpUIgiLb2k7
2rF37QlUJ2i9cBwe3z9A7crME4Q5UtjtDxDsEgqIawKoLBjTrsjWTbKbc5i0
44Pm4b50NeQ/0x6E2e6nuNCBvjtrV3tHsP/D7Txe4guREVxFYu78eh4Y/xWI
gjF2YsLXkD3WZE/WMOoImmFdQUfCTJd/70gcxybtrzaCdAQp6LsArt0+aDxX
xVjvI+j0hCEf/x4Qb1D3bb49MZdT1XMNIQgFEVHzDo1qTaFgQp/xhEH1dDW8
Soll/CWJpQDA0c6Y/I4J2h2BWztRtroSN02d5gtThfNosp4J0dpfeGr0pa//
pGUgX6mKNW0twaih+Gq5D80f9uSKG7OPs2hAZB/WSH/B3tFYgtAtAYK2QaiO
3xqCipFK5Km53a5U2+J/NVW4w+vk5TCPBt579sPXxkCg1TW/+r8wSXR6wPeW
aisi/1Iz0KRQvI1GHExZ9vCmU/ntoN0sKCBeEWxrM0B8D7Z30Hi0NhlAElSN
U/9F7JJtmbQ5lIrALHsLpt88Le/SwN29PLbdnoEd6zaqNxmqCemC/Lmt9Q90
SoDuEW/MUSBSNNGyjcOrmk8I+yT8GGFvM/qt7ieb2q/aEryp7oIzO87FRfuQ
GOW8sP5DXslQijLfELmBBNfR3btYf9EIa1Aw8qPe6JLTgDD0nIdRobToDD/o
RSUC+70R12yFfTaTBXrwSuuUFvshXMq/n6EWbHBDQlkxZ2+g9Jyknu6SEj1T
xG8lpNNgL+VIqa/tD8P+RV4NCXU3TeImxa547XhvBVDcJQRCm8njIvelhHiw
IAm6GLRFoFqGAErm/XfE29Z367+2QTFG9C8oPUyxgDpvVsvQD0uQkdzLLM+n
HPNQT8oRY/GU1mivg+hqWPIEpk05J+QdiLpSgvVLXteSg7XttCvMgOxGJZiE
T+DFVw/z4tPOLrwUB1kOXhBw5ctGlwz1IaMY9rXEEHH3s6y5M08I6INpzZAa
vXnoG6Wxg8fWD7raO6bg9UTtKvCJmZhap2dVJlfHTcGLIJCqlyWnrGAx7AA9
HQbAboeYMIn0Ms7jIP4FwiJj2J6SItXdyScUTGaKh/utMnZ3FercD+zSZzdy
HH1EIB9C7eRzFIXJ6Z2QXCFo+Jrsisx9bX72HinW6q6djU4to8TLR/wJddOS
UcBX9J7VS4QTeWhUMJaqUHTfIdc5hPK4uQ263DH5SWrl1F28gzwc5P/qYWEI
6qZ2h8F19GG8TwshB+aylcxCrTfCa2c653yRw4RhEWXcByDn4nFmsKcOtW4k
ZXuMfv6CyQdRedRiom36UbY2Vu1Cm/CE/SeksfaYg4uZoLUd5VuE2MBt7wBZ
xwx0JgVDdDAalN3Zy05R8R43cf8wnxiS6MLEQq8vLlaWjtfjPIuFUBsmWsOX
lbpozW2eIbnASOVjMCt3Qh4RDcX9Rbq8JJV9Ixs35+qTjLJvPbrda2RbA/jQ
mNRX7WQjaKjiMjk2dTdoC74tzNDVjq/WXC4B6bnHJy3e/OmozwiCOp/k1AQv
gGKMATeFVs0K6g7Bl2ujC/ddApJc9o2E8evSutDxyDotrau05XG1OCjc5E7p
wXlN2KUxWU7KuEc1hnTLPLGEoVeemjjc05NkVJQv1SFwW8j6psigwYzI8Pgg
m50sNP5TmYe8gRm+m4NhchVfuNRLFwfJ4zb7HoIKcSkwoI3tHn109ec6Adfq
puYV4orBjYPu8exNEAltY86MvW5F0R/jm/P6w2jQj3Eo7I4kVQmJfoMDYzQZ
p06BydEkZTRfG5zq8KhGUS+zSvI6eYbdRuQ1TNQDxLzKkFVXfGMMDKkotgp6
7W1zktDgS0SE0VpUXoV0+MPWw9YRx9uBMbKlo9+ApLQF6fJtjtxhDRnW+tpT
25kxl4DMetaun2ifHxtGHs614boclaNRTVKvC97mcB8X19WSrjaurtejJZGb
Ge3lwMyZBVQHdUizapLi+oMm22uq7+KLwiItodpyCdo1VZqXyWpOGiUWWcZu
PuC1fQlYNAVeMecZhjqMteFTZ47B6QWSClzDRALYWhc9rHeWdZFj5DcLAKv2
T6GwYG1X2PxEznYpu5IvM/w8YVNNByBElFaaKc9hmX2CtI1s6YMMMchdp4xQ
nCYlUF3aT8rJYMvSAw+KwFvnZEeElPeviqhITqTw+u6cKJcYsixqRpTPEya9
kb6UUKUfF0r6Zr7wvqrzhrxcTpJzllS6JSgru4z+PDW81YMyMh7L6IcYfJMV
yKM8Mm250ZVGP5rkvFRRRM0avlpOryEP0aQgaGGuSXSNMeGbgiCSMw58mBbP
Y+I9oiRXjQ3x+0apIrI6m9tQQW2ElGbLKq1kNMlNL46SRctL/Uynl2vvs0g+
htEXsOxWTkVoUTQ/Sh496oZebnvQm5b2LYn4biVvzQSft/f2Ar9+ZiFACSYi
zhRVhZeJCytKOQh8FhD5xQx1YG+xQ33dMF6IJqRVJSfAM8KBO5+vUb4HaTcu
d1EkREg+E+Mx5hGKYZH5vDfzMgKqPZGSq9IIjpOqEjExY1wpFe8ucNX8YFVq
Yo3IgOK8EOpAVK0dOVdcq/Eannd0jSMDUjRjzr/ParpQGg1+BvdRwnQ++lRj
e3m86OOmdltpmnY9BFDxG6Re4d99pewRgA8Dq+QtJpqXebMm+DUhGMesmRWy
8sTB+GonEGdqu8YPjcUjxGWD7MM8qwpL+G53dlAFNmJFJpf1TkFmg6LAv2sk
nLcaTuI3+u5CvY3WMIE49R3QgpoVJ+rPr3SZkl6Lx0o9bZvJqUBjqGX6L2T/
NX0DwZL7zDX1HVyr4zMwHWyd6eQQJQRd5xOw/lAEhZJEkQVB/UJRewYGIL/K
QoOtSjCZi3nmtlojaP8LWBPpQsOvb4rSIweEdO7GUjzNCTJi+zLCtTb2WRvg
o4QBEr/5JS+TcuRE9DRDX/zPwbtUPTfaW7fIAyvMeC1tXYER3lwYaFkIm3C/
1m8+p8JfdC+9Z0lCBN6TdHdHYpfX9FHDasW5OLLCNvhUnyTRHu56iS/xKu5w
rjOBQypmJKEtlhVwP+sfjh8ZF+e34FUNfMj+6CA5rnWQy4qrDNWw3zg26HpL
NZrSsTKE6JAw7d0h+MxR9K9/BZlRx3qiuPjSVKygtZPWMjJLkXwft8+jRyWg
krj93lHF0jgMrXmoGCDpU5qtNuk3anqGnxxGN5L1yn55gk5soGccNzF1GCku
TJtrRRl72GzkGtwZluzWL562N9+0lXXJrrWwYcjVWFCWg+0kJ/gm5BHjvjXM
io9yATXWRwLYUfa6JLkz89mS/Vxe5fYNzD4BmsmdTdnsKc7E0fUffZc6Y0uA
1scBNtj5HNZQFhwv+rgBc+Fucee8FD8la7U02/7MQqQ2izZZW4VBs3JgrEoS
lIXz9QF8QgljcX3zb1RHUdRi/Hh2OGKYdpjKz6zyCgsmgLMcbKUnhUQ8pyty
RDYlr91Q+rgBxpPLn3xfKxOPm2BY79S5tm83Q4lh/ql26kDGiXHLZ3wy6wYp
1j5tKHI/+rFMiUVwDK6WcOTJek7Z9/DPQ3GuZrma3WbXmSD/UL3V+Mpq7ZJJ
npbtACj0l6zUpqFgMnY5qcgMZryFqUzpo5n+X5O2HV4kzc/vVN7I5fdlfAWn
CIfIic5RHWEbaasFDVPbjReWIC4O/l7t7YLfNcFf0OJmHJ4PRaKmlMGlJjOx
rO+kPDtyavNbkjaIfp2voPReYEXu2RqinR6SY82dPpC/bIbV/IyDLngsjDeu
9oTTHPuM9Bcu+6stKX7zQn9+o1xJMXxJZpIYfM5I9hNt8F7GTJn1s4nWqDsw
r2ZgCZkdfMXey2u+V0oLXLXXWPM/ce1OJjwDIeDrtQMCBZV1Z3tBTejOMKcf
zRggmCc3tz8gyIrfeDogmGY7LhK7XG4E5vJ7Yg+atjR4GRBaz4mc5iNMhjzm
M0AKYfBqTC5+VSKSUafVi/n0dhk4ucVHEeo9ehLI0qL7Cb8QAgYGLDaQO/KI
aDTYMymyy8jEXHtf5W5urXzCOgIyofchDuucznC0ZekgRdlX4/+MmI+Hji3K
/osSOU+M40RnKpVuGHxhw6oyHGBu2QXmLeInFEuAF3OJzz0eOCZhJP3iUlVL
rFM7Q8oLerSrg8rxndFhiECSAJ3BE2QAF9xjKPq1+7tzrSOWw+qfKIhmiVQS
i6ISPhSH7QoqqxeQtJtQgMM07xx4t7EjsJTvVHh+Xq4QzC3DtzSRoEhRJchs
/qjTXA70SvIZy0oe/CBQflJX2WtQ6sAGAJ3jPdyL+hGzKmAJea6XEQKfiqtd
INKu1vhneqrMWDP1Z6ux3ZtDKHmLulx8sH3E8Vnq83FUZYoM/qzS+8qvEKNj
baSs7CKaZCN3XREj/HgsIRIvzVKo7DcYSp7JgU0OLxB+wdQSV3hXUMS5j4od
5q85zX8O259Y97ds7iXP7MtnoUJr3HcCYkGgnhJx2zV7azY4QfjdBVYXln4A
jlJM5E1mgdqTkmcFVqPICbJyPV06TDGoq0EMQLfy0NHVMjhdT4JfDoLbM9td
fHTQwsU+2SED73R4VCz2vE/72730oVTGb4FvUI57QqpMGfcTIaXVTeH0JA87
thmaNlsXvnCUwwJ5phE3ZgE8Ue676XJziHJOe/dGn7/BlMLO6suJ98qceSvI
AKlVcVoBahb7lMcC+PCpHbT7Abndu92IaD7ggaZ+dKRrF10I8PXleuCuUSLD
R1tHXJMCAuSwVV60wQZIvc5EHEtQqf1i06eNfQRYQNYMeZ4brMa9sUxCGclg
VWV087rhwxCMwn8bzhHlGBPCWI3iZwtGmhTrzJxxRbMwPqnPF9jmXEIDn0ou
7XXKN9kphGAbfGCnDFp1GEfXLdIA7sdyyI0GNf4butzLJINgbQOMSyT8m3ER
/MwsYitCUnGysNk2EAwrAKjvKOTVvm2vp4GZ8E01pifcLBNRRG4eIXJF9D5v
Kz9vqpr4pv/iFj8FImuDQTwJs6wqXNfDdDHyWc6/FReyHn55kIbi/S+u5p8Q
Kd3L1Lq629FWUqMflhIk0CtmRKJ1UxZfY6hj0hxyzE48T3rpJi4TOzMRamI/
J5qVqR+/dw6q52jmwcepHCQMARYM8Day8xUGFoew8uRiF8lnzjXORjyWLZVg
5EtvPlHwLkG6KiwPbHrW2n0EwYJR1Is7aM3C5LUs8OT/EOup8G+3c57XLwL5
AvD7H93ZakK/QuS9xfxaXi2ri6aV+YZLZh4BCYVP9e0ZrdOJCpPO25SPt/zc
JXR/8VthB57BP4WIpBTK0sWCjDwhdp6JnB5xkXhsBXIRmQ53Za2SiOUSvdDW
HzJsydHzdimFY9A6G/H2zQFx6YTk7i+F/GD6eFvFV58CWFKyVtQmkv9+wWsg
BeKB0TOrbhU+LjavZi/ddW0xaSzBcCQnlbfHO8lB7O9GnoCpKrZBFNN3rSnY
KNJcJKMsv8PdrnMqcOFKW7BeryMXip4KNuDySiSzR+TAM1RxQUZCnVW4AT5a
3TWQmRGUBsDy+BP6yxlWJQsx+SGCxuIPsmJN2Qh6n+br3nPQmqe6jtvqLvnk
Jnm6vn1noespwcbmIJ+AKe+6t4NJxUd6vHue59KAiE984bzbIQX0MDYik/GK
RNdkhr6YeC5uGjpKaWW5XAS+fpIEYBFzW2x0qrCVJMUjibZ1QCDE9/F6FzRa
ATdHXAmCmh2ERJLz0rJrkFtcXunz8LWKaQdQ8f16ptWBgSA0TR+nn9LjuYh5
+LjQ0sqAyxyP7xaKAh062nul/MU8+rTpDCajHwXSm1s/O2emqzELdijczZWb
1ofcBKOXY7hF0W+aresRpgAxpQoeUjMXCSdfI2vcNqaZ2OxwsUId0bsLVtMo
hhAm8dF1qP2OQMSWFnN7G5Nc3mEHbK60YCWYaX5FoO0oAITMrAa972Gv19rh
gGT5HnVQysqBoTsQxXmV9jl+loxZbLpz+jmCIG5jOsJUshR04UeiW7rvvwJ5
VwQ8itDkNc7MB7VzbYX2HN8v+Ft1xSrIGKEiU4JQpxzdyC7c+EndYJ6YXgu3
c9KiyDjVU+vSDzah9TjtrHIoMEPN6Pv1RDqAhRoexGtDQ6+UnjI9iygGmJ6R
33Li8BfRt/bhKdD/i7NKArApZPIldh5l49keYO0ygVOfphluxuqZ3qNm6VT5
HDjgs2u33Z9uj9NNkE2VXwuoZX2XpKK0tl0EGgJdY6mE8Avf9TCj0qgfaMOb
ytP8CQLjUHW9MKbyqdwEk2PaPBWG3GADoCW19JuIOqNQdFO/C42ZN97CAwCS
j0RDpWv/YmQ9djaCWlNI1SDrtaEHryYOHpY5iImY7tUOEJPa8uB35jpWRGfI
k8vdES9lDWe6npSnX3PSIrLldV7izlUWwHaDKqdWEDB4y8uJD1AxEimgGzvY
9Y8je0a6OOXBemrzPyJxfv2ZT3KGWDTThhhQzsahDOFeRCFR1PoGEHIQyCYP
GzlwSiAry+k4VxM6zp8j8frjWF7X993sTyDKRNNUT6Vt3mD2O6szlFa0niuu
F4bxHGXH71DfJA+S9uLl6xDGjqCnSXSotqQdgmHXul+XLhkGyfNHQ8AAXJJz
flY3NhPFVa8QI8WKiaKABN2myyGYPi5iTjZKyMZsrik07B/iD/Si0+6XI2xl
BvcFxobnRp0eP52iGXHbImY99k6z6lpKJQm0UFiEIcQ7tqnMdJiW++xhmug8
y/CCwrQdaA5QIfqUpP5sZrTRKOetGcQKj0ffFu3W+XgaEdTTSLvEg0/FJN5G
19dnNuONmmjpKQoJb0HakQswYNGPVLLkTLZJy4l5zkBM7nRZHzVbVH9SXldL
Ws79z2R1wCF6TvsZTgjzJhi1wWlv97Pl+23vsev0/Iwopd1cPM2cPELiti0q
ucE5ta6CWjsWkEEQz7/zXO1a0MaH/Y28GEMsXn4o9Ask7K5o+21YOMTf/3Si
riwIwQJtxoCqSrsEbWTxA5ZmopSF5o4aXdR4TeaMJmUltKrzJguvR+QblqaT
RjffxBtszdmlhnEQh1zR9DCMVflhbyXpL21cgX9/gJ28ALzCNrcKaqVAjd8f
X7sbGHhIS4Idj+/HeVPn2ryw7FF+I1T3AJoFcxeqbJBp0fiiz4m58kXT69c6
f/Bxhq1ALHxnjLkUg3xc8hqLjqwK7lZw8oaBHB+nYFpIAGAXHeX/ERwVYbWv
ajjnOlBg/oog7CBcKycAQp1fj/fpTXzbjB9YvzOXwC/45ntJBpcvx2TmbzIS
DVptbEBirvowQLNG3uNESp27RgK62hVEk/5ugRa1hzyWUNdSfPS84axA6CMJ
V99PpksoovyaIQA0r4qUQziws8VY39u9zPJnLpxvywdFH68IFz/CjlwfiniF
8oDtu8azl+pHJVMZpBu4Is2H26Oykey+2QGft7oRYVh0Fx+3ky0Ma9ofoxev
E3ytey6IoZkQHvL3sgnfnpvXAxt05cxFWP9KisO0l0kidNgNULL4N8a3RvK8
BI5GpflUv+/fOzr0t616IAA7jKTwOW0Jk5N1+GdJkUUS7XNUvfuoCcrTvdAm
zgp1aeYCCTVzcxh2ZuRvmH6p4YXbIWi5n4l+UCG4YK9SZ4IVVOd4RCG4BcaE
NmP10VBC+jGXjxuSuuMMJLyDi5CvmauwwNFsun79kqaU0Buv264YnrxGTNwG
PqsG2h2alsKU3Vr5TXiWXLUJtVyln/UnrAxe+iaVXZw1QgAw0f1Y8TgzU2tV
HuJdJiW69Qqan0f6BEtKQxLOPNao4b6fpvku3IohfiOm2WwPErgDG0Wx7vm8
/qCq7T81JTNvF6jsR/5lZD/+PI7GC0poWd48t8WZLWYnP9uL0EfU9cTkLvHf
MCGR0jMb3x2Gb6vKgqLPr3H0GKDEbwlZuNABijnJ88x00gIc+O5EFeyEeJuf
Aq3cw/03d/alip16ADggle/9y7L/+6a/78hjv292Fj5oDG6lEhwyhyTI5AhJ
d9YmjyXAQpDja3lEahPw+CoV4hgLsyMaTR381sjSufJaVfoixnXBFAoRZqYg
9TZRyTNxxmDBDM1ovPqwVZh8IDi5L0lUnbmPqJIysLGTEnE2KTBKOCp8e4U4
yxBWHAj574emWqwRKA7FC8aH+RNYymXY4oskq5RKPprB66GiwK35F/txWABS
UEs1QTeNAWwaEsk39Kz+9/j7k4sJ1VciEMfLn6AV11weCka9F0hN3T+Zry9o
zIR0CKW2onFij4dxewtBe2vZnj5Q/r8p5orWp1xsB2tgATaJB4LkKMvDIpDN
d09RslO+DCVxSKGtkPfEiULrB7xffAH3mfzEPG8GuDqzOyM0nbGOS6cCP/hg
gdyq4Bjw3jx84BPdH9fyRMXZD6aY7iQZyz3eR06qfGCvSW1QfcdUXfLhmAu8
8vFUhPK/VMc075Qu3rmcdofXVRnX4UcjEBeUde60PDVPNnRdk89LbK3eoUpk
dYplLXOx6qHKSHXBVD+217vVmkQHlBq+aczWusGn6+9ae4AWvBDtCvyVPTQk
m39VZ1vcKJvuHRdW0tIiZVKktAS61IhOjth5hbFfgP1miq2tF1VN9qXPipPo
z25FPV/3w6BbfgqqYGeapW/LwubBzAB72sqoxMAg47V6N+q2/mInVnfcgDIW
dQWw6TXyaoGLVF26UlYuIjMwDsPN0OhPLQd7sKs13t4JvUo/pyedjyJnuyXg
Lt8igUkobJ0tluItJyLDz2lSQ7wLU56ao4YCqKSbbd30a73Twflmz1LvwE+o
DxCT4sw7RO0KmVjYX3Nj6XJUstU99OJ1FCITQT854yq1l0BamodWs4UTeh5z
79nWDiI6D2uZnoyd+N+BePJyfc04G81qJZ0SVpoxD93wKiNprSyLjQERZp16
OR1XPXORY7KOQCTtIzKitc2MjEntcVr+UrMCtR2w4SSfI9Zbg8FImKv0xoTK
7ncF0OC2/oCMQLhDtIVzh5L5Q9/8OOUG/T8U0IE1xc1KFl/oPfWqtTkPzuyM
j4TJDgADqdJvhmUo8KcRHcwxZMWAhbKdQ6x/8Zk+0ThAYapq7qAghK28sJ0O
yHf55LYvq2/JUAaOv3ZUpeMxU/O8XouLTZguMKijV8WsGcCXzIfJfLj2/cK3
zl3fbueojHPQqWcoStwxl+crUAfm35oVlNP7eYZQS2Tw0DcFhS8b0JkED01P
/Q1Dhk9LgroqOTn9sZbZRTeaF587CPrSQi12/dsmBtSPZmXd9GNbLg61l5EO
WGuAQ4c+tBPakI7rOCxRDQp3wiJMm8+bWwC03vhNIS+KOPlVgbR+lx7tSqZV
q3FRIWY5kFmckONHil2kPZPgXc+syb4/1PHqORXFvp6ReDJUrL+UrVZb441l
d2TXNnJv4X4ikwVuaFXh35zLpCLATBn7lK4jtzJYlARC6ImMPWSJg6uZxlHb
i58FUiWUaW0TB+2kWjlHuCxDQe0m4AeFWPqmknDxcPcjf5Zirf+eixVWIvMB
y02ES/UbWOqyWJQPD9vcx7oS3O6W7BC2pd1n0past3mAN4P1Fs+8V6HREshh
ppKrijvOOnqgrH0gMFyiqeNX2EyinWqOj9DKHebtZtk4Llt94+o7gJ7HNO4Q
VS2SYy/5Z7ry2qzUilxlCmlj8xWDmS9EY4ASOdHbscjqJiIJM8A2thIV7RG/
cdFYPVEVWiXNvRBo1IRxwiD+KGeikQxflk0Q9b7u5qMXKlAVKMhrjoH5Gbv1
7ZnxpBj3iaq6tyVwpSOfSghQFAaO8yudypKAZW3b+UCZlU4L0o45Kqvimqha
Q1aYVdUrX2LLK9M4Q50+4/EoyNmK7PeMOCzBWVrDWlz10QBkgBaKEYVS1TX3
N0HjDJQ10pCvuaxzNmZkewtCE7WNTr//Av+4G0091YOY568K1olXhEJSWtjO
P8AUrrV7zhMxy7gRbFwQr6W+CxM8ZV7a/HP5AeN+uk4vsbsvQdyY94dY9oVX
RlefrLn7LeHgNaJF2HfOpFUfqltub45UllqkEQPyHOAKNQguy1ETLL0pG9V9
EHKV5f2eD34sNYN0p8jqzLAowvFyLVSrsLnl8q+P3IBlSDlwDmmmBDVwWboz
9NFgUfF7klZZfKKxOU700MiQwhHKR2wVH0T6y0KqNr/AQmkTd7Xs6UzFCX0+
f+yEl/5IcIltOeKbxQKx8ZnIcEU66AK/9RigsilXDa5Lak1xOVyaeE8NpnPC
/jeoY64uF3N1pBfuwh5oX9QWwnSpLYcsBWYTGcmhGvKTJmkhkbrJy8anXDOU
Bd6O8KTXGclEVbPiM9wtc42n1SkBvND/UNBvkSUkZuSJmYGzioS1ByPL+Fjk
rAzY9PFN6Np1ZK9Is1s2GHLo6M9iU0C2a5MiY3LcXAbuM4BZ5rwVYn7rUr8x
+NbdbqCg565It3zGEN6k1XTKoG+JJr9RFRiLLSdtvzbDdgBrGlgDmxd97uFG
dpOZeWlvr0A8J7rH3vS1P4Znq97TH59Qb+K8jMQvqVXrr4v+10mJpFSQIQCA
WFuH19ctbSghMNf31mk8HmUHQQTkn/K97Hq9YGThppbFiygT1W3X1BreBb5m
qIgLiuC3Dl4dzIATPjIY5+AG0tSeaBCxKwwQ1qcl6pYXhSXAiMY6vI0efh3G
g/FN0mk/+pgo2/W0idr53cg+jzeaCrtGu3z7OFlOfI7RynfQcJK+RboDJ4r2
rqX97oxMUnIexpg8zPKkxLlu8FHwB8mt2FRN7yrZGtnwpsT2LA5HVD9vldSV
OHCi/MeA84v26nF29IpRCbK7NFq+A7BGNlFJzSL1pGPm9J7BO+WPU0VQHXWR
Lpcmam3LCMscfuoK7chPlHsNRE2BTJ7OzONCTfm0i/sX2ajARlEsClvG0ld8
XLUnG3wqvDHRJzwleRyoLOxEcqKSSZABWID77qx/8jiMVNCCe+DNFFXsukHs
dNicaYX4xcWe5FBS/XXDU8fmt3UVPekkGHz2SDTtQkW8OyFnvTZ67Cs01sEi
PVyICZsJtI+dSJ+IFvRdt0ID6k8YCdV1FWEwus6qYHxL5o2RriSSgtbUoS86
ilv+rQN5yxV8pwUs7Mv+tAvVUJa2okfvwhsv7Pf0Do56qVtJ6L1NZQWBNnsB
RbQmFUgHKvYLTlrBDMA7kFcyoTfyk/e1HbThD8IpR6JbT7jrChStrQkTy4Oa
j2ZXNi6RrXz/kZNmcNkU2DycLTduQ3zoAxrVT1e8ty4UA2I1AxS9hSGJND2l
L9Et6RISJm/4XdZ+pAXiIxLdxJX1d8CNG8lRYdUUQ3hcwAvX1d5I7jWdc2f+
9GCrtziatdOR5ujwq/yPLO/3Ewe20j6EveYWjZzusvWEnMbxisShpc1YF3JE
tb5H+277/yM5xywSclEJ2Q/8hGHC1/vdWde5SdKTo6R/0dMauTzpWJiInVYK
Rsx7nMxL36946cxwLQomWikvPrbKDIidDntI+/90z3wTCCosgkRKpvHy5wCW
fYY2o4u1EKjbuVpAGQQcMqvO4o1siJaX+smx/gp6krPuPcyiNxlkc592AH/t
fWMHLJhy7zq/sY3j/qcEPpOrW3Weq+Vm9dkesDkbgdfj2OHMLq0QqvTxG85X
gyACd+OqPCRsYtuNIgmUJUAqJSdtfXH5t/DPh+lgfYTrYY9TxqGMF/q9yth1
qLaX/38T9xk09PaOPx/DQ+4sWkRJbLyHeSrpH/MI0Pt8rajjLR1f9793/COS
BG8sF2sGn8rEVRqEUgF6AySBD7ybo1yZDthPRvdIH9BNvbr2eXn6DBYjF192
deTEDkhGRTB96YR5LgR6INesoFs60a7EQDvg6LM5+7nH3yg8foz9T2qUDrKs
AlOrJwk62gwPCaWeyBx7FwpBaNn7ur6zxd7Ae2WSVO7VsU3rwJc+pH3+Hxua
Nt1k9BNQ5A1Z5Clk1Rz0+XpEaHa7rZu5ATHOOTc6ORy3anEYTcI0FKsq4BEz
o+D1PXIQZg9GrW8NSkRLWJ0zKYMnYyJczSEWRP1pSbMmsd3HcGkkiOTflxlw
tfv7DW66O+YSkNpxIXQiEAu2iKrfU2YLuxIRHCyhMhTY0/pBZV4pY1tOGrVD
eAnvmcIYD877/97J+PdY++SZnIkv+/PuQCMavR8ydvkrlbePNk97hKj/NaPj
NMqOnBnoDdXMsNCP1xkZMlZ0Ik/EBBKtK1SYZY9uG8zH5YsTSTa+hhOMOvMT
DNmLBpmjY6rhVKonega2MC1yzSdjc/O3HOCOvRP5vn+sTeCAwXtKMJtND96C
VoujnzZQLuZXxF0vGxZ2auZhl+VRlANLm5zODps0GLxRuVYzENUR2jJQ7DxM
8kmHSl5Hf8YXrVfU762kjm5ywHeXOzSxJvpozDiTYRnSYcsPm9YG9VV6HYvg
73udhDBKDXq84nqxrDtjnqwxreFmpKH5Qw0HPDX609uY900w830mm1pR7fg4
uFqUT0uGepOVs2Cj/FIHYIMEdk5Nx34B/g46lBgSvJ8UCZKPS6mDyN1TcJK9
45Ia2hDbixtwXQvZAiPhff6/KtOF3nTNXirr1CHQyQOFqSRgViJfJtfMFrlV
eeZJNUd9VTnEXvkrPOCR6undEa36cmEAHPz2NPeH+0NugqGzI/XBw3/r3WPP
lP4XMh6XsXMUx/6PHhvfpbasNFW5UJBqU2Vbmbbq1HNP43uIwr7qEbSQQPuh
FJTHZZLecBmnKSJL1jy0T4lEIlk5+PZOryBIj6yPkJTX9dc31CTIOtru8sXU
89RPYIboxvSlLCu/Fd2Nm8pRiBcywj+nTLLOr1Q+SsttCrVKs7JwuI+TnMAI
6rsJHLvDiNsYDgckwPhSczG3mlzS0zascCOfXQiQOWbt6C040kbDaH5RLBtE
x+YQNgYGP2wD68o99QYWCAc3rUlQ7bWFOWQcOEV2MgzIQiNQHHq+EBkg8x0c
Iaew4UGGqcat6G+EUgbNe6bV/L5MTpD0jbvGjzAeSB5awAbFoWft7JZ1yxur
TNXZjl0rY1Yp+mcIvag1TjwQdej3YsQoGhmgYOvummrWJSw68PpxmarUtadF
K1aQljhrJ+gCBOXYO2LcQFQgk7cXcX0RkZpxtx2ikLI30GidwvT9bbbSPRww
NOQXt9MmcqIuU/9M0Jzf9aIVmZsdhnceJDD+isQ7Ckox573QoQx5zdQFU/Hu
P0paXuV5t0eZB2GmeSg4vPvzYv/2/kOIWS3n0rqXycFvwSWXMcKCEEOu16Xd
V+ciIY6uuon+HJ0Mbl/O8zT/PR+bA6xzrqdjnC0e5MqhUgHOtHHm66+9DBK9
7LdqRZBicZr1B6DkMJsJVZvB7JbBZzMJyrWLtZOZwyeE5LVt0M4IutjAfeII
Ima9qE/7z8D7EDqy2xjSSm5jiEnqjbcp9eYgxLyyLpnN2SA4KzNS/Yk6w11Q
vNLzdOX8UWTAAhEhiWX4V+hgUSXtkEdWbPMCcVSPip5DhyC252mlRn/EdXO0
KblRLM/j7ZPwUgUzyvkCWzIUfRX3px52sS++41djXR0E4YM31lsVpqFk4f1C
dExKaLejgxhs6pv1llJSzFJuT+NL4xelY6W7mDydBlixGA4dNNmP1wvkgt3s
mV6/DhKz1s8rAuD7ZPh4zpyNJv2oBXoi4AsP3Q6rJl5S1bX243g1OCDRjEaY
IMzQFadGGWtCqEykrcxYb9GNdglxnY3blExbUy1dNR8kjQgJcHbuOi30blHV
BbqT1bnqbptUbT7UOIj9RAwiFJE298gbqXyN+nCAbwaYJYuc+Gc7iS+FGU5u
PU0+DHXtP2sxrFIH2hjXbAineOaiMPkWHnyqd/K8G6NqnyC/yvuji3S5pITM
JN+p4RG7XmTqbRrXekWF7w+3p2KaaUfsZzInGV8/Y9xfCFi9o3uhTGqIfXrg
ru+uwCa1fHUKFi+lwjCr2CtoS05E0IE4xOpUZ9tsfvmGDe2JZIoZQAOcWFbi
hkR3lA58gWxnLXmHI1yzBnF692VzIlBOHO3Zpn0rjkZS9XoiKNlz/b7TJKKN
szFOoE2eD2Kp4oBUkhl1RWpSPJg+hYONfX8gk+CIFbJeDY0rpdCHROeNCgfX
YS3eamRaSp996F1s4bcTbyHGP5OqbsfXhqKPcjoBhcKwtHsZLeXvCJ+4EkFc
JumZwKRQqTH92t3g563lgvUqbpS0C0bIy/jVDDjmE86LgTrYQpghehlvMR/P
ZOfvqvrKrZHgPnM6152W/d3cOtATNM2kEjg/DzB3Zf2KdZ4+sBCVBn/Tpk4x
j53j2jfXgd0D7BW/Z2elnhnzdC9XYcrgq04bvPDkArs+OcR0S8cRebSoex6Y
mjdNjWQ69AUOz7jA2PxA18ojq40B4GT+C9W7UjjDZf/z+jH1x9Fs35xbZHa1
t8A39p2/OAYpEgGHZdNaMwmZsDRxzzlV5xeojkpu2fgLtywLQz63lJt+DFHL
ovcogHY3Bd4Sq8LVyIz91CSs3b9KBcdy/hwhbkdGpAwxqDZ3liY11D/Lw7DY
SLnwKTIy5wm7/frzkbJB/bzN2e45bHa3mQvau3q5ln48R0yMRZpXJqY5awZt
o2Z+d6Q5dnmzltNxrOAuQWDbGIVw+ApGE2qVHPPDhjXM3AfuqsIFhCFLWKMs
qBs4cCQmVRevUCu7X7e2NxS130TXr8xWIucwxQ/gQqSvXcEntLyp1c04SMOJ
9fU/oydck1JO6QMICKzEpbAE5IW4iZLxcpc23X3aw9BdOrAs98DaBRZvalwW
FLqWq/gv6Qlz07vOqVAXPQ+uRN0YqpofzF8VQk1qIyB0dlhOtNqgxh8AJUwi
aq1uzzhzlXzEYJWHA46ArlykjFeM5xpY9AKte1VXt/3U4DieonCpExOpyOQx
nj3jSApwIcKFTBAjBwUK3Iea9p3abro/5T+fb5rLaAPwu50zYYS2VADKiQxF
Ut208xRZjr8Tm1vhcpOVD1nUg9ExymRJBQxv5xJ1lhAU7wpjyZkzlpaOWc77
6Yo4WwEFVBJznign2uueRuoWryjCAf+kL4RAX5uJkSUxwlhe5WSqTiM4HGjl
3dA3gvs7vV614DMroyosYAhz9kfLqWg73EAMWYL6tSUEU+UjWnaV4oAmTeh7
0Ekd8qSLEjSOFa6d3Eu8vWmsmH7pOwGjfgegtBi5V+XIEMxPp9HIr7B84UNo
RBoQsUQ3Vc5ruhU7jEg5j/f9FgyCAmVFdbDC/tLBLSX2TtMrMVOo2OlF+uHo
HBRyTF3ehSXOiw+01kxjqLnMUMgcu4ljQ3y6Ep04XH3Swky6olWhQPO/J7dl
zlCZjpYhdQCxYEWD39l+qm87ig665HU1wU8Zjv+bauM5drFYi7VSmRpR/ome
uNS0kT87nVMRNuHuhHnTwKapfoVWna/f0NJZmt2EguZs4HD3uBYH6vluZopC
21m8ZD5EXJYzc7RbYs9GlxO4GBL+SJgxNeDX1l03RGdR6WWffx6qK9tnpRSL
cukjItpQbYdg1pGNL9bY/gYumI6M77KESK4yBklHnZ/Uo5FjYysqzuKfGF4P
Dngw55kqmqKEsm0FaXf24N6dxSEiZWNgKG7Tsm3t6zZi0RV1kI/deTLQXNM6
hiOGqRRtmlBiY303JV0FZMfQ0JgMSa1bqdJtfw2v0UsNkjC5vTp3TvNH7tZo
tRniK2i/htaicxUSeyvaXm/GOD5qR4ZYQe9oC2JXIiE0oiSPZzccxZPnp781
JJT3ZSR7uIa6eVRhuSk1eRiW0KmVfLR7rRg8nx69xt4it1Y7DD0S1EMT5ZOD
SWni5PB90jKKqYNEYgxPjYKYx2939OSH2uEBwV3E7cRP83INqzIdrywbI0c2
2qAlthwwVKbmMyJleCJNhbEvl2DALCH5mFmU8uUlIVkg+8oWrhZmjN4WyVlD
2rfTqH82eo9lPneIsVmUUIl9Piv7nBx1qAPxN9f58BFI2j0xoQNMYDWEl4Py
UPp6cltkvib5wJNRGSftXgfQ4F9dVrxrCakBpqW3GAl8EElSy4y4FNuUU8sR
T/S40HBneBy9X/c2SNaqx6slx5+RNUpGA/GuleydUm4XL4IKSW/078MjoItH
wnM5G8+c7hRNgLHmi0xnJhIeLt0qI4qcfvIzlkA07QWv1KCQ/ZaFaKnxREE9
FZy9NYXsO85sRlMwjLvpGUH5uiAs2yiyZ4c1mIFZ5BDvA57SfIZfNbJzC4Dj
0BRnMOmWGZ5T2g8htdkmzGL6RgKAvdSRR6Rhrh4kh3LILqncfR7CHXfLkH+u
JFJbC+2Rblh4Pz5abV9fdB7NGGxlCKl5Rw3yx8GDK9R4LowhKvUL/UTA06LS
OEszVv0ikFwauQuMUoTXvhFwm6pzann2NKiQSplNHPgE1jyLmTR5OUaS4Azs
LcOvXa0Me+uCMq53Uu4Seyc8g1KULwF2LLFmRDJLf2rejCvJvj9xJOP1TSmK
MqGnUPktV9tnsGFxt5vavDckAzcX25C9UWa/nF6tO33QrS1ABUZmvhmsVHHn
1XUzSJgEDk1KXy+wSArAvfZ1ZBcaxijVqXOTI4AdNr7IL7rMdjVBiv9EXDI4
6x+k9SoO4ywuofZBeMK5On0lGplj6HxEXFJSSG+6QgzPVmKF5CU5IcV+WWaL
oNaqyobMnj/lZY55q73BsOuSkemgt3/LsUeacaTi4K+hpdj649Qc4w544YRF
HmgZgkKJpi08CSD+AUG/u67GRBvAvnoe2joTwaIpJCHbv53s3t5MIVqpz1OD
+NklgnyCoe8IeZFlrezNZHkTlom+3hnRNlLDFAcWGJonNqq5vX9rJOqWN2V2
873r2AlWGPLYjZa6RWO85ErfEPDzEF9qOi3hUSDfu0GRUwl2I9rdrVye8hN3
uWv1Jun3fxC8oufavCl5v8qlJ8wHrJO5pDy7mbkJ3oW2oisKFmp78W3KHVIC
jiQwKKkN6K1aeVHndlu7p/YVkpWe6b/Kxeq1YaW80+PIdCK9K7rHrGXvmBrc
QyBAoVajNrT5bWNvrdgchuNAMvBkrUh0caWGZ2HxurANQV/+TGgqWim6LWBW
FyTaP2g/gd4Dzy3t3Ad0nH0rY5MWiPqIuJsfT5+fnKuoyANuhsH3x0s3+kCV
jrbBoWau5UxNd2ExnNk1N3RT+bn5hoQyl1eq9Z+oTa3eR1xJMBNgF0g3eKni
/AYcpEnodOJrrqNQcTpavqx3Y+zbcbqKzvA1ux69sV/pu06CMibPXNkWGEHN
4NOc8iYUu8XEV/tZfbndFAmb6PUnolfdhhu/T8MUC3tSbQKkG7vIBokXlN72
vBytTOXTOhq7VMPhq/BOmE5sVyozCmcR4XAYFF2pumeuBlnFOmM4jcDaUxYH
fzP/wEqZBPbleOqOD0vWuTkGHC6PS3ck6KUPUqtZlxUwZbU5r2DwaWrnSAJI
kwoL1RAl//dlAc1+0Uj3bMOB67jjXBaYVcVBvPkKS+l9TahaeB5rHgoG+dTQ
lMrCN6VAfr4W6pA/BAIUBouWSPD8cN2XckVPtTXElo9vM1v9LiOgVdJVDCNZ
msXOKVuDnsk1aTa6+IQFlcKDwug3+e+07dWXUNNWwlo2IxZK6mB5qbwRZ23K
GdwJLq5rEFlXg+z2u6W6Z9Q7q8aloFLove5pgN7YXTEIlpr2k9tUIF+4BR0U
ZxXkIlazARcRUo1hM66hudCSbmdv5rqqorYi0aURjYkTpb8JNorKwJcLNEtb
1urvXIfCvy8F9doFT2YofuNHy9UzYP+gweYEKLfso/J1pmmnRll2IYgYZM7f
m85efkq9L0VUB6ENisJHeUmZk4FTuJenE5porG9GLhdcsoJCaG0irkumxOyV
UPtyPcxKW+6kcTqgzBYxejVyAcPv6SxIGwXD+EBhu+4sv7ebqpTLPHogdVek
UH7FYABoPvpYUi2bK9nXvHsnzL0LTsTgfysShVYNXbxUjKzhEoDG+RPOEJBq
kpDWNkmRUHQMeRKxfSa/bH2JEoApORsPWpB35XzD1QRbrGhGrjG8wWrGM5YR
pgVsVtRroZoZnm0anHL9WLX4JKdrWom9I5JWCkRc3nMUE9qZ/k7gVoR8rZcx
+JwoGHPYg+AU7ypyKnkISUJ/UNA5Umvu9M61ubbQdblltHW72C5kaHbovu92
DVAIR9UIEAMpasme5zkqACAZfBE65f+dPNnF8jnhipg1J+zWuCNKh+7T+uAq
x8NqiX0QDVbyY1htvj5gdfuAOyznOOCWY1FtMNp1THpY6dRlyocFWzBQJ/SE
vsMKlvhi+fsl/OuKbOCHR1yc54xCOiq+uoXwnMu1ucQI/xKrsfQ2T06uOzD1
a96Rrgw9dqbzAlTeitCF7IcYH1flQDOpfeSSNWDbrygBLsEu+VjLCpZNU9so
IPUFKkGCyjnts0fdtQxzljqbv7GzcL97uKL2iRwOOmI6+z4/lJszc2212pva
/4G2UzGuQ9B/eYXJjog+rblgMKazbZRGq9WgBlFRThATviKdkLi8n/kdmN4t
Q9dRtpT639bTQFkRWucJ4+l97A/tFXlCBzKMhQhHy4EJy4AQbpqEpNDVW1k4
T0fXpwuCgCNKLr2XDQan3K1Vx97iYmwYT7BWe2Zz6RtFm786SuE8GBCH1lfv
2bN1OIIDQ2O0ulR4x4nEYbNoWzN5zWCVcUbyw/x3Zn3dTx879vpOI95SBWWq
hblQ4ugDen7GmFU/N8f8PS4GG50BtukRO2MsGNvViXI5OcZsUH+0o7GX/aRK
g3LrbPQ1ZIqVyc/kDiiizy1RyLEAiXJKFOZuT4caUVilbcshCE0bKWa/7yyj
LMmkRj4gr9vOWl0eHavTJYwWOyeMuylczK/4UqUW5BcnyNMXzlEQsZsmp/aA
TgnR719M2APySzMcWEK2HnJ7NISAgv78Ux1dFp4KLIiyJ0SSrO9AL/OA91OL
Yihe38P86gfE/Y8osFqsqcVbl58h3pbdXelJ8W3g4Y/kyIxzZlJADtGiy9h2
xDrhxdcQcNEwLMroAOdhGYkLxzKX0VKpVhERob69xim+fVdDLQfjkmi7CH6l
MErXnJhUNhhgzw2SmxKb993hp/a+YiBF6ccoVWhtkku/Ue5yR+HcuOJVkrLw
d7Ygzkda+Ag2fjCk/UNbpjzjPgeFjry1WXlhi5AtyxLFXTXcjdBuXd2yJUCU
F2uzu+/4RNVcfQojUt4t5EfBLQPhmyuj5ueRxxox2KvhnA2oGRKf3cWQrMd/
YYM74uhIffcOntVv5bkuSx6Q/km7TrJ5MF4sHUvlb1GZlVlU20ZvwwUTsJgN
pxViO4AF+2K+ZLQI//BTFBVGF+rBGi9/3J1oXQfaErR4MjrxdOmspO/53b0V
PVtB75wf1YGUub+EREn5BLuIXeLXqcuQpV/5s18eVeDC8ReTJAc9ZJTgrF/N
a97WP0X34uhitT4PF/8OFjRcM2BeVadKlvlFzczSzBbBVwC91yrt7pJvBkO1
X4aOJaqWQksXhTDfbRs6PZGJv+FGBhzXqBOGtpcXpIZRNH0iLirncG0P4SAM
D29OX5TmOSVc9vJeveiXZyW34TYuLkqixFci38N/P6zj6mAlGBaoV/GDYNgL
d/nm2vorii53MxyqfT434BI5zGphOt+xvDJnZHeuSINkb8vE756rmCI2FfD7
GjBFG1IzdqJNkxUpyXwT6jCdelrHYiL1RNgm7vXs4kZheLInQQ63kBoFN1Bm
ZI5Xgz6d4hF6K5pb2mXl+OQe52XeSC7OJHtGw0BOTYXNqd4ak2VX2ScnON56
GdaSY234eWfbAVI9FJVygZFLWjTobtpNp70tM7zaxvXxv+Fdag/+lNG4ol/1
zWUimx/9qRf80bHmSrxkQgXdk35zIHCjxUJnHY089TJ3HFEE/fCZ1xFMnben
i3X8Ml3YnEzgedObJbjgbR+dafA7w+2PxIBkQMlBygFqh5KqlGeLCVOpxSxq
RM6wSgS08GU4ZagYK9S1aT5sHJFrDSw8TxCXhszAQVx701EZDo3jEUeTUNix
7zHmZkJmw7L6G4leqQ7mdKLd8b1+T43rJoazcrzXXCcO+1zzcmBUS3/UFRYX
dj0nPZUPIdPqdpZVLaP6p83/GXRlNWdTufPHIcbamf9DMuHbF0RxyYlk+ZHk
yUoBMgzJBOAb+4dbbTDFb0b4sMgspN7CLoM1xMBOoHWa7SFNw5dUSRWUr2hQ
E7R8wkvN6AY0Rpjka6ac2WfZQ2OLIdtzEx7J2iHCt2JLnnHl45jWuZBGS6V8
mVOGURqgULo3hkTTCZZ9vTKtQKiE207MeOx4kjVRqV9ZELj0J5Q8RECy7tOi
rcX182Elcc11dnQzW+qAvJrdjIk13p6RKUI7E9bF/jif+PKjfxxdIx3fope6
LB5fdBh0p391DkOoj2vChuU7zWITBWQLcVb599+4LX3LGFwL670EEH9YagsP
MM2hI+IDrVOhiVBU42dDL9ncdr/4mpiIp2yL+SYa5vbHvH2UEbRut4MbxYV8
FLxV5FKauu+7LHKZ1JTVzGwCY8WuMgqSgKUohEO5IY8T2Ki5jU+lQqx//R1C
ZrR40A8tB7uqHQcp08uwPtxHxuBvk+x81koaLWw72boHDYiBr4M7UYLmEdN7
z5H1gKs/DQ1Ds7Gs4wxsHgdpnjoFAhYXWwHYEj9BFT3W9bUUvoFlZf7Zsjwv
HMQ6bbHZzkfU6hAkruNfZqo0GS7Awnxg4c4QZgYZVmLQKzLd77Wqz6L4Bj0t
pQD9zzr7tkxTmTvnDHiiQJkXxrBBJeFN/Yq9e+88Y3RjWHD4p3H4bKx0vWdo
3Xx7y0YFR30zviUTMDgMhmb2mXM7kfb1eAjzKO2hfVsEcQLTHL/Vr70kRx9u
/Q8DJAg15Q8cWSiHax2P+fgS7DQkVer7UbCwX8jM4JzOJNzDh5pclznqA+Wp
ifx7NmJDKqcU0DPxS6k5IDvl6Fo4eW30gv4FiBt6pZQNgBilbM4D93lt5Hau
RiKOt63GH68YOzyN7t82JaKZlT9FfkFUzeVq+nlFRIyABS2OblGfyWyZdIJl
2Exv89//xqTw1jFtVVKKPx2ikGLsxZw/nDLbtDonQZzDAba5XGFr/t2dLdjB
CnBoebqRpRTNMuKZuhCGkhcAq1UbfCy31NUzEvxpmqsGONQ0BSbPsf6p2DcL
PlMKmnxsmzEYY0fapaynjKIzA5pRfOPW8h+kBqh8aLXBfu1aEivqFeLVEc05
aGehcXyW+M2ty6d2gqe5HZc9LU+7Q+tLjH5uPRvVoww9813h/kQTf0gB2D3K
nfPip84ll/EflZ7ofV4UnkU1h5SU9IoZK332XVAjy/VVM4EKPjiu7SZmA6LO
ThTucWdixcO7ad+WAzdsPYDdTSz30S4QqxKTXjDOJIRAvkX1U3Doud1tCFMx
dP7CyzHRrDV6yXNlc+LxpEH/gQvJHnlelz79N6SbOARV28dhRZGHNINCtady
qvdXT+x/86olu/Nk6JgcFuhZeRWMRp+rySzT7JIW3sh98pIlxbHrjuE/pfVf
O1FTeMjdwDriZkq9/wRlVXuppoqlFQIRVOOKhIDxF/SlbZ+ZJYHBwY2CIloh
MXinStowic4KjootvLDh3nG11IZitbijTcjRHuHVnTtw9MD4fLa81muapH9q
CftAs00hyhotFI9D/8Sq+LelL/sUiTplVRqSyzvLV1Qq9NodjdCQLuM8smfa
wNK9cm4I25RIso0KbKQAmi+C3m9FB31GwA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1LjduoO7cbfF0CcOukG4WcG8bW7tMEKppEgbkqI12jyMsL/tnxtZTizg9/KeNcv1eG+cHWNvzCbn9B7ONmm+fKKP/fFDyWXNyYAViu5nO8uJTQlfD/ybo3hsPN96mRWAqtIckZ9v5L8QUaExoKxYX5741c4PZMsmItG5s1B8eYYV2lLBkYs9Cz24oyMyz7hULn1IvazyEO6E2l0K4N3x/4S87iUU1tNgbQf5rZngBeRFMDW0IcC52HsKFgTKB6zAhmcGpBJFhOFmfuiLwu2sai2DhIgY2QZHED6euTdNbNCbhdBaGDXSMlH1NdGKKKoBJmtI5jKzJo/i0jYalDMw5QsrdlLx+0ofcHZKK1U7sprsu+VuDofCsAKBj0ArLKoh1P/eJ3XeTiCFq3zKmx6PKp3ThYjl8weDl41o41VvNyioCoinvSMxvYQAXj/4cUC4Rc2Y8xQ0gTIKovWKBPRNKa86EC1/UnyumeBpa5lLnYrYFsD7SQC9KibsaxVDpKPqV+kmQHulUG2aPFU/9GXwCHLLkvFq2qDuKn51+LR1T7ecRIfEIaRpnVu0ogIYKXJ7sdtAtr3StEtdz5bf4NrcTAecwGcN+nOvUQEMnxUITDb59A7n5KqBA6qeStOLUxRAUbulqPj1lZ/xGdJqk6OnQ/8I+IwfXvvD5tdAdaV7D5oZ6EFBrbBqoD4TE6J0FhQ/4i4LWKAPdumh3fHAowI85oCj1nA5g/xSC7pMudt6MymIw7abcSJcOd8D7y52H8wB/WiSOpMPj21t1qc3FQbU6pu"
`endif