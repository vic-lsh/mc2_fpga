// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zohHYAU+f6Bmwp3tXmtzk2oBsTzwCsPnm7pbS8UIaA2yEQmTgfRmeZuIA1Wb
7mdUxUUp7fydy8IHN9z2pKVlTInwfhodJohyp5KZvixWHVXpIyYFJyOLZefm
2zxETM3Z/SBk4M5rj8U24sA8jKWJDT2aVl+U7s0u5Gv+RgvhDdLA3SdOaip/
WT+Cg+62RxfClSTUIJZZqqNhnn3wNtb+gcmBQYHXdAMpZiXeUelzwRZ7K8fU
cgmoDYBvk0sn+QmiL48tzTusHgIDx578c0OAU37wmdpmHPQtzUjFImucy96/
Kl1V6NAw6mhjf8jACwa2jwc81EgBWglMQ8nlzdCKdg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fhrD6X0dYkcLO1Ev5ISrbEu91uDl1U/xFNBNu5M9j1F7A6+lely+F628AuZc
8pJ6rcONDxQlUHajzVmo2HsH9OCwMcTl9/OQW+hA9BwjSk6jbYYHxR4/5C2j
Ia5WJGxi6tJPezDezOFuZfuYdWo2aFW3nHbfQLw1qhTjMqReFw6PSiD6A1ji
O+YA9gZtB/EVOHFZNqszG+C3fXZVr8HJZuwMtFTO2BET8w1BOJGELjlXIwl4
lx/Z6UQcRA9q5i5ErMkyQXNzrloj1CNGO1xA0SRCeFsd2O2A0rQwOHGhDQrs
6KijVBY/ie49Gw8sbI4mkVGuulFKMnWEBDyoSWBPxw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q16+bK+nW39JQz8+rF62b42CeSRQw2n/eBUKjJ26qrfjwEgOQCe4cLlqm1ea
/dUSAW+QY+eiAKc+J4Fi6KYvF2Jr4baqnjcFGgBsjDW6rHLyTJBRqpJvidXw
vPA/yzIod7UI5LJdBKwW3qBseAfbme8VRvFDZt+gvR5Fq1Dq4qY1bY4+icBb
DTGqlO6dXOV80DheKMG5Bm7T+hasXLB2eevNUhkSrWkrJIaTBj5xsVIaFuAy
MZ7aQ9J94yDg1fQZ2xUhqDP52hg+dQaqqGK6ScYmq80m1PMH6fcltRWnWyAk
rqNy0WIYcEIYi2h1ek1q7ebVpcsOxYO9nToRI+tR6A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mEZhL6q99TfsiA+Et1PXIsrxYuwXLqfwV5zv27jfcC+vf/ma+t6/tp2oC2Dd
5sltKPWttarLHJXHcsRXsbOO3ud4PgkZQE9x5vVitNFhjtC4eBqT0hvdAFti
0d3otWbI3JdEsjgtyvNli/Ufxjl7PO4fjxLIAeQa1GdnXt4KxZwpMs0o/DEa
9bOLVTZkTsQpnnuZri/tj0NiYBT+sxsLzA+Ng7Ett2HiP2i8bAVp2RAddSw0
uBOcoPFxk62K3TasujHgUVo69ZOhC21Z6q8s9TUf9OtYPgaiVzYMoLE85zRX
Y7RgL+07FKacIparmC42CbcuwpOgZXeYep3OHUA+Kg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fHfihRBVicy/8qPpkdJOlW0ZSNUbHUoxs/x8Bg+nW9WzaqxCPZ+xMBr9hmJo
KC/7bN+5ycXCcDPp7R7W8loQAerB+/2BAnkXIfPBKQx87ADPWWTS3hpQxcuL
RvkvWSNdSshy/eElAz3q7EpmvemnD33inkqoBFEmXLt1FwydLH4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Pb0gzSq8PeR+4BoDpHYp16IYJrJsrFgtauSNBX/CZSKne1fT4Huapco83HCS
ZLTAuolAASo1drKcXFKrl+gSllWfjt4cOZgrjuA+1ChVNwnAI8eZPVkZFECo
f9lMVvzcuiTb6SPFRoohnOV44S6KFiu4lQgtAnYKVNHWMdTnI/l4gKpteklT
W+VPh/sfYfxwzWBVIi9uFQfDUKcMM8JCb97gpYbGGDG20eEmsA9eFYPkzOoH
SI4fiwrO6aA5tTMJZSCvng9XTVlUZx09uZYMzc2VkBF6JjKfK/+ZbyRfgO6z
pbP6kVX1ZGPtHJsgNmeS89cZXBR7VCRomkKo6WCbKZDIPI4G/4IOM1gkgHfG
igdz1jt8MBWLCgYookygvCFDroIIR++owJYyBpXYp2N3l4lITSMxl4GPJ8YM
hz6jUVdJOQjDUtJkr9kuLy4ijch9WsHjA7iM6P1Wpy+4bO9kFLc/h444JUSh
MQ0NunWRKqGPemHvS8MXJ5GCn5fSqoWl


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
X2VBa/fLvCghY7EuEsWeafN+ONbsUrnrwlLv/MpeXXCes67QinIS6oB1Qu9G
v926eWeMrJlmuT740sIM/jnTp5AXk4s+2IWP1BwXCOWCl2bZFCAWK6dBaXEe
XrW/0CZlj+Gspjf4NIITZVDHTG2sw5cHbaO0QihkWAnqmMfRWA4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dmyoD110IfbjM+x2lmViNsrQib4LwaVEVsJb5xD4wcZpk/bNaUkSBLXL3BTU
hx5paTKkcJmmJsOwz/OngJKUDGZxRKCio+CnkpCS8QNq9KaOWEEPH56WY/f6
1EIRCF2z5BVCvTYIwCAvqpGkr1+J/ZgMk+VkI0IOokctV49DvcI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10448)
`pragma protect data_block
cs9eJpeVrCVLs/wqRcsryZdOjd8VNO4dsrEurrWoVATU99TzmIveFrTpLjZj
TcFdGMn9wRwpbSh0oXn4bmiSX6qO9LkfxQE6V9lmSL9ZSIj0V6Pu/1eOF2Os
YiguiwWD+DlqX0OfmF6lnq1uClBfmyrB3OBDPqZ7pH7JW08A+0/axnrYjTV/
zosmWT9Y2FM+wMUtm9aMhT/YeNShZV+nQ2/4uT36d6h6YcxJgn1IMWQSwlsj
FZOuTlJwb7RKRtsVzKeCRFBu9MmEIBSVCG/EJyCmoZupHFuaDU3Ny2vW9fpJ
9C75YQV69NTASQFY7T7cS/yPGNEw9vBgjm6i3FgzazxDgqL0tJyDREDXA5V6
Ud29eta7/UD1hEY158qekAvyBXolOLtF6h7ejmhoS69ywRmJKc/NEPp1DBHH
eBS1Hd5ME8xahBr1l0ujCJae/2Lz1j13TbPSAOhoYWAHC4avCIgmvryxdl/4
Mx8Ygahfa3C9jONlWYfgIetrIFCeqyO3ekWYuDz/bqj09mcx+I8/oqLOs9LO
ZQ0L19TGhhLio9YcJdDO8wPQDEYFddiyXGP5chXVv2ICpc7AHGkRIHZxdzIo
ZHcjfjWhCbGxxCZe5AEZJtWWOeewL0VIHRWnTKxQDnhdOCSz5beryO6Op9Th
Vfi44o3UBCuZwDBKlWpokHnu4AsQXfkWRjc4MO6IuinW6MPRekbbuXHTyujj
nsIh2pR/CPEKdbZ6lQ9R/NrcFtOXpcnPMHFD7tGRJ068PFzsk4eH1cSXgfGX
Z85hdImnQV5rfrTg8zfmwY4IzWX6o4zjSWh8yKqMQRweKDkLiQsj3LjOZI+n
Yg0FKB9HdLrmZ3DLC9UEfBCHKRuSdVdJclA9DKGYR2lN8n52TuKcM9rsxGoL
F6ug0UiAjHpu1dxvoN7XxrWa764b00pwML9FUHrYEJrEQ5cv7LwAVFEv4K9b
UN6MEcncci6gKuaJ9oTTjbX+VKsqNAKAaxF+ajJg14xTFDgaEk9RH8ZOMR1R
00VakMhMdvD43C28EY/BIfOkfLfKXZKcwlkxQHJV4zsSkfuJn6dFVOpcinCg
gSqZmOVbIu6cDJu7lT69r1NJ2ntmyNRSG0uTQHArTNfcMHtMfBNqUfOcltFF
WSZe7D3ppKWc5D4jB3Q+D0qoSDxDCE7wxuoFbJqTxqIkmOQc4fPKzIQlmfOJ
w7elSmFjCHR+V/P9KckKGd5+vZfsnPp/KlFt+0VxvbeP2te985E4rdYtkqyd
i7IvG1cwNaTtEcnT7tKWom4yzBiIbEdnqus+TerwArYN257L+uwy5D/KhJLU
90P4F4t8GPVFBlG2TB3RawlxwcsENzUOW83+umwte3FIBehfKCZ1GieY+kJg
NGmMG6eO6BPCisgkgKaQaAM9++Yf+KGccjU45eqHcsHVa/EksywJhSXRXl8U
hji+JkEn+E+KlXvGPpkm7Y26euT0HWvHG1FEQ4hzhSBDwfi/SCgFloX1R3k0
70GwWh+kOVVUeCd5Q/4CD7aAqYW20/BwNvXX6Frwm/O8B9JE8FDbOfhRCxAv
jJEpBYAVWUiIxOi7BFjllW/bDFYXwdZu5dYCzRQl4bXjFQN9R53xf2H+cgLp
l4rf3ZiU58eem+z5+a54/5By1JPp2ypPVHY+JSaE8mhcPrsc8I17nY4719EI
AR1KcHdIBQMxrrnDRLWjwtTSc8TbhMx0ol2BKkSYCyYJMX5gbi8WADxu1Frm
tNMl0DaSkhyPb6lUnsk0Qq55/ct5BiesZVMQvVn5ha67MchZI7a6lMfzUmb0
GM+pX5Df5ZOESBc23CCkrxnePGRNFk9KE52tg4bI9FkTbBSlUU1Y0rf8U8Qa
7Z+7i48bK6qlvgfka/3SRsMWqDIisvuBmc197cowX5bPLUz2c1+H6U3MiFyz
s3k+PYwFr+DtY6jOjnKWW5b5FU+ybAOj2Y6C4fQBcvGU9bnOqmuohYgohbol
9uLhqQKLv3VfXt+VMcohDE9PSuPPliAJzoTcWZLRO7ewOE/BHEmE1iSxtJwt
5Omr/0+0dOG12m92Luih3bV1BjlA4tV7xzohhfoHYVxj1MHmhUE/NIhth2k+
85ORvXb96hLIyVqLgtr3F7VqigDzF5ToPGN33WeJoTZUEEyRxdZr9uRvucMP
e/El0ZuyqHbmbwYhvgPYLmo62tB1jmfdoiU4xEPamVIo2/vC3O5VOyIJp83o
Y+ANIEMZ7EDBpUvzu0ay4u8IyY1vkPf68phSclBc5cYnOtqzU2+QDSaSDDUH
0oIERaDWzxSdaeK8U7m2O7xri83oZqGfkUE9xGDqZvAFNShreVoNfiB+ZrB0
AGavi+botlBXoySvjiSOBbvspsQ880gNa4hY2HuHnnkjc7PRDy+ewWNIMZxq
Z3mh6azUH/bh2aXaw03yiw/SLgDPo+4TLypkmfwk0OUal4MSC9JYbaBdelzW
gYglSwK7AFmdA8nrqJ3Kuvf/exQgDQuHWFfyNXXdRCVqghr7eTh2fq6mLBMv
fti4D1NPmSuryxwL2cnTq6InG0V7v42dq8vxfbjblqMh4K5QHCMclCa7rJee
lxFeuIuupjynuqe73YYVdnLS1kPk47m1mFiVVvDEsX9CQdUxizx0EY4Dn1QR
8ynRIvb8QF20Va8ICqc4iYxJbqSJu1N5y8qAFPVUiPuTEkXHjQz0Hh9xhR/H
A2d4Q96XDFQcwt/38BgTUvAAymJeOXFenIoOhoW9HCjbEygM5rjzmQvBHojU
KfXXzwrWPbZy5ahkGtm6Yx/Mh0GPuNb4yJatgyscqTIZ5GHZtd7okS7bKr/1
14s0X909rOfyTRkassnQgvv7GpOwklHmOrGLpuhlQr8kHcPiDXna+OZKMzN+
5WCQFKsyg+l/o+6Nd2tEBelpbu2fmU/PoU+R/nxbWA9MnkdlTIROvXc9frqq
DdFRZzK9Yvmry8n36ecQ+hjG3iIGrq2aATXyPVj/uVrSGn3xN5DyEvchp9dA
hj2WyxdTfrG+fTTM1Ue4uCyaEaT134KFCcYyHHj81v5Eo72zlJr+bpnsI2Xf
K6iaJQUmpuojmqM7mr8oMFlMNNwcwsc+bzpsf8OTDblrnIXB2/CPCu8JUdvj
U096SsqxZxOzAhWDj1O0rB75uduH37CPcryukmZkgNnJaI4AJY6w60j3f72W
uEiVUf5R/d6AfShvoDovlyzzfC0RKCGiQ9EizqK7iYIsNnUWUmx7j9yzTQIH
7IFlhYSw/2fkvL5fWPto3z+/W6omfxGkYYPZjyOjj0HZFIDLdQyN7BpGvsdB
zAI1NQE3g5EdXrvLAbK4BfK3pld+q9zFcwa3SMjI47Z+LAFThlWVQdsBFBwa
SySiJTED62/ErQYVs7aH+/zPN0Nd5W2ht2TCb6VC+TzpxnstuKQbuRCXs1Y3
zmQRcWviOZUiYDte9b45ecn201JSzIUgKk7o+wQcq6+qxkZ7MFMOhVHPMJfG
2zwsDsC+i4RfDNwVZNS/Vqq7r54vLEjqaapPQKvlbUhipSyD8p7Xnvr96c6U
l3dh0xOc7pctW7/8YgS3eKFTDqvpfaH0KrtsinaTAZmoIxi6BxF2Fny3AeT/
/07IhxijuKgzB0mTgaST8/NODVj1INtu6YasxSflt1fibQ2i30EwWRskmz7A
TGs2YZbn1IZC+KVBMnx3ZRqjCMfyQK2b73VL6gQ7Oodbqo02OUKiNTnaVrY/
OYp6B740tWfe/6t1w/WIXViR/h+/9zMsdNQM3F/nazdncDvjq9FS4Rk9gRxv
rpg1xCwIIMee2cfnZSBWd+TJLHMJBLJZbxGpZA2rwNIwHAVk8zsEefcuSRj2
HnmmoT/ihjcrspvh6lPSCIIeVo/x3k/6GaNEqlZaz3HPamKWPBXBHwwsoAWz
+qcGZo7/jZSZlIi7lxTr3dstzcjmjdYm5K/nL65nRS9Y2GfqYsdpNm96m3w6
slpkqvnQ4gCpW2iNV96Q+RvtL3gm1ciRpsY97lPz58U7iRxD/VqnPsQxOwRG
AT7eTnBAJGBX3ba8KD+oNDPvsv7Gqz2I8Cwoakw4vOlW3+8w3WKQ1hH8qC54
tDCz0G/IAAw/mKtNiNN0ognQRw8N/NXyJAveck6hCetfBU/ZCDLNQPBZMqtJ
hAbxqkvUHH4SQBFDmZc/I1ULWX8PrZhie6X0vDmV5IbJd9cF7LLxv59paRXc
apyVuwb2kH0l8ET70pBSCHr/5HAqgTBvbGywerY2Vcvk7t4p9wgfvYsgDsUa
bjsNWKO+HP29aglC5GjVCdpltmzR2cEXz5D5qeRtasyIoKsV9jaxFk/F47kf
JGXfeMfK328y2+7Xrr/OY94t/w4BWB0taT3sSi0hj8DDPpBvVdai6g3QUbls
adenI8Nh/0KiVHMKYbgdidTWb4fYj7PK2kbnkAsRATQS3dmA/2b3a8KvTjk5
OLEgbq2CZc0vW+eUyaWE+8Irc40d+/onQgsN1wk3A3Ts7lZTTEU8QnBx1J1v
qO+xkxULGt+ncR7ZS21Bf1JGxecG5Ug9bpMYNPTtYVJk1AM6IgkdwrYZ0NqB
9+LGHJ60pnAgprvdVif5F9QG2dxjS4xZR5BhXB8ajlJCPPgBn+LSvOXM/LiR
gDHfkwZLe+/2SSdi/YSjXwZl86Sq5lpRXmvagq3xBrH1xONcIE6UjybvK5rC
t7CDWd3pnoUqgII+xMxBLrkxLpQwJCja8R5iVG6qPVbcZf+aySVqNY9ZqTbs
rwyl+CWAjd+IAVU0tbKPmw9I+E3r0/SACIBean279tDdEvN2kFKlQLAqiyPP
yDi7EIxo5M71vk+UyPV9U8mchPSRP4tLbAsPCuVMjh0dtOkEJT3V5Bm2FyLl
4BsgjLYTga0Csbf/LxbwHdISASpoMSSueqrqDde2ZMbDzIO9Ex3JDg8DwYZf
skUktVyGQgVYeH9Xmw0Hy5ALqIBWAXoEtoHDZKnReQtbfxhAhMAwOHdUwX78
W8NxLA1DsFenH2+SVXQFdcgkmvDMabrTQSUBhc2lcm2ojrTOtgfEVPLT3wcB
BmRyNDqdbvsT2MsKqFB0BeW/9WHdWUpARF+s4nWhfE6YecyzDoNMLLQND5Pf
nXOXYEUmg2WxyXhNERy/ujpDsTTESxcNu51Aa5VrPPV7Dvz41Bf1wVJtNknK
AgzZs8bfnhSlhYF+gVKx8AeDxtVotjbfgmIEoJm29+VLB102Lo30xRsqyjb1
fgbcztubhlwTdf0NKXOodJ0OEijj+N6+pyGt8+BBfXcTM0ojNdU6/ph59noO
uoU75gPQo/44Oj+B8Mtc9D5DqH8Rt183PHJua2apgFpOm1ZJ5F5H7kwlVbO8
ElF4+83qUEU0dj/gDrMsnjLh09frRqSNsPWNEhclpy0LlXjED1SLCPxXziIm
H3MCpWsLrPuwLgtoU6pzk4qHpTzRcpFglUg6nZqXYd0DqZmpx8JvJCA6rmbb
9b+qhiGZIebpqRt/bw9Gqq7hnWMG3/dBCT+u1OYp8XpMoU78ELbPi/dtthDw
qNaT+hULvs+Q0CM5lIk3SmPUz1gHti5ae59bCP6efNigqQBdVZ6F1hr0coHn
lzc4FcFSGEms9yLIQA1tPqFPAvIIpoV8eT1MhCPvz2uhnqInOC0KPYV5J3lX
K70jbcp2SgSYLusZV+xNhEPjjIYa//m4turqH04EC2ZeyGOPcl79gQ+f1ilG
Egx1GTASMNPqffKMyPGCiftHRftmC9EaMnWmeu7an/BTE17+qYscHuPDOxxN
sYZ5h4U7OBprHAcyi+HwqwNQBdtQK6EibTIAh9B3B8dCOeR7rcGgkoCyl5Va
/O36lukFF01umLmcB/D+hJHIxpqTBdWUuhaJOw1//pTE9epjvnYc6nfUAzzP
vQ+93CTeFNvzzuF8ef1ALHz2iN13AwGnNDvKPzGlXmEi4w3p2NueKK/Q4xE0
xAYTz6LADIWRx8XsQVrr5RhTshMTPtwzt0BMeyf/qNip9g/5xt+QsHLpjpen
2OSjmaM1Pwkd9nhrXaVbx3fsAYeqXBVVKxSYgL/YmLpmlLqrNLFJQirxD/7J
0q6HlgODQ4fSPS+tqp0zjDzL50zdQTb8G9O6aZiHkRfjNxQUDXvlRCzcKwH2
JOZNUTcpoG6vGGHoGBojIXgCQtf/Z0ekb+/2E/0Z05QnMkx5VPWmjx9bMfaF
8fIEwOpl7/dhOLQQkZNAvEUohcJ2L+AuDAHHmdhI2ip/ptvtRXUs4wCH8tGN
UZ7rGns7RR4BvgCEbRRSkwhVoU8HXNGKt0sw8+fYTO0IIAwSXK+b2NrVp0/I
dypa4cHxA05loY/kpqe4ZeIK+G2Rl1IK/F8Yourgm8udCT+Q/95uTV9mL3+m
rVs1wWJLh9xXaRvt5AnpgERiDt3FJFRlo5iG2T14GU9jMoZz+tcdp15Zs+9I
GitYqY/F5NlX+Y2VqalcyQtHnt454kWAgzutvs1zIo4QDqZNZnubNlgfEp3k
Kl3HdDynS2gTy9hkU1cDZHM7zDFZ810wgrbhp6GUQMFU4CIm69Ey5BiksvEv
Msm9wnjgDcnjlZ0iNYo3JPi7MLRW/4wXDEESZRut3hjlKexbPbDXRGuG8we4
6O27zmFH2w2RnbCuBDWqE6tNuVMhA5wmtaxOAc1swsLdy5gRToECbRaTaJyT
fVaLNNSOkfh+iJqLzJCq41PeQb5sgdNVSNa+UPIZHgaPbEO3sw2u66qnTfOv
Gey7PSnxWbaA2AzDDsVL2lI0A+2dLh/iUAynoG0+iXgBJ8YFaKScJkEn/V/5
pKoCduxL4D04LFj/NTDgtF0RgC3cD/+dxpNb/xZYozX//HKzNPYfrEb3sI4Z
pGnUSuYF3EVVjCTeDXkkA7KvivV6ILit2lJTmjb30PAUD+oowEwN4a/qh+6n
9kqaOYv4J4T30U1QJ+1pB6aDgjpZJtWj92+WaVg6pjc9gycw4gieC0fslqM3
4BSZ+1kfk0gtanunH8qcLTvejhSz6TLwsxBHrSdPBdHZDsQOnmyR8td1IIf0
6XW+IKwBSUugHo+w8K6fZRwToyjr7nYBncf6J5pajif6Uzv/OQqKSccgHaDH
eVdCHOLBWMDokxbmi+Jq3BiqIJHZrvvPjmBglDoeN0B+pjISMjMWrQOo9EEc
6d0Uwo9IaCSMLVYYqROlj4QGaw/PUwzQhBRM25pS4DD+J4iIeJE5NC9kVMs8
f9mXIXvLsQRcDTI2pQfLMbO5s7ApyKDqlbCok/hUjPgBpmm1qIRKXk72TbzJ
JdznRIYkDLIhIgID/CbkfYsr0fZ2zYeWW11UuAgqm9JKh5jw5jNXvlUZLity
n2OYRJ4ZLMfpxQzwD/nzDSzDCdMQRW4walMoYxmzekMS08EdNr6Rvs0XVd7p
/s6JvwM9pE12hobpt4f91Yw/Gmp6ukDTweNZVqdOQIsxL+nKgQATEd60n50H
BjY37gQG3ww3rXi7XGeXV8AKx/rOHcvKSKIeilq5r2IG01j8K0C4KKC9Sszl
WlRWnHgfTAOCDqkDj+U2xD1cyguUwqeyU1q9goCXkSFQuswBqlMDLxt0wAcw
EUY/e1l1gtLNOqGdXSKj0d6Lzzb9kT4tcY36iuwL6bvOhsr7A3WrDGPalEz/
cI7lDNRkwGhDCUlxztWDfdWy9L6ib4u4RV7m8pHhf21I/642bS48XpT9CBvY
eqkSTZzxbuRkoLXMKHUOFXvf5TLrMbMxT2F7MaWeVxYjv/ZlxdlxwlJCwrP5
46uwwsblsTbxQlFmrZ6QvgBixYpJdHI50vbiIDzhN0lqQjTOGUv21BFOtYaN
6XBRNuYUV0yRUzY5wla/9IlpclWOQwqnXYkCULS4ulhBJxz7Rs80fhxXU7qq
I7WsoaLRhe61ZZ0UNoiUsx6qnNcaB7XWTXligCBVeCTIeyqr4D8CTJvtKQJn
Q91+0zcx0OrM3d6HywzqyhGKoXSLZBJFBvN68r5Yg0aBP/jv4LmTzLQ9mtk4
bwkGX0/efNDegcC+BQZe2uMN9Y5R2uAAE3NyPwUcCmKmUUm74/MfwdZMVJFH
HbogsyLFpCys/1yUeA1nBV2LTl8/JKbYoEeEmexbyAU1fOn1SRzvXWFnpwuI
hgWj9ctn/YYt5e+cHPa4C/ODSzz1H1GcE/dtAiRWD7RVwEnsDJSIwpMCtwR/
grobMjuVWSY3SpVAPemxfRSbokBe4QeoPasmrXJvComzXdzfGus/CeLnmkCk
SpBbsWNN/X5MbZaD+3yY26CTipbHa3gb2HwaiO84MBHOYtJ+/K/XRFQur7kL
50mOB3IbXU/K4cH5dhp6Wpa4EiW4Svv58Qw4kf1KtTBOVaqz3n+lLO9JkCXS
9743q0TFlxsuvid7qh14aiJY6KcKg67SlhY4WFEHdJG78JllsBGFquNOpt0S
AKWYJ2hr1DBLZwerQpsG/CdeZnUs3C2bkvxrGJVCNJyyVO1P/54nDH0bA4We
wESkM9gKeYG/XPnNqDWycYJhxS7OsR/gxR6ZN9E6uaEGr1MgFik7OXsTOs1f
cl/1SRqyW5ClCt10LB2tPEGq1bSJUofI9/J8d9ydEXhNhimOKogJPhut5TE+
U9zZTVE5rIbUTpNpfSwKs44JstiAe3yZVrjF+nzHP9bBZAUDF/JkOArcT5fO
QFZ8/4ZRh1DD1XopIzLgb4QbBPIyXWYN5EzXxwNmZxpau92KanbIJMghHW0X
PdIlknCCysJDOzSa0i5GzeUoRz488pq8qUZ/LqJUdu3Mq0CjfVsTVjDBeMa9
JUE3wZZRa7x4B66X2mL5A75zdgEBsbnDIFGr3k0cMUpfg0ZO1ouKkqugBeON
B6J5g+dtr0UHC86BnoM6X+Gd0FB1tDeW7E1yaeZYsxAgmq02Xikrd/+l+d1O
MW2Yv9aoXkbhSReqtjHvOABaXq5AMmAi0Adm4s4PnU/nTdNeeMq5sfncV+Jb
rPl77kOmgERQGa33vsx9uiWIPeyNVUMyRej909CrxIdmhw30EHVjnZrYAlow
vsmlXTGiG6CV9lm4KzsMPHHHn5EpDjsPBK74gnfi9/j+/GsSS3qlDwq6HVda
Wznmh+cXEyozNsJ5T/nPbXNc0ECWwkCaDmMkGwSBF089qtrnfd22IFA9d1KQ
8HtfhHdx8dqaWi57IH3gu4AkKSGEabl/ux33VXcc8eMJSJknyTnC731/pPcr
I0RWPlChoXm2feKHs0blfsu0SxGfU8xqefzWd9Xs6sXpdv+SHaqleCs8fu5l
wtTgO7ID2gFH7fC1+OL0gSz9fLBRPnUQwK7IOczpBivRFAR0mEpcKAyGjQ8S
0n8KLqZndcAkjJzqYXEMEGQLmQhvWPO+/oBm09hmuFEJvH9xVay+89EumUkX
1ggshifCkxsxE21hYVWAfJJtRUDNHcDDO+Y76iFKBM+ZnhVhQMZtK+GbNpvb
5Fn/NN1WFCWICEITLtUepsGIjs35NlsJ+li63srNlczm3bXlwLs/tpiRYPEE
9/FPbBMEF01U3907ix1uIyk1ODLXXk79K1g1OT+7l3BDt28lXvIOzRJZahDZ
0EredzPmWKP0pbURhF7T45yq/TrYzdV7Fbptku46RBRGUz7Ve3gA/m+uCuXY
2Mk9NH5ij0avEwmc5dz0vWPx+LVmklleW9Mutn6tbD+qgiWjzf9qhjswZami
2hv/Xz8EIpPpGqXeNsCWDtAgcqvQAfdbVeTTKmskSf4Bph2mBPEbEapNOhaR
6jCxoHvT2rYf+t6dejaeAt/Mh+SuSXkxBTQPu6T1jaS+mMNCitWILnMQfv51
C39Lah4iayCgMXdRVAa3LEucOXR+XsWqoQu+Gkb3T1sH/wAS6tXLnHRoMTMx
sN5Q8HvWo89A0fE9z93t+UEB4/N+Zqu7FHGgbUS/Av8c5IoMkU8hJe277llf
FHp6WP7NWUuPAYB+lhZTU1XvWf5miiW6LJ2hcBAc3lAIsjT9j49umE/ajvxu
ULXsZiW/1UetItmdRUwgPtKtmAWe6dQMyus9In5eKiRsLGkw8gco/VX0HxUJ
iphOkFsRkxyznF8nBXB1axrbCuO9SaKWEQ5HVvpNZu3l9WtxvugfLMjRYDqz
saL1IWxpmRs6e/NvQ0RUnu19aC6IWu7ugFPpwlTALCMQZp5stvx2Ue8qj77l
8+OLr62aOZgtO5CAQGJxZcuKTgFevEnXndg+9JUe2TBgebgkxe6MOypX2p6H
cxwNyR/LkloQ90CdViIA+YW1rvaZOVinJ3dKroEOeluOp1CnTmfsQE6opE1+
hEN8Ki7zYxVC2b75zTOUGAUyl73B+4h5E995BbjKPPfsvkCnFr8g2ulfSvJG
cw0dhWpap3ZyNG2suPAGGobDqmGDA9qlppV1IU3uEoVAe4ssxAlztPsLc74N
klNy/3tDyI7lyh3lHhFooeJBZTt4YYeN6VbAz1Q0br+h2TKT/nSLkHk3Bb44
axAxFVOLbhhvvT7UsBNrNzFG9iKDnzKWqxeI9k0dBdE6VdJEUTG3sdMCWh/2
ENSgxh+nlAsyIgqnH3BaImsZfYqoeb3MmTOmAuxY8p/g85P48O+7rU6FYCRb
nO28c7boNhK/AZT0b6mpN6xwtNe+Hqt32C9RJf+qLzjvd90iuBOhiAmv5qg6
SUxw1F+dXrVqSa7AI69nl9BYOSLdUOtb5or3KeuCpsO28+jx4x7kCzSXIEra
Z2hZPDg64xhujMr9lfWBDmDzq/p2a1d9167QJu2fvJEMYQfokkfJMsBtNr7J
0xCbQDwkaVDxD+5jG2y28jFW/9A1CX7b0rYnop7O/idTD/J/mtLzptU7KMhx
cOhH/JnJaWlptQ5B13eAlOIZgMAVMfPtgC4QjNVWaMzXve9v1KxRHcPw/YDh
FGkxq0T1HghXV6aKZd4DsI1yudxu2JfPUscbayitN05N7yXlkZiWDyDeiOy+
Qj4sInsreLu1RdLahgV99Odh/ocHa9vVi6TySW/hGrMmg976O+7bVZ7l6q6J
TyQOAyBy6qT6nfjl3H/QXh3m9XiHZBmrq1pOJ3onAWzBt4OnFbNGvYF6dEOF
xie680hEBAWl0Qz4a4bm/uqNL88fM27DaM5jGN08oT662ucP5IxldZ45dF4V
kIWyyk4Ms7+y4pe4SkYZRRKCkY+zJBYYu5Onrv3cVafKaGE0zT4pWdfMb0HS
tMzZ/UMJyJX4kSTFCRhWGBdQq9JpVSjxD/xPMcrA/8MmMKbPyc1cBm0uLl68
zBGPPTzo9DbCJ+sFPPCrAJYBHEZO97yttLy5+UA9GZW+VUhcjLCWLu49aYKJ
hL6qjxj9ry1dwZ4e9pQ1UrbUBLKY6lHNdKvgrKmbu8PA8zB0wI12ljLju2XB
8bdowGOYEO/GV2BHta/TYMsvUyxkA0C6wpG77zUMRlnnkEEuDgmMb6OQnkzN
tAP3BHxb+1Yr4kfgLRkuf/LoYtzZj0FZ0ezDBm95uOO8UEmlq9CmdjWoiH+n
6l3QvvPqbpkseAeP9mFRVwOa3Zh3FNGz6DSZo9+RjhMIp/Rtsy1NG1D+ktAG
pNeRxcazfWdM350xeF+ASe4v0aNk8wJEfp78wFKb/FLZjoB6oJOkHdQtupvU
4Tny7t0yN0XZ6hC2/rd9L3Ben5itkchPLeGO8xW/Z0Ttx7QLtCDo9gdm7kak
SIMAQR2MJ+VD4Z2M7zy7fH85HptwngiWSPfN7OlROO9kZ5ZCerSdWzjVQu0h
/2fm6VkTLwVSNuytvBpaeNScdRmhzMjXA79WRExOEgV7Ne0CfNYssLUMRHk1
cpS/QUavWGZ+EWRgoN8KInYw70bLvWZI0vcpuV67IrN/EvPKKmADDx7E9qnx
IVPeXscdGfOdkKDgSWwKN6DtegMLwJZBGkKw1hSMIG84Ln1/R762rJ4RctTp
oHtwhzzAg2qQNCZhe4eN5S6UGvim8aaYuJrXZ1ZBfXqs6jLWAeZVUTAW1I87
YCYKO5cb+E2zP1ZZTnXTlPC6Ucl8UlSF6JTwZ3SFt7+504ZFxq1YA83+2M1V
CbOhpjIr7si82rE6lY/F/h3c09etOTO1ptTvO7OhqIUz5N+lNFm/i1A3fLVE
H86N5rraUdBVRTvdbc6NZYtwqianoLE3oG9NdeSLZzYHPsg0RNQGNh0TW2vz
bxjQgwdDsm+BWueZwEtvKow1SqYiXwaNnmav3famvANAE4okWSh50faLRN4k
NxHlcR0lpV8QEcCkVuY1mKx6ETax7WZ5X1MtoIWOu9YrhOppkf6h8xwEEryY
irdG3jFkccU3l18twmZCTro1krgdnBJjccP2iC0Wozc7oEC3+HSmbsx7T60j
++UwkU+GIWFPPUaJi9uK8uM1rq88zTeTU/iNBAPGgPcY9cvqjCozWdZBRtl7
es6a9DVDA2MeueACZzszD6+3rcYWn+oOHPpoRnzRsS/NzPpz5Y/aUC1WzS+m
bQnswIZsOtuLeuoMIulTY3icNvxWJMwpmjzcsW3avGcWZNLD++WVOocUlcG1
e2+b/vKXxcHjaS5z0FdDxiA/cuXVQOoHAvElfgEm7McXebz1Ovn0tEbaw8cC
oWBOZVhP786FLANl5Rj6Py3jkskovj2RYhfNBJx76Kn9BVrlwPNAxs+52R6T
bNUYhy7yhgHXr+M7iXA2Ms1fEHCb3nnrLKPCJAOd/kkDbjybngRHMfb6fjGn
F0pedmGnbPcgnmh0ns4Mt2u+8eNoFcxZKg6opOwmnbwZc/OkP1QUdxbZ0Idt
ES5/epxVP5hmdVVWNNG+z2/9uv1V++ksQ9ZmLapB9SUBDRO6poM98Ts8bKTD
JWn1bpOn5Uuarhr4gx7fsUEnXdMPEUkbaLA6WQeBhRA6Wwq8qYfip3p3U1BB
l3G0Ot09fKTe64ytWyaw/iiltF+cWHC8sALNfiRbFTsiGWUvZEUBpe1W0Xrt
ngdaKyOEvQmrk88dhPrehGwaEiGI1/hj1v7BRQ8pscIJ7aQ9r9xL4Hj3YSVn
ELKqhW8U94t+Jm9+TACx3oFvWoX6ro4pxEgywJ+QP1A8GhNKuVa3QsuQ89vR
mK6xg+On8Jf/hRPuowknjUeCNCR6m19VhfyEw3xfxwF3SSHxLyenfFfwNJbm
4kKZqx2qIx5ew93qY3J+/fcDAx9XQ3p2bFNTMhmN7BiS6Z54ADuCICDBJVmz
N+0gjwgaKp7gDSj2pbhGKvKQnHaBLrb/bobYXO31Ocy24PdwCRUEIKYG0lnA
LQO8edtm7qkggwNdAiSLPCJe6PGjJ8OkTsU+x7kHnqV279ZdKS64ZIsCkvaQ
sIhz5Y8gnRp2VOrQBPc/pnh2mOu44x319NB3YbnVvBOFbhrMgnjLMhWeZZiW
HTT2zDOdQfmTtPIpP1JX8KeD5FapC2vrjgibGEoXGeSBKMFhk9Xn9Tv2O63V
A7oQ6qed5RTNdhxKtzU2JPAATHmyd9czHsYogDTv47EFjZoH/aTPinx01+q3
CHu0zw6RNkA1HdON0ab3HgCDnvOMR+Tyt46AbcsGkKM+9qXWgcqPkqFz9GnV
yyaKfk0qSEXOVXdDoNkA+wLkR4HKUT8BwvBaGECbHyVN8nikTVhmRaP+GGNb
y1TpNplyVOuFo9Weho+mKsWzZlSjZGaiaGe3XEmJl3ktaUQ6782RGYTrcclq
GltvmORFFT3iF/waHbpKU3KA5hgNi+ZmZhb+PGh4WiUiEBXJAOT6zVh0qEZi
iavCZTYQrHm8Tu6ZEKnetJa/AyzS+mJNcRbrib/2lPeYYBHDGWbc0RA+DO3P
dLLp+kNrJ9nnUEY2H3ySbFhr9TK1ltRQcPh4nCtcmvpjYTiMUoQluh6NxUR4
051g3x2/0l6w+enb7QmLBvPOu1k8dQWVXvOb2xsqFJdaLfgtIvKwDtcIeZvs
5KXMDhLK7sp0/fppHgpkNIZVbE3WTxgcqG4D+fR32OkxqEf5SFpIfNcYFbeQ
xJB6v/wyno0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpejUCrXCERvfda4UnGTLQfmABSG4vlWWaw2i6sBApc5v/6RagmsOYEz31rRlkrimtv5NWxUmvT1FL7YUnIkRqVjhVtkJudkqkHw7idiXJZC2qoyOUB5hvp/+J1eud17TRGiQPY2lTgtwGM48H4mWwjTVMTtDT3Aczc1Z1z6KtR0wmCMZ60k+zY1lZO21vK1HyZ4n6wDEHhcwsZQS/PWZenLchHtMHBfDnEOHUDE3IJE5IX7eURlCQJdEXUwhN2+s7JSI4kM/dbWyGWqTde2K35kcG+ZjC/sEisE5I3fRbrwEI/4K9UeieLqZRMWrTusySWmDaYo9OOJTFp6pOjsxLAQm+g/r/UKbi5hg7SGz3FEy/5wflceM8VL6Um3gTldUPciezvCfmHUD9NpPBkL/ky1hqtvyUynFBdqitwhM5atXLUU9go/oTO/2PGv0ZtSELFQZGtmbleRmvWCB8DbT2ulgjIMpsviyEprEF6Zc1a88sWAXjOFJzEfsDpZZUiOaLiLwBR6rpHR9ScquO/CaZxfiOWb87fe79gL4ZbEsQ1TfNEvvOfadpCxpm2jES8/uVPwDB5lZ0EzAPlgl2VOPa++zlYf+nFXBRB7z4dKdPVeltIcXPW53J3NcoKMsw7n1rZsB7YIDn+wpRvRompRLstNjWc1ch2gnm1kKTwY1wWdE+h7jTIHEstKyj5uxSavA4kG49Rj4VG5v3S4zov8OrJFh7MMD7PPLauOfU9EzRvSKORNhX3u44hSCIWQUDJwu0rmMbNJWKw0Cwr4SvELIJVNj"
`endif