// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vN8/9AhdbJpSMkPpxu12VE5h5FazTslZvWba097Pvn/L7wMIXKSPX/DH3uNY
Qtdo38t8juMTF1nvV70VzTeXZoiOdLXnxm4psf1hw4SiMUXuBcHkdZFFvi/0
LpQPwQpNKUyaxJar7OVtYVRqX4hUZH54OxpqEneJRKi4qZL5cxcokyLRte4r
zvYT/3ogRGmgbjhHoFzbkII95EdCYg1Pas57us7AoP1Rpg9WqiaYyPPUsV2i
U18iBTTkcXDPakusA5lImfByHMz3cmFXG26gk/P+8glMnvvt6kX7b7NSrlEj
V0tM2qXrWgL9J5kBT+YRCV2mFoZ4QXmTGh2jzXR/Uw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZocP8U5Wr73iAfs8s/mcDW/EZgDTUFxzZjOD3+2UKgJJeEiq5aoKVzuszkqY
KPBoTCLpigDGQn2dxEk7vexzZTkenzN86CwXxkUCOffh4rgwTOG+l2h02S31
vW6jwPG4PSQJy7/HDttjO//8WTXZWsJ/rFr3jxgmSRUh9IC8JM0gs21GTcm2
nyzt6vdRS/HenUmBq9xD7i0diGR+14y3VMRfCSczTIM8iL7OCanJtgxmLOkS
VeqKPw91WKZBRC1KTA6XWZ5pxoVPQGE7SLAfbGZJq87tDjsZC5rGtsL/ntfm
UkDWaBJHXf2PFhIQLNWszJUhhJqU+gGzl/B2gIOVmA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uEd5nQGyt/IOzNbC4OaLaRJULPjWFoKGeTLPyKbN5wSCLeyhJY+iaN5O9qBC
WA6tbtPsaLBk7dGGQfDJt/wGnHKQ0QOeE/f//16s72ssjC+IQ21wEO469+PF
Ze+JTirDsCjPkoWE4pMCJDrOaT/8VOCvMra5bG1Kr8HGaBLOVpviRZJcSbr7
T7aLpKdj61lQoy+Smh+uLv11KaV52r4CaeSLAKJ+bPUDyyFuS1VcVG6XaiXw
Q1TCsp0gLKNGIBduZEh5CG4dUXYSuR6ybthA3qJA+CdqRd3zwGpNtwIS3dC1
pRafdla3MNshXwBSRi/kXGCPFxab3H6saZHJDR/vrg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IfAG4lKOWiluKvJEplF28oWkfRUQ8QPF1BIyM/gtm7l9DfljxT5huH7WRxyD
T0U2TGzGNI2fPLFDo8snAMjWN8ltAHnqTAdE/TqK6W5Gl9zLnCMnxpN42ILT
xPwyk4l92fjbfW8jJe/ppiF4bqfVmOaMK7On53kTDaW2ezSyhtBopyoGYNT6
dyPhuNw7WVHEpw4lo/hv442TVPReh28xpsOqnMqqXR8JmSKW79izopbDk7Wx
SsYX/nnFD68AcE4BKHzNi4nohXgSQFeMHX3GJ5g2wDjaNDrAr6cmbLKPwwn9
aNdWdVgEhAm87wg0RXgpTIWQG3VROLEv2dJ80COOjg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eOfXR/h9GxwqzSvWutQZKPvMebOnsb94j/0TGgsUNNJl2+ydpAkDRxhX6j1g
T4VnNqp8RFKr6sXEuwmz1NjOGmXbZnqXZ1HZrcxfpgXEOxot0Qdmpr7jVf1R
t6CO3VA5WnP08UE22Xfox2wPE7kSgK8iJJeL+7WJtSbQbU7eMWk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G+2QPhp6sm5HZbV638YN2SM5Jguap/Xs4sMRCcpGe0vsOr4G3vzx/0WjrMR1
B+C86biN/cAH31bddHicEhzcpXCFwf4JsNO28gWA/6b/jDs4IlALXxM4YeSq
H4O9Tue1NB6TUT25eyMzXndGCiLgaSFhaAznQx7dikVDLQUJRc3gkO83tFwd
Ivk0te3OkrfxtVx1Jxo8fc6TWwW6NUURpCRMKdjXsHY7epAS4zdXV2dcQXHo
CttALkhHCoqle+x4RZQ2fbOh9DEYkXTDC7cZV7AusAvjDm+ZGvMdOOxks2W5
fQj0wYs+mCHuTEJM9UacKvxfIwfdhobSAXN+wrWe9EY/+Xkj5TCAgiT/lDlA
H/0uJDG9lOBs8ptibjZjdJ2INpB5escsi1MVKGBKIrvnXEssdB5hzFXoZVmM
dDV2Fdf0524d9i0TxwWY7aCI1VArwuFaCkwkPgqsrRdvPEGxUc3Igf0DpcxK
hYcquCQtxUD5Zadl0to+gL6X/TSoSqje


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H0wbnB8SidrLIIwaTCDz+SgPkSpOVPmU/Smi6ihsg+Jm4MYTy3BUJ1vLQBas
/E4E6m/25muqblGpsR/iNWZv+oF0kLF+aWoLdZyE2UfmV89cIbymNDcwjzsN
HRROV50HM3O34aEwzcB93P8Qj9WGhhxhx4VVMncTye0q0bd/pP0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E9SviLG3wGH5cBc1wWLN5riLEeHH9PTf1w1F96vroSOcEx6oPU8jFPiQJnkl
sZK2xp2AZIm4T7iuEUxNOFqT/1wG8paGa1EdfYE8FxqCYFkMSn15ooxt7PmY
/xOPp4UhrRqjHequ1wU72Ers0wdUXlylAm4Z+mUgiI2GTzslVnQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 25728)
`pragma protect data_block
bIdotfOeOcG0+Jo1PFR7U8Z6cCUIEkrSyrNasiP08qK0qxXDVAHFXS9dVind
QKJ3wqArnFCsB5zYJPv9Yaky+9hOTyUNLdoD9H59MkUuKGJR1Vafa7QlxelV
KImnLgwRDAXwZLD3z23zS8HjaT0PEoLAaWih0g0ud6lGl7hRmzR4TxsD5aEs
2MHOBwsAV48Tvc7ulhKbXQl1RPNlfX2ZdA40K5r8z8U7f9zg/1//I881xb1m
fvOAwDOfrszG8DuqA7dqtO33JkO2kADcU3qTHK++J4b7TqJj0QmjZh83g7d7
YQp7bL2R4Y9E5hoeaYRMBo3ILRwIro2pL1YOjlpCAjAyrZuMVaP+McZu+B+R
zBEbzAXhSatyTSLkq4F95ttX4LLFZAG5wgpPfSM+AAJ2Fcbbr+sTifHkeeAJ
cNBqOrKYukoKLVGz6jxK7KDSEDoiSJzTtLJcmPDk2LYMUplHDTsbmhaZvD/F
NKrwJb/jIS0hXwE98JzP0HDHXAiRxIr0HXY0DEupWsFYzjVipK5n9YQdeBGj
YuSQS4eULI9XmsHskr1ZfZRamXwgNzG1qqB/wf7XmQp8EMCSXuIfqs5CI4dY
1HR3xDkni1Dg/Wn3fyelpG/ed62bnrtW6O8E7SrUb8pqs3lv5NVnZbLrmQ8E
9mZAB3rku2X6wD2EXjr5leyfyavWlVuLhSonlzAyhN5q2v6sB8XyoDPykMZv
ykIOumXaWADbAAKOEgny2/xpvMatmO1zOZWnVBcY59G9EhpCjVjhoF5unrwG
lhHQ9OdL/+22no7ux7SzIoi8VsLTA0B2dC8mkkpLhqAvOgc/sHnlVFEulqx/
8FP//DFX+OkYHrciMgtqheGnjghDHNHPHqhY0r3wpiIYC+g+CSeIRySSq0bt
rvx5tfL4RNUk4jK0HXnx/5voVPUEeEJBd1iNcIhOWCFA95TlS1Mef/iPLqxe
/2gYSItHeR1mYR8/Si3gX1M0PsnRvGqbfgASM0YDzOd0TChYxfBvAR/Z2Q8P
eGys09tBwPSKp1qazd9bwldiLqFfFD4rZF73rBH9gVTnvi//Ginni07fiaNS
DH4XYkz6xWJ3ufDekjfGVSIHb9AogXIdYGQj3I9MYa3NOJDxbzv5ML4yXggK
jh5gP0qhCX2Q5IPntFh6TBa1UsKXi8714vSuVcF6ZMdR/aVSg5fQNROqKuBU
eemedvxkJ6LHYSyvY6KC7femS/L/ecFVs5v510M8qRBgEdmhL2TRABRsQHoY
hIuRdr3rVQ+PwL7n9deKqIVJ2rZ/TrRvL5Ilyy0S+DgFM8sp6xvouIF3r41J
eTZre5ZsNfPa9m8CuGGI1sU2kXpf70aA/U1lFf8BQA9Yd1xEyLP7a7tDS7nY
YG4GfqCCSGArqLh26C3hX+e7AK0IJZmZm2TUAtPZnOEHE1l5/f3b4V6DX+Zw
erO+p9/IyA99KfNrDxBY1++21e5eli/gPNEqMtsV5tWBjNQ25wWq0Sjfee53
d8IyaEk90tdrEkwYFROvy6XkhiXb3TRWieKculKmxeRVwvuA8I8Np49YXlRL
ysCnxvIdCjv9qpJG8CwBFiGl6XxT71s73svA3HPp0fGk3V4EUR/R9lSya4cG
AWPBIFI6d4+tlM1BRPLM8L4LvUgL886lRKA7hfdQnFeHg6R38eTITZxIMjEe
QA4DQ5aU07DbjzBNezvq0m5sjv+qu8IV5e7LLeCcadlph4+Twm+HwHH3qo7d
Mh9ktr/yxiiWSLEAv4Iffzs1QQkph5wBzXQOnolTfHyfTtgqcqrsHqmuTCb0
kmYqusD2drSa77c60VqvWX/t9rh334rAajwxjsHOWKy+aRAYuLu5biYOaPLZ
B9JUCq/Y7w/wfBJeZ5pGJbPCYOTKJO5pG83fS1AMkZhtWb8f/EPU28Z0+KF2
Q4gXu9vMfCVXYSXhxu0G+YXmw3TJMK1MDJ6uqTCttLua5XRDDjygTAbHltwo
Hip0ESv5NNLQu/OpsraVW2hJVnvK0e9gbW2MyNOhjhzjB9Q8kkDBGlKhkUx2
XhakIlB3OGzYAFRR6nZPebzDYhzy+0teAXlgj9FhUPmiI2dvoVHooSFXU9ej
/a6k4YNo2fEm9WboNwAhYZGYiJbHLiOH5m1yyKuNlT3Eb+C6wNCH4hVMo1B8
Hasa1buYbd4VoekYjMKQv/kFtdRGfoqjNFk0qqAnZmOs+CRjP0hA85zZFHfQ
iW9gKyrFyVIgoKRIgRjC22PuvB0hZoTFOUbQ/RPUcTZT0SjRRy7otSZQaPoA
Pb9fu7ndaGck70mGr5x3gX2Dtl6cv+GVoonIfv0+Yjteo9t5ReJi1RE0ymwT
sMwrN9A7E1RU4XXt+PNZgeQNhnnNnAX9pPYaRSqASci9Z4Fr0IwyLlbIT2f+
WnW9QPuD+lo9/KXbKdLH9dqZR7rDeBPNqbLbJ3+nJcpD/5pxwGaXsjfN9tAZ
Dme6CQMbP18o4Je0RZeISTgZdwvOYAfed20vPd6srWyyHbVjfJFCJniu6P0C
fF6TbdYAbmyDGql+FHW7f7eO+BiyhHCUUyJwkHqRb0iSsoK8NyTv9e9wBPa5
7bKbJ0aAFCLLeRAq7+czX1zDX+iJ4oxgx2WdBZTOziyuvX1MOTNSLHeVnIyL
x7HhqzbOw8TETnHTkoBWYjAtuMlW2iFBeSouZmwtqTrAcCvV2qfksK1PJDDh
cFB8NDDlaLXHzhqz/0ZTSZLKV43Dq0bljq4FyU+qZSqkUQe0iM6Hl/JRHKgZ
V4AZMiwMmMT126wquCLyg2tO1wk07PX/4kFTjLUikOwZKpOdGfRN/GUJw//S
Ey4MZUgoHJEhdJSfggy79SX6bEJt0i7770WTlTS+EWvTU+MKCZJH9hTFD+G+
FzJOJ9FL0A9pobDe7eA7yeST0hPUGg9A920qlGZk9oIdUi7H6VlWOeu7xDYa
f0WZ21EHtrpimjPSSoogM3NgpSKYXTO3t0ZgUO2/v1m8acMo1s+jaAXs9nb4
jQwBieoBP6lqXi6r1XSN4z9KwcNKrvl/f4TNcwDko30bfwNBuS9o1fso8801
OtJ1IeApX/c5dp6hvxLVh4AsSAJq+8S4nn7QKYYFDXYwsYUDNpIWFJ1BdzCO
KI5Rm9g+D+BOr+fSVOQK8GxhAFYLN0juUFx80s5gdcEFruwx5+d1NMmQuBTk
WomV1kCZ1fiip0J+8/ZxLYcdIGnLjg1aL7Vl/bceIv9o9fu8ApipiSKHJe7D
WSGio3t9np03OaKWxbMOHeEID2wCHz1sMFkwIryLzGuvtZB4x7I4h7mDEYjD
tzeSU/hoR4CK6TVhJLTF0DQoiuwFgozajfr9HSwCj0Q+/fiGRrKouTcd/U2f
MTTh37FOmuoi/otcm2npE+wJyvVkiimKMxSluCRfODYoyjXZ6AXPwYHDyRVM
D/Lv062v4qU4WuA9wfb88cY9K5ga5+A1rqR/nojcXeKLG36nJo6PRF7IKcPr
AnyrFLsaxtDgnrI72FS4rq3ZC1qnXtSxtW6ZJNSdf18Hj7Zx2/+tLCudBrZ1
l7Kljw8egLAvuoaYNUyxccHi8N49bCngZoLZmISneC1xsoz7PHQmsNKQw0kF
/wa2eN5zgx6MsC/u79YNvYW9G6vQc6FBzHK5ROflzEWuHP1xuOLpGLLlObSP
MT6Y8bGgf61v7FybYW8LPkMduWqGUNrNgKMm/AoFUm41QGV2iZzSJCw4L+6p
Tp5kkD9W+QTQzXMaQw5tjS21qXA7K4rvp0yxMvAKjxrb/DN5j71+QHFsVi4+
RuWCQUdpuwtzNU75hiXrDq6e7DGIOMYO8gtDOIrBadyRC+9nK2GLQGkfweav
ySAenXDdT/ydAisL7HDbKoMDTLdVlOv/9D2JKs2EZLfIMbhi0NnwuLnUp86m
g/4r4zpINMesXMGmtUzEzP1+/KozulB+8MjkhHPt5P/50GiQSjSwE6ghyRcY
+ieuTVSaZcqSjODjlD/1qMUvWg0u/t7opp36kpMf/Zl2bRmBh3UVeLijNIm6
qQ7WfQNblKA/v5YBO0uEThjG8iqfOYbGe+7Sqw6tD7v/qJYB5NctlXw6vber
uacap3i3gIywY4xanE8e3PjkXnjhGjmZXWtL9/NGqnEaRoHDRMh/egUi6T5Q
1EFUYZQ94FxztPUm6EqNMGwDzALPtBsfJLacyvBRgs8aG+M9Kb+f2w0wWpTt
b+93+yIgQgp1wOZWyPYFtnTCQD0C6v42Cn81FInBQgscNDp5SG/6e5OvyD+S
deQyoVMvumWrJMIZE9VdCDQAjxewdqAFMXpxxpLHksJ/fM28eeGMR5Yc6byB
47bwwDXXsZ728tFU0a+M49ste6kEjm32RHd4IMGcJTwAAwzvNVy6n1qGVwvz
ujVUlFAc0qfdQlPki9MtU5in/JchB3Hw5q4qabeTaiqH8xrSFsepeil3CpHx
XvfETJptYMjTUzeJ/9QFJvlevdshnGgS1LpB+E9qsFk7ayvkfyQgaUQXrVwu
f5d3Jp72D091RsGHnqk0X6ef/AXQkC3xRzPUVl98r+lxYHscGcL8M1fKgjF7
eBBLA4PAePJ5I1CpNjgPTcBImRZJiCitsawezb7L/gfT51odeMWe4Ad4qKyo
GUnHRTnrDTcxvzXbFrzKTqjC1vJ2JCzhQpq55CIsl20VhgD/u+zDKD8nfcNP
4GspAjm3xkgdIkp2Ejbk+7guqwxfb5u9i+R4eiU+36JnOu05SgmUdVlakmxZ
fD/8ra7eln7D2kGwsbh8g3+quBO2e/iP2RwBQFvuSz3KUCYQc9hMRbglDp8B
ZeUB5h9gE8rPurKJ7yGSe9bg2BiTTxGH6QuHagZFUJHJ+lUh5hdT3Qo2BIZx
vHl3BQOFwy5K0EsiiBdDLBAk154N4s7QnphHe+JdbHE1P193p3nrHWhNmAoj
e1/I7/KAHAfUyLnSSwi71+RTLf7T0BurFxYovGSyAwktf3AME8Bn93CLPG1e
61MQ/hqhhF5g0msslzCIjjxPegb9lBVOdYr3uYBLSPc5MFoFRayzGl65jO+q
FzR8rf2nqNpVs07/YWtnVkOLZt9ogt19vFeAxuEHivClw4rdoGO70JVTAUOH
Fb17K0ix9P2FMjkGTFDTZ0mf/dGAglFky/nvRVzSXY6HCctXPW2DuPZPABFL
EC/44fqZHekMAUJghfwXZQ2Al87EMrAk6FpJJVvBugbzG1txQnQeNoA6/I/A
y3jwNPt7GVMvm8HvwQxVy0x2ImtX6WmiCaycHnpXtvQD+cZJsUHEpopE0ptt
1bax6icgw/+s3uv/OZER4mWBKLnqO4CwRfY6/rNoQcv/yNvwfpgZ0veli0Dd
oqoyz2jUsdujJQO4tD0jnuCEmRysRv2y3LcEk2GJyYVDA+ZaJhelPebMNtVc
vu0OFGioKlRG9CwEk8GO7zi5mlHEpxtdxdIjqr91ED9ATq50Ms1YSXElDA+z
zEP3n6Cn2G4g/lskzWauyAebJqxk6jXtYX3VohqE5shhUOAcc2Gy2uY57e2o
r5a4lPtNPws+TO9I/aZCsPgtExfNlvFVKIxwuEmyRzkvYEaNxHt3zJ+4MvmA
MfZWvJt9tGDTT78P5R7+WspyD4jjS0EUiXDgxhEXKTPklDiHcHv2dbledGnT
dUlJ1nWUsDPHHcNjjUWrhEpS4UQQE2/laE0ZVj5B8gw5M+Id9UoAgz6Hb62x
PEnUl+bIf7pok56CNlOx2S5JkNJX85rcC20e+SnSlJWkCjSNM0+af7oc9D09
ARiQzfkPfsGsxrnaL0QY9LIHRY9yC2eVRw8CtXN1RZxIopmqwc4FMNq32jyb
5d8LWmQNOzk3AncoDU4BHLk0c2/q7WY9+ToozmgxdgHYJlDVHz94PbxfFt6o
dizgjpFAwMI8mpv5VCRdmsE61XRXtkxnsEC7PVZ/x/4eviqHIfkfmr4gMhwy
DHh5kG4QeQJMnH3kTSpmUKOCioyQEESBp7gOnD4CTJIKWU6AUgkN4Tki8DXz
Xb04Me7EBuhgMKW4dMMMSTBUei/ggZPGGKDCskemRyixxBpJmC86UHFrVtFJ
HnFPPFYdS7We2SWZTumzl8Q3p7+mwI+UdKLfEZ6RAMNQNUcMdozgKOzeuqUR
ffSMA/z+jFWQWVyAEeIS0SAedlGV+0fAiZ3JoT2zxPV1RHmAd0CzMvpxoQF7
hU8MwWDPcreIPzgBti29nd1N/N646bdGJVxPRD0+buinAF76zPDOTo8cKUCr
f1I5rAzVSmrHVW5DwYhnll/4Hd6NHSPR82piiN7qBgFs8p5dZOUHOon+2td1
askPsYFx0yU6nyaDeWAf9pYpMYJ6Peada2JLofDTmqiTjkNVwI4Ylx5B+AcE
1eY0FmWNpA6grR42CORA6h3e4NNUihp1XB9/Gooz1qsIZ/B/wh098N2YDmme
C8K9J5ob1+6Pjuy+QZ2DL+3sdFtYyZtSF8u1Jx9O7LDxdoD/MsDoj/oNLcQz
iQ3pstIdiDuJfOo2xqf+IJzye9xRCi00pewZvFznQ1jbLojrijSyw1JMoE9R
DACDcGR+MW7MQnlRNgQEHMEY+7hQCAHSG010xE4JmNjqEv2CYPujmG/iU1zS
oEBjEDYm500Hq/Gb28NN7VRfs6iIeoFYhEC7neaaNVdywZ1Mb0vOvcHaWsjP
VqWpVuQfAxKpgKTyJvgUg893nmO9IZhScCQBh5ZdkrTgdXpOg9gWtKZVatbY
Vl3H7dFLwcfeLBLKPDLxmW0n5/wAPfK9AoTI8bt+oGlCqXJaOQfVFt7wn9y8
C1Y3MC45FxCojayEUYNQeqfxKXFqVlckBPWYTT7LB8hY/k+TvoCehjwzHgUQ
NtHslua1Btb2o6KcmrSlj26SDBYrJrtL/4lfUKY1iJn3p7V6scN1IgQwNV1F
uaksxxV2VSkcmCtki9BqRHo4r4gExOnrkjTJV3qeeYT+H5seZwx9xQm6fQ1/
vb/tXdgdiYQhBi3/b5yLd9L+ZadSDI8im19PKN1cZyrb2ew3b21j1PM/2YZg
R1ZpY22EIviS2MJ6QqTm6q2m3Dvpbp9y1OI98S0szWoDUshqNjdlCc/wqkHq
Hrb5lSdKk1ji/Z2gru2oJ+ZAkeOFLf3nBQ8TFOzD0c4dVz7djkYjyw0m7lXl
5AcyfwAS51KyCK3cAPcFzfRl7fxIInu2BQo+ZtLgEuSaXAUgFPSkpO2Nxhz5
86SLuxgi15WE2wh8f6KiVRIvV206l07rM2W9SO7r2VRQzqt7nZQpgiJFHKlS
IazHQ9hR86B8yTzYtpwOcUJ/ShPyx3ojT82AAopVhpfl51+9KCreb5efVIPN
xBYel9ZIlbk4bUfbKnseYJBlBmK6q4qfyvlSdm8fzySchjtBSdf5/hJgCFIK
o2B8VjA494Ewf6btmj/54KU+ncLPIDY64yofYe9Z12LS4FG32ZEmEGHUphh7
JOfQ2KYI4Grfnxbq1WuFdsssIsXNA29yb7EwGeHWuKlhyZ0K9JP8w8ULey3r
EkECHPNemCxyKILJ49KV+RgCJhjkaIEDxKuKlRtarcoshLOZNpl0br5MhDhh
974rKqUuassj86yPvNHThJvGaBn/D68xNEhLCSayjX6yBSCeL5W3iSuEhdyO
QRAilN6A4CXtvfR9BHvSRFYIVKYVx6iasrI/VZDPB4WQOmHJ/phLlxNcJyzt
RfF++CzhRB3RsipRMgzcRZjkOVU6JERTBbrghR9W8YUjNVepG4Fs8Rp/sS6/
7Iddrbg29+hHjAgg4VnosnWAKQhiObGsB8V2rAER3sSL2FK4aMOlpP97LJsm
OtfK7ADsWsB3P3HJcleduz5VnZFaAwYLf/V4ZiPH+/qV+mKr4gMXcl+wPY4a
gYtfZK8b0EaN7lSEO6ieLsQlbt3ZGiR5ARIxyM3V2MoKf+kQN0th6/LHp2MZ
K1cFi1a20EaEyXHXTx0plMEJUvJUI446hVuAHPKYu+u7+EArW2aZBxDjzOVx
7utA5tLgO9gJ5kebmH0EAN9UV02DuAv/QEBMesiFb+hOkPPmayWbG0sUPIps
TYTuMbSlEA5DnPZC+dk2djjxANeLLsBnwJ5g/w+vsnMTJgmP83xP6mhqv1bS
JDZP7q7+qKrZpx8oWK8Miy+BbR82K43xAf0WHK4QBw3E24l4hV2kIbF+byb0
bpRMf83bLQf1u/Dlale0MVx4NE3Hc0nMM5cTe4H9nOKqQA9jHG2jvo8SI+/Y
6Q2SINkdSboVvWAIiqwPL72KzwN1EqrmMx/zglHJX9JYRY96CAJImJTOLhIa
bNw206JBlPO0/lzHdiToW8cVPNGZCWVtNDosWVt1pj1e/SquF27Z6R+RZr4C
uOkA1Q3QOypyh8pSd/fwB69mGYy2J3wCpPzgNjC+UC5BE++U+RkwwWVaRnUl
lgRw7wG7W4uzVW/E9med07xwNlziwxK5P9xyt9RG+NT1Sp4JXZaj93SNW2J2
013lJ7ly7+HmIQLsldg0xVT+vSsQKjxC49lYlWq0ysdxW1Jdp2isIvx8ftdw
08z4RX6eyovDiTMxvFelMLHvfaKTeoEAq8AsMjN8JaI2cXuEdQG0uSyPnI8e
UY4j9MhMGMw61ABin8Hx31cTPC5iXUXgF6eeU/04zeyj4fy0b8O2fUl6Hx4f
kkoglNUNmfOp2wbEQAwuiEbp0BpLBOJIRH/PrhBk6rDgWrK66ez+taMjylGy
8I8dZoeIZYsi2XaUWYT/T0ymUULMpxqfRK4GhjtVqixXt0jkg6H33I6+7h/Z
IHZMKXy+RDWt+TlIdwxvZnpm0Hs6nQikRFL7ciezDZPIbs8kPsGh8tJiys1o
88AHyiAOX0DF9WzWauEXSfZkd8H2XMztHkhQ83Cq/6npDI+P6ShJe3jRMYnZ
H1jg3tPFApmbcGjEl+oiKv03SmhbhyA+A5PGM/h4Zl98cW8bcpkTbxLj1M9E
FoqTMrCNX1TY3vI5GqUpxeB8Aa/+r+sX2n3LfETCuPnzwU9ImEnAye3tXDc/
5mVcrp8GCHX6T1sClKVsDdTbRoEwab4o8i+7ECQJFZLT1lokrEIYPyuIFT3N
V3t6BpWvbCFdiR392sounNpLaH/2YNssJ87+qpbBydBRb0Kt2ywyKnDo4UWo
9EeUInutP/Iph618Pb+fUujScWIgUsyjuZv2AXyw8lRR9e6UXYVL7F94KKBs
xPagmwl+uyD9j5uXm8O8CSlIFpRDbHIRw5ThrY0LQGTxU3Wfhme5eJbO1Vdl
rQv8Z4xGdKDQnE9PaK/2l2BBrOTfoLdZ7FRdbSE7hIgb8S3/aCsDmCrSzwqe
hbbg4tOtzcFymGQZ+UgYIWgtfUCebSGDv2eF5CptV0u2JkFl8+eVsqhpXK7o
ExCmbYh1Pp5c4t4k5S/PMz6+u9stTaLbD+TIzhhTpDSx8CebY2r4W4C7Oojo
zOBwXdwa4ZL6SSvdW7JE/5iOvOO1vcwgarseRut2JwKxxcDxK/aOyhEfHdbi
QgVhQcad2QSl3YkqxVtsMzbc6kpScFoAzw0czWpzImPKt+G0xYpImtR6FO9A
1SW3FO2hEE/ylyDkjFe/WxcLQ/IYEmpW1k/7CPt4DLG6BMrfrL2/wqevnaKL
0xCJWLdayNfXEYZ2rWHc+qoINHCipUfx25HeCQ/mqAS04AvD8jAbnK/RnBPO
rQwn9ibJlM2LjirPrEq51D6moTEpEq2eCA3u88ToX/ZYS4w7AP/GcSS1wz/T
9nt8chfNpbmg7egOyYzbD0gcz1QbM6TJeMhgNqBHnmXkzrSDGmLB8ORwXQFz
I1lE2SwMC+8nyQxTLNRCXT1iROZbNwTeeJnFcyGABb7m09ChM36PG1+DwqTS
1jI7fSBFcgAIBFjpUM3TsYPdIYdP6Gh4/lk7krlESn0L8Qdu6el/E03wDpEA
vLwxfurhRmoOJqfAGWF5YB+9qc7jlLi0gvZvaAn9WGDvG4fsChMqDDSIHTdX
YtMxPoSw7mgszbGwlcwBIS+QxCSTTcWUtrfbfPiIE+mEFEBcAG13Iq80C4+N
TpLKE20zK3FQmnEXynKSxTj3jK2Q1QQD5MYaSp1aQv87qtSUwF6m7doYtXcq
TXrTayK++DBDlyWlD/sDtB1WmWI6LB8yeUAxA8sOx5Yu7c260yqG4AsrCnBY
+oCnH6Cin/J0jp609qsIt4vnuiV2Ruwa6znM0n8DTNOrLlAoirxeLvcnQNel
GicpJzKmiXeZ+4iGcRE2czpqwYuwj3vIgu4dmc/kesmWp5AbCJJcjH17Pqo+
p90g14wF4Wsb538l02TH9xbYAXeuLENCORispz4cEUwx59g3W9F5voTKPk3K
hgX11kWieqUao5hQIos3ikVK1LlB7ZmXAH/Uduo+bKt1gB9A83N7i0DGrTWb
vIoMZXoycgrYpO1LeOXuG7+nWAKTxCQA6qkRiOjNGC8Ro3qBGJVpmdA8xWzy
HQmaEkHJV4ArM5n5irksvZJtGDptmt4+bIj5Wa9LKHyV6cqhPXrkSI7ag4BW
tNo7NoWZhA0Kn8IlCY75u8kXsnyIHxFvhDCmBGXw3qTgeVIr4jYm16Uxz+zV
POf3WGrqc8LT1Ev2N5+y/lw2jx8RgkBHrxnXDdaDqxb2xX/XowBzAEa35I01
qfCDrHzQvIxGQN7Yz1qVdwpeyLtdAJDQSjc/8D385aRFlqy3HGCMAjg0iU8x
MEUg9coI7vJVuGcgExMlciqtBgTRNEeBZVw0a/r8UOPEfxFKGReBoxonIrOq
kfAS0FJssmtBr+UcuEiGTDsiSmwh5PvHW4pc8ZhE9Tt3w66hE0YjFak+riOa
1BKYOQ3iv4iNs9biz/LwWg5DJc7Dg1uV0PwG6X4t6ZngNqAP6a2w0va22BSC
aXhezPma6KoKyAJL3TlD+bO/7jaVPJtIX5r/AZY9zn5ZehXaWonVkTO6n+3Q
KvSr49Y1s9VoIz+FxSpWtEyXtW9icyw+40sZANyogca+Yw3oj0EqBgmyIHOT
4BjuaBdfL3EsQpB0LJoo/vfnKmN254RQP1CEqcClvCI0IcSNbDY5Hv9vOIj8
adWsBp8dWuV9lfK4lZcDX+aW8K+SLvSP6nuPGBgjhLIdFgCzYW6xbWWUzT8i
zlXSCldJL31kIvtGD+P/jqtSESBt1BrnyevFg5cCnv6WGJVaippod2PntbZj
U4CDXucTHCxcqdEy/AQrhahI+7Xk8w+7jmRi8j7r2zqZk2nbHCB1EExnkYq7
TwyxL9Pa/4ov85EOPtU2T3Qpgu+9NuDuQuDouRa9SHWuri+C60o7Jywkd4Fz
IsTq9TySpn5dMZL0buJnHxcouOvuehv9U+RR2m3u20S1cltlyUpt3lbkk1RB
LwUnr0N7OEMfc0pYAsFyntX91dXALp00rgT63Oe5f7xQeRrerrgpq9lL+MUB
LvrL+Gi9bA92NKLkNtj6YmysxBqP1VNkUcU5MAjuMBPiwEH5/wkYYRhomHp4
17Mb31AI21S6bPqIWfmcySuaXFa4DEYJUiGYxgsefbGGxp5w6GnldS/rlOWn
5QCTnio7z2m3/3rB3BzuzTUwpzQsw1T7oNBcfqmWvUVwn2Hb4b4sVhG4U+i2
fQfknR9rqG3O3bjy5pWBlmFNXB5j7bT187+qphYqEriDvvM3dcXmZMHL++RV
eDwE/hdhmOLfBskgld5dpAsluB+T8epZdX5O9lqB9wYk1C7l4ismqNQ+mYOr
42pH3ljudWTLDwgQKHvkpj+5Y1uhGbzA1IyMcicv+eEyFaC/kdgzp9w08Fqk
D3rsGS+qU1Nz3oxz5xhCfygLqY7pAR5iUfzt+8UougRbNBMiX6P1ehpWMYW5
3RrTWRT8UpjCGlYb0g+iJShIcnabxz2gOSuGoM4F4o2nT5pPCvXUdlaohtfg
lFPn8dI7vadR5DHO+ptSkMiHabT6EmEnbS6YVKmel7MgDwDJNadthj4n+NDv
OKzwMPvFbRlGe4jrpEmmX4STkpCndL+Oh7FuLDWXtYozSN1L540ZAzvmp9mT
VUPWiZoqgfBP/alFe8zbzUUOXlELfpZqZr/o3gJPbQIup96/8sM/UZm+oult
1CMqobkRT1TvCrJfFSlg8bfEzNjEqppG+evt1Wkj7Kb3rO3us4+dEuajwymq
a7klWTLYo4gNVs2IvjW4G0Vk8Y4lVub5/n3P7eQrbLbViPiz0dEs0qFZQt8v
uu1U3GqB+cLuGdXKQ/MpnlXFe3kAGNtA2d7366WSxQE19Jyhn+5fQG9P8Ek+
6jL8xmx42ohwe8WGYvMHq+nt7OIaRA7hwhAKiBlJA9CtlSdhJJ3NxydCU2g6
su/dWLd/7CsZC+4cR7e9cSf5j+O1k8vrcmJp5K175i62ZEnsC3xJNp/VZpaj
SB5X5i9BFVTdfMMITO3Zml3C0Y/nm82zQb9yIL1JJNgLpkiADxk0qF0BUInU
f+/pZont6sU5eT65d3n2U+iYZlKrNGvfq3QpfW1eB5hwrJ13LcAWHSIIDh64
hICeS0ifA5hztUMEKgt0FTYT+mKHp7+iteoB+/4/R7AuGMXLO5IWAyrc5sfy
s40o8HrRbb1u63mcM4D3jxGbLdMOjCSScmH7MC2DyWg4XDOxdl70H7MwSP/o
uAyKejh4a3PKcMtU4b+qnNuf6MVilvK7nbfcSYJMCTozfyIF8gCnnqBDVS1q
HYCRJjUVTYNHUdmJnln4wtYArLj25XaS50dcD6WnkYmnA1QtZfHqomf9e7CS
TAHRy42UIcI+X+hkxfnJM8cjuPaHUDkqzS15eh8MqK+OMOalz/3Axpy7ZZZV
96WWY5I0zrUpMeFpE/8U74e0xbGA5GBal5fay0/7B9pgFwvZWz8Yz153cHdg
Kvg8JS84z2qSKygmtoBtm3/TfEU9sqdv9ZT4EiMnH0/PBvAfYwddnTRfipG/
fobTuuHG9SLaOW/2yYz83FOql5rP1HcnWBfN9QSJ0MxZUrtEJiuMtoxfMRbJ
rhtJXe3pJb2nFtgFCrc/0m8hAX6fHghlMXA+ETxHcACVtuW6SQgjpmdUyUth
uwQ0yxjgZoFq0A65BqiKvXUYKzQ2mG6RfG0lZy9tQ6HBhdNZsL+ovkfUn3P4
9Ja9+BQkW0f35FKqjVjx0aUu4WpjzNv+4wMZstgCktXQZ2MJ7JMQrhl1P/8C
kweMfVPenH/KRgkgL9RXKzChIIsdExQc/r/hlKUDihwPd9FvGwyzhTswT0V1
6QuBKWX0nitRQsCHzCMDQZLuKhSXeoNO+BkNw2cdn7OrTtYOmZG+6b3ZJ557
aowvkiQEhfz1CAT6syY9+M7x84IfIzYlCE3rexNFtF3uXwXJn9/fmtAKHMq0
rV7UBlXL/ts/Zyg7fmH/F5qMGcOLUrkLjRAXN0xncEqSvWV1n4E2+ttJdgXE
BsSYojICS91/JQd3QquCfUAzFSlZTVi6VYNbiz4e0u6qb3XP9d+KscgmDsqD
flcFIe07ppsYF33HYGSTrAS8hgYp6s9uW8Waahkmv0wQvqaFfkKv1Pzsdmlf
vH1fEN+C2MmEmkVp55dBTVpt70SzoQZ8vOhDEVK4uOgInp0n/rbeBeBCkas2
5+JcVw2ui5EaOaqR40hSmBsAv1GcxlIOEFv/OlK2LhxZZ2cmH3sudFvo/ER9
aB2JIENBSqmttfasXNX6aYUG5SsdXmws8f3Groy723cBuNcWvSMrvraMd9a8
IB7ZyCUOb44dtvsvjh5VJFoJePm5STz2FlGQfK54XNwp3Zl8nOtlogCoYbsj
9O1HQiK6/5xvfkhsd/qo0A89ooCWy02mjU6B0lIoZluNvCDLQfzuke1i9Cxk
2Lf6d9owBHSBPmtzPnXaoyLy3ZCjCnYNAVUd2GXEvpq4swrG/IAWb5gZ388J
E7W9m+bXRj6N+NL7QMfHZce3ql8iwHj7pKtlNNIGf6wVHhcn5W4V+/wrO3cW
PuJ0XwhL/gaM0yPjc9XoiJrk6g7vb5SoHEd44zz8757QH4y/S6iZd/5svnjc
84hl5UuBIojSiOt04jpaeZ6qxL0ND/+SFB2Yo0rp46f3hgZC30kyluGLyPfT
rnk+Yyyfc5sYANCd5DHTmcqWGATirmZmpM7ghcHzDKbIhOh4qp9reXwr4gTb
yTVltWIbdagwVquwQQMQ+/MpVjq6IlKOD4P040x1PideemgFzbvlUk6H0zSN
itQDH63CNKJX/BlRdicTqJf0zZVm431VZrgkamM2yqVqhvZQokLvkUCVaYf7
Q1NgNVgEG1MkMy6pMrpjJny4+o1hNwHkwV45BJYbGNeOiqmFmWMGHDp9xkPw
rE2DzZM0BoZyxAEKxVUrlNlH3OJA3qT9RzbOEAejD5OI7/SrQL12BVLMTmLU
g+3kGabDzfYuyw9wy9AArUxuMjSdLaQRkl8bH/5bjFUH/LviOIg5kvvzX7wu
TzeNjZwfENRnfgmh+oCpMnogXpZXZp0iyq91Gnd2TV5IYJXSFbjnODNCJyb2
VN39N+3C60l+8bByQovkQoytkOLIXYmK8KhElwjmtgrSDET99n5rqhbxYt0X
ThdYPI1mIfUaZjmQfRrsccJ5dPaskJxpGGQED0h65zrpTPFC2Ydoe/G5fsh6
LzNM9TA9WLnzeqeS8qx0LcZ2MGN11Q+9yBu6kUrV2xNfLeh1SuE3Pre0P/t0
vFxVXQMwUDrMSL1c+APBX5ssNM1PL0nnYUk4wt7zEtcEBEQy8B5m0r3b4ia9
AxdykqXguSSJlRANQC1MNumZ+xd263fdZyOJivhY6z2hGKk39uAhe0Rug15e
Ox9b6BDp+8XKBGM7Mc04WALtl17YEO6YmKzaSmhnSiSek4JovbEeeF8kT5fo
LbQeqrVIDodqMqYrj3HKahxzOpeEDjCAFk6A0ltL2RFNhJKs9cXNBeiRgHDe
e0DIhylMGTMIxM7/o1Mb7MKIs6yAxWmDDnAc5QarxzfnFGAs+mzCiRQ5RvIX
svrKYwUUVqfkyh+0ZWHSaqHqkfFXcGt/2NicnJT9p+qARvgmgJltSMaWoduS
ku/s+UC1GUFVNefGoe8Ug+ObovRqLtmO1VdhtCzp8N3ozDnqDqUttTHXHHTh
FbtfaI+zAJnTK7ZYbcMm+OOgPRE+x4ieJXXyW66Cs0jKA44CsbD6Rn7H9iRb
+9q/o8/QlFVYlb/2hv9HlMklFkPRI5FUKRkrOivLeBONhcrE+aNCdNhlVkh0
52755dKn1/AnohOM6huaj82oCP9qas5YcbAjfZiAThlkuGucxLCheeAkzfTz
0EtuDhNZOFdgt1rKCKue1QfCev7cz6yrmSvrJOvUqTULk2jyNC2FyH3W5Je/
2+6zTxyi+7UMnKjIWU1pgdw1bWSSg9qRc2aqICsoJyajaSEbEHhx0GkIyP1y
L0aUvjDeihNuB8TPcHlJ/EvDZZUyPAyHx9YXvmXPA1KpzQwtEBbwkbNamcF0
aREc/18ryU7BVHg8GcPpQqqdHyQ5V92m7MtGSi5fnwwlx5rM4vV5sctlppXe
yURfw87wlleodCkh9jGvqqpSDnrsmfr1yihq7nPzX48YxrR6R7ft5qONltSX
LZML1mykx1lJi1i64TjswAlB3ak8UI9ko8JgMJHJZZGvmv59S8k8pb8HNBFn
kKrjO6KmxGy/L9B3JgxW0auYD9Y/+Bdf1jnc627U4oT0y7EM8277QkVKJy7T
nGzX6P8od8wxiCPUJJ+bVp/k3fGzZzEAgsMpjXRw8L8CJHxCB4l2AxLu58q5
pMIKhn97zPdbwY1XnStxmEm1FUxgIhpWZAOLllSooKcbFdM9jvjEjXTWruKI
fgjKbAzRADNqo34S2qSeRXtx02+qWi1ic8j75etGPyfJR1FyCd+QWYadqIXO
27UAVxtVTLBk1YdginjOMPzec2dCYQ8C4t9Y4TVAnumNvnEM376H8NBp5/sx
H5KoikchUK63UWV5cJEdbCGPBX9vJgqDtzAfvflWDrfgKo/C4YTuoRy9X0PM
0tlRid50mS0oeEb7+tz7XBqRHO9rLj/1GmA37pVyN3fJFA09bln91Lc0P7q0
ywAiYFiHDI3O2F3msxTTyl6dXQYzxr9U5/VByjZQ7nAu51hfOUKHsfphxN05
EI/altDvfgc8zbBfoGqLynhYBb279CaHzxBqjN9rd0SMz6H0lw8I+dQKoukr
Yogb2CsFtx8UoYKvBBZL3AJApBgCdZnaH05yto6SGhHTpkESJzCaQoRkpkWC
3k3BGdN0ZdNJM9HthIKlSK+17JRGFjGEA1i+dmHAaRWI2OBeG9B8qwJvYUE9
vTAVWSo21anT09tqn2U/IMsoUJDo0YXEWNCOA5EuBZx4CtoFVtaht7GKYmfj
3sqq9RN1Q4roqTlIwnpxdCW1wGdEKBTJHJ2DeuO5q+wGQd73PGi8JC3XN2wq
pdNf7r2JanpN7FOEJ1xOAVE03Qv693vYTEhv6LLLKY80ckCpRiV3BezinXJu
Z9J5kh1PdV8GeqSqj4NXoaYSmkO4K93Xmnw/NBEGaqaQ45cWtf2GcN4YORyf
R4CPS7rmVUnbDvsxSdkbZKOvc8No+dssKWh2YVbAtoaovYYhG2K2oZAbcDYA
hrp4C3yG1uoyRcwEw4hQOl3W1Bw+c3qkr6baNkkttdBcYGQRI8jLJpkfIBSn
lUlHjlWv8cBDi1fUBXEdYfzn4CiazChrNP1xrHhSJzLMZJ3NKvmjV/BJ8Mqk
wdqTN3S+qnT8hcpXMRTyHzZ0tLaF5RHowHxCQnjwydEq2/h9T3TQuNTpsLcN
MOBk93wx1ZykH0c6uVvTtbEsnxkJGK4KrERAwJaQUM/Ia3ENCIJFMYxkQqzs
0KI+QAoZ0KI3TMxsrCJYv1h/BrN6btcGbaPUJo8WMwpCycnsYPq7LAdD0yQR
wSfRufP3kbWfiNV11Ww8eactgWxUp7VcSVu7X49w82OFCKZDQzLQ6lbF12b8
C5AUO/yGJOJfY8/JTQlKAwDC1R3i2EVv1B3txTI+B/XOGZonDYKL51PZT77H
onLdcKCIFn667N/p5ra8INLIzffinwOltl0BKgxWN5DdCU1REgDJZsymIDgS
lAcKePM3XE/mTl9QitktD3rv8Y0uoDNDcTrDttgqHHbptmaDh+UJIv6/1dkF
Rdi8ze5pDNK+dCOCKO4qdS7sPLV4zKcdmubL2CgiwUdY4SJMdrrIysaHO8xc
MN220dHmOxyYhx/+rDaly80gI/RHno7WIeRlJgOZRX4W37Crh0pbbiD2TQNC
cizYgmCq8OR4LZy98sI3LFlwEYwmCynAvoxYqbS0kjdGKBlse0VPeQzqa+yl
RtjE0cOxKoc0jNYoZuTwfqw7kT/eGA9E7m5U5JwNzTeOo8G0p8BsIkY42YHv
BhtrRwuh5B62IT0T7+H6MBVzNsd0lQuOG4Y5iJNJggyupNspyVwhpLQaEXmX
tqZ0POxxunca55mjSuA1uzVT/fH9/bx1KWO5lpVKyRQkZ+bEZ+lTDfZpR3gF
EpsyAqU/lhjfgmovupx4NSNusVJJveBfVufZrB+PNAbkTU4sNmhCl0ubH12b
zg9Ln9BD1G+DxV2snRoSnmybjGfEtwNS51TuTd4BJ4OJ5ZFGfVtgIUF3y3v9
ugKDndqf7zpolL3uMFdyMEuK8b8agt4uFynVPk/btCgzC5CDayQp9sSHKTVr
PPhlBeUhbCf5ixXnoMdMzbEuQ+pPddWv+s1x/5E8KR2rrD9To/emU7iewlxv
J2Ve9SG4Swg8b/TCBW8hQSBsToYmbDGh2ExQ9UP4yQ4YIGkKLCMWOoVCbDpR
XhmYle+A1/eT38ni+ZXP/c9A1cFeVxVdQTqtodsQxwtm2E6D6Pf8/aaOoV9O
Gzdw2l6LGwXyme5THFuA4/dhlr1pCM8P2bkP81sQy+03WJMJDz83w55NyDzc
e7oq6xYY62ShfKUUfzw0gj0XdlqnR1AH0QVFQQ8CS/ay7NUSAImgSVDAbah0
6Flw9kdsFUwBwnAc1OqTo1JsV+X0rzBHYTjg7JfqZfWhKoQZsBwOLs0zPK06
Xes94e54r/Azd1klpinWtZ/yM0/yplNCbl68NxG/b6RKldyzPS6Y8XVTvipQ
/1pY9cdq4NPsSVtV8oGIA8LKT+F3gIY3tVM3IgXZXNKPIqJbzFhbb7J2cz53
S2cfx9OpMng3O0HbNeDw0jeOI8bvBs+mr0nSFCdc9OVmYCCw5Eiok7pqibD+
q88gvD1uizX6vg4voa0tyst6hWyTK0xTkge6sFS3BG23Ra/39W2t8bUXy7//
Ml0qXIohaZYML0cdktWeTSSliXJrhNftvlp+sL4Y9+g6xjVMCFRtttI4MCcP
y2oClLQ0KH+GtxNCUs0AIeiuzTc2YExFEF1jvWNSKp4Y8nPUYgMFKfWO6CBP
lNbytS2y/zQTIDnUhLUrL5KEIh9Ylooz2VTecYlWv6AACWUwSmY8QuKy2Wwo
gPmMSkUsoQlxfTgFZwK7d8XzE3eXyVYvdX74ABMs7ZgWiW0GVmcocJZExjFv
iVnusclBqUquG3qQdh57HGl4a/AbfdKNs16piBzYLDhyMrOBjp+CTklnX1W7
kYHF2Yd+pXQhgkR1vuy71QFw74uAonkt8cya5EcZLu59zLv3alDfteCNSxXv
EVSmJq0aivAuTFlT/3mqAtuCM5AIdgoXBNnQwAwgGrDWNFbjnXQCjqKFtSsq
okrqEQ+E5rUpqJaulWoHNeV90FaxwU1SiF0yBE3NODm4paNbLLmOjb8sEEqd
Foqsqz3x/D4pTzaYjYdxG2xAzBbYt20Sp9RnQEa7iEoKKYjWIH/UuJwuV9xM
gxVihai54R0uV0ygfnMBiSztrpC6h3Yrl/wV0qC8Sl7JjXiPQC5efF6XvATk
7HIrKgROxoQo+vA9Syj0X3UWUhesVtMu9WtY7fSTrznHwWhsneU6XXtCQTHc
afhzeGQobMl3bZOij3xz27WMjrvigImfqqFVN+h89mJKGfN251n2+7hA7Nu7
RAL4LRtDtcdrGMQF+ZNSG/nlZZCR7zfbtJylSk8y454IjHH1SdnOfA6evF/A
kNTEH9QgAdvxU8LK85GoaatX2zTJvyJEVGWyosovYV69OkJ+0OizXu8rvrQ8
2EKf1T6gg5/O/dy6FBUNMS2gyu/OWr3WrDX0i81jObjG+ICzYpuyqKhm/2IH
94asfXBp5BCjbBgC+gV9M7aSwsWVwqwwZta9asbYwlJbLI13PEUXT+RrISHx
KAtnKOc3T0s2Z09rxCn7GsKsPdWFRJjtXGhKZu+MgsuWszruUzdEr5adZAuw
IJm/P4yQpmKRFN8rARRRN4j42BNypypk9m8XdW338Fg9PWW0hq0s03+gevmf
YqwTVwFuZ88cEQ9uAOH32HbK4XeS+P1igr/GoaW0UJ5fTHS/9OAVvcnXc9Qu
pKENXG5rb2fpYxwjFQpt64Fd0REblmI9XZSpwruYxCrSiOCah1CkxzVfNK4z
lMsR0FAvLUtWElyKZ4oW0q8CiODFUKr88n7bgdAPv90AXZhtdQ0gEA9zso0e
Bkv30ul1JB+LN7Xd9KxZ9AyllcJAO+YgcJtKIouT0DJsNLxOUfSGGhTJ9cXO
/vHqvVEDcxk99jdpgwLHnXzj74hZykCB8Pgqj575QaMykOtW1CqpwNU+cdhZ
yWkYCW6H76XhdAw5kq3hn8SixKu4UGOUOB+0eOqNsMsyAqy9awFWYLMdF4BX
0jHQwQnHlO4o5og4MFmw+7Vncttc4+BpcJEgUPASlkRjm5YRAm2ZUlJh4GMc
Onj+y/iGb3zU7kQBWSYF2MOmf5N0WjRl6x3n6W23vQJrpQuYLkQIQPHT/R7Y
xy00/aiJm6Dm+mofLw8MttMcVXrnIblqMK7p/W71oCUsulSff4t9s3vmVz87
ofZHsegaM1p3SkD8BP7QMBK36ffwPm947l7O5KDjnd/US6yDFpuJauPvLcxt
IxkGnj3Cl8i3vIFhpR7GqrLBaQiIbyQLU6d/b0d6Kni5ug1L2qjg+6GIh4dt
uvVB7VQz9oL9I6apEkMz8TauK3mhm8Zx+cb669+bY184ji7ivXLsJ89vQDJW
XVs0lc8nL6de1s8aCqdbfc2u2drIq3oTZtSfxLlI7JoyRxcn5g/ygTgiWqNE
FIFTdkM+s8FX39Pc18j+1CCbBLuXiE2sbbDiA0V0Vw0dmfdZeBt6E8WmFA39
WgWQTxACP/1pfDLOYMZUIISEMU+0LR5yvR/Ki0Uz8Hg+cFnXFl8Xvk1skAGp
Bgbw5iFOzFJpNRHqX6IJp4AgVI0yZOKkYswnWRwXxHQfMycmTRrp6oZrRJ/Z
9shkVobhG9lXoX/Wpi5EbEsAa8oXTq/c7AnYexgLD+UQEDe2sdA6rTPQ8xDp
HXL9AyNLhN7Jq5ew/HRt5iF4IB+flkOdyZT77+LE9QPLiM9PsAV46ldLwoxL
8zI9tfbYYG+JCrt9dWWCJqEFBNe8ElcN12o2P6qotPahbZj5b9C2jgmsIyuB
vvLt0Q1onRarkSqCv9O/s/tWnstkuanGceYd8LwfYlLY3qGIhnRhS20dozbe
NKclJLm33cUgmxSI0gmF1jfDgKEG/XkW/uJfVqbUIoyYVMMyDdoUp2KOfJ2j
SuBmhxTf59CADQIpElHs8PXdU8L++MRerzwOyfL2iTTyGCvexKMU83NvFvoM
IhM7G+AaeVxiWP+mveurAzlhQSeKK/0Hmo4vh48o8JCxfdLzXKfatrQbMKHN
lIBc1QqBhzeuvOK44rwklAcCi0mED6EzGfuCQC68rwqpZmaWZQSI6rj/zsVE
rD9SpY/Kf7D1LhjGw/v+ZIxP56OncumCErcVZ6DDtjwRFCqeh/ULvoQOHi//
dBHSLJpUPCsJYpoZIDL9X4uOSUByAUe+X+Ru+n6MIL8UX4iRGTsshrQ6FMh+
EiTvsQOeQ+TOfCQlefrkO6xYXkToRhXlMZcVzTkCLQ+13R4kkBicWQEHNxeg
vID7eZ4RiCVCJEpCBz8QesE2HFZN2VC54y7SfRwvL8QcQMHeARaU7olysBH4
tMF3RhD+vzF/aAFN956HtJzvFFw0At3KW2qjuNK6i72bwM2KRsRCjPQlIq+j
nom6Rru5GZIE/278zybO0JNwFWTqTpAVB5Ea1m9i2ZqzZauLty1ypsFOpWKt
n1Mbpdbto967rP9vvZ8QAhOpYcCN5ye6d2g2FZUY3gggTljTZ+yyq4vYRWOI
TbosLagJOnbu1vnqkFfSqJ8F15au094f3z227VZVPYTJyduIE1iiilsF+rvp
6R+bTZVD5rIo1NeUqxPBYqD5OqmLvcJZjZNIcDbM7ljgDc/pH8Y/IhKLJodf
i+gr6UG6+Rp3XNwFE6WphJ+i6ri/DlJIa/3gg05ESleJ6l/jYIHstqAS03Er
6YJijhXJE3nYubhYXvHuNt2NR7/w9oqpSBfe+boA4r7Tkc8pArHzwM+jIItf
U8oBUrmYKauJPs8L/D0jFltgrod6GSiIX0tpr+ntYIQSQWfgWukx7PyQjNlx
ECePk8V05RqnYuybOGFTR7nLUQX+uBIViWEtt/VXm7bx8zW9+c7CyK81bKyJ
6yy4xwU+dQa+AhXbIdtTqY/G4OhJhrobFj43WB3LU4X2cmMvTCzaq1iDcXxx
xd0nSFgS2wr164Rd47fEfjpipMTpSv5g7OjGKBvyge06WnBXumR0Z1z+O74p
2LxuSMS7UuBBHPPDe6oyE/QVmDRHRFrNcDR6wcFliQKNcYCYA3Ue1CD565MB
V6o4MaawFYmEv0oVUekZ6WwhWjy46On1YKXC1n4MTH828adaeTKfEpVF4x/E
2+1PblgdHYvaebEhl8b1h6DZcnmz26h0Or6V/lFBQ4Y4hUj6N13zPI8y6nSJ
smPTv9Xi/CGbpzBds8mtWli4yUZQvWA5HmFYnC3b9XHCAxoewmVjUn5ZYLBX
DACFCuC27U0hxuIeidCaWce1m4Eq1Qfq/OgC4FoQgR3+YfINWKSwrSknZ6Fz
9idNa6Lbf9x7q2zM8Q2xrBId6VkVabYkaO4O3HxVrzOSIxY1W1xmpEsMXG9L
WXxP+4w+5K0MPhcoKyeCu03F7VAr22gpY/aNZ3sLWe/HwtCKKskFrG+tYJ62
g1kjRuQheMZbWhWUhKGIhfeoY4XJk92A1Rhc0kgR7Ip568AoyoOxg961j7UB
28iA4XgJgDJqsoWND8J/Q8csUW4Ql6TNlWj9CP3sT0OukntkuLGFNlJetRgm
IGGM/O0qI3L1etvdmYU4XpvmtG00GtoSgWDVEQV/8lhrhCs36xGOa8uI8sT5
K7Jz/IHEc6Ly+GjDTgrfmbwVPUcb+/KHzGpWh0/5aQRr0C5IbP1lgEiWYzzz
OYuNh2doN4cyj7AGQoRCpLHWt96cTb9gDQH5C6iSIzXicsskD1SoS91Yp/yL
t7Rrha4p07JPT4QBdr62/8UtlyQfq3QjJGgfw4O4zKloV3HmYQELLZv+qTBW
oQWb55uoofc1XnpbyPht7n2xZTz6A5Dm62TloqtA0oArpWxrZlEPZgrgRgqH
jvj+bVMI2/VRn3VHKhdzcOqRIIECL2VPrgnZCQungvIYHTMQIkq3NiPfzTSx
8V2Utb/DGv2CpG2bhAFbb1uowdl41135CaA+SXrWVhQLNaRE8qkhlT6U5ss1
36CJLphovzm2zbnGjo9oZ0JA0vckfVPoQpdV1c2MgJYxjuaIwwnSkkin0izL
rHINHroNo//Jp1Kx4V9H5PoJS+QGrC5rqJTtyLYKCf/FLl5h9xnprRvED82/
bmAVbZlNlhMzRxVu7BRj82YpQ9UL4OdLnbQvVQ9NdEkMz6bVkbzAsc26q4in
VOpXTeDTo/0+Etaj2PWXMEU8I1D4x2vODNpK7HkbssMPpixr18JPcbK7kHnQ
H9nfPyVJqnyZtGEtDz5hxSCAU9xw6XHzvBL/Aiki574lrfs3etLkWci++Kow
uaEhHmTCdMl9JZuHEm0x3/yHiwaahI3Xd8nofG+qHZEP7YiQy+2FWsVK/Ugg
ERCZpTvN2C/e0lfFHbcu+tvH5pGZW9XfdUd6AJQwlhdkYlp6M0xmLylKV1JV
3lYLCKHnanSTOjNDmhn34eL1/NKBLtleeF+tHvCfLhUeJknXW34HRGUVdRG/
8gSQGizyqosRfh5w/GQI+6eB8kGAcH9Y823RQXGTpQCrLx/m493Y2DsS33IH
j8/W2+98DKzpXfVVKaRM8vkvAOXwxYtpGEZ9RrulXzett2sR7+43aDi9I2CT
vt+31RCozp1OSaG2Cl5IJBFqEANfMc9+dZ6bdFiXKdVwkAo/fVODJ94OyjwH
wA0/NVwQxZ/hrFh5/CVmX150G4PL/x1ysx52VlgrIQPamn8Fw1TB0zs4UZ0U
xiEQdH4pJtG/+773l0k4nBDXKCY+DUZGf5KD8AxdEAlyjzoEe6KefeSnSOX+
QB909SJroU6e6yYPvP9CzF6fQlgUagTMCU1eKQhGEgf9u4G9j+3j0mb6HI3O
+OpI39vkkcw0KlNOJxjgvZOhQ6w6A3CcEsfk39qnONrMxzOWrkR2gKs0ekvP
znayOnw6liJ9bFydI3wnwt9lDuX8NkHaIshvTK7grGf0O9DErPtABRle2OD4
bBqPOwGSu/FR0WYOZT7fwTJO0kYWifl/4rwrJdPb/iL13Ah2kf4BHKqZyjLl
xkbwtbf1RCKA9l2eL7tO1Mv0hMWdSxqFtA1rNtNkWNMpW99zhwBU0i2+GLdD
+3Ut/y4NFRqyCLHpdx0j2jymIPRcAcyTtfaplOo+TVpX0nLy6M45PTEGP57q
Mfgm0w73VcQGID/hz/yLW/kCJgWhayePjGScJG4vr5BTxOo+WbRHg4qDlHZi
N0akocGVqEjtG4YXOJsXQMWTfqFFo8+wxbJYqnUmeblcKzk588IeFoGOfxHQ
hWaT15Mmda0Pep1qQ4SRVeuCr7K6zG8qzdZduJr39USdTWiUsKGScVTVE9Ka
yNulKS0vxp6SIDCpAOgatEmfZGyLVhfmDNcqGXqeFjStEV1PBTkznTUxTYKj
uXwkzXLEumV/WptyYhvIlJ/K/mFf8xtOQzeXSXxsO0lkcCZmsr1wesD068H5
qXNmX2FkZEw6S7tLgwuYtSSX49s471UsXT+8xrk60QL2xnRNfmPHglRbF6fA
+oS+wXic7Q5LfUmeithInAol7NhkJvoe704286nEAT5DZgeAYkodD7NAzlgs
q7X7tybqOnpODNojtMICNhp/3RJRrB1m9OxCIPENN54OtmKChY1ND7pniSXA
dIDnBmS+yVDjJoJLm9KDsVZuPWjQAElFz2bpxtpKLJFakV8OSPNziPiyXFX0
FDzzBkrXQVg2//Jq2kmlGn0mA86VFld7afbcjqNQqHAnNEDNDbyoDutQ+p6B
63IqXLqNnye4jqLSI/o6m55QEvKn2cbryv2uIUm31C4trj2/XIIWCUpmWnE4
nqRXFwJRb4rSzxp8GMaozIW1Zn+C8Ojg3v0CxQTLmSJjmYFR/zL2l4JA6Hr5
ViaiJNNWGVAYXpoG24H1eIWXOaKxyBZJe1zwOJx1C65gymDmtRIkNKXFjwf5
ImccdvLBCOTmtNmh5vHk8YJjMXMxYMGOA+DHIBoED6yaoeNitjx1UJVovW8Y
XRrfhCPowD2KYZ8g1R0DXETf7KkGKx+GZ50ui9cDaneE7IL8vYnLuTw9X59x
d8ULZQHL5Q1Rbk4AAk3oN2idNQhMUPVWt3fWDHl87jDguX581YC+72WyFKpE
hcKf4UL2uPLbmABq1y+e4JdInP1VAoOnUUcdRYmAnlGdQ2/62geh8kot9HYV
7Qr4DoEBq4YHvFFdknwnWOeY/YEpAbM+aOl9ek4WFRZ/47uIU1sCQ2Kv02Kh
Or9rj8qjkx/XAMsiR+LR/hW01SR4RJGFgN3Tzfnv79NljZdSx0H7L9nfPrWw
v8grNBtxDbzSfvd/Os9iYKaJYXbCVkMFMYlrwlkwbV1bvXFFCa8PB++RBcvk
OCuD1QF1es835QSLkBvuTFqt32znhNnr2xHuvz00tNnO8FkAzAY79T+199GG
muENGAS//XJXYvPyfDLBTYquNiJ4sdAM7ZLw04sDO0V4T04WxDl9B1IbG14w
Bvky2pCayA14oA+YeKHbCK9d0cMtK8nIjZQ0sCAMXEmiGnLhN8C58TTdk2uR
0czUYj3AdbIL5uoDT9uLv+7FPQEYY6EtDY5HZmjVbYYaDB2qypbx73Jaylup
rpscxxWCBp6b4SpzMa4518pWsTwVvbJ7PTMWyaI57SdjRDTDfhcs3PphirIA
hZr/brXrVgeM6MUEcqs6w7xoxPwV6CFByfd9cyLoZNuqgps0Q4sdend4jkR5
69aR8JflOiockQERWM0JySQd+x7N9RSDlVE5lRuazOub7S405zVdDzJqPHTI
YfKevoTLq219qtvDgIJ+w8gIYDQ/4dVteA98be2x42ur1PWD+S8Qk71mkwr2
sL/czbo/1Jc5ZFSHLBnrzM/vZ/bVOt1QA0odj0zL4BPeB0Eb6srG9TB95rC/
aasFNuxJrbR/ABn4s2OHflAlSJ0DaMWvVn48dEdqJGW3exaExRrzUXshqhpG
U+R4w5OsxiuX7U4J9tc4N/di3QW7ou5oZioSKEDPJgEQqgzXQR23vraWFR3M
yd5V9/1Fc0Wwzp+roU/10AZTSxJjd+CvzT+b30HOFLehCCOgLOUCOd3Sz+vI
SlPkueeqmVDBtFL6nMLPdb+QAthUZuURZQKwu0lYK2s6NHjvhNtnSLdjMqAv
IOp5WuKo+BCmSjl6/0WQ8pt3C1MYzWI1DuIjZ3N8kNDHaMX5MsmXrdmpyxhG
e784gAxp291bNgB4K7Nnf8POE4WBDO97MWWXkE0pEurWmPvEc77YOec1vMDu
7su1sNoOV572GmPUz8U1NKYCbGP4RqTTIgUaya6NfCc+cch/x1Rc1sHWlUQZ
8yofOObFdqw8uDeSYSC1LZ5xGHaoRGuV3nsryfkWVBS3no51szmuS/J+IkE+
fqwK+OROEIvPBbHavVycDhne97O5k46XxZWfqEHDhpQtmhrY17cHWZ9ks2ZQ
va0Xv6GrkSFr1uUSQ8pYs/Xugle8VqZDWaIRsQlPxufQqA5wXjsjHHuX6WdD
/7di0X8f1Z7bdZ11J08PGKVPc6k3Oj/yoTRlAWzKfFMX59qyalaEW0yr/8z+
uGAB6RY3440VWr3hFftJTngSmy/1ozRPD3pfAWJtqjqRZ/8kkjr9og5w2oZr
oQ7pCS2y+7rs6pZKPYBBp4iV4BDqxxJSRrv4JSnj6sOZOJPusUpfebhFF0M+
6OWlJu6YaIwuc9wYKc2bIU+8tRmtU+XkL9U1icqunGKbfNIlO+Ld31KVcj0m
PFfK13gpaaH7wQN+3WHeIcT+/hvOlwauTwOUc9kaRZKxjLtu7It6BuKCM/hp
fpbweq61HefzqwlqyroJ0dYOQN3VvdVcBKOzYnoIAxLxUyYWi9rawiP/LW3u
NeOF07LDVpZnq9ljhBMPtQKf3Qu0b+MZp5LtWjEGi2CRpunF/+Mlz90a6E1p
cI04gtlKmC2jOZ8zOETiPbRPLmwdSM58ABYMj3Qg9oAt36u14tzjI5QWcEi6
K6zzL53OpcJEzIhCk6tV/8XD06eFztYc3FZnxH2XCm2XgJdPlpd4m0+Z7ZPg
Adj1xH6LJRd7ccdAWrbuXEvbJhh80/KDq2eElsI8GpgUuCGwTg1FZHzHH4JE
Etl+vcIt1vqhv3X7KZFciuj4YQmIFds6ja5GvtURMTC+m0DDMAgemcn8LWB+
JRe2TWXZ4izvp8Ov5LxePE3tCbzMwgTCdbOwcbd3Y2Z+2TTFCxiqz+6R2br2
Tg4yuLSUk/cXkq8jJN0vqVdUEOdegw76wus4s0AJFTqRbMdN2DY5cbaTO7/l
WRyo/TDHM5D+B37h+5fhX0TxfNCHYZ+SJY+XrdUQi5RNuTPrEkcveknQSMFN
WuhLwLe4EMyAN9BdiMuf6VXIdd3PxKbqbNzyp8RWB/I8JAbPAdHxnp0X/tiN
r/EWcvNb2fNvNxC6OthS3sbL/B8L/xDGnrDuicRMg7xg8Jfb3KGYTwXu0N1I
dFBCTbsN+8R7446caSSidd1rz0bv9jicnZSBn8dr0euZCFcaIWP0VmrijBAL
LpyL50zv6J9FfFFRCs3aaQKQNIoE1fU8lX3GVAZCbjTK322nAScaL9WOG/8x
gbHWHC5iWGvty6l+ZRgLUPAglic4h4tWeQV6r5dqBmANfh/ybZqalS/vD+di
tkLzvoK7Zldd1qzI2uNvxlliRPzC1kVvQ3CBM6PT8uCvoJlUJRf9ZRB2EoZ2
KkuVN6fDAxUSL4BMunBBycYqZc6NDk/GVFybVAkLwr2SQeKHyv1A2SXv0MrP
Ofh0zmmBN0INLemrzePdBe1Hc3KmsWIWLlOy0iO/s5XTP1tWkM6lzggdrruW
Jm8fBj37Eg1zNe0LcPZhmEKN/J9PwFf/o5pt5z0pI6TKL6WnthsqkKcCh48E
5e5neZ5SX3xbwhVvL/K3ER9eoRqnEIh3h11zIkZBOmh666rVm9WT5LmZGonP
iFMCiBEA3r127Jk247tiw0T7dqdWcmG/nrUWmbpv5wCsfa5vh5vMjt3jKuHN
Bfqe5okDQV8WASgel/rnnNRvCx2JB7EVpdx0Xt2rYubfWpWb8i71B5exRmn6
ec2M3IQ1Vwrb6lvEp9w/EWwfW4DbIwSQkCG4McpdlTQ1tVVVJiJd1iTzvtEa
zPvCjHeU2S401FLkXt8QabiaIECmhfjzfbTriW2YTdUsvLHnLx8TtHrojVtT
O6QDzL18kM9rnK8e7/ks5SLvPVRW0ntT8RavotgviCmn1qwk8zAkQ4TjHNol
3k/fp+AcQNXtkK/8xJtzABGKRhp7XEzhRkiIPfvPzYp7ON/tvWThVnXEAohF
qP7Y2bX82cvS6q8+X2Dx2mI1HLhm0waFOFKYOQzS6iCsEOPohEDuqBjSJr0j
DjByodx5hFCcgTn+A4qt6NGf65BCNa42dgRiORtoKFOnXxuwNXqF0gaPTCqn
X6zGM6tNaFuqE8kSHq5ugTvsR5Y2IgRW/I0mQGx5eUhTQEVJPrlc8pG4O9j+
rFTHaF9eku+TUb6MZSEfD1wM7nt5SsyI99saLHSWmw9La8mZF3qYHN/FyN0D
87/NxgNyzf1YclVZ6YmyeAKqsqh6Y0UpPUGv05qTovYYZrQpsupmaOEG57m+
kVyPqSOjzAqvg1ow2Cf4em9DjHVDkABLMW3ywhaF1i4TD0S1Mez2r+tqt5M5
fhruCGGWO/ySAvgdB+L3tBVHlvqS5Aq7tDEOVL4Bwer4ansQSnWs6Bu0t3ai
PiNElifHa3V4UnqTKvSjimYG3mTfMxsri0bVYMz4Vgdd/agJd8X6zVfjAeOJ
Ig/umpcveNQtyZwrq4W108G3htVMm3zEcri0sp0SwWPBzOqF/SZRNCWpiq15
vxpHIhmtrjaMwfX1AVCIg6tOu0A0UXwhMEnUMJckJFDPtHktMnELkm+W8Kn8
QMP+GJNW7v0ZQI7YpCsb3I9uyx+5qJh8RgtMuSOUEHFm/4PYb9XcmzRqojGr
1TwQuOYzjM2K1dnM4gZVMSktNP93uG6FyB/9Oaf3TyRVY2tEGdopmQFpF6Xs
lYM3yFjlWfBBcvBHdbFkQNcclrSIHmpbNTBmSnlTn4h2i1SDpomIk51GepC/
1kxt8sNSOJUolfCn1KBXuO6c7hvKHWv1eIlJnVt7ra57zIYjQIPET2+1936G
MZAQu24bMTHJHOkVJGyAXyJ7J6OSplH0wJUnYazM9gV3lIJT6e5dotE1lICP
19zvppyO77BESM3x/i64VydX+a1D5LfdGXsLBmZib+MB4V+ANj0lVhhVfGJR
6b/KTfcYKTrBiWr5JFloi+TU/4S3tC3nXgE5SkWCQpXfTGi6qzCV7CO6kI2z
3jRvwl+THXQrTIOuXlfi8y8jEJiL4kxKYVqwOZjZWzkoTwavp3S3dfzPv5/w
VLfE1hVjDCIMv8ePQ/Qc8+etTD9i3E15URFNBYZyT/dE3nHCWm9EmCYxC7Ei
5mOW0liQtKm3/7EWPkHeEwRNWcrYqfhDGjiEGt1qc2mphxRAdIDqjD/v+Hzj
1deDqSMhQnJVqlMQmeEg1ghPYbqCITh2bVb5XocPIxI8CxtabsnBD+AmzsUJ
AOSy8sSkIXbaXuLM2PjXIONsCUBvCOLVm9QQzIzA+WKzgjH43B6DcuL5w3UQ
195STW9ubpxKitBK2VrhBcK8fdT6kal6YVmsWv2DleXgpuLW6d8X26eozIcR
ncytvxapfR+Iqi9olybvel/GS8YzR8zxYL87jDBOhlU8m0HysS0vz1MpADWA
t3QhT3Lpdd0FIXuogWy5Xn5s41MRHumNfVSkPrvkQaab3dTppngs6PpJ6fb1
MDqPK/Y75bidWDII0DIQAyVIAig/h0C56vICOHL0YJcMTThvx8xrjzPfn2G/
dyHCBMY/TYvmVAeSzwGtmMoP/GeXCiLkl3ahUa6pzVulSRtUEcnwYlK4c5ag
ElWCGhIVBe/NOY8kUr9rUm4TdntiZfQRm95T2tJTobLhMVlnI4UP0MXsU7Pf
yZFhrotWSt5MgKrnyDeNSGy9E2eaibjcVp19YAR6mmFP5NDK0gln4DRkL7h4
v4bKqVExwNowuV9/agQz4eqcHLXhKeYPj8zYTOYkoxb9vwJtCovko5eKo9hM
K8MfPX/FmLCuI53shOJx3usc+F8Ub2VkKhfu5nLWu0ret+mlNItOzRb4EONf
QcG6O/IYQESzkJFuy5Hx5FR9rt+mVBL0rOfR9M6tv8pxCajZfTt6nN6jp3Te
IBfwqEyXMDWr6yyW+rH3xjZ7ydK16F5Kte++obJv/5dqbxzB/CuhTSQz4XiH
or9/WSUHPzj5ys7UIOY4q0FcpySIq2YWEShQFMUq+UOh03+2JSkQUb1U5OjB
XjjloGwGtSyga7CABjqtmvfN9HT9Kl63oCEwDKXFAKzKpgZZpwCBijG4jy72
E3Q8T8kO9qqr8Pm5eLmfiQbhZRtnkFb3Kv8fASl6UZbcxGLY+I3L9WWYR56J
5or1oIzDz86pxGJjO+OishuE8n9o5ia5nOYy7ppOa0U75Wzm4tcDZH0WH+Qi
hdrVFooqChY37o0wQwfQb+WkWVqZaIaMh2SOsU1TodaAENUQip8LZrAEgwiO
IcWHYMFDVen4BI78DScIaqbspLZvgHcjvu7BwYj/XMvDmyRrtDNYkWEP0vA5
X5A/McRSTHcMnf9h+Viw8b5AArOHPQBVHGQtuOXu9mhJzw11wU+Sq78swBJ2
lRSI5OaJUWp95PVzMdn4UwH+9AjxdqF7T1N91xRIgLDiq+HFLJUSpArUemQK
pBj+yyHW9tv/ufoXaGkAgLoiLTKJzfIVlW8ytgDvOHfl69aKdw6RLlZcNSoK
aCrzUULC8U1HL4PDfKDQ2pqLPStf5oX4SAZPXRt30crqpFBOwb5hwZZOuS1c
m4kGhVpiFbfXXesTimh1aWGG/zvG378MXCoqk45VKCzEYRn2U/fALTSfpncP
N0hBU25dDOPMCS5+6NaVSjUEFhTPwaMfNS2q/Me+OA1WC5pprgK35tuRjWlA
8/EnxFsZyFUrs3upvknuuodTjXAnJSx1nadzt+nEIY8KFSyCinnYkJY9YJv3
mH95G+y3Ju+LDj6fT9KeYS8Ruz1WLYqKtNRf3AGiBuu/AdNf6o70MdICdixm
OLtaGFcxzFeBBQ7QjWzFP2WfS0EYDMgzJ15EgxpsCa8tZXG+jtEHz3zWSpFj
5qNPkxVO1AAvfP37RPDoEIXToxzadEDJYMtYVhXO+sYxNIMfK+C5I0APPa4G
zvfWJAR3FJZ3qid8ojZ/WJIjFyIND9p9jV2NJlSbwhY/eN4WYTM+rSWQr1Ul
uZdg0ofGtGJxp3SGNt631i6FrcD6oPpc9elFqaCfQ4cuAuDB4lBIgt1ewJAZ
LCx50RJ7g8ZtWY1VByLFWTEADMhxunA681bJ3vdG7RP7huNfatVq1I/baVNH
i/tPyCH8noY0hIFegOLh4icRUE2swJped3m69i1GRj9ao0hibxLHj/qshXJ9
ykEq+9Wg9bBVAl0c7OGEXf4pnBKxMDMNuFI8V0R2ws9UBNwmLXolnF1ZXvEP
Hsx989696YzAn6waZjfNoOBGz7TwZhsRa9bk6SaEMXJhH8HGevI5K+qbCapJ
/AQUAS8TdZCrZ97YsnZuAEVsUibb5mQQZSx1Gboiov163+EW+68ecgdZN97B
TPo5nCYo/qSw3X7EoILja3X3Bnc+wpN9DU/gqBqciiBvxHkAJUw9FZNiItR5
GsvYgVPMhk0jJ8IwwAiT19uG6BKQxgm5RrB4lB/zucuw/iqk5OrPKN7l/FAf
xARuEfcQcfkfQzVH1hHutymX1YjDDj3jnWvo3xSwmM+VBBzt8u2/U3ud53RC
9fcMX2C3TZQEADBC8VnfBt2lkXCe9D1aOlB5DAIMX7LwS8vYsCCghoSZVLIy
T+SQDAygb8L1/pL1k3P5EqmXFr7Kro483AxKp/eLyDWSLzWnLeiXBntqOQNh
N7pxLNydcPO5n05YDOdLTk6eu/+CqTAKqlUwEw4KLqjk8ZG5n4EzxWILgg8m
29RTte7Bi+L68aVuPeAbGIZyEoPjr/ZrUnBmlGyCqTkMMPebnXwUuPmXpSXp
l0jxeVHlO4Pd93whyMxkHeXYbq0Ul68iAVAwgIedcMwS7Rvbl650pbcLuyfl
Vq+ubXwG7GmGI2fQ7vB1OD045StGFoCrOC5mzAzSVKrgTo5ZSWqf47+YOIQL
U1p/gnYqKhwkme9glQ5wU3ODCMi0j4WJkSjtG9ZMgDi4RdQtR9QDhu2zs7wk
i5N9qN3IhHDv2lFigiwm8oY9w6qoN6/vjkDCcy+4K4CiGRidhuj6pcBtFVCB
pav8Oke1XxIep2PbPlKIghf1iyQraLRYpSaNuSics39v7SGbRP9fG3PFBNVY
ip+MiKcCPEG/9zsjxczqdSMozQniyfM8Elklap4+QJaC9o99afaZ2SQr04O2
Uh54aLVelbQIG2KOQGSt7CBTHF9/Ok/Pp6JuxAp2FkRCGkPMDaEbB1M2+LB2
uS3kjNOZJH/DSABixim4TvvZJEUEx7rQaz4HvRQl1CLLCqIwhRn/qSg0SX4r
NZFhk5UUt1pgnMMvTm1uUI3HIcvuPvoJagBecgfng/RjOdXVcqjDfU0swAAW
kSg+ZnQ7hYlcVsAq/EtnrWvkLRo1jxhP7tlzvJiBSLVwBZDfF5bwJT+by6E0
gY+kgDnb21D6zI3GJUH2eGF8YV2FPbj5ZpTY8Lwg7WY/ix5mnLiL2cHjxeBA
VXgXWWrj81MT+sJHhVZlDEt6MK8gSlDGwmcObLozd2C4I3mZopruTTL7NK6b
2erzDpFj95eI+mRdiPdy0Cl5xOAa8HUNPY+R4IDQKU/slIHj5ONazpoIz/zY
Q8Ep0ah59QbG+Q36lpuzyc3Gccx4rRHcXQMVXRszNO2TXEVCgicsa9JKq220
6gLonodAgBX4VfibBJttI8ujwSfh/I53m+feH2lZNyfTEEYQNYnUESATchfs
2N/zeY1OIwhbBorIrQWAqd+fg0J0iGhXcdtQmwfHRCDMAzzaP6p6UfTd0C7M
lRqiPS9daCICtjkiGD+GbghvVSGgbs2HtAKIAxYJ1zBYRNHuNG/rKzrEhHAj
STpQvyWev2VAyG/QJeUtJnCWNVO7gtntCmvO7l2OOFjr6JvVDGkQSUI7AZls
CmFURPBhwjXBRYHeJZBsf5Zo9qaPxuACUFB+hKbs0N2TXI88kjAFrqiig1W5
FlQfNpDs2A74f1Uzfo+sEAnMHVHp9PcMMi1IMCKTzkJ/pszKH78CW+Fbc/n0
/43J6BJRupL4hsIa4nPlzKPPbMLsYI2CMTlF/UAcZ8nfkP8oReYaJfWVEAFJ
fgavSRGzJC0Ve8TqHWofk2zgw+tbunrPXOhmh7Zt61sUh/3vaUjr4qXwtOLC
fUpNYWRh3PtxBXrgWjFzq1nYE6zDLRr70kP/2JoLZpCu/dOZK9Jktg+fLDXL
tX2jzIjLzFguWz4Ijpsop8UwelU/2rE+ji/sZ8l2YIaJzYjjRFMGfKESPIsd
hYKAsPUn9d6xQNwkhavLFr03qFkkIahJFmscdS5Vj7aNKCASxDTsIgzFVUnG
7jFdgjCYOaWae5VWMlS81SbEUl7z10Xqm77jNs+okkbDtvVtNzbyJvgFA+3n
8jo3yNxur8xuPtJuEe4FnMhv6iTfCoGzbXL39IF5UaDGTR4gVR4gG2UszUO6
mfTmHrARye1dY0jYTOHe44X73qo5cGZWzr2CgUni6c2seGksi84SiU70Xyym
jFwP+WqvVqMfKGJZ6spuxqYHMBPR7dd8oHVo7fne0bAKNjgQbsMroElnN+z2
quDdPyg/1vMXL8ITGrnywUD/KmA7UnEQXlZ+wi79mqo6mXCngFfipwjTdUkl
DB+3cLYhsjTtCSR7BYjNmPmcE26SZqoE0AKrkKd7UDEJnqNcHk2DBLMOS7b6
FYgejG+a0Yg7szClwmMohHf/Xi3H3wEVS9SD9przMo1mjSXAEjcg1ycTRkve
ZTfHbrSkanpcKWrbHoFabD1HFrYQmCgx2A+jPvTK+pIhnV1WPY2l+GiUnbEv
vJvjRHdhwg19VBT9MR5gjVrM5E2meBhZSDPWhY2D+6+iSdxgu+vK4ErEntwD
tpGtBlrQxoqRwcmsspnU3SKXU/omTKZ/S6YuzIdx1ikPMNmbMXzQOFZuDCLw
fvM7iahdQyrSIShHMDGEBQnsLjMgEHv99Xag89hBnwfIe+li9dYL+vB+M5u+
UdNcHgXtT2l+Wugjd/Lp/E6hb6ywSv+ilrXIFU99SFsmajL7wo8ZEyYRKJ3y
t6cihsXZlZ4zNUXWiY2EhOQfqAyQvYCPAQl1rgOtpxnnzttcbzA10mWNyrXV
LJbUlFU50vLR7boVPVjhJHYO5hMCwHQrR8Ab6iLfsd0h/Fyu6Q8iYVXccMMj
QqJEJUvDTY2Ijy068nL8RTIq7F/YjV1jbJ3tf7ClVS0WeHdtsBcXXbHfb259
XbmrYRRs0r6dT648IFYitL5zAj4e9r/ywWZNp4nz5Q7r1/pWw6axfstMcpMZ
y4VL+H6HtFRmOm/3iDABz7OVaJn/hhPMIKJSJF/hojhOESC5BLf1b/8g5GH6
cdSaMi4W+2h3wpuoqJ7bpuYn7xpoFtS5TXibPVBiMO4qy5w+7ZkLZC7WP6qc
IJzKz3KlTPq6IIYaIULUfrqprKZy4clQIhpnbaxqnrXo

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzddL2f5TAmViaUvDO9n1+0wajCeA52FLfLxYKF0oe4GLUUGctq2o1HdkzdcYTyg6ClOOwZ8lUifbwiPkwxFh0KQB/0hQeQkaP/IaZJ4QL/aS9SQfte/K41W/grWAgxzI0PKLk7/AyWIW/fyyqMmcmmgPHWfzi38KWdaJ+x/XlMaei9ITWe4+L+aYP/3rmRDekN6pO1jB/8dbap1wklb9DaJfOHVaQ9psIT61I577JaNJc5/yWWYQAT8foU40/QV7QG68OA2U3zNVuhFRUlnO5CvkVAP/lrp0MINn/XKv4ZUD2CZFvwCMxtXNTnSZr1FQVlIrEfTyTHJkI2GsEu6IjkwHnxGaVr5XZhY5ex5QwIFdYpjIywvcWrRvV10/7UhQ8HZkd8R4c16/7h/b7422RfCBMh+y/6kHeex74xty2VJ8D/lmUAYRHVwyNykpzSHPR/xaHy0+E7dd+KD8LZxPZu2EdkFVMkj3q7SNi5775jJkjXFlFYkiUyZcqds72UZBkk524Pwt+lF8fL07V+fvIf2ULkPGXlIf+2PUkKSRSbjloh/sq8rNrKX+vEbYSg4nH9Q03dtC5eqLTXjSkg/ZU8vfT2gkXBQ+9suJY93BdJO/THcSRhdahLYwz9A9XtAvVJTJNK1vyUHhxymdcOSrh2/vq5kPnQoXIR+bNPOYS0M1yQTkq4+FvcKgHCxJYrnbANmr2TZyRn3b+1FzwNwremllO+NIDJaas4w+WI5K144jg3Ckfs7wk9DcK89G3llQmF+oZhJW4x67EKNO2ccyBgR"
`endif