// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l+fkWvLklnqC2a09kn1gdgsgiB+3kD8RMu5CiLbSyCBglZqB7VEd67bL5S09
K+GhB2SA89kFx+M5vKT1ktW86k4rckKN3jdvtiWCTv+co2KPgdh9eFCtQ4y8
K4MhXFz08VJk/BBD8FkDMycVYn2Wv2pDybIw0q7hv8rW1apiaX6288h04KIN
X9NW45wL2MzlMTmXJcLAnokyKijKGw/8DD0oyyONdMvmxKV3KpXb9whjiH/m
Lq2YdAY1kjB4O6fQFCeV3D/5e9llAJVf4puMdqNxvZvaVegujZJGWVSkKYuc
i05j95ZI3vo9Tj5hDHP02hSESoSwNN49G9L4ENZN5w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gp8PI8qH41QCcxC83Hd7nLxLFWqcb1rV05wYAIqvR1d0KsoSW+gtEopTnR7P
9tB7CEEf3O3JLWO44BEwyCBrqZgcZxXRPWQdmGbZ7+dPQa+emUi4U2WCO8SO
Hhi1iTGFe7MysyKLPsIXnf2cL5eVkTM02us6BRTFjy1snI6uuIek1Y4fqB7O
yVSvrCKun9sT1UBDenFT3+2/5Ram4HUHk9ZIFnrx5+bGQdCgdaAyDBtEvobH
VqIQbOy2GlHAVcyaTfcDxEJKWyVUD6yG5fSSEXll6uej/Xt91UKeO7B++0TQ
UJGuvu5IRNnimQBqwCnvu4Jz9lMB8BmLek+s9hpD3A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cz6nHXACIplv2TWfr964lwb8ft96k0OA9nSSgdHY2awn3W9JtMa8MkbTlCjA
jUnzcKOjEM6zKWGt0lOKtWdy/Ocyyh83zIHb6uraXMAKcADAkfT7Y/rKB2gI
H/Fi9nX0qvqtZhI+zAff6k3ITy9jNEKLrDyojOjkPdTRvoAfKyxkas6bPWZ2
NfwV6YEA1Of3FC/JSqiBCGmTuiOpdMGjqCM7qiKFVam3WFHxufcYWbgttAWW
m2oInBkVfm/wxz5VAdoydU61UiZLCj0vBtPlyOuP4W3ryxCcWiJvhnZL2Wuu
gWDG42JVGEcFbxDqCru44/WFURM0qtNpVGMf4/7qPA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DtI+HmlGK7IIOchETc+y2XrIo+fHX6vsBU7dmHqnJs5Lws95P0m8mKMJbtt6
oMVN5clXWv9/o8vVRq1IZVfqBnKNxl8LgrDoU5ntVrmwO3EDGPtCFmi6SlLU
GHUHm4RbcBjXc3hryGQ5Oo1USunsD4TWqX8Ch0nlVPaJSZ899br+sLaYYraq
LT8Jc8K94SSA1TLCftbHf2JDfEL1A9Ni9Ioap6UBTb65R2PFmLLBsLnDZ/Ne
eFNZJitagGdq4KrNq7xfgoY/Xr4+kllP4bf7oSVs5axM/919sbnyNxk6htAy
y8w2I3AYBfKOF1GnsIM6TgYYsbrdS3UIoKeWydl08A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LhaCD8dyd9AacyjHQIOVZnTFgQI/T257zpSIOvBsxsgh5dchVUwvpe8cYn16
TWEio/e1cpNsLkuxJoGaCylYl+LeCu7tr3RvhUwfexwwIiLGnW54fZ7qNj/y
RnyfMoW1dW7viT8demuzhRTegBdeLjiSmGmDcUhZuwyv1kqYFto=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rerY77IclYxuiRfQasVy5cWz7njjPPaWcuMcLy3eC6FTmWfvxFeXrqCmiWbA
I8Yf2cn1RKig11tcPvRteOVyrOPDZUlG3Hr4sNVWt4Q4yNx36vEcGMYBAN1S
FCngH2xQEgErRjWDiDje+U4l3sLC8NtRW94Jmsk8VfjdCoY69LezzXjqHlAa
dyIgKKXwqDaAuDMktWfKE2escCDMmHxot95oFBteTufdqiCjAP1Yxk+LixZB
HReacb3Ohaw8Jywb6PmT4lnNqpNwfy97HQby3bopW+406OaVQYd2eKowD1Su
0cp2Z+GijKTMtZs4nXVIAZQmN8/0gQdXXCi+MdsPNzQJg4KPJTv1nRwJNa2y
/k2wmJjf4hE4qUJmkPDF3T54cVp4BE9JVFVsa9HVYVjvJOeE48/uVIVYthiO
KO0f8HqK/T3gP9TEYfxsoj3mf8OmiXJh3yvToHyJYa5NIRcwS4jlbAD1NCWA
KHl314fnc/9RTU8BQT31TQ6cwuvrMURh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gM0rMmszcONetrqnmWdbioQEOwci91BWLrwVEQ0bG/BC6wWfeOCtvpfcJC7z
KjvRrfEqI9YM2OtNbawS0hCHy2L8Z1BYFnsf2zKhDQnqgs/+QWsYTGZGiqLw
H53dikml44XxfYyKwZIxL3hbIjWWdvVMUkhOLaF//spJS/PF4RU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Lpj9VmdYl1vOpwvfnCcaaBUDjMjDph0T/RX+80g8OWGih3gqxNi4Bdw1oVL+
DixplHrH9Zb6BSedpYW9WTPZ/uUw955wlMP/udOTiAFRme2Ip4JTSzbjKifl
YCp9xq8wtrKE8SNjFnQH3oTUa65cVz981sBW4LJ9aCOZ+kfHTCQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23552)
`pragma protect data_block
Wgsi3ZuM2S0tXZaJGBCiNCaoSc3sCjZOA2tKut0o7YiU5DrxoBBm3SDEeJL2
hYkQqQr/S9p7XULrbnY/D7STB35CDiD8YvdXgtZMYsijz4sge8cuh1AUOwWY
0D5h5iMFACfdoedEXqnNyBG/FYWJsfdcHuzyRrMP5wA+9VMbOCF2SBx/Z/ul
NICEiGE3EAN51XDY3t+v1+wuY75n0iss+QgV+/VMESOEG6jjCNwUdrD8ZvCB
XIGu9jEj6kBekHZ50uVOGbt3EVY/vXy86y7LmTRgm02ho04axB7iDMjhF2wr
mbtGbqF5eTIwnIoiQOw1/UGYdEOIQ7B1b4+GStzvMIpUV49Ol5635MhV1Dk/
sk5/pGNOsIj2ZfPiQPycGN9xeKPz58fKihRBiN8Mkxg6f7OI40u2zJxPP3Cs
y92+BzJ3PodvfDoJNbDgvZ6xDgd79TLs9CjrWGe9kMTMY2GphBZpkSjzcEQb
n7AeEnNXQPlofnrQxTsMg4dgyx+Iob+tzFQGxqaGt2JLD3Ql8RM48dzkON/c
+kPk6T6ix1UsAirk8O9ORkOdYUDY/fUWI8TIz/FaPpjMHvshg0xvSrv99dJw
C8TGsoOYhRTgQfyhUFdLBtdq8iK4KGO4QxcG9cN7GWBM1wJlaORlIlvKKHqj
1C4ZBz8lEU19pJVcQ41Gn+rVcnUOEWZyjEse9xL0ZfwFr0UeX+V3tQnw1aiT
7EFg5RJXlJoUHua6cPnnmArdo5P4uoFVnWHC3mKXwDFAc7nc3rtYFgZzyRFd
lfqDTB0fT29V1bx37ytYo7Lch+F7VNDzfKXlmsiCon9CUMkODgqmC3fLG+GC
dBoAuKbjzX6XpyjLEJfUvQBbWdjjkf//HW740kea54ryW6xlAvCd15FAZ2fr
qt9iyZee16epW+4TrsA//m5vc3YjECbskceA0ammMEpfcim2HB2DHFlraIha
0acdPiwlxrLSAXpdZ9CqQk1vHZk6kQ+FXmjWynHH+1L0v9FYT14ryzv6F1wL
fnEm5eBVzO8om0i1ZTT4BanFirJeb6efpK1MSlje5aGtL/HwmFnlAG4F/xuM
ea+F/Yhk6Wa7y5S8AKIY+Iy8INsaq0wEZMXc5ZCvOWnU2o9tFAdAWx0AOU3D
//NRTXC96zFnmiqEpQTQYEZe/CrUxBd3oYx/Rf+1699V0cDhimZMYeem7k5z
R/dT1JTq60I+c/i5BsJdT2sTVSH/zzB0VbudeqbTg6aRHFpIJsYVO2P4DkKh
TJ8mn1VJ1Pm4hIuRDOIjh0iaB5lKMAxw6FDFgYBHZxGHgg20X+E298S6daDD
Z/CHTWAXYroTRPeSZgw7FQwo+w5QiQb3NL1GAQ8QZpEp39eOXtdrvJ5a0cqU
HP0CxfiZeM4IaRBWh/khaBvVR584Q7kL6dwKUem9jOUeaQWcRWEOs2SrnyQt
jJl8Rms2uRblBo1eQ5JjWpd+U5lwsWqBQu6ZkWgxyTgj9vEtYST8HGfRpHDV
j8098QXltypK18fAyOsxvCer9Tj1Wi6cEzMKykpFPQAbe4fX/GA3QmCplXwf
Fk0oLBUTmZ/Ci97qIT1dVEsqdCh2IpoC/BTfN+MEqcgddb/fD7Bhkhux/KTN
SVMxd+bCAI+1TisQqaZKOM6YpTekqrvVSHyD0+0vJdR/OS1qfKcg1vFjn+wZ
3FjVvVA7H9axwQt1IBVsY6j1Nr9I9daMfZqwTd950s9ybLnJqzrHYeUfrJwt
EtKHCQ0e/oNVStKQhBVzoHh2KTzihY9Xj+M8amtOHrka2xLwKO47dIqEDH5X
QjGwsS8SY+eK9LBMS7HPB0l0mDpLhDP490kBfdhLQJKO7rKgGrw5D2DmGzlw
dRC8LQp71G3w9mDSsTShcCEgAmhVSQsGduNh2oEadYNx+no9QygqnLkyoSEl
uSO75SNIpTsP1978heXGJWAo3mlESV+S3tClaBdqPMG0/luff+txgBPu3iXK
ApCvD/ymAKj0XprngP8BrsXW+1jjxtwGgxFn8IzAQlQL/DfTnDkOcNjXaKa5
WICgoMvIg3cZxXudxMSDeMxmcbTlUHVPxGp8g+lGbbriwTl2o/YsaQTPfXrW
dFNPkjLUvYkG+SUb4BdpV4PlBxHxpx0oiw/W0grfdwAd2Jegj36LrVQ9X+4T
XPX/YECd4NcdGP0nucx7OxKEo9y0D3lqSaJeJeGi/K1d2dnvA2x/Fozr5WE/
su98e8WpcGbLxF9YE1XVStg4s2Nc1tIOxCJjTyfIN07ApyOcWjD5hyO0oybJ
vDPiq+ZSBhOGsbZiY0PbZMxIhbH5GWiZOIWSOFK4Iy8iZUSQEwFq6PCGA0gX
RzrKKtboRoqiqn7x0K22d1uWy+MFxphUac212uJh5sVEOlT+IrGvCy/lRHOR
O1ZJST0U4+e/8l4VTw1AjKa6YQnzJHqZVYyVOJf0TSqZ9GmKZ+OVbZ0snWvA
Ok4b2smfKxW/2z1mC8lYgN29yhjdpEOfuRjPZB0ScpBrPo5hbLMQdrH8R1YS
0tXaA0dzetUeKHednNAwhzp++SVSFJqwdicNYT8g+UVfEUJQnyWuX1PWHKtY
jQUG2BlgJHCfDPdJaaKHMN3GYM/YXw1Y61+/RwifuEVqJ5XcOZLY6bb0eyO4
efwlvTlhkS7o2E3Brc4+jxZHz678R/VlqEr0ZqMpcKwWDH/WG1wP4rXzNIG2
3nPmxqOZ5QKxV9k1wYqdTJUIZITG6D1fpxXkuS5JqM8v+gQw8lNLSDsYJiyN
HDQfY0VoP5akt9tJ7Z1lI2KLGAL2g4LXTcqTkFyX4cB3mdsF+pwBxT5fEiSv
L58JLXI9saxVBjSZyLFrhZ731wMr0NU5/e07gv7sp12ognRc4EEbQq7zMbZn
HzBamFKAPkxJXy6hVsbIUJbDMeoB946vMGUx/6H903p0ZfOea3doZBVc27Of
4hkAV9BT3QnZwVrnxeHAefdw6mQQ2lMluXOnduMrJYQ785rW4M+OhBhLgfX7
cTyye2WJ21GY/lpXtGkBpmW1cTy+VVv6nl1+mfx/5Au54F0rOkmtjEBezymz
Jy7b03JB3Te4PnxVLV2MKoC5A7MruEoUnw0/iu0emro8r8+GMsXuHiK5/CQy
Ajof7IPOr0lRj3dk9+/a0rNFl9JZEAIsUFcaU8wyZmD9/L8GdgIhcjgUwpGR
02Eoh1plXUoDxQNCVNJxsXoXslxOB1fNq9Q1/Q3y8HQ1ASDBDqcaUFXxK9Ui
Wa7Pk6k9kJv3QoOlXoTrPTb1EXp/8gRfIlZkpawxNmuffsRH2DPT63B0GtIr
atHoLHt7TE5lnM9LvwCZ1rRO+ENhkQl373IZYc62xoSKyltGOMRMW+ungux5
Dn9/LB+N9nwtsy+zckVyA8c2U7iYtWV6L6esmsH8nEnwMYoy4DBCuybwF47A
2LHqVTe2+RLfqnJsw652BcMurvEUqp3dOJKUbBrWKvuYyuX+y/RlYHMeO2Zk
gx1TKMD2D3fIAJL13ylzwr5mBnJSSOPjY8gFYGePgtXpjJ/NsLbpwMA1fqgR
TZ62hO9TmuMJBK4Ek8V8WIUZPQ/DTBxqt/8gswWQIyJvdPw1aTmwPgNQwRBD
PChSxQMh4ejpBiVfKS/SQupUtbIVP9UVEsGp1EgHAY7+6F2GAzSG2s9+37ud
tmU2AnJHj2CVd6AxUmhnj/LL6SGf1ApysrrqhagBcjMHbImys1pawCCHTkjW
w69uvktoW1rtI1duso/5gjaf0r1CUC3HSyTp5xV3fRR0DVZDneQmSUFvzOxT
1iXYyqtMib1inPP307x0xg530xy6L8eSjCn/uDGmcapzBwzaFlhoYDKcqecU
ZVAlqoa+aX5d+9y07W0/gB/BhaO93KOdIGbZ/bWuIye9y23VJdnx/YI+fpko
/qUzCtA/slJxVj096//gCDxRX5LsKwtZO0smfyM0+/jbbl3/sCtgmC3mE88V
2yX4E1eQQaRXP2zsmWDOP1UYcuj5/W+HNqKhT++6AZCIYz80mRngoicXdmsT
WHymHAGV7kaaxDNE3v1uyMiDW4t3VIxf+t4BQNasG1GkYQrjR8H0dXhZGeiy
NoCSvpwkLMycsWDJbO0NLWbP/zzoQOeFsouOxM+ipPBA5CawKgbbKTidmDJV
kc+MHjio9foIHuz3vYlx7JndP/J1BHaIPNhI3bBszGnaPdpKWRZDjDmRO9z8
sWMrwka245wFdjsxq1NOkdaAlEbiom/byH6fUBfzs+9EbgsoGRGThBN4l0KU
yMfzAz9Annr+/p5EBGOOGdZSWBHkP8zajqblo7FEuguJXubaEfIlTSWJN7Pa
zVit4K8h52CVPL+zD9VltfZLC0JPj+q5s2w57rDA72G7YwqWhqEAK/Bw+Taj
HLJRJ5c8zp4rLxkVYA8K8BVM7xQip9hhywpPFPXE3jLdohGzTNzf5gfEfAhv
9rmCHL4VpOvwJTpoHPS8tS2J8Aiy4tB7RuJk6a/wR1oPNfMZU+TdvA+7c7S5
sNnC+uBE+4SCaqcaNlRIJhjYi7EWUeeerDtTUu9+KCEKgkeZA0CZNb00ioXI
CJeGxiFCoXkmUgH8Ko2xBQYKkki5SrGTDwEZZJkho+NzdeNkp41tghPacW4n
RUbeBv+JANSvxupYkvz4jq9GwcXveaZyb6AgW+0mPlkbPLkCYERhUx0JhJVt
GTe0ZMY/VopSJnh11r0pnu5oXFMskl8U0geUMbtmNJyWvkQKb7icuLpYHc4Z
2bA5Q+YqWJeHxFUuVXvXcTpdNcQPIwIAkezJwR8AVOp0mccd7gGrMSpiHZjZ
VBiHNCcRVJRJQZ0/ac36fw0tF/BiOg1WLVphBE9eB6UTpjuIlRdNiGZDVBi1
H+6R7qCMwIHP90d0o33UOZyyH8dYP9mbaiLgx8dvJXpj+D6CzRStniPDnhDT
7wmSDPDNN85sVuiNDlOSVlPUSRJLux/NL41ZrwDnivixemBmRXGdRhkUAr1S
MeYM44HMucbXYdKg7akYgIuT77R7/WKwSUlSEzpkPixPIIueFKVMYUGixRd/
sm3WZsjyy2HDae9gpaptNL58LsBNJT0liDnoBypvQ5SpPfnXyiIGSNAfKlIC
R+N4MIw8XN66mMEBAnxnrYHCB/gTMw4eH2HpVEdjT1Saklm/YjVOmdpv1OlV
UkDWlfRIE3V2CVCl24HChsw+pJyzw2gpGUbkB9YvOWZ4NStO1LxhYPacx0z3
u9aDYYvPiMZ0N26ft5xEiliUpzeSANYoZ0WegJbhoHkDUd4LSZQPvsZwVooy
vdEMrvanXKt84IJJJWwRi0SIkCtLV0CY61ceZmrF0Tug9vIyvFDIMnMjS8b3
qCb2W/ZLDKrBC7e9n/MywjvylYA+F5LOkYM+ADz0pRG1/J/4ujehiHVuUXP5
c3k2No0tsykgkCvSztdJ8ddctD8gyK6BQr+y2tTCgZpf14xwRqdZm+jkCdtJ
/f9Q1bit6d7537eadlRFdGKNNcGtv9Oqt45Pb5FKay9H+AsaU2NXt8JoQDV7
kk0cuYRAM+t5tpJwCGPBsKXk0yHFIIdrv+o4et6ObEqZ3ykVwGhQo5IndMQh
oZotw7iwIp/ZQm3WBcjZVGCso8kMyKWTpXOctxPkSxCnDt9v6p63OONshIOy
XO5VsVo8LNDcdn7UZ+o01uNjUuISDz5b59dI+lXV7UAQ2t0F0nFQVZz6EZ+t
EqKQEaxublrPDLjweToS0IPTTGnL+bItdBG7MYve2r+rveJXSCigldcFHp8M
r6HikH78Cy3AwaqAtdmKm9NKRrFwE37ItJmRn9avcAQ4Zq2Ci99xNU6uDM5X
lq/FE1tbebfhbNrZYeaDT2vHJbS+e+pMztol+Ifv8Z/EhnsGtdvddNtovEHt
yDRDvIpFRSqNs/PoEmy8UPzewc+taJG5EGOXtoYvtl4eGl1qRUNTSBRu8U17
DvQMk84SqGd4Q7jVw8EE+jcnfIAXsMjdRZHSrHi0J0MSpOKAcSDOpyMRNJAE
/Bi9W+DVmvq7uZBpB+ez3S9ZEBPeamz8MgFoDoLRpxVNQyZ1/Ts9d8VWPrF6
ZEIImQ605ANa6M1RPZsk/ZwDi6UVWwwbhOOKYaM9jOd0JEByaMTSrBvyARek
EijdPMEjYqFback/ESZIzvMrOBIWnVzTxCINpwPfnolIsQWafhKf5D99mZoR
T1NMN3zbSx/Tya7Y8wUV13mc5H6xXNli3sIq7L1zsJMdH5SwyjeKRRxy3vq9
jok9+3BD5vyNE4tRxmBjEeqrip76L4VPsHDTWfjPTf9xxfmLVI+n7Lo7a6Dp
Ptq2QxyxQ68KPdxJVrlBPhH+7E/+6lqQ0IgBoxPO3nB7/OXwMNgaSAMCQtNp
cQZYNUsLTy167gCsB/TWtfvZRX1M3NiKa+fgwTNYMt3Yn9ZVFh753teG/Ez3
GOvOuqIGFlPNC2x0DlOZxTsEYpa7rA2TnkBuT2rLqJwy9FuBZ0FGXK9ycEV3
R/5R89FkC6mf4jBLqwoC+F3BwuAbuvW+bCWRZ1dMvR+I94THycvLQ8RQWbXZ
xX+Cqfyf3JJ6lBCwsZCzmHLHybwdAZp+BjlwV5G43aUgErbW8g5JuSOE9vVj
K6yCtPEOdlN6y1gmVTkdGFaDLrV4D3Xg0O148vLfWY/wIb4f1lePeAtWNEdG
fcWXbo5Ml8u6xCAZXiUX+uSclh14Ven/DbfxL7tb3TyLt1bOgyTc9ncMhCLj
iMR40AOAaO+ICAX4g3TntRjl2kFRuAH4P3h5viaiP8P/PBKPkguCmt30QKzB
egYHWpVxPkbKOUs0++aFFujmcVnDoDhyXlVUGFzctVaKVUtb3ZZaltlrZ/FO
EgRH/vSaEIR61PT8DJm5lbBV3iQzac3up/DcafyjyAJ/n1E8DI8b+DOHXnLK
UT3xGvx4QpWTug9SOtVL8mRfl6+eYacp6hSQxli2o7Uk/ctApuxb9bmjXguA
zOwsiQDwRf1/d4NcKrL7EP3h5OWMKlKRSsEprHRvmzucEUTX6pFpLVLcfavm
fR2FT5Fw3YAbGabs4tIHPd4k4zY8beUxbceJOOTWGI1JD+MQ22E9UFnBSSbr
Wp+DUBCZzwpW7RN5PvkVZzaeUljzHD5buujcyfwJFGssLgXjW4N4Oalka32r
wy5t5v56hgIpKd/iaPXbWvlMwXtSp+YUdFOHMFlTwdEiFPGMj/WrZcEDx+Oo
oqaePK/1CIS6nCNG8IuoqkpgCj6sAzWTNmvvGC6FMS3gFnwjg7VWpEUp40KW
wPh5VK9J8CmxgDwNp9KS7W8dhAMf3XF472lrtTRSWz1WIRJvgyKKVxLCEZKe
7slxtQTvp+OQ49VnEbBe1MlujhsjOCG9mZs3SquPGyeIpDC49wrrguOd4eQ4
/TOXV0x8MFtXGHbdpAiyiGiqp56DFdQfCPDjUmGoCaPZs9qDpt3+KUWB9u+T
Kr/ItTtCyZ3bJfD1lqamTEMn5Cs1tnK1k6f55C0chdQOuerCzU90qv1954sv
PbLHMgEZcPFrcQFtCey64jjjWbfonrlGsj1p9DFscE43INo+wDBqrU1FOETy
dAp6gHoSZisZlRdE/JRKcWmEXgbojr9zVJwo04Q3HxFoVDHmJrZA+l4n5NrC
sp9g65PumGkDikUIV+oYdTp7f3NCSaupGL+0co14r6ns+G75hplc4gSofcNy
Me4g3ZFPOaaHP7IliBcxm9Ms1Dcrbv0Wjb3GYEzDQUY9DpA8EWNNi6A3gmD8
DgzDXtQp0FLjjCIwMmKOX8C1ApyWD7QU67sNI68+TX1fj7mKjSQRQl1Q2Qu5
zgXNakVIbLmJqf9T8Df5xmc2t+f4Hw57JafHK+AxH3qaC0oae2hsHy8Ikf7h
rJXhpj+TpzU0vBnjKwjY90f/iHOnBVO4hLM7W8dguPZUvQh/75Sdau9xLhdj
fNXNE1j4vtOaIWr/yOQTUDqAYDNPQWQcjGuhiipDJilWxQbq1BmdXeTik7Zh
7ivRvmDLcfzz0MF11oMY2g8FhD/TMwPBFkxxHzlvVd6tSlIUOSCHjX0aCxxE
sHqDldmu4CanMTc2SChFtnBjc5AWl7LY54ihTY25gLTvUXncXkM8Bqv6de0l
d6QrZYCwUR9QTkdQcZfcBaTy0hN5MKYKsLsnU5WcLW4ObEJSDhToIiAq44TA
2pzrpRVQS2e2XHBttWDx8xGwzcDQagmhDJjO2WPoDlxWkidUr/pjTLsrduLN
ye7+4AmRpEFZExR11sAmt4LcDVYP4IJKyDYvGC2IA1Ve1pb+5rj6M+D9Xk6L
F+xXpxIu6pphYQqlX5bgA9aTzmhjvMqKnIc9tBavAxsbLjRkq5Y+fWaAhea9
uQApOrVofascXdUrYMYYeyqywHgfgOWuH/bakDMyqGCjTWiY3tKISaWHj/yS
xRBCGut53XfdHhBBYWQVoPPm5n/8kp0IO7d5nEddgNiQC85Vsom+CCbygNmp
gGVCWnWEUPhlv4DZICmaSPYDTWItZESTMtlGS68v8Fbr2bercBR4mXeOldAJ
HwhgFBHQ2Ior4REm4xc9hKmv7cooQNWcD2I5kiyIylQfrm2xh2BqfaM1X2dG
El/mbpWf/wFX0OMG55SiRzLrQcSFHfPiTY4Va1Dyy5ilXR+n6HhIO6S7HRpR
9ZRHKyHaZzPvFOMFTgRlJjb7qzjYCRvGUx3/MNwKF6tvT/WGveXp8H9Rb1ox
z3nfUIM0VpBY2hODDcAJG4yVXgJsY3H5Oe+BA3URRapTa8P0qm4AmROUYA1H
BALtwAo4hofCGqgrji+P0CQ24c2SaqeN666/J2/ERAebXmCcHcPsNMHkzG+8
oiJdnmhxkhAV7nTBo/sDUGMGZK5qkGey/0R7p9HAuyj5eJ6JzcII3ezD+cCW
nVmeN4HtVAWzV0beoQ2kNBQE8JrOXYUZG2GSVlO8DwMKWdOF5Yk+Ppb5YjoG
Q2BivT3odaEV275spF4pPsD3WRkMhOXz/EHNv7P8pmCuO9HbiOSF3wLSdoNI
hik97m/QFfgSXSiDGOyF5uOp2MBtZE22W0vJ0WCP4TbAPAhHsWIGqkcdzxev
TA6/N1z2BlI4MnRpHp44jQ5uw3BNU3DJAdlu9m56MANiCRkewYsctBN7XHjy
4OH7xAICM/9rqPD5+VbiXoGH21/JlpVocDEnPnOpsdnY/MjL+XPxy42Yn2Yb
G+82yEGTlpJYIh77cBo3BBnKvWXxWanP/E4VaP4FNzNNFnWSqepD3cxAPiuP
oODK7UWD12f9tNE9ymwuw8bGWtS907Imd2ubkH1pB01QOVeonaHL9FA8aF45
fB22uhzKPhEsR//xMVi9evLVWzWv31D3r53CaMriBFMlGhIeXwVPec0qDK/M
21waMplappnumvw6Nq5njCN4unahHbIiACah+rnE0FsiYREtpCwMa/9KRRTH
vH+1BgEJ7mgtzzDGCw8daC3W+WHBJarRbKR7sBIkIggpWlfJbAFNnQ+dTXQ6
fZSU9VsEllY+ygT6spEvRPukfjtdijfA3uH73gcLN4qXbpB3iENcMOaFJEYw
HrelV18twhouBrz9AkmSmQ/6CwaPYP7Bbj2q2d93xz4l6RrKNboFkE4QNhLh
FasdruQK9Z73Hz3pircDOvwp6UotW8XA6DVIHV5CzUJCukEd9K2wamrjmK/v
M7lmqRKcLEc1rb8vXA/Li5Ayq7dGPou6nfHnmwDjGiw6wsZGgLpiDtMN6w/P
oKbR4ITbi/0rOwNooeYRAbUK/Pok8FdyM2HvGdOs+zimJtn6j1JMkpQXs+yF
5L1rSTNoAs5hFBMZtMSwAQy/3cx/fIor/jQ7wQD4LXPFXcCmAr8WhqPbs03k
npUm6u3uCPjdwNU0z58fqWTn/Qb5Nzgce1DoekiHSnunhjEampqgAX+Jh3gG
UA6pk4vC0sZIpZovZO7Yvqjfz9DhHbUsMD8IXrQUrDxzQDn5tiw4LEFVgqUh
ZLsLnJA32HCZvssvsOKbEX95q6RNIRnrS5dfTEikZ58O5GBhgehS2wXh0bvR
BxPX5kaHCUnBITSfpQx6iyPI79Rzxi2IUj1BysYK5SceyggSQBzgW+5P1ReH
6aPXJcuylifgoUUrgKPoIiyEWJxHK6xvGrxUXaHxywIbFLF0b8n+GVsOcwo6
pfnfmsLrWjY7HQN2M0TGADqUXBIBUf9FxeHhRYlrKmEav1vODEMGU1z/R0BV
om0ZIBtUKlwx3YnezRxOaYyw1FvDrvN+8p3cCQo2pDey8YiQYr/i4j+OqcGI
jZqMvHLzu85Pk9vP6lI81CSJtZPXXjirGURRdqxgybZgllQYVo+DgOIjmg83
KDxuEXJY/sc65TXb97Npp3rBnQjFafm7bTBNL0rPm/PANywtCWSlq4n/VEBh
8s1MyEyIV005FexnYhSK20BDQ38/pfl/16aWpq+2mBAWPxn6tFV2/mvSm5NU
//TjgWF4PVDPpM4hD1CmnGeJwUtS9xOcJB4rzvvt3jk53Cd9XaEd4LuUiimU
++uVeLxXJiXVGIsvT/eUK1O/rQhl6FxtAi/Ltx/WO9mYcis3ZFipihdQn275
hTCPv/7JctbLag3U2ieOE0G3GC51GpAcBFcuMwcsTP7fOnmdcPfYYyD16mtH
iHZ2sfTvmE1JNZCyLq10cqsgWKAsZnG/Kd6VvxEX5qSXWfCc5FMfb9W1jSzv
YsgEDNHlQgub5ZxNuHoLOmQL+zc0um4wNOJSJhKToO7XgvRchWVUAXmubhZX
ODwOQcWgEwRvMJ6EIgSPbBFHIkDIDjRjSzSiyjx06LqTVHAt3FPnlolm1pLN
Zn8PsREl24ynZCUavVmQVWpUpKFcFRW5/XExXjrs3Uu0JLJymFuxGMPCM1QP
dqylvwa2HkdTqFZq4d81Zr8GGfAMY4zynjczLLttdp3z2EyZzqSwJVMHYT2o
lMvo8m6DHSLHyr4qIbW75MwT86e8SxOm/JW+HRckP5UZwOTVxOPfvFtY1H5m
dAdZ9xlp4r3PnDNqLhW4a6tlqobsYwmdUrMBNasRdhvfnj2Qg0Es0q7UBXOk
FKIrNnEhocrfPGYd88tzaJnSk4sQi3J0v5fAFgE1H/mv6aWlmpZSF5XoOKLw
Lq2JuNgl6+txQwqi/BsdgNAnS2vQODUkbXQS7lfDKujZRuFbDVCmFg8ojhEw
hYmkB4L1auQFT6UtYaRlVg7wQ8reEfmbUdus94ePV0TXp9SxYBlLAtr+808R
PG2zzDh4F5ySHnELPJvrrhtyAz65qhR8GAJcAeztCJO5Xo5xxB6yJG1758CJ
ZjmbRRF21SvO3rViXcgxsQL/g3Hc5fYHGQw/li4A42W7cNYFyCGuk8GNMGrf
AXBBEQEE9yGHFSyMZhCpK6Y02encT0JOkT0hx8StLudRTd7H7zw/aqz/wcMe
pZyzupDkYK2qhy/sOD6F6t6g2WZJbZcKot5yB4KeMUkcRnLeSyLcyRpWhRaH
M24NzErbQXkGKigiOfJQ80FDstCFGyWS5V2vGnU5Dq7dgDBuJI4+gsJBmCyC
ti3Jk943qj0oBscCAW8rMxXsWFc71i9cdsiwYFd4bFQMHm/pGWaNCIO8He4i
i/xjZxT8hSkVoIFpFOKnowh6iOdS+Px9oEldavZ1tKFI3gVjo1mYwYAhgHDq
nydYGZKCbffyyXfwepbwqOOJDhrK/uktyPWKVqzIfzshz25EvXXsIbB48i2j
Hgg6e1arrcVuny+ZAsrHhHVo+njC35d1rVH1YFSX/+tkKM1muddOwAGbIG99
LQF32ilnshKAyRDnruPXlrZaBlvgLsSQPKoM1zBEFnbjXRNrsEqmD48hRD4g
vFEXfMmbhX7P9Ju4B+yK++Z3KRoTc3MTUDP7xrhIzEwIXQhqe+MGMisduiRP
fWPrl0n6Topk3fwE7XLjslMrUEbquW6aIrMZA/2hH6afH3IgmOFEID+aXrlO
i6V89Dihl6iRx1NJeHU2aNU+12J9rja8LTwaTbAzZ/kJuzDEp4rtB6RLBU6h
u9KGGoIa2x1itI9dsZpm8qcZ9q5xpsXaR3Y4vIWd5ddbDArARWa8wv6KgmrW
lBLTSFGHByXlTgJxlBkYyG27bzfgcjANMj1Ify4kqNpZt7Y++WZi/M4XKu6K
CkYJMn5TPISzDuv9ht2FaZ8izsRmxtSMZi118ccIatOtZqx2PuAzr1n/mC1D
3R86T7PnKGNQ1my2f5tnDyhVbT56su+2Hmgus2oitL+7iexvPUUTlCeUYj6m
2MpjxEs36kjv6zvsGN9g/qe/p/imGGpUXtKuXXG6LjGq1DmAmtusrfKF+O7g
mKsuuG1HfRbEbEL5EGAVnblofMzipF5xWQFStSbjAp9vBwkcTHxBMntuOY1o
xPaDwfcr3p9eM6wm0yYK15RRjRphA0TBZ0g+JMD+RK+zJTT0QOr9LcWypYqv
MamzqLsxQIpxMlE6GGpCcRCD6PdqCWlMzs5LA92d5mXIzF77YOm89w8MM982
vrEnrnDDRW7i1rwsDVBYnw0FGdhSlqhiiajMd+XUDO662nbm4+DNaCRECUkv
CurY+glVbqZ5aEtrodzqzAykRQ4hC51V2FNPGJxPez740InQCG89T8mSBmjF
NUURH/dTqe6gtzDVjO/PWAW92maAijzFXrPcGrp2Okfc/RIUgkxTXbmuVE+F
V4XGynsZ5l5HRtAVZu08M/p7xaCe9wgtrEBEHp/U+TSkYnydZIn9Y+HULE8m
PSG2sGj8yPavfASiG9lgj8zefL2bw1wxXj+Sjv0ujfnoQxl+Qiuf34vmewgF
oEqTRbqz1I92k8i2KV2P14fSuy4IQWZxmTssdxVPHi2EmvSQx1N6d+biXRdE
+irtKohCHa02sz3vM5YwQX/EeYbdtQe2+Wm8ci8i8ak3IxjlzkQnE6RZqFuB
NlVTC3Emg+8xkXP/CbzU5BF81bSuPj/uks9+UqPCg7e6AijE/hExp1L1rIsU
vjiRXeeVC7ueoagvaSQOJSW5IBofkh2Sloa6iIz65ueQXUe27ERsRQZ6XuRv
cPUOM6XGb5e2vW5InDStacgVJC2SVOs5CsSOl/booVjlUtVB1GpoYTqUyDYQ
OBMrTNykYrddZhl6d5LTSY0g5LQ0PLhQ+H1HP23RmItt89K0I++w+Ap+N/Gq
cB/10YFB1Sf+RizYZR+CloN2yDu9ISUjOO7BjAvXYI6vHqivv6fc5csDM2Pt
UzSAkQU/g0jzTdZ7CbIcnAiWiEc2Xd9GxbKv1fv09kSHcCacPHb3/V+Lhq6O
lCfDKkGDAoHvjRPLdWSMPAjRfevU66G/tpuJ79WeHz9oznTbMB+etGsoV/0A
ksNNs8IpI2I1y9PTKhPiGHWU7USpnurUji5o6ixqEaKcb3pYv3dS5qtGG9rP
WwhwmV1blB8omoxNm27BZXHxTDoSalQanGngT4XEAZXc4QPeDiVGSOsChcta
qOaIj5F6peNlk1MNZQj6nht7ao5k+67k049s+5+pLy/i3WbwB2RU0p2EOQUE
oFzZfDA4SIyr7ntoZ0Yojx9DVqFHCuEImlO7vs5XM+UtRKv2kIo8BfwVMELH
eW2Hwh/8+hgPCSxYGSzDnzFwcK0gHFgmV6Ro8QXl9r4UlofppZHGdObOLUc/
63NKTB0Mi88tajgDAmrY6+2X2l7ktKSnBBV/gQORGqXVVE9gmqA/SVfHz+2F
ziul+TbM84b+XLEXNzttLZjpzpZqYOLxPtBqUuvTKACW2H4jNga7oObfd2Ph
wJXakSGpot0veYrN1u+dxpFEs2dMO3FhWi7p6G1jys98Bm9ifAbCalhxCuKa
6dQZ+P1kC2FE+qQzsBZzSFd/k/txXQ1lp4JfKfymp6aiwG3d2eaGA2jl6Hlf
HUMw25ZxZ9RvO9XmKpJ2d00HA8uuGwP3IWJ6q1zHGNsFWB8LxazffPiXaN9S
Kca99i/YBsb0bEKfMUniQDEMU6P6eUj0mzMnmC0yrzKUW6ojmhE20xktj9Xg
h9AbJrYGcj6qE2X5MjjtJK0MiQU7K7Mc1xkhKNDCJ58PK7hIHHoTTmGBEXMC
IzQq+LIIZVRlbpN6Un3JZaAY2J5xEI3h/o1PLRvOCi3m0OPiBmC+uU4Fdt1L
bC7/RvxhROS+4xWfn1tHRAc0WH4zUlVwsAgosLayNjslwW3zF3L2hKQTUGex
UOVsgtkIr8JBWfG69QO51XrhNUb0Lb8Kaqf+MOS0Nm6TPVxfsI+t903/aW7G
U+u6h9wRuuHUXTh+YYAhCrTujSAeLZRuXuVlH9hSjY9woJ/A6CjF5TGlbZtA
ebWSNKBXS8/DY8t6hZZ5zOFBpO5gBa7Wm9aZF3gpszhyM55qf6KZMXTdafJG
0lP/fYmSFd/6pes+ycV+rjcReVx8IhhVaOl9D/RJKy+dIx3O3M2nVTmL676i
/G0W3nvHNdZR3BEeB98AyW4/iEoFAGL7mDHNFGGxk7vJSBpVzqMSGTt0qMbO
n0T9fh5ddQmlgZ1ehGikUBVTNAaxSLUHq+eEG2bVxOLuee5usuaYSnmJuNqA
BtPD+tlCWOI8C0uw0Ysgtkar6BdL7h6t/JYz8/JUDgzmwDlFQNkSUh2JCrue
GrozY5WuHnuT7i/H3zJCzraO5qRqALU9B+D4uA1R3DKwkFHE2jNgUC70rKdW
ZwXnWPfe6K9aLi2QW0W2wwB2EZtdA8MIlRlHrdGfUPxP/suK5LUsw1h8zDKQ
It3OMFU7xR2tAXf/w6HUlEi4fkbulCuqUoVCwF0RPBtO7Woo7J8+cHLxwh/8
tfQbSBRL+srrSVaUZ+qPfoMvGyyNW964QbzQsL83HM/6+Iub1lIijk2iRCiQ
nk6uav1PkytifnKvLNXGdg8UoGpNQSE8bkGnsnDFYGbOioPOmaoQxCnEtrfp
BLE0958wvrbJ/2oQzA+mAfkcMOUPT+3VNbLOpU9X6ooUuLRzH9hR13WNikSb
hAOhHSagMqkoUl49i+wjCrs1xjDcMDw1yvybxNQ9a6SiSk2Sc5VdCNHmBFjF
rac8bjaCO7MlbRWGIPJTc9cFqazseRaWtdbdwaQGLYdDFvsrJVhhlTGgSdFR
ph8PzEadaaGfhqYGWiliptZDxTeAUUL/5Bk+qzSJvcXn5Xb0o/JNSF72+8rH
AIhhGoXwDGAk+kre8S4Ey7LIWKXgCJwaWze7Zp4I3s47Jc3d2yQmtDxe32hN
LgF2HsKgLWq+7OEHywfxDk+If819B3qQsS0iO9uM67r5py8jZheITG+O0ScB
X369/yypFmiHzw02UmdCsrA7GpO/FxXzvUZMAewwSGrXFkK10JDyEb4Hy/5z
5n5/3pfn6Hjucav1MSzMenuFTVhWVpfMSvz9+rh6pMvTObnbj7t+3mWqL++M
d8TV3Y/Qv5Baxrfo8WFS/8hbRNU6UeKg53i7+ijGHEUrLv40Cq2RKzW/M4fc
p1IECacclJRwW4+DDIzjwJ5ROKxFJ6sTIME9NtAe+JOntz1RNvkKj+eztbsG
Qa2jePdSvDJ1MKTAd0QDfyX6jZaydTZZEvdWTV5vANhgV71Y7/6N4JcaPWTv
CW/MXokAd5hQz6TAEZ4u/MQxjRHXyafIOTaeN5+jm6QBiOg+5DlqikRyFF9O
p+s/AXGsGeBOieniNqh1QEUV8dEWO19lKzJXVl8YY3b/0U9gk+plhXP/ObU1
cA5hu6oHbVkXJUu/hPFwRgljY6CydExiUmEXTUZMOEnLLNFIxuoJ5K53MJyZ
ap0lwqkhrXQKp+JnxJSyko9NZcqUDAdRhT3xJ8FwLMwlXedEQcO3uU85XuWJ
wvU5r6I6R3qxHQGC4avi9fnJEzW9JZvPq7FQF0BXl1KECwwds/RuRlC1/f+q
uAEMx0sedNKiuiPJSSvXakitmXt95Q+2gagqosuK30OGpNSw0pbfEmk0wOxm
/7y7jTp0rlsLVopdy24yc5rC5vVGn9pUsoacLYoVUuPKc5Pw60Xi2kHib1gS
nqPUeuESStSwyhIxh4u8CYg1wm3uclx1XAiLcf9V13d5rneqtoB85MKb9Vn2
qwOcFetOP3ZGy7mzxAm+XvYDibRQ0UdO1OgOMtWBJOOGhaaj9iZKMHR7HgV/
U/CyePlzHoRUzmw2uuHPYxWOntL6VAsngnI+4I9CSdMKC4oQN1xhHijcSJOz
FcHX4daXv2+Ja+A36Eed6Ez81E1jq8kbbZEYfI8UPRcy6IrkLR7JbpTOoR0j
ya2pRAbPdSLv1CgYVtCgoTDWWZqh/d6mOu9phyeean9N04MuvihtxtnHI82W
EFgET5XK6BZ7bUk9qNMrfMsBs9HRUyhDb/oyVskafdgCBCuKI6URp/G7lnn9
qN8IvQdfA0czHa58OnxJtrcdxwSxdbGVQXzQgoO2R7UUY6GWV3RUnpobqNcv
rnj0629WYT5wmLssZ6fJmvnWZGoEjBMWb2W1qjvq/k9Q/fa6ROxOyRkrjCo1
EskMbjuC74fcf/DU6Pp24X6vuOb+jhc0Ha9TE/Jt0hO/zZhoQrhJO/2pvvpr
VT0wtwLYm5t0pMOjV+MNTUDFW0ZF7F943/lF8R6FZ7f20EUiMLd8P2YI2C/g
j+20bEI6sgAY/5mFB5v5cPZpOSC/zjhexA30zCPjS9mmXQf0woS+4pprcnRB
L+/B05aVW8nQfnf3uGSZiet0bNDVe9HfYV8fUVRjyavW2MUVC6ovfKccsfUY
yMrpUHFMt08y1g++d8whD+IZezITK3RGo9QcACi7JJt6YycwpQirlBQPQktN
/UtBr3Qu2oWDHPbJ85tV4A5/Aiy3qmXgkkH+uoFw/dZc/cM+P0Mm098+u2g0
6Eu5RxwkZ2TVtf0G4ZIArf/xuq74Oivb7kCr0yosti/3We4gdU2aLx83JHVl
jhKtkTb+PxvoYi58TBU/TjpOYWZYG9eHEwNZ0eL67SRBOPCEr1o2tQ0VxzDg
LPDH2i9buzZSsxjpE4kNfZkqtmq5UZgYPcdchZcTbiVD+RAQF/eDNz8WJI6g
JrFi59moSXRuumG1DVnG6z5Lyp+0RU3v8hYJR7R3jfbva+1VMSGRokPzSSeq
iwaAbdnASGuy9LxK8RVb7OQodaivsb1WgIfAXFB3TNEstVdu/7CqKVmq86OU
3Q7YWWjiTQABbeis0rAEk+qtLoDvI/TGT7dk4f2GLcNMkL/mR2a3n+O4V/oR
HjCtJPr4zhilX417URep/0TywnDR/vF5FwWlVuWkyDF6bFdTUrJ+YfTWAdoX
k7Xssf46ICFF/pYA/N4Gb5dmFTe/yfczrLGSF9oTNpUIWnNmfVvnWjQnZYhK
rfG2jdlEOsNRWFjoMn1U6uOnEheMMpr/yX8saZxB6LJVt+iBDFVPsABATP/P
FkTixAevSJybxb03XudjMrHod5E6ecmy+bEfYyxZiVUC4nvrpUucROkDpbF3
afdiQpnuyMrjKhl2EuVf6/FMpcsR+7fVftkL/E+Jwvh4WovQCadhq53944GK
paFoPWB5197n5U+5YwQRlXDU7FtbzM9si7uGQP1QBV3z+43iBlvrrnq2FoLG
swrLWSwzbIbOjKmDa1zQdYx+8XqE7LtOvsp95mRVcXeZfCGjJTp5olXuQlmn
tqbnnEhzwe8aXbf+r8eb6Ivr+E6Y/w59R09vuZtGsNuhtqSSU+MLd5miKbHC
TpEH501yJp8uFQbiSvuzRXunnlNH+Xrw7rpGJhHraepleBuM72NE2+L+l66s
xCeNxnsRiOsEjF9QnKArR8m5gWrPFiiBV8NWTwN10pukXrLmujGk0lSq+c7V
vjehvwEUSjFI5WfF0D6tc8plLQ/ujiOSBFXg0M74+lk1W2ytr8SIaNHCOFjX
8rWAdaHGH7PTBYK4dDe78xYja7U0ZdBOzfvKiWIqWnkyxggkYQMcidHUpNfA
hFXl54rr5wO37mTFhyrv5rYVVFM9oLkh3jQkUnKYnV3YSE0riD0drDzlvx37
+T+AmRiyMijk8IZyuKAVj2JOJ2+g49KC6neRL6oRlBs9nynFCui8Xv45BZMx
kw8KEOPqGSr6HGfucJy7vCkgRtsp9MQd+gQ3T8S1W1ERqELGl5we+muoO/Qb
TCMq1LcFw6gA1S+s2cz1KUZn9dy2mhikcG/HW+1QnmC7V98v4zCxv/I/U0up
6llutIWeFRHqa3f+O8y97csbzGmtyPDQNRS35bPzhKXMpzisqQeUqYirV24w
GaAF2+7sVOokKbxlbQw5qlfMEKstSI/y9mvnr5xYpU0esB0RR9rJbTFNKu/Q
D4wRhEVBk40RYsEdn1GS1QdJ2STrN0ibYDYLb7iQFgNd5gQpQzqBYqa+j2/O
rDCdPRl3bSkAeDg3BwfCSWU1dniJ9HNl82B0SNC+WzfUE6HK+9YHWLdj/orB
Vpdur23z4nz0pW4/HAeGlOW72Kmyq7jEfBtDFq9Avu30ShHNT45mzBIuDZgW
brdklbHcLS9lLuGMj5y/r8C2m1TWeTDKIaq+TcVDpLQuPCr2qBQSbvfJxK56
/LBYgo+XqNWzF1yW0rsq1JeM4So3LF8KJuBRDv280maNrGOSWwUTL+3YJt1A
ArwlSEt/soD8zKli/q0DQLTT4CYADNuhjbGTJvzuLOgam31pYg3yE2J6Kk2N
fXl7hqlrHQsGNsG/knZ033OSNj5Ng++mck3boPL+/bn8knG3rxlfmKGFni9u
aoKV4Pv41ZDHONKpCorSEbudoGVId5AEZupsFRavK48jfqrcxjNP5MzCKLH8
kfvfTrT/aOSYcA7h7INlCQLTnni1XQUks85OHcXPhYy6tQyCnwd//x8/7aSu
9xpPlieolZybicoRnPPgAHkWlqAsSCXM78M5jh2oY075LU0DoPGFINYw/C2v
VZviXf3SBNKd/mDPsi4/WQwwWPZomtDcujhxlhv1zf6YDSPdtg1ckh+MjAPj
wYoLXmWfTpA69tNdhAdriSu7Vs2dqNVSYzBUcOCnrG6rhYrN4vVA8PzdnQgK
8H6uwZY6hMBlAuA/7xo6+ItXg0EvcaiVVNMbAYM5hTL6spUO0A1L4gmJaTIX
3fis0jnl4l2TON3P5AY1ps9QNsW7we36RQw19P1eKrZ6jozRGehwmci32K7g
Awv2+kDhvvc8WTzmb8RGQK+FJLefwyKTNKwCETriYdFCBKyHKveFaogo+G5m
JPfKq3mmLXwRwTIIAUrhdICPIYCxJi/sQG+lwPp6hhvMloGDJCdOIII7I134
IWTbaf7814TTP+GePWaWj2e8PyHyKKiv07+QvUryO2Xf3o30RFnWT2vuENeg
fLtqIo2cEDQUAB7HK7UtaBdCaPof9KZ2NX+11OmzwGHKOug18WUC2yYqHcO8
m8plNY8MnEob432pGHHBnuzwrj5XNMeIY6M0VK035KstTzOcncTObJPjOCL+
Ez8gkPST/EoIBHv7zaIfeeb8aZrosRt+onQAAoILnfxHeTYlrZygo7UsM/7t
ycjCTpTtytwLCjtIICaZGw15f4RxUogr8zY+0Bb7y6XOf254ATVZm51Hq7fF
8fg0i4Fm8a0WUA4dixHR2BOXKu4qtfx4IsuZL58OCJZLi2dLLqI5jNW5erR3
JphXLSXF3mkmqKYKIz5OXMGOhhZ+nvG1u0RBOb215PUPAXchcSuX7xsXmMcy
kb2/yNF9rc5GSGMNtvUo5ZohJXWfPRuH6WYnXUbfMMbj4ow/KHmk86rQQPa/
a6VtVKZVZp+fnUeztht7DLILOmA8PMSCdNW7P9O9Xau/gqVLjCin+SRwLySb
nK6FaSvJBMzu09iB/pCPAbXLSEar5zD/TKScX1X6voG+lfo1bjyENekai6eV
Zlm1RUY7kyMClsO4LKpfgIt/XRzh1zS4Z7I/Jao+JXRgMR6W+hBNQAyVz518
5MX2Th6KYaTezYLqteiHXhNKEUjFjIDuxWRaK07b5odfQPHgCGBZXR4xC3td
tjXRcT+teiOvyX0GQElWK/fJ4ayiZIiHjDUvfr6ZN+FGP/+Ex3G9Y7LrPsqx
B5/SsJNRZW+ujgiNFlGWr4V5kAFDdRsFjSHQGRDiQHvyVmofhSSq3eDDWVfD
vT5DcoGANmverwv6Fegm0VxzWwZhlZ/0kjqpZoHDr5AJopcS6+cO8GytAbHo
tGqFC2mYKFq7Ff/xME7dP0ZukN439BBk1xifBzFRz2r6AX0aIKQtdfcCfPbQ
aiRbfjc26upMmRlExud3ScW7faYb9zQ5fgoCZyBXCZVbgcmVhzZeS8UuUPuS
NI4gN2J/0QyD6F9zAUlyEsJusN7vuUilCG1MALJQTSgLCiFWnItX3q+WL/Zo
fGGhQa8lbc88kuf39wHb6EyQYH6H4254XYjdqZDbpAbc4tauzeptktZB+NgT
pofV3qvJYoZl5udJIsTGUUe2mze2s710Jve0vj/NDkhtP9fov9UT2DPrMnsr
H8pxyiIe+bgZ9YP8HBIeP5wDJ8UbRFcQ/8kaE9aLPwbPN9psGsmdL0XHvZN/
zI/bttmO6h+gh0NEWk3GhM/H79k7Vm3hrQx2X0gK+Onzoe8ZQ1+MswbJuWz1
9ylJVc+Ybhg51a/yzozgVQfToxSbgAByKnbveMLO2X6gAzEu+Ct8Q6qNM97B
AKDfVLwtWOeD8JKBkklskZtswBi4j0wwlJWvVvS36eUbHHfCPEE8wwVAhhGJ
O81w1WToDb6gTjkusoWAO3V46tZDKZnfe8BNSuouRkUjXRvo9EluY+XMwpuE
hSbilfN3uCSgEO56iuwRFJTeVmJD7DfeNrKekx4lueoFtN4I7QFVj9BmvLOl
AMMAtWrVzl0GFqvPyDFu2DXOOz97SLESVbydFWGeAUkQYob7n+s/G5SHRnNm
xoJyQ1umb8WcDv+cVQS60vDFfL/WbXBXKfVA9B9vjiF0VO3Ys+N5LuEwfg9b
nIeG8ENRIkfrPyDQLzuTVn58RK9ZZownb6DHdmlg8atmllphTGJOn/ZbLiJx
keq3FhcwFbPDgh0yfZrvIVaiVT53ykUIp3q6dWlKJ5aPiIcm7koWv9/4lhXj
x40+jeiUqPYc1xaFCkJpZ3/knoYdZ5eCcQnnM2w/X8gdTMm1yO6IxttcOXov
zDOmrwissRL3f1P45lu22X8zpyIDHjIqgDwlHvJiczgRmehYeqP3UOKgueMG
pdqIXbO++84NOR+/dx11RrCi4jOkArKkoZDOWMx8QraLPQ60BcKjYZokOqC0
SNG2OMbQOA5HIdsbd6nD93OSE2isuZnhxWuxvisnuAUoUzVuPsDWu4gwypeG
tvBWuKaHpW+1GX9N2gTxIsBBQYVEjRHRzFKvUCY+TWL69ATIOdxuHu7F54/c
tx62cUK3nwSIzj7abUFnjwdujjP8TOeJ5D1YKSzHMhpl4R5PTCatZvhjatfm
5dwt6RLXmuPYdiWnAR4Djb1P+Vyr0WfCFgM04Vjp46AIXC0YmOaCFNCtsqoe
9vbR2k/t1hoYrsKz9/lIMK2V/5TYFcAftN50t5JO16fkDxL0aeKstpRCqiIP
nY039RxWZFDr3r+QX7/S49pDR4qf/ByScTfHFqAhTldsJTmRnzeoM3cZQ3Sl
0wqw+IRvr0smHwYp8g0Bjnm1eMkZIjNI39INQ4FczQpW1mg1EBS9xnFrzmzr
ma2t1Yjv2pnAg+Kcv0ETgDrkMx1nRE3VrbQ4Qxx0WdTLZ8bbDKaDYFQ6XPGA
xfqyBXejEOgtn7Lehpw+xYwWND4ZCSbRuyVIY7dZAKz55JP5QmsaImOkdcNs
Y1gEbaSvru2B8DkNYi+J+NNWLZL/8S3Ao/bcnxuWul7Up/GjSaQZ8F/xp731
5zdEHwFNUI4TkEJlMFsrZA7aj1MPP0gwbcNsAmfdnH2WSY4YhgHqPL8UQgWa
gNqwCVS4JpOCC22fZMqLayZArlkCbsWxjfc/TPNfPUioOtQZyz9PmuKiRg+x
1Sc3wDhyxF7TjWPDW5aJfPTagbpyaapYeHSX/vkd0VTDrLJer5qVNKlDIXJx
Ak2Tv7UzhIDTgWu6Brt07BoQdF5itsgGzJrhD/kCs17MwkrLyJRuIx67MXH2
hyHA3zGl/3cjjHv8CIKiUL57DZD6tVTyaRXYCdiKq5rNePocH6HRNHIjbYjj
SEHlftxFJ6zRKKSrw12GTLc+RznxawWH9xFzYFJEOA4sKYwViEzlY+Fjw5ME
awUHwMLRaVB6hHpIeqgawDDqs6G+yGJAToduQF+bQ5ybVlkA1QMWS0YMHky/
0kKhZhwnA+nntX2LeItzqrdqqYNAo1Hp7IiJYwsdQs3bUQ1ucz+e7iEDnStI
bb6NgRsVHe0+IWqPf387WcqO+ThvuzyGD+PL2hxxcbzNLbUvnAOgWdXGhEeJ
21W8LRdFN2oxL7MFCP3lbVCLw3kqzk4VjLEdHCZ3G9TtH0THr3LCqMpxXk3O
3CUqJLe1XQAH9cxjkBmSO5JhGHM0w6WHYtigPJN7fT7ukoBO/wYtBXigniA8
exXHuuDqHWQx6kOVT9FwphQ25k4RV1IzY3DbCDhkxolvvCUaqbqog7TFtQrz
Q6bWXs3DjU6+h3ZjBPl80QpGAuphvcFWcH64NQHWjFhaQJUl1FlUiK7coFbM
KuqOYQTCO80YLsmcO96d+Z2N1l/0L0sJ2QwzVf5iRMke/7XaMroWWKEsAoVH
ZgzstIK++RprjmgQVWZgaAr1s80hq3mkBZl6fzIy5Rzu5dQhmpl/agcYdWRW
fk198Jz4+iGlpgJuCGdaDWw5NoylCLSZbuLCFJoNOsbh7XX9aIzgrIIdVUCo
Bvupwcecs83c75B9NQxH/VxlXsBr20odBpagWVzXbRgPWz4KjnSWIYtGytju
i96OHUdXUIwsebE9xoY/hRj4VsO0cEuYRPHJ2ANWqacP362XbhS8dN962waM
43TBcfq7GpnltnnGH9+KCS3OlQUo1N8d3+FEM4+Nc/RG9DnCgFNOefAGGc1c
jsfYDJu5fbAWxw4IvJB+C+X7WtKy6JV0UCLjzNtfL8b7ozVTU6MO60+Nrygr
Gwai2Y5+dw8fbbH40/dK0Ob1SlyBCz7Ovk0MFQWHPprpqU9pMAT0iCNDylRq
MzQL0P9UuoGJmY6zYAeNbgbwtJhsrx/TIA5b27UPsQybS1Ccf+C+67gyw9r+
XsCRcW3X2k8sh1CvtnZ1frrgaNhtp7AZazc15XZ3T9oYHIXswhRFFA8fxTmU
dGZ+EO24aHwwNtKEk/8eSQeIKbKKLvSEz3eRhHmXvTslFY4kBaxZJ/cK5VHu
TBCj0V1e5gDJuf6BFXAYLVBasuKQ7/pipc9FJ93i0ck4gp7nn/ziR1/7IG1n
4aqw//AHobRfH8mTjKg99VzRE80TwpDN9Ul1skkxqkB74ArFSB90aXz2lIWl
l7I9/hMPMKNnTMseQrJOR2k1svzvHdNKdZWRWXuKjtqdoZ/ru1iifMebAtgj
H+LSXxn2TbPAOE2KRYqnAswyuCPJoVM43NDVY+cq63OsMgvbxsrSkk6EzVKS
ckZ9PDjTXGmXJk0u3BzrWHGQA7e7n7ij2FKTkLsngm9XV6qtgO8qqyQOJYOW
faWlj282JedVOfcPMDiIVn6iVtjZuR6fLq/fCGnjnbbGewYZ+iWzSHAOrT4T
NJzceoC+R59MEQkRlOXGUCNOyhk7ZhnIN/tuuUjdD+sjTUt4XoU/k0uG38sg
QT18qlFHuaj7Zl3LQ0aN0mnmOuhpoBlRjw4jdfWenaRvKzr1lPJcn4PgUo5L
56kUBnefRR8E4/0iGTGlpPC/H1s75bB6yeGbomIWs9otmv8blxkRmzmXrNn1
b7mfVvl3owIEoAIcv+r/5TOYtNqh7pKpwo8oe/0EfyrL1U2Vd6C+9tpLICcs
syRFUANP45JmHwUIPPbXhxeFFOTYjj//6OQ2uGu/YS5yj//mq00+gd3xSJJW
ne4uwHmRJ+FFC0BlVL05q9Eyagh1+XByZInCG4vDz2JBW093H/HzSWrqoHD1
nUsJYEdW58uGYo11MSc+5rwXRJQun0c+9vk8S9j6zM7xCe/iifP99QgDqyBI
jeT9zqITGUC9uyn7Scas5Yg23E7lDld4NvMh2hUpf18Us8RhUEA16axKKMIe
UXA+uQM5gtS6SfKhT+epH+iYRHGKVhLk6K/hj7WArK2bba1hoAD/XEOGRxgC
reS/fiz61ahNlzgEnoihb0KJy/jVlZJiIlXN6agt6fOBVaZ/H9R1lT44Sz6B
yRd6mlNO/un3i8rGZacYuz36tVBqf8FX/H1PnYUfn2QNAHSsfEXaAX+ht4jD
MMWkVKFTduxLmqksD1WIZKOSx+t4ScF3tRh7pPhUBIwaziHUZonI9ZkByBWV
0UVgpAsGhobmtHfP1pKr0akJvlCd4aDErjGBS96k1+4/kMRukccBwGp+pjGm
iGkFLYVNfWTfFpTScv/NVTZIoVGfsduRklYP5XhWWnTUh/IyNs5eVO6FOuu+
vYUy5KmqAsFzicg87doNc2QDdpFfYx52Rqt39iG7Sg0vkF96frgbmR8Sschq
EH8b07igR3wAeZ6ji1B0l5vW+2KyaKErsZ+s+Tk7Hc8VkTHA+MXE703rfh/5
6Xp5YaimPSM+YokRWSzdovJWhpHRPcCd9HjpTvnhY/tQzCqD3h9UFJy2GONT
+UeqvTw9klHQWKFEo4tUEr1u0JLAy7/kVyJXOKQNEQ3nlrbW/j/H8XPVjPjL
FelWlGK65do5R7LV/NwX1E5GpaDgFZDuODBNzOTxyhTtmfpiFU35yIKa9qIF
xXp+Aw05VlwDwe4jTeK4Fio1clUOj6H3+yzowfDJFQgW+u6XWS5amz9MriOh
oZtOX97XHPnfCfg8fMf8/uv3k/l7ykl15/X1uaMW1AH44raTqFnSxQEnh8mI
pfmN0dQ3Sgd27QVAz8zXXVapXyo0iqzxTdTX4yEjSTNMmWecJmzlEtOOJDBk
Fnl+biUcEIgW54H4tXTALC7jUF3Iorkr3LKL2qR4AhrggQvntP7eh7W4ut1i
iKgaNFUfPt6DJiGPCL1XrcrbLkzW0/JTwUl5RxKoIVTfbknr7dzNntsGreHM
30KQYw635iTVIq9tcFWe3LfQ0YBnduh4FMom7RAwWMYeX5L0SHP572tEuPFo
cohKLgWiYHd5hJ/ClsmL9iKXgaTUW4D53Ef75ZwLedabolsKcDYb/RQN3si/
g/JhbBsq1h+/v2ze8fre5nyeH93W79WUY0pBTfv9f4vAaICNh73DHCaQBfxL
goxM/JFZ26NifoAbfi8ui0DUX7I+L/B+B9YJEd91oKzSWBliMuC/b0pHJWzq
05eb1pmuUGRGd9UNtbvENsxgiyvgJypo/He2kq0c2f2Uq/lhesieZt0VH10z
3e+x+KEw4H87Cyof5DdALlUaAELNfvn69Co5+nXFBl9zaN2UUp1hs3JGHM6N
lOAZIp9GNp0JE0bfFKrImjAUJ1c80Q52N97zBqFM1M278HsUnVp/Hzduce4j
An0n9Gh/zb03KguTy6NQOJHB935UCOdUO1q+3h94xYXOYCpd/3FpjS+GJSou
QtyYFghUdDEB6508fukuIkCJB/6O2OaE27frwf1039pLQmeRsyoXs8mDcFYp
om5j3zJIr4xhuKjFKl7dURdWXymni5ORZj2LD40O1kfLJsaN0RGyYXtLTGlb
e0w20t5ZtWVzsDs318wnSCqUx2L9d9ytRYpUJUrwbm2bow+8MPNKNLDL3R4U
DM7jbcN0a/JZOqCeDLv3I39XVYADoU/5hlrACqs+5ca4aAniPOs/2y17pVCu
2pdbnq6opiwFWPVz+sT4sXKiHxkw8kMT5zNZfBIcsKEKLDrX+WSXjnuNEQgP
MIZ5NFXMb0Zp5SmVGZOSZHatKTqI7gwEfhXqqtkmcNPUln6SAT/Ws5oQEHvD
J5y0I9XYm9j1GJRP/CSZ4fix/qR9a2K4LyIzshRhtYVIC/3XQgaAv3YRJUOo
SILD19NInrNnDunf/1HNUF1oZJcRaINGDqn9/N/50wgHKzC5jq0UrXQAYJBX
RMdQb0fsLaEL+LEqYoabTOAC3Mb51oy4UEnT1Z6GuyHW6uZVHQWaNtg6N8+V
waO2Hn7NAbjJLCLLNrIii9Et8gGoNmujsNWRq5MjwxH7Id1TzlAuHTDg3H0K
QedD6jtYjk7n5sMP/E+cgggqp634ddmaH72G/AMI3G8R7SJl+wbE6jukFaDI
ZmVi08Zt05xDNsmJ38HivIOi/2JaWPuS+5G971AtrRxTSmd5uKYo2VEMcOEz
iP3nsRu/o6F5hM7JMXG8wBTUuXiqJJc4J2V5JalkonygTprK8Md9i1brevK2
DKRYnXRuTYleO4VNiE5Cj3UDr3Fd+GrqaIOLW73pw9f7e7m+EOAs+k3vv9ex
M+YNzG2efsnq1j6Ls6r5io8ADsxcbZU7zjaV4BFTa47Sa4SUpx4vS39Wf4L6
nyibsORcFkr0xJ8qN8YShYXtQxRBFIBs2bFOhHvR9UwyU5bhlqEdMBIpzXWJ
Ph8YWZpo+Pa/rDGgKVt/pIF7WDkFt54lkmvB+dSg2knunIZYLcsJdq5azO8o
Ox+0kNM3/uY8zvXvGN7sfBq8yAbQwytOFS19mY1591m18vxbW6d9tcM+t9YO
F3z1HPZ6DVB4p0plxIZMLPECAVqzTSAx/UMjDe+R5HV/f6hJCeAe5c1KOyxu
5r3W/CDjZ/cmdHas/GSQwGZB3XIyYYH3zLefpvWHbZ/7kFAqhe7IP328FF8f
YMPrUS4o5zbYOAax9nN9phE77JcjGPEHw7BDGy3DFG0AK0YrEkvpWgbR+4y7
jDcFNijRVpSHgD08vavr5/kDhvsM/kZrnKCyPetadMW6BpnFhcc/tO/nmt4V
nK6M13n0sgaCZSn40CQHE00YhGSFi7HSJ7Y9x+5xd0VJtkRON5l6g2TaB2X7
NfVShe5AvFEfgNHwyk23qyGyKk49ecXzdC1AL5JbQsyWNMv8b00IdDFKrDdG
wt3NKC3Z0XIVROBjq5neR5D5ilzGp8oExV9jDtlmq+fSRse33D+848FLM0Cs
qKZykipLXnmSfOXC+P26fjPcu+PaAJJWT0pfoRsFiI7hpqyj6PuSP6jp/acs
S4HV8FmPjBxBBqPDbMoPd3jJPeH7T3i7wH6EfV3k0V20kC6A+bUQNCzEB66H
ocLz8cusLjIbqBseITW/QnKSFkq6HbPYHl1wn2N9MoZRxNYslfwTXGNZFHPh
Ogg8bqakz7k0riZGenq/5c3sf6bwjSFS4pBeWZvZexA0On9fn/Pv9MFddDoP
Tw/dsLwG+oTNcaX1PjRncITIoHlBD0f//8Q7eNVk2Igjz7XZDS6Iev8Q9H2F
l1jy3vnpQ06F2cnOZVnPSHnNGODD4K7VRazHRKW/1OTC1KGlPxSmwI+BN2qX
6dkdJAZbx+MGhXXEeLTrN4WYJm4iG1B3cQ8oEdVHuM9TF8Q5pSDhMCgjt6cy
0SyK+jrQW3hOuAHMEWKzf81srf6dRcUF2uBNohZCBI+qmgknS9hxRLc2Ljvp
NlHiPJpgQz/GKhY6yiRc6fUf4p9osHqy4/c+4LkfATHwp7I1ElmSgcbHUA9h
fpejlxHXLR0QxtUCOQz/O6X2kfGTonbaEx1ygHwSQi5itKgP/xL5kiuidYp6
KynZUjPkhslIkIc3a9SLa7my7e9gjv0eN1JhTu1GvXKT8dCeVW/Z07d1khAU
WCILP4E9mAet9FB9HqTGHzTAeiSFXqSEkw6XiNA3Zt0AM8cH31SzgTmmg7XX
c5+o3f/NlU+4YSBkYvHrx/2n2qi8/SmKGV23zJk1qRgUemqFw4AD1cVaCGTJ
Ov+ka1IAK7tUdGX4t9rnDkBSseK1qQQDUy1W2t3T4+mHKMnohFJ+tb871X9m
VGTXmFyU3/CRjLhi+NauZmwRHAryht6chu2ZscQZFiXrbcy5yYJXMYBLjaRS
On+akUuWcTRoeaQXVFXhvh9Io1Q14DhMXb7GYRESs+BZvA4+q14+SsQtEiyj
siapZ5/ZoEp4QvSVzSWBM+4qslimm2A+0A05zOk2hBIa72GgVj0xn0trI7fs
2NTe6BhUjiLvR8GglHwN/hN9qnMlM/DUyDgWx8HZQljA+M1/4/VzOZCjiX9r
1DuEbyN1f/JD5/8UWcg9h/7KBsbJBtRjBx1X+mBPJ+sUUPsOLzob+TNxdOKV
NbWg7K6fIAhuiNZ07qrQ17AFJHf4TF+KkMzdVa0IJWU8204tucbxzweXjwG/
BNFFtDxYcdHFtXM9Ib83NyDwRetfko4Ll7iPkJFKct21l2C8llF2jwd46Raz
178gZW6fUB9t3IEX7wX3lyPkmqRfNF9HbN+ua6LgN42KSWTjBdVvyocTv/pV
r0U/VYW/qN+f9f2YLMRWd6fTmtuBdAEyVTkzUixge+Z4bUR+2tz/E8HOG2U6
cPdxSwTbkmfr9KDEorBUCfRekcNUD8kLUlxjdBV6PwVgyVhMb1wuSeG2CT4k
mpyksAsEzy20vswvQMnGpeRokH0SkUcpJTGjR7vlhkbJBL2BVa8mb2aKo1ou
vSiDa4HV5yx98EjVy7GgEjAaRwnIZba49WvYU64C9wma5BO1E+FRYduOXqzp
ttPHHZrrmVZ5HQb7MdpSc+JJJIEQHK/QkwBy+vtaZdV4OfPWLNTy+EV4jtss
MqtEgqR/Cvold44cyyKAnzXTLc91sRWNix0JHO6v1V94iaOakB2VyEPL09ou
VXsbf7VZ967X7RLNkEqMC/e3VsyrXLQWiG4xEm5H+B+DPAlxdRVQ6+zo7WXu
KCRtPiffTWLfwFZhCBiDM81UmhoRSjlJ7tfO1HzBrd6kNyzloZ9PKLzqD7VA
ai4CUdjaCSnYVijjZsw8ron9lMzeYdkvb9Dm0r9XD83/RVkOeJu7D+QNnqQ+
X2/rSFT73TzXqQYpPnToS6I6OMRRB9OysMMn2cWoqejdh1ssoQIjGeESZMQd
yg1ADImgDB6VC7QoPRrfrd7Mqzw5uNZyHycjDQhWPVXuSWXJPa3LfB7tJhCd
unOpe+8YpRx4rni7MsNQSkJI9sAL3aThqFf5JpnbJmGvtomNvCJe5ZSnqgL+
D7Q2YXyNgKqbtWNLnhV8mBMYbtDnJCZ57fwbMhDYjQNMM7RWedw64zjUx4TS
S4iRGU+xuQhSXlAph/Osds6BoNn2SZXxerHeSJp4tEMXV1D2Ajm5+dIkLTnr
8NckAJ5qZ6409DdhAJfyKXJz9Z7snAnjxSGzj8DWQG/U4XtWKuKVjpP2haj/
gSqZh6oOXQeSDZ1DhZOV1RV2IeNptHjrIgCxvbJSZZA8kVU6yw/W9FH1NMNa
aHsmY1i8kbGWCBoIYYQjwV9ZaPfpdm/r/DfHXzkdVnh7wxPSxFuqa6DSrn4O
ktZBFPkx+70Pyg4rouhhNcazrmIqDV9t3vroh1hdNCY95S+gI5Rajku7ZWNg
Cwn08FinyJpyCEm1ct1tCe0OL7VZsC8+eZ6qFAc7rU1SJf0WE9RVkP28q4vv
aBXK02bamsd89OYz9O1dY3ETJLdb0cb38vD+ns4YsTiRm46baJFkSZ4uIOYI
sCjeTAeZqj4S//jh0IVm7k17166txYcq+222+k5o6dE2sh+l019KPE1JqrG4
uckZtyAuLQn44WUGuSqda8i9FvlTGyWr+ZnVY0NT1Aw0xKbCUbUzi80ITdGi
Jyk46B0zWIt2a7JpgwUJTmteoxCdIXZDnp0I38QWaMgW8/mm1HXzYRrIP6Xk
Il0a4eRwlNTOQZ9P5dmGjnWcmtxlehyzpRnyz3VIbxuZVMzsJ1GVqLSch3mp
gFdokRkNXjSTZ1DhuNkkouP4X6YTmSt0n5WKwDInFGkFC/UGtgh711SxJclM
2AQC2LcptCl9PMp91TVs1h6yNK6nU4NT5yvzqBzVrtFchTd6xJJaNtf+ODNf
J5CZLmxWemCy/xPauyyWRNWb1gtXGS4JeSWU0Xi9tJQqrefnJrmcupV9Kf92
Ts/IzHm2HTYgtmeCMMkcWNufUvLpPt5r6Re53VCPIWwwWLMYxna/jdLljlhf
stBzc+47qBI8gTxgZcXtF3m4XZjpkGM8w8iwMcnSlCUZCW1I7r/VUl/AbeSP
xE1tknBq1NYAdFef/dSd/SU8yOis1wcg3d0mXkW7oeZlrAIODXNGWDWfkRvA
W9YGgru3PUKGAq6FAb6UwYVoJqnipZ4mSa7oMSo2j6/m3oHcu4IV/sf4MlUM
w+mcCLpyPf999fxedFAPB+lRANdhbeMySdLHS/2HSrAIYRK9W4bZilAMMlIV
TJsXK9qJ/oSIPnTopApkXyz1YvsXo6IwCJjBHtz3+0e/TGewukI8xX7m7N1f
BqJkry846xozWsWxkAcyGEcy/eHR92RoRqQ4Hb2rbeFOFtcjawMDbF7eBV+f
uzcUe9Af0Oz3EwacTdkUVHaPYk57UJE87gnprW2oFeLEuMgmJarmqmW1K9yU
n4XXN3ATJRoqF3UZmPOWtR0GrFtRIlot5L76PMQRjwOwxfgVKobwR6cWYpdj
wzzcYw4+EMs3wFQRb8mEBB3SVKKf3Q/Ryh6UHq1l4A5mLd2rBguVhqLcSc8P
gr2OOWFIb+oYbpbqArkwmrggrJli/jtniT0j3t++YackJSM4o5Mhslff3ZLW
Ncv9TvVw5RYpWj1PWMmxA7+7OqNSfZELRmsTBv6Pel8zenTuGOnoaophxKMg
aEID6Wf/8JAZ4y/S5eZ8KzdBraBGHfR+9Ne8GaXKLAzGkLIYRXeWeJ4volIA
gh+WOZRPqji7nV+gfi+9j1wokpEAW6ecHk7l2HI0Is+xNdhSiwJbqdGR1jPg
zaGhOK1GydT07kyIhWJyzoS/tfqkLcsElRt0MJUup6AT1T1lytoM/2TzY4uO
H+pO/8KGuUtDXrdt9gZlMKUI9zCz8ZPrrtxoCLbEAXI2zy+C6M9kvy1AEayF
yP4j0SznOCIrxgYYT/sTJL60U7eySyqmL07wtqr4+C/Mv4bATW4h5N1ORH8l
cybf2frHVTiCUJfY7o6nT2K6m4KlNB4K66bUDxYfavoBMm8lgs94xBwSY05Y
cn5XzIIgmglXWZqpKVDulUguHLtpfRG871sIcH2SWYVKXRosyhbh3HsoCYKl
TWxLPGE4spIDVNcpFFPwqroK3HAyeoBZh88HTDvEePi7B8n0/+VdKGBfQ/Lk
hb88cjoL2xtUP9K7DZkpi273wAOwRGPM3LmuCO2vP5NdxbvimPc6eyFFzlO2
VaNu90QF0LRDyeX+mvA/k7xBGRD549g84YnsKUJUcohSmHs5KyRTBV2i821m
nCpAvApgQgVizPXbkv7Mj7hIk/2hejXuIdrRtQYAlD0t6De4MBenW0j8IkkA
qejnyelyPPgq+HxCT0QCs+saD0/15j8xxBXE2eJ8jh7ML1+efDiHiRI92vYI
H2GTNdKmqB4U1mwjsX5+Zps=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qQbZfD6zGrZ6szh62Mk8E5LI9cBYmyRm+TVuWxKVBJT+g0uMU1kzeaxNcTvuU89cvVf25sHwHy11/PetfPHAXz4qQZgKDRybOyCREmT1MnHHw7O1/sMK/ym18bWDtay6xD90m5pI6v7BaX4Jndn9VnroI1hgd2Pi4/sZo6TbIER+UN+FMlQSulkbNz3cUYfIVeYSiHSBXC3bB/fRl+y9ElTUfUbD7vhX4+5UOfKpzUnz6a7lG9CRoGgd695ruKDfr9NvLbTksHTdbKaS8Glr+b//7BeXMXivnfI3bo8++yTbtiqALRVZuLhZBC1Th5b3QT6S1/AUapgBOs5AIMkbDetm1PYiJqwAFff0eqjgzBNkFlDLR48ZHvj1S4re5tEbubelpQWN9BzauqGnS4NWCECDcyHJkfK0YVYJwNdMt2zTJAp5Y0bvlt3W+VnJvATlgxHNELn+CI5/g3ZySvD0y9+BwqpYxXKGqp+d920LqBzs8j88NAnQ1xnDHNw9r0OEJ6OxKU3HUWVprAZRcl74n3rreYt3saoHUGkX6BWBuDJqNCiSFNt/SU9n+a7Y7zNznmii0cobH+I9Q4hnzQt5453AmSAqrNOvO3bUDcMaoSpqE3Bate9KLbyz2e+LUcNrfKSPDvg/iHyScDTLotRXQgvmYNjiEBzPZHIsk/gXwO0tVwLJ4TjGP9Kj4408PtGJnrIbdkzh4fAJnSekEN9bHP2tQEDIXnRfYGrTftzazaqwDkMgLn+CJrPQU5SicC1j+BBmTq7cnrPumR7DtVVFn53"
`endif