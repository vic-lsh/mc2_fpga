// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UDWsNXzMMxO24t4Jgh6KI/a/ckiL88G0x5gEn+vPGETaeh6eAaLB9KR6+G0q
3jWi+53LnHkgWNz4RpVOECYk5Amg/aJ3bytK2f9/+RyNJ52XkBV6c2eWk7Qb
R/Ppj9/EvsASeZBb/1cYYmUD96pr1So7bhqksWhB8xB4ib3daGvNA4pM/tSi
5QH+oydTbUdWG9BwKU1zb/kgqRIkdo/jfm6zeH6T09wpevwYaeq6zz1NVveL
jJHSAdPymEOkGr5Z49pziGgt6OmQzVNIcRyFy2Wyxcz3jYLXxKGUolRTFaG6
TZlUe8EIfnaKQ9+03Y9kH0UVcjD5xTafKkkeuvCdKw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dt/7vpd5Ke6yJG5R5A+nQVuyMQhXdNpN+naDgV+dUMQHvh1XGMZEMnqE3iud
Q57GMOLcFF3UIiNKHHC7Z3ZxU7QwakxcOOZQNqAchKGLFSqCeZ1uqcD23Tac
3/iFAluykAiU+BdWeonwj+dkLO/dHhrQcIz0K34Zre3MStAAzweGDEtRXoHl
pkvkFbPtEyN8JJHdmrPo/m0hrfND8DG7qCsQjYQeR4cwe/kQxp8hqbgc95Zx
SzXnezqK8AfYoDwurzgzzcUn56KtA35U2eLTJXozOzm5kKeNHaarf1If3KUh
Fy17zn2+clsZe87xDrIvGlKS8N0uLrOpBs70c8qMwQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QQjRv5TqUrff0DBOXcocqRLNO2bX80kpCBlLdIftyBSLamqSkMD7LC9Hfxdj
9zOj3S1sKDVqsS5TU9v2WiwSaVXW0AwTiO9j+6liVpWUkD7g83FMwIp9DUeu
suh6Nkjjb7aerTvdLq8vrYOM8qFTExLsIsCA5/6Ka3DIjRKJN2GTPN9AlwdA
MMKWA03tuQyszpI7V4GkvZqz0V8TuiI6zElAoBJ+SQ8mRmwMLQ56wcuR9phe
/GBGArWbWj3y/0rH1gvmahh+PjLNDJtcvt5I46RCnAgsolj0t/ziKMfGIUDA
dOzvA61IvWde7TdOovBdpuGeAfQvU+xMbDti8qtZcg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SMGzhJKCgTiUaV4bla7WF9xwpv+U8RywESK844J6zq/6evAidDIBYwpfuTXB
xtn7Q6nqmeQhUF2CrjH+C6jr000ERRNo8R//Om8a416R4BmeodBTlypaY7Ay
CE7ROsH+JYkdXmXO183E+7vAUDsZCtu+2yt2zSVFSJy3iHsQtvSnjVhaP2qn
yN+G9eMGko0GBSPQfTwejo0Z8xMdpcaYQl7NQWNBPVnfoegWpTZF/4R8wXJP
08hW+B0G4mdvqUQTX0wtE/1MFm/3wiPPx/svSu96FGWfedU68YdhCtSHg9bO
Xt32tnyII8ExX8J0gGoo8HROb5rRmJt90NS2+KpoFg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m93Tols2ZR/wJrR+SUjPDLRH337nqFMxkxZ8Ol/wWSfrdjD4cnnqLDPLqLMM
wGiB/Ivfbj+JinEjEPboKyfQUZYzDdIXvfBLNGdUjn0jn/34GAlTRLDV/iA2
vGusSTSxJ2JpJsisYD5w9963yZcJEFa6A89tmmKjjMKrMGjP2tU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hMkhOFD1HRvfLi5eJs2LJlPWlV6zwecCwbE7/GTKcc6KFDKrEg+zCKqStNjt
ZgvhhcqUDhEjznLo2/DRf3ZJQFE8UJAm6kFWLjW1V6eJeYU9VSGPyOcd2cfu
lL7kOzjsdsQA1cY6YRitR/WWEGEx8+ytzmEtvUbxGwb+h0pDPQ6MVo2DEzWc
TuOrbnRw4mwhHE8Qkg5qtlWrE0U+NGDUL6mmcmcLbprpy8AQ7l+XxgE1tVr6
5IhSBABw+mJzZqAyhScgTtJoyxg72hJrj1MQzZHch8WRASl78CGsEEih5i8f
Nd0KFbF47oqxOHx1EbNsUlEwS1izNsaeoA/U5Ab+npnTQuf5PEs1mFGtWq6D
gdyKJv8poqIf/yKx4BAbDQg3+PhBFGFxen+58upbJGA30nLVMRYWrqQOzkye
1nO/RoOIVnTSqG8AX6J//T6i00+TqX20GHSHXUw0Qf6FGb7K/Vdg2Z9uIIZ8
nuKWdOs1+fEe0GxG+x3J3SkjcPg+n/az


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bnULmF8hYfR9DNw43PCfiNiR+m6CmjEsD/fDToxrc1Lyby5SclNQ9Oj9GHpx
5NEv76JbGcuzCIYUKboUMo5OQudAloxqmActUFzjQ8ooTt8TCB0aTtafZAsA
pIWK5embTPngmrXt425gypx7sDXH7vmkYESWObYEl8agIZGWrCI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UFNFUhoyLH9UwgN95bMexYtORmJdbQ3gWDn0Fvy3RJYyXdZ8Ym+zhDKz/lwP
OM1EXx8fvmmq1uEvMESmBNmMkXUypJbew78QBaoWSm7JW0g+GfolAE1dp49v
pAh4h/4o2T+DK+xVmkaHze8eT+KHHUMNUe13fbc1egYgniYPn6g=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6096)
`pragma protect data_block
dwfZnr/ateTar3fA67Hc9qe2OxXNvLwm9+anUkwODK9Tg9uk9v5EFcy8iPqB
2xi15Fiyl2GJLjk9+E32AOrbJXveny7500wdhibtQ8sjq7oHLO1c/2r7G3fY
Y14pGwl9q6cA+POAy+VVAjbDSEQE4pKlZazgD5QhPc+VIIvCtdSNC+pponpD
0f8a2MZ1a32LWMjoxvd0jmFyXTdbGfGrbOYTuxppRaMmtGW2/amvwzV7tDIS
Ktyxt3QP0Iuhd/JBJsJrTssrsjHeaBY4XNHbMutbAel+TOoqthYbu45Qysf2
ayJ8RsRVTVAVEYtPkJueHwmDmr/XnyuXAWFo27HVJPqNfUDm9nS4setR9QZ6
Fy21USszxDwq6JygpoYDJFZt9WC4C9feHlHBxrUHzXihZlSb+YD74jCjR3uI
ZH4HMExvKWorQUT8WQU+NYCU3DIgA6DmirIkPGaScnC/wKBDnybfUZX3l6co
DwGD/zhbEmRBUUgE+kEotiBWVEzJSecmwSUPN8nGibet0QdwzVCuZ7yybdXX
7qRftv07bM2Apz1DBc19idc2ZEwOIMlh0NtoYlPudQ8yWf+vzbx86v0PK1Y8
2GPrJ/LtF0dblkA+ccurwcpzRjniaaERxcFxD3FXRP1I5uyUlleoo78fuiqE
9w7EpYT3b2UNwtLO+iGKgthokingTCOhlt20lhM0wNM00XJU5Yp42v/oxAgU
xFlOoa6tquxsNK4YvGUoRwG9gmemwmY+IYfruJTXHpLcDnAOvOd1Oj7FfuXl
h0uJ+Nq77f3Y9mVNxRyfy8FCU2Oe/No9dS3EJwTgzvpQJDu+hkXotvldVd5t
88EDNQfKm3vv5t0ihX+jDI1s2zQTVPDvZ7lcIaBZcgk223JZNKbn9sw1fw6/
MxJnxrxGrRSX+fWHhfQdcT5x+Khl+O2Gz7qJqv80Sv0I7k1NvlvGmYWWrZbJ
WGl6csUPUIdlpPw2nc+7PSZxYv8Y8iLSqyars/IEavPeKpsg/46xe+PBaAH/
CRsCTyM35wqbq/swxgDTyuyFIuJp/7WdnrJxOXkEnA3bPEnQ8RyWKs3nnVqv
m+Vjed81y2Vr6JQ/eKrQXy5nrMqtcJv/m7H/igRGPSef9b2bJ1lI4EohDtBx
doxkrr8JPq2dViifeinWJ7YNgMZvzL35k23eBXY2zw/DaSOgdIN0Mlw8bS7l
e7FhgkPdPC7YuyANzceLu9+kpU7Ivcm4Wvs2tuljljkwCsGEHb9pI23sb1BP
npB0MH9gaO5j2X5q4DIsI+hQampJrhN19mrxYumE5DdfPBGpcHSBU294Vs3i
Azbyf34ugHeMFtS9NNnnuTaE93DzSbvvqcEc3PRXRzzPdtLrel5blLBpDrbQ
JlSjM/TvXRFvAzsdkqWLNQHEVep76kXrBwtZnKHNldQqlg4zWo+chfIqD7ZX
nYC/y91kgMwySmd8DQ76fkzptSJIHB4i9BWc4O6eZ2jg1XSY0U6Wk3UiLwHU
0vbF/E/mgwm3afld069DgPLkElOGZxMpLwiv9vb9EnTmrNXDERRfLzMnM1qK
pnwmgRV66yyOeyfE2oQTBQwc+nfFbeJV4x6FPoE5rIFaCOLV/+z/voJgUelg
WVaCa+/FLIECiwMwksz2ykl2HcHzNa1g1T6XbFLNXZbqCyvM/Cmhqbka7Cpa
YAeUlPLnrVXrDRyb8pRtOM8gW3W6TfNCOz4XzpwTTNk10yHRCx4Buq+WFDsK
BT/dO3jJNeleNWfF4jB274uGPOQQ8PAH06vY4geP99ootqVGhBAudy0eRZhj
x+L+RwvPy00dKoqdegx0PoAf33Jti3FSYnD7v88mY4A94SCscJ1HbPwb0QyI
+M9aU4iPMfF4d/TqO/5Y+g0Gync6d8TlvSI4+eKHJhbWKbUeu6Mwelh83HV7
HnobS5zECdl1kxJMkoXsU4v2JanZCJH5Pclxbjq9OfmO+tASwc9bEP2HE5do
3WpZXVbhoL7lLArrVnLmgcV3FGT2+XzoKSYFusz6JhT4km08XU43ITqRO4Ea
roTIJWxf0Sm6stBqleWzjLfafTT9+ody9H8+mjaPaHm+An0124S7ru+UoOVs
ht8LDYM291XUJXtD996oWezzxg4E7gUReeWIrFIHix41t6tZeD6b0Kgalm9C
NCxFDHfQumCqw7yhYT7sHjnv7FjjUUotu1Ldnz46JscaFPsqv6AiFFHUsueP
3mp89ZO8lwOFcSBYfFq+cjsVW64UGRyyt2cuHHmGk+RCUjZkMvedrA8PfcCM
ePXA+BJVL6xwox01nb+oyioHJvdwUCBFrytnTQah7MNi9BlI32+6WHRKzY6S
okHN0fuW1qnp9v5Ya2cdmYMgz17sH2X9KtGH37DoN4xnIlgsxLD+tp9WuraG
Dn5Wu0XjegUJh6tAeCBEc01DzMO+3HTYMf3etoc57mVW1vdhauQxGRtqp4Qw
aOHsQ3dOLaQ36jsA4IIFwYvnyHJLgnVzskrq4QTAE9Tsv3f2/HjN/20BjLyB
oLCLminHpT5w6nQhUw6jBfMo3Uqd1Kzbtgp+houGdr5XLhUzLYQTNT9GnFbh
OyoPX3HVtiYpGgsrWjHIz+BDPpbbluj9+rmu5K7bx9TTLK3Xz/ibEUAAEXBC
L32ml/yOOiKY9mlCxuW6sdro/2VTiWNYkX9d7qXZqBHNTGjv0qLbZlpXhZFd
zDhYzFhZ6MFZM6rA93/XYkH/HmBOwSHSMnZ+Am6xMNNMEzbfdQC6QY1GKYWZ
gmfP+YOnjQmnfIZT/DKoZCkGjzCtwb79+5OdzB53UYQNPEA4RZNpkqStoEcL
ZA99ptvbw/jq0tslYM9EVfZJkpJy32eHS4hGgD1kxAQDO8SAg/xZnM8YhqlZ
G5838AJ+fjfia4Yrn7Bn12M6abgP5Sf2M8OAa/ydMd+XR/9sER7iZdrBUoJt
FDbVI46bSrW2xDGQCTtEIsLBRBnbNk+If0gOe6jnSb/njGKY29KM63nk0g5U
LyF5K3sXMw02bzb86QKMX37CC2qz0ByfFHIeX75tqM1J9lkENAQTn7RJoElz
PvKb6f5ilG2MkRxGu4ewNEpCP3h0X/L0o44OsMNnMQhr2T/Gcm8sfWZwMzvm
PFTtzJ4gtntH8t04mDISycxNuBiswyMpk90BeaOzRBqaf62iHefmrxFJFWnZ
IWql8NE0oUgFo3ei7XQUgOFDp8cJXYLfm1yGjs+rzj2uvxh0tbdxPiWKMj0/
0KC3HOdQTrfl0ahgFX7GXbrqQEC71vj4iYBfGFws2w9wpVgPw1tNXUdqGb72
yqXbaK0gZKBQBGilurL7uXiC6QFGM9FQo4ix1eL+9564/5HXMd7pEQmLWyOA
QProXZAgBCtJQ2/MnnzLhwLVThzKuVLMLCoMj6yIiCAcZFwIvzRoz2yYPUn9
mHYihoAs9QuSrJSKcjbUoEtDZDTQqWHtV+g/qLHk2+9waOPDlxKJzIz2LW2J
Y71IlpRoOckALAABeNFNNLlkz/1vQ/cnH6G74Wvs5bkLeNAvC8nHZo/hVTqX
0h8wzegpkhFz6PmOnb05HpMP/FHpHDtfFxIpCC7DZyS67BMfzqgNyivciHLT
kgTeP0+gtlj+l95g2gF9CnZYtN4aqzKHM6/sLmf81pf5lV02iaD3Y6z3Li5m
31RTPHQejTPUw3xuYlmsqyeng5MjjxPE+fyTJzMQC33+uo/Vv0ZL/V/LX9Kh
kstlmnvVFYYwRJ8VgYaVNTYoRdf9S83R/VoNq07MgvWzCZ3WyHCoi7/ZXXwU
zIIcJE5NxOwtH3mR0Y72EhCeqdqEQaR58vIe0NUie9zhoubN31MVqBtjnXsD
1REvujtqCvAJfHpEwEbCA0hYjRULvW/DZ6PnqxlyCbEnoGNxNzpFJn6JZabW
3y7D8TtmEb189izibw0TAcncEb6nkovZ7dKn0mwJTj1Ludzt47KYsbUd+Exl
9kfx+AAHWZt9eGsKzZBY44b03iTK4Wlvp9J8cGgStT7FawxJuFkgpnfdSdxV
WncNc8jav69Oe/y2qAQh+QV/7cig2188e7d74XcN6bFhYGzLMUdHFoUUVViU
ucfriWH9EH192xUYNmFnRwYAnSvka8QUJY1uft4d4C3m9J/yVVOWTmR862Cu
HbjlOdK8ilw/W4an3QsfWxw46zQwODd2gsenFAfs2jjiJJ0H58hnMvZ56c2v
kchRsS7QNFeaf/BC3J25KP5wBJJJHG56yxkh6AdLdHS2m9ZrsgBx4xVIlv5g
aadnP3phaqNhx/HiF9OMz4ubq+rtO/8daivvZ2ioBmkxzT5Up9+ESpStNyOR
5MgXsfVLZ8HjNKe0F0DOvhFvsWtrynD002LJ8SlT6T+RO9tIUygUQU0rq2lw
W2ZLcuVJLP2R8mAwKnDvs+9jtNj0OEH1mq4oyTrgHSr/PmCuEhBMc5pDQ6Id
4ibhsgl6RCYLtt1uYyxH/qDJVzrMbvh7G4rYdKu1Tz35SujtZUZtxg8xD6Kr
tTwj3KBO+CJwuHQZsvGYrxmBnLOEs0WW6fHvD1cm0XIuPKH61/QXSyvg2Ybe
uaQheqQIgIYNNF6Xmife7esoYJD5pMiEjdgb4iMtfat3UFlSXKQx/ywqzwZE
2y9G3I+zBaIqHEYhX6WKpaEvSnlm4un0HsO4ex4cQPBacJLz7FjLFDiUNFRR
yKGAfqW87+JHuH69PymgrxKx/Tw7+xA9CFLZGPivtP4wj3mfWM8FAU5Xi4CR
VXo0EeGdaoKFFuBPOcy4+IwkRaiaUuVMPK/r1v3L+wvmverwM2FH49b35wLj
wGTx0f4nvgrourcJLqLwFCCZ54QN+AUOrPdZJ/MqSjFTxJ7+q/n5Lve+/3sB
u6eFp+zrxujj8gcPAiCqM18fbNLffIGBSItXhnyMcEWUx3tRxUPXmDLs0g6j
1xTtAghLu/gthP/0akc1x3EB3K7qBeIAH0EcJRJhTGCA/FLwl2KWP02coEyZ
IiQGRgc6OrimgxCqFR8WhEaCXzA264WcTlzpO8FcBstKMdLfWhfDRvowT2TW
310z9BC/by2uo4qvbfzndl36LmTTQKC1EYki8iTD/esSWcWReZAo8x0OONJw
K2M0rkgUNSKQvepLG4SKB0/VStkIYfPMzaTSkhR37DZ4nfZ70r2h8xCr9oVD
MeP82TdLYXCH7rIl8NlnKuCz2XTy2W58Dq5wb862/yykkpNdjhFVLj6T3dYk
aUB3Di9H+WdMp2BO3kziRkwUSJukoSUpw/fTCN5YkNJ4TM04G0elrm1yC8Ca
hqgmk/ar3QhUiXM5idnYQJeHFqBII4eArVTpcLGR/BA9wVowWRyz+om+wSwC
ydgnBdBayTk7EvcpTpsyDk7HYGFDscUGlymJ/Y+jD8ZALnfWeqThRk2t94kD
HSgRvBy/6mhOSOMv7m4vH78YgiSJ55kY2u+bXmtIYbcZxs/WEUKiIc7yJg1w
UFAX5kBoM83Idbh51kqpoILImjYDKoPoIxdTrnSigZMmEffIudOPrDmSRX25
g5qTbKY+IEXQDGOdi1rBz8bAVEiO7tbeU8A1THoum/6D+/l4HaiVGK854rLJ
edSnZbYLlfcUOmC0GZkZ9mb6ViescIIWumG4Zplm0pwNTtZhh24wnVqNyGtq
6aV85l2ZRS3ERNc1aiIrjuyel1Th2e7qfHliFcyv+P+20cf+QcPMkTOp7gZN
xCoRYwdL2ffxh8IFgXZYJKkrCzJOc8OC8wbf28mKoBWUPfae0D4VNUqlUcd/
qBUPO8RKDkLYqjI0axlGIzjUReQhufN218CLsXdIWew8g2eMnH4pTN5zK7UI
qbtXcrhsp2c2wLmL8OTQLth58e/Iqwhp1kfNQ1RnCfOf1atFjK9nR+ubrppI
YXjdR3xpxIkK7vvILpU5YtQdTu7+V7NzdVptHXv5XcIvECDX1dJFh6htxQJv
YPceKjIxr3lad1srXpkbfq86SKvBOhEyhY9w8PxiKdL2gQU8N42jL3NZUKHF
+Bv3WmGT3rCONI9LFDg9mejCOKkBs1MBm5Ssn0rHc3Tc8B09iO75ypJywEh2
bW/w7x5GF+5bpniudycs82oy2JYw52TBMJhlwshV0ivYushedq5deDmWf++i
yZeO/qDHsAVbl3HMnnzjcLJJN4l7hejXPR67SXsvH70XpidlodGxGlF7PKv8
7zc9lZR+UsMamq1UAXAzcNCotL2jd6SZO+ajBny4fKIrG5c/3QqubEZPy3zX
I8g7jmx9jVhfgZubIVwOsXF01pt48VWwqXbB4mFedck88da4a+luNTvw74L1
X8qYccp2Ne+iq2LwUwlo49Ztm5koHrV35wILtvv2/rEz0ts56tZ7+cK7dewO
NHAmQjokQxWeuW7YK9RN62E+A+enfayFunJugMV4HFNpss4yYWAX1q+GXuVx
vKyck2els5s50TpMoSJW7fGXe3dkpysk8BqZkpgwOiQcjUyaY/7zW/lRcaBt
zyzkxFqfTG/FQ33UIkbHOef3Fv1KPKxMYFAE/Mpkf6wv5k95llTjWnZ3adt+
G5SrEOl/iUxqJoxlZBzQ2y4mH1sZPlI4HYBd7051oqSbXj8I5LW3E8B9jvLq
5b9sz68+KzuzOiw9sjxMjIE4BOLomdwbiZXhe7RB/OCm4UcCbn8nkzpYUrvK
ylQ/5EPDhOaozYZ/NYL1fh82yLqy7ga2RAgf1XN+gAJpgeU9SzeYYWURwwIP
VKi1zUMNKJJULWlWy9FJkxbwf15AU1YsebcS9Nv5dLCRjKcq4wRieAOKcC8N
LWAOhZxSHY2bWAhrkdY3bLbxxKPoWopcajxYzCDyS4nKx6D9YLi+dAkqB4ul
ZfgdS2uEoJeM7YBFvXC5NWI6sdeNxoCnBkHrNGnlZ4jW8KTgCEI4RZczUkq1
YiiE178sUXksBbAXLUW1ueuRgA8MnT6aRUzIfVM4y5dLiO7w1D71NNc1QvZX
yTz4gTkfR6qRed7eAu/sLFfHJsHMLDwj8GJaBa48RyJg7VJYRueFUwwpOjHg
WkBIJCsn9JrCwa1V4ugTgu7F4Xk+0t2EvVarqo//+fIDyeIo3b0cYzxTVAA9
odhVckC/9S3ggc+zQZzZe8SB1Of3p+QqCT9OPX5F/ondLvU7vqOvZUxZc+lY
kHkyJmvXLvLN2ssD6TjQlTUX5Jh95Ltmn7ij4Jjn+pt/QjziJ3EABB/Pwyji
DP3NxAtPPYwQonW2AVighsS8u8c3ewAmGdbJ5TM42It27aPmj/WiucOBxcnA
x2cqj6yczo/5MgKxNEoNTCWBhUNWBX5LY3usR9HDbMxOnsvIvoW24fJOzyCj
HTiI1/oSd47qZ881xypd8xhUuXhHLYKQW+P9disE5UmLcMg1flBrt25ZYPQy
H4Qi9XbPYqgyysniwIt55Oyd2NMf8d9Jq8e6A2/4OCsjWTzRZxDTD/ha2ShU
BvlKqnLCvAnAKaIgULnVBqNb7T2As6icSL4Iin9bqtFabasZmjFVjz47TOYu
/HZdhXpdmJAweg31OIDvLWgFd/4tF+pL0CIteDBbfiFBs4sngqGnE3itRZSE
BHddwBRbNp27mWa34lhp8GLNITH71Um/4/0XdazJnNcwTx8IUmYVTZyuNjNN
owHkPsQjb8Vd8WOqxTEMSm1VFk5zSwBzghzrarZnotOhAJeRpSLQFXh1LfQs
NMUQ0Dghszpu6VhuwGVLq5c5BKpWhKGO6GBtMRQkAfederpsln3eSOTMV62g
hfcE7w+Jy/iAsFb2JGawSew5d6TeJjkYw0IpJ/9tTUL7hA3/g6/JlAVqQSFW
fGU9Hv8SHTqcHtVbdbTrNyL9DuFs1o7qtFBxVVxuW/l1dpB7euesGcSISZ8r
KejupWY3b8X6fnwKOkmDhJdC2cjpb48xyWgAVeweVt5m+DqlDIojQop21fcV
o94lYU2tOGbjEeBNATUMoyUzEsOGY6/mDJ+beH1WMSxKmB2Tv9gts8DkG9/B
LXVZxssGF6xJSDDKfEWQelAVQgpNl2Wi5ApHq6AVjQPG/zZ+lU1UuAEJ0+Ga
AGOlNAAuZZ4z80gKYx5HfsGfqOXUdYHBBTjnWGBxf0km61GH38aT6pWubdAs
Pmp8u0RW2+ARUeCxs9+UmYa8aYe3

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeiY/kN8ErHSwkdG8XAuxGhAAksWR5h7pUmqvU/QrbirhDJg+2X0WNhTntt243yzSkz3L/yJeMFn3/9QKZBsd1/eoDRie0umjmog6vyn75TSRgMgkvMbvPmWVhui+EYv1rHpQxUpNtqMIUHmwAogfeg/mNhETyLmacr/uqVoUL1rRY6mqpHNmf7lx6194lJ7qWOwCg11srwfRvBfv8O0y9l8BVspmo+XQRuA9cLtYO1ouea6oFXf8RV5t+AkC3FJZdKJnb9XTGRksVF614JNSj1rLbl2qi0FQtoi1VV9WDbqEmNVvRImeGow8e/h2Nvgms07KuWK9kVyLGC9AzUzA1FYhsSLZzjyg+QV5cyj/QV1ANjZQnsmuduAcgDSSWvlzQ4FO8KLzwOB0jzlkspDmuwaop0JDtpW7PHUp9uYh1E3X6sPhSwU7CRUdlSPcpawH5adtGn/041WtLsComQtK9Lt8vsBgidNPowDxOrxz53AaESZIRhsLAn/sIfQAXgaUakXF7QNxLlDKpBBpzOLUyL1XVb4/blBqFm3mVTwNvrTO5V7RGV1g37OvAMlmSobRRh3w0ldFLxb/IJj09HQ05lfMVS4xd8MGAl203Sm3itlQ2w58wHodQZW1lS2aL29fQl/d+TMjzkUXUVlapMZC0s67vzHY7ULtImrg37uurAE239o0D4IDZdVvCVjfqK4/qEiXpT83SBXpSh2kIWlDh5EPoyYsdeJZb2bIdoyVb0tP7TgYXn8iRmSb3cFLhapUnP+k+S7R8UzyjVfn4en0nAv"
`endif