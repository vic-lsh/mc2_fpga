// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CWIDq7qMeVRXx/VrFQqqy9Bq2AC1ZZQyYym+TJYbVUNyAHAp4g5Bu4eq6HV5
oIyjf+GhLepc7aawccMt10mtRWWKb1adGMLlE04YZU9z3BgkhZfMQH7U4SAv
e/iC7yTjVnokc67xnerNNo8aCMDzhzjIKNVAtzXKptP6N9RPgGg8Y9UKJbaH
EnGAwjfi9aKgiiBisw3DjQbPkLKxnGEPWfzIYoVIS5ptOddaw8mG5uLobMNj
j4yshvuyjYrblYUEOE7OdRSDYdc6h4ITAEDwS6/RRsDp0JummVDBACk2HxPX
STnG6BfDoLWUTjZcRS3YWRn2CZQOTXwuhD3ECKAZ5g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Nmb75MbtpeZDKbvY6bWkpACvfVwd9JlpNy08D4Oq5x14CfUl3nHWxAmeCyO5
rVXXuW2A4ZsspegOgdV2d9OCFM/vT2+ZBbnb5f8sz2JptrjEgkx1Hoqd7EvS
lsdzajexp4e9NvYLMeEV/HqDmqr5F2tk/BFUOsagkd7xjbmMUyw1r9RUVoHk
92iQJJuk9KrTNrlwA/b+rIrkr5+H1J/leZQutC0BHtpUKWTuKjs9RnB4pQjh
+SfaalS3gGdpEth/AmFzxGe0vJklBn8UxIiILh9rr/z7geaxU5NWltq7B+GJ
dsDPB++GxZ3b1TwmNoec4FdH9QlWP/cqoXeCyyU+VA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CndQkiSLMZ1J2RIVssgoyvaB4Ejm5+QSRs1RhxrQ85XOLjvmV2oaGrfyRe8O
23kgJzLsCCYOKBRZj2HGiTdwL2wQ/F6qtO0PMmibzOvTB8A2EAaU3HAwBGcf
RvYeg0H4URnf+KIWvT6aSx/i+87EFX24hCxWqXEIvwbPLodIwj5ErFQZzKz0
Xm57misGrR2MMw+nKalcOdgo0qWLCn9daxoApgEC1xfnXTdrO0JM08U6goxs
Rt9MW/BvCkVwSS8TTKy4cuMM9cvp2/kH0CmmhaYhR8mgUrBJAdYmLuVlA35k
WygNttnu47e8OOZwrcMVb3xn63RbtC2+0VkfvkYiFQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mbihi4E/igmpVdyqBtb6Zzkw1PbFbH+J5tkZCP8tIc2jF6xzw85FwUlrJteN
vm4qmRvh54NIr0NeiKtJC6m6hhFgrUxvDZFENhsYMawcJUlWI02HUonWVM38
44Ww9ysEJg7b2B6Ib82M+2dk6uz5D3casbROsqgdX7ku0T0vIPYDhiI2s6GS
MSkQnWCHc1SfU/rboqkIXL2RBbApSOxm4oD90YLn+msdxirOEI8EluhIwQB/
XrQ5RYMbXCtVPmSBNNKnTIoqd/JByvKDhjAj2/2oNTwaSLDCUNCvD5Vv0Y17
oK3hlX3T6vWngsQL4dxhl2clTaqIWzVjr27IQeGk6Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZcQ2Dd7Kc5g3aQI54iDjiBeTis7K+MlTL2Hz/psSRf/lhF1I7AeOiGgQBZFR
/+AYtB9NpTbXsclU7pz82DwlN+RVMbxdyC28SIhXjomrN6k/G6MuvXwvzWkd
ETyIRIEtQ2TIFS1n1Nt0ac7fibpN1jdmkbxINGYQVY7p57KR6u4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
STjsm7fN3uAiGfLr26p0ETrgj0VVBv2rTtRB2x7gki+hxFukox13DtA+Y/C9
8JLB+RBTEmjvupF84Ic1nOgA44b8ioqBhLNo+n6JkWnfDjsHzDKkxhN20UTP
sjbI2YYLcOu/RTQ0DUMLN29QuJDXT6bnnU86Fg8l31bMETkF2dNUs0kl5MTj
GNq9+3zs135dH8s0v+01Ht5ac7MfTLXafBvQKFP7m7zvhYhwDGmzLO4ut7k1
U1TEZfucETz3xAlyqW10B4UNMxQGhmkpa1eBwZG+EGPbymER8/9u9NQZXCH/
VSiXS6zoyAXexW/nk158Hmo9FUKxmp4JNvsakZ18u2iw5bQW8+7qo7QrGhfk
Jv2crc7G7HwfMfN562WSQX08HlVPKoGxM+SQvHsO112bsIhAsgcECr76sVh/
TKoPpyHPZZO/c20F/NSgh6groMnT27OMzjT136BTpqjlbL/RogGzZ5qZbEBf
saniQXy8OAi+d7DbcqOEMx3aZRcJqbLF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DohIPc4bFDliC05hJOGoH7/S9qD6Us9PjsTGSpPdzmtEGkXPMMUB4uX6Yw4l
UW0XsE70NUBsCxRh0DR5VYyZblWyOqz8r3jrWdbaC50aEZ77wxlBzIq2n4WD
CgeUG67hRmI/nLAGDxRHvhEnQL81eD0mGzKLlJ5CSuOEEcqMX7c=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dgO1oYwmAeZ1/OWoz4mAcQ4zoamz7x70n8DUWuVv4vpayo1DOY6MYJQ1/uH4
u/rbHgBrvcU24XVGSZgJVry2SSRylSwFtn9LzCVCiafqzCRs7mrGWiuaKJc7
gTbRaF9eHkOp8ptdSj5WFh73bw+1LAgBiCEYVdnuXyDk9HUUBg8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8656)
`pragma protect data_block
jKLephGVKDwB49dJIJgvFV12xsJAFY5RUEBCyZUWLtS8m0GNOqoNpQKudi5B
xitPvk0okSyr6TGuwH9lgU94ZzjDSM6cnPwDsdyd3hc/C+TzDl5vGnlE1DHc
T9Gsd9NfpViW5ee38JX3f+oaYpXCR16C2v5QolIjKrTLl7sbDvUi29G8klUW
yIlV7JILrt0QIdxl+B3rI1HMXqHryPRMq8hgMJHxL/y62e0O0tjxYgkeo20a
aN2nkeVfViA03Be+6WitsmTK3Icwl1F1O+kzlztBaTgWUvIQ3E4thTE6OlDu
sTW8FqfcRFMJcPPuM7LUrrD+7JhtfL8QJ5n+SXfixBTuHKIHWhdKXyb5CEhn
qdcz0KWCJzm0Z9B/NdkS4hC8hnCG9NIU0F0utN5UjmbF9TZ3IOpRYOwJClu0
5LFpJTW0Tgty03GI9vOSM7oxwKDFMeI14DkCmD5Y+QMzwFB7ekPn8KK/mXZY
KV/j33SrxtyOTMXc9FJwumFchdNjH4IXolZdTuGmfgwEgQazfY7zquYAlRIk
u0ueik9aaxuWq35nWjSieEhQFsKLiz2wWMoWbmAvvD51E7vBrwO6lr2ZUyL7
OJ9AJ12Rt6lPnwJN76+TCaUhJLOyPDqEA9WFum1ryrIFw0y2YVqu7hWfgASU
JPOJAzdQDcZAD4fZlQcYUz3J+wU8PVPiNN0KgsKYP0UbcgCTfruFersZ64Sh
niFzZbq+rcVNIIs0D8sHS6wPVgSRnGIRja8fq+M20Nas3hmeGvoxu2A5GV11
7mN84b0JCTzj4sXH+Pw1SNX7CephvUnp9OhJJ4w8+1TY9FyR8EvrOT5L3tyJ
9KsKj/D32/cw2wI2TcLR7GREczmmta0x8bT3id1svTpjHtWxP0d60f+Z2ww1
oRn9Z/DakeLfrsBkpvRDR1+ekdf4QrvhVgmyn0uV8sS+JXwy1UQvjAb/y+0d
dkj9V0jPIz88YjrXVeZz/0vaNgJBdafbNv6gpQlZkbuawPyUDWZ/9ffND2dp
8wXsMl4PQ5PID8kQdpHX74MtiIighmcCz2SFZCsmcgBNX2PwY3TT2bLugKUD
Qg2yxii1mgP+9VmaKGGFWAwSRJmAF18dRNZpYDWiXHknoWhyLKqyof41D2ct
PpLDJtyaDRg6Lxx6H9cOQCuu7g33Fco/TQ/o7P0x9eSR4d6yrQHMb1FF3CQJ
HAM2kChIjBJhT7xZGXGyz3Y7URWDSEbFW0TErJ/gqCuibnqwPNTEsKpXEbWN
udlkVhEdadD6JkAOJGRFqUzmbnZP/7I9bvEUARR8DmPlIy1jsjIP0SXWwUGy
vjPzA1zCOTPFSW1Rj9sU7kaCqwke4vhFRoEpyj4QST8i0UeU/I1qMowLn2hr
swqxIQqsWod5YadwZgEgdCK3tcB8SGwB4bkSTSiuWOH5jSDM5/6sBqzf527Q
phS3bFZMyq1cY7EDNJK1zcwBQ7Zplh2/rgVZYfN/XiROdhxIo97FwXLNjFjU
GqV4IiAyW3VkgCrCn0RYsDnR13sQpL2Hdrw0vM1Ynz9xlRIT46n5ljXQeY3y
YYeSy7ghhD2Twf7p7h9zzcbkbsjw/t408sGOMjX/BEXjk8wiINFa9idGIKs0
kqZUmzVLhAHx9JFaKPr5OckfT6/ak39dgzlt8JYdL8ND1eyE7D3l7PW85aaz
rdcpsZZKaTTjIzQu+n5QYwqmA2geuwu+nIBneMPoMmz7ef8OcmRlex1SuO65
F3ptg1PqXUJVkD8DQsqlXvVNEHle6Y+AScj30htIp6mpqUg0tPDbqx2+WmwN
XCd2qxpf8itDdSDg1BbH8AZN+BVY1551ppdeU1fkLBOyt0PKBPbukecMLSFA
hAjFeu1WLDguZY0AQ+wFEeO5IOhSYqDZBGtue79N7sRFpv869x743djTNkc0
3orMaHfcoZE2ufKRtXJvT1IZD4AsP463J+nieREnfZgxZAoC+0evkb1ZwUnl
OX5uzdA6ZtPm8BtacNUJnVusRw6catN1PurGsACxlRZXPGdM5aDo+UDARRYp
sCm+SXSEkKrz5sMeZnrFDdojcQUVboyou41jkMQ3ifDAlg3ZejvivT31214+
mNwZvLEcXG1mTIBD2AV2+/6Kx6pI8YJQK02wM7U3QzfrBNTFIMF3z1DV7Da9
Pl3tHEEUUP3ft2LEqzo4lH1HXmKh8/bOSiHGNEkKPJRmS/iUT2igL3MeTa9C
CiH4aUuo0w14Ovb0DhnrOsNgN8Lu8FHgoQQNZSUeQzxCZ9pin4WK5MXa6BTf
55/TCYA0EoFaJEkJZdQfUD/hF1vWgxLQjWZspMZoPMfybRJVkHNrRdvvHH/P
TXnZU0usEQlHqHQc84GJmlm1Q8gTwpLFIbBYk0Bw3TdZalUYeVEArhYXvygR
JLxfd1leDBRJezAZAk0n+3pWUJlENaFJn2dn4dOsClbBVh9wbSdGOKpkfwxA
sc2UHKmccWbxmfFnjMXQQRkTo/gP27GFDF4j7ysmAXLE20GUS+cdiv8EQciN
We0IdAW7PQznGpZ+BtmF/mBnh4m5NnrRX9lMyoCk7u+FPXJS2aIfkjgjgVsU
SQoXB3pyhVogdmdVpdrVtLExDTeIHkCzBUahyuxw+7dM2DZOSg9AEWTd0M1S
Y3E4pa9ZZ2JSIyYgmVswhp43bsYqE26P7sCubue7LP5/8Q3bES93GbNxtu6U
7geOu5Xd8X3umAwvhX3DZ2nbvsQMSN8NfTNGSOlj0k/4nsqDS1fsF5MyAREm
2R2BghPRaIebuKGJ5xY7KGGd6GfZSyPRKa+/jvvPj47vB9nmpfWJgwd1DfmY
4cFoY9+oal+rJ4DW3c8FYuEk6D4tHcFfbl2ej76FBtoZMqFzkSbiNBz588Zz
Fx8ybIbHu7dJ12z2inXBXDrrvBJImRT5F+W22Hgf0kzfg64U5OjAuSLtfHUR
LRz9q9rwBg8XhkdCJi4IlzAeXYQ9oeBhjuEKvUeRh2SbxvM09sK3wwK80AWc
EUByn0FqIkqmI0+mFLLEcke/tjO1AbuuJ/2n43+Md4zw7cM7s9anJ+/6+TVO
dKYKUrgSIQJyU5ID1TLGs6/6qQuj67B6OZFdbPgSdtcINM0KDgbTdm2R3Kqy
OL5f5cTgiSCv5waDdYpz0Fwnt9I9N7H8FgH010yO4QFDQrN0dTQ7lJQ48NiY
v5zmvIjpuezXa649TdZ78TCARENpJA2Fe7zOlYXP78jV2j7o4sVfRwz9KvR3
5zah0J1XA2SkVpyqoi/ByRX9EOvf41swuWScBOyYKKd8Hf+YpE6B5Vynml1a
tSuIFiMHOxBe7sLZCnDVWtpWNfmfu3F4AAzmPibVU9vG03YnEfCx7m98BO6Q
n/uO3wYz45XlyZwvF4U+fqttRrn3qmtKSpXqoeydgTE7i1LzY/gys+pAQGiP
e+o453ltnHhjF+n81DcKbRdPY4wTaplfqHyH91hViZ8GRxS1gI+joqL/jG48
CCuvKdL/NleY9r8lxmvE09jmY2bKhrstbkTGcYau327OeVCrA7S8j/9abeIA
YfyaPSsoMcTRx8ZE5urB6bz3yTbyUgAoL5EGlWkg3XQd5Bni0QIsfyD0WIRA
BcgbDkO0sN2+dQrKXq7zwoQabhTCgB0UsaE8HPmS5xZcmblyBKg1zQpeyTDI
FU3wh92Px8nVO/a6PgjAXqDJbx2Il5tdlw7aPy1c3AAoCbuzxO09EaLz+RaX
ffRdXqBKftZCj49kC31d+VLXtBHQsfSXN8U9/QwC71Aa71Wimzpi7bCOYxUS
VOHclAel7YHXlTaqozcDf+cA6l9jcU3TmZ1JXiqjwd0YkgNcQxQ+7d9qntP5
W9kgAR9nkNszvaSHlTarHzVQmTxNuk8eyZGYxcypFGHnkjV657d4MH607hIB
MWbVaXHnomn4yFPA3DdV76pNNAI8LYjwWblIUpAUQ4EoPWR9L8Uttuva4rk7
rsAkZaTgyq5kvJqvwhosJAHBrEed5c5wtLki7bncMoa8Ka4i2pvlJayqVRf/
ybJy7Z7B/WC7iKsRclS7R7u4F7fc1q7wImCphXg0yXmdAPg9epSP6ypAZflk
U91nVOSB+dZSTHxCayODusIKBHE9PpVOlGgQMMc3UIiF0lwnOeEXz7zrMSVp
8dmmGUGWoE4wDf22qzRwrMeleRaFSy1AnjnTx56ITvd9Qf8LXDDUlPVxaV6s
aoLvl1/a0N+tRMuw8XtYWiJ4swFLnmA5fdLSKWpjjC1lp6BQNhvxbvavZJzX
bsUQxABsfKrSD8weUfKnF3m6TY3nMjZeUbedqu2pq3+erRb0FnNEL3NNqvqy
+zxzNVcoqJF7+oGKLjcQkY2sLpmRIy2zzUJYnicmGL7YV4WNBUU7bDaRmgv+
ZmHVWcBdz9CWgEa0aZ5hdsGGJX2vTm2G2999vFFj/POFJGCN88srf21pz3NC
DhgJPfriNmob11VT1AdRf5+L5yowM4O6SEJw57A8YV54GU/EyBGpWC1G1Kq3
HD/tjZtQqDVQz0PZwFqbqTEosBoHHXE9FQhvJqBBSYkJIdAYE+J9IEOyfsgG
XHvaCzg0aRU3dY8BsaPxwzEJgdhCu/H0cAmpqaYH87gUVJZL60mEPw6h0jhj
puUbEvi9dDEOEwg8qGO8hUxDz14BzS8lbHkox8e2tyVkJR/yNikRPfsVmHOe
lFSBobBWJ2qxovJmoiLrx2GooXZXBAYK3wRMymyOBM+EfO7K8Jy5Yb5vTzKJ
JVZ2ZPW54d4+ALpPNZhT6FsAEBcWMFU5/F0ZAdgrrRQzjHZdrvgIUYq6uu91
u+CO+TFh1R63f5NVoMpoAQbsvTiVGeGMPzwWqv8Mmo73n53Al90/SEqrPpjd
qjAUDb98EQz2AhJbzQuUDNLEcBrd0IFi1YnnPctneRHDum7wCrNIApcxRhg1
4qwXrc9VWXQAtFb6ZC6uuXmNiPjMhyuZgNvaR3kIqg0vH7lCGH0EaQ68imiE
5LB8+56pvLJ9DSF4iPixs1VN9dKHXlwj95mGHtuLQVohkY13hqz4hODBRXvD
Z7cws68kC76+EMnD0/dwMkmbqIRLcvZfgRGUWau2aX8NC7M7J4ZarceCc6GO
AimA7DPiIwmDBLl5znQr+A5Ftz+aRlpXkRXw0LE+FUFgHqcrHxe+nKghD5Td
mAzRDR9wefzoxihr8bhCURSplwn0ozBqZaUcjsurDx5OV5ubOJktD8AF3iqq
9Lfkg8Sb1RGwL+lSgHkNMHv1zBSZhCY2L1afYTh+WXIiqqvA6uhMk+kTzMDd
dyoywwuKWx6oxgUlfDW54/fJkfkcewyZvDOWYg0+bEEgYfhxIIUJYgMULZ86
1P9c+iAZt+At+nVzEn7nLFDNgse23ZS/Dv0BYYrfGD4TyyOb6ncxzs+Sky2c
OZIREX12cAiwwBER17VbqMIE3/2E8XBWrgtJJ5GkAeXEaRodo0Lcp4u4d3eC
4GzFFrB9/q+9cP0AyHfeti1b7qbJyBoL86HIc51r5GZBX6uijznRlJp+z3u/
BlVi4PnpkA+moxyJTNrXrpw0fbK/zgAYyH51EhSXi9NVAJAyigGH287+tCE1
ppaeWpMbVZ0J2zZl3qf8NGvJVhjFT61OxpSPO8gyB9ToIAYLvEumRcfQUvlr
tjdRXyYz9RekybbfHGcTAuYNN5KHNwAdrNQ5LS86t0k3VXO/K8PkHSANST1V
9gvRz/Vz7/mDGXw0/c5Utt5xhUKLBCZNW0TlkDcIGJZGbeqwmoxiUbG+QE60
SkBC3IM30irzGr+Aq4thm7R6qxorUdLVjwi2RSyIeDq1h2otdONuw4sPObG1
BmPi0+Hp1E2Kw86I3C0Y6ydftyVqLQee4BkocFrePITv5XTTyIR9KcZit0Qa
pWtUhjUei4gujZviM3bzbVgZewBWWZmRMntp7RDMxGPkAQU9+9yy6G7a/VTm
WhjoBxD7J/Mu0YBBetvEB0FOnCVCAVzgr+24UiYvLXgBYGbOo753XR6n5z9G
7A06PpMVzUIj4N6ZJfzXMPAF3XdeLOhGcS8MGnuYNUprYRjTw1YBTt2a9FVu
6EDAFMSzmjlreGJgWO+fPfhWyOQ33VcrMf1j2xEZ+9BteXPjZXzoi0HkNKb2
I27J4JfPq92YRUVW7ts1BdsfXGzZ4x8L9mS5f6dlXX1yY10kJx3/5H00K99U
c8b+JTKl/yZifPGw0OzcyMxf+9Vf6IMfKbapGYkvNT+4iQHj4a28ru/oJoPU
WymlxmXtWg7BNTYX4uWQ/LW14E+GcK1y1JbhtFMlzJvE92vaTThg4yQOCbrH
JsCTthiR88PCqu0E2Qf/KbJ8Xbpa+0TlA9A832oNkL9fQ5N/sb76oSFmX66k
YPG5wyxoR1SiJvUlh1yGK69yI2vVDWxUN5NRD5Ugce6p/C4gfLagYz0s+V66
V4AP/0vytVLS+T/QIHqOLvxCIDnJSiFxOx37mCB0dzd0SgPtXB+K3hR54kVt
R0dE5hU4XSWQtIGp0SERUTrYE0UvFb6n0q1+Xcb8TP0dXIzyCUNKpckQ424i
FHy52wlR0JNzy4dqyPUMCD58Tv5U3+QsytTTzA8qpNKSicA29TvlM7PeHMqD
HLhyC9hkt9JmonyBonJF+XKxqy4Yw14MAwHiUZ7G+my2Cd62muT0zbYdRb68
+O3n1q0qZxSQWdMl2qBAwVJiZeCz11SsY1MNUuA2ExQKfc5TAea8HODj1LLg
R2eC/t/J3gXcWkTPZXd2hkGR78nqhel4UrwwkciYsX/l7q1MrWIaUy9dKLVp
fwHDUGQdikeu4ftipJv7nFV5ntGNClynT+6FqcLN9tMoIzkGFp2MGBDvXw/D
X0ojWqzmCqw/0enUf/4RoNg+9wRupBttVEjlh7rirroLOEWq5evlYcQ7uzlL
BfR4JYgLfre+U6gUB9FUbPF/MMZB5bWECVz4YdvTdAcCxV26UvHyvYEkG4r+
rkkLflsi15JfQqcatkADO9NbyCoqzYg1fDdXU71gQWzRItNzyDq2OxOVix7M
1BOBUinIj94TWB8tSKdy9T0hzvvECHMdnttNekDGuFFwHJj+rKv5M59GuTvE
132TTxSNshDDmhNtja7dHDxvmou4t67KV9xDHX1tQr+UqXj68sgzQddKW/CE
utWxjpX0eX+Of8TRQoHNcMWn5NEFKctVV5mY4XUlam5OS+2hah3Nk//jVNpV
6En8FUSdUEReOKbBnsjO130j6XYvg1mg/9PAAhZmTVDAp4hoCFo/ze0GqLiu
ysGO8nBjp3PkBBUfjA6afLGnfjT4UVcpVpyaGrcfRdZ+S27o2SNdvJgj0JH8
noKBAJ9SxlVB0AMMzt0LcZ7PmMSAIeTVKOy6LxrvwgDIiZhWamYEAwrHsNNW
qGOTnF2KWBL9xHKIpJ2EIiny8JtPDaBvYXvVRyvjoqP2glEb4ayuPpH+PZ6B
/sfttZMXDDeu9xI5OixGQUr9C9tH5/RPuUHdDfx7rl2gFI1FgrVequWqa1Vp
KiNdTf3mq3E/MWv7aLAvoKrAWW0Gbn0Wu9TUIlxsGQUSfTxfG7rMuY07hZTm
CVzV5bLrmwAXdzEsABC9gpJIb9F0foFFNybgVybA8+r7a9bT/bOVSgwdVjli
mcwFqZFhVCpokd9itfZsFBxdFBoC4ozVWF4kvEHaU95wOom1sufXDRBcDhpY
FDcl+rmuObLVx/l8uKqVuSt9u2Xm6nv5neZEFoszQDOw8M/9+7yTIAslWSEM
f2YLsVHVHK31rcDp/FuFayiIBnuV2hXj8fPhHGwd2foS+V7URUCQW0kktZiO
JAbMRUrPzl7jHfgPEvIMa9EsJbUFwIbsJxniOIrCvibb4kOeYu6M+W3junDZ
cnMS68dntuC2ZHwLRpG6yVtbNUSQSSDRwXNKFmlBwiKQkViIdoA/5hNeO6s/
fafGo3DCcgRm85NB86//4IHl4mIJMhtk0LwQEfsLPGUpmtOfyfq0UvV3icgO
8rpsAx0r6aFCse0ckAurMrHA8WGQou3b27+lqgJRKbdFpWZfJyNDusnqgixB
xcR/x+Jb+SBeDLWZ4ZZJC1LVpR3pnb9vkjxH+jOA8ugxcaY3W7vLkMqFchyl
cC2S8spUfwu5DPlHq3yMHZVcpYzBHMFMT57KyZIBBo2fd6ib+ffyezbSg+Gj
1E9CXgESexuz5wnn2iJtLqsDGPCZPLZ0Zqx2qCi33f1foYSbelusNMYK/3vr
//osIIwRDN+S2NH+cBtL8kMSUhmgqSPR6LR12TTy7D7rXIclFC7rbSCZl+DH
S4pLUbsHUzsuQTWDGAnWri37L1Np9fRJijtNAFjPd4+DSJh8OdU4jpporf+I
hPVAiz+vYBZlB49UVKzUlH9Soxd48LBx5IPUZdntELtgAEAeuKiVneg+oYb4
R6DUWHOsGupAfzWbZ3syyYrrWxUoASIJ40cgwuhP1aWQ2QwRCxylbW9KBp5/
LVsngNmZ0Z1EvTxtUhvwfrtoNk98dtyxCiRNjRybqdI1uNVQ8orVlUxQCwL4
CFM97yUH3iO25NVapKTCGk0Lksdbgn1xmE85CPenTU/649LytbG5+dH5oa3o
Gm4dtFU3irWi6NmWscmLudNmcGrb6eCF3+L0rXrhn38UqzU+1dxYl9sNRTEE
6UGfBi09Us186+8k6Cob2AyNYfEh6lLvwYkjU8dRe5DhjSRP3XsQaqULXX5f
8nLrSWo7z1tQ8+bJsK6GZr7i7ZuaHQATKhTFlx0Pxq7ZE6w/C45EsLeR/KJK
vupDftGiA+Pnihh+5fE9ynhvjlel2w9+qoVUAgiL6V5Yk9YoT/ApFRmr45Pd
vDsdmxMEXfqKmxt6EfX4MAl6FztKCUpV3Ho5SwzRF2Bbryb2rBlAlQYNymTV
H7RjyEUl2mID5pityn6yBhGwhg1eRB8IpaJ1krjdN2JFct0bJ4iHdcRR0v+O
IIFmnA5ACfX9dYlz8zRjjH5Q7Q/EVRxbhC7CFFu1A+P5Gm1DmOFc6iqOfNM7
zV2dWX0cvcRK6f7qvMrN2l5VZJyKEJ06b8vGbyo1KZH80vXOgt8c+n8tVNI3
TphDFJ5WxwPCIAaci7lhkE3V3/3s+lEmkaciOC43JMKoRafH3AU7vi2Q7YYk
Ggz2EENUH2eJL3WmggImfsgt5J691e7/l3KntR++M/siNq22Q5ltr7AHlbvk
0OruG04SGNhHeV0qbJm9SArZVztQs1rL2FEDIt4LgTdaGPHSXCtBgSgjSuIm
ENZaoZl9atHT/QcJu9agCHSwkvBm5joUp2hPE7o674Tgw2mVzSAZhPuGU4xT
q/kCwDJ6+HM5KGYxpCPxvVS2wghE81NGshTYFiaGR6OprwrvYtsFrWNy5ZUQ
8fct1jp11xKV8HWRQfVWTeT3ITsVFlMitK7cnPjh+f/7pfWlhJtuBkaTaZC6
grKk9fxkkS4oEcVm+zyZcxJUQc3KzGR7MRzelhYUjQCAkOWShKbHRPAM+j5w
VZU4Jcq1RimgxGtQoArq6AkGD44Z6eu4iM+lXVkAXEx2bKtNh3gFQNFQd0Zc
HZVaa01LyhotSVQokSGQTwUTOja/cEKL5RfGdEgodc4Y2VjCxjzrmMlU67Lk
cZsJ6qv1OXduhdWCPRWazbrS/bDfKnPhnjva4cpGviZHBeMsr4tGQKm/hAPA
P3cTj4m6+Xw/ZCg/Em0QfYQV7PkPRzdgEuLcquyBIK87cXC+6dBgK47l8XEd
CsjuHac1B+4tRPWaX22YcR2QakHcq/euy6tlH3xfu1w10SBtfzf6JUdoPo3J
7z8c8kojXH0QXUKShBK74/0BFp/HQt2Nnq1QpnRrzSpOZTqbyRY4Ow0V23M8
9ENng1uiFZHD8eQjebwkHdnBhR4jCyGrcOKEuFP8vIuc5NyeWM1Kj+i0k0Yc
h2xVE30c9wvI3AHShQo4pzk1OPAxek0avRF7o1ANytfoJ2mW9VL1hjmd84wg
QeNH7/DY+v9eyZFcfYyFTazpWpe3nmzbxmLmNue9Skr8rpTvXpOEFrcfhDSU
H8+qJsYnYl7cs7AEussZCnE3rP8w3zl+Gen8kHYBaECWHuU/+6qmR4aYF4cY
olkEm31Amx8+0f8PwLLVOkxgNghXcv3Z5PROmnP4UkN8jYrr0gseczRX9vTX
IH4Wfb4BP1ljl2HQ1eim2jOsqQFEbrHoIyeiI+pD2lOz7ieJdHjy5XPRheft
O4Dar6GTUAqJMYnStoAoeinv3maqV8C8rRPTVLHssjn272Ta6n4+1UQmbZoH
dlRdWtVR/ZwZceSDh1LG0jW7+vSJLmJIWZfgRbMUoyGMRuIHboSrezEaf8So
+MOAd+SRWXC0etBWajFALzAZ6j8FAvHrit/UvAeSeGxcmlh1/V3cdkTvZDC0
hcAgfE+az3US8zKYZl9slPPn8Dl5dnLMHXhxoImsGZ4VittjydhdMbf9fuN+
14oMA4cJj/vmI9a/ugTLQzVAGLsk4LTJrvnogMl/JTq5HX64H0L+SZL/M3Ew
fYozEyD8NNmIFcWCZSkBrlMaEeQlcEVRTm8cavlNIpaFNVwVr6OA++ElO0Ed
ANVikQN+kwlQWNAPkgwEONkKjr7VoSf8Ye97P6Cj7qpxUQRzAE3SCudUlVCV
R1r/1k1Wj0d7ImRd0H01quKmvfCfUt8AjaPW8kiWQvQPPh5EvveeExrXzMKa
+Xx0vxkU9v/+2T+v5KO4FkVqG+USlmJWWQaPNg6Qa2Qgu4JCMstFP4BYmfaI
uLGfeyfZJswda9BTiCkKiEi2+AV0c0cHAPmfSrVIGLN3n8YY9Xww8kQBjUNm
Z8L6VXhdf5pfy48AqezuJVYGovYsU9vW+247Ta+lOY1kh23msy8CFJmbN2Sv
dZW0SnU4jcRlpapyLJCo5/qRlH6SNc9p19bShraReVgtIoP8ciqzkm1bU/YT
iLq8I2vKtS5nPsFV2TEKSRbSqcV3AtDZnR4caSK0+YhJK571x9wAQ+dDqlCB
wfl9Tt5NeNC1cpvzPTS7r1fww+wu3uqIbtezNpsVa4uPxe0JWQCznxXUioT5
OsDDE769VW7DYahJYkC2KlLlhYVdPNh1YGj4+mVTV5uYW68sw0K2sXwb1/yA
+WGqTkNr5lAUONenOrowSXNYAPNDdMODwHccvM/xCAsYWE5f8iftmJdVFvKN
S0nQ/+Q2y5hRIWz5pyXNPxHekQn1UWZmPOpk8pe2u7JkS1Yqhmq5kZe0FKOQ
r+K9/retIy0eieoaW0NnpVEW9ynHWD8LttGmCV/W+nvfK25Rk9Fs26tFw1Xb
fGR6WxwaNVi0pSy6BG/ukWlBw5nfnhuSSyTqdiJjQF2Ys7O8MXoDzOhamt45
FvTZOhP1jy+7A05QiZlUEFpqOnehJs1BXEVoPMc8vNhkGUfH7ZTptKJ0m8kQ
qY/ZRovPl5O+lmZYlohFKl6AQtaEROum2gawcZ/no4famkAZxZzSkbKJmxxV
kY0n4MsO0es+82B2PdZyOob4qxNuWrN0Bohb0/cMdl/LDrFPXuizIpRhvSo1
HEVVyAJmVEyrdq8gWrN0rg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wiTfTW5SpF+psh+h9akvUiXZp9YoEQi0NNLkBdFOAqEdUFSyCPwUWsty3I911yUt7rGRm2/ze7XtX9fdu8cmYu3+XjByLoFgX87lt184AuZJQ0SzNUALsXJJ8o8CCT+CJ0XCVveiNl0v9Bd42uS6DNo7bD/XLtwgACWGXdK95bm/tSeQf0lNKq0PIsIVdLjn707xzytpei3/wmpLD2oPs9RTM+JAgJZZcaYh62H/MkuPtWTUuuCZwPU2TZyChFb1IwGbTx2ksBq/2rmO2PPtLdSPOY7JlIP2J1OeyztalFXUc59WAnMg/vGksiJnZi7PTORkoNnsXFWhLZrcxUo+HSX649ce4DUPXTDIcyJGofRay73MYtNbJ/PVkT0B8nRr2T4TUt8nVjZ+iYwpKYTTbkXFIVPDzH9g5+BO5EYvLIm0QnEfE4fyBozWi5SeSGAZGlUhUyG8UhkASX4uEIxHwAtO/YnqvwQcW2ITOgHRPRAckTBfw9dCCbGv7iuOjwGJZq9V6xi195Aau12SiUazViGq9Mvj+vI0rqYxQhEfcvg/CFCmPjlcojuPQjeLxF6EEIYDYStmcTC3o6tbzdXnRhrnji2fXFr2iP2IeJPGUw0osNSXHOMPK/sJNe3QYylSKNjKSi66er3YwyV1v5mrmTdQdL4ukEm99XCb+6GeC1MJ7/8MahQHMdoDNnc/yc3Hqurg7N9rmqQuvYO+wAduePLNkWvoBHRkmNw5fZmzmLS6hKn6YMuDvfNT6+b6RnkV6WN9+ygRwACNDud/JOMjxMz"
`endif