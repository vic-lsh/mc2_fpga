// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iWYRcaARw6IBGHGZKnJtKvThFKFbNkEsYjqwrdbJBbdh4qUbwjySvneW4dcB
vzITrzVrCVgIP/wBLrwTakALRNX8smF61m67cJ2J5yzfUlSCQiPJmxigkkEy
Q79UcuTrUXsW6ECo400SikjHRO/tT28q8u1Y1leY7XLSpF62qi8MeovCL3mt
rU7uFqmRRrVnQKByiaI8V/NxcIe/pBxUnpXLugAUCAZsGuKpUjHcsUb4IeSc
YqVmsEdglAX7wZ1UhkBjcdDetF0HTZs4siVgXlCg2PPeI6POpTwyWMrI2YwH
c2SMCyatRHudS2n3yCyvlELstUyoynGKmPSx267UmA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g0SJ3Qu/DHDgTMc9zg8308EIAcXddwzp9TJwAZ58X1D5VZcMwqhjFRH065JO
oBQb8b5Pw9Qp6hw0QDOfw3F+bME01E15V3r3DmPWQtxD5XaOM91vBG+OCpsh
MguPtZRnTGbo6JZdYn+XGg2zwgNlB7jAs/6/ClYLRm+13EJdYngt4my29Xmz
1Q+MIXAXigeYEMFVJlhJ3VOzAS4tg7T+mKuIDNSgDS/Kklslh6Bv6UPje8sY
9s+JHLPigvKh/J7Q+0RMMWZZBoqzEB/0jHevAha9hfiVW+W7/9HjOIuYKLPn
8N72VqZPAZbm7596po+rduFEC4T604A0R1GeE8aZnQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G9Mac8oJPIM7GlZnKQp5PqCpaU3YxIWOEU8bWK7Ec7QhNxNbXnoW8js2BGSF
0CirSHwUBsVbhnrHdgTQxU0LvpwKmD3xAQJcBkOYm6Q03Wc5OP3kAvYtAnCy
cj7sUR5VB/VPe7XbhTBs8FulgEm07fF31c6u2HFftyNd3TGGNnvy6TtjsE6i
ASn2RvhgBiXW0n2yjcCrw9FK+hMzxFjD53xPWq1HXOQxsnzvJqvKygzuMQPe
d2YrkLGUgw/XAu5jfLDRsgbgoPDMvemQ5RA3xmPlk06Ms/nbAm6tr+EImx9l
ldb6K+eEJyPbkEYNbNdf62e1zgPljuifMlgiL7VOZQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aJ7wlaHGlctapx8WcBJOHFjLKy8f0ZIweJQWExx11mEskyZPBaBcXctDprWy
javwL7a4EhXsGIy4MPsqaGaBBmH8tplemGDLX+2mi941A3k9sjY7OA/DXqK0
Xt6xRfrUU/Hl/pGPXFGCbBjwR6a/qm6hW2ggznq9KEM3ZDF7av31Mtp9dV1W
BiJzedcpeCdpWT6KCtOYLpLDACocprAX0aipjG3SPSfMRZVMuQZk2PFOBWKM
Ni7/Pj3SnbTFEbrLEqFKW+ZqQ7R6kpAPHFB1jCsJJboax2xmrTMkqr2asG7T
z6nNjLMfK5TzJCGLJG0DycIy5VpCWNgZuuRwzJItRg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J+wOAbse2ctaw2ZNLoLsO0J6Vr0CWlweKCOUZOzKlp42oXrRRwVo66frfDVq
Cmzzp0E6jsjD1QtEoOIA6yed9nxSTn+6/hmfHj2FLzD6HDmC+CbQ0rlLpW4W
rA/OJVAVNSCb4luOXx0F1sr8ZrwP1rr/vhh8YXDRN0hJOXzJOkE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NgILu77U2dASnNZxoEH3VMO0Gb56vPIpgFbl1PVX3qDvkFbEiNzvz2Vwvq3j
nHXS/JI4wEem7Phnvn+4Jj3WygOMJRNROW7uPIincZKWurJ3BOqz0dWcFKY8
jiAzbJoh+a6QZdsBdC2GcsWSF320KKKyrs5oLHMyKXF9/mX6TxHctbkL7Zkw
FVSHSE0+R31HceXR0EgjtlZIaDW0tVimeekeipV6GY2GBTWzMT8ISaMPrhlE
FmGW3IkPFHTeoPWbEsX/siaH4ScQ3rkskw9tcWJqO4VFproMInzJttT4GQ4B
uQkIOBgW/XjxnO5EXNpuuOGW3R4/ImuKSk5/oUq+17CeOlzaam4YoLKeOKTR
fcF6Mnb1TRYU+elLu3tfa3H4qSonXXLIANjCFbGyeZZwl6JFkffn7UuGMHaJ
JW+XawNOkGcWStD6BoUst+HF66wxiabPzBHjJkL2nug7dinjz8cX3jwGUEmZ
cKVgQL6awO88fk1pKsJwnUXLSevzOakm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NNwqdV6lgckPsj5GKa3qTdVs14mi1czOn7n2/xnyh/gbNtIE31iFWfYdPDX+
34tLUmIOtADSEJNVAroe1Xppb3OoOa4/rZ7ImRQ6bvm7mAgt3j2qqGdjkGC1
5dvpbUoK9nT/06x3QYDgeAGtrY1Y7q0OyqERXBeBBe4aSpf1VZA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bcOSdeppntAmeYjXiCUNk8/yu9zflWcnhgQEr+9qv4EZPmdBwI/q/geD4Xcx
DcMvWS4YRjC2YDFCg/ajcnerT/cEqOUXib5uC8796pAMkNoTbME/JLRwx6wQ
bh5fq28qwH7vrkV2OCzO8Gq2nISj35oCaRxNoi17FYhPf/Tmbm4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14544)
`pragma protect data_block
dpyZJkIFFW/8+3E9SSx6wYxhJvOgqCAZ7o+U2nKlnARTsNBq0WLAU7911Kg9
X3ObdreY9Aeg0nPkFl5SB0XlzAgM+Fiorkhkg0qFK8rp9nXWn0H+FE7rX3uk
dkPW8PGQM+2VaIdGm5HjE3quzN45x5nFsFa5GFdC5p2R5oFb4QmtwHEUi39i
GnY7oHrwCLRsczKUa9vOOxFk8aVLRBYaMvVpGn0dw7fJyFs3rNHku1XT8Rp3
f0TBomht3KqVH2S9Zruq9b8HsDv61+7RLuOqLI8S39x4rBQ0gAd3UZrfSAp5
OVzbSrDS4HaPH1woy149CUztu2TLv1PeQcHiN30NMcgpvYD3Izpip3D6stLj
QCvgYZn7yJnmgR/GNFWk97xdVkopOwbEC0FASQZ88F5IULQ1NlVz8G2SzTIV
BrUFLlkuqeqGL25wsrgmlLfrqdD5losIhQSXXHZILLgTGXIWxQlrzlCK4bZQ
nvTmcXcD1z9nFCekina560/cjWesjiVwi+gpWRhNpC3Y+fcWRYPO0/U7CWrt
FqbYUPAHuUwomzs+tK0uuNfpFOLLJlEhiPQ4lP1HfEVnCb609kSgbuWluLxT
ARv5r0DcKvTatzFmLpevHVv14zCbMs4Y+f6YRJiQEg3eNHFFEMCAEwoyXIl6
nq7d4sxw8rzXwDw9eBuxKM9obKbPELtkCjyaEsi/E//vCnxEtMV5c6e8HmK/
dQ84v3feI/HECz5m5qx1nRJ0FwYuqNIBUtGfuA6WndGvdGGTPufG5FLytUiY
4KQ7EcPC26dhsVn5xgNDMMgQ6pwS0xO1FNRdDyay0j09lF8k33Et4/DdXH5f
2f0b4eMVyeE1lrABBonm0ws/rheknf1tESe7fju0SZexYzd2XPFr5vuIFcsZ
oocly9PfJeb7JH6LJXN/uaAxqJPZQbazD/gFo9n9MZH5+fW5wJw0Nr3/XxWm
bcr7eJCxBq5qChuYUeKHTdU1ru9GY9yfvDC8i4QY3g6VCmZ83iAVSBgFvcVP
Gk0HkUFItg6Isp3eUxFV6PYP2lbNhM489Elyi6foYcRZY0o50z0YoKFB/tzV
/lZRVBSgpsh2kTnHeZKmuR4hG/YIfGW0n5tPw7X6JKrEhBb3FulyOzlN9yIl
j5Rw2wlBB0/7UAJC4MNHq6lf+xM+P+Xx6kTFZsG5CRAQgZrxcOitG+5qDpTq
EulPS25laDmpCmkCHK4zcSjYmJ+fZjR9kwFop91vKY5Tg1lQrBChSYeLAWdY
Mir0P26tgl0zso7MDoXrLl4Z9Tx8fL2L8dM0i9lHgZ+Buzw8NT/qBPPRPEYJ
/x2AZDHMZjx/OH46UMgp+pQR8M6zb4zeb17S55ovKLCJte+coKzT95roTMIK
Tc71YgsLRKi3k6vNtdfUjO4POFVopy5Ks94ilPQZjXkF622Nk3x2zHb5hqzI
qYuTJnU9Fo75WAwAd5qoLZmMMoyRF/Z6GovJRwXyisk18ejvCtgxlGpijPbp
W0tRbcbBZPwAoGdHd5PmXOPVgStxzSPbwQWhe9sIYPf3pBsRzrPdnDLZ62zM
tbrhhLatf7XVK1pHFQ7IrTd6mB2YCoDSJW0yq5AAFna3oq0rpssHBy/BDArU
Nka0a6wVnh8CFyl45WHqidFm3ELUHz5MLnHxeYzLtGB6GmbCPKxDXVA71R0P
/aBEwoZFB7zBgdFvIA4zOrYvVn5SiGPDNxkRMInOBOVPdMeLwR8U5AyUQSUs
I9/8G9A4d3qYxgNiQa4xIJSiShzIP/HzQFR75QgpW174Ue2jUQ/fyJ1orY9e
nJg7jUr8lxOb8B2aaanjXzCPpy/io4WtCI04XdFDYF/9Zrou98qQYExM4Qcj
wPwDKXXuhcUOqHvaUqhQO0C9EeR7FdwLx29gHhaaCqMWb8MQSDSFNupuRYRj
rvNF4R1MPo4k/2IKhU6MlBtWqkb8vNxaFb4W9AU16dpZg4T4HHpmYGmVAw62
UZk2nLuHnciyHwsSNCmGqQS6CVU6qYoFbW1TuUz6tObykhdJljo/Anq1uixW
pv1tRDXIqFyVxBDCZVJW1AKrNx0Icm4pRB3panBTO282D9i4172awVLvo1u5
Kf4qlKakCKf+QltyZIP5FSW0C3+8NxOy9x/qIbn1XKoFMIWTYWEjGYC7s+Bg
KoUJg3CQCK5oGsd5u4N+pC3XZrXg1ea3ADEfANMqKExyfUx0UQAX6xPt1zJQ
AQ8Rn58peDEO19WhItAKfQH9sgTucLdzynV5FM0AC+hOoXe/Wn5Ec+9PR0fO
OWzjvPZqWtEnugpfUVWa4kabWw4xuko0CBDQ7fnr8Ey1/ngGZsrKUlAhHK40
GAaN6R1JSVrCw6oIh81eHoPG/pDLwg5DeUFbQMuAvHB23bAsQRsW/Mx5adrI
zvbd2H31/d8ryejyr8UFf/J7pWrbHRLJhBa++jePlF4Dt72SMcezSCxKf3x6
xkSJZW4GkcvljmroO266fV8Po+26qzFyzGQIFOs8byVg13k4/uqa/o42BzTQ
V7peUPhQcZu85jPl7Wjdz20TppP+rL7s3c0JBWtOtWUbg1EwL6fhTknVZdIH
SrCarJpI8y8bC/Y3bR8zBSnwn+0aXOSNwxi4y1w1qJiShog0gmdNJRIyqzNi
YnjRd3DxDlEpNqGTRPqeCN1IWGegaEoScnpyEEqVrFWoTrnO3XcqBxRl42e3
9l6b7o30Cr1Akedpp8goFkFe/u57N6hlo0mrFJ4VWXSXAOJebt9lzzNv09L5
In/BcPRI7VPR+cvxPzRk2XH5xvVNwJga5Of4bXdiRkheR0DBfSizA+0Soh2F
19f3vI7cwAlQKZPWcLZUybQUPDd3gZ4krbr5414yja7MbGlf3eookAlbjCD5
CKaPNgAxuQ2aCaInb2Uv6kMZjPP2oalFi8qE27drxNqOuTy51NeuxHCfLKcX
55eRxjJ2uOUgmlXUx1AqzYf3/YGkLeej713T1GnrTrZGW4nvtxk7pd49Ci7F
Q5CobFpYiwrlL4y2i6N3ES4ug1ASEbMlIUnXqJqLxvbdfLrTp1b+YvM6tqHm
n1p5iV7e8t37NIisgGv9Vmge6e1QXzopuIckfDpyX8Q1eLf/P5TFDDjH1DLa
JH2cr5vS9DDdtjsfMa+4O076xsmdWL+WpXUaxvqQI4FcrrurVtuuJ/fGDJSQ
b0YNRnTUc8Dmp81Mac8iHPnOFJv+C6LW008NzJUq/6JBh83nG8n9jMIbAcA6
s4OlXoZsrT5uGt5+xrQTDIUc92uasU23IcTl7paDAzgbifYXGIm2wbhVeSmh
/tPJ3wU79ATUX7QLIiiTTLEUh4VOutJAtOTl3n7vYJqw53rctBxWnOz82a2l
TZ9t2aVa3K1RwIMBzq/tF1xtDIAx4fmwNjVLrBAsztHwIU01gcK91zarId1I
nhJ/2LprNrH2J0lN/J43a6D6HQT5+qjzfJLsawZ5VwP6uonTV3LbEDyZfBxH
qZurno5+T6wjlGi2NxbFEuYC7gBJysvEH2NMa55BNK7JPGWh+UA7ViPyPjCX
7CwF4tdxt+ayqwiOWk9epkiHcQI/hoOriqIH+3zrl5GpAT52JwyLaKeNetlv
H7PF+gfe8f5iU7CX9LZBaOy6gzRfH+MgWf9BuR7WgjPXSWRjmzOkdFVFi19H
6cQ9iIXmBU3ILbLqWC3+wKN1Lja7QZYTk4cGExf1wXC5uXYJ4cRKGYDpI64E
UEwDsr00/svY/Q34quNBvDWwgNkUaJ1EQIOynXjKpXv+8eLXRXmd+OxbmpMu
5wwK9EohZY0UInmE3C0QePftKBwubxalkSKd154ar5g8pBV6hBm6lQlYM2/9
1HVQmiY54Yyjtovf94n6pMAoQgecZWOHvQvnRS+eRRpRVeU9bju5zH244EhI
lFSmlLTrZ6mZ5ApLo1asiwphuGyYXhuD1nGFjSfRc4rQBWWQ6WuYsr6IG21o
SwMdj/9AEbt0GEc5b3NoA3DA6e666T2aFhTtNlJedYfKz7PqlMoynbDydoEj
q1Pe3WBqRZJam5m9MZVvfhp72aYcvMlMt06FI57FtH39Yhjj19xyOoV3wGa4
q4D9gjxOkGZbcXUEwK9pCS1V6C9KdP+DrscnVDBHjFc8Bs/fjyIJzEMvBbRe
4hipVUbzgsAyTztdgh38VTNymG+7GsgShlgCq7FJaqm7zqV0HVr6afQQwarr
RJOLflBvhtnL/2vD2BaJvnAiopN7hA1Rs9N73WWBTn01NjCKulJcZ+1j439i
A8WjLN7Lnw/3+JkDbOjQYmhHB1hyLpkIyKv9L/+TyAMRSyGCaIHcNy2iusOt
UWzS/iQDCf9K/vVSvD2jAX0YVY28ZpeDqpmtn2Ep19rW3q8HBGIcjfOjU6fo
awfCXrOofhwx1rEGwuPcZmjrpjyFJGk5F8VT14O4aCw1BbMBxAAWwqipv9Td
j8ZohjRXK7vY8Q3tuu/rD80aULYyMsiXwtqNfD57on6JsuGmtu+6zHrLG7FX
Edev8u/TmfD6rA5mZMfFJAE6llnNEIdXv2Xm247w4aR6GCWyXCh/uLHQ3AYc
HF5gcFet+dsqK4iGkofOugKKhFa3yuDRbA2QTZMbe805Sh9ZUriVMF6tbGTe
j3OLBBewpfhARi8VojNDjpBwUAnLPQeIJTfPS9MUCoUW1c1b3lS4iRTythS4
L7Kx6wJfcRQGxHSNQ/nYFEVoji+yfPB6miHdHNNoHOoDtNtabvWsqCs9DYy2
zJr86TABXOAfUWzHfpISYDDD7+SFOjw7rmITLP9KM4L4+uctqlZKFd7c22RL
R5oBknnWJje8arhcjwuh5AFsdXtip/cdeMOtVDYPsfQfNCaMVwAcVRXhyj4L
gJvkBfFaRRLAYw7dUi7ki/DYHi8NxRqTUTKX6smF2zPok9osZE7NeGoiN0FA
lcznJVeZhq7nJxqep1yFhASgDYsGeSv79J7quBWBTEZByeCA4tf6/aJAEvqD
tVF6CqYMbEh0pxYX4X4zAlxv1QzYXmNKVvqGILsto5aMWObocbttk/daHkyx
sXoA+PIsXtD1j9v8cXJs4O5LfrqFYBr2ObFOoHxGH3fafT4idClru3KMSnPp
ocbr0oWKGl64XzsLWvFy1xl9EokGO3nrHHrik7h8VqLbUUDx3Ju9KKppYYIw
+Nm9auXJJk/yhzwhk67Vm/2EAYrvA3tBk8FUa+5K60+qTH3rYAqNqCHLmrbp
/DtAHo33WY/9HG8dffYMX6CJ80L8jU2AoGxYS3GSNRScf/DpPaPDsE9sLxIP
6uwqU2WEt+QVbnQ0E7+zGHG6vOY3UtJqFL5cjH3xdZbM1TH+5nV9ovHcuAoZ
CY5Om/+oijLNO6/Ja06fnn4szUEQerPprN36qLkasyU5fWucBZW+GCnYCshe
JWrwaLhXrDsuCpALegMH/abpc+6LjS1Ee+pXhv7lup53975R1+z4i3XUIvol
yN8+TkoOYwPBjJJK8XrhKEOPm90n+vh761+IQfnzuTFPO01K2egYRPAXUZbj
geH4rdLoCXtkcZIijAWSHpO7N0h9uC/et3VExybC3UHUYwbB+m4Ibg4aObuw
f1rWZA+3IpLksOCq7EfSnNNDHboChvOxWm9R+C5zFXE5JEqISunuw/1EwFSZ
RF5tOJ+RCedIfaXoRNcux7yg6hmKZnmSrzF5IpN9OzdTWsjkHcHH/AQdVHFZ
P+daVanPRAnkH+a4Td0QTLesps0BW8apI1i3W3cFIUxsl2iLI98IVqOHWmLY
HbGFaSFSfCFYBA5QM7tXOQrVTV+2gNm+LrTC97WmPXr1FuGc3GDfCUNAqC5z
1/J9FSKeStX2tyePfjiXAzBo46rrdldsq7BKS+zcKKvNcRHscJnqBWjoZyni
J10H6Rrhs8EpHkAG/3rdaJE4+WiNQISADnk2RPpEXgiW23Ov+FzS1YYidEZL
1ZYGSTw57qcigTP4GFhcmQThkxeNlf87aI8ZH7RcQ//S4gFPNIq0MavvH9oY
jS+cJA2kzGtihtnLWN+Ig7tn1nEn4CczlN7oSpXHsRMcNrFQMe3yC83O8Ziq
WsVDrJmFEWnCqxYxrgPtiE9tObncMs6GYtSCc8Vbl0tWFCTH+aGs6ac63viv
kBoOsYYELESzAcd3HPSww/9nPzbdyNhNXFyb8EVyM9CNn+BRP35K2lYHg5ST
hGu9u/Q0pTjzGez29z9mH7299FzeCPbvQcwfpeMrOlrp38KzuXU+cN7ruj1O
5HC0zbBTEMJXoc3VmeoQepyflOxVHoICs2SGDKxLb1G26kGzs3C/ObBfFJum
fKWvnqNo2UQ30lLAWCKkE8Z886oA4eQgRL2s5YpJ6Pt4Lnl2zMXRHCBmfRPC
m6X7fM/kV0zHDLJ8hkEoz/TwbwWu5XuqsTWcShVexRo2dNgg5vdPE06bftPL
trA1WHSLEWX76Z5pcfL4AyUDe80pCxb82tIpx3vPLxrJUdKjH8J2RKp5P730
W6B6mJ6jtbk8G3S3SupVuS8MqYUyOm1Vy7GCRW/w/X8BFKoLMR9FXXykKQdh
7N8zMOhm/7rv96Vcrc7mZKMjpVCemFL0MnOxMrB1W4d5PCvCsKdAgwbHYa37
y/ZoZo5+YlOVdcuN0zvP0tgUqcemE14z8zscQ5HnoEvYIvjBDSwc8tRk9sBm
/6Uk6octLDw1ahGxgmCoBdWN6eyybG3YqqkNu5ZkEEiG//OH01FH43S9PKPH
6mwbyg45bBZKcpFIbpS0gG19es5AFF4HOGagwRwtKArTriFJg1DtsWIq9mk3
LIRN8kWJrtJOsMXQrNt8UuVFwaxjHUiuFQXhcgwOkr5d6iT6elxIz/b4k7Eg
/WW6pnRqJ8tjiscsLx9mcx1TN7Ugi7K9mSc0/GBIbk2elsZgP139K3hndIxM
emrUlZHz0tiaYQ5QRb06U2/tIgAO+Od8jArX61IsfcP56xKSSSRGw0iAPeYd
uwygcTk1p4ODM3x7G4O7J2Sl5+sH4Cm6mFPr8hexzffWzwIIWLMERyJd2tyz
owtHzJvkHvAlSCmVpb1cf0DfKddpVneR+Wiyi8EtPmzBFOgAQD58ZPvCxmmA
W/nIkcrQp5KcU1Pw8Ye3XhBqF4qFsjFBewWqyfVKEDxh2UFRAcfXI8wSsEVU
09IJqJUdk2oCR4ptLCU6S7nasqUvRpGUBqxcnMb2hIROCVduWb5Tq9NMRUZu
7kVFesathVwvHrSNUq1Q0115z1piHwxFQLR2xeJN62OGV/p6GKA3ekABVt7c
K9FshSCSQYXtICwbgFBtPg43cmE2dKCo0xwdtFIMfQ53x5u1JDDwp91r/4e7
mH5oTdfLffITJ+u6CqHUPDxW2P/ban7HE/tHmKr+O190UL1Z9Wn5j2Mgv1Zh
KwjhiwIEGjoSSADT2632rjBhwCKs8zQhgOPjBBdjBmPARM/k89nOdCA2/4jF
jph5nnFzgVsYqW9vRIpYvhDsGlbSS4XtCpykDhmcYcI+QLvC31H5fmKsGf8+
1bLcy8/UKIAa/6Zc2buHSRE9tNCpW/sTStwVWlJ6yVza/6bt0UhT3ROcefDi
lteRXWkNauahz1WvpzpU+e8V65e7J8Cq8kYvEHRqT4Csl7AaCQnfmTamjmSz
uuI+vQ4TkerH/PGz3HjK7C/aje6OUhZ+iGapOBN4Fvb1mXygSoxSX6GimJId
hkGKjRgr90pSeUdmo6J9Ql3mKym9tE76JZBgEJSd/zWY5bZ4S7EofCMsv4NK
FInF44FSq1lXBBAT+2tQ8l2EX79E+0KCyrGDS6Vct5Auc3vHg6HAjfsfueZo
tlErAm6FA1gsyiyKbCYXsTNIWw1kvvaERh2y3HXMwD91fENVPnGX0Gf0424U
KRKVbC2BcWF3qQPTSkReXge61ZVHmT+FprXHwmXMDdGBtc12lpsWavdZhr7D
41X+QGxY+8drp620iI2H1SYnbS7uHB3iG3dCl91uWOFzio3Xo88IFmS4i0el
cFiq+KbTF5vhM+90Vfk5At6WPxxtcrGOWI+ET5nDrx8enxgrUqQlCnHLajIT
NC1Hd6gIfRkHLOpxxKAes4v65sZPwwpCO/CUZ7U3iG+QwfQ/bZC7+EGaHwql
PNQgP+C2PdW3mTLPBNapf3Ng7TpHjY1zmz2C1ieJhjBtqjr9r3aUFxhCqsKZ
ac80vzS/WBfxbuuNOnDQmTxB48/U3+wef1UmQhnoCvOaD06Neb5keFSW5AHR
/KyVz1TnnjfjxeCnMGtZ79Y8+wmwYmwuMzBfB+aF+eony5JL+/sB9YFViQLZ
VJAposH+Czu69mrkPEW0oT9d/EJbgcQhy6czQWTQzbrNnLzusADUvV2VbKWy
xL9rfWxp/C46FdZcZ5vYViKSpJ3cmYUDcN3W1Ffg0H1/AVBjijOB/kKASoHY
XflKa6cy7NfdiFrusPGlaiv8rH/GvF4PE269x4GJd2PJW2F4Uz+k/LOC7fCy
MrVRg5yKrSr0pszy7BYLbd2UengSvg4VwKQ+DDeRlG14sKp5QAgFSO0h0Pej
FWV+GHKyULAX80DpnYF+4DQszn8bUBuhqzNn0TTVWTEWP36xhXdzA3mxfVWo
+gYLWragFRNWvdvULSCMPSlQYd3btJ+uRxt9YxOtXaCl+0DKpAntQJm7tGPM
0/KCn1ldtbqHNpEdQWTtSsXEOuN+5wXcL/HCBsP9KyfNEPTJytLb6fPx8S+u
YAvKsZse3JUoXvBtn+lIiTl6/Ep4KewZhPeXMZzcO5Wvfco/ms0C/EvqpvLT
dbJYSn9JUlzlDalBWhTeOvXOsnHNob5X6fJ6tUubhIbRZFoRGMozxmXuDIRq
Xo+yxJJlJd4+b+bEB+KEqh+6ductARHDC2WPM/plv2LL4UPKlMgnOsoNFmmC
Wbd8LS11bVCO0ESnjKbm4vbkLzkwqFIMG8YdXU3YKatarUZ/MXVusBb7PsvX
bZ/OlFWF3gIs1C8OJUH4CNklmVxXstaR5m8lXrytpEH9DH8tFrzfJ2Lw1AwY
eUadjtqhuqVwKl3QguVR+s0qxpCESJ2VFssjDjXcta55TkRYc+YHfX0dNZQW
b5HJXota5+sMwxT9K/WEv6IW9vYJbofKhBQjcn4LOJwrLLlnKJWs07F73Cpk
Q5IOmg6m+bgW73BoVo0n3Opo+rbec2hET7OOrGGW+P6vowGBBvMYHR/IyDwg
Loykt83TCvtUP3jWotywFIhvHVBDK5FurjswBaPPH3i2tGZ8m0moyUP99c8m
sYOiG4TZ5u37pixa2NrWSphF1oCKzrmVkGvkVYwoVDiQr9htgLvni+m9iTX0
TGUrO7I/Zqy+DiPXh12JJuAUNzIN+L1eTPrafVQmj2bAdaNi/RUUBeiQK2MX
n9kU3QOHDUcewFmSiV6bXVJlemR+j+xSaD/hAM5bvh+Upzz/PHtPCo+1fAld
5/8V/FIQ5WJPYzUJ/8ltYTTmJY9FKwvQdabwXcnxY3K54c4PRznwXvkoUT/M
zHnfiD6s2qHUx/Q8o/mWaoZeMzh0vQbcB6YndgfamMYtbm8jgutNtWBVf1jN
EH2SxiVdTBkqlAQUSrRdi/b7R0+ZTA4TLcC2Jg1nxS88jXZWL7Sj9SEWBTXc
nWBR2r3dNtfsMGo6Skcir4WBtDoMvUH3pu4OtO2eBb8Fsza0TrVEkApJYfbm
BRZQZZXq4RZrykP7+bIacjtcFvJc3peTr4zITYTnHwL/Qxb9mXX6wnRe/1YZ
bod4TU29DvCgw2N3d/W681bc+qVnfXSBUU5SY5GwlBOwZBDWP82QhhUZ8lqx
J22Fga2ZcjCmwEIiv764AAZoqEWWWqFW0fC7SPoJ1X3qeYBgTUb1VDKDLUNO
g/i3kSz4GKYcUX3pNtbTA+lw+Klal1HRiN+avDVs1lZUt/mhCroVBWXZi1LG
Vr5IbMOj1571M+GbrNdOFU1iya8vsxAsVKtEXgyo98Mzbpk00EQfEovNo2+v
WRUWksmSCX4fIWIrguW+nGBFVSCY80TSDvqRhMRB340u1YcNq+/QzVlHYEyd
H3H55BZlGsGpZtzEpMFs4W01F1u4/4+W/rg5Kd3sSPGCu3pzI+IpBpiN15tN
RXcqrzK2QQkh22YeazL+26urJ2uPBYfTeynELd+ijlr0QgkWpHDz5lrln16n
4XLDARenBOgesIl+cXiWobL1HSl3pNJejuuVzXCMFtsY4jLI7uIU4gg0oYNa
dDX2fLhW6THRO5X0/ZfceHKW8YVZ03ElH3M8BPSFuDGE0EO62X5Bk3Yp5+uD
L5dm9KUIu2MGRReKYzyJa017BNu4DPcPO7kdT8xnXXOfXQqBrJQte57A7J47
2Jko4QswTE3h7wNq2qF1imZikTNFUYnKSiR73PLFKiYnFYi/QfmhLaWi3dkt
hkZEMb299Sx9KC8tcmWsVEE9F0jTvnI7v3l39HOwblC+CHKxVeEciPDuOT2N
fH+Lr40K1tOZER1f0PSWIJFKe/p9CLRCDYA6auJB5+/SbTx9AnL5BEZz4/S6
6I8sCwV5tTQgFA3HAt6Yr+xBunNIrlOS2U9eFOs0k/Xfg2U5dpz+Ef1ZPa5C
PEp4ULzCJz161mP6iHwnsuZaMNf8qhOXrnIZW0GRodEYlqoeHDhJExxKoO7v
cwl3tBRQ3avmZEgmVBh4/yXldT6be5HQ/CPppzNG0/awo/An6NvoKoW+ORik
mYLJ3w2fbOEVqRlt2H7Ulz+VqxNmyaFFiZI3kuyMF/LO7obhDtu/k0OLYsIn
e8nefAsuwhxQ6Giv4eTKnUogksqsZxz1vdpLF+S3GtYSeCqxwqQSjNSpniUC
qmqAIT4Y8w6D14r/kcLPzWxO+BKBbx+bVm5q+KaO/UzjvcaxRdN4uZNAwqp9
Mv/wOyq7MGrKK4bNFBUyHnJptpSMC6+OMZRRBzmtgYSpO0sNbLiiWeOmZKK7
AU0cdfyE+O8gG1RWR7iWEE+Xuur9u0CkcC3MwMsLHUDgJDDL2tt7wKceI0Ez
bCKHx5IsMLUqh+fx3yLxIuR8YG/+SRUAOCuPzTvgjnlgmi89JrxooZJ4iqxj
/C4Ul3EaGY17ihde7mmSUmNIO7tvfsS9vNEejPra6lR0w8bTc8v9jWga2Uhu
q1Lm8ENPAVPi+u72ma+ATqR45O8AoKd8OBJCWISMZvcUd9j1aSs323WKhTin
ST9T8Zzukre8R4L9IcadL/GioYusSqiUGXu3wIb1TLh/ORDaRpvC4ho9eBw/
QY6rzjlk3M54sxlxbMgCkmXJaVbq5NzNwVutgCGk08bOG1B9+Xi8tbukVde4
l3m/qgNf5lsq/AboBJeyPLVCiRc/ss2XME/a/1/Q8MuhTXaYT0ndTf9pvU9j
co1Ahsc9uJ7eoAFPcogHiHrDxa1ZH4mYU5YaDwM6BHAEs2TJxKaeKFHX/rtx
6g5NDfrMo4JeRbXHWw4vYixAyLNJ4Waw4zhRZcLGSjOiAB2l5u7W9FDVHKNb
L7iWi9W8fugT9/XfyTOaJDM/zxra5nbx1W25kzj4Wa7OZ5pKMJMYqSgBKsdu
5K+QKOMZ7s6JEovUESqnyDI2iYZWQ4lH/FxFQ3/sLwBQ3pxJc1wBJUR9NcJg
dEtl8YBMO4Fc8IEcPIr0Dl3GqtoyJaxasSSEnalf8UBcbtaGYmU6VMRiq9KC
lh0I/3SAHeSJfP4xbs2YEcwUjlaDsvErHQobahB0EZKNVcWRSk2UBJnaKRPM
CLo2aCqurl2Gfwv9d0VboEAkYpZAluawJWFijiEEblaFsnIeJOGvSN6sB+8a
wBLAzrv6XQ+q06HmTgSUFEiMx48L4J7An4e5RgIW7g0TAYOc1vx16Wo3Bagf
Pl4AM/DENc9ugoiY50A+59OWO3Z6EP6fg0HcJFp02pZRRpqSsV7jCnfrNzyI
YbgYkjoWeHqizqObR+1qZgAjxNV1AUvzSjBWFnmA+XNhm9OmyDZ/PuMgKfvB
06hL6Pc1Z/kUpbXUKpg7C8G8TMegrIyIaGJG5lBU0VSl90oJNhyPc3NJaPvo
5N5jJpBNn9mESm3tLzu9MqCOWvOusFlGPfGgpIMnDrzs7gDpWiKBPOyQXXau
BLl4/xKDv+5JnXP9nWyEmCCAzkUUhOtKh8no/28GY5PGC1bMtWny642zxqzU
USZ9aNZVouWm8KxegSsWGJfM/oo8RwuDJJfxJKYvX+glhqT0gnq5uwOSFvRB
hkPcjk8G/PxG0NYuXwFB/X/nHCS8m3Stl1Zv5G09C9DXMVCqc9vE6I5u7m44
eMrNMxg9nrJYB0agHld4YfwxjvBBvQwmanCFfUR56F8oYxEYwKBBHeqZbly8
q1IN6oV5SaY9sUSiGes86FsS30UhwQKRayR10UqWfl9b8pNXkRYnzCV9HzXQ
JeXR4mHpRLsguq0jUYIBKt4FyTPa/zfp/XZoOarjSl4Gh+iIDFeuuhEzXrP4
1qc0HmGbMEmWYrWW2XTx6PDkqVJ9OCGWU+68PvZgJMhyEZhCd2YUdLiSrEN2
4CuIfaFmEOYoWH5GRQ3R5/1sRGKGrF6FYKbuJsFlVMh6pxNS+RtG4DQQyMQZ
2gjsYad/aYd7gKLOQbPAUIH1UZOlMthx4ZPvCQiiV+4XN3xaui028IHl+Hut
6AT9YS6tPu8daGUMr6iDf9dExct6zlOoLIAgAKxG6xucl2SUACRjrkfiYT8H
GM904qAktwi5KON9HHglgupd35nyKBNLizOT3Uj3gwxNI5aepnMuSPjJvQ+Y
lyVkuzVHWlgvhC4qeTyH3mplj6lHdvIm6lsNSHVUBlUHuW2TscWAaGM5i5L7
L70h2G1JisF68+9EcL9HaCTWYyq9LwnlCjQhscCxqd0fsSwXPz+EMYh+YWZ0
GqfmCkKrIeK00NyJtO2cnhSsjD9fRaczhmrJNWvHn9oboP8XTETUMxu6ZA+Z
QlrByd2SlWY53DqjCB2orLZx8Vq2rvIA2+R9A4EIeu20En29f4j+8hGQEtj+
/Y8s2uVar6PcGLEOAmeaXx83DZ4Tad+JV4XBKWtMjgWX32BI+L02BzSFkz0x
8vsOmtwkmkb9I6UZh/lLXqwNF2KlCm9HQDMV3NKneegNvliQ3GGNw+7rNfY5
9n2Ec0LjybzAAT8J6Wb3eeUU9bJRQ0k0DUuChlDI9BshcTs8gtFYz2EWamZT
16T/t2rQdUYPz6WXlGE7n9iHBozx4cN+rx5cJusfQxr6P7Du4kYSlVaOM2ea
e1PjMlgNFB3MGS6LFXzbod1fApz5K4QTMAN7PMOtRZEoKpw3gM0DKABHcP04
RbRQMi1xsrK1K6WJC0MoZHZ7Te0SQ0Pd4HsgNWUe5FS9ahpHSjZWo78Yz7Dl
08plFCMZ561uW7zd2RUhGgKcYm42gdQm+qt3MVEe00WU8cxTBx+r5Yelwsip
hqxxSLtc3WXPZwRv/VxOTCQOn57KjUq4Dsn3+zImXt7Fx/62nJx6JpUILwRV
Lcoens6ibMhn1K3RGUAUj8sOH1rmQ4A/8UNvE6Dhy65d/Dest5tdnNGiklLv
Yy6B5jgOhloSk8B7QMuSqAqCfw+e7LdXsUGj/tfBPVBeqaILySBOQ3SxOeDU
7N67QEdCwM7xnw1GIis6Jt0r0CinlvHlwqmcViYuO+/02Ki7q1yKiRhOpfnl
3Nn2/04iFtk1Obb1r0BwPuE/UBlL7+vn1cW3aXpQiIFXrgDfo+xUq5rEi70R
kOSRByWp8I45ktjeix8xQGY7YROnWvbGdTT1qbCMip4AIRWDL4vYA5rx7XkU
6oKPoGYtCAROIFhc5Ora2HmTmSSOXmQhZq9X8IMhljA57a7TQIBZ3xj3mH1g
jK+uPyajD8aHQt+NyVuwxqqkTnalP6JcVFesSAs8bPuZxJ+w3pTuehMY/DdS
2iu7yqkuV7VZtzhyF/i5LbcJxa1iNR92vt4aj+LkrTf1xSEVsliWx6jFa9Eo
McHr8gfYuoXL/ZVEQkwH+Whbvt1zu5wmCw4pAuOQQH2mmNUYIHRrBR7+85uG
apGPaEvvCiglMfxsTnWuF1AfiIFblVUwCz4ZuWk+vDontQbDT6er+lvYj6aq
KRZmW3Kli2ookpfGI0413fYQoWF5ezNX/UBERnNH9BK6t8zD0BeO8a53swXZ
q2vpPj3IFFjheip3BjjbYa2RfbFcd6ckX9jz4tMBZpoeFGHYS5l5grpuEH3v
h/zKtc3wN4HucsW5DphcuRQlXUtv9bUAadvAJm7ZM/30JPruXNYyx/qOjdNK
7VaEUKmPTkTJqkJIogLKm1450J4pkfYShRirt0Tl+5eRovgINHmLFw57k0zD
XXX5PIgvuERgNBe4hvosVbgErUmZQSrcvx0UzDxsGyYCqwQCXX6LoT7kASa7
blaMCBQVxcC0+5ZCkqYNUH0Ap/N/94ayhqQfUT9LWskp1APX5Akj5CXI73ys
7bqytsGsN8dCGplPk8XhxUoJgTfE7nbyOl8MkKulUUgpdEOEli9sDcTVrA+7
wOsKZ+qyUdFlfwI/ZuJWz0U7oh4sv6J5pbolY+WGw8j39zqGunhFxTGbPZZl
v7OrHdd+cifpgB9lCNC5kCFO27g4xMtqVzZ0Wi0qje6zyEXdOWKlKGhWERBf
h2pb8MPKiwWG3XZ28fgC9TdMF0exZ7o8oIJX9FzPSlxF3U1pWvrzls7EKLR4
8IHAEB0ukfpy0U4lMhhfo0DPv9q8fHCCUV/reoYFZ2Tx+N1lCaVunIGvWHKZ
IXy88nOExoO2n/YlP1laYpZiIo2RGb3/16Er8RDAcqOUcKFmMdFB7T6fkM2b
xq3k8KUi136XwJu8eBh44nybAMIv7ih0tEEA1S1ifEOATBYBcU4J7/YlV0gR
LT0NR8KF+5XYRh0AOsGvFhsHc6N/APgmxM37IgK5X7Zi/jlL3HK+C2paor4U
04s/g40IT03WZmaWOGTobhixbrcoK0V9aeR8YA/YgcnQEc+oeY+hhE4ywdd8
SSgyF2NbUEMOrxWDJFzGuNx2zWAnT8WMeMG1NAH+h0NCDNVlfhtpfepJBi5/
sOUtJS1nLmCEPMVxs1GrxLp+TfGZhE3dwmcuqPu9IRrzvSD/UE0djvwQiF54
Umux4bLZ9c0OzG2msz2J/o9SyuL/Q+T5s3MEDCGU6vRXvQfkrNHnb0yBSTee
5W1Bd7Rady3HzwJcoaHkL3Ud3w2/7Y0r2iCG4Fad0uSOUfyyzmsC2B3iEa9U
aoYVSjK8Rk5dR8PwON38Rtr5NdeYUD2mghjx6MD1Qr+clUOB3VpAVKMWNHcr
DKHcC3Jt+ydRS0Q2gZw6TBMo5ikxUEkW62RYsb1fHHRmMv1etEkBSEcCLfJE
YAS42C0DsU+YlXdm5tyw+nxnrHmJD/L3gNbCyFVDsgL5MHUfSifQ9IIrocp+
UgQ3H+9xzeYl9ulormq7f8dBDKSDM+Gv92oqYM5C1hcCgH92c4IpnqbZRlGh
eGuS31749jO7aW1/UhdW3eUYCKukoHn/BdSwZtE9UC8CwpkQbAHc8uaqrv9Z
NR8djFKhaHbd75dL6x4cBgDgN4eTvYw8fEKJqsD+3nYV2p1LTQjXQXbN+rNY
nYj8/1jgapqGW44HaLD0Pi5G8Gfmo+ZegAZLh7mnik1+IaIctjp/H9hX7SBq
5KMcCWMCE1OshJCMNyAOwVqxUccqmq1LvEAt9usWTzKCKA0Twt8Kty1nmnVr
CNUdiTAooN/8GP7llbHTg+Tq74ShUkL00h2OqUEitIQdcO95aAMVaL0mnBpW
U0dyqxOS3zrrpn58bYu2LQvTZ6rAZEwmXureVlf3hImmzP2Z4rLCkmcZ5BSC
wKPrlK/NWmC1dV2qWRb5r5ju974Sje3Kznrk4kmx6ETmBocYsqpUlee248R9
vgsBiCXhxsVqW+KtsXPW2kVEAwAV1TkMoby5Triyuk9jiP2dwU5/bj1JFADq
f3isCXXKAR9uDR9x7O8j9x1CpAuHqnLSkewG6gc7XMB9dVRaIcM0iKpm2OUA
UatBMRVeOKqnfR5VOZejWRdGp/G2Oe1TIQ9RUb9mvqT+HbD5czht/33jOvMj
kXrJYCh5Oj4t4OxbbSiCc54cAUZqD4xLZzTUuswfobeTCAJzS7J0+P/ZD0gZ
O3X5npSsBa5RG8HAkUrsloEtBUVNKw37g250eSDCHe3qL6SAQbdWwDmi3PX1
NrDog2MZzB9du3N2/g1UZpHlhYR7HPS3400FUUPqieLpBhNdJHpDLask6euD
gEqusxqKLVH3HgBmLoxUpuxx96PtxWlkfydXu8NQRguLsz9x7y+JVZG3PGSL
hSufKnffo5kTo4vxFRpl6pCJxYF3Dma0G4dv6q2bLmjQd6EAFz8dFZqJsaMC
3kjMp5EFAC8kDnlEAFyXG7LgLN9ghYSLNtZA/k9b9M74UO9eQOiBuYD0ALPg
qaqpNpJcCA3XlGis4CxVhpuIAW8rNj8HXPiVjiIDLZpQTJc891bOARjLVI6S
ziD96X02/e3021MsYHTE6MiKYhDqnIGRAw3ljziL5H2aQZFAOtV631RR0xd8
uu8aunkRzburetNuVcRflB7HYTsVlvBT/B8QDOZdIBYq9SbaLDWjagoFJEFS
onudlxasC5+EUWTdWJtxUWqSHgYC4w7/ACztxn7b9gUPEuwJmBkyS2SC4ESw
11TUWbfk4mExS1YY7wLxvg5aK7qtfGrZsMaZwb77MVz/0VOm9Qh3yYA4VQwW
2NQzapRRm0xbMc3t+COhYLMpEtGXFxObGMqVUskCLHrho/GxoayM8HFYQ1PG
kMh5V5OawsF1VLU4CAxgiLBU0aemufwzBEmhnyY28FS2SdNohxvzr7vAIjS0
Hw9+hXlA5DvNQ11XyHTueq7ZjQQZIgGc511exl5u7udtZhJ5dmNn2tNluBm5
ofPyuvgXDZ/9ARWUaWTr+XEc6pnTxJko/ZI9YuBS7IdtfSDG/DAuW05xoZef
Ly0CHcVNJY9s5ijBfyKXE/VY967aLUV+JkUbl9x9DKRER/emYxOcTRv5fVz5
2UYptXWxv5+YWGk52jzs/0qkHeAFBY/1rzUrMuXqoSrMDi/gq//W0aOdmK6F
vmJHzGY/rixD6sjIkLGpvEVgZIKEaBDTyECH+LSYbFSdgfv6WHWvh3wKSoeN
GE/BR8q1DiTNx0vBEsKCXTU2OXmTe9cBZrbd+GGqrVZgczInUOxz/KEdnLg+
C+OywnH0fMRd3EF2MkucRrJn5It9v+Ru97l5zMtk2QIwARIY9SxLzk0wIYbg
AvJm29U8mDsB3LS6FgyMbkeMN3UXExIk1C3hh+vKzjgxf+7ZnwqELtX9n0wG
QwMLLeofbm06aya0Mud5c6PF687Ow+lWcNV93ewwaYpxHQWWpV3kbn6MvBs3
eK84ktCTmG1BktmPqB7ghtfdKAF2Xcyo4TnCLqnHS8QwHKk84cBd0vGRXX/q
FSQGlHpco+8Q+4thysDrQ3kFRo5BysWc2Ie3iBrg6SHoBnUj49cr/tDP0igG
dNXtP3+gtn4++CTiVGJV6UD92SX+rv9cfqtue8qK9xMw/UmR4l3dluiEIZEF
PLhKiZIprjKGAiGxTgsFEwRqOIYTRKTvQmgcbBkKalXuUzgOqW9NyEiAhGos
hItkTiLmF2H+3dOOGSt9sFuuTQUaIP7045TaAAdo0JLXrmwW1+/IgbGr62xE
JENKQ2BBTkK6kO0nzaDcKieHCZagwZr9JHRAAjA0Xj55UExOhgM212KO7BEX
dGWkK39b4U1EByTpJbp6EDC+YZlskgh1LfBNiVyBYQEeZVs4TKHkWXr2yUH6
9s55JT1xPk5gQVbK/V0mEzZaI+kVvmYi/6bkklhChFxVDUflbft5JXToL/CV
foxAlRu5l4/yoBdPjMC7mYNl/K7lfVbXOkVT/711+XzXVeqNHXDckqhoLFWN
ObIxs1QhpDRgK2NzFA249pDzFIX+P6kLlXnCzZ2njMIH0bned5iGhR4E6no5
STIsKynW6jFs4mZOXUlvUu148keH3y5toHirOdTaPNO9dLpAFp5MMwaPNG0a
kobzA48X10bRzU3674ttjtC909sqMc7KUQI/qM0J6jRpQtICqaTow7nbU+ZX
ZR+rinSyAtum6IHI5IA3Bll3p/9TaUE+3OsJPtpnsEn5vmV0/tw49wjJLIBK
hfZmkF9sPcTv9I2mtr5FOjOhbhs+xGQjXFWtoy5ANhDS/mE4NkUThSjCub5b
ivV0u2jdQviR+2OTl0U6cuXE1YMlsfAbGE0l/scUy8R4L+A9BGAj5Gz5WOnv
TlwVv/5IplOD5ufMRQifi56t6+E19oylzDeOxLNC20R9cgV+Ydybc3ICdcpS
30dAQo6GEmVn7Rgf4CGLsMBaOmF4bQPu0RCbAHsnlaxTmIrr55r/U/hW9x41
JOCBDRzlDiPR+xCXIgpTaniD/NFGrk882dAWuMCQNQDkrG5SXfUl2Ht080Mv
1vF6K7nDRz45ahLA2jCU9tzuwWMXfJ9zNcIgsfxVZAPX4kRNQ9hJowJ8hld0
kZjmhifh/H28gBuLBro3wtTgQ6nSav2e57Yywa09qH9tLeF1OjjYM+b6ipPs
6IRtTTCW+GjBPp0BmUlNeTV9YhDZyRg/cMhO614AT4b9VpaauPpsPwKrBS2K
P9tNO+cAUjzvZAta7ckRI2YQaYzS+e+OQH8amv4CllDYDxp7AwTEdup96F5U
1j6otDr4wjC/llIfsj5LkvyOmtwe8fLahldR8YvFwVRv6z7n9z0b0hCUDBMm
MAzxy2aNMP0AOUhvUPh+LxDOIS2PSp5qInJO5Rlf7bYdZCTSVkYL/GVgDzOy
D9gfwF0kwu6To9mj+Ro+5C4FQFRb175eT87Ff0X6WWCrJb9er5PcDJjYJnT6
6/T087e2qTB7zT0dKuqFrUqtkJjOsPgm9MEgqOUMXhXJi1PoPx/Vw3Wd0MKD
l624y995WUpS5OKtWErjGuxZwsAMIqUkRudniWEb8cGFTpTKZHztqp6lKTMX
vQk2/e0D2sWQf6uZfKpWuVofhvUpH3s+xBrjPS5DfjNN+oFQORRbtFiyBUKR
dD9XTcyUvJMnj91N8HsCEVYGdfBjhPiCUYHfrmMNKxqHaApR+Ti/8ff8KXIZ
o+vUIsS9LFRDqShIZqZgIaBoSgbeVGcye19kPmCRuJeFfXLIzgG/S7kakj0C
8cPlMHaN/haFnoU8mTYZuorzEUcscsjfv+Ao5DalmTHobXe6RYGdMZ+CBAth
jzxzDIoNvFu+Y01G0imy0S6r+CpjN8o3UWdQrk0auGvOBVPye+N4s+eNUmEQ
b225XCx9SMtGGAcT9vstid7tI8NPcTOiXZpHFzJu5J4efgQxny1igF+UVX6u
sbFOVFTFzBp1XeA9FGECi4C8I1yUcW8iYDNhuteqemHFBdCNgj3t1sJMq60j
v6MArryn72sa

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6Aro6OxmWNBkKlcs0Udm4ySRINTXYHmF8JTFrCN5CZ8e/3QaeZb2PmT7x0a13xxACG0hkSppHCGN8BF289IGH79VPV1qTuVowA5vqSr45uWCYvSH+2GiedBm5gfpT8QvLca9XeWY5N4uu/2eIGBgJo7Www32JpbSe+bG9WUHnSZzH+OsHD+19k/CqV2xKrgXIRsmTz17obyOS8mRhxYvHGwB31/T4ti0BXolGkFA+VjEwIDwaSZfQdZCCj7Np0xHqXKPZwRcyqh0cdP7Qqd8IalAnYXClRE2UAOV63vfnlruxeE7jHZTj/qUDZcpJn0gIp+9PGm9d20BKY3K6AIXL2D+TAFJFWE2UDfmZjTR0UAppgoEOYadR526PAV732LdtKqhgI4sCs+BWyxPdkESx+6VejOk0bOqFe7/RejyoWR742Mbq6NAWYzTYTkQRkJSISBt79NDpRiVJpfuRdDkcjaB3aweWQqPhZk6fS8ezRikP1Vgg0bhiB4RqEKn4PBxt1a0kMzoqBpSDt+sID7CodQoLden7V4qsm8/M+LIMDOpLjYFRJsbmlWW55LPIowB8hkpV23yy1Frvu4CokAfiWcrEJKjqnOMuRsAi/K1oWaOLmqQsLC9NrhtU1PzBsTVoq9emAjzmbPqjA/ZZS5Syr1kZ9+iZDjvF+zpU1n8YruCe7SOV99SBZScLyKY6/GTPX6QG5v3jLc4Hsf+WwGe0QFU231A/LiAJLAAnkZjy93M00iesp8BBrBvTDfLIZ5j7UUf7pKeR0B0iMVHRmFK//Y"
`endif