// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lVpU4gVQEZSwVZflxiUA7LgdZEBVA4kSVfJBB/N/+kbfj+Cm5QxnvCm7wQqv
uMAGOEJPB0JGAcnSw/8mY3Vmi9ld3h/8ZUi+bIoKpeWwyp7enfP5nzifCrUV
FJSv2/7fcwVQQy3R+VCDEIx3wzZ8U9QwUPX5RriOK+DMDVmpq86WW3dpNqfz
CrHJmsmjYBlSpFOCmEMbwfNSTgpLjvepvuKWktXSXQCq7wk3pen+oUP0my75
xRFR5keTNMmJ85EUYHk6WVzstmFHmFdRqi8f3jSFCHg8L0xrRrJJx1Y0/A0A
/JNmufoo2WjX8jflYPZJb+obojl/c6uDAAL0JtQoPg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IoYaN6m03XUgJUPzNV0woS+53VQKyaj9ZgvThCMOjXFtBblRDlJZVIso3Nq4
eWcOct6IUdJV0v5i3Y5ELNFBDIgtv/iuQIaKmRDNBmanQmNhK3WrhA/ZFcX8
U4lshenyCRPwQzMOUM8RT/xrMkrlwJljmfid9oltj2IzEdoudS3YRO2Id582
yjye0Wx0tMlVXqecryBtXi9wLkEQWccL4MGQOCGUYTNGbG/5cynPjYbcfIa/
bZ/95t8JASe7bWd28zCcsEOR/eVRMyOA242qGPyq2BuTCLJ3HTIBWRzIY9ec
KrlIhUM3kmNJxb51saXd/RnIZM23PjT4upzZ3UOQuw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aI8UjEeotAxctAxtR2m5z4PFJ5hJwx52Z4MAv0UhQEyuSQmD0oPuIJg2GESI
FHHSjqyTtRQ5ZGCjdkyFaRupuTrvVD7hk3QoEqC4RpI6xTcO08OXn/ALkXG1
gZWUHjaXi9NMkMaW4DP6lfgtiNOLLg3eVPerLGOFAAUotecvyWBH+hF9YFWk
gcnTRPkqZIJEzBxXUQUNImLMpGv4CXut24rW2Yo0Yagn3Fv+hxddvr3YB3V6
2ALNowcRvq3AMqt2bNorbQasbwDDFGyKMKuUlmSP81bHkzgfYttuhjMCTn/k
woqHL5tQFrdYXqCU9skz889JUV5Pr7z9h2EgZjCtkA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KVBt6VXu6V9G3LyeORVu9FwnXL6E742vbDdHvQoWk5c6G3ipB8pgd1XntaF1
FmGY8/D+xf5JQXsfgFJXcFTmxABpPxavbW06aACwRAEGGQO7EelNNFNMGuWw
LCBBl4SJs2ibBWU3UcW/wuTh3sLoXwTjHNgWmnDAdFqbrhi4aHfn861Sh4hw
RRAICtPZv9JYZDoma74qu3/dlrN7nIyToflpyZk5Eb5tlDp36QH1a86bym4T
oGq1FWYRFdkydbFw2RC/+ox4RKezZByGsL9vlCHsBwzfP5n6+cRFrgU8xH5N
lI9T0Bh8EVxz6/5ZK0/vuevM7Pwt09R88MvOxwfKpg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jsESK8zQldWFZaPeSFaU7VfIFfHGi6F9yw9oPjgK8RxWsFkExLMthBoMFknH
glEreCcufTdp27Zaiuniom5euf5DsO8Lbm46yXcTS0SshpxQ+wOzuPj7Gpyo
KX09t3iw7gVFiKW76edAvD0o3HlF7KUO3ejPMREuLkyvR26tLbo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CCZruaGHtAiYtI2n0JFXHOgF8iBm23KHQiFY9KAngb0NNZG1B44a96yleFdt
Nf7DLDa3JLCJrNV8XFxSW5eEqh3Pxb4mHXxtA3ZSNxHcucb2MyiVoUcy0WPu
oVmxp0AHBYAdmUsSPAH9+FKNtMAAyNsjC8925ZL0SvAp5ycbMeH04W32A3aR
AfxAo9LlPtWs+6RxSl40/NUR05SJeLGZkJGqmUyL3r/w5TJySQS5Lo24q2WH
Drh8AIaGMDiZ3gVbtJjiWhMGDKVjyUU3roL/cQyl5SdKVnwdr8U7FXl6c6al
Opqne2FrfeZhgNt5C5rBxbWbZ8orvm3RJ4qgwUmPuaCizDgksGMc5q62tzP9
AbuFLQFqvjUAc+gYVJZB7E20Xnd3N0BNXnk+DX848EGJQfYU0XFL0L0qa7wJ
gLAk8jY4J0M9R0L854HvamIBDwU2k6eWU8qhSu8XbOGPk/Qr03FW9RyXcJWP
NmbZ2t967Jhkm3AdVFF5L5wQGh9hLAUL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
T04P22OLAE/idFS9AKJAgR/E+t2hGXQ4RaBpWxyGKVa6jJXMpHHyChZTPxN6
V+fQGAw2I7X/6DhMf5wsb9EB0lliB51bNo0RlSCKEjD5HN/0sEnp8iU/PFfg
pFEdWJoPH1HSE31FimuDmKgb7+R41WqEoKXAf4gr7ZAzpJc/EfI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tl6N1X85zbc7lWSJ6fP7ltTe+kroXQ5ZcrQONjGjvvfJv8dUbZ/OspnAXZXg
CUtJWkY7yP5t+7CIV+DMN+vUv2JFCzQWyNOo0SpTp6xbr0ru4YZ1iDBT/hJ0
Bnr+cXUHE6hKW2oXssFS1bR293jLJItySWqBJCjDlFjjkUwt1tk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18368)
`pragma protect data_block
IX452EkuKSqVjYi7WCQ0KsQ3gbOq2zT3UKNaa1ZLawvdrwXmNmkwrOdY0om8
vPytWjwxAAgSCTSZ1+A4oLc0ZtiCUwWI/8x7zP2mf+EmJdv0JuNpP1GCzZ9/
qtmDFncxWH2uUyBQAwXEHxcrJnJybYCKHBlakFkmNosMY+34bjG5CCt51AGO
Z/H11noOeTXcsiJlcu+r5A2itx0d97f6DykKtdrTq8jBXupuPYMgbGG7vt09
4ZjHVRtniJ1uTDcFVsVpOFVkviKxVgiyqN60dxWu6lJGW+RZTjWn6nvF+Qi6
BeBbVXWbZUI111yv9uc24wQCg1FoomfLIiH8uw28ZRL/dMGLg5CQBXzCT9wF
2bfQOWr5OPYnsyirlL4xAz96d8rlphKMdJWUazxrTe05ZkAe5caEX8nLHahW
OtSIhxGfZ7HHp7EYcFAXMMNXVzyfkARSSVs6rua4aP8hQWb01QPcZQWG08qA
chhc3s0Qo+7PLrnHhHN6RL3Yjp2bstyZjvBYzPnBjd6sZo99GjczE2EQ0Gwm
BVS6mviptG6CfETPhdBlO9dxAKdFYjrXofTqGoJe1w455m6CA+j0+X/jhh8z
yBLRyLPjKpmjyVGmtAwuCl+pVPymJpqPMAkq/2AC/vgrC88OIDOzqzUxD9yb
Ge5qkfH80pLcVEOtAegNuuupAQ6FAoAOM8rlw8tu27Vpx1RErfP5a0t+l4Sl
WsWlz/3/HbpyjQZCfYZqitV3m7/nllA1S9znOZbaI/28OoBa9s6PIpdBTxeF
MOB6Vpb4BfX6rZ+mpGeHTTRtYqgapooGZ/O0F6Vuri6Jw1YDS9ZKrJqjtteO
t88w7yWDxipFfRJxJ4zlDhio8KJu2qXVFzayOWrd8Ums49movmIi9THNq6B6
MjAO4VrR2Sitkcvo/LOoDfh6assFxMJRN7NxguOUqQTDOciqMlLuqHC66Zih
IxFcgVF0w5K94AMpk9UrFmJIDHuDxQ01s5MxJ5g1DxFREv4DubQSW/5v42Ud
L7JA176hLHqgMUV3ezMpFcLXOvzU8MQdaw+EM/0yomqJ7gR1t4SIx08k6H+T
A9QCRVte05YnJcpccIvH4HznCPqKKCahtplRevDOP8hLgq4f+TFRapZCUzwI
aUl2lx1z9zf8FMHLN4g5XEMZ3sOmaQORIOjQE4cOptmb6YwZQGTGHX1mMCTJ
DU2QbI8BQ7xKBDqh6GLGyEHk6p4kvZdygojua3h6KclZISo89hWbb6ybpiwl
8FMEkX3sKZLWTbH0WwJEQfHTd8DHlOBebtqi+N3ov0i83Cv4cYDgDUZPMkjX
1hRtle/4TMR7l0RTPKC90D3Wmi3OFJ+k35GbTE+GhtUMV+fXBA0QEE4HDNjZ
aiHR8Rsd8/SDXr6Pf8+rI+v83VR3BLaPqNhoDoFx8IiotgFLK8TCKpwP8BUT
BwQ7FCPqlau3OaY1uaJdjx/1Y4NcLjsuPfm+HwUOs6sZPla9QGhC7EK6jUmu
J4OD7WuPqIx9iXf/D+2uOoyoUh6luNC/zcj63yiQ8v1qPoY07kZO7/stsU5H
yPsjqd30J/UtO7K2ssTVxzPLacyTEgAiwxOS0VYRLW6uZ0oOdpz3KEJ7MZ49
fH17JoKS7jvAFKyZsVFIEO/z7lIzIiMO2Vf7o9HJ62MCfu5Lp9ikoTnk8dP5
iTV59vY8bn6sfrKtIdXoi0oxrVb8JbAkxOgEsm83O2vpqAgCv4vlyVtiz73b
v5mMKQz1+ADTVTwcgNpW6qqgZqatO+8tDKfNBEl18QoLLx2CH7TwhfIVlKep
yBrJCgK9VvVt6U3s7WtHhjb0pnkreubAg/pHA3/7s6mkJEGoN+wiQoYMyohF
+O3NVYszCIRF+BuhpKlegv2jdwk0HnVONciaC9rtZEWSeb74mEJqC58ojiv7
JDwJ82lxdRiNBUynLvJJzrZix8YDqo1kInnQpJDfVChzVWP7pw4U59tHNiTL
ptXBTSlaShOnzi5b4MXMPwVO3sNFPPOf6wnRiV9Xa44PzWGdi08WDMO4ZJg3
JRbeJ+kfzUp7+4orn3NOXjILRtuakGmO2hrwgQCduJ4l4/MZDGctmfTeaI/N
oGU3XrMam3c9IKvc3uQ9jTk6HKFdVW+S+HES63WGHMPcl6eWjanqy1KCUBOU
g2I6VUf+QfpNidf+0jwT29y0kCjtFAbtijIk+Yp4Ua8rDAfDwq0QNd+VrGmA
CgEp7IIzpXtrDOrad3FIsezoAOmvvqH4BpBZ/8jnjG26qOsecn6MSXOxTPMY
D15PBzTXJWAevs146c6xea5DAGBoAuEHaSrXw7CJnlO/udwWgnu7LZFQ3ML+
vbqcl+7IjrbrsVlkm+BELrg2Jowth+yZxzzxoYnumKz9Xe09MTnC5SQjeLa0
uy9cYbT3gIdgx70eVfPs+JVtwgCYMCrM50Q4/PbVy6pXoWpR97acY/itpXQM
8F1ZgfDp3MNQIriagfS2FubJ2vFlWs2Fk0Rc9V4ytHfZ9wBlR48IZJL+KKDY
ASie9wPjyIz4H+z14sU9NTkHPhb/xxKZPPBZPa+FOIEQgxCUp6b0nqWY4vwJ
pteHTq4qhISNZO+6lK+gS+SFGJ9SUzLPVNwXTyuSmfkPGNWpc5JqzCUUBpIK
4WCBdyHEmWugd3aE9Jez8Oz9+orvmcjGxlGIaoM5CFEzh5jd4hR9P+Muz6Vl
/fxgjYTk4+vZnm5euRmVUuWd+mJUXF3MCDG9JVi8Po5djeS0ha+aA1VnzNpj
TQx1oyurxmy49QzhxTF5wkJKBiWQt4Xoej1WPlc1tDJmwrM2gm1epez385MF
66bCqrnyaA4rH2wqj01bxQGtaR0DCc6eUzL1l0Amm2TcgNXTi2CyAewjPbsL
/cSfXLYoC7llrjtZ/zlmQD4GbN8gXjSQb6heKQfLJD+IDTml7wF2glywerh5
ip2pgy642THg7kwZg4Accrxxk7tRFR0nqgH46jpWHumxMRa7tKXjXetK/Rrq
/g9Bvu4ruOLVNridWsmE3ejzJItId4Q7lE+5VvNbv42BZjbkiaTSNQkhC6pB
c1M/aIepuMqXZL76ROAMWsOjgUbPoYlX6AiJZdk8HitjJSwQ2/vTHhzhnTVa
3af9VT/8mmGqyRTS8v9h650BvxDLn7n3Fu35w/inHHmDf2zKHF0d/Z1nDSr9
B3kdKvKJDPAebGJCjjmb17JUlulZvhTQD6Nj9MdlV52nTbBNyYU+bWzw5Vm1
kDGP609JogSGFJYpoFf+Wv11XxR/YRB2gI6pfFdvWQwaWFENEAF13Y5uAtlA
ajOoADHRfLcFPYyXpNUlVt/S+Oo6f8wtaa79tIBDVHD48A91fqimDiqN60bq
ZgfHdlBwYlpvSI8Nt/qQU6rb5IZe8ZqAnGYOTakbXcggcuFCH19JdByW86RP
nUdC6KPc/CjQkijlSoDeZaKugfEMYxjpxSxWGoCQmT+gOzVUigY8min54ZxQ
cMvE9L3DYUuxSN+YPoFhzbPGa7+yvBbvwEcp6DzsSEhxrKFY4S9YYpgm0UOa
oJLq+atz1cEJjAy3L/psMa08J8/j+7vI+LxObL2dS0h2Ev1jsu87OkOGWfkN
bMAPjoqqfcITOycPGKcdc/5PIazlYYbfeCyV+ty2DmMhajBLKuxzcEWLSKtK
Dl2QS4Jgxxwy5NFeJcQ1rQtF5bhJy1xlKQja5UNMoR8r3a96xZ0GV6Vupq8d
RJ6xVipZp2FF7f9mEu4CLZzyfe3QXx1+AtohHIKVeqRm0lk16Q8Z4uFTelRg
ZHidrYBRDuDE/nVHwNS3mQyeSJoD65xvAyUIz9D04PE7xWniTv7O1zxrLqX4
bMhHnEi82e5DCng3x4PfWnpEvbRbxmQs4War0TUwM+6v7q2reGcIS5vWpblv
G7N0LcsoU+u7xYSN9fG4Z1L48tTEcTcVUiH1dcmlhe/O5rN3wJhsfZRtmnSp
IQfZ8Sgl136GIRAmO27ILbp4xFPXfj+CDdrDSe1J1cTN2ALB5tlJnuh2O9L2
MMvylHMp5gGpMfwX0Y1j9uMajWyfBsL8qnKsB/Z9LcZ1pY0kD2JpO4fxzDBD
5gvqkOfw+RcIjI4NzxQSjQpy6MoEalhuoivf/lr8L9FKfmxlXsz/fdNslihY
IaGOeCsZoWYQ7F5g++es/Q7exHWWrUqR2juhtLFmyrFGp9tQRIaRExUeiola
vWfxfKRH5EUoi+hz6/vYf2UfXndW1+ALCxb+SvCs3d+wAPScv9rF3a/mKgdz
7LaZcGoaVw8oQ83PZvqC6XFdORtgxZYsL3XshyiBaN3pJ8wezB7+Yak+ulym
q2Pbxxuu5EEVe1ECtR8aXXebvXTbjn1ACoA99Ow9DDXjiZoXK6xGfa1ecz9C
0CZw0S0G7Y+ClIubu+CyVIrCqF3Q0zo0JK2fAfYzoXVJWfdjMczyxhArzJAg
rr5bj1SfyDB8CC1gd8OFF8tkC9GhZVvprteM3hClkMr6nMtBqq2jxZGhipay
MWP29l05VdkjNI9AI3XwXpqyfV35bJUvTK2TlrUiWO1gtq1yD9gKwOJh11bF
+Z3CRhotxuKDG/qfHkFDkS982Bi0PLdCJWpvg1GXvx4uWNIBwnYaH9I1kf6n
fO1+5TVEAM3Q7jojgsrB3kIIQQwAWlZTg23hJkizFh4p4T9N1HsHQzraYgle
2t8iQGIyz/XFsVDzM63ZIx3jPxez7yVBuY/P+TUSEyBJccEz3B1Umw0dBFSc
PcxRxKbNJrd3Uxb3dtojUNZRhRjTcP+MbrGvv2nCkkEdfz52HMnKrrBsGX9C
OvKWHI1Tn7IR0Hdim6087DkuLIOz9EWA7OctwjoaZ6wpsuBZINT9Ey87xJdc
PIdel8bK5WsSsyoXaTawg9rDAcFq6UtjbnwX6QgcinejRnX8y6tK9kVP3BEc
ti0zSDZ4ql4cI9WNR0YIaup21YGqSXudxMvWVFPPg2uxY1MLSHf8GBlfO03E
PWuc7Wxct/hJml8YywoftRUmtXLfa+8L+xYQ4RYMR27g83M9hfUH2YwyBQTa
3UXx/4z4hE9LI2mq8leu1yxmO1JX0SXytN3gFWGKxnTo9vm0myx/gu1IAJBl
skELthHjEIVuOYSnxZKR+FZbobfXg+yzesgEYC0DHtU/gGY0p4Fl5SbUS9UP
N5GgS32IhyXA8td8SLhTtqfbGkQVSDuHqz9iSfyAQMV9SXOnS4ZgYj6jFQmh
dsAUXu7xOs2hOByGE3soJb/VStB5jS7bKQzvp9XTH9frCw3OV0SSAXSrsQC7
XbjmerxOJ1DJGDn8iphiV1b1XSadJSBUHz3f77hvY/udhbbdup+cAFd5cMrE
Kqfm3lMLjTXNAbpv7XefN5cDeA20eaSFe3JdzsvgKfTEe8akfhbrgS5IHeF2
DwxEqQIPuQR11zArx+mUoJLqmvxJ+NRwpzqXHSttrAo3zR+dKvWvs1OfSGwO
mXcgyqhQGGv16E75PBQ2rv2StukTUNHJlJ4ioI5cFz/F1lnEfdB3pkfDmuMk
hgL2dq/sSnUq2JMrdkVkZVi9sMUAREtY3RxIekey1zJcKDJTTCaSWEzJqOR1
/OU0q0E4XEYQ3s90hBRXasGrA9665ORbYx7EqMkR70ANaoCkCuo2sGrUMB02
I2KVfkFBq+fDZPp1IDxpTM5U2I/KJvB2+8LwCCz7NImvG0j2mpcJ3IVTBAUm
YOtkZ/UITLNG8y42ifgmsFoYdON1iClgKR3sxq00FegrHqMDupYNZO1oiD3i
oD6IIsvt3baU1RIhFahGGUuAdQNnq4uGarFUVoi+teDQIYXfr5xKocIW0nKS
vJeA77jiBUzPIdK0X9aoUmL3B7GKLvWTReko3oWFIUnPX+0U1EXadHdS4SMJ
D5+9wdTYyCYh9DwpkNju6OT3zWLysNlYhkVesYPFZqfTUh0rQ2yKm1/5WTyv
2XHbTLuRO4tpscREUqzYRSZ8qy0AbU7EBY2im6B7yuMOrx588/fFqYMmdxeh
Jc865lZ76WVGhnR47/D4bzKhpM38uZms6HuHaKVGpyy5RDK8C5Bjth1RC10A
MuaiAQ9ahaYTtQwOU5dWOJNL7OX5RPWHZp8AGtFScIzEoK8sNVboBZAEdO2N
iihzW4nQ3HDa9fbgBFDlKxZTSe8OTwQo8wLR4Vgf/ce/SEIL6u68Mg0+rpOy
A+brjRU5Yn9FamqCZ5gxAAzNtveBYrIISjLMOBBI43D9pipjfR3TGe2ThiyW
irLultoLmHe0lbqi5rrm02iTLQk18l//L/z/MLpMvtMdHxKb7LivHLS5s4pP
vZDZA2Wti+lgDN4vHJChxTBAw9OBfO0J91UV9OrqZQG9GdeRjpr6VpS1GSFS
3oOnrzVU1tGSX9pl7e+ESmYWdTgoimN9XuwnxF6sYs3CXfySYNPazXMAYOBQ
NscZcKFmUDfWeOyjNEM/RHverqjgaId05IfN9LgHES0LuKkhq8Oj3vnIwZUl
UIqt3d9DbVWF3PdabWgEKXJpuzjtcrM9QYVzE6JVrZlkA4hFp/Pk0yVU/qor
9D5TTT3ys54eFZs4ihwnoIgduXa/fwu/nAt+g/IvACJ4k7EpUUWdsalHEPkk
SzpdGJxfpP3QLC8XgD4n71xM+DW6dyhpjH8g53MTafAKnGb37vFoxEJUiAei
VLrw4cBeOiLX5zQS8tTvG8JW1pHiZluxKjuWJ1odhj6MsWYDBdLsTjjTihMn
VxYpv3NWXtmI5rrdu5OevTbFOOM1mh+ACbUrG4OpacntVrnqtKRtYputXHjP
dIXbvEOvJAmmz7SDaXWBZfEf5zkzGpsvIU3dHvZx22yMPifO3PnY42V30xuy
CKo1lD4iG/5i8mvBXhF47SBOJ5ClFo4z+ehFUGeFNZdZlkWufBg5mzlJOOy8
B54Ece+DCxIDHp6n2vFBn0ounauORbACVE4EA1rUOmbeD47Mo6nriLaU4U5n
Rtb+b/K+XmMHIF91/aI0xhoaGgIDtKeynRswMuVfAMXqqIR6IqPDB9IoV5j6
SB7Y4uaaGsD8vP5gfzLIBGnNLBzqAlZADGor2xYEFKm1s3GjKEwkUlenblMz
LaMask9HRLkBrsJgm9V3wr3vXJuGWeyoYzZR+WOIq4Qk5cB5h1nkDxoTwtjd
hFT9JIr72xM3S9RU23DC3zZFykJ/m1x9IQTZX4Bw4I4F232xUN/xU0fH089S
lgGJEh4hRIKKUEz3ZOY3QT5/uSoScTxqRhJrqBS1TaBRVNdeVmzX0FUP3k7s
LD3L0W41pSt0IGgkHwHda5DY2B2jzcbezfEVJQkpv7z/tA1OZWPqSLOArxNE
3GlRWXQXmhuaY7i1+a3eOvPpnPZTv0vuW3qXNgVt0osTaYG6/n0Ccik2oQjq
GpDax211t9fizwrBbZmSyv1JlgTnCnAdPWpTkzowF2cPPWp06scc50CtFreO
3JnJB0ksIISJCdwrPwuKTsoLnXnjuGh0mfakkEJQv7YOtIva65C2Z0Z2QYv+
4x1tPbxP3I+Kqs45AtQZkcaJ0G6VsEuFx1pWasvqSDO5YrPw0i58PxxLjgL1
gVOokeum+f1XxMMjmcUoNpwIp/jRZhsd9sP1HxE6CSnAhVBJPGDi+voOQVJz
C7xmU0Vp/ZMeCS5YnytftS+CF3MQ6IAbaYM3ALjA8jZYL8Xvd42E3/CEJEwr
X7VYUmAq9/KC6qe9GZ+dS/8G5lcpKUqE31TaEzsn/3zb3FUr42c9/ers2lKo
xaCnFBpXBUSyRqN5sRcd0vDS8wj1g8nuQy9U4/gTqrG/ZhsNt6cq2KJzRfcS
aluGCLaYyn0LQNlU2/43MVLytHkdnCznG8RnKhYJr/bLOp0bYUo2iAOPX4Df
6HXCrRH/LOasO3QqaMkzekuh+Lwi7lwPB/+i+aEUm2mNhIHHdwHhD3mNfcqc
SbaegmxYqTVocQbDmTsls0sJly/OYz5ZHp4S2TR+6AX+wN3CmlOjcnOl0d/X
j/8iyYSH1zQGMiyWMoEetBNq9X4h/+WL1xIMDdbKUUcOFTx+iVqcV2rqe8IL
No6+6UYn93MAuPNg7K3h3ps1Lbe0Xrngfy4z1RF2oOKHVifttsGXRQOciVVO
nnU4AiGILHhmGzRCx7CRCTbKMzm6rVwHZWCcrIVr7F/1yzfjm9/f9xQrPH/6
BU1OGjrT+8Qo13h/ZTKug7N3LcLKpPyYyjlE8/Hax0z4oCDjYEBfk5DWKOCZ
b3U131CSxuZhQaF26BNFB0gSPvUnkoxKyaOTg+/ZVYTI5c1ByEspieAhWfu8
NCOB96MWgLt3ejX/lWsKiXhWG4gPvRpyn+WSIfkhQYSPnhlQpHt7rTAftxYF
YTJS4IA/UEnFOQOlOksAykxJqcT+iIJX/UYMTLZ5JiFpSoO8JkRhxtTTpgBs
ePudGduceiZdhMagBMh0PWfWulgOdATF++s3eXKvoXTHARfKhlAm6sCaYx2q
5HUSPKwAmHw0+NyWwqbuWt/abv0HdeanBxb3jmwP4tTG926Ba80BzM6AJc3J
FRAN/UVxivRVGf+dJ4dR0x8e7DilZ7TpQBYYUSXaLtbes1dOJ1591MVvLsu0
O8eYfb7Yq9OXkPDh+X+iDe4RzT2UOEuFoU0QJku+nJ30hhAViyvQXS1uKqYU
09D7Gkkf3hOSWjC0NuctB2qnUqCxriUZZ15xNyImb7pkwHoccnIdo7ba4lnF
bsqbjy7esySc2u8lYg66pJ/HSaVWPwEyqcQFTuckkiwwq60JBjO/f20qtEp+
SlzexGLxyffF8NeD+wwbKcF817o83LcRqiJnJPPxF8k47URJs5UyHyFH3hjG
gaydXvg+yiPr0zVE128mb/MmZDRtGJm0UxMxthLrz8suLXdTTCdEJ9m1Y2S+
fhbMF1zp+EGBs35zM3cDgUCo/gdD0sEVFBnpaOhojocE8xwuk1OmwNxfAJyX
HB4I+6BoPFmdaLEuvHGadXuVZcQYJaKGl22TE4oQUHIan1/7wYtJL5LLSkci
KCf3+ZSmVR+awbiE3kRMDenIKcM4e+zWGSkdKF3Nz42K+VbL8KQr7sjV9o2Y
wxfQjIjBb0wtGicAtyhECsw3uGSef8gRqBcEeDXdPSCBkG79YRlXsQVo27XB
y8+3DL7KW6V0uRmhENRqj6cbxm7PtgjUZCO2AApjWN6C3+pRK2S2v38ytcBZ
8yghp+iSNqb6WmSGHIWUNNkbhTYdu8vUh0glBgpNEH07A6SCgC13tchw+h+Y
3ib7M4dUfTGhxZ/c3huQwO8viBjd4g638l/SgwDPTEIG/+AwsDo8OrFtUIVR
Rszyazak97Q3IoRVTwt4jD5QIGcOYFmGwP4kV5Dac251XsdkE+c3sZuO//Bp
Nr772c5roG1QdVx8ni41LPThFylCC+guzZYckIsGiAID75a05uLsDonWXhmI
gu4QVod5/yNRLGAP7wkqmPXC0ZOMfS6CsSSa/kP0DKNwgv6Vyjk8Fjthq2GZ
RFbZLRX8OBoVKKrwPQx6qbyxF6kdM4Y3PzD1PmTEVZaAu1dRiIAQdwsA7KTu
dOuY/Aqj6hSWkGG622ZyZxSeOTZNBUDy8Ds8skUfNsRn9M0gCWccUWsEygGU
iBoT14/N3FsJ6VRT+yaE9gJsPPnNc2W6iG5YK06ZNOxAW4L0kSONrFDnbSb+
RNogHl0/7QlvGoWswTwbJj2Bq/kmW8xSsnJAsruHpQEs7smlbU1qcr8Nffv6
s5QgaSPcI28nXPVBN9lR+gLWS8rmJqlFOfU+bQpOPDR/H6qVNejJlMwKWRVx
Z2lJR6nEP/W2nz8ulSvaiAg1uOeou1ed6ozwvLE0cATj4tczfjFiMHZ72WwD
pQxlTUaFMFmHBBLYfOoCUbnz25RDw6jSqaQ2F+WH7vOgMivlCv/IjHT/XyUm
syEC9cY9WDMUn9gf+x+twsgmcrjgG2SpdgUvvWoorf4eDjZLqNve0zbHRv4Z
W51cjg/RMlLVgfaaeEjfN3YUjvZeK+vdpm/PUU6ebuEpRYoUEMs8ndwwMSPD
FU6WlDQoDfiDxviE2GP0CGo2qNOIOYKflZIdKWMvF2MfZW6VG9c/Z9n0c6s2
pxOMMW74ol3+RhGqQF2wJdJPVLS1yMO4NxrBAwoCObLHNb1vzcHtvnRbwNmh
QUqzQwAaU41+6mr0Jhf0AgVqR8VvKTwnJzVBlGAkRrBIPjd/4A8TH/U524Hp
7groV3H90rx+jDV9U/zYdIbKdv7lwTMla2FvkxjvVwXOGuZQMEmsWX3iRPjT
BIzJxYtPw9rETN2uclyw+CLHvZRKhKb0wEOl4fK6CjGv6u0tX6O+nf21gvaa
JAlJOnc5sTVBRfL87FZW69WCaOR+ECbSwRUe+VHhIY0WOGHMqwNkM9NfPb5z
7cS8XZ847FtOcN98WoDLExAizcoFwyQyZ9oOnCkWKfhm5pfCfE+JQXdre0O8
TszgL9gMxfuHGdE+ZWqUP4AaX2+dfz/j6HlcSmAPhbHu3LavtT3VFrL1+5Tz
PF1/1UQuzralGIEaynZrJleG6xWinrDG6/LMruwU3i5bXo8MNYSlSz+thEkW
62LctMLPKYYJhTorbSuYHc1vfY7ik+QmfGoK3IVo4Jd+PMvrSmRGjgv+Z86N
9z3FBx9g0JGVgL2rW8Z8O2J34Qb9WBOWEVLMSGJpk1q07Vjzb9tiP+jRTZ1n
TOTbWum4Yv7EKLy/8vLyonZC5IU9VI1QpNSQRPPM0gOOzSoXxaV40qEuHnZh
SnQKXfEFDuKTgWwDjgKxko+I5qUtxGaWoinvHUAgrkTOyXSYgI5C3zFWSoHL
EX2rWPPfKwKxi7RQ+oIPNBd+boKjMM1OBSXIyb8Vru+Riw3KS92BXrGbijiC
p1ld5wdzg9br7SwtxAvSOwapIYH+hQFo+zuIgGPcZG+C9SMsyWhfdJcQ9acp
Gr0C21NS1JiGnAApvMEb+HhDwKWyppW9z5/QCIAWVYxqx54H739tm665XCdh
E7kgxEV7FkqmgWP4KAMKgjSqZ3RlwkhusxNf6TfdF9t7LSquRRezwGBBNoOf
pE7/8gfdTSuwlC4UZDYisFEzjsAh6quP5SpO56InLkdPcSWyRZCaPaq1HPV7
WXhsQGjZGb3ZRbAiRbyNCInLuqMnWAzeCXpX2dtS2yQfbbcqEUSV9hjujvpa
nVGf9AjmhkcftJeOBwjlEpWbF/Hx5k5PgleiZ05kbc1dZR65zjGfNGOZfTDi
qf5G1XjofUUkOPy2aUNEm5oOSS68yc9NA2IRKR4vbhC7wACXw1xNrG/Gckoe
fkgt64o/vDXjGlONjS3nX63ubHMUCQZ9TLysZ7vn9vprtUH/+7irnpE4D5co
oKGMQhjfekqfAYROt2eh1pikxJpjBg55vZ68+rZyZY+n0p/r7eEQWQZwqoyG
RiZxvRMCnjN8YBjcEn3z8a3obMJY+cpVTvdnG0UG7+y8uXosjn8I+1zH6VHt
tIWF3AoEtuq93Qy2+dh0j8h8n4ozJFXklWqGWgkmrPrxpTGjIrvvS0wy+PYG
SpyJR4waFZNKm6M5FpyD/c25Cd0XYzpJH6UXFUwTnpyX2CYUj7D+5x0nj8wq
x7l5XUXA6mmg/MnQpRQhMHN9C8hICC4TPM4pfmlpGEU+6Bw8kPLyJRhsnTGC
k9KDhhO3E1Fk2fXp1rswmoOZfdS+PtPHDA9567Qt4q3M3Y+b/FM0+wpQY+rB
qLvwSR28GhIm8qeMRb4j0DR5FMIRFg+rmRmCxUMT7t6+OMj9Fd3A2tCkT1fu
cIeOs5ctSU8PffBHGHGJbMtE7hiR3y490wJ5C1FjRtTbrNOQbgeY0dA5ws+q
C9UNrdjfp8C39bFTJd+Ud0Ws4UfPhxTitNoLqpqRK2o2an96zPyuuuBTpqlu
rXrZ9A+J7hcS98QbQ2HWUvkYYYiXcv7HHj49Xygz9K8KSmxoCT2C4vJ581rK
upnxHyvjhyRN4nTBb2OkThL8VduClUnamOYG1EnvVrBFmyHlY/TWZX0KQMQE
1J88jOVA3eKtTCHktsCUgYmw4BBtWrju7pZeNj1xVZo1YhRjHqD3asBhCrir
WQCDo0cH5+stjLzBcMzzC7qVn6tykYoSO8HrtNfpJM0OBwCjSmvhAT+Wpftn
EzRULHJu/azKgSLGizFr19f408eENU2FQ6dpM8r6iJ98G/h0aubFbn6QR5nK
xtsUh0aMZtXGp3pI9s64+2S9IsZCY1D0YK2C1LEyM+Vg9uSCk634C3oh+pb4
wJ1ngu9tagKtOYMoQy0S9sUPMlhvDvjsW+uMhBm0UkyW5MWxhLbgJVPJGptY
nZTVmVWof9RIspBkBowff4wQy+2nuE+PY4V+ju7O9STqu5T40oYJiF+iPkTv
mkQXqAikFY6h/qwxa0ZiuuE8uonZpgVIeHqpAr/QwkIbWhqLbZT6wqWMkpdE
AjBxlZz+T63XprcEXGXtoMcx6Bj0Zs4hVyLYalShemvPpuuCgSq8Zs+expIy
GI9n/uKSJI2n0ahA3eBG5n7A2rleWrNUtEnvmw1jMLWJ9/lmGbCJwO23Zr0p
TYpZCG9N6cTYmuKiQQY72JYNb23T40OyAoxDGpX+PH8W3OYDe7TX2g8xYAEB
73vpLeCXI7SJZd45ix22MUO7shKEoGsIOwEEZCY2lHBQsK9LaDD4AN04lwXI
gy5QlYnW8riCl3Ses1322eVpCuMnwShx3uZ/QEUJ+cjWRMXkhnYXtwEgro4v
OxNee7qo5GHTkOLPNZErRg7RIOHbzsqTnvFY74Br48vvtJmfapm6/g0DYQtU
hj/cWmK/e/Yzn6axX/oojctKsl6aFcnKNJ2vy6lHkuH3OoxA8X0+QR/9j0hk
40Rj5xbTPoxxfSVHxYAIDJdBjtTWqHuX7FiPXIltXJSo0GInDidvoiNeagkV
upg4FLCP1y7PcUXkvVuwWe4KA8V9I/44rcgU1xa3pVBw7wylyi6jmBNxzdjU
qh6MZjCa39DMxflW/yEuR00w5FMXYWjAyZsHptVaJJ/NADxizoiocsMCwVDj
Zz636AS/z8OEbcujhTYDFfARd3kcHbNSqlP4qkWewlqvbj6QidW/9vb+oD+s
Ml+eT4F2zo9+YdQOx0OI1IKvQuyDc9XvUCCe8qkNgY4ji3ebnkxEI5U3G7Ug
2ngDWN0FZROt+LJA3dWYpZX5DaZaEX85urQvGj96HoNLO8iaJmmWgJarwS8M
g++0poq3Rqro1cizvITgSL8/XPZ4zuURQGiieiIaBshUwCNhlAferpCSltoN
uCHClE7+olrdTzIjhTD5PysG9vXNoqfwVcZfFMayus/AQod8VYsgkC+YWU/u
BS7t+NfKpmrcvx1a+kl6Rc3dGbT+lerdNlfQ9moaxh07TRyWu15KMYImQSMH
OCs0Lfznf3JA7eflpuQKBzPKZwAAMIm2JhKj3yItSC6vybrPAu2ThKGdFtHL
AzsMgLrAmENsN/egCxsBhdU5iKyKjfSN/GIm/YesQmyWuoV0/ga5mwVFX26/
2NgnZ3CG4t7J+75cM4YhP5ia9NdAoaCHGQudtpD7bnf+f794EBWS/dlt+0C5
dRaIN3VHbCMMiXmp0ajqGDxP42nVYiAV6i1hOoJ3xF4108l19Ts6+8VmTfAt
F3ClD54HS4/vt7ZvjM6kZGw6o0eyxigblR1uaDKKH4QmeXNVKRe5g5DIbztk
BotZ7Tq7vCyQ9Jkc9XXKOMrj5z+kwqM71TSTUfL5cPvU4YrYuZwzJCg1Suca
gdeArUCUY2liKVmFnatjHx8+du5MtjkQ0jmjxdsh19PMedLvv8h28QAvpemx
P7iq/s/zzx1eNpNVTdv9HRusOvZenuj8Cfip4be3jFsWwgkwsYMcQiLDBylD
lLNqTqonKbOGKJOm+sw2LRbG4OMwCsRRtzRcxNgz+lFx5ANRzDQPjcUFOqtt
Kf4gCiTNKWRDE2CurMPWgnjzuKGpmIfuOVmduq22uCI1OqQpgVjVtipZQq6w
bjip0z9MB1XvrR4yAkhbDCHyMcatafdzvW6CDlm984nUXT3NejetNG3XF0Tp
ggaLMs1l1v1s9x8UdafTfXyRbyfP3rDw8MJ2rE/I5h60/URkDQggIzSNylWk
YqhHhWhIAlreoimqa5mMbmmjgZGQkrD5WZCHHntHFNAYF9oZbm1pcE4EDB6K
xJVwNzUrBt+t2J4W9MBSbMF5jdeK81wWrGC4I9ih4wv8JlJEM/IDPBZ0ZNJy
YWbyzSm51W/hDAsC+HFDgHhwZB5MHXETQqdAWIqDhW8GpR/CgSHZ/1nZ3M45
KZKoq698IdAmz6nCi8yCqR3M3RYy34ReAH1joAu4gA8ytSz3Eb0RpapTujb2
C5ZpUpRXBP3cFhot0+4d9IDPReM/7jJPbC6hDsFDMv7qNTmmXc9DG2GeSRYm
F39imnanJfVUXHRtI2PhXlZwXXC5AkXxQAUp4gUWY85TTRfYUgWrC3qYCjPT
DoXp/u+GC8h4GTkeUtpRvlk+gTLKm8muKn5Z9VIKWDlw6MzmP/m/fHeP7t2P
GZriiUUZGOtPnVSBzGVXKZloTF9s/ljjBrnGg6OyWVwhzeLQYk4kkLUGHYxC
fWPrpSWY/CJnGxHwWwLgrrAkcACXV1ifCRrnrzz+VgZTDP9vnrnABkXl8RkY
jFK4vm4V6zMb6M8mVBiPqL0t2wVVugVUEs0dUyTFg+HA0fHpu+AAwx0soPbT
h3AnaTJJLcP530StXItoWDIuYl+yXKrU2N2lFq+3mg9/946nsEyXYv2CR9KB
dd/EkiAskzL4lDlpS16u6RlTdkvahgjKI5Lu1PDV6GJLGBe2GvI0VeQnzYCi
/3qa0y/wlj3napuBJTDcCI3R1R5WJpKBvEeuSb/xSzxYZ7e20ofTvQ+TGVQU
D69NKoe8l4dEBkCmdbNV+5IpMFhJgVaTSSQ2IdinKIZPUNGLSFSdgq2LLh+w
W7f31s5SDA5iEfdLThqUMLvqpRwKTj20S3wPszCZATxtCeWgGz8TZqf9t3cn
yCWNG27Cq7OWFkDSg+CcfHCXusHqrpJw954ned/upupNU7FUDH5fLAnATHSe
rrZOcAzNMIzF6DXq0VtTGP71kGoJD3lyyyKT3STLPSWrUTnMi9UHP3uyCz/c
cVj9f+j3vGFGkMjot9+eUSE3mhH1mOnJnaR7ftoQmCocvM8KXbgPpreZJNpn
w0QSZMwOgrrXfIfk4N4vRnIjvxVJw40iwZWDlBdKlZc3HNp5GKVDv0O8Np40
eukaWm6vN/ASAFSkckT6VBVparxgr8srs+JZibBrepyzhEUfJFJHQDAHbaWp
BvUcytmylQ4uSfz6wQNLASXklkWumd1OXJKyabg4gZiziwrkpUGwTUy5+MHZ
ibQEajrtKchEa++5QK4s9SvOW3s/ELwbTlSkDByIMrJYmS5Q98t5iqj7QK0x
HuQR2ObaYa0QK19hNkMc/kR9b1+AwupNVsK99AZtHMPg7+pKxNg4undfSUWD
ismHKINMvQSiD61lc4qw/P/J+pWGydFZ7daAvZpBXT9pNRtqz2cSDXmqqlsR
LD0JBbAkkHvbwdmSRI2S0o3tLloZ6efCReETUx3jf4z9WJT4MUr0ahnAV5PO
19jdFJrnQXXo8Msx4rE67giX0zEb7TtGxWT/hjylhCjvx9anR1nZgmgwMe3A
hyOgI4dmff7KIDinlD1/S2SNJ/WwSXXSoN0JswFV3SZfYO3qxt58i06SdONk
VyvNEVsGVFoOcwJSwoawTIjIL1Ou+0rqDoSiRola1gH5b1ysX6+PCMXBEi9J
KkAXati+gBtVwdnlxo+KCJdTNhQ2MMPQXUbPRcz4/EL9yrMnrRt47Qmk9p9a
UdZGppE0AtE3QYH4RXyKobRLimrlbBWD1zjjv8rwJH+DqwPh8rnspC+V82mb
DO6gS8E3Fc20TvyLEgkR+nXMBEQiCoi+IGmIpaZeVSpPeBl4rznEMyrlrh/y
UdGSF79aPtzOP+B8zq2vtxE3fsvruW6m/ZIsHLZjxU/ggXD7Vnnieo2nlG6U
ElewTirLGsGivuGhbgNl59XQHhsv6jQ2u4jIZsuthf+xiW0UI9brqp4Qiwm3
BtXJxK5c6qZlU9MMw3dDf0um1WvCW2UU200H1JaXRn1Z4f96BXBnhq3BFrBs
q6dNaYj3wZ2ZTMWaY8bURcbmWW7f86zmerMta8962xJwIKuGWdmqR6AIleNd
9pGjhSCiJnQ4ul6bhNhiB+/XRT90gASPbu8kDVVozViINTPQjLTsQIo4Xifw
5vQelif9ZuM5ZXEzU5sQNyMTQx4J+kEeZTir8IdxecOrfJFU5SivuE7KuUU5
qe3bUrmnH5EZPHEJsN3cRrQ5vinAj9Ahi2WQ4QgyXXOBUM/uw62mFbDF4tWP
tHOfU9ZMqUVFfPrlBQk+RzpiD8wcvuUn8M4BAS/S1xm8ijlyFzoViQ6SDVr4
disSL/xZcpN884jeLSK7aReJmXt1rgPgSX/figJ5I+5f+OP1UFzM3Ruy9/NB
45E+NAb3eWamGx/Ry0dNiZK2E4ZbifNcYfn/qi6Y2w2QK/ojFON51Y+O8Qg4
DGvogXfcOGt6GnbEMAgg2CSfD98ojVj08lvNFq6cx2xiEOa+t3f0vJ9gTTnN
e2JxJFuQoF/WDx91/tAm37+VeAhG40hjlBDDj1NGRiwx5treuHYQJUO+TsUI
FxRaiV+M05SAmMcLRAn090/VABmR6bg4UQFDeYE/zWG2j3PzlNerX83pGvLb
GVq8LVaDkNqJNJS5nvOKWW638H8zUCr7vn+otouq5VsBjJMLkF62G5Yrx7YU
aZRVaLjj4nyOfpraYBUEENlUCkdy9GiuH7kG+NEH3raeIvtn6SskWELiZOTK
YWsJyDIZvKYfhVklnMG7tdneAye9lU8N90Clf7/7EHQl/Jy4KU2dSiDmDqJ7
RAQFpooJOw085B0S7My1oroRfxfD5aQSaX1K0T37iHWsRm+dzeDiwBrWUtNG
LJSqySAxEVdklHMitJ0yPLLytD+kg5kaGUuY18Yuvu2zs/sHYciBT75wGDqp
+a0xUeOjTwRArSLMfsq1+k6zrMEdhEF8dT//v0CEPNMML6vHLE75IeNJ7wc7
7+TpJ81tpUc7l18W7i7zhyAToQzAMkYesCGXLPSmjDqHc0/bZX6MfHn6NdDb
/a0G1y496ZNc0XWWqMpR+I/97Fb3euivjR+dvLcEl/Azdkkb6g7tR5cvdOxI
MjL/PY3ptQvJcShCp+Skiuu+wA+/7Ae++ztg5stIaZRVuYAteatqd/CL2ygb
ZUisqfEkfyhyU/4jdKwXKkpLLK31sKrZoVTgt0Nglt9vlZzSAffDmHXhuCMs
nXvs3zK9gyl8659HFcNhtAnLV9n84GK0O6W8CD+naVjJUSKDcaBqXdr7lzXj
+toigZgRbu2c5DxwUR0onhXDd+8C/DB60bgWYaJfo9jjneyu9+6xW25HBMMQ
+DRBHNVK7QEWQEnXkXKT006DMC8WQGni7B6/y17Kwt7Hz6Z1X/7Z9FbE9J79
bpVDqe8TFAAun6ZAf+MyTv46HITnjhWQH9iITU7iGfSy10TqJO4K14UBB0/Y
5RWV/7vJq48RZVk59/CH1B1wFpRH8FP4aqLGTEpJIe1SxuxJTxaJGiepoP7o
2IqNYb6Zt0BhckPMu4rW6ms5P0CVuqwtEYvhF/L6GoxyoRv3m73cqcbMJ8BZ
YInrfylKS5iY9RkphlsBRlGR2quhf2kDBwLANHd6cOHmoqtTQNC5cSuG3qo3
mBobVCSGXgACZp+ahbXLxo4lKNbizwKa7TAPz102+A/AUomveXMN3LWGSuRj
Avrn3sLyrfuPNoyUAA8q5JtU+uIQH7z9DugUdgC9UhlMGdYnCHsLYN4GM+DF
p/046nMDej+kijtt6AKYo8QAs0iinnoLFWaOiebI5C6vp0Si/+IvO2F/dJsO
yEtX+UyXBDQ3bcDkGcLS/njIVb/6XGk4hFfOsOVKjQhpdeyfnGIzOK9w+VLp
Aq+mMpQHceArDCnX1YfLbInucZYijsQ+lERx0yuSXFtvlla4y15BYJ1/SORu
AZR62l1peEbwhcIk9eYKAa1kW6+gJ/qhAnEbOzOOUG97XnK195mUJvHsKNV9
eOOf48nv+klFKq8YnBtxkKQeF0MdLn9lK65l77q1J8P8WzOiUxMLMZ+hFJ0/
HGyyQCDCM3CnW6L4KA8B1ICQfRTjPJ/OV3VkbU6gNyz+G5E+JDtslrpqW+tq
bmwd4TKBJleQD46RaNfuGRk/g5KUTsldiOZGMGS3gWiJq97/n4l4MsyzG2xH
X8n4upIbrozDZCOezPCoB5B/iSkXYCFXoFqHGAubin37hzuW2+SAvAZisoKl
MdnWhP+wqvO/fr+tucpqtWGG/CIXtjza64NpszMMB0XQm24C0ghz73eYMyHd
U7bxX/G7GhhYzwQFKlnR0mFj9ARhcO9ojYg9MT0evJZ0qIhQOYRMs+w9/gVx
tO1vKfmxCyggaQpM7TTFfwEu17K+4AQLPWrzvXH4pIKUaw0tcWRe7KGeIUGp
AANofYU6L7+qG3s/VnRlNafsaKMlGcCDeoSmjcZGNN13w4/d6hXqQoTpNtQx
ktbi8uZ4JR9Xyc56rxsT/Ot73bAVlDePY5irMut2vpRb2Hmw+uITWt0afhLx
Wb11Fr4LpI0WiuEE+R2jzSLAcBRYbLAjPmSelLYj2aJZ1DTz5An3ko7lihTC
lzoGQWx1EyPV1WSu3dKgJsrCfyfIvglGiJgo05GIBbCXBFRAaQKFRoexwtbl
vtL5HBxrEosWNk9A0JEek/b8gX7S1Mtr9PCb1nxo4pBu2IEcK0tzQN5IIZEx
5fdm7AjlrWgC9TlbXYTLAk6n7JOoNVX+Bzsy+0MDdqqz7ZQZGmdmBE5YZhZ1
vvWVs8hTY1z/KiUR65X/RKuzWrfhehcNL2Pvu4HTMdTcxC7Xd36ZaJWgWa1D
/JZaS03fAicdDThwn5o8LEaFYufyq5edv4tyWZ5ailmj3dQx9B2J6vM+pBER
x9GGCGsJiUKiTl5ew70HChWH5OjsCTk3QqWDup58yzlqVQyythySHjnobXFw
QTD2s4zogtGsj9uwo1D6t5D5bdk5juMg9gQ5+jzFJhibrwxKFaVkCt6BnvxZ
14MHuj5kuxJerQzKfSSA2tkmdCxs/bXI1XWk2DxhOgzX5zsUapTA5VuELlFH
i6oF5tm6dbuNQhDlxjgNKD8mfkeOflrHdpjAXVz/HxJnJxN0upCZFYUcRuJS
8rVx4JSSWkUcowASJJRCKizyH7jhtnC8vcGDjz0wR58SghY7+BMY7qfigOVC
YifvtBIuxDU8TzPxJ4hy/XoBi5N9jR3p3Gv+PCN5ENjw4xIjBwmVqGHHETnU
+wg1qDzd++x6rd5pdbXZ1vMlbXQytOgOwfhSHm3RsHDJchYYGJwCRioiIVte
RrcZWEAnupf3Ku4wTY5HgzHwZ069umFjdrynL5JPuXbxPn+rFGH6WMaxKaBM
7EuwIIqDK+6kcrmHastJPcO9R0+H04i/Ops/aajr/NleDWi4dxASTtMAK5P/
LN8PeMtycfhTe4edH2LMfljLGD4FSPhTc3kOeysEB1uFA1ZED62ik8yK/J7C
23SaDKJjgdL+2qiajpwsjERt8l/Om9FXThxbczduAvtB+rQ1YIEGG2yX7Cfo
hzSp4GL/fmOQmM8C9SyfCLX1KgzRNFGbH35k1vbvxAV3zL3MpaoXGT9WPrIr
RI3KT2OQ4PqrWAFfcuRjFyI3tUtLA+98P6w/sxf+7ttaRkRFvFUNQKDJMA7E
DcIhYYwwB6r9ReTAYqDC1iy5g2crg953CrLBrNbGvOkx6U1Zi8As7Fx783Jf
Wy1fQKNI7Qwa/EMEDZLdootLTOqvaDAtF6vI+N+jdQDZ2cHHUhjiujXitxUu
lT7wrqCu+n5yNxAsrr95iDzDFM8Oi6X7XIXLLQWlq0c2tUhdn4Z55ArNthQ3
d3PUKANRrp+ph9IpF9cDpBEqPwhcQ3qtPk/S5OrxikvcLgNxrho9ds1zVGka
cYkSd7hBxENZhOppZ1qaAQ2pwIxMfNEzcT7X16m4IJGCNEpDjktpgX8iV1Wm
uhBjlLWpKh4jLsJd24s0NsdIqD0kBpvRfpsG3SdeBSsTtHUAfD5p+VVwMsmM
Pg7iIxMtXnE6MTuCvCc/+p8JGJTYvOrcLavZ1X2soRdKtzdIHDVA5Tajzra4
8qZZqvkPdlDcgbNPxNOfz/jaqw9Efj643Ht4X+EiMqCFlwTSHmP3rWUDxF29
nvFeuH4En2cu4v3hZnRMLPARHfj5EF3wIg+Ivoct2zOSvG8k/iexTCNgZHFn
XTUFGQ+/beVxSF2YzRF777kYBMLn7poSMsM2yz+VQNxXkxvynpkcyIjgjec7
Fb3k4bs2zGnPdOhQjLgq6Y/ktKFSZa9xQbZb4dK2Qg240Td/7uKdQe0lvDAl
r7t0oSmCRhTfTy82gPtMN5T6V71GjqGVX8HZ/FMbFcGKm0rRCu7VnHFNb7iB
xQxIrxTKlqx+uRz79xlIeyl1gjuFCEbco9M4nG7SNNpxTXdoLAcSPwBxikTh
AcDjMAdGCXVbqdT7TlPuwqq1adHf6CgyXxzleRHuzdvIKShuLghqbJpV/7/7
UZcQ23H+TLirD2jUcwH9mUacv2OwiFyEP2on8NU8KgiOPvJ0rA3mUrYm1AVl
RY8RpF1hy2cT+dkr4dfJRKSOSqX+sxKQmV0scRbIGoKr6jtgLzmkZV/Q8VJZ
rkoxgKyPBnrUYuEnoAtUNqdqYjY5lqefgT8hV3XFL+YQPtbShjZ7cRAZHHcS
ZvMvwcPVnhPUVI1dIAZwoD2+JyTOqV3sJyhRMwm7tiDEnWtd1i/T6gkFLmYv
A/QBmqJevBqXiV3wyyk5IN66FjBpt7AinpPEJ2+F1kbvh3nNAVTIXO8x3VK/
xLsgOqfRAgMjO9tJr0HzvsIm+CnskykNBIAMlntb1D7+knaSI5HZ460f0Qfx
WcdXuyq7l0qbqs1PGhwTfQB2hhHe8r2P+d8zTJDFqkcjzO70LE9tuboOfgiM
p3XbG1+SOW3RpHf6skONnZxWYkM15sEJVuSw/ybFJ3pWV/g1lOcTKa/wckQx
gRz2vjVH8aILM5n8PGfOk+PxA9JidMeyU6nAY0sjKDx6skQJ2jGFG6H6wJ3K
UorbrKhNkIsfAnOqcKFVI23TflxmuZ5Bn6p4MEjZb6JwDMnyF1uLDaXIOmuJ
UhB9HmlGglXa00FNSWFdF/2lRxjXlAWcaZ26U0QUilGbhznZC3KOyN2qiyLz
GrOCbwkroCFxSPKXKZeWPocEHt3Gx86KYqPODLZKq5Bt/+C+W6XOqZelDKxG
uwd6JA0RSiC2wEgJrGrIVD4uEnQDiVmdJe7+FBjo3NShYT9smjTt/m602u45
W/67wxwIruHr8X+gvQ73MPKokyIDlOmusOjqaaJ6mn+zJ8fbm1EXAuDWo5hl
NQtaGJ8a/er0odNWqNFqujHKQBVsznumoS7Olw/SBLHTT1Ge8SZeLbsts0ad
b/ytBPIidTjtA+cK4uoV8D1PpldHBOApE3aoXjdhUwNaz7hlkunhuzboep5P
yd7efgzskBY+Ajht2EtrBzs+nBi7Io2XysNka/RJtzitN4H4Q12yDM++0LS/
ieOrN3PXT2GC7DkA960GKVuMRNasMVP4s2lWYbZ//rk4CkifkXz4WxSX8pID
D+nwy2qiutWNC4HKy24dvCtVFUIHVHhZX6XDIWuJAXMb6FNGtLJlRDsc9fhK
FE3mHhwQNELyJjS2Pv9zOdZfl9BH79aXJ1mFzQ+3QXL6G2Kc0uO7WP/J31Pv
RjopiYyiRGCkvQeDUHSCk9dt1YlXXAb48seTLEsEfYcBFWwKZUKRML3zauir
qWbvDT1qYZF7mXW3K31zN7SiHlw95nqwXbq7DLeLy/Ix9pR7m1RNNOroZM8B
A+xClulv61CNUm2lF7JrqC257Hf7pJfgG0sFtdDB2mA8mQ6W2vzzHA9hERMx
QE1VcEZVOS6yCmAN3OUksaMcTZtD14Kbdd1BosqKtChwziNHBwnEjew+k/hb
wnFKoII+AjIsQKc8R2UcwXBmwW6ON34MJZTm2ny0EHYGQfp9dTHLtHtRaeZY
kIXDywKjBTNOf1c2AeqRwSUdqTtXHCMq2n2Eu2wf4+/y/k5kO9DFH6KvD9hz
3cSdwu3Rfz1wCKgDBR6awogE7Zh01eU+uERhdrF2xh2NNtPv2MHNyR+zNlAr
VLtLZ2Io4JJZtvR9++UqO99l3RQ5vBJkjoB1VK6XSA7SdMktsbPSQRnBnTt/
ALzHGFXEiyE4aXa7ZUrKHfYtNiJaQ0nI+JkniI6luhcLJ8Xsw9HXuRiC+KIw
soqZOyeJEBnraTYS01QomXBMrheqn1pXS69SVi6F4lpy/jmjZnm0PSRPaDZw
l98Enc5LPOoh9MC4+7udyQlLgOfl72pJZj7556H/THqp/X3ynL4fPSSybRkO
TXjDd8YiZg+3gfGn3l48S95es14Da0HUQeTVPUZijsjfjMFZN3m3G6qReZmD
VZ1xFFGxYkH93tKJ6n1Z7NNEhlYEBfIIRzmchV3NXlb7gDt5u67+sUgah+yf
IOWePIRLesM2We6atAaSblN1r/z4oKQpnpKbb2MofG97xamH1Ykzd69BON+Q
8KZEP7U+QHRTqWfmBf916OT82NRyVWbxHzCNR1iVGUQ+fAAhCMo5QGG8boK8
QEVAX7Hpmz2ABqtAA1pQ6VV1HjP7JUTeE9RTlyW/t9uQOdJPszaAjt/ytGeL
VoYxCrh2kvad0uY8QrEKCh0kYIVXv6oZVAS1U3jkaQhS0c0wPCkKXcekxFPh
RSj1DgbroKHTqaq3Ui47c+6hu180V17pjTR1v3f0iM4YDy7d7sxU6PcnL7mD
FPSewfH69GGqTvX7Us5cpj9Re+5ZZ1ywblcI6KfcHxbc6dd92sxRwjWzpNLx
WPMFMsV/IApxqZ3Cu6dTf80JXn95qSgxvMXFUVdP15r1DvtlhNgzL5rRj8st
h+16By02cjG/XvewJnLJedHu9mglFB77l3VShbEornxgzIkw85UvMu9G1flt
zaeI3PeZsV5oFBdVls/2y/9OD7ioYzdkJ/7Qg2go6Etn8daA3YKpORr+TUxL
5aSNstvGWEQGAP9svU31FK03JfI0rmUo80SiIFSm2mfaBnjNb4WbNFVuBN5z
MuljWHvFQZGZzRpyQN00yP3hn2oABSMkEcg/D6AxFdpTmLFTMIEDrIRhdkZE
7KUtlFEVM7FuVTsavqC7zNxD8B9CPfM+q2mKfamNOmJg4qCQCRVdn5/I2cYI
PgsbEZHPn5KH3OwGR9/Ehims2mrHuo/z7E5oLzt5Q+MsIn2pL8Ulf0CvyWDj
EHWSEk5Evp+AsgljuhKyrO2783sW1a4r00FZ+hYjh3mxATZFvftONwLR2ZPR
dUF6uAIkWXd/tYUBHY3HfxX9aPDUSMVDMV0TmxmuLCy6F11fu+3B08UjSDLf
uAOdPdm2cup8Awy2laXAxPi7l+rd0nwtcFLWFXUBZ5/bBEoyBf/Jl1FE1/2r
748LQcYp0QbJ8zYRPW8pzPbfHDFLBGdzT0q2N76tFn3Zl0AeFLIo76mT3tQQ
PSmsZQh5RHdgNDFafOTL8p/c+3fSV/BCghxqJpGMasN70AHo4sUf90dzIT/W
hSUK9t0pnU4nTyzMWPy9gQlx6wongPyzyE2k/pdT3l4F7Nx0oSi1SyhKsJdV
tt8+bOcsnV19Z+WLgRrDLWzIzonyoESBX5BqHTcnNgrc2z+NT3nl1iIEm/4E
+CGfcMAnARhXn9eCh6CIn6JixhuDstb3anNwCgxHYiWiRXyV+ogGnIFPkke2
B+0+o+6brtfZxy289jaauNEqThX50e6maSXCcAkrotzJLeMQmcEQqr+TupCZ
Y85kLCGngQEgHtrqSjybU80gLZEi3zs3uawqoN3VwSLdCJ8VvGdvIeFxaPWf
irk8N2MsdAjCfm5z+MYrdk/UpWO9MejHifH/sGml0+aRd+sVUclDoKQUbuPW
rOweh77CNoupqk+srXqWPyaBtONXyLpufMXbQaWQu4PRez/BKX4ieFN5idL/
2lIUNb7VuiMWFXFZJ5EHtPT5DLpjtkCKB25Z9o9sgE9SNWtsEe/jz2udGUFx
9HtoPqpvGr0NpWfcOfumS+/KUPpH3AMcG1WhPLRIxi9K827lbXYBmHw9y38L
y3aeFWbxzExgSJSyx3/yoC3ySpLdEb9WYJLh9wMALfrXn2Pl9hOtWFhv9nQu
fbdiWV3VZLCIWm15IpwZOnc9fxoUsyLmiXP7CD9HXGxeE3fbgWsdd0euzHeE
04xG6j64c1y4ifwli70P7RxPR4aVO8D2wKqNPdrZrSuu9WnWPAOairZ7hHpM
XvRDsphofqtpTfayPzCIg1Grk2QYzBA5Fgud0j9fuZGzssEv1dcfYCackOfc
tRKg41yCFlo=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpegM8/Fhn7yYYrpu4vpNQGXc5xjfIKDSaUXdBK3Bn0rv/Xd+9YtyRUG8e6nrm4xEkk5p0gmCo3rH/498HFllij5ZaG49cIx5lqDj8zje/ZbQHhRnTS+sYbSlPXPxW3hH5rGouNE3ALaC/p9fw4Qk+y6JwD1KiU5Peg3jpD7GFeolBANR3jCKEkIAbJUUz2+T/e8WNO2UYi3pq3lZsow3Isni4AIEOPKB8DYpEW9XaLHnG1/ruWrQJ7O09ofTOSFX+3JVJawzBbGOYGl6xvxfS//kmbelpvtSSWQksri6R/5nW82QTePzNv94n6Co3Hz5XHmyADd4a/IoQXsbvdAFRh7x2BsG4b767OH/QE/RokCa1CwUaJK9pdradEPYQ/qkyA0/wQgXOxBqoCn1+tC5pPu2jjBdEITkqVgV1d8A2alBUfEHWCgn6Jxi+r0i0M/ekRQhNR13iQrJhMJwdB59XObO2JlAmuuwO+t3jKPYn1tfdNaRi6q3B7oIEldvHYsReSbbBkgqv9Tvz7Wfr+M3r6L+jcWygiIjkHX3SAsRdnZPsQax3Skm5cj0SutoNoo/l7vV0CM0LeBMLDMJhEK0fyV8BHsHEmqWV6G6/0BxE89Xo8Xwecd05cQ11ODaKi44GC1rIW3snQPKJQ9iXlDx8IuVIUe6SkVyeioF8ci/B3cnVosHv6Q0xIuKRRKESU28k4tmB0xkFdSVDtvFr1Yz7mYeInj30/rX9PuTVysAGOixi0ZYWKtfqiMTOU/pJ7SDPslLo44XoqLrO+N2TcW6MSBX"
`endif