// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
opkmcxzRHLNac7Mt3nOuDuJmH8TJQhHv+R0KNu+fQ9DcKZw3tkyNYNbpc+Cm
yAxqmX6MNMQDIT7SqzDaptQ+1Rnl4DTisjgXN/1vP/O0ku4fyz9QoOf0qsQ7
/NemSK4v06CHQo6F3p/28A6jHvvW9Z+Hw+vCSheUtArhA64MgwpfT92iTTQp
EFUq2JjFrgzfRRS6J+cCJUXMIBe3oCAnRKNuIsXzo32dc+o8kSCG97RH0Dxp
rq5rFWcq7a7XSuYUVsBO6Hu9UuutPTbJIF1gWByIrNKT9k2s/zQoOkc+0rJE
yoZeOYTA5J0iDI1yiuFeuvVdkV4zDVVE76FghvXmlg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FQ5xnt2ViqontaxS5sHjDsp9p9HDoeMXb65V3LU4Wyk2h9GFP72XaNH/TrPQ
8FJFgr4zAV+6kjKBCYPTGqekq6qXFNE0SXAAxUdcdKBFyoTTK0p9ZhfAKvtE
aHHfxJFz/2Gpabb3vRS/Xuzd6VDHnqwl7dK4e25OyfHJrCMPpstZbuBn/WRa
PjVsxrTqiwWY/JIwDKYkILTwARSAUAqsr11/h8eHXoxfsHfamN9LCuiLSOK9
DCc2OieGrOtu3yjz/4dnhGdzsNi37F8fkocbyIku/bHPk6/ZUaSEAo31IZx6
XuzimZ489Xwwf0I8UB8wS2xqTyu0+7y9V06tU/dtGQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NVoQdpyhcqSvacNITZ674RQkzm+GEGa/Q1W+koUeEQGfFMKn1eKDQ5/7E2Hg
fnNrgQ2nTEZ21tg0BA4PxIXrBf0H2WA51egN3jeHwx7DF2iFIGIxAEceYL63
qt39L+YDK1ryy9TO0TLBtqib1qX8vqd7m7IQ4YXleFUtcsAlK7fTFyCcbkF2
xlAti1SvtsLdBiIvFvKfqN9+cBSTJLq4nAIkXSphVE9Zcjz4SZ16d1AxKvK0
xcWOw4jRhr9sSChQUhiWvDc7hiKo6/0DsGZ1+9vuA0ulubrtf529lcMAdBN0
Nme83IJWMAH+ERymiYlLLUTL6Q6wT2k8dkhOOJHclQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
USdILXfnMJh3DC8AHk0ASmOImfQ8dNO9TufkO+USH+DCrNUAVlOGAWA4IxCF
OrR3yeWuYWo9ScqqZswoDpnCoYz6QYqFf8HAyGZdjW+tojf/+VxLZotkEl9n
XhjLfK/wb/ZPN9DTNBbsysHtW7bEdgtB/a0IYkNUS+v0l4RZjlDafZqDZ1e3
rYGiV8YqCRG/PevPGpomRGqnMuKno3YFJBf1RR8Yog8dO8ynKwOFtIYoNXm/
tAxJUsOxEMFPnrOdqH/gPydS9/DncHd9CeTOM24PN8HBCLL8u+wFoFL5k3op
qkoKUkAe3eZSJ7UBHDroco6Q2wuEPKztertQDgccHg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TeBCq4IPetUintoy5kToKoouebuavripd/Go4A8MeWASwZNmfCpnweBANEpG
dkTiWtMlFoc5k3ufTwjH1QIGKF/CNOHnoyUGiBcQ0TiaL8feMD8KWJmc8VtN
iVNEYdzKJejSQttAbrmBQkEG9kcnb+sfJSWTnZ5jpCLLq50kSvo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ksQsiqCahf6JnyJ3mQk68cOUIhownedIHAh7m61Y/P783q0lUrXm0tW6IopI
EjjRMGURfa+B6ltaRq44DYgTb49ZuXvEf/snxj9UGWgZkb4ty42i3fawyRPn
RwpeAmJ4ymM1TwevU0b3JZsbaYaE4u+QrvnB1P/n8TVfcMcSpkrGMOloPklQ
VJp377yfE8uITjoR/iToTbFm9XKlU8rltkmODxln4DX2cUKPqDFBxRApmtMm
Hs6FeaHN0Za1yND3Vp/CVl3xESCwfS8QBDb4upYj13G1O0UcSlJpZo0HKwcx
hUa5In8kMRJQRoQoFfIDj+ILWlSm6QPNT+ZTOYpSPerUmv9X6Dk7kumdr8QL
/W75gHwKiWPOVXvY6fplw3YVcjfewQI3jy9toTXfl24jl1p0P4ZMvyIKymX3
E7ZH1IMkt0mwhS4L4N6ryNQ9lWhoMeVaoXXgmOY4qfQzhq3r5va3uFw0fUfP
JfFGGGPrHZCg7DDB3xKjMPZ8vtQwrdfN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j4EIAYn5BYEtSNqHF82xkOscSF8L/AuYf1w3b359cQxX2xKabSe9zErrRvg6
yhCoN7SUBW1ruPrHgREVcGy0n3KoaFaO4xg9aqtHS4VDUuZVfwt6ERhgklNC
CATC7FwGy1uI4PDuTYbwdiKYDnD/Mnpw610Sgd3aS1UGyQmLIdU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Vs+VmV0XuEq1aqaVdenpT/J4+fN/vaxxSpsHlZFwiObOyeF+Q1Zyh5K2zDbW
m2pJAfqfXNAuD8nVgLpDOUg0zioKQYF6/N0d397Y1xym4SOhneHIc8cMx9sA
is3hfL83ZeLc5Ev571sz9mfVP80gcTKUi89FSnWcEg6nZ9D+aD0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37104)
`pragma protect data_block
X9hi4LbJpWCYDe9GonbJxmx0zv2VU5lc+aMt3koyOHNWfxiYjwwLfrqmEigR
QuH+GXV3sAQyP3MTsHBvrDrjGoWtjIvmEIfG0erwIOCJNXa99S/Fc6PaIbhA
e9IIm8PNBMbTNGYRobhnEoUHGU5U364yhnnsciET3y7Wycdb+968CHORcKz9
QgTrwcm0/SByKAsv68QPlGlQyxgBRbW6+Z6B9nrpLr2k4GEb7eaKn/AaLHop
bVR/W6nUTP61PCUq8QEyck5+Q3IyHr8rQl88+Wga7SolEtnigJTi7tz5e8yK
lWvAJk/wikvs2KMP++4XTQJML4hA5T4+FqHSteJH0jPVXgps6IJUaogOwvnx
5q59I6+Evg9GiY7FO52dScybO30vP8NBvj38IVIiC6YthfLWIPNNLwQJOWmg
qNQSibzFJcJubnW+xE7CxPh/UUe5OBdQf+aMvFXY8yP8L4Tc6XprkLNH2fEA
ghmlYZDlcs+QrLXmVfkO8rnGuM5k9dHRUeiaISrxxLEFDUOq2WUocooZR6B/
IMeK5OQ/wmxCT6bZQBXS1JC1FZ6oJZc2pMuJwSGjZTOXwwkyVKdjGyUSJN3Y
19QokNhuD2HaK4bo7aF3StDFnEKVdSOZqam8je7RIVQJhsGaIX7cNd2C197M
02tnvVo9qjmXxZGKmbHcG8RtWzALDx+Rv2m5bynm1zGaaelaBgRt39zPA3Bm
PFydMCxALAX/4PJonuZ1HN50YkNL1OJu69hPWxhxcYLULiLC1U1Y1+Udmh51
TGjcqG50STxEpdIoMHsUEKSxJszofiK+4uEM3ZZCJ2kdTJP5FplglHzDnNGZ
3C6UEXeinrQ7rBt91nH++Nhwu0fOmknk9Dp8eRR/jIsGWn2i73R4Q6d1pO9F
15tCdJRhiNXUkGQz5pdvLZFqZGFRgD3w0jdHoNY2u8BpB9GOg77u6Hy28dAg
mhGBEdqsZgIYNbrLNu3VloGVvV0+txZ6hvTbzjSkMPfxkzHfhXf7SkoHoLBY
5jRZzNhbE4VrYipXcrh/+tkl0XY36k4a1ZoCyWT318HaUWr6pwXWoUHq/vsJ
Xw0ieG25XD5zeMmL0X6EdOz8s7yM1sqEkihq9GmTQTBDYnnYgz07qI3Q04zm
D+cMCykalsezWX8YFK5haIEBiK1HmBpTlHZh6hxWi3006l++UZOmdpOIfsch
z10Ldl7V/E4IoD1MMqK7R/YfOULlwhjEgxhq0fnqTD5MDalY7uARkzJPUsjB
p6vgrwvU+IrY6Aaj/dmq3kuLfUUqOdYasD7nXLrIAUoR2gYqDjrJoqIDHoF2
uk+dsbB5Z33m6T98c0/szQFV4L2usjUwNLcE9SsbpZXHZLtdzo0qSwDWphAE
eWiBkh/E6GjIywUsAltd1NdCCwR1tnGyHRat7xkHtHthcWNGx3X0KG6Sm0WT
sDwsyj3Z8LvfKFeu+v6Uva3VV5VtDalH2a9jkrhiC8GeneF47ZAZXq7PCiB4
XMCNNkBmpTpDIn7TGfrdUghl5zmbyL+lLXTH92O46+wC7k+Dr0z6mqFRLmAw
8pA4RwzCdLsk0WKST7xZt7W900ANoX3Tr8C2rQzgmN9qXFKMmAqqdPWCKTa5
drBvAi+3MnPMh7gYKnVZVdu/holXgxgWvA/h/egD3SKg8RsX12B92dxLRzkX
do154Z0BN2rjsbaV4o/VyH8vYp2efnXbiFKH2P/aQSUEWkEEXrK0nbwrJFga
KHsMiegdlxFEdzDA53adNJ3SEyuMT765BzaMQWpgDpwJNNe0cCBuZtr9gM3U
TdS0G6UlZPGmHg6WfLhxwsS92rF/43Jl2Hny5Fxq6nK7q+6XVnJGyt4EB89k
nDcs5r5OM6aSH7sfoFWf104hn+uX3m+rJbTsVJkC4mgCfvzOZprMCcTo3tK3
bd+MBU6jwiyS9PVDQ1p1+5W0raehxCZHza1JaUUr0qxJwc4wBMjKwMyJrKrl
S1vakH9yXp17aUyNx/znWpBJdu0RTuxORxFqyznuAoigkj3BGEYfsrrYw1m5
vrrqVYO5xYoENkrcTNmBrtfd4VhKFQXOzZX0Syf+adRSDBLwpQ7uT/HiufTc
tT703R99i6DmuHNLyKZLaF/dmHRoW2rOlouploc0TfWr+Ulmz7GVBgdc35Ec
6uY4u3EMyzPT5H40HBqMQFmaEgb5Mc4f/sqWB4zZRNVg5ntGUkcik/DiNNbr
LkY2Fy8HWGcleC5F5jpTwNKYuvm2iGmsT91HanCdgbBFelUWqEBhtIqR2dnR
OR1ZV5zR5bTHxSjclZurCTZfTVttTdPVNsbAroxp264xOVRGG4AOF/c/TyMG
o8t85f/vC+A+JZCKRpVtW5f/rSt9bPbNT0xyvPItfoMMOzAaidwpdRejmhza
usmmxm1FN1EI1qcfFB3fb/sdB8waOWaIOnCkfy2uF4Ly5Gx/CK/fa93FBf0L
HigeoI5X3yWwZAfYUf5+ikwfvju0JNMm8OeAUsn6KFjjlfxL+tEhpQFxX5Ux
zxHkKx0wP6RjdQPi3exh5BQyywODO+xOAlQUAygQVRC0i7ArpyFs2OoYWYpw
yf+yiwSrXLkPJvsZ2GRxDvzjNnitQIxz1a/73xgjSimaZ+jfsl2tcECnQ+mO
YShv+xLv6IC2unbzfN1orJBvWihyIV2Vgxye8d3sbsNc6BXdKqS8IZ1eo+h2
4R9oWnjs9Qkx4YAhdKZSUk9Xw9PfHVLFcZ9O9vQ4jSiURnJ+y8mQUg1WKHbA
CIYt6zemDO5AwU9kToybelHybGwkZ44bMf3yJmWj9Pe3U64vQtHzelzCoksK
oTnVN4Qq59KIAMCO/JAnXNZ/ffynRfiJn02iWRIiKxXhNL6BtEpuGYla1QFP
L1LXtvLgfw4Vxiqz5l+WBlRuzkHGm+N3hJWMIvujsT0s5SZfiCeGTeAPJHH0
cZb/kgpE3o145r/jWvpgMF8JsoUdXnzxa+I0a4zhyUHY+NiUS0DjWckBxPbb
OcFRDEvxxn2TAudVi5iRI8mSUVvOHXseBadhibMwI137F2v6eIjhLCIzBPAq
+56g+VzhXg4q1HuCGXZ5ZJ8WmR0yrUowlUfxPPeJHGIcDrldBgVyJ2rJoksJ
q83VX9QsGA66Ujo7d1SI+7fEA/+UCcpggRqPkhQOCeJNP9uvEYKUXiEx7gXc
YmrHYkpUpkE1CdELIMjUTJ4RC/FsxH7S/DS013RrrvDptUuAf4Wca9NbvO6K
zeQjGe+ZTpaqYbiDBMf/5BKrIy7beK//tyuFxLCN1hDJ+9HEyZYfMcwVsd5S
56hmCx6n4r97iihMvCkFqeImgchrlaSzjEr//repLS4Lc03ybs+iEtQR3HI7
a4MaaCQoHGZD56CXNWPD/FBfRMHRZO5clj1wnQujEJuWzjvREDvShaHHrtf1
sasQQZ+pgJh1v0eU7sodf9FN9MkslC5FCEEDzyaITuKrETTVnKfhlQ4rsJJZ
dTByfgUzze10rSSb3o+L1/4iyRRX29RE26SUCxzPsFaK/2LyoGvQWd52sik2
0isWPZlRXRLwIQnw8bYGFJH8enYsQ8C43rnI4ncZ+RQMJTU5hLReKKbfZ6Z+
RivaMbgHNER6OzjwLeekzLEGZPqFRXfzROxM03M+hLS9PHSNsvAbWpA3j2X3
ewIVUZXXlYHSIMR1APsfRks0PDPUwG8SRwUb3pQVb+VYJ2r8EiRlRdTk14TW
y7hKgIdJr18JfU3KLlzTwKS/D+0ddlRiaNkxBtYXiogFM7KTnpKfKdkgxesU
SMdLWYoGChtbsEFus17GcflpDLM2NXYGJFs/4UzPfE9rP3z+e4gzgTd/XRJF
6Qyr2GWL9oOFzF0L+8/3vSRRI0gjAyftXIQc3KWvvBhYEra62cjPfFShHq3n
oqvAqmmg/nwsDPX6oV/k21KW7tc/slW644WP/l1nPfoIfLVlmGKRbEuJn6Wx
e1qJUAcKLIFFfWOQ/P7iI7hEiOBJuAxDhIS//kUZH0Rx0GufhCBzy3Jx/BbH
aOAJwM5PtYDZGiXRWMppHfgbVTHRvlvUGZKTb7/S0bQONOE2WbbeKWwAHRLs
PcgIAyeVTniS0ZfIGmOM4m8cjHx+lrs6S95j4xgiP+UBcWTpl4hpvLbIAVTB
InsssVMiRnqvOEff1rE76T5PKxqWgNO/ekK4tQpJFVXe9r6N/hlhRVhzdYtQ
sIvC5t/HHqMMaunYajnMaCeHBO78nVuTEWetyfKsb09Bmnxl8NjMak1Y3VAZ
g8p1EBQnscCxHq0QwnUMKiLw1cHPwaEzNZEyXx3ti3lPJbiPhmPD/2SWHAkT
I8L9nB25R0HhSdcxswk/XyeEXFv/nK0FeKjNhYJ2vg0PXxhEnR9oeI8Wcy7w
/SIFFZYaJysiLrGJb51u8ZdKO9P9iT9B6rNW0BTUQe6KI/Kh/iz99KcOK68c
tJwnkZq77EzjHIMAbtZoNd3DuICnKOwZViORZ4HOvQ4eKBjQjrkFCCbDGfSl
O+86uOEEIIlPjNeS+huE1goo69iUOo5yMCIhtsl5Nt/YVBhYb28cwX0WQPDs
mC74lLukfB6f0ZTIa7VzcMbu6SKV77wuH5XcpkK3yEqZGlwIKQmF7OWC+FGD
a7SofeaNJanJgowuLlQrazmz3TtEzU/zBJiLM8mpJ4ybWS0AwqJ+opdUbyP2
5geg4831+hmGljJZw/Otw5cVXK8ZKlJJ+DJQfUV4TFSaaYg9mKuBmDj+qtHU
+VQK3Fc6lXjDE2yUUlzvR3qujJ3J6Hj5fVYaFlPaEnlfJ2Rj8GgOJxFHpx1/
ojQVDPhmOJqIwwwg6t7dk3aatzzsBBdwORUo2jIVDRQEnHIX9fXaxHMxrN3v
1jxQQFRAMEQZ0WXeipVv3g9k2nW9+bBTy6EwI9dbMljAo+6Ni/3NwNahaE0j
thQOwl0bLgS1qjWRjSqtaaYV29M9MFMT7ZDlRXoJSHYNV0r/8uPxIdIJFIwH
Z9FyNS0W6rLtvbTAVTv/4XX6HZgd8DOpdgwMJe3o6ABOSYen3lljNlBl1hD4
YWT+KfZNjCkwcY4XlcrGaovmXubExjlRYVWmf7xnoO99HHP9lso84N8omt7P
cLCv5q9vzL/oM13XKeK/bEeKwBgpRk+OlZKj7brPDxwbRhanpSipbYQlrPET
09N2vR/pJuDG6I3kBZbwc9zC+dXiLgmeGIyzP5l4D63g/vCIhw8TPgaTTkB1
Yxj28Hl87fHQ14OhQxgK5XyD5e1LcZCU6LU0m6r/gW4gVYZXgWLcGh0j9jFg
paei4/0OAA44iUWD5Xp8qRXWp+DE//5dPwkQY4+s/VzBDIg6dkIOEecmAXT2
MG+kZtbNLk4VSwUOwlHP24LIrzrBnsh/vIq377ujzqEiNiaNKVvSExtvmY4q
vjReTNgW+KWQi99q95X//R49Qif0/vbnk2TTKiulas9/2pl7Oz2ycMDviapM
nNhLU03f6x9ws62SXp6ObxqJAjjAHz7YR0oPOsuCwGdDZNWreGqnbd6Tiwrz
BwkMJRa2wshf/dts+8nx7ZHvrgUhM3UTubrLAKNQRQ7QLixSSnzCAgFltIDK
V9/7gzqMkoQiTHV924xbn55J/LvBiieyT1ERBX7jRG/1IPbGOlPlhvLhhM5N
ANveur1rohaBVFVpnRNOM2IwulQldSHCoBUROWiG/YZ2uA6bVgZ7L/P8DXg4
WGvFy76JGJdjyGsLdmPS9L1st2qgwy6Af25vDcNw/qqcpj9Wx/ad5T1XebQW
lV3pX7sa9OqvdiFOfWpxG1t8Uz8ANHQKCdNDoULXXENQIUSr3pt+5t7r542G
9nF/i+uKlcVG39D/RD4rOAih1xz1ta3lI3XG1LSxgpqcDr2i/7c7XCNqa8eP
o921Dyuq9Z4lKde2/1KOK6DSjt+dJ1RJxbdtXFe2NScmeIv9k5tm/RZlYGoO
9Lbooho0nW33Z9WrLv6JIeqVSxohyz7jPdy2yY7170HXCGuRWFeyWC6QzNpo
MM3UU0qnnWxouWenICv3mZ38iIKMRRyT4dtfOdp5lkiFl78hYuR9f20V0Pca
Zu95NV1vI3yjC9hOdj5p0UvFhdjJIKM2dm5H/ZWe4c/8I1B1B0vagfCYOl4E
r3OCO9q/XdPBvdBAv0VHYeOXAAFXKPcfWWFFJXzdPr1/nRPLLlHGWr1deb8E
RcnitEeVugXQjzCfYiF4Gu/UKRVv+EsoP/2GjMs/blm83QnS+1CymKRwcrge
lYc9ODGG1LZF8HmJO/AM96e+be+m456/9Q/eUlnqH8taDaJOKiMic7rWwaUZ
G8/tqvBuk56YCZcuWsbEzLN619h0u8hImj0qW3owD5Oiqoz/zWWyce7kjigE
KVjMp7KP8mfzdrLOe9LJuVk83l8a6CFqf90Px/T/lor0Yj7uoCE0qIg1wzAZ
4ezubFG/RX4jotBO3siAW4bga8RkRVo9S8I4Fl5uaqvL1KSH9ySyMjg26auj
FaELkOzXzNt7ZsWNg6b09MCqG6p6oLd9sdT+AATjEhZY8sstnPtYQaTr+q1b
C3z9/Nyz7Bs/rvYm5nqAeCT6BQMnEWwhxUDPdlTRQq6cFlacEAChnsG4gGPD
+VCdJfAQ9bRcew7qELncqjWumuxl0xeg51DgA9n1Jxt+3E9xNFBlnb+s3g2+
Fn3SUSO6TNmtQTl0b5in6Oa3fReF8p48qvNC31WJanMswinkD4F5R15CTL2d
0jnD67Qjk/YZ0gCG58L4L5zJ7Qqq1t994XzzfgLYj11SGP/5PSF9QKRiA/+w
Gi2wjCpPefZO3lYPGyh5Ds0rBVdimazovVeulaU6C5ACkyv0FE37WR/1d0QO
ejtmF/Dl1xgw9bPvyIhG8FdDfg9slNkHNvACDhYs+pFtbkzLsaw08Rr/b0Ie
132fjOwja+/6Xnxz0eAqyybrlCYfEZckVo/UOqrG+jSpr78RHWm/RSuMHC/w
YPha2BXyTy4zisO3jIsmB/DcJ6erWyNXOcVD4mnuFuhnDEIbnkSU4GgXmM39
/DvjYa6c1tWWljq0GbVXYR0btr5OJGn1S352Gslfd2lHVgCznYQIUmirS9hA
tQl6Yu1fVakjGbjFBILvpov0w5MlffLBMmopzWOhuSCokTnGeuMf7GBWCGfu
rZIpTrkJMLhCfKTP1c4i4sMxONrzMOPGbUyGDtMDCMfWc4Lb+lPHPkOND8xi
e3sl1yIsrkOM+lejGsiNwZY821x64Cw7IFQe5VKbrRgcmhxxbA8l3ncT6hQO
/tnFqRQQ+UxiEdcoUgCjTK9g9ivK1mMUJCS8v0VXNhFWuIUFsEPN8ZE6kw+F
7yZcFtDjBeT8jqZFjLjWFSuxDcRsuPB00PHDUJleVnVBczjsdIk+nDsb6gGM
r/9BG9e+P1GKogjyeuaW3mRW9wrGtR09Sdk+qlbw6X+lFU1edWTmAy3b809y
iZk0Q/3C/0TRiIoxvwgFREN24bM+SDACacr12Vtg5heQLUCH4FSbcBfOL5rO
CRF10cMVufmBVr3NtvjZXFeMap1s8Qbc01mqLsxXGcitKfLeqih/YblpeSVn
bOvLrjq0JPIFViqs9sdBlVx2I7UfGDK5OVUhfa8VGoRh9d4agU3YReOn47Cm
3T2HgIEATzQ1S46Kv2oxpa+br6Bw4drLGMtIcNj2Cbq+kGOtRvU9Zd2WCPHB
lIhdfoBMjQ56ifOIgN5RPnSD7AsPB65LbFcdTLizJjvBeGPCVETYDg14S8la
wfL1r8KH/eeYnocqZamtkuScCn0YmTGSh6MNIs99QB5xeAY9Gui9sDzqLMP6
6RKbyFYn4deEahGSCv7q4pjdLwHYP5XaYO+IxDwtpOki+h10ywARxJTN1i6U
eCUi5y8RzbUL7RlZvxdDv6ITy+jlosthwkRm1snJltuQ21u7teJKpyghNqEY
nXS8wclLItjR/iEjQwKXwoHhJxyaGy9zEPHf+5o9+0dTsAL35FtiORCvJMmM
2iyUQRE+n7XSrBrJ7wkjXj5c8Y/bR6gLrFkN80T6ptoW2h9v1c+Y7eBQ9TYZ
Dk6NL7/ay03MOpcZfBCO2EZT6y9u/rcIPx/klFsQYWafUg8Ek+2exIoAa2ra
2Z4WmisaBuRkOWzNiPL698uhuv7Jh/rk1N69zQtd+CDh48eOCe+t+jbksJ+s
qq8k8iSgA5LUjnxns1gvljCZum220fZxmX06eykKcTcHErE3L9+tjLys2myP
wJmySTNiMyi46NJ/kySn+mvhN43KrkFrpQCEore9XM+2BJLZT7ddwAACVVdv
LiXhBsI0C6lzqrLvfopCJ4GFG/8tpMIz6XACCbx8PEveFx/SDJWUeJS3frE6
4hsdxARJ7kgU076qqj/ZlVHf2owOncRPQ67GO0b6v9DQNAUug4l9RWueI0l/
JI8H1NBME6MtnrElW+IrvnlX/4HR0wlTT+QuzT4xft1oq2XFiN1/V54meVvM
DlZ3YwtSnWYbxftsX0NN0+pTLZdVwyDAneHPCmWdD3crqateTUjiOQdCK+VJ
vlzH41ecAW7MJ93BNyojF3HhfqPnHK/DEHf+IAXJR/rmoLAIkkVX1ZQ/c+8Z
SCX5J+RcwEh0aKCV79AFLmqvHAmop+GmeDQMTOgwuJwG35DxtMm4vqhAsOQT
Xacb79hIG0Uwfz1KK7P9ahPVixXXAR7gguxWk52UC4IwFWJYzSankSaKkf/S
z6vPvHmaSnN8mqP4p8GdGDwvFRCvX4eayVEGfbi3Uw2KXRzI2hnxfTZtcVuf
Zw96GeOQ30Sp/ckaC21RSCQ4KC92EiHCBHpvsIjRmIpmYgh/yI9NMWAo8FK7
AD6Lln5tT6TO+Fp1gpYIIvyaXUztWarCj6RVWkq6MnfWaCDFRQ9i2kr7KjCC
w25g4t+YTORbYdKfdL9IUamKRCqDgUb252lD5n93pccB+29SGjwy5aYVIz+o
jn83qV1gb8NIOqbAE4FKHxuVeBNBsn43Nt34UZe8h2tU3rVHf9tcHFGNW/RT
oPpyLAgU5PH50lzGABQXeDTfo3wJMlBhLayP3bQmPTLMe5NunbsZHbSVER0D
MeHDSnpPFyJBEPWE5KhjMNxu4ZAjmKJKBoxkD8RDfoCg8BKAq/BcIMhcXp3g
Mk2uz+lsCQC2tRPcZtZ9wHXhGMW5YhmSUjgNTbXfkQvY2RbW0HKJm+JvsVHt
OzwwJmVYKYh12FH033eNiXLW+J44FN5j6IkaPK+JRIPkYkAwB836/681ftp9
h6GPekg7VbiYQImxtcEe2HryzDkO+l2S4nmZz8mhw36MtmkE25pUD45kSN+2
w6ne8UA6xk0csDTO4sg4EXlnfwchYD3ResvI+Azu3/bNPA3Ja9UZK6xF3MiV
VxB+6T0E1+jfh1kU5T0jnYmexUcmP5KPVnYefqFkztPXeAj7al9YRkPYrjHz
z9x9pqLR6Pxd2VA1doVLSL+G0GRPeSeDIgnqWeNPeg2HLD1iQ+iMdDClH0Wg
PrnjECOpOB/IkkBKSy9EfmiC/HTddpSZP9O2eee5ynCERURApd94AFL3ONE3
vuw4H1AMcYn//UTUDj2P+XZaOkBdJwwavzPQRMf7OzvN2iwfYIJbLpZBnJ1Z
y0RwSzMSaKDWkkWK30LTKwuPDMmpWfutP0QJ7C8wUHjywyiB9FVzvjSlzpoU
GTn3N0WI29AQK/34FROa7hX345Y/L0YAL1tAu1mLRYpk0413KwGbWnjY1YZL
lpV7CcRPUHgP2nCOP61NBCRZZLsuWCVxYY7LUQF8E/Zd2XXi4FIzsAa0YIky
R/wJg/DaH/JG2TyZtljoojhpWB94dIQBG/H/J3ql5FHhZ/MXWVq3c59BIo8c
s8vvWmNERCWFnuiBkTXEIKfN+xA4R9cC28dlxl5r1KyCKmJ7Pm9waoPOF6sE
w1HPw9WOpzJP9PrN1OVBAjHE2TAe6EjPo0b7TLJ/tMUv/QpOKnxYYw5y/l2m
ai2VnkMVO4dz4Sykb8J+Ekk8HXtSSMnflu7VKxz8/mbNdGlE1GYwDPwBR3cs
ObctWdtHkiWctDa6SADtqU3kPlwFbxhv9+cJ448we03fCxNXyk/H4V9H0sE9
RAJRixrzuqBjIY2lcdr+p6x+AP/Q9kxvAlioavkmTk6sz68zHp8uZ0pSlb/Z
qq1HL5d38Mh9EP1S8+nYgtaqZqRII1Xs2NNoOn1nNhKISdGFllaP222tOkRf
+ogKketw2NOnWQWW1hL81oY4NTzqlNmt3551KNGJC2CHT5QF+IkYR1UErxYh
KKbVvMHHoVg7bGzEO6CBoSL7POmF+OqnF9iuGna2enqdy8eNFcCHauOBuDud
zxrOyojRSzIJ/84dJkObx6EqcnI7Q6xl6NSZqOIPb6S17VGv8q0zryt3Kiuf
0cDa1xiFVHtsR1ZWnymh6IJxmhiHUEshoevZQ9RSUSBpf2RPPdcKjgvk/eq6
SSA/1K0wI/f3mC0syVfBgnno6Jj7ht6aCtKrYXyjfe0GAuBTwHqcoKyoFIPB
bk34yS/t8UURdwAB5UW4BCCNEbM+HZ0P3LJ9V32CmeeNZsHeuaPOdZRUQa7h
OTxnuCXZU/kYpvbwSbxSEcBSkQ3leTAm8kQ3EZ5Tw2amJeTjerQjpiod2VCV
ZwsJB+vLvzWttIF8sz5z3TvbR2/YMk2p58kILDPpBLgm/WdtKZC78oBFg4JT
m703NsKGv4y/vJQ77MXqwigFG+FoBi6v6oJbhjM5lcTLBN35lIjbNAoo9Xjc
fwXZeHQXdgHfyQmCj/9ssK5aCzoa3MBXCGilXp64OMix/jLHfZqPKmNxYJaP
Vkp5zTYCRnneNSg1nv3EO1Mdx5Qx0b16bmCAZOuC5cwYp53o6NFWi4PVlQuy
lqnPWCkK3X4U8EEBM8a6Mo2wxUeCyw0b3JIwHw3Ljk6HvKld4Gb5DOTlmf4E
bDq2+Z0uNpRupFmHJ5oAykJ40c902jr5Sv57JKG4T98jEnQB32w7fcxwb6xa
byIgvVNan2BAZqbBcKg4ePRnr/5E6tb5oWrIauYghcCnRP91/LDAW49Bpgjc
AbzmRYi1ZKozux47aDWEuTuMVsCJrQq9SSlfqVcN493dAG2Yf8wMzVI4jdKQ
rTGHGwjQ0276jHOKsEemRO4tCnpk4ASNmtpBwD0pJmnyU+Cd8+/cfvXx36Rg
P0lWR1igkAI925hH3ht+i9mzwiiP71xzyoZz/MRUTWZl+Yge+nQWP7f/TGuJ
Mb7+sQIcaWNeh+YEEFx6HJxzKRHnNqeZj/VmtY31/6/pDhi1U+Rk0EkphQpi
ACuw5a6AoIJvdpaQ11gEDW5lYYhNVNjlNKltKnYtMycJio6OAnFV5m7xW3XK
WYZZACORu1GkzsqcJS44PlWFfMcfQDmcT/e0rmdGskPNdYJHVo11q9Fj1m2j
vgqVQHT1wmUdwofzhmsCHxqFMRfLpwpbcohuFwryRQMLQpsstz1XKJfWFIIs
z/GbklDF8uHkV/tejlL7kbT4W+W3wSrGvaUI7mgIz7u3TpIbmrzFEk6b3kL7
Lx9qVdfzSDI0vmivdGasQG/cO9/ZBiXQJwsF3xw5zPhxDFPcWHm0ovkJcM6w
D58WBRboakpnoCc6dfK6qnTMRA7w3Uop2XsVNmB67dk7P4D9lPVnAwjL1V1C
glEB7lcmWOncBz3OBTALBG91xrR+3mNJyX3uB++qFILv6d/KyeD6ozkfAfzH
T8V4HGWEhRhas3V5dsjFQG7ULUTAWrBmOKw4QOZxbx4uwfu4871dohl1ptYf
o09K8f2ujoUgBdLuMiH7yq/alMqm+zs8VbHWKE154HWFECPjiH2MxXmRp1OW
W2vyL3V6l4oSbWhGMxZDDjkxKy4M7ty323qsXBI9jC+DwS+Nl/2zdiYrJtVL
qXqnxB6MpLXBC31Hg9kp+y4xbqh7AeQgJCJpLVZCvkVvF7sFEReKX6znG67u
uEeqlSW2eQ+FvuL0lZ4lZ0E0rmJDtX6r43AOvCe5+bQ2gzN/axzK0vtkRbcm
q8tnj7pMhNw+xSJKXLNJp4dRAz8R9Bg1ZBqLhW/zpE4cJ0xalIsf1NHRgu3S
ZENFPYxa1rTlYWQnOWIPMyCXRBT4gMHWxwQnjOpfnISh98Qtckn6paXatagQ
Mhm+r68t20tc5KCuPA1QJye2BFEIfnuD5/o7s41CpCjcnPLupNjwsF4aJP2r
G3af7Kr6OrDmFT/6vdxYvldmt7hRHsaUYMaUFjIcmdg6yWdmorAU99Mw3EDm
keigj70AW/nnkD5O37d54RbtU0loPgWmPz5NZSbuZcmu1tZjOy+JTsZFSrfY
2blVmQ3qYq1XA7PHpEYcg6QhP3dR6z1CgnvgV0DkYRGUzKL0SFWIYPjPxTg5
d7BGRnNvSN9gWhlrS5+FjsYe8WO8nlDUgwDqTDL1GVXXbJGUZiuZqymN4eEG
GHMhK/ea2bqj8SN1TkZsKcSXY3MBNQuKAUKGIDti9NXIYod/cPBmZl75zqfG
To0uuCT15+MgYgNCngNbT3jWdNWS9GaEnE9lPZkldpLugIw+24z8IHYV9eFE
7LCBPKOPCZdpasWCauPXd0fyH6Sx2yBQ4exCA2vpAxOjGgafpQwlnKr+riaj
tWq7G4bA5iJ5oHqO4gUdgRKm45IPEVFQRqfpBl3zVppKvDBFQRy5VYjgBD1I
/2nRj3GHgDQOgG2Hze4W+7lmEm27nuNbfcZSoUSPDXrA/mII6nH+g8f3gtL7
1nKocGWjyeeQ/YWV7cFPaWiCOICXm699B9vKHywyqaux2LkXCw/cWi6qojMr
hWUuJlletMCXm5s4Q6sHoaRNKfq6eBJ/6AXlJUVqTRkIS6iByszhjAPiY5Jh
59fT3HzXVE7CX3CCHggJWwTLo8q8JPObXqv32bZfvphXa206Ueg9+4TmdzRT
hhlATpn3LWOI3bbGCVJHq8tkEM6tM55pOSTVO3/csoA658I+ehH24qtfJh6z
G1x0EsfqvtvdJP5AFZILb9PYlIwghhAXf5T/HH/5Q9xe3wQt1H3acYM82+9W
royOh6yEUWC+Vfs+4ou/DclF1edmGhd4xJEHRYEAtyrg38/p5L5DSTKLkCrJ
t/hEQxifgZQ4Jwjv0u1oN1Us8B91JucNJtaal9dXP8g9FKZzxk89Ovz8bXOK
hrH6duBuNSdfQKO9R3junQZQJfPQ9wdBbOokd5Yfk6N/ViwuEHjAXG+ubQi7
x9T5EVVieT1FvJCDR3vjNUoeA90PskedYmzPQa7yEbWoV2cEX/jO0VSXEoHL
a6z4gv9N3c/Q2qkcg8Jw4wRDs9HVmWIrQq73+ECsV1aWUg7l+6Sc2QqJ2s+S
6n8/7PIOD1KVNNwhSRo75pNuoYTdHT1EBceqL5/C8tZCKqCkO6qSyOG4cgH1
Cyc+qAoleQ0G5kfoggyrhWRhFg68MPvcZTRNXvTmqTw/NFRXFL2rnMyIxjfe
ic2iSjzYM7w5Bc97035zAiwQ5RsHhNbp5ZxyKtRmPJ7rWtkhBAq8TI00/yEk
vTazHN59bS2L2RR/5uvtu1KYB7Td+eCTrs3OIBeMttKcMN+enBYXUe9Aj6Td
/XE9t3+CDM0m+ViKICQGqeG6VRkg6JDpJVAXiliALSEAYDxeiFEG342Usjvj
fUHgBqnA1K2pGrW4iRhOTDKqAwr/RvvKXp1siZdR/RAJaO+c9YaXURiAu9Xs
0Xto1OsegQpP2SG40YWnGQcZqaJdRx8fegGAhtBYfyN7Plab/xNgEqLHc4DK
FvFF0QSnDxAAXqrxtVOR4Q4GiplsCmkG46S/mcLmZrBbU0zuV/uDYJFeka/m
UNavhyxmx3ob31LsFpFaWc2g8rjz8Yr7IXRR9f71lCfKGdEz6KXdxLBHzG1Z
XLu9sXWOhCPTF9YfGFb1djMxv5sqXeLrgyF7x71RsRMLKxJYKxytaPKU9MGI
8xF4bboDXgvIFVF2ga+M851Dx03a8/mxgy3/PFuEzJ+PFQmDzsKc/VYVXGBT
H0LbiUpa+3v7QQZBsgzWQc6AF7RYYLLKeHHOp9ZVMuD5WS4PcD8rv1bqAIP/
cvLvnZm40WpEqmxgWw56egXbesLT6nkdNuwl4EkGiHvxnlr46Z6PyHfvCCov
XRB8u+wfSC7gOOgz5NzqWIaD0iKvpF0uP8iCBou0ZAiRtau0yW2rw2Y2ZByK
w/a09i1g11nZsu0P3izV0p3NhJ9nNTcUE7oP2WCDOV6pMI2N53VG882PuOqF
G78rV1TWvLBq9ARxo+WojfVfPPBihPRVRb1O7tKDozmMuYKI2LkARot9cu5F
gGShRhLPQqJNA/80eWc+IqkXbD1GTFk8AeQ7Lpp/dq79EMuuhXVBQAbbc499
jFO9puXHTTm03WojfG1Pfq2RHiKn3v6bT33DgRiR7p9KWU3/8prstJMHEBcq
HzkFaAV2z+67q3Q7Nz4sQH7qc8IjFT7/kLDabzVdJkC1cw5yi5mdIGisl3+9
LjCaCDjOTKaKIxIMdSQ4Sy7d4+81WxOVS3SYu/oGHDgKt9+VwoGpX2K2nooR
pPPj/rbihWGSeptuOaUAA1IepOkI6zLoO7xU8RJZN6D5MHUXjvCcCuErFtbm
IuabMuCAqOckUBGSBOqAmbU7Mm6QPkylM+YgaVzdZteuWSK+RM/RHT0LLP6R
pfsmR6Hu3LD7SRT8UgtB9dMl1oCe8z83ldBbu9VAC/FlctuaUDTy1Jfq9+gx
6jLwSokNpas25bIYiDdsWzNYM9j1QVS3p2VvsGot1vjufYfPjn85dCnUyj7j
5rkRzNq71Tj01hEGCZtJGh5NXVGlFRhdZW2k49DY0TmSSmBXroGCIDTrX3I+
g7m6qEwkY/CUlPRAePJdo/WVZp00hZKWV+DhRXLV5K5DFbgIkSuYqrNb8DLb
ygXmORZ/ZqmPIBEDIPvn8eUeHQaVxT72iZ4Zbc0lULgnmVkKHHl513WAkwT+
FWwppXtY3gxdy1uQ32ObNjGAQfGKpLtdk59FlkguUYK5mooSuiqQstU92VRW
dczA0h30BfnVetF9mJoD9odPi7x/N6nwPpeVxvdVz+0QGBu3MJolg8lryydJ
fAzz8lzHRdzVbMBJCI75Nr2nxd9oZwEjXZ+aRu9e/yvN11yZGvGHNgjW8QKs
jlT8/gCH7+mXT0B0uyNnX50rKM3JKn1Qp47J0Z6lueiY2PmQvCpl8JtS/9AT
3EuC/WfycUTBXSGjTqL7TQ1nrwLtzsbjyTw4gQfpROWijlP/tX3Fh+8RjZ71
xi5A6TCeL8xsMAOmdSyMglcZpkUItURa2OGpDHVUva/eaKkuQmP3CIDshNg0
FU66vSZNoSnClIgWlHAdNZKil+Zn/7TaFjHgW+oRx6O2z1pi9kG0LvtTbh1O
celQGnmUo/a4RE2MJ0GkFhXRmWZ/Xg/eE04ScY2j3D3KoR4ALx4g6kUcS23C
LglSqGrABSNK8I+xRR7Ydlhjvx3h+XvP8L5ROoiOnkZlcJPx1J1gxwLmMbve
l4y3X1XQKdNjzVdlFl+iF7JOyQhFAJWHezUQjndIcIJsK8uv8N+7htxOp/+v
M+nW0TujoG1Syq6K4vqAHyBz+qAw5FkW5CubBuG/S2EfF7WD0puZIOxg3kt0
DWIzOoZBlFJP1ITP44NbW/C6XgGkEw4ni7WY89PsbB7PeFADkwRLKTLsNaHD
mhhVbfQy2YTPsKNECXFc7fu1YVhFIgojinNVVl4lcYtnp+ZpdA/jL40yntK4
kGYzkgIPdXBKBf2nLZoZTh6Q0EI8j5cDxbGiEXvDS5psWId/xJKNTH5y/9xR
vei4QuuP7+x5DN8K1NKqo7kgbM4/lYaURMS9JZCp/ZD53FLKOW2ZXKmQzyz0
IIhRi3p24kE5oL8e6vnRkFoqqLl911SpGbZ+th6CDVSrDa11YGCaxUQxhO+M
PO8mSvVt96Snk3+bwe7onNZ01CI1c6F2RYVOuTQ7GolKKIDWWqqstBQkmlJz
kLUybo+Ug19WjaB4qD2zfRIHz1P1bVjLPKuaTchY/bt/iDHupuYWi0Q9zWin
yvWVUgWiO+0GgN/JKLVxGDOrAriow5DJXDjBGiSjpHKuoUkdvgS72Hlfmmbi
MfZfSVMJ6WlUnO6ykZX2RCc1EfF7UMST8Q4BUAan6+aF1V5x3T2vR4jsCDVh
jYN3ELXM8BThImOJOhM6CoKsfAMuv0GhkMCHXjz6Hj1n2ZtyjIqcXGEXCgpr
CKJRsRlylf/5OBIHWSjYrtu5mBnANMNa8DGF1iFKtCG/SJhf2yeO+mQhTTsL
ThGdniVVBerXDnWH7jgRw4/F1wo79dYq6aLH/wXQBZ3tBcAAJ3E1qJeOGce1
dAkk1V3GV7oiHmI5iuU7MFRnH8A5js9fS8FCtzUy1CIEGsTL/5qGNGytWOZo
A2oucBBtj8iABeAnpfRi/WAfhzi0WBTzGkkTBJGU4VCh1bhsLgXmyWw2LddA
dwElb16p1tj5LuJ6Jv2UhSkgutpqE1Yunh3jXpfgM+CjV7TmPtUvvOTLNVp1
V+m5GeGu79FKUYnh6XTSvDLDsjjknbBUB64OUBEk4pUmvXMk+0ce9ibc5j9Z
SM9SDfbu4ii33eaoJd33++iHfT4P6tXJEwkW1sfq05rocmelyHqNcq6zsCv7
PGaOgVSEZgUgo0acjOrtAHrKdwP4Yvdqt9RTqJWp1uC+J8WcxVMSXUrKhwFR
ZEx5Msj4cUfrYzDNobMNoY9uX/uZNudvmnlwJAtmr325mFlEoUHNndOT45ho
nLq+mD72j0Su9rHH3VcoTAFetp15G8QcEyAgIMvMN7BNn8o8TWVM2TIVWB/L
N+udC8aMBRy2EoWt0dPiIUa0lfZLSJiYGyy1w+2ulnI04US6ffgAQ5AG7aKP
/LwXLM0+w3jWMJeWeuTAgwL588yGR4ue3BaOn+YwZh5iFuuB2egZ9m6X55PN
di5/+GgBjI3MDyBvpY0BgoY+fSTmQN/pMPJUmALRQwjV/p23CMwh3zZVKMe2
dz4OjVaSqHKJvDPEd4BzUei1pz3XuTATYsoD7lQZWnQBFuRIJl1WnrSrLhHU
GFV2Qs2aFWhB3c7trhKl5aOKOMKM1bkHFIF9td586WRiBqKEa26sfhwWiTAp
Y96osZkPfyf+dCa8k8esQ7xtQWYcC18Q8/1k8ohulEIPaBG7onJ8t52ho5UO
UIEVjDN9ddq7XFPsqZ1M/U4o9ILIbFi0ai9L2M8BO+/katRNQprgUwriRXba
ohUYtgpJ8Gj5Fi1zoyt/IFikIuL3S/zCyH3zAJNYMrppQbKBWIwJmFgXCikR
YUxGIB3iBkhrggM5z0P4KCayZD+9KlBkaNlnuxpMzu05enYM1IxmcL+zOnId
k9wbQStfQEK99LcWogLtVhl+zW0lDpyhwh86W8Twu8cl3NtHX8mVYaM36HGY
x+32K0C8TQgl+7vI7duAly97tT/HBY0kx/TXCSbugzvkgTKdIkiUnUDqwzWE
V17mKQS/y72ICa/uF9AIO/wwLNuvGTyx6N2+gqDjjn0EHYlnggLfC7zd562f
UypzXn7NahfzqeD1WUouOUdqx97fWUZCe5/1xYSkYNNkN373ndU79E7A+ISV
XJz5zjxrdaFu7G0dq5Nd2T8TiRJz7SLXKSKI7t1HDy8ne+Mc4Y0/MeRUvD4w
RMyap1mpX290ovX58Eep3taYSGvVmByZ+qdWFms93WhWA+/EgmvDuP3ggreq
9/FMwGHC3l2Og/ZklQYZKcy1vqzeejIfvC6/buTUG2PsoqI5nO6uNgqdQHOO
nj3IGksCLA4MrpV0fNX8mq/TPnAO4yJ76sONRYDu14faHxNI8RM6HO/JGsaf
U64VhmQl016dwkGoBs7RhGxhC2XtGJlYbxin/LfZJIKmhNk6KU7kz9dkkucq
z8fNsjZrO//UczGbJYq5g6fooh10FgLnsuBnBrM5Cvbz1nRpfAlm1GWh69KZ
iXJgQWDugmhdInC0s5PPF9RBjJlwWCdVUrpxaUoEwMvLcvOIkdX3q1ks3n41
HggxmxkfxXSoUNbKnV6JDwA07sX+pC/ass5AoatZnv0OcIq/45f1g1RcwgCr
jBY0BiywF4deksscPuHLeeIfujEFqqgrgdxEZMOij/NWG7Y1jiZdWwYamupI
9vcdDYD4+6XAEsa+QVMwO0aJ6TpIN5xKJV6r26HgwKQOa1Dvk8ZSfS/qLxkV
kheW2f/+EuwjpUUwWBRAP+l3UZ+Ax2g0Ud/v2zlHl8VaSQYuttsWvHAatWXP
Fq8xdGQ1Ld4lhaWSleulowX7Rq3f1k/CDIamEDP/P7Ax1v1rUbHmmFNfTbkl
9ks0L4M22HPRucWRdtt+tC2AvNVZN9j8Hp+Li634MkGBTAbSAgM349KRD+v+
C+2csMp6Ei3iNA/WHAHuZsXD1zDWi/yjasAzLbA3IY2mTxZfvrjO1cAG+CNT
Aoj3Z14MYTcV8Go6mXLCmRrQ3hawAZuamhS6dSyDyeS0MGp/IU/b+d/Pio5t
AS/grTWxrXxfcX+jaueLnmEHP54Ewkv9KeIi6owFtrdj3e5ctlMk5C/4Rw8c
C4KU+qWIAeWFNuSnyDnRaOg+95R88RdSd1sRKQy3vZmysAcgus73mKtWuhJZ
i3tJA2KFhp089Z39lNcW7l7iCVwie/SJuS7ynLxQclhzndth4e+nZgRaWQ2L
FPZekF8cneQEkiOTFZildnjVV8V8ILxlY5b/AT6YuDj+bqDPefz5wZaFnzP+
PeLtHaAAWsXZvBRhCLo4LD8W3NGBgkzOLbz3N92WJvJvskkh50H6O6po2QVl
VGgqV2lKwca1lJyPfzKqA44nH+wkpIigynoT6Q/IW/o2Pdb2zRf6gJPkMqb3
+uOLyZ5BBDsZXGvVHi+wjtHLWm5w8f6j6fJbYQcChN9x60R6e6QVIGSRQRx8
oP2fp8c3ncUlg0HIPXXv0Lnyn2XaoOWkm2CzUrhW5blR8mCJuTXklzvaOWIx
uDo240M1w0MAk8bMoe8o2oDrffBgVqxkUOtUaElFY0PWzfbMFx7lhQUBoS6o
9tsNW7eGcEfW7VTSuGCJ9HqvRZjf0pkQGB9FSqjzs16f/RzQst2a5faPmaIx
4sEbTl5ZHDax3y7rKBBADU4nLDFy/OSsFCd5ogz0kCzJUA19arrQpRJgjTSH
/Qxx+oLk3BxvS4ebUaIVBC6Lj+/wThaBqHE3gZuUS07lcyVs62WXYTMyvFqO
ZM8ISNQvkhIk1wEP0vOMl73jU3NA4Mo9bO8HLMePCed81St7jMznzJJuV6cV
HhodfbASqTdz6ENFBXydXBhv4q7JU0zjRyAYtbZ3dRrp2oI7vQG/c6oCMGIr
Gz4258wLaEh3xuFDqiU9uwsNNZRUOZynh6uvEogUYIYoojzvucztLA1yCXCo
LuSsMzmP1EEQQ8FSNDhKnpR5VilzCUXiX48UZNlsj3n2CJyfIlZMy4pk4HZd
ML/D5jirYvEhbzKm+g2wtHee5F/j0AB+DLQKwVIF8jpSxM8/QfpnvFaEKYM0
muaBvRil8Xd2xTmj9yUmOFEjNG4Mgc0zuQXfawYf0QaHjPEhFT8c3HAXncak
SaWdLVVO4LyBw1lONvJdqAdy2Lib5Ay3gD1XePN6myoFrldTkh0ZnT3p8Okx
yn7JLy2BGOstPv+pRureg9PWBJ6BJc57bIxVoPnklBQGLgBQOXf7FXRb6gk6
RpMmyNtL0OQybTTRfIsBLXQhbHzNG+zeJUcHMu73lTxRmL8vK7zO+3lAsnrC
1TFUkzO1IZiZy42AZhmONdUpxHPMu+JBbL05Joq2UcGKCwclZO3lDOVruCVU
EeXMzc/CBl0RAjo33KzfbVvsTQ7fyJLFUyWwhWtxdpCjy+urAV7gnUlTjAL/
tMWoqae15vEWnP7s8VW8FM4/v3vbtsOyGMuBVhJY/VTk5F7JcelvAb9dN/3w
QoaiUOixT6CeFpvV4tB9nVkdSjKNXTuo9hKAWG8eews2OT6mrfJdi3+QWwzb
mlmFCQRz3hMLpG/WDZbFHCKBpYR2ain8hvL8IW1DQ3/8W6R2XG5A4gQ/tJHi
SEM5mOo9bxmYo4eP50zm+qEibVjwovxPjiZxxbemEtS3qM2ZLCP7oUSx51ef
Vu7dZZVoWSdno4T/C8wD+Pj7iHXnS2JbTkFM9IoE1u+N9rbdoqIttkcTthE6
OKEMMm8s7lEhs8aTn233ZMQcZWfoUXlp9aFcZbfBMzB8BnCc8wGZS6eGs4jF
eIfF37DBfGX+s6oiwaKqy+bN4veBr3lVpH4Y7lDcWvk2kEM8yBGmFu6+kLXS
O6CENYWx5Zavvx9NpnYqJGczDg+nkMe3r4GC2N/JdifOnHoUQuNPSlzVU2MQ
rm2Z0EXsmLDcYMi0NKSvvRxzchYt9NfO9coSR0xdR7+zzR6qou3jtWf3SLoo
ncgr/lskUUvnlcjNOWpj6mAAROhiAJGZedOdB8zTLwMqWj6eu31Yu+vCmtmX
5IOYTBMQQA4wNdipeX/jDfqAhsviU/e5M1zk7W4L0autWd07uHbPd0hs0nmU
5lL3C2Yo0zJv/ogQ7bg5W2sv0lQ8MvnmLfCTtbr2o46PjQWy6V/6RSwc8msM
PUf59uwQDlC3ZFo5V9u+gN4900vdu9hL+wk1USowaBo9NhRLdR4v1wPzdB28
X6E/vXO+0ZMJ//9faiGeJXHJz4oqJqPELbZ0EC3b1dApPCUbspwNuq/bJV0q
p4aSuD5/fhgwNy1qpu/qbnHZW+TJBpfxM/rlSPrQr0H9c11JA2I8gP8c+gSo
pkKSEyKs6hNZhTjqibqw7vdpnsl6lN8zU2fl+QfLrk3UDGCUVN2eeEDvNTwp
e31AHfnUCY4zE8YOaBpvQamHkF3PPI8IR3XIg/osHijHz33Zc06k8C87AHK5
wxvT8Md3td1iVduytfp0hEsioAnAesOO70ZMgDGzGGDzkNjK6A+heaiNsmKm
Y6YBfPYE18nbjPx0k2YpOnV9LsZ+eWHOIm8d0DX1je7QYpUvjsXTHrUdB7ZO
dnQK1HIensTANcKw60GYnxM/FnCbiF0aOpn5nHFvtsAd9NOnxLpYNnp5Tlea
HFNUB7G+GIx8kxCxqzWapgT0uiajdpZyh5aPPM2G2FJBMEM2eLslhbs4S+D3
vMTg+mJPvG9Nhe9JSJOMxn4nscmdfE3WPG1SBHic8jDG5+mFdybmt/vgCi3U
JabneixKn/Wi5uDUb6B5v12eVSCXR9BMPjQe+9QPLrKgZsC70t2TYNPsiGR2
H06LbLcXCXdWvhw1ofwS5mvbocuM6uuf+n83uP0H8wFsi+E1v52YZPx7h3+K
MQeF5s8YjtcxWnXx+TGTe147A7n+qvakZEQHV9P7RGQIml74QWhMHNdS+l76
YrGm79ut1zffpY0LqH5ATettGVJQKV917CVdnzroBKVbiVOLNR03ZEaQbgjT
mvymuTJOlXq3ZS31tadkMejQYKrR1atLLvoZO9sm4EaR15efLvMLxWnXUA0A
iBnLPHjZrlVC1VnCBGG+q+7Gs8lWjRYIdK+nj4SJlBX7l+I6YApDIelIWh6w
82ZmX8DsaLRtJ7BCsl/3AqFvPcL/sRq1v52UZkiZOGxe8b3z9sTEBh1CtDw0
C8XOqDWpPfmUB+fHcBwiWAYVOpZ23ownGXppZ2yrYdM0c4RZUuAKzDJ51jyr
3k74uB8SFILCPve+WdMCwSAxOjZdzXZAhf8ySGe/LKR7wUTZGkktP9T4UPxm
dyBA3UzL+E6Nkf3Jw/h/0/HB3wjRehZYXVeVZedDVDaRH2v4sy5IaP26v6g6
ALb7InLDGVeKTz4vn1AQZMeK7zdsuRnzklxkcLxSoDY5Qhcwdoe2QXzCKuLZ
ygUehQ72lniTXXP4rHqn7q/cAXHC8ENei/fvfrNRh1zf5Mq25QG0/4U02WLh
4YNWgTD79tZ17++81Rb14gJfosGJnXHHc5aYQ7CjOnpdXLaAeCSdIkyr2SXG
QH6qB+mK2WThpVcmQKcwHxBnf4E+XZVZVhJS6AvZADqX6EtyuWJjKLLbGZhB
5f0gg6lpZvQFaRtWE1MI8XJKJEgjmKW211lkRy97hVaeqgm0viVTvFl7BvdR
VyRH1kEJOPd0dejlteMAUUYefl9pHwO37bcB69P6NSkKlfOEURhuqCLoXgtW
AzMiBLeabptBa9W8F0SccAgkl5ki3kD2fK7v2tY/Gnun282EO9oYjZnPeTkM
28mjRsl5xuv2m3+OiY37dmKF19YdTmKUKXfDQBVyJ9b+3LVEoG4uucGJ93Eq
uyiY0xhCS9sHjoKoh/FvZ4o+9D89wRM2KAah+/7erVUZHksSOet4V6Fh30kK
BP6uueF0f6kCD/YvtietNLU7dAXLu+z17fZv7VgFrsf3/9nbYwsRxyp4kfWg
UoTUNKcFdUIpw/EN/yx2JtMW0S/QSMMv6RnEHDCJf4+9Z53b6VndmzpnVpF4
ckFcGGWFlM9jgGKPHpK3MfgnHkdWxqUf96ptOPDVGZ1IMWhsn5twi50MDKjt
lZtiolgaoAmUZsl2PZJXDtZbtGE6T9YtJM1QOo0di32HvZQ0d+ZIKvO4rGmR
C6NvK9ElBevf1+HFyoHVrNrVvXTj2/Jc62sEFOUVv0Tri/PuKlGNmGv0hGlx
zYl2zSheiVJtiVPxuD/MJgVPpkcsmUpTGMyMQuKPyWYuXIdwjTcx0VE7JhJM
fc840oDcymXZkIR9M6FiVkHiNfc5PouvFtHkipTueRH+NDSTuTJ5mDP03eCc
TrNUtd+p5+oR/jbdovt3fPbdoesuay02o2Kdpi6NxGRh2IIVh8Sa9wPhVFXQ
kL95O1AZOIE+2WqhLFOkiGy78Uy2HeyYpn/yIpSAUIswT4BP0/qY5fXnC1MH
VAvLzcpCHmXxmchAZyhkAAEbMiYrqL66IkFlEb4tKmAM7/yQROhfU+gBgGW/
w+hWdSOsiLhtEu9M+J7A8UvYd0uq8Ghp0bw0HJZzffwBAj+AI4iHd+0HtRYA
7ft8gEZtvBy7ARiNOokR/daVkQloAfp/EtIXktuUaXOs1Ifg0JNXnRIgDed3
ZYWKC/ui8oxLHNFQlr8EXNzx4DWsya8Okmb0JH+SVHwSDFFYF20bwJ6eeNn5
BxUtvNjHAFzzv8j42A/G4+qWpQ57Vuo5cXHT4/VVbQmA3XTOGq7SKqZyhh+X
D0HUr6MkkY7iVQhk4eszGGwcllEBJhyHvZJ0UgulHO6L4u4k8z+qb9a2fV3X
qicxubke1eD3t+jJIv6DGLjJJZrkdHAreMOggemabyO4uzbZDzaWt5P16WVG
4ljAxOGMDA+wyIm03vTXrXzdNqsFDYEX6+5zhPU5xT1QmKgyhTeq3E+h2M/C
5xoqv2ZDGPhcXL73YHZWLvDrnKM5X59wqPUNKH4vfhKo7n8ik5a3Fr1z6sYa
nzmr6boaZk2hTUI5rFlpkgUfobbbnYRm+QCihtNHVdNQzH/JAsrZiUGQ+5EW
jYp3xd8MquVpPAYue4FIF3Ld8mP3E/Ie2ZBhQACYbTH5cX901KciluT57mrC
rXOp9vMdnLvyrdqv49+NmAFGbwOOMhM8+TfgUeSm7Kwm8F6sL9mCK7uQx/ZJ
373EXte0tGCgxWzlr1GSE6//2ROhPMh6xlFL8lQ+KDYmxmGUYElQ3at69Cz3
THi+VH0I+Qoff4okejHi9zZQ8s33AlZ+a1E5GzA7zOrtjGg8TyE5M9flwyzl
M2ab5JgSqFA2A5CEW19MB2Y7QcpQ0E/1j0ANQTBi1Tuo/trANH3Cd+AuQP+A
9RuQnuR+ntURSL5fLbfX3VrrF6QTODdEXKlItzIgJyLyKmuS28HLAoofl3GH
9Wp+orACsHBQ/w5bfE7jBytvtvFFptHiv41rN+cYwZBXU5ZPWiYMNUy7G0af
CcJ1wp1PeaqaoZ38EcXF24GxKNE6y6w2ER7L4c9S4b7GVMVqLkpSoGTlBVG8
mEXo2U7pKxpkKXBr9PC4CahTMX9HvCFgVAHJXqksA7dXT7cHFrdb3hfqCiSQ
1lTgDe7STQ82vX1YXygrSomBMbEKps9RyRyiYfNwIr0FsxP2Kxor8SzSsIGL
zGRMjv50iXGi1b0xKGh1DKgEybPExxlmhqpwJKP+PxvWbcWSIRcErTs30aMK
Vs/+KEd7wWAOe8bvkEu7HE/dTrGGWExWBL6wGK6QFDs6h++xwmHC1PIc5IAR
6RLvB+ghjkXDQ8aPqEz/88jBs/hJVestHXjVoyjTwFBguUslahhzX0xX6Gpw
HUem1oybom0YSdrpSaypIome7TVjqOxz4L0qikzCJ/xjILxqZ6WTV41RmbfA
0ynJQkLqdmSGUdtno48sf8ZRCdJg+7F5O/cZR+Wjr19ANGf/t8GutgjN0zew
Uik8DEn0WJp0WHl7qu0CrDwlh5M+RMz9aUfADDZ6nRmcPaa0wF8HA+FC3UPa
pUvcdhwY9FQwz41F7NjY4SZPiRV9lc6OZZtAToxwmWEFxmu9ON0eZOslZ0DA
bmn83cqd6G3BM4MlO+PZSR7olkSUqG4BELiRMmDT4M80HCXmSvDCxVWhaiY3
s6MA+rcrNdXtVPlWoFaQ5LMQBmuk6luECfpIh7TE5J4TrUp7QWFiTM7p4YKA
bj3HGksO1p1Tp5yZKzjynFkuR9G4MFneyfOKPtyRp7iLL1h8iKlzi3QvTFHm
Lt4z1h4FVK37L4HeLqne0y/B1b8CvW1EW/3zUTdpTNQQfglCsWvkAtAmhjTE
45OCbzGHfQ3kIbp8Dr7AnnUJJM+qnaevR/tagbwoJa32bcbJR3kHap5p1PTF
ZrhV5CngGH2IvmnBKhs0itBWRpl6p5Ske3n43oBsxXw8+Wj9eFFWidxwMf02
s3a/jyfryIOGK3oSMhfz28MPKOAXjfsMa+fmgfLmkGLO37/eldWxSsbCy2ea
DSNjD96CaXeiD/WKeiOFZBKZtSEywI7JzR/mjxQY9hPAWuDbk43NTvwPKpeH
Kd9fr5zsHNfPsM3GwvKZ8oJy+3iJBq+dTlNJLP7U6V+1MlM4MUrMFaF8NjvE
5jT3w5ZRRSbC4+lP1gFGk1KX60uL2jT4GQJNh0HqQd2mId5Sa/G7nSKhXZf7
+xWQc7bwPpEq8cUenZV994y6rtWyPja9NTq9VzwGOyqF9ta81KkUU/G1P61X
AdXLIW2q+ifJHvdtw7wxHU+XGhPgQ7ocZ+Ayo61CtJLfSH6fN7FYVoU1aazh
tsWwptrOKPhMgzwjvP6k8eOpnsod4W1ALVmO0OG31PR54Eh764aHAvhF2uqx
jZRDSn0LDIj8D3Pr3Nhue2C13M06ZjBCgrT/L4DqdGrpOBQZgmEhagpBRFp0
vSsnBtMEsZoQwu5mXMG0N+2qLI2RaWRP78L7NKahdgWWTH8sXww1XqyMdMNM
n/h3kdVJ+70vT9Rs14lw1qSnEM80R2q7UitaLy0qdLRREaynejc4vL05zLfK
/+GGB6yG9cQj/bRiKN7pxVk32xwoUty+FC6Aw/cw9Vl+UINquky2LhxPa88t
hSkxwhsSe8NwulVl1Y3ulbPmaPw5aS8YFLfDeEIHVig0ShNE7nfZV/0XhgNO
7I0EMCZnhQ+Yts4KqK4jmvYrN6QqNXc83+3rAygEAbulQ7roMhOJWLOiZaas
vOoEYGmPE7NlLjhCIYjgCFjMBXgqsKQi1WKKEIaaq9vmPILU/IMPwMxLdijl
tlCTCuXBiLrTDiSwKhBdJ5rAn8lbII/rxxLo89d/zj3YgpAdgsMsxZ8Hc9Wy
j3D/4c26laZJqc3iG/wvtSPkMjyKsEU/rXe5+QpHQl0/Q9IUiALZZNnChjqH
V0GzIqDaae8lNhMX+l+n+UWO+gvr+63Yr2Hv2l1vtePIaZJxQUQNg4LyiUmt
RpXmYNicOVYTpdyoHVlp3b6LqfxZvOlGtQJX5Z42rsyxosnfJNfVrO6BPSuO
7xfFZeF8B88Br6BvG7d6Qc52qNKflSQifsWpjsLksM/l5iZXqEWUYPMzlzSz
M0fqEPrHz3kgSJnwdpoNNBPTSzEp4Ti/2bhl9TRbmKONboJHeVZrFgoVukuT
VMNwVF3qA1Sae+nPJdagdq3osEWDsXBtMoBRgz9nP7r6+m/y3ayeDBft2NLB
M2gLsIJfp5I8vflSM1bRIGup61kSvgEdgo9dCVWrc5w7ay1DLOwXwK7psxPd
JWecBwNxFFu50RHcn5wbfa7w2s8R4CKujmih55BYH3t2mwaqSg1BGDQqskjp
nmxPrssKtbPokNtFczI99dtyUksYMVta9jwIgqSo5NGl4UVyntG2gGdnsa0N
2DBxtld7HBK4Euf8gAsiir7+oIIDz8zaFcnrx0nRHktAnbj5LXVvZ+hGndg0
WAnQuQZUQzWkvPtEt4SIHHmYhTpeREhGqMuvQpoOC1FeBQFiqedbjJhy27MM
VTaOGAEFxduuEjIAr33R1wDPGrHDR19DbeTbUEj7hRPGmlrc0oafgoRqCSgw
+zcWx7l/QKesINaWuka3Ni4gDzTowglOZZeKgEJD7Fp4jZlUE9sXFF3aGcuv
1aPriZAz9IfAuDDIUIGfKzgiHe9gk6oj+6KiXZd61ZNHphinZnkGUQVnM58+
TMGEpWPI/30P7FAg5uguUTe2an7QcgOGEeDtdyg13WJV/ZWIOCDmFlun4NE+
J89L1EFTNXoZuVKf52GaAIrgDbV/MDFo5lwjfhLOLThWePfO22goOtc5R6C5
ZG/GUKzzwfzR0AtrpY3dn7blbHl23od5OCtkuf31dwMScOHneC1TywZ8+S7c
b3tFQzZuq9UcsXFipN7Q5o0jo3InkIBDND52KgmIMEPijNf6p3KwHphRQhD9
kEVZ+z5zIrReR7sxMOYwYlCRxgxFvvZCVxUtQeXHf3toVuiT8ainZnLZXu36
CXH9GEqZZwR7+z3T7NafTjcfC/kurwIpvMQZNAN4QNNkcUbr60DTzYqc/LIu
yuFgmN1E54k7CnzBbXNj217MNIJplc7lGs7NhKK1LcRfJAUDSkpqlDACIlxM
uCijzZaq9yVNG+T+9u1VpHHdX7VTUYElKZIf71p81hPqNwRskeOZ1/BJ8Eqz
b2BLIO9maCQRC1dPKvgJ8kIZYiq3Oqi/AxExGSvFt59OM6vdYGHbvgfnjoKu
FDnOkbdy/ZrTUZq7ltfo/Ar0a/ueSkUVIlU8/nj8XZXckcvowYa13cqwfHcC
tgTM/iQ4pcj+BEPBXETZzMPe0fw5Yv3ucdDfFOFrxNDqIt9/xxyw10RNFdD8
SzcTa7iCy7YI5urEu6kcZnILjh0H15rsIg/BmVZ47WrU04aO9EdB4FKiYw2m
kO1M0880R6Zg79etaP86UiVl3xhbeB0Rq3mt/sM4DQFksmnD3T572wt47QjI
tF3s4qLUOH73T9NKvDVp4uQHp9SvRmQFa/t8pjqwW/4Td15V8fO7Pz8mlttd
8J/+Wrjs7lTnuklQIom4myiBMxhFu5GgIsvfAESpv5A8fVbYs8XSWkxyeHXn
q01o3icGuCewRuf8BjxlnpDB12qwuzvcYzrQHNsJnX7k3tI6zcKVyE59mMJn
F1tnBGciB45oMbXeVLR3ZuQydG0iqpTgnhi+RyAkYGbv+E35vmbQn60Y4frq
kY98mLKvNkJWJ82BDEfk+RR+tDgRxerebwsj8vy91/f3zT4Ed0ckbl5rIFGj
5hgH/8zmFnPMj1S7Sk4pTSFsddRP4xn+q07JEyOhcBvvnLYTiGW5IwwJp4KL
NvEsKMo6gY5Q47lRYn6cEBp4GE+VFtFmXCyinNx2vMmYD+udOjgQoNG25xFe
7kkpPc5W0rUdiDTrwpY9oVEJfsw0jBZUICFVMcZeqlLoTN43/mzxnAcVdgrJ
3BQLvawHJ6kRhhvPlTY7225i7vLSZOQbXR4BHaAJvMbhB6iQmOhQJTmCOcIV
fasPSAh+F9xhGVtOpvqK1VN03KUlYGhS+UimVF0RL5zpE/bBEYCSiUtyBFlL
F8wcuWv/D9t7Rnt8tG4JKmWsroZRfzknGusWTcouKcQf/P136ek8gXAoqc6Q
PBQMBJdBkzXE/Ug5OLLmWW6mV8KDI9qwhOnoWuqFsa2W0JWkIxWNM9p7LpEh
A0uxqXjun8erG/qrhRvP+jHO0rcBKrhr6LYM0rWjlIT1E+gIBrHimiUr6LVh
Gu0ostVLXe2AUKd6JabXjy0A5pS7HRW2Jtw/V34SY20yDi3ILEeRztkTOoCR
eTMeS+ISB2VWLMaw5Y0nl7OUGfx9qg4CEcwYeB/EPM2IXsAk6i89A8kIJpZc
4ha6EelC25rFAwBqltGeMQOnrtMnWwzrfiOtr3GBZceqDL+eVv0991kfwAJT
RXusVEV0ncRZUIWHMnhSFVvnWEpZ39MBMOr6yGMbB539rS2d73CNsDllzP28
j41laP+XDDTG/tbxPx2/32rNsa3CNXdxNH+/4l3tjnVjilIRY2sKAR9wXohY
vJHKaAaregsv0/hqpKmFRTHQ4GKr+QJOcgX67wbNxwQR88CrMS5Vp/czCmX2
AseN7DKrbXgF+9gEhmy/S87yATodyXVV06MKFYocdJ9mmvtzeyGoh9H6JfV3
ySDOxVWjLHhfQlHOU50Fx10+ALn2EDSUL/rgKAXc2QBmrZcqeztD5e70gIeZ
uMYFqHeJE32BUTefFEw+e3nrayDjp6Z3i/teef5ka6wMaul1GTLToaIGxdJC
8baAEqkopVydQgjA+8XHMD+/SYmpPoy8Tf/TW9dYMDyRDMMrOt8aKMRGLn+w
PF+S/91xp+xwFbdWqHuqQo2yYyR/tZiUq92zD9BnmSpdEINbXw2a/Y/J/hJd
fhHMzxJHALZQsYPRyueGgt81hzorb0IoDIA1huGnFbNLlD12Uo0aFxUmT8a7
uUmZ2x1CCTnvbGpDvfoLxFOHQE+x10rE5EsnzE8tBBRDJi22zSbe5tcvvbBN
r2xOaYH6KDBnOMygmo35HWTnM4gZhy+AR/lZBgtTz22v/8iOQpeNJzi2GVrC
65jTAX/kEYPbl680+39J5T5SnBcyWwaLP0C0oV0rBKl65Mg9/nBHVuSxGbEC
o+pGduE+qRQkTG+V2q4mTtdlmn9PCNaH1Z4uWM7E1Q69wDtSWgxKd5sk65bO
jo0CP0KvV1ZSpyFRgc/8n4+4QmR4FATRKGAfgfB5xs4FYZAkxyotycz2XiX7
3Tyxc4Jrm9MUfCyju9TpWHkFkCA/UvZnOPAalwzsQ2jaJwsxTO3gf5z5PmzS
SAptSp42m0wxdrb7rq7zCC+DMpcSeK/DtCdZJ0Yp41D5bzKI6alVsrgqVjRW
IYbYArIRWBlH1ryG3j9O1jSl6Fr3W6jYzu4Fx4wM3Mwv7/6xZUWMk3pU15QX
oXTgPkPSBKP0vg7g6GsmPAZ8dTEKg2nqPAynNtgFaF8d889Iex607UmCDPB6
XGbkpKfnYOrs/nSaV762kXhz4BfbhJhdhNRsirZvOC8woKseYdzRof3HvoKh
sUU8bAI8g0o3G9eL/wjJaVunS3JHX3nPVCuR8wZ6V113bK9j4SSQYy6aU8Gy
K4uzEKjzkbtUGL1p8EBsLQBtAvKHeM3Z2zn7GU/AIsdqxOYeEynX+zn5VdPk
w2rC3j5nLds1mNotWvRO5kZ6FZFQJjtgkLUboyBom9PWwqOD6rxa7culHPjt
TShTvLtqu8uPOtBE89TQgmPMRuJlttAVbY/nVwEDP+2zeWdJlMhKY0R3e74I
2CPTwkSf1Jdi54smJ0XmvJHGwzu/aErlhbEGOyPxICrZ82X2WkD66XH9S4Qc
4aCx0InEYyagNq0JQXohC0Cih7bGjQ0xQbw4hq8fxCmUEbJhPLZJLNX15/Sk
qAYtzrK0yJSfMLjwLeGThqj7L2xb3+1A/e0xmhymMOBAlSn2pet2dVPIIxLP
v/oWk7tlm7P1JyATL6MplpkjHSozCfF62t+J5YjOTyURUx+6vUGWZxoE7QI5
QMldtgDhdFnc8KilTv9nN50CONDd2vL+d7sj1z8tgey5j4IjIxrubvr0FdmZ
o0XwG6JAWVtUiQYU8DmJHfu09qdIjYRWk0GXlB2ND9kvupElg38AjllfWHJe
id24i9uguOr6IWUu2BmHLp/+kpGccoXhym6zUD9rr/9uQq/8VT3GocW9V8xD
Ruo3IoczVrqym2YLLMwd9vjVOSmXZKn6s2OWYDN/SJ373O2RjuzW7okeGCQi
idx8Eo9jtesQGTCj8vzDl6emYDSy405F4Z2ITuwzFebiQ5bpGo/j+suPI8R3
GnPV0PzANGZYj62pHX/AC0Oy9318V/nlIiYIrY+ZjjoOGA1tncn9O4dUDoUN
BQV0fkabqRdlrKpQOAXv7yGOLRhRte9Lan/DBPffo04Y2196XwA9nPpiqeVt
/Mvk4EUh9HswR1gNXcKxnOgLIcB5z9QLEx4nbiakP4ZKPOBFuHPDO+Bp76VN
KdjfBytAaG9x7AOoE8Qffq9wzgAyZ3ykB0GnOSx8uTcQbaA2La4jTMbVf6gm
Rd6bGoBak5bN+jZfkk8BwCWXxNJuWiAO32ALoGkz+9A+8dec1mG+YXWmv9gv
0giAj0OaFQ0GImZmuOYuX0zlSIygDR3D3vf+Gf+repnWm7R0SEfcrsSwPNnM
S6oRhZuLBdqCZKmmAO99yL7l/vKN8i/XGV4suu65MaYaKJUdIfT4miaj2EBw
otx9nQAQ8rxlOVquUtsANIqAohf55WZ6i+ITSecJ+CfWeDkCskEo7zpdIFPD
N/QTEEzT0pl0SUSmbBWTaWVJ8P1BbvmlDho7I9ncGFHpB01ZXtmz47g4GrX4
i7l7GipMXB6qJbwpjAM2NuVDqObyOuUNoKZAIeubQCT3mXlId1+HaA/FfqlW
pX96NmTcgU4ZGZy2n8GOlWBHZaKM0RcUPGTkzSKJbbI368RCrVRXp19aNFh6
V/YhH46MKzTLT3j8xzRaecIp/zNPwPPeap7laIHmQfgBWH8xw+DUqGBIkKss
CqfPYK0Dp0kCLr74Ve0nspewg2FwYw1vb1Qc2navb1uNLRVmj6RlkPyJdnLz
WD+o9qyWvJacSJeCVlWgPhtp0P4rfGdnJBbJ+W0DpTM5ESSjl1R/CmRTjdoY
obFDF3k5s/CYkwofC81h5x/2CPjpHilDpGWCSP9rm/MvtchJmFE1YZRN/Djt
vbyjSlyIBKl20OqW72BQZVr3bIuqPvjidrPQo9ErSyT8k0Kw0NWYhFExR9+0
N/pQU8XPeExFISIBj7VUnz3JWMOHK333na73mu0lXIRaCKUpDtzsTeePVLob
VlYQ4h1SscQ8lvZ3R9FDvXRK8oUL+qjP5YMvCCHsp6K49BkeqxCdIYjYCM6A
ndyVaZzfYrLQZMWcxEejhfMB0KMssWjnbV+Vxazan9jxYBchfgy5iGmbk4RP
Ik7jpgaNnNlps+ZiqZNfhRjt32cnoAINGoQhbMsD4Mm90zkwgAkrlfCRk7GB
D/flsKDnPmGDbd+Y5we957vFKIOnZsnJGmarmSpQmZ3OEWwyQFc9GVwKBHSF
hB7+xCTyEJIVcBnX4jw+0t5DKG6TG72EYoXTCt/oaIbGE7pZybp0FvhmvE0u
GMuXDHdx3iALP3x6/yPPRmDh41sryI0xLg8Lgl7u39IbqS5mFo4eqSezex1Z
38sFkyffIlsErrGqZ/I7YLPNjJETk6qVILiKguPGj5MyIiznrPA02XT4pp+a
QFyPpcZNTXocF6tkQ9hyyVy8iCVvvVu0a6QYatH8c3+3ZxKMTJmkUp1zuTxI
+pnzDw6qqkzl+pTon9OH/uu4wDVeRAcXbIXLekg4I62ugZd+27Lx3pFSINmu
uYIL/Q9zUf2p/UyXEU+FR1uqLlXGSjFQy6pBPiGugwGvMB/vUYH5HpxK1zCY
6iCC/1RdX3AxwR+kibApjnollQPuQJMc/AioTcIKlWvuAgyIkzMY8DgJnwPK
FTFSQfGGloZ4uvB39+exUSVQs61wGdGAUcfLrEHp24LNQzbUtECEsvdyJXkB
yFLgJqqwRZdShBv/WYzmkTOT3DnXCbtHQ+3hHKQN1RJmTBJwGojxMcOA1lJE
gQolr4FTXDwp6IfcGecoGGZZokX2o2S4/Yywjra1FRArGckIbfIdXiPosXKa
sYm5OCar8RVFh6TEsfbSNUR8gBdcO77/vD3eXJT6beLmpoYV/9JvW4xTkEiu
2PwP+MRAJ+VFMgHyUuKWGe+3/B7ft2aQhRj7ur9/g2fXGGjn/FzBprrgN0Af
sdTfQIRbKr7/ta4IszA5rAuIxU3r7PR/cluQ36d5EMXvF8qnABokM4pn1JZw
8Ic2EQ89PFswDsX4ezp+v5efzWhN+w3UXGWXC7zdMmW1HwHWZDa8dKeYs2v2
SnR3YGLJq5UVtt1LNMqiCJwwlggjagR2Ha3je7X5dgP9aHSnbprFZitbiCeB
FemKs4CZFQfMU/+jLxt0t/9DjUdOaUc4fROs89EK6M3Ejhn68WuTnh/lp+pr
QMS1imETWKYkIGZqYGP3kBFfRLIZpRpcsC4Vyg4gRBJhpmc2WOwBaUt7cKb9
mN6NA1vNa4J9Zk2LqSD9Tjht2RJy7qQCtBGZA0/VkDYNX6GSSRlWPSWfowfp
vl2X368AVqo0U7u4EwZHYJ4vo78IF4WKA+ELNYlZQNiEgQMP4Q9zn1GG7nXz
lombNVyHuR3gTBz8+y9bR9SjHzJRQCPfVTZf467u/0VDFhLwihStbf/H2YIB
WVwF6uXmQpvF8ne1FJFX2CQFSquB0SiMQgmm2LGFcfotbcFSM/4VmiwQGsL6
JXa9YVd0JmS5b8cq/BzYqx1fFaNlojlGuBeTqnTePA3CfahBES9Izs7nQLCg
T4dEqzLZ5H0FxJlceDzeC92W0Dyze7v5ADnu5KBSOiYV0Bho+jsKvhohyHsQ
4z2eMSY6COn65AHggX9D5ntEzO1Yt4W4OgsFK04BThA9DuADKymyJjQZoZ3o
15+GQsWBscTnkE9LWAmy7hj/cbm1FzFAyg5UpzbjtV4haEVl0zEzhdQwvCfC
uLOi27hZvr2PP777noq/cSViYjsVuzp9hQnUI//ddahZjbEHhK7ds3G+Gfcm
4j9EcUY1pG/FwlE+cg7ojvCrMNdPJNE+Jk9ctWNcOGsfLNelJr/h02yUQ+5F
ItCMKQ9g5Hq+vDapEsyB+jZJQY9z0px4Sa5dnVH59Dhe19/T3WyjO3qVgK9H
ydEXZZelEg4FMOQIW6iSUkjGFe9M83CNaSPxmfMyqKO1BoBMsqF3dbeUe9+Z
6AfGe5MyQhlPQv8yRZiSGGY4bUDKxq9Bz94ggShSEN47ZTGlHwxlfYUyOdvG
cokjSa+BlZK1Pv9XX+YNcT0fqGcFPBOQtdqQ3UI4aQC9uCpVhETvjo05EkDo
vM0+xwPfGMRI18tAfbEgGbUsEHwzRQO9xO5kvZ0nLHOiRZQYJFNW/8xPueEG
hTEHQL3VrOta6znoHMsShUKtgMEm+33hhUfJPXsAfP/ZhsnwQzpzM+JlwfSj
GYhS84000ly6Zn88Igx5cMP89ju6BUtpMBrhoq2rLRxtqwejo69Rf4YeLR4J
MIfq9axt58NA0rUqiv5h5E7KhfTfBuH43r9+nGtJS6PxVsqaw1oiRWnHyY9B
bf5etTMMC97g625UMoGG9MUenAayKs/WHSCE/55cEO631PF6cHkk04TmhazI
ONwMM1/kWRS5W6TxKyNqG8hdl6h+v0LMfe8IQkeqcgqBdle6DMOgRZOIeLDV
Wt64RcZJNy2tFD4TqbSPgF2G/OKgGPISN3Pqu2NdKcfqmws4bnbrSwBoB71i
v+EKuXWG6nrUMvi8etSmpsdq/MBdzwRJS0PXBLrZN4JxCLWHvpt8B+D/UBWm
avN/xo9/4E1mLVkihFgqMHksbPvOGZ2YGittGB6hJ04NpQ7qSfCEg1F7fO70
2BEbuZTDGXd6RxwLH3vDpHhQjqer5hOc1JrQAigeJ+vyomtlzybeJaZ6Y9qa
LqTUvy0ebkCuV+FMDisoXIYhmTDZ7i3do8Q+q3fQf4b0AX9xJUxgb9WYIXOi
FD++5MK7ZOKVSOze+9OXh/u3F5mtYePYR5K8t6BBgduHVYOCzgRG0gyx3C1X
sHUNc8RusrPWz2tgDiSpfj4UBZWbcm56FQ1HpoccIpd03n1u2EZ6ag0lvv0q
BXIkg1B1kael46FjKR7OK1YLyLGgI4lEmtTJ2ZJIU20JM61gCFwIPbm06fTI
0gxKvvYjzohhiF7DTMEKTcb5gtHUVvoSwpB5hQEDLLdtFvaO/mqGbAdQT347
3shqwHlxJulTr5nrmrPI0mNS3/9becSzXRfb4o62wPIRRrXT8+YPvMG0eXzC
BpEpMAzzpkajSCR6dbnMr7LV1Mr2N8zTVzzayqSCKOnYoSIiR3Gnn9CQbn+e
HJ0Es62TdKApswIJyQrv7Kl0y/oULhAqoBM8Y0lzOZ1T7emuktp1GIS9m4NG
bQ/xJuHczyYGks/ekQnWNs9g4f0cPrbzrv6laiCOhRVLgANKX9q03+on9OiI
YIfF0B08QmS2bw59obSxv1agpB6TwLPCZrWr5Y2UL9faDn6ZeWyNQga8Z1GM
d5VQB+dokJl5r+6/HY0n4daRGJsg3MQsFpFGROrWljIR4wANmTaanOb56VVj
ZiPKyPsrVl9HhPIa71JPTCpVueY7G82aeiU8fn51IkwEUW2/tYhjmZq0eOfl
WDTYcfmyJu5rVVhD8s8jKe0KRVa4m1/8WPsojG9sWqXHqPAnZnUKqWwTHlyh
TbLo2qDXCXzkfWEnVwb0eX1Pcjev9fCYuiU39M8E2m9xdtzSxHqfJX4v3brW
+DtPQvHOXWS3s/vGCOFxD0RXRo4mxuzqXxkn69NddZxlLioPV/HEjd5Cg8TP
EYMt/jM7LQ0jd2c35Nwy8a24uTIV8Udm4laW5c8em6QFJDOxUY0ttk7xnNUf
sY9tLOeRenLOcKJPghc67dqHADFGA+iTjBiWOeBTcGDB+ylXo3Sj62LlaSRo
7g0Wc1fCQqkUD40MQGoYFF8uOMkoZP0SJbt7kFI4585eR9LRd/LURioBoM2H
xCA4fSQs5GyHlXEUIisErXuANepqGMNud/JVqLdncmBcKTUEbotogQ1cKnpq
8XA7ZwozeZMG4yq6o5NtbSAegk8ieb1ou0EnllYNX2ztstkpJixhx2scIkU/
TUSfyM64frwkvNO9/6qfpCgEo+djpwzjwfFjZca2oQ8kk3hr1zslvqVxIR3v
OX5fiHB8byuS6P05HCP84XjYRBwUTvN+AwEpJYy6SCoEEy6Ynej3milqu5pi
gVhFn9co+dvHgH3mCyXlU6FNS9EaCnHn0CnM7igfJUolyIgY2gk8FnHBBKRK
bRGlK+DfI992UMUWOkkKfK4l62YAEvEAf49p7HwwWrlpRG07aF2/I3rgeLC0
DfDSOAcwyVUI3QrZd+phjcwBM/Gbtld2wquDxD8c30xXkRNDDym9wzMvO+0z
f2UmFEXEr1QojZfweI/CXAqTyz9NhIM0j39v/qBsSbyuV3uEX2S9tKbQMaNc
B2Ja7YOGXGfwrWkhNwNkwu1O0XaPOsd35UMgmXWRgofD93bu/6uD2EbMJHaU
uVbcFUxQpe0PP7WO8Dn2VcWVZO0CUGbXk7Mr6T2dxSGlMRX7W4IbGoKuJEP1
RN4oaV11pjqQVU5RGgXy1W/q/e+n4OMQVF/xo/TCRdhMWgHHNdFsnXUC57GC
pa3aie0VO0qKYyXASUVg2CJHnrPeg2nRa9KrW9hHtioJm/IaXDkmTqnVnaU1
cuKJWrD4ke9vEoetk/GomsRduN4P9LOlail2Q3VyogbH1TYakMvpd37pqzVL
l8Xhfev3bl5zcV25DqYe2gEYOsEkdCd+xooOfv2P1pGoepnFBSIeCtm9H7tj
SVRZO5taod/R+alDazZFd4zowHlvLBK0dvGZM5sC0mtbx9yvIy3BePfArqDQ
TGSHugLIwMF2cWsqiDQBviUigUEMRzT+6NdG6TsNvDdtzr7EZpuxqbo+T7u3
AN1Ra/yXUDaJKE699WjTs6n0rPBa4uylMZDJFqi2GoEC/QUiw5AuCASj9Cbw
fcIc3rS3tRNXVyJz+866HaerED6hRhyfQi0WweoIg6UNVKO48wHSl0eaF7oh
mYddYqPP15vLkkkE8HWMASt+Ybj4vG1z6GOdGBhW8EGTr6QAvAiVPyKP36m6
gMn0jnQ3Wl/ZWvzFm7uZfS0gEPdegFKvCdG+cGKMtGUP6/oGYV7VjSqMX3Jo
Fckrwbm/Iaes2zZjmj/gdSrSEwC7CKmBzl/B+4GOXWKq1teFY5ODtBc//suM
BDZEUaIOPLSGqNMgj5N7RIyjpcgmyw0OEykIvqG7vbxoReGSCzgUCPM0Kjaa
ZBcuAL7ExYWDXGU/cCvQ9/9Na35RW9ypvwFG7ZOmZ9vYKSVBLK1UqZK2Z8oC
SwC2NkYnFsS0/CUiq71kyUtB40M3mpNZpE4CZbdOS78UVZJ2irwVzYqnI7ct
8fUZSvaGaMm7B217LwDdmNXh6rwAyRhnNRLe9hLzYhSRJZEoFw+99vEA23wP
lwunDolJinDnoMrI/7lthMqs0NqR/tC+WQAOd9Ban2xhGzK82Tuz4Wo/16Ht
QvJrWi2ACptFT8d+JizQcQbOU491RrPtsPukskTlePQwI80it2G7ji4SgFy7
iAidsW/SiaEXDyoyAGdI4c1+k3uTDoRL8UJEdXyyuouN9ZYDzZgAw8JNy2xu
Af9vJiy20uu40NSmm5u5Dq/W3EYqyBYWPKWJBGCCmhSsPVJ2p/iDS4lNR7gg
sYRaJdKqv6Sv71dICZ4cByvo8Hum+6bE4R2TixTWMU/nlxr1rjWMSPzbjWFO
PPkXrnb3qPw5nvcBoIHEkeGj2MuxCb4WCgLqstAbioVgNFIdqqc9vCtI4+Gn
KIN5u8KBuSzsLL3UXg7pp2L/1gxkCCx4oGcwhFuL9SThBoh1AS/f4kEepSpn
KkElb2GJa0O8HbTtXEPEpWosLvVM0tVmTLykRznFtLt4rz4xeZ6WfpT21ORK
OhD9NTss2iTf96+YthP3IRRjS1WK/WaaPiP3GNm6JVvxIW2pNRm9dnUDDqGU
4xVI1wuxIWWae/DYSrzmzOAAkWCtxL8TlZo2+fLWmemWPZa8K6ZinAtvpeNS
aoZ1pJFjaIJI66QBmSr5V9C2/yop/VVNrJk8I8uQFb2KlAWkrwloehdcGwmg
7nc7Tjb082CsJTlanqloAfHUqKOcXO+noYCNUpNeK2LNEjP/rjXjfZBlzuji
kQ1E4zlgDTnMHaHg2pB7MV7A/SDjB+f+d8O2OvbX4rZrlCgT2y+CSYvxRNYv
3OIRd+iHiVgfBb7QnNHrf8ggQfnu49hKCAmMTXTuGF4DWkL/RfeJa3c8nCRL
TbWLJ9wb6ZYA8YJM4FHvkftja7XepgBEqn4ytnrP0mZkZfwhmLCSajvzKOLa
LZ07iwEbDg2mX3RWgg89EsxvHZ0jUO/X87/3+nc3YlTmSt26SoTW8Hco5k/2
HqsyFsmJsn4Ab97+rKD5LmHNxQaYKGyP8cXXfMe8c3CNOxVS1DSSMXTEm9pU
aLfERcyJ7mkHYD/t8gr6XgMs98g2R9tKpoSFv26vTx5UZwMx8jCbR9Ee0vmv
dW0Lz+5meeR3viaw2he5whiiICWjINkde1+w3wrHOclRwVDQsZSCmTP0bzy7
5OHmKeQJJVY4K88ICrSPM6epaOb7VvV7C1WzkBDID+3FLpvmywZ5+wX5/ILH
ASHn+JwFdFmcwGGddr3WNf6UeA1fj2OFaL4ZzFOOuIIEvGSCe5nEgROfFCOB
f6imhdMsfQIkb92oCYtXrj2PNxmq9sEcQIrW0uzV04juBxe0+f8p1bP03Mr+
5X1o0JjRPUk/BimjN8PDs0BMkTcRI5pB3EyUMOt8GQFkRxPJRj7a6zaGfsI+
K73Id67BMstDJ2rpRBKO02fdnotPLnOSaA/YzosK3KKuWTmdNLkn+5kB97hX
P2HT7hrIt+0yN0C45hO/SZe9zzI3j7X5neprOHtDrpdJy1ncloS6no4+Ykcm
KWx3WKWFFJCcS1tGa5vSXbgdW/+NPe5GOsmd28gCVPeFJGwD66Ga+ZCpFKjK
zij/z1W0LA4inzXjMxJMuwz/Ld6SvMFxeg+Zi1fKyE9AVei0hF7V5WlwAabf
JxzY6QzWvPlU41TmOMY4g++5cUpJuKeilRlP3pwYGZk4BCc8XQBuTgUb24ij
o4q9HyENGJOg9A46S8Ekzq0+SIu2pQQxBjR+fKClcoOQbjCGZoBIBkPvAhOB
hwMddg/F0Plcr/iYdzFIR+HO8WjWqUt2VBDMzF7j+cqc/aoRDo4Q8I/5G3EI
FOcsoNZm8jH6yOhu02nRfpsXQzXzqsdN0TC/69jUhYZDo2RQWYEiOCpYnn0D
cR//5yarTrmVV6IdkWS74knZhtvB0FNVNWtc6/izuzhVH37TLNXzjaBBuCCH
l2KjEBEsvPc+RxhexhXremmhgOtqEw927pXO70I59imgKJh7Jz//9eAZ4+wl
70uOebt6EokAF67GCtCuw5rOtl7Cf+OZgpbEja/neu/kEYlwOgm45y4pSgOE
sXyU6DdL/YZ+exgbuV1fLr8FJL+X+KAYUuKFq2gZU2Wwd9IraGbvC9fr7TXS
oVsGnH4phj+FSOZe2l8kk4zmUVimY73m0e1m5vmjEwMJq2g7KuiquKfogkO+
u3xwrKQ6eTJ67c6GuET2ZDLFj4encAc0w0ZW/NgVV4QpR0cKg4afvATVEEj/
cmlx3fzKC+KyeeSTV/Ngm4Lo81B53MGJbOWP/1Oe4bIQ8wpGpKyshNVt0Iqz
RB9YRLbLGopvUd7qERkXWXOX3nq9AKb4E4m5V/vLT0gdmSJ6XsWKNF3+o3G1
lfAM+8939y3k3arMIPw6RKdc5PL4II/onWzxG1WGfJm1wqlQHz2wVF6VdSHY
mr+qAlEaRjdx7FyS03t1oBxZJxDFtrNxOwJwnxP6j4TqKnppOjQ97QbEhRW8
Dki+aFnDRC7ygKHJmrg8UCXV1yUJoGLV/DwCUqEidjsNr0vJng55bQYUQO46
U99jkRetXqkIsWezcBO28SZWBgwnzkyrjOwjt/vUmcIpKhdCK1uifbT66V5Q
htEZMBSQJ6iKKGyHAyMw2fibW6Y1o8VnnlPB6a1DO1ACB2A+NZqqPZuBwFcR
vJhRXxDg623YHtAeWQTtHtwIIPA7a+hsfxpsvYtYlsbkbTtv33dIC+FjhUo4
AsfETy7ZRk1o6n3PO9n0hrIcroEObjxC0rhFG9XNaimMcM9O44P4UbofFTRU
czybcF1WvGH4JuRGAO1kEJDTwPs2wHxCxK+J2sVIxSd5FAqrgbJ1KnAituib
X4dOhPimYC5OCQFKOiJWp4+n6+30xeKLlMu25JHVzc4bbAIBMQU73cEmWBhp
HWRSYsNqBHDOas5J5U+fvb5nd9RQBulXdB41a9sICDUhn5+4JogWs3vX86yr
TWHtCKuadbBOqD/BVaA/QI2fPWYeuQ91dbzkHux25Ba/pRZVwXIJODpFTHf7
e2ONCAMqRuSvxZ1AKUL7SWysNMZv67R16Fh/D1ym94XSzFEvYzTVActfcTM3
Jqjy7oqM+NoEamOCsAb2BLwb45FDDLGmAkMgKkFWepiBfMi+LljnT+LdnYnW
DpXdjoe7VKuhoSg6dApBcCnn8PV3wlbgILsWwEleMzj9er0ukM/BB0I2rARi
lIjCzNhBh6qn98g1T+sIHDQQ/KfenoGVpDIlEw16EtHjChye3qP30eNCvNFv
hcT7ySc0STdleTDQoxF2+z8fLx3UDjWZgM4qwxZoalxX+oUhT2pt77IGg0Mn
k0KB1Lm/9R021uAev6W1FvzeKL7yTm1XBC4Ih62iJYYQj1tyJ9fGYf6qZsi8
VDx9ULj4kEZbIH9MNpYV5nSBT/9cWrKEfS+U8inhXjgxRI3a1aGsK9dKgWRx
xDiFHMyEQLm37O+xhSliOmnfPpy/AroeyrGnPLI20ORxG1IrugcmJ++djAze
iZ7q/N7LRhIadka3ZAxFj1970ks3abh9c/oxXZpKOQ2mcBRjuRGM4eBY2nJa
QwJcTkUmCm6GfivzIMUE4uiUR9mpO0yBUFbwZRw7PbWCBurVYax21RKFNcip
YUl208Ih84GBlWEqRdJ54X15ko2AiTBHgEaEkY3XSkvaWWtecigTJlVcWfwY
QN70q2glr8N1rw1uK2C1C03gqA7rKOf0AKN+xj7wHdSKkk/9OmviHPLMQzfb
ja9A8/FNL6pYx/DXpLuyCV0yfc/opdDFjhpROpVqH/UkunVTWeS1YSWdnDJc
U9lenjb1UIPvI5xIT1WWmA0JXsbxYp76JnARJOg3Tezp2FUUA3/pmy68n2fe
cYJEcFq7xj80nPS9SQAGGxKdjj5W/LOpHO54CVmeNHt9NlDobneQgvUbbPQ1
/fZuQ8ZEZAPsarJF38p2ZfgFwAlkiPu8HVBAxBN+Zlx1oidv/K9WLC+jSJJF
2bCiUr5ouA2lORoL1SgRZpI/GFNI1gBHy6yygtDlVY4y3DM3Z6lS4/zHU+B3
bFkDKefqJEP/r8t1ypCo2Ys+1dWztrCRO7XkDvJsunnH+KTuB+gK5/C7VvU8
52ZyO/xntEap8W4EOydC4jRzGNfqzhsdifvN9cQtY6Jp6QWdMO6J/uuD2gRD
ed+Q6LsRpHVfk6kzSXEyYQXReyjg5SGRK4lHIITXF6jraN9WtPvQKYh0tdE8
ZJq9pJl+21ihblowdsduAo4sR3XQv/dF6muJMYyI7nlvRp7ZJGXZo+1vhL6t
KZNHeYHhoZYiTM2nbxH8W+Mn347HH4OqYwQ/NOLtxjZcmnHST87veug5aTc5
wnc8wK5YSwuLxWxf6Yu//o98dTvYjr616v6ojoDughSuQfs7LDurirtc8T87
PP5Cb7dFV15mqb3OCp6zwA1BTImcn6Bqeov9p3OqfQPyUW8jeZCgEsgaA56E
lIZeqi/b24IczkC+S/2a/LuAPnF+/IN7SRoTmXWrylKpAmSmbR6UonF/aYTn
/QrbKIMFwB8QZCeQ+IbDuRwmjWfUlFRiz4+PTwSoM/VWzLcPT+ksslWjy4hi
pZIU8rYcAm5RqyEzHtfXTJ0tg4xqvGQ7GX+teXnY7FPGT6RUA24yPbn5Bf/K
qbJtotHlFufY5ZElTca+eJ1DsSdSoYJR3K8/U11phczkhD8woNYbSAcJ7Ni4
M3G/rTfF7eb5AtL0JZ+eT93NTqdsvplNpfrThvv+9XAx/sYyR9mECk868VfP
xq1o+nctwUd9LtOoMjDtAtldBlOs9LhWgvIFMRAuE73s19wXDrfwOtqidMqy
GFFdnx7sLFEc+i6IKlczGsT7mxXVAvmwrlW5GrX4ugXwj2Ed36IRD+oeIBDz
w6dQFZ/7RId4N5X9M93VnLXBp1jk/y1iffhDns0yd5KJUZXnhQSpwmHJ0Zns
ecyoXOBmTT9LbIc26uuLuSM3Kia+Si35iP8GOXQ0n3vs7DDwG8SiuxZqkRw1
G+BYkx/bWUdE4kluNmNcMKKtxVqgncsuhKFg+SOH59ESSfhhksaD6vjVGfaO
R3Wgio7n6QeLuP+Tfhwpj7zvoJJyE3KRzTHSQtN0UOf8Hl73yvuI/tOD3n2N
9lcPlP8E7vZW2LG6TB8Vbaie0HXqOMOrs9FOuo20GCXssSzNhkJKVd4/EusU
Ei1nMec2slAkTF9lmnNFsNIbqY0iqc9A9rDo9r7Ny6mYrUa/xp0S23exjm/i
KDQkeZNgmOymlpEXvYsvGNA3BTu8BuP34LkVFzyyrw51wKUMJSCl13WE9gHy
4mrAgEY/12PZN4+Eu72BvK6SNYmNt87fMG9IMVR1sFIggAM6biD3lvA7zgfy
3FZdMQpe9fT38uAHl5OqfqvqaqOlb5WI6a5v27uvzGcnGH07r8LJgVV4sJyQ
gLRy8MKOow1Rz/4KWClCc7gGW1wiKJxPwARbMCCovxr8xFt4kuMJYB75uOev
PbTDPraeh3RxWxrnHcZaTfo/ypLUhzJXBE3Vpt6bcMSp5Yf/7xbQUW5Cf65A
hifSMY5wojywXdaMKEw0UtIdcNlNlsolaysYkG5ex8kXnQJJX0hRQjp96Yb7
QoZGFb1KhLMze1s4lGh/oeBMUqTgdu1EIGpqJ/qBgmvblzq3C8XjseewJt2i
KZG27kTSoVJ26g6j0Z9W4mx7JIvJq6pO2GP3Fo/c8hKenAaGXm1kSuU99aYE
NGsIMzUik9YjYF6qq8WXaMeOebaniK3NHs30IYG8y3fueeMIdayPlBIxyzGb
S25CQR4j11GOkNIR5C+dxMVR9x8awaTsg6suokh2Y7b/lDBSw3QnWxQShA/J
dFcNAxr2xXXOl/J3YY5o3BfHVbT6lUO0kxk4PX0wiU/32X3xdQ+o1+lQ8VCr
+ifluaiNNbBOlEFNU4Hq89Ozpm4TZ17kjlPwWoOlugnbAoqS+12DlKzZEfmJ
QW4ysZENeH2ueDjonImJKH1/hIRUHtNl3Wvz0NWOwdB2RkBmaqKnO4D72GYG
DYxnaKg1gtNwYZFzpPejnBuFfOatXaqIYwbSVT/7K7OOwXrD4uPQhjtd6DrE
BRF+geRovQtmZcIqqZvy95S19Y3DzI9UfkhYhpt9dWyNOjjTi7N9BYkL/Jox
rGnGi7fGj6cCocU3HNe7E21epVPXkzUAPaFVxQ790AsrTDXOwAl+cz+n/9VM
IwX4dcUDB/Q6Z3ZfCZ9LJcJeNN+j9irqAUgDimoJoYAMvhK4A3RLQpVge933
FWwcXkF5sjk0y1LTMsi+oQYzLxXoeZY4XjQVl4hCWob8tgRJNsYJXciFezKv
57pG9kfVRzt9rmS8st+tPvaqDc1L/Wollw3VudchLoxaDiaK8N4a/aPSyabm
4V1AyHqul9gRsMk+VgqF0TopXoM8VTVYudmeeQXu9H1sdIbUymfyylaZ7b2W
Z2rBMoF/D/u+dXM+ArBk4MpiRKU/MD6RW5381GK/dFBDaXL1R9shrs1w4gEI
qk7RHYO+Ex3JDAY8ExKoL3OO2pDN8PVbsDM4ywI776gok8H+3fKLc7Yk1vAT
NIrV3OZWS5H/Z6JcJ39+illlVusnVVwmBLO8Z7rxJgqLQ/I7x8XXVHpuKQXH
4UYA27hW4yKMkGDxOf3/VP4OMhC+fFN9rTBAnnH9GbZYqgJg7sRnfdaDo4/m
0IMHVKaQ1neWnXixk4JdlY4aWYYhz9IEo8zQAceVvEWQvhTbRAB2/8aCPQ1f
qGToPhDcBTftdzTM2ZubUTg/kdWlJmOAkU84y/LkFC7IrF5nUpvqGnf+z0vu
0RuEUsCXAJT8z2uwm7FvWHtnqASZGgn/lb+EA30QlJ1513JZfZJ3vcZjh3Oz
QcJrLBTB/jPZPQB6xQxXlEcFa0PCsB9XIQJJRxmIpK/Y7E7ZRIiVQ53zfjjR
I9bSPdb4iNr830UQb7eTcoge10psCi3V3BcrDhcywscYralJYoCJOK1w8jVi
0qGVCoABQUOgLG6tmQ8WYa6hikOSiZsbt6w0krnzo4jywggUingBLTWP/j7O
aGiWQfF6/Nr4gwOlXC7MH5wBXWgnnz7Oo9CKpj3fcjCPfx2a+Rxg4DBQEFGg
NVS010qNz8+3CDGqkrLi6Ri4bkS04OH8sCCzzMkIaf/qeAyPC2c70PS7/jke
kQoSdDyTehmkhcLP4FCujaoTA4YZIuIX5bsirPKqc/16ZBKQKrHyPsvmRbKJ
RymndLowKZxB60q25Iw9wxlmk6WauTnobn90ioJQgfI62s5H3p1BowssFHzf
B0T9mIHZjV60akhT/12eRkC3ZuL9DfvsyxB7i6HjS3vfen9T+JoKXgOHgxwc
y/EY8NcpEIlsWZfd7WwGHS7mxLFxUHdt0bONxG2BiVaLuoN9a6K0D9qKSLoG
TpDMZaCX2xzKB3jvUom8lmfjTK8OpATefcDCnUcQTt+I4x6TXEVSwrtMI8Ya
m1imVh7tnv8iXtKUU2So1NIB++uTqzbUQf0rZgA0L3dIJ6TGFtDbvsP9fKBj
vwCfrA2rufYosvyxwXqYRHdXGF7Ux5UhLBwGtSEdc3AqRY9OU2vDLut/eVxx
F3Chkcgs1DXZg6KnvDsm402TBa0Fc4srRozGRQojaunmpjqqdtCFrnzAxI6F
b0aBqxSLa0PClY2rIwXZZusirytIVFYbnba6DNMtFotw/8e69ff43b5MAbgy
wvDc4qfkjOIcfw9coP0kOBPx1S0J14ZlGsUWBZxYdZLcpGEEbVW9lNgOwmsL
zrmJqdd7vDS8af6P7LMkuZrMremHwcQilAO2ppPGVpdNnOkSnCVy1Dt94djK
an+y7bXtwhHkcOcqqMVWXOLoaCHqrs9G4BoPAXn3tLIseIA6KlpiVRK7uATD
TRKhYIGR+SNUKnjw1jD2GRXbodyXucgYavkj4krD3S+RXd6z6GjwPXJwCRia
KQIZBHlDkkb3HZ1pq8yePhfKeLpcydd0iAoduuGVF+HDR1qNF5iZIrfpBccm
7QsJ4bJ3sXJNzubfvKREzFbofOvMvGofBTwIOKeiE9fJCBCSETXCBQ8FHAua
9wgFyZBKLfd7FBJIIli8Mgy+LRKz68jWtelXZsDjZcoJlvDi36on7FjESTqZ
J16XlPLS1/uxUOGPQCfZmNZqFIg/ucH3NzIKO6/3owr1RdclYR3DTJlpddNq
tbpYxUSdo87AG9m1/3r672KOUzdK/yqmZtgGrpNJXVP/rlFqmAQQHxQY4DvF
xAokWqT9mzLbae5OZElqOvFRPoDwacYumjcoUMYoGUZdjIz1LyK1uaVNr9kP
m/S7MZIZKlwk5Y1NovodXYWJdWOt7K8DjoLpSnJJgRCm2MXe594VCH+P7ubi
gc+b5n/8b6/2QPTA2c/ObXEEi2L+liUpSDMjM/WQCSQip9gnAYLKcrGvruv8
YqX+frbrDKCTrWZXN4AxQni2dqBxRSu2mTQBQ5KkiVrybTIeySbjasZlPpnB
tCohGU0TBANJMxWAQSnKzgSlCextZ0GpFpFnVcoh8Jyo8su26cbEvNMY42o/
lu37CIYxWi/5RDxbtB9vqz2IRH53vf3XoAFJQCUZFBzFFvKr4y49Pqks6Pnj
MmhcXyu42rd5leb8u3Fb7P+qT5ITi1P8v32XdHwg4q4l8Kb3Bvanfhx3Uwka
g3rCeBP4bC89cHwHiTfGeeug/BNVqz+mAxMwQLpYt8R32EgjvxkqklQ19ANY
anVZ9Tfweq4SXsi7C5NMbkt9M0gNK2yotsFugOrmt4mdlxROp/VpyGU0UWRu
MTEmG++1SgB4N4VF0zbusjHcCxAbm9bd7NOwepvIbCqUuv5EjSZFI2dIPjkT
4U66E6F4p8p4Vg2SwHqWY7AhqOOBc76W619qNM1jiNpyMRz4eMVAeqX4K1o7
vsAWD35T40nDeWSqT10hgAHnHwePxuDZQyTYnNnW7OX/NHh/9icgCG3+2To1
nvkVlNMmfsvCypocCopwzczv3ht7sYoYZ8xuVXfC6BJlQq+o0gUMkeTcwKWG
MLRc8iA0w/ncv29FckRejgZPrX1lvTP3xqZaVeoT2BSFo1vfq4lZ/0jYGM0o
04ueHdSaXB4aJuSCdwzYaassvyRM9fqopxY5J90djnYDIneFLuKehps2AKa2
MDfKO4SefDsDypzWOqv7LQFDHNVYgKj5rAmCE9myZhAFwDyKkrvN8BzYhkuj
8P4WkeiqIzelk/9+k5K2xKjyuvZiLWW5Hi4xsPzhFytrSjoOxYhUUq8x55hF
BQDMhKLlrv/Y3bIkwgBxZmwvxo/KlGD+jn0LHRxeJIh+pf8E8OQXIb+T72Qg
/rnbrhdrMnf7SAvAnmzHfMJ+oeFIeLz4K26T/HLk3LmF6DrgtVQ6LQ68taZ6
rm0RnnxPJhFpASSwXoMPXQ5lv7rRzGZ7BnM4+xgKQHaZA3mRdQuANdR1Xr9Y
GCCpetvQCIrKZr2zHEtGRfnRTUXRgmbsuYYTRmex6HU84tl/ETut4mwxYKu8
ysUchy9oO00kMwXunQEGHGyE4UeyBD04QewzvPb3s2Yy22xRruYFMjFGhje8
EZyEfoGhydmgr+Z8m3tR9nmo218t0XFZUxbXn3dEu1cD3ejaIvWk1og+8+ex
pfqVTCVYjnN0w5u7DjCEN4Zr61UmktqXD6FNqL647xwwvRaYSnubqh60hMbU
Hc1jJOnNcpUlJqXrTA9eEFxnwbmtEeNXVd+jhQleLblSl+liAS4Nchs3YEYP
9+AuarbUVLmuJkh44wFGSOjCZ59JnhikXdTPi4cME9giOttT8uuUGWY7F9sJ
OqExPw1QanG4mS7NwZc4pCtkAtBBRmG2IMIuGtw2S2Gdk/bzm/4DEXW8Wwxt
UrAyyD3yIjgbuqCHMtaex9ZjeYu83EMAFsZG+svVHwCRt+828DVQC/T1C1Ki
17i+1sfosyYU3eM4xdB/1ErRP+Biu/5tvwj4q5JOznILrh8OjqhaOCS/K08M
7EQ3Pcyz/XdqLH6C2WfXPbUGJhyJQcIn/U+GobQeds98/vC2ebHQKX8hOxQj
pAv2ANwyqB09OhBZAoP7O4s1mi4q4CpqsWddTpYV//07YYDjmLw5/FQtSrxY
XNeLNedPcr2dvo0J7iGY+JlHsXenmdqQqHzXVTYH5YXHqL3q6VYi3KZxA5tL
B1JNoVu5mkcr3+nWzIpZ2gWJaFXjejo1VNhEFczZhtgpH6vQ4kbjYCJXYC4e
9ejlvULxEsTZKgmAPnY4B9dPr6lx2P+MWRAZcSwXjgWY/w8lupwHt5llUvFS
eqw33XOk5A1vdYEMEXUv/jXB3mDGm97Zzk9FRe0KGjhXCn5SgwRrnHQ7yHfa
wCZKZ8qdD5/Tf3xNaA+VWOIzAutGaRbhVd0zkoBfBC3x+hQR32ovWrLSwBcc
q362YRYmmEPmToro0dFweipG+gbmSjFSQ+3NVOQb/RorUkevh1FH6HJ+LL7i
NgRuerDJumzXiYXPAFRojGQQdC8zBY2ApI8XFDImAEnSNZO1cbwIUdcHYT3J
bxwInNmSSbmmGRu/fKeVESOKn6n/g0S7Hw61USXVm6Mm+vzrQkZRBUIcg7RM
AYcuReRkx6Nec9LHGev00XXzBALpnHUhiLdWvuSKrNrWP0bMUlTt9vywvZmi
pzKLSHZxF/ilJabnEukwwkgWpwjLJq17Pm/76kXApnYu6n3ZL8XXBbpIuXcJ
UQ32acmLaOmwIYpimBQuPYQ4PtIAdPwIZgoD8q42GWNuPBQeyDZ412gKaqY9
dbP5KYevxGN3s1ylkQNjVH/TgOPqOxfYzJVbE4A9Aos+kKi5lMMX1jEpwENk
itMba0eWbQ0h7NoFlIQztqQjfvuYProq14vxJNb/wlIC6tnkEvtJaouinFD/
TbFoBJ32gmW8+gxdb6o8XGpgze3vscRKcQ49/F+6oB153YN8SHbxv0jvdN4O
5PDasN4KvYQvaTLtTeIi5PDw8/IU91OB6fEjnsNTYqefPw9dApBZoalG3YQC
EtIpSLlK8WbSqMWQjk27xo79ILLub+xoCf9ws4WGRy+MHJquYtC2V0MgbQ+D
PZbZfYxCnF4mM6fYecU4SDyq/ShfHVIKEactEYqPkj0lrAU48C4vzXh1dwZE
nuxM3CkgnCArZXU57A2wbD0sYLg7Xr96LP997DY6lIskuopaNWMxxWZQ9d89
O9QyOo5OsUM6G+PYvnNup3ABd9+0OgXkPiKL/49Sdxvkppe+nT8Dn+gSIW6n
YHCHK2SVqJ1KmM1BdFdL2PctFwqUxeK2se9QVBRMjpZnnI2fxiwfuqVju5Pr
N846D81+QJ2/GIJj6DyAht/Hv+rURms3L5DKE9fWogSx1y+upx3A1RovaSVb
EGJya0muhZJCxgG3EfFyxlYPVa9jDiPqLq+0QGVP7DtrO4aJ01CZLTTt3Uug
S2VSrT0QgEcWQ1FmLW9evloekhp/UT7ABDKt7WuTm+nJrb3NzORisvCsSzZ1
XS2fSGWS/pIOzQeZsDnR6n99djaGpC8si66lJRsfJ3inpahLTJYpPLs+ol+V
d1fnw99LomvCXSbGY4dAv8zhd+B2mof08Obduj25tvhbUur4e+QmbBfZrbgF
lNhGJQZUkrwR4bUKVDZAH52AuSQ/bVBr5f0awufACSYLZJh9O/So+vzItfUm
cMnclMp702/Sg3jMwnixpb6INTGj1+KH6umIVmZJR21dBvRfXSrvFRfmNL2S
pEmlXx2treVZt9Hnzipn/cY1c4eD9RWv03tdx6Bn+s2EFzLZxcpKWu0nagpT
JKnHBG5fSn8zWufTMFrabfQHpWdPKPkYu68pNMxSEEONWCQ8PdhDDxa/igEX
DbZuw4eteKzSg0kzeUj0zyGVKcokDuLROmdwDHu2EpHVyaPjNPDlllC+Rwlr
1hbINU7WZKdNEMIquuZe7pRpTZEhllpXAKLDTD/MIea76ahhD0KCi6C8EH2G
qjXJ26MaGb1YGAz6cYOqxgklzGndjWvgkr2b5ugThCFvgxqemQReho/7GcWK
y+VkZqzuuHB0fCCh5XHDnPdOuMZiTIeC2Jhuemkcz7eXfWwuKm2O4ArHiCyW
M+zOCJrCCU8AcmhKAXVW0YJsKgCXzt6Ese0EcWXqSoHwD3pBDh1ObNR+IaRF
q09US4G2ibsNzWDVqLvS7noKBjrU/ifUDGzR/VsHKs/rod5gtvoWBz1cSVrW
f1VbUt/G2EXE9NN4Dx/fNP1y0Y8ZwYOHbdq/3IshdYGAfbEzztYjhlR408Zn
q8zMMTmWmldDw0ZgR8N9vcQI1XgZ2oa8pKjNxrjGRatMZ9Zav2ZioxSLsEkj
HSRAg4yJkN8ZmwHFhKuEc6DM/Ozmm7+t/RSopU0HKFXJ0MteQ7/J4g6GukaI
2qZkBplES9lwv34cy+UOzTMWipBZXCPD1k4mjt4oS8LxUvH79+rPKAqu9LOE
EudDgm1eOi6mKBcAIdQorIyfPKvLVqMLL4+cvEGlHHT/DPmuqQpSgpyQ9GAG
Lxu3diIu5CZlsvluiqI1EUo7wRU4PKLIeK0cvBLSjQ8FgQFaojzCj4F85hoU
WsKAOOzY8d7cFLKRA85wIEcqbk8PpchNNHPTHZR4f27K+mLvaJKFgyIbk671
L+PCiKjhFDsgdVzM/kYr8tpfFhmBcjumw6e3diAto4XvgDUY9RFfTVM2Ws9v
iM+/KYQFH49pwvrgMySHX3ZZ9Wbb1Cu4D5pzCZ4ENN3Anpds+4e9Lu/oOSSs
H+fIDpdAXUD3Ot8Ive1CD2mW4OB202CGeJK0/VbpTQegQXfchoy+xMOdYlyS
+gk4dP6TO+Lir+XnAd22Ul6DlSAEUfbTzYXEIjs9Z5Jjxx2w7rTwxyrJCx7e
bIvZ0UI4T3Ys7mJy6tqgDdHfm30RHZkmxms7WnE8KWVf+wbaGJJFr/kNmwE9
YUi9SJXP32AZ6ug6dJ2HV3mzjy597Lmb

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wgPrtZ8FCfRMCPnqzG1pp9F53fNaRRLrkg6o8iyb5pQCdq73OLjN5/7wIxOv6ZJ6lZXM3W/LwTMZrhe9u9P7PHMBRs8gg9fHlIeZpnCap7u+VpQrnPkHswiGnC62aXQjHXkfhEO9aPUQR21UitLPH/KbqoyuxFPHjkIpImYogSPm5oOTlv+gOkHLIh2qVdhOULdYZFWtl2a6lX3ivVuG2SVYMuI7Vt0ZX+4Sq34uIPxXVqKz3AMKMTM8FLjbJshVC0KXzl6LSscjDsSUssye/J1bzlcszKfqN6ItepVMJbOhsW0NbUi3loNKHRpsVRjSVqubzwbGtgVr/O9wJjg8vmedeTn9hGleMFWct9yfdHTNleY/nFYAPaA8SVfMguo7OLkBhWTw0pq0tlcXn5O3HeydCB9H0zERSkU6U4IfafBhWm62IzMNmxLvcKoqwhptKtxv5Q+wwgZWyof4LMVmnahYGAZvLHJH8Egts4cTgzHaXStMXDMaZ35u5pTq8SrpwPzJx12YUYYvLopaAH0NWc8JuHenLsBNNoLCNjOAlJeGio3nMuptLxKFF+RBayeLvWqw9Fj9seGinBBzd0VbUp8dVmImxZ6uKMqGtKkQNKwfAZhZ3YcyEXpO9qUZsqbPWZLlvZUxRet1RZG0EHsUYyGulsYijXJNJRckmiEAkFQHZTXxlB+VkA8Zz9a8hZ8qTtNO28r0OxhUh1IJNP0M5tV6pXInqSzgx+TzIaB/NwTj39IQRkx2Ey8t1IcjGx5YlsE+WyckyS1Y6T746mH4e+w"
`endif