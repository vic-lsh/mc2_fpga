// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AQN2QyJRvZf73uAjHn0tPBvmDwv/lRuYLBqquhyMNJsPBjKlF39NDkea8yEv
hbkn1S6iMD/Jn+b/iaKXIZMb67VzGcQJSbn4NvjDeKlkh5vNgTqU+ao+ku9Z
6fNy4AxmG60XrC59LUlV8tNTOozn8cl1627K5ga7fL5XXH1cL1AHbSKgYrhl
i8sUBaDSICWnNwFEWfFi6CVubzTu5dz9eCHcJIzb6/w27avgcbU4oUuP39GW
D+DnMFf36O/6ae7EKojXg5wFwzju98U6QfVqvAX/F7FWlkbLgTxzN1josMR+
3BAhDV9VI188C8tb3DbamFrP3mBV+tU6TpOIxC8oLQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IGbNMvGG3GW7ltmMBytg2wn6GTBJ1IPnfgGgia3K0HWi4bU33svwr6suUymt
QOt6mFRNuM75t8EnUHQ++xEsTgSCIjeS08zlvXhN9AWod3UAZDxamhJ6U+j1
AGzSCVao7lxHxccaJJPrplf54wqiYQsdhRU+sBX4PLTMHfCBZxhnAtExGya7
6/0kqZG2PZuF/r8VAOPmlNXTP2yY8o5fB3qFizoV4Xspdgybj0//FJoIPSrk
7gxrmsqRzIS67tn0hpW2YEL/OPGRoVYJGIxgxTUxOhVXcYRCgG8txiymG7AR
b0mrSxm3e6ayeQd7TYfGY+KvcR7fganVMsbhoId79g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uBAwgizs28L5kbXCIo34gwIiyvMhW9eyqq0zckBbemLVqVtT+m2iLa0hR1Ir
7TeOGb9/0ZSoeIY672pMtp0z9EbGdKTyBdElOwH7Dmjj1TTNBaL4EbZja/I6
V/Sc49+hpFnicnX20J7bLxwCV2gQgPsfEEstosESFeCtaMxChp0oCCuk/qjX
TEJjLb+TtGtsKJmxGUbiPmiPGMGJVcNjnHTAvOApj8Kayd655cjK/2a6uShF
bpQ9WrxX4OTb9mAo+7SfIj/uw6HVmQj1LTPEVhQyQpX9sn8/o18E3/pJthqz
gIwaLi0a9hguwMyGIsN59Fk3XZCMEn3IxVBlTWTovQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Kn6gAQgbUQdjFE0moOEfjatYeYWOc3XkfK0Z1MoNfh20N3BA7mwTfqw/4+jf
ZjgbO7+DH0zYrVHKUpZBFzpkvfDhPLWjxL3QikEj7q8EnpEdIPBvgjjU83+U
5XWzlxZ7OrP0q0uWDZKQuqOMqAhkdQ1mKBNZkYHqVwP1BkWA5FOQwLrySijb
tDeWumlA2/zO2dk99V1HzHAYTRyh2XAnfdF3zMQgTq2Afayv4K4kvLrq94A9
f7f9MhDCiveFRxawjcKkilYSuIZP/K7EUOT7XvVVP3fJqKjCghPjvk4fImIp
1eiGKTKpcgVsnwgtFPCaceYpSmFXYK4osKaMMxqtjg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VwBT8lKnRG/feTSJY/cC5BtcE+YFMchNhWOilBdpWmGi09Ia+ibQJxCLnzJV
kNAhIn3oxd/zq2M4J/iI6l1ySG3pYo4zK64YQGxH0lGs3K/9Psfpl74mb9IB
x1e2Y1zTpJ2aehRylYW/Iw7uALEBarkZ3OGuVwDoiUwloQU2PyA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cxu6f5Kp0JLpgjb+S6N8COG0voPSbA2WO5fH1KuHTXYw6SQbCloDClKlFhgE
fOXqQYAFv+WkzdR2X0Hb7ORYM6tbVE+5ZxdBH1sFXyOofyQNIa3K2TrfrShU
fu0XeE8X8jYeKGBApG8wkLX7cjPqcNTb7BM+jTKKjQJ/sKG5eX5r1Tk0SOBL
jmyqkY5ClS37cX/HGXhz6dutRmZgB0883AFJcACiNTWk7ck2MBSnI7Qwcb7R
pT7b6KEQjJS+tgeZjd1XIP8hg4Umpo2zxX/+TefxvGjBAr07PLiRpiRBRLWw
h0vODwmEXizMD4D89u60iI4RrKWj1aQ4vf/cFnr8g7QGxSfFhK80k65zvZp1
X62KFNDwq0ow809NdA686Vtbts6SZ0CzyU7PgsEQpLhQkdzmxqVwxCiSrCUF
56OwU1FeSSPIwO8m61rl4rhl4P3fKhrg7UmJZ/qiXArD43/NOsPxUoOuT/IJ
xYLJHjePPGyEEwD8wkYnn1SUL7LQ/kM2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rCE1loRBfH0jqLGom6D9sDrZAgDZo9Iqx/XXo6m/Qmxow0MH9YAda3iUJF/K
7LBAULq+fkQ9mCVOu8+jRTf330d9E2g1UKZVs5EKXo6HIcE0ZnXsdiYEAjcQ
wGzqLQChzA9fYhdOmmQzYCQzXRTH86v+Uk8wvzsDhZqCJHjLgKQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EyzAE8ZP7V2dvv85RREro53j1Smtsuypj2aVMT8PEP8gi7iDntV8kb72k+QL
uV/O22EXN1k7G7DcrJj8UsamIc0iI8tCzlnTe43euO6CFz7I6A6EViEQqlFb
DtwZAIavjK5dXJ7QqyaxsMWhAhZC0X5yQKU2OnKYDliEh9pwlHc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13792)
`pragma protect data_block
DHDdm4gFSrsOGhMF8Jl4YNcmAV7nbi8vp2JotX3AQstv9Qtz6WgEjm1XLzn1
+86w7MVP3GgTXa/ZxIy7cGXfagbEdDEIOMzsOw5Men2HiRdifBN6Gv32gnWi
mX1QXAfsDXQ+/jpnDNhixpBnVcG1+2db5PW949CBEXplZdCsB+TplJM5oTvS
/k0qu//TjsJZ46QX/BJXsCOpMnaLtmXVgeczFDONB2krndyZsQO/XQTDED7v
2OH7rQ4FBZv4Fqd8RmXaLaKmD4fPB+r+JlP2MuE+c0o1vy2EvnOUyZDVXo9f
PKzA0jb1RKTO14EkEZlcssl7a1zC9zw+HRaionKWsAT/Og8TlARvzNsEDtFY
6ZWl1jwf/71XW8E+wcGHJhmfsu2qBWPnm9Ay8emayeuaJTOrwI886Knf2V7B
vlkF7iGAxJTFxdkoz+P9Hh4onf9euoB3lLYN/LRxtQWaOVB9TncqnNhBLAI8
Ww+iBi55H9fpgtGK9XLl3PY8N2lH9Ecn2m+hvfoPyu17QJDnITJnpz/OftEt
zw2a8FY3AAspe/LpbtdE9A08zyMSA4SuVYcCWVIdBwSQqYmaDA5ndSQ43vyn
v+jBxa3I6O2W6Rci482iqtjtnM45gMv7GFh+eiMUXhf+VhpCTrR7i8Vtoa9h
HqFE2ubVEstX2ke+tr+KlZL//wqcs0Vu6g1elIB+bzznZOYaAeOzUvAZO3yK
DtEnAtCR4uEE50dS8bOpHJhj+fkahhHhlfAX4fhjXkj8Aan1Q/taINCK+oZa
HO2kKu6YQlmSppWhLQ+OTgdos49664u/919Yx1wfcJPGFuh5VaEiqqhxZbun
amdGpWbMccfsGnW1wCAIbmmJBQCFcb/GzM+ujZbVwbwjG6Xpuh3GPCjF3uMl
1k5xXGfoJwWd8+lYUNhh7WiO/hLkYpYizWcwrPCAMsMj71SSC9QzzcLYEDqO
I8yEckJUXyg87D65umRmQhFshoRsCZnzeHDOg+gtwArQSiGNHb69gOuUXjny
A8WCElwoFHwKJ3y8fRsXLs2yPhZWj9hsMD3YYARIzjPxJxck6Jpw+ema7GVa
giQHB+hm60p2tcGsv2wFUUfzx0Ih1U6aa1SGv0A9Pg3ZdvcoCtnuDw65dXgA
IXMlWfL/lwdmMH7mZKRhV5emrEvhADOpIKu1xnDhu22xer6Bfk+WpAuo2taR
c7rA2D7auKJOA6D1fpp0lrjwW9Qr9XNia3PIvH64ut/Ipf1vjXGA8nqDLx6N
bKd7V9NqS48raKcTEIjQDCNnDNe96/+/1cwiaMjy8aJdcwWe+O+17r8fOEIk
TmGNtXuDIO5gur/4e6MIto19/22k91YU4LL1dq4clk0iaRc6C0AjW62tHRcD
LQJq04xpGSeBy6IY+INMIV/PodjVTXW42ZJ8Tspvj20HiM+mad+NBOL86HRg
YqqCT3ASPpb48FxeXZ4PpXnerUGXn28kv7MYWrNqCbQGoNQZ0gCuJ10vSlDI
NbiHSjDY6b56gUufEDS7eTBBRWKUmzMQyYi0O1TCRSTc4e7vWaaf2XgvLbMN
HDoP60PGJzqOXGtAYc24HVPwdotqmcf8ENzGtyRxuvndMP16JuufsmHC4/Zz
HLjVIlvSqGiftT5hBcCj35Bk4ZNb8ep5YRO50KGUbqYHbgMnZ7HkG8Ri+cAC
UoaMYEncEBmrVhod4Xv5yfa+EvRazZoLBc/wrHx86JCrqH68gTsN1wdlYHSs
K1pb8yLJRxNjTBa48uKAp8J91ahgqD449EEqhuJMDILyTc6rsMR8w2zWQQB2
m0cpOojcdrQr4mcaxODt2j2nXXfwPAZRyCMt/BjxizQZgx/y0jvO0OhAv8K9
u2wPk8HdF2ndSp4iNjWYwT53gdaCSLwrEtmPDhVMhH8z0Jbnph60l53mR+gF
IfME14vkVhcGQ8Sl/AARp8YjOvrYXy8fPTHGQ15BGfvEsblVR8fpT1/UtXLJ
pTYT6kHjpKvj8ngRgSg1Al8f2F5ktVkhf8j+aFYbRfI+Ydz8xDJHufmAblNN
OCsC9yVVWXjAgXU57OAzpJpFiw+itbnTzGTVzSOjZypqdkjLkloWn9OngGps
7hUysCkaGBZwBj5chNDHCKKFeBe433+kDlbunmDzuYAdTWJguJScybLTU6RN
1Xdqv8c36PgwAPV1awOzEZUE0QMzjUTHLya2DPVwrnmTP2I1meBe4UvCv5Hb
QIhWdu3U0figJiP1gkfPcIZRuLE7u/SWapoFY1vhCWunihEKYo5iGk+pFgIb
1AixKe9YPMaD1O6QUuVIHNHM3Wdk7qG5XpoMsJRuL7m8yi4qqhsEQxg6luZj
M87/erBmJqo3fofMJSG2RoxEioUmoZB7VxJmhvF9v+bcG56cIvGfZVdiOTqR
OsuHxE8V2A8aNpp6eG+7hxjENL0evqiETyEcaH/V+MJK/tSiaKHojQKfbA4e
eDS1nDH6JEwDRXQqV5MHBi9yfF9nsdzNEq88YdD6DQNFY1IkVgfmbcjbAX2P
6KrJ4JH65wGNI5x3vWwy1eui9m5TcuH3PLp0K6BZguT4YRuns7geNoZiQACU
+fAgk35iv7F7Lh9Uc+bJopddb/0e3FB3iOpoDMKUlzMhSBNEJku3xoSkK+zZ
6Yvh7uyZJimfwIpp+6A/9D6di6CM3gDAG6gp7XwXfGZW7Fqqv/O2Ioh9LrrR
l8nuT0DvLKLYM0AM4+tqbo6IaGoOWZfin/kdNn6j/kZ51CI9tG34kAI8VyHY
AHhcxl0+Z/E1x5p83M1f15CSLICO9UFv1s8bzeZJiD4zHS2EK2CwFNJgmzif
Ng3q+RghwF5krG1rfaUCtP2j4HMafERhuIDqYb0JqYDJM5FQ87bAwecVR1v0
5MeNpo9/6qD9ppQcmQnha4d/IoiuRwNqyBFm2guGi/jBm1rhiZxOw9t2n031
Ek4dnkGoVEkKJUEIj0ahXYN4Gx5cYFRK2IYFaYix9KfC7gEKpTlO4KU6GHe/
Zf/TuPQypLu3aQ9AvSscoP+e6L9GRX6KWrBHjslL+hljOZXNDl6tmzp5rHb6
5GnM52kTSt8dpD1agvYbOd0lcYjw9qRO3UnBo4Buume0bYfbs9P68uauU5EQ
btfSU2D8/8b75gv0Nbresp/eY3DltkyYFhHNfW8Cpv3JWVdHVkR1i86ZDqTd
6YLp2YpAIEG3YoB7pVmjB9cNEhfq1Hxl2AYkjT73RZAHRl1/FtbB2LLyNGip
vFxNy31ighD6saayONcd3HzP6e3MN6tqoeNIk4aQD1q2p7KFwEa7nI0gpcBg
UDyTAPBYC4si7pYaTgM2Mssg3vRly1mvaWUFiy2CUEwJVyfwAwqgwRek+Tdt
q2sQBhlUar9Wg8/ClCLhpA4MK/KmatrQm2d5D1+bQ0IRNZCApDGdaRh9fR1F
o5UdTNxLReA9Wj64kbjmi+AJ7YGmCjnZuz+yeWeLexs9pqifRW6Z9n1xHalI
TtgwgFE+n2jaoT+G9y1SnuIg4s1MwALAmLL2zS5Rc6A4d4jYSbQD6PFRiTN6
drJ4dkjCxQB1ZVXGwQE1M9Dqeb2QP9L5DcuDexkNrYy91DnUg5xSldYw2Yno
VCLE+xCLXX7UQQmBhIplJ0aCw3BtsDmFh7ca9zeDAWZ/4PEYhdY9PXFqPVdu
Z4dSqL1Zjf05r8IRjG7FghyqNgJ9oQK6OCNfpwrzmWr0JjXlQ846VAG94gX6
BVR6D8OoX4bTsSFibt23HjUJUkGz1+9+llklWch1hsGwG8I+y6ZB8CnIBKmm
Ctz/aHfIsKzOkYSpyCYLFUKrP/pZpEGi2nLDtet9ATQuDjmAV1IjeC8dkMVp
3pdYRWyDxSnNEYFAXJZeQp89M4iLYnqUiAKnUycRmAaVXRUXe3WXT+6krUVD
FOC76OHu+TH9qJgWXsCNI3XUR+CboEBXBC3mDh9M6IDjinDv+Q8vyAIlj13I
0IUdD3n1x1vjiCl9LDDGoc3aa5Zkfv7BiYhkk+Eq1CnQCn94+TFIRFbsZy/J
YdvX8ueJQL7c7Ex+X+RGoB6rUHPUUq1eiHm1LF8zmhIkoADFRnoU0Sj7RS3a
JDtzzkBocZ283u6ukSznkaqFKS5D4cJu9DuctCOChVs/nkMxRLkVKqle+iF+
E+LkVCojhS1Pj9l102R1PdFCCdZ8bAxGy7BiGvVG6TvnfnPBucT1bmIB1VOY
DuCpzuE2MnEs5/m1WZqjS6HVX2hZwFsl8Yzo1C+z5ShaqySlgQ3xH4H0CvvK
+8BXXGYhBKM7ZZWoS8+qpo3vJ/Y7B1A6oimSv+XCJw4eBqZx0YrPbb9bEzYm
MMwAq1RPi2cZSmyGbdo8Y4Z+tuuHF9bGYl3PrEbI9Ynz9eHJxq9RIMY9XJlR
N3AhUuav9Ig2Kat9Kft5T7+8U551SC86roAxqSjqZwdfcxOYMPDzNmIfKipj
WVaWDkKcNYA5wyWsaLfD5BFt8vyNPUah6+A3LXzz/pd52SlK7qxkuTkdyKsg
uzGihFeGNm+dtGCuKqkVmgmQn0tUTNBiWXmpck5sm5K3ySyps1KzAT4a1I1T
DroNx++IasslTTeCNuAodStyufJOckU9veb7lkuCqjvdNOh1+9BibRKeDqDo
L+6hjkjaz1MzhEV1bvoVL5JHsPGMONrG63WnW67/rj3KQH/8zPCx/zsa2nPg
U9M4dDhvevjJwP/MCfe+9HjKjUcpO/hLHbeMpL0a2S3SvPVzQUHxM5uq5V6j
86xeTYLmdp2ZZz2zeL1egtxfJNF1KZmc97ChNI6Sf/6taLK4axxzJTnBXHe/
ePlfBZFZl+KKI1mYW/BptxznadXaVwpx/apKoqEHI2yT8zU+lTfrNupEvZmm
TffmlKhBn+Ry8/9D8QZltehKlLqrEur2hcBcWdLu+GmJpibpiR6eLs5xjhkV
7ho/d01nPR2KJRmDRG3KaqeLAfmydb06lc6BifRNs1qvyjM2L5jkItemVS5c
T+hbLA51gb3V72c2rwUq7Pi0NeKbaYMe+UXwykQAEK4Jfmuqb4FH4rhcHNG0
TjRGDg/TmYUmT2TtIY64dlt+pFONOTuytJDT1MC71Ows5D0vJD8xLC4WSDmz
q1VxIwkST9ypPddaXn+RXK8TPh0YmfxhEMb8f65jZyCr4iXtDUVZVr0W8w7H
pxcZTtNXs1d1cFyfv5bhiszq5p6PySk94Y4hDLsxG+83fxXXuGIVAozK+rR7
r5oAhdTWWjJS0AuXJ68HQdQfWERa5Sr6Oh6+W9lmuE/Gbwq0/ensvKwFqiTQ
sRmShwVqhZwfey6G2WeoMH3RkRzQvW21VMDcCHZZbB2tPsG8qwgqg7orRLd3
9uMIz+zxlWyBcrCv5ImcUQlsBDvDkJDTIKKYLcXvNRqiMgC5MpLBECINs9m5
N5xwsAQegptCBaRXyYtvqf120qBfphJ8uTDy5scTqbtSN1DZEs0Ykx2G+fqt
wICEMYrr9m2b5ixtOW5Ce7ooJcZ3LzTI3n7VtPpqHm4K+rhZNfJOZtJ48Iru
dgiwQWHjZ2xoUXp0Uh1R/MR/VsR1YXEwPTte7jYA0G4Nn9gdn72LQCD/dety
c3yl3i+VSecmS2yoO5aL/W6+9y16R202nIrn7xHpYcm2J7BngkNUgwUpHTDK
0dm3CeqN0rNClJAZke/hC4IjEpW3oB/JyXvUlCeP0d7ANRJbWKf+ltZWsYIo
ytT+3AuJ0dVWPkive46NG43MU1e8oAVF/GUmyZWyouwroI7J7Fx5FZVpiItL
C/73ajz1zVKr84dqr9Ks6nXEFNUQRzUn7wQfLFZTzLHgLo8ZyVb/QIJHix10
L21ZrW4WZkjp3KmmyW8Ld3EgIK2pcUIJSx4qT6j9kSZln9k7tUJT5ZAfYlei
dwrWQTmYmVTLPYMA9Sc2Pq25F1E+tYdmTB280SCaMT+pLskU/t7fMseD2tL8
LyuW495ouiNj8c1TF/NMMyZP7NqAFtOqUQt9MIwsgCcu1Q/dXanezZYCXJKi
RPymc5IywEuEf2XZc4t/WyTzsdFT71qsztGjtW3i+039xcMapLKjE0j+Rh2q
+HAo33DKJNLsQha7rUcnjDL7aPUmTB1UmI0VXAkKRAZRBPBjU+iZoWgnZKYe
6wlIM9g2cgni7ORVMhPe7TLvPxjP3+MIsxJn4vE18bUWTFpnfuM7X5NJsOLh
dLdLcy6KdFmi+85cwDWX+ltUPBLcKtJ/M74M9Q6Jxll3uZb5i3ktiBiXRFLD
Pq0UL2+kpUomdVvDU2NRXN7F6mD0ignlC3PIYctJZToRHaAPWAmuf3MdTDy3
hh3/kMZLm5fdu0G3ZRe4BwQsopxZE3KGu1qKuZ1b+8T1USZJAeRjAZ8HYl78
UO2b2W56FIMRWbxxGQpmj8RhEuDSZGCFSnN4CsOLHqb0hUeoTt+ENFFA1mk2
0U+G/jyefVUbWt7EhbineRL8jPV5xmR9aVr2Oq14RWvx4lHjyRZ51pJUxQoz
cpofPyZ9f70tc6ePKRx7pvGDvL7bNFM4Dqhp4lRhIoveOSFTcODt61EvAzeS
qU71qxDigayzD0C35xcmWkIrXuCWDK+QhTj1bB3NvaD6qVScvLEsOi5+dBjo
LwVmiLBrt7GJ/M6Rzy6uIX76L5mKwzlTTlxt/dElJzvffaxmlEAZuMX0FOxE
CT8silfj9x1HqBkeJWQZXHrFd9/X+EdIINN3fiz1M62QBtTkLbXdBe8Kli53
B1+2uMv7QO5cVddugFddx7Tskk8D/noTUBFXHbj7sGS+xptUe2aEgxCmTcJs
YZ1D29gHHg+sV2KhKO+bwpgFIGxhlju6lwFrURMi58ZA/6VXvumHf+3gtUXC
xcYjFtYkStllGJ9ztvO70zk3i1NnsdMKx5CVal3EAjEnNMG1pf5zII+YhL2f
2iU/M0bokAU3Df7r/alayv38eiqsVTM4wCosRnIo4K1Pk6WVcYEALYSUOSCi
QnHq0keA8BLzGwf6ut93hdjiDoH22vgcYdTq3VgvnTsJ4EKaCnonSSWjEluz
oDz1ES419O+0oPBRlqaL9U2AEnoTIB8jWW0LZ5GbcKFMIz71WdU5ZVC1yxIs
ChcGmiVNPh9YNBfW4pSVIzw2zNBi+9H6coG4nL9Rgc2J5jt5QrxXdoYLvZZA
dLb3jhK3ZiY4kkZ/jV5zcCdfkSdmWbNw5JrVri9nRTGQLB4NMyy3LEQHjJCZ
O8zbfFtPwF897cEZfoQS0b9mrUY8wEzIFbiiDbqkHKSpSCKKdY8l4TWZB6Fb
NLUCDUlOosmGBBk3sLwzkBxxxYyqitpzuKSXCf9zv3qFXC8ZkwkZC6vBWEEn
TS2SJMOCv0TEHk1Fgi5bYg770JUcLLr4xr69t0wkZgDJeglhn4JXOHkkzMKM
rUNfMdmQQzZ/62kxL15r8xpG12QK+69VeGPn239xa8OPUa/3JrKPZfmmz6tr
39tUT0Ooe5HIc9bThmdctJp1bohLeQEstiv0n1oD3pLeONQgXO5XRtqE650J
O8cmRJYMAVaMkA9rjQNU/z26LQePP5ThnyMePdmQzUrr0qcn5ibyTE4Hw5qD
/5nLfq482ESNccjKd/t8qzLuOlIJli7ef1zePwzb9IT1ysTK/0gZQK3u74la
RCJ3meigTWOhPn3IWmE0eCibtfkYAf6u6la9pqYl/a5QlaWH5sGM4MFrusy2
4NUnVWJt2ax6NEhwTr5ncSF/GRTyWGacKjoLiyrhF4qfTJ4eelJ4GnU16vHR
mMxXwQmTKrKu702ywI2Jp7SzITazA9Inipu1I0bJo1fISWTMnb36ZC8vRPnv
017O75BBFwYGAcc1E3yY+PYZSgzhy28tl2wBWsIa3AcO/EorWHLSkD6NmhBO
FhNV99ExUfDvt5/myGacGsL8dEMA9ogJwchOYXYsPb3B9eORXEd6Dq1fQfh1
27eOSkaIgO2HNd6PCaO63j0nKnzHrQxZCKrd/IBSDBJHN74kecv9HXeQF/zM
LpHfSmI3PFBco9LDSIn/qJFBzAvcxB4JFUTNibxq+pK1j5bDfBl3ePjDWC9b
ASODMhmGAlUx/PxFvJ+Y6JHVH6xbOEaRxfraCZks4T40Ha2161B3XR+pjokS
MxvoCTBwx4wloaX3uR4AwIi8Tat6Yh/iJUocBWGDuHKlSwXDEXrLu0tDhDdq
tNIa8JIc8WbBWFa2Msb7RusSFykAut3/qv2SQ5SaP7m11vPvkrMoZIRzDFaF
uFzP+lO9i7h1IWpRbMTqA837XrAmxCIv9ZunJ5OqjFSo5iQNZ/iILkOnEw2o
Utrk/7zlFtJV1OK6tw9RGQQanrRW3eWZhouDKk07q6JLJsJkE1ilzc/+a9Ho
kkDw2o4mgHugGp1BZjVd2vY4f0Qg+BjyvaHTEwAZ8fhHmlvEimPic1xhjsjE
cfqAPSNwzwT1sbTtJTkn9J22ObKewM3q2oqJiyuP42i65sDeSi9rALoyyVbW
DMc4HGExcI66yVbu0/HKzn6ar0MmVa6JYIuBBvmwKizTvL/JXvHKL7AIXixT
WQyXYrPp2b+1r/3Wr0j50kcSiFgzOuTgHOH1GoHfEdXe8NpckRsW6G68NohS
kiMA9Kscv7vrxr3WiQxsz0bpDeC50Hxg3yOnfdjgM4CJmdpPqxn3fdHcSShy
qSVdUoA6ilvY9xFBOIl+MQftdat8JIyws9nBXBtcjeCu0DTi3fSInfQasL67
zg0pCyuUuVYV882LyzmRup3/Uv14htQxA528uRbuWyw75eKC/zUo7LznXvlY
JoJPuEiUBsrXXVZmW8xSIlp1iVW/IFvRiboXqNwpG6CRB8QOVM3KMJB1VM/j
p59p4oTG4Cm+x//PSxa1LJCyvH3iDN9rJ6kpl6sUgiPefohZE8mCSlW1UH/D
RfC/KXZM5eHOzHCsIqV1kaXdPNCpLrB91IZuQm6gt+EzvN2FX7KDejJKpTRU
oWQ1AQqczH4/4gwU7nA6T0h2nv4Fp0elSsHB4bE3mEnh568k7mYpBarLkxvA
dRFayHUJ4TvK3h//SJuhfEeupTexntOPlKDo9F0esTSmPz+TzPWTkPmFx5xV
+7QG1YhnwsqI2OQXtccG/LEXs1WscCqhE3K4JDrXH4slJyqEVzMrPb3+nP6g
c137adVRbQrb35KZn8Sc+r4/SZMh5loyZCrvQfDn+HrFzAgiZZEyK3Vevoov
pUe9joNLTPX4N/jayH3FV62MYiZr5sos/BwvIfuU/Fgq6qDgQEqjyLGcZ+eU
w7iMikwhG9n9CKaAR5EfH9+4OHfz627TfHzGwZ94jwBSFlY02QyVBn6AnvQ7
ZptoBaNa8ataKtgDRDIgYj1IaWivrF8bG03vyKcO1XAafqMZsRhNC81hDmwW
N4nuHNPK78PrvTd78jQffA4kTLK4k1vjM7IkjpcPhZkOk6NMBW3x5Og8zZOj
3CzXRvoY19QFjFQBbMlHrmDvvFBKJ5qHKuAovCLR/cljcV0WRw93ek4xtKFg
PFv5iaRQh/Ku12VDMqv/7A2lunMkI7Vxb1WoJ6/mzk3Xm+puzmZjVoBFI40b
XeBmlkKJ+ZsE4Y7KlvcljLpzTVHbr5+d/cSbXaizeEkGowj7ZnTXWEvFQGy9
wXPKQ95tvNWJfpePgnbWhu2k7CD9RxCsmf2NrT7RyBsq3ZrxqkeK3TwkIgvT
obzQx+ke1IULwMEzLvbL9KKVAeB+xS2xao6F9wprNCTzCFDdFKEROb8x8+jB
nRz+BYtrt/gN07s4PHYB33r2CJ1pPRIGB19V6K9djp44uwQpJmKyshoAJ4+z
RFwDXusIg/fvtcZgTsCj6HN+RuS1JSIMRB9Io6EHDc762xanJKPRC9Qp5cJx
6KcE8NjOhRMLSyySI2Bj8rGFrraFAikqz6ucJB2qCwhqEh3nWXkq0TbPWZP0
/4MTM04PvKfg/+aWxDg1j0nQ1b9VKiNNmTSKflC6CX2FCJm2lf7AGL9mlkoH
boYLWBJNkDEPAOkKxXtFqgiIDwp62YPx3NDhMhC4PQXJ0qqbhiPqgIx23mkj
gbdH68CUW/uv5JfaTW6P0UOPOGcSSBeeT0R3n5P+eSL4RsZYhwbp0oQ9F3wF
cwQWFV8V01F2nC9abyx7S/4la1PJc9owZWENf1pKckuE+iiS9ZlwGtEQj3Pn
hOQLJwxYuPf+3qtMLk8lEjUi34zUnzEsYlsWXIicNFsAhHNN9C4uLSXA9Cv6
BT+Et9DJLOPBahyoU/z7AMOaKn9qfZZ8emiVjm5ycSrJAqtshvirZaObAe3K
XKryjPoqj/UR33dsA4m/VMtf/80Ud/2qjsEuDWKEQ5Lq2qWklPT2w6WyS4iw
aqagx3bPap5sPA8L3qNT3gALCqyShCa0q01wbrKz0vGsGCruFYDPXZpOYYwA
7JHrgphiz3UubBeRvxZIM75fENvod++RlJJz5WreVLtykFoieCeTIqVRfIwF
F6w74NTgg2RPUuw30GzluDFuX5goUFmMI/A3XPcPLDv3yUtZnnZu0+t/41/Q
+O/YBcr8O+AWVt9/HTkftdDaoLITvJT+xCvdvNm8n1vFOqymaKu9Z4Vf/Tda
86YwrxffTsYimtb3wzk82xy2LrkaMiVXO4ZuYO0qq8nHm7t2Mz2IBc9Jy8lS
bhl/ZKQtNvmtVv5hQrXkToksSO+kphb6mz07Uv9wwQZX+WR3rac3624IEGIP
aEgB04LErXzPEpqafvrLyKjWYYdRqaktXiZWMn1vw6Wjn9o3XMKIqJaKfgOV
CkFc8CfPBbdf13h11DmUXx/YzNsTeQ1IZp6kooaPMBZ9MbWMtwxk0D7cg3g5
h7j0QE1fDnpi5OWbJ1IyY/NTWTZ+NEfJGU6K7wzCssB89KE0MqYYrGn1ujYI
zclAeeXYquTP6GYF/AKaIfv9NmQUINEuJOUo6eRS3H7FmDN38/L9xh8qFm+v
mNy90kOxIj6d8WnHTp1cWlWrkF5K7atAq2aKQVhSZ42Rlunvkz8EYCrdfm5s
1yYP8s1Fh9atzaqRWwPz0IxjraD/G1W8KWKxz7vI3ymANDEUNJKInS+u0H+0
8nutgU6VpokRiGmBEkRnL/15zujoq43LDmF7Fj9KwMpSN8hbmgKIeSLhea8v
F2G5WBYfLiHhBLp7ukU/j4ZYWu83gtAy9veOIkUjoL6lhXfOTWl0oE66570F
XFTNIoqAzfdYfZvii+a++1Ya9kf/WtmaERt044p2/lkjIcFonKe89C02aWcA
48DODn1BE2Nur4SCzD98antGXmiucxdRGAxAQdufVN6SDOnK/+HcWmyfsOI1
sWalbRrW7n9n7MCeqWoyYldoXePaqkidRC6FoC3stF4qgJNRzAUOmbdklhhn
XjbEqH+CjgU9ORJfJu3F8IW929d75et/wIy/bpHVAcz5QfIAiS1NZe/oXwzn
4hlkIyHXcY3lrLH7gCTNyz0hXH0dHYy2wIkpB5ucioe2umnwFd7xdfF3fG7C
//RqjnVVNDp7nADGSR6SxznvXqk+Sadvvl9tWz0kHL82Qv8oxWSzXQuZh0aK
va53BJOWmhKnE8vWfNoZeTUiLVft/WCvgXbWR1Zyxmiy7sDvmykTjF+v19BQ
SauJzxAh1mfRBPdli09w2ljcE9FTXloU4buBLnrlXTAYps5O175rwCAh8s7f
B2TTvvD3mzey+w372k5x/2+4ZRhlCX/Sr/B9ZCkv2XB+jRG31N2gG1YFUHTZ
6G3JJGmWmE705xaV0j27rmGk3CKaAq4vYlP1VMvF/+BFP8EeklJ50SL4r4JJ
i5AoCYvYxfh52kwXQYa3tFT7/F1wQZG7SSmM3ljJZhqs3z6ok02oKhUTAi0X
rd9/mIZVtY9T+LG+eVDj37toeJU2DDhRlSRG4GHo1thxf/TO6sIPYsedyAej
l3bQC7H/bLVCf3msBYXrwAxjVQx4dKdbKG5hvEQfv3ioWXPlInkHvDKpWZV0
Esh5+R7/hGtoGgmru+CpijjIoYLLEtHA3npuRCN+iQ0rTE4EkRa961AIoALn
68ZbHnpdSyERCww4r1xM+0hH+PD90/zW+MfovOc5bD6k3TGQ8fDu8uPIADfE
y4SqbZjgOhtgcY7qq5TEQnu4sv5WDpsJ0KZoxT+MbGHKqpW3ryN2IzHhQ1k/
caLUMnD33e53qmkxF9nU2ZQvIClu7oiJlKYKJgj1+a1yVbcGm70Ze/7mToCx
DWulygs0f49nhzj2poeddrmESF+qctvmhd7b8lU24hKIazm9Jf+YrsX0sKPH
0ZcLr+CiDUtnj2WycC/hjOkJwgEmBN7OiuKU8nz+Jr4Gl3dbUCUVFdfNCQk5
Nt8jOz2GDZ4v3oCty/rI2P+leVk1wYnXh7TcCTkH4o7GPOL1kmI9Orv+OdGP
8rZFSIASyozwWHwaieX7EXKcFrRSYua6ak4ZPrVHFB/jiEl6Qs9tFDYLW0+B
/HWstKDphrQ/X3hFjfGJtkwOxUEn+njqTktXqKO+esJaOxSBySFotMEJL74q
b7mmfrA9Mrj2XOFcrkgbvyf+NeKZhMg0+GH8VYQr05f/J6cioY5ZjLg15RoD
rhVQubVG/ZW4glFsmHDxX5xHC+oNkx+EXje/fSzfgVzv0URN5Ov9PWErjPKZ
mUs2G4+aR54XqtyMhmAbBpLZOXGi2rEnzyoKXkkGxiU0ymnkrdCARwzJKEoE
7Hw3XaZlE1CttyURmrG3/Zx3jp/GQEngO8RtunqOqd7YzJnGSOoaYYvVCrkd
OwhyqhUPNcvf0RHi7T4u+r1aJS14uj44us2YNAjpoh0wWdxTDXmPjKSJKLEZ
tPycSesiLBb7ByXM+E0gR1KpdHGaKTbNhNj5I2gJtrEbnEbN0hSKOMaUqRH5
31qSl2WtsW64k1DVp/iOwI13tHJ1V/a4H4PgbF659XOfqtODFveDU/KM2arQ
SV0hHWbp9I5ZVDefODDuxf+Esdq+HR1D5kaAyet24/hQoVpQseiQnQhwFRWB
xXRpk1CwGVmZ3fK27j97oMl7xo8bFE7gYRuDOKDxvpbpZIKqSTvrJIqeLKuw
Lm5lGt4ShZ5EnrN5gCFrN16UQYT5N/qLw22Fg9L4KLkVQqEKfWz/zgVu20ao
pLWIGJIkVDGMD4RXAxwN+oLPNIZhnbJgQeaINJlNikNP9iee67n7x1lgmDlN
AEFkDSrTy6rB0Anp5zvNkEBReNRF3rF46wkwy5bPeFVpaa6Okvdt/mrP7sx6
GRteu+GgfTybRx75GaJ6mzKC1kdSrrztod1fJCLbuLzK/kZbsEK6HUXep+gW
3hOtRShtaja8GurClz0Zziwfwclo3t88ZiBMY/MkoKmfLa/JzFUCOo5663dT
fnVAb6bLdk2CM/EB/tlCfEexPVtslwjNtJGoUozCYgSqGgf431p5ak5SEUwE
ZYnNyjzf6ulg22sLQ5xLjw7meGJ2BAPIO0CMEeCNCez50swBYLHjmKv5/rzQ
G4bci2Ydf8O5iI6bXyXEL10CBjQOSxJiwnvt9wkeh0rZofzoxV2iGL+M7Oue
y3VTH06sequguJ/QFCtX26ihHRw6eBvTJ0fRFoGG5HEriZBhUVRcnXcbAY1V
1k8WnpqWntK2VjUfveIdi9FDbaXJrqcsTfV35LNt9jMRAdasepqkdU++zKnc
f/KmRzLhVdcVQGIATftf+OuDVZITQexMhc7+6UT9O40GlhXXnpgQmvG4Qz8r
pN34gNgIAI4pyYcQJOdLv+KsU/V+rWulBixPm4erznXf0bs0WhUqaLR1DxCR
KYHrCsm0wEW82TU5pnp8yrJAxXkTzysKL05+P2g4zTijZaFLavDcwCHXiWTn
mpFnZXmVigvuGLWFeg8PsabZXr6RcQYMCR63/xGdeADPo4krO3SUOkmoP3OO
wk1moWCrdgLRu/A7XtElvYN+vbx76CNmG0ZpLG8kCk2VABO4XZK5vxMUNYhR
T7uoNux9zTWa21mSo9VRRpIr92FWmYo27pnW21eKIyZVjoIKzYhu5z40DYIV
aaMG5DgI2RJ8MVI9zswegdDyB0mOVz94X41TyIP/n8KAhfG9uxr2kT14J8Cp
UBy3Q6aUES+474YnQ6rdxy/O3J9D7jO1RCvzofyDz23iiLAH35K6pZ7bqj1C
BzFyhe19JDUHy3vrmGZSLyuPz4yN2FqBr9hchDG3WRCeo6IlzJdyQaTsm2NE
4n8kyAUdZGHUfxzfMmwbZYoYIG9nGX4o/qKc6QM6kiY8HUt64ghT/+Dmvw9y
GlSJzfjSTwWSHkkVE/+iu6xCq4uoayWKjzJBGkaEdpKGPb+0SDZRFaueLOZi
bF6p5Lm2ELeW/Z/5EVSXfICM7UZ/15o6x2CS32iCTxARfdwwzsO15lkO8PUc
bvsCOy9U9qdIpOtBlXZaoGrelyXSaAlJMm7vZJmvj6em8Xw9Qzeg3iWIm1Yi
6lxzDTp3hzsqL8f9fuH/f8jESqxCT6x0Z9P20EEDzWwbHyHDVeW6h4E1aqOw
jT54pBMzIAZvctAYQCZgrILs1slngbv0KcMSv29DbzxnS0hoNZVu1Tc64FOi
7TtiH0Rgq8xe3+FcGpHUKrxTGdP/Nk5wvLjO7Fq0FTfPuIwKtxi+gSaggh2P
cCBZ01u2EFSS2BvRDQzF7X2qbaNcIKNruWQiqIiSevbjLL1XFQ014grRv2sl
w3uvBM6cu91w2oFhWqIX1Hixh/41GrlYgy9pu42w6KgG0rqxPwbi83AyaA9M
+fg30Q1cZZoBdLUCr4RaMPyZkxOTdUAHxH4IPQ35gvjz4A3NCbfKWMC86s70
6j22d2JFotAwcQw6Q0eUvGg1q+2pvpwwU3i+Nn7mGAfD6B/pgZlQNSEK4kqY
yrWTANaJey5x5uslR1pK7YqZA2DMGHzitZuY4Bd7Ag+CDBi4q5FNb+Meh3ZA
BHbsyRNJ8GF+GiViI06AJHvT3hAI+9norI1DOUcICl546uVFSyBlICt38rXn
kRUmV719+sxlhKEWO4lBRn76jSk6+rme1Com2raaQiRvPcZET8Meo/w4kgY7
xuBino8C3tu2IIkW8tlwemKMRZAxg78CMSkcS3VRIa6/U1SvLkiAHNfteqQy
4yzkp0R6LRW8sNZ3n/jHmuonUy5uv30XUhglQgkldSd0wqmYM4TTpJ6AZpbb
k6LfbmM7bjCYbw7fupwytjozJmIEzgGjm8HPiruv3vCVKfGihIJb0PMZmm8M
d4gwTH5aabmKNyKfnd5MU7TKI/ScNzEcaaKh/pxqTpO2RM848V1hzAawAUe/
egHiRA3wMXtQs+MVy4h9BG8LIooLuIBFZ6NGhER2vzYS+83UWRESw9jfTLDz
3uMD03OGJxUzl7EB59qbAgCcjMGWI/1Vpk5U2LLhQuYP9pKFaZ/IKlkfMTzS
yf1TM0NX0tL1kGwY2H8ZzlMrMlfcWfVMZ1+V0CesoYjRed4xGJOv1xOWg6Om
Nx3BsW5C3zHFaK2xAjuUPU2P7+ThJnVa3MVSVCg7jvpf+4SFEi7N+0+WHloC
vIiFwgH1cOES4e8SeMOZd130pHzmYk1cd5sef73Af0y6MeIo7zfD0ym+vUIS
aOmPAiK+oA/DrmWUKl03swG788l8upFOGZmbXPIaLcHkGDwR+2VxXZhFxOyP
vUltUlWZT8Ac66ld13r25EsvNTKoBvQZKg92ijxSBh1oEKmH/3iFUEATGh1z
AZFW9FGmL6iEIBD51ApAEpV34wJkhp//bXbg0l93XXcl0JENdbG66Rja2Zw6
BvOOujQD1lWam9RXbP6emJJ4Pn2GiD2V8XsupcJMGOgRwf4osQT0YejgNEFX
4gNus7u6UC90/5SZtInRNzlfpSbVWJK5+tOt7T4C/tPIggYSVjZPVjgljcx3
jlL8Q80XduFs87ByKL5x1VKKkFLScan0wVTKgfh1N5QoTo/Z5LuEuT03N8T5
Frn+pEwZdL/lULJOby+LZx0xK8AR7CCHmfrl8jVEXsp4FZ47IzbEoGSNqdno
1EaxXpeS4YQQdyAHdnOMNw9GKZeatLgDiuJr89nSM3sBuB7EodMAfDRbSGtE
2/xrFJBoYaP8t6zK3ioKtkmJVHrgnS1sIA06xe5FAbyu7fPtLLJuIGSYRpMF
4Jz2/lxpZUPlYpif0vU2SmyiVD44D/ZLA8A72d43uiw6gyum1Adg/FdbsmDT
lZx6v9AjUfAlI8CIkIiEUIe7b/fqnMJ3G/mM4LzXPpFBN0GAt3ll0UeiOi9P
VARJ7ezPFlVi38nEGRNR3lMNpKtqlCte7Ga2o9dQD6QlKYcmlTVg+iCh6fBp
yDxhqb0yTgctGdT6BWR2wUG5G7XzVaJZDyFwhenO5BYSly0mqIyBKjpIwOuE
ek7I8cU+7Q1NLSmzIVlAOlyXmFUm1D1aVpmVNoZ+JlAajkxi3ufdSdCm2AH2
QQqllgJevEnbIi4ux4ERxslNBJxiTSB4hkUko7vDpHTJzfXZ6omEx9Axt++n
0AOtMl1jENu2AI2kFpOprWto5CTe2bn6QlwYDDsjJqJkQKXt4huxInoBT4Mi
p/lgWf6HlYgAmw4kIh6DXcKpqawXkyCAXTu22Gc/RfDhWhUIn/bJexnlfvKm
j6bXvsdvPfvS8sCFF+dGSzAfkT1GRA5EEars0BWCC+jFncFJS4Lx84jC+GYN
Svjh2jXsfnZ7Od9Wf7Og1OuNsBL2nx7pHpFfhy1f5t7GwIZMQFcm5fRESOd4
3nlOVjURChp0+IllBDElLmBRUzDqzPu5Nh+HJS9P19XMZV3JzyNl88Rd6uT4
s4D9J5RKX1k78cJvZ3+V0zzN7vUZT2YZThvKkw1uUzy2oQbNz0mL2TcXC86P
ydY4T3L33cUaMw29WIfxQAqt+mNmazUaLg+ucRvjp6BfDLt+K9QxoHTABPwq
9OTre3XUF7zyieVIlXIQzRm8arGAFCB1n3/Af/bT2Qtl4PPR2iKHxGdsLg2E
NHPX2darHhwEzgFml4crkRFI5htp3EEDcBDClINuMJF4YA4AETIZtFpaj42n
mHO5zSpVqZxSwQqNK51MKj1pU4cUJ3+Jl3ePsUamxo1sfIdKnpzCk36yayfp
UpH+3gzZ7NjyNJJBnrGG5BK5KMduZtQP8SefXApqGZMcsPqW635ZlCvfYfv/
pqVbGIMdPZB0FXzE7lG/bbr/ti/kaEEiyLStq//NJ56gs38PdnB1P4GelPzX
E/R+UJuJkxVDWYKbEi2sdkutpKubVEl12JKcbTh/SM8BabCRmN9pCDX9q+ki
Uw6JRH8Qavf3rMDUOJUhW/DJ8U8+652p3Pq2ZEzNflYF7Zp3F+T1rVzTZWWc
XiKHXMAj3WTofMBOesZa+z02RzOLAmUl5mfOVIilEJF2M0mhiCRsh1Z/Ze24
BfBX/d08VtqpCU8d9NphJtqMyBS7elUhr8oRupESrmZwvRovOnmp64VJC7z5
xjruG7/+CtZJfutmcJSX/2gGMkjRBtHuGnAcKkv1XOgQ/l+YFzshdS9fTohL
9pNrndIuvVvHPAdn03C3q+5wjh9HiV1Cgdq73xh597ecOyOnn14oLIXWVBTA
tluco3rIiVgyPbhHq5OHv5WAOJnFbRthGWJ6hNm+aHKPprfEdaZ602itfFuP
PdyssjRXjcCNPFlaJ8p8kYydE436kT6471VBX6w+DumOOLnXompvYyTV8TB3
GvhAyFEDHEWXDAejrvd9/DvS/Vp30Aumf7KCFWxqfKZNw4wwMXhaAeY6fUJk
X/BhZfaowoPaaGLiCipZZChF5AETXxEIWCydAI1RQz9j1Korlce2xo3XIId0
vma3mYFoSb584PTo0Jka7wHmudHrNZYZItqutR/zscCIymxENprttCEB6+SH
yYNOntv3N7N/Lcn6WtZa2714QCr/TyJQ9JkXngQfmSiWjvKUbUbB2FhPaUId
99n+BMRCCQWcWRxQ4WVo8tRXFh7wSAHgkZlL5OlgJOHMQ6TdtI5GjLa91SPT
U/T4fkIqjYED9ZtBP4HRgVJB3bv65WerMvh9tHuWhKcfnvElnKxNRR4V5ncB
yUXBrnRtPCEGkruUoJ5DvRZZOK8jv6JXtVkrC6FO6XMRZSvjUo3R+EuuwHyC
0VxOWVchggAb9fLZGLiUeuw9YaJGsfJYQUSCpdtuw+kezhuyXmPKOIwRlb76
kOX1XAUMLigNwABaG2r0jchTGCNdmSrlexiisSZlfjVx27P2gmBebx+p5uqE
3+LOiRnNzRc90iakOQBX17RT9tLijAX3RzizIqEII56RlWp8AdatgSAVIqtG
a5EXN8X3JoN1Md1V+yHsJIIhgEJfXkQPezmPUgDiEuEOpSvBiEEAFtxLl3kJ
D96OTV75im2juhRcPOvsNPr7ySE79UJRLI5s5RqFgbakO9UhrhBRjc3xS6N6
pi+YqseK+JYao2Z8Ki+O47dCz0qq6A==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EotmfKJtNbGf8C/IqDLAmcht0fDK3SsDpLKF/Sw3j/TPf5bW/sCo+DPo5eulatZuvuiFpFtcPFZ9MM+SRxMX7YRvn4dn0kPiZhC0GxDkDuB3Iwva3pDo4UyEv6GaJ8fckIiOshSFDtH3GTR/DpapPLuqzCqiKMAvHTeZNwIC9XpCyYXnw0DG0O73OFHz6N0IJbqV5LFmOF8wZwP6jDbBb2RbwPC34G/NeXRuPHQOzXeaVuPgD53v/WHUODzYfzqi5ry9oW5vKVobcKbCT0/MjK0fO5dZjrFREmN4/an2hM2h8FwzJwxp2kHDf/wc9WzlhgZj3Sg+1lvdZNDHS46hAjeY69nUi4t0lcjiZzoOKK2aGFsZi81KdyhiyvPm6hGjuCpNNxQ3nHAPJ9uOWqn5DLE2hhfnyX4Vuho77Z+3WA8uPOmLiwgbn61R+yIG40loss4xZkrkFcqg5hZBy+3MBrWXf/CvhI6NpFdrDDbQdzslNdd4jQ5ORGHcKSigJNarxIR5L84n9KxRgppBTC2w1X+LL36oj1EfJJSFx1vPDJhLMP5Ifbil+kosh5qL2Gu4/ISI15UsHRjfnm3/x7uwttl8wOm+vZY84oZZCRv7fRmpJPuQksoKc0q2DMlyeNSL7SRwaLwm9S+k9yuxWjCewoLGo7ZPRHeqHn4svfqLSU/eOIzR0QStpXq/n+zHtN0JJFJzRRrED76PRlGP1HqPxOr7c9mFPnyQMZ1oANiGWEIIT3AxaeO7394NAFtL32x1UXkPUAq3a7HEOWEx5Vs+lMa"
`endif