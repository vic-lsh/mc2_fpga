// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BgrrfXQgH5tkzL3rDm5+F0gYsr9PC4aPjXgMVwQnsyzVfAiQ72Ee6WKCqrAs
rxMSGBaaYzmznaSUbkuOQIEK4QFGCnrJG3WgGf6kHiOZsINDwtpXgVtuKxXE
RaeGdFN6ZjvoX1KuI5GOpkD2Q0mYLwag2vqx0XU2jLUfwQn1v7DVV2mvtXg9
jrcredEGxv8ODGcX74dhz+CM/uaidPl29KzajYfiLBsmzTJr33/gEULnsfwY
eTxKw2Mx2E2UfBmv8U8nHGDYegeAcWQNHrj9Qv+AR8XTZPBw8J9jF7iQafCH
+SsltB0oa8lDYE1urWpSogykhy11S/TGybL89H3M0Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bKxZlhLht0w2ASWDsSgmP8aFyGjpj0XlmUbuLjtAkhRN7TIdPqjAEAPhCZFg
ph6GlMOykp+smt9cdhGOWDNOnPXQ5Zg+NKVTT5+/dGoZBrNRXxOVcG+Me6gm
uyE0xoYDC8XNXC12PvU4RktadhEwkTuJ1sJH8oQRFp4njVuT61tT1HRea0gC
EUTgS3E44u/brqe8bPeXSTmOnxafe7yc0fLXomKmHVsFLhKspdvxZUUFNLPc
yGeN/1bJwZnR0DqWINPSb8Do/zCad1zoywEVGYLlsJvbWPH9n4bdvKiJUE1w
6okzz2fYq+AaakkYax2zm8QAzkD5hhOaJnABAMhGgA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gOQm3o/wY4JMzYM2/VuDJuzwThb+EOYOFKe+JLlQ30T3YvoGPlxK4NtTLqEI
bii6gQYFufgt2+0UvMe1TcxVpmVAp8s0WWfmVXV041p7fOExhrb5DOby5g2s
hWDoZNEv3oLhfY4fo65NcGzL31432tOjq/THJG4HugybyCj41/PUxU1awCk4
szTbMrLr0lLPr4OGU8N8IjNoUA5Xqm/AectcDa/z8muR/i4+T7lIfgm4u10D
1Ak39v93y1hU3Pt39aX4J28272KUPn5L//Vo0Hc82J8WnmGCPKOIepeO66Oe
LD19BVmoyxlzmQ1lM7BF02d0YYW5yJZ/FOPCHYFw6Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R4q1tWEQkIQwNH/aHFzTKLo9Z45pdGwkfHWTndh+bsDFmJkpO+fhHQjQIn2S
hDNi53Yth0KGEyq1ydavIJuClbmx3SGr21nuz3wikYvFBt7ZA7kHEvHyURPW
ggIB9SqJ3eBwwa9Sj3CaFGTSJMRN95edGze6Ha6Evy4qKKETo3wDsvcidzyB
HKPxL9SjEVb6qXZOtbA9Zf4C1RfQq7uddbCBKTvCbKCF25IxcIgydUskoL6P
UTBVbmeOcLcz5YSAoetnr4eqkLLdEYXrQcnBC1ewVh25VnIPx1P7NJx9v2iT
LBPlAsAOVraPwRrNwUEqcWSX8OqFZHCfRJ0KljJHyA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DzAY9x4JjUMrPZ0NQ39pQUiSnHbdae1LvOCR8GX1hliC5SX0CQ2pJr8P4vad
sttbfNi26BhqgwVcJWQ1XtHOfs+8xS38apI/Wt325UZvhni+k96JCIChebCx
SG5LZ7DqQqD3TikFs4D5Bm10ucHGLRm+jsBGZsU/P+y6ExZQTyI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FTn8lQoi8Ziu/F7JVJWfT9sBrqCMjS42omqvBMx3YdwpK3PWTl0BSA8clUvw
8VJ4lS0eOxdAQ6o9lGfDJwGI/V9rAQ0vXoXU94f4QQXHWidq8Rp6fLQiJR6Q
x7RbgPMPVXS/ErhpwPTql277SBSIqsuPEnS1GmtFtRjmmfo57YDJ4iHcRx+t
u56yF3RXoaiK5BqhegwVVOauBJ66bd0vA/KuAvsg/iElI3VakcGszvgRaqbN
dQrkrl3QrJlTgM+iiO4zrgAzd0apYOCCT8XgqtvJa9coBG+U2wgbwyMCrs5f
h8H5onwhTfjWeNOKX8g7I8E1nrdR29FABcgr+6rMWzlpV1zdQV+D/XXhdJkH
zSmRLJnqNGmR5RspdS9mE+tan1B8UEb9yO4OAgoHwPkOERNf83CGSyEt50o9
xVRJ5YpEa+cUnvYQYAOf8xQzkc7GMhiTKyjw7hU9GmAg/3rxBUd1wi+YZSTD
6tQ8rEk6jzxAUaH6ydTbavajBVACR2r6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BSK6iDxiz/xHSobOkPAtR/KD3H9lTSGNJfIJemroc28GqZljO7/57HpmCurD
e+5TGyUYtq9GCW2iUdFm4r4neVL9CfKcUtQ28YDhV2zD/sBBVw37ajEaidRX
JcFNK8fP8szn4CNzpsLsEHJpNDC9wGzB8mfqF9Nd82SOiS28+OU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ib8K640qZC6LcmYJfrWZzQzis1tkVO5bEmsS6EA2842PF8FFPqtb69DZXki2
aBAiHYKyKvyqtDMjmIhtq79FNzgzpk4tfjPPdIPj4xuoWMfDRrDBnwq2ssEE
HOVs6+ECMIcV6e4BWXVVz7JwqZ1noMmd7HAdfR2JpGNKlLmV3oM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1344)
`pragma protect data_block
qyvU0GuXq8lNZ/tF+YjSKyhjCLxX0eBgV3BtWkcWPCxD2PH+KJ5FQW2sz01e
d1GA35HbLbfSDAYB5dml3NS/Cy2LdZfGW/Gsbora9Fy0ZVMUYLxYvny+mTfY
t0ox4ExoifftPK4YXswrH9qVjQQuZ1TAHiQPGK+d6yqY6IxYgW84rIJ2zNjx
fKzGtLExsBqXYVcABq8kV4CEmsCWng6bEvM07iMH0FJIKReOP3Cyke9LM8zA
KZbo8D2RHAFxqkt3xCkVCPrwwXAGOQ791Fg5aDIT7zCuZc1xJsqDgmwpGKHN
JHWu1EEvTLW/Qz8VUIkfTRr1PAVCIiwRMXWRfZG6boP9LfWcl6GAZSMRwypg
wm4QFjdAQ+8juqvLb6edYYTnBaGmYGZjRqIoYDuIUz+YH59F5VHYRX4XDniY
+2OF2Nc+gXLHlaH+AtlK1aFp12o5jHhbsMDVZ7B32zxg8X6sZhBKU19OvFBz
zrBVNYe+WrEQqpRMo1yK3mrKJsgpT6n/WEHGJmwp/fETVsSkRuEPssHUQ+a8
doQsRW1f2tanw4i8HYaJX//4aiq7YEKVSyuO+FfHBP2H5pZIHsEgRzCrvJTb
JCEaUKe1kMsT+IS3txt0g+F0TBFQ6W9RQdRs/mEuCG4GldD5uA8C4Wmhj9Vl
YqjVtyjJy7OndzghrkLGw8/fMRpNkCTu3ZQOB7Lf7oLlAqwVxv6J7CaqP/Sl
fkpD3aIQzX6SpNFDh0fhZFjagUcDIdRlLJLZHOAj2W9ecjXhM9IhIjEBvy+W
hKfD3I9hLGCf9nILbxFGVeg3Mb2wQclQb18f2KYZBOrYy6/sOEfEa5I/bb7e
VO4fAodeU32eLu6L/6TcsH4S5Ecu3A5Vc1Z5dcVlzC+dSXQtfNVpzVmGxPgi
k1Mq/GLI/5so5UMA15i75amQc7mnKQ/MFLJsw7KVlDq+t3BPX0yHL0mYeTua
2USLOBPL0RVL9Gn7YupNXKAOWfB0Z1FNVgJy3hLFrUdGK3VCKoJBOSZW6TAA
19cewi4UNYGbkqjZjSEgBI0QjnOn1dLgeTMw4QwY5E3xIdyQgBwg1pIK3FdA
OkQJ6UbqClaEAlm0MalerVlDnd+pOJqjlgoGrANT/NWtYGaVJlVgHuz75ZEr
fNRSPa+qZgTq3lzuaXUMHAnTmxJ23z/hn6UzIm/Kgebcv+0KvjTyKXggex1A
XqgzPuKRlMUdh7zOgS/T8cYj+sb/d/OJjGuYbfANeTZTj572KoLfcueUfCux
gXoRUDjhsHYnxsu0agzwKqBum/YeMjMKJDK5NsLD2k1BO/MSHCTxbv2pbtNd
u0QICPY5bAjg3jWpWfAh+AKN1XeBx2FDWLOZy4XQJ3f2yuvs3uYXT+HhMTu0
pcc9vlV/PgCNVqX6BAY0I6VJXb4+oWWqRU7XqodcJMABICi4Lmbel4PjyByY
+tF4uPEG40kaRvb3bFYT4pRJ9906M2g31XGfc+ggiUICuXAmsq2joyNLlWEu
Hh9JA4IQcNiHQf1D6SqbUx/l6vSC7ahn6mHpZFtrLreWjaTVikm1gY41xeVB
/wVdyniON6QerSjxJldcCQ2aVfDuYPCyZjeWXXPU1cx49RZtd7Hj+H37PiQU
tS4PgoTdu8AhloY2DYXxVvYSR/1aoxJ1ZGJeowIgjkK3b+LbqGPyjLFFTmt9
51NfYq6YYZ1wlVS+nO9SDFNgM1W5Qyj2crtYXSsx4eCosvDG57h6f44K6A2J
D/RIDuk+ruIHhAQpLY50nu8D6FQUo0SFg8gmqPFTQRXtKCgTeNS9

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQozX1IV48geOs1ztMTFUyqI7KJlLZQn9s7xZolrYNH13AcUcj4i94p/SNNvWSvB974CGoR99dNN9D5l6SjS/wn7UD2w6kC38Uf1nt+cub2E+Yj3gr8lMcbZKlrmEUKEBcy5MxCpKcrjbQCRk3ljCzferrUNACnKr9jQMushsJWzwfnevIBx5QQr+Q4pliX2w6pLtdSqFsGzkKgfVwJU9aLcJIs4nDk78vPK6zo1DbaWt3eraBvoUjpFH1D2PpXcIYaODo/+acCoa293sDRb0dzEg/YqbotnTPZB32rbu/i03gnSkDvChmqgNfY+gmBGYaul5xGwQY1lL5QBr8CvInFZT1DmqoAzyszVX5wTOthIFaF5qIOMe2TrQMvt1k4Ga363sNAj7ruO1XSarA9w/xIl5CSw90xlItvbZmP9tpx7BqlCorNWESxkb7EEiM2/E/zYI5xlQ6pzNl1FIdnJhlocdagqSC/gxz9NI8Z9+u7FfpdFUtOwu8rYR+R8lW36cKPCXvjNNIuuNYW9V8/cuKFeknvHU4X6VXe2FsJb55ORPdMnTQKBLczufVYtlDl2a1md/G1zNdPPR61e0L60B7Cf9xQd5vHFJJmohMqJkDiRT3Ltyj0/RjDxECDPyKwwzeax5sPuuyvMvQLQ+4k41iy1nBLYDxtU9bR6ZEDwgz2n0OhFuo6kEuW96dEe7BTrm3fSWB1hm42k9HeR/PP0fo60HF2MfMvcld6pTzyxFjxraurDbLvJ9qRCKlaLj0GIbIOiE+HRAqctNF6hbbmgyQ1FZ"
`endif